-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2Tt+0l+DX+3ripY0To9ImItXoe/M3f6SnTnpu4vxtCt6SX+xeIoU/oaLkb2sT2iN
UglAwSNpy4bhEAbil9m9gWPBDHBLMgVIIWQrcET47VeIl90P/u0O7umM3TFVe8ic
nwHDp5TUdEJxZMiZk1DdG0YSUxGDlwFfhZN1ki2zx8M=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 19904)
`protect data_block
e7iWg6chxplIttLBKhUTFCr4B661JYGLpObYiTFG/Dyyrtyh8Nhj1BnkAKaEX9Fq
3OoyaTYgElCn5OLBv5mHjhUGAyR/mGepbdrtsBcj5yLdjIBCrzCGToNVszuuHI9k
8gP0UA8LPNyd1gTlUsTrZ0e/bILjXTl9nNxDugcB0y4sdGhU9G3gA+8WCbh1JJMN
JHer75wnDvpLlqovSrOIxdrrO3qIHh+THRNwv26yr00KEtEy1BhqzYvJBOOjrfRf
nRyy5g+z3ET75/UX6EBG2XN4nvtRNoX5SAiP8500Rb4Y3meKxrJnIwFKEE2H6ODq
lmVGIAM7yssnU1Gk/5poUz3SQDu3XNhbAfgCUOnq0SPTmuqhpxyV/qC0t2LAktEx
Oyj7t+XIEjqOFDx7uUERLQeeJfTAMRUsjXlNeDM64lidH0/PJCg3KEEobiJ2dpEH
ULzZ7HBtqGH5qrvEexo5n3RjYrDUk0vRGxIhllTnm5sYlGeWP4n7/XQk6g6OGnnB
owFsFycqHV5QV1ABvNKIrNxBlOZHSn+a7/apHhCrxrHlda5N5zu3V+Euxrex63xx
a/97DO2Q/zMg6RDQkvq1wrxGQtWe/A9OgrWHnqY+t8Y1HF1gV55A9xha6ls5VDuZ
a9Jadr2KGwwduGNK+98rXrWB+2i9+09JXBbWDmG4vBwPoy4bi94zDqW+nS9nd1H8
1D0obEDuECkQ7MnJvnWNrr9zEwXfAYGJfPgjIBwL8Drw06YOAeGUcSrLbSJeoPwA
iqUOPIc/ZLlW6ay9Yv8GRHAjOrl9jsd7pLolzVZ6TGTTVrBZ6HLjTVVR5iAS9rTL
9RR83X9BT/2bnwiUQEI3jWAo29ZIfax1IJr4+ZGjnrIXLGoDIutYY04ueNUETJf4
euLc422hZ/GntrhxGZL311BXCn5kR9WKU6MToKquQc28C6HOYwC6eV+mz2Uxto49
ZuHkSf29lPnnqW8M4Q6WfAWWVe/TLeJvl9OMXI5cCqJKyDT76wGFnX3qgkjgmlss
9sppaek0yaC6foJGPPPYEZRWAEHXAy6f6X/hqWQ5TJDGdIrov8dmoVADH38AE8II
CL3/pCeBRAteWoIkK5SH94A1aL0k3hXVGMFcixzT0vHUc7FgDBn0tPJ3tNN02mxK
n2N0JC7o9pvHOnmk3YESbwOZ0i4gLob26jTnUwZhYJiftoE2/qeYxXQzeHj6HXFL
+m3ON2BVr4MWGSunCzmvX+eSR8QyA9GQobKv+eaiuizR4S5fyWq2VCptxd8dnS4b
EX1tPez89y60QKKsw+iCIZwFIYZjOCiazbCwrwnmkgPLLrVbNMybLk783TzjouVb
Y5WGR7dTMQSIUVlcTNPjuPAM6vlh8TyIWkbcV4HTWFNFwW/yJ1LlCOsIdTBUYGyP
EoYkcuA1rLSE/+DF/OnTk/cq7ZX/heiIZeVyYXLACegoKSg08jrJhOVOmiM4gXhF
EO5CttnvTFNhJvtj+8z6TUHxzQDMeEl4TBLJCUE9ONaat9D11n25bKu8fv3s+n2v
meuKQx7fi5CPtOfPXc6DxjPXvazsK5BP/QOLMtmwmEizlWrIbjwUmBNSLsZITlVN
ug/wwkRKdhwphWusCfiT2qejR27CIkC4Vbs78LjuVwE8COzLHXm819WcKL5IG36A
mrYxrmF7qB9A4sws4t1aotBw43MOKY6VssPhIyXC/eIsuJMPeR4RdUMmHTfI4xif
vrA12dqsEw6VZqkzG0vskrUgBXKmW62+4dWgI5tKwYECve/iOPQx3SvM9FQxO3EJ
qNxNNH+XfyW74Ya6J3jVbl5E1x8RMdt1UXwaVKk9UKcrWJrNxFBdt+uNXqjsPRHU
gkq1nnu6yp1ctJPiwToU11srvPWRCIjfM0sAkVmpnzuyFsjh0uK2OFPrUp+QpMks
F5w1w9CwoLGsPzfeHXLHhuw1pKGAvvqH9nttUa0HJpom4iignjPcymo0JF3Fjpar
upzZgwC+8uOrmrxk+WfnEsv6kWjORk47A31OyMGeN7mhXH9yW1ZbFvty4418fjjq
8OpsZFBytu4BgKJxPTu0cihbvjVsAthmwuTlqH1c9fzAb2jOuxevZ8o6kxZ4rY+e
WSOLpStGqjN0zNEFVbn5bKJxdj4j2XMCUbsG0WueNb/yRO6rbJQQwbzlGLtS66/7
BSQRmOsob0SDrfrw5zxn0wbTGadP3qZoxYMMvA6ITYm/6AbVkKQfw2q9ei/EKlDA
ZS06tNx0AKe4YAPT0V95EgT+dfxoLox+LmIoJqDbF/0+8F9002d8MzZv6H85nW97
k/zt/dYjNIumA0v12z2GKCrFswXtceRHzvl0WisNK3E49pxKXkFSUqleLQ3w3MjM
khy2GSE22frI29CWICAGKqw5q8F1naoqU/yNqVAzM08uJFPJfaUpS7k1nQyQ8MZd
r2Y9OcYVx8Z0j4W2hnWSZHr3GOAbDWtfufsHk/E83kkFl/2CQFKr1lPTrpq25UIa
+5/eS5jtpsquKWuII8yDE7SSM3f9hnbdDNBOBWdDBUuig71s+Kagb8s9Iz8A3N83
ByEysHUMMXH8O7/GGFUpNXdNW8Px8hH50FqJoMvBqZ15uDX1hitG/w/zKTYB8Lmn
himriHTnww51VzzHVdrXmFaAQPi5i8rIppg0L3XuNzpZoo6oWIYE1rPkizoPJZcp
5ye8syT02NPBoEVdspZGZY6bkGEdlSP7lPejIrEbqhT7POek8PwlB5WXiy7coo+3
HVqQsh/POtgU26Eb+xqwCzxIV17zEGJMPLWEfMClexq5p8RWxZLPgjzzlzUkelQ9
Yc/B68AlpDGLw7IZIJZclP1tfwahWiBr8ciJikncGTsl1eOydhiYbaGLcHc/kwtu
cbTIe1cISKPvsDXCtDr+CCw/No67dwcfYUmxqodweNJiverC359zaNdtnTZQZUli
EWyY3T/+KLU5tL2Qp2C52gdAeYUxY2T9ck7/r0BoFmzP2sBYCKboOxNNtfQZ3mWD
8pPP5eSg/jBrdbzZ5HWULwpI5JywBSvqpA7DweGlrPqAmpExkpdzUaOCz9wl9Tlo
A3dy3X4/eUPTfeKOXri4+uqJfYR18FNuJTmoerKrfO+8PtO5+WR6vXzqPaCtdeu+
42sa797RAAUH2Txbrd7nT8jc2/PUmyOsWi9ZnJ45QXrXJf5sDxsacPwr7w9WZO8O
kQYOuR05woDdR6v/3/i629uUprWSQQxaMuZUvAaD15SQ55nkXQlixXKoP1oFcKQT
oIoEPoTQ5z3X5/0SiyOoQeJyMc6ctA6X9tgy5Of2MqS1od6XEf7MLc0gyCLKhXlz
O0Fp++7NwevzGa3zA7s97XxRxjd69mHJ8DXnD90G4FAageFgNrJ+kjddTAkjSeBK
1KJO6JSFG4pofiTeEADWeCnwPN8L/rd4nmhr04/nGi+rSmAbi04d6eTjmmg5bPs6
bwJN79K8/yJsHmqpUhBYeiMrO5CuzxVqRJG7/HP1JTcmkJ0g4VqR81f+QjTjQ2aE
ZlRio904bF/k/jKl7n8jC2ETvk9YRQnvUSGMX4bZAgpFx7eFS3HhgZjCxKyIpEQW
nFKsfYmjqImwAtqegd9rAviRk5vPP7vlIZE1nQR9K3clh5cSzmXD4lepOXdRqcXr
YovR3wq3Agz++20mlxWAJ1Iys9RJos0vLUISXZcAcvIbXNOSEMETRwTFuP9fw8IZ
sn8+EEq+UgCmjzuW6/XaAelN/zKGkvk5AwXdNSHJgAXNVC+6bkwi7oZIuSJpE6yN
AyuR6wo+v+0JQYmicmlhdQL8VdMwrr+M98dOq92mmI7O/+SopyWOb1P3gWcMZn2j
kWZOyIk3nJRmR84ROlpqOT0IP0AGtudmjcmMBS/KhIV4kcHM6bDLJaYQCIFxdmi2
N+dmDB6VLahhVQIAL1BXX0I/OobJcJoUxuJBUVNPZcZbpbF4OQVNIjqiMObArULn
vZgJ1Hap8rlev4WLb/h8CtnpBtFzjg8WecZx8XNYHtJfIp2zL27d7TKCRPrR+nlq
ZPm/2vrwU1nc3xfZqByWDVgGn2L0Q0PNsBGiaZ9YNlC2VqEz/8kQxIlToAFBEm5c
6il0Beorcdy5qCzxhFqKWLRSyctZUc/ENr9EN37/Xiin/SaXGRb5Y0Ocbn3rpDIR
QNSsJDu5Uar5pPBpTBvG8Xf7lqrpPk0Mmfgk+fkPgqJo/KA4TErru7q3cwd8NeGR
f078+AC8zFcM60UHAVzL1TM3ISUxZH0CMNPMXBqMg7Ss3cMwcsfXfonOwge/qVuG
ZA4RqqwqplOCaS+Md9d4Ykh0w3idFg4ixRCVxQ1wGNihgdXE3V1pv2IdXZEkr86O
e6M3lidc2SSFmHg//smp/x4hM2r/d6gLSNL2ENy0KVbF88rdO1FGGckGPDOPUtRo
qN9CexMnZPyiyoVucx+eZz2DkbKTXAC35GRiAlqpjI3a5IB9ysI9/720aFdF4ubN
upXReByM2Xef2S3fWnkxQm7hFbHXDoMpDBYeJP23Cl17gWUY+iQHH8xJFk93glVC
5ky4cjqEerF/YgP1YP22oH+lJ7Z34zlCra1ShKff+pGa9IinI/WKfRsCY9MOnC9D
WzB/Ql/PUnY5NSIzX2S/hR7i/Q+U+/9HtiUNhDazLzMbL8GIa9E0ZSdSKQA0M/Mh
IRTQesueqHAMiFufq5EHEYc8CnOpnZi6rzGl4Bggvm0UN/iSEkRk1bMniuV2MuH+
9Sf184z3RcJzjf5c1yqvh+xqrtAmqbe9Bah6M1GjVDchL7BbiqYiX6ihoJP804Em
vN/ZhizI1Tk+cNjMgh5ZhZ0JzUsljmS8+8NAOnRt/DlZBRzwFeGYwnWrBY+r+sIM
kRICgKqGuijEw2pLo14C6zUnKpxZWhHhwUWW3wYeoHQ/olKywqpkI9NBentAfSeJ
LS42lyGg2/fkP4T37po+vDQEqviz9cN0T+a9y4SXw4d1IA7ZdtQfybp7tCpUDShe
JVWZJA4XvybzfrWgtryy580QsEmB0riz6KUBviZov9tA1i7js4oP9PuKm30GjayC
I9sYNQ7vHvbMSv840wpV40kad5eIQVQ/X1F8+y+ACD0V5j/wJYs+Q6C6bF8FRNth
k8kJXZm2L81bFvaCupdG7kiT7FR2BlzmZUqdORIqz8agL/wgcvhvrZQooqwRJk16
VAHNKFsxUf1ZJv33yddrwwscisbR4h2CEMZSIY38r4yRzpxHIBHTcZWJb8LmMhgK
soHaAvbgy8KTj5JwY3E1QVPIahMxRPptXHwES6q5SsYaLgwm2NqwA3MzLFtpPCFH
LPOeiOyJ5QZNZFZjvB52eHyncdDRFldU5X4mM0KHYSaHh6vNBxhrWhUqx4bTLYNJ
deqnfeSkJjz2OD+1SFJTK+Ep8+UdsvWwHoWoK1wPYPJfMwxlzzlxsyyozSitj7+H
PmmYK2fe1mIufeCaMcaV6P75U5qS1MsQUX3E0JGMUcZSVVz7d6padzAMI6K1gH2H
nYxeBZaOJW6CcHLhMsDReWP2L6C8WX8FA44a8CqLbfb+bhGmPiht/XXlq8/hPJqE
4NlOI6IA5ZDWsD31Jr/OtT76Xot6LXiZOZ1ZoMFsyAS+W+i2u5rgs4/q+VGRI18S
QsMJxNVbL3UHZC1cEMWn9V/H/xUT4ooOzgaDJZjnvZCSU2+tefK7Yyan+jV+jYDX
rOJSl7FQZkO7FNEc+jzcYB3U6KFLfyzxW0HniiVTBhpLJ65VJ2dRyRGQZACxBsKJ
8mqC83SXmMHqRiDj5LvWkCBEtIyODeWoFFw7g88+CISktIsp2XsA5C/kR7cMIv6U
tC6wyHDFD1/STiFD5ZZbrPc3gQQO2IdLvbaMLvWVGK5Hv2fRUpq5yplckEqrYkky
IstGg9af6F791PrpVDBlhi4HjBNnPZvD98YllKB8ZssPPFm7ueDE5MKCWKdFPmzJ
h82BO7+NmseaxPqVpiuaNtAvl7UM+yAeYekhZYM0wPfXpIowNQdbCsSea4TNK5yO
W0Vr/s/BN5q45eonLVY67ehEsTqFA4kWU6q6GRstspA40BiOjvTYC59VzotgI4ur
uGAWpIysZGnQ/70uIDXbgflMOQNFQkl6XDdfCK14RZ1KQViXT1KK3TlQbnyDtl6j
k6kQkcj3TVCwxTRA/9jg0Co33Xj3k+yRwp4Q8V69EE4P5+HiusVbDS1hVfbguJNz
mZjnDW9bUItBf5btESTFRcQiUWBwoOAwNLrlrgKj0Lg+1eUAa6TI/LS9DnFVu0tS
mJryZ3WXstLOkQR5r1EUk6h4envwtimHToEKIBSR9TMyu/Dj2h8mxPM5ifHwUsaq
LRfYa1ayGFDsn63I3cEG1PR/Z0FvhUs+K2YZuQQ1fZGXlBRn/YlJR2n1c7yDzCHy
h18Eha/8iLrGZceEdg/CypuJaIw2M1sYTjbIvnLCgio2p7Z5Op0wmFVflFHR8uB6
elNvnYOrBKh4vqM9mfPVRuB1H2M5OpUT6nIHpQ+qo12K8lAUf0LpGCVJPZz7S4/4
924Uv04Xg1dYtUcSKqtnrrOejKV2e4wEm1NtC0AJa2NwxMmvHMudGYwyPdL04Tkp
a/NCOPfXk2X8wdxJZsNALgQNhWKGUzVjOa2B29IhtnDRMrtbbJPoYHDA5zhlPffD
fznd+HJb8ZV5Va3phR8cXqmMdEobNDmY4nJjqOM2I5exd4Bt80ly7f32Y4DnV7Yj
kibR4/rzVHRo6x5XlltPv8hw5VVNHxSUkxELM+qYnhCshtpGIy/+sJpb76WPmA/C
0qEa1JnlPcoerZM3tdk0YY+odhjjgHMC95M/PdOC1zvQP0AuYJj+gLecA7qSQoN1
KiZTM+cvAsJ6djPEZYQZHZO6TalCeZI3VAu9y9/OEUdSLBP8JNIteKr/y+h0ytB1
6J0OiWi4IsZ4A9n8FCxdeagjXuW8NULoA7n9/hkLEZPq48rMgmDLVXWeK99zw17F
6eqFCGiRwbwbIP1QnsiNl0ywxXahtodEui2VSKG7+KuM4FhajKOxwxudaWYBJ2Ct
d7ves2VGqXuN4ypsulzh9kCLHjCBpJxl52CaB5rmG++H8EZ7oPW5upGg3vKPY/t2
DuYsNKNn/uZepn4asS4s6u48Z6EI62yk8HDePVgxFAi1IW0Rl2V+FBVou4jHOBfW
f+4cm5FtJSn3hOzFkGwr4/8ZB2QRCodVtkPJzhkQX5SrZJfcV3e/RZ9HWqpmVxy9
vxA7y6+jNhMXv2MRwQDJ/zZxiKwTmG7Q+xmA0KpoFitZsMwpo07iPiz9tQzUVCOq
/l4dsp0BKkhWRUXjVT7a1zbH6bB3z8z2AF+nnSbqXySWa+L8YcjEHCYmC4Qn4J2/
m4jc0L8ei3f3tS0nizbopuzO0mL0DQCf6yYD1QXSZRRXuNwOlNus9bE/DGk9b4N9
zQ4Ug9csa4LsTh5gZE9pP2CGVj2iwGVGcJkv/I86V9MpYaUtmgaR2XGtYWvmvPqN
0dUqUhu/rOGXrWwIvSIp+CbOtAMYbK8TrtNWVkuMvl7POHDINcMdzRN33uwEH6Z8
mKSx0MViajgVC1UuiyRFfZTGlvCxfImoGe81Cyw7igkSkj5zs0gbMVDpRGQal31J
zxD82wHl0VquVsF8H7kGKggUM/Dm+EJpgYqLOgvkrb6qe6oBgdG2L0XJgtTQnR1m
thAOCijOANDchmD3W/Z8lA/vEwGFhV8rFWRNxsH8sFGkzchjqTIB6JHrbyP4FyGk
/vRIocamBHvwfjFocl/bVG0pR7np2HAbL75rqZ9FpzEppEH+43SbG3FX7ag3V7mY
SDAsxcUwzef8L+cKHx6IG0A52DNWRRVokfDyN6rV5OABt43FbgAeK6eMf/bH33nb
kZRop57qwy+83zvOxc20Gg/LUcEQSPMer47MyJJ+b04dwmIhD+69rLKgEJweP9fY
sEDBT+UontmNXaCqmOxsuDj4YZR4v2KeNVjl0VeUaTHoBJHbqFaEUMmW2jnaILG8
2UOrusuWYwdnQxn84Er886VMH1h15PAWPHtHya29EocBS0VFzbX5rc+OaeAPM+h2
tZPmi5SkKA+fpbda/7TbyunlpoFZVnkSldOy7GdE9x7KGN/Es37i/1gV7VI22deU
iuz1cnAcsXtv1lQEVyY9uvyKlIU59D5TbJun8PAX5Oi7RV52piIib8mqZ6rI4P2u
OrPh2kMaL568ExJsMPcAFtsFFJDRJYav51nsJrWLGlFMGX/7vzYDmjPkd/bu/vKx
s9Cc4tHN4xrZ2LyXG9/3+3XRtuY2d5be0mBue4qTPQA4Kd30/Mk6Lmdwzwb9rFDn
1rlEZawKzkJqOLUe32GZlI4CRNFhOG7jjsLlNjHRR9i5uXNjZTwfyuScWeAO118/
ClnAzbZBwKhaKdOBsa0miTvz+tu+ExY/1jwhhdwFNkyw8Jjf4NZwDY1/jTeT0MHf
XzbbQd4oHW5W7rOaqMJKNom/Y6BaYLgHceYn/RjAB8s005onyzjf2W3OcoyJA4Sl
YadEneuwD20yD4cfw31hmltHarCkyM4J5oL5zsU+QLLf+aS1Z044Aleh8M7ugk/B
4ykKr3ZJeYM9uYV/OmdH+Ym/C9JcXHrVWU9rhks/7iNJ31kL0xZWFi1u5go958mS
cpZl5nLbKoaTBE9ebBiwbmkbHEaHkyfpsPO9Z8pTPNEuvV+uXf8acWo2gAj/U/pj
da+t2bjSbfHS/FXjfrJpE1FXdoUdup/lostcx9OfLzEZ5TYxiuc/n2W1dntv75pH
3MYjDkZjBuB/nF4PHIia25Kdfbcyt8qRoNM9CF8X8bTpabTI8Wji8Lui9KkT5wt/
r60Nla6cjuRVYejSbz+nZsCYhky7V3jnaXD0Rj72T9Lus1f3XPAJRqFBzW/fTHxo
eHMOvATLX/Kaq93TTaKrxHD+zwuJwYhbZNwJ7Ilmg12ogegEj7s9yxwQFqhNj5bQ
w6zXEe/OprM+lzukMgxOVjqDsVoZMLsQGlhuxjehCn/ka71TuK6Uh3smGsogw2q1
btYPw6BUQzVomk9VzI1oQ147L6CMjob6mL/JlnW9y4H4geXnzXSQZqwN10hkBAw1
KM8O0Qw7tQ9rvPnESCz/rvzJVVrh4zoB39GNt/ESKGBBnGbMI1Q0TVvotbkVHALd
i/Iiomvwx45U+zN9vogUpTTJycCg/zhwSI3JQlaNX2Q+zYik7b7AEzUqnH0OHpEt
RmVT+MEG3BL4VApEaph1G9Rq5KUpk4M5+B3IjI6UuKRZIUWXGxmnD8uOfw6wS6fp
8EO+9oSkqkQtliPT2S5C5VwwQSZPW0Oy3Mgq73L7rrhC2MmHpk+/ycVGoLeaa2rR
XhW3eqzkHS3Mxfrev0Uv4cOQGMuSw+2UHbhMaQJXBQPyJLKJwXr8k2vxUOcxdqxL
wxR/T08dgcIzC7oxWPLTdfUnw6Fc99XIdeQPcbq/v3J6pLMzi/ZTwtQK9TmsDpz6
IH6zoZvbB3jXtB1HvbQPqGEfPGJyrSE0/Oy73c93X4sEyMJbGru25tHLdMotU9Kh
MzMOgioWyzjPqthh/zl+OeMqHYpijMmf/tjFWkumpR/2eiNaVxjYBHI2SZNdedlP
oeXrnsk+1j4dfR72W/qErrYY3k/TZgU2F46MsQ7iHztZ9GM0ANVyKGrpgmXTOIUg
jcstUeyw8TFGMkqev+D9MXf5PSyRzI3d6oLFUtrfMwWBK3SccCIdIK+zxa8Uk2Or
XhlDQDX0S23eUX7s/TMYLlMQQkXasHEhbxlAGEiI1f+NyVyH3sXCZB0bNAMjQix0
DgquRqgdTO8fF7BcIGKygkjpNLNNYrHcZxGeu5yDtce+KoUE1Omuuol1cru67Obq
4xWBnmMqw5/6zkz4pw7EWHEDFHgCpizpTK+fQD3xaZISEceGsU12T+XHiBbeMI37
urq3DwidE5vqzOpRTB1Tp29ArcmvG8fgpxtgf0Net7XaZZgsdzfLtUI/w6sFUu94
48XL06BkVtozCvrfVJGktWPIKISugvAzQFFqGIAIz/q7vfQQNLdeibj7pZcHIhPW
b0+Y9RjwUCxdGDbzv/KVF15fAtmIH2TiRUndTK7nLxSTy1OH1S6JGPNP8OyTPEay
ODB2P/o5jP17unZsPXv4BsEOiqtu1DDN3St7a7koO76Lv5xxtnARn0OjcuDvxY6e
PFWgTzsAvyzredrejIG1HTUhmL1Bno/hm/h09C8dFULk/zPVwHbRWdo+TcL0oG3l
UQvBtOiFg2Lt/LhjyiP/okiAUN3OKYS/Noh9ahEFne0rtiOhbZjgk58UYNVAs0YT
U8w7vq5/H3fAp9BaLDN8Wc1dUdV9OQyJqNsPcFQBKjcKgowtKH5lbTuURF4Cz4n1
JQnZzmgLWc8RSsgbEFfgCJShrljmV0WtVXvLvHpE95+6Pb4djmvIEbXYmilap2A2
ZPANcqWgEQm0G6ruiRoZyfq1yoHpvqZgtLx9mCPKpthllarZsPZemwLy0+IRDahy
32h7MzSfJ+WYQogDzHbQazjKI89geWyHITGqQIb2v88G1R7r6RUtX0qR4sR1XyiW
cBf2SeUStdwRzBUORU2ExUHW58Ie0n/dZOTYMafMDS/tkcUivmWskN7UQT3wKa+k
v22MeKKbgNDBnjtd69PRWArZIhUQkpoxgFoNNM+pZXa61vyCI6DTlhf/F0/oUJPm
mmM4/GQWvqTTJqwjQ/B1ODJDPfSAlnJ7f2jdPxnS2Ch1NNRRIyyYihT2qA60bPrE
rjcMMGE4C4LpO3R6JJoO7tXdwpgTyVRm6gzERgBnOrMPImaFF9sHOefY7lqDFOOF
zptxaZG1s2UXBYmnOBBirzDJN1hnlUu5IGBXFrgA/PJGhYG86Fk03ZueEpm4QZww
P5Z5KAZC9iDJ3Pt9xeo2yTbDC6c1kCEIK9s67rIl/LLUAmQ12lVMBNT5ZsS7+TVP
adeYo2/HsyizLDq+J+6ONzn1BohYnoUH1S2dbf+5RxfZOAwFd+XoKBcGTnr17Age
naNUQN08LSpUpOgIjuJfltFLAn2co2OoFUpVvsiRfVyu4ql1+O155MGE9YtiZiS5
Zg4RfbVd8qrHTJZ0QnENdOLAY2HD3lGQl79bHa/aEcVoZJutk3bWWpJNPwhLhH0z
LJZ5XkJBefWwsf7AQKMW+s5Ol8dAPUjN5Cw5xTNrqHR4HM8NrImyciCFQcNEaX1F
FI5bxE7rkvoc7VMdSG5TL9CA7h6cNiLZNaptcL2IfiPY+yZNTwy3+BMNuSjJM55g
TxtcWgVVV69KrKS8huQm15408wWlIbEktuFG4udBWIMgY9+rnrlmsxhTvmwNBds7
9Xuj5W4cD4qj3WhWvNxfF6/VAwTch6Fm9Cgs7vcSB3dTzbbWxO8+GfuZCtVxH3lk
LGtvAm9NA8lzA43Eu/ne1WGpg5H6utv8ZgKKPfPOaKY7NWR7CTb+GYUNHxc/rZmS
9bjnSveBqjuCCXb8T6co1vSKPAF0PzzpAXJy2Rp2opMQzId2FK29LTmGDp3FvJS+
WHZ0uwM4MzEAeDb8xQEFPiqIiwrmjacojzQjL5vxvjs6gaiqS214RZZ0atDyCkNG
10jPli2/ce3+zz4DhUC2y2EWDHPLy78zaHVL5GUT5ZAw4bY94StfLb+H5CwU7Puf
BBeGlAxJElA65S3kO59L42lU3opE7VdwNtpcNmQMjLhcaYHzPN0mUsOrJc4MS1lx
G2cqk7xm/KJBsyDW9HXjYGbL5McU6vnasnzOP12hzYIm9NTKux20A2IDvtzagri7
BmVGtcpYWX9KVQ32FLsVrm6X3S9zeVrB1x1VdOI1vmgSezGGLoriYiNVSa1CaY60
wKhKjG6yNavCzaxgp79m4A/SiRhde5GW8La9xCkJDkJBujesSn9/tsSfWepxdqsK
obnyodpibOixcbdEuVddxlMUF1hwiFTIbCURIpAVG9hFb8DySRLIdgcSO7zgnOXl
wNFiStLeyxP6hZHsQ/Vd8jeS/J0GY4Ck8pt6QgGMohO4B4OXFSoQJYEPCLgt/kBB
Su6lr7DcyHusI+UZ4OgAk+jLTuztQ7g6+mpMjxKHW3mxSmnN2lVzmmt/ZIs2x8Yn
Aw37q9LCRu93oykHwdvJpFEw6NuihJOHiII0EyHqrd1N0mbHgLZR3ogZW+9gPRnw
SSMx43zsRDDP/ny62SRf3TTHNwKB99HxtS1znShAneT1D2v9Y7Z+clGCAxuctgDa
iVw2yB3VaTurfcs7B3Ol/IL/j/B7hTNkOuwSJBRxT4i2ygepXxLY1NQGLkj2pAY7
WcOJ51Luh3Q7bzk5zHRZXhR6jftC2Ia7Gut1ENtaDPbAsXhXFPpysdPe8835C2yZ
AM+C5OjrN8lY5nIp+OjMlCJQ8boAF3HSLrVE4lC/iOGxXlFjzawb8NAWlca1/Gsj
Jd9Elqm1sVwQIG9Zexb/1UHeRMhAdGfynpswhaTQoLYulaWZyEcU8HdTXpHreK5d
XLW8d6V0Jhx1NohJmRoaWV85pKqDlfuupIZGH1g4f9HtY1jHCVfCYG66S228H8rO
hlao0K7NAFBV4Etn9fpbAaORtKsryuylSzy21vHOq9SM77M0ilg/UqTGS57DUsf7
3rI4XBbGIK1SpDVLRzCPF5MAyqmDJ41k9U/42IW19RXNxUYHrk3Df+u+IUnMEaw9
kW68yL/kQVL5109W8ASri9NyDDn45AIK49/4JMamR5ndQvK55JKqT/TbKEMPDQen
pBtBys+AdXT/cH4KSAkdgwKZ28ELQ8YUbC1/P5FJEAwYshXjHu99jZVwpiLYtgAU
A4ou2I9pL4gDW2n7aE4TUec9QR9l+yyTgumBilpZsj28URfZlGgZt1RuEr19Zs1a
8W9w29FlaxWxdq4bHB1swDmiTFT6q1R0oLYg5AKP2sSGjmgsxfozeC87/DB5lpl3
lL+zUvLL5FplhQ5xePOCrcx7mCyMwXApO1c/fk82lAabvzHdwD9YxbXogcyOUexI
QruVNU9bHgfDLonHiQ0QViBeWOXu7MKBGdM8iLOE3jfalvAIsUDH7BNesncDJCDg
IxtivhZBBXLlSjBLgWxPBUz4YRPBvUcj1C5PvWjtNrSwSEnHLwxxL2gLR8x/lnxM
41GnunOTZGkohc2X7Gb1gggyyKU/N+iW3Y5E4TY031n4OmhxiSINYORElb0UMD+4
L00qKEzCdoY8CfvsR9iZD/11fDh2wy8I0Qj86zq00P/5rCwfrIwDl9o0aFYba44n
8XsKCc+ed+hT6VxVS3nRiaKEgb+v6G+fbvzffyS/3H+EpsQGIXhea/n5fuXoYrXR
1KpCX6VGzuQHF74tPu5a5ldGlAzp6y1ktRZoY+jvvo7EZUaKvjJi7JAy1ktsQIOr
Tdf8ORPhLfIuxL0/hnXPiLPYqOOpD4HQ8LTuEOUn7k4ngwDOmthbvTc1AEcat0fi
Jed15ZZFDXf8FWB9dHnuKqaU8csCFsoGlDRaaMenlU3JBcrywEZ4U5BsRIg0nJJv
VvgfrpMcLetOir/kjKua6rF8Xgl1jeSUAppzxkGoQy+wCDm06jcpmyT4ijbDwW/0
GdnvLXsVVidVpMK+LIPCHPd5GlkZvz+7HX4sy4Wl4OZpOMq3CQx6X3CQDhysjXfv
mGHuiQ2eisq3fk5rOKsxanVQpSas+89SuUna2namhHumY8+cmAbqzXqVTUYd68H8
MzdJ4QyBVJMXz9gV7Jiw8Zjxu1ZK2fv84EO+GzwSwQE36jnDIntm/ryJlI5sWk/h
y82OOsP9HB+RImnxw5yrpK6/jzI80PEKuQW54CeFyYeP1VfbQovllNpoyaJbMbCK
EzGgXReG4IVjGNXM843CKxbPsdxmTAmSd6nr2nWkQdGjwSw5l+MBO8ysSTYb05c5
pscA7u4wFT43OoqlaDR6z7pLYKexsv2KZayE5ODeNmsOt/5OLX/96jIa4VnAcbHE
fMAmwd7w9PwL23l2phR++kye9w1KmqRInBYDECpQOAEs1LAIlkze+OaSkACAaAcw
Kst97vJt4dnQMfRODdrLEBFAyKULRXFowzAtUznzFM6qUjv5dduw+xAEUd7gaXid
9UtJNB6dOaf2iwIJsmsEaf5jEWzhP0XXgL07rovWE6KaoeAXpXHPsAEjlv0fny3d
m3mEVQklZ+/YbuZOmt8G6XGf+mUM7y2mAe9mh6R0BlElw5sus+i7e9GxyPiOnXVD
fAFceMBYrRXRAcGpUdG2gBhDFeexQ55CcKJGxeClOiZGkNrTwQLeYNw08GYhZQUk
jtUJXCOyO3Vby5fttSsBlhdd7Gs+0JoUsCcrofCrWKMrGc95NLLg2pZm8WjO9tjy
Iv7fbemF1lEFPq+pTcZb18WhXSXJlBukri+i9JoaBp302DLKWqfEUhZWzdGDpU84
lXC10kkLqXVPVhQKuLbUR68cBFYgGF+KwwpgDf8hW+9u6a/IHdWKGdjKIWmSxaTJ
vpL14P1FQNY2rDrRMFll7EvC5iV4h8OCDBSbkkoD+ZyekoE/ID6lgoTbMFxapWYa
r32SOX8p8nhiKRr2X2VM1CzplJhWwhMiogD33Uu8u5rr0FyrtxuEI8B8d5rfiBvd
Uowa6fRWlb+TBYIIkEoVHYliohb2SUg/yK0jZZRcVqlsJO4aKz5ig4fANmJTZx15
1OdHo352/PSrKm78t2R3Guclf4nXE9j8bMjpE+l4V/k7zUaf6/uZFs0j0rB6+m+C
NMA58/gLDj8bdJYT7Ouufu1ysk6QmcqI13BmLKFFYgGVmBt8ziHrUeH62kGydPLw
NcMjO2PnNuYssfmjsBt/V8DSVGP1s51UuH76KmvkGUVap0Kak6n683nEdvfThGdx
RvlvYSlEf1fPfgQUluBzESry5ZWPWr8jjFmQgGAMDm9ie4FJMvX84vM8BSMI1Dnk
aimWbfELOGcRnginUG1AHz/9sV2Zf9NihL7NqMKuhyuoCJgQdyvsp8f0guoo78HP
yiTn88RW3hS0/N2TIp0guI5eYYHVX9NJQiP2mLWJNL9otwLrwALHiEpxAaCGkl4i
SafoK1t47aybVChjQ7Yveb5JF2DKPfSH2hejnCmzmwfWqqK2clln3AZp40NKopTq
vSMp8zYExhRLCKKAfmazB7jo1Cm9tlr7W/LnmPpzTJdpAgUIaZewB3g3X+L8DIdp
sSTLel8I82LNvL5LFr4gRVlf1maWjBp2qR402W7BGBni+Rbd4ezioLVAaLdhacSP
EFqNihRvaewmAUiMwkz5EE2SmjG9S1QSFexDGeHDPGuFKWsNu9RmQXv+EBcr65q5
1lqoXHjGEBkhGMGjIH3+O45pHbKNlf/nBPiRzqT9vf84pZ9wvsP5U3zdimTjSwIb
1TZc2VENbRsowsi0kMOcidTqhz45L4AkYUpxcU9obYB80XygImEmT93DKV/AQM+S
CEKAWgHTWcNlyh2lR9QWn9WfrhpzfuXm/mOQXW5tMlMhSdU9QxihlokmhkY4L98l
jIvNQLTwvikiWuVXDaxUAfiXfM0Cq6GW75X+1VmPq8vdk5fGeBxFnmh/Hz2h3lPK
EZFNRd65vVyFU5rtTL3C77z2lDLQE4lFbXrVrkja0E1wzct/eiQ/MOL372INMVtO
D1Nd+LlEYA2k6Fs/lKiCp6qPgPc7a+SfBnO7OGwOuK+bAkCU136VGVAv6xBPAygO
A8mNCUujACKH+wN0OGaZrLK4jXp8ErGzPi6jL+tKgFNcwX17FC8TyJ3dZ4MzOOIH
32x6qmULf1Xb1kGZ5phiQ8rU5x7wyMEjmmuo4lbpZULfg4QTdKRMixzbFsZfD8a3
3IWwPtad6f6lSJwc2dn3pgCOPEFgE6+NoVUvLXgOgr04LNpoA+oKzaXCoKuhhLUx
xOaFw+8aJxvYisk9IvmQfJx5vaXOhyPIlkYR2RnnQyVKo7wqCXIh33ikp49vOX3+
d8JoWsyCqV5sdkZ8vItcHLQevQlRUyfqbPqRhhLaZ+Q5cKAMZ/7wq5vDi7iaHU8W
+P2In/VK4yAGsZ9A9tP87N4mFLadzYVFI33ZagQW6bme0UdCbqoZ1aIRXcSL/zcP
gDHRpJwQuOUyTdeWmKYLUhm6tROz+M9vrBW/DfwaVFVzb04uIiH+FpZIPxe3je+W
CoeDd8zicHba5qlQVNHAAkaoTPl32P1Ls0b03tV2J9ss0UOSeE8Fm1i0M1CGRt5G
veJRgPUqnvTveX1BMuIDf7d42UlAg75upbu8A8PSXY1DtOczLcAhu1EzfxrREj/f
O/qX3Df5wIkndlRAt3Iu8weBbVu+zVV5PxXloEipGk8Ah72E1oTbZm+VS5hpad+9
wTYUNP0jTMgF2ZyBdfnUt+Y+chDeRy3ZUniB5mEx6NwO9dZrLM+V/rG/g/1QtFyE
h1Cd2yHPAAfiyfeXkXuUZzPUFv3TSlCQd0kUsAiJoD9u73x6fdsdVWR26ah/NvKA
dLZ8j24U58f6rz53F7oe0cfZXYVwZL+sAB0v4h4lNti82DJ9+iVkWCwRC7PKyBVb
EH5oouc+35r+TDk6te/pMeb+nnReSONwmMLY9EJuGbl2WaDdezhlrKA3jQI4xQ9w
yzB/mF0GGNLdLKCjjFAADdDUoEb1psKC62ZyqVAyO1HNBIx+scdhrXPh933r4GDc
v3rm6gl0j4dPhYPSLxcxPlMLdBIeQoSd8VK62ftz/fcM+ihP4ObWhtzEK1ArYBRY
wsalG5qw3TSXGabndtTyBbfxZlaZJMcSxujqchHH3b005AEPOjfoZstbiWwoB/Ii
+s6eMCNtkeRNK1jvE1y5TcUiNgG9DddK/ipUq2o1LIXHFDTqZufRiT8e7iuyKZBg
la8Nvm0DG9qfjVkn0TDna52pjGFD8hmBuygBpW2XppOh4q2kEDNpi5EWN+lp8/7I
zDV1/3s6BHe3JWK0EGzdz2UipEjuqiQ9TZiWsMvLv4HAqweyITdhC6KGfW/e5N7r
Sxa0zZ6YrDK9EKK5hsUQZiwAeb5QzDOf6S7EtLe6j+ToXooOqDiRn60bZiaRIJ44
P9OCd2FLaPJ48DMzMvzCLbIc+8e535QQykOqEOL1Xgm9kjIArAGBvdVljYHZUaqP
sD14D+gptA/WdC/mYlT+EW4ZXFzJ+MMjHc0j5eUt3hVGuJFXag+v2bGNp1DLT5X7
4ol5bkwQQcQjclWv1q3K+ZulcMtRA/8oxner+GvcrQ77iQoxgAtTve2OCE4CxmBt
k69fk/i/U0J8nXBnCJr4pbWCzfiZAFpBv8HmkPUUcBDKkRfZw6VmydlOW/bCsz9R
9np/++pEmsafJjLCUkmm/p+34LU6A1AB98tzcdmFCW9CvWJOvizgvLdYVNI/I3xO
Fo2gQnb3jk72ukMVecbAgAyq5rlu62IGhkhiBwIuqx36HkFBvUGoNBAaNjDOmC0G
0bQklnKg2zBvbC909hki6PrxpaR6+8DrT+mTcVevMcmb15hc2bWIcyYY1qiQTnTt
t5Q/BOC+M/Tx0uTTYvBGjhTNRU5V3cPkRJ9aqhJA4Et5cHo558tHibFEnjqSvmFU
Yxl7WGWS+kwL9u6EJzKGdQuQWH38KZZ95b9H/mHogfrzTATIL3TPQ2aCvQx/l/mh
FVwR8v/p4QSptQHfhKP5jOKNvkMLK00YKw7EaQpskRFNg1vv6aEDf4souEJvFI5z
VSdGqJzit2pd6HjRv/u/HrTFETJmcn717cZJRwr3vbZoSa7SjsicZ3LfC8Sup8Xl
sTU2xRFqzO5BW5mMPhRcEA36Rd1j3oqAzKDxU27C2MZPItzc1VQPQwJ/at3AgCI2
BEhdm7aEEh4+di78Rp74Gato0twxDxuzTpWL50+iqUwlg/grtJNS9c0cwprC2vzx
hM+PHZ77JSkvcGXENCG7o7V/GNve8Dp3BhMtZlZJVLiTJJYXz2Bz3buqzfZBHCfF
p7LhG6B5NI7IW5cBNOMTq55vnNqDszj4MGT+Q6xlF1tWFEFf9IMEuSfqavLltupA
JrzqL5BePZeanPlbQ0mpHTFmTNGylE0mVWxWinm8IcIZQKjclwM9c4K9f2nFZRiL
PTPrU51ac9+tanbDeTxRgZJIbBBpf2FuPzhBd6PUcnilhPNp/a7LuCm8OJ0Nc8ML
9JCoKPdGFApPuC0XaRv3bQE+AYY4ByuFzvnXDJZFcHNLTqqn6s1H4Hd3PowiEFTZ
lIoIaUdmdA7LF2TH6/Kl9ofqHQe3ftROgHp9Byts66aoPNCnvhWqsKWocGykfwhs
hU5X8gdZbSnt4ZdovoM3ErPblQMiUac88BTbJ9oBuNySjwmgV6/OKkFA0zkUzBns
zSGg5ZJaGeHZvj6O+mqEyVXWveFgrygTkuN36z/4H3Wm6tcrD5AkgpycbpL3+Jga
1h+t06Mgs3N3eMi7LldyAYBmrK4h9fXYz7SUf/LyegWrtthaHwbwpzDOJVqRXuah
96O04En/WJfLzDeDcsHRP1y2MD7bDtt7SflQCuJtUY8dkKTpdKiJM1dWrcoFT4TX
9a48Gtasv8KXQ2zOaMcTpLOQGbV/xymV9FFu90dL40DQ/RVTPI1DvfLT8ZxniczP
k1kLvtup6mB5I74QC0Qsqe8KpJmOJFej40OENaemUw83EgjICezCXLezLx14naoa
Doeuh/ZH2Wk0bjiKzRAlxD/2WOq8iNX/+85fiO6v2PX2SCRwRU2rT55wJjL2Rnj/
S2ceIsa4oRFZAP8aLTQvvgsnnnvl3I7W63jWPeoxjcuiMbI8YUuwHfaST+W/tyq7
vHsKojwlBzMfYlUWMesDkIvkL9xBpgCUkAt1zj6fdwux1TkunYTKkKhUx9OZ7icB
hM9gkz3UZa4L1zpHpkrHBwxnaVPW5+koL7FdX3f6qo4RdGEXSnSdwCNLp8YG9E6f
b4IrTpfec+gt7v7Vi1OYIxo1x6MlFmBAU9DEpTrQ+RE1HGgocBcS+uZeoaTvVNVs
38KKejnxJC5ZJw2nFbK1b/7dXdlFfDrY0us4xyGGP44Vsk0ykmEF7lickeq469xO
ftFptP+YSIkZPfLl08OCgMvsSO6GMsnr7Obc+XRtcqVDZF5/uKFuR9yloOYhwiMR
NNs/jFSAXkLAps/+9eZyV7d6KPQT8Wjm7iSCtQ3exq0tRqsx0KQQeGUyM/CKMZXp
OwO9o4nFFSyepTsSjd/TQQ0WJ0JzSy2qHCXJS5jKPRLyBgPw+nB2FCw+01DgnDCE
SFrO2DWkPUJW8APRs02nmuwRCnW9VaxZL0iBgFfNNRMXboeA/cbvz710J7g7YBHg
F63jQBHnH7XboBfqWrf26jcx51aR6nInVg/8RL8iA1994SnJrgNlgp+kCs+DFQ3q
5ecmr1CbxisgZCGsHog+R1Kcmd845WaX6MUP8b56v3H2l21WgeuNJEgUCIQHhT9l
ncwyni3AB69kEsbE9yc/nzkWv7NoFyVWP/bDqBrG98lo10frjZVsbJ6G1Ab5ZLVW
L3HEC4vwV7T1qqy5HhkaLgOe+3x2iLJMB2hg1bbnpjB1oXuqsGu90wuitzJmSpeD
/wpegOcQ/ZklD6mQ3BgxgNrfGazt2zksXX2sy7oX0IZHg8H3n6RU/it3roWK3uWa
aOrhpNPgZH5DlCZ7X9AQmaWLnpBEFDImMrxLATblCMTKq/BeL4yraLUYjfbJd1PJ
MvOF7xuXcsX/Zw8A4wrwJ5UiwuoSZ9Z5Fd/Jbi3PnhuwNTIuIIetBWVe2YnNbMNp
O3gikCQrjLQ5W2jjud7Y2uIYf4SBxDCGrV+MolpDZ8lSFlD5O2uYDZ+QLJvXcrID
TLz5Ur9TtpxMO6w48/9xpb6ABOsyb1hGEcNEb77CNdpPVfeF4rGvMdSFl5ECfUOQ
fSxf0ZjIhGfPZOmIGbRb0XN4oP+o0dKSyFMpy8NxfrXf9L4xv7hFo/q2zqHh3m2w
qW3Q4AFEsqD6J5mBmCHjJWHITHmsudpLUI8+T08/j7cAsZJxie9Z/tf0wojzEf9T
KncZXpxwBpaz2Io8h0lSvsiVag8L0+jKHIbUXb57RjPLDL7wA/YB2dY10/Qv8/gQ
EF0r0ppMTblT5b7rBdcIfD3oRSAahllSqeicc72T2eziYvZs8s/xl31fqfaJwMBI
GcdnDt3gELalc/GL/M9O4qz7PfG7FNpubqe19mnONI04SR3z3qujcTIrRUj0g7ti
yE6spisluG3AUF3DMbgucFSY5ucMF7VNNiYUcoXI1vI7qx6tgFJjp4hee+vAVcRM
EQFreLcWCr/8IjvfwmkdleP7gwYy/I/N0cPojrIYuRffdHdnM5Uh+qp2yG3XjWLo
T0v/cndOI43mO65P41Fyw6cBmQF+93jFs6dvQcuQzZzf64Hvm01aOlsUCh/kt0NE
1gHBrdQoKyHrhnjwC/WIfPD5g1mTEbDKGnzWghM+teKVimWnAg/CUrYjQ456GpIv
dNGhn0ZKHKlePYq31gWNh3jGQUKhIwejT6Ftt/IW19wW0PZSHVenR64gdhPr+ahE
qLdVMcYL4rKPpeMxhgU6lKdyTw6sRFf8va1T7619MdcwEDkY2Z1T5s+TCJ46gzQ4
eJqKKfbpjSBcqxFV2O/WmdpV71qCBC6dNwKjiP6xXZOSP4MmXuLjIvW5IypF48lj
QyDP3uxigbwRDVuFNb4dXSTRJ+9yKLdp/w8LKVSLimta+uvrzrJ2okP0TRG0Gx6E
CeHl2JP8Z2RddesYh33IsBQmIKB7Q124/GvlVa7kCyJCZs5doUU+YHSK/PccjJCX
euoliaBJX21K+Y/QW5EW3Z545n9NjimzsSFMUfgK5HtMLJz0/XoaXTdYNqiI6uc5
yHi1VSOYsjDZT7JjErZQx7K16I3fIyYXrOa3k4Xgd18H7ZSF1TDyP4IKVF9C21ku
2zwQQJjwt5mOIqt/D4gYsXSnV3n9LPTSa0zkKcghd1sHhMsgyLENum+g8lblCpLc
STjRXq8QN7MGgHVrZu0nqzQu/U8ox82xxPzM1z+lWQAfXA9XThcnPwmE+PmYH1hB
C/Y8rKk+o74hNzSGbRYHnLKYZyglIZV0sWYH00wZ43Prg47ftgH+huAm5tryKxtr
qtijuFRxRRCZTbsNym1hC9HTfH079mPfkOX7agsGSJ05vNgtp3gU+5FNOEZ0iDTu
USbiLTvVewthg2TWWgBsK9dIqfkDGVyaJd+IpXVBEIzLJs46ti+kjT/7f+NAf7hK
QKfDfFUn+xhp/Ru77Ww9oLI9wCe406myV9+c+WsDDIk1FC4oPqYIH9xHZC149Agj
OlpoBfllfWIH9OGrbiE+dTsLSzuF4nopzxq2OaJu7t0icAqQ9XtdDFeiIt10VYMO
BVb36bl8gYJ899+OzTxnOC01ERfvFwm+3LS2HurltACNYk1fOIuCOlFqz8ySI6Cb
W/pL3uTJQIoLlN3UV9+qijIjp9q+Ls6tRnYGgFITxzPNQuZ3TtndaamsHXAuipgc
sFpTNNH9T6xGP7qd2FfnfVmbf+bFZ1f54S+d8+whe61YJMJ/+Kig1fhc36+EVm3t
gLwh+E5adpef5i1sVLz3vs1/imiB3mlfq3ME1TwRuC4QRCYSbHDdERPTQ39AZL4d
piG6XYaxeC5Jtskk0v45j2WU0aWEp+9EjPxF97P8fzf2o6kaMsCxARRweMw7zeQm
OP7KpVXgSa5oINH/NUe98khl17fqa5Hwu09okaeTZtPgKQgcrhIztHu0Zq/IABN0
Zz8PmtRs3vAJm7ZSaHtDm986jH4dMNel57qaY1YkDjUCq70wBh2GrRg7xRtrBvAI
FZGWstJDkc0cIBQLTJF8Lfnc6/kxWxEZ1ptrZtqJP5vgPnctHjBdOqFft9HUzWmb
DLiOB/GwES1uBOCJj0aDUFmlx80TwWDbbXeLVC1gb7Fpc29KSUzZDzN9uhyakYIr
5lwyVsAgGIZz6jA766S8moNAn834vB5HNz7Glg4eiVaZiaZRCt0w6AIk9pmVhgz+
SHO1EtmqOHq0UiibryOSl8nqr8LPVT37A2NKICJJtCObVRUIWHdUUsVFkXjTxCWS
6eLYTMJXJHIiBi3zmkV6UN7vjZBeI3VG6Cvd3vrdejURhp5nqml+WohFJzhu3LK9
0QV+1UPF8yAQS6BBH+lzeKIvHwIICxHEXj130bH+agLaLKkXC7vTRrCzR4lV6Ezb
upDrDdiOT95pkLNRrhV2+njZnk7wD8RxeYBivNKNxtQ6L635Ds1uGNdQhcz7JLP9
rHhC4gkL/IidziZ8q9sJblAn7EpVFMCBOrpCJF8rObuwVHhdHKDGku8yULe889o0
b/B8JvdjjyHDsdrlXwPpHdR2SnqoF4m7wkUV/i4zjLVtOD1TBjbgV96xCAVbC0nk
r5J4GMDkMvX/Kc4aEpDPcW41JUnYwjMAvIzFAQ94qTNhwDux01SvDyCO8yEQjc6+
XEFKOT/nCT6AVqwWOhUttFmvN/irMWACYnBDfxOiRpDcONYhRzlcKPslCkrGOJzq
dhOqPDKARHPvWZ7MGfbrxeN7ja9N1EXeT0H7MgitOtrqdYQJdNPOjPY4W982uOhX
GVZPrI0xDduNxZs2uP5bQQTS2DpvXl5kLg+EMLEnuytUswP50rNwflQpHfbhpYQE
0jjHme1jBzghcJyROkgzMK6M2QvceuaZmykVA/F+3+L++e/d4lkFHdgP1dB2UOiI
KB8s5AzzewAGdxjPFtQibjBRi4iH6Uo1FSCmo07Fbu7UkA6EHxVQgssOq34HZhdX
7U6x4MSmvpMm5kLtgln9JcrDoEFiqWGe5Z3wSq4YzNBoAe/8BYqM1FrIUyHDQTwk
UeYaTwrzphOHmW+92xTy5NT8cM7IOkMhjEIEO425mioX7rRubxIjSvprhdRinO2T
GIdLoIDPd8PrrQt81zfg1A6BpzW/nj8ofhbPglhTZnKiuFPYaFt5wuVpVekSYqNs
QWaIrmE4M2dzaW602ZP+mJK4+lh3KrOYEBxGjhsCnAO+7ui7KjO15t87lrzL15sZ
fVDYvcixAC6qGiwOWd+UhEqe4emQXM2u4rGyjYz4+hMyZIYytvIg37o45hdVfcl0
ydtZvq8nxH72EZBIj54dkM8qaTJspycls1XGVHUlpM+cj5REshY61uZ7XezTRnIu
oD72gnLKgU391QLYSrw8+ieni3V+FCU9OWrq0g0FVNy16yIro4PbLDMM5UosGozh
qmzsXFvCU+JRRM2a39ECKdeHvTtlt20kB8zG+fg9T288mNT++BpV9kbMspsodAI+
yPFBCCE71OGhX/ytHNnFYgH9NS1HNT2LSGwiTan4gYEqZDr02l0PG23PQFNM8rVL
9SJA/yEFWVciOFxFKAoBMPVHh73iei4KWN4BT+kJkifKtEN/w312Kc3u7K9qzeEF
lGiwgqNNG0T/BXKkQ1ywDKOOSjBkt+4u1+NTqgwGEK5879ghxP5jfWi2VOf+l0nb
nlfI34N9hDz5OtLdHX7/Qq0uNRss8sAAD+bRc5lW1y8tRuZumRe9GVKcdnIOw63a
VCAVIcKkenJ0u9cVHL9Y8NAXO+5hUWd+oEND7y2jzlYYuXCCyVRc4ZuS0ibl0yzt
wQP8nbYzyEswQgzxYcJWm2twCwOekqWUkLXxpvGmBBk/5bdm8adImtJLMnIKqm1q
MlPoZipAoQ9dDdrx0C27S0w8oUbyMWxQBZ0jsLgxmLsQOR2TyzoCavkQKWD+Oil3
w21Z4av/f3VLCKFkqe5kWgJej48X12/zb/ZfuONSNC9oVhpqJOy4vgzLzmZd1URH
vdyk6b26UKKXB5pLnhnybLKMxeTUPTNhYGQ7Bf64KoZgj/aDkISm4IrcIOIFTGpR
d+CAnc/kMf81OoPoYN4LZK2zmK/alaP0Ypbu50j5RbDyiv00hCm/PiTFAQHC1RoT
NkQ+ekUtDyznk0WcDddLUJp0fIYT8HaywnQQYrQLSBIv6H1XGSHgokdjPWdWj5Vb
OTP1H2worToagPTAb0Iy9ZUZP641F4HwYuoeOmXx1ZSLIp2yjdO0E/qh1EoQ3j4F
dbyupHkDtxAcbG4cJwnEnpcarQ8GpSe+s0cVXkPi/54cKL2Z+hzOw3GbfaynEBUC
Wko1UrP/iKf893g92ia65QMTmAczSpF3H0yCDxZFsIcLS+ZodJbMBmv8r3PavxLf
0uc5a/caWDd/No+hFUxFg11X2TAE3QLPR5Qo0jXXV/UgKUrtDexToYDPuIJv8kZT
VaH8sk8MqdkzQxVy+0Xm9wqAGufTwYl8SXapSOWP9XLz2SyOxZ7GooMfebJYK0cH
paLQJB67SXNZZ7bhXv/r4t14SCmPesW+qD5wzZYcZLHTMHNYjiV9CLqlEks7REaT
P7Jvxy4jTzuVCe2uZU/J5O54exUgSBNP4770HFzfuzORH/8KeEdjpUua7URdQA4Q
KZIt9AEKBsRk7D8gqIvYdB/Lw6AQd+cvvpmmKI8LeEs+rVFuskS9s5kXm9acQTS+
4eQK/Ezl417FPtGaBzUigEDHRrLkVJ0OKNZfkU55/9KspTF+kRDyf5kQEHBYBdH6
nvzWLdAUg6Itf199KdAMTlEB4Ce1mhdk6OZbHOi3IlTkQGzJDv8MGTJSaVS0cejO
ANERCZl+RLQd8eBwDGi93RgruEe0f4yNJ9TYd821rxz0COdLR13dwS1rheGtrWx6
LCdNqGCZQLDpTCfywWtsaRESC5hhtJYyY3TZud0MbYSNDTTAypO1UFGlA9VRDkhk
gyFADYl2OIieacUikW8zdAhrMXPyIKWFsc5lWA6T4bVWQFxP5+8fWwq03yR0V14I
DMHihZdcSRS7iv0Q5SZF+9ohrWFX7sjasOCDunEG6nkRfA3UheM7JDw0Jd5Avh0Z
2I2t1971K99solFOFKMeDaSUf3P8VbRZbTBQ7K0Sxdgn36mkvq9EXq6Ct60OMjbM
0PvXxEjcTK9an3/dIlf7408ULmxSk9neKcFGpXB5IgKB6AIs6VVXMjrsY520Flvb
SmCajdxuLfXhXe73ZlHMl1FjCVpPAFm+ShdlgeG47SxroCHBhTgKXTSL2HqB3O0b
PQTQF/DWPQL0VDOVLq+t6+6RThhN96eXzT05owAvWDNU3sRDQXqH6fFElwKD4/9A
BYW1CNwtAgcRlE6FiaIlkk2orPginnJn27U/Mq2QsYo+43y0iMfC0AK3wcM67T4h
CavAzTFSIL9Bip+tFerK1jQYOc5U93Qex9Z4DDWBzf6ZwBQFvouAXumuLu5ZWpiW
ecGkJKsy3mK6u12wqAgJSmb0U2NUzeRP9i4Sblnm5o1bcflq/pVt9S12k4hZKHd6
uWh6kxW26LiOSKqhI0W3PlqQ3+klsT5Tv/NhieBP1fUVM0S6c40XjCxEzD6Yn5F+
3z3XGUDbbM+LTIlvz8VTbIWxaJzsah3HgFIiBsXsb8hHO5EgomhdRMb81H64G0gc
hpTtnjQdYUf0UTjTzlVCExDKJdODbxURaA+vWfjazZ2eGE/On57YdXVfBJ6aexAr
Rgdj35YjqgXi7/Tk4Ao/Xrd0CF2R11HjWHuTe71I8awWv+SEzvM36s57xIf+akTS
BV/Q0QWAyZ24h2ozjGooZO2Hqh24pdXq7SEtA6fVD3/Q+F32Q+PA8LGqSC6ZL/9X
uA2IgS68ZpwOwjy3N/2gwsm/VMqycx2mjcM4ntjpHpl9LfjeAVI3nXKWY6ncx0/A
igQtJRQjkjDvhfXijJKCgR+a8D44ppZH1cjbc4A9bSMGD5PGDiro3sD+dHZB5Kfr
tNm8F6HOjg1wZcgbQAAPB0x90sU8+CvA/O1eLhP3KmnHzS5b3NwtYihoeTQubpwv
LbtTYWuPov+kbnpSi9BJwR0du+r3sh/lGlhBW6q2Yj6VRJpB/D5ySCCXBOXcVaX3
vqndwyXHgm6eoNISyn+x/AQsNN6RNxMusR1/2nYHEIFyrZ3RoYbZ/d+vtwIpLZts
yaZMC4oKjkpKedEeunodx4xhxAkKL0P9G0dECaZjLZs2IVFKldZa7tKpuKqwk3hK
ptYXh3gPE0HM18bsbm4WnKH2fjpbot+86NUydbcrMfK75nDIm3c1arrVueHBm5rg
JEFrfALan+93TXpHcojHz6CZx75Sa5a47vha8k0pUgZjgZmbK0fW7+NosXOtPBwx
QdOsK9cAcILMP3gXO18beJO8LfMz2XWZ61FZI3AnzvfvQhYd3RIeUSBZ8ycBaq3C
gK/8fapHZdbzr5XP+pT81kipSNosT9XX6XSStH4y9rGMbl3l9j4kiGVMSHl5S3zj
3KhSnhWftkVtlSYvxH/SQUaN/0IQ41m+Aax4t6tCQRoj7l/H5sj7P1hYoiOLmQHU
ufJgpPI/ak4DxTgHLPyCikR52aj7G50HL1FmBzY0SH63hyk8Ma6Zoh5i7z0VK/Qr
oC9Of/UTKZRKk5hle9ZkiBGKd5RXBwAqKfLEn+p3NNj7uzSEf4qyVWLu+xlvSz72
DegXl9wZMQbTgZSQcqfnwDbqM5lEOYOLp9OEYr5IijLGV5SCimNit4fu6IV4whVo
PHibYy85XzHyckpW0yRGS/IZbr/HwjrTrVw/kN6yS4o=
`protect end_protected
