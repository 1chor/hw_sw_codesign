-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
csRI02LQVGWgJnctHnP5/aNoBklGMKZ/LHVJa/gkbSkzdS7DXN6XrmulLexnc89b
LwFx40Of4+8Xe7/9VclwshObg8SwTvvX06aVcZcfOCia8ELE5aeAlO587jyVhT6f
tDqbbjAg06pbtJYd+f9DDXGq7B3Tc4rNaYVsyVHmICtbztDnVbqyqA==
--pragma protect end_key_block
--pragma protect digest_block
oIZPop6W0IZW9VD/Y4ZGE2nxjg4=
--pragma protect end_digest_block
--pragma protect data_block
b446vqgAMBeXJ5IJ98KonNwQAG6nBexAThspfKNPkG/rklHfMqvFDGJizyvIdAzD
hN0Qwi/xc44LL9rMTBmvr+SwbrWlmkPVgiNfvzSQIk5/y7026ltA2EoiIOKFvoq0
TdPZIbDxC7zzJtuRvhipHpu/4LbucOg27qdqsTZYrHVlGji1etnBYFws19tXIded
P+9HgEBtv3ARtwM0tR2plF11JYZekhnXi2QedBruW6iXL7hlJ78A3DZ0VyjqnTfL
BKoZvwNHh8RMknQGplLDTui0oNvhX1slqTD7JDMICA38K49kvZSO3g51GOn7atq8
TeqiWH/BxeS3DokitVwq/5KNGFQ5w/ZlC0DS7Arf1KupEca2UUB0nczP8rq5up/Z
adiiCjYGSIZ18Ys0UYp69QZOw6rCExDk9oB3tZk1kJbErW1DdssrGZLCH8/1n5wR
iRfZ+/M7UvL9hh5lYvD62++qdkqPBc9yflulqXwnDuWtVHdws5ZrVXgLRqB+YIyz
HCzzmLrs86wQLmOUumm9+YFzzyrU+fgO5g0pprmv78bV7tT+FgGUqRzYC5IcyKAD
W92l/4Y5RI8Jkafkwr+BXXDf8pYp+uuLUA1AJmN3vSgH+uQbsHppNvq8RRWwjhzK
i1rnXKQKjxqhc8alAQMKCrPBOenMWKJmg1Y7mqhuP61q0mLFdmFjnCJ0kFz5Q9iF
M3nuZTAxXoBk51GEJ8+uIOWznvfLOki2i4GUJV9NRIRvFhTGug3GvAC//XxNDVOS
+WW5tpV5Ab9N5PFXFNSTJkBYBdkGNKNJzFpfHaQ9L8+TLNtEwkDbLvnrsA3tS1FA
Fkb0FQ/cJTta6tpXuDiYRlbL/dsNkGImQ7LRTzxwo2q+6P1P3UC4N0U39XK+b0Tq
sqBnJtWw1pedfF5SEAlVJPEGzm24T6lx1QFlIu+CrsmZ8d8E1XLP9GmyCtHLPzH1
4pvBhRUt4X8Ma2eq6oAVkEbfnGLdOPfo8K62+bV249Rmazk8EphqiP5cphPL5dUV
oVM2fSKSkuPmp/zazt2WtZeqL7MpUxAfe0Ln97VY1RfwBkYnydy1cYIr+hArAjPF
IPNo7Ra0Afi6Ds6b1UBe1O8kZoV6s99jYSYt13Aghp9/lrvMuuJkLgFhKlv7NaNK
J0nGBKgdSrLSD22Fmc1K4ijytmJe6+hdajpvKQDUewAdISR+qql+Ai5xGbHXlACc
fQLPcNSOmdNfMB8t9V04a5T8maRlw/yyIukrUVBXHeIz+4qrYTwaSsQoSK+H/61R
zviRWbgQyTYuMIhjohoc6I1XxP/1DubH3wriUiqURZF99wp/n2XFb2jq/ckqfTKy
tndZilTcNLI3qea4Mj4KqoLY3RM2EBPCdg3+/JZkddL9AWB1clwDM7bNvIZLoeif
mE+vw4KBa5DjRhT3tZqvDm6Zk7XadSsLzcVuOr4U58EUBhyS8QpSHv99xT3XGu6T
H4xBmQbeidNq9w0hVlV7jaeS6X2Mhe7ZaLM/0SnJBh76+L1UD3JHJ+KZcdwvE0Nh
5s5Dfd/SQTOl7XSMPEDl2VeUmkHjmXkrcR4UsG3vCW8tI2ApUhynkZZ/iHoaBMCy
7V2mZVzu/RdOjJtsgGheFufLRNK5pjrf5js3nTzOxbOgcMZuglpwI3FJhsDvvH3e
jbHhArhlXKTHX6OZzMV2gtYpqLX63+pqw4JHNdYYj6WLz5OgjP4CIU2Z1jgXtscP
4Rkz8HPB5KkL2NUuEHgC3oigVrrkmcsrw1aRJtrGbGfRF90VNJiqrEmhmcLyLDSx
v7YFl+6yLJAX+wvWGM8Q7uev9vqtydpRUtRWnDmgl46Sj+xxT+fNJfGxHd/9qg0i
CcB87FJjbRHZgufnblXyMKWeO3fQjpBVD3A5ZCXELpfElwFRD5IdyjXTJddjE3wb
cg/xIbd0DRWzIj7YUiNClnHC2ypoFagaazOKAnKTJx1/XT9NZX8rV/RXDDoLfhnQ
tP2hMNE9jP8w76mH8zG7ddac8m/mgbH2GhDdh2HyeAmOfhpehCfuusOizBWG1Twd
ukJLnFnLDzPd5pmiw6OMZ0tiG5HG4IHIsDFlXkT+DGOBJbDs5lIMP2DEPJDYFOwd
s64YcqorKq375qlNVE1D64RutIwRBn3CBHuak/VXyY9r3uNFwuKMWN88OtTa7CPm
GK8LAuaFg2GyR5+0SCQHzkCMk9WLWOTO4lApglg5eI7vXfEMxfJlY3yrdnBlH25Z
ciEIjT8OW3q1nk2qRxT+uKX615m6PPD/5iVrIsCN1zuuIhkJ75/R7mi+AJXMwQq/
goLUgZR17Yi/cnuo/n/kqUk++mCIcM8NQkAYk2EOS38NeMvoLxX9EZ0xP2SatPbF
4Q4ZG/iUCVSKnF+4MrIR4rQbu8bdkmZW+9zIuAu4tNapIy0035RPZ1ojnFH53+8S
7E7OzLi/cFnelQXLlDbsDdQ7y5oSbagal/HN91ZBD2CicbNDs+rft7djdBW+Raz4
otweK+ki7efyToN+dc5iFCSEKBsDqn97CgGgtdSfUDtHKcgdHP/YJkiGYk5XBR0X
XE5uQc9uhGEeb/5cdjfurrqrKH52Dfa/FOEh7lgJ2OIqBOPq1U5IGS8KUYv8UA8B
GudILF0Hm5Het6h9BFfzzkfliKXsYPKo3hnGnNwG7whpXn43//WatepEmybX6sXG
0VSPGF2g+5FiGPR7SIo1n4/fdif/JfSKFi3rQFSnLNPdC4jgr5l0/zgGiyvLj2CS
Lk7DCOcFZY7ONDCYzJ/KoApsOyCm3DhHwBA0xqcQQCqkJ2wpXnQa7LIOerAcWTfU
KyR9VUQDelYATekU85Rs9diXo1ND4u6GeWKcWgshJvGO3FWQckFYbDJ/qoFImCrE
qmh2fJEPSeDiEfAfW+9MSeISQJDxIgvsvATNcsZjP1sqKz0v9ZSshNtOmLTzgWEN
VvOoQ5qa7Xb7UN48rj6QeV/5DYk+wUVCEGjYOAWCkmUTe7+JtRdRyBi7bYgdNL2e
h4/PirqyE8MIOvSlYGipxqhqnZ5jG0dI/X0g4oPXJgrY5WzONJqC/BNOocMGSXVq
DKC3KjGk/UnnujYVWBohqnyFHlSBGK9lb0E8E+jkeAS62EijGmJaCYkjkl68JFsX
IdY24FcdpqtjpVD5mDlNa8C3i5W7rD3uTEEHmyid8tcL11qLIhnnlIX/QhcSXjm3
mM+5YdI6ETVbITeuYGVFUm5yyQVao2yS5y5YkAlrA3FX3q+9kTn5BVjCLuITThB5
SyZ/++jitTk6kyeNh7RW7gVkfFzphrLUgo38V5QVQo4qwHgrJA4+xxqMdhlKOR2P
BVXHHKf8/33MZWQNMRXWwycQLS/k5qXOM0+63g7GNzqDU2j0+A1b2BQDvSUPmZxR
p6Mj6kR08fJBcWQwoTxL425PlJsrMmd3vpZ0nRU6G5cV6S3wMfue+SIobL+HvGCW
p9a9z/1sLeg0V2I3sFP5ErkUYRVvjrklV3zmsgh9+sAc7og79IiEESPLM3IAjI03
znkbI10L5ECRV0QQuyBwuYpdDVE0MJg3SjK0bpbTfmjlQBU6bXcw3hQk/dk0QeQs
QLhxMW+dAfCr5LImEkw7/HorzZGajslSi6MQMrG22c4vO0uxq41UoBEj1PFuuRvR
6hX5MKz5lXWfRIXMRJoX4rKAyKbAVhLXkRvsmefRbk40Jn3O81P0Y8Nf9iR+UCob
Dce2d92GTD+aHkiXojabRq1kOKNcACoT4PT2u0l1HuLChknZ034uSKUbJvNAebcg
Mt4GwHq9pJje2JMec+qY9r2v4loVHJxkZH2nROdhz6ivaIYkFP76moljE+1J37Ca
SJdkT6nIlrCumBFnjdcSfXO+psoBwE5PM6o1znaoOaBy4/3xXKQPuvK+O3I+9nr9
wBz9xpIJel5STDqVViAFhXz9ZoRXLfpOB9hWWxFqYWyW2UELG94efAZZbRdl2GBn
Eqym6B2h9XAM5on956RDO+MwajcnmAxsayI/nBHkOsFiqsHQoFmPEfV8UWqeMnUY
H9I+mHGQYq3UCYS3rwN6+hozOBCyq9iG62Wsxa/9RAKa1aHgaeRBFgqKShzMvGJT
8V4+JI4i6YcWKpulJGHyb65jCOLC/K02k3xboAam2gXL/w2CmxayHQQx9xy4HrbI
/Mri1ES3zAn5wBugXS9En4bu0J9i5qlP6ywbQJJ0akS+s2S4nhyB94l8oUR/cFoA
RfeCSpAjMKAqCTwOj+Mv2xpp0QM8bWTic2vsoFnLabnjwALwSBdZeC5FbcEaDclx
ehwJmuz2VcEXsTY11/JS8yrdsz0qu9awzxY+GKyLJ8J0md50ci1woaDC0WTZnXA/
tBh5V0/e9K31P0Vg4pDcub2Vo4BhdWUPcblGFtMdnfyajT130EMuVm8u0N4LgsRw
CRrZd1mzpp/PZvTsdhqHxRQ4vfD6jS4hHBWUQd5uGsCYFbaONomfv+UKmrL6Ammy
UPOPbIhGacbjPN4cB6yhm9xwIA1JaGzURWlT07CleUfkjhA++ar1ncSORQTHinix
vVpO5uZcOhRmtt1A96ADvSsqPaKVXQ+iSw52+XTnrN+8o4BAdpEkRWNYUhUqkLxY
+NtkCw5IfEY4rzEQDOmBslGb/8LLshR8gbmDCl1fhXogfoj7/pt68to9H0tyVT/0
hDgRutRSjMCW9mP3/y1Ipt+YBEF07vpBRNNqJu7axaPXFCpl3ZJXq8aSNLeyGcj1
mKJFuN2hvBTnbgODbsWcB9qF3DfDQ087EmENpIABBawLyRtc3XOLhfbUNwBI7Lan
wuS/ciMiNcsPG63/BzGX9bc4mhtbC4gk2xBt6G24uip/gBBuSS3jt+lGbcshsfXn
+ecYCe6sezgdG1GBioE5flK4HZs93MNZQsnL9dus5xy89HpGQopR+uiecLDWODTx
w8dsWDP26m0Q6IgBGyhF1au4JvmrEwWDdHdGLZhMiVfxExmYVeCq05iAjQwtuYNf
uhNnAY3jkfMFuPDikM67uMwv4kXQqD2F94LSZajtPlvl7nD4LIb33tH+uzQrvXei
5jAbbbo6pMBRV46CyDAgi8JSk8AYpuAxYBiJegzSpyPjHpW8UIvgFvIHDxCRVNYV
TPrEg5gT3vHHiMYJvFUdJejrT3AQec0MWatU6CJ3UK9Mr65cq4zJQ0EgDSMWheEv
2TmZRtgDLm9/Yx7Ta3li9+CZqDWmosczJkPMVgiltyKJJTl6AODOiz0z7qoa8vAP
NbNX7eQX8/mQs7dYyYiyiwVrXZtTTyBsNBuEIWbTDKYU8WEP72Ul2rcnXO0q96ib
U1b+jFTT8sFtbQk+1VPdKzOEduIqtHIXUVt12n8hHCM16zkgdvylz7638/nZeM7W
o5Hd5koQhhJ6x+v1IxtvK2JFr6yS7KP0GtWHIw1uhzX97T9Mu7E1RRAQKBP4Eh7Z
AxE+QZk7VWdpMEZOEXUjG/4Om7R3S+7B5t6/E4UEot1Q5jQt05wB+jlLghw/xLiw
jwEX7ublzN3HjbxtAEj/wMuMYdG5Zxhwws2D+pDnRlPmFtCBPVgNvOOmscvpAJmr
iWt0V8SY6hpjPtyrC6mmpOePKO5u63FoPziaszx+lP3C80po6VdjX0Osvd8OMhC1
yD0f7XxCBd2kYbsufVe1PF0T8KyoU514Pby/2T91Ne1G+iXSFrQy/xqNceOEHj91
w5Fktr5Y5m0CoFBCtSXtEKypUzhUh9189gp+6Sduw1PzE9uIvxUjRGoEe+Nemwhl
5PUx1WJ74AoyUix7zhX5GI7qrQMi3V35CVAO+DherXwA2KLPH6mvnLAhVq+ObQoC
WySXkJ3qzcrv+Z+9PdHzhi+cXc/sVD2swCzanLE5Vc/tEcgw4xAiZ/hSzPniJvU1
X495khjO0Dxa6Zjg87N8wvXlEwKZRawZnVhgDeXbJDrilPEkd8kubPQBnunb3Jfa
ROEiX0yz1Wul3cHtQFz0Ls/fuEIniaWM9iK4gCRjNhQUW9qk7+ZPuEt9TqEooV5u
1tOMZCIxGwnsqohHjT5jOK++8YrKpmQKVOArH8Q0JmTZBW20/rx2tKqmrABdMhka
kWSTYl3Ukkow1Hul7H4lRxBjkOyl+b4abMMZXihCm7ok4VabMpXNd39W7cZtNGNq
MjRX9+Ht5neS3UKFEbTKdhf4zwcSEdRj26QjCUXkXBc99p4jr5yWWa+njeby+NMf
rpuXao++cdCpcI5h8h/5ZbVXCAW7VtGu4qoAWyCZM8WQNus0o5DNlL2YkxDX2ihQ
b7gw069RNElvtA4DttqsZwVJjotbM2WB/zZq1HToNBu2bIAasuFORn3nAUnKo65T
mVCCA7dA9ex+FCdfJTgIvf3gXy56Yf6j5ewmLWulrQdrO1QHKlKBvv3rfG8UBSQg
QOw9BHAWItpjUpdowvIU5mShp4BbxRQ08fyGnD/wC+wbeVKIKqJirX69k/Nxx2WR
UiqmvQpyFsuK52E0QebtQAWIQaY+aDfGbHQIpy2xvUup6Tc4g5uSy5PpLWNNskDV
ZIAsqvlfk9mE0jh+mnDPRGxknMjk2UpqrF55BQijAu9/I6DhleXjLgKkzfHzExQs
rDLpe3dtlFWLbvEtdR1FfZQsTX1rH/5apCMgfaAdQsgXOtSbyVI4cYHIP1bArZ2t
CDDG2H/f+DlmVkwtrabdnvUVJRuwAqEul27gRt/XudAsAB17914fXuSdX1Ubw81y
d0R40GUAp1j7IrICFa2vux7AWzEf+4YIA3h+QzrZ4ydZMCIvjSFb4SzNO3JXaEwM
FnCZc/whvKLLHloR9cj7yq/wauVzYWyw8j2r1h76ZG84/IBclcT4YCTOWsvVurcF
ND4ycrHE7wBMQWPHDbcd1zWE8URFpZL0u43uE/DAuamiQTNBRhBiYq4GSE8/GIEV
qNXyobGzPI+O1larJJLoJXH8wljrT/z84TClC+YiFbLr4xAmNQBSlXdtOvub2HLi
6HcxbHclDB3hKus90rg9SI3fVCygYniaVVHDdBswFCJpTK6jwdKImU2qomJimnA7
McgCSJ99awzZVsHAa8ml8cjLnD2ul280F9Wtta2qt8WweskTnGKVILlQI1sq8f/f
guSAb1SDTRAaNAnL0tAmXyFHvsYufctzIHty+hKV7jDUQz+gaa73CwD611UpOI4Y
4+O8BbIbRO/N7vFbpynsdByJtZtEqxR/8KPxph7nOK0q7+4Dw2ykPcLoEaV3X3Hk
fOdRzp1UxVKM+ACRD6p2aFbw6HPwsJu531SbN8Y+E34sIYxUPcFGSiJaeeW9hoaz
XAXJbQFizrV1OuV0+iYXAUBMoO0VmUAoGBZUItGRRvyZk3kUz+jjk4dOcLFeLlz1
kzcp34n/dBpDGZC7E1FwxU4TXIW6DBjsd9/HYGiEfUA/1UN7/mSd1mYQVySMZQ5C
dEay8NPpj3D0VBTra5ctxY0yrNMx6cH4Vp0SxPIIGiKayKkFkpGof57YYGCImYGk
FKEavMHRv6C0rvIKMvN6NLeUn1TdMvTAq+AZujkh3baGLQ5TLecwWBy3N5MQ5jK2
R3mY+ydj+C1qjunnsyj9OSMZtdkovPlCu/0Evovt6TUBr12o4yCkoOiW0QGZF2Yx
JikU6JXNXmpH5bRmtQTIDZFZaoapcnVCPSARuCEUVwVB6SVX8l16tRWSKvsmTM1f
47MdQonkgC1n1OXbLLizIBSZeuLZpJo27O1Z+pdp76YymP+rDyb0H2Z6rnl9DGCo
U+e4rXLfmV0deXgDNeCMPtCufbguXQJpYDizaLR5iyS4YoGfb72ayQI0nQDHEKGn
mcx/eLnHJTvxlavFQ+R212juDGi4xfoVw5ZSnhmaFJLj75pzeZK7ZOnS3jbf6Bmm
ZjRyMDCJmImCyUBpc5PCOtzBMranzvlebd2DuXJoRTR0HqahvEcthPZIgl01fgqN
u+yqdizgFDaaFQNqJXtlxLNUAYbvfFygwpD+BGQXPeDOTMetiGmgXZmAofSnmIFB
MXELqLP6yNLxC/27vOVrlXIbAXB4SrBUD7MNMmvMmzrnTQaP9veO14K3WgfYFvYt
XbHPbr275HnNzRP0gWQVvvwC9i3mWC1cbdfP+rB3BtAC++6jD4eXCocfPu/iD395
tL9CQ/YjLr2Lm+MTnca+t0Mi2pzIOoW4to22vBISQJ775lTM7xKjEa++CtfIUIX+
z/X4aMhbURODXVcD8cBeIgHzkB7h2ladrFo9cMGFjZAhW1uZmqHDc2q3tVEnYR+k
OW6ftQHUAGDx+n3y/S9Iq0R3XmLuixmrotgunm2k/B+5EyJ0cJBEpnF1KACbE82b
ltl38FVs3y3nOTT4Bjby6BRh+cxSMD8RCq8x9a2KlvY0V6rwpi17cbfz8CupHQSP
uPPnHorhg3HS7Ml90+W7iXb2a3BEHGXwghTEo1BNDjs2xUbHULNhHDSBFSOMS7t/
3lIBif8hjAfbHVdpxNrwBC2ubkIshHlDwhP7f0OI2nXvS7+xEpnwPqnVk71teUVb
6Amy6/ULh+EdwvGw303AK6mE1pLFV28jOQ8etJbMVjPJrTVqITGPQT9nNDuHhxoe
i5A+6SjyP8hvj7KTvx9sudw/lOq2b9N0InWK8z+nJephQnB2zo6ZXjOFnd/0mj8M
FQXuAal6/S8tJcmATF+S//Ji5cndjT+0VxUdrPCdITlBxH1QI+edsAGM2p2oO42f
MWStmS1AGZHCgcN+rLV/52xDXMpRR+UDXaF5hnsJHvhoQVKUVQ+wNcRMN3Mkfhr/
ETQqyr3cNh+pxrpjWnwUWDMLYkuYaYx0EwUWsGsRNVG6+fOm7A2wIey/ZZ5OfbtO
iz49UPY95KngaEJkt9FPWSLMvRxfP29bNFYg2/olrToQgq1PgNlQUgTjS3mvIbBz
YSYbro08+DcGdCDTXRVCgGr+0Jp0FT2Ivk9GtSGukgyaDks9eWwATXyK8ncn/SAA
x6+UJzJppil+nHql695h/qOOE8Bug4TANlHqDcmdURq6SQsCRSi5AYedSYozeWKp
Ugtq+BbqDEQYgoPZcMk73m/1qb017vEbb0QDXj4WkA3reN7SWBAK79a6BiYQzYHJ
b46lj0SRkQ0muD3j48vGiIG6MlpXRQN3xOnOUcGwmP6oGS5jV4xWekM6DTY+d5mc
LjQiVIngiYBHP3jDkiMmTOyNiXDgHSPRkFYuXpUzdY+QhCNbA8rdsBj/gkt2i7vb
4LgAeU5TQUntxanmXtVV2Eg9y/U1RcZFm5rBoVeO1/WmvyyWDW/0Ex4ASuqn8KV5
O9vcoBcHKXr58/acvpPNJdVjNbyJyOeXEDYoJGPg2VDIyKE7Xu1JefftCDTQI3iR
C4IGFbSaoBpwZjxM9qQyJU/r8lFZB20K/5l7l2/pzCePMwVWaT4zNIX2Gq/Z2E1o
9VJcSr2luSPKO8STwzSl3rtQ2Zu1w2uSYKdE3cAYsINt6HtJEfOWhgNvEDVkVQ3K
ktIo3Vrie2sDKhFJishccYRaSH8HbkKDauc8vka6Qz7BoXJhw+ZOYH2FDq1NEpLe
kly1RdUmqwWXRMbpA68mnLxnDy3Ga83q9/YZPbRikEpm21YegIF4DwfwwPItCg/A
iDZyFQl6BKa0VibEI93FU6zx0eiC82A5VNtLiod9uJukApLL3AFnSXL7yqAbK3F8
ZFfB3rSNTdmhBx7DSXzK+qSsuTAutkIUOtqdU3GtIp30x9VHQl+vLk9LwqZuVpeB
pICxOr8NQSNKSBpF/R//aWmqfq3X96l3oT2DprK10taVNKdRzYL2mBBgQPuUbg7e
PnQxG0dIWc6wFLUEzdo2MbFVZFHL7N34x4+LdorG4726azS+prIv0DEIpcF3aBzD
00g6duep30rnx5ppIOeNb6vvkylH2CRA2q9DEORgvJkjqKq2IL1azsy/gA7FXmk9
CRjExYi5usmlsKKEa09d9eMecufVEh6KqJLSasOx68DFEKVEIn5r7KI9I50eFhfn
EyUGY8DP2HLFc9GuP2Qdm1X/XcxdoHxRY5Ma1dL2vsy0q0tBMkwTbWSEgkxDcS4J
diLnr7oldFSInyiS9oCeBdAigE2GkQEP3V2J08xbCoIWHR56EcH+eNpGxoOO9eXt
4PtIIHtucSFWajXkVZrkCMhFB6gqgEWEYcJH8J1VWYREG+sHYYIQPV5S5Ac2P81D
qQxcmSus/14aXPHVIzKN9Z2Ee4jCsZrBfVKc45+bUwGfkQVAGfZA0Wpd6puXg7GZ
hBsc4EztZlXYpzvAuhj8nEy0H2UB0UKaLBzurlEuyqhE8swFRaMqtWqU9mIkljRw
m9M5U3S+hXPwkCC4QN9P20xymnI3BoUhBWM76QBnTzrPUQZq59ALUPdmaqPaiGPT
8F1ZS1p6utgDHCJaWp+LGi+RP7oH+H+gA7N45th0mYDAEq4j6yBG86YrepPdz8W8
emlTCt4lJ4CAQ1hBMXZhh3UAANTHojRW0JrUZ6sRQZnTL/JM05JrHN6VomZGAIGy
C6WJGzhCLKIpRM27Xjuw91sUpKkdNBcAECB7rnBTa1UezGHIF0WVT6E/kEdDz/X8
Ac7H0/YmxyXkQRm2E7H/z/F9ZgBcsx7m6QXnjp9KTSGEJOUkUxaB006+iinw1p8S
vBjd1W3m95ZpST5HODijYKUINnhZrxk6tKjmjn5sqLq623BYsiiBu/nXKEa0571i
tyRxdFg5ifyH7DpPWPK65JYZ39JyqniioJYU9N/OSF0gzThTK758YpNZgE3A6+Z+
ybUR0WL+jZfkccLp8MltOSRsu4FLcapAcmHtNFr94TEls1/FN8cvr9G6BYRcfEP3
TiTPZFDYMPYgd2NT2AI//Ct+EL91Ij3TZVNDAIapdKdkA/J3t+rwh5r97QSFcsKN
Ce+BH+Y41p+lwXoJWvouTkMrp+Jk53eTpFe8yTY078UeD/Z6HaqIT8JUkoVXCIY5
lYT8E+JyvrZYuD/JtNbkWTxAXOZMIke8pY2F2ttfnudEmpUCM6I+KrW8GgIO9BKW
vOqozMqtpBKaZsngNOm+RvpRVSi1PVPLqNU/TItKiGxdoqED0jFpx/uPYaK7Y061
9pmib92Ggi9kI3rnfF5bcrY/oG75sYnAYa5RoRU+OaQ060t2PyCRYgHzljxg/ac1
sBFKqmri9sevYchogDCStXU2k56CKY+fc3Eg8bgBub+vxDHw7eS1Iq361It340gM
2/vZVmHnvz3jS4h/BWn2AJ+6kXOvB4bt78x0HwBuc+37lPc59K6xwYGbn1GwxrH/
UgHTfhKohtIvsTIHNg9MfLwMc5jJl4SgKJqNoIr9GFSiZUme2NNLQrOtvayCqsSB
FfOO7QCWfnmC7s6ciTEg6KlKGiSPdCbdhPyGqCqassgllr86g3m4OsIwFQD7DzAQ
Cwt1kh6x6XqBWkRCbJqGLiW99Y4jAhm7E8zijUD3fpZhe8kcdl8SoIYIJMafi8pw
ypHGcUXM+GK4hzNdZsbajjmGcce8W6LBJJTZXhXtP6SECRhBg3O9bN1ZgB3uQnxj
83Wsw4Dn7cb2ll9q1knObIGuuoWJhH26iFdXcNN3iTSPA2VlhmcUmKn7txbW9aN7
U2tgun2XgQMnuFYpYgHL45k3UrFop8/GgtTmbkoP7XwqwmadHtyyEoMcFUyjhXvE
upAY8XOdx7vFpZfU4qW7e3Bc7TGFuJ/qvVjTjk2LPyrM3MFeHjjEG5pXenQrXYM3
Qc7s6/3Yet9BW9QgF0D2Ya13jja+2Yx9nl0QuWxmFMkgdK4x+PqxqRGU4WIX+ZfZ
P6+SmTU2j0V0GSgTsesDzpGd22/J8IbmTZIiQoejniC2ilUNi6XmxgZ60XrZy0Or
KDoKuHiHw2MqDE/+bXafNUF3RTnWvSxAHTBfuq1x75rvg9CBHgpRYZ21KB/qe0Td
xgOqwgjRb991PprlOFuV9oDs93xE8ewZnfwayzpSqrwscuuUHy3GyRgDK/cVzgTQ
ou73OWBeKwbbHfSXkqKswnvmM1132kRH4LcIKMTLH/GP/IwlTluEZvm4ykVZsNFx
NikIU8B/Qm3XzBoJ5MNS01RBPb9AXc/dmpLEE5idhTZ6frAQJzUtLJXD0bIkHY0L
BxPRvQluuo1Xm0JNUIUxYwHyYlNXRUSckpbVoW6FqN2QxvZ7UNVtqPHYsB27md7S
KD17B0sZkFqzCqsaf7RMO4wNXhDXSaiKADZDyiyGPwQXtf9s00+OUPDOSkTSw9Ie
cNUEz8c4/dppZXr/tJpbVckUl+/91B5cILZL7dMph3EbUpBMrA2KYO2RcKTbNwKV
5RxIhZETJNF7z1yGKgJLa14wbA7JJr286fUmWv75B/7dFI6hblI7Le/BipBJSQ1a
z+csESWpy32Md5yQPlY+FLbtXsThVeLMhrcqh6kHH/aHx1Mlwc3w64fZA9Sm/w5i
W8wThJVZXa2SLC3NmdE2Xdkvv7/OyrV7TXr+7d6poZ2QZ6zS1dEriRuQJKPcd22Y
zAgGbvyuopPWSVn9WG/xsevcQSL5PeS44QywBZ7YZLQ6r4YA8U4zKFZ40Rk5YogQ
egBNOvA5F194ln7eVSN9w3DG0JMymU3udmNxt663pXxyGBvKQxWwrB90YDN/edzW
YIm3lmlaLZap/HRuCheoAH6fIgJeZ8qALUOjyjXjTlYJTVGcN1hJFh32MBowGIcY
gIH6XqbLKR2EGf32tcnKut0TewtmvYP0+7+Cq8bEJDEoqLA7Yl4mAAe6Iin3IexT
7QEdeQj5iMB3WW6iEuCRmjX/0aMO1G4Zp4CMd+r7fz9+loFiT7GmFz6ISN7brPxC
WouJunzWrRuDSPU+xrdEb3fW4yCMlrPqEHwLHq/8jj9BaOV7op9NEHu+o8HVya7l
MVbF0oncg6NMv2A5gLJfPlTH0jJRINsMjJVQddivnQIkUkamJyID90CQqoWPOOtu
qfah7mz+ZDBzw4+0L/PrZXm9Xj2lFjOurGBKW8cVEpHCAjR94rf+IYT/OBvVRxzx
0IhNmRgBx4zdisJP9sukSnPLRsVE7rObLripM0NOlGxF1a/wTwhx9S8rGBFoESnK
TcSy1BaW0+TKPN3+efZuIC+WnPTYKUuPvENbFIzn68+4BTl/X6TAjIXA5AEiVCpo
K0fDJwsZUcqkY3oDMWg7g1o7CIgM1362gmDzKgJ2JhLOXeZXbWY5crQJIHOhhL2x
H1Qxuz48Aixkhmc8P5QfFaXVG81LioivvhZRWqVpcq3VBJ/u2RgavRX1/cEjvdEt
yH7TNRKcObVhvP9izz8mSfF0P+ksiZACLcqKII9pAbmLIVmorR+msQfz3Df9d3Zy
yohXqldv23wHQX4VrzSbpU2iKo+2+rRZpbhfnQQtJZj4Ze6UhuvnF0mCApdzJXKQ
x0bMhy1wkh3tSsnRbYnWVCcyvNqcDIPlePHxgyF42dokNQ2mY/HWEuOqq5cdBQFl
9iiNcykcBkHtl9yPE3zhQRXJGPwzu/XytQqP0sB4PhDUVWpl0Ju9vmBjna5Npwnb
sOuVyZ0o7b9J/6viV0tVONs6/g+KdqexFeIntLRJgihSi65wPo+uEAuxnCnO2lZL
z5Y+IXSdNNFZR3XzreBu8IXyXMzU8jeV/enDaeQm7NkuBJXxLhzY1/pBxr/bZ25G
mjy5f0Sq7n3HOzSAhH8Aix+rDXyfJcBglewGbhiJ/VdoVU0CU/W5bFX1I4BI04br
B3SK9CDDtod5xAPl+FJ+U1Z3/n0Eq2m3Aq0ZghXM2p7MzLh7FSrZsH59177qir/t
zDnQ6TvHaHVukP4MAT6F2ucJ8n2U7b5aCMJ5MOvYoz6wg5fZdEoeQ0qo0teqL5nj
ilZsfn8XJzaLPyGwUWdeOa+QNjDPjJLlhBqXJzBe0G1K5WlthVU2/Ml7gtTjjK5A
+ZPbla7xDGbqPytzLKc8O9/db9Et016FJa3XS6eYtLFBvjLpunupWfKO4aiG3vdL
UiDOyg2T6J+BnL2bSrOBFQ4yqxtXuPR7M7Iyl+aJ9wkcSW/AqEefV0lHQh3NmDH6
KpuKv7rwgYWwC2QLIVKqrTZWc2VSaBEZ2H+eMbLtVbOfXVGv0NbqHDhxRkjOFZfR
XBVjiNb4HeGUY9o9NDpVWN+2Qrp3EOrU+1QtLtvLypVWZh95Xn0C3i7gIsEW++4F
XjwyK2p6xF0MxfXnaRSGnK7Eym4VIN2I7S4fWH2upJgi2FdA9Ed9vrQXPxm8edgH
Xeo+4hB1+0yKui1W/qAl9lqA9lO+832iENPvpcfoeez3UVHXvXsRHIyFOxVwrgc9
U+lsk7STpqHIx9L1zf5pNTGJl1rCUYJBV0yU28S6uO9vFK2wqHPwHOk8s/5n5K+g
kfTJRvpyVkENW0fUHA1NVtjGe7GfV6TRSXzGkufJM/IFRHR1qmQOdTJSHoKhzcrz
cUflPE91rhng2mJ9UIR0nffpMnYnn6DbnNGRdiYgE4OyokVgcjkgiT8H4dTJtOOC
C1P5QhIkL5qNp8bQqS3rph+DkfYI1TLcZ/2P/hLmmMs/0oZPhjLcEN08qLAHIZVk
fnaMZsxbuslc31ZdQafhLU6DnwshhnA0S3QS5HhYyvM66cLohEPBC/s8NMo95HXg
eTShaW+v9g6ABJZf3cbqZDE52zwQpsg7ghcQm6Yi09izNkAuu1y+pVKhsSCI/F7p
is4PaMkN3827fB/896aJ9xKn/XV6JK0BOKX+PTxlKB+qOT6Q6oTiA5i6KOB432BP
Py7+qbiTQJ8UflOwCuBv1yWqui8r4c8cQSfPqxWFF+YwfXeWaKX38ywHC3z3lIAI
v+bESg0P1iL48la7KwtuaASaY2HEBWv4yrJ25swkYluuB1Tt2YaFlpplpC6ZsC5J
IX/OWHmI8IOdwHeuO+cKF5427117C85FLps56d4odXiwVA6t4jSxAsx4RhshaFAM
t7JNo07ggebBqwBmmUIytDNKZ65ThvVLN4RWlhKyMXQNKOeah6Admmzh5hgAXD2t
gC2yUge1SNA33+dtC303WvzbJfMbiXOeoExIdi3YE0mIlx8m019wvgoxov53hs7I
f+RBg+n3uUh64Tisl/hZpqCA4lsy4owq420HBq4nscqGLZTbrPcypH9f6hxaJwMZ
XjbWFWDAIsXYH0bOvUTqY1ub6dKg7qSmidXF0oexI+GMKMjMSDLEILZUMVrE1Kwc
GweeVKVFb8Mz49iw15rR86xwkf08r4C9ecyyNo8/ecwrErVkgbL5j+fcM7xOCgkE
DeA16aKvu7MYKTlEOlnPT0FcPBkrLmMDSGF63tOBoc3GmsIV8sw4NDhvG9SLK6WK
IRXBfaIrF/D7N7xKlb/uIW/6BRVMBBUcaUwK7IpGIl3+E7fRazTm0y85lhGbegJU
unXbzT8ddjZcVMae5r+NDNmtSQsswDFUvEEtA2OybQk9o2vqDZ9U8A0NBIGdAcuT
PLwB/fSmkrrVMX/SayrS+NprE3CnSYC54TFpBatjsAzKvRCw/EVyCU86xglU4g8n
Y4TKwYuG7IfY/X0jKpa1j+6MMGr5d/AFwsN14gxt2UP53c4uJZAiKPGfNHYXZ8a7
8WedA/MLjGcxzCyiXS2lYzIL4BpGADfnocvQQloUnvmNV4LBt8RFIWwVHsvnZ9qw
aX9dnNNW9vbOwrU5Ut0JbuxikMcFuccVZX9jFdnFWY4YJDcuXGZREZ12N1Cyfto/
k1s26xi31vj3BmQB2L/o0iW0QHYe91OR/Vsq2vRqZ4XUBmQaC1yXhRdqQhPJ3KnP
mDP+9XWlZl6XCMwn8lCaZ5kPWxqeNV/Tti9eXmVm4NrRFsnyzfaANLHaCddTqkIN
7pFCS1wm3SsvqM5tzYhbM8VN58Kw3AHoNK/ZJZFN88ifUZyqTl7ft4jn9cv0hfpF
fniliJJjXlRRBKTtk4dL4hMfOE7vMaKOjv9eGLuRcnpw3UkYB5+pJgmXpW8x9qWh
rOTF/Qlasc9vuC2AiPPAMYeYyR7Hju6SX5E45JN4ZUtOXKnElHMGCnrcy5xTU76b
QYdjygayizV+KbHnKEGc1/93tlovbKIvWSZLxKWVCC9Qm6JM/H1ADfXyrWGRg/XS
owumOTka/I0mchQOuPlJT1jbR+b8Dj8Q0BcKRMSF8PCG10Q/u1mITB6V87HeEzI1
x1Th1+TG1tTKKQ1kRLvO6cxjUpW89m57Tx4rEtB+lUO4RaSxexsa/pPQbQry9Lnr
MCyt/SuUf5/khGKZmXMGzY6n63ioN7DLj5M1NJlGo7gL91UIkDd19iMOYnYAZpqs
lLDEbD5Hv+kWr6ZgGcQsklgpgUrKrjtUMhAXEAmuRBP6DVE+BI6FnuYkQTdfJpqf
X4kvl04v/IEnhIe1kregAs+nNTJ9Dj0mJ4EVphPg3MoXzSgCq94SMtf05Q9Lnnr2
8TsN+MwVe5DkDgprYqtJX5Kqv2OJA+zqwvEHhW4Tnag5OKoFowNU9uGcnfa45PKo
TLlR90xbv19GM01fatc0QWQ8zYXwgxtIVG+nJqbKdLGfPRDOda3ItKW5dxbRVd0U
1xWO6A960gs/FOFWP0S5LNj7vOXIo8026koVbBQqABwRITiuer9c1cmqhfx6NWjC
y++W+DRoCYBWfN5i2fm+ct7Fn/SosYseMYJ3lyS5IyogT42dYE3r5a1b7SOdJqZE
/aqDhSNnGEoyAI/wxIkEG+vEu7LTxmKA415souNl3h84sDIK/8Ttw1dcP12ifgSt
X1d/0BHx/2UoX51rMZXyOjhrF6ssBcQ87xJ0iKczdFY+3wJlQ7CBO7t7bsk/jk2M
ssmMkKN7Kpx27yG3NuRPAoqs37CNUoD9W4QucvLJnq5uFkLtZYb/7wLrzLhEQK2B
+UHF2WuRIadbIkuB5G8esFds/mYV/YVcIJPfbkTHs1AVcPnoaSwFGZgrfGtdX6qZ
rSFql3mxcu2eCRY5KhrSVcoxJzyu+HCvhrsZR/uCpqRTnWw0CyR0onoKPUocZUwe
X+ESCpgPVilf5MDOIYMLJnjUoaxzaUcI4avLKbxZUUPj/s6STqc9FGACIKla1sPn
0Dr39C4xH79xLpNacRpNfvStUEi1GNHfCdAeTTiNOGCAqtSrUTdZaIiTRLEBT16y
cuUE/hInK7sYbZeCD4+b/2WqSTcYFQtLpLX8Y4kfcrHCLz+W+ssr3vvDxczDWlm5
vq0/nSut53Ie4amQEQOLJQnlRa3OhCu4qdMl3vKDhc2UQ8uYmYrf4taR2njIDNcy
D1XmutS3vgoSVWLlNYhWlVL/ELvK9zZD0K3WeywDXqC6pKIZhmmSgA4CJSrTh29G
ATFDZx9TtLk7AwNBJEQo8+kjO8s0lbBjJ+c97tDc0YvtHlFz9+3kcbjLHVHjKlkU
BvkJsg2BMdxwZ5kPs+Pyca/CZSXyNDVeoLZv+Gg4DlPGv1EjzMZ3CM/g/ky0Tu1e
RECXghr3BZgQHgYfyX4C7Bq9x7ehP7c1z6KFVJFvh5yZq/NxoZRqVJInL1KYb8WI
d2+30aySNwNFFZYPeD1nukEEeXDr4aclntmKigehzge1r+Y0KPesxtsg4rv1aymu
kp04F1kubrlneA6tU8WZhIYUYEsqE7OKJF5gUkLr/Ft4ZJvFftTeeDIbZk1LW/3c
b1QkY89zwVS7HE/82a7OGuBbTSHYdmpLm4G3+ZQ2BKdP3ouyRF8THOxwKDSPAgE/
GKTruXjBfeqiRs1G9ALbIZFGpq4FWUn674kQErpUuLCoRZnjEIpaQ842boV3czNV
Dh17IhAJoWJqmY6Vg1EEVjiWSgzjoVJCY7Opi96A7q40X33oBdxGFEaGWE0nRcU2
4jE5Owa+w3M7DW+JjwcssPPanhfymrHqJSBm1R6UjK6jxJktH/yGeMMTsSVYsviZ
v/JFybkRBH+IgB1vYz7fDWQXrUB899m8jk7b+iFeCfUfgPDpcruXYCGlIeeWCWOj
2cCOkG8Qy3ABUJBkZAh6IBEeWtZIKjZ3qcFMlv0hSZLhi5hb5fErTX5kJctBMyEV
uuUDpI1s03Glx1z/FsTmBq2mLkRUqYXXb7ajbn0MVZzts14nWc6YmQAfCNLioJ36
QUH18EvpuUfXyJoY2x/Vt2Rj+jCAFDDPu0V30tsXgeZDNdQ1HLNGj6go46Y7+c0X
SzHvgH3p7N1LDaB4ijuYvvDhVkTZyFSlNrVnbLyEsd20p2haKRlN/x29T+pDlvEt
eIp3liommbGSKR4r0bh8O2evQQ7MhAHC83hiZJy8TUCaK6pllO1iP2U1KGN0QnvP
8CUu2CBHb+LRp5O0XeJ84sUP1JMb3JXSJWx4/DziGgkuNM2hhggl/5qLTrRtIF9p
nel22zo5BXVoXpXs1g3xLtnET9pS3osDlsvvfRdnZ/mG2J+pmsNc/KFyUUGS64k7
EEHG4h8MZxif/LhnxFo05PujieHANznR8jJDqMXlhyoFF+st/Ev2cOFgk+ymLvTX
lK36o72a0ylYQecMz0jbXk0hM2stow45p43zt/rFaX2DIP4xRF4hGmtaUv4wkAWp
JdTACceoQB4db3MbVdSQsak1wdXNDr5Z49xQT3QxhFZIkHqhfXJVwOhv5RFbdYCW
7LCH5sx0CSJwbqCs+hEJNnY5O4d6Yl9CBDF8D6DjnyRzlHeZpN1e/TBQ+O5XJ6+5
/KovbpcHl6wkaWo3mUhz00xWhQOpPHTci1UokSei1rDxhtpXyAmaPGlR7Zlso8WF
ODS/YAm3LeSemBvUOGClH+blEafAjUOXErtpY/ZZmFYMXOpixhioepD7muSk5AH8
BqHya2IDIydSLvC5GoZmovwPT6xmRqKMwjpN9tVHoWQTYf/OF0gNRT2ZFfcIx4If
mlfF1D9EfFt6NnsRtnVbrzCboUQjWNvxVwBqwFR+evFAkqbcDjFEA+yIUXZyCZJK
N94MxJxcSc3QPD17EbVu1kts4Tve4GvjmbxwNyochzCV0oYbAuGXEGr9qBHUhHh0
/cTNmAZK1cOjIvsl+07MI46tsYTtvzs3a8+RhqR2VsJ2AK9BLMPggWUnFIhw65XA
ojqOXvP4MpD1l44kb8Fv9d0py7EXCj223Tm7e6S1FK7iRXK1Z++uZGlMmSk7MVrF
H48sgqKex47HHi1Ma1LeCbUKFPBrZnrHb5Lg1RIhrn1n1efEsx17KU8DF5KeOaTl
TNpU5z0vPqJMdlw0Us4ssehRnzIfB5YgzViuxNCiDJpdUNpuy5K09jYg31trRjyL
Avk3b5zc3mtBBL341WggcJTfTVUaeL6BxBzIgeb2Mh7UBop3QLiB/X1eeVUM6iiY
/H4dSVN+9bFr0Kadx1JnLCf7BSdamBzPIWX2ocSdGSlT33iqrqrfhbMyyDVeX1hB
hi/nUsG/ZiRwTx8hqU9BVp/9LVKUqqOMx3A9Q6F/8Bw9u6hZgi8jOvgD8u2GTCbu
l8KEKwNmnYgvsPAOzOx0XfRSEkvXb/wloWTbuJ5TjXZsmEfs7SiOMhKPW7pv2fmu
6rmRCk7l1xo2SSDxNxHog7ZYgqD/AjV/ECvyzhEVDdg6DWhyovb7H2K5Z1BWumds
tSn7DQS8VI901LkJM8OlAzpDAd03s8nLbTQk320zlKoOMXDu8U1p7wOYLQmrumrm
p5ANMdE/Qld2W/bZT26Cr/S9CdhbmVSEBSUEifnRNkUxaqxsavT33gZAvMvadl8w
a3RhaFcInsGOdxAL8WiNfpDWkDoVQ9qtFckWYGpX4AV5KJwZBQf8kp5LKqSXooaf
VS9slYrCFTCGeUHSRdnBdEalnRNgDJbGPAM0pMpaez+/nrLvs+L0AWDT5nbnEkFO
+ZLyXXpA8mpm3yeZC4nCR62NK8iOxtZdVUMNOVFiYtUdcwisVCHsWOeT4fDddP05
fc70GxIpDgLn9KfZRZdPuke5Xuw6039FCkBUkK2kIQWYmEflu0seZLmMNsXiJzRn
oEURJH2ATHHg+Qteusm3+iAw3VAtv8pTojslNKDwfKNN5R9ywfNOF3Z6woei0BhS
Az41V1XUCjZg0YN20opPFlOz9Rln271CLslIs1YoVMR11Jr6Y8wdR4V8wmlC5Hin
i4rs5NI+nm8PQTXAYzNAa3C8hY4wSqWLM03k2dGexUqwiKLOhP2VyURYbqudUdHe
o+9Ub7+cd1N4+wqFZEgdYQ7+69ZUVeT9/sdcBr4cs64Egiy6qUeu5GZWnTmjzSKf
DMaYUOeWnomBhsUrRmqLFVrRoO7WjM0GxMBacGEnHihD5B1/PP2qqnadTZjehdgw
WsndnEkURpni2CjKDeyNXsmOi/xJ7IAefv1J2FiVfm0Wq8mmY9Pc/PTJarw0meZf
CbfNJLeiBSYvBj9vnuPOsrlPhJD/ypi7WW5q8wesnirRzG9TvMvULgm7agsolyDM
FR1KWPQDwZnQhJ9Q4LWeKjcV1Kfs73KgkUV9sHDFk+xSNexAnC0Y+MbAuKzjMFRc
j4czS27sZlwZhi/uGcv3T/d1CUdVFIOM0+zhv5sxofhcw49URS5cf4Xf7s9HdZTK
EJLnDvn683u3iLZijF5oRDnH86KikPDMtYBTrECMHbbU3jnDCOBhDk7XKRX/Fakz
xBd2kQxHGUs39uDS7kknlndS8yq6n9BVVuUoh4SRN4nrvecPd5umV8iPqEKDrDEF
XQuHVcavijX8PPHYoFw8ZNgHmBLFihAPqYUFee+JvPZ4Kzm6fb+9ZJl5WvO5BqIe
gPoi84S+qeoiydcGJx5IYkUNkjKRV59lsGauU/js4wapDBVIgxCVXJQxRLclV1m2
1UymKVbkE2Trub0fktRs1TnGDf0tQuWwXG3cEWgc1E17EjMhR3n4oEn3tdkIdo2W
dQd3wIzm0+2CspZoVZromd6MgK91WdVWCE0uGAc7II1HMD3Cfu1sDouRPRYyP6Pq
RWqUME+5UGpz6w31Ca4RQH9lhbr7o1BIqwYVypiYQpNB/LMSHZrzs9Y0hsFKU500
DO4S+FhmTpi0dtNB7sC6ef0cilHUKTxSEq14u4fFu1vatkQ43+SF5m4T/J5FPimE
WifxC9JppBio71mc7LsZEbULXAGH5eKYbdPAUm/+e21/yQ0aeG9inD3VOsYWw3+k
r24J03Tjb1rfT8Pfoe1FZl4RuLbQWd5DQpnNjSW6vwqDPgBXPDcfemfGX+GaJBqO
gghe9iVZ9DL3KP0lKlgZmMy8Eqcqj2322OeV9OqChrROLzacE2VzKKdzZPn20b64
SxmoyYBowkIJ0vxWECLSujz1q81JAB1agCFyZA4ysxyjAJ/yNNC1n3taleukR+6o
nKKZw6xje2d+QAdLFefk7iInvLrpUWz0rJyznqSpyvRoIbY+cdNVleV9oPE+J1Yu
t5ES/Qv4dX1jtXOPEbyYss7bfy0LixziVYP6KoGe6Ckb56pc47DQLdrVytK3y0nD
QLH90R3df9vekDZ2YEa1ObqKUwx+ySli3i6j6cBwEAJZk8rIw26vlmfa0L+LPcSl
IiC4JjWgsXSxQ49SShPyNtIRR3wD8Wk7DYiJkOGhMQ5b72GNR5Y+94EtA/jfgVqm
JH0lHGFS0kkajcUa90AfBINyTDoGQke12jEKSaYlrfLP7wMleCynek45anOH7fep
kuPYdfvTr85GUB4Svu6hUFZQIwbAt4EN9ZsSSKiresLVjPNDAjLDmioW5VCj8mWi
783AxmPRJtjIlKzaVzhkt7U/UgJo9y9XUVIvkylW8F9qjlhGsQlGr35S9AtRQ8kI
kXjQABr664tXaEudox2kOZYYHpe/6QMcSz5C+V3lfbX57g7iAYPJDM1eu3XQimMD
H/1UfxNwhv6BLAIEQWhXLvRh1Punrl90b0ogAofuPh7FWLGX7edUr1BW7YhDTtjZ
rgLBWBJSp97EV9au5AlO8e3KxqfHg7424IErun5ZdwwbPZ8zdXm8d5KzdKgy/d4r
npK12ilzTaMIOlsAQgrOnUilDKpSU4fwT5DL5POQMtkuquVp17rWUU1Viz0q74fv
W4Kt2fm89BQw1+e8fNDFFlw234j509voFt1o7nY8i3OhOdJ8sGCe0Ct7vJJ1/KjD
Vti8JrmYARhwxy3mrBJ6GAPZS/7H5abNiXtikrD2J7/zXNtMJbYGP4Nx/qQlcgSe
Qr/wOQU6pUFMbnnp521+IXsWeWbwcicwQ4zq+e9UZb/7CwO77rkYyFe0XldTMCbm
g1mvGY/FtIz0whDDqIknWeGeBZaJBfMV7ND2Y/QEF/r1JjpKSYQ5DUY5pICMop8B
OWZi7fa/ZYQYgQb4n9+Z5QLI84TyJQAr7EYiPEs+arDiicCRJNvvR9Rbf+W+nCUB
25FXA7zqCD/07zElFFwmKqKE4WBUy5w8k/e0z7eIFuGuF9uhaRwQsNXXQE/HjUlT
VfKsD+wcbcxUfJFsYuE5DmR7mCBSKmfgn/884y648UIl++leIyc0iUNn5Sd/aEev
P004qBWsyTyPVnanE6DHdXXPG22ku/AudzsYDVgLOYU6Ly4hFkT4SU/9QBhb89uh
04UBYtl/68kKVrYph743jmWSk0xJYLrCEIsmt6xuW+FuLF5LKMzXek/xixCQRWjB
Apye0YeQo6TdeWOQ0n0Y9s+bYG1RdJc4HK726vPaEyuhBU3NAL0+tyxh95zModLv
vzM4Za5wVCyL5lOhXxjxK6M+4TNEollHqtJcF9qYT3RQXZLdcTRvE//sgCC3+b1o
jndWR+ZCfR3K5u09mNSw0E5e84OijD3SDRzGt+xrHg+lFqyUcmMo/cDFiKo2Q5qP
nKWvFHnpHn/+JiXBiv7l8R4d1p8sBZQN3+c/UYmehrz7YY/brB2D3dCmbJJEx+vD
mdU/iRQYflgtZWmUlFgGU/8J9fcq2rpd+G2NcfBYSd27nrcCwYkBjlu9UjEmpI9F
H0ApjS8z/0fxHtx+KK/4QJQ24uU+Su6b7mUBNdybtmqot55CvhZuMBMD2DI163Gb
S4RvCq+WjmkXqVcBRfXnmp4FDbnwq7wCzg/n8woPt3HjP+MicpXdUgmcfvP8PdZk
5XSbBgJcnxiCpiOxVQRKZ1sbkcQQvTRG2VZgyj7Ps5MeaVFOJpvdeCqfXAF5+h4X
XPMPeS2GjK4c2T7EYhxym8igt80D5+Ltq2kPeY0LKQ9A6kIbeB4Lv6JH0p+eFnI8
se/gW5k5RBGbWW5mceE9cv/tJoPaLz6m8d7MikrKVL5MeV2oxxhohOJYOq+Fcaz2
DKoIeNSIj7OpxLQftsJRZBRMtIXv6yuN+gSTxtmEYlUhQpXb6Yqhev/Se2LzFE+n
4BnE7GNmIGWmQO+zExYj3DOKceL11MT2zpHPe6OhdYk8N7a7a+B11xJ63MWX8lY3
UnERGloEXVn1lJ+p1UW8oL/Fzagu13cXSQpaymrO2PpatKosIuv1SR7t2DDY0xlG
18qAV9qnfyV8u1ZMKZ3dY0tKyEuAZHgPQacBHk94uaiaFVcSSOAEVHS/iSAY2woz
HNUeW1DuIV6SOQyOQB7cikxsduNSKVE+E/gHE3RhHNOLuwpo3onXnmV72d07TREe
CIIsjEt9oGpiKjAcVslspKxsZl8YxPze+I/o76qnMI8EUkj5gCx+w0JQtaq2HlEz
qH6X15fgdx1omW40lh+MZL1Tx+sn7RGryoHGkMVxfMHYDLYwPi8abbfAQn7jQSmQ
XNPG6HiWvezhJ6Kb+UVswUWeu4hS4n/zrlAVfOWwoAvwvSPNe8Du5RxmWnAVeK9e
2lRZz6wqCz+WKVKiMSOqO21DJvOqVtfuwcYkXXX8FF4eKtphHzzSxWaoJTYj/dyt
+P5GO8kqFzaV5VkaxXLsrbmzUMOOKJ5bishXDuhIZ8jqzKqhmulS1E4AkDSdzMFG
uLWJuSoCXPvzMt4d3ZqiYt1P8mv+zeRMHMB3w2c/k2LP99PKfT0VaKFvj51VKTEx
RwLVs5zPyNAL3RP2hS5lYJTZlILFtLICbudS1PRo85HVDm7UIQdDr9nvawof6ZqR
BpmjGqPPKUTZuH/HF37jkKGWP2pkhLM+l/xP16ZXy+QSh6nqJIfz7DD/pkTMtvb0
DEp73WQjyRHiOGeFIoZ5HHihJt/yPIjePaitRXK01k6w3opv87eq77wNfCzuOtFX
WJ5RPeAjv44icnQNP26O6DKrh34Yb+iAkYx3YjMHiU4XHIATJ1tJIMFyE89vruyI
BdeduEK2AJBQNYWZn60487al0RsGnTeyrZfqNX0Hg4KXRlUZFNYeMO6Fz/TqjeeV
rLwfDtOVuMlPvH5zaFYy/9NR3/XX7UV0YhtUyfB+muDtpWkzbl5cJLgizqtjCF+R
rSqZu6BOY/6ZMT+0mjRzH4FKVpEUDpDNFdZ/aTbeo7GEtClaT+qfC88jxe+wbxrt
8EsX02MmhFWe10Sf1dLDItGWwvTqvPdz1iWXGZqthY7YHLNUw1DTnrZkPU16mdwR
03rRSjAUvobLNz8XA7BdXmYudy/m+IsVaC8Of0PnMSO4CX2Ky0KXlkA4zhJAuHdn
mK+LWDhAd2QJitcygAu2GEltLgEQTnIFdSK3kdp2plhWp4IF+mCFjnz9J3z3BdiY
K7Uq/XTeeSa5Y60TmuTJvenYtPiGsngLFFHH2iY8rgpSQ7PBnTVme6FwN2M4aCS/
6nv9ZLxbKkumOEIQRyLcgiXPmJTs4adOF4D2qFsEGKP+KpVjCsaVT+ndxBVhYu6+
DXRQJBCx76cm+gSjxF7YCJHC8uSZN0K5eXRIYRDru2qMErcCUk8Mzc1P7OqSBHVR
/eDU+3yfBSB4Ye5x6E283QVSHDgWQdHjhfWH73s1Ll0B9/DMIv2CQt+ncUQ1QhgF
CEeonx3vUkC+AkctIX4yvX21jSVG7DPtsbnlbcTQdKBbjzz6mDm2NadNRPPED36W
rEyhxp4DgmQqLhnH4b8PuroAbFWPgN5Neq1oyoiTk5FP1odLmNmjsdJBsDdgULEC
kGuLjMapXHJ3DpJZR2wpsS3CMLNufCOhp/j+4FsnXNLDDxb1EBDx1i7t14/1DMBh
w4lvmdUR+TZr15+I5D2V2gN5FW6c7ZKUtF1koSIAvyGK2/YS6J5NQYX6pypEKEnC
48qcN4ixy6z89UREMkE7C7KaJwtuojq7gwUioXNjHgHlk2YxWUs0+ah1LnZW2kKy
zeRO8a/WeVe6JI1PAfaoG4ZjZv4CUd13JVcwM1Q3a4po7zyv6IyD/52c99UzzT6Z
scHGWCPfW03SSIJyYZIZe2qlPipWwFgiRlgMuvouVypSDoQ7//M8VgPgO1VC/+jW
mADWL6dZfXVc8vjABHEjWxZWdRAbv4+iUbUlGHjVKhUR7p+uJebufJiul4FY9FQm
ahzuVP8c63UdaAlKHCXy41xpzYr8xQgTFH8kEo4z01W6jZMUsRnRJB+bZr0K2206
bAGCEi77UM70aJAPvUi3eze5K/a9+srOV7/2GCy6cWeNWfN0xNKBFuFtByFugvK2
EOb+EiSmfAC1Tv9yxUut5w8DMMFtnfj4h30ZD6oJlZYYQPbMsLMaR7u9kZ5oMwBP
5RApRuZIqHdXfDJbwt84PncSFiIpBxm2oYVTLCDr53AczztlMcr6EZgaJZILQCrW
r7Cu07YfzGgR1Ct7oom8Q6FjcCIE0B1k2L3UCD0HyrhQ4BdKqKmJOxr8HYUWk5eI
Q9eEoanY3Xdi1yPKkI3T2la56vhTkHtikvqSwLs6Bv7Q2heZ3sEcOI0l39ZGXGTW
l37Puy0YzzmwugwsEp6ddVpq7V/5TvrLN3/DgorxZ6ObFGeUQjBL9CwiVa0c06Oq
uxvc8LHZt9fReofgNd90EzvCuslRnpnO384Fi548j3HvaW+HBcjFhnAs60tkWqX6
CX09xtkm1YY0bJhVQJgsk3YqI6lw8UOtdCio0mEYMq1zVwUg5sJa2bJYJar3gEWR
SOoWXr3K7aFvfG0tXceYxUN1vmF2Zb1hp/M+DojGH1qDFb8Rf4v2Tjdwl6+bbQcx
GkH1ccNaFZ8UTZbwUO1rFxLZMqlnOBLRnU8wwN875wBUGYYTjYFKtU70iBzza3Cp
jOaYWr+osOAXXv6gVeHZm8skF6LKIJ8Q+GziDov2dPaVAVrOH6S3LYll+lYQumE+
2qDowWel3vYSwXU+FwCebjCznbXMWSLwu0Bhq4Bk4fsS+C3uIQzeBqIiPP0Qulaq
hVhH8tdWqPvZAmc6HyZp2NtXyV1abY5ud2jyDTXyHeO2CTfwuhMi1szlG/Or1qId
uMHjof4cnsnX/+ShfAlsXB/Wrpl6N/pcENTTXYY6xuvck9IkrQKPW2E+mWtuTt5S
1HVJM44LYcqevIEGRObq6vOCqMtYa1nIwur78wUvSd/iJwXztr5FD3w6ylffyRg0
CLrUaE4KLCuBgBkrDkwo+bi/3k9fzs+81hCqbgnM54A+K7p0Hsf+4i87sffvFHVT
7N9nVL78glJWwNSR2mFeKm5fYoD99tJl7pBI+5SRVbe5k2EzthfyD6kZy24X/D9A
d7Sb+H1Xzr/skNzOqfMKVG60eKA6Wx70sLhGYmbcQY9n8nWB2dTBRTNiE8DNLvac
ZT8CJIUfoOph6trBhj6+de8msgstWKTSce8bS+cd0bnsiaNG/5DPzkE3GhwDcjKZ
uq+0iC06ZGkMZyZPFzLUwH53ZWzVyyEUI4hVgTdmfk68jLBxCnOT99dslNcsztXt
RXw20aolbZ9jfjU9Z5oR1tzZ4mZzh5D+9r3iUev4LOk4PYQIFapwNNyg3YVbei//
aD3FWKFAulAbrUD06Tjm6GXnJPJVO8Bb2rIZhAgJxYEmoH0atF7GGsEB3Z/stkLL
z9BYlmedQRyWtB+I6MoVS/PHWotAjP2lwgQLLRFzEakYH7p+T+l+MIWokoIgscgO
4iHxXL6WP2ImzpA14UUQJXFGehsBqX3PhKuNwZOR/9XKb3FvEGw7bUgNa/BnYO7+
zeGisCS9Ex/j5NKizVWfQ0RNlN0/TeWcTha+3LfiwElKFJopGu4jNhy7+HMSTDEm
zQ19PEF5S9ZgHatiFi9bPZgVxNpiH8XkGSU7BA5+nR/8Fqwrgm3MO+1+iMB0zFa9
Hkid9D2zewe9l7QkkAOuNrg/9ABXuOtgqiaiVfeajE7O3AcKvUeE23mbFFLXHBnt
ipFyIAeO255YDmukQpyFWlZN5Eq7mfdhzcC7oyha9BL+p0Efcxbl5XjtNLwH7asZ
qBXYSx3ylao+iPPaNvuB64Bbinyjp5sjt2ijVBE+EsI+dOyOxXC0waDFV3miJeue
2U0guCuUMoQ87WVSEiADta2Hl73ay/uh1Px7PKFacJcpq6+PZyFJuY877jM2pxOV
VK4USUFyNKOZzKEVZZSCyegVAUm6jLQO05Xw8Gpzjl5yUNSV34bS7KI/1vS+eG8Q
sLz+xa9OYGk8CD1XYHbbCshwy4K3ni+X9utvtqS3aUHvNIfcye4VZiEbLyHbKwjW
eyfKJ8wNJhbGcEbIVE1/T6x+DxHNLJJ8mwWOMJq5WcOvSb0h9TTHN7T06Jrj0fTh
q1IHFLlTGl+wXVhyhFt9tvCZDsiQdmw3l8e+nrehq+2Fo5ZBjSWES0MzcJVIyVWY
c2eTu/6znbggG0PdE52HiF5ro37+jD5g+QnsJ2H5ekv/g1FM6jjWJdC4yyn/2Bnv
aEDEczTCjhAcoWWs9quK9+0ZTeJ3EgkBO7Y1I7Nahu+NN0yi+2Hzb/S1aF6BG7KZ
L6F9SD5QnTtWXM8fTQsatteAWQfCApKdW7kDn+HrtQUmAL7pgScQZxLNa3aMxwg5
PpxEXGt91EOBMEgCgLwPsnx8xtHku3JdT2X0e9IDK5lbSlxJ0zESxurGxcwsxsha
tNm/EMC3pYqZkwwqOlevOFPl8ySi4FGniMWwV13TV6aZsilgRojZOax72g7eodkf
SGqjQA99O0CrVkyMlz2+xjBdwXQX3JUodOyx0IBB9otjQZTk7nbxSkMJmasVK5Jt
0plG/b1jakTQI9FIqyV+3xRNiLbGjYCSlsRbARI7bZ4eSF7Dt2HbyAiv/TgTbDnx
iTwbE2GfB+hnxeyN8l0P1yhBdWBQBugFHOVQWaObLKsDV22to0eP0mQcb3mCdXwF
6PZy43e6LQSsTWaxROTcmEhMYTZlhcMLZT6Ib2vSemBkvvTtqCTTZvbJtOxeGtAi
AKCvTA0qd42JBIpPY41OU84vwyjEOC9+ElXrMiL4mbvElCYNPtuVSM/fBub4dWP6
+1joXcBgvDUdD/3OhnIqWjKI6fszDb5tARz/LwFPGO+RfxxL/6WWFfgIbQ7WmXWU
2sA452FHb9tPW02Gg2lULN2I1LRMMfiN9z4SLAv6kb1EDBH8XascPPVJFBdKO6xU
jeVxu94xoVrp8+looYFNi/dyCkijnjdduKTKozRYLYmyjpS6Vg8orgsFhSMtbVrj
7yRHx0dwItJGddSCZBRnDmtSygrySkBcg6AEdhEcgzxt4ApMQD0xGtqPLkoFQT6v
ogrx7DPsPgiQmvReie6ogm+3IFXSFtDmlg7O8Wia/ZyFeblo5PMngC0GrUUBpKw7
cPp175y3kuQFzW+twRo9c8oxVk1kZSo6vPAJ7XbAlsQe7Nem2TPjxXLRanTbUj6f
a2mjUHXn04pE7gdvIQTiYEOuYchu8JtTEGwI+uwi2eW2knVeXLZDpXDq8fClaeBV
47kL5SIjyyTUUeiKJ+Uq0BbI0LwZmGti9L/3NUW5JDWAiQkzhfXATORRthDZ2IMf
NQ4fMkJDUO/tW7zwUimLROdlacQ/vjk8Vx5ZXFv/BlEgtQi5RTztEiwKxs40gfdF
1gp/PaMLXWyFnsr51TKC48s3Tn48QFZ3Ko+EnrohDAKuNUjj/TcBsZhl2+Z2/XwA
m+mxuv+XXKTFyaTVUwE9UhWnybg4E5fSDwNn/6v1uzmmrHMX1RLCI5AFTlW1f5dg
aenPN+L78bvu4axoB/eQDdqSnLPrDivez+OxWVZvcq5cEZuVZ0QuCZAmcDFgbXKJ
kF5AgaHxfabCPXGqY2CwapvuRVMJoUuKFCXsqP9dy5b05sbgnAtBaaWLLM60ot5D
rHsSHnoRcwdV1g01xkKh69UYN60s5DkEkiEZFjoxt1LKDVZMRl/O40TCtgw+p1zy
8MLDJTo/L2MHgUHS3EV6ILbhJJsmKITJ01SajHNatbmankK8losKaTRd7yWeHP7f
2kzulO8nt1VHUjc49uee6oezKIghoPsd6MElEnqPQR0/GwQQWihxpwkR1WEoefEl
WAcUphiED3d7H4gFziWB7qAe7tFQHWVjxB1Wplz2zci6KLBDD8VEKPeSB+E4IaWw
UprtNMZ2jLjXMtksMwMCvGTqYMtJp1cRK7qPuKrhh9olMBsIkpP3PyfEUmnnbX4w
wnGWQRGvBG0ViYq2zAyC9W0qGgx8JpcmOfvahV1ldrk+Cy3BhkLyfM5OY1E6EvoK
KHan10T9Q0TNa6okJtcNcwK8lB2e1+eTS3/cAVwFVP2s9ZnOAHS6BzCxUVsDG0Xa
BtweLnQjvUgIJlXOfQEwtaJTMfnPGf1QoWsjsdDhWWqPbnhiFYRy0JewsjzL7T+N
XBtFHz2c61LkGFXgLf+h60dxtg9H+54kxZ4SbWWbzcRw9LKg6oHjbk2XgaNt2E0c
XunfUj6YaDeNKKAgmQ2gyVZjjtUY2pCyFxse5/7sL41hjZRSilNwKnl7BDpNjdkw
mDATN4TH128/7ppe+S6onT36vdbFhP2gkL+T4imfFpwlAFJpZfhHWQ0oUXGTOdfG
d5bkM8whbUFqshT8N6XaFWXN2xzhWhXvoxVvksZgBiJyVLQ1xJLq0PPLxFkFOR4b
ku4ZM17ghNaZVCofVsmWGIb3lF+vh+k091XrhK4ufKl1G8rUo2g9E3fNPlYMrl3f
vrWd6L1TXGKwZEliZCPWj4WzLOc9kaQWZwK2i/CHmimtWgJQodyH/L1v3AIbqXtx
2pPqK1ky02rgII48RMgm209Rc7uK9XkuRABrHCJ4LeZQF6Rr3FWrDZUCAbL/nJTt
ayq/OOd52h8991MYBtuUcL1AjUYeXL48ryUwo4/PNs4Q9183HcXgXbmf8vNg6ppJ
JYLM51v4z73TmwuPx9fAoCmxQXcYWyuHLbtllqkzi2ZmmznM8jYQjMC3OkaPn3yR
clOvqBs0cIjCQlnZJcg/8dKByQNI1W09A23xx+HrIWvLGZrJLz6jSzULy1AUpyCN
MrqCtQGFS3sX7wB+TdcYTcHN0RMPpEA4MI/nevxh+oGgT1lJK0QgQrRE/3/SrO/h
40KSIOwGmkb0TZnx1QSFuik93gHdiSZhMU1BLEVxyxf9rfK0fjoF9UP8Kds3buj8
7zENowe6W5HqWSLBn3hfRruOj8rQMWO18afCHYfE0k3p+3bihLJ6GxsFLrqtqTYk
WKEoXbPV7+zeRYp07x1ah7nqcOE4aMmIJTpxOyZCP7SEJB71MbT600xCmUzA5aP7
KmfQvgrMJSiloyAnVUbBiBfP8fPrEtnDXZWuHNdxr/u9bhvohQ5hgoIUqDsrIkNk
ZZnwJET0Gpdzbg3fQCgrdInYMN70u4yEbmqIBMWnFDngQV6wLp7SpAX46+61oDS9
QEzol6DNULHu7xnqmrS99RCgIEl/LnnK/T2m/kaOzZAZJcws1UsdSnrfl4X2NJHA
bRWG+MaKj7Jb+1XCOnG+s/lamhtTAcYcPwVEWzITleNuaAy6MPdnGV3Kg+Lwm0+h
E49PUptU8IdtIkfHv/QtcuN6Z9biUDsifTjFHGuLcCYVfLi1CjJWX5mXu0JXzoqQ
8n0ceEm+KQ/iH0cb2aDKvoe02PjY+g2MwR5l8N5rSrJPbAhPIRfbh7M+4HCSGzBX
6933wB1ChRwDFDozlyMyuZXYDMYpiTDiulU19NkAqro3hrc+ff910iDn72wD8RRJ
2mO8glsb9TWFRwyNFRm2qmIT85t9qPraSDORsu+apt/HUGfxJCKU4E+0/pCPL9sr
Un+vKmdmEqJmvt+vJaHkdLXLjGAYux8Q24VOanYT/yo9MprKFyp6P8C/GgmGuRME
INJE++K/R6PtB7cX/RelOCYb1tKBCSe3/ST7r40t2MzRAcxCheQkSIUtfq9//Y3O
pZ1kG+L8pnTBapFYZOYZPNgomzyoTVOb9uiml+13Nwn5xUVCW4L2WhVFL3xqBh/d
YGKTiZGs5nYSSldmfm4hYOOSu4xDg4eZWpjmNH1GjG4GTKaMUhLBWXWSTjACFrs4
V68kBcp/Vb2+aWKzCJb5rjHEoZRLbAP9F3y1J8VjP7n9NFsWqIpFPeOBGKUXNmVY
NU95rS4P2bMIhihaeUpOrcZwxSbgceKtFQo283zPpBAlIA//uXWBvMxQaQR229Vj
T4P3dhC2eWA7n0lbT8QdpPv7wd6I8Cb78JAkTN43lt4SxyjhVhKNOTpO2xgMbciH
7IFw6lqXiOsD/yuWEazEja7N2/fzUZAzq9t4TR7VKNuKCzi0JefQM1AKJBI4Fntu
r7xcysCDTSJR8PQl3RX0SpCxPQwV5UTQ0VjFYHFSeNb/EyYp2hG98NBQVNRMMQBd
d9RUwM+jzVv9R92znvVXrXmkQgJHwPZU+ozmf54g30z7cH4GtsAHuIJ8938AhTeG
r+RJYLUrq/MEW5yDu0DPALw568aL1crPsqWYTxNrLBmeOo6IOFyPFqQ6KZiYDP1I
JcURQimIuCrlRPpDYzHz0QjhLGrP0lniVFBnCoy70i1hsZQHlI5rfotsh3dy9yMo
D8mkFhIp6TRXXSR2L3kSkvIuhrALOoTb89ecx+hTqaz02JQj9mdgKmRUKzxojYwL
XbvGoEwYwHD9sCrTqnhpGa0s73wTrDo4GTS75QL6FMIGZ+usbtf9tm80D/lETxSc
lXhOwh/uds7QGd4/qFciwYYiPdeyKvco5Pfvsb+1DB9VwPwwKr1dFH22KctzM2+J
Czb/utSR2mzc21+Y5/P/wkDs0enHm+SA9JRENzPc2IWQtKIMCgcF2At64IDqBj+O
zmx7wM9kAdOnsDxO9ZCjs4bSDiwB8MmUyDkn0KYHnofoqzfuKfJunstHjFmb37Pu
Gd66X0yIXYJKXqiuBxkmqpEsmg5lcFd2XcR86EWHMfkW/nJBfIRfUiBrfs2XlWFi
lJ8qmZEtmDVEF5+BI1Pr3Nq0RTcTTkow9gdOtoKeqkGOiLrXLjNJrX5OzzQ6fei1
goyBt3nZe9UWVC0oN6paf0DyRYxdJ5vxXUSmnLRkIjf7WtCAQWKp+jf2AgVwxzll
fB0JBKqRMbu7tCtajyH3nibTEVEMUVKaMPevcnHDrOm9O7oKGWsKN+5V3OA3N5aZ
PRoA05uzRvJTgM9FApMWqn5zMEgXHCBHo6+nIV0NrS0V43aE5KhyboS4OVi0WyeT
KUG0hhxY7JVChI5/tHb5vTecUnuAKWughNAqft/uVnJXXetzyKVLNHljHwKxfre0
KjPdCQAj2LHhaBt7fv4CV4KUxxk8tOe/PR+HIl/XANsLNLiYJzD+hsWI29YXZ/GX
6abpRIUGG6FKrXh2bpFwRt5GB2NZckbGAR96IhNpf7WOQmt57h3wSV3D+WD7JMqt
E3WlS1HTHchhffjXQES7T3UJr+J119E5FpFm4072gHdgBxeZdkDNTe9W/mTahGcS
BEg04TX9nOBWLL73Fo1YJzrKWBzqm8rq2J9gXE+0k538nbfJfkmcksraemh8e7lG
Yl/hOjIywbJHGAi1DEnyrFVbWkfZY9IhWc6bBA395LzyfzuI/z2JH6piVY3khjdU
PezqvsmbJOPksxC6kDsV2Aa28PJCOx9wb+XPl60AF8ya9bsRVUqZkgghfm791wdN
DklE9YxZimGFk1Z20yPm01ziCM6Bq4tQ8yB3PjUYs/jPy1DH6S7NoNWGwNQjRFhx
hLVeLa9wOkCevzUZwj8R1eUrDjZsAKRTy9XhE63m0rKH8t5Jy5KEFHvSpxwvBtC5
zdNyQ5Qq7yB1Ypqk8OaNK5gORnuLmq8fsrntzsRZp/4Qsk5Z512U6zwMe+8tClef
qFvCPoqUeURBsIyNT9DDDSAYhzURLt4Qg+1lEwIR7BIj/VRYRrZzhUti+uorqyGg
KipyeiKnYqL96nfA0N8RRu1VTOrtvXOEzgv33+J5SKWkuQ2MMgT8F/mc8JpT02p9
+tip0Z7hzbmolSENvKvxUvz+NMvt8SVoeLo1lr8Le9VvSvf0hgcPR95llb/WN7ba
I2j4k7rZSWm32BKmv70ACYJAWYj9nt4V73BX4Ibe1SBiNFASfdE6L/SSnwPsQw+5
wgBszLkZOn4xKacDRjpNviQiBG64/6SNEq1AyHSpjwjWnPlEUREpPkvO9Hp5TDgK
/E+/etsXk4SNtzBvwHezSmsBd46uvxP7TKC0QVD9vuewHYRSFjVQDYtiRdkKluM2
UZw4zx1vwsO1cY1Qk5V7Fk5BUA2Zj/BrRvTWzVnnePx9HYRukzQCXZ1o10jly2nZ
eNzV1DVtlV/ufD5nIamIsH/NRXbMhlBE9obr9T+N3vl3zO5inZnJ4Ycb8RPTPs6+
LqxEl01vyPMlEG7sUTmq8L7PLvSGSmlODHlSPlKghHuucUSnb43tc5bnfbAg1WiP
WOHm9NwnERpa1y2wt/6STgd4i/ubJrzf8FmhHI/HGw8GnmscRAIiD+0mH0JRaHt7
HuUytrHHKELFGlbCBOMSrHLdLAoxb9nRcXIaUQqwU3sKNyRtYnDI9jFonvaGKL/4
VsQONP86Rmb3j9nGDAMSoTXCC+3JaD4ZodGTLUAf4BKjAMPyhkW4xr0hedTwEJeo
m/RYZHrNWyU5c/GB8Oo0YzUjseiOmxVQGJkvwbxbjGYnvhO1cxiY4mpHh3UwfqmZ
iMSD7KmXN31uRHL0gYq7bcPHudwj/tAuzirHJrgwlJ+I4Zx+vAsXYk/viqqt+1+H
izbRqBUlCp7UW500d6cmLoVhAsu1s9skZfQnzg03u1a2zMk+hllbba2bQoKDXJJ7
y+fqktzytxtzxHZ1qMfOe1K6Nnnv6Kn0fuO9qAs2U8pCPjB8hTYOpIsk4HV3oEF3
uq82TEek59fRCdFSKv7YlIvpXYhWlWMC+OUN34KPiiZKmOx62fnl2Gb4Y+x6Xgcj
49K9YBkIPZjODL4qgeSXXcZavB4Smx1h+94WuFaaOPtd5/FXwfHGDIXX03OirEcb
CSiv7CmvNKrJb/YJb+37KShNr4Y/n9gXNMD89xeZ5pjJ+MpTFASnbf6rIW9ccrif
jJioEF9jnuCAddJJeGS//t3cEN0GsMX6zlREGrAhE30TpgGJbbLStjVD1znecMR9
3whzBNlOsOlH43YUGsBd1QUTm/ZBqAfDWDih11qxDLI5tQ7KfqGLqlWRAW88kx8n
3DSa8jSjywWlltXrr2vNHVXwMzyqNVmPhCl46Acjq5KUCz9lg7bU0737zeN7/TrX
1ibdbTwttlMqj61POkxC9eoHJKT3VMlkGtPVI5fDHX9u0p37x8/peqoqJLQ8Yr67
1UHS0AT32IOcbhthbdWCxsER7jfuHM5lOTRfPUAHAlBVrLFAPmSguR3HRe+3I+ZP
NxUzlbCGWFuq2KaHAWx6tjVzLh+kCelaJbt8NBvZwNUdXf+joXmybaNdliYFYzc6
o4WA2uzhTGGkzOhfIzsrVBBiPhNKoQIlswMpD0vzFrzjl3Vv8lRSeOn83QHNulmq
OUuQxNJ3BeolWMGGAIE+5BWFOGcxWeyhASkP2xjjjXEd3QEmmL26kc4gTv9nkn7Z
/O+aeimCiIjUxU8dVODSInx0xuJQNxhou/lfKYbqNXP6aKlBJGJB6XkrmSRQEFe7
LbkWgnw5omWh8ZmZVi2HBUEOmbyP6/aMlkltrGj/PxQH+cfkQNsD65rM4lIxtSlr
iMT2tAdJJtlRa8gxGW1I5Afddxf7kZ3A9k8e+BWlg1qmVWcG3TKlyp7Zd+keR/R5
zgy3Ckle7dy87y2bJ092KA0zzBVHDxp36MAh+OVRwDt70OPkNeM2vaMSfFdH5vtF
Ouw8Bp8hOCMsMDRmiqsJqZAOoFfRZfOxzFFo7EkbegemSnOIVM9Ampti10W9GumH
yqqR4ytdHzoxQPjTMl4oXxJcDs5RF+foNwZMX02dJBQCeQtCMsvFg1LeEH0dsNRF
XN6N3iwbpXYY6jVbJVJD4w0ciRm2rMH2ENtJalKtKHZ8u1cgrgz0p1QXlMr8VmKp
bNnsBDrHerFamSidiDSe1YkHcNXxSrMPexaLIGlj6dglpX6MLwCYRim09BAodwMe
11XEvg0XO3Dad26ATQ0/Vz3dWaUqWlWLT4QBr50fPEomAdkHOYkHNyN/VAzB176w
d+0Y+njFSRbzDBoeD4dEoW8Sw0j8OXBEmP6JAvMoKAZywL3aoqC4sFi8JvZh+xtF
wvuLArTX1G3iXuM2MIabJXaTRqx69/9w1Xp12HvBB8BP/aqT7HoWz2lvdZqjZ5Sn
uTokedcbqHvd0LDi017W7Cxy8dDjqF4dCAiZsEAc0QB7XB4m+LXDRp0htSjTHCyL
nRG5IBB68b8N30G4vfvtgPYmJ0dpVBQ+NI62bFOCaOtoNKtIuPr9u/6YeSEwCcLu
G+2LkFvIORELUfGhSyFjPE1Uo+TuAnKLOV3zMbsRr+oZQHl2+np7Klgk5+APkSmG
/SFPF+CoFYd5/qQ7ZR96lSUQkXgm+dldaiXouc/OLmeSGMoO2qqT2jp/8mr+q9ei
Z60qrBXFhmrVCapNRO9/B/TQX07jsjHwDY37Xrr2RU95rbhRXWsl1DlKVm/egmjO
+C0OWoNMUCjRoNlYYySMcmgDPeP1EWfQ+zYTFinl1H82O2nZaicoM3Q2cM8LOFDK
N0OtfSL1VE+ET9QuDEyrmhskVrvmbJCofwWF88oIBTw6is8mzQ2PWTi3srRw3uVT
dpCZnqYJCi9zJAjo0Bn5yvJ878nglNvDbE5XLM+a+gnUSYu+OdmaF2AQuStH1034
w4T2YLsMdGb1YtER0M/a+9i8Cwep0c+MPLvGxigKXuoqIABh9gOFkzrIRwMo1GGz
eB/PpgrlIq93/pUzatiuO9pCU0bEspGHbkc6a1wjoUXrzlTc1LaMxTNciVT+G/xO
f/RlEX/fFbHPjWvU+fpbIuwj2LeGtLskwZlnDsyUBOt/GkIGdAdKvWbmcRvN/CK9
9PePcqyTbB+3aKadVH0OIrKAUbPu8R7HCoBYij29D6JABh27HoQz8tbw7CUjdSn9
SOpoL7psHgBQ7WlSCwaoCW9ZgWgZ0+XDuRiLAklhCM+6SFfz2jloq6ZLW5xD2aMS
h8IUFFqGADxq5InabgyewuzLHYz3I87eOg/N3N1MG+sLwBmUAHvOrJZdgcieR7E/
7YTGt7vIW1iFBOtg2o2lteYkZXyDrpdP8Lmx9MwS37C32Vlp4mjrKBTGV7sCdX9N
Map1z2aC02uzmrARP03ndOpTotPYs82dkoewQLTQhzfTsVGu/um5X861dV4tau7j
4x9ZNl7p6+1K2wQyAPpJkEfGRd6ACfBeE7rhsjVvnkx7gb6gYk3VeFDmT+2eRlX4
orH7/qzljKFBj8VxAxYKA/ItSt7s/ZZfA2Ck5v0OKompu/xmdNZGhBHSC1U0yAjb
AZ7YsFtJKLjJaUoqPX5i+dDRtVHd/gXLVr2Kt3dSV78/mcTY2qu9HWSasCXuUSEV
3UAI1jfHIefIn+hsrCo43UQ+YX4RtkauMBK7ZF/41deI9O3peKUsCKWjCQMdOkO2
OpkoSGIpPlQOUoPKMYMbG1f55zJkkQ7B/H1AeN1HDp8WefuPnSUYr81qOpX3k1EZ
GWtOdaYtyq0x8qc30q+vPR+3vnq7lciajqZdBzAw7rBEmNAf2DC3c9WzrKIMp5Ar
uCM81zHY7wgtoanc+kPkagd/4rV6IzKDw3Dkt9CLMvP2xBF+U6vv3k5Vbdj/zdGl
WUIFf8NYpcTRVENPTfBc4xRMkzSbY0gyIsuuU/C8c4k42If/Pl37GHwWhS3k2BiG
mCt2EC5gHK5rLeuZOAjiUVqE0X1lPsmMbdG1NshHUY7qETW2Kn2lz90aOqzjj+c9
6sBx4LgcC0UAWJUvzJyvH5cwWSPjdDIk63wIwQ9Y53eC1wwFopn7gECca5Q7jFXE
xoB1NRs7IKjVLLKpNho7pvWaGsIglutssucjBYxIr7TTrUQhnmrQ0qrPgl6RzMFq
DvY62SrAcY3iQn1D2tr5RkoUwwxWQ/5SHGtra41lMKSnzaeEorkjXh2wezhNvC2a
9onshLI5scC3sjFHK5cDxbzkBKFYc6gQHkdcQE8WabkgbyqPe/PrabuWm/1smT/c
nc1PDJx97S+UWuaCwAdOjKUkC5pIYDWdfWm1l9o9xnGWPnygEwczIewWdug2W3nD
CN5aAGKR8n5dPvqmubD2Owvp5NKsEQWuJrv9ffH6R5CXzV6TbqWjuS1CulaYVX7/
S3e61olsI/CnRub+GmQOuCVNf2cSWRQh572cLCyH4c4O4atVdk3CPaQhROg5VF2F
ZDd1XFXh5KZsovI01NKVCrpe8Zo/9VZ2xqx+xKEQZDEtADAq1u30sleBZVnppQYW
AlcjEFnCZuW4i9XKwnH9OgvX5h/ukZQejs1tov/iXImSibL5NRVWJD6qUPtffu9F
/Bsk90yZ/tCG7ZXqEJXF1YmcD4KlXuSxK/sQ+GAp0GZhqZ+mctL5tEzi8w8eCfQr
fMpiGi6tk/m/WTkr06023krS+OUDylaCgX3yaaCFIms9SoxYm7skb3TeRIOHAMDF
B5qdbL5A8kUq+hNznqlIIDFV5+ucTVVRpw2NzZiyIGRhX+KC8WQ/YZCH0SWs61BW
1CD82sHlnTaHBdAXZldySIgQFpWOSDC183HtKXajab0tNeqaz6OLkEfbWcQi7DRA
StLarKjlMtrKPoP7JgCcqaSp/3DS3zayVjMz7oiGCZ3XXMJtVJkxbtvGGvbizfUO
zRrr7hKXLfH0AuE8FiFzJ9Qjui60B348yywVnvGErSAjFPBBxXRrNLBCe35ybTZN
+qUw3hwlaG/4ghFcTqYyhWJKeMw+FRQD5FdmSTC0wwpfvOONzWVjpgNETH6wSVaw
uxxwGwbVHnBVEA1A4qJtOCHNnteEZy/7TaqKtXwunbNxtKfKcnRykszxpRvU9QTA
1Exhr6U7ttWgFPXl7mfa2QCsyAxL20xVBZfsLmMZUjzRVeqdgd0ap8JacqzVI9la
HPjdwN5lvG8uPvF8J1tGHBO0VZQ2dj2b0Ch0sTtFljpQvupJPCVGpJcdz3k7Ta9A
vbT/xj5xIL9p0dGi2hgIpDJXH2BLy9Go/AdLLmQBn9GJi/CYSVR21H+0RvIFRr45
jLb/iRImrA+H0bwemx6EpUyXKBMHHHRl1WeLCzviG9uK11MZoxoVAgizzIIXAm3E
gKUHsasVZE/U5Au7WyFq1q3Rto/TBs1NYguDu5qr4dF2rxV4bq4nGDq33zzcR7UH
e1tp+1/LHnc4zMv6k/4gzCu25Zqev4VlqqYiG/oiCNAsv9WHgnYIGdq93jZ4yaPx
ARvxnPsQNN22mQDuKAKk0cautCO53BD/UoqFo1iP4Lc1auS9FAuYKK9xjQQr7ALX
9sxTXsGJorjq4M5ihj6sUNR/UnY4LsPi3r7VFgx4buqYURWIMnjTU+DRkqQNdbia
8bGt7oy9Azas12KpDQNqGsEPjL/CmGTgINL3oCDBvCxXT6aXDrHkzuafVY5KjOdu
JTpvSx9+h4bfP2oFoyZN95xPHuox48D5/qz4kRHG+32SZUN5RTwxk3CwRuRjaqpg
6jiNqmtjwGGEcv77NKt1vDGAvxMd5nPDDW+rJ6KpqDi26FNTe/W5SC55xZRslW9B
pWc1yyYw+Ow0KuV6op4XTSAotO956CIEFMR9OqVTEngD43+rVPaQVIwh+LWJBoQB
KBHuBLtGEpCQ0r8stvRjlrZ7+tlVXvCexSE8BVdy2yGg8rQsG5N/30PSsqCYHg1k
ew6RDcd0e0YdxbdRsdqRWJsucpbNFkUvnpgST5jEn4M4gg6IHEoAoyrn5ZhR/98+
7pgvNKXWCpx5bVOya3UAi8eax6OufjB4s4xooC7tPPTsRl9gJBxbC5OvAX3d7YAa
WtTqyDLB0I2+CytbJ7/VmLkDv0UTMHHzhMKDzb4kf8v6kyB8ENuWOMCfY9OIRz8j
FFbTdTXN9UgaxwBvZYAbaLmE4HFo/jV63iNyitjJ/gsKChnSi36zBftz3ib4b7Uv
LUieaDQTBECbs/e+5A1r8c6ewcmTg6ShgvEHSXHqwOzTnr7FffMEmCp+inFWkZXf
7uxcoN/7Qm8X/AzLpWpK+THvQR3qmh8AuqPyfwacrXymGLtFRTq96IV/qT+vvhDf
QiiIqEqjH3D7aCqMRNB7+6rAx4YAqBfcFp4f8j8Rr2miIysCrwXmIPUNnTjIH3n7
ogqPZB9lFKVl8k8UMBkzmJaEe3SiVLLuLaSpQLRr41Wqsf4PVm4iWq60uvtqdFPr
JFQyPObIXtAfAuW4lKDIVFBxFDAH0BQ0TEW2+tUnLKCyP7laTtfnX26yQIlO4scL
JBiYdjuv4dldvptNkIbsGzah6MIrz3HyK8fguwomofMVKwZQolZ5AtjpRkZn8X8D
SikV1EHljaLcO+KwvyBl4yKm76gKdrBvFGMyYRiVxOUo3S+6Ea03uQZYm5gfDroY
tsgDpvuPRjYlL8k4eL+EUcHzAEJ630kUzDBdJNgcNKnMBrMHQzmALza4FahGeTpp
dSH/d167+5FnDRZLrsOukAsT7+l9q/P7HT5cbD7UrU7aT8Fhpbjl2IFN6RzQwjcw
fyPO1iiKBcbDicT7t2uZvPB4ci1IZ6eicoKRroEGJTSblk+xWmQZSbDtqNYClYTZ
7UU+MOkmaFsJ9DU5wd4E8H12KgnC/KOukbHM9Te52Yz8fAtvWVSyyqQt6Dn/W3sT
0XQwk8bVcXubse8/qXoENxl9/63U9OktwFA83HL9Q76HNu2Cz8G8vVS2W2oVLDPl
dkfsDwlX+QJ+MKT+shEcQoytgQcM9pJfEVwqK0NP/O0ZiMPclQzmBjz0Cj29C3km
kxigk2lNRSip8yX3Z00kFOICQ/cVIedMVxeI3UOzmIMiSoLTEZJIWhAjglJ6wGNJ
UDh1pEcNbcp4r8eCqj2z0w07ku5Dqc+Xk+Ux1BmbYbo1ea4k/Oyh5WNctpT5JXF4
BlKbwAIMbG3wY6cIsofm61wrMhLCHjLjT7VlsH7EI9xwuUEICLZuBieyhPeWK6mi
NyUM2FPtII413OEVqzUNIuq0nMZU1AQDxVYbozWcdZrd/p/bFzcuMOORBqpUTx2w
6N/KV+t83fMdrAMlsaZPKWYsLOSDzowGMsU/dSr4M7dnZetYsdOPOsXlP6YqgNAs
l4kfCaFUw7EDeyU3jReBIkPT9ji2FxRwjn05ni/yQI3RaC20eU0jytPjMOWv+0Bv
Bdx4Bblr7SRcKhzTJ44KbKA9iWSsLVce/pZDBLswggStYDw2f3FFm9OYoyvw2N3b
Hy02nxXF5Jsc0dr60BFA8vMBDwQ6QKAJC340T9/kfPernSbNeOhITN0NPiD3J0VB
T0l1PeqVeKqDFLsdHlUbNnBYoQcQELRSRwxU9NBrOAp+isBIt5LFz4WQ8iTyg7Y1
2S8oTAMCiblxe+qoT38BS/Li7cGD781xrFkWLA4SH2rQkn1KWNPU4iTykpL5T7in
7OPnxkySu5QMFrpZlWJoe+0k9AH/UrnSI4FvpzmzKl0OQQh4yfj/ywQz6Apy5XT8
xMJ6D0PTu09KwKNl3JIoMiP4x1b243K9ZsiOLUoDW7kz2HHwW7zZcFtHqq/EL5kh
vYQQ44IJfC99paYG4tAgg3EOgVAcCPZggxx0hUaeMjj6MaSTNZft9ir5lnwkI5I4
ok4ofLWd5GIDst17USPqiq3rySEWkZN3BRjYDlLm/YVU1ValLguUPbbXuqu/q14M
KFCDgCJqx8pCwxoKhhOK+JTVI/LAgSHrE8/PCNRfsRXJ+R4oQkbfkwl29GLzWSyr
StsPR3spok1TUCvPGMINw5vrSJ/2X1tRZd5cxZKrE67SjbEOdr4kM/IDlj5669A8
RkZRPHmtDqJyZwGLH0sLrlodOlyv2cBNYm3z7gijUTQoxqvNQG8oKL+cgDqRURPg
fOaKdixT2a4wmU5+MKp/KWTS6ZS3KDtk8oBpOSL+MwV3YiadtO1q7KByHsDCLoKM
SEVd9oitbKpWo16/LdWyqn5yrQZly5EdQvFU5S82HHfBOaFrA/70YfeMCMbUOR2q
YUZdxQM1upSXF/iIsMCZbXxXFHgNC0c0FJ4VHmNi8+meYYmSd6IgTOXp+t9WBfzK
hyHTfQeQzkaXVaCAsYCQ6aILrs1kXOdW69Jj2Y4K21sTm6weo8E/E4b6sj3kuI+0
TeApnsZZn4l6T2G0Q6ZiVxtAdGksfMkivtTD7Ypa0MMrPmjP+lyqD28QJZXmpPgS
n/2/dyGikl8tsmgD+mFceXiXECef+TPBLH6hpXIBUaufwi6Ky9K8+DvxIY2cg9Jl
O4rloyRZkdeOCYxFbrMDKiCYG0EnvTcPw1vkccZEWdh1VrJQ9bD9hpslWo3BUfOm
iid1RGwT9F0l7iuxGnrZSvKQZeYgk0s1DRDjpOj6+xJtmxpmBbw/QEvPtCiwzldk
hzEJGP6GtIF0x3ZKmZGT5IbViLdZg/IfBRgJpshwBXmUSXQLrPlzdLo8SjIHVSQ+
G/N21CWWHh/DhczwUX6U0e6LhnLOmExO1laSefkNZ4XPGag6olqZYfJyz2QDDAYO
1nE9egUpxtVizWSL3akYqvH79wnTtg67p3S2+8wYtSJZZ05xSPUt98Ttw/lsEj3d
ZO1Ws/qb3A7lqQbEQ4qlazSHNB/AniUqjKejN8VrSPgB/ClPsiGjfjs1lf4jv7k6
K4nMZYJ2saGLXAVnApB66cB9azQkMratK+KVX+Y+0nLfTVYU+kcWoHxUhHW/NWYd
O59Pk6g4wU012jDFWZl5tCZ/b3QFV9E0hw7+EHYAX0bDRn9hzz7v3/UGaeHBr9wj
5BQKVYji+n4NNp9V0b7IkKc/NhF0aU8tcGlUF80QLNaWiqvZWP3fAtJZY9EN5eyI
lhekrFykZ97U0yJwP96oHt4bctQT7JR9WV8T56atx31kZLQY8yT2DXySrY46IfR+
LMDGJV06YwYpSSPMbkf66NtH7TalJvEr/fKBybuke7NMlEOE7Vql+S4DOLc8/WkA
UsWNJT/m95nxnalTkGXEr3bnF7D4fgDtz7rb32ID+sM3tqqMbiPIXT2NFDzut0lN
JPDx933iSOQAKQpzqfScwIdG9Rq7r55Wa8LRvwIjUUxj0MtZT3vcvEZ5Tuebn3ny
Cv3cGZ2gPN0hNnS6zvFId/d8vCLVYog4dBVBG3HdJgQ333K7c7PO6c5IlygQvwLJ
xjVtojFuORP9Ni7bbOzaXacPnX8MYNEj9zLeWuUHeH1431OpPQl/TX9AjUkR6eZK
j8DLkrEJyXUzU/zKw1lhMcepbAv+Br+UjysQhES9P61TKzF0zAEKDLx0tw4DmUZJ
k8QVYs3h6+oMmIdveBswPSobPdEmNerW2L/ulvYd4a/5hCvPHNM0sKJKFD4V0rEc
SYd/BN7FmbqkVU99AdbPw9d7o++OUGu60GyVfvTj9eUZtdqKa7Ts/YSAsj8jPUSQ
La22JZHIUwdwbJMysetMXer+QIUeHcWbhyebzn+DhdLdNhilfPpl1RvX/mNb1yns
w0cYs6HN6BhMnyqOmwKezaQs6prpjnQ8G/Dj4VIkvPBvvoIJ29uABkk0vOKiIjC0
txivX9BNCzTVz1SvscsY1pLE+LK4CY87JiXE4V90wBGHzAtF2f+JtYfh/jCal9xM
jygAxi6kF0JeoBTYkR+7fG56IOfI28BwY4kHzPuEMz5Ok7AcYCOuGS8Yb+05RjR2
wrLKqeKDUPYt45DmcTCpsIUt6UeeFiV2X54rQEUv9nNyKebQ3fTEDoCOQqoviXtb
0r4cF7tzTRXl9voRGIiy8PguLBm8lbQrZ4Q9C9oDz3wTbNZsw3Ko28Uih2hkDgfw
5RtqXM4U0R/OYJzDPB1VVXADR4D5H1unl0BVqtZtl+CZgJXFdUiQGhdENtDWVVw8
3mx0KaMMXxHPZ7KYg92HUJpFzfE8hO6Vl7pjgJlHxqdiORD9AAaUTiVij/zN+S3n
TggvCGOD+tR4HWE9yVfRC9+Dkf9XTaB2NJosKdMcXbYXS52zeTjI8qVFC55o3U9a
9MS6OsxgHcSjiIyQjanhLndjyIJS/ciT4pFvTpdBcqOYInjl4eI19fE9VybEIXlC
W/Kabo5mk6UELVikKLeEJY2y5ufcKfAO9n1bA1KNYtrHM5nPjd/gXMckZc/aCWwC
GZm77LTgW00J2WItvQbbY9bQI/B723JTn9yUQLtYe3dFUOMlXVBunc+r/Dram9j3
zd1VgBiXHU6GZoezU2+VtS5o1xUAgSfnnlbIW1c36d12N0/4gWYMTJZ19jIW/BoW
hYHpBJTf52vMEsykJEC36kDvmK+OV5IuezliJMzDmMoM0gSkN6gmgFkW2xxfajQt
vnsE85G6T8harQAVMKMSntMkbfVpJ6mW70G4ysa3BNJEJPVRmXegdWIvdy0CK/An
z8QO4YJZadDyopPkLcDDzw6N+Vcjm8nNBkIRjK9F1OlgEIJxmN9QtTa3O/qr6pmu
uFyzKcfeKqNTpb4C6J562fbwIvo6zccy0O3sVBZM8hxDVF24X3UyRiyUVL3LUKh+
3AhLxhwR+MCGA2pN1LF0/AECZHBKiNOviiJIAmNldlvidvbXdtWCqzK5TFjdGzmi
uw/7IYPm/Nh/Lty6DHPQ5NUb2XzYVkLrBa90pRC72vUmBBXbyqBEDW3qZJrF78Ke
7kTasHN3na5C/gSeGHwQJKr/DP80f16SnfpnUfGnutqtrllV91bblHTOa7p+TNhl
x4yaBszWjdWO4URu0SiNjAcF6fgUJNbvDVQVB3pHsr8apcm7Uu26LgSZiBUQbODw
D2/UkLd6o+oPALzTW7yd96j6uSN7+RZfw/XfRL/M6Fw1/Hl9ySXbg4PEB3E3dQxb
l3e9SvHHq8jslZWgqiQ9fwiOaUbdSxB+ckZ8gfdEyvG1WGirmdZmoV1stC73LkvT
QTfd5ZsOy4KFrSijdwfb3aosexZ2bbXonrrCM8kbYiicWArYrkznDJae1UzZjKA0
oTLPswhbpJ/4zvU3rtq2BfINJyN7tg8rzbxExwb+ZZbRc1+lSZiRx/+ibIZw10RY
5PjV03UfFGnvE/rupDIkJbqMh/HCfp68atTqAqN27qHE+DvEDmTzav4XdmonUYXI
4JzQD4AC4Ikvll1LCuYuqqa6Qy5By8eGDInGJEKzGVDzeu9/NxKtg8Kmm63+Dsme
pq6aoHyCRH9nFyvvFou59fbiQrq0F6mT3RmRwaIpdK3z7s47OS2hSTNnFGKieuM/
e+e+kw91OvOQN6TQ8X2DzQXJ51LUx0yjo+lHPUxcN6hPV0EDkHLZSRu6SsHCmyXt
OL80b7qZiUYkLMxnRaviL71Me6MqneeNrw370mO1D9gdzEjHNrL/lan1/WsQ01YU
64XYlm3nC2IOY4b7QfpakBsDxt1hN+2/+uinDto8vrmukO9/vHST/i8N1TlMiWN/
RKipxGveU+aaC3i5ARvZkdI7AKTQChBUsbPiDOurthRZevDPCAlsk8L9lsn1uYin
YTzWJX9dRWkn1blenZIUkM2zuK3Bx3isL+ajMhBmwn0V+3zmj9ics3UgFcuFRvPl
JsSFIK2n/FoxxM9j2pv4nXM+DQLgYabcvpyQTu/pXCISiPJm6AlE09+lyJpYxsJ/
BkIEQoWhZoVqB6KjWLLYE+Ucty8NbCY7S9fV6K77RSLp/4eXNsHIVekAbEW3JTo1
slEU2P8yRQQnhn/9q0Y5eajqITwrCXlDtDRScfBzzczb1Dta3X02At9AXDdF4ZiR
bsZHoLecatlC8a1WtmdMeh7gUgyAPgLOdLT8MRyLKo4MCdD4M16iTUBjWlyN+/kH
OKE1iwCDgniGjY+EnHxiYcYk/S97Hje8SuyGpH/GArj5+K8a5iBy421DWj1CYAeK
fq5/fz4x3R6+vR+HgReppRQLChNGXL/Y6OObWegJrYzcdmqmAcdFAJm2Ri1QnO9d
xrfpvd2TK6VziYHXvntm8AqJrAZWjA6m5N118+NcYrn/G9Jfq0RQMwYqjAW5cCGz
jEbpuv3ezN9eVUohaCb9QKYr5uFMlb7YDfOPkmwe1QZ5lfpkIkiptVEuUPkJ4B0l
76bHKJLEsH5pqIPXKp1WwCIzuz19V2Owyluzm8xjHvkauzuCZpIoHsexnUvvgMRa
4wyjsf3KkGwgA7zQDjx4ITbRE2cukrrEFjySfDfoEtYPlv5fBZX8fIlPop+fRqNH
S+W7x14+PIwzLQNeHM4eXh7/kAJnQtN1adm/eBpZvW9MIb3ySJpld4uTO8J8aqOi
RPXWxhm1UdlvbMU9gLa1xiHYWmWeMVDYqOUCdNC0KviQStZPrlbGf83EnMaWplvg
ozqkY28s/aWo4Pnbp1eR2QhJxkSPjh74LfNQCFPXdrjHfwZyhUURkrLsJGEa/p1T
bLTW80MzJxhsafrYyncfL2C8wZM2QLe0341FqT1rFhDBsYm9pMZg2q2eocqmyRos
VNFlbVQmtpmtk/3LspDJvo970vJju8iKRvAHvsIIH8DgalUoxC8vPv2D9iYQgAYL
QIvZ9Fe5tWnTs0o+ulBQvHPXlhXDIaxvmOgMGgFf8hdqs+aOsASsW0+ifOkxefBQ
+EGVw83aqHnCiSl/Y9uCJb/ktuZnOey03Mkb1EX90ha8940FKzcUSnJjaRtpWZnF
wCYH9YvoAD//wWH/rK5g8tOipcO6riwDOrjyzcx5PuBNVm9eKMcCNZNw6u604raO
bEBpl8Fo19VzSBz/A9j1N1x5XISv76lfLnAapLrjBXn1ta9TPjqSLVf9F27Iaveq
09utREi0jaWxkUKJqNMYi8C8DK5SgPbji2jqfiXxl2yGfPdPeZXVhe6yGByhYAvr
DQ5bmF+tQJPedGmkxY2zM41X98ajziFYh9r+qDutsfY+ftSX5FZ/7GqXPom6k/qV
h+uhmjKkFfapO7EwnXG2wSES3RzYN14GGxIvTq/ma8G7OVt6SUXbiVLJVS9KwUzK
oyGIIa9q6m7MPAsdiIW3FXy8G21VJy2zdxGgGcNBZMVE9bRJnUwicLT5RYHaW0ir
sXkukBdqIaz0ZUlKVz/Er8nPwZT3bU+auO6nSbVpocTYEo7nlQfvHQtaa20P8mYA
zZj+T8Dr/UD2NOecmRcYpjCNs0YoaMPE7KkPHAzC5QWgvaS1wa3r44KYkp/DrUSb
6oObL5szdsDUFVA08JLOKx4D4IYm/3aqhwUgP0SXxt88V3jHEk4mBEsBQxEK9ZUE
1td3jZCKu7IHZTmshKIIvGl+um8QW6gS/7BJu1Psdrl5A51pdrkgUeyiUh1BfmsW
ZM1+wA+i3mimOo3vTJGVgKNvdaIgLgFf9Y2MMSqS7Oehg/K5NHiTwUZpkRu8SUdW
jdmfcxMn4+SemBFEfebMNECiPIOWk4Kzq3UBPhawsjgDd1JTtGQJmTpoX31YvAub
4F2tUTt5EZQeDRbqfolcnm050ViOnLgnS1WrznRLwZ8w/WPxG9CmEjnRaMC95eKR
BCf0QRY+Ek9btN1fIAtqslowDVujJpkOp2+dPY9GOZ5pbMBN3YTmQaOUzBgl/hLB
ls2q/ppG34QlLovrXTJ7pZwtjd1GQfyQuKrwSVYOm8zBC8L/TgbU2ONKsI01u3Zi
jkBtqzX5xfdnJkWbAxuSjy5ZkCdVq/ca1LGApBb2X+l4jr4qMV7dXd+v/adj6J2M
OfPVBeftqgldLAcQQucO2765pzl8SSqCQopmrTfFj3R7kRdcc62Z3a+jqVy6/Aws
/5kpbQ9azAaOABRSoPPZ2cZ0CCQ+FTjdN0usB6mIt9dV1GwJk3+IL/NO2i3yyrvJ
0bRWoEAfMSuW8ikL87Gq3XrzkWkRYPCHAaJuh+goHALTU0C+/oKw1he8xGnBUoX0
f1wrulSumCWvswi+Efi/eP7yL+A49M4RwHNn3aqqQifKrdAv/QXIJueNC6KMDtQZ
YUm1bXMHSKoyKPBeLXrZHbxdK2+WYQcoeE1UYTxRn4hdGZNxF7+BjIzN8k2dwp/U
+To/bGYRftnLDvyoARGzA3ffXrt1wD4eAuTS+P+k5xBBGZYesF07neIDMD2MlWaC
y0HDh+SOdIFLRorunjwU8Sy1y55ITmso0FspKNdTlU3IP9SBoAQHKiJt3sXLB7hl
dqXirCRGCJXdwdbUQ1QvR10Q+i9uaq6TWltlWYcT96+Ws0Hrw3bEAOdZsu6Y83rT
4MtZmYcPtEeczR3eKI1TaTUc/zElmJj2NcunWSduT7oHpXLobsb0cJiDeGOIytq6
RY6HPacv6gRF7ClGItc01OKhYLgEw5yQg0z9qV6uR+eUtP1C7sOr6Wqy9bM+KymN
Hyb5yknWcDeP3ZsJW/Pdl1aSHi8x9Tn3F8xnApSR7t5KEMWmTqEZuWCat1UoqpUO
34Jmz5jeEddtAmnyrIiGrCdmU0KmKA6DjX8UWztwTuUmdYNQZ6ko78pb2d/+LGfB
saCiSi0hm+rCNMH3R+b5r3xSzj5qLLfhFQngcCyTBhcBcvKPSdIkUECrTdnzg6M8
MBBJxuSd4d4l62nYwQ7MaE5p5NEzfiOVCnGPtBlgqFGViXjF80C+/wcZDgnTXjbY
Q7rEkG7K3arbyIyJT/rmhfoxFlNq9TJzP3AIc0dGUeOFizMDALMkE3qwdV32IAeo
kHvRY0pwPITRx/Z+IcD+URvhy5Dc1QFMsWqdnVqlnjx2AVO2QFOfNVFjWK3HQiwQ
4QqqZyzMi+r8nNGAq6dBlzn2gfPvQda0Z9GS2jCSeW5u1JkAprHYsy94h8F/pkgb
4R5MLlZR8CC2c3koz5+cAAoSlyOQeh2iv/F+YHvJ6lhAn5M7Iz4eksBgSFtO/MhO
0RcQTcgxlnFOnbX1LcFgEd9KYSATtpElEg90DdHlDqTDcMwKPOg3eSZHeE3hKXg1
dJO2/HBVciIzOc7NBIyn7LYomDvoXhjJOoD3H+ojeo1kA4vORJYVkWbP2fVleoaR
cU2ot8ArMXlSrHmnmKAeEpUPyDwzeeZCvQEDXer5PBK1XuZ+q5OAdRxW35W6Xt+M
zz1Q6StHxeWVkh2XcVxDMjnOQpKZYSVV2Jj0Co4JYoX6LL4dCHzo40H6L0g5lF64
geEIG7iDnfwwPQSwu4k94zlr0FW7JsXjlIyP4jyHyz7OSK6ZEKRg1eiNfDKu3lsR
58vIt89rNekUrHb9XWsb148eeMT+yX4SCKEzWvGB2p5Io/4WilR8yYa2VzPuPfws
6qJyNyRFWSlrU8FMC+2N6dyYrux2AjJ1SQID5uwkr55XCB3fU/St6MCxM3Z3d+qR
xs8NYJhwCg7DwMmg92CmM/CJAgJ3DWud/Ho0CwdWM+x1hdq6O/7QuZ1ThFqiTOZA
8l2AydGW3Pme30CA0EiWvjDc3GelA/XfWeeToQqjliRheG74pHEulF/jifJB8jIx
7ZvaeUAugEO9PcWzjYaO2IcRiYmk/P8OtyM30V0R8dK0zyDnecJhtXKwncIOGlba
Cofv0thn0QJOQulC8L02WYxUQw7fbkLXZJi/LcDKp9g2TyCbCfJAfeRozGqXORZ6
Py6iafb487x9Lk8vaIuWxZQ1RCNHNa3R1AbEx9d9ZpFZO3BqDvUsFdRSefCUWyPf
8CzQo9akOtGQ2W7VNc0lbytUmmi7osB83OnrmTk/OarRQ6GUa1qJZ3GCgUgwpxjY
XJXqOCqCnz/mF1Cek9k9eKSbQ/c+53T44xV8WgD9OViom3UydUIbN21WRDexODSA
eoM4+rd3gu/K4A1Qd9MgQUOPwh1fE74g24KvKD9WAkKuBLTytWNY659/LXm1hQCw
17RPd1gcyU93uFKTwulD/6brFklNT0ONLK5W4Y908/I507wBFIjS1r81SazJl7lR
sNB225km3LJi2ITDSB5IRgClWc5kj2xMAAmF4I5tu6D3bPbieo3g7j68EMe64TOW
WvTK00SzXEpNBu/NDC29UsBGhuRQKACvMFPB40qOhR66B+SFkJuWvkE0wa8oTd0N
syNjFHxosRvFHhKOge5SoLbptLV6C+0V+T/XGMsCIv2muCU/HpHFSHqSqTRdkNWo
SY/ZGOD8KdFCIeq+oV/MVS9hbWVOPGxSxeKfJlNGDpvCsGSJ9SKoYYcVFZsQExH1
8wqeRbxuXR6LS8pgYgc/Gy3yqHcK/b3AltV6IaFqttsg79kDVLURwpglWpt5pkmt
Cb2WBxGG5L37JbpmzPFPGP2pkPuEnemgKU1QRDQILKmlwp6Owcfy8/4Hw71pkefp
1dNPMkLrRhfFDS0tJz2QFwXPnVa90tkJlCb66n4PgwFkZd0Z7eDIlwk7LAXIV5Di
G3vE0ttqBlAZhMuN3h8xv0oh4k4UD3ZPKRbVL72PnBOiBUQfAIURGcu8o9vz+XMo
H4D6gMqc2DgMorIMAqH8GtQ4IPp9vE/ojbUHzeAUQxWv30soFixAiZoS1IFlXA6u
vhkm5PKyHwsjR51Q4xbTcNKpRCyJ9qC2uYkulxEaSJnxRZnwMCwsH3qvubX+PpGr
L7IVMINckzNfst83eIPwmocbJsgY7BymilLCNcsuRMYu7GYxs9pbAeNrn7ewdgbt
p3u17KmbgmPfpRqFf/7byryMoFqaVNJ6ID36PC3+8CpvO6y6WXXztiWt0Q11XWT8
az/Sx0oR6L4IV0HsLkFeKpg+DnqyQ7DPz0pAKm+1WYAFnHgoSZ025QhYPtwk6aLT
qK9m3wta/us2GCMM7nrrvOEXavslBKnnN+qEoPfvS8nm22ir/9iRoSHHmEc9zmjp
MkvDnCo0xGBctqQmVsRUQyHhBZsXZF5zogPSdr8ldBlHZpE3eMnduIVC9YHP03mY
oEbj69IIXATNCh8w8hVw61I9U6Xmmqjelz3/V+pUlQKl0RsxMiSbpxQU90XRxLDB
xVUU3PUY+OiGg4yvwgnfbr1Gjc41AxSrryBAwK+KQlO9dSYhKp/GHYoBlrfGJHZ3
gvZY0PwbePxDPUBs/DZ9oUaWGP4cSJFRdI5Koy5unS+5w0Q5+8/Q0ppnxZ08IJpa
Rs+z+HLrf2TTGrArKCdydrfjZSWBAKq0u4JWocK07lA7umWN1cK96TolT29gFAh6
wdSJbNyrOHPcB7gNdyUsuvN0bj3h6m5/j3X0OyAqsC6AsCgtFC2RchHFMrB0PxCz
Gca4Yh+AZ/uSHBE7P9xqxM1CamhWsgvjqnTzJDDpVs5ag0rk69iqA+fEVFcZ3ioT
Jt4ji41Qn9XH63AHTwBd7hA/L5V7ziI1jdUfGan8HVgVWbVngMMuKcoyri8EXvaX
vccFtCg1LX6qrCtUmpy/Jo/2ttmar5RRAS9joavaj0N47+HgF/xSpaPhH4MaIfsI
0K+aLnRCzettkaaVAP9bDLR2q4CFaeFoJyrsy4Ws6zj5QwN93+Wj1pTKA9bGjSDC
HjqI7aPRjfDkneBVfdIEbNv2hkW9k1+mXS7EGlYgAWpDvtdJPpQkpYJvUJ+pG2jB
og5jngZzMdzMcvmrSX5PjBpSPp1YhMoR1lOu4lLVQutVegdt/gZxnpvwZzhoa8U2
vkV2aorTMfQYoHU5m0IWQhNTel0TngtJqttpceDBWa2jQLYaZRa7ruEejK5w23Jp
qT7+z9/uihMEJMB+u3yR690rJ2JqG8sUaMn6EKDEujm4cGqIJP1oDujcmwdhfFM0
2t3WHrdIPAxVJtUsOIDpIIoLqBzbT81Bjzeq7FWkKZOtNCsejU2qvZjnlVmAIl9l
pgU7Pt8aCoJYQwVr+HIkfR6pFyUdzzQ/MMo3ADD2QFS+BlMHEujTNIv9j0OBeN/6
UaGEaAILcqlTiasLRPEzXa9qgV0yIlb/2En0/Spq6Tjss1mczxN+aNBHy3PbKQDr
DLQEB+sZXEVNe+T1EFGyjGoeM6Yow/iIauSxyUU3BoiMtXuqtc/mS6Z3wSiMSStZ
W+cMudWi7RGoGhmNop5Tm4+zmSMHxZSG+WdNSqjdMk1Mg0WFQrVLetVRNIa/BbpG
2KsDM/WuL3ha+DTSRnjQ/DPSQIcrSNZaH8mqkJ+TaPAhf56GS0042VzfR9zrRf8O
T88XhSKs/xRpNpblp7SaoZPOCEi3Dm6e/O4F0Iibj8f8afPj5w3UMe2ehKTyHjSr
ST101rzNSePuSmu7AntcGGELmP5UfMbLDQ1ZGeN00wNLXJUcp4Up8pQ2LlLuliTE
/mCGGH0cyVvq9s61gXIVB43CaikBY8yd/I3O2jJJoXwbEXKn+yZG7avCcGqIs5+L
H8OQq5FFqvmT9A6sM7Zs9vD0zqg0bjior8g+U1OqGWqd1bHzp/oZsN0E1ZX/jUUv
7XUyMI/le9eI/n2WNgPd5DhuECn2f3V/uB25qtZpmoIdy7OgfoCX6pZ/mf7HUZX8
mZrnPMEG9b7plfyYxODQETseTUOcRTyZO0qFI5sI2AQeVnTqUVdGe+w4kqFXptpY
t7IJRL8Qn760ea8T2K30o8VIE0I88sUsScTH//W2yZN3mcE9GaYwtls0Nw83Fwuj
H4zslWvEHlK+7bwyv/gWrLR5Lartwd6cGPFF78yOk2yMFGCTGdVB6uRpkPy2baen
OJNPJS+mFXX5MGlO0qbowTqDt3WGI0jOmF5jG97ZDjT52WI/L4WQgXMmPoCH7lZA
OdsjPyOMf8IKaF8gbsxdJVr4qQKt6kMk78r8oFCUp9pVEgo3fUizNjd5l8A7zOfz
j0GwrOOjxOQc7O06m94U47xCdxPGNwZdrpet3HOteB2fcfPYA1OJHtb7utgarj75
4vXrxh5dWi8KkOBWDBZfsfKTHVxiantmXx8loZ3CQPP+aX1gwhVZ+iMCgxPh1xhz
BHYzl1ZMA/iBk49bFSSo9Qn/w4V0XT02PeADxvcb/Znv/Bu3+Q2c940d2zzm+IPr
Qdc5OvZovaU3hYm/mQgNLq5QE7SE2OkpjQKJQa4RsmX/wh6tYuGoId3ait2jCfIm
FKSTW502SIqseIZjysuR6GvD7euK9pyaV85gjBIr6q21XCvcGj4tf58XM7K3E8I/
6MIQo/T9h3tx2XRBp6/IHOmLShGaao0NBwexr7jUXileJihKPfjcydvWHHcisQpa
V8w/w7NManXCaV1btfk7bt6JBTkdSOLvIbOqdmCy5ytOTBYIdSWeClqHMuslGk7n
lyDCiASfbNeMC6ZVCpv15sR3DH6K3mhu9uvbec2sB9xlfW3tYKGKzFquXI9UMyjV
jbvTXNfqvZ59HPyUvhl3TkZzpOM4rmd7ezYEnAHkeexzjLEvic4Hal1EjUgEWI5d
FW6MN9tCkHf/73PxT6G7qfAyMkmTNcP3JUEmJLeybRZMskKhJicKBfM5npuOWC3J
shjTACfjpP2ZPwCzdEL3Qce5DuREU3plr65mjDfea0HbB1iNKJ/0Bc+VcNaGGWuX
gjIzvVMS3dHkFUWe8DDZwDrdFX6jMdnVlFOfqeQ3KVNEv9j377wZ/Eb/3Dfvpe3h
Rt5bAldQfP/ZTiq08a0BRiXOhs0A1C9AhcmoCTi6TXprIfD3Lht1TDkvfQrPBiSG
OG6bCKP3pLk6xChoV0RHo3jqIk2FJ8dl+j5c+QpTMAGniBP32tu1orbKGqHaPTLN
kQyCjFMTGt51lKBezoE2ndr1fjB4Z6dTh6zChmP0Xf55NCkG7oM57pKvS5AhFznq
h0BqQTDqVbtIC4Vg0NBNF6AFMaQynJY9j/UIapNULbAAtrLA9izhteDInSt1ceAw
73rHt3uF/Yme8lSkYXdUM0wMbgecVexoEk6Bag2ponFhSc5qU9na5diIDZEaEL17
8Idm+6AvVJBlf17i2O/8e+Y+J+laNiQtjuHVlbiOrCcui9Q4JqPq+rrBw6bhdslD
KqW0R04Hh1lAmnOrVJZO5/wp0iY9kGumLzLaxJMbkTQP8bndpmo1ycEq7cB708pc
Ml1uPZ3PeDQfgT/Ll56Lw4yaceWHNaso3r1H9Sq/7zEwrkNYg+X6KBnvZECWRZZ7
n7MX2AwHyrPd1wPDbO83B5MflYXV7J2cl/0pS98Y59gOfNt1KH0cejVBK83ShJ//
av+7b2I99J7zyeuE0A1ymCd0WFzdUHq7AU6e0OkYIgaULzOS7XzKD5ESSA7KFZqj
iMncCvqyev0V55z/Gi+MZ5TRSxuhQTlol60atdoNotMArKIkoBbscVuMTH68dxg9
EttLuFeW9zKE/Ioje5yyYXQCxfKlqySOzvpEiRwPhF02c3Tkv9v7TGCjj5+NDpXc
GJ3x+4BJiiFjChOY9SuF7uke1Q9mAWJ7k4R5nb/AxHk/U7UfiXRlgAuKbfYbW2+z
j5rB4urcFBlyyfkKRdqOT7Zqd5RchgGEA8272AW3pZY+h4RnyPzw0sLUX3XC/Tkt
XM+WY9W26pi5dRlJqjQei6IhrQhTp/PsniVhqHmOXNhxhS4rHNqLVee2gKFTRwZt
3VAEBLS5UTC30vFuVf20NHC97mHU/aQZt0ircjMY6Ycbx1e0sg0lcbrb9FuMuwkj
VoWd4B49lVz3fNcMELokLjI0Jqu5ZML77ovkc2sXtKXlNEAMdifKm0Rdast8Y5Sb
A8Do62ZhubXbcMkj7zTZWB+BlG3nFnTclQYpO8TN03wxAHUg8XWsPgscIW7YPWUC
ADmT0R/jAr+GRNngem/7PNM9pTNiOiDMBvjuB2i7QIXIgskTGK8mJ7sDhAF+tsLc
zERgjhPPd9eE/dWmwftTS6ojyaZhmKpK/LYU0JdfJUezUlMNXt7CTNw2edU9kzP3
qeECKvZrPlZdR8wOv3m64AZhF55vzmVW9l5SDUkxCUtuNzOqA9PW7BDxqOzeXnHe
9K+b+PIuU7Ubajbld5oeERZDU39tlmWbl8x63JY7H43ycc2M7wcwzuExpBOdL70T
DSx956u8M/2a7nZo1GxqtGZVR+gv6/+rEtyw/3BlchgeaRkRIHO21imDYWmAjyFZ
0Ir9oMV276aUmvU1L0o0t7hG8uvGTJPVHFQ5vmxCNxQCTaok4xL4cz8VDzZZIyPx
NpHM3h1Kh80ixOnvtFhv3Z8ouw/jAM5HrcAD8PqxPtQTUAirTJdQGeAuHo0gQ3AO
Kq40McL7KoDIXqT0RKxNlZljZuQGaJscgVmOGt3F0k8DR4A580mequWbFBPp8JmQ
dGKcYzgBsGGdTX+xlRhcqlHv6f/8yJE2noz1UwiiBX37hBBaVHUCyXTc7MVMNS9N
5m0P1B2hduQTdAdB04HAO9H7DOy2RVzFpa7bnbmH7+dF8e2WfvKpvRlmPbOQ0142
P0KzpgamLSYwJr6O0g6D3XPmuwUj3f8tB163LSDfsEgm5JRZdBcDnRlcVz143YOz
jXAjeAw3QZL3xLaejBkRA8fKTrVRXmEcfeD9Z/6wyX6hC6qaJ0P+RCugJxsI0pGS
skcd10pPwTDZHNn59NR+Lso0h7/+kNNikTY6In15nLWBXL2ci49P4CifzjJrRhig
CJmlA3iOmMQ+Yvqe2aoM+SvVipwSoNGsURZ/iOZftt1ZdQAHLfT8ZLUs3i1Cw0WM
GnVV2c5dlQyjUTcRvSXgg2n3wfIFjEq73k2ABkEuezASZA8Ew98MrDOEFm44Tozr
quNm/ZQOMLwy0knGnfh6/2WF+N7S/2aUMy2HmyMU/ifqiWUHfLIBVr5wGtQpC7o3
zRdnEqWhVAXE4nehZiFODuNKhengNQkaiq06l0pN9XcVoGgrPqvvGAO1oVDPHlBZ
xAkJ6p1ZpyjT+QwfiL7ihamsqGnZ+HWLAeZvpoBC4InFb2j9htO/sCFce4pzAhyT
PiV9/3Z1QIVjNLp9MVt4QPJrRm7r2sqEiufs7I1K6CRINYzX4jPNsGkdYas5tNGa
mgkgyiRACMt51TcO/izUk80D4qi8W9ImtHbUi/kcUgrFlL5bEtx7BKzMry8++YYd
oaEj8D+O3Xhvu96Ww455oZ0QN4qlmL+nE3cQpAoMwlatqjL4mmDPiVGJ7IHdlPiH
Fv2ZYcSHqMcIYE9fIt5TYdhG8mb8OMTsK9rCCTiMriHOMuVh+8xVIqnts2ZnD0bI
1tNdpjHHpFAQTj2l80DWrAtO4XwisWhHeJV9rTD5RX3MmJio+xzCLer9taxLInSl
MVJjnc1xb+gUf9sEOuW8yt5kBOnrUHhHupgFd+TV/ehZqtII6uXE8hgSp4+GoPGg
kMgslzun32hXRM/1zOnEg8M2qZ9o5EhOukwV+kK1zgUvhwIE2bdStAJ4fsKWNLoc
+m5X3ycqyBe6WfJzPkhY9ZqrV8hCM+ihYFamLRRvmO9KnofcxuoaVf9OpnHrZ4A8
Qrc41IH4EvBlA7+e4Fg++INPQL/hldFi3khBlGmKWY/d+fGSL7K/kJmhpcAzxRz3
YQXwQklUElE46OQuhnUGB/3t/y5559dHXvDi+hsfaFH0lAE+F1VfNGoxfpZjb8pz
LNSTVr2JCWTYzZIn2fGPh15pSlbR1G7bveWJs2r4eKgilBOI9/sN0ros/Co0TtNh
lDylcPC+VBqksSJqLtdgu3l0XNHEe2aAuXOIAv/n5vcu2beCIO1cs+ENHzZ2t5j9
8P6djQSJ6XtA+do8TR/6T9ymje+iq0HYjXcsY4rCpNx+pkHZ25ZHJiUpf9sV9KZz
7njbcAad68P7qb0iWRt+a8Rh2ujeog76I9UCL30GfwxwGtS1lkSoiMdqs+6FOZEr
aZAuB5cLOeGoyZcUhqwX7FmBQYd/T/YRJhGX+eqk8gKRAhNxi1K6mzSVmbzOERxW
vffY6zZHXLYsDRg5INYCqBRB2QoiF4bq9dSwXedfPve84CwViPWoxRwlIlWEUtQL
V8CDHHizDKWReVw/zlOunURtH9Isw60Mr5r3Si+jO3ScaSckWgymdw2SZ0i8ptfg
YI1GB+YofjZQDad9P7g1oTDQdww1LKaDG22KtZNo52LUCoYS2Te5aytyUIfNFPoY
bVt4L3JQArmdtG9rV8q5+BrIpzf+AHqP3JPC7vTAuohzQhupFaZRYp46OTfhHnIK
wzw7Crwdcr4c9nCs5LCbZkUpJrO+LwDoXChz3HRfhmcXUBJciuV+i9nq5uyLH3sh
1Cji5f4MZjNlXTmx4/SU3omQcVXheDaoPjLxj317RcR39bxqcaUQXOdFIBC53ZdW
ZzjKt3zpgiD24cgaUqpywF7gPpyNBUuAWuXIijZUNZ8nsFMxrA8lTeFxr/rIiTQl
/OjX+PZNxfsIhzORv+Rn8v1Nu153yKSdg9UnW+YldCpICxinwFWcvg84hkCkJmj/
4FsGRkiVzxGoVUthq2mhrdlmlZNssUznHMwn+89yHMUOLHyvgT1GsBF936BYmcCk
S7b4OmH0YQzzDZ85mjWMZe9lYBezb2iDMo+ff21iY7/p17TW7pSPPsifvEe8H8rN
lwrIjinwfxGQSNAh5CCJMLSxyB3LWJyhbyC4RzUlpEQmQFDGX1vhnixiHRsl6kz1
3doLJKHQOC/ipkNeVNG75VVknlw/eJyEoQMd79lkR+WU4OT6jzC6sP3UlGEF5++s
t6q49EXbInM8EF7E9JqHe10WubugxXGqz7omi4ODtlyqEnrraGbq+6JjTdnWKWaz
p928e5mclOZ9V07F/MGiXflcXJiCVnjZ8XI5E5oYh+xmowwNqH0Sg4mvnxCzYTKE
COg6ikFnj+uux+p+BDbJp8Xcq4jtcpnBstWfQaGB9f7h1vClnr8hZM1IQuqFqjX5
pFnItrPItCb2sKT7Bwiuc1vrncQmBLLiI2qvMOa8Q9bQB9tuFeE/aKaw1oTvpvAn
XKmkqWRZv4dCspR2LYFB4jdjMkXVKmTgstynZl0uYXO+gHbvRKG5mRX1c8peI6DQ
TljktLqqESqHlW9B9VI6qTn5mwaAf/NoweOJBkkcMppnI5/PBPVTeHloSsSlSSLa
DquNGgmQHbcbVf+pE0qTeylHN6qbJ49dH8HoKQNq/JMK2mNrzbOt/SolPmIABS1r
T+g3SuN4UhdP63TQ1ZNyLNw5xst9004Jym9TBY3/aCdtQd8OIqfVCq4/Sbfl7n0U
kdNSETX/TnciOZMx86YrC8CvKqEhmDdZgH6wjfH50BEbmiA9fzpRci/SYtSSgZhw
uTlHFz14xDekElm/lGrkdBhwoKG1LRfPCBh4o5m8iqThUNriQSD0PeNCx7scAhBd
dQiLz/zVkLlC5cnhye6bWAe+Nwqafk9JEAWQWgUb1z6Nz4KDRLLVvPJHIVx2r0Bg
CVNRnwHG1hQd+WmhaoBLZ10kEWFeBZ14CdAdkvyQhf8IUAWa6zc3qkC4vE0U4t8b
7dVqaBd8jJj/5n/GSK47WfhLhvyb1//jpluMwW9Kk2pX4LOOp2Se5wDscOY6e8CH
HlRhD4u/Pw2BRuE2RBCJ5sMpbkyBISY9a4VfH0KlPGeKPCw2WdkL0Z6OC84czGkw
Bpu+TV7tZzrQ3kfSzM7ca0aGj4VQYYO4KK94BqNORSfwa5DvCsRVYp3zYBA6dBKw
RHOeFWgnbZGkpPE6Um0kOtXF7DQ5HdW/BgM+jmmLRkl4OPH5vnnmHKtJYrxYSiOt
ytEBzRNwFm1zmHc2z3YeZxRVxkPFhW1iNNo/PNFluDLdEIE76D+RCx3+xm1H8+62
cy7xV+hlIAl9J8WJdSJ2hStFEZCBSp+gzFqeiX7j5+jViUDNm+s06iWZ2m1Vy2ZI
gzsWdl0thG2C2R0zp4Kt6v588NPBzAQpUziaw810+fvLtefAXKDYYJ+LkL3+JnUt
k9mTqAewANqqwg1O6vWsCLXn4a85nVcKCEVdQq9R34wS5nyyUxSQ0R9UNDbPqVaU
qmuLfHNCNF8aQDp0s4/8DZILaoLfbVFcM2hg08XY9iEhhRw5svMuyUT7svsjiTXq
IYtwnBF7DqQicX25q/9iDrL2uD4TuRi4H/f11C2KRGamdU/Pc0aY961oJevaDgif
76xoLi8jeuG1HSsKLD6Q1Ifm/8E97NMVfypVh9IAg+2LE2GtnRfDl7OqviUixWzq
qXZeCRXHbFdO114wXcgCVdE3jnVL89FWEDgP7Ew9s/OQ4Ngfx4C4kGFjR4dhRAlL
Mulor/9ixZrQsRLl70CYvc/G6IN+GLqpHv+udYs7MBAPWQkCqizyPUs6h8me5yFC
njiDYAQS+7AzR6P9+ENQu1STs7aQRRbbX3ED/iLffZjv+6/A/RcZM5McGw+bWMot
pEdTr9ze8mIzJruIqPE4aeiGlt0B+DTpQmA5ZXWNz+gDajcKb1g1fboFtqHRTleq
fDYOBEdBNauIrSMBoJF7ZnObJ48eiECGIffOd5gkFEZbJuhxvdzgj3r6DMkYj7Sc
pa6Od8Jr0IhqBQ1k+gbEpqOoJDd9F3OmUk/kyg+GjRrF1WJAGNPK36ZjrtEShtmQ
m95+F/kjdNNKujuiK9m1Vat6F4GnG1smgkWtZXT7345lSPW3e4dsbWyNsHV/Kr/I
3k3MFUPopA6BOAovJDLewGcoNZ1UoGtz6SFncBCIKrZET64LhBZAWnhOfMZPXONv
xaRXc0GI4PJtM4BF53SL1Ew3qjcFTmnvZiQGB9T2E4OjGhatBCEg6yJD00vRyJxw
FJrxH0DDzeN+rQbDpk0sh8bUMMPIIzEt24i/w7o0kLum3/nRxUjjofS2TUinhHBG
nFq/ErSEFE6E8Qfj+QyOpNkH5xdxK93yrINjFChgyq/8CxZcnNr8H1EVgTV97dx1
QXU4n4Lety7BU/LFTFfmMTnnYosXKBXZ+mPx1748uV0wXlQLhiCVW1GvTUkAz7h7
TzN0SyMu6s9pbmNVNv8F3Nj2WRbcCGNwtsCdJsWhHLHqM8n3QYpEyK1GzQnnPgmN
iPUZXb4Yc6Masy9kOnFmSxqUWVeEBasPQkDTj6LNPX8PIT0td2A9OrHJaPekRTIV
VHYEUrEva0D2+WeANPOe6NeKSJUr9QEXmSGZYBcuJ2tRiqjN5MM76WZTszZcEaxd
E5tt0+VAdI9sfGJJaTaNeg9VhBgRLpevueprFl2DYwQIyT4z26MIus8AXaSCBQpq
cWxqg0vGmnMoTzRw25836wYFSrxjc+MuJTuSxpHLyF2hHxsybdaoo4P+ueHbhOfZ
eqznD2fI6wrMrDg7Txk8WQ60Hnm6MxNja6O09VdzYYbALCFrGx44dcWAt7lxO6mE
Yfn16w40PTDN8N1KUSVDIc0cBQtQP7P6+4enX4WCf1UOhTaDP1bFPyJ6SLYWP+gD
RzrPeDNAfTgOAEu8734IwsgWeIH/yGsUmn9JNewltXKCrLgCUJUCaHsr8L5MCpC0
7GDpz2AhYQdiccQDCYmW13WNshqdbWkZEORWf7qm3CYltOlf9a3V8ww9ffKfKpWn
u0DRchkfwGOKD6VOIwvIimeAGYIk/NLgjTLX4iWxeYSk605mOdouG8EhJ/H7yefj
QFy/EWBjLkay2MCsBAWdvFJ/Dv7XdLWvYIoVPgq4goLmQ2tKnf5UQQ6lomQzIHyl
RiiGGG/VqxvUVFPmjaLVuLb+ka0uofFnNU0oZbXYg+MeqKxinWdG7WEmK7VT6wKv
ZMemmnUXuQmmsqGuBhPlqpevbIWHf+UYfP6aFzE4idXlfpGwFkzFV1TCfOsHwHnQ
4RkA41IozjleB7LHbu+r43Qipk0EQX/b1QInFjtDk1J4i5Oz4YMgB9rayhMNM0WG
IuKIiJh1dXV2evDkFj77RJtJ+SxQpNPhJd7JFxlgMIG2MFTgMy+WZd1iDvO2wuFm
Iod5poVkEzdZtjesL/WsX0NAx7O7PIU84Cg+8EtDAkRQhg6BMyQcw3t5IgwOrXZZ
60xLncZy3jpkY3RdcOzKfqXF5Zq2EWr3u0mOkXijydzstlRX+PSqz9+4uNgH4xUn
DMax1IEjd+ccFS85NNa2Kes7xihzlsCmK1mGuCHAfro2l7g8lUMcws0SOWnNs9pi
ZNAhQlaqiGlX7k7r0zEiX6MTiRuwRRi3hD7do4NzA1mXG7lltrEn2HmG6XCUj8zo
MFpaUY7x5VJ9BOQZeGiHTry79G1uaQdRNJyni4T/GF2hBcRBjk49+GLVbMPW50ng
64ptBIryG/opVoHMnsFtPwhJ7G2lFqNJHmoaP9t/AgLLd7yELtl5ekMjftsepSGE
OmmL6uh1qXPozuXYClaHeeNq3whNr/EgHGRjqbeeGhgBEKtac62/kMjcCeSlN6Dl
wzMoyvAPZ+L69e+OllXZpovC2+1elFdq9KrPzu0Aa1Za7JZdJsZn8bDCfhX87oD0
9fRbHiEE2+fTDcPUX4NVhLiZFDSJfeHDIXanPAr5Vik3TvGm8SZ5EWOA6nUsj+kO
Xb8nG3HkViFACjdOefLwoAqOfkea13qg9Dk0QwYvIhOJjWeHm1eS8GnvR5NC+2HK
gDRXr7eDl/6FrCD7wB9ZqOA7lI7jMWjZwVHFyYCkkoFIX3CpnxCVTqfzckykoxTb
VzAqgIUauXa/QNdWmzv6VqtDzPBhmznnz/cZhccOqEGq9dK5ZZAnnZAuRW2M/YEk
xhWviNdqIZDaHKJI01jD58oTpYhdWJn5LTWA3h+o2sc53Nr2TsfY9f2CmiN9CQUx
BNxMm11wWJD9QVz87Z+/eiGLjos+vgNjY4iqwUqoJn/TUEDLKtjvNGqBYFuwOH4j
k3Z7evpzK+8RIj1qA4Oa4sfrcjtybGq9/RaOXjeokzCxm/IzRQon6FbuGsE90Fd5
N5RgM8efQFzZEY1q42pNR+00Qv7YwPYYfqazHpQORfCpp4PyZdkLMVTmFhi/dSwv
KlS+5nofboOogZenp/c8l9NlUsyvEhikNA62gtdBBbKW8URp8ztSpci9ud8GFG1G
s0vcj0PV+DOn2StiC0cNH8XZ/rMzOSmAOwUTQAtbu2mk/c5t3Ju64Moxfq9QGaa7
YghBi74fC/BYvX5mxbGx9n8D2aaaojPJqVLtmkFn5cDqQGkCne74JUuIBvlug7Vd
xH8Nl0YH0nBkIvzbn9PAwydld8Ym+lsd762dZwFMSGhJ5tLTfbVzQBPneRzXk1Lg
cmRp60PAsBjmaQSrR0Ci5UspMYD6PlMiWannwa6BCRyVAdYfuaoxfr9enXp7LWoI
qdhKRRYajM3p6ADYOe7jDXxy2i9Ljy4PU+edJuJBLbBz9z2lifSRHLcgIfEedi8W
GETpU/7RMXaKg5Z3d9l07wlYxpPm5UAhRAuUY3lWpwFiciJwABSodRjUGdDOGcFw
Qpm33hKZpGKjpgm6Sc0ECe2qeilwggFtWI3mpoCHWDs8d66krXD6DUMCgrcofC4K
1xOPZDxEy7BhAvLlqXo161X+OE1w7YyinzCSxo+b5Mn0O8GmkUWycHedVPjGIGkJ
l8MN6rVK1nGjFZ1EYIjH504Lrg9DX+b04ZFxhBJO5dcBzFO5UPApxo9xrIzSbNef
Xpa2IKjNN9M/xuDCBpVydDIpFtdWlYIgmGeF+fmB1yuA3XVMkpNSewDYSCenLx9N
EG5p2OTWch/73upyQwTBYsl3dWJni66atn5RsXzTuEiG7/8ks10npBa97iWok89s
5khPC/9YqcnyEQkyStR2O9HAv/e67dEE9IvDzx8ugVafCgb2KKFQ98uvWwiWSPX7
CYg9sLnxSGR+bQo6xhecrfqs/0YdThkU6Olw0mL5gZOOnMhce3H6Yahe2Y0S9WRZ
4notfJ4SCww+mH7TG1fEagGRkXkOon5/JNo9Zg2mrlhiGphdWaKQmZvufINox0s5
6rmoyXxsWSQC6sTcpSX2C80PdDLDNdsmj+1QU+u/3bA2Topa0CpsjmxRwDmPnZkS
I5ShXITA1DDCI6DmwEuZwIaZ9Vr2OxNShgXDCzwU4gmjSVb24D6Krtw7izuSUs55
gvP35NIy8Ls9CDxLnJjjoU5OLWcmVXzlXac7fZPnBSbOlSal7+3BUOeuc0J7B1T4
8796/xSE6IN7LUL7Ihw4BLCZVacWkjZPBW1/wbnGc3U4V1SAqxB5vqLXfHxq0sG8
Y496pHAF1h6+wVCXObcejXY8PoJ9XtS9AZvhz6xD/Kc45p2kVbj1IE99fASqZBgQ
ghJNG223p5ZYvtP/tHcDbpG6JMlO2qqkawMtdj4SVM1lGYpt2MJN6eK9UzSzE8/2
Gx5W1RjGHG0DGkzhlma+AIn9lNc9pNpoYZpp9hIQrT/VxdiSpkFYmEoTdl/e5z+L
rySVl231RtbwMicWHD16AO7f4hyzgd0ez1tWchlzYL4UkjUoz1dwlSw9MPrzpm71
Y4o8Jn9nAwJ4ocJdYdY3TfU/DsaleRmWfehAec5X5snR8bfpQ83cbqfNJGWWRcQb
tpT4J0wNGHcSGbfAcGCfKRzuxGf3j4uRsac6OCdHiUQCoHgwo1xqr+a7mgsX+EkH
OchF52+2m/G3daWmDJ0qomhGV3SSQ3SFOSxWBZNSHb5iDMQM6HiyuvXbLlgW1sNR
gWuTR0OOSIAZObFaiL15xe1tDg3waYpUglHA6P594y6lCjWkASMMviPXMQDgXZKN
AU8q7AYJ9tHHsr1DjZcyLyn+AMvWX8fIsD16PioGZbT5/Z0anDeUNMmMrMlVNx8z
ZmFrxXmy8CLFC99iSaEmMaBAlp7coc7l437oYntgKRg0JeGfZrHdvpXVjbAgd065
IZ/sCtuPPdgr6WloBnVyjG5YwIS7qZyP/CrYG98FjGPq3RvZme6QbZeKeAtwJ7tp
5elBspJ+OCIUf9FKBwKkw39JLyOCeUQTtpSnCkdXiNRE6s3Mhk4rTie7RgmN4x05
nSlutqbxWC9rPMzhtCtyYQ/KrJLWgOLgTyNwPjfWZsHKgQU9UZQSOE0JThKIptmr
GplZezyGscAMsphS99PnmZrFHQpymygGADifJyYtAavI5En1sNPC2T8ILhNrSXCS
tRNNNCNwH0JIXPfnDpZgY9Mde4dBTQqIoYYhYh0xvq8G9FfBDeOFrarptRQhNFQQ
WJfIoEUdxcz6ZxEJ402eZ8OYpMBQUEiuM/AYfCbV1lri/onTp8AQ37woxuurCthS
6uttaivJovtAvH34yL9tcUsfXoKwiZ06CY7jRwc8jBVETVDzvZlXzOpL9tSo6Cli
fqWJicQAfdj/ghQMJIiLKbKA7tYpKeNSODl4D29Ncb3k1s2YUnD4Yuv51UhQ9EnH
b/sq+Z72D6c0eXfQiOh1JYsvoSGrXip2bRIe2SziYdWSUUqbpx1eDaW8hAAQJmk9
1pDmfHzUn4V2uGhCgpbegHnV09hF8SUCUksf/yG0Ohm9lqRaKpdpUFy8BHXYqAE8
pIkDUi2KciQPAV/iWscOto0d8Q9yZ9UuPrIOivmNuXDwqrs5r6Zz9boecWk7G/3e
0TGVXMOiluhOvcVeBOgOvcdUDXqIE0ZytRpBz1NYK1694VMfGVSHPH0Cu6jGO/fn
45k+/C67nj5p7KQT83naMv+yj5L7KM81aB3h9X9izRPW2WPoQ4+EEzITB3Etjrg4
DiudFch6nMXz3enjDDLkZwgvfUk3/mEVHf4TOzqvWM8UBMVJaRJ4jF7o7yF49cni
FM8HSUi//uuDeExCCbfcbi+SgBxT84o0fmSisKO+weHWnMtuA+e/SAkx3WzSu8nE
FhITrE9qBmYOZjnbIslhKash8te2UB/WphoWmig2zRT/bGXvQKlTRWUJZe9P+1Bs
c+gX0VEH/hnzLj+4QEi/QmdXkViZVSO21mbjEIJKEg6N6NgFvMUGZrNM8wtzkMGx
eqIgKSV2rT1jVZGVMddAU7YVLJuaFbQASjmApWKDFO3VccuyFAolWjZ7qQ1VS1xO
HnckLNraZzivd/h7hiX4ST7xa071e+2Jt3PBvJoChjnYZeID2ftGRCwagOxgA8s/
kfw/wvFLAQ2VQBJE8JDtt3EqTNvVOd0kBl4UjG2TJSyuybmTxG1LfNV8l5t1cnW+
upgKw73Ug0WbWise2TGUps6aHE7+tTLlNZTLpri3hn4IxtShrnUlP8C0d4Chkgs9
sIlnduxpoQZSpUWInC/iUHi/jYtVEu9p585GdbieBh6DU5XmLYj9MW/DPag+xsby
4HbEeu+6F61UiIboOJ/e5gZHm3CWUvlhQmbrY/lB8i2vaCqelkXYX+Ucl0PV/mlG
1bWuIMuzwafAyvdYp6bhLiNREbzHewqVBOey78Dnfy6W9QDqzZMnDCkqQGKyrAkU
Yw0xWj47tRwrY8vzRZLGxCIM2xVn6OOL6BXD4g9z/nXzyFWrq/kj3WfP9Jd9k9/w
700tfD6UqCVLebQ43SjrKPYQDCEXmC9JCgqYIoFDl6jEyBnKZ495JnVVCHZ6P0sv
HFbvM+MZ6t/RMRKBMJLeoHgw/PXDTuTkmIbzP76JmN0PCjJ4HJij3/Oz4mzi0MfN
rwIGP65OfVPBdBzxAKr+LntTzOv16uFIkXzS9/bCevv91iNSopHZfKnQzO2yJKD/
2ARxa3t/2p+X0PpPjnO0BFKtiyAIbjCsG1jGPk9ThrnCUfsIhn4s9TNLj72TCnAZ
1impdUsRPVHFhEkCWD5gvhi2b+d0kLOlDwCuKVCI4FzIuMxwcKpTwK1lGebwSGhd
ooyNxUnqhA4ybKIRtYF0OiGEFd1L0CwxyAmZpWFsQ/e/G+AyszPKkGvvc28TYA8s
bsoWrT+YPb+rgPjTJFBCPZVo/O9FLb8tA3vBV+3yrtriaqbdhSUlY6lF/06hYhyl
eNonbRtpIRUZc1sZwEF/Fidwu2VUnLOD6pjMmVt3cR+uMU9B6IN1hQNqbmd9bXQD
1KXqhD8Ni3TxAC979/t5qUTBlunhPf7i3hlew7v1HD34a09OJP50ItqrnU9FPOWY
yzrb25oX+NC8nksmsPhZ17XA7DvR1VZ5fZTSyeDHaJvtfFISQSd52MLixx96yrbE
28PP/H9pSPARSRlSPStIEOKkPlwAbLNnvynIMs3v4qzeTRRg6LPSpg/YUIOfnD4m
b+66/yi8TqyH9kc7SIjGMf+ggOlOgRSZk+MHyroJxNcah6VCJkuFdDLC1rqI3VCP
bzr33CM2X9mRnXiGAzA5qqxp0sC+zCoI3glU4iT+bVWnqfo+f2yzrJPEN6pFk9Ow
jtKwiOpAvstAKUW92yuEGLsQ1Mea650QcbRahJtcajGjf3iA380Roc5ELd8Uu/bg
8qt+XZ8LHdMXeUevKazgsUKE5vOqMcStbGT975QfD5t914TfVsZ4ocMVpFkygRKy
z8yNQr7HZUCaCW2J5yD92CFGTl+Lq3YzWvBATWIrCDYfDseeziW4gT9FUt8fUy9N
Sw7XfVIYnQXXYG9UoWVweuRmhv653OG6rx2PsRQWYQQVq2Ze0GS7X/9S5yIWwBjV
hIbH7NL92JHlnzwJKUgsbNYDNWpx+44ro5QVdozmVU9dbubRx2h8upsdzzDB2575
EzZ8OpU4cvtA9YronNiJZEI8LrglEnb1+caLaTyhmdYjFpg1ihvULifmcwV1CTjJ
EvgcB2rn3ZXqINtS4yBX/dxX1nf8dehIuKMUPSKNNIlnitwSRQl43BuGqvok4xuP
h4xX3TdUJ8gvuNQLJa2gOVzzOLjOiO0SMUS+L85GRAYjh/eqkD4i1jnjYF4n9yMj
DZ092lf/ukjNw1yN9eqllYmnRYdfg2l3HXNLx0vNgEqKhtxMBfMaZkSV1iJ6WPCF
t3EZBxJnB8GeKluCEHnS1oVWU5Lr0tyN9WH/d9IxZG2BJ9eIXozMH6L0TLNlP3CB
0eAXmiPMUIQ7iEy5z/ygzXfgFGzSGegAK7reS3IFRBnvWjiPGUsY9f/vStnCiwJT
urPIgeKj9GMvY4GgmUs2zPXDnIG/UCmZPYu+Rz0m+cGn9ZzZInWd+QXSHxDko0r4
v4hN88XIVLPXVh8JJMq6pRdMWHsNwql7zfZUKmG7VEWXl9ZvKDKRQ05mcGk4QDvp
ojl4E2Fus2CQv/QYvfagpIbFn2I7PhJ16QxRDnqEemNwTLzX+Ihx5SWX+qXGoa2m
AHWVv86SZ/67PG2j6i/OwHSBu01G5wmf/DAk9lvG8dQTSb19hApHSwoBr93pr24C
tb0HKk2N/mYwymz7aidTkNoCP9NPvCJGFrqo7Mu4kLhmtN0D5Bqf7ohleDndC734
jv+9guggCevRHO5+LRYwM+kotDHsQx14ca+HHJHK/jkguv6Lwj2u/ZzGx9sJY4GZ
mM8jXojjE6prua6hWsk3SCk/fKtSNc+oQEKfJDzVyVS71tPDUPJwXy4ximEW0kRI
Hjbz+O0dVrrVTLNRSLMkuwsRvnuj8N8v0kqKMpd/g3IIEVs2kSV+544MUZnbNvn7
4TzC1xEQ5Z4ZqGV7PHO7wB1mKz8gEi+pTK7QA2kfqO5qq4RNtlHKksrvKLSKGYXb
CfKv/Gbek0qL3lZJj1FV2AyxNOjvQf/DDNovePOK3SSQXtLLJQ8DviE8V1iSGf0/
dnlXanYooLv6OenEHfe9ay/sKqJSCXdeDZYU/qW17rdmLraH6Zds0cbl9en3EMVW
8CPUyuLigbcgDmM9QruaLgTw+f3loUFgicPDGQ2jiOTq5gKeDsCkap0pWxGCwJx5
MVrJDRR1I5Ye5Cv2wXuSXU611+oFnF9Z8vZ2xAuNrzywKvZVbuTReG2jCstYOsug
/pep3wDPoplKgR8h91qYBXf/ShnmsF/ZrMQRwYhW3J0zlTnd8LevGWfCHcXIAw1N
L3wuggeylrou+wGiMtWeRIxMnupk8LayDb9jlQZjIf2/aNy1UDaV3QhA8CTQyXfZ
eVLd6oHl3KPKDQqt0rERvvdjUBqTCa4XVTZlMguQT1X+/DnQKO6C790lYp4w5f6R
msa2/pmiF0RziJ9Jpa9Zlc9YpOnMpNciHRGgiP4ymbGAYPLobYxhlrEAcZpXPcLq
/0NrQqc7jRJyle/6gtx6i9NM02v/1H3mO0gqgHpksdS2VlzZ5TDo3qXeV8YZ5y4l
BBik7OrEAlDiH2dh/JxXWtg2O/i+IoPA71bFq7MW/+M26Pu0riW01GNtpR9YV23g
CwFn5TL3yAFLmD1jyCVGlEvIi6NDWfVvFseThmtQz4ISdKkrPLN+v6IGkKEgZaMl
T1rHL4I2IJ4CILvBJOaFq/URipQcuW8epbl5B67tpl/y0/KYfUjVpRnpHFmg5Zc2
EkfGANFSV5ZlR3OxZZGH48Ice74Ow2BZCa5yWBXniDkZBospjZyEMWDUEfOfnADC
LwqhKDapJQ+So2UvuQWF9s2aji7/T8xby1aT7quDuAHSOLclggf/MZLzrxnWjBrD
Rv5RKZnjP5RUTFWRIsX6/lMObVAeJIdxhAV9jbY8KeI/+UdVe5idmwnhxaujOKUV
DEKNYYCRX/93AsI5Rito2sVt8HhhpzzoNjdxNyZPq0AXcTxJS6r2EPiRi3LIuhYj
+84HF1B/J0FVD/HorrH/WL9hUDi1nmh9c76mJHJXFrC/5ASRImu28B0thVW7Tlol
2Cr4ZaYeiCGB2DMcHcbARWixEbX307UgHmcrpHXew5ms05MBJFAeZAkK0MrJURWn
XQV+Adq583p5d/Rv3lkLVOcv2bhsIpifMnE6oMRMxqPROdomo0koQug2rPrenSnD
SfArgiGkF8so3+M0m4wDiLvuu3JWnY/yfJ56SdN0xd4VjL+13Nw2nOkk6DWTQsxj
IUa2CzwPsmD5vZPDRtpcAVkQSMdSLbfnw28ihm3UXkBBs+pPLUAfA1i8ResORiuu
kxW5Xxk8S9LrPveqpb7TfUR2biDZ/EPlI8ShmY5ptNMplzFZxPKiNnzAlRsBN7rP
YVPAoOSMXWQiN5+D6WEe6S7Ssmj700uQJ+m5FHn/gUbI0zvgbu9ulOBXAKDzQQBH
GBkmrnkchZ8X06Q0PtRML/IU85z3DDC19VgdECuOjUThDNUOjwaCLBEk0bx+xJld
MahACKr+mxxeqYqtGqf0EFQsJBpIIsYuW1TdVVLx/veet8llEW+3p2nXg5uOq4+5
4HsY/BXkG/Yrl3IWgY8WG2hADC8hGO5XsL95LyDe8EIF7OtCKUN/aNY6hQgSoiL2
azB6u0qVMDXH5xVdORAK3nRz8UtcCIVqeZBawSJ0lJM4OfDEnfVD0bi4LNA7qyKk
fw1gmJ5457G29txvp2AZ9+49NKNaiQYx870lCHUzTrpqyTAlIwlNhUhcUr3GB1SP
o4d5ZDF1qiCCWYPiN0SbqetDonmlPaigqaUOaES0sfmI0fla2boIfL7dwABHADLG
lnlOFhxeo88Z7Vqw+mjH+ZuDNWLRZtlicOpGDXO2Qjp3bcW6M3bChMirYmdJzFyQ
7Hhqp2IbGTFonh9EFarctmKJa+objHezvg5usAiRMpQXw+8MkxIgM8iSKERMDrXA
jL3ztF8VEwxEDiLHcEMXdF780CzhO/mpvDpL3d8MzBIk5JnYq8hzlHzNy8Bxmwl8
ttIvIdaDwRVcJmr0iWG8lHmxNTbKn0iX6UG+P8IdAz+IoxbpnXWePB0FJ7IICGWN
hnET8t8swhm0wAVnoUdA/Zy6rV7i+Oy8/XW/dkpEHq3G9zxU6WFqzmuij/R+BfA4
uSqMrW0jA4OjhiV8WW6whBbjmOM3Q9CnBbeEC+DNMfQLvORKeEVtGs7/LlD2zUKg
gwSZ3aqS6gRCt3gvrjstDzPT75vbDK416xLW4W3rpIUSfCO9gVaVxXDIO8Oi2CFj
FfiT/SBAZclR5ESh6AEJeCL7Lv6190Lzurcno1VedJQoGFVw2quD2epUww73vm1H
ZZPpj6VknOtNMhR9SlU0yp6/lsJZ/kA1yKdt3VD08iYuoJxFv6yzb7SyBBTPQRr0
zr3Vn67fs/gHhCXaKGUUFuSerOhUFeJ+96nNL6rbQwS7WmdibzqxCg+QB4ilaPXi
TXPk1044rx2HQw3ajkCRnOdzacTzEAaI8n9+79yZMVS8LTQQDU+cb884uGPoJeGi
TzhTzEOa3GCjE6kva6B/jz1Bsmo+DaOyVkfYq+g9vipgkWecEd4uosjPaN75zgz0
CPQRLjobguzSq56hHe07obgv5XW6RwO1+Hguw1+uRqAe4mJESAzLfVaxjuNaFcXg
kcm0EigwawAZ4QiEB0U47KrgeRWq/kV/iAbcYfEq/LynCZSqJxXJs1AbricCnrmK
hOJ+st0P2S/pqgmM1k17Zc4yrRRWQRG2lm9mrEge8ucIymAXM1y7ycEBjmDL/ng6
O2+dylvdnfT+AbDulDpx5Dg/i03Z/nX4pzlQEPrmbUQBGAW02svQRw/FPHfPlr9N
mHW5UPx6HDRQ1/J2pguhsvT2kSvg9pIdTf8xkwc9iuO9aUQHZiZkaGGBA+35dl47
IJM+an9HykWmsyztqR/WSdGbPhOSLEN/79XZ8t0nHgUkb7QGNVqZr8uY1W+Cr/cv
yq5N2k7Du7hBOYkQ30obzJ0lFFkPWmjHxacehL4vQHIwY7JXL9KSLp14ZhGcpyv1
HU2FTaCkHnQVNYW0EPuRNYW4ZjYaEiuLmLclZzmmxy79Wzq4RrY8WpheYGegwqy/
aIy3/k0cbOlZIG956zZc7GOOV5f9figX0qG2hzDDaLItqmRJOs/aEmeGJStWBC2x
ROHpnp6yz7vRREKpagLkQwzrz8EMj6quKgl953xw/5HY+EEItbXhyv86xq4ntiKG
TLIjWpn5U82SCvKzKy1tDfH451mxM8IxcR0o9qmSJ9uzI4YhLW/tMOq+x5Anfn4w
Z7ssErADl2scAs0kIEgOE26WA5BFA5rLr1UtGmHZV98YjIOvyiTuR5VYKcxfBk6q
+ZFb8bYH9drapwDUHopSukbGxYm77yfqfbpqzolcYS6RY1yQFBAUYxIP1nWnP6US
OVasLCgQSumXa2HjGpJGV1fGESMreWJ7NJDpFgmDe2VsQS+GhdvckfSODWXqMdT+
kiV1EKHF4x+B1zV1ufrtsrgjDYigFJaG51Q8k9Dt3nHkqTqcWgX7vK+r05o5s7qX
d/FwGB/tUzZ3B2pDIPFyaFIocmPA1kx+hS8F5o0smjt6yNbJiJjPby6948hwb13H
A7BAqEhCY/RHFMoboyz9J35SZlfNkm+nV8/BjdbchYu8tWLuHPm3o+K3w38i3aPU
/cOdDBu+S2n5tIr8tlC36m2crF+AvSH33Gn9NqZfYT78Y3yraC7uwQB6wT1cC9gJ
cYoZWSNljghUn5S26+P3+AXVdbgtA5mKMbQeiaGBU3juur3Epq/AlxMNT5Ija6s2
c/otBGBlPE+3GgRaxpwgw8vcFvjqUmOzGWVTWZ5iRlMHLHL6yMTKdHOel8/SQyw0
6Moy7oexErMEeLbVWUkhPRxZDqnASnjCcEEKdg/joId/uu3jgb/Ioq9OePumC8ba
vifCjaz+Dwk/kkx79EcDwppomZkq+mkMebr0bbi4PN7cApn+zaAPB8++XmCrFZNr
162Yx6HHZJxz1RctzrbQT0+QWmqYdxrULGGT+cjNBAa1Rp9J02kUlSKRGjU0LLcw
xhSaQ+NDkvJSH/iNkuEaA5gx9kIGwQi2onwXiGv81uXp5CKNbxt7PRjSmBg0MMKM
lDpn1QemgzpNZ1BYUm12pORPz8pZo4MEv32D9cIBxdVVTv41cZZTFOghfsVv0rmC
l26m1RlwBglY6Ww/wVzIoS4kh2eoLflxR+1mrkUcbNWaW1HvciA68RyT+uLu2jXh
xhTs1FZdSfTGzRks1PC5bIaFiXmQseWb3R3nav0tMuc4bUCVrhzgkNz/72OnlqfX
Dith24HVsC7F83yofKjuD6ggNM2uevZES6AoUmm10PYMUn/oevSrdQrJxdwO6BVR
Pd1kg/ERv3Fw07HKQO3+gX1mkHW2tdwHepQiC+ha6ChSnIVag3brO0Rwur2iVYPg
6B9MpFRyRbjINjJIyr42xn3p5HYXlzi6/bxRjhx+Dc7tq7dYFYUSlOrlfOvWT+cb
FDgBPfv2rIKPVHlitnuvkd27ErmEIr/qdcRsf11t2bcZDfZoVhEU6NVQ0TUlnWn3
wNB47h78gRcE9szEWMHgCKTC3GkLSWYrxwnZown9rFOkRZ67iLcFciLBswgwMOcX
gw+oSgBL/piSzWN3LFj2A0EUaPrTW9ifV6eYKTaEkiucABk8lK97YqZAvvS4ZNhq
rY4ZdC7H9g3XmW0bC/RqFY3LzLkuADhTkLYMT5KAwMw5pNJkjfNna8s9+6KklnC5
alSrPZWB3ssElNqgObg30fLT73/YztcUMzXD4aTJEYJVQIX+p12xrg7fZXLycggt
A2MViX2MvSJp4p258J3BgOzgodPPdfgcKERT6uHP+9Hx8qWfSRS47rX/CFpmdmHW
NzPWHpm/ZiypnlAHk5pjNu8UkdAJZLUy62bQCfQ4cN5uA1SQ/kxBtAyADaPpC148
n8hWXA9pjB6d/NstidWAF2wxydgcbwnYTHfm6CACZStpFS/aQAZioI50AOOjz7Lk
IPARHxtm1W7Tr5qXd3COpaZEcXSk82dEM8Qm6qD01Xfriqxmqu7J7xCcQdVqRCti
lMf8W0FEJCRbKO15vJypiTkOKhKJd2wIuJFZrYe5wRMrwo8yCbB2cHOkwJU28FEN
pt6u7QvQG08AZQjWiAvaAytD6VicsKLGPulFM4dSJhy0AnfMgzR7OMaP5FJL4MtV
GvnvcBd/Qm/Uj0ULl51pQVg0YFaGJzhqHI/jN0lAIULP9alXiSaiDp/W/d26jmw6
gGkY9o/Md8raE2OQIKftx7tA7r2HruI6rn+cMuXiv2aPNMZX7IkXCLOSbGt+k9hG
XIM9zYuIWPSvwOUIkFin11GzhjF2vutNbUO4rY02FFGMVeM/9aCIJkSXuSbkSWpv
bQPJwiJF6lSAdj/3gKeFmHUptnsx5LmUj1EWF7j4F9PR/wZ7CZW5EWu2kA+JluAj
V607n9Mx3SB4OC4Rm5BPQSrsIR7uBp0DX2ab+Nmvsw6v5TMGTSgvUslFAZKIvd5Z
r3q7QTPqsCF9BOVhcCBTmVuhq6w3iqKxNfTDhOQEgwqJGgY6qhvfO2/XAh/vNxdt
B6uXW5zjQGHHBD9YlX2PAoM3seakM6BJmtWW7WLuIFZFcWgPjv1HYT8zSdMSwdT4
m0j0jSdySYiwcbIOj0vkSFT9bVLwlMcIdDradHF0EgtSR0JwDH658xj8W0hZjVit
mYaJbRcFUiGP1HzplZ6hMeaXXqjl2VwkSLCziyXIUdh/1+kMrCvABrC0PuqW4D8g
n5CEWVQblXgMZZhD59U2OFss5p+BA+TIEc0RMHMwY/eE6dX9OH8syzz1uyClHFo4
RV4k9cM407wAna/qZFh+JrEKRWwmmZB5EMc+aWCFf61d/MwPjdsQd2os0sKKINF9
ski0TnfP0gfAdzyOmXQdgAqCSgGEzT2vumxxJs7QjTk5nw2lhOriYK8JEq1FM22N
DBwtYd8r1D7upeX4RkSC0k2h4xPGOnWyyFYIZPkuLLnojmO+PjHEqdMNM5bxlgFk
L6cS+p9VpUVJ5YswkoVHrWX3uto1LCjWnlbSc7rlvPAAglcEJftGnoyvcYq2A3TY
qLCZ5w6JZxVcl+MbU8PbXUS0T9e9Lp+ogTPgZZXYpjaLJ+IuSDkLd3AgS2HVBsfR
e3Mp5NujW8+Gxh1CUczXu3MfH9rm3fgw6m65yUNRuPnGycpOUrHJL6ZvpR2KDCIq
18n66M8C/4pMnmjn9dvj/jeMkOteANIDkt64oQgf/zqZl+PCmaiENWKnF3gaRybk
7r2DBPvOsE47oxb3pOBg8iCpEmPtYPz1wCO09psbW2baDZ1+Fw0W4lKdHrHgdXIe
FWgDAQu7aaVGbMtRWc1tbQfBf2W0XoJxHJUXsYLT1kZyM2qgPX6cgEY6KWdPwmgY
vdE5AFli4fbG1kgHR5ZD6y97wVtxUW79PjgVdE51ypwU9mU1TckLTyJIMrGCEWBU
5w+ricW17IhbaMSTqwxyZQxdSVdkq7i16JGUE/svrbfYrrx62YCXlG+GYUuhuzcQ
HhnAOAdoKOSrodLkOPD5g20E3/UZ+usyAOfceG19CBNi8EVjl1xtGctqt3n/7ULT
ZTqyQdwyOzrjKnaEEBxVi66uBng5b+yHtvj0hdTk0qJ2hiHMGOf9Nb8pgfPjeOj1
Jj089Ve6Dw7t1CFjI24zZGjSxw+rVPV5KwOjo8hCrI5vk+OE4nmBnmv4u43rW/+o
fcXkW38ErTQWI7wefYmzdiFrSf+lLupCj4Izji4mVvo+tbbGU5n6G94QlPYRzn9g
8x1xyOBAw/KJM9fl2fEPARxoMsma/M5vCB6QTz3/obeVPx47p7fGCL1X0pXMCHnu
SuX26TaipV95oIgCItaT0eaMTLSSlbBGpkQRrUDEr+78IY/YQSfaPpzrmPvNX/14
8pMCaY72ffa+jxjjSPp9ooq22K8sjoKRCTqRA330MsEjgj6FoMIw9/XY2Ngwm9K7
AkzJfk8nRQovJ0HXaOpPiPQb6bVnpiuXFBLfw8y9tVC4pD64gVJHfaCEWBAY8P5I
/KyWR3u8tzmPhLQQhyoO6GGd1uwiWvKkIe4UColgUKm5W0MW1ZSOZYGman/j4Np6
Pz1X1DlE/Z/1KDhYpKolG2a3SxlqJMunfsFbcxKN0MdhCS6pP2njB++8VmMOO9jw
Prcf96rEcLdRWQnVOayTfmi8QU+bh71WxGiaYTtZUNEOQRhplEKvGUxFqdoGVpln
CRPAXeAR2Z3J23Ou4vvqZRV7NrZcZVK9sRul9gtGC1VY5zN/6YCyWkZsG4SC5g0G
OV+gGJKChbqH0oaSU9bc8gQA0JkiWIn9tYTlNjuQAcjiA9wwqQN5d5Ibq4MfuPfk
/OPS3mPGxkjto7avy8Z11fJiZMEzdXdoBaohGDb1lCYQRA3wIZo8sW7UF2+RrS5C
wKsuV7Ebg68dM/qxyGxvnus2qNl0w6auWq8+CiRKj+t1xRbyqKzHjTShivmQseBm
4udU3XU9ENbGyxF9lhIh87HQmb7LV3+E8MJnbCtLiLTZK2sAIk6zkCFLScUnR4u9
xZibT7l0xaK9zyEGTvTbEZmxVflvJGpl1XLh0ggG9CgON3VYrRaI1/ObFqi9upOQ
IU61MxJ8XBqSMJDoE9B9N/4iLymyKoufYrWLtXfAzfBGrrOUAsQ6JeKozEDvvtKs
io1rkBb12305XHwWqeAVt5CrWqZwKeSCGplEJwUcZ/dnxiqBimu0KsK6cz3CWsak
22SfHoldFdK90zVAPq5gGoj2a0oOcGwTSHSI1yNgZF6WfxyTCDE3oRhlQB6b2bsg
yxt7UL8pqq3FzqiWiz89nFS9drwxQZH4jw3W+xrQ2q0bZ6v9lJUYpNLZ8Q/dKfKZ
DXeV0zse4N8+VD80kJ0joCtd/Jg7yckubJ+78vZwMg4/OgLcNvsYc/qrRMv1XkTn
gYt5XX3uKdj0A9TBJaLijC816Xg8gWVMK1QlFCYcLLprZbL0Uk8lSEleaxVmkS9i
ueiGD5AJkG8cbiJeu4LgQvn2iVU+cZeBohXGJ3OIHBgTVpSXMd8/30bZca2K7VPO
vl889L4RUAJGI2eglxrFlBv9P4lltMDXW+UX950QnQxB7pNDqHxX9GBOuRNW/qpH
DsTuMiKzChRZyM2EkWjLGbqWnA1+RqlLU+bb/+xLfXaD+O8Nqg4AD5q69nyfZSrX
iDxWdgmzAxsBmoP1CwAmE796npLOqQOEZZmGKCjJQv0/Z1uSEFynj8iThlZwlbE+
xVE9QBGHzvwiiS6IzYifYhnc0p04l72PoC9Itj5eSrvAzNdlHI3wt+pAy+ZPEbul
cc5Ko/eerpwUsT+JV7AJvtN6hio8N9vdJKmb62wT//y8OYnguQRsOqWOJowRF9te
HbelyK1JEQatwGJLWRchM8pMDha+fXDPlWOoBH7FQHjXYUo4plvTqbiPLrnYVsJ5
6oNyRiwIZsXE533Ej8uSgPEgjKTACyMQ9BxDlszKJlPwEIN8y5pWiQrhiB2anwwG
IfVU0qFqflZrGBwfRWfXiB55tBhOG6VD7wA25Fm8xkisA/JRdH7a3SLjSctsgX73
+9b9dozmOug7nTiLc2jfis1Ta2ugsYlnIyw+zNBpYAwH7nVtuKPhiUy9bzlW0Nd4
3hKGZOrBOdoS8muOm78xL5wTx77/vI5uSSwiOOSJJFxcsfM/Cy8qzyie6GuTdA5R
+uReH06fK2547dVth4WcSZjlX8dHfB3VPTpsv4U6w6daREtCbmPCbuwKIcP0VzGe
TQq11p2bJYb/BOtDdfLLpRhfOtPeNKrySV3uD69fBZmY8y6t8cWr8BATLaBh1V47
ptsN8MYLxIozdsFCwGu58xPKe+0os1wrrkm9NAS5BsFVjLX0R5B/KNOC13eeU2Xc
ZmkOBLnN4Xr1/ZpOJNLRl6AjC+ucCN2OnnUl37UouSoMXyxJbxH3BWZBRBdVHhEn
/wFsVlLJgC9kizDwD2+I9dscATZSV3DNWdA/Na6SheB1aZLUUG9GOTt4wQcK2VEt
mv+Q0KjVMmZyMz5hxu/X++7pykggf0mVp94jOP1sclg/cjK1pJTj0FPd3ijJAGY2
+B+8errnLgWatPKs+2E9HZu9uy4D+zCuFCwEDnmhsEY6BOt9Ge3TPAx/KbisfcsJ
nubdL2Xr2/Y7lsxnBXVtQ4ypZo33kG9tsI9ZOr5G/ee+xD/OveoPZBlsieClNVfR
zP4MQfSaCS/IW9NXOtU5HJISA17zid+ClTuM2typoZzTe8xNS9Hrqk9TCS472NTU
fFuapCQCu3CUeMWpuTfq5D0/5+mRepSc5n8dZ1qYdWlwnKpBDxhJiwVb99hgX4PS
g7NcDlRv9waRautI/luzrpI1FcE3nxFJQZYukgwp/ounIybaMDuVxivNnpMKNSYx
oqfdmtSNLCo5xWcCFCjFgtpWYqnhm/WSJSzxdLsW2QJsQyd4NrIYUtTMQMMhwq6s
vvy2EhF3lF7h1LIevAqzrYFwLP2qQDvDXs0pbOQzIH8k6IT4yefifL4fP06ZDq2V
1h+titj2aVFKI3LGJcr9SrNmL1svOsBAssCyojyuWRFOnZHVSVlXe8nplc3uVtP+
4DF/yIaqAdgaLcDHFNe7vXbCu8dxs42RJTZscKaPy+IUUex/B+uQfSXEAoPf/n7A
wOK93eSb88Zp6E1uh7e5k2rnUTZRz7LjW9EnTPGr+ekETSWTaz+owYpQA8K/Fx8B
AqXFd8e/CYHUwxb2PZVinlN6rFVA4V6wNRC5Xz6W6q98sC9ms61urNQ3sIKM26o2
wyKvE2H6MZgvQPOXEDwEqolzATMPKATgq9zPuip1Ci97mjZKYpjKx+VuwikCoBgD
Awq+4dRACJUGivD4zHcpc+soEeiKMbT9o+Oy/a4jgkTKoTUneoRJRN/zOm0+erjS
dRgcxnM8Qp/ttEjfgn76V65PUd+ixmI/CDY4V+znY/Fot1JlP0hccGOo7yxYyDTB
AKks75tHqLgT5Pcj7CCY7G2nKUYmmcLXE8lLADInmGaZeuHAoDXq/ZbUCKnCrjV7
QprA/Da+bMs0jse7wSzYoUfbBqhfqnyD6uIarUL4cxWPLLmGBnW6530R1Rp8JIaY
tUThaR7tUHjLuWP0CN/MLIsdJGbrNbtd8Mr+i2tJjfz8/Nsvd9e2IEkTt7rCm0pz
YLIWvfdroOrAH8yAfhSDQp9BX6qnCxDhl2at/WL5sdyWJAl+CV8hSflT30eKVxPY
+uR8lhlj7vIQEigOHbaOmxkGo/trvqx2YLOvhnh8RJx9mc14Kc921nvQW5PvLjmA
w1tuDiBBtuM8uoGACkd4Bkv/Hebp+f++7B6yiNtwjBCNLX5aFyQkGKjMO4LlkcOM
wmHWke9VS2433oDergth+3ckev07eN7wzbwVp2leXmUNc+DovlNCTka7cjvomt/T
+JDj5hsXmJ869hQIqDtsUcb9decWhw+sM3ALF40rZONYUPWAMiK3xXXto5JQxCVu
5bnNKkcjPQvnz7D6ZhRpb9RkXH8INVOgF1ZSdZGbA2QZ3MVUgC8lGoRRxCqdda2G
BHlbUUtv9jm/aVsteqqlGiQaLU2nYG3Rzw/xpoVjzQMW6o6W5SX+tITPCd+2KDPP
DOI1djUfrqeDqUEP3gEDYUepzr6vIrtqZE1dS8OnB05QYXrm99k9iitSHRx9WAfm
+g0v+8k0tk1w4bBByDzRmTxoPzLxiMCGOZ0kgopF1ndtQm+f3Uk+aqLQk6o/V5yR
SGE8w5hh7KVnqN6BfgJ2NHBJQsCu0r9DHiAn0y7QLj8igYfWTWqmBm5ZcuKA5j1d
gukpJ5P5c6hga3f0uRd5uWe1R4gM8oZMrD/ptkqkWJyO3XWo6S0H1Cwg5IIMcZUe
rufs1KVIUpca9zDi42ZVSv2XRHg9YukCKdHSMOaKb05kP1bwi2pChKKHmTtVQ3DQ
YWTwFZKJyrmcDsIUKTkXawUD+TygvlQP3eJAy8Lb/pPmXvmkZTmWi3k4OZNDbmdE
8ymnNEpMYH89mk44S+/bXUoZVk2ZmK9ULFce0s9zlznzoY4N7Ckslafu3Wppy8SW
nC0L7hDiWuuZAWGraweH1WmunZR6Xdt64i3XIujTpN9YobTca/uZRnO52R+eKkcZ
EBztNsxwZLedUjOBCtwspvfQJt5hLzYGoB/6uGrzc+pp9DfzbQh0QokA5qLCHR5r
vEhNbpZodd5ldaTb8i583OggroRF3ebXzNqUg0dD+f4lSZwbQOwCZlw62IPDd0S+
Z8XkRb14+uXgEkk5RDgWopM/BqT0HBuhCDqArSwu7xP0TuBSTJ+T6+JYlcvTUI+x
TuUhNOVqHwv0vLIwJ8ry91+K0qKJfY6qmIzdA+xQvRzL0TyNHh5YL/B17PCsL9wC
DZCTJdDFUYmB8qDZksurHZyQmRfqrtUTIdvcJ/ivizWWVY7sl3JUiZOcvKIog3kS
ZYXQQX/u0nXDq050Q/zAQxbV25Mcn7xIlTl279n+Cac82h9YAI1xba0OUf7OB+K2
ydP5htHqUyl2CuiUoPoHYYVhWIpHDWx0oKhZyAmWizIs2ttlaoa13F3zcPlvAaed
9paSI+A8Akxac+X6JCeKnyjyn3857pDJ6Pr+syNjAveE95kvlOl/wkix75KLSKjx
uZJDde7vSCFMaGrWUrCV2XVbRYshK/f/0S3kNgwu5GOHivMAk14n82W4aLr7zANW
LjWyP2jqtkqnAOzP+aEyd7v04CqeXpeiGU5ptGsZuz+BWruj5gYBIh0BaDFJRjKG
BkqW0E1jt87B++kducbZZS3XN8j9VEZPiukFzG3Sj5kajL1xFVqnzf1SBIL8popj
v3qJT9rpxv+0A8C0uS29qtR633r1YqH6of0qeztjJDZAMvvs+sOMLcUw/JAX5tBF
3qu/NDweEUI3Sz4TaJ4mbL4QS8805s1lYrJc64/5PuvXVn0NpAE2qKSJIsBZC2hF
A9DnBp8lqtR82/Q/xpvFtQnsTK7G2GZIOt8osMpziqq7AUy7xbD5/sQWw2JD3xTv
v6X0RLfD0rr8j/cO016ROXWfdn4SqAcsfv3n5WJNkkglKljzkQcEzyCdupKy7u7E
B0xaTRXiSLxa0oU6U3sw6EwZfJqS7KNBZCfG2hD7Uy3X1xSTtDzh4bKZ/Zq+tdQf
NipxY3qZcgGZm+7VSpA7ZlWvMi1M6XErMrnNvf194poW/53ePGJg0UtqiWaNdiwg
pEu3s4KV6MtMumF4wSPnqXmcMEWUnjEvmHzf9G8m5sG2AELlSn9wBcLxbPPmmo0H
1VB29Hh29BNm8B0TZCtYP1vA0jsPlunRyX9wWaGs823PLbXnaSkSNTld4glCqkTg
EJos4iN+Lza6PJ3s3+jBiPoRX84rjxHFadWTWD+QKcv5DCqnvBknTDAhJoY2NN8H
mVN+DhLxmSNPBOhoj0glyIogkKxD0tbV/oCHJ2d0IZRVFIxRGX7F/8w6EvaNKLHw
KZf61ZB7LZun9kavlnurEJrm3LnnXrBe/9f23zO0DPpIGgaodEDEgpebWzL7FyWq
SfQvmTNx89padZw5Du4RZdFpzsE20rsGBfCSzG0DCQJmIiYZ6iN7oN4N0v1R2izd
rXC+fIhKxY2NegNIQaxckOGZln+h5XW1FHAfvDg2HAiRSxdEZ6y+Gnfj0cZubdQP
kQvEwXr60Wg6DcjCNr15rL/rd8DHnoRb22x/erD2AJi1C6xHkvPeJoDh3tJNu5nq
wJyWZEAyPM85Mo4wEmajtMk3QOOljhKGvYTm4jzUOLjSevWqJajYD8/IEXZXfUq9
l5GxlR1hQ+2wohb8NPVOFiNl7+VIJs9m5m6gjws35cn5VwWRxZWBDp5sPgzX6c72
bmKkJ3BPFtiuxcMY2q6BIhc3p80t0aY0d1RoUCkU1CJygL1JhpHxkXVtJ+xS0lG9
BLalJolm2IPsorZXomxdZvP1ZIosjcLKpmsVwmqb4HgIhZ3fzqpJPEl6qn1L3UWv
zCYCmFbJjJeqrwK1Qr7yb8y5hgY49jWcdyBzYGzZe6Y/k9iOQ0+5ccqMRYaQrAem
z3MWhAHe8IHdhz3MfgLiI7EhzUEqQdL1bFPgN3AjzNPNQJL1LV5BKIfTGvDxRzxO
P2hjQEOBnVey4ynMDCjVl5bmPPBVN9bWvsVuESR5RyE75fP4d9qUlwtjCGFwhCay
XZ8voCzjIfCmz4Kq8t5o7OAbpT/OG3p8OV2OSVKwqKuGcqssw5iwjq43FBQ1hNaP
uqMULx0HBqYXdW45FGI/qgbxZuQedIi1bndz5rpotOJPRXBDvqys+hUJH+2hGzaf
AFL5RCCxDTDmtN27OEcDvhxWrDtujtWv5fY0Se8TToDBkZaTCkRqQZTxefyMKQ+7
Dbn8NfhrcITKZwU8HqcT/Uku7xZnfX0LKHmJ3sREJ2tsORlUmB2SkedneNFyZUyw
omAAXqjnO+H3LzwxD+UyCaT9E3X3bo1FB7w5GLb5yzgH7rLIpPr6See2V0AogXir
dwZeArIESrRnzE2ly6u2kVZeexO+y/0T8Kn26Khu902hegyIAlzKZaVRnnNAAaY6
h0M3P5FFLNCorJ07hwdEUt+CWIhHcMc/mJd1wLAKrh5gLILTfvjMKXBtVg6XTWEb
qsD9x6ZOlzAHNgQJw7BEYdlx2MYKFLh4Ajhs0V7Hv1dxBiNrbqA8WDmjVdxlGPdX
WVqjqVaJdhxbyRPLeMAoIJ5oT2CtRDD7d9mvgzpi1J1suXr9tzmIE6PbunR+nitt
zbUu1vuB7b4uWhBIaktzKSeBPuJPUCdPjuZAa8yIU3KqPmmYoQT67bYBV6ninSfZ
8LS1bppd+ogNpcNoghMpUfRXTzdTtRbZc+L3jS+OQsZ7SaAF/DnL8fTi4/Q6ndnn
KwUNq4n+5lYS0ZxvTMaOiASNUQqGTSKWRFA3/LyaxkT337mIRIeHa0Fk3W0ueGhp
RmYx+haX390BlKAA/hlrXbSA3hFywaGIrTXZaifREQO0c6VIDNUONGEj8dzXCOv+
TTIFqkqRWzGLZ4aIBTZnOpG8GDtZpSrSMSrq3nhTTzRC5vbTQkSIRkV1FjaerTbW
IGXzeJ/pz+6aqa4C2xV9xbVI7kpGoXG2u7GB5Zj7A8fUNHGlOz0StReUbaHXOdYv
LTwofC3eAJI9a3uRh2FLGIveQiI9j2PVeDaplTECt4TGTkxuDg56Vr2Rx3wcdI1i
6eYHFRzHEY/i19n94lnzkRO1E5Oq11tBLmyNp+FT7mVi3L/SWDHixYdolc5qSZSX
XucDnb4/9Ya2qNyGssYCK+Fd2U0zbXCy9zBbrqeegs6HwHSv8XnJ1P7LQHHkQ5Tb
hXTIt2SCSfa/f9b1pzDyiXQDdxdTFr4VHh7HDQybFAgFh+o807spggV+dkTztYlU
lo0eAt2oDJ7hFuacASQ2MNTl+UdU7OskGVUpP2go/DH5gB4IH1EcjgcKKh2K5+1P
y6hgFgfhY1dI5XT7+PXFdajyima33p7BBvJtQUej2/ImcfnKUDFVADHvTKjsVQJf
pEd7x2YBDqy6SheVtvMK9F/H4modqPyqQGZkaH3Ujgjfa+7mx3TAn+R+mn8U3yuQ
JyfLxBtEkGQC+9VfitEGSCBZBS+iz+dgT9LM+eOKDegkhDHy+bk3gZHPqepEJwGi
CugDhlHDLy1hgv4BWobjuA3Q9hkdAXGTx/mk5PzmYmnwU/+hhQ5uRZhdtYlNel80
nnKpnDIKOJuabTpF8euThMnEcyPzsW3n9YvmFmk6LIssCiHNWh5rO2YlZcnlHQ7L
MYkZua1LiQozqSvUOFbH1wRH/+T2iCyguv4TfKQY5BYttX2oLRCRSERUooBXOJzf
eUoGFHgvL3eVU5zNAe5UpUTrQ7jU0sxyGT28xCiiSkj/x9yQMCIONi0LOKMbjDPG
HUsFa2jELXjjtwcM7xZ4ehV1CVta3XYL4z0AdI+RT5DxOieBb5sJakEubTV26UEu
UBMldIlReXq/8MMTMFHNPpv70TvwmmjGy2ekvXCZ2VUieSeRHiqw9BO6aqyf2UrB
r596/TqSghIB+/Ae2jJIFCh6j2CPiRisA3DeJZLEAmsNu0EHBx/B0hYiiRuBNhxP
F7617rMR/gxd2D2b3HESmttq1yN9gKgr1jGdlY7bzGFHwwlw+ed7VET9Ie7Qt/4G
Z9bHiPfEghmmXeSb83e1TYBw9BYHcoeEm0ZBy4hq7eWvaB7p5PyKgWeznnA/C1L5
7+49+jDGN1hDSFe5LE3Ms631si5xPVIgzA5Q+ZYyQb0ICUu2BxZnTwKEsX+JAdZN
mnck156+xqoyovB9DmlnTaEY/YugWDoFRGJNRH2rGeUWaFFoKfao/pgzR/vv4xvM
uwZjIG8N+NWRmDedhWqUcA28TonECA4gRSTy5VlrLVcbtSdlfZ4wkil5OLPik2hJ
87XINDl+dXfYFfH633E1ZykOEDqyKTmZVB6ucBx1TnNQl7dmG9y9dTQbhr5dYkaC
SUDBPzsxp5T583Vhdz4vYvo++kzdHITpxZySZhUFmF2DnTNikYgsKPx/n9a8iUBF
vjj0w61zS3DaofA1x48J3PVKe0booHE0VVPGg01hscomTB1oR3uawZVr5SXtpwrW
biFeBFCA7HygDYt74CmUnaaEBMiRSrNaI7vWmtKnhvJM/DzuDvqbDG5lm2VK05+C
aW5ptkE/usYR+L/0EKwQQI9FuUc+MjfOuC4DloWv+8ZdxxISbQC/+S/dxlKN8zmc
wXWMJpiTgIwd7kN1JC74nk+nhAA8COVScKsEbL8f5aq4OLqFJVy8kJJc1gP14VfP
jyMR//JXBvYSAl1ulO2CY9+fRrnw1hU207wiYwvaq0Pg2BtjrAcuakn/q2yMmVMs
fKSHJN0G//FARhgxNazENKfuqcOKj6zFNcLcJB4nI+uFUhxQn+lniHpo2oJhWn6l
garG1DHXfEJ6uMqlR/xIr+FFwWSj1H1sleKS9ZXl1mf9dGLEWJ7IGjif1ezvcTGi
R5B4P8KrL3i1hEsqG/tjvf7xTfEHkA20oweTN+ypIQulhFC6Q9zyPcGrn5myhm1U
ws1GVW8i+GDUv5u77I8rzhBYC7HHnsIKM6ydIObNxvY45iV7NyiHuDUVmS9G4/i8
yV1owb8DCAFgn5ExS8mHCCCtNhsXgZTo61HCQ++04KE1234RJRBd1ATxfJVs4jR4
jP29/wQY7MlAxqYbiiwtfUpdSNzVFq18ZMfGqbteFykKRbNDxBc3eP48+2lDHgu3
ZX+D7D4r8xzwYmX273Bm8/i7L9NOrh4AVWsYe8OI2aTTGz3o1o9FQlmrDaqwj1N5
uWGIsOmZautSZEyAarseHIojSLNFAa9X7ngc/b6Mav9wye/z1V6RSLDUyplkMwDV
bagdxm2BCSkO0t1SsZEsC3fmhwDAcLHLDR2knO2BLz2lY5O6Cxf7ediGIeghPkzP
YpDH6PnptyztvkbYqxrOBVYR/3vaSuZVp58gKYBtTlf4AwLUShQwqAN9mtYZvVvD
VtDRGINUPCOmjOc40L+nPDxqkiTEMSjsSZYPiWOPxcWPXX9Uu+Sh5ofk9JcCKca/
UCAKZ8TsG8WaogzskWwWaN7XAcozO+BUSV1Qxy/NyrYWyDKFtQF9gP7UOerLvOt0
27i8yY/uf1SlcNHURAnlrr8yA5DrfYYrMB/q8qAEpf9J6KmC1KqEgdCIebPmHVDX
9FhF3Kty5Sh8dRhMEhE4uRLOUe2jqljfq0AaAR2bU+qLqBEuPsYtCyOfsJ3izWjI
juVDvfr7kYvtJ+E+7+BGKUNzsXA4XksAd0O+08Wwpm0ui8CrrYx/WAUNX5HszvP1
5Ph1UKsuNCBo44MKLd74wFLC+PPnyu47oZDphm1MklnyxSkHJGn12yJ62MNC6UUw
MqELHvfiSHSK1+l5IgMtnR/G/IB0oXhlcmrwUHCqQREws3sO/QuJaCaJUIDBP4zL
Wef8ifF8Tpw9kUv+xAx8trqZuCxp/4NGTb9h/MIaeJ2wGlCq/+jLPJAGoONVRW4x
Ta93GQAbRbsn6C/Vyjtlo4nsK/+CgldE0IO0Hd3rOaf8Sc6vteqnzWjjQZuaUqQI
c6tp5zMk2OV+/74mbfIujvoN4NNHPnllALFzADP5rRxzs1f7sq6wO59Hcl9g5TZV
Nf6ldm1vmPkLvmIxPha8dmFxISQjjlzIqZRIQSCsS6MfjChpoaj8vbs8v+xMPSfj
CnuPpMzdMwXaFNaOiA7D6Cgl1/ztISgcBTycBtp1v9jRcji908MZzUgh3N+3Ixq6
8d5nfazfG9uzCDlD/q2FbAdZtDN7nEmxaTDrD4Qw0OQKbje1WA/rq8J3N9crUI9i
l66nl/ztnam9cNRMKNE7ZxZ62FaA5yxXjb1g0em38GaJdGsT2oe0doBneACuE7F0
dApRZZieQyPLX4tbQUYdfajDL/QESAMFVoz7NQHkEMxDT2jXdFojzp5HZlZ0ukOQ
4fkMziHEV4oS/VfOlfc0SBwYPujl+1HoFVMAMeNeCKZHiGoXCy2IaNsFq2jSrFh3
7w1jBddq98u73BoIFNitON13NOBbBvFSW9WDE++ZY/Masq3aCBCFYZpjA+eyXd95
o5TrtxYZHdSFj4cbzX6uoAQN4m4HIwvdaMVAYG6nSxdd4pQ3oVOyP7wLk9IyjYax
HBFB3R8LYh0PSqih9T3caVb5uEabm+eYhnlNB634j3y7nYzF66GJnR1UXkI8hFC/
Gcto4BugiU19IiwKeRo823l/tGtBU5frnv6IzyrpkjaaU9V/0TbigJt+lZe396/t
r6ATXxD83EJv47a4z4hsO5GQHzvbQ+Gapu5GG7tZ6FXHCou7MBYKipVgU1rMDS2L
rc8sBnhuKVqZ+oDQo8w8S8/oGGwNO5h/ZxF8jQ4D7t9Q7zRNK2+5tepXQQzWZ0kF
DGeENaIL5jaOlEH8Mn1HwUrUPuXLaySV4m79No5aREQmIqUG55Kub2LP+qviiSUM
kC0m318sV867Xvrt7PCCD04IRgTU9mgnV/G7fXlKRs0wLbVGjqCiZ6Dd9Jri5YF5
4Lq6uvbEoOt83WYZfwheGo3tyY2xtBNBA/iQ5x8fE3iuxG7Yn/IyCLBnN29oResL
iH574thicLdAdYNU3jUN/Z67u+doJOtngYkpEM5Et09ojkFpHlfNt5jZI+stflKk
KeMEONZdE52cP57iTZjA4N0gsS5D0JJJjCsagoIYP02DOGwRqmIiHdxW3pKL/S6H
gNYk0R0TEfn2AKe3X6REgQ6bg651DmQz4t6vimciC73JlF+86BY2NIVNwnMxYWE2
GkBLSGWcRbhxgRnGL3+a/8cvCTy0ZZbT3FtSFivu8DtE9zllAMexG0R6AoQiZKGh
21iPLymCsnV0jZlZuwgCCONau/aLhGxGOvGKRuOPknq9Of8Rco8bSz04cHwJOsj2
O7rYkBT9ogeqUzfZeBWOdsI1nlDSstZMdTf0EYBUR5rhv7x1GRqr00Au2wxLcWVq
LouaWghuOTSxwy2P6Lh7hlAGFpLMRRc/V7CDAQVo2ZJsINq/H1CdajnJXa4KkR44
SHTkGYu+EQ19JkbaIga1wu75Ty5GKhthWrBab2/vLVxYC4C0nCD1qqBkHCeTtigS
ZZTJ+pwShSAMLjKALBDxV0kcYQr7hObk4/W9MPqXqibvXwM1BuMnzL38KUX8Mpj9
BjVRgDIH5ljBRSX/kv8u7GV4PPr7TcNd9aSV2nQwN3q8bJ51RHqJreASpMEJPmAA
pHQl6y1IntooCUdkulmpqsG8yniKQ8gKzZ+cMX6z34vMEAzer5bANxkCoxW1OLww
qF3h8d+Dn8ltFxc9r9fS14GHRGFKj9qVaiZLYKZmHuBRjp4Cy03l1FnVfnxTJSPg
yyDLkoSxML/EtJ9dH1DsmlwICOlp74g7HvcrvOZ/PCShA7eQSNmqDfSROkTb+XnX
3GfXGOoWTRV1JErpA1vZ5gkjqNmY4lxP4/XNDa0Y2tjnvUXapbLWKlN7bHG93UtT
Ha718xEqLgGGAvAQclb4Bduvq0VhD01+OFv5N9M8QJex7Y1Ym/HtaGpNeC8sMdfh
F97+Y9wvh5CCSBRtIQXyPmMTWFs3l1bk4DTl8Cm+irTO9oH3IWkWuFHDepcETKFh
fj2Z4o/NCV4AGy0ddk27fq4LHVbV13ZQ7xymfWDLiwOuVGqbntpiq/WrLcGFvNdR
X7W2ktXq8h1mekx0lFr6JfMR2e8LhKXnckGRthB3sI6MaGA8CrnvTtE2gCpp4Xd9
u4eaAH0vxEIjcDZD8/Up/7eow0e1KlNOv7N/aPUvFEotfHxa5UfWAQOuRA+BNKBG
fTruS+UBp4TV2FZtRQ5gbbnY4DNwch1v3IRgit7luFIAjwq8fIhlNeoIS2y4tTA4
XmjYS5gT84u2dOACZ2pWJVd6Kfa4e9/rKK1vhmjD1pS2mQntnoT4f6RqgnupPS86
xrOhrz2/zyImVU6wFG6Gd5pdZbqzs0j5ebpywHo0Bol29gViw8dd/BX1nbTQBfl0
E36gAx7tDi/R4waa1VyDB6BUd45lwbCToGTiqGPzRnw7uzBJS70AG3naLIA+ybEU
NJphfaOhAIfnHOeQ7ojdOUN2tIHrf5+rZY8XfCVmPnuK9iZcDXwUbQfFIs/GD9Pw
4KB0TK6kuHby37AcTtS0VkU8eyvlwVAJVuvw5rUFmrX+oMS3VHubdoH52D6gqVH8
EwqKnE6Mre5u+9WDtumRHBRa3Sf3JR4IblxEeetpcwaMxi246FJanbMrxY5RViFr
sbLFAg60eprkajgSxC0fwH1xCD5oqRxaS9aQqiiezTXChLdAQRqqRpiqMxPSGGUb
aVEIR3BatS7NCOmbfvZ/Iy7cM5P9R9ggqe8QiK70tofel4KqUxREpsF/TJdBgWuV
3UfsIbz+yx2RavoIWHfdTToW2FMbuh5YUeZRTMav7RKrYsfgpe0d4HpgD+lQBsRG
H+vKGq37CD7jzP+pdrLq/0TFyA4oG9JqNSLr4xD58zMTzROFhS+mLamlRgnfJ1MQ
5lUcefrvsVWvK1L2GHdNBpoyaGuRtn8L+eyGHuEg7YRMaEDmNdP9rmRRme7U6wXg
L28j+KhtAQC+UrfTYg5CLQeunic5cI6DxsFglhQOcDOEeXccWENfsZojd+89y+2Y
0NvEmeOe/OLBtJn2mzqiwj5Sa/vICN6cqvs5dzG1Sp6Ld8twD872OQsZb/qRUAB6
xgajyjcAuN8HsB7kJhAyYJM6n//T/9X3Vy83Y0krQWrJSoF7r9M0GOqwKTdGSzE3
iOi818ZBcYovVrUNtV4ZdkQ4YgShKmZGZROiBniFg43r2+7hXRUQLu/tOmTWigM0
GTQnmjYzfbanuZ1J4PwNBIPLNJJnLFQG3x8qjHAlw0TqGX1UtcQmkz8Ma5P9goxD
NP9iChxY5N5PrejWMztgC+MsvAqdV0ee263wyp8R/m5uCyipu5r7a+BjQOGyMmk/
ZC59KUGPOXS39no18NCE4Xl7fnUqW90Srwkbi37UkMX00GnjuPiahKUMS8VnElY1
0D+0CHXm2ORC/PNfrIZFlsSIIK2N5uCAsCT604OTg46SdP4A4OKwEasXVD/1apjV
cG0KWko2I0A4gwQIrdttmd4G+pvIRqMMHKZQ4kFEl+YlCgJzcrUoaYf2xANToSBO
mzLzP9OJHcbtXt4bMHe77v6gXogD1ajJpfi3FkKKeoEh4xDa7edSu1dkPANbMX0z
PEv9F3FM4A/9Uu3DuXV9HEfFve3CCXiikKzAg73ZQU6H3DWt4dkkjmbcaiYz6cIb
0kZ5g3L+Kot7O4/20UIAItenAhoFmJk3z4i20I3NQ6KuW2l5fJZPTcZTpYZNq3XI
1Cn/mGucDNZrRUFh0789KDNrpniWxop0Svp3sEhWnYt7VbaKnVdhQzjNNwZ1XkZd
y5pNzlc8knjgKou5Swk8WsPbljRxhdiVm0BXOLn4j4fe/Hjt/sLCfVjrUCPeYIRs
X3M6PYaERvnlzdf1R9q8JmPQWMRh192sKeXmePbacCgSxxr2haOpkxlJMkSez3IA
bbG4kKxt00A4+NeXWJTRbVfKaOBy2v60TpYBtr2NI3rI2Ppt5deytjdtC4leOr1G
9mZarLSmgmx3hKtRSEYvhoX0Afq8t4v9dYGXih+8rYr28Yy3xK2aDrpXgiSGdosn
cXGoSVXebMQ1i606bZIryEtx0qqj4Aq50KqKOk7gNvc6n1fui85w/1MYn6CMBqoA
/9IsnKQjdZ1Jti/O1Hzy/TUIv9wxkR+CqHwWppOuwF/720ooJR/dKu/GBcJzjw+d
E7/jq6l0ZH7M3riNOVCnWpyZlORF343LNInbflaA8XRp6QlVvZOEoe+TWUdQ9Lj0
IOUl/oFgnu/1N8meipCuSkmccqi4qz3GXrdOw5xXBt2g3kybCC9yelU7gL/B+MhC
mrtzxIWPPAx3rMZxTzZVd+MaEoVnJhQJ/x1Op3ElFlyTho354TIuUGcLMq5/3eg7
vMPTapPTRkTeTBCkxN2926yERnpjKJPFOCVkkAV2aQ69mIVV3SEjsN0Gchw6UxBb
g8SY0WdzZm8tVGL+qL4C49uHKCFfRRhRWN87nNW9L6kEd5Vf5ZVBgh3/AEOhjN86
NpjAhqTxI4v6njP+NtczhCq8qrgd27cpjucXsXSzs7db9ObKrA9pdQbWlnuArM8p
XMaXT5/iKZ17SFnHHXuwRcR+JysoQYOWLjnNn41EOikA8+Xi5ciHX05bMFY++Osw
IQXvXkgicMKaZispC6TP8tYgvmi3Vu+DBHPGVxDbhT09EZU3nUjj/mDdJclkBwto
+GLpVHqSGGTGtH+0DSFT1+vIP2eIUd0hVFgDIUU8cyeondOws5wxS6YUIlocfpbv
ayGDUSGKD8gPCorYwETFEeGr8wyn37hPizsSW9YHMzXOh7FxVsNZp0uo65srYtSX
uU6x7LHJxmgyRVh1VpnztlcVA2NTiS+rS2RZhlH/hWQnrjkvYFdjcZrxxr9/wqxS
QbpzE9CHG7J11FDJYmlc16sEUL83keBMMqECA5bIldKARePYIoiw4h8RqzJvKwJs
mzDCsazPG8zgI82nala6KOYvYDRyN3U6UdKxIoe/lv/Q/XfGzd8yAw4JNQj6H/gL
sHWllN0aEoGQB6djVSTEX8jQlUvI/1IBdQS9/htAsEdI8eN51A0TZk/jC8TQLebp
Wqq6tobDSsPKxH6qWQRiLhiHorLIx14+a/eqdmTjpku5vx2l+kvkEkVEDC1cnT+B
IhrNFZBOSAKTFm5Ts5qse70DSWJvvXdbd2vWtOZ1fNAr/4FgDmYEOyzIXIGpxg4J
oKk0rsC95x23GY4xRq2DANvgXBwMxDDgceKeOI9w99N22m/XYMv3uOTWpzKCw4dD
OUFdJaFfP+Safjt/EKJXZeIRKgnrdlnWkNIdTzPAVGPGhgJZB37Q5Ps1L5qBl8RD
l9ZNqhks7uEz2cifMcDnjkpX89SVCFNWFMS7XBBk49TlOFks1vFehI5XLBG5QDWu
m8pritDsyEYOusNVvTgOYERIwD02CB77ux1MPHvMVy8w0vS7Y4uylbqR6k0j6t+C
9N2+VTVoKwVL29ZKleC0Go8fBBB8Ev6HnQdr2XhhrenS0pcmup/wB9Tup90rbo1p
FI1mTHshgNe9VaBpTojdeFpj+uA6S/gAyFpcSE3/q0t3LPimMCC/PtIWDuV597v5
Bm8RwY7aXzDfzXYntaeanFb+b6Hn/nIizQgtIyCNn5hKsc66TJgkAtgjVAlSp+UA
gvMmemaijgMgDHjXcsAZB42ZoHSZq+a4bG2pyiRgzUxfZwV0bwclxTSJV7JVfw6G
eSFuV0BTcB3h+04qb20lQ8oYw+l7/Q141jUwOPn5+BjrJVsB/3akhk0AU2UeX4qp
BnXTuGJdAfK221VooDYxphQroZo7yhZk9tDX4g3cNLUIL3WP2VbRTzwYwLJoLy+p
YdLhfhvwpeS6yRBnhi9zp/Zhb7k/z/j3vEQm6TU5Iw1Hn6Bq0X3cVVvhTidwp2es
hYiCIyHuDYOex1xQMLZ7B1q5Cd6PRIf/mNy/+nL4Hh8p7F5wlSQCimR1B90wuaQb
RZbrKGipkX88ZlsPOAsNY00CQYxM0ZqqKc5HS37WDNZFV7Z+WYdN9rNNZGpSymym
SBtYBrdOEkyb9k1/yNEO3MplNLUq830zaMfTVev33EkKx8nVAR0T+/zWW/z7EdBB
Exco80cUGFWU30HgUng2YNGahzFJsGWFsWBtwokBy9m1Al+IrVf/TKy1LC+i6ZKe
wY4+pqhAJjsyNhDXHjvvQHWODSdAWXtNAWgrqJJDplNLwxMOu/g7bNj0lGZAcYed
faFQVkcgmGhm2OsBPpk6rL0NUJHDadyLW4n5jRLU+9ts6l0qoUdL2zNBVzeQfd+V
IHMsQFtcbTkijbqDoGlhci2orbOi4Z8EcNCyT+WNa7ac3OJ+8j4RI/oT8DkT+jKg
gC5ktvQn0D99S36MkfFvhPSImqoXl0BXe2JW6LE//NK6+Ge6HIhl0gfHSgFsuogU
df3UPfvBBVG+tfuexd9cyWY+K+Q68tMv5uVHaPLRk8z/C+52UxkbDEWf0P7oJs+3
1OUHkxCbXiSBeTsR/sQfa32U2jbS8Q1thl56U92pg/5HjQHmanN78v/MZpLGjJT5
pT6Yei1mZwN+L8OLOz5EJVBBkYFmY+NzXGfbqwtu2T7VIS4teC/tponQhn5RqB5w
UxMP6niqtHfjfVmoYDzuO0UJRIrGtK9+iw6cWlzDAPOPlIOgcCknIeiYWT/jXjSX
BjfKIRaU/usm0QgN24skQ5eb3H2shRiSCwdmjuBgGqt5jX2dAoDHStbUOkQ1JXMA
nx2SpytqwcAzufqlXqB2m41ucfnw/XpLXZnBg+7OPYFEkauM0HTwmtWNJpgR/9V5
2H59Rlvj9yqIm8soM4vVqR/7949imzFBzMD6//kgIpT2dEu2jDhWNRfi/+IEWY0w
Ol4xjbu1BG6cYI045FxM4ib+xWXIjvemBhcsgVrWVRPTdEnHFgYM6CFzde8ol61q
BSsA5G5YCwHAYu4ONSGuvsWEIp9KHX7PXip+cSxnC6laOuyLewJFHpGHUWTSmOcs
arFBaSjLNmihBOmAvFwba52vgfU2etbi1CavZ87MdFW9wJbdRD6IkMcvE/0w0Ki8
+heLRwG7pBDEV6Iqg33/YRC8+ZPJSwVw7Q3iOlbQkfbulGZKP8F4baQjjH0wvKOB
Juc6rWaQrM/smMGyG3Yau5oLy82d/03hgLloCxk9Kr7McNXzGDEo5qTLCsJa25po
vKzTc82Yw/BPeQWcjDTdLlJF1Wri3g6nAjS8SNjmahsRXEFpuz36/RT35cHN4z9v
v7w4toLCoC+Nnx+PGC1BcOIfYnSW0dCfDdNIFcs3/J176X3mFDdokxuDQRzbvdm3
BmXxCtyzX9dcWkpw4PRLBRNxa5wWBTvuZTcRHCIW7Oy0S0ANpxSGHKkXPoB9CSse
V6sovumXIAXby620LXCkIPfISmsnMSRWtMKUUlK7iI4yX03sBOMMevjftZkYjUbw
wkNAPNx6v42VJela4TQd38HRZL6DSI1YHaEHVIc2Y0wGFhrJWz8cn4WKPU/LOPx4
piZ1H+GqQ2yDj3u4+x+IpejKaFZ7E/VSKWK2PryB1P7BqbkgHilBGU4WWfFbbiWV
cbOgO6VyDaa4mLsbGbntgtjg/IYK/wSJDzepKGDcxNWxgatGEQ3avjfh0+kHqm04
44ULWyCHbkW4zYTbgwv06L5u3sJonT8JwHWRP8ReTRTEUqGu7nk2PuGVCd72eYhR
aWZqCMnAHw5uur20OGnjSKEc/JwvBCGDGBZ95U6heE9NdXppwMlA82E/4eKKjVkb
EZOhBM2PfGiGjwHI4N6bIpE6NSMcJgvyRfWJezXu5F9SRMRuwpzFSvUe5cA/6b46
qtKd2e0GApM3QO1tTCNQvZf+TK3e+QSqzhruSTN9zmN4e41O0hCtsYe6jqfLfRbb
YoQiKi+M+5JZMJ3AKNg2dXkhIvVNd8yoxsnI3cnU58VCqkRE6CYZyOb8MaP5PFMe
T0cIZo7i7VSXAD6PyVMnPuP3QUoPgEcnnaATkuDc6UmYAaxRwNOBe+iJ27dpuSwt
iLrWRTu57tbbqGPIWMHt6xgIqTrNuPVJb6Ev9jHwZYtJzn/nX4DanbZ0QL1tAHvZ
x32AzhunTAnCFZnIvju+VW8PMu3gA5nVU8PylN9/qOLG+c3F/XQwr6V6TWiy9kG2
K5EMK/DX1KjFY3FRiYbzfbX+Y1xvUnIidgd+eeDqJ80qcicWmP5bMRomQTo+Ao41
p0Tbd9BgbtTo+mmtnVzXtMOravQv+VbCGDOhiL20fed8piZo+N//p2p8pZUDHILa
161IlCB+DY0FatscmQFEBQKiykZZBmN0N33YoPqC59IeaOqa2Rc2S+5G+yfZ7h56
lbYan56ZKxEotydp6aka5C4dvi7d0AEgoWajWKlQ3wyYDwWk6rhTjwWTQ7xML5nj
1WZdvaGKOK4SFN4cYHk8fpE8wl9XYraTukQNVVx10/GzFPXaacW9XnPC9i8bxHaB
E3bxdtFzJyS1TlfVDyk3N9z5U5K38IfGzUkEsSfyQj6N4S00Z9UsYthMw5otSMM4
ngnI51WGl0VZ2XrU7B3UZHUhRLoRXzOIcZ6vZGPsgb8yDTGdL7+W5tuusIjAgrsC
1tQ8C5VB2pzCvtAtbwmkFKMP4RtzdxZInr1moBad+xm7B9KfUO2f4c/bW+Ix8Zu8
HtoUZx9wKwVpngQiINJO1eboLVu/VIN3Iu37uR9bytqEkAlaV2qFZ+a4cMEhKj7i
Z6Nx+MUmqfGRpiWgLRk8Qza1g2W3vpZYuh5ABKPzOfxZJ8qyctx+p5b15APvmBDE
Fbg7IP1Zma/wjHMjGqUXHZwgeuSf3EH6G/EwzmpOhAbzs7567ZRBHVxxT+ahkxia
AbqKV5tG92yl5ifFs8PLnT3Gvgv1kXXjfrXuQWImeum08DtzOjpiCO3II0E8sGmT
feV98wQdrIZWZaUNql+Z+VTwdRbpW+lWKXpz5coCZjYdzOsAp5xQm9ywWcKClW3O
oZhgqHIq5R7kYOUivA82EdEGwB6ufUCZmwx812ImQMsf32rJm5CAak3jy7nCe6SB
D/U6F3HWWSP3WeovHJ5abGslfFCkcy+6bGLSSDKw6Fsiexnyo2LHq0ny8vuEKGMT
x9wzOlWuJNMri/lsqQOIQcZXiMsxLxDmsST2/0AqWOnmK8TyCn/2Tc6BxG5pnzD6
NPsdJ0fUWoRQQpMbM0+W3vw3h0ecsxWEoY0HE9yJ4S6u7z55Q1BmRc1Dh2XEw6ql
beydXzDnNpEBxilI67AvetL8oR1La8frubvkG1JRIerrYGTY+TT6ZCt3khWAeG7n
hUetrTwSlWV3ymfHX+3G2UjjTXbHFnEji5Dx2+a8iw1XJZDgA+zC59iDc6PLNFEg
K1iIxK3mk7wYKwuEMqskiyncc5DfEFquH2enn9WYLRkuyqKjPOX9JIBiNJTMNHvQ
S5nDpGRrSXZKQJfJjTfE4xmC+5fO0k/78SZj1hWPejj54blFeS+iecv3dZyvJ75p
IvwIKGbheU2BtruV6wVIn5Hd81/0QBYf/wKtGWOtM2c06qVzQsnOszVEbkTpDnxq
lp7FlDTYj204LlX1vkdpcSjOkcJiJfb1j5FUMNK+cWdLxBp2Jv1aSz2h7OmWx10v
OIUCPZwqH2ReNyzUVK/qivInh+htvNjPkiAoeKS49SyRmDci6ElISI8uyzVViK7C
uJTMGpkHbNe3sRiMtPZ+Qj9+INejkdk8/pWyJKiOQuDmERJW9qZLAA79cbnKtiMc
3s2NLNCznZmdXG4hdrA3W7YbFwc9dy5rO40W/77X7OFMeD6e/gDvBmjWj7F4APM7
eTXULQgFW7nXtWZbaWa5IExhIizpC82q5Jpdys4Q1sFbwVCsZOPgcTvsTqe4g6Ax
W3EQWVe6t4pxWFOOe8LsW5Ne3Acpus315a/zQWDZjwerX1eyATtr6Ay/YZiDineI
sS3Kee7vhqgTcfCJ/alqhUp2EwzfWJFKVfztVT0mzX24w63m8O2zBXJDCfN0A471
/avOeBONcBvmBQ0zNzNGamfjz/YmrH57VXYV7BZEzrJKG/9FthEPMtGNoZc0SFQp
A26U2eGbdy/TQv5mDFLA6AYX6bWYPsddRCWOwV20LpGlPkO+/D6NR9eu1kYW2LYO
Gf0dEc1UtNdO2Yl1da0Y4/yi2hvaZH9bQTsVUAqFi9az5dbUiRw8Hqt9X9+eCmWm
9I0TPjnKbEc0CElfvWQk7EaJzjQCYUfUhXSB1NnQhvPT1oht4wlTkf5c37ZgbA5F
EyDNb02Xyy/64MbZCVntGqsMZihJNb4ovDYY/lby0e7Ipk1G9he1KZyBhHzRSTp0
tSecGaMDPFgdQRq3RaXuU3SCt3Woe/jWG0f0A8Huu/LsmAIj2rr9A5YQzh68PZUm
/4ivttyzaldWjlMqzR6S1UB8MaozS7i68lgKvucz2w+7DCwvtAEcjWr59OwHsqAT
2X+co+1l8xdPU/DQz9Zan1/sQjPN/JeG7ZdL2uDcxZVzl4PITOGBKo4stBIxLULA
QVJ3GzOeNJ4wJCpHd2z3+HgCN3vn708Ub1zQEQ0fM5SbMlnH6ZD+kvoutBGjfgIm
jG1KTBVFmm1uxKk8AGtGen2YcUDhgJOuUbcX+Qg/ke+oVBVYq/BzmMxnLJsEmtef
SCJhmhvbBwdV+KHKGJrmCEuxEXPhd2E3yWgkqDQqOXDNfOPyk/kyObVdpgW28mgj
car9oO+jNmgcjxozPLTX8DiBjQE/mbJXAptZBKHfVPHjwaFJNLZ0dylhy5FAFPlM
H3wUugDn6rueKHPVA7i3dP+8MAON5yt5RYs9JNTog9Rp6G3br2+OrFLJwpPmbx1i
BCIo7jgEbj6toD0nUBYEH3DvYzWs9ZEadkOkExtLoB1ZEcOeW5Wt04HD7vYZCUxD
SouUvc6riurk36qaa1SIgpgokKrYhEEWH4xsV0wbZj/K7MnebDGDwj2+uE0ZtRTG
4P9Y5uxD38RoAceRza3rnW594+73fc34ao28imfQ1iw8BUolHYD6HQTmUbcMF+ze
tBQBOdL2uZ8yOUhZtwn2oUYM3AVeUtuOw2pK8Wt2QbBX9MtzMX9w2+f+OXcjLkGo
VuOvVQKzjQljpACNbr0QDJhNfpamEmLRZIZ9Ry6dqKvZ/19eE1FxlmMMZQwqzRYp
MC/6gEWg54AbQRDTEWSbD4x9y7N5D/23xrSNvLh9mnfSWwn/FSHq+XkJSLvgl0xP
VqjslKAxDA6fr/17M2JLAibgUZXdBCPDEG+mskoOs0sIWHWDlh4yt8OM9MxeNgh8
GyePbpZ0aDxE9Ls3sL7SiSbGl0O3VaIW8gsymJavHzc4Ht0y7I2YELQOACf9+ahw
BlJjhkGxaCVzMtQ0i/R0cFZYEUEZBc0E7aBpyP4dUG9puYt0aKpA4SOIJc24M2UJ
l3JNNhiedDD44uF3a6kxYU5FN3pLd93D606zlq19Lrzs2xuIbyDdOoIcb6fUH6JG
wQ0XwqtSEhx7SsDz7dkpV3OO3HdSGFw5TTMXIsor9+215Fkh99X3HGvAoKyI1bst
tT+kbSh83jx85BiAExKjBiRUwpp9Ze37uovLekiBs3XUPKzfRxF1H1R3l7/I2s/j
HpzkSLZYRLxK8FtO16opbBNXgCt+/Cgp8FpEC7mmwNVpkUlQKF/LKGrSd2MfA/Ia
cL8w3wgziwNLcPU1viW7kZWNSETJhB0Bno64BcWYXsoC+x8LBQRIUzXfzfbBp13g
nP0Viby2MrxGMhawOOnG+tY5irGXd3StwSVzZHwvTHfclq95rHmym/zPc2JfcrmE
v1tiApHP2c2W1bqZXxT8nGX1aRQ4TNuLo2SV2AZwXMEGeFVyzqlSpPMsDiPiBcvQ
DAlzeGcov7aHYTanLTRRmBr/eNkBVVNlCmXdqJM+Q6F+nFaTvu6W/T4MVA6kz0FI
tC5CFeubyn58G7JTUchq+LJLkEQWaU1ZRpfshIU9wQ8eAu/fP1M+t6VsyXxyiZsU
W3nkC9n8EY332Flf79xLMYTgqGayiX8/I42OCLA+c2ERM8tlcLBJFoIy0qO+gu3K
RBZ62VBwMXbf9VSYEVkbsyYglKneTdIM6aJp43VAyNNoF1WCJ+uW8Eiwm1rNg7E+
mNxjuv5o4JNYJ+B2005SPFkeJa9UfYbdc+BPFyVVDZKazNH2eY7wYMv88laCAj2U
5nDRf5e9DQRJQpaqbCfJHfN/RfMFG49UggsmQtb3oa94r9j9iTzuyWIYQI3OlpRc
2TaII9MYlllqtcNNmlZjZtxbQVT6pnDxe7+v9gTRZgAMb0dJMGTTgqo8zwzZscK5
93YmHUvu7J8trxRXNc+mE96CK70G7p/PnTMDOFtImPb/wcQ3XxFo98yBkb+P9BGM
lGeoV8LRRk7pZSp/lY2qAZyQno5xOKau6A0sTOLH1cQrWfGNFyvzSuFp6tRgrhsE
9tP4x/MrkFkVyWkwVpx3flCqydTJSeWM76biI50c51+1s2O8GW8akQ5brFpyieqi
YpTrvVTYAOHgINKV3BVBcYlxHr+oY2MgfQPdY7hie59uJgUfuE6rupnLbrUUe0eq
14SVBmKx0OeIyjzTwY7cijgoCl7rXGR1tnui0XdqukB7nFgapcenD33sQ71xo1Dp
lXj39Dx5QdBPjOhG3a1LGn1iinvEOY6wuxD+vh6zC7zjP4yrBZ2195bCX9Iv2yn7
v2Q2gfpIZo5/lhQUDx8HGKcaz77IFn7lxhCANwFiOP33TocD+08P7+Jwfuj6xkRs
Pf8ra1p9x5cnHcXNRYoxvNvj3CCj6ngPsWN3F6okGiKDp0+r/4ilm6GomOd/teKi
8f6JT6H/tJjW399uCj4gMtIqfaO//1LNoCzD9KKjLYZoGnQzjE4hrxzKRipEx7Xw
v5eXf3wETujCXkyXT7CzM4/k7Yx0/xhCriZNFbpzEKd9teGsZfup5TlKYY9lhakD
/BzUKgoB5iile6cMhZxsMXWzu/vhQiADPVEFiBuIxVcGg6hD+6tOEgqkVG1gpTsF
xffkidwSCOs49+tAkxc+jcKesfjnJJizOWtYqvzCWjl1Y/pWkB00mxPSshUBO50Z
MxOGWTVxSPd/AoOmihRTdj+416pnCbadRQ14N0qnhNQ+uyE8tGxOYZ82IzFPMirf
7/1v03+CfP9xCfGyBsbg5nArrGCvEoIHuQLBNANI/LdtXEQtSk8b12mpVFSd1id8
j1ZnvfajMfpmS5dYkgaTjBQwuWwOmYHKYgYi1X7dnNg1A7d1tR34lskz+j+fmAy4
8yCxbZO2+hhaqX7tfaTFlid0jQ4w9K/dAEarnovTeppmpl7UXc4Jgr6Q4ktKsvd5
s6z70XA9FUYyj0rzrnS8I4zbC2vxkPJZGz1ik0e837rdZlS/O5YoUUHowMyk70P0
+zzXWV8gTla0Hayu5wXDBuH0yZ6abuHE9aBhKDoCiLM2bDp0C4mnohLO9bo7TxJX
eREnQAyNfjfDx5oj5UmKOshfDhgfmSqWisWhs+G+KWtCi1HAMGYpEwjgldCWRL6O
jU4vyGPqF9fn3HMYrnWvTyq3JLr731Un6LNRGUwbvIHO7xrNce2AFae/G5gXt4cB
49mcyq3KInOOJw/fHBIi41YfnMpm+h/hvKHmpaTKLVmDtrGcQF+m7AIGffZTh6xR
erQsO1M70HGJhrUsA5vJEAxD00IlEV7ycq+rIy7628a54644X+yuWlY+tDJCjomq
My0mlBuL8P1rwy7P0FBZ1eliM198TIUSG2ZxnhH5fN26AqxBh/OdIIwqHIXYzpwE
qqumi0TAvDF/vtSAbTRaCLjBStMKWxV2VyuK90WSqrCPF5oOMZxRYSS86f7irmd7
LnR6FtXoKKCLbyzOVKHkNAv4O9XHG/y0hlGVhXXqdPRm8+TCkIR2iJ/FZKrMgKnk
LJIn7IbJxzsoNyPZPLkJPkPnjpKu3Cua/Rt49B0++jmPjsDfdFIpmhEO9IMplyRS
fdZofBOsEV/SIi7Ca6sZYNc84T25H6w+PILrQL/al0J/ULQs29LRAecm5bADBkq/
ZkapSfjm5ZbPzZHSTzNs/WnKC2tPb88GoIOWT+cgCct4OvMbHk/ESgtOsPtuyGXq
c+hCcij34/HA0SoQRHs3UBdt5qDopm5LO8G0z1qjM1ftCElTKt3jWtC/L5UZMaK/
CBOpcpJW+rXUF2svVGjUGRoTxTXrxaWg88r4O7eUsaxk7grAg8XF/udjJawIsVvC
+k993GupS1vmyzq9G4Oye3oWwqKw3G3907RK6bL+7QZwtoy6b7g8ptMMVzgkZdVz
9rgEaDyb625du6ZpfGe/nLt0fU10HOmFB5GdKcI+x95X0Iw2tx+3MuR3kD1gc4sp
IcCdqQe8/CmCeNQisZrsDW2FrmL47Gy/XntAY1O6sdTWYQgsFFirbMvkgfbPv8ED
fWPFfiGlIYdYNeCabWirxJgYugZrEX+FrMar/aQKlJ84WandwW07CQP9/03B5mLt
qPx2GXnLbPjDWOHSzQvM7WiPXZl6ydvDsLVMWA36d4KUYW1l9tEAxng9m3FsRbbQ
Yd2pk0k49I/zbAswrX8NUNdyFuRFane+H6EcJEqVvA0FM7piQxlZTE7Tjcw/J4eo
mI82dhMa8iSI4oZgVi05VWkSjIowZGXs2dXdElQ+bQBK67ZNAo0GxenodCNKgGqt
bcBpi9G+xWgm5eLSywJMSgpSm7dz1VJc7KWfD1D1/CbOQYl/11HDxl50NGQnwv2S
D/XANrk3NyHN4oB88jiirT/izo6Rf9vyg5SfvRULtj2S3JE/JUowYDcUAKIgHl3S
SaGT4oeAOICZdaiLtJiGOMxkI8hT2mdNYIaGeViDD4SV6D8rZ27M5oslNt5jHjSy
JgorAvXT1x0tO2denwKes3XxAK3zqrEoz/fPyR6bTsT25kHOXM1HZcdWtawR3R/i
u3CyOwvHdl+C5sDUJMVKHE/I1PkGPf8DwOh/R1Q7rABCr+DBEq0Sfo604oqfgsam
tNPKk053NRDA07iQcZvJDFrcTp1HUbVwmoAzDSIbVrRsxXwLNe7pUxM+LWfb2Lm+
sVD7flv0+Ts46TT8ycl63JBq4agN3GW5LXtcFhi/zafHjci7jKcin9ogWWFAlsKU
aYm2YjfvFN0xNCHkmFKW3K8lIiofSAlduMtv3NEbSTtNi31DBdeD37eqXeMrHjrm
jsxwnTpsB46CaK6qVb1oBnMwedaowSYVEB3Jp1ghrirY3rfmcB9f3/Vs+FVUBTRE
EVzoefo/2UQlVxelp+yo12hegUrBjfZBr84CxypSgjlL4I/AhjvUmq1uE5sGsrIP
ghYib9WJXMMQBviI7iTZBe16/fPD4diz1oG4pfhLCy7AbZoKuGYpOVOsidZe65Iy
5Pog35eeLyCAymGGD0WOb/dZAQ/XdyiVMzsWfUapxPwRByS4W4CXWb0KxArS2Qlt
5pHgR5zN30BMCSeUrBaJwpLjT8SHyT6IKJGtcbyd2vo7jRNLHhxtqQxzQ4FrsNrr
55xKrVrCSRFxzioWp9vwa2kLt6ljXYBFmf3myE6AMkG/SbaajRKFsEmkz20rzJ65
GUV2eJObODRXoG8PEN7jn0oUigAa3d/l08TcB8g9ZxqnMZ9gnno7v+a+XtICtIM0
MvGnxxiCu7xZ81uCVf2SH4QfiS4LvOVJ1Wo2Eg6ETZPmoCClRdCHjzm5i+Pb4FKx
d1peRXfPuPyPQ/HHwYK9UOKVnRjioqKEHWp63fKRJPyyM8HPf0ip804u9P+d3v4+
p7TQ0WEeaDtFxbMj48LFPvz8Srn/AiMT85VZG/eVNHJvGQi30v8Fxdd7tmvKvNeC
1LOwEr9SsnbuF1ilDcy5eRaYHclQ16HVhGLC2sJDuCHWqvyk/hT3DWXzfQksol5e
OJxZbRCMHDhzGvb63uBYJiUp0yb4lM0jGTmCz+xGPBltZ3evuGrdL9oiagiXE/Ts
1BsGISQoNHNe0ElPG5ysZD8A9bYjaabfHkzILl8G4XFZFM0rq38sX5Td3CKSIdhY
O2zhTPspvewb0ACmy7EDE+KhVSFExOo8XgFaYMhSKMWImXaqOmbBzqjulaK3GTg1
GvP2GpsJhljbDoTC8AaKMtO1X2aIZCc/w9H4247PBV1ce72VPH+fEWM5sg88Xs4X
KbSpXrBeyNiZaXf/vQOkyQ/+ZKduClqNFReAwdAayLqAxxBtRRG/S20kqsOUMPpZ
6bcrMbdtpJon50/bpbHFfelwwYzxpSHklbjQ1KyTuDKC6Q3ZGOr3YcHA3X0qnjAR
0pKVxSZiUD+Kjx+ioH5qpJ0VQSq5xI0RSXOYBiU2ceDTOyiGkzGF5HkjmiuSOXgC
LJpgQTKmx/Yi81PJEpNBfrANKS+JSwdWIpO+JfpG1ZyleuTz0z8R132Hvr2CgLaK
3OPa4LzatLxCzzYgT3JOkIodmE5+37fKQFm6ioVaoG20KcXf3GoEjKkbN4QQY8yz
gMkBdE3Y2qSpERGvOmODxYZR+dxHyJahlRyfnxcScWy9/F8A/UsIvJPC/DYMBSEF
XxU3dJPMWvICEH8uRND3li59B5xI9FuppMDv1gLmd+3foDKlvcESsttUJuyRl3qg
rIrdh38q4S7JZDoR/6UTM6EDcnqzwVZD/b3KK3GJ2bHTEwNeqk8PO89UhTF+m+eB
uKsdr/GJVNGc8m0AgDcwx7YcCQgeO3aFhXdOX6j3drB1ALWetPv1GMP2jmb4zw+L
i5zACqMxGu5zVXl2I8o82JCVqHjlYBIeETuP/KKav0CNQMKhWacXHNEf+kRhJP8l
/zzYmjK2YmXfkhD2fYsIR9kcUlX494ZnB6DUb0eiwUod7Vq2oLLUqwRIBdpv91WT
iE7cZ20H+dSSMwYBAQMX2w2NgiAvagM9n8f/ilAtZ0auhGcxB4A6wgcP+CLYYfeK
OXq0977spbHhNyhqc89md7i5o2WczWOv2Zog6GabarVq6knuFLF4ANU3DDZEVMPr
Qz9ihfWpyO3XGxBt4+ySjhKI7If6mvh72YWMIvq7WKfMfmZY4RCxay3M8r21vUmL
i2wSr5n9yxm+zpDbBTMWXp1Twn5yZpPl15987AC2ZYmHzUDQBI7A2JXITOb7F9r0
C0YKrnZL6LSXesQQz92siv2a79AyY6tIUo3FZRkC1lI7qQ5pg8LzrQxnHMt7Ms2y
OeeOVvZO9QDy101ZyGagryLkc4BsQznTS1zfvTN8TFHhVqHBdigHgi7bV8jrTp26
JY6OOnEFQuuoCj4TU9jIldkxwqOBIlxX6/7TieNH6CSnWdHlfLDUe/1hc3+x/Bvc
DhdKypl/Lbfq7hkS6/xswDA42YQEzJ32kaiEZ4eL/eEPhdJu+bmKs7royOK3TpCJ
wm9l+8edyKmLYIm+68toPt/dCSDdTAyK6U001Tle65UCOTRBNUO1IyGw0O+AY80j
w8Y1byMNAWyFHRzsFU4d8qyXmS4ijwKIk08W5z70Y4KuLclm5AA8VEh9AFnz1nr+
nWS/eW6WISWwrJMnh3N9GIItq/1DGPnFdAnPhCHpbawOeUiV4CumHVx93hp0h/UO
R0bsd5JYNUAkJ+VpMzgCIv1UQWva+ZTaqaCRXookK8EHQrV/4LMOBejOAf1TwU9w
i182I4P30u14zfrEW8cjZ2tehG9m2yLqAlnlQlJojoyiUZzUekDLMsFsiUuoC5Gs
AGovy1cTc06yrIqSvV2iCcdQRs2GUtN+7DbfncLy+wpT/rQHvv0RN+KpomzR5pIt
GoO38DkZh27AFKzttthDUeJKhapOHEFI8gGZ/CLqIzdBnKHAb809XhUBXCLhiozv
Dq5+2Fr3uDF/pxM6mZebg/gT9rTjW+xEq3roA+TLdNgkno39YFShHRJBLOVqkVc1
zlh8yMBaSMI5sF1beEiVq/qfwxKuHSF0eNMq3MPSEr6FG4qSs6T+G1HFDR8PwwQ1
Ge6NgwAanuvGXNW34ZH/wwWXj+RMcYQ7LnQYjDNeEIh6kt4FlYTQgCfChBY50W7t
JcsArysPQ+8aCsGt8c2dtcO6VBeb34cOx+FpfREJ6HegXnQhb+mK1sjjwZjm9ymh
apIvIUBltnEoPr5Y6+czUnVQudhgJwlBfY2SnH31KXvJ/mc8HEqfcXeDJ4upgdjL
3XoLeLmE3W0YJdrBJVHqVGO02wcXNigOjMZkRURHIRMnnNZFrzJ3cl53AV6lSOcg
+w1lONlN1LCmddewPsvpuyyoRPTPb/S26r0qIEHkBk80nY5DGH2TH2lE0cKavA45
hA6BPChv04WUkKNh9EH2f6aRVdIHstemCwmXbFwR9aqWJnWptGG2o3HaopKgjArT
XUgfGiORaS9l0+yiipruO2zG/MU7ZZMMtPUblLmXH2e+ifWZpwz94rcvTeT48AjU
PVBmiHZ2QyU3jOc68WOoJ18+yYF9cCIxBnHH3rECNde0abKlaVduwix1/l9PMPxY
RxVBpOdmqaqkYP7B9vh7rggWH4bTZ3EDDypzB55gmK3YY7TQoyqq82VTYtI02FfW
SxiDz9UJApRAId6jTTBcyjKZxkCSeoml2BEhIlzF17sH8tZUAmMDf8au7plJqOWK
Qq0iijXnylbhndGX16R/J5A34lxE6ZyXsIPmR7ZUQ+j7vVUcNJuxWEdTRe0xjHra
lFdVo4s74lIStR+w4QRCj7jaK8yqp8URkBjB+VjUNsswDUgQ9rHE2+z4TT+UzZbV
zCivuHOWl8KwieNlVUrlOSpbpngJBJXJ6cW/lII35wOuF+HqaJ7nBUc5lsv4uWz4
YdXbblPXOF6Ql5gxPq12KvD3MPHQN0qtqkVtDUi/7fdIS69iFhYV+c6dfv/CLG3D
bxoTtlJhtuaJXXwN4Od64oSBkdLeajUe04E0SoqnFlvCD87qB/WTEfyjuGUf5fnb
gwj2ew6L57Um1VL7co/Uk4ipLiD989Rprs5wJ28wFRnOS/nW9NNji7+kLwP5VGGt
HvMVuX2xVqytBYv+b5EedvcxPP7Uk5/wmZtdotAFz6yq8+OsszyjZsKZyRNPDoZp
hSnUg+0PqR8kvJJZ2vZ+SoOa2v3GNEOEQgg+CCQhim6JCrTG7oS5+REKHl/ZOazW
72l7pUHHjPK/0tGf9YeaAaDzylUcsUE2y+1qjUe2C2NfwikwnLILpi8Lr2s44xWu
y7ejSfd48piy2XyqMEuR9S9u7aZ7dTfG22FL0JaSoP5TXjm03lR7onrrI3dlGtg2
O4bq2xBXp35ONyXAkJw8v3IuMqOwKTDVwNLkxvYohFUqY9a1lYVv2OyzwxB1Ax+k
8gwgvjU7YOdxlZtwA+xl2AQ1R+Irnil/W8rhyEdqwQ0YCm9lagwwm4RQdWHcFc8I
09Hr1FdnPrAIioy6PSs/evCW1YkRVfbM4ExyzTA9pHwDl9IQLS5niQIf9qjepHLR
g00hIRJHmWHhJUqRgTedQ1LKg12w3scT/DrMex0IwU7juRavW5fYPD9ORsAOhWQG
aqASpjxlBnJmdPf7/xyMEh0tU3eUb1jStvU79AGes2+Dv4zJ1d8GsdGCAc9ZQYFy
Z/bLKpJmsV18+ckImpy2WO0lOpNRbePo9ecN67C6DtbpkabOO8pS8qlIVq+Zjpng
IkgN6WMTdwjT8E64lGEAbmrLrbCO5Tiwg+hCOS4nZNPs+Fwt3ejmXWpibqkGCTYt
6PnbRtybAlETnRxzQffe/CPPBKITT8yJrp9ZPeF264Yh4r9B10r4uWMK8Tv0g4ac
cjNyTQOz5oHzQm97MM3d5hN2CEDqEWZWcrDVS8s6Qm7A3TSb0CM2P2N5f7H6JBbM
E+j3O2JQzSQkUFw8mhAriyrqT7halCjbvJK/6NCP0CQN2Yf6IG/5GtdcLmksxTyc
rU0bbsgG5B9qa5NnoJaCwuCcYA6N2af/V0DumMk5tddOuOx9ImDeIrmH7P0SZvuT
MPx83fLvEVj5GClyzVdHoKvna3yd7touwgacYIV8RhbSsvP8Hfu+OBy3qU6PVGk+
pKOplSixmvwCYwy9kNVcIIJbWxxiTtbTJ30l9ueVZG/cwjR8Q78+vVtHgGA2F2k1
qdCm61JIHIcbVd/ybHVvbmBP394NcgSYDOdKjTRRt3tsRA6lLcqDtCKhV/IC95mA
GQ6wq0/7W6QB/XWCPCaStm9YQ7nv3N7jEXA3Ep4aRfPgljjgppg8sQYOP2oM68Uw
k2fTRAOMrGB5pgxrLE+KqZqKuNXoRaKzTxYndw2UA8bnvHnlg02UOi3Ri5pTI9O+
ZLbJKT+32Gn0eL8oDKL/y0bW41AgqNVkGa4oZth3F5/SMBUw2U5z0ew2hcqZl25F
L/CbshRCLxa63UZWFnol/bwnfd5+NsXh/WDmI6EOnpe3K54AVikPudxaLKN51nf2
dpyhG93vRjihPyWDJjYndbHYQnKknKGJb6U7xx4h0hz6f3e5RgepPpLj/7MgRrjb
ARPmrLZJ5x7KUgQQP40Nv1Fj4O8GpQKKAh6w0HLZVRTxCISffbpbH3Nl36I0jFHs
yI6F8DK3Lb8IExZyNC0TqXXlbeldjrphkgN19Fcv8Sj2uxh55tfqs+mSIs/9Z9ey
0UMEZ9+qcvkiIWJqkQN+INGmhMidTndm6YJnDvu9QV0S1fAy6UhyCS3QahSZY1LE
gv7vYVMv/zThaEo7HoCk2HzUIv9RxbUx/C+Aw+lcEInttMM1JCeNKq8pSt5hsHFY
meWFUUpLv+8NuhfOt4zWFIBWmJTHEKfpKO/mHLwPZwkRd55VnwioUJ2An1H0wI+K
G8JBjWh/qXdfvSHlOV3ZCqjjksaGlyu5w0BXBL4Jfb/obhk/ESVl/GZdfCTXCp89
aA5nwB6mTU4ux9kB2wVOqqXRlUdbTSqoV7XpsLl0G2WKdeIu+pxvOC9zUCWzxcmb
KKw3AG6CZCfyD0Ay/OdnnxpaknMpWBCtXwweKFyEIkCpH2ZG/87SUdMVo9l/8ulM
/vYxPBfL+DnY3EBD4s04Drcgbc0dWeJYFoLfsF87qhL+HO424Ri7hdnb5rJqd0xj
TRuImWspBp7QwESu62RrcY6xLmTWK+MxKM/VK2M5T9lVHjyEdLlcZnDO7z+JK0Va
n99347b+Sc2vRIuoVIY6v9pbWO0thaGODlMLnzIZjaHi0EKCKVJ8aHFGE8lIcUse
0TvqcXeg/6BgcRpU6X1ZBByWGTLZMS4dpAYIDV0dz74V0PpetX6VQEJWsLml/qk0
IUzdqoD90y0MpPL5s+tpHycWd8DoMIr4cLyjjCXq/Xz7kvaPXtYSramU8DTdTZPo
m4xud7Y+ShmxTeyFKU75KG59OAWSoMVYhPcO4yqEBKgl8bK2lZtOc9583FXPf4YP
G2ZDw5ewJOYRpuqMnCaPJWDzliyA68/kClcZ4RJ7GCJ6Oxe8UQNzQyLVgC/8WPc0
R/aJ9C2Y0u8GVphWOhPgUMLvkrdDB9l9KyjC/LcyLQgopYkpgTbuvPY0Pnjt7Va9
IZIAq1lgamVU/NoUhJZzLEzPrNYLRtoCD92kECVSd5QWYurZpyHeemWnBehDzr6z
gMbFf41QVl/GDd7D0IYy5fdp6FLnjXHqtMkhOUQ2r7W/2piduAU0fZELts6GlPCp
jWn5vUVSxfHcO/4KXbOWNVhM3hWbWtxi6RCH9+0xIbuJBMys1SrEFJAX9vouRx6q
deslzm1VLc6hcSuly9v1I2M2gy2pfReX+zLKGK5S9ORhcYqjMl4FcOIlBS2O7spE
wvh9Po2UsDoFzDRcb0Z+stPv41vOyaG7vgO2oOr0/qjSjw6kNoAJpCYmnhpRKAFG
aJShzbcy12zokGseogVJ9DIsG1Ey1w/fOKpDoknX+U8WBmRho/ETLxZ7xnr+2VUD
OluP+ZG/PWJFv+3lCOk4DngJokYGiOaaeKJp0DYdim2xqiR28zySCZXjjomC2AXl
jruzQqsER0FFW1l9Z5dCePRiBMBsBNWztr0zVRdT7voTI3BMR+MxhovNSjMxVQ1A
Xqh2zhx1rruJGt3Y+ElWuc2POVLuQmBbY1Fiqbu7ngsJ++mpEueBzbWav5En5XVb
+aJaGMWgil+x+0jSeAdSwf8/6D/ugjR065g0CgcQo9rnWONsS29BA24pIHTiy9t/
M9JcxIBInvwwFG/S2HPnFX2atsKW69F2kCiFhy/p1rXn0r7Sjp0ueQQtOp2E7dCX
Y9i+w+SLeDAaBNkN+QRDoBmC36pQV6zu3FoKR4zhFmv8h1ttZiDz+ywgYAaNW19C
uRWWZjte2nUNyPNrOVzPWJOAVnYjgdEdC/04Uj1EL1r2iUPCE/Wu6qnvK4u8W8L1
+MUYxp4gGf7/9+Z1SOY+oYVTb9MWgZQNSiUg3M12WxUa1uqwmmCr9ppWcWFw/GQC
7KasffJdZH4zlTqbeYvX7B5N9ovtJ0FvI6v2jJMYu9RdUZwaLtG4hxJw4Ff3IKne
wfjXLxzLslQHPlkiWTFFuxWNAHityM2FP8tiQ8tMM7/QrDAWr/NTlRvV6PHe2N5H
1VnqGjtG3sogH2o2m6dWweq6CNNCiv/OZNXCsZDMEF25tJBV1P/MIozyum8uiWjk
EYJRBTuFAi88dtK41bB+RB1NfKxyKPoyn6z0ObB5DkcZRRfshBOwEXiR0JlVkjcQ
kk45R5R65kBqq5A1IozHrHpQyYfXryXfHcdcclZl6lqfwmq5nCzoG6Ff71Bjd5Y8
SSj6dWTn17XI0lkY32nvocN4yf2tVjdMcJH1ObE5vsC3lg5xsYkcoILARz4A4X9f
eBwoGW6nn4paiz0Kzf/bWVrxngL6nyOcctdWMGBx6jl9wVe8eT97ZXuYYGJYVyf6
XQ+yStdx1u+5Khk+HeVtB6SPTRG2qrwJX6nbM+zRLG29JkUSg5WHFNZ2Zam2Jhuy
7NeL8b3MN+ECgFElmD6S9rpQJepYi0DnEiOz9Q0UHpN6Q3uHDNqZiHIBGhlPkt7U
t1nJeDsK6gIhZWiDlDYS6VCSZFLr/P10nWCkfChFgrYWNF03Frsr2cUg+pNoqwSu
44vozr0j6ZXkUK9gSYrLCQbwra7glcc3sGOucmaaqoqKzszHZiIMVEpNxUmerCSj
wU2sG/PmVPMQbf2aaSz3uAZJ2dLq69MBEJhcgm4oBwFxzgzAkPZI3aTMSZO/1QkB
XVky1XVuATVBUsuveWTi+11S87eTn+5o/oaUcBy+H+9UyR6PbaHo+vWgAg4nRr5P
q3TPe0rZf2KESe96j0ak5z0TexteyjewcU3E/EuYzJZr6gUuL/1bkdKs/C4KpbPf
Y2JZCneYDC7hJaOZ9Y8g0GQqEkmAg3oWb5vU3BNf6CaSI1pflplCt01+rRfSzThz
EtzV4GbMJNxT5tLGvPrcsPnr4aiEBBsRBIyzuSsPfXtCfVwhXEhamrpEsPICVTqX
5wYCk+HIGnGawZqsbRLnrVj3b3PPASKBMgH5Z6ocagwqv6DT9rv5lf3O5reuo+/e
7ALhm9ffPj6QCmgpoRd2W0/iXL3YoMV66cEHxEpDUZ08MeKY33LVQyLSwI/GSTm/
yadbPYMYtiQbjS/74mizz5Xq1u8pJHNhWcrQKiUxI90XlvFXxM1LZ8Fd9xmHF/28
k7NpEI8mtdHhP/+MStXDA13xyCvRHITA3kbE5M7PJeUXRzARhDPKr/nPEv7U+jg4
eg44uWt5uJcmp2pqsgeZM7Ul251ObGX2sR6JzvCPxdwa4HRoW3RVSeyjpU7aMtqA
CGOdTjX7KP5eLZzY2KzuSyjgyNkosQYAT6G2IZxb8inB+wS+QvblpNpFUXVGWMqh
t/NplaKUMiCeJtk3muBpHt/F6IdjF8MvG28/Rlrl41VJKfLsbeqk00acLhoP37G0
C8srDkAY2tMfR6Qk1vXCR59aj6kBa3GU7KRS7xrLMV8U5g+g3NmLdAjvHZPNkeZ/
IW6GRhQsd2FLoZzmuLh0iwyvCa65/JNLqlFL5iDc2Lm9m1tUipiI9GjZtGilDBso
P48gJk9V1j9mW29qyneg+D0R0YT/iA1TY2W6fl0wijbsy4hUeuugyJTZpDY8iyaS
ArGffZMeB4cIthIbPygyfCG6aguru1FlE9RigyIRPcOOiWxa5VJcwmC1V33qnxbI
KHN+HPOnVEHpx9FlP+zDJf8QZJHvzZ7vCbUuWKmskfSUOO6O3l2ZA7wcHB5UvBtK
UUwM+x9KyTrib837NuxShBigWkSa/C1IIyZvMhyVOFQbFQa3Hu4q0wh++Pvbduco
5c39ZIZ/1PmbDh0adHuAk/VGIibBV/nD67Xk7jstZmW99PDPCmEi1eTmjHGrgHhJ
TPOUHBf72qYfc7uPk+tT53fmMjSme8hBYdCZbFYLFUbzjT4Uoi2u6Hry17f9miqE
tBzkQAjex+WuNjVtlRhpvjYAb8kbz7lbIF1YFIUskJf6bnV9qjnA6nc5qkMXoC7U
fwUntl2ZTONQc2NuQzRV12+ozjot3drhr3MXCOBvkoU7pIKZs55VznquBqs4QvBJ
Wg216woull09SHwBPybFoUyYlbQWBZib+K1veupl+vaDr+J+cQyyH3HVlxL+LptC
ISVI4ZtVWgFkot7bUpTRpf/dZWg0XH1vmnk9uQYHsJn1iVaV3/yOaBEKAlJ9lNA+
ZshNjTGg0Ui9e0lQXvt4eGfZcJ1OHQRks9zYffa+zUfWWPligEmMiXG/NIj/hCI2
4bOJ8F8SBhECgLqI/CdEiRF4xVxLcdfimqV/U/lntGpmKadxMgVqNH+QCZEw+tIl
00l1BE1FqGnoqWkIBhpFiyGg2NXgay1ULY2s+m/yjXbBIHmWsSEWu7+qHgTeZ4B8
0n79mfXLyf0aNSDPZvIZluFj3DxWQLVjxjfHcq1shi1XHOcbYLJ8bBQVb86Ue9UG
W7ameqWjP25EInYlzAOGvloXWYfC/JuflIkFy7yeMPbJCyUwgF+vDjs1OvMMD2fC
KBdyaNLUn2HGT/h4ZJKSjhht9E6gH+iIe2wXPZNLw5fkG3tG7VOPf2KHHE9SvK7e
bfr9jVhrvCuQ18asTyyJfZzVVLI5YQX7GBZ4o85qOn/vcTGfK6+cw16EvuQ5yWCP
3yCUv414ydOVmKtgntlKL1gWcywYEqzW/wKtic+kMZafPNfXMrd7xspWJvoz4zKC
UdpqgMjaEEakpf7qyBO5fDMXX5IQySnxz9UZKCkMu2Cc+3NoYvxJ5rSES+wh+0Lc
FiMkypolKEHjmNRQgl8t92nZzFTV6/wuzjBj6BwtwsJP+I6NQAY+tmDIzYWrkMcm
0W8sdWhjZ9xKMO7zu7WWv3YeG5rogiw9sL/WeeKcDmUg5PncnoceTOn/GS4x38/k
QrwyFsnzGQ+iHl1RniF4FazqdiuBo/V2IejqnFHH/4rlUIZTSxT/aBssoBD7U0py
/ZzTENswdlEPQujNy83eDwxvBPVJqIAIbcufPw+KaumfStHF8j16cT+mArIQd3m9
mlHjJFGwCbm1GFcNEF0IV8Uie4ktvrmO7xwvMXkuLX4QclbYC9HHjQU0Oj9fmVOd
aWoryWbrU6sllSdYroah9ttRf4PSYtFvxKjbMarI30Kjl8tJbafF8e/VIIAMvx8k
NO9WSlX3cAxLyAt09pGf0r7i1h0qHxE95HFWnGc2a4kz7TL/CXgmg2xKDlyqsXZz
0KwnD3hSzyE0+pf7VT6F7XhV9CWQcqXLi2LRbfgMscX3ktf/t/srcOcqhNiTyG4r
GXuxRS2GvmsWx5JGDfgGmtcFzA/ZG5zuWU2BlmoOE/nlJEDW9ov8/CW9P5Gj9qwB
C1/IJKU6biK3BHuxB9zkLVBTSCZzjvDmWi3bcWZ+wp0O6WOdV/pZA4xnpCUpPm0S
ka0R5tPsZmV8i9dvrrWpA/H4AwMsZh+HcY5BhLaSFwAZ2BKz+GRqfoBigy68+edL
SEdXQuyHPJdcUEV1fk7jNHL7LPu1iF9WykbG3j8U+jUC4u/daz1OSeuTOIk04xLZ
lPL9D5D9iH00fhVAwr0YX3TTyuxmlKTwPOxvu6BM/miU+wlUtE+MlHRsaGIxmhBG
4hkrf7ST7n6A5Yj2N/XGdXv4jYJpO+GErv/7qmAJO9FI/hW+eIh7cQnougwwSQzn
vnHBM+8UBAiInwkdFukPyIuHzqrL9FrnA1DfrNPgr2H9dp/ZARWNGK2bJ1aoVmcl
M9Jti/v1zD/HKAc+4c4H6xBSzwMAjDdU01JULOyCzgCl4/NPTulzrBBQiTpsgMYM
d3VpcPnLqdyctWXC/PluHmHyRtCjOfMwRXf4n+jZZe3ucUncBU3C+nYewcNF/N75
lLxhX/IPJD/PkDVS80v3qDMh8USoDIDvC5hlJ9qalYWcOerP5FVx1ezZfR7hPUyK
KUy1Mrli8hk5qM4AhdNwhsM7QvzbMA7nlp9QUK2lVuC/rvrN9Sc9LlIna3YM/Wq2
eyKzkvBBsL9zKMsg66VNDxB6SO7URJ0SwudbwzG9Ch6uvd4XAvfhqoghYt1LdmN6
M+1l80gdUz2BEe6XRT54SY77OLaj7OMdZ023994O1UEV2A/Cl22wUzQ5Ng57LoUs
hDeTkTuC+SGn3nx7/YsVWdAdLxxzBqWpKei2ymXgRVgBxIU5KBEecRl3TUoAx00d
4q+iIxefGslj8zjem0j3MU2C6MoyDRvHbnkR6/6jqeJhOloL00P0kAnLCCBATtvz
3kRX5ohfcDxyLAxEZVN+6XyY29ePNJKQBYFD3c4c9ri58ggoRHqOYrDQsBPbBLe2
EkMOPmsM7spkr/K3wUcHxXqMd0RlKM1Sgo0yBPQHxBFs2qqmjdftp7SbMuGX0XGI
azOk4HhAdd7vuUDXF6gsr0UpuiURaVag09ePxOd0EiZ5OiMX37mV+ghTxw7ipPAJ
KJhoB7Dsn1LTGym+SEEdXXI/Xx/uqOS7LmBwPS3vEMHIYdAU/7RCmzuoh/Up4JSL
IoAQiPZbGZQ/56WMMAnl8m+Oy6FFJE8627WKRlRrXLnHNOP8Y57u7Czvq5ei3pY+
3wNtkJ++D+0HerctYkc8l3IYu6YvR1TcFhcT9y8zQPwm+kjffLDJuTo2jEPWtz6T
QTxPn4wwc1Bj/BlIwI3mx6RtoN7hE0A5WW9Ybh9sqb2V52pFURF7eRp176Ll19Ub
x160CDzGyXvoEZs6halHR3Rc/8knWHkIzEW3R84omNsMtXTo0nmc835mse10/CGc
34OqXQY6EtmsXLGAZqB9ir+HTF28L8A57bfvSmVN74CSt2RyAE2As1ItCizdzI+U
9vcKfWGcnsqBNIrCRZzgUdKKjKu17CtDZKxihA9Fj7lYueTjGVIUYT/HUfCBchgR
cAdljeYzCTg5jcwyf1Fc5C24rF7DYBMS1pZdhN0H66uQiFvV7MQCpgIocAloKbkA
6FxOAqBYEsxgdVDggIhyGV45SnXZE0SitQ6H7eZVMsN7QouOC23efTwriMjXRRja
5zE2A3k/aE8W3rHjcRUdzz0y4Ofz7TtIMMAY1sUFVvupik1M1AgVMQ0QwOu44k5O
cKMxbkHJWwr6spHzZ7KijnvP3A0MAH9VNOTfaK7GaTasOvpOUsLeizDuTxljmpq/
yP9iZAdJuNx2iNVufMcMFTsWbb+1Z34O+e8QbwkgJotr2gJj3XDK/vO+hPsa36Hx
mjojhWo5Ui3cz2m/5kR7I4oSJO2M1Aa/h4d12pyQLR+uMj7KXkrv7tb4nZO/Jq2D
+S7Mb3JowQUYYwJkDSQeV9NlnbqIsKc6bzob61cTLRdPlg/liqVlqMqJiyQ8CWJj
p+u6svWFQVkjCtpm0v4cu36tfoTd3/WgU9m6IJEPQiqTC3T8ZhRWNZ7AwzK/v7K6
xDLJl6E6gCb0KSnpTY24Z3F8vyeqnXO+jOHgHIom8RzR1JCr8CWuWb++vOiv0hNV
XITZCp6tQwVudj4FZ/apN1rhB0y64IWadj+gp/DgrUEJ4Wo4vgTGMgkecyAvtmmO
RsCaf1pGVbfTo1wai+EnHufNuU0OfWB6QMdmRJwQz9AIo27IQZxa1Ke8mIz6BjAF
OYTg3FxRMAGYiM8x38pqsT9A9/Jr+J7gLxyAU9GYjiDjPRtr3V2mrQeF/RJRqzX0
gmnAPHFuaRb2jjDnjis+bXB2syvBn1A9ByUsrhja5aXMEz1qyyHJyXvdjBzPrcvP
as7FT1EMm4tNdw+zWvqN8EiNq7XrWNkr9muAozNbDYFE4yCNCjN8X0PTb6Rxn96e
1xZZclAKhslYkjd8+w7Daw3FsV2FAQV4k71GjrdaFOJVTRu197w3gDDrvh0D59dV
HMCEktlmocRCl1O4gX7vsOF90gFDkvKPAGOb9K/+dajQsguCb8J72jlBWW4ladlo
GeuflOr5d7olMTqhZuGeRkEPDNn0kfSKaqLB/wqnKFpoYz4D0b2j3sGb0Vq3Jhye
HZezLKodwk6pWl+K/sMJTc2We+BE/DOYsBHMQGgw7oe+umL7sh+MxBrBNmwLIshS
mMcFUV3CH1W43NbDuRDSTVRUE92dwOLxJx5uTnPsbVfcwRmhw0ic/ca9GLJlIIle
msWBsQ843upzzlQWeKjvGFcwe7utkD6RnpElWBZIjjVCUatkXq7lJWj9mZ0iFQvx
IzZCyX0x+bReFuHFy61dWdRC65/fsT/QVdIOApqv4M2brxHx7Yvu25kwd7mOCB7x
yIi1t27vJezEjWzoWjRb7aS2hji66NMmq+xjNvmQE39FO4X+ivoSuTFohSsoBzkS
Epx6I8eCXFemySwFxc9yjSPNuRxgEIRPwdVvAmunr+g99dA2nsS1qqcTU5VpWWzQ
rlIYH09byw18L492eV1RW5evseS5nxWi1QTRxyY08YVwDA3lZWiUoPPLIZ02k7No
qu4MpGgQr80r2vGESqxhbiIdcXlhQRZ7PYM6FOtPbQRQMjVnFH2K9hTgNT70vJWW
Fl+7w8Czg+9ABCZr3SxUvPTEIyeA7pfP7VQgFMoeUrAHzCmmu9E+yJWFhre/QRr2
BSADPAR7ujzKs3EIWBL+RJ/4LJCa7gt4MLrilPM5xYIUK5LljEe7hPsx0xqSc+1p
DjWpLPYOGZJUlid8j6QXVCdNdK2D0uGMiAcaP3f02D33w6+UenAs6hmWowaugQJm
MrVWp0EG6xym5ENVRntOj0Op2HBhDsokY/aN3EzNDH0WsexqtbNnh8izwytmnlg+
bULJvtfadIsIc2EZ0uKDammQXKclDkxTCKZ1Ayh1g29NshU3DW4SFscVcBDHsyKM
TdKFZ7e5HSYH37UWL618FT68AUe6dZeXeXXZck4TAJ/xgxHtOnSEnJ/YuZnjDuan
sUgf6ExeKTXhTi1Xh66f4kuwhievLT078kWUaOlzNRk0YLBupGQZDUSVI4rDFPKu
votsPxlZQ7ivYtaMwDDgr9Ed2uURUdakbs12YV8sGWDVsEZM79cfQA4eU4aufZhk
KPbRZ0MayOONhjokPMAR7k385FpR7y9KhPK57HMbyL5qTQGNtQqtD11+1AZB7Iqq
1Z/3qpfdsQxmsfV9kDUFVWvTsqJtmsjmTb7nqtGiia/9nfpzf/ipel9TgoocQqkE
eVg9AMdof75+AEo21MDLDjYEIxA2tSXjd9bAUBE60qwfcbic/3ozXNwkxM/ypz2s
onh/8IxpDCiaioHsYPb6DRBHMDk2C7NIf/IUtT0UsUmFZtIymz/qHSaiZPAQ+2qM
iOcsRn4zysnITZlHiHY6YjgMEDxKvs8dyG8txaIWg72dlTG/CwihlveA5HMrnrXS
6n9FlJ7WB+gR4t8200MnKb+YVwzNgVRQpzIEVomelbQXSN42CTBLZa+bAcKYCryA
zWKX9XN4iCcj4lICEIJAuDjJ1qs1Bn/HbNfCObHKYB6MTfqkXHGpBy7frmNXslvS
BB/UO36OW3MUv8/9l8UT1TBgEdLXAGPzW0x/lvMa2z7k3rHH9/DQUU000S8QfjRr
eShGeBSeo3NssQEvizjr4mNC9cDDGnwafspLqoFJYv+hs8zSq59lvmqy2JTMPfxV
6dFh50w9k3LWu2SMKie2nFDFz9oVf8wjGgHdUWR6NrbUGmhQ4X/5X6E6mCTBETJm
/+Fx26mcIcEwx4b/4pMGQK4jNbClujyj4SO4HY3wopj/mtkhKQPHM+aOMnrYB/Sg
PCt+2LJ/EwJLONBoUFJU9XwZd9L6wgHdwZ5KqogMfaIJ8aItoEn28zl889+S445A
pbW4rgSOFvvXjVR5wUbPVubhSCTTP2uLvuksCTeG0KFwqy93LRfF+h5tXZu39j+m
ShK8hMxj5SMA2EvwE8IPTwwjHqtqE2152zyd0LjGO8ZftvfFk2IJBhyEkVOQ+nbP
pPh6MN6cl6tkqEF0K3O3NR2dHwwKDhU1alzJgZyrBTkIVz0O6I3rAkDiCqkdMwx0
daTfmTRpQOJx/+DaJOl1ggR6VAF1JQNi8Bk5RKV/HWNp6V1YpPTUVkUmBVDsjsg3
iWSKWqtsEu9aaKroChWzC+FNjL1s/A1Jk+5P/6q84cbyVeGTHv7/SFL/ToO1gvbL
rsxOpxIwfel0vmyatjSuHUrRIF8pcKem7ng1t3KiIVfmKTUarUKzECp7dI0f2NLk
upYhzr4ZSzzHKFeZd9Ri498g924qOSLI4hW91B9TqzKeUbKg2/9jWSNysDiOtKgE
TKiJsU8lCTFa5MVkJN5Zd9D57vsm4X0kcUK7zPakalYSUTUnyYESkNUfVidNE0G1
s38xMfLkGIaU5rQlkVZZHok/T+WCIQiB9HBGBe9BBB3GaEYLU6EgldcEVWg6fiES
BbZhyyzxkhl5S6FoYILcXTM+0vRiuZzdJxCSzS94pNNBlCc/wE4CZypjr8rSgUk8
JK+vS4Oj6ZeULBIc45UXCFLDFnMi6jx3vSzG+VryCI3GEFJuRUIyGVtKjz/d0rsR
vaap2XOMsGPlEfb7S6XrkX5XkNpZZ39Qj7FaDheTsh6UC4DYg4r5bALQUd2PYt3j
kDWs/OTOE6rwe3CIoClVVQFo1mN1XulzTiXFqs3ML5I1nQw1WcAxtdOl28h5uZnE
U+MuOl13EDf/y2yDLdE7x77gox7eu8demmX46qMz3sQBDeEvjuf1ypKTWM2S4Hik
50SI6tKHyNSbT+EAyNWGb/dLBIZW/C3m6yaMb4Du5/W5ak2W2Zty0c2QXmj8ec90
jtwn/zZORzKeWlUDD1eRyljknc8b0fop2Tcx0NEv3FzU8yEae5aqWtbFltye0Uuq
A7TBWmqeUSqQuG+61hzHfoigvGPBHYVowt1RaAYIyx1Qvo1WrQOz1aDl+SuvqYb2
qm5q1rO0vlq0BWzfR4eoDKn0gS18Y86+RgnifBcVx73UwTLG0MDf4wHcvsw6Ctfg
8VWh41xfFtJihcwmDwMHCgePx0QFsv8ceMc+DY81p3UgI3r9QlyDvHivu7KehVGw
rXhyUWoNauua2RbWPePxUFIeR0GgT2Ypl5MiR6l5LgEGdpm5eCSyI1d71lKKMYKa
2PKliB0AAvChdlRgTM2Hn9pMVGuMnck3/1CkpZS2zA4NfxF8A+oLWiTW8HfPfx8B
bmZ0+ZMSoRRjNsLt5fE+I/bV6ayShQvjoH5lpMG9Ogo5BKmrRaNBfwniIiz5GfRq
Ca7EUfI+75+ghsjqyFEdaoJ559DoiYPc+Vy7GRHz74cNGTdSumCdURER2ENaLyK/
8+VZj74S/wiNPVZYwcjts5w9qMEdh+GwOBul4KicOmlYuAHImwRFVTWCIzNmr4QO
VW24NnE15HsWQwRcaHHMYjToEgrMeI8CQuWQg0A4SNAtQHX4COuUqCuDts3n1ADz
TCoeEouPAQkMLUvnBAnwFRkCqmD8nOwBc3ZaC7f/Ur3sjSenIc0OKBxDzA1zy5pr
z2g2ZkYMJu+aqduo0RJH/UvUVGbSzVpZbm0PN5byRgv9w57FYrY+DnuNKviKvQUn
+0HBz3XnllpkCszX+bfJtoS14/CI9WmYBAd/A1LeJhEkNM7mWZeiUHd3lcFy+7Mr
3N0Bz4mzXLvJRgl3d4VJRkx7kfhWUzr/+IziTBrFqAK6dLmV/z53a2N4+xNmFSKR
eWvRbSxWmCdBsr9yEXHKSk8nI/Bm4/LLWJe7lkCyR9oxnTLCRo2BCXTBwo89akjT
wGUfnKjnMVKTmjqSEBlzs7cgV5iB7MuXmGJDJw8jLVmHFXVwL5iqmPwAqmft+82r
o9uV+hzeJY23rEzC3w8XIgBCLymiJjsLT38jg+iyEGOCi0kFvvBc7+ouRvPoqLwH
W/+2WQkaBqtUNjjju3KKu8Oe0GNd4/Hsw2/+opIJtmiXmogmSXtClLTC4OgWATCB
zalwtrJTLxAzVNtDJGWkMsw7CjQ7zLvn/Dsu/8vMxPqeNpEaF9ZvRvzhlk2Mmo3K
Tq6Xmzp5lMtmKRY3Ty0N/KjuHhHF5R+O3EcoYgcOmeLWUe2sbKzSzpS0Eb0IaFju
xuux7HsBWqUddC6Ke2mRBrp7k4AJ+YnTGReBhmdxCu589oBL0qNAx+4gGfCISbob
hIa4pBpOoG5qRthNhwhenVTGA+GLncPpN6d2qBVDMwy+UXBXQpwst/LPgxLLsTX5
LE5RNjGCgJLvftCbtpqiHxtov5v6MC3lPjZ3czSSA030Dh3Q9WDxNCBBpqxKhjVc
Hy7imwdEoQKcqNdJh+IxAk7Cq5en+2E0+ToUi/2hHDegHFzXVl8On2YZ99wNqgRO
GwGYA5YvR4znfgLkp3WvpRzm+gP+6duSXaIpM2jlX0oTDj81yo7CFphmmutoxT06
Kn2AwJyjXLcxOcBIv+IVInGUQDU2LkaXK3/2s/hO2C2lBpbGL8CHB39zjYtfhbVr
tNvra5jZPtjutURcM5INP9ja7C4ytM8dHcypVjwA6Pw7rNGyygZB4TIMlShS/ccC
pIR4YMlisMprSNWffYGOyfoulNOO9ZZNuMB2VUvyNwFpbaToFbslt3BHKvf45T9P
gi7oqclbb9sNtm8jooZCPNQWffDilXDjfy+3sVXeV3Z3choJgK06mt24R8TynRyV
NsAtnxi7bDiqukEfeWLiqmUJ6diNE45G0eBFb2gS2HoSAERWtCOsosz3QE+jufNu
advVujYRsDuV0BpN0kdrawiXKM+4oeci86wQx93HTiOUikq+GIs+vN+3Vrw5FLjf
U5SXwF+kVJ4z5O6CX4hcD5nnLbHmxfZoiT45Z51s2FxFwJjjhCzpI82BRvOMcfiS
JCXe6NTzIltzYVpYiAQrpCZ2c3u69Vl8vjnoRL0IBFS024KadCZ420auwymW+vqk
JWUMnZR7qFnz9EctyTcx9L/TyWSp813xCr5T4U0nsEo8vr4UaVgP10Du7kDt8Ekz
mdktHhMhyUdKjRmpkSRbZIqJ+7hPG2U3cV0A6AYCUUZlq4dMWlMIl0/7T2Tx5Rqz
y+gqHYPvBcaRVt2gHaemTUE2JvyMVJUp2+ULyJUs9NO9bxbkJC61RM6/sQSrUiss
CeEiJSeSoUiMERhMl6FEfKEQV1+WKd3fJnpAChe3Mjg5/X5wk+ixqY0ortUgHOtF
ktaBVdiwOEnjwa3IAGiH5TwFQfBVBgeOuIvkGIjT3DunULgZ+1EnWsLnv3i53hYZ
YXX8zzpykDtHUBOHxvuTvjJ5ByH7sIlRKo5JWt6oZp/mSdQIL9aok/UjZnJPxA9H
p/LH5y3AUguV8o2AyqBTuuM3ZIPDdtpmpgVq7lvBOPDslsXyyfn9SClOACksJPU2
Rn4mdXNZghNdyexwNInt4wE+8oGcIq1+v/BaRiYiQkqg7VYc7l6drMuf/xSKg0er
BOLnU9LixERDX90JH6OYMiPVKxQPNnNZ12lMPN8+N7Aq39OLmr+m3Tc/3sZcJsHW
fK98RoI7TLswaLvizSKSXAmmi9X3DUhvp3LVXFUnjmvM/4YZ0Q51+ZDYkWr/dviB
upnaGTZXK1PAKaxbUHpT/yrc26e7fgSxeyPqkxXOTIGsOCD9eRoEu1Cu37AQ0KjD
irdkUULEHjR0/9wJqW5p+3ghtev67G3tw1BM5ephPt6GUvEF64Oz5f4GulwfVuWt
Hkbx5rPYTa1giP8myIGlKQ4d4F9BFB+r9Fr1gYmR7dRj52Y2qodmiBEIlgraZt95
2UV6Jsnuu0ok5cH22/eFvRxSriqqIHkEPXTc9//zanObT0I2wBRAsbVyIWLs/h5N
QJ4wVIqXV7jFvZa+IBJhg796OQT02txmrvt81BpM6MHvd0wrZ+ZAtW5fSC+Aa9by
i/cvRsrwG8551smCcMIxs732ffyDUiMLepCP/ypjBn9zyYR9cXxH8sCec2QDzAs/
NMdqzjydYywxbf3bgY6vb0kWhm8dc2/L/hXa9pTF2/yn8Dw/fbOJsPn5MqfoCYAq
Hl0e6pxaRH85wK8RzglKGHzVLlwdlWCZPgJ8btRo1y89O1mLNM1i8dnXrBLpGZ+h
hF+6J3axXBW5AhV4YFwmzR/0Iqi6XbcLcYBd+7/vROXNFzrngYjAeJJhSyxyFF1/
v65HzTIBmERp+PTjTOvAawZd7kQhaPkGFf8QvD2gaWLswAWHaFX/xsnPuk6qVBgW
47j5dstVOWNufYR4UcNw0VIEFlkBMUjJWvyCpZoDVddmK/oQ5/Bi5kA5qMdWE4Sl
o2eAqjHRMg9ZWKlrz8pslswXaUe+2P3kDjdQ521hbW4KELhikVqCMbAP8Bi4SJl2
zaMR40zXhcxI0AepYmcdc0eAYpvhiIrRNw9VrKDvDbnVLojxImfgXA0v4aeha+Jp
tY/MIYxPI3TDrNddSJNqBoiPsTORTOY+twfoyeQtEJhkRQyJSIJi3mtF1qLpSXkY
2IQEKUQx8zobSxOMTbS387wbxv416hso1kshK5C5Hm5QDYf+qipPxrjBkpdTPuN5
N4syvt2u4r7CJkCzbRI5OHp3LXW4R8zilATPcNp9plGilp1eUbcvi5UkFrcGY437
d3rfgmvtockogdT3JL5CTskJ9zmXCuS4+S25S75NQqQKDgcVKwBZ/PM2OfhOfoES
MLTqFhckL+JQsm9STsTHIJ735mDrKRvUhkhZg9U2kh2CprXWL5NveUTI0yKx2I18
KA49JuHSwpmkYG5jbbsx67wfJNR9lKPaHCNim/V6ws1B3rnDp39wW8mL/HxINOBl
4wkqXTrkRqXqyhRwCc/I6S/grs/2SUso2lR8sgItiJhe7zW/gHVhU1FALjmk5iZM
yinKcXuqLSPraT1Q5wUgtD+QFR2Wf85MzpYGiHSfM0xiFR/MvIsFAJDlGthAUG3I
tNpLSygedWIjvPlfEULI2tjFSz+1033rKQRfzdOIu2ceZweFtz6c/prnIwJ1Upnk
Tpi3L3XYGhtSiu1e8XmanyRrcGZ22lMMC8MZuOwqQ3aZEcPYgwdfejgPq9Nb9hG9
d+T6du/eNpMYZgKr6pst2O7YSdL4BmiSS8HQvUaRn7vDpNdgY5qB1pb3lzFWgPbs
Y3jqbFXlZqW+hP54g/fAEjOloJ9j7fVA8wO/yBXi4KQ8Ct09ZeBDlgE/s1KDlWas
PHUPzWWXIADs2Q02W1ywrGsNTFUOhr9Qu31IjE0Y7ciwON9qpudNRPa9R7qcrjsP
ydLhl1tWl57iP+L5relP9pVfcwxyAq8wP8GbP4T5/na5Eq41k35McLVsnlDJigHT
oJ3XnwDslbHfc5bE67f/4JShBSETOyVm6Hd4F9VKVqvD4dVSZK63F8GHk/bGXseK
IBeeZeW+FcHnsUkLiykrwtxEHvWWV5pC7MQeKhk0pX0NN+ymSlzFE0RAUzUmXni3
cyIbRoKzMcbBh4Av5UIc8SkypdO9AfFiXlZsxPFjSUgs5CgVESw8+O6jb5Hjl/6Y
ACHK31yFTIj4vX2wTmuolWcIJkTn4Gge0hNBFb8z0tHaEXIeHcud+gcNW9IUtgTK
vVh5FVxMEt2mc5ZneuUd+wMPWYRH0IiildZnIBDWurYdY2pB70K92qJGzVLT/KUe
SEAz+am4hm7/h1JbNzRI1j7Yg48opCMV/4ET8cCy2C1P3q0Xk5FLWPKltDBh8iN4
8+B0MkSQdOFrdoXylqhBZDET4Y1TLECybrqLrU13iMaE/Q0PHkZnCEh+GIMTqGq2
p/Mmw/3Q3I5kvul4otdqeRwFH6eDX9OizSb4kWN/It24uH/ktMVl7uyUhf8bwp6i
bXhtA+g8j7ZxoDTZRnrXs9d86U4WYaZGx0HcnR83aO9aSgsy+5+TUz2luUTg3wDm
oTn2yRK+HsVBt8CTLWwRE/XKE4V2IR3f3uQelq/GaTEt9woj/vGOjzZ8srP4nJEn
9j8lCl+mmWQt8ljKOegjDHeLinDOMwddWN3cO+d0rOfrHlGBMQBsZi0OWFebPohv
OaihaJKDYHrE0lokb7r+9VBOtjnBWd++lqpIvB49bxPxMQ7FtC+QW9XR0m7lWrOX
oSVDNj7rx81oYGhXh+4gwR08m/yijRaOc5NHvFM0VwKkhF8COA/zXOIeclFORUgY
Ctyp6PLps2wyR/Gt7hFdK7vnhh/ZMZOacf8Fp2PClle+kHAucdXk2nvvp6GnQCSs
y5LKfqYOQgfTb/IhOt7GPYBkE9BjgYNkoTo5+HCa+NUgwTXunPSvhaA6+siNM9o9
+4eVKTMZyuH4/F/GXgm9qJSW5bmbOlGUN6c4yZBojBDmPIDTdVhH1Pqpve0hAx3c
BySKn2T7Q0be4OQ8ZIo8rPNJP5Tn+UTTsFoGUYxwtYtaPKnPnZ9Ayuxedb72pVkH
KsUvWcO65Zw++ObwZn1iLlSaVKKDEjaxgHvR6QE8Q0ldBj+4K3kmcjJfGcny8HF/
LmpxpGZc8YDfI7bA9guEEGIYoxUK7gXm4gy6diryqwX0VW5ykPtLX4x204dWgrvu
yH2owKdSaB03uuFTMW0AEA6tU1OCDxuK/Z1p3VAEGoVCjo7rtMF7BS9WsnBYhf2P
P7RaywS0Ihj2Hbv6XCTjZT0s7S00YDIKudEgxaiMgz0y9BXMqjnvE16JuXDzJqIv
tnEIgDf2+ACt4O3Lzv2bIUHw/+TglB1iO5YnTiYJEPz0/+mLxgrpSKABrndO+WoM
Pr5u4qNBxzzdA4P446pQ9wgfkqa7v8rNT1RZEskJupsF/ZA3spAUGG6n+jaxbds8
ezj+0iq2ijSCS3XfZxLVinSSTicVn/kxGLJ48uL7sK2F4bp0MoGyjZwvNvq1uxEy
dqnfVa9c2ZUixUpIiw+wmBRT1q2vWQN+vVZrQ/FN1ryI3rGnMxFwJYei2J7mQhNh
s9MlQjE8Z+GCHu+ZjSEfzIWOmmnkjASSx4cwi4Ire7QgwWgM1ok2qZlQKo6+SSuZ
my0h1pU6qRCMUYS4FRfqoLj+YHgrcWESnC2PDc45tNsy5Q+R2R2N0zr0Ekhl+1Ct
XBArdhmY0tBY83/6wz6026rgr+EImkJtShwrQo4Oi/+3x9/Tohmo9LDEiyKcI+x8
x6/rf09a5xkIEsTQ+jM8LWhkd41vSW/TIGfkckPxlQOIhKWZ5q8H+iNeQ0qupj76
IjXYqfuoAfNMytgxOiKNmOvowRp6suprJwpOe7mzfB/Rv8QkLWxTpMX+XsUf6Qd9
Mg9yCWFrHyZocObgV3vQ/9SbyMOFrxqhdgyKCIyBRkphNSwBXIeX65jnytrRa76b
gw6lrQN7E3d9Eaj1aFNfVIS7pNqOOBX7L/nFeoNyJkpPNurLst7Z3qV5LEsjHOQg
Qbg9QEu5Yh0QL75IlImliVkMohEHRpHINLHJxt5hx0t0a8sWHubjnrpT05sAEPVv
Q9OejUN0PGuxt0tWDiwJ1lT7YX+w5vu18whVV9vri0/ewjeBB+hEdnaDv45/N4zC
EhBzIytXMj78bhiraeLS4JqqIm2OpR7U0Wxn5x0JmGS2FJMdsmXuDBqP0RhYrsJ3
JrCtv8YchQ2lEJGtw38hQi4zbpdEgrNQfenJNnim25jzRh/zZBPSyBlDEJjWcRZJ
Ve+pE6sgaYz9DQdXpKrsIUf9w7o7YAqqYR69EKXgBrLXd3PmmONp3QE82xrr91Lq
fXXgOvV7Qh0IQB+PX9PH4dbtpLqKPPoNvAZWrsf/CClY3e6MiCjUsZFjPF5Xuug/
nJQMRMT2VRP+TJPZJC7C/PDq2n9AdMvgs6FueAQZKSKgDhO/wnc274zmrWv4Bvz0
IeZWQ8/Iy7BmUVyLCR8Q39qT+c1Z903ibJtkMEwBSgBwg3vdQK9PY4s6qgF6JPZf
AkopxZtXQfWg/8XHOhmdiWGUvxL5py72LS2MasFKDFWvyurCS91QnRxT/02HOO2O
zhqsYktOlEGRy+mWFTppUJ3yAHly/bVxU6f2DAUt7fz4K7Q+n+mN0Pf1fsKkND7Y
h/OVJ+7ScbowteWdFsQzJhvI5jWeUn5HuiiPD97hzrISZ7nG9MRe/mS/Ot0of2tB
KZ+nbp9+nLU20PwvbJGG/1N3fE2zmTYBNic0ZdGcY/4ueK1DBEvgP6FKvAhq9bmk
LITN/6mMGvRiT6jkUacPkLJ5mWXoYRTNiOzd37KIjo+Th6PM3l0n3WgaNnNSPWu2
48APvaxfqmXtrv7evd8Rg1IezX0x6pPz+QBFMbqqcfrZRjTRxcmTH/OkBcnOPXuu
XBWhH1oTadePHoONnGQn7oYvzAH2yTEXCoEPWWLp8N796Ry5QIcfqVcc3VVMjFif
TVdCKtpsTO/ILdrd/SnFB3MamWH2JdqHBe4UOwC81hxAkzEShoV83lfkGIgSltnP
oeT3+j6kyDcvvCXFsLN8pLHD7HFasRy/YTFG7qsYNyDfq/TJfmUyBFooqLBBOwGR
s16R1hxYRTaPp/ostWC+5LkE9CbBXUN81ntASu4PH3z5q/060p05LIvVLkn/brfL
tCBHgUgZorbwrgeCBXzbs2uViiUF3/b4DP/hjb1eMfDcZWDROCoVGgZHt5QSmNnr
iASc8tnn6UMwfA5K1adPsOBgbsDHvQ0f6Ej+0focIoNtP83rq8RnlXIATnG6s3No
HXdWDX698rvhofng0deWGVNy1RdtiGnt8b2aHmdqBCRWtbkok/eUI7i/N1SE12T5
ShzuA9ojlzPFnWNmr8yD2dNadHenvDuPypUEyCsFdHaD0PADP3x9mIoSOrMRfxCg
dLob8grcEs33K7DPMbVGqzRNjmtgVJvriDUvtZRobLFYcdgrbLABCzpCOtxkS0gS
VonZaB7ZGnz0tp83o6kQ5s9hGVbNTLVE7CRfX98JhJa6zF37OXQrPrDGcpoLa1oy
I/XvC5FlvVg+1IJqSB9NIyeTzD3MBxjZ9X4iTVAz+nQB4WpnWK95gQc+ljNhNz2Z
DvLyEhI5cpaUUx8dh61BUJCxCrKvaT5M+knuJsvzFr9TO9EJwlvghCZejw5ef2D+
fXFccnorVK9jQL0lo/6p3aq1PHPqz8dkh2gnJ4hpLdnmOx4VbgpUU1gkMp05G1PF
lxyjjPB0Nr8Zl9r0WNjP6J0Aa1hMEn0ce/X2m9ofsCJ+ltlIvuCb0OSdbqVjfX0R
AXgMdIMGl15eSgPdNkobQo1WEjmc9cioR+95do4B/ak+Axvu7dvl2gGaatKNIU1V
TlH01dDLK1P03zysAciXGv4IXtMDfp0pabcMN9M2h20919Pe4g8KSgFcqzwSoB/e
uK1mIPp9XR3ETYJSAfVUTg4qoBlOWTrR9EjI7lNpM1LZSrx15OkCZKgJ0q5dWLqE
J+KcZSQDKc1/vrrK8d5IUQijED0/Lvu/x69QUqTRR91pEK/GHCMexR1r6xNUmi+L
qzfyVe/yOH6jv7eDAKQiXzryEmdSmxN4DlPGscCv8SPpDkLbxgQeYiQk799MJPU9
GIyAuGaY8cals4XhqGvQ3el7ujY7lWy3PfBomVEG/YWkZVKJku65goVBmXtyiJwO
/VlcsjgXwJMFVA3H/t07I2VzLcZE0oowbiDaxUXcAv1SP7l+goYc0suiry7y4ZlC
R7wVmuiyrhoyBD//yMWsD2kBnJNz6kJvQFNg/YgXpYRtdZ3j3YozW3uOe4cj1cNa
imfub/HMP84lQSS6nzaBHS9MnxJz/nVMJck5ReH9fPVBFdwqMkL2+/VAcwKHsuqv
VeILeE6apNwXE4jE6cf6hELcuq+H5NBzFUEQmt9rHlUHDbLvh6pA3xw0vzDX0Tbe
gR/5HzGBN7QYQCmknxhjupkZM0F0svgxEiSWkGQvWAvNSpTgXykLB6nFq376LF9y
SiNYLNKVCtbgfsgJkqHpHmHrGmCQVi3vsUGr7HdRq9ohOhVu2+Lwjs06ukWYsBxj
2lg35biVKwAJl+JFN1UW47F8+MtJJzMISUV6yjYTviGLxUf0yLIA6CP8zJlN9ihI
ZB9O7ySt18k1yVcQtkeo6SIgPFUgRtRAryHOTBTPAjgSL5uHiMPdgvzMRhVTI29f
T6EX1yym/aRzkE128rJO7LWZt9L3YUSajUOoLq7PkLXlaro82vjZZ6d1+x9FgRqi
HFwV5NzW3ae/LFeu9h6mpBaQuVSdDMc9V/AGzA6lweq/XogiotyqajJrJpvusw1I
DGbxittr6GqGriNkxK9mwUh1BGvHWLZ7acodLbHGS53fnHI/rUjS8fsVBBGn7rEe
m/y3yjDuHZw+ZjMRcgo1m/WP9nI+5N+FwetgPcPTLe5oAaHYhYoL/PkBIC6JqsEz
nbP5pLMZPvXbvl022/kPezJaiZCCsFh/UEufqAEog9IuojSPx4ezL754rWEQk6WX
4kw8tNK9dV+Ey4oNWa7vCA5LkuqTZUtL/ZSSTa9YMN9iCj5A68cbuB/uwvEHkKzU
hRlyuSDTRQ26xvou5zZ97WqR6yqf4uAJrlFPRF/42L4RIQYcJiR4sAJu+wIrLkFb
etKojsY5KwE/Onk2B4G/D0huZg7Lb+brpPDZSdOyXVILvyKfdrfmutisnB3Zx29K
3uCZa6VeXdc3i1R8uews1A0pBbHsI//9wOAddlGmZrrB7mrDdhwOp7lMdErAR7E8
4Fa5Q0DEZ9TVMXo9SOSRjc/s+pqY+hzbnajw3Q8ouanywEC4DRd8J8K5Eda0zHeq
Oih084u3lQ2TNoeCY4kMDjHnaLUppzaUXrqpC9ADFA5Tg1f/qlGTfYY63BVSZrMT
LYcZBHU6wW2vB7Q7fKUOVEWP7By8WvEgNJezM848IyFiV4ogcU6LVFKlYiWHrZwi
nzsc42xsv0Q6TbeLBbaDS4tgUkKvXGZImbV4ykJftgz9i3FDbGipCXkibvyufVnV
oUFCOfH/SSZeDVq1BiV1W8w7vCAyTAmHBWOjOpjtzxYs3ZKjbUZtamU+zQPkLjK3
TTj18zZ7NlnbELplYn4T6MK42f+RKBknd20s+N6VFCuipBOIECwjT5p5b8TEaAZ0
ruiVkILDJh3n1MPrO2DWXyglOZGwLBDUo5Ew1T2OoL3BJJxZmbVR/TvDU6zuyBQL
Gib54FzM17oPsikqAbcXa1Ps/PTHEkvU1HzMY2Ks+a+sGEYIvu8fTN46K24TcKfL
Rnhdi7rHn3hfRYPIzApMSs3zXDONcixtxF74A/YVT/8A7fgr9n6susBzL/d7U1h5
ASvw/LA6MrMkIl8TwlcOcesk9B7/G8v/rXqo2WuUZbde1HvYu9A0q1BtPioFeiwp
Zl0pF0jJSJC6Ctu3RXZbg79cY99D18i9kR8a0ZghnXyrpuGgT6xVTXxpk05OK/es
svGuU5j11tDrh/w8tbQS+5/jq3ksMHUVgtoq/sKTfMMTGGdWp9nIdKg1z3yAOIKT
h72rxD50Y0JhWXPz8U+bML6Z4L0F3415IoHpyLzFprrvDlmqABQTWopeAaFzi0fO
snzyKm1ekG6jqhRGNe/5QpJBd+zXwhS3OodxuUW9dXUlnJvgVKnGvxLP7fLrFd/u
4tUQNDkIrfml24Ln5x66+E1G9MjTAaRAT8WF4o0LyaY+QuJcFw1BB0UeCH2pJCLG
SOo+7uRNGgIGigC9p2fFy0vFP+AW+RPlGNv6XNOo1Tp3qA4wtJKc2ShntNYrX3vq
nuHSEZf/3N0QUOgMGZpjM9uDMSTkwHGYgTZHRiYnkWdFroEKApdA+b+n6qnxRGGk
bx3+DorTcGdZ20UUzHNjtvKVNE3eHn1UtteWXqGi6tZvUvecY32bB18Q6APGmFZZ
7cX5Gw2z62zUQxzvKa1Ui9ZCY8ISfl9pkAVPglr6HOCWA1p6C80h9R597bj/MSOF
sv1SWIJ73HtkK0ehNR8xjPn0VzyT5dSJzfxNN2DqGRtclyQP8PhRBt8CBdMaAouV
xIQSv1gftRUOUsXv0X4wbCcsX6dnUAEQxQ4/2uGpj6GA/tkM9RCx49i9g+DGxiIB
Xc1cb9b8NErDeWqK0wZMyKt7CZRIq4Yb0DPpegYawHdi2Ros0/+77IckWd5bBGMt
L2xshznk/KLxr2yh+l1N+4W0Ha/G/3DB9LRAk4saQ+jQnS5zhZXbo6qUcDEaUGPP
ibyHqxw1Rs2VOC9NqTn57ZWtWDhOmLefgcI4SCD1048Dj6ZaoMY0Pyok7FJ4Twwy
5ZPyQWUPqPM+UubaMgsdCT1UtBCi7k8jPyjVGBfXFbhC2Jm8F1/JH7Qs0LQh0dXb
sr/e9pk6HSO7WbnU/28D6z6fucZrwJyVdjrJx6kHmfK96YrpOKEkLIjXpNRJb25P
hVzIx9+SL4XIVicDyTyArbJ6rldGuQNFEI3//u/MxvP0rtNkDdR37AuBnmRAd4pv
BCy2Cw8p4XpGisQHMUZE2AeJV5TKuacW1bAKwgffaXkVMrfk5kFccs6MpW89Wqqv
Zl/C5t4+7SKmGiy0jnfEIOYx880KfNrY7ZZ3P8N8hh2fF//B2etSVuoayKr31njQ
H9iYAVKjJWdBhWbgkmXq6pxVDKS2oK+SXdI6qDA6IBgak6cnOx1wexBGz4wxYCj2
e+YkVPitYWP4vTs7lvyAIH5yHNbz5/gDG61pJIIlfm4/iUpO+0WVKj6SxoFopniU
tG762Wod2FZnOgp0FKU3dwqxQtyhrOo1bKDTQWziZCSKzncFkA+CHQeJZuaoe3iH
S7kzJ0fkUxwHAvnQFwZleil2PjICn6y1CW/ElobVtJx4glc8oy/lHFJrkpp1IEKA
Gg2aWCr9SiQ86Ox0EYkuWnR8eF6NsK8l0Ga+haPGhqfP1jy1KXJeLXbQjLyibioT
MwoDTnEdLtILFkGmxSyaT0YKoqevzVMZuq1QN32sGzSNHyVsW4xKglw7K2mD1OQ0
oiQeIsW/wnGgaVt1rukmyIYJAXvgnUlmMdfbWOvyy7DBDSRkUlKST/2wqEUrTLMC
42L9ACnlor+PQsSQx90qseY4TSpYmE9ZlsVxdr1kvS/AmGRBFhKnoeL4spP3/0Xd
yvSlU0d/rm/A0z8RR6L6Yk6qo3adLAaEze6VtJwRE+qwakTRubzhFR0PgqfMzcoH
DjpYAv1KN7cyXht0qfx08VxoCyA8bvWFTMPnkYrmfhUzFDvEqefrjU3n1YdaRuiq
L3NaZ85dDzIE/Y2qcCWjC2N2SNR1kkceCwh/qFmgieBP8YOxTJZxHe461GrbZL3r
9pHXWLaDKk66eJ+VxfxzAGq5o73nhJ17cezYSOwnzJ83OsyjoeuIdqiHci4d5DwH
s29aCcIUvEsuUCJLowq+1JeNNx/GCsa5lt+hdrUVIy8VrNKO1iJ0dorfWziy/0SP
WRo8HF+RSjjHGxELnpmtWz/jKcoCcVKUqpY7W4mB8ttrnddq/u6qJiUTd3PPlpzX
IxItWdMMUyuyc9Qh+PM1zBJsknoFhH+Tzgwb5OovK5KcxT5u2WwajqPS0I5lCchk
XJcmeRICElLc/u5qX6k2pA9tS/MvZpr4YMQXXoqMrKAFTlSrheOFJhzdT0lnzKgv
CjkL4PX62Hv3j5zO27bGk65K87t7hxdVE8PU1uyXUplRL35piKwovUgk2RsvaSSM
p1Ro+pC/nOKigViS7RrKJbusaLVN0cCQmCqRsljg6mR16NmW+IbSVAGW+PQ1Ir2R
qRfIsV2N5izWCwUO5QIeQqAf8GfNgyg76LaJFJ/DPMKDc37pYN+kkhIOp6ViFiDI
JsKI//WBVI/G1bfaN/Q9sYHrR4kqFUFGRllQMABlbOHddvl6KTs/WRSw8PEtvdtq
wCKQbBCahzCMiprfPpu3llaAv/yxk3Soiq83UqhukjgmiIY1IQvzY4Mt7l38HMC9
wx6QXBTHrVP2ud4b/iew8TX1fmAdlzPOjy0OlncmQCeo31Cs7N127yCgpxiB39eg
q0ON+Us/AREUZ/QNjn+HNvIa6B6K9jtIXwB8uM5FuKI7v4JegKiL3KW5kkC31Nt/
G+yC+gska/4ctDMbGJq3BrCv5/qZx9ZoOvAu4BGxuEGRLl3OSe1JZbNbd6BEtjH8
kR4Uci77RxIPV5XzVdofHef/ojRvpZs8OK05VFtiW9PGGf/xJDDQGDO0rNQvJztQ
1Y8/j8eelW/MR9DGq2EGnnW30y8xQ5qz2jpEieldCR8Kle8nCZY7cIklA2iwuh2X
cTl9NktlM30NehZYyZBPyqRdCdErtr4w0QG2VqhJT+5L1XvAsteOtfqtaDJaxXST
2A5FwZf2/pLsBO+ccaX6pZyznwhfmDQG7BvHqPDwCcCe6ftZDNl7nu2G54lwhHi2
ncwWo9AmdqUH8rRQB6ILrtnhRaW4fuPVodE2yssKGt7CKcnvvzoDfiujucPjs9OX
+H8z/7djIGTN3fDvgobvnqREQ/qWiPuIvCb9gaUnTHidTpl9MNe/ei3uKptlHkhY
CsM/vZlnrtwUcQP2wzhHz2+CzOQ18xSt/TJZgnYR9kXHi8BEkJh/ArTyjy2m8E0D
xuEctFynpDfY1A3GXON5A2j31+hdvK2/t2Y1HJeA1+hsqTbnuEEVuBNEQhOmNxBU
MgZeMh0whIWhm+SBKAMi9O97tx4Cv0zZfoPBhPs/hBzQepnAW70bFlAz4pLgPhzc
cYvXstAwGwRK+7qCOthnqiv5ibr2kDkSj3U82W43s1kysL2uR5xF52fSWIl8TQPS
HzvsjqqZ3mFJVJzsC3FI+e4sMI8vG/9XcbHDBdIKk5/VtFRMgyd4uvhY6ARqhOKD
Ij7HBtVJZ9nQwBDWP/l5mDjnz8o/1hjEN4I5We/a7CHJ0+ehxlG4OOx136x7BAaP
wLIGWtUM7raTpq+RUAijQCjSGGRHvmi+2w+zBIoUncss7fsVak+ALkgPaRiQTkI+
mJKyTtJmAK2ZlcPPiHzCSHTXZHZxWZ1gt1sKa+l7apLyD7YuVAOT+ea7xOnDDCFV
l0jxsDhMxRbdmX0Qhg87Rm1gapGbqFUcKOQPTadvF/PgGCqANktkEp1PuSpo+wbl
UtDfJ9vzuufLu0S5g6SRXtBg+WHWke6Q8Hv6sQ5pJNjeVqsv7m05XrILJBXRuAVj
5I+RtoXpNQp3l2yHsl2JYt/Hxz10lyPZlqTceamyPn3Q6Q6C9MpR4zzyWIm/+sUR
Z6kvdhIoK2nkfkKXRMaKVqOeMC4H2RxaqW2Z508YaIcgfs00Nbe44ZzBl5aFhRKZ
ljRskLe+uNuaKLMZCpSJdbqChdAt8BS2ATXQNI2BRS6pZUIqO2xt2XzpDkwo4nn0
5tkUyTA1kmBFc9UCRugZDgzltCTwqWQcyrFhXys4LeI3aIRaSGw4Ft9wRqw2mD41
52EOfI11JquFMEmw8tzwUvdre2TMSl2lCbLv1J4fo05JfnitVNgX8S8mxpoQfv6V
DomTs8ORzvQkr9UmQVtzZnw6SfIis+woUR0NloKhyCqzZSQhmH0CVpaBpxnhSPy9
50MZ8cQhQYJjjaycVQ9LIfb8ccanASP+ubkTsc5VylBxqr7buv94tROC8rXsvEWZ
Mn/j5OUdjxldY4zShneCzBxO8go6ddSEKS8jkGtuMvT7B5jiKMBxiEAryzVKJj7g
nUwaRpvS4jUWHkiFRj5DDnfy+9hkU7g6MjGR8A4BZdHCbMKpKDtCJQUdwnx6LiT2
JDYK0SlIph5pH9n9YG/ToddqYTinMb8q4JC32iHlVH190yMvZwCQqVV4YhOy3cyQ
mOS7bWOsK6Xfc+/b6NpcY/HVsVA/z7k/0Kgs0RtW/T4MxLKB17aedWbXywYa7kjq
MHM1biZAREadTinVrcaE/qpK0NV9BZv8bbkmr/NUnLTkizFjndZc+ztuMFXqh3Kn
0eS/epi/G2lJHVXwtXx1q73CSbFNQxC46clJmGul3c0gFcMetxi6sXhIg1NvSxFt
KilAn4N4lIOy5Lml5qn1fKu4I/gWCquZd2TM0ITlt02w5gzZrhDJMNPOJlS4Zkd3
MQznyIjOXbt5HArJfTPF6YUNElBvYJxETeKRrL2iVK1rYysckoeXDluONzWq4B8b
+gg4zeAdnQv8h7gRH+LzODuk8hIEVitPA/f50ar8w8p8PMwf7JhdFPqzwsCeBqbu
Isvs/ksA/gZWdiEs8FTVTN3aL52JcpAoqjpRH3Rftlmz+NppvHoYzG9WUK3uqXPP
nqTQAkSNqiJhoTSmtDceCqn2S6vBc8npr4UBKQLGEJAxOgOI/wUaVo2/7XO9eVRO
s1YIP0FiV8kXGmz3nm3iafAesQeuFgKI9gSxtHsz1lsWioCRUnPXy2he2a/2fc7c
QFBUgvoePtkGz0tGWIy2JzaGpzaKy0RRWzCISlQ8P34m1ntuiPKnOSn6kow6Juod
I5sMMKMgoCBqbLHy3cIJle9uSsjbQofeAInWPWIUs+WvBJO3myVTVePp719W57L/
Ck6SB2Gg+mSZG/j9MZMM4SCoxyxE/HJE5Ta0ERvbTlxIHOhK0vicXBXAT1pcbN9g
MFBmsZwcJrQWz8dWx1sGg/tl96FT5eAZ6VbK9PF/AzWKMN4gSvpn/i4oRjyjD8mP
p6KDIivuY6EyL/OyRebbWnf8YHz1qjR2wMjwC/VhDbavX6JSqIiJQkQcglrahcqZ
ULYkpE+cDIWjIGMYpWwqUxRwFgzrvyw224F6jklaZWm2j2MUm7bvp75xkkka6OPr
uBayuOmlbYtRGx+CuZLVdV9diNzGMGJY9IkFb8K4WSwFhFXD7xCxmPskhRdzIONS
Yw5yeC7oPvFEnlAn7m279w+aYdqwZ5sLHwtXn2yIR1JJTT0KE89CYGL+z6B19ON3
gWJA/B3Le/1suMg9g19RAlD2na3pLKn+slLqgnfMNzqrCY2aAKaKZY4PX0JOlvEp
ovqfpyNoJVl+hKKaqZhedwJ5+j6LYdhZ/R7Iu0vvsyRcjPRkpbpGoYIggaR33JAv
e0ogrz9Zmh7U5O/2Ta/8F4IPWLT9tfyrEK2aj44CPOQHRFlp4yiSDYemGUvvteU/
tGnCWMjVmDPDfrqrn8a4md13+z7yG90hd3rC7oGxRfQo/wIEYwTdoNUrxIAAfrX4
mwCUF8P8ddyYrwgpy9k8dcXpkQmFYxw5mIkOh8Gr2tRRURu7vkaLhm51QEuQoX00
FWo2a50e0r8tXETBRDGv5vib6QK9iVoSbRQVRXzFnqAFmpi6rpN95lE2OV68AHiR
ZtbtGqx6ShkZQuqoJBgteu8PCB/nhVSR0g2ejtEo7d1D2LGqmMtNISIOd/3tq666
M3aMcJGywcStPgxmsAcp5Uqo7izwptSR1rd/fwasoACEepu3kI5BB/pjlHqSNNpN
H7UiWhmzj3hT/9Va/tVpllP5OSFFRb0U8loiGhR9IkAij1SQTC3s6G3I3+OA1Rww
6w1rj8wBCfQtY5abY0OAZQEbLVOHlDQzFmg+EiZhxgOygCTq/Eg8u1U3GMV5T1+c
qOTMFHPnME1abCb8rBkEkbXy5w3Ax/6H5im6IIBY593HWsEwh02yaVFhWwkiECFc
xNHL3GQviIE6qhKHqAgLIAA5XEm0uokA50SRWv0WkcSUgQgsA9TeG1+UO2OOEc1H
kqY8XhUahGj4Um0twySYVfNkdNpOU2eaTrshjqFe/HQ5rRi64dhnyLHIyqOHavrF
Ucwb+dQcuk1zr007BRr9LlFd6vzLjVgPppqSUQrpR/xTyQuSOUP1fv7d8anq5vnU
T6ZvH97lfft8WmZnv5aY3cMBGFNYDtIzVg0sxAbZRh+JfEv672OW/l3NYFHLAYom
UZlPs90fMomUUFJLdbHsnMWHWV/0CjfWVceW//p17dTSEwh+ynTyGOiQ2LpoOguV
LG4o3pWwTETGopgVdsPrzLLI7zD4Ykp9eHCnbuQVD0vgYBFzHAU26UF6cnVwhBlJ
P1ZSglPtKlqBCY0fSCk0M6ITEMC3I2qg+j7u+v7SnY2SmyFPLpaTsD4+F4fOUYH4
bV5bGBeWbMw9bLwzRCEDR8uTy9AT8p/hTof1ttD9KJOt4YjcTJJpPaIPXs6kEj6o
ghz1hzBoSRVsJshqPwF+Zo4clzkkjBaKR0TCd92olvT/+5BrJZx1evGzJ52tqBct
Vm1jFHIVXAlsxy43gFfpDmHtzQ3oZzasRTR6EhAHEdmYruFu0PEMBrU9Wq6pio81
ESMznRgq1xbcOLgZZTOxkneA9Pyd3xEypEMZNEb4MBcbtKFFDvf0FcKyyhHD4x+9
dm+APNb1NvkwzMeeJigE56vzDTSYYb79uSdIAIulZ/9f2w9u/h4Gdk7tydqt8Ewp
zu25EczgM6UqXDVWY6aXDU9gHhclnTiqHn9EIpT8ayv3NXB+Qm4maoxGkgeXeq4u
RkpMSm1k80KI9fhyAJh7092eglxCZXrrNeuTCnA7GofXxKN3mB7FP+b/gy+G+Hhh
T5sSpVuzGwzzu+1GJqAxwq7oPn7/lnMl1q0aoAV2LDxJlQe8HBzcR7M5dvNH3QO7
papUKL5FrXkGqv6QdjyAW0WOLjblvuiZzu6ISkYOQ8asZVtCmZYMVo5cqpGrnz7G
V5jADp6dSsIZqgOXZRPeCPNaLQMHlOu9pHYlfSamBPdbaLVToyEX1vUu3EE7RWKF
EegRDu8K5kqK8Rqp33SK0xfciHt77fUXOEykwvEGMNSJMG8yeUIRO3BaCdPTxjaa
e5RR+f5Mgm1wEaph1TN67nR/WE9b0utpHiqfJ+LE6j5mLEFjxdNn8A6m2ANQ6wTM
z6Jscl/FuNAi7JVZQTwlBa+R9s+K8HB0xIlJ73H7iXTJRD24XCFEywklRKaunTCU
FuIBGf9gFzmKtqD2vABm4ARaL/n0mepLW1VISkhOnbnm9dWbxEZj24e7JrAp7oGH
S2dih2XazDffE0wCbbA8JuXnWixvi7oU9ZI8rkmVk3uIk99n/eTcrr7wTJRXrkOu
DqcVjdb+RVkff13eWXFUGiJ7ecdvRlD+E8TMQg5Zh6QKtKzOXsSkl9X62v3T0K7S
K9+tpP0Xf/Xwuh17ibSfntUjSdNZ8m7Wy7hbV9U6JjolthLSEMarXU4FrzpD6AWk
HZLhi1hxXO8t/1otnTUdrbwXKLUruasbCe/ORQlBnThzc+bLhHPQKsfEGKhzq2xl
+eGIFtlnSfo1fNI2MdS0T0Dh9X5M536WikQJ/weHP0q6wjH8z2sEmgmpS2RKA/4c
+L4U+RJ0CNbpUtVZBKvqXBufOWTQO164ErSdekUNYiHAY90nOYlswycWvJ9CZ3xZ
amNVck5W301gLCUh7Vn45ArG6bKFQaSK/ddLX/wSeGwK3frEmhB6/225Far88qib
xDSCIa30XI31Fqaj+7FYuQfWP7RVkvckETarQs4PsOjANFSbezZhtbJEWCGvcE0h
JGzFLskZFcsr2TfVPRzeqhh9ZTyFGpuZ1ZvQcg/YOrP0yGPKkUy4ZXS9URRa2Oge
spmOBhRYjRCVUUiErczWHymgan3HjpMqxMiINFTyVdbJ262K/GUn7Yh72zCP3NsG
kkSdWjbQpwt7Q5FEMJAK6jwQ68Huolj0qt6x6ZBmSV8+xwLgFkuTY1ziVh8VGeK+
MZPR/CqhdHlWf1AaH1JG8YWIxO/lNOoZ2nsM2LxBNzFmPrZ/ihe2Bkz4WxFFKjzj
MK16QRwFvOzaCMIREtcfGsOrkVL7QM29fGSzECA2H56UT1gZauE/VHARhS85EvP4
bkLw1nxImOEjhlq9fcJQWrIINupB4fnCYm9DQ7lPfc7vn4lUp53/2bS4utlICJHc
3z9RTtZL0bCUYkidF7fb5HKWL2V2uBW6g8iaxQijHjc4ThjmcEyXY4UgGc9w/oxK
/4eajjhftkxNsWW+9nyNA3Ulfx9VBZPNOFHUZNsLFw8uV6lTgwGwG0mVZtqGolvo
osGfmJsCR/nRr8cnJTD5N0HufqX0yA6IMyq5YEus8yiRM6Bt6ADrVV7tLZrI20km
ZRLOVE25kklSEIlrWdNRg4yGF3x6oYjsJu1MIKF7lA1tLl8vAeB8DOGxjPKAYu7T
NNHHkfp/1wFYB3um4UbdItws4oNM3jxGPMngruzGrlLcKNd/5HO8Y8hxhs+CggIK
/JJg5hyf4SKcljvjyvBITYnJsgylBiOANEjoODcBiyRvCLlDWtLKyshkoBZVbGJH
IXG7lN7jAyrYrgxInQv7UqO42OmbTtaqK3FxzdzS3E478iG0bnp+5Ghb0bYUA0pN
Wt4oiZHNwYYfiaTRGRRfxlxH71jI0Bqw/h0BcSv8O4iWga5YHPsNRtdvsH8ue8nw
vUv4ZORWmj37d6LJt7/y4VHNWtGyIdRNscaBEEFY1VJmkqNZUPqIUOIFdIUtm44w
sX1CKdmrqWyoSIwiwkEZpK/vF7S2FM3vAuYwX54LfTsQ49DhFNZcPQGcI2UnUue8
vwmZCkI/EtG5oNfs8IZvWk19uLQWG+bhxPOxBBU2Vh6meAOCIGj1dP/984mSJdhk
0xLZMCfeN5X+3hhz4/HD5voGcF25VWtyc5gKrBCynQ7ebfuPldjPMOsr85YcU1Jr
E+RkJGhnAvEzHHzM8D3li+y1clpcjWOQR9v6f3rX647DVh48MsRgaprkZ2w4K7rL
aYUzcjCaGeWxmv7/lEe9RE2Qqa2pfTILOkIK2TKtySlHhH/jp0qLeqMXN5MubgOF
MHqLPxbO5nXlcp1hXBfZtUPK4rFpzCb8k/qox+u0q9LbyaaxVyKfGOFxVt0VLX2F
zXs6mlCv0nHfvYGaJLlEiEaD0utlskxI/pdAIksI0N+Cds0kQEbro8wr9WYbF+fF
TNqU0faLpE5UTroQyRTTiAGq++Rc6J17yzEZv8nPoCGESDBUsjoxfT8VkPaFanmo
JVEwEunpAJ+9sxCgFWvpu9ft2ZmnJvQGcntOR4xZvoyq/q8wvFw5qN0Ke8q9Loom
iy8QH5t8wo/r9FZYxg43Q18dM2tnqVdA3znGdGPYgoZRKAlaah0rEyFHR3gae+sU
CdFa0OwU+6d2hehUqfOLoxaFViVC6lBgwPwztwuFYagx/491XJ095qOBts/E+jIJ
Bn2jG5zDJpB23cTVVyd+xjCGxznWHfxRkn/BZeg4I+073bHI/dDAL9NwPuAd+N4a
J76jLbKUG/0c/13H4Bs7rPhML5n4lNJZabRsrzpt5xQDQEcTpC5YHxYMP5k4QiHD
905m+PEHusEuSO/Bb72ahkL9w2L7+igxIl+Dm2FWfo6g8vg3nR0D07tWeHcUXsHR
u7amDcWB2e56ZzchjEzP/QWjt3bJ6yMGdvQvRijcZz+wTj++bX/9AkQuR4kcLs+C
Jk8ng/ks3CCwjwawGevV97xvmlEZPZCtOq+QrtM4s6djrkDtpJFfSPgCcK5dm56E
o8Verb4xlsQ0QoaRgoykUebM/K2bitXXxGjQEcLu3r9BLSmAqdYztUmjvO0bT259
AFdD6u2WZVois2D7COWM9bNTXulzlnKq2UJbHnb+bBK3e0+QtvGH668UMkyg6wwc
CgcnApGCkjMdliTIkV0S2sE+zVx0eNwjCuN7HlN7kKe2pAIUBwoL/Fr9jfXj55v9
efn8zJL10Zllf8mze1iACia2preU2v3jS+trt67bL9WuByu881aes1RDBDE4J7eq
n32CHNMZmiNb9f29JhxtdvqbMmyUFzwzT74c//1DYCA0+W52h5rBmHZOM/e2GBgW
8Lbudr3GirFLtMYgdNt8u7ugcPhIRcVIVaAbSdh8xm//SiMo/7dNEgbUb0AFAH5L
PxqtOVD5kqQDSG64glnDrEfC5tVrHKi9ru1rONVxeiD6ovpkSa6ID3tqYEOBkB6w
hUabyFsaXsBGkfFTGAqkmMYii0aWSJh9JneRGh7Ldvj+sY1pApSAjld8OVeKEBPt
OVw8H0RXex6HSZLnkBuwq4hFbThtglDXuvXwHkVCmMEVunoUqWqV5wTuwLrWk/8Y
hn30BqgdulB/SqFDwjh8e++4uhu1DwOeB/TTMooJUgi7l3gB6H/dz8pcN89NYVo1
pPtVbUM6DeXNKt39DodEtgcvCyy6N03Fn+NJ3W6eTechCrfqeJOTWWTEePQR317L
FGVw4hrXy2DzyT8YDlzIzE/VMiedFr+bBl+oMi7sOeCrmobYN/Md3SrTeHFWjnr/
mE44IRGW+UENp0S07EXrA/npOhT85cNdgg/QGvpTUNldP5zFZveoAVL4eNTpArgZ
JSLPbes6mWBeBoisqkNTpnJtTLVaB9Ju+XfDRLD0aWIwDskba6znVUjiarDrt53U
y9bYrrE+vFwbQquC228He9t/bIsbD/RZ9Z/nJo6lO4Cx9YKhTiX6W7H5o6fW1Czf
JMCqgQVIFNx4kqlpmU4t3yWgecpgYDSM0KoBhvzRI1En7OJrbqex9OCkF9pj+Ca0
sgQgt05aOrodA7FAHfCO6R9EDEu2ms4fzwzsVJ9j0QYg4YX3CKyZlZMBXXsxNu48
+L/ehnbzuzP7HXIOxXwRsyfOoz3VnLupbgzfWnSPmyoPml/b2g0bqusbtUHkcVY5
CnJmwXmPccLhBphLNrr8yZtuvVn6Uba2464aOAa/WAK6A3ig27ij/ZtVDKv2ckNx
4SAwU6RV1uBa5ceZnWdl1DSEPCroHaESn9A2FiPQqM/f/MAX1Xlqvs6loWWdRcNv
7dUEWA2ne23adoCP3uhkWMu/LXCBt6aOw252Kte8VQztukXck1X+pKCx5GRIEwJQ
0BVX9+VFdskp+UFr9F4YnaGsuYYrYG4WgbtfhyFobd/0pUDfvSFESpzxQ/A+2Iz2
JjqtUfIFCJaTTe35mVOyBevSJFMnueobCgvr64wjPxyjBsCvqEHZCk4OMZv3jpgS
1MimLkiJ+J2Uot9jLjGx+XliVOKh8//lPLWb1JxYzD6klQ+gYIW/eHjW+As1Q/aN
lTO6HREdu9HBuUXgbgMGzhUgGRjJDbU3sgO7pDaqlj++7PnLioFGcZc/wDtNd/kg
3tFp+MGostMTKPeVu2slS8gY/izKGEYdHrQ9aLWynw4qsi1iwyW5H3sG002tWLzZ
tvRrLx4ydxwzMNoW1V53EpYHnmIz6plJVA3dbH5eu9YAG51USsNQCCDDsVAhpuGx
V+0xROvfkibu2K2KRLx1E7Gt8bL5op0nd0ZB6xi05B+2rXdRSFwV75IP54c1RE1j
1FcJwRKJjFc2i2yg6RGPMDyI702jMS3A94PfMyVxgJDb9P2D78Ttb/vjvE8nXf/k
ox7HhnI0HxQWLqz4RTN9Isol1BzSMEf5pd7YhkYPVBOv+YMxVgXrNIITLA+C/sU2
Kr30ppU6n8cLdYSrX5x0H/chPYnUdhPhSewJJk4J0pNEd3hAQ4nOZjot3bWRJ+jx
HKf0ZEMBQUaIk74KZLlpY5QpNbpEtguKGli1RcfORyyGZc9Bzwv58bedVidNofVW
m+xxy4FirBzzq6ZGLh0/fcIApd6cUI0FSVr9MAsKY6njbDm5yV96NE7Hps3Wb8cK
Bl+ZtgFaUJA/XGwuSVDs4sRiRVp854EgI5SmWYNZxuNu7Bfn/tIfdweOn1Wk2r5L
rLjhtUBYFeQ9BjE38IAVGgTc3mFjIp2qEQ2zckekaEzhqt2billW06+cYWdA/hL9
QKIdZqSXFtNm1n/lwYbWbZHLp7z0IpIiBrx3X9+1FXq1gjPkG/7Px52LJZRAhOuZ
a+qXIz6oxjyrmya6QWdfyqQqWFp+A7DMESHErSkzDUR6DRPnLkdhf3Lp+sxAlnxK
EXQi4luhnKgHQkR9oL+ObSYwGQQmb4r5vDHIdVYF2DcZpXQP3gQJmBLzyupAGy+A
678Rj5Uz0FzbNMpIhzwB7owXM/iofcQXh2a1xR8fd4HMYWT2Kp/PtneL9Ccqodtv
ZKU7FSv76CnUwG+UyqZdxg8sOOdQyi25+MboPQUB/0mDUYHCi+XF944HQPPDao7m
d0q3XvSfpMS/sD6aqnFjMH2p6HQpMwm1CI8rWEbi3HvyxnpEXwRqofzZjOdr0MRy
wY5NYJ8ssYb2de1ic3QORRSx/hTCS/lHfc1gzJrLgRrLoIJSY/VDZ2N4AKLcYWOF
gfeXyntVxqvOyjyC70aByw1m0U7R1zhHVf+wUhveFV79UA5h+b+0KM5osqfs6S8R
ZLcGr2/hcOhLFYjoTvkAYc7OoYEFf1KhYyx3x2fxb7IlCPcg3PjrTUe1EqOkVa6B
O24+DMZDObhNPC8EafIVwfAgbqFkf50v0JS7HCVhKd7Qnefi/8zeUQOtd+Wh2yMw
SxOGSDHFlVgyfyEvswq2LV1xYTQx8Vj8z7yMS6V2vNIa0Rj4Beuzr0sQX7HDCQyj
vt20SMhEVNW5qsLBAqDjfviL46SLkvZKYPnDA02T7oh8HoI0YWG4tIGK1nKZPwbt
6yko7ZmfwIccDzet4fo6tQ9Cb8txVuqOmovLZSslc1nwhWT34I/tFpUXV1DdBX2V
7Wvfdj4eCdYcBchAmKe+cYy9mvDQCbKQB2HZbWLdNEJWSPjHkFEe0iLNixrVPNOb
gDkq7eq1pWRNDAHJ9Nn+Eyt+ftn2POC/qUxAI9h2L+tEgbqIF2ukeZ2pnyx1RXK0
Evw+ouqnAd8BQxj4UZaV1e6BFn48VoYke8SsrS8kzJ9OuyazUxE9iipi3ag72lco
2oZaq1mOcmtQsIhn9gn6MaO/qjvG7348qv4r3jsub4ZJskTXvT2aRTlwQrxSOpNw
47f62fOoRxdxcefsvOy4WcBJaIqu0M1zmMYriR7ABrU4L83xsAsQkZu1ZAftTWLn
Kn6+GrZ6CqaaeI/0j3DhoBFn6vGcQ9Tt6GyPxxyOWH46HpzRJdasTrCQAqaq3nhs
iP2/bpaZQSRi8S71KSLAipRK91xHJ/fSLynGsR6UyLo3f5/8eU8GKDeTulihK+l7
lbBFMANYOFmJTJJEurWjUn00Jo1J/46W5nyM3RnN3nI/p6ViXNlKVrsMPSk8Hxzh
ns3CXqsVf8cr+gGSs9XXe6Tut3Um84lAIwoRAEkw2XwYwS9MmquraYonsfbOuIsH
k3E/eE75eeathnKIU/UYhXSrDduOvaJikr3cVlE66AUd+ukUxC9d8abxh2CqtQ7s
AggHclz1/1WrbAKwqQi3RZ/WCtX8gS5ti5+faPikexkV4Bh+E8soV1uswFtF1KmT
o/EO2Pyb4nW26E9ywB0KpfZzNeR9fj8542iX+wcQaxMGFmnmffYC76lMKD1MqK0e
BQ27QZl/Dms7ZLufFqcv3ARV0lALC6cfiWMNJnzFfwo0GiT3KpzR0ba79yeUDH9i
8K1Y2F/rbrfSIJc65l5eKyqLfPunuonjD58dN8ImCz8FbRd1w7DpvBlayoKwIiTF
7eomXI2bHJyvIvKGh0gpLJ7ShSm8Ot3DbeKrgK+8WuabJJXbNXhGyXqnPoGF6JBR
Cu4MO/zEwgZVh0wMrXV6XklTDMTdy6ZUUWM1Vug/0sjJyDoA+1mRGim/bIlkGV+X
CCuSBtPDNIDc9hRmI4tH7KguS4sEi5ycowGIYDQHT19SjqalIAxnXo8dipLi/TMH
5z23TtXvmmeefyrclhN++n03z1DwMDv6yIoHUip8ZX+36x6dFF4FcBg/Qv4OxkI8
odl8w3dfC/hFO2Xr0nUMToxQSvAqxDV+XpRhszLBfjKjV9PRohV88+fSt2cVopyB
xS/R5zktXG4LV0p8YcLtKqVeaq6ZaDVxa9T1nthTJtCKKEZaiBS+xjRYR0wG+KPY
4dSFRX/4AOzl8xFcGzr9xuVSp4MZPT9Y2KWdkuTrCTmuPnvgn7e3clOc/j9Wr9Mi
tKAsHJl38pTHiVCB4rwwFNjeR7hpqczza5AfmaWa1fW8G6YjOxI4UFqfzdfsZTD/
MWE7FAsaydynIiYNbzMcRsFBa/0TGXMmgLEAJppIrLkWbGWNcL7sfU7bfYxMEjEd
BU7qoQvbC0ey9MX/oqX2DmpWDC0EXvIX0cCFO0oKHXv5pfK3yiMucnzDKJ9p1MKo
j4bcidTWeB7QQU49cvyi8eZxCZitw09pLBRh2OtAMWc0fnm33iSIc3V0EdiejKEh
I4RMlV4KLukvbmgy7qYbGl+j7/bAuykG9nqtyJ7XN66qwKcfyYO2ig/bcCqLLjr/
9jy+0c77GKLDGGWnHz0q5oXgJ00F/EgTNtsicM2jckE3UALNCCJk8Dtc53NYgEk7
OAuMP3mTJCq4ZB1Gqe4yZJFrTwMvb2byNUfdY0dLs/H2oRo3w/A/bhSIcbJ3N6db
069XvLDz4tUV++/g4x3J7zT2BURivn5VeqZsJuSvUBn6uzPQhiBkDZbPqcGEeYxx
QYUqHmiuj1aHGSSwQOo/xRbbskTKsCNId2ZZ6gzJucNDG0a8W/gS0w3FfNqAEpsu
G8c4mUv858Jkcm3kIdMKMyZSDjCM0E0h0Rn9bHPeqr5eiyExMlWzU66Wdgmta28e
MY88R4QCom7WBt3XUCJagkh3Z+6opYS6joKUpeR72cZohCpNLXtjdDHiB5Bea7gy
o/Ngmn/Y+98eNLRb64Ch+V2xovBXq/HyWPuF+AoZ3cx0WDwIJQmeUwJ2OBcZeeG2
dlBeDosGF5AXFdrjRO0FSPjqUfevWQvBrCkVEzMBJJTq57QvxViZuhd0W9c+EDzR
vz332NDZvPpG5XUDVXMK6KdmSsBE59jI3FK1tySyEwUao2Sn8eWFHLwOZH+OcN23
Z7ldL2uXL8uzYR0jkVea2TIgzJ5p44X/XOzmmEjnMGWWAuS0oJcE+ZTXRu/Z4Sps
T+DytbshubyDSXYCCi5oMgggKSSqUaLuPLlnC6MNjGcTQMhokOWZKzKq0aWOAJFU
y0QUYVKwScVTTLG9Zyq1N54SPZIZKRejCAezFy9xeBv1D8/cH5z7PNeOxYDskSxJ
nodTYulxV0p3Dd7j3oaqulIZEgDNqVQdyZAtHwuc4DdrFU3/Vqk/jer//brxT/yH
q1WYLk4osKKPSDxm/nxrfGcG47tTqa+uk8FIwSQTKNcu/y4973/93krcx1pj2H3y
jBLAtaqoLmGsL7gj3uajLo1POhgcigC9msbTh37lQJhklTgPU6pR+mkEdqdGxAqH
JW6LxadWS09BGtguHMuHk1N36cnaISO/73JIU8FKKXDtdsqTeMjvc2LmVHE4UvNd
VoTyMz+QU3TRnoAgUgVzkLvTZcXv7b+ZbhJrsTPPQ8zkn2/VZqR0wcwj4TQNuoJK
n7LsTXeXC8MCDxg1yq3LT6owifzK9dxp7Hw3AqLp3eQt6oF1WD1+o8VZAmpMMtV0
YgmMp52PHLYo7RQXxGQZUXLQ/uiuxFIyCqhiBTHfxwtNQIDifTAWmOlwT6YayJAt
LVLY3q5NewDeAITAzWWDIjRl6YqzPPUR0nx6fSg8MeS3sCwDEgoZ3lNtsjO20MSg
SA0VUdksnDSIGvqz7+f5DaEY8SY0a0nnfqlg8OHLSwlpXZzRARrfixQaDA0w8349
v0nUj7o0uemeGQSYDGalaGyp+Xqt1Jx+Bd1p1fR8nban0Y4MRdMVqIwbMb+oqw8E
3RAyb/CTtU3Qii1qDHEPhVVmvUcRLDqoZd+gdtQjnbCWM7c4t7eEH0F6rXuDV+/R
osS+siCr+vmlLwmttJHocEE1Yt/sS1bOQytYsGEeF4LY8SyCbuaP1RqsyqM9OHZT
rz6FLKBCXrm8T4xWq3jBi6VsHhgcxGhePB/ox8ekQZVIvjkA5y+DBVnsFuxMAyrq
NzOq7iRWNqcCvnWyDMKuEV+LfJL7zTL0PilXl3T/Ag+NgxWk+VYYmkA94BYWEESY
ilo3Red62OBaEOXHIHLYGfjmENKZBJqeABacF8WLljZD8S66rKTGHAngbIzbI4fk
ZML1EWVddikdJ5LND5xte3ILk/U/8Lo7Kg+HN7w76OPe9EiIni1enq5v4agBjzAO
XAHb+qayPGRHbE5hkT+2hgD/IWWY62ycAVUdXQ1YmveX+T/wAo0efnQ1Ma+LmKZX
NmuMlGnd5sBeDebvP8w3rn3RhCbJHCnP4ureH0+WdGEjTCRb+hzVAj10qA8lyHbB
PnKOs1rLkNGMchycGbsge+TlrwOqMXQNGeQlMmuQvmvq1uhjd0PzQ/PjXbQAOdiE
bOuuc35KCOymCKowDLjfh84Z6+sZW5CVy1bv/LSEIj94xtPX+S08fsZf1pelnVv9
x8LugqScFF8/+jWijef1mSoxMt1mABVTZcakY+5Rw8HN3erJZ30JaLRtCHFvc8MN
UfWa7xdJcA7/dEZ3FudPDPAV4kLyK+n9+IxWPYGuUQTJRAOed+6V3oOVARoRCO9p
5evJNmK43RK1qXsIN4dVsECinnVVS2juXk69EQv+CMLB8k1pfuHOR293HRJhVepA
RA24RCAaZgsmfGIPwIukxmaCwqO9bbW0XRHQcZ+Ft6ActHCwz8zCJoOwBXTqDJAK
y2xhR2T3AsMdhPJRNYqbwXJPa8q65BSJObFD6ySrDnM8tGDODgWdCcH10Ryw2xHC
PYeZGYSAMITQhh07zjEg6K9/4EHminJ8uc49D/vBZqYlj3wbxmy7z+PEswU7ga6Q
KvGNR/1Ew2iHUxY6RvGVshQ2rU8ZpfbOqxSEVDMq/lo188pipmGNIa4ifv8d04iq
YXd0RLyzu7+DfVb287TvVgpbJy7McMImFj4BK9kKF3BK97BGmvlOJoOGVnk3SYe4
kDzv7fDqxCitgTpAFNYUw1v2x387r/g8UF8glnYKFMiTecuDX/+xy0rMuWjNUjTN
384kANP8xsIMqGiqP7GY3naPe3iwxZ6Xw6g/pg0b34BUDla9LWo8373v5tcpUf3z
4RCOvj2cSTYfLkQjVOgCuVCDLvK4oeGwLEa/4bjibVFK8PJzoJJguQwogzNMi/I/
SSqv5lAlQjP3rYgeOAwzjBXEQVsATAGJDpBN58GlVZAwRpYunMtKfZL5tn5oEHKf
zyzZcAwEwCGxySUmj6V5AdpiQstNoULU6Vt6Upo9nA4U6riswkLvn81dfKxE684m
xUlzj0M9BZ4vw9TwpzCkIKJQGniteCBpkaaAunGWXUE56A44vJJ84tN8s3WSTvb+
k03GU8knVD2s3HvvwBjAXJKN/Sv+3NpTGUg3B9/49HOQ2+PP4wLr6JRm8NrMHnOS
Mgiurp8yQi+7R0S+9CSNp6GSTPSgkwZfmRnnV2c/1wRuLCug/CE4BS85q3vfTJri
QgQGuPm+4t3Jw/e+MpwtH0b93TLhy4GnBcFLiDlr7DkBNa29h9Mf6r2x3RN2yHiY
IX0dB5FoTurO+DeLPWDrlot8SOV2chTxGYOHyE7eSM4uf9GoGB+hQ4H9gB91TfbS
xfQ3ed7nTArCvbHjpOqGqVrpqZ6FLIun818tg3OhXs2/9Eexu0AFG1v69eLQzzWT
EV/WL+Nv+PU/wsJQlUT2znkmd9oU2vzjPfMRqLmQqlC4nrCg+FwVUtWXtot2GdfK
ADNTg+U2vhhkWuu3CLRffi0mHo2chyVxZSL2vbUX9ri1xwGpDTPoNZOIf1RFlKYi
tbVtrODiGvjnT6ehi9/zDpMqkJJEwpDCZlVuDPWMLFiDXHscHZY9IHKShMKv37IK
kW1NvXQGCM/ZXWsBS0jROh+K3SrQdodrnTchKFx3USlYNU8v3CLwbIljQmzrvfBX
qYtSF6apzRkfJlCOPFUiOlH5L0TaJ4T4i7+gQvwwb42WeFSE9br4yRFLMcGo3bPF
yyKfI+PyOaBFQ1fKJLWwzjFKaVGMXydZMIVAS3W9XT5JZgABQwMHeqJcPrExgn42
CR3gf3V5KzjSmF+KfWSpa7OF+iQ52MRw41nN92mhUZJNKCBsPEuXjkOk59AH4Lfs
QOrc4YGcl/+wHaiizDskFCm237R/V0KcRCDC1zcxcT4nnoWoOobC7dk3VRm2+vxT
ypEhi9HkqXDBOhsCDNJ/vB5YR1NcGdKdCFanIkBSx9GDutOYBMURhsxbcfI9lo+m
q6paCPj5AIzz5z07dnZzSA94KbwSXw9M/FKDBtTqvpdzDScKOQFG+dvnSk7JyQLR
8Wo5bhVJFed0s7lyoXK5EgLigFbwZdG/7dacMdTVC69XD0SXiymsHbvsGdKVJ8if
t2GNTKJHTxltTj+N4t86Q5vUTsIIp+vpT6EvvjF2kjVReJUK3XatCBsejYrnh2gb
ZUmawDzPMba0U52PmhSWCcBHZVCncic6Cnkh+kBzbam0cpYvBJuJ+auWIpjaICCY
5U0LkFx4RQh5/l9Qh3+1zE8qKj9KbS9xHX9BSHpZ4RY0FU0J6XCdFsF4MApO40L3
q5zDVjJLMOCvqe278HdFhWsxekPd2CmUVWXkb6Mo2gs/JPEUeeCJ4OirMeSF488J
S2RdKXy6mUiNiYIQORT/GNpYkKvqtZQtrMuCGJh4AKGRuc/Hk8L9ZsXL/Govoo/L
v7yXDwHzSfkvaHweZ64Dh7M+T1DBO6bhtLZjcTENmDg0yQUAyhSxOZErz5z7AYD3
lbszTl2eDGoT6tBPMR7LMUAtvmta6krexvdi8CBQudhVSThqflO9P5ilkmuHfu2q
6SKZMn1xYWW9sGf10qNyQBd1ny0MEwBFmP+JUQrc52qkkHs0tyEB2JVkVUkxavK+
3ElpZ/WmAk+uSHR2Z09URscGAbzr8UMz/hUK9wT6vwvWMO6rT+piQ5d9UVU/yLw1
kx9bnFkU5Puliu1KDFjje4ankl6SGm1irYn/1QhqUDPh2m4CDritG6HIrvgbGDxw
6V0XbDQCPdQjT0xqGvK+9um9Uej5WC/uf336Z2wnx7gN7mpYH8wClV5Eh3RPpvU5
ipya2VaWCehrMs/2uX2JKpzjgpHy4VRZWTNL5jcqPRKjZtLfegXKAUg3XBqGgk4j
cPqFz11GNWign5NtD9x0dcV0RGJwRy2h1XVZ/DOlWnhvtTUJYLc/xmpf6qRIWxdD
1QQwO81kUejs/W1tYPyNbbMODYzHSb5ds1g5Ok89wz2d+HXdfXUPkrOxzJ7sVCSc
T+N+R7G9tUG9DdQEp+WNOL7kH7VG6C8h8FaePea+7QEwGETqGXpCw5iCPs1vcwgW
M35rpHUi9bw5HtZwENt6yW7KOL1HnBM1ymTQw8RairfB9LhQUBkngpoeJ0hBQIdT
XrjVDUzy0QKTkB32cXQD9byBaFpRi33jLst9ny/xaRp/smVEeGThld+KIvrnaZBb
Oo7blQUfwd561h5DMEL6ohsZ5QfVIO59rCnw3lThryjviokM5hS2AA+/wAe18T6/
29cTC27eLKdjqcfNyN0qDFkWzDnODBnnGzX+yZOeXAV+xm0GI9Uisji2ZxtfKT69
E7icTUYkb0KEZ4hFyLaKlVuDPbWFbQ9khqkPqtrj9KVu+r72oGqHIkKpG2GVZqPt
29t3Gn8lCG1Afr+7TQzlqPFk2VJrqRdvtO5ZhwjHzEtp2HH9udDMUw6397mAERGo
x//j+DFv+ZfTomBmVHgkSRuCbQ27z3D91SXyPULnDWxWbJATFJzIU1U5aEOtby7F
a8RczM1evhOKuUFZoIxeNxA90dPRkYGuG3tsvni3QJ15D4BhBeZsjcJfLSO/x8Bc
DRVKmVF3qEyqNE2AZX1eFnXVVOyRSgR8HsoA2r+FyukQL83TXCJ3ZnkyNNKiNbdv
E53wcf4jhlkr6py5twZmV2CKUsIb1XMX+1XXvlKknZaccMrLNEcyNHwmkOn9rCQ0
sf9nHvc+L9Nxw2kjGjjRNGQyubAovi36TsBW2V10TYaHnnOpFbXsdww1A127QBpr
liNTMwKsZGFPCQ2gndnlhWiiTXDtdWTbF1VUUXVvejnbALGc5GdmbCOO9ErGcHL/
YdlSBFjcc88ETgjqbzian6GkwCE0tzukmo7Po7Rk5o3CxV59aZ58mo7XF1JFfvWs
A+dntJBJhIUS71gPW/+fHSHZALWzUUTrwYC+/kEgjgSs09db43mbaLLLMqN++pD9
rMkLp6Y/DI+G5eOvOGUBZGdvOMv+as91WvCMU9evo4nr6xM7LsjOxaaAmDnEWjqR
uM9DDfElIaTdlq82tc26H4ZNw9rvX5ULjR2yxOq4oU4QxHH7IyIk2oV6hHcwGF/g
K2lW1+/P11wWtKi4AJn6A25qlOiTwXxC4vVD1lVYnuE6YHJS/ti4NXKZcwuRHVhu
CdPXyXXc+Yg14FB5eYAPHnNr+BwRA4eR2kVBTC13s7y8TGGC0QeUpoTvbHoqULxJ
nI2TyfTLLvBhMJOLyP5EsU3WG1naausIhajLrem3ZNuu7D/ykT8N55kcIPTjrigq
+jAH2q884ieETPt9o3Fts0yJUcz12clSM+hV5sqlQLJZI7erjrWxalS3GKGHwNB3
Yp5EtZVtodLG+wNyKC5rBiwtnd+h/j2zJQww+luo3jqJ1IKq+N1BFK3lBuI44BNC
3gDxL8RKRBILHemas8LnZlf4+zcSvvAJvMD3SKLwTKEg33FhZnr2SBPn7ThKIdRO
b643Zyd1SSKsxrc8RVKUJvV/IoVwfJasS4/wJY/Tut6uuQQuuQfnVWoIIRwzGGMc
74Bfmp1gNpRRZG86mnvrjhAOOMSN8uNsdBmU+7zFgikwPbfRsZqImX9lPT4HDTur
WhI0HGEJEtPuJsBnc6Zpbq+Eec1ncndTccAEJzX6JqQ4skXCKgxVSl0i7+nuGcK8
xLPWwTwhoaE39IRaAafGhYwNCFZ7ALIxx94V4a2l6nJCPhUiqpiMLY0RuUnRhmBl
IyA5EwE6IunGHOojgYRx4NbIuQ2l+jRPXrUCpQ95XYniR3cVSY//7RxzEqxvwt/C
LkV1L6nTdpX0yMbToYfzLW+V5eI5ZbJDzt9UoYY31IqPwNUgcNuwmS3TCui6XTT+
Y5bg2Bq2/baaGStlcUZtNGgGtaxwZy7mZmfvEdgFvR4+4Dq46wyTajdwRdN1viOS
RPbXNIjdqf2ou2H9iYUh8jcrtPwHWlqY2OWhdpNPa9J9Cr6rRrV6lJU/1eGZ53/y
VEnYxbAUvFI8T5oXHDxOk7gO1cNWMAi2spzkjBOOjP3hJFJKgE8MAztW+AUZM2YC
8ijePwN7SCtYiAF834SZ8xJ5wgSQHdBcKJ0OOZOGvIWnrKu5xf2eOOe3bATji3Sh
VyeC+XiLWs3/lLBXPn2TaGMlX3h/JljNoWLcFFWHQEb12F6FCyPTMQrBFQPVRCpt
HDDlOY911XHr47pIIScCxQIdTmeZAd4KGVrRz+VgbsfYvpNRvv1H7RwXi0VdhlAu
m0CwwbXky9FNzbzuq/yxRk0UwBba79AF2+UcMPbPuT7yjaQU2AOWV6TLCnbVnQn/
ltOiM9qptxqa50lMZopAeXaO+1TqE6cIDYE0o7CXgYoO/e6H99CPFNvmBR/ovQpX
zvHnFOqZv3G7fCKpMPVDK44lHwHu+YEq9EkOXtd5Nuohx3cegebLb7JRp51qq0W8
GfoXJuvEH34tqX0DV+NsSRtUBbHWbS7S7ikfWMjF5l+DCvA6C9hiBQpMJKCO+Htr
l0wmA4zt6PektORmz45kX+OU0QlzBGZaORhbSbAuxBJn2K9Df535VMDBgBmlcBF8
ilhlhdG2lbkqsNX1L+HvL/7C4eUI2TGioaHXRV4gBQH2EXyw4RhB3hzuMZwPuZMT
rUSOySak9b4kaoO3jTz9Scq1+yn2eeX+7Et5rI/JKO34do8/mh76dC0Cl7zTbDNl
uJgOMpdP4TjVK7egEPckRtMmbv3henhZqxALy3mI6gI7QqlTF3HveE7Mq4n9MLFq
CUG2H8c1MVqko3aOsCUH0v/r2s1KeRKMgrMUpgZdsRwnc46y1/vr5QW8eIFf3phn
E2RNqTDEdvb6TiLgL5DC7615wFZQ3uv1remtw17BLXeMMspg4CpY+OdZ/XNqJsdp
Lp+5PX7j6ir5H0W+xf79SXapRyceKR4kWgRR8G6ZJih2M1WgV6Ewa90TiYY2IIhC
mK0Nq67uWjjueg1+d20ia8ftJUDSFU0n1fXRrNEwytbrt0Ryqa3ptxNIVzkUNyRY
ES5pe8zN+kzN5Heq6diJ2Ai/pYebp5cTbPuqqynjYTmdiLknZehZy/MmntIbU56n
4zVAJS9VROlsP/cwTCLqrpj3HEjUEFYaZHfQgdXmhmBs/8libtAPxLuQdeXsWvfb
Y+XMAXcg/uWDSSczepwusVJHT/CRFUWnWG7ObHkais9dlbRnxApojWiKz4rV3u11
8wJuV/S6g5mA78gv+bbYuCOo7GKs4kcc58tIUdL9KjHyiycv8nmj/OdTB1NvtjY9
ouwOvDD2N2QXjIiG6LL0cqP0iWnqOPHQERHJWrDXu+jrLb8IClnb2DGklZx1ijSE
e8QJq82d297YLrvcKuWtiMG+4ibZchDouNMfAYFRrOrw+Ow8yD0oZhB+S5A8aItx
fH8QPSJVrZrcRJ2VYAVOHL7ROlYpMu+0X8ezYG2EoF4whw0g9SyUW07Ov7jO6Scp
9v/gSBVwQGakdg30Gpp9DcCLfnGAGFP3GlHW2jSv2WXpRsCLSR2XqiHSjyz1pK0m
uS1p8851vqaIr+D5gEUghw0oQ8IWmBsrfHQie/82IKWFk0/RQAKGsmqYX9rZML4L
DkSokW97/5jehNVeICq8DtZw0L7GGZi51up4e/zc3X5IcZvm4PNmN1WDZY5jCsUc
WTvWBVhi61KXW0yTVG/lpowvo4LHvq/YtFslul1EauKF1Bfm3Ru8x7KbCpVmdowJ
C1u409Wg8vGgywDHLzVHiSD2LnyMcbIh/cpS4jYkpdo/GvAOAUucCNmM9GQqjWoL
lblM7hW8iRkIopmXs4nxbGoNeY2SivrcXX5gt1fYiGM2wG5dMaxqoOQDYAM5cMM1
d35qhjvOBYGzve54oXwISHb2evydMt1dYRl+VkdayWnpDXxgesOoCLRW9qTACS8w
mSQGMZf4BYPadMiEiKcl9URbv3buSq+Yj70djbO/+EahTZqspJtdWYIqdGmHOudz
DaWomFRQ+qwOidRfChZ+0e9ZfkHylK7/DE0S0w8HzLUZD2uNDhPw42ldceDGOc0S
ak0jK7TDaCMoqvULCsUz/LDpsLKsa00U6Tni21mIXL/r2UN0JHWNWgpkaqXnyk8A
AXEJXluYnt7TUxJwtZAnc9EGTG+MlHUS1qbTwPhflBMj1vnM/YZ2w2Ux7V0dKCnW
We/Vb/ofrpHeZBb3jmoDxp/5pLLyoZJ0vlDssC0MCpZ/d+jlunRfnAJXjCISY6Lu
PqCrCreHBbyXuN3x+3GXm3EOtNKHVDuAogYFH+nTNwRuHeBrxlJ7bpge9PBcDRy0
c9JAmfwyppzp2wZy9+hGlGndx5ArLNalAju2G5j0jXENRNDrLoW0RinjpOkKNtZX
xDOmB+Lq+/x8F7pUPwEo29DDtHNPFAwqiYQMkWq6XaPGTJV2S0vCe2atDCMSPtEj
iqkH+/Yui/GWeo6ZS1BnkAYZMw5ZKYTIg7hIgzI7oe9wwuCiortI0WKTIdMSHcYR
cQjkh7cXbGwmmf0xlC710/5JN6U6TB29vOEbrK12vtrfkh+lOT52KlXErf0PJ7kl
xMMSyIN8VoUCbxbXSLeXpLeQUsRaDJwcy7XRJVYKtaFbO1i7+qXJ1v+aVgKrKlZA
jL6akECk0YXgWM/yd4bRNlg2/SV/YaWVehiLzlnEXTYHfD/ksERw2FIwKLyUrrir
moEjnRr3IketLguTTMm9vTLpXNIJ6aMzX0fmVtDH0vRskinBdFaRG4x+rRsav1+O
xDIMFE3Jj/zItUUi2RSnAQ==
--pragma protect end_data_block
--pragma protect digest_block
WDCT4cWCAH7Apd+SJvP8+8JO1Ww=
--pragma protect end_digest_block
--pragma protect end_protected
