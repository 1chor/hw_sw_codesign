-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Xq2/HvL9spo9DaZpMFNwDos0io15+qto8Yd6Htfqo6saw1Z+70ELdlNV1yPoIBHa
YvLrUndlTTjFJpqTYD0Qd78Iwm3sHahp9FK5nBxhZrsrUqoxCUrvljmv3+JhpWIG
m3AnM6FIOoAZ7dl4oWYpqbBEcTwE2KlKNW0QFZknqOc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 29214)

`protect DATA_BLOCK
iwK3yzK8Xd4vAaWx8TukCfYf1DbpbybSlkx7QiikIrwZwT2zk4DrlAnMRL1UwO8r
kCpdga8cqw3Joaklxfoz9yrNSptrqMKN2yqyRrS/l6ltPd/4izJ0BFtKzkZDfSC5
3cNK7UUFD06nHJSuQhSVGoApbsWPF5H0K2ZIKgz/7IC9nMwrluE8Y1DQWVlz6WOR
DszaBO2L0z18H39hNLPsK3/gj0OnjgRtGmqBjwuyK4eivFq8bm3uCp/mE7PXPbxQ
aBfoMpzb0Kc4kRce7VcRkIn2TfKchtoXOjSOKDU6de7zOO3tKKJ8uYzGpdqs2Sje
v4eUjy8nsT4RsD11PNPbmxTvnWFxkPDGLVg1AGYEqjlbSk3rCVI2c5hZAvDdjYTa
Y1Td+XMzvXn/slDIxJgJFVh8K2prwM6uXe7/u5EIC/xWF6kXBnSZm1qcyrbLm9TT
/wn88AE0fEEohmdSwoYW5uxDwHWQVmyub8tNlZRz5zJ08uioCjNnzQCl9TpXjiGI
Q006584z7mzlls0dh5nlz3EGIf6sYRHaGlcNt4iKH+dgKPzBNi4NfCgB1Ak0nrEf
P+u4AS0bKfuEFFajDkY8B9BQslsBNt6ArZ3ZDsP/YH3UzaUOTeBtHxOgmCIHagEk
DQwyQm2PkuG4bKBJJD1TliPjoB/xoEG9TmVWSSS1YpfqBmZ4xHwRe3IN2a8gXQR5
bSpaWJY4543K5+DejsnWM44Mg8I4hbkhyCt5DVV/olni47s6zuvCmwIlpAol/o4M
PC1Eya8PMdMdyh1O8EJzOUo5Z+raexdDXF+m8DMusTJgr8qg9DiMNhsNasbpy9Pp
6FNaG5wtAaylTLgnWTfIDYV95zrOtqL1w4jBH++n1vrDo3fHLLvBmuf4PFVRvyIj
bnpxLV95ijdf58YJwb3n2F/XeHk+0pniWJpd+p7WEMQtyj2A+MRoyKQenqTQ5852
4GzcL+RHuR6Um5eB3PTQUPSczbrFWVzlnvIFlXzXEhutcp7pGoYq3KN8kNjk3LYI
ZYEL24PibzOjckAJ7zJQHcxgrLiyllofnRVziJ6NcoM6AELlQsHx0u4VVT5rfi+6
3WldZ1JmeKg8b7NTU9JVC8drc2ihWaawXyKkuTkYjbn8CwZwM8DRXDPPNGZslK46
4gBJaJVRrzehv2VUnOEE3Z5SovRlJl1thCpf2OntBENizKdNLvXdTjflGkzlorYw
6KkP3f/W5aDQkz23UpM1RYo6nIurpoEQvW6wWnWYLUn3ySFicXJByBhW8jEo1jCq
xcz1BsZy7nZJWQIo41hMTNjQnUw44KEL6hAcI/D8zvluDL0UmBNWN+kuVgKlhbpn
JK/+SYj9qAADqCjRUxAm9ariLqgh6UyOsq1HEA3+jhvh+dqv2akRvEnmLX1OhLxT
e4pK85ZLaWBfLkIrq2/+P50Fe9p8+7tKkIKg7X95Jh0sgIYmYI+QT0Us++m3bivv
8nGXYtiSEFHMGpFg2FcyXv3isHslyTpSQmdBWlBsVgtU1MbAFrBQfLFpG97aoLfw
4J9z31b6uOrxd7h+fBc1ic7nMnx88N6wVEekuqHbP4nS5wcPRNhNvcMdxCBwd+5k
CgO/r7Y1uhmdaKdfshh6BzwlzhjMyRfH97wakNiuZccs5U9Afrz0zuJ2ISOgieck
E4eW9y6+38RVkwVEf1fpGa3UjpF1MKpCT6MDo+q3JQg7xtMrlgo9m04Tcs7+Yu2h
oPUmVfamARKwZG6SGvNy2GxlgOVuvQcQtATZzlYsi82iI4q6Igc/p6yaAIGIdR+s
7nGWWVwJQcndG2ZM/dg/xKSaipTKr/Pd0zmOh0uAGFtwjCm97p7ZGObmDShTfgq5
O3Bnl7fBFkmyfHqhP5CEasyj5PcjfNlchx5pAhXRm9m77FS3cYjKWAF9VzN1gKj3
9iHG7OFdubiVF8jDLAAoPfd+tVIwl4PCHA66GmQtY8c/9SfAUs4BHHMfIlxdwmPq
ZjkeltQOIZzrH3EU43iQ+HY6nbsvyFbcE/Rrk3+kkSEwSPgoot3xD9dEJkjpRBDs
bfW8cO3n2vkbo6+l0eHzyqzo31tPJB8LNnaHcmN3yGEP1cQGxf1IoHaMY7PFD5Js
BEeAg3TUmj2YiKE5UMZQUQQaNLk0LoQxQO12eGbJOKWo7LzP4OWxjbh/lbARIxQQ
g21n0qAdUsLOOGotKMPvT9+gFWzVB0dN0HNngZ/NhmebfYUJpiGwFE0342PzDpGY
Hv38mMORALf9aiZ95LZh84MyrFJ20SLaROcEliyYMbMMXsFis9IwTiWGuSp6plNv
qyTQte73bIGvix3UePC9HfSNmrY92UWAOBw2AlQPhhWTmpHzwbVfjJRCI88tHCrW
mHaad3RpIu1Vcv5kt19JVdi6Lb70vvFThyInJJdq7M3H/buXVlL5tKn3rQs4S8tH
EMDzu+wwYBKrCFiTSWDGuavdQAi6kaFAdz6CenGVzphKI1O3fVyc5R9GL6DGulbl
ApoWfOPJEooS8BVqnKKNumdzjCKzsnakWT7ZP5dUY1oN/rNJuhEuuRHEHoDs/XJL
7Ae+sGaVQVkDmCo6nD0+EmbR9umVaCqPXve01JDR0/qgFsRSw7qkSX7HEqOCrg7p
Xb1eaBsbm2aUQMWjo4WcFmEjBuOBzXMeM6xAMjWU9Q+1LYjCMzgxdPXQMvyEoXwM
n5ONFFVyALcbKIjALPYg93P96qHEsTwDFMbHRYBdo7JAkkIBk6WCdXaYf7OJlFDk
i6UwLSLwNdDmEak/ZLjaoWyB5YYH78csi/Xqw+6CjG1Rc3uRqyusElHtNEw68J16
411DSVxLiULjrXWLOpewpM0VkLzos3Wq6MOuByUOQxhGdiKgeyDF3SpsDKO3Y3D2
pZzRzZ4fcUhdgwlr3mPTprRSkbfOd7olYVVSBLrWsomPWTc3vDn7olW6urUqMFwt
6M7l5EVFadE5FSYAgAXalxLNxBTxvH3IXVbKXDiRLc2f0JuD8isFTctmnzmXRuDJ
Nv5J4+j7Cf3abIHG0zvi/rcz+WRBA05bGKO4oOx8B9zfuOXvaVi2jnFirBlWOuo6
7ajTl7kWVJzWkw+NpLHTvAVVNsu8YSSKmavf5YvVrlHU9OsGjnqgLWCs2fjxj5dq
AqXXZIDdldH+xUHWmAt2YwCrIy0u/Dlp/+Hogoncwa+aw6AZL2taqbiarbf/zdbd
rLWA6UILBId4pDKu6qFC1MmL1OreqQFXkZOr6dBCOkWmiWQPlBMT4b3MCatZwO5J
PaQ+TLRPmCfoDbVTr3M4w2TeQs5zi/045RAFdpqLV5sWEVx+iPfHHc6r+RtQX+f7
zl17l4AmK2WZghZWowaB+Ne6qWfiRnI3I/YnTPXOXGAMFrnMsyBOmCOreJ1KdE+f
1/rHIQA5gIWeBoML8JBRGBss+YnzWVMe1bHCkfRAR1H1uEAB2JaNPA7DH0TNkxhB
sqhh2hgqmA7tT7BklAUZoLB1RFHJWmJeHi8YZ5t34IvN74UdPellnt3n2qTWhowb
/GwXaJNRFNKxuJTM8wM8n3F5mipOCpD7iIQG2y4C0oNo3EzXhPNIQnrvHPkUky9o
gpmIsSHDv6y4hGypyQPRFbEzRFbYBONBfAlsrkRZG9/3coIk2YZ1zwJS69OxkOnQ
7uNf3Y1Be+MvuAHa8mE7p93eW5BlLvAtjADiH8OnbGFlWdJHzt/ZPq66nTnI2I40
Nxhjsz3dWVmb/DRiDjQ/LsuQyuzBHhLPnP9YUEkDWqNJMUfTRvPPrHiM6QNx0d0h
mUv9Lr8HNdUEXBihDPlcw/5oI4+D4NNJ12fvckjkOGwyMofOT7QQZzqUms59k9eX
tW09wsCTTU/lET2Z2vwQ1tuE68a09h5pUr4df0UArGH1oW+oZoeWaZcxpxjfmCIl
nKCjQtHJCuLb4nn6OdxvmQKf/Cr4XfvWdiEMdIMOu5d1WQrtl7gEZtca4E+yvvOy
TtJlCGDiURdXJCWp3xTvhRcVMXqOA/B4+akc992dcFTOX7LdUOFwkGranH2NECNP
u7rbyZ+MqHVJJDzcBdMcn+WajguGIoUt7a0weh6Htvs/f6kQrHF33y3bPJsW212l
SMRsO4zir/m/umayPIdaGifAnStp9P3aKTUSdUtZ5FNz/wHo5swNF/f46cK6uQpJ
Qxnl7DMsYyzfPr9yg/BZNxopylrWpZWE1X+ew0EvtiNukAgN+Z1W8Zwy0A0MBbCB
2/EuhMegWC+IuQm5Xv15tmYLPNsBSgfXVn9B5nT7Opvpwe032GFkxmezNlLPrj/c
LT/z3TWRn+08UgX3ABy2qFJe3YkMYtvB1I0pkHow3Hje2QtsSzky0oO7kaSvX1QA
gAifD+torikbzLeNro9nX3cBc7gPZ4SeJl/jHERSlM8rcgGi8fHtkuurmyUe3sWK
Vc+jWq7Ne7EfWv+DkbsFt4K8mPOTyeGejM+ulykbUhaZ1l6TK4zvMNNugTsQR0b4
EGyPGYKfquVGtmFTBcjXpdRghVPwhsbResmP01Z7LQkS9lJ+gbjHt+CoQjt7Mr5y
HElGvVDwJa4z1gf2nPAzt7jBHydPKU+fa9Kdps6E43gKaJPMwWZNESofH0gaMbEL
j+ki1X6lKRGWVtuRbiRBN5zd0XRhpfsLxmUjro1fTp0gPFcD+lPclmS5gy1UMsky
0dOCZi6YheZi2o8pzXj+6UqwpXFUcwuR+vtzjdgRDsy3ftTUtjZU2NmKzmi4eY7z
vIQzhh3W7CLcPGwjOnPe0NH08ZerwitDddnt3UyF2j7WQG79yz/sPStlhEGacygz
L2MJxGvmfcyxAeK2VidjaGeeK+FB7QOM6Ep+D+x5m5Zw1pMFQAOxsvdXboi5VNRu
hyDso2wcrKt2FRzYsG/XqsmgltIPMrjpi5wpC0dRAh66mCtKsaJHpxzLmgWfrpnV
2BQWx+Z5fw0PKQE4y0yeNbWHBwSw4PiwiYxR7i48yDzP/b7xgNp82YLe3UiL8I72
qfPl3mgBMMtQamfVGy37WZLTR7NugridmT0zYikhyRYCjV2c678VUrSA6qWuzPWz
cPKR0bOR7z6qB7XwWBZQLu+xqwgpRKXV6PZ6moFrHORLojdygVM22ntVtNQSRRiY
1JueF7AHJpH/SbxiZzbt5RQrQfNN5LXqTcOhHPZ1MJklCt0GLjs3CM4DBl8CgJYT
wN2O7yymk5DSR4985xI1nSFUCopZkMmfMxFnRV3HOtHXRtP6AzXY0qhVPyUgD3Md
IcVzALjedsED8IcgttwzsNeTg5fVxkhJwvtcSQsmeekgINfN7j2bjCHRG9OjVdVP
geAbA67OXWvrOUuaZjPTO4WrwdQSDjirmW4K2pJslxaRRfmcxKXvwEXfAuFiWQXV
OvA3BedBvscbxkNuQC4HAZtVPYeAAVE45BghVFWjTkBjab2oLMu9uECL3JPN25hH
8PEDREtSVpbret6jEarBQbGiGHhlvqPpj5Nn3gPsmoLhDJBg5vG0l8AHNVFTTS+5
TBs/pg54/2fd9DI6b1bAbNQMFWt8jYTBki/l7NSNHQRvnWZmCnyUhVtKkSw5asrC
Hbnh2tvv/3j3q4ZvNatxsF+VUJxzGg4Omw8f3AahfdvVca90CtPeLrAJGWJuz1up
gEdmiKPrEu9CrQfx9PHXfagfXt/JL/PnxlXCHdwczj+CenD7krtfGR7lY9sU9DX+
yJijneHvCC6FZuTr14lAwervHh46nzE9fRRTq809g+gftEs5izBitREekEk0TFIN
OeXsw5P0Q7M4PVDVMGj8+KxlzAIzlwPlW7j6J1lMqQN9Wu6WkqVKbnEsDV9Lg5zX
DBREDZQhWWGh1X3YN/q5heAuqxYu82ZLBZCngJvcnLi8hRG7rjefF21okzzcGrmu
IKVy1AzfGZTCFOB7qoYS875MEhPC5wHXdN70g1xrJRZhE9q4e9EBirOMNJfMCyEI
nReZKV2xs3POJuvYGFAHf4tYwnJBxKhiljCCDvW6qA7L4oY0YdxWwruPVk6QjsFY
6+awigpFVVZd7cXQG62apPaoOA2fbzXWsmtZrR0qAM2HEhHPb2Gnq9LWOR996HcR
gZp6pldoO7QN7kFqD6bDRg7kKksRgTdpff46qSETphEMDNkZFcZeqSAvOPbgjuCP
Egb0Bjup19UTX2YcFndL8u1x5SOqDih5ocarTVnzV3tplOhklad9oOqJT7vof5Iw
u5Fyd1UYWbRVzHlB1FAHY/1L9KJ2Kjy1fgbHNSodXZkZ87X0ysF2wxCOR/5LcW57
/D1BPe0EbZ1gkpJdxkvNjL22ONYFl3d7tl61Ux2O9HVL2tGjp1VQhyZoh3Y3Pj3X
9VPWuD5bZC6uYGMlDu8VqhW8IJijWKL1d0SA3s75aNGBGVz7BCN49hhcmp/sTDJe
fdbCMKep3Fu3qgvXjNbzo5OgVkx+oP/ew10Ij4vniBpgKSkVjMJiMihWJA7Pv/HD
at7k/g5qx3Vh3iVCq41vvsgCeahy3YrVXrp6YHiLigF6Q7q06SZdgZc391tiboC8
oSS0VgQapi/fkjEKcDVkWHat0DltmThyIJ+c7LsM+CPZuYN1gQfAGUGQAznk37vW
jVn0IoILU9X5OvCrnnvfLV0ijxkWTOPOwGLSppzkorqIl6tBmeHRBtLDFSDMoZmc
T4da2HQ1Z5y7L4qTjHP+VmXuBtVo5FZ1YHbA4qmFharIrWZc1pj3cZUKKEUwh7qt
j+KtejcmOSsoiAqy7HFMQCgAPnwQueKf48va0ESUCjWC1jf2pImJTJd0RJvWnLES
Nc2VSUandDvxUxyC/XRYFBLwBrBnp1ouD7Fcf2SplRlbAQZOiHeHT8AQSwLPR42I
zplbh3B40xCZBCASg7UFfe5C46sbdsh3MDzIY1pligqXrMGAJKlWSawpQ7ZHeaWh
dbN4d+CD6AkJ1vQmOPc0vQzZFyAEoOcbAnoj1LlysY/QhwKPXKvwAZoH4qZQQt2R
MreXz5yNESnXR1j792LgykN2LgT+Nq6RCghdeHLGdg10PpQ5jd2LQslgve8f6fx2
0jBsbE8dTn8n7hAw/r8fVZqT16hJ7KRv3tYcTZ3+Vuf2/nYzANE66svhJbUxrnil
f9VBiVHcyLW+BQtx20OZv5o/fg7xqJvCqbpF3yLXtOJQa68LEbAwYHL8/CdNZCdL
ValnIhs2o4aJy0JND3ggQ4vEaqyPR12kzSj1XwTW1IBtw9ANFlyecIK7boRUSiOn
9PhLio0gy0AMToUXvxwR/UU41+ZJyRFZqSJkLHnoEEHvexsfbP8TG9quQE8kMFRu
wV8a+VeJmfC4NjMIQkCfOtaUbxnTs3neGvxxS8eyUx//znfJetCFdpovTEmMaFkf
gSa5WDI/APrahk12Pz1f9zuoeYsfMFdQSuB9bbccNncAtDgGcdF/nB0zISaj2avH
l7ydvUHnDQCaygYnr8H9aMqskPxWGexcLCF3XG7T6xqdciebe1UzHnp0vIt7qTML
KbC8q1sP8/3hJnIf2krVUTyOWNnKpfWWANctfQ0FYverWDdGts7gHBGbsiOz1E8U
A3/Gma3DEH0maQaYyvUxeeUm4D/nZxxDaE2yfWyZKvYkG4iE34dG4gu2ckjg5HjM
cZSsdeQQI2MbCVI7oX0d+ogiGlKg4MH0YFrCi+BHxhYnnutbYiWLelljlvGFvEG/
zMC4CEU43gR2NOMqy05WHxvFFoXj3SajLNYWsiEj+OB5kMEmTqgq7WSUBO3loiTa
c1bG6MB2LBCbMEstk9Yboh+lNjVGciZGXFxXjeE2ypQiYj2TmgXZAgUG5bjBRz05
PLQSWpqiESMaCDiAdsJE8rtaupR3RMontxxvAoscVZPhu2FQgGOLw6Lxutxw302a
Mv3ByLMHTcGHg7IOV6Z+ADzDmEgsS7t87oonNbiYFgp42dSWApQkcXd0ua4I0sXY
8Q2Z+8B4exwdTkQf9q9FDchT/93HjzYHY+E4Mc1O2g0k6SQjFS+WOyF6ZOzXbPh1
qITS9KA+JyCvt6RXWelGCKyEkK3pREBOsmSvqec3gVejQHs7yIPNCi28Fn7C9RXy
XCksaGEwjSRgl5blaPStYoMROu0lx6CIXO90IVjwrfeF08mtD/abFJyGUBLlvrkO
ijcFqTv78llqz/Mb35jLStoDDRBzMaRZ4jjiqi6jKk3RpRfypWsYq5Wcl5tgWpit
8Pyu3KUin5Neurb+vBtIAQsJpFxF5C543pCtOhu8COCrIZ3ksRg/gP9wUYX1bHX6
ivhXMGMV4Z5pZSRAVU18+alO1UA9x8LoSAYrOlu7OZDB11QMfIEIxkvdU/WfNEzE
BwTWdvueBHQlYK72FHSFcUdbt3HtH3ihKd5aubFG3gopsH9YKs5rIsBy3rQCIOOk
UXlLkHsRLH3TPmrROnoDbNDfUeTKJR54A1NzE4uRBX5wkkkMpijv9NZ++V3bqL4h
p/JZglnJu6M1p1PYwC2b+18GkcVIKc37Pfo7l5v4Wibtp563uchMTnfGjnix1tBp
Cu94W83wFV0UmldB9d2Yyy3xgPCqwfTx0btQYfSY0SwfmqV165MS7RkJcdQa6+er
AcU4dNM/+8aKbO+3ITu2Lx2l+NjB1iXZsxLLSlHYPGqVCz5lGZKNEL+GskeDgRPD
QGenlxcetINxNHXkbh241CW5AhO4GKc/GdLkymf2IQqI16rXnhUY/ttSD4pAhLNm
UBa5eaWXEFt0IEsgpmqyN1gttQMo79HSckxlFdoqSsw9zCd1bUMTbj/2NaWItWRf
bh7ASGYvqNt6QJxD6oXWvIjPeoM4z9L1DL6g+rFwAat/1NMVXOWCALd1C0eFxxOO
ecPxHk3r0VOioVpt3y28MzAMAjnimxqNeqicjcmpm5JI4CSXsxTu2+glyrYfe6L+
K5NTYBOyIY0Pv/cfCMD4gDiG6hNqmQjPum90APEhma+DHT4gDdFgT5Q0xzgxBdgQ
Q/fuLKU4ujTczp18vpS5u0dD8oA48U2axWDjDH+gLUn2RF/Ztk358OGwL1/dGt5q
lajEzCYtJBgT75UUZ8o+4/DH32uQLXyi8SVF3svsqJVL702GXZz8HNSxgm/Y/Czg
v8dN7wjSqSRhctga4Pdb7KJG94QzJm5epnK0ApHZaFiSoIFZtCU6iH50WL+UbHkC
oOQdAIcEEzLPPaIHYAaNrXjUnb9lst6ESGb5iyREFj7FxGwf06tqrFC5GcX7Kgfz
ZXb+dsO9L7XIUHjqwSAqkbPH7n/fFiDS1ApEDiEYL2y7PpQi1JOczqxvJKM8Kr1f
RNn8w8OvXSqpixOlGJD2PdLFLdEgnCt1LofhmHJ8kgvRW/xr9atjoxwzdeFeSLtf
JLQdlQMpvaIRb//RRSHSuO6ESkAJXmDP4mjX9SBTx98pEDR5ysBKvaBQtO1K0Lzf
UEzW/FawsKfKXn1rKbCqkNkbxuFX2qjGUA+08ZwvN96OYTgH61k7cXEBV73iMPVq
YPgek9sZJo55E0pvmINmkbgAp6tGXv+1SU+mffmwp4w/jpsVMyrCSodolkAfpLIF
Nf+0ym+IbxwrRwFAbjVsSLnvHy281CvsMx4RqnY3sXNK+OleiK9vt6EI3lmUkb+x
/aqKPJbQdOvf7c7UjoKMk8qu4q3AAkMhAffecwnTJDVK3zRSi5+NSx+dSuQkWZ2z
YdqbJnAz+OBCDNrAZeolvTa+cUFb+YtSjl2qSHms4IlITKzK/s/zjLowFRCDthX3
W1iARIkhLJdWCTwTDLK+UKBD24eMBPxxiAivfb44u5U/G0AekAwWOgyir2t7tus7
pHemPWjG981MZClP0cPfGrxHQFOMZx+WK+bTAb/MAcZPxtHcFp1pfgXEHu//d09j
HIhoaIcG31jy1Mcij6FxG3yTxK/vLfQhJZzxDimPPQG2UAGDhsoGTr2VxyhTFU/0
dzAgUzPbvON/NTpgsmSaPF5XneP8StfKuW1+5M2IJO2NJm8/wMYK9t8MH/DdcO9/
38OsOuDwlrdS2NtZGcjsseFNmZ/M85J0I72va09XR4wedtWXlpDpVncw/OUN8Pmo
s20ru8IjSCoReEdxETrOG+cwIf6MKE/5FarmPRknSYyK1a0tBsLKTwtZAirg778E
ejAa7dOeCgYL115g2FzNhfhX3DczemVgQWYkuxjRJP4+p4nh8J6ME+ZRlM1xTBow
Te1ancbjZYpRqEarUL8cSeSVK85qDBCao/MUwdC0spwzj38ILnMUsmlRUaq8AX79
IO1K5bRxyknlQ2jKgqsdrT3Apt+DUB5m+pidaDMkO1u0lBqPlXfjZk+4WvT4RH+v
RqXAPczBV1ozuMgyDKGHo1iKDeghoExfqVSmndC4UIYSqgP8cn6V47cn+XbMpgmI
ON4peb3VGpUSPBWMKyJlPfPUNRSybHkmbyy/BMehbHtr9asJpKM7Yhr3QaxwhSKq
RiZwYla17WQbvhpkD45eqdcMsvqS2gR5Ng27FPHsEs1T1VbjekeQt5kuP0F478An
qYpn2pogRwet3c8PJ56u/I6k1+w3gcn/k0IPxFYcuJVeDiD4wDmQUFcR6FDI0fAx
7W86+/mvW9w4NIm1E2tk3OBThcKW7glnx4Niqm3uJC8cAdA5V0eUDuSWJ+t9Wudy
ozGU7na2sBiBJqIrh2pOydLmPWi8/HR4arNyQwzp4AEZ/7/BbKTBR5ABLL9u78jE
POWO+5CfRNflrDGwjn8z904nZlvN5zA3uVdOhdQsYDHAPJillSHJ7Rx3yLVSn4+3
8l50ncA1nQs0nvp3rfhGnmtNTSbiiouq10WlEnHoT7It/QUa1YOcnBAI5JuKZ2Zy
T3J9kQ99KqeO+HYZPnrtqO5jWupeUAA6y1o/UiNcLpS/1/i81sGWMbDmsV3dW1Vq
ayYVqAuKs1B59Y3W8NzrvK7O4o23HZhLamisucVXek8UZHg6pUjWxasCEU3SHTTF
JUUPxuBmZ9TbZ+yAndsshcD4BIWIGgsDd2NIklrw2jFonmBildd8XzEpr3pN/w8U
PmHHdycgrNETjP4eYOjc/9WNeUzluwqyXXJ+lSSMLtqPP3gwL2q1m+Hp1EtAnlWz
i5WMt2QTMmtKUuqyfydAlifEaQ42GDCc7yti/803GOLM9fw2GrBvrtdGfob7PQ1+
hr1r7KfH43/89LTNUw1nBNhlOhnA15ESzu8Vgh+bA52Uq4CsT88ijkQ0FRexUd4j
YuBBmU2f6F+Ttep1Mv93LFwYX72mgD/BQOrJ+J39DlK+B/WK1FESjA77pQvskyL/
J9jN/OFrt/2IlXKf/In6wlEhBK8U2vZFfwGYU4Cs6ZN4m4DD+TLtBYqKerL0iAq4
RkiomWEgqJGS+ZeuAPMmMBOqZ/F5Cbdd2aPgxejPskDnsNqFmHAe4J18KzyIF1a4
Dt8d6QHoojRxeLpmtPMYvdimSZi18ZI9TGzRARO8VTsWRGA8x0xeSc5YReBwK5Xl
qLCluNi88GaDhsaV/uyTEb7x+b33sSzHz74CNBn/MikKvgmyA1uKmSputjkODHcH
IcXC8CbNl2ngLBgzbzTjyixEk0Jw0TCl6GwGFSVqXmWMUBd5pc8hfVNmW/KzsUcw
xTRAcEjf9A5568tCvRr3nDL/8w2yDAMDJ20Xfe5ktfqOPh/ZllptZvbCc1wUw8uj
mexhbICMRSGgWvy5AdiZOiK3M7UDjo3I6VBvtHiYX9mjcf8p6VmeGTKkgX4TqsQa
CpiR9lIDIf0hvuh0X3j4JcofoWG6i/6hBsOa9kZmQVRLaBizKlo35DUg5L9vyE5E
WgfVRaI+tLBNC/0Xf0G0CI0j/8lPSulUOpiCnZIWX2CJNf7QiJbj1yHpWOWe+Ro6
1HRv3tj21Jbn8bNeFIarvb1BQ3Bvl5J1O6TI0U6sGkUUVEjPasvggxM1S4v3jAzU
C9sNfQWJQUvAI8zcxI2AuhOmW5n9GQv65XfQitGgv/A4YOMadUtBiearQupxltuN
Iynm4dIZoTgGI1Jv4aAUk01jnTaHRahV9ALLuhDrBFmGUoocy/Eg9JTUemt7SC9A
VsWi50bPlXo1LbXt3hQQWnRaT8vDVoEstGMgno/zYSPsjQI888Rtc3j062DAztef
9VtR9vfLCxs7eLi27cDNAGic0K9JD9UPdx3shbxNsgLcYdlpYXV2ykJg7nT2gYLT
1aluV8jgeojNMkttPU6S3x/o6aIp/Z/1KIua6+Pek+dYqxytoPB+3MK2FGin36t4
sdIX5WELh5wOa4oYvNwQi1sopycemncXXC2TKmNOvN556Fq/PAurofjfD+vmrcYn
he4TASUaXqhkqdbZYGPcdk0LISYmQSfe6RQIbKWImNZqttYvFZbkMxDruPz3YTFM
UVJG5NxbWrlMmXscaDVvBtmED3pRoJ97OPmNZ4JtOLW4wWus9BLRB/y+9UAcAQxE
1MuSIoC43lZR6XEwmaHhGRICRbQC7SK2fT36oyvuR1wH3d9w+hLZwIobnuegZ73K
kC1Jnouc25CXZeUOwV9SSzOnu9i6IlINOqNqmOQU7Lr/Q08UX/9CUm2urpBpZbdq
1s0NXqNGOK5LFt6tVm4I0rgV5vaoJViD74iszyGxim4gFrTRqo78QD6dYjqhj5AI
MZHXkBGLr86gX7NQSXkjLh/WCx20qxi3cH2LnK+u6X0cWp/BPWPWVK1TLmE2cuaJ
OnnlSxnqPe9ncl090KYdNufUHoEwZVACs6mKkTO/cNcwdxY0VVDocGk4t1MgBSL+
zx5ho9Gf/SK+GVmXHjqXHU4HNNjN2K8qBEWXFcM4ghur+rjFleHlCQVptXhxrM+I
bbVNMmaw+pPLQTj22fNYcl4ffY7ePuKKgvh8wrFE6L68j4uki3z7khiUzhaJsZjQ
r/G8hUUKB4YinLJ7kvmIkudL3WEp6McoII4ELKuWIBjUU+WsUFYxfjedbtlSlO7F
MDCcvPPrVHVevuJ4ZOqWyBGAaf0njd/fT4s3TzOejYAe+6CIwy5MfEME3KbdtXss
SjZhh3B1h9LRlJ+d4x+ySI/ZRrTLRxJSR9OhbUegda2Yn2CcX30a6GLcQbcaKJI7
YNPsZ9COV6wVcXswLNMvqmnvjgYhhIRvfWEZBtivVW2U05FkGA5pR3b0U5uDMc9s
FBXXovpcZUSkF4wFWhtt70GKYm8ORqa5cKKPVgH6+DwvLwslm1ZlQUwHFCRP9WOa
yVmOEp8nDXLMhnwKsFErRN4q7P3b91SEEysbIzHfMx6g05notOgw9K3V6+tma7Dn
8rYRNCC7a8hD+OWPL673CRWuNnnFYk6qbeJ9HO2bitNY+FLnBwnMSwGF//Jr7Hcm
+TWl5uyinaIkTW6N4ftqpVH/V5i6dA1XDxhadFaLbdKiiwIQGnOGUhveIBHW+VVh
B1aZV4poFs/adyBIX0jClqPM7U5y6uHOWPv3owLA9XpkNmNkF2AhL1XsjLBm80Mo
6nM5OpoHqz5WvcVl6mNWBFWdSnlgWRO01emV3Rygr7FHOhKg1PcpVbn8U4VmScu6
R4PRvaXk7MUT42XWYf++AHvBZ03EBaQ2lfvKnpw6bqDT2OZ8Yue+upEZwYR0K+Cs
xIE3UFceRZilchJiQhNiSUTZK2pR5Xx2Pr18d4OZyJ1xvR69uhNPRMz7ZTm+Z29x
656Avhm7SL24wn4TsjHWQ3M5uomzxEAwVeXN3MSr6VcHh4t95Ds75ADddGkP20OM
jMZ8QhMfiZBsDd3NO5h6/tHUyk6GfoE4se8pZYjHwvmNyGQbEZslJ77EnCV3S7ze
6Dw7FvKZChVLKBSFovXJyAR0/QlyYsu5or6LmPrP0nCvk+LP0qAFvSHLVNd9hZ/p
rTmVdc/TUpn/+b5DOVLjtJbLfaczGXIsEkI/I8hPSyyRFWGai65EaUd8XgWYTeie
THE5LtcyDw6wbKemKQDDfHR1fGzG4V5zQ3vJdIsjUw9KK1NvyakHevYE63Rpmn+A
JZWVomECdGrfaN0eeVvmZXrh0QvQ0VZBqdVTdU5W6qQEVXuvwMIu8LyQCbNJhqmP
i81hYMw5M+EcZ0r15GM28RvnaDp8Ry373c4W38MaBonnxpFFXojIGJ1+u3jv9SvY
tvsJhNwrARdGnE8Vk2Rq+I0+YfJqXDxQgR8l68a5Y4HrUDWbGV7+8rCVpmF1kluC
4RqUUIzHF442GolBKAWZX3Q+ZGGylbmSNNlhm7XpKhNTO2P+eW14YlyR/Zgz9/Yb
OYtueYoWv1AdqLhtRPNUzQy+HCXzb6Eq5ZvbMZYqhy/Df0ne03EjCzRGhcivUaRV
BOlQgJFl/6Z/ZSOtPL0SSQWYzurG5SfKbBfQ/9qK5PciraWN5SZYQaX/7PLrQ0qQ
GQktpl07l3XSqn+uCx79pNpxlbzNJXanQYbmDzyqDyuLUq15EzHKTgfmCvv/doQT
TUdZnMpoRkHrfBD+M3q9Hh9EFZN2T1lTOSlB/YIc90xHEBAXkIRdELwrtUy9fb9j
Y7QtW516T0+2GSXjLv/yh2CP2uQPsGoTWkJx8EGl0QNTkDbtKrm3JX2gGnBU1z6q
3gBECXw0mGWHqv2ore9me+ilSdzNiOg/v8GlAUXGJ9bewHc9xLEs6vHmPzjbnZiO
+ZZ/hJiSa0BlB5wF4bdg30rZlyvoK7lqu532eKDOONAJZAmGe9DJN2r3XIPlX+DU
nsFBPDyXo3KpmzsZRWbhm4TYusrOvEIJgTyn72NAZh6fVY6RQZnRFh9YTJJzMHQq
f5QiZduRcuLN6r4MPlpuod4CdI8EGeDTei47sWLpNTyYtKzy0paknM8O22Pq+2xj
N35u4JtCXwzj/OdfPsZ4/05cC3iAR0bM0OHnhZXh3LXdL8TNpc7QwukLE0yV4KrD
hyq6VwCPEv7wU07kwSN7fHuGf+uiDHVMF2mILlnDpAupVL2YnUXyWXrqKr+b1kea
GoEg0vPTQqyoI/SEZeaoIFR2uWai0ie9sq7WYo27iuhnzCnLGxL7Ogbd+LwhGT4D
FE95eVRZOMXavtXG817APkbuxns8u1hbewKVzbtD/prcfwHidJDQiBDbrid/XmF6
xOvW6KK50lXy4ZXmsyL/36gEkuzmWuLaMH2ShfxBaxwyFeWlDARFETvH+fdg3y1z
kthges2kU5xoaQdEBoADhBuphME3ISNwX0RZEO2AdaefhxWh/Xmyijz8mYgJgpqZ
/JsqHi7gbSeDurIZ8ryKOXHXHa/GtuvcKmTCOzgB9oIp1fYxdud92xVBECvdATFJ
vEJSDn3p7Jn0w19qZifQ4WoVlSEjuEhT0YVM55b/4EnBSljks5C8NdlZN/yVnsBd
wZ2BhmLwa873kSCyp0uT+FHt+CIVnyQOBhSjcysxiaYbJmv7+PhwKpDSaIW6jt1l
LjfbwvGH36dUaUsFyitnUDvv70DtHSbxponkJpQNAhTIfnf3awXF/5CPpl7aiJYa
gSnwVuiuycmIOW52clj3nv2lYhELtR/8sJ1Fw8+9edviOKOI0BrIN/VxsMi6BQkT
SAO9SYhAxACYS2rtQUinOdF9Jy2MEDP3GTE1ZP4KScLlT/uZoWj6pAIiBkLAkKeB
p9Nz8nqypc0RdWr9AndcyXeSApeEyBUSBDmrI8RgGcZ9O21eRvl+M7kaazFGL6M0
itfgSbGCrYkyx8qxAjg+hZdzvkJjIWce9PIl9igr4DUHkVnEy+V+94VKnpgeARFO
2jkb0WnjHQoWUHvKGBOTr/L2RIn6qopB6rYybgB1yAX8LBOEl2ur9To+5ytsKiqu
BSBigRhEXpuAdwpFI+dI8lGQIMLTRByZUN9O3vfkC3vvJGN2HOoLH0XgC+uWyJ1Y
vQiHWsPLIJhdTELDqC4BBLV9EZV6xEuRcUfNmlyWW3/h1GJIhF/NhV8QauF/OwXV
Vy3NRkqUhLJcdtpycsH5rlpU3d1pu5sroVKhaC2JGRKPeI5QeQjt1S2ex9gjKbRV
OEw4vlLkNOYtGUJQxXxNhCD0a5EfsdgT0orQ/loBGqbrhF4zuqs8m2YtS/H1ZriA
KTUYE+epLWC8USZRkqWip6/NkmZYsjmvTlgL4o+Sc+raXR/Zf3x0kOrfgI9RQKK+
Uei/GY63h4zcxiuT7FCVK15e/D/h+wOd8BjshiT71OEN4MZzjwD5IEXHAO6HyT8C
Hh3wWt8MwAA1sV3XQx+D3FrdTuSH3eCB6wDF5KIQeO/eFgnVXrzbF5St2e+hgulU
frV7SIs8mOJ1D7uZxGJTS+OXCYnfY4FBXdRXFV8rk8Ey7wDE9NIeBXt0j9LZhTJ2
uPJtkOJdd02JlKEwwADaszZmokyUiwz9JPddTPPcGtiMjlpsZBWKyzRKW5LCWO8X
W4VdYNnlWi/km1HGEpGW273bP5O3/XBhlCJpuaCWgwnkJ3wOIjn+VXbj8vQUng8p
re82/wsQ4byy+Qmquc0S0/7jZ0GwYSF6tIW9SNITkvXfGzX7oYf8P/Awy6nBeZ9d
RYy4x4XRR0r7dbzjTxxAFi6618m1Q1Ky7r5HDPxCcntjH7I/idWi0wTXsG5zig1p
JQPemZkEKZzzSg1lAzGSae+1BhDThaWx3HjXL/vtfVva4OJ6R5qIPpEIUpKYfoRq
e7BbNHlDeNZznXnmzoNUbv2i5Xxnt5upWxiJXauF9ZRiASQfSqNdo4qvPew8r7z8
u//4t5OCmFzuSCol0JI/K+NOhxeZVcI6UVCpt6gkK8woescqiHWWV3h90lvcgDh9
MxUjAkx10Oko9SLXYVb/QSonVMZiIp7VHQ0KdTxpWvIzV0dkRMQ8IcrDZqCcmKKo
qvfWjL0Z3LofowcOLjFUj4vjoQPHq36WXmaeAMVLHeoFxkOP+vj08bVQzST7PUDO
oXKivuNd/MrWWucx2LV0n2qCch3jCyuAqjhdNbuHA+mshIFI7Zmw9AXMq7pQ27if
tQccxy1w2AtaevPO7q+F13ZSE7/ZEXGPXxAENXyfZQsr5Cq7uwCkoJ33xA9UIKux
IZZfr7zLjsEBKYXJqyLmYeHOvQTlaMlvVG50p1D1i6uHwGbePCEcPPF6TpnttSAf
z0t17QfSf6zG/TX4nqXrHq105fKFRbrXKdMIg5DYCRX57DyE//oZkU/uPO9kY4rS
ziNrbrEKnfAcgkeH3yW2ci/mmGjXz5z4tAfFR1Ww6hiF6hZA0+OWu5ZtAcGF+HU8
etOWMNcLDnn13HSZG/6TWEK073HUg1JXVDcJ/lEyagrIrjPqy9YBcneQ6z0F6f+v
Qw0225vxW56tgwIjh6L+RiO+mHKHXFq/l72j+LQ7bGYuZ4G3DgsN//06nXcZBGEI
oQJvOhFsdrtFIOxegX2gQ61VF8mlBER7KfO1hrPvFwJ7cehaX02Rpb454PtNGtvb
AphuqIAqam/QW3H/wAHd6K5Ot2jb1+igYsfl73bmdLvEISOpNHMd48jOtVY2DYDb
7+0KlE9R1OLhYEcUhPrfCAKl1jwdkTOfbxFBDC9tPUZZzCcEgP+ZT/zVkRtZP7jC
ao11ThTh7mLgAhf3lsB2zwlgwslk41+Gs7ttpKoy/ial3zgxYyHSeZBe9m4Dm9HA
e5aWPZ5fdLBE+w2pMVpINnvaalaMO49BqFt7vp2hxALOjei7rXRH4ux9Hqy1WdaP
PgyiYQeHdYMoTsnSxX+DdDcbji2yK/l7NbIgq7ZPfO8GL0qTlPrqnpiWqM+XFlug
Ynp521VLyLG03/lhX9TpDuPStEE3d7y600FufHz8TgcPSVnHkpczojw5dfAyPZtR
CtwyGRyVD6C0B+7kekvOxj+/eF6tlccwPMikSKtDm8GUYViAjrZkZ15X4/AWL6Rp
43XMlw0hGOqV/iz/DcGDeqJFYvnYC3/kBmO6nSyrS4M+odpfRLsudHAdG7xtw2FO
lWjXAfjTG82HTqn4ixzeHAxFRc56Tm2rDJ+4KHOTdcDTBuzJdsRgBinEFznlrMPW
CUSqZ/IAoTEx2AQo955ohPjMI2D0iA+hyycgXNgYJTItxBAbY5BjFcPkFqUJQrNN
rVsHe0K8lnJTGwHjVh6e0qZ0gAmrtlBJnVWxv6/ZiaTR8+Z/8t6utIT7AKtB+6s9
yQ+0NsKQ3U8EoBPUtLYZ8FvgXatIL0HHkb8DJ2nL+uEZbb+/L4Zs5BBMoH7ZdNCK
V/F6JKIkZbLqE9s7HKU0NlS774FXhbUo7AZuLDUtv7Biz7S9bgomM2R2iMLzwKJL
h3Q9h/jLOHT9Ggy95MmK6uS1Q6N7D1JZotv+bGuX0nyQdKMCrdradjZ7j3UAV6rr
nsEHTf2w4CKqDCAZe88dp03wm7qL5jCzBj7Xk+2puWmOxKSqHXN8dNytNpsmr1ET
Uht2MgNKu7dibGDZCeRdOuYK6S4ef74ybL0Nv04ALbPbCnBMqDAh9sX/lUyOdaQZ
/1ou9eBktYKYS25ilPOh0e9g5C0IbL00ntT4Wt2ZQaDysBfdlPv5WQtL9TkVew4s
qcjkStHQFvRCBLkipN68S8h/RZKn83Mg5pk9DCRzgHIErbKIIHayIjjt+kH0LLq9
Dc+N0u2+neBPaOWFt+pu68Sd4rKaoBjw9xm2uzg5SeLO410F+TX8Wf36f5T7nHTj
FDIHDN+sBYe8g+gGjQp+WjQN2+JrpZ7IwRp8HEvV0UPYgD6A4Yhjs+RpEylB5n42
9hceJicneU6wqxDFewH46qTHylhIzjFmqXtd9qxq9Uunxnk61i/LXgfljLDrFYVv
UdLvyd3i6JTvl5RdbEvLZ+zFol2o9Vs5mP9b2pCMXv2HdVLvMpiauygPjT4Blbwr
yuaQb561/HgDhFYCu6XVf4CTrzk+swdwr9UEtJSDpfZtolReVnESpNIkaqXB/TTq
eAOh3L4vG/doUshFYRNlb6RNNikKNqtoh0m1r03MCmMC5cNw9Vc67LEw4AaJ4p/E
xDErG5PHwjjAOsmTEdaRIlOK0mK0bigS8Xtsc/ASI/YPLqQ6QFdUtjr/H3xVwAGb
ujidmigI41vpXN1DWXVZqRCtneGB1BMZ3TaFZZmAipsSuElKrMD3SA8MtiN42J9o
00jPwcOBMQ/Hg/2fi49vHy7GyVO+ZJyUuTfZpgiOskKy8YWooUYbEJPe/XsbozkU
WJX7//G3O9XGV1t5xpXKcWxEfuGnY9pxLFXNry57CgO1JUWzKDipDNX45E6VL/3s
sggGI4fx+F4N+ANpBWB2HjuGk50lWSL17WciEwKLloeRnFfLglO29V+f6pOSLsNl
ZI8ezfW9no9cqmFOov3wDsbfkLL1BN0tYbzmCUSiZY/iIlkVV3YlyDLuL9HFDNo0
xmpfVCzUWNYX7V6mk0cgwbhJrvPxzqVmvz/xyNy7zuvTBrg0y3pxS64sXuOSGWLJ
j8TxuFs7cO56l9y2QwAeCl08Kn/2HbHxxqXQ3nQfsQ3oiYPYuES8p36TRy0mHd8Z
sW9gIk1XPhMJ8ztNHaXCYzavT4Omjf11DBROh0WOnN0LkfzPoZj3wh8s50Bq6iVf
jUtMCqA0NlfSDVjlP5ZrTThHI/2QpsRGUXkK1oryncSiQHkNblMXvSwLALLvc0PF
3DR6K62utrEUyzR1UyHo5veMkz7sc0vrF3x6c94eiV7nQOs6RYLxk3wMZ7FqTgtQ
53wtKs1JmhJGZufWsEnJ6uR3EheN5HAgtiifVYsAmvzb6t0AecwanmXSubT6V/4S
F26izsPPSjSiz6REsujNYbNVKCpBT8zvb/apgha4bnGIx+Inc4KmxJfQHRVFWtre
myWTOJbs28Sk0apNaEZPW+OX/MyBuWPoS+Ay5fEz5e9F1YguPDPtfBbtnvWNdpvU
wY111o62aQzH97lp2phzlBGgU+c+hgPLjWEhKhs2rD/HfdyUmZHC2AjqUuwz6Yax
sTgTQ1rKwKQi68o/7iow3Prr4AvYKoro7GrhU/GxfyWPj8y/D0RdZMgiPFM3aYJ6
bU1m1c5IlCiO5PMeKm6jtajWuZztfrfn27csKlLeuoq2bNY/oyB7rrqPDEEbs89c
hi/k+EU3aF/PskDe0uEKZGTLXIE57b07tri1hdJsVW/1cZa/xrZ0wOsLVpNZ9Mxl
YEk9I7USsmkrtTwe8xMQ2lwfBXVZPYUUzcHyvfhGXm1Mmw8EMTSG/RtMDA8vjHBv
2K1QgUdiDqC8dVZfwOpnej8XB9i64IZZmeoiZcX9nQhWUS63/tHj8c/e+dvkgBXv
d5/ued2sQvzaatYF+adtjpdgDcpcgjDvQQLaLKtwdd4NTU/BiurfgBe70W53thlS
3RaPBu20hArGepKRRUAbNf7OQToZFK4E0nWQgW5tcYnjdzwEghw9fxAPB0xFeYV1
zhkYN3UmZ5a6F88nNYuoMtLxek8lrEnr/iwbBRQkYtr3Sl97ru8BBmx3HpQkDVG6
gxayA0bMwH0Mnawdyp22o4bibHHPqV1Za3IjST5mfdgsthN+t/GfKYJNz28QJmQF
p3HawXSyulIAdjYDJdVRmLP/3JldpqlITAYNlb8UedKngFe55FEMzSgB+3MDbe4X
7mQ4YEpr04HY69T4vPn+JYBKWXlsGmA1AI8R10IM61x2lHMpVB7WNUTYFagL3X61
UCjFZkBDZw5tubmVxuAuMxfkMUUSkRhg+MAuCQGOCEey11jUtllR8jLywIIwaqaI
XQgnpmfUht4I/qV451HpYutf5/L+RzkMrLSug89ZoGbH7A5EyaLIg5qWQbGvEmJB
pu5RtZmjrRqdwBMe8Vxojz6zZ+Jum/Zuc4ASQOTprDHlQYq1tQRKPJA2og6GZYHt
KJWWHiHJ0iAiOiswurnWyxls24bLXaBKrdMuHIwwnqlziIEcx9ZP8OLiVghGqj9i
vYZtYl+AOhTxD0ntyRqc2KGejBJ9j5BjPAGd8TSaDxxOLZlskhV7BEq0aslysFi3
gGgWoUWUh5v62Fowf//gOKLhYUQSpYZRet7dhunzRtbsYIWQPC/X0b+7H6GjRaJo
e7tftegpOYv6xdj+lLxgAEeQsyhhI5u0Ka7ypBKYabo1+29PFKyjQ7Slv5anuUEM
+ZSXZQ/sVa6g/iEpABbDbY9ie0bMZFw7Pi6EpchNUpTOlr83r6sd793Juv7pefyR
jrZEorPl8oOR34yrCtvuHkW6JdVtXoNya34+LKrwBSkCmR0nZOYHSVgukq7tPVwc
rHK6rhHgJNqMvrn1cc83Ut3+5PKTMnESehXevakQB1Ij/jwnXTHvDOMJ/yoK0pgt
mkbMEVPl4Wixwfle8SOsqjupNrzAz2WCoql+n2ctPk1Gkm1JZfOcqiOV6Aw2qeer
r8BhqOAucKHnQC8fix6ZBgNO3S0Sxz/EDkxkauclKAY9OJa3TnLc6bPbCzA/1yAV
eNUro/MSrIAnLlxmOWT/z7dEXSHzOVUKAGeeB8ivod0h4+TwtEtLBmF0jpbGRKU7
L0ghX2BAUXChtm8CbsmSoaUSoKGLZ5wfo/urMqziggXiW7/edBQkWIqFFw3mKbv/
LLvWQGU9CCcww2kGsx3gQk8Ihl3MisDpkxend3xbGT7TtloHg+MPfiXB6xBQAWik
+0sg5vjI+vL8XzyR5VGlkZ9mqOOdiIv1CJQe+HbXZ92PQe2xPmdoy6cjdF3BbFdY
ozvP8vbwojNb9lI+fwWR6GbFc85k9cicjTarVxuYw4a/NU4YnSiY9JPkwWQbsdpq
XyV7+56naaCCKV+c8Vw+g6uzEnt/xeBMDWl/nwhNwvbAKKn+7DDW0JD62LfuVaOg
sezrDygIpVUBS/M7uUe+cmcmAjwUTvwBBmHy2hZH4pSLS12XL0qXWAQLX/BZckfy
jPhTcexuNHGaC49l1CIVZn2zeyC7fLRbSRXY+JqRYhow1Im/zTofSD+SVGbtoED5
MI+rC5TlzlNd2sKokYMLzaaw+RniKcmoVdhxLr5kxdKwUQiOllgSHLjAWnFMifD/
jVMFn8dTBYf4UygGBX+3HO3rKr5TRjadLge/wOe6m8F4xQe6vlimhM+kJQ9cKMu7
hx3I0XJIaAz4NN/4xIoFwxrn+FT8gD+DKUBP7dah2tCW/AtKT+JRIcHwXO8teWN+
rP2ACBfYag3kvtvJBsYx5OYaTSYq9W2/ahVdRLC+QqvhrBB2kS2bCGZWXW+QCMsM
ufzuB6IZ8yICnBxt5OqeqS/4aZ5NJ74uhp9KLHGpWAJrIbmy9qg5dQKf271cF9Qp
0XkbVYlEKZiAyDPO25thad94vCKLjyMIhy8NKhBwgFNlIDCGAVwFo37wl3A/h6LD
6goYanD2aartf5Efa9y8xd7YmlIOlc+UBuR2dE/SC8EVKniBJ2PEJ+Vj/hvceYEs
0Pm5BP7niDBspsXiPz5wrI058SW4smevthArreCToL4JGV/8r1sS3xHVvhFxduoN
Yva8jJgfkGvVO4oelwuiAcRQCR3/qzKMrGSaVC+67k/B9d7p330w1RLnoYXiClZZ
/XJKN1j7qPTZ1YzaXubYFHU9oZHMxj2kfnUpqw4sD3unYL+PlZFK3/0Pbip9XJgW
sypA90snUCSUVIQhnFX70to6glHubGQJiaO6idkWh6yEs2H9aExQiR73zk+wSos+
AygZ60c+bIUdW52JyP6CNHnhjbdgO4ysuGmBeR8+RisCx+tHrzMNtrKUoGhJlicV
ZPrHs9KXRLPwzyc5G4PfACLCKM/908pHBHHpJAl+RFMqmzrZSBIRunaF9JHCRMMR
1Cvndxt8F4fIpHyfHMcTSzIN9RFWMAy9lPqVysMu5doKvI2kM3JlqoblZ7OjTr83
IIg2W0lBS9B3v7Tt9BTRzvJ47RvKzBxMPOQ9/qgvxY+w0rg0erWPRQoV6Lx2FoYL
cHG4RidJXoDI8lllX4sfF66WYPkSUTBf0dRr5c91DQ6OIyxddKE8yzxeyI93mlg9
dDPSIusOdOB/Rl0UxfVsi0lc2t67GK51ZHxbUIhp8TZJAcWN5tYB0SnLCmRNgnq7
t5f1WTk4xa1fz+48G/kElZ8zo9OZKi+OoCft4L85qaRseHIXEElt1kAocrOaLzL0
owB5Q5sZj/JvfPL/eXXzUSN6MfhEM6PUTm//lunO71IMUn2V7mIruaZvM8dyQ1lP
Y+nAJow0w4+6E8zE7nQXTmENmi+7Ae5lMj9J6DKIfElbLus4bu3kbalLBrA3XCfV
pyzLiYlSSmbdqvlDi/c4hu5ajRYhV/cX5yDGJDK5B9PFgQJpIWCknQRUIGDNSb4c
AZW7bibAg/v2QT/d1ukRgsnW53sNc2oCzoUwVuArAsWT9TeGsEBDlTUAnIMTm0hg
oMIe+mbDjMgLr7KQg/k3Fsn446WfrrySOvueIZ0VdRr9ohhfe5wa6JjUDLx1iYxX
dBiHg6oaJzw3OmX3KclU/f/1leB5xJpaLg6xqvNY53P2cqv/ecI/jH+FqULjanqt
B5PdDCB1QcqdyNaPUVglqUi2CltXPhliHieCJym3i2ju32AhqAuR8nBoTrs01RaL
mkLg7QxY2MxrTHn7m7bWzwIm19YWcFYbBeDZtBsK7RH91qP4uYjbb5NQuQ8tyaTQ
0xWZDje0n9JNsh1ZIWqu0EP+SZENIGa1inN4CvTCr5jLuo60N6/Qj2VlGbjHa5hV
VnCJuL+b1emH8SmbLFVxtqY579zKtVADI/GYi53vCKwBMB5cv8pC4ibG8Nmv3Yyb
A8h8PewfHpJc82n0/Rm4LR2PvF7NczXfY4jpDMcjEoiUW5TSoW6Wjj3q2v5DI+4S
UTYDGC6oXkrJb1uUDVpWK1XjXMtkFIXkjqL8MCcqpQ4adOUNHDo1ye+FF1IV320H
tIKAKYpI6wzp4WlmvXmx5GaLwSWU3j8zvjJGwQ/njg2RV3qFzc0/eVtHlLetAzFq
0clzAWfOWk45Uxkw8LrPCeFoUoNwPI5T+12Ki4mI5kmuVAsMS6McPdHwfd8h6vyz
+bUH9jd8BCPrjTsuVRYQVNIkOdvd0USUFrYbwzZ4Xsq+acJICll2+oUoMtiToEaB
THLqEmqvScwEgLVmN/FO/Fk040X8N8oItXfVXVleYb8ObDdSDS3SZnkKvOVBYQcq
JV0RVavJ35b6Jwm4OukSiQfGwgCyWiSDw1UIOicNTU3jS+JU4LrXMUn0cbJ59Eba
Imnw+Aeqr5Qu5KPuOcthYaeqHPHTfUFljzRJES6h3IIhWk5kflw3F2cLlGStvDTy
Uc1xpkObzsv6BJOSt0bdqYOxaC+QWnQwxBkug6h6ldTkSJcovDXAvoWsS5bl+uyf
AEKyjhGLvj+rxXJKp0YRP5uc7S0p+s6EaEjBfqZPisUadLQJViNY3UnKBea3k3xK
y5t5+ph9lYvAxjbGytvYlF1RNMrXN7/rGcKOOKcUuEaK87a7YhOtmiv0XEPHcLg/
T+mRJab5ej7rvedMoVul5k6jX36HfEVyhE89PGeH8UkzzSvRAkjwMciOT1FczXpD
woTpa4pIq6ujHRim8K5m40i4+xsFLtwxnTBvm+3DnyZaYXD5AMbl0dhWRsNCiRgp
jkz1IDMP50u50rm/GKSNV+AH7giIL8X96w5AvDLiGDlNaFGQT8DaQnwTRAYOvq7y
s1OQhRNxrXY6FaOoe41TBTErs1ihUL2Nbdi1VYmrWQuyMw9Qrum+/tiFniW8ehrg
bcCqqqudYOpRCd8TvDnd2sMnHzn/TpKXn2Ubh/W9fMEI/5xySa8ydC3aSnGkimYK
wgzm+IKwEUX38pBB6p2FdTRmkHwrt1GegHD/32McQAKD2ra7tWlem8KHBN04yzn0
dSsa/8z9HZihN09gxvPeynO4ckeyJy0EyBdM8MYOqY66A88Mx829Qmg/RfPeSbii
S3wUGalbcBxuAUXUbvQ/CZKPrY+AVtYL4rI89sMHCTWzx8ydYzozGQx6Hxw40FW0
+b2QSv8XPDtjLa02O/wrBQqpmPIUo6hRujhM5QnjoWvsfwvYQahMFw28z6x8z+pF
po2BAQFleGwT5D7PVT8I1PxHwknrOKd4cwuxn/Tu7380z3hIMNl1gMK4jucT7lXQ
QImY3DZUZJmkmafMIgCa6cSxcUQx/aabi2syTdD3bMrWj6PFwlJ+zhWdau2g4NRY
6fUvMFweHGZAaGnV8Jr6SQz74N3MJxnPPTe85VkZITJgwXVag5Z3dQg9KRO3ZEzX
hiumrM+UlkDro5Qb1scRtWxYWIHx9bGP7eqgpFnTJzUzrpOLkfxSTFP/n2mJvY/0
lRKUzfZfOUaU+z6HTPV3Yukqp1wNKzUrgiu9eTqaIglhLR+01PB41fxSz0Kgo+ux
PJe3ihSAABH/tHHzZk6Un5TXM6Gi375jaDy7+ABOHVrbr38nARFFMy4jmEH2PUgg
KCzHSzex+EZ24UexGgUqojjE8eQyLNLfM6Vux+ra+LQWwIJVX5MZgRVF5Gmv5lzs
uPMNoOP1g03YtbqpekP8Ed50OFG2FvCA4Icmet8c9x5O6OZoqmALXJXC29Sh6v38
zGetkaXtuk8CAxfXOhYAYc0Wsi6iuwcDEVqcKDTMPlFiBS3NjYlslrU/405nqCU0
cX/e+eW8KQ8wdFVJdU9muKbP5jRhp36m9zSv5xuuqTKKNC3HXrWe2oSqtCtgXYyW
XQic+vU4EX7XVNT9c/Nm9/hBmrCrsOHn3cUvQvmI9nWsriaVhc9ghSSWehwX4/zy
Mk2ZepzFvFp3XALgFHx5duphxcPMX4EOB06SUYGQZziabT3ErhbacZTW38OqL8PI
XQPzi5sW0pCFtFTYREcacWCy7cxfn8H14VnO1/g3ZczNBha2lV98Mej0hGCvy137
nTwUBPgDOoym43ej6LwYExCSwB8jVeSsVxhsMK53tHldOMCW50487S9HMIrZ5VC3
0Yrn+YyOh8oyfAX1q6IBgN2/ab4di6CMq0wtPT8Dm5CT/K9+hmJVMYdY4/tUtCPH
8KwzjiDGJzZkUJkpE/n0ismUHpclX0YzSL3pUckF4tr78wbs/Q7oCp5hZXi3AIUM
myiSQFExpXAMMh1im6g9AwvRNuGqEfzMo89SkSparkCGwEvthHaxmeNbool864ic
qahVlT61ec05NNmQvJerrRqgTrf6711Hp/6xXqiWfnkuxooGrrQ+YVsPC9Yd8TQg
fwnNtjMF3Kh7ldh5O4lR1Fx8/QD08bNGyT9IyZusWhOxSXgYXPniwbNs9F1LmTm1
5qbxsTzk9Uyv6TyPFA3P21wuG6LXisUD4lSzh0rjK4V4NNslf1EsEJHZ2mSOITFg
MOlzubaIO/ooVmJ681M71RtG8WzWQD1Up/boBXkrZYFErmyCyGg2tyMniNRn27s5
UpzcuAbaXXBbKMyQRzyv0SiCjkQnzQ15XUu4Evy7QiV2YBGC2WsonCHWHHuqUqKs
rTKo5RuyvoyfbQk3FYWDo68CAUKqs9BPehuwqE5ANXH8QxIcR5GUExa4xPeH86g2
8iHz6KLOH5WT7wpf1cvW+Bo2wllGbdfJ7LVjE1cmHwBYbiJfnVB1UDeIhotHIhU6
BezpsyLdmHnvsjXF/9A9Jj7Dus0AlsmrDtXW64MEwWob059NgNK1lUVom/J/7Oxl
G/khOYtQazhhhtJ+JiaxVTYlYGuILgjDZPE2421Tk9d9yBxmx21Kq59Mp3c30XkF
fOQrZszmPKjngyW5tKBWg/jis2oiaRa6ZCJGwJFciE1ZkSQvOk/1F4WFN9spd9k3
X+TjXabtThOqY9jVnXnzi/08gZ1p7A0LisMlQgQcTUR/Dtf88ALvQ97GOlfPZHaG
glVmfISve9HQvVTV0hITXyE2X74f1nfRO+xXKXsDtN2UM8bPeFPxjszcBDcDUcZG
ZOp8YdbQJOyDU28JjLLyp/mNRKWUTgRlOGEb/FRXdoW6OChDHdkiEEKPu1jxgpD9
oXSCm84Haa98C/utARX3uhioRv9BaGrU6UZnFzuoYoEd14iJtV6fC4A4NBWxNU5n
VyLF7cpYbGpZQ1mXhnpfNgriiUohr4a1UfaPRrhjHOIxFm4dOxp/94y6WzpGpQDR
ZcCkdhZ9dKxpcIvvpqMTHagisfwfQQ1LRRMegCL4tE/VeoIFDAtv+kswT/yi9QEO
upljfqZv4j+FJ1D+W7H/3gDNXQsAj6y2DW0muS5gN6MNGJQmP8rJQ+ARmRXO8CJ5
vzMB5ks6j87Ofy+ZRsQPlOgn/jbW/vsV5XKOwB9br+1+GFiJuK8fIDfMxbJq3AlK
iyXhSgRVutRESC6weCgDud4RSBJwAVHfiKNsWzNF493SnLpFOYxSOVMniLT3XeiK
URPUoV3d3HrDrW2W+XKCebZHqqDyvGA/nikrX88TU+bjJ/M5iRLg8tBoemTdkwQo
itHgdwdiZaK1ww/4sQd85AsH84x2gEsUqQIBEo9FLYcULVgHfQrtkeMTudYbZGbX
MlDHHLWsYacGotSdJe9XBR+Su/2RN3p/2IcOCDFCIgQZ8G3snF+NgDO2k0RaVkga
OAuyTgXDAlJKGQiXKnkD520js5nPzYUMXP+sF0qpXNrxyJmKDcL18tnHvgrX00Pa
INY73xt09muvuSp2L+qgaF+xWBWX/5ASmtIBG7tKl26VnC+zyIU1bsuS/29Z+Rgj
WgWUe7ZTyEDQEnNnf62XDrv/gIAf9KKyFFJ5NuvhNPFxb+5BoDCRTAVHF4Gy3oal
90G9b1newmsxSWx603z0lb9MLGkEDEViw/Rpxo5usczq2hDgsVHRDyX8rydFekPo
qcVTGFlV50Gqjg8bFRbBt6d9q5eZcD1kpXnYqoHLD5R9AEpNKz2k1NaWIDgdHDcZ
H2n6HS3WjUKbo10jQqrBWxzDpSEx2RYuE9WLZN3uIy4VcNdj5kfuNqR5eELBmGbi
DUpxYC97X/bfN68k6zkpHCD3XBl2utcHIU6NXPMXZn+wWbSbdJMEUXWlOsh38ONZ
jbFgkJNgMSOiGGkKRjxprgAOXs7XU8DeUO5fvMX+994zFYppp8bP0Hx61nXOGY1K
4D6OG0vm7AbaWamkGJqlHvvQymvGgobJGM2u5dPVD2RzD4ag/+DcRf8zwvP+rNsZ
AIjiBB03Mf/nfWdZMVy9SRcAilxA17V7HU1JeNZogzDkjXSZpwW2JTcB/t4B6W60
07Q81xwTE8nm/nm2znICSOMFSRCwnh/RXOibgFUAcckeJdplf5V6rdQVEPfpsjfh
iTowXMkKvShB9+09a2bA/AchjhqmbQKs79GorPuk1MnbCEVnfMDgQoHRLQ/GA0nV
n2bc8n9IS/UnaGSCcmTawmw6CS9lqEUoSlC6i/lexPMIznGgCx+ox3zKOAQUFF5Y
MOCUcGrfZaQdot5LaKRxQvr1LtN19hKLnKfQ5eezs+cn/cUhUXeyjIDwY3nnKrpT
aFslW6XzNaaRShvHnf4ivrjqyXN1UsDTd4Zk1Raq1uBKl6kETnP/Hrn2zqsJOi9C
n11MbaEFWVgIspXJU2+02saffJ82x3gVibTvBsWt1Dv4u5lyH9g5bJciX0M7Y2Ks
gNd02w30gq4bLRdDNjR1gYhehPISqBfOnfAgPhvBfS2YUZRUSyKGh6adsxEgJpkm
NqvM0P3jI657bY4uLAagKYECjIg2mD+n8Rfk/Mc8YY/GK2/5NR+KYCbpkVPJKr0x
ZSUjGCA8ms0aztJoko3sKFArbifPvC0adpVZCAEdCEx7xlz/dgrP6gyzw84BvUZM
51ePFmyqVGiFB0H/QOUjYN1VfSOT1aIRAqj8TtDpeqYteiYVCuciGeQTnc6Ezclx
m4FRcWz2kW5cnm1EaVTJMHHnsKKU5WxPc3jqJGZr4/gl+Cup0RieM4wQnNW6s2Lf
mYjnp6TT8nyCgKa2l5/GL0WcgkZrTeedfC85qCXd6ThC2kYkGPamHphK8Y2Xq6oV
odtV/hZjKbdAIQWgq0xBqIQfYXZcTmyAq90bNBTJBzAlk05ybf9yuSHgVlhYYpYq
VwgUG99mtWfrdf6gj/1LJuX2yvY3Z22OaNizvHe6PproVco0p7UjNs6qpLwqOD08
rPtS1+cGKFZaTfZfDWN0kcdcQBHu3ZdWq/W3dERvJMaQhI7/ykB5mX7cqx0VgDFQ
3KD2NWmiFTOBVPog2EH97/1JzCJZ425DodyFH33ghwkRFjD9cNS0TBYfIQWVNNCW
52MLnRKkDswa5VfYzY8wFb7RESm4Ea4UbDbGmFbiVsQamzHVtdkAUf0Hsj3eAcOC
cDLnVAEMs1OUkxX1+kCONtocaX0z8eSF5ntyC6xBdZg7p+RaNwP06w12JqH/Iu2U
DK0IMF+KV6O3Pg0tWykEW7b3E9P47q+2ZvgHVV2ubfla/mbFmyYLDjdJUojZAiOC
pr93d+6ME4IGFGPxG3zVfEWq8BEL1m8VQ7BWJx/d3XmSeF/bZic7BDvURCP4uwu9
eLRVIKk0yH4O4Ns96ADyZjsQ7et1aS8aaFuSqMcxwFDAvzKlr5aYvx3/fldHtENW
GDRDlprZe5AnPLNG0HuzHnjmRo2yBUtFlI6fYK16wWblgnKogJkxKSMzq8NcaKfK
odVslcWcbLXkYVe2x03Xy0OYtVltTDC1idr74HugyvEZWBU3NjiWlsEqXWYqmxTl
iCP9r7WyI6QGJuMnr/6T7K22yPNGvyKySoPzzRqGIWDhopyne9abtXWXd/JTVMLE
fZvlBAsqzyVk6PzRGKWFkk55lVnNxPa1N49mxCcReBqEqkx5gaIkQFDUx4Z0zm1g
mhn4NTc2ksdl1fKBo5Fi4ZpagmOBFnRzEXwBLHht03ZBblWtfu0vZv7phop7Ozfn
B490v108ivq5y+nxH71gvqj5fY1q9OkeqqLIWph5MWcmrYQEicIymLyhEFZdC4Cn
NgPA0zRmND9Sr/1Z3gqlrgMGxiMD6EdCFcXo6NEAcndaRTvkCt6GBhzSR0VBXFKa
SHTwQaDqs0jBCCGMo8t3VdDkpk1AmvdqTUDL8+ncVnUkpcZeJQnAn9UauFYamPfx
MJJkae63c40OCS0EvIrVeBkxvZy+yzyMeixt5HaysjGuQeTGXT3n1hPERaZdTk43
qiue6NXfAcXTRTWwMlj71+9wXh1TiML9Zp2dEPsfYIbFbEn5LqiCccc37TzjAzb2
8Eb7aUmsv3Mn+US6WjvgvdmXJD4R5bjvFnXTyQl6xjL3f1jFMywa6hwk99hs+qVo
pdsG6bCNKyaC1QgE/QDQ2wInar/1yJGE1SYy/C3isUeePm0dxonHyimlAdfW30YU
h+C6JA8coCEOgLuGk71F3Ie+vyNydQCQyT1cKo/Q50ZJW95q+R2z/jKatLlKCdcG
IryCoh01610dy55Fzc+ygDUhUn9iBGk0rKRsQHRYf3bIomicBJL8lVOwL3JkdiOZ
O46Nwtu284Que/a0n5zgFKT0f+xECUXvakQkAfAJtnXCBIrwsnhNvQvVu649QvMZ
ZzHF3jZRjcz1Xe+n4ZrSdnR9ZSEIN+tzLLNscLyh/sAjTbtOFY9WGQzW7qqqFP14
EzVAQTpTnMVAen+eFIx8HS7FDk+zTA1MqRDAW7g3dDbe8SvWx64J7brR8h6oPC17
IWMjMSPK5oY78LUCgKFKP4Pox6/5ztFf4orgjBd4QvAPn0m6j/bjXbhxhHxnY6VA
vMqnU7SWc41Ze6tpWzqZzuDmdy3etnMIDHRvB4EJrRtYTWO7OR0OQ07eMdbL8cb3
SKhaQF14oMMtK3XXNLsXkcejfbqn96fnrGv/S7Z1MBhIAWnd+VWt6wvYFHRwkqrf
QlatWyfhKqdPurQZb8jggla8ByAkxA7jcQ4j7fzumGf1w+eZulyJ1bxEG9N6rnoM
4BOEJPJKj+xMGIFPF+9iy3i10/6YeB3NGY3yoLMQDDbG6sRe0NJ/Ph0O9BX/OBUx
2pQzvXDeTi8IGZfUdiQ1dXrrgEF/S7LpI4ZKrCPEEAUp12JXI6VbhRIwr1HmElKo
83mB2910EIINzz67riqhkQDNnE/TuYFvdxu3gQpB2SgtT941xUDt0bdaYshE7Qzb
JNiW3/1BlzYX5G4IyFq8/Fvnz7v/2hC2/iHoEPaJASz5BnXuU8+3B8z9bGsiA9NE
IDGFO5dSpRR6mFP4wl2YYJ8VnS46Yz6ljA4MiW+TnZVxBQzeq7kfPkX/+V6vW6S2
cyySBXW0L4hrzAkwl7yi+CPOPtCB3Tk6CmP6eTTwzN7ileqWK+i59YG2nplYZmZm
5+8WhnCmZFeM0409n3eg75WlBJsX3yS5drcvZYmHxEOw38DfCtn982BV284gNPtM
24vOnYIDJG97q1BeJ1usAAMsdkqlcySIkByPOeruu1eEPUT8K1TgEfVjj2ocOe/e
6F6mfAH1lH/COWdWOAOYIzsAeaeI71rx/T/zLqPZCCwZVwZcO6WUEZQ0Ukl3Noj6
aqUhvULcUEDq8b/NuRraKk4iaZpBnF7W3wFrCD75HPVYPeJHDKEklKFsfsNbiwhV
qaycBRtve/HhKn+4x+Bmx0y2BUEQiUQiYSq1JsAYQAyW9WJH9AZ5u5q6xuPLWeTZ
mZyXdfh9VX/2k4/aKEXBRulIPFcu4FXzIXe+/168e2Ubms3LTheb+1oHNG70k/ph
Pl04uigHMQQ84rUc6flM2sROqfoXsBT3JNj3IbtiMqI60VvJjJhXivWoEg1onDH1
c57n65WJV/e1OLEtZSUL6c57eOn+PhIYmA2Ib4tpR0bchz0mUz5UknHevCzp/Yhb
VrJThXFl5sh8GWLzyEMF9PRZKrazL5haK9ZjzmriKbvKu02FbALgREgqxITi3I1Q
AjylPX4Hj2/ihQruD+EcNkCoaMLFTC/cKdFzssuHJu76JcVNMoTm+2IsikPwh92N
+OvjtzF5nXsuOM7Hy3Q16oV1cfhpCgW+cWoSIbVA1HScHdEIGv/BpLeDOvuVM49a
Zo30pijB3F0XlKdVB8YNHOMiZpR4edy74SkM63SX0z8Y9uhCX6xbp9gjTW6AJyJg
Hn85MfuZYyD2ZhiLxqiqnQF5ZCpUNrJgKnZB3wiD9Y9tv2UkI8Vu/0idqqMD0coj
4g2vy3fKzBIV3KRD5DR5zbcGEqEdH9KBw1OT1FoC7vKDS/YWG/sBsq9amdvRbO77
w1BPwoYDAx0R2w41+G1omjGH3NgopIp0k8Xu753WIyPpaHNONpJvPHiJ1LynBmME
+FlMOfDUXb/Lce3sUS07BDI0yYDXpPi3bqKFlWoD0DlL7jdlDiMh7KROGOvqQoyb
8LTwarqvnBiOwDM4nn2TAg5Q/ml/1Jrpamui9wjs5IGQp+0SNtne9xWDIHzDDvfH
val+F+1t8VpTXNQDn+wiV8QRmwQHTgn6JU5SK/OfUnO2sN8dh1CPdfixkOyK2TQ0
Gx0b6jnIF5AMNr9N0zYsLdW5YIvNv6SLl2KE6AVCAvG9fk6GE4wOiARIwGVMoBLl
7Fng99ifWb2Rbveno9bFiu8tFcEsmT5T3dpOfC/+xvW6TG5Bo+GSIb3+VZWHSLB9
02R8t4vV76L1qXfmRlLa5ld4f1Yi1xuK9t6ZJ6vgRtJtSIxKDux8g34KbkfXSZHR
sSzFifx3I9e46Vq6rmOl/RMypShzk+6WKshWmrbkGEPP5l6+cuCF3QqYlnJLq6Bf
kZclaXc9UVvs7DlOTlshFJS1r19fNN84r9id+e5SnT4/X5I9L4croafXTKWMFrJu
ukr+GdRHjr8MJpJ73e9RVn2ho++NXRsteedzV6Gk5sNSrZfk6wsOhGX0yYwGKcjt
V8NOLcjsFtU/EGB0i9zyAr1/CXQDatC92gaoGFWoC7AvRYZ5hQ4XilIEOS0Gwy/h
HC5019IbMTWLfELpn/kMUttGg3uMj7P9PvdcBrxzOQ0eTCsMQW/F8BZAQE0dpaXQ
p3FVNBgDqU8rf21Zwxae/uh5nlJrnq8UE1CnQ8oZnFxPfY/Tdgt5M3w/PorkzVWQ
O4Dxt+Rk4Ce9kgGiEebFo6hhaZQyzXA00M+RdrUoE0P8q5zVoE2ETV+bpeFO9nVp
JF7YL4ZVkGHxCHFD+Gx+qumGcMuyh265ZtX4zy3gYov8H9ty8cj+FhMtLUZdnLVb
yXudHv+dIfB+vbpGKj4EieDnZKsxMO0l32WIpddLUcX7WzwmKzzpdsxyQKq02Sjz
U4QWA4wAWTjUy/kLMTnRxPxTgrlucq11dKVB5/cLS315suwUdT8PsbeIGM1GgKXt
MeFswf1QOcp7+s4xA0pgMgmy8ofOAkn2sCbw21wojZwEd1Svpa7nxz8QXWs9GB9E
pALx8SWXeEaxIO4DaXsRDbIiejnyc7mr8xKok3hh7HFKIQtElKCP51sCssuML3Ms
X2OUanPkjDdPY76Ou6z/Ftv8DYSXfVdgzG1I3zzHSeqX2QbHvmx5sUkE9eZcf91r
sc7HyzcPQkJPzI4PlL3QNBaw6bYEiBdkL4PIfYShuAPWQDSfwUOZJYZcD+khRjly
UUPoZQ021Ss+M+OrHdQCihkPegFOdwiDDcejfsfXHn+V6Tg3vaNlggMc/U7M9dLC
8BWzNcvADKAmunzCO/J5/WSkdQlLhVJR/ZP/7c8wVW322mjjO100ynu2UYDdv3nP
7fVhd2ob6YJvV1J2ekTxEBFc362o9ucoTHY7fFpL4xZn8gXQR+vt1ZxuUIGyITUZ
4CJ6L4N/+nAqzYxKaV8Pw5dxspIaBNR8KqOGjb+1dwqyZ3CZl4Lv6YuxhZ6Io/UR
+F6eHk3OyZ0hCBLB54+afA8JfbLTLKST5Zv7erFi8U1Knbu/mMv4knjA/O+Fg8A9
pkfPc/405t2qh6ZU+Qdl4bgFRL5JZrdl1Cn5W4CBPFWbVT1Oosw6KoEGF6pNsnHF
2En3Pm0V4Od8LVKHHH0wNdOkuYBvqbw5LcBiWriVmwgGnwbzAU+mAyekpbdtAtWX
1WeYopM0F3ziBtMGD9oFQEW0+56xgYMMPs2Qn9dCFUnpEd0F7BVnpSXtoK+CI7BH
JY7oH8rZqgpq3JD2ngMKI0RWOuHfidSgaX0I6vUSm20o5ojPsULtVlTQ+g16euuQ
qDRF+xplYzXgJDvh3OT4aKbAX68K6ExRvHjM42vB+pVWInqpywVyv1gH7pGGZokq
l4ICSuh3yyR4osnQ3oLz86Bw2lnczEcAmvyEmv/8dxhPsXGSnSoImE618hHLJr/1
dnPvT0rs7UDJKkmMYBsFVxojlY5m+kO1JriZquBBM5Gmj/989OdlcBjrSfUpv52n
zV60z8tTMk4yLxYOLyxvyjUfkLds5GBF8OpiwRl/oJR+3qYecva+AYNrlWh50ZrN
biYhvY/I+pfwRC+vYC4sG9tFIoLeO04OAHDtIz8+A3rVmzp769HT4Foj0hq9djm+
v8taFgnPohkiQwaa8BEYcR9HMuFNaYc3WgRIU3943sCaWsYDjITlNr7kkOtKVxvW
f8P6Zuc8TcKeB36+Ll/y/LqTDP1YoGMPJUnP8U7LRn7TdngaRaXJtPwZH3H1l8F7
hDzCbOGrZ5JyI+W8HiqmX20hG2JYmpMlnH+wpPxw7GOI56vglK4aXT3y5aCUw8Jg
wNHXdOOBcmsqj5Yu2WHt/MvXpNbjPtYoF+rzBnhj8PbzJ+hAyMc90XGJm7QqK7Rl
pLzzHulgyGIT2bhR6ntRfrH0yUAMW76Umt85kOhvQwUgbYn3mfrI2Wj9TNzAJHd/
vfR6qeO3D1QkNDblA0wHHoIvsnK4Y7B+RPeKxNQPu9zJdoO4RLe8GE20RfHu8SSt
5Xh1UVtVQ2p1YFHf4x4d0ty1PFPBHMPJHGK3RmRQttMz6Yf2bmvfl4gn821yc/VH
oMnhrlWk9RwZYw6JFijpvlA4rg7RB+t5TATZuB6dj363xUq0Sq3lHl1zhVIqv0QB
Twom7D0jJBEiy1xnF96avm3rtCykwjiMouWMAVAEwRbf1b12fhQJPwy9Mnni5G+L
QMTI4VFHUO6UT9+evFkswJzpIAiDrPzgP6l128MjB+2YIQmrLL0Td75jLOkFqo7C
AEKIA9NxnjwtL1IdtM8/upr5py6F4VcPB+QwplXeIvf/KUEN2uzVvOn8SXX6p2HJ
KuQ5VNN8TEpkNjh8iRtqHcg86/EHdwzZHNiZQJVNWgw/8nvVgbkS6P3lUfIUE8E1
qT4s1YPzmOJgWHAosfAdr1tclcmQFzciWLxLOMSdj5Hkx8hSJ7fVkqsKiWwwc+Dz
/eWWq8XatTsm7YnUz4KHV2Vtyl8+yaZIJMJNVcL96RNIbkDshGEGZfOfUK/v0Ibw
DPHOtx9MlM69txTiWNsSRn8e84UeMqBpHakqkwB5F6f8GiAOWpZUqLf/X3o4QztP
gDvtJHxa8K9JYsJ6arSGncXg1n8xOrMgJX4H3XlAbHAm7so9XbE5TfUED/SpLRR7
MW6Tfck0Ap4XiMrZ4grDlvP09MXGo7VgwYJMYAn9rWjpSQvl2DRnMN6vwy9PQ9gJ
ev3SLK/BRUBzfAC7yvzWkcOPvWbFK3Dx1l0TaJ7kTEvL4LJZfN9B9pULTZoQkQ0K
6QBcXXCEa7Dlo4SBt5Bejphjj6mxOTtn+vapXPJYb4MUuQSMR46CFS3lhpE16C8l
ajDGT/qvEWTvjNkmwwx+13SU2DCV9hZeuGmWwOC5r2OS48rsEu5V9GM/6aqehgj7
IotBUh8VuMywdbdIV/SPfO4SetgmstlDC7JLPdNlhCdKi29Gd2bPfTUurIyPtUL9
4+tb23lQ5CPzP99H4vsfELAFItWveOqsPwhfK7CfRvta1NVPV5m9G+2VWrjfnEZs
vrqidqfW7V9eXPbFc4wAHlypjmwKyw1jCtg7iE1XpO4/7O9wzb8BQ4d2YWiE5LBe
VwtDBY2ImnNC7zIDySnyp6CsknDtm2Aoxj77MS//M0L45IicBjfSGg2jxdppjMTo
TFqQg7a62W2iqYBuwcpl1Me7J6NCzKHnDmIoVUmRx/5+FK6tkNUXgUnQKupItpYC
cZJnhOsWCTH0fc7UE9KGkpQme6JW9gczR4HiW5uWWCUnmydxsqPU60Hop/buemwW
Lnw5ng74PuXV2jp/ia4pw/SlMK4STHqlL7I59lwJEEjiO9fKZUrw+djKA3RNeVJN
6PegcvnHv8at9PWVlW38+HPxeJrH8K7U51PAvPf2CEMyr4x3OpGIfx5ycc55nmG2
HyU66z2k91o3HyXScNyDyLjvPhh15R+dur9BOfqK1GtlNJ+4BOr+fbFvXeHChVnP
VMr/BMIXHgKbqW6ZYPXa12stSM37g9q0WC6RThYQEJT1TGpHzqXWzemK+a5pCkqM
csVJLwuuCZoF42AOkV1sULPKFX7N5uMftkD9bK8XmxevuAcHg1YDN46dPELCutfZ
/SV6Vj4mu7AvPjwpmCOTpScSs4skkxdnrppgvCTpUEkvOzUojjyMm8kxNCLqoBWc
FUV2Zfr0PQHi7j2UQxvTnB0+58KKcewzoMX/lZe9YZwcLNokRS764QZ9kWLY5hjn
hXv+82GlEDwSSj2wHtndGVYc40HO4KWGS1ABBIq6oCiKTR/v7fiFdjjn6LWtvryF
uWVdhuJyvqyc5tl6IsXphmE/poo4N+Eb5kzEL8c/9oC5eYVN+yjx75qvAgjvG7rb
FK5hINYxsQazjhtpQpDOLZ/PfRc/oTHNv1KepEsclikfRGue7bXrnzHXqgvoQqzm
kOsZZ0+YvQ2htLZAuV7Qg+VkMCqG57jtuGCsS6FkJ+PCUMG5mTw7YXobs0kErWf8
VkDXe9e/jKUhxt0mhvge8QPUgPW9ngF2fM+sXWSlM4So/nwEQtOBQr4IavFHq1Vu
a3Dvw9Efq5/dTWtj+FfSBrrU2f/R9zN7sA73iXuNWq7NBWiO3naeq/30bEcCOuxH
eigJSSx6ZSCOjjZawCtdDo5WNr8lcIkrCWu3uAfdJ5sei1Dz3FBf7t8bKiA1wk6/
3cLUkyHzl5RRq34abOb4D2Oboy2xxxVcEvv0TDXlGpGOb3AzCOxB3jgTks0nwkxi
VTO1SZ659QxaoHtpYCnt4HhNM5GpoPFcGJb0RA1ordlbNLRCRM6l2p9UBc0rsWZL
Pre4Yb5sARJpaJNx1nCORAanE7feKhXlzRZixWZ3mKhSY2fxe5jDxiRnb2qfCNIv
p4hR8JEKL/AhtQPFXO+wbBHgHnAvaPP9I9wZ43yKkfY8qQ19AkpPhjcjIhRufwdh
GwUsxwkL9amu1bMTpt4TPmuNr4Z1lHdi7Qyl5KDZ4yuvk4KO/AQKTAfDNFkiy2uJ
flwP9MOa2TzOWvHD6KihEs7PTdmE75ic2j55SnpgeK/5hb/Gqirpedy8n3vtO0xQ
W6QM+4PSgwqfNK6RAZaj3lq+09UBf3KKPiRtsOhbwevD4J6Cgrv+MKC93FXQshJX
4qXfKOfsKGTjeDQs64TEg+ludmlMyGm+wFGxQ9GYHEtM9s/WJk7GBEGiaRZ/6cGp
7UcICe1orSVZla0k88bwig6p25NJpRU/Vnal7uJMbCSZk3opV1pxbWKquNovEDb/
XqeggRIkkooRNMxoxmsKAe8L8+99USdDPWm4IWqm0W6a1gQW1MjrefQ/ivtw/cYZ
gkxeFinSDRxVSMtmzXXzMdOyFTyDhv5/WvclNMAsFmDHVXUksC/XP6A3XSOAQ+hY
GRX1lUT7bRWYaPM1MNBt97dPGsMQk3fh2YxRvwJRczd+rCwPCjQqoVWz19GL5WcF
FZ2YPUwnLzRw7QiccrjOREEL4+cN6HBEErSK3lRo1QPeppi7K75M2AFIhwBsS9jU
92RoAx+wdC6lNuxsQkxJzeNmModCnwlDHVqkTFcr1gvUwlz1s2Tb9NLd2JcyPTly
ZcwIe3ASVbnCOcgPA3jYQU86sCRtlyuyZBNUmmMJIxb1mYW3uMtDMXHibRcZ1qAh
VIteJKyZijDyp3wLnpouswN4Akhbs7WSErl4FVLEva/E2hX5+q7ZWWfpDf4T35JO
UaqobYU7E5bkDFRQSp+JECrsbcTJRJRIpdbAfU734nySJD7xYDJFswDcRpW1LgX9
VYmH35QrfkhztKXlc1J8X97TIpAWN0rYNRBhrdMpyV9qwIRRF1MMJ24R5ki1aPi7
/hgMJfWGccQcvBQnO280WFJ5Oreqkc6G8098VqHbbhRcjtme2IWeo0Z9RHqxl43L
F2NbD1qnPe6eW3h3xMQDFL/z9MjYXVKI+yaoA57cIJqFE/nBJGXPP7eDy6PIHL2b
AIxD+9IjkP9HZkz37jEKQZBYLMwDu9oasnHjwQd8TzgzcMTqxjndqDF6QWpaceJ+
dtaQWI/PZp7k1H83Lh1SjVGHizKbB8/Srhr7+hF8UzcpKyI6M99enH3sKxrPz4Ta
OHKkCqUXD53HE9eb4BvFiPYrzcL049mSBq8k4QBQpM4XbP1j+g/lfvlTgOJFyn7m
XU2YhfyvffIdqn2ZI3NLCGsdb2Rf7wSFDOPKU7I0mMYbuG0jMMD3+XBuFiq0P+2Z
PxKXoYYq/3O1/cxyJMYXB5zXUsUF778TlL9R7+0GETbNrgK4KKYCBXt8HARDua1Y
VPBNt+E++pFeRNxHR7eclO5pZStvVBKWUnbnalwXBkPFl7ZXYG1+tDygnyByo++4
0/tBSTbOl7sve/JCve0h7ZYiaM9dRiYuHXo9d06UA/uB0/KPdsfVc9JcUk8ExyVb
6wvtIgtdcag30O+4883uop3y2vAFjYH9dU3ITw0hDh9tMTaO8Gwe0q8cfxPPcJSE
BHRkw4z13xyzD8s/MjkGxKZ3kP+M4CtB8Qvb9qYqzF1hM/FMPRCMEfEN6fpblDEu
XCEBdOonE1nmMOqiKrBjsxP4MhEjjcTbymsSA+SDDlxGF4qFClpm7UeEFBaY/vHF
HFrX+6TPvIXRTjhweBi9TAgpbDuNLCfD2LkwpSvsr1LmVfzwsHyZnuDhWL4gF4U4
qoEPkaIZrkNTXnlcYWQpLb5SvB4UhVHfkhSdJvzEhklPXkCR3i5UIcvpJNuQlVIH
NWoRFkrcAdIhqxpxpAhq99e8hFWt5yB2qVselDYpROLv4DWZRe1Ia0zh5nibp379
ImpY1KeJ4jdPKfE8PNJMQhE+kQUDTAgxyl5b/MMxOQ0zfabElSWeCI777U34GAIy
`protect END_PROTECTED