-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
wNQHIy9ugBo7iQoguWjY0m8DJVVOfuDIZFEh7yw4VLyng3jgLa++vtGJ42tpA7yl
FgLGDee8M1kpgtYYr4QEwUYYJ7lWS8kRy1T2RvE4bJOnIAjczK+XoV9vXxYjR2W6
i2k9m9fdfMHdYgTB7zggt90mwZ9iQOWNhcLS5FSEXyynNrqa75agqg==
--pragma protect end_key_block
--pragma protect digest_block
ZhTokptSF0XC/YuYem6J79gWQpU=
--pragma protect end_digest_block
--pragma protect data_block
YIx4VRt4kuGhL/DnBVELfMo+pBd4lX0LpEkL+hip/TwA0RiujHggtCT4gvAmZnqF
/wlWGrWHo/7PO3t4B2XxhsogeqI1Gg5+PkQBCnwDAAXkKphqoshY7e3p9ChtGMZh
M9k+WlGQcxe9N9qWA/kD2NQhJQD/NEGVuVtY3XFp2rFU64263o+0xYZbYchpCMfn
Xs4erUstqfah1EHVqvKP/RoWLVGmLo7+xfWXB/PQyjbrqE1yxoHGv1cxOILJOabF
ze+DKUCoa7/6x/90J/UKQAC11gRXd5J6aispoToc/XuMo2vQ+6mk4Svu74gY1itg
x537bpurUtRcr8zBeN+1ZAp59zH8PE+97VO3exWNaKJca8Op0kg86UHA7SJMFTZZ
SNaZuK/01oNHC4z79Kt6GgmWzJe0Y2mViVPoW443wikF45xD5ii1glCJCXmpgGLF
IqrcRSyIntFdg6xMtDeZyNt4b3mZ+Qzi15sqMGDK2TQcCwF5ZZpTuGRZ+jwuuJi2
Lmc69edGIMuK9Jjn8JEPt/R/ltsJrjOz0Dl4EtTW5UT4wZrz3ftWCD8lQPXGY6YR
dso7oBsKt5AH7SWWT74V2EfISlqoFpiZEP0kIUqm0wrIrAteolrWXNIHmcwQ1ArZ
llXJgAIYwQ3w9IAT+NGhAFCx/ZyiyNANoixQHw53F6srMbyhss8Zgkk3sxJkE9OR
7boyCj+fnK3yRT5Ic84aESs8RcOhBgJ7TuNhFgVUhMZjvrpVGLDVKKjVW47hd5hB
10HBtgY+E6KxHeyuUxeDGtpeg7r0Gscoq7sTUD5+Hrc+zVBKtDTuJ7oUluGhUMI9
SKqy5VM9/T4/OXXJ9qbN2O0lPILs+xWuc5ehc/MviYOR7lMfCoBtOZIMutGzICdK
Bxnt1Rj+WFEdNs3qCMcbtKOpiejy2rFnaYeCrtLD2irjS2ai2C+J+Wkr9QRlc4Gi
FjTucFO13lYUThD5+C85rllZKcuZMF2MRz2LIXrcbqAlJklbRO34FYd9H0e7ljX4
oy27izGqi+kHTVBkk6IcGCDhYNLw94SGXJQDeNe07CT8mlYG5kIxlvCl1RK0BuJy
X62nXENiTGGDOw0uvY6cPLfpA9m5UaC91ZZj4QvJ6kHIHnCcIdC/AiAFJsZe3ncA
bgVolRePkQwWoMpiTUHqkxoTsWJS+xYY51VxpnvxfzkJwK/aDRW2zX23WcO6oTft
urfiZdRu7yF7BafS+MN0ZKC5C1ESj8vKwXFV2dIyuc6bhCcbdU4QDHCUo0nTnSeZ
ikDzU4DipY7rgJ7qWMEiSfXNFCA9lQj9dTIoDXgOlosCwVJfuH1EVbwX8SUF9eJP
cwV4NuCBpZhomSwAum0WdB5g9Nz8tv+gdF0XYxkyPPPZO7GN2OpjrbdOy+2TUZDs
kvNYx+mhB1o8+8Jr2twTO8x9wdUVN7+k2TYNLiPdFdgBl1E4Z9DjOGC0pFEBBhhY
Xzibh1e+FQQlx215EQG23mISnDm7vcKQ1hsPS7hgylv/TxyOa7yjtCzoLqnnXFr6
dYMG4I3n+AAf1d6M4rbWlahbtB2OL8tBUYGRAh96sCCLXBAptAjFsDj7oDU6nE39
F9T3yuz6VFkZHmDbvtpj5muSb9yTJC+68JGGjRxKw+F86P17zeSk1JRDIaEAKBdR
iukbSK9uxz1fCy+s5o2QTrU2ygPmdKTSEQFLRXTLZ+nJkf9O/rSs0A8mXVYDlN7y
Z1thkDk7ctwZvtbi58GH4Ll4tbuJEuFlbrmtL0HU4i06UC23nmbtdap3ts4M0Ouw
4OytOG/L5RWO3KM9/sk9zSoeuc+LgIP1UuADLjPmF+N5nIt+AX5Xrd3R1mP5m9lw
zgDzuVyvtqOSFpvhzZdVIdsJfbGucRyj8GrCvKyS5gfScOfYAC5I0KtlUPzOeC5l
28TGQyOYxwpNjhyGEJTvqG3Dh3JWol2VDFR+51nuEQfPrEqQwN1Hb1QQZoppGzWU
E3UZHZXLLRV6VDX8rXXv9q1TcssHE/ZrMnhfug63WEp2G1bB/e+Fc0HugV/9FOb6
ruhsypenjI62sS63OjzivRMWKkCgVkEgCFNvhpb03tB0nXxjH3Uapz1IqSOU+SZu
2RMgwXzG4I2KHCzHRXalv6t022Ddh8/JnerhtJNYD9ZrDjqrupc0ij0Wg04gDT/D
ZULZ3198eUgkwGuj0ogvYiUgNp97P1+QpYJb+aWsZhzDJUXGsspQzub/F1JFY3Vo
akJ7dGRHqlvXc49LVc82PgpqI1YszGlDqUdXRBUjHwHoqddP0THHzbxmV5Ib9lh9
gQd8XELgUvetiJnSz4d9svTc5+IaNP9I1sXcDTPLf/MKD5Wzz5nnrP+KbfXq8jXR
SadENArN/ywf8KM7FWE0jb2hhePIkPRoLlukw5VOyFdYZ9D/JNeLkO436XWJdjWA
BLR+ZKFODT6CLlDdhCrdggUT/VV2URr34RySDeCgmp2zPvQN8TLHfYG7A+b/IQlw
hH1bFCxRNFFCitIGdJ071qs2n5YZfF6Uu/0zXYzGV19AM9SoyZrcARBCwMxg5Ksf
h1rza92P7ay+KF3RpRtd23N5t4HQwFnVOU1/bA3y7+adFK7RCojIsrubcFpG7DmB
yy+TOTPXCeBFnpjus2oZfYEZcrz/MrT4ISjZZSu9svwflvw6jMOKgPNa6ETiXJ5S
mDUYMBwmHzn/3bssKfYJUyWJ+25J7oRJA71MGtAWuk9s9LeJeK0PoymjzvszpZLe
WvevOTRpiEQp+68mnHVuuyNoIHbiWuUO+uU22H4fTBftjwbgKnql+CHLx7ZbnUrr
m33wrifE1kTdMlYvdWYyOHpizufxQxuZTAgxKYk7xm+rgA/587133cXA6QK0SljN
A00iho1PWJ5Xg7YZN7SXAsyEnd/u0JPuqa5UwF6WM/kca9JXCy/dMeX1pCDX44l4
wg6dJAV36Db+lk/nQcn18aAtYdCVfSWTZevFKKi3dMCuZ9XQa4AcWLRyag7pVlc8
L72fSOu7HDpZhA5l12gkz/MQDRePRxsXc3z6qF6v9SBwlgquMtt62vY5AuqGH2jb
+cCdF48ghxgI3bG2wX4sc1lgghDJ1L2ZwNPi2JCmsWKFiwi2DA1cPTcfl+XbFW+a
YvY16K3iXyRxwO4bpRXxvsID3cX2zyRvyqKxvNUb5dikmbNJ7UarwbfunQE2l6H2
Ol5CrRCEt6JQ1sJ64zY9xMVV6pXqheNdcridg383Q2pesVWV1paA0quhSxAsdtvB
+8T3FoqNXsoeUjmBsluZgniTk88fktQKEgC7TCO/MC7Igq8r+CKWYL3oRISiGux2
DaM3vMyZm0NQJyNciDE0a9J2CaGfedMlUF9IXuiIn9W75exLoMN9ARHgglqha0a4
piNKoCriylIw0gatksBisc1sBpVTmvP0v01roQuXYxljm16CsBg7QJF9dtvRuLcb
x0lwfUtCGUie8b+FEByO12+phkc11c6Flv868JjClmOpNuRA5UxM+gXAydJwgLwG
yR9cYDirRupr5fTwqVycPG8y4/rx24fdUPwEqB/wQOv6rvHktWkYz3Ng0FFt+uvr
K+bGkdm1l0uePRRI07VCkLnmLMH1j7FylV7/Nb3AmxuFRpHijCC3qlXMocSd5G9y
PlTXtCH4GF6hOzRu1rB4ReAhjVSRCe1aS8K1k+xMICH/h8msuHElUiitA4l9RTWg
1IuqOqgcs6dkAPjwQ+v5io5I9qg9Ms00uJzUV86VpxgEWuuKEhOMTtbnjrDRPT+8
wofy6bcaph532TeuGVHcgr4t2kskZ/VHrNE28i4yN6YVhg81OEZLJQX6iJRDxEuB
UpPrMXMZ+tE1acruhLWCzWNmKfx05KIFhFAq2LqDHN26fUomPqC/ckXwvGL146Mg
NTnpialS3lhNOuykkHZtlMgC+IAtigsw2syFV+V7jnU8tX03YBU+qPhVrpvObzN4
UNrZf5Qlbfg/jT5SkSNLE7+mueVLgSojI0Fua7aKkVWx9XkxqZbRXVgCEE6Euk90
uxJzFBa29zjpB3YpSjgjp068hu01hkszG4j0faB4f6aWBsHejxFCd5C0piraqaY+
xep7CHmrgwpsWy3TsIf+tS6Zr2qhIVnN+BOHWD+4odBaJSddDwAcjXbz8xt52+gs
Y8Q2yc9yHYJKMVZTTRPZValzEm2w6lDthyb1SFtvvyJcsP1Vt07SbwLYF3+btPV4
Kmf4Yd1QMBi8CEX08ZlaGlyhsSR6Z9wM6HfFj/wHJi9mFaB7nMe6SuG/0qq3Vbl6
RfYlppbXD7o+iLCkwRThPW5SHd+dwgKo/4iKDAHlp6LOOBOAqh8bY7tZYKtenKOY
I5YlI3ZMe5GZyqqLAs6UgnvxXXZlmxVCt25jmcQNYKuEPuKDnsZczAjq+AWsG2dM
w7sFgWBSoiTou9/ofcuWI+hWGk0/GnuF0RMahSpm1pz+hms4r07xNs8ol/0odylA
eiiaip97gV1kuJA+FxciiS0QcKNvVMFEQU87NZd1jR0Qpp4zeJ31gmLQuohJ+Bf2
aWXfpLqRKt8Tu3k3qTEhwyI5qjIpdvux2hQ6VHtNG+SAMBVkgOqh6EAUVE+9vVjp
lt5YbeTUSdWe1KcI4G91QFETDDp8q697wR3tocCeXgZ+LnthYLkiL65trMlI9nuS
THAPaW2WLfk6wWJuVPEGesLUejdv4H+WWwXkTAipgJ6vYgRAt7u4k0DJ3+w6TrPU
rSBLGg7m5SAA+i4eTNR/YdPIfwHg2KRndgFrm0y+4vkVUwC20u6xOMBpy/Ci6Fh+
ng6y2E7jAaTYftwVKKTFD/FivmSKYhrVzMQGYP90fH7SCArk53DIVWQa1ac0fB+b
zQMgR3XP6Jo286bR0u2p1TDkF2RVpl6fZ9vxs+u/mxE+2DID/CsenTD9KYXY3QhU
jjea22cShzUAlachLqe3Oz2ppEvRPnphNh7OPPB6+1ifA+ex5IkG8u9JFNEsqC3H
1u9Tclm56G82UgZBi+ZsLl8IijbJZY5r9ZhsFfaKmtIZCGrhxUxS8wXto3olAdN2
1aRCrXoN4N6ODxsjwQm3/2qs7gkQJ4EJintEv6iH5wlCQc/WkGRsizIcCL5YUFQX
678XrxQT7j9EtBtIM14GGMyYGCMdA1Xxy+ZNiaLmNa+A1wXasPEYStd1V92Uux25
065Koo22xSfd1T+rrAAQr4qjUGq8jtc4GczSZWWLRHTO2kRcyu5r3F+fNc/xDWQ4
NdcYed7pZxUzKtSGDEJnSZk9wzYnwo8q0cVBCl3qb54r4DeDH/Dg2h8D9W1kxk1F
m3T35njaJ/KwbabUcs7KBRT7wigvyen9bF5x7rRJAYheYZVkiQZytedzsMDZNelR
iwJp2XTsZrQ8wtg7ieg+w0tDIhEYHm/0tgouJQyepoOGUv4AmkPa7XFhsOBLvCVU
kSj9z3mBrjsrISCDf0OkDpIupTrZDcb042HPSc2YJNiFayTgdnaykY8YFOtAbBxh
j4CpYlDcWrwCGOarc6oW6iyqHyMsKYYptPThjN9L3bu5duz8W6NKCJLGHZDgT45g
xofeVgUdZF5qcseqm4WmIxr+rpWWb3cTe2X5ayHu6xf9jn2VCGLeYpgewmffzgz9
RCT6YwOUqsM4ClMkumfjXNAAHx/YsmYVcvyWmDHVCTEIHg3t0QWm1MicZ938ws8U
JjiKmARyIJV/uUnWSg0mt5q60gPKfttSjymzmIyFT0nBNocqciYokmU5nSjPV7dI
x1YHDPvXZFNXXGajW/9gcAYuwzfssT88avzSqcpO43PHxHw4WFmYsowWeS69aBq3
oz9N/xhAR8elLBze6K+TaFhNolaS2AhHWo4F0osgyWBqQVYCfk9F/wlN/XYNJstH
jX+fMe8YFQHCMvGkMDSMSF/PN3XZAVWtYHAFb/aTJKfh0oXFadzq4irCgZMZFptL
a8j3qC2TsabJ0xi0iUOQnVtX8FqUnOEP0pmSGWO8wZciVuBF0tWZqPR53HK/QVdx
Qodp+1nCpNu/cacaI/mHK0zydvuUT+heXebkLMyjI1fBVVOGP4Jq22J+L8to/fJn
tIzOf0cC8NJtXMs1NqHsQKgjzR9l0rcS+114R+wEdudLCNlBlJyBvemrrwWDFe9I
zY+YaBdyTt4lbKp7DKyAx8ssBERzSTtpUkjRS/l2zy7/XmV3RwcX/7xK82I/a3pm
uGpjYZ4pABZ27x0UVQ5g0nOsrjBWdD56Uo4SocDNw009V5XzEHEvV2e+G48rRC+O
O5vb9u6me4uDKX7S53iCdjQ2Ldt/YZxJ30XqMBSRmqaTQbQLcvNlALzfl/Vqjgni
TXyuJcX5+3TPQhxXV/QekksZKML1zdNRYNtIr/euCCfmic9/xiRenKR9vpWzCQ/i
53lAsWkVlbWgVUaRrpfzLw1qkjTuP7LC0lyd8X0FyoUdcS7pc5T2prfa/xBCI5j/
GVuk6kLH+irhnbS7IIIgv6qpqAPQH63nfFZMUVeK4fFADBUU262ShT9q5CFh1d+4
4zuWRIyVoGy0z475e+s7ceZGylyVaCEF0WVqfaX5tmN+KT7mcnER3WFSdto6/Z/f
k9xxdqYAlf++gg/LdLf2FucDaOZCXf1TOV4pkfWrA/m5s0+FgYrLhSPF9qnvvkMz
vR08DR7okTu6chY4RBVu934lhE1NL/Ft86aGYADeahkfY3SQzI2z9IMsrVx5L+GB
0WuNcAsuCHLYGy5HbogT8VJd62bZL6nkDTCpE4DGFwPTBZb8nESnubq1PT4O4JWA
vt17LWrKE62C5y97flZchyxUy+Xbw6e+JGa3mjz7at2TILL2AbbusVKJVF1ICLj+
kFLUBmMygyVoehdCETjCAImFFrfxuzScJJiqR4Y0lYjAeNDMA8J/P0igZustDJBg
PYlxJF1+3y4GMaEhSeAO84Mn2jBS6kgJciGZpb4l1m0gVc5GdeyxHTez9bO46e/l
8Ykq1LA51JcwXbYXKjXjiJmr7LGkyTgBFJpgkEYMrAeMLBwGElbrJljn2GtXCwvt
P8M3rMtltxWcdxqrru53kt7mAxWVAI3RbE3kzXc7XKfJd6by3TV3LkGokddRL0ZG
EDZyZqmPNHj0qFDrmE8gjR9zscY+fVb+4LNswb7u8OUuydGFsDAQi+N2eU900RDC
H+/iBp7jssfznKTuCvhb0InAgTyZ7OREEK82beFeFDMASFOVSzqwroTdZrlh9gj0
LGLkQg0fqxxL/KOCNJOkuK0eCep/yWAG+b91RF5rMdiAcOeOmHAnkXDHI8Bkdom1
W7DTHRMC8iIJgbHWxjzLycvAmuU3GTNqGGmr1MiCGXMn/Jo3yvDuj1FM3UdR0b1u
V5FPUxGVLjPZfEtuVT6sFRm9LAfae+/Pgbjvcd8Ktvmw5DzzVJO0Y3ewM2hDbgoU
tMc+hl8i56aln+/IiCrj8witHoxtZPKxoBR2F690fDSIRP75IJaRxQiGk37AfKP3
nVxOfe5AuJ2xAAuBGlqyB9zYYcBnzRjRsOayQl2vboFPE+A7WJd4AZGUaZCIvAE4
POqQcFdiFwvMBNzuKNDvZja8vnL+V0xV2mcpNriI/9a9RRAAJMSYWr8WftHQMKCJ
PWgVS8XD51+qKrubeL80o45Bt0WZFyuuK8nYUpbksMSzIsJAAxd34JK8U22kGBpN
Dy+hjEZ9OEcUmJuW3eOZbLJejux+gtWyhWZZhmzONU6RKf5PaFfYWZ3ha1kXZsGg
WOCQmwgx3NgT2dRyKQaVMZlCqQNgCRoSyB28x+Wlcgr8rsAD5exqYmRCUKENQ5sB
nppvjxd10fUj84SgXreXWSvYDVQ/AIVXhYFeHovsvWjtP+BGfS4/+tgX2yEw66gw
g9610XgGQf/LALpdgQAjbM5Me6bhCGaaFgCYZ2qhW+T0paQZ3NF00ZwoEzc1eOg1
y2vhUgSxBJbJmVkIXc+AMWMHlUA9ZNggmmQ+gMwmWz4qkebchRkDY/f92gEBMD2K
UUpqogNwJomJq9sbZqoCuCiRj/LIMRYBjVFQZpu/UJPRPy+SZauyH0COUf6yqqUv
B254z4UbOn5+i8+67kdKB/oUlOD/TPOW3Hl3W1mwbdnLg0PqoJgMdurwlX3ldPGd
3Gzdj+ZNkDVtiZthLmB9mVLjEOmuauMI3+s6/YkVomevPQJbMitkyj/+RZw8u5KT
aRhXQAbAdD3iSp6eWML1iTaoKyMD/ZeO+1t7WyisEggncbbMs5jGrovNjUgnBl0y
hAJzoE60FBnS1qxWnqwCCaLPs1AaABarPwyIVdRuofgrq3rkksty1HuuTiF/ppCV
qsH0hcc3CmJnjb4KJfLIpomwScYWHN5SZmvpuoOYTt7pQaOVz1dzMtXxnAHabYlm
7t+V9dpom/yErI8sQUnwqGi6NVMlrsh+ZWl2Koe4n37o2OTljBqmxxC89b2CrWu2
zT3X3gVKS//MP3tnGGsm2g6z11sNuAbu1SAlOCxF2innXY1QJ/BxxvQ7u8kf12vF
KBfL06uovcnJ/HhaA6HugAX4o338yFeBvJDZJz1GXKcpY+ATxem7moOJ081bzrr5
tqMVOqwoyZi/gqWZrlvWNMRBXUzEmJ9fN+GHe8KmvVysL9b15bJ7iHPdc9ajt/5C
bcwlaTyBSuyEvP5PJdmItK5Zl6ZNc5Xc9wvorhIfJzYK2MMR5A2G8RLsS/4rSRpz
yqn9KQZ/2Z9rH1usaZy33OniUp30PD1ZXZ1EDfDPRp0JH9sN1NbDbqSKtUobwyb9
nBMsdfceKKzFdHuLTrUrVYTBat5WQInQq3hxFnn9UA/LXvppQA1yyrC5Oi7vvy81
B/j1zk+9JI894z56/t4sMTS+m7Dx2J+haqp2RBFc3Stiar2asvBTFAtiit4L1Gqf
F5+y8ObSi0RB/Mb3DcwjLr5f2yK4fkSVSd036DXt2hCS4JLPFIMot7V7sSdNyG30
ovOJZVYkQdgld3YT9hK3jo3w6f1pKVgjYMJ/BKf/3KD7BrgtiBGjF2doPa0fpVkh
PJMDx6nR8e1KO5lLCFWyDpaaROnSPyt7mhMeG95lhUKGGf8Cl8pzR40dvuTAg0T2
RSrwaDBy6fVAOWggYd3+R87g6ZUz0uA/LN16v6SNBeAtRfWHA4Sk/dUwVnruwRXK
uSXvUG3nuwz72Q9hTexg0G8Tp2w30c8GasrXQKPzFZErxCOFdgAyC2SOGoABCklJ
TiCF8iCI6/9iiZJB1hU9sgqVdpJmjFW2fnTza3VSNigLNZokH/lQvOC29ll9CiBK
y63AmB/+cceAwNDDDSqvtgexDNbTsUtdhlrDttZfCvmyjhS+OhrHPS3AdMpGC0e2
W33FQ5R30cvCWzClAummntsh7+wwICBUrzvlgc3Z7S5bIPKGV5Qa/lPnZXA4YGBa
NIe8Ctl4kPYhGRXsUYbNJV+Qxmxp7Y6KYFHCDFGQ5HCsruqWiJVJhPEGLXcRxlF+
ycjxt9YLq8xmc7myVdOZ9tIkLfwQLDMQDSNbE9Q7rdUA51IltahT0K0uBDkLnHb/
0YCLdp8xlbUC+QN1Gs4H2722iBz7RPfe/my1izQSOrQL8+3KincP39Ty9cJWmuHj
32anW14gle7wK34RYm31u1IyjzAGwXCp4YLdSVDeDC7mv+YlE9ebUJnvlyPMlXZz
gfeKsG5eH/Oog+20nj2aruQs3lONWE212YH+COabFTZJ1OHDfHF2LhUwJMoNVB++
RcncTMH7shzc5B5mC6oGxn1uKU1shmVneGb7cWlyZTclhM+BSz8kkrdbpG2tmmWg
BfTFQ3Q/33AS90VZJJOtJPgqyno/2Pc4fbvmK4cvAwhLrab1wdrmIpcDpvVgswcE
ndNfLL4cfEGCEFPzYg+2kiyn45GoZKrYLBWzhueOuqlk7H5SMKAtigU8oLNJg8Yl
wo3onL1r6ayXo/HU/bnF07m0yuqkoEPjVOh36PDmIV9p3n+qckNlrhqZ2Bh0OqDG
WsO1fyq9JjPbgy8A85i0eZFx+7hfBa1yzHLdixvJmauYQrQ9yk7D5V8GqN85mFD7
Yn9BKhXrFkkK/Pi0ptyMJbTHjPzmS1ozTdW9SUyHtWEUvAiH+jqh7SLaCEOW/TXw
0WI+GHKzYlBsQNs53vfhRoGj1z5dp5MsvDBIcsXs6oZrgxOnxEc9mL6i7FZ5zn9S
2cu+n+Z93D9Eq9hLYZIV5j717ptj6Jfr5kuONVdfcNZIKJwPYdBWqUfyiVvJV8fL
qyDSIRfrYYvo9W9smS4eefSBd8D2sw3IfIrgkOohoZtxbpZ91nu2huI6QRmJ8mi5
1ZwWTsEucpYAMHZt1EGNK61auRlkDzKdvXSFL4cHtSVcV54jQVGSZP1DIQEj/sAC
VWu/TCNqzls0WPpTDhm81OPFmwCnAty0QKMdPQuwGrwCICanhsMFDAUzTT6H3oKT
EipvnTRAPAZydPdfwR/xC0bDxkZUBebvm84OKa7xQyj6kYeHMQwvzdBZN86C/wLY
bi8VzoxZ/p3oTjUxC3EEXsIwVIJ6EIoItaOWs7pSLVQ3VY/vDFB9qUTPss0UveQY
6BDhNNfJ/0gcRl0fR7v3EH3H+qMuRokByGJv8+FlZHDpySY0iEj6W+nppteO8C3z
sGMoZRvBeteOa1YpGMIYN31iH/j9FAuvliycnpdWk/3aHzWeICRTa2GVpUnsjtOh
dWgv/XA4QL9wr7auOhmGtjH0AY1QlduJ+BdAim9bnvvw/AcaTtOBJ+eJL3yeL0oK
AJckklglWujnTlGogS2cu9Ient685JUZpca/idkoMDSAKmd3xjs3OpMvuIDpUqpF
QpKE4SRC+/8o/d6P7c747Xb1zEsXyLonO5g4xxSbb0nQjzhHw7G3l1JkXsFVBWkL
QONwfWhWX6YObrXvoFLhyNideXV2Ki2YAN6PEosRoB/0LxXMzIjhoosnNWh2AjAw
zbtC6LDCoOZg8gT6a2QSpFFXUCGisNVbi9Dazan2dujhrhYALcTdelBVZMUTGWBA
3w+T7Rx6VlrdGHaFp4R1qVPCjfj/+t6rbmgwKHV1dx2hm4Kp4Sn268VYgtWg/LJa
+KOaXSQ+I0ksQDvsFEvxWB3seTKbF7U9Gl9CX1ZoDv1CEPz71QxqhHJzRk9L03Ij
JPCPZWlCNw7wQ7TTcpG8qs7goG2Fa1u51Y6fSYSdKV6W1gsNaxNEfLSa2PvhRECj
kzJTbaomGNM2JeaykbTCGvbpB4kTJPP+Prx6SqkXVzdWdzRK+RNmzrX6OtlAYfMw
ZilYsSnHhroEhQJI3Fcb+56+KCf9wD2BRsgdv156D8lAv7EWAQbnwwRrDsNQBeIC
xAIYGDVG2+LHxrZ+OaFV8Na8sr0baksf0zu3CyJaaEmNg2YWVvdauEV74xAq113Y
kmHMshwhG0Vyh7QSHXchXkODFGPtLgrPIWXAC92WYXKiSSt1On8QJeRy+7PM2Eep
IWJ36VPg28AQbNIZ4WbK4CzgJYx1JVVnR5zlOkH3qhb0mj1s09GamyaBKt5v0T5w
zMvNEiXygnOAvpkfavptPgF6u70e7Kz7bNT9L1BpPDfyMqsFAuJuThTG6iBxnSMP
S3Dy5sX4g9PbFdLiGh2GCnlckDVCnTcbQWSvjPfsqRGN6V790k4INEOc9+BHFJVd
ijE4gQvURWYE6xKAyrmiVy/iGyy7IylCi01lfidpe2nGqr1K5HJ/L7Wc9RrCiNN7
y/BnzS+y/arfvcfX3Xb4Gyelm+0+k/2VzC3X2ygC/6IyZUplgUKTRrQco+6qQgAJ
ojiwYiqSVSlLK82OtYcu+DjlkTcEBuxdghCMXJ/9JdGRZJnjH0ZBgadBUIkEII0J
xbekDh17TR80mAybcBNIGAHXzsTOX6RzRyU8m6rsxnZpGi5gfJyQMGKhxp/qW86/
sgEKr2U2nWwppvv/Awc7Nh7LiEwzsWVgouhd/4Fw9b5DA7bCnd509007vntpvKUD
xaSX/m9rO3Vc7D15HsyjMCE58NCKfjPJ/Dzg8cc9zZJj0tdKYqE+z2nzkVcGmlEQ
QU4slEA42ioxJ6Tm4+/iKYpxmf8moZamWWDKPM7BYhxFPoSD4s4Cq+Ri7/jjd82R
pyPn1G7dQo1h5o9pqwO1UPR97CZK43wDS+ifY9oIgiqvCenvQsKguTgSMMiFuMDQ
7R8TZz55tfnxR4mZY7mNPhZAwG9VDz31z/XgSv9ZfPC2qQt6igpaR7Dfrtn63nPe
RZjrH9Mt5ussn+HaJVKogpTMlL/GFTnUJBLdiAMGBt7GwVJ2Lrwql8GMm5DmZguS
KQ/gUIjgd4bSMEZMj52+83FbU89faAkn3qx9tgDNTNB8BqTlEf5usrkZ9bZLNqch
+SLwPNpcHR3BTajj6znDhvBA6uiTOoi+UTRsx91Wu0YsR8DmAVmmLdAFyPC0dDWW
ppyBsn/QvLjj5yami5acPiorJsMtdTA3c04qBz63YGVwvfgtb0ueFyhAlE9YrSZ5
WN6qL7csgItrdVg1uxgP0qwm8BQ5vT4vHczNjkZxYIN954h95anL3uk1FgTDlB7X
coRGhrkB6+jkrA8b5QajNE38oqdA+FJlXXhDyd1gJw3w9bgN3eas+bxruGf6//jf
4oUgP+v83VJTNta1PslbSoILtVYPhaE49KbU5R3NID4dk94lorw68VP2EAvVVLai
YEywn7tDT/xMjYsdOnNdcv4B+K8nv8drZVuc3up9AFOJVCtUn5IhgDqMdclALIdh
jCnkmbQQPBH8BmKZIB1Sq0qRE5nqhrCA2AqT+ownvDhKQkxyJKwkSrh0jueMo3UW
x0pJx+JEvLDQsWwpwguEHKF19Ml8QpViz7xTjhwLFMBjP4TVKcSe6rnyP76JeSZW
vG788j7iPW9HIYIkw8DeGlkdBwYbWvtPxQNDbiyTN/VuX1RSew+iVTYaY64kArit
GSA3mYwJa9Gr+478Ft8xZ1yxzxOXPwH3RRGIC6cRp+7/5WNqn1zxpzILwPLvv7mQ
9gtPNxgckWsBpS7Wwqqto6IzK4mD8EjLk2WlP45iErUV2ABPc1YRzkbN7lIv+T7K
ybzJhpC0iLwLAGdCvHHtFXYAkIlhjWMRH9VrWkOCUyHyFGa9s8gB5oJsgjwgk0I0
aRV+aMnpj0WqVTSczCXOP+MMUTtWvqhHAn3bhprOGAn9IUlPgZtAuMplhtmh9cWI
w98CEsMNlB1ltB4YArLHJQ8HWCUF0aybGREr92Koi+mb7vFxMe0s8AorAbAATYhw
pTXeFlj1uc0i3sODXon7T+BcWOlu8+4pJ3okw67J0GMIh/10Qf5pZgEE/iJU/QOq
6yLJohPFJF7o7NPQcvyIhOnzy/ToaecrPp/chAwkUC49pwe6kjyw8+UosJwuLa/4
4yZvsqYKxtMOydw4Hu8xm/BoJQNT+gYezhTU8n6JCF5SlZgybV7rNc9T+vJ5/U0q
Tst23REKgTdDhZSchSfkv2MK82LGtPYnuK1Pjz8+WZDQv8+t+jyus8Yfiqb/52L7
iM5vD1AIFTSYVmdjbvpvM5ja18PwK6UhylOOBRcaEFYmRdAIXLk5XrojrWYdZH8O
wmi5Um3W6zQjXaRcIFK8fGTHRCgcfnyM/ovjKC/g15mNcJ81/CGAzLr/Az64RLAI
eSPgsMA1WW8z6DYXcnYRyaPN7yN1NRfxpXZ8rWsQtNKAV8WeFop2YvJSzrRVfYK4
YB05uu5HxGiU/7Pfmsq0eYPpOcn14Yq+GHBw8LvI76Jdcptv/+bzvc1EFEC1S0w8
Fa8tz7xIhv60bnCSxN/TR+g726DM+eCdMxF8wPN8Pza5rphXOfJ9C8lxdD+VAqKj
CdGfQX6P/zrj+ikf39vAYwwN7ZlM1+LMOm9r+PQaKsd9aqScOVa1HdP7tf53/W+k
9v3oPUZIKPOK+sk51MP0i8wdlPkYWxs/SOe3RpAQPiUot2Djdzdd6N/Zbp2YoU4F
t1aC2kRgQe3a65Q5nb+ajrUtdA30d/dnvk3wH4Nodei9+R5nMW0a93s6vK+aJ53/
shK9QzJT6uXtmNndYfwR41XYgnamb/bu9Lp64KX9genymcCgAo7CppRA6VhpBG6m
vHcSy7WoV8U0LsLBdjuU3FvDirMgyXXFWZJq8odsFMDGTppKZyBRHWGlW5Ey3j5W
SoKbIpG3z4W9UpWIxA2m+Dm6GKDtM9S8JWyHuZl1zjVCjx8IBGFVisAABCORQgJK
bhbUH9F1Dg2xaAJQStcLBUwtofXThggKP64vyzyRl+ZnYCV09F9mJu41PubD0ArX
zKoXWHglS/UtDSfreDVhD5c53GKjyBKdgESnW9zCTIT5kpMYzPiOV61Yxltb00Wg
L6YMkM/hwXrFvKZ/ceEsjLF/6HuB17KYgHuM1I3RkNPtDxj7t/s37OkYbYv58iXZ
KE8P1eFBPsik3m/zeMZiOVJ7lIcOZyR+PC2A/dqoE0nRqhIYpgaTqZIYjBMt618p
N7Gu8vfGJgRhuOqAQHirqsYVBYC2Cg/6gFay7T1K7favFIwQ77T/2zSrkvyoSBID
T7iw4VXcI2UOrLXCN2vKeWiDlcYBefdr0meek0ajJ+5vIe1QefDlGblTfSHHB6b0
GX0ytugnkW+gwfdxnLZyyyf2cCrZ5y+WX1xCHB9z4KLNcoB6Mj41YyJyyY/bhbhL
8qA78WOCZ+CSrC9ZZ4Y+x4LPuDtOu7UNAwpQXlj/Zu+l+FfhPSSypLwi8Sw1Ttdd
KwvZQmbC+S7SHEpmvO2fvrY1HrX8OvmNA56LtcE8Kd4is2pFL43ICGpOuBHH7j/D
xk7F7+dfwQ4dM1nHhfquuFSNwf3DvpHPN00yMwxNt/lsgt2AHFqwr/OYvMAo8o4Q
Cx/JX+Jy/sDkWLFN7HKYpg5iNDmMfUMaPAvmMnu5ZgXibqvHLbNBB5c2/XGHm70M
nJfhK53yx969Zd0/E3/PNtXBhRgxJBvuvC9RMYDZc/EwkC6R3tepXA4zqwzm9C3k
Kzf98/4k0I7gKZpnyegzKLChCVLfk4/j0ul3O/4VzGj06uaJN1LsxbhqOwWhAu7q
thWVn9X6FTIx+bH9hzEutmSL9vEzh5NR5IE83eCk4weheUH0PPecPEAm1/azH72f
jaWRttSqZ7k3qucekeH+tZsnLxn89gL4pGtfqRUPCUvumytdVY3tFJhAMBECRV7/
vZixBmya9SZ5lXmMR1tL+bh1hhqYhhZHcBvqGaqpYFMGXl8T8Su5wvSrM7HDrA/a
Pb9wCkX1P/Xxdd9D9q/XEvAcRhdY/8lPgEoxu81F6k957yvhDDhWmsNSL1OxPk1b
QuJe9LaLQtTY8dSoH1Tu8CdGtkCoV+EQwheX1MsOK06skzwcPu744b2DpWZeGx0f
EtJakdRMhDtcKlyQ3gLq+Wkzx9Oz7qdxVb7xRvXe4+soamkzTDkL8NBP5c8JnLiW
TYEkM0rUirxv2BXXnclTnuKkUFVo/K1d+VaaRDFhbT59n/aXIDcNTkKYFxdRJLGd
C2OgKJsmw+GMj0+5K/ypXMmt1jIk0qI6rKOtUlYXmqiKfI6HNIk9kFWA9bzl+sFJ
Y7CsG21axVioAORrZHosBKjaY2giEgW6TlkO9x584imqADEXBWq16qxw3KsJ99AG
yNFWLc4RVwfHcjVQ4fbd1H+UfT//p0JI/N7dqAaVfBSUTAhCpsEioo+TBmcjB0je
D2SHbLbxFwAzgdi4PVCV86e5/aFWvF+Uw0+feg2/h5cUTyaZKdhr6otg+Eg75ApE
8MFqHyDWtjBDGI8Bd6HBmXjD/YVrlNQ//cdnk0pCEj8zKmw9X+sxteEP0OK8GgbZ
97I70GR0tYSC6MeQzK9Jcdumb8KMnvUwGD6hKbjyCyAibmnpLNLyyUEXXkvYt7Cj
FKY1RuBU1KsWkDECZEMqrvoapZFM1sbbPneXRONba5cKt9Sx4OzSv1GVtxaVin56
GlucDgEzP/a5oIUQ14MgznOP2x0Kmk2Azxxwqkl8tDUOLsrvYQEi5L9jF3VB4+HG
QdC1qNb/ISTjFZ6j6vwRmRWmDvKrrSJqMiz2MkLRcxFgtx4WK8WdLzt6WSP1s61L
dT1O56RUhBH0pRmevqDIn6zwldqEvt5r/HNKz20JaEIMFqhIITfMmUZWTVXsRQki
+9T+wkTpinLpVdH9yWu4+mTlGnWYbuG/BH/L/9Oe9GQgYQ95C53SLo1Mb7cLVOrk
SPsNMvuHKxnhQtJE/tm/8T2uJ44UFInHTssu/VPdY0jGYe2v2vTHDU5Md/fKNMEH
x8J7dKmACWDza20RI7C1YWXq6cJIwgke07rl3gLvv7Vsqbs6MYZ4bdQLxvVXclo5
m2N1xWFdAv02cjdOe/g2h48IDHSiJHQeXGT/9HYIauywRz6Ylgl/0yXvGY94frA2
sWPLeDJQeT3BCPflIwD1khj8ryhwxjzFDp5/pO3OaHvoBC4jCv/FljQ6T8pPpC+Z
KL1XLhbR8axf2njMbEifZb3uImDYAdN9uMK8+vHfxbB16n0yqbXhKXYyrZmGBbtU
9K/Iel2iSYdCOVJ3Tso+yudB8LWp9EG0rX/gaXSyWiXZHUo/FGH2Q4OnYBFLTMX8
9f27lSddjCafYxQSwCqRKm/DL5L5emo1r9UteYv3c5gzzmoetDLzWth7q2b6IVQk
kqury9LyJD2uDtUm4yTXGFsovKiMH2DXwlLPZaGqwFPXuSj4DRLaDzO/MrbsJ38g
xp+5CC71Rvu/LiLrUgXPLX1cYRUo3yer8/5LzLdc6BDijYNmJ1IzZhPF6ifZxcGg
Ho6Bw/ecOEiWe9dkerzG/PBxCxQ6Qvg/rUoF/ekzKFj2G0LdTF0ev7F/QyjoSOXB
52azTQidBoZ908VzblpqhxojglBWR8ytayI0abskTJ1dVcTdVr+h4TwqjRSVwm9X
57V1JUFSWrofqF4j5i6/QEdOR95ati+eZRHaQOP8m4wa4t4ZTVmT+TV51b+xSz73
5rdLyq0bbcPi4XntDHY8FaMJ1yU2qlmq4a6uPUu3PhelJ+CCtfR9wuarWg6zA+Qy
QXy397sZP4zabrZJm9Koq0YBFArFKEtED/AkATrd/Z9tNGxfGVVnhumXbnkIeeql
koHgYfaN50BpWw0bhfeLgldIO28qUwHcYqcZIZylzA06NnKeq+VOWmaCMwhKZpEp
ce+mC9k/MC8/6XQjK9QfThbqMYPR7yH5NckJlj+u4YGzrAnJ2xQ+XdjGZ5nyK34W
qaApHsZiuAB5a3hN/s7hVGx3u5iG8NbwM93+J353DcYS3KWRM9Vqru1FNDPZceXB
nhud/0GNF19ILFl4Ny0TE2kuP6jyHzqvlpf+un8lpn6S63QV75L7LgWk/9JWNeyM
adINGbMjRjglnz/og+vH28+8aRMkIBRmfAzrKYIIMQCeIAvkOTJTzd88fTfVRgm2
dqnDISdleoUwUo+pv10EKPZMZrWox9t/connl5mmDlIvE5ryuNMK/+oSOoGEooVy
WFT90DlCkWfrIErSpYWIOqShICb8iv12lHef12tsl8OmV/XiP4vagu/a65cxnh9b
kqB5Gzv/b4Wt3CQWIhJF5gZyCgfzHmwKEk+ohBnY2YL6HBZ/ZP9dQ5lDRz5aBLSB
MDj0p5G3O2KZX34bHSR05OiQ06lHyrukSWVlspO5MMTp/TyYZxF2mnl1cJz4ZEMa
mr7wagVY7GAWsYmch10NzieKupcjEJRWdi1k1rXDMlIE3hgbAL2A4ITrExehadF7
vrEjummhZ/FRZKZ80j3JNaloP3LLvvz4qWKeeGZ+PT0H9SLmL8bnhclQNTQxDawI
yXe7StmSWw0clTG6Urg4Gp06oCZUDDifkvesx2AbsSt2Fhs9WEL5gVLjMlBTWuFL
g+XcP3Q4e0k1dy8r4TBHJoq+VY6ExuoiXyU79tPScn63sXHOscYyw7uuis65MEk3
4MmPuELTjF4/Uk47KbEn0k4TvsX81qnZUN/Whf2wW2PrwLRbpSS9cXJBQitjG/HU
OCoEhQ+LpMWRJVPU962UB9lajvFD03CvPJQH3kOvTSLUdcezmAff0C1FcH9LgZKW
drC87TbIFb5deyZvH7Bc3iN4q066p9CH0148p9qFE3wZt7kZZ40lpEUNeCuX2QJx
9E9m0Asc1JIaYHhBs8hfeS+l/KlPeomFXZjp4Mx20uSXCG6jZmG7LASVEdcCc340
9vcFXSNawFPgZWKmT7YN9gy5379Njw1yHLYuMWjFHs3T3Wx8aInZdlkbWB2v1/Vl
xaoxM3cL9HzhqffvZOezvJA3MMGIsKYYV9uxGfKb8u/oQTYJmmE4+LZU72sWy3+f
mfFtb8n3WKuyP1zn77CMVPKKUrTSh+20cyccslYtLK4q3ywyZvp8CI+rsLvbhoTm
84XBIhrwF+WtZgI7+fR7CLw5maGi6e7+jW8jA/JzmD+Vk0/CiP7nsbRoFWKGXG9h
0MCevEx/UfnFewcPeRUTA8q7KdVMx44WKMrZM17lxgQdE9Ug4ArP+KEXp8VdI0hk
YbbOpTtgDF21OwOA5a8lQlTQr+OenNU5dntXY909XxEDV/rwrHIJk6w4oCP8nVRO
lf49vAC/JWz07rQcdyMo5RLFqHkiQxFOYwdPtPd/3+PGbe/vqp/K+F4TYbe6bexH
NFDy6OS3jGkPM5V8HjISnQfeyQnBkX7/DHA04IzovJsUMogGgytOvi7sf6fRN5Ap
8PiaueXZZQAQqPVGasr9OZ3PZUl1XNRR+airGg/bdW/zguegRKBhBL/Yvt0Wm8GK
hrzsUtWUN3ffNCo1GydMAX8rCZgwMmeNT4mkbz4XDEAooJJ2Q8uSUzKMuZ+d/TbP
EwZKIaNYW7g3JarytCCr4GTPBpo5nIWbJAwov7ioBORgv0VaJPnCkRFt2OenkcBO
+ohXnVac+26DFj+QK4a2yuqciJmMRbi4ZvGYzlZsYLOfKXr/wW8czHpEuaDs3vIi
0+WGzGy6p/47g1rh8SbidgtjW5ySew+7YRu6L/A3iQdC38NXNGOI1Nm4AD8lNIHZ
oYPojE2Ks3RdwO3ldthuLZO63TDTjXKzm2U9WTELXWgevJBao/yuCZo73IBOdrM4
fIL6m2hArGcI9VtSUBrvCYyhwRpczPP4lYK3CchYF8wmXpUaSPq4s1/J0TgfRA/4
J/usvU6paAHirUOe3xfzPccQiY+/mu2nnZOQMHdwuDbkKLwUEFU7YXIif495vSFD
BYQdRDNor2Uh8OzmcW6r48fIXG1KqSNSvBJpeH00rblj9QKO75b7UHVvKN6hkfio
zFYgfLO4vkGx3rkHXQH+K5g5vExHjs6zC+dmuUe/2YR5EMnIPHVR4KEFNV7XUZzo
l3We4XCHMjVP5jC2yEMyM5B1CItPFKgKIOAviXrjfcyLM4HrDiinbhvpFZZzDypa
yAfYplZ3luxODG6LzcOTgd2iMwLhwipyfomw+TFSszc3GpSh7T7ldF5re+h11CRZ
53E9PQbeGyrimQ1YKuuweT8o+Be2A9e8OOx2Bhsi52PBlvot5lQ5V0LG48t2B4nx
7muPzZDB7wzm33lPTnUEiVVPSjw/1TKvS6rqhWrsuRBdLb6k4/wyuNoI23JCkf5H
3vAnivKTVOP2Ao7EryrJbwelPsTgVQxEAX2cgyWQ6R9zXI6WxvMU40QbKcjO6kmc
KIbHNF7NA3rtiZcp34fXzISARbmyHsRi0ACTzxUH1MvIslX3GncWYhRE1G3qh5TV
8Z1mGT7SgsfrFBQpbX2jzAEiqZVQXE4DP/xx27ofGNEUw2Krvnm89/HouxiF/aGX
OdXlxRbN4CEfsit7EAmuDI1EUs3/XAsl1iPHhf/mWZqCfe0TQ0eN8uBM+VyT+FRy
nmI4SKFNN7EoFcK5QJ4GwUUbLpWwhgaOQn6XnRaojVyQvP7Q0hlDVkGP3WA+qPZX
6Fgwyyn8j5NsJ1MpK1FPoUnyUjDQtEbNZJ5azV92ds3Q329pyPPcDsnK92APoqOG
ji89O+FklooaxZ2pjl4BZoJvbP1Dq0eXq6v0qzSdGR3qEWgpS2ggl6nIu+gp4Bbg
h/xOGqalInavDfmF+OUEAXQGW5y59o3UWzhj5koClIP8Z1FE5f+Tla0R/i7QPOrt
/XeCoDZ9y1NpoS9GVgStNVfbOQ/pI2l05x09DQQTAKgaN7bBu6IXXy9obTxSbYva
r7cbfGeytC5CjYieCMpeoAq8F7t0yjNpY8IhOrTtJ/1WrMBKa/iRrG9k2oQ3s90f
9ZXJw+cGsjJ9K4GKOZqXuFaVeAfAm4qzNwTJjEM3uAgTXNJYrPMn/ksIu0k0smLI
WvOsdR3vcmJSH3zdM/9adU9sH84i4kHoMNJvfvlhh+qibsrpqXfabP9Lg8zXAf/w
Ej7x5eFU7OQd7UeNzgRNb8hRxAGy32NUvLKBFkz6OY1HNGwnDWcU2JqeCiMV98FI
qkoKuv0czywjECujJcdh066lqFhk2iuSPlLFMY3+vL57H69dJojvPviixPrDUO90
K8DV2FZ3feNS67PwbVLSMdD3a4uVPA5g8v8fhcVkltFW4GOH7Tw2PTzeIIsnhC+X
t1w/BL3hbDi5oom/qUShs3+XJ2uhEBsrPxFNN/7hqqiEzkC37JZNAiqRYwbJ5FSx
V1kdWS2z+dtIVzUzbI5cpzxklFJdet7GQH+qDOEI2JxBCU2lxRzmmLz/eKd/cIv6
IeUQD7awcWu0UqV6Q6hR4bwkZMmBvmR++lXoQEZe808UrQ33jsXMni04bd3YIjQ3
FpbRiSW8sr817I1eRTwrw0B8OQM7iLkFvefVavC05fNsXvvBJLw2CGArA7HrJN9r
MunOk3S5RhNP66XPWa8Y54O80x3lQxAoviQ3ztIMsNp7wHE8wzQhDgAFUrO4BGt/
uZcWosvALqvrBe2o0oOvzkgnGafb6oE72xGW8/Dm6kFtJ/klWIBgFUzyU043Mm3B
OZc26Py2gALtEmAZKTjrveXVP3zxXvt6LH2jFxzKnQPv1PnesASGPz6KGLDTw+12
HtbATnIDnntyDRlqs+n+olXKx6a6ZgonemI+ZW826+yCbuB/aiykKY+M47J2Bo/f
NAIkcwaZTLbcWS9Ug7o5vFxP/vp7t6iFsjLl4RCgoD3Nf0bz/Gj/GOC1rO+kA32P
76tlDkBnk8VikJOdT+ejpLPig49hdCe0vS37XrfMN40FnPpoPXsgDnzK6zYpMHpg
xDLi5tpGmgBqU4eMWujm9cHQ6h/B4L9089ep+ZOEQALKrUdNPRhPjapad3p6vlCo
MaKw7YK7PBZ60u08J8BeXIJLhgv8NN4sP6RXiMx5WiNQYveOBcxH48TGrBw2nBxB
nm4gXjAdh+bsg7NHWQvnbD6elAcFw+uJm5cNIXGe73gId2Q8Yy7PPFDy4eaqk2uM
tnIx5Tikh3VQTsPQqCu6VI00QP8Dzk+d0cEvO2grOCWgew+3iDk4xjL+Fn5OAyv8
CZHLfsrdBrZnUN/Rck8l0hr+o0eH+i3Ksx5mH0HhCF7vRENQrSPo7BScBqcqQYIF
4R4mWPfrVleZGIoDx19Pq/FPC7rGjVvnblT+PqMgPlMHux+hUB5IA53rOT1Y5Qpt
+rw2lXEsQQVmzjuP3taJyPyLvqMPrmvgOid6B0PLCCOZx6px1nVE/on9zqxbn5ER
HBEgvuSlbBYmTqz3/ATl1txa7xT0iU5fKI1iCE8nKVU3D3Tz/cOkMuVboFF1+s7x
qPwXkk2xBkIkhqFdxNr+WgSrShSrzyhFfP65RYGcubdQf+HLIEvtmeJzsAm9Myz+
06Ezw7K1h8JkBeNBvTNfQhpDryD8rcHWXSe7OtkYvMeHyGs/dYrMVt3MkaYEaAwG
ARfdK/79NhbRCyXQoWgA6EzUvQySp2dejZILZzj3qq5NS1yWG5g4JMJndrPVt0e5
tamgWyzK5iVCBEO+kaDpQcS+SrHpqR37K/iKd79pSK42uuiFfCqvh2tkJhVzto/S
yclq/+pZURoJzBVrsFlA26D+KPXWY6aYTjJoeYdRp7hw2AzA5aIUWDkqbDhgUQst
SLol7ogzhAxP/KDGN3zhgJaa4tI8OxV/mfTHVdk5v94m9cJt/lrIR9DjPetlvUZM
nXu+LjCHVqq6R8xNCVBsxRYgxtSuHj+SetC7d/TWtwFlllukfZ5R8cjVitKbyBCJ
zUDu/qn4aTTVbG8OB4zgOoTlPVHS9zVOqfNqrQQ+nRZjhf4G1f9zGBxDzVztj3Ik
YcjJHuozPijcvKOmNlUXck3h7IAIpoCt38vEreIJgzZFYJbNFUxulK6cIt4h8QSq
aBSMnUa8R7A9DYfyAHR+Gxuc0ixFuD7+zaKCYLpDzFFcfv79Dh25J7ecVOWmYDGX
khvx9oI04Aq0y9tXXcBoyiKgFnyXAUZEeIjy9Arm/KLvlgf2EXRpMU4J8STBe1aY
kyZqKpG8YKZYm6/n3pSOSDqqXZOW0FXjyLCVc0HUCox1XaHC2tnG8bfADZmleBaO
fHtYpCXUwnIgrSeVrzKpSOZGF79bRZAwm8IofKhPW4WfTMjwsZrc7wmwFaLUKgMT
MnJu3Ggai8iobTnoXbJ1j3iOfQZgSZtIY3F0eEwO88FqR/TgyeNRlq10amjY2jqj
q83AOqQXCVMu/8JBpHB6Y+PlOkmp5w9Csdr4+l39b8JKift/ObHyeodIFq9yjHq+
+0/pDV1C160Qex4He6nedOVavV/32sqZXqrNSzy78YkF7x1wRM9813XPlJfwfVJ/
bP104xpQhJxDQ4/OlYLGg5On9pB3yiKoPBhrWCLGKpmLx0vbUQK7KztlBn8iooUH
N4bS5v6QwWYBlyLHj2qrG8B1+oFx6XyajSs944twjfQi5dQreHBUHgxy7g2lES8f
iLelShh3tRAjKEYwdXJbhbqC5klb0ae1EoT2JFikzeVlqP6+/WELIW2YtJXOkoo9
s+tsppqnJ7DO3r2ZTfXzHvailZgT2AGVb4yMbP3IhBpdgwGodL+kcp9boTSQ0+0q
oWLgCz0tqVYRj6gwvgU5bnT7tBXDXww7YlT0ZDj96/b3Arp2Td7niyZyqoWTsZ4h
0Vz2XM7dFa2R7j5iFECb8080OhWCPI8Fy5EiNiSM+d2H93VXZNF8ncrEWNguIKHF
qSHY/LcIX4yEJaF41xyhMCbpR1/HGgY3+7lE2t15/QYrp2vo1qZd8jCS2WNueDem
ALkcDE03MY9nvnJN4xO1PdMZnyxOqv77bnDw+eHqY6tsPwefw8S4BBQ5BiLN0Pel
2ECfzNyPV3/UFMyuJOY2bbyRh5oJ+hiY1OOv0XShxssZ4Or8R7cEF2tT4RaziT+A
t+iRLeT2AyWqtkNRKuOZs06kLeCzv0XOfNeFZ2EmS7NFjO2KeQinv0W8NVpuamSd
RmxZ4/xT0EBVukjoob5Euwc7CHKnsPHghptfLclGLjZYnzAsLq+ckORoYU8MC8iI
Ctuyz8CrmOXBo4M+olWuzowXoh5oFmzfPW6EFZq0JPMDtii5auKYKXdBeIJh7eZJ
n4NZ55wb9MBJHBfcQItnF+ewZVF37t6fJ6AfYG/r00/6X2Jt9ciNhFleBZzmF2dW
YzEOsHYRlj9ZBJ6UyRhvWdIIzkTVg8YDenAaczscucwOocIjUiNVAVvkihuofIkq
twoPbF0+MWozNVRBfxYO5NzZKsb6kCfZEFNfMOyGg0/N40an1doqd4fNmProdsXo
sEF8QW8a5NQ1LWPnDKc+ftfJZN0zKz2T7/balAfM7/Y27R49qisnIIxH7Yf4W6Sp
pUtXVgQNQDC1npo2oYzp9wOukKkKrSPtkBXsZAxsSFBzIAwkRJCJ5JpTjOJKK+O8
GbhE+n1em3ikllrQBf3XhyLlPLX3ne1kn+K9LbCg6z5uDh+JSFLIS7j9zaXVCVCk
OCnimTib9tnKKPwOjS86nanIj+Il+Gt75k4PBTSj3g7nSyDkDC8J/rkkL0TJQaT7
fttbJ+DJnqVs0M3Q3LHo36Pe1GbTWYoDF+YrSyvM9lhElxXdwN/cVNQJiaR2M1GG
Bpos5JaevPB8QsiauHswNlnmPmG68TV1/P80tcXiShvQWsDiFEeqgFwdjip5jrQ9
zFWFx72CywPEr9RWhOPiOT5YxrBheaXt7V/DTFOxIvaZ2rPsi0rkz0QLFOrPK0Oe
2sU368GP21bado0AbppToOJRlEUIAh7WS1C38bqb7rygl2JmkFcZabXzzcShy+Cr
KMFrh1/giq7gxhnD9QfsxJ4SrlX+UYXKVP/PsqXTSU/Ol3neWoPGIujsiKU0KN3f
3JsStuUoZkC8sVuNivc5550Yy6/Oicih+K6EdSDzF+HInWXN6+4UuM9daQgdgiNp
yOIXpHOzD36xZSBjFVFZw/oPr4G0m1oa8++svTEiMOECeG20HxLXI19w7+4Vkboe
mqa4xNxIjF8H2opELOHFGTgEIsZXi3+GLFsvlbpj6CIY1ch9cS4jrBxnTfFqzz/I
phZzBC01RB3XYs/6VL1g28m4+jCsROU/6a496aKzZyA/+emWXIQxybqdA3QKY0me
g/hGqc5qrPkb3bgD/gegzrzX6Jy5PXCfJOso7hRMrYtR6ojosMdiJ3ZVAZ1ULPYS
lJd1JhYyzCtjZneSpiIKO1psl7x4ykW+gApOgnBbPnu8bVoFM6U5MU+Eh9EJuHhB
IRrJJ1UhgIcyLu86TMVJ6m4rH8kfpb0QeML1Y83tLxuXN0TJqxJ/9uBe7qwrJ0RJ
Ya12oXjJYdNAUY/UtRXRIq+aLgWna4+e6NLOVFS39y7YUPvAfvtJ0xP1SyAzK+z8
8SuibnvUKUelKj1F+4wVwS7DuzYdtiKYGWxYwSMv5QH7O+/iASLQ2IdfS1sQqPnf
H30FrH6qnMJUc6twDK4MKzky4CXXGK9qkeAWi5aAeh5M70k261mT0jhdwvoDgXYv
i0xYHvvZbdPrJnE6a9mgJNNNF6VJoy8jY12GGNm+BExl+Tt/Jj6wiTeFB1CRCk35
RQWFI710V7LQZ5vo9teJYVVpqOQtV0G3s9yVUrfYMWqIiGGNPk36W+WLvE+dyeOx
vOuMZtEL+Q7s2bLo3O3ghzxyMjPYBEMlWAlpoFZ2T55ov2heTVSIzDkvpTRST+kX
TFj6R88r7lC44tGrSZzGnW4NzR604hFbkEghE/WbxW5Z+MzkuzKerEnQUX34kjkr
+H6WfYhUP46rihODaeZ6YSW5q3z8JzKgUwl6vNA01VCYgMSLwfOvRf1/8r0jLM6n
hCvfdFsoSmgvlAvq0A+s4zgPHbl4kYaIUPV8VTS+MJEcyrD/D260nUi2FiQmomVK
xmObP0T6qDPih2sPqLR8Xyg3zNcACe7EgBiFmctKbrzsmXAoGAtPEzVcrnHonOL5
zZvdo63w6gC8nu93Q1tjwUlW6Yqbhnx/H54sE9uiTqTxG3osw19oJS1DscTpMc0g
18bxo88LyW1XNyRx7nAWcUevzemJleljaqcGEx7fQIWibLdXFW5Jr5ZK/l76lzso
RTzk/h+JwLF049olSQZx46+YbAdOEKf4ytT1WXdizi65I65A+fMhquDE12C6NB3j
I4XtpmUPqG9W9mJqoY8kjBQDehuOc1uBARf5XQi1sFMW9n6NkCKBlF7w7L31IPPz
iSducWMN41uB2v2eYEwO4wM4DWO39JORXj7nXooWVSrb3vQM3fPQN/LxMtqHGxQf
8YrfmubwNTBgeiYsYmMWPe+BJyr8m78+JZJKYtCMBLy0G0SD2FyzODbS5tPIXnZL
SqMgJS5pa9eeeHROZx2sfW6b4lBQ+gyFs81Rw9iV6pU9QrGbDbw3L4L31C98rNlJ
tJiCgs/0Wc9kOyEmUlkoYly1pn2IdF7z/tNY+rmeMZNJupltSuKy1MdNtj/RC8zX
WiG++zaCy/LdQFEtQM2h+Ky4bzV+gLYjw1I9280CXdoSV/fo97IZbDOjLgurFbgV
hokQk4R5PCSQjNg100k9HjhCsKuO4u8F8cTLMzOO7k8H3UfSw0f3bbkujzWddi07
dYIRe4e+cnXv1/cTht6+0ZFMi2j9Reo3CIYT3nIdn3Ofzoycvvx/4e9ueP0wUI4z
lk8Z6nMQyNOK94hBjUZfN5m+ByZgx92ivPWitg7jwuD1RorGD9obXiHrXjFG3bZW
9w0qocNKNz+wfpUzHspsLA6I2gfqwEd4bdHOOl0wnlMa0PU53gAXNMBs14qfMjOW
Gof6gldceD29HPv//iiKsOIrB6KULvvVCQxKfAVhi8h3R6pOSfqwanVvXUpPtVnk
UD3CEu3pRfy1JfdwrQ+9aqYrj0tDJh0BedqOIDni7ScgWyA+IgXeCwA4rL8c14ZZ
Ps7T5Edn3uWFLx9+9ZWrM4qH+EylARjj7H0WByK6CvoCpgDEoWnZUFYqZe/sXAPG
nY7QAZFm/DF6C4CCxF2a4ZaGe+jPiVuI+aBHD9mJHiTBkYfV3F9uiD3yfeehBpD3
lbYpK/ghR4Fp6T/8TquTgrTvOJcyK3y5JB9LjFOAyxC5BFd6NCu2z+0KqAMg9xgP
QyXuh//1+V2kLSbjojnTe0xLlrQkJKp1lXHfECwNEW0Bt1R11dVYm7dBhxU/Pn4T
qU+j8SzS4wXT7hyzMLyAEteni5Xz2osfSUvlYuSqd9XYDeeIOv1gvCzTnGTfbyEK
v7cyvhNLxXKiHDsJXM6L3WqhRPZhyMrMIkRtTkypbNbFwK/cGuBCV1eHawSWYe7k
uRB9nA5iyoTznN0pEwX8Z5/lJwh/Wn9tjFMpdpxxSBY8IOHc8wxjY1cuF3pQTgRq
LV4AlG+nhGS7fwQpe2gdO3L5rH6FJGD61XRJxGzKnMsW02iupviOMrU2OQNAtq29
+xxCGfTEdTmC+/JaLXUVkOPMbV/Zr5O7tcNs7r1fNLA5CGjCGezxa/3IQK8gLzpn
ZbN5sBzNe2xW8NRbjUkdiUuAO1A2SUd51/KF7R2Anfc0ueQzy2RQ1RWSxXxOl0Kn
EqTYx8daPh4yA7z3xRqPEkdT4RUOhaXEPzRCQDJuymYiojzRLRcOg4ZnXd0UTYjq
DLaax98dwr1gpwWO/E7zoy6F06KQL+7DTDvwg1v1dDE9P8F6JKbfbFny5hIOHMW9
igN99bbaVgLN4IQABDZSwf4/glniGE7UwUZqhloZecHNxXulN0oHuyIlZpWWKWMW
6l9s4jHWibx+j+X9FffYUp6YPlo6rCyBN9gp4sdTUxPwp3xgzNUUvKrlHYjQMME3
NH3yN5xp9DeTvthWC74Qzkump9HjYZbJjAAd3K6oYWqY0jWyylMyegSEQUzDstX6
4pksTMgxmqhWuSDlD9aO2TLru5IVXFNkc/rjnkfhU/0=
--pragma protect end_data_block
--pragma protect digest_block
Xij6UtNqfh3Utq7TnZ0NNEO37ZA=
--pragma protect end_digest_block
--pragma protect end_protected
