-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
/zsMLsNBuwVT4eZuN0D6LM7cz2f0WlaRbrgpUXJC8SzPmuhfbjkMTv4hiS7aDZHu
FQX00TB5vdclTGFNe5nlwn1Q1hJpzTsNs0mRTkrOmRtRh/2gptWSHvmKURprMVHP
nnH4cUAgl+3tA8TUCk3cHyGCIL3vu/4hhbUYbqlbfwA/vKJmtx6nKA==
--pragma protect end_key_block
--pragma protect digest_block
/lkjoCxVcxhcP0g7iHhDqpPHuUA=
--pragma protect end_digest_block
--pragma protect data_block
IS2F6+FO/4jmmDlcT99SsAUvO0UFOgu8qvXJU/ezE4BL8fPWNsgL1E8DbUMPUHgj
/wJD9mMbj9RtsDtTQVSn0hMeow0+zq9YG4P/C+tfVrFmNwgUWL+88f29uK3EzLAs
yUjfvjW/nwe0koOHbUaqJXAqoV8i/t+bqVhJzCwY/10I1sctVpokdnLl85yhzg6A
GRkNAruql9s6d4pPxg5nOe6Cpas5ymEJN9jg/8WCpFZQRd0h23LAE/uqJ7vZBG9K
x/mozwTJYeGcn94Hn6l2Xk3x0OlZxHvekIr59zVpzL9eEEudEUQKE0VuTjaMKWPb
HbF3evphjveXWX+CGYPTu1Ky9Mm5eusL8ao503OWPbu7x3g/lNFfyY4WCrWKt18O
j8YvRvXZLKtHqJQcnhJu0Xqp0cTrUpx3UNqmThMKOUW080iQvCZMC4kbbeevnSWg
fSuBVOR59Qsfn+jtg4aEfnPPBIOiWE87KKR2LC/N1Hy/tltC4s6Qx+ClebswNACv
GLGii9zVDItwPDQgkj5Dcz8Zo3hwNuZbrD47h2c6PHgCptDhD4A67ouIekCZKTze
aiMOmO02B1sncNRidL2eO1gNkoEdC3E8tQRcKEuin7up/4N4LpfIx8veDRHMjQ3S
lSq9vrMcTtCzhoV+uroHcPmq7bWG0AEFPY2GpRX7jrAgRQ/S0dmEYR50Sy0KTXLM
UNvWwpl37xh8Z3O2q8ynIhVb8ACHTr1wpDvhO7Ag/xV92p2RIW4QCsB1kISAH/oE
X+FyfA6QvjaI1RixNS1hYBUVOCVCrwAibN2BzegTT9F0zG5lKAFY7aQkau29yGLG
FwcbYFa9mgI1b2acU1HAepmK3intKol8ntDIhphzTtAhsOrkDuv/MqTMceDopwTB
A1TuAgeu+Q/uY7BE1rgIpbZAQ0UVFRZ5XCyVg+T9JbSETPncz5iIW6a0lObl6iEs
TnNE9eVTbGmgluUpjReXtrGGS6bmj/Mf9USWAiUCJPnjOVEN1WCK48BRxW+dHJkq
l57ipJozlwNl7YuHdk+eTrext64hjnHT6rWuhilsAf4m3TpZ0ztPIWJDLmHp2tVf
rVppnfULMcwLBfqX727mmPsCNXZwVL5NkyIOLEXZ11K2zwYGteFs/TE+k2aEmkEX
cl+zJ/R20DCQfqfwxkis3zCMqssT2MDmig0dhbeJ1OMJ7M7GUgsbuZX49lpV/eta
xmDbaLtaoXPR95SbSQGbzWidEj6YWITa2MivtYhc47XLb6n1eMP+QZkD6jRCA7ws
RM5fcDOXfCWEnNBT1iqiK3CstmxIM5m+kh54jzWV+wksaWS8Tnfn4UUwCsm7KG9x
VssH1WEeA8LypF59j+EABi1CrVbUfubxOjJ4gLNMwWmaDJ2OjUSQBZjoEILXNyPU
AX6HivCJ+6rMo/kQEd9OjCsqOxDkGeWm4wcnFph2gkVxfRgVA5l9ooE66kExokqu
kP7nhaoDkR1Sl5RS5r4CO1ZYvB38PVd357TpSVwaEu/olzDyQCHxc/0ZXc6vmphR
TpDQ8CRxiMY413pXi2QZ6qqCiBEojD8kfSgKxCvFfU/IrXxO58HSk0Kg6MdxyMOk
XlZZ2qi1+drJjDxeIwF29Kl1E7P08vKZeG91W/NDFSRVBxals/FqxELG+L23tfKQ
7vrkLaE30HuJvcieMqngNXS7SEi3AeS3HiV+23B9vgiDcfc323Rlt4SBlDOaK4h8
MlWmIYYwclAf57un5wa2eLQ7ECYJ8nB3lwRJm6AvyINwdtdzGNhs+RDgRwtqFKs0
ZNKd7Oqut6AjZJtFV8VdLEaVSPqTmJ98fuUthx0QDMj8N8UGIXleYvuyeQDe5q3y
fFmNjJ7BWbIOZ1oOh1/KXLABClDNG+8usRQdOjdnR23QkjZZX/ahwol43t3NzTJa
4hH02WZbpmJGmpqov91k3JM+ALfh/9ldMPqlNqwmsONZ5N68NEdEkoLuBngmyFdv
n6DNi9KxNzUs9WFftfLOa6ZYtFb84YxG7g3aVyjrrLDekD18kmubI6kiG7llxsVx
8TmzrhOZLO3iIylpekJn31XUIP+8rEwHV+rawmROxWTj9SLSFFYMEhAIzQfhOfCB
WQU4Ig71MqiDCNY8S242dIL+IvqoNcgNs33D65dgIYlszuTs+ab4gQSeaRxxUvFm
iJyP1QRQPhJV2t8aV0OBNZd4/NFsYDl+DOhIsxrqj6eMsx1zGQIjApESuTa3D0Xf
cYVt5XdErQTKFnKBNwlfCNA45TYXU62D7M1THdAR46YbH5FP736EO4KcFict1QHL
0PMP57QGp1WzxlHgPyLHcPsFJRUwVlPrzMWQYv+4tRg9qbizSk1TqLbjq54i6m+V
WpaZPUBxffD3xvLGjE+HJzGq0cC8jSLQkT51WW1A3M9nsjP2G8qjH7hCS+36FHQ3
hXqHxXrauv2zjII8C3h9rdUjii4g4KIKxxNF+7lFla+0LRZDAU1B/v0ty6imNUYn
6iU1OkrJYeQrjL3I/YGdwnI+TmzxlQwPEeJB/HaAIw6HYAnOHF1+Y+XZvGirJO7y
x0DKblv42niijz6OUnsbbgpzpTwvDRCcHvNJY8X26xWcmGndJpCQl5hm7PZ2S9aX
aOoWtXk1mzazo7J9Q8KwvXZr3gzRwIUVr4896dMVb3sjNjRdjjRJ+tQB0jtB73cv
cq8lzipo5nJVkza9znh1sD8uBX60ouwoZ5JuyAurfKlm4Ahp4CH6Vz32B+xOnJGz
dsn2XTiHpWXLKvUXVjtzs5TOucY9jqmJyPrqaUcjwnvT5uMm3ss9HTrSD3Gv8ALP
P883ruTlfUd3kiu81sei8+qvv1bFMuBntzkwpBO7A060DcE9+s3N6EiOgGJ18vpf
7PnuUImxk//XMLq0wcFFizCRPv1y8/TZLcf55UcUVNxzNhNwoEBXNw9/8pk2fBZg
CdLmZAjgqkoWDDkENBy6ZUm/6UH29i/P53FUwndK2JbDAyu05uLheqxu2fHUrWQy
yH8oSRNKxWVJiaeRoZx4yhO26YkA9OaCDHQPTFmuN/HZLHyOSkpqGP+BftXCSjkD
vSbyqmsbykGhHpwX6tkeElhbfX5dr2I5HUbge8PqWE5+NTqtHrVeQvdfIYxMcegb
XOpHlstGeQz3gu2KOYQR1pNScyzgxb8tsqimVPQE7RMn0ZF805DHn3PXM1vmB/vw
yfc01hvdCf6GDXmntanPf3P9ST0zRD9i2TAJJviRI5t6tkZD457pe8ZPA3lkd49o
T1g+iqhs4go65Hw8V1GWw49WRQAGT+UUl21S9wgJuwnf5csYPRAxr2ypJsojz7uL
0onPWuDogziKZsPYEGbaWLr/6xykKqieWPqVk+JY4SJUd5OnuFJFG3BwpYY74OTb
H/or2ozy4vBrULvMJzGgMikaNfyZVOm2IU2DvUvNVTC5HOSmZtzfKUZo2sJAQPXo
MbJiLFAi+neL+TiXIW26SD6h8S/ApCPvj7/XO//U0pDZ9m57Khh8q4LCKhLEY8KT
lAk9c4fP5MojUvHFznsSRQHgH7Qi2Q3wBR2ZqZN+cCyHNen8alSZ1kjhtZxmLE3S
pCfW3xpktpicSbJVdMpfKPIcj0KtAUyaTWkl29UeTFzG1ysOhdRxil/jj33xobXX
oiYRf64RiNinWvbdESCdqvrNd4xM97HiSjhzlqGClXl8hPzA0BugeQG2BtXk3dJa
Qy6Ta1aP9N6MAeybx/Lwv6suK3o36D/zvXgw0bsqpc5+sFPiv+mIbGXqFE/KzMCP
w5djrqH7qcaUNcbO/0CC1oakqcJQ+GrmgBk1CsnTa+jzXenOD1AEN9SQw8LDOtd2
aQ3NW1CWZzpgYGykCd/vOi29ghqd2LxBx3sBD9aQOMxfh489/XWD6OzTbz2d//ZF
rGzXwu0qupZ4MUvj251PfSptQ38NgGQp6hGcuNl9YR0ZiSnvPs9HLs5lWXY3b0lD
We8EIOsaghkIF/rjeGpAeAvQy6WqY0AreOdZXdutVdbLKaCMqnM/IWhmW6AmRnWy
3vcwJ+7ZR7b7i6CClkYhtxsOIfKENGsIR4pzbg7cbANXATzaCRuBSPnlFhLrIf/i
SDLrGaEbcgpEtDAtblx3e5/CWY8Zk65UOpP0MaXAUaDVls1bcdUBSvxXuQ8BLL37
sVXSoN1XG4NgxEloC7E0ZaMYSNSAFTLyoN/dYvMKm1hW7CEkcjp61HKMTpD4hD+n
yswSW19pdwMO/voAayuFZgIsh1Nti92myy1KD7sCW6LOe1dxfwZMEBu2dc1U2JPR
73jsiz81/hQDSmyoYPXPL/HtAYIjZDZXbs8bj/l1AKYJBIrSBcY3QyoszKMVqT75
ogUGyTGN3KCtsqT17SCIYh9aNYVqr9qcURaKSaUI3zMVwB4rMYZ8cTXuUUgwgYvq
9ItDQugFxuFQi4Lpi+3sru/Cd/0CpPTar3YWSrLM5BW0en7t3rRxWswwkF/n+k2y
wT0BWvIbF9lK4U9yIfLxndkC5h65cHd5BE7KGO8MHcFijt/uB0KMS0aT1U7/1G60
egn1W15bTar38zfzCjOmskkSkjJWABfiuah7Pz7Ex48wO+UgzPlmGR+/ZBk28iG0
Dj4pW/YjJFNEKw+D5p2IarxoFjI1p/Tso65exG8tbtMLGClE3cuoafNRLoqfk/be
TTaF2EoYwl7utBUxqVRjRLLeOq6Y4WmjfzYGvJBVN3zCieoZc8dMfqrdEH5qxXGC
JCjPTJgrTboGDjz0aJQNWVgMusH3hQm5H1oboQQmIKtuMIACQYCt/FR1ThaUK/pj
ZkxY7F1rqWVj3ukM0RXrJpWoF9K+c26zjKZe4dMDFqbsjnI/giE6vhG+GCFrAZ0g
EXsD+ktDs2Uk1wI6mHXhniUsha4auCbM9zbF2aJXjUe69CFeIGgpFeHLzJiz7yfw
Cw/YjuJPUOVTPcDa7wnufGqnmbMhK185oaBZJaHRIk6g4ykduHTvBtzsFQqjt9nl
DdVqQKffATk74lwsWNDj2s8TNKA1QO1nMtPq2iCT+7MZyDzfW/XgieZOAfVW5iW6
PIPUFUtRPsGGONK65P1VljH5x/y3EldEHAvISj1L8HTs6OapmwKFpef5xvf9UzJw
RnpLYplFWxleNQ5ZrRB96XgTffc8X8cDFCdGfyy94IU3rRaaFz/TZuVY1hmDifUC
h32pT722b8bniZr/KdJLt1wDUZp95dWBNLruwJDOCdvjV7i6xUVigZ6FNFVphELr
BN9GZUUJmQUKGMeIFmGwyq3D2MLpXjJ1GAWzaJcJHBWo3ls+AimL2E07kJ1yEpeY
oQf6kZER0DXNdxHN2dbWwDt0UpwblcF9K7R2jzCce17qZaWAJkO0BdOh3G3uyBbu
WHc8wzG+lWzn+s1VRRydvcDCewehI4LIu2QTyfYgpiAeC11rwahcUPFwn3WMFruW
/AfnWw+wzGNIfzKYAfL2gI5Ypww6MkwAvjTNax7PSH7yGuYYjorX6BJ7dHmEXL5X
jxxoIXK9hUuHTiNh/DdUa/8WAlAB9ezEPNbaSt7x0uTz0gmSvMm0KgkGViXGJ04P
WmfHs/4K7w0HqgftYawZJ4oE+5v61pgtRZgDGQi4QGZHg+Rw3btPl2weV2AMA/Mi
Np1zy5JA4bSxqRXwG6+G0BfP5/rJJMDxrnXn2sv0Hb/160nljiZZGU6iocsp1y9G
5cadvfgA1evM4craPZfVRZzuL+4c0R1Sldngw1JAfCDedpOycN4bCQP+VCoaBbuz
OtGOl6EKJwBWlWj/f6SUP5QiRpH5vye6BRietxslC/pxrdZqirfUAH9+DybTun0y
+Zlk7aXoLiNDh2F5HDWyj9aGXSvp4PUNCRbHcDQBFKHfQQsgfXj9i5pgSyBaffZD
Kg9wIERZLvETnkJwoJe8q71DYs1gFs2j31B6OJrpqKmOegWo8L9/ms+Vogj5YJs+
8js3D3LQ2iCOYPVTA/3E1BmGYUCXKUW7vj5MWfVrkHyYIxB6XXYVtkm79EcgP1+S
FwfptOqJpasGVkBxI8Gn27twHpdtAvU5MpMtUMwsX1CL3OagoyhBb8WLS4UFwnz2
whdqPv3lPoy6ij4IMI6VbOx8JCNsEGDymNma/nmVVL5KqpbVE0MYvJM3G5S49Vyy
F100sLJrb98NUpWVFKgILbpO9DlchuBBRZdWChi0xHDS8njvWa0jrjlheUQaCpye
Zk//1Sc2dYxu0CbeMZNDj0PXjR+qHaKC6eZRne/Xp3jPu9uoYnTKeNkbVgYatfEt
OrOjMfXOACNGInpjr7xh494rIjPrQiJ8G6He125tBkRl+Vso4zonh45Pas92oA66
kPuOv7XBifQ1RCYptc4LIg==
--pragma protect end_data_block
--pragma protect digest_block
T/C8KncII4yU1QXmkCqEza9eAns=
--pragma protect end_digest_block
--pragma protect end_protected
