-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
h9c+mFpPXNTlJ+l/Si4slAGwasxPaTIIcMK5NHLzKQ+AfHczXDq0hr5gIMwPQpM7
josVWb7lxp7PJmHrWQg7wuBd8vcONXB6QLWErQrOFH6H80E0W786KPyKkRPaibRb
8sEHhKR8F/3heFgs5wn24JPiG9WBOdWn2t8W+MW8LV0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 111940)

`protect DATA_BLOCK
VrkMMw2GR7UUg+L4PYRhXN/BljTlFdbBTg0zynNJ6NxiZOHckQ1nxft86VEgjPyh
v7cOlM9e7ms8B5JXkAvOpbtZVSB3H4dkw0RQ5QgcEIGAuJEuRtgQLBTyOe5mKKbH
yOFXBjaXIkNgVaC3Mj3g7GGdV7c2pD6po3frnU5+gQZtqWZlaQ27VuSqLOVT4mQI
oM2EIJd0KOfZy9d73bMOJjMqyct9M8cZMA2SVfvrENF4LVG/k1roa4LKEFqXbeRi
u8xP5vqDV7/ij6pfmL7N0CIzdRNsJ5sWTwIVeuHr0c/COoW48cMpKHhmuWUYMbPJ
XZyjMsCuyZpeZ3Y17d6EFlXTXUQ29ACXjY9fW9rN9r3D2RGszxs8xe7G4P8l1bE9
ZI0pWkSpWYfewOuPaBS5wBYSa9tzYStusluaqReStb6lDMo73QkcHYW4ZScrP5b0
cOk1ASX/XeRs+OUUZIEMTR1jGxe9ReO86SY9E/qro50RRCNQxGgKX6jsc08jJF+L
ms4DznrBj+cHoAmgsqs/M0S6xAUwFK8xJFDf28W8NLblUe/NoK2oyk5/ZMCCYO9B
/eRac5Sk0pG8IAIGfAdLFYdiEqunlstRPl9IopcFD+UaB12ab+Z/B7+4CjWeAU5w
nD+TWe7raaTFsrktcDXzVarQHLQTl7OzONyVh1pOx4vKXAiNiAT+WXXT6gk+E7Uw
wehMpc3MEn1b8nIjhXoSNFvv9ozzRLTOkXasn25/+WkUNoEzyupulZOpo7u0ISCe
3vLKAejh6qZXtJBG/L1HU5QfRBr49FFxsyxACJoCoTCYh4rkYjHuJwb/hpnmNv9l
a5G/ibpWUA14QbYe5JiHTjAkamHcWDGksIZUucxUhkAW066K1GbxVR/rk1hlrtXS
KDI9qkOHxtG+am/ux+IItQVncFjd8Kw9vEJAE0Duz8fMy3d0Zxc4dbfsmN7AGMYb
HUaQEcWC9N3QAbIQXQCJxTR0sSYwLAlLst75crXEIW2B6NUo9IqfGOGk7IJVok15
Es4X1Rw0wNISyB72spu5XrAygQAIJBbcKLFhAx01PDasB9WBjFZ6tkVZ103rokQ2
ZvfZjoeOLVzDVjDitZDpTBOTqZcLytRzYfRZg6F+U/fDTwUy1Nm9VXy9v2yGjOhg
kDCUK0spTpsC7dxjhs8n4zWg4oaITPqhvuF8/YjHejHMSJZbkqa4igFFkRtCb2Hu
MbPmPzE4+8L5uMQDrHVUSvrFRPzlLppChoAMAcqPeoSDH4RK5WQQe4vY8f6BSZOq
Z0J6ueMSCL36tVEKNrHFMMNOxiwp1RxscZJFCFN8VTT/Ak5ODNs6Spk7fjbxIJVg
VW/chgyIB8AFbt+q5KUEZh1/z4WwNB4qET/ZY0MnRVGKum1CSouaW/H9Zp2Yng/B
DCjf/mdB0PfPOzAECmfFzeOQ4sUXYU8ZWdVAIJRHjgtNM/nj7k6sUpE3e3tbBvRw
qiizOdGxHLTvFgreVmMsBz3+DIXnnKCYZB/CGtmQsoSewTQaDjVhRKWncwGkXgXk
XM6BOfLx5H6JKh3/WWGsS1A0QQLeI9Y351mZce3AywcZgS7kWTkmpewtLh5iqvl/
2vDpztw61slJooUmd9BvZiDCxAxIfp2iPrJ8g74W5mjPjBbfeViAmB5Ra0CgMwkR
QDcyP06n3LBx/e8GvrL9NhyBlF5dbCwK7ozWHGACzEofRqIr5F0A6T8TZl26t+88
boMFMitplty0amGI88lTWfJ+GQsjlTrdnQG+URieqpYdTtGJzWFMYFIXQrWmmcZ1
0UNqJcLx3Ys+WDFFGfKW2hObZj1ZCE6rMOjqNl/1DRWL32XtrKX6cH4gNFqXOHS3
gKgkXdFxVD2ieZxgTok1n/bj54R/nUpASr73xIrybzg7JxPexbHhEUTRqARCKKoT
smaHpQMG0C7mo0YGwHVCBNLbUYpR6AlhnKP7HzrS4xsKjctPMHO9uIC1tgQ/HvWe
t7ueD3tOxCEGFJ64IU1PYyMPFZO7ZKkSSIblDoxQCNr6Whr33pc2SyMcGeOpHXKP
qWdPgtEYzgfS0pw+OP8KhLtO/tJNGCZGN/NHRveus6I0B8TY+VMLfpenC9Bw58L4
kLJFL2aSHgQqlLRYO5JChZZNjUtnPiIzLBZ98ImurYEfsEEgrD+BOPyLpLTWytB1
36h7nGv51wKkZFzSBUo6SLRcRwsINsXM2iNoThrL1A8RlkXw8nmKuqbgqvOpYqP4
B9l0izJuksaXDq60UZVIRWS/J0cikBSp/26jxYOu8JmRGpottIitruWVKFCjrX97
mYu4Bd1aAe866xm/stCpWTSn5rhV+hKE6eGOLY0lT8dqzwZddlEAuWufYvhAM3j1
Bs4D+zyuMlwqMS2jylODYD6EGbu5zLEI/em9/zMDSDLUAn/kaAYAl3WCNjBXEusK
ujNDYbrpWWngcn2KxOE7XKpJIGPcR8aZDKAamqzPxXlupa14lgZHMbbtOrHvzhpW
SciKVN0Sli85aUgBmby6TtuqJuokgH6ZHqxGVUEd6DzmqBWv2aRsY4g5JIi8iCy2
IMYTKroNJKhR7EgscmfvBn9/+PLuuR5SjF/ezZLHFa+Pni07RYlg5P6O5DDBnX2l
+Tq6+JZzGuCc6tXC5qumFvLIfICRFqCB9xPqlm2/TV06+inGtBblrEG5HwfwKyjc
Ec7Ih6y6FCfOAH+mBRaG/B3xFNFXGGdgsWc7DNqwa3O9hvVIVuxLefZ9e/GfKWah
hq9ldK0YVnWJMKJpZxtDQzg6oYOuGP2Ni3kPso2qrlwS1meqIJYPgVgd/yqdEiJr
1hWmUry3OZAmQDwO2z+TxXM4Wuvhd1OvQ7gnPp8d1h79W7jvaCfpqQP9wvThtbo4
voyem4Nj17aGyYhr1Uya8VCRO/JHfKTgXv7Dc3vEz8MNSALH21K/pk1gSIa0NcCo
URvBTzChgxJcFYt9K9qw/IT/CndhQM+cNj8h7vs3Y5dfpfgRoWsHVKYA3N4I7axl
1Ex6JLxIw77kDj4DDNDVd9aSJlmYSPuzVRHkuAHweCTWbn65blZvKLjzuWLMdfL6
Q/jShQ9nscHYNzw5oA7n996nq2qK7rp56iYyi1gQwLp39pTpnbU5XWD4DidSkTgB
8ka1kBkSzyI7Tq0/BZrNGKDw1HuRqjjFoXHF2Mx9gE27qI8besHveJ4hrrxUOUV7
htlWb3Ka9PWKdBnGiOZWhUHh9t2R7dDjKBPp5hXAXiZ7Bbpkg9KJmE1ItYN/4pDo
k5M+WRQJmVEaHfmkne3SnnZSCDtIgQC5lUJObsKwhMCpCNpKqSSGzYPf14kkQ43e
NsVobLi8LSObaJwtsTfvmKKY3HWDu0fAk2rG9euuDRlOJDT34KAedO5NR+ziTrR/
9kgh3Nrr9Dul2FD10QaYLulKmB+6XxE3zrwLIME55D3k+1Y2eZUbxlb+lQ+UM33X
9xxFQJfqI80HdocSmg+aQnYgeSM85GvdhXnsMNyBoFifjbR3XdWm8W7bbEB/MpTL
f7ocRpHg73/AaQwkS16WrNDWHrG9yBsMTK6WAPbQ4xwBetkJVeldXG8GVIz+56jV
k0F2qsTMmjFqAF1Eq2F8FI/IaOST2vdopqRNVgzickRsj3wLQCRrRcJPl9vLqP7X
OH5h8SoQLhPX9gUloSIAC0Dagd+sLopwIRGcDHi12yR+iafPyxYGZrO6OyE2ZXxB
TLeMPLLwblzoDCq7rnXcGWN8bHmNpiJMuwuqTlDKVZwtHAOhph0YmMDDApZUv2QZ
5lGD14RHYPpEaRdEZZdeQvXqTtrevLbVuc1OulIZfCaCShBjDoYwK2XwhlCSFwm+
6uoH5jKUO/tKqHkTOF4LlvfFVvzrHG++a6kSnpqEb2G99lpW1ee4XY7RWINBMfNa
L7F4YYQlDvdv/ONni87DcUawiRBGZ9VqRNkxIJx3JoCtTPtXWtERonlu5PkKmfyJ
ZOvue01/5g5Xk8CkSf0aUR0Z+V5sby+wBiX7YI2HFCsoSSzWBBSdebmQz5ehiwnw
6RNHVWK1czHOK3qIwfBgEjcQTb6hojSOGJkqQTIciwngoMXoL8oi/sXYaMrVmV3W
qBXoEauxmR3y6/NJJ+gEOTS2AhMDW2FFor0goWMe9EH06M9Ufhj9/i/5UQVN0TWe
pszs44zIJIVS2RWmt9+stmnJZBGfFPv+KiW1gy4iEO3RM2//crvBi07pl8ZvvAHG
HNbbWW/NKw5V5jXUH3HOaD8Aj7mLJ4udCzP0WxXZxMhSbJ/w/Ip2hcwvMGkkkF5x
+s7TnlNC8wo/QBFDHcNGiPwBhMpmXZo3LXi3KzhqIzTPG3KFWlt521rBm54WTnCZ
hneNcLaHasb+QjQW9D49v0IpKTrSrppAwP/cVTuRbH15H8+9Uk+Q525KeLeXRpoP
S+2ybWYy/dy/gbpAe4G8D9X4Z6PRMCUlf9PBn67n6Kbsnc7Z4bNq9ds5YmL6WKc/
hNg+NXg+o5baYteHiCx2Ga7ozixrS75B1BtoJKdhRfjl7nMYayUSD7Y8e8DlZcI8
6US6vg6/CVW/x3tY0ws85MRHn2072a+1tGV20pJ33MnHALgcAoqb81z2q5QTYWTG
WTqm0Il+ZTPphyaUvRdWSD6t6QwC8GE/EE6FZZXl7nmxpMhb1C8ivYeoCVf/xx6V
QNjJ8nj6f4BZWDPAlZIEtwx3bDGtcVfF51udu1WJWwJbWiO6g28bAR9HnRoi/Aqh
bKrtj2OxCJIoIzpsu/mWV/2VEmrH5KlmGAKmm5l7A4TqfVPhGSyo3hcGVzy2lj39
jXgmNtO/I59YSzRN/0EEcR0ki2ijTbcdzaAkfDpZ/+9iFeuevQV68XdmAf5BeCxY
e2ND+UH7hd53Mj/EoWhl2SaRCy3F7XU1G8WL38DOsIRYtHjnargbq/kA9MWKa8F5
q5CujUCKonVvDFYHYfR8mddrLeRvnuTbvVUvoQPgqh9XXqCk3TLIM+e4OPDOYgXh
hjyeXkGkUgZS8fRFTE/bhzFPUuH3D0SioX7tEVRLfuyH/dJ4+Wl3B/h29tQ0AxFC
gbjKsxYRqzuBhrAOOtKDxdla5BHiQ4BtPE4LyiQ7A+TnbJmpUrAI9QdVgHRAgOBN
r00PQta/nwmay1A8g7PX9dsr5jJk+SZjhrLwnLRNu1uHBk0d7gua2Z8V7G2yS0re
xK7GJz4aKmLjvgXHTh/J2W0tk9sF/wPFMUwLlIgKH63S5HJG1acmz95E+17+ZGur
XCOY+xlLZ88T59GRl6bQQ4G26sz0HGAmNrClLek79nCdXY/3JOlFVaIRksX/CnkZ
aheweRavBm6LvQXZKOAx4Cse0s/esQeQaR9rtdH00iOtpQ3/6/pSFDfNR7EgVJic
6sETJCEr4CeQJl2+WYKqz6KF1+86wisEAdcXsN9LDS/sCtOz8n0F6X7EiOGYb6uk
ghHpVv09+KWWqrZdz6vZL0iztUJvrw3ZvRzM8il9v2GWy8jBumtTCjA/oBDarSX/
FYAv8wyMvfDo5ZMjHXE1mIgmHuKE7ltql+MJB9o9VJCxLfbU8UrsOyaDCHa9g7de
xFH/mLdH92RluifR00dJ0fE82HlnCqlk6oZwZgZV0R+2qFcOLMdQ0GXijclbVfiU
l6uUomHGgZCy4W1ebCCYeLF3nYakgoSYZdN0CXGet3fmP9HMcYtuP1E/Preoa38/
NfUxeLlhJ7v8Zu+7nEl6zmr53VNQue6fjWPB47sqzrvvZYgb1fYdlHKj83Fh6nEO
IUnFGGVXjp2HN3Nzq0kH88wE+Xf0sOLpnDIgTzjlTMFt4t4wJNwTvb/RqTgYQWYp
mQlL43Lg7h1RyUDLhKxrwDPJi9oLzvTMTJx9LfbSo44lx2rOFHcv1g7m8U57m2kL
bL2qedh9aMrm1hkmrjjC3AMb7w5wFOewOFdEGgM0si6POW8G3CKFmT+GYr0DJ6w6
5fXQqfCA0s0xe8FNU7iO5Gss82O40V9EdTfxvviSP7KT+V2udlAW1UV6K9txz0Ow
9av/wMC5FN7iUw1UmLwdzoTmjCOj0LxdDLqBWbUpPs58o5ycerZrBM48FYKkQID6
7raAEqRygBCkYqlCwtNguGauifhrv1ari74g4s6LfU+exJ80h5N+Z5scNehQICQT
evdyHp7SgJx/kuOF1AbbO3WIUa0OVuY0N3JUD6WfQM3y6Pga0Rm/WKETAz+Vbq8G
5bdWDJvn8GiM2dIkxPB8sWlefnAV1LOAo/A8MGU+IHRqRzSxGrOBrcfqSPKRHpL9
QVqAb+5dhUgZHcj0DgaJhzhpXYujnukT1OLAGgvgY+eDpqkLvD1PsfHe6ESH4vux
230KtfCKsGMdAj2qp+1E3f2ioDluHPyx6TRrTIwc44lBLGRnDbEtILyqy04A2gCf
07B85LGoPZndoHpnjcA3ohltGxgvhWmomuE1dqb5Q7F4KuC4XK/h9xnXoBB+HaIC
GnN8cMs/0F/kHJtslIvXp8UxwM3qkDpib9R691aJvzNfZOJo5CWrVwcFQIk7Wy5c
+7f7kxPP0HOWnoq1qqMoVLkmxaGPnJYHQtrKmPYzyphwbjbOhRHEHledEdh1DEh4
trirwYDt35GK/eu5kJH3XJWL6cQrcuJ7quiTmNYaZGWKBc9fCkwsV2MATjLgSHJf
G7VatZI4TUcViug/Vvt2pyio38kSKT6ItfLz9hzojxRK41YDh47iSCewFPeskAhi
FPiTBJGb1OaICCWl6Ax+r4BUo7cpm6hoOoLT9KnWI/QfLWzG/3VZk7EQknngr2qH
TlzCqSgeZiPFSqiETAwLy15cUq6HCS/cp8M5EvPvVGKH7e7p//gabn2MBRX5VjHq
lwIgN4TEwwvsdtbXXcvByafGzcx+vGCmHxmKBzeEwYnb6VqfTV2ekNnFrvE5wMV7
tpKZAk3xFzWa3Ar/8T/3xjXTd4g/mCzqM6ZOkKAm03jbNzpRTqxp6SJBbJREgINK
2GwDPTDazD4SkYsJyMZJQw6WggWkH1q6keDFRiPaNvgiqm3TtUeSpVeMu0+18SsB
7WRCtEaWusSa9LApNReuy4y34yjtmoXxHfMkw9zJgIx4o1ryNlyjR/ifWNfbqPB+
wWvoXu+qdrjaXguNNEq+UeDQRPAhhMGoTlmcZB4JINAEuVR07abJxk7eeYYxyyYa
QSrdO7NGUCDLik9zMQrCUuAACBKBIwpL3rUWNhggW2JyphCWTcw/8TXgMwSQiJVM
iUWdc5ERao8jjrbrgqaWTRZp4Tgu5nDOzsGHlhrs3sVliDdRyuWHN0wHFBXP9wJ4
QdVhXd2qDZB5xjJtR687PyKutgZ1BHgMMI/X3LE/VUfrMgsL4lnOBkrhuZczocUH
kUm+lL/8BwDVDpijNYx/DlGL8PF3DDE0OpsQouV5SBPGwYLvnSb0Ta7P8qtfmyX3
iGor43QIvtGE9J6pW1Ht2Iz0T7WjQlUUT7IA1bu3gFib2NZpF0n6FE1bQAphRJJw
NQoXExApU/AS9cRX50w1y1OtQXEC+tZhEFcU5CMYkKffG0IBti04ldAWyvPcuDZE
qg5Z3V2yHA+LJJCe8mKb96tQFPd6mABBrrGwJqhi43dwAIPbwYnAkcLKUFJkhnBl
Axz5x6BgH118LALWqIW8jHiwFmP0QyWT1DojWRZfCIRwNIWz9vvR1mGNdgvTt3ku
0K1rgsAKbuEywM2j+xryFd2W0OtYG8vAsRH9HMBO34EsM8+MqLWIV+l/OuaUl3Xi
gUx0712IYET+oOASjN1ssl9pL28MKNg/Qy+eq77mu8SozxTHCewWhIo22cnfKC7r
xqGBqgybxfRJW0f/j0CpkKnsKTzGSUTyxlpKbPA6S63wPC4t4EJmzA7aM5K9FRBe
PEJylOCTUdoSYZE5pSa8ZebSvs+Dgtt69rz6TRFHYUVqMQdwuKh6wlS+qIG0ufqn
gMDzT9QznbqssZZAWp0MODh6FqUcFyba/v+dDRfppEIqLdeZsNLnqsBwNhgcUNtV
h14Zvgng+DEiqq6iYiOsm/6xTQWQ/R7Hy1fA7viIMMMa8vyAbSJNYr/gA/+52O/S
oZ7ZYMA/Tp0PfVl9099Iay4nEL5BlIVRqaEV1KgDi/o6lC5xszDcGA3GGzAiVaOq
xcNNjXxBrM4fiUhQvL+Y0fCp8ixSqdoWUHTivDjQ9vvPrVGRF1mm0EzxA/ZsMHtq
o/xSzAwU5/AsfnGQtYAS/8oLI2Hr0Cd8rOebHn0+jryXUR6UIlWOb9ktW+t1FpGL
ruB2zlkTS3OPZSjplK5Y2gFd1Sq7Esur6jMjECBEXUytV3E2frLacyJ512AM+Gc1
Ho80q3z4jI2WUxREkVnKPCtvv1cWxsYlU6WdP4fWlH4UM4QArPI2k7MniVWLRUqA
kLDM0o/KH9v73hxrjThcwXOTVBTuw3VlDxPWnKraDEUCNdPwWUFohYQqVno9oQrO
fe70o4R9rwHzfbzblqQ2Yh8JQ/Dzb8nOLsSSnRRrAVXtbhJ1koMQqqbvjvJ30NSu
0wpHl5CG4wqjdG0vPgOIMxsMgHbIUMcn6wU/DFDxdtlyO2pV5Q6ud0Gl8f14VRbc
4jhjDFxZ6KQIKPUwKjOmdcN2b4VMKvjLXUEmj478nTyjTmtvgVLETfV10aq67Hso
JsCBb8fUgV6sd9whBRPwkcvU5cH0wIswTxDJzo96kD+tWNv8Ebb2s3EpjnV33g4Y
ndFKCXq9YR7jP63kNXtRq9ACzEyfL6lLMhKRwmMv6d/85E8SbgnVRPyEQovO/g0y
vrf0R0zzdF9+52OqVBsCKb3hR6vfu69gUS6DyW3r7F0DtMBAI02Xd4EM4bvpyqC/
v7kzjcqOzcYLIwpgPwza0DboLAN3AJA4UFj5dLXWeqR9bV1f7jend3IbYa0o/YIf
Fd47Mr4FowN8BFkb+dSzOBSAqp/lbDNIYYXDKzpIbLIk6QGHeJ6n/VLyIw1zEv40
6mu5RNsQmuZ4dArraDq0DvJ1i+SCgRtRslmjVJx5EoGu1xqzqO0eLxhfT1kPnrhb
Quxu0QSv5IWE1lqw3zUw71dNJ3f/N4jIzSZX4EU/FipWM2pWSxkPH+GgEarOq84M
5jKBp/49ny5LIKvmnjTlErg1B4v0Q1ZCh2+AfD3BpqCXsbeGd2dxOpdLVFNQUTfL
y5oge4v7Kj1p0EhzjQ8QYWhd+7N/cVNvWPysj3LlPbrAvcyAs43hbolFMcPSltv+
xjFVi1TynCZ8q218xMMUASP/KAWwsdc/Mi9pKh3A3hePawNuUekYwl2qO4skWF5+
6c/pSQrFk7wo8ER3/R99D2VciSw7kcAdBGABmVxZCY9GzcEJ+Jw/2HsceLLN2Wkt
mUDxL54H4ZT0O9A5PDoYCODNo5TbpPvvYCli0PCv7KadgkJMTrmj+GnReWIT0wFD
wrEm6JEiLIrxK+bcoRdwjs1acxf/m/xbQoSVThMvB3uxv5soUqGrq8bpQRe7G/mF
Ped7Ird8w5Tlo0lzu+1ULaKKQ85Gc6JrS6CC1Jg8gtDAA9WdKnezDx/ANhZ0sDfC
SXGn1svfVEE3mMPJibceys7uGvI3KV5DOlI6PpgjEKuLQXtHkj1aZbAVbngzeYnA
iYpg4PMW5ZVDliQTXUdmDauty7z04pp2/nJq2+fHvXGYe7oNRHG0F5GdLiXOBQtc
yYH+k21HcOsR0IcX1uxTaynf3IlzGMlAEk3JHaCmWjBbwzA+MyedXwONkdVEs+lu
H6Ju92g2hul08j4hT2uzBoH0hzNnCwYhXs+VnsUEuE7m6yx23SN4vBkMOPHKudb7
weS0o4nNgbA0U7nb+sr2/FFqBmymHu3YMpk7ilMDualI5khphprDKWgW1J0D8z9y
gtYeS7G2uDnfv+iTfrm5XvIk3huUqawtC45iOYXhCTSvLA7jyWOgeXa83jAoeK76
pwo7zUYD+Bx6ONYNhIWhE+a0AmuYtcGT4wLZ5YVnOad9JKH0ecTeDFo8Zv9/L+Eu
P4tJc4ThgaEH/d/GYsVZJnV+uUhJo+1nIK9x0cmAjaHbMvR05DQfIgP3zrek3cef
sydy6QePFemAWYyNxKCHX/8Tl3CBfqmmK4hCC0f1TU/n+fbqwkdApDdg7fytXKFS
LW72ji8TJ+Os9Bga7p2R5/ch9OjBjub+qrstdnECDWRhjhCQ2LI/hUnLjmsR+3KW
2bLrOfCy/Np0s2kF/BjHfGqvJkiUYxTKeMLGNSkOYzOjKc2NzhbmbjlXBb83Zuat
kyefGAYBzC6x2aRcDBkFwJzjX1RPFY5d0PrrV2wT3nqVlhDDZkVihfNJJ35f13Zu
kOeAOnte/cqkvPQ6tAXj2IpI09h5DDPcxQkYsQfD2bQE9Ple7YiwRfelPBkEEpIt
0muqAMAomOf6VLyAOvApgmrUfPN1MerMFmFvjncJlSNmg9ukYMBjv3fbB+LRPlKs
gUbIl1TGEfgryzgxz4HU7AM8mHxCX91ObgZEvrAyrKvDnwjH7dAPVwDXEChoRGEa
/pHi1RkGRcU5dmufrORycbYZatDEs7PxImVST8tukdVsdmYwIzdgCKYI2FLdHDEo
jwgKc0uijAfi34ZE2kIn59DDWHFmIB1GAGEZBE4EvvzuGd7XQbXOExj/4/rCm2vC
VQyLL3IEjvjUXi0Zl05TCbkdZlwZc8hXR4zShxJEbwavBvXpGC3Xuep2dOZc0gNt
FHDSfaKU2kRXzzPf86quG4P8jXmYpHCo/Pp/LBxOyOj2bOSED6SDmVv3UnPwGG+P
zKB0IFiHaiogfuxMeknE0EKblUPOsTE9A1kW5LbHo03IVZSNSK36BRpd1jOFBh4g
wRbmYiXzLPzZx2k7XO1GDuvp/FWmctGxu6Ed9eQAFbbdg+TPIc6W7fpwbJ3U5K7T
pPIe8y77ddp82MW/9E48NMOrZhwFs1yAfz/BEobh7ah3dczxH8UjoJcfA6Aax2AF
n1QT7lsUHBut0cg5aYmO/y1HJ0hjEXrWxkkFfkDAUkEOvZ8j0JZw39kz7RPHthh0
XqObyuHrXfyZceCpeQY3mzsiQCr0s28Ti+9tRW4Ptm0KL5jI8tSatUzP/K7E1cXC
x4maMDVRalhTupagSMENIt4MM3IX99eVCC6V3E+3VTs06Qj30Z8/XgHQU2dbll+4
YrMFnR2jJFl42VB+ZDbH2FZBJ91+02yRLDUHlp3gUC/fREOkEwIAlelqJgHPiCk8
SReBUWkGCOkbRXgQxc6EkVOmer4c6NvTOSHgni4iD7CFAOnJlanUeDAGH67nzlAS
FTCbZxMIIQ2dBtC+PlZ0Wiairp843ldTF+wfxofXeEH24n6rPyuWgjH1JSE30fik
9EecOFUw4CaWPU1hwjjBjiI410rICKh07ajt946MqDw7L3uqDJLRNzEelusmtQ8v
VTXHuKi6LnsKB1h1h4A1mpUVUfYC42vjzmElqr1cLb817us1SlS1Qj7bcysAXW9O
kI7P3R66HVid5EfLCkhrdtFUc5O7nAx632IQ2dh0zx/IHtVtxsy82W3FKpah/cJt
yRYeJYHr96BgYTm4PDcwjAp8A58EjsmMR0r/95+hL6SwUpUr5GJmouDS/+qwNGNy
EblJUxH7fFLb/5vcNfZkYhVMQk5N6zG37ir7d4iaGDNtQWCLLEzU5a3NrYfRq1xu
KZUQ09Kpejq/itXwRVNqJoWRHfrIisHp+OzDFKhNoqtc4VKu5xnpbNcDNMikmU0q
fH0U4gdA6cBRykvg+8xeqhX4yKdmZHERWaCyDHK75dvHiFGGnRzLtVBNcqqxyIcB
ViKN7OqTULjLcSI1xNHV4SzblvJkSf0h0K4skvOyO+ZUIpu1AQeskovZTlJNZhl2
3dl4XHvonY7keRgJROnd8yWckGXVbnYMSyoM+SDjs94OLHTaYVd1QKmrNI97lJ8W
zTl5Q7rKFDwXAD49Kg12YrxAiuROb9ghrCbmIpBcoB4ncmizrHUYouH8uHM5ISSu
MZ3rG4Nl4R+KOe5IDxB0aEw3jDxjIBl1XPPkdyGgtOYQOQ3W6MWy/ePUp7F7f5Bb
NuhAJIyCJ+4cxijnSeL4SocB9fXXZC3dYy1SmeE1Rk35maLPpiXGX1ZGAzfVnrxs
w9qTvbGa0dYD8Eihr87NIAcVirEkkJqOEcA1D4dhs6xYdrnj7BPVw9L/fMTrm1yx
JYilWrQHHQHz9kjuxZpHSLSHvVg6bk9qxWYKd5041ClpgJfJCTK9bnGjvJkn+Yd6
nwfF8dS4uU4Z3rHkvJymHInWWMhdBnc9xzkQwFZQlV+xqqu/WVzGhDbasjCbp6Y3
BnJ35yCwKxxRUCbBRyZ+N5IOMwMUSW9l+9Vs/kQox/l/wvztjg61/xH1tLYOK9ys
krFouocc8JZRJMH365mZ0lp0l/Vwtk4+plfrq0XMNgHwK3F5jfuDmqzqxwvBfYPM
1RMRkNK+WnT4VIa/Z7SAHWuQrZuPFmG6jv8+miPEQyfV6lp8e4Lu4KOFQH/gA81e
3ri48Wv1ATCD9EgAwJeBPIk2Fw383WRzTGxBcubWofr26nn194jrua6cIAcM9DMN
wnkLZz+6wbSJq9DEBu5zdIx95UPYjpoKc9ZjBWybf7hl9PFa5ekFD9afwYWv7ihY
q6GmVw5LPB8gXNEfjB3Uz1/mNCAmK7LDUL9ZKLJnmlgK5fkxNE7eslsTkJnJHEt8
07JZQQgJYCbcTXMwcMF6GVKJfo/Pk8KPZ57htdQzHh4wpB5jADQVxp6MT41DxYRk
N4KOF1Zod5s5K5skoqh/a14gtA81rdeXMHKeiWoeSHdHlJbF0ipIovJJkxIS4BKB
ITyGqsxfyXZ5s+1X9EMAiDM6MJl08AwJPAyeyDA3WXfiOX8Aqa1xoj85lARprK+c
i5X4/LTOD7BDksfm7k8+lVLmy3+znHdC99gNWUPK9hzrnAZOYqEFbryYJJAO516b
+8q/t1I7lS6r7jih+gGjh+3iRQVZV4R3ADvbzaShwgrxYhHXI5+8CX/UQUktmjTx
RSS9CAUlcWvFewcyKU/h7z4HDg7lEPqIlOYzzqQ77qkaMUXBbafKmRBpz8JFQbYi
Bjmkm6yFk8bs41V70fKZkZfUqwP2QupqPphC3TndVHkojJF9VlvYv7VMUDFcJdcB
JttFdrxWR89NXKe/QHnz3MbVn310UQaZMEXHfiqilz8BnDGtR7J4UifNVzy1/IJc
5i4ygXaC5bvLk5tLa4HslBGEoAlpRAeq4wH1H495h4eHUBr1sCwntE9FOO29eQp5
/ZqQlexLgQxcCbU/kz3ikLnrSCkeVT4fB8xxior/nu5DtaJlLRq9H+951qDoNU+4
WooL8dH48De/MWocMgxL90fzwPeqGxgOw4nMCXZXi9Jy0dkZSKsBPleiXFDXtFLN
PQQsQwZVCoLyPDtoD48CehKb3r9/97338dy57cHYrVsgUNcbnHSQUmQeVz2dksoK
Mdkqcf1dgUMB22hpPQCIt4fc6Aa0SX+dr6SOZwX8k123FoQzyA2vbZhyhuVApbk7
+ASe+BLuUgo8Lfat5P37z4hCueTfQxkFIvajNhj6nZEcy+rsQOXJnYwX7Stv2ws0
htUtCoVvuAqPgp1fQROqfebDO0+en36Qm3aau1jY1V40I0oL9m+E5tRhGHy5jwQI
nrLPUuUfnHo5oSkn53v9/+QRI7RkSE4kXJ+DkOgVBJrHbi0Cjz9mCJtcQsCpc2Pc
6joYvg6TM853MsiPYpaJ0EmIqK5dsiRvxdkPBkvQxqYYO6W4H6FLvMs9toL9VOJd
1h0UqTby/oIilj4yKNm8dHE3H+rwdv/E3LAKA9nDPG/Iq3JIa0+4eCLzyAWG+iN4
Nbdw0vbLZ4EeRef6my12+2Tsp9ZELAMbjX/8B6SCfBLZeNrtmzGoRjWZSv5i6dI6
gnbfx4iWVRaQRv2Y5T80pZSQfWf3X3gNVH3RXuYtEtImxme6CYpgozqiICGu6oBM
vNiEyB0LRm8K7Kz9jYo/2eFS83pWbMnROj4LbKeww250aPaipqvAnhcwFSd+i/sF
YSdQAh1fL5JyZ116WaKCKV8x+zD5ORE6zWLdhTo2Uv0XUXpqIg87cvjQa0lPqPdL
cA/IhxFW7bNdj2ahl6rVkvzIgSY09TMgeb0Sm8/Lx4lf5Ar1uzhRb8Teo9H82w97
a+K+XpSyw0RVsNmRsOQXx8Wd5GV8Uhvz6sigbyfmRI8OLFppJwN/KIpc0gpvCNEo
J5M81CvsTsR5YKGJFsCSP5/HP19cW061wLPHbe1nHdpcBHyb5POsa51U5JSeEhMx
Tle4E8KcuoG9TzxrCNyofS1ZQzKTIwMoX7nw6mfSrwcfayx4oVT2CsWcMqbezjlM
swwllXV2L3w6qV63G1n013VY0G5dXJxrZ7Sx4+kyMYJ54YionRXSeBe7nWKIAbDm
mzdVe6rTp5iPg4BMvijubDrz8RiybXf3hgEDY9DTe7ly9V1wCXFk34Mr7n4f9yu8
mz5T1t+8C+eIRLOB0sV4puDi+PD0J3j8CGrunRxECnCHtc1IQ4tWmHfT2pxbRb5B
lR9oAlOWHXoXaSEOilsoNTFQB4uYLfbNFU2O8oHCdPtKx6EfT5D7jWuUv6qgpw21
xvWJQAH7gdLY6FUqsm1OpgyaBoMpgYcsMmaBdWd71QmbVt8qmQJr38D8G1NH9+Rt
WmFaiqO2dU4/5KE6m9yQAuxExMiWr7PwyWybRYCMGemstyJqSC1ZoxgsgUdkSUL+
VmOS6t4XQI2bnzKkKk5CRPjYQFoFj9AsWvmmATjE2RXq50Vm+1zAmg3lEVpKw8cx
eUGlPQniTJBF9Fy3zh/GB+kVDOudOOIPNhKfstFL8kOaX9LC/HqrNxMt0y4rIqpw
dHhYqJhCIpwvCb1BlNkQGCXXHXJdMbfa0hgQ2t72840Z5bgrr48E08GfoXkzqDwb
Ijsxq3QvW7R2p+5ngl/FjCKzviTtDoJybk87+AAOL+R7irDKtEFFdJ64+rbkka7Y
6RDHQcf4Z+42r0C7tvL40zvk4piOXAprlv4O7zx10RDqnas8R13GXQPTtYTiAWU+
EsidHfDd7NoaL4WJR0YWNCHnEglIm9sijQAaCJNZokKUUIRZq3kWsSmhMnJLOCXk
9Fn0tx6LL4P4z56F1iPj5Oh0vuOo24pQADocmUTGIyyNQw92+e97VAeyE8KFtFPp
xBpED2gE7Wg4KgJTPXeyqoWR74n5DcgusoclhC7Lb76Q5jzXwckQtGO3XJcb2IRZ
QTwHG397ebFM3wyXBZr9QIpVY2qos2IW2hAnlyUu3IIWjJqWyEnfZFJ2YHOWwoi0
n80JvQWlkvk5kpEnIG6EXCwTQ6We3d5qGDhZ0uyvaVfUFAtgLjubilGcbJrezxs5
7YQQoKdZXsoDX3XTdWwrkBSWhydzcbOOQbzzGHNgpFndOXRVuhAuI8+q63l4HLm0
edOS/xi1OKs+U8X2HoS6Jqg7jaO9XlmJjuRqMCMH7DamJGjxUW0K3p8yuAme4PBp
PgY3OMr9YObNrwqrngDtA2lBJtRT0A3TTt7JSWJaOh26ZiFQrLSPt0rskLvIqkBq
6aRFHyFr7SQK2w8tDEUfUkv9Wx3pQSg03uH9uB6czULCfjTSLGpxOfm2T+tg5KaD
rkunplrPQo0OYiPzrXMueBpZ933Aa+nV0yj4JPiotmaW+onYwOtHpBipUHJ2kyLX
b6ZhGvOqZyOOuwUWNB9ibsIdeZGGUgijuyddJB25D/UkxGntr7m6qqF0KGQDWqF0
OdK4KItQUiu9tIhwQ7Utd7ZORPNI6ri+85OSOuaUN8RHz/bfPDUHcrJkAny19xFV
PeJnpvm6Dnx31iVQqLAKgK4V83YZW46LG3upclCRU3YZlG78YcDIG4MK5RGDMQhQ
6K+QwPMO7Nhbha/tM3YE3bGcHGvzHGyORyOLb6t0ueSVQ3/WL62U1KhLy4nIE9k4
LTiQZOlR0HuB1I1JYl6equq4EeJR8s9N94cvTJJcRqdYKP0Qv2LP9/BffOtONazL
LHAdF+EQbzNrUAB/fIydtnlN1kYUXgTvUyOsOrzrTlwuibXBdaLoGz4mV7U5lWhu
NIm0rOYcSu7qQJIZ99/VKXW2f10r+sJx3UPUNY2++orR5TeKOctcgwNvrAJpaSc1
k07GyXxLglHQ3krUZqkKjmMSyWYOiTHwG/xs4N3GqEMUQflvr0JvYVtEFTY6xjJO
bNNtIdjEtX54Wh+/E5osr5gfSo2tZHkROxlndBn44nSK4/2PoiDJ0UFkfkx6HT6Q
CgY7Q+iaF4qIEoiUuixII4evfWATBYuiosiDLA3q7lmWMcl9T1YIyu8WXONwlh7l
Uz3dH4c+odkMe+TkfKHUxkcFIjDT8jj1X7XmCDwTayJKMlh0C/FZYPpAQRuJaTZE
rKQ8hHmWlvSY4UDtIjvXqv6bGZf71NajA1/L3k1L2CHsKMuzJIgpYG2m1qc26y0k
i27q9O6k9tGLj6ozkDHjFYv+4qxzMBOElvfeaUIFh1BRRDyR+o/guRcAqIvLJyaI
i5mae5MT7jQckuGGaiDQCNNXcY9J+3n3viT14V0o5vUuNEH2z6IZx7Bnq0rvU+Yr
KEBWnB01/ta4uTzw58hyiAudvuLVM1WeKwTMZMlU+RZ6lonhs5gM5LNYC+tja0xV
C6VNHtC7WDGFzf4cXDQKOAC2ogXgu1bdWFIJrpTfqETQcCwHwr1IrZ+sz+WsTPE8
fMJOplLzWMGaPMBwSY11ZwbAQEUmu5+yQN37MHIxAP5HF0jgeejunOs8jVcBYA9c
miHLLuLQfGBvXlUooFOF/x4AJsk9uHWosNRkesTvouWZzSGTl9RCAqCU2Qke+474
ZzLxO7aN6cSHWO0H0Z4csq651ozX4vBJ6kjOVUDCLzmfPbbe14FXDybqlW44MBq3
slF5dU1kaBvqUzrpuDlexw9mQdq8YSbF9dmSVmwcxu/+TBTsC77c3KDpe2S0RZ3o
d4jHbr16tzOTIJ9rByOw+OxNoqPm66EALoY0amQaJASWtu26eyOiIPCDgTA4Me60
ixBMEnyb3sFugzZIPbaXAPYjcF0E7Y0rnd3cH54iEm9r7JFzpqdq2D5Jv3PsVYRM
udyBUvkbg19nlyAEZtmCFrQqNGqio3zHCcFZHUrKoiHlm+6B8bMJzhrRiVwlWC18
0N5oRQnb4Dj9KY5cjqrPGNE9d59eslbv3yAZsCAYK0834ZAF2FIJjUVqosigqyQ8
taRO0/3QyS8ibKd9YIe9HfcVIHD6310d1zJVxiw44HYZG7Qf4xhfWM6d2pI7XgMJ
MkWkqqXKspoKf/lz/iLdu3R+eiXIuKKnABejQN+w6kg4kByo/Dp8f26eGXVEqep+
EgdB6IxdpYsXsaSvan2T0pAExfAMjgWlUT5IeuoMwym4n3JLjHGxsFoMJYWDJwbf
cXaH2R+YsNUIzU0lV2YYSPtnZDKR8bSpXWdeMf7TiXAD/QK0u9AG+nyJeuqCVbBT
/ButBxUZdyd954w5nW8izugFcQQQjff5yshsCulRZwa6mm+MihSUoICEkAFzSJ0A
y8PjZttDOts2lcpIxuhF8d28FuxnNKNbyFNoucW8IqtNhv9M3UKiHEbB35ebfo75
k+iFatAbWzczb1urR6aB9W3BJuJScQQHvlM46aTaI3xEoeUvp+bGGZKQRR5RpZZI
j9vboXzHQYMI6rCCgpjU17wgsUcZHLxk3YPCS2HHnHoDt8dbvwSPSafpDfOhFAHr
qQn6Oyp91H7UbQdht+mBbFuQph9EBtXL6wos9byRL+9sZfKoz/HBPNbNkW1n82TA
eAtZBduGYtaINRTjrTQLuy5HkcJGg4CwyCmTD2T3tSfG1aT2fkVT9CNwOZEdKaLz
9uh9CfGIqe56erlIs+t5GzCfQ76ev2w+azojhAAQyqfRfKUQw81L15A8dnOwXLmq
yK8UONks2F/JkVutUMnflltLHPSVQCHNCdHb4jBiOUY8li9y+hoKKEQfxW41nwz0
iF/h6kAZbdo4M4xa6ZU/+TUIdWJm/ODVtbwYRXZG8VePjd9FNtX41/kcUWPqwHPq
OBKcB+8QVmVgJj/+wWX/ZEwxrImziJArA2FFlRshLirhblEpggZPTaUb07lRnbah
W/EXPjGpc/Ob1G+xSUHmxMBu3uhEjCN1pZeNhnMouhpQlk8MGMD/S85YIgPJqV8Z
37K+SMDC8xPYWr4sACCR2HUQMxfGZH98PGtPaZJsvtkT/E8KPEsgMTKqwL+niI/q
huAZ1obZSnErVXk94TNnSTfEAfZED3HAI46zYmuIAHKbl5F7iuBLK5aTbOyi5uWL
nXiJ3yi+9PlyNwLv+zSYfOG7XMIBxEPUynxrtRlwQVhQ3CN2eW0ZYRbmGCU8+xQw
xmq1Mevyy83TsKmWp61kYrZn/EZWFrGepy7MndGKFXgJhyHnw4Jclg+OfWfvogfB
9bteaRU6QRvxB1CpipPQszSD0vXW0z/MQrVatZNrZXlPrBssvfnbABZMxiu08p2p
QaI3d58b6kl2O+rYWD2ph4Uv5rgqOE+H7mKVQGXk9ZOvqZTgNb8FLzwE1cMYSfPu
ncgUtBcQ9iwCgQQwZM+SstPVrFcpWPqqui4laUI0eWjdkW7qwgmiNAhL8PI50j11
Kh5xnLjdOLIqauLq/aO22F+47WkBbRQAJLu/SRy+b9iEaQxILNicwNgjKTScqN8X
wQnye2lvcMiYavIKCwktmvtbKzfwS0IQz8ru5HH0nXpVEueaEi0SlCP44P0EMgPz
odI8ZMTMsppgon7oS+bvTMvKjSg2bMAfIsNzy1kjP6YqCyka+BrciF8lOy3k9cTz
//Wq1p+EEURRtfHf6jEEfRfqHwXeIhd4ykKEA9lXd10tOr6tIQBlq+/zbj0L2DMS
g6U9wGE6MDRb6bW8FIeoTLIrvBPjOO4FlGj//xmwRO1MaqnLw/0MkyKe27XNk2Hr
ZVhvDVJWa9QbQ6UlEjtwIDxh1sk7doIpV2QWfReCS+yLaQE0+HnmnGBHemWx2JXc
3Lficd9IIZGtyyw53hLMhksheyQKOgNkUgqOWY8zmgrw26bF0oGutqydpx7h0tuC
1RxpfNDkiKZynNRwyWJCUwbH9BLs6gLF+OFtELJHQOBpvWK/WLcTwdzhGAFEja44
9byqPojtbV7qsyjERtUtULEn/i5b7qfzOl2q3OVtwkvPu3VtxLy1211HjT++d+Id
4kOifBjojKXerickE2aOIJ2Di81jrGPY27wqxLnRqdQYkCQS/OBGQO6t0Oyu0dqv
pcRiO94WbrNPeEp4UqUG/UkgJiwSbcMqLR+4X14VuwYiUT/yJGa4k1FCpF7qyj07
QxaDFiU7By/6E+RpO5q+TfOlw9RCt+ZJWNxB9Njkmh7S2LdRmatItuUP6hLt+aQh
VyW5cmprnmcOIrQRQNdXijBa7dhtqOS4W4x/TPm3Nlhof6WEAiMqwKTRJneEtwFm
41pcTIjmi+vZuPsjmOq+zH2oLgqoEfLc3zbCUXqHePIaA3D8+NBCTsDUUfnpSHu/
i6kypE+IWJ4q0ByikVdaazWoKF3NATQFimPDBTKIyAlTyBd3lKfWf6z3/vMrcE4i
jFXmGW7LkwTAH7xqoxN5T+zQtBv4PTwUNGR98sm9iQ9/C738tV01N0QEbTrmbXEb
RBr8cu2cqNfj+zPQkeZ8EYwrHFPxZNlTo0EhZSq0RJxJaZGypC1pPH5EBxpfCJez
KTmz3uFIoJp7FUxSnrYtwdaW69Ac56pVhUBslrU8LF3D56+PK1AFZdmrVMy0IEEF
/4QzicbKfcrXlCToq8N/6824LIdymmh9hPuNKPXX8jevop09HRTQ/QC0YzkFAj08
f+UsjoKvz1AOt6LoJE0OIZSnhyHQjBUKmyFldJBPuybIk33veifDe281mhgAia7K
9qw8471lB+WFEWT50GZZ3XRjZTjZ6KE0Z8R+UdaSaTYkhbyZ5557koH8q3rRe4kb
mlqMAvO+aQhxk967l4+c/BHFBEOkJsScm+MHLapr551znkyo8inlVwhv+Pi5qTQS
1GejaAcJ9Y0n5KAh9Vnf8yKaaBs8I3RrJN/MknGlZKWhfHnYXtDPd8GDdX3j5sUi
XWd3UBwLjtlLNLoXNxZ7O6tXUeG8yM/HPy69lloMwdOHDeZJ2fRE34e9R0JRgbC+
5z41sstd6IMs9W9n1Yr1S1WZ3CY1wKjoYlGJBCf2XO8fKwhJyL/9eo5h/Ne+rmGt
zu+Gp8/0JdTp3AN2rL8QKXT6htz7VgF9iz0TuAsvvIVqPdm356Kt5HPGwYnLtAAf
3sO5+Kewtn4gaXZimi4bshjPsZJA+RmSlXSUbDI0GgqEba1WsEQ1j+LzkVvALN3i
9MrCpMjJ+T7fk2FhsDhr13MT5CR+HPOEUiKk3EvL8mHeXDoKrFltJ/jq9z0hMxGf
wydIpjeiVPzNZnSUnvzWYDi2YWm9v2jEKmMjrNLckqiqJk4eb5rK5skOD6+SnwUF
t/+OB0CPfZ4v6gfzMvbKFJ7nyBBImGb6HAtJVAgKCRn5n7d5R+/x2/e5Wk7qj6ET
vxWjo6dju+sgvCs141+j+i4agPGWCt6UxRgiFULHXKZspcaAAFvvoiDQgT7MR2us
cZ+E6o/ggbVObIEZ1r6mhCnfdcsn7xxzJkQhJMEaX0ityouirDgZA0WF7tNDIlhl
dq/kKVz108+Ud7Ugr6ktqFcKDTq6GxVc/yYImBzCx66E5QCX6aLmSkoHyorJXXhg
DqQfuiR1963Nu0iZcXm/QZAGRr43Zm+58Gz/RSP5NMGuyrL3Dv6dbphnDA4bALyF
K5UZQEApn5hh5Q8Oa71V9HwpXT1w3WI8XBDC4S9JJN4Trf2qASN1rwuCop9SX1fG
ADwUUMppgO59ZeQpBnShYcftuxJMCdL1TiKcQs0e4hSMT0w37dmTc/FNpJ/uB0hS
PdYFfiS70bijSvQt1CZo27i2ckXPJ2Snrwp1LPJAzZJHzvmYddSu3w8vIPkxrZXq
cbLK4zp87monHWFDlhOqfGF92Ahyw4LFcE7/3z7mTKLBOVUofolN8JPD5PpVT4BG
bFNCj86j3PT3Oqkae6uuKb566W2ndYGfOKHIdA7h8TXJa28NVQC7qp+OYJNu7J3l
OMNMVxgHvAE1E7uhjiaWAIPPtlMKUcz39G9aTvbiOUDPXWnRljfDkdDk4B+LZqYy
oSFU2YoN7ZR3fI1FK5A8Wt2S3RpNknepOXq185QHkEo5rNE7qe0TqaZYtKj9nB9F
x6yurPGte03tKIJA3E+Sr4GdI/qlDiLMX+450XOz0z+GrVli1N8BNhOzYdYFSk0e
rZLxaYroIZHLIGJ+NO8d0XZRuItm1VGM/l8KditS7bZwbA9Qk/j8K1aEI4CjnksJ
BYGPNmb919cyuHHujXAjlg3ak5y2stfwqw0Bp/CIFQvNK3jzt9M4ryMT9Wp+UhaD
3ClDpDg191MJu+zn8vaPj5Jb0SVRGUfnERzSlWynuzYpSOZObIwWLINDRYVSucby
PuWvHkZhbOJksiVh24OWiBXFtmcHfHY2VK+rWaTZonPaSLXjaFuUh8uIyubbyq/A
hE9oM7DYAXzxnaqgMksoUdyzqMrk7IzyDUc+cEQYgHc/skEPqreq0H+/gAsYCe/a
CZc6wCv9npQNcIpljAM/Au5NNxoKYz3NkAzMjE9EpIifEj7Jre3A8zHFbj9LV0mX
zNmgcbX8yoBmkxJoz1zGNwPMa2hHPI2zV86qUE2NUeUGlgbabkutgI4Qo9Uz74Mb
H9sCOSJCoYdJhu8bxUsurUyNaY8Zc13xs47e2ddZZEuPW8HM70Qib+9Jdf+WSIft
B8Z5524TQKpzBqvH7CH/TMAMckS/el3uvOe0yxvBCMASpgwBUCi79oG/jxIhE17t
8BI68MbGhtfZAElg9rcur7xImRxlpktyCAmHotZNqB9jn8q1D6ZWWFTDxglewzAU
3w5dbfBQamp2veCYoH8TijrS8lDxo+9ejhXgAPBWepyTUxk8BV7xWTeaUBmTV5Jv
eVZapOFINZqwlhWwv0DdfQxs46D9ENQkPHU3klDBoFwuiBayVgY96S8prrMUllId
WfShAt9uXI7w5avD9kvnP+o/dBOzbYd5RH5mUke+4M2res/mkXKcvRmnmTZpPlsu
qpizlxznvnScLneQ2hNmsGWhvXf2SW6xUijmgwe/eBplMe6H+abGXckbjf6ek/C0
XYoHcL3oTaPoIYSBasR+fA52E+5Fe6QdIvrfNPNh4MtMrnpsWtVuMfXJUw3vHCtB
bd95QylH4JqtIwKCDOVVvw7srX9xKAqMX7PNBsJpmT+8iAEPKv3Ea6QhkmHxNedG
G2pjMv+55vbVuCgxlrRB4Gdx2OrfnFL5+EGMZjOYAtPUmW39zNieoAkuj3pkxGJ+
EXUGmUB5Pwl/jbhMcjujNlPBGpACB/zuA76TxZFWSaAP+mLLdqwfG6horg+B3fNu
10SP9yzdsPAPMKEzefrfpaV0gz+OaMA7uELq8I59TUsmtW/wF4fjtjqWF9PlJvT5
kMNRHU0QqDxuF+wlsyTuPW1ZiWt7zYCxwfu3BlKAdfwfpKsEK24+xif7o6bFKQYR
xO9h72dBVizi7uSd7EHYWSerMPDZaD8o6mVfi3edxgd8A5FQn1SekUbzTDl9afEN
199YNRVSILkt2Zkho/e97G9iHqHI2MWRnMkii/TCK8XiwSd2ELOd5IBOb0AtaOnp
rUcGcJStmVv7j9DHenwEdPOsKyY+baCQoocjE657wEASh0RQ0kTFJlFZegrCA5kQ
Tt+lIZ9IWc9x/7Ax8+NmPvDD/5WmDo/QbXFG5Qql+nwBjm7hpCNwAXaPcYHxRm8O
RYgt8qpJIDwqUPlimyMnxSDFRK8S17yEkpoVczOYD0K0Ulb/Mac2vQ//RCxL4yBY
IuBvvpisQkRVA07ViLA0pvch3sIY9U700MBjqAw/PTW6dsdqPGq5MCoszcwaisPQ
xmPv+ZARu0XNC5Yrr04QVeuLJZXxTbIIzsHqwI+wt7yxHU9dTBlyLcq75hzIpSE0
cfkP67P7IMbXPP0ARrbkZ2BCFNGm4HMakenEjnVgmLznYKUfxUIt8v5oCwzuX2td
2movvBMbqjR9etiWfHTG0nRMJeTe288uv6kow2tt3+AgjsZYCuldIDUaDHsLUVqs
hJPIGfJoCfSgLmW5w+RCCZn4554M3Ge0c0ewHjANkqCDGwFFQsDKNfbN2N73ez5M
PyT7WKPxdfwI5hLkir6Lvx38fYql4WTgMOe8cZOeAeWZLPH1NEld5OEPjJW/AKto
7hqotWXBL3fq3OCwRpGkAW36jRjvSrJEFgEQEjA9uPmsMospLuBSN5dKSjGI1FI6
fAhZy3D207eS97ya7y4s1tShqmJMvg4kfCJzAb19+BvymPeN3YOC+ZxSn18OrDw3
Q4NRxrBRJ9c41wjJsOXDoiU9lnC21VtcSX6V4RG/6F81DTVPT1o7oKyWeAa63/Ef
SOjzKIYeENCfeqTCpOapsoTLUC6kSI/2MgGlJme7q3HeNhKUtXsTofFI9Cqekb0u
ouivxp5IVPJkeJX690Gr7RBK03cm0ZH09wKUFyBxGRbHwRZtRpLJ96mJIbGJxpfa
5n/Fcohg9T6kZe0FE543WNhCf+HwkIFIc1RQZFfRawfne8YUHuLP+0/z/6zN7DuD
A5yG94B39iEnTJDXBpRQKbqlF04lgieIgKezxW3J44By+YUXR5jducB3C5ZHHOFv
u2BYwDa/4KAUVfT1C4YwE/K/L801u/mxDF3OWGazXm0TAS6l10z8u+maZw0wksW7
jX0K43xjiO4pV9uPey+ub7hHdzbvBqCMB8QhMdRJxkfuk+HP1CUnO6MT6vrdmiXP
xyUcZUuxMxEX21ehrGV9nyY0jA1ULYECc97Y53xRMIS6csdTdz5Uvquzy694eOev
4XA0DBkrY0MKTwQwb07ufBWglQB4Yz5AwuY6iWLJnrsHYN9RJCxsXI/DTlC1esGt
Q5DSfYUes1AFSrpCxNBQdM3Qlz2nlDgA2O1khCsjem0qs+TO6xz6+6bgL8FH93nW
rMb/mDqHtOEYPlTjRzlYdpKvuOImAImATJHPAvT/01juTsuGq/v6ryRyshn8ttA9
X4Cv8Vpf1b5GqV/7VNbt59Rhd2VjyZ/o3omFIdbMNn+H3olER2PLxFTDWda/LzvR
9wdJuuSr/Ya5c+1LrHUIeBgcJXvDKr+Hobyb6BjtAlkqZRUJcWI0XMe6dwmvav7/
9C7bP0F1H/Mvpu39WT2/t7Lzv3RM3rIgQLJHgzK7L1UMzXlcQWB8aYL6nc3FMQ7n
K71kuJvXZYjzXYq1JLt4V+7g9NTD9gf7l3MvLoHNOtpvJCYLeMaRH+T7xZPiwzDw
Wte28x9Ik1XQ6mpM0yncEpxHREJ07W2ShZepjZaN5wrW2dGG6MfZsPcsiudMpLKr
A0N1i6ZSsl18QtdWqROCB/jDj8a4XA+kJ44qBSRrNdULumq69+8HdmY4KyBeeAkv
ZatILg+mAx/Lr3L8EQSWNpcUdV0A+GzM+u4rxpn96wtpBl8AOwwJwbNiqr10aG8H
/bbw0lKyF9xrj0QqpfOxT/HjCswNHdCzTdc/I9S8vDdb/F2iSs+KrKY86PxHdHz0
l6d/egGBVXgrjWjsC4i2I1IC48uLK80MrF0l37RYLGFBEV1KfxZhFSRfgapiVmnm
cxpe0DhRZmOqvwwUavbyMm0QfVbFFcPCuVu8ksSAbCXOX8zUPeqGzGBCs7UqLqTo
oBUmH6WKoE3Hr1Ct/1XXEftuFaLx5UUgyMs2CcF829mUDTAKRePImwdUGSz5P86Z
1yWZOzfMamcxY485P9zW1dHfZr19FjBe4PUzgti4zfPL3/K+0b64TlS0/QwNV+ec
6HY4uIphQoybtu+yk24WvzXOIMHK3rSKVuFnXxiHOsBUzf2IC1fSyQh8sNTAEn06
tNhgk3hh7dm8FrQAUPTA/cLzdfUSXcDc5z4xgez4dFG1KvRQeauTbo75w9aZaDQ1
9YKKu2zbo/BBQnwYjfLwAMbcuAgcreSm5Iqm2vKJOwlJaIwO1Qqhz3G204PbaD+d
6B+s4MVYj6hiXveiOsSdyaXUBCNpWg7IaXMo5h2ZRBxWcdBiAjFkrz8/38OlYu1w
BHsDojU0tUsY2yQ+AojJjxonlqROEOVHCVwE/vW2V04DdZSac49LsUcZVAT7bspO
0CulDdgH7JVme8bNrUt7IPv4Sc+H+EVSFphWTMl4mIlDars+i47z1BQB/57ucyjm
ddejVeGwhGYt2qlPUO+VOG2+kMVf2Hw2PjQ/CpmAAnNUQjCgc6m4T138pUMxgwmw
3w32uqxLLpXEifrXsg/tW0dlNTk+5raBwJow5seN8nAJ435AOmkzkQePWONI18jS
4Tii/BVbiuPNGV2G1DSG04Vv0XOGP+8p/f02eN6oWINeD7WgY8KReEEy+v/B9Of5
B0C03XYkAuteORIXB32QtdgB8IMYsHU2jsfXMuDigxTGMl04+fBj06T/rlos0xMx
tS2LgVrh5cRZbh5lL/jJR5gOc/Gil++iRG6oIsBA+DvxAd0RwUaVRIBopZpkccmC
ZnhOrfuOT4TxbjRzeoU7ggZqHarrjFj9BAt+nvj4m7zoGJAkEvbxnRW7gSeaDqah
mxTOYUfzQEf0IbcylGWt7yf+n3qSLugM37Eqn0shl/qBz1UhI+DPRYLtLFPkmHyz
giQHX7Chw3W8M9xibVkkCchn9RbNYYjgJe8AXFYvVgmaPoXLjVrTXorvUOaS66fP
Vlp+gal4f216fgFdshoeO2HhuKVitDmhNIxTbrH8lVaOjAp1H4V+Vv9DwAejiYO3
khedMiYh0JuiAyumFiVLEs8wwbjNKSyJl1MZMYWG4J2BgZ4AOxGXEDnoN0Tpx5ty
PFNKV/ePlOdIz0C1WNb+P3dHMjOWXJkA0qRqMXX+L2GF9nO8J1YbMojC9Zo/xOTv
64OTLtZ7BTwIVMsbgH3wsXwYSR0sb7fivLXsHjeJ9wOg+Eueh8fJZuSD/BxX31Za
7Ci06au5W6mjeyf2vYLqPCy87oi4q1fwwlnhkKwnIrORq3lwshvGLIS2ubnPWx3/
uOTWSF3aRGS0AJkCU+UmVCRrcqGzylMJIVSuDvIy3G1rleffp9ctldYtQ2GE5N6V
sOrqZsENdjYNxV7Rg3CS0n61cYk0dCRpM5DPDIiuMx0InVhMsbfDjQ5bXy/arTRb
NtejZoiJIw8xqgdLZ6xR4P29VZItpehnlo5zYz66IsaALQLb+0MpTO6JuzGD+PwT
UMFQPjf0dJ3Y8l8DE0iE+CO2qfNsA1dQd+A/bHlqW0+NCF8TibEFx+xLr5+92ZKk
xm956eMOoCNU3GJoov/H8dRWdezRtEnkAY5uXoBPmpN+AGkP1rsGG+JC2DHQKwgz
VnqvdhgT3m5CW2YUILEwJvF5ZwuDFGCqtbX7dGZSlObQhKqKEnAyBEV0YAjN4kNL
J0W1ku7qjmpON6CaElAhQpQ1fAeu6vppWe+eD5NoPdywoX+CMGuqNfEEkC66NQ75
j/xm45DKUqp7trSyvsQeuGlzMDXn+4JhYkUFS8cAd+Da2aT9/dCMxTfxhrjDKV8D
xNuMbWJVeYvCkL8d14+GbxFW42jSC11uvcWODtkBU16T7aK3smY/Rt2eLNE1Kxzu
Gp3cl++JMMlipCveN2lYaNdFryUAI7iFodDW711YtBDggDiQq99EHZk2/fyUCJc5
SQASib8VosUo0LyYSElVxCW6wbzsenqCIsDseMcblYTXKc8Ti8DreESg0KlyR/XL
3ILW/1kYKPJJ0UZ4K1crTkRG+pGAoy4OH9zDHVgrpRjUduw4uEJv+OFVxr7uGcAE
uU3Mv6xoF4+sHW70yQSjjkf8D69nJspmkcap5E+EYunsJzPH6xv4VN60FZHJdFBF
SALHGRfPDo72j5rx2Hk/iRg1H9KK9oN0IqHcJ68uzfyBf5oJ3L15xI6mVID4vYbY
e8Pn1RMGgxJhli9+no8WMbUsLtpA6XkrPZ5ptE5RRNwJHWNRhhmFeS4HA7teW8n9
422+d8eFQWV7JwuPkiHqvhqyymtiTtBuKJtISvwuibpXo39/dzTP8ehCyVTtb4hH
ooiOsbgY9Ffla2anf0chLQA9dpKkS3XYltYmbdm5WsFBAGGnM9w35w3eVvKAMysf
tNLGBi2J24iiCPcHZAypX+bqI6kHixKQBvcz3rUqAVKy+ztSYWbp32PReyzO6MnR
LRKa9j7CNneGkEyxlh1bz2csCRNB/PVFGizi6qpIGtlZCRKgzNqT7MsLuVo5pWy2
W9ezvChVNyffCscWGSfdKp0fywEyvjwWOsTaVlaiGHI9MAGonvEGYILepn0iMlKc
ZGDf2o404UTcdVB4/wSQaH9kGZME5A/ue3oGNE/qW0t3W9+2lS6/eYhhS2jhkwaV
lkEL8t56nkd/39G2SnhV/8DgC1Kvc3VserUHLbiqUni+QZGCSFK5wktWEYCWRA13
C99bwnWHVfXTN1R8wRUMug0ZTQPieHYgb/acZqS1/k1JkgSGSvF6KKUeFulkZ6Pi
OvqJrkc49r+udL8Ynckjn5sLSOR4ttLZNiQDY2Z3amctmRiP8dZw1JuIYPEiYcbo
af7hA0Ts+kb0jDXOVtu3cvzfpRauFt2nHo/RC6rezH+HV4ojqR1doOzYe2yh7QZZ
ZjQUD8EVnp9WmH23G91JY1jtFvFu3FPpkP+js0jRi6WVLj75XMeBaKkpTa1b5kOH
9Gqei5UTJgNlcvzguYe38hR+kXnbwqFsOOL63y7upuX7or4Px77O5y0JCmj86EFW
01v0L6N7yKWIKzQkzGXg6HIWXQf1nSGn06R8wWangp4jIy7uzeww5WBlPGYRRJXd
eIWl1we8stDMTbL/7JVB8x7cief2Fq4id4njun+vlxCxB3EorDaalb0Zjb/ekrzO
u6N9DidK3pDrqA6fevD0iC77/c8bb6R33VF0TON+ymKS5u8IqA04b1Bc50q2C7db
ZOh9NyQeE2qwH/qawvqou6yNgglTxGcxYnD6hsyO5Zrqu4z76fpsSF6rmfV9SCvJ
2XNVMM2oAst9rN59ROovbPVQBCEQMP7LuALxTmkb5qD/zeCmGeaBdISFmYChBv3y
4aPpCeJ61Yk/vZFr05xbL7/CHC5tTWQHf21Q+VUijhWtMJ3wofN1sPH9HE5g9GH3
O89GuFcvhQH/yVt4fJTp84wLYAMYNOKwdBvqj+hmmKGUbyr03GFErw6vU8A0IE/6
j7vwOhTbEHbO1KtIuSA1Pf+1ODLsj6ax9p5XB0lNPdnBH7YVsxwtqaYAd2oEZXjz
AqI51+As/20CuQAlN379wt67HA3fBaxRVZHBhjMxBWa1tOEw7oaxELCAWK+tbluZ
i8e76dyouvxcdLto92k+IsrjVWP+mAVUcovUR2bpz77HXmmeQDpYfjuEDaxO4wah
YinlBwC9ewET1mkhfza7vQhY7S14nrknXCzYCCB/u03FvmL44bw0VrJkdFOVc4kf
8KPpMFx5j2UAnrcWTUI1WmKJhgTmJgWD23GhX0ud3xgftmdB3wnHn6vOM0bUNQHh
kwX2OYKVJkbQcxnllBPDqH/PhiV7VD/DL8gn59WpiAE5Uc3Ln4XVBbJAOyTdKZba
K0f8pdAaF+WL8LNM66udHgLwhSEWQk88fBHzaAfQplTuMfFFb0B0OXxeiDp6zKel
/orEpatggbus6J0lGrPVXW8pMhX6mix4c0627p8utY1d18A2rthfALhUJ7wPRm52
KI6cgs0Ij7kH33WFtf00R/HWs6x5GVPVJAV0Gn5LrpQXPJ/sekbsQwp0QPDMQrOi
caO2F3fvaRud2vJkZPEZm4+8zZdPaEg+aF8s8LzicWdDmgDIHwFEXHqAYY3ckowI
qudZhFfCJucnuoqFno4RTHTa0QFrntEYotzx3fJ05N9AK17lrotkY6GYK3MqXQ5H
/QWRzq66drri7QXlY3U/+bPkyw6t/NgnWFmy8WKpFn0rpmVbanU0U6a6Yiuwu6mz
NOEGmlmpMUbrGEVGy+H5SgHVAktkFp6rfcdAWe2njRPzw3pyt8k5QU3/zfQ6G9Og
uIoi2k8jmJWeaNqSWfSQm7oxUQGhYQgeCBE9RVhttgFFYpETghrV1JTFzXldhYoT
S3hUPHydKhHfJh5FA4KSfqqI/agwtGJPRuvgNDvYikB0FUr3HM0mekb7D2I1gi2O
Ry7MAdURrLglpePAnthg9p9WLAol5GJyqBpaoJYysbTUY2/gWeqjq1WGjHpEopp7
NavOfUgQ7mCLhBygxozUdi02tTc5VFXQZa1DvrN2vqY/TbXg7VahGkrvIHKkcKD0
0XKSlZGHD40qhZbZSN2RRHYJ8Spy8wcyTsLU2TWt+cFQC+tZ3lcKYOVKxN4YZI/r
aZ0A5ITpfUPqz/B+zxipuhGV5Y9iy2jt0IxbSGA7ByO0QRJG5pki20AlYwWhBG5A
IHP/umbOQw7OTcz8TKteG0O7GCKHX9+H3idLXWw7yNqqvNzGt3dq/3f7/OGyNK/f
B87HO8+BdL8ESoSPtWwAH1ZS38ipG3xURWnwIlfxYCXXb19fkGkcoq6LdXgob6VU
cikQiPTXu7Gq6fXDb8cksQ9p8Py2iPBXGDvR3mO/px+e7hDGPzM+k7RKkUI4hH8q
ZF1Fb2diW3gMgfMD2JeTFlVE2uya34HFeUgKuiiymoY5Peg3DnveW+OcvYQ5sOdD
veEDewfDgzI/1Qn5FszQeWvP6XExKTfqgJw63EMzBEOImkMSDzUS9HQUxzA/nyJN
aICdS+AMDWCDQmEapG75gX+UrLJHfYpmft+Fcih4dO3Cukcdncw+HOOjuqdh9MXk
4zPrrgTJwKL7TGFcx5H14x5pmlUOsBSiEGm18XLO+gG2AjM6bd1Ro6PWB0K7s7CA
Vssmy1UoDXlSO1u4xKW+v2U/aEn/PJmOPTPuQMlkTjG1XKRPSCF6yMxEryhu7ohA
x766Jwd9Us//23DOsYPrYiesDzpPanfEmDZnIQmhD6jesz7G1xyRpdC78YonvK6k
rAEpg1hVTPxZ12MO7K9n6bf+7Snh47N9IUB/9g0MF9/AgMGCPdf8riCnC94W6hhq
lDZhNbaEP5qc33WBFQ7ALNp7pVBvYii3waYRm36P08fPShhERcP/10ZYi3YhBGdG
brvBkW5x3XZWHNu+NXDKhXUHNURzgxKMvDBXqgQOg/w+WMMjPovSbC8FEiMeRTBP
wcYiPmtYGhCNxF31XetjX2sPllTUueNFfKjEj45181/MdSCvB63QzAIRr9AZLKpi
LUDemsn6D3VaxZC4SEBBHNTF+l4bCkf9ZakVVIu2mQdVfW+0K21FCYlJu2hld7Ps
VpGxxuBIVQRL9naO9l91HAT6i9U3pxK1L5dbIYY7UfnuD0Pp5NF1yJLJ7ABnYNKO
zAZIF3w3I6Ui5USMEGU2skWpUNh9UhIcEN+kTb/zzooTVLjUTsbJ8QFQY/omTEg2
c81Yo+dbaPceiLaXyAq2jUlUUnp8iBo9znuhDAlULMRct5AnWd3taEv2gXiH0Bbd
tvXiSZHuyUuDAYhJ6jBzCEg/l4Q9WfWdlZjJ+Ia+HwS1EejMxHPT/XQ6Ix+m4IwH
EGGLiF2rt+6Z7hErBegXlXK+/oGxWPPCgtCorD/sJorJq0GWNygeTbsAAMFrvDju
VTwBOU22jO54crs7g5bD9sWd2XkHcuFNBnlMNYTr8D2ih92FKED7ebNK70Ran+KT
69MNCoZQlF7QpmWD+0X4P53JaK4ZprL6lgeTPVWLxu718frlVc9qCgRPJxGq5r1F
NMZ8asB8KJPy16X+HaLaDfXwvK3YWYLP+9Ld8JHQJxQUWisH/2TLDCXFXvL6pUqj
8GWNqHUhf7WgkryUJpMFHO1gNGmZX66dS+9WxIrkBv0dNNCrvXpJcky32ildgu+c
zWBPktEnjRBJ36NxlAZA3R0ElRC6VjZtrPXWyYJ2VKDQZNyP+ME0Nfk3QHbdEZ8a
vpPsVTG9le3gnAzMBnVkYqImGGM3GLgno+yh/0TmiI6PPpOKmE8C8yrUyyn4zgH5
oy/nRrZeN4FNClGVvrezSIEmo1vbI9L9Dc3Ur6o/rGhGj8osRK0SBxquLcujrTET
elTTSRrP9Cfq7t1moxbMx1/VNYymPTl8uh32qQVlC0WCXsUrykZ6iByiXfXpNfgj
avJw1Z88Xrd0LJBtc0rg6PnXsQzAukQhX1uRcAGisS0yGEX0uQJpLPBkdvwrN248
02Kinc5GF6HvbvzLk3fW7P3QJ+zp/gHpI1VHbyPTKi+eHLPTH6HEDtPLhl+WJX9q
QzI1mQZohzQSO0ueJI2AoIy2kt+nB0rPgYDvwbwGwBdo8hfyDyZy7exv37OeajGx
gEEw8olh2glgSsyN55wzVQpxeJtJiH5TJbbL1Yf/ptumc7TR0L9TSu/AnLoPVB4k
ZUoruN7FI0K1CxA+1sb0NDHv4NBGspZBalakybvjlDVvBj3aJhagReKuPqKvlCBo
q2di99x1PBT+RlEgBs+EcwCTLBWAuW80zWNs0Fl9GdQ090jD+8KfkmgfYLAu+24l
xVzdPdknudLo0KhtfPYe4b8gkVp1yNA+1todZ/fSA2nCXQ99aBxOSxkueHNba/JW
pAzrwCF+MSHru9N2+Cn36U7j7iZUkcLMseW77K9d1reLrhgidAgznMx5ibakyf/w
aFdC3JzTYl7vVTiLCgKzmN72QWKijkXbYIDXDokCpWBl3J5GEgun8E5Mi5N30F5d
KqGUEtdOE+tHujIwwmR2FKDCK0ySf+sfkKGvHMTNbOhwHr3Rl0wJil3nW20RFQ+i
ZATWUVqIlTlOpFIFnxuQAA09aWs3QluUm9RTw4ptGU5UuPy09MxInhCq7MojyVws
d72UihiWsWbfzKYCltrgtLUk0f8eU4kZvqBBUEEJA+HMX8zF7L3E6sCgEkwrDOk3
jtda/zYAgwKjMB+ijYjc4Vhp4PLxPEPSYLslx1pfr9IKSPxDlcrHyxfk6QoD8Ptc
tVhCypok3XAfgBqk3ZJQkvuoXkfx3/PogwUHUcRwopYNzg2KriAjwZWVaWYpYof/
Y6OKYGAcVIDrcXL6/GbjlgygL9wxOQytyEYYuEP3wJAup6abICFrdtFt1QP/Z6X3
nLGz/cqJJOoMaZY1rSrYyaGHjibRLYn6QYgjnHUNj51c5mWnlHi7kcVpFCCKLuiy
oB+VYAl4U7AUr9IL8/qARyo+cAEbNbQmXvirtSfY8rSrfPgbDlbsiIQE7Pvw+8Az
LKfV5R4GhHqW1BbLUYT6VBZTQTFJZXegU9IGTXSdeW6IuZNQS+tbM3BiUoxjePFL
OWPoMzQV3bwg0okYdFxAFvmDplRfAhq32d3pmGHWWWQ2YlMFJCVyjtOt0epz6wpX
3cSrXDgxuoHtKMz3b5HzMAYMBUmQ/FHHRRBDPnJWomXcHhliDxPxiK1dCH0FSqei
32Xr4Egt4KleLC4Qfj5GNEyGrSlJgwi8rXmKw2y/2u0vPUK9JguU6T1W0ZpCXRV/
MO67/vgsGAU8zYUXin+NkJSY8Yy/seazJU+b7m4PfQkIcm2YyIXlaW8HJXrzp2D2
6ZalXQ2p0W1oS+6ElMnDAz3Pl2pCaqXMs5V1qm9H9BheSIb+Zg9bvDMCdfAaByj/
GcLK2bEIG/cQL9dqyIOW8a6rnq9Pn0448Jv0awYHxA1260FinrjOzBUjGFIcsy9K
FlF9uu9IXD45TH7d0Y8v/pbWAKdSUc8qtPmPn0r5dt6WQi5IGiABAXJiS9YkDjfS
8BjLtWsrsZAm5pU4MwaPsPyEsxeUTeSBd6mKfx2rxLUgiYwUQHcgw9KHHobJuVl9
1M3f0BjSiJC64dE6sEKn7vGLiIkluv8D9UIv5+XGpe3UpF3qHPtugUpoKS2A2W2x
pwT6+NyrrKbtAOOmVw9Qf8IHdsg3vyMFz3zip+FmNRcfdD+38dpWvfeLkoV19JI1
LUVKTKPCqdJWWBezQk8dh3Agw3Zw+tBF56Uh22aSbIW2h1jzomd/zpUOrcZmJAPz
YikFC2KFK47wiZnOe9CPpw3h9vJi7ZrcQfcyLiPVlpT5tl/5r3Qv6pck6+Ez4kI+
QY3aM5ik2mMrs9kQhZoeh6ZnYYTJs1UnygET+6sGgiq5eNdAgrDNWL4XG6otjOCq
RC13x+puZCt4dvBo2m3oDKoMg2Fv7KXFBwKaA7nbaik2Fu5O+1cQjF+DyYMFGcf3
I/ZbIpgIMJRfiG0YWaqlHZlGr7v9NKVp79Bx6nHiXM5HZTua+WPKMbjC3yUbZx96
GRiNF//PNJzyfipuVel5A/RtENgwseBWteYGB3UpMkW38bEVFIVzuRgAV/vyeFHO
CHNjuLZ1Kdw3IO5mupE13LVwrip/mAB/Nk9MIAqS+UpxV7VD6BkE8yFWtg3IvteC
gA50j/9jpXt9tltsLoHD1U0C/x1dsfsHAwBYP0yovb6oSC4nX/1UuUhwuitV5VRV
JFSevZ6epan7soXz9BtQsegV/fstOUlUPIHWUuRI3WjErX420NDStL5/dIUEbA6m
WJjirJ3UC99MSfeMPnWGEhtbOQAKxmROEUsJcSHiidVC8rDE/oibZO8YKNX7DO9u
NhINuuEAjQbe0dVqqN7lwXpgPf/gwJgSq5Hi3Csx/Cf+wKQnKdfqUGnjwl70j+Fr
kF2MZLImacSH+DTDek6z2XbQhQDMWXeS8nUA9xirFAdYzvyy3E1SH59vApNMT6He
KPHuJ7yRPWpi11U4w8EYt+wMsWtBnwGUtZis26jTr42ebufFfqvuoul3QPI+lydX
zuXuZkwsexG2+feKRiFaUQ/7qomupfy4kYK+nXBNUsuuAXK/vcZ0BS0Sai8FEZ6Z
dtp2+8r7XvvUzr+L0dh9ZrQYFigMlt60YUZSCG6jQR1o2eTuqa0OqUqOImzLFWOy
kyuuvX25TOJcgXEP71Pc/8HhuRcMsO3Zw76IgaA7WqmfmyXgM7f9OGuY43oIt5+w
7gKIOWQsToiMTW2VYtSWTCtAaXl5RHqLLWFJXaB70iPyXHtY2EodVTk5XOX/t64E
Rw402DFUBd3E27HFjtC+Ha2fM5VOVoYrO4TW/XGxciwVyYZU9Xkio3X+5lj3QdZn
1jbT+RN+eYGvBCReFek46TdNcHgyhw/eJLbKpWdaF75RswlV+OZkWHugYvoCMEJy
DSQTvu5JN8tAmsU8KKf2yKMsWCC/jN5c3esbylMpGfNT9pqQr8T5W1fUKwkRazSw
RM26dZzoHwrGbjaTfnOc9vB9ImK7PE3y9L2ZgBYhsmww0Z2ImvSA4DpOgoVuuQ2K
X7BJ82mGRgneVRKkQ+wPktU0LDCius5UB/vKzQzdeXe7tIr0b/MSlOQf2r8f/n3o
2H8Xo5idDgF0K3kv0d4qv11l0Aa2pwLYHY7ZLJij0eYHKUKassi5uKSpIPEK7jy2
LDJuknIbqda8Gr8usp+7A70IUylqToriRrDlctYFnWTs9VP+hNp7oBj5U9UV1jnq
/C8ZpXaLzxuaic8dclHCCZb4CBqk9iR/hzal/nB+2+mkl/BwtCV8NyFJnP/1GjKS
JYigCDrqOw7lwcMMVIvAfps40kOJpRvBhnnXkWnRlo6/NILtPILsrwojZXmVpL1Q
/JYO9OS3Y93eBg5eP76LO24QZsLqpQTebRbTceT12aa8Dpa1YqKThiOPkCAZZRWu
xHKyDtKIcVl4qCNc9fACHYmiQI4tV/YO4Dali44ka3SjnUV3/lis7AS6qNXZ5sgt
W8zJM2WkkiPlawSNjVeJ6KDAlsDYFR5NrJrzk8aKJeP5cb29/Z2yUTwGlyyhsBA7
NPe47qJz2TzSFnoGjodHvhtiecTVNWolsVdO04VgebBi9AelvkrHDd3LBr1XkIHc
RmXk4ItL8i2eHLsvfwP7wxGPaCRT4MahlMLQJiBM8037lb98wUpotYYn8a2QI0/f
iKQEywlH49x9P17+8Tmsv4BlPSABrmpz3w4d55bDO/C7WaZko69vnujb9JZUgKug
01ryps4GerP4+X8Ky3JEMbufHyxXjv65IZVjjecIOBD62pI6GAp8aPWiasMsDHzH
G2BFqdepOLKFAyrxeXcqvMawZgTLdWAx1cH+hDni/BTz8BRmP2bX/1i8i71dO6He
o7TAs+REbU7QYzhtyoldONoZNYSYKhtK65Q6QK7AQYMqCoMOU/+Phi45+naVdrui
UQ5I8cA3Ar+nfRJ7jnQ8RZ0XB5/4Qs+wJUa5iUNmXhsjDYwHT0r6VkCHmp3NhF47
Q9hp5u+zlozyeJ3Sw79YIbj82pzYkzu0DE3vGeWDcdWnRERZ3mX/u2PRGedstmrf
NwRt6vq9uEK9eFqNwSjX+/7BOBsWRL9wwK6IjnSug3c1dqDJ7kafRmYTGoMH3651
q3Q9/q49wESoOmMMurlVvbJIbXeGw/1ZRGImGYAz4z7J5YUQZyXsvXcG5VnotkcE
pEw4wKTYrH34EtYYK0c4IAexm59jaooSQ/+DhAKwMnkCGDCjdywaXKDDKZarDKOO
u7eVvwwVvJaZeeO8cDA+UHy1rr4NMvlj0WWGAEYxk97+F+QEFsm65uTzWCc58ru4
AYa49yjyIkPwb1sR6JQEqyTCSqrAqZOp9XQVoo18l54yAkFQj9IstDRYc5IkJr+/
9l7+IlqE/gQjH6hN+f8jy4KuPWA80GAcwqir3FLpZYupMO+9/5N1sHbVbRIwExEs
kqrvbISkEnKgVbO+MmPv+9pgA2JZZWW0wwEHrRbDkOl3snqL5n6SwwcLpTI9rgR3
S4eAuuG6fvJNP38BrgRPh0UljQjKiagko89q+sKWPEGdkV9qJA1Eoq5u0/feD8bb
Xl1ULNlvJR8qyGfWh9/vb58WvbFP742UgVOcwfM0Db/3kVuZAXBcawBPl19IEVRr
ka2vCA68cVqxdG2gTqhe3Jq5H1yff1FPFU7npOPunOz4xmK44Q6XhSDX1aC0drIl
Lb6bp+RT7PY1oatOw96QxkOSRkq1Xe1ZoZeBa5xJ1aa3zXVp0apoNrwfqYrVTA8N
BN99hwb9U3j/6+rBQAu6rPq+orrY6lrXlQFCg6CfanEPMXRDzWN8Td2HtvsOdn7M
QIhfSp6pkbldjXBXpJBgdozUVipcyiLww0Fza3t9So1JiEbMvwFpDzkAmckBUXRP
s1WZH4hHxXsANgPoTL1TdQtC1wBmsQQAZf7585DwxRSVbywxhC9+m0toswqYscdJ
cP5i4eOJLy++9Jrd0k4lEfyr13ovFdl5zaUwCoulKHhcKBHjAwgtJfPe0pXa1jw2
SURJhyuhUqz4GAbNawHaMpBaHM0+aa+tULgxjuqzSwwqNPMsxo4xywN4b8t6esi3
3Jhe0aFYlCfs6tLVBwggvW787wuXwvezX+XiMQc+hNwhSNxSZIlrmjn2pxnWciUc
hSf6U52UCUsi7+3x7JjO8EqZpVXfyGpOMBomJfsAP9pqKsYQcxtmyi6UmLMRpNsH
oZKg/m06BIGiRZsX3IrRkW3pJ+1dzSIgooO+lj6+A8Ii8QMP2/otqr7evMS6p4zi
7qmCWfKosha7cQCWIJJ2EYEoJlP499iDo5JFuZg20r4a9YaeF5swKC7guWBx1gp8
OBVE5siwy9bre+JI5yqlR+mjia4350Il7umbENJk/QmWh66qe2bXp3M0tikIh9nL
+w7JoEAU7rJsmKNZkrMHHdqYZjga2PLU1rk1MD4vY45N0RPnoxhKiQfBajZffaR3
j+upDelxpiOgYW7uBkBE2zOF5rWiTGTo44DNfa/c08iJI5/wXKmpDaWrFM6JTWop
BJJz8eMLIQcnyJOu1wjIWpbBUsg380yoD4fc+6mRxQeyot8PAkJ45Vsg0eg3zjVf
aDhycuaoZXmStd8Y81filVx3iO27QfwjEy8nuN7+p2XLIUqROtvKqbgPsAcFPU0Y
va8eIIPfqMaJo1gRycISy636y7BQCCQoXKaxFDCaydl4n549T0qbgw4IC2u2hCZA
WLmZDFg8+w1s8/Eu/Mk9ZoDxDCfcG7ECLdNXIdv/i58sNWUZ6uiD+5GS/ILtRorl
w93oCf2KmFpMIScWAQDQRmykj+T3dn3bQxz7sD7IaQPikELsBnc+RRYYi5QLn2dH
YThHoHqI/ix4w2IUWb6UBvGlyMC5FhQ8PufGPz5HAjfllLenc/dmqw2Tp3jIKtVa
tHSbkZhTp+xVKk1R01C7cwwR2JrONoQnK9IfiSOFgb9p9vIJkSHr5v5ugkn7I5cZ
4kz/C3p9d/tPhwyFZ3AHesEItiX9ABzBxj7HQ0LN1fFP3xL4Vtz4o4+9kM4NEYJK
Liwi51++/LfMjnCwxtWC5JgtA2G/HLXvhSiFMlVSGQtE8BZCQuSZaCtnlhBqMd9h
2F+JkdbiolfAaKfmz1o6TTqNks5W6ZfteIvNTgTN+ZXbC6BkCmvj6a6pebDLvqGv
nmOU55nwzZpBTdi4PL0ofIH/bUc9nC7mMyUdZGzTt4INa/w7BIKIFCC5Ff8jDGhN
x1UhICXeIn4exZzBeYeYyp69iQclC+KbCLL6Z1N7Uje5t9q2XOGX95WEeK8QKv67
4xKN0nPeTY2F0PyakngqIJ59d/whM9XvZBfZ8HzjnYpugFrmWLYgCGFfCl/DWM/T
e7gjozlZDqtIAKWqJLWVeZz5Fc5Ws6VIvKiGgUU86YcztmQLO2bp2gK+1edXTLUS
V4QDfiWvMP58cQXpY1LKVsfCJ2p43nXvYSZewjlQtTT7o9tVBfV687kDgJ+Ak/4C
NCUhfgPBAT6G6N8ssdVly1pxlHmT3YoA8oIDXwV9JdhsENPpGb2nHau8f1VnqTQ5
JE+IqE/JQDpq/KIYPdhzAnC3SLrCUIN9AzT/o8JRqhGXOKTO+/CtLFE/iXGeA6vs
8rdNYKB5EWUcjssgCgGs3OFViKEpGtZJ0MVWZ+pl0jgQHOq0sgGfpRQ3wtWo6//c
z5fowE65DsQThFLDd7fWOXhcSzQK1zOa/MQad3B6NC+CwDrG2+p7fEzTrPeTgI2I
y2xThwAcT4rsLhjGiq4bFuDhgNBDnsmZcxZ+VwUDATC3u+IR3sS54baGnYI0n1L+
nCa2e6/y7d05b34Yc36PxB5xkuowDEsobbrmKupJdBjwauQH9C6KCZEOq2/q6qO5
z2onrcoRI+PZZFL3wEZZVJ0SmuRJ0/Rf5sTDVTEEmoObKKMgDPtmzytx4dorjYt3
kDAse9/lEhH53h6IryroAu2V+oQFKc35gSy+XrIae/A5yTv1eJELreooNkybIcZH
XB/GOIYgUWiyJCX6L9DE+ITvsNCQe0ogOkSINqWgRtx87B062KOYtFjiJORfRI3x
h0RKw4WKH3mnUMu3yfb02yu+irD7N6UpenkVFtaKwvwuNCP3LsHdzMw1Rd2m9Va+
wz4d8R13RXS/47u2YRas9dmxCVMQIm7csV6FhDu83LtKdzqgqUo1F94NmpN84pp2
TFbZfbkm3+TjJNYypurgFOVEHalqwJamJtvIDa5o5nXYze2oyuUM8rSNRCKauJAW
UDvEUGMxPudqCyuaCdC5eQ/dNkcNKLm7vopOPCPm3HDV4FLJ77wG+bdZc8NjVTSs
7TBYDYXZXYluUpIP4R9ZH6nykLl0yE93aBV2ju+Cwf/4k5IJpYinl3kFUu7BtGA6
BwvGlo2iNL/vrPoGqx4hj8vfWYBfME6hZdmfYlglLG5e37LQKaIDRn6RUZTVfmq/
E7EvHyV8StYODl5sAx3uxdVJqAhAcsiTw0/DwczLlMvXO2DBSCFfmUxNdtMQ25s4
Eh0qCnZuAmqYcg7/GZYBgLBwObt9LbpUfpBX0VlXIhne6GymmPsXKNWZV2T5Tfe7
nDXSBk0HjhwC1uw0CkBQeOZmIgNv/fPkvXTLx2LlZHGCAkDhucOdasC5MFOzWUaG
zFyUj+0BEv5K1ldfIvjhbXY5/OsDJHRxjnXvzMzoV/N8kk4EY56JyyjqtSZEc7vq
FqJThkySIVuVSAK3BVSUB7r7EPv4PtYEZCRYOPQEjnmZxmkXU2V9KPjDhQDWyKPe
hNCcS9XgAk3RJlY7bdcgzb0Vl9JJZUfFLo8ATBotKt8aVyx87pDZJqy+PpmKO770
ixq+eJn3jhZipxhXOCAtwGNuUOAF0ixmYQKGcKmxjwzKnsYo270gTMhIXRBlKQvp
67ownEIlMkETimRhGz3YXoqUlL9OiUs2FJAlPmcop8ZJJt2PWCNHbIasrxWV91PK
Ob3gzuX+096Lb/5p3RsVimrpRGI3tscBipa1SZtghzmHdDyJTFhMrhVrukyRi+T1
v7Xs4w2XhpLqbddZeZRcwJzdeSMaq7drepmP9nD7EfyLg6f6TuRbRRpjlZCB1eXR
YmZ1JxEuAH9gNOwDF4cmTIZ99OpPwxvf/VovCpry75+du1wJDiTzrSyrf256utwO
9LSR+CG/QmJH6jaIQ9ucxPvXdieK0aql9N1ms7eDE0dqpWH35V2hhOyo6d1fUTjI
LZoycGQtGh/nfD+wISsCbQ3cN9zZhiZhO0rGTsfHb99k30672xFb8urpi7s3LZa9
5FZLOzdQzKT4QTgL5NCEDTvhSRsbczZupZ7UXL/SR4xR9ij2p9z0MZ3pse8j2KG8
Cfl0Z5vgenxE1HHdh+N1lihSCy2gV1/GhEpGWKWS0b4yCj+XrUBHkinR1vcRlBCB
wj6o+hijXlg6Hh1PugP9W6WN60jqppYbgfUPlX1qFoAlGBR5pZUCZ/8d4yEC6d86
lpCEv667wktHG1cJ+ow0HzM6tesK7cVUlm4rPVrDSEwK5v28r69kG3chw5SvZWnJ
eYRuKq3GxHO8fDQ7Kbd1PevMeITrI7w3TUl5oY2UEz1VYRfn/vfapS0ooiamKsfA
ErckAiOiFaT5MA2SZpa1tQZMpUfcZlX1DcPPxvG0LoDoPGgXXj1EE2uEej645sy4
0whph7JYQz92tXiRyldzHBhkuV7qY05FI8zj7dx5uHD6NE1QoLRKVa5IsHmFL9QY
4rqJqsPD1HKqJJyEv9X61/hnx947zjPc7OWHq/r7P5VgIykRIyL+L2GnwCIKa9XP
G7dSKl0FbBt7VYUdh78pPjIXpp+JwPwDVL2tDzDQLtDxXAJ1Cqdpj1TZW/TzrCrF
L7mxT+PKIB9bTR/dmDXPYbRKqn6+BDKuZlCA6NaFMeugLuRytN12qVNsJTXxYE1I
T5YtYH+zqGIxWc+6R/0XX0L4PwuXH64lwlc9xGQJ7MiB1bu37nms4w9z8cU/q12o
E7gQIiJ1jKDTuPSHD185Q5/T9IL9kLi2MOVEWJG7nOKt4Tf2oJPV1JJUCry3OntD
gv1KAdvv8WPjUzQrbA4LU0I5mJ3PyOTNx4qdMTx7Yni+P5SWMRuvFwgQ7LYqIP8B
gtj0zZcAzJ47uYwanad4SXlDMrRKhAU1/t5nrsionQwHdFUjZ9ZANMaiDTo1d/61
YuFYKu6i914yNwrTJpSSBRQd/Olt8IodrHDN+TljdwINrD0DKG6WKry51WgIwyba
sXB99+QAsDbBoff1PM+kv7UiS7lRva5trYph2DTJNK9sEhxKzf7o0GeYXF/FAZkG
q8NE0566KTLlz1Iqmp5/y5QbM83y2htmvxkZciOLVTVdmv6b0WJvjMh8V/Sh9pNG
94+/E37nXLFYk/ypsG+KKjQSU/QWYGUPrOAUOJBj9uSZBeOZtvWxRXHLdrWlJA7g
X50SROdZy1iwolhkUUPDCPFae6pOFz70hWdu0O161s/SPhO/YNbcFNEF0ec+jqZj
42waTnNvRkPenYgWnBJpOGcjI/qnRxEtOuwZxhN7D11S82ia6GXa+g3OMdCuvH1B
8UUkSxMryq/zTl1tcyFdNhgR163/46aniSXnnZsg8REaLCSDY1DAp8Z09/NyyW4m
wgkO3wTfOYSrzgnhGUX10F2sIeUSrII9Aj3ewLAf+cCgPmTZQHLeGsBzuhwJhhLK
H+zYyTwFKTJy4lkQ9+kq30aX272rLZDgIvNen/fBEg8F8eGxA1yd6NfaiRQB30NW
J+qrORz8Y2ASpErBTG0ZaPvPC5yFbULPO9N2Y21pwS7d85Z2WUiS0RwZwIq02/BB
ySMlyNLPVNaWgf7bo+QGzcuV/fUYePgP/JxMzpaCx8i/IkdQA2puz+FTv66AlKCk
hgquuZCKPH4V21B2HdgJBzZNOs0Y2mggCzfiN4jThYWCNGiChsREicvpqZottdbQ
cAbj0/pqmZ8HFJUyVIIy1Q9NnWx3nZeGpNF/r7aidg3rCu3dqXyKEO26eLWa36Bh
Hq3ItZBDOf50fZSG9ThxxM2wH5nL2Oc4yz+Z1d6HFpC+lOqiaLPTxpy7Ef/1TE9y
AtLeFInXDlVsq19Ud57DyfW4IfRV2f8LmsjIP1T/6p7TBtxUMV0zxhVuzAOGqsOe
Q0st3yLuhcwsoNzvGl2AzNPTK0OjEE4QRkIm0HkUxqmRT7Uq7lWL8kcW+dYaWNlO
glhin+rI54PhPPhYx//sf+lBwhvD35cDkyI1CFa8j30wURfIPgFNyFSRs3x+vG+y
yPsE4BL9meVJttxZh0qnB3lJ8VlSrVwdug0MOFmRPGvu7v4O/VQOrCh+FKAMTlDD
YY426O/54/Rj4Zqbczib4IN9x3WFrn+j65pWkmJN++3ct8Qs9alGHWutbwOAGic8
5eQiZBVKqiwOcSHD7kLr4ocyXpUhpm9hOeQIryaWFKQAsyp598SYvjVi5Hwlytg/
12rdYdvPbP7VjlVsYXTJBbyX9U5UpWxd/f0mGu8jnGgsrxem3KGzkcNEOlIMDvTj
cH2ae1+pIoOhc9MBaQbT5iMwD/n4fThcBB/qjzwiAug6V2q9aK8priA5m3e3PUq1
mXonFH0AY5V9jPtZbqjGAxOWoAnz9J0YGlLO2NYSSIgoKe0L3OUXrDMs9MykItTS
QN9aJtVrGCILQ/R7NqF0DPkYVQ5VwpEro3OT+XGJlhj5yn7XuBClJiGVCEkd7npG
JBTCagkVod1mHM/Y+NPrG6QNTmJ/gawjwd7ry1moGD9IOBz+ivqHmuuG/lvA5RcZ
yUt1z16VEiS5CN8VwUlGCoX0CeMPNdUtJmM1S0gNto1HAerzBdDTKsXsthiyNMKc
XTcU7PLVB0F+ZWPkEkkixRXEI2wVX8YBDN2t6XA5QzpGSQ7SnfvBg8d2JyBBgwhB
pTDeJTAN0zcKS+Jv1NILOmybSZVdIbGxYmIg1/IAXAjMm/V/VW2vEYml42Be4d9e
WE6nNItODiEpyARoVyDsAmtm1V0kcn9ZkiFZZDN0kR7M3jUZh/JHK6uCv0vl16pW
JsyuAAqQRBjepgvhckHIBylJEIGLRk1sakmq2s+4gf1/hYDHaYs/E4vBAtuByg90
bdg1aJnxKxQDbr3rj4Z7v9/MNSj07OM/1smafxiFNz1QBos0NB0eYa7hTNW+b+U8
EqF5AUvk+7wZWvEUlW7bqM+Z4sCHuKLITOjD7KWEypYzCeMuep6RIiA9SetwOnN0
3Ts8iFGb2ZfaS2uofHvuNWOXYiG3Phqbj9ZjwVpdcP90A2YtrwxQbcsiNfYxBB9v
kv+m3daaN31OFSROaj84l0O2BBRrY3glqTVxmruJJrZ63Gbrwx0sPtj9nNRq5Z9r
fcSCyZpXH8bockdgVGPYBa9FLGbR+37pLOYaDj6Q//EU9QgVxvO84IaWXTsSYOQu
FO5xoMx4P93wLAb8JgfP8PYbRAQqlBVFoV0vMjeTF95Yzn/5bVNt1VPzhhUct9Wl
FS4aaj6+CDagAOPD5CQaRBF0bjIWDxA2urmw9zdtQTx9d6ZeJZhhwy1igITFnp3B
cNagfR5T1R16voR2GqXxUg6sw8zVtgt2B3tSmhxtsGlTr/M/zqKye0QJG+VwPoVQ
m8f1qpIZ0+QmjyFSJ8oV+du6gttcfmYBLkHrSIDWZKToEHC/UeQ9eZ6LM4U1oe54
dolweI6mYvPCfmtvtKLWanYd09UTuqq1mPz+spj2ieu45nDWoaDCZlbR/V32nAZ1
gxy4BEUE2g1Bu7m2IZMJwVvm0hNJfDpiSxjjZVYUBCh/e0GHEw9nzxUN0Xcn85zb
HJ3vfxP+QHeQ10jbMs0i2JZknh+SDVyIxshl1W++9ED6Jc9JgOvSeevaHXgVxOZH
72bn18PnntbPdfCT1CkBy2ew5HZyjD87yCdXCO9eaoYWCnfLDmMp7GB0X5PFztYT
wNbTMtGFteWLWl5dEtp+3mAROZcCkEEIKEt3Q4Y5U3ArKYhqweY0SuaQSwr364YB
x1dDnf5yvKgIq5cAWTLrQgcD4aysszubU4y00DsbbB24SIgv1N4AF8f9yW8TkyVE
Tg1cA/Kz+vREWxU49RqbWvcW4JJbbhmZdPd0ho2tH3RRJaScYLGn/RYDrdWtB6PY
34bcusUaedHf6L7Xzk65S9JdQRt6SqFNyE1N3Sseo3rGbAmI6SexmQgAlLKH016X
QjM4Mk/cIlwDmprTwtMnI9AIs7zfjgwY/w5X9+LgveMeSFJ0VQEXsxkiBfu2PymV
m2sntzrib/cqyg3jv+l96TSgP0bUXDShVGziCXzRXS1CHw+vm/T/W3QQlftpa14C
IPJZxvQ5ee5nb43h3FMUVuJrxZD7KGNMWgBD7GtJlllZELrVhzpDl0106OpcKFCa
96z0GtjW3+zci87qbAUvpOL6Ze/oqBJfO2U1kxbjzDWfg+TEA5zBpE283BGflI+Q
cnNn8O7ErU8L/TCsmIoHYuSF+OwS1txPokKJeqKZHwFJLgF8yja1ymXY0U8sy8PD
RQr6KflnO+Mmde4lDjVLHuz1TEZXRJjCaB9RuRpglK+8INxVS7vsEkmIS11Ngf/k
dX7+lYVb/9op2wfwrIzkghBcMszjt2nMjcd6SirBXZXPYnXr7cboIW1h6vQAEQvw
OrH/vvZa7XPpX413kNZRwCdO685gH16FpHFIT/hLWziObuXT0cj9o+e95Wmob1H2
lnQ1dF0mqr2syPl/t2jDNCDhpbyFR23mYZ0WW3ADDx+PeRJWb2JQ1bOlXWnB/sV+
/pvZukVVuSS5DyO9kSkzaTB1vh9IDrSu+TvjoFXoN1nwqOtlmwq6ATyfGw2wVyet
JCbdupf4u7Wxrj6IBJvdPL1kcH1D7w/WnXD2MUMvMc2RpTo497wV1cq/91dCxL4i
cUDY3jiospMVBrDivwEBmEPsSjg4Avt+xoVXaT5yo+x4lJx+pnQNLOSxmFfkiX2U
O+VTK47FkEIIJMQIFCKM7wWlIElIJNnVwTKGRzQftNLy5a8sv79pKdLUGzRZPWmP
NZUQZLAm052BILtxqNW9G2hAUlVGfAt6docxEM1gIEcsVVFkVxTM3XPYk+MeCaET
ncF2hDl8YTAZ6Pl4TOM7UryPQfftp4YADUtJAOsQ5hR9jzNdpkcMH8BlY+HFDYAQ
YC0pHQ0rPf5BBlr7Qh0y05dwFi4jdn0Fhf2A8ni6I8xUGZl4QUE5KyBiGkDR84GN
LoII5zLQvehWf+XSG1NOD7z/SbwS67jVRPVJEiMIS0jtDz4zki4WCymxIqJcHs8Z
wioyaDz1IRloB0LlSqYgqpQLyDUJ4FMbR3POqfyNODUKSPG9uBG+MvDxOw+q5pR+
Q6ejwXHSAOLwQyJ2DG9AnHmJPEBbrqxb10Qf1yjcmjkOGpRPpv6HEx0sXuWVphme
6ED3zhVCSYNYeYqk7+5S/PUQrIO3AoS4WX/01CFZi2ZFefnuRBLJFBm8wufhbivM
nNCLM0u9eQmKFTmgvzsAi2/apyjCI+fGoqJaT81vKwtwS+LVBeNvdey91bGa2CoS
ASaIxCB38qsyYvcfn3x4i3DxB6eJI7cuo7D1W6NUBY1YDGE4GLVznriQnRgf0okA
G2OS7mwLOTGEiPYe7RiVovy/PI413mEyBjVbMz2UsQm8p/BRghcTR4vEPmDJljkf
AukOjuTSSxJTLgT9X1XzQBBTcunKKVRugmBDWQhD7ofslVI/MSq+WdwTaltbJfnd
VqPVZtm9xN5gZFcrnNWxaJvrLGs3q/ao0K8GkCvylnjZJdGSdpMdqjc8n0jSVzrk
OW3wmNdH0StULSD6CIKjmYLN6BNZ3eUZ+3gptkpPIxRfQK6alU0hX1wzUFdsbukc
+MsbVt0C8JBtw1v9TahGl0v3CjmFo0bMieskmKJVhv75bQZZK7BbpoH7XmxfS1NI
PJDja4/J7sSqEWhWIFcKFBYBLeAC/P1TY+ntznVlCi19fmRxFiBkQ5MDUtKv8/0A
s0gRhUBpLCqLTfqUYN07xXjuVaqTf4XGiQl8O8WdWH3QuDqY6pal9FP7mNOo2zrr
GRRWUjbfn20YMKSasehrVMv+CD7bv3IcvqJcOqWE5q2TG10kdHh0i0uTB/t3TKIn
nA1HRGPGZs1IczzAPmBG+XegXF/YyzydYvJV36yQuQEOo6NGE56d0t6FiDlhE3nf
4ssSOc2UDjOzIs9kUoVG9I2hGf9CVv+xEbqS0hVp9R+HLcVuBcsONz43EVJHni7H
FelKWuviiMQbkYhNjjbBCUzn/wFU+1ZznIjxE+HctR8f2bAbxkbDveueqnuZ24+M
BuUuoYlVqN8GwkNhfL78ksBZ8ihVUqsgQQEUDDF1z3R4faksAL/7s28nssswQRtG
UFKQ6AT4s1BuPphAFIM+u/RVKY4PRAbvzwv54ClzmsXaJsLIGBkmhzLYCQ6sBSzk
I47U8JKIrewec03eIXlINtwyThpAR0S1LSuqZU9W6jcEoZ4GwYCrapAKRBj0xXQy
zW4rPuz69wWLzSRJrxhZjF2V9pLPdDOyD3kBmUp8bNsZXh/GsAMnquHPjYQ7oqLc
9wc43pR1apHwdycIKKOfNewzYJD8HjwS8cRwFRQk+osJvEp03C9UIzl2B15FSTiJ
hWHOS6a1+kd2b00vygLltTmtMutoyl40+4x3TfNOdidmMm8l1AETLN/nK8HH0p3/
sSA8HGIdMESHcb+wKF7uLPpzPurk7HOgMp5qx+zopZjHWCyfv3qN6aIOaxUAs6d3
73z89je5tjjV47qZ7VQh9i4ZlRo9vpAyPVKQa7+G37MXnZuOPtE6BNpwRsxOjPZU
up9tT7xbQB+3Bu5rhDryHN5FrcDcIse1i+rWSdZY2F85BHVWBTj1Bvi4ZHGaOHxn
eB5op8lLvznzDFzNv9PVCle4RdF9XuSYGafryyL+qoRVD3Iqy62LXw/t0WFLjLoE
s7/RhnfrqeT+PzI3M3GcUr9XMEyF65jFYiddNmoWY3l9kCQROSMRrU9aGWTQJVcy
tltEJXfIfwIHFkBxAbRsV3pxrlWYVIaUZGOQTqD5ekNpodcG+HdKxebnGOotBMss
OAnI2440iIJNKGIL9H8QFzzbO5hXKALN23+lNWTqB5aikXxuHIqKtYMA4thN64KL
DTgrP5O1wyEtZEXCZb2DBl+sspwkOh4xAMvJbkSwyl7AjPCPZtBduTalWa/wvl7B
zuStermWXQfXIMAVxp/1TSwRfFRM2Gv92TFsSHug3dZbCwy3jKyBjGnfqaVNf18W
Zu91hoiY58vk3cvT8AQmPmDGtpeCbo7LiI1enQnR+XQXVwdGpJ4iKZQuN2YByr4a
60Gs8hEVQwNPABt1Uluzn1mktwRao4UV5y6p+gmkIhqgakYoLEbrWejKyHMqKf2r
AQemS6lyml82IuxDYgh+YdIpWcQoIsJK3kZboEk6EOzSJyy9SwnAqvHRkLxHDzcF
AXAyKnyFbA6Lff8x9ppPaposNLHBJCd6Hz9LRjhsuqisjo7QBQYp0R/jvxuye/6M
5m/zaSpWihcaK5leu1ljKLLppSe1MDZ0neLLlxInek2CYfdfaS/IPu+qSGLLf9Hk
tITaAf9qPuQj06fBXENpQH/8f5DjtHIdIIwrUY+rd3y0nNlTvERjEfyKfGmsFBth
YkWB4pt3x9fbBdYjUUZa5uO9sXxYgLQU1dMHPXHeHSc4z+VXi2rCfFrOoSN+WQdm
whxVRay/7T+kToAM976WHTySofYhxDR0sg03tCnR1rcV22/0UK2DaiEIAwlJOjWj
ZjQp+ryrv/6NJCs2K6yC856D/NAQEz/b9tBQSlpN5Z6DR1ZShlq15FH8OPzNuiDI
22Tdrj3D9ce4VShsPamri1pAhvRT1pLjtAMksgO2Id5BY6MkX8O7SDIU8UXMT3mR
kDYlz5BYnqQhag6rL4onzbIhcf07/JiJZkhBayUpNLfpLxMyHB3jDFeumaOx1CIM
ndb/NmFMfPhF/NxPSrXANH2CAWkAtTOXRZZltK6aua0YrSRBQlEky5LxwNMw1swa
xCfFLf0ui2aTYwGjvkUJMVWtKMDmlsTA2/0sXQFrsBUGFva9yELYsrXkQabHGDq/
FekNQVAgjrkyuvFa2mwxGk2fCcq1GB4rDAedbOayTouESzXIttgf6VY5oCoXwbGD
sQyL7duKAUWoJfD0RRVIrtNRLUXXo7LSWyBwPXVHU6M0cBxFydh7F+Sc0xdFK0zd
go+dF6b291CKqQjkpHK9f9Rq8l13sGBQJgS4vzqktFvQt8zXGXKuzJayZBg9GGDL
yiPg2V6i+6vd8NTCBW4rOcCrD+ZfeOFi6J49W7jDajpPPTNQEghO6kQ+VSVt40Rw
monwXcKiN+TF1+0Y/Gi/XslO8osIatQ1mnEAM6109nF9P1jn5615T6SF6/ekhObb
EJxW6bay8BSUIo28DoTMO45GoUf03TVURmQri9In5sFoIXRuxTHKjjXJAiMFUaZ6
4z4bOWpAfjrnXhLlppZzE9KrYDZeQtkzhKgT1T59wfBeoAvagu0LfkmggcXwPus5
CYKAGuaj/7C3MP0DTqrK25vWAOsXjAuSSCCGntf2WX6XrHCukgwL1XhYzYKM9jXO
wrdWYXAK9NjNRnNZbdF/E7A0y5gW4EQ8Cs3KZhiaNwJlpvSlIrlmDcSe/qOVteXi
+Th0Nv1lE29fTVYB5QO1vwQdbrEpNPbHU+bugLyeYcF+VQQ6F1UQfFU5qGWOd9cI
KtSGM+yiRCy/b7n5OD8dFvf9VpBcvA5AjgrvvrcllDvyRSwaJX+WzCArm9do7gsc
EJInJ+PmJMGQ3AONkTpXs9iE84klkFeIPYIW2VeBxrjWDZqlS0H86a1Zfeg6fpb6
2lI9hWcMEZqR+J5LuYBfNFIyjREbEEyXN2/MtfZTmPhsYTfcWErpeQ2FnGH2wMAG
2Z0nzW3HzbqG7z20EbNbHfGD8TpmUJT+e0l4kpNiP0jKYklASeS80VyT6viLKhNc
gNe8rSMw1WXAtOQOjB5CFs7PORfYCVuSC3whzka1imhk9vKP3XOZSpW2uagFVU0E
FG4HXlutFGI1Gp63sJ/ICH94zoSBA0G2YWeRzriAOCFClQTO1JgiTzX9vK2Og8wW
5wL9oPWhAnKMjvlL2E/nFlHuMf1fbGc+q+1xGATMIx54q2gxB1XA4Z2SSsHU2ynz
g/5Vcio8qygjHjddGipiIZo3nJV3Eal0uy+pKEPyxyixf5BTclqsDpPyJyfy6JSX
n9rIgzjDJX8yZ9/Gb8vB9WNgILzUfmJGqmk86pcEuMBFt+vXuJZvFH+BgMbasqDw
fBSkUmqOyUy5zRdARVpZWMmwFAx9sNP1wUAVbTEeIzJSS6KaJt2r1CzAGZP8MfgN
ib8mlJjQt7ZXsGpA6TGxYZiLss32VVskAh65SnsVJL6w/0BrRT24soy6Iay/TPoq
phVmy7F6OhBOkRgLPsI190XQ3E2BNZw+pVcC1rIT5oHniNk69cgzGA1hSKCFOdLZ
rZ9cMJfjCwx2BSy7EjJu6bg0wiPgdAZNyY5kmEfVv+Q7nCBfhYL9+AKpI7asRvUC
qGTPiScjP/gj/n2ZX/LGbtQQrDHwrQmjtZyLK85rSLTyy5HmdrpPZEPUTSinsMF3
PRSTk1mA0zA0U3MG49Gj21Pm5+HOvwihMKMzAVRh38hndee6XTRpzG/1wg4YpqTq
b5Z9d8uEoLGYnap0ubX/VW37GlYz4aVUPnfa6JvJFESJmZ0qa0h1Hlvy02SvE4eY
J/wHc+4YApWhK5hzMXap5/RHSYA5G5N3JNBircGSFYhqT4JXYadAxykIFaftBayv
X06jxX5mIXxMa42eMvXUOFnMaFwwC7FMSDM1vcoWm4e27DWwqBljpbTRlDQBN9oZ
e0ENvfsPZFl3zRiidOMXZuYu85gkGDHqTsQZd+axmBUV4ieiDlya3smhsXiZX588
bNdNlOoUfgM8ZWyZUdAqKiZkQWCWuCjOkkeg+qaZbw2r9tJpfnVHSlNvEZZNT54M
I60dyaSwgacw/I/+FxtIhL8GHSgZuXCzDZEQEW58m8q7iX5UF2pC17leIzZvvuwb
cTc/UDZJ756JDeDDsQOXNqgEcTRc+/eg1xx1rXcyhIbEjSucgVDoKMo1u7Y2Ghre
fJ0cAWHaKhaOWn07bbMOzkaMalyH5zqPOy7jVZotTvpKCj1cF/d9i+UzJUW0dqnM
N+nVvthhQ3RBRqVUlhFe6uR5pB7drYMgWFKRkBJ9x+02mQW6Yz9w1carpiH9DOa2
gDqkuLK0O2OvjmDzfxkmmhBUP/1yV8cN68GhiB2N/mnx1anFtZuL0KvYb3aZCU5w
kZTyR1w1NHGDfedURe+xdPM+t70kuCb0A02yCV2zswtwWlsyjeFX8gSz/RbMV/RJ
SVrMP+ax2j/ZE9LKHPPMRAIQ32ht462HHEj6cjLc0vlt17/7BYJ4ajdVhkarRT7k
vSSSm2DhfE0YcLHD+z4nOFHSKSorUCq/wPbkPsmoEIlFbusHH5E5IaatEWheMki1
0X03NLamus1VfAJhXnU4nujOH9ILMQS63HnjB5vYQP1w9saGIrTuiuQ2RsuPRPNu
S7lZ+UXVSZqZ0uI+8JC/nzi2yNZpppehtFuFTMqrth/58gD+fXji01Cqa4c+gwz1
Xkz/k3uWjmVWFq3B+2DulgsaixVPxh8nZVaOKpx8XErmDqfapyZOKuTxhwbJzu3I
vCFHB+i0ZwBGkew2HeR80B991gc87OMN1gFoZ8DEZMN31aWkCugejMb1leo+eyuS
uq0yrgp4srjhJQru86cGE8Zp0PBTGqXqzRDymtoyri9Xj8woB+mgO5kTEydy040e
AZJ85BUbU8+CfTe0zFrOZw5HsGTzxHNKJ1HrBtRxzcZwW0GfKnDE7+Uaz3T4Vp03
Kk8OmBe7r2Th9V7aRUCDj+uPcgfohrtytFQM/luev2P7RWaxSoH+iWZm91euzMwF
7lzEEzDbnXS5Inj/TrZJjcM1qR7AZ+qHrhvBb8iSTWhGWCDQ+o7HXMDCVdE4Lu9T
SNV8zLly/MebN/40TgMqx97Yy3VYcZvMTgYLM6vswieuKWXXvH1BeTnqcKL/63gj
ggHJBo0Q8zsoF9DDBPof5CkMdJwmGylHL8ZbGA1ujBekJt/UoKGgoMN9eHuwlgAn
pFFbF0tIEEtnlMsOlT0IxYfIUv9CqhzTLHQ6lvDS9A4alYQMnrXooJw59+h5onVq
r3L72n3rqaMrP0sO9Ukq2kqmS4J+AIulDLjwjke6w235JNZPgAQS+/iBoDtEmGx1
KjXfOuOkD/lZxcRz6a6r13Gadypxa3ingB8jLFdNoCyY78+xKbvSHq5GMYKVnAKj
rVv8dVlfHptImhuCyPcwo7XCn4t5sZrTDgbM/Tb5unQ7bCzrVUXco5lCX03Bqatd
wN4gAPJG91uZYSOa3PeeWK9fQpeUtvt6hMt/ZsuO7kWaWv7SOGugkdpbTfvEMExv
j3/hYaLff62F63oF8k8i4HB3Bc3xxyT48EwqfZnwRHEQbiqN8lNDx6haPFSyj925
AAX3QJDJ3WaQMsY4G6snejAUuCVujRLcjwZpXdP8T/bUCQUCPZh76dTGxe3qZxNU
k1z/xJCc7OeBUHtmJjqVffkPiaLV8DX+SNNwlBi0uec8oY460VG2iAw3DPYWKh9X
R9Wu+pRFFrsohYwEGkWyPhY5RWjppoqAxSXree04+SMOqd967Bh98jv9Z3a1joWh
vv6jia999FZd94t9FP22AdZA2bHN+JjO73UhAQJ7XWXfZWZVNXKhI1eYnNd6g0RX
eWuMHDpQ4J6rWlGbSFOW76DfqDWmqoiCT8rndALEdFaCXdhD+CAO/hInf+WsArWY
2ZJgchTDdQ8z3eqU7K0xD9oJMBvgScuy5FRqpsULH/8nLQc/R7rJ7vIMGD9CkUzq
OD+xZv3X9HlpuVlfCyYb24ftFzPT9HQgrz/VTQtyUThNYc128fRQym4jky/EoeEW
w42smY3hj428f2pCSbpNEwJMH/jgBzgYNWikDJe4QyaU62CXDbUOhlD4+ZxOK9zD
k5zNPR/J89k4uo9EmzoxdCIZzIT7BWWzEqMU/PdvmP5czB1ipU83pltAet4ji4u/
JafwjuzH+3FjXnFkvu8LP/MZHPmr7XOIIIll3yUT419uyr9kvVqxSR/4X5PFfYVL
7TKDNbTxbXj9eiPLMHmwaftCR0yO6SYRYQBlcX3RZ0GxBVjt9NGxqgCRio66OqQ+
hEcbp106371aPI98d15y+wc1ueWg3/fQWhrlTo+1QeX8+8CxImX0h/6bJ4e2Nsw9
NBdEmBmmqAHWz95IbhFvOrS4Zj75mMMeojp3sMkkxZ2arN6qyQaOmBYNXVVWczpm
7mVM9UWIMntBTSMOMlNu818YeTTPZluD0D+iRhG7Pfuy55+NpcX7wddYpSS89KA+
3+D74YDzAnBhlzSmyQ0eCoTHWHGfgt4YRapw44M1WLfesZ+TgwQZKaUlCPGuisba
x8V4SKSnvRP3vKz1Rxuv1H9Z4togKV2hcjQlYzC44m1GdTvNEvYmB3aJscCjFotD
ztd9CekPHQnRbutxx6LPqQ6Xznbuo0ouLkEf3gFPsoVu2VuQurIhnopKY51XceTI
nJp/iLfkZivQFTPLq7+pX827+ZG2nILEpbkBdo5TC/pQ2Ehze2/GzHx41fjXp490
+QjDL9XLT9IaUVHX2PsjV01EPUEMz3AqB9dXaSNwVEQvY+340qHOOaO45z0XeoaF
gRggqbUm28Zw/zqbOQg4tTO4FFgP0wpw24aIRPZpj0lOlqjuHJdMg/oDYiO1ttUK
OmtgvhFiQMcMULoWdp/igrqNQH0w9RW3nCWLA0oDpQfdTCYSKl0SVt3AFWkUgVSj
bMueD2XWGFEEebFYjDSluM0e+lCU4m7fBA7W5CWkEw82dpYNsw6P3ksd38fLO145
O2z/1LcTbb4dHb2Gw1SZnvXJyRNruiCnYZV0Op+WDR4yugk8eSkez1TPzn+iJpU7
WTs9fGllSXqdzNDQvtt8Gt+5Zk6YTzDa9iatAcUaxj7zh9I44fFDY8PAgtYfIllv
Ld7u2BU9JRvfSCLEeCxQUREDCYV84pRwK6UQnqzyAIHcccdCCeVgeU1/Agoalv9n
khIMGS6Xk9ySY+vJyJqsu5KsTVlrUCNw6q22CSXDqWfuJSlgxmfwyNBoRnN8nA4v
xeHLy58iJXRiSqFWzOqwWyOQ2hQQrw410OZYhChTJk5B9myoVA78Gn3JHtgvV3ge
ytAJtW+nDkld5ZmSJPwuME7jsJ3EmNAOON+kpHcV12QIlguAkvuLCp681yS38tpN
d5fMIQJ9iAUaGXbo2kAFF+f0RVe0II89nw8u41q1thCNGxKymP9LzGgmbtQgXUS1
s5G4nfpY+eY46mHNZeGrOBu0zGA2Kt8lzmVgUMItqwVe4S9K8oGbnDZ3gHxKS9JR
aaUZJXh15bhjMpbbEhMsx9dd6MuKePcdLCyzTBq5Nntj3U/i5hz8mktFlXV/hDkN
buNd4XJNO/fHrRUvZjjnc1D2xzxKgsut0AwwMNHk2w6gB2D6/l3uQ4tRm7sLOejt
Dfahd+APXHT6AuXnvqBQ/HujbX22xvyjIGPtr3UqA6ujcacMrlpuUoO/DbSa306P
/VJYiNH9BoEtXqQePqmK7N4SeeiiWJp562Mbi15ICfk7kB2EsPmn0pAQfP8uktxd
WdHSyCuPoimxEC0AiqaX9tv+aPeUtgzbu4l+n71WDFUzvOnClTg+4ZPRqAPFVtMt
6r7q1tgTL8GMmoLKIKghdb9AzxH4m4e/YhjF8gbGMRPfSAJhrMgPDAETvcwGmFiT
wa8Rwg/8DoufZY2Nx9mbr3XSCYBla/dbxt5rqYkwjZ4ITWZB6gHus+x9PtYYZkor
XDN7bbyDHHLnmXHRNAt6WvvPY92NuVJOWTZ3LA1+BKJtsy7kSHvPKIWPTx47EEKd
dfCtv7AFjm6kPFJR223i29iHgcgGcrB1KL+2Yq5Q5PCaqLujJ8+M2M0KM8wMOSBN
wqCn9Aim0qp09CzVTU2gukQASu2bo7wh/q7gh5eXB00WrH0Ajy0plu8fh0p8pNdy
qpZc7+AiFzqJkSTkQkvRN3aMkrg7KRfNNfyaKtdeu/r6gR8BBKo2LQmDYB1FBdCO
FsmBs5Lk0goHBKDucSd+YRJtQvm6tF2rfJJkeAjxVBSGFrnCWI6Sv8HnGCgKol4p
mWsuxJYBmDc7yC3SoZ7cvIg2Aqlb2uQNy/13xY9JQpZoT5ggwe9gmfUrYxHrdnsT
pqaCKcsq0U2yRExWq0ZpQLM0C96u28eXnD3SUdJNO9MsAr9OkglDPMg+PnkBHM8M
SIgi9qaSH7kjWBsAlh2hmP/vyZUU2YUVi4CjGVfqIxXOirZM6+GPxRxCAM8u5u0W
ov1X1XTwOsd+mx11VvZMG5Qmf0VCHjLAxwrWITHYBcpyiq3mDdCnmsoJ7vuplcLG
a3JdXYGwwevtHXpbirhyU0LuqWtk8WCw9PI/xg0kr/Ng3XqI5aAe6/fUccY5GTZp
g2U/ZQ2oDv/hbQJUesS+BL4iTsfMQQZtRTEZBgLxStQ311tM7HVKNDUs/lioKxI+
dUkriCSX8Tp8QUsHzYZXtd5IXl5T80IMQ8dkaHrI0N6rcwN/kuJtWnqXnrUjzBT7
QQQNUp6PsjFLz+IQPN7w1zAURzrI1dube894T128B9N6FJL3nVfs3bWb2rNKw2OT
OHRwdYINd3XIWtNR+lJHDRCVKdIl7EzQ6kQVQOuQ5PxIQuCMdnfBjn7yAJ9Nr0lR
ciCN5MzclF17cUnAkMBrdCt2e8aldfSZk4v/BCoM4f3mf0uCOZ7xO2enD8zZub7a
AVduL/26RAh2IUswWD0sz3ibubE+wVAs4uivPpQqkevbmVOtNRYehM3zZkS9CLNE
RjzUrGNTmyttEq5BaqSxhz+Q8l7Iu4fxOZ+IeeI2UAEQjb5IrBhx4shILwRL1KJa
HtN8qbgT6dSNbbKHs+NnYbE0dVThG2zQ+n1egm57ld8LYBAmqLX2rjTlMyKRENDD
sIU4Iy8faTzxWsYvy86jKwDDrjBzpWjRXo9q57ax6Hbsbc/5C+os711p+0y0VH0B
kQ5NfiWjszQMr/XeVphVLRtHNqgpOIiPLuUeg+rVZkraNCZMlHuF+WjPRT5tX4aa
RY3h16vRVVeoh0IlT1rC9R1lTg5KKNrPY0rt7g5BGlnqEtatPKPEvFvy8mprSzr1
HRmnwNRizwrxvbo5PpoGuQHupcQyASR8R1P2aj6ZIPdaRXorAbBl0ApwhG9wM9Nr
uxETiZ56omXwj8hmdsrXx2e9S1x/R6axVWGA/MjoTGBeT/K3+BaOioukT/P4hQXe
nkg9jAJpUnd/GYxZP6+jytEO6qam2YPzJn13ffAWPZYQNahNCDuTG/05NZSlLDsq
w7Dr5ESgWt20/98j/edbSNTdNrf1vleS/UZDoB/biMFMf2/iGBE+Ln9fZjpdWlbZ
bGd1KjEKaJ7xQqHCwJp+d4moa/HjIGKEYJdVWUF+Axy4z5BnO46IwiwC5xXtP++2
YvfLg0RIAj+7jTqy9wfMhL3+RmrkTpwPnzxAw6d43L7Q1JK86/kIqxUoajc83xoT
bQVmNbPWExkKH37JSwGqebcSpbdnQs5YDJkRxiIqXbXNZ+Gx5L0onZp6dIi5/nIa
5hi13KRI3e3vlXlwVDYfu62jcnWaQoTWoFE1iM6o6H261RzGYAAQ5Me98z0VxbTL
IZDGHEeM3XkkDN3BeJpYK+DdhapxCyI/H+LRPtSc+P8zSxT5hWqg+JvS6jkI6Kkm
gj2eLTP/FeYkgjp+tDH2QfMqZNl9xL3lUlusySM0V+oRWsV+rv6jbCZeZf4HDEqB
t24to9HTJcWfJEJMx78wKOrVOYopDSUzCKxtxNlxw4LicRSMD8cBsphfMwgsN9mO
EQoiW1AlZjCRX9l5kXfYt6aOZvzx0OUInH/whowodbSmKg5U9ZVp3ulWiZFsBQm0
ikLiOQ8ur3BFSFulEfKf8f5oBKDDZt5LjR/XJWiLsNZPm5UUVGDz9pouTrGhpRrg
eHwadLqaNR/EvAXP1ZKIR4aKcnnH7L92u0InrT5hVBU1euDRPuvnDlvscUMiW8kd
RTSsWsAVQL4cRjvLWUc/Buov7L62WwKaLARrBae9bu+J1dyq3LVx+PQ0Q67XvDUy
3BnYk6NpSyIP1sICgXad0+66GOb6Ixt2R2MVGfLUAa3lnSw6niCBxXAj50Oswh9M
DqfWNmYKLzvdRQMjfCoEl6mAMfNEmliBVQ1Uwhk/Qq3kXWEqpJfXNq6sNKOJsmrh
cjj57F4rHlPVzYDyGAa2JzDZRkI8oztZKxxJFmztcukln4/6ICdsGXyR4Wd4sV0D
kd4yqpSJpD/WvZsoLLc7NAn2mOGr9oPhR2az/Yss5gXnnXf93v9V3X0ldvpY9OqX
YFBTw2+FUf4Sx3g9mxX21UWaAKnF4fh6gVDIucMAeNshuoV0YfudnSCNWCoiG3Lz
k2mH6Ad+O02iwzjz0jt+oC3EBLXKrK974KjoTuRlM07AfYqpt2tMvqkULWNU7+xs
oZ5OzRPDl7X5vneTAHtoXPokDkJ770reGv8tKfih5Gg8NGHerj4qJOhhVVhA0U8S
/wbeb/iZy/bJ184EpgpXf50veCQmPI5jFddUu9MPyKClAKfOc3dCn5g+af6gH3VE
dI9PsGkT/1US4f6+JxdC9rT/ENtG3paivQRbYSyNKspJj5XYz8VT0uz0Pwr8yThE
OT8kYqGTXQ/uOLOqJoyjP4ByGjHKeXTWJsTdx8olUu6p4HGOi72Xp7Jb2NPevqO+
asSMIsrrSGKzz+h0+Id1wYEmokWXfFjMgDdbnHWCrcY29fRaGfX7hl3MvjJCZzxy
9YzfJriFllFe98heHylorse4Huy5hxoglw0+KVJOUOdPPzbZjVRrK0azTEEO9wBJ
vOPkxzVFlbbCJJnwRywJwhtOwTTfTy0EGsvhWKIzwAwD8Z8Nl9xhBwVxlpL+O/Sj
RwtSIbGDhXm72DD/537LJbjiUmyuyotAkZHdck0c/yOVQlO3Jvtu6GbqcvZxeVm0
51WTGQyac4GFBA/m4xxvVr5ioWBSxhL294s6RJPlmS10ZaBjAi0qy/nlGEOjvTdO
gWuEyadVWUY6mt6svs1TY84ILpjIuJz+A/9o0A/V1Sgzs3xpD61gVzPFanwfxgUQ
xdcju+EWuZsrcBqQYYtmoZ8eTMsju5+mkB7/+3MgMaTr8jDftcM8spYgcz/8BtIL
Crq4zMWIHGlUGb0Xj6dKneGMvugIy2cLXoDVB+QEy39P7T79DjTod91+YhIost7d
H0OeHAbzlyTEtnp9z2lLITAh1c4qmrIKebnojoleDSzDhCWwJnIaL6Kail3/yOdh
QZn8BNU1MlgId+Dv3vdMQa8uPxCRRdKmIokGLlfxI0vvrLVXixFr19aEU/pLJqTD
2ipKXIRLQkZXtUkiXCvD2MK+nPWIO3f5YuyRRxzSYVURKzfolXhubnCKzXaYO7TF
2NxoSRwXnTZtdWKSeNrL3IIeKyVsPUoDP6eGSLHMxCfu4/B1ANG4WD3G+8UP6NlA
RvoCT0c8wbwifPk1QlzLRFmk0Eos5gNo8hOobjfbSxceUMorKetbhaWdnYRONwB9
3cprjQAZdUecogesH4/E+9J2LHlXJunGW3GJpVpvkkhaURkXtq2pdwZfsBLPnJxo
fcjGUZR0H1/NaHnBJ1ZvxzVhXPtryfF/jqgxjVaabrSjHKqBrtUrAe7oearrYzOd
DLvkD0irFuhUoqAgle8aU/RdfjRrtVhpmJlDobC9PvuXnfKdic9vYwKCXUYUWLkK
amMhC9Fe1OqK8k1Ymb3ElZdTliJpdSF+XhYjQKYp6qFG+hiGDRhNd/tXOzne/bu1
c+x5RNMVdyKVa54AjtCodWLwx8AO9Nv94fe82nWe3+/J7WNMOpspy/91cocpO+bH
33ny03AWFqI/k9lPsBSti3MpOERKeWiglBtD6WlDFEPkwz28Obtxnfn0yhwPKT+F
wv2Sp4uj4OMjnY5Zu+FXg//6Yu5oEN378VBz+MwN5P90u99g7VOEiS4OwdgOlAjg
Osr8nIFhZUUIGWh857zNG1r4CRo9SLhaudZ5d56yqDs1nHzIMbLpTvCRDKgZDqTl
oDCwGHKdu0t1L9ySZmfflTTAn96MwQxqZu+kTi4xCuf72RMDQUFZK1aUV/2I5Vqg
grN/g8876PTgavh2Hlu4fCUfthgGx7c/P9zl+JX34HiG70Ze2eUzumk3VuUeiJe+
PJihJbq2shWLkY4pTUWhjjqnwS4JmxGLrW+1pcRmyi3d+ZuDWSbNQuHM3hBIrOdZ
QFfu8Ilh1UpIcna60uh1ZrtH9lU5gFnEZxcosmLbTnKy0d5w5N+pP6O8eJGzfixU
cDo/XYlCQcSImdmeuqpPtsbGiTm5orTx+JGRcLdrjYlcZifCFQByahG0lIexWtcL
2wn8m+yQTauN6EhqfJg0TrIP0xsNcbJiQAqs5H6vUN1qTfxS+3ad/sV+IiT64teD
1KdEHXc5STfqmxMhsgvbJzexF8KfIxJ6/GA28/EESJL5+6Jit3e720ZdlDrgpGNK
WmZXmv3TD4CG1Xo02BS5djlpzwgYRfmVhz7Pj4DUAIrGaQECtW85HC2UidAHd46a
72UwKpMYdL7NKjQsaCEc/f9A8VSNi0h1kirf4wIwzY9SD9jm90vQyjIvkHmJKITa
vkQgru/lFhQKLequEkNgO97Sdayk/M6hFImZXzhR2bUbs7RGygl87m2ZC6kk8LNF
/zYj/a4O7bIkDNBc6Ri1IS4MUlEVYbLxifDa2QfBi+tMwTdZY67+pgs5pAI/mosR
lJXLbNVyZM4Bw43Kru8s++tQ/c2D9LA8mjdBsHZPgifrCiRbBO9bod10/gaVt0Ae
UA9LkN+bhsuQn7C/basFoGswvc8tkfuuhh2yTfrBVt7p4LPeZSeDuaOatYtYwXlS
zWnTaIQHM4O5FqWYYLPZw1Syzi1tpHBMVu0DKsP1FdHqvwA0INqrjpngHkXW+SVG
bBgmlEVc/EY9NtWBAISlDp5VmaTFm2B8I3BV9m04wCN//BLh2Ktna5MMyMZt5ldK
rsfTJlZm/HqjYcojJp/WkhzLk3Z6ikL/S5JV9Z+VtBhKYQjpo5dyidH9P/VtNrxJ
afonao1VOtdcuHcINRxyx1/eCMFUCUUwJI4uqdkxLiiCAkVceAVAQPXpA83cohBI
N6+9/JSqtaEAEe6ya5KT7JrX3bTZEbV11e9Pm3UVLQz83Ope1qo1MdjS41IPYOqM
5hRltKqWOURJA/B3Gor41PRQ3/U+MOyozTROCz2J4GE9wGK7VEOta17+Q432C0Nu
LTzGgP0h6ypCYVezDX8lC//fFOuHOtyMxJcrCgrD8YK4T4m2oObs5GS3O6gmMRkK
aAnOm9LKCvoYbLc2Hp6Dw7yLbTI777xHYXvr7hMa6t45u61R8KRs/f312xFzNMgE
9ZIzdDNw7UOKVY9djKkletszPdPkalImEcVK6pdU8PEffPVhsR2H8HNszu0QUZ5N
QmqR5+X2M3Pd48jXbv/L4yQ2CfuadS8ZmRmeGR0siaOUbBPUL1acI7B1icHnSegy
aLR2FswO5DzXYImTaGDld6luw9Ud+MyCx9db4XPUkS9pg1v2ERS1ACGv4ruTbhAn
kDkfNFjtwy2Oqe2WyiN3gtqsvdPtaJQRDXh4PjxtX8cK95PFlLaJICBxvGGUe5ov
W68cT9l8834+pmnki+R7wKIga7BeOksY1QszJTuuU7hU5xS705iZPa+LvVqVOWfv
Z0WgMcizxqC4tbrqRuKU/gdkblqEAfFFpBw3i4yArp380kNwa3KV51XbmWf8QZTW
0IcpVtpLK5PSrE+RWwHdlAhGGxe4AmR7CtQoFCRr7znimIDJM04ANzotW4qxLA6s
IiygEHrJmhnTXWluSSuMC0Kb8CfOCI3UaQ2RULhBIsLu/MqJ/hTkDBZjbgrz52Xv
TWxDRWGrzNUTSFTt2UDwGHB/YnnrrkF45VKSTt1q7FbccAtJJgvMJOTEVumioxZ4
55i1c/tvrsQOwDdjl5TDe8AbHs6JTBU5QQ98qVB8IwJ5YNvQtK1KD96LCQPu0xXS
+ZNckbNyOpGCU0wNGYagG/Ri92wT/hdiqO8AkMBoUhhcNJyfLS8jPiL0v6yM8nkS
gIOPBpHINiHgBJuLGwaPPykrpldSn7r37qUjn4KYFXxUSMddbffK6lSgCqWrsRRP
5uwW9vI3vRP1D+lQQZ53iX0g+ukm0bA+TKvXqefEeE3QDDq4Ol7fCIC5eJqAw5lk
cd+sDmeFjivmxhUM6jPgNWdzkdbo/YbdS2YY5KkTzAXGn8fwPjWmwjw091/4eRoS
f3fqAQkZBgja8jN8zy8EodZs/50p8qpSlcVFtDslsimxbI/Tb8sZvuMJxq2W1eT2
K+rQe592ZAmZ+LlMx9HbxA9pbYOJ4+tcJ5q29wiHxLBa4SSlsF7fstc9mXZuTU9+
+3o+SZd99SEfeXt61VH8pLevYF/bwmAqpq5UAdO7U4lwxeYIxWiRgXpfR/7zT8I5
a5jRTW11F36TSch4xKLu0dAd/IAWJYVH0fZeInvllMR5WLsSgyy5gMMLRQzr9tr7
HifDPxLN06iHo6kfF222LvTjTD8ITtyZdKip09nMEBFLNC4G0hQDQ+X4VBo5pUvJ
2EDhK1hHDiARQCq1taib55Gros72kfKQ3OlGtVIV+Lz0LrIiH43o8BJDsI1+/Q6K
fLUgsnfpf43IUhgRmvamamNws7z8mHBpzcwkj2zVRfkw8WGfOTXh9OXjyeRUffcp
OMGeLO2tXywHkP1zcbGbWMEL72h73KZJDxxY3Uy+ASvV22TBQnoM2VQ26nxIxCPE
Cb3MJUiVYvOGs2/zfw7a3awHfC6ji0W6syy97WB8DAkQF+avQuBiQqLq2erJdHWN
ye0jReXnUBlIvNWQumxe6+IVoORfA24z8B3xXLy+TirGX8Zl/ckUxd5FDLop82Is
wFY7EHtCXnuk8Wmd8nRARFxPE4+AYD23Raye4SYr4Ew+r9O7Df6X3qRFy95e6PR0
vO5KXQ3MiLWT33UZ0xYCXH4XPLm2u5mzWtK76jXOVqXaf+8jaGyKTcKZGhZG1YZM
9lm3bO8ml1dNjTU/Ppkg+ApTeYWyR029luAA7QbqEZPDZ2mf6rugacszUFUIwoK3
NgG1xS7CBSpc0ZnpbzFycpFpWJiQwR8mtVitQdXjGF9IvVSwwOlCagGFHbD5Lec+
8lxpoyHlp8oRNXMd8dfsmARSER0IH+jbFNjo7AUzvt9OruVe7ZfSQuOM1oZmQvMH
imjL/TCtRTn6b3LH08blO2QeATuqfGMe2G4QlWFQdKGUy9ZRnwPi3zIc9ttoE/hw
jQgNZ4oaPqKAb9I1tZd9HTC+i8nsb8LmIOuQUmr9B8ptUP1UpF4HUQZkNXi/dIhw
hA05bW37SrkKtqfyPWv/EglXAvoosnGNK8a49Lffyd3XKao9BSBPonbWl8jDPo5f
+EZtQlG4xi06mamH6SgnQlBEayz1zGKaAirsehuuIxDA7VNWZaVT71EQiiag/l9x
yE8Xltb0DVshePk81BMRW/umoVW4rWR7e7O72wDav1mT9swmj9SRyW5J6msqS7UC
lW7RB1pI+/oNQOA6b4noQYXNWwxbyt74/v/LVd/Sr/MmZZDQpsKBrjUvYhPj/oHc
WrxvPTE0jvuqBGIaWQQaMQDn/vLo0E17KZiD4XiT0mu9rw7BpnCAZ7szKRp2scHf
J7LN9IQTTDHDSzC2kGNh+afjUIwGlpx5vVUtwpQkno61jGR4BbW4yF7XJ/0G0LkW
kKnz6xgjipweq1Q+4Zj1QWNM1u8Bl01yEHntibGWwgPAo7Ua6ycSov133cEKhLLW
WnMvbavRRzodd04Hbp8g3qSw8mdPM4Hc1cXUuVlEXukyO9W2UFI8WKBZ9AnxAREg
BYL5aiTFEzsGMDFYakOJlecgHVb9GMvH1JJSkJy/+sn8PE0WZtl/5LFeZLqKTuqN
Ym/UOl4J6nc1qMh6xRj0fWNFw6cJmNF90MyBtq4kzkDEZqrptJWkFmRrYQv4hdNu
YtvA8Nw0WmVZ4ZWPLOwtLJhxza6khK8Coom0RkF8pGvStba6YShBeuGPPAoVPwT1
HAux8cDUAu9D+G2V95cvc3hjW7cSThPk1JpEM6SgPc0TNuHyHRf90TaSSLaacSvX
t5uwEo6xkZTgu6l+JIiXjLSTq+HX93QhJrMmh06L+HkVSNlMZuZIG2W3+Oj8DPyI
mD7rU4z3lng/lk/SMOMIe2o3pvlvohzeXhkL+U2jXbWmrkDnybzb03uodmA/CaG4
gs/gQ3FZtw0bNgQrJMETOWb2+jXdmCPOxJsbFjlRDYauvO1Y/xhmfpNESdI+VUKf
GhMz2bND/+idH/I0n7FzHuXRjy3MOjE6n+m9Vy0tymGRfGrs68CZ4wPNCBFTgw5I
DtObq0Pvf+Y24tfLwwFzKePrPijxHqP1+8FdwSBxMbUjfIylaVTvaNETCkYaFUAX
YEnXH63CBGoIdIJnjD78XBjMgdv3HZZ8P8yqACJITyenb4fq9GPK62qlJZLdvnU6
Rv3CQt1PwzEf6JDVUriVOB4Je3iaye6yazg/xESglkxkXbyLv5AFdd/5ZktEBWQg
KQQEjIqntIMl6GqGTIk1McHTwwRJmdVRPoWRHNlnmZj7ohM+e8yaINqZK349cSQ6
uG7DL2gPs3QwSLA4XInmbeH+2Km0PuxCeYruJkQvFdcz7d292sXzkfjNWSUS6wPA
2IjGMB6VZa8ELF/8FDPEKsW5G0b/UeWWs1cLie6gVawhcJtcreVLrXo0jnMbSfvk
iycky9njAV9lAdSsUNdvDiVgplA7GUbeV8/zcdUSoCTAZu3GKMAbyL4BK59ZLnzq
UAz+6J769TUN3Fwy0wbE8txa7FtY3Yi27hGfX1E0BCXmQkv0LT7m88wOZX1Frh2S
LpHTDUpAE/XUO4rA4UqOKj4/XutxLVnw2jA3yJwnEn8+eyiCQQ+wW9hH10WtgO8/
ffurTTt7KTlWxlqHI1YBm+FLwFRE9CxBjX0m117iTCRgH6ClH+AVIhry0yja1XMI
dz0lIb5tOzt+HMQlslF4UD1V4s2VzbtI4Xg/lgRovkfXdm5TY5+1hEcBsoSz+Oxf
X+x9/yTbqQQZzZQrI4veUU58H6QFVvhsjvtO4WE9ieQgUlOYaGHMmhC30hsCaDeW
N6czbpTvSFBvhGXsO8ePKx1+RoOWHcnwEn942KnpWkcKpfPNGgaDCHfXCM07Qq8k
hOlkflSS3AwAHVn5ZmQEWpfABWOcDJNqlYi00twjqIrpxyk76ornMxjIsg+kUq89
wKgdD0U1gHRJfC3t4yz1RKjvmUYfJMYwcExk5T9kXd17k0dmFtMAA1D+9zm3fLOp
X6004WTIMMwouCcGpHWabva6OFGzKl5kK/VYD6a2FakwMfSddg4asDjfonfsiV+u
/jwwKtdmKh/JR8QT/nVs32XWzO4on3OKT7E5+9oM2ddF+UJZBl6zveUZIBCKE+Mo
y+4kNHufsQsdvBbaRWb36lrqpRCG+aZyfD4eMkg9Ig5at/X2EZDPmUkCoj+gY7E1
4Byz7x2UM4QkalOU8J/FhGvdcOggyvFQkB5N/0X0bfMFEdF8xzjcYqTuoIfHfO5o
53HXfj9mU9srJXVgn/1yvT3Mz4al5KD7XRo7FIFjsFmHdxY+4qso4+MPc3R7tBdf
Axf9tLYwRUhKiywirMRfZ/rkkNiQD4FOw2wV4fn72WVjNhKxjdl9FVLXTXU9Sayi
lG0QynkCZzSRb3u/r3W41RiL+kzfQtxK33KsKFd9i8e8ImxHSfe4nXQOdd7iuQ/z
gVR+iZ6Sf5fqU/T8w+E5W4tZZwc/Rat0E9gHmiL8s4VFY5cVceinjqQ/nfBLHo66
IUGoVso0iJFt2Wissv5nf1sPyB//A1BSGyxVqvDhXJNW//Gw+uLamtkhWfoSGS/x
QJnhR3v62Yyufb1OXz0uYa9pI+GxrPGYQrtYtQE3PlRe20E4ECyP0WnJ3SD2Ihmi
gC/zRqd2ovhJe2C93N7vJxvNPxEIPPhTqHRluX2u+4gTzmhT+C6U2p8vrGpS9yIu
mC2KsY1QAdU0rwUhPe4MHB0/cfx68PzGyt58rf9ORAKDC73n444v+02i9v98bmyi
ZcTVgugeySa5Dld7H6hjdFbaoZ8w3pWuwPTLSqvVlKHYr2Wd9hQt2JANMszkEZ2K
KEuPpkUPaoXR5HAlvwrBrM7IJzV/odZrK8LdB7PdRyo6AR6emtRBAGUcCZD7x1HQ
l6nrC/sLyn4W/MJ3R7SVKy16tCThVoN6vdbdabD8Br6M0A1jxILnHSdJx0D5a5Uv
KWm0zmbIRUIy/FPo1Pih/c0Q/JGuWXiw4CjfwytgOwZFWxkoW1kCxTl8BheSqTo+
y1jASW89CjSnaI0L1vXQDNuiAkuOrsL8F5NQFjr4Ci4Y4kKf76DvqZ0wNV5oyhPC
Zt5VGVjPUbF9qWahPUIw6+QXfzkzxfKUu+Gz6mI9ZLSyR1EFiUMr0CafQ2y2IEgu
kppiZ8xTNa0K+GL4z1mMov9Vr1MNO6Rtg0jHNUX3xfdqMc5RUHfAlOypV7JPlGE4
lhGUH5VTXTvPtkqcMivqfQ1RlTwAXndWTDfPsObuN8NfMCGwUyBfnAX3U+m1zt50
ujT8ZXE16ADhoeOlJHc/NLNHApn7xzvE7jA9oIkfZXZXck1THIIN7vbw5j8+Ggiq
oALq8iurAWlJzm1dZNuLo5ZFprAlE9O1oG4PFKjjALqetUMNA1OWMKWISwX3vEkS
OF78QzpbyIApwFAwK+zA2prtvlnu9IcK6LGfNljREimQtzqYXbcPU1U9KOxuNoRk
51wO5Zu63hC7bTLiX2rWobTptKFMggf9Tx9SSwgWpzbzOohl9iL69VncEjSFu/BP
dvAN1dWEfvXWRivu4em46+UTs7Jl6cNY3WviWfuPaqo2J4BaLkQ8aRZuvy5PA0eJ
AZJ95cS6TnVEnQoJkxSAN2g09oPgdERZAG4ks215Zj1rtZtkd0MgVONUPgLmejBu
a2/i6GxNJs+or7a32gA+2qOT+I2q16yCkcBS55qeC26MUl/goyAGKflQYfRMzEcs
GKycaGstYayTbmTva0V1piRHC6Wj/LSNJMQThuO5y+I8oedEyUFBTa0hs6cNZwX1
SQAB1bwKk9BDxwJUNEClXX0QqjA49ECMTrnh5rRlUemH8nlPnlI8OBcnZrunHBu9
SW2eWjMDd4RFdaWa2cVotk/waob60wk6uktzlbmr2aoZDPVgpnfdvcGtsqyL+ATW
dL+cDCWXwpCvhqSXEfRliuRLZ8o/66JvxslANDzxUxUwtdUL7CbtEOpmUf8FT0mj
9n834TGLPERcKWHaTe6BcFb8tVsC6stWUmDmb59PfAfAzSKJZVorKptiuSJ0P/A4
Kwd7nYmTrBaluEleg+oOwF2gh+vbtODDEHXx/frrUQa2gIlrLVPs5ZlSW2d2yai9
KQe7+ODQOjvku9pl3KnjocP7Kci6dwrIKRZyzrnb4+svtIrndx2ZbbDWGHgFidzX
2f/ziSZZKybyfqnmJMp2fcxFkaA7rAc/5QNtnBiMxQiE5CKDycZszCWojsU7gHEH
Hve8X0ddG3XAoTQ7VJI7qftefNu58FFISOfanmdhghFxlctgBR0JPM4SlzdiEqlW
w5L4qJVI2g4Mdx/kNcGcuxS860NmMeymglyNM9HjA1azeHnYvPWq1olaDODutgw/
00Ha4GWBqIiQ+/WKqZ0pFVLSpBEp0lWWuJcMRmmJuSRMCfaWAaQBA4utEEVzeUkl
ORbHhqFGCsBOF6PM1BwP1pgNmVkaPt0AdYOEXhgMDsR+aGwpKxHX68BvAfWEwslU
UDh8F9dcpMaMBNJb+6xCHmxOm1U9yLyItnJ9Jf89A8/zw8M2+7hfxbCC6Xcl9ZUt
9D2Dc8z/gv0Or9cOL9emu/MUipukeUE0lWSnhDp7yaTLkn7MDQo7BZXaYpFTafm8
t8QWGDcIj2Bujesi6P5cap8ZHoLxdTV/wMi7zjInV9UVcgN2rL5I5vc16QZyvA+H
djKhVS4nX9cQGJOiUupfa6UHAzbCDU7IRgHc/U4zPh9Z6XwNzAkw5bNGP11PDoTe
eg0iGk37CCdsssQ8q7mXAXWqk+4Sttrj63dFwwR0t4ysA5ImXwuqMK4L3YGVQ/Hu
8Oa0nWhDpmriVXVLEDyX9QRxxbQu6a9gfSxBrVIQ3z3EDcKh51G5uuxB5x4p85TC
PfgkwylZULxx/nc/zPLbSz5ong/SUY5EPEe9m7a88CRCiQwE1IqR+LMldZS33uar
PQCNk1TYYLi19HAWQ+C6gJYdPv724AJ6K5MEnUsLH6Y0xdRChY1gxImqLAxyV+/m
cdgFQuzOoEWlC1ODTvHba2Qff5Ag9PZW3QFRRgaMe25Ut9RjE/CVAC55c99DTn+Z
KaW5xm/Kz1K4Wy55BiOhcepApuoMARaFoGVv9WhTptv657sAKZUVr342S8WRQ6VT
dZH0c00e1n47us1kiPwZXhmeqgfghxhnrc6UDvAqzcGViV+nXEmAnuttwZz4yyVp
UOsbWEipyPRRVk/VFWpduvBixadl+Tf0j+W7gtCE8nZq/RcNKOKcYavAseYnbkq3
97ZPU6lkC3/KqKAHuqyGA2/Ojrm0Akc1EPDcwwmmY4GXOccHQXraZ3avnDB5RuS4
m6/7WWpJRgGzKnQmKTqm9+rmgUfyimCIwVAWbFvKMpD7Bi1Fjrt50wk7rvOdb1N3
ie6gCyUEYOnxuQ6nQ/zPhQgj7ky2hLz44eJhE4CXrHiNvPQaojglDOSoRL0zaXnK
/NCxHDl/9Ex+19Z9xCfw9GV9RZDASRZiuEK4ds+iXBC4tUyHx5p25Y4JcfObn5ha
eif9dgP48Z4YD4ZD3zd4YH/Heo3I92BBojodLuCrsRhjKHhU3eNl80iVG+Qv4rRT
LJkZfnWf25HMSyZDI4/5pC6YC3B5TtrYs0g+HSbC/1JvGKFeK6dw4Y7YdcDpsrtM
fW36mq51zgcRmRyOd8jksFA+NE2KvL//gdSwdbOhSF6HeH80YbE0Fb1tPLx7WUTb
7cS40DrTkpI2pKJDXsGTkCwWRWpHKlLe4M4xjD3PP2r/bqMpZjXCD3+S7+owGkNe
eH9TER2BfOSCebIODYC3YmECuyAqRagj5xMgb/zJxwyLDcdrHq1z8fCbJgfpUccn
Xb+bObz3x9IF0LIYdiBvHbmmV6M7Z6szzK/WbOg8OdL0EMI2bivQ9L54wzQym26u
Ar88j82v7gAcGacicHcHR/BaVN6Rkk78ivem9MNXXyMnfhngGfizPX5VasS4atQB
nKWnvVZrFaOfDDysYXhT+EoQI8Jk+yzSJHLr9lpgX4bC0fAHOK3HFb1ZRjlqKMc5
SOQeAHui4Yyxk/nzn0GKNgMjd7c5iUl76fsJpN9uHy6FXE9NjIq/RBK7tOnft5Qn
aNVv8Th6qVhpWobJzYkoLHdI5u97RiPcd5VaE3fofxv7xd98SMG34W4TXdgOiVSK
4FxZ20MMysdx2RyUOycujDw/w/eDUQaZX+i+e/JzAuGDRxBPAdIzAlompdHuv8aR
QdEtuHB/XcSGhtd6kf+LvipcXnGdVpAG7JY9SbhR3aOUUW4RrBzSi43s/+HoWGOy
nbbEecIgXcBPS/yBIpfn3hRL+30MOrsLByVnXYx0UC8J6Xv3g/EQTEiBiw/70xi2
xS/7VzWVI4T5w8w+c29rsig3CiuFvEu6PmdVqgI/pvjYhKU9rske8dxtyTIh8VW4
STuY2NV/CHpvFzap1FWaEcg9cirG2rB3zpxLnTK8kdsbl76lwRgz+vhxSaa47n+i
RPrp1FY3q0izCkzs9slcQMN3tr3he/zMhH74XFaVrs5QaEoauOG6q5v3Z3jfPPmm
wfu3BPtMTfiJbZMjLBFMpQNPmWHqZhaUNEQpTc0dUqfHJELJWFDJtwJBsVWebw74
clP3Mr8BvjaQ0fqS3Zz3tE9r1yVfRSYqQkcdPy5QSlxVdFUPKbEjwR5AbBTtBLMC
/gPmp+/siHOcZzckjrAhdWwRJioVkGKcVWf9G5kmeDUlfKudMgNRJ4HUIm22MFD+
QJt34SAy9pKtBVFjZ/X0HCl6/U5vnGNsRX/qBDmVDymUEHXj9rOrzsyl2M1UreOy
qE8qwT0dnBE0c/s3kyCBcMeqjtECxPxdVMQgmnt5qtwlxAjr6ejRQ5SuHMa6ScVr
WAyb34XGP31ABq9lQOl7avLZ7m+umgMXQ1XWaA+TjDnT6qp09fBWn5dnDuZwuGqi
LNE4FjWQNOL1F8i34Y6XolSGcro0G7YXCpa5UGxZrUsgATqjE9qkuxzng5BicfSO
Ycr1E8EVuQLlBlf0sVgQ3fMz3KUnbiuAYNdx7RHyMH0110zfZjF7nsJcrBozeKbr
zgPFPK8bITDRLmdYHuj5qKzBzkbKiTEqj+WLUo3XDJobkm+8WD+tcr7ka22zcVy0
aeOIPb3QZSvg0ZQ2IaLRYUz5EM+M2qqT4Wav94GxXKUGGHNgNjAIIKkKuAFl1btj
9HkMzkDKqVISunbPodRUX+3ZdLRYVjbMeULFS+3fcTQrehBrFT9XxHOZetqHNRH3
OVr6OAPFM8IXQjfQVJkgZKBWfJTvXWyP+xmbNxAbQel1m9PF9IlpQAku051agmrB
BI7cJpzgRqrCd405TH5H0PE1qyz4hpxXE9iF7JBXJqWXf6lmS823BqxILjj7PU6w
LOrIXkj7X/zmqWIAh1X3oqhwOIsctnYvD0hrbwhiMRncCmG3FSpsT1ZPzP50RVJk
nbVyWUVldkdu3/A9wE6gx+WeyPWlgpzL4x/HFQOl1B/WE/2W/ABEqOfV0+/pJd5R
cNXaCUe1497RJCCfJYcmM4prePLl4m5zS5jsKdBpIMxsPYHl6Xin/9bcrKN44Tum
NjwZbpQmXvijxgsJm9YkvPtCkZkIrZ0ak+fJSg6iQ9/98tR2PSJpO0APa9muyLUk
HFzH1gG2mAuvD1HrCAxfNOcJDSSWf1gvpDCwJ6lp+HzvLVT5UJaHyIKzjwwOcqQ4
jTVDfq30+D5hRim/m3Z6eQroTKlKnvFwdmsx9SjWHOBZq7/Y/KGwgT0/gIDBMqka
gCONRJEXNJ/yCK5VCkGEheu6eDp/U3bZa7HQ2eQRYL3zUcFzWNj16rBj2nqTWPTr
/v/0YbR8gzmYu6gBPA5LEGj7QzSMaaFOpnHlmbabWlzDg3Q/cD/sWqLjriexL37t
2dFTaFIqM+pK9z7tw3ZrH3Ks7HBcdpKnJ5PiT40q2Tym3/Bp5RE2Jk0XbsX1jbnB
j9IijK6N8yESw1ehCZiiZjGZkbzvGZuu1An4JiD5JmhttPAus2nVT+7FOXXNVPRD
lbQRJhsetrYkezmuB8gkEZxHV7ikGpa57LZ4oRs0q+VQ+AgGaO5a3uc1B3r2NsRm
8NK2soRZCJPlTRmiU27MDhAoSIQg2zwpuMEUb9Y3lCHwZv74jU/0ludOps8EBPQc
Vq+XY4zhg0/1jHwuO76fNrBq9uOyuhH2d3LdfSP9sJ2pX1DJjXwg8jmaq0blLuZJ
a6CmHb504NP1uhg8NzNy/d+ctzbtoPIxtyfsz0CM/syap4nMz6QxjE5NxluBDfSp
iGRvb7VGnbb7g9UbMJ6PollOH/O/8PpXO7fr40jHK7832PUUjL8VWhFxw/I3W62j
jt2nZ0Zkib3EEFqWBtT9TSnBdKlHO8Py16ygCN+kLHgvYjemgAJWqnpmA5e9Vbbx
k1CEGlqwaOvC34ekD68QLbxkuMMzErpKlUPcUsBJkSFmE4Wx4a3+AIGRfJJGS0Tf
Gn4ThGnl0XwrfeLh/q2WmN3XyhmjGuW2SGs3KnGWaTPWimJKeRIU1GJRqolYrQFx
VTZH1EWlC1NkCB3pM8V/7T5lHPPaD10SEx3Q44lPw2e1P/qGdHS1LjP7hiMumJIg
cUBNTNFLqUqV4vdi+vRPJXv41dXq6yJYWzI6kkneoquQS6UUVK47yFgej4oE8P1Y
rRq3M8+N58ZtxFCLzHxSiKN1uPl7aSAEVOUI+IQfWUtiRJ9o/lAVMIayGbHuVgDJ
e/OYzHFXR6yhbhFk0ijBc1o6Llod3qWsVC2B+QUMUsmiLhD/mcTOjtJze5Zgv+Zk
GkrdhwGwGWBtWFEzvuDeTuuCzGCEPObi+IeORvrJFV0VtDnkcG7D/tYevJnFjtuR
VMNwmXz70B/isTvGCPDEZhxwa7/KqG3DwkEG2SGjnAGkyWEFIr9OA/Ho5FtXg/9V
pctEOsyvz52g/8s3aK6JDgvDvqT2wJrbwEYbWuJCus/Yj5m61ZhPJgyzTouP9eEi
y6v0AZgVkh/jqLgv7Ngg3PKh+s0JVlgLNzmTvXCJ+PJhGU4mzUCW1MUVQt8tXrwZ
i8g8teO85s6HeAj7FT50deYZ6hgI8M/ShqaOon8AdTOu9OQt0nt2kTB1fw6djS85
kL3NY0ZFZtEpsYGA0VC2CrGXNmJcVdC/s86ywJCwrzt/hiT2wtg7q6Y2D0++afMf
p4WpuNMoqFzU4QxYo7Q2lz4MUrRhSeh3DnxLNIGLzaGFTLOKueXeyxuxaTNCkLQ7
ADA+2qNNCcfuhWdvNVw18IR5HYGq7oJ3iUNXHALalnJ56qyiSgSCeWpTUsFcb6l9
6RI8K+bANVuBl0ysgI70M32Ylr4418sl0AZuYdJKZ6zfrBDkAfbTf1ZtjxJSDJuD
gFzEBKhFTdWoS30Ye7AwNpA4auvOCTyu7ZybONr9D6c4WA3AFGz9scSLgUYwS39t
Aprpa+XrFOnTrM7uJIJPguFklKJXcF5i6K1wMdEqQ6VL/ZcxCkFjyrxFkTSW5EFV
yr+AJiKvi9kscON2lbHrHbb4b5J/83cZ3gMfI4XpbtaUKMRkFNSbkJPqw8by4Owi
5Ccg4sJ7B6LbWWow02hfySXGHCXmdk4TJkS5uoBYLOB3F8X+lC0d7sKQi1tIEX+k
E0In+B/Vi3OWpwg5GQqWkfVsH5D2Ve+MWKGax13UM+XMZV5zPZnA2/INihVzHQr8
4JyJMSkaUsvzy5w1GXZMMG/c7VpAkazbeTp8Okf9zAi3pbU2jPfT0XEnHoAxgw1H
88sDe+k6sSqSMZCLvzwUvKz11o4Sems0dP1hKaBffmAW6CGOJNmHtOpLFWTu+bJh
GF/e1teDJWb13K9RrvYmzSpjELQe4kRw2BPhKbL/aTWN9HOixPQCjNSN1JLcCkov
JpE81XEFo3FOGgvU8G2TRWHWDPMgJcbfWIIm3+J5g5We6QTLTEqtUeFVXdsc37JZ
V/vBr8+7bypcQfgemAQ6glQ/l+05HwYk5ZMCc2k17eCYUYE9SnM0Iep0svPw86F6
Gva55YGBOuhFXW1ix1kPLVodYH97OFDE8RnP0bFGNiH7J4JlrDrSk0TCvY2qMs4C
xGegXbbb2bbOu0FHahR4cgCS6xfPvuK/5y+X27BDqMPvggseJjLUL/4ZvysBjZ7U
npbjNmImzuP+opqO1GWHxE57RoX6KnJLk+2XtsLE78Kh5rLu1S5uv6YwkmeH5p2O
vz+N34Ym6lDafOO/ZjOrDQGsc1TOkaEN9jlzNSyJ/Wu/HEvrSBboXUx8BCE2NfTw
YDlx0GChoJ6Y8t879hKexAOU2+v1Jjf+0RSzYXSlF3GG5n7P42FWv+m81KKVX82/
bLBTxLDWaILBpR0kOq1Cde4cGCtfeW4TyxghhPpEeO00Q0kJff1K+zY73ujktuxs
Yr4pTxIwA3JNrLphO4VXYW8peJWvPIt9CNeOZtJoovg5M3e2tXFrHTFfp43Bt1t8
vP+QW2vC1D766yEXiPp2j2siQJlbeUqt2qGkK2RlNHPy7vAeyHqPCd1G/66TUk4V
L77w0JrLxMHyiGM2yZmhLCc13Yt3UUJD67sTZxwklMglU7zZvRqwixJEJhYyS6jn
0DSmYfpUE4wLRmo4LrbpTimuLaKRfWm6mqesWT19bAy3palpAk5o0ZaDsrxKdQA2
ulVJ8reXmrP/k8+Pg3MYjoLB+kiL+0ijCWvazGAKEoqWeMyhU9so7N4w2oSVPA9c
ROe6ZXrAkvuGZ/TP15AIlDFovUdUcgcAfj9g4Xq4we928q5kuR7AQZPMVvh6wvD0
sXq2PkrPirsFW51XFQX5lOxwkz8r9avbPn/4ibeRPta3q8oj76UVZGfiktwyUTit
+WZ29iFQWjng3fz7kTIJKH7w1z03mCu8LgGSkkP4/1E0jcclQEZkCw6kgtLSQsyl
Fe+JmkXJ3GZJQ8j8bNw524zT534IVKRVbC0M6gMLULFXmFBT7qttOpAzUU9gNUk9
JMRpw8AA/7gpZZYJowbNIw7dFtoBF7+Ie7qIUdY4t49kEnz+gOdDLWd5LX+uTjTg
X3KPOYd53p6rVm8CKjdls52JenWJioBrnNkwp5hYAjiH/zyNXyAx/i+d4bW4lWdo
i3UNZ9xL377INzaRV9KyemZ24CCHIXCiB5qUMHnBLcwTor/XUS+QkEK8vcyBlPgl
GwOCfgsQI9u1NYGuadVYmB2DtWXfMAs9ggZqDRp4hsgtSffB+DKUjkO+aH8CImnC
u/KLFGDc5ZK3ZzoMCwksKJav2tw5/BotEmpLekMtL6u0gID8eD0tiXa7MEp7qxaY
45++/bBj6g1qHJBy4GyNc0bogpM5ieTL7ebod7KC3fUCz0c9Sij49RcpIvRwvBYf
q5JELhT31vnylQLBfJEvhfORd0yLx4JWgJpxdVkYwfc/C2icw+0YG7Z4pVN1kR+F
/KXnqLHpC7mJ1qw2RPUNJYMhKFPHrm3s5LNkhlJqYLbjXBtter977lnBHyPDQ3Eq
9ZbW9ziEaHvS7KnExpLOQEG1xTsVDrH3lCpbqaye/+UVxroVCm0LuLsmEhiCrIeL
1md4mfYTvqyyYKoZNFIE4fcn+QpbWnit37d+uzDARoJvxDwrrOZFnsNU2irmDQ0J
shv/cd6QqlLkDDP20hUnYCCMuiQjOXbj+eZyukzWAfR3iEsweT6uhuOueSfVkOYG
am2Vk/Dct8csMUfHDuXDoTvgfSurCHo50GwzT2fdK2Ky+G47Z8mlDM0gUh/rDeEb
p/+C6PPqOTDfZMYtSU8i1E3/I8TM7Abyb4UXaN8Qr2Fe840LmyybFbGH17YU+X73
ffBm7lxmqALq6Uw4Gy1rrfoBZTw8zwNZp5mCWvihgJTaIsvkaeLQqd9zpLT4Gw3+
cPd/mkDUkuJF5bwsnQsNWbqtQgzKE3I6yuTdR98V+TmlPjRJsB+izHx9IqwDF8tu
rxgz25vvERM8AtNiZ3ieNjCSMZ+U1GmiWZt9zJibAXybDATyDoA/V2aEI7I1DLgO
RzfHMFP+Q+K1PkvV0R1hcREkzkIbUlGNrU6FsPcQHHj0H2AruBs3LXrypNE6Qy8e
/lRccS7kAmUzalzvYNdbYxafK45wKG6GkAR19bIvG2o2cdjDbS+5Dnxn727Ewz8N
DvXo0UAjW6UNmIH2Bn2Db7tECWeOb36wrFY7taLqRCdI75FeVvIvg84ld6p39uUY
3fsp2RTvqKDRKmXr6h2z23MYWZY+ik4TamyplanDKKzUvVjzZs+vg6usgBmwYjcu
qkCKYTwze9SO3alRYC8lQjt1QfE712YxiGW1O421wkqoBVoOrXuLhf1AzbjbUq1k
Pg03oQi6fV8xVgNIMEDl13g0K/M1WbvJ2pJm13jn/0XI1LkZqP+la5G2ER90hSg0
n9Ocjdg3c1u26sUQ+e7FD1l/VI3kJnshaB96R3YqLCPlMxgnswk//n+zibAY22FK
gNHkkvF/GSr10dbYuPD5wYDxIh1mziKrzNsskHVzS+Jp5gq4JKrF3fBFz6LCcHjL
8hdHE1joMQOMkbSelgjdpSlA1i77WevGGGdGIAv4ehPbN/piwWX1hJ0ivhDfC7k5
diNeBcKA309NmxUH1frQZ6auE9qvmR0Sl7u0tKxYuwl5NHM9dXUUR6AzMEnyLqA1
u4iSn0jQWDj3fNOO/n2sdQl7WVQkdBKryX7ZtbdtvxOpaPFNva1GdojZgL1ceyYf
4eAwiQU4TE6tKiCCNf5owRmnrHvySE2KWJtM8LwJFMZX9TfUKEJmWceDvLkJ4e6c
f8T9UxrgWv5scw/ZmETk6zmuBbHE7fADMjkGLMYlCbkoheLvyt/hU2aSH3HVY+Wj
Om4n87+ApijyQX/BLvI2PM9vuZSRPOaW+hbtOQ6yDN0PWxUU/EGEKOESKN45M2+c
Qk7yTuQnnIetkcdCbI2sg9u+HUIvTbPzTk3oLCczDGdkehTXNcDcVuZALbQAJTh7
Q0dOvNQD2fJoz/vP682RPsCJbWGquZmOSMkiNX/kPcavGQK81UbJIVq9tLlkPHae
qx8NZTXQja7y7JGe2jNdHkJcbYv7dEq30p0Hey1f65rqSw4jckf1N2Gh/mgEtD/I
e1iJ6zl8EUNroMIpm6jHIN95G6abe/PVBhveDgLnNuCxKDT4H9aa4BzzRel8qjjY
OBAB5YP7UnnAb6z8swDUAbU+iHu15F/toAim/xHlm5Pi9cOl3TYkjsdjNezxbc20
kwwEWHVhQ6Oudzp4y+s33JooqHh67p1yPKwqTVrzkjiKUGrVL6MS2szom6OVDCuh
t/AlN+Ha4/JwOH7OmLNonmez54TzImq65ciFmkurr21z1zYZfNr5uPe1eCWyYlPD
sibRNJUeTOLNuiYHOxhdfZECarspJiB6uE4z2LhvsxkV6r2fZA6YnNdql6a8EjkZ
dl6Jb3vp+eklu2QgF2oYP56X9rG1AQurl8C3jUw5fvACaYBBpkYWanu2SRBWetaP
Lm3fV0WKwwnZ4D5qofdqAAu5X0ecRoQg5Q2q2RBEp3lrggAs3RRtBFJQuQJFBSHk
bqGX0IToHgF7P+yVvAc8POgH2/QUarlJCNfY8nqcfN3o5Z9WN72a1q/QBZBydgKk
aPRD3I6j1w1Nz1Wj8i/eh7enMcABFxs/DkNSP710nwE/CdneYyX4bpDxcMkqFTto
Rn3hl6/LIhhPPcSuj9eXqt6higYBPaMHSM41t1hbavkFQAvNkhKZ3pXg8jeX4JmH
WoX0u8J7ssMbiw3s29HOj8P2JDbZK0wLeRcIzTG+BdywrGIuJQw3A0LhkQb2PhwL
lOulTs1tdmo3/ZVbXHVFp7Oz8iaKqVa5t1dDzZv8sFPnVFrOpliL24oDhjKZcxxL
SvDSPCV6pKQMdnVM+SaEKW+Nx1Yhoq+axlHkPK86+qZDdeh/BjEBKsGHHQ5Hu4SW
773+6NrkIkFAQSqd+skT9YjyME4XJv1JjTjSyW3Up5YM9L2RBoO0WX2WnfWn7pet
8ZC5PeYlGVU5qPfkkZt5OfNNM+wIzU9J/pqx09CaN5z6vjXBAB3YrHrmxUl4QcnK
KlAE//zX0nC7Mn2syyaIu7+1jfSqa60vddytg9v6bzQwMxX6map8tE2xuOaadDaL
hb8rH6Huzo4rKLzco5aTMgwQ8BaThjqe9Cr40ZCfG/Mk92mi7A55+Rp5S3WSLC5t
PwRkdIMUcJN8LtDDJ248PxaNWTK2aEumhSa8tW0UyXiUezOq2pzlK059GfAsOWiQ
kme47/qPj0D93JOf6oz9eKYvyOso4nvg6pidQQLD4TP8N0xT5w9abBKSmGDPE4C+
FjPF59ktOtKKq+vYg95vjlDCJeaToJh/B8/oGr2SC4d6GjfruYzmvfjzwvX05vgZ
m2tCsA5ZrISK4zYQvoH5KWsIXddksGkQj540DeiCcKf3vKr3z0J6jaXcdcmmfFCD
1eU1EQ4jVz2IWEx0XdbwN8qmmuaLchdRXWoO3+DQHBWHh5D3zIR3TbiRi8u4vsPs
4ywYdKgV6hkXurkoThDdkRvNE9x8gGcBBIjWGl9d0b6uOz+jFFEudzA3we0raa9d
cSbIF78u3Gk+LEglhvdFXZB58knYqC7l1i3vDXpl/wzz42irWY0Pv1BWkvzZkEdA
ygAB5u4F+WbLof8MOyLglho2hqGwAKQov6hQqUJWTiOK2T+yX9Vn+oDnj2Gg6Onn
7o1ybMd+FY2JlauQMJ/wWmQ57WYZwAb+ykk5zJEcabfSVP/qmn7tztpQGQwpXH8T
IoMqsm6+6QzdkguZndMHR6EmE9r3F6OaFbmYGjsNvZ+B/TCzyc+c+bba3NqpMYmD
078hHcHwsj6E45Eg6DPLLlZ0MEgH4kJUCrf58k6oc1+wvygy0hacNOZFrub39W7Y
fJF6lDQrj9fK+rSHhoqj0Zn9vslnjLv4dt+B7PKf29VDICvrRgIM1/AOzg8E/lMr
Z8nsT+EpIbqDMVTkkqyjZKlZGDgwD5YeFbbsuasM48j3yG52m+BYCzTyWpQUOWTi
PjCk2umwGphKCHzZs+X03EfAJ1FVxCwYx/3kjRS1FT54oCVzzghETWzmHE1xnD3t
+Ojk5lAVGBf6s6xoOLmPCxBJWs+WCQ30kTVZVSlAi094pP42LfVxkIdXgYnEzOhC
Uw0CgM2fRAaoVZ5ZqMy6M1SxnjfxMKmp8E1i1g50PZpTLBySTnTbZFhnrM7AlMri
knrw3rmNUtaChEHZwaRU26rnpCn0ppmYy9tsDPFcqxShFB88UpwNLLZIUoJeR+rT
KghEwcIR0u2ivZKMTenwBIsbqCDWnSJ1cGhMD6bphexSdG3WXlDw7GQrOE9nNXjK
OfIsWLDLom8vD2w73J8mqmBV9tiJcRq0n17/Wwrw6Sicm6AcwumPwXDezbYOGAYD
lDyTEb9eDPev3RRw+WtvxElTqjWjvzbgU+dJdJ0UeKru+gYWvB02RsC50HGdVOos
3DRBdLuK69tQEKQmt+GypTp3B30tAvrIswcrUMkqMTRC614reDKuADUBqkufiCyw
0ixoL8D/CncFIKHZ8FDPQR7XfAVNVm7MGOg72PLmAkPsy4TC/HyAySfAqdh915pR
zzOqkCN5kWkjt/BogO5ISXEAQcbtoI5nUqAL7wzP4ey1PdiAA3Xy/AS9kUjJLEJi
kABty174c+5DlqWvrKYgV9USCdkgwK4eiU/wCnC5XUZWksxLOrMYK1Vr86e9Sriw
tJRBQjJCERNzEuaJme0J+twPXymZ+uhR851r3wbUSeJd0BOetkxPqLcR6/c1q9ha
379Ag1AC2rQgNh6qtZ8VdzQGboomY3i7LobppNI++AAFnqr66zKgpvk1OOH7eju4
jb+T4zZMcuVdTGzjIKJVEJ8mj0U+9J5RNdHSbaE5XREWzw2XrZKT3Mxl0nKXxVQg
XRs4adYGawhn5pzpfo4hWU4/iQQcZGKx6aQzg36FjOFdRt7JCmeN47RdIP4I4J/p
r1WswQdkTX/xu+0lViJnyM52lQSOKcvtPvQ+OlIYEp6aU5XOEVDWHn/oo8Nr8vNE
zdG4628rX2is2EevBOU4P0VeKbUMFq4SkwUYcDLIeyk59LkhrJgje1bSDvOKTPkX
1Zz+NyZ9a4ox5htmtPcRx9+QhAZ6QY/fBHqdQE7f0pJYpp4EoNMU2jytwvZKIPVH
8S1f08P7JFtHVGP5NgUWgyO7shEXPBhR+DL/vpsQaxaViKQE6ZtYGzCfasPM0q0r
yTml7J3s6rNd3UQZ9tJdE/Qjk8PEZf2QpISYLlZ2SPRWIOUjZQXRwmV53WkhzwXJ
2sikJOeZ/u7U0KASVeOPalH86w5BP8IgEOUUpfWIpqaPrKEJZveQtuN/an+NlFDA
P6THOt4xLdVGS3Y9URKN3PelFaguys5t9mCwS5MDcX2mFW1dtjTOmXPnrU8/vPhF
GdJgMYilGFGyZMF9D17dLHhOMZJjRd+YvxAdG8+tD2APflQAuSyOz7tgw4P9arAw
KeQqMhh7higk1XcEfZJflXZBWA1PFMxdCBn06VDEn4hqfmPuJ5JLIr+cC3JkBsx7
1nPA44bl0ygOA/8ALlSTIUbHcs89iZ75zXgCHETq0ZzorBhzmO4WiSECDAkqowZa
tjeg6fNxNm32eiG7Hm2KUoyF2VjX8CZHLEMz4YBrS7G4F5A6IsdjWFqREXP5PE1e
EiflRgg3trcdyf9bIS8J0qGCs5cGwb/BH+cREb+mP4VMAqc4FZhNORBQqzL0WcBd
sw7IfVZqalTBBDmn1RourRAOYvYW+rElnI+BTivp7ZAXeJcaS4wDRx+CW4Q4/jEM
CvU+EF080Mb5tBPcSBLauMsGdPFuZpKjTXavzZwUaXlxFGwCocuh6Zn1TMsq4H9N
McrORqm71fBxOSPjHfceKUeyJ9KYQLW37GAoAPEtaleqoOrqPXzaT2pLSrV1tRuB
GShnbYrXlCmwqT4PNpnfB1GZmW7keJMzBTp4t4HjrVxiKFZS9i8NOQJ+QPfZx7hn
bnKKBA6rtcZX1wY5UpoUV3dvmMCpacuIBBaiETRvFJjlqMGz32qBBc7iS3iyTRha
Ge6AtU9UFJYQhvRYVbDfgMNX9bnFRndrTHAuVym65NTVYl97X6clz4iqKoUebbp9
VCYYkggwpyfWez5g/Bn3R/lXH7QR+Xn333dUk3FbQc56ytJPp9GiIhjbpQRgS7CW
31gy5JgCe2lurdUxdxameymEzbRqyUnrho3KGGFtcTLh0mYG/EFCjOTGh4FLFbO1
G1l4aIaFoYfrAasAABkSIPPbrqPLZk8p/9YScmm7/S1gDzyyp/haDpea3tdoix9e
oo+6a/QmfmO5/HTHYa4o+r7Xl/Zl7l6dxxz9M/giqNaJhJK4NVO1AcN9BEwkOj2r
0bsLzDqHIyam3B50IkJD1nPv6rPtV89NfwKLYduqMSQRLr4O14h8/bDEcTDy5zqS
usb9IGUFI96RPPnJGqBdHWILOj7Pd4nVg194EP0bN/+fowFjuhD/E3O3RoEelYcE
SqDPJWhAuOyC12o/0I3/sWNluI5k0cr8yj1xCANsmiCbJ0AVYxAu1uDWbFY5QbDo
MuvkZMHSgXhQggjTugktfqp3T8TDFp9V+hzNep9kyiKSQ6F/lxQjMBgJqTWHihQn
nu7AXHtEozeng6VQQ0aOtRf54EvNJtelb8/MH/17camuVJ60JAsUO6bba+9kwxvP
RwrJcQhUWT6sD2g/sDYw5hoW0r8xZhVXfkdimgUKazqFbwvdbZw/uOOb40i1AvK6
HWP5mSAPV3eZnTDFKNQvmYU0dvILxokfSq3T0Sk1gzaNOpftRovFYfb3GH7WewAu
NuWBXYCL1YjGO2vWGqS1njornw6MhTrT4SmWEN2eXZIPUO5pWFT/GsDlWa7FB5HV
6nhJpDDFSDPtiBCWx7i1e75tegHtLHL8lxa3/MMAULbBQdfyN3EPsE/HMce7QjRA
LTHHgNrWTbsxFq/VMUIFabBkm94uCIHDJU5v3T0nRlpDrcuzDG3Z0HA2IFtMvQG7
QmOHrhehhbN19GmCHMBvu3/alMsdbLWvRxtGlx8JEtoKn8fz9bIBIil2eOw2+Q3d
eHIxtsnDg/XbT3HTa9oXN6sS7N/631geJcqUTOYxbgF35fYYhCiTv4sYvHh1kBTE
lI/FIuDxC0886Jyzvxd0WQRWWT35O8F5bUTWg6jbezLmqNmhr72c9hpT2PmDyqtk
Zs2VH62m42auLktXB7pXBnGpLpFdSMRh6O1dx+JWu1+H7HQ5tPDczWfY+20cbJHt
WbZ9IHhDztMB4lufF+zq3DnIBXgvbnwOfJtqH31mmRzoF0hjiQhhmjRIVh90I2LP
NTkqR5Q7oBw8N8Bad54/dbddyhEVBoYR/O/zl1B3yRBUR/8wfT74pPD/FNjKRvRg
Lk6VcmFUSGJsWOL1MQ6nCqehOZNb1p4AlIhe4gGUP1TBJasrGIXu7sqDFJYhlpWh
mdTILKx3l1OrqvzK/REYWhGdx2Bz49iNEZQLHccdPWNqK52d4aJXpv9FGvWb96iu
2snk0ckMdv4Rd8h4HLQLD7Q5YwQ1PXpq4GeHGExGlJUqfUI8VFWaXbmzySpRADgZ
Ahjy10EAitlGfOTNe7w98a1kveuCDOHoEVPiSQgugenWo2F/Ne4OLWN4egmfmS5n
lGmVVM5C7BNN9PhQubou1yOvUfoOKMGy1khUzFHMdTCjNP578l31qkEoQOsQk2Uc
H7tUFF4HiFVzZBY8+rAOiVnFEgm8HpEcbh5FfRlNA7jYBMr2zNp9CHHhec9kZFMn
Jj2j+3HyquvkkOgkxMAS9ukTdOLGP9GBhPCKuu4eYyG6CuygrzGQl+rSv62+BPdI
WUR1xsDVk0dk6dSLRiTdGzQ+xSymF66gUh7xceYoNG5vj7f8moyWDOqMMU33u9cU
Qr8M0quRyuQYPQ3ekt2cdWRGb/AktaKvJTIBKTRt0br6aesdXM/VgoVlZoReOQkz
3F+e+bsoaf/u+CdVrVgFBIaOmZTEXZbG3mGpC422aT9YJEVUulto2j5u3v2LyxoP
jCkS6LRDCZRki1AKMzu2NLg0yGCeOyBa5nQC0XM0tsFMW6veKLBx3+l/CinblxkU
P9aCRdpxocm3GHTd/Otsec6062MMZ7rGlKLHodGlaroIb5p6PW6l139yxG5WXaf9
4T54DOteoxe5BeqfqBLN8uSy38hcjkkEBhPfLyWlXhc2wbt+XjMZaCn+tKGNlBVG
TLLkc9mKZwvpjnXvx+ANhQbKvG8QZ3IhNj7XDn2v8iudKq6N0CBhFmPSBE40sNh6
zyaf+hs87BHHuLyOVY0+SBCdYgH5d1qsfoBpATzuRBz8bL+cDkWh6LsGFy7xALdC
AMoo+DQTpqwbjSyt0zaH9zsw536jqXr1hSNk7+FHAYUfczyAycIoEEG3xoab45PT
DNnEvRIhD0J36pf/AnDfp8upiQMjLUT+V/LfCcJX8kG5DraIbjfdPObgeZNYtWFE
fh88fziAhz00Mlfy6UnoQpMGNhnCWI2j1zS/k0ixmq6JjKWSQExdrIulh+RpSgdV
yz5jWm647GHCMivPVT2ofGtk71v04yyTjhpZWFxHvQieMLeFCz3frdowXnZe6Bwx
nHf4aFAOoYv6F366LM9E+mK5ife6QYgIzPIJPjJ/CpwqwWNBo5vqrq1tdrdd8x5o
3Sy22nRH9GWfB5s/KjTtL2qhGkjvi6LhKYJ9aftW5/ZqMAMEU05Sfe/JAEGPoDXL
0rEi/oH+u380nteQHhiOvbbBjaWahgauu7o2//+QbKchGmKv5z0P4UseduVShkkr
xBHpd4fuU0GsTOBFljUJ+64FvN22qFCSVh7zmi3+FPAUQR1y3M/9XE8x8Ye0IF21
136g+BdlpxIcJYEVK/kzasxFC7gW2IZXu46eUEoe5CAo/u5eKlTCBRhWi0oF03W1
TqmTEe0Vx0WqcPfystXFCdKO1VzpMju0nRn7klyKwU5enw5u2aStuvTWjKeJgpph
3STgUmPDHUYftxRe2LeuS9HFIcxjjig1JunaYVsigjdfYlEcoLxpddq0HKr1tP1x
uK6ub1KTp5rpzyqyVFhdfsL+CUubzDPRjjj8ZvwgBZHSaVWsi79uxg1cC355EFgw
W4fWPzLvFZGUZ7HttdxbvX3d3DE0dYEQ0q5X/xMuoIE8N82HWrBTpNFlM9X08VCO
XcRiG4CJvzI+dM6LQnLqpA7XfmlGQmww6vsNbZizJGPKyUEabOx+9GvYuXnc6l6t
2C2iETjMG2Kp7CMc8DR0mJLzDXPvz9YZd9I+aeUTwh3OtPl5PorGinn5vf8MEJZr
a25XaPXdLcQU5DZieGIt2IXFzBMqQoBFatPtjftog7GkBEQ2Kr3N4iRTYrrCVAeY
wXLHAZJFRs4W8pQEhdoaNYigZcxydLFBp1iV6oGvTHl0bD3b4ouTpcAFHNtEoEqw
dZlt2kq60WsjXMV73DUbhRe8NYThIf7IBPL8EsD0qNacHmjcocV4egOKDEXvS3OG
mdYZ0X0RB9u4PvqvBWcVGw5kLsP7UXAGe/oepBD18W7LuaKOFrCrSOSUKIAqcpAd
EUBIqSvDDZMYAnQSP7b/4XzZnD3LBXNP7vukfU8jz3NYMJy3uDdQu7ceaAKDah4L
I6LdgKOJUW4fPoqjdP8PeVYJwzHGNlmQ4mWOFE5Qn00ZVXAuM00ziumupnSSkk/D
Yw435kQS3YgqTU8J9qMju2nBBwqalP1K9xrjikY69mcasCrG3k2lLeTVJMchCe0r
f4pqxDDiegI3yh9xacImbuIwYNfpKc/GaBS1NSr7gZZ21lwiOFAslfXjJoQ7coF/
49wFmXK8WvyeRDEsh7Wf7VlBbDadScDWkkMg26Pte82Ebe+uk3BgpJRUuDWOhPNr
nLg/LdAih5MJ2pCJhj3SlchmWnodxIegou46rM/YvUJEQkhtvaL5UMkCHcUvfVUX
/sla+vgRt9pwRSKlc61CBUjQ1plLbPrO0XBCSB6mo1V3seu5eH7sPu/jLwDjZWk4
CW39AmA8+hDIyHG5eAmIVu7aeCuRtJC5OrpbXXJI8j8ItOO6S01ckYA3Q6rKpIvF
/++0Wgk0iDiFJGxr9z69vzii51NOHHFxo4FC8nLjDM/4/n5DpULP06knuDBkK/ni
dhNR8Wt3VnQkMj0310E7fLXrBuHJ572n9Pg1112YLJeMceMoKJtqYsbKhM1mUlkw
+IhshPiFS56mPbduhIeFiAVYf/weXf8igOiLeNdO3Wfz4Lr9nISBhL6MGqClm+1l
v58kZSRUENuheisSq0/2Oiu9DIvgGNVMv7PFKjCk71dBgy2ExWvzA/B+rahBEpM0
/FnHoXa1s4udCh6OAUH15xoRcdwvIelWptbwBNVcp2AJMNaBXl/NP1hPjV/ZA2ao
ce5VFIf8oWz5VwWsW4veamZLE53AUbViNMOPtdmMb+cyzw4J+HKT9JB/d3MvLW92
Cd+CyacQERvluxCHJn9l9BSw5OO8aIUyPoqOCjvoiySJw/G9XSnjzmH0xJWChLMP
zhOA0JDddelVF82VtwYbrI5utUvfkHZPGI2DogmzD34mlpkYOMz7SIxYKvowYAhl
GDn1g75ey4MVBRCRUpFoiq8WCFmolK0mWkaoRoeCr7w8iYVdXTIiVEr5qCoC+WC4
vLgSCn3olcP/72oYzggsLf8wTytu7VcPEmP8UdVtLObSoSwAsrMU0E8poCtpBkgl
1gYwPSknRe1CRZUb48mGAQy8SG1qdJB+gMNkXoFiWCMw7eaTGHF6j3l3S6rWyP9d
wIJYVCAGwU5mPZ57OqPay+IjZEFKbG1QCDjhxUxbtqp18SewnjgsiIoKD4vcXac2
5zu/a24015By/ev2+gt19cAhwPpwd2Eg7YIKq10iqMBY4LUAwOMSsNoTOElAQXw0
oAseFTx8LAp1b4uwMyL3/w23kddnytRai5tFfaq2/vDNGLAoWtw+3TyvELeGrTZs
QKfHqyJ29ffBYNC+TXr23VEYyD3fLiOcBFy/Ff9AgEZaNju5511JGLjbENbvMSvD
wncWgwidxYUSlxLuh6SuGdUZbZO2i5wtWlYUs2w6inJQXxpQ1smfooVWV2Ch2rFf
Vm0G7y7RaNibLfQjd5yX6497gJ0eLp0mUAPuyOP4oCK9zcWSGRBE2UwU+KzYPxXz
t1PI44WtFZGDYOBPCIrBx7oPQJezXAPYk0JmNlfCBYhRrno9AWrUZuYgrN2npKVG
E41XE4xC8gF37iKz1FTACewgz+gXQpmMHvIwWeitPtQRyleNJhbxUP8NpipwrIbE
G+1IGfWqTUevrIqwF+D7y0R4uDiMgFU03+RfZXoFlRfwF0RDi38+qpwP0HrC6rQm
egc8xwoj6dWPwdCIEORAhKMDOW8+qi0PqDnWbuRYGLi6eOoyiSgoTIFBhmcj2kpz
ASDAcH5oSAJVV+5yD1Jo5KXtGkE1uej+B9NYu8vCun/raRNqkkJ4wG+zNlMKkLRM
qmK3xx6ZHLSSFA0IHPTuE9Qntn/AgKLr87SdYDh1O1ePFFVgsBiJJTK98YBcWNz7
WQXaHB73uWQoJrsJ5gjuSO6UYlNnLwnknhVs8VNCwl5jKWHdaSuuc0xIz3kN0/Cn
U6Ws7x11k2g8Ai0ebwjA+s40vIaw3VjE4IdI0W7W8NwCdMjlLzFhN2Q/xjURA1vP
jrtblZqrOC0x5lkOyZCHv/Jl7xUMXe7lyi8EowKqudhI4VF2pmpNIVmKzdjk0OEN
th348b1Ve5dhsQc+Y41M6AcpPpZgUJawzHmD/wfjFa8hDOvqna1DOnC/N8DXQwXo
oEjTLKVxPSF2+u2pKWX8NNE7QEfDPwC/6501tEq7T+OY5wmTMmqjXXB0p+Z53M4B
u1pgwlVVus5Fc9iv1zkR3dHVRXHeRVBV0jzzzJqWvWcOMEaisJBBAEuJ3gZHK26Y
njmq0RL1cEBSlpcpzgU3Bcapqvj64v+jPWg1t56ZXyenTVrKMqHb88wb10G0T3o+
dNqKJLk/abYyNaOGIgGlRxha+AJ/o07g8lsC3sxxDW1sy8VBl0hnVIhUpltU4bmP
QW+03Bu5Kr6xSmEY5stSF93Uqp4I1v0as3blG3x00xIQLsw1xneFyc/5GnDXQ40v
SIv0WGKGIXnGR27MKCGJGSNm1uoDPg+bnTmfl7wlL9ceeaAe/g4WTGBh2D11YuUW
UwO7O25HXKIWXm9ZdXir2pJgJmJAaus8RFqzVxo5n+LkRAHr6k/rkmxdZvWCs6bR
0Yuj9iCJhKm1f8jtLw3JTFC2di/4Az0eaP29EvAxUqk650IEy/CGrF9M37vDW6OG
qJipkxxHyaGpp5A+7s6k9Aqs1os0Iv5M0ijFvMD3Z1WDtcSKNy7r6j8RBDSkBmyf
P7+GlrS/pPb9YCv5O1ppAzTmGmrfvxcDJr7QjMKiXAeGipc8scbVryY0sys9yyFU
Xu5p4UyRJ9ld71ZTQhpl7IDZTDB1MNgPPGw3AnLZAJ8CVeQCQhgQg9W3sr7TBfSf
xzW4z6a9mvbVhK+92IFriQLj5RAa0GAqb6BbSS5qCN32sWIgJ01WvAvldP5ZqHR4
DT4L1u8G/QmNLZx3aksgC2cMHmCBQ0fmTtyH/J12+ki0BV+78zbe69TK4iEdVhSS
BTezSR1liCYnGVsXJK6ttLB1CqJQJLtaSNLB2ienXuJ5SgDn61WAv/tEAQ7er0xx
1XjXQDDd50DzxMSY5ZoPDxVn0+69fgpq3bBvFzalu7u5vXFeYuXgAFwj8SqHIYwU
9nIvJobBunvHmhSMJR14lUSaGaEpndJVg6dCMOpQTnhCfFIs8vt8u6/8BV2AlC7o
DK++CQMEIBEWit6AewsFFUtFD+ZL1JDEsSBFARxDHVeM6YC9Q8HoD4rvnVPi5u9B
+nmksmiydFojV4PpUTvTlMF5qTBApCdwifg8w9hCVC3GSmJaQs9BxepOv6Wu+771
f95hyjtA7sMGK5kRXLeg1VKja+EK9XMqwUpnemoRn4+ZZ1IyK+J4xr2O3tUxdcHp
bQl/fDtaXvc5Zo+5xLhnbEehrm+afQSDSkM/nPAANjcy6+QK3xt+CeTZlWzjkWod
6u3AAkVC33In+PUIPSh6nD9u/YmD2coAX5UyUQm+kSkOWnaC4lBTFoOfi2JIqXQy
Dt3DPrwu7iozCUngq0zMvfw4giBBi9GHgGv0MUc4cLJlQyH2/JBgKdns10pRYVYv
/iNsw6WjJ2djtvZzOMCbYFHn9WPygCnHlGicWF6Cc28TEoCmR2k6cnIdCt+4qBLh
6UKeO/HwGjfphRlAOqBPWfWYGwSwpNgOwdHMTNikH6s9xp7yuRATzNt6U26eVbgT
+a/RrOHxyuAUK/FrUc0HDibBw2FvTIG+kg4aPY8cOwP5iqyc5NAakZMtqhL3NH5l
Dc2qVognY4+VbtZ5JJ2K+p5Leov9SXRewSWGC8uJicJZT50nIlYj8mcfZnJK7jvO
oBPCbbMKgSly9pyX+tBbiFyh5KbH2b6LxIAoJriqS3aHwa8AUnjnruKNw76qZlQN
KKYkJ9v2FPBcoD9J2vMSvyO7jC4yKZX5ZsHCBgu2QT+9+daAAeMW1JBhDZQVCHns
x5BBVrMxmzr8hU5zIP8CDoTtXqH5FEBfWsfAiioipesufoG0QrV2o/YkCEFYap+r
0pRTTPdjd/pZtIUXSONZK6oB5/ZwbpoFp1u0RlrTujyUeHbDtXZr30VQr8kIHjnF
As4bNA5NhHp+H12iQBadZbHeMcGriUnr1C7N2m9R9xNR0owGLAPT0QYwY3I4/ktc
/0k5OM9zjMJb0TsMTIB/6RFAuxg6NjESBoh0Q2KT3VZdff5P8quwvgexklEbJ366
ticYN29mBO3wmyTC1c/AHBH5uUWdLljh0VVCq3jOlS1IZ3JKeZ4Om2pxW2dQFgg0
8p1StgW5f9yghlOtjAY0mFoW7yBfULhtOT2z5KLWVdY2OXJBkcKIzjbTRWVxBSQO
FO7p3B4NAhPWCFii24/+v5BxbLthA+Px8U5RwLxlTqBVRbVAnwEf1KRdvhFXOG7T
7GK2zA5AUYFRGoD4r3J0YZd/zm6JSZ9OM+6mHjwqOnRwEG+/tfe/TeRi0TNnQ8Ut
/FYGb+uB+A2JPiMzlGBdIT/t74WDD9Ucy2l/l68AzlgG0nvPrVh0GgJh6aeD/n5y
Bg+5ufqzsYitqoyCbuRTt+orAUQ7IB2/3L0IJl6jib6p+7ebnGxoxLOUWO8zSweY
QOTs8cRSnPx/DPrcnAmu34R43hWIPPvwU2LELY0PSvuUdKQG5z0w2egQRok5fQNL
jmokWTGa8fDzt8BxrGFQws+3gcCKpVBMw1QlC2i2ypYClwALw2OvaFJ3rNOZ/uqJ
BS9NGaR7dqb+tjDmJq/0XaHKEPobaskiccPp+x6L01HzozUHI6rsqnvAAE1TGamk
Xk3VMiqBLFD9UueJxyGvqyxpy4EjeV23Xws18ucPUfv02w9F9rDJyz6ZS7Fu9w6i
/8VHevtpdYF6ttY0GafiVeX6B9C0oReev8Lz6P/QMv6d9yXCJrkD69bjqIEuqkV8
SYyq3iepAr0KXaFBwW0082fhrK4srfZwM0oT+v9XlCNKPQxn1RGpY0F8J956U0Rl
OWuDasLuUnsQ25vMfq12qS1BojJwek9Ajdft/CcP5Vp458uiUfheD8XJmi+8WV4b
aE6Z/Q/QAYJPFf+oczKC90B/nTfgs7z/F25LCC3JqT2UiJ7dg7uy4oBIi+Cl4k72
LZpKOIiNdr/AX3988YrHZWX9T6+rLVPHG+Z4yontNMhfpZ8xKgBfZQT4+en4JXdz
l6KXmhmd1MSbwWcrxTPUX3WzUNo+uYLXucmHYz4GvSFVLSPqt5Gt1s5H13/Yil7l
AvC6vh/qw6obeiZ+R8vanfhCF2SAvUmpbjXGBXCxHBTDpXkzW1Juud3u8P7sEw/W
chBjdmNnXSHqZdiptdD4SmkcGM38jkHdn50i8AGexT9X7Ov93tEdEjU8NLA6Fhkn
7MKRIjIbVZULcA1mT/q5ZjD4a8mYCibZpQVWyqZbxrFy+XVfmbNlKX1MXjz/SoEG
d3jamphe657ImOIK7LY4osvzScUn22sSbMdkm9WycwRrHlIf3CyiW/ZGMVVNC5Sf
xP9n+EwWKlHnQ4vcZf1KXLhNoFiXNE0OUK+DTdeHYUmZVijsWXqS6s+Pjmoo873e
+YwZ0aZc8w8K3jsGUo+NIC52N/jfDR22F6AkvUeIerFs7ocZyS9TgZbdDeuUkKgB
/fSpGGrTkyCXTC/Ny94bNTKXJe+dxfOUUM5M+fqiEqMgj0T/WeHI0ys3aulO7suO
i89SHxvp23ZyNcMyqBZxdac2v+MXi0RxxMz5INBphpTQ0rsjjsvsDamEpp7qBXhE
McPLRwNHnJMMhbfsLhaYo8i0OltxqD+vpNPcehnp1K1bHtiWVTS9m48Kb2vqZNoe
sqry3QD0JhyTDeXr4kK4f7VsNxn8BLWbUSrUGMCrxLVI/6PzFnYRN9cZHimPZTN+
RbuMVpTXufuU94ABOfTgGMt1FneFiXEkJdFcXCZZcgzxWGH3EyYxbUXM7Lfr6QGK
Q6WUP62L241Pi6EvEjswH93doFQfouQJo+SlHsxaG5l8rr/LsDcigtxq76VTkQpw
vf5wZmAaZqlxIpzvCiT93x+S4wAPxQZ+V2lAbNQOCMiU33mliSQuaUFGp/Eekz7Y
ZpED726sduBxcWQk+fYgcb7UCz3dX3sEwOo8SZhYBwNN1U82Q8q+yAMVVZ4/BjDV
ck90yVQkr+qn8TB54QXCDk39aD7LU0Sz/b+9nNoRt68CeYhHBHqIFTvFRrSvBMEO
62TXdreI7YQxn39autn68S28OZEGrgnNjtLOvQRdzNyRsCDoopnDXMOvxbpITDyu
eFjNb0s/GfQDvpXePu9fs8bTTQL0XijGuY+u8z13SmVIaEEVyWqtRlzjApDkwojG
FmMCT+wX2YicyqcKSDnlpBQxOHnkneYzzyqyrS8TFaIwh+EDgAnX6d7Tyug3+Gdp
wnu0stWTFd9hiquAvhaIByVuNn5fF32ZEQZhH1iIM3gpKcMUfMhnVMSv5ddAQym+
mC/ND1yVmEa+v53WqhjlSZmFa4WsqNqjTbL2/2ke8U8HJGFfQOnOiPOc8zdXW7Ut
nQz/D/skQOZKlD9yLIZ4lGiHMEYP8WIMRmsKkOrO815otCrkiY8p+pCywt38inG6
6Ig6r/DmePY/UQnpIpQ6cOQvtGheZViEgl98V1oL/XQZSFavtXjhSgMnB1tguTvD
OW6paUXtV6EN1I933jMSbr8MIsgVoXig8wFTJgyv6B4IYccEuoQd28zkpzpD9nDc
3NDmy5ETwqoeXi346X/Z+dohbSoQguydukPFTKgiU0AcC0G7tS1Z1s9g8qAJU8Dh
jFa6jwvMj/es+4t/Brt26V7fgnkTlJnCoomNuii4IxvIENlB5LJl+yp0+EefXyjA
H1WMzt2iTOlutITyfsiZNGPqllBkPMC7AACEPJF5h8c/i3i1wEq8t8PpYHjl1ZI6
C1pDVmQmSA9H/HZoDNr/XdZneeSm+7Ul4SYst9DnnZWexRxyBhdzkcYTleZTz94C
fwQDpfK/XzQuF7yp+Lh0hsZC9PC0DNbMMM0ZH3ik77fMvhwpZmMSBxzaeCsJBymF
o2PGPPEHwDtkVnnsJGdsdXh87gqHg15TiUEfZsszFuf9dLnU+QPgcHEVH4FHFKv8
ccKBDrJsh8iQC/yb+M5DykPGACGZ2FHEJ3PnE/dpCXeCaY0UrtxCp5bABelt9AEX
Kjsn/FbzqQ0PHNuLS19SpfPvlC13jtap+ECi/76fP0Haq/Eqesl8ThM/UAwimchq
jTV+S/ZvVOsi0uIk6ImlOZYVQGojRg/TTbUFTH5rDVviLj34YujkuyLyEA98nlFj
La9i5gp8Pkyp/yOT2c1uM4vBwTZR1GOiuoApjkmct1TMpwsVTp6DSwlZ7UxnrFM/
6Glwg+G14/4tNJdNamfdd94RaAk2aK8ocwSYquBQ28CItQq3N2z7B5W1U6YcCTqy
HXukd5iWJafCUa1LSrrNSZDQPYZtn58gVX2RsojI7+ovyJWkLhK9BR4hWmAIZvfw
bbotjV6gELOPjr+y9gOSJreR9HFuMrFIUrbDrQGhSaZId3QpG3TFw7Mbym6FNQAe
MABxxJ876P6tOOal8rRLxtOr+3j8lxCr9W7VHWy9NNs5HiZDrNf4zIqU+XCBm8BZ
PvHxjisF+oNdPnWXZknnePd7vyi4wjLamCnv3jMPNY+3gbQgsBo+G1gfiF50aB5N
MBzIkBPzbZAjRn+Y2n5G7WrqbmaHqTZtG4+TUSnE3l+3AGD3WXyJOTraciA12y4I
m6qchEbfmmfT+LfHaGao/wWHBASrKhdR05uy7MYV2P0xdbrkkOFyoP8QlnXGA8FB
KHj8rfWsj+o+te6XtvSdKDAb6yIbadCXzXydj+gbSE/5qyFcrFUsOjoDEwQucZ4v
lt6OI7qjCiPBhWhydNuNHTFvDf3IyCeghma/1eJtBEHdXb96QARCE/CKgvDL5iWQ
u/9jq42l3cApYIgDvuEHDnkRTZNHqDJSLN+qNwyXAx6ZvQj5ti72iNx0aAJs5djy
LRXwELPlaKMJZKz51NOytawJXRPbrxQPdKCEiYrjZd+J4e/538nOVzgyTifIX3/Y
OOy0TG0T4pCgPW0snA5vVEW/tcEwVkuEwIVtpLfbdAo9Y+bb2SNFlwCqnbQujbIQ
RGeAJJ6+pZ8Vgn/q1B3GI6SPNMUFVC0ea8BQUy55ncwhjMZ4xiOMka9U+rtT5CtZ
7O1HFGWgp0A6+HidxeVNf1C2pi7P6GrDG4aEfPEplB8NrwmDApH9enyW6HSK2EjM
Owwwkq0qwRJu9myLHGHOQSZyllVcKY1jQwHS+H6jqN+O0GFM7Zx4mX1mLFOYPtYW
/7AmhFnWZoY7FjUb6AD5dy0UxixVqcpE5466kSno5O9qCirwF/ZpK/uEP6mWfKyw
chVNIiZjTpibGd1tEnxEjrHvIQIIr21ydtYuURYftB/FFyOFY6BBMs7AjERGhD1N
i9bLTJ3Q/RmDM3zHum/SHPGubixBI3w1kxikDdN9Phak7NF0B7lClwqnToiNodD+
UD6Ed3uUxE9qAyWp3glecFYJ3OnPKatQ3CnSajjEdL6bsC1XJUGeI9BkwLLebZz1
lq9DwNLqzJXC9hI7Lxua1xZj/OoeZapZC3fOCUNrLKKrFd4dYqdZbMBBN2aV2rwY
yDOFWCq3yNKZ/0mEqza/6Lje7nxHaOFoOD7dhwhbTYmzwAsWEqrSxDyswiVfpIOu
UbaGKYjTQ1TPeJ9AvUehOTZwNay2GpaTPHNZpSR+iQqPEG90j8zqteLVbQjVVnpE
YHfw8ye1481f3Vl40TGGxmLSzlFkoiXMeAqjY5jYAyxXhpdC4ZMvrCTg/B1D4/sH
YrpYgga3Wqp65mbrgRjxjdhncTh6JHl1HIfVp+4u7EjQI/MLtlrwUfsWACsMutDz
InTCA3IxC+FPsx8m/Hu/StbHa3Tp3GmEbMzjw/V0AAL8B3BU2mn6LRuLg2d98ib0
/x847Ft8cIFMazVGtkDDJ01s/EHKGTl6ktgLtiY9oxqESw8kM/dN9t/ZUONE70+4
+0tEEFwRe/dQUaGk1ItySme0FK0pQ6kRCxmmEbOJbKKS0vFey/U86J6zCRon97s1
VIzhTZW9c32LWYwZTh0ic0kWH4AaAQaSGATps3OhHPWtDSAl3SGvwg5ACIceTNpO
FwhEokeNdHFUa4tFZcv/dOl0FzZAanMqpGddVckla9hzC9v2LEMxQ4Iv5LgSD4W6
vcr3LyT7unmIFFkkR3IoUIFf93tWH+ExSXjxhEcc+5IHXffmsAPOOuMSnJOzy0eK
Ps/+SrzxZIMfbnbEL86kPbTS2rEhOf+fkhYaJ58b2dEJIF8DjTEowoAX8neI2JE5
VhM4eOg+fszMyt9bYdEGoTkHQiVppVZ2pj1ZNJu8U2Fj9KAEr4ifR7B0fcRR9H9u
UtkrGZEGOnSyDWDRc8MWosbqf9wLnMNBNT5Rm4DJRYmpnl2S0x9irSpeKPEG2BUi
m2g/iyGtf0yde3WkonttEHsYNMWg2H2o/Jf2Liw4yMjXUlmQ8CUiIah9MagNWn0D
4iSSoR8r0UtncaFmdIAXZDdo6vYuYLfmXean+F64WegexLvtKKqGlu++ft8Zjt97
xurl0ohlnciQWkDqo8Uud/1YcurpvgRcFdad7QFc4k2563Tr53J78Ktht/+R7hTn
V3xXrfHHaC/h0GaVt+GjbD4QWmc1kDd8/qMYdPqqevwbacOyvgpY+5m4I58e02zZ
fknKqr8M4CRE5ZAzrzJIkoPy+dN4+LI/9kCFuAiqbMZegtYudWrePJX2EFpwmhI4
/15CTRyr2Wp+LND/Ubgn/mndtd8lde/6n1f3z5zZPI2xvm2tzhyuFEbaXVAQ2cu5
sbX4/cmSgfKzCXolUHGmAQvZ4oRaJMrvD/KDTw+GF/BG8Fc2cWRQzXHGId5RkDxk
YF4Bt74M26sfGjlKiwC0ATkueQRjWlS3sOxEY7VlYOF+4jgRTiyHk4w/S4g+w0VC
u3ZuezyBxlRNAWG7w8uLW3EjGK16kfh47Gwy7MHDAmXJSKrbTJB2qRHby6nwi282
iIGVxM80Aag3Gr2iic37yqCGotDQygZqY9KDKv64PH0p3XWWrbBTRyuVmU/EsE8A
V7C33t+XYkca0ewGD2u8Wucl67uLJzTmPEJuAREltb0CTMZKUPUqsnP1T4Lfl45S
1kATws7gzZWu3hgO6GbC9S7NqJCZZqDzyCCHBAhBLqmZLA28qcI5pZIkPuI7orZJ
LPflk/X4VK2phvn97mWttenSuHgBFs0MnGcV0jF8f+dhMd8bfxBNSY25fqZFjLIO
MeIclZgxD1tIEvnlQrHS6MQrr5xjAcwPEyS/l1VvOlO/GNspjvTZ+kw3IQWWs3lU
+NfiDAiNpYEIcz62qCIf1rEpsy6cUytbN70GJkOZuZqmAxO6S+gwln26kQHT+cNt
Wx6wZOt82fnDHuteCiYJBUdHgIAu3B+AAws+ktbpnG4v7+FFDeRwNXYyda/BTIZt
vREosLWMzB5lTEa0VRf7Bvl5MZAyPdGRrO+RmlaanTo8hhTJsGB/zpHPuQ5vN6Ie
hBmT8g+V8OPpl+yVpgwqNSnDdh+t04dhMF9jVSdJpUKHl4yFAtGopJDoC1RA6p5R
WAGu7nZGLUa1sujKteEYd07zRC3Fdi2vVWL/L6JEtOoJOs14cNHxyLQAsa9DgKzs
LhssOCTEXPKNUI0ZGG7NAMEDeiHQiwv8X+MwKjv8lgD+oO23GQ+RxuLB9VQn+CfD
I49fv5ywEvob6V1J71dSdfnjIuweXYWepJw3KlsuoIqmojqfeVdjCHmZB9NgdSRY
t4b+qGdGKbNC+AH2B3AVdNfjt+5ZALjvE7nweWOve2N+JV13Q0o+pSxF0eVid/ly
V2bNlWhL4qF7r81VlezJFBmTAa22yvMVtfVBnAtVouKi0ZtwI6R3HFssMwgiCYjs
KJFTKrvJfNJTmwteLF4szYbdTytvFQeyw1uQHGt64ws+kdzbTZPKii5K4aly0N5p
YaTzPL+rW6CjK7uU37+I5m46ktiChkpNOQz1lIs2DhmOo8714ASKWKLnUKYFt6Om
KYA6hDxtUiGDwhLxItDS/KlUTkx3UPlADmqQsRcR1SmH/DGhST8lst9Qkekrckga
Ir84ga1L9+dvG3/drEcXD+/cksHV5JhGM0gROmeOU2q0ah2vlEkbbA1TJzcW2Mik
1rL0dqstIa2XTrVGAgercqircrUOMiuSfZ6kmeeoFNTI2GdIzOVZ3QHrEvovdpdG
uoWvOm2UQsaDxTiOhz3GAaqHa3MeSrDGV1A7wRXvzRSYYEhu6tG9TJE79Vz1XEFe
b1wxvarH18SkSJCMwCz/VVfSFgFU+xwnSQv4FRQrXiQWuQ4ciu05V0y31L1iffEQ
FoiOe+z8N8TCmghDx9w0YEBYj/Fl2RnFhP9w2hot0FSIwArj25mqMvSUngnFo81Z
HGZjzhJficQWkDtIhFz0sqJ+rJEoJ/S10cPrqDoN07csucw7P4IydEEsGLbF9Ivx
3xR3djid8qyBNUqDIymOmdwkxm8hGpXmQjdaTjKCzLr8p7U0dWvJ1W0Y9d0tnZl1
0KIhE0TK4bO9yZYnXdV9rQ3WGFi9wnLQrxW0FI5NIDcFNyWVCNB//TPvj0ng7MNe
jFP+BCOOflUbiSSwiZAEGhRAlVb5VmAlxSr2mn0cCSCNWDUuEaMcclB5l5VX3w2b
WLvGqxLo6YLex2n6iBOQ0sw/YPDIxR3hfrevx8wv+4oBAnxjifXGzVx6USc9uxP6
n0np7LXAnhrfwuhhBMMuysdNSttyF9T4YVUgjTX6XcUk6365Ha8zJBj9nHJthq+b
FHqoPqj6gLNiOgu0aPfJvcufNhibtkIRMk/shkNCto6K2SgKcJjDXy8/Lz+X2/Z5
q76xVvgV6U34yTD4azwC3bjgT9EjgtkL7sJwv00i3y5oUmjryqEcVkdQf+f9nNyO
NAhsgrhgVsbOqeH6GhR824xF2wjB6bHm/iiLVDpItmX+VmNF20jtEONy2URu9ohA
UG4IztsLbIyKga0HRUbp6pM+A+uqeMA48pzubgrGmLG7KM2U13bzEkPM8ET0WRMT
vCnMKumq2XnG5QSu9ChxWVZqphsc8Gqw3lmalGERr8XIP/YsLG3u4rLtzqP1pX3J
dMzJ2bF2Ot2kpE6oOULokvIFewGmIgT5XLCYPAna8CUUlYVv/8WG0mk0fKKAMpC3
/EltUkK2E2MJ+D593ETRWoLZKi71qSa/1Z5t/1yTmTx1Tt16dtgYPwxtecs4oatP
cG9F/fhwCmfeFZpfh0RJPRlhQJ4tT5bPV8dB+C2Pw8wGCijYU0+72alTgJoPeB0U
OUCOOYMGeWN3KBoah6OLBm/NBsApXBjU8HKyTmJ6bXeMPsBUiU4iuKBVMrhPQHNI
/W/mHJWrRzR3wJ5tTB4WuBeqjhPKqEsGgJX84krNTLg+jFNiFi/LdRtM+EM/jn3E
fD+kezWsmQZM1orCB/2jjsaHoOp/otpXKj2Iix5hKETMpwAlRmqw4r4rwpU6yAF9
z7lnWzn/1veaq6zMvM2KSLIV1+FHoZBNUPx17MC3MsWhPdwTo3Ip9XlGIUL+BOuZ
1LlYx0vjdMJmSEeEMXnFSKN+cHfsv9IKupddzeSUFUNr8Y+RNU5k8rotvt3Byvo0
IkFKojDmbYGCT7gKCgd7raYtsfqx6nwp/cldjgh9wq0bbot0Dhqm8+vM/NVZgNSs
uWHE6nKLBhJQp+67TAYN9HqrDz6KKFHSC0g9klcg3inbpXFgY03s8t2ldzPvXgDX
d0/H7qQOwJI6qA+ghSHhLilbMRkLxm6Rtl0jGFHcfrJk/QNDEKIgJkptuodUvRz4
dHyoPSLxr2W8e2CmQLMD7BU49sKCq7SfTnosQ9/bnZgBeGfEdxlQ6xg6itqB8Hwv
vv1pWVpV7H6ZSjzOgyAnnm2eW5Z2e43VQ7mQ7fuhkh8BhSFMaqTlYeb7afoqpoSg
KaKcZGdpwGXNwmoqVyots06OpJiB5+WltwVl5CUvyglauhKsqPmiYV3jIa3N7PlS
qrZpSBu4Gz3DEmgFoebwExTFnhlLXsQzFzmLO+yxobYYf6OGlUxULhX0EDG8hAcj
Ks5VfyLCThZ2tpyxKK3kH0QqzYXpjUdigmWZvursWZn1oncmFJ68jRyKrFHFGT7J
qEFM/kLZf316CF22LFh5dwByY3wAImF4Kv4rI51ACc/+FdTj6S4kNKa9EaC59cmH
k3G83kcQ2ckdVMV2kGXppmEuGAiyslA53F6PcifQmru0xM46P3qk8NjWiK8+mhBO
XeI9doNrPLPQQjHU+4NLmdIqRZqs9bGbNti6aGcyiWzTkHh3jUO7GHiYP5iTzxhx
VLUQ2TVyqnsiwauHWdtkjMEQmEK5dnsYydxnWT57Wnxqe98UWVCavTVhbi7ITAxr
QCgD35DKBOGeSUVbAin1X9a8JuwVelPJga27O/Wo4cskUwAYUaks3eA9ZywfJuNt
DKk5sXLV4BAwgn6QLHxhBYhRoVw9apRBkPCF+ycEy37rMgHQlgsBjSxGJLvu2gHi
5Z1RtQgSu0A+cK0Z2oZ3OtksHoSmFnIMJVF/z9IVbOgRHV5ah8VQQXmfiU4oBLGz
0/DldE8ppbQwb9NmhpbK5dD7rKQ8oUESi3TBbi7Lq7wdBMTuYyS+YcqP9tUDF1I7
aOh0a8o9QmKe5Vr98EkV3fgQ+S47D6KfLcssJe76iqYtMCqVhbQspCW6lq2OeO+K
8REN86REaWgbhnM0AvuRCugD2HpOo959d2gnnGaiPNBXPSK3XeVTR3PHzn8fFb3O
oMlI9sjRHrlXBs2VBaWUzLHNM4AQHa3CuPmPfXgL85zfwa3QAdjtasVqw1CQH7v3
IFG7yNJHGXJ5lSn+k1yGQZb1UtGvB182a1mxDu4Ul9d5BLgEgMi18Udh1NRucAJE
AiuFs734wKprKGFPiKZGPGbBXzo1IikClXm18bg1m5EkuuN3TRmLFjxCKZ7H4TJI
Q7MTfFTtU9vWxV7trlE4uhguyiBLJX3Ky4Jb31kwb5V/5dKB7G901OSsrHhMPXaD
oKQV3A3ks+u7Ut5PYBOUvyjN4BrJ5Eu2ZFPXEJ+bZgfoX4WZ/+/30Tz2vi/cbVmM
LzPgAXLlwtZ4sM1Mvl3SYvDCCVYhlW+trObqXY8bP0emjPXv7gjug4z1kAuPPeLI
biEgOUiqIXSxMTLyMu9dFIsxpTrA+GceMCBPgOUz8vSunbiMkPzI4pHqsTbP64Q5
aT4wKVg2ST0V9k5qNxX3ClPBlxZeHA4QktWVFKhiIAhoYhWgZVecLvMhSTAClQP5
D9vyExxxpNq19PUAJsNzOPGUI9ZR7jQJh9Luoh1QIlFi3p5w2NxinxX5ok0OnR41
13L8As+5HkyGnK8twddWmITPqoE5t4xF3UbsDQB+QzeueaaWvaV1JbHfvI3k3AZz
oBlBbNfllTr9mD2dTcGEKtuJxhd1JHNwql1cw8QeBZPfqlQ5hzP7fqFsKRNLR7mz
E+sUEI6bcnhdsXjDYa1ZAJ7fbi+mC7EX7tZFXdOH/VI2hFf7WwJoRe162JDNFN6b
zrzXbDJzEgOZVecprHnMd06n2uGBvwbgoIJq4Y123oGN6EbjS0sYo5RP5drQnSW/
85G3S3DRVTE9i4RVA3fnUuOZkcVWeGBSMwSevZz2ub3VDMnhlOLIHrq008hN/uKr
EQU0hgSWo/6uDrB0Zlx0xE26jszw8ptnaMtPJVLpCYeK7Rup6sTPEt/kJc+BQAYv
FZ0fAzlhlqtAhZOZQssR01M2ZC8fhBdPm5hEmOJLazvq4C+9xvz2qfAZzEBr4oB0
v8KuAPuWcn6FkKPXCz142ZrYtvPX58w55GdfTDo8digXkbW9dDyTPc3ZWXLM/QWo
p8qW20sX0jArk1STiNeiADzYSKzxlEtXJR6/cmjPcK3cMJgLjDzu/u/GbjYKgDnv
tVAFiB7elwvJSb/DpLQfXnCoWNp8biwXKMuOQwlT94ms7NXw1SKtC9YgXahE7acN
1+NszrVXorK4eQgcOnYXCab2M7CkBeffin+zwLJg2Ayqr/VjnfoeFco2NMkcfewk
DVnfBgo4FhECLipKdRVRHN0g8UobjBvd/NSoQaEzXtCIoeqdaodCKwc253e/ezPy
AhANvfxCX3tQrWLmaEfpzK5hz2MAi9sRjjdVqKi0XKYa2Qb2KOzlDPDPL8qKjhK7
jWb1qrV2IcirbAhxd27uKhm1ekn9B4UTxe1Plh4vVbih3wnpr49/vte6zWOZxwR9
NJDneIp8/IGCMA/x1xXqfhrijD4v9nmcTkNSjkPUjIG/Umd+OLwo1JUUmO2e8Qnf
ggYk8CSTkNxWCnF2JI0mHx64w3E8lNwRsylVlu0lXPhcWj6UHWoIEtxzBgmaQH9K
yK2S0jVtd7d3pDM+ZE3jFe0TRH1bv9mbijvgqIM4ce/NhcE34fq7E6AKhFVi/4gy
OZHcE2noFgA7bbh9svljujFLomZ/aoToElDbRzIQ5oYrzp8xvbey33XgKc1AuenC
9CTiYdrrkzWjk3qn9286c5yH37wlVpGZZb8ZdQkj/5gtpl0BFKoZYFodb7nO1ktp
EJ/KqXsdIw9MI6B6Cq65W3ujen0Fh2lz4kvGs3WAJa5fQRa/GtclYgMLBxSx4N7k
QnqI+gi4TvoBxKsFcYA3e/2kMhtkl35jYFlh8pWyQOxCquXAOUvI9GHKQwsDaa5X
koatwpJfWErL6GLK/v+LxameOSbuoPBqRhFBaDpVxWCYHezM1rw7gmYmMtFZJ5P6
4gzaljcPJVj3wm9fXWYG+eZFExTaCFKPYamAhJhq4crsgWiEu3cjBKOrQUwBdksW
sEj0cV4SuQYjCQgFOVpEjQhc9/FZXokAHFRh/iPCdAAkrQOFWgMHvKVTWs+K2kMD
n9AK7sCF90vriHxFXUmMCFB6SCXch9FQuA02sW7BJPZ+BKyx4s3uL+UPEiy3xc/L
IkH6nKAHb+DHv63sZ6AjM9L7eJrEMjLLEloP0gwhaDiVkf7XY2jU5Qt4sw2kiso2
77X58fgzwpgHXHkM401w2b2chiXFvLGSEuJdZueAZOi9awRtIqHoFnzuAXmq5b87
jdExuX+3O8dRHiNX3zKeh0Sweg1RAQ/KRuavklSR5lpXhInuQy1tPDBwxvNW4uxe
glRhcqbu9YF47MteWfXwAvFsGTs2ZGfalJlsMWBB+WEqjEYGkMdaLU8hpFEKDdxb
ppr7QMVuq7kq2OZc33ReQ8WJjQ4XnMS94zReCQTEmEJvGzYOghRAtktQt8Aepcz7
ULeMEohi9T9AqLihowZBr+POsCkCsRUr/JWlNWlbn5MyWUKy4RUJNUlwtkxrqxfp
BjhZeWKU7hPuevkSdjzCer2DameL7eHGuVWDbClzDDsVPDwFlw8CkX+sCl7SG6eY
q0F0dpPPRmBjv3042b6sB642dvPKWyF6QTxmOPYCtwRknMP2cgaPAV+JutP6IJWW
zXJ3S6LILRUvijl36iC3+tQXzWDDRE4LCsa7YXDRIusaVWDg9UbpINSKIO1t4CGp
zzJjqylm2u0HGGC2nSD2ji+HytTxePXHsSWXKZfiQQYrEJokgtjvd+b6Suhd+2cX
a6OA8GPAhDko3hFNa+xd/5IA5X0+PkquFPbE87S31Etng0vTZHGdHnfh4GS5YESc
I4xm7N7iWh04T21fhMI3Yo7NC5iPYt7WAa2QoClXo0QeT1rPqZoNtal9SaZg9Iz9
3VA38ldlS7YCefTlbCeLlWlC0MZzbv2oRsaRUVLu9k6lB6qRwgON/I+1vMAI3CC9
qjJQbJojJg8uG0DeQJ3k4v+D2vfeN/eKY9G87KUPKX5GBNr+yCGKDejgqThBPGs/
IgO/5liP0knUU1r8navtTTXGHaH96M7//PaOSce0g31JnNzmKebE2tekaRvJu+MD
XPoVp23wdgDNZQdT+t+8hKo1w7Ejs1lg5gIPgxUAoHBcMllczVykZQVcAWj1owrq
FluQAE4d590kxuUYwRgjWAMVSC1WHYfSFYIJVNmKzWqDRyYpJvNPYRJzngC7zM/a
tUdY8mU7jfM6tuddf5esEKx4qLKUDq5HRGi+gQ8GWFpT70SgxvhM2rfq8dZJ2nFo
rBBPaRsQYWjIjylucH7BBeJiEaapDR2ooDVpVS1AE/shJwiX972wV9VE/m3QU2kt
WFH3EDGjxWH7Kx0BtU7Jxk41wmep9CLgIEXmoJx0i79WR+wL019K58QEXJ4+aOks
Fn8Ztb8bW4HSaOqxHCLqG1bzl2DsZq+6/i0j0yNaFi3d5Q015OFIiuVXmYhSnVyY
4atXtrbvsDWvC5k+caJOPoesedsII2minnaTwQGHoiqlDFCD6Gzgz+igp5epiuO8
p61mPlES7MixebbZMO56quiOAbX1MC6i4PBl+EFnxcDny/3RVpyjykjOvA9AVVlt
vUroOVhWsTCa895+RIkiuZlEcuIAOmQkH7uo98c5FswL9r0gSP9Rs6CKPhgicJtc
ESek3hO2plaDx+4ValAkJxzitZhSfYp3ZwsRvZUN+RZAHkTtwNNdRPhelzF4gjIl
GN0wAFfeNX4ZtAIGQ3wJWMlFjpyAXAqoRpyvn7Pbf+AC1GN2eUVYlAEZ66oh1Om2
BSqxCdeCWuqAymL5hk+u06CJSiNyFt5ZXlBNrXNLqeKz7ytH0+6D1mAisx/LC1d/
yE6Kg2VqIzGgJGNgXumUFOApcJhilFxgqhsVN470vLFIlXMTY9RxjRXg+7HRIE1z
WaSNWec61yEvqqKtNuhmfAYr88c3wGdpl8mZuPtNxXZ2jgltp+R+QXxyEGegsr0W
sjA3juTGA8aBCDFh4dJp+8gI6L/n6S3rn4Tr/cjukfIRhWyWw/uzdBnN+y+JkpUS
rbNQxJ5Ed42gd/gpsNsRO3VD+7WqXiTN3f0ecDWs/5igMIspYl/SYlff31J1+eSm
FkDE4tvHGIKonKEIGTjF3+pCV0XaCOtrKfzrpg7Rdem/q0kxTUduo31CDg4BUsk6
3SnYvMINhChlT2bl9hHAYBznktD3IcjPqPpcqXPCpBnUNee1teO4qLrZxSKUyDFW
tZPUUzKyNfLuRKG7OcCK7amp52FG9IVl1P7eOJBE8lxs0U/XWkSCxNUgsGd6UVtZ
vBUU0YY3cnQKZSKzI6Ewd7JT6NrO2k6dz8NHIh50zKv7GvjNYQk2cz/qfenH/IkV
cwGRip0fUZBmLW2HKkyQx3RdKoQ5NUG1dd9lcnb61KO6sGWkCdvfguPfh+yuc7kS
95B3U06ThWWyqbPy7TFEXagWnszzNGc13V50u2tQ7BRx7RPioTj7uaFei9NKyFt8
lgC/h/QsLYR7p2/67O7Hh0qlW2iu4h6S7YeAbFl02c1W4Q23Gdwbw5IMpvG9sekQ
zA75h+ATmmid0eXce3eNXYPwWa9XBQe1mqqi5MAUub4sepUEtzvuWi0Wq8ro9XmV
Qo6uG0bDmGI0RupRToJxEF/hcjCulKaN5eK63XF1wcntKP/Z1w42JzQN8CinS3EB
tzP3VQafomd/+wguVFE3F11cb3bW7CDD4Su15GppZd9PWgEx6Ogg0TlY7JdfAF3f
lmzye3XtxrIiFvw1Vds0JAtElh0CN3Brpzir8qnWT+O/KDVkp60MxI1+h5GRlQ9G
L1s9ajwMg37ZqOKJAuyKsVgc2CGV02VgWiv4g6kCyZI6MZzjzTTBHXyRcFH/2R+3
GQ5fm+6+eg4/NIFsUfIwbFkLvZ7dPFa+2lCNzO+1c5kVsUcnONfLN9KMTnX03AFc
DnGtxerfq1Kq2Bs4VZOOfdMugQQi46UFiliONmzAY7fhBqikbB+hWsObcne4PG6H
SXGSRj3ebPIOjznP8IIDu92FScal/HGmJl9KxZ6oYPsJpUXyIiS/MiqduWIIUD7X
Ft7MddSPIwr2ERT77C8cYEU5SSTK/L3a3nSu9cqhnKYd1h66GP3+sTQQSlUluWXK
AySsx4bhkRlEV+Es1l00qRN4NmhxRLwiVjvwFXGkrLQrNEHdZrYPn4LhE0ZCQvVn
IhXGL6WBiN+9gsX2jCYl2pTr/I/nU+yDxkuuPANPD/pTTMetdRBLXODoAC31Nkap
IaH1vnCq6rrvsbajXpyotACNAsRpK7Cqd+Cge2AozpipHxE7ef7iUwROneToZEgT
TTDDgkDi/vBe4qUt7fxXzlqFdzrRIYv7iFs96DUfS2PwzUhcIG/ErzNr/0CCUtpK
lCCa1Fxp1Tf3cQC9LYamW+tp/8LqVh/cWJk/ySHk/7YVEC/bL+ssnQ4aKMxnXhlt
CwiBThjD+Pmf+BC6qvxSS8caSRB78i0qrn/6nbylb3+6MYttYXBPSfGMlJtRbrdP
GnLlEuHBUkEBkpxHFuxhS8HHaYKVd11hzHreWVlQhAC/0in685Mm0gkwUhT1X84Q
7ESta5JQbBLKgb37+pC7aJRCTDj0S4Bzv31gVBosKn5Sj4m8cMy0Y9+aFcYmEVmH
lzLxw0Q8fxCeZ8O/WJaLVpWQtQjdsNyUqcYoj1dnjXpfr7JNUM8e3rvpEGQL40qo
m9OI8XtY9nCi60VVXd+Ccho/sQM9gvbjKGTXrZZ+DCs5hsfmYprn4ikw70YNd+RH
r8ke0qE0unee84XP2/ODPhwiqhaE4SX/E6NNIyWjuurIfKLf4U2bhiyI0HAwDzX4
byfC/Lx5zzxdP/oP/EjhgcH/GUwyCwVq+dBJO4e2ORVceN79SExSFguIjPmD/GYQ
clk5eNRoAql/c918V3wWvVSlet1dVvSWkMk7/OqMfEA2KWefJUR+LIpw+VH/nnm3
2Gw2DBw1TDM9vQqkXfC+SH55fCjDCF1R0tBjHgg4KBfYiIv/JRz9LXxlmMzDipRp
2h1VYC9KoHBuUM1zhfKGnHBpdFgPq2y2iVsrQq7EOZd0zSbBmg5EqDT+ZHamdyVA
ErjmIRVkQxoFr8rvJisS8+Oq1YKFwEw08AiPoJwQMPE4ns52bsFIB+vS8vs1qSLr
QoPAmZNNb8hw2YqBWsvrzbbpw+CpfPImFwnSv89nPfUBtZXGdLlkJ5Vy3YjbhX49
9SQw2ICaktF7qfVaOtGqLIXrQdaC3HGOREePKgiFxFjAiZS4yVUfGO6GjsvYAeie
R9etOV2bCp8E9701fwVY73mgqacUT257bWnxTcb0x2SasEUJP9AroEF5vrMWI5qJ
K+7/stNtrLM8b70Q5dv3UqOeuQ6voxWWIP6n3GdtvFAuU/D7GJ/eT0w2e8zR9VyX
GXhhxeQGO6cXUbYE7diboTNEZDuaS+sMfefFXGnfkSuI/z4Kz8jxjdNyu5849iaZ
dj9vC1oTwK+r5luTECCCwASNRPpeOpLEtY12osuIpsANc+6NKdhcsVBNXjT+cKng
fFayq/9DdSWndhilh8XsCn7hdksPYGZQ7ZeEzPYncx/Nx/uy7OahqfDtbS9hpj4C
4K71CWDQzBgg1gteVcbWHlCDAO5izFPkQsIwydooEuLBuLbpRFlsRbEo6JwLijrp
0ILU/oCwYKK2bmw/s4lbW/jpmU4a+hSbvpt4P7luAOTcSG8WPRi1/LQvkfq+YP/k
Q284ymZjisckVnxfjnQZ16VqWO2BDY15zuXYY3CegsupUnbzgsJMr4FG3tXWRyWv
wXPXkLzgiWETTPPIxKyorxDXX5p5fm9Kow07/K82XzFO+rR0R+cWjUDsKZXFaW/8
37mpaIkWn4SEwlhqHS/iQiabntCNfvQhQ7U6BeYFH8iuJ0SqM/mdTbwdN3S1+5rT
9FoZccetQoV4QTU2fSLdE26jTfX3KnfAAZhXW3vKDuutIBUCJaF9TYASJ1vf38df
U/xgYQ4hohZ96AW8lIQAKttrIjmWgy2hqsSTR8MpVFlxqrZv1P+8l8WMHBnSrD8m
YxCBh+l42EFbKIHkPKgeDjYztaw/9WSYK3/VaMTiJqQYv4uc6bPWxG7BAqAjkBIW
O69es/iSsGPmfxeKUW/7i6a24/m0r7sj9M0ynQeeBWt9Iywerz34MZZ20oeUqHwx
0FdcnGGx51KwjUrZQkh/QGspMjUGti6COCjYcqZBCklTu9xla+pmI6CbVOAmxYyk
WgndSXXcuWv83k5DgzIMTqWwRSuJIPICdaOQI1bcP5SUGHn/uJoUSUqs/8rLT1QI
9Qk+9oX18kmruHuPvhEq6O6DZ7gVQ1SxkR7xnBwl6T2Q0HizK3HicQY4c7cRNjzj
nM9NQMnWSL1gWdkqJaQCL85oHykY3GshJao/RNRQ4KZ00ZLmjVYY4kYVcTeZKSW4
0yVLf6gG9w7Rlul4COQBafa0deNOU7cYfrRaszK34nAFkEUlefUZXKyTpw8OL85U
AglN5Qq0ApUG5i9yF0m/WrR2EuX6oGNuPCv75MOkRZTNhwJHbd2sa8s30XDirXaw
ROsJEIJsuCuNRrd2OvSaRNef+e0giEKp6A8sQIg4R/xI+lkiTE6M+XGh0Zu+dSow
Jr4si3FcT6HuqdEF1ZFY5Gy6eyK0vCmK7gvq+Rk9xVA5VFgY0c3l8f0cfoZO8mHe
gv8DCWfqDzQMezE/S/1edUziLI/6Kdq9v2Ax9/nTfVaO3bhunTVrRXT0ZTZ6q/Ke
XeV0xd1GAd702ZQWKKtlVqP6vh9ClymDcIcXQMKyfqyk897/HeeAtvcaL0Bpp8Yn
3563XQ3nL5sKLDX8ST+yaQ0j4pV2hDf/RslScJtc50S9PYqwcIyIK2ECqwi6pTAa
/7MnK0EZUjKP3bP8BD7nKdzp1L5X7VfIQ58nUeLlWizzr4KNvIElcNqtrYn6qQt9
MGHst3VkixrmmGvefFFEAs+OkQ+2rHdNQN+Vls8tZEXYrjvonORbKkWUO0eI+uyJ
6IzO1kM/VxpKLLVF0L/1Ooh6Wn+PmkpFMneRlBMvhUzh7CR+Fx5cYFMITv2Puqnp
30KpJSkO8NhJM8ilVDmWGNOjnyepH7vlOfaesWAzICNl9Cw1LYTD5ptt8gVSvjfd
XQSTXzMNcwXJkPj0/tc9LCRwM8jr4f9iFXH70lln4fwJcGHI2GKBBYwHCmx59Rog
IHaib+aN/8GmcZCA9t2nwin3Ebe6NMcFMZQo3q66leBk7CiQO0Vdr5ef4jqFssz0
LqMwn7MuoZgp93Rdq94IaM+kjrxyR4gTFAudY9gtu8gAgFQlcvmnI5bcXNlEBiqU
e35azEknAVrsDjWxk64VPWW8COoTlf8P8r6BzDqGJToS2wSpP10x+KculrF8Rav/
ifTo4lJpnmTWf+PYlVqurtQx1ea1Y8FM2W/eNNNIIE1K+awBS/6GBkXiVPHt9nJk
3XPAWUnkSrh5Z23n03Vac1uIq1nDPSLsLdVA8CZ4eHmq2h9EbaUtNWRASwbS9pow
kW6LLM6axdFCGF7B/EDohulisxVdZjyWCN6dVz/iqB7r8r1PeHgONS+MFXy1JXVk
maUvKtxBvm9o619Qd1k+1HJElTVE/jlHx6TjVycLXq4lHN17wl4iZxNtAqpW6ooX
31CxcF2R4SYhPbpBYGB2HWfydCPmRuY60beOy/Okxg47FdFaZuO5wXoYIONldj/X
OjVYJ1uLOW6/CMkL/aXNXuIjJRAgSx/q/TYApoRre9bkdSz2XH3NF1oSCXKceONO
JDCEMHsXS6Dgx2qbekjKhxcoArlDAog57epXRw+bjq1WlL/Eo8Hwt46xhpHHeNZ3
TdgLlZWT+49T4tk0QF5JJYaUvgKgC/wsKUNqwwcDVoFv9SIPQbDY33Jcc0SiPXYa
o/KCOyPiCCOYlBXMr7K+fal4T6V5dC5jL32mlvhDcWSKTLrISxtbGQtn3VfycnOi
Qz5MEZ2E/Ne6auEcQ2LSs9N/7P8a3s9X2b6U1qUGTbnqPxnxCrJDomTdEbrgiY/8
VGWsWCN0jYZmRgnKIZ2VT3map9w8xZNXyhRlQj8yIyf0OKR1WgFXpE7q4chTerLA
3//wAop5ZBQOMVyuGHaZOavhSuYML21fT+IUp2HaP/LN+KzsdZfBahC6tc0EDWDm
DYRvtn+KVS8hrt8FwV7YDaON6TuSqjO/WZMEJ5NTr+uh9Q7JcOeRRLOEfMfrB3SJ
L7UabeVLxSmpa+XpXe5KwAIU0diZzm3tg2QQ02fG7AhbvbyzpSIwZhbvFIFEiz9V
Y1kzQ8/R2taAeHeiWeCtXysFCySPFPbfjv3heS9xkPC211jYH4NGcFw2W9kf+P+p
AnP3N3dDyh+nBrieQJD2YXBp+PNENWQrt3J0P+j52ii/ejjyHSLlcKvlw54Rp+K3
sC3+uWlVR0i21t0ualIoKn85SGUpsDVYQKesBvZ13uzP4zJWjFwryNfCkmhNzCXo
RGKENt3wqCpdAsxv0mY4AqF6SWhUyDRcFYS9TQlSyHujGoV0lkkTEa19y/nmceO9
YIIpx2KmA7ARxDk28aTLzIC/3/xw4s9fwA6UwGXXOLR4gAz+vNFJzhBnkxgJ5Bp7
o9/k+zD+Fu2YjLvICWB/pUL2xae/T+WqGjWoJen6d1M153tMdRlaFunBhq5zg9D5
vgIiiFWlratKuZS3v7q1PB26ctpjVdd+FFUWcpSe4ggfHSIOM+PZymn5Ewt6lUW1
wwv/DoD8rWln32DnZm4A/l+Qw0HSkzJEJ8Og26rTKhUJ79AxO0MQsiAu1adYJthh
C337nu1Qm0tK4KSjYBSQjXS2dUmW7FbkyudFRxAkGI3O8QYOJyxWnF2ZwsRmSImO
yDaBw3NHErIznoPuHyarCgwfN3YSyqunx7wlG2pqHm6nytisxcmn4ssblLM0mq/8
1xViIGr9PCexmfO89hbTKw/0f9zHVHohHwcPyHGX5STWSF/dnK3lpEJb8xhpS33G
DMPg0mvEg7D+IM9OQVdf9YKYzcHAxqyXpSZPFMxvnyg+JLa5+BXf+Wc7XFfGOLZj
/txMhnd9Ozw37jfk7P+aii1DpqCu0fwUa/vEZoiQO2gNwTGfGeTqAvKdcE2jxdFM
3A7UfracEiYzm0XIs404rJH+yO3WElwUCOx1TcHzUdldiJKD1mHznmc2zhtt65tN
4vFMsEAjtM4elkL8CvG9tPwErtTMlbUrePtbvwSAQm+clDYXhweccls4mLL9iUBg
1TQZdrtPZ6/sga0L/sdGKBifIF/n6WJnlxnzwhurehuPHcCgI4O5UCfw4MFJ7TaP
smE7PqWXcorYr8u5SXsgyifP4U6zG+oar22+BlFfAAlXBYCBMdelbhrR7xIxE7lk
Qz9VnmAG5QLkHhKF6irhOAXRE32ocO2alFA/myMfm4MjiVJg9MbGaRvJMECjUv+Z
wqXkr7HLImq+jRpBTfBz5ALRjy3EA7aT97emZJbhViSKhn/fnzUWCjcd+wK42Nub
TZ/A2JQLyzrKnIHKx+DDdrol5iHEDK9IzBRngxyegrCSUw5kMZwhY2R5Y70VLhNo
55M1R7g411XOYthJhV2C62rVLMEQYzw3gkAav7qxV0QOZ1fF7k+MmGR9C4EbIZyi
mhwyNfH6AzoHjrgPmXnyWZu+rUm17y633+Wl2/3dkiz27ty3ab5PeagSJ1J0DC4V
2QHLYAIXndvDxRe5uJCltMNKrXOPHARb+beVkoidYh/kh7Mm257NcCHbrPAJM9iE
QOoj0mqaUbub8sDGf31/EV5W5eAhkYeyj5P5BX335bZsiGRoKaLDwr+Te1E78o0/
ATMoS81ejuq+iD55fDqnj30yvc115sUhSW0gijLN9AudOpnV5VQob8+cz3N8uiz8
q68sPLS+H8pj9GqN27BZxxfya4w2dCufG+QVvGIq2oX6uKs989YEM7K/CcUWIwVT
Ahpe6NTDsMOIH+nUnq2CA9p8cimEhktkH05aoppu7UpdfikB81Lcub6jmKMCwEXI
btj4BMp5yFMikQcbfcH80OLNwJJjwvUB1t7cWNXdGbZ/gTPpv9Mg3xridFSH9bDY
06xv5C/rTxtjdd/th+zMYg3vX7NAegH96Hx5LISENIye1WcK9K5eKRZNx4MCCfHH
jHGL+mZoudBEZJfZl8AHLyoRSBXZJbKH38bGkWSYHIiYRFeehOKu51WNHXtzJgzt
IbF5Vs6AtaGRNRWcsGTXBx1Qr2mGriTAtl+CMSTZNQfXtHblTMEb2bI1WIfbVw5e
QtvIFBPN4F47RpNI05mOzbnlNrxJkLRSs2mC3lKprBPrmADHgIAU8XypQ0PdNHWj
CTnlb2yWA/Fie0P/d0nSQu3vMxOVjDcx4nEy3KP/dYSNqXnpG3SKcT3T59QXVStk
/8pm0+GZm2ympPSwYT3zgNw6aYiQhjsot6WQcwh0JtjLYiAa0NW9MkLZuIlKKz6k
9QjgeN02VhbQbuXqI2RoeGlE77cz9ZM5P/eMNLrruIZvQAbZeVddTd+QAuetA4sn
88jQd578fbrEZJrbdv+xR8WVSbZDqgoUKYf+VBvJo2AWYDPH5YJQyW2qREpDx1k/
mNnzKBZkevSW32Yu7+JhCXp9REcZZhppkVo58HCooLYdQD87gDF5jq/TBYaLzhYz
urPSG3CeTlEB5rTnQ2WlEAjEWIBhSg1B3aYvmO10tuGEacyzIhK5itwt/3mUrBmD
0eG22E8sCKfX+/2KANgL2BMGPK9K5OpBO4qPI83f0CwMgMWLTnKd+baXmZ2W/MJF
fBjOAWEm1q45iNFesem44GeSjZZ+q/vCjxRL60iVuFqDjl/tAfjiunJ1Vh4ZOeWy
X2+phGen47Ik/wV58C3wg4cqlgei0XoQ1Bq4zOtMZTbfjTuhcnWb/Ny4RaqT09EW
Bcd4NvyC9StMBd9l+5lDRX9w0HpR9lqXYyKDyQjRBsL2B/9s9m2WkfrHie4oSyAn
jfmgpSNwSlwQ+3Buw+1jpMgIk6kunHlU/iJ8plQXIpc/LZF3ONmGrW/bOamaBZyY
GgPi0UslOGHZVeOA1xNf3O+el3Ocf042gPRl/Kf93kphee6u2qL/EIMV4xMEE/2r
Qe13GbeC7UGSXFbnPdvfsEmAtKbCG+Fz2YRIXmRtWi0V8v3CE6Pr8eqW/EyUT72/
g0tjKlnsox7EBtwIMNCblyJRSkprci7zO0y1SWWjOxBoI9fM+5IA7zgF76wYFHOL
S/n2fbwPXMOcRzAE8AVSvwVIg4uL2AMFffiD5NEa9B67YJ45rlJvgpVcwcjmW3Fa
PEuBiFEYk/a9eLrghrb5+3A+DsTe5RTy/cCV64j9p7CMJqSNJax8jE0BEVEEIBZ5
ZaR498bKCcYK+oBFmylcp1BwmigAkTgRjJIHeLPJ+mAfhidFziCxf22C0Lq9WD++
MWuvCUX6uxbHsoB3S0ZnNxxnTaDt0RWy8x/ZDQWxGs+Mn+GtNxrVYvrfgWQQ+jy1
WK+JA7/RXU8LbdQinNfT7tbvv1n8f7m1Wq073xDrhOKw7CVIQSLO+laXTjaO20Um
sDqWDGLmOOyY8GOy75RtTnATy/Psm+DwNszgA9vsFPQ0wbowlYSyBvVOO3m31WwJ
j6dWfILS5B44DZn7EepZjFUX9EBij9RimJBThoD1x8pkPoZy6cgTlC2N+EPwWskm
uelaP7vnaBtrokl+txwRZ0a1TfuZXS66MIfwAPU8sAZcf4gtcLC5ILXy3zzhPCr9
qpuOUessUdy61jh+K+Jl6+eyDHq6Akw5r6LBZbjmjPWSy81jcCx3rUrt4Yg4Wc4J
/6RKQbHLFGlvRLafdi0exGDeMF1Hkao9c7Nu1Yx0LjSZIip1tjET3HIFphikB1Lg
wtuPXlMawStEgCgnBrvU6/AJZQG8ERf6JC1qljHJAvB2wGwtZccHjHX24EVP3RbM
zcKi1ai64QgLAL3kK2+tkcnUFqbpNqI6Mx0mvK/KNdraODH9MsGus9hH8xrhqgW9
HYGAie3HIL9+EKz/gobUD+YnlP3PupKjTPTxl5Xm0u09t0jhaahGul/5BNzvTcd/
bstzT/yT4VcQ+KQvmO7o9JguFl2RL4dMSKTjg/cjoC1Pkyq2Rla7a+YSvM7NmGrK
awUI2z9azyj3q82c2Jd4dWjgtU75jO+Mjb+Hb+Jmk95TDOC4LBbveyzAA3/xPs/Y
R/iTk0lzID6KBEG7ul780ZlFDKHyc+n4DS+8B7QMXE6qTNStO3wJnqRY+Uwg2Uve
XvTj1gY6W0Lx1CBdT5gOqHPWkQXQ7L4WrdnPMfN2Ox9X8XL5tNNfq8iFlOoOlGmc
tHKc9AeXomN+7Qm4Z1Sk8R/7b1/jXSfZCANC/sjbXChfskqhPMnnmpx6c4zeTcZl
E9VK4YeQS9i1zUvfbDd1YDk1jHEh2TEYvsNf19cbH1cj13gQ+Kh04CqAVfe8dtaD
Ka7kbij6de7gEzv6p9Mv3EKLZQkl1iQyBHSWXAOI3bhFkUsoI71tpFePmSZxNh2T
KuW+1kYlr/loYXBlymCmDCFuOyFW6pc+iCNpgyi6+7bCwiQJbl5xam76iI9bs7Wb
/iojaERTOJeIFh+s6rwsdPIJWEpWO3eJXl8XJ8xCC5JKGGwumIvw28UNOhOA8b4o
N4PjhdzRNg5GK7LCD70Ai7AvqtzT5jb5u49HxiCtnXqcWJB7DOOWNBXF66BcwG28
B13feX1FBBA78jDDPrxdhpiRT7cux41PKEWUdBXXYMYo/bjVLekPJSj9vZ216HYY
2lPwFb0sXGAiuYDTOBd+S0N2ka/RNAmXI9xLkvXN9xMRdPX6NXNCpCFnRdUHPF6r
CtuELkBX7RwZK79m25KOYEJj+PBdfVAJOok8er/rpjvbx+Et/Lbd03nnSH3ox/+P
ecPi/SitlbyAVfVNLOQTfPWrni/yZqf4WSGMwBXI6X0m4iP/Nnooev7/K0u3e3zV
UpwD3wqZGs30rYvvl/zzcQXhnl+JtsN3m2q/m7K4LJ5DQtOrbwBGcLf0C2+By70/
z+D+353vNb6afoggWqc4Gh5nIrR6RiYiy9FdEB35JCUtzq9Mqy2UTwtuuUPwuudJ
zU9ERYTWUDXsu9XlpJsjsqkmdqX2k1GGPd5XCUsg6xMlx2OwTGl+5shZ/N3tVtNx
zNLBXsxicPOe5r0L/FNmiRM75o/BiQmMBqm3L2kEZCvQaxJr6A3OwQYaxgN9QApL
OVuoCZAQfbHNoVP0Gv5cfnolHpeKXNF2pyH+P4oS0DQb6JhH75FN9OCsyY8Vp+Pj
vnH9Ya1vJ/vlFJ1lXZjbUVyx5ZVtkv7dvycyXKX5iEBtSd4Ez9K7+qimvYAUyLOo
xDFthc9qRxekcLkva63SCAke3XAxxxCOjofMN6zW/KOlddMswiVqm9/jH57MO7eD
b7vcWG8fsvx/gUUlZEU1/9UujDlU7YvDej9G0mo/6jZ/u/95U7g+PhG0qfJVAru9
1OYlBgjdH0olqrqsSGTwC8de4MH3cZNuM7l0FkHdALM4N9BZBTDNdv4kT5OQHKws
DQ8fRw9GGn0u8GG8YcP7ojNHoqfD3Gdkibp5gCnVQ2QnVHXmauG7eq5QuA7xe7F0
OF/KwyxlMJkZCJOdk3xQefyc3tK5sREJiSn5jYWFzmXjGIXgKzp/1H8ZIMvRmAt+
SDceQEuVxxHqwh8YKnJQZrsJrQWUbEEmA+Y5VhO0S/pCfl8/GcpTovYM5CMP2/RJ
JFOePbNSFoSTXWwWcleEU902BMACx/ocNb+4ASWHETVFB1RPdldMLaOmN4aEwNOS
Eg4k2hTG5WCN/iT4/TEu9Zn78M5eI0YR0GoNKc+xt2W4Dl2BsRFatnX9PVS8b3L/
BJmaeLfESUHzdV4dvNltxlxh7d/WJVQDXkNPNRppI3844NhMAWHvCHq8OuRWlHix
ck1+qO4EQuJWsBdhL0x3Wf4VwRsX4Xhrg8CwLydRjk1SuUdVg9hamFZb3G673I1e
bsv/z5/kNOf4MgrQZWpv9rqkYj0by0oJlMoLBOoZg7Tg9rqLCeTGi47BjZmYav1F
8HLZoinfRsfqLbKrceAt8niF97mg+bfG1XmW5pOcyP3wNKMOaNTYTH5hQiCONuQE
B9BMhIOLMGtj9onJOMakSsusd49NJhXgKd8vnvbh3jOLtKsYki8JcZz8jBHCjMqP
6ZzCIobj/8xNhGmng9X2aOGH+1xiSXZw17R9zSigjP6HiT2OQf+tsvNnpWetvmOO
/dzz+mef7UcsZQt8bEZblew7yKKSIdgq6lRUWdLg1VYZV3cn4I+Mp31t3/JK0sXa
qNn/u61WAAekxv5gJB48gux44igYn3Ac39P2U7XsrjsVcwVXb6MdPUK+FpUjtQr+
ys9LKqR960tFOYkbALlnaBTghZgQat3ZC8HoLKaHUpi9RajtrCcR01Yvv62jeotg
ob5P3RW85Uirzwud9atD3MuIMm9kb0Dpk1ob8QDx17c233B/hJcAk/ceC4nrKJTZ
6X8LBzBsQHWmLMJG4/Bb9useAfMEG25Bl8iYHRGxWpws4qk0Sk/uHTHs/W8nAORJ
ReGne47PNB2OZLRizSPPE1tO7PcZPmr3d1ywiFxu4MbfJMJkacg876kOlYDqZGpZ
IDHQtZLJoXLIhOcn/SfqMtorrM4yKdIX7rt5BDTSlFPniqlI8OLXFEanw94RDCte
OYSDbzya4lfT8zxioJS2taXZsL5eJe4vOTK9rzk9jw2tj1Y4iRk3egcECz7Rhl+w
vZCF/ILIqTYvR5FdJ+cM/VFbpcmIb4eyTzewfqpsonlAuV1+t9dXW7PTJcu6jYQF
4hY9bHD0ABi9QtavZnKKp+Z7BkUjsc8ATdAW+8mmE1w4XORniZUx8wncIcAAN04A
2e4lmpD6DTdrJYMS2HjW3WwbTr5tf5xpt84AVXpTl5vDyllVpKFVLuGkNuKqPEs+
jqKm5UpG0s+0/172y6M413cnVU9XpXWmdDCi04yU6ivUj/GvhhfDJiZMVSweCoJ4
JM6XMeI3b0ZHS8OgpSWzJf7fEs5siXq0q0VOj4EZVGqqC7WFDTR8SnoXcP7Rxizl
ooMt8zlGqC5wQ5qk3RXvSrDyDX9ZH/8KqF6S5RK3QFYhcDbaHKmJcmcZyMHrJxZr
h4SERg6j/LO0AN52C+3uwi08FSPP1xD6Dk6OKLOq3NYNXPj4TO1T3JceLDUCFvf5
SHNvvgl5c9gn99xC7VHvmbwQQYaqqaH8a8iV2jY4m3njYKeOuiOmMqLx/fU2Y0T2
JwzTXn7uelgb0tcLWdjOc8QKnmpYg+9fTL1pAVj6Ri6MCKd+hEIg/segfFc0PDtw
TSzNA/bOErMJsP8qzGVM12F0ha8MRjXvmQhBOrNtJp+5jeDnaoDnW+0xR40+oYkX
vYv7tKOY3tg37ghQyHm+zzQI9eAA5PaVVvI76xHLfuEFcdh1ypa8Yp2AFbaTnCfD
xQNHLZCG0uRjydxR7Eh9X2LadTqzLAMJVoO3438QFpyfuxUsULWN/r/z/a++BBHd
R4MLsI+wFUwQHx3dQ5zXTUtUISPNhLfi68PY99FT2cMcOGQeWJAXexeA8MAqBIkH
XJAQ3dfmxIdSmdpHKHkhIUBTHgw2SjiM0isXHQ00ow8U3mWj/ZuWROdJVKoSvU0X
ZiWNea4VDPXapaWHxe9rfy33pJv+e2bXJq7Co5I4lsr0K0Wrn5bMw4CPgr7tu1eG
YxPlZxHKwh0G8fMiRagO9D8bwiW7E5zXFJ8OZphvCiye2XS3dSnISO3Zy2CPpq7V
90nwWs4Ljx+VMO2DGuRbhlowqj7egidNkhniMAyky3ShdjOh+f01S3ShPCvznGCf
/7bdBecwQgEm6eCFcV6BtoXpbrkX28udZ+HB3KXa/+R6795kakLXXsQB9oWx6c6G
jlG0Do+DxE7S2Q/31iVzCQFIgDnODd4wMq+YV2MZdZsVuFPcU8oxZbfZGNzXhumM
kPYaTyE5+hTEXPsgSK8Hf4zC3FQXCwWCwwh8nsL6UiUOxy14t2VJhxD0JsVpj0vx
REdf5YqOMCkeVAn3r1GL11jlNxZn8viZgPhNwE2NppK3uf+PKeyALCFvaGuiqfT9
7pdtq++ht9VBifUsMg/t10tlmsC95+W8tKp1OmyF6Ef7K5FMnkN19TMeUIkrpBMm
1aSds4Ev0CyTb0NSwLWVn2n2GPW9klw5gDmigUF7FcHHGt8tk4ba8FxaEMpfz8Ql
+FGPABGEVo2sjDHDUYAyEUCZpLE1kbcTfrUYMY2QJKuwDIAyCwSsmxIO6hCvXIA+
rEEiepmjR3fevaMwQ6dH1XNuTeeyI5qwMJuDUjyzIET1AAvfrbLaW5gSidjACPc2
80FfCB0Yibn+Q+Ok6juqhvqr0XfhWaLykmC4eL8BUisifVP4zwjrPdfHV53AA8Je
wx0GIIRjNpu+8O+iJ+fT8A01MwIqBoBYuFZiAa99tG5wW89zdOhWpFUXz41SvoXy
c4SO+tyfM9dmcuxpLVilncx55ru0RknhIhb7JGRL2Y9QkitBEGnUKTaqp+g13vkl
a2ker/sn7Ec5X606IdBibJXwcIuj1b8YHVyLzTOOJvlmFhqApg+5TLs/Je8XmjHi
n2+EiE8DGq2Zyv/AQbML2cPduwHMq7wC9Zs4eaNTZRbnsb+GsfQr8HHkf8uVR3Gx
ODaIv6Si1U0lQ6oZlGaJ75E26vp30io3WxOzmvj/clj7K8Pjcrv0qggREnbxdig7
zgApAzTxTq/cbcy7yU6KdQfuHEhN0P4HgIP3YTTBIuxX6EmYlqiQxxQwuMahSSF7
7RxjvUEC211sf19ljmEwbsl+N4YO5oG3hOZ1NrmtkHOmpEicfsuSYd6YibPoyxaF
MLnGyWBlOwBuCj4syMfIlG5C62gTMh7eE7PFONohIqDA3CxyjhfAhxePCtkN+ynq
UebdUnREVbi3/JobSvbhnECoCpbNkcUMtYkl4Y3v63SzmUoa2ZM0OGQ+Gjg16z13
wgtg25r9bbYoCWdEDyR36MZ36OSHThHNJ3mFyrIWMnq3P34RpQuoCHG+huxh0Y0V
ZPHM0hdj/+3ootHjTWqy3BcM/iPjGSaqeinx+HR6IlaaEd5LhlG9dT+zufoDQWgt
/o36STEgoTx7qNXVHAHvVZXIKCvD2mX7RcrKeW5DfnTSq1/U6F+JN0YkMj7NICuP
qmpPdnPjX57xymNbxh26c6EG2OQh4qeHJC2eUbaOILcT279cRE/Xq9M+THBMp2Az
bndc4f+g72sr7sYi8iw9J5EvdM/8mRvptwY5Yu2zKvVVtFxnz2GudM+BlvqaCF8p
8hOw1CifLj6xOSuoGyqEzzGdDVJzEADhsZE8SvxetwIZwY4tdB10ZPZ4hkPMTow0
MJCx8hvJXRmH7t8SDWUwxDmuXqZD5sptfuD4nrsuPpI4JwIW1uHhE7sGEQwtb2mk
fpcwTNy0eVy2xODARSr/3zy0Qtu8YtTCPUsQe95ZOzl/4xE7gN3HMT0RKkHBK2sC
gtUB1L9lodE/rCFWLHp+A3lOerUJgV9bGIk73K3oGiaof29qPiQE1MbM3oM0cVGZ
aUID4CVW+r6J5FUXk5RSl47PHLl1P1gCphI7QspMbYtDUfnLoyaQPN6Z6KkQpo/s
t7BfJkZiQyjnYqiTwccw6QMQeSUF7fwiDeB0CjBDdB9Z4VJdMt8mqYTODNZ8k0rl
o6n1lFAy82+3n7eOYeaP1FWtfY53+Sip4P+/QfJKIm4xWB9T+TvzN3EUCH2Ygx49
Pi5hKfWB35BZOesLrcd/wfC2nlnd5aCs5VhOHiUdsFq5C4M+Pr/14m7LYyFLSxAo
M7nZkH2EOooR2gGng2uSkaBEfMYzVGRF02+VSY/skNk+ZooGyyJ+3mQTifgi4xTz
kWjruEmkrJkiFxy1Pu8x4JPAGHWs5EeL/HMUGqezMQadckFpsWVRnnTZdndr6J/U
5c+n9QrY/IfQDkXSRq5Q9cOocgZ21/AIpeN6ROPw8pVVt+UeKaxF2Gs639LXOSbg
rzRrfyCGRfbXLwvmjVFluwYPtADZPgV84OBoWrtmgamb0sEWebPcMj94uSlyy9no
y4R0yBO5I9U1b8b/OaewdAe4cXf5hNMlK0MmvV5O5/6zmXROUEvlV6Z9HMnJ30pl
fpdzeXRSi3IkaXFgCHk0Xc1CIUN2cbYsNOKZC3aMK5oCVDVWcAjX9PjXySf1xwji
c9zyZ+BSxby61NLu3+xmgvEMVeMSe2+dnmOSw38GuJ+gdDPV/fSi5mh2WAVsJU9Y
LmgCgoluQ/pzhE/wRsrv64IzYUshsukW/r1tODcuMlLUQopxmSc0d7U36VL2h2bE
U47+XGxJXENZ3odBivJAioGZBiRpF6td+uqjBGmDeTMPOQn2+EYHJ69AMSVo6Dho
WcPqo+5D/Ns6Ho7lC27pUUEF8qT8mmHXyxSWeKEYaiNd5pER7AaebVoM+NJfO0pr
J33L8AsT28R8MVintrpDq/CoxRf4rqUeRcZqDb9EQzmN/6esKLkdJLyPzBQp2edK
WwY86/YvrN2O4xCDhiSHrzr4J3FwVKPyTYQW8PgvquUbXs8Z2xVwsVZ1jDgcXN2G
Dm7EOkI4OzLq0LW+4hT4rSnMnTXLNwh5CHAz8v/W3MiR+laQhKagXzXDDzXyn45L
3xJ8GNoV96TILevtUO/BPf4b4uD4HN5jJWDyg5gUR0AqmMooxO7JElYRwHyxw6oc
LfnuD5X35UmL/ucI25l/XQFPy/sA5CfMwQ2ORivOfAhw+DgXvLjMsWbJ2qZXeMCJ
4B9p4ALxsLvgq15SAjidpE6zqKBa+aa2vppbUUy/+TUD+hQD53uMPoVQBKU00OmR
KXQfilLgEQUygiaae9IkYGnOvpRr7kmHiNGyiFteiPG6bZqQTARTnoqTiAeyQRYJ
Wwh5SAFRTWMkJBYc+f8h/5EBmnGdHTbNfFAOXtS98kK7OX2bAvy9JMWv2bOBonsU
798CQcOOF3GImtlOmOCmIzbC/TGdNK/mUVG8Yph+fl6qmw0iNeswvn6LWnxhnev9
QSV31Zt1mo8Eqkx2sd+ik0LxUOboA13x/Fktf3KCoCVEaD/cwzX0M60jS6qDM/XT
fPWaxIg6teySThq6kjL7caORnVMZ/odCS+CJUmQcISmDMYhNjduqVTbS7VvTgE+T
hSVAhk/rtmGo7p/n29i7yOWhbfzILVx0apel35AXqxsNurF52SfTCpYMUPzPuS5l
GfvEjW/Wh0P34SN65/0exqBMhlCt0BXX7IO6tD0tsxjP9qPLf7PdNB0fgp6MpW4l
T+fwwYHsx8wqobjzxJGJpUMi5NusoAI3DXiTQVm4ePzgSd518xGJjYflV+hWE9Ce
hFlYtBIwOuz7FuDk2wzUlgpV9S86MgCTsDrV3pa2Y02Lv1NM6c267Wg24OOPQVTQ
2NdGOgUBLYMob8YdvmJ9JrwLauQnJP/SD8gBH+eaepCS/s8Nw87xxLpd1AzDbXJc
XvWBvqbg3QvrD+TR01JmgvEX7bXhaAfIaqrcTQpcY46zWnkWtdV4EF3yZaT3iWyK
pr9q5oGps3aNU/uzWfR8xb335Ns6UOd7SsRatlJZuod1wuY1Dpj35pVf/G7Ezer/
zHIRf7Kd4HJ4np/NMcZQI0ReDiirazgqQDRc9sRY3zU1dTIBRVNVEG28hPZ0mJmb
XeDqiksi20rc8Iia0rOGSnnFCov13I1GRwhStxsErPWy0Jo6qVvZqQt17ghsY8xl
N5qXeWoHlEg6qgP01xhvRgJM804dQX68A3TRC9W0XMstIHyqiSO/bhc5NOJKjpks
en8lPu/bVrEMH0Q66yrCnq/SpfY/QJghQ260SP8DhscBSKsuTXlwjC6+/2NV1QrY
O/pqY1tZljUX84GeRIHH6YAuMYoG25YXC/xSf1WyVWP6tqriLiCD58ptjW1rfwFh
HoqtQKJy3ZARGr/2E/KH+eFxZTsUR5S3FgNJDIHLkRjx3xP4krOo1lHVOoJOXI67
S/z8zPQcso1aajeJa4xcvqZCPJOehC6o6PndcGbP+vKJfONXG6PogH+4+7Poe2Ad
Y6Ls1u/wB8qJ8zlVsjAC/pi7BLq78OHlc8ycT+T+BRJgVhdJKucqBw75uE9mk+9s
EuhFJNntYKSABkw9RRYc8GEp1WrkOqWLDqFqyT/I4rhEh19pNFyiOJywXIp9MGKx
7eLOwAfJFFZ3FFtz3uzmIVX6zTbeQdN70CV4G6xw+uQ48znCaCJd8o0/47SXZf6N
w6lh9slLQmqGZ6kYOEAu0VuPomuOd/v0BZ+v2QIHS1k8nNwGkTc+5H4g2Egqxldt
lMOLlYVGUQpYjz/8ZXCQ/IjlhoU1OdqCKac0xfyHuKcvt5uUifUFmabgOEclBf16
i9gE8NU/YM4MSHm78TTJPCljwhGXiZ3rX1HvLWM+PQzWfyrLg4SpArAfQlyHgWvc
bihdkPakglORA4qYDSJtAJwrLSq3IB7/MaihOLX1rL6YxfBDGPlnz6UbcCut6EfW
shV42qPKtTPubKYZZRAcLe0bGvwMRDUIwd5Ehyenvu8mrsXrEykvq/4MzSqa+Pe0
L4GkKuvdl0XOcEyA8HAfeRg/8fP185SUg/0aC8kkCqwedL8Q/sKUFbHqT5xRX3RY
6Exk4cn2kbqSoB6TBUl22DpBoS9XmjBrKiFY0/dOtlnpBe7Ps3ER9Hq7Sw3z2q2w
KiJ4uCqi6dUFub1IdAgj4skFb2+klmGtol30lrn7aoacG/pjA4oBtVMa9MS1wX+G
TNmhcq595vUA8hd2Jj7oq/JvWfEHZjm2EFFsec0Czz4pj9qGhmVj1GL7b6YefuLT
myglzQvzz3tKrt8Za52b1BtVUuU1Ye7b0lvz41up34iIOk/Q5Gi4uCjedZmV5+oG
I3stW595TC4PknUZRsCwEIieEbc+ykfZPxWoUJJmn/u/bRMnAsGMa28rcXSQnNyT
xgz7u6yM+q+gX/LR8hQ7RMxwNFJRiGpKW9D9PEegLHtETxgdqlsYYkw/WkxRvWsO
ymzkNaKkD28i7rzw3SQ+hYK2vkyjc3jcy0ob1yEE84oFFq//PQj91GA94GoIeGHB
QdTQwcDg+i71rIKCP9dh+toH2GT1KeixUKZjyXxjbZ88b7DZe+d34lg5pWY4dbQI
7fz1oJEf8YqdHxAVeA9FUUFv29wsZqLIHXym9kz2uh9g1Gcxph5Ki9MJKH2N8itu
XZesyFxz+GnwitZmLNeikIKTSbmLlJk+MRfIL6wdKoLdP7boQsxK87Bkcba16hyk
LrphgwL2uF9ujbGTa/6aztxCt6Pmg+Ro068cVjUofvuI3r/mX7uI4SuEZtWjNAio
vxYvX2fqoaSJ8N1i/xN52yHM0GHG4WG3wc/s9ccUCMO6OVCxZM5fDs38Vnc6y1SW
nwuK1gHeIyMZSyeFvkvNRbfN0WswMjJ0r5Mt35LJGCW+pEZQDbLC0cZIf2jPyJom
g1GiVqAts0NTQzXQy2yjTI3qtowXoZCq/IMyeXJ/lmMhjUQNNnHpdxdmmJyx0m+c
eWCbb1VcTGLzoUY0WXnrSSCMq6PGvT4wjX/56ruj4nZAsaVFMW9sq9SqZXlDEsnI
DFUFmQ/9L5iFSZTMUvnCKEmIfje7plv3tbIDccvevFFlqBcsozX68TIVFtAPXphw
09gouYZSVVxoZg9r3dJMVTGIH7Zp8SYLRIUGS/zwg93BOJ0RMWqGdiz+4sl4eZd7
OHS66ihrOkgicSFu701+mQaEE30F3Qwc0Siv+ATXhKxvsOf2A5IEtzAarXXuDoSy
hCXvGrcadErurPffWLc1jMhfb9rfG4OETHXZ4NrRSFWpW3c+S6OQUPhKJNlS4X9D
lsn2UsaVeNXB2PUTrTNfOzlVrGj7lgFs/kumvUVOYv3Ye8LVIphfryEkX7M+wByG
+G2OSQ4REaN/+/vtDeITICI3BFf24z3wMwyREpgOq9m1K4sHn/tLOYTpVJ87DrVW
HUt9a0oDHp//7YBhDqfljT50Ow5iKRXS3RHW85ivMZAzE7Ph2jsrHJ3lLiYymGsI
kHSTRaDBbRYtOy9TTCeWwJU0q+wRf1w5+TG8cCsct9BNaL1cGXzPChzSNh//+2Wt
VdX7oqDn+TjOQFJvvpJ2E+3pBACEJrLvb9nzX3yzg8FfiMqle+CcJxUEqJOHYYUJ
gaDNmQ/J0F1VSV9omq8sP01ePYhgSgnRd+v8a917IrZPkrFrLVUbDWVtv9L8JatH
nfjayVxaMeRURDChufBtRCnSFlDKJthII10cYSFfTuxh1nLuLwv4xfJBi0RtnaQU
NfTUypr01+kX8zzheD/embCBJDm8VX09f5n9E8PKFQwGyUP88i3kPfnd57UoyUXJ
vOWrmWy48Wf0/nQ1+mn0N5X1S1gm8jpnYakJUmZuyKrD0AH4EAJCqiOKgQY3Vx55
m6curQL6JjmOthH4trGO9XchTOe3o+UJgmWw2OX3K95rClLZF0mNlK8K55TjgyiM
1j/sF4uKTLZIqwFVZxA7WlDjkK2+08f/yRM55Glgd7iozF7BgknUbd/uycqwBKud
hvwp57FElOifa7cFr5vlV3/wP7BU+iFVeDphcP0hygnIDD4IcKWHAqYH0hWkQYXc
fcNk/5WPhHKg7izcA6st4d3zPZqvLZbfsbXy4iinnWr5XMTUq4d/5gGpr5ZiZBdm
YOVezqNY+wn7vvB3bRfgi5ZXNMBpbAB/8qzTdTEAVFLvZTZsSZxo/TLG7p/EZBhy
EtgdUmkLB1HnOnMXKiqtR/bLVOBB0in8OIDmRHbq7WG52sgVOfyE27xXdFDVtRlh
Zqb6ZdURGrMnDPUOUTmZkB53IcPPrphP3Iah0Bl06mpiSU7Epqo9VWSZuEhd6o3Y
N6E/oI6uGVz+yXpPvdIeDGXOScegex3GT8R5t+NW2gB03+EuBlyTvCpolcfoiOU6
RkLkjoyV5I2ximOpfBujVbcLOuiSiWyYytbC1zfTIWfJg/yESY6wC/X1YRvcigxX
cfB8nHavjzehnGfLy2+2C0MA7BBOJX85oPEFFr7+KPWKdVhmuJ9SyEBXfvA9PdAN
OzWi0kQPUaysKIMHnK9iybzCa9u2WafSLPhrQ/sh+7Dnv/6cwxTe42tu1J2BbD+d
VH6OULqsV55jbnoRidWqx2BO4rf5iWh/EDCB4s6PlHflcVKQbfLHIxbTUBObXi1K
Ihp9+l+7kBZSghGM68ZrXH5M9uuIACIfodKIwVm+maJ0FIfhCUWXMx1RlIIyCj2E
u/s59q5j3EurJWOLXlxl4cZxOHs+BPhj2CFsaJeJdQF6Sx4Ha2qCnm+QgTdiPI/3
vT8QuCeQ7mne4qEOuB8DPiQOHzoA68/dBuadunujb12BZswm3Gyxuq0VCTAAuItr
R/3p2+97xpri6X461zIIwPr/opTEmkAqu054JKzV/lozJK/dLADelqEGF5KlQ8tn
FWxV28w4+H8/qMKAYjHzsoNNCOGy9lDPiARq+tsnpR/rI1CLUFsBaSmj0jvTgLwy
3DSZTujG8hdcP1LjtPzx0PKbSpsyQzUM+0kdXi7oqmpP0CA1lFkn78JXknmQmXwV
qvgbW8nUUM+HfKCfeGkg5f3WzqItuALO1YFDjFVonLl5q3HtdxRe3tTupRp1fl0x
AlFnWF/yDLJFTKJ1t/GKxT8odu7ryr765QUdrYahx5TR+fglzMC0SaNU2+ICPAmw
BJDnlOeguJqCAUHqMubq7Tk+caU0xCUAMRgzyY/bI5GLvlXw2QCOVZS3NCSk2qez
8o2GJ+S3syrHbW/j4WHevMR754EHkzx+ShlR0K2eV+1qRjzQnh4qeJkOnnnod476
LZcPVcFabDdIufZZD8jBGkuWHOAq7fqDGDLbplOV2g7iMtGu4LiSrLTr9aD6MNd4
EGrohuLkbMNesoRF+blLeR4E3PkhxfYb3cTrgXLeHg95/d2O7iNSnPT1nCBL17jP
2R+a4LvEfMY4bYU8vUqNqBR/Z2EAdb5i9exn4lg/rEgBqjmerbAqyCzwbwgABydp
34xR9wNBSkFaPaNTowHhFIdkNvOT9+/LuI8+xcm5SYl4dm1G7vAvJTCypOQ3Wjdy
L3TbdjKE2mdA86xN+xmmCekVZxpQKQK7qmf82g0VJJk/WRAdNAB8Bk6WVTP8/GkJ
Vvl06Uc1r2gQFY65D1DijfP/i2/baoWUWnvxeVlcd7tGHb3qdkf7Wogr1ya+aqfD
vByc33W1UWB41EUoUAiqAx6rUeeP1wcduCAJba48RFRr355Soq2zumBdl2dnLl+d
kaxf8LHy5dLO4TC/PpuUWkTHNt1XnkNhV1vhjRvEAmFxVtPhWrsNfav2QF55jaju
68AIvksUjiGG0H4FXlA+I44h+maZFtNS1a4ihS5/UKlUTCu4ABsCEHlmcNkRmG9X
RYaxejEXIplLzvCLYHjzn+EkzjT5kBMM43NnKlivdRNY9esp7IFFlNz0YFDWtJmF
FU8gC4YFVc/J1ccIMyWDsg7lOa8YJzCS2Cd5k6sx1bVBAg9RU0JESO9cOqndik+c
rfcb8zLg5/Tq4kxK/73bTPrtbe4F4eIl7PwozVSZKpTjweK8IZFAAzxfeeP9//0a
EvbEaGJRx0i8zLwpDlGTrXphk5uwLd7VOfzT2HZCfpIdMskRxmfrLKmlav0gklM8
ZdMI7saBzH8lpolycgWAapReQCRV8RxoGZgKc+Hp1YsAXPm7G+tI/DCqVkp8YPy5
Kj491RGGx/m1jhqn0njO03JJIZ2NaHKcLWAdVvpGIxcZoR0GeW1RdWmIKmn7ki69
MGO0WhYO206ysYUrQzMh6qtzpY9noDRKdW4z2EGsHbeWhc9Jbw5Yjzfi2JaF0jcp
ctYvflQODDV+BWuAUiULhg3Ojmj+JNNux2gQ69Vn0zFuvYjoWa0p3fqOQhtSzP7J
DVqJCnQmgAJWiF9fhSA8zSIra/C3r5RsfFs/hqkRdsG5v19YjIBqflV51CvJ8WSC
k4d7Npkf6T1n7Vz9ggmECiRX7Ld/Px08xEubd8LaO488iLPMyBu3arHxSQv+Whch
Ez8q2tz+9ErN0iwdX16kN3ml2JxAaaDrXj/rfA+jmHnLjJAOavEK32XTNdH1N0Bd
l8LH/Ca5Yarmd1VWayM+5J7FKlEXAAp+28JbOFpT/ixfZ0uFQJ/ADF901rImlWfQ
FfupHWfPzJm0VBYgReQA2ykfm8DEeApxzqCnFQFSoY5LqNQq+yuJShuQT1PzaWrL
GxCodT7FW6rAv9Y1Ym4++hg/muEcn4Mg3rC3rv+RTcTxD3wbg/EgsC0JW1F8xJYb
Pp0gxwig1zUXohbzX2qjWNjGzx8Vi5rd0bpaChAT0DIP/CzsPA0kAcaUs51W8OvG
Fz13oBRFvQTD65xJkaezQzKRmSfTqIPFHnwLHUnGnOwz8Aw0g1jHG1N/WO9zx3EZ
+Loiol//lBtHxo/dW2svz7ZdL4isg9b4oNyQrbMpRLfdUt3qmGL8XW8mPgma3qqE
CURvuR63hlngEJfcKddBb3v0+x+Sulc9oYrIOtFcm+S/Dd/bpkPYMVBZla8U+9/U
OITrOrYrV6vyivVnwvF3LHlgl4r1bJ7W2jCwBWUnh1gtNiNfVj4f+GPJZ3GSjv1X
0ykmKR+Hbuian75jbRYEDv/e3YFWlEaoRWrugy4WOVac4YiprhZ2OwBDTDMLtJ3T
NhuwjoJTZO3wymcYMHgnKRE4+zTKtFDn0ivi7H4iQnP9AAped0iNduXrtus7/8qF
PIvV5FnwpVaYRH6HFnaiNf6CiNJwbaQjWC+VIsKNen3oaDs/+veC4iOE1WWjF+Tv
p/6a3KqhQCh1MgdZQDg5VfPsDBEaMsfsW0WxlF47xiEEtV9akvy8TKLYTQCuIGsH
fkrunucdRkqHfO4SnPO03MJmz9dFl4ry3HksEbHv8H1PC0qZT1Jc1Q/XdFy5C5Ok
P1uh685+aCYQsEt9vZZuwCZ81CO3JF4XhQvIAIhEgg0RYtzJ9wYhZ6g4J+Slw5Ce
2Aof+92sx1y9uuahi7BxYHOW+jhl0Rjc98tbEpoNbwBQ4e30N/NQGJuBmemPbxMe
1xbf0AIBie+jAXzj3v6vGf6i+KxQmxDW/kchFMjvdH2mAqEx9EL2ivpscgYN/Iha
SrUCMN6eWdn5IFxDCdsjaWOpK/nTmyNuwrDlMnDC5pyBdIKsYkEaciaZJ8LntMaF
zZKp39xLHTWLzfwwAszIw4VJ0v/UvYE7n2Rg5vzdkzgsOG9m6BAIrFbMN35tXDi5
H7N9kggN2ru6N4NNVYmM6e9PRL/08tjHXBo/3qN2oWw7SXAeBgNu2jY2W1QNHZwy
wiAGa/29VzVopLjbNaKljno2PSpiaadnEdXAHIMOB18ZXWrewbuP+jAsL1khpebG
kJHW+DYL0A6dyYFqkE4jz5eQrVLU1/JO9y/kMFz8ClGL512tbTifmZMYcbyL39t/
nsj/f4lx9tBTRLtYfQHUKjDUIWxPm3ItIsIy6joKRLTuxSEStBBdbB0GGQD6RK7V
+IljH5K39kvm5rUi+yW2FDJmjUH5QCNKsTIYRWTE1nkLBNfvSLr9gFElQ/x+4U4O
gupr0894kx0udLYpqlHqbCzZo78vrcMCyVvGap6fVRcTgXphc7GQSzVoI7cANC2v
/b5ZM4LOOHhhY8hY2j1n4IpVfCp50samj6l4iEsesTROl2Be7hKVJQf5DGUJ+0/n
+ZY+w92Vab21ssJQjDeljDrYfuFHtyaEm/2UPWR38s6zlxtruZ3VCPf0+Ab9JdOu
tzAenOWJ02G5qBYZTLwAGFjUL9El7YgvIjFth4CS0ptpVQars/bNSzM2odQmTBCI
CNIrtRJb+WSX/WH8I1QcTeb7tWr/NuksqQqf8n8t2Wp9zUd4Z5WybKYKzu/z4c1Y
vFlnVatD4Yh6D92M+FJ0wcor1Nqx3m0k53/tC8E/d2kflvNINg9utkLFhwjQFSmD
xC9XP5l5Lblq/F19bvIqRSityRlLzgkz/vchYwsk77XPe6vWn1wO000OnOE7o5Fc
TurqtAsGluQGBMLRe8pgBBZLdH9rdrC49UC2RagzZi5slQddcdpoRZimb6YOLgAQ
S0npiDUn6vGzpqQpZpRUJjENNERpfK4IBHOCNNN0IMLuXih/zfWt34Lw4PO9cywZ
OZdnV2U3ZTciuoG/3NMy0ASvaybMKrxuIns3Ed6+hJS9sXbesdfOJjwisV7mCDve
xBO2ffG5+wEgN3HEwhWVvTpwAI8ifJyb/bqYpQYeBho7NOajiZZJ3Lp400TAsJTJ
ecjYw8Abz7MuVQM561QadrQfaIAtzeTVVHXFAXJIs0GgWeGrCdob9OYOm7dUBm/9
pTbXJd2rsx/SALBOj/CkmYDw/CQxvyVFqM+GtaVfn2n1TxYySupo37JjeUwkUVRb
A+WG7YS4yZ7i+yRqIX1icocTKJD3jSXWokCBl0WVGjd2nHKymyQHQTRpRJmNTG3a
d0gLLtjF8Yz6a0BM3O6ba+o/4aKjVYKz0PQlAar0L1DFNrTmJV0ghoQTf2OWEQYq
kd972+BIvUzqeacoIEZFzZbHYp7EZbwTfTd4S8LfK70qKlhqYMdYXq1zu32rwRpV
fzo+a4ylYB3iSI3188sFAYOdUqYp4b86LaBzwbIQM7C3S+k+a+YgEQgUs/3wD2rh
gGZG235SfeqX0I6BDARBEre2T83uEP/GYCb0/5D6xzhNG6Ezw3YkkA+fv81ukGTo
BFtC2Y6/6yKQAC7iG1QNm6IziGWCHSHyzESKv2tz2AGXoicymuTwRdMEW0CxuUPT
zfjLYcdQVyKb/gPJ/QF/yzZ5lajFrjKiDo7t4e0rUXMWVCGIMMqD87ZI7nkvh0vP
DGD4YIGDadVQQdOkXgAWfyfyGvNZs2ftODhQSLdRusgIcXLEgMssjkiUTVMRxHwZ
yr237vXrFotVCHpbE9hcSjRDNYEdJXdHk/W7ff0Xcwr0mchzkUHqrdyLJgWdykOw
Y5Doy3tS1dnnUaAbkkhebySlzH16QlTUsWV8OTixjLnjAYZYXr38s/Rs/zyybP4O
nt0IJkf6pZmgNrO3x/Kbp5Puko9BOBN121JgkSm0YMJc6Bsk7tbVC6GSjuvQ1HRK
/iF+4cImlLwbKPrziKhF7CzDhZbN7CDL1aqiHOlXuYsB5vprbeysoWtrUShU8d0U
+J2B77nbBFxBU29Spc/SWH6SKk3H48OrQG0ju7HXbb+503n3E1zUxWY8jydxdgSM
Ca4bZYCAeDKvIWU+SBNOA0uirj5dLZDs6UDuxJv/qumvZ5rJOaLe7tG+eClfFZrZ
yRJR70zcR65lmoyJb9JmLD3je0sdh7eu2EJje+yVAiWRVV2AdU7VdZTHjlqEfR4i
x2U3vbQ4zyK1sGZ9SjZ81EBErjcz6X5UyWYCOCyY9sXyzWgYqXWlg1gGuH4tCKoM
CinrxnbWcZ76tUaaN/eSH7Q76J+EKTL3Q1KcHXIjhWdJOPT9YGdaO2ifysenlhuM
R9HB+e/X3lxtq7Oaq7MTxjtXcSmetn4QBWHx38jWxgN0DfEY05fxTaQfeIVZYejF
Dl3MtPdVPecUi1n+ovJFTdQvdMQSTmXcc+lsSfuPRiqoezG+zxwE8FkHtAJCVSe0
R8xuteiyBnfYBi5JOJxgDXQGBSnW5blK/XjRXdgBGLg6r1/je/u5dJeaWIzYN5bB
t0ylz8o0Kb5kpeV1EHwLRnDCo3YNmhuvtesrmwslbsyBYBfnhVPHNzz/gu73eOm0
IRHPSkMoZKqPid2aHgoXehfSL7I34HD9nK37CvZCuh1rXubiJbTi6YmyJvypASy1
jmhX5LBMo4KxttqCjkzXh/WwwB/OsP7Q9i4Ja6nzgluaOzO2R+uh4RnuaF8L7FTz
KX6kaczz1T1pHS9es71bcFcyKkjYGe2bslezsv+xPh90Z/M6MR6B8TDA+slOuLxf
KyqEwHDG+AY8JUnxrpY0uMJHTaJDRJO/G5AE2yr+qzZPeui7EuWmyfvcIa3xDci+
fTrG7JuTlG4VuEcDOvrAl0tXuJWaaXNzAiX6MqPQlRq0z3qOjcIl1qJmSvX9lHC3
wHObATuSRU8qXQJHBXUAlVFQk89q86guvg5B1Efea0RZjA8ynK6oT3iQBb9NWLeF
oIt2qaoqtTBgHbOwYqpBiyZ2AKvJmqB96oFxvJsjOXEc5fdg6a0cLl6iiT9No46d
taLy++xTmbzCt+ALohrZnPjQDGdU0ZrliYBFoyPu3nTcdmtPoKGKyNaSVr3ODU2s
a9OQQ8oJE1bfw7a3YjZD4sBQaq/rWYQ3wi3jy6cxqBm+Gb+NGfCBxfi42pYxPIG1
GnG5xD5aJ7mhw3Gh9h/q83HWdOuFLMhbph+qK/kYtxqyTXc3oB7k7BVIYdUEzdUc
X3cVYJiOguoRTn+hDDgIHcwDLfJA0MZyhafcaFPOY1kUIUrw/3uyjYx+5qnMLx2c
/IFrtRZotp+w3dPInZVBCwO2kQ/zNQ/tgrDOswD+EX8u8JR/bTuFPkiUJTVIqLEc
oahtqQV1tkPyZZtU64ratPjWkcjL7goIMzKoW5xZDMGkGZ0mT23wi1tvIxrWZlH1
41vRscWNPV2OQTNvWzRskl6cZ7iEPrIK+zAe4TtZjUFL7meXcvYWtevtMIWC0rFH
DrMGu2ub5j35GO6e9wbvkd8re2lIiT0tiIV+CHnZusdiZ+yayoIn3PgIqBO7cXaR
5VUg2XTqFIBZRZz55VcL4THUvDVGe+I1/TOP4UcPV9j1/AluXxgj/eX2+w90/Xdu
EFfng0Jwtgjnnf208zoNAXyat0Jyye/NXbAEsmotNyhwU+I8g97bvafGD9/Tc0Cq
TNDrx129n1NpKUjbSIdVlq6GWnVei1dOAbkkFUV2EHCXPw5pIhQir9rWpCOQHz/W
kWRpYKYiwIwr+x3RYtrKYckEq13KFk/L2mJ8VPG+pEpBbVvDpE1wCs+LrQuzfjnt
/V4/lfJsnEW9hp8LGBsqSROM4DA/aT1THCGDfAxoEYFFCmODoHruq2QlhOCDcHXD
EuQ9ebflIaFxrBZvyp8R7nmdbQSeGAKpkA0BzZ6mB8qsxXBkYCmb2+zGzxbtOKBA
wXurv8iLI7ipd5/VxdSC5620f7srD/VIiUVgm9Pb7iRj/Tii6aHsrYKejg/YH7nW
9O8vfXLC1KwC9ApEs8/mzu+eyDpGPD06Va5gZhtBndBWiTbNG/eEJyEWZCUeDrGJ
xOiAYOM+lw3v3Jb1BdQZI9R0upKUYTZt1R9Y7SE02X6OQllL1m34vtpo3pEV5fjE
kJn4FtYOyR/Zop0ryrxi0XqRZ+ss6KlmL5yaYO99s2mGNtClNizTvkDvrJFQ0KaS
euwFPwWK0Soy+Z6PyTtGDKbJQBLnjSgrZOrdFd1xrJvT9oj49DWSnvq9tPlMt/a+
1vbcCvICRcVaRORDMnS32S4I/stvCeiFBQ+ocyJ92o9x9Kfb3cu2Nl4H6YjynUTb
zqO8GISnCAXzFBA5zEoErxgLrLE39bINQYA46nPQ7glZP7OODcUe2KDiLP2uKwkX
ECUuL3N4i9/EVR+FDurA8WxRpgGioBXWFf4ya5nu+FTPuZ6H1otgEn0l8AYeRePk
2uQyaUR1zRdGuCF90rAPws3fyDiJXISVC2/qFELS0GWuYeLPFXC6UhD9TmM70Ot4
eoUGo/1v7264dkZWgitYGSYIPPRtsAsWnIPYZdRzg2sRGSTcT9YRfws/nyKzO4zV
xZnku/+Er4fWzZxsaWGcspy/t2ydwI5Of92vTx4bSe9ITdjpHKKCw4Jmdc1cV612
KEQ8jY5vdYMUj529jc88WKbfaA3YpSSotB4PVmckF6U40vwhEKw2RMzWwFVq7ze7
sSLCJpuquOqsM41KyXt/6W7Oj8oGrXgJuhrbQRW+r69oQc2I6IxIA/QMafIhjCYb
AUvDzEjph/rz55Gn5VlY2ZSqGWsRJrF+KCdyzZOdXJgNYO25paZCdR1SOV8r+/hX
jQInFWCzLnPU4F3d5MRwI7ZI1AFVp6FMUpHP+TWx86W0GeJEYiUtK3umsexC+FW/
5ipdWNSyBX9KzDLQ5Sg75wHmsR3IAnqX2loE5fp0mHlrpZ14TdjjUpyTCAXxg8qM
7RY2I/ai/5JQIaHZcWZ4SICcbZxz0/IrDCuyrnYb/sBFRhoboIcNLfSway5hKCWN
PVD0XY5dlsNi85armj3F8mzyBkG5jmgwi7kcHNENBxDCYRk58P8EsopUKKAyPXpZ
EYHxbNPkgQsjJGP5A/WsNi55A2ABexh+5RE6iyIa0rO9t4kSKwDE5W6YCK9Ey7OH
iDld2pPqMsPoKtmw1Lwoj6bv5k3RwVSLLve2F++KNcuQedCkIJgfDhpQJ4Xbjs0T
AwHOZ2L5JViOT/RIFmN4INrtSWaZ6iR3bQ0Boo+i+lCqff+55HuRlyIwg/uAv3sy
NUolEXVQe4hhtKH8Q6EA3kstoZyAcPxWVP/F9UZnnrJlnjnWNitl+JCFxXNV96Tm
c3El54OrE9E1WLBJMuKI4ZYX2r+WDoKyJQZZ7WRfEQuCSqM2FfPmlFMDcK/Zta2X
jOy+XMBjoZxhJghZw4U/4ovnos93PdF4lEvwqJRhQQtep/P692/LC3bGokL9wAiG
fzKsYkI6fhdVJmzKrZ33mbNb8RX++EE9oxMMP1dDb6ilaOG6/4poT97SDwEF4+x4
3JMfk1TMck6DIkoTFENrnPiYVfFP0+zmIACgYclYwb/LH2H1NfLQ1vdEtI+BdxSI
gC2UNeYAPiACg98ybH6YsipkQHKXMsM6PxUMmESyCCAVkEvikMWHvzRdla3VuMw3
ofnI4fKPxgCvnOdvjtqx+gYTyYuVVdKMy+FzcUqzG6g69C/hKTxRM/ROCI+jawKI
IcH17NxZV8icx3OKQ4U3iG3k+xcYITKK/zfRoBZ/VDOIRPoMadlsMg3wmkbABgMJ
45nwNoRzCD7DBUMtimRhIz0xnXowB+VibuUv9q3x/TkJOpJd8sCqmrudPU90CCKv
TwQJ6XZV8MzrnaNOkebcwGhOw/+2H/Uhz4/aA5BKQyCx5vHZw4xbQh9Lm5F81a6T
6D0kbW3ELYxhgkzONK/hvoYQ2t894JlLeR6QFGRN6Puixg5DZR0dipB4NjI6+tk0
eP7F6WzGRB0AhPXLCX8N3ladR3nNs/gi54CrgUCxmPPL9DtogNE5Yzk5Z9S5s10u
0LoUAMTAYdG1dkuHdj1oVBQ5p02vV3ysNhU+rZo3gBYlc6y01fK0ZX5ho3uMYEaW
D4cU1W4M54o0qGER54Xly/JfgZEA4jZUEBsKZc3D0Sc8mGe46VgaaHYDC/EvrtSF
fp6HO3nmHLpL6dT7SvIY1sXiVJ5n8p12H8VV89mS+PLsZhKPGyfgK9zSj4pTCH5t
JyvYClpQ9u1gQEmmaj+L14eq/VdQ9ZGJv5aE8grP2UTBnK6Y+eEK9mrQhN222v2R
lfKZvm0YyiOjiXX83TpkaOBE+8WJ5CS9mLX/2BcFZDbt/0Ec6Il4+iUIn1z3Onk+
Tm4zy+tT/GhHPtyrztWNZwPbgZb1xMFGIAAIoRWIE8I82D248Vt3ZDfgsy/h1Py5
l9M5+2kXn+sj4hktIRcZFB/WrISo11GgLWKim6k1E/CclT0obndYTBC50/pWHyx4
+/oAMtfcIf2yQt2yr42ZTD4/Exi5LhQEgQV/QftQkcfZzf16J6Y0fExh5AW7pLJF
bV4/FLEtPJ8kMZf37+nfe2v9RFL7STKl1G50z7Da27Z80686ftgSB/l8KxGv4EVX
UECmWRPByEqZXDoVh2JW7rUpwCU7dmVmmksqQQYCMDssN03+BJwsgdet6ZNIRJud
S2Hr4N0FQeJRF8SzoWVDafDt4B30f57qMGC7ISjbEtcmfYE1D3HuESnu4ibqPjPv
aDOsbOi7Ee2h8BQbdswJHYxAZ0D2YOirjYg7z6TIOWLNzUnMh9aQr1ddGgseuOkv
paaN0NhvKdOvAhjyEWscosJ6VmcoZefWTH1qCXMp1qsq5WBptkXtca4/D3LkJIQ4
LDxVQBPo8m3Mz7U4A9MidVEX78YFFgr0hnePjkD0rI6rDnv4lL3Mp8oPfcehTQD8
j+3sP5FVPzEq0CKXoXfZkTJriiBWaHXHr9WdReGf7XwwTr9KbHKMfSZbv+MetLNp
tbj2wMqV0tHHvC1bmW/ZzbKhJ8e8OuLf6aXtVSmmiBDgbs50zENdftsRxfKQBNF+
zoLXv0jm9wNT/tIRG/36+5uQGur3NCPiZG4CWPgho9Qcfs95CKFDDDnQNYMAefoY
sHNCeZmNRZkCawimFKfbHojGgotJz19okPwisZ1tbKYwGxJ5yf8p22xn4Y8Lzw2j
zQRRsKrEjX/zCpBi7UFcbv9deHuqjX5uLyoBgvF9Rz5k+lzwjIsJ3KxKW1TDp1z7
kMCrRJ/wHGNUMOAPY7Xf0TOBgT7poPEb131abeL4fjcUah97X0hgeCnAPqm3GHFu
aRgTY6daEBKARgmCNwmWgyGEZdu9qMI4FJEeC8kCFrFDPhfG/j82VeFHDs/9YdXm
2/x+0vMULNxsM7gIDVpctGsBRxSKsovJ7s9SEaC8ZZ/NVHu3VuH9OTAI9Rnqbj09
U3l6CEv+mTSVSsPX3slzph2eNVQv4bUbvidVPGFxTVfsyBKu00VW26YE8sBmWYp1
yoydJnf7nnAoF/x9Y34izVlft0vpa+oryk3iKbp7SHnC635MiAUIc7tPYIz9S0P+
BZDtNNlyRrtTMFK+qeJPSVSkwjaOfL7h7MqG3HZmPj8bl5CqvP8HTUozFGkTAZXr
JCgjKSDus0afnQQK/Ld1h1hDLMtvEEjikkN/uwSxL+tnKlC38uO/+mCFBG3VTdmW
vbcpRI90BtbaLWI2qR1zik8vxG/+UH8J9d/0EkvJAIRC7nQerBNAAEqJPlSlleA/
E8vkAy2gT/4mczMTid6tZQdqWrEJMMdLBO/tzpqV1yKr47fWUbXiqTEH5KRjkcS0
Fsz0iv8Gr1sjKWa75LrgaIoBXadSvWqPiuuFumzhkwWZAQgEqgM3RSg5xNVeHusD
ITM+Rv27oaJQI5WFEvAQ0Gw0T5Kuhp37bT+0ZBiotbObauAiMcSXC70Fk8gY1q+R
glGW3zjbxgQJT20FJ5oej4NK1mPabcR7ffh4yShoWCZ2xhyI661+n4dUGdpuY6ef
ZZcRrHNfA9HY8xT+ONhvwOzUvQZgeiB5SRRyuY5CLcCbsfTDfM8bUOD1XqhyDy58
HbxDr38JxrWjLg4iBnd6V02bEmjIP1RygDe+mzErm27zq13o8DGYI3QNKdA9Vg3b
obYAq5Ba6kmkha4lB2a8zT0nmXXDpq0wYeWWdbjTeyq53y5/mM9eZL1c6TU8lGL+
p8MUp/wc7+ClNmaqYXVS2fhYoeshjTdKtW++v+vkJtD4BeUHvAr9fqr9hw1ktZ7F
6g49fuiympuDYJCHjC3rT9e9bIUHo/zv5P6nUr8LE6jjrfo/wVhn0V3bxoRWB0zK
Q4rkcxy6+IpIYMqZR4AOjCJg8huAdejq0SDENqxwuINAgud3gMhCk6BDgEXQ8hTg
t4SDsDjXnGJ5S8ADLtjJ/hMUQTysSpEfQR5CCRsb20R7jU0YPckgA954vqoy7cZE
v6HGKOzbQoyJRoilDYv+XSBAk2d/tEQxedhUmY9nBxQe3EXrVXLpvSn6Seo27lcf
ke7Ppx2tXU/lBEWn14fWyTkfit9PKMXxhUebYQZm+Z+1RqvLk5ria7P7Q8PK8rE2
r/Hzhd+9+HM+xduU054MaKY5WEqQ/DhqvKYBEjvy5iNLllFqD6A6boje5M5M9kGA
saU9pd6gU/AuJ/p+azMIejBjAzAwJnKrso7wcVvU359uoR3e+HK4S5/qjeI6JEhE
wKP9VCwc/CpjWvL4Ns4YOJpuX/Qa99lSP+aWZrhwierQFsLqQ2kXKOpluc3Kxwlb
3LQHiJOe5WQQZAQb7QLInCTr4nvTGENp8Ne9XHo7E1HQ4V0hTzCn50MPSfvc4X9J
86FCGVADvzrYypz9GyBMB15gTa5SwZmmZO1+MvsyVjQB9r6ZITFXbiAEISHZaDwU
uWotoefAvs1yXXqDZ53TaXJWys4RVN4iIx/5IrPP2BIZmu1769RuXqBn/Q2xVdZ9
xp9OT168mI9hJDxSG6zo4b+jslsecrk32NI6djOuGYNAbJ3EHT9oOatH0az3dbDh
KEEetGTXgkyvS1OB4+aY+5PX4YkerIH/rik00nrk60cIgFRwTSWAVC6oeBVcVz38
y4CL99dXCMojBC8TQe9eb/Vu+IqpvPWmFvrY6bj10fj8Nnp9HR8Aq4nhq0abR1bX
EUpWjpVO1fFZOTS+HtI1eXLEJSLvlFhG0odUlxc9q3i/N7sV+Gy3Y1h6GPLJYbXg
od+dwjXvDNZ38ZsGBM3tkVuDnfR+IpyVNapdhpb1lCvH+d6BSVynCIvR/x3RTXgk
PJanUK32r+WZrsHoITzm+8++cdT3zvPcuJ9EDVEXcAVQ1RfMk4r/OyDxnBvB4ni+
PH/HVrk4LYrCfo45ZfkbJxA62hp+UiAQKe7sBQDs2O7w+JiDlusxiD+04edh8a/D
MvXClScKh/vk0V3G6paFDYxMsQWO3VcTBKqZgUAFZ+gLdeZqFaBU6pQ9Vk0TuHMj
YQQB44WUtvJH2fxMm0CsJk4V8ty5xLrp3kGZmNTwQECRAArL5V2EUxJ2ha8Fudy5
ayQECS1dJInqbsDfnkhJuBoQmRzSummarWZhgoQenwKDiJIbWcUu2XLNwwfRovpH
77lHuJE4Mf9NGvxOGiS3WYmsvCoEW9OuWo7bZoUDHW0rISbAjn5rx/RDzUwQ+A5F
pXRNBuhY+lP6EFoporZgRKb7N/6ztYOYamloOABQEgLh3BK9pNqchpQU4T1ECeGj
T7MC5GwHVxt2VsXk6MPnovvgaFMbp6/qzSNc+g3So8hYiiCBDQfBOyDuQD9CPSLr
CSAaDECLvnZy3SyBkm5Vb0y9epOH2kyFYTLIsmMI5+jejyWhlv4Y7eb+tXAGpI6f
aloiBXhEcj14Du4kmq/Cja8gqRNTIPcB5RePvM0lDks5TDV2ioPXy+zAcZh0EOvb
+DahCndUyG4tkBSmmpTM9ccopUmQnerajDDsj47+yv0WH2HmVjUK6iPn03PzxFBs
OMIW0Zaw+FMk9Xn0//qGfS4BGEGYG0FvokiMktDmMlZYGTkdwMjNaTTixv/PzSYx
XrLiqmM18t86tJppY2aacu94u9cv6ebkr7EUzxa6iYF4AMVzRfhhxNS5dWc6SBaS
SpB7RJmLY+uvWqTdVQevA7xwyEZHYpny9V9/h3atdKBDayGjZ8UmcbH5cP0DHB36
ubdsvS5DQv1UyJlKpIw1gQfJOrXOyRqg/AYj2fRzdHdPggj3q4YErsShCJvRM3ni
Er2lCf+h1x3hfmV2Gmc4SdQMHN7TEaJoJ7j+/qwmZ0wYIg9jhSAwA3eauoxl1x42
84S+E+4TpRaF2U/FJT+5i2qk3rO3A5WjJg7WYdNCMyx2VG9+wWtLR+Crbwy22IuB
TiYRyrjCigm3JO5dESV0JYYc1JAnelqcRg0yy+x1HHO0RVoYLn+cpaZQmH3Cd4ju
8R7Irou4JGsH6xhD5V19EPDdBH8wg4xILPQSn47sISxIlAN1Q/Fiov3IWFj665T4
qGZ8GrCzZpu1sXRLCO4v5hNJobxwsbGflBna9spbL7CcTxQw7w9PiDhqQMunHWop
eRjmevR699/yLJLThZZk+xl+9Zjp3wpIUstUMnddJUj/5Ek59KTgAemfkUQsT5pz
aJCEivx+jZA0FHvSMz35m0L0lV6KvvFHQs6SMIW2bpMD9XhVxqMVG4WgAvRnL1vO
GzMrxNZEU1qEpkGiosEOwfv7MviSkN7Ys7nXhCjhEioCOOn9Dla0rMaJpqpNXpZo
cdrxUFICQVNFFScJLtlm+ourYYHGJo62IvaW8tv3LDIBUrn9usuQrzXukGomUZYD
m733UDNA3BxdHedrJdB4hYHNef3tfkG+hC+DxZr0zIgxVUB6CXNcjDBh676H30kO
2w1YXaqfedIw0nTQthMgEnmpYMjVK4/iL56q2RNfXSoW4+6R9fn2LvzIqU93f+JZ
AMYWX4ZW2v9qaKcSoARL8dn2Lv8kfLJRp4iHgZeyHowRgHGup3oNi2LvYWboc3ic
iOUdIKTCzgi4/dM0zxyyjGujeCB/agufPdwDG8JB7dcwUypNhZ+JaU6j4yz+yX2W
8lyIKDkgNMN2ash/rtl/DI7KLBbCGAjvf+mKdXZV1vQboBCj6rXGNjy59SJk69os
0yySXFAJJi5swIV5uXE7w29276iSWvvOM/uK3r38H8HJYzVHrmHFgMU6XWSVCyV3
1OpM+pr6NaPfNqtq+hNgdvaZsbWhwsywOnAapkfckBIOnYB0EoLcDj2ZkuUgMU33
QEyh1e7e6DiTrPvuXhUT/Tuu8klr9dFlqR1jYRLd/T1W9BXoWyNcYQ4G2KTmdM+G
qoDMTDJMDNe+14BKyj9r0HAV6S0iofGx8+5XBRye5/gv5P02GHG3ycOeOj+5OGGl
9M+JSLg/HhDZX1bYUpqab8cTp+CZl4+daOpZtdrsdE7uGRgg3wjIATE0cGwY3moU
c+vz93RwC66bdxw5SO5u++3SFTLxBIWzdM1xOnkp/jZCfXo4344LfmKFAf+KwV+o
tOBq3ucG6IbsNxObgnNAeZ5g/IKhS9dTQBAFwy/3zsl6sZUeCMPZOQ97VGuCRa24
aDpmqYt+p41YWpVslLbPzEhFv/GHc1IJZPvh6/N2fnhNJ+fKYclfOAXVqKOEOhLV
UDS053ZaZFatb0NE0Hnn0Q5DNmgtALQ1Jz6MIMiTeirypI/bVQMLpqwnFWnvnApx
lui5I8q9bimvZaFZTOV0dpoUiC+Xm+Py2LfRzY7TmEnoXNcgvREnWgp0KZOiwB5J
cAMtiIcH0GjNvLzvktrg9a0IhIT1GNefUJEVAYo4UBblBYxptWQf/qpOPpq6jkDa
47rR21tOQ9B+KG/JfGME5GekI99uHjP0rDwBltns1XMSCin1DBfTA7WaXShs/N7B
AkGKDfQZSZItUrf6M4HIX5upUwBkh7v/b1x9XjbdXWLzKX47hFw+lhPmidkZPk4u
vK8jD77bsrf5G+Y8jPt6vObA119a5AI76pIjTN8t0mmsg0yLNgM6YgwRYy6fU25X
Aw8Ji0zaRjV5uWt7+bda18qFbwOLBHF6cOSP1rLtkun0OV/l/5f10uuZqfRrpyVN
PLHzUFtLfaA8/4hKlkp2uvDD7kWVoLDXEJOD+ZRJsKpdGeRNU9Lv2sCEnpCOl/zZ
W6DYlgm3e6FK6/AuqF4I8xRA1e/GC6zifgEW+mn4rQRGtzyAh0itDvOyXn13g48Z
chxa99NOJNUpVCYVqKSmLLx6TMLykvK9UrHV1G8bwbnSJC2g5mYKmwTXrGBfU6L0
k3yYgpHFTyLlUeCfkbRjTj9/SSg1gpGY5pg06P5P9SJOzaq/3ATqOzRXN7nJzgGU
mXVUUPpHUO/pvfoZC0qXrRDZ7p4hMyGupbYgy7pqAXIIiyBTbCTc6V00no+1XCWS
TmES9On/NywLVW7iarqJfU0/8Wfhw4dDmDruBIzaZpu19p69moTVYLL92cIHzkup
UHd7xqPAo2fQdXYDgx+GGLEBVI8qUGtvIEzcbqFQ4/C5Fq2ppGbHYrpfT3+EZn/u
HWOREc3ta7vjoMxTLtqKK0UFi6CfgUmk36DPtrT/BYaMM+0p4IHb5NofJZI+FdnQ
T7vnC2zSS1Hqr8cPRhqqOm3wltEmZ86GRx7eZoyrden+iZBcWRX4zGWlOTfaQgbQ
rRSiEDfWtjn2mUe25S7VNJfaeuypRvv+59grENdNSIKIU0KW4XAU+np9jElM7QjY
3TB21H4Syzux/N34P5ESr2c2TGEqo+8RFc9V7V2/PAlSIrN1KLtQVw113PfcFClZ
KLOiRrOU9qvEowHQvIlULe7GYVqjNhOxQkjYamgLiiDsoG3XOvzkZDX9CHgAdbSL
KF5WyzpHPjglnRVz1kW27cs9/fwNKXAA6h925WQ3r6DSa8XAuRQRWQyJCEwb4IZQ
75lzRgp952S/46qHpEIxChy8S6lzi2aP7NJWXtmh8jd4mcP0NJPxxx5Vbqqe42w9
422DDVYPO6BErxx0q3aEV4ASTGQqhX70KRyjsWUVQvo4ysZHVfIdAyPl0Vf7hSGb
ZMKrN4WIXdrMjGcAQIWGnXTpDgzkgyLuJLq4FFyJ+a+d7xi8cGdUZ5PVrNXV169s
oUsLpczM35FZbBrviaQxMGWjfS3IvDtD8jMsg4a1aDZr4SLbYKEDczyAHvwSs7dt
nK6T2KS5TLhnW77i+ulCxrlL7O7EuJ+m4BKci/MogplT/d+NcAX/gfPqVqEDODSv
MTRgga9wa0gOjyljKJ2+022uAkTCcE0N+wDtIUDTifO5t+hedtAqRHS8+a1KWegO
igQgCf+lOkNMgcA73pN/+njpHER3eoDTxVhLPONVRQODe89Fk6nU2m+1Ygj+cFx8
t5AIAGKoCGeWYZXfmjtXvSv4n53b/fuGLgu/ibUdS54qL3cmSeHGgFc37v4Ot0it
UWGy6rUBffoeGjSZPZFAUvdLu3v+L/ttDndKDfm1CTdiYzKanXXtB5WCECdLf+0Y
1LLHM47djZkodbJ3pu4rM1tEvwj8MQcH8+gdZ4u67S2BAdtl3iadE5lrQdTOnGTH
aWV7rIK6Rbb5dF9ADs9cu+uVCX/Hw3Z7g6nKnrYKmg2YSx9Utalnqj0LO4BOjcJJ
hXwomjFvgfAIubz0leOVnn8IMGEKN4EKB1xMf92AafogJei3rX5UCYdNYyNaxnGp
WBK9MwRwWrt/uFOoDWsxV9E7WnPLZUOUWzl4bOeU2NLoB29cMF8+P3drC5Zn3sw0
D64vkL9JwSTDLzqyZUs15RyqYG5EdjQstbujPae8KgPlIfSbuftstBaRN8gjAAVE
XvawMqiPmiwZNdAG7dhhs8umKUv66UMSFSRHdRyOyHVGXoPLC0Tp+fFDzNCoBLh7
Qoz8Vf7Y+3436UiPFtnYd3ecaPEIe1d2X7j1RqxKKVjcep5IA1GYFotZlrqkZlgg
/4fK72eIS7ICE+0fT029F6xT2lk1XBHFNpHocwKKtZpk9RPBZgbVwoVkZCRgkoWm
4MWDrG69D98E3dYn46J/WFYXIhtHNrf5erSJgmehNIMZFKfO5mpEAeq+FcC66LK5
8aD9Uy3DI7+3ALmKT6Kt5Aymr6HOEQjowNxyi3cW+Fi4wx8siEageyUT0VG45ZTy
wOqsLZ8RywaW2FJ1FTC6uoyYyJ5I58EwpgPXl7Mx6irPKkvs7x9qA0G7n5m81XY6
6zshMUzMoMYvCcMBSmryZCcYm2JjJInIAwCX7AyoW7q2qAmQ436LFeDwSMNmvLnm
plURHBq9/nTEHQMoNsBVGaqXaj6qMXfynY/AmhjhPgs/9h/NectmU0TJ5C6PIjg0
Aq19y5Yq58ooRK2PQvtHvXZ/18TBFAeqJchrPX6u0E5GLNPfLNggC3zygBZ8xj2G
lRv9ax/5dteQi5BNfrdNXplxWS8khhoFDZweHLFmRAQoq+ZB/776KiAZ4W/QUNr6
1fccwQzqybFLqcrSm3U5rKDcITZzCgQXRnTv4KYR7P9QYp0RyxrRTq6y1aIDyHQT
VvgG55fgbkN6tboXpZhbeXCUaCFm0mReJMSQlLRai2mlKrSgjdPGdOsRzBLW/R/2
4YaPxtKWgO6rBAIrZg+Xh00Rk42Y0o6g7Q8PSz3/nRCNWV8G+OdNvjrAJGyw2Ohr
PovrcHE9HaXrKRltLtGQ9eQq4qjD5EognCXCZR/p3swFUitJO+xoE+llU7IYF2bM
DmIweSMGM9Z72OxlXlFk170XjUV5+ycC7432AvQDU4SZgl/I825Wx/340WZNG9ZA
Vgh0wA7tivPjLV9LO0vt4y7E35ykizo+RY6fAKoeYkLod/DMRwzhw6bwYqyP0Fk6
muOvDK7PvRhjyCaZZ9h047IWClEf8ibR+gIyzdZzL2RKwcoPuBQlCyfCTWfQPFRS
3aX915FROqjUQgBYsDIu6eW/TnEiOI9rYN0qLWdTP8UEPrqnOZGZFvuvs0BkKbWV
IDm4Wxo0PNk2UWnpGBMmDY0N7do/xjScwEf9VAvfGE/jXJChhZWPNwC3PCUKmyy0
7AilvgiWI6X4bxrNt+AMGx5RBZUflhx8BXmybWihuULRAcq4ffgkj4vsyVTDWB6v
2WU+cEj+Wde1+tFtzL6VZR8HmjN/gkYx+07K+k88A33jXZm7g1zlbyxWL168vzPg
f8xQQJJmPN4AvwobjcfahholgtH8J3XgKrvEtKi5ZMjfBcW7So3wiiiyPoKStHOr
wy7Ycybc8+YLGwhEGZwPVAaU6sBUPHNe44BkbvPrUUQWkc6kAsW2JaMaK2N6rajQ
+Ny+mcWTTDq52ezzcjTWl4HYF1Wf11BqToBawlewD4JZXjZ+e+toKC7iBGEJFXUc
vqSloX6nYxqYZbU7I+qZXJg8OxeAElw0l3BYn/QyfxVnhw2ymDAzll8TfTNn4kmp
DQ7nzdGSN+SpFUvwHiTz4JWjckJMMeRolA9kKGo2c2R9/TjeztaoxSgGSZXr6Y0z
WHe32Tml20i2iyvbpKM6IK/K8NH+KXxYr1l/1A2ZqSZ0UE6bAWnkK/Pc8tL/FUYw
uaMl65jAlWVjK1YnqLjgbjZi+392GpOQmGc1EqsBj1FZnBgBY8uIJcg304V67nc9
4Gse0qTWIVIFsEfjX9QwR6dL+uxv7KOfJbJ0YCo8BVLqX1OW/V11OgbZVOuulhyf
5WEBmHxQLNih6PyB570NrRync/rx8QO8yDXYIpXJNq/RDTc9NoVAOkTivXVsE+Iu
w4vKJQH3DV6WoOW6DbsIz3+FIdIZQlwO6n64lFaXxGvYxAjmXs+2C6DzNyGnI67c
U7xeZNryq6z8JduFo10j6LGBrfCjrb+JZqJNjwUAtTpnLnlcsnRwwN4UEGZnaX9F
1N0JSsq/+tyEUmjR5Oi2IjBT5NItNd4vHueSXj4uUL8ZBYi+CYMoDNs3vJe0ryXh
LH8VHAOpfqZTJj1b7J00Fxh3+Wwr/BTpyt4v2A2t2vzaOH+7QUKSPwcYXu4fsb+A
EohFrdToqxduOGj/2Cj/BZtmBokvT7/TLFxv7y6FKR2YWv/nsTOshaGvXCSXjGZ3
xik9/t6bvynEnI6rOksjzyfaK+APp2AaKm68QSj59wPvq7p4B9UJ7VxaDXeQ/rBi
Kz590wCoJwK6fyvorS3Y/bvGi6Ho7OIF1P+a0fsJppKVOg+fOJBFpz6+YNZJSJbQ
LehygUQZQLJYWqOUqOX10lOkbwkvyIFIw46/x/B7fsowjLpOSKR8JFlybk7eRHZY
8FoiT3QwYPtJlr2aOAD5hcKsWlv4IlyB6Afr5xfaV9V1aYxJ0NPH1L+GaO7gLFNg
d1oINxK3pfkkPQn1ZKlLiB4UrnDk0OsWkwe7rJ4nzK1jcGGjk3nOcBPGQJx6YYHH
SAuSY6HwR9lVtAsmA//XdHrL6yi1D/L5x7HeollMJ+s/O7BYNPBU/sXq3cXKl8Ix
6XAQK/El923oyMd/U7hmKS6//8+xwUkl/yICPe9vDxcepH+2UnPHZ4hfm5QWi+8/
ZJPLvYtrGn76WYDlrA6WHn0JgkFl+tPoK/afFlGSKc88tlCxx1QHRu3KQd0n9iO7
p7xhhiW/dWGn2wyIGTjSUxRR/ZGhS4giHTKt0g2ZzUwVsS5OStTeUXK0P+Lnx1MV
Vyr4ksE8X/Vg/45YE6XFkJUPYnvh8R8XrZR5DJOK+Pdm2bdjk8B1CleROhu/rLG7
HtRTkeccMNlC0sg9MXHomBYwuEypv2T4EPm3AUH2aEJ5UL9TwVCGYElYX1M3JsHE
q8mI89QvWkS3jdZmaF0OnW8QbaJ4xCBF5bpvTizBWS9nFm089HmOurbSPJTQCZ6E
qMM0W3H/UdW1Waep3HXk4Jxp15mn33MtXYPQmi5/HZmmzY0L4mNGttqbUf/xNV7N
We6+QxHrpPXAqX81lztTL3rq6CrMnPfwFXf40RA+zV3GsMMKajrG0bHLS0WYaB1g
lg1kJmA7SANQ9wpZCiBSuAFg6z2TUQoBv2Tm+CVfqU6XCwoo9H4AEm9lxY74fDzQ
JAwfqLNJIgG258EhMbgaQu1kQSy1YwiKP0vjOmCZsrns5Y1GdOGdsevkQhn4WGkR
NoaPuEnRvk+3G69CkrGCWQTqt1GzTP6JFwIa1vHpmPeEnszU3byy5YtOC4qz7+nj
lXg0zPrUlqN67r94YMb3Lhct5wt4uXBfCBo6wrdIX124uxeLD05gklE9C7ajuonD
HddqHBI/TM/UqOXbR3IpRkLZ0Ecn0AS2sWcpWCBK1jm3JqJmDIZ8EueR0uiH6k0J
F3F8JJAwIU68voi/NrC9BkRP9s0rGbEtEetjUrXl1bfo6Bms6FmJU0rhpFA3cun3
v3qL90oh469gEPJfDlJpKK6VEdOYEvwBN6d/XKjkZbhRKuO3cG9tNXYdUqMpwS48
GDnie0E301em3VXivQ0AKhnhWH+Ts6L8DZgm4aaCFNgK+kjV48TDWD/IufMqm749
LeUEEfY/eDubRhO/UgAMLu8R0LKiRSPIhR6tW47D+V9uonqOiyPz2Uo37WaaDNM1
KDVnQWefHoMuS5+LfIGniwnTGvvnVQd5Gxh2R6B5jBbGYKc0MmEwR+9NI4LfTnyX
7DVfwXOqby+g7bn5zEm6r4gFfSIl7vlsWdXDfeLb7MzMoY6ghdyRKu8Az2cZPhMD
6k7GIs4LS7MxE2xfLDNyr49DouMaQRD60d0NYMddtu2AEmrjJBZPzs85qww/lQ5h
Zm3S8bPTrr+xFmO6B+Z2TdwLRdqiQ0fEXQFwHvq8CbA0D986XAMIp7t0nywcmWQx
VHWKV2QkbjlV2/4j+3tC3jUTQdLJFI+TVwHfyA+F2o/BcNuABr3dcsN6PnGuLbFw
eG8di/PCM0MukBJezDrTEwBG7UI1Gd/ccPAfpt4s3ZbMZ1gowrjenFxQT/P4gDdJ
7THIbPsJ0wkjaVU5gtEQFjoeAx4SQ4Ms8pJ/MmWdkQa4S+4SEvBN2ZvGV4Qa5hqO
BrAK3cB2bJkr5Kzi+Cht/vQIdzFTNxkgwTi7jWXzRoC6Yhv01vIatmY5oWv2E85V
S9ZBYB1Prm/EdRiNPangeGKd2KzM0C3KbN8U4C482Qr4DLhBijg8/QA8gAq+ugdO
OsSySt3GfxtZ1C1HmquCl80mKn1hitKLi/QFS95HfBXyf/d0Rifckb+FdL3cy9HC
CDZWhqaz56kxFFPg2sSiqNoBZryHMOvcCTl8us3GmdE69m+Z3tW7uPDAt14lTJkY
VVmusEg7uYJ9uP04g33RVV+vERlM/5ob4HymEmWdG5Z5I4rbSsbI8llW5E8Ykc7+
wQCN+WAwEDBhBjMFqm2T7nqYX+91v9Q/QSPtBUForDqXEVK/32+noPQN+hu6MYro
cQjaB1eDuhkkngmJCoQ/sshYFImRWq5NKmbcmVb4X4X8eY9CiLlpVW1yNSVAsJ2Z
CfbTaNQ7wqkRWfFGHsfLjrsjdzjttPFJRCmUNVHFBmEbo/yfP2u+q+VLGRlXkHH8
h5ZFpKhUBARFs0CJMvQ7e4alf6bNI4KD9gs1x2LQweSIVez02tDGAA6huIIxWNxl
cT+OcvOYHvzco2OJXdHruywkWKPE3l0lJZ7A7/SgW5AENsrvdaxEizr7b9bl1G6U
rCgnlUFVfCtCMUjZEp9I01+2f5yiABSe4h3qMgv/mLLS0ep7TFatWUQ7sptRnmG/
Ar/sPY97dC+eaAoyiNmHO/INt2L3nID+66SS5ESTJzgtkIec/TYsD5VR4HSnZWEb
Y8eAGyb/0K+4vr6bHx3kgkFb1+nTMcCf/HS3QezkEfqFHnlOlnEowGIC7CgkNx83
CkX3/tCFV9wW6ws1QAfuk8x6PUINBn4hHI1IgSAsWZERhJwTl5+n7581QnrvVuEw
uA4ckOcjnd078Ie/tjRQ9JdjcqffaAuCxBEwrFkD9+ufY4CXMxASzhjVmp0JtuDm
TJZTV9GWDx4oSEqfn2Ev+ZIiBoMzDeXoyNigzwdR71iz/MrA+uCZu1GHTaVpC95/
3SKJew2/klzS7SDSCrNzCku4pnYzHNDASWM/ye3Xz3INVQqwuUA977XAvdafUtFu
maIoF4iKBsfwSYr3ardYki48kv02X+R9Pv8FQDMnD7/4YFJKZFRS2gPa5i9xN8wg
3jb3by4xilsAqX3IMxezqTkSEP6YgcPB1Nn+zCHTdDb04LDSw1XHctaA+wGTIS18
ktedDMOeRBikrKsCF7jINIct8I3rYnVT8i1x5JCrWbOt/wWJ34qOmrQB9LtSsQIo
b0H60Z1Q9jvNeLzS8uJi85HZGJRzGLlLuwGC/7sZ8YGQrwzpJosNZUxGA2A2SkAD
y0AeWIGJvi+WMgZJ9noNVecb0EXnHzB3Fk7o2arY4aUFcxoAhm43K9QtpbjCiCEm
WWxoUEyt3LJvcIJruXmzPWMZUhJ4TBXwbIbhh4OLr2DLfNjftx3nWKG4gxIKrh54
ilbjZ19KLTam+nhKG3ePSbiMd+iE3U+WbrMTMRvt6zCbRt+U3jaw65heT+rp+vUG
k9ZBwSEpoar2SZf94fBNv39nS2A5fykGpKO7Isth4PC+Px9ZOWPs+GK68DP5FBB4
kArYitmYN6ZwelGodPdHN8QRUkt/r+gb3JvllppOC4LZsmWZLWPWmSD1c9PNdlQ2
xuZn+TQesmG3gCxFFCTqK6HSYPV88dEUex3wrL0o+0N7bwWKwQTXcQyBOvnCOoLC
xo/8Jsm+JmmfgUIngdK08JBwZlOh4gnWzMVwUpEjI9gkDw+vaqvbHRJhP2G7dATn
eMOIP/qZMk1v0ecKNphB6IAB4fTgH4XkuNi6plnjDoX2XFJNSIyGptxJc1ZwAnsA
XFDOkuG049wce1YpCgZdenhzTIL+gbmIsEnLrB0PF5l0+EbfgbdmjrBonC6dR7z9
A15fzKW1cvHbNO/cXJFkyad0o8s6rpqKVn+p+oMbvcd5hSEihSnUfEN+HuTGUaop
PB1tZdyYvFFyshBm+TiX2Dd2xdyPKNfi7K0WOj3z4rnzTfycPlOxt9ql/sdBeQ7K
WqOiZ5cb9KKruC1DfaaBm5l714Qk7jIvf2Ql1N10qgz15bx7gZOpFBNUBLpZqpbt
tzJgh6D6SaxiQzCyGXw/tHV8vztS3XpduIkWs6WYwAawf1btnF+laUrLWPkp+PTa
yC1X1f+IBUYJT8+E+K/GTOWWQc6m2eOy3nO0MSW5K9uQ3/h3bYnZVbPnN4kBKibA
dgSHvFsoyrOfcEtQMgEujug7VVi0RDxBQY15sOqdUdATB5LHVA1hLpNlGi/pr9vF
B3Vr3/zd3VUlfVJuYgrylGdEu1d5mul+HQV4P+S8rLpyI1P85GZw89zTKurlk4m9
vB7pryOTapl9WabwZOUzYNxquWpA/qrMl/ZvxoIT97EQ+bF1EIJQTW1TVDf7N1Xk
oOE9+W3V7Uifb2+sgqX+d8RWwiyOGu4WueSMG3h5B05Cn59knTtP/PU0dr7oBscj
EWs50GRn7XYe55WppWVPLdJAJ+rpJNKP2nKkplUwGqyK5QJVlpXTz9NvMzqchZmW
6DYuvgmycR3+hqwjwicD4kshmyKzkaSfz2XPF3qTEg0wPbNq/H2lEAl3KYTzQ4+E
xkcKfYJbKDOnuKE+prCin7oWMcil42R0R+jOj5u4ehf0sZarSj/EhI8Bj9DeTHp2
3IcpEANeqIQggXNX7kAVV8nByo/CSALKD/T3kOuw90iH4eQXdxHC4/PbS57EurGq
OLZjA4R58h0QxVQCdp75n1pXx1+XTaZ57heIkY/IFP/nKg8GLTzDhkT7Zt17tUM6
aXBMSUpwiQcTImBGHswNDZD8yju9QDKRo6LMxA/7mRws5KpkC+2w4feLORmtEYp/
oV/L+hQwv9N3AToGA3wooV0CCZpLS9ojgrm2QbgiReS3yMZUahyZK9pINYCp3GvA
m7wCPMFvgr/dhnMFkBajFXPYxJmgQYnYWTansgRDQ4HjNC6a/YG1jvVGwLp+nbCP
1UnB+qjGj6utLtU8EUqzwq2RFw5FiIG/ybyAMeve0kt+FrtBkhpmtNmjNwYI/2we
ii4n5VKbFmRAtaIEA3pcnrxTGnZcosG9XHfb4NxdIoeA2oKAO2JmbaXgBgkcou0t
78TInVfAEYkW4Pkrt6fOkcut0APpRK18xTUzo+CzvkZL2Vs16nGDU6V4ft9hEBC0
tXNstDkRv6mNNmJC+nkY91aFPmGTCqBoQE8ZlS3/DRQpBHqFjsFInK7tjQJcxkD/
FF/glANbgJsLIz1y1s9z6uL1viEQb3LZPqYkFmRtpoH2EQL9gc30MPIZ3s9jILBd
NfNRmik9SsMhXRFleKNx3VMR94eeHuujYzvuxVpBV0GiZJjfaB6xTTIGniQtcMau
uc2WUYLGDtZnjfpgpenR91IAWBhjd79qyWY0hm7nXtGpbHDw+7FEygHE8SCQwjKk
3Cl5/xf25L4kf7x4iE69WGlfx+3a/6RXXjSk38j33/9R6tSEaOuco8on7wI9t6fS
EBTkmiHZNbrNESFyf8xnFFSE9M8UKGL/mKd7zFIHQBbUoxv/CToIHSu4ZXhTXhXD
XMter7RjWwLe2rPRTegX46VmAeC1+jyY+ocgEucMsjbbnbF/CJFiumdxEwQ7Ay/P
MFPkatJ0NrNBwZ750OzfVbl9o81M2zl/gZx+Dyc3msLm+GN33L3cKgLGLMeIUz3i
T1CizMsIBBZT2t5tbnuDn7peIa7HECxnWBJm/EPCPG0EE3D5H0kAbOvSoUOH+H+X
LPoC2joElEFQje+DGNaDvXqd6DkO2rf2tmh+qYzN5+Q7Gz4X1CWqDuIYKq/d0DKx
mHWv9rFPAay76Jq/eOc8hSopiOeUwh77nlULNwNQ8hrDo4E9IvI1Mg3KJN5TQ+QU
kUOuayC9m2ZEeaVvKs7ZPCnStMklo/y0HbwtaiT4EwuMwDmWxL4/M7ckDr9M2O3k
wlFI6gobxBDxAEK8hktWdu+mQCH6bKwmt9yyvUz0+7zIT8mrXchzBHYqBqPJU9wW
jec45QQROxgtLmyXUJ6llMFvLSsDg27x737vcneJGb+gX5fNU/Zb1gokZwC8jxVS
lDe+Csjw0XrZKgrtRbNTpEZptUGg2hv47KX9vefKbbKNePpMg5StmgF+3Mges8TJ
cmaXLKHYIBzT9NSldHO4NOA53BApm6iZLJ1ArqqOdUcdWmpYalT7vWYoTXgR/6N3
iYe+6ga7bwp3DXhGdiVeMFTmlG9LIEtf7Y2X1WsKf7jaRI586es0CapeV+y3Gght
qLXuxLQ9SSpTpoBQ6HS+QHtWPeK5nbPe5A6sjDyW1eup+PJsHHcnJOd3MpCjn/Kf
Dr6r/fxfThZASBdmtwKEjU2lwQsyDKLKZJvPV49k56AofWNeu3JFu6CokYZmsZ2k
W5maW1j6C0RgM/NlD/17k/icG6WZ/0tKmySpv+GE338vt2GlyzimIgJzLZZQi6JI
Jn0R/picA55JWVd4+0VNnrkkglS2CO0VkRp5ddYVbFz4e7E/1cH29KRnU6Kh2I3R
8EUg3GR+9KawhvXDHKukDqspURnSiG0o8RCNx7AUD23BbWRodn4EUBY5SUOGYVsw
HlGkBE4PT7/kfWI7GjLCVlmV1wRTfX2p2iBLxkP7GDknQ1RqnfXu/VfiB8NMOu2S
ZIVLud5WFs5ohJpLRNpSvbdAuy5Ig69Qw5DUFX/cNFDJ/+6/ZfY65fJAo5oXdRSF
iEu30EKSEtQ+3PclWOlNwrUw3glJ3yungbowt39wNzcdHPFcaJRu0LjFkRMGEAY8
csZ+148COWiq37FqiTbQ1scALUN45eecFFTntxNyvUcC1Op+dPlrBnCX310Jg3Ot
2NHLBSpyUZaP8hSWjo9wf0eGZUU9QdBKAf1Z69J1f7aBBsYQ0Xl6AA8UcQjqScSu
aiL+ufxoA23m3afpUYMzn81JYu9f8S+LxlzDvt7T2eAnuU0eqhnXjSScm3mk3P7H
L6XvmrwYVcAvj7Tc2uLKOMvzH1278lDk8S7EtthXMR0Ls/rjjTp/sXA6ThM2ksZH
ULXxvTkRS6MuTCW9FDY5Je4K7hcHpwmVPhuak16mZQKHPkSgL+57nczb1z78qkmI
kPIvHycI4N3ajQBHjrIHf5zOBiivjTLAgJWCCGp0OHb2E3ztqjQtVdBZj6vq6J5k
WjkbIw12AIdu79MCecnytS9qnJ9Rpz2ZT5BNos1W1qEQQ1CcOoUcV+PekOe+baTb
8t1lwpF5iy6jWOV76SWVkBo8Ko601Fp1LSn783X626+1nnPFCKs2gheRb3i9Fb+/
qIEJ0/2DlMFKAO6v76Z6zWtvLAHaWLm2Nb7j9l3f2/ogM1f0YgIFVuAZ3RhOmFC1
DHzqwQlhOOr97mrEDoBHkABXkQd53TzgDHQ8n1aWDS3TGmSizm0LuYtxVq7vzE1Q
P6MD8NcNi8EXBAQOffmK/gD/0Z9uF72JFRP5zV3tf6GKw5sjvCjLw6LrYmzv+ZYz
KOof6BgVASeaUEoDFEGQq+qfIlJcoAaLOnvcvkaGCYZ8dEUeO4tfL6wMmuk8lLEY
zrRZci+JZ4o9Y3QBnBNfkRJnsAujMdgzAN3gDX6tqfiKfpPezoKijM0Ra8W+RArH
NrSOa5tGh4k3efsHI1zJ00n6ydYO81c7K9i262oSHdqfPreuaLgTX95cR3dmSqVd
J5Z/yPJ3XqSdaC3rVwTPNZtY5NHZ9JDXMyfu1/0esEIlX9bYhd4y2IKbE9DDJ7LI
Nw6mkjsj127bZq3Z7leWXuGqG+ND6SGnH95jPcaXiFDWZjrqEShmONKHdlMq7Zj+
NOrKL5N8reA+pqULp1PGPJ0LAB4IDgUgBPpm1DHBYkpssrMOwMN/Z5BsZRiHvG6a
2wPLLDnIZWaZ1OwyRdP99a2oekoR/b1pWubqAJfdABjO928GvszeEBZDiIjnXdDe
OYjaFmSxyfcgXelA/xhKmij0zy2QHTDabF27avu9gRmCTt+kt/rhEdFxh4lB6kVB
AXfk+56C5n8MWXvzAFdaLRhq8tGgJJxSwVhnRrEcvOQYUlvQf6oUvVy/UNi/yyqo
HZ6GmWhGUiFeznNHBsbefszQ0LyzkrvzvgF99H4ElR3d19MGGOHQfOghDhr3bXlc
RJii25VNft7Xn7mLra89RD+/UkbrgrxlH09q//8hS3TBlPL13VVr78h7aIaKlTVV
YxrZeRKudjdxkAOQ7xWS3APxxU3g35NqGMd4YRI2v2oNaROy4IfpED5210acGihF
5cx+sLIVaBYcof1i4f6aimn2f3yw3VdKX1K16Qr1W40sFabcIoCQ9m1x0v28ELGV
sFfYiW/TOvG5FLPXmdD9hApS9dkUkprj6cbpm6rGcUQP7P0031QfTOdwgX0GoC3W
As+ViBgmnjM1U+VA5qJxW/DpAbXiNcI8AIqzJA1925qdJtDGwILGb0CgRl+DM0sm
K9JcJ7Q+KthF0AhUdR5anAZmw4xkyt6PQgYfLu/qdBuowdWm7cM/sLY+AIq8fr+Q
fNKBX5syZQawRq9ovyAYWw8X8Mc/3i4+NcTbkoaBWymctMicDCeO7EcGsoVn4tw5
ehDv6re8Uuk7KHc6bGOYub6DjREV9dR2VRBhVGvl+c5yyDl0AQkr7ajcaDnDJtfO
DfiTTt1/tYrR9sxB40muxu282eM2IP0Jf3EnrZpeW9Jf1jtda1T6cKx3uIifyywf
rPqoYApqVRGBDXKEiWBZq6aooeHQS6X19wDQMRdvh+8GE4yFm4Bdc4bdi+meo2Ve
uoaQbwT43h7WT1hhxnI9mbDg8fz8wr5a8eiXU3NRXQR7oNJvXUg8gwaO36o3dqcn
42Au7Ds+HvYE89sJ6Gvab8ramc2QxovsvHg6cm07BG5SM1kW6xz6oXIus5wpvptY
OOiz4ebHqDRy/Dy4ab5MtkyuhX/8USR2xeB9K6H4BOppd7jPpfjZawj/nccJeGas
y76clrTbk89y3us333dAlVnnxnKgtLKE7t8kMK01LtddetTZ59rOoPWLbUhO0TA5
1gFOWSAw6pCF/Yka9CpNyjSKIJI0PA8dDNGTyPp2/I+KsvoTScz8F0U8ReWDsm3N
5icpt0BUAyCalp2D6onyAjLY31k8HTDBt/Lb2l+yXIP5+qQJtJRqzEf4JEUFqI8J
H0CxbJ9evV1b3YLpUNL+Vepw+Xe54S4aEDTL6anxFpx76qx/9+0cr+8QzC2bfO+Z
znqYykWct+uvG4d/a6aet0CVfODvp/nXkrsEYG9qAhdMLpk313M2Cqs0bK4KsYlJ
jrryBu34ADEP0s9sqqJKUUX4J80hqkWDrsTVNZOkRghjRIr90LCXfrBSFvL+A8QR
GWcp8NWc2RQmMnwn+ClfboDL98WIknph8hN/GG4MJLG2W5yIp0Gr/p2mP8jhwN/B
VTi4grztVJSGSsIXhkK4zMWAncnyJwJQlDLmLX+MhPaETcLdhmx1eZ1SEWMl6rwo
SBkHD6U8zKI5GioiXLUQ/13++Fai+3KPfGhWEmlqv41EEFdz9CgMQgvQ2X8G87s/
PUVji/EIqCV3LvfCcapRfc+P/UjXtBuHROCzRpYW/5qiffrzLJMnUMzQDQ+0rDX5
Q9lrPCJOPZ3bUMbkr2LgQlor971TS6wc6pKRPNUYZypRQAvI1BKnktk0eCCb6I4e
e8xESnm6fHZII1PRV6z9+hRpvvdRLECnwM042yPAAL8U+FpHh3+HQZu6b/+E4HmF
9xYD+sILz37rH/tKUqcsn7lGvdX8eKy8ZE+yW5uhBriT7RbNm5AQJM7mW/dLmaWF
YAT8piNZlMbaMsRAeHul5DezxGi1N6sZX9dRVN5cjG+2X8lzXTPkW7xV+IpM4D75
XmPFNHYdXZ7Z5np6OJrCvmrKK9Y5Y2iSViNPKydOx8lH8jTebfi+Z0YTVspS4IF+
OKykSTTv1YTTW33wLJRP4qaJAe9BC2QRzW48cgNKzEA01ENQ1PMOQHD22M2sJkxO
iUuFSIUxUzX26fwutFmdyBBDZ8v3qtFNRmk4rtB0pWc9Vc5g8o4CX1wyYnTMECLu
QTOaDyaifwg3NNXnswt6LopvlU4ue3EJ+/B6RKhGMGfhQoIHf82OfUxRYKOSAomZ
GuBE75lrCGdFdfcqOBjTd0y3FQMrNANbcfaAq/sbNhJ7dSQb5RT2dbMVw4BlqyWC
VL6lEr2VQxiWQkdANiFNwb1Hi1LJDCgWnmf3l+0HE3oWax4s/ixkBVmL9LfYaRQH
0Ed5rfNnCj3cJ+V/p3Q5Se5/Y2EUC1d6tpjYtkC+qWUL5Mh2DoLjYhHgRB0D+1/f
znLRAqe7+zIDZnKcIxzyun08jsXcjBFarYVLL3hGsm+8DKS1rVFGx0QRPi9YZzy2
djD5LF2MdOJbF27aU8jjk9BR/77t+TW2mPcoUnBGAHM3qDWMyzMxtP/4m/ejbtLM
bWQC10gfh1t5NoWDSutplMUv4Jh9wntPfNR82NyWjIM7FGD875ywvn93AzT81YN6
T+qlx7WLrIBYfbXFMCYf5sqvKnyuPHDMXDg9AKHyTZXTIpyzTZgHrfy69DCqFLMS
/ks/XyNOviMHEXCj6N5KaDgVVzr8LcmUGJ6BGzzzN6ntshwGRE1BwUnH+SabIxU5
6R3D2U7KSlnlnsm09YMKC6NCueTp6SSH/Ro3FZC2iw06Z5LVeZ2e6Z6Z9T/ymz32
COk5pshoGVPAl68Il4nNpZ6duYVVRCt4XXPZVX/6Yx0=
`protect END_PROTECTED