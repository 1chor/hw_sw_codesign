-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Tl6xBR+CTPyGO/1cOAD0JcHyKoorq+b0VNDu3ocktK3yU1/UjZY9ZjNxFde0zJlb
l4ZiqKGKkz+7dJEF+fzbFIwcJEKRDc+NgQWoC836gtrUnK0gB0h7FZYQDNx54gnq
aRi5K17UYoFSBhvosYgdY6qf/cEl8rSACn0t0FwRXns=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 79872)
`protect data_block
3uJfB5ie6me29l7tl/G1VHk7hSBYSvKqFOdeXO5GG6d27YJmeL1iO/8FzQGZbLNs
+4W6XHBiQtDkq0m3HemVlQEcVsjNHCZUWjjPL98eEsS8BKmdN6EKRKA/50AuISCG
L7lcYT5OmGi8PsVmPYfSGILEO1uNgf0U4Xf+lEnTTvD/sfvelwOrdKs/GSuPWIQT
b+vHCcuLWtNy8tNjbrdgl2orTezTAgrH3kVo5XyUhv5QD/NTrj4AIYZaUKnczr64
CPPdBTV88bBuNTJcANlP/Sc99BXkPRdFFe5LJpUNJpCQioIS+AboyUht+MvgobgQ
PrAHz7TzjBLHffscE9SC/O/NZXYPMUwghxDTiyUTYeKh2hgjpQd4qhzfL/SOrX6i
PmDqdT2SQB4I3zT8kUkvZAfaonRsFuH+9WGkSRv/7zVPelendYlRxEtTcB3yuPYP
H9mzRrNWKpqw/XjMGBG/wSjnSwHfkICShFM4dt0S68LreZy9PhVF1C3eSwZgtSO7
eI5pERRhT9lK7DM77qreiBX1tMzw4DplrpmGFftxcq8c8kA6RcMLRD9XLNC0wJmk
kfYiqW5oaTwvZYhbyAML3pbotWm1c5SjI+HzNgTDlC054ewdYuDmF1fmSFaMeES/
1c/NB9CnYtkNEw1KfobxgsPmHWx9EXvMO20oR29ghIsfAKwBXeMluI1eGDUx9Sgy
Zv4OP0fZSX6izMWZTsOzVX4IXr8sDj0Z7zzJtw5b/Tt2r21LbdECHFD0FcX+sOM7
JqMenfrv21Z+XeGJ+7zpKgA0hbl1TaI+TKKjz11ezg3nCaLisefx5dyJ5YQV9hha
cqZqQrHgkyGk44t9u4kS8BYybY/PeMXrOJWfggI8zhxa5/63Q30w8pOpDrETr5/O
CkEoAeGzXyikZEFIAmiViyD0HpU3dPnY96apTEQp4H0dFLIl4BcQC2kXwlkE3T23
FIBcwLsiuGvYEj0hth1aB3VlepVaGjv5SrSBkSDpwB6oPvzDJ8qE0X3mfa4fRqp4
hjRvzY1yl+paDPkLAjkGRxptH90ELwvX6PR5F19w5P9TH9coo1G+egNxdOVTTU1E
9/goARQLIXhhc9bNiYKIgRMyNtFTFJUvN5JBm8oUrZxhRyPFGtBiwP4Bi5whNQAh
DzEKhpKvjpMbjjzY/tPZZyrm8XbMOM0swPnFH2+YUo1SEV0EL8qw3Eequw8h42Qp
iZCGBZ6UrVOl+w+YpQMXKk4/kKriBeqciVlAtR+VXeb4XORPloCqAOXVtGh2+Xd2
0zhT4d3pxINLdMXjY8wZYoIYovTqvWuMuYTs3Nn2oIB+z+HSlLGz1ia0caiJRyCA
QjClsbzWmB13w/McQhnGNvHUfuGTJ+4J73xDToMgAhXgKcv/v+6hZ/s/nnZxGiLD
MpONstrWTfgEqSgsy+DHMRb4r0+KaoTsyqAmGJjfx6WZIOQzD8aO0t3lliCRUZzC
T/qjPAIjehbmngSfRSfinPdUQbfA25Zcm/40OCbl/aghlX6Q5MhzQNVtSk/EVXSC
LSC/+NF0G0LFfPijJ3T5tZhj8uww0gFwXJ3guuoDHXOHEO5HUEildliGKy6u8yi9
Orwo1A8KWPrd3DRg6Mz/N7YjZsrQMjcclPxnputrmST6J+JZ1EkNLPoceSbMcFlj
2h7B1KcGoooLH6DpdeTyV1KtlGVANWDiwdcYWjgN9tNGSZ78LW8dBtiL+QW73kx1
O3SSrMZmh9pNVTAays+LKsyhzPGbKVeI6ODKvkVdtiVWIPLZO663v8dsHdDrTdss
sGqxOHOTaiPOF6jshwYEyds2/tkeuUNPT+lM/2LErSQejgWi2nzszwSOaCQ9YWQu
zZqwYIHHGv2y8EbWIwy5xYZKa79vbv4V9C2x3ChPq6zbfb0esnrjiTAtNlc+8rWJ
3XHG+eFWGO/Qe+sQGih8SkPXrhwrau010m7Pp30CI1vOw99Sk9yENVKeFQ/JSgrO
QYYiqya+f4ybAatDWUd6Wt4eQMKEldPQ80ZoQHNjdAupLUqw2Zx4Iqw0U3oXaxCG
vlUbr49PL/YYokOk/2HC7y8jXlEjh/hJohYUN2VllGSd6qt7H21SRXDzHbwlsfHq
7sbNJKSFRu4HQ/BR/tr9D+1Um5eZbNhE+T5V+zj4wbB2OMX0wuGM+A+zNU+1Q150
GRXjg3HUc4PdtzaNuIecwGhT8OFf1vozW21Y2GZAIEip2MPjr5R44EEeWcH4yODQ
DWYgufuQ1MqKzmFybk7zIbnexvI5hhiN3GewqJBCpKp61wFIdu2zRSzSRPl6Sr9/
8gFYHanFb0T/jgwGImVQelmNq+5Q57Ttefbv7goQK1J+221r67JcrjZ9P+vc7AmS
yk1SQAh6Cn+1+APNKvWk4gtIMnt+QRZXgJKlpFMOQAU2xXJsZANPkkwpz8YjjK8P
LCNG1SQOZ//sl2yEPtJ/Qnwvdljs0BQbdJK9OApG3MDm51nyqhk3efg6jfiRACOJ
ZDs5XWLFgBUcwVKz0/O/9nl5yqjHyu5xnYm+uuF/YbapM6OEJzbosGXs/GaKAyUw
DrP5F2L8VhzLaNAQk2oNeuGswif+MQLFF2/NlmyYPJpMh5c9OzLzDxBOXINWehNp
TYGfr+5p7NZ+wyl5qhXd+c1ZM51+pr4UHycivq1g+VLsU6LQ1FADRGGePG+hj/0V
M7mX4ebxa6NfDcZzC8Q7YpKIfwkk17xfb7cEG2zjCasHeUna7MlV65wXfiVymVM3
zzoEP+bQcsGnYeqJH6KXncMy+xIR7fX4irtzL0U2k2Mkrh3B/OKifKgthhD7V9OX
2sUNTg4i4Pf7nSmWW7q7MPFCiYE7U7cImGpITsGwWXQHMEaYN1Am7uUHJH/ZKt1P
kV6nm7dRy6EUaItuseZHxErwMKgYHRwgrKgasSaIHQrUDzR0JQagTciB079JDrb0
B6eBAV7VRKLmsviT3Y8pEjjTjnSnJuicqoBS04csmaA6JXx8o78PHWVIroqMVa3R
15nQaOGuAO4K+bZr6gc4aGQLqLGpIhWaXpxLVT9sGmmnqH5f/m0HgBDEgqGRLbyp
GeMWNM4jrJTRpRDNHi22hRhwgH2qLY3Wnca2tkIcfl/CZcovl8W4BGT5LGAe8ezq
GHQ3MB7DETfL6x9MY+b7XGOVscFBH9qHceWeg51Jb/pn4mj3VF1djbgY6R/uIUcB
1MH6Uek0TmMSXegmUeKdFtQj5Nh+8+7XbJU18HWwaQkmGch+dHXPwvmEyFbqrPF4
NoL0LUEaLIpmq8GKI7Um50hTVvBCWWyXRefNLqPI//DhgNLQt5MwqYmPh0AwdsA0
9zcVy+8ZxT7UKLYwzxe15kfZjx7c8jepCx7MVqaorfQfAW1IVaSdF8MIWqlEaUZU
xrymJ4DPAsNKSiPb8HBae4WyHCvkRfcuIGiE/coZIxXYg8+QymSqHE/dUXPxRlmG
9wXIMAtC9iGxU6OXpPg6BFWRgQ/YPuy8M8TONVuoYqgRc/U0qgbT48SjD4BwMNuI
8PuXuIiAmdDbtDy0mt3hC6GZtdAKr9hjUYDWGnZAxKTNpUhtIZo0jNUY5dTiAT/X
jD0FL6w9ofCd2CQ0WfRVrXupWGT94G/cQdQlymPl6OZ4NTsafLBYm9K5lS5UgdQa
+Yz4TMhOYF/iJ5bxuG6I8voatB0OHz4NijvVaTsyMszhqUpMlm6N5yYSQwJqbk/6
SMkxtDTk7WhhuQ+YhwGRlNbxT0eDYT//3m0+LMkxFmnEXeI0bjqjSL9llCJktUGo
H9wroBWfz20LrK0NsxL4FzI5G5fMkO5C3w/1pmSgX/fujGUON+DQVvnUsNOAqzuZ
4Bozgc2vuUwDE7+N9Iw61c5BpKy4LUIkfEuRXWq7QXc/22riy2bRU2k6H18BI13c
cFQxNQ3mK0k3hIR5spZuntCsHF6UirB8Zt5MjUxWQUbUiKX8QuWmNDSsJHsdWw0C
DnYQJacrB8d5xVMwrhUjoeb1BpdgRLVXHy0Ock2axYQGhClMvFK9f2DqFN3MyOeV
buNkGqlkjLDKHIleXIbZfVgE1FyyK1tnEornqtVOeRNHmzuhxVbBYO+C9wXJjWeZ
m4dz/YLiO6Rn5Fxw8q5MJU6usadKgRRmKMw9VRPxdfa9NR9dhZ5Lt+IxKT12oUmn
QSyLMT8GjPmuxO7KqCusMfYRbcYC0RLXLHVZgfKim79hLC6qh0Dw9p6nE5+8jrzn
y8qXT4SqzezsKseZAoVjZStC+Gdsa2adlQkJjAd45H9C70kX5dvgsfoWd/3gHG80
3R8DALWQttc9vvIqAYAjyAkY7I7DSP9ZPu2fatf+PFm4YKwWMSg/CWw1qDR6GYFe
gjmup32tlNkwBSxeaKwOHQEWxYWKTO2Yp7iSHfbNy+9oPq7NNj4VJsYpC2gf0a6m
OuNeR7GWLRYpvfaLL12v1j58/1XqlcN6aKq6OoCbndbgZAB8nD+gyfijrEMDNK/k
1ZBYjlrQvycn+0e+PTTN2yz/k43ClD+HQ6VtHiPBgr73S9su/k2rSMYiW4bilAof
AdQzHekdUiSKOySsy4dBvNCAO4Ih/UWc2iSKAczGxgVk/DQSH89Xf+ZURzwqVjEq
Ita0/TGrMiYe5XWkFW5oqs+GWCDsMqahCkppvPfNFXOB94Qvjz7nncEltl0QgT11
O4TjFeVEuHH94R335QrK0uxlQOe1W1FlKCAdenMw6lNTSaTQkRXPk07ujZjbqRH8
+fgaff3ZxTYnfAAhWw4ZNZf9dG1GxefFoURD/s0G7mwCL8Lxgn5OpGpB8RgQww3Z
7NH44wRk3+gdDohsiIfbhq1SfKLPdWYofuZzv3kH6AI+362Y6VPD5GYhI13lchUS
KGP+zdw3y8yGw3LpYC3GDaiy6IPc+JeKHdtX795T2qoR5I0YBH/Ed8JroC+PtxzJ
WqjAGZQST1kSJG1gUa6+B7H+5vAB4RFEgZ9zpRxmQGZy8g9rcaUxm3JV/LNCrgXD
NmlzlVsdjmCthLOWtlwDbws1uJTlbUlAV/994Y1WtvoV2UKkXG1L/ASjQe8vzMld
c8Hbsm5XC/rtF/8AW1qXHHog0sxNletblhyXi1Ic1MxbflwmAhMvExQdUm3I70YG
dM01kwvommWaZN7XTWj//2uVT2wEYF+zeBNuAT3gtp77zbXHFPvWcdLcL2m3BTK3
9dqbIr4Ehlmq2IHC+F8L6zdWnw5TfdfrnAnjHcgpKYxkxU0f8j7AtDv0MBaATKMs
7w+0qKuScOk8ygBV1TA4CVBpHrzWBEO41pswcAFfrHgoGTYwlcXC4tPQ6gtYis3r
cgQKv9zvtj4uVyGq4ri+CAI1AFrWas8UnP7rxTGCp+qMNcduAEumhJgQVUngqpIl
c51tndNMz8HG53bn3sGvMLx6VhIE53/SXxM9u03/WkjXuj1X6cMBfLgu3F7WcM5P
IeS4EdhWhQITM5dUAP2wecAYUUCfKGx/08lHy1DLRkRqEQz4ljoSHRvK2t0JuEwb
lTxrN/7ddHVxjX3Xwwwgm8IWAGmnlktOwL4tFRFE8kiZIiXUjDyRYXP7qwubp8EV
9Fla3h0cGG0BeR000rkcYa8XfkSjt8sc4fFLNi1W5IRndFsG61qncVd1DHFPQpSa
2YFISj1XVAGfDA1PEyu+ekM8J5MvleLV2wn2wm1AzMcTPpsKcUqBRTzMVOXd3SQJ
S9S0IJp5EKgQrheJZRtEUCvXu8k7rkJWWW1bV/vZclGbrMnlv0B751xnHy78Lys7
96as16yX9uPG4EpD9RVSRn2nqqPMtkN6UySlxXLY3Z66YoivO3olMYJcCvT72fu3
9kFSaUT6tggkK+789CZwipZrvmJCSM/kaDK9AEbq2BOtOQ7OavkVwYA4w6L0cr5T
IJBeoY6ho9z+pP0/8NcP4p+kCQ0uCAY8duOkqV7PjER0war1uhWbe2I1O+qZmlJ+
EVkvAWx9tGkuixsgqaUXXOfcm5gD8YijpYJJluBw5s/Zcbrhcq26XfZl12B1VujY
iYjji8IZvwWUDsuI3+95EJauoEwPojYYcMX/GKMijyLHg58pVjktwrZJ+FAGSHpn
83MryFlcoIOhar/3qyaWb7tr6Ml8WwdmuhX6H91d0FlMn4zo9DWDaZJmPzVzhnTt
jbLAhbfLbXmUFBqPFZ/ATa0GgsIXHWnvDULvjIdl66rCviTHT4jdeK6Bir2S2kxO
BUYpdoLcF8Ixt1o5EyTyz1ZJLgACXqym/bWPEKtMnjd82H0GbvZRoMqSSVEN5YZQ
D9xCm3TKQJ8aA+1xaZLOytIXEOX+7ZytNkhRLyP4eVjaZUpTew2PboZV8g+GxWri
Afc5jLGkYME48boTvP5ntr2/A14/1aQOo9lK0G5tMpzeJmf6VgPpFz9fmx7o1q40
CXTdZj/d3eDmOOHx29s8a3+LXWmd9arff3oOCsz4XguBRJi8ItnqF3UxpJVqAeH1
PAWCEnN63hrT6NGRvXGCEYsEdTvKEejGv6u8BeEplu5eFZmDr22njB9VPNpAWweQ
kiYoi6vlfEPF8YJqLa04fv9d79khqDn1sK+GRRscj5smnFmTvqbG3aq11hHXv0le
F3cG62/vYUoiIy1goSs6CI8e0jOK2xIuoH0631ozlZr1HErTSpE5c/1WdYOJjW/1
Q+NXbxVGNBUuC9Spx/E9vZy0onyjQGSKZw8+GajYY/b1fKPBM6Y/8O3CP4rMFtyj
yibvdoXt/lLH2k+PU3S576XMp0nDLXvLhicKUtW0FoW2G/nA5i19tDrTQ8/vKBvS
brHlPqrzUwgpmN6QgBBKhSaJjoPDAvecB6xIfyc9Y5ukC5YwLJTox9b4g5mrgwRh
OFGlo9uaM0xTfaTkRoj3NVGpKkFj/1jDKkDuFnJiNxxV0LPa1aoBSFWtgXJBdg4B
8RIy+4Kaqw4tRHoF5DuCtch2j0ljpTTSx63Z96148bILmI7fJPbLbw5EgzIzB7zq
lyhTuQ0imEl9vEhXauxHyp3T8aWZC335OzifDsFB3EDhsEs/NFAdwPdXImhThGvI
s7OccWPgMvupevLiE8yh0DIuPPZGPn8wBdCNVuGOu00dhgyqLWvV4Im8r9bF1sTd
ARK7uTR8EOyY1fl+g4w37Z032EhcCpbKdQm2L4LA+eE5JjmOoYWOImj3JJycB+qv
i+jA3RNiYnXvwCXBvDsUvP7I8bXtLwLOjYzyE+awRjvDgOrPqNIkPEp4whxxGfje
JQYn+IgDXsXwp9oRCLzZuvT7/fqRwXjL4KY2essqFw9aVT5R5PslQvuPhTImV8DW
6c2CD0S8xoI5s+XTzwib/+HtRGxicmvnHZeBINmb2mSb30lyrZkFYC/AJLK++fdT
IoENY+pGulwWjod5lPfKtrc4EBD3HdJOuNkn+jRNQx+sjWyA8zqVxd3pHKV5Yq+t
HsX7TLoPVuWJySuGDdAw1EDtEOslrRGvDtm6AuZVdMEaFKdRvIiuSuxluqgrsqWe
CHMg2UWxHgGWceg/k2YVtcjF8C0Y9FH8qZrz9GT/PLGXF4FkuEcfKQnqWIDtpOXx
yBuzmj09LvgPNdrEb+yX0gdLC1V1dWfV6w32ycwwjsrR1l08AWbbQAO5m2ZUG+pt
FU2bIXY4pBetCiRWQH0IEs+KRCZLIlbohikbVR1s5V9Yf6NozTPknSapHhQ5t8e5
Ig+8v6rVQTe9WiRJZSXxbNZWzFuVnGN82qjtKZUyhzqSI0iGWsUXU8J1ahifTJTz
G8Tx91Cp9T7PyP9scHnG9gL4mTE3EISbOy6yo8aeT+pi/kbcZjXH4OscLLYBfu9U
F9zw/mSmGyFOeLfnwE0yFm4lswpSW6gZ0XVD0IC1dVL4d5Y8Y+vlSPASGwvFmkYG
ncg9OdFfUhUQZHuqfh15u6P3mDB3etoqqIeKUk1V5c0z9e8bDm3tOeO5EY1wbWbT
9ACFk52Ggjfvvo9cR4R/1pHD20tRJ68bjFXoZ82l3HCwexVa1YI7Dc2u9gVEJ304
ADVwNugWDVRiQrHKjDg56fA/CH2FeKCMYv8LE9Rln52z/4uYaMuUZ6PGQBY0F+A7
mQfaI/whRQE2MbmrbY+w6dAtF/DGI1Y2H8TBcrqgM8e067Gg17CHCW3CAoi8HZA6
5JCHPkVgqCQX5aZZ01hXr3Jx9cOhI+mpfQZyj/jAiCBSdKga66A+N5KMUS/9jbqt
yptPJZooy3fifbjM0RZMOo/75u9kcSf7aR7UdLSGTOEX5gSwtClBSER9W53ohR9y
i+7+Vkjtdgt+qfvLGVzzO0sNnbIVbSdkWEAmgeHeCh3oy5rSEI57KU9NYjyljs2l
ejZAvaq/P3+d/iFl4J4MGC+192YxHeP2gSGjTinc18m4y++5RRmRLIUbh+vCe3My
yzdzhU3roHWpvMmjHJBbEbFBwIYvYM/s8mjsi16uUAqw2N3h3qqBp5mPAXE0B81S
b1bxsdJGI5xCRXxctCB6/4j7k2ISu/eij7eHfDqhDrqhwt3PIoueyKjrd/pjvL/H
ki6oDLGVKI0YJ6HK4Yw3BkE1Tm1n7rnki5htd9d6P8oyOW0usrlD1ZStsGjrFqUz
2K3Mo3c7BUYj+5hdxFDuBEjcT95qmokC4NQL8J27HV5pTm/Dx4GLPuohRx7SE/RN
UOpltOFg0kqpqeAMxgeZgKKNzK3TuWsrF86mGpXPmLNpwtG9gTmqindHb5qZo0Qq
xFCS3k7P51glPrIGmjUc1xL1xHLEQRBj0bJG3JDLjeFPwPWWBenkzk3W++wwGKM9
9Mt0xwJ4mWbxxbYzYKZwFfUHuHAHLaVPetxO8jkxpwhIbv882czI8qoTBML3qis3
6j0wgkFjJIrvT8+A+2dH6727eIsef0bBAcRvZ9tv4ppA+b2cRVBnpQgMRXzUiTj4
UzErV8x7lFoJQxvSnCU7coNe/APRBf7ATAUGCIV17HDaoX6tcWofq7RlsZV8g31w
8y29FkuQs8G+r5+XtdLstUhk0lzNDzd00T2MhdL2YEU6nvFYuRKFrbHIbLIaslxP
Omy+5t7Y0Uq50ZTtS5JWGabUlJfkG5LndtiEXYgGHbhm3cAAcEyvOKfaoXPT0oSK
EuOLeQ5o/cO8a3Fjyb/kKqVTbmbPD9q+o9UeMAiKTOvtzdBhhhdoiBXIuNr/351Z
T8b8urTGzsoBbWXT3kX9G53D+V30zkA0U7NzWMGmpE5Xg+qNkVfAOGOs0Kktj7eG
A3dDvMXbC7E7BAdeX85boZZjYsj/pub/IlHVIR3BcN2TZwDrBsgbFHmcdzyfcuHi
kb6yqe/X6sSLOf7hLv13CxL70wUcK6e0yyy5bFmA6RGq0cDzrz9aHflswf9bCsGt
9DJID8Ldvcg/Kwmxb/g8qyb1c0MQrb2IEfDrZ6RyNDeF8u5NQoGSPDu/+dG2g2Mh
Y8FuJD3eN9EHUYUJWRuHcmDHz0OL6So+Ng7Vx5rSHyAjQa1UEvfTor5qGFPMgX6P
K8w7iY6eRtW5LkYO2TnSO+eI028iwv8gT9johbc4M+BCbQb/OM2iArDP+4uXpdN/
9cMiq3UzgpJWJNaAylBAoWVLF6TpNRXaoQfmyvjwvI2hyJqdOApQabll8GhrGViU
gjNAsB3C7rFUOIzkqqHCzp1f1YU5q7sgwdkNBOdAJWlGqmvVx1GKQG9nGNLMBedo
lZ+rUJUoJGyS89V4g90XJjAc2myA/a4e7P3sbQvAVEupjK+wFtY6+JVRyaIr/7t8
IyEYYw+ZRqswGtYn3mvJkSR6RWB6b5x/C6PuK3MB5VrcWNNyc0hzOn4UX9oM+cIn
i/0fRr5cBKNhhIWzdYErOEUQuoWINHbjpPJx8j4GUew55/eFdr9bw7fs8sbF3A7y
bAa2HsqSSb9qiGIYgXVJamz4gMyvmQgYKtbfm40QqLsT760xV8sp3y01R3VGoz60
25+p6u0bVyHVN92OgOJhDXaNtXXpOn3cnp2aEwstdBkgPcUG9/8d/QJ2JtDJV/u8
q5rnswNux9BKzIHmH8u0FB6jesW6uYPrmhZPYAV4khm58D02xJeh55Kxyb6zjzJw
c3MIwlfk+tsw8g40Pzg3vMIIRnDltI1bD4DO6NLMcYvftRIKcD/Z/26hVxVeglhV
AQraNW9LpbMoxpRxvM46ge6m3fgDKt9Y/LL9LKEWUAHkVF3Pae9dECaDZo7A2Uvw
0DfJ2WblfdV1YW0mrb66JaGLlGm97SzEG0biL2DoAE5Zq0Z2spEQrFpD71xpyMzd
Og2ut+vqV8lOWnxNxEIDEERKRGMfXB96qp5skJblVs7ppD4mKLGUc1BwSHqAyST8
6RyIv4htjFYyRKoIAjt+cykxOuYf7EXeABlSNQ2rzjcJcdxrah93PLp5yFvtY8jw
zdkMbOASE+1wIhgSuGJCKtALVTM5W6Urce9OUQ3hEWgQ6copL1skOwBGa5yz+mnI
To2aMD6BMX+6z/dhrnzlmWgJYqvUZvgk89wOvQciapWnsVpypADc6gnMw5JEZHpO
uGKOHbl5hnHed4869ER8PzXoREzxwInx/6/DhA40At4FuzJDWv2UgemxS0ZnzX9q
PdaH28u0T2PuI3cReMRYDtLWj0QYsbpDrQl6A9d8Ynhd4QEJKXf6PdYqXhwokPtR
VK98JkaTfzUJqk228q6mrdwgLkri8OopIsWX+QAu5gTmEvqs9fl2Q42AoAYHOEaB
lTijOWBxIVtOSQkN+sRP6+KZAhVriJgCeC60Rrx4aiMoRM62Ht0IRdGmtu1PIjY3
HlTk5o6qx94fQs8+6W4gJY9K56EnwNAiAy3iXe8VU4LKkqS1eeLWSiyip9alDauL
CuZuOOnBGEwooP7SP9QviW05+gPBOlAlnnI7XiaxlxGNDikz7IjxAYvaS2A8QKAm
DBQmtjEl3my85w8ZfVs/cP2nxlADUz2R/NucoRPuiCgsH3T8X5CTPzlypQl5ThrU
8wsTZO7ykJfVXLSgn+CCKeWvMLOQLclceRP3ANOr3+IsqAZwqx4/HJriJ1I+SgOw
/lOZhHnxju36SNQAMgw6Asq5lcEpvWvBW3a9nxzOKxy4s4ATda5fRKR5iqNMKLi6
G1NCfedF74tMS+2x+x3sUFoND130tGuJAiYFQRN7B1n+pnlyWS+tYUmpcnRWL3tE
NWwLLTTreDhgyQimlz1Go8uSpSpXRGuRlzXMkLuVUnblXzZt8ewAw0I6ioYk975a
fa6YxI+bm3t4eLdLG28TV/55cNXnauEjdqvITh5GXgs+NhSm0vUrq0yKAPJgGXeD
hrDwCwFUJrSzTBq72h3t7JecIYjy0YMr+Rfdg11ZXB3jErbo/7ExU5PWE9gCqWxc
BHy1e4NBgqlD7eVkTNP6Mky2qx4MIWpOoTDxrp8Fy8cpBAwxHsvkHLGp1p+RQsQH
EdNy5gYqyZlyeNPD3ULyGbwRUCVO2rm6TTYHWQkL6kN8A7PoaOd1EViGFyuDJMDg
bv7TDi8/E+JJccrq4VLYZDFglUKRUjINTXbGugMfUM5hDyuEE70G29ruX2gFZKZm
MW2FJZQbwvQSNc5ykbrI2fAjDwQGjlXluSoKKiYsL20yUpbTxrGwKcfLSPAIVaiD
Da2emTDF+ylm9eeazdR98KlGLL0DKjGJzov/IFk8VuSbeDNi5gH/PGP1cGh57t7l
OnFCxk7wG6GBGKtNbKW6SYvngjvtPMdYgapwvElZBh+kiHTG4/CaYz8ehjczNRl3
/L3yWg712aSci8+n/yj5lm/wo8Y/aaQoIQVJw77Tkjc0CKhFAdbfcrINrPttrmBs
77WlxBmpcqqUMKNyT12a+0zI22IWwiNJepMPs1QOFWe3ovUoBS5wNE1ENp+VYwYI
3EGPkJDskZjEwxNQYAMPXKbR/ZoFHeeDEo2fj8v66xb9hZxMNat2OlgnReNa3MwU
5P7uAHBf/E/7bD9ggCgDQOaXryO8WajLrkNejk9nBQ7cy1uSsK1goiE/ugHJdMve
DTPgkoLXjeiPqKG3oBKl4BjqYBq0bSf/qCqv7Kkbd57R1faVPpPxTY2vMEJvvRGU
u6MWEhkdUHOf3hmFompXPulCihmU0N6kbVxWUnTbkpx4X4N/cBnqHMuIR9WXxTlc
hK9rMMYvD/z7BCBYKR1cmMwhyFx5Mo6fqfeI8qX0AHMBC8nQEK5tdfLeS3tFfjxJ
I+DbzdpF+MDVYlJpJn/jV454DEawCoLzA8aGFWPBV7/p5TbQUSyCM7Hths0IesSp
CumrCRjokMuNr5hSK2R8xLdQOcnlPXs8ryGYAdBKuIzD5v7q4OCsLCilfsrOCSE6
bBL2NAdzYxZBn29YYx82LKm9yMNXfgu+LODdyQTWjdfx/ChU7L/7qGGCLEJTf17H
Foka+GPKnMf61sbwnW8ELXo/VzAIDm86er9qiB4D/Oo2ncbsw6/aNHh2W9tawIAu
xwd+VtNDa4hxz4KPqXf6UbGEYm5AtNEXEZgPScPXz5xqXLSlZ5QdlrLV/Pgaofw+
yKNheMVAJaOIQWU/kSQlTgA+P/xsKcntaxhmnGv4dk98Muzl2CIvR2B/VFNTnYe4
CIRbLnYxPSjyQxOAC/UE+Mhuth/0LK6ZkPO06H8MGQIzRjgjOchTa6A3112BwitY
a0tmY9gahy7G+iHaMiURZk3YS7cP9BrdQx1/FRxA5ev0tULjnI8uNxFUvd5Cbwos
yfCQbM/U6aUtX/SV+L+cVdCeOGIVuo9MHJ5j9++I55oXG1hiPZa3fuVzbHE7tG26
qixEOxPIxlUmJ7j7FnYug6jk0MVC8fTRxPKfiKnppMlnnJy5abKMM2vNO2h3VCMv
0yAC8LHLoNXcBE9QJHLQG3oaOBlRah9H7gdXCsg1tlKMZtivSU3wtPlWuW06fjKg
Apk+b3q7q/OwvOp8Maf1rGg18vusBjGHVwhnBO6tLfUgvFF6HoIwIf0r6YLSYICl
sju1gvD72PdTFQ8CFVUUWDp/miE/baFcXMwZX4q2tyEWNyisOLOlsavPETjcXR0O
/nnrj9z72opbTj2G7KlkYpt8p29mKOPYHRwrMCRzNyiu+ArqHjwMyd2OKxVFxf8A
mFYsos7m6dEcQWugG9HFB+Hz/QsYI+TZdxNkg4jklt63WLHLzow1qU5DmhINZ40L
PrJKrPSvLINPc9Ge/0WkwC+3FYpzfWsLnxWB3QUUErZ074IqkIyb6smNffJFHNBU
iHWHuHoy4Dbt5awDDjq4GiSugJyWepQvjhezhfIuXv+Dl2K2PwMgNsSK8LcvxgUR
P2RO7vEww7w2xBuVoans6SP15ufH3NtlWwYZXFPM2ITorN8RKt1biMV+9yWr03ue
YlCJSixr9NkvR9Qm7++dmzAPQl5znLV4ct+IaNWIRWktS90YavwyVbOWgOe9pYrD
vQ/OS2Hk56Lzm8Ryk0Skbp5208sY2kJCIPQaYfzV+bNWkuiwlTsTtC0XFml+MxGL
ruziuNuR7UTq31pUXAGc39MzKqMt7GTXM84L+c/shIT4saYgAuEavURL41yy47sf
I22eKPMPPn6gLyRiZGG9m/LmrlrG61yIy8b9OLd/3IhwFmhjrQMnynWUT15Jel/R
RtLBEkstYhvtxL9sI5bUgcjHvuntGoEQqcoUJO/z7rUPwe1XPrmO2GYlBS+J6UIq
uNKZYsSa76HHBhIo2F4UGb6SGHyftlscpNVMvn40P/I6GelIRL6kQrc+TBIlIpV7
pcoZSeycD7bdJc5Xt96VpGTJejPxxNGRK8Hj3fSsE9Ks23ZBTp0UadIWUWCcx1JC
bBNrU7+mWkLqCj/ffNU1qWA3olOAm2FwX3++LS5GgU50+aUaCQt3Wa/+oLZCwzOd
JQV2900h7zH2svGylwjXXGkfafrqxCZec9IG4NZuLzw5D5M21ul0+A9omhHEoak5
OJPQ7TkXaBZN9J5BZVw1uwxLHUJLMuylsbO8wWUedcqrxgZ2pxWDKJA8/Ca1X9yh
A/AYC9QzYKYQuJc3WI87m/QQFOxqIBA4eKWQdVd9qBzj70gLE72sNVVXomu/Aq/r
OwpIlrWjdZM1G4lwwFRpa+cND6/mn4fVOOIlGEcE8edNfbeVOI9DMSkAQ6z2BoR0
Epjrcg/hxoa5mR6vcPvT+KdZ+3YbTcVxQnJP+kR+T2UJrbh8HeMbWbWxlerew63I
febIF3eRIrWJOGyfY+yYXgWZVKXzrnX+xZZS71IOXclEe73FfgMfIwEKf1X5E9EJ
jjutRk+G0CQEmCI1N3JOanfqbFKFunahZngqoJCKlP4/K9M5jOdYx56xZvuBNRAh
rSUg4+l65Zf7rzsK62W6ygz0YLZ0YyM+ZRUrjGzhZi0RwL9O9ohYs52psdtPKHxT
qr9YehaOaDA9cNKWwwSYw+MlleLupbNRfdahxtm0KrN9/cWgTjj0aOf8PIfFrmMB
UPOgnqOBKuEAOEb2sTMJ2Kw3w+hYhtw5HVdPuIfSV1r8nnI/4vshGarCoUYQvJYv
yz6JOZmaC/+5gju18JXlMeGxxga7YW8fqlOsy0KIQOLRpgyBvdvNvUjTiDFeaszr
LRntHuXbV6krYpo7IlTYZ6mGwRpOYbkZND9V7vb40DQfhWkDNm2XyrPckkrS8jt/
g8QmVb5fu0Tjn1OYJf63MsyjikIv7JvFc4cJb/wFYYvg1eDCrLOwVc2yd+yjFHQe
okIlXkn9jKS8ixSCA6uhX4wJVBwjdFrBCHJMJhWaQRGW04vipicgFXkNo9vL/lsB
+grOZvVcR72tLNoS+R+LnbkVsZvz+Nwk/q1AVaNq5lQpfBi11XLYhfIN1svJDdIj
1iMEGpq84Ay6z2lvlM8NzYjM5b2r5DrV7JLjVkJWF0I511mAu65/fmW6jN2YHyui
J7lKIaEJQyFYPWu1B2+JoTXT8r4OyIokitZ24DFJbeITN13+UXneFEaX2Yg2qmGO
+nYflOQ1fvDyE6cv14xxiAOnKp+dj42h8WgoFZJ9KmH+AXhPVNDY3IWiYH7rTT5S
+0Z1JCtvBiAon4I9dDUDv2iry2nzkS6zLGVNL35w3XDiamScroBVh+cm4HDcVOLs
qk2izdruQZ7rh6yTZwHW011U3BT6C8fblyJJqpBJiWKPSfQdvyAmvtAkbbiqwNud
+9lodTQL5rKRl5jNyp/iFJchfMEGbvWrYb7E7U7muQULOIsRjBI8JNnjH4Bk26sX
iXENFiG3O703IGfyVy2f9C6CemHBHe7URlbCYxvQiWLviMA6nbH1RJDxfMmmGK5L
9s1F05S07yANbk0kFtfFs8SmNBjb0ePUxKNaEDirMVQ71U/zJfqZgNWZwTpbhVXe
/svIdwqiv4IzKtTc+FspYkIy4ovzaxPswjT7+YK95sWxPS8VtQGrQH1a6N1tn9Nw
dfpt+6MIoKSbOZg91zJi3YGEFM9++e1KctX66Tub+5C0y/9x/k60iYl3tYFQ32Fh
YhRz085zwVHGIwF2XqGlkNbjGVAi6myF3jT7Gn37b7nZ7bbrQgfTKFW+zH0M5imX
kpp3HLAzqjR+r/vh8rdFPGMiBTfwwUub0JRXO/UbXUS75ZNEYcGZtaRP+EiEztx7
hU6MCMF6DINc6Ubzd/q3OXmJrfB/TIwMdZ9yO97QfguGN7b8G0Iz1pZATX2DVHQk
DMdOaFIrunOvJqwb+ictd0XZ29F8F3ZZuu6zDVnZNNRuw5mULRffXkcChAMwR7OS
xwH3/jGbaqemt4FtkISl83Df9U8s4hHJLfIAf9smBfczW4YYrJennIh+ed6fztob
NY+4TnprdQctMhfMMdTYOxzXdmZd2LpNj2y6cz11YcaLDxulA+8Humx6O+WnizKT
1WU9Y+vjlL7+7h0zQJzFtAoJ/ZbCqKXFISQB4LQtokBo4eK47xVza+dlrzvsX4mp
sVMkS1zL26dE6xIQa1F0v4EQUrDFA08GwP92djpwsx7lbmaYKQ4kkMPoNicbJ+9R
HMlmzfJFPIPHPiZqoGLSQ3bHBoFqtvi/5+3wBepJI+BKwDcHUZowEXx5sEK2NbX9
xTISXlVfPoekpPnjio6ZdHf705yIXm2PhwpOmwI7ANhxd4ZIcs2Ee4WN55YQXFQJ
/x8POOccZN+jkBEYaX6WIJcwT3ItEbG7bKDofufW+z/ZxnUvlZL1rsgzR16ssjyl
SkPAaeulmUU/vKDXULFfv0O8FZah773jyUp7gJJB/U/EnP7TqCutPcg2XtCt2euc
ZtYzVCcQNE9ZUJUN/wIjRbwRy/xEntOPK8EU+X/hR1UxHBakUVe11Gbt1/G8ESUL
HCLMaXEO2zsUd0cZhesulMPp3qiebkfGwo4FP+OTFdonJRUvKldDxIIYLbSnqX2g
W5l3fSIsKhjbCwL9WdcwRR19Vu2oR7sKQjc87q5pY49fssPHcx7SEEl4QKFCqMiJ
ye9ANz18lOf/BADIHrcGwtkOcm1eY5dP/PPKbDbXtN/ZCKbDSn4k4ZGX3lVHwEg8
VcDlfULbgiUbWKAlCJNPV3/Awf0Rc5wFjah3Ksbt+z1Mpe5xFLP2v8Zg6rRmyjvP
PmKwcKIYRDNYKlWJReNxJYzAAq07q8lUzyUaHpcZw76i+7tUaR+hlntVDQthegRC
dcxZ8OYEez9/SVU9rwqK0D1/VqknmLgGhxluWAR5MEb1J3OpGflAklu+fEesPVm4
w6rugiU4j3FIocGlnMi+BN5qHCdMZ5WRmDk6/dve6vUMN64skfmgQDNE5Uv8tWpD
7+qUVlT6wINrkSZkT2ZQajka5WkEuQWnfC1HO5aXxl7Hq3QAx7wlf4RX0pikkj5p
2Dz4ybtHPKcN/czck4jZyQ5HppXcWJ87OqjdpcJr0FogNPakxpdsu7k5lsYHGe+8
d5wHO35aP/0hRL7Wecb4coAaigB4aSI5iJDWY03j8n7VazZYe64ZRnN8tWQsjGOv
yFdm4L60jdRnMUJnMSDqjdhv/zhC29SKygCc4x6l9P/ff9nrsq3fIvp1oHE7A1k5
wu8Xzwk1q4Zrlp8v0c0FCDLf61ljmNQNNNKvrny9x0/0lSiF+w+WRyO6xVd1iW2/
xUWiuQpn6Z6kfIkWPKYoZnaIr0peWVLqKD/K0PFanv2wppSPqbPhEPVtigl2LUEu
i+bD9Ey+dXLn2CPYi1ompjxhFnh7yIqycbCvxEgC4N63LuPZ+v9vhYtmS28R/6ky
Cr1QhxlnHMR1r+ylGoUtog12n/S3z4MEBtClMLihCparNaz5oinC9SOUqrWynUT1
mAFHR3WloRIja7+TNwGRPaO3xK6mSRj+XVtTMJxs+Jcn2cgNnS6cxTsbHAAzkVSd
v+aD1dzqSGm1hLTKyVb85uE92Votzv1t2PAdBACzn6li8pDGlLxdHLuIO99cyu9c
eH1YkSNVcEEQ5plp3V6VUtF+I04fAS+8Frk372dwO6gUV7aP/Wrn+XBgv21v5huE
3qJrT5EhBjbn3HC2OWkYQT4O1JIfywiDamcxxTTOD3Zw/r4ppIAz2RRqL4w+WOM+
Uos/rx3grhNwaahTSPqUmLwNXI+7Q6NESSssyjPE9tGogbQrv0QNWZfGMQjfBI0A
VUxiJRScoTFq5bVryXJYI8veF4RRtNosR6aXA6EAAwAvPDa5xUwDTc5U5q6yA8vH
Tsz7B94msVPx9316jWhszHASk/3YTnKKKHMaa3R4xXIR1cFwNG9DKc7HpHo9zc6p
X3u4OQbjJALrJ4QnSUuflsEw7ptaV1h2ufveq6BhKL6YlTp7YUUqOM3bpALTGM3p
Lakd51nV59i0Suro96hZD8Mngx6RqUgDFhHbzd9X/kdnzxtfWa42o6iijpAN69Bg
N6smYwHS5mJnIuy9dlst7rnsEZ56rQBnneeE06/XYyab2vY477hZklXkgMSUabBr
gEjULSd8xF3/3LwCxlZQqu42m0O4oEK8rzeI/MNJnDqm/wyx++9sHNyXC/QKQn+S
lyZuPeqTCLczcLDZTtVm/g+oIHwDO13HwQiD7jVFOH6e5GpQp3alP8cJvdIq2Lxw
E53/AMhl9mZkdILNSZCgAq/LEbjplWtsBZNGTAq5mL0mC670y4q6PWar85jXUlr9
5/uZs4p4DjWyM5yQ+o8coPFMw4D4AJzsAa+MBkKMY2vHuvZqRXMi6tbd+ly1s4JB
gHP/HuncviVMCjk+Yz9tyisG2+Dk8Iv9wc/qRMFeilWqtwrMELgIsD9YA1IJuDaR
ygwVMD896CfcIxNQksFLGqQ2axgrA6INt50sjLSiOTAHcjgPRcTJRiAHS8hjHdkN
O3CZAaN7tZuVyz8FcFcUknpFwXK05Yt4m1oOsKpetalIFpfRbRhsYRbbBFdbMvz6
eRf/1drPeqfrsb+8caBiDDbMHMGQqv6n479XAyRYejzmzTC3GmOprZS7F16DQ/Li
j6JqMD8O35wALiZNnBHIbJdLdUL2jA7yRiO3YmY422lEFlA9gOW6XWWJU/DXWL7c
DRDGdn9b48vAlqxf006zOUkq2IYoHJM84Y3KKljz+Wt/e1VpNQN/aACjFeJIyu5/
qVxc3OLy4dKRJzj5PMOzddP4s9yTgvXTzFQhu5t3IAyueixi8WdCzRoZ3Z7jIwa0
v7TVOQQ0KYQy0+wKLrKE8Mjir5Bn9t0youFeJrZytZVPKjuvhNPnqtEbS2oCV8rt
/l7U13MfKfBCKQ9zA38tznFJ883fxd6ZY5d3f93B46owpcPUX74mEIRY5B7SY6mG
DmYfERkLg5lbSU/9ZVaCGlsYJ9BST9zFG0WNEohj25JbySarkcDTBde5anv7zVa4
ltk9bRdVYvp0U+Bh6jk6GeUCJi9Nx/L05Y5B67soMfN4VAh71ORuTXAk8lhXvvAH
kRHNnE0qUaWv+OMusIR46syRCp2CnaOfy9Hlgz3+Un+JqOO3T8/Z0nYYGwnbWcCW
rs3YRMnSsajlGyXeoh2BkNUgVHQSS+LRuoHWUXJYOhdmDnoad5/TokIbTyDRJPL3
BUkfTV4EtRBJqQbkvYF2/gT6tMUKQDobgc+OduMAaQwvtsFtzKcIic5V5YcMr3wV
QpxW1q1w21W909lQ96ietKXOigiPNW800xBnpclCgWk0DMjuw9Zfbr0yj/Y6yxaN
nKLhscPXL4jlpbDZAQ3yJUPyD3CiqU2m4+qaaazxeVFenURnucGO1p62YjSYlWkt
zNgh6HIboGPP+nMVfVZzwdxLyTWD21inP3XDu5qLtJrnHAJqCvMCaxL6hzuBwqYt
s1BdrGGdMvOoVa3iExe10j6ZMdU4Uq7d/Ne8qsXjc/1d2Ks6AuAPrTaRRasUOUha
zU6hxCiyKn+e3Gn4JgtHAFegLyOPWxnH4/9ewVGOJQH0eB0+YtfAmUTtsCq5axFx
WUPeLYZbynXK1gQYMHCU2YCThb9uwvA5IBkHKGbARsJ3aDhWVnCVGKGOVrrRNOIQ
9ReYGM1bIXZP6DrvEOOq6zp5yNlXfFZszvr6QwsLZD27x7rLJTHEb77L+wIDOw2W
fyEC1mgIvL0a+ODjyyyh28kJne4Q6gn6wuQXX1nCSnZooZurT1XuzszJCOCdEmsr
UvNV6ZnzqRO5nXbr9CcpCN3FFztPEkTgWLdw8DwUDzMp+eYLvq4iSyh1sIv0EGGY
48RmM+nH9ESe9nd/LqAKvoZUduyQtXFqhtcFeKlJMbqi9CtuBsoruzkNkHAwJAgy
69XTF90Xwx0LzVhobAMvQqGgNxBHdJQDH0HRA7n35zC6MQZVwsN4lJiLsdRVX+m1
rovW6cYZ+0rGham1yMVsA4AQq2At3uKo7yxajZE+8AeKJ8CrSSw8hJUNK3V3QYix
TqRK85Cj7X+vBN908K7YQyLlCNZ32XiagTnqw8X9UN7nBTRn6IpC1ds3/VQx8vU3
8WYXHYx6G8kTDAJRQVjTjJ7L4ntOYSRCWmA9kgN5mC+Gz5Ss54ReG1AyBd8B8TnN
bnUX4P8xxbDWrihk4cjX3uA0Tw1mzRsfa1Sa0SkMVcvY5RFcbq2imzVwj/85zDJW
fQBB956dSKVwIyKXSERD3ExSCxItZppGCZBYwKqbsE6h42a6lH27gGjuN6o0XNbV
Vx0bpKVWv6pESM6oYVpT0blK4RmdDcHm/wpQOAsynbzu11Yc4eegkmIPgNmnaQ0X
PlFgpZRPNyYXeMMeVFgl2wVkYbrsbLtlO7M7vYaAem97ZCE0TCSu+UHvYNVdmmNR
T/7LUywdN3+LqEqWlUzZYXwld5u1YHMqJVGWhFw8j8CzWgrqVqWp0jrzjyZeztq2
QA/n59FySUXTpBCHmrXZ4PVIwez3DpxD81LG70/HArmMNuq0k33S6qzyy68CgrLn
O66PTlOJN08Ell+5rQTA8gDztOdD00SDkwPIQ0lAMcQq0RWij3cgsrXb2h1yf0U5
LNpKr1jvrFB3gACyDDuvffkTttfdjn/frRgaVmYO7+iOvAoZfbHwwYmX111ELiNp
vAew5bA1QwxOB0NLmusgyOdVlGzWlTQNXs2z+O2EJPIgdKJ3hQnwZEAe+HoLeueY
7MmZU9auGeVdB99VSSFnjC5iWRNsz6fjRd5lZlbuDZiuke/p+kVa7WtCgWEhcqe9
71uNHMFXwShq/8JpGMuiugAj6LUKnn5LAIt6MhiAG77ULndJ6dOmH07kt+hEXazq
iDkVE7adIv/7HykfVqMDoQb1Zp8lNkDjQXaPsLf392d8IeBIr45iwNN+gLcd2M31
rhf/CRZbGDPgYToCcxEZB4MtO2L5Cdh9Z7F4NtYqZoCZshphhRYC0mJNJs4f8A/O
E0vKlnrvmO4/0yxC71Ftaa84dvXVvF/3qnfVOhw2Xb7ZMtRw6ya1vkvMOnZt7XSR
T4hey9YbkHYy70mwGgZEE0DVJQ9BDGHjYxvuiGhVxPy+XW/X/nnLGs94Maxy66sv
imHn+SzXKvH5HruRWoJg0RLfsaMxRQGctkicCo9905wRit8s2VAPurMzSY366ur4
6WHqxv9bF6V993PHmmjKl7ahe8MVMxLN4kutByRSL9afMU2PRvg82w8eE5gN8Ul3
GrCNqU84OQIQMtZvVTGpOcmt7tlSYehoMr8TTAsYTW/xvBBhzxu8QB3mo6wjWwtl
cWF6hLQ7pU69CiTsxevFIot6LaKc55ae+bnOHq4Eq5TzOzA6XHRJn5P1TPx5GSF9
eZzBm83FA4gYKhQ7Qmw4QmxkC6GfbOy6z04GVKQmEVRzgKmGaUaSEdZlkEN2PG1U
8m6cq2MX/r79Pi+F9qNcZ/bRBSdq+ZSoBSgu2XjpNL4alUVZVFIN0O07oLsWxtGV
LFxmi48cE3qpDVotaoPoYjRO+uENoQB3wsvfr40sXJVK6xVlC+6ME/mfNPIWTztM
YYuI4DieiInFw0Q8pSvCw+/RApcOwlEmWJ3qveuw4cZqyPbhrKKQatdO6BBvF3VJ
GLKVEdOOOhrBikwtuJr/G08bFCjTVjxO98CrLcPpF5LJ3ZADouXXGaj3Ftakagzd
/M07tqw4Fi7njGcxc3+t9+XTdNkYH5xOm/ZOmCHyJ7JVJ9wklsuBRxumaTcSSt9v
f8WpRlrUjq1S9aacsn5j2BAZb4ORJXPz3PbMxvcHL+EdPc8qoW7yyI9ZdA7wSL+2
MAk9m7U8kEZ5hNJJVx/dDUnaR8dXW060tuRfMw5DfvxeOcfOPIscRNmW/gY+E8px
1kmev0p3O02ofNUnl5qnIdEQHvv+Wy1W9afPD/uwpwYBJtrV4BHkUf5dTUTn9cbX
ca7/LSAkDOfvQE/ABJFR65gG3f0wTYAW2RGIKeS0auFKunTBOKbb36MvFZVSdd41
J69c21rMlAawfIuVXpA1LSvWKf6vCiDPMWwrN4CAWPzq52HqYVqt+7lvb9sgrfMt
ThgnNA/Wfq2/ythWiMr20pTF2W2rB0ZcN5/6kDU40692hhsPwzLKhK4TX5x9HUU4
vtDllv5DAeVsulJuUEKrJETiGMvIVRFP5nOefXzH/dYf29H8Mby6Y4NpY4EmM4it
8QBc7g3x0XSKYjdNnm9ppiHvSYAFOla2U/N/sfoEw0bV+zWhBp1d3OfL+gY+I3dL
TYdOqxHr5KiEbtO0kRzcbzk+dREGEI6r6GtnEFJQzxGPPx9T/zVz7A7lQyTA6mPn
nycQxnJ3zrNxSJ7QqX1Vqb4GrqtODKH82Klu898ZydY2jt+GhAwkEES+80EW7gyH
cugH3/ErntFgBJmfm/tZ7IJtdwcu4bLGfN2Ov9N0+1u6VfMzFwQA0Z6ipN6VbjF4
jWDu6HEUWZwHM1+MoSA1WZrGQj7MJ5HwuoTtMyrY/tizTadVlz6wgiVqROef7jLB
P3BGvH+QSwBNffpu4TgdnqBcHKfeV3NaPKOwI1Rzl68kPk1T0XXvZwHdzeKVBTqJ
/+oK0b7Tg97+JHmMK//mKTFbb/+3EBYRZt58fFc7X7w68cixT2/8aDlCJ3Ko2FwB
b8MPpGZGoRkXJWwI25PNJxGQyRxuD6/HinrgHEGi+T3f5oQCFFe9ffFRdAJtnoxT
SgO3TZvWliexKx2z3XuI8mCwC3f6NSLR+EHCoRhl/P7Om5XNNBbq9d/vrEUbJ2V0
lbbhUW3mYms5qSL+uMBOx/JJGJFYKi3ic2Qbcwbc/g2K+8dMpbZKOBob8EiKuD8k
jMsKprKC99FLpJ8uqVorCgibtg5HOpTpNePDY6A8c1uJ6BXQ/wnNmqUYwGZ4zKfT
CnJBgD+v5XPIGlbgl/lrHRKcux8UKe99zJ/MyEQ/5iApa7ugcQ+v6lWi3AxYe8LD
QbrtIFTSsyb09dV+aqRgzaa6BDsYOhs4GFjaRpbUHkTMeTqRSuAnW6tfwuS7Fq7k
XztR9Puq0zs2jP9nHv912upPWIQjBWk9Fo6ZpcTLr7tUco3oowwm++ikFXjD7S6w
v6WA2dwuuHel2YIJXqLfbxUlU1IEtpawl/WHLBD9Wy6tQIDtGtdkzYlThA6zWKd7
nAlJ4FTBIXCivScZpbO+ssiLhzI2e3z0iZlPMJbWIChDwIT7QIfcjBktPk5QZ9LO
1Eo3UWpZ1/+wdULm5TaPQuYlZ6grbzxH8RbB+NnEGde7ZMSgrMyXsWmFFpAKmnGc
vJkTjcmtc+eU74Wy2ozsRRF4tS20cO/Pm3OmnVZBWn3qvxYyyVLdwLLK0EayvYm6
y3YDCrE6NLfuppYvdCsauZs85hW84IOyWCC3iGUUN2b0B6gKV+3+NC9VhOVhUu6o
1NWDbBZQGGPzT7XRmB8Yt1WilUV/rzePwrCRv4B/wvVAjP7eWvzoAucuIE/25SWd
xxE1Dk/+8juPvTC8h0Ust+1a0ady2QEDzqWQNOuhKaGlZBb1oD50ZdcAyL0qX24g
nQ5PLvcPA1eIYRs8dp7U+4pRLt6GepK7x8AKspSjyyxRju60qKAY95sucO35dRuH
s/2r8nggTBAV1pCvUkLV62rKvseL5x1F718ms9BEVk7Wv2PvDWth0yNbTRI0Z5tY
g2mMIG00OD8qGsLsi9iaoSHIQe4U5RRQeHPCHHfEL4ZMTlkMii/JEKSub+9EXtXb
uhsY8+RXuGLig4BDA+iaLqH511ZlUkJFrtiGxC2GzZUpNpxsF1AkWMO5pmODfnXJ
JD9c36O9Lad92VoS2KCCFYJ4AD+dwuMvqzohgDbZE2FMSdlpGyfVS4qt78jcLD4K
/Pp72+n3L+mOfmr8k9Urh5cfMLNXWksm6Rm/WzgU77WmORMuHDVwY/LRVQxprx2n
DzYGB6/ZSSjMca09Zd6OKnow/O7HhVa+5Oh12g/38RNDaqq+wH3gFntrsxIVqy6I
ej829nn8wcPcgb+biMmNsTZ3wJ95kxZXiPjTOb+TA4gsL035i/M0ZATMjU1m5pYz
PEYi2va+3AuNsdVTZJxr9h3OPEjSrR9v/S9KVLAJhFGtLe/FSjrAaxMRNJlePjln
y2zIbj6ZT/Lyy33aFE6OOoc/Eq+oOKDckIPjXL4PDf1vxndrftTBtj6VKMQmVF0w
cyihk4XDJ7LI4I0VA5dfgCE4gJKWG/l1TY52yAwmUPu6AG63wpMEhhqvsgbH1Zus
2hwPXrj82CoPEv2x9qFdDPRBQZxYggzew0zZuaHx+pvbuktqRPzRLOOy4IC3y1He
tNcHUpSRiXV9zinoyA4AJKBBcUt16uIiTW7CmF6MH/oNJ+SLyWNJBj7dQkOAa/2h
gSILFgGt43dQlHPEn7Yss3ziumEjOfqeoI1OTQ6pHq/gJ2vUBuDf9yfIizZNAmtM
Ons6QefbS9Kt5fUZOtPE2n1Jl6+Z4vFjCOa7Qf59GuI3e/y5TfEWuxbN4kmnrG7Z
JMHDW5nWu4kj4u5LE+RuxyWJ2Ixd1sPwA3vq8WMy8iTI/sZc59iTGU7oknW/TH7G
hoBeB8k0adZpC0aewIQXJ9CPDU+H1aFX6ZhBvY/QXVixoYyYbBRO0XExVxbUchqF
1mxg19/1v7xeDE09maKyf/vkVBjgu81KGm8JyO9qPxxTjfzST0qGVcGNuZz9Zg3V
VZ6Yr8mK4wVOnDdUtvAnX8cXOe6W3tBWu/m4rJjjHe/creBfjeIOVlr+C6yufEkQ
PaR2JTwzNxj18woYZWF9OMsQxiMWYvSfC2QFIVVVxNJXt6anZR2iptmSEZQl+6W9
WLRqqNU58lBgV89bmJ8qkUKYws1xXYG+6JDCb+SIn/VFQJTuf/Td32lHwqHXitRY
fxCEALg1YidB0+pt3ql3lii/HJqFvazl1jzvge2hcsQLYudIY+to3U+FdSWIwUwm
AMP1MzhKv5UQM4CzSfCHV76S1nBwWs0v07h5+R8ZVIHPGOe0mawptcp4dVX6LCqC
/LjEZ1D3IZz1yjAlfzArijFlfmYeMhQM7eOuGIP5z2N9jH1C4VVbXzXTkphLyhIA
Xzn3w/nq/f9Iolbt08Llc7SWjuMk0sYS+ToETW9odPwu/yigQQOWQ1vV+joGH9BO
mmUe9L+FIH1qgd+GQtM69zLRMes2f2bpejLOs6Q0w9dBRSeAjkUEKoNAXu+rN7pt
yOm75votAh/zQGwJYPH75cmApTJ4BvzCiB5D9E/sgfXhkUtEfspy321csS8xPr6Q
iX6Bh8z3yOE/RerAc0UXqI0GMDwxvLFOk2ERWeFMwujUyzYZ7vutrH4Qz4+fHQV6
R8KOxGYWqbqDH9X7MJ+MclPlkTZxz4PVCrQxj8BVWREpBHdZoo/F+9fTYCJhxZza
Yz2dmWyfQD+sLTaVb3CvoFUbZtyph2aqhoQyIeXz4lN2k4tzM/rTJbDsfr4VSNQc
SQvNsxvbkfndPtmMvPoWXGgpJDB/qkjUuz+wIDPTMk5ycAiUtXA9OldI0T7LTKth
51vESYRc1iBvUQhZpAUNmTz3GSXCVIwgHYucNZk9PgYz7RYe7CVgnB2+jx5zQ2a9
NQIK09z+ODyh7fWKWhr/dg6CystlCAf7C7UJsh/IZk9/LUn8/s3VJjDt6ccy3+0t
UOynRDlsItvtUYzBLfe80cZwZmBVZU+e6hL9gEOlJEq8zamrfxw9UHod8Z5Bxas7
wn8DYuLD/DUfkMp92sfI0tRUYrfOSLyb5OQ0DoAJViw5Qq16vSuyxf49yOfcBuGj
WbdH5VDHGYnrN+RyDcU/xvlU+nPLI1/Yp1T8Ghzz4cFSbMvH2ZbKax4UmFQ/4bbx
2VRZ/sNwuadY8ZDomEb2LC076tuC8KaSie0MMNfOFkPSg1jYxW+0Q8eYRTzoT9Or
VsenD/7PDldl9TOyyQRHxWw8JSivqL69EVtgnw+bNiVEugL5vKkvaIfeIJV5RBbE
OjLDdLZbb1WOyleH5Qwb/PMJsSL8eoP5cytM+1Es31ZlHyeV9xrV0QsYty9uMOxc
vIMQEm2yy0RhxaIPeDqIziD0jhAzlafQ8AWMt69pC+1WK1KLmXKRnOJZwwPMKrYe
rPO/g2l2gEquVrU/VNo9MrZfCsQJ8Hhzc0dJyt24Gi+JtbUKgQ6KBWru2EZ4/GHf
WTWNTN+nNSr5WQBVyVsR+FP79IV2fJRFNlnqmfPpqKK4K92ru9XQLnbmA1crI2Xd
jKjBxq/HysB5kgj2ra4t0FK54vUgdOPLbnINAnJQS8amrGs4Ik7uz3xtxyxgjL3z
GzrJF7w6y0MfJZRapfIP/w7of1j8ZRon8eGhKpyEY2tdgBItoaW93jt/7weNRZIC
wQEAxKrzxqV62DtYXBs/TLAoTzozLyERXzr5PxUOoMrWqau0lqMPu7+sIdeKimjt
g6gNQlxrI5rQDI0WH/EhcX/bD0ynqBdlgmsj1IW6hq1jRFfO6KNMoRK/54TJGP1i
AR2HAnouV2gPFOObscemfkzXA/v0CuzY2245l4icDZ4jvuLF2gPPfd2QnbpyCex2
Q7kLVPYcZ4kMcQMt33ZmdufxU0t+lX4NsFuzYeW2GvZ/dU6/xqVmeq+x3fqWD07s
Fna4yWCxNDxZlL4EYRvmowncFHsOqFUbtlyiF/UYuFh+o1pGNrdFjgwCkfaIirjm
t5DdXoJXDxysXsAW3vNzUtnX8hx2mKduH4Xc9efFnZvdcCtqj5W6qrqflVXH15jX
UMf5nnYv/7kaURwivEnBi58h7Eibd2uB4UAAXECgnOKM1PDzFf1UMizINVpaJXkG
68UcgF54Y71R4BoVNKU4yVDpY+o2NuvjM500+vxyECx8TjFhEI1O431EvIh5BJkf
dlKuZnVAt8RbMstnDtFd2D/xE40M4k/yTHvDznTTALuWYJ8K9Hh+QR5VdTqkoUnP
E/hA29l1w4fWf+iDZXQnvYreog0nrqdBb0BeG79LcNu9hrMtOidATYw6HGxGIbzf
LdmxFJlc+y1iLgtr30RCaWYJfCiRDUquPtNli7Z373rn3s4oqDS6I0XvR03g/cKy
w17X6Wv4vFN96tg0L0u9wt2cCHZxIlr4395FoozYFa0IUBoaxoSvVzMBzBHXx9UI
chsxTIE53bFYKSSKoMdr5Xa3HJYFcZVjThNxQiFT4WB/oSt6n1Yj2LGUWvkJfajD
A4FLvC/k2YBBPlj64HoC9SavDI8ll29+uixsQyBcrOHq6GR/5ut6FEL3BaE/MmYA
jpb8RiuzngyRhc2p12uM/PiJs58ZYHLyE0CPoVUDigqLoUZ9qjLZYn96fo7kWk2J
bss9uZ/yqzbKfPplyFDtzApg/Az9wO7kbUP4UTToiAH8hCzCwCTKYzjEBoVIn/sE
0CwC9vhMcLp9mWXeEG2aCIJVoRSPNertXnaZcuVnpE3nprn4VERhp0xX+x/JCS60
Doiff7GLnSk2aKyI6y1zStoph/OfR2F9+74g1+2SQoy2vpdTqem59oBLnm+g6XQO
rnqz03O2dJIS7JwH6AvN43cwccmLvHw6zjnKbSju2tygR7vjvtRQdkSRBELKABBw
7PZDcUuSo+3zdSkw+DLReIHEWUCgVqZUPmJBeNrHVN47fDSQ0FUA2hEbV2809Ynx
nAjK3oYyDB00mm79AYrFC2HzczgmdX/piQnwL+q5G0qI2jtuTHB2EsZbXTZppA4W
c72cEVMK4IyeGbce4MI2kqdmQgghRptI9iIxsHCfBpLDKyedmHiY4pDerXBrqtfe
z5u7t+Y8K2Tn8E355cDW256zl2ujEGnleL9OVfy79IoNh4PqO7jxQLAVvB8q4cVz
VcbULLENNjJVWdk5SxzVueqR/rfjDHO8hlPMR7vp2++sQvAT2t8FCOxBf/Ryqtao
dQhMOz+/20eX3rIMEf7U/dfq3uIRozJvHpd869Ava2r/0itY2+dQdFajDek44ZBB
/hPNwVIsq4we+c7S5ZjEddZML/Ffl6VtOvyZd+EklWV2Scolm6aoAjNWIlGVdfXM
CzoWSe9CX2I8TwBXwFRyE1CVi5xdLIlTiIXZxCCgxG/in1wRK4laBfABOQQBkRPa
pbpqEQRSmuM1dxrtlVM7NDNDvdmNqw8VNk/4CQTKqCw88Z05qzyAUG9ZKT8BhB8f
ICjR6l4tsa18S5sSdtxNZJfodzA0QyYwKEgRF7LFad2j9b6dA/dwoRQDrT3MJPc3
v8TpXuRxhEA4V9xpTDO91z+crJNxMFeKjhEbt+bJSeIgG59nVpyRgDJajpmT2Q47
3ywJWXzEEMAA+yDFjNHs5jnBwMwAdATQS4wcSld/oEIRxEXrEIKj4fXzK2bN8SpA
oK9oknKqMhCdW0pCeKRub3yL4vbTIuSOCU1kmECZju01viseBw5DVxTepk8G4jmz
8LG3g3jkByK73o2FDww3mNyO4s0RbSGcjVDEHTRPQ43tioO7qRRNJETqIGaG4Ndq
YpIREnK+M8TmAFUxSRnHcD0YCGki4zxMPSO5dl8rZDnktUdBoRJxi7bydIlfAvuq
J88JsyqO3i1JbMwoogCDIVoNz19kxfkX0Wz8kkDvPWsMxwkGSJ09Q3eu+5i7yh6b
xNtr7ClpoubksvYWK+JXFP8zfKCB3K4ETNW1zHgZnB4H+s6ZTCkHcQ+/4KvbOD88
rtZ9ZXknrMN0wZubtdRN5J8fiMf+rJLge5QKrB5Gam0vgrrCmSQRR9qKZqPR7Rl8
2mpKkRUrUOpJVIxWClaT2d0UTR3FkaSfWAk/cgHJJiHnKhXHoLtTK4nxlbuEnURJ
iWmqVOtNuLU1lRNBdeLYu040tDZ0sBHci7wrQHMxPV0FL/M0RxiQb4Ak5km2L3xs
pXyTtEag3hnr7F1yA1iJoFYJtlKCjOM1M5PPBspRhUyfqg+yyNIQKmCCTz6xPWBz
AhMGTBr8jK7Ov1fB/OsspO/5wb4ubE4Gdh7wRDDZBSltWBAoYeNOS2BLU5Dfx0nH
arhngmYWAzQYsKCLeCOTQPU7tQhJ6rTwcZnPd2Z3BpufjWgtcCtkgaydkRELlLaw
aQlqvS8pfjkd4X9efoYWkopwmYOlwOhMHTgA1PiZFUnnxou4Jnc4+B21EomnMmG5
wM0DRZ4vpRlY2DC7tLPpuLAasgg39u4octliinXsNipgwGNKYBTFIIEy+BkTw5GS
mXKnuSmIDLB9afrv8JOf7q9M3QwOpJ4yVQJ6i7095oiDHbSKh5kI/2yQeraVXwou
r1WJfkkokXEWJVRsMLy4+vMGAW94q3gr3ac38RuCnc6bdqcNAnT3G0hQb8wLlpRE
kpb6PIbXxLFW4c4aVY9QU3+jeDXYiTP0rUdkrRhikJhTHDkWQICetclV7dMvNFil
hdvkqid64JYdfnoUMJ4LmJnFSS7J+glz+g6EEZoyvQwRvYlC3QSVx5CuoEgNfj2u
ZXL2R7BMqqOTRLu94Eium/bWaSpIKkAdE9s233/MwIF/apEhboPmsoW+c7pGMGlV
i5zY0xKfN+2S/nLpZBR3zIufp9viTNVo9/UeJ0cIBHQEsYzGv160QUrnjEna/cS2
cUwYOuHh7y8/r0YBD8/ihWDWF+sf7b8J40UIwvGq/5dxnat9y23ix3xE/Y2mU3qY
hWQA0dNIHxnScRMNv5Rmv132/6ZxDUiNuhS1SlUA9QYKlCh2EtfKvK38c6FvNx1F
EB7JqJb1FX5Pa7PyqXoQoqLkrDjmAYfeksafQTZ8TJZMGAUdyNN3GJy45HVRLsS4
u/OG5DqNqAoMQc3E+PZhcsv4aRZ8SVXZaPba1AyoRRe93Qzee2EwLSo7tI07pmF8
9D4PCjm2BcKSAF99dDR5V0sd9KBHhiZwEFlsGE9Km2kTRh0gBsEDNREztiM+EQ8F
NPZQ6UTeV5Jxo1RpUhNbtmiFhD22M/alT9h7v/5Y/rwMRN9fffvwb9pKlx+c8VQk
rSyqamiQzhExj6pXXmwPwP99i7i0XWGtVDSvtGBeye2yR7wSKPvQR/44fzcnsDIi
BR7BGI4JKM6Z+4gi95X9H6Mj/atZKzHUcHGqRyM00Wc3sM9AkTmAkCSh5F6+7cSD
8HJZl2qSQYwUV/AJ3z0Pk7QjHqaIDQ+Ra9n/oSaMXGXnFkmI8AXhS/c/7PLqcGNb
YmIRjeGFbO2MsmxMl+RnMAz5Q0Bu8Ah2uQtrIv7YQMcbIObbT9JWU0HPp8r+/h/1
WEAgQxNQunDyqQ0EN9nl1Pi7oxSl/Vft4uiuRoKovil68opx5IP8GXFpOSMxDpaq
NyCsU/hP5A25h1KSSffsYiA7dn6RcBfEwA3s4s4efBMfmJvk5Pz5Ny7liCkt3thj
QmVYVk8jwpxwofznbplx8lab6lq2s48PlyONJ3VOVc4V9otYIx0Uo2x7IJkgL6IA
EoPB8/njijB6U7+2ketqdaO/T4TEyXzYTSwstyPnnzuKsRi1mVaAxH954OtpuZES
yTu+woapq2+vjlR8N1mUOH2Rmq0r0L5C0zEIBO4bdPTSJ8rWTgYvnkdMJTothy87
UKNpo/McAn5NtvTYpOm7wybStH8QjiBgQesTzkUekuvKoGEwxosPCI40d+3dt9Nn
xA2KTa3O7DMd4sQ1wCk+RVhEN+DYerwV3qqtjTu/aU859O7rZ5Tgx9gSaBjnoyq9
7DspGOCIaqum9vBfrzOHtNgoHbftxuXaQtXKXkwrMPFuf8favtcwOLodnvrsTw0H
5RBjaC9y5kA9PhOmfY/pq5cevEH5YvyhN9tXlsS/lwO2e0zNAnW6UtNE9aweF4cg
EDEgZL5HWJg3yweR2B5h4aj+x/5RK2AugkEM/905Ad1EO/yI0vJX9bjeI5B7Pm6m
W9qoNu56zkFsM9CbMI7eiugqneAtrm+A4mYsoMRjvJpigiUngFUHCSz2K0QPtCxa
oMEB6aW2oKGtES2PZb9HZGFsn3/HaBHBop2Lpf7ZaP1XHqyyAF1uQGSLLQ2oq1BH
u3ChDihgp6Qwo40pXncIMB6GQsrMfy6UB3z7cyZhpbDBO8fVl+DhYoYSGZGS1A7h
03sxSAav+Mi+wBuAKJbPhGimO6awhtBD6ORPl9VYyOOu4nss7PH+fmDrhcStKv2i
geXHQZT/nk1t9x2RGTaECJKxAa7FJu3fcfqkXCAjrP7KMUWVr7ovKGq/723mt2e9
igWSPuKDPVcAhcMJSaecaAdEHWMLdx5bguPvNng2IOnU1BLvnfGQb92RrqSAYEsX
QI5LMgi1D6gQmF+h2PvrsKnZHl3FngDGtUygDqNMCEBWSyJdVyyhq99bdLP9weuo
02/LqNkDs2cFTGg8qt7pgki96mri2QG3l3vVFr+SFy8lrbNZRRZOW7h8eTPwPu6o
JOnS+w1qSN/tjIL4AGsnN2ytm8MCZemJP842aGVzygLXfau2HtZVe6oaKm1bAYJE
DmTTQV1oFrlalJHkU0S3hKyJ50hFse6KFJ66JEpwX6dbCKJhAJnw1XLa5ak0HU5G
ur8gZWhGPof7YfJvLUCD8jnmrd/7nJE3mJhBNepzp+fYxIrXw8sOuXlIExF6n3AE
eHtByloDE5psrLlYB5+MB7oY+YbMZZY+3QSagqkld6TYzrrzPt95ZoLE7NZByDXn
PhRumBI43nwd6Rg7pQvtfTpBLRhRM9dE+d+BrZsbPC4psZzmXuoz9mZQGSEkv1Wl
6o4GISBtz7o153pF1xkQRlPAg+qNhjRCdSeoWi5WRniqRz1aGN42yj8GMuUt5iPH
TTVvMlPslSqRBT+3xAi1iqsgSKURBMu20Z01mYBzZuIbvZ2kUpHs6OuUCyG1/TW/
frY9I2AXtJ7cjx5mBGYbDu7iIeGf6s4b80YFQk01EYSZdp8oENKSsZz4YxHSh6d7
AmvMU2SWbxl4O12BpfAf+y07m1gUPvpXa+R07oKSjJu6mOn4TlZLHtg6zDP/08Ys
W2eujzF51cLF8xqXvsW1f4IDqJ8/coSWptM/UVZZMf6nyA84oh0oZz6cPsCOeQz4
fZJPt6zC5bdf326dO0UR+Tm5ACE9NWHIPeQBXP+KwYY1/UiDPBpWK7Um0Tl3+n8J
C2GeJeTAujhtQ74wskZ+YBxqyfLT0pHLvgl5lfJvQ0142ZFoVvnq2oHFQEVurSZE
0eegvlg4dgR9/rU+HvNqVz4ERGMyAhguk3TT19O0NFHtJf6LN0KgDghmxsrxM/SV
NkJ09bBJszeAGYBb7fy3hG1DImYqjCiYWPwn2HOt1VQAIjYQZj0pWg1VoWXM/Ehj
okjdp25ElrHMwMglGXrTbDfpiQMOJt47DJR9X9/+zcsVHcSXvA5XpiMgwS2kzKH1
kpGjubmhSQvaA26SJRiILvegx1qIvr3nvbZaEsez0gOYAfClpoix/+R7Q0UqzsdH
99uK07v19qqVIumLok9uObPSQ2eCiJ+Kv0sOqwslSzfcYglquZXizDG2wp4LXTwX
qWj4t+7qu2ziiYJK8Gxs9cT9W2wWjj0+k8Y5RYdzq+DBeYWU6OpqULp9WylUlV+c
ZHRHxCmbaIw9FTM6GEq9dxbqgaoQN8IqEO02EFtjCQ9Z4B+XKcKW3GCy6t2YsTUt
6gPLjE/M8GvA3PTsaqfsrGxlyS2Dt7lDINxm9fJbDrEyPZb5/jyEzizxlDZfEh5C
4VSILMZtTJKhhDoTeRoaU1QfA+sOH1vcg1MvpgmSHmPVeWzXrzVGwgEF3u58ivzX
uowNFBa9FwZX7h1PWAfGt4RqNv8Ek4rPJwxcO/US/QfvBWngXtsXgJQ/9aXLSXyY
m5rPVketDrbLx1rqFrluOz0c4TcVIT3+V0UUbk70pPPl9Ou0mYyownycZd2grXu4
aE8f9qspWp0fO+f8NoJ1OSVxO7nq6ysFBSKj1mu6/UWbX+oWh3CcUlPNPPoTEYvs
89/58M3YsbeQpI3JuTlj5l4lRCorI/si3TWKBJtRXHr2sWqzp36td6c837y4l3SB
jSqbhGuMPIHhbxkuMIT9tvTRGOjANKT+aKiSSapF94OBzBpNchwPm1WB3a6ehBX0
8iWZDgdGFexRNlgJo2tel2FQpju3RsejJ+Hq6hJpuA9kwJlR/A/dDrXE+iYpgZSh
Hme2PxP8XAzEXp1cmytHnif2N9p+QUrvqLAuKPfreXGDVYwYj/7ZjJaxRv+vyDma
DYknu9p+RJQy68GWoagTACK8nL1Be/1V5jorI1duYbxXdDaTJszljOUbY5ICKxFP
VWS7Fa9sjlRJ07IS+RLJNgvjXxGCiaQm1l59WDSw9FArzYMDjPJ9YCHVTjvL4TX2
jHMx/NsNXmeCYxdbogxlppmEIos5jRgAJoy/gUmKoJ3P6WjBH2sbS0pk+GkUI5RQ
+5dzyjG8RnCIZ6cs+AtCyotCxc8Vk9eOAW1Tyc4sU9Bu477lnU5DqGA0LmjVboQB
Z2RjqThJ5y9gyHY8hz08MuiDy51MoJW6PIKh2dooJrWsfzt8KcUeD5+r0IpDkeRh
BpCH8oBXbkqCANEfAy3p5ZtydZy+padZ0IHex2xG/DHc2QI+lP98xlhOBTKnSg9z
++bifAUdWnUGspUYlVcUeur6KeltozzF8pe55CCNJ5Cu19dvZEVkeBxPNxgTHpkO
d2HhwOhGuAbucYdR3sGoJsBHwhJK91PExTM+tBk4KkGa2/wogbWBvTksEt20kBSX
VAJc0+ORGzeTNxffEso1nes7pT1HmNhBMhWoKovzeBRi4cTu0dZoqL54e7mcyjaI
6WFdRFPv2EtR1QrrcinLNKiWfcbPtKaryqC0rdXrE+RCYqDoZgo03/4TTvfyueXx
A+vbifZGAMYh3d5N5h7HPfHejQoeEWZ4PUCHi6DyNqf5UFixPtCoL1EB7mmzMIgW
UemS+Fjxht9lesbWkIZOi788zri5xQ1+WHhRiEkFuQwlCJB+omEUu7QZDqEZZn/o
J1LNf21ICNIUHEBmQz2imWgsdttwGwApysXYac4y6JJjQFsI1PXFOxPVw7TlnJwM
P9KC/YHssqYDoyVt219SyrUpV5H37ez5AiUdMVUaZwLROzsHmmTaCXfpSb0r5/Nz
TYzb2YEBA6P1AK+O3QlBhqrPkdLnn99enW7z1HUGw2pN30ghtumT+XC1TYMqe5RZ
5RHuzke/W4/zeQUwBpgdeYtS4taZ7D/pzSIKU0CG4f7fJfnOkxWY5oq6VYzhiUnj
wOjK6C7aF6XAxP8T0VDkZEtcCDWh5cFYT+i2zZXQgmcD3CkTJPnY/Qh1cNectl1S
dbiVPvq6DXs2xVlm+gb/fqdBxWQlCGQfHgPwGIV0mTmD9jLpDmr3xNfiDABZVZ6f
MJhQ7T86ejbjNVTWsstJCmTiO6C6r5DZPOFB9iaQDMvWfANoER6r5peUSFNivkdX
OvZFACqvBiQVZlTt482TSXfoxL8wM5tDyvvtHtgaPN7/Ivj7IgDYbgE1ovvvbtgq
GPtEaE6wGVgkgRX3kgGkCV4ek+25RVRuizthAx0McN5fdy8POU0uE2az4oidIdIm
OZCO+snhANvVrmM+W5mv9NVUYwQDNcIRRERYsm3RQk2ohQdbFjUds7bUZYSS1QlF
KZ7XJI/EnHTavscoGn+bh7Gc4M0R8sZSoSPImnGPxUgZFgWtS4a+lqFp/5reHLt8
brWaiG0ULnXQE6TY/Iu090atUkI+lrvf5U4Mty8Wz4w71+A3751oAoNZZVU6aeUm
RDJ3meNjvtHegtQcEVO8WWxB7ziz7M//cEie6EQA8ZT97+/XWnIbSclL0pyi5Wzu
wbRlqf7syUM+tGbwSdTmScc4sFBT88wttbzR8hPWJ7fi8ndtTUZWQvYMSKswXszA
66bHQIIyfnY1MHNZpinR/ZSNcqMRQJPg7Bsx/E8qPTI2a3T7er9bJ3o8X6TUEOv/
sk2U4bHxvevHtuinccrU5XLarBM8bbtwB6tCoMkb+EE2CoyriDYldS5iO1zW0/pX
r54dP/D+uonNi6bnx83PkOv7mSDu6DXjzlaroqLmMl4yvPIZ8YOxceLcWXWic6h7
SJZgd1u/CGnpGqAxy5l+kah71Fd+bG3ROpgcCEaMZGwEsS7YMB/ZrXVwe2/fnoI8
iW1uJwstZUHrqjIOxkAr2ch7EonZ66D9xcMOuaCKhWBnEgnumrXWrIynt54i32Df
iFqpyq1N2bmtwPeWg1NbggkiQYuhPG2eV1NjpwtfPy8FWqj/BmGH/MaNTQWxJNZV
Kx8WX+7y/0ktBgBmqiPWnrg4u3IQMBi1O9/EOb8RXqfmU+/oATdjlKBWGi1PJG4j
0LDotwQ22me0FRJ7fqBpRQhCCpetRO536JenSn4gCLgB0SEu1+U8z25fjGuCrIZL
wrrx1ldQD/Sk6SwvUdgnn61xrIUothXyD7Y1ZFemCIdRZxiSbzHExSY7zqS6QUi1
VExnkggS7Gfr7ZlMtPvyna0ab4AU4sURrjRHFLJt2aWFvN3WEdFrw+dqAOPi8neT
DXvehwwztQ5By8J9ShLzau/YExFtv6E7/yR9Y9K1IVfxcZHbo/4FNHhcykFOXLDF
Deqlpdwm8UdayeRB0mJQryZr/wbsgvkq8W0ziBscrwcaim5myFdMg9Z5uctiBwCd
Kv54s3BizKO29RhqUz6+FUzcs550Ro8B2vnhjHCmrW8pPt5GoYOckQ/MkzDU3qJA
4NZtGc4+Xy9HEGLrtKFkqCUXRfZRJKQERNyhpkpgl6cdypIUeZnYa94a9JNC8hjN
mFOWrG6H5zK234a8SBwgIPXZS+8wm25B1QurBV2CcnNygjyrQaJha/sDcSobRu5f
7iGSI8LD7Rg1/Gy022Mdhy29GTYv1MTkX7KpQX4aMsWCQtdLU1PS17eNMgn+O9Uz
iHPE5dwFDjrZwvLFd5vG/dCL0+rdy8Hgcm+0JXky4kE+xf8lSbcTDTVooapNvQWe
saF4fya3f7W2gEUMvRoo/1IBg0Dg6FNaDKXXqFTwgWIzq3febYle46o+pTPmju9N
Zsxfr1kfaDzj2m/YQ2pxbAwnvmHtAKjoxAg8Jaz5VjgTEvJ4sNcfXUol5y7QcaxL
Nzx62Vs0ra/yJe5+5Owjox2CgsH69gWdoGfSaC0n9vaPFQD9AwB/9pajTUMzzbtj
rUwM9pkk6BEss9g18y27fcj7wJxUSgFuQ2R3eupvas44gdjPsJ0tnacrla+9i2hA
aan7HBXCf1BMQGlpEf+GIe5bs9HeADWrIGrztj2cXSbVzE2GawzPzae1Xvzia8cl
W657ZtlLLdxx3SeSj0SZUnK3Galtad6Yd5zvkw3Z+5a/iSwM03HUs0J6mN3wgXKV
COCAj4BoaoC8oVBo31m2C/N3sobUIjjjGWiD5j7WQouGCd7WMSrDOA6hooMpIRi+
AwdDbEGQmsIMSCXPCmj/FFIYHpHJl+RZ2YyhAxUa14pV9+J5THPbih5TBKq0iSiI
8UNVvuZr+z7qhUBoHiO2KG/AMyfS2aoFDXylpo6/4O3sBx19zg9CjLiPsbBgJP2T
+wy+az0ebzaH/tWKSACA+TdzzV8YE8DbIawIoZWmgYNZSHXSWEOMH0nfadA1BI12
cBxVQxGSKt4fPMst4BHiYr4B7xC4ANgOmvSo6gFUp7xKpzAaltG5MUSt75tMmJ61
gvwElzacincnvqY9rGEd4bHiD9dHl0xhC6iaeVn4R+i5tVKvkohGIvtIO3OhQZpN
L7gMx2d1wUuMAVCAStwuNTGbEzL7Ap+xuGDhf7SULRVLWRqnY5kr2IMoy9B4bnte
DMfDirm4V5L9dlxMbpFmOD0NrSFcdb3PyfjzU5JuP03zalVu5SrfTG97fGeVWxVy
wEvk4vKFYQ5O+Cr+9gyXGLarfWAtKUktNU+FQcpPkTpMIcXVvzQJT5d4xKwFe3jH
BsFfmahtVPZSoxNlMkoIrjEfXqq9kj1oVhJLH9mfTD7rKKTbjdPxwqWQH21KIFeC
CBdwoEe2w5zoNHKNOdbPFHbE2hsIttaeFLYst1FJcNGNvO9PnMHKT0NiweuNjI5G
h3MF6l5Uu0VHwuULN4e6cYLpgqJoZBdkor8a/Ww61WQrTP+YVvBx1u1H0u+HVfIX
x0B4KPNl6KnKpzYH4bYKpUgB8Wpt28gw1QO3N+wuf4baYq1o9iuTDLlL6jHSTheM
ODeW4uzav4nFA/LBrOMpcb3simBqrruVehY1sRRMoRwL0Jecf+jRzzkJIP8xDbFM
+PqOwSwRpFt59UDR5sDik5+OvqdDRG8/CJgVkdgrn/BYVV0RvFOlghdoopGqqKWu
tHccFhc6V7wp8xT+m3lHsHLBHLIgr3uSt1aMjVzNIcRyr/DikEZTB4E1mhHBrq5G
9bvMneR/vpoBb2CFFdV3CSWf8I8Vp57fmg7ro7SwupJeACT+4CPVukobZC3WeEq0
9WqzqtqWqoGBcIasGFuGaHfomQJ+kOaoPs5H6KPFFohEmYkuYzqC/eSsvxXuOAl5
tNXYZVBvZBNZDDzacmghafTMmeMV0i4DTGh6Rt7SYEZpc/E4P6cu6dLYDz0Dgq98
R6C9FOKj4tRRYC5Q9XkUmEuhaj7t3reh8pwIGXFAXmaiGeOLSu3EWlr1ALjtr9hq
n02yhxwJ20pIWGSPzSPeLN5rcKrevSC8ozog91gxVj/C8QpA0aH84WFsXWDX7jUh
Ar+lsHFVxrwx9cRvroTg6K1OmOcLANYQi4d3YIASzBrOEnpN3maXU2BBEj1iWKol
7GlJdY8Ty0HwR+Hp3EW8dCPRYqtO6LIdX9L/a8IWdssy0nBbGBpTY8ntxq3Krp3i
oPuKrj7T4V09i8TBVaykNfuRs6ubdYMCa7r2UZdYQ53EgZYYiRGWzx2SZv9FHdxw
AHoDJIjPUsZBj5nKWGuVbZ3eQPY1UAgNLwgv60MM62svLqdnxwEpUQ55QtRWKyom
dbbEChd4HYq094X3EawPLi4Jtxkdq8fC9Twz5FMnd9q8vTQbGWQ2ZJHrYRtcuZAc
CiORhL4uRKyCwC4tf46OYb3dr4alvNPclTE8rTj9cJsUK0HwcM/XqxPk9TLbpHVi
NB4DeoxveVFn4zGWw5RK2G+BY/i6Sjjpc2BXYw4o/t9S5M2SXKYn/leQmPR1Ewr5
RYSyyVxSiAGlMJTO2TgF54cw07jui0/JOPmaPvsYiJvbDF0M/JL8FWyfU2X2kTgq
/aszO5tVTcwvUKSSmsE1nfc2WdaF6UCf44r10FiPLO88Sb1iT39RWaf9KyRs3XUE
+qJBgXFPqillt/QLPwubFNpalqJ4Hx3FqirsB/HuHh/WCnrzjFp+dzYvrwhRg52F
JpIMoakVAdbj0GDbGldFT+uICFHdJpLnefKbe8IquFDzAnbv2oburxevPLXZvtkY
x6wqD04QhzMiCtwFMoXPidkMgrvLJG80HFdrt2JnmU9rctN8Hm6iaUpwMuaHLAD/
yj4fjwHFG0SkDW9AEgCYnBq2ub85L72vR1xsduXDi2MBrji543lUVwlt5jaKwWEX
ULMrr1JdZJK1XkL7UFTP7t0qY1Ph0PU9xcoE8qLHRmOiNp+pHeH12E5xi2PmPZFx
vLoXzn4NosOFVvFSHkGiXllB9YYmBpcnYkGPmu3vaK/OBuoNBikpuNzAhUuikD1f
Ae+fPx7YjeIj3Grle6Rbu4CPHK+i4MZcAy7th1ta0yWne2VJfSgBNzyZ2pTWVQDF
lJbP4yr62yS17QThPcseit/oi5eByV043os/wUVI+cERolawR2YiBT5V8jo0op3N
t9SHits+Fs4hXYzg54Y19jVMca1ytAFxwJFsWbGOp+offMzwyw89ULKlZr4qF/ye
MpMHYw8cCPPL/OmHItG3qijVXvNDzvSTIrMyWhEAbxi3+sVidmFdTV3ouDGXna6b
h01eCcDuxmAAka5w/Tzy8z0IlF6fGblrFL5VZ3T/2dXspC1SP/FsWCXna3D86G5D
ET5hy2B6Vb5yoOpmlOaeIIT7EXl+hRX0Cr35b2Yg4Iry4OLQKRkLYlzmcl0aDWqN
RoHvvzhnfTKTS1RanjV7fbD8c/B4+ouMugdgdjNvCzZpepidAGzLI7pA9r0yuW9/
SSEcizRWL6Ti1xhLrlNuPepm43cSB6vkIb4izXDmQo1MyAAfmXRVS6vzdwA+5Scf
Hj8j5OLAWsBZ2d2L6P9vdsr+0Xiv+pUbRUoj+tketVJkhV3aoAc6ZNAZLsO/bcbR
jsLW48FkrCyCRUDBZ88Os8bIbfWY3nWgp8Q8OKsUSSLyiZHb0tKoutmIw2B3BvQO
qoxyl2cCTPlxK5JhiTM0LG+heQ1KeTDeVCFNOJI3O1LbLswRTzE8AGxjF6VyOmVU
Llw7r/yY5bMAYBL4ZwAlvXYrOQi9UzvFKoXG1hUxNWc7y0iWqY1k1zke06nF/FDo
JCNPZAI01FOV+eHlgrhjdQSYmOIoNyivRfb4+OZr6pfuvC87NPBltPtzWF4GZHto
kJxyyIlGPhcByECmOJnoxnIgUNf9c0Eh8RwaC+YYsd6uJ98qosc+SM4BZExCp7SV
r2URPKtrA+bzcFhq4zWO+w8jXCFbl75XrINhtTwmew98p6evly+Wyt+eGVAd3zD/
ImkvBQ170mNwLrsozn/VBbxdsPxUPfP7NQB6n3oxdXqLD+v+Ys9CLBlbzKhYQqzd
YBo00voGW9pzI9r8QTHw2O3ZQzKC2JzkbfEliwAF0BbrR3pL83W3pCwRLAuKwpsT
jMTy9xhe5HkU5dwWlg+4+9nEHEVLGcig+fs/acxI3gKpPfMmU71pCKEhrjvbWKZW
2j8LUIEMxuLa+UZiaIhd9lf0kXZeFNdXI5Urim7Y1gg/LqBv9CmKQjRHWSTuz/LZ
bdC3NlZLpw7FewJ5xIA8HJispqsoUjmTx9FWHMdXkT95qC0FXuMUxENlhZxSffwA
JKbs4qwZmXkpOcTaEZ9vWoCbJ5UgpdlsMrruuW6k3lGMgftzVg16Jp1Ns0refvjX
HphbAYP9iuQ8al98iaoD9WWuEMFF7c8tUkb+FEg9vuA39C88h5ZAu390LHz8xrcP
/AGnguIoMDX+p5dcdBQB4XB+w0fJl9L+zXbP8Q6KCZOeNf5ekrqAVFfoW1Dowq1h
SbfWAJg3eGB81i/rxJX0FMknXyyi1XlbWdvA+lSAqg8SquSJHu3yK4TXplkwlBqV
1f3mPze1pu+hOlLxgT4iw7Fi4L3TvsTtDXgKWLpM1+XXi0Rq0eMC5djkv4g4aXuk
8UHqP2tGFn2rv+MEyPB/HwPheGN14/TQmOzZ7DZW9yqoc78g+caWtEHV+5zcPyue
FfksR7ddiRMD6JKb6uViAr1wZ7JcV4xF5TQaDgdp+8GKi6he4hl7KCeacALZ926/
vWrWcvPib0+MK9JJ9KHPwgQXuWVjZfZOZEFYw+RV6Lu/RcR/7X6Z1eu5/Ef7RV6m
iehI2RQrq5KhxnQkSHGNjuZ2omyfwpB9cgDe3nc/D1GRiDaeDV+RWiIYoFSnOdIj
KQp2StfSDGbF3vkR4Hlb+goP+aEJvXZiumKLrTfUZq1MWYfCyAKZPfV5UCrj6k2j
C6OD6dMCsRFJLucdE1cbvdQAidtRiQhoCsXNJkJuGh2nFDTj76s+WFVgwg6ndEMx
wUNFx87QXVUYEZ2xf1fWfLylnkvhD768E8ovH7i/MpgdCrv71lqunBYYygsvbQwX
gzx+NY++nqdfHyi4RCjjhSIxdftUw6468owPv/dthUOvVN7dO45DU7QNjmCY1Uhg
ijMqD4qRlMMDD5au25B46uhqhaZUV1lqmYIbWHP2W/f8I3lHw6YXZZcgvWihH5ju
IFd2ZgZ6n7XHjcBKMhC24wnij8sPrnIP5q3NnE9Dj3wNwmsDlSaAZUs7V30YCe07
1g6hi2na6cUlAZlnSB0qYkVSAdT4S75VK5sUqQ3+TeyWphXae9NalGAzwLXKy+0W
BzkMrNBa/ttlhtzd00Q1VsRWDovBlIfGJYd3OIWfwAWkoi1JxQmqK9RnWG0KCrP/
+YIethafmkQATSJlB4pce5BylmR6Su/wnwOaCYQ9nGR9nhZBwyQeVn9I9k8mdqob
HmBXmZZ+zAc4n1lFfJux815OT9Ixcu9P+jsXi9XZF2on7k0pvGkhQwSv9b+mq0zT
5puJXN5qw+VrBpBFmporQcW6s8G4wE9WGX+DKnSJFty+d4tW47L/ny1iavAXqTsf
pJWv8KleA0QeQBBLGvsDDrK/kwWFllg1d2wS//u5fLPoTpzxnKCLShqJwotrUFvE
cv6s6uAGJuzaLI/V+yS6tyYNVUipjVgYuqXjXMfbTXezexKWBA1AN88UjDeMqGAT
UdB5fnT33L4m0+YL7r/O4h2xceWoAW41qz+jU7402Ry+g0/zX49JqIlvXEweyLES
rp8OG85IrnDVnH+tlDnHi87YwQ99EOuZ5N+3wV4dIJLAjK6TY5AlYYZf0pCsNMzk
JanKbjI/fCMae1RaY9WiMdc/s7u+SBzeKIOKd0C2pyiZuxsiY+/8nqA5Vv8cV6UY
wuH7voLiR9Y6cWo48/JqDYrVpv60b/or2NQwRxYVZhFWbL/1T7vjuOVhg786Nx8O
JptkmDZumR92wwnDuHkpsr1aho/0xi0XqJVkGfvZowpAETnolGzVp4UtE442Sel6
2SPx6ictpQMP8n3iFdOwqjuO7cC01jKsmBpYgemSxJ/w13VpG/6gn6TqXebuM21K
tzYa3IDlR7KqjvBb1WP7wt9FM27fVNE/xA/Xdj9iQPIymmjNadwl0QuLarj2NrmR
P9bssXPiYM1lCdNmZSEj9xOrRJGYqK8aI3P006hTz1twuw2eB1P1LUGKZxFBHM7G
/xHyejD8LO+sG/TGWGROLM6LwgpOc/M5igEntu4I3ql9B6NALuGAqoIehCFflAn+
lW79kSIqlYRupefjiO7js+dUDmAj3av0R0IvzxZA6FQkNRHvbV9yizLYFvzUoLZ2
ucZCNNw4V2F+JmK5RtT50DZu17mXQiLL7utwdNMsqJX5EpnuCVflYeN092w3C3oN
ANkj2s1mpwZtel3cNuGybcIP+duWm1E4o+2bSEnA3EhaUnXHzJSWHJGvZYjzpvNQ
5uH4ML1wVTOHPWW0MNQ7wZZS2D31/oAExVDkxKqkz9CWZZvwAPMHxbsiQR8SIAAQ
HRgpm+7Uz1Y0i5ImAjCNW9LfjWWuQXXDEs+U8UM+TJUu4I1CWhutWg/BvyRPCeHB
PNcbOhRgGa6DawACON8+avJ88iEzONsVeTDBLVTEo5vpfKyrqTHgp5EpVooadaoI
Vt8RtXTJzxMQ9c4u6tYqqn5fWFtCkE80zq9aJOgu+VDJCK2M7NuQoFW0Sd6FI/Fn
DMJDCdtt/KArpRD3LgrkPOvibTEBEvurMNLT2hzGiUpkHn8XR/4p5RoMsuhcxcgk
+L9ipgfhkeKC6FDKwEhvFoi/IbZFwoRgF3V9lZS7CBY60CbL6I4sm9X7p/YNUa1s
PFn8NFr/i4R3sCQOLDqO8ETWCDkN9QbMmDtwtauDmGHNPxCaMSmTZsLrryZDvBTL
EmRCvXYpNwIKtV2hTFRO2qe74hz5SNCxFikFkQFhgw5CKKsELftpN9SwjHWKIwmR
pJ6kHYP/xwiMl0G58qaJcS/yOetY+0DGV8P0w/P4rBlJoT6M2/Xl9EJLmy2MSdXa
8jMX35gAYpJsmodaIkF/TXUrFmDm9akA8XDv1cyYLEqd8yNTxDOK5dzAFCBoSqxa
yfxFP5C52Tgeob2krssbCcWCq8nSIXrwCY96g6fp9GiXJFSLGl/IRZjHRS/JHgtL
q+Ki5tsmQi+F6k5t1WObxVhd2AMDuMOPAiag1fzDzZG9IFqFni+2H4Dppzx3/XDN
m9Ic3rKNlVyFEbolCf7972c9Lo18JT5st8O3iY8mn403/orOV23uCbG9dJbeUHDH
zAqcl2CjnGwNy8j6me4gmZ9e4OE0uHlkeyx0/7zI9rf8A7H4pqBwjDGZyVQ4QkO8
mnSHVdGdiddni5YCgxbwHicaZ6paPnX8UlF60brwySNY1+Y/GGkBkKwfoxteoPPj
kciNTjl1YHKaozT7mlxSmtDJUywbcoECUPfSamVPPsML5NtoBHXybdRYq3uZD3Jx
sNtxnSbIRYlBB0+bqd1u1b4kut9ZqWlS5FqhTd+dMxoB994MX0hFhBojm3JYC5x3
HakNLCueC+Tjtsgkx/zQS4N3VD3h0yiXvfQTtEUfkxCTVJBtd6oganCzX1hM9Xr9
Gs/8LEvvq51pzD7CcERbrWGaKFkELW8cDzclb4j2ZLbSqAqXTifYR8ydKrwv0KSx
LPB2cugLN46lprrenZxi0HfAiXluoNj1fhysyVg5lyqdzeCf8PP5+S1rU/jajr6t
eqlj0pKICNMKwEll42hAETmPxXHLNWW4qMz/xAbW814faHUZtpmkoxFVtqMGUJKu
8T5ZL5GaeSlk0MJK8c1JOwmyT6/HlVHzV19scLDXPjMI/Yhd1lDtCwmbaW+jr2eD
87ROI8W/CUb9mu5XydsmnwCyDxQfTl8091mkZbfvNUCJQHDfhowlRwcCgkVeWunO
UzDfEZzfnqkKjLoU9Q8byEAsPltCHewM/UIkuRkgpdQKsS9RZQllc2FkOzDsmHc4
dlchwQGFecYJTnWThf+FE3SrEDAoc1+sFYNG6oZIfCMeeWpCn0M1M96RTCHznPPe
POdFTj/pDWzaLQKklk5WPYOtWbVXTWYjIhUpSR085OeDoKF7Ixzkyl7eu+y4mcG1
Fa48g8R+H+CqCPsSrA5lHRf5ArZklsKEr3ERR1Aot0rRg5MpdzN9sxHbx6bu5zpJ
XSvEs5fdV3BhQgro9ahrTHBE1iGy6ZWMhTJo8m33RnPc4HmGfHq+vXTycnkWo7J+
JUg8tVHfW8Sy3X1QtowI3jsx79NiSnZg6C7uvfXeSpppzXReDAvhA8HIVgRl9Fyg
6/H7HTCDqyEyR0xdHbqy4ipUbCkntFwdnn4uNbJ9nIYGDXQx569Sp7d0uBpIuVUH
omtqTEr5vBzYivbmlmeQmJ7qGOHNs2J6hpClkNpTS1qq+leoonyZn97AOz80MANg
5+V60dml09GcdJXEoAmZ+KzFRghNddNXiK06gi19tuMHsXrzjXl9jDg7FY+hXYnA
34YgyJgVwfS8/RPaAgHm/LcoBdcGLOGFZADv3/grj7BqiKSjhAFAKH4LlR2Xd9HQ
1dJAbMcR1PLd9235pQEiojY2/rN3o5UgaGExRoc05YBKG8dTebWZEUB+XWO0SclW
eX4OiDkXEQDNKvs9XPfriSxFQ+OwqwaE1ze4dWdFZKd42joUicuf4IFSSMU4y66Z
JmDiZdrtsJcNP+xpySkuYMUBFnYXO7MH1cYd7e5gaT5NpuagNb29o5lA0hFg0P0y
WobSDXKEoa7fd52en552o/PFiCUw+RcHotze5CqVkVsq19PAl/UkPQ8ZZCvk/h6g
NycsbCRjma2fb3w2zW/BSrggxGnC7mYZLpxylDLcvW2X/MMShWh+5H1DOtkYpXoc
5ZGJCiQMq5K9R6hm4TFh1RztWwDcPJD6VQROrBwpkczNHMBMEODrAs359HWGsTuJ
yQJYTh5M4bhL7DAEri6AU33lBG7IXrZkGhv1xiNRMiQEQqQSxuw+9SRcRMDkaKOw
xzSNmLUd4+OetoF5rzHLn+R/JO4n89pURHr3TPwe8GTMbHkv2xQ73F5m+edTUljD
rZVKGVI++wQlI6vYK3csLvfpCA8TW7ohlgiVsB5I7FTy6A+owjDF1JgBrDwm6+0f
eBp9BWM7lnCGYtBjcjkWUuuYwHBGO3sVOujARlNDNprRMijNohqEHUWozKls31Jb
wCogynhky26FO/UYhmQbWi7I5cwYLapBrFGflUuJ0drdTfhv3t/1YBFIlUsvBGgg
OR/GQmzHI/7H74tNKIy9LZQL6QurLXeFMndRK7/wUz5douBS36GKAwqbq+Iy/JCc
ypG69H5KNICo4kqql5azoBAWEF0dG8T8yRkKBZssiX8hYSG28oEX1q48cb6Jn5cT
wdQYWYnv8JVXEfnDVEv5zyaMCHW2hGrSOSDU3m/rqZgGEbLjdbPA+CBbn2R2k188
8+TkSzCVv0zy4LxhPJjWgCCbyhXsci4oWtmdcfotlm5IbsIkPumvv1H8jY0NWdla
j4fOWx54MwJZUhbLLi7PBnU8kFEVnnLaeICqvhPk/3MppfoEHGw44pkaUA4eeRBk
HduG29xc5v7+xc+Z9cW9GgnVzjwgY1VryYXgsVwBFcE5wFB0+MZasZGl9e+pptVm
R2O+yevb68Z6t0QxnFCqBSqK5W0MKL37m3syu+uaA+Br6f/bYeqykVzh6GXlXGea
QIWjKM0Y2rpGYFS0y9eR1lr0V8Eckgr63HtZo0HHhV0LXTtY/THCWbyaOenrm8o2
hm/RUI5v7IixhepDA9yJhxQz+xrNAm/i75uBhf2FRSxk6fPShs21vFkcFn1G9MX8
tm4s5mRdeHO6P9AO3FTk1wf1EcPRFepxZYi7p+4HEPfzJbOf0D5NVvzJyf5RlBTo
bwErkUEHs1lJubg3bfQ8S8+DtAT5sgNoY4Dj4HzLr1rKGOK/i/96JfyXhuBfbnCH
Pmge9+Jk2h7Cq64WwO6gmCe1bpf2HXMJzLiZIwx304GWQbY5LxWKVUGEnJ1sYnjb
3T6PiMSkp3FHZVbcm1WJSdDn3oepnynMUH0Xq2XGilE+qr1gxBS9gBMrxCFYxZdM
ShjZH2ofdZU3tofHW9aGFyhXieflqOsXyyvkc+3Kg8usf44Mcp6dcWse+7XO50zy
myXFW6vWaFwV8rSIsL0rfJVASdI7+aHSbNF61Z6inGN2WoxY1usKCWDbzIQfDaDi
EpcBPSw7xYICWKG4Si1Rh5WZMwTyEZrLvOcV95puWDCdwwn+LjYRhZC20+B3IMOH
Nur3fWBmWwHywNW4V2mJXk5HXmA1q1Erv9z1EaSg7DTU8a7zkBskL2RPPqN7K4I9
ntbNXODaDpr3nQgSSaYZjLy/LefWDjsP+2SCs7wzjb8SOuRzdtaud4YKuCXPjWlr
zfv0EG5dUwMIfaLKYWhBJxJ8RxjP+u6NifeR9fmcDQnF4UpXKSSyrjV1samlDhnM
lkqMsUeRq1necwTZ1MH6n+OrT9NqK4bCAVXuheGZrtqA8iPak96A9bbRlr0jcAuE
48QRgcsalj+hSYU+R7YQWZ9EeA2t/CB9Ky9l1B+N6cfOClHizSegS1Equ4ooV2MX
xa58xJn15jJNmsQjlaT/R+juSDh5j5wxHHCau6wgH612Nj+U+7yl1Q0Du3Wbk3fy
DMVOLvIZ5zT2Zq9CI4hBmioPxG15wcV6nCG9fTRR9Kbmw3KKwvwh8lA0Qzw+hcpS
jMIW6M95iKDOz0HHerxSzKubVN6bY9Nq6DzZ/8g7e94bGXD+77ix19pX2kELNwIs
ILWOAlsHOLXCx67/L0ss+dtOlrUaQkDRC3tmS1hwXYfBHjxcAl2KFEVDJu05xYXv
bDvS4N7KfxQ8UrP97FggziSgnIGb2nPVHKB+DR+GTM6aBI+4kMJNcVi1xNajrZ08
fSBvi/XbcbHYR+R/wf4w30TCLS1TiB84L+iNJTzgFbau/hGy2yCyWhj3pOXXZmVP
2/OR/asbK6WWCAc06sgDYNKYRELNC6UMrWwXcHw8bjMAu+yQMZ9JkhFJ3CPSXcUH
OwsIhxOTIOBS+fggrfU93dkja1ICAS7uwcDing0JHF8kT83ykRjDWsPOpSP/+4iE
We1EI2LuUk0Mtkc/o2oxvvLwgnfrbyL9xrWXPqKj+oKq3frKlvWfN4RRTkT3EnMm
b4ruQLMUcgTQkLKulNuIByDQvqkbIPQZ5B+WOUkrRNtufhw1Z92z6jOqYyKuvNEx
lqE968kkBqStTov4+2pfnTSQKqJlG4lR2uEODbc2Ym+/GscJ6vOd9rJ/T3QoDb8A
jPEqhHSFS/viAkCCHFKQFRQnwOomaAoqX+j4Xew2Xd0VkkvL5jBOq9vRLwpIK6Z1
SHMxcEqNILl3fsLlyEorY0+tPt8CZNRVMFYFpxzSSSha2YDguciF13Dp80PdeKRG
lEL+2c5pnU8ZLtCHwo5Y1yWU9XyIhp1gbIjFQ9g38cofJ/PyCPhY9TVG8bifeRl3
YVWRrHHK1a3tG0hAOGTZRf4ZCKPdvtHkIenAl5753IZsU00tfebYm4PFDiW4dbo1
yvz6yOG55W/01a5y+lg3CIYxjuUcLjd0PCe7pgxxZYqPNKC7oXUjNjL1OI8gI4yn
Kp8/E9F6AR3xwYfDz9dve2IvDV5hI86lUbNTuWxDCj779/DGn3vUNheS7iMhmFrA
Rc+uSat/MwF+twEA1exdz3N4zUsMSzOAez0sP+NiTQ3s7QZ4yETiD8XoQCKPo0Xo
Hng/fZ3aee3wm7Khb2RqWo43ogbKzZRScEmUr8xyiEZn04YEqYoXhYNTulvdpkYC
LaWBLL0/dvC2f4S5v6SE0/HpuuTwMryrAd8WKpryzXJOIV2YxkWhwXHR9nixlf88
nCmbrqOOxRShW8c9TVf+9+Fez87iYJSe3OT3YaHO36+TuUzy4WHCQrVFgJl8cxIk
4oSax6SK6Su1aYTcY3wvoclFafhVotI4/oDX3XTy6KkkPcDhcfwAon9ohqKtcPT7
aCWo9L5b9PJV41BBwFYY95nkINKYdv9QgizCgWvjQmwseC3FzhLLLA/udAtFD53h
3khL68aep9OIJDtjtY/MF2n7LAVigJXNw11azHMYwOiYgzBMM4ellXErRZBnw8BX
tou9APUOWEwIRjkjudXn5sHhhkIsufss04rcSUnNr4g6RmEuYiKW59bT44l4tIbD
b9kw+ExDKYv6ennySQ2nAw/gwDF4UpjacNuk2KoVWaPeOsEzraRtrBJrDq4f2ikL
d3EJLpr0R8+oeQQA3jBj8urQoVhzQa0jdnkKZqrYPXJ7AEbgiryL5AhNjzJn0Os4
Q9WyBzTBjPuMuiCOu/7ObsPwhJKWHPejnIa4gAssyvkzX8wqapi4iJJoNNh5muR9
X8wDhpmlaIhc913s4xKac2390yedIdJuw0nl7MlsoWkfaYc4IZNGeTAVatRSHiSp
yQn4v4LMtbhVgtBAr/AblE1d9maMkS6jkYxbjwugjEyzK0cyMtN0+JHUUN9ubIkH
YefnRAZKImQG9FqxoCoT6ZrAEeHXZqupq4BZXUZXr7+RurT7gu+aBKVXkcfE1iFd
vcxrs/+SxPiPAxAhT/JXZ+mw6VfepCy0ztUjqcH04ryK6EtuJ3LwrgHb6EBzSGvn
OSuk12G8X2AePM+etDsqGJsIW0Q7PdjQnf2wDG7FnwARCNEI5Orot9/wXvNfLT4H
HZ6/bhlaUapca4zoHNRf5nB3ikkIW2c/VtaSCECAQdvym8eUlFfgxNmGeBnf8zHe
0YCpBjzMBxckEHe6x1/dagV/dEt5gu82V5HN1zSZOpHR/+nNuTua4n8AuBkJQHIW
OEkC+VbMTJwFobPwCRW2C1xG2Zb9UHRrl338Dh8+xB/b5rT0Fz0bnhanWBBCGtXB
t6AtaMxhEZOKJL5jU+cM3Ccd5rGETubfAsaDBt30iAMB2jeTtiHl4OBfjmTToF4t
ELmYYPo4HwdIsooFCMQPn2xj407PCE8AMBbiuTKCzpyyp7uhg2D2o1ZM9RhUeKAl
hPuzw1FUV/TNq7GinxxSb+j+Je+zQXiollrjdEz07mUmbJGc2QzmvPm6dQVUOUNL
dA5VoonOaXe+xsoQc7yLOANo8qYWWNCq535wTUtRT7k65et2ZDzsVNU4FMhYYtzy
VNDVh73fHD4i0S9XV0k0wYGUNVyKgk8qEi7byeHVPCTMKJAiOjBFppawiQVf3uj6
rsrbZJNWDWHVxvfZFrJ524p3k8FN9xkwMiLN1WLbVTY8suYPOz8wQ5nZbbOSMTU8
byE2NzOh9BAGoccd/1rXMxW9PzxFlaeryhywzcnItr/rxI+L5C6OONY2l/0AxVKa
FGyrF+8MF78u+fUvGwka3i0t1qgVP00TOIVnDb/emwFngQIOBQ61gkG85PoN+EgQ
ybYRp9RxqimjW5DvYu8uZKGRcnw9m93tr+1piYEgOxAfcY7YN/IRO5zRBbIb/usy
N6NlZiGFEfZNXljnS4AMcqUk5TPHW7C7Uua5aGz9J+k3u7KOm/sCuiBl686movYT
oFJmgpVGLYKdaIqI4HK3zHCh3d3ZELhVFOYK9GQV4fVuAoAUc/Kt5IKbUB5gfdjG
WwuY+FF9M536fDgHj2AYt59QVfd1KJtEBAMzt+SwkZyl6cZ1Sqx19a3UMSPkmPIh
R4XSEanAA4dSvOdOhFRMe61OMraI6zVt+kEAbdh4dXD8i8rjZrdKkMolbwsbnWom
pIhjb+SKJLHZV9m/5rUYnSoHZWrX6lA9sNqpjsR02HkLxF/qBfNXKWIMDJd/m/CK
ZDXnW2DgS9/OnvFDh1a+MgrKDvhibNj5ZrekRueAtkw/MRdElokvBuTuIexiIUVl
evwxU81eRSvVYYNbTsCXGYL2NOfZFxy/YEY9qJ208RGVtvPM57Ox/mKDd01ByWwj
T1bHRchOZ+y2tINfa+P0lbX+z6NEkY/mdRZy00/vfwTPCVkkfk/Jcddqina5LUxz
zpz9rQCj/oggVH56N2vIjIvcCjZswugFiQlom7SpPNHJ/B96Y0URRcZpmWBaQEGb
Uj+QrM2AGgAd151B3A2x/xkLgwzgc2E8YV1fgNMiUZDFWb0WS9UpJgtdHlG8BT3U
a4HMQZ1MVdf8tsbg9kkArhxFAsI/XUE/a2GXBRWx6ukknuNEiYUlIDSw0MfQmb3H
DSW8bmuNbuN2a8euf9wGNLo7SavsGZ+1lS8KWUFkwAKxrW2kyhFH5ighH/76YPvC
BqBYMVGtVLGcAMHiWVUgzCP/Fgrvc74Pyfz9NltQkVZh7yJgShumBVvQS9QqB3My
m6/oBJjh+567G1iPHWBB1Yxbr4twymAuhPW+DYLpG6zLYfGnIF0qG1UzGa9PjiG/
WfBhpT7BttzUytuaXy8PQE01lgf0zyUC7cQiDcs+1FqJUH6bDIpo4bgtu4oacxYL
CO75PkbFihymRFRVnWI2VxBbNKjOIaCEfefq7+jWhI3x4dpVuF+uHDc6pKTiirlo
xcKSBrMK50qhBaGckrGkgrQTy242WthcVDdt/hqNQEiWAiWrUaEwTxhDYpt8Be8F
8hehITg2E3g+j9cp8e1XRjEFOqskXzIgOofoOe3YVOF755qch3wWpB5MI/uCX7Yq
MriFDHjZfGaDJGjql3BmXgme1nxnIzKGnaxu/VcOGIgI2ZoTHoVk2TcNgykj97dh
DpqkHC4o0Jn1tEWKCifCMuz+hUaZskVuyEd7UpC2zldMOCGctdQiw5jGERiz8M8X
qJaLXQH+pwIb1nMEN6GJ6gRY8andmUde4kSBrBkMxd1ncsHHPJcMG6vF5wTbL/GF
wm6Qx8z7uoJTOZQ079UVAOtBVUfqjGig05femDreBRBm7wjLJxpZEYcRpBkI9sDk
RIKwZ3GnuFoFex4LhYPIC7VDTjkmZPl8361qlXEds/L6ydnde3hoRBcf4bpdLIwN
d2kkfBcLQlZG079MoH/1RTB+x7SSOw99XOcrR67wBONsZ3nDC6evQJdSVQaKOKO8
Y9E2xsaHEPwbakZvq12a/49ofsyK9TLtsS7paGx6dMQQnQyG+Fc3lU3M1F1nkH0j
GBHOELHytDk4/Vj+t5g/UO0vbuuJxObqEsSbYoUA35bSAw0VL+bXDdbDZKsclyz8
eAlpBVrx/CVml3M4M15Km4jsJpBB+mwDBLw5Vfp8/cIqE90y+87OdkTrJs0rd2Fl
u7FI6HeSFXR02+CRdK2JSwbQ4sRGx1sf2NkQK5zegu/NyyJeK5BS6/SjPTzdOXeq
JB8nzf8s1zNamEYtBQ0qFtGOrCb3yj1DUe+ltBsxR8hEZR13vyNvw6vajzTbDqv8
/hHuecNAwVdl2MUl8UCSyiAg8XYbLUNYpvaqb9Uj9iQ6l1ZVplmao7bfnWYbIrgk
KSXOLHvjxy8lMAx76KzQ5rOL0CA2C2TEJn8T5FW0nXMJJ0kZL2FhzgBPm96AZjY+
6Bs46KVKPdCSyJI3XAWxCTEbjqYcggO7NDARWATFDIRut5XCsqwgzWXJPreXtESl
PJNib//PZeuzDPuANl2qsVNef5LKcOZFNVyGA0DEjEGiAky48xiXL+PTVvirL81u
SSFS6pvK1845VGIpbFh0lOjto0N5OJH0e3piNYx2sn9dNn+FJipjgSArikHTm9j7
xqED2inGrpAGXgC/1Q2GDB/wBtAgN8EItIqd/gy3y5liau7ADNVcOzgMd6dd9uzl
aUskcCR6IRsJZGzxjFt/Cl40HZzKE2wlzIPknbijS3DRExzc4fVzSf+DsRsuf/a9
VrfrgZ05Qk/56X5UxxYtaV/A5U8moj74z1mVymB23Wc6prKV2+Q4o3rxYfj75Aad
OLUAJx1VgvY7NI7fSssGwfwWxTxWTcMCKpVwJULQSln72LywNjiyYL0jnsGTnwVk
09m3+3h9GVNEsxTL0H2wnKRCWLuQddlB9u8inXfD1lcw/GtBzHDWkw4QPw9y2lx3
EZTAMjU2RN2pwJkEz6FXYfez/u9E1mDlE8Sc/Gl3Vn/2W0Cxd/tFdbjadXVxVByj
j+JIUuoycQAHJ7gHj5PmMygzmB31Tf0zgLywRBjaLXBt23sj6KTrTx1EoQOhVdql
Zw7i0kDE5Ecpg+zWqUs/TBlp0CF6kQFGoLBztSrB399rHM0MvsCAtv4FfkjxjyGi
ecEu2U+EHVeNvTXyrvNN+vgnqjr4UR4k6XbEj9esZUo55gXhKMzrXKawSQKpOESK
xje1Lrdlp3yUVt3J5WPyITCg7hHNhQZCe2jiMv+rSQuIIugJMw4F+vI3g2kvWsuM
yJZE53jk9+/cMr8W4c9KkYoKldFgO4Q1OaelGNHLT5XQvEkSHcTjbb5meVZES2bM
X9+Rt9g6Z9QxwCdkvjJiP/k1XYMgh4qrgIWj2d5iOIYs6RZ9HBvPcQq8bakb87Vp
F8jXw27XJnKv4lPTQaZ6IK2PF6LMWn5Kkc2i3lFtSpaSHfJKcQKW/yXwrNHs0nfO
LGopgrevRbaRZ8S9v+JwxxRmmh2DJprAljs75CsxQFR7o4oKCH/ytw0AP06G4HsK
Ov2rJewkB7uizFMEoPvtHZQ/F6QuXtFe+lzwzc6OUKM2FDnxKlhopFwNtRdT77Sx
0jlXSsdRJFXCqD2S2DxO95lIAfkuHCKph88PGRus7z2G9razFpSrZ4QW6rHbMLR7
OLmXyXX0vr8GVNFheaV3Ypd6p8S2713TC8QvNdGE0Y5umQ2iuXIiB8qlq8RgMc3q
G54CjGDBKKqlXgBSgj2Kg4CEueSfsaC9M4JZXq0guROya/04ic8wgpWJdT9UK3uh
J0MDyWcUh/SLDZZEdWZGEPxlwniQalBXzjnp8txp82wfw3C6JBegBpjvYDfz9VLi
vfhwqOvOk0DBT+HDS/herQ5Rwut8SmC40dV2Z152xKV2JzKZj1TBoV0l4LIMMDAK
hewDXOE9RAwewdzAIKDbLwGduOgm4Bn3GG62QEHLpPa+vcO3PhrokEs9RP90RsAp
9QiWzMbD+35So1I/USWhP+ERkvi6gnucDQ5XmNyZBcldElVAxBSmsNG7Vx/5Ff11
yLMgnD4h89W0WpZOipdh0isX5JSPcU413CVAGbeHQEA94k3xTE9LCOTYA8xnbSb8
ldWTbPnqlmHF3qk8IVY0a1jOda1znJba+86SHBi3osiTkt8ibK2rCs1B1tCZP/aV
dBzmNlobv4i8hKa1m16rR0QvmSDwxImYVNvZQ9OU+uRrUfGvN1zGNIDBko5DoScy
fPT+59G+va5xDUQqcIqXbbuU7ERNeHYA4EUZqZOjbYd2P79GDNH6CiJZa4lIMXf+
kXTwPvnTD+V6dSCuYUQxczNWkEj4E2ZxvMhOfDyUWpXODOfn3EbBdDX/Elz3JiV4
xozDTOtMpSB29SRFnJK5gx0gYmFj7JVG3+72gqOZG4ZOs+m61Pc8SZLLcdwcfseO
9zA/FxLJYXgcinly0kkW4fz4BgL3LpVx9bJJT6zXPUlIC5GWKEta4jKW4hpPSU1e
v0JhmzGeOJl9t839ciaA/z4Ijp7bbG4VK0ET9LtTKCIWn70GMEB3s+yA7U/H3Fys
vtzabFbSE68Am6IRAMWGDFmF0b17S3Yq+MrVy7fsxNmgZRuTFPodLVOSyxCY556O
yL8aZyHIv58b8zJPtjjnOJymbaynHOb//9zFi8HX77ruj9AdBH1RZ+KX7UxiXOf4
DZcKVt54saTiuri0EYxSDRFqWf3fKNDjoEzTjPMlkwuhA3bK5226ksbeOblWDHbd
6zQ2trIwZ2WIE18k7wyQjWQVHobWSoHkQOltVTv1L7y3ClJ6jfsvpvtjZA66GKDe
SRPdqlP5Hd9SD1Id36nJ0iVrTkCbvJLNqIeTtKWKxkk4yMLQOJDFHFRIAG+9UiCN
iXxHUDUtbsaZOohZ7XMUTfQ8BqNHcDl1qfRxghG/xM6Y0uYbv/shJGL8uSncMmJG
WhEbOzBCrZb/Edofr1t2gsMeOo1xypqwuIkxgAuieVMGbK7DafButlQJJ+aTxiq1
jup/85j0J7StRxPzkW74HOInb7cPYGbIikkFoz4Ckxj/xXdku86UULxB+JAfke3c
7S126lJBg0CMYtdj3GtGkna1AuFZ9wy1J9UIJp1nuJHzBaHJMRKtiOca+POXktIT
94FIX5q1wjPGHpBtGlQfe/LYx/50C/RYyOnwPfpj3h7sj1HxkfrkPtmi/dHJ7/9S
C9Ps3/K866ZNqNIO1d56pA3QsmFZENtgUGXSYvj8Y/NAci6ZLAsxmeoz30rWZEax
xh9UUnWozk+jeZcsk54ZIBq+zq9cm2Qi6gA0tEMgbsJWcDYCSWsUQoqgmoy1aFer
RgoZXgN8/mcfi8PZmD5gZ9dRXOGPjTVG92nlxqa+OiDV2JQ/oGlSPZ8Lgj7EuVwa
1sCNqvf4BROWjUHpdU5N+YCnhJJEYaP6HeiOJTdqJGwY/Bs7qVQsuN38Oif3q6gm
PXNY/XNTf05xoDDSOWWe+DE6a/3o+G+nKK0GflCUPyXRJW7XTUob34pv0kZXckbT
0eFsVnkcQjDHqxja9y80KtOfevBpm9WQY5LMf+dqXxzqDRVYvQi20rMtA7SRjvFO
hZxKUH8m3Kz5FfXxkOGq2LjEvTUzjOQnpum+E28Y6ehGTf3TlIySM4A7XO698tWM
tsK3opEHQGKbvCH1xD2g9Gd8dryDBmnkhTdu7f70dV/dLDg8RONIqPfp4FYKvBR6
nmc3Ma4WkglRtlI3Sa79+h5/V+LeaHCdiDT3NlE5DXFy+tmycpUIaYo6ntzpflLW
BeFY4qlyrZUte50rXC2YLKSxxpWWwbP1syxJAzu+0OBxLck3UxB9syFoM0z4yOx9
yD8A3Pt6fElCAk/JAC1kMoDwQmVAIIF0cQzc9RWtgTIVF49XzBfebpEdPwZRVUUd
pm1vLU3i5teiFBdkhpbXbdZqNMe4Yn5TAuonF8il3QYi7O9Bi+ruJAVrZvThVxTg
WuqzHBAsLxbkWTr1bqpYRT4wj5Bs2z3mgrpSZDiH9To2ebJkQQRKaM7KBe0KdRxa
P/FpkrmG1CSTodlW0/XMO+wslRVHl38CAu+zHS67nVg6d/mM0UdF/Og4fuR3RcfX
eQTKM94r/TsdfOJTF83JfrlaWP2wudtSfvbWCs+kX88H2uaxsj1NGk0n76kIn9EG
jMXVHoWSlIoWTLvb4x/L9Z7ic1ZIUOsORN6yCVRlAF6MecYCdXCHb5A9dOCu4m5T
qJ1HmXEqP0VxPg42sMCnaRNU8WSqdjGcRC5W+5Q2w5Tz3yoCpTSI8EUgsVJCm811
WqtqiE6rasFJntaQhGpnFq13r8C9UqG/54n5jDUxA4CLdmSPJjdj+NUPfuZSnFj4
4oH/KWUkns+QDzFVe3VbHuRh3N2+d0Dbb5OLoYTs88XWANqI4TNPGG7ORmgUStef
ByOZWeBby+SDWtguwbeKxBiS2hdIujrFJuiN1/CvcoYvrHiuXNGu8kzhVqTPwy9Z
dT2VgJ1Q4eupNgaOkNdE4MxHL4e59twcyfsBDM8AyhV5yUVBlJwyDtpxaBZ2nvrw
zhm+yTynKuoKBI+DKx4jEikbeuue7Ur/T69EMr383zwSA2dacemydAel5puPE4xa
0NTbJWCPBECPs9KzMtXD7ZnIenOouMdh5coqiKGw7fT9tpA73yVCQza1vHQMZvOG
EgnrrYVGm04/NY6+TFp3akj8NW2L9yIzdqyfgCIevsg2YLAR+Htbzdlmndw0eciZ
rwAZeqs5UWuzs6qmT+v/aArN8YHb8z1e7fhUQjBNamaNsh8d2ElFmuo3eZQPZSJo
6CuaZ0q6CBu9teXYNTgAWQIpDh1s0FZfnbhJzcT2ppy4ASQ6vjj9QvRG9+8VnOxN
+tgJ4l8jm3zXZneRlymOdoVcdQBz6cfKVF4y4MmQXXTE8ShKLHVQEk96Q9sllLFo
7tZVH9tbu7S1o91hCdqIAPECbLTAu6du64CvopH7pWQZpdSIO9tCHd+KGYeRvGGr
TTzpYIOXmES1tDb2qNpOeeWyKUvHRduXzjWqS8YWe5K2okZXo3OG9Mo6yR1NTnoY
JzhgSL00/I2nVDKCerXnVLDN6oF2FY2YKQkVqEt/3Axcm4girTIlPf4Ao3k/jjc9
5ceSb4YXgLTeWI6YOzQSdPog66H/pmq/CNn6KoGgcDV2OU3OFF6dhrtdWzcMD2qq
yGR6q+/ANHl2nNqVfBtia0JCtmI2tT9VK4C79UV+OTU3ayYahbRYBqYtkIRy+feq
6WqiY/gNEFyzNJ5DqWk90ATHGeIn8+TB4aUuHcwmhsN1tRLWsfj9oV1RzX46TNQO
+D41aBGNV++ugp7XbH0cX5912nIYCtseHZnDio0so3V3jP++DQhQv/dEAb5chxLK
juP/SNUkewUNcaZrhT0K24AaoKMT4Ane6Q2NzaPt92cFzsWjh1NMtOMw3QobVLEo
OJLNlxl7SRSyAKtTSfoUGWB1PjpfUmnLSdTivZCnbeylA7arqXxFwil6tKReMzPm
xMT4lj7W3xW/a9a4Qb+lYISjzJhXMJvV36qQA1yASiLDWu3ZqE74q7Ni9AjMhPsQ
RstcXXadQJK/cWLTudbYNjWJeC2YBcmSVtKcciP+nC2pBlkj+zCJ9IFAuzMCHCrK
QME2bKl1W2blyBwyd/RUroYRuwWPo/uQai4+uARsVusW5j87YIwSlLx2ZgeXLc3y
LrMYuvRdpYc/7i3XPn2qxHMnlLl6v1RW2SRNVzIpLqVxgjUQuBGB9kAy1KK2CjJd
H6ZbHDhW48C1cqPsRah3oqRujqX7XjtvmbeYC4fhgSQ85NYPuBQNpmwPzU2CGc38
RfTHB/bJLdabTuuOWY0OtzQklvf5dKV5EKlP4xNheNFkoFO0iHfi0u5CF+9gfpoZ
qInZfOBLkPFqBhpSh+gYXIUOPz+UbAlrgaVR8epGMACHEpwiXXRyl5G/o/os4NWP
nYz7p5NbCSxKr1xeDtJ/4yhEeh51ppXn/egxguslI4u+akzDhjfEZOEwrnGZ38Nv
u+DzQUnDCbcbmZq9Cko06CPzyP3k5r8Az24GxJ/CyO902mluuHorsdjdr8SmYupi
1L+XUGoXIfY2gL1eozGW1bJ0oXmQfNbNY8VA35S6r3KK74KtE4Hylxxp9LlguCRA
FRl8VFxg9f9hckP/5e2343WrZG6IsD9Gf/pQJx4zoQXDK1S9Mju3C/rJER1KxKF5
vg35+hCL1BCkG/MHyOLnhRA2nn54uSM3mPW++SpXEARe0SUXBji4GhWCanuq5WsQ
T0Zz4YNaMEm/N5QOKD/5Vb8lke53Y3GmkhAdu/+CEvf4AbT3w1DAjOvnmnVI0P53
rj2nQafuGHXj4k5kBc+gyspqOmQEDG+v8BHR20wkUp7elt4srmEpmWXXD8DwkD2Q
TWFKlX9+uygMO4eoppeRqwP/lKFrDejxG4lZZHDGDd0CjLI8vApsV1GZiHZ/jFxg
Wsrh+q4hy6GkKRP8Kap6EU1OJ2UyBwsL/YPHpO870ZwuGuLxxSBGsntL7D0USo1L
TBfTrvyMKgaaC7SXmVAkNm3Az2UHHOroVG44lVDwrQIk0/Yk7SSUu3vubpJlLDxV
mhHjN9gSG05MDBSht/++4YGzXq3Sd9J1lKOa6CDftjk8Szlz2ULr13BObvc5KlqC
OPg5cCV3GoIPW/HNvG3qDg94azYsEanVdqJ+Gz9IdW6Em+0medVTnlmLrJtyjUBx
h4mu2UH1ZFVZeHwxAHRA08ZcKy8UmsAJfYwSx7EFZGZD22fofG6Daks3/L0DbZbM
/8HBDgGxJ9pOOPvtO2ayNePIg/BcqKslZb65p+15pSHPLyfCsj54KPak/wEpsgfy
EkA1KjbGNb9fRWYldDso13ynPqFnaQquA3z0DmWH38uEpeX7U6bm3wPcslacwy45
M4sk9wIJyzCvcqUrZcLNIybbQt5Oo2B2VqCEAIwOEoDlVAUHIP0lPAppGRvbgl/+
yznsUTcikXRHIdfMBeBA2lQ6BqXCYnNndOhxLI/fEnnNXkBW1RXP3L4j0xUPzgQk
N/R92giGUfFpb/jhoueeeVSLCp/Z5ygRtpA/h0diI5Qs9yxCZSVysLzff/k3LPed
ZDIJQ1CvyGdbm9u1sc4puSFPbGVADrQmoeaBdKQ/GSYPnIQRpXMIYZbklcXTocM1
crwSwOCq7E7qZryKqDveq+nGzaS1sKCY8OIF2uebcfNi/WF6xbozD58ml0OCgG1K
08wkChhHKeUlFxbyDp6oAfcf7c53uPOpFUemhNSJm07z8suP6jdA+5Ztu7+6gaL/
jzvdJIof1x93XkT7DtOQ7T/uHkkl0AUsgRio2uw/vk88imuWipl4l7iVES8MzFa2
/WukZRvZ9MnTegpRr5lGFNCzdCMlhGRPLApn9iaX1spLwoGjne3tPWG4A6PmxnqS
A3GBP0p+mtomlhb8sumR6ywIYE1svwRrbTMDx1Y4fmVoZX1WcZgJ1ZkHi5ZwYWcq
Pffg/N1sC3+NIlo6NL9jCnBVEdndc0eJPgGsyc8AEDY3fy8xjNdzsqoCQupBPTS4
M2XmfpCNtmdnTh5d1Duw4irJEPE8sD8gUpfoCD2r2x1RZswLaTxnDg94Vc9aiPvc
mAbDaP12LgIobj58q/FuJH96TLRD81Kz/HpvNFRFNeExwUXbf9pihe34ehN64F52
aG516PnaeORQwzR6Fm6/wOI7p61Ak9PdHBcAo48O7TwS6F1q6n33ZyhQKMkZEUzn
Wa58clUuTNcr6cLkl0u1QpR1/ZZpO0SQYj9khzzcmFP8/hfgn6vxmmAV+gtCh+GU
6gO8UOvJ3u7Nh8aYwRO4zY/5abXulyAAvMu6N8GfGj5l2BYoQHB92/b0DXezqSlf
++PG/KoJv7sa6CaYyzTPk1NM1NPC7y+PJw/+K+TnL1QfdtnwqLgAc4IcyJShZkP4
03qwB1xYHo+Dy5fP+1J2wfTv7x8e/z9kj+Cz6vqPleNwI7LFcCpPiDJCyJA+hEoA
jrk+ZHWFfB4Wi9jL4O5sAwVKfq3uN3K6w2EdBkt5nnJwG/lVS6WJTqMo4bCJTc8u
HSACioKEfsne3v/f6ayIOInXUg0VDAeB5H9wZr2ch6bAUAqwJ5R4bITJfdNe9sXd
0FmnTB8TzpXZE5a2pyNadnFVYuRzGjmC+wGcpXfv4KkCqqSXyWn3oldt3ZYPdf9W
Ph3LDO3Z9tH94vmcXU2DbcRfYEUFm59Z9Fl+6kTlZiqNfUYV8Mg9DoqpkU85rnPH
5jVRzi3dcXiJaatVyBV1Fh1PMuyaD1+rSmyS9DeaqFQGXKq7xEiA/6gQnAqSrb0a
MOE5iV0NMCCkSGPajA0QbYs+h2gY8NWw+rCWATMo+JthYz6jqwMjhGmv1jUokKj8
JKUYAwue0ag4rx2QDh2b1/XeOmp/n+0EXZUrynuhB33c+Dq0Y+SPcRPNkhUBNbgZ
Ppc9HJeJgu3aL5pf2T9TTbmFvyZ/WpEv5t33YJJ+4qR08GJMLNsGD2oTe9P7dvVC
P9Ce20f/FHlegX6cu0QM5tRmz0dXsuLv4ey00tuzNANgzaOX9tR4sDPkpqJJRjlW
KO43n9LjwItgrpYyG6yKXCpArpng7R9BEzTgGlP3T+an3gi7yWO6Q99/RqJI1mU/
eY2u53gxSIE0BOEoxFUPBrtAk/r3y1hUTyahEjdG/V8whtDmt/RBS1VZd3favSZp
zFbBAVtCxiL9Y5W5us/LJ588y5qypdOEnMK4nNN0L3v2ZIzdeWACyEwMKbepJW6j
MsT4rofTF95ZyUiuEhK5MDnWfmOzSMKtbmLxFPT47KAV/L4lsnEJ4E2bw25M17T0
+Gn2Z7R2arE0PxW0gBURz5W26A+qu4nnPYcbwEfui4YTXhtI7up3vatuhkF622aB
6j07kc15KcmzqxHf37wBgAqE/0eLatAfyJYZEqmIsfMSJjvUrf5ZePp6C5akBKXP
vaEXHMJioeeEdsI6PkmoLC++Xi8v4rF6R3AQ78AjgaCrZL3oyyPqS/sm3Ec9SfgJ
RpE6jxm9u6qpLxiLWSk1TNeADBeUDELarrZjDCISucXAquMmtNIfslf0AvZyBKa7
gfJLbRdsClO+al/aCIUyHQy0M0JmDV3/ynpJXGU2LoGFwMOfijGC7SGVvtpQxB09
hRPlMdffvgrzNfoUpmgskZFeR1F1YhXX22hFeFpl7GpRG6c7cASEyjzqQB0fS5ar
GHwCUeYZpWW9yf+D2pvx9vdCD7CWo0pGeHomilVxpZ+8HqJGIc3eTB6TBIcoOd/p
Pv/5xM7Xmj2Zztm8/YGzHZbHtm0J31MHokLUeGMO63QepiAq4liVoM1/Jz0znrb3
oCccYouclO5P3NbAkyRTl5wrLbHdLw/PcoBajYnmXe567VmOrKW1IKZ5UzR3bwxu
kcR+ASnLr2iogFF3BeNpw38p9jpFwnZhoxKzjQXJ3OMylig3XyXRF5KUde1F6aVP
UNbELrzskqPQ+n2Xcx8jxnpe3BDe1StjQUmgn/cc0hqCL/d4AkmWcRz9xyi8ajzq
6WmhFvV73sLEC2EZWmBuaCvgsdGW/b+8xaXXRGTPJuSvZEEhA/wg3SIBpFF5/YGm
AKhQtyDXG6WsMVNPXBe27tZp85R4ZlkntcVU3u/0L825MTxSTKnhfgMnxr+rgKgu
kFZ4nvnlwLhcUEzfRtN6DIGcGBmEiAFqEE/OJg0j4obn0We6RDtlGSj1HMN3AJJH
bKg5WtTdunTQudd4dp0LTKKDyK1BLcUbp+jKE6Jcx645EXM1AF8zuDDUh/JQ9NGe
BIpFl/xqZ2ejAYNlou9xW8HIQRNwg8JKxtXsr9HOmzGIrbrB/L94OQP8Bv62nGzn
j4Nwb2kdwUKzgXJ8MV/hmXTYHmm8VBsHxF5gTCPw+IUvUn+tFMsb32KhEaVcIUeU
dJHVkpBEMDEFtczoMYy8VCuAZ0EgWlTVfZOtuRQmhK/fNShXs6ViafNcAAKCJ3Gq
VPIQPRAM9je9QiKv5l0r4IUvb9yudq/xt6G83glQxlfPjYGXkXunKwy1CNXzksFd
dPdJ5KEUPvnBahWKiepnubCzSNgkPK70fSmvDtfoygZ2O1oaUs7NksgA+9tByE20
J9LujFmKO8qWfzwu7IrqTaYDOl1ECKN0LjF1qb7MsJUHiWTjA5JJ9SEO+CJVZwYT
+63pjYnD2o7EgfJU03Y9TlRooqZa6bvTLFmiHSA56N6I2BklNgpAueY9V5pzobv7
wsTiEhaR0wfnEdBFRwieQ+5znWi0hFkZvAHPcQFLSXhYjliLNvdzmkw5ZPF2lbP5
vM83RmvUKm5gX3k4qyDjSEV+2/AOdhcXUvVPOLTk5baZUDEmeoBdSUkVKgogT0mq
yucTTCxPGredrQyGR3j+EOoQmgwT66ASJ/uuRkU6UJAeOcphfIE3l37azG3Dojj5
ZBE7UMEcTJgryg8DG4++bnw5dRg8TYV9mA7KQSVL1GT4QWHqlBayl+BM0EfyerXO
BMroLDUzsGKlgRv//qyaBJRQnTWqY4IpYV4ge5MNpEXkVlxiEVZUi0+okqCIlm+m
qyEaedUVSOk6OosKkEDgb234gV1U/71ey+Nw+q/xT9EvkaJC7d8BPuRShieDjlPx
uSvKIQrgxzXucxTyl3Nv/aNDSUsKatflZ7IebUELCCywC+Y6IpLaJ85/kY77r+zN
wCuBUX7/74nGlObW6DVe3qjct6sytMW1wWxEsMiphv48olELaLwtIFpKIcw9CFk6
N2Q/eqpGRBw+mclgOhrnfmAeu35d3hYR6oaSeTgHiKOwScPHwKGBoBXNoCLeHM9K
ZcS9yR1dIyLZm3BuEdaG0ExNPRV8IQQ/i6Wrad4XQD8Ps+sHU7v5hxq6TusDSEgh
hrz36H9Qm5O7+xUUmZYWjiO459QeDPupNMncZiSWZagznvs9eUD2DrVVovCtlXHz
y6fAQZdSbEkVtPnH3VMHyzkBkhdtMKeZ2jBfDKNHlpyolqii/U7T5PX250lLqhQe
o1HkVeW/1sMIXL7TcW4sRd7Bi9V9CqPinaqUagu/+wItX7/A2l6byZ3nAOguMU0Z
JzX+dQmyymsxi+PyH1yWXTVvo5v549PJOnaJu5tbZs1P92iyW4QkfFbwbZDLtReJ
4FR20g2PAHG0VRgYldN9dR3dB7KSyHGIQCoqjb1knJil/TFHMhS38FFyKqSoebpN
KR/ycSSq8eN08PyB7UVqGJsed732iqQQG8Ze6GACPptTZGqPRv2KfM/6c6LOhgRJ
U0lktaTu0c2O+OqlQZ2b0o6uJwW9naHBNcCBYQ7r3OSfbsaiCLVdXeVceVOYklNc
aqZg8Ygs92uT16Wo2eVUu9pn3mlm5nLdFOOkto4w8aqtf5FCuM81Q8jHWysA1hco
YRi0JepR5tPL8gH8yZHtNa/ecKUlmDyGTLvhOrhoGI06eZfDhn5VBaJtzq+2i/Bf
V7XzHiG1tJ0yvGi9XFMFCu9me1NYuYHMnDynM7z8KIYq99sxxLamd245M8I8sUHo
EJ85JH27xKqfS6l0VnwmFOYnKkkyi/b9SPp42Za0vtMTisPrT3bB2xukEnVC14N5
cN/7OsHUxuedDpYf5CKFDG+P0ln4frWON5FzoCl+rCRO/P4fGEO2MpxZCBvsibbx
o3msE6CdzPIB3sCHgPG2x+NwVQ75U+bkV6uGFuG3xdSj9sUB8hAQWT8b7R9t4VV+
0/xJiOPgv69pdjiNgJvnpcE5/YiTXPuyjx+4MsGZCPQDOderPFiI+w9OEsjJkTPF
VEqgnj58yA06RkANHuNyIkz2qerXlnTIKK7u3hDGCLz+1YQ8MyfHY+2Z3nAeCpEO
X9NRnNOB6lTX2Hf1MyqsbBcJnie83nSByzND+oXfFXE47xq0ise+BNUUZ8y7RyEE
jNL2jqbv8gxcmGlxQ1/SPhRuj0PTcT5TQcJs8XJkNkllSa58oea/69+KY9vZEDXA
gC4TS3j9TX698dTyC/jhwYUT3AwGvMf9kAriIEQn6DiRHeABsBV66d7jSO80rwlQ
fbyoHFbG5HfTG2dDg3OMym89+w2369yqxDly7agClvWXA1R9qy/d3IrQgaguQynr
027v/4uJwr7GHqoylTT4X/xRlAjB7qU1cJ9GN2QyyfnJG5aMdeE2MEDxEIH9QvJS
N7W2hfzcRfpMpg7VW/4SfhPid6KSiuaQYqy/xTb06SGShq49KjkQEopAf38YpOtq
inh0QwIzfqLP1NmovApPOM1wDhCrFTI+ddIFBoWBGmE6uSvUoWBDocpzAg+AG6Mm
TA5hGb0C17F+79gNpFofAnpoeDYJ8lPkLoA6UtigjPOgWrN4dZt8t2g/MWYc2xgi
IrseNVeCBQP2xJzlUmvMJF2v2fRhWuuD3+BlBo62QI8w1O+kBDa9m/j4pLxqqwD0
wrckwZ3F0g+Q9rTOZNFOLXrTftS5V3ZHNDlAxkr6pkv3aP9agJTJU9I5oc4k+WOp
uYQRwTODg/LI4ZeSbGIpQLxISh2OzpxDqkqnsJQ+T/dTdCd/z28BB6hLfVUShvat
e6qUSREAuonspLLvX0WuyLQ+V8ktophcJZOn8RUiW+4VWo2eWUv3t6P+pUP4zt0J
C38b3Sj1xrnRAwQYS/iztNllGBNPzQlLvE7Tu0OKxZkTWEY3gaJcIhNPlpopBfxb
YfwGcb2u6jnw61jieKxbQLVZzbr51Cqe5MnIatgF62ixGlbOoV89YcjR6uTnb458
NaaEDodPCfDTGhMfWD9AiDQqx/iYNzqT4tcRd8kAmLmFbMw9CXeR+MzmAvs92uEb
QWHqY3aqd7QIb8haB8pd9NYMx+5gyvEEIXCOd/6wBJuOf0+4XuxjqHVCateM9ibw
/2GU9EUd3DHFj7f/LuBxxg7KrOuyVJqhdHe/67WoQ5MdOHG1emF1W6K59lC/gvM6
s1huZcx5oiLSiB0amvzl9dyYpycly/rVaXsjaQ7Z2ER2j/zHtYYcBPYhj59m2FMM
7mL8VFSIT5Rb7CkP5vSyNxz5mUk0KIdYn8DXSa4R97TKSqjswrq0GrgVZf9afZ0k
6C+t7La9HaWuO2HjHD+8c/2ZaE9wgvAWygvPmVcJIdR1IXQj7jDsZn2l6x1JhtMv
6hbygell05IDZn2dkXvLvLiUoq1nf+mK5JRVGuRRzA6Rz+OPWzn0q+lPsY96gyib
06Fxob8rlthW9Wc7JjBVYoFNbITpXbvhPjhSRm1FRsal17zTiniZ0BhFCqIqsMS7
R1XP9qvBl6BxjuAatKXk0mGID4gQF0CPjJvGoS2NZNAzzS9LEADo2FZR0Krw3x5n
JwWJCYt2hrIUBtNfbrzUKbK2HY7gaGxydwfgzhPrXW6qYrjxoO3GxcDPQs7mDIbg
NEByyBwVaCp5foEuXO3Gcl7s7HgrVI88SAwtIxbjrTJyO19O7kj78ZBGRrk2eR3u
h+ibXxF6jrDkQh0JjPNYzJUnBpK333yOy2bDQCRyiMfbh7tTWTTL+mUclvpGM0oN
6GHRi98G7rCd5K7YcCJgmHKDlMqEuI+gzv+C157KGTK8/2RVzCOrUc7QaA8g7/GX
y11/PCevwm/PkhzRgWAVi1zTgc2wcFpNAG1OXNw2CfPJttWPSfQRGc9ZsYg/WMvV
+i6C/HGOoowoOvRGFatDeYIEtepdEFGL+q/ZILSq5bUif5p4wmIEkTdX0CtC5nWf
3H8VSqdfQCMiewF3ojNg9YnBbDPVqLhFOlhshQNzGJXCilxL8zI9WcYYjbcDRmK5
E3EJlA/oS9xrIZd/XT1gXktJBO2btavaVcwp9nkBrWwOG5RLkc6C1GB1oVoiAn3U
0+xTWFQU0faLJDLSNMOrflMD67axy47IASDkI1mm3qsayeu45yy8nN3NkUmCJ31D
tlLzIvMHy8YY8FuO1rTSFtx9QJHCuk2cy9nf+nG2vi1InQJeHBEyuGQrNDmNhy6E
eV4RBJmcEiy68+dPQ4X2DcpBDfe8VF1YxVIhMAEJzH7ic6azpsfBKoG33tSAIsDW
I8k3x52mTqBa2esQwoCVaMaqmxyKFUuhpOtOfEv9e1hBGybWu0Jh2buhWDnJUWXU
B/5w6Y5ibeND3vNh7LgUMB/0yc/9bP+4tWkSzUD1yOidU8iIAZJOJaXBgeg1h0Nu
utosNpusQ4N6eysxJ/ez/+yKnfZvyobWM58Mp7+WXDE/KK9egyg/VxTSbQ/fFXo5
9PTgSiPMFbh+xC+O9LKOGYjGWz57CE7+5tSGEARHGp94fH/hXLFmjBKAu1w5hAhT
qlZ1sNUIri6Ios4ECOSSlsCOKai3puWgXEVmoYA3Le5Z26u+xQUoNbjhEzQ9AD2j
5fqG36hebrS1Zj6//VcBcLt+9ha3d94OsCNmjeAZ2MdSiDlPTN3ytE+P3LyNDu9W
irbezQlQsP//qmCgmgpwmdaSftmBGx3kTg2lHkRu+X76NTTLNhEZBEqJb6I2qvMu
k7g7/3Bdn5evTCpKEnyMu2V1TeCEVOk8wpuT1NYFhfrSFJRU9pETs+qq8gzKSIyX
SayWJLaGlDgM05qPljUgtV4aGZmHYReH5uRZTqb12Yhlm8mUSW9ClcjRYjXj8wq3
94s5JFzp2nFKj5y1J84WVbIqf+pchjPnjC0HeW9qYA36jbC6JUDa6haz/RfzOw2/
zLmczioK/7AuYNaMAFjQ8lfFRaizS8vVjw4MxpWIsf2GfuZtppyEfnQiIoaDsY6e
+vFcIZiunUwBb1dDzPYGvd8UM61oOYCQnIVcCmc2m7alcWKYph8k0SOJiTxxIe/l
rpQ2CjtADQSTFsS32OoTEGaCRN3d6UczZvQ+sEvCdVAoa/JYpN0v3JKpa23lMRLE
YMsgQWANPUo0MqEuuwJi4+Wb5qIumn0yp3DkOCG1h4m8uRkiD3OB0QSUZYGWYUmC
SOp39aIUMJHK6cFNmZywX/7YW/0o/Pbhr008aLNFRfcUlztDAV+DJPKWYbrLLmeG
5ld9Bi85VlWmpdmDDrw50CP+W/lc4qwRMnFr7vmHpOJBiIxmftu+9E5+iY1FxP7z
PzLMK8L3eBL05vwZv6w4jOmi61Z4soJYS5GIxti6+LIFN12tvtv1k+GbIB3abg3U
qvy4c1z3dChD13HLV//4Cm3oOs41G/BQ/+KTYW3T0FVAT49rN99rE5aJNHXbfm8M
WHP24ENOe1IlrimxwCO8Sdhxrhd03OD/H5aDvX5XTV8qdedLaPi+yPAj/ZIHT/56
TBPr2Mz46vsGomhw4MMxrXdU7ZYgPqxKh4i17Y51irAUGeYYs96GVMA0l9GHLblW
qB8H+OcKx0Z2ARWi1oO82OnJ+OlPHbiIUQ1i+IaODO+t8krf6f6+obwck+p9zLi7
x1rb23A8thZBoQn7jLFgngPTrUPYBo3qnhweWBH/zBNQ/CBSuJoH1E/xit3BomqY
jSM2amde9Znsrvx9KspV3Cr+MtkSmZzTL4ROL5Gm+1TEo9eqlGq+vLTB7/02PH5q
2PTJSLKxyo0lm+vJ/IRyRxzakLdEhBSvnpdRAP4xMN6bFx3cHb1ojA03Repuc1Vv
vbt52X31Bkb6I5joS/Et+WohZ/bumtX51mSuWrGopBpIuuYV/JQOnyTsQ5YAVUM+
wB6wepUP9EqhaEzOMXD/8gxHw6p7n1hRrk49PfWuTyGcWr2qPDEu15HVCXKYSHtc
mCjooHV2JudFsEOn8/6VB9o4IfKAx+ZCBeaWxUjO4ejx38KJ9SCnOHSJxjz2L8Rc
QkS/iPiqnEpbdHcrZnTCYg94gh0CZZNB2nip4G07y08KBc4JeSajEuNKkFWzEB8L
yDQJIY46saGqkzOmaguCEyWmp7I3gCCP2rUR7hbTnmLIno/GGiG9XfjNYwh6sCnf
kz1ziv0Xzt6bueDJrKLsyx7mjxYR8NtHJkcAZUj6mXb+TTaXLYWH165LFq6ttNn1
BkHmdk6UBLyuKc/i0qrtqzWZR07xW266sucVtATCad12V+NT0Ke5/XP7P+ZRAbK0
ux0hLNEo0eLvni0QxnXz/sJeWKVLDvgix4GGfMPDu865wcQoNQaw9oOXgqwFvVH4
FXohve5bxzc/kVRjYq6YJIqNApAD4nOCdJh3RVjQgIdm91RTUtf/Z5p+7fumdZ57
p3HyefIjO6emUG0B/si4qGMC2TDwzNnvI0sOYpzexsvQrvLNikJWF5Cqwghoq6sN
0dYqetC2c0hG1z+FFAHNvib0+nr3SJA26/Kiqqr5vXkpLe46yC9kQ3tzEoJ5s5Xa
0I5pYYwrplmiOBp7P8c+sBK2fKdyUUbZ0GDpQLfLjOuTgxuDoywRvgNXI12g2CaU
7ma+FKq89kl8ORR+gUZM5HGHbeUL9fEWi+vLXS3LgtDiu25UjmkWrAs2F2tsXJWZ
h1dzfFiubPaOBChPF4+QzYKfsOOqNwYg0W5Xm2iC9kaMiLnce+mClOnsjqeQTQ/z
WbE/q/qN6cYH79/x/Ffdl+Z79LbrMmLQIrJRiPNygy92gxojsoyz2rheFFO6ScuI
g0tjt+51uLc0ZZgzgmKI9Oi7nzP+p6dOWV1Dik5DjQPpXDe0UgTeZlCQVo+f5q6O
ZSBTBMnLAPcj+O8yVjv8hTcK9Oeff7dB1AhDU7fKBqskBbtAethSmDmiL8FfEp8s
GlvWL6C/eSll8vkya/2Ek/TrXGOKk7JiC4DlUjwNFF2cJEnWI862tbdqw85mpf8a
WSnzSipJdB8xja4IbCaMM16AF+zp/k0hXXF7L2DSj/4jUD/n0AZFMVTYc1n0U20p
oH1HG76PBnSBQWkWZyobCJBxFHHeQ7n7FuJj+uQ8NMEpAjiCDz9C2lOSkBXwWwVs
jvhZ8JzKpDp25hCWXUg8pY8qgIk03rwllyuSpfgQxNWcMuJxVo/Fndi9/i83gava
xN19bGsQDWyPkdunxwl7iR/5WvYiffq9qyLeV8aWI/lnhbzx5OcI5YlxcifgcaRk
P1J4AElbwpUdsUiA4XQdQCSciwNfmu/1keJTYnWdoUSGo8HdfrSse4Sey4UWyj4i
ZI44+lXR2sz6XuX7ViKxksJxVmSTbd0xer4WAfrP4fc3MBgpCDM0DErLVyYbYM4a
AMBmcUHADdBgHVx9PmSxAqwbZ0hvo2ZYr18Ho6FJO2E99sbCYVG68p3XsihKm01w
xPuOcYIa08K923SEVEC8IZEyfFwB+Gk96n76VgUsRqq5DQuuxWijDvaZ6ymXzXIE
pOouidwXilO4exFbTygk8WaH5/IIoI4TCRqU28gX3rpmnFrAdLCrW+I9WF5W1Mum
0cZzp2W7aPKbrApCp6SHMXk0ZqToSZxkFYjsdSMpoSWoDSYF8okcRMKM7NyDJ5xd
LFzDvnbA2yk0STP/bTsLeLg4HcLBJxQHv78pmHlMjQd/NmeadiN6SyNAyJkdTyIC
7AUy4OnGlaEPs5Ym2BXBdYvF2dwm8/CCCDgoQCHv7rEIIobMv7jKer3stAY4vfI5
Umo4TrM9p8bHB5oHBKqKfgukIMp3kUJuQ5kKdyB1UNVIC+H48ZmTwCVRKFX2knXI
Vx3e0XFivng9QVnbQnMNu3QaRvrtrS3VIHFtVJU9aogGRbDHNHh40Ja9UBEFObn+
xJwuEKDyFdhK+OyU2HzAtIxSVsTyVOaW5kkTYA25bIAYg5S+Vpb47J3CutrEgKyb
L4QwDL8iMh+Hh7RHFtzisCjZnGP2FJG6O7OFOPwcHDuFoUDP1h5xjMYRsXcLTZF3
TahlKDVpp9zgdujzPZpiR7Cg8Fq144vzbfo7iHomGZyH+tlQSPSJDS5b21FWosA9
bCjkEl7hm7yC+6dd3PmE3qVF1JpDo5YZIkaTWfQ50NrqS9HjcHYp7FFcfJK9lPID
Mc0xAcXpc5GDN57qcMuMQ5JD2IXkFiqCmau4QyvOOQ/FbYzm9mrMkEfHpB/BZUaA
TmuD0JMf3eD2SNlwdQK9jI4DPHSHTYf2uprXPPElRslYG1ujCc3zhti/QVRl1VZD
JZPJQlzUDQIOi/xSEVfQZLkaAu4UYOvXsuPcq95XEHFsh3JZz7+66iUFoeUWCv5f
4I5lUdyMyPMWZZ/J0mlcpDuSR1VfCzZybfK6eAec3MnKYiByDjcagTUhXOSJ6PbW
tnOd5KFAkKy1maVgnBODIcxLiQ3zkxxLndQxH4gfwpJAoBSyhdL1/v7M3HNe+rod
r9DDphM8Bgs9J7QFQz0KSFFjsZLvqMWv93zqfIzHuh/9G+MMF3+3vHaiZrxjJH/Z
y/57S5dRY5u2vwMgupzsVMLncnID+/ZLCI6Mr9GJ8fq69BOM7HP0kNIhw5nXbQ1Z
0WyzSR48yJEoQNrDJZf4O5g+aOgxbAGJ83RzvAact8FpDJWC2Hacx8z7m//3EZuS
dZYadKm+ZlESCiLTst+8zQZTtRYBvwSuXNQadARYZpv43QR0GnjOkokeez2G9fCn
mhB/U/YZQxQdGix5xxwhXD31+axXyS7a1AiI+nEIRTJc2Wy28fPfTruk069XqUaP
IgqOZ6fuzURWaAkrhUcGWLy20uYKVaG6Bd9Bq1yYJOdh6MCCu23vGBCdzFAI6AYC
S6lGhOa16PEg3M+lARu7LlT/RClAboWia+oATmQzFCoiavjhq/yvSBkjVN/BKBfk
J21ocuiw9e5QIHEzDlqUz8wyXTp5kvapg2w30FuaVWpLGI/Fv+k2OO8Z+5YoJW6k
bXP58wy2FrrO9ck3V0q5eHpjDT3W1+2K5d5ScFZ66ST8XxsxDbVAfOOMz0uy6DBh
mQ6FRWDi3O+Rqm1THl5EiOofl9E/m3w65WFZLMujXyxCS9Q1NmXFbWj8TCY6fGHE
QgpnxVp69/jqVrbgP3LoszVeibyIgJgvQ8YH1a7QU+8MOHtUCIF9saI7qZh2FX/4
KcTxaXeDp9rc6nyviZS551A7Xtuhn3uxiWF7u3aT3t7yTA3hEp2Nidic2WB3aOex
i0QfO+NZQD4LhUG9wqJHhWFDnSYP2NDHeKxj/9EixOLEb1LpBNSl7j19UX6guiuB
+RYIHxqs5aLlpV+Rgu0gKuO2TG92JwDoleh61dAt21IS+ce8WiLCcuWjUHEdj2Gc
zX4Wwt/lNEDKSjmU4IoLUzajbkVm1bo1UPbcWh9nAndpfchplFohupsUkspeiBYt
MmQPc+G23NFcZLVuHZUF1lUEy0CMVAc4eLWuNEQa7B0nZRe3IicatQD7ePZkLecO
L3HWC40V2yUvLCYAolStQpMATP1FoMOHJz/Mu/dVxnyNgztoI/a4mu9/eUHhnStD
XXaGY0zTvozI6DO2nivyqe94hRufa+JQFKJJcOQKBYm8yXQtxBFfspKFQ0X38uaA
ZgwsIzrme30nml1q4GmXPMCC8Vw/gI4HIyFEIN3bqV1NHEdjGA4lWIcoaTqmsnjg
X5TebJ/csx3+eiYxWbXiR3rCl8+xE14zAryPtIvHQzwO7pc9UV6yj4+dE5xCm6qg
scQSjCRKm6BoQoAXAqFbHsIwtISQRGmD6KtsrDKmfmJ0zLXyeswPHAvd9nXgalXo
m947rDupGKt/iLAW7Zy8sFch0a9xmmaoHRGFZaaTXvx9l4VMl2282CdQVKjFsh28
m4+If6coSszDcQaGGAOYxI1UgfudQzFkN205Axd9obhAaqzDaQEkJG7OSqHPk/x/
ohg2kfPafaB7ZKGQdJEm9HLvxYvruGUra5MHQzu2M5I3MfHFwsjvWghHkNQBNmX9
gwCe9he4hCFbWxmq6cuQSrHxpE6P1o+mm6XnqQ/M7CddZSUmHjLHqEO0C7Wncsy1
KpI2cDkBVmsuI12siItk4pV6X0Dkaa1zg3wOuMEkMcAZXFUN16FZnAj0zK3VpQKL
/DpjAZNss81gJoIMLErhDpMdKi0Gb09az1sda8mZ7Vk4t+NvX07uscxwYTNuv+P4
E2WMsc17py7/2SOSFh97uHtVORd+ZOFkLYEsqRRTZqOa8zvOS5uV84a94bztYzgu
ULUotUxJ4R2GiiVai4oBEGO5SjHhEu9vscRxLFUsTmDI23wjTBGKL9JmwF2etcIG
x3k7BjMR13MvrfmkwYyXfmoNkRARmcf+3uJ51199OFX3SXEyfSPqdqkM0N9clft4
uUJ63s9pmFZNEvi+VLJVGZMOyR7gPPhfzCvqrQh75LuGlxN6cUp/up8bZ+xFmVPt
A6d1cD6U3/QKReTIzk11+ffDdmT8l7Sx4X/2yXyyCgUpjamJKb17DL/w1zZi31Ex
CYOKBwhAHM1+dQSeBu1VFU7S7COr4BE2VmvllgwTktfVJv/CQ4KeRXnMYe7aeGHH
pFFPSlsnWg/OumPs1RJRvK0A7i5IY8V4FfQhy3+zHheqUNAFmnsZBJ/povZGiUgb
YD5VLslWYB1fmVidC1F3WWDMyblhe3i0k+DfRKAKOouWlXFVnGu4mOuR26/XNbZs
WVA5zzijHd8qk/5sPz2Jxpw0dK9SpC1u7IEyyruW5eQMd8YOOqmxnVr/hTH05mD5
qkXfMb7aOvO8TkMfuzVzx26othEhcUSVo4eoMVCf9TKy+xRFgLqDZN7nu6wahg1J
d2ko9YLPxjacrXdLCKX/9dO+SJ4yytgcej9CBE96fOVzGTV93gqDmFfZnsgB8GnP
AOKvzEWNu49TC7BaEQYwgs1S/1zohYZ5VHPDzTwXHJSz1joRVIWmr6q8xaMQADgE
HQo8LorlBzYa1LtZugSWTBsOy9dVKv1rsmPY04kiyRDzYW4BRc0Bj8Ub10vKZdHA
nTYoI5NcPxHWCckNjRjlgX1saV5Yq2qDiwFCdwQ0g631lKNhRFRaU1jjhrgNlKXV
wY+7c6vC4opRly6SMTBFad+TzinY/Kcju09PttrAlFr0B4K0ki1qSRfr7nBTdaUT
KdULQ2I5hbVQJb2xzJcwozkeEhpCZlge08w/1INMFxa1ZlFZr6ziN7v3r9Lxqpb0
I47Pq4zXRwa0SEjBx5+jXoLbNQYMWOADtO5blkp1qgKRfxVhfLOdgrPwWKODF5MM
RrtOYTjjQGD2FH+ugBza9yh8VMcekq0JsBFc3s3UJAUiFcfNcivJuhjtgPNAUj/0
yvLuVfDH7vGvfqGjpecQ8tT+Zbol+eRw1jRKu8ggtSv2WesQE4q6vQ3m4KheBv/w
xMynwWzodT9lbQ1YAjMG7urVO3ptFYSOwAJ/MZhMHh9GWBgPDIzP/O5Gjog7kZi5
XGsw/DagbnBlcPyJE4guf6nkCTgosGqYxDN44nNTKagYcGpccf8XraRt3JH2kshq
8rGj40/TZ9WS0ZdgCmu5o7Q39HJjmPSJ7CJhwPiMkWzA3v5Uxp4irEiicsXzYadT
x2bdLG1+h3TU4W31Od8LS0Vn9K3Him5AzT71hWML8BUyD23x6gbFHUANbGP3rWe4
t+4BJgzcMxC6fI4xODWFb0YR8Sycd0VUsWLVxaNLmk4l4wS201AFvDN7wgMoHVQp
pXSVaDMM3PxMoRO9W5GBVQ1Q/e5UDDcp1WNtaSTWyW2y4GS8d+7AWK8QLId5Xv12
tnJeV1a3dg5cVeUk2n+9/XQprn1WPF71DZLxP81WDGY1YGHh1+Oz4RQ0rRex56wB
VQjD4nyW6KKrGudTM9U7UOAkli7ifrEZP4PRJ+1wAiouIyMlNRUKnHubJ6bE++HT
DOvrYtkRApt0ZvwH//96QxltkeMTG8m2aknGuAfidcQhvgs1pxQ9NBSe+FvK8ZYV
u809yqZWwuDaOolTzMYFch7jmZK2z7IYCOAOH7hE2UQn3aII4X21XjgTMAEhGdvD
azAy7erUaTFlNQOG8yPLUADgYcq5oQ6gGRstEoYjazOTpOkWAO7r3LBOOuHZKvQT
wLDfVjPJWVnqBycblMzQqi1KZbtltjEbqL73LaxTCLkH0zJ7WG53cdEUIzGffOLI
2yssuz6Tp4zZ3QQsyJWrZ0FPIeBBj4cg0dWoQ/PazN3pusGyQ7/tBkEFfsVOBOBg
rxGjTUunLa41LnjHRD9DlkoIOV3hssf3GiKS9w3i3ZNFw2K5SWqCWwUfeTHZWKWz
keCSXyD5qxR+IZ7Xr3qZ5LQ+xcU8KJX1VCSDjzrKH2+MqSH7jhcmnWOQ1dIISiRg
rjn4Do7MoLK8eyoAcTmWje6vsDSAWnddo6aCwiXlO0XiuIYEo5rdJb9pYM82TQ8Q
t2UiDFYYmOxKKLdmLi+yV+sf2COZ7Sxxn7tpE7wNUg4d7L5qFSpreL0Qxv4JwlGQ
Z7cqn+uh4NgpbzxE7ZQ9Hur2+UEYVEe0zG2tZPzK3a51SV7otJk57JohIdGxgEB9
dKmzrJnxGwHnOwzqAd2IURQRvqMFSrRmELJI7ZRAJLKWGlGtQv53mzDCwHGdqZXf
DkAanlPpOCPp+mlywYZgbyD2IYPnJQMYa94Wl7t4mqqz2DrrIqp7vtD1rzzH9rtl
P6t1xF3QygML1eC+oEC4vUfufBZscZKkrJfOjj4thWLx9RSG3gElfgYcRKR0C9y8
vcKXwYETT6kG+g3nZjabPwsUMnztLihD+zgjaYeruFzZYzXuJbminODBxfIZHTQy
1ry2AqtS61EkF7vgwPV4N5oPevVRzJZeobpkvrm3+abD1qeB7BoJBngvnx0AkaLQ
p8j04NPRQu5Cc4fSZ+0Gz0nIGgFswtF+Xjs0PUhOKhiNhxHRbzu2g44hZ0rBzb1x
WNqUFsoZ6FVskBaZZh3I2zLNxLlbdjdFU5lxdYh3RKcYcTCfIVGz84SsTUzhjGiK
UQbNuyoX+GHknKA+0C9LMho+laPKB5RTh9IQOvkE0tjljmysDC6r2eD6vZKtm+FG
t7JUe87EqKj6CQsznoV72cJU7GOOddk56SWjnVqoQGD4fmJl0kGLKGnxXcQj6+qY
PZ967DKKE7CANUhAWZ3tZ5J/GxLa5wyGwsiWURLSVo7d/jk/JyhgiomWLPos5ooV
RHH0wiEiURuIAORy8OUuli7vj80THsZBXrIWdj5UOeylmcbNi42BxyGrc8I70Afa
eeX+jojeh3hBz+pbMKD9gKvTs7RwHMkKn3cqqg39fVgjBz/BljAwWP6Ev79GU4wq
Ea8+oHkixZ3faLiuIC9MSIiikW3nLZpf9ya2YZI+BQq+HI0x/AUya7Vm1vNPcH7n
ZYUEnagtMtxAIqUft0/d3cFZ1B15GJUaLpxYJkXa1azYJbZD2IRmy7bAjHROMdro
qnXjv+4Ohl82kCoLVUbGyBTs2ghM9ePdjoV+NgSlRAseRnhDkAiukAszfdDXW1it
Ff0WESAjCAq8slh6Lku4i3q/+bXTFFjMpKg5IH88mq7f5WW4jIg3tu99ze7YjbQE
uWDB0skeM98G3FLxgYa/5/4nqNbnX9teia1qQbO5DqAB3broIxoeAoY8jGnNitJY
y7C2PVMqwsPnw+UZEP7yi6+431/h6ByrpqLnFI36njeVchHNgn+yOvkGuT0P23qa
BUCU8iLEY72zmpLVneJhIEH0sXXvkWfxhdCc1nxQm5Zcxpa6HFMLpnxPTWuttQEj
ZkXmTAo8j57lXQHbWdX/ktgnOOgbFJ1iLP/iE5BVizpiJqMlOdTOtg0Y7C4SjiMj
6X/C7sQ9i+1ySl+xDTOaJcBDzYcHb7EVDpvAT9LluYKk1k4DvHJrcOfpYS2GhP39
+sLGLmJpAuWDCyHD4+30x+8iBOkq0z9/m0b0iLLU8QbHT2MPwuyh3kMXkm+Rre5c
+3V44PtmDE7QJjVBpLbv7JrAKnkJP/rgH3plPvjJne5vlmXesk+qo2JKVcX790cg
mNkMJtRN9kRdmGranz3Kf72sAPi/FxzqvZOt6EJm3NS787Pn29Nzxl9liqYYi/+K
Oh/PePvR4ZqNiGU1NTqDDJP72rxQknRrH4/0/P0wZMDFtKhxvMMscMaWXcYVYJsI
FvFucmvKwAZLQREeNjKiKNQzaNQc0zXwAtBhqOMl/XGBsqfUDhIo4IyldGF03qJD
X4fX8LP/pKPDrlo6h3NsS08dGYYnLutaQre/ZVdq1IT8BsTjsjs12a18xeY3umQ9
JKZMDKez6CI9J4P02ORUSWli9sHhZEgacwyut8OG4CTITS/L6PLybs9N+v6+Hovc
/HSGWEMum8Mm2ji8b4GgK1PR35z0G0FCSYYh2jzFZT1uAt2s7h3pDxWMhP98THaw
+sOohwoeLD+dsxoT7IwiEcZRK3JGE0zu/vHJEdSZl8W21/qVM68y0ihdUfNe4uLO
rn+oIlCkw3oJQEZMwVgxPmboLP9dGWwq24tQLogBnkJ6uF8atByg5ygbIVraEiGq
jiAFqGeoupD7GEzxZtGP//CUezRHzD8DTA/TpO3rN+Y8Odk+mylduKzmqceBzh+x
jVV3GSIgiEi9lNPEGatbpKM0jabnDMD5YZpbKlIAMLanSRLgguApcQ36JZH7ewMa
0zxDRWoejvPApLZyE7THhFMyCtHrk2CoE5fsqVOyDZEVaAbXnTlXzdRGTguaKqm1
apZGYvE6QoVw9vtofUMdy3U64SlJlkL67MLiE6kt04z9NVt1Vd1wKDqj+47yI7zo
nEvCzBzE4HgZfzkTcswavqOWE/0NA+eXfmpUAebleVwS5LJraTuP6amhVFiUokd/
FFwbCDPeXRJCuV51yzi3aZqjUCX/fmFcIkMHfr8nfLYiTELkJtYBX10iIpWPCUUN
ofC7g4woM+nmhFs/FiuDBVS6Y4fdJjZG4eXfcvUtY+ExRc8NqOdq0KJ6KaDtn8xy
gYuIP//H7eSowdi9rs7+t07qo0WHYhRyP7ub6bIh+ZlzT0ewyMXqQpyiYYAPAWG5
pQUuhc1k0F5hdXfC7pCBcWWCDv9FmWGofB6WnXZQMREp4uO+YorPpHvplWvEJZwm
dFirIEiVj4iYaItsyT8QC3XN1DAqRAGlXXpODihtRhHxU3flNxDiPwuNOAYs9Ruj
BChFBqlWMPfMO3Fb+2rPyzsu5+VAlyQd3eOv0NnbY/Z7Qxq3d91/Xe9UiBmRpZPJ
DqLYN7pozw7femZIQSYjqZ6ob8lY0yZCCDEJVkcyaAFjB2nUP+y64yJGID9nNnUr
Funhr5KhkEZEBxbRVHFeJYVeACMLrzPHNdkAjvJEnuOEV4POrHVXrEnEYKttlrO5
qKnSB/UYsU18qgjaTNYD03QL8G3aUmOrI61vNlpU+bWrpWDEgb3LUJCHh31UlpZ2
AiOModdIRPz4NlsBMIcZ1+Ie0p2gWuqRnc2mPRW8nHLuhkJdUM1NP4j3Ac3dtwkr
Lp4eFpgVJ8Iy+MavhDxOvJYSDVPKScLPeDnNU46Vq9JZamxI/50wBQft7aeoMH+P
5qJWnwImKRhUEknNrCxWybsBaeVVnIGw+FjuoAuNpDliJsPt5L23+QzPe++dvogA
ARIwt6WWLO/B4mJUzL6Q3hMvLMX+o7QL2vUj6XGO+6qIynIZBbHEG8u7BImnJdEu
2nsMfAYux4XNXJB/tMDq5amTXKzAYAOb6VLV+A9J07sNcZJx/E4xhYqOfGpF/+Wt
KqV7Ra4DYTqbHmG97eI0AmW8wEnWJ4Ecd99tT0hHEVEUovlBDuNnFYgmISaDRgSI
qG1tbgoWEzp8qHuqTOdtg7aryapsVx2mYZYEm5xFRxphCJbCpJ7v+fXdaWMbha7k
PPrylcj9KHNRUJWB78J681kp1Kv3r6spdF9WVVFUDlMDz+L86WhP6YU/dHrg84eT
6bpX2AJuU9du9ORSWzKCUb/38lVwre7pJexaprpflLwmmdDdOtOt2VffwM2of90a
YnCdzqS6WaG8PP0oLGrGJPWcq6GVp1V03uyIC87U7huS7PtC3eL7gn6IqG02F4br
/MCNhPt8FceC2P0eTWPqTi+L6Ha+aUPagNC11HfFJdE+X0fSXhRyPWezgdAT9HUs
y0TdPJnAxFc1Z5LUIXgSwXyAYdgW+Bg74nV0MHzbNQ24jBB9jJItZlsUIl8vcBnT
yWnHGEr8B+NLA8C/toHd1msuZHGoS8VGnEWR9cjDl8XRTCbT8n7bI6PM49GXKp28
0arw3ormJroPlxfHIbfZlvBvFmnsm4OGFPwn8lQQWq+Y2GJfOQ/SpD38kFcHG2W5
phIEgqzbLxAgy5mYOt53FdHd4X/mRLS112rz4ZAGyRQkQflzVb+m2RpUKIm7wcGf
YukkejySF0dmjqfjkXsFM6KkvowL38WoVGzLzBywu6pugGfJaLPfg4kVsIJiRrZE
ToD1rpPZ64z8IjZfJZxUKUZYRZvHXcE3q6lMZ3UJRgbqv9SFXit49VDnbLH7yK6t
bTPFXMzwEsCsE0NPDnTR+gGHJhH906nmjkR5nxY0BXZnhRsSqwjLdEm8+lAwDxTN
flqNAlNL8aDrUZMtmNlKZCwsBrAyHcRoCAjcOtgcLCZwB4gf2UjD64t4AtBLjEB+
Ft1yK6NOu9yY1i4uziiCdsMTI7seEU+E58NtZsrhlv0QminG/KCE/vZpwAq8ZV5q
1prkV1ec8m+s/PjK0qMbSIoOkA8Cr/Kp7AGHck9wVo3GhVQ0fTtMKbsQTrf3wVF3
WpkLua0WsCtvqKfkpeayIE9fu3w47HNGLh4FM0iHKk0n1KzekaX78blXFZUgqjKe
Ld7tE93KEMbZXvhiYf3ABfSM29NY99rMm8zOgD5GRKkDs/AInuY4nUzY5jCzUJUA
10aukWxUjQaJdgp1cd0qi6yN3U0ELoecA8+1ylDBTYpJqcHWuYCARv//vYlK9hYZ
0Z+U3i8NZ1zTegPAkB1r7YeScW4s/3Ix/4LknZ/Zh4Sy6J4jqHfCRmtRA3t0/xE3
rgG/2zzFD7T1iEruZQ9JA30JTPj2W1DA+aXJ9N/ZQ66eVRU9LzMlCptLPH6eGt0/
MftCAJoVpor1vBt01Yj8b0LZ+BE0emE2Xolkp4c5ow4GoHCV5iywI1NOssCYpAFI
0c2J0hZKB/m/SAuWAZZpLDXPnl0kGLKB2Lod2gY/L8GZwbHToW10W0BIqFEHG863
HPMqjfvu6/9SUZy+cx1TbFwj2NGe0ETLwrp9/Md4UFSjNzoOEagrOHOg9buvT0e0
Js1uM6ZXZzaAz5Rt7xZ3JSlDOSl4ge00mGBILRLXGRoe3E3aYxn5P1Kh2cycXdPs
XfNuliGSgKgAjMlnKATam2+BPBgc52wcgRlzhUxBKW5RWUbgqNSNoaUss+/bEETo
yHDVCn9/UmFC8WjVBD3k052bLqDIS6nMd57H/L/wMnJnafJ6rsutcx5hb/ly1Zxk
dFTOMu8qEwEI/cUIDqFk7dCxxIWRoaxiFLm6pwovk6oj7o1f3TnzFFw1Nv9gpICQ
a43yJ8neHlt/uWD5qokTCz55APrlv050zTTQlM+zeIgu578OAgwRlIqgMglvj9Zi
ljs9X3B1m6z57dZDWfxGdJmTlkDWq+qIjS+bsf9xL8rFQ75AetknfsCeANMwDbn+
QdwOrpjDsfUIY3rj/zCx478PCJE/aEi/Od03NgACwisjRDq+oeG2TtxQvwpe3DwO
4WAzRer36nByG3mgmNRIW1cJPTPdsGPThR6HFTUNrB3mPhffrwZEhkWo84aZaPVS
Bj44lW7pyyyqWn493zNaxqC3f6u54yD78Sn9Xt6eknKGbtIoUYtyIY3FGHVKgORj
NaogBShQC6SXhGiOTh1bwg3IIIocc6tnJIgc2NyjaiHCvvFAJLuIwrwhaZr8/fkl
wG8YQ4BN7GO4rrOp4nAc0H5viEsA75LUdDMvtgASeXbyY6l852GV8l0R4jk80vHq
eM57fVOwQBBE5M51GfJuCT4KgAIAblyx7R+BUYL8RLRMMf586iPD44OntONnWyJO
OhdLNvqObi4C6rvBYcfBMyyVsCfeYAnQNZYsnNFmbsUGO4sKcW+22rTdXaAYLK6T
Z1SH0Wqp6aOGBQrP/BxOslniaYqfQSvu5Qg5FkQ57GupmouFInRVvAl893K1Tbhv
cM6T7GengM6gBqJfNgq8YvWin84tG9O7KYNAqvU86H0EGwN+y331uxmq/H3AHrSD
uvQgokDZ09cp6VCgvsOfE3laISIqvUGyCSmC640dc1Eendbf/XDHkXnt9WKRgKt6
mWjpn3zK9LDovOjBp03u6bCTJ5QgUkoM2LV6UUdlgebteL3OFA6NXWNlP3gz3YRH
XOkVNvTGjapJR7om+d7xR+1A8qkQ7NzpeHgBdQDP9ehRTCgA5w7K0FdFrWYwKt3K
H0IIasF4GtkYdTTqBiM7tv0yY7tGqZKkFS3SPeGHZ58zmkLnasxCJsRsGmDR/aK9
emTaUfv68UsE+bQAz/tZcPR/Mh6tZScpDt9dNbs2pPs3ClQ4nxU+CfwjjMcqOhz0
sFyFPIZCAs+WCCrg6xDDrLy5MLxisGXU7JZeODq3NK/APY2rQifaRQpD8270kHSl
OwxyCxVSlgh6Yzh58w1db1PzgCi1tA3+09Dl6EBB4g3EX4/EAfquA97/G8D1RLWH
p3YTiolkTwUJn79cvt2UrHKyJkVvhW7TposWY3xA4242xpdBsc5zBBpeEji+osou
biEtN+Ca6v0+upQOG30DQi0oeY2dAtZPpaxjgax6Np/AaAXalT1RB35eBaLNFp61
VGzfYbhoUJXcWKRwWwsjl+s4exprFrWNx1jCx90M8xWddY80gC31RKoNNMPqZlel
fcXEPk+r9CxxPs8PrmbuxEl8uzfHD5rulqm6OKF4RkdXTbcG4Tjr5TH+w0FupIgo
SFzFjdhhaKi+wx+cdR2Y9in0oTRvBJehBxInAzkVIe88r2WeKCh6zbq2LlsJ7xka
HCNqISUVghkdYldvK2ILBHhsfS5VemkULHPxNfhc8Ak7NAC5CctOv0icithssIix
X8OJRYuaSBwgvOYQm2YNOiPifTKhuJor0zLB2R72l0g+eL/x766hRXSeTCQWicCv
e1E2CP+ooAMj9TjDq64Sfh/GtmgJwXeXnVF0SWDGyzI0FvLFhFkoRJATvA46pe6Y
zTL+/+fQNvI28Frzum9HdAts54HhQsxNuEw+yhgUNsNPlpJM36QjaaECS3q6W3di
asUG1GShQUfCMKyeXhpjqJhkS8zfxANeo48it9tdnBJFlQqN/M8VuXBJLGowQPM7
YZAJEMLf6b96T0GPOe+bOapW6D4MMHiyb945bnt9QQQMTHyvA8PdI61a/ZQEE7hC
ehML9clqVNftG7VhYyOFBpNxrgVd1lbKygrqJ03z2WHMpJSB/ZUeD+kw6DR9x2iG
PZxhMjbgElkpNCXIAw8CV8YWAUoBCRZdPGR2ne9/rNCa9YIP6lILZyz07nKBGsCJ
pHq1nnrWd7iTmzQp1Q0J9N8AO4WcFVQ/f3VXTB3OSPqesfRh3BxHjg+Bb1UD8pkh
4EO13Yrc4ANYzT6oDC9RkoyIVvUNs2SlAi/e4aYBHTC814DkMcsZ4sEGSQW/hf6i
VJcuxtd4H1Ey2ZeiFMUWJZkdfA9woSze/06z4DBC++jxrNyu09dLd4/NcKb2bA3z
4jAy8zGYpe4j0q0uOdOJosdtiUGCsarDBfxwZUqVN/Z7gBNsV5VCgnRs2xU/1Odu
YuKDio1euL5dmK/HqxxEeDHktz+kUDr2QN4DFGeqEjTooEdPqiI9IIoDDVzeg2DV
L3vwdJ4xVh5ZZbEqSHNxFQ4tMAgZX8SyBcJJPYLZKlaecBj85+R3wml6LLS3GnE7
KULUq1l2yF4vTkayXaANDRrkGY9Xad8aWEgAaz3noFWSf3Hagc6rzo6zIeQMpJk5
NNdrJ7XSfdIJuf74AqoWKWaLBBao+6Sax6LzkGoQM5DbrsAVxNuxXo48i5j9g/sv
QOBfxyI8N62sLhXLL04rJIFMF3jL09rT0qTAnjqIPU1j4TsW5/2qDxXU6IcW4sPU
jaS8kEIEmlY88Do+EXsR7uhdfoE/dONpbAaaB13FrDaMkEM6zUaGByToQh+iRBLb
R5guYsm4g9Lk9CSu+6LbGWu7zVepgHoH2XlOp+hVKK24lyQYEHv75VHd8zmqbQ0c
ePmLxmv+ftXOBEuyhWRS267sThtBl+OTmriiVOQlhixEOr2qECjiVVQHAd/h+AhF
O76j8ZZUcPJ27WrLgMhPReS1UGPTCppLsBoXPaWNJ9pxdXJqQa8qE88Mb4bQVnRJ
sJoNgtWiILOTsJuLmbM1avfprpJ3TGW7iCYoHian/cXuWSHeRZQPOfRsH/DmR1uh
7GmmAaGntirioklypvAOokNhGiXvvY9ejtegvhA0wUMw0y+vkuHKhRCt6FNsIn+8
E7edHSLRAU/F6zQVYlmgPdtDfgZDuqmQtIR/wBrPyAhXvOa6PtWfylhboF5c961S
GR/v1L8Z/tARBumye6gUmNbXVcSCSGxOb91/xFEUCYInVmprFRlX/K8s/nGNOp76
iYdGfA6QNhGNnghK40Z3UlGfxoX6rh5DVxZDONARbNev8PKExwUrOA0qVr4t6j3A
fSzz81/Y3lG5EeftgAXjI7qxs6Ak6IXePXHNHQzRguWxD8EiM+fiF75b2L6d40vz
SS+IcOEk6gvti7AZm75yi18Hk727yCy/KhV+pfOPO+PMQZw8Ff1gUjxrNkkK991r
9mxNm/gDwmB2vgI1m7mOSRtEd5eWSa0qQ0UyKNQPlOc2qeIv9kBIZsb+NjkPJxbD
rLfgJ3tMqlQOO+ZiyC+Gx+GeVocjdVlNvwMD5aLSLHIgZBjv6QwbCQATKILody5s
kM2gelVxgM+2Q7mdfUAtbvuqC35AG4CIHt28Xr4FHng0Ea9Wbn1r36u1p8/13v25
padriv96II1FaOxhjYmINCiuJLYlosjQjT7JG+L9v2vFUYeEZ9aF740h0BW+lM0D
NxrAQw743iGVcOjPAF4e76iB2wxPHWUk1t1uQrrwtZN1JD1nE7fYlvib4hiRVGPT
ArMMKwR059bk7XkSKlrwFuQSEGP3yi4KtWTDzbHG/ryBCQLPP5XcczRUTAwq6Luj
TLPDJ9qPC9lUK7D/OHfN3I785ollhoPCvPcoF75IFLK/nW99+0dBFXhf6qbSZwq2
CxOLoioHikI+TJ/nU2cfXW/8URJN99kWj5/yaPdiFVxmY51EC7HVIGHDhDmjmoPo
4chqaphSR6ghaU0s/q3DIgQAN6G1M/ly2GernsWefPwsFF2rv8lcQq/uzYQnHCZB
rqxxiprJ10bKYfnSeDdR2gbx5WJcl9Qpj8tD96faolUIbmzGvHhqs3ASDGBUr896
C2aKs6aTBJtOvu4d3LOeQxiBxxBq7amUGPNGB1UhkAWgLhBl/gxoP7fZAEReKoqo
SqXma7dMBc4QysnUk5EDbyPKezUvEZzUA8EaWowdJBQVC6NbuNo/0gl+VQqo35Xf
Kdodmd7/440NSgragMKUsOJ2BijK7BVU89/5mIZsHl6J1MxTRa7JkpCqrQ514xwp
+HN/YbiDnoqJVIwIYQ8dEdpuxxTV3q4xiVUjUsrMGzk2DzWlOf3NgQtI8XKsR7xs
vbhMWig9gUMSvWAFyiO62h7tI65mnclH/bkJGL1SRsn5YMs4sr1sXJ0q6uneZ/bu
oBN7kikPTmUykE9lu4a91IsdvWuLsGcZUaelHgBwU6dNbFYTTGJRx0zsqqIZnlEP
/FIaXuA2HUmSxde7z+wbIJXjjoniyUuNyQJ/U9iWN8s1ud8SzHZ2S+X/5jnhWEDF
xIyemuuooB80RPoGsj/u1exsHXIhwYYCR35pPuJc1ehfNXBwK70S8xyjYF7p58BA
f6/W3Ka6fBfVoc1sK0+mxK4rQTSHZEXM3LCMqtOU/8MTaLZNaqb2FZbhYSE1CNlp
bu8BG9hCyJ2Gmt6GZf4ZaPK7tObC0CxZavqcU/nMKBW4sceV3T1jCDGt88Yl0+Nm
0Ery75CMZ1szwSjqFIzYuelBXMLRiMmvm/vxFSRPXiRPb1IxQysmfp3ElGVTC436
a0+EIGofZB9nHjKPhuufBuPBec7Xa9ANKTP3YNfJdDH3CdCHUWNX+KCYQsQrWhQD
DlI1l1EoyFn5T5yz3xh0Uezd/DhKz9daO1uD3ton62aR80WVfAkoS5Ro35AKq5dl
X+vyFSv5BIxBR5R4ZZWVIq/D0bwiXLp80uDSPIyZc231x0JW9xQkQ744moRRmziC
oAlYtPw7fthbua4PGLjcBGLITrB9vDoQboLGLBlFPClJDIV1MG8duvycSovSAQpx
EbOind3zeEinG/NevPvAF5TSTDqgq1TQBxoOcY5Gp2rKvwbgaZYtZHe6ZGo749aj
fBdueMtYLxaY+/JXWR1n8NmGg8+BkdKPYi0jiCVAEdZZxCXEgkzWaNYNb65CKZA8
zlgy6pydthckr+OS1XkMFA6FX64wFMjJtFSFzt9bff9pLxZ9qU7i5KKqXjaCsUf/
1QRMprh+r9sMMXhOdVXcyxFhm3kQNkwkM7Ln2RmINQ6tKfOOW5jfJQ9McVDvITj0
8nOPpTY8dYwK1EAV25KwLmatuc6xHVoleWIk0bFREPShp2lV67M0zyrqmuyR2oNs
Xl9b2oZgPhV5qaoyLsrwSfF86Gp1Y41wt+1vm1vUtjtQrGS2h9xJi42/GzxxgIgZ
pDFPUJ00TdZfJGBp/BThQB9zayKLybPeEj2tx4Sjfrv7s5BVOkky3OMqMGkki9RA
/mbs76weazE1NBzoTJgnrA9G96X7+rlH5qOkOnMcId//Qo5voLdmljmq1T/Ft5DK
x38QI3u4dkrXkKp8g2BNA6tCG8lIRZzN+H4Oc78YJyN8ZW58p5foVB1nEmA9P9lG
baQyKn4vYlLgmbBTx9NfBYjuDVIvpStAqp3xptOKBNK+Tc0BIYkKyrsgIgB8F7nK
wErnpUi7KiEN0UWSwGOl8JAzCfOz4NPaqFgpoPcgwEc8JTfnFeYpd5Ut+tRkHRm8
3O6gGpVQwqtURNMsIuG5H7oKD6cH3sRURmwBPJrD2yroRyXTLTKrs+SJ5uO166ta
ms+Msgn0fuXok7N7IyPUW/MLi29esqAVSRLJm0Kd6OA7Sy/9OeRlI2XXiNuPm+qh
3HxoFQPmUI3AhUWG4MyzG7Av1FSq8KMptIR+NcZY94Vhfx8gspkuw6uj2948QRbJ
V49yZ2ZnfqlBN6r2g64G/2NJKlU4S7vI7TDopN/rIfvjvKtemndm0lbr1bv7v66Q
lnoVu/LWa5UV7iw/k5cWLjpLoz5h0YCda7ZaEVXB6aKtE58Z/jgsXKElstoCcsAJ
CTu3hfygPz8hgXMtYRG/SxNC8rf8I1mH8e6mW7ACX9j8GMPr+PLiBfET55USkdmO
7QhVHpsKjaNU+u00/ttabQTH8AUYN+9ugdvfzXsZzbcAKTwvNdwcN2u1XKEpnhsO
48hZijVBPHu33BRzVlOjg+sugABP+zGk3HnBIjBT7Nt9CEw0M2W0bk42XFP/SF62
KURiMma8Uc7IdvIBYVjzeRx64DDKlxWguRhKPE+DL8KDzcCKUTKNFkJdOcp+bJCR
qLAuNeKi1DohXPRrB/aZi3a4HlYXkrwDcFo/BLVc2woyJ3nSa/XegkjgDhqxNikS
dFbcUzety8PEUd3JPvBeF3k0VM4V7OAlp20y32v3x9oR4hTkob/q+QhiZZ+ULKk1
sm/vdRvFETytW+OGkaw0JegHbUwVHliWZpvh43xvzhhvTZfyzw+Y7cv7YwnyRseK
3leEH1gt+OemTiJhhR36B85l4NQQQz6xZFpXZKtzxOzFdlQxUClpGimhw85ij5Hx
M9KaKcLfby6uSUjLQC+LRqTXjsSTKSyK4qJ2r+ydZwgvvhlzhhh/JcoIDxd4WEZf
Q5c2EHOwAUS840pX1jCAOqh+l/pCehB9VxWHqYr/ifHANmWZe6pQzMAhhZVmsMS0
xyHgLim3M8vtS69vRhlqDCfP6C5yaFJt6jVIeyfDElXcrTtBhVrA37F6ZiYE5S7U
+PaNYF5AxjY9OG1zk/5sJH/G8k+DNlTivsdVyDmHPxtorUvHeoK8zFUyD21K+AG8
2kjDRFlyRGNKROE4oRw8Zj4YBIDMxXBfkzf3EfKCj53q2AedUhBEs1hYbvkLg0+2
s5gO7k3co294uhDsJ8idukYTLzAQGpmaDcxD5MmL7Ti/J2GgNTjq4CKTlFvU70tC
8ymd3WEsRPpbeetvJZ2oNKW4ov+3Q/ubl9y4DDvo7xfe73XPAZzeJZ1TSox1aUjm
Lu1lBAKA9t/6Rc1S+GvDs9nibTKxoqlnce3F2Im0eWrGCg6KqvktWrG0IHItJFn3
DrAi60BHGz/TWiZBakJk4llsdsNIoHfBIz8hBxWmDsWbLJ4r6QRnNqJ8KdUsn/IZ
D4/BmLw09eCuKM5O/bN+9ggEikeYlQyaUmQCYbdGP1F0TVnvYxT2JDDq595ftYc3
p27a8nrDKYrkI5YjoeI42FexSPWDPmiTGajdkKTlGT82zMfMmnCpvlVkg6ityZej
VljMcTyL9IQ6sJ+/jDlY3MIHpax7ExT+cWBDD9HsFg/7lEkxqwwpWxXyuth+T6QM
Xqa+eEjkSOQeTAhW+gF/d3tULOh3sX/ZI5j01jNQHPr5jllaoiELZBkH3TPwueRE
n7GCPZO9miX31mW+ZBDeD1lfj4GAWak7Vqsa5sanVcK0XfnPDuQdqKTDjx/LcUrY
0K8Jpa9a0jceJ0cr3SzRenU6IkjlvqfkTfKQaW36PiFXd/Gt81YX2fdaOcXnsGYO
onmzoeD18x+YsNPYqfE/QsXp6rZZQ0fK0bkKHPYynMG5Ub1v/XhFBK5BhP1WrD3Z
e4uV6tM+yepSNphfcnWXrJFwom3Yw9srBWGCDT548XXRdXttnBuLFdh2gbAEPggc
O81BGiSvgAhxgW4J3+AM1ULhppixhBTi1y0R74tOYH6Rsnr4AbSqcudwXEea6qKq
94db4H1RY8m2pEMenmw4WHLScSNPOVd96lDolfy3Hh9T1WIDrGekylWwaPZGUtcF
3YflBsmbtMPDZjDUCNFtwlbehaBfweDHpBp1/qVP331J6EIid14SPYB3ezhxg1i9
czXsdyZ9q187aP7TPuUe9/FADAvSfbkCjQbN9gXZbf09QM7dLycLfaltRc2CgkVd
oXgwBXBtlMJCMEeTDOUtcnoFB2sxj0k62LW/fC226p4l+P8kTVkCTuQsNxMgaX84
c3/jq807uEummQQA71eqvIHBy+giV5/H8pufOR8NGeGuYD7JD0YShNqrOIDoOHR+
Ny+/UXvK9sPwstZpQ5niUSrK9yLrBr7R+MvbsXFzMv3EcOdhb0zGRWS3dQ2mB9UG
ds8GW5G8hJMiMWySTqx7V73K9Z+Vp72Cn3WZvpIws9LRk5n79QNmFl3TTl+4chId
4PwBtg3qMRyUNn988DAS/H5tWIrkHIljCcuazpWuccO35V6bCxuBd5w/3k4Sucx2
/4uBvsN0tmHy5nTsgw0ZxZc8/xFjbSPwF+T/GM0lj0wsSXL/9yHIFeo2VjWFS7Vo
ePX1LZB+L0bMG/ziYcJDsWrt4/y/AI8bNvYcKGdeD4HELeFCNqa9+H6E9CBt6JOl
EuNG+cU8GVSajfm5N+c/5ujxLpOOf81BOLjIfaZjR6+HUak3sxohLylPiEWH42s3
j6EA50ZbV1DrDj2ixnFdVkjZOfP/ueQeWWLIYBm4rFK03RqpZQGq9cm0qY07gL7m
9mFXn7XifFCrxwqjnqC3aoEj/jJ6u55ndqkdELwF/iGHv44vK12ci9s8q5hTyKhD
t/yvlVIBRF7+sawMFE4b4CC3ScCfjvaGQ0t7gpsp0X/SLGypvzZ575aIXgDkTp4Z
esh9B3AVQ1HuZkicPxf25TFoTRg09EBQrcpFiSSG2ySdAsjQreA8PkJior4N2ehw
J+lfP6Z+a8NjXWMz/rUulPkKhieFEFKQBxVY7faFnKHR8ImfqUImld8tNh6mbR3v
Za2oGFKKDoAivClSHGhSR7atc8diwlNfLSLKVC2SosCahjAJqRW4ZRe2Rdvp7oCI
H83d1DInUlE66GjUWW3BE2EKSDUKyZJhjTnfUzIHAINQwQHebWOOxq1UG1Hli0QK
Rzz9ge6fPEmqguGhZuxMqJKGySkbY+jfyyV4BVjjNnsuAeXRNginl6ay8knicyWV
H2wnXB3H+E16+sv2T6dYWr4AnJN/tS8nfSGpX6cXWrZWWEgoL7oDBvhSzJpRlVwm
ynPGTCcDzBvzRY+fqKWf3MvztPzvNYuhM1ZxHdm/29sBgssiN2wxVrq+s/QP7iRr
y9eEIiCmGq9s75wNNOG6JhmeKjC+ZnuvQB6Qd8aQkowWgIfU/VE7FoFoWqEsqWHa
8W6GekuxekE4RaDhSNTohK2/5jlOHBpaj5SMBZK7mNNdOanmrB9H3PBYadhW3jXZ
4yeLmRj8SNBvJ21woKQEhKFFYb3Fn8gueL/tF2DPfHne2lAGpX/Bj/ZbLZGoTIyI
tBYgkVS84oG6eOxTdkNxykqfOb+Ebie+0OLKLq7puIEkCENSPo/lPLE7Ej4bDQhl
eCcl0b+7QrJw6GKoc2QKnS/ivK37EeU5oMDSpoLnlYwOnV1S/S3opcVi/QmZR/Qs
iUmnPLXe6t1wL9kmZq+PIlx13e2sLjaYswsZaMOd8umbNK5A4Fn511dGXcgWx4lh
fH5qZlXG+tgZ8aO87uLnhTOJG+JcKcXzgAlvZr08SIE6ziscNmKAhYADNByiCl98
kUCocAJk1VOTtHJqGzfM50ZbTGs892eB8DtFPfzK/aDj4islrKFBj1qRKi39SnFb
UCtPiSur3byg+7BbhZOlpWEcmoQIVj24bu0Rqdogyw+7NoGwbXIDDYJd/Y49x1t1
a28AMVXAh24yvDgSalouU8lrjDIILOuTMm9DnaZI3hRA+OBxQuIphcKS/UWYR643
01J/XrJzW2QRl1A3GxXIxeQu8HTc4nd8shU0Ej+TjJMAg4LteaLKCxW0x1SJyyfW
8zhxM1IMmVV+o1PwpMrqPDhy1cVfve9fd9iXurAQr92AaWmaYWpAR/CCcmJfTB8k
7tIE195s0Qh91jYrTJ6D+eyQ23Zfn20L6zxZLm7+/LpchDAnelzuTjcmCt+ZmpIe
ujEUGmFeppkA228fhij8TCVyFfbrk3o0GDIm/Ctcw53DuVdRvnVdNaBVetSpuw0c
GqRBQ2kjPaRmzoIByB1i0/MMIUHRoZFiino9gw7IB7A05Hcom6MqRizv46bTw0lU
D2IGqDcRMd7P2FjJHAq1xI89/D8iiBeqERzvR3x8VVZmgamGrxB1/s7xKgEBMIZl
Q4Zp3kQ49iwHw2TqHLy6pDmLqI5BCdQVWOfD0WdCaaoFFxeP/OqeQbXth+9mGpd8
lmc64f9OI/JAuN8FO6qL1PY6LR9KHpQoeWBleLsCZzggbM2EVjLIpUJphiG1Knkq
5s5gRGFsarnoTea8XARsSD2EAPiFg0bGCraNn/gOhOssQbbYmGE/UuwO1mI5iX8n
VmafDFYQXquBja/NpvqaraX65teHpOWTk7jXkWFM1LgK0BguTnwsBEQF7ZH10fW/
i3uD7naPurXpNA0xozcCA8XKbq+IbaPOmD6EKGyMW2mhsdhO4d7Ipvld14Gw+G1a
7QN+rzqbBlS/aaA1S7anvX9UAKmv0IeOsIMbNBy+p49sYkuCK1m9yK3T0nEuS3mn
WP8DQt70rG+IXsSSgGql/kgQhnHqWdn+21/1YxGMc8KQf6rsX0VB8AdCpKGOjWf7
gBCX0eOr7aBHSiPTj644DQu39ZpL2gPmDV4nWwofxUEz3MhIQImEbzlaXenyqNEz
EbeOOhVk6t28iNujEn5X5RFn7xrCHZXVJ/MzaS9y2O5iFHnAZsvdEBMX5CRUjhLl
YBrl8NSyEDinhTtTFMjR86oBlOP4VvxPGJtmq60Cx3pw/Y6bOlnQCwqKXyEdXGnJ
0MzW6NfI3+Z+EttARXiK+/7qamyeXlwN6TUXJkCf3BISX0zSoWkX8RBlpm8RHTaG
N/mwbgllkPyVeM7p0cdlwqPGermfj/TvnRXveWz9rRqhqi7CKaXrjbYGlgJcFZuP
C6QRKKZintRZ+zzz9XO3eVYOtKtQRBYq8UBTMBQWkzuv1n0U+eOHHPE++HVi1vVQ
WJmthXj6WwMo7FRobM34KZKb1U6NZYEbeStl5Qvkrbdyn9oMiqT6mIKKjeSZJXOR
CA/A8/XD8eVB5EGClA4sIA633VIJqB7AjuCbm4FjXXRy+a+fzSWhinMrMOO4XrjY
kiWzIPEkIwDZ3ZEVsVRlJE6rypLln1RwQkKu3pg8SJCFVVn4J9D5uRHe5TpSASf8
65cBOHerQdipXi4PSbW4u5zAAybFAbZtRw6Ik235wHdzh04k8EOA6xNBZeMlDDVb
NhWDG4o2HrBf6C16FUPFnmUYsG4LHLnlS57gHjqZFOsxxWOB/g+D9z47R9+aYPAj
Q5YEqPp5TYOQljqhZcFvCfGrnOv35rI6gnzTw37W4SJ4tChlltTZ2jc0qqL8AkbY
kQ6k75yusyp6SD7rXiuoO3Aw3XnP7r8vgmm8Jk0TdGC+aK8HE98xXpB18mxjLQlf
bpHdTuxP+XNdFhDIC5izk9r+x2F8EdGl5r/+mjwY5NliuPp+6kehS6xytOLdXDuS
e6wALu/LhKaTQaS/Mj7cBwU04w4VfrV7JPAewhxrQEgFIPrPhXyFPLMPwR/jLa+W
zTcB0c0LeF3ltgEewkY92gcwVO9WEPYIQHIAyr2ya+9VTL7Bd3uXvB+xelS0gzUK
t0Ad8zTOkIc26TFIYLxKQYJ8CpsbfGtZ7q2hrysdg8utesEPwwY3QF/YVX+bP5Nw
iO8ocHCyshHo/6qJCR03CYekMTct+FDk0q13H1uBuOG+UU6sU1Utvte2g/r0fVo6
NXKC0JZz/4l99Vl9W3QCqVwl/3D3bwFDayoFyGIbtwejTbY0ei5I4vwU+9d48acx
ghJ7RiraK5vwUrj3v/9u3dmm461nFCTMdRO+Om5Zci3yxgYBzkIYLSapUAQy2Wck
XIMTOahhj0yfkj3H+hAYgO0z+IwmSxH6+S2irAaYvS8w3rSydZclwmjhROEaRBi4
3Mdc3bOUCfNxdPYhYvcS4JrC5mKeBbtFx7iPK+0+/xuznBhqAEy4BP6bwVWhI/68
YT96Y/+JPdyVrzb/NNtGGALXIhxd5+geAtaDIv7CH4tJNmzeruyKrMFkqxBtfkfZ
TDPl/2qlpWvJfFhSkHPawEWrqxGNdUxtD/QbwtanoG6eBgd7qzo9ksyOyqyA5fsu
1ETHPA92aOTKCxh+2hrXGjC1b7mSClkG44FMsrqt2L1djNoG4x4SW2LxnPmfe6/r
2N3P67Dyc1LZzk0kNzaqIxoFkGnvlRN+xqb2d+LxwjXPNUKTyTdS2lbnfa28cssM
vw53VgepZJMcfseF1zL0QhvQaTF8Qmi05KumiL66rdnsU9JccOY7RtCXQE8rh8k9
YWAlFLneAaDCh9d90DYS9Lff/eZ/jPLkMYoRAG5T2/GGr1TURyylJjx6vM7i2ZcV
n3bOKFizW5DDumi6exk/yIq4FTkMFDd5cOqFro1bWoWzG2tBFegSuNkvL4zFrMAW
pCS0+uIRHfvcnBr2ou9L90ESX2zT5DQagmgRvAI3gi6ISwzjdUPBTNjAZMgeM83l
YNKyqdKRjBwkK51n0YuXhy/EU8GasqADmVjsIHdQz4fE7ClkJjFSIjNiv102Xats
c9jXyHACGaGs4FbKpyupQv76r6uZiovHvY09wfCLmgUk4qN7ipUo7quOMWSMpkTj
Pq0B5TzYODH3J/tQ6E3BfJuWUbUahar2Z9D5ugjs3fF/qOK/fSUsFfG85CQlg+BJ
U2t5amq/8HPR0/tEuctM4EQ6pvFXMpdgEZyrSm//ML07JmfUIQz2kfe2ER0c0IJR
cieOuYpO3b2qDadaK3FmCJe+kO6hLpwe0/EiVlLjtlJrewGPiIVpxzV9qXj5ch6i
Fh7U26FHRcdO1YLdMH2+Ct3aeoW5h18NFzip3JEyuJkKTqqXf+KZNzNpNLCMKniJ
5kw1Vf/PyY4wAKNN7G3z0YvbCCOVNW9U2xeivXaGADlIPFi7NgSQTRCpbrygjKtS
5uVIcuwf6ahUyMTF7i1k8s67+dGbKjoTdb06yAbKoLzjNVigRUUGvo3dnownyP/A
MIwLiv5vUYeZbXc4zZ03sp25q/EOG5Wb4qrnLYQhPx4x7KgxXQZL22K9gHWyY2SJ
maYrb7d2g+PIaAO8VBrhyRw/sLZVIQ9p2mAClCHDFe4PDbYXjNLLJ6BPJnt3ZSnd
2Ugl9YEmP7Ocs4y00NrFTydzvG+pZJhDlcJ+dRY/kHPUJY3nFRcF2o3iJxgIMDgM
mIhtfUF8BLfVYOvJSbjsO+uWQ8V9HX7iVpYH5+8CZxEzvkW/G25ylEI4gBAqfV2r
fmElkBzwKIRoVNi419JuN4/I9IvelEZbNJ3X/4ajB9gd01QaHUPhECpl2Efy6gVN
RTmpk4YhEk4n+wQhQm07aexsv2j6DLf/AHh24D8a4bMvJ7ePKFANg1jP2mtWHcpI
Un3TXmES08Z76ktW0pNxIR9fRv6ZIzII/JKAFLuRSGVnzD0Sccj7tI0zxVbk+bie
pNTQhZ6WUOsGesnuD4LxrVC6l+wBV5dCmyeyhIKooEIAhaLRHoUbInVUCWUafQLz
c0iTfRSjSY+rwr0lR7wLlurPuCpp3msrcVprmiRDpN5xvIjG4h9PYmZJ+vXKVAB1
jCuW5y50MqcJ5oND8Cz7JB8Qo2sQFSgS4Ed4PGAOBEA8u2Bj4sISdISMdW762ud2
pY6atkyGB7LK2ftEo65OcQACNxRDmBLHPK8mSz0H1KZtppeeVVuzrsJIXwCxICxQ
Yzp9xy4eTSM5Prhh2MsKGDKeWbunXIh43DKbeiwMs1T9gGt9/xNFk/+RYMekf5me
NkQv7fDwSodYt9GLJpLpCoJPS7/sfFXGPEfVcHFtdhVQE63WRaMuNX67I45ICgp6
UaMmvCqFV/IDVu3bnL6I0MhLRB1isq+1mgCwFO1hloqLzXaR0mROg0bDetIb8GKs
cMFbbcfkc8rpIodDyA8IYHkgPBJKlX2fJhzN3BRJarQXctCq2bjDI8xJw7yivW5u
Jj4hZVOqa5ENSkHF4Eix1gCOJEhknWYDhViXh9m+7QxD0IHJwJDnbZVKcI/PzxKK
WWrWISX4XTjJhUnRF4jUYfgU/N6SgUyG/EVSmY0F6R43wocSgKY/xWfjDBGPs4Ge
usyj3y8i5NFQ+uNXkcEYpPGe1iVEFcSVCZxnW34aeGPfKyTYLB8G0a89Dz7y1I0O
SBxOH6ZUUlWA+OjWVI+QdOG6Y+foyvWPQVJN8Q3OYLRWYagwi4UzZE4aGnwZZ9c3
OhwYase/A79eccbtKmg1Yb2hcyzj+YhSYvCHnCK0Fao1W88tGmeC4Q2nPomGzb76
AH2FmeYWFV44Lh58pijIRuwM7BSQs+q6rsr+50zF0qRZMNkE1goTMZJ0E+WuJBU/
NTmu+fBGKCMdKvrzLTYnjbFIIcf9/tQ87WkUWf260imEr+A9jlSOVRZ9cbb99/Md
0tGv4k9PDA3VaV+lASm8k0TySuLM6psBFqoktRQ/a0i/wnrChcBeKFy8/wWPW7R2
mmMg4OFSveyem+zYa+Q7ZALKWdsTHcxb0ju8foTB4ZaTcXX5PpyBs0PE1I89GOHQ
IpjreBF39JVBqyEZI/eiwkHLpklkQ29329q0T1c8ICpxesl02BCnGt39WRs5D5dz
zzKbBlUxa6vTZIhj3I/fXJU+gEMKFkaHddo8TyjY3mPXtv/2mk6B+5h5t9cvRt16
oo130QV1drylM61+Vak8HQSRv+TeOagLOeI2fNvGKbcR0DcEyN7tuyS5uA7kWm2H
Ha1eTiF8UZUlidKky2f6YLKBIIohGDoGGODZiSkNPUeai4vEIP7hWii49AnHR9yv
rL+E39GwjEfdX5mHW57qeorbJ+Qahf0Ctdzr/e+s0rcFDLr0hne/hzQPcB/kw8lK
qJJAY3WP2BEQG5KwKIjA436zmc4Rb9CHRvNE2jbnaGkb8rC6PaiaBwMGQwwWKYhC
4VQIjipgjWibqF72UYJO+Dg8Mv4u6JshBHVjfn0FHF6C4SKz/lKYdaDBMvvhS5t0
EPVm3afLhxLX7uUDRG9oVNmdvElIBRC7BDzQC1ANUCQbw3qWawav1jTHOADd/qnI
YGtkAvUmrTvWEy7amDOUJuNxldcySL8F2oZB5+iODLKBJE7t5C7AM5vXGbnv1fJW
XD4Hx3BWhmhnxXCrlZwDpPOBloPNiLETbS8rXH/yvKhMmotbRxACG1Iqc217X/os
u1yfaAgOOWwRMc7ig54l6hK2N5ZJ7my4Fc/pQ+qk/kR0tGuP5oqmKuLqGgC6MOUY
mRWzuF25fRzn0Jw2us8lBm/jLy3HksKV0zwKBXsScXfwyd+lp+MPk89GnXokUfdX
RvyYS/KNjXRBrp/eNGAiZLEs9scCkT7IVQ9IzLX86P/80cgtzLGl9b4MCSZvx/Ff
SXxJMTPhnoa8Hi5Qj0gtJj9PyS5Vw2YGz8HKLCCylKioisJ4LGFlOlk07RKnT3oc
gQ6QQbJhmoLbHRwojuI7sTC8rFaqPpsiBnlY8/HvQQpXFSVm2nZUiCpeQVNsP64C
VyiYZGiK67XGUdw03So352clB3SyHtYjdkU6dxn2SFm+WJDtHQ12lsvER/JpVs4P
Ceo2V/oqxWc17PDTvFYbs7SOzVUcsvbhBTVQezmIvHpvI7OiCWxzUtQpX9Hi5tmN
4ooCEoWEGhbnHhTqYhcp3Kw6nZqWJM5l8bpqVbuVb+GcoG66TPfVo4u/ie21cQfq
QnbKU+CWRHXvw3qE4GlVeWnIxIAT28sifH5GCJJPlQHzQlKv23c+u4MJv9GWwL8f
LTlIySYAuISQ2TZ9ZXDhkfc8f/q2P/PR/ie6T42/HuRhh+CRjYRxvBdr3GjDuPmd
Hh5zKtc3VlobWhso7ytEgZbYUjhFANztaCC4Jn36vaEwlbNtLpMLSOHjhU734x1K
RA7H4aohlOrruRKwhHCYADGl8coRXYka8ns5d5ONgY7ENVFxaHlZGPcvsFocze0b
kFphaEzHR7hR99pYJ0evL+aQtrhjzXDdLzuoqRMm+Y2IlO7NvMiUvg1nhUIV3U6v
l7YYphbe483i5Ndi4pah4n8fSRHMi71RKvKBI1F7y8Eg0kJ1OL40C7KHP4h8cL2L
dQM9bq5BhMU4T48lNSCuQsqolmFvaiboH6wCB8Z2RhsZgeDT2mGBW6JH9gdDqA9/
hTka3HrBDq91kCrl7W4vvqGvJu4F/kWsxgIJfuLWLwUvZuxPtKZuIbBPIE4NjLh5
2hUH7YpYlt1WR4iDpMxTFEdiCZ8of1UR4lQVbikdyfEQ577xOjIYvX7LHesAcvOn
/+5yLKh8O3F7lkpehwgOww6zNsxDcFzLqUCLC1NhRCpIJF/x0jea3UJZLwtzsDX8
nWhBY3MiJySDadiPdVZThvHMbklJt7/HVS6EfV2VUnbEN1jP/1QKBV14RxQIZ+T0
MioCryZLXjPk8bIkqyOTxslbToqYclmfp1FLbam+DsDtSm6FRZojFa3gm4ruECXe
hRlFVM3Vxcel1mxDmRR5FRqPHVh3ZPPBPjecTQw5pnM8swH2LxUFAE2seKp6WxA9
113WxnpAnTTOllEes/yrLCuVsnbR0d3IBcXaXQaqlK8zeebKDQ3hicGu70Y82w6n
+wUDqWIYC2LuM9sxJHg0g9gc9SIGFZcqcF2HNmq5E8gxVzqRowzpHZTysFX890QI
nEqGJAd7PpwUhPAjnOzoglxtW0NsTN8leIn+UotCFdFat5QWev5FLQ3pkcUNhB1h
2krSH5j4fQcYqhRbLTKdtOQeSgg2e0hlKNp3Kjd2eNm4ImabFPCqqVkBCuOAvqC4
L0wMQFJpgXDsdgFOFFnJvI4xJ+gmIKLyIlAW4gO4AwReadQcAaHVrqSuQ2zvdo6t
v21HkHDUOkaxywyuERWDhddRo+43FgJO+2915ZPX4NhM775VvRZRksIkXaEoTOay
uvWyWyZUcgJ3kCEYlRopibpZBSOvn4Gw4vk+1LtHUWVoCtRZaMQ4o+Fw/IQE26Ed
INAqAY9v2/N/pxC6OLvPZy/KB/1ccueJz4X02XmWgje5iWjbfX/jXPKpeCdvq/4j
J8fBzVOWqtmDcALaa7Vn0Pr4sv29UFhjpiFxiMzxM0bhfob3INatm7oYr733AFap
Smz+EJ1BaieWV/hH2ujEV3Sz73ErpzaR0beSNh0xqiSmiWPBTWVyIlqAtcHm0wip
dAeg32i/YspCI0MEqvFC8Gk1vjV/d+40IYRBZ56Y5DrQ2uo1+1euNGlGZfcDQWmw
0RQQFhg99ugdYtZNe7JymM2I4OpV1Wvjtfbh0lyRt+o+dHWDWb1a52oEs1o73ict
muTuUwsEb3+V/aGjJsVTkNCkVUeF/K/QEl1fc7C3Jcru8BLjo4M0vF/QmssIJx9o
Jl3EUOaGX5w4/q5d0CHFte4SxAUXxfk/A+uhHJYNuuVMpa9eIhDHUmLLDw7WAJyK
zGam5BxwSpTTa9MNIU4qscgwhr9Y8tVEc/dmdaQNew6DXC5EgRVrlUqQVfJD4ZmW
ANhGuSXeYn62UK5VaQHzOiPZLhVs8eo8cEsZoJF3xkim5ZD8GPa2V64UR+s3LAjt
H2iSMyIqPQzQutpg2Km8bD7L5mtZ530666WOgZY7TwJlNZ0JVhLzJeLVj1+KVKR7
vZeAD56W8EeDgAqH+4YYtWnMkmSssXdAtqVrSK88EYase0gkQ6VD+iYp6np0IwTT
zg9jNqllZ5jmp4p/Vam93H69xQJr9JmboZ7l+tQe11O0YmhdIKUiPs1yYrI91anF
yP/Do8gKnJ3hkMHWerouYCXU3HEi5qYecWdlX08D+9potparTh+++VgvsriNl1Qb
/lNYBBs6Kroj7SI3JwWF2Qp03ErK0xTKWjvQYuz7rzRI3x1lHc2biU7+bQww3Kg6
7icKbHIA7hOf6UdHLoJ8LmAgD4+zF4q68dKcoLoDIw3O6lklVmrMl55ladvadTgF
zXBk1V6ewlqJcJvLF+NLNqWPuQlr+Nox8lvys2zR8N6NsrUXlKixZoTCbM1+4SEx
D1T/oW085rof4fnnkN81sXFMpQEMYaCtg87RSlJiK/AfOZ+DsIXJ/ySdwyRhTDSM
+Uz1PVG1fEV3PRHpJ+Oz9nQJKO4/ud6gAqtO0kIfcFspbnjCRoXyUnvfzNn/5/iY
n2gbdb0Ti/njBMhn5jpJjY8YVeusQCPLuOeW+aOIwLVT3e6u6fah+cLiXL2Ka8n6
0QbypghHaz9BYVvMKB0W1qPERcWxvWZmUM79kzKJzcU2mNsToCn5hptHncmFM5kK
pOa/+0kIFJbEYDvfLn9R6/RDSQuHjErDQUd5XyBqTmifvHTRGB8ivha6/rONSSZJ
FD6Jbm5M9E2HHpKtffay6MsYlESVVuSwX2SDGBY52447qJaUW+PEPyASt5DubbyA
9/Wl9bcBrALQRDtn443fant4MXteaFGEd8/yyXZWDnCjDeT0wJwG6HtlWMYkd9+h
M6PMxQdeH02g8JyrcEm7LzvJA0kP1ymJAHGyNk+L9wbZQbdUa65o73KeoF17S29s
n1AkMVl+k0uvs5/r54BjHOLWDZPq3mBQHpjOL9Chn+yYrNuBo5XpBj0kQpos+ZIy
pZBo/tisYb6gEVG4CrwAr7dsNpaNkzZn/ued4siqmDMYgaJT909bwxLfisu+va9r
BFCOD80iVogB7FQNPTqItQD9xHFNgD9IH44QppuCWNzpaOVeeOCdbKg+SqWpsVRP
Xkm5GAqM1odEkOtXMFdX9imjly2S08hHT5Ya8Yu5Bcqvn5Jf2C9aZxqTw4PeRavk
OzSHj0lSy4AKSC+q56Fd+25u446m+L7yX/Wb6VZRWXYs72QUH23fdMIR1+rOqlM0
dtEyxkJ8EY1JtbF4rN/TgIt3R857aYLZxyyBxjCJsy3VP7PeEZeC6yOhYDhp2Hyo
+NT3Pya5zBJw/VC54uEaYJYpedEajnamKaFadVzN9p7vc7Xni8Ba+qz29bx45IZi
sBbbXWNPR59lOWY5S0ydkDhGmX1rmz7FaXXndiNA8lp1H3e57U9yKfjoIv6xES2N
Vnkl/VDCMIKD3W/r03efPdQZ5jk8oU4d0HzZ+Wp1BcS4Cea+qbaPt+tRT/inoqrS
grSvvTPVT/wXW9Du6nm4xoWtXEm/M1MIlCLmTIywtuC0fT+D6NWDBfe42iqEBB5a
/grPVJDSvsgDWegllDo7WyMcctomaW/vFHsSpLSGf3lzPZTpzdbxQnD2EdGJh1z8
FqA1xoFuCOAOf0pxPfEe/pynW4Y6KEINbj+0NFLJKp5kMQNDXuW3OEewwB2jkvY7
fOZLWzTolFnSJqi/wdixdF6mWWv/NCbFyB4qhsHZDi9FW2BQe6RZBZHDx1L9BoMz
9nUN8XmF/7Gtl4r75vJO/ThRAX0TuzE23bIu2+tDUkPPn+DfZM8PeDM2jfsAurC3
kAdopH98izeX4XG9J/0cJh5PSlgJD3vgwdAFFks3G5k/tYs0de+gXNWd9rbrOYgV
Jld7ABCrnW2HLQ/Lje4rPWHTCikc4hgMjHMkby9Zs6kx7bFliTOMxvoRUF4uFiY8
RI71c3Bc8TqfdDskFOM68qSeGgaofwPdFmzW2O8uQYbbtaUUHPHOoOmDUDScPZRw
AhOixtzOyUbFof1kSUl/0HRHIj7QtYZhiWpNbb0eU90UeSeIFIuwCwKHYy5aerFI
Ziepp3XNy+ycvAF0iB4ZKGEKuYJEeYEYCH593Qg0qc3eFthbKlXd1SLjOuychV3C
xnUuqCIg3EhPkM2We5ybDrgptfeE1pQJBX8l7aWP1EP06FlDRFpSS1wSwjvApGD1
qdMJV2QQ8rqOMKaDItxsbSBYDtgk/u6/fHjVnyCszd+FdWyQy8XPEUaJyeelREf5
ZfxLFZHmgw3LllrIUkLKk2DcJJk7CGaMWdWC+0w8HQrbWWzooAFp9DU0ry8R9m/X
czE1IIRYy6O/hx+5ekdumDgbV9rKU6gat6PISwqrmGox8xd/t0dVSOg8emAujPth
jOvHmpxe/rsHH702ITvcA/mPD5+dMbe96SBwz+iluVgoAIJd0mN5uGnAgcsYAVZS
uc0kP9qQqI0TMmcKdGF+i4W+FKxex1mkgsoYUbie0i0RkxzsrRNXBgcAoWG8Ru0D
w6ANFhUJgNV4Q+fsL4fej+v+siz3K0izlYCUP/eOnNAujkeTmA6FsYTAgYsr5nY5
Qj4XyaTIcn9rfb9wOlv6oLgazkgLYHXdlaYGQVV+Td0C7oylIqG5Tvc3Skwmb/fc
YNgrBNq5U9kZrba96B4pAe28yPhpfRe93r+Fw7GVKBj2i3TYocbG/zIr8vCKjJNn
OwLKHz3Iz6IzMPMETgiIIfgO/dckHeFv4pvX87KUkjmAhivevz+qebBn5g2MBJHn
joQYOkltFSQzkM9RhpJxsnAbX3esHS+qTZAjfQ4mCtBH17ebnaJTXEcPpmkA6LpD
Hhn4rSBs9d7MT/UjH0AYl4kNYoKWrxdJS19aAzUECkg/NGs6olR5MtwL61b16ahH
KDFOOIkCLT9CDXxKz9zIegIWTXS69MrtpMH6p4F/epDDQpqaVTqUtpJO4BoUxbbP
1tF/K+fbpoMCKxb1kj/tdnp5qRpTg2bie787ktD3SJHc73JsOhbk8vjC7UYQ0VQD
6yEqRd/gTGPb0E+NZ6vgpgum9j+PtyHulPrVEXNfFMkln/gLVskkagAuujJHe5ab
VQvOF7+aU0ghvvWawdwPnJQazVmvf8M+vPxdFmaopGeKfUbGzKL4yBBDbdIjBrU/
EfsNIah/qFGoJoUsQNmGCcxkzgCoA6AdbdLlN7YdYLCkrYXGkAPU9ZN/AgDmWmhl
4f4/EqMtQsiPzQ98qiEdnAZkT6RSqrBDDHgvvCpEdBFyZuHWZ3NCnfBLhu6cStAx
SK0XHamZjE2s+V8cze8CjGLWB/akzgxNJ6oJeYRYKPi3Nvstd9gc/SFg5aVohCgT
ufSS/CM03Y9zquflnGip5VaO9e1copRTzUEX0OCAC1/g5zsMtFmhMO3SRttcd+KR
L+DvNWNYcnZUgOPca5yWOPIPlm3z9Ll/c4fdE+kc5Tmjq5AWgotxCQo1nxf7xRfp
MFmNhN9/yY454z4zBVSuFcsuI62EUa7bk4wA/kxsRlqMCqZQNIBjXv1HWUlXEJVc
hJCAE8nPMXw4Ail6zCo+bnctN6ndK74YrCwHyir3lNzI1hbai9O4pTtfLl8Z9yGr
PECwmMicd4ss4k40rebDCACV5cxg+UE3YwLiQsxofXrLqEUNomlVpntvl1O6vr1G
du4iHCGjTMCz1gahV8jei6zYj1FtyOiFW5Rtf0H3Udc3dFToPMnjiaybn6xpeufs
I8NwuNLjGe+U6gWe9XmN24TAvL/qd+tHr5Vrg2pl758cvTlt8I8qKwegnDaaAsBR
QSIlswLI4tuAdkgKB+pQx7/xOEcWWp1vUloZw0rfb3xmb66SNziS4MogGBD7J/hS
mb9nosFn1eJyumsbrk3DVBdZyppoIK0cd6GoDUH2Lym1V1T3UpmK0kDJZYl8JuQF
uMp8aQP4HuQl2Kl6x5xv0qinbZUojvsOVd81R3XJj/K2v2e+Fyn7oTseKYAOK/8u
j/WsiSgkjeIyyaYhMoLMqFn/ri2tSi1rjmfK1/bucm0uCGalussyYgz/F7PbjTbT
WpRZBLEl1mOIQ79Nq2y4Kn+GPhD46jIYtsI6nt6T7uuRC0bbwnPKB1HN4SCe14+M
jCJJak3JuuzUmu2Yj3X1IOovOOARpJtxVTFDQWOoX1FXVxIwFUdJmY5MVZRRn1V/
mAPzPHfrViGJTf9afCIu6DtArNjUexKYOD778lR49u9VA05GJf6/aHvPud6LNxzJ
/FfR7nV6WAvcWIhyaRVM/Hh8wiHRbs2ya2YUnzDQIzsNYdEnnACi2kGiFll35x22
5XhztqBYBOt/dLIBoPw6YPUrSHzQ1mR9fj3qhfoh/5X2wgwj5en4n89Qx57pPzyc
vj+vdnF0OL+AYa2i4Foyng5sQ0jVCf4L4FIICCGxf0SAkMwmhDEBTHGWmxJBQMyt
fbkQOXgI/515njAnr/Lu0PgRytfFGA25y45l0Ycv2PkDxEzsO/NMPTpEWfk7xVnq
s6qaB9JsV8aM+2dFr/Pdlr2bvwAFeVGl12UGSOZ3prIFIx5S7qnzVq3wGKQ73GxC
UDIgAmGg5J3xyd8EmdUJahuBVECNvzPrTSV9WWcbf5WweOx7Sx8JGDHiguCFf1Xa
yTKfosAO1KHNM7HBWH0KiLH2kXMxQh/SsMozHq/SKveD4USF81JqS/zFEtLF4N5L
AedKMX4XGnVE1LCDWXo3HuCwdAmPCM/31iCnCJsspYA7ti8pimqnc1W6axFWjvnK
p0geph94Vp9MrU+wiis1jG/e+PAgNp1qJqCgije5l+QTYxZ7TzHqmK8YJgrZrYPx
OWU03sw28BnOHonYxcV5GdavN4XSHeoCn+Xo9FbV2yeT9/3LaYRnQS3gAJN2rnpU
xdf0vvjhQ/qmh8VJo+QhWIo2ZQl8Oz9fHUOwM4+uIItppCPiXU+LYkfhbZpM3p5X
Zho3z45LvnUToO6S1sBb0OjIwuYUUFd8DlNl9TptXhbhXSFIBRphS0h2kAX49i3t
nHxFStBQK8nSQMxxtBydhBkfGXaf/Hsl3QYxtSiXFCXJg2XDhZwcWz3CyHCYtLTD
peEo0fVg6iywW6HCSgkpNDY5xk7VOb84M3OVswJicP4o6TcOwAgP+5iZhQNkojmE
UG/6odQ1hUlSBuj+w1wOOPKt0gEZkqSBusnKwTQUyrDc0u923rHSEQQE96nnURn/
Hz0qWVsDJKmX6lO/v+2nRDp6SLHZQMa/rk3yrw+mnLWNLhNuIK7Cf4+Q7vsO64YT
rj95eNQTsq3iNi67dIFrP3mjGCkPnmRWCUiZBLST3wZjo8IizRyYj6MDe5eLtGeP
GqMH45vgPjHuLwe1mUg22zAH10UP6Zz5vof7kILN/feblCMgT1agMg+g8EYiVmqH
xjIbu84sqOi/zyPqJfyJ5nw5C+uiXOu2UVLkGlUa8n5DjWJNqBDgetO0bSstO/do
pUC9s9dPj+JUtjQ9Q0WLiH8ROzlhDwwv/jckYCK2H1ZoEO+q97ByxeyToMepXxaj
tGhn9pR4ZUW2IrbR5QFckqkfUfqA0Cyua2WEqV0u/8P0no+TYBnHqivaQa3WlQUv
nsjfTsIc/fXm5qiZueJkR+eiebE3xRDVy66lF2mgE7Am+sB/PZZiB0HyEVenh/Oy
rrjJS4gdDEFIZjhGA/8uDNJCxTpklUg4kN8nuOLdSy7ZOPqLvgjBOZFsWK/9WP0q
QmFOfrAaLhq8tcDsDWZLAmh2hGib8GBvdyAUUSNoVxJtHq+iLCemOTYOyz+RLndo
v5dogcm2nTu9DVO70M0qubPd1E+hwWIWxNu4saNvw6fRVzU+fMqnRAlOsUPYv4Rz
nqKmBYCMlOuUeK5q2A2aE5JWUUTl+DtZyjKJYPbEwg2n2W3YCbKV4MjFAnGr/fmW
rP79ADSbXyCx/+7W4VePy0bTiHmAJU6HfuBvOOYAsbsdkzY6ZgtHNOSr1q62KgBz
m2nKmhFGJR2+0sPDUjJWvL0Bk16S0x068TaUsJxikjPrbeCFum2H2l0/COwXRYwR
4yi88RlaYCYsiG4e2kQlbZ9Jl8Lv2LNSFcsVaRmHRyDiZNJ4zwiQj3PKPR5o6d+K
AgU5O8h/8mo3Cr8oQP+cqJNSAE37pcCDZRi+DLYRMmSIh/S8BrHwvmagtyZ0KJYf
lQ6BOqcYGr/fwGwi/W0wLmPrl8OJLOZj5T/eABq5Z9o9/udCrOAkFZuGItybfYSr
I+Wtw6phN/fxJeQWhC36wtX8UwwrDnwkePydUuPSEPF8jQZU5U21pkOkWIfo1DkS
mg2UVE7DuN+2XBqW4pp9NxMg+ugsqkdSHvr+1KR4Lx9kT+TBfT4hWg7a5KSPcvu3
4SnEIXRj5Cx5saWP0kkrnfWgGxVo1H0D/TWLJ/d/sEdAYAtXxJAa5OSFtlrufsSe
YAppIrEHauHV2FhnHKAdbAOlHCtGTd5A+6e7pZEyWstQXua5TwYiipWb0B/w2iag
GB1y8radyt+3N3jFzJvZA6xF85/caj1sKIjYq5g6n4AY+RtUtpb4qvtMgGg475BK
A71ZHgt8lt/InH3rSpE5zr1d8qY0Fgw4zcfFEfIRP0VMDRcjdnlGNBqGdWzb11Zr
17VSnGFc9MlIT4PMeOxdZP6hNCEiivfICFxFJNAaCGVP+BrkFTY7i4zIN/X+8PuP
gfQHbiGHVUXsEfEqRnDSoRP6dRKrhaYmeWXb/jWEuz1DQL2LZPpHCTtQHLr+S1IO
TIy/qPkOR1vIAT6x8CWVeLaVD4SXqGiPvrz5BXi3RMfju5OM5XR9GYhbF6LBtJfd
7K7eABWYjo6g7u7r3K9h9fXqXrXfCo3RUGs5w55id91pPGbVT2txrUMxMi7AkxJ0
0M3C2yfj8wA9rDge7ArtB7VwTBWSmIG7EbERTtmEOXDqlksUWlBfeFsivk51aVVj
GZoMlGxlCl4bgG6fgJcpSpT6jy+z6A1Y7j2Tr3Y/KQMv/oSKOF9Tk+KXW9bkCTjb
M0l0ZWjl5NGxyt3T13Kk9joi/NiamkvRKG35hpppYqOxhyyXF9Js+rTMtBcoey02
b8633sqFWXpzYDDYodSl4hDFN5VYkB+kZx+za1WLpsReLjMoAuTkhy26aoaoE9En
Qy9lR6Vp8x4ZObH3VEZUo2qcq0n1MOrJiZmwBQYCzkHVkwD6jqTS4dVN1L/RJ2oq
znti5u9Z1Z5y9SvF/BVpneEHvGHIBmS3fPU2HRXq/YA8JqMNEOP0ePfLJ1qYiRCH
jM7Kq7CWyHziPnZOwqFZqS14dgLFtqwMGhNigS0GR74GRepwORNocpJ1ExsYjZLS
eFeHHNOXwCsEZvkFoyDGMtFVsl9e4nknevw1kYbLO4CcLSZJ/0bbOB4ygxP+niKE
J2F3z1nddyjOCMNw4OlSc0UJHulOJ6V8DMrXbWi1F5HFjHfhvv4GxhcL8R1+5WJh
OeANt5Qo16nHi3PqKgtEnQUgmOaj/+g7Pi6nlFksLGObmdWGfVM364qon6OwZcw0
vgh2M32uIy8OV/uPRt8rLrBCZvK5vMrXSVAYTXCiZUTd/t5WYCYIk28FCfVAJitd
0aHTs12t2k+FEuzv7PGNEZ71vLcIjOkbuf/vBd8jBjsSMqOoPkfbGhbNcJCqgHCR
Eae/vL/ptdc0vjnA77p/oQy0nQSWEe6e4g8Lktr+TBftsM+RcUWGmB5Hbxqgu4x7
+0T7DyEmfOuHL0q1pR1Aq4ZQw14KNNPmn9Tnj2FBv6Ctyh/t4kUmJOiSijxIUP7X
CMuPRPRrJAM/XkPKv7OHhbr6dPav/5AMQsvZW1e9L61vHFE4LxjcnTicwwCHVnSd
MWSvIaT4oqtYZ2Cmx/0kPmmCAjmbrIT9bAkByhj98xUNbFnFfslzBwpGi6Pf1m+0
PFQUWIDwsGPdbt03mhThLbSgmBAaK9a9iEtYtaTdskKCxSLBj0gCx/PrpPi9aYyg
ILVs9nDr9+PRH9f+t4XXSyAJ49phNSBL41TjqZBCMIJ/su+wARpGzZvXvF5NizcB
w20xDNcqxe+9SJ59CVg00iD3ysRP/jzmGR7+v2wAvA8pQRbpNxA0iyd+66VV+MRO
ZZjDf3D3NNaeP7lNugVXq+zBtsnS/p+IjSLN7D3y3aDWgpwz+op5AInncNte7Et5
7+bM0ckhK4pFiPGTbixZT/GK9jMiy7RWnp/6TR+BhOcGa/VnYE36plvO288/XMBx
yLFrD/EGsxRIu325kloGd7Of7x1lv1/eH0+U+gGsI6iBJtulzJ09p5Cn8l8/O5KJ
P4mFYRrtzz5qm+Mg4RS4+oZX07kplmG1a1W0jPhup/XbXiMgKI3shb1+fkZCIT0c
4jiSTdA2duXYW1gjeWhLesYVldla8fTRc4dEcuiVi8rxsOrFsPf5Bs3UddId7rOL
gfFTzC1zJkQB75QOGFr2yfYp++8X4TqQ1pC/JcWcoqi729g2qDTNPkZb39YbKiYv
aGmPhigngCFPfrdh8iyKjdem0PMvfqj9DwZQDCJCThz/j5JC28Eh6axY+R5zK4OP
EPyzhnc/bD57kwLEnMubT3xjPoEkMTAOY4P+QXO0xgF5pV2e+0qDi8VIUIQogiKx
W9LOLVx6hQCuC+23rS8LwqeuVWfv1ut2+EHlyz5hT/rR24MYZHTwa6RSr2f8Vt5a
hiaVzsGmv9wFlEJH0v1QET1stbM58F80EjMscFI9nwME7xhd5onZ4YTw28tyjXB3
rM+/pw85cbz5KpEyPH80iVuYoOvMJV/5UmDgfRdXYcK+2OBAJTR1UPl4GgVzbXjd
hMAh90OnfTzv4+rKmQ9XL7vV7+gCexAw5g88z0ce6iC/hx5/8dAZZIuUbtwLPaBf
P289pNEEtYnjGHhf3Ab8ym83RH/I7QW+RfwmR9jiIsB6uiqAsaaJ3B2xUlVD9w8N
LSxE2iZnSMb3VOqUfhAazXJZFZAPmpW+8xPtxkS3Ej6UAYPRsxZwc5DNRjr32ukC
QuuPSQLl/mKlY9n+/aYj6P2ZTHlpR2aip9TccsGOv/WNbxKciUdl1W+P6a5O79ne
4r5N6nxc3tCx+Lo7AOLTJxx5+i6DIowJ+B0D12dQs8F4KtyADElrus9rI/2kHZy0
5dTQz1OSSn6KbOQnuxFENL2J5BwNYkdw9a74JGqG6D7/ihciRICP4h6cbTVJZrKL
8bg/hKhDykqNehpK0OUEuTBToxvYI1fYbmDVY/4u5I/COctYB0JuoQBfX1bc+Blv
fzo9SMxicx/ZN6uwGEskHM/vwReRxCUq3fvPWxxYF/lCoUhxZTLDaxLjMktN7DNI
ywZnJMjPv84JIL5AkLnTn+BAGAw4xTH8j3deWfywG47WiQ/uv+CnJqTZqaxXxT7N
BYTHaMgVQ7ktfp8PXNLAyJqMCHVJTp5m+h29rY4WCoi47I355kUKSpoXqQHwm0JP
xLSczHzRtc6aCjPoQnzrIca673uXK6jYE45e7Rw/qVWfzebF6PWXFdye/JB1/zLN
tL6mka1pvdES9R/1Ydw9KXdl8HD/YfGSssCoTIvv84l1v4KdzTR/megLqS5M1pNQ
n6YrLV/RZMSsNpXgmqaFtf5xKowCXWL0w/74EvKbmd74jivDUYISPBLX929gJyWN
9YAzOY6Swb7Gu3Jxq5/XFW0rel+Lc87NG68rg68qChHO8UPJhYdH9ZxUfQO1ANGv
pLYDbKaTi1bqST+H+g2aT/+3YffOyefulYxYk0/gUQNACFzjohk/yfwVe88OPLoM
e+s0A8CgL3negjJctSvDXbiIXzHnHgjIhR20AAS1g+tSYY1wsXfzjaBltsFc+g0a
5KYQh09OJFV67h6wLoPQqnab5qUIHUY+yRznbeDomQZdmu48iPO/61n0Idmpb1MW
Aba8Ke8KRwebLmYLg1XhPTTRoPh2L1bSah1KxDneUNnAdwPqagNg9ubl1J+lzwVd
pUCjsQtDojQWk05696guRHvsIrhu3yRF0mNOD6J36wbmLI9vFrqM0ggo71MBFiKr
An1NdYyk97rUEEv0XhH+W3nBCiC+uEoG8jq2FSz6tk/idk76jMZsnPZg8LF1btL2
I+KS67ZZhImJi8ObeMuaSORMpOWJtr1iG/TM7erICcf3ll+WLq/lNWfoOhciYJO+
AQ+oYUPIssMOYj63I7iQnpek6Q+4cUSfCQbphyyzhipGwm4ldSlHjwvNXz74ko+k
i100oEh0byBrDDrX7car3W7rPYO74sjw5gZuTOYZtVP1Jyta/I0jwjENbXCJet1s
6vM1QqWRbsHOQ4yoGr9szJoHUY7TvhPh9oLxiwisBffQbrfoIUTpKrceorB4lIPT
UEJKKBMfW77Xe1OfzBNYSNBtrZo6GFHg+7mpqtymOmt7X5IJIPjFXxPBIzQi4EP7
kYa5JItowUG4hYop9JX5qt85QZAZDujtMqXnCiM+MRqIinnkZV8K76Jvl8WoVOBx
DakrvuZjzTltsL8Ptde3r3jKn763YzkpdWUZbf3yBiXgxOe7BUZoIhwZHs99dlho
aVHCnJOhEXlaVCkd2PYCcGzaw7WgHN43crz5SQS0RZQ3I1FAi8VBJc5/VXxxZnVl
DzrxFD5MRmSJyXPO3qyPuUSMJO2/Xr4yFlHRpQ+CDd5Q6jYbGPCNDpKsFStSL8tK
TmWdVS949qUqsX9NbO9QdFNdfkbGPFgWPnJNxHyplx/47poX+2jUUo5p+nahVeo0
ot64Po1Ca+N1Www6UvpHeN7infwpleuEY3AOzCsJ7BlIr+IbKVkb38ZhDpKNvnlu
azGHs6WKPUvHqYXRBsgRe/xpiAeugGXdoCDMeRlsASDVWMYpbG8ZlSUm482pgCTT
L5RCauMzzxB3CdznXbo+4Xf4Ykqv6ETtE+NwhRCdB9b9hIoaZV56EPhTnJKakK70
4ZyocIs3hDcs1shYEoKyJiqPJmfreQ6higl4talLKYKnQFLkrzULjqHBAgaBggFo
M4yYC6CGqPKPHBkFkS73GXlH7pNQMjJUnoiAqJEgBhkZKox9FfXM+DeSIvCA0ZFu
pHtSBlhQ+b5zHqB5zfdOATnNdAtwt5RifVcS+9zVfBLseyFQcl1RvhxsOe8VvGM1
EnUaJUA6uChNW3WKJ0ZZmK2AVkulW3FgMkd2DOwGi6lroI9JjZI5BxiJ5XXy6Xqx
AF+unP56Dp9Py+A6OZSN8v9gIbzNq/6HcPI12DTFF47TkNZWpbSYXmZ+OOvwaLhD
vJzt1FoReuy78fSlqHNM5tDAtolrcK4CpHjEQaiXwKD6gobWe9+/61oO+v//pA2Z
BomQrSa7Gzb6sL7CeOLtS+ImU05cNhyf33a8Nhwv6cg3NjDwh+JZxnlWJ+IsVcVj
5KKKvsM4twO02NTCndzc/uZ6HftM30/vVyDK1XxFuC9NCBAAZjXeSEcSVaHWpn0s
GNyKXvMd8JUQVgxFqVRSrLWNM3x4S2jU/L6+aWLwCEA7cQKOKtFzuoYmirV21lZk
`protect end_protected
