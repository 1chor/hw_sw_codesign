-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
0QkmCVyVrr20eFw3xPaz+OfvZjakkEru36zZ8V4F9NAA2CKArgsR/X6BS7KnMQHt
sXKQU+y3CljywqS42iBQYtpgO2q9iG1w0kbSsLi7f+QdFDPtdJBGpA+NCewaRRCn
6ICKriksLHsp3F2Ht2G7fjLmU7YbQN+IeuB22KtR75U=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 45984)
`protect data_block
dSFKbkORgB/VJR8DbWAvG93ySlrdvc3hhn9RC3HS+tbFUpAIw84Ej/P+Azt+Ls4E
D7ez3ac5H3xiG672N7fTsd0pMEW5CaI9NGayfRBNC6Sk+sI+yJU8XGDQREnPSPNC
ak5TK70nsSo3ElLAdAXhAagzc9KvR5hZpBeMsljP7IMVArkYP/o2DDYr7wWlHdVy
uWF/wMf3nGShLIu6b2TkuxwhgscITR0c279O9gcs5zB2/QtSt6Ss9o0/dCeUv8F3
xBV2UqXV/llPfajdnMI/D1rB++7AFaehWaRbpYok0crFusSAXHj31+/K4EvAQF2J
C+iJOayGh8K5mbPQqEb2bGTrjjSco56RRD8kwvxZNDsCSK5gOlEs94t/lno5eIme
8eNqTdmqcpl+QqX3tsdCU6hlUT+XgFjahu/ZxwtlIz+o9Wjis9aEtxiAax6EyfHj
BLEsWMcC7armHEKgHO2SrnJ6Hy5tpTmHzKAJbWhNikAghr+c0jYT4aVHTaXF7cMP
YflHvtg9guVV7Q4+0uzs1eg53nmpnMDHDdkicXk4HXECoIDVq92h9U7aYR+OB151
+R4ws5nosWFPnQOV8LQJ4K8w79rv2WWO+Fm1ywr9/nC8xpSQsa+zer5z+662dvF7
gKc2RiBlkCZ1hqFRR4yb8f6klnDODPJ3KBDePQpMwhKL8hbbKi135ANZEdzwVFun
pWOS95FGYSgpob4fDYcMpiBq4/6ZmyTcor2+bwKQdh4nEsm6D1x6mTUUgmtL0VDE
1HYDDodCBTCWUHp3WgMM2YhD+MLk36BJlGAEUEGd9mK5nSGJMtjToCyG6FjRpCSa
MOJk9RJCcSPbQ95Hfc8wCd0ugO14+H8AwOpw95hz+kGrt2gy8RJLD2tY3GC1SjEO
+xl/f7P+K1Ee6cuu7vE4qiQbOT/gCCYGyAybOdudZuIScDfzYadURevywhHurrJb
rj7UMTCbUuN3ULdvy+xo/ckGlRffaXo6HrbRF69J79Lk+uww770KeLRtAWEOymRA
0fJexeu5aqBnOiHgT32rWHVNIOkDbZOGgI/igWaj/VKXJ3q/xwbxphQE3jTaU5+b
L5PzmATRCNh30xOf2wIoyWbu1HZg6ADBc9SWGLIXEer9zsUa8mlnnTu8m329z2gy
13lLIAaF6YfWZFIKOUaQetTJnpXzv1kCvNXOVXXH+lKxaYXRLSfeLWKrlkrkD/uG
MQYgdfXWmKyl1J55LCrnd/QXOLg1pcL8xyCJZTv3yyiyex+Y1M4pmXLTRlaE0SFm
xZR0EjmKLIceAGFGDtO4L/pBINu+MY/FEZqIYOQCOjsZmiARcVu5FcRO1t4RhEP/
2mm3IPMVVIMEJPGUaX7vdlJOEbr7U+pCMZm9vpMYEglmWqj+Bqk816q1Lzp8cmN+
9PsB9NTFiwYqqbB0n8BF6JNO7SYxwXSqUv4uIDHiiyX490o/6KKB6fZi5mt2L6zj
MEh+OGgb3/lkmtcqmVTLw6rPNKNyj35hK+aRbesOAUR2pvWelSbHvERpBjOL5jVg
yltUi20IgPg0nhLr8Xpgkt9cJ0fv/k0g0gQZHbbf0i97rLqYeM90Ms0FryZQ5S57
zbS+wKSZsUmcKMvXWyyJNnoopAmDGNAnn6sDEQYUgWrdctrEc+Hb/YyCy5fvniQV
6cQ8VKAgN/cSrZWGEa0O9QmEq1eIRt7jNKjCKQ/AAt0Sj+h5ivfjYw4wAES1VEQ1
0zfJ/3k+Yax94/OF6qBXSD6x4yjjQBnf0nYhpzHTw11I6VDCPFn4E2Cy4d+UHGfU
peq4YM1UzKfE+Uv036WZJpYsjxmZPNOo4znNdE+i9VQ8IkGJMSdgBfmZ3bM8UeSR
fIc5qYfnKVfUub0byLAnyMAb3+ws1mgdQjmh2x/cfAxa34UGwwm0/043CzNTDB1H
RgXE/3KOM1sHY/uZz+tyT3fKwTMlDWy6nvQ+M1VvBMZP2JMI1SIRTKGotftd9n5y
17GqiSucANFiK+7JQEcinSihuiIvfAllucBrQI37iGiPL8u27yiYA/4Meg2PLm33
DeDf9xcWmy1Sgweaa54YI+vkPxbetWcCh4cVQ6hRKEvpzbrMcykK1N0WnOaXtPI6
z8ZQN/0VfUkWxN+a7iZphsibgtQHUbAk5WAm3U/gonxZN9h3yRgXUuCeF2HFxjKd
hXWug6tzptAG1+UH6iJRSftApRO0A8famLiS8e1zapZ3cMJuR3HaZdDm/JnJBn3f
rCO/Pqh+IsGN1CddD/SMHiwqpvHvw5uo7DXCq2Y+H0ASSq7Qp3Vsqv3l2MWdO9D2
DWTqcC8PmDj6s4Cd+kGcojppfDJOr3k/whea4h1gwJI7+CKZgsSiJ3QhbR8HH+SC
gmhb/IiCIm4KyYTrVPOVYc03HN2LQMeU3ZTJ6I9AAJnPH/YVA8QOA52PuoruyH1D
9IuUrZ5MdI+0y2+WQQbTJi6BShWZNcYsjazhogtO17cDDqysU4y+VMwE3YhamxFQ
VKClStV7PwXCsWGv7xQHo8QZHcFACzwK6/QL726ykDzcK9/R+LUe9SkS07koqMRl
KpfK/p38dgXDg7g0uucOZU1S+bbHdRirt649LeVLeKPkemf2Hm3UK/ZQt+a5Ta9V
U56jrlcsbYWW5mALwOYCU0vYSK0gYCkw97YsVffQpvtakiTqPbULoXlmw2eUZafl
ztJGJuVc2Ny/EL7Gm7QmWODV20baFN+ZCG3A78Nr+VulXIp48kCgs5wPtI6JWlyD
17AU8x13q2x4PW/RwaPVRjb6x6Gmv2NmzZwnLeXIUHpUXV6Of6GF4QuiHTQy1V4T
ms/2Jd5eJKKsgDOnlMopM//OBjtDVOHFljT2NWeRaDVDbrBNqtUNAGvYSzO5NxxJ
onn8l6M8bgDJZxks7Xmd9/nLdZQ9YwfBgxxHzE2NKQilDgz568XmO5paYxN1Pb+4
uH0LslsnTUsj/xi0D0Ep3sqVFCBQ05q+UfYD5fE0AXLTzyHra/a5E9Ns207rqmlp
rvmNbkpsJWCM8OUYj1nLeRp+qQ77yfmJk0hrjipds4wEGKIfOqqZnms4750lmK8S
B/soWbc3ec0hXOxYOCMSo0u1rFOYEkBhBHK3tt0muJTWz9GZYEoWKRHDuBW8iQIQ
s1n1rylg2thjkH1J1t6LRSxRH8k5+4yHotN6GvMXE2Vb6pddEsWoSY4a1rMr5CfY
wkKSFHI4WzSPpgnzNifLp2KwMs+s0Pw4KYqdIHdG2a6RmqRXDgXBpMmO4mIrVgWN
YEwMjY1Ae3pihC+qGdTg6TCzX/r/FhnklVT66vfF/e7kWSknfa7/ndgfRhBu9AIR
rsRpCDNF7wlEl8px7OYKR+fUMlv1PJbvv+BstdXqWNy+yG50L4XQoW83fPZLpeHH
cOCFVnERONlCduihZJ3MMG/foB2OV7um3DPfcpliWc7/59cQWFKobtZ6tGpvIlga
A078i4boZYb2D+r9vNY6cydUZcYg7esP7WuVxl3EgIV8HtzPUQM2XNXQYElk0Oie
NlQ/hDflYMPnvtH2mzUX/3LJdjQS86zLE768bSbbask/ZUDANnMuNmEwAesw4rDs
rnKpVPT2GOzpHHiKDjOKqIU2A+54Wtzmye1dNufU7yles1IZqSIq0Wi6CgUPer5c
OYB7+BvEal3vDTDgA/UQRRVfbSXMu7eLLHvK9O4rbxv1bxoznQJYTSBXDJdfzPIM
htO0tO27c1mHbqvoHMghLog0NDd74cATJrB2qNlBNO8bCIH9cVyL+xS9LOvKbcPX
7o5ddSFjzmtQDnNTD+9EbM5fxkmz6SVWS1Z7C3g1v2Qvbcdl8lajUtUK/MNF/dBx
yGOkNsFzvPgThISizIXXyOlP0EBtPexccp2fbOy2ewWyzy4CoS6Cn+8GkuEqqDSd
qu0gTMFWCf+0/nOlsL8wY9fKBjgDEpKpRaxcDsrPptaq4XbIEMQnbKe5W3gWk2Sn
IlpfyrfV+xzccQhTtVNWJh66xGeX7OCGZH+hSHnm67+G8wdyv9PU0P/704qrmGzf
IDR1zlVClGDP91gFeVP+hmMlsyOj6gtzbUMjCQ39Nc9eCt6UmMWbptmWSpdk8DDD
Ol/ChqS/4udwhNEBo6iIyQ3nOiSxeYGEryl8kya8pVIwBZF/BF7W8Md0/wO0u5Ig
oBr8K4X5u7T8srreOkXKsOcE3u3E2xEjh/TVOWkou6uUGV6dc4Prh1vTZLZp367I
FOTu+fyI5E40FIvTdzpOQqQ+YPTG64zT/uHsGZNRqXs51R8sR1nuH56XqSIlhcAv
xo9P94DMyalyWP/V9u2sdt8KH1E+tkboVqBaywyzDZmU9IPvUHh9qsKFJJxZb+jX
saRT+ZfhXhuBSEuu8LrY8QKc4gC1E4lx7vwYZhuNQsYfbB9MTEw3E7qwQ7DaEnri
XsYZbmXgo5ewqVZGcQugh5EppzgjB/sFUcSjnL4tidrPsf32yD0J9lU+Pw86y7OT
U+i/GqFUgS4Pom0mBWamjibnQ+RcBLUWnf7BoFB8G+0mIZb0OqZxVLhSmemT7olL
q5xsiiE4AvFhXuGXZhMLz4Dyg/azFHuveTGnHLVNrn2eJxrQxwpGtiPbwzSFmjAj
uIBR4ARSBqGDqbxF2LfTg/qIltPDw6CGQXcuHHipnYVeIxtd+I+dPE98IxjAr9UM
9bJCV69wOn//z5WISc/rVV8ypIKv5jIURVrSTrS89vt7OTVpfoBefs61dvVnGU1v
dL66Hnzcst0s+FOdCoMAve6U4Fs69woLpeje+ZID9Cmpd14tX8BzWPpMgE+sDAv0
5ZSJV+ELbxHHJ569d/ugoJ5UDRa0vC9Kzm0Dem/TOpNmMSIXYGPXpnlslwqdlptw
MQxoQndyerc/ZOQvnGsJklJ4rIjn+HxWHgKpBXXmXswoUesGADV6/nENLdvPtg1q
lsduM6c85dng9raxIKIdcac7zyEObE01VNxpWFZJMkQRPwfiRCbhCaIR60VrIbN4
zib997UOZc3Qs7rGLmWM2h3ez4SAL4FnhrAuGk74dpI5IZUQ+yZdEKoarvj7rLzU
jG1XxBiHk9A3RRILTwZ/NgNy/+dH9M49oZBVy4RQ363exMg/fqrH2EFOaIymM9sY
rtl7yfmJBt1wJ5MOxESHssqsvxcReNwGBlZa3zj0mGrhele3FvgtAtuX0YND/jGN
mB9REF9d1JAHQuDI+XeydmCEU8MYvshbgaiR4nRGykbW1u5hR+hNCt46SY2rITQe
2Xx/sgDEkqffQhvFKbHZvgJKDzu3JP8Oe+vxiN1uDbLQg4XxdzZvScQmGPKCbXrK
gwv1cNIEHfxxqvjHdoPRpuAlck34ZqXEgvc/k2oiFAex+3Sb09dp3aVcu9S6gejc
S4FSD6ziwLYEJbJJ1D2pz6Ae77LPdSgZOccRgpTuoTIfHs/6aojTfMcE2o7tIBjo
e2uhhiJneq4iQlOT3dxwqGYcYmzVZeOqr2Ydg3skkE7w1Gd+flsFO9kSWeEVBNA/
i9MfPCfjI1y2424M9lnCp+q+B3VA2GSf0Z+bPrxuhy265Ayi7HXtDk0ehzVWt5Ij
4H9PZJb9dNBVl3x2gBdJWP3EEvNj1RfhGw3m8T4sTXQKTSg9dukqDncA/feHJyF6
XHZcmw7ZSVKsX87HeDatxpMw6rdXSjdiSOtE3vOaYcixFegrzBjQK3pWz89xBEf7
Out6kFMnk8N9VSCZw+/9lKUTZ0SnVHQLIPPhL/7SyVUvHFnZ1CtYX/oFX7IxYtZE
5UedAYh2QU5iOxH0gSLmdhAelAZRmt0+Q9Lwvw/m00jhO1nofLnPPNwHAYxkhNNy
UnhrOJX/JA4R4YjKVv5JtABmgLiXXE/JgarqtKJtOqE8H+Alk5b3gweI0mMVl/Xq
EGA0pjcvOI+qFGhe3H60UUT9dS/OFxWtqhL6OGLkuXNsLutEFDR8290xQEKRF7d/
BLJJgdvuKhd645WilMqgmkkLqsiEtrEfYn5tisdglMOZVRUlnx7OvzzYcWG4BBjU
nWHvfhM0zhdKK58VypW6FiWAN5LkXuGEvnW+Cb2Ov4s9TwZ+e5UdDtj5IEHLVXkh
2rlVXzKzAcJNI3iuSvCkjwkgKxgXBNHBnDShvxoVafJGs3X1GGry7fqs7NeN6bTh
E1+fQ44SaLTgDdh2aZU6kxcMj8XxoSacLvbfK3pZvNqtiiY5W85aNMTnU3T9CiGE
/TPYcbTlcdP4YEzpc4+Tq++95rw2/JwWy/vxIn30IQRQinuDQqFlYXUe8YN9/lYh
dUC52+CvpjSKd9iWI1/mTJHyMkwf64M9+0KalLvohf2tnsJxcvYkUmsnDVWsAuA9
uYWEP1NLGGZIs+slQKt8HOerWhImwdyfl+4eeAhqNaLGQdTGYPOyiS7Jcl0MhaXa
ZKmddVHub3TuZGb8kbROCqVbnuxtKzO52+Plx30KEWSUF0bf4zaL3JCv3MMPS7L9
ivUL6mIxiDViEHPMSwb0XLjSr2X317nqAi1aESMT4yxSaXKL1PheiC0GlFG1tZ9m
aSUapJMRxyFc+n7Q5rMPrDRnvZgDyCT2Q+O6TEx9yuFp8rklgHDv6d6KTvH1I1ju
dDl1t8Ln5ZiNYpDdQDti50nYZywqVsg1bo2fwxuIFh3+hXkRWsMUtYFeFLvCw3PI
uXaEIjPIdM8nT2MTOBME5h3NB5oZPo8QyHcgbRaxSvxwJSUxHTu7ow4MtJNu1qam
ZOBDrX8CNugZvc0DO8i3t7yAT706R7LRYGa3ECtdXQv0FrkAINiJx3ftyyQN1J5t
nhGJA77Abc+oXWbC5tReSyNq3ni7EwWhLr/pDY0buVzdhilLiK00mx3wvQdsIN3o
b4BDR5d9s2jkNJVacSfaxIm1+1FQzrb+E5rGc3lXdMNTEKWToG5uGlz6jIl8qaSc
wtBmNYD7YWZUFF3lylKLty5jMUDtfq852jl2uwZfQCZwQhyUJmhmheaDSuClueKM
J3mmd+yeCm258gXBXZIEKhAuZZYRQE8WgY3EwYhaQu021eodwqXVKtQ4nPEmDupf
vOdBTZ9f/Nmn8zk27FnMlx5Q+JuyrgWZRAQKm3NK8CzzXKe/eGW83ZMjrY1GcesC
zNU+KzHSujEFZ6wsMFw7fx0+eNRMHjeay8RTytFHWdJFkHvGOhbWYYCzh6XzJCFa
R2nBmNVZCpXOgo973sjLhUpbV++A8WT/MS1NvqaIqtR9Y3yErSGeOOUHg4fDmBgD
NCfE8udwGd5UXGbXab41YokSqELjRiwqajHpUCxlKP8qMkYUHO17YR658CCOlMP9
Ul7l3ahIdzaez/lLBRTTvYkkLRRlaFhC4C8QSYo4+Z+Ey92am2c8lHcuOXZ4I01b
j++ihzzh6Lv+wsHAZ6xkKa0LJ/Egs4T+DJUxd+I1To1BW36MRjGea5wBKYih6YNI
xyVVAsNjRY8PX5O+vS5SRkGX/Z+6ZfLyV4ZIv9dMESlkd6RysO2CcycHnb0qrzam
twb8BTMK0ffq73O+L7R+fCY7uM1BYefgo4MiNNvWzu+EI5HJJY5z4ZPizXWHdPIF
G0ofyemQ85xvxRnZcWkZsuTjOlkKmiaSUfmqwQnAoUdJurzZsctZDO012Q0Q5yYn
w6sqGwSBS9r4oz/DZ1+zLZ5+zsQMqtY1tkcFBaK4CnHRHB2GGC0V9WFIvexBTolp
RRHb0PLUjbqiZLVKrx4iIt9R5CRKMDfysbE9VtNCLgbwwjSYMoCPKpRu+8JFw8CZ
ZTi8AF+FZ6ep4TZY2MevDd4WAch0bQEXZAjhEpvwtHgvJMAx/Uug8vgA511r2gGf
G7uTeMWMhe637Dg2CZjUth1prmZUHl6tQIzO+tConHj9mFOjDZrftgNjtWli+W76
RTyyTg72aoVROLdV0mLM/PFFD6f5R4Ko3IUyAtUBnA4tXYUuCAqxZ5BuB+7HyYj+
HSudIio9psdWJdMkzR56DFFcTxkDkNaXIzJbSzwgdGsDmt0zxGZG/5YcKJbMuF9w
r8mBivJ8m27IS0eCcuC/NTQLV4EwNXDuOeQN0wYqCFrGb4u1gnxwowNzRtIuYBPI
KyakmsOlyG9OidMRI3ksXvFz6e9w7ks3ro+pHjkQtmT0WAlwiLqhl2DwAzbMWAVt
8bSTrsiZDIDr7KshUUjU2ME7VklBM7552wrxPuxXtrlzE6JPnDrrHTiGIXa7B364
PdXOCKJNS2E+qQeeufhLygi4EfYqqSNdBoRy/K6jrJHN7r21ZgKxJFuLzBryG36q
gxJLcbWah1uj95N37V7CLtUb0LYkLTDzvcFjYQJoDqe30icwvVJ5ObuXoiXgfGIF
82hMB7oofq4supVDVD8MErGor64hjIx3EPOVDWouLNlJlph63fCsXf0+NyDe3Hme
wmM+GKRz0q7687YISMraLKEsphlXB3EXlkXxH0mAnByiDDdpLXdwmucJMrlYe+SD
8dEOhkWceusR3ozTRr8GOJZDrRjiJajs1J0zvmdqPsozr+owT7Zox5wbGJoeLF6V
tUFsXxfnoZGVUzlehY2eTVKaNK0N0vsLyF4r+m8iMIpRyUbQihZxjEe68JXrePwc
FKn9pYWSiCpWfbQacrIRCIig9uV3HgHR3yRcrQGftr4ZWxkcst5+0LnCj5y5HzxZ
ltVnPp7eg9p/HlWmzWim4D/UlA59zn8zxESsV1yrwAD0o77c2/ciA8FDZCQJHIWt
hmNPhCQy0zJEt0mlUzOdHmZPEWVESh802B1NEJKmHA7yQ5K2XlHywdIP+YIEQXxR
Tp0U+QTOj3hapK4FEXauv+qD1Di+va7flc82E4pjwZU6Hx6CPSPU1cAb0jsGjDGt
CzqjXgpfFfVTgPsFVik0rSGkfKb0MKfVNRXh6XYtQA5nsuFxLMXBXjkkpvkJm54G
EVNWA0S0gL5kW0Gu+0ppZFKsOhinWW1I2+2KbMTrWOMCGm3p6mm4OwgaUnlgmhAu
wukE1D8Fduto/5La+zsM9RKrTxmj+JkbLnLjth9Sjfbqy0IiFBDD8OlVTekXYvkz
WhM2OJCmFGqXp7N20a+aGdmwV9ZzNqZ0KiImeoUpxE96lMbq2PhYkyiWizjOLKvF
acO2H4HcesLRQj5+IgkmJEzv5gfOnZFLFJSSv4GUN3HdyrWwRHROBNKaFBqR5Wwy
r8QB6b0qDF0S9k1/MRdsPsMqq103L7CtoAvFgs9yyjcs84PB3srmTjf9mQS7DghD
ZWg0CKVKZ4z6K0fewvtVhJR3TgqM8MljbikGAqc5ES/FxYbpcDAWaqbZ8HyrOcuH
jOagUloBzz9KQIgoE9x0Bj2XkO/VP6CjFtJDU8AL3mvmgu58S6YYAv7IlaobJvpM
lJtF2F7sJp+BXtILGaR+581sNSQMJXjBpaZelzxN5P0AxkNT9GahyTD6c9FNsIGu
GcxqfTrC0Rt91sKGnUaiJiIRJ/0aeieUNW36zxdyhxkTXyZKY49yHlRJ3IrF3rQU
q3OI+tmLocCHfmvMPJmbg0OnHLoQWzfk1Lmls4QBo+QT7TvAMW1QsLLRfLIFmLz4
HdweK8r+24pgscOlaLc5EJRMSTyYTcN+8DhA8Y4tW+t8QkQ0dhwnTgp3A0Z1Gm/C
vYPIKnFMIlYIMnkErcKHc6Tdncl81Ijy0wpdm0eneHPFVDjxM/QzSkJinueu/pYT
GgWraz4HR4etlkoFVx4VB4w1KWSgv2YvkV8zr4k7n009D0pWO5j/AWKIlD2OrjdN
c8Ql9c72PtJV3z+xBuJaD05Huo+nM5lOSXtBnBmJksaD/wCx0qV1JvMPkaKvgogf
MO5O/cfvy1cTqkYZY40CdQVQBS5HgxXR49ju6NgarW4hkFpzlCDrxX0wC93qWGkX
7volDO0870h9ERdRpu3u1mWc38LgRuWY5hZ+mOLJY9uRXCu9/071St2rpVzU8MK+
6sq7HZ/SOKBdDUZmBBjBvlP8tU91D5jyg5dDuNPe1frlyZiW6AfoU9p58/+Nj0p+
FUAoQqj9CMubND53qBPDo2CEGcSizIiNu2ITGpH7YnhpKFphbqZ+IawbQeQ/rPfx
ovMTdexL8ag/dtWvDpbrasbSXbC21Zt1SH00qfyg1prpSVQVJ8Dn4tWBlym7qt9H
Pn969IMgkdnYQTFDfuGIOLmTg0TQzKTgXu0TnpXxPqnXqQ5dTEQgx+KjyKyI7Dj6
bxZgUwAJvLE5zRJ4q1DfzxQbihmWvDLPRJgv/Z1BFmpfWVyPq8pAMt2fU7XzVivh
iUwdc2qNRlbfCaZR+opHowg9hWpO6hAvUaPCFxDzvl44+8qirBF0CH1K8RhCCtHU
A3g9rrIdy1FAT5jmRMFpm6phBwIIcPt3ndHaMUs/VtVYXndVCFqC3yEc1qoOxCRM
0RMTwTgjrmAFcZLeDHVa9F/dDJTCMnaBb3UFidsW34veEeIwSxiPlUkVM/BpaE7w
M1+/b2tBGPuu8QrQDFtJ7VQ3qR92/VGmhqz9WgZp0yFzWYGf/nMFVTbWZo7WlM9Q
Vr54jmUbf3cc7Qe2DxrT8OZKWTkxnCKugByj0zMPf/5U44BFmxQzZ9Cnu1np8wci
BfX/NQfkUUqTkqlsd25fjoHxxiHt69ddtjhLr6//ER/BJ1fYFPVaIRmMWZpmOP3T
OjNlIdq2MgLaEwzWVgIDIX28YxwuSphyenqiNaZApMJsQ0mGoooamGCQY4Hiqk9Z
mq4RFcjj/yxfRoLKYyekBM/p2SiTO6/PLLGp3Rw24hrURuhPdkcM5BRyG8WLMvjZ
5EiBVzMu3kc8BBRda0eM+CQW1MY/t3B97G6XCjSZd/OP/giAGV8G/wtqNlFbHEvn
XGTNCZWY3WZlKsA4tJQ5qvM4j4X8Kuf0RmTmCZ0kNy5q4aW2Hm98sg75StZA9bUZ
bxR6rhImiWJGH3pdlDNzmofDTVsVcOyvoxO/lAaaCtf1XPt7E9hCYU3I1uyhD6/U
0gTn58QOxc1uT4IRRBbCL9/p7NcfXYy+5lhlHs1EXMDshfYPfmK3kcV3GjvP83iH
OjOf0+8OMDVyveeTn39QwyZjSIXF01WLREk1/jZ0iIMm+eKHswhll9lNJ2TNkc/+
PdfbVGMOZFqlRbllNcMalC7n8C5sBTvJPOiCnFfMulFsoQoT+/5/MzPbuKtFzprG
Dn29afMwiYPLu4yaoSSGUxFhIZiies0WZrPi6vTjElQNcRBV6YMrE+v4UGpvOvHl
L8+faxjdTP1ZTciE3WfEmY4D1XTP6CxgQWsHbAA0NI0wlvnhtkvJo/jAwdtHU/Nz
UEkKIr0UonuV80mZjArZamkpyaG0peY3l8yuSy3aZtPkkaDTe35daPWPdIpGa1IN
URdLfA8P0yZHMgB+vqgJqDn6W/agNOgeBTTPd+vuvQGrSQvs3ZzTLMiJnuE5E1sf
6g2CkhIYiZAGmHVFHOnZd20B0h6tlfoV9CYvbGGp9dVKsFVnnZM45goEF9/BOAxf
IslLTJbAt0gmwMx/V5oLV5yk/nBThQ1IMUd0/zcY0T0xZCu/5DOvms+JwQlE67k6
RtvriSSt5MBExa85S5/POXVbpDMTFXv9S1lkdwozClz5fEzTu1B5pQl3knuqNiZh
ci+cFATxGjR6ZI3ZvNUjZpUqakgQ3/wnKHV5Y1OPeUUQoR7DZa3DReisXlFgxqr5
vrUxouapmG28tm/qI+lkuyks2A49gjxSwffc+iJktgzMk5LkYp1zkiWtpPz7AebK
9ytisRJoFt3PzB0z/COALLCDsWHxPdv55Mo8FD4v3eU1PDLohoYB4f2zJuYlLoSZ
IdEXEEp9s4Z6saGxyWhItE7sOK0CGyYr+xFlJbJXLON5O/hABJqeAsn6EDW3auOl
v1WvGavgQCZRVL39jkPie59LJ+3WSREY6QUmzX5Zy8o6HUErwPXNU51cUc3wc0YG
s2+wuq4XcJv9J0t3MHoIAm8u3qTDn938xgEZMh3gbk0cmN1Zxj//899vp+AxWQoj
TlFDV45pYmhasiKjd4ygYISpeYy842wGwqwZpyZdgkf1IDfCumutL1XyPqGTQUpl
wV3137r62OF6hcrC5uqNtZ7w1LDgHQRz8oZi9a+iciBSecJNMAiLWj+xwXpTr3ID
AS5c/wClCK51Uah44Ci97FE9X70O3B0S9mRCz0P9RAcOBfHF1nMyDG+iScO5debM
58eehkF1dSyF1B1Pzb2y2y1Z+IG43f6tvd1NEoCnqlNH7p3sx3nyCLaTZrvTera6
NFSkh2eJNVblnHLmt3/DaPxXn/7ojbh1NMq9rrKQdrAWCNCQZXJOdz3hfAZsh2vw
722hmDyCvwdhfcYsbN5sv1Sj9SiZZgyUnteJmSkAT4uKXgHUkhPy5ynJzMw1LYLO
OykYH870Ago0fbCg3g8EiLyCjRTkWhUGkENWFu58PtLQSc4+kqTrpTV33Qchx6iC
Iil7ZTqTJwcyXSZlnPeMc5CNT6+h1bcxzchhUM5wjYIylEQrNjFsdZi2qipohc0v
ua4Z8sPSbt5RHT7/whBaGhtSLLBedUpsAQkqfyIngOxpybMJeyczrASQ9WLJCTs1
nbBmyJ9x4gvl/csoYJ3w7uPXgSApif2/NsZslluQpAhQrEKGoz+ywsCYNTFmWIE8
w6C9RG5hzK1QWz38poXY6RXHqPkTjPStLK5aO9lLK/Bfkrn0W7HWM9JaRRDGA/x5
Is2SYNaK/53h0F3oNOuEjBiIvYXMpsnqS3pqYAaRfeQBsnOh8PTP994zJLJNfe21
B1WWuej37dfwrv/IjozNz0UL7h0kYTDo2v3BlIXUFGXlFyzymhxwUo2ok6xp+Wry
MU62Fbabd0RXq5Cosr0MpZj6wdRUD2vel9Gro6XYl3Jz+MXmieElMbaMa6HuQgtA
vBVwlY8dH4Ev6TNmc+2OpIDP/F66wbl5QWmb3RK8afcKFdllnlaB129FzmzfLpBX
22TYp1WyT+oh+VRARZH/Jh/cCX1S2COMcS9chhPgyCc1pqvfZBKfk06mORKOd91D
yCJY6+TfxJB5aA9rrFB/V7+rSOh9JByyy69WFfewLd6AnnUEzpjZtJzGyxQeQ3hm
+INFyMFTUQYcKO4oSoYoMLdRED5dTV8/bIJyL5uRoG5WGM+PwUtl5ClylXagRMB7
jkvywxKKL0lvPdbqsZLWepyXUMOHAUbXIu+jkxrOycBiHIbsXNXHaA2WvxIuR+Mw
DvO74muPXv+QGlq3F7vqY0JR0cAEOn74+p0tLT7/LHSnQoi637Z77SG1uaHy6K2V
gUPfdkWBCkQ4sCiybcV+9ATTdQhr8vn7iT1dN4WqLrtz7FoZWhrAnYWQ/EuUhcO0
cOHAsDVWk1pcK2fFZ0E2iDByLiff2e22SxtBBbTfGLG5/Xqn2yBullS0d8xbCPw3
IKRuXs9N2IJP3pAOPMwGT05wmmDYLS0dYHwY4J1iGsg1Il7GUkB1zRsrzwTkpuRb
/FNqhte8M3mOSsu8PyxAmkclXHTEfevThVh0l/zl1rauZ6Rm+bx3ezMNSVvpuoBG
EIAflLPkpPvDD2w9SDZEWkDMcc4MQWKaH8bxHhiZ2BXLjqvju+11AzGMHgDiQnAF
h+XhaWRZlE7Q0szQL7335PzROUwvYyXcLFg2Nt+kgpsFMZDBYxQSpGk+hQm+k8na
NXGB4JJgAtsveJ3eQSXYf9FP2vIuubmDZ9qxfh7Fctx4Kj+hYDM2yM+QCL2PdflK
4nG5vEF2QTYO8ZKGZ1wEjGpUtmMo5mzmcN2bXXCUJ2+6HUXVOOV0OiyaWgIgZUj5
hjB/RHRDDrIYIQTME6lHcSM5aoKoPQkHK65BiMqcFR+cM2W6UErjVBC9m9Tlqsbo
eJe3hcKVh7vkbZUWWmf64GPXIT8ZE+zS4gPlO5JoKvxoQSt4zPcuBUuNX2c9pZrH
g3WF2GTD4ukMuasGiOXq1PbpLTTDnV6ulPHb7uf7qUV2K/ulUV0z26/EywaVH/bI
Ka2D/VPUu20ohy/bWuFYQfi19m6I9LkIlCWz6zXZDRRC50+nxiskkAPY/rfvCza2
7be/LEiQGylULG51LwGtaOIQUDZgCrwF5jnrouiQoA/H9vnTfeNHv+m7fNKyz6Ta
FExri79MIF9XY+VFcJakGzcMPCg+1e99QNfheTNY1FDwac60jjVBIHGAU1M6OTVN
cX6XmoW06xgicYrOakNnrpiVc5VhcuwnfpG7Lm/iEbdWKbdzF/jSvjkKN4ArVZ5E
gwJhP7pHjTJBqJ7btV+yGPp+xawMEB2vwf0GetzUxCEnxeGaF1SEqmYkBysjR7z/
YBYdyWbvgF4PjDfbfKeD5Ob07wx7wNx3iyWxwNrc6mppjy4kJJya8ekX4BBo40Mp
pZy373+iz/oGT8dOD9YD17cdfQydMF8zJXJcUWYMAizXH2U7ojIcIQoOxaG60jsR
uNBY5fT9qYnDupWVY4kMLnNrVdjBrTUrryz0V74BnIBPDFxUhY1CAG7fPO2VUF9q
ybIlgD/qYdP6ulWQZQBbGXo5gTctRUeP7jjKki3YGlopW2n/n43iFySYUlu9KXJ7
L45aaTIp+pLp8SXryuQ9U58CWRZDRqRJZRRu+AkDiI/3MoItkGbzbyMCEtf+b4Q4
zxlwGDfE50yLoguMW/aKsm5qwRT+aIbzTvxT7MgfpabdryG0XwQmoT9oijQvOR1f
l/dlg0+0mY/jIV90kT+qJOphDedKcUi0rfe1qyEQCXba/atTy50ISVttdRbjEE6j
vNIzQQdZfQ3a9863ZxU8DSvCzGVT9LezfiH9FFDnM2HiJkOfwgVtdKgS7B0VrePF
Q7+IlgJ98oGLsYYOGofJnPutZ+XPmEP127lfrhTzDqdehl1oJvaMo45c/jWbZNos
aqubrry1vddQUUjj7w7/zv3MZL/B84p+0FZ9h8G9GRQmbtKtb+WAbhaGA9lxlP5g
DYyurPRlTZgjF1u5YjnMyfz8TgxgUGgopKWqfGBiCTXR8QrtANjVRphlw2NLldlS
+Mukw5u150Ch1JiGe1gHtKhe1+Lri2i0WLu6ePi5otLJr4LPAej3OUidGhE9ExRW
ved5rWIbxy/XXiUNqHPG6i1F0zFVMlbfNcAyLD9XC8lncWRbnH/8fwEWu0z3ghLc
+WW/glLRnvXUGR4vCk+wGSDt8g1ay7kBgX61tuq2WXBPniqpOK6cwbpQOazmgHBK
kwpl8S1Uj2PMT0RMocILob1RQzZrJBiGtZdmfLbq3aoyheyERNexPuqgLJ3Dt+NG
0gUuit6kVDypgJXI944U8nhTbhbWWfgz6aSKVUCl1vXhAtYWFTYpFrVMiDW/1Kg7
KuAYkciQxq6I6UKYQ2wq4Y6KZSyKP/YEySoO6nvjUqN4ul6G47sDUh+KSuCzx57k
Js3amJHN7YNcgGjfvibCm5MyeDDen9sDoExEXHB8IisDcjBX6OAm/Y55/K70JxYV
fDAnA8UgHoAy6uCfGjNnWwe5lOU6u/J2G6jIwMw7qQZUDiXJDwRblML2FV7eDgC8
vjXtBAl7HGxgVnTOqmq4bMXZAli9zycHFmTFU72KLsRq1W56RMxqkga2tykJuUqe
EpTwKfHX0a9mR7KpTDPt1JQW6pR0FabIpzS891RfxQMZFKj7Jkrp5Ip5UzHDEbEO
J3Ff5+4I4fD7GdW76/jb9rE5qC6DN6rl4ovv3uqntwgigkwGWvec5Zx/e90DEHid
wYI62NjIW8Q/EG4gdfp6CpQu9WNT76vjD/fN2HXCZ6WdXeaBxPw1yJ8TD8T/+ii5
h88KMvGC2hq7xYG8JjFnHrtMfuxEiJf6ctzCMTIpdD+3atlf/tOkR6LWFZyGeq30
fF91UCca07Wyx3G1AM8VpwqWsiCgZtZqEBlZFoTu9RMjhPPgSwfnYa90KDrRp0EY
rzRNSWm+VkmkhmEWk+a5sJio5hfqgKmlqMJ189N5eou/JQU0VqBMz6d1j1DKuITV
eyP/zbk0fdqIm0DYEC7AZcauXzWOPktvmsQg4MOX5KUqPlic24PibcWcgRNkieoi
ZE4jGukDOfVO3G6h0X6hpxRuSanbOBpxZ2hR2Zya2w1ZsFR6C28gdkgLB+GnOGbR
JpgY4z0YxsfFUfWB87IEG876DzBJNL8Tkfe2SQm879laSG08nfFEJQPS2dwayOWy
7yUaj0wRuF37A03ZQ5OTKF3/mAn22yozJnqze6pwjlzGadQdy8j2WUSjL0Ti6A2j
bcmRe2Jnn4GQKbPqaXjpKHvDZGuujkNys4ciwW4YHSQ/PdjiFeuREwYtkUpWkOWZ
u68epRh4Gl9rx+m/DsBTX9Zl96S6hWqHxiIFac5Zb1NJzTWVQehBenVrPY3VRcb1
b4ivB9+CRWCI33rb+yHeuIMPh0X+0UmmfSQTHuZVqGmadhdOHrKAnGXOgyDqewGE
MAHJX5hpdDa0njARk3+WNjjpt0aqPeJVOgQzvEXXiL0nejEB1Ax61VZaLIaUt2+R
0SSth9lBdYbJOCFfP0o9TZYIvHPET0GagMWH/tIYR/3yY8sGqAWnqdDIFc4uR/N6
8jTP+upMAyoaYJPLfqv+oTkfMGLpeEc1j/9wQkOHY/P4ziZWGi/sOdr1h4EGT7zg
dN0dDbvAeJuS2aD9kmruSiayN/9zG+6a+Cz7E9nzIhfFcWflx6DbAFNAxBM1hdKr
foZ+hMRwZ8bwg67pQQSLVcqvcMg6Dgmr8moso2u0jnyfw6vCQUOFjRQ90AtUUqbb
fr3hBard2WlHXriFkarM08ul+FJAsjlaeV9U02qgmW+NcYyiVEpOPkE3IdDkQ9QZ
pHddzFumktyhCl6rZD86mrv+G/VYrL4vTFzb5fICgyZAxLG+i5nweB9UKVLJZEco
OOCsOYnyrYPvFAb7/b/Nf4o+aHHsn75HNba/i1lVhwP8xu5TItbCgGJ9nM3leMKI
TgHBSXzPd4+V2FwEcmpqhYVZT7exG9JpdY0Hk/JNOSjdiPkrE+xYjFtRn9MWtJNV
wF6XgM42SDjqCVi+GkeEXv7MKMFyeMsikHYG1Ql0tQN2Wz5Ix43tLxTWrWTrlmGK
9VeYt/3G0gc7cFeDd4KKpPAb8XqFgshWgnCam3CVP97yqW0KzRGALDMpJwHtG7FI
eGvxJKUkapI3M3JPE2BIK2x6Cf9te9FCrriGWaI/Dx9/FiBopOHCRkhlJQF9ZqVi
IyIT5wvaavm3XWXWXraYEpCclFCsPq3RLNj27lfVB+FJQrOVPEbA2cj5u6fDWYUo
bI73RsYDULNprLSZRm/ckWffbAkeTVBqLaeA/WOSm6Ql4MEOdJVfPTzpzpgN29ko
xCio4EYCOdPMEhRruhkdsaNjlSq6MMM1Y0AO9zb9CtDUP/+U1b/GkPGGiA/JaTMD
FEnR1ODkQ37dnt4ydHXrkfXCqCk01XNRUERGtsx0iB842AMtNDSYL5e1EC0IKcDl
JOSkbAPG1xzw+DCD4EAiCwlrLVjw/tBxAOq9/U7TCA8a2kQm8ZGqZPNSl61ryfZR
Ua3bQfizKntooRndHtge1YwQqB5oM6IKYUqv4YTFBWmO4+Vj2xldUdOlPe9tMY++
1Pj8y6zH+s+9DxHuOORyEBl3a4GbcEIyS+EJ12D9EgqhJTM4/95zDGCdsqEO7eix
AyPDKiGyW/orO3mgtLYLqWo4fXAFMYyBWVyukX5/bfKQCe71/1mO4RNZ2J5vOdgu
T/k8tqcSkRGnwI8HtybR3945MwcHGkXv4Xajp6xv9ou9bTv8laW2pa7zn5RRBd2L
gHEsYJn+W4ombnS5yBu/PeNa4Qw2zf9z5Xip4KctxCE6If4eqD5yPyTyt01hk2+k
XZqcKN5+wCDSmTcDF0VrO5gMjXyIpIxXm46ZOfNgA2t/aW5dJhaPYYQuppgNCFnU
rfOPjb4U+dPM0BL65oqawPO/zya+hOeLWwmtJ2AwVKh7yF6UaNkFVNN66G8+bJ9u
Wk4HiqqCte7+KE3dytAASbcYpg7GA/gwhhOl9Xx+cnJEjtdh6oDmnKAZA7qsT+F0
8qdZ8B2DsInXLsISYUSQAGgoEAt/pPV+rB2CoDTdULmmZazRuTKIe3B0ofYWmoRs
zQXXRDJY46SfvoiIfqEwB+QNf5Je98YVP5EYl6sGYiNMbt/Boq0kq2XxbF17vWWI
/d4dDrrqSy4ZFo8mB1dR9qMyXkMk44a8N4TGmP6CkMISfPj9OB+0674vhxKBmdoj
bZa6aKPu1jh4iQqNa4fObZkcYKkHWZEw2JdxagyTAuiAjYloRzjaGBPbcnWOmS9e
/rGHQX8it72q0adQDk0W/OZO3JmpluqWLXbek50NejJnkQS9cawbOgPnqVNI7cfH
0Hhkx4eAXBBUt0ML48PWVSIrY2ZlaEk5Xmi+1Avt+8WGoSedey1ithupWDnvYicR
NeAlBTaOhwK0xuG3nmL/iRHcevUrOgfGqgLMNw5FkgRABMHksCQNww3w343pvgl4
jWjx5yA624Tw9megNyG+gtXGEeFa0vTVH5d9ET/vBKWRL12b+Hyh6dviMYTFA4Ev
vcABHIpUSsHuGynHirSY4+ftLHXFU++ubpZ5OERIjFip37Y/xiKmZc7iIouzYFnK
FxVByj+OvOjlvsULU8lWePY484g/xlsdbf1PIP+6DWyNkaIyF0m5o2+9Auhsz3Mm
WL6kjHhdm167oZ5/HclL6fPoXnmNCivO5oMFf7ORLXPnHJY+jzL614Mpwfg3XV09
ApDKORgfTLW6nklG6L5MVR313S96K6L6cZTC62qBHEfrJW+AXs5KC9Q3jFw6GFb0
92tsbP+x97ydc0a0PqtCPMkhj5QsUwTP0BMZFSsMzHqlGDWwZnudEoMGJNu+G8f8
VT7yYqfW49zdMN6L9zrvJbmLGyNJp9WLbyeNUxdEKXUhOJAUJL39/g97rPx7B8zq
lLzCCEQ33sSYd0qhxs3HLgdROJ3kkvqoScU1nNV/6F3d2T2O6013lrIunnIpVMRD
nnI5eUkIV2BQMi0I/JMwgPYNWkEpOvej+UGEHPZhvtspjIOFuQvNQyk1C5IVm5mk
Wjvc5xyu6wa/d8sG25sZIGWllsk0sAXCRkHJsaNJykFOdrW6vStvE2+1e7ya38hC
k2xf5DnlU+DkkiC822ApJGQlZONrrheiktyKGDXdfCP1q6nIsbDrmaIKX/aNPZDb
58QMgGwE7do6C9joBo3eRp+6a7plzzm/VzmujBArR0fDuVz1HXHrzDWktqp7Uwo0
BNgjsLCVyeCig6+JoNfbIiua00LX2AzghMtNfFXoLGDEMzNC320g8586YFX543sx
ahrP8hJvNTkbzr/9wxnj2yVjJACRsiTUwmd737euzIOsv35G742edo8jn3dQLLK6
gQ/5RpHPrL0TyOCov+CNP+veozQ3Vmzrmfm0mgCx5QyDVigRKuv/59rykY1brQ1e
5DLIjqexu7/jfq1PKHgTxpYS0pK0c6qDRgqqkllPb1cvmoyS7Bfu50fXSr4osRSG
fT5Ip25gVx0ZxSLrx1v11vmzAZCJm/AUWuq6dSrNuoVd1izTw5eYa0CSu+i0fdYa
FS3iA53cwnZmsKzcGlM1+4qKjMnKC3Nu9vigeIkMZdW1V5QpXOCSn0vmIYzRyyO6
7h1JHIjCcpoDx8fT7TiqvxuzSNbEHdxa6YpqwnnhjKSI7mht0iM0K7C9zqEHLkAM
FgSaZsTFpQRpz3Jod2K98aT9AjZuIJzAe3rVajjVhnMn8Sjay1iRton0ysORGtij
VTorC37ydFK+zZQgiU4D5VRKgYPJXFf7y9pw0htmkJEe5DOzNok/Ak/H8vf30gsD
/tSw/20Ss0A9GztYqvLPgaB4l2PqAHAnPF7sjcXR9BV/hIqHdKMWGomv0GzCh/34
wlT6nATE5K1jNFGXZF0J8Ow+lJqm7DkpdDgOfONF1UsZlJLhz6vJYJf9BzCuPua3
H7IefUFjLjuT1LbsnA59euiFaJuXpyjXq+8BwX3LGl0/ruuM/oybgFlvs1L1yael
r0Scd+zVcYVUbHjILkjgLArnnmdKF4ga3giiQgELnOk/YA3/NU6eNXU4d3G3BxLS
y1i8R2vruQ+3vammt8cTnQZ4WYq2j3UuXahc2OPGQWsz6DXWqxlAiGgSVyUoAEzM
/c3ONaSHQRuS85kaHNNAe4GU0Nl0QaA0yQQP6oHRYpgP3lXaYPwJzhdUsPxR2Ko2
+ZDQJdbMMm7u4XMbKFvtnZdPeopd5wsGgnVbAn0dvqsQWjFW9WNdFHw3Z3+cS0R/
jPia8YYkOCz6ILmvORReBFmRC6t0an47JMgLDqkhAu4agFD0zUuiQldvy3FVoG87
awRAkg1h3lMDXSs9SM/UZpE2qFa9nISj5ZHNWkTYl916gtyKsHNZh+KHyGJYxEvY
KBgOcZ+hN0clHPuzBtbk1HYeH6V2Y8iHCsG6BgbHavnVwr9zCiCxGQ+gW6NJrMj7
v5PCMVVQi21FpeZfaE+bzQukVC/jKtoVotRVOTTBNRkC3dRHhhJOJOBO+Zjg+Xrq
AJX7iN36k8aQV69pIjeIb9mi+nqJFexqff4EoyRS7O+0NvMzmesjD1BmgGEytpMk
k0aNwBiZyOt2ndu5JlGIW2EUCCNmBPGryquvz5ST5Nd1qxvAtqx818KMRCWFwgs2
qv/ss7lZi33MkBp9V25AmrpEQStARWxbMaxXYPKdYEmoS3USKaMFDy1BDan9j2qK
ON8xKfA7K5hQYsNjMJ/3DdV4A1Eubgx6bJ+5fDEhuS9Uo3RlIK126n+G2/76NJbH
WIVAbtyjjM9iEiC/N7Fj68SSmNXZ7d4b0P+WVtgLEz1QV/+1mZbjMkBiDQooV8fh
UDgWB/gN4Fnge4vHcDqL5PCRLeB1Y/GIMziiEVgH3uXsnXRYSeJLIX2PFajcXAVD
JsvOioKK5Gi6w+AcmZetqKnBwVQ/gmKlSHhjTNjiA+fz0eogIs6FXx2F415xL4zk
JfZsc30QMkLCrXrnnMuserIVswbW7ZKMc+Uou+doUZGrR9jnsp3hGy2EbTDr2MUj
d9hWimAxh+xjWLpgccReT22Py8Ghd5YknL6KC7UFedaUFsefo/omuiWcZ+4Yu6lZ
20UkW/eogFOVrzVT2Ajnztyscn+oQXQqKlIVD2NQBQYwSYSrMfjmLwLZOCp0OPNv
ROI46QIWZyrQpoVo0miZz5pYDkv/mOpdxwtv94jvMe2Nr53c3YbVnuLfcLZHu/Eo
wOtTVHoWr9t1m7zqKDNGBezK3PkePtfKUq+LUqrOyNpifA/de833NAw+PYgh3Noo
KI7b02oLf+CvRmAgQY7XkDbJd1SQW17zzpq7pcCzYxWEcpbmDAx2LE5ARBFT3+YD
/JtSI9YwFVoWG7FBUhG6A6tDFcHKvCpeugMIPblXHtQJUAZ6hKI/sGL+/Pd33I0S
hUMMM28wmBiHMnE2LrRe997fAFkZgLq63EChnR146M/aDyiNNQjrRPzfg51aB4/8
60WMRQ8tkwyp1xwKl9forQCXh+wDfjTxLVIPk2t0NJisYJOiAFZfp8bwfVusceKx
HWELh2/JVj+REU6e/Fwhzg+lem+WM2VT9qKNaGjcejuqQ8qrPNulDYYAmPYDRGJ5
pvwgdYbtQZq2702tNOjZ1IOU4SXY1z8s06XHG99udw68IR4KOUDcZEP99KGVFdfz
oxFX5RpWYsgajjuPD8hwQ8UN4rHXCaFjs9b1Zy7SfF3tqj4r9fPsd4P7rS9VWtMB
NXDmSeHw5ydfZNmCe74znO4NMXrYxp+onOLW7ZEcI4O0zBSI9rRoCSpMxjOsNlCA
gx85ftHnu8VK6oDpEd0ibsf/ZWSIPN/6t7UcO9/Xax/EZfEHrl8sGoZkXUgxm0MF
luaDwNhddf11uhIgQ+Z7whjnfEJ1R4lssyLQOH0dslDkhev//6C/tYZyyo9arlCp
nuTYBwB5g4vwMIquRPMyTddekTDrs0LnwRaxecPoi8CVWwZglyEmKLw+ytkH/7Ux
BQhQMDJmbafygrDOCZCjjVDkzS8sXHpqSfLEJi7o0L/c5DSG43ktvlyBB2QamFr+
IoeQDPDskqJb2blOySbIUwIY6buoQwIOBW04+OpVNJOAt/g9MZ+tjb+APGI6iVWk
7JbRPZfk077d16XNTaqC0LkRPlxurHrQHJDYyODlP9502V9cfP8fibT3WrX7X55E
HOaTH7JrRwgt7qtdQXmFIQU9qG2PMEI6JZbjUCTyDNhmGH/JbPL7lcLkq1HMs4NF
5uZDxdfPyAum4p9Kb8SOi27u/Lc99eDc9ctaIl9COhQH96Txwy4wzO6snBhXKO8p
19DQOZTkDVfxTc5KwE2k1wZ9dXyhaLE/qgP8/kPO0mkmrM2VF52Zy6HqFL08eB4i
QGT3Rquf3U8USG/HSCaauM8N9x9lPqQbjO9opTAIXXiMmUYS6f68/n/9dsDh9z23
LEuOQnw2AHTuVtqi9djtiOuTevN947OjrkJeNe1Vo13YFJvwiuw7yJ/9G7xpbQwr
2iECUpjncaWrfe0z+MHPjMLny/SYVsqutmprpQc29BHl+s0K7OJ6/rv+JjJIgR0S
u9aUg2QUqNEPiJwIyGOBj6Blj8JS6AHJfUpJ+0iW4MrmqYNCOrxOA2/4Ii9WBe99
k9Clnec8n/TD4UHdO0itwsjuBy+yLR6p+l+Uj48euDPPOiJfXC77BrW/yyZdBMMz
90Surb3Udb5Nz10j5mqnOll3ShLXkl0+Eg0gsi7dlga9hI37H8B8nN/QQ8C42mrp
S0XNRCgMxnmS1h+dcy1WfFNYqn2vWNK4oej10XC6lkZNMymWpZOng5D5XzyIRy+X
hwRgMJy0SpjS0NppAcIYdcpKxDPIql3Iix6JhPjSF7CC4zJqD7kr928wWADvqdKi
q3lD7XnQ+zBBA39xh3vi7OQQtUYoEPAvdEyEefwt8H0ZhykF2FjfZcEgsE4OuzC3
2pgmP7zJ2rV1jN0/I6NBa60wuHSItnh2qvjeh21p359nTrDlIjln3OzE/WUaaELp
HgDPg3UxJOOwPxfgkqfA2dBO3UTt84cwuWV89Djm8MEWvqllCB/ZrFQypluKaREi
HHx6Jdm3awm+b846RBlZmQC3oCqzItZGhMbhXNPi6oVNQ15sp538utMb4f2Qxfmy
XZvEKsIu6obf3BACj+DcsnBzgpbx7gtwoK9u/0pmEgd3jlnN6BqTYW2vwOt6CnvR
gNRiFAcZPzSzXS3j63Q4ePaa1Kyh4hfGDtYPAwV+Ok/OiXnf4roTzhgwZEpT/Jyp
n4ZidFPG+K6PFj4jiVKUvPgqwjdbqC6ETS5D2ygnjMmdciTUDuHKQYcnDWhfZqqt
A3bU7H29Au9JA7A7tjHjLyzmcSry8r8sfrwOriEZ2MLkIFYE3yPJ+C4uM22TLiBU
zcSgwVHX/jeM6O9XWxsNAYKDaVV82sv+BDYFrlwX4EHNW43OiAzu+v/ntsC6OaeZ
4FkUWL5KPgzh28tV0elRcUQ/nScUYXNC36904F+/GFP4QL8HVsbAeiTSRxAxx5bW
61LQE6Fx9cbPAnu1Pe+4OpDfiDoXNjFqbs5xJw4VADE6N0ZWNHVWWOw1CI2erbG2
qkMMdIgDncsRSgjbeHpwcaMW+EJ8FWWla6iGPc6jqsiJ+/W0wUQzwmAkTS0ylu63
R6tV8t+fir1XurXU3OAgfItzSrBa7v/gQBfBNRuns5Oy2zO/zXJ0b7i6glLzvVkU
5AC1Z42Fe8XJD0VsFfOk1rDDbT1AicfvO1rP3xqyPZAaQPtyNdy17fUSgfx7S1SY
mkwxE1budBOQeQpEjPBC6soh/Zm8T1VhkSKw4ci9zxMDqVt0YE/PTAjRRxOyYrGL
menu/PNjNYy8wCXnMsbi9bYBtI8/k+C25fYjm/jvnKqeIv/ZHz2QnGD7ksg1G/Ks
4GgUJ6+Fusmig/qKKx855HPQ3xyjcH1T9NbNlu9ieIqLEgBafB1VL/z40fy26vM6
bSnCJUccP1zDDJ1T/l5XopqQzUpBRUmvv9cjrIZHf9/KI2PMeH5QgCxScfzLuS76
3nJvxkGjfjTSClzBhz1ZVD3BGtwFrw1/R25ARf5GN3yiwAbXdsmvIMB0MabeVD8S
ARt49FWPsi0Hqz09OZJ0IwT4dnWeY0rlq/MMrVROK9k85XPj/BUDRN//8xaTlC57
0wtT7X+JhQF7Ca3WxtSLFHYbvzh4FfFrcGfhzQk3cdRi8Ux3rJq45meTut+LWMSL
8CwEN5v28ToAqdskp0O+Ru3IvGulmuxBY/FgqFscXWGXJLjjKI/pBYxmIBt7LeY9
Xh3P0qyzCJye7v0C359eENU2eoyJ7NUBsyVGtUUVYprHyZd3Q0RRecmRRd1Y9le/
2ad72OPsKH1fXjkf4sww0Fc10GljIvq1/HBJjF/zV7aDcK/ALYKwRXoyfX2eGR/M
e+9AR3JeUspnp3CwH4u5GVyPVr92NhNM74YkIYiJUFVXgLHlEw2bhkARUE5PM2VZ
7CZs3KOgR5z+cCtcTG4Ty/fmJ84tv05dDmmtySjEVUOcrC9qM+GjXHFEIYMa5ZGR
aI3wIu+WUOkriQwJoobGBuwE1sMtDBZWYAIyBY075Hp3ccLnfYARmk50tce8Y0yc
Ib2h11knMrY/FHeabJcBgQesRtwDwnIZDuKtwK4IBnptzO04+CM7I/45XTVWnCde
bybar3K2+O/PW0ItjZaNH2vjQjLcSamtdB9VrvXMAqVdykGl4TwEImqjPj1o8J89
+tuO4uR89rp5Xxz3Vk9j/3JOlOMlVwX8af40nFkB2DCE2ryLpoQRgt9Lmu1x4212
UjTh5KWaxxALd92mWWS2U9Lf6TIadcFfqYrcNKS8q93XalRMwJ7WnFTOpPUNXOr6
ZUo3qpHyO5LHnULm3FPfN33AYEvoqS0TzCwwitdBdeiAE3fRuH16buO/n/N+7TuL
yXVMLak0yR4Ec/nTHU37nzdON0CbwgRh59lXWZp6Xx6gCqgM+1r/T5CtT2zWyeFp
dy2Y2f/Zak8JrUgCBO/b8IA6Mh+VRCtIG7+FBvwssJZHxF/qz3et+/EqZq6RRSkk
zywPnQtUruidRA33bkLGzZz6rHA7TELiFysu7gLe27ouWJL3+NsNYvOfQz/cLzMW
+k4Kpq42n3XqqgFW9JKggNwubay38keOOOMxTtXL2ULSbrVjM1BFfNWVPeGDyP6i
zvdcFN5Sg2MxZh+5s3ZoLt25FMwVjjWo6cI7syeLtGtx3VBh+IkfUoJSDLGV+J4Z
Nqo61lKGu070CdBNy75CqMcxp+2VTIax7Sp3v6VVZesNVE2G+2x5i0yPnece+jYP
Qar/xXod3e+GjbSbETiZqSLWDOw+vPsxd+FyviblGJxRMZ90uhtsMAWjWvxs5pYZ
yiEABu5xBNMKOc2sWOFkEgEyEZeww4tE7R/0siWgTVrtPbwmjZSiwomi4E7nThWV
52F7r2vxwOR41tzNgjpRfhqEag6CKRALWDbcC+oE7NaH4YJVv7Om66Y0bW68QQt1
WEmNmddDkeC528+PeaaGJRQLxflFBvq5r2GWc00SpXYCnP1GDaPykuitMakJKVZE
fwNvj0MPZdXcZEN7GT0l2xiY5repE/eHk8W1rMhNyOGpR9nFOuOdmfpGdBRKO3BQ
fvAtFAsHJ5cy02jHjr8dPqv2gt0X/LFBp+8ngbeHr2JJUkNGioMqdb4LHYuKG7Gj
+c0euLsl8SHvV7Spn7qLKViYA4CFUe/I2ai6N2DX0/ksgitcy1I5N+ZFx6C+sLsj
AchQ3pQw3jC3KA2bdmcI577FN24NtFYN0TcIsS3KCgFbSy+ZoNX1e7buXdw6sJ65
wZIaCqf0sty2xQY5GviOAErtPiSY35qHisZY+ToG8j0YSMaEB3/6BLyp7P0vwtRu
Txvp4FKFVSqOXpOlmQfkMGszRRyow8g6UbMdOKm5807ZEV1gEEZrVpj0lq5aRYZb
6JebcwQ4zaUXn03IXwdi9lxxq/iQBqUE+CeADjNXRS5DxIViPGkd5dcrBCJ4ZEH8
PxGNZnzm3WM37t8PDSCcY9DS+2bueuuEQ/opIr0zLCi6ogkLuVYWtWDyErnABZj5
3vwSKod9iAgCBCpS/pTe60eclQT/988TzfVpEAzthCdfqhCyjhF+9c23/Hp4uqK9
21f+1Qomogma6ScWBOMf28w98IzF4BzRyZ7W6BRZfViZ83qmrC3vMjbNb8yzimtj
mmX6zic2eH1DAYzbxo3nxh4YddVfWz0OS0jwZoL3a9SN3aFrV88agDQSt4gezTdT
/D67RXazbVAB2llyDgiYvlLMnylgd9YRHcczDTNOeZXLXcuqMXBMl2zuMNnnCjJs
32KxlOx2dSsBFca6x8WEkHUx1iE62tt9IC00rXUDyuV/uc+ZHb+Eue0B6k7xZPk/
qny2y/A9MbdiiIdyb6npBxdZhdZpTwZ3FUl27V7c7DtfbazWJJTPzPdj/w+LeiBR
Ax4MVcGdGZRojOljv6X4DPsLqw5vmLaSmfJvLGirdb03b0D9Z6HSIaGPT59ohmfb
ijmlPq9jMemFcXMZ7U8m4MpqKyH+1bXROWShpHBJwRw28EPl/cmk8lvRqCSHD6Y3
4XhbxAaGHh/9pl80Ld1axzMdprno4OKP5WI/TtsbJ+nk80Ek8RhAyE7FGPS4NSiZ
FkGnkTbMtEFMopaEesy8P1uCprVEE/f/37Vdfk4XwflNn95UIBMO/pv96N8BPyZq
1h9Tm6xIXc2tJuY0rx/ir0duDWwg+C2T9lS+jNP0LpIt83R3s3r1JJLWz7eSnyeU
AIWvE17FoLj/9UrMrv3FUF/Q476l/pttXDCosprkvsHZndzseGULSVf/Y7smrAfi
v+Uh69fzwKijmYOZkAgd2mmp6WyGkLClTfeBqRUmAb22RTdeP13H71qCrZyNurSh
4/QV/7VN8AcUan8Wl0RNWoh4BjcEbhjfcbyWJLZNQcG0/pKMHgMROQktJpzJsG37
66pN2B+5xAlMW9Xpjvl0oGlVSpmvSMSAlN5D65v9nSpF1FpCdNxHfaiqEkibLKPA
DoIvr1cuvKaE/JGkH0rQgnaA+yv0Hu716wV04p5b6XRvvdbNJPaHPysVX2/pbiuT
w1yi+6ucOIBmisFTivzL4VvVIIqwUyZdT15pQ0+vVyGvjI0hmp/SSa0BNu9l3Q04
8UgXUx37GgC4NfdTEUdQIupy/9dDx8cw7Y1D8mZE1waN+ZyKwUSNAVqbJIMO8dgF
9LY1oxEG95Hq5kDH97iUk4DwhVY4s3FXKgSsfoamD5HBgZSbRzqO5qFxDfzJDDwS
6AR5C5z8ZVLA9h4zlGRyfVyI9NJmzX9yTF0K9ZuzuWvHYM1rtM/GPC9jluRMr55P
M0Ru65uuvbglzyWO0RR5FC3GWhsGekg1it58bEiUi07H4JmuW1dz5BpbGQ61DaDs
8AM0ZEIDlNb/+wR4+ctCjz7GuBgoDQHq3K9CGwh1gIFRVaL/aFZdDz9vZuI6Mx8F
IcicqCGrt3zUTNkB6olPXR9rgYfzWweR2cz9OoCzi7y32YCY5It1QKhXTTP85f7c
A1g7GS1jaf7xuZk7hJ71U/oB2+Q4Q1r4o+nkRgnaYsyoDwzCRv4B0wrfWswU1Aij
sn4rb+/NTrPSTAaD9GBhqn4REQcNpZNq2ijQy/UXZq6MCmvspzLu2gLQQ8qXd3p8
4SbxKkUILlXMYKt9sTZhdyFToSJWhXdHTVON9j9SYQfoUUiBuMKxUngW1cjvI2hL
QpLI1TFbqrxaFwTFo/2GhPPyH2HA8vghRi+GID9m4/k+kGHnpAOjzXmw1f6qPKmT
Wl97MAfmj6/txu7KefiLoAGw9cGFOrRsqAjwHvgalO1tWncwWtIahJU1Rc1aYvY7
7UuXl1GCIvgpJVwHUT+TrU/LgOqkUQuSgk9wt7L52eFLXSN+KsA0gz0ThVplxyYx
+//RlbPSl6Il+Xsrj1lxO1SMbrty9k9FBxIdUAsnphgXFDrQOK68/ET0u9aaH6nI
OHkgJHbKtoSOE6UrQ1TwHVlQjoD0NJsp1Rnbu46cz1qY8I+M1V77xyHgpPfVLXRc
EaoLOxdiRKJqJtdCd9Drz8+J8+QVXuF5gDgLMmw4yD/8uzvbE08oEYXXpPIUk0BT
p/z6CzBKbMGgwim/rlTwTWM0EFfOvVWvYuUF1ZQWIp0RFpNaDepiZuh/kBDBsTRZ
lSDf8BMPBrLMC3bGrGcBMsBg1Of4BO6nWXn0KKjA6ya/YBPCzHGFF9Cm/UEHNx4G
wuAcwoWJnmPxQ5i5wdl7L0Qr+0VY8qxxvxtGdh6heF6UJYN+6lS9hTQeFtReqUC/
5LGRcc2cagZSsiMB1PGRD0Z7Ebqklxx2JAB8VPMppMNQQGfV5fJhbRJRaV1tYxXb
VTymiOpOez9nj3OKgCeAATea43nr2nSG3KZXcwwqxJY72qD45vGCHE0sNELpG8j8
a25en7g8ye855WwrPJof7lBh0U9sTN8Z8zt/GuuAEZH5uR3j4iOzX7gS1LxWpOe/
adlWxtmiSeq28cCva5eLEpGodwBEdv3lq495uHIZUOYj67NUHDzXhV/tWWNakZhY
GixNERCH/TrO2W49ktECwKEJlSixS6DFo0ZdjDBKXXkNw+Oq0AENMUN+DjP20fQP
y9cjpR5ENyiBPr/axPNgO6hURUYgQDZ6Dod6CK8gs6GP33KwceXqTlm4mwjOadyL
53Bn0AzZgg6joP4snX1CYJd6XZoXv7nSL4kSa3Tv8dpHddyrTP/02yQ0oqKmYm12
YD33SYCMiqviBm4dP8F3DkLGekncTHNmEu1eJdfY/dC17YXKCa7L2kkhd3m/lEj+
e/dRqDlIvng2DeuqIb5l6OVVumOXNkVx+LNhb6oH2ZFr29O6PVwfMKsJrJ8vSYQV
4BcYwQpn+Y4YqmQ8hYkzjUcQ8DwCo8on2HyyAnIdsOLFM7CTEGS2Ja8OaT/cfAiy
0cbLuSCRICMgbBKlNvti0y15V5QdlzlYCcqJ8X+KnpKi6Uto1QAvkgQ2tsT+PdPs
r5OOcRcRCLOdA71hB1wmSvZk60zYBiSCKRa0eIfpi2++i6K6m7DmeUyckyLTxjbg
qt42tZ0shnZrSAwQeFCxHC66086+l5xFXJCD4HSTqQx19PH5ENX48M8nhECEa+tO
bHmBoo2OE1DOqXf5Dss3wwYmuRiYkS2FzlE6MN889SfRoaJevO03htfKxlcGb/qb
DRLUbm4hZtw1Nu+NX91B+OtB0XB7CdBJ7twpnjVkgBPQbUtkPcOds89JHBZizfDt
AgNESXrsXXfS9M/FiDxb/dvatEBi6Au1/2vKO+Nwt0OqO3OzSCVWHX7i3k5mg/EF
1U/YZw2Z/yOZ+/Umco2S8Qsl3MdwMxFOeOEfGJk5HKxpXYu0/1SjqSsix8au5zyC
sGV/TLhpz1KFLqWRhjjVKXs4Cg3gfMDhDLBlKuslcKkHt/nT7HxnDB81Akmdt9BG
hgCvak76mRFmrH/qfisiNFUu1F3NRUECKJW23apXYtL54VqSiZTfDTuMv2DQXbOS
QaEYa0qIFcmFxkriHPcRNGwGjXdY+tOnn0g0kRbJtXnm/U5G56y4rQ+VLmXkqUdB
bzoM505Ckyf6n9a67HLzS98ObbDWNqf4T9ZqvVQm/h9qRkHsrgwAK6rvQvZeEzcG
UBQ2djqnVZk9hYPXcTlZPN+x76KqCxGEElQ5VvYfgJReB2A68bksvrZy3amBxxyO
mzFaK3s6WB2Gt2iwIiG3wSWfcVI/dHh2JTh2soA8rVabwigozYF6zFcSbZAyGw6N
XEvIpfp4LjM91IdJoE8dU757Qa7wkNYLA99zRjR5vvzs3yjKDFlkXGpCpeYZ+pzk
sjjQgYY0Gs5QBdYltN6GacUQk55iRTVMyvaNBXdXJj9Tu2Sswl4xMilJICHLmmYe
P8U5iLAG+4sAA/KhJOtFWAuhWxuv2kEdRmYEXhS7Ez/FuOSbt3E1jt56Fw+VrrwN
fePLCmPRBXUuOtUN9GuANRG+uxwdTb9nh9kDl3aFCBhofukgBnjiOr7bUWJP/2Cu
/7fbDGGUNnY5V9NuOo2HVDbCNDLXAH9qumUJINuIlYFHVVbzJ0eP4c++vv85dk8H
Doc5bSBrYC29nK46ZEN6qKrGVApyArYNySIrVj6AAS8xhGTWPZehOBx0FFfTpfWh
Ln68QEHrCmf1Z0sMlw/7ah4vzd8Q7qBQgPfM7XCX/C5ZCz6N0fDpxtIg+vtQE93N
623n6fRwQSPZ20CDFJjDv3rGFA/vVIOSJlckqcGb1uPb1XWuQRXGamBbajo7LZbg
70uExAmAHg6frnUW4GMtF52Bk4dsIY9PZODjxBJL8/iST4w1jqPPc1ARaAJ53grT
a1+mCgKuj8lsaJJ3ZOph9Mc72MzgAfYLiVJ1/YpUp3PD36aI+k38vPqC/ba2CUEC
l3qHlnNH9QYgcBDlrww6xQ9orFz54k+5cHqNyt94GtrH578kC4N33TJKhW+jGNXO
On0S9K7/6bGazYfTvUcPVsFIHzLODHYgfBUqwuxc3vp7IIwAPNoqROmDqcHe+9zB
ruTS3Ca4WYfIaNUfKQE+2//Oo/qki4dfjTpWDA4Zo9jaklJWeayE1mAqsmbCAPUB
+E7nu6jWf7ywWhIgzO6w3GyMj9QIRobs2kMmWvmHBZ5iOl9/weDDqQsy6mmX8c0x
g2eeZSxKS7xf6EQKP0M9hUQ1slScKqB+icD2gqIB6hDyvOznFNc/Al3rLtU9yAWT
kE1AKu3AX94xvdCG6oAwq3kIfHSSO1XoWSh8WWB3jHE9JM8vA50aNHmIh6PdCzQg
+9AT/LoNyzQlwlzwarn++i+mQOyd0VqfQGzXNv2Kaw2qs8torHW6LChehu2cAFHF
pnCkIYAkJxbODLN66Wck5rMEoiaxytHzLHHp5QTLDsmTqt/KZ/0Qqv7RMFfKEyuK
f5VocKXKP5iwWNhw+n8lAvZ0YQXmJdsOPnZnRl5jBUsFJVqBoG9cjzd/XTv37VPc
IFWSORv/BmXdUhcBx7cmCkXm3X6DgaCZUaYv6MJfT5pdDM/7CQfQu1lNyO/iwoVu
4eMN43v6jojg/w3CM1k9/qYq77tpfNfMW88YD89uC0I7KXt9O+KwahCM5xf4ViJs
JbF9ZUZSxW2avq9lri9c/2qbb9PfbNUvRs0DNOr6yFS6drCLWWDzj0aaYV5NpcOp
91bP9oQwPGm8hJiCFInk2RXR++AZvSAYejHvE+RoeYyF8VR2C1JnBZCl9oqIAqhC
c6sbRyyWpWwHdU/7GWi6jnRwFu9kdWNbhmV0VicrrR4NMWuj6sVVb+arZwe49KNZ
FeAw+QJ4L9KB0zvmHJ8QJXW7kqYrdRRNkUDc9HTGawWLAt9/RjwSkg+Xtm5I1DFJ
Tf2Kh0/VVP7OtHDoHe7EzagsZmCHv/J6WC4lV5wngpyGgZjDE/NPukqL4kOekd+T
NLG9/dGeteOgcX2KicFiA9D7IBFzv4ZjnMxB2uy74gtkjdjaRYcnWfHSrlcZkfQj
JTdww32b49d7ZbKOS0OYCAiXTzJgL4xpAaNroU/Injpov5OJa7EheSVTjr1d8DkC
LLs5hHFfkhLJrtqF8xTi7ylH/cBbM4pQz5ZkEej0sslo+7i0gaROZ8uVEKNK4qxt
JbZLZ3PSIPXzwGlnFOZ3aWt/O3hpdhtadb1tmHmH5i5mxQqWOGW6XRdUDYPOB2UW
nczwhSVAbgPCzWQkbXjk5SG//zXAUlBPgigqoM5cl3g/b1YNfN2zlSW56vX7lZ1c
wg5XJKjGmEV1ozko3vHCLuFAZ+JUt61/leoDnlFcWZHHqZ9xXAmXOVBD6j5kooIk
DkEE05TtZCCr8cfPcskmdXXIYvjdB8jR7p3u3OvbjqbH2Z8gdi2xPKPaUMZkgMXk
BOFiSCCstT1YJmVIOF/qxi+v72gdhCfUCr76qsFgSZOgyjUttGrAD9b4fuWdndAO
FCNOvH49kliIO5dKMJDjz+nwlJjXKnafHNIyJn1tsRaaWZeL4bc+zjRuV1bjk5Tf
nL3J0ASfo4PqyUAKNhsNf65nSTgtkH/e960asXjLtfpK4lru6d/Fh4CyIiAdKZP6
tPQJ//XL0VVgb76fXAV+77M+KuSuY45n+ZR1LO8VeYpsd2fRyIpC4ucy2l8goo8Y
21J8It3pMtrUUJJTZy5b3flZC4PR4KU5psumjebeYwr93EAfzSYj32+7fLnHw/+O
AF1MID2HjRr91MiByyGuY1XvPAEr9gdJvCMstv9kXIdiuKT1Qp9+uY8fiv0uHA61
Z41K6c/UnBAgKAvwRjT50El/ArP+dVN/K/scDQ8kWtW+PNyuGX/CFL+eGTBqgc8U
GW6V6qnooM+fcUT4jfmXoNZbLLkF1GX2IDTCVHW5vEkPNGXTTT9uBW0m45BdaoLX
uNVOzWIxFMTuB8cUCkheiCke+Nq8GyxWyTQNWlUw+PN3mVSQDPi/3l+tXazYnP+T
65IkNVOPo+UpZYn0UEvkad6rfNfm3w8jjWt5sUDs8sQtBeeDgqrSJGkKdAIxfuso
xQCZfQlL8limtcMbBa5ZzFFxNoZ5FnIEA91fVRmzTXYVpp7u2OtZPSURRhLf7D+k
VdfsekB34Y1l5HCcWG7p5dAySvXo74Zb/o0e8DeK6/r8bCaIOX/wsBTQxjd0RloG
nhF4lEXVkBU0FIAYvvAVRGu+kZDxVmIFJbCpWUESU0hzzhA9TP5/0ZUhR8N1SIv5
lFmdR4VkjcJDM7vvcdrDefSo0gt7FdGuoXIyhyTnJ67owxcoYHI7HSJgf6RiY6f8
V6qv7ija0ioQ1EbL2nm1H/xkJDQCzOkVjLYUlBc3idI1hNi5KhJflhPgYlPe3xI/
p6uPiqYpWSWNIgib0zEeU/Becv6oU2cnyTjTaUA/PrbmsKndEVLVI/d6E1ETnuZy
eOFGPSlSZHdRDP9mRk8X6NK02gp0YQneF/U0sPvuQ4emtRQwpBYFXs61ob4Z7CNE
Chck06V+5vjjlPaqb2lOP/kBHqVA+WyFRxPRk9pKVlv6NtifNLR8b5rFXrc6Yerj
gyLTrfbT5Z0jNHFA2avVbRSG4qaKkAp1n72UfAEEaIykapcZ5q+mdp5D2goNIrFe
vjicvkV4Kv2kiHEH5FUuwC9xyPst3Yq+/yfKO4OF0dpcbxPvflXxj9Q6TrxKFt/z
rI2F0uoNepROR5QyVGaHyb3pZJan1KIWKmC9RXb1gukdYwENWghbPAwih6YHZmtz
C8yfYdb0T4f1+9KbPy01ToU6r0BDE8FJj/i6R/+TCuFLcMKQqrtWvOtZddMmQXvc
pgn4HiBSQZ/fzhmwpKNJAtD3/A/+XRpEC7/v+94bgL1neCxiAOgPT9J0FpbgUNJS
0rjD+GZpNjZjBoFC6cVbzWsOgVujrFYcUu/eWPT4ly+DSgnq2QO+e/zLE/WCMemd
06mhsgVh5LdljZ0E6Cb1l3i4j27xG48GAiJ2qKmK5JyCUiGH5yO8HJr2fnMV4P5Z
2f3mjsmOahR7E19/jI8IH8YOfp9Ehj4c1g+5DWeCGG5GtKLaQXF/V4jHvBaADtUH
kr7LHOaCbPW80gTDrkVKdtbkCiBbzI0Qpi0x3cllN/sLyardwux/KXVp/500nA11
+Mlu1YttX3w+xitSfSk5+/+99icvebqZEgOMGbasUhYm6IlzExErsyK/9G0akI+Q
37Y4OezI9sLC3vdf0fqAB9flBpG7zhgs+80a9g1AFunXcrnIDq2IEOGqRtN48y16
uWZnvuo8E7jb9bBa1AF/3lhmrnL/zb/pzUwaZGDrWAyX7zoQVIEoU1Wt6PA/cQW2
kYHiEhSbDUO3cIXfi/sJqUdRa/C4sxO4w+P9fseTedqkEdrR3vIZ4owJ7249C5rv
UaH8HI4eBfXRH7zWlFkS15utUX5+opGWk+BUtZ1/ZP5GqvUnykbJz/TD8CGeYEsA
bzVuYl3tujFQrq+2i9iaBcFqD/P/r8vFY1bFPIddkBpQIFsMz1RM5g/KcwMlFe/I
ohOd1E3LB+FPNJecNYpxVL+ZaxaFvHEy9/QAaPUhkyBiEoWJzkKhqQsuZt4aQRny
e8aq5HY8V2TPzAeim6slQXWE9/6kUhPEiBEgK6JQhdKIcTooz8xEHZXQuyCo/bFu
r1Ri0Tf1PrnwLEtKYy9P2m/X87ySneSO+GeTUuzIk21oLtxqekGVUtjn2kJz0WYk
fTrfltEy+vU5TM8VCYf2adhzxPgZiCOJb+2wSztuu9+PlYG5sFDIHJCyzGnALr/N
675U7mM9AON7yeER8DNfEGRJgLNqcxF07nyd834UJMUDS6P3Bx1L5cUuHbG/qQcS
dz8TccZOGi6h7yOGCMmCmfxfd7Pnza28xW3kcBY+A9qFN08j7oanfYSh7sdPCZqN
07p81KHBKhWYnBQs8piPakEu9HqNj2d3UP1x3bheZm6Xi0G1oVEGbFYafNAadRYE
PKXvO+vAGeXR/r2OC25TNEcrSoqV5m17YCeoN0gYTWc1TxQg5MpaEa8Ut/CfRb7j
Q00at279hm6jcBMmXq7nAB2czh28vBNOI4VtNj8K/uXHq+J/61aU6pQgAVDIsLmd
QqXofomXDnGeh6jl0kc9tj8mJX+lBh4PC5fFVQm4bTbMnWET4Dr1ntuap1ZepXlz
aVadNt4cQL/GaLZBsr8ML2aHgRx0kEXgUdysnz4pxptvCB0svXEezqf9hxKD/zdj
rWwJSEJ4jmi9nG8ZKADrjQ79YJzJ68NeJRrd95JXUqPTTfcmWu6bC3+L0JjpkolX
RQfhDA9elD+apyTHlxAYn/9zBEJL4tGaypcPi7pyvJPNz4UrOAu5FshU3w8vPtxw
ltw7rBZXjimJ0D/yy2SifQaPfHrsqZVXOsbUYaA6XKCYk55t7XMlP6NjleYcZ8EL
YLzW1oC+y6021z7kPjBiRHR6GqnwGHtNa69L8fbqRJnUW5c48KR/jCWjKPKCM2i9
EHr9XqswsFjfcyixrAafzFDQsR73PzextlYG3yOGINqe1mbRZCQS84cq6Cre8P/z
lOiXWLDVQKTH1UCz3iT51eu8ayfLHLAcA47PjHtryagYomajhWg9xqbdEid3sq6R
7PX9udHbpYLPoPAKz1IWvkJ0TosG3bpZ9rb6F3CosXVIIJylS44txjwuj3fqB+/3
GcaPsn4yqa7ZCO0NU9LxrxDevT5Kdwr6eYTSfPpGPy41YFyi71cy6Jgxl2HEuG9c
tQV0h9IzzLDDVz7bl5vTN61CJyCX87k377t/zOyUqlY5sDAWJJny7QrcULITMS/J
Z3Xh1AeyqOo/ht82KbEXCs7vvh/bjDSVSTghUUO+Sauz/AJ0B8DQNHjvtQtu4o/K
u8mEVQV4v4Z4C7G0l1WR5qQo+2yTKPvUAiYAwvXPLkdaG4G62zWBtCdaTHhYRrq9
wxLl2AC+ZeMj6TFRaZAHBuWZBnodkli3bOw1lK8aYsDDNHYtke3uj2Xr6nR/1K/G
XXUyknXlhCa+lCtbj5fdd1oiv4+IHM/nAY3SZOPIqsac+RLPgeYGcViOEQkLZsSI
Z0tDLfwDWK/f2u1gEgHBGKTSSWiwdSIMFX83ItE7L2acuTf9KxYG+vQ+e+s5/zVp
7QafcqJAeanpigXMqhuEQLlqn1SR8xwPP7kG21rpKCmoHeTExgNwjUu0wJT1uBO0
8oU9a+lmOQDhuAPy/5NjbBQRPZKpL0Bn0raL1EAoDlNuSYSuTEHXS/Osx37sjxul
GBfFIB9pot2jNCEKohrsJ/U0SF0UThmnHQx883M5G0F3v/BzH/5qSpTPae699h4c
a6pz0+XqAYy/467UO+Q8Es2YuTw2ibAmkHt9t0k4YUuqH+fQ4Npg87KxssEwAQL0
rOBJf2tTeD2OMiabExG5lVgRNNfkhGRqsBeDwRRTkq1jXq98h6IvVywoJ7wqRA/e
8MJeCwRnTpJDNnTv2Aaj7T5vyXY/T2tWfuTzKg7PlQIkzrv1T7Fc6rddY6c6bZTd
x7kkBoaRrvTpr8d5ScfWHabb3TW4oLkMW+wKBm/5ZruNlP+js/kert9y0OHA4geN
tJb//4YPdFqfi1nNWQu7ox2GUyyrORiJOj5Prr100PG+DQlv04bkFiAWsicERq/k
boDspSOd6A55hHCo3oYnQzkm2smcL5+/IaRBrlDrs9uGz20/DC4xb1yC+6yaktN6
zb4kkElqpSd7PEn+/cGQZpPr/VpclsjzW+TuLiiK++qt3mATcyop8+AXPF2k9rwn
3SKQtFBNzjDmFOldO72pLGWQr09T6T0zuHUK5eeeYRBNoPC7WRpd3sFpeUp8aX+6
fwVN2ce/ijKnr7xFQwqRVlVeDScgq/z1tumnh+3clPhGxG6uyS5yfx72RasRt2so
qzq0ou/SPiID/RQYW0ZHZj4Tae2ipfMYD5eUB5PGiazJ3RO36gztanXrlbqnPPDq
S0dSUwhwk9mpyGURXZIz1LCfZwdhqlcras+iW2RrHDOjSvqNrQyiGAKQnXQFiUvZ
qa+n/BD4wn7YHaGVYXS4sqB70c3S/e6yoy+T6O4goFqGOpIHu2+BVftWIC7AyT16
ABwpI5PItAb5FAZI0NNGF88on0grg5KuaWjcvpHY9Z/VnMBImoX+mwtL/K+m1wxJ
0qFGVU1yCEG/hWnmCsyBGPjr9muV34inuPz1gQCnV8xC4ht+D+IMAMQe5z8IKJ6M
32fIe6MQfL/lkZuTKp7rt8Vmt7aZaqdc+3KYyWAvT0+Op9JEJONoDCEkH6yQEiXR
d56ZSvhB9ojfN6vvUU99YcCoQB1/SF1AWjXVx1iBwjU6DonTx73WWjHVV9mtsGAY
6bo+sopZhigGunff8ZqPtdx15ABEDfmbeDnsg3nThu46DEfaxpQzVgl1QZg5W46Y
q6RrYQ/c3mTItuMC/YG2XVcP5N4D9KHFg8C+TZjbhLDEqlkGEopz0INqg7jVYoVa
HTOe2cDRjhAMl0Fhvu3uaUAZ4FTONcNasF67M81JBN2TJiezubz53Uy53BiGDQ+H
YaQdQno8xZIqttBt7TPAY9Xei6XyUi+NQMFEx5wmcneqq9KtghN1MLWtbfWEDU4T
Qf8WmKqGkkPUi8b6BaCEriDExkgRv/HGO3i8lDn1SiPyqIPs2wpJPyCmKdVIKgGS
S+w4S9kHmEbRnw9HK3Ciw6bMQz/Iye6jH8rOkQCsqVUCwtOET9W7v+9/NkT9GKF/
0H+DNrcCR9rQaiRWGDdSmF4mFA+WPVRqNku1hbw651L0L2kqk/DflqjWNfmnoWen
83xDmvogeWfptAlREcW9G4Dneps1ry0pSke2mTbzo14DZqvyobJ2QLkInqSUQX+z
h2OQv+4AIxJg3muN2rvhA0IWdSOLcmG7+9PMPZsJezJ4z0kSuAsyvd6Z2PSYd8XL
thP+MFGBg6ORQNTtJr/4nBy8YjCbV29qmumRZDF+LqlDkwgPP0RgC1K+3qR8wVJ3
qjbv5hYkNGS5s20UdWmCteeh3YCNRUYShTSqeaV4gRAj1ysYgwji/d59YTb5MzYw
aBT0n+h/CKOkC83MOcvPiwsstuwxxc+G4tFrfwlBm1kQrNNkWlLiMnkB8MFRf6M2
ydbxRDwpQUt3fMcMmDnA4AJIseHlZGUBy5yCEFMswyxKYXXxnBPoHmaZ4uT/EQeo
lEQvK0O9mvjwdbqVVPtMizF0m0XkNIjrMvrLePGQCXXz43Oc2Jv3i33MN3/w+lCY
H/eXXYeiAazkBfghPgw5SFvbBWLy6LNhrXbZ4JiJ8eW2hRY2YT72B0t+H6tJWTRf
WDm8gnAHjxxnKg49/B8VHChlFB7BqsccSxl0RJDK0JpWw7WAyfZIqJ5QjflKPFWk
R1ZBoFX47HVyDuJxACmSGFw6/sBmW1L8NhCPfwO4QY1CMn6PGisUs4EaaRfxSIjZ
GETxYORKAm0YgCK0w9tzUjbx3i4kXQmQC3M8QLrUJi/tzNGswGOiQb5aonrpDAfQ
oD7N4fL6I+raPSBcGAJhrlc8oTTvCPjTfnF02L5qbzOtqOVMfHu67W0X+Tamtiya
YXIA0r+70/duXK0WJ16LO8F1sMTGrQaLqmANpn/RCnuHR2u5QRRyKnS7RTGi3LPA
g8HFZG4o5vB7uKwwWnXy4rIN9AHBY8Kcorr+xqajV5Tsjq6vT+NkOwRg/pEDLftU
BRSmtPZRRtk0Qg28x6Bw/S+6oMboVo1haSfF0PdI0Ir/Qezykji+jOkRZhbIgzvR
+oZwg3QzuVXcnJijrAM8GPUcZ50eG65OYtpsS24zk8mkjv47iSOBMXyv0qVJraK1
AL7RxpeLlP7/RVCwboQhOhrf5N7bIk5KL8zb3Q98hbyGha2FR1UJxO2+yhZHCe1v
3OatCmp83UT18C1RzvngQc92+XFOgfPhW1hZPnAgEtMUAsu/pvDLN7DxDHDlw0eU
Ves0CRrKBF5S72o31OQ5ToiShoTUOKJcXijUhgwLlcIqRbwlCCN2k1AagtYfJblB
BdlxnUNp0tgTZx3k+HYOS27CYrrAd42ja3SzNbPok5Gin5vMiLrgtDme+saQGc+W
Iiehco9nTeufkn0e9y/nroNShqw+cEGdDv7YtsEZPJjjsfYLjyaIYH/O9PNCc2BL
ivmifwA9jkXMiJqHrfGalFJUCPW5dqrGkd38+ueh8EqR4rJBtLo9iXTqE7rrVHqr
8klIYgCHrIw1OqaydAGYxfAIAfgjAjZkiMS2TtW8CdkAWoQrWwqoBtIF1PHOyzNS
qNji7D1HdMUNInuH8MtZPM1wQEzizjtw/6ZB0k3hMHjxpuB4DbX7k7gLcfux8SZU
/aMnVCpfkmqMJMcu9Yzw2uVxSmOVctli+YtPzlwt9I1LhPY1N9NvRIxbIZUtsHu/
T2I5JrcXHmH+7Dqkuda25Wx9eAKBWQDc42un7cUj+tDeNCPq36s7mqfKF8Bj3h3r
OFRLeeTVWzO6vw70LM5JEhJRvCUUEWSP0F1o3Qo7VAycA918vGr5P6OumXhqz5/+
b6kxKxke00m2jqanpIXO/5i2onCxGlxTbnu7yOscQUmfX/YqH9voi+sBoMAxlnHO
1PxHSyFuPOCgJ79otZKCSV/rwrLvK9Je9wUO9zUanbtbztsIFqxfSTfMNL6+h9g1
moF5ZXgIXeERRg600okpXFTDuDluW33ljFGdA+ROo+X72EHMLaC1dPbvuIa9c4aQ
t3OyTIRc5NH6R43xKqL2PUjFzgi1COVO4VoiqcUYTBX6mfh50B1GPj7gQQkNZelO
LAoYggBP6FZBqxq64R3+EcQYtZHGfnKhrLJVhQ33uSIIHPl/U/Gq3kYGeJDmNlno
SmX6QM61+zuAYfh1LmM1PW93gMoBwZpjnQTR/LEeddvbeSKjfhy2uA8uwtnShiPS
5FPZjE4beXTigTPQe+QLJtT6hIrGO64b2ZaINlcRKJFuIR6AihtAD7F+SsAlf7tX
jo7XUntOYjm1uzNakVCRZuE8Rv2kmcA2EPiCp4PA4UT1RfNnwJJKdTvuidanLvKT
ACUfGkN4Uk/272HaVg/PQdykQ/byS8tDYZOmK7Fiu2IXVpWIgu8stTIO5v+xqUmS
xPYCFeXCVDsldP+2Bf4QsyFSnrdbMl23+NlgvmYyINv51399ZlAsOWEyOaTJm520
KTQf5qT7+6rljAjdxV2AJWvSZ81sax7GS1xvKr5NIVEfB9y3hgxdK0xf/cFSvtbQ
TyikhijSlBU/VazKGu6gVVdMjMHOLqKhIFPKVFgrkmPem27peCr1grys9irNGMle
8isivGiLG8ZVFcsBCbimD5YlwhGJhVxgX138ifmNLCGVIkvkfOhYpJgBUjwOalGW
rr0iDD0k5OiA1kw0UIHbJVf+saK6cluEvATGVwiVsSQh1klp7t1DBZjVjJBDREq3
w2idZWBCFzkNszGzh0PvTfc65TXVT7oIYXaIEBTtvuBw0jhOwDhM6hluhxVfzxfx
edD4aj4NDOl2FpBT/5gbWzdhg+i6xKaMbAxylq7E6uifoD0uutc/r0p1p3d6CsCT
88tZpuxwrema4koNcaKFlLLU9FKUweTqYVLAYZ4HWB1IfJxrG1xcP8M3F0B4ci1x
kOU35elRVbF/sONRx4Tmo550JoQBSEkkSpxsPlp/e3pktBYoFAnlb5+Z/f+nA935
WU9i84gZo2jLHSWIGCNqtmYyb00WInvGgIb/QLuxTjq8aFZX8JE6Gu29mQ9SFJCE
Bnbtq69X39w0UyFfyvLf7sjSOYVOdSSrdxwBmJ4GBArDtMVaeH5R+4gQtUai5CEQ
//rbulU5lBuQOyKFJ0LGyvzKuWSYzQGugPpl9lsDSOke1KZKRyFsvDDvB3Wj+hAD
+ARVQQs2qbeSs5Wq3YEKT+HMNHpVRztjeg3UqVLWROKpklw+gCwiB67AFcMxROE9
lvCGSvJVyvjs+7vWxdTmooatgLMgH0cde8yuEhGKHFZaw2Q9XHQhJHCiFU0ai60U
+Y2ysN77KzJnuOSx7hl1cMpwgAzmLFvefLWZPORA8kEeul1o/xW4LwmlBjw5Nqkp
uMVsXPHk8/RszNlA5s4c9hEjpLJr4pgM5NFOSF9w0Zl41283g5JXhBdDSDDhlc1h
hOz209AWSvXuoo5inkK/Cn/VUqzOF8RVRYBuZCXQrd7MnefccRKsl+spVIl651nF
iDjapSd2w4y26GxOL1+SikINyyR5KbRWstyAJmC2V8VzYUO85sTjJ257Q6V4iMQP
1a9eUNnN8i5UX+blnv8Pth2arApPWowzP9I42/p440/lPLiliOA74v7+5yNpTlzy
9fpsnhBQub1s6ZzHF3XioPZxlRIQbrQvTqdFEgjC406Huyd1D3fDWz8M4I9tQxDQ
xccxyIjjl9VrQVO3TG84+mTYWNaaLfOBNEomEDym1EhbB1szXZeebBxGNv2M9epW
Qn1ouwSQPSd7gl/SZxkFvEnwmqA/boKRDpgqfHhuBfMlzdkhxdIDUWGyNs/amrFJ
qP2Kikl36YfPvZt27s3qLk0bICI7U6hNpTaMpolTkXS2P+udNKPu5006ZA5BJp70
/3ODk5l6pvM67stP8xQgp2TKtql8J/KoO8e1OXjzG5bMKm+Hz98cIWSiDKWtfbhC
g4M5UOg4hm1zMqPRCRiZKA0+IPUM4mo0V1rqi+fjJfG5h7g01EhPSyvl/79/k1Tj
sIPL8svCcO7XW7Md8Wyy9AmCGnoXDnAhkFkDFGghjxdYZqOfApKIlRk1virD5BlN
H5hAJBPFvTL8JObbxUGW614CtJUkJqGDnIGfj/JwG++/gXp8tFQd7E7zsnPxsm5v
oCDzjRjLwAnVMvpBc9eMlUp8yN9bOQB5JJdbh9k9NEn+RvLF4mwZhw5jPUifO/IO
79vctcsMPoomxGFTRdOhogPULd8W2nS98W38H2Cdlayeo9UnBl6H+L3h3M9pjRwn
6UtVSLA4LZ7n1n0+e5IxvWAmiD9fXwKJIMqN5GXNlz67KRNFqed8WoH6BrljTgdb
PcWCzaAhUA0+tXIe1DKE4ciNiw0Mr/fsQNXyE/hqTt0y7Z1CZgiAP2OulAZTjaTN
bJBRO5593mb8i18PiQ2ovw4xjcGNJZvosuxfkwpPDm9f6x+Mccc06SV1XN5SFqE9
hhUSeJcQcneISRiG3I48xiXYJpLr/x7Uj/gSnpq4JrPHSFVz0AnPD3FFcnZ6cs7q
wDg+XDrZB2fkME58Vwd8SwmFd0t5ZtM4t8LJwgdpW38etv4wS4huKQ/vupGa8PoP
uT0I51Ptk26P+V37QWGefV2i9fbNmkqSV43CPEp2el4hijPkPfCyGeGMKhU4zgNW
Tek8/7i93uApPb0ZWCNuvcQQNr+nj1VWqQ2GHWijdORnLMn/cKsPgyLtC8miBEL5
vzpbm0QxxLBMfSrn/5d2Ddwb71AFFP9yi15B0/9gb1OMesZ3zm0N+pxsoyG6099E
LjVN1myFDiTsEpUieSHxiInCE6zZp34RG14vIuriszRre62a/+OMcX5IiU3sik50
X2PxsG2w1fyW8y4bPmYg5TQAP7wx9PAnFB1hCA5zvAnMrCRHCiKymqYTWnyHXEmy
Yvr9/SGf1znVO6sTg6fhSsL3AlljEJnviGs5yfiD2pVBIFNfjAegvJu7GWxkmrdz
sazntKttAKRakxK6OwgO2KJ+DOVUVeldAewQytzBEciVHZF3puOE8ggdfI8DF57M
rN6GevGUmQRwocKJc+pRqeAlbQifO+crJ+IF48wUILPcyyHYDEBHHdvoe12hMTTo
Y9OHLP/8lg1JIwJo9+twGO96k0saB0/2tv5efOXD4NGzAYVn2Eb6+11A2AETY0jE
yqT+rlacX9aHLabNc//OLdoZ5XHZBjMlMxLK5i/2lDeRGvuEuekjY5Kfdtq679tM
UQzX0SDPg9o3DuzV50iOUdSED3aGV87MNI7XQQc7Lnr13pzznCU6Sp3msUahiS2g
IqXYtROV8F6r6OeydnfOGAIa2ClfvgE0gsIV1Ql2v/LPhnqpqEuPVuDXqPZ4iVO3
FmaPe/+g9uciBLK4QY4bFF+BLf+PNHUOJsBlQrp77KoTwZ2l3DqjCTm09MtkuauJ
J/5tHjIVRzGtTWcM0VYi35qHSB2afOMOw2uXuNulm18KB/PcVXdPuygWJ8RNoEsZ
A7sFp9ZNOBlUaB/4GtCfTrdxTp2QyCbUaMGifcfDevoV19fRHomlcuNcycXENb53
N2TukOTUMqfpj+qBzq4+9qdJaMz80eVLBLGzjbnw673cVtPcHPciOW3in14bYrAb
/qimyFgDK/qoOh0IPKbNFvptoVEaHSXySZULIUNfLqT7jpNJRhNxdTg+5/RJ/Szh
QH8QrtA5taRU+MAr2HWk1PDemHd/yZaN7EqypSi00TzgFXYe4Z57gWmssZYLOm+H
QYI9lTNAGIckGyh0QsdDnNMK63okbzh5WKdihsx/M2QIDI+4fVFmdR0bJBgF1udH
H1164LyL7cElqjD66CSP7tz67gDBzw1VJ6Wwa5vrkdheQu1xdfMWyfZwk3QhDN2W
WQBiTfqa7Zn5u9vv2zWeueeLmVTZeuGdBhcvdvRD0TlXr3undW0Vz/xgfa86yJAk
JKOMymaoQ/whs1dhKY32H1HuOPCqW4z1iJ+2M6XJ1csCwNT6oFZjgn+ZOg4ZveYX
9Znds0gwqS8Pb7gBd6n/CfE6tYs7W43E9GOSKhram8bOnuQVvAGFoH1EVhlV1GGM
REXP9soFSC3dw3bwJQkRJTSXuR7XlaIww56Avid9s213GTKSRKeYxMaHsXcIwhYZ
kmhRxatiG/w0MBpMqGcvF44pH5VibwaA3cAavUIv0xJ3zeQZBc1BOUUA/va6x6bO
BwECDVUpu+McQtLZsZR/GHewW+BG4ND6wJ8bAeE9iYWFTHmdScTR+zOePYCCIxtl
rmw9SWQiaLWLXSq1MoX+qTcUiE3xYYw9LO5VzGRdsyJ1FOmbUDjQ1mjiDfI5+E7V
8izuE6dUjhTjdVvr7UqpRj2Udh3GhzCA/iv22A29Uur5KTdbLI4O+Tlp68sigrOj
IyZYAMwQq3ixCBH8zd+KFsMYv1nNLrBYZM0isiQkpdNVUc907hj67Jhs9Wl/oUxJ
lWNW9YF6s2t9DqoAP8pOOvZdkCWYPBYrEdTHWdajS+ZIqb6lKEqTr8StceCOBTbn
9k3BK0T6je51yIwhHjF5oQkmXsLWzjCcPX7lhDu8MtrCjbQzfVcvzqqU4lXoDMUF
WUnqpOPHuot5F1FTtSH/FKj7ap7LPEz8aurALmzDNo8GNH6ysnki63nryMU9x1WX
0yHAeZ+9n5g1VnepY6EoOFhWAmFYMZWu/Wwyfu3CTrO6McF8VG6xYwzLdSs+xa2o
mlTom7xAm4nDjiUPNZA15ILHL3Z0sdIVfzAdM/qy5ylZyyP8/1/HZpnXM+e8qrcG
69d7zbMpV7C9Ty+83FlvhdZSOmOtHQXdhJkFFpwSkiRaKDv5exp3BHMlsRyYd7bn
pg+Ud1Kr0oLnjcFDovpog9ugYZFzKUF9yp97MJjN4I63p+IAcx0553RNE09JdEcn
i8gEvU9yU3jy6ElnY/5IzNxgbmGZYk2dyfFNYBMUjlF8ttMmwvA6bMrBoZTy7yy/
P8lxtx8eW/NTj1zbsxfTTeTJRNaMtKkzG6u1P/4xr9Ds4PW2gjBL9bZqlcpGnUWU
Uq3yzBXEJ9Y4gUX1GOeb0I4g+U7EfphWtbTVXxKHlAzHXyjquG2f+hlEKaSsFMXP
okmS70a9Y/gB3qQYh+v+PAlOaFGFucREfvf8u9SqRAUrNma5eQDCNvD2LBw8P4VD
LXe8SlSkZP6eiflPzPXn1Ck8ea4z2LyPVTlPHxX/DZXixronjEpA3HAFpHwSj1kV
K+Ljrt9lkzSihbOTp1ZUCuchIcjffRv9FIiJrVGBTthGMNVH9bP8LkWj9CDT5cbr
/chR1gzCwfP9mQwOMdbU70AYtirE6Th+MkwVEZTeLNgM5Jlcb2qs4HBrWgub1BxL
s5+at74S8iJ6N5qiWy6CND/lhWpBezyLEA/4xteZJzCVjjBNQI4+WHnMtsDDKxZ9
j+hwYJMHmCWEUYcFBCTroTDIkkMBK5KkHz4MZD8IOdIpNB80aOWzQTNW2tKOYaGU
Ou9g9Ysa5JAqRxHbvVm44GznkiHAePyjvFke4+hWsG0y832U87mH0Kfql7W9Lcup
1LD/vtv8l3cQEuoOV27oRuaYfn9ye5kYzepNWpn3bcey7D45dsVMkBAew8KxUl1E
OswOSYfQ//HeoUOC1DWB47H0fcCKd+GjFGUAMqdnOlpBMjWkn3rdZ+bl5yzaL+Sf
76mRL8V5KVbPaXmWGl2Wam1Kur57a4ZL8kR186IYhWwqG4ZlZbDDNk3LLIMAs/pv
jt67Io3SSV7grkEowcWNkxnBQTiFW/OC4YroDQmPCta06pjS6o4tgOz/jukUyiaX
G3qDyIOKLmATPgUfNNbD1TT4reVn1G9R2OJogLIithoiIndFCitIMHvngYzvTxxH
W2QkcasjptE4sTzhlfdJMmmEv8Xh2T1/9Hqekitfw1LXWjry4guWar73I1FQXjtC
653UptwVu1oUpDz1SNLsnXVV+42vWkleafBlf3p08naWlKs2pyvI+a+Drz37TMXH
BEJNaiE6x+bis+LeZHU9LcdMqyEg+UJj71BgS7Ve5H52Tjd87l44f4CESFFXmQzE
KLjs1yGt4Qc0ZRiGdTt0XXan87CMUAR6+3Q88MI5t58AloOf1ewmUWffJ9b/EhoN
927CG4YMrlFJISxe1mvfK8K3+iJpV5+v4lmaVeJB0noowuNJaTCcCuF7qm+BXer6
f2ywIeN9SmV+nkfvIvtHxFD7aOQp8nZa8GuxXVlMxGQQ++PSQXb4c/iVZ2CEfV7x
ND75rsrW4vEG+WONXrisE47nOJwem37SgW3QzaN4TiJP6tZEDRLtxC1ytfz/R5P6
3TMqnOK9dfhgxj2w4XY3x+JJrvXitlc5d8cfUa5qoxxAuQ7A+SJqkfb7uJ7W+YYO
JMaWd0BWXAzqPIgvupLMxxtsGj7uYawCR26DvQ05XzpB7CyKxDgBcxQF5P0osX+h
jRMg/WKwVmE46U44Irb5/RnQ70oNSvH9f7I8FSKBhf5p59UppmJmVZuieYyndOj5
Lcy0KMNQplNhXFNzMN+lyCtRF7PNSL85WSQiP8OEzKlts7UXDT0avzHoflcgbsEd
Rzw8qWE0srVV7xql73jiP3QoADYdIpfX1f7wULwZ6IrR+ZZC24gKxbRv3TF888mc
RNz9H/+BJz1iAr2prcoM7JkGoWHHXopFf75yoZdkFJpEXlpa0eZRiIJZWwI+A6SI
KmS42qopc0gvO04+Wxc57jeLs5XyL3SPrXqSilifsXXiRMY1cAVzboTp/tfL0CKV
B8KILzE8YwFQ1hKt8fYSt5V4ukcALnr+lQeogFNxrgBgQTxXUtLKOfKqg0MHfRu8
VPAXJA9C1DWUqqrg2LPc5bnOa8J+IJciDhTh7x4NK97zM4K3LA5uQCE7L2v7bb4Y
wEnTxsc4RuE/9uw1Pv/CBH8ooKM4QQscyTVHYqj5C3Z/ZgYlFVy12HUYjWY6ATD4
Djl504GCTcLMQmlL7xIGwW6oC4XLhozoMJ0a0L994QJIZpDYRkIR/6d2xZJVJz5p
aDTUxfXH3cSHvRZ5WgNxUQlInlad9e0lEIZsnnP2v8lkuyrimqo9+Rscxe+1EicY
jY392OQs01bGuJHaFPt5zVeld4ajAQMpb4oEFDnTz7CgA/iOrJbyR7nzTbYOT11M
otEyZDYGIJCKniWhBIRlZ1A87bGCe/lJh3j/WVeBGdTQ43ndeAezO+cda4SFEk2B
+Ikm+/0jTMi9x703EWrJlLBdu/0Oako+qyoKwMoojbdoEmChOCkxM+tgAPZoEop8
zuy5l/Q9j2WZWPuMaMps8XzSbFTyVmaML8BL5u0uskPsbXiHl2RgAPR1ogbdU/E8
Brg8tLbmRWZmgImDyDD5rdxHcIYxg/wMnNy2ycvqghkrgJbyO20b0HZkvnhC4K2W
rZnkcT+Kf4/ooc8vVz/g+FEE+TxTkPB05oRg7b3aGXJFAw7viLJqOWFk3t/UcVEy
UiBM3YqHDQWjFlAzhxeF7Y77Ih+xGN+D5XW2qfV6+dnC2WiDaPsGgvukBtTmBHSq
vC8C3l+OsJLSlKSh/pqPWm9LGwPSeSSmRFII4t2TpW1SZmyqUl+THDR/+jH3GXr3
GTiO7yFLAQMQ7F4xto7oRu6P1Nw+rAerc6y4Lg0oOHnzEi88ZkgAsf2ORfRmAKiZ
C2UQF2CT0YQhZ2y/teUfVSMCA1arGprr8GQwotjQeA0GhCb6U8eKnvzb/eDc2KoN
OBMJeyWlJXSzTG16uO273aB40rqe5rWM04xq++DQHNwE7DYRB1JHYwwitiEVituz
9+cQcLSlknsyZAEQ6dXylju2DByvj/YxeiwQhjikfCc74xv6NY9rSCkbE0/kY9ER
grNdfJYEMGntRjmUY0psvYcsMrI4m1ikcRjQHsBWp20ww9uUfXH1n9EQyT+uA9ZG
NSM5NtcLqmpssx/H+5CQ1Nsjz4sttnZqq0q4ndIiX6plvI/oLf5pyYlaBwXk+iz1
fV2LpzEJpHpWxsTI7fN1BWUpkEyqos2z2YVf5AspmQOEVlIPXr8/5uDAABcwGkhw
u1n0V0o3+nLgjQoFU7jQXdwZ5gkpWMGB6mObgkh4SXshu86o0heXiYotER2r9c5p
smVnowIjDp/40hzAtnJh+MklJIL9lR3H5qLlTfF9jNt4ymEnujpAEMTOPSP1bgSv
iv8xK3qAraiTxIs25AgV8Hw39pabrAfy51rVztMUMXhi3oKLl24yqb+SdZNUx4AT
5edw22rWhUVeUHNt+XqRQmraEuuPaYmBbmra4TPP1aQvHkTiQb6+iCB21a6u+UtR
wVs3D9tj5UsfI4eveQdec/vnjNVm0bnEZ6EmNJUErBO4Uzyu8CXKvax5rScUukhr
ehNhT8nurQVNfToK0pI6Ah/pwa91EoOoesUz1G362gOIaRFsEPF5bmpPVgSV6/Ge
JtwD7h06KtGI8Vq9MG4zd0OEsbDNOtMyRIDD6nALFAAlgFPHhpSHazu6wTuo3zhf
VnTfg8cip1gZTB+H4pcaEHdMb7XtAOEY9U5fYjyT7i4kkO8x5zdZL4sQJ6C1XKdo
6Biz/jtxyfqAQt2VGhiTjt2dhGLCrvUrp/hvPLN2Mfm8KeCFH36Fhcej0MR6L9sf
hbCc146U8dcMTnX1J7D2qHdo7wCVfruHjlI3xUgHwXsJDDHeK4QXel4KkGdiIb8x
ytCQGsPJ4/IDcm77vaR+q6jP9dTiJ1bvKMprGKMfs0UbCA/XBLYb/CaA7jfIbiNo
3pgNekkwS9tEak7C2Ho/2r6WNKe6zdBBksAc/FqgGqiWXMwDpKjl0R2X8UwcJ2R1
Gz1qoHiLkORrA5WVZ7+G9PXEcnNgnO4s3zNHTQ2GCJe8gT3/0f76LvM6JLvCBq+1
Lr9oZKMA20YPnOMWReWmR1P3NFuBr924XxGk0hoj4u8P6T5Go5O1JOlrUTUpciTu
SOP85GayKKA/vcwW0hEt5K4SwbT1Kgb++JlSEP9Tl9H2LVhgqv/cOn9FIO3tMj5n
hUwfRR2bIULYsCwRy4475ktL7cHIe21yBa/xzYRfD48zPvmOszZH7MLoFrxhX4Bw
b5aDA3oE5/o2c+z75YRkHzTTtw0R0Inbkt2dFNuI4loOlaCAD1thl1ZayS5fA3Qv
jWKjkinxLGCQNbet/g2rjnXNpmah+GtaWSqJPnnLCIplwrgSO1Lg8t/PBmdPi/iE
xikm+LQWTjkDP7UTTjv4uQl2vyi6Z7mFmXC6c6hfnPLA9kY0K0F6DsFwJMckuhMl
7nx8QQ3jEYKw/Jl4doRi/vwcprido06vPP3yVJ+Nq91qn+CTk1XTXp0UFYGMtGQr
BbpQELpTAc1m7CNi4u6jlhsNk7ya4ejT7npv+8c4FpqbLoXTGsaIaWMbpqW40FrC
3jhu77HrfrcorleZ26tOgTO/PN4CKoS0uXbnh5KQe+fSlJpDl2hqAdk27REXcYsT
xR8hGeMFSRuiUY23wpT8cSrdJtkJvh8lJJUF2A7FvwdyQVcz7l752CuWJD8H21k4
LIhaLj1o1iePD23vWVItvYdmvETawzbENbQ0HQJbh9q9Co/9r8kWSCZq/dwMCzK9
I+ts857/2NtFnQ3LRjn2Z2agKK+wuXgfEMMkUYzQRIis7rtApr5pEPxGR3caTky6
Jdi/p4QhUIs5UR8AUzUvYEczXVgH3POnIXf299qWGKz4+GR5a1fiIeRz7/+Ahrex
4Vzbi98Xj++kE1mENvou5uwOUW69JLU1C1bepGGtjg2SradsDuM9u59CZc9w1bmp
pYF0Clwm4NfzEq+sbRkV+4SUYyAo728mv95yrDAqMnom+bknH0BnvqCkmyMPyhSo
mcpLL3wCBqhjN8WXLXC887fDFwakaZ3E14gqPocPNl4A7YGHFheoS7mhVeWz6aRv
vL+xq8wBim0PfqQaxyK5h1ZPQTi4A1Nfq/UPXa3irGyB7jU1ucFa2mdMdXt6hiud
9tRZGQwl/Y8p5CN79t+c72/BXh5QaynlfN3M6jd5RnRjX3nhsCpTX9aX0hhTlQCd
LK+f8Xxdnw1+oj7jEvSXH8rYPbnDOsKvcrz0DxUVEPqdVm/DgycmoJAsLySOL2AJ
mqxuaLSOXlGpuO3APpXbLS17/WcUr2bHgEY3Sbi5g7poPwR2U57UY7wmGAdY9oRW
1zSZPd/CFxCuVeBOWrMxFSGbdhQ5te3nU84MsY3R+iUs5cfqOosHSz3zPvTd7nil
RPOsYRp6fPYcKlHrgp0KwMOsO7ZLc2D08dYkHhfa6Gcd5UFbMtbmexyLj3fRDLgT
BS9MbOWP6HUcgtMEIJvuevj+bnca9mL5aWM2uJYDjkan0Q14zjIvo9TJwqprSl7q
1fK12scZXIITtsmLO6OwoSi4kjC1QP25DWC2eLVepNAqhHgconslwKzEEtqhZIl/
rc/+LEmAFbARNzYY6c2zlOVjhbJqDF2EcIkEtaf5XLVGzQR9SOg76dihlmrpaRpS
7x7Tp5GDM5l7FYro0ZGVTuTENZZ52SZBG5Oy5rV4JTgwLhFkbLEURNvRZBoLZqha
nrxspRKKwjhUapo4bUR+wXUlT5TN/pikpNeEnzZdN3biEGv1pYTYuVnvQRRHuCQv
DCpIPEUChty/Dxzd1lDN3AoCU0JsNfKRujQyQnsmG2vh4LL712u5dgtoo/utDJYX
8bmYxGCrnwPfgBK7k5njCK3BX46vMR2aIa9PE6V/ZkP4eV4zVvKVxKqz5jf7Jg/a
IJmBf9fnv8gDqDYd1551mvmKu9zDfdKgjAqP6bwO/qHrkei0ei4CmW3T2SWjvkT8
UtiQn1e/WpHnuRh2AFascpcngBafLeSLK/n+F693LY97ReWytvu2bg88FMFxduRa
ku7z6+3tx8E0WkcTaHxaVB7pzZeVcXBC2hIH/x7xa6jaz8YWASoSxKaWCp9nIFij
spE7FuxbSvBXn64jMjh0+eVh++bvP+IF/l1FlT9P8qa4KcIMO+nI8khMCQa9gokU
zEE4ZYsTh5Sbog1a6WF03pRrNVX648K1GKn7mCioAUmHSIcI0OJukz7LMZF6egFw
6sZE7g0ptZh6J7inUJWFdfuEThJgAXSVDNIjCvMbNVhrjPrxcgBb3wBVOTVPAgfN
kEVrEkTANl9wxND+aAFkhsNzi7i1ZaLYasXetL+lpLgs9S9v/yoJTTlIGp7PnHQQ
f38UXmbywjrKSykWdKNLWIuqJYM3Vyy0HWjMK3UvXrm13oIx3XuplXAurjEYOQ9r
jDgfPuZS1RGBEd+Rb/Bz47jSGAZqxK6IrO3tcadBPRC19yVGjXkDe4yfV2HxOsGY
t7/waVSNnETXXngfYRhOvrsBkbK19j8s/RRXkYSXKIijFm9MQpOMXlcKey9JC7/g
ZWpDlkrgXRg/XMJjjnzL4ZJkEWkLLQeaG65NoLbfO05NMyIvjx9j4RP76vdqiW5t
AMVfLWwpo0VBy2ruvhksSmgS96Yu4xOCuJk//T+Ez1jg0hhsfqi2ZyFt9htiGeUu
8HTj5eyJGFCKlV5ZqL7+tiHhg9MU+iMKJcfjyjL2MpjFDrvw5JUXbxFmE1lBLmHV
QQoPHJH67rxn9qbJAixPH5XmWAy+SRrUcpCdK+5ZKHEs+IXmqEngNu31k98ExJ7B
g2ruJFaIQtXQMtZKiRc9Bu1t8pQ/Yt+4szkaPxjs3T6kqdp4uPffr46kkxlHJj+e
UuFIPBlmXtH4L/SaN63eoB57bGy6I09VpWlJpX2Ldoci2PEJ6AD6SMtEIWljZU8N
ZRbPnRP+SVcB4EmRsrx7xq0ooLA9sQ/SHNQLd0ZOZuHr0oROq/VgamlFAZtKqe6k
z6zPZ9EIK7tIATtJZt2r7esCrLdmtoUZIdXfuNji5egn1WlQEwyE8mlp7qucgxpr
HwPZL38U+4NtzDI0+/9i0WIyDh4X1ExPjACLyaBTecmUCsdLkksXnjeNTvoK9rju
kpw1cWERMvJqMVpRLiH15E3q+UN7ZYDmOvJAi4q3wNJR670JaJp9ykmlMsfuQqp4
WIGUujN8SCa0WupZILJBMQRjH4qjn93x8ZI7Yv/loqShUAQqA0L9kVHq7PeOuiRo
K5XLXHENMQxrduT6QjlxbEqTy3Pl/spGaTURsjlUSixIZhh0CYQbc9H3BTivPtPF
fGezyZY4NFMcWxXFsb90WtpMwfDOXeh5LIfleB//eFvXbe1yKj2d6Rdagy+f7DLW
IOWlEPOJSefA+wm3ghB2IPe240jk5FdpDqCGSjEIwjjnO9p3tRnJPBj8dz64mBdH
U+/+s8kuPwjLyuANTgIRDNYEcOT0xNM0I/ONwHolkTTue5izrgaifEWb6rNF74c7
LTv1eJ2Ry8mRXdLpfOgqglbUyc3OKVDyXBZ34IJ6L7jpguv0ZL2vvGiCQ32FPyuD
wso0qs7vGqD7nZCGpq/5k6d/9SFyALyK+IcNEedVKEuPfTa1khdwuRMrWr//U2w/
XRJ0IqeWHwUvqnP1GVdlzj6t5kKZz7QNf9DsZ/ok+i03FoPalJw/K0hDqeC7umYB
U/L8hAAbhtr2YdeheQK4rI3dUyykCm9cvxuJDt6JybVK9xMhc8nLSkx7mERCOS81
PsRPnJ6PKSqJhX0NS2L/mf8Rp/goVudIL3wK+uFnvwr6UksIbi0xqJJRqYpN78ZR
B42NN4cuyr58HteNLv4mxP5DuRihK9a5k33k0PCSGH5iwlNRxEwUEvp34XBFVK7t
ggenI3XaCeKgqrfs/3h8wKKeJRRVdFj9G8dSnIvIJAp3KLa22c/iSyCOsY9OAyrh
crgjEbNQOTkV805SU9o+6EakkXY76tN9bFECecddOycsMAtQgBLSOmGgzN+RP9wP
kcldsWwsCsfL/CcBkZjk2ACTKgLSEU81qKi8st5eLVO5/2fUGio9gi4NxEC/sAg6
SRC2HTT811VGpJE6hEgRus3r/9MGS54MVKtyo1M2zMO06kUI7q/LOmjVquUIrWY5
a7Arcm0L2GLiRdOpHr6RIBRuWroAMaCYBxRlQJWIjMDOHpHbkNJavZxTTDXdDNvS
wHFAE4lJ0dZKR9puuXVenxVEg1/tGYHtSfyUbBPelsy5TJok9jXziTj9nkOzddow
wfV6m30I3LSk+LmG75UfiYMD11utyQo19K0idttpdwlthVFmmGTCfj+UV8ARvLqO
eIrZcAr/DFrTVaSD1PTYcKfnP2HXr/C4ryDudVjeu4AWNnhJXVktPBBq5Jq72t7f
rY1Gl1OdaWCBUGhigxOuCDXPHCY5sKd2oOSpEpVQQ5OzF8Ua4OAQ9uYfX5z+OJov
zNxnndXrp9bm06leQBSAtYtcvoRDPUDbqJtE+33JHsjC3XfBPGkv2K/WPdkOqrzC
2wk/F2DEqWowlYeX23g/CVxLUeUK9xm+ta6056xITY+/tcZ0EYwurEtrKXsDqWqP
sCnt39mCAjGFzm9oDJMUKxsM2eUDlqRB2wKUaSBeELcj1ngAxROiu3x+PIHbi1TF
GIg3nDgVqpVmt3EOh2JoOoQ3ICz8gIjUiM+u0erE/eZGs+j/JQOomreCqmeGGX2F
2ide7v5aXdgJc4vazkH/kkzD1xllABCGDBfbcUVLKtIImSL+YKKt/C2dYVsUFdHq
UpdiRp+K9BIIjVQe3tJY69jIcIHxYbAufEytjCc6pifQBRbuodLe1PbCy7WgspwF
cp5b6zxiDEpP8QYwiXL/CFN02P7B524JC2UEMHCL2HjY7u5FAK5/QLmBkzhkIrwe
dWY8IjD/zTfDnVy4WPpCBGdQ11b5gl73K0MKo1yCoYdxQkJyrFPTNyyxqdmCglzc
K3nQ81YxMTpDbduj0iP/yXbUqFifMifleWEAuz5+GzJcnIxgoKNv72SZfv9Xwx/V
3RbEzvpVi4K2RY2/0mpnKwLJWLfyGVJFBbUbpJgOFMxSgpsRKEzXhBvbN8uyjJxi
RuARSsEnoysgEVoQqoTxdo3VkwbUc4W9Bcfan7VU+vZ4sa15DbOdwB/UWNAUaOJS
cThbBk8yrT0mBu++qFy142cR+18Ab6j+YKOJU6Ci5Kdwa5vy5/5twE8bvtYOzEhb
BUI1nzhvlzTyQJQqXdtBBSIF1D9mpWUnSqx/zRVdxib47KvZHI3gwSJLylZNN39y
bLEwQjHpDksPGIL2u5TfpBgyA0CtlOcPyE7nBOLt1Y/fH2J97LWHUAEfEOKrqmyj
bw8eu63w6N1sYylalsXOc0LRtJE+OQZkMBr5XRK08SYEK0JwENiubXYL1oa/Zdy6
2iEc+2xd7KiocxJ8SVEgnR5qRnES/3RklOi0CzlO3oN1QlkB4PU0sV0NagFf1uDd
bB28ZxYY7G0FffFgmetn3HS2DfE1rpMO741biyipTIGXjWiEDFz2MbdHjJdZvtWY
8JvOw8EVqKZgZaO04MO5fs7V7NlsQonlt/USs4j8cIZRUa+6LEK7Es08d42681jd
sx2J3zYsEGjkw6Beh+NfSkKlYDMl1/TQJuB+8It+YgZ+mgRNYsqHoSMb8FU2V5IY
Vq9EHCVUrPt+OzB0jBTeZOUpr1vLdBD47QZfHnWMRnuFqTCugm6Pv5CVRGjzsDFB
6QUcKo+WZOp5XvxOcEaqstk1+Pix53gJHPJwu1eLe2KBB2PzMbE0iFGEg1g4Mt91
uLJcwnlpKY7AcICoZraqNVVlMdVvHw6p/836GUkEv/8K38yUb58e5YGNArjTsLje
jyENbsjrVKl4pUbinYuGOal660oSG246IVSwU18nP8new6/aRWqD3sGLpyXe6IUS
WwGbtD+/S8YHTX/0OZBgv1oHrjOQTJlvWQ9VcEifNVL2DOx9GKmYt+puUpLJ8WPE
g/yn3WphJ/fl2NG9eC6Lk6b2Zhe7bY4HuiKvQvmIfDdp3vj2rG8Au8ASKZ+DV1Vq
WvhQni6i/X/93VDODFt3guxMIhH/k9CIxJ/qeRCsmg2cAF+y7vGyPZ0amwDBw4Dg
SwMZUoWvSTGxm/BOpad03RRFkNSSZnbJFSrEFOEx/fBRgb5IlKk8u5/hPIhx4aPC
K41Hg7iM9UvM7Ehf1jvda50+klryrGPP9InfQJZqTPMy+V2aKEgR3XID0tUfoCzo
RboXgZE4ApjcTNxWwSfiUtO8nCx7tEbqjNqqNsF00ogS15Vs8fyz2fkvd5u/T04q
mXgN+SSyZudeHxYYQOsHFx2ObtC5Foix1k0dc8szFxBdWLKfD82wWlUoGARzWAQE
gNA4fOHFB+W8sERXmy+9JKIXobxY95df4aWXZmiL3YMtXnWZ1SARy96PJ28jz9UY
gS2ATe7OTQ5/nlPryTB8f8h+HWWthsW8y4wy2Ap/zBsCKctzJ4oYrUyTCbqw9J1o
LxAGH5D2TdzRx9CgVd1ZhyHO0BSbjjwqJs3EkrQLuTCY3/hLPjCgN6SmMZ2y978G
J+y+iOBMyF0BhLUdqLfHnZrYBq/LXizI1rixqE+c/RviGf11cV04aODas3TE8tZo
3oHhS1Xf6QU1V4NHHy24dDFpSlevX/Ed++F833anPk5H5pyclkUC1/Oot1x43Mls
Krn1CUEIym2S9s1yuPFHgvSXTcSGb2+QkCRme61ThNiXOl9dNyYgO93OirYiGtWD
kIEgWxf+tRlBwUQDw9P6vRfvcV5s7k1HS587h6xTRAuJWVWE1hq6w9Qwd2AVlPV9
wnehWA2p4zZ+3mRwUfwJqsZFkaeSP1Q3/kWgfVGAabd8/Dqm9YP8b6lY+xd4YRt5
afDvnQZPm5AJpKo8hp+CWVI26DklxKQdkzOD0Md6orQvE8bCFfOse3z1ayz8G5ie
bE7AVIPLU/Tz4FF33ruZfq2YvSsRsPFbaTcrt7MiBYUT4BPMd26//d1qgV/9rhyo
lu8iLIwboxE27EPe02quD/qVUa/iHPZWWceBKhGIsi9u7RKkWqJmJxhOhCTCspeT
npNZ9D6zi5hFIknQeNtvyLX9ng6akY32TYEJEEeujBTQN9Yq6WHQq+MEdcT00oNw
tVdFVONSqAy59Um94K2ZzA1KVQYvz0N01z0SGGhTPKDAH920q9a0LBTsA1hSaJxK
8mcI6bB5rwuFBXUwmmnOlDk4bkET8L9Iy9C6/IREtcU/HkKb/uo5yVYmlgM5oOzP
ucmV0c5tnp1FydjL4MXWvBTUuQ1rdQB7NvzxhyubXU1M9Pgz+/1jCVtYltZVPekv
2/PBRa4JhKP5EPI8P/JDnGGc2sGHIcWCLAhm1NX83iVGKaCCGE/WVO/A6dKllDcz
Fhv/DxNB6VbUrjlW3Tdy2O4x96KPF7x0JSYKXswLLvMeuEVsa2lqsYS8wqJLmbXV
0HjgqQ3VlsuXu7ogsv+WpGP7ZJlOAos/VdqSsHz9xtDECdSo1hUPvG7Yzck++sTs
pC9zSNNev33dAh3LkFeL0It8z9dSFZv4HP/PZd+qX7AYtu33gIsU45+Cu8RSUMK/
AFDbQfymQ1pIT8Ufk3ew7vim1hHhxbgG0WcUXbur3u8b3WYB+yLjxe6qo83ud1c7
Z0j6U5Rhu878v3gvZB9jrDCig5FDx+m/tDFr6FypZY76ogX2glMw00K+qfYTttNK
pqQ3Ze6tCj9h5rGevre+2kBRiIOI0LGW0CaYqK2U2vXot4dm1jetqx0dppBbvCf2
SYgl3DWhr5X45/GfAk2spEKKeGOOah5iXc6Es3bvwJh31AhQcGJqjcPUlYFHISUB
wETaleL5xqZ4S2Ds8kyAyQMqxILZCr0NXHvHPFKz1gXbr6QgfxRYctnb3BgJNgyA
cN87zhHyHBA8EBFekApS/nmgoJhCYQLXPV6oS5a4oLoy/w7AsbF4c/lv9JO6Kxfq
aSWS/mWxbw2o4+plCCuVHAWnEtsUcBtv9QGsJAS7stFjkQsj+Hdabj0gacwYxRwR
O/fOnLiGKHoKkZ30wREZ4dmJoOFVOzy+1hsb5HNBX/ndFThBOyhot1cX1ZASGz+y
PlHDfzey91vwjM0V+Bp5no1EJBTmvQHGPUdkgExLzikS88MhysLJlVYWKUUXQuLC
3cDTOvEUOfews7axs6fU+d60vkDAxuY4XdhWnEkAP6f6toJGRGWQMnA5unOaawAn
pqfQCegCjftrmZY6zCRnEq+wQmFu5G6B9Elr59u80YvWcmLfvrxwshInsdMUQpT9
J4pTJYyhG24E/vBhJta5xVnGrXcgQFpza2COYYKwaRVWexfzfoQ8dCvNY3HN/2v0
TBx8Epo+PWeB0JmVbEn7t6UWA5X1Ey2EBF31RIFPVxd2+TUVhi4sz9NiQt4USfQy
qLbiXdHnWjWZgMdXH/pKb7uhj7JhDUN0+4MmHlVsnbxY/w2WcN03+l3GNNvfyVnG
cRrViwzMJedTSzfWoeU3M76ZfvqX8sDg+7ASzAP2NfGOMxRbgaMISEhO9qIL6PwL
uEXS963EXDjlyIJJSrewnzNqOo7tnuS12UpiDmj9djzCwH+z/RgNze45flM81CXA
7ImE4KDu91ElhVkOjI3z4AbWeHpza96iOgFuz6WiDsS5MoP9uqVoAawJoqDqITT3
nAOzseAED7IZ6t9V7aOXjCtC2REQyHCKlIaQBrgeMef+dl+YGGh6BgfOjjBnwHch
mXdp/hHFCm7E3I2/9PwUrvhFhkjspwzZQ/ccEAd6NftF7ED9+my2yfY0l4x9Z/3m
TpbHt8A3vbsxlJbnk0jMpWl1o1DVQ9/LCed6G3AflMQE/DB0rYOrMW4KPVZmHwVC
FWsLLCSzO/3NBY4okyb4bVeMVQ0DjheO1tTJH4oGQ146pWmG47DD8MDp945AeWh+
BWX46Jo740UK3+wYE3Fe1E292q3uUoU+2JLHMUS/kKxhKYQ1tEMCQQ9zVIAt29D7
eBxC4mlzI9upwDRwYwU7FNl5DcbsW0LfcphT784Kf7lltwSNaeSMOrqAYAFXVGqb
iG7s3pmZuo9Dv4Q+XQ7N/4iFrfRpezcT1/SsrMcYDpmbGKTBgc68TnQqOo2/3Llr
V+Y+5ciMKjCB9SxavPc8iz07LSTvzzbAgEAZxtnyEcLjk7k0PEtMTZ+8OeExVvq1
QeH5Sg2h21R+0KgysPhNjAAZWJ7kJZBWThs1pn9GZYQ3DEjvuLQiTuN1Cq1/7AmD
t9phIVPwDwRPG5j1vxx9hNFK7h9913EhsOeQpeMukmBWE+fYKXp2BCaSPORBd/AR
g0IbXQKJzjXCTrJ/d0pS+heyC3ZrUb5PelWP8J+8mjBsJAghxNyaz4Ejq0BOkSHx
pWP9++V9vKkrb6MXQmORXozWcdMU0VROkGR74AcJdU3tFUbtpUvyO+o8WTxJsv4x
asNK1k1yMxE+T6I0q4rQxcPt+WrMZ22n0ZiDY6rPQFM7x+OBousmg9FllH6+ZfKi
ub7TmxOg2XJrUMZBxAa5U7h8oi9WmJLkcqvBzCXWZaJvVm8N7WklWkbHmocx3+mG
8npSywKx1cujILNm3ROt+mXwfIVN767UCm4CcS0yvoUzbV2ZnZzx4WrETFMZi4CD
+C96oukltfs74bDrLCARBdGExOWHs1zFKPDdWmc4CXTvAok6halljZLPsxqrnTYH
7OqlE0qfIerD1cAB1vjjfaPgu3PqryrQHI4DVbAb8a1GxQc+afn6kk6BZyqUlK3X
yTi0KwF+tWcxFxs9oQhy7MEQtv2en6yjLUlV0lx3Be7JduID6XOXIl/P2sqhIlNa
7MBckWsQNyYjXWYK10ibu2ccZd9GHU5CUONmdv9+qPZkvLkdDT7LScsqb9veBi2C
qxKORJaVQLHYkCD9gN3/eSw58KBvdk/LhLeqQBZfb8p1zhcm3+qYN/qga+79TMIM
TnLwJeLgW5tdbKtVoOnnpqyHo+8ISzm5F5D2K1zwLcx6h93Gae3wCPGbCmA6szYc
wl9rs6WPfsH+ajp7uJTgHbehPka05e6IMc5AnkMAahg2d8zNHvBKgRHnwY0sa+8p
/xW2/jMA0AcVrylAhTbvT0/qN+5fLVfuZxjDPl4CffL6Hv88/P2BzNgw80xAmR8J
RY6CGm689DPh5ILDX1quudjyBOscL1a/tGQmMOd6DpD1M04sNB9Shz7WYDfrAH6Y
QRYbjTa2JeLetgNf4FAj/KB7DSBKQmvNc22DW0t4r7pyke6okF1zVdIYo3pIKWLu
MzKofM4fD7lDBeWqQwGWOXpd7eQO0mOwn8ynpMydD8cKADXdYJGyE/yRujc1nCIO
jGD7HX44PHJUBsGmM7uqxujcZ+pftS5ne++kp3W81/BJr6fXykQamHbmEHCwqTsf
6kz5oWOPRG3ly1uFfQxnjVWo2RR6yl8IIBAiN5jmkirXmAn2ns8GdW4R6kfAjJe4
4V1tyG/c3rBQzC1g1Y1LCes6ZLDVvrNCnGqRIAQxIdc3ROQwH6oMzTCwnhjHWxln
RJ1XIP45wrEjTLs87R1AnbhkdvldSsMWhq+XnUTwNCAY6k5OIQOQt+wwlO33NCWH
B74i1ziWem6YNPeStpmsj9UY0+D+/vWIwR7gP7at5GrZK+ZxScxmIGuQlQAnR9zo
S8AJb+XjmaA0umnbqtRCnUa/m9S5RroacBaBHihyvBK9rTCdD+DVIVMhUUVveKcP
nyojhfIB+lk3XpKyiW+alVVLCakgwQ25PktK1VCJwxXN3LxJbbaol5ul5G3KghIf
i6FSM4H0QM6JVkLCNTqVM7hk+LJ2YJh45o/T29+FnbTnxEoVn92AAMtyRh1rYgby
RuFqCAg7tPZW2iG0nbiYPjFmlyUJ04afthWUlQMn5RBxRvqxQGeH5NoDfUTBZQ3w
ezCJ49BuFhCguc5gMr7xgGm21LrpXBpktQcJK5NyR8q32KNXBML0JSzj4JmeOFRe
7FyQCxvXYenPVm5a/jtTsH/3ohxtoZgoSB4Mb9OFTgrovbo5k4N1tJfgUpPsT/8K
9hekP1mXTUs+v7EvdXrUfbZz6qt/lN1wuO7/hYqmkadIKkRVkYe4RsY8UgKLDNIL
cgnHw6sypsqzGf7kAhMjQKJInBk7X2oZv3eU805FcXO2stPGdep9wLklRrLPBkWm
ZaQVc0CCl5T+yUoD3IcmHQV49OlgVKYUtM5BmvQkcYI+9MONipATGCKiJqadbumt
Yti1p80Nfe3LGmXF63oeM7D8iT53sDhC89PW4cQlurWd34RSLKKzKMh3mvn3EzWI
XlzAXfW6cpuIHu2ySOoq3UnojpPENekpUFn/5/NOAz6XHbFwTjtXKSge8wS4J1ix
el5ebGgIi+sd3q3659zfk/rdGZbpzt8mQLtcNBinDP6fPmw0OIBQ21+gZHdePOMg
BkenUM3mpQo/n5jeyAqWO5L5xPL9Mg3XJQIYDLp4PuV9o7LAW+eimiI5BDZDPKdN
KnSQDtiv28GVJ5zm393jrM/rBMv+0LgTuB1J+Enwrj9IrGXOkNB0UhZ+3p7PA9RQ
5qzq+aFy+o9kdFjqZPZrp5tikoBLKiUPSIEy2NW3ia4axzwpLv/4XwOfyDjb5lw0
jeA06y2zLeHdS1Bat9BxPOn3IchFF0WE8G0/ZUYK6wKotSXH2aQfTVX3lPDpR/rp
tQ6MSygEOkWW/wawGwZxlnpu8SIfvR+muLZTlofNGhJpnWXvT1Ci+ywKxSxNu8CN
UwgjtODu+rxFRTw9iF8qZLYWN+kcEiaCh7Jds0ot+D0xqyp1L2DU53pKl/4s7s63
4RLKTPbMECa0Vx8oh7RFpTOplPKu3KtQl7TBmzT1ZfwSAIrFPrfGz+/DkqnbDgYv
akCohorjpbAlsmOfkTbstF2xHATEtXTLMsMpk3PaA14Bj1Wq5VbFpIg2Ks7m0rcr
tT8NzY8P3iQV1bLgdbYnS4eXLzZM5T3YCKk1k6BoeCyAWNTn1P5Cf0djhiF+C9YC
xdwT0QHTdTFVQI4haryVFIwx91Vh9wjC1+1B05brg4F1uYlFsJDRIBQPbs+ilrbx
mKd8PBXJXxCWhX3wflPe06AgRHZ1w99dEfhZYMrfWq4WieUz4K7fdB6aboOEBNUt
Y2O2rRQIluDuJtk3eVkufuKaQ960f8xWWYV7eqKPATgTeuy4D+NRRkSB7M2oU9bh
D0z+CYwCxqgdSarFXJTAHuVuxGs75twl5UbmqrferPH3T7Kdua21FH2qRNB6I3f/
MM9Igk3dR7TC4YzSlrR9ZKdWjuy3K96cS7ifoTwhuC6bA8BtWsVRRpS36H+2VXuU
RhfVmue4ACbtbcfH75J9ks/84/+Dq8+I/SD+M95bGJHhtFEwiVyJbAhpxCUFKlC5
rXNSaH7bJWW2dfFzBcxyj0x2aEuS1PjMGCAduuqfYOpCrKonpuVcNaUI6KsvS3PR
V+t4JYzFYYQL+RtxnQCLwTHr8WtWA/z2Wl11lOgubE2KbVHw9Ze/lRTDEoAVkR7x
inw/U2PdfuW2f84WrEISTa2V57Q1RSs4tnCZbGOagF1HoRe1ZP3WTzIIAdYwQHz6
Y8h2lWXVnRwsiwSBH2TO/ybFGcX/gFqTC4az809ynPAp9p6FA1i3ZOXNLDxMGhMY
Kb6ryE5OVKcil6DrtEcn0w4qzBflVEuxgyFCJDwDxnP5x51aKK3Td+Ui6wMj0yk6
Z3a+UExs6CZk8rTDpLSqLA9PuJmL8dWv+dKPlgOKcera0P4DKQ9Yo9Tue2rbnccn
ozwfLwAMygFFUTyYUQIYlt+/0gMWgiaQDV034O3MTfIcB+gIi7WHaTWBkTks67OP
+U3l7NPalkdBRCHF/w4+HOFlaBl9qrtA0YeeEsxHE0vClxIlQm031kGBNe3VglfF
q27IxmIyvqX7sPfA+8IppLNdLv2gLuWoozwBlArG0+Pxz033tSxrLme/Da0WcsLq
2hFxb3oqkdv12beDGSkzIsU8uhw59ojR7+bSvFRRsHGMJIKZV4fEX4fnc9OLgdlj
ryj4G3pKd3LuNui5W+yWYxVytorQCtSXV98KR6iLzBU0P/bDXZrKRultoq6U7KJk
Xpe8QKnt6PCgvlBMnuap2Z6iVfP/nxzG4/xCJ2Me9jYenCUwkOgy35+t06bAU9MC
MzVk2RLRdYjULvE4NsyoC8MaIH4pSTuN5dGxfPbVjttbG6lJTjM8jtND6ny5tAh3
eTq68rtizEDKAwfzv3tErVvI/KY0ZjyrB46qxV5kIS66xAOMZg++nCO6YTo0S3Id
D0bPEWVbWll8bp/CFZrcfPLotWKBqhPZoAr7z+DFcDK/EnOhE8Vjb879KV/GSawH
`protect end_protected
