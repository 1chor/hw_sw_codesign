-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
4UNd9QJiAJZFxp04u03jOd52zaKsLlEuDDS738dAP5y4AKCo8M7MVXfc9+SNiMdg
4tfbWm71FvNa+j2g9/lak+wdRJplbFoD5vgcPKhqdVgy+xc1uarBlvhiA6e6oWn0
DDllR0wwpM+pMAu1DBMNyCpryHAOgQgsgd1DQXPtLx8JD1CHKdbMBA==
--pragma protect end_key_block
--pragma protect digest_block
TmkV1EBey3YaFK7vtsP9Akn5kkI=
--pragma protect end_digest_block
--pragma protect data_block
uPawWexzgmsu42LhI5vyv8Bbp2ebGUznyWdiUQWumf+Fxf/EVaKQVIiusy7X5MCJ
KgdfKz7dSe396MR1Cerg07iUgZf9RuIpT/cF7YnemgZsiSil0g93+2mu5yvDZt8Y
POZq7/5OhKzHDVIMlveRqT+e+y+ePvXn2tE6Wks1hDFV3MdHACQ8OfFpclcilxLR
Y8tKn106bwGI0geR8+2JDOe9auijZ90M6Fybu4ge7U1wxAWxasvYcP6GtpoSuzil
HCZ7xeYbwHlvc052SR+2UbXGeb+HCWPJ/UOCm4V9shddR0PRe27sPYQbiLE/N7OV
DhlvIAGqKEXMCst9Fs+bKV0nsl7CISGhmL28FxmPrXyd5U93uUvtedomULtWcsiA
5IdJsu5RBCgosbJSFmdbpY6lzWexNAnvzo6Pfs3rOb9OlHU42YNwRdkk9d2tIlkc
7okGmMX1WDBUbKl/1MNfqMgIBMeIoFgycNn2A+7Gj3MQ21kCiDGjwqINVEOZ/Ja1
0sgd5HjCw+22fPP3jgyEPfF/lVaTTY/lpcFO/be8E685klZphkXivPFgDVnuPwLW
/TM9X3JBIWZIgd1z4O0MHABf/wTWNuBuyZ1UCPQAMyie5lWM/WW+cdRFd8VTPI6a
3hHsOMo3iSe36bhkSqeTW+w2kLiFAcUpV1znr0ph/BuxAZiyzm5K/EGpFRGoCm4o
yJsX4qHRvCcCR2ug1n8xhC6hBzLNjLQgTDHxcpuOoQPjGmoVTSTQCQi1kEJBSCZ6
crHm73xbyx3um1g2jO6WAs3YEFYzeQ0KxUz/odq8G6jMeI0DZ5wb2av7IptFTZiM
V/Vc9ULYFioBjwuie3QCIaZPOGZ04RlUiB2ei1qX9Br5ufPO/0whjwebvJyMUKXU
O3IOzUqaUJra/tUpydP/GsHTEaFXvdC/qU/3+CghO0g0JHdK5I0NMnsygqwOrA+f
vBrblL+DdVNAbbXKay6PKls6muHF8NpjhRyFEhtD92rgrnCYr9PNTFpr6JO7L4QU
N3wLEeCu6yjDUIEVDcKJNwchRnYqZGohTV0BGV29Q/H1vU1IttAeKIEqSR5QkWIM
Ipnfm9E+f8izLAK9YXAbjns2rkdE55X0fR+mttfCR///Eo4q4f+asrlSPDGtm8av
oHeXX+3oqi6Rq7HsI9nUHEhUk6Tq7MAnd+HAWo1Nx1pwiuPLzYJo2yq3/bf/W8B/
RGni66d4Akwn+0Q+R0VBNQx9KKIzP129PvO5VxkkAlOvL15jp4jkQUuKziRAVSsq
b2OIylwqQ2cyzQUZs9SMXLmCL5UbQ6+t4LGIdr5g/ATzFwHlkVyo2H/xPhsSIvMD
lcg1saCVN4HTA5XZMT5fyYp9SWqjvzgTnQXc3evYnNgfEiA9c/xj2nb2B/8F2h8f
eTxjQGLq5H8SBPAJIbYHVFutGMgwrfatyt3H4L8AuBnfXl4T68N3IuMdGjIxZUJL
Y7tsmCmmnKwjKvlBCkVjO4UAAkWIgN8yAIVoJAGRQGcrfOzw+38II2AB6GQpDMBo
U9bjYe2zfudfchcHsPMo7jlt3Mv3Mz2rOJRSp0Ro+BVydPqbz1HLrDkwghopiFUc
pA62cLSOTP1rrLBgtsret4fn3SX3Q0ernzsSawfuPzksgaWqCrsX6Qtz5kfGQVYM
n+OuV3NXl3CT/XWAB1AXLCtlNPP6MPqsEpwodmF/ZOEXKZacS83GnoVLcMDi1sKL
zCEBT8PgUWx/59XFyeL+IR0N+nqNUCURQxN9ncDgJrVuH9h1b8XZr3EN/GtyVPWZ
gJ6GYlqMaRkMArCmJr7RDSPQx2rkaIpYF7kY72LIjarxqttStv5jIKQ03O0R49IM
hMIndKcrTOaEzcCZTU7zX8Qj36WsqoQyFGMDYT9kmwGCBuRnbe6lDMM/fFobVMdg
CkJP/y6hmDBCj5RYaNqsAQXxuD8MagmuDeq0h3ZzfsyX4xZ3LmOceNXizkyRdtcc
PmFB42Bes5MfU2UdTYq3k9YPa4tP4SK2RRPIUcinVHX3qKdczss2wWiVjXC/bUAa
vPlEDW9I1TEosPbRvb3001WN4DtFwsjkqt/Zzt8L42r9TcXs6ixcWWP+7SWHIRj9
45eWtS1UQXHl4v45yOZDCh06Txl49kLR5hz4GKgg6tnxYxIcNiMODa87tPRamnt0
3V3M++aDJeovEKB6HLpPuU2H/V0QxF1XEu2Zo2oMUnZ/NOwLWPm/v/9iHVKsSjqP
OLD3rx1oY5Rw0la2Ud5Q/7tbBXXtMNf8Px5JZz2WrBSbdjNM9z0gUecHVOujpMFF
luzw7cguHuewyIMTaDq1rlf4yMlx4KEqA6e+L4sbq8vaticgVd0dJzJaW9OKDpSp
+BK+GJYubFKFhUwQoMldE8/1auFX7AmB/WDRusJpC4qJ9J/MJ1Bz2XuRq8obeBVr
223XOSTsUvD1V8o7N2kTMolHsb0iMiopF+pdx6v6KV92niyaAkeeLm/wGsuQf/UM
+eOJcdDfme85FDhUdGorsc0inVgRZAFifQOuu7v2qqPuIE7JwxQrsa+cbKw0o7D1
mFKdt1vfcuimPxyGHjVd/QgClcjc9EaW/hllRQ7GqOZ6gcsonQvDgMk8FcqyADIl
d2zgQa0pjkn3k41EaW3C/ikPu1/R64ZXwG/r5C5oeMBx+hVXvlBKw3yhQfusW1dj
jIpH7B5HC4k1UynWV6rLSfF4XRRYuZ493iA6E+dW+8objz3IwZWKxgjdEEmL7MsN
htJEU/y/mjnuqjBzaOPAbZVgXaAYk05Yc6UQyLN28QUnojRL/osHqcJ6ruFk8Vbo
JC7QV2ElcL7/CtltO3C2hLbPBsoIM8KFyZsryW7NTYwIqq9WJG+LXqZFuvNLUDap
ro1hxUCqGL33b1Mxizpmzt7QvJJgDGwb9u2jn88y9UqaOJZT91cM1LNBazpm/952
eCwEh4AVdkTs64Ne7kr/gT9wZvO7gbk7zOVMsmXcsFOnH9hIIGaqfwHeF8taw6cJ
BrxhrWqP3PaF4qme6fy8zpK0Q9w5EUB7euy/6Qn8gjku09+XALoz5vnjHnebKBWI
VQZmnD1Dmdoogx2BvvcjXpTfSOPE9sPzO4paYxKW1jxil6w/KJ6fiF7qUJlMLxa1
e+Pc/63tfQbPWzbnW157qvnFjIPHVg1ysta8v2bwERWNkZ1lqU83yIQKFDHkHmKA
fw68/x/a0ABjdeqcfjEW3bwmsnLix33UnuVaGHQUHCuf/WinyA1u98cUwxlJ4aO9
ZQNNrRM7hfXMBl36eNFv6pkzlveL84ggoA0gZr7akriHMfK6HtdkRSt9o2yYclAj
HciB9BSL93YSjkqIJRbUQ3Q1RjWE76z6miYAuo7hVph4wqa3jFuyzXI1K3WSMOLY
uY+81Lq4GfZjhDUq/sVo6yG8j2GOhymTotRSU6IjQSpEZbbiUHJJngXVmCmuv0If
bHm/LMUfNrRl1hXB6rVv85tkD6ChvigsIZhKVKyJFTj4tsxN1jnxsOl+BKZIaGAa
4w1NSQKpsHgKB4a0279GkaQrE+HYldCCu86Q1suUKoyBFrUo0DVR9cOxCiBgW3un
5nFvTXGS+EYH3a4Vux6skSZNVYw/ZNojjE82EEl1PcAtfDHbxTGH5XUsrs0HYKfC
2eL6EAgWGGOaBprK2fZRhd/WB9IgyeD0ZXxBvpbYkAZ360vrP/xj5NMymNEfhJXJ
sIvHVwqaoCHpaViirNgXI1vW814RO8S40i/DVVbjM2bJgwYz1OraDs5wKG7eWu48
t7RtztGygT3zODDGzgVoS7TCTMLv/tioBXgIQMzdoUaHB5yWCPSW2KRfc8WkG5KJ
F0aTIzIWPyx4SLFmRJ8XxFpx6lMyZcOdmOko97RqPIJIxQ4ztRDfGe+Cx4ZhypsI
5S8VaSr5EhmrdqE9RMgfQcUYHCW6SJWisDHXnoPOGHnOZfmgs3dIiT5Cs/f7+HDz
6naWREaoNN77sqGvRbA3nYBnxFDe1QmO5LJ8Jc0GSP6bL2DRcISDFD4vAtVpB1b3
+kK7rJm1QKVNXc96LKUZ8g34vNczfmTmMl2qBa/XEJIw3Xtt3mze+5uz3xqb59qM
vB3p5sKBNJLI4QOZKTD9BXWCPd+WexEBvIS4ZS47bKBAhn9w3RHNSBvvHLXGTxC5
BfxTKGXM696gewMpzI5Cj2C6JTT2BAtfXpKD165S4JdTZoTY7bZ3r5d2yzkFTyXt
GN89aJwalJFqGXDhVjLBZM4QGTVQIaws96qWNyz/PkLBFhNoU/ILtwZnMRlaannH
8heuj0nKsKMyyYLnHzWPqFcMmNE01X+em/qbkA8ixhDMsXhXGInKlFE75Gcopug8
J1rlIK18J1kNm8k5rnMOYr6tA4YDfqkd+h+/yQvPSWa2TSwa81GppcXy7UoCXfsD
3kgV/DGTLGBDOszU3fSyD9KHehNBCpunCZet1WomxPyXNegZULgUjhj2vZzs9K/2
osPBBsbQurE/uz5UMN6rAgufJU1FNoQDveQvOrNGLDBlo0ddUUJZiurRN43x5XWX
nKkEKGeeyiZq4B+OoeT/eXjsvF6+l7t973MjDGdpw4aKjngpmYeZ13Tha/spSz1K
m3BOcnGGMkR7Q7+gmJE3JSZ/d5qyccvGyeyn+V2Dm162YZwnG8Nvys5U/DCK95mG
FddEJpVX5S7E4yGlPgQ98AgtRYzkN87+AM1Ow62mU7c/dM3TqwzwYUGfQNGQUnmM
Uh3Iz6JUWPpmjeRlFdCc0V85YNjnFoMpN+9NxUxLuHt3N70mkL0EydL5rit2Vr99
K65A3zUHiJH6kZ84Woo4s/CnETg1MloGACcwMru3CLZ/FZ1kki1J20w1SzXbmUuI
lpfy6AYpf6majE6r51U+xWcf/ZyxKPGUFAO1ibpENNLJVZ9VTBg9uyWiLTpWxQf0
UmX+lEXdmu7TlIsGKIyKxQmmq0wD4cBFLynbWGLEUIWzO1uTEZMSfcoA9wFEqvTS
9mlE4CihsWlt7hiFshINvb+Lf0OrUpEhBBhtkHoUeor+7sfOE3NJiI3qrlwl27N1
K4nE61PZh67vfNtiPRcIJFHeGuTDjQZppieJMeNj5XBalzhyxSP94LD1vUu9t5uA
eJFmvC2hkvua6WTNBl4Ug6AmXcrapjyujK9kyPlyxMe9442MX3Moe4TScH3fa1W8
L+Aa4X8lNpeM+KlRQym19eYDeoXEPslWOmr1tvzOuD4LpYYb5jjDNkna+OE16tYo
k6FR5/c/El8ILfHVWDa19nrHd9EhniiMEjW3ixGVZ93j4y/92CF2gXnvarB4oMqq
Yk1LNntpA884Hkkz68ZQUypi8PXT2Xxol2l5gG/IKOwvXIzIJTbqsJN/cT1kYmAf
lHYpbn8j+tHl6T+el5GK28KKQ+ot97pK41NsDrh/d3ykVzhfSd5+5PHwzIHREmBV
g7TSIlzP9nqQoJE0RvQxPWJ5zb5bFIilPhLKF1/5AwHsi9yhdZHvDP5Dhvketihc
FFf169QBNQaKuKsXRco/tbv0W+Rp44mybclW6vBXXHBG8jIkPkdupSOoZjLz0a9D
9tm0nyOZp5CdxMHdTUWK6500r6YGMulR4ifMJ+veV4He+x+nIus2OKra++fv63wc
FmMHS6IDvM0XD+Wp6wSl3CpLTGK64fZ0AO+NmpYCMlvLd9Chhn2Kuac9OdaLTQVC
IpVLsW/0HjVetw54n1N1Z1JHAsQ5Ui2H3H7HKPGmymCL55LvMPqzh5ZpFS9kjQlq
foh9DZ+y9cXyMD54CcM+0K9E+xfNYAK1PKJvS2+32qxs32hxU314fsbEfAg4BBsx
49fJH3AkZg7BXMSYyQ2fgHzxut3laYRC+m1IF5SHDRE487CNyO4Co0e+c867RadJ
QDKSV9Vs2edKd1q8sOGOtbCtK0D8+A9rvtvU5Rz+D4k9+N7eK/YIthb89grodPJC
jMcuojaOAQyfvti5V9nzoSJZIpPDFuIOsAskhPfOCBxWrp4yiteadUyxlXSb/nAR
r93dRbgsvxtHOIgfbn4JLS+0sdGe16qtj6RYuxWEYrWkFZ2tVbiM1M95vIpRSdlf
fiPP9sZ9FQfw6/YJJsyv/gZlya3LCHj+c34TaOL65gtF8MOAGzhxP+93gktyy2/d
6T3Ek3Z/FG0+aLjGF8/bXxkyZVUK2MqrlnYfT6fssjojfXDvK2MVeeLuPzQ+z+am
8sQiEMIrcQFrH2mG6kF7BJIL/9n8pFzo7TzwjLgl0G2PSDz9kC0QTfSR4prxj4Un
76jkniiF+y/QISgO0fAUg4kTQKWT32Wt+4JcqPgkhZnfAd46/vWgmAGsSLiH7IF3
i+pDSrEM/qQI/3jtXK+rYB+IMmtGte2ZKKyB1EHgmu1VWc0JyBRmDWoLgAhTfJBi
ZqajsZMwwZgtcHpJojW3gdzfFvz4XXoq/n1YSDfa5O3+FWyuCXS4cPVMh7GFvr9Z
yYaas4Nah9YRK2FdGXkZFseNL+d78HDv48YonhEdjzdNTaTGebx7z323ky6ieuv8
MGn4JNuVJWdee5DPqU2Eiqzk2JA8A3A+WRl94hU06zbNpEdEaUisvHeZgnCtkGOM
UIdmE+dStPLeVpKhh6eukcH3hGbv9+fpzM8S4hyhh+KX37VmT/J7gpFKLDfMbNDn
PNlTLzVbUru8s11nBKef7KPkP29kPDHq5BMesI0CXoP6R1rxyF8FDaCjvZ2rX6DN
zOzTttplrGcFY5XFQbGhiZVJkDeDcE7j5SoBZa1lmojrOgAyKZCRw1cBt8ml+imw
qPCuR41Tka7ZUMS12YyeW64zyfJ1P9q9EmM4h8pfeHRQdk+gOCZzJZHBsAJf9ewn
Y4xo62F+OSTNdG1kUkirnMugQeELPAD8MhLrxQ0V8qerW+lzYkb5QkMRMYIin344
KjgzeqaAXIundockh2zW6WDZsprFPQUGusvgNpb8uPYj//dzSFG0J5s8UqazN5Sr
eHq24dc7nkelWm5qWk6PPcUMLzFo0ExZtFOflxuW94VZ96t9CK6f0uIRbj6Vhlah
nBseiALMPmHT9tsdUre47WqwAdERwG75pegMFZI+kB9IvcW2Vevxyn6FTcnb4XfM
/8GudnwzW4+szaWnnK2MRjzPLhc9aWV4/G38gABcpZO2STwu0PwaKGqBg1VG82r7
j1W1xal4lQRX3leYxpBE+tNxMx42xHN7iZcDKIIHP5gVdOiFSm8UMQuM+uTMOhSo
/tmEvdk+i1idpsAV0YmtKcUOjTYg1kysCVslwSoo5uekZbCJdy21IuhlhdQ8uoBw
3Y5pRzR2v7bzCqF5asq4C3jBlAhAJKaiLirrJtSSOwO29zxMdn9p3xrQD8fp15mb
MxIOmzuCuRItbbwh/YYwyJtWA/aJCdkX70x3A31CrpQhBDhkyJmlfU67ckxsKAUO
lTBhloGc2Tz0z/JfF40PTOs4FBphssPkR1J9R9UZ9xdWjQPGUFzRV6qN6ZxNuM3X
F6giT7ZHJNJf/Uj5QhtmVqQowW+78T6ARL8c/iyTza3Dpxmoblr2JNpAfJ9wJosy
XCi/snLmLjF5MQAUt4mzyG8xQ3B2I8naSxwLU9dzT31/pDDGIQpdJbtsD3JXrL9D
ywF8p/FkpSdK+sgNMh+W98jVqr3LVgOAWIP1bHvdRaLzCFhkavxBMPpz5xrMjatF
yZPyOJty9EISlb2Zl2XmPGcL8q3P0eatD33aNSEPJYKo2fh7TMuGv1agpjFk7woQ
ohblCk3/xsjiX2I9KAHC94NZ8IsW0iNylfSgkVs9ItMF8RVsKXWM4M74go/zzlic
EL4f6zlTxabNdKGzRhYqa6MEtmkTW5raEytyr2YwQHhzj0tH72Nl1WFjH9gmeTBv
2K/hkJZTBUuL4syAjt4UVn9rDgJvhrRZRThtzx5vxnj+1X7ipzSPR5eIYlkRFLY9
3s5qIOLap+uwVt/DTiXuRa6JQY60gNkUvYcPrwWO1zkY+a/58B+pxSkYsXeAoIKT
IbIBGkYXTyuZaThVV/e4qI2WAzU+GIk3VCnxBPYelNshKTZFzlXMqUJQbmj/PL5F
RdijICObt+NG28kkwxwUz07ld9QqKeCB/Vt5ASpUVoQxNGcQCrF9eAH+QFmds7dN
tYVQW6XvQcFm62xgoy0+zjZYE5LZbIGJDN30qK+DWaEF9HHiQxKhASIY5m3LQupG
VHtFfVF5ScXYQ3akT5E3aZtPpW4p930z20q8Udsq5fAm9vH5pXL2+s+f8mkZ7Bdx
/aQKqsmxODs1F69Q2nwRzuO6BAdUfixL63ly0itFWTYT8UlYSgGQKgmdTXvr1amY
oLGhlO8edGkEdzkrAsD6J1YU/qTNL2kiqPOcj7Gs6PG/7ivzv5UWPWZPhX+lwuPz
id8TCX5wdAk1DYCcycvFilBrivDxpYd5pak9iWZKnO8Ypum3l3boZO3KNEDr6Uub
xS+HlsLpNBV/2Fk6oje+8FCnopVDu0JYz99/prVgc555Yky3PF7TM6dsYbUbLChF
j6QJzXmFfPJZJPFZQMiEpP/ABmFiQCfS/eqsVx0JT+krn9NOp5v7tA059epvr51c
5oRkxaA9KCsE7ey0ydtr8+plsy9ptr/v7TgJUJfCdzHNNbGEEyw+eMKXU4P4rJnp
qbZFGqV6LD+DRWUCCCw9xwo8B2EIo1f0oRB06GLzDVZF5kiKV5Gl57quiR5caMwY
FE6SkVJFZvyOl2+VG+JCnABq+7zC3QnYSDuhVafyoXE13ra79oKKx7QQ3+cgSJZM
EQvGE7UuMw0RdxhctZ3o4ueblIrnKwE4MsMmTgwNLCBBOyAuLlTjU91K8Rbox74q
zZJ7n+cMQ0QnJxHEdHLu9bkTUPG7IuqEdpBqLSFFcps7vtHV6DG5mCL8KPquUlsu
I2dk0rJlk0ewzUd3ro5XjrHSOvaZ+IspVD1564auTez4x5ZcSRM7nb6v03mplLvq
Ye5qqXDEKqk5h2XCltO55dUUh17xMilNDvDZujFAFksfMSYZPgQhdGMnVZg8YZLL
+B6IOB15ClX/ODjNnF+1NejeqGStol5eZxzWLKw9hZVzL8amjAZrjnvxmGDzJtS/
1U3DlMe3hAh6mOQvAopcaYqq9jsu1vxhNXH3Zx6I90bT6VrcdDMFmI/sUdaYQ0l7
qUXiZXW3JXglTPzOKSFNb8eNSdUz7tog0scTugrZ7cTWRE3bik2KTT5FALtwOOJ2
BqNmwY92zsv/Tdgs1Y2ZuvePSDDv8enfq0WMDK6eXfVGW73cebMonAh2ugd08EjG
91v3OE3Dd1dq77k5sQUd6J1gYOngDQ1JRqM4FqAAO+WFcU6HxY8zZ0hs6c0uMSdW
0bDunFdEWsA/GP+MOjC172Pww6LT6QVSKLX9ECBGSCbzI0uOwYuFH3tSuWCGb7jf
PgD2W9RIyUuv9VeaUR44m3Go5+j4DyCFAMYyJ73tJT5GuN2fkPURpfmBJAYt/Gyx
ZGc3vYqoPJz0TfQJI5vui9fWQX6vzNQKb2gZJFhkB5pfkVGBQPGAVo7Kbv7/0XcJ
lXsD+XNxx2SPVehbOrYPLQIqWgIf2VWQ4g6EuegKMacfGi4lV+kWDSg8M1hG0WtX
fbf+QSNueo7ntMqF1S14+KZ8BNGhawShWF62ruv6nbjSW03cyAYAVoBpNamJsHPi
LFD86EFGdbHeCAJKP9yDI5dVB5WnLIcWpYRMylPcqiYFershpyLNvjWN5Gs2nElp
BnsueGoUjYNhM0zAWoctZ2aIOx940lEfBLOQ4EAmgQLH12KKId9/iJp6CpOL07N2
QrVHB14Q+3MS9o8YNYjdQFuR14MpLY6HUBptQkY8tOzg904Xk/3dvziP7GWUbc9t
6v2ng3acQhroamIPh24KGum/StRPXSwGn0RJCAnWRMcztULT5HjRTh5vQ261nuYf
wKNUHhzUCfgM1/qol2Nymy2T7WngJkZfZSha5waRWgE9MBCLOTd8KMVaab7ItDNU
HTJintWGIWXzCsrowFxHRnMmyCZdYLM1B2dd7HLxsZ59rMuyCCRayqiyQcWZKvXW
6R+JBNrQez8aJPeTQx8cT2AEtl5W15B2M1pDdUC1y6uz93FPVCVdNg99chYiozjn
Szsg2YGD94eMwofAkJqJr8s5r74JPvjrGFBEwV78x6LZVXEn+Cq8/Fo5vY3teX7C
8fZvfdwTYcH16YEGvUflPMSCrLO62aIloExR0VpsNG/2i3XrdK/0z2l902YuU8kM
Lf0uy+EW1RbjksNF0UhOb2pdQiz02VSC8k70Y2dIwhGVJKdd5KEQZFivwOoDOMTf
g7A2NkVeZzUlX7UwUfCYQHOwjyiOfE+uJEZxUXrkGEzeQIEMPvl9JbZ1/a1f0wlk
Luxs8e17mwycWvUMJ7JyKND8Ir67+/KMAp9FXA2QzcgXjmMvo0Wttrx+SsSLKXCO
j1islQ7gIZQ2hUS1dbgVx8gInpaohQ8gKnevzpxTJr/+P3GNVoP2rWiBoeEPEYyk
fa8MLzcftTfSF4Hqz5p/3s8eaxI7YrX5iXb32hhcIEi3Y9+NBs4UOF61LjIHs4qf
ORh3eYxVqepy2Z+cZOcPw2CsWdGZwxVZzgsC24rmmX0dhmrtE8gabRy2xJws0Flh
8TDBrGlDQ3ZR7mT+74DA1uEITb0XTKFWxKAN8EIyXUyZJwdB7VVIr2mbT9UOp9wD
222H58p6pGSSMI5vZo1+YruqQ49Acjnde3oJep/9AqnzbfAQgXa7gZV6l6usqQMg
vtZDgQvX2cd49TTfn3Jf/a98wAf1ZFdvVBzq2+q8JUNV6YdTBO9lRyD9PWwF8QdW
HMaALTNqwcHGQXT5nMZ42g2OS8olipl9DobZxw1+dJGzag0MRgyXkiub56zDTM+i
UsKJ8giMFcO0oBM1MzoYUs+z1vFhCVliHVcLLY1BAd+LAJTnYHX/Zxk+uDHoDSVG
KeX7FQ0KcQHmudwhnIBFdXqK9ta+xx0YMfrWsvKAQ8QvNv8qtggtB051MgmMDGS8
MBTaoObRlRCgUr6VIh78z0ODpHqnmd9UUmcQAVawefelUwiST2d8JYL/LHIKNvGX
107vPI77FnRxCXrHNTm5vppt1bvlNF5c0LW/idlD8DTNr+AAzTCuwLBt0bC/rFIm
oNVNHIGa9m8Lbz9XvrXwcYqn5Vplo/sO02fMI03phcmZswalPHNqU94kXbSuSz3G
WVOGBtx6NIrrTlXSEXXTKNjIzOoZz1uOSfIK56LMwE+CoPj0i/H+vfj6Q/UogAPm
Vv4OkLo5Ylaso7g5f2tQgWOE26ZpoyrnI8xceqocf6ZtKOGDzLEQKFT6dvzN8kXX
6R3n8lHl1XYKa7JvFkgjk3HxxjHA+DxvoCdknL/jPbtzbKV1sxErupTygDYdEuDG
vk3YUsXGcKNQ8yXz2BYv9wHqzNXKALazfAS9B0/0M7IuGCwYo7dmUOdA6562zGBk
OPlOKtBb+z2Od89nVgHtOnX1NH+YI3s8FLb/5BsRpEErZP6+3vTR850L+0eW/ry4
ucW6h21F7HCTn52Y9qFEItC0dccF3BuHKneXzu7qQeSK3XA8hinUs/GWrD7V1ZnV
Gvm1KlqOjMR/azULZUlkynSluFxrRlwFsnDbtyxVvAPhHr553r1TA6SlBFMiSWSl
wpUGVAr669P02mUtlZgdpnJ7wJxaDAnl3S9ripUIpzu3dstQTsvTN4cOirApAz9s
fTA8JJwFtUJO+a/gYzCBSGlVGbMc4IFOcp4EOOlldnJkyx93xgytft56auj3pAtS
b7rYYPSfR9OaO1zAcOiNKMV9z1wLmGMYH+Gt7sOMNZQ0JprbCcFAJU6+WSUzMFpy
mpS4gKZxv+FqPasK7UI2+2shul73FRTqRnH1PS2ID8KqUeiqQwY5y90j1fLw6FX4
DhMzTaUuG2AIA3uZQ3JNv2tgH0X4xm0kTTcdPmWc0+2HqdG0Atjnoc+Ys7o816ED
nm1wItnC2EAenU8CL2ZaNC7tacWM0/99/NT8EIbj0eG9QyPCQF2PENF5zUwpFDqP
ZN67CeevU0/oJHZmpJxCcnHw0blwlOvzcwZu+te9p3IX4ierAHkryttjhXSo4JH8
krJl06lv3XgV2XKc7g+KLsBk7jccxQbIP0c5MYtY53O5MLelVbJiKSirUimbuGVf
d1fXyhb3waLdcQLDlDS0TTXbiIQp3YqBNSjiJwV96+rgZGrtVVhxTxzt7WwlJYhd
1E+YHczau03OFSZElHu1F9vPm2KOybCllOQYAnuKKqzmX+De0odhj4Hklx9fN06x
NPuGugn7KoIIGI3GWPrm7Gqwshv2iRcUvVG2h12vtPrkADr0JCr1Ey9wj+ZI+bvR
sCuCG0MFXvxDcaJztNxfBSDU6P5sG48kvKDvpP8qT7QtSaIF5NCRHNNbP4Bc7KxX
R/7Awon/h1JtftFJc8RJMpR1sI7P5O/bvwVla0xP+LmFpUAseDf9t/s8gPObhZy1
s/qSAoPeibnj6S6D+Oi+DLwMbFG0cWProGCr61KeVY3ZiKUd9chq6fi829V8BNkR
f87t9Yf1F+X7brcvGOwtwPs9Y0c+Sob9F4/IaiK85q8vlqIHMKw60GWSugkN6/ct
VPUIDtn4X1hFvvZ4bsDWzDY5g4X/WDRMN/Jl9DR2so9WD6Y8kNN/s/lOasHoLAbK
3RAGtwCNcMORFJjYSOc6V7u8klDcZEjuF5WIEBphxtEjEvUA3iDwiI4Fu6mmWe2g
MZ63bUuEpEO/aEulYnKLxL2TcNqVqf8qHj2FRpl5H3dOZgEgoPBBulBdKxiieL3c
aM24wHvOKUS1e6QnkuidMV9Mg2eTAa9A+UVn+eKueaXPWCL2F2nlUQJpXclewXit
q0TucI4uvYF7DtHOC3B2F2iGMqULTI1q7FSDl2ku7x4maO0CNrkgX3gK5u9A/+4z
xlFp48Ez5RwHqPVOEpa2/ItQP65dY9b34hBhIjqJ+aSDDpEg914Ciz7tyfLpAsat
ZlLZgFiRnHd+lxVGjHEdBi095u6VpLZifoXrst4O+l7T9e/KfYrxUDKP8S6Nutcl
asIy6EmayNW+uHvBNe268VytGzHly5wzwzrDQb3y3XrfAksYufXNgtyZxhLULx6e
jbBsVL7+rTckYiQ+HYxI7bkPkIooGrwMdfsGFAK4WhqjYgALIehXLpfvuY9xogF4
4MSx2f0mojc+SWypP3mDs+sdjLv0k4JBTmHpOuV7SaJ1Z+XZ89S4qj2xP+tbHlYS
9CQpQvfL0WpEveepPmf03j32j6c6s29dLnAj4OIhrc8OC4PPm93sugpxNQlF/3oJ
xXHCGS0NJ8PVgsUo3N3ZmsdtwTdLntMG9ivyzSx9IXN3/4euz8JY49Vw+2yYrS55
sCtz8GoNJghwX1Y6TkplRIz0SkyjDx7U4t7ilxLFaWoR2/prh6i/U8C0h9CptpDZ
+G5pigAWKbQaDa6zEQ+IRp5BjY2hAHjB3371D4FZrHpbkrYHq1xGLsdR0Q8k5rn8
gCRG/ZNhDxxgEF0O384QV8l7Hg4nGnwmMHUbD/6HBrBJPuUILY4KjsMbsNlkw/jB
2+V/ZkXIV7LaEl6tlp6Tb0p05T3gvMaUp+eoFIXbfwC8sZg1/S5JzIZ9ELdHjArR
tHLwI7IKXksC99nBco0s1pEGuG3e0ZH5Gj7b+4oEvRPkSzQmkwzPMTItOYc4yjTW
nZMhBPvM574Yza2BZ1W0DFGAUWpUTfV3PBBqEDDw8LS7MiCPuKYqgHSVKlAGBEPO
eAIELMZoqKwN4gYCTqcgWeXXMMr8LvOCs0SdfVP0Ra9+nOdEiLOSB4vgBuZtqsTw
0y3ZTBtRaA4cj8FGVMt5PfMxVVXN6oNisCFh5vEyQS7aDFW8NMXtBguSbCsTN4uv
U4A/fA7cMZj+uleUA2mCwSp2KobtOPd7GoogOxv9iGCe5YdootTOj28JlgdbUx8z
VFS/Z6n81jtGhuZMFtXvwxva65+9TGP7X97aoPx6lbP0aZkK/KemI+Va6zpqPi/K
Y25wYRfr4E6yGOG9uN8XKfbxjyrFUAbXztOO8deHc5v5SIHgNZtI9Soh25TuWZYT
TeNn9Apr+oiGVy/M0SxvrtQUtBud4EbsHzR6wP7TFKBALReNz9grgSAR8SjaNvvy
u3I6K3B/5jva1EZfK/unFtgLk4MaPsmo700s40/LOrS29kcYi6qjXeMvJXMfwYkF
qcMftRL20BDzLwJJs9LZiVDkZlrhUDhWfXyEg9ZNUemRuHRKVcptNQz/y4mPkIKp
c7K3eBgMpJ1RUZ+jER2pSFOA6+QNcoTDYy6apIPmH3KjpxFHDljuW00XcMdQ/fRT
/hgNY7CyxSHX4qLahSb5afuHFb4c72nyk/Z8motWWo8oK3quG2/GnNTbEu9ttpYQ
7Z1tEH0WyouisOwL/u1PJNsaR/jrt4rVkgKISi83+JS3M+nM/0AtJTodCsRItnn8
gZXBPNZjtZKE0IB619m1k7TnrfZyR79mtgA24UUNllLfwfI5ZBmcao6xnmuCw7vR
rncuBBUBRJexJIdSDm2tViWYN+twbRGuClDfvoFD9NnX/2Z0dmCj15qlnnWm7IzD
k2FSWP8fKVR9gWY/e3o2xtyBNUS3V+2sASGDFnKNiiA+B56IbC41qsnkObwpWNMj
7k26JAFVB6bOiSk/0qvbclYFz/IX+zuez9YcCbkS/+dzA4+2ZLplD2naPcdlw0Oa
WLMhJVPHR0mktFWsTBtO0yga7zVFsjBAJg1eb2STdz4LJvX1TVyEBGcrnPbHswgp
kQIFXE5RUQxglkiwhGrsQZMIaA/4k2Clo5eZwPLHy1ETLEcJmRpKXksmpEkoJK15
EOtQ1rdMTg8zwWrjr32OcCXbMCY/Jh1A/4HLB4fl6xV8xalfo03calotwJOdXHTK
JQNixvOx/mQUQE1xDVeMsY4snjrjYZ3YR+YtbqVrzTOBw4clEKrlh6O8rkCUwMZy
vkNueltNX5PgkRo0IPBcxsqft2wG0NT9iJgio8Ber++Up+n4DSUXBBzb/GI98L0H
ZD2cjZxc519m9HGoUq40vovZbadxp254p9kKMsO7C5Xha3mbX5gtqO41PN8pQze5
cXm7DBEzicdlD/pjqyCstuAxnbkRvr7wdOIsBnazt0BFMlSLRsmjXtcYzXjPrSKg
DUgzfjIlBpoaMvwxAZhakuJDaopMIQBMo+p9i8jH4UtzHv3YTpuxGdK/aVP9XHMx
AeA15PDtj9rqNjiZYJBB9e82zVxY3iAH31rrWKblsL36eZuQ0ILV82yoy02vW8cu
ofzXTRTY16yJAafzA9lTfkoLLK97890+EjEa/CUVFJvHqfc/VTR/5RrU/RRGe7a/
AuIPWtpAusALsKJCHNQFxgHmoubMLXkGaBhNq9XT4B8FvmJ9LZzNeRG1E1xr11zO
xevkSeE5ZVWgEBZlqntRZeN4wRdVIsliHav/Auu1Lh69azCRA1xM+8u6ZCl/PFj5
4tLROtlmZgrvcnMLYIztC8zdyvNY2r7HurgrQ4Gce9CKaPgBEYNO/jGyijfmY5HM
6ged7+kkeJ7sCND6Zc/S9NDwNBw2vfRKyxqkgfxe+hORLdRMxOBu/W6SoDYJ0ArR
sj1lWlv41Hqfhd4UpEwxvKVX5RH0SdB0mwODvQ9t09oIy58kkRVfbk14FrHn4f1z
Jcr43PPDxOSj1LSr/UiV36eiwCBaq0XTbgIo8qCgW+mA18eVIH5vTS9qCt8KkLQQ
zSndAhZJmuP+LkSbRUn6S8Q+KALR3METOdHQW5UJ9RAKpYw5+R4oic3a2FXo+s9/
Mb4dt3Gj/3qd15id0Ul0W70Oxoke14+kWoPl2UfQ2LybBUv30CflTsZUxjhORw+b
dNcSLwPYX0hEzm7Ioc24fBarRA74+fcPC5I8xInAUQ2EHOy0BSpM0IUNhDPron2w
4VVjZukPM4Bm2HpPGiMj3JqzOr/k0gi4iniOxbP8nk+MNsRe9HQum9ykkaKw+lPv
jech8ewX5fYo4JzGS43o2E5Q9wtPrQxBpTgWxdqTAIVpVbfe18dsTfDvi8kl3gLz
G3kH9L+jVPI3d/ISc7c8FIm3D+oqzLgYqxfpgIPKMjCjWUEuY33K41nyJaTBpRrO
t1EEYcPNEbkJd+2dMEhDlQgzK6bgnA5JUiE0MnY7XTWCTacKXSVBAQ+JMNvUWGB8
jUUUMitVSMDTl0pkC9uv6snQT9WbOpzq4pVurfzZmozvofgmUc/iCPnVGMkG8shd
CBb7VycgHiKAHpWtX/JoIYY5fV3lHpbYnr++iptARLklTuFx2eaWEyUZW0w2UI6F
uhFN2bkRvNlXQ3R9zhgv2sLRxXFeZ/v7fjGs3w6/QmPu8ZBRqIN/hupx7S0c/eHL
Nlb8y1jf/JumWw056qYaitZ1VJn0txvYQ8+o8RVB8MoiRR/eqYvrW5jb5KtKX12t
bbSXJYgYj5qOJIcnxCU4DFsvKHhWjyG866/U3T96bsxFP7nxQDj6x4KjCCo0fzw2
vpot915TzU9ugtoD5KlQDRiQFUX6qSrR8NVlUqjyAxnfF+ikCDj7NsizPDq3zS9A
EwBN87b0ig0KPGS0PBJ3cuBW+p5fTCxzUYeW4DiYj8kjT4iVzwcpumgtCGGft3Ya
I6kqdl55DI5JhuH076yMWTldb6SzVo5NEeOsJ7Qr47fG658xLljIiJLLZwUkd1bi
CDMcWbswdcyphob4wGXAf0JZH/M/Nm17EBejLs4lrYBBpf0JC9STVU8V6saJtAQ4
094WBAC2ur/tPgR6a2bqE4A2xdidgOH+UOLJ4+E1aQ3nLcH5HzD3vtdYXxDJZaMo
u7XaxqF0tC9Zll+gKJPL8eEivkPh8NFhJI2BGND2yUolzvKH/39BI5ae15XmtKiO
eEbJDnteGX9xgEcwd/uLsD9fhZ2Y2etKATvgB0GhFVWG8cs3HyDzqnRqLTJwbI6e
h9qsrHnjFQQqboiqPjDGXSr2Yn/e+Js+5cw8kisg+HYqPoyxVSdmR4HV9X9MkaqT
YfbBue3V/uLoCo78MfZmh73/jcydcnf1tom6BjGXsTXOLOuhmLv5FDCahkHvP79W
eun05HxofZJrKj3kZhHWN7TgZqUzpNNuyKdLDprg1LYEQf5PnWAepQ52Z4HTZ4vQ
QIp8VBcUw0UMJ5JRq6E9j9kn9Op0Ovpw6EJNRGcyKj6CZiiVjm8pxg4ObfqvZajd
mT8VE1Tts8UgM9i8coeMEDttQkJPkcvrIKP91CD6Ho+FxapKmydIEs6lVOkywOlo
txLhM6tyv88A6ZP+GS0I6Mw/scnAtMl2tg3lNHG35BTtBE+P1378jRnb6vZl659Q
fEu4i4xJfKOaQUXLW+QPOMBT3OyYB/L/LoecYoiTVb8zpAypQgkcJXgRt/Bzc+Rx
HQmLJv4g8pZk038Sf3Ku87jR8DZ1PFmxVyMpY1ox9AJfqEXnZUNyMgAhUEPlQWM5
RqZ8RVLAy2P6T9ZsCg9ChpDiVLBhPYfai2cejSC6/tneUBaUbN3K10QJExB7TX7t
TywHgGC3kykwWgKatoFQEml2YJAf8Brv4DZAPjwwMzRdcGRZgJiv2/gUgXKliQLW
8qu0LDNkvZWr8A+w/S39M3AWvfQ0ejElbKbg/uFPsUGFi69o2eymp+93kCQl4mrb
FKh/FYWAafWZ7wU7qnt6Ry6wDTGEonXwedo++Q5jYuso40PbNngaCeJD2AtuhsdD
QiaNAcC2oHbQVkD/nqVYlgV2kM7UNGY4aqjRXiVafPH9E4zk4c1OpoRlSLyE1lFk
exztix9/eCpXfFI5Gv+1+rrEyXu5MlwlRHxq4/LUS+7wnRh0iwSBGuyR1gXZ8xMR
kUjN3aKzMtIIQey3aZ7CbpzXRNexnMLK/RhksDy/Wom6oE1MqgYeT2phaqP21mP1
a7tg8vI06PDiAKEJWL32/ypKDCEHwoHhUmsqsrm9tWtIn4NGHWQkJGXib4A5rQnr
yNclufMxsXVqBwoSqBpXEY4TFBV9EXNFYaH7lzOTiV1qAlQ6LW7hbiq09d0EYRPs
1X+Bvby4TTJNkH8XTC7KWtQqNlHPY5yVX1yfcJsfy8WFXzTX793QKEUWe+GVgCU+
HWeQivYvI5tdccQpwGHpVPZT+XWeh+qtWLW30Q+9HgErl+ydFFSVA2pSOqso3WtJ
Sz5Gs7P1E3HVBbeVDHqUxxmdhmJK6nxSLLuWo2ffFDDrQBTYs/hdohKsKPQPYB8F
l9S9CYd1dZANybhnVoxojPp+VXjr5t4vXIWCzWOCjLvjRFUT3D9tgrvlTlKh9AM3
2FukKwhlJqSQJz8AIRJ8ceomkb+r6HgwPeEiSgPbgchYj7Yt4UzQoVH2EUmuXuIS
OqQJilszI1ZklO4XbjkK5DE4UlaUYfwiGxF10h0az33YBzm1gh3+gpxG6wctCo+C
twhmPgGSIyAMpGi2W9IZ8+aSYJdPBMFKfyVi9RCmQiSiiWo8oAGqvMnJdNHh3OND
i5Ayn+blH/G5Ha6XDL7yQ0K/gxsBDK4pmN9GR9ixh4cVi8cS75VbIbd9DI0Z5Bdb
4MxVyrlaxFJFkjqQXFghq+nvF7IbmVtmvW2S2k00LpJczv7rVCwHz5rdJn9e//t4
D5ncn2dV0EcLhl5zsraIepUqj8MX+V84nG9OLfPx2MI8dI3bQL/3xFKRT27hiio0
5Y7wuaw9Wzp20QiGPJQvzzV/z7ZGw5IH/sMc4BpdLtZvSrjSiYXAT9LcTMDIVZ4v
r7JVFfK64bm/e//El16Ektxjftl1oVZRIphM9w1MCf/2Ge/kquKXD50au5YydY7G
S1hihY4UZYv0K0QXxgf0f941tt4JBrCuZq++sic20oYt8K5RVVfrgrTYlyO+KmIK
oDvrypUwlyLN9ZewD4W48p7+rNdtoSmnxM4p2A2sf0z1JfA4Otxza/NkR5aRd3cs
a6FSKBSjXa7r6PTJ/CLFGhUFhhANemgQr7BnwjaywxR2tVOGjIaCL2dV370ttKq6
mOeKzhZ8MtOlN6qM4wMhs//GEyuD6Kd2spdbkV5EJLt6j1A3qk/fvlY3v9ddo3UT
o1mADGNEeFnzm/WVGx4pSqmJ4HPqbRbXTkOgYCRC0o+WFRP3UIwTjesvye1UAZhR
nnp03OCeKgVmy5Ush3zdY3/gd0lVNmo2SlBiBoClMFdzyoDeIQGCuGdfz4oYdX4l
ttFsffQWvWpZf3Cay6Frfzrm67akgFNhC0Vf6ISTw+c44tTKSHYgVv4CR3dt40du
j9UuwdQ1uGtuBEW65fS6scC+xBwytnRVZUvxtEhdIWei3O5gq2E1HBkKFUSySUjC
bzbFsy53dvT5MQ2W5rO/+bZaY+BgufRizxDvpgHuWGiylvqKAnMgziiupzrLgpfo
VqVQMx8YdUU92esn+WGlNEraRNh8JM7zig9Zxrlj8f6xzFTytVtwmmC77Q0gAGve
xQ2Nw1cv/Bo4xyMCg+b8DNBA5wkdhRfNp0Hk7cqVhQVfF/P7dxbMb9+T4gN3iDW8
0QEXrexX3rb1Npf3OLbgPsYJx/C+8Csls6IEyfOry+Zk2BDREFRha4XhB+Zqq1pR
E/R796ECInHxz/afcnqw1gZER/JiLGzXKyZd9CgRdGQqcSvH+8zCvC95Bgr0SWke
c/v1yfDh0NZrqLMeEVn9O0gfzWxIZkIH6KthP8psJCVha5obCiHhnopidb4CiIHL
/luSMxzBPjzUu062Di3MhP0y+GfBsJghoKFxu7KCsOJ1deofNOQmIzyJvxVGKLx/
REDQzmoY4CZWorltx6S7XJ8U1tXy8X/sJlB+OMtNyKVrNe4O2jFethOGqLeyAQzM
40XLQ0prntfbwnA/uX/v2FOgw9NBblzPtrwPbhhqiSWAVASsHq6U1qMb8v4w2FQf
UeXM0eQQmqlrWg6AyJ50yn7qtaNMC4d9DYOFjY3XdokLOGEilrwyofJjI3wsdfX5
uSEsUvw2V29afo0VZLcwZEdJcOz6oswJj+tjzAjELifjC4TWjiNFvisPHkPUaMsg
J8ZA2Xmw/FdgQjzxgK65vAO39O3Za+LrzvEv1oWXPZKOeYGl0wBRH/nHyzDoWPrm
HSB4VL9NPPeKdyXVJtWcHgk9UXvagGGbcIuha9Vg1iI5JwjMcDG9R8nK6ROPMsPb
70x0IRMh2Gtqb/t1mV8yJelofiQ5pNcYJ2ueAqVPaSi0hwRATlyrIyWOBK1Jkhry
6tEOy0gcNM6MBqRyYCn1qocf56aaEM4VrytSoShWU6Tw2LFUbilUKrOm2uAGfKPb
9Jf59eEmmGmF8aFAKG9fJIZJl79s402094Svtzd1jKszoASnlY8XJKlojGPy+nhU
Nd7sLvUm6I3gkRmIPsiBAht6++mzsFVa3R7QjmyGHxWwEMdvPBddT1YQmNKotqHL
qaEZhc/GT7fM5WToJnkWdXMJJ9hMO0HhTBV1Xk3B1j1IyYlnyyAAxs1yKrGSJGtO
lIdCmiEGxszn/WWrPUm5PyErG778RGyR85ggvOvLRxxJ8HEo8uLdvANEQ/6B8ozx
Uu6Ogu5ei9kHPfVxwrcLcqFAouAqhpwwj6ZXIKyCNW62DPBPp1wdw9UV5wemZ/WV
QbaObMDjswHVMz+Lz4ftH8yGkff3KaiCyHVHAepFAkVjRwnGV9WB60IJv9zxV+da
eEfhfZpmm3nSC8pd0iDehi/2Z33yrXsAyzUiKI3Qr4hzPkG999r9uGFgHErclodx
vlT05Lfz1JAPTjNRz1qKmDg+l+Wh9+Ys8tw6crEN3PNdbHMokx4sfdeNB1OTy3K0
sdDOSYEk53Wd0ng5509QumUNSo3HrIpWqMt//ctIWTEBmI4Jq/GqvmRkytbaQVSm
1Trm5h04IVMvDinxEaed2LxRp2HZNwdIXd/uflUeiwxkXIyhemH7rLcJ7a5Aify+
DC9kVnP4nkHXFcYKHTPiCbgwsYuS0Ey9ZTeysF4NoWtnFRoj8ZeQhy8nWGpXgKk+
3GBx3G7lUS+UyiWx9QbSCWnIhN4+sR8CeAPQYfYPD+Gj/dCHp4ngZmaZsN19ny/u
06gGBqPZZkf6xRwJf6tZyCKrWp0AFZAzIg/kTt0g55BJzC3EhrixR66hGVCRj+rr
AK//D92LLdllVQ38I+UmkeaOaolbE4NX5cSNXWJM0BaR/W23NmbtVJ+S/sWWJB5r
PMLXdG4q9ZeBz/bR8R7v8lC7ON3IDJcvUA7vbnCdStBnIqcvy4KRG0romq6yQ11u
bZNCKRq4LNAV3EwEqOcjI2fzEuP4uNNf1YUIKMrpL63bPsKIRfsXy4xDafEMfx1n
28HO2fiaaI9ACMuMAJ1omQY6/f3rhRBt66RIfkmaoMuxSagW/HRcMPClNlTpV3vB
Nau7QlxSF8QK+MI9aPreK9qeNiGIA9Y4DBCXXpNnY+lkmU1eD4AhQZNfayfXB/6f
5FCs2NsbSfXwgqD26rO61JXm713VF608rFdR3Ey94c1Mx2TKRmiyUo2e2HKaUFeq
rql7fglLuyJgfP7tF+0yyCEC5hSUWT1QiUcQ2BKAQrE+aykkQBmFSwSLPIYqtqW6
UBfiZCYewydm4p/gKXop7ENx+EoLyhXzt2+7RwaHtorwp4azoT+a2kBcLKKOWzDP
o+kqTbWmTOex8jQYhP1egmujwRViqeieLpfMTEUAzOophplcWc0Us4FZxAEIbE5h
UJAkrdY0cPiAxKsetvDrr0sLmzCcfrFTHg6rVkG79odUTfky+ZqgCnwBoLudlQfb
gz1MVjH199vxI8t37ztgei68drA0D0NLm01nYcFlPz4EIE4zRKMQMpTSdO8FMvaL
7qS2r16Cxp8pH6TAtPQv6I7thv6dioaLeD7lFdLSCORBQ5wBXcGTU1JebTOq68oQ
AmlL2T8gFTAe4CuHuGZcDoGyWovtbCBpD1btRsZW8ytgvcy7LsN+kKRlSv2QN762
3OacB4sy2c/Lti+8yeDoLUZ3vCxOgAVVWKlvx6kAQ8P1cnky+gQ1KgIiy4r1+cfs
TQj6PnpzykabUOabqJWPwThmnS7JoIT8E10mR/boK4MH0j7eaighXu2s7zu7h8nS
Lk09zHN4PAohGFDHmwFjt1JTl8IdFugJr9p8yoGL8mVzwG6ZBOVCltTm9h7oz6aO
8U/Gny9Whb7VoaL6UDEHAs9xLQG+3/xe9Y7Eqvv0QiKqYf3shMrIdhUEOnSxk8eH
Fdy6fgakVv97VN0AHl8coU2exP6TgrSuP3HWYqdAG21RkBXmhJ/ETQipvQF4+hb8
7HZcdyU/NMVBpWX3I+g5DaPFmNTAufMvtRf8B7h2WcvgpbdnHyhksQ2mlMMzBED8
Q2c4JlQ80WW+OtxWWBg7Y3glsP75v2yPlb+yKwsN50MPjA17+l7IXBcrblfvvJX3
jrJi+yazFyrJPRuZVyxBI4C3Y6QWoFyXFRluVCXz6S0BZsyQC4s62HE7NSh76TDM
uLehfIv67deN8S1qAA47rkLwPvSeD7elzm1grxS+/L7N6xqKL22CrO5zEhRAGlA9
ZYICUwbDiVs67jVi5yNp04lgEjK794QdzEa2V1peclQ1yypa42yRPVLoU2IVOSxr
yB9udKlHmNXsEqjCSdi1PcDKDc66/3DKW/kwcMm/jIr7Zy80DlW5fPslTGqrEDCe
A5Vp/JijbR7regU66P9hBoHDBCr+f3u35MrLbBtgWQG22G1CPZhTqkEi+WBiAelZ
v3T+KSF595m64vKa8wGFWFpfHH54yP0RvVbksO8F+kLut+bqEkAS8r6g8ICzsAVC
4llDj3Es6SSQdx/1zO53bvV/Kow55TJE5W70wQ3YutCs/vUqd1B2AMhWFa4V0Z54
38gU9pHmqxV9Ak7MKxxVMc6y0xcIcievFVmt6/A7+0aVSl6Jay3uonGfTXn3cqNB
1y9NpQbFhUfPYkGGHTUWtD3YfklfDzBr2kQWpHsYnl7ivXRZue2Hv5RTiPuZxeAX
IpfsRaGuCTsicbKhWrajx3QJ3xvtg9lFenJ6hycTELcnFi2PpSDEuo8J1vTCWaK5
d5GpXDvPljQO+I+jGsGmVzUIcmyUkWPmmWwE2rok/5BPqZmze+iWEj2+ofGRYkgK
AWRGuODMs0+KWLSSmJCz6zMTnSPTxkPJJUOdaekrefNRojd401m90eFzWZuEfQD1
QV09eY6+yfk6EZIJ96NsFxuskDwqxrFQcvvO/ki9FTOXmkvy5JDlY+fgsHu3ynhW
0sNN6TAYep2hZGdALan7uqliISrkLrRRedTdO19Up2FKlmhfxp0k1RNxb/8bM+4v
QOU3owXJVvIjsC2bCQ4FvUyOp0KLsVaFYGs3Ozzljg6hbku5hNfgS7tf9NoH8Yum
AVunuqbkdEAKDTC2HhrIM+WjP/W/Zl3NYoTh1lYSZKSDecE6FRcuTXzMrOGZaHtL
8NrVJVuz2CLBBB5LXmsHT3OwklIvSH4UXKpG75q/sxqI5kmZE73syWHYtsEe4uCw
w2FdViqgzOjparDGbCtFgP+FAmzUQNXu/ne5i20r0FJyLufKs3/sboNq/BS+P1yB
cLdtH6eNDXbwIrLYzjPjfl0Mpn3H3n9ipnqjlL2kmWSfWJdbWVqkbLJbkhU7APqq
Wo7Oo8JWlfgu3WTdvyJfxtcyrmcxkbNiS2/JQrKhvSVopIOV1weNLAjhcXW6phJA
eDH7e0HHh4bEqeVVOGmm63jyPRTWUVq5qSW4OOokyqro65sZ4cRSXR1TSFfkyGmy
uUpCNUmAqxOxuIwQQV+fm861x2hZwPmrA6zc+jHyDuuOUYQYELfXY0kmsHrs7siw
fPOfi4L7MArwECmO/gQsEaj6FJyTJICsDnrpGIgOqm+yhMAUq1xG/JRl2iPdUMVu
3HnhoNBW9VM1pmwynirDQrEL+9EuSXBjE0SGuGboHeEu/7yhNvREbN9rIXFMSThi
qWSzg/unG+O7fewyrVBUb5NbtqhXvwSlmMYNirwn9Sxxub0OdNVcfSXG3+wTmfwx
U/zUE07SjcPJtXqP6IBAzV4bg5p5dJhqhs6czjdf38+SfjlsuqCZVC116sNogGNW
uR2aI2MKPerlYHWAVODNtkJocu6ymtsxiuLfj2QyJ/GY34m0ib8/Ceooei4qgo9+
C3ksMvccLQqTJy+kNKVI8tldicHKFteXTLPjTTzVdVJ5MA5+nSp3NgN5kEnp3qi6
9iagr0Ya0sx0b4RlN6rTXhYlCAZRMYlZibyjaxOPagad/vMbRxFu2liKdCYeCxnC
rr276tovwWfKui7ojPqyj/d6GCTz5dBhCp9YJCIewosDK+6xbxcdMd+5Bs1k4SLx
/kS6Ba5UCJTVIsMaFis5LJe4YIBz9BSGEXOhmA/5H4+BYQLsGa65xiw7g4LJsAZh
L7hUgrjPqeg5EmkXrjWUiPArap/3Y/O0rjIp5lhS7LSgt5Mb43Jd1b8XIJJJc0LP
mlS2ImmZva21sEtYEAx3CVcgePlBhEQhBrKndXsouAJVcnNIeQiHmAcRNlZHyzkM
ogR1uhY15Zikg0vBXdwsYjz18KOeNUFlbyxZHddrYHSPDUCOdih86/mufjigHD0o
Q9Jj8vYnFFq4fzjdV0cbD3Aj324KuFK3W2UePTdEhE+oio6QWBBHxyTtVfIFjXvU
XJNufBaGimeH9AXBYSvuZwQjsDaPlCF8FUgw4XN2RpHkF+exvmYeJ74Weuw3h2Me
qKbNNGO9KIZ4lRXxh9cI8v9L/tlVuLNdgLHr7fYFn31jQB7rkmXi/XO3wi/gib31
FCyvW2uLbYedQ1bfblNhTLN84iDXNkP6ZeKRm1V0kqfy6t5hwZa6Bx396vbU0MYe
UnOnfsRStSgC0afr8ufFCMg8sRH9iaNLGmOUrqattXeWUKwblxML4oPUQN/M7FTX
tCODJuOvndG/+s61ORfa3qA1VG/VcNX3jEklR0JTOqtfa2IHAFljauwcACyEOKOW
ASi7WhAXQW+MLRpmipXK429pu+2ycVIrIdO9HfVY8kE/sqWFaQ3ugQYlYW92/UQl
nK/ALpS6LtfUtxg/KLorPFxqqyZjMvgY/LSMA+rAicymYU47pkvw/TuQ2SQ6ECfs
BlDknxSX9l+eapu6zWCc/sdqIHzEUrxwvuu/mp899qXGFcTMpAE35c5jx7DrIOJ5
yqwpCqXWRYdwVGb3YHfQQmWHsdchO8W7osJRvI8ivPsGIUWgXh5m1x2P8IOvGYm6
loIRt2l0KB44mE9IrldEHvzg1+PHX+CVpPKN0OnaezCcf9Udjn/vC/2NxwCMcif+
8WcNpO9NstSVdRF1N+kyJbv1SbxOcurVVgVz7ALFNmYfl6ycDpATwCO/rePUjtEO
QXoEM85I/Orc/nwIGWx9AUnE8UATH9a+gwtGSf1PwMw3+5EnRNo+gz5ghsUp8Btv
F7BOdbk+lNYx4IrBD7O1K2PokxAIXc/MUwVVcddsNPu9+ZeJmBtyZ4RqVJkpW+qz
3fvKLJ09uxAWFQZymZ0T7v1efxTg89uCkKuqB3xrXaOV/uHW7xgAm/B8Q01XhrhP
4tWOgkMg06x6rhN8/Uv9fM+DFMpgtmnWdw9/m+Yyl6EtzXwXuIwPxaDO7Q6r9MLh
cp463tIb9vuZgsnH+U5e5ouw7hefviFM2Ore2rvXCPECMJPpAC78vHQVZMQOsIwT
10ZqHb4gAKDTZfjAhxqc20HeAXSCc7uJrmV1GLCAo4dvzk3KUw2ib67j1QPo45RH
GlSJDgelmaHg+OMthMtGA9jht8vwIc22MQvhDxnJ4oTPZ5bZynB8AvfNvXIoyN1J
OU7oeRE68NzVqzwAj67CtwfPOcnF98nxDVPKrLexGRcYtzl9GhNiKwcBileht3/V
0XTI6Mkks5TyWqEPOZ6GNg3MsPUSPbeJ8NxFH+LkONARgEOr3CkoouwMZPo0F+8A
aYuFjAsYdo3hIO3QLMySVeD/adHkskfv1vkD/nyIyYlFtQXKmNMi2bRj20GZ7vUe
pdV5L9nwI0oi413Fd1AlAfzsbolGozaRR6/Wg8P6wzaJdbVN4DX7Hnigw2Sw+6Ab
x/8O7Mtrzx6MjI2nd2x0kqYWtOCVOOBnL0Fvwe9+6Hbzlk68g5nktQrqBwEFWCoB
AqunPU5zmjswnmGW7GtnKFdCgkcP7sI+bL1xctj1wy7tbXJEyRx71JlkI+lr2WHX
Y16cXe4AiTROj1wpAZuvKkoF9wggSCt5h81x5CW0B5NJK32ePnzcjB4IjAk36fYH
cKvU0XmuGJ6R+/kHOB9p4BQqrOFTXlsfy8gQcFq44PsqTtjaf2wdxynvQV4V7YMH
EMUOezdz+1Tk5Nt4W+bRh+L2ecB2mLI6t+x6bqddkEC0F3kmMpCxzwajh30WReIq
OLMAqF+t7srKkyfC3MhNW0150+EneGBCS4pcBQQgdwBLFRPl/zDIQwXcgOpOV3GB
HiHLeNDkDvxV1j2AZcdnj+4QgaaFbJQsKfhYrOGqMFYxHuHyD8KR7YyOS/VdvSnG
jcshgKHL3OkR4sP1krOWPNve5LhsYiXBwomS+SAFkV1vPC/icBdnZIDBTQ6bxrqL
HCxk+sPGOodNZvhc7oHSFdw5R3pTtmaTxPXyMcJDeZjJtHbgZX4x7Eseqj7uKlTn
ZEmIQ+Wtkly8c6eixf1co2zYBqCKZRiFXP9yHR9hwEwLNxxmQak5bnGiFVw7u9Wx
FBNUxWyFxRo3iYkzs2h8uPPRRbti8ReNqZFhifV8NjJsS3+u118U8WEg/0FJCnDt
EKDTL0cilEJOTodXYeHM7Bumy4g+x0p3kF5AnKxgpdVuDgu0jSgT7lCgilEsOZSh
BXdzfF4pHuMGATCqGJkB7LVX7W9RJS9HnHWPICsb0mUJOwEJJk8Rl99y8Hj2ZtZH
pnMWoQDFjNI0ZxRceqUvHdTpZabMDVs8XAlxKCad+F/clf1ySNAiwsi3Klt/pELc
AS9EVVpz30nkwNx1aHPQT1egS4RPUtm0tqGtB2KzcxMRs9ygYdkTfsz+bDT8ja/r
szduf9dfrk5jSBsfbI28seh6tcAAnDCpRBuBriTAKga5W7FzaIm0c8V6Z8IUkgIB
S7jF8rfclcP9VumzHLQrkOmRTqaKHniwFfdEPrLwm7/XEyGBG9BH6RK4k4F1sQHA
nuXe2MzPnMXYhfX6qA50T2mFP+BalpcfSa9cKR6Od1iBmGeA7b1Z0t7Cu0WiPwxJ
k39ynm60JXQlGEBW/3oEg7D4qIvpbqIe/bth7Rz7O9AkKyZpZR+kGoAaqtGiV9TO
i4JqjgzPo+7DRitBZPV0J344C5C8HSmw85ZSPRZMJx1k+TPrqw/dg6wbpwXmPhyp
i9PajiIGsUIrMaX096lePLeNYHUk5fpbFtgrZNhpKbZeyFEh6ygy5KZo/xyiO8jB
O+tSsCD04r0qcBH7McOtwZ8XkReV4cgFFJtRoKZQPiUn161VgvOO1snSficYcBgX
TZrZw9HsVtp2gTe+/wAgKmI51uYkiuOnFgoXm9UWAwEa5jGhJJzhv/mEGcEgmHKH
UhZutYmeENo4OJPzuVUqzggzmYGxooeb58g14BIK53bjFaVQBstLTgPAmtYf7n7I
WvPn2KOcMd9yPOuJ9JIXQmSjFDv+iWy2xSKv7SV/tqocaldoRaOGDfM8viGjvedU
iOObOS9bBxwIXjRp+07JcECtKrWfehwl1qPS+JxPaMzEcoHrEiXS+ped6h1m9+jH
eC1G2WYjnEoy4Dg4q15T+stSqDx5+vBD5GXTOdFlvbcEVjbi65sedqiGNz//0K2I
XCkow5OFSNCUHc1pTT9y3UYPnB56S+g8Ba2mQHve+c1tkRwHOVW1V3yFVhOE5+G9
ZpBDNeQgj9mzwKdfJ4up9yrpPGd0CfQcWS6/WUcqXX10ibafsthY6fpzC2y3Nh2Y
umkk2yotfkUHtG0xQ8dspTTNV2GztyHpmxrDxtaYBlnOLZwDoBxvC+RfGUGPjUYv
oEBdEbguLWYul2hMaxk9+IbWoRHT3HjM/6WRciTGtI1y6qE2L/5MlLMRm05YywGv
z//KpBRPDYnfro1hU5ZugGMFLtqVQv3DS3l5GGFVBhQozNqgFYuqofmj0tcCs+Hu
PVAZ/mYCNWR9ohIIsTfaE8JEZ9lsD7PaivD9VYMrnzjIqdQqWIzt6hDpof4RP+5S
TVlwtSOViHcnYBsqbggL21dvn80PfIegMLNkuLwRGEdHOk4P9fdJ/xbh6+gBkRjQ
6HYGL1SwHLzGVVqcJH7G5Lmc/7AQ8t5/Jxr+iVkT5OzQ4yzzqYosI1jAW1ZgKx16
lgxGo1KQciSJVlKEEzaHoDf3fVq5KPKELkwVZ19uQTWmY+OzbwSI1t+cKAPOADiy
LWxgQCyMiAkIDrLKOqHcFCSJpumLcq6K4juZttrtghcLt4ZpsOG6eK7HtXi7DYU5
dVQEkY/Y8h1ZB7DLFVY1L6CGZzaAPk6IN5CACJXPO2rr9POu+KPFTscKUtFYMfKM
i5MgZaf0VeJn6IoBlLyFiDCi0Mz3pEnmpa0LLqEfR9Oe/SFdkpAGLYxyqC46nuPO
w7tnokkUHhOoC9XqnZc8svXf0ecTT1RhFUJ6Qsq0pl6jt3nCpm97f9nN+zseZvS3
pkg5nzDKaKg8FlQ5UDZFwNME5WXJnA2wMX4SoodZBSs4ViEy538U8Jk0oFmO4GJy
PKc1VD+l8jFv5KqzGzH5g6CWB3Ja57d0Z7lKmStDo3F5smzlcxvgAesPkzWCtP58
vtsrVQAdxEniqGEvw0vyx5eivH1ck4f4dZNFfOVWy84Le5V1EYSgDC3PG3npqWzP
ipXDwOn+aI2v678sTJ64s6H+LAz/qXgX2ulLj8nXtIpv0WFt+6DLGPXVVPus1IQ1
8bG7wulhGz/bA1nT1QTWRP74TyugGn0m7+ppkoiBsqQ/+P6HlMlx+qixWxyuU4S6
ahDMRMWIiDzAl2iEgm/F8iostNY0FCdKbwkxEGM/vTWSEa84PlvGkqkx/Gk3HQgD
PVLJovwtt04RcO4r1orY1ehfsOsx8HH1bkrtR4t+SAS6yDs9nxdIoomVUfcId7e7
sTxKGRhZydqoLbJmThA2mPMabJ46NHCl80YqyL8J+xeVG3oMNW3qfjjzWC++dJxG
hiYm/2r3Rk3V6h4vMjUGm6i6hstkzWHSIOO5x6QBIs554AKVSa2RsWg31jJzfzWR
yynsRpWe10arB19q1K/99URQqOqyfxfukzItiWRHLRtzk+FZ466qDgZhKqb78KsB
vZJHh0FgNmgKJ8I075hsT5v0K87+yNKBSPII776G9ej+uyKWyAXz6Sby3GuUEdny
rwaZHMogOyHP3t1P6bI5Ippwq5BEdkhCDvbzdePTmQ0S+QV2ELj9Y9eTQLCeiozM
0Q68JYkC1Dc1lcEY/4HzGFO6vGX3lksxIpJDDsNzJamhPWwx8pO+gjUNyfEdiVm/
RjBoDX/q3xsgGllDEqKgVbzaf0mSMZThrpgMA9WaxQk7CDDUvhQ2Z40rCmw5blgu
Nz0Rs/UQP/dL8wUsfyWYmRqWU3gMp4woMKUKAMexp8B5Pdm7I0oGLhyu4oFlk47A
vBK4K/2JCiw5yAsZfNiGWs8s449bK3chBupcBozGhWu5WnXplz+7FBolT/1klyBU
GT7sGS7KrMS8x4vjH2y102zCNUHBcRKwSk8pBKanEm6RMrvSOK3ncfWEd0Yw6hP3
bw9DDJwXA5+gZ0GI2KUXogoVOy0Hnq3jib6HqgUEcDZSyMrJKxBLK9wXtDLorfzH
ZX3+WYuByGfD/LRkmpy3L+R13yXe/L9GA6mDdkOlVfEbKvrz8vKffhzeiMR1t0LU
a6P0AqA++JMgAGMhTfBp77gy8RH3HpK7EiXmfJ5SqBwfAF+3F3Fm5k2TvS5A40O1
ZdSaxmd5VzujvtyCHvt99g8xE0W01EaHnQgn3cEeNd/pPp+9HyjZ2iPn3rYQzlz7
fVPvfIh4BgZLR7q8a0ro4y0TRe2n9VdYZq+AUlf3dR7Ynm648Op6G/qqB+HdUSoa
ul5LH4A0O6TBFfcN5lT4CX2CMMrD7VnkWwk0glT21UIFSJVYgn1bDbBbyFWJjMri
O6TCV4FuztDZTnBO6Nnxa09sGkLNJ7R1SM/aKN7ij9hZemDh/PzLThelQdMpHkB7
8ssDJl2X/tf6CFEw/1sgGJafax3tuOUDWJbXGSHbtPNJp5gogI7tq5BKuHuPqpn8
aUOAjLTTQTDuP0rYK4wrf6A6fZ8JU7gGkZQmA6XU7fitAkNu0N+2mFF3diWrhODj
ZzrXsn72+VOK1qpFkXpf+UnMFDGUF4ZKl+Hcjv06593l8RJSpNRWIYr6s3ffn3KR
v6Q0HZ1rdddhZzV3MtGUz0KOWD1bxzos6EhZpmjUPEDLVY7DyLCW3HNhm/5OHSPd
uFcswTnkg4oSu87dK3Lr2PFL3/pCg/LfsD9SlMhi6sJVCUJSU8VBndH2h8H30UUt
GmdjuleRFmr6Sb9vvJ/2JzV7Y3+ApznemWuJLDfW51aOBZOI3oPdK8QgnPqMJt4L
t6qs/H8VX4KkEONn1LC+2x7Rr/MEMPOQ2CxdTD4R8F0CupPeJjNoALXR4z22WMXg
YBCR+ze2n8z6B9O7nwhXKzKh6IJqoS8ZXGbB7r6OaINGtqfPWl/ITTe6POFa0Lt3
y0cBZDvXDnm5GYy2jG75512Xg8f3AL4ktK7zd7vHRON3LihiQbK3oHzyu/0rPEeV
MpCCRYmmQy7dQ2rR8H47X0xZm+4/1ZJYqfvKbsTNuM9J1lrB7gY8ZwWcKPuyf9qm
kLdmhYSS0ebYJeyANfCkXSkzLQwiyTw9QDVnbNqVsEISADCYMxQ68SKMezk4fIRS
pVq1ocX2XqUdi4vV2rVEnzAoi4EPQvSnHqy3fKJylIyktdKrXcEfoQoG1eMbE+yj
6c33s3Nxk02ZvONvt+OGNLaSNMtDw/1yAH9IbbnWSGba28QtrkKT7bYTKWKMZ3Y4
5Pszj9wvlr/eXgpaX1dMNw8u4WDXfLwX3jAu+S3sLmIS4B3ZpjznBIAp3xExGBiq
NvbVGCWrlLAfdFCTCqprghvODKHEVHabeSFsBtpFuh7ouZoIT//hqwmGYlBOQwwn
5/YNyo14L0K3BZzfjK4sMfjr9vWwgJ8uTBXugOWlTzcGYgfSx+iHTMPHnTsGX8mq
FygQIln/jhj2l1QTEoIfHlq2GDJU/AxNjigT4c7cNCy5g80oYPUOWBWfU0fUqfcV
jeGFU4C7lnmwWjq5mOnO0UINoCFzXSPCBTnihK4H8Vr8QYoS+SAtFrKz456JluXl
WSTKPXzF+HG6fu8dDPImAGDkdKaXqVBgzi1bqb4OE6L2tk+O0JZl9tHsdjMT8hNi
zmGMFStDS6QFiAA4v/80bzlAm3BVEuioonk3Mh2ihqe+mYo/nF7enrIHBpLTQ8eJ
Tm2YQFbtxZjmKgtyti5++x8bqGO2UJU3Hq2WkfS2Mg+zcgq/dnHRT3zobbQgXVgj
lqMjqyR6YwV0XrJ/AlJCQVqk3bNsmOyD28sJv7ihWMh01NlTW8CRW+e34eYrZV/Y
+3jeExgI0WgNV8oWKO8UEuFOZfdkagQlJGLFlsIYF/pbdVX/6Ie5Ri3Z4YhcchfJ
ne9NhPFTCTofdY1qjtOTPJ5MPbS11PvzPGilHE39lF50ci8SXP/smbpcUrjMgdef
gCX77JTh0HDyPsEfT0F3sUmH4RQHAhOkik0mq8wo2HCjyelbx4dbF2mV9LrSsrtX
lNpa9B1tRhhyrHuw0ah+Jn8inG8uLEGacu1M4bo4U0oT0eHDUy/Z5UK3eEDzjd3M
SMoPNMdf0HOX1lz3BJlPxFUNyeI6SGAfJw7mGg/zjMUV+Oudc/3uLw85cd1eOqu4
47yrD1DSxBcwkgWbp7AuoVlGL7SLiOWOnVHlnae8tgU68xxACCzvTL1+vLeJUj4E
+WnjvWu7p8GoDAqvKk3C2uoz7l+5MVvqWpmWhPLDGhXtW2fA5Yme11mgzZZ45Fob
yIwhNNyfqUYrijT6aWxVvu9y3WfBe2EiHQmlXZtXNMx/+JYnLfreOML6Z5uXjR+Q
8lB7aZ1QmpnyMCkS9SJ5ZdoxJFj+DcoHITdncsAjztI+aiwA24p+cqmPNHO3fbpj
ofM5MreqS2Xx6ilbzNm790aNqOjUGcyddaof7K+D0iFL8ajIxUnPtwEl+P+vNGZQ
7sTY1J8sL2NpC++yD8ekKT0wPyxOUyuRPaMTbHvDIUjhuX36iq3hms4XNOIO/2IV
0OcptaHe5hRocJLQ1J2wMEekUcnH/gsV7Jo70jWwxthUN3veeYpePLoo2PC//Ibu
ON1/uNJ1+5PzDMquW4nizZr+Gl83KsbC8etv89oCuFzfhS20p8iUcpzI/djJjBg/
pBJIh0df7vzeLdXVZm6dvI1xFdVvoEzOp9j46tBz8wbKVRtB3kMCf5YbZfPfZXiI
LcL70MImmPOcQ6klWq33OcfgMX89U9527OesxoBHwU0MZ6oW+BhSjQ719ehiBUIw
Zkk+1IqsPOSdVBA35x+LOsxNVGx5jsT/nJsJHP0b+QXhv6ttOZ4FEycXFiO9p4Mr
Lrf93Q6hTt9BgOSoGZmcIWvtwAoccOubrFO+nTNUKCnWwhWVsS4dgES+31snF3sB
RXOAZw35qiNQsqFtbRdS/qQPcnjWnbmw67Si6RR2j0ibps75PujOVm06089M2tJt
smtpJpHK4G8nIIF83EgB8UH0EbUxHjXsLbXGpflW+I1uR4J11SxryypN3O2r5bNs
ngk7DwRXUIFug+4F4VVFlPq4bKExmAcbcpctYVNzKNHzMXwoJzr4YIzi1wYg4ylg
QiNEDlM6YGq/VmfVP4xETIeCb2FWklMRR0pY/Hn/dCZAKzVL0v6sp4SKz0rUH6RO
tIPGXnsgEXIobUO0PSBGhZyI+yGwwAjnyA4ZeFa+EyXmFdu59qKAbNXzvFM3fzYJ
NU6paV/N0k1uUf/JdjwKVTc5GMP/HDzPtOdGrz4tLzc7vxfcQOffKmGAiUIQwDIn
83x2pwupAz42CBl7gw1C6mSxM78HIai5l4jpL/cdxU1R4cmPBz4Djz0qoJkWW0Pu
ebvrD3YljaqWuxZcnEsMpvi+EIcfAMtf/tAZzfSiibnxxogMAly6l1LLE82KIqg5
1/+lJ1G7yWYv/yE7z9sJFzJQTD42h2TFQg9DM96qSKPqKyiN3BMRwIhoWu59tqTt
xg+x+JQxG++3/2XNT0ePBbzjBEHs26b0NSl9+KOef7sBJKj+b3IASj6AI5m9E8hV
H79WSW23iK9bkII2Ius35KoFQf+xoPw1RqT2WyiNQ0jftnASIi8Qux8vCBSSFPcA
kQoSbmoeQ+qVyymf2eNTAdu3pxEJi75bW+fk1JrG17EkAQVOlk4q8yiMx3C8+H56
qLdcvDwn0OGM0JlutumzEVD/CBkPr1u9f6XsJmftFaZ4Ac/M9Y584t5CNR+YtoTW
yfN6CEz9BYHkzWeGkU/6iKlCjaeJZoYfobG2raV1HdQMIAXxEOIAP+VILit4wC9A
rj57DlPDi8IR56BAhhDYJbbECQgV74oYiO4lrOqB8glcHP1EBOAZGC+Q4lhponey
bEo1LLouA1+7tkzuL2fE10r5sTiVkkgXK7sVSaDsGxOlgL1k/QzHwfepYTdDnCL2
Pn76ntcno6eSZCdz1Jt3EE4TIu+IuGcR5uNgOYKV4qzMSpDcjBJwc8Gd3FHzmfx9
pzq9WRY9E0SW83YA8X29Y7+QH6jH+OqAPOikNXsR0neDZ+XEZRxSbU0ym/NARmBR
swuCjTk1Nf8XQvYqBjxiCyR6zZ19iSlLG/i1wfUgjLV6CZz4h3Nsj37Sqmeg+x9O
iPGeYhtCjD31EiAUKJDuC8c5WoXH7vwAaRy28/bLRll6kjJ2Jq/Znrp/TV9lXi/a
WN72gO+rT+9odhx6Imrr1+Ui9HDu8DkFHtuutOP6Ea1xV9Ty8K7iDENe2nPe02tp
62uobjlom2vEbSb/r4uu8e8wDYEU+0sgojSlu7HdORei9MTxost8zws5jruKiVx3
TwsI/s9RAk7A/K0BjswHByvND0GoNMINnf4om2SWLIsFjEyDQw46XJe8Rj5jjZrr
tQNu7uxhOkik64qtpvseA1rnkKkgQ33qb3ZxuHXcxvUa7WlYwNOqBNBZPWDgI3ut
WRDUEYgYZy4VZ2VA/dzRvgqNjAeADA6ewunI8azb5uHBQ64guWRe+cfh4mtwGIma
pmWtcuzV6708tgN0Q7w72DalbJL2b7SvAlI5bpj6/ha9cnHd6Gytp/w6QNjNrDsu
2s05lLzbRrmfgsG7OjwdVsFaAF/9p5HNme5vrRVvJkrqzOuxJijlroKBfBNoawdf
mOPGarebGkVrKrlPEB+3QUrV6UH12e0ORa6gEFGDh8l/MM8s1liRB0VUIJXYdhZj
WzalInranRl77bhWXPcKSg/jsSIT8Ny0bVbIcpRG8XPxarzO8FM66GynlEJm8lEp
ZDB50GKiI6OO4FxpWjKzDjYqLJCOdluNEyPJUlKZzuVbrxF2mceHmll1TiG/EQP1
4HxNCg58qDILcaP9S7X1UKgFjV6O1MpX0RIHUbAXlKk49GYtMHVb3vYY9SjgrxqS
kbPQc/8VjxwQtpzT6pBfrSR0NKt5b7wZp2mVwBUdik+qEo3deoFcKmEHQB7vQNEx
cf01amaIuUUau02riu4OTh6tfYfSxgRmeLyX6rgAVEd1AKk+2kXC18119iZPnx+U
RItvswToUyEq4Oamw6I96FuKtyVWnOCsIYDLEpINO0p55ugTKRqMKBjBEnlSYjOc
EgA1De7rc/VOYiZfqfPofgG15xVZOHDIhScNxQllokpQxfYdMk/evdu0pDF2GCvw
t8LqXWi6bDQJcVG7Gg4sD2ay85JG+PMpMi3haclCFaGe5rrJprV04cwHTjV9Q2ZK
7zE7E2xvh9MnY4Kpe3hLIqNe7hjKFee84/plH2JNx99Y2sI983mcWuDsXoo/quMY
fttuLUAQZfefOLn2ITaL5vcqI2Fo9b5pJfW1jGTixHN2o6/0pYD28UqlfcPFrZLQ
YtjKYEOGgicMGoZyqijwCiK9Vk81lCzIISnGtZztnQJP8ZyWI/QZiv3aDV0xUliR
BgwPDsQ+UxV4JOfkE/QEBGa33wY3T8H8rwZV57ltKJSvDWQyKEkBin07WrMQnvsv
VO+P69A1hvSjP5jY1oKNyO3XaKhXFx//0Zi9w/eW9o9qBCxbFN6euJ2mylLWDYCW
7tbHEsFEF6fqmLKhDh43pKUzDTKoqrMDcWHPfazAEP5YUVi4CGvPRycN0Y371ixA
pTzt0Rt97aWdsJYmnIA+SP3CG3VcDBD4seTTAEvFe8TnDkWmxYEXwEaVoTdqYItE
PQSwLK2ElTopInUKMvobof5ji5yokP5sUsITK/Sjp8NcPLCAMU3+sPlSx0D2f/S3
cbYNy3NdqO0fy4T2ZBMP0fS6CLp3ZlGJI95IOBqFYCTwm7xbh3nHaVQRc5lc6gEJ
AOhthW7Lyu1BJhYPPMJn+k/+pSGkEDx1ULK2NQAdIVzoS4KhavBsbxlLMzrnSCOf
IYPyX7C/ZwKzTPecUA1meW246gkYupxcNyFcwqIBXM7xnMcvXUJjt3oTIMIG8Gdt
i9dBgwT0StExTiQ8pG5JnUh6utX6+ze3tCJLYril+g6431GRiKfV5gunw0BWVUgd
z8p4YqxTnhZ/F2mIHA5opZw9jnXeQKHZlnEZmx1+0/kFV8Fwq7cn8lKS2dfOReHD
DcMuqjOEYqM7iFfJpFx7V71zkJmF1a6L8FTdXjIKMF0x/I6dpMaKrZPZ+dNthE41
SicEHQRvSjuAW4iGzJ9G24ToNxyiVGkBqGyTJlyHyiloMiN9Rw067+ccowNhj1Ms
2yDTCsKwY9dkm2o4DPUdB6HETXnj3sdKYNPe2LlwSg4bRgwbyfqs6slZpK1Rs715
N7Ud0jIYuQkXOg4IR9F6m76FHZ653Ur+nOwmpq2zjT0DyUfCd47XE8w/++f25UYB
PYVn20781IrWTmbiKX48+GRfbusJkxYvtZ5pAy2OP99/UjKzFyxpyWdOH5fgyUhQ
rGW/FPx9Gl26XtWa7USj9BFSEuQqOgcokfx428VBjlOlhIoYMJagQbce6IPnlmER
Q4K7cxueVxNtHPBjjcPDq47QxWrXPHQ7O4Drx7fmwk5vBXRTUwg1zwCoP23HvSjA
DWtiLGBzPyAOHulC3Y2IbBeIoy4SoDiq6sHAeO6gFiDh+co7AwNrHC75x9cCZUtM
7oTdgBtA2yNAPpd6HubeW0EA9Zd46cNA43Epm+bRXtM5IBXOS8VlmwnvSh3cKgjL
BF+VKcZb69N8+bJkhYxTSJvFeW1IzdHaN/PmzPNKVZPRvI8N6Xyl4EeCaaRFpy1E
aRgyz3ZzPd1FWzD0a8rnCoQ05oWakUEVMBcwkKHi0zq86+j2WE73DOC8SvC06X26
CJkFzTgCnFzRY0q6xdvtozGVwJLivZit8bKfr2vvu+zmpHt5F7agYmq4E7slhBGh
U+eBZKQjM1Y4DiB6QhasQhnJsOstiNab6gLfKneXA112qy4ywKt5gMq42r83Vekb
JltOeevgYzIQZpLetejBAArA2ZDOkH2MAocCg9OZKBbhzsgHvxnAnDNZiQ8pUvJK
1E5F95h426LNIfd5tPQBLwtdJP4H/3sXPezdFkduo1/a0+pQLCFYzw/bZC0sr68m
+mzb25OQd3mm9EzU1g6v92Zs1a/tUNunLZ20WY8SgrmMNcDbA/cJXyx3LKnjSGdb
hGm8DaLcLypQDeW0uIli2exG+IUhDpB/7IwD36cAeagv3Qv1WYglUsHya6xDtlns
p8dr6yOi3vViSd6uC0bvVS8C4pD+boRZNbU2fwyvW0E0Ia0ceO4WrWHaWtJi9e+l
iNJVI2q6y8x4RK3lesHA8lHW4jcXU0BlBh6Vh3NwmCZagOH1BZwRDhdCTacHD9RA
xUPXR7oyfw9tNJjKVrOUbqEesg7jwqpHISGsDE7cv0/BTVffEyox+orjkSFe56ys
RyUJO5QXYwmmbLUO1sOePo4VtS0Pyu+4j6dai7dF5xIjZ7TByW6z3Sgy1O5wSRd1
FQKe+fOPYNIJMLp0FOxJLO86Bu6Fi7e/67+uot9rW7m1ymMUXzS7fbkx+FAItDh4
g2UqknpKKVHBTx3CXyPeP1lp8npEWONdpOhFzdcUxCGsW8bfQJEzDkbLhbG+CfNP
nNTtfFakPlAqL6g1QCDceUuVjIGLF7jAc+G+Ki9i0rQAy9OA1mE/fKPnltAvaueH
t114+SpOA2YkZemFqtcDXshQ/0Km9ZdLlVzRnP8wqSxaz4MuiOLpsrHsA419SCRT
BUTYLDyuYXDK79+s44Ba/NWX5eD0PAoQ4v+Si55FoRz7dRwZMdoZcENP0Zh9BQta
nHEZO+NUwG36+cIbsOjhMWWloYfajsYFN+Hb2K6S+pwsOzC5XQjCx/vTrN3FfU9C
M9VJSyqDXpqyA/CUCMTi21Dgc2pkP7nvMdGcurfyCrHhCF1KzqXNerArfjV4pXej
w2jt6tQ2ljJ4mVjDBRZzwheCMlEgFB2xsw4Vk27cXFtTHuZCtdD7z9z/pMKVkt9x
Ux0qVnsUEXawKRIKzhq70GUU7RneLFc37/odDCjbU+2nO6182TLiU4MBn2CeJ3DN
bcGQ63I4xspErKORisSIXNIR2H6PAnm4mxD8dFdgZ0gxTZtJoJdaOH9SenNJ9HDx
9k4+Sco/yPqPS7wIY4FQndq2ip+3HSYU3Q6A05aXg7/rqfvXa5BKq9CwbqEvNnqT
bNS9TfaaAa0bYCCSY2vqWyyXd8X0unBrUFQn4Ilg/jIaNgLca51STb27xrztWQfS
h0gK+SEs0Cdf9Q5hThzkRkP6URPyxMYo9sNV5oiGODvYcXH5/Dbengu9bZQTxjaG
e+gfvBUhEOBzwhfl1MSkIcnAuvi+l7iyqZWCcFeU2/+bLzpXf/AedFYxu8eHabMO
yuoGP86itCeCkeXj1GLDNoMFqmR9deQNdCtB9vx+3zFqnetCNIesEEqUMmNW4IIZ
v6pPg30MoUSdboKmy92gg2n/H682R+xLhzwuobE6eKS9aYiYd/EEJQwqL66ZKuXj
2wCff/h9LPsqqkqINgSRNjiKmY44xfJbLN0vDWtdWvkXPSOVHVn8ca2GffmArKsp
gXs+gFOAy9/bhQwLCmVeGqa6JRfIwH5/8XMw+kujbeOZbQOAntIUQ8kvjzIjyEuF
6e3T+HpZSjeapt1oxBwtYxsjJE7okkwG/T6yKPJMVdOWKEI5cpHkE7tKk97T8Fiv
XjpmEz5bvtKBzzWhMgB46JmWOMt5k61PIU07+B6jCQmbIoecrxAPe8DTLg3LxWUz
JAd9TGckX2vQkMGDmCRfJQ850+D0ydzg6yWx0AFAAO/cg89AcpbcrKxLFnTfmBY4
kAN29+xG2SE13Cc0Gu/1UGgStf4NBAT6VIddefJ8VpNyINKHsw9QkCAgCMgZbNQY
ZdHArLGrofT0Egl5sflPva4J/IOCoSIejx97K+G4jVtRoA/xAA50Capv9ce+SJTv
oc4tJzNliU9q6x2zh9247eSGeJ/it/HBdkPV2KdOPkMn01kr/KgWcl8PI+O1udZu
i8r8eN0RVr2Mwu2C9XDQN3hqr7r1lxO5i7y1CSlJ3ii+vfZ8HIRNsmCvWWnuTgOa
OuCoiGq6dM4OuU7mivXgqLX9uBOUAQWbeo7kPWgvHXVk2gjlhbF6TNoBstGsJClV
BUQYV0xSMsI+uKAd3vQ5t4Jav4DHap82zQj8+/etgzxQFqUKLSlwBSBYLzpAFMuA
G4HTO99HulMhIi5h1eIVhLIEsiLxdxJHiWf9CvysykL+NCgFu4j2Z8I+fp4dhVQg
C7zHPGrXcs7zhxKkZsEcj8C0m0oQiGji50a+o4X7Dkii6mBFT9U9vVozivG4Ctdb
qSutLIGmsXNvavJdDhkHmnSdB1MtNMdVfiG0PuALQUL/EZ6hI8rD4qZ4bQ3xtqCb
n/IEoOalq8L4ZTbQothaMFF0fpEQaUC5KI8h8goZVw1X523f+Ac6LKUaDBBz5hrY
UJ7rvxudNdR2C+61mkXo91/V6U2xZsRnnQLU4caDSdhFjp1Wchdq1L5Wx1IeQrtJ
q8QBY6gVFzwt7wjNvlU39pqi0LL39gAgA8WdyyzEWNPkSD5hS8Bt2w31l/1OtSa8
UxGq1IhHGKihVlxz+3KxeWI7JzKhrPD6eRQHcRW4NZVgBIxTA6jNAdCXhtVn9E8u
VTf2Qv6SSSLeaPDAJ5b42+rIXcMFv9tzepiROq7emNOGFdkDg6MM28j96enzXVzJ
YIblyVIK2daHtGugXqGEIdQaqzB8vv1irfUcWtZtVi7/S7JfYZuGmSSeVDb4D8Su
EPPGwFREfXrkTX4OqVOiLlhmUOgEZ7QMz1KHGUGwPgDYBC44BphuoA2O+zvsrORs
9V5bA/Oz83W6ziGIq0NNsP6sRQr3aPNaTApsg4kKct6tD2hqjd7UtT4xV8kjWiVi
tB3wcx1FnXz6IK/D94Ro4IjhGZLgTrmQZkswPi/wtrp9sWBlHRY48gvP7sOAq9d1
uLhI+TEAaK2XtI647G2vP/EjgLHQRPAhgp0RfkEcjurcMgbL3sqQShvFDc0iyUTQ
M3RWZaq6utnywd/wKbgQFvy+2M7+eYoqdDAJaEXaaFc2L76Byo5frxhU2pQdrOK/
mBGsF89gHyEJ2+Af0+Yq1ax72vmyJ3tBcefzVnJlCwXTMEMO+gx7LEn+L36QY8Pd
Pj/WuW5HdzFqXNeUgVXdeg920PTbhhEc3cXmG4WYwJnJvvw9YJjwcgFq2d7gC7OA
HHaCk8EwTds04PJI45vSvjSuGYf4tammp/k44ShkTHh8/uS279nEp2uQXDX26j25
ciVl5KA45Y7bOTcQos+r+wvwxfjMOLztBr60hxMv8/oh9nvXXt/clyxA9H5+KQhD
g3LVXZw/wzzyVyGacDkf4DajpKP0b4IElVrs5sUbkvWCtTPUPZiKRT/5MaFkJP3Z
5Adi28iRwe6dT/HhjpHPM5xF9kh9pSrRF2tAy+7/6Y2GEwJKnqfVqqwvbavCAb3m
JMKZdb+MibJj+rjfD/l1t9t0H2zTrNP8qDAUT0iTPAuzyVDbULm/zs05BBd1z1x1
9Qpe19wm4sscFSuY1dmRGUVwzBFSgUWs388JRSipYlMwrxXusPsHvMjqLCFmxH0f
M/kzf0GN5YCDu6xFOiadqcWqwnfj3DHMV3znL4d93GD0r5NAUsi8KzM1Zc/cWGmy
uelb2TwPj7Fp573LlCh++u9vYE9e911HB3q2KB4M3aN6OTh3ay3Iyun74a3PU7Y4
ReqPtLg3Jd+L0CU2lx6tucyo3Ux2Sb2/2ipM/QCAauxUAn5jywPqyG9mM9xArPJ1
S2kr1hBeeOIFN9TshdUQBiILkXlI6qTZycR8g4ca9r+SZxUpxOdSS4umjwt2CNEt
w0dYDTF+Ha4A0rTqoMf3/BBHbYTugEYiHxjr5r/ya4peMv2esZSW6zXzMZi+dFWN
8QRntZjFibMNhfxTnzoZsvpkrVDrGd8FX4A/7XCxCirgl73Vu2ns2R3YZiQs3Tis
RtpmsXDboBkiJ/ktWh6CJH8ghLwu1DnvzWsm/zbjwmP4lfuJtqnAKNSU7CiunRau
D1vPzVxvMR878mi2DGNimWZ8xaUkz1a7Do8JunM0cdLwmnu29kifFWITqGkrPTVK
NeOZYcFjg0DR6bdS0kDC+UiFmRShLfvkMyyZ3pwvU+/R4WWx0o/zVx+rfUlAan6U
E7+KU0OJd0E73IteVXz9y5DrMaF+qK8y922uKxBZBP5klJZ1Vae3cj79M8uS8R7e
L+WdCAzmSw7J+Dci4wGfVcOPoSnwdDl2xPpa3dudC/mV4g4I4lxpT2t7NuiuVbMX
NeovtBqXMkew44cbyKZt/9lURnW8ezg8e8+Kk7eVmIYoRbfWAXnbJZky/nV5uJlw
6eCLq23aFv4oVT+ghkSkIpbPIxqjxeEiaysdiWTGR9P9NfyIGVVuspZE35oHHkwO
Nai8/gLd9zXnLBDK3UKB6ZsUWpjGWUIo7OZCZSWFa+YrN5P/5VBLjBhbcq04/SXy
14vsfMiyqlR5M1Gio3eIrCZMntMOompDwPbR7qlaldfCm9zM45n6xe1BuKmRKJ2S
0MO5m5n4sCdfN7UcbcdNLR8SVltM11PVenZzAStVhvDbf4Nl14OLsnaq/MLpdQHm
DWLJUncFZOjCvTfYbbsHrzPZ1DkrX01iaVRV1JapLPUItfdVNbSt77txCqIgyiZ8
zBnz1NOAZbMcg94WuodF146vuEsvUPSU7PXiStFyjaKzBfGOXe2eNb/NCCE7aR7L
dareS8Ly7mC57YHnXV8Y3nYatLINBMaB1uN0vMLFuM6ySv1hfSw9juRAb+VfTcTx
6OXOBA2xiqsRuU9l7KZnh9ewAyDEvyky/0RMmbejADYL34qznmki+oQUThWL03DP
MPEhCMSSZlQSFV2HmwzEmKb1VLhD5fizXszqNFFTPRD5HWFf8AWgWGb8UD3iG1U6
MfENhtIrpTXcO2r1hQ3dg6A91Oov21CT9oeSaE4WtpDKQEmsp4ZSbgOybGpImfeA
tP0uc/Dqn6jzMMinai7F84P1ssw7SA/s5JbXv6BVBNXs1GCeNA7qzrUtQtJn6DLf
qljAEAslyOkN5gprlOHP3dROivvZeiRBOGm4h+IUtVbbViOdGV9j7K8KJCYiSvqb
EDuo0r/D1dSOkLE/HGhKOaYp/CxsBm3kMuR2dL5zLVCOWPHmYeEQ8Wo+J2dcjadm
UoPN5/cxs6vqBW1HNDGG/MRtjq6MnHIrs0e83Si7oiAQiFZ0Byj2T0/oTviken+C
sELM2od7IyBNqGcm/cb1nPMTOASmbEb5eNiFeO8LZT8/tP8oxrwBdCfS0wqnuP3Q
hp6hMd4JflX74zsFgoEh8frv3bdMGed/rQzECFhozA2JmLmU4asT8c1Q4114veeo
eFOne4hwgO8/4D6rlNG+jaCNSgnq0p9AxkmDjZgumodetwr8hnI3n5bW3E9omUHi
GrZdy1hNMUjx7IUFLXtcpLdpnJjxdo9icuwnmDjYeWPN3AkWgAHAlE9tLoPrZy38
+wH3zGdLYmhyHT+RxNRb1fbF1GmpAgB6I9Jy6swiG7JXb1EYrabw+e0rMLYmMNKB
9lDi5xFaF6rd1MIIT/IQkcENtNBzrXXUl1mt9u8AbzUKVh8+zZ7ItagsJmRswybs
NPrHZ96nCWe4JmianhqXOHhy65DzYgKsWJvn6uPRBMF/MBZJaq0llwCPd4RcWxQ1
9+tNUA7iQosmJLmTzjFGdasbe6Fz+w6EYe6tRCoaJUy65+HOnJDK5eCJTy8Xh5kQ
bYFWX1R89zfwq47d7cKHOsCW6j25faGWDpvQHj6HOi/F6kwxW3+F7NA1kjJiofYz
WDAWudlr+YMQLpkDjK3d5zZjVtD/YV22brApv3j2I9AT5YrbcC601BseWRxZ/hER
S/o7x6wtEwZk0DakKK31RcWKFXRqcNWMzkjOFkRhuCSvXZ/OJJsRdrk4CvHr1h3z
KcQDr54GN3Y3q9YoV2bgEDUZZoA+ZILslC1k1VjE2h1qyReLGi1akZloJfpQ7RLD
ne5G66iL4GuPdhwAr6oSybLgd2N38Cs3enNF4zL2d6KaS2mwtbOWfB3uqL1QPDL4
DOihs4Ed6xiQWlSRg7pvcL4sJ7kGxK9aUIlJzuHuzy5s3fkBmARV52qkLDmnfNFJ
YQop9m5/wDbLjPm04oCcsdZ4PY2RWDD+/ai2GxSFBieRCTdNixXb6WVhPiTt/irM
6UFksG5zRG3I2Lq6nGdoj0G7p+Zatix5Mub2HElsYbqqEMTD6h3SYlIUzfmzNHXx
HL/doccsy+C2bJM83cRP2VJZheirgIFXDMwdeJ8FWv0X8M6+WTCFtORzkDs5Y6lk
AFS0M3VQJHDig7/c5MVXSDOP1x7XYDv+4b8t97JEHrg9IRut0jLUO4fLloJgmipn
ZKS2ishlLfM/5C1nQjPPUar2dc07GTiP4BQjRg02hbgY2IUbyswmsYIM9L1RYaC3
VymZFAok4R4Guio6bf3BPWa9+b4D+L2SI8e/+ZHdKE+hXsaqu5uwqPggwChuQEpL
7Kw7ii/Cy6JQZydc/M8umj4Fk0/JSfPnCBVMvTf5xuaqy0aQ74laqnLnZXdxrI4P
1K13IPTVUNVJyBIftj2dsQ4NpAEhzGjA67C3x5142gvs0fpoA4sJaDycsnw3oaiQ
luiGVRoYmbE4YbB78Wn+S5UZqiF3pwMnoUFSbl8zmz749uw94yzP0tgR/PisU1eX
FQ8PtTTOwYFlSWLLoetF/RQq7k72WVzromnTYc8CJIrBhmEhVKygpHWllDjt9xNs
q1GmQoJZD8U/mcZ8UZg4ts0gJLHc8OwS024zW5Nh8G4PkvlHv1hOoPq+GG2UEYSH
rvX/CanoONnxvq4x4oXZXhuiJcZ9sosdbSeGt7t0r1TIyB0Oal2pcvbNuMnJj5iv
9LocOJ+Jfwns7hvOnKn4E/Vupblzfuh8z54yA7nZ1KqvKzBmXNblSFK/fV0eBva/
k4mI+NiMmHxtrk++vvVP2uc7BiT5e40RuBVjVYXGWmyxBhzANRCDIyncr6tMdVfx
3oxkUUhLH3GAddlJWOKipQfpU6hxFxn7FmHdbKxKtZksRxv9uvkVd+oYOtZTTWqE
bM5uxPgcUjLhjiUqaPiZaYHnCegbUlaeF8unpzRS1AO9CYxDJOPPxKhNeK0DUcuc
HdzCjnFGNzNwMr1s/6VSmNKpkOU2ERb/+GH9Lr5WtM+rItIJn6p3k4ItJdRSzM/c
Kghb7K+5SpC9Ne/TPkKt5KPjM/JzCJTcm0yiIEdOBQh9ZOI8yDtOcV0aao0bKH78
OGg/3Img2qFfIbPvvjglq/QWmUnebnmKc4WpStDwuA7vyy/3eEN1mCvlLNtUFiIw
TAmI3iPpVuqnlvPAZlWMi3GBbc/GUahTx9Qv+RdYXVYHK5cQ6r+yCgvc7JMQqT9k
OQ9ZcKaDtWJ9J1pgXW3A0+7DY3LS2qHX53HMNPW8CB8xGQIaTAu9MCmnCE6HoD9h
tKMw0fgCTgZ1Xu8K90KbHgoVMtbU5qyxemsXlzL8Ju8f8jnpqSZ/mmtcjik3gZ3B
inGrmxzNnXlln2nEekACXGS6COaS86Mw0iUDnr0Pzd3TaLuXIFiOdSEXFRmlJq3T
qOPjaqYPkpT5aNWviJ2RSOaZQSvG72xNja/q/qhhJkheJfbd98jXvFduJGkqWS+7
y9LzfUxJzAeAM94UpVgQuH43AMDUn3x5FIiL5lcnruU9Z5wMoPEqMRCxELrpzTgm
HG0cJCrSP9/d5KSdephryUjxyZVTSrv32N4gx6Z9Q7j2/SZLfnaSA6gqp+UaS1RZ
Ke9qoftuVkOgbyY6E+odXW6Z6tZxSfQo0OKnleK89mKlsOnF1wgTs29ZknyJfRW0
7p+PhDbokQDkWbrd8a/J8DdenSDb8yD2FFG6ZuGJct6bquAhJSj0lM9noEeST0M0
ON5ZvF5ni0GvFv5mYbNm+q/L83izuFvXTGifp5V9W5Piz/FANLiCNulGBGjVjyZi
8XloPT49o1TFvkO0rtLMlMkboSZM2oLGIbE7eaK4BKtF1Z0RtYQdDyEZVZk2Dsdg
ekElu+ilm2INcPyw1iP8gRy996bY/HxGpvnbVMqtqLydSaaT7xpqYI1uUhNRkJB4
FPU+Unk5nJQHE5qzvxcgvR+YluKgbSjvXG/jUQIW8zWNEebjqiQlr3P6Qof+B0ZB
p3GdtKfp/CJ76ByniY+gzSeoJPz8GRP5VWsgr1zmzluY15L9d9CJ/31YLrM1DJbq
zrAOwzmziCqSfA+O2ewsDirh/ixgX8960/T48cHyiMab/lQ23HlIfPF0N6zRc9xy
v9+ZJbDH4PYrEWG0Ot5ZdJdnaRF5VtKTRdTw4WG4VJJw2LhIx13lYrKFagHaJ0oA
ZuonXVCCtvHWE3fZmF2v+e/W6Adzyk6Xyyt2rolnW4V73PdCLNDUrrSHog4bEiWJ
nrQfNL+EEcs8+r3161THrF5BeNV5T0XNFaDqKiCsY2Dfh8bJwb7VeWAcVFNXs6wP
3jc7yw3N1rVnVAiFJ/XUH993SaxkA2t77mNptRwo0Xg3L1iLB7+9CirjuRJFYN5r
1rAiAzG4Qg72B3nFNPX1qIzjLPOXHaPfpTlkcIapS8QiatIwy/yadiSSaSeJB5zK
jK2PbJl4CXhJVvfE3HGFpNUswOjcyI22T4QWVnu64ZQhTgbe9S/B9BEN+wXEdzA3
6OavOlOobS+PnTWI/V7Z81uhZZc1RZeP6wY6BcAhOKAmMV0Iz6SbbFgRXqXYNWq7
dmSe1NbUe7+ATHaAQhMXBspcKpeH1dO+JIXg0PmdxvuJJunS/a6Rmpx+hWqXkf5l
Xh1C48M94rM6ClF2OM6F1m9VuIgBIKTLmOTMmC5uRjG+w4gLF9FLk6AXdUAAEWVI
mtayZjR/NnL1/7qmOf3wkiaVUHxJVhCLgTztVMldR6b9fcLAknDt2c99VwOFqTqp
Qz5wHbJ4U5LNt3ReXTFpT08t40BJrFew1zz5k6GARA1qsDhIhfjp2JLEXVj9dZvL
UrFJINaVzQVan+wMF4NDkt80j+4fCnHY5E2ghgRsqaWKJIdYfBHf7v9acSqgeTVU
lFE4+1AclO6fSsyf9/y5IBM+23hJdtVGVsjQ8uk4yhXG+Z94zUcmSksxRTX7tu2i
zgLxHbm+0p6AiPdRW4vDOLGODWOCTaqsyZnREoY/1k8li9/XGgGTi+SiTLWPnPLY
5EwmO4BE9CqfPUSIsDVoIlP/pOTvbIKX+vyO9BPJf1K3gTBJ9CAu/Zdakr59xvfq
nM4Obdlgyi8YK7jNFcy2cBUcWXG2UIHqIlW4OL8f/DSYqzTseAeJKZ/Zk0hNneAQ
osrh7ir69+AF4k6ePfRd0U3L3fHLrbeOxNKUAOfDLMirQoXwtWDndT1MIAFKogNj
KcI/0C61AjaqCLVtXHSXRc+u+ufyQNGLYh0vh2ZeyIxKC2uw49LNgdbHeFv0OUjr
9RKmVHR1nRO2jUDCFtFKAn7CI0ZqgruNCGlwdKSEkk/Q6YIHnztgXcvFAR/zrUZy
JbFPU/hDq93HgpvUguYqvnnRVmR6yATDKo5eR7h6xPGY03PhZ0v911a71wH0WrBy
7Qghj0NeVQmgsnNPEjVeWGvLYEP0JW3xr3XZ1dbTq0U0JN2NuhB79fnnm3l0k4dV
U3Xgy3qk1lXRwjBoueXrgUoO4GDyae/dKVq4hKGQYWVxkHXD8fsncvJ/ds7R6nPV
kTX8xNIoWBQ2dKmc5Yzc/CkTYwn3vx6Bx/8RtriANTaf4Z2GNviCJVZRR74sODBj
dw6qU8VhL0p9Ceme33JjwT1+t83FsM/pTpJ+KexGxTmRl7zU8q85eMSxpBTq2Wpz
SwXURdWU6bLK2qEvIwjHC9afsP+h7AUJL5nFVWTEanBbDIuH6cbHwYArXTh8FJvn
j2GnC5ifRza97DwPnJmkLh/NHIQr+0D61f9mmoBzbYjozR8DVnspO8oWdK6XojtG
Us043lBKDrY3CGdqU8HNtHjA2Be5G62awHgbO+CZuWicFRBmcNWgfP8DqYDJuQa5
JeFmdgdfxZBEvtr/mfvzGtO09hwnCGWQsWQ9HFMh0s/WhhJ2OS8RGM9YsLHJtppV
IW0/4QtAqNKkLxCHRLc3fDNnE2W9IDq3ItZzfh0QVj0NqMox+US1MoDoRVB9SGGV
KCmFtelAGcHbwhWtdgBMzytz8oMV4JHh7scRCisuKmcX6ydxDH28b+iONFii2CUe
ofEDcQrfN683KBPvjg378mr8P15/r9JJjMW6LLIHEMmK+hzVzvjd64jktrJAEkOh
DqgIgKpDnKPQ0gwyrPmj8T2L37q2dZ8M49a7rJy1hbMHmtorHtVKD7gUi0C5zUME
Isb/Wm1nQM46jxPrC9UrCNJFItW1rZ2zDNNOz+VG/fAK+R9MyaLXVUfy2mqaxIoh
vbD8rmqTy3oDEoRkdIT3hzDM3nE6cIBmLPiJf225yjIJogvUHU0zzeL3AoBsUV09
PcpSrDd//mg0TEiD710XUxv3Eqbvr/B1kJDwLJgr5FMXHkZkzumR+ORYz/q1x8Bb
eloufoxPIHf7MDk7DivCfE/VUWrTV/j5dLUsFUGRaktjOCJYQMYZq4C7255kGVyK
lHuFmJ1lRf+eDdyY4BRwIExFMcvgMxiAdwzB4znreI9XoOfMDPhikzuHSyFq+ClS
uonqF35ZZ25lhQlgueExvS0t3BEFB0zyIawWbPD29d2yPKJJYfd10oI3hjzGl8ht
BcDoJtRT7J/5d0Nw/0ddgEul7qTyZuDpRoWZljb2r6KaaDKYSavfAxnNJVzaXXzJ
geTzUG12Xpd4jzmQ+mmxAU/V6/SchjSOuU3/6bPyHwmNPsdkHUkwbN1KIJIbUkSJ
MO7M/5x+A1flRlu2mj0khhHhuG1vUw29j1O1+wik8/eLKFa450agFxj/u68Cb1Mn
ihkIlOjaGfy/oUHmI9NLgrWwj5sYi2IG8GDqy8SyYExhSIQZ+aGlFE0cYAzG6xC8
m9QgLRlDxFeO9dIGJzNKmmszW1EhQwb2TEZkpUr9p1lVlj4PzKfqVfUOY3D4uNMc
jhXeZS9En2AKHKDQNRaIWoXPOqRB1cFa9SgY+FXln1KhKf7uAvXWJRoLO6DWDE58
ni8R7gW0MYzI1EK3ptQBTarMS+iZ2bsWTSTT2OULgYoZXtdl2kex9G8ZMfM1FKLB
7w5abkX6nd5iLNcnTUhapwy5cNtEY8lB1t3eFNSXOjmzG23WGu4A2Uq4hL2fvvyp
+ib8ThjKnbF78m31haVOtmkhyIAhbHX8ppLKuk6f6Wgl9RWZLHboFgW3L6noraC3
2bSwzdmQFsUgD8yV3MNT1mjom8LOJH+9ShoESJRDRg/ni/cWqgpQJnU63yTzYogI
t2zTXJdeKxC44XYdK6DT45Cod4lGxi9yXrL8nkjD/IOmAwz8a8MJixgbhHNiuRvE
VLGQx+lqsDdFE6WU+paqYfipcKPDuQYBzkmuFEYSc1Z6QXugpdn51MZVdwxbzJ+s
2BZOPetptD3tQvhibA2ZFVI2giSCO0cWuxu7GlHGI+JQUay/zZXK+Z6ckW3VQlff
OjhA/+AvN8TI38iuM0BbNPT6EMZHOIGLjU6KIpW7JGsUyyN8czR3WRfYuAhFfypk
dnZPU4RH/aE5oRBAjE72AwcH+Fsbd3+XKpolzRAjBbmQaiT/HMta95wAvKZJnSXD
3NVqEYic1DzZXEQ3x+w1Fi1STYoH4gC4wtsW/vZeHy2OKrHi4C+OIqAmrOv3NBAx
qsM0e7Bv3Mpg76O2xTVHOJBriUwOMcF+NUYdMM+tRkWw/F3G9kYerQZjarzZ1XYI
V5KaW+gJaZK7S0rVSevKEexBnd6Q+moouYwxhpTb8CbWvUBpYnQZFmL1hYU6Pn6z
JdLzDIy/WjtTjVPkPnMFxzVK/jiTbbDFjDvPerPshtRQJVtD8cZXXx3zLG5l8w+C
MrEhBwdpjCuLRQnT8Gb93QyAxS7IV4HbyeHpguh56Bx1JjKyZP8jx6xJap2DuR4s
NfJ2tzrocuQxxEDzTAJLNq4TAY//ZVIZlEWmlSk5GTNllhyi+XRkV5VR+hw1AQw0
6HZ4RJm63kcJo5Nag7v/RaELnlSpggJ04/uJuFa2z6Je439K/x/i1/LE9vkyTSnI
CKPur7gW4MiiuyxDCDb0KhlB55imuzDMIoV+vT2aM1ubGDEUFg+9fZq5oCURmavn
1cl2QNIHadvTbDR5bhZmNUOFu+QF8NOn+e6rydB5HaWtjy+fLNUJ1tvRQSR/P9mM
VfbrmHba4hoCcnUhPZlXVeDIFHC9Lftlfvyg69M9jgxq7VtME4yTtBPOQ92ikPHE
rKHsvijrrdEG8b7CgCw2l6IjLl3IGJ2uxeLm7yiVLnJJ1QInM8OLCX7E/Vh4u8J/
6hF2UvwcgVsoCYIp49CqxcXh065npNBUDyXttymVXgdQsbQ5SE4iHXhCTePeelU1
qWYHHWnpByRP6jocHZ3Lb1s8P+aIU96MW6MUCBj5mVpEaiukhdiJPjV0gSOuheL/
DfWfS5x/fky9mVxxErGD0X47Jbnon7dq1GKXx1JzBPTuOqevptsH16vBesakdyXq
d7TRhJEltr2wlzDf5evhy3GD0TUUHRPeJUKsGw/XzQn75chHyVWYPa5IH9lbkNtx
Ut7OOyWW2kwZD5JLsZMtAWD6BOSX0YwSPUvr0gECk7HHY/xzs8O0LfEMqGHYIrSf
cJBZw/ZG1WBPRjBn01MnvSNLpAhKh5WXijx1D9af7nCSvknSXYlfTscZoyEN3q/f
yw0RN/8Erv42sqO2rEiBijBmLUIIA7VTEss2RO59P+N4G5MaoMody4YZPWERk15u
r+Q08RTszKYHNS3vMYTX1Ft9p9gxeQDo/YBB1spRTUBpCu048E89bv7RVB2+9w9W
gI4dOkmNPJTgbjmM5FWBkCmStCBv07KOCehSVdLv4B3ph2tyVkPCmTS0DclWPXJy
c/i7M7XeGq22Rz5TtSNB9vR7jIJTOCvXpGFjL7b7O30Olfo1F5ru+tLtg3wrD0m6
129Y6T8KOjIzLeQzH9THhf24IHUTk6VbEAHCmUXV3WW1RipYlswzSZvc8AifU/k5
gubWuRK+rA9Bg2gjj7Tzzwfz9la6RiKW7Kj0c5nwn4s/KfRULh6C0LHxOjlcwmlC
bRtKKJqYfiRiE/4Y2AO/8OFtfhBkOncou9ASuoBgashBZu1Fomc0WtaTiwG5QLPq
7Ey37i35tAo6FfEiNHkkAXqcLxrXIdWuLLU6Mha3QprLmh7Yln+edLvLZEu+zB67
NNCeyGXSW84d7PchmBkz9A74DQ9sXiVdu35DCtwyOkbDGl467OrW5yC+nMaSTYpr
K2aAXjxJBvV0mni1JqvtY/ImSix7UTyIJutmAdX39Rd7jChRw5JY+ganP4rZknE2
NjBZCJcYac+w3pneN62ee1aN42KL5r4C14ajFbhm4h/806PkoAD+IBo27ic9l5u7
SewP5281Iz/KRLWFftQdSbU1zeMn3G1sDEcW1NkV5x2gzsBYT/N3S0aZydoCIy/c
Jjsw7CfDdqijL8WEObLcihrAxZhZ82ldFkuvH6Ts1/1ZRGDxk38UstU/wW9Tw7Q3
0SwBdj1CuM6RJNjTrNeaJGCIXaTySZKNTEr3y8U3bFh2lEXRMu6jVOXWlJ8nXUs2
RXaAyVFyAHWjzMGXZS2xJxGHpvHt1KQCt5ukGoYCqPeREUFjcdYkRRI/D2jWeKYd
6nad9/59YM1h//r1+vmepx+4PuBtjXI/qFC5hWtDeUuccz21YOMUR3quWx601+Ee
GCfnoHxl8V4KOmQdV1tKbwunes5+3ranOTS1aeE/zlBsPY7V9g9BMgAjrkZpvXQt
YjT4/xUitH8p8cT1PzaiFXrUbovWen5IshvaJfoK55BNGOF2R3F/YRNwTcujpAk3
Hy1chJiaGQA7B2RoWLu/KuRuTP2Q5b+01SKUhanJKNiEoyorQldOLHdX2a2z3MnH
E5AtDPU9UwZ6GeVfnk+OpEvSEgoc2FHh/ORaU5BeN6wjDkkzP4w9c1EWo4jC/nB8
pt9Smn8htrKbwjNYNoVx89pFeT/cRqx92QSQHqJWrNfOJhv0aVk0berXeFQq1Sed
vCV7StaHxQe4pYBKZ++UUu2Zq6QcIGDRNiq9aHcasqaCTKPExmhXGIlL25yJWoq0
oo8eaIomQKRP8kKQB/r9/jz5LTavEI3vApPHKuXRK/pJbYQiNJzBCcch2xSde2gN
XJYarZ7xpirZvLDgdKQ+SoSndDBwhCM/TWV4F+c1QxNwoL5UgeBljfAMpS7syphy
sxqfloqjLr/o/8HkdrfDYimbQyKFWIhePBenkXgzLZqugz+YjtPXFwZ+Ymbp3eAw
+n3B1CYJgSMAYPphYdY8DZdKtjHEyZj1SjkvMSd9xwDA8e2pxxEdApbZeZJwFDy5
x5q/ScBVZIH3HZ/t4MiBESbo9UNs5QmiamKYxfFqfKU/FeuNJ3zSgpymht+rgEY7
HXd3PdMSkJMIVOXu99YmQm7glIUNl46AZcZaXeK9pja8UsFlN+LJF6/Yw+qPvLcc
JD7yGFbGjTsvO5QkkDRrkbG/yLHi4hroXuXvlwi0m9GaUfSqXwUZteEB4VsJusWB
ZcyCidOtGExj9gO/3AzY1JFu7CFGuwOy51hpmvY+wldlnL9WlJtMxt7uADEmLqpJ
x3T3EYepBRpYZaDsuXJrobt3IOOV28QvzPwh6ipHhH5tYoCFIs/ppyXbBwubTUhQ
bUxSFGbdVE6CERKGeyDOXCX794Ph3uxb19oFotk36gZT/NTXn2aV/h6TZLkAtzZI
uG874jNJseFBe4VLIc6YbmYI/qUIdv3gz3NikSvmOe6SriaewNLmhI8YodwvKhZy
GJ2nfIjuZGlK+O5dx3ryh5X612L+aeTy/ukpjO91t9YC/qajwf3q0BRjMseds3sa
P0vVT5oqymA39Ji/9drEaNgkyeXcXqNzHSwEzdcAmKT7PSP6qtCi0mggOm7/H2Gm
1FEfeza7tXzjbXnRDj/8J43oW1aP2DWcatWyyP6gfK68xwC6mCLzMXBzWOlJdF5r
olBO69p34IogqFDBMkQ5Y9puHRdQNc3jdpFplvLWgetVa9zVbrAOBt0Qu4pIComa
ZRqWUfoYQlIvcoeUtWSwwdZSFerVBU3/Ru8pH8UbJha+ri4tg9qp0wDGwQQfJlwO
2wgTjADvoslg/U4y2TmGNU6U4E47QSd/5V3BVNQvvqlvEPniFd23Jnl/fEvjOLMf
AIM3UBssJ36UDPwGtwwXyyHqcGto7OqJCnJ+FMtHczwL6rISk3mj12lmUpqJAeqD
tIM5A0xXopHGNCQRZ50N7nBl5XsNy9dmSLjmtqMREMUeq1Nr/JcMmyddTK+ASgQA
jOAwUp/pi/O1sxDwnT3tCkjXbyN78dZjNDrKyp3DtfN0fs81ez+wrEHOIH6xitM6
UlWSlLSWMvmPzYG8lJzb6Fb/L6ydvE7a7MZHsi+F24bshgkYeCbOnEv0jkGWiP+4
mgPrAWZyGY+vI5fJkF06UCXIgV/sJMDPp0oTv3m9LMR3gm/y6oaLvrKgXyTy2obn
6A5+p96a0AxVf85eNtRqZjIX9S+nFC+p095HUAxpe1KAgSze1JQ+C/xwj3ErCW0C
p7N2YVg0n/VzD/Nj+tFNPZtG9yKG/XjlGqIL3Xm84MBSphA5NVZHJ0rSDbbpGzLP
jn1QyJSpBHGSkeE8icVIbDnp8UkmaBMBRnJ3TrIrMp04gItonuN1rq2yuzcJCUsp
GUCowyr9shL3oVpHeg4l+Z1jMnDSZB8dJB/c5o9r7rOrG2o+MdI1IK+bYR1QpLTf
udsLrQJYx7BnGzKgfgpSwtrjnm3ScacJD9A3sMDpKmL6QEC8MsVgmZsUDwn2jd+v
x4w1YPsXbzY5bKKfn3W1Lfn1lW85FZPg2zvfifJoxLDLOoGAmtsxfa4ZqpLCmk1l
6FtaxznDYkEnXUj3w65FxZ80C8/kkfaLzdefOXyaeU+eWzuDfNcgP/U1z6JdbO0n
uMdw7h+izstCjN6qD2VyMFUsqzboVZgZD4miSUy25fzkDklminEBAK5yeHu9tulG
cjALepjViwb8KArGv3DAb/sFTb6ioG1Io5bfWutbKdZNyksefqPYCtQ2a1Sg0it3
zfbh321b2ZOWFKw1K0NU/wSLAiov/cvhgpBK1HzbdM19BsygmP/Tl6Dr9DxXukRi
B7tvGk8iYHAgyMqA1K/jFamN6km0ys2S6nX78F+LH/Gqq1GX4EapAOD4zVQD3mCv
jhn2iyKZWS37A0zWp032rkHvXCn0O/u3H0JxkcMXKRl7H3OKEEySThM7258rS5Za
ajE5auBLSgz9injRLKeaAv6c2tb0R9LmV7wLoqLLBeqyy9qkOPxUOtMrhvUlw8NR
s0jGT0i79J2jyc4ASxjqZF+Fgm4lRtDSFhkta+PTrjXidZuQXL7l3naShnJCV1UR
8ThK/7nKwQHVPc3+lb7LcK9XhIE60kvu1WHNFrOlL7Emm5nzQHydQGEpLKLUvCXm
554PPGs4JrwmEMgJXguJq2zffgQj2Ue9Bfav4D93+2mo9l5TnWMmMoPH09WmM0ss
P29wLGW1s83Llgtnb864S0Gx9Wq/hS6cksfh5Ehw2+ShdXVTTOdIuPs1efYgdJYu
kA0d2byHJCcWZ8EYdyhrAdC5KRWXjlnCf460kORTKpMLwV7RUA9Nvi2nABVxh/Hf
e59kCWINA1q5ZUCSWLMGjzmB3QQsPSj0w3gi/QZcAJ2XjhHZ4LVaPuBaw/uFPHIk
Nd5C4zEYcIZr44I6ugJCStqRWqj8rjfLS7HxyLItZBdSlS+Q12e/Glytfgln+OEA
d5UQVgJJsRcUU0jHvmDKjyrnJLZugoU+qt0lYf/YihjbqvSfP8o8AJwB1J8Semsd
jdpvwbdxRNLzKCk32WYEFONkxcj2krvJQG+bD0RTdhx4lNLdTklf5mSf5DI0pZIB
m61qzyAYteGwGH4Ve5pqu6oNW3iHHV2juDCKJ5RA9nB4ureUeWdsqhVDhMtemeLc
P9Fu4wWLeIZwOC95vFAl3W55sZNh/L8g94Gl+k4k+DpNz3CEZ9i8OXxz1qtjw3sR
AmIN3iqBy4YV8tG9a+omJIcPZV3GxxUAf8oUX/jjZzQVLCBdzaehuTos+qlngq/i
UTVKHsfOM1YaGBRbj+POP7wxibEEXIqY3PVML+djlt2We1ZpwCBmOTAKIFa0+Jlm
c0pyHGvcATKAhVnvcuQV0Bh2wiDG2Dv35xfix8RQ/p+A/hBuJ2ibtpCU5h2DodKG
JkO1UgGTewHugxDSGsvXiSzBSZsjJ5mIucT+jYC3L4EonefH2Lb5QaUgMeN95JlF
/OL5AoWzWoemhXxPY6oEpl46g/tokSCLDY6yz4RwkWCg6m6ypEtJe58bX34L3dfB
F+YVE78NFajTw0cDKUGgHQ9aSKIIkvR6I6qTT6cSXaAJpWCRtHfInh+t6SMHood0
csWuIa/3uC/7jh5l5g/LcreO4tYcRctP83XiuXJEhrn37W/PbExz9YXWFrDikYUR
HRUURycHhMWFea0yxCrfrwE2Jhm2lb168vGozXjLHfPLGb6of4WSfxkadxgohK1H
zZoDePoZD6Uq4ULadFJ3m31rk8sQfB18LgesYKR3uXngGWcSb0TTyEPksj7C4HO3
JKKzAI5hUPK/2kBDim1jTxnlvoXfiTNllHe2ZjDXeJsA7Ngo6wG496todLBSUDsl
t7YZsFGS8GRmBr7i5ae2tgIG3X+fAVUP9ns5MdcBldaghcE3cMCveN4KPcHo0oz5
n1shlpUbYVDIP6ylROxTcpDvluVySIJmcTjI6cibtZ+S3jfilVZYOUUXMsD2c35V
zk4QML0rltIzM0cH/NCDMfOcKMO7KdWC819MxyrbBLqnSNuqRmMllFllurKxaiOY
DP/V+WktdFUcUpQyGTEGIMOI4SOXkAmQ5A1zya2OFS3XjaWez+UiroH7tiBWjHiT
Wzpoe6V16eGX11X0XvIQ9w/UMaT92IyeXVDwWq3UuGXnrPS1Vyb/mT06wydgLPLm
jt4zxBvwI+8+PkMz5rh53dbtrSs4h63AWvf4l+Bdz+tZIgT0gAhcMYzRtXb17Jun
6Ntg0qtX8i8zybO6qBBVvHEFPG97ONZ8TgcaKs8JbE4S6P7TFuIPJOYOY+O1avrz
SIW74Pw0x2OFRBoKrJVRqX8qTbXc37XZnfylJwwOFNWGMwhT19PGCtYn8FPXQt+j
czn2ZFxf/K9ds10WogkziL5dGJOXMKFtx88Z+zVPB09Ku34csUKt126EACGO90xU
kzPXFe8axc4lbHpmfHV//2JIuGYvVw9q5P4p5MvWJNa2uV/whV0K7IgQPMv4s2FD
ka8qyyCCvOuKkislGvPEBYPKvLvczEzLkVa3Bxd9DbAEwT0P1B9JpX0T/jRIBFcj
AHcy1Wz0EeyHFCubcbwquMVqIfzJ06qfsaxUU29mAOEix6NBRgkZhPAqalVKNqj4
SepfItz0G0soIDrGfQbJwuSogpDsWoargJNigq3BkTzPRICO1Yv7dgrfS/9aoM0g
MOXW/vT0fRVcJbwXx2WHqtffCU+JchGEIuCIMV51YLbm9jVs3PoC+YE/6CAzZEXJ
OpovrXjJ/L8ltogZ+LH7tVQ33E/bIDwQN0ytsF1XKxav345HIO8pGc6yRvbZHIo1
vh3yJD5+6UtQFMkhVIviovmwDdj5oAcXdGJrEG/XoIGduZT+tEM1qHT8NMohgiqq
e2G86pCEAm8nuNipxT28xxyRf8qN+dE481hjvJOCaDcckCsBW/Iy2uT9Q9eVWzoB
994ZjlnHgCHlvyRtU1AvA4Rj0LgEzbmDKgjQSpZK8OCIGYbWNajyMsPfjZ1ibXTu
RCkTq/zN/twgoqtnYpvImS68pB0+afXfrW1MsX/9KdRonIHjE3Sk0bdFe6Npaepb
ZX1on+8LHLXPxmzWU4b1mc67NOdw+BcdrX4PqWC0Gp5sk+Gb4jsMnOa4uDxVkC9d
7CfOggCkEfzofvoWQg4QPnhGNjAUQ6CW/ZC/5euRo0QqHERjQA3xukwLsTWpbkCo
19Zxu902hMkSluWrXG/Ie2WYCOXEIiUldxny3xJ49x8TJwg6C60n0w02r7ErmLok
EuN3uN9mRX7eP3gCL5h6hlyYxFxYDBtL+hpEslVhN7gN3V8iLEF42rXrQ9uX/WsJ
aaMcg/nqg79w7qfxRNpICBc/bqw/WOD6Q2DSQ3ZmL+L2mukP1Xm5xreIclslL4+P
RanY2H2gEg15HPLTTU19OpQQt+HhWd1DruxBvJbmNyDZ9RyiJOfi5Uj8xcSCoqSr
90y8CFmZb8qSIjIhPUs95/Z60D8x1LEhalHpVbk1GTNtjkCQGL2VmsQ2TWwzJH+/
BQgCSgTqVE3WlNrDVu315mfEK/+myq0TK0eHqm1VTAiH12pLRsLK5/k2oyWDDIQx
A37nrhB2lxr8KyheKqTIuNNA68If+bKxLoSpzd2ks6cRDIuPVE7CkYWMp5TOfm78
DPBeI4UIOUKTXAIijVnVCkF8LkumckPQX8T6REdyMxAzyNPd6+Hc6wDNZWW1/C68
akoUJUYrSl1dU6THKuoKSaA/7Fq80+HMkufwLX1m4LeRrovBI9KTZwoC/HQ9UikU
JMhcoLLzCzfC0fxjZ907cl2sWL8WqzLP4FTAOa2hImQ+XHym2JHulhvDv3MvYZvi
ivtPIiC82d9pPneQULr0HBxAwcjeNQK0Ne76IZ5LF/vsibyODHx7I/jA41ZHJRpM
0zruwuhI6SbsGiF67j9s0zrXyADGuejsbFvOEF0n6v+T5FdwkdqxFbFFlpY6QPLM
ZUDpvirsjj5NvODRsVwxNzOViPiE6a6rASRpJ8eglirD2Z7Ecn7dyQ+NjHS5gr0m
DIIlqoEl6eLcl+g1oxBpFtUQdSzlUHKl1bUwC4UEvoauHIZ2Dol1GEd0RX9nIRU9
QIN46YbgBxcc5Vqiip/t+T4pafrM73KI3E13C1GqRGcIuo71NUo2KMDbRUM+VJy3
yHEbkuoO8O+FogsJYsevVABIfsb6sdv+kldzCNziiJyi9I8P7Omy3Uve76uUr56x
StzK2etkV7qaeCMIZFOg1dbv5KKLGR0cSCXZyq6cLur8mHJLB70TBAezzGJVARHH
SdOibzxAZglBHAyVy0b69pLRI+DsjhSacVQNx2EqKWXGXPsJAvU9J67kMcgFahx3
/zRIt+jNghuONxKR5WHNWKxFq7aX+HGJjF9IzYihiqyA311adVvuyjNN+IQXUkgX
aPcsx2ML1bNNfXlisG2LZYNG2z6+OI/dIMIBt+zHUStwgRExdOtMIqRjs7oNLN4B
wPHPblhRhWqM+6FQJUZ410dR+v48n+brSlHe2oeiRqcUMB2TpsBp5TQfUEyzxzTs
rdYGoA19fq625LFefK53ORp5X42C/Yyy6ThGwoPniBalet3iLmQA3dw0NnQiwVFT
20vYBH7LkLcpvwz+W1nWSKPCN4ALndQe2ad+IFFMQujjxF6Z1V3Ydql1e7+MH/kL
NGrr4jH3M2U+S6wqiqn44LaAtygDj/fgGDJ1yqIrVoohFhxWDMSOj2RJa+6F8lZS
1W/5+v+pBRKLPokfdJRUT/KanhNd9ji4LxitKxcTZV0j8+mnzqLdsyfQpGJEgRz2
tqurhw76wHS/KO9MQJfKZEMzwFYZjV4sG8U1HTUbRT1jNJggs7o+F33DCJQ5e4Wt
dO3PxaTjm6xXWgK7tztYjXZ/2M0GvDKkpd2IH3azHYrnMGHMGaXKmi5si0NwI1Zt
sEmVfr1eTr8/MQdykSD0kE1MiTLgfMo6MWbko7poPjAa2Q7lMJrd8a+aYw6GHJjJ
byUUZRgLr6sybTNu5HcuIziWLY27DwrHUEvWRZO7NyGh5/NXTR7GjFMmOXQYZHzb
S9Y9x6gqxA+Bfomtohue95vzvmkduJRT4KJhEH0Q/C8C8/kK8uJjzgJscAc+aLov
+eQmRgb+66vd+05cNswKByHqK52xXvFFCRWcHngrFj7mp66EXDat/zd6RxXIauAN
VeVN2nmsbuSK28QXNe/D6uSjFSSGXbi6oUpX6uaawanlBFm7asHQtbcH58TOBQXF
jf5f/iuWlc3Fnv0IATUnVbSSVutSs1bFf806e0AOfmvc12g05OM7h1DzYXuIYm13
++RPTsDaqSKLPmL1HC6013GJiT7GfDSKRA2qyC2ZhRyol8AAUdb4HfEAm8Mw0YJK
p3Fiyw2CJUHOpO25eHUf7MSyj9/9qcBOknLGPXNUh2fRtjFZS6GNqDAl31o/hJUk
JjoHazzWDNcQIFZaAUlfQ1Djd59Hiah5Ck3xWEX6SR55nCWO9xmTbx00Tdmb8W1L
dSsFXP5Har64gRx6rPdoXXUfqVwu0l2brTBCrzdN/Te3ri+0eq5CWSHRurS/hgOQ
Q1bIjxIvFRyLYEddQlvWPKLoAMdLWkwvoxNPBPoTps8Nuhk9wl6q63gIknRzNIpo
0vAsFWMrC6VUbvmV/65NCujHbFfzVnI7qM4MEM2lZOpgz+3CGE4yNCXKvNyYkFuY
EfdkrK/AHCm93iCQbtBDBQz1h5lR77ANv+mfEpxmT9EtwtrwFoloAfNArZW54qr4
ZW+0Cs4WJW9BBC+qRoW0jVHHC5fA0O/M7DOw5FTA4h0zUG72UzGwOs3/LetNdguq
n0hXlbjHNYX4s70SBUMCyOKwjBGwsQZ6fJZz59M6XW50uITHGrC4wlkTNLydZnoG
P4gcATiWg+UW0zSf8sofUgA0ZK6MesxQQln+cfhIxj8ZrraDsX1YxGqTrCEWNo71
fA1UC6DLoTYY735kv4Ri9VMpLCXXU9C9gTkyvbMAG/RDTUAcJNLLq8DTwbiawSaH
avuhBYIv2AmJT5Zml/EGBSursXXmzKp9I70uxL3HsbqJSTZaLT8+yvr/at7VqK93
dK1Xfn1guOAV6yXAoToi2UuF/UYG6PdqA7kvxrHCgfsPiXKpC7RJucLTu9GDSBAx
zD3vOa+bBj1RS0x+TjJfe2Rt8eLA5V8Od7rXz4jipS57E+ExvVQEMNRd1UZVrf03
l0NhxhSXaTp9KirRGNRjmCa7ByipqZbPEkE0+6Kg/5wP2HPVEZENpX5A5w/SGs0+
pfBeSJK7MAsPqFCfR99YrB2znQYa0wlpD2VyjYjhhEm+FCYDN4h80q/qOWnNrGhb
+qauczvzF+IVOQVmHks+1umyVriB3L5fItVIpLlQihOtzist/wisQOJExfUwVC/y
sbBRtBOSeUix1oct2HXuS6hIU0BMsfh+E0YZ9K1t3vTFfatcPtOUTr79yksupj4v
luZE52hw/apHOS2PVsUuh8QGIqo57D2HYSLQQ7LVjdzYhDwvNm8wOBZxoIhWEHJz
Vv7meHHZrKut0ILa8h278hLstZK1tZH672jEIwJDvxisD/9fOb1hUSUOjI0W4Kpy
EEL9yfI0qvwjdDRllHqOq44wzdIG0W4EO59GR30EzFPT1f+0Pn9lCb9M/ntt36XX
lqcMgEXXIql/1SG+O5eCfNaOm3fYH2Xyu64Xu8n9zsiPL0hl6vOrXSxHecxNGWs4
2ns4eXGvX7cy1mCHNHn2aSs7MmHFbiCIenJRoBu9HAOGrSPPII7fhPnZtaSnGyS/
SzdX3z08YtYeTbOlyNOGNJE6ojGotyf00b4knqcsQIXH1FV0hFaNe8vMClt70JrN
2LZ4cjqcJhmHBx74s22RkeEYSIpAwhkIvqpR+mdFf9oyj+OlzlOOZIrNK8XDVbiK
paw9HQdhZR7XYvEishEqRZtzZOesto0SxoHQkxaT8g+qVVspzPZrK+egN1w6itEA
EyM0EGs715CNuFbVUX24jujpv26YH1eVdoGUvu3SNHkLBFS5ptqW8N+ytB5DhkmT
TNMF4m+1PMD0is+eFzZk2A6fBdPxc515COHvdwIFxJUYEfHYbXl6I4RQAIGkmiND
CGOtY4iPy1qRR405yvBwLI6DG0O4iTVg34fnLeTLYxgsR8YS9dePH5jx4MnVx8Wi
IU2s/YLW46fMGy7MPsQyc7FfWOpYbr8SapLOaF9GUvIS2bkGRN7AB1n4g8Hh9ndD
oBeVO53ceGBRpddYffgaY6CmU5cRy0Lod07MbUxZClRKzt+ZxY7lvMZBgrg2plrN
Elr6zhVSKgbRJaVRoPb7n3rQ9ErpiOfN6Iqebhjn+21mLY35JnldFNVI1xxpe9Um
wmS8HPv9WTkqqbr81Jm5D2yS+lWq/NnsDCIIQKsSaUbMoZdOV9dJe5nhrM31mGQH
ytF3iLKVZeuDJnBsyi4KwSWptPK/hlJNNDnF25EQ1k2hEiB6Dx5PkeS8acKArCdN
fMbjUAKUDYZaZ0UG+6UFReQD0f5vBk35ZRJDSwGxqqMLZBscCvuYHN1CWVC/vwyS
vDrym8LVLNzy1fE4jZ08j1qbHAfS4PROBEr5jNePfEvDvGciGIQ7uAffIJdXaDta
4c3DByetrjoZQHegl/rv0L9aYKUjr8kUM1Mi52Z34ivKOfLHF5dn66YmlL3zhiPR
EqGVX1A7KxEYH7EZZ3bndIBGlVgZJzwHxoTH15ixU9mFv8Nwk7g+Eua38qHWTu5l
MOwGS3ERDEZNMb3ZBDocNsonxRx/PfFj0sohB30T8SBdoxDeg68kfhYpxpiXEE1J
kS1cwzb1engULrsA0ZSf1lBXb5r6YR8UR3qVBeC5gdHgwPxSNPoljWkIQzV0pq0i
hHvm7v5a4TcHq1yBXhS+IEX9I7Y0querwbotIvoQivCaiN7LoD2TQKRq6jrbhn7c
hMnmZUYMTr1irmsYddfwN4yt0NHc+c83NSwXsFHbCiQszs10M2ECYTC68kuO3JFD
IOfsQCwcK3NXVC0Lwh9dwqRAgnpMAXYP253VrmW8oGZYpO8ZbJZirvZAvaJSUaRa
5tWc5yaXK0qIBl1lv+neTk5yYqHT8Mtp7D/DDH0bwxy7l+7ZvaU3NK2ZgW0vAZV0
xEKfTn0BiRl4tqu/ezUCb6++uAFLJkSRYfhgnfWs0n18dUpp0Yom54HJCgcJZsef
e3cS3kSKPx845PzKPxKufxOgM1/ht2Gn2QyeYRHwVP2XbCfenBg3lmd4R87PvRf8
0sCYn+VUJk9ufv1T5j/F9Oox/Qm4m3iQplCtXTZRUS3QYmLV4VJ2Uz5TkSeIZ/tS
dRxZS9OfwVSgBtFLDrTm3Don7a5R4OB4r8GcW79U3++Tt2RdSm7My754QaZofYuM
TblLXLTYTye72DNrd8owabrMLp2U7xSqqjU5ox/d36I13NwiO3Yqk6U6RcX3KDpS
GYa5jBVMFSPNeLnx08sYf6jE+kmLbVndvQQwqYd1qyClBhuo/wtuXHloOVmd7P9I
YVnZq5ROj9oOXYBNqWPNibd5eh2siPE2pfsfo+bH/2/nZfDpA9iOASMQ6s0yRoLi
hAULyp0bu5WsOs2L2ziGUvg0PYOHiEF0vbBcozPsyAUMicyJS4TzdvcBYjF4h8Qw
h4+gzWx01oX7sxP4d7TRNc9FAm9EsdrX2q2lCws9dzMHlnZAKMIs40NJHsEVdgSW
4I5BXUwsVMgK2HSqXQDxW1bMCtY8JN7bf+EhrklqLg41OIJAoQZKsxEAJ27JCpN9
0W9PFgiWP4ewk5RH6USK925o3uYHLvuciIYfsqPqBUtqkkUy7TGkPWI0rPt/QO5L
joI0EQ6FTQjGofmgbyyiDYDRxSd6p/FfP0mVuL2I6MkO970LLsOZwrKvfPUDsk8o
8zsVqsXrVt346Wp4htLAapNXOscBHD/RbTJStGx/4zpBcOjo9DYxU3HMhE7KXJdr
deNmAk/pX1zPyrbP1QlWKZsmFiGnLe724WG/Ulucsm4=
--pragma protect end_data_block
--pragma protect digest_block
jgFZfRU9MxkxiI+Iy0g0741dtxA=
--pragma protect end_digest_block
--pragma protect end_protected
