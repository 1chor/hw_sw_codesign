-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QDwJ5rd99Tb2GiaBbXVsKvjQ3RgMIGNl8n6m993GfOkeUaIh4HeJfKigKxmEih3m
tGt+5IcTjDtsMfg7N1gSdsUmNitT7aZRb/Wkc8v5L7KGj2WAL6zlbd4/CTAEtthD
2Gjv3oj/Je/zof1/kS+6Cvuu6Al82wcCgjqRhPyBIjc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8143)

`protect DATA_BLOCK
FS99zdqlxv9najWB1Lq7AM+18JXFaayrzndg5Ssga7TnIZIiSmElgTfv9n7vPkQV
ONiOwYU+usF+nXlXxWDhUHVjvVkS/XZKFBEHf60UjJrw1bMVXha37cF2MxYRiEp8
k+McPzZdDEviOMO2+jtvmqcC5ZX56/oAtJkxO1ApBiZv7P1EGl9dmUrtOz1vSeSO
NnRkpMyroiVSK4rDxrGzh4ZALL0ldV0IRuMc3oUtHuN0ys8+n3SnB7yxuXH5iMzt
2lnpLIC8DE99tdgauh9K8nbBjHVgiP/Wuq79d02biabiur/VH20WgTPn0Q4iIbGY
O47/Gt1p/k0y1QUFZQxhKEpTS5gtxmU8V4idMlfwvqNLGSf92/2cHfyXVjXxcAVw
Ik/XuD2ZX+NqxWZZaTUhQLieZhH7kJ6ed9t4n5ehUMTnf8xhXdxbh2+KfrLguv9v
coz/B22a9gPCj8YEzAJgtcGD/Mjs5dxfuxfIgf2NNM0oev1WYfEprTInk4Rc7aBx
CZf2PFIb/2Lv+Ui97Ha5cfthH01KGZCpyjKfRJaYiCRIvEOLDrij2flcltxXWWTT
c7J52xKQ4DZ5C8mrjDwHxZmYEeI8gpMiXvq8LxEmGAVNiCMwpXkgiZrSd7vSgRPW
shJFUGVZRLmtegiK/8eBrJ9Ff24/Gpjyl3vXheCxLLAfDPhyr+SAAXwMQdg9uJLz
oR6zyYts2HDPIZjBcMBeR1fsQLPoGxa+PLm2Bi8nx+MmlDm0EMQ1mXx/MnFvllB+
N156ejsJOVGhfSCTpwYZZ41tHoJJecPWdMYia1hhvOC974bRbLz0+QpqbnE9Vtkl
A3gsRKzOevDaSOB/3A4/Duzapa3B+stVtvnK6Od7dRxLY4HRz/q/IHGTbj7kOILz
LqUMig58zdNx6/bcpKyFmOXR5F2Er39pNeE9i/tPgK9NqTyCE1N7ZgGYmmiRqZUN
X/I/3OJTkGr4mMH+HsGm7BP2NjDJdE8KuC5mouo3zLjKErlnqU+zjxdsWiYIIaXd
2yjx2hRLBUy0OqngaroZCkm+xNIv4oA+k3WiG2wKUBYMVwrD3RF4415By+SGBd7r
T3LHO3q6t8H3DBPWatpdpW1DUJfZMjUD/XFylI7SXLpsS22wxi7JaMsrRHeh86l6
O7UTNxjLjbYQ3czhI2OouexjSo1NTbw5T+9m5atPkNjhN9X5J1EZie5il2/XaKHG
VfXIF0M8Ixf+m7ExOle+RMZxrEXsaAP+xaDGvXlmCPcyosO801hVPSYQO2Lk8+32
syKpSzbO7b/PfcLVwgnoGBc8McG0mYdZSNU9QCeHwHYhmBhhi7SGFqrRyMcm1RXs
Lf75ygIhA3e31R7n2ljCx4YdQtezocockWQqREjauZ4UGW2OIkFRNxiJo2wY5iDJ
jXPlurtGTNypCBLyyOJg5gSrSUdvC+5kua5lNpF1HOVKtD07H7mFofmb2NXxtonp
aMRFbhK1e7sv/BsGY20dfuTYRhc6XLoj2hHSFbvLBweEPS7vvFPVR+6CGGv5lUjm
gCDnadqeMUlmN14whOLR71nqV8SblZPlAiLHwVDnjqfqAZaS85U6xdgQEkF2YfV5
HglMxFzVgnAQu+hA1dIKOl86//5URav9hee3yeyTcxIqPI6mojwuXnub+I/3WmXo
+fzQ/gD+1W0CNKS5t8XW+cp2Rzg0aUR7fTCrZWfWt179+KYGPzKz9opqrN3L3jeu
Q+pXtfHRBZ44mWNZWr3o+rG4VzQDCenUHR75Xraymm4kmDK4ISPdLJLl8UOJeBKN
XwP4iayocyAuzhm2g36CcC8ncsJTycpOsnQWeFRDNh6n3+WHnrq8sEI8jyHrYUDJ
Z0FHXCWHFbbeoiRkcs2IwwkkPDIhoaxRwZz2pplUmhLCxq8Pou9etjjaL7XAe5Ur
PgjiK/QYp+Ruhw5l30tQtRJ1SnVaUReKrhL5QCpfYRWdJ5D6NNmQaPwBg1bkHaBb
7HXgJJJyjOdDVIZnq0PQMEJDAqsA+8nBlzSv9aLOcUovdnzCzt8wB/O3TS4SiElH
GpHytaW+QnhsNDjYRHxAdhwzrZE/gs76yAWU1z6iMmHgLaRJIapU55R+IJYTuntK
m1B9WGIxV2nw+Fa2FwAU+QTefIAYSYCHJ9Zx8f94m4HNHk776pLj0tuQmIil4Xc2
cuIzY1/2TKuTEtGpOvEqQmhIm5LVEuWwhNsoio1J/rOq2DjQaaqRT1PUxrHamome
JgMPwqTFUWx0/ddg6ZE0ITiFafjdCSgOQz1kt4yz701UV6P+fYNUY0WLqn1BCwcC
GQTQ/PIVIDdBxYQ9O0q834rezabE75ynC1GaeiZlFn0N5+sN9t/kO8YRWEfWAE56
CaIFQqs5fsItEq2YvaHoHi7w0ihb6M4mm7cchDMYJEeAIUoj+KJaeKXPLl5NcHf/
vkrDlP83orwnw7PhG5SW2SBVkKdvdlSUe8flklm7wToTV5cRRFTnq+LVeMJJiHvp
wy9lvkfroVweNs6EEI9+28OSVra86eUhs2UikoyT6rV0NkxGAxpXAkVJs4JRbnrK
+QYErzMipa0ql1LsSbhyep9gGb6zoXMPrpkiHZH/Jm9YQvD0RWEI9l4NfCrYR1po
7ZGImTLkTpxgCvGnmuioPKHkdBHvsfqR4vgP52B/l184W0iRH4m4NEK2NYTxW4/T
oc/D8pZl+0EAr2Q7GHgqcFDCxc09lQQhEWk3AU8jLmctS9qNRy031z4b5UxlFxfQ
FHO/Xn3tOITDVy4Rg6xZiP5LLYvkauen7rVGUhT5paCRO/VHkybb2SmQhLlWJIjM
FcBAuVlTapPJXeIolfLME6vHb8M+gzmTFkvnor+jPLZ1qeSG/nAgMZvy5sLqImB0
yoSnbbWgBwv9u5x+1vZBl+c+sgV4A18t/9QKOszHsS6KBTRZf4RcCL92i5wvlNrH
mbg2UorcMZhZjaKBnlctJbgJj54Dlvftms/GrAnI9l3SNzrXaVr4jqZNum9f7Rly
W+/SyaS7i9yDI+5pjHCRM5apBT9eJeP4/asGret63QaIxr7IbMbbdlgjmNZp4OrI
WGpJJlfW++9vABgny6NTfbyNYdxKnDCBY1jBh56m7p3xNjgOV+x66OiudU9oRgFd
180PDkDpKz2JEC508ljGLtUj24Fe36S5iowCVq3OWHK+zjJg8m/jvOPMHX8vjjnl
JoN3NBpgc2yV2eYlnMPAMnKhV9kGr7RcW3vBvOsdEugEkkxsPjWLAL7Oy/nZRQ/I
mWXZStePAH9MpCDUzRDxGXDSASaXqJtuMieRxXXFavh165ZGnFHRCu+DK/BRZVoQ
OLkuKT9EEOo3gUZIm9TP3hi3HZtohRjjbuuMvOqLGK2IKT5O3UgOzLRdJ8QEomXh
mVx3dQaPMHWCXAqML/5lDNoV2DvAK8fZQwZFEct6yD63LFc0wRjct7OP2WNM58Hl
dD6OG4QMl+LNkM/jSTrpd8EwQtcLvCJPI79+uv+rI4M9AMxqku7XW+Wem30J+iIG
Z7fFnFf27CzyyUEZzAzxV9NI7Kh0EFe8NqyrmgTZBH3DeE6IwRIgYyWhi9URg/XP
1XIemF3PjnhnXV5Uvnc9zonkQNLk05gnfEOOEETJ+HGYXThX1KnUzEaNFMAZZphH
VaprO/WvM29lSuHVa4TuPt50uX2pekKUl5SZdN5lTGisL0jBh3bvbuFrXX9mXtwW
OzGjQeK/0AvQd5ump3Hw9ytN+znSUzRbP0lh/DYyz6Nl4ig1hq3xlokeHnmfOEl/
Asm2ap1EeXL518RqiF+hpHTuqathYkzNIA0vreWEGj0MswFhJr3we6iGl2AWIyMV
N0qCNxwchWtpkXJqE6Mur3Qa/zG7ISK2PmgfW8SxVAFzhFUs+S/PvgDwOjdV4Mda
Cd/Cu7cIUSiRd5xLDVn4nnLwOcT5qH/L8pfK+sFH0EKIQAQt+sf28maZsLUZgkZA
phzQXj/ePGrYBH6JIbJfv3LrYg17V+karBV3/a8F95adp35oqahiI40q2RXyMHBI
FKRq2kr4CIegEy/6HU5bA67Wmmn3F8c+0TYZhnq774AoO86uHG47A9F9J4imYpyb
gu5D+Gfp5Pm0KY7LS5EKAKTL+NOnzDZSKqUcoQqJAnFWPgMy6QlgReklEUkcqpv+
fJNK6soAGIUYRixjFAuTaYXNc1rKD1F748y4uDp500KSLHUJiVoJrQYdu08SLwJD
oINKZYsCYWGIGqy8rOSECFuFUhNlFdNZVBZijvWUF0q4ZR13+1b/QOlUXnK96sNQ
5Di9GFxT26n4y/1SREzEl4FKCpn1rtFC+Wrv+qGtVEWiLEpyzTW0KOCDTEFvAe7G
/q3Qn+1UQp16ANUzrzPXNyexLi53mrQvRTvN96xyXn19lqGMdflSu9sZ4yIZNN76
QfTT9+UcHFOApG2d3TkzhI9YqDJZDBh9uj3dv+kfJaNp9pfYCjL21Cz6toGfFpH0
nLKzmKDuSeSBQOJbOavw2qGf4PYgpBYGFrmIyVcMte0zWJ6k4CIt/LxkdCg2p63e
c0KqPJCi1Bgy6riypGpViAuwBcsNuuFTaWRqR9C8lABui1CBRsLkS5qe7bkt97Ig
tTCWw2aiUlmcrqCr91Dp7uAVS8D9298wVeYvIeUEDxYKU9dcrEGcif6/XEw0g/nV
cEWucAwBjyWYtBZo01AIqymiRVWaYnnjGVqfIcj/QZAzE4Aq8IpW4hqtcLsx+GgS
VF6CBtVwJfSxR0dJz8+DxoxoEsXguoKzB4tJ/aKSdpzoIfbk0jkSwL0ht2TsRsQQ
N7cY/7TRtGGVlsSOBHKoXwZzgCaYUkQLaR/ixFD5PTCZ5KTqb5htfD+SJRCNoq3p
WyGYOqDI/sa5shzMk2Pf8G2/6vMm+5MSNRpocSqjxsknAcvv6g2VJh/FfSzypSLt
1tQslEs1HJZ2g35E30UE/oYeA4edApYX5nrQwKpO79M6c9XUR2LY7T4jdOpB7Goz
DPGxe4GysB1zPtm7TKFteypmchqfOMF3DQEk2kGvM5VsaRbqC+coGaCEqBeZrY4e
9vcsVoAV7v3YjIRL9/NMD8CED5xVf5W9YPVbQdfW9B6M8/reHOguHuC89m1q/bDo
w9Nrtm9necJSUdx/9yWbrwhR7BS55zzGRuaFwsTURI9EdJFbA3IxeF6Cli7PIT11
65cDxNhGWCcqls+UxJveyCIKK6v6rcCEi+2A4D1d7Bcd5Rtbs+qdpotDyU7vCsdO
tRmwSIi6fubBPp4coZrztxwScjDhoGKXeyHQ45Uo2ZLa3X4jJjgH0bvgDd/C9h/N
Q+85OJTXP2pCqoodzna8gZxC3bBE1vEoerc7F+q3C1b4Qw0Ho3Su0/jU4pKay+1d
5vdOWyXcY+gc7T968wk1tXgztzbNhf9bXneAp61FJxqMkJgS/PCfmZdkkaznCgpC
NMcUeUWp6sGgqFtQKU7gLsbb+HCXN59UN2pYzLdAq2U5Gwp8Mg7ownjN/yYPsMLm
Pv6MHDYpSCvxETgCCwU1YA2h9jyhFXo7OvWW5Ds8IlRMOUk38a80JCgmi2uNG/Uz
L+OTMgj7oyrZyvUTFpO8JzD5QTh1XePZI40tT/3e5rh5L27pV4yApYuqUgb8Vb4R
0NEdc2d0SiCFkytKhcrmeeprgLcI0kyvtSpEaJOL3R97xRDGP1kF3EgXWuSzquC0
Oto6AI7CpKqiLGiOEIR2UwZPrRaebBN8Ulmn8djAajxDffaiAEv9laZubcG92zJo
4hZgGRs4AAFiDE+GoEWYrnIPVfGewrv8R4ifvkqy3Fs0vitWPx1nSInzdJ4Cg/2S
bISstGUYm2WnmToy3jjPFKzVldQ5LPJCGZEYr7HqQmgoD99wgzdPRrWVdHfjLVZs
Bbwwp5hc182BOJlXcAz8BmUnHvuq19gP7b/Tmigem0GN0e1zJ2qtWZLXw0B/fgAg
UIWQUAstjQkeTKNd4YARZPwYVzQ702f+AaC5z69XDReG5XMQPGVjI3pFdQS9AzwR
puBdJ/tW6t0hMSeppIbJJv512SbRjx7XcE0DH0/Lwu9wVRVElcyPtJ0YMjR4NUDy
SEzdXdOVtfymLMru6UnVIrPA+ocEKmT+rzn071+GpTfvWHDbveA6iRVKOYE0l3wZ
B/gQD4cE7tj512vGTihLaTMffGkxBVDCt40dyPCcE+p0bWEz4sdOwUCpZlZYGDsF
pMGDCV5VuDCsmzi/vm0naIpbJyf0wf9lKnE1FA3B22WOldG5g5Wt0ajaOLIGXybm
Hk3boRrpNX5dgnWAYHwfPAHUZxuiywK880bCLTlo/BDFhUgqDOKRr3jtjXIMyDc9
o9Brn5O4DNzs8Ycyx7XALzt4jE5VBON0Rz/iR4VEtvpKnkH5bHFYg9IWc7C1TJe7
CE1060kY5XeX4k3gj/ICYB5I/wLu5dX7Uv380TRi3b5dwkOvV4i6sPXPLypLH2ru
byHuY7iGAEcO0cUeygEIuypk9H692s1AF2XKZy2t8DVyeuvqo6Y5natCW46XJstW
8Xt4JFdRompGViQHw9D1RCwZ2LVctle6aWr67wmEFi0E27NNoU2lwZ1N1VSkN2OA
/p49JMTNadM0FhR1uBin6QPT2QRhJjkKK27Tde3fj1FS8PhT3MQHpMvO8iRIxfK3
Ywp0nj8bR3b+6NQQVebUkJ5dzLTjgNN/4TG8/b0BCI/JCg0xs38Fm5vAVgtKyhiB
BS6eG0K8OuHsll2bGrxpqav5jTfVbRiHHs845c3z2XWIlUIv0e80wM2jepuJI7kI
cF0yDNZlyyAq2W7h/a8OJKRIfmxefBApLPcR9GFOH1rCrrRoaiklA7fksSMuDIWu
xabwYlANFZGLKWGT+aU6aG0WKSM1mCgJX7ZfBYmxVxGNnORtTdljXEskDH19R3oZ
FJ7Our7tgVBL0FGzFuY2iJvTs5HNIcirEc9zGHPggcsVkANgurnMGZkervz6aJyC
6ISbLFYa1JAmbWijBeNUrYnGIUI+lTKG4f5rmNbReg6nX5+XygGRffwIhOzq8R9V
xYzcWZK8kbByE/Si5JUiPt6d26NK+chKqdqee/JjOUNu7U2nz0ZNvUYV8L1VBAui
iSPpg/u7nFczUdy8vu7hZG7ozVh+cGOuB9HEgqfaKuYiaNBD9lT7dEiYhSU+B5eo
JA69ItfnhXvpl+LbgVC8/PjehzCKu21jSQpXAecsVCauoxrM7skJlT+zVQI6565P
uhwpuqADJJntIUdVmS3ZvA5UI1dlUosTsD4RBoRRPJe9uz3pklT7NDb7IqLThSD+
2ayEF6py1ssQCtkEsMDIvIn69D7Dg9yPWCAUuZ5XIVWuMB6KD0g1IkKz7A95jI8z
sV/Qrc1Y+pKnkbhDvdnSNqyArVTJUcSkZKOL8qalWIzA6MdB4c6gQHh+ji+9TBxS
yukQFl19fPRRETSVmQC2MRneQ7sizWPD71ZK0mo/tJoy+Y98Z0q0LtwN8JlnBkEu
l/oBIuQT4Fc63nWMkX35i+ELQLqw9BAdKR/c245z5IAFr/uZrnZxPBqgyrOwZYCN
D+D4aQ0lhRzWTRDcAjAfr1JV9gw5VwFQT5JnHF+k+FtvdRmjw8msC3BLMe+PuU62
t7F0JwTu3Ovqsq6lfXj2N1IcNnltBFXnmmSx9KvQqwQsFEgAX84lizA+nqKAM+hZ
5RnGMuTis6dP7RQsjIPNpL1vCXuKxVPcOCZbi83q90dIdTh+4TR9YhpMCkLBq7QC
DTpOHtMUIL8jEk4aayD3OOcu6mXTHzM3SxCf4RBWFnoI05ZubfMW6s+YM6l/Fo8S
R1JxX4Pndd9s24F2mNMawovT0if1iV1eF1J07gb7gBIDYxXBQvoZ6gn+vuMyAJiF
Og95wp2E/xiwDLUaRg9SfWNZDFYdU2CLiftK9Ps5tET2BVQsjyxPnhsmtsD4wJq9
nGsag5nWvKxWTEpxlZPE6q3xAgdr4G4ZFy4hePokxvVm6mGvGqHgY6qP/OROcNcx
NjmgepE35+jhNICUpWym755+r8f76PQ21SQVhOl6aQkInTrmSHVGHXrgSedoO5Eh
Snfv1Lm24540qsbpO43HOSaO+LtfiVt33C0DGkk0iOi4gB22/+nH+OrVOBPlNUJU
NhwrNJjzomHnXlbvi2h+4YyS1ZYjdH2S8b8STGaEi0PhKU5Hx8rag/hHHY7ONtq9
PWK1KR7yqqZvuV6xjSjh52sevy6uA4MMlWveQNhgwAIx6rRwrku88e0AazGwzGgR
GcqR7YKmDuT5oRmcUeOxokpLhnGmWp+en3gzVCl9y9qhAQAWzQxPOJuueK9Tptxi
jI8kMTyem6ytGhmIAQ/NSAKRUWGoeWwoq8C7h6fxyIqtgbePLJ81FmfjmwaQLWNj
RQcddXBF9tb/teC4F1EvR1CLuIKfGq3ZsQYuwDFho0HdjR1pW/eSDmZZmiiwvdyW
0xpZciushvILUeLJOOB1ckrC6+mMimAOuGXTUdY2fpOwgR4mtvsjGm8Wv9GRDP2h
G+cme6xqcsld8r54sia6ZCatK9pu7QJZDza40eyDZ9JhW2ob8At0vjuJHRfzpAJ9
7Jt0aQB7dyz0TJu83R0TkEcXcx466PoiJUURqhA3nXz56cWtm8OlHg1O45KhpMzq
01nYPft2NeotTaqc9pdTMIPhsja8Q1d2Hi3qdWDS1utrr42o77H+VJXPUAbxsjjh
wjQ7L/l3Df3+gN6ojULJjdY2vMUerckcUGMQoLJzRMKIHj0Odp06i/MAXFevSfCX
J4EyOpHQwLviO+ceI5lnJqXFPZA3Wyy8w0AA0QLS3LhR4CiO7ZFctCyO7Uwe0KdE
FiD7iN5FPluxF3hHjHqcxY6SWelsl1kzqv9wQ7KgUMNyjq4Ldz8+2eaO8+gilLc8
hA1GSDbUtapP7SUoed8zEbWAn60dNmYTtvWi/GAlqPrbpOwFlc99mhzJM+FlbZs8
2eZmNIAd84DUVwJMIiNSidC40hhjbtaFeXcW1uHwkQ4YbNDxv201panmIFNMQ8Uk
4lZsUqpujAsNnAQ5QigX2Y97fZV0B82apyFyLHGkONu4tnnXb3f/LPpoKEs1D2DP
c5w3c1/pHE6ghdgTfnuiqaym+XvTWHi1GafbndI2XTSmZetHA7MLxWl6yeCCZfT2
CCuFDhohKdEsLz9mZNSej0I6kvzGwtAxkJ8d6zN4THQ7ibNN34Xqdv1bHI/Q+3GJ
7JB16C2SZO8x5CRmm+bdAvv2UbiCKwichme2p819ejO9l9XQvSP6ZNOXNzHDQ3/E
gkMW/bvnkC4NkfSLPz6LUvEZPdrcA2OiG9Mo6ElI+dPBnAGrybO+IhljDqCsuLoa
5GLFwqlkMs+yQ507cQzxqqwzBeqYTSJ8D5tpOk1aSmi/JoxxX+vrG8xZXYAqA+TI
vjTJg/Bz+FwdThamClg6jbgakdUlwWvAhfCty+PzJladqfp7FnJgz9opXJOFs2WD
moIe9pqBNtuM2vkTN2ZrXrM02PHxVJIAkCI5POXLDWAkFu8oPubPStm1BMylx9Gs
FOtw7GC+48BXCw4cq62nK7p6RzrkoKDnH5yY87PCPeGnnp7V2hKHWu9n/sl1+ALY
5SbfADjdeTwLC5RG2uO2Vn53ulFuTjjcKtstB8gIs2Ko4cEFsOPHyHvQkbwvb3MP
UhLyiT/JdESGnrcqqSjBg39BWlKLqMc3onDR+FkA4TItoXzN7QuY6xFJQfzFp7OH
UoTs+pHbnlXYYlmEyWScE/DaAMHssRGoLIXXRlKNMpk5TtwdNyjTxdTaFG0Wt0qI
2c+g26WpDSExAgd8ZKlHVw7pNkLzGPF1Io59Vo6XiBuTq3LaIKE9RGGUR5bl9w/n
1KsK6vBzbS+sXHIsEqABY2C8PHnSMLVV3Hx5hNZ+mbWlq7vgpU6UyEtLlSuvzI1W
LdeLlFZdbLnE8EPxKtoiGeXbTSt3MdemZ+/Sl/kuTKXoDgR/oz8T84Mb0loBuuFg
jlH7yiSepT3gNIOG/b7eoipxPcSeCGi4aQQgZo2uX9pirQhu1dDsHAjO3B0CT/gR
/jYCRA2D9uSWKOQ8GGoAmkr813BqmccKsqVCdA3VA9wvj4L/XXYoQZhl1V0tPN+l
m+MFz3iyv6xxiXE3o4i4P00Oq9afc/9se45UQHNYY8KpO4cj81tjcD/JyWTNpTQp
+sYoQV6qQ/xTaRCcjVE4jWvsuKM+aYBrBhWG5Z3TRaAGIScbCOG9seVAw9tKlPbf
pJx5Efd0nUSQdHlnkCXpNg0kmqSYaACIwFvouxTqvpUsLkDTIQeXPf28ZnvlJhLh
pPjE/ttjnxDjrzyKgWB4JIZcikpwxnaK6XA8yLSJQzbYMGrhEVuLeMAGevFMHC1r
F7o5TN0YqclZl2jE8mct0fkC59Q/bcgRAs02YtmpLH8VmCACXLWT7npVYle82VLL
ZE2Zj0Q/cKW+ruG34BGaCOQ1ctVEpSlOPsypDaPytoVbAiHHx6AqK6JU2BmNo21v
2eaRzIazIAgpahRH1A3S1NYSPtbauMgI6iEOeuvNw7rMU+G++6+Rj4ougG8MDIkG
ngSxhKFbSM01yJwBsBN8oAYh+38UOlEWgxdxnHbg+kJ5W7gmwec3uV4oOg8LtPKu
wLTMI5WRfyhncTME8Gq9lJpRFLs8oWfS848eqP/8pLkcIheN8LH/X9c+3Pwl1UhK
9T+J6+x44fvRSQEFTBu5kO3kiS9A2JqBoDi/qjD7IS5vtSyBo68F6uxhSnsPtBGF
9vcvCkoKMggqx99dX0IRRh26rdGwiQ1/o5llFtFZHssx1pNMvo1mkPTv03JrhbbG
VD4FQxP6sva4MDqA6HDAgbJ64wlnLsEPY7ebJx2tGqDS2JUe3DyTJzNYaaq2rxjS
`protect END_PROTECTED