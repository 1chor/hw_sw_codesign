-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
RPVwBiRk2IgM+P+TnjVbNS880+YUZcqF3BeiealhEF7KcTbrdHtP3MyCLetbkdDe
1q98q4XsLZg+rXB2Sdde9Tgnhak3LNjoywrEbnA8zvdjVSak1Hcltpd+ZRmQz2PZ
ZDAR0wEDuVaocQQyXAFmkwxnUYL35JlcikTpKIbhzS4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9376)

`protect DATA_BLOCK
Gk4KG5oH3JV30b2yQ6+oqJb8GfaAd2uU3dk0Ean4rz2ELZ+ACUXF/n9iVYNR+JfE
Nebx/O4e/GkzfCuGvKhA5ozVbOYWCSdTRK9JjUvVAtY3x5J8S0ZSfLIzhYET58xZ
4bHdC/77LlEK7B9VuTaIgPqWrUYOd3DBp+nEcFjT+rJk6QsRXg6VTYh4TEgsvq8N
gLejol1pQ3WlQyM0+qqm+Bugh+SDUZeBrN+URxwQqMLUB5VUVbwqhAgaeCTTRpEg
iHOCozNW2IgxmhwaJ8qkGgcsiKo5LoBU8kmJFfmWkKpAEXQ1VMto/pBTiax8wzNU
epfVsxs6zSfK4ZFhFK/cwPsRS1JYvYixr2xYGGHyxzJZavoGHTeys6oW7tbo1kWh
ybuqldzCUqeh1TjLM7UkjKKUDrler32tBxx9kwyZE5VGxf3LWYykr1s9S2BLtwIg
myPkfnnjy65sSf/i16eVWf+4lLT+BS3f8PeAWD4xpLX0xATAexarFtxEVkfe5V94
pkx+Y6WaM5IuT2ARiX3cUGGH1/2kzFXzhk30qcmYcNMkMlbc63HeIUXP/FDCVoWA
JtoVkXXneDIOccCqVkOsJM6zgow5DJjLbgJ7hbnUUlhbFNhUToT94d+YCPlnEjt/
mGePaKuxYGw6LZKPrt67bMu5ZnPfhCelNGw4eVb/zESipfYUZrspaSRfoEXVpde/
GG2R6NmIs2EJnFCwhdfMIiWjaoLDV3uVNBRw55Q08lmsfumkBWr94fHV9gciqA85
cK0+9asWLOiAYUTuf6HABGrHw61H8eH9SiH5wJCmodj2zrvSOZK8u82gX4sgn9vd
9zaCpCVb07SrQIiq1JrfwAjWk+JlQKuFajWJJzX6RAFu6SrOYq4DI4v4l3PDdH/f
iKAQVzCS7zLwj8ht+wNAI4WxvXmxS8TIgYP/gn1ZYl3INv607f+3tV2fFTt+bWgx
6vWhgPLqW22eHgBOtO57Ux+ahU+9ZwUon02cwszSWvyzFHikZkceaZoIYN5kAfvb
0mxvKI+2Xd3luPkQzc/gorCfBxw0zV7Xx5TE9SfO/Iu1B7vcFEyr1kLh81FPdsxp
1Qb2BvthWuPedwThoWqO4GGRSW52fNCwhEnk5z+ecaOKJkaMRy8EplCshu12BdBX
l4hDj5OIXZK2Vp+iazW+3Hs8pqu5l5m/fnisKn2WB7q1qxSzpm9tDsRYkyxyDpu2
R1aUA5nVvdjtSptRxYonz2lGvDcQ5BSfS+sihQdVnwVhK7axAHnOGwAzqVaaL76g
tEsJhrVYDuaj2fiwtP1SGtGcPrfTekEnOV8EsodM/ahK2QkRPHn/JqMVWAh1tKDw
e0CK5GPJACCD8anB4gt49ox64D8ehbpwPJmwI3IVXCvMA5JDOcSWj7ISpAtaYQp7
mB9l2OA1hJeSd00ONvwwTyfYu7rfIPnHaJDEYqp7YJ8E/cZVaFleSrnL0uK/3+6+
l0TCYUdVht5zZAnzyywe1lTvIyC/cKMrYmgueq3ayJUVbituDUq2iywiccSk8hs4
IDVu5oyKIR45Yjx1Y5UEQFdTX5AB2rJwrkqBagINt8Jqg6CXx+cSJzjoV/GCNC24
9ZNXCbqdme9Eyi60M5h1s4U1lU1tcYI5tn9Inw/++5ooBrnWx4AZgX+eS+vDEWsV
Pe2VbxZorY63k32OPEkjuCsoPl0bNFirko/j0gO2BrhM7ZVcdEP0MphEAbwsE4Qz
2v9Y2rVyU8COj7ZeC04xF2z5Chadva6KeBHB/lyGI5h+k8IPp3XXQOmomOZXoUs4
MpGGO3XMBKaVK0NYJptz6jtNaRTUquR022WQFUBd/881VFwVsCik1UP194e6ye0P
YXOdqiA/pf/q7Mta/EyIPhJB5/cF8mP/6DZ1vL0vNsYZPnhNQaEOZQlbEI4aPK7K
Q8p57I6yzd657YUzQrL9ZcSRvN2TOyX3659zyl7n1faWw1hQqei76fI65kVjzCE8
Xc7YxLpeUuzxK5yRlUtUMm+PsW3L1NPyfUQzb2XZjG/D3ROgPpHEXfGn/aHKVM15
YOQcTb5kObmCYW1SlBt5SYL/SGHiDf2+3dmG+V7xhFN4IPD0TMyvjbsNQJ/Q5aQ9
npiBtT5u1kJDU5CCSVvZLJmMaiXOYhxR4I75/OeAkhm3CSQsSo/GBCuzS8ZFmLZv
+cupvMoEgVbrWkOFJD3xQ3BCNY0G3TrtgIvZ8te/fkl7a4j4iSETic01B/Q4eygC
uHpRy38o5s4O+tii1xx4ppWrqxq11TiPmEDCFznhiA5PpLqxuPWQHyxtRCQc1NJs
FtwTJ5K6jE4N5GB9Cnoft+Es08cZTSnOhwo7PhBQO4tQf9ZTLhZ3SzxFD/dWjSEt
gRMiElwbYrEOk/R7NWMp3C0R1ef96KkFiK//JBuvemSqeLsJafdCALz6eemxWNCb
iFfNPYm7KS1G0gqf/zGafFhQHL2bKzicgkSnmI1WzVJtFgvUJ9TOXAuDDFpq4982
YaTIuqi0KWGLg0N6cXcMNezZJEMydu58lVQcopjNrugTMeR6BZaVZIKosSU452XO
xOpqO6Ez/uXfCS8jGaHdiX1OtpOhhoMwpL1BA9CenerYxsnsj1qHDYaEBl1LWQnq
TT74DBBh+ZUXKFCehbTjSX/nOT3BnnVZi4q+AD9ygdkPWSGCUqq1er0qrWP8Bw4z
siJ1OLRxKQOM1DZ7JHyKw5tjM7ZrmsoR2nNkNEbVj+EabYgy6Q9dtqGzOVLBbHzW
dZbza5Q1TsGgm25iiiBs2H1onztYVwXIVvuC9t13pULZtrkFcVwhWRmgDfAMONY4
RPhlm97SRaUQVI4qlshzYkR/jDWKxcZAnSa0TMpC8TcEg3JsP6YXxCbwYXGYWx58
QW/1Eq8JRmM4unYyYqzZEfgIafBuMu2jHrW7X+tkpNHaOGyRN/folDYmFjgOBlyR
DfXNPa4114HWiOVx7LImSjrApz362xITQP/xPt9anVOSLWKX6G0Y1jKg+DCX/cvj
9VnS1LNpArXiSIMetMFll/otF97HBT943Jyv+EN1gs4Gq/yafD6K6+gySTRiwKQ5
2pjrlxXxM4ePGPacsPrDOtnJ88fu/LLn+HI9xnZutLzLe1rRK75tP0zmEDnUotNk
Kbdy+nGpADW/wG2HiaRigNLaUZg9kwKsaTKREr3M0g/QXukOcXi6adVbu4N63nO5
Q2U/nh21Pxq8piGUjfR9WmDZWAltZBz2/fpEQmyyu7lHDH8QGMRYePPoANBiL1gZ
RUVaNNRe3FWdLy9cW+9mkHmVxLDUxcUTsSYAs4hy3YIxnxgbIE3YyePelogkU6oI
B6DhppWBCKyBjdaHguUsp5vKXB7OKOWtOQJpr09dNTnR5eRSP4Dtfno42r5J0W58
LnFtQJHESP5fE8fnYX1g+wBSFnpAN7ack1ekhHAiZUroYdS+fjPzvqoc5PGFjDy9
I80BWMal4N/IBOAmI14BeobTBbsk/Mz8+lqm+6KiVe5KXBvQnGSvE03VOjyeYIZN
AHxJtnE706+HGmoGL3VAOstKK+c4VPupZy4Cz+7VtPFDXORoJy9ZkltCCqVhD5M/
NZb+9BigND8xvH0Z+EGWTv3gP96YFjkuqi2zxj2wW31Pgd9od4kCbTr1s0wGnhQE
w68H9OdDBp7TjZBguIw6HHZ7bf1WnMmm+HmgxMHR8llHoO2zq6CvF0hjPQ4Qi3Uv
8c97VLtc2hIQn0lh1uadGXv+W103IUjxUMgg6Qtl66LfTj2WrvZNCu1aRISzKNmZ
c2GNU+JlzOmTHrs9LWgTYl0wf9Uhe8QjB6T4LwEMhsdWwY5+Bzr+9EcjzUK6nDkJ
uNuwlmcSWUjJgj6dZk0aiiP0faBjLsl3DOBByYRzhdxVRD3la0pELTT/3nGsOVcj
b9C6dW6lf1yexvMIq88fKsTuArPUwABnEm9h/Yb90Sr4prASkXdTGu6up6ntEuOL
9RAyiitkH46QNotj2lW/f4xYNG+G9s6/bvG00UbCbws9M+xHsSR2VWA/c1550nUv
PKJE5HLV4Gpu8NQ24auD0zDG8SkbczpvagK+tMiGiBwz1mLnY9JVBdGCeKhQqbFG
bH5vljCz1Gr5EkHM/idfAhUslWxLsgTQxVLffWsLBwmv3gEYYTCyd3iSuv2IWDuC
arh3cJmALilLTKpFLE0YsXzGaFdTQgqfWNJVImu9TpP3nc1oZ552b99klRwuyXcq
SMW1XKgFoVe1DCAuQINa0it5VZLvTUca33tm3cWCBHOZuaL9Y3YYvHfgpTAcWsfW
Z5lTT8IcPdbcWCu8N9/b8zXcuwH8PwcInhxdaE23eB5cTqF8cg+m+TwNRAgmEL6b
00dq/UzQaGYZL/7zQ3+l7o+Lu0F3pjlcB3n3YDwudXs569LX0u3aSEGoLxK9UxKD
TywDRcXgdNfebn6yqAL0SZps4QC93tYD2mWF/R5sOJnzX6GlYKpfH3sua3Z9o68y
GHFN4wpnBJJwGGrtAXhg4hFn3AwBWoxioo5Tao5O65/Lwe7tXyF/pgRXD5eyJDm4
MJNO8utAoXCKxJdg9nR6mznVzLHBBPlwMZP6vLz2laHy1taOcfd5v3t2RnWcr9t7
tVouontI+c0XA0bVX4l5edX65OJxUVFuPiF4vbKbZ2IIGlukRkQljxlHhzcgrIzn
iUtyc5NEzsZbu4/mbANyBAhZbnJ2ukjiOtK6n2+1UyyLQY6myTrkopYEvo4xllIf
uPOq5vIuyKl12q34dJJ+oITKAsK3oQRI70ae2lYyq6ceS9eMStEgj5IUGhXJx1lh
qohtLBzSSfCeZjYy0TvN9GY4wHCGFHQ8nH921evdK+vwn0NxbbaWFsGIc1Mvrzen
KbFAO2vp69pR2x34s0toTAFenq9DGXSgkYUTqpQaqh3gr/7/0qHX3ORtxZc9OnhO
JS1pxlbHPQaAMD3DopU4TOe9n6ZhvdBKvVIrq0wavXqWO0/arGai84K3ZC/UI6re
SmZH+gKmFxajW3Nz/OD5rTsU83VWsbd4zbMcDsa7j++QJo/bclnTHblDTJdC8rI+
DsStzfc0QKPRabqy0Lt1l087mzqdQr7ZGFhhau6D1VMCv18Fjt4ActZS8JQsuDx8
rUiPqnQKSMw3zXLUAiiQPo5EEYg1Z3EsSiqna/Pjz9Y8JwMw7VGmYhgTzDNjDohe
zSHuObFf6vnQ/GzekI6vq+kjha+i8R2m+mQc0bfZ3xMXuoNwVbkVTAmyZe+0kJlm
qSb+MP/YmZM1TmF5m3LmQEXbeBhCbrTv3U1rmYFugew8qEqZ+gUBPaTxKV5Zp26C
25YRVOBgxl7HM3NDyv+Y+V/v/CTJUDFIefFPLtkvfBFvTMR1bbqjovuNypn0LqsP
6RylsKPmUiscg0qF3FVVCD+r5IwFReAyJZuIevNok0M7hSRbF8uQswi8MYvsaJSZ
CgDW9IKnFkj1lly94efoAJqJaDuBnl6YtsHlg7nnYnjWvG46J/oYMGQc4rxdQmuh
FiUI7IEyU4XVYLSlAa0/wZ3cRczjMH1NXRxXg6Oxy7IpOQeoG7wl5ghX5XZjQ3SC
X9yzdPIb8K3pINz1efcdRFEV5/BgaF84AXbz2P7CiJh6062uFD/7AiHHKk/CYZPe
0hH4OT3/v4ZU6uFaIBf8XhO+JcpYzd1XuiwJpp5SjkX7jpLBRdrPs++doPuqOChl
ZAuxi4V83+sTyTkB40Kp+zoCnMKEOROArvr3hJB0LIEwX/ZBOtNhD7fQcJfBNn2Y
DhSXUnOMH0ruycNbJZN+kdqqqI0KHkFsPUSyeaDdZq8VPqj0bXJSNKWE2NQACT71
J8MGb2IW86CnTEsd7Y/LHtijpR117UhrTqOINs88Towe+x6IVaJU91HZhMv8bmRp
9c4caHK2TDB9rcE1FHoGtmK2TUD3PyHMf4SqqOVak7B8FZs+ofDOQcy9jRvQztIe
bHw3lQVI5V+pDcAUEpv/VYp4GfZ+o0G/x1JyJPR1InXPzbIw6kQ9KzdBIxmWLTGa
zdcKNGPteT9hvLQIi42kr8hbZh6bEc8de/f3EXdVE2pZ4ULV40+GrVUGExGZrDEN
HUd0D7DzAEsUEjV3SNopN9mD6pbVHZFAH58Ab21HNP9TuJMafsgz1EmIWjsZ3D9/
eCJKC8BR8xdbXc7RH+diJEOsuFx3zc40zAW15Wu458/tq9xmDQPj3UgaDfAeluHc
swhPvcmy3gKGyxdxbBbHK4r/arF4vsUQsFz33D++zBboyPUBTrhtCksj66Qp2Lym
vsbiGeNIEshnSFQ+iAbSHojwwBM+4xOgPgHMorOMsIarhqksluX7MXw/aFzXChMA
C+NmpYTWIobfauOgwvCKQWiobRVYdFmVqy4UyboF+dZfIINsaN9lEedp+SxXsAIJ
LgsbL8Z5ueSxJMJaRNkgoNA6HE+RMe8E+99PKWqPKcRBg4oT1Bt0+d1cxT20ZzU6
ohX6MWgOu8jqkGC6Htw4kKtmmvQSTsQK/IjcDRz2QWw9/MTF3Oe+Cy+mn+aHaLm0
lZTCPkGltwKzRq6ZJ2m+vOEj/PjiCfIMfCZA9qymReuYetb7CJtS89wS2ILAXJ7s
kPiQEljywgX71ej+ic8nyx+z1fg0qBS3iU8mxDnsxHFcGvngKLYiD6lynR3jGe7L
9JzhzYAjCt1JikE/uMDOF/lylb5H9QIVzWYuus++l8qHWP8F1/qHM7YQV/Q5fPcV
XZnjJ1DbZWIj2g7Qj6ZuYETIKnJmzoKVwV8kkADF9wOVugEKbXYkaKYp1qAwrK/u
P8ArYUs4rhyYeuIFQK9UFJRFpPBpG0K0Jm+u+O/pXHYQ6f99Tmigib/aTdqiUukM
NuQigc4CjS1oRxPHsP+QrDcFvIfKfwaCXf4VgstzsqwSwuipywVleoMQNnbwbrkf
wuWL95sV5CrG/Dd59d6k4dnyjvNXnKM9qYMcYkfbZFIgAUr7GEuUjTIknipJTdNM
Q9uC03Bji1VFsoXv7DTTlg+vgMq05IqAPXN72SVJhQhOHMW70VZqGO865Bi2AWTu
8iUjReORDFOHntjvsIm7YhZoFPDScB16VWlZ1C+8m+T80R4QceJ23d3Q7rQ7ivaR
0n0zxyFSQYH21e2gANzXrz3+sr/qKUi/r2cHN8axhr5glaeQeK/ZliIbYNGnS0YN
PQOzxITgB5pLJ2Y/P08oZEFCN7TJH/J0/bRq+K9NkYvTq5obVIIcIMHwzCV21fbj
nIZNopDMxGkr9KUB5gnp4HgikVM/AwaSy1npNMg4OfefulcL9G7G5A8RudJkLi+g
HreuGM2Y/l5MERJc+9+m4M7gC1172p48JLMtXBaS3FI0hv5mYaxWKvhCjGXw5+IN
G4uRjAZAjrN5RBzLQIOkFeRE1pjEqxUenI5XWSx9eGOI81FjeX93n1ZOcy1REEHE
2XdFyyrQ7XAyXErUP+rNspYBJkEaLl64pdk0rP2dUG0o914zbLCaAf23eErFsusm
JRrrlTUTGZX94TLoRyBzU9Bn7KxJWSSC/FhL6gDXytxsOyBcOpvpuw0mwswA53gc
gjcjCC31EBJfCKvBJQBje1eVDyRBhk41fWAFGJIPaHq7iYmGT/o//0gtiFDAklvU
mm3bAmd4UpoQGJ6JxrKzbKHF3Q1Mb20tFN68y3Zmjzqm7nHSxOYVcWkBeRRlyM5G
g8V9LN//0LzCM//LRhaDpnLGRPjgkzM5DFazmiuDEf5+SLA1QAiXSk+I1tAUhiFL
RmtjLJk4SosgyFdVDeUoqNKYfLg+N7VgtISDAw1Le/B0b2Y7+BQ9lBN8Tw0E0G8s
XvCLaSFItGZ4l899OEoY0aBCpwy7K/ZNw+vDfohCODuMio+OJfF3mvpMEAGIvWAj
vET/oKIeshihURcBABtxxwuLDXCcSLiD73LbexH/IW2Gi4WjKg29k4aQiag741jO
Pzq9hxCn8qlhaoaRRzdjjCGmYoc6d3JPQKJH0pwySu7kzAKLOkgaRRoH6BWd3eaG
C7OzevtloU9P0Mc3nXd8k4FheM8xY6ZiLLqS/T5fpbyfBdbRJSW5UrRcyQuKsYMN
ItxN+VGe6t+Zj94z2SvRaqoStYoaPsfsh/ieiR4t/I7uAArxRov/dmdt2e/tP6jf
kauQEcb0D0/ygWKdqA+ez1vK8JSc/UacrBp6fxydPoNCrsWvtWPXeD7EjNGuMQ99
w9lo2MKuHp9AAFh3v4wbhQPVLq70XrIm2EQYCV/ZPNHeTSaaAvBXa2PTkpQ99G+p
iNv1oV0b01p82tnJzkiwj3+ehiY8TrxapAWiWIVddzToxE3oGoM8WSv1QNZjyZt6
/1cAgJihXcSgZqXeQi+C0X2piimujG1wPYSXw5UYGnTkO/PjxYPmil0d8hivLT+u
59uy/TaKueQIUKO/hBeT1WxZod1iRXvb916qOEDMzauxmxdWT+BJ9QLjdsvkMejr
vFIowlpGMAYNZqMW4UvGxO35FLZQdmRdAHnySpL5UMxkx6OYjd7Yauiuwf6ErbVr
g41QF0Tc6F8B9+CzHbKcMDyd045yJierYWD9A0D3rjVY20/oMJ9kGVqAYkLD4b4k
apxQD+BmJQg4uWKlTC1JD4rvihcTFNh9O/hlEw+TUD8rW/Suli7mICFIk2K0n6b3
aznh8WiY1g3Qy5uYd4udrk1HpSV5JQ0VNUiuQnqbb54/XH4gAOfacsPvhZnofRa5
bsOZ4fnlgo3IbnRAfP9n2oNrcV8fVwAxZML6xHNzhSCMA1a8R69fYO+fHNTqFMzn
ru2DAP2bH6Lu6/tKuzyJMAFO/w1KIB+HOjg4FA4AzSkmeAofxx5og+uFJ7G+SnIM
MqpwZwFmxFxxFIJskgFsAANH9drzjqX6LSaTCyNS7W59qoRD6t8uIP+OVMU9tRFS
FXb9X+I4QtNa95HSbwP/0Bg3wf+Y/71G/VFBBwo1sEGuSNnKU2wao6fZLiZA+bo7
zhMZPejcN99R0OsegnmfYn/66SicCWj+db6ANhOH0039ECQpIeCME2TuQtn+ocAD
kpNrwW+cP/Ie9fOuNKj8zKw5yZ7xeGbfBgMS1Iz4EqLDJAysJfAtLW5bkS/+sij2
gSEn80DbUSu2nWBMsk/TtYUlPWkRRMXZH5r5bIQaHGEcPI++ii21mm29CUrqaiMo
6sJyQqTxqyDi5sW7Y1ojVW5H4jbSlPPzSmbVy8+yp82nJYmhW5Z4PUQk1phshUoL
Vl6v6zyeQVx3UmTk+qE11epjS8/TMMu806l1vIWqyxrQVXFiMZyZfb48mZgVymPw
kLsPMtdmPs0h4UiBWUyaGhwifYViVMzHxFObz7ubE2MtT1/Qlir90CuoB8ExKr1L
08WOLy9RSQP9a/CldbJ0SquWzmDzfMC01sjlzrmV9lpgweCV51LSR7PPO+tMMimD
fiwR9YX6P9TAjh8JE9NbA9Fzpr++IPdnONN5QxzqdRT1oWT0pnradoAbTKKK35YT
wL2uFGnS28tLPPa6y4wyzty8/MrOwHwusMhlGxELmoQa6mWyOcPruJ64AbjtbKIE
pxJELSDacf5g/6RHYQZx87U85bLJ8Mt5wSsivXly9zIGjHLbybgOLb9g3THAZMh0
a2UnyPHes6KjjES+85F9bFHse74FTDojEAMt5UjxisCFA7V96bKuuo8a7zek3Hq+
A6XFSG4TPzNT5xaCAY22yuCPDjF/lWrFmE5fVW2gGGLqrTC+qSQFr/6xDBtAgGA6
83VIojb83oPGPdDHetx6Ikow25sYQL6d5bSS216H00/eTzIehCT/1jvV4CRJPXGS
t72E0AgjDalIx7wnU5scXoiYHh4FkvEs/JXsnaWG9VdOwZfs/kcx3I7NwpVQHgWW
Qih7apZfkfb359lQA1ZABz/75nlqlWjcpzZb/c40TveFk315L5vwsWeNo5O+Gt2M
R3dfR1wDKBVgMp8MVHnECT5hjcVB3zgaCrcvM5jayS3fsY+++rojPGEnGBD+le+a
aHcVp28fN4ANPYUWZnZMa6CrRYKR3Zpsteb0ZD8dJPs6CTKJ/By/HYpYkFjgNzDO
o6iwKYDagMcGV8oeq7XMXwWYqrqIo86KYMELTfXtNOVjNOiAnFQ4xOdbcLmAiKbS
3uVbA6VW3obcencOGGFFTjy7O7f29LGfKNNjqIOlsgoyTUrhia7k9t9aK/gA+sSJ
PoyIHCqt6FGZbPJ5Z5JrLuPmuGKcsUduZrUMjXdsOwtC+2l194yyt/V7TeMxIcPR
MELKbb7POyAQK+QLf9Y5wFl4hxdUFrDJ0PKYvmiGMJOQS3J7304FFb7Daphq3x5v
pZdQ93eYBtXHwBInBsOFG8E5/6n4qCAFMVXwquX8XjG3CBHwTTL6PIU5gxYOiSlK
gHMT5g0dlqnkubeJKoXUD+VBnlV08L2m9YfKGK9+8txUgtbEvbTnxS1Y5BIIORKp
OrwoR7P+4iK1/fPu8N40tF+ucXwpLIZaQ9Lepplop0axFLsIl1E9yjb148tCsDfP
jb4A3ObMSc0YIGT7H5Vy3EdHisOLqA9Dxb5C+loyTQbMkC+2Haf7mt7Orii9m36g
tWFC5POlrNgYgnykK366LGXJyqOuVNvvCgRmRGNtuOJiZujkN34ZqTxYqjFw7o0W
y9E11wo8LHJEs6sBK9irGLFjB+kstHtCHMHUWrdU5fdC6hZ7DPd654khL3SwTA2B
piMQkk/T7rbOdni7wU4hmTjA4QS6YJH3IM0P7lkoyl4qqx5JjGgVVhR/GXNHsgsB
XbAy3ihSqTH5X6K69RMGuTZ647U4oSVRoYcuFqTIKTFEjTNSPCrzUSF9yo2BnobK
oiKq0y6Nx+QPZyUf0nEuwZVlzAK+4sZglqy79GDz10jiaq6/erYBBqMf7m9yI9IQ
qtuXD9/hRTkPPlnEvhXduNBBUWO24p38EMepHJ+1OTRn1v5N1Tsfv4eckHTiZNe5
3bHXWYN0Z4Ld9VMvKGQ6gOc/R1wS6QYnuDSqcv7mU5GplwDuL7IrdTWK77RI4YoW
7Z/IBnEXpgZLJYT5FlHLxn4SwaqwbC22Hqvc6TmRS+m9NoKdso3+JUHutmaw1iXs
TcPzurQ0Wiz2LHFsA1a6GGZZaJazCE4n7D36onoY54SMY56hbuLPLvgRWLmqv/ul
J8w2gaeMfFobBSGoj6e5ywx2nY5RG5vVYDGLvxiLYt1iYD8UPQoLvag2Y5bByV68
5YyJF2TxH1GqHj/s23FQMjPDTbnN6WIfYWt+WuEw7xnQH8WBsqkELGhRWbEPWw6F
aSr1Boqw4x6CLuuZEk8H0tmdtcHsuMxtQwGEVq8IusNpH1I85MIBl4uHF3IkaeLl
Qn/5QqpbJQfmwYKW16nbeOLAzKs1dXb2+/ZR4QIXmAtOH9UoYpURTiEAuSBTCShy
cK3TYrxejLACRNdc624zLqOW9KCJCjvxy+uFA0GrhRcXCzkKIG6R9j+xFHLxhh+S
2VOyXlk4CBW73X3/hF6406q91AOXarKcfztrWkXaJxJyPTtFr8TdAv+ZiRh4LQGm
+FIXqmjSggXFMXV7ru/XuXmbQuRqe+iZp7dpDuy5PayJq4WvUA/XEb5Ksp2/LgGW
uTHcMqI0XAGgqAfIBwQ7H4+2rvVwbnJi1/YKmVQJEfLr9Cj+veX3CmGvnPLqC9OY
ZXQrUadnB3qqKPb78GHn4NEcpbPjFy6lOMnhaoXNU5Z3FR874DCNGSVoiTA7lZ4D
F23mIEJija1wEGMc9NVdqSZLgDMY6RuOBlwtc7BNsJ4BUdc0XWx+Y5+D0aH4nXxa
QPBDExLHIup7Qc+ZlyQCHwKNTWuY73Sritr6bxjXKgvbfjNvsdu+Ly3STbA1u4C8
akiUphhu21z9v/Xt8PRrgFIJiVMnuQByW95EC87wnfP0kMwgOOv3PqRxsmwOsWh1
882Zc91vt/ieUCEYJDAHXnblKaJ9Fat9zMcONymj2tOektfW9hLFrR8iP42DQXHl
GMv3R2dxC4yv1EKv8z+M6n4fRlyM5YZYJRkyBO3gCFR8Lrb/xXN/E2OFo0q7CWvd
hZdwxSmYBQ6PHTFS/5PZF8n8UEP9pGXFr7ncrSbX8RbNGTqCHcVL3/jCyMgJkOx5
isz+19cIdj3hYARX5N2Ia5qjMeOHFBcgpBLm9LWvpR/Le4spYSki1ws1l/pykJWZ
5ZhH534kZON8S47bVR2noD+Ak7IKwEbXFDn48n6WKPAboPwNy9u7HiHujRbp3UuD
XdsFOGMd4na9IB+mz+C5+DH/Q8yfMswXxxTW18SS2snbcnmioZtVcROv674Wm9fh
iFsFd7LRpBVTUJ3+71layOnKNoz/YjYP0LnqVgv4bGnmWqS5MBc5GVznvkELcQ76
B8OC9lup1AeApnxbGqITmik43P7z8Fq32yHL5rVHJg8/9TC7AZs+c8vQHh5eLXnT
XvWc0TlisrUKy+TCuq/uOBPlCLMwIRPRQwFN8wm/H962Xksc/2N67GOEW0pMB1tV
fTW+AY3/y3Kc3veXuxqBTajYsXRFn+OHSmlpOv1ojcC1Uq3JmCjzFjyqQnXl83f4
`protect END_PROTECTED