-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
b9qph1jivF+teMctjM1zTDsmdyDcgzxI1V+o9Rs4+dL0AZFduwop57wJBpfOcXhH
foMGVznBSRvaUEwOmcUuJHiBCOGEWSb5CATtIiIJYKWQddP24kJYQcWqJ9w6g2+I
Uxxo/GcJAEy4+XVx5SEw/BzSxaHdGIt3JqVD26bJfew=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 12517)

`protect DATA_BLOCK
+8iyNBPuiuAmFWHKkUXm7kyJ1Sa1mHDLgbkPJQZxnmPd/2sOFcmUPwyn2sfUCMhn
DYP0m8NzyfP7VhouZwfHO7aWYSP0+EtkoxgnlnNtb+Ds1Sk6XRiEXV7w66m2AnhN
Ii5UGKB/jaFMOHVe2vc2U3GmNtN7cem4ArHiejTyjaAgA9w+3kYECVaEkBSOWrWI
8ThNBHoe4TtdmEPvSl6qtNuImfncyXTFIvVw/9L4J9HFjZSm17hX4IJr1vELOtKT
wEHmMdWzPKsr1ZxL8aex6fz8GuXm3ruRuXjbYzTaQ6FBPr3XXwBA2bkRP86+lMH+
yR23IPaTf57bR6D3+GiVpllA85lbKEzYGaRA/Rrj1DGkCoWqOjk+swNo194nczXo
nMauD5KQ55/BB++6w6bAkCdTMCqWRwc3WVvDnsyZ8aa5oPdoAy7oz0Tj31aF+3K8
4A0bcrt/7q8Zuk8ZLAF6N2/zU/pbicvuUm99ygV7Xa3ysXDXvwMITC6CR5bTfWRq
X997nYv+F8odhpICXVyAEFOE2b/iTqKUYsw5ZMT2RVn8v3Ht1XYwoEfL7DrZ/7fL
VORkLYq4JLVYDJl+qX3584oq8lXObjO4GtQn1IvYnTQTOwpgrD+XNF/tbQLDABt6
WJzMSQqot442TPVWQ5z9uPs1gXdYdFUP6qbntvg3fjy5nnkqKqVycYHCiTq4jT9F
FBo5qU1U4Zl7wgD2TNbZlhThltfoWJ0ieGuKrdXR0+GGUpyT+N4aMKkOmaXC4FpX
/EaVpHF7DCS3IhRdfrG7cJkUQy51HMy7Jy/TnZMmLfd0nyiZ/7o/vMW/wr0+ZWAQ
HI1kW7BHPQ7xRu+yasx6c80Vigi4JVzgAQvm/zx864o2qnAqPXac0SiwmiQBN4dZ
fsjAQXjNuzJDJvVTbgc6RtgGUE7i6L2V6Y4YcgjlhDB06X6BkTH7LejAJ6aK9czo
7FS/Pj3gSPQZlXMGJdIZda+MyDeT5dPmY7YpiHeuIvUHRsRFsJyMWCc9P4zuOwZC
rohSIxr/pLxRc+/xQIdmNF9py9PTGmzpqTBXnyRMl91rqQEwnAXoqsdCsVBv5A0n
75WDGWj8w9dRzsCNxGv4WqTNyu1JyWHyqCB9uruyrNHJ/hJw4ABl6FLze19oDFgN
ZXRFwUNSaLbV7cgcYgnC5mrlxIOBDDvlUy1SoggFISOaCUSUgZyUUiJYeBHXdyut
anyw8owTww6RV/YrBnbVB7VUt8GRk6P/KW1CmwbOZ9vF7ZZNdOmDsuQLJ0vivFaP
ZHF6htuqjblwrDwew/G0t4fL4LrzLTIS4XefWGB3F3vjDkc/2Cva+nNyYAOjMvNb
/xW1VvOXpnzgzuHhWK7fSZyORI/oomTphldsq2NgXhzkJrFNOgD4Yczb4ejLSdzt
IISBthU9bU7MY7Eng+EIKDUbQSHEQtlUuE3pmt3Nh2KGcwSYbY1kIl7RxTyOx8/V
ggg+ZxxLV81j6KuGR0elptIhC7KTUF98KB6UQc2vAe74p3/5dt2gOGEc/65ryi+F
5n+bDS2LNXgN08LraoxsFTf43xA0VXHrmxaNI8NLyC7aVJ4LXUmBLLR3WJIzje64
sAna348HFQ1erOk+Ae+co4CG59Ug5c5uRQXgzJO1Z2IQmh0ITEjNQnPIiHif/71m
eUUlmzwenZYhhGxOPX50jH6l4iCCxd7lQpLMpNf0nlTB6QN24hY5fJCd/28HNx/J
L2FRYuP/NBYwAlCaS/4oP6Cg4GR5uymjxRFo4OLtQSnbOLChgks55U+TD5R7wDXe
5fXqnNQIzcXid7V4ZlD6WnsdkfrrhJh03mUYH5s3gay0aY9jOG4gTxHtbop0kUnU
9l2Ml2WiQl2ZNtUQFADq4mMfivK/GrRC1jJRGR0q0rdvnFCp8GmMSb5V5JSkIAUv
l7IR6vbGWQvzYattkYTTPnMqtfTKCMvnr/aTb03BgxSWKDJ3mFAhWafb4OS9cbXh
0psOCVN8FARf+VQRsEbKezTGymY6fJtoh3uM8/MbZAY2sExtrvV1CqxPNxi7khSA
6MLoNnSR+Wr6pq0HqH6heno8vmUnHFIYdOSsaed/lHmTrWtSNaMXq38+8ouf7y2w
6R/opFTLagzO4uUAm8n0gxNv17fmg+reSh/zgOEklDe/y04M0W/QfcyhzLN2n9aD
AqPf08VzhiyQmEn1dDUIAu8KyHZCJhHEXLpi4ZbEcNm7i6KGhUOeUon1959gsMrX
wvIioPPCTaaVhhRkzmuzwbgr1GlMedNCb/utnPt26LPZ4RUU1JtlI8fnRsysiSHL
2ePxm3UOBogSpvU61C+d9SE4+cOhlvWFd1KnUL9a/TpwwCQMJt8m5FZwF6wTwVpL
jeO+uU3PWgaUjBkC/7dqEXoKXR2EPdsQ2sQUSPN/cuIONJCjDn8t0wUwO9nJ4amA
Zl9TXkc1mAxte+rp1NFauYKhBFfY3U2L7ESx7ycNRQGFjISictTab9tdey5ctuTq
bW2rykeVA15HCHwzRj+/rMOUDtmutUJIbqFDFU2Gi/M0Oe4hNZ8xxihTjdZdWGAX
zZOAUme31RVfzMhBTWnQgPa48j6sLTc4H6BTAADzuBpEiu8hT9L0A0w1FpDy2Cmc
X+Nok3vYrduQ7m1oqymugB8UUuAWaQFrUV+VoTVFaTUj+yqF1TPtZQf+UC3d1Z1k
pmxFr+zBr8l/EfoqXkzGCS9WMQXv9kSI0Bbf/Ig4JmTXD8PKMDkvUEEC9NY5SnB9
cp4IT8IuElpNTPUginV3G9SnFr7gp2jBxp0vwoJQXovs7qEbGBsLDbS3x1b/0Q5t
r8SPMLqkRhvhnT2dwYe5bME/jsGkpCyaaAVGJgbfCYoKgbt5kcvrM4H0OfuYwGYn
oxEBV/2T5keS3QPa8WV8pkWI5+dWPkBQh3Rs/CDYOsjYO0RrEOQVs7KhzMxSqBqR
3/lF+7O9YB5s+qpC3FCe+Db3RpM0cqJOfkfeCXUSKKo9lSrdiCCIPznGxn7MzAWi
eOJui8q+/jeh4FceBLHnA02M5umAQP5cYDErdFoPDbVDQxQX9Lv3KnVjbwulo+jC
e8CKfnxaMY/MK93ARdpxxBCi/joAdILrCCpUIDWFh2cooZ85ZD7jyzjYXuKdGTFh
91GN8Jl0F5ovD84/pq9SS8A0AbtZfJyWX4BDwBo6uN26YrpR8cs+BxvSaR53ebmz
B8p6K0QlqkKQr65OK6/XkPQB+gJhdmOr0rhYFSOeXcaGwdxWTuQK2/BPPqQkugxu
vlnZQP63h3y7P6+6/HVdlOhI9XFq1JkcHNleHVvPHLMoGrXfVBnpFd1ltJjQuHLK
4ml06Ep07QJrW1we9E2413+5Cjx9IC/8hnRGXkL6rDvyJ7/f0dJsx77li/HH5J6T
isokCO/cKSJA9Y7HhfnS64OeP2CSsEAhUNUZqfpIYmUIHsr0x27GSPmaFdiIPryW
VRrBme9lb7kIehcgiSKqWfjr7MuEPi7QS+LSlLi4Y3q8xbldNliJ9TE1oOW8CdfW
PwgFsvAmU24Q0H/pOfbWyEWfkYjrjeZFk/GtyhVUg8nsSGXWuLBDT1IXV1h8MqDX
4uIiOZV9OC8gj2cyCH5GqRtXrGys7kmh6Z3GU5V2hHlvqLxotBfIfRRYwbizRAb3
6uyGoAK2NVJ8rFAii72Ccsme82XkihptVo+mILMDKNPrWnl/DRKOp7aJ7MtMgKhK
n7rx4jIofzJj47HvafgbMi2avvvMkygJjRCHEnO9mXAea9KsVc07mSUfFtBEZ1Bl
PYT7sX8ALj8t/sRicom0nPvDZxqcg0XpZXt+hftwJhZaE6yTJvckF2vyokqF8hY2
xDzbKE4fXCrxx2XIazLB5f/Udw7vm/PKodrY0rCLa4Drh4h4e7cKTziaUzdyXiFk
8UFb6ut6t1vsODR9PrtWPZS/1imBynF05i0VAuILMMEkg3lY77LFNEktmAidfe6A
zNDG1Rydvjw9D/NYoFISx0gFehvIE0HnnSrPGVKF7rxag859cRsw91EZVyGNAzGR
Tec2gG6H3INraMcavCUs4j0vw0tsBPVyPOwwZ1wEiBYIfI4i63ZgnhK8gql3CPim
+zjvMiLR8cjvTFuXcJcg8nlUVCyS//zp3ZDStIj8SEo6vUgDLQVW+cG3bZ7QZK/G
Rn56BtmuZpExB2qt4whYQGZE9wtvjQCJ9NuQhlcFyzhh76y8tQ/FBo1h+ry5zJmx
DcNqTM0L9k2+93FJe5f9qz3To6tMRo5lZ6n83SaeOfX81yjKC+tXsMflx1UsTuc3
W4sJweGQMnGOfcJ6JkuVz52/dM8hlgYRyHQnLgHt3CS9PO8HK2W0xd24zSFinh8L
5astEV5JAN49M4PJfRVw+3QN/md5eGtGHb1grFecUS4WYtafEIzXfgWDjDTHIX1+
c6EsSSoIlGD8cROpdok+7Q8wQ77tfolCxl9YtGQqRqRRPI6gKXO2fLY2z8wuSaA+
U95NLddnqdJykDuubRZOv1VhGRovWdfFTBKf5FqIhN3Fkum3t29J+FbgsRCLjEnC
1guCklplhvf2JPQ5KqSbIS28rzV2sc5tQJ4UWjd25dog8Yi6b2WPPK3zLhIaDiiC
k/vm7cz3FGIjk7ORh2gpmJ2ttxYJHJzb4VKcKwQ/bl/8ecUS3LG5UcGkf5c8kuXi
Y1AQ3CyoymiURnoak75Wwqqxk2y9Vr/G592P+0ZF29MRrQ0Lfq07gAH8IOTqaXMM
uY3Hhq9FLv0lRXDXH9n0qrEr9hKvz8m+kTHhwfHVgXBX5zvMO66OF7cPta5sb3g6
10WQQ2a1RcegJt666dYEbyuIlwPpX67v7+3HxFaGoy9lF0OEszbKXj2kVlg04JvO
9oNjaqm0J4Boxf9AJdS5CjV7+ZXRgCCZJ6zNTtr9t8ryiXkyhZOKEa3qCnOVwm0Z
EgER/THqh5jmOLSeeQaGiYU1nJjXaJCC/4+stSc1jbGZK9z6C4EUWyNIm4qV8Tou
YxMa904BGJKyRjfTgdBfXm50jScss4nVHMG71Uc+Lzo3o1gumTz5AMGEsG5nGNo+
k6yghDkL6ezgi/IqEBVWSCGp46EwslS9lFjC6Pewdr8CrUBrZ2Yc0FWGxOMzLlxZ
zEoJgn3DCMecEQKN1P1JMQ94STwcs8KCPNSI4y7cpKoDcDfpfDs8YYQ2sCdz/o0g
YgCB1tbvyr8NVS3zKrU/tAKs+CADUOvpzGnFWDukKHOwmZa/JK3Fa6mSTuSFdECb
iVgPw+aKzpauL69EBNoqrGYZZr6g4fZv67hcWQCg1HIThBwcCU9fWdQH7ouvEQf4
1hWuFcVMUGkxYg+8lGz9/t0sPV3Zwknj8k3MXHvw2pkxSfA82ozVrlifykKEpNPP
M4GbcPEHFr+qSf8+mPNczlhU8wWHP8+eBLsJKhSN5XUUgeELU746c74esrxQZxXH
nfN0oa1XZUxc9L/HvCPQcNYvSb+HcpzIYcg4X7nFR4EArLqSD0LQrgq1197wPsFG
O7ktJI4CvUAebTBCgv0v4y4M9PGqT3BJQ+0cvYYpnXzexdANPJiJGcrqBisDgvPc
xUh6twdgfCn0B9s2nfJFfcI1zciDXeAuDRrxRWZWj6yUiNI1hFgkOk/hXeyDNv+s
nisdKcTuzx5jsaLHG6rBF+IXbZvbxCygiG8gGP4sYLeGtjcZ7tHv5zqqxBAUOrUN
nTtcm+cYWUfikrz1LeBG0+cNECUJzJ3Tu31F4uzvt1dcBz0x4FwnVcZELsym1/wq
tpB1z6Q2w6rrJ5Fv4ajP+s+6ZNRPN6RBGes6JNOWn9OJjCk16FUmQHyGQAY1XyFu
m5Mx0rPKJy15TwosWLet4b5Pm9uw8P5UnyMMFeXg+1C8MHsTByjuERYk6Ip5DPUc
5ihDEf1q1GI/wD28f3aBRQkHFaqRYS0QWfyPvwUG/DXDwWc1mGNvnaIzvT0uQ5uQ
6jz5zHp03c5ky10zFqYF3K/ovN9CZOPslPt2QrdrkwJ4Gplzd9biv5GbTxqYT8fs
/0xHoMT92asgqgFV48v+dJ80MwPSTFnme3FAGbPeSivG7jyr9HYJs8MtgLXl8/j8
yW9PtalnTbGDsc50c5kAR7igyGQ8Ag7tzywVCT69lbPPh5Ifklr25IJZRh3vh+ml
SjQesOg4wnJtDJLXG8QeWYmDF+SZrizBsgV6etNds4yv7BrEUdLVSJjD4f9kbzHx
IeKspASRxtQGAyy3ChwZBTKKvICEsV47ecsvblWWa6P7F1sJTcrVw1FO8zN6+8Sc
cxn1ViRacNj75hJwa5T6ts4hGoLhvoo3L+tHOQ+j+I+EY51ywhKVMCvQNxTX565K
pClaeD3CmPZLazBF4vR0SVbWb/lbZ8f3kBi88igJ/clJrCkWq7iEoeDnz3KHZf7f
X1ltHEr/UmFwNMnjlDR1mB1+LWdsTGUCx8/rLtcRRakzg4LkWJ9x6JCSJI5Mb2e0
0Ykc7XgQXrl3pCXVmlm5Ai1QWu+vGRUxqXtt2FYg6jAXS3VqNn49bGP4s7VOmNI/
H3KGY9Is/XnIXj7Dv1rU5ktluXg4FYLktHBrWu5OOnNSLcvu6Do/7SLNCW40SIE9
ZxdWdGorAMGAA3QXmFrq9zX7ol4eTm7o+KGrFRGHU8OHTHmsF5VPe8ERqKQxFhYA
em2IvZWWiLA11WyBceqA+uJPFI3TnGMp6PthImHGst7k6UgTQZhzas7t9RLNWCPV
AEz05/GPYyGhpkIekn4rjhfT7IDas7TcW2wYUPi09jVjOL6S9b6RQYfMNlZGVRIn
zHtJra3YqWxMoISPNUBVdHHi0Puoih/czTuj9SuLTsYfstuO67TkvLNYupuHwBLR
57yIhjInis+lVqbpZP4pfCxw+57ptKb5pShSrDoAQrGiC5Nl08NAq/2IBa8Q4ify
FGzr2KcU9i0KSHGbJHofW6Lt76ikUWU61HFmDqeg5OegmTbZu6HZb1ANHx683cQJ
Fz3TJv+4XRw9rtptA9UUb9gKcv3wLWvK3tpRHzZRqDUtjy0JjUJ3LN8RmM2Y/fXW
pXV8ew0TOKupVOmWvd5JdlwNZhv4SLe1V8PMWrEe13DhddKuY2RjKCYPUXLLs2Pe
oaxxp8LV9+n9Fr4Z5gJ8A0Xa5wFgOMN//yajj5n4NBoDBV7kJGbNmAcBZIOem28m
LobpRwRiHyXcyCv6W8ze2Hm+UpuQ/gtokm3qtYps1NZMRB6WKfKKULw7DrZ4TGeT
dKCK24HSjg6X0UbT8FJ+UEIsLblkj+7L1+bVVw158fmn9SP+DzxKf9qAlhIWr9Es
J77g3kk4boTB+MCQ3a2wJM1PTjf3+L7DLg6RyxmP1WPoFgpDIoeDyPqmRxrUCZ6i
6JJ70Fg73rVz8yYdiwaWPH9zYaaUh9qu9OxGSdAH98rx5QKonk992G2+nIBw72zZ
pd3O5KZQrf0JdYWCq3OE+usF5TIDKLsl1m+rN+7Sq+xFD95KOyZuQJQI9m28RmNW
VABEibnvBxsETx3Dw9bSbxcfjVVIbKV6A5m5psOOMCEpvp385iShyy4BlTB/RrF/
SNYyL7mNa1Jb9YwrVRv8rHE+7n9VDf0+Facpj7GFsyk0djPDc0gxHsZ2zM9yv9+S
tHWrcGPz9QHN/PEHbAe3+WkW1cPot/avFzOiXre6CChVhAcKZH15/D1I8boCJkRB
+LOWUR5E8LTODtmMh+5EdrDDk82JWmikECUHrkGMx66UdIdFtjdXEdWYtoLuoQY6
DcdDIlbyZ2oz6np0wP8tPHSCzvLVD8jkFCUq3dQ2QgGpCfh2dPkerbFfOaKGXuP6
Rdj7HVrrPArSzfhnPHjj9asSmCagFOV99W0oA9IyakzVh6ozWVLQ2ppza72dIFz+
BzrTjqvWROJJMxEkhGfNZF5ONx48tkYv7lDfq4EChnkv0S4dmJLNp7xwqgzI0bXZ
JRdim1z+FDhoEb9cPyJolIeiAGXOKJWojUxr80goZW6Oy/jG7pkrjt5FnhpSJfuc
DFB7eAs38YYKnSs16f3bHIDOl1ssep1pVcVCRYqqayxz/hbR1gBYzHpmAf58CEGj
Adi0TopjZCGPMjus3ZlafnNPFCLZnwqahjS/htLxN1kbNJ93QCfsLzhlpqVT57fU
+32+FbqP18wt87oF8j27L944BebFi3APvrM+gn0UkxecKp2zdRcpqp6yvTeHc3In
ZPHLUgSBx6AkMJyIqdjIrTmymh9Frh4fH/Tr1fX1OGGpUSUbA4nTNGSD0rvDpn8U
/yXGb0IPRnWiKsJ+v/Xrq6pc5K8UTLsZ6VmBs6tbmsRu7eoBjBrAkfnL6NNCZ7VN
4yzWycm0nBu0KcJbgPhO9Pddr0xyn10MKCNE8JoguN5T3B80QP1+5ZO40jS7aSan
DjGkXPvk4VuErC7/iI0ODEH+JsW9QokMcsxzRI/9OynqdxnLgIIm1MkyokpsGdPT
TUDrCzoCiIA+WMuXHst15vycAL16HCCamFEnnl+GH0pA3D2/dap6rvMUv5pbnP3z
hmOZ5ZfsV/0pw8YHgk9nC23zUarJ0Eg7YORZKAUp88FVQMvHwrS3T3QFrN3UUmEn
YhrnUala+TA15XpZAztAH8fcGI2yBAJHilzUlTLIHX1aSHsEmQCnN+SSxhYlSX9A
hD67ORETTgw3AOl8IzGaZEg92zndWdfTigW8dppmDIMgJLsj/4TnbEJ7r40sprs3
n0REid2rVdwNDRQvO7msCEOLktFCOwGNdO0UcP5mFPuYCqA8sMZvPiqIOEXwFLzE
Le1U/OgYTqRdKbPSYvRdZn+CqCbYkpGsXvzDJL4yVgvijyvGHa2W0xPSWgBfzRaM
oNtiY8cwUrA218PAgUpjAbQwB5bZBktTQCyH+JjJdNR8gaVmB+41ioXGx/y8RR4p
9PG8mL/WHRwwYFWSk/ej1xi23jI6qcJC6kmpBpF/EA+KYjKq+TwBAAZ6MZag7Fl7
b+X14fKw0OEj6kTFY5M1NmuGSysea4BViUwGdVkGJtErug7be/bZhqm9z2jpQm9W
+ZnlfH/0HtlxWuJ0osdrgA/fpMK27pp2u+mDyOuIEe1g5Vi2eqHzcg3/JSFbTDQk
53GBK36cftY4N5pEbhHPMRNb06fC2imx9jVZVR4GkXCcSfLgwsX5MD0eY/7IWdkk
nSqEKx+14v5aSTnOjaqPEs8VmfjcDyWAOCq9sgq1YyImB6DfSB+O+oZTz7lRGEFl
WEqXnhHI0UYrnswcWVK/TMHEBssopSyUJwYeUus5EhokeH3zc+VuxbDuG1zQyPPm
QOi2s9KKPP8USX2uPS5o1zItMYzNSpjCTR1I/H+zPnu0ioB9RmzCZ+F3GCDzRN7h
9/xlNs07IiQrIab0DLkNaueRxjD5/4+rCSjSjgL260Qu+BbpPWHiEMjKshyxUJE9
51VntQxn0bvbf7ckiOwFsXBN2Ge14x66Du1H+qLv4NGbUnYX034MCaZRHJVxjIad
rKImQ2BCIgieeLCLrv7UHzvJLEcJTUbhK1Mt/UHjHoHwK44f1Qa0Yop5S8WqmfI6
viqXU9i12kKiUzIfSlG1Yd3g64dCQLCRi378sW071VsAkAXb1X29JujleJIuVZS3
fGqb7aTaR/3wiIUqir0UTx474TPXsze/Bb2VoENqKrXo68NFHHPKrFZj8M4P2Ixp
bWw4GnaIDhIlGxE8FUebp4CdVkCftH/HFbFupH1APEd8w0J9eCXJ7q54eUCndRvo
pLvXBSBuThiAGgj5SCycDf0aG5FebcfcvFeEz1gnQEqQDRLjLIwGhyxZVhNP3/M0
64IehIqikLjQMxVulnG8/6bXKH+5IA+jAMaLwaaTBXelLjIgKSeDuoVVqX4P2zaw
lrLVfxMBvF1hXfZIfOnN5TtgH2C1CW/avETzaiYoVObQmn/LaQncT74hq0yf/0QP
Irh4Fmu8LD88231+mjC7lzqaEjQCq7+wLo/7vbQSbwxufZaHxpwyd+fdt+0q8ne0
byhkqSX8lrK8usvsSvL2svMlIqbrm5HWHKi9bm4dI9yIGbCziHtKNS+IfOJd5htb
SQK7xnses2WwU2e2OXOL3FiFdJqgeeosNkuY0nrN0b/zLCy1zZGbCQ1i332cV4Gn
cjnUFoIXV/xmQnvroHOJ16OoAi0xtBAsRjQsTfvhuqbCQV6Go71rKvBwFVYRSo2q
hnFAT62oSI1MOkldmrK69BFt1G6jaNWrEI5oWPcrd9MRszuSUAlc9pSgbk23Zu+R
dYWCmLkqj1cB8Nsf5FM4shn0pK12Ak+1TBm8HH2zBpKPWMpkvVjEglyqlFHZG2/Y
Is8x4KuS/SemdDHJAV7LA2ncj9Qi4Y2ZCj4hHq81HCMK+W3huWphGvN2Wywt8322
eRc4acJAQzQajsb5WZ3so3d3Qrrs0SkOeiWoaI4WRmEtCyhZZ8E4vYyge2ecmvBe
KqHMkH4ZKi44zHIhrbvn19jxQzrdY3IbkYh4LBTlHfY6u027VtEm2qAoFsw6XK25
UO3tiNb0tVFffq+V9T0VfC1mmgirjc435nCs4SuJZvWjUREQrTKj2Wg9sJx0YCPz
SmGt6ySK9/9JmaAO1dIO+vwb5bv7ZJuDvEHesRCPnDb6zDd9qQAioEGIEbd3NXpS
v80iswX4vJ6zobc0dDlovdef5YA+R7GU/IbMa5Y/RCus3y+4i7yvtCSJGhOsj3yu
soTLlIYIEskylZnGxpCx+9IOIGAAHBD6yTWa+ud0laVskju4xe7jzy28aRwcZkpG
b2GUnBgyWBS6meZ+9wBQTTZf0NHOeDFwulI/YPgGIfKM5CR3spRQ6ccZ7btnVkKN
C8Ys/yddQyV0nkdNGJdiXBUPebSvKo82iwj53+LkJWllTI1JHedslksmWKs/eW6F
APxFOOXgT+rRSt61i6yZAZQJPe+y+VBgVFYjV9wDtACAkFibx0ReKsXtpD2b3llT
ecbJUafRDn11h8F7u6T8kcl/+S/SO78LR42btwJ3S8L+1FeO9NwUcs28Y1ObctB6
M/uQ1BJmeu6VEnItck5Y0IDpKyPKu4zWpiGav+dK+K1zcYQo6rKYauOlNGosVew2
x1/zm6aGg4S7KCgX2G4cDmNLHfkgYaPuClF6TEQ16Sc71AJ1Md5Z/mMXqdNrwRMg
1FbQZSW0huVqxNIhpbpbxbtaTQLuuF7bCfmVFo/8Gbtr8i6ZVwyNRHe2WXVmMxlb
XgCKoojR4c+4gRXk5vOtA0kghRo0g32avJmtZ3TL0GBw02+RXbrfsVgDbP+zR9yp
XyCko8wzM4fPe88oSKrN07qGWCL2Z+knE+Q0a/V17ocNFicKuMA29zi6aVGgZiQn
ij+F1mFaIaiTcFR3xXjpnL8SY+U5v+kqWFOqMjRkJSR3t7EvBs4xvw+/OkY78OyV
snU1cN/ukDtTnF/8Jn/tLopz8cC5F3O/XYWDIg9e2yJc7qd3IHMmeK5Dtz+LiTRD
ZuVCS7gSVhVxuJLdKH66veTQP30lbLGOZvePr2xDbtIws7sHoWvnj5d9PH+q6r4/
QTNgXVaIsO3ljDt56Qkr+kPRsiLZ9eYJX5G0t1ulRRzb4+I52b2Sz5zfZaM1eDt+
trtkKi5GzF7AMzKMW3wemP+S+XZF4df+xtjCyYWoAkDtBslbdNgrIS3e0qAMv/GN
e6cteiX6VQBVaefuUUQOB8tUsk4ESDeM434K7ClAbe9kLT45T1ntpKEcb19klBvO
WNcY/e99zz/cHTYlU6Qssvub2OI7+JPk6XVkCccPuHUcl0wLyJ8T4TNSp73Kiz86
c37CWxF1N634lwuDkAoDe+EQtT+1UQyLTt+KOzZL0tKfSvrGgtqjrrJwoLmU6do6
YH7G4H/7DubYxGevF+obro2j7kuykp7w0ISkzcsd694EJJ7tsh1iKbtkXEPR06oH
GB5Z0CgFpE9jnmiIcpfHwRMhX8SV9CStmx+isEQDVRfd9gj/CjCCRPNZ/Dn4R0pL
FjQeDdISDombDVXX1uUYWq+k4fXlP/Cq3pjIV0FkCAj1z4WoJ4Jz4g7fYtFov2Uo
NWEX3V/NXMBOaX4mzm2y8BW5efT9GfB0QyAkiGF9V+jIEC21ExHdQCM2scLuwajK
Z3Ijvp9aAsDG0I3Njo1axUDpK3lmUDSNuQFZaJVTKQu5VYyF5U3Z41qGiJ94EEGK
7Meh7LXKV92PIQXnDa88tSZ9BRnw31fXpLZ/MpEo1tBZ6ejROXiZMBA5JVjG9+5Y
HsPoE+r8eJMXpQA3CC0HQJvHMZyi76hIu3MVPaR5AOyzU7mxcSwQXK5VpEmHczTx
JtgBNp1gXGlczKSwkgZrrmDbU1z/+Sw6945VC+GXZS+cuR1+cqY+2GH+tiDquoUs
oiHk94holSD8uJ3604NeQzs4XeQdBk8vLJ5UppSMX/Uv/rhKGo0rkJv+IryculGO
Lbz5GvNn2TKRtIi70GDvnM00QkD83j7vSVjSbwZWE1AJOUfRVJWUyVEz4tUsyw8B
7kDIkcXkNqpQPq/PQjzxOjIXwEjeW+Bgr6n+J9QoPtsHtWdCzjre+oz5pV1mo+Qz
Whfs+rsLkDymgDvYP564u6+RjECfW6pb/ZZiqbxrm07SvbCgvtwX4lMJ/hkisxif
FjgwjfhBqESCvZL5pKsljR9DY8n+hnXtLcloibF5hAwH622WpseWGC0R/MGTwvXQ
lYEV6noiynEE6SxLlOwOk9E2BK/+A4sx+dR/qRmsWPlrZawhsSBOdoxO+yAvjO76
T7/t9SjSmPSkNWU4HWl7X4xW18sRtMPqF0Czq9vYnfyrM8HDg6omNGsk5lnRNX1+
pqohUWEoLuUX8mDBTtGc4T2uL4Bj1v1LG7oMZoCRh27MeOoyB5NHP6aYsHAdvCB1
NXHqeqrUVyIS6/UOEuRuIpdvlAZYHZpEJp0tUlenPkTDm/u+VaNdQptedOGfeOwC
Byd2ogjBkKyMA8lh2LKnHBlqwrk+yELJlL1kJ0kotUzCrq6VsmMDP139gp2Y3/o7
nPgNZWN3rHMRysdxx3vnELGyUv3G1v/Q6dCtJT/0NwEKFuce1m2sY1W4eW1rFJDu
iv06DR/frLRr3IJ5H82atbsW4QovpQ7mjjFcGLHnwtX1CWRDyoUNb4pgBypF8xK8
pY82QB+8JNPUf84ykV6orfd0njfUPaLlKTO9cR3jpkygPWw4HNh2D0g30/srV4Bp
p2MPYHpxmgnq0nNwWCxD+vOS2c0GgdHHvA/N/j+QSoYc6QaeOGpG2SUy/AlJaMI6
KWLUF0eI8y2/kKiJa1ETuQqtxL3s4CBAc1ZLGz8VwoF2bEEytqV41s50TSL09G/q
twEi9Tmf/TMhXlx2De2+OebMBxJF2Q/a9fY6IWugkv42vX6Ekxvq4gGENW1nuF50
mwy1WKbpIcErPM9asYq+kBGh4sl2avgpaMeBB+sShSlSD1Vq1t1q+L1OHhL7yNFG
R+jnzB4IHSltx5lbAZ0yNo20FrfTs6IOIYMEhIIw+b9DOAsO66wNR0UcGTpxR6w/
DVZgX/TvPVmzzHz4b0vfQq9Os1SqNiqlpb8E+5tt1dIn+MWY1kAQrKZO+e1YrgPZ
HVJfMOcJbfLKxajziptoo0MDgF5WIwnzi/hApakZi7RW3BTVuuX5G1corFb41ZSW
3zaDQDzhDkNG2/1SHtEwApmVn0Doby0yrwK8R6DO/xjuy5XOf0+z+Xi1dgE4SCW+
zUM08QU/1PbjoDPT5pX1KqBERZofhSr+L5GJu/n445C2hcrpnL33Db5En2xo7K44
3oEMf87Pru2jTuiz4/+I7qVF4X8isD4+THUzruPlrfq/4JZrvRfVhsP6iozJqKBs
28hZRykmsUgfRkL+u15BD+scHAIEecXwxWDYtMUDFAvCv/7kGuwMCLFVzvTssjDT
mbvfbb+Gqo9ENTgTNhCWjMM7Y8Ffx5LjyQMotS+yjwTONyz4/vVEyBtWuzuBsnll
XfSwiS8PJuvm5pKsGKip/RDlOAHZzRi0ZI40nQ0pViTzIOEmKEWXM+qxcVyJ87PU
RYiVNNZjP1Cwd6EHNRS+B2Gts4D8g+0gCuhM9D2uToypr9MaVemdpBWY1suxN7uI
c91tyIhUKRtBYJJMxh07U29yXbHPGT6t3LqshyuzJw+PzP625PKD7xIDRMzundnb
x6uz9ZtafmWnm8HF3TFuOLrgkfEd6v2wYWzGc1iSXBhLX9ngFKXG5kkJ4NcU8mIm
6b6di/NXnEJRt/TEpNSx3PuyKK5wWrTzb09xbfcLnAbyXrprwEmBRdMO5WcRPD7e
bgRbtnfUBvNuaTfQjkWoFx8aRx9CpIdkPmlKzGL5hjmXOdcP6wiVmkxfK3UBMZqg
/D308f3unBEXdFCVPaDPP83YyCcoVKliNeFSyf+wmaHXBZQga5jCiX/d2jV2KTpa
Jhk2inERBu/XcKmoRzY2HlcXTX4D4jDzwW6UXWg5uqiz00ML/CDzHGspe2ymSv5Z
vtcK7yQm93q+ziJv79RlSkAmC6RwgGjFzNLZJWTl4X2chfggsWxGMVY6dC3zwTgV
JOq/rgpJlPGvUbrNz0KdZrg6wfSEXdGkm/HTLawUHwjfLtKRRy+d1wUgKCdp8xZk
L/B+raCYo0E2KMQzBS9ZnViogzMUViGoTv1afb4Sv1UuFnIkzfQNRI9qQAbBAB9l
XeupRD1p1MP+QkE7T++YJCh+ookbeTBl+rXrn9TE8tsm8Y4JoySufxQVPA0rH7s3
bN94RfaEzCdhZXVuO2cCSQUNjla3DpmOkXUTf/zRev0hxfQBqyGyRpM/nUVCUYoJ
JtY7mlGUtlev6QjR78ctgYV25Kh7ZajaKFcxhPnTHv7d06xAxvItMPOKZo3U/ZAW
NrMjU+NuTj0lO+C4ipPzGpZUVWvg8DTTIgiUJmGG4HZiw3rcwsaexCZlrI80Bk/C
qO/OX4DkJBL5bOm/mlvFnVmFdgdmSVsqE3ON3Wc0Os9437uwCBIBU/JOw/jIak1i
Njfv8euXn/5V9nDi2nejfSOq77EW19mHex8ZlnLEJNZPMBloX180BIbJ49zknnJc
g65zmz57nuI4dNEfzLaZ25zHIW/z1RhK51uE9so3tvN23wWLQXUFW+HFA5rv0d+w
nyXlxgxp/MNFa7s+CbgUvXX9sWuyq7x+njUT0W4m7wvOi+1xANpbTIX/0NKa6beW
jSSiKvcUEEDS1GCo7qx9rtudPeRKqPtulqV/Zcabxk0kxoQT24MKLWa67pilx5u1
6B8xP5T6XqtX1YhGlMwqIIm+ojpqmrJ7xiDrejQ5E59KSSLPWtKNQZZK1+Fs8UHr
dBJOZCxMBQlHavyy78/GAUe3hlEzshkzJpB463VAfqbrsksUaW8And6UeKyVTuwJ
5uT127BW5M0BMUfn/icLb1QFueu5N0akZ6Xis0YnwdUophK1sTu7XX4RuaWm7300
kfm4foWVWdd99QcFN8SVGWZEhPJ+eoJrU2/oH6Y9dgqVG/R9LlF5oa8urKEkosJ/
eqfvSAyR8DJvdh1KJnPMaQAn+0jQt+ob/DfIMkKTPkbVBpIJ7dWcicxnegsUZHfX
x1r2SJ0cJ6OcqzqkIUosu2kZxrPoxPrkk8fW2XuWzBPaOOoa1Q5U2z3eBAkcQqZT
DIoxmdg9DqkLDNVr7SuZpddzF6jZ5KtMyK4kRbePixRb1s+irl+Yu/YPZUUsmVV+
r3d7LCmR7AopVd83vW0kSt9Xaxm/zRxBR7dfIefWljFJ6WouGqcbSNEpJ0mT3NYw
3wD6IDPMlqwBZSvxS2+8M8w4K8aZ2IiXTuL2FUhs7OMetPFt4rS99f8Jpeq4IdLq
px+bPljmdM1ePPZkRJQwi2oTXRqibuMMqtlj6jnfSRrKw11j+f6Ma7SxJAg9jCaC
UGEO31BpA1U9vsSoFDNSPOoE7UJNQ0SbTqBe47jmWMFeA+ZN39Si7lwF+pRFjQXi
wTF15zRNjaoc9wRnp7NrFgWtGAmrxPLvhbTZscX24/lZccPbq8BWOzn6FvyrnG5N
3+WwdKxvUYo/9RWuw82bVutSag4yUSm2iBruR2UT0dcEJA9Q9TLzO5yxKXFVCer+
S4F8lYo5jf0lNfunHq4rYpb00vYAQXrAZ+KWbXK1W7vDi3G/lsud7ty9al3fT/sS
TL+RIw/0NbSbRDLMsTEsL728r6OQrBe1tPIL3wfesCmPV5PaIIdiySTAr0IXPk1P
NkqLQw3uZQqoGXf6Bm3nV6lixm8l2LZLOR+U1oZOj2qVHALnctu+bB8Dok6R+QxJ
h2SyIeFQflnZWOY/QzG8dqsmM5ooARze55uAfzqyRgCSOpOtKdmK6ul3HTyZEKBH
pmknBe3hkU3c8FxDozTvCsZZh02r9fKsASQDKJz8oUzZcGJFWNGPXdgk8lBZs/OT
gHAOczHpw413I5+Xq5uW6R692NqgvxDn9fJui2nU4b9Iy382IKn2ciO0v/T9ZWkN
jbSA9mZ3YHPuusjrUAJab9vpx7n647q2JGpTH2jOEpk4b1Q7dNtLYjfS62tcQd0R
HodABKrKLLVfIDmyTeWUrbSpmdm4FdyQNKvVbWyBqdVj7zdDQwzYeQtF17P+MP2P
weU91ObPv4Axp6KCfnaW/XtuJ6AtzVwXECJl5b3lH5wKnaH0SsIJt32PpugcAPVa
vVOIC0QZBMMGQVlFvXkPOXDKzK/hygMhaC9PjxaE3nN+sHkqY/Xyu/jRHh1bM/7x
Kplg+D0PnTuIrTf1NvO4jg==
`protect END_PROTECTED