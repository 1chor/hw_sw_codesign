-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
D/DTY7T8tuFmjm6a3/bjWMlwLqpMIZ/LW5UOQ66U3k24JHKpe+gW0VmvzJljd4au
CXoIph8uijw73ewKumdNY6TaIuLmB+lkrMYWyAvZb15AbMkNGTAOR3rPWvAnG0ap
TyVP/vTjA/LxFfIvLoWJzRs+ooCTmj/g/QCgcnNNM3Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8605)

`protect DATA_BLOCK
rSH+/XqpNXLjTryMzE+G5JEhFceNejWF3L/tT9mc74JvJUbZjej19zXQPQurIygM
Q0KnZVac4OKvIoAU9Gj7Ey8MXP7mH0vgq5ig4r0AMsMenlZ4zX+9V4mLyAZ5sJp+
yr/eIZcys4KS5ARA6LHrjJsyeRVxR3zCZMYBFolHIIPxs/RAh7i+0DUSzcKfUOBL
n92867S8bkpO6cHudMDOuCEAtfGx6oHmPIHhH7DRH2sO4+OEyEhAIOnCzd56TCS4
F8XPZiZH2ttaOU/IyFBkh4tM0mpTtrCx+0QujkJi4QlyryKle6Bxz7dCUV3lLMBl
nqC9a0XQFbxyA0nWEzWVcZ/WsZtv41Ii+rezApuHQ4G8FvEzoNjQJB7qYzKY8ZvY
FSrv4n5F+MIqSwB2rIkKeQElevhzWDf997ygbvR00x3I+hOsvxGpWblnLOvM2Ljc
I4v2dhHB1+eTkg8WVzni1fKKkP1ivqFHUqX3eV3+ZQcxPe9ZntLYFfiSlRkf/E4a
r0Y1UZV0ao5xUoDjY+55L/w86XzQKrQ9X0sGsKWOujWsBEOp6sL2QmiCPdDMrvSv
mjitTJQTCiKYr8yuvyKoKk0gcotg3JCN82JjKnuy7n5tYjBrw2J2JFuvry6VR7lx
Ov5efaltnvL3qcMfVFg9MEC9M9higPy1EIAPQwe7q/AlX3ROqJDBqCnTqKg8iuJs
C+qzbXHgbOfjIOp/BBNLb+OZ+3GTh16sH9znGMovK+SyKE0McHsghFWJVRILVgJP
nbyCRYek8ZMxRIDBrmXMaI3slLevIMxdlWNCBmMe/biz9tkakX+TF1me/Hgofvwn
jVQBZtiRDty70QjB7XYv7WoLHbRg0sx9nSdDNmm2D95R9xrvmZ76dr4BCvinH3GR
UGE8dyEXzqzbANWucaZeSAGvbSShOMU2CSOg5QE2XeXag1cQU7ze7WMMgDeka215
2bCTAttKg8bhZSfVX4OlQWmhYgsClCqZJaIijgCeKzMLq6uhpBP0I2NRcQawkhBW
/WgDWOCnWCKdeMGOqnX2vIWB2I9gHQH/uj/mCfbXyy/3ZfybFPPIidTfb5e2MH1w
TV+PpCxT30y6F/rRItaUaM110v5A6I/Fel6Vz6fAZyqPCMfsLWE3y4/FHWS/PMRt
lk0mLqVp1N1XlLFN3PjMQ+zpT71SEJy0fPXKs0hhkvfrtbJ5TlE3RPcAAtQNwq38
AMCqOeS7+uR+Jl3+u+Sw339F7s5sh6VcJL3TvjfpJjLC+9LwjdbXkxKSqpV5+KbB
x42jYeSwcocPpX6MF8B7L42oAxEBR08qBWoaoEpMuiNRR6nW9YYv/HxNoZ1RFCFT
CSV1N7jMDkc7KoxLS+ytA/bCv5qHdQIuAozVbvk5WFFftUQaRQmXV3Q2eGwR6Jz/
CM8FYByNJmVjVP+uUVUM4v23lVXyZ8z214yHdppfiuGpID/ndv2XL23Mt3EcdjkQ
vblcP4jP8ahH8hfkl3a9hnSAE3A9PsRh/3NdI9dxoovik5MwwKqYyRPr6BPDotez
f/HOL1mOv06RUnPDGcsV0h1bKCnBlLvb1j4pzSTQqudQnbsIlkQt0Sh+mScxJn6K
CSQZCdT160T6LEvyQ+ePsXsLUAF7WuM5J/XnDJ0xfg49oyrFi1AIGPSL+MziZm9W
dkIwWwP3YAfskx1ba+GGFMzkM4ekuqiiNCyP+trWe2BbAkdlVumGWQzt7BOm9frh
VnXL9U4eFHieOCvuB77+6EzNosLUsJkbukpwvG0iOpRPIsjQm6iq6GiaWURiD5Hp
XM6PdezvpnzDt845MBExkcM/8mgpzeCfa00w9XSNsHbjR/fgtIR03Y6ME9w8h3QZ
thzbTubhI/uZKl4o9jXooUCYRv4yi/xZ/x7MNBlV8RD5ucuNczzHyQVlGHC7MlOC
tWvXpqoq04d7vl2N/a8zOr/46H06FskxaHUBSbYhTHAHl7PpJApDi0evOAFr5Uby
PxYdLsWiSy/lNiIjQrsZy7Kwsi8czj/S4efEHonjKhhhvnm9msx3dyyWQJFgupi7
eTIwYppywfeAziOtcnXuDQT3FGGt/WFe++Dycnq6DrGclmb9/RXk+NKeL1Zz6/82
0r5EOfcqX7yBclmkIPmKnJCB78tZPt5jX4bEY+OZ31vUnpoUR5WG6IXWvx+l06q0
fSYkJLf71oWsO9Nwffg4JK5CJFm8hj+poUbytBXLA3m3IWug5cKGBDuua7HPFdas
b+is5SquH0prUMNeiv3Kmy6Dsp9304fy3mG4I/anjGXw6UCVD9cFVUAyVCdtL3vh
mNEKwtMJvs/fv9B0OG24DNv8//nCSC4vTKqDczCILsh2+2klI/zIzC+4It62rOt+
33OK+u90YwYU4jSjfodtVRUrr6xBtZx7FEN2X3/yfyL++kkHgUZXGk+1POfuBRq5
yI8TdKyRerYxscX9ZemXccL3yOt2QNgv0k5SfIjMmb2Q9h3aueXcxC8VYkisPTur
k8pyAVx0rf0ERNwoqZhQYUg94gA+PM8y5H480UGLh6hoMY15aRhVjgbXa58WRS90
bFpw+hdFPJEZ6/GbdSQIp20DMFcfBCvk/xZDQqFERyD2MGNJErrz8oj53vGQtDRh
ju6m35PjtYYn8r93GFUkEPRay9Bi9hcsCmNTnCI/AEdvoT4UkxGIAFfgJVuyPo0z
AuiLEvMWqeAReu68fupXChZLJQFOrQE6rP7KiSHajF3/NnqgvM9NCvpicbIFFGWf
e5wk3qspWOF5mpbVsiC1cIggTd+oqxwOtQwssPiIKStPLMwg+jJNRJEO69lhp1/L
56YPrQZ4YThbX67XXV4Poa14vYX8ROdrs+LWXve+c1xCYpi4r+Rz63HLOh+jUNh+
u22yRLA0/VQG9wsHsGfG/pqLAk66neF4Ws0dYPSP+8FrbUDxuoATdFsSXdGkZ7dp
tTLO7Mk/3zh6KHK1xsHh1WsOJHAvGOaHKiOonUIqUCk0OzOhePOWEGnPfRDL9EV2
ib2jla0hDFOT5sj4+t8IZx+O1HZ5B+gr/LnPbplBThdEaBiNZ5kqLJ9kPJLXzhQZ
x9LppnSKNCylPeIZCBM/eCpIZR6tk7LwXimnSmqdjmBzCygIkAohZoLc4nK5GgtL
jArNWz0/X0etoHcHtE3OrW566r5lbNjyVeRGJylXtQnq9mngZj61Q+vv4Fg3SNk8
xRSFS91Axcnul7Hdq0vSV0Acovj3FxDi9489ZGDMEUYY+MfbYq4LzVvMWQ+4w21b
xrcY96FLhsVc1ps0jwqQ+PrKO7uEIww3pyCKq2ZQk/8lSN//nWCQ1U53MpFGLvq0
xdQr5aqg64l0C+uTo0CX9gvgOlaJt5zKNCIF83pA7hTPr5EHIMmSf/wmnJBxJiNi
Z2GSY/pYDCGBJyUOzdo/z97VXs+Q80KxAju0lmu7b6SSWpcrTj89OLd0rgHrtPSr
YArnMnNu0hwaWrkI0lhxDiB7+UODnZ2v5lCwAFlsAL8GQulxKhCUsg9ZgWfHAXdJ
Nkoa0xCDwZLHb4JBxoCJQ8R6jyg16ZfpGzTkN0dRq1I05+h2K6RSl/Fp2IBarOkL
iiMLpalKr6OlAj7NTh14YPCZ2hM2jpLniEkc1hKW/CpEfMNVCg1x66M0VGmrrBv6
LIlnhPuQYF9t3Y6Y9t52E9J0UzpJqRS5jyUNroSFYe83TjexeAFhAkJwOXljYPgh
/gTnd8kFBS7pP/rpXDFxnSq95BSz0w2G6HfHA5RSpCR2iiGMEQ8pxlhTmd2cg0b+
v/cXo6L/zlrOTXEiSfVLPkGPvi4PHGwESLaUYMOPgls9yD0PpTMSMSBC4QYNqhGR
Y/bXFdT2GvDa1oQOf5uNcwJOLs3gUG4fj93ZSE/JZRLmMecwmRfM9b8k8o2rN6eA
WGPsIxSPjfK6bm667GqGOxqZiSiyJDMzliHSpJD4rI1ubcXxQFYbyQebpD++aWhI
oBACbq2i3W9ZhRPeoyQWtDYYrl3k42erWy4NQzKlZZQyng8af9u+qMunveWkL9m0
mA9LGGBmjZNHlCwtrB2W7XN3ZKST33Z6jbc/+cFUwHeoVtQp2vB4c1q+Y7Qq+Lyy
rcxbZ0kQ4ApG3o7b3fqkhNLuniAh2CNOTYIoCCOV0Yz/0gKtitfMsz4ju/OfrJ+G
Gfh/q6Ef+jU3YIIciS7qiDy/hXyeQtKHhkOAq2fXAtzytVXNMjXXovQDhs+eDvW0
+3B062lrwjAPPKG3CrcoScUNszgqPp8f9AsWo3Vi/pUrQfwPV4tBj54Lj6kjVlCP
kFnIq74ItHEB+bQNug5nqU4prIdzNZxa8RjYL4B2mzfS2Wnhf4/mbQxWHA1/BD44
pnB41Lj9mIzEe7/ZW7APbDFGpxf9WrFeWeKFgW1ckIQps1LjDLBQCcHDNtm9tMDa
IIg2HL45eblQZVv3h2vsBVpyChMI4NQUZIJ47T0BFUkSfr6aZOshyuIP9pZBFbLm
VVP/kHOBFK8IU4ZeMtfnAT6TJ0J7DvujgdHWeS46Je9jAje1jnwz4JCUSu7CYx7A
xwoi07oGtG2HxopkLujt5ZGpg1vHRYUXSDs6NjppFkXV8WDaWxBtP2WerzzvQViE
pdeVUKg3kfGwPhD90/+Bq/79ha7PpvXox5ESHtpys7E6QsyklfXfVNkWjRrFwB1o
CElZi4zXh0+cnLgvsRGIX0SIXqXEty+4ho7QlY3OQorDFPXv5JyO+paQSv6JKGWm
YFMbD4MriIOnbM9TERACjsMJ4xFrRL7AqxEBqDac96A6QCu0KeIHa66QC91TnSud
9D37Z8KJt3POEykYcEVumjADlpODy7aJKik/YJFPujdJ/faEvFw7Xan1IOBUzJ8q
bQJiAXPTuhR8nAboZf85Ux1IlxpdwAQ5Y0n39Tyf4huApCkVhCtJPMBT5zXKSjNg
FY0iRcVkCWQ3tAhpu7ZlQqWhbuOGI6zwxl9J3Re5+4A9ZHaR9HtIRjW1iiBJc60l
LFvcMWvisPVZ6Mscgjhf9gByo57h0xlw6dNQhF64v4Tg4mCTpqBWCgmwNCswd60V
tDUMCTzc1BVWpHNAiQnkDELxBaYqwSInayHkVAouS7UMGRKlxOxwN5Fo30OtrR4t
OgoW78huibtZNkaqPf5/ezfhl8m4MFt+p2pCrJGnvgu54bzUbbH3TjFUQDJDrk6M
rJOIkNUr9ArMu60Blp6T+dP6h0swyjQtzVlJBZiZhNcZT6TR5WDfALuhs08exU+W
GSQU+cVrTMq4ndNJiB8BU3OS4wZbnazZzr0ONZkMb5NU9c48yf3Rlmvpou/jrV+5
3FDjaQq9sz9llsTF4jxZ4TqBnvGsIUaR93thQUhg3qPFIeLjZFVofT8e9tUyjdsU
FkNM2yZWXAzTYz+1GUlHnNzBdDyZUjbczYk5Oqh1yMezI19/b2EuvFbEA/Er7pS6
VKjRMa/y7RNowIT5WpfIaczK4umTbZN2+LK1pB1zOzo5kTqTztNhszCS32xHxfSR
TxwOOaZRqpJLOEVQo3IWjgD3HCyuQwE9k1MlQh/geEj46c81x77qb+kYGDYylAiQ
3wR9wnIKIGOl8OQpyZ0ZQY67xldaOwcZy2Qf4H/mvOxfnsOfTDwucroxLMO924E3
yZN1QS0WyD/R9yd1vIlF3FftKtBWPqJeoWJa75Wyxg8YqeOrBm67t51wtkJM3bMI
ivh7OK0yTgifnVIcEwz6HmJcUNfueiNvoeOnhMApOYEx/7CJHk4YpOXWD/1tJQCe
H2kjpRgU74lasS4JBY+74DKmZrcTtcOoa1CHpe2P7hAQroz9X3D82geLaKE9fE0t
RGaiVd/vzgsjrbo3CH7O/APZSnRKswEu78nUKSKFp43LJGTLu06KAbUY00SnUIcp
SJSQ6xPwluj4ifomf8V4jsTg+/ngPXY5YzmiDLL9mzOxnRgPHhGbjA/VDBj6qb5d
44xJLGLfM9dl0oKjxfm5g5hBDGO7J371Lyy+QCQ8V2DNxH6cbyVnAbYqpSVfaUdr
glDzAkCWceV3+939mJOHJTyl3kgFtW1bpNJOrwVHyUHKGGdBH3M9bvYAyuOih5ij
q76ILb22NGur1SUX1tntOX8tFPGPcWIo+bsWrDe2ir7mVTfcHCW+ZyXFq9O4Kh/L
dxqleyuK2UAj8t3zwoJ984H98wtCgH6R2F/xKPk7SzruBpHutbDCbIAmU4o1XnsW
xTk5wx76IK0B0QiCrbk9GM6uCMvBsmTrrZi0NV+F/i/dY9P2jijPyJM9Pe7dAzVj
nUCCvoIFXgYhs7W0nFWA7cyCK7DhMxDQNE0kHLBQhNY5MOOfB1TgNBTGmnmoHBnF
UkHNiESGkqBR6SJMluIbuXRAEvMmGMa/XXRaZ36duM514CcwAQjb7/0WkVo6XKeZ
RUuv9YyC/RP/7UHTIjRiKOGV4/H0LqQpQBkcxcEkKPss9sQxa0Kxij2UnVHvbpQh
r4mjqmOkX5Y/IfsejU0kUAtdy4PGpJaRbjfP46eIdTCOYIXtOsYj3XNFQ2kdY6oU
ZQns2690K2mJ+drd6RwWhV6j/jSteElz3VcG9YcW+M9Vfecw/JpLCzYH0ZvljhNi
GcgTyG1/WhKuxXRoFR3fJIyGKvzr9LTeRum1E6Ki7llqYVR9VQYKygGXfVbsNdZe
8YJ+0MMt10cZ6vyKLmv5gdbF2vZ+b+PN7lpWYhSX1+AjjHXxlppV5yIOf+VT6AXo
Pk2DuOxqOO/l9gwxWiTPkpX0B2rHr9JURSNQeNfgGnJhp692y7+tv/Rps3M2Bii4
yTT6MQqh1Y87q0Jg6TJYn+MssLcb5bi5z2icy5EniOBo/yP7/dDhHhf3P/0YF1UR
LDg2AYbrkO+CeExp/vjo3nX8Ry6bTJA/JNjwO2RSw5+JVuwqsOfn2ESvVFgt+/q4
23rjbWTZkA/SxUToOYdVuAn1eHIv5dG778XjB3lhkaLcrztaHeIKiM8Kbrh8v+MO
5aC2HHAOjIsDWP8UarpJcf8jembnTRSxRHSsC0U26d7RswP3VYHS4HC5uMjP3N1K
abj68Li7YOJsiWi+J4x+mCt+oPCLLRGh6ufC280mskyAVz05qDMLI2suMhGGBBM+
mvXZJNwzB2Nwwf64PtFNngHt/+C5DyCdbYDN3PMMZgwhv9oH5cWhmQFsgH/6jyHT
7FqPtnQqTXqmw/X0ouJj41BRiAd+8p5ER0vm/fOtGSpGBy5ruldAsuYY4kOBkQUg
ZiUjHsRZ2aRIIDWaWG0reTZ7EIXQucHYE5+OQhBiGFhS79F5AZ7/AmzKisXDGmfA
GTLBOhW9hqERQQbXIM+Ue28izZqvHg1f1CXPLom+jmAcGIcmm+/qUXmuQMPuQnhV
iivLQjd9uUo36fzHNB+u5ctIJEVphyFuDAtq3pvHXM6v/8hI1ujjtGAFtifIb0Yd
hvkL6tITamqOSxTI5eyuXnJrWQ/YzoLveQPwVdphuk0Fc6O8JIuHkDYwXHKk7Gv/
aB1L94vLpPApzidia6Tn5pVLoRAVusMIJA+yLgkLNRUE1wDGYAMlYa4UuoekwBUW
iLdDJ9lSTacONzvv5wPRJQusvlQ9B/xCXnFHYBtAVN2CqmvFUOcRw96ckf8cX85w
928okzsyQ7zjQokHNvH0wnRTe+VYAILFmaXfyIannxrufy7jqmfkFjIHaFYO3rdw
jZKVqlDupsLMg57qaYSRTvxmESG+ooA6Y9tYt6lKVKqbk8JYhTRH4UKa/Q0huTYU
53gpVh1+gwWPz+k209wz20lxokQJ9N3CQYtZxzL28dj1gjvH04fbgwqwPwVcFac6
YciIlwoplEaZvNjOIYfi1y6peXqv0rayBfbBKaFbs7v2XKIOg9xA4G0t6bpBZYsB
s5dsmqIrJxkD+KIcmwPzkMyB05oJaLeOU7259CnDDVeu5gd78euGmFQyjSD3w9RO
B8Hq925bKmCKd8kaSd/ulz17XN741IEJZKyDPTW0JoNPgXGwj9Co+9l+1YJ1u3GS
lc2N3woHXLXZA2LjmGIukDeBNTvzBprKSvr0o+wxe7ry07X3qtLhYpYWAddsTeIJ
62FV0q2p0iTAetfpBAHUacCmrSxHpDwOCTP4BxZCRwOhNxnQIxGJGWNfWuhww8Yi
VqVdnLV/KcDOmkdhW4G59VOeDWlL/fpSrLQEuSL2AP98ikV3EfFKz057buNnT35F
NjI5xB76UXSGVBiFU2qCbDCWx/4n3zQ8xx1N6awoCvvR5jnwaWtj2YRTtt8hY4A5
yTE5py9g+8pSqAXEuSlkk+7T6tMfyEekT9xWsy2nTMilUk5Lfh/LU+ruLM2zRkKa
L2yX54+Vivzp36vTyUWf5XsVvT7IVb8Yc4S84dSp2fw2ktQghriujKxRmT21lyph
pudVt6TzMVeJSePY+ScTbCH1GLpDkD24/u8yIKQ6yw0BTJ3wU55qrZ/IRlw6R+8T
wTMcVjxKmWNuVGbSyg+InBNTze2HzRQcL1C1ydGIOFKeU2Rgx0L8YmajdM6bYV2V
GeFKG0dsR/BZEaUD4E2FRhE0Zj0VsEiqQyyHC7vHSOYXD7DCu+6atSf2/U4DXqpD
j7F9qdDtcDhPk3ymqe1K6GkH8oedjL+0LC3fCsq2pZG3Y2WH1Gl2PllOLfHzjIjQ
smaBIIFwyZ6b9/7z/nMb8m7xnf/Bx6D6O6GGClN0fhMHpCRNkiCvy31Nfl1QuO1F
IN4QRn6q4yMmZglEhMDMChi1HbT+qNka9197XDtGfZVAp/ZtztBHWJUj1k9P26Um
weRXPJHEm7UVaUrALWZsb0/YE1GMc1vDaQE/OOMMGA+F3KWFu0AY9xYefk3jr5iX
fvctzsQn3MGyJGUi7toQYI9F7RSCVqctcQYKGV/pN/j+AwCcSeq7Y0bPyKE4LqvV
N7JOjyuJByuhyAu4Hs0buZ6kBsxGVIpk4TrkNwxldvVwQXMUnk8Vm66obpVTPDuj
vwzR5Al8SP7xtYH2Kv5lsbGqiJoi2wfSpn376QeyOlwFjffbBz7bikxY2RDBEdc0
B61PiCD6P7GSvklfva+AOchM1jjkgbevNZaupKOZDLJ1wrClSF3Aa20hSXZPqqGF
SPd8gCEl6EF2jASo3LSk/4gH2pqSIW1r4uwLafk4dMqfKY/8tNJQddoraSnqeEni
kiwKnLZSUvkZtv+aVyjptqLVlzM8C9u+V+r2mvDn5eSsqJ3klr0q0fn0XmS3lLei
hk/5Vjy7Kk4phfl3Hg8u1mkgRgrSyL2JjSks8dC4NhOysBgN1129akDrob1Sfv23
sHjzefgzbpiK9LaPiAc8HWt7gTS+ebwwMyyPNoChwmf3JeW1bLHQsiVIFOuANG13
2cy+eOVrwJtes5xWUv9DuZg42uoMFta1DZj15ZRfJQDFHIy552l/Zzq4L0dAnit/
M/oz41DDD17JyEhf+1w3FyIzno3FJRsY81ZXnsAaD2ex7Dybgonr58GYRvz/fcJF
Frj++9WF36WvDFNOKa6fpjsvJzvCzaozdU3jq5B7LH9Ud3wtry8I5RXipyjE8tRI
RN+z+tZkJIa4pWdNcAoWgftmBeg6HTqEwJ5kw+AAVugiD/3B9FaokuCzJw7N/ZSP
BuAc2kEPZrvL+vpr9Kt6OYD1n0T2jOHI67pkuz8+4sfhvFivhD28HPt/xnTe+g0M
Ji3qRnlw77US9R2bXC3Y6dVQ0smhfD6RDW8Fnk1yilHEJc7AZ8isYdk7ej3x5Kam
fTKcXfvwvCos6lgZmraMF+2syxD0YMGPy0mHKyy0cmo/IkRJZ/8a1+oRQM8qSdHD
TgB6ziUKXgOEafCaHkRnQDOOijE24mq3GC2yls15Yi9+j3IbevXcxQIZyS6ebcPZ
qo00a6+nGoBFF86WoRfFCY2nSWZIAwj2tw+lAnGKO3wO+/PZX/ZL9yYNHGMJ+Kd5
fb+dxn5RYm7Sw4P5MsMoeMWteNYxKSEaRpwdxASICnTIMbzLrf2cqAJPLNWt6Ted
nVJ+SNjPFMha3V5IX0cI68EJOkxLaRvseNOtZF5nJE94XEwjs6MxBp/kE0Z8qBSn
H7zJcj+ETsDq+J5Xcrdr8JeK4gHfWyOTqlpvcNXXEZEQAYvkGargUmmGlwMkDRBA
rp2LSYz0fH304cev3gZprVhUGg0qCbewWlx9jBunmtMgO6vzTG5SVAvbKQeSWxbH
LhdBFJeAq253NV20uDKT1AwYaj6Wc1gpGNu0gjS2cvc5gmyE7WPDJhp7Qmxlu2jm
sbAGNu2WIC9O41BpA012W3YNMs4fjXZ7ypotzI1B+Q2v4+Q0fkxON4bKu70Uj0t8
qff9IxYcES3+Q+TEKiXDRz3HnqIeO/4ozvmB06Rh9W4tDRmaF7/xBXZNETS5PtjU
W4SMq4hRe9fhIlVG8356u7lIVsxE/DkvQ7pxQfmHandk1Rpy3VpXsJV+S56DLW+7
o81+qZLYwamxWJD0A9lVkhxXNqDV3hXcodQrVqakWlfqRYWXalIfJK38nAwz12XW
AHhEUPuF++7RfXh+3eFxvZDBu5i2zlP2v11a4t+8reL5ich+N1yetQelqEN6FkZW
zRwv/3arxiJpLannkmtEED0OvFHmkpn2+UJHju90EK0MPWG5vUY2n/LNPguzDv1A
2AXuAdbsxmEPr3mP7A17RZlsoc6YURvOBtibaEmD9CNRkCARCGVRKTOkpNYDEJfn
VYicFZM+Wh2tcCAnlKbdPn72oBMSrR/H+F3VBTzcAS2DK66NOMTMF2QB5VLYGXST
su3Gv1PW0JeAgrnt486EPcPCfhEWxN/fW30r21nyYMLGzhWvDA1riVIigPcMPxAJ
sqLwEFr2CTgh+UJNGnJVef/nLLXFEbWcuzuENO8ZQIarxzssO4D6zRRIo7r/e0eC
UJrvugZgVZyEai2xv3nWgtH0emcpWyEk5iDp2FiNDZgju0aS2RzJoobJlJN5dVxW
JjB+2YFpAps7KTkEAM8jodIt7GyyyX7TOUQylxhPN4wsUway+wlIQIfzyj3JXOZf
lvAmp4bCoCv/gObUtQcUg/kKcsHDOSKtHcT02Saeh+hPWFqKGdhbeGiGuNQHWuQu
WWu+/m+VTKnv1hn6LjFEQSTXqZE+q8P1NUgFqfxLd+38qxxNEpLGsr8Z5/DLSb42
67UVL+kQficb+7aNpLUUArH8bAsb6MCIWLw0/4pcLkT2jVZELX4lrqxobEBTG/he
a/3yL27bAG+lUECvLHf9b5LFavbFUHtOuMc4ZJQe6uTVu+U57OqCslqYweMR6MfI
yHCnxVBXgr5B90UexbronMNSIbS/fOWZn+7eJHHG2W2gZs95t/F2a5NBMo3rHWg/
cDIa+VM840Wrqukm9eL/+utgBlB9fUnVGinwwK5B8ylkHSMgU59Je8vrhrIO1bIF
FK8l9RWgONEaGUYObfRR9DkQ0nTmYsR/giOJ3HShnems9R0nnBXE8ArKR4HLR3jh
6zeqr9S3Ic7F79sKdUnWtbZqI4jgCkBVQCrbZAr1pf0=
`protect END_PROTECTED