-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Tl7Y4IrQqLr0EBQw895qgW6jqGVUARPXiMIsRBlkrxJBb+DN5wGhbPKEHW+E4U5Y
TPoT2iRkLFDeWTox73fkiOjmfsnMMkcB4MNEEkIBZCZ/pMxAlspSB/EoJ2TBQNh+
YZjYf9bArsvfRgXnyyt/BRCYcRklUSjhF2xjGxlGIuc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 29445)

`protect DATA_BLOCK
HoU7cImnrugOB8fOfh1pZTCSsTd6wxaw96RGXm4EKcX4D5GKMhQIJ0tgc9Pv3xrm
FCDzu4coCz10G3YmydDNnEmNSQVGXmqK+OZ3FBBF7a+Jr1F+42KBuGqPyH4HV3JS
hCwx2DMhNJ/8yLyOYl97LcfpfyeTorF4hScCvyxRZN5Rnm2fNPoVkFdoKEtEEM9G
FAJkbEck5CfleRGWQRxtodoLRn6wHXCZiBwiKF8fbUnEEkZeSslNYnumNcxme08T
84YI2MdLXwdFmCGU2aozYe523V0+geYGa60L8T1Kw1zCLcZ+r1vON8Mjs0IRpiIu
4l4HJQKVaLudtFxZ7+3ZEHn3TbjqL1cIP3Zt6MJ5fpMmt0jw1wrRzMcHUvvA6J4s
KHaykELgkdazL7knFiAqeI8R2NdAZ7P/6EfZ/okloeGu+LIkFFwbMZTQznFnKw7M
269LuXXkR/Hp2j+1cThYZwNRPO957I4POORkIRFaFULiJu+vNHzsGsmkpiWIqyhP
VHC6LzvhGdUX3TgUsu7a2P8WmKmY5yn8VttAKoRam2Oo6qeFfc+YaW056vTALg6N
OnvJA5NEM2pYraJASRMpgbHTXX+GEP/p4IO6ARs3plXIo+1jrBrD9XwnvQIZ4UKr
ouv0aOBbiY8ZFFNcqutTFKByBJhSNyg8l1rx377ez+uDH9k5Aq63KVUM9SMK7UDn
kEvGZgk4bHQ3xHoNe9TbShbR+GpVqMsFAANB9NqQTBbqoD6Ag6yIxNJUQunpCEQr
FKYwFM0hyi9liUyHC/n6P8qkdo7uO+NXXLh2W+w+GQuvPi7V6hml9l87mgPj80cx
THvf5e/d6FPhsZbjS3Y4KTPYwVG3Xmlx3d8Hj1bp85nRKc1h/aQiSsbmkJElXdGQ
fk33AI+X2ancOyr3sfp0e9L2ulr8nSD6LcpgAT4FpvM+Jpu6fJ3ft5WbA54jHJDK
MO6nG/fn0/3IBoUbk6VhQ7C4M6wu7GqTNNuWFeZH1xqMiYL0z7AGqnloE3gBL02n
cpr1/wDlbvHxRBmqWU3yI/NsbOmQX8FHn4BhWrizYadaEqAs95YFpAmRDkAXXgz1
j+fQAbUFtJMteKbNe5h1sABCUjJFf5fUb7tifzq7acHPXgrgbGiUuYPqd+xsKtog
IJeMEWh7mxY4CezI0FTOJIjz0CO31SCBUg2S1SDMw+ijZbtS/mp/ZS9dcKHdMlok
/szaqFzB4bqFo+zNT2T/+CbFY88G9U6dT46JBsJi6HwXL+ejzaxUcQOGCXYGUFJZ
Wnm4/Qz+gxhyDOlNcx6BBfWN8IrB7EJpcxBLxr2pkVECOTVydZD7y6JsVkKquNsd
G4VjohVnNcY96Vd67G6YyUveQJUQSExV4S5DvcgDxUy4nUhk8yvDqcVrrMnJ8oNJ
390d79AZoySBV9CqTfQsenNchcwTXBfVhawkdr50Dk+NlRoP2x75Ap/zvjHBZM5a
6KZCbypZmvrN/U3fxJ6Fmv6T6ymaxsHXOMQf72TTQwBvvSturPw01Sop2IDX1JD6
QSoEOwN4cHOq13/ydkPmt2dv0vAPLPk86+eLzudMupS49IBKXKb9Cu5jrSzSTVNt
TJQRfiPir8yJQWbukynokygNR15qZBQOmEe8TO/XJhL2XCrnC9z+7uIS4pCrIKyA
Dlg1DpmUR8gTfDGA5uBGmionqS4+/o0jQwMiZ1cJ1kkdXLNfuZEBJGrJb13JEKWI
TG9BYOMEqyUWPkzxjT/JlIycwsSxL1EFcQ4luFRoqE7kdRguN3IHxmGL0Mmlz2At
+BXGa1Oby7SJWMe8SSq+1CDDBgeIgojPrSIi6td8tK8czwrggd6EXXAFLqjuhLtk
gJWLW4T4LApegKXyqu4STuHexAzExuxAFq8s8lwexT3Eh/+LRGXa1dq4iplV0PSM
MQBwC3nCBC+kReo+HI9fISQt83T44magIYXfSP5Wu1+MRcmATFn+D+cQwAvglFw0
PwVBhdwWePdbpgUM6rObfy+S6aun0AIg67aNbid6GGxTW5Xy7e6ocb2h321FXryX
5jyPLqiB+mhte3Rzm9mEyX1q6xhTE/KrFNnZ7PGizm4ZQqvBbyhmeWfOY6SVvqxC
5HT9f4FOXF7vtkpk/4r4UlRM/Rz2GteyLqLqrkxfbrQBisNb9V9qDHK3RtASbdcj
GBTMQnAlG9yhWTcQsYfOQUWkSetCl6m8K+IdNN+mM1WiWZnZXqkbw3Z9KNvrhOaD
YEdXGQFg83gkyB9AD4yKu/IjPoNBZ/mldp3ODihO16nPEfDcKnFP5DeCLo0s9iKT
NgbxGWTW7e9N4F1NPCsoHGdi1zm/Lb7N2c2N6PmfnDSJqpFYOhr3m/OpNevRbmYE
mULb0na7VqvkPyuZjieMtVckQsV6tRpQQUdSs1VZ4NZp2N5lZqFnbBrZKTvLSRG/
njQp/7qQ6gA/fKtYE78IwxhzH9WPzltKLFf1mfzSCGNoWQGps3jcSt1g/wi0coyS
RIkXvcPFrjltXEpLKgBc1u6bjwzVfIp+8rJ71Q5zicqh9obPwn+0hmR0UN3QBbFh
K4Szm5+mDFi9UWYRnDDHbFvurmo6hOUZNtvJ1BjAijLGCzQ/kdR3mNeTusV4giGv
dkxKz/uKWyHrtW0GhkbcyrUYwUClytZ+ed+jQaUXplIKNCSydDIkWUg0BqT286Kp
8HvEVsAxXzQXyvdDCGsBm4sdV7Sncewux9m+6HbzdCX511QX7CHSZAdsMZkRDaLE
Xck/zsmLsvy9gG+LrApsk57ZE8tDXrRyQJWxCDblQEf2YzlHVOBgMb/Ffs8m6nqp
MsRtiWyDij2ERj8lesj3BPyapLiK5cYHD9mHEVyKnRFNd0yQI2GgGS4zcs4mt/0C
vlub6mVSzBe/J2GzkBg2n9+pmMnxr/+wpIqN4CaZwGQnXqB5JJyjJSlddodOSzEZ
OLLynf2I3MmdF0Ct9j2Rw+bNbQv/WWDU2ZRffdm9VMwWN8l2kPy1Mmy4o7s1QmlX
IUxsjC77kUj3Iu7d1FXMxrQeHUdaRoVanPeVpltTBqOLAAqkLXHKifrGUMpLLpiV
nNqOpk3HK+NLrC+f+w4CBPgcP5sZzsW1ghcjl+Nbnp3XXMGgkMyVyQaU46+tXDhW
a5UBbiSSgZLw2x369w0RjHXEiYFZcTSvd+D8/f0rWeij/gBUFmrZt+uD25LINklj
ulbQHRE4v1dkKeEUvOkV/9BsGtQsmmUH+2HbfYi6UPFnax/SFTvVRGAcuwp2mfBS
swkt6rQiVHbWJPgrarw4j2Wu/Xf+1UvKmPOtE6rpQSejU2Bau5enpFDPOl4AsHb0
6XnULba/EeeYrdhqu6YBWtdb70mb6QSGoVgAsBS5wbjKSATJl3qPuDQPPlWeMkvF
FPdTkMYsuRH8jZCG6COnDxSyhaWkOiyiulVW+3pVLdzFt4sgqgxUj35PjyBGLntu
QibStTzKg73kVgz9NKGiq7BtmTpAhWySSDb/HLULmjAyJLN46KY7yBDl3Ik1R76Q
7ur1+9hts00k5ZsoKbmmn552bGZpxKW3Z0IKnTuHxdSzh3QgrFPtRghG0IgRMUlw
s3KtXhauKvtSMIldZgOSrNltRtd6TB0EboxgQidGsZw67tmHEAiaOCOaITYqTZb3
L0pjRnZPiZtwkufaRuap/IfEplEb1SJqqlMfKWmztJzHTTeASFhr2AzE8/R/mogo
Y5rC85Pz1V+YlVofIAPeGVHDSkJLzNbG+6O79ikOzH8t1VbVhRovbvwSE1+n/kSt
RB0ty4IKpgV0yEApvzFgnw4NppCrJB7t4Kp1t1U0DK20WbM7vsNDIAJixLH2ljIt
X/jGGoWoPLugQptZSROrg5LTMZWrPbVTgfdMC+dz9wu4JqLUT/y8EdvLl3JbhksF
OkuLTxgBfTBOziR5gSAwHen7Ni11j3gw9hgBIeT69VbvPoaR0xnxC1cCky3vRZSE
qVw2i1axLbwKFOYGi/WUWHGSaepHl7FI8MFAmIHJ9LsuhOjiSNS2xvGzW75a/r1K
kyn5sRLAU8ULCFOvlajZJSzaUrV7nrpqmGNdatnciR3DN2yruo8lnuoLsARk0BFS
p2poE7ruDHsQK8YaQGBUqXPVMbxn8CG4BvONriXnHaah7Xkwq9flaak7Sx/wdGKv
HSmxBMcAPFuuZR0I/WlYn5bh7WjuSCG2GzI798c4A33c1jfZCxm6a5LmTR0UMKja
LEyoVgyFJZ4mkUu533y1HcgsqJCyMLD2kjrGmhwUmsf5LoAL6W9UuROFV8LZcQAC
OhbZlusOYkLyOEUfYRuWIpKV51zgArDO0/QRHPcotybClofyefn+urr/dEw6Kwk5
sdYhyCRYiWLbQbuzDaqQ6ghMLP2i2H08+GTh11zkCwmn3NbUB2ecUEM17FlIdhum
p3D1VsajhVMyeqYeBXIEWBoJoZHP9n35p61BDyKN3jaAWQqBme++rJ/Uirqyty07
1kWuuah4HDVJ9cfo0n73gkzxpbELlYlfYBlg21gsIzro2gUBh8OZPO5oDIwHTBGA
/6riNHSVv2bwTI0DecD7gd19Qg+enHORKJi/wBWX24+UUDSEmRVdA5Ox3bzvbPYo
nydrwqxFaOkzXpUhUJJmh1uVBGs5NTOvjSch7ow0R9iW3flsFli5OkLPxYwWN1Ka
ZSo20owR4t//5vVmcV2+UgHvEfbCX0zzjmSX5k3oWMZPEZbKLmjI3q+KuGIzK3MW
LdxomQo/170zoi1RTvwaM1tyex0VH5VKzNWoRoTgzKXcSnis5bbcopq0/tv0QA9j
Dh+Qit/APEOvADhO7uOYibbEcl7HmWiW2Pk/xICKfcL9v4tjtd/N5lipDJT+Hc0N
Hcgzovn9j/FaPvrpUHe6sGqLDVD+z5/FP/bi9ImPASDKFMqx+pocngMPBlN6j0zF
jjrwWVQYZ5J2WYJjxzhOztBCZ2kV428gwsQCxbVaNFfLaN7u1QOlZAWS7Ld3z1wq
P/N7A6K2MQS3x8ye/qH9cAXIWtIH+vqVEXVMun8VilhFF/WionDSmd/CsFouS2Ix
OliMjVbLFUu0giBptFWknsH7cMS4x727EKyykTNWguampXRoWDelNE57U5IG4jua
ZaFm7XZDptl8iSlJ/3ZBXJpU3p4DSHaDc200do4Kpxhw/pgYY9+yPeGFNpONapEf
2ucNFJ8/MbPiyN0JC/fpQruvkIP/umOAluvWS/R6QxVk0TmOOKdb+/ZN/B3F1s2J
V9DQxDhEedaqWqfHQ8t/NRCxp3j3L1IMHqWyNJTUUaduYDHp1e2VGNIrvOffeTQI
//bmTiMOspsPuaVbNKJcIWb52kxM16SHuhOz1mas2Df8gOnqq78i6A9G3weGCGsu
Y4Z2o22GF399QKRhOyGo+fhP+1sM7j0ZP56gkOG7MG3j/Z+/GaJgkpU8LGJri2Wn
SnJlQd4rod+BVRv+XY37KXxpRHqrGcSlr1LPkfPV6njUx/2R5Xxyyvi9p6xahUpL
a7c21yDZarhEsYbzvHM3V6J8b3lFcQPnjdYDXWcFkjUXPhIQ3uLg9HTRs6tiQt53
93zdSyQzTsvvW7w8x1mrpB3hlhFp5Iy1kw8kh4SaVKLSGMR+G7mNFO/46oBN4xV1
yRgsIptdTpXv+9YcUeJsWnSd6K4Ir4/WU6kINv9W4Q9Fak51A0xQ0DUqrO5kDali
35tqllFljyLoyNa4UF5mpp8vJBvJn+c3UmvFvBYv3HKoiZK6wKNoMIkX2zYVjKFU
NiIiGJXA0XEVZ7cp333fNuEOUAnF49nfkndZp+fRlLiPWMc9QzuiyNfunreH+PDR
XEmeefh52qCDelXv+U5yc73tYzzS7DFbIt3IckugCqpt9/l8MuqMYHspNkvFjTHo
3JlZxdhpT1bT2Qyj+E3OxjzcTTVWtNQWeuxKNSD/1EFnWzfbARa7vWy6KIE0BcJT
g3ysc8MCnIMdamRQ7O8S3DZYaCvuFxvEvFEuzORWk+9s0ldl5XTvjItF36T+eD1G
zJkgmNTRrG+vYt6NGyzDVlxIqC5T0rSo22DKFolLvzqSMKRmuSVgnypAj/C28z3E
kJ0x1fEZzF5Lh/lC+1bYJLqiF0Pi2oCrIuqtQbBskTrwxl8MJb6OFvN5BzwigowS
J3frOFzWpq4IOHkDVYlnwr+d/BEUcAZh98RwKmT4IOFAxqooiM28YJd+5lMyfvgv
x7XVp/1VRqb3Vyve0lWtgZijx/QnhVMjPsp8guJK1GSOAqPzqMYRal/FhHtNduwN
LtN0Caes327e8EUs07k97jW1cO5u00iL7Houdcj0Q9B+a1iFGmtsenApEEkXvV9Q
SA0bhKdjUqN94fF3HIPoQv/RkVaIFPhLaWzPxhcEjnelxM/u1UBZ7ROOUBhIoAUS
NLOhUu8fXQRNh2XTz8tDu/xUc88YEisNDLos+tKJTJ2b7N1cjwI3LbiOGvuZAM2x
TKCAmwqiCSz4H9RXNMR/0EbvT9DIgxfFc4RYbui48PShQwWr8u36T0n/T5JGPdkv
2Z0sWYMQF0uIfqTLmS5J34ihCn4HDKQPiaY8KoHthyyda3l40mlqbjKm6ksOxIYL
quz5nj2Uzk3sZgE+MEPtyJmSv6wYf4JIWPmK945HgG2kDLKRzdCzsVe28aVSh28A
kpEuqho/NUN9UW/1qImRUXXckG5powtMto0qJ0rn4dpruPLPpraXY/hTHOk1j266
XnKGycOHBdOQ1CEJOCfwIMdtI3Gv4M8A4PS3a6ssaaDGQW9E7MyX0MnXip5DbysX
ihXit0DcG4XzQ0RjRSzg/RM7Jzw4CfXNz8gQMcGLO6tuFdMd8WP/75GTi4lSDbsL
XAYt1oHexnS+U827eEeWOzAsPkI0YNZYxIm4Ultaoaq7KrHg6Im/GOZ1qN+Ou7Ky
wvLN+CpxoW4CjSUgrbWEQEda5MjsSzDbEPb+NLzYOZyZsx0GfRmqTNHUL8pwMwVK
5zE6p1RdC5s3iqXBgEr9/wsIB/pILMbklPTrNRFJ0Tm4hfXqVHE+V525xn1FFavv
C9Zh6k95ETdhU57YXpStMItEyJjgmTE8t33yd0/AWrJ2GU1A5h0Nx1cNWQ6iaqwY
BjptzYIqvVd5UQUjHTZ4l9HEXBYIAkmKWBLWDWBt8fXRD1TR8ZUxqwXSoU8ysCja
w6jNKJCf1C8NsuUAK056vH2GU2fedGeBi057KKsqQxZE43PY8V8dWrFaI28Nk26T
Io85Si56xfWkHl6iMyRvSdHWIaKhEwahexY5p+XTThw5H0K7/jCGsY7fpcXD9BN2
fO6pXOKq/GIcOWgXLM3hZM22h0IqgYkKmrb7Y9b9fmdFo/z8KnsKB6S0S0YgbnLQ
9lFup83YkYAOf0095SxRH51Y9N9Y9JC/yQBz2uK3h6qoFH+mAnD4TLlNtHCICnjF
lTr65c72ZxffrZpO+HBSSmzhjogqoLJ913L1uchCmH/ct4WVIGF6/SjshVy2lw1i
e0/SmIkR2dX3WUa4vs97F0NTEohXEoiqbLLZwcvQeW59+ifU8EEV5hMuGNcrj3Ms
Q0pK9QdhR5wDMd06h1cYhCQTzoTLjqFjEXcII+9W1Chq6HFpPCbKPf43M7QZ7cPq
RFHLYOW0MWSTQU0sNAOTQqMZVNVys9simeuiBotM4z2HwXIvFAaJQq1fRLzvCQgW
fi3yvXeog6oDCerWhReS+kGHhnp+B0lZSmOoIOisw9UAD/Mk9CgV3qV/l0Yw/rlU
yIMC1bjnahcB2xMhcCJAS90fdsZ445ZDmlP5adJ4OXTux8FMPCxdEZx/faIM/M3u
XwkJUPdaq9+CYjNU71/nmzIYV+wuiROUMvYmeOf+3yKqZNeUCc4b+mnnkFl31ZNq
8iwGKwOaKtCY9DHrPBsiJGZKk3H165kr3O6eiM29DGLBlNCkUv43fZKMiy0EjJzw
FY/kk5hrX7kN0WIb+jfvLSzOmktN/nC+huHsctczZdFSImimpaYvt+waQwNyI6lc
p6J1+QHLa0uodH/p57bnUIkPlTlLkEXO4NsYMbW14WAP9H93lIDJjwlhcKsblVsT
d2h27L7YVAfhRsgvbmSgJaEW1wzxEjNmdocP//Hd1S5U+3ERkigDeWeQ8jZzr3gg
ot6pk2q+tgJoRz11HeKFQVYn3/8gRb3ESvf6lmwh34N3n8wKKz77o8OrWWK88UCg
DzYFpBjD9O2DIa5CMk3cXhM8OFSFxGSifNlsIWx7535Cd5H282TJwyJjYRIMno/v
RkGVJTGzzavV9ejN4iaiJLwegSvCp0RwqrKOMdPVLQg+uAjNokRmKoMsA0n50T5K
r24GzGQoZPHVwK/Ecl9ohvZB4wOh9F2AbHJ8bWJOwQx38ihfKZxvLu13SlQJuvq5
hFQ3naXXSYIyKGmiMtsFJx+ckhqxYL4fa/ZiU8iqh7xFCvbe/jHfMYwSMdbHYLzk
eAN5LbZsyHDeKouc3W53opDgzbJ1+iMv1dpuILslj9i61iP3YetMPGXiLd5zv+v5
3ognJuNCXf3EjFqTAwuZ61OQzxeN2eyBEqqyub3xAtZdR5+t36EKOfx745R7hInI
PFS8MqiNb7aCu+ParsV22iC7eevKfqZcf/MNKeJhiQjP4LOSX7KlbXQh0OeGzskQ
uRVXlnm0EAiBFJ0QgflXNmjdkYK4M4BiQKT7IZlJENiDO7Uc/JeXQxfZqbIeu4eN
MV7kWe80xuL0ZB/4+AP8p/ZvpWdwzvkIJ1oyttKyKWQQ+Ws56d0pEMb8AMUxKojN
8DKP7xFCr9uk9OVTdTkcU/spkhN/heJq8DKRNpW758lC7V/FGPhVw1XhXPftgN63
RpTblQmzfjzjXVWKU8VgtXOjlXZAjZjPgxRu7XAQfnxbhyK5awUnfnrhHei5Bl4l
II9EJfchXyewumrCjIedKNX+cMu1zyizYGI3z2EM47lUiLvUlVBBRkd9z7fPDAHY
9iXUMf6Q/RU/jqbj9iTntcDGqZU1EjrCXDsGYiTKjai1MojSUAWblFInOaCoECku
FED7WRY/LV+OwRod2xxMOguWBR/sO/JA/GbE2bSwChccc957froEp0xOkA3Gpr5R
ZuFPPJGFKm8kDcY0JieJYsEWNtzqfBMRVSbLHWYToabDTa8ixOq27MuJIfhjIyoJ
TmwRa3oB/3FVx8vY1mUJopkBIzwMu6fhnBa2tKzT9e7P8AiGDWgsYSjDMpRCDY4w
merMnmfINYP5apGxpLAhr+kRpLRvdZXdsjBsnqHD8YhAgHths3hQplroPr7ex01y
U2XKsFMX9bYqwz9m5v6eCo5Jo+bl4BGeSu0WWzqkWIWhXVheusZNdggFWmXWLQu8
UL9oB/FuDCJGs5CWqoxWSUoQ3d3h+hNVJyWT54MLRogY+iM/bM1bDrHSB2iMe3Bi
oirxgoqztvtV6PUTjlSVZJevkp4UkdNDTAI/RZVt1UspgjEawptDzJkmhorSdlRs
IhEwMS665FWPOwpD8ucAavngrMo53gdcaMijjsVvY3dmbqpG5+LGVLZtuY0CJ8QW
JGNLp5s1GWVn8YeURRHXYTzbWjop/AYMgO5fl1HASULpYb6PY2dWhnhZfloYbn1I
H/1IbUkQ7sdnY3jtkcAxyzOjsjjnIycgs1UcpLzA/oYbvz1lv80AQnLrjX7Exqou
q8hstp7JpkN7gK4a/phW6WflkIbxN9AZQhkXH0SDhcrA/N6M1CtLko61a3MoqH0q
XYoTzjlmIff356Wkm9q3kCDlBeM5gE1f8o/u/ivJVzY89usekFCXvB/KO+FM+cRo
PZV0VdcbJW41lAoAQCd9gJ2qacOeDuCoSlM9WVhSJ2vN8/hYpBljL90vQ+J6K5xX
0RizGEDdu501Y1JgqtiHA/cKhbhM9E4jvkO4fe+zMrvktyJHWjIZkNcEWZ5re7ox
K3CpjTGYR57l20d53n9lsffByLYF/u90FFivRL5Ie+I7h0CA3zJD36OU/PjezDA6
pvsrsNQ4lQpO25Gqr5QT9Tg4ZkSnk6feGNj6sWnvbAJPQ/8R3V9G36X7gFjPOCrB
Gg0SpljIhJWNF/MuaGNE6To3zZG3YJ7vkwb6X1Q6wsV+3njwGaP1hNdFSn+c5pmf
Pf2pj6jSRHxZy3DuW1WKxRiM1jopzqsMe+CfIZithzTDfmdbigXbSvBRjGhI/twI
/9kZgz7wlIvDxrgPYHP3vbGcRlNnUhPB7KTXXdbn+RngDJ4Ze23Q3fPf1old5ujo
K/hS2p6Ao6kCdD+b5GgTIAJ8lMSF31OQfyo+DOk8SIK27c241EUfNJyrw7Uj6F3S
LDi1FoavcoXTECFLzZMyjsiYQCiY6RNc29N6rYSshBL6Kq6F6JtSztYVJlW0Rf+G
qxgDUw8sgqq7AewSLit8yG3Ku5Vp2sbaGexOpewAa2fkgS2/1jgsVLsyHswrPpKA
TkpzaEdsP8ck78WaJjJ2FQPEaIsVAVMaMmHxT+QZKusmz/rDarHUkpbGxyygHKAw
tZUWXkWwM+bC5tsICK2P2O0XYDzApHOYkJ75R9ALS1DLPNcqsDsZdBuTmivlNqAj
q++V2+n6JBQui5XPL5k2A0HnhMZbwdMjHaWtQVu2RfcE+5rTWuLaH0EZwI2I4f8K
wFD5TqVwYvcZtRLHWP9fomNHJYGYHzEHKGGgkiTmqt6Ax3QCAE1L1/KOanKClgZ0
dYwz6gm+rtIOTBJXSZwOnU20WVg6UfSWmh5JmUGFJf3t8Uwv/0c5nFv0qf5rEiBv
yiOen7VAB0asZcvWoaoQWSVY/cHsNv3LRFIEkgOU60NAsMHgkrI+Z/+FKSuwL8x4
bhsy0l8Dtoe7OZ1pBvuo5WRx4vt995uTc23c2fvxkx6kj6VVd4jliFiSJgCuO2fn
cEGWEMRvmVsVCrFZH22caZBPcDqxZvmkvSoy4RuTOD9dUdKvUd5OzdHgFOnKsUga
HG5ONpkBZHF1I8PE8W0+9NlXGFvWx/okum0JU/SA8uemK351f6KL0lCpGTBuK0Ne
ebX67LSWlWqn2inrB72iLmOLV2OaDY7o/R0QxKmjhOeRk/yxYZqoHIuj4AJO/Txf
oKxM17giq4i2BVMq1eXaPbQ17PCFKWSAXirPSjOH5DLEi1G6SnFD3y8PhyWw4KLG
PylduOg8KI0DTBACSV6/fxz+68LE01dm5IVzixLx7J80ikVDux7qkWB+wUMKyjqW
+XtrmeCYKgeVmn54ca7Asul22hRTsp6aZI+bJ7xs4Z1KIxv5N6ooAfoxdg9Td8C9
WOPeOKc2MU/9gSVvirhUKS/0WXnF3Pkr60wHtRJmQAHLOn/C130liM7EHrfgcXEr
zxOdDS/KGwIPLBIrxw9Wkwi2KkMt3BwDOp+XleT/PaixCuOdFDXQI+cRsODG0p+1
GrTJU45JXcdd2Itjaeh/tgm2lXj8mvHbENcW1fZ2Oyz02YrrrIBFwWniXHh4tZ5c
Mz+GhQGQoZZ9m9t1wsOaBYOr4kT3Ugnibi8wXcgCS7QK5WYMTA63aFQoQ8erLqWa
iNLM7wjbCVRhaoDHx3Xu8e1w2KmBgrG542rtLdijSUE3zWxUcXZjKlpSoJwklzzA
zCUd+/aBYsIFQpQIR1tboPaJvhCu/JIL1Fb225dg4sty9QKD4Rjy1FEeXN30+oE8
HtZO4adaZAm/LRMnN2U8wuKxhZmFi4yxi1Zc/9cglyLOw1x2M7inmGH45yMX0fp1
0E+CxKEnuokW1JdXnhIwZBGgd+hC7Kejd+GPKz9C4Y5ErlooshJMm578kXVp03u2
PofesbdiTMsgPX42zJ1NCPPdXUFO2hnDuLxGJeE1K3cnp6FkcNLtCv4sFNgQYr8a
XU/e3MwRNrR4Bwss34hY27pIkRmjYjHHwv3I66DRyK9mldhpgHbkpQVzFDa0s6rm
UOP8crh/7XZKdXp5TQgxCVwGc5GqtgFxZU5jIcXO69w/7K++oJ565JscMs7dJ85+
cctVwCygqaDX3bOinmxeIeDZAhUEXYeXseh0FLUCsoRXy4y083HLjhaKAPmy/Kkf
zskU3F4+TFKv3Q3kjaQoKQRKzADOsian/bbT27j1BUX3+0EFSdZ1bzUzhkrbeUxg
JvRwDZ2vp9aSq9W8Up2tZwUiyzUD90NPgfq/tMCsV1FOhojv0zcTLAkZQy9AH4z5
2Pgf5zt3bRkgHLWpgZWRoGa3zt9fquSHVxSrO7cbtT8QT0Tm57VMIojewX3xt3aK
MQTMkvnQh8E6k7i9i5nsnitNQWEKGRWtSv1/ppnuLe8UIZy0pQpUAdzZ6uYXh21A
eiKffHEyMD3vswDxxW0qaFrWhEOfNeuZ1umpNHYA3haySHiUsjPDDqE+qGVG3wz1
j3LRZQvkE1UsN1PnWwQmsLICegRrwe7C1S41WMN4MdVAlROrVXPuNIpJKdJ5LQyd
CIrpuCxE1XFCj/Avn9bLU4Yw7G+SrcjrTpqQMxU9qZBRHHX1Djz2XLsOni568iYS
lPP2+otmFxvj19kKjXJI25YSxyth+pQ7toNrpTiDLagxvc4olMMj/4WgdprvoybS
Sv761pxMJ4ab+U2gj44O4j95k/xS0mBELhPGY3h0kn71hVeC70UeOLfhjtf7jghi
QthP1EA2GKWaGusX/SWlcoa7IJajAq1EoebWEXGUtEOUwaLq1BMSck2Xcq+/NzlU
XKZmPSs3iCzLV8gFjNcoEaTG4qUbwUb1pqc2vxseeRIAVcHWcIRoKNJmNFyprM5g
xK1ohmVlnCwRcK36ddACAHWXa1MfSQMQ8ICFKu/3yFo6s8WZkOByus7AZ1tpSR3F
25TIIA3ts5n6xj7pdfV4H4a2gPiD3clV7tJh1ylOWPW0KxCPdkLoeQapFpbXRoAe
QHs2I2hkbMTc82R5yWZIEeD6723eaIlLRF/hfJtDxFAPJQD4Oam7WlUf/EOfFZ/V
fBXksZpEg1A/yWOz2X66+MgmBZUxS72lOGR43yBUfbFKSpIZ7QfQRMS0W5I8q8Fk
H9/rXr9eT4HDtpwVRhC+H5E0QwmlGx3I7B5PSUPa7gCPY3Wf6AmB0Z904ezQHFdc
F3lgB46eD30rGN4jyxVVycCi6GNoCQur26M+hiKkC4kegevKyTppTJ/EaOTcK8y9
JmnqojaPC/+hSVwyqmeQkrXjL80kf/NJZ2wm/SGsPwjMgWjMsf4fJmVn7tB19djp
DLAUUnQm12PGzr8xl87ZbKnHq6H5YFb1ezXTSPtKM42GiXoqCQKPFpwbmklOq4DH
mDZaAu7C7KrxUetRsWsBwNPzUh/3G2DZSty4IRrO2kfcicVkuc42/bLQHNhoLlwF
jtXX6672Z0gh6/MjnhYqv/7zXaYS255njtV5ezLXJknuEE/7DFuIdEd0pzuk2AuY
2pKVQ6Rs+gtx1vvPPGiGESsUEQftuDP9FnqoCQ3qEyzyXv2qSWxgc9y1Rf1chxba
7BBSe926iHyrD8JtDBsXxAJlUmJhUlabe9Ap/09dvIlxhnPZF8DSD+5SvHrrfpoc
jHZG6Kz2X3ZCr3OBvbWrAsRc3GXgQZTQVNQvbMipLx37PadqxNXW+zACq+wr0j+w
4VsYf79FmMmhYlf+Sdf3MEFgphw5vdYO4vnGrSIot19M6XDj0/L3/9RCLAUc7Y0P
WGzKaWpy4LSrtc/2oYRYFSiLXddBzV6r8K9JpPs8v/cvIxJMgm2J9RQL9ReMyhBd
tWQUB8gxst1q8sOtiyse+2ywznsqJFiQ4TFv6g+HxiV/vtXCLADNMXHWKH427tzO
cvynQY6OQ/cPNTirH0uh96mbc8w00lTm1YdXiHBC9Qxcao3+x/wN3LhXmUnTKFZ9
99hoepXyGYrzdPbfHf6qHOTsrN5h3lWx7K+lnVwDBnVJOq7rDy5UXnetuMgRvkaF
AP9J8L+M8h+yH4vI4s8vYFrfxsj+aQ36jJqVyYTy/2QTyzZVFTzVrmVM+UG2InQm
c63GXwsVR9fBzrWEprSJl9YiS1zQGyZXV2xTeHPJY2BdKWpsrdpC1V55svTB/EMq
/M37DRHcdB6C/5qdr7KRcljZirFZN1rD04k+J67NPJMS2fQVVa0cbGEiZ6RN1TPX
Wi1VFUs5F+oRDvcuhA+yLET1ud5L12q1S1295I4dA1mX8tZ7tM8E01emSbY2FdJP
u48TJUIawUgpdf9299+bWYFQ96tfCsoUlVcEc9U/WAiqo6/ZIrnCoTYo+Et4Ln4b
KB+JKR9+3wbdv9ABAWgtIiB4C1UceATB7Bp/qdiH4vYDCII6FKtDw9CfEnRb2hY1
w0Ahq8aZdlolWBmVUFO+yQfLewlIIbGSlPHUgzvHKvRxrJBA7QLzSeMxSQRHtplZ
x2kY6tMgnE2kxI0mREh058e7W6UXA10bhon/IO+VruWIhnVLMYA0h3qh2Xzl/stW
T1F3AXfNpE+aXwBpmMzuIKoX9y91wn8WevQe5QQGPKNWlNQkq9Zkw6xxEKrqHSD/
dCqVZgQPG4Q5+YazTn6Gt/pPPkE7sBWOj6t7d5w6Ulhh8RKlSyC0BZiSJa7AQHG2
8W0IWUUaZnn2K5JlGn/4iy2D6nMhzxzCh53gP3ojdVAjtcTRoJ7YBfatIvEsNknM
zMF54NTvZaEtB9A53GExBi9nOHyO5FfdMiN09K0YPgKUeidLBS4Z2WhaguJpMjdr
zxlrYxsWBXhemjcPweoNHMtgk0rsa3YiWXtolim0/SlC3IqXlGNnyb0zlLhlA8zq
Hvzjd26V6Lpydau5QfYBhwkeRtIvd0goBAepp0dliIXsKrmAg530yE2Jn98I6Jw1
bj82UaIljo2mUaKx6aQx/cua8R1ROIhXxX23qygzOjoIrtYu95CTEabcRlmD97ul
PH4AmtNem9gj5tQBtzp+tXX9+4QYraxzwWbSZ+gm9+IhT2xijmM133C9iJt/JM2O
s4KrZttPYVLtkztkK3KN/RXOodVMkRbjswJjrkEioNe3cfFiNc92WoKRi2F3d+eP
0FrhmUtsPJnFtb/wIXM8mbk4S+gQqx+susxHISx2tvhuDeo2YLLLAa0S0F9EaFUA
f/RPz5sQRl79kwWWoAQO5jPXHNA27DAgIZRmUSYgpatLVuoVpKEKXXTW54b4q346
iQ87bRIccL53QbB3SeE63hLgf/x0TyQ2N3dIMU+5Vknw7BJ6sm8SDjeYD+rrFjtM
5N54pFPDMzLO7FAGsblY/7EQy9bumqPyY1pNW0w6KqMS775LTh79Br3b9nwZyuTo
2jq9+P8zVcYpLnFlKW7aI4orNvK+xNpG+rqJZ1fGTxDrbFOC8ZJ9FfbACd+0V7Yl
pWdigAGSWOkS+uODGz5O3AwnMBJZNQQdvMksWwni5gdJS6DbIEF+Y3paPdH9+Mrr
3GpK+oHm5aO060CPJV/Y202zh6E4osiD1KoWWRLn/3EWFLQBazll7jnCT1gBeASH
DoGAT3k8MeeHE7+3zURQicx28qe35pC3poXSetyWjGI4PrEimkJAzsN9LCp4zzkT
xVWH5Z8b+gSnCbLqlgGVJFiFIb/QKj3edBz68JtPzCNIVpE6/D+r97M92Si0Pe32
QZTk7nGa0LD7hL5SFz9wmip8yeLpLV0h3SZbnvV7ODgihoukHGwbhMTQ9dye+302
BI0lsP7utQhDPm3XAGCEMHeRx5G/0gGSGzR2aeBe2sQ/w/Rhi0YKKxRhvbOxxjkz
GkvZhv2p1Uh9+WrWvkoZvrHI3FlnrCk+IT35be23iil6wtwCNiqwP3ypZzRvh0cl
vQI2ZQe5BuLs2ZwcwlUqloh4SisA32Ry5tGIGfBMLS9rde47dDq7REyDkxJ//1cb
/oMHvXDmVb0WresTqyhizNatpdF1yCWWOYns8vP+r1BwU+xGhJ+KeHnT/qbRQWoG
CB/Sk/j5rRjWIoxLPBfntcvQqTElr6cwsqt9tdwKbvADMk1pcv6xFRHajOQLIV0l
/Tuhe+gCoBogUgoAc4bpIsMogtzUGbluUgKr+rOAvpLIetuMOngLxgob7JCR+5XL
GLqO7ximfU7TDb7oiUcNayDTa7v2ahietl1y7WgKQOwQHN+bl8BiokfNLxQjkMZn
seTfpRtHtHbAaGqOzoKLe5E+Q/1LCRyISCAruILJlWbFpEeGZKv9gNJJkDW9nfcH
ZQADCGRobUaowmgtUYw85RndKBfdWabJB0ZsNWGcCM3+GfMAmnicnGUFsJDpON8a
z7SEJyzbmPGYgAXKWJH+p5cLge7TJeou9KPHhuZX3h46IqsOUJYUMXyNvedfAMr2
3NgEYPUxNItjb8tlEiQQ3j6CHVTSo4LcPTYO/n3d4ok938tiiPwf7aB2z7EpAkGF
9NgsbBHmZCCujb30JTopu7ZHhan5TuP4rOwQ9Zmm1gPGn4aBkUpp26IbyQD/n1QW
EwnexXdCcY1x4Bkg/eGDfQRlsQh/IIAnw1nLkKKjQX/sW8jywnyOQnaYn32hdNNT
T/HWuS4GLiCw+6quC+27M1DQ7OO3GqECPWXr9ABUKCVXUULj6JDTntYrYNHisfpl
JFXD7BxHPyjWXECtt3hzM0JepFOl/P088JQBBS9ZqAzXK5yvBKufKllDmhlnLPig
lMBMDdeQlm6QnZmiRffTfYXFuFoD/8mFW2H86ZAo5oqYVNWszGwX/scAhfv5GAdP
r/94zkFI5NKIS4zERLmC9M5iF5WaTnpUiwIIvmVZQbQEnh/ns0cP8Go12O/SoHkH
2kfBEPbqxFsM12uCeVsiBqjh/upPelBlN1fo69Uk9N9XKQCw88zNg38nPSlMy8xs
gvLRmj7krxF0q/PrJ6L/6JdHp9Z2nbjaIVyq1Uk/nrIYWuRlSxT0csnCf+NbyzTU
gGhlpNCa7VgpKm5EVIw7VrBnGuJSHKQpKJT7JBLiK+jwdRyKkpY/ECORyBbeIusW
aeS1Ih5jOPGZg2sLk/Y9GoVJmR78e2ed7H0MDhVTnbWX3YoySYMf4+tcUpUca8rB
+EldJfkRL109AQClehy5GehPLFWuh4wtb7onu2BTso7s3ao7E/YX7AYuNcSa+Ppg
ToqnNJO8OfsZR5nIMa4qucGMVZhahnJ8X2OQfrp8lUbY0t6mGuV4FO2cTsAmZJJv
hDugMBXq0uITIiKN2DYzzeFhxeFOZ4gqhMEiWGxDlv1gQdDJd5eQ5W6E5Cs/1jvA
nHUYCWwVDKaQWDSJuHEtfgz6cpg+Wu5d9iLqanjK6rjqAcle8G8T4K8QWe3b+rKg
5TZ8SXwhB9vUmxCX2L/VWfBCiEUSw2XkQOT6DxdopHdDdlPKHiLBMVIu1LBlJaHR
KTG3y+fopAiwJlK2+NgvMr4LzxNi8u/zsXNZm82i5nE3TgVFpnFPrkbQ8EUBDk6S
CAlN6wtlEi/Ra01vXJOb2BHQGC+S909vXh0uN7m1RahPkQzBhmjl1oeLcnXvM96L
w9irpnL9oHWyFF+OcEuR4bm8YyyiKKE4flN1TQB6iOkOKr3NQGzRnEZqOgNxBe1y
Pd9FLiy2jwFB7C3oer3FYisDFS+bCQUXz+TjWmuq/wYKeA/10HUjCpKfDO65+dHq
oGueImqjUZH70uf7DzTMYfs8uAuOTbaAtCoHLA4e/PPMY4oePNh6IjlUOdDNzjl0
bp/wez4TsNwsxlvIVFc3Uh7IL3vwQ1MkUUCqyGs4cnqqIdTCpNTaYO6VGYLVjIV0
WJt7fGLUxjikM4mcOV3tVuaXnqW46NGMorlRNINCJYZ40Nz6zo2b5bUZkF/uIkbz
z8LYdd9CNVNz+vU8OfzO0NQmms5UAO+yUPEthS+vW8fp0bF9X/E4jzTKMOj2ui3N
IS4skklJSLQ0ziyVjJBJQxJ7l/oz4C6XRRn2oSqSoobTJUVQryTFpdKhAkIfNXHP
B2YT6C1NR1OBdcMRm94cnEbvZed9Dc3awhn8yAJfaaa9VcaqMZvtfYwZEL38ZLXX
kDirPgsCWduCl+zCA+Kzn0KxfzwVlrb1UUbQIgu16ULOPauAIGgEPa/hp5HcGO6w
novXgI1uCPtJC/wKYrvzuGWna4Ch0bnCM+2lZXZ2zpvV0dGHe/mX26je+N7Ke0Ix
0M4WHfbQ7njI+Qqu6Ftb55FOGeHLSNlwOBI6nWBQJcjGF+uZQaCxy/EqttTqPlmA
PQYS2eK1odag+z4i5C5uOptcFeJrGrRzFInqADVocskUiuCImJ1Q+ggOYUbz5NEN
42aFxN5rXNdoe3LQGlvPiwWCcOgvPOD4gwCVgHg0dnVXa+aDVRKPaGNzuZ2rZUkd
Vm0N8yjv7m1hYAroYmZHJ0YDHlW/aLln1+R4Pb4Rw5yy1FKNHumOXRTI32rdea2L
FZqCvXZHPvIzMpLw8XcHDV02tadYcsUWWNvz/iHYJ1ha81Eg2j+3BWcXVjmOI0j+
DZI83g5aHyBcS0Q0npLiIpV5v/UGOTgs/duJb4v2Z9B6MvA6JLPtj3irK3NmZJQl
ahzAcPORNx3q73r5W/WXpPDHX+FwNi0BIiMNOQ40eRnlQGfJVbHV8cmB2JpBqnp0
IGYZ0kCspdw+7D9tfqRbjH0WcTyCL57diDFFRNadYLD9/TDsfGKcbaP/etwlIqzo
V8/sJoKTWAatFeZK1aOAeUJDie+5LeRp2IxvlH8jJZLVDJTuMAk+3RKoOuCu0OfD
Awx5ZPGltrVOaDiaieZ9UyBmkT/rBuHHI54hyTwMx2etkmqd5Idmyu6EMCvdLFC6
Hx6061hUreC+bW5Xi/PTmhWu/MnR+qPP872dZstne4hQwXSXbDaeGLBC/l+L96mj
7yHHN3M9A8GEkPHYKF9o53hVkIgidazmYiXq9Qt6ovCrrecjfq1z7rQAplUMQ89p
xpVhjrQ8sc1w3T84KVvj+LPHI7jg6zEYaZBIuAjGfQWLbeb+fnHPiETkUDU8Hw5R
c7usbv6YcSk38plbYCIjzgKe6C/9MhmwSuJyf/zxZu53G+LLcYHs60Hdx1/ZquhU
CdS+n0bCzd0pbY4XV4eCbI976lUDimtkObQHmQkGPEcBYHDc0F8N0hSk69PixYku
c9F43KRWzkGxFGvFUtyeUN0JA5cRdR+ZI9JVfo0aZCyQCBnwN0pT7MrIOCfB1lgd
KmWHIzWH32RodOa6KmI5fb+5H1iiExrRa/4Gu5ufEo/rHdDA/V5DceztpcGqY1CY
knkB+iTsy7BrhSJ67vDblv7j8KWtmrL9M0vJt5zVqj+3tO++ArUgTgyCiQBLYH5b
Os0ikLoF/weHf0ECpyHeBxfboCHQhTygYt2VvLR2AU7OrpUIVX/QqlUnxcD4q4P8
AyzH5ZTWZxVC3ZkZorFdQWcMwU5VGfJHwkydC25lKBVl2Y08zdGb+Fk/OuKFZQ/V
oTEg9yovJvm0P9ms5SSfOtnCgijfK6EdDRhTEOCQN9KnSHb10T0eZ2fDqzY3VhBl
qUjccTfIrJjgJMyfxj2IlQ3tTmiwSSsE590wTNkUEm5vfv2gKqWs8noRpMkAmWxa
96J54y5WPdC7esiqCAc1JCRt6HinctH7VIBbvxcVqGv/wBx1AR+NFUjUPczAnBy4
L4MunlC0uPNSK+x5nZeISOApteL/Gu69j/ovza1cnXw8IwzQ2BQIcDIy9CWzSa2/
9kdpjbsMrBLl/cndnwOQHiy9fYE1eLyJa6naGCwQlqiBkQ0jpk7OphNyoFehXlXc
M6rTeLW+NgGjeWGmNpILRBoVncjPekyjrNz79usR80AQYnCkmjv8fWAURNdvDbYA
9Hrp0sh5TGUUn1PamOuUiY+3/GXsSnTudQyTjbZB8+WuJ28qrB0cNpTbCUSi/Egr
oLmHsKpLVAnSzhHRxNhNqPATUdpeNva9d/8eBlOXy8EIqbDLTH8j/cKKCkL/1h9O
om1Km/5YBMm68PbEtcDF0gJov/fqBQnyXCIkde06kuVLunSq/o/1xkak7uY7L4ne
9vuZwRK94t07XqSMl6ocmoHQC5vLNFKi+RzFnmwHdfMeH+PDz+HC2r6q5d2vh14R
cR4ZPY4venLiZ3mzVeS/zJ4vfKzdNYm9dOOEYdU+v7X7jHQJRKOem1bNW/izZL5+
cAN+I9XlKIYNtqXO3+xbNvzP2WjONE0456b1U5R17/DvkohEzoZ46nihCEP2U0P7
oYQHT9agMGRPhKf0icOYy3K6edV8+vqPChqt/Zq3BBlLRQ0ZE20xcjDQg13CtUp0
FhE9gSTYZbrCTroswdRxBk6wR4+bDKTDvo5j5f/A2TRjNhEm4VZeOwGB95pw/bD2
4N53EjSfislD04BfKRRUVNsGVRQD3J2erOfQbcyf5Ur4Lh+YVkHlVFNUXafgAwV7
K81jeYMbipyggeSAHVqsFtVk1SJt+piPW/s9YzjHr+QyX8t2PjZwx5rS2qUDkAyt
UT6rsgsqkURrek1IuxfmYzS5d6Sgkj7QkGf2jifSLW31vtpteqgclNn25KUMkVFf
JhrEKMecKnaNe6whtG4NFkpIAsosXwKgzYJIMnGepN7TaSgRK2v/414jtxMLJw+n
wV7ziaU+zpSECGwCOKqtbtFaMfvsnipv5UeuJXJWB52gNCd1Zpjf6c6pJ+5pXBQ1
+RTwVcVG/xMvlYV1JHVOcht0Mjss7x1lVc50Ba0zyt7y7jrI8XlGb31Vccxv0GoL
MnQ03pxbg6Q3oWLCDk9qUwVrOmY+G4D03uu85Hf+uy6SssnumMnrSLpctg3yDYy9
0bkQaMhXk5sT+x2m2cz121pm6YuG7P40jZqb0VmzRir3iaxRzuaZhw9B9Unq9Cor
pZBH7wJeR5A+2Bo+iEg//owUR4pLa+9gT/ybArO1kLalqZecDoLvPODXJ7F2/fir
4ZGc8jXKRIGZEzlrM1ayQnzBPf0DeBsVL5lcmpGhTavbUWkvY87Xo/0UVrm/WzAG
H0A0v3Z8PexWFaed5pz0TM+k5+rIuoiL6o5+22UfzV+Ynmbj/ZH71h0CzVFj+Wt7
9/AckI3klsbLKCbixAWdwqaOLnHeKx52c4jplf2HV4/sdP4S7+wt8SkeUQsT0SlH
z5eRgAwSBpeTukTu7+xuijYRXr6/+IaXXkg9y0bRT5eLvPkEwR0Mu7GsTjKFNCQQ
WE8TIiABUxSb5QgUgTfKOJVII+nyaF9mwmYwhKvzSuQdvkVL34pJYyT3JELUKHQg
QcS2NJ2oKATmE8TLeb9/I4ilV8tIDj4TnVuJbMLs3GT68XA7fMnAeW4tim/Ov8LW
YJWetfAKWgp7gwqbFPgkAeY8h87tJo/43bpM5b+eEaeknpS1b6Dr1tBXB3pr59Jr
FOr18U4NQG7QicdkyW9V5QxYa5xDwzVE2o5sDm3IpjeGfKdaxwKsvYq+bZQH06tC
6NfpPfd4RaZGV26HOb8W3B2rQtwwcbNB/TYucGkk3jpVInoLc6CpHD6l3GwxdWx1
8VEnbNROfnrQ5g9AsqABd0l1O+Asu0Q5beQzwVgANmVnkIoEqHa3H1Ku+UrFe0hT
WhkoMpyxgES0sZIlVR1EGPZ5USCh1Fny8XuSo9QKHD7n+GVgAU6ggZqXiXZiWIPH
XUrYbAQGTUdXrWxnGkvXr5uKRr28zQP95Pl0RxUD4SnxVijwcI/xie6LcAQ9T7PP
9mQ3E+Agk1f3bK+IihFiVg1B9NtbujW5nuKbWaSm+68qYRo7O1j5rXdCio20nS9c
mO2DSneZbOGEWuInxT9kbnnbjzrtj6nQsiU+qJ8pspGtb2DEGJZHzLZf7jjuU+hA
w9hYCIC12JOsU14SCrIWOp7xPBbh/JDvSFZ1oAp+ncyO7zi3/WUoSWCysQZH3UZW
RGyhLsWMvjadd6QspxRxEtOej4Zci8Pi6gvRXTldpQv9DExKdN5iwSwXkehtJ+ly
qnOQrPzLu8UbKtEKvkmBgaz58kGov6GeZBlAB1OiNbt/rjCqgK415IBKHdTZo0Y/
h7SYsa9krhSiWM6QKjWwezNDG3hjdC09/jdh2rXLKfEqJofnjDFoeSwsgcP321tt
s/mHK1UQ1xzAuMOeOZQtvLVQjIT4fuMBq1S+Oe6/lyFRl1oMyyFqz2Il1xdZhVvX
jFlsZB/QtxeWAZZFqWY95Qjs0mgRYcXmesc+z09StlXpdSyyTEI0oztvkLB784/D
WP+pXPufThlNML94yCV0RZ/bOxZk2p+IOwjBJ+/lJPXXAexf3/aWq68WGQPN43dx
fmODBV4QB0ZdmJCIYxlCIGx+Q2BuB+gQl/Qk9Z2dOAsbejLXPFmbaSrFnVlKi1Qf
iYSKFmgrkNc350JCUnyLLitsl7vv+XurUH1J3s4f3b4EDA7ZG94WukuiirNGEwgU
vECCkhAhZsq8phTk+LRLWvewyRVb2GECCw2s5RZc6sErCVNdNyJjkshWFDap0+xQ
2Yh3cnwEsaXFdkOOxJdrGbZs/fR0dmZ/2q3pWMMPY4vcz/3AIrD6V4Smg+nbXub1
4F2pTU4WYhSb69iEpNRKZh6o7qGaAJ2LznRnO5X2ncVrgSHSALUie863e7wyPCY3
vf56N5Q6GKVaRV+EilUN7Bq7x2WVctlEHq66CN7FQNB1bdumlfBSXEKs9P5ZORgf
GKuKFsHB+6bk0HhiBfeRlzdMFEpExCVhMIm+ldU7soRjU+1FDZ1SlIBFSivxCjcV
oBjQ0v8Mb/8sFXqCbU/5UEqbiBGzkne5VmaLBLtvhwQalCJh/FEMWK9gsrTFdNZY
y3Q2Z/QOjLPqBc6gd90JmS0pk/8swmwcQ/rbID/3w0PAsBS8+oxZlBe0stdFmVcT
NikN3I3wGc7QcIUwLg2K9yj0IfGwQpz4D0rcsd8F8Bl+sSN0BvWHo4fhskdIyD9i
8s+Z/Ca4QH8YQhWtceJAgY05K97//3NTwgzLXVWWpIlF3oDmhTPGPG2bNQSKvB+9
GegI3sQZGstHid91eu+ZQfulbQr29QXZK1lP0uHDVhspQISaAG09i2VqcyXEd9aD
mB7g1RoA8xyam5BLx/GBc6DXbpN2RCb5hmImH8VVVm/yIBlNC9ZgSiFiGTqAgWQg
r0CApo5tZ/BVHNdUY3rhtuEQyE9EBnMo6FfsbTxteRaVL+OnTTwBtG8V76h9Z8WO
Ae9kpOZ0wfAPKsACEla5J+UJRqw2aSOcfywYvaPGFGBtHya7b8Ri3JOt8Q7IOZDx
BA5iNqS4xaadDzApu2Px7wzxeyRM42QfXN6X5SMmUzOgEYI7rSnK0wQpSlV1n3iv
4Jdf/747+JEB19rZmYZsbo0ydOVYFN6LJhlt3cAPPv6NEmxgZlkVH24M9n5BXJRB
xQSbnRvxVtACsBc42/IWzmQ8k5nXXM0T7S5TSnwlyGtNM2zeibh6p9wpwgMpSOeV
trn8Ld3QntQ82+vPO92l333+QjPf8skmQuXutAZ1CQa6WmxVDg84ko+4iFVUz89N
SIkiwSosZ5WYJLV02qTJv9ZVT8cACKzqfAU/D0gvqThKuapRIgny9LFCJsgbesfv
0xB+EPWYk7Dkm0R6lOq0RDGBNiiRr/2+zReW1QPv6+R8bobXNJZNSWfp0J1N9tkQ
8ReBzzoF42slYX0Ko+7jPjZkRVdCCLtR/Dm9aUA7qV6Cmp7pabekngxjFQ4H0j8L
um6280KOb8ELeqYkiHYHHM9jGiZld425eLp/lSBOBEHHKIeVr7exWhh2fW19BSG0
kW8aJi64fJA/hxa7g/INHmbPzojL/wKLmAP966jnK9dRhwgUp4XcGCc23K3unius
+gYh6NnWnL73z3AnlLsh53p+a1NEF/DmU4wma1MAymZwbacM94po5F361e8QXd5+
hhD3/6TyJlaOZmGoKBjajT9peoxjh/rFfr1IMj1oktPQOLJo900+43Fj+07tkHw8
2qB6nXgHHBQdr/Hj/8DomK7YpKSrdbuqCQ8wu/iTA16fvy77aYdqraFdqK5pNL0S
fvKRRlLgoCJzJkq24pcRZmwZRzTJPR9zoAjly/bqUrvt9SRfVQ80WtA7Zp4/uapY
3Br/30IwGt1mQUK7M66W3pqFPXY/EzBEx4zCCGYPCoSrdx0g4u/pHgAhIWhOiLMX
sBVdOjsuPNeQ4/y8K3cLcQc9jkZWltJFo6rm2VrISz6xsdmi1dfr4G8YLKF8hQY+
s8YJLY6wbiOUBK46PbxxYUnYrbkd24zGy6IIxYpmuxdJzefFQYv4sJF6bgJSjkGJ
rbr9n+3pcdrqb5Gc/Ggipwq7O/T1hkYaANEZRZ/EOPPWPXvNqsgshvzfcNNN0nNo
S7WjG0A77vsvt3uQgZd2NtKPGPluGnoPmHz6e1ilA8S/M97MEosquzxWJgqbIe42
DJQbHsiEnoMQjBMZ1FUrIx6FD1oup/rTgZeQvBQcUVxlx2qMi7sDaSWhwqPKAFj3
iaZ/WKzAc64rofkpZw3HStu6diZU43F88VacAqSzEG76X/rkSZCk/iajk2MhQ00+
/NQVgJIowbhfJ3wo07qdv64cIqaHzdZBa66mlG89FEAtOTr2zBLOTiV/HvScTpEd
lCqHFc34s67YlPfKaHAPQC1TDi1CsI4sWpOl1a9H84G0hd/zkukTOn8M/FEwzA8V
v8ecmHDOO1meRJ9yHzitykM0lwM+n7Fam/cC3io58DsfeuFkHNqxSTMsfFLKAZm4
7Bfgs08LHxpFgE3yWR4aDa8zK8OpkjLp7h+k5x7mI581ijYqKV8Cz5okVqeikRDo
X1tfvksy+r7amiTr6uTgtaHMEY7/wJuIKQ/jBDRRY3MI0iPrQt2l+HR/V/2oPxqK
bvaiNhp/SIdcbh/hdIo5CqY5RhMt5zwDglvk11kvc2yFgaB0dNaCbm7z4XP+TbzX
KfUcHaPsFDtUhMRtTRB+OspWqYR+IRrIc56QfqDXqBa8OF0PjmjTr7gFLkzDgvge
G8FIy02H17bjhkmeqkG1eKOg9a2/KxfKaxFu0aosstBYNo2bGBdq5cft1wGLU+4G
ChwcOfE6Ultb49L4NiLshp5UDBCN5ngql2tf0jYInQPKbQromfWJBDXK8tmsMfSw
T4yqPg4SbOjEzmyVVEq+r5rZb86VsSPxYMiVGdA9ZqDcF5bWOeJz4UPv0aKFe1Yg
/n9MCvwEOHs3IOO8AyFN7w7+HbkdXqNDyUh7lOrLvFLoI2AHOr/a0U4Nf+QMEQCO
VLfvn7+vl5+YA1povQ1GUKbmb8ScSZcSdgD4yxuIt8rETmkQMWroF2GHP2PmuvIZ
W3f8xnF8T3BbKPUsIErjGsiR/SpMuTMsrixm7JN0xRbEi8XLkLmUdcJqkuDPbqid
YPL4uuGzBHfGCq0IJsZ0RJQ7Y7ou8SzNury1tddOLINJl8SFMrf+sdrxbt/BNqDC
XlzG2AWn2q6l8apupBf1V7ITNLpYz6+sTEG3oZbDKxRMBm4+jyegj7Tkh1L0JmN8
N+tS74ZAVuBgANb2OOogiB/Tqg+cgrozfWqf0a/zLxakq1m1JrZrvQLFPWE/tuAN
QWD4U2t5D2n5qEvKDgJdv1XzTpqkNRh1dKo6vgrxzXbXSBCu9jDcc+pCvHCoRYRK
SJGZgOfN4ToMZVez2o1NLZ7f+bM6Z1JMpN3R5bXlYH8UarMq84rFPznLwbwccmRu
lKnkJbJNuieok0jheAHaEybcT8ZdzhNTt/Wn/shJGAlu6fZQIehPBdTgJi9rG6Tj
N/Vqab5pcJd4Ag4KZ4XAlOtkcPR99BzH4fYLGz4L+Bui7ZLXfccFJxUtV1XTYk4Q
FVTlYjCY/8dMgsPiP7GfdDfYk05KymzZ6RqaNgM7R/N6zvtyUjzzGPL/FxWJHNlT
6r7p1MPP4R0+AejF8UnQqjH4kHocIGcW43NDKyxRh9fecF2DDKpD7L8WYR4YSkIQ
8kYBL3F/0tZBvjSpu6rK5BkPcb9dF3hALUtO+5nZy764nWDsJ3s1bXZ1TARiJOvE
/T+KqveIeUnClgv5s7xFfyolJ/+UWn/eXushMUhOCz2PmhaH0ZqXNpGprBsNug5T
Us54y5n144yMYWktCMLWsaNXhk/j3pPqlF7zJ6i2SAjXyg7qsMdPla68ioBILSEX
XZC13cPOTBWlRCXMfjddEGzAi4cCGyXP2dD1q26Lq4WiAAzjVAs+YtFcXw46T1RJ
fp9FEIgDQ11ZY65MNJYxIIn/mYcOeKTgBx8puZjQwakuGGo5X2YOmcDDuvJN/3+l
t9MRpUAq7vT5RhkMXUl9S59hV9WwQzso1spvNA8TvXWBV+C7GnlSKra3LCMVIt2C
oTiVx1vggyK/zJ+YtFkURc/zEQcxYvYyXcFBaInFhJEPkxVWTdV+NjLqHYpPRoPw
qShtbNp7Kaxzv43rhX1z1Fza5dby4n2U1/ntRboVRX4E9uzjZlc3Tw7LfNjYokA+
v+QtUofG5VjwK280uBzlmvp8PriX8QICif42bonfAX4/tvYq5cy1m3LnqT7FZI1W
QBrnI55gLrZGwH7UEC4QV5hp/VMJ2Ax5LLwAm0NP+WA3GrJfG3RoGkXkmpYSzDX/
SpilkvV75jnniyUvY5Z4pddvEdWsYhwml0812GOMx9DzrHVnhxnR+bMxC/bIel71
oASU4um3yk4HyPiLiY+hV9/dwmlujnPpugG/Zc9Cnh8I7xoY1z4os9B9rTcmmCUd
PzJQgdX9bCIb28whA18IP+U/BFi4Gh58qZgd8u9a+NFvCBagYMwklyHpw52BZ+wa
z8Stq/j13TGig/PR0Ck5khtWUoA0+pq4lmaDpOzBcFbHI9kUj2ECXq9AHjOA+cau
ZyKxznUKnnzoArL7LIvrK1JHEmwxe991GJbC12Z8Y0REP8HN+DKurxyxK4HNDZe3
jjFBWnuHwim116EJFTVlSJeXCnyqZXFG7Ckca5Q7EUCLaaxD9gvp/pFb9v42CbgN
1XybpmpXcAgrGaIUK61jyTJTKoOwQDB9uXfROpZRSo6DkrRuELF2BTFFborTUGUP
1uM4BPKpHTvG2ZIflQcLgZN1OasZ6KxmVPhJL3pMT/IncC/HnlSZ4p3QNWqJBQ/s
2rgqRE+HJUauusOO995XQBj7twW4q8H3S48UiH0KQ15fspTfrKNBY1Nt68aS4AxF
JnX7l+YGnR5507hMH9NIclH524VfAwrh1aoPervMkAdhKIsUP0bdhuTBQGk5jNTr
BNfUz5X2LKXn3E+ZsWxK1wk2nPQ1aGHm+a3Ddcgg+fce0QXkbty2GhVfmQb5RP8k
1iqKRyhEhpFTswalNfayoaPx9KGx9tlB5zhtEXajVUlCdaaRBBkb4VmEmbPhku5S
++7Y4fYWyGJRSPUmOLxxxRa4eMDO6+NaEGap9oDzYfZ9ODSBanO6ULA60HBJfIf5
QThJdrEe0K2W0qxZl2GDsrZGn4ht9qvS1/P2jng/Ymzhqjou6ZbrIfDzxJjnI7Ol
v1lSCqTcQWs1Tugh4Pc9s7Rtml8Z27ZQ2vLkC5luKljFFzwX6j4Z0ARxdZcdrUv6
ZLbrYW6M0ksZ0KXuT/7Us2Lil6ES/LEiAghnEF1yfkTOaOe7xSVbGma5iIt6rDWD
U1KF0NUqaKQG9RXT3m8fKfhZwBIQVDANY40xwBUzqeM+NQaYrE7GvXpas3kw2ih+
qOZO569t7YimqJS0baHZOAsHYmOqRsmpTyGqGqjVMdloF01GFhN5B58oWBrv5b6K
/uz5DbEFs4+BoTLwqUxGlcY8ZXqGZ5EkEeWSeLZl5YsrcozBFtLJ0THmUvamPcz7
Kk3Sjw0cR+ENZk6snLsYAbIwH0JqkAu73ehTyyohzBIl1s9bddtI/EbDBPdGeBlt
AXj5ozUb91rAeWweBQpN2fF5fkraUiTfMlEjdloaapYBSc1/IerqwfQiYCqJ649o
GDhPzjV/o5ejNtSbzDvw8fFLlF19fhOerrBxKSVi1bClPuhgub9eRalrw2mH4nah
y/qmxsze3w02mtpyWWBFc9URUifLzLgl0eAS0F+TdwgQ38TToJWWCJ3assy+DI1y
6gDoF62YzLV1DFdh34fwIwWjr1qutZ+52hziI92CDt7L6JwrtfbuHhGTkoiNEEq3
uHvbcSKpsmGp2T4HYiGqMCDMTVsKfiucb1XyU2L7+lt8ZJzkTRaCMmPHXrbqWtVX
YsV8AFwGhE3SY/tqQx3HdDjIr06Lmq/OC7f2SdbpunDKrQD7jV6Oj7gfApQHIxDH
jCfAnLzTriGou3tw1IZiiVw1ytHmaX9v43m109BhpTAWJToNiw2EFywAHLMQ238h
5HQvXYkJCjhoNqKbBnXMTQG+vSLTkYQd5MmkuHeGMPra4DmKFjEGE86aDcdaWzUH
+jIyW996/ttRevNqoMIUVUY6UtH+y0kDdDWNpk2O5+fbspxU8aJ52b5vlkQvAFVb
Y5tthIyoxK0UfMsiwmYIhvE73QpdlOgDgYQodmezEx9Us4WWhx8xyQ/Pz/Q3zc2/
BBPSO1nlfB0v/UyNaCpNh+Q+jAnY5h9eHeazkZh8mhCHnW5pr1S/AklixdUs0j18
7M0F4XzLDlShVZxJBbh3ZUSsXX+C9wsJgosD4aNK1sD0E8SbxJJDeH+IOZshkxLU
meujoA3U5OT6DETnLmQW201+WoMhyE9K56rxwrq/GsO8191DnSpozFWt7ajD57sW
LcKYfRsX4Mbr0Jk52FHuUlyyBJgU1tQabe890eHp7wfdl0FuYV+m4quheGtKTQgr
l5RlAaD89ZmZPzhlcthGLbFvPTZmiynDCZ1IC6t6kC/xFfDyDg3K4G5eLw9DaHnp
m4Wvz+9ki2l7f7qNHeH09M2R83AJ+Xlk0MEDx0XWn6WQwRlt5xR07cXqdOk5FBVz
PoIBdR6MF5hwL3SXcJNYVv7z3wDtmPDX6gsGUGDkjY3KY7s8Ym2frXQjBIsH3Wy9
TFIJDHwhYtkqORMtoREWhzcTI4qN+sjvYr2xSJaEYIk4/5dLRawD1umhuKKctr6C
E9/TbqAds8xiDh7OSEYfnyutZksqWLL9JrlcGPAR8ht3xh1MYGNhSpecCws7fcEa
OoD9VmV3bYZXbK1j9Cd+Fp+gKv6BBwFoJHWM4hhACHtM/LNEYegRsx681Jz8IUDo
iIbNUsot+JNqZOqKcQgQ6vUA0xdnbKP9nEP+wV5U5sk2WyUX2fSLSySJQ315zjl5
H7PyxLM2xIYo/JcEekMuzISGedcpz3zJ5TVjA2SW/8b2CFPJqrd4xxi6VUXC9tGB
lmJmMjTAKAscuSNMvF7gtX+xMlyMMAbigAEtx3MU6vFhwi7Bmhvng5SN/4KGBvq3
76aOI8ufJavxjsNivuGml01fBJqzUwCPE+ZlVlu1c4iNXSyreJoKWiLG+Agzh2vL
fi0gErjWYcr+YK4RkfiME7CDtpcWWdtN9wjz0ozSjiliKQSfHpq3jHkAh0IrI53C
DrPmAjAwcfZElWJAVHr7FDeKFNGe1QCTFdew4J/jb0VsVNxhvjMdL0woZ3o1jSWS
jx+9gF7HXbWoqAdmYnXprP0RP0wpf3FucFennyAh4iPUJm96EVEmNoLJ+BYFCgGh
BPy5zqt8G5zoTzFQ2FIhJbV0ZdtbHNb+PtxdueDZAtcKLiJmNlHRUK8kAe9DPlfX
3jbP1/rolrmYYti6b3EOR+E2eKKHZse+IZl05qfzXhaLXfYrXhhovqJhQnW2BlYE
zpnIuG2orNMlx2FViNYy0mIhtXwdo3v2fjiJnJIy5DlksJZnnW/cSU1mliNlj50f
aGDX26Bk758c/ciwcdwZX9t8/sDZ6zrvDSgtYOef4FZ4dGEWQEgm6nwHjienIZJA
k/sV5BZTyPqW7tCFrMiFnwAFpMdh00jybZBJh5jHNO2+h1vvHN6HCqqXc8Yx/78T
m5GC/62PLVqpf/9vc0DmpUDwKYkgS5X5r0yVKJsGXc3pCbjpp90MrlfinwwNcrTa
QX6WWoIooUEnOpMY8ts661Qt5YXJCKOD+b3G6oj0svQQUl020BjgwPSg4XQELpvu
XCFWStSjjmjNgZa8J08Ybbo4DFZ0R55SDEkxhhA/gVqls0ZqwI1HualN7DICHJDP
opYWWBPIVCvFHdQoP7/tQkWtiGPWNbilzPro9wCWprwuFXnvkOK9qCPLECQwHk74
UJOP7l5EsbBYwOJEjdo6E1B4R68hxqRbKv1zQhRNkznCLL85aiSbvRE5u7Iu1k25
+vS3O5xLMc9MKwjIIqxMZPR3EjJ3BjcoIfwDDad/6t0Tmmta2i3j7BFjrKEq3ecU
K3daK0IjVZd4HXw/cMvgsjcpOfBzS5/hHPOaNbV7nuDd/gS2Q/kUXbV6vwvZy6kM
mltZBFYrtPn1/fPuMpElWMNV3SYKHz5bV7Z6x7TKaU0dbixWJquRd31bOb3cKZmp
5+4efMEupWiHPayHudFFpqAI97TL6hdfFu2ktv7rMbmEbonY40h2/dzFfVp+0+HV
bV89Ftf3LC5aE+n5gvl8RwVmICM1MDQb0KhmxGbqH59/zDRFQPaMJHPLz/GiJmcE
g+mSqUVOxso+/J88wfb4WtZ9XuF8MjvD6WL7doVlz/wiq2SPxlIxDsnMLN7+SVwC
JRfQT6k4KdaggLcBU0lNN8EYSrgah6Z4Yi7UlNSfYMg2iY/5gS2/Y8Zmr+ioL6Ej
gMhe3KycWj9BP7EkagoUDzCWfoTCKKX7kobvAM+HHS/7MQtLGOUh3anYJ36/yEb2
72ywJVA0+B3VpNIyac4068dL3lN6Y/aYzLG/U9UdOoUu1Rq1vIVPBlWknsf8LR2p
pUTaZ7LLR8yeC4tt5FAcuoRfAhaqyGp1yhRVzUGw/wGncPcpICc+XqU/Ze/G6ko0
kuwDKyxHY5x/Bg7YLPIMuEx2mtqrv54LjBi2ZeV7K4RF2/vDRwDMuBHUH8EeEMXA
ydWslDA6GjpkZj317FrBpiSHOdpUvGvmMgU5J/F2DG79GbVOijL/vmOTo7t976xA
Q1aIKo3S1wE+0+OnBr7uadU1A454NB+1TP1r7IMukwWDjZlnh+0nE+0FHU0vugLL
Wl9RG8MWG3d+Eb1314KshIUl+vzHxIMheNyped42KWS3oJf5Z3EterA9XEhFaP/F
WRvCeyRSYAxZp13y+xzIIst8g4PK3TXuSKz1EzjkajWl7pe88NgtHKg1LcELuOnG
CLYtTfE1+atJLkTyS6SvxeSDQIGw6bzuwyq31leIKem1t41VGmwSkQsGW8Cuwok6
xsDrIROcXf/sO4R4omDpyOG6I1tuZydedshQdEqP9Oiq32zz/8/t7yi73FBb7Oss
WRHFs8i3jC/hFCM5fC3TwauIGju1K8ERYBlF0kINbIi84C4mk5o5T1cEKOLTlfBP
NQHqahObpYZ7dZpA5Ot6lClkcps2Lkb3twMEQl3/DCVQn00cE4v94DxeE8kXpRmZ
cZaqnfLLrFmHfnThBEu0oRXJjW266ZUO93uflYJUPRo6QXBmyTahhrfmEIw1vLSQ
AkEATr/AqeA9phrfZzrDiByXPQHaaplJj0aeTp4xLB3mjk/OA2A4kAlWAeLi8I/Y
+sKl3Wyk3nGxMf+Ex/QwQ3J4WPvuDJyRsjlgFPspuuJrCtUeRz1J4YJ9upyYD8wy
dAgaA+Y8qwBP1nUaT63QXn+gD0UFl4sWAX7owlfgKsoR0ViNilxzDJOfLsovTB9j
fPjFV40qjXN/MI9xwbwcOr+ldds8MloHkoe8v6UsX/pChE/2MBXv7BVlRfUGu+lH
ikNO5+2PewWHp/9vOOcQiwy3hY5Ctp/QrUdhkteDyH6iaxuQFeWqQSQ6Ylquz4fW
8RWJB+CCVDUYZuyBxX4H/C4qmuXkzEiXMvu/Hg3iUO4VhXa0REfTU8jNv4Vmc9l2
Fcu0MaVqT2QYZfS+ftA3ZTkaXjmOJ67fMwaOkB2ICjmEdgu6LO5kEeyW00hk3Iib
BBm3VmQT2LhsuCJ5G93WolFgnppbFqh9Uu+j2dm3Ps+QwIhyinfwsiB7R9vLKIda
BHmSZTiY9zEb+716M6PVtixWiwagHTB/viywsJWYCDFotbNzVg5AMbNK/S4fkFDg
Bb/g/b6J6zP/b5n+7SX8YgiDrCd03PDisxH7siOl7qlnh11ip/YwRGcKIFX9tv8m
SRQ94uE1arK7fWGvJ7MBfAiHxIbVKzSzXoCuUABqYx3EpbZuph3ZuVnJYHvnFTj1
OJb7t2PrCBI/qUUQw3v/GTVfoR2EDodY/5SSfWzbVFgAAihaN1BW+Z/LwmPrDlgN
qXV6iAHcOwdNpt39rh9iWR6Gh4dEUNJq83/TFnHnmNL7fj9X9UyhpX2DcRZMMwPW
Drc0nmZKNnfKrOaOrXLEacgC8UKFfNR5+dJiqwRub2oR9lknxWpdrOEeLPNksz7p
x/+7bbSETcKJhdrWKRNs+ZS35znlG2+C+qQXt3b2CH/mksrVW3YCwywfPvX+WSHN
DgjGJmofGvFCa/GDvnuXBKemo0Pf2ikXWlz8jgBTv7poH2UboE8FQLDbg2mTIVyk
LpuTpFxiDCKStj/dB1K0lx8Yf4B8KzikW8nd1bmDAvP91NqpR6hdNwxNUGqoz79k
bjfJLIG0AOXBWJp+wakFDuxkbqL+X18+m0WaoySNZT50GtnUe3QwMYumdYMknlRA
m83ycWV58Xm77j6s6wRt4PdAigcKH3alLj6xS9Gx0kuHuSzgT/F6Of79Um+xytE9
wJdYLad3xDiZ6YvvDRdzFn1zIyn/3SrzCTDmShzuUmMji+Qa5Oc5gzQg+AkjoLSb
3qAPV19LvXUkmor60lK/qEn1hPW7nDZvVpn8/0hQvPwmyHm0Qz9joLraD/eumOzr
B6Yh9gDhP3sTsvlfKcspFu833hvBcq82YbwVH2IYPKHt2TLetB3EGReupmxA/3dI
v3xJQXwtUof36xhUQqFebHXSCjF3Wh+3WlRqgNfc12FeiwG9FdM7zzvb020iZ59k
gi53Sc0hw362uEWEoC3SfoXbD44wx1ZP5tE4N21Yvn81xMzjuZ2JXWxUGydBjVZ0
NvGn/mbHE7/PFIK5J4m7ZtT5ZkQ+Bxpifm3yuBM4FR4YYAj49xCadUYrSG2lj9pp
XOuVa2Wt7ijCpwSsRyz5sGSYEC9QeLApV0U74sb3jtwifdFJxt5x57AiodQNGj58
hpha67gwkjDOpuQqjIOHHAlW2szO8MMGhcABXB2E+eMUe1tq+QgSWur7i1Gmx2Ke
Gmo/mrINpTRPbflueERKTnK4qe/Aau/Oic3eMLjGjMu9PygwcxrgFkE87stooKwm
RL7Jt1qPzMoVdJqzWA9lOtzjr2t0TuMfcZbgTVmAWwn5vsmc5BQ+G0KhPfJNOOQz
v/sBIenHkFS+oxk4lnWU+KYU6Ywyy6Ac/GSWlOYMpvozIltG5YdUH8wrYGmFaHqu
2Eu7KPCVW5gVJlsO1nlLAkeHhr1ZjHZVE2YgZQXvm0VIQQXN4KIRpsDkWlCAjAjj
XyPODMo9VsxdoTPexJDLYOVFyOAEQQOKdtSmnHAyNR1ByDfMErdicmUgE3Yn7Y8k
6csWM8de6JAmBuTJBZZl/+YXW509jQhOPQovt/JHc5Nu/SUv3Jg3Tr+25sqBOS7F
zF+S/BVz+Rj0eV9wSi5dfjcpeLhSL18AJlSxDgaVbEUSZx+Hf71a3tEx9GRXaTbb
w5wRgqsSuYw+JfMQbPQhhuaODjj3vdoOf6dNxYWRHl8SH3AOFPVilyGWkLCb6eNl
wyyFAOg4j3DjW2TCVf/hSyOSPdU5n0rge8KpnALSNAolE3huW4v+XLOayq5gTkSA
o0Tmp8MB70ukv+BRd1AzkXaRk6T1g0KBtyY82XQyWkiFyn1ej5CsYFz0BJBFLRnZ
+lmF6dVYZST2rG/8dAwISvRX4quu6o0yfyFxrbOjG2VxT2DVhjWzKHJlLto3YN1K
DJQlXz7VkMXcrMI6JYZ/Ck/wPtj/0hhfLd0Qw+BJnmv2s+JUru2NOdi/3XG1gc6D
Y8xj91JXWpneMs2Oenmk9BeVUoktypO5fz72Xed7w/oMx/AtUAj5x0t89RIFzsA8
qfy8gAPr3XZ+JKM8DIqFM5PRWPlVunYLmuSqDNyBCA1kUbk5QXii/WkBBp0yGM5M
fG5aBxo5McBzExzJA34dml5cjSi4/gecB07jOByVkI1VilO708wKjRYx25KTTGU8
b0Y1mHqF108VJx6WWRru0ZP+SLgzPIF8Z+8FojsDjSO8xNrERbNmYYz3eKNQvI3H
Vyx1KJN/bihIYOGBvZnDeKHSCRJni52X1bLezYYPb5dN+6eteyc02HLoUvAEQT6K
XbevUB66Do7ojygUjvPMbfCgzIET+y7oUdJY0750j1A/F+ZxhykcvoF2CRni4dMv
VMmZmSSQBHaDSCOU89n129tc7Klm2867iKMUvA/8Mon5d5k70U7gtzfMHYUgylyT
DViQS0O++t23uIRcOJMiLMXN+34LrU1BBc0+ygvXrK9vV0R7BUV2stYBlFF1Ro1S
wHXtL0akGP068BEionPElP0yeTc1wm1vu3Ebw6B0VIWFcRVm1fSStQCKIttLD8FR
cuokZuHl4SFdRMm6spM7QNknj9ZOqpPXg/vgxB8Gz89VfGZFRYALQKL2sN+Tpmt/
PZUcdJz3ijkeXR9wN3lsxFoxfgHm+dKp+kNkVu5gEMQgYLSldf0b59GMLbkiLggE
lJqnaeIKgfim/8Rn/Aq3f2QBDybqDnJwSprmn7ciUss9yszF6pUn1JeMLorFWncY
qFr3vuIQ7+OdefZ6+UsaJnUsYVgaO8KLmnlSEHs9bdVLPr1tAZkLHYkT8FnW16C0
mTFe7RNr3TZoHasZdggEC7OF7IrePz8hXez7x1xu9GYYSfNqYoTxC62eRe1hc3wG
iJFIEzLu+riipw9R5kgjsp2jVYtGHeGJOHVDUOeU1XIuYO6HT70nNEMoqqbnY0bf
vukc+GOcQyNco/twqsZ+I+k/h2ueueDOJIcLFdBFhr5jsHUAX99YvUwSMi0iAZAf
mIOyQb3dnjE7M8GrLnyqR7s639k3JYRJJm4faqiGhxDCgINig22MpjbrdRhD4LAL
7yo512Ck/IeYY2dgkPztjRol157NF35zxXAf7B7tEmKRKpVsvJnQ/cinbr5/QAp7
6ZSwgqKLdXG706osj6xyE3x+YMuWXxPk4mMrYXPzWqA2PzvT6OoFMpP8iX+PGVKd
wgHVVytmnXPYxQDeG024wqTpgSJMZ14PD31/bRECWYeAplM0Y8T3hxYaL9EuA5pX
N1fQDZ4hsI0WSJUu8EvHpaEcNLa5vLJKgotso08z6r0Wi21bEdSjdqjX78jyZUQw
iPwjw3ZhSt2EWOChV9yLM0e8hEr724/B/pJ+lAWJ+cRiXfDAnx3gyWYUz42RdXap
PUw4VBbsVFvvkbqssa2oDthAK3rK5XEH+EPqqc2ngkH6D98rOVnurGwqhDLTpwNB
9kQtvjIXmZOYKYflZ6qLUKzlcLWAoXTfQoK/MgR6thEjLUzknA4i3xWmoRDbDogR
J+1mYTODtvdFMf+BXObRWzz1dKie7rYPqn84oSKTC6cQSh3h0gLOhEJeSP2m5loY
v6sMN2y9nOWV5IPa8OdaXGGeNJOy/9UgYgWv4SfZTlc+cWVIf0hRQdIj+gTKrmSK
kAiTCgcwaV1xy3JjV7ef2yN2h0PrzazY28LlnMv0U+UHim06jkn6wq0GLDHHUHuM
Yt0w5avkKnp+D/vYfQnUx6YdcShNinpWxfr9ykJhtkANUvE9B0mFrrZXbjYZKb3m
k18lJI98Bb1HUCefqESwlB1ggqEexAVmZO0o/77a/FQQ2lXFTXjlGgJ7lFCI9BYB
j/CJFP5TuFCGCN3Pw4aXXV42IBV/G4PpKpTki03pyh1NLnwsp82jXqVvGgclUe+B
Msa+5hB8fJg/bol44QDlpemHJHFIwY4KwpGDczew5baRrnUofgggz6Whq3jIFC/Y
gIUlva7cQOpwcmcTnnYMJo7bF4lkhwrxpIuR7rcmOmW1UrdOW5NrzUA3xTohbi8i
kBHOj43ULFV6P+1ZZ+Avd92ZI/S0DOJfB/m0Ddsctqh9IlQfbDA0Oqs5i11r6/V2
t33BQsrrwnnUo1fFiOXcRSP6TSRMPMBI315U2eKHpGg0mAGEg0DlBqYMex8cHZxU
wXdS7Jp+cvJoYTGtqZbG7i1BuajfO9SbMsieznwMVOnpdNfgwdpmp6HdLq2xJo+Z
zlZYFMaK5yBBatySoOc7BrOZKIBT6wbaSk2vY3EqJxgZkbw4DQPWB1cnMSr4eAfc
AFTs5V/xPpLdodepj3yya73jk/G7SouBX30zmgCCCNYuUnDvKImSM3BT7rDBfSWV
l/Cy8DnYBmz4aYf2SshqqQm6epYcflaoYvkP6hufDqJh2EfAYehrYwp88DtLO4rb
QayYi4/xrhnh+ORM2kdYRMqBi/M53pBScNhGIsBHO6Iexk7cIRq0w6v763DmRq2Y
6qHKMXNCL9jjEFdrfNsbw7HmRbT5gYLgMtXhOUVVhNLGog1e7A3vUhcZHpRC0q5L
qWlNGEFmZZrdewnA2BiH8oH880F3AeEf2b6JyRgjJC9gUP1OM6bpHBKoyGcGWTwj
5e3Wt0MytcuZ9GZg/IKLp6VjZrkrR/uVDcBq7vJrpAG2ks6USmQgjWCM333tuGLJ
8Xidf6jmpI75L9jL5L+h4W2inWvK3GCOJQNG4QJaGhiPGJ777kxz3vc8d/4zte/d
sTFAgu0RvsBidmDupSbo9OjtUUdodkUuw412GmQF+7Y92L2scbASvqxuXGJrjtV3
6THGz6ASTt2NfoaNlrzQL0SDtVCtssMiMZC2ilbbMCns0EsitxjcukHpjb+L3bSE
FHNz7hgqHQ7yxX/1jBegDdXyHzZ+8FULljWfJooqGCVw9UGCuw+pLBLTKYh2rbhq
KSlKEyI4DLnC5ynsMO61VlNDBhhiYr/Zihkd0mNMu7r6otreOWAFb7I1/u+YrVrm
oHsZQTuzfyetj3ayPUco27qvKSIcJaBFwiqkqJRRsS7iNKpK1qEKci2rot6JmKho
SOLzEjO5Lq4vfGow2qgHMkF7lJRFuyapsQKy4lbMY0laEQMDputrkvVeIIMWolIB
3uMjThGrpDbOcJKSIQd4sOmMhaBOZt5rNUKzkjAhbAzilGIjKQBp8LeUVdyYJ+71
Tyn1JyGK04h3WELIq5Nyi0HmStELUuCKlLtNHEnxH10Tyndo5mN2o4Soihsy/i+m
gMCRrNBeUO0eIo5tAeOzC/+hjn7uaJBEWMgTZfzk/A90ZBn5ch1rv90qiffTuhpt
gSW7BVfP6PoZBbcLJvVcNnbJXdJJMw8ivRMeaTN/LuYP6ctM/QoXDaE7drIzIhaP
7vnxmHNI8KA4HiArJKVAKkbLVuuQ46kb9GMwTwz4aPk+nahhTUg34kt7Y7nuiJMn
DJ9p+6DBsXsKXQyuVFWtJ1f2VeW47Kw8MkpIauDRzs3dCaJpRsPeKQ0uC4+7cuQA
24VTDBB4Sm04kEJQSBsySsOZD5nwCuy8P4CiF5+KljcxZGCoOLfsZ9AUYptPgWVU
E3KGf91CMqjlI/GCSqVf7NTJxSPZcMEkSsq8sZY4YJ36/4WPOqmwBAEx5CvtNJrS
2aVGuHbK/kYcWh1qXJNgPa45OES8WwjHIPJj4qoaJ+E0J4PhgXgg6lGKsqIp1QR8
0zTHoGijS9lgcj06BOWtACxQLa8ME3ALWj17Yqbw0u19yU0nvglYOzDY7BJXVabf
PkJYQpnkgubWwR0jB11PFGpiw4KtMJa+JvaeFRob+vWSz2hfRjl4hOmnlrfxxa+a
M2yJGk+mate/sCn7D1n2Mt2ItQLO68YzjhJeOIILOTIn2oVQkj0cLDFdSXFMy0/Y
mRjIeiQmu9Q/SmmnhtU3ZW37GyhFgFuIfsbbXD1Dxld2bqjSY6JOFDmtR88pt66z
PTqrLUIZhtcYnnNEgRvzOiKhEKCG3VnWS6lSjU+jKtO2PCJfGplCasYRTRA00VKj
yC3N/hlseZc9cu4znuNvOVOLBbRFbz+KKGY9XVnXiNzPBn3U6ANjXpPOOWha+aRI
d103DnR+bnHoxFmzL2GUeWx2nyS3HQ8TEBdlOAK8DGo8b5nZQ+bJNaZFU3kqWbbU
qMQ3+M2Ka7NA7gQj3kNe0e3km/zZg5S+p5/5IH/AHrzG6gwXK6AD98I73YfGybYw
WGdGGRQ+w4eyQEvEbaNuMsjagSDHdc8HTcp8pTV4GMTJun3z1XuoSUmDfrlBx7Ku
ED/mNXAeJlQUY4b8ijKPrVRHU/WFupwPtTSUQydDnvKWi95ELjsH7OH77zFSw3Mi
g1+ulu52cIWbOpPfLgUAkPdVgjWFBKEETn2Kqu0RofTcW1IJW4U/lJlrIYAWZ5rN
GLzrM+AdslAJPiQb0qGBKBwQZbltYp+Yg4x7u0E8FcXKQUM8qpTW0fPVxgYMSSRL
LIwWKpty+X2QCwGoZuCoAkbsx9ovSMDN9OBaQOAzud8q1gfENS5m04SdpyhRVdeR
8l2qgSAEN8JJAj1kqPYQYvn621bOp5/V7eywgd6nQjkoEXEwAufwF/vtNCZA5EK+
gQtGF+kzs7knOrl2m0ovpBQHcG+qKVtK98I26uOxJpXbc+y5Ajq5wUpIeBg4vAYJ
Y+omVkGJkT4rOGevZvLOSCU16BhjalBJk4QjuOiKyxOCEwCezuJIVipfdDeKsD2r
Uni5S8KWIjUjmx/P+QEv8Pko7Js63SivzwXzxLPT9JUORY5QA2xMulVxzplDipEd
HxmZLlefjX4oIkpQQ7ACKfFib5QNfoRCXbcXz3/JE/ClWqNGWAQlV676zJXEmdSf
fRODLgHYrX7yZY4jh6eiVr9Lf9/n3+998nqtW+Bn/LteL1jaCdfQFM54BVmh6bFm
FlsRGSLk2K8cHVvUbz/nDkpuWNrwvFWZ6E9dmbyNxIi39Ku6elR9RDOQzCpYVjNr
XNSxlFC9k4/gEX9V1fjQ4FqbaUJkmuNhuI4xtLFL7qOrHAD3luNljxZZbc+IiSD5
VlTGGW/2g2khuqPVufnxQ0Y8h6CqzL6jicYUe6jMtax1a4OtDErjYqXlk41Krmrk
/DA7X8Kv5p0j9CiH9lZJFW+kgKkQJzEIh1e05rYu74/AyyP/SG/jL7IiAvWhzB6C
7yHJoCB2jRzHE1gQDVh/TD6f8RKomvkTgLlQ0a3E4XHdF0vJ0G5Ct4fjNEp7wida
fxoChI/UJKK+6VkgB7tk5cSGTim9YvxoygbU9ZJjnoKv8GBUmME3oK7vvOElj4xP
I4hcnn6LM5ic/iKhpb6OsreVz38dXHU8IEJqomttpD0rO5WqNI3GrvytFaTwvS7z
9DhS616eDa69esvRWsyV72KVbQPRAHrGH3p02GUHmb66SajmxUUaBLPVaD5NryOe
`protect END_PROTECTED