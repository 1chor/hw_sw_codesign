-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
E9Avc5m41HlTUclEYKf+q34GR0G0ZzPnvE5gmG4ZKjdaDHsj2c2cTQcK23xpTbyE
bwSO3VV8sSdnkTkZaJyJw47aDo2U0jHQkKqCHEcXrM8pBddpLG3IvsQ1mSd784cD
Ep/8M63gBit5HsUJvvn/XQ5MDK8io/+uPeKoUpRFVEY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 14240)
`protect data_block
3oQDZpHoepScC6D8pelQyqUlFKd7GUE5zsQT+2fIRiA185Md0zA8QL5agkzpHMHY
XysMGcN35yqmCSTYTzl+msMqsOjhPvIsHG1wuk5V/f5EvwCOhmahUJjgI46GQT6H
g39VxN40MPPbP/PQ6Lj7+10UduyLdO0bDZPVocO4gy6GQc8WUDqzSr0DnMN6oQtb
SexkI52J/UH4zVHDS80gjpdofjqUd4GC8upjtAptzW4ScFcAoyuOCDGfeSW9uTL8
CRV6sJ09WfuuOa/9KOrBr2QZXhspphih26lijsxFqV6s+Jw39xymBeBofi3QBAU8
GacFCarnKLJ1fMzmh1MD2CoO1GxdZp4u+qx49j9ivIix44DLYfHgnsz/Q5r8uP+G
7v4RyFIzkC9LPo9bh8AllaJXENUYQwkoCh9ppF5u+jfG8Nf5fuFUyYIwbpxquijJ
xZQxoK4SxIhrRBzIEV8OK8JhwdcjeeOwU4QaJEs2KI2yFt4Xjc8NAb/J/PnEoKcc
GwhJaxDuTCBmwbPtigR8KmwnkMBHnW5IcG+OI9s08Gh2PHlwfZHcMLqX7BNNps65
hfZqB8ovR8PDp6yQwroI+l5TYuxYhoymsvPNubikztF4wL0MeWpeH7VTb7tZ/sRp
AyU18OBbhdGuKrL3VBBzRVyGpo/00806PwDO1DL1QhSHVRfpVGMoXS+X/U100nMu
CXoNmCCZbnU68pJQLPP2pOA95/ZAdLAC+8+sEW6NQNO4sJCLWKod9pSXgrZD5cHP
moMy8SXdrK9Mi6Rm5kkDYX268TFyYhmMn74AO5pq3MO+niQmvFL8bhjbTcbk93CR
zwASGihU2gTlxdkCNLYzP39eEddT5D9UBuwjxStes9+uMAKd/0ydVIC898W0RonQ
/Yv4GYSOQIiyAIqHLwqY5nLIFotMqG2FjJSyIzFURz06chcDZQfeB/nuem5xhV7L
0eWVLRKNkFJRpyuAruGxMKd97bAictrgGN5S+QtvB6dIimRpvEhAU/T2vmBBV9VC
hW82b1Y3ghiSox1ToxzyxCcnWw5LuK+4/7U+z4jQhtVXZ7MCtkgyoyvIaEdGra9o
OuvC2OLZ/neOkdRCZ0bFDSkekBznvcslDlX4/nynydQYN+r2e7rEu64WXHSc9ZAw
qWzWIAFmjP3WgdTno3kcflv+5BPdR6Sp6vUlCgZO91V2Sdh+HCZUmfXmn3a3GYNQ
khqLHZz1OPU8j+6nkP007v8CSqsdHyFuTJSoffjCrHwDKMHvQiJgSPgZAogmin+h
+n8NEZ2/CmPDlwljecKjLfCSof0ETpz9TtoFTj5OhpZzubGZzDszoGQNFf1Me22n
Ec90b0Jn68s2VpMlgZjoaiumSZ+HlVsxTXAER+RUyKhexlWQEcO8kcOcTIrXoIHn
X1BPj/BvUldLve9eODdiSEMhTlcu89wSW0KBIjQzXf9/bDb2Ve0gaQ2GmeNLLsPN
uKPTiWlQCGQPfgXX0O533VhX76NHA9Pn0ZoZQ+xS1zOUarpFtWOkywPlly2KuFEy
eQhH1t6ndmCZ3yKXhFK3D5KXeJG3/LDRHfWDYer/yP2GjiMYQ6lb6QHx3EpXY+Kv
p6bSYZgjrNE1biP2JlMnLBHUhSblTHF52jYzC5+ni7/H3wmNwM/OCd2a1HQ6dq8z
QkRt6kLOP4ag2VMo22uHBaumvR7Zu7ZMq0nt/YWO0yCq2XdiVaLv12iRFFVeyhQm
Wu2EMEWjdQXlNzLyesSJdyzeIGppmJOEfjP7z0QN8fr7joKaLMxFlcWU9ZGhoziF
oyIfVDNLUZYFyT4SMPo77qX6VbUJVY6lux4XW+xvyNVztt395EAGZfOKrHCsSvZP
usbmgpZ5+7AtLO+D2MZ/FJkYOnecRNePYyXf4ZyML5FGcOLuS2wyfXjaV/lLzds2
v3pLhNz8NdBlEAtToIe0fvQL9xIcHiNvJZh3dcXOxwdBN++lDG68pIS8Z/S/3taL
I5kVshAsPFXYyCNAMs16KSYhOYweI4rsx+lvsAlSY2m8MmNRe3O/YOBwtresYY2f
Hy4KGt13tiwnIeENxIBAcfNjAG/Tuetbv1+4tjW5y4GWHB/xMi3CacnJVAPjzU9t
8gxjrYnMNQp5PIUmA2LwhIgUuzYAxlT/ANsnDSl+JYlM02S6NvqooCBildx7AxVZ
F3G/zfUN9v4/8FCJBBoQFd9iI+PKFYyuWWLb6UgIniTfK4BVZmfoGkfPVpKlcwHL
HBzonsha6cVwAoIrxXOtngO37oO5k8T3ocuoCus56mY8m2HVl1Depf3ROxAiywO3
8r8H64ljEdPwqPE45RqHBp+lKINGpcb3aIdQk8MI9u1BVorUDnSdSSI7XMgB4ZuA
noxWtP6kqePvZBVLJIRip35jDbUHNBtIpDnik8dDNouTNdtk/Iy6CO0NHXJPGEzq
vlzYKs3F/sg83RpXVO9aOgJsWXE6pGbThU4ASopI12iSfdKjcDN11Fyn3aRheZPA
lc3t/KzxmlVuddDXBjvIgemRUvFnVs5bWBTi73xlZXiK3WXl2+J7sOMkOsTJ9tWf
K+wR9u/Me8afMiNF6FIonI7sXtbH+3ThmnobAVTMmP/W6VJVP94i8GVvE7n+8fOn
APs3PwGieV8QeRjdj9fi8p4ZpZsOzO/LvTcL3sfr1+b1L8wcQoFdOeF+mBICeL6G
esIgGSEQqx0zgJpHulI8fiOO+U5ljWxyKow7aVOCNVeRmnrvQ6xmDCKeWJ+SMdGa
8T2y8w6QYIufVAtoQlKbAEFJFu7Gl9UGwglsnui/hf4k/O54uOEkyEWnJhkiN7Dq
SVdMMbdM0xBZNe/qHtiNnTNiAR5FZ4V3137zLqH0bzDCmrK/biLcJBadSgoPy5Tk
WUy7ZGiQiulDcts8iSN8WMbkpiVBC9Q1LJcwS/yvi9LJxxMBNVdj5c+jtm0hk6+M
NLdoMql2mIMq55FkzwlIM1WstccnZ7qYiLPBrlUR5S2udiFtuOX7sD45bWaXIpUs
w3oM3HfjUKquyQwpDW2NpIllrWD/m+uwj081qwOtvCfZItpzp9QilVNQ+kJLERT4
OyzvpOLRyUwhGvHQMCOhoJm1Ab19uuqAlqHJwxv9ydtXFDTz55esiyy8h7uiDsqy
xiSBDRGalrq3SIzVLu+WHWEFPDXgqe0Z42U8PWUobMUtdwxyw8Esfl8KmBPq/Enk
EOmgV4oIE1Jj4PoaySONnAst/U9k6DfsTGEDbJiOjCjjgDlCayBd1KnLZqHDvNxN
BK5dyK7VRvGsmIjDLSn5IwJ3brX00Kluw2/EYfICscXrS9XE7Czwo9zkpDGm6E8l
U6QvL8ei87LAsQCcC8ftFxavmf2PO6jpw+dP+nNtXGVLziDsdEGdWrulBtwxtnAP
ppjMlF+7c/9Ev5C/PxLm8iWngZmxKwUlbNnzWOPVS4hDmJM8310+bHbyelnpFzGa
4fFSUvTzWRfJOieT5TErv+H6wbpaVLTREk2rHL6EXOvzBKV/Fxp6wH3ELEeuZlnv
8oDBJAMaiE5i/dVArWhLbGaoVuEvoEX9ycXDPq0S6kn53AC0gVozw9sInI7KYx2p
8unKLPmrLuL50OgRTMwO7Gv2J6uxg3Lv7BzmU1r2c4v4/icWrDwWAOscdevBbfII
rCI0YAjSd8QxAiRbKVqmskZPXP84J8jOQfvCl2LlNMOq9Yqobgd7R0pnCYXCSpQE
/WdWSfMGD8G5ryGKKrf9vt2Sad7SOvEwxQ+W/aHvoRj6KQtR/sX9VDPfDY6AO/Gh
2Y3JIA0coAdPqG5aRJveegqJIWM/AkOg44Q9aOaNr5foFLutpSWtWLArMyU4hlo9
Gsb23qBybxkiAhJqfzuw8kd+nGNucxxsmE9XqKSwzCkrUOEj9eIh1X1JIkkw82yA
tAB9xQP9MZKXPN0FYDrH7dHVtab5Nh21gtpYx9P3gC5kEkYqKMkVbfQ6PmZvs9ok
s4Vo44LVyujboaAxZNEoCxwevoSDoAn0ziV7QrWfKuDbP0IVEtZJyj0nzTZ+tQ1m
LNkIKspLGPU3iZvdTTD54uyyzLdhz4CfzmaUyXp5upENQqUgP5PFNxqpOgSCrs3X
NZ433HkkXeVO1uevINEBh/mHwN2EtzjuZayq9BDUCeDJhKedPATrtdmxluj1L4MH
TuhVEUOn7BI2ZzTjZFSetVxhFMONm6WqIaIM7jQuKNmCgF49QwWcem0yAXjcSMXk
SdzKE+7TgAfyupHj9l3PD43nHcNo5s8h/7/d6vngyKLl0ecxfPUQqdp67MGifxKL
KE1G6QlXkOXTZtyjsfgmvloHDtJnnM59EdflFx+LhJJL8E3tdhDQR5KcA/vzWlwO
SqwI6jP6NB/VFqb7zdxFkmoWlAaSkyqUJ/GznvwLRMvmLwdn1Fg9NnVKOBB+IvjR
KvyamIuheoBmpAHSJSuBT8p0olZhNCysSQ9AsvQ0AREixPP05/hF+6VZDdWjTFNt
hSlzRbDRoOJOlbLeQeyiOVEQCEjQkvKSom7+nJGQLmWYs2SlWyaykE3mburXnNs6
RQgUHDJexmM+nKKZgigB9JEEUxDE5Vgcf2gF9Oh/eHH14WtVpRhmV5ZztJ135C5X
HNqyqUltNDG+z+S/O96VH5BB+vBkqEan0TnVS5C6dtl1FmsOQWWgC4G4LX4MXyiF
iL++ZiCORAQ0zM101FPbOHzWRqBMFZ8HJ1arYqrUn9hp/+Z2S9w4YHAR80QHglvN
M5acZR6V5aKUvmJTuH5a+ZeJzGniULIKD9cA/X4pF2+T2Ml5Cr12bapK7kazSfm2
7dIP1szt29yBy1MCtwYRiu9Lv9+oxA1uLUDyjFgvXt4jpmYaVcNVXuGrlX59GF2e
lRRUhjTP+bst+0eldSedc1BVydeXSS891mlEGkhtSrntvmJjwzH6WH747b/BRYLK
4jtbeH7vXyiELrGe68P7ICAeU2HhDoQ4X/RaegV4dOhOii3S8DoiLRK2BzA5GOqp
Ef8Lqi9sK2VpiwpgnbjXsJLbcjwWogXiGsyZAiMr3A7+tQprZ67HosKobg9JTHOU
MPyduBCuxxVqcPCRIf72mitDY6SceLZtUmaFb6OxMIjvtxwrYKeqIN1IS1ew6b/y
4nqr4ZPBpSP7dXXKIyOgowjcpaYk3Ltk9RlwUn3uymMYNDj2xTciigFtRTdG9BB/
dtqtPs9zlcE9w96yn2W5snx9z76tp36Z5oU5fsS3FRZ5wm6Q7S0Y23D32gLzBxl1
ndOAFwwEIXyZiJWNnWJHme/nYgFcVxSAA54WNNTCs1fAvMIFK8RhfdVGQU46EPgy
nQaEW9TNgVbTMicVAaBEDzEEV3TSm7MWVpn7dE1RtPwpfP/DM1SC5uKaJZFCqB8u
AvqM3ZZGlGiFJBXjmRVKlHThbU3cGynJ804/z+aQXpiwxQAPtmZQmZDcdI9uqLGk
bSQnhxcPwC2He0X4tVehjTOVopkp4gKOnx4gRuusJtvAuTWrjjTVkqFT12Nu1XLk
uT3OaVbvBuA+4FVr1tacmIqauKUOzDjqdvjyoQY0PioDboRwwviHVCazx8aydBIB
1fY1MVdDTMFILajd6gOIBe0ca+6XPX4/k4gsPvPQ7k2ENgguEtSok/7zPLuNtLVF
k19doOKC7m+WQO85ALPSQEPp9RyO79AOhtU/eUL6K70TxlSPH1S+TwpxSncvd7VD
jFAyXnAkdq/+7weC1Rx6kde56dKIN3nbixcN9fzFsVL1q5qCArmcwfaZpENvc/1z
6cJQwHewv/PKJJptT1b1TtfBdk4f2tNhrHezOfLWoeaYkzapsJokJxQxcXN168zN
Sx13xay1AtKBj4o1WGqg+x7edNcZEL9O8ZePCktB6Q4m3nRecAdxX6D9THtVZxEA
THt1OjAIZoM/ZYoYDaCjgPS59eaifzguKZosiltafQ2DdbpQOzQNY7bUawPMeZKY
PpLY4W/u95LQ6YcY4NfQ0GS20ELRDWBemXfNUSv0WF9u6VS/tFV+ZscyOVIw9h+I
cLTyL740IBqwJWAqNH0o5tOo5pWMHlPisUdynOD5mATiRTM+UsO2KxxR5MAasTHj
bWbMPJDv+ZXgWtaUvGaFib9ZePzxiRSd0440NRVxqoM3vnPkcMOSUew2tznCmAKT
weAu+JDzJlZuPpv+FmcPptAKzP8t0jKKcB78sLlEEO9aNcPVjK/O4LnshlGc2+uj
8OfbK6UPaZCiKoFmorNVyN4e/GZn2D/9YGOJB9mZHMkHqOGMvYNOTeQocvrYQTdo
SvRDt5ez6S8V2vTSw88ihDFRqJQeOcO19A5ScgP0r6WDPugkSEvCHB5W0zEiJqjK
dya4LEbri14uQ9iG8AwvnwB1pxMsivzxK83d0z5BxTTP8X8CD4ZFMcQamW/Nao68
CKpX8HeEzYUpoYSHFLAGnHB409T4zWwtk46eXLgFm3Y0PnEcIvnRxHLx9f96pUTz
kkwmtVayBdZeC2PmC9oUFNuyy1OO5CPr/O/7SX4rEy3sSG7lnT7nhkeASvMXYdJQ
ThZf25ecpOwgJyu5sqaNwJUuYUXI8Df6pP5nFaCfFY3/zjv5/UklbhNS+GuVjp35
D3sBzVVOHT+im1IPMLUic+2GiHVg1PIFYYr71rbhkBHIwHS7Fa9wIKPjyluIYVS0
ebW0fC9ZcwS0Sdg4+pcOv7EJR7cn/C65wH0Cb3YXZcR5RtWzje6j1gGPsny+UuXO
OieMEZ0VoALavtpoSUpJetbcOOJa3ouH2UgVD0dYtsv2LvK/7MARr1WEg3iwsJWD
7wkOBwB+kUhGppHqC2I4JXUwjC+c2Lw0Ep7g2mKPFDnEN/3TKJ+DSE6aYl61C8jQ
usefKO5jObmsEmnCBuOJ0T5CSBxSlK33J2eecJDWlubJ6o+LX7Svlv+IJSCFwgO3
9ITbm34e0HbjYQOspicBwtaVLKRMmzWm73sswEDHkJFXdO+tZxGJRHiQtEW4Xsr8
NwXD4jnGrq8bnBECPyvoBL7bM5fxOOaCAPM5iyUUuZH7fSM3hqq4+f9fJcBN4USz
U9ULGrdIvJMRfaekdQnqwsH1hCRusqi6EtSfQEFat/XkVL3n+7fnXJvzVI4GpByd
I8RW0HNvp7cs1WwtojM9AkrtpOLGQ6/QljCwDz0NKCNKHg/cCZ7Hf8tk9irh4TnT
5OX2qldfzdMZEfYRF7mboO+kxsdOewsafL0ihjVwdU29AnYDV+xJJUJePlkMzENk
Mbm4Hd7qFUvxWq/4l9W1nrMNGyhX5AKKE6Ky1Vu4dfsdgZWu5YFKKh/glWF3EsJn
wiRH0Uilagy9OnIDXYMa7Dpy1W3xU4FPk7yT6BuNZhWkjME6GeNv6Ad/atHwVxWQ
KdeShyRM3wBkaX9pfqe4JQaBVBMq/9zeSi7Y5Pl0GWf5jB7k6pYtgIVLlhG9SbAq
qjwPwcJ3DitDyR2j6lH/JSPd5DfhY962r+l+tZuQd2idOgzb8xYnNlIPgqlmtGsB
ONk9c0RsH24BUK8Or3nZUN8VE0P1cXl3owyJm1uIVoHRPY1MXj5XgJJgTvReoJgL
NpCKL3d5mlXiUVQDuq+YQX/Vw5RdjpddaRfWuoTyV+q8Jt6pbZ/HhIwme3GZsW3Z
p9fSEcazkYKI9BSIfQUWBPrJuBsymDOODwY5JYAFVskeggQrHPoLRaFq2Nmr0+I0
LS1DByrnR3IQuI5LAotzNNJ3ZUADr531zG1VBs9H+Z0m2bcV10Er+7LA8yE8MckU
jK3qwBa83Bg7p+oAGQGmwOoEUSnUCEDAIWFRw3ty67M5Wi3yu4Xr5FywOAOP3/iJ
IlfTuHVQL3yWQ209a0yt9w8i7p4Jm0WbgWNPzBZjF5ULph82X7bBxIFkfclXnVnP
56RDL2IxjB8mywIAePZiGk3a4VXFmKACfHBAZys8rXSGYyGOkD/lvXQViPXnScIc
3IoMQr42ZUs+7gGPlO3wfAsYSN09cHFLWJoNVW/1kw+/iEhp8ur2YAuEfRkLyAsL
n4N6b/h3abHuSd6DQalphlZnLQ+Wlx7x7oiKBe9AOBVLqSMYCEOzYeqfJyUWDMto
rSJWYDZ3oT3v4Sv/TLFS8B8Wh7lzv2S8gZ8o3BK3OdPsYpy+sCqHId6ADw1nvtuq
Kr+7FBRkCZwnz+StC/1zWng4i/Q3zYG7uNOHPARkvvqoe5p9bLFobMdQysZxquXe
lipTZmNIs+s+jJdlvEC2nDCoidBPIh19AiyEyl3VGmfiUmYZLdqheawBJsg4M7fx
LOMldW5hNA65qshFn0sHq0ROhm9Xuv5gaEAmrh+VKW/uY5L831v1wugjmMQPXWkL
BAOnSOR8p0ru1DYzVbLGVoSK+EDS2SfddYWFs+O5tUFJK4CpkWJI6SQ1/e3dotnD
6LmaLvAi4HaWczd9bkijLQTI5Yyxxx/s3UTBLPRRZNqDPzTFF6PLibzo8S1tlKXG
K8n67j+QR5OPoIevZ6w139TbwMyu6+T/17D6K43w7TjxOnhFHhZ64rxNzW8J1aN2
asuR5yirS3C52FAqMvUDYK8nCSvIUD+wTv0Pw3ILnKZWU6TA86uU3KIdGMQc+BeB
Cc/3hA6Z5MzK6SBA0m0YbezhOmcLlzGJlw9PNeHcblkiNPDSWSivRrdciFSKhoL0
ZUhMoN3QDUMdxg+ehR/BobTUedvYgVaP2ahhskHkRFkc7FNpH1WyKGysE5M7qL/u
5psStJhpvKzLCD0xGtqBkvLhgE/vB78+WacVjsnuntUn1pP5gSLlWW6k+ygD4zSH
IPU8f+sYQOcZY4Wsl/BPmstrJjcDncB1aKfCLazNf6NMuTXl4B57tE015Sm9IXM1
/tKmKE/IkCQl7Pk08ewkvXfeIdsbwag5sPMnYRuyp7W986wnwXoI17F3jKAF5ovP
HogOv/edgE+QobPdGqVDXdrqfDRws7AsHTrSQfoY/YFuQG7al6TaBA8wyVIpKy4+
1CeeJo7ukWheEjOnbOKT8yStQgX7zTjUHBZNngcGMjjLUDKzcbjTYHON7S+5XocX
hx+QVW5rkjkuULr5PJvBJxEGtazKr6Z1ILj3WQxlPyph8Xz9pSL59pe/F6olKSLx
6oJjONr93xecLUohw46PBVKQLYJfOuuL4V25r+9clBbR7M37QJt6u1j+3IRUjLR+
OMmNXU/el0z6Z5TgzHrv8sleMosaV6OPyu5ej6LOXrGCbDZzTH+/QRchKubTZaBR
qWBygqwywkWbRa/NfBu5+zgIkRvqLlZGlcsYoORtpxruqRbvt7oScIjGB5B1voJ2
5oI/mMJTvZSMxR0NU3COaMUlawaWo3GmkKbPrYcQusCS3Ha5uKWvXEJiIH8koMQc
0Dg2BXiE4I2ZArDTdNAJiI+tlAiAP6FmI7UfWPaQmDaV67zsKKUKqHYVKe/B1ksH
0Ucf7GNY+ocqeCyDD+Xak6ijMM0j1ZknvWORXETOgnFKz8r0aRkuvP4PiQTCv2ks
ZMBm0dGVcZd6XDF38JcdBgZ2bCyX5xeG+yNM7xIAXCs2PzKKrm9dwsYpkgIFtPAO
uWSCLHui7rNEntYY/H7xuvV2sPH237H0Q5TtzEoGLQxJRcouEEb26o6oaVcD+KKu
1wnyTcGAzG20u4dtYcYY8SV0RBAQfgzAzfu1YhizMb2cp0gahk4dLsGA3Iv1fvX+
xtJekD58TAdZ8MrhnOzeBseK3pGmuPr9lZ8/tBL3lAwJWY6mXMSk46BUn5dCHGOv
VvggCOOapfHvY3pNi55SNCx8XuAziOlvJPv+L8jVtnAtLwvGCr82qENeaziYT2ef
ABzMeUCglyByxqKwfFPNfNfQpAfiF3M81uXOTClmrNYpJ1mKqBMfkH63BWcvQHiq
WZ9buy9fvrleUhnWDC7ExYtMqH6xeZb8HAyt57Ypx4FU2lY9K108KAv16qRRiIzE
k8hbvnCuDWQQrfgXwbjNjEi6sJh+M9jDIu0L/bHYrjF+PpoCKwSFOzvl6i7fx1+X
iMLRawUbr5M/neC79nfffSyXzKsqtTSJuaDz7D8g5y66uya+Jlc8JtAevOAL4YMG
vGrFOxFO3GPg+fI+U0I3VfWBUxScWhYzrmpipw+IfpNezq5wx5V9SFCfZeaeOrVo
9FZrhBxL2HVfA6nXzUqto3oPAtW7Aickl7BfbKg/VKJl7WpiE9MXiI8rqHuL7ohw
+MzK6EcZ3xNJ5PuIp0FEAnENhG4Zh18korjXvfFdyFQwpA+T254jo9Wh7p5jOWuO
Fv3vdeSqzNuJCfq8EYO6PfxIF4ZXyOZN/DBZLe2FA0iGwreEIP/n8TLIm+A0lXlb
BBGsr3VvvsL8+gjXutHiqLKWyDG8GaeSsGCRbqQ2mX5HfpKx03sHjWNdhFFxkHUb
BiO6i0MT1y6m+pkiHhSwUy5fsdgJRgcLrtw8i/+074HI8qu19PxfmVnA7/6YTv4A
3G2oKv+TbOABOVvQiPZlBV1rT6SpQXhHhOJLji1Mk3VUjDrllq0VVpVZlYa5Jy60
7nRptVkdLEQWf0wldZ6om4Z/scVohS3LAOGd7NCwIhIA6viOl6TkT4gRL/18G3q3
LFtZ/9fOiqi5BxB5Ydpds4O+i4T90b8brsxpQh6ywCixguegL9a1WfhYj+Y3gShg
EpCx5zWK97kBFanRDmHxsvxSce1wMwQxriDWx5dcJIB8aK6GvYgbDHqkmgOwaCU0
fwqUPt78Aww2de79cK2DrS28spFQ+8PrE8WnEEVo64dW3HykNJNxW/zJI2GnNwjc
vAqIu0VzZRPhPPTzAQpiMM6+qAzdPNHBhnlicBXIyktnuQUdblYA9+ehKSszNc4E
56/RMlXVZee8WTPM/oPFiPdmQgQGqf9mWBcwbsGHiX3RF/l4XZF/KmUrL9LeJ+EK
tvmDXA0lqU4Ow2ivQojdeaXrZkumio3Kiw2MRjurdchZqElu9BnRL9hJOyJZErNn
z5tLaigPBq44lIdlJMbk5ApBXppsJpDiBGdHp//oseqDN06DptGlfOC/+Ng95xr/
3NloepVBi/nZ6eohQCOqbj7h89e8IL3bTPEasziqZSesHj1c8JtEBxnkPV16Dpph
joXdHe+0b3UwBF8QAOk2DGe2A3+2gP2ZEEkeHmIBvhOqO2zqU6e266AewfzkQ03H
W/pK2641lr1d9H3uqyvcTdTyva3yLU87ymJSKZCl2UK6iAEqyBdmU/hfLhT9NBn4
P7uWabff2sV3QxR8JHHifpa9Y8EnS0535OkVyXhb6VZgcjqXRXfdLyStVl7/Gaan
a7HGtNU1Spi10W+RdtxB63EoTd5CTfVT1z7LDktLFwy/9Od/tXL2jKG5Dn4OmoEI
zji9ftp/I0XwJvLRuv/Wvf2UqyFVGtN/AQD2omNOnEL8anVdWX4MFyOqnx+gc4Zk
0em5cNOvTPF4FGhfWk0W8mE41HlnEjXlMIwLerf+5J3XeRiEVWoIZ0ac0zS7ZpdJ
lzKbE+mFS518kcGyJpWST6aLEREmOvHLqfJHPMv4AN8UCFv6+THq9+S5L11QZzNx
+EqrQmrWmc2w8PQkU6hXPhstVLd2RqIeKXYiy9KqzBqdUBRj7nlE02XpzgtuZ1H+
DAxbT9Oh/FO+IddxSVksaAq/l4w+v+FxNaR12zq3PP8ncDM8ulEOdPuGbFZ7sCsu
fmv85AqClAVbBgjIhE59HWTVcYugsCVBX9fjV3ezDgvRp699mfxEno6G13iEFu00
oHH2JaUTBF+akbxA4BY6vmvyZtLY6jwTtoKU4pu4R7DQXUQeSjm3D3eCiS7yVBfr
lqpY6/WMTsqjdhPatd670XPi2CEIchhwSvFgKvySk74oEpBCTIhOXvbzqjWohX/v
G1gpc+Y1vsy44GKadIeOAJH6MFYdXXAzBR2pC7jIeFae2kVU1TNUh7aSpTAedFlR
TTqJXfGvGojfBU08P5/u3KW7a8zDLCHgWSl0gwOcLiMLEagDPX4AcE8W8pYVq/Ac
C0zwoCYihss9NQw+qWxbrGZS7y4hJEg6zLLKWtgTci+cxdVpf1BwQGyCvZfXSpaE
kr1njJSSRQ7wP2jIk4nwQa2CXcEJEv21yMc/CZyCHe+euJ6Wr8BtFqPlh+MRkqzb
fADjSi4P5lj9aUK9XXevNPMPYO2lqcdhLZXh04kT8f545ctMb7Nw6fhjYAC6z0sO
GTKJXqrsaqLJKJWcWHkV+jqEXpQKVSXHQncUhl5Za77NEHCZNi977rUNqQ6/pQWV
aVLDre5OS6WvP2PDz2gsu1Xh+6aZB7b6187xTPcjpXv5gyw7sNGQu0Ndi8X6qAgy
abzeYBlEs+1XR56Vu08VWfFjAGj/z1TR/uv8rjdWd1hQBkclh3NhbXhT3xIaCSsK
4KCxo4WDUjlQLKW1t/QvHlmaBCPEMlnBVGVnXZjsQxt/cLgkpf+MDkV234OrelET
44sAJ+RJzXaR4sAi+nzKSVfpN/EdVmos7HFaydS96kBhiyFZw0Y5uxjcYsAh7yVK
v2eMLwFeUIlhUb3GaLyiWafVL0aq64klhUYVNd2JyKb6kNh021kte5M31DJ+cydi
VlEExmLNxEHdVEdXCIEsGB7KzrUrs0wwhFl5AU8cdmwo0iDAN8mkFX2Wul46Sb3K
4ldEUkPPRV4RNkb6KsIUm2FiW9jyvED14CSryhBMSBKxkpyvB0x7oGZShbt3H0gk
oZLXv2piwMxFq1t3UzobnFzsoagDo2v39pXxW01kgYquAVkNa/ES3TqMTeOp8TGa
v6dpnKPPpoCbpZ72N7No+hwGAymeuUlQKgI0gDscRP6rysRN0PCUAGZ6AOlnugmq
23qnyx8SSaNkwDyYMJxTsNAQPRGlbWfg6060Pz0pxx6giShTRdGQcHd3ZkI+TWtK
NMgq0lGeYLrc+BlytXj3r3o4p29vQwoHsjX3QNUnR4EEngmL/OoWTSmgF5JzhrCK
I4LytRcTfQmLQcvQ5NWu1tRC9k+bxKld5OE2vAqfpp4rnRmb6b4do+GIbgUs33uX
JTGsSJDgtRR/F86doV1rl4j+OnQhrWLX6Ec3u/vXVRhPCpP5WRVx0X5pl09IvNjv
NYN+xxK27kBaNqbsdEtFF5jdIs4NnT6fsFThaySMBFhfQeKQqdiAAq/eMdcCngZq
zfYdatz/JKhJl2mWdYnpDFKP2kNQPTgcPdHIxz2xk6EnUWjjJZWRhreL/1dKWGTw
icBcYOsxJMHk5fsouxMxAFq8YNWd5fO5WqNygqseXB1EJclS1zm3jq+mnSSZuLu6
JOGfxEmf9V62Z4G+zkdDzSRg9qKgaxLQlqEbWmna6qcWJXAXcd6iSuBvSG/HC/PA
iUNGkDSEHCZgzcH59xXcv7Poia+np1gjj4OulL6rQOW1LUaO1uyLCeTzFIUNX9gk
eL3x+Y88aWS8quEvwtnF9n3vSdaDj4y0ebewy4VivYflzGUGe6efq/FhzZvDSXeZ
SQVp6n3vgxcwx1yrzwQRlwrwbeTAibn68PbhxITkcNFFYcw1yP0N9Fb+TMzwQ8MK
ZDNl4f/XJlVXOTPUGNhNkeNPSNoLPmBmpJYerNa6RyR0/aLmaE9g99vyqdm0iEjl
VTqEJsItsIFOfTd2YCAE3V49mO7GnapBacRrDHGYty6kJlk3mFQriHyapmtS/fBy
iJc6NRFnncojds1wN05k6lLUdSoOAG27UwjxagmfZ8ZCVlJ96p/vvZZh7vaVeeQJ
B2CdUFpZCcduQ2s5vj++NQ918dFX0+/JQdyo5wV1K7pn7GkUrUGhNqPkl2VH8ko3
FhO+iyzMt7G3HGxiyC3/Sqb5gMeCzpA75iHFZLCu2I7e3ZzHuUFAI6mM28eLPbc/
ty9MPU/i0mG2W0BfcKtR0DtW96+3irlioK2k+NuyUDff2o3xZ7vKd+1ejNdMcg/f
0+0sik45oMb5Bt0OM7qVnbuHef/dQaDnawlvdx315Jr6vzer+IIkaCh9thCZfeLB
KYjpQyvWi6VCChYfGs6xufFGbdgTTeNVhIBOjk6pZ1cVwKr3wU2gtoiFzTLBzZU6
U3ZZnyhhrxu8DrlUiDl4egueYVh2hMhHe2iHN9dZvqiSgGrSAiHujPAsAXAmmh3Q
2fwJPQKYahzlBVmYzFiRUiXAStMgNpXvaOdkonxe+BqZ318u2vmUFmyoWwjezXlj
4moevPOdo9f53cmUYykvwVnomQuyw5Z4A0qcKoaf6vGCUY3OKI0PqlgfcfPXDPTx
6PDiEbxnPzWhchIG8HnGHvGBfZEoBSTJfnhL4n09v7KHHl3QWNzErjVrTCzr7P0N
m0cvKLKE2xzil/DnP2prgwCWaVLiHpiigCYAvEO5bsbEBKwcZXwQ4IiXF88uNGUq
nYtzKqgAeBuDbegGyYgTTxt4qV3YeNAigLXpJA42e9etpM+1h83DsYbB7msuJA+P
2xXehCgBcuwH1ngZoNwJLsP8MRbk5FT/HXmsSgUbjYRo1wQZyVuasYP9KqyaB+y1
3PxRN44IExcGpajCWRw1F7JECYJ4ss73RHd5oKatGcdoKomll6puA8vv1KXfi4+6
XlC5yMyyZfBH9H9r9RfhzXUpziX61kddcnX7ejlveWXpiQ16TzYaIE7Feas8yHhB
6817DxS03DQTJ5jQ3Gr15ytgxQP1OqsO4rzPap46gsFEczKT4cuC1m/8vxfb6QtI
h4SarrLTinLePsM3IIsOIi3HpGCej/c9B3RlZiTcVOjHGEKuq0JtLBvNZ65Rtn3W
qzKt0iAnfXC26+SJYyUPG/AEH0+zasgEm3INMO0NknGEhlWLraTu6i3394nxzaMX
i/bWzGquVxDUkqTOpjNkNMrNU8mIIdBwM/JLGlrse9r7RmB8SM4o1RSb2u6eT+F3
qjbCT3IySDi8mPoq2J8jUwQ57mT3Oo70no/bjP/KoWLN1Jdd46KKef1R04t9vfKP
4/Xt9or1X/OBOck7ITDbdn2sg9lx0kl7eURLVZ1oMOmlioZdBh/dy8+04WmaHkl4
i/buRO8TaKVJNQgduQ70nSbcgxPr/NpNlRNjLbo7si8GCqrMh+IPYps88htKLVnn
VkIi3+Fz8xyDeInVpSHBDa8Uu2FOvDOPUvOFSfNF+SfVWJPHXgWVlgyFpJ4XlXZe
A1+oQozc+GyVMWKBKYmgqyrqRLx2GcG9pZsVpnHiweMndlgMM1nPg6/TuQ3h7Bmb
Ah1kd4QqmwkqLhVoSmoCKYMZjQ7RgI30SK4Zfuabqn+pajw7krZxbqmRCe42twUP
9sGDwUrMmTm8oGPsZbvJSCy6Ngrf34K18F3GED1rjC1gZweIPySxuTaTGeqMQm5v
94g3MiY+ANanwxz3OMzK2chzlvhP8Wt6mkhDNWVtzT1kOL8y/wITEcI2g8YiPGA5
lRSIy0Ro2iPFacGgXlrZQNEACOZuj6YYb+Xj7hdmRO0z1l2Eu9RZUxVCM1T9LSR8
cDgxdSWu5M38ka8vUKQALsxJC0mUbIAlJclRTb8yDBgJU4eBsaHWQpzNNi7KxjK8
hpUSaJm+/NxSV6Qi2VOysx8Cwt05arm9iV0pMcYFwx6gtkuRTuY3keflmXTPA3CC
mnTpSBINNPU9CJrmUuzbcab6ont/jHOLt4/4uBiH5DfbmVlOG9kKDVw/0oWF+jxf
Yidb5TeQ04qG9m537eihdz8+QpJJGPIUsfIcL1BGmt3MpA8oAncKdG6WbXC7qTgv
FNJcFaXMLchIiqnE5eACHPxDeV6AdDs+hFe/DtAyPUugpZwhpck0gTeX7/syl62w
zWocoYzE8ZqzkFRwPxLzPkTMgEZwNiIfP7P7zR8EP3E7G7u5CFGH4joCof/f3DnI
FugXpiuDwV7B76CPRIE7C1G+1LOnj+s745WhAh/HepGbZJTr5VEoFkJJ4librmlh
HH+pUPfeIZm3Hv/ternfhZT02pKfHlMXAp3kDZlm/sLL0HvCksLjtX9KGbd1SrRR
84m8hfmLuOFuJu/cAtPOFjXYvfCpMaq7a6fITmxXktkYdjXqCxdrRMiHCO7nNvmK
hEs0aUjyCAa6Q67tHTMLwPyWRlyHgEANes2OMKKwUnsowFDnw/o02zg3y/kbPIJY
RJxxS+YEYswFfyyFu6wpVt3FPDm4NOh8X2hERFDMwll5wh/0XHyc9GsVQs8VTa+A
O5T+3O+OYJEtDk6EIO3jAoJoliKubaOZ2jymu48SAxUlLxCO/vH+TEVbYXZ2OTpj
MkC5IaOsEsdmcIMGrdrAHZkaaQmJTUnZcGjOCzVXR7u8tVhgCF/y6qg4ggmWWpTP
stUfHzeasL2qEMCHKksUDovieSAtP7mzVHiYMtwsmVQDBiDo9/aZt0IwTSnGnXsC
60tq9T4m/SrK++MtsgmPCUi14+GHvsT1vvyfhi79MYE///7lh58PyBfSihtbn5uY
zB4I0VXXTfGrRbZjdy+zgEy+ds+DZPftI55gr1LJTb0Fj3/BUtcddd18SWRex/B0
LpHTfjYhCgTAaaF6BqrhcKPtpFztmAP4TUmmBrJnqEPtOfLZx8xaXU6wAUljlK0w
XPVMz8nsUcMllGtkQA4I5tkr7ei3AmvIP4L/K13QPI1YSsmUN20n0QDkzuqYT5Sd
fmzFw+pPrEuVqwBip9jNl3OpEO+vrToIzz5o4ZmYsgQAbU4hjs1X9ENFtEYhp1Mq
4VzFbg4VgmcWfRYKMveKM1kf+7woliOVl0YlLpA4wc2AHGTI+tZuUv+4RTQulHlc
KEojnRaVByTW2GHsnKKJMr1zuFZ1jaUdWM8BSYUjr1mQlsYFoefLrdaHIuyaAtBR
Dj3iB/Tg0IXazTzEVr+SjrI1kGiVsrQI1virbdBHvW9mSE+toFkBIjGJpyteh0yD
yC6VAMpTnq4vz62OgeIY0G+UAsOQGO7Pc52QAwlm1Wjv0XuTcE2ljX9vABYltjGn
sfM6qNo/sELjrxrQ/I0Y1G/fav8pUUnNVlIUJlSedO6L129JEfB9S/lSmaZLZQmb
tSsBeenjSI2y1EHimrgtTQFXFfV0Inb0F+QEgbF6gCAaGyQVmEjRBQqItH0MkOFJ
Qhcsqfl1FiYr+zPuHzZ79oI6ErzVfj1o6wjDlumaQEypjxORMybXyyIjiYEtDxuo
N4r69BlaZuWxdrsNLlfmesS6prY+Qywj+S3sH/J/ixxlyY8ra5ikBrSY4zsD+pPd
wS8yJqGvTvRmsLee0QCB2boztf3oQu2eAvghY1Q4nbj7V9+fqKeve885Bp6962fy
1Afn12IEoA+xOudUHFFFPncON1HQN/eZUfpfO7Ll2ZmVdmkhWoNImTL+N9IiCVZe
jHIWFsdLRzimW+CuXaT84DDbSDtrizCLRq8Lw1JL0clnov8VMg8vEpXLYUyX6HRd
KRqfQRAsx8O9ggR1T1PL/AxYk7NyHRWSoLC/2Ozn1y3FoL4X2j6w1rRw3IQze7zF
CaEvTRO5PfRQR5ArDSYXL/wSdqOkqy6lUgxlMBIWLhm4E4v2dAmkN3zSqhy0CgO1
kcam8ylqo1uGA7LgQvH2hDsRwxS++68H82IZzPVXERavbqOxhi4qyuVR93aiYPiT
UpoKHW+4UCgTkKDYo92bf26AdNV7NLZ4gx2gIBMj0Yp6MWT7ApKNWJlElkJ4fRdl
cliFIEw6N8eG5M3dfs20y+wS+WgrDSnRcrfeiM3FGJ94dA4GT4Y4icqSG6+DCTmM
svzn0lKbUiLm5vV/Sk0MlsSAcHV2Q7KsKzgDAt18oDbsjgFnwT5TEAZm4SvL5qQf
7xw6EMVas145diax05Fh/Mcu0l8kaFhURY2N+qykEEVslkqoBv8sKfvLAe1VkEcg
hc7XM5+MiCL3QUwlZA/ELps/HECN9Q+Vx/y39qoqCNMkN5sKl6TQ6TMNNnw2eAVN
i/GgBdLnIc2BbYQjSWMM1IWQCN3sFuh7pSOWn+JE4hc8uEzNeylAl+VjcJpRR3YK
P2B6EVyokdkbPsiV8V4CLVJkkdMUQtXz7lhxmzz/EbY+q/okZMM35YGy9MLB+9MS
C3q9FhLAsp7YdGXekDetC9tWMEzKmBsjTXxDhNb+2lFjFzZVjBSL8ULwo8SXlTVD
c2J7oFGaLVnlvQVrc6D60RE2Df+hPGSd2hmm1TG2ovlYxSlP5SdUuREk/9ueu+/y
w8jeB0YK1RNMRPswT/eUyzY1T/SozYeTdlNsi7X5bL+CZMVSgGYn/Mw20OEdDcTt
LtaLgZ8r6v4mi4jloKOsWLO+r6sa2f6opNKUyASZ0+IjMuUR3mADy/UTu5BmoDaw
TwVfOndzsESP/PDFZtJh1YvC9jyJwule//nOVrWqPoMTJj3uaZWu8jtJwFCwuHmM
V2FSYOIgI7Yh+LQNQYN7L+bbMZyZBVvsihzW5SHPMbY+QvRsJu1FmBjeYAhI/Ume
jHZUiSAsA8q8wqxlPpVlVAbsyNj/LqJARfa9o+Z91aOxHWEkduuA79RkXbqAhaa1
TbHQKlFf+5nOetBMtxv7Fm/FXeAKxMt4dHBHxQ9P1bmC8EBMIjs2siOZ7pE+0kib
kOeS4V/V8G5m7QJKDi1pwUKwVXjeHlYTrOQOt5pweN+tHgjl+VuBoxTRJG8Kw1iJ
agNpFgU9JdS2oHrXKNj6J/tFkvUZFBbLUhcAchb9x9SatuDl3AtRVOEDF4LFDYLG
Rkml2Gh83meHHUVh43j4gdYR5kaYik19eD0bRgdxTj92EoXjhgzB+IYvnkGxHvvQ
BMPgPznp2ZCt0/Sf8tboZ6HXoaMPz0XwV7rTLQXMjA7Tnt6I500RxnYEpVovsuaA
bjzJ83h05pTPNrLMjv4/e87tj4uJx9Ql4PsOkokrCLk9sVKHMXGhL7XdRHWDY3lg
rhInynYMHRT0AYjhQn0tI8OX1LDLhVDaANu067WaDrBJRjO7PdxoupuiBt/DdBWd
rf52/418xit/eeZ5OQBOgz7TueL2UHDsmNFBC75xgrwMZNouuZwlduxNL/BBr++z
oKP2G0W5xscygtCZ7M+p1XS1yyARzE4yY1FUi03GNmk=
`protect end_protected
