-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
oRKs3XsQlXbSTsUHQGzm5bosD823ArMcEXMfotxWuYeDRkw3jv5xg+qYOvciHspb
NhGo3DUv2IaE9JFz7EkWsCF6Zrgn/ugu4t1FMDo4xjw9o3NnMBv3tSNloHfLlHPV
t4lSJVgBeg/He0wSTEmbVAEh15oWs8OzVM6j7WhYVc3lYE6og1mnPw==
--pragma protect end_key_block
--pragma protect digest_block
GjjxqV9S43UPfraFSwBCHOZDeg0=
--pragma protect end_digest_block
--pragma protect data_block
tfxTA/Yk0nbivBN2tz+55tpU/wgckrJ8nLjCCVUgCOwUut2zYqppYITmhimOo6Hj
0Bd0CgRMEyRT6/3j7EmPVa+IkatQ4mX5QldASMBGk2ZqkxT7/bR5z46o0foGGPKQ
kRKONuK98QszWTN8bttUKh/KeGucO96DdwRhs3foMJUz8tfwUPJ0ThHXkx+5yVbU
Fp9A+nM216+GCDDVCmxMYdG15z9KR+AxGqfdkSqtj5D1NfShKQJ7QBx/ct82pIWZ
8ujSD+b+lc6wJoHFxnxFK1IPWgwnq938v0l+bm9lIVim1BPq/431J2au+QMDurZX
wVkYFY7uFfz09AFUdWd5caabG8YPZ/fr6QcVDuzHjt0jmapPMfP3BszsVRCRWiOV
2Hmza0hb6+45oJ/F9M30/YweEEaWAXnM1DBtNpGnidbjgdnSYGhtd53cV/q4ODmc
3CJHtk36yP0dU251FTG8E6cqBujVmRvGO3pejlmyTrbZrRT/gvma54rgSCJIdwuV
RSxgfhsaa2APDUMrcqhAuJVNLN1OLggc9BSbR/xwtOmGhrES8w6H/xvBBh8skiGP
tOTwW+2HsfQ55Svcspz5ENle6EeClkGPCMa1WBhzVs71dPxwySV+QdYAWiXqw1K6
IZ/Evi0tcm6zDo6bvSW55mx/6/3QhgjtiF4jdzJqPEc0WTXOuVcoHmge4946Gikc
l5gyNFyr5oyTjyPOmgdq1zghMoY4z/iShAFi9aiwOZM9F/7ROQdIxm1BtwiZuOLI
NXwhjd4BbhHQOdU+eRufx3DLhPk4FIh2TPDcqhoXXzmsWuOtr45Do8tMtl1YXUxk
zVwiPq9j7LLjdRiqE6D25inr5FcdZxZUI6QQXuesZZA4WvCcUSAf5x6gkdF+nOdl
syYXwiaWE7qx2mQjZhjKNi3yck3ChIAnUMa8X1gODyPqIy0dLejMgDn39BLqgvhg
MuAqjBLQS1TP5PAcx7xud8jGt2Yt9SCwuVPHYwtqLpcKc+vnk69J5zjIClB1PbjT
ISqHdG3l5mrRO5iiI5ZjrY+/YxDxhbQtNwu/6IYWjR9MVKGR7wl/z+IxMXSMT/N4
R1gtwFNcrerojFtYx6oo8I4nvpyRvhTGCTQUYfCzcQxqfI7s4jSl50N3W/CQ2QsL
mw4DfdT4kEY+ljzTIxuZdilNKjPNx/POdzvPoz/c09F2SNovKhEBwLOBTExV+2cD
YyBYd1pkCyZYOHDlhvqRuCJ/JZf7BBUBX0dhyn7YEWL3g3YUXTH2JPWLDh/E92e/
r1bh/kdHMV1r7Aa3Bd1JLXfBgFX1xfJ4q2cau4FtNatObEPxpbrgR6rdtWYYNc6w
3Aeduibtft5LldmkiAdyBPMA5dMNO8vlKij4ATseLeU7EmVP/ML5mQrddF3k1rtf
HrITfrpLlYjrcXHxi8O1eWsxX0EOG6XhyGIm0GfhBXtfGO+aqm0RhFuMWbbZx9cB
m3Lma0/fcilKiuYt7FxOsoKhHvcx6/pgFpsSCJwxOVj4mNAQq0/bcCDob6+KvQED
noaS0z6ExN+NRxiZSkqQ/oLn8oWcpZpbGK3J5naQVw1TDUcBXGUeclhJpNLgAk4u
UIIgzmLutzekzp3jdkZeXU/5V55Lc8Z/D8iMFqjQCElHxkPmp3uOcPAMJhxRduIu
Vi5Inh4mo1K4p1JVxYNPEkyDYoQpiOieQZJpHs4dN2qWMtAfLZGfgoH7X6mpoJ9v
gHtUe6LWf/r0ksYjYoHR6wjOJr3BQHny97BuBkl+FRA8H1VnWI6+zVMRmVSQjzbz
NDIiu7dqpPEV86Z1sT3zxoilrQHsxoVFxz637vkOzdztrXSlNF3M+vZWteCpOe08
fp6WYqExL41mxZp828BY+vxUi2vl66fI33O4XZwlqdV3QrBOU8xTk0SObxR0B3qI
Fr2cLWOjoIXtZGq3pfTi8XiKGVxYowL63br54GskwvLZq4mVDW6A13Engtr5Lh0U
dmPjA+hUME2bZpyS5vg+xRSHtktJesGOgZ10z9qxUbNGLHSUIWaaqCRJUVrScJlS
evpO2FqzBDd1cJxFuxDfIG2n3HJme4Hfeb01qCvytJPHQ8UrioU1M8AOR+LMbfUt
SEibaBFXqzRM5wSzDYPVx/6pmUfD4vQh+6fheO+l2/teS4ZhRcMC3PQVV41h1XCE
4SLTtg7Lj68Gsf9vs81Tym276fYlbq7kU0QlHtO4q0MOn5iXxnpk1aIJvD/isNk3
0zmov3mPIiGD81op4MSAipn6t5Bj2eBMwgTrK9QFfUVn2NRqNb50Uj6Duy3OkbBe
ay2eft+mTMzyQpxlfJkq2vT4VNWhF6YQx5WuH7o/8G/x3fJRliCeUZnfytRXYV5H
gh1pL4VJXv7yXKDdc6y708dmMlgw3phI0csT/I5ehJepDu3L3BxFaM74rflfhTuE
tOgfo0IRl9eG/Gx2HuPU6UdY2UnAGJX9RfJP5Wq6AYqhjOE6KG12sq01OmbUTPTG
v4zHJBuEchXOOpeaylyNhNqdSQsVK2HfgASb8A//2MrmAG7+DjHyuCWqsFjcyMgO
Kcyxl6jcNrhjaYVQaEYneMbC5I3Liwql06KT1koqivSQCvZWSMgN7XT23zOhwH5y
y2yMyu4k+Jc7ca8rc9aGN1xw+sR6Ko4Emeo4ZFlTl7u7mPtn4OJgYweKGdWj/zTZ
D+uJLT4SZPz0kNTESoo09eo8afQg+IPh+aALf9w2jMwkxU2B9Yy5DHv1KJDiJuUl
vkJzV843F1PRhHRKk4MLygahKwhDmXTsvZF87aV+PKKktcWeePsAe6IYl6chw6EG
eD6hzrsP8mCjgsfpDtHtjkmEyQbquNMvQiceRwnltZ3+HV8NdlUJoVTb/xvgi3H7
v/zU49+QLOdNlFIkWk9JCrYNMTBhLOhuVgM+JFcUY2m14Y6t2eCcLDOK3My6rL7Q
9OG/NtStG2lehQAoVNoc2toU94Gl7M1thAEPc6Iza7x+3GkdI6YoHmPByBlbDbPF
Lk/kvwO1flQEOgo/ZqiXhPWRVJspSNgt61f4RYxQCZtXW7W7zaD9l+b9groPr2lw
Y3BfJ4FOGC3j6qA55ocGVgZ3OHz8Brs609LCsetpQIktWRHc1p+xf4L3qUK+/Ato
ds9l67BZGnCk4K+Aw/E1vVXcZBq3HGGjtk5OkRHmSVLTrcVBT8LND9kWhNC1yDxu
McHMgyCF6XxIMra9S7nUCilozuicpApAUQ0/z4nGqohv9jJLOXLQ4/0+3tYiq8Js
94ODvQ7vpWYvEA8eroWFB/wZwb9GxYoYUHP/Xl7SBDjH99yCWuqjpLZFJVUepLUm
0I64sPopdMxlPufNTlZl2f6xArhIldHKlKD/ult9jkeMjCwvV5YjEsn+L4YZxhPV
Bvuj4QAYs17Q6r8oejFAOEU7HwFdMBy0Rb81FMj8qtAvASZQXwMSkxtd5cNRK/bH
5LalYnDtsUnuMEPea37PhCWqUy6ZmvM7HmffAa3TgU1X25TLjKDsWLZunPTSxNK9
42b69Z4zLdkcOgpjBYlEPeGvv1lJXr7IBOWzfEHKl2ixf/IScFwUTRSdgCIA6wHj
KHLmLHa4qHnMboW2TrZFJGR6iHZkeGaCJG0qoqYZdj51Ka02CTppPHg4Kw2GIW4Z
QWewfT6Xha8owypocAdSYDq4Ep+9sd9rbaN4QlGAwsTcvFNo7E6sCPVeRg44Y8SR
oBvhH4Va+t8jrQY2CxaimjCl3iwClBASMIKwt253Yh1QSTIdRf/Jd/JpVtqfXakH
YtD6Mz1HUibxmA8+CmHsM5rxCKllrGaPVsn4j22arCuuO/upY5y1iqEo+RvbFEQM
GDVoPEbk4Dbt7ZI99QmDGxywa8FCWuVEb8z+NgX2OhxMg218pt+roN5UFx4Snw4Y
V6BAX749y0Ugty0Bou6ULBRPBQiUbwX6jNPayQuYnPtOIx0V7DnZVyCpEYi0/w0e
KGwnDYSHhTnwXFjvqdqvHYZJjGZZQx3pkW4gOFyvX4gJoFbcsXjyhgjFPsYRFQ/5
fIidMrDlokqtZwDjylvCq++ByWG+vBbTe9mUClwKWEyydf8JRTwy089Zh4KMQjHY
rYxFlRCyFYC09ahRR0scFvXQiWQ7FNoSwWRtfz8Lopk1ZK8c1hc/tpn/ptsNmGeQ
IZFNnRbQWw/JfbtK1lHdM7Dm8D4yAQsdXg4FH8+t0Fnfnf7rA6/mBds+fSi9ezPf
SLU0uWuwPnpEx3XqZMJfiAoiLSfAZ1RuINix5dJvhseds82wlUzcOi+q+fOmkZNq
1UVx+12OEYkfMAKojMY69IbtyXxWCcG/d7N0LzydoJfjS6q1YllYIMjBK78Pd7DT
Z/rnzmiw8gwmMOgAXM7cry+YTb3zIEIvsUlIGgGVBWPWPvoXL3p6LStTeZFhUEch
S5fXUETqKM4ZvBL6HzVmFtfRg2XeFgIrATPEDbavc1XeONJ3+c5O8Bl0pvSHfbNW
GwqvBkX02b8DhyfImtAazdVWTSRTNf6o06fOt8Rq8ZdD9yh0WZFl7t50Qnn0vbh3
yW+U//AW5I+XK/cveEe1Q6Ply5uHhYZEJnYFa4DDYOj4eCcDj82HJudOJyo73GZQ
5lUvsqujRjL5g/UNY+sNmnzekToMUICCtExsdR34g+pKJEpFXocEg+VKaVJyUSES
2YXKDAbgacaYSdRLUj0piFbFogEzpdOUAgliaSN/4Wzv2S5rlsLnDoBNhZc6bs2+
QGLdBP6mpOg42D8VQ68299BneGlXPeOGvumA5Z3BDBdzjk/IthG6GP2W58NA37qp
Jf1ydvmrrDVOlY3tokwkOXizqkAOilviZk47y7AaxIvaihX5iITYMIMxSHeGZ4Gv
6it4qEJBGUz4rU6pWDM8hSBfDLnBmj2b47PyXW7G7C+QHny+vYnPSJ3ALAlV+IT6
suj57S3SNBFi95RntExFHqzLwBUQA6aZ12nXn6BuCc/vRJXccnU9Rg/T0TSxvPb3
Nk7Z5wH36oYOolYXT5KjblAycjnYUEm6YA2/+cfM7Jz2/F3sQG8wJ8VX4GxT8M9u
w4fNJQRk/7ytehC9JDDn11C1DGU+Lmn+oT5JISkBZM1yHHLY5DilSmOz6pN8Rd7L
tE+C/RacvxaESpOBrdazVd3/m6Q1AACEML/48UJJHtpDk/j80ZIGtXvaXwdM0t9c
Uedg+3Xk1afYPBVF8tDSfhsotvLj2EjQz9vZIQ0B3bwadhNd2/Gehv7hiMw/nLBx
KBu/s48Km/fHF5NhObUbR7gJAupbmfEzxOENSjmIqHPahR5fyzFxCrc+6X5NT6Gg
d5VV8zlybTqorVSQO65uqlo8E6J60gChm/V4D0/MwkiiBYextKjzvMi4c28dSWmR
bL0RdFWvgTRA3H6SjGtPQKt7PyXAw8FhKnDdfOBF69GLxRchrT2sI8FD+yCvHE2j
PbucEuQxe9M3GSCvY/rHZotc9Flqc849DYmcpSS/IAETP1WaWXmCZ3eqdr7tSCmh
4SUNjvD0nkP62r93GgZfch355C1mPdjQUFFNYQuha/Cb1RI8+V32hWIZuTgfsSJD
9K+W3cuTVcuMg7MSVGgKzcrerSCL+357ZWcqI5Le0OX3yHCBzUgygwKFwH8LHc6l
j8iajCq2sSTGakodkCpqe2lZC9zSvVrXvA2B1RGhqq+5ML4IQwYbpcBTPuXh6Os5
cYEUGUe83WhtDcIxihyYiJHAWZrIqItxiuaBmG8RNiQDYn97X0Tjxcph4u4bVstH
8gLtPAlvkso8Dh8TAM68K+q2JaN1sZrsGnXERcR6Tgb1n8nfniOEFL8YAafVp4L9
vvLAYzxTFPgpjbqaRKU/EsX8IYMl8THr9+WkWhq1mAiMZRZ3EtVoA09PWQ3nAKIj
C/VnCDn2aIhcyptmmMi3pWnyyr+t1JNmQdMC5XF8CK2SEocBqcU4gvBDhFiHiIFA
l+BpqwX1UrHnhpViaZE0pMrQ+1L5Cnaae2ILxQ+myReqyaBv5QPqtExpTwnyBHod
w+sAT5mLF1xHw+dPKlYKwlHRvBr2V5Qif66rRbnFqf+VcIRbDw7sSkcOLKZrUwrE
I8HvU2noFwhOiroNx9CjfYWj100i7FeZHFOsTZ+A35X+7aMMpWD+Kc6zm8K9Mnnw
ivV+q057s3E1WBB1Culq84fGg+uGAV/q/VQYp5f9YGD6A/kvNU4NJM2h0ivJ3XRw
CDvWeAHsOE94jZCOMxRSYrCFFvNaTKGePIJbk4kt+uqJawTohiNEc1tKPWDwdFkr
dweXsyj8+rBgZtXtD7oWxQKTF+oLtlLPVnt/2rHzR+FpXxZ7t8bN+4gCa1x9999L
YtEZ9FB5QrgKRO6zYVwNThibtdng1OyYUonaeydOZxDy+TRtarK1OtBdSax/Ocav
9vrE9u7AKOIJ0DB/88zG3zV43l+AnWxBtOR5qVWbGI/YozkTFDse9fbv7yddPz4O
6gszRnlYE2om1XxmPfYGfHc1wOX+v6fKbX7wq4dakcqetoZfWyJN2rGxoeC7FXK9
8ifhbSeVbA+F6UzX4cZ9zTFtVde62xrXwQBQdN9cF+0Jy+SPxAv8/phN2f690+/p
RSFEbdJMMFdTj13pe2VMUWXCkefr5E70nAPRaXfXAwnL6cPfkBu16EShMr1fXHyw
RD+71DnkjFORWmDRraTzTI2qEArlFpiReLpVKtW259571dzS6nnBpHsm7iQDBe6U
ZbrRGxSKSNrCCLnT4A7frMVrCG1LO3UHJq/rYT/B2lSebl+Agmgx4fGqGIBMWN5v
aoBW7iHVRy89h8i9vToLphevuz6sjVIU32KNCwT0hxlKlWUXplc491Xl76Nr3dSf
RUFgsoS2n8KPb8sDFrUnARgop9mryC0P/FOFC8GkCkAd8QyHuRflZ0e9X7ezBWEY
0KvqTxkbteeyKxYxmBecu0JjlMwamz6oJ5wm8E/uNZNwU19iFKaWCsH8l5wLLp1J
ROJphS5STie15QCJFxEOLfqnaSEf91gwI1q7xnk4sNgYD6gWTgVRykyze8gcnwv+
dWCQLdrKnyAQ2XKokf+OBlpN2LDiCKx95heqWfnv1Y1OCwBVn05UvPUuX6gweLZA
2dNild25vA1rvmDGC8gKtgdgn3ESwhnB18E9L7IyRRBGNO5sq81PoUM4KlyNLBLw
GWXiS/ypyWrdmH0vTcrN0CGmacCfsXkrdCxY6t96Jc3ZrESeWFL4OEkNGOVMQu8Y
zdIfqmKuGdfdx4n/X9HgdKlNcOjDQ2vVWTi1Wr256LdZW5UXyAJmSwt3tT9U2JQt
fVUKsIpt5kZLP/JwBeIkJHcxNSpmuobXJ3EtX30KMJ3c8p+jMQI8Qu7PH7qZR8wS
1GcvDw04tY8jYDRCXiAWftUmdP/vyCwQ6G5pnU8oXK48keTRbQtAmz7yHf6oY2sB
ONG2tBHCBnr8w4W2Ku+WDSubjwxWN/co+SCDC7CpAriVZi8xleNTSGI+QqM43BPv
BEyT1adroKh1zXMcL5IDl5IcHudpNZvLoTCrzaDSFlslxp8a/KYnESWSaQcGtEea
IY+V8ua6sM3y9rFeb7zmX51BCpLgkcLqm2INpjcPSn+9bRNqEcdczNdTUkugVkv+
ATNYgCLm1eui0OwRumfET9WWJK9+B8EJu9a+Bhg//+7V6GxHPEA5d3BTt+ISO+mV
1vsb3qaH+zDiVtIvSjubxpbLdSuGZDLQPoq5WFDCwnGH4YU80yOM3zgNmhnWJJi9
J8xuOzYpRo8OvpdhcIWUi2K4RHZAsh1d+oWtG4+wTixGuOW5bNUo0L9o3o1tdkO2
erSSD0vzHI18Or8ELj3UGHgUhsTbBDcMGoJfkB4zEKqDldUdgoodtbHokgePADQp
/x6018CLIqPWZ56MCblQ8HjYt/GYdrUpgdmpoopw1s4MceesWptj8i31OSJzgJsF
+u15eQ5ghkDwjBhsZvgfJHg5P9Dg+Mj9qToHcTlF1dy1h+3EzIJgNfeS4DlIHOnw
y5lXelCZBaDhIjHm1DdfwkGOcC98/cQfaWShCLeleobvOa8N2jXlSaAHPmurdrr9
1TiEKEIqRE9jY5n/qfhBmbJ6VtAXpWNYwrgvGyIIueDo3RjJ3zFUg2TO13OZfVPM
n2+lIZu4pYNZ85NUyhQMshQGnxrk6nM2HcUcJnJ1w8aeLn1zjmUwThPCNoG9dGxS
aABm/C63wpjEBV/sFR18GdsK7JoDhPTFGh+pZx6AD7tJv3mvDmGbVgYS+yR60+Vi
Bp68qhiOlf0mIs5Zu2YD5ffxESS08SNGWbbeGE1q2Wd9dtCePa1DYUyK+7TztnPB
dPnyfu0eC6Zy96QdAtfZrdNKQ1mWBHBIoL5YSfn9aimMk2Pj8qJG/OFILOsykiFs
Bx6ZpKa7I9YK/UDeEGsOeN/PKW4HVeVH854sCnoeKVpAwc5U7BMu+jeDFn6Ahcmw
vdfatUvHvWApJu/X7EbxtjfoakBC8fJjsVvmRF6LRPc2Y963obR68gsoxJgPpkw1
pmYkvFB80S5yQrB3HFljtBm5a52f/pi/5Ev8Ww/7QJnety8LjDoTCj3JlM56GXAs
+hjDmP9KkbxyUlEOlNxA5Deg2ELEnYyruyLtSCCDOp6YzrgCMwPpv8KCbryCk2aU
0l1i4hZXXxGiSLaoBK8uYAvwMPoXHPBvRxDusu5ALOo2OE3pDbhEH/uMSHgB0vIr
w+ujziVvEAkD33cFDlnLKXQlPu6ShOr73ZlJsMCjujce460iYMe4njaUfLyG4/GD
4D23s/tZjeL+sRTZwBhupTeW8s3jDarhxqLk/+s6zLLg2QYFMMQTR7eCeLNh9ju7
CXc2f7Vka/BVQJKIyH9tfi+KL8GjIPGqhATkTM2eEX8C1FDepGhgDIt61SK3s6en
RuZdt2c9qihRyA+XuzxVevOn/3lMjp3JdAnsvQmf84NJ3XPEW6dVI3T7QvX6c44q
WWFemnOuXZDCoucYjkUFKAmMy3htM2PtFikk9D1Vs26jxIhbstsF2xs4HYtCi10d
CwvgjQpp1Rig88nFY97Crf9ouj3hkjmJCir7TMzq6E0fr3IWm4sKtlr2us6HhFrX
7bCDUNBEtIFQ9vMoXBCQu2AT1/yMotC/NxfLrHUYzkORp4XKc3ieVHC3jP1uYEaR
SAzBjQm+n7zCrXPf4qdS2k4ZIHP3xw1Qq5d/kQd+jHvE3MVIyLVYPY1zYBSQd8zP
tXa4Ftar0m9NjxFFD3RyNrSyvEJe+g3hPtGtXKndmxnWmZMYc9zs9Lg9SbXSIDvo
2m8C3jT1pdmXSLE5OfIJNZRwOmse6tGcDhN6aOoLS4TzWZuZeWdaekjEh7SWu0mm
Hk7CiNXLiz/wU6U6fxDIYcCTdXaYCczFtWr3GUiviTcDB86sEOZAxnV6l3vLVQrr
cKa/s2LGnh5GAEKFqyiAQ0kYzb8vW2ctXvdslrDNHE6edeQJALr+wDfYlx5uuBkj
OhZta+SpAO+QF8R2tJopkPQMBaEDoDwjqzFUassRJNBwDoo8EcyPMZ0Vwjd1r9gv
3e0xJy1bpYR1f+XXEA60VcJ21U9//VL6JgjTwp37XgCmDn18nOaYKG/7KQcrytjg
ptyl7hudjdqO5N6PhuH8Z1vRWSwx4zEpaHPkKui2ikfgCnLOJyNUn/U5p+JKGcP8
wSXfrdLCvcp7yvmXAYixEWLsDaPdaIbm+WSLNaUPNZMsC3AIqFPpVyKG79Wuob/q
7OP7ir5lmPoZqOq2y3ffXStWqm/t+Q2mktsGd8ErfIUFo3U9oIbTrRAFhOuTHK2W
t10Ldbn2Ib+zoV0t+tbszz4Wk8qlK9I+h2D6yQexz4Qb1ITgwQhT+9a9dBbaDhom
BolwhGl3yy58nT8s8AGm7V1QcxsHwAJjWJRwOY6Bw2IqjwDZ+miGG2e4T86cfvf6
CO+65kV7Cz9L61nOPZHMnoZcI6vI9L2ZJ/5qbJelLohyduKVYcc1mtOUc1XSprIS
z+C9ILvQ+g5u0arcqAI9wvQFx+ZHaj+CUW4f6v2KOZoAzLAZNNgDsWbv+w088VC1
ce4AGQMRT8qIpLJxaCPqeMgWtF9kbyJ7CkRiaX9DRLyeClq4+JFjRIBnGoOeVf6Y
cyewRQTT3MEg1zCoTcXgADjaSqXMA8jn5chrmvOhtzezvgbRCH/ad3ziKHCj5o1W
vZtA9aAO2h46Q3UvzcJKlcL1OHqv0bmmguLyzf2TSbBCKHYwgLO5w78/8YetOJM8
G5qmmIR6AccQ34XUtgZr2HBhfHH3ihvBQARyoG5+Kvm3APBqIhDonjcjIumLg8e6
lTzSEnwX/6vYY2qlFwRzGfK3ZWnN7ZujWoyRiQ4dwHzq09QONGlvMQhkoFUzTa08
rzbiFb8nlywmdVPUP+8qjTx9HnBWcRIOQWUWJyjUN5BmNcV7O/ruYCSeenmkGJ65
gFWnPveLiz831fQOl90goYVG9kWUFPTW9sBGwfEvKecZzf1mvcUnLkgvgOmxNIFc
WwR7yVQB0YUTrNL95E+78hpudMvfVGt8yuvYB/mWAHqfvhmjb457WFOfc0CuJtEM
X5AOWSZnnqxdM7SsyUfJLatbbYn3ZlFH/uR0e5H41Gh/vLihw0p3YkNjRF9M2w75
M+3AplQI5kCtYUVtGOw3ap3r0xdVKSI14XWGd7mXfE1b9Gz/kPgHriN1BPDF8dTS
n/MCn0kxtx2iSNoaYsUoVjYvKj20rwzTMmmxM+WJkhtNA2IaZAsxavgemwySTXfC
Ybqs+clf9m3YI7NMCOqLhbhcOJTHyGvv088XLqahr2IcduD40G2l/8+V3gap6w4E
KP7/bdH/ikbYr50HOGdB3Nj/XFwlLVv15miPvACLGD8blVuvXUeGSJoTsqopCdYr
Qv9vxWlVrTKbk+8EQnAB5Q4FYEx5MWySvp6O5rOma8pd/0uDT5BI9Hj7MSPoJY5V
JFVjATWK3uHLtXURuDe9hkBLZ7zaKtSaOgGKNW8anPOajZ4CW4KRNADdON75qKCt
IE+Xe27rWqHYC7D6cnnaPweL6JemI0iPrLpjxY2UBapqt9FaxoqXtcFJ0CZ+Udy2
gyUnZYJa9Lid1Z+/L8y5eDRAHR/reXo/cRhnSSibXGuPhbWvEy/cLSlXjcGO/Vq9
hNyXp68eKUDGc1KnXdKMVcU2QPJw+f0+V1a2ZN2FE2BXcF7ZAI9qjFEkC3thE17E
ti4gp7jCmkkgbOrF5dcR5Mo5R0ufM71Yp5W/dD3TwwfzDuNXUbWqFge8/P0iG/c8
9ehwvZod0Xs0iaXgjw3yllTkE3tg1Z73LXnTW4o19Pru6Zc4vfvIQjlzJZHpLmLN
8Sa5xZTEnxngYyjICmoceHk9p7yVsqSuTYfkluG0i5X2QJayu41Le3d89XUXaCFY
G+8oR9IZZ5KEpX4G5kgc5QqENGWJDdHs2Mcn5MetEgM1fQIOCt2dKoq5GZJUf7rK
5NROLuA3eg4PFXDahxlP1ZzbBF530bsSt7XC+s7fX+DkBV1ZgVw5Um2uDcWF551O
uvkafRQ39cvP11CMPE1E8F5cuYdC0zKGyRcKIV2tojh88J1PexFz9aM44rgmkvs/
kEu8QX8Yf3lEPjag2qZeeYb/dS4lOjcQGcG39sShmKHla2tQ1b5Q143eDStDHgRq
K/cDoCyor7BFKIhDp1h+2BZfuz7Y22raEED420MfwD7Q65ta0d9I8YISCaIlIyfM
UbGPdfSCRzYBhzCgJvtgTQpJ56ZezBwlAIBR3RrOUtTAJORhWw5vRUbA6eAyCImo
JB+wCCM59U4lt+4nZF0Dn0Nw8HFRdW02x3dVBkSSTHCtgZMyTnmTxV2An9lKpEwY
HIiiDz+9A19pytl81/WzSnfVkE8YOoHHOOJQvhiwDLjNtorJNrBQ3VlQYYyhF1xx
N5XwZoWqOtM0tjoxKfoueFZDbuVDPHbZc9Un2wVdgGK1LAcBxBunp5KDS0cHp3sE
XQVoHQ7AfUBpzyHo75giIiTEGxSw9LrFoUOofwYz8tw/zraQNkHcJuLAgnR28N4B
kBFl8fs40QcdCXIjeo6j/EVxsGFIk89oWjApmpMvVr0uC2hEjPPem8ZLwEQ2VDhh
G6X3SKIOLq8J3x7MeFidDlzC1MIJ6in3qGEaezXDy9B6FTkPXE4qIeAWpeiA3Nuy
Wn7yvf+EeqyOII/LutNAzkWFmth6npQcT0BAAWYMmI4EvlESTfZPmS8qytTfX255
OVSmq3wEV/sCiVNpsxU5dRGc+MY8e5iKZVvqxbFztzouRzxbp1240yGom+L+vqoo
rec4uKk5NRIpA0zIRdc1b20vN9Yu6+JiXxz0QzoWpUTo0yOF7R5BGnr6Xau0/tXC
6nJKrRSAYkmHZWL/j1Vt7loKg/5H9iJApytMTQwsAWRHK6wmR9b6i8C8pHxDR0Bu
3ynEyHGvLoyIVUys8CfZgicphRCbkvdJwGMFPdp6+gSRKzrVkNS7ncmfw/zXXRbY
esTR45RJeQ/uBL9PpiwCYlo5fyECWnwFUvWjzF6ZQx1PO86g+PHxdqlUi3KVuSWz
yoXDmkz08dJXg8QM27CVQduiSJQ1E7GXNMSsNDvepZx86XPU0onSUQK39s9WS0cq
JZo7Wg8n66E4YeYYdCSdbXlUv71aWSFG36S+sxK/3oMwQbr3lbIYUQ4ZlqhFzK3L
jSXBWiiNIt/kKQVe7/+O75mIO1sTK7nnj/wUvh8JI7wo4+KaNq184FION7KQ/VXK
oYKemDCgt6ucn9dLL+23GRO5SFP9SZ2j6a/2PosyBCb2QMlcLbBIIlDjKRurUR9R
27pxI4oRiNTNgR5aW2PiFxjXdC/mNpB2dPKREGDlGevPHV++sE1V4b3ColgxQJuG
UVyzXJKa8jNuIiTrFwPfhRfChnsxA5ZvGQXGw6XAhbwbuhr4D0sJlH59T2XbK23k
bUebbWn/1k2Vvef6tWwNvSjvFkNLTW3djj88MWSGbXJ2FEAvWKQgNnXAVXhpKCZq
wL69+J2viNm20X5QRLBQlbFAzirNkZxfnIo/u0cNVzHVEHE9U2Ou/PJdbJHezOoU
qifwMwvS5RGqQdYvXtfdYMXCuEvRyY0QNALo3hSjyKwgSTW9q7MD+ghy4C1H2vog
qSmlGyzpc7DHfC1C1W3aGPZ5Aq2v6EQjrM9CyMX8D4VMYS20sdoCNs+hOnFdVDYq
d8rjnzhoHsrb6H/TVdlNEVYJQzYQ8mgLWEHnj2CZnToAWP4ccocdbMLlZlr6xxeD
QQkyTRATLPnAaAv8jpDj80PLrAHf2CEd/ceDPxhXJUbam33cIAMZebyuZpY/x1Qn
K7bsPrnG21HsPChJeC3UqzUOPPAyHucqJ0pAGuF2SwUj13/32zWTFeKAGZ53WQtg
7APoNRfOGg6CsBzy8/ItNoZIiz98KNumiJ25wb/e7lMWPbpBIham/Br8sdsFYAFl
nXUBmXKNAQ2jT2J1evPxg+5m1ckIrZ47t0qvgD7C4AbGf61KPm29HXLun/R138N5
eThQ9NV83potXuac/ViiWzTX3G9JATkdxcmYs0pnbZS1fbUblBrpGa3w+XKzKY5V
his+zwMNB1a2lS2HvED6Lo4v878HOeCP0XdP3O//vTccfTy+LpPEEJNwMw8ikpKU
DEcAZaGha4zwQTNeWILiG5OYJ44j0mgFRMXDCJl0FgZXQM3KBVky+KIu+2KG3Ouv
KzCua6SWQEBjK4kcDn2VoJ2aEhGypZetulmkQJAReleoux16sSsSw60Z7P5mU0q6
SvqpW3D1bpVCB23vQNUqTqxMx4cCdS0ePGaSrtodznj2S6k9OzgeoTv1BsZqa9Ck
IPCCrWzuxkA7eV2ke6oldfc3R0NHpkdzt/oAz/+0lHleZi92I6fZl314aBVgEa51
Znakj/nyrksaBTtZsxQqEJnf4J4Y6SYtSkLy1jMgXOD4ZKB4mZ+ajBI0ZIsDG3Ul
/MPUkh25EGoHx3fXyACNm0po8A+SlBe5qcumYWqPCrfVnaPZqggEdMbYWHbX97ty
9a/6gmJDMP+u3j0FoDoLq5qeghTbTkXhRIID9ztP3VDgMKwDPtSeG41cyKouf6Sk
+4+CUOkqsgfJ2J5a2uQtpJh6TA9X1kNqM2NgW7/hP8FYq3RAuejI+HB+gmmUxfae
T8DA4WepNkIcr28vrxWDM0rMXv3yWQrLBZRBtu9Bko/eUwOGfiZeq+4DWAuyyiFb
Gxsdz7uDcjdd5YWxde5DAGPoncyAaptqZjBpmeBX3Tqp/YUI0wkRTpQrVhrzWhZw
y8B4O3OVswibOvVoBvfedU1DxLFHFFHSI/ZZtgZhCrGGwj+2zqgyv51batah9VqH
w2wVV06DICyOXcWsanFQwY4UW+vLETsRT5bMwN8HB04hVvo0+EoQAeSFmyu/Ryy7
pmzlkxdE6YuDuc+oDn6rHgkMrCw3F/Vps1JnvdcL0cNuJisa4WoWJeOCU5SlnsZQ
KxDfzi8GiX7fC6Hb/2HcEeiZBoYveHBrl2Qt6qxa8EJYDjSWyf4vI9ElIOb8KUNT
Qg/ePj9/u5bYEyzh72y61s4qGVb+x0orjfmH+5ZDrvumxjpwr1E+xLK+F/MpOEtu
6MRC7lzgvb8aUUF/w730cVwaOixPGK9ldtCvJrmZWyqF+zJbvQopqumTAZOQuQG4
Cr9K6Zerda0FlMsd80quxDQkoZ+CqtXBv9tj0AVxNCJxWXO0iZUJluPdZ8nT7kLK
ZEpY/33hdrJtresBKX27G7To6oZD37C63qHv0oZPfs+kSEZA7zUgBgak22UvhtdH
uaOOUY2yQVIy/W2hQuBcnDjAlN9Ox+RYShK4f2kFUGoU4TLId+pqLj2akP1/nER6
WZQnR5lSADfazu96WdneplIzAy9km20oNwey5Juh7A3iCeY4uoqTZIaCCcPXwoT/
T9NnT6Qgw1gtQ/NbL+Om1qbJE3E3oNSeY6NyvnmYzmSpAtImEGIW/GkyspAIuFa8
9Sw66A6ta9gGNTqUjX0ExZExQ67SMF6Y2ems6kpcTdtSYdlld97Wk8A3QKGCuGD7
5xUi9hgp3hMVBK9OVoEBjcoa0BmDqukdsO0jQ1kUh3/e7RIiBRy9tGktNlkHy3Kg
1HfagiM7KYC7fCKmIV4JB3U3MSB5b8YXxNmgWCe6BfvKL6/QFj1zSEBH15iC/vQN
Al67u9a2iWveCkrEaJTSQRytS2W/J/6ptKhZsht6hSsXk6DErt0XO5AFfsV3VN80
qjRpz7SSlsrQuc+BddF3Zz8za7f+ZPc7WKwD2faYiB+mhlvofnCcQgosW7/+7+hy
2EbyiRMPIsucZaYZos7x9DbsZfXWqcdFd8g2wnavWemghNwSQuqzxogy0xnPYnLb
jcBrZWSkZJnjQpM9qkvdJpLP3iOOEb1Yj/XT9a7ejj3fRy/SXeQR+VUMooGeUC0B
OkY/CzlfiwBjY7azQlmQwHtUaSGRVMoFxkmr0oYJUQqiqzKuEPfJzclvf1ZIiFjP
Ep0QGLeHA+fMdUL4+t20sHoa//mm1EWIzJYJXY+ZhS7fqUbgVe0w1+ZHjcEP8bWp
rNpBhEAF6kQ2snhdRm0Ez5gHcachRAbi8AF0cet3/U2zTU0xnskTt8hZvF642lvc
HokMqnwR1krW/x9Hq0syXOxhgONlKElNJsEavMAoVm458zLAh+kysP+J3pORjLUq
jv9oGGJ7dP/52QzXB6dXxFhAiTYsYxuRg8khQLvOeEznpmqfuPkKpUYK5Dxon85g
CcXW5sNZ6KlFCmgxWsuKWlu6eCHHglcZ43j7JwlS1ZLJOOpxZmXhfnCQt/Dwr4H5
FKKkGByK1q1AUkR0vR5ZhhlxyFPmdzXG0frAwxnDMR05+DunNu82GrpBzfsiCkbA
4IHK11FJzzAULHh2ODVsP9Zu6oXUJRtCdAs/FdNDzduc3pAKGOpRM8yLiexG3lUt
YTXuKeZh+iPjuEJTqEPxtkxSxRnFRcbggyK+5+Cjfo7FM1uc+bOBBzyNBD32BoCu
QdjXve+6b4qUlkJrthIzG6lbSJBv9jNWxYb5KeyjcDegtwA6dgSccHC25EGovget
ICeFAfgUH9RO9IAMkVXE61DODGUdcQia17SqNTVoyNjwm8XVfWo/lQzRdx4kL5bq
HfUfT+w73iYlcjVIrre3KFoavGHCgm0zK9xKC5PBd9rlPG4QuYykwRlMaolspX74
4iykH4DLZ6/T47/g6fwZhhgzb+8gosE2NK9kFRtBdo36QUMcUVL90KjBGkzSzaa3
EruZjRLMeGpPVsjMEEqBtNzEyNQV3qHCkbZSB4aIxwjNKKWpJVKu0/xin6vRzbGY
eNHnXbCn65JUrdpU9Bv3mt68JzdMnsNi3UWZ0HqAFn31NJRxv9Av6SBCBYAq3KVt
uOHPYeUz1aMaiClcodYbwT527K6qRZu+npYc0w6nT9h/0IBAk21ABvDwlBmxbU54
X8svXJf4nQZfuRywhMRfDmxluaKtCLItvJNy81hcRE5zocdFz7jEn+W2mRjJ+qhb
c13EMXxZ/QEkFlCQHhY/OXpEsfqIepelQs1SHvREOpsNWY4bEYq2JZPG7oNohqlj
SRwRJKxQ1JmrQaoTUqDT29MRR9ymm4oH2xlT2nK1Bj1ulfM+DcuPIDlYbK+TNvWk
8zV3cDpW422XNciJDrs95zfxf2MsZCRxk8R+Oplxu686xYaaAGi6t4z9i45N5LpJ
nYr3DQ9ZGYlmplDzcoaKKt1cs35/GR1dOwmq9ivDzOEbW2/mgEUZiIHYWKruaVvb
STVIridDMXuoM2G25Hr31JNrkvkXiEk5B30Z0lxU5rL4+VMhPQaMK9/v1T0ZofEx
0zrvDyQgfr4NR5+PdcUMpaRGi6yy5o0YVtYniHnpfyugMqCq8Zohuni1plDMX+Uz
ylHLFtkqBt4XnbxmRIgJgwnyg/iCWPWid1T4HDQehLIEPDgQF+PfdbJpPuzLpXR7
uWHQRz0785ZNQa0u2f2StstWpb4f09FePB7B7AgK4knXrEjHJL5Q0ZRrYBV8j8Ar
6NQEyEBLH/4yblYs1QBDEnvNFmkh1b1GPn4/CWD4TY6L8M1oPfqGGGmmYhyp2hcd
+l2XgM/Wfrp9tzC5kz+aAM2bFMqTBBJ3NqmbgpsD5ocUpi60U8Yf7pMMAzuTR/k8
8IzcW5ABHvcFVDHCpt6YNZSJDEETiEiCmPysa+v8UsKctkIxv2keLOWun52wL/r+
kqvmgOs0cXgKlurEWNXZp5L4aWf1u9nmXWENsofCRIvuMy2bieM7L8tvKhYoYJgk
g8WkwIC8Ua2Vj66lSB8Bt0esVGp0PmSICaQ7ifdkpRldBcUb0TsZB1OydxtSXrrZ
vyPCb0RBtH5vR1gUsJdadBBRpy0vZ7FnegrITGaVRIuSfiIikaV2hbenX8OJnM0e
UPuwo/+13Z6cVqjkMyYYVzV6RdaQU+Zp/K1fCMQff3LKUTgQstQapr6Z98cNbDZR
cZhwz24DHO9M24l+TucM1UGJQgnYkc7+Pvu3FX/kBLqIzHc+4gESA75vXKACxkIw
9BbI4uve7KZZFOorImRPSPo9a8qZerO9+wLuljg19oee8zKGnoN8bRab9htLbak2
S6xfYZIH/o9XC69HegqoTztNsQ3J6Qa5UsNPufiVABN1QeNz/ay9chG/tHW1Me64
DVYf7As07lCBWygth8v39TKmRWhHLFVQMjEX7vHwcHAZf0bhCSlP6g0RkelYFFcA
WmrG5eo1BYCyEenPa7tTiAYccu4Vh5w/uQwjFxhMMP7zYbMnbGn/09/opYrcoXWm
KcZhDf/jPVsEftpbvnAgjp5JKMKS7vLrRjYWEYJ5DDNk4tgHm2Y+Tkz2jL1RYEX8
0YfP/qW0p6hf4P8Qela+mCzuHpLnFC8RPBwKgv7bzSfJQVyULzyGHDJavJiUTMRD
OOh/IuU3+W/TCi1CKR7SD5Gh32Zxzl3S+BFn1siDhEVvs1fNUH/uxyBc794gv2l8
f7CKoJMWFwSLhIAqZ1t1AJKzq/nzxDDRJQ2KuS9CgEOAPSbKtLqtRv2uNYD7Wr6a
EpKDXhaxYy+RCUInmCbAJMA/fabU27l/VgGcYyZ75p7t9p7xrw7pU6CQwiMiNGtl
17wRvpBG8SE92G4R5iAIMI2GX9nlbmxMlbI+DpwgQHni72rBFqAwd75ijteHg/te
vKy/q2EJbCTnWMhT+rWBWpcmhVKbP/zEbpg3Uptpky/CgkJgUe4ehLHIrNgeW5Od
/VEnDC2JTp4+Iz6AoXi134ecF8iixj7nirEcJ14s0reGwdathb+Epibpj3GzqeVP
uiEyYkqiKKyrsRL4C9rREqGJZh10uNuFbNC3EYhQ445+40bzQH9IAb92kaiCt2K6
DfmYye4pYhAvwDxV89S/n8E6laAzYmZWHjn55kM6+Ae1xsM97xA6HOo7lG3wKZGX
ROBtK6cogV1PVT2HULCZEyLk2j1lqO29IMDCHniS14xDvHDYy2so2w1GUkLGhl1H
Sep5Yjbk9wmJxr7MKWX8YMMKbuV+T2++Chp3bp3JmHoUTFSL22cYfKrY8IdUibgf
OYoUsc4v3tTKyMY5pJegswgr/RAG2Q1ujsQf6HtwIcGjsEvImyQiVVsG53fhEfot
ZOTeAdOhq6Xfrt57KKziAGsWvRHD+sfctK/Y4yu+mzFPub2k3PhjMsOwzireZLSg
sLDHZkqG8hd+2CFrpsnCbsMWqcSJMnGdgC43bwzZJW1+jePyDIuMvK9U42GYr6QR
rCTAA479AuruDUzIqDFPSk5rjNGE2f7BbvG6gD6wrcP7aga7Mlv+oKlOnjJh6+1r
msYZ5HEJNKHzEyaUyNft9PLiRU9nqMEN1n3mfg9VmraCAdvgNevv4rznL40rUR2R
go/piZbh0SM0dzhXMWbrsnVrj7sXhn1CwJxWxigdihNc1BwYfkrpACQUMhAh9b9P
PdERVy/ZQwHm1FfjB65dVNwo+uq90rZYhpN2ZM/E16gB79GWP4aTv8bpHgR4PMxV
c+R+7IQEYe4hI7gphpUSJ3ypXJSxYXNzQiHzpJW04wrVAt1oCTPKT2fGJqshQRUF
n1I0Kk15th4h69M+XvySLSDQ3r7GAMclgnpVU7v+ZArIPDdAywDvQLts/i8JTNxw
wczzJlpRQWdh9+Y6He732n4ibM6jPeKTg8OHqoKxcuWBb1+Wh1bey2HQICT4P1UX
Gv12BLBLs4YpiTscE2M0RbNj6S9anuHb78Z+fCtd0xTHIjOIjcuBpXAOpl7urEYu
tAopjgE8z7Jb/Xd/9zSAWLtgcPKNnsny2E8J+jURnF8x6u84EGdNQHzVxKIcv8HE
Z1cBQIKkyZ6gWEGgqUcDfBpGNNdEgEI6TzL0AXVMpDtMOx1umsI9c7vlJ+SzbTSw
a9Rv9vTh0/h3LFsTCg/j2Qu34ND8PD7biGN89JdsKbgchp5Hjn4pNL6DbVOJ7D8R
7ay0cjBld14UZGRjvk3xMmnN3rkF+GjezIYxp1v4MH17Ocj+5S+FF5cAgwm9ecI6
dy/sdmjumm5xzL0gZFmG0DfpeZe6Ab4pO49n20bff0WBrq3tM82OnOD+Ihz1xOvN
0AsLMSPYELwnVBiug7l2LlrhGs9GGhrowYIcoTVW499umQ+ol6vBbiOjM6j1Rr4/
iMJGu97fEtAByzgucaZh+YiiBMEZ0Er+H5gVsACH1V8u9mq3gwA61OwWAPkCh/rs
Oy6Q9Cuzrz+M2KbgS+2idU5c5C/V7QCWsPqs8bvUkTR7tIjpetMBPcrHrXHaRGQM
GFK6XQFbFVbglDluxz/awAmsLsDvpb+IbG/OkgiZiR2z6r7LWuMOjTg5pgkXeGNI
YUSRuZP23YINYMeIlIBQ3h60sjH3Nah+WSMMdp5TBx15DfTEAhc7LOFuw/HylTS6
G3l/VGa5CNifIZxGJa61xE3ExGTRqifoNY/szveDrt/Fl4w0UOPbtTi+BrdJFEmE
bMDrUWro4bjoaAtcxYezkqw1iZBIPBAuP+slh+SqX+b9C/gcC9gU1DFiYuQqZ6hM
m/5szS2jCmKu61ZANuKtN2/UIbkO2TA8Cba8xwgDjUAv9LWRhytpYlAAZSoBdfJ2
BluSyTokTVChr+wssj4MZuEW8AO1sknKUvRx8/SDNSr6nEMEtS4t2uAq94fwCxbd
i6BDbjOhRRNoLQZzTgCQ8C7G+N74/6TthOctuX6Qyi5P3dgUUG/ePXs4jzgpory2
l88uzyaLElI3heIqi7x36jLWZ2AfiTILSz7ysC6o5GBIkhdGpK87O6oq1C5/ziIc
vYKcBmRmkuOrfki8Q5zTQDd4TVRg1Vo2fLEGkoWTlqsccwNEZ4XDYiMm/hNbYVAk
BUDx6YrUwkkmCJFJhXaZ0RvyEtZ44OSnGF+8mkjnrurP+2jxsD0AoTUremI5XnCT
1uDI3Ala23KjJ59OlGQwEydaBs05NdsQpt/euCPiKtrf1xUhNtHoDP9SqnPQ9oHM
DNJjSgZ/U4Pr56JfY9R+KjMBcwqw3Ny1WqKUrTh30oKb1rSjwZUF/9NbdHHwJvE+
gr5HYgQErFLZlwsGbvuQx9+kO3wD9OgNB1j9do6TIOTKiVWOXspk25Tl1ovhXa1Y
EnZ1bl3QFDZxYBwy+ULGZcqnCh+PoHAFpFre3dHqHc4qPqR0PJynmArpAWjbWOp5
tacQSIvy12H/azwXvYLDUqtPfzDPXR4j82sZNCmJlz3d46yoKUPHldn3BY/1drrH
KzivdGXh1nkxjnLhImun2oV+TyVSwwsjkve5QcO3c7ystzNFT5x1AIm28ltXTdE2
YNDxDWHAL4bA67fiSNZ+30QewiK55VZ2jGgfirASBgx+P9cCPlVMkT4KUTWhcd2O
ldgVWmh8j6UwH24VbSaqK9R1228WApBRbOUrPQ60g3CA+XVjtvd01DtVUzUeDEna
szZU/4fUkiS1DA22Gr+BAvgDZGPuKdVYjeVHP0OT5THTGRan8Cly8nfnfjyvoUGP
YCDrrz3DydtWwx21Dq6ZN42j9HRu2vRtyzvPvR9Q4Fp68fSXgvZSrv0feOAuwMyc
yy5gQ4W9NH2+M+wNGdYjOlGR1eSSrFvEXQYXOtAQqVsrYfduXPuD1i28FONFNsx0
yxFJFTRxg1fN35d//VyTxfkW2uPbGL3oCxD2GPtqHr5O7JrmU9Q6a89IyLGEIFPG
vKk9yWNT0D5wEHXjMvO5wzIZR/9CDS6soE5a2KBr+fk9xKe8Xukk6nIvNpQ2LZqu
04Lb+pFw3HU+BvrqI0HZwWIWms3ILWUq2Esn/VwQl/kGXLTwWGqsoTlP6Xn63jeh
HRlqkmgTM07v/tJZUqkMf4wpfTKYE8TiCHNyhdUOCGlsTs5bEC+wzFTC2y72iz+w
9CGjHrc8avyWcYevyHgic5LvAa838bhU0TtzbshynTJ4stgiN7+DmJX7D1rV1r2w
Zuai4X94IZleNbASW147/2A2MhioHIjytoUsmDzt4sWO3xhTXaRJmhDQWNP37L6L
IoMqBMnPG/9LTiM/MrCx0/4DXkvtIsD4cKPhFoBHYZq9jSYalpAYxSYz0+LxiYV0
qheYFSE9Yig2NL8iOwILZA0NM5HjHfrqgrCin7rePdWi0qA1fFJqVB3Z/uNSsg41
IrCOaJ8bxVhszxjTFOxd98Himj6457iLoFcKwxs30VsYaHEYvQYaQOuz5AKo8+hV
/0mw5iY8Xw62vDj9ih4fT1LCKKhWslXoIUWlZLEJOcYUDmJN2+BDl6A8B5iy5MJC
pn/+zlV2O6tQq52FYWCg/jQKczpYOLA/RVLdcMTT6T/6GqjUWjwJ0RTOtB9/n78G
qBshFlg3eXm51fOx0zI52lXWr3/RJvO4JZVSPA7j0Cf7aItyJtBJ5fLWu4S8WrSq
kpIlWTz/zFOQ2nk/rraXfupTTte4H4TUE/UROuNyIbPsXo70AjGYnmDbkavGEi+x
InFzOafrZZcdHdE5bylmM2wj74RZOUsShMmd2k28wX21EThvXZjw/Q/6sUvlOggS
Gs6ppOlhUSkmw6rI+cjcbVozmXvw1HrSO4eihru08qcGNUHcfiBaaYP24VkQBWQ+
AHxNzXryncEDTPS2q+7yLvsEQ3fGcPEMvDOyxkZvqL7PJNY6N+Jzy+JDMphzfyZ8
z3Lv4QOJS4mU8sYjKjuHEph0M43bWyqcbM2nLYRT7ZCT1crwS2xZpaVqHU5H2YRQ
w+7rx3Xx66MOXq4EzIX4RQsiuoKYoj+D3fqKR2Bvve/lPezlc4VSN9UBHQC6OD2l
xt0/iasxTiBkcByKY09h3gtd3ah6Om3MuSVdepud4dIbE+1cV9LpklAXTn5TzxOX
IfZACKdoceIcXGQn0kXDBziZCjLwqj3rZQlmSM5qbrW52SHBKKuKhfl68VZoZHUY
I6s6tYBG2ttS7+gwKfWtqYKIQfbO+1E/+gqkVIcyLCI/OSG3/Fg+0zcaGlCD1s6e
VnmP3c0u07nDYeyFKY5PmwSO9nQ4hZaZt+hulQVp6uGeh3HplTrD2v9yzBLQcJCW
rkyibKdup/+q8Dj2yWwO5xBt45XKXGKhD5xBmiKs2LiQYQvYiNW2l1SEnclmb3yP
QxgTmu8rwLkb1h4yaLkr/4cuB5Ubcmjia/rv5gja9xDUna3R8NCJCcVrQP5146eY
0iBLvHbIniAjykahhDa9fOujQjkYUNDawMIQztfEsS1ZrNQhp4CddGRb2134kCz+
Y02fqaPrqo3CyRR25myEGvwwsHFrd2ysApQwkoMhfY8eHTuiBFCswvOquN0W/EQb
GagI62+lnowZ3/cHDYRo0Wzf5KksvalbbeI8+yWObG1Baz1v3jgTijhNNnwfQM10
Tmnx04EVT8E/vnUw674lSFMXdDZwV/I2esyRSg9FDBz4BeABSmON2fmS2vh6g2ut
ZQb+sbIqrFoF7h1mi0ZfJXcNBqrDElfH2LQmsi0vXmedLbKX7yWxYxDZbei7jUMP
HZn//ldEPJgBZXi/zLQXcJnhLdtG7eaTLQ1NBsZh7QFPc9kHcSSGIiBpBNUVoO+Y
ZeDjVlmej13FI/Ud9uiHEhYI6on+78U6eRLAXNZEtQHeuX9gGTI6M0WPz66QLjS5
v2k66AMzg7BUJahKvY2yLA8ZMw5JPlyQmibAZpxLglkYgpVA3wknTdofJBk83E8I
WZE5i8rgCmDYsKZzN+KMzq8rR2nHA2ZJiX22URv53sZ76XdmtClHJQrC/bplEuOr
HOjFW29zFcs/UuUsVvm+/5R/9vhU4sTUYAGck2HthacLMf+mo9TlC0FYsx56Z4VD
zL1J9iI0TQ2tUWRqCx23se6Sc3SWQYoa6j7FSG00oFOljNf/ku6FXeMGAUeoWcip
AiTt3TgE28hJ0Zg7T00cnR865tCGhVVY+VIsObYBs79rZX30odYO3/rgJHwuiSfl
TWQdIrimpFIVjezopf1ydx8l9ebsbYZrnv/97iGzKVUChLAJ2YxGXFWb6Y7N8CFd
vEKynfHzoXhfC6jATOrRpV/Ce/8Xv4dAwJPKgWYa0WCbbPCxqLHsj0KJlv5/ZkYw
+tN+YP/2576Wz3lb3kqZgaZPK7ykLfkWVvou9en/dJGvfNHxMr1PjJVU8+T1A6FX
Svgu+CxgI2pXigRsS1IqDYEWXkusW/aaq/5f6LE82crHkNa1Plc37mGRqpDxhe20
qGpQy3nIsDHnCx2o+QRvEreeHD/E7ome3ObIScPmnNMzGbAhTiYrphmtk7T26jol
PtgHu76tMX/h96j77YLBVsjkMc4QwC3finVXi/kUOy3hTn0Se7JoRJR/w1r74sLB
NX06oodAELb9NROw/7NsXxLC7Tu/5OXzKI+GO3LQO8Sgqd1PxFzm88WtFAqZUQMv
PThi+36ujfBXXGRhKji9L4RTqqu0P10Q5Zt9uRllD9IanxuGU8qEA1nshyq297Iy
IuePTcmYT48Z47BU8AGmV86ty4iZGANRiAodKCkk5pLLAdH01pmWjFeH7oDbCwV4
+X53DLiDz/jIgkcD3GakeVVli/b/ZwRfn09KI2kb5yCObA5DkQ1kKCCOfKj/SJU5
P2EwRhMBxDhrVXDg21tjYvSuTthItzxP5CnTTK9PkwfpPx9kW9E7uGIGzFIlCX0P
IheqqX+9D9SYRoJLc0/g+tIMHIcGlQhs2Bej/T26an2daPmUtGUMie1Rda0JgQm1
e+gbzfuQQhkZLU5KxKeEbTSkjofuSJnISf0NW/JPXWFRKpx3hjJNBL0iHBP92KPF
9Uya1CE+UvBOQTlkVqyqOdMKo5dmvSE6/dErCK1oC4BrzZ7coNSqO/S6dGmzPPOi
PeiqqMlcOk5IrfLk/UqHOv5TfjUBRm5ilhAyr+1ROKOggjIdugM5kU15Zw46TWGb
1XxH1ILP01z7rchjVlBMLezZtx7ffVtRop3aCZrop/8qm+3JCtFiEnTAQ/MJRqBF
frWbam0X59kgqIIHJKeWtHTiwT2CX4cmv2IoFOKarrMQndlzo3gjOHCcEOhN0e4v
65yZn8U2ECheIPDR9eqZtYix6V3qmUjPR2y85BHHxs43RB8unuYFSmois9chrp4A
3VczkroUQfYv6HkD4IGBBHvjTBe6fYs7jYsTzkfhFt0audhBVEArHHHeiC/25ChU
QtKRXwzz6cxH03rUGFhjgZxs6v3I71m015zSH/DOzdG8FZbKte1Jq8nTbYtqyhkr
NQ4shIQqKsy6NbpIxozHZKecFK23sbeV6CEmcfB6dLQwzNTSSkB+HNza75zwjQcw
Z+BMlBcNaDkCoRyi33AtB+RiDc0QmTppGsCeMdgj1DtHvOSXD06+bi96qVN83igq
B9avXhlU7QOS/mqEfQoBbbJEDBe++b6/6dVmMOFfvlrMHQLt76FlGKp9pm2ePY+e
nhzImE7pYa6qYvY5xBlMRRbmrGfzRis9TJYXmAjCdd4J7qSFUgwLblo7IX4vid7M
yn7Yhka5X6faaDrVsscU3RPMEP+4tlsmHcmgmW2xU7QcPfNgiu76amtMp7CliOwm
tWY+aksnZgQvSEWLHAG7/f3HWd0/ZMVaEnwRSjhjy7oPfZdLSdVqBQQlUQGS75dK
kIzJzL7xw5qJDTIx45Sd41qYVbx3aSSGe5kcWehdpztaq5salGA/acCgbn4F22Xr
V0mDtTETMeQDgCNA/Xs+pmcCtA/H4ujDMdIpsorrlWj/9EidjQsJ0HnZTH763gs6
pwalXpmJcvL78EXrlD/lF7rrnOFAJZPqSVSNtmO4mGxGI+kQbgwrcagiIXRK9nt0
midfZHJznyQUNGoJAEWwxgwXLOeXxuNjEwuqQRM4umatSR7880cx2QbBozuB96wJ
ofmmtTAvMMj4SjW6N27+iuridE36RaT1jCgpWQcgzUMKGyd5MfHe14MNGuMGZjzR
0sd9IXHGAkg/ZsKLUpB14pNXwuOfD1d/rL7o/DUUzhBAbb5Gd2jue9kbQdFnEVuG
OUVMf42XM0Vx15pYw36nzReNbgqimofOj770W+u279rLBEEbNhc67wSb7YrklmI2
/9pxrje4QDY5KgRK2NdQBOj1k/QK1nUvf9Y7R62fyHLv/PX9BkOKF5vzHtBOxBl4
TZQCo2bBtz1cflexkYYFaEua7yV7haTNp95UAWsHqrbqdxFERHQs6l9vQwObxQUq
dyTX5wY29BBy04qHtJM+MSBBP2QigiT2+2TY3SaL7COjZhHRPpDBUVVw/MPv1Akg
miCnR1py1OiATiqCzSiah9rRdqiAdMgyjq/8NOuKCfiySXD/9WafJT7ZbXyRxyAn
xGZEAOifdK4MO4Bt+StcX3o/GXNX+kyx+cXE3ZREHtzExdGJbuhgsIIxFiGu+Uli
1EwLG0X+nMJX8PskrzK1KH1W/enycHmtPEzpVius9NNEUJn4dGK9rVi2DhjVuBNE
3CRbuu3SrsvIg2urUDXMYhlRWOFdMViOuX+Wdc3R4Mnj2wAJQrtqGMm9AAoGEN+O
UOqClCgmrmhUyeO7Z1a+72eCzY06nK+xIeGQhhhN4aEPrDbZ52srdopGU+ppukRU
/hiKny2bAiawn0hUQnxLjlolcCvRaod7BbYNEjc0GwYXwZjolnpCZH1BTxSa4ZH/
Ni5klllYOyiZ8YAZSQog/QrSZL5xgHrAGjGDTNznvIdEmGlvrrZynwLOxgicDOUQ
WGmThgA8YWDcG7QtTgmu9YUcfLDXAPTFDLDEc4mKXYzut04ntA9CtrXFLXJAnhYY
OR/AK0CJkl29V3/EuuvS/+qQA4gAdSTsHoWdMCXz2pNJlvsq8XvL5+p/29Gpk7Wn
1Cur8Ae2NNdEYLYplYq8S/oHO3TIO43yjjmqK1KVAY1s07x41Si3HnXva7SxAvom
OQHcHL8oz+UjWhJV0A0z4B3Q0s5RHUIbQw5TH4Wus2qtpQJPFDJ2JYkCDOmUJSMi
ZO2szqffSSHCZNQYq3VS1dix2DOXDDKbkPPXFjt4zlg1OgTSUbf7uGgC6JFeTL9X
bjC5m/dMmhQqO0DlizQQ4Bcvfu4QK5vG4vf7wKiO6I9qNXAZKTS/54sV96MA5nsp
lvotiqUx0RsRItENr8pLuTxnf/hMpRWHlR/mLPzhBa0oxN/+lq9Iobk7Qa5opsTt
p7PUcZiJcD5CvRQKZ38+Fmib5PH9f1zablHmPm/fd9h89Ku+zzVejYK9TmlJRXFT
WAFZda1T+x+FZxXDbw1LAkuxkdvzrPRiDMoMt64mPLVJUEUGGnkIZygHKPjV9su+
1Zb2Tb2716NDmp0Rr8VNPPsZw2WlI8gc4RsJPrMNyTytgAZA5LvdASlmBDsN3NVR
dIcGfdHud5s56UHzAbGsgHhqU/4M/SeFHNg/W3cX0EI8S/E5hYWgkRPyRtMgNi40
n7X8C89EBZbb1ODarQ0IXQHE7MBKMhcwIAi5JI4ubzcKV5TmNKE63Y/Zb+HVyesE
1c5r7L8PdZMMD8nU+ihyDNxAhP3YUV/ZNqbBxjFy0BxABKZ9KMeZ6CbdBxKmY1hg
8eMvoWIVPpUl61srovFsj0mvb03JGYvElSfFZHB6y8bovyYIwEmAAbWYlDIRd+Vd
/bMbnICdfIucx4QONxg2Y0vJF+ffWw1/2P+yP76R1xkE054pADWFLTNT413KjZg5
x0vi5cagTOUpq0XC/jDDdGBTIQUmVhrFS+noCaiIGgSpc4p0gfWKr9IzSiYZFCe9
BsQsBEpM+EZhP5mPOUvUZUugta8w2Wf5pxP8eZ8LnIdJCMnwRgUKf7LY4QqumKQS
tQsdYistzrO5x+pov5dNkjRShreoksQ4OC38MYTC/fNtvRA4iID1kGLQqbtgxsaH
C3/6YF062AkbhHLDbGEHvW9J54q9izAbPlHYv3SKc8g2yX5CqV8RyFrwVCyv7kao
j21KOKTraXFHn+KMrQ+zGSyf3oGbB96p+j8lv8WJSa6hYf3f3p6O6OUiL1cswuwR
RNmhXSMe7zLNqj4pqjTOqep8CsI9OfoDv9au0+8o2qjkEUDkgLndKafKV0sejkYP
AngWNKR5LeY2vG9zD6+HM2uluulPDE6z2fZEDvlARYz8CxozDsxqzKhgaQ5Qzgv3
Qj8mcvXa0YG2QQEFgHLps4HCdZcORd/2PK5Ncr5yoH/w7b6s8wFj3fmrOpnWRuoU
VMsx0baO0hQ8XhFlkpw9KN4mgcD5ruwDCzvjDmVETGmdhqWFE+PSmRDj8M0AFGuS
6aNI1oyAn/cxi/2rZFVUOEmyyY6qZGOyGNUXOehZIeSRxWLfE1zzEiBsJK9vkjhO
pxCAKdGB/PwdcTbZqlI04f5hwXhI/706mNrt4w5vBrBdh2BctEXJnYURoj2wdywr
kYNtQvnawioWLy+whtGqyh8b+d7QqreKRKWrJLzys6yfr1ANWHNpWi98WrVGxkXV
XKvRTUnSn9ZwQmWBp1MZFUF/UkY4pz+57YSFp+xL72MTbvJnT8E59g/yNOttzzTp
yQtxlqyZHBzasOig3G8DUsSYRd2Ds1Wauw8c0MeqAUZnUTp4nJBhIM1wH8W+BV2F

--pragma protect end_data_block
--pragma protect digest_block
9QU8lfdWZjChGFRxy7TbPu5cB1k=
--pragma protect end_digest_block
--pragma protect end_protected
