-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gn77er10B0kUCI6AqxoRPRORX3AeczJ2jS15mHewwg70FatFnO5i7JwS1TIEJeLp
kEHbPtaqRrUftf1QmjzFj9FhxFMXVJuqqTpVKjCn6H0lp0dBFXt6+/CtME3I535y
FfA30YU/aFGeMGKJifwUitXLCTo7EgwgtyuTIHhBQa8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 111438)

`protect DATA_BLOCK
RAltELNkr44RbKW4JZ783NvtAT4nSCVEbmXiyIxctPT4H+gvIcUD1247D1C4ra4R
ZQT9xDkPB0c1MrxypNXHqYrhrvUaVUwnCIUgsyZPWuRalTulhXLWbF+OnBPC7gwF
MoASxVSz5Ie22bl6gqNm2aEPkjjNyKSaBs+68iF25JzS+1ZcAvfJdN6m/nV9S6Uu
R5RY41to2vh0wwbDHxdf+pXtS1JWT4euJlfJz2EGN1MaNa7v8a0XSZE30DNTcmXq
Js/4QxXzriTAySYlafbh6PG2roapRCMGBDcF6nd2wUtRt0ebPCVBSxQFWjsptw0B
ul74FXMy9n2GGKXSkEY3Gz7MCKiuUMn+Z1YTtdEl3DuNsAw5DG39Iv/JajEYPa5r
KuSajTtSfn+IIcQbUQbR9/oB496Xzikuf5mV9t/QsWlQkXnVvjzxRb6Gf9b9kK2D
4e+XfQLRQA2AkGuvHoMcn+e6bFRjWcJy/M0b4tBHON93pCw03MOX97yrkJDDYpC4
PoMJAXmCVpOQ2zP5kaE3sa9UmDJlCwDg2yQRg9YCFUl7oV2vNzg/eGxUo2H7By/P
+9giPljgQarfHF2D37APM5oJg6fEjBiXztZpxl13WXy1HG2exv5t9VTNsss1Ol7W
GNVbaRiJK4y3E+4jM6M/BhnL800fIy127sw+5KRjk0sl0UMEltJLqnk6okIsRRnG
XpplEvoa2xNQqr4ctq9t3eAqXVVfur8fBybrVJEeTD278rU9fecYlIJX8AJuY7Em
DxN9/WxpD7b9nfhipEYYShWbHX7mFL/wIjrNj37mY/f97Ty8z3/KxAKn6UxzZAdq
t9AiAWORo/bfWC9PyyFeFAJHpwe3O9B8jt/tUWvfJ4VGWwARf+PFBmmMbiyNjJgz
8Z04Zs/h+jPEGrnMXCroqPMhnX6e65ylyNMKdaZGtLeY5caeIpYLLr1+XdNwTNkz
D2QxTAGw2dqoDj+8pc/wGbCdAGhlM9Untdr3u9Hd1ekXlfosKRQk/RBdssvonqJa
8a7sjGwlxY49UTVriWnZHMxQ3HNDzkC+N2ROCfLI2fjC2GMfK/CXlXPGHvENpD8Q
zUE2tga1MYglSPZ8nMQpDj616OdQ0dDIt6buEt1NIQ1J81MtY450VblbrwOLF33i
b1Fl1p736I1Ke5R5PcG1od5B+r5LVZ5tO81WCtG0iPavLBzWNtEJAlfqkAyB1wlw
/ZSA2+cE78F6Ub5Chp8Zdd+LSt7A05aKbUj/S81XAAEBq551DARETMRIPMIYilis
6Maw/HNWrpF7dYJCkWlAxb2R3wWV3g/pwyNEFU+OTMZkdwyfI2snE0Xfvf3rVtAK
xL2h4s6BvuZbDS/d/r+alJMlGubt+g6YUpaPkYerERtu7fztbReDfxS0Dmdrtkdn
HXpgNiDcMl1YNjC0cck8h+J7zkpvEk+j75KyrLbFIlY8F5mbNIOQmR4e4EajRNY9
rAQpgF7tJOtvoEvqhCOUscluCk75G55IpQLJWwYr1DmJjtwHr5id6y/StAmgWLCN
/GZglq615OaFPjAl8I9PZCDvlVrJFyeQ7Otx/y8aCpOnPoMyKjpzobcMw4p5nABg
yJTtKJJZg+q9C2NefZxex9NLidINLjQxpHWjklWmSSwFiCRL22TMLzyKXPufjIEd
CUrcCmoloTBcZStbLfbAq/38gjbJtdir5xfgzHaOiQ5L1p+xu6BAl+UWfsMyfe4P
WnYqFGt7Is6GCjbwZnsx81yD+vn2t4dKK8W/ADJsKlH7/uNI/xyGlv+mtdr060WM
rE3Gfvff24UQsuuTxAJOzRz7p6kQxK1QA7O6CP4IDc0mmAZSPQoQXImJH/1+Hh1n
VOxhNkgxn4yGFPc1WAguf3jrorfOq/lRuI5MNlBcRoePtLTpgPCmyNOHRnSPm76u
O/dMkAqufV9tJEi/qelYznUmbFj2nFbQcXNkZpM97Q3GdZKbUhpUJfw9Nx9sT0Gl
JVhzx6fNTLleCo+/CYeSSJKumYqQ3YvUaxOxoTTyAzEyi0D86TGdM2gxQAIYgB+s
qo4wNunnXRMreKvEPhjmUZrGCtguQPFm9SH2eQBOkyAaC9jLBHomYj2W5VNG74OT
3HhMkD56wKZ+BDInLtKsuETJWRzG8YMOpxuiCKwnM0nrEfkG89WidghqaGGCuKKv
Nwvk/OxUWwO24TaDF2K2w+KUp4/s0bUt3xaSJ72Z2zTVx4e1WCMe3d2RHO4fzC0R
baMQnjbLT/mda1tmljESy0gF0FcXpkPFGVxr2hIFFFCOnGYzOP/IKlQ35Tr1RSwt
RWsr7YoGnutMolYj7H0YU6iASYTYXd7JXryhN4fMLs2b9Ovlqyian8YcOi7TJ5y3
EgONYAde3zj6OTS8uGe+sdp4dQqKoKE1seOaJNi3IkTgxFQbGehXLcnM+ptA/iml
cNwtblbjnja2p8ZLF++oXYbbSmMX3nQSaXpRH5XDy/HFMPvciTiu+qFeCz4WmfZO
sitld1xmHZ2owndrYXt9eE5VXuo687og7LJrJp/27M3UT5RBDw5znAZrjM8yUdNU
XFYrfWGkUIQ9Gg7yAkG0mFD1Q0yw77RKFUVBC9PJIGXZlyNso7BB8kr0QDfiKkqi
7QFmfaw4/J0fsn4+UxgRZ95EccrqjY/kh309G4FoDFXJ362BtyBodOuTKVf1CG6U
x1EBO/WnizqIlwi2qw+C1BhcXjPxlU278kx3u0d+YinfJgGLiLXp5PxP4eUi07pY
ivmOEilbXGL+1kYOZXl6envS7J/hbBKheDC110YHZH7+035vfRh/U5+r31+WoG3B
pmts0J0BXGqzlcjF5vRlbSR5GD+DkGvrYeOZubPBgYLIiZOrxaqJFAo1Dn5263ea
Tkfwh6/YhwGbXf54CYSo0l4RcDzLrFlAQQNA02Oxr4xll4PJzmFoMRnAu9twSxbp
lqggp5N+wEkjdfLR+5NjVKzjtjIPOWqwzZvuFMKp85zI0cJ9zDYPTtaEiid6BF+E
+T87390Z1Ur/Avx1ON0SbTIJUsX7HuvhJcNaYBrqgJbF4VvLI4cFd4IMPaZg1r7x
bToCn6xAsHc5A6lp/vBy4GL0dl2mtXGMKrXU1oamSuoPlD1c0eoYsc0/pJ+tC4Xj
V/d/3HZA3IHer9ULqvJL4UsNKN7heuWy+VZ6YwCNWdDUBB91FLoqxjAslGxtno1w
V7fVKGT8clDRjMGsYVtxJzfUiUARcNzsnpbmJ/XAmTG9DcR1HpQGxGD/W6iOzJp3
KxLIJEhZqJyiOnb5cPmDVIEX8r6CDvy8WPDp8tjh5UxRScb8zwwPZAi55vwWvq5n
LJUWIb2CIPl3G8up74DOD1VkkAuJe+AoDPvEX6l5Zxm6BnQgUYVyXI9doJTx2KfI
Sp2Y3EE3if2yG+yexx1CVSai0E3+HBlqsmXHrKO/1Z4Ip7IFq9lAtfxpHmpXIPSy
xhHWTNUWrTI32rHm027DkgAaykEJAazZHlGIs1OIJ4mcC4WFy3IY1tBk3NV9HE+f
Y5535CAt/U51Mscf2Tg1cgWBh6kx1UI6h+W1W4aTccglYcZauQO7Otjp/tuPr4pT
ONyGNrXPSECIIswAaVNi3k2Y5+GDa+ty7dS24M/4vcpEeapIUaZTgNLwC443pYnu
jtBwtDqbuuxEi67V5N/OTfrzLrN8RsCcPtnQmKcJhmP1sqaKAkIRmLo0XIYSxVQ/
+iLkJQB3yFRU9kxi6zvsygdSooutTK00OcW9BIiPlKBSuE2uJAIRp3fXPvOm0WrN
nVNpWmvlu+2pOQBTG+J3Vx5poQKYwTsz/28ksHacSJmI1aq9tbuxl1LV/v1mz/o1
Z/uSdxjhNKmwyvFnAAe8cJ1H96Rr8bCtRTTzToCEr/9l7brERssmBWG1rcs49FF1
nTiMtZEByqPDfru1hKjn7ARjJIO/RvCl6jdgUJ3muHJRtAtmhL71hQeDfcofU5pc
SiNIQKK8ItUHKWPWBM3+iwAC8v9aPpA/jwyHLzcRL5RY+O0NVV6hnN3nWSdY1Jew
mkNwvZcKk0dO2DN/OCiJey8cgimJLIRjw1vCyHmRkmH2Yj62RSFUQPnlzhyCNAV2
5AqsrmP3UCmdK38Shv6G12T8VbSfKdgANP+9PysSaeyQsb6jOzYyyqqd4+yQIp4t
xtfgYfsiUs9phtdpMCuJCYBliZXHYB4wPxmgZGMGD1NUV1ZOWMcF0egn30GmWnpB
EFansEsAs6/YLpJy2Xy+zfXvQUDPj819484AECVmQHopNsmgwaTTr6CESek8MDmT
oG6XxetHK5yZ16/WM4v/x8HK+6J4iTnLNphMmxgl/0whoXmCMXMsxefl9+euIIqN
zP+mTlcIVvaZnvCrQMYVLGYhrtA3RhOE/a8rPX4xQbDqmKAjv7+GkF1q69qe+kdK
HKl5wEnsEtQguIt00bUPBx7z0xcYtnpqJC3vNtfxiw+uX728XbljoDxpYdJm8ikD
DlMiUvrUFovJETX0lOhAhftaEBa5M9tu2rYHoyy3PZC5vPwMtnlsuaYCpK/TBRoQ
edPl11aj9myxBGxgjgYsBUe9UyU+Czxhpa8oqHy8mv5qWuyQZ4MQ8OI8V+VBwdX8
tWW9aDHDE7wHfEdNch4eGOBMJLBVSlRDCT0QytXpFBzv01Q08u7XKJyZXSRzr1Ur
BbTkTD96BEZnntmvW3LwFdzyRCxWNBWlbm+iJTVAoqQxovdPkWSeRPiNB+CrT1Su
Jtk92Gig4OPtXzCxpcDd4jJgP/25QoW4SBeu1BzHljdu5Dr1DuJLKSGo1WdiewBi
a98IaLKYOii92hRvNhWmJ6d8Om4F86P/v+bVq12g5lv+SGMau8MT0UYGcafTkHSu
8/aZBQlYkWUob4rHFpshjka0At0TMyKFZtPCOFszA29PuKaXN4NuZN3KMutu/m0i
3dDp8YewSj+GBc033bkPx+vhpNgsoJdhH5V7oFixfc5CfzA18Fk9CAaJVDD8Dk97
68gV8CzGrEYLr1WPv34+F8QDQ2y/i6WN95w/RVjpVvxi82B/quoI6gbzfh5z8ihF
ATGYyQV2iA4Jqec0I5H1jwMOXHvET5AWIMfCE6nKkTKpcuiYhZWg40WD5Qme0CKk
DPeuda1PrHlkuLCsbrnw9VERb7fl1aW2jlpHh0lCjSeS5muYQGexDpZ5OEmhjmes
fKhMzptElTVkE6Fc63/HSv7kBE/9ZJ5TkF94fFALRkbxS6jBo1Xp8QE+17lmqf2T
V1QVzhJUyug1GmAzrVIODjEixFm7FTwnv3AffGOjgUk9S7fUilzUJH1zAn0Ai7Nm
mVZrjKADbaYrs29zTBa2NO3WIdDZz8kNkAn1sOk5c5Cbr+G0G7kpMN/3Y+Bg3aG5
3OXQ0e/BAIZh8axt7VMASQM/oK6yO/lHMauLRpPVudwRHW6A84Pf6k6tyXSERGQJ
QvqM3iPIRcCoZdQGR6VUsBY/Pgi1YoBhPZjX3minjzXoc8tdjcEPeOLR3hiRQhqo
1wR94pH4jFpcPV6u58i8YepRpBPldDxMEwDbU8QplzGe+G+IorfaqBRbDO2UKgnl
GWceltoPiDHQOk3HvJ1kb32Lp4KHS7UBSuNIPtOQdrMNz1RWuAuqdCH4+0WDfp6A
Jiu1noPIhg4JmnjaiM6jFAxidt3Fg+X9XFm9EWW71tyDbyGMCpzgAsFTW00yHIsL
93bhdUEuvqkNCYsmLVV4nVXL4yAujbWYSzjPUbETIZMRZWz9NzsMQp6me7x+A3M0
+j0oUXgI2vrEyW23gn2Y0FErjKfqnv0zdQhMxmwDhkMlsaSGsapjyYCnDc6OoHWL
k+V9pnGbR4BypoQ1uYiUNnteP7RxzdVut06YgG19DyoVlGQAhoFfhuBw0Kfs79OG
RiEdSSgL3BnKkFi8PcHKrw6jgT8gKszPbn19+OnY5tJg9JQpFeLKQl5hK1PMWHTx
qcCpc+CKSDXa/BAMDQYdNa7F85T6SaMovTRxcAQ9hm1jAiT6qJ+LKewjeSN29SD4
B9JnD/ubWZgS9XdFvLxw5sh8itQzSIEFEFezXwqps7maF5IzbghDX+umrdxJOiu1
4yIN1FqJ1AUuj4neZA+5ydJzeb6LmU7jptwmPGyb/eh/FJMBjQR0P7dfFNtJ60zf
WJNqwFg7tkk9IkQMFLI0AUgEyVvw0ReDwlAt30LRRO4zd6DerpAiK7bX/bfexKIT
4EvHqukohSuidmPcXHToV9c8ZIO1lkZ6yQ0u7DBUX6EU+UBq/+I8LRX/qqoZr5/Y
Ky6If38qTUWQP2oiye+czlFJxiOeC+oTk4qchgyn63tXA8KHDA4jVxUvY9nhRoAC
PS6zE14//cG/VpkzT/mSoPq6VnKscPYEm6v4FUIbVmJUp0AX1OYk6NSIcyi8eUiK
0j26byOLgL3los3j/RHPhhSaWzbnGeOMUTXe7Zj90GYk6nrk3VmD+wpcw3Xc98M2
BmzPEbLQ3JueOtlKf86QstFtire4SVO+BQXZm25yA9vLCMfwI+2YmJRRM6Ems7sm
H4NjBkxMynZFUze8w0TCwAk8EyABgVGS+MLmJoo8WKw3D/1IA07Mttxjy7IOaSit
03xsmt1oRJ0pR7+dDK+L9cNV21Jq5sHdPjkPFzWKi8i0PM4p68MCdSZRJuIsgjYu
ORdMQMk166wUP3YVNWzvDehbJSL5ZzGoHNl94DBAekseLtHzSe6EmS4lpAfG9NzL
0/kWkCLD0zgXj/WLYSqCZlY2TJJrHmKtkTuAzHufzGPEAY9bDWNYvaxV1r4MXuSe
ZyxgH60veMZip3+xw2MWWHV3peryFk6z4mg/LMRxaIlxlQ9f/cGH/0vSCO3jErTb
T0IpJl2ddR7pFdb4wPsKkrqg39giUeYas8r+F7oVIoUV1qhHQVXSERS/FhLPBbYA
YnCjUemTK8bKqBjFrF4vDYhnBnh+UniOD+fqnIS3nsuTZCk8fqFRa00EXk6AYdDS
+w2ovc/COdXpoaCytAqh81J2+BARDdd7NEVHZOCkK3DXFsqoo/38ZCKfFrldV1HQ
2piARleWG5cuvY7nCvAFBNuAekRHJcJZ4hu+cWGTpEZ57n90IAyEuyWW/kIQ3+kR
746WEW0g1pCkV2uDn7sVjw4QYI/xoIgF0pC1CBRCvapDITBKVey4qXgx2C6zuuMa
/GXF6xIut+hUo3PGeFiRsq3giTB2w9zVteN4YkZuEKHuCgBq0Nzqf+JXuTT792fY
XEJ1xZZq5mN2lD9r4sg5IPEQZD9nvKHHeANjHbIjXxP7IXEENoYIzKLZGZv8GFV0
9OC0OBu9seYv5Dmnoia0V7MLMAzl09WO9sDvqgiX7ZUs7+dndPhEiwOHhBi0Crni
ZIcQqCTgT4/Ywy/hfmgaXJzxpkBAsbh1VhaMtbCThOuzG3TywLMylJGWl95zPmZK
rRvoHBL7p1BoqtYXinL8h2GOPnC0TdupBPHftCde+CcITlZxa/F5xVi3uWMK/rY5
3lAKkQ13bXXoCi6GS+IyKSxufmm8DpHgXXaW2ZK4k4Voqgd9f4/ersouIfQBGAOG
wEf7pDXmnbsVoN4QXqFYNiq7FotiConRcXAmI27zSGhkHvylbiWe5WMEUcWPYsqI
QSk/juBl4VHMA1sYg2I+VElKndN1Q1k2kLuv0xPo9x5lf1CvCRnyPxUlPI1UoCty
O3T0jyzhybnqfoMHuMMEKJVcQKCG01ov4IHFTNAeqLKmuR7tKjzPzCbaZK5rS6+9
/bE97vUsQ4jqKzkws1ieUsDiPMUYC9Jy47lhDWbincB8rFpCDcJxWV/+/FHNBK7s
up7r/DFQJuLS7zR/i8GlzN9wAld+Ypkw8GcoUsLqQHXn+NcpNAaSYt5Sa9Ac/vPW
l/A3017z2XY2GPm1WCJikSdHLwgVmMQQchC7wzjHCYb8KCw7Du1jmtA+LuLql7JG
e5xKDGZ26RLNMyMNpyafduOpfgkyPKSgu9jiHixwLRfuMKXwTw0JshGJt+pPlRw1
9bTFbxu3/25/rejdBwBTymTdPW/yPTJohMSVgjm5e72EgBiUdQg5HcU3paF7acTT
Sb3II4PPVGJUhwBsI+UAvZD4MUPwjyzUe/tqef+5Xq2bo5ApnHCuHpPRcd/U5y/M
QZUL2IEHsIJ3HbbbT6EiBaNVrYUfpcKWoydkILdDloMf7ImYkxfe+KFeZOTK7MDs
vw0VwVnlZhBMAc88SAI6UTdC0YK0jXQlTQkZl7d3HyUa/lPThGnlNZ4kWPonRFtU
5bP9z0TX0E8bzY9tMRfG/oWUpph5Rn19IpXcbiuv+P/7quuGeglD1xFMKVYtTL4m
luYrcTg0mpkL6AIyuOYyMMCtb/3cEPWc9CJWbWEgXT/cmhPo6S740zchdPAjN6Bq
FidipADpbn6gFsVWCIgen3/l7L0NAzVJsWfhqL7oyPq5Z31IdLe2QvBAykMVlQVS
q5oevGLgLPWixhxiZiLMsw3yL6WRdUz+GbWsjzSGxmr0gzyUB5KdoyKJma7+TlSo
M/rGdKdyQAwjSg0zNgcujilKmuh+sNlWMxodAojGQnKnrbrGecEAeQM9Giv+h6TT
ldwj4wgQ4tTfSvhwpvZtyeRqm++7gTHhI/da6OhlFLeh+katLoTnapiNXgMybcWm
gJ9C+hRd97PjApvEMz7VAUdmrJuFtWx5DHxoS7mnnYcekpfLh7Thh43Pyp2klhzq
3FtuFUl9x7DLYkI6u+l5Zec5UsoskaaTqEph47W7mb8IKXF/C7MTMburKCimirAA
VWDYE7y7VTXJrCBu464OSrScpN0gxtLlCa4Vu2Es1b0XBc0VLzhWEoR+eNK+bGvW
Bgy2SDMDVR3wfp9BLQIigaoiGbbquRUj5KM2R5b2Rem/us6b1Vhyy6Fw+YIX9APt
zDdwGKRZDiMzcydz+KCDK5q0pjmfX9i7dt2e0h7cxA1ZofAOxDDqthHqSIrZKI4I
fOXVExVYB6BKkV7eKRfzDpzinU1fxNjG8i9DmksFNEf2uJfpdS0wJo2MLRChHKOZ
MAOYEIxslQjQndCVMfC0En/BevWqeRjLoQjfcv5Vtv9B9VWkoUU3zR4x3o3i4Y5S
eNHSuvbupNmN9EaZfb43B7lARoJsbTkc+2ay6VJYGk4AuDO10aV5gwnN+JRubf1b
StfG6pPutahc8uKziGTZxNhpB6Y05P1QfgAZSpREdfAsbh4FAN9ONVzwK9rPQW3L
hh2aUC+MVOOUMEZVQe0c5+XbQg+v0aIg1bSHIADdTI1dVX1itQPPMmxKDEIl+YOd
j6WwFYMmdv4rO7rhjzuC29wCYyLAs3iMPjrx+S+2sC9Ik9s4RlYUhFyi5TYjmgdK
lMz6Q0stzrqKRo44uuKV1trQFG2seItxiceEcni/t48JyJKOmBFfaLAROjy6VMUG
h99ZtG8+MULfzKGrAP01f05zaJgY08v1NJpDBk6aRQOWhWMGOTEBfqPCtrZ6Pp5c
1DwNZimvzKzb//zEtkrMNORDEQquJGYLiYYW0bt197p6nzuWBO764toqst1cSpdf
OO/x7jN1U8wK+vkoEQe3DSz0JJGL6HvGlZmKY9p5eCOUQ1FtTqTWSHPXdXelIPT4
ZXs57sRpwSULzU7YYrXPhpR35i0qcRlCdD+3dNZNKc+H7nitg1rF/w4buAGwHNx6
qgHtZPNdwtzdobJsc8Na5fhIRLfvmmrWM+jwgwSBhlIZvybVFSEikbAW2v4qxdLT
tSxV3+8hlSIRmL3WpTaDwIcrJXJL1HS81Mt5PTOy0QtqX5isBDz5nHr6H3ccFizd
ERu/cTnRa1cDGJiBicqMjum4RCn62wPImWAIbhrnS/o/v+X9+lIWH8HhSrYPmiqF
ZsI/0YGnNn6sORUpzz28vCQawsTXpMvu7gqTk5LR1XDIKP+zr5RNwD0NEKbzwY82
HzmD3025RlCgkMc7ntIzeTuYW5zyMDTh/Vw64Mb6AQb57HVq1HrNanZNz9Eew6We
Urxsx1Yy3gZKOBf04gliEzTWZQLvi68YQraVf2ub2O1XiPCVQ51NXfkrc8c0sNzm
PIWZ2AL+1LY2e0bIldtliIzqlSDhPI4qssdK7CS1ai/98HGa8gSPZdN8BWUfgoii
NDqYxyCQaNRCN9albin2B0sXrEdyZcqUZyPDMrNqEWwHYjxpOTRhZl67mSJYC+MG
aKv75JyLUd09SCHlsHdiAZvdNobb3AIZX2auDgig6T7z/xBDeAKt5GMARxtuMvqW
yiQBtQJ/nJ+1j2ga1jA+K496wb1mqex+0rMY7sXxaMgXYKVsYPD8T7VYEtiNBP5Q
SIOTlbtjRD/fS6BWeJG38PCjy/t8StKjMUwaw74B8f2s1EDEMIdZwNbnDcfL79uS
yhpKOD7PW5W4tIhyXiKvPSAjGjhsG1OSezizepmvlYxn4W0jjOLDOiRSX3+nIEVe
KzsaeGowuVdnzYVR2XUnMRuFuvSMJfP4Y6WXPdj/+fUKlfW0/hNw4OLfeLYYKa4O
Ef8bsIGxQH5Z+UQCgmCtPs3+1L0+ovoZclJEyD7PRRnI8Xi33mBEFaGWiiutXsfo
xDTcVetzdWIaq38F3vb8/Y/Z3d+rBUD2iUlnGR7LIztIPzcTdTiedOLpsl+0vrqu
Uyil6Mn/Ctt9kOC0GW3NHQwN5sqD3gSEelTZEfKMroFOuo8C7dxtem5FL7v2NgfQ
xMHWXuFtxGNyLn80FqN63eCmeRlq+MRcMrlnMu4zHZky6Czt6VRm6RltLjwactfM
S/D6A14JTr9VQ8OIby6PWD/4ctnELgtAItHkSXL5f+cZMuiGw+dX4DRqDOh+FAHO
TJnHTgMsV5x7dwydlLsep6yWsMEsC+RWTSms736M4ADHQm+a0HA/4muTO87ORTsD
j8iTIy65Cz00IUQf45WWCIPIc24NiiR22rLbNNXdcIKa+xjujMJ2o+9H9+ElWd+x
bygvcXmll/gmjPaiBKfo1aJvw5lUFjALMP0G+SHN6xbeTmRFtqgQm7E3m/cN6Exc
QTkf4FyzBssfFrGQOeNfiVZ0L7/BNaf9AIljS+bZ2ABZ3r1A+9pFlf4dSSCyAPpp
AJxazf7Y1Y2UlWUySYpY7fgDspZdShyQvv3Iw1IvbXpjKa4dXBJNXf+vf6Nyh1FC
FSk4UYZP1joxX1vgQgeNm/EhJb1DZIfgymKitWXmTsw/uth4FTIqOxrl4Xzm1OQn
ufv+lCJ2+GYuzsnhBc6kn91WzqqJE2po0CZpareAgWvyKSwl6U0Bsb0Xdpou2Cfj
710spt1PYwHOQ40uq2SV6gvNv/oDWzxSfPCNgth/rr4qVhXHulV6L08cS6z7LT+g
WDO9a0qhsrhsyeFn0z36pJ3pTyFiGzuQUKPqeRlIaDJiJsUb6bG6xRQ+1qWl+c1K
zVrQVLGwNBSfGZ+o5sFviJ3AunDqEvz1osbRZA/OzG9c+xr8dOYIrzJEzlb4vy4N
+g0an8NyU3EzIetz7Dgmp8buEoJUp0/8wOQFqrVDbUMfx+IpIQOP8GN6ZVXi9wiw
CLmeTIKVSPofBJ0H9dVPjTqcPh8ShojYSzg0WG+NxUMZCm7DsYhO/EJp2a/MgO04
AOWhbReDh17WrVY/eHa0lGCzUcejtjbCkF8Gx2yiioMZMYkJsYwH2lZoCm/kOUV0
U/VKeEBI4aCI6gXaZRizllDoTlMn9x+/Fs7zPh3SsU70o0JWpi94fECDi983FWnc
UUi7Vg86Ly2zzCeK2wHVno/H4+8qrepbE8kkWeTjAp0W4dkjVTE4/NqhXjSj5n9c
+r1UsbkosPm4cgIMcDiUomgktLp27gR6aa+TpJR/7UvVSGWQDgOI6Zilu+YQn1gp
WjxT8KSbsE0OjikaS36IYHUEBaVBl2NDhWlWvq0FzVLvMVPLab5so/KVdW/kwskv
7sOhWJDetVUdVhIHKd+Lz2Rmmxyw9l/VH/ymTpZPdQNodXc1R7dkXJUuaFvQ9gbP
fQC1/F5oC8AlVMLS8yA0wbFLVc6w+U+BBUv5PS9kdTlnYF+GQC6hVDghNeFyGBie
pKGNoFChdbGGprh2d4+9mRUf8Ym+LJCS2FW4TJlkD8x1Lx7be3C8onDsAz5sUnKt
mnhujdkKoFzIhRo+nS7YW2Nl/cpca8OOlrAsdvlEJoqi2KLgUkkmSYZyVl+aOVi6
qufoC83H49bPfOz0ItkauhyctnNFbpodleaZYC8kawkHDrN9mcptKyUsh/Zyy4xm
yNbEFqIOQ9AyacSyfBJQYfjWH+18YGmQZKjycBx7AC3LKDBqLfzJw90auKfEiO6I
FPO0peJji11yOUIawx8hRkxNFJo0+ksGC74Tm0uUgKpvuN12RhdLTfXNxKn9Vmxr
PmRZ3FEW7DdzXGRj5esrVEiCV7ogPx5VZv9NA/UO8NFeLHX9MbafUVhZKhJkUWJb
0POThMKCObLeKGGJWuLIfpkPCtvoKX2FJPeqPsIg+Yy8Nj8baGVite2VYBfO6FZJ
WFwHg80U9TKKeIddDZ7cYXAT6tvc3qnqrr7f2CfE14fnBktzCL+vgPfG9ufE8469
RAXcbKHUAyHJnNUdZR6tNiXgYQeHDqWhOdtib74uRVGGQ6Al/kpc3nlwp6ljbVxY
BlRgjpblgmLUcMPJq37zbPY4IxKYPW8CrGTS42VkzzGvT1JVvqE6SiLZ5upsoAC2
hAugghTqb+rSwuY0dv+U2iwdOBaMBxNzY3jQKfKFOrGpGx+9Z4HFxyVgS086ct6U
gouDIERo0NOXfpIEw7BsZG+XVnBTA+4hIqeI5A+r3DFLy948PKAoj1PZn5dmSn8O
zYpEd+QeLX8LMaLlWhD5LpR7rC0BtQwdiMoYVR+/ObK7TrAqrpWk3Wqbh+i7ekjd
nEP65WJ9apZt0f3exUh568qpz6aKBssBpt5zFL7nlQ5wJxsb4mcFkWowomsEq3cp
VbyM8KRPnOMpi1SlI2AZR/LdoyvJztxzHRMUjAVZE4C54nKYblaebgjljLMqvrtQ
sG8oYc2z11yjyFgHNkOIU+wJCGy7gun6nGR8Gy55Rkp6IY9i+LIhFANVw0TNhRtD
osHrc2sUFO5TQ0FvPOzKVQPWxZZ3LH8MYBQ6XGZ0uIA/GQvbNknW4Tm2K+gkmHfr
KuHJPxa+l+SiBf3MqEvoaLLa2LeJh0tL3A/+AHwDXoKFiILC9Z+kvZFBPKOXlbjp
NZ2CWMMLuj8mWUpU+Knyxa3FRLLeTl9klLuDdWo/Mrr2crVzYE9FxBCezbdvs1iS
UZaii10PLKGRI7p89POYk9Q+G8ztSK2S+KGHNuxvBco+iGXeFfM4vVtVNYXS/580
BCH37MZgAlZL1J7SltuUmllOHRU/s/fZyy7qQRLd9SEJnhUZXkkGBfz970EbESmS
Q7OueuJZi7QRZ5RpdcMKi0sGKH22IIL4d0N/fYQfk3RTTK4iTqyytaE7WBvH24f/
eFg7zZwoODyfnK3qbw/CPNZU8W9nNHEEGzc0cdR5rzBhdHFelSD9g0ANWUmxPGwA
Yya1iT42mZ8tSpfLx4s7HkeKpjSa3U7MRr8jgeiWRJ+/GOL3/odG/VBpAa07nFOY
sgC+68t0Oh4gjfap/Bxr1YjhZEn1ujmrqCCQJKWLKaAUsoI3F8lCJmUv84BeyTYs
+NcZ8BZ9282IfUU2/KCt8rEKJkn0KEvFUIFGt7/Qp2epUe3vZh61Ph7vMq8w+CA7
4CFAIklC0NTLBl1OfXHFiQvxgNtXUkUqpKeNp4xI8oj2ptYHKGLOUemqBJAyyYbt
KtwynNk1n/TMcZjIhtT6rUBaZk9sL5nbScVdhbvYDbGu7Awb2wIPsZL681DC9EUY
04X7mlmFuOLX/nVAek1mIIVT8huHoA/VBdj9ITaZwiuHap1WiGU6Kx+I+Px/+6F6
ZekD8zDrE6kGQ8fvjK8RzDKnwi9vZs83P5QMzhnZd5RLMKYGf/pdDASkUIsOzQYE
HCpUhqgoLvmJfLmW3PC3bmGM4u0buto7TrXFbsSOsO8g/b5XOLxcbGIADz0ywuRs
9QuU/ee1oOmdmWvmQSm0QcuZ/OSe/9PUxuZR44mCKrj4xWJ7TOZE06heRovQc/K1
tibrR710S+DdcTV1ISl/a0gn77ELNZEOlc7k6/DsoRNjbB9baUtIrAxteMsCLvAG
oyrTz9oWhLwpsCmEEwxCAXwozKx2mKUrRPtPXMlPFiDyuXcPb3wF3atQ0FwkSiHz
Ov2F1dou/dIloS0D7t+PXVpGDFIMcMUEkkl/JRw/w/118i6da/ZNuis1OOZwXnTq
KRarsGboLOOivcH5K9kwJJ5Pp4m8JMsQgk0OK6GmGJbCHWerK9OSCOAXQjBoiF70
5IER3P2FRvCEBC5AorsIz0vVOVbVqdl4+L4PE9uBF8b7Og27THD+PLvPGaBZMeCG
HEX8x8Gqm6kb3WYHs0f+gf4nxQELp6W6AC59BKy7szslF0ugBvM/cNhNXFAcyi/1
pVcLH4hAkbAYEHNf/dxA//EDhX4hr8/5mrnCIiR/398+oet5g24hdOvCKt5m0EQ/
zNEDa3kNlaaKJg8svqYqhZ/zyv+v40WmLEsuWpVnrSqZEnzx9dhpSG2txgKpFax/
MK32RZqADrpBJUbCanFc9fb2dmFgiEIZx3Npd/bOcHo09Ov/4iMJR/sVfPoOYRc+
vy9t1GRQXvjuzFq52YZ6NAt4AxiBs4mcOuwvP8P2xiRC18i8+PBcok88oPvCVeWp
m2CdiahvTrJepzc0z52NSJlpCQAJfClFbyVj6LzdC1sRfkd7Rc0/pSla1mqnNCyj
TPzm65mZIYS4VhmeyhUTjdiODj5jPO22gHNzAvyTBGCz9F/hhabgNKEtpfDRXpRw
NW1TqtXPKrf5UEO0a6Qtl+fx30P6BN+YrvBz/PmkwM7wRDkbIoNqJ6zWcjOgjIop
H4FdUbiz0rH4CwKspQ+T9lWMSLYKCO0SPPDr4nQDNvE8VAG62P9NDXwFe5Tyi5qt
HR1Nmm+PL8avZlm1BoeNdMxTnsRmfpb+YueZ+K4uIJx3AODljuNN0fhNyuHqhVR2
+P0VW8jwgJ2BZBJCcUjNpAK2o/GET/OjlNbD2ix59RzKv/lOJTyZf0BWPa+0Wv/T
c4sCMsxDRdZR/xIUKEFzTfNRw7IheTETlPbojOE0rFiV+nKm4/aoAbeK0A5np2ZX
1+Ic8BjbEDgH6fKwfs6BCdjZkrkgwDqnrASHb+se0kmC1QQQGKH8P9K1u94WIw0L
mG1zATzW9voE5RX5eh23qo8zwGrC2+sF6PxYf0b+xTUfM30Bxj1MprOW2zWMUrey
5PN8sywEUTXsN9qqeAK+y8jMQd17FtpWt/lF1J03HutO+wCLnjNSK6Q57tFyaahy
tJ5i5SuXX6flFQk8QlQZ4aRDJaFIrdFe6Efwefu6ovx/iTyoF6lZiBDme0dZJr6o
qNRI60u1FmXhAPBzeF5mO3EzqxpD6piGlHTyGX4R363h/FtMSV2ZzMiyi/SQd8DU
BA+DU7soYRQ+DZjMy+9TDQYv4ync1As2znb9sakBO4uhR+ALq/1vpKBDGvpN25/y
NZoL6EIKwrTaoUF58rwUmDnffuxxtoLR3Jd93l5ch+EBnSaSnmBxrk+w7tykOSmO
RjqBjja9dPu6YFJnORshLvC/lGKr9Wv/3/0pzD87bW2/Orv3a316x4QculzvP9st
uEVyeFAvH0YjzXze8jG/yjuBBco0VwHkYBfIWQa/8gIVN4gNZV/OwsnFTvBvxYGG
MwPyM1PsmKrCwAmGMzOzLcmebudw/PGA41W+mo9IBRQRh5mKSEqgIlgYTGM0eozx
nbR+AU3ycN2T+M4KXKj9vzNaB5j9I0+tp45IUur4TEiRmaxd0MEnn7tr/2sAw67n
qzRHi0P1CAPp0T6GA4DqQWNnBLMF+eXzuRZ9UJJPpXoudfxqPOkmOEGjouy83JXx
24ZXjBr3c/W40NZbRDgN5SuRYNqPZmVpKcsAt0lV0fctFpDs0eI8JG6kuA9s2mXb
8JRHUl1AF1hiY5jIEL9ouAyk2VSgBOOjMUJkw8JMo2//PJDTY0l21EVGVTayf5AB
p/aUSPQgJxxBzOg+XBW3+Kb2sbit3hx4rBVPjqkxWdtYszQlDSfgHOTAl81JM+Ld
xYmrDM3b8fYta0EvXvecWNLAiO5nf3/xVFS0prlAbyf3urKUeoWjWnnTO1IGEKQD
sH6wh5x3KtT6rF3NbYpa6qBcOjDZcBh435i10LRCI685H50ZeQ4ZIpXFmzEPqpyV
UaCZjxysg5Zx+Phkinb6rkSAUTUr/cjQbQNPUZeo07D13IEc2rzjqIkAgsnTFA9p
CTwJHYtjq9te6Cx/Wa3y5wxHenDke60frvn4Od5D6qfN1rmRmmACLEfaaYo4I5tD
VPyJD/oznlen96zDqXZ2u9Ka+GKsq6TByPZCpXrgGS0fLIo8EFApA+37U655kQjM
UkRO8NwwlxQ0yvqQMBzNamC4n3Jb2QOjOHsL13O1cUA6y4uIUF7CmSID40y9gp6t
HVl//D/yOJS5jGHCxqzgsf+yBR24ksjF39I5Fy36PPuPrVoPZcV7JiBL4bNE75oY
nE9Laqx9uN67dnBR21kXSNtgxfx0jAg5SEHscrQkQx89bK3dDuNUsJb0g46WHKmt
1+XYRrS8IiA4GKycxAFv79iqHUG36tig+ahfAzoRyF8QTvsSo6ZQj8IxuFH88miR
2yAJzz7D4k1GhIGq6yi2wP0o8Uu10K7QKKtSuB6wCZ9R/LQy+E46tq/hxg6OQFJm
Mgn3V8lOykBqwG5qpk+5ySNi3W+Vg6+ZdoklBt9VfBcqfVbjiPXEQajEm2jBcEkk
x9VLX6hArqe3Gqr355NPhskyTMdVguF/P/fRePaFpl/npV1y9Q/Ak21gc50g7Vfq
Ws13zkVlsjArYKMWoTaenj1jE86A4wl62O9XZrJxEIzPEig4NFFBeDNtZkfcHKn1
IzA85Q0V8LCJRdsJtvS4j2ko1P+bYMoxaioJvFX5kiWABgUCP0VZT+gtGwDuDkVp
5QW/DnGYTB+TaCXpyQTx5ptPO/C1rboQju0NDhJtMD8atsN4NLA3h/K2oJqvduuU
KtyxNXrGvCFQfwmcBD2o6VaDZ8JphgSNqVEN0IPIHtqtGCGBM1tS+9dmwKXiRUVC
6cX2ALzg3A1kvNtuCgJkbiPQzys35lIKgPC9xOLkdS2iBWjzVmK+Hax83eOWEFZM
vjsxXfjwG6NIYPRWuNf00oaLudhMdbXB9XCAYx3ZBMF7mkCofMQ/Op0b+m6NI4u1
wysxVFXAfyS+OF1NIEO97dGYMzx+PJOicSEeXH8KKNn+1zbAzLNdIprKOlRFELOx
URh2XzXjE2i9C1zgHM1s24GrKeBQDo8akuAf8MCfScXF8v48iy9p6DyJmMCx0wy6
RBk5k3KYddqYsbXk68+d/MIf5V/WuyFwD3O3kdXXbOOVc9nEj6/fJjygDSW/7aeA
FZ3SCeiCeX4F8L3lv+O1C+cNwbhjyZFWXOCNDdv6Uv3pQbeYu8LO+YXaXrOiqlQa
u4NoKnTa70GOOcoB0Qsb/IaPwdjRBjRZQIStOVubV9rUC9fIbGPw9yUBvj6sNRBO
MuK+P9/1MubpYhv29Q4WUlXhtq0J1tSfI18zUJnJvID5bdjAFOQT0LnsW15i5TuK
Ez0FFYcH9MlHwjltLDQTuHDhGd66LTac69uEEM9XbQhm7Ci5dJcIkltTCMSp+slz
98HXd1JIYleWqeybIWcIJ7XTZGUqGKNEeVwFfRWQ+wH+rjDZAcox13KN53WZndoA
GyyXiFVGbo6UfLOv6IY94CT1JMkxRP3moWpPfZY9xBQt/vbB/wsTsfWRu+SnhHsS
yzMml5tOasQlNfLAQ6dk7eXtEIjDK9QaeWnys/Sn1ZkLu/FAQWHKihHEA6xlTfd9
Mfc00dv+BKx2BATU5jUbkog7nQUDUZKdzE1BP0PyRz3fSR+cI/xKitNYDs/B8kEp
xWlEgLgTnusXZHvPr9/K1/NcATATPVEp21AKTw7T1FrqJ7SsLIR5sDnmhV5+bEqj
snyXZcXG/EDH/by+6hUW6uyNU2i6YxjKB+vLJQxtcxHzoGU0M7hF1hPnH7AUx1XN
ZW9ci/RHDkz8WITVb+6O0+UEU1ztprazUxO6nOuZuLjDe3E5rVSuMndORdINSQaz
4qSd8EWKt/O6n9wgKKJQ9b9oEm+m8u0U6mPyEMdXhAlpHVb1kDdsu4cd/hyI9RK8
yhKWOmj4rV6kafXuka855CmP11uaTmGWunb375mXNfekN8K/5AUihLouTj7mpifv
G1ffNVVQuaMa6EBzJfrB9yFZIpnBtYvinmiZxi8SHXrsMOO0iqp/3ntNvfEdVGJ3
2zVvJ15TRFvFEAgTlgGBoYTh1anaPseTcQAg1f5SngOT2iErnBt4KpQF7HQtHQDB
BndOa7qsbLjqn2bGJVh0fRwBjiwEXGkvnQCSiRUFuV6k3sh0T/PYaIVuMSYnhi/0
BU5E1g6J5VYOHl+5yFhfyT7af5nbGp7ZpQNYFo6drm/kRdTMs0WfiiU9ArHXPrFO
G0tlDNjxfrse25FYlGYOpcwvy6iasjKSS0QRbsT5xphJqQIs7pXuPRjvNMpZJv0R
LTibItzLf2uVwtgfuGUoxPY5lUfL8hwVfEzXkqG9X6S8VRnRIw+kbs+5kIDWM1lq
js0sAQRxuKi86YF0W/x8SK3Bx8vE3sqt+weE5/Autzu4nzCyPsO4Hr5XW+P2e7cX
EF1jigcEs2/fKOK1RfzHeAxxtHIcK5JdHaBJOpynzgfbKhqvf2dmmT3xYxfzwP1E
sZ3NwJXnoNMUaCaYXYG7/jzj/ze+yzYKalmRn5FGqj5ze/51bExDDhP5glbaHVZd
eCCR0RAXdzr8m23+Yi80QDRLIZgartSYSUTNtzFjD+RPYNOYmW2Pn+kMp3njm9Rz
k2ydiSwditAM0M1MVrag/JpnFtr/8/sdaVOs7Zkw8CRKxEt4165HB9nVpYkCENdv
1LAbZqbEhmwoGdNKZ+dwN/besv5wDd6AzHJgayJmLBEs+Ndg1lcrTknoCCuaFAwn
jWThLmwHei7f/Wshr+lECPo9IlYxyBtvHRGL3carkOSW3ljpPLHvaho+GRpLp7gM
PNdlD8cZqTn68Nmz6cIFmcXJ5rHzuI1SSK3ux3ZT7aW+idn03t+BzEyXvZ/mpqPW
xU38eKzbIUU+MSV3d8Viiyo+tiiGKbNfZFvMpGe8N7t+17PKFtN9550bhVx2fjuq
HzFCFxUiz4KbDmqJzWWGdBMYcjmkNYMwrNluI+NfHYukoZ5dQqEnEOR0Kwm/R7F2
k3FBwiVOLEGolN1KlvTveC6xfo3EyVP0CnC2KxlgrM7alJ5lfX4Vw6l8cM2XhyzK
02kUvHb0N7XPmLgk7FdnV/qO9wGz1IBzgj5tWDXx9S/w/cAlfk0jDBz5JXKXBt1t
baY60LonfmJAdFutj/6XuXAsHcanHd4LiBVeYcIxZhOoeem9YDzb859pIC/4yXu/
aKXa/GJPBGgeJqS9GJdzFjjLHQiTlqfE5mQB48hAg6+qfzhDoNymnlhBNW+plXat
75cNXxhyaOfw0kuoVEEoufB0JuiB1M0mfuR4ZnlMXO1QPC3AJD9OcSBJDbUn4tOC
tcZiVOfL4YDQKak4NI3tZ5VzwIwvx+iD7g0JTXXrM7bl5WodYffWvNWZiuwkFQlg
YDW9hAXVXPhdtVqQRGZJSD4uII8wR8iWKQC3x4oWKANlficLlQhEEH7+ueNdyVRC
ZdDXhl1KdwDSRuFQca+LXTLd4AjJy1MJ32a++z/XKlZhvE/9hGP6D6Xfu3ssN5QV
s09uByv3BUpzLDD9Deh4pCi+G2Xxwp9VZ5ZGEaucXLKkBH9LStgXH0O3bOiinTBS
y8tYlfkxH/OnXY/15bqEgXs1KDJc6pP2Ih3B8Ab8R4l62T94eGBBub/ZZl1pBiHS
U4KVDI4d53av762PutS2XH7pv9sH2LkEFSK0HLG2sG55nzPTe+0uJvQe3IXgGMVt
c4q3UjqWzGcrQh2LoxB6lZA5nN37zoG1ORGhZ6Rh/uE9X29c6UMgS2AZhTTgnczM
eKh6TXNveGHfDU3mkx5qpw7pl2U9UcDkJ9w2GFNv5rBbDiw+oYeGdnAlbdQdUZZN
S2h/KYC5U/p7P6xdubIeOQIsByW5cifPcMcrtkTvpCB/8N0gL4D/GmsPO6jjWyjI
E1jUtyKqDS2Qft50Nvg0UJmmPH67lolpkxg5I6lHHYLl5bok7mhe89NHsg1WEBLF
4E8ns3Lt5k68BdJYMHtfOijsH5+7kot96eQZm972ZZCSoeIeKCvyz/SM2hqpzy/C
6v3OZyHZ29CiFl83gTM0diqc4namE1Vs7wZ/vEfyRhwEYt1771I9W3yRCW+JbnH8
d5H7HMkT1ivOYr7br4TIY3xjh11UWX0MJ3xXZMdNz2leCTjS8OupiANBfDyMoiN4
zyQb5fFRjuJ0IcyFTEzn8yZNz9IPqdtxKUJ+7PWVmqMxXQbobINL72hLlUXceJ4q
oUhLwaRlPe+XUuGgqBR2WtoeVGJVGxXix6RRgsE9ga0tSV8dctjFSZ8/T0dmUCPD
FJ2l9MF9Vw3hydH+NteYSkrmNO0acDPxuUYlUqRVSQqalUQzG9N/B8g+b2eS5AF8
Mo0wm2dmy9bwb5xQhgUY+ztVgDUJ3CPMJLDGhYOqHnUZ6JbwXytiGI5Nl35ZYE3Q
lJ5Fn8iN8ytidwUV6KSzU4Uc8JC5vYQ+/28a3OEmxDpLK+Ixbq9xU2W8E4QvVw8O
JK4N65wvWebza5OfINWbG/4JKEpMs5NCDHXwpCvWbzqqK1IjarGJHzq9cieyt+vQ
6IHeMeriiUPZPK5u56U1ZMvMHocXMZnGvD+E00Uf7rkwJiBkrJxxEb3b8obF4YuL
kkfCDSxwVa3TiznWLgS2EXO4U6ftNoy4vZn/2KHSA2ALSc0fg1DvdTrhwQyB0af1
YuYi0E3fqcUo0tZMRqpemA4mndfRpdNhUKOwVt7l6g/4TPqkPCi1CVGoLmSx4c3z
D9gCRoxuOzIK+jvjZJ6NnmaEAOYiUxRsucfKB3f2hObaTtsAmjhKC7sUMjosfeAx
bbNf9UZVBqwDVmJb8IzIv6Vs7bmomVsgRYuOB5ZKYo9kU50udx+1VbmQv6HtDZE3
FgoImEi8MDZpP1iS0nkNbdnzMHLjQEYBQr+Vu4k0QBYrE4m63peJGg0UgKN0LPi0
XBNRjKDYwWtAjSEZ91h/ke88/lugEwalXhOcnUSSK2Nc2eXXXzmEmbN5TWnZGkeG
+icvaUAVhqYM7gjMBEYblVUFOX7mUHYQEwnn2nIJcAGiGam0j4CfsFfSB0M2d8ZY
wFF16FF5nX7OVhKF6wq3xiAhHrF7REx0CYPg+QOj2kN/CQcFXXYNW/npJsK81Ay9
dcb/dQgbRQbVSwR/wDBrgLP6TdNXDEhiTcAN3tKMeD2lm11GF3jDkoKIbQK6ykYE
6j+FabCfjI/29SMr3Lg5zmEGrM95jMxOBxqBNg90AA/lc9P+9LBj+fKEWr2rS8HF
RKUA+XqONLrqyHdNhI3n3QPw7jjWrq4DmIz+uBVgMI20cvYjs3GCmH+3+4PTUm7S
NpezBYkTc4qHoxb7s4wl9jQcx27s7lihE7cKw+FBbxFRwGU85YNIU4dbdHbFdt6h
lRNJP7c5suCQ+Ge6SbDvxjSjsvt5hwBKBw153zpGpX3Zx3uACbJo5/RPAceBWTmh
7h+lCyej9vLPHMXpfCxx1X0S+Nkiz2M4WRywE8Z9QWJSLlmNJVN7Vu1H3AJ2xVQn
fhILKAxpwW2+9sVvE+lHBBr0HAhU7h428vg3GUi0VEJI7w4VHeQew/iX4dR5BLi5
0DmGSO3osdhXeLxCn6ZpBTQgzh+LLQlG6Ge8lIdUv1jKlFg9oWkvr2yu4XW0QHC7
Vh1y4nE6oe3eyWxs+IOfXMzMQoHg/qur60a0vm9kjJi0HRJzKs0KFBn6rA5QyR52
fIaygkgI+tFsC9IAxXZFPR7zGBUiqPfxzS2UkF7kbjjllsHNe0jGLdX8R+sTWRrY
gqBTde6ZxZe40ZP6OziMqnFg8djZUHrNFOSK1Bd1AtP3UrhEx4BWWSn98DVhcjoD
vGAK5XrRGM6u/o+dotAILy0gJqLj/cwcnTCRWLcDlLeptuDDWj9UGfxKURJf1p9D
2q32YJXQe8jubWqVLEc01ZWmt01UjYhDZLpzF9SbldNkeZYj2H5iLafeS0ZkGNo7
t74tENKCpcmKJz5iKTwKSH9jwwqXO7nf7kwhENNpgzy+kzQcREnPkUkZk5yNMGD1
rIp2q41G0QnlulHZMSX/H60CSyLbWYIbI5HXY0qYgYEw53hSDDGaTdUPDWSjcjdb
5nxpqfKsU//FgY5nC7TGmi2dywlWepDirBLa8+3qW6nvXxnpvnGhAnCtzTLtnCK3
gdNQ9xlRIfeXw5dJoSoui6vmkC+KtdAIKvXsT/s03aZkWy6/lk6vfUv6qiEfQbNz
Ia6RXDfTEkEozCLAPtkGxrBkrZE+BgvchW6Ld9bKbo3ndbuks/q1/PeVxjb/sM6r
I4CleuDa7Loyh53eg7hQCLMRJVJCK/mKCRrpyuizszBW5sqSew8k5ap9epJe/u+0
FE58tu0UMvO/Ekh6NKmpkwyNd6EuL7LokJlunjgjidbuWVnLzcDmg6J3+PJSYZum
8Zrnd/K6NnJY184s1oFU/MYuTNAsFjpYjOLTcMIIrrAmwAgcfjCn7ib/HKNYgkc9
N68QtfQu7FCDVyIuf5c+jhb07S09RpFMDtMo6Cv4DJNYMvLQMVcKnXjWbqvUJWs4
+u+r6H+zzHqtCFZOmAuCYsANgUIvji+5AsU8pzJQOan1FWNFTWJjwgP39gkTZHe6
v4Ou1Xtc3yYumYqWJa+REYkDlklPj96N2dGXuyRYEoeGFDUbGHo37d5hk2MCce9L
WtcopkRyEgsx3x6/mqfMc5UbKpwBgxk0Cc7lFv0cL/7yreR+pld1Upp/L3Um2lGW
tJhJlP3o9AhYvaIfiOHN9SRfBkQefi5y7bSxjQCviRJJMBi639FLcckosj+En2oQ
kp8nai/Bf/Yc7W3y2iRs3FjAx4B1VnAnAZ+TOiLvi+nXYcSyATMVHmGN40QyBiW/
hwOEf0xmJO+eSBLXN8zvdHgCUoUf96BPfeP7/QnMeU00Z9EWTvhNNpZOnL/HIarr
L8d9S/vp0EQIuUsxeazMBM+LcuXqe0xwS1YKuUOkYnhLFauPjQUR578lxvIXmcVI
f8nna0k19lKECNe05mJmbkg4WAdM9E21kzMqYB5ycdUov2BUzlVzLWWi2GHBt2uz
jF2z4T8Qi+q9qkjKHBs+qqG53z5VXN8CRRx6W3KWT05FOMhzY68Vzz/71O6NkbKM
qz74FQv04bljjU4h4Xc+jT1fGSjJO0nPIuTnjgEFmVTWWlgi2nbKhBWbSva2cyE/
V6cuVg9i1SLRkF1htKzjtexqTlFfIALKAxw+ylRgETE/Rbyv3/qmcHqlPTHl6h3q
9RWkieFf9g6fh35kDAvRbf5/1LoZRBWRotOkjoYMGMqUKZk1S8PVSjyuc3rE7o4J
rh9wy0mHSyuaSwMGvkPwZi/BYfCEWxwYb4TW0guQoKT1PAHpaGXd2lmNJ/cw014m
WLLjMjAkbYLm7EsP/jU/OMfeUMx/2/o0eYNoBCXYPkg+ECF8qqzLhf/VC/4w0Vc/
ntBeBSYw2cYHiw3Do4MKplo59A8AZ314bQ/Gh5BHfKGla0ayGrOZh7iRt1Sx6Mjh
4KEuf1g9qjmkIITl4WSYUJOGaP85Snqo9IgRj9QfnDJFSlPo8JpVR/COvXIFTbua
ccn5Eib2vbbTkARiVh6RPmdlUS1ozoyyKdGdMjnhfqemTFT4baz9+ujTYsNxX3yi
USttnF8QLL8xDAdBzu93Jj8zRcK7nqEVJgkKheNM4skT/R+s7XKIGSAPLSPg2yj8
tJqrGb7lOGLSU48q7aEJNQpy7Qu0mW2IpNXXl6eo/LB7zdCSJqdhCabUtubpY/+n
XSx37QB0nssEawUeiX5L8jGhhUOl7dNko9kPr5QK4ofKEC9W8YgJyScnAzD/C34E
6s+OgPgIfcbw0K3KqksdqVIEMYWP0zqk23E4R8Y4FF6J20St99EGuAbrgS0ME2Tm
wik7zaxtR+40L5U34fjQtXsWQlNanMbUUTOyLWrqrOyETM8NPqURV1FMGaKXfjz1
ygotoB2aWEScZCM44P7YDF7yygbV2bRIhZ7LQEZvtCMh/5+hCdn67cVWALeKz0iE
KMys3AfSmd2EejsSoPkszRrIPP34C1rcCdl6pPW/kZH6MMXYuGkykELt4R+zW+U0
ZvFPMBLeIcXB3fpSOzxknXhSO7VP91TdqkHhIEJdSdqj07dqOUb48PhOkGg56/yl
kyl/9oD28QXPQTzlNLD8/N/Vw1Pp+dxRlUJZ/wt8afhZ+NnfRZ2vq94y+D0VB3ri
3LmE4h8fJox/1NDSpB/1bAOxzDm4aX+hIq0c1+hCGmv43Q+J5rxaJ9420IIHQb9k
eECeZiaQ/F90JA8MT4zGdJqUFo/qh/KgnvTRX7V569G9P5VPZjWambrWbKTVorED
ROKITwDVrh4EFuCj9kin5cVKfDkV4d3/jl4f2wXx8i2vjYHm69CWbn7GpfOWaTov
LqXnvKSOc1wDnbFFYn9o2UEFbmdDwf1blfYcfvp/oAlnSYNymJoQA+yGhVC2LEz7
pr+9kwqfIKnkeJ2M4ep7Rhqij2tkIl1biPO5qaefn06wIDgixJ0qZvw1fmUvIQAl
gXfybtP+1dWIUIUt//EUG7W2X/+zD0oyOPAR51Y/3fTTLPZTlyO15eJzZoeMHh5j
ckoyln3K66IlJwxgwO1fUIq6gbXu7aFW608yRB1SCdVQLv9+qXwGw27oUscirnwP
wBfKLcLJgGofGzNYf1DlFhKnKDPf6EfRjOIxVMN+jofIfUdTvO7yf5Cct+LfWig8
0BDtbcmeoNU+elWpsMoZrACvpThBZbnTw63nM4lZ4APX8QBx0B82mZnFi1wYgFtX
1j/lG3nnCV4Zqz++vdjCR0I9Y+q/DYihFSA2lHxT0NeKz5R3JHV4HZP4DnnhlSYG
/Vqe6W/+ZCFhcWtNzN/yA6+nvVW6DDoaObQBOAEsfVAhiGqgMV7d8bXNJGLprnUL
xnOSiqKCd53EebsC2Dw/s1ZzV3fQrqju5y/XEM8kY8B0S6wdywQueQFoKV3VBes9
qOSUVqmkjixF3hpsT9xNkQ5N4X7JnAGfpVzkP4SyId+WFagqHttqTckUraU6oy1s
Cuv+2B9NZJV1nqNUOTmZ/2WyKWmMCJ8rfmiEHLu5qEdM7WVlw/yEx6m6BHLCDfju
Wafzhz+41Nos/bsIf3M1Vr4rN63h5QAhW4H6n9NJIXp674SpVVGR7WZzQCgL2Lkv
LQWCIu/x9YbrLPbX8gQcoBLxzq7cFIqDjhZLRSw1aso+XflimXo0gqFskW6sBc1m
Z4/TyPXzhNJXWDZmGQAv5WDLyVFWvQKqVuGyjIIAZ9oQW3iu1c7skr97S5ZIgPYD
qJ1ebPRWU6yRK1ps26VL1aA1TmVuxEyPcgfrvnXEOQl/LOYLAVZyL06OJIyUHOSl
E51P+6/888FrDU07lCc92KWuMwHhgGOVYrTWA2TFbXDFq+Htz7kiyoyym8cgzv8X
DtZBe09FtXkCRh53TACqagor/C6bzeJC617aH3QsOkXq08mKmzoI+kbdvNNnjbBy
3OYDhowG2QUBcO12jPbyDKtGpKb8RkG8eklmK6P8A+PTKED87Y5FQ1Gkfds2wmSw
aweALRMts6iJqDIl0xm5Nrd/rW/CkHpuLDgmf1QJcJsfr6LbodfAZUfeU227blq/
3XdgCXqMz4PLTHk9Nt0Do16RJ/sa/wVlqpc7y/HXu0vFJDd/ckwVaOjdAH8E7PG9
+FCqYID8g2yHbTwE5VY/J6pYoUIxDPfBLB315l2fe4fvGRiUpjNKG1xucGWj2/js
mAajgYZ8OfOecK7PP5gMpF6EJ71ciAeIyRd52alPI6H5/A5uda5pngXFxBibiv1l
9cGa6fKj+Xp9WxBI86uTgOQA1AZfZrke/dPzEDGAfh40CT9KaMTcnzQh1S4CEqUc
Mgo6zR//P00/+q6EfBRNFnWa60naAKMNY5grLkFwXdSNibJjy8snClw1c2btuj3q
H88jnsEEhCBQUULZRgdZOK2+ZLSjeGUgdikX3js95p/FvRVkUyLU1Dbeaw7h7ty+
QflNgxTMYnTuXrUv6k1unG0GqV9hXmuTvdt3lseSbyK80vU4xh0tdXauFbrC0ICF
8Q3tRSPTgrpsBVEMaYwczeyC2jBhKVboz+a7SROZDQkwg2l5nDsyT9Swg0V9zaq8
Z4x+jC/QfFwFxsi66yKlogEvY9XMBxXkqAVWmQ+eph1kdXiHa6Kpfut5JQWWTqef
RwEM83PPTX+cCltvpcKE9C3JBDwf9uvFuQ3yEx5oNs8pBXS51Yy6QnroKoFrsRxE
bCKCC/rPjuyTc2984RW1HJxC2Mj0Lt581XzhYHnpo2zmzALCzp1vQdLV89lzpN5v
DJaieZml1Qll5Cjlte+QK6eTrb2Gl3ei7yFOGZoDe0UJcqhysJoe8WsuSRvUKg/c
nBvSauQ7EQuYoXgJJppQU4mqz306ZYFx7Yw/c7riMDgEDTXLqS4UtZMDgAqtX118
dTRrllpQU5JgFruPmJ+e93gq8Ejp+ftsiZL1bQuvhSU91vzumL19GomQ5ZHDjyez
SLOswIzzvTj7ui4QahrJaIZsdqiBELztdI9Kq/HySDd1KLprihFJYOiOj+p1jQss
zJVwg0FE1NkUTIk2VJJSMGV4SBfbO23ZG+cdq/xu0zmR99wxDYp0B/nicriqu5Il
D8wKh50CldmpIEOayn6ZJpUih5GKseecxkoZYt7yzfx8BGu9ZfsmBMM2zHw/mrhB
Kfimt4oxHew1g5+ITZv74R6NVoi0IgYfpk0mRA+hG/7DVVglhUsgApAWnpWLcH9z
wPcpeDVZqAH69wIPFXtJiZpSAHXouwT1tGq5RgWXFI30rHZWJZpdxMedT3EUEc/7
8JG9XUKR9OqILyJ4wpLSfBT+dt5y8oTXDNoxn9z8NeuUPLIYixviCt5dxrpZhL1G
N5vwDdavVIVH2OIygL61elagOFS2eknxUfs9ncQxChLr5sp4awTN08AknW91iBEH
uT6TADonAmKfzcowJ9wHy2A6QVxXoj86UTPpXJuO8ET/GZeWo46Ur4jWadNU77ar
7o2Wq4oc0Q0Jo7kdE9HjyVz5mNdmlApS6t2Yg84qZtfYad5h3MdDBM3TK1FvOnYc
H24RA2TysSSoEb8aOsd7SFEurUAA9PRb5TYZrJExHW+fuMqnfYsjN/5u3tuuh/7m
E8uhyBgjMgePN6/T1Mjv/nUs06GKKEahViTzLcfA0uaK9DRGJrCaNh/psQdUoMWR
TM0+U3RllN5oXKb1G8jQbPfLRsec7XAs4DJfU/nKTvSbbUDYi1r23AGcrTmnuL7i
4w2+oWxrcHgUPipF44SLOIR8qQwEWejk31RHWMSBw85xxqC1gS8PTSsZYakryluN
AlJmwDyBRuNyb8yMg4NrEsFLGmIi13UdtKOond225bSityfMuqqocAJMk/u7pWsE
WA5I19M+PYI4/eNOgYhkSpT8mO6d5oX+FVhL7uG8h7vZJYWbGwhWqjv3JSdEEZad
eMNpFrZqwX5EfFC2Bq4W6vF/q9QFU1C5iJQIFEsJc+oqhimE6E1Ei524kJ4PYw/+
BLUjnvs9+oBBilQirSL7q+E4YumT4MHxDaS23h/3+V0QYcxqeH0wW588/EckO43F
1o2rphonXpq/bSO6kHIX6gS3MtmWuwWDQs0kjyc4CKkht0k9UbeSjIMS2ATRfcYk
+YbnHMjCDbwt/kFc6Yn0IaITSVVThotVLgqvQ1NiBeRYrtxNiowcnmJWdX6hhAUH
3BGMxsdK1JKTQ8YnWq4uEl3aqrI7ssEgSiYJkBK55m7WMUs6ltrUFBvIo+TTDXyF
xasG6LEmnvnTWteTt0XM54+MdRJ379Ct7fSOI3dPaGGjhgzmHfMXLf54OF8abimH
8PF44odTJ0yVHrrRMUVcPc9qxkWvSOb2VJlcqJPCF+6RMZMpPI9E3W+5xCEw1rkH
XkUuMFj2+HSOoNp7BA+FEfe5b0ZZfuNrcWtqfGDfcn1JNqxFhSCGt1r0sCi6wEFs
GHm6IkNoQ4A3QhThMjr3kjStFqLFDPDase2t+sfe94ob0AaRAtD0rmHiNxm8yUP+
zd+0sbSXi/iPcJjqiru2EAp2bdE0X5q96wNb2xVhnNbrVu9Xaw8mHhOxssASiCbh
s4bjqr29c8+6ouFcNSbmnWypT3zDS+9XVTknDEHbqttsSraKB8gCEG/wEdPQ1+Up
MH5q/dBIpJGTD9doEfJ9RcKiljWktta+aKajT2Lz0itImGrieFL9IL8yKMu1a49O
WstT0Fhw7mMUptsNq9GPrcP/5KNXJNu9gIlA4paj3TwqQHdKunAY9y30QnXY9dNQ
/UMkvFnxcLhpRWwwxFyDdUmO4mq/KoNjSNsFmL3d/0oDlhpsDqV+PV9ZFc6GcWHv
yGISaqX6v8T+ebeh5tRzZ6s7ujKtyifSVGwoJUJWZUJK1YK/j/bcoe47YiBdkw9c
286cCPSNaoTb2fdoSUnVhoPMt5oF49QR1BaE4Ns9x+hFUFiC7GIzwXnlH5lfIIZI
Lk9iXnBUSTr+LANjEMtwySLnUVY46ZDlbAmxSb7Cl8Nu4lHyxxL/LAJY+9Tn7+km
S0NcYpL99RwyZZMJ8OoFOPs3uPiQAbgmf30WGc8xGd+3I2sa6THQEqE1MDS70iMk
HSolPdRZk18u4aGgHEoolwKVRZV6lx/yAz/unt5nSX46dQtSeMXE5XvDGzuyw3Tu
kIhria7//a4qjr5Pezu/n8yxleO80g4HS+MkPr0xUlMe1LKQ03QmYmqniEhv7Jk2
qEBEz6Zd72WtJdIH6Zocz3XlSRCRSbRF3AI8HdW5xP5DIAoz5qMzgMTARVyI2ybh
rIa5ulGSVuhFlKDOdRSd0UZHDle8OCevBpJ3nXgS4AhiheIyvnbScDJMlGaWeJNA
GRQpXfYMCFjwvrSBGE0Lc80b+m1hYzP9y7sEM+hoR2lZw5XHpPdkVFZ5lkRCfNH/
eBYaXmnMP8B3cFHLln83jS9PLP7V5xdKOxry35OTjy6T+VRC+5gC52HpXXnM9IcD
hnLZX4EeM9RIUDHamH0PwxnkjuwQ6RrMTYB4H9j3Xn8vAZWQW+K3LZqbu9GxOccY
rt6vY73NA5ugmoZGX48SaV+VUosyYxTRK+eoFsAaN4VQC0EtDSeG7ohxUEiqg4p6
T6ikWSy6XoOlvtNLTxeU/uaFqycXh9byHi/jmFYYmzSEIsc3/DW5FbOkl0QP5Y6T
See53XtvM73Joe6wMtTPSoyc0zBRAGTtKJLkeQZ2FiOmeW5rfYxfJ7dt/5rjY/ob
x7Qsap/9+UHMl/GyVrDTEhxvGS/A/nRb6VJpHeBWEKQIVANGTBx4s72IAIXmd8jW
ges09fGzWFx8PgrXT/7O5tWXspdY/+BUtg094SXOk2/2t2JIW0Jh9JM0BO25sRBO
Nh/u4Lz7xlKIBHRbnT1qfjgk8Nr5j9Y7fVOmqAJol4JqKTTPgBAv2GzrtqJlfPLH
JQkoBYPhOtkcSomeK8bIj1ST/FaL8Ss5KBv4j+YL9m+zw1Kkvhd5ZhcSiWAiy89w
59Q9YLrX/KEORYXerSU0201Ph9jBKb1v/V+Kof8OJ891Trf4f2y4LaeRl0TUVNfj
zCd6kDLQmvqmUpXhI0esgU4rpcdzqKczXDzoraDubjR/UVDnCs6Eu1uLi3qrJPZg
ReFSRCmBAPLsSLgpb4EyPhZn8iFHi+kahIgJNgcnAgWkH/pgucM+6Pd5FKedjnVq
jH/NguuFdLZl4vY6E5t7gzJyJkc+Q/AOYKzNytNmCY1NLkXnGZttr7A0n4M4RKQs
vIG9HrxVLGcjaQj9rLWkIsKULxyOBIpgXrb7bWEQwBGBMm0lHL6fZcy0mkh6WTPQ
wWaFdU9N+1KIQvJ00tLZCzHaq8G8oLDLf/XDlFuQq9beQlWH5qZBFgA0Uf8T/6C/
uigPaBI/9QlqBQ86bcmnPPPZz5jnfyQoJ3EKm7LxKU9ihpSD66bR03Po1zD0aPrn
jiMqDI6TFw1gtQ8PlmNXPY8n9DNBYs+La4NbNNJ9YcdDctMRBNGQA1Odq7SoW64B
NOdcFO8FnyxsK+j43tqgJFWgc45YKXJqdzOyWpzFvLqUK3uebQ/Kz10lcDWHALAc
4a9BhGD4oLf3vP8xmcwUPNXW9yLrZ+qNbugZj3q+rLc/646swW9f/BVgPGAg9TUg
txpPh3zvEjU8l4o0JobXwmJ3LEKe7M5nY/JHzkpOI6CeMHvlSLy2G5GLqyr7jhNQ
fV7waGyTlvXlRQjyvMqudIDnwOCeALMcbU3CG667Xhakey1k6LOMjK4sHvsgfPYF
AU2078oua78OMHzDl4ihU/rgxGBUUwKR/InIJD+ljHwttJuO6zK0ghE9YRcOR/qE
ymHl5Rq/ONKC1eqDdvrcxujRSqJvrcSxDurKQvbpNdR2unwgu1oxfmG5wRNsQ1Lc
wWTxID1UQa5S2oo6aCR+P+I3Oo7Mkk52qBgm1/lZ9o2Vc+t8ISNm7u1NyoupE8H9
nMxUJAzfEdSwZQOK6jvDOnUJBGuOtII+LmbII0xcHnJJF+B0QhTimwusjIir+djU
RRVydgaCAZU7xr8t8s7AAPbLNt31GqtuBZTuicOZCOixFxdOW2sxd3wtoBQyseoV
E4QJlJITEX58HwK63tevhhIVTCdUgMCBDvXufgSpcZ3YjL6fJDwpc4HrlovG+5K6
ZOL77oGFeVVe6WLBqo6rHW59Ast356kjQ1YN6BgGGKVoDLLI9VnzwArNfyMq6kSs
K6xERBIGNGo9MavdVxoHDOhxvCO6/F00RCryjdyBXwiYtWgvBl/9aIq19Ncw4RJn
QjnBGmH4P3em4XA4yjAGBpfOnFRY7ySdywJ1DVUKsmL5/GRX8Uo2+7RiXYEcaPST
p0CaIKywpjxmfZaMRyfL2Uq9ksZcP+aYJM/W16bPcptgZ3jiEOwPZBiEUUkn0gdq
SpU1RRfiYf80qjpoU/sfmUvvX58sAuoUq0EX7wByBCEItv05Xyj8z64V5VDHC9i5
bpiNAjNNTR7nZUHpykHMK3Vgue2QvbcX8XWKan9FN2XkJGSWTn0UVfEpfZ9401Xz
SfYR2I3s3zNsTFYNIQim8xzc37t7QpPWbb3lF87svlJ3pBsOBl6OfIuY5lo7L9rx
MbfBQts9erOUThHDLAsv89JpQ5nUiOEGLYyHdj5oP/x4su+RtV2YchXLMEV07sj5
sB6EYagca+1j+AfeRc91vJATuMIPX2TzrRquLj0kAuCAZi/gTxPBPhovnsRFIAuy
PX97UeOVpIyQW7VVhshACrEAH6bL3lfEGTkp76am50idL4G8NPGd/kO7yaDRerLy
A7VuMGVEqAH0ErKtsBJHglN/TZE3wXYbRWXS7SOMlZqUdhshJRW5akLSOVQQyx2q
WexLQz0L3R7T2BQ8c2jIRw934zPhoLg9jXL98xgluvHWQkBmzRDUr9AiTMFMy6nj
4eWyBIsAJZDTcb6DVIR5hxz3XGBWkrBOmAZ4cVyEMn5C3HhqUE7Itsh3zSdjblQc
N9r3LKp2S6ZbmC+OG9JkRwlRCVzJJCq8IT29lZcBAq2b9D4UZXQ+OsCUMcQATQS6
4eGRQ19ksBmeW4QrBwQHu5+zSjpSv1OLQOmU7DqTQjeWAwmMZADVWVFqGVaaF2OG
j0t2uI9GRaQoBTEXQl3Ig0th+QVHtcPEcbieQSBPHKfBDYkFOIX/Q+jJgSGpDtxZ
9yV7AOZCm518crJQseLclcjuo7zDpcihx2zbkUO0l9r0q7Jz0bBggb9fOWJxBbJ3
zKGZiBxAh/VnfL5pgZn1VJ+HZROH5Zc2ysTq2jrG+m4mSqg5M/EABx43JDaKFU9F
Gim8d9qPElb6XpqD5GjD4+fSjEf0hP1hpMPlrXXF5zo9eGDIWQPMaWDtOtmKe6rT
aVQNgwSaxRRgdmhi3WvrSzkw4ktSzqvy39hjN+0vFbXhtjrJEmkctpGFiBk4pUUb
YvkSVEpCoQXd/ETGsrcblUo5OQpNsxfyiujMfc0//+syTFb+hNwteFeRHGRvfrQ2
LQxQVrQd2d0NSzoVqfC+/iZhGvW2P3a05jV3I2JgTjiWKhT40Mp9BnEOYJ81Ssgt
doeo+KMPm96njbO6FrexuBTNUvVH7uibSjx9zeJjgfJLvimOkXqDnz2L4iawX5nD
fjSREDyumXTEkWXSuFxcGevxmH3doufA+X0V0onIFmTQm94bV8ORBNvcVexOhEPl
FXJBmVJEGmYtSNDUtvTKVWZmq/NuOJMGmwMPftEbaFHeaxJJvfu8wtFG1nXzrxiH
eley2B0f3gmQhTS9ODBd+BfK+VAQl3Y+8TXdnDbW7n9FU3yHDPYg+XlmR5bEAAXd
QoCVvj9b1zEio090I03cFN2WIBzbkg1dPVnTC2fjQEZHUE4CPqXwFRuqM58B2IDS
+kYl38ZIjTupK4kU4qCwN2PjocB9KbTqhxDrzSohCApSRzqGqO78N9aRm94FRAEx
iQ/uI7mNJnp+3sB9G6ISZSqPxMeiwF1OO5xfdKkKcYLQC4V3bEFFYogzjXf0D7c+
rFZcfKOh+pmr6pbk/JBfn9hvMVgmnP8Y02af6CvZJsKAVhj2mRLPTZDXIgr5MQB8
sW1n4kttV5vOsu+WNr483IR+UmDk/Io0n+OIww522cogM3RLwUGEB4libcFOhzny
JgWpLhDrRrYcD2yAMnaJGgdtMZb941wgIHy/S7+ka37QOVfmPWWgjDfuwY9V9GX2
Z6gNICBll7ES0RBymhj8sOdKu2ga9zEDSnUqHBaQAWSK1LOeEbQ7OULOo3s03/wl
T4Q5lw8/q745HlYSCRlJYt28sKelNjZ76ZV/zaKUuO/Cf2JoQIdldg/yz8gJxOpg
QzpDDDce7B0ZnVynUNyy7efIxZXa3tmlxooCx7Acz8nV9SVGjzf5U6+E0UWtcjoO
zC0PV2mYgVEei29wt08wIIrztImjVF0ZFqFSRAQa20SyAiBqPkSvGesdhL8vgVGa
2m8iFhiR6T+GWoopZR0NZ2TTwVsplT+gRW8tkGCiLnqjN69z5CciwxRcRXSN7RDz
6Z+t0mWrrKVvGqzsa/s0y5jVkvez80pT5U4gw9HTZYnNNxMiMFl5AnzqY/ysAcQM
1uvUU2a8Kc6iXWFTq9oS/RuWmRV8d327bLBIg/uRvUH9X24Juz+sGrd09CD8KInW
JJG4I690u83BS2J5mhql+htO3MFwwa1LNr2fXZUlQI8ABIxuKvDl1cHpcwR8kSo3
bkiEBqjFbs66qNSowXtHn75Kbx60CvQgn+v0JE0kXJ+XJS6Mt/4jqoD/nLgKcnHD
62QDntKLU1SPffWSIccz47b4BjnPgs31fZm/Ji5lUDYQlmkLDEUWw3tPunf41A8y
54xKyLmjvymtf8wfKDM8dJsyCqZeDD8IGsNJAONw1wuzwBQmPrsiqXmXyx4/Mmmb
aKovcPhLeYFxfddYregj1lUOOU6Abd/Sp9c0gGa2g6BlckUxz5hsLNyLFfMngls6
GmKMIb7bl/xPygIkYxr3UBxqLtHcBKC5HeeQKFEzpbOunsb9BZtePpkW2PI4LnCD
rlhwOw0KYSWeLt3N6mghQhpjlBdOhKMCiFizjC/kwdXYnqjVxELWTjqbuNigjK3y
tQPGY24SFOgaxZhjULqpnzhOEI+mj7P30ezUKYnD+Nd318KdqE8ITcUomCVySXmw
9qW3GS01Ngg7pTnb/EMWsony9apHdvEv1qn5npM24Z7napLz5NWnbOhzKQBC0Ouk
GiRs8OZDVU7nMBB7ERcLnO1J0rhAIziKNDLCReR/93+tqLYWpTzidew99jjQZxYg
yuZF5HeQx0sPuVjb0N0idu+feo50pUKxz8G2W3EjXwaNHkFj0O4Ktsvy8Wpyu+Hx
ys+VuDWAtPmqcqC/4Q0DittsRYPa9twvBcucKkg7ONFFP7Xe2xTW960kPA1mTA/S
bnkdhEUhsn53cP0LQGnokH9fPKk4XJZhOZXOe+ZLH+/3zGhXdBzxLGcIJvl5rFWR
4rWD8zIgdugsTod8weFBO+o7zCewY0giXEEn32cQTXGesfF93rbj5ie3eqMlUkkf
cZTyMOm5upyYeBWh1iYufLMU0HQg3l/iIBam7BLAbsjjZBh6iRfzofmw8xyXS34n
nh4WO//2+Jk+puI6PnB9yVvkUiyMuXO02PnDM1RlDV+gTNZhZEbzv8w1NE5/pyvL
JWuRBBWGkDbtZkG0yrALnSlRzo95Jea0GMthJsuaGT8o9OC32KvbaK2rJuMaUvZx
E4odzNkeZJZGSpzpwr9NcLfrDDTlvAOSoSNlu650Q0r30ve6XyhYwHqMvTna+T/o
pS54f0oCWtzL7VeDK8lqOUa4soU/thj3Fq/Z86IMjMzIRz3PorCwTLf3KKS+LGzh
3aw2gkkVmyHMQ36Sr8kOlzSXkoQ46FZYUDktRGplrN3pnctqQdF3SUuaUlFyReXq
09HGexkzPMVpEWDeblUyEn1v8JVLndlAAxoS29YJicj7zXBDQ7egdHl1yzrh2MX4
IclZq+zBYwEFNZMK1jHSMdiqldaOpETyvp+/pXqliruS1puAfd3Qp99rqMaoP5y7
VvUM9cHEzd6H+cMW2LXtvwuNEJ0Ba2kfb9Huf3F/nJ9iVu8Hglhn1Y0L6MKvNFkJ
0wSc6mQkavNBlLiPTg5WTbpgyVzdUNH704DWnavoxBeqdj8q6TgXmwSsezZoSE12
z2q5CL9TmQ+iHgkuL89l/Nye7vA4Pqx6Pj4D5wrJ1uCcygtnpJScpUILwGQsRlkb
2TrhCyP3hR1D5YQRL9sW83PFnz1dY+o5Phr/GDhj10JDMML6BFBW7p3SonmcknEe
yw8EWabCvB+WVpc5+4evRFCrOaN/GRCEGwsb+Gs0QPMtAHVjSwtfVfASeFNmDm8F
0KR5j0TDbSE6CGgQaNlo5Ol52bKMQ7BImF7glthUFS+XfvQ4KWA2SG8AzJtOjPlo
RHzylSe7F3lsrfRaOkRGK6KKuGuUGrK9aQ+83Fuh6gNej5E+k9Yw3kz7EZwp/V//
5vroUrZSlV8agUlWkY6+cj+klpmMAI/InSvsmMzbSeNIWb5BT1EDQdqxp0JNy2ak
JKkdYObDV5MBk7cmacSTKbnfZQfU+fH4IIDnDmtdljQEdApwjFuDV/HJkJZ6knXc
uOc7UZZYQs3Bz5C5HEIp4SiLrBR//tz120be7AXfiYoSA8cR8MdO5cHxOV17r5z3
EYAbb/itisoe4N+9zOEIf+AzwjlTG9lUchonc2kQuFqqsI7bF1/E5WvrVcDqxtXh
+oJia+hIsvJapVH3vQAu7A+1rsf+UgOaquFAcjNnTe9NT+JMNv2AVRedTM3iljvk
qOHlaFK04p7ERHa99RjI6dnmVjRI5BjUbTPgJwiH+1PEdyp5HzxokQY5R6kGtCYj
10UWFC4SzXfRc9FOZ/m/KCVSU1+j4S8f9+zPt7YtG6XBq0GWur37gelT8/8+TPLE
TZ3cHOpvSu8Q1adQCDGzPMe1WEfVM8y4Uu5kEflJVa2gsYpcNeRKPQmhGy+Znz0W
Sl60xFERRE7RjIV8zUVRaCwpUGp+oGxPZIRNHDQXyQGgtRgRDunIhj0SjuGD63dg
Ss/eR+SE2BCq6p4gHs4/d2EAtnuj+qbX9f/D+VZzfbuoKZeNvfg5UvvLaoRL80d6
nIRAkIuqnEnQEhV6gTLiQjkJIPsZYOKDwqwKN97Q/vpwPCjJ5bPOcX34Dfi2kN1c
XuScvq9jngHS4NghnyxXnJ5gJRav5BFKNWalmVAS2e1jwts9+dIcuCXj4Lp6jBmA
EMART2+Cm2KWdz/KyfZeR8E7TWkaWffDoW8AEYL6l/GIl5hidpPBwtdpMsYX2Anr
iy+7kz6CXsU4NPPzaz6uB6lp4Ik3fDyrVsnnHKqFZg2RBfWhaEqM8WeyGbqIwNjZ
uhK75zWJvf3lvLkRuIFMQUVaayGKWWiRyj5qa2Uajz6iDcyNcYSiGCU7W6ffyUbw
CXFDQaSbmps9cFVJGnwizad2fy1frsFEvVcFffwOvREp3U/D5ASTMDii0cDojvVj
i62zChf0igwpOvlAhnY42ydWzCGoaEzCQ17HYj15/MJC6Jahfq6W5Q+8++m+RqhV
Wuj2KViU7Un+rQ4/a/phJuwZNMvJi0C6xRoFK5piyPcladVoRFH5EIvsKLATPq/p
hRfb0h1kn0rvwJM2Ycio0XO8s2YmvGv/1wZRFUjW/w6Ve//uyGuftDPqdBCCy8nh
LfyGekrhUtpclAvaHCdCVRANG3FdE2ZfiUTx3zIDRE7D8ws/lP/eK6bMYLVkDlYM
6Vwt5c0yPIpiIn1RS06SzZcu6jL+ngxZVt4E457dv2WMMD+x6bBLN0M8cRU9jjvA
SbfQr7zFWP5t1OsnbOnXrIRBxFjrEf5YELP7Y19kxpRoP/tGixbyb4kFqE2NvqnL
D/DKGZlnWz2YOypQqO0Fj5HJKLauvjRZUgnsvLgoehth+tdarRzWQXo3yyqTKN6S
xyJ2M6KhqStd3A9wvieQ5IVdufDOYvfnAjDuUrjT/FRD9pgCQ0mcXrx2tyGQdRDl
ItuToAe1lO+ZTm+WCGx/uWu1CxqWOJxa1/afVd0YqAeEIxAX+rqbqVNpz/hmbPOZ
urlrVF4OAr33ccLN66SeRzWM9qtkJpJZcd++L/ajRw8Z3bGPR9lup9aMasvyBuH5
YYX+EsDD3P+eP+OKjcYkwrQVs3h2irsTLwDOkZzEzTO/cPdGS4vCUxxaWuX7aOlU
AplWJouIM8fQ0T4vNOg/cNABlwT00kRTOuuDYAgJBNtMMLmpztnYe3eSuySlYBso
TyPvUfq2zrTZxIRwMSnmYVeznjZrayTrvG7CDwdXO57O/f5PaBXga7dqmiyvurEe
4tUCLu0hKeQKFt0v+x31/r+fobUkuo+hZia7zyP4rD+9VSbc5F/UrUE99FfrHKQf
sR61zmopCktCovDDFEpaOEjKHDDLpL9ehZttN1yoZ1rUvA4f1wSXrLn3pJWzK5F4
UlKzL2LC314mky4umyxpBoayGdq6MZqzYsM8jXa48HIQpKmDeQWBndTA+jd3Qm33
7rgZtfzW0RTt2zgMh7F/30xDC7POSpn2OpTS4MuGCIhCC0eLlstRD4v/zURoRE0C
ksWlexbw8tfMhO6Y0g7loWFQh/CvEovCNIiuTV0/eVis0TaCA0Tp6aXGEMk2cI6J
CW9jML3a2pv2IX5V543qPyf2enZHkCQva/EBryTK0N/pQ0R7D287kn/2vbvlLBz1
CFoUH/jYu+WIw6WeVUxHmZB6nAE5GazPZWy9L7erW4rC5/PHtegY6Z6Tp/Q8R3Xo
lItjmbkbAOHLtIKDtfil8cURxkYXYBUbcMQSKjDSOnjzm5RRzfY6cseDGndWqpxP
g/9I96qdh0GZkhh7BohVpuBlfTla6o6AEbvBmzlFrf+dluZEVVfvhADCit6HTjv2
jzkugnN82j0rUKZ/IiBfLo4OyLyHRZFUUqfvZJYOMuEz54QVLsVOmw7xOAn/TuiH
dgt/JmL/CR6EKdDxOE+sRTZ3sqqGkiaoyfyL2mbOiqfGtwk5Dh7ZHbXULblFt2AI
h6aWn0WRIbmtXeGiDCz6eEG+IwkLl/nEXRhHeH7lCyx1ZgmF6LaO3HxXRvC5HgDl
Bw2ouAwN8LHokXBGNKi0qw2MyALhPp1wrJTdWd80wbarY/Lxfcnne3NqaO+hl1ai
qvI98t0HiJtXBEAZg/dDBeOw0J5wLMMiA3cruanEsAY0ueCBHMVNkS8TBZ3zHpb/
KzlzEMSGSQVVtnWpNHGkrgZLfslYvyu3c3ci5vjVB6zJPyVEGR8Tzj4PajbEtISo
Paypn4tPsAtOR6HcKGoUTzis2Pfz8vSeEWXuz5au8UiWYqtE1Fnx/JRdcmhm15BA
41nt6efIltm9hQf37OmLBM+6F5uLaruJfsQZTShDPkG86NGv5euOW7eE5TRwTIMX
MWzI7zfAfi04mu3NxmaggnKvkIr+vacZNVJdzH+sOObmST5Pg6drKu0cVBlu/FnU
PUa1in5BTEH0XEEHe4jzBbIxWtiPgkbV1YksqJIx1oyCzQpep5RxCuYCD8GPzuLO
Xo2IRHFJ56TF1VZY27P2BFuStY69fU1XimxXEdRSFjxWzmgThakO9uUsCS5NUXJ1
09BzsIVxJx5uCJe/vjkAYhESR+UKpgkFhWsy9Hm7zNTvlyeN3+w2ndodUYx6hAQx
KWB63a1EK/iXg9SuwJQbRQ/2mf/hkbldTcwc6MT80ecARkEpOUdMr//FJq0L6chf
IVrfL6Kjuu8ed2mLemSkHkWCBZmzbaWPKKPL0VqA0sumHLqE0+gPrqVkC4cSvxu3
4oQCGJ6zm6PP6a4Qg/O6ZzT6OCnRb7S6M/2Q8Gwa0h7YjajMrF1pGFaJMWHa2EFc
wroFhcJy1Mx0mDh9t9rsYaHEp9/0zyQEshnCVWueFToWR9U8b8j5IFqxYyXdndYj
wS3iAXl0uSYqrqxuD9nM/b016vAk9ZGVVC3Qso75lyjPlw/yctIfbcpSsQo5y/dq
uIyxu+a1ow5FaEQfSbIAFN6QJGF/ALMxBWeTtVqkP0AdSgk/fORodTL3Ojz+Iynm
5pRz87UiY64LQ7QYBohrqx75RRXVAgaGUrvNNMWq2h0gF6IRYXTQ0SfxJeM08Nf8
WfR0uspQ98HnBaoYz9hWTARGkE7hb8zRM7QTP/iTawQ4KWwvEsDCyrQvC8kegbGK
EVyKQxO4WIiKwYJ2y/M/Ph/90Qx22KULCS3zuCs45OVWl6NibJToGzoW+LiKH3J3
C/4TjXwQEeizkrnqxdbGKosczB/FMsX2aRZGMOTeyLWGOfRjFMC+jlyJWBH2aMDi
7bMmc2rns39P68+RaHRQwFkOB42OGckFinPJ50o5Sqp+KVRJcBWY3YTy4B1JD16B
c+WbkQZXNKGc8dRpHwivUnVpWZ1Pe5+on0iOHt/StiWUOgWGxslsjkeACJBZU1FT
zNN3Rm//2zT5uqhQZIVMqDXBC9t21Tciuyo5E/0RfKFk2SJkTdvf1gPlfwRL6TGl
tAKTY7EjubSPd2ajo65Ww0phfu+l5fpHq/4ubZyoNk+MwIFl8z82Vv5fuzO64HUU
0gdKD6nPJKM5T5+djuPLnUK5WkGKSjLiPSeJkJyEzGowKIqPtqvBoqf9OA9WeQm/
Mxq3AkHVrxd2rXYGf0oedRmulwa7JCLWGtbAhjkOiljOaZcK0YPzzlh0oNc+R53I
IOdz2KIZYysL2H2HOgR/vSFPh5KOT1v89+YLOx1r0Q7+8uMGQJc634wk0jCGI+qx
DXYoCEhsXJR/00l1V/9mZFvHFXNOYPvC3dnluJGuZqtyYHtX810LyKiAyHr3zCcv
sBXFnHeRGru04NllL4LCKOw0tGR6JpEmK7dCh9ItNlH0J0s9WD4p+c3Bk5khe/qD
jY8OkEvrZlY+sqXU9d+V9OYL3Y6cfW8dGHXUSXMfj6FvzjTUJxSSWZs2Nhzmlobw
T5vn27UOcfdNjRMFFMYWlnJH4OdJJrCQ/+qfZeeXdr2NxS3KUVrRL9BuzpWtgp9P
zLw3p/CAEdyq5bOdaSrbXgp/xav4FDeRQbu6sRQqCsRwFnsm+0+JT9zD+fAwYUz3
3upgpdGy4zVaWLKBqBKFY9QQuvaO1YzpR2yGmHW3uZXsgDq3MnXETSlSIIPuqisw
muXwOTgq/4aWrYKF4Jp0dsVTkO9T6npOFwPmqXzevJRG+iAKu2MizLP7we4ry0wo
msz9qlGYjTCqBDAn+tls2WjqUY6QeHRQBaYR/77gFziDt+A4hUp8JAiBe8u1kNVC
DUfORLz9/8uJA6AhcxvhrvE0GirZ67tlJyXRnaP6tff0E19nVb4uN95tOrlh5xcZ
vS+kI1fpSmX5FxcqWMKQGZBjJ83ACOtcOLYio04ESpSoIkHPaGVIQCrtAsB+iroI
GYqgFsSNpUWT85rtgmvtCBQTKxmi/J3I8S4xNlr2hdoc08rewjH2vmEQsn6TDYbY
2t1jDvVo+9uchKKQKTJPvzFKkUkg+Vgbatcv4lMcZGQIsMQqJh4WsHwCIYtJkOS2
7cmP5FCorv2GkEqTScWXwKbbjVDhRSA1OAHd7xHq+NklyQmDSjksgaq1R3o2VVmi
WyZmWRutrfqtEBTMBJai1Noume1etKm8YHPNw3Edu3WFkCgUH2H2mdcSH/xc5Ld9
GB91mLMZvVMasJHuPboaAE3InnJGEYndm4WlzdVgdgFlb6/BbPaowfXQmBXhVsVJ
EQLoq2vrL6Y+YRUjvbsBpV3PTxH7h8x6QStuIqmqaZ5JRZ6sxllFD/sv+tjRhBXl
voxK5llR7x28oTIRlV1le7JVQJU6s6EWYM6Y2wXACDnK/tfZSarlD5Yt1aH8kxbf
kw1jon4GUJLuJgMdstanw+dFC48GVIUDP/oWViEK7qk175I8Ov3U/JEb7Sg9hKUl
t0CBMM7TTiyDXQckzJMPUlPrw+68S38JmuhzbywrmObZFJ46BsM+KQyUcI0dlYb2
my/FZElZvy27DE6zgOKOfIq7n/+2bZL1ZTD8mTYr5piVUWqzq3HbaigNDa6Dh4zt
KEU6ECknUUyUpRoqYTPimN+lvd536do8+syIVHkBDdAj+jGbpiy6wBvAd8j4Zlx0
lnLa84W9F/kKxkzKYVYl5dKj+zvm3gsmR3yIZTxgxqrpoZimODn4stBzla0Fh1DQ
feTto0cYSwxr+TI7D7yxxT5ccOM1EG2wNUS5cQLBd5eJvaKYwggM8nZHhNejLoIj
bAlRXHSTvtuaSM9zhYna4suMGfYfUDUmH4KNnC1mAvAJuz0yKriRVQrPOq6J6z9V
ocbjSdPqlOajxgGp6UpMJr8u6S65ZLIw0Q1Uu8vbvaAXCH6I4lM2ZQ7rK+aIHFZC
kvJOSqqgMPyb6nyUcUFuV7YNkH+OmDT8WgZvPbvPZBd3VySIr3PheiITrZZOgNrq
t+j9zHBnE5/O1/QhySVTsROzCyHNX438h/Bjfux6fuFParBSCDaZ2MLJ6YZ5DLfB
T56tk5nczvXV4sBvA8dvUwrXQvGLlM4fzatGcfnCa2aK7NtMqJKz7ISkPf8hwoWa
fOji6Uy4VpnPD684cbv8nNQlbNfSG7jCsl6nBBio6vQ8XyrmDu7iusM3RnqFLnFA
yHtInYvuh77dnY1fOOPVhaBMPR+3Xx9Te9SIEiBjnMCZ8rA/Z3Soh8LRduooyjKt
TrOhv1f7RVAsCDtCcRP7NI/14uCAc2gQiFVkuYVB2VKG+iC1iCHXzKfKROQJodyA
E6/aH7ApSmpt2pQEx0bZgzQ6+P+WzMUjjRMAMyt4CnOsSpCSWO7vmIwtNBdsmXn7
85PQt4wy/fvsfIJvMt25vGJeo2gG7/VsA7JksL5yvo6H7WIwo4Re+sdyp/w6kvYg
Wkn9iTarK11hBLhQIK9QUU4ZCi/8YR9pMTfi4XaJz++SGhm7/71lerkyLbuuzSEz
dEtrMCl9Q/eilCEaRtJsGTWHuq5BNWqAvKXjrDoGoOkMxUlok1Nr/KkVizhJ1Cmc
TiMyvQxXhZyAh72fRlkcF8FmcMRO2MmW8C3PHWwcGY4NskRRwJyzSC7ifGaU+gmD
aT/K9vP3mg2qK+ONdJ1roWl1+7a+g9j45WZqsqvUwEevAklZjmWdlIqTWq4oIHMp
DFyFbJ8l4xmfj8ng6xduj3G3IemAkl3XiurBYLcQlC3m3+UnJ3HR1/3eKbfSgpp8
CfqM1J39z4V7FGOjMyGER1WF3q+55FQC2mPyj0ZHO+LdaXz5IKyIsyfzetqDotHp
VgjvjWEu5OphsyMsELRaDUe7le/8bqUWk2iJeO/bli+gdu8HRIGwsovhqbTNycU9
2dAHQnUB7Ln6bL+2d0fttFUga7XW2QzOVdnydjxkdqubeawPjCS44Ox+UZFBmGJi
5wJUmWjaRq7XmoZFdqquCubX2/TmaYyoaKXjyM9weBBgvMXMmlR1KFdX7AojBcFN
vLCqTcZeDb1gR+dgf9g2sky+FlXgMqXEepcjJ6ZTmbtqMHyYd8nE7oJqRwsRuzPd
kNfP7R8X3MleI+TQrPlF7FsrH0LKEl+NkYOyorMVKgz2ig0m0Ci7/lQCTfF5z6SO
4Y8DPsICDLr5wVqQfwTYGmAWBVGzF6IIuwo/nOC8zB6ip5xalXMQd6lUedZfhMhQ
qMRxHM3BYQTgXpMAenmbe8Hj9HqJc0CKXQPlNj7J1Q58R97D9HbDafZv4zkfBjnN
0IEfjXA/uL0sRJy405m6NziL5ZQwrAGbQwORtEE1fpPW4SbgMMJstCaLbXHDnv9x
udjIobP/BoFzm0oSg3Z29M92vCsnnNclnk4Y+y/19J2gjhQ/NnyeXIiF7Cd0Qh7A
jK2kR9gIbR4rc7rrQzPE2kWw9NcU2j52ozuiS+m5jtMdqIlrA17GtiuJSxx1eh/w
phoRYdKsbk1f7h+XDuUPWKXPL4ulGxTEP1EygYUuSuS9fsQn3rYpj8NqaQLllu39
Yp4MdfqG7mIrtsFlzUzJEnSg1rfVE6Y9SoEp2CM9jrMO76V1AC+vUEtcxwbZodqC
OcZk1eSahLUI5+HJB38Qiw7ehowQNSor5N3Vwl+izrXxXkYCtO6+GoZ1DjSAOy+v
288G9JmtuSaDRxmlX9UTASUg7bNhYuQS4XuDiG/7lGfNyYnZRdGlT1vB8O5qI7vh
ve3I0B/EVFlxPssrd5wWB7S2kCwVmGEwRkOf+Jsxe4AGq6uITwNwZJ9QoBIFeRmA
0xv649vPws9AdCAzlxhCcr1kjVpwYoVH5K76d+7Cw+hsNAA99JOKsjKQwScQNKVC
ZhvqZAWMvNi2GPXHlHJJ0170D5ebOdQtaO5JxlyZS1fCoXQh36ELs9OpJRyK/U8m
pofx5OnryklJe8haM/uQ9hkRAZHT/BvrnXEGBUKMV6MkacIgxi2jqBnJrLnObUos
AlMGHfUfMoQ7lBSR/AQnNzIHgHPmK9PtCV2OHP0FAyPL/+8vH1mx5zxjfJhMUQMS
jy3u+stM0EIHrGOtupLvwVMlKZOIcktMB71wjOlX9D1+2pB28Q0ttZanYP85iBGf
lvGM0XufOzhOJH7M3CUPJ/ZtOQvtVAZFjcwiySYd7E6ms3fr2KeRENV5iUi5ALrQ
ifQoFLhTzGr3fveMQVapPhCLM/JQIWPr+H36g0LvMXOc9/TeBKJLpAA8jQ3ywBcR
LsriLbRe8cWwVcm8J1CeXeNOCuzx6pEwFgeVjpJHX1CcCdrNXuZs/txjVMjPAeVc
P6yFWOF0rqpMinHefAEtWp/olTMyzWUmGIaJd8h+Ht/cFKYkLFZ/YP3ssBcLffoY
7+iQFv53FnSTD5sxRKT6iq65jUVbT4wwQYvtIzh44MdI8KJa4HEF+1/7A4Be9VMZ
MDzF56m+nctVGPX3iQ7qxJXjkXVSuuJMzP7eoLD3AZcCxpQ+ZJ9mdVxvd2nDszxw
evTfar+6nHa4Hm0ObNwRiytusqzTNuvY2mKnS2GVzSUnEFF4VMYUS9SdtGLpf4Vh
eatrm4JTsBP/VsThnVeZ2mZgULET9MDw6j4C30tPKkYC/WVwd9ZMML709ywZ+C/1
py9c4b6CDtqO+ls5IL9QcVghpzpoVXYSBuT9WXvyEu5TB3+LZcfoVT68fz+JTs9P
oRnXCu8hGa/94whSVJtm9ELg4rV55XhVpXpzQfYkGELflnq2gV8bO5a9hae+80oa
H1UNusWBt6pilqCj2T+JxxJy3Eub+0AUBzo2hEBxHwkkIsWr4d6RqD7/E5OnyMS/
NcZgRybjpK3i5D4Ax+39tv9fjt9Dn92idA8tXsDpgxoQNaGeov7gduqfccSzrgsO
ml35S2xOFvLkRxxrKOGpxJ7euonWbvixKKw/LStrVeM3mjK7aNeFgUA+sAgo2Geh
SsmawCN51TmiGCJ4CvlRV6WavwTumRii25WfIHCZMk+S20JrvLglzNGzHp1R5r3X
T592ibVo7g6CWuLXDPvWJkjya1EfwbZrtaS8XiJ7SNqegvFqapSzZ9RH+m4NdbeA
L9Jfk3m7z9G5I1tyK+IXHZiXaz4oL8i9HKfz2xHwmMNqMOEB9JtRE4RzEDx7QEcr
goanX1xrqcs3eYjP/Vp/4wAoAJZnw7xJYuwcl0rrnpOeRxitct1JjeyzeUMkDuP9
ZGsMl5ikFqGoAD/Hw3sRsBCC4A40USaQ9ZA2MNP0jCmbDk1PXSWhz9879sx+i8Fg
OkrtWDOnLNDiFMYvpRHbqVxWQ2/FqHzTmlELta3IeSoGbwIHdc0xz3eUvee2GhEI
EC47GEI1quNlXUmZtJ98ovZTMBCnlCo0BlqS3rStsFLRr8U74LxnQ4TAHrjgSrIL
YhwsxlIASgHrcinVzp4pPJZFOcqltYIuk9sLeXLKoCzUWzcsh/fKs1fWXSF8hgZ1
/1W1ipZbfd1XdjLJZWGbHSIkKI0fQeCUPCv8GRdz3eYUQKbxnDRXife3UV0ROV1E
oEOTTe2qWlQG0WerhexV/u5WPisWRYcfI+mtROZgo30725ogodNK6Uv9101HbZNR
0wkxrMU6+lYo1vgnjxoNmaJ4iE7MlUSQuBdMnhicZZnFRIdPnk3QOLQdX4IW2jr1
BCatxeDTX3JJxTd+h5h68QegQ/EiljWcHwtO7nQF0Um2j4pZavcm7Pn4ICxTWzel
dJV1YYPosrOQaOLsnwqg5+uPurSY94Qwgv+OGJLa2VDg+yXu9u3DLuEKdkGKrqoQ
W55LEQixOeJC3fsdWWQ+C2vnDkkI20VGmyQxqNai4ZfxKeMlycS9R4Z7pKOiOe6L
QPD1lG95/+2BGoQuPGK+eSyHqjjzef5ySavocw8qGtW1qLZeiT92qyxuFc6UEs0f
8HPDbSF7xLxQtwUjM0VntzLS9b/h8Z5+CP7bd6wR8AUFq7vx29Wu5wHYJ8GXXiHr
CeNaY3Th+zUym9AF7jzxA9NGsllVFRJtMUwI3SE6gOGJwPXU2x3dihcCFz57SWTJ
bTYQOGGU6RTiSK+lvYvybei9qqGbBsKYN5FKAmKPqXMz1aa+oKVyp3XepQxFOXXW
zGuLGUtM7DZZ6uWH/3n+d8p2WlitdTDw/NWQEdps23iMd4HFIYZCfzARglOszFUS
aels8EMLYsZZJFmZwhq7fd2o4aXr1WTe4i84TyCl8AMzSApFcE5rTaBXYaRPcS1j
TXdJxYLYzS0DApPxhaHJF2cbq7l8ggBa/HRPlxUiBLGB8rG8YtIkEYR4xkafIia4
7ySYGYz/UW/MEhPgJGj3vUzklfH6Th8+aYyoepbviSad5d5VGVGnamICB3yFTQV4
u1JPLRYpxnfSrqfjnA8gyQnjb3hn1MSdpVraCpCCUclWd7ihwOvmjbwE+fYrqexS
Pf9e8LfF8mlj0Xn7GoolBifU9wxUv9G3nmuorWFtHFIBvMSP38v8OQKeBOLVjRM2
6Xdnt45ndZkXdcjgcfY7vyu+9wZxYjeotb89fNDesg4OF2BVerp1DMOz3ywauUGE
HCJeNs+9MzVYkTa3+m2kKJb09CNmRxd2TMO0dV4MbUKXtqoGYhkFC2JSeBU+/Acy
Fjl+l7OcNEfJ0LpR6zGrfKi3YURj8BFAlm5dzeSAFmeUAoAeOmNH5/jS/5wBX0cB
kPh+jpSfj/oAWwbDIaqnReIOAvxbQUHyzJf/9DoeucpmoZJKAZr7wXUAU1dQqkXo
PDcgvsDTkcxoqSN+pLmxKg5RJcA2M5UAtWoRtVKohoL3kqRQNUfBChQfy2XfkgQA
koN8Ydbmo7OScq/PbnDUhYz4qekDS6vcVMdpXfF+7bSJcfuOVqIfSWXuOzlttRvV
jBdWoJmM6K9gJfQz2oUYgTMGdrlgAiogtZ1iVnfu1ai4hGhjrAujwqAz0ElP5A32
CmFIl+Yw0M7you3s5KPymRU2TxjhoKGD+pqAbtnJ+WK46EcK7yI04fB3B2su9fTc
xYcRmeyJa7mV9NhvDFaAdWf8V4T6ERL1NNgv0D6Wfpx2Y0OE1oXCzPcHzTzPmRqI
OetzdJoV9I7byvKLI1UVr8bBcQeDHnIDGHHwdu2lOSsd162nuGEgloEBITBQ3rQe
QuNLULMbPBZ7tzuouuXMMzKaW8iEETUvTkSMobMTqbs9fSTLRMeDcyVobMGtNMIc
5XyVRq2Ry/Ju49SxccJN0ZICz2xXOIONJg0vuEbZhMekjGu8p+yFPtWafp3CSrkc
87A74ch24rSOMe1LeRpQI5i2SNzwXMhn6FORl5SyhY5uCHhxCMdpIN2VnvO2G6ar
/9Q+QRk/NyN0SVAEdtJplnsEPqQ9XLoMmfqZv+qTqjV/kiozkf6p6t6cPm5RpiZC
NnKGp5eOK7VDUSTfvHPpoMCwKkXOUW0vKzsY2IyJ+SafjAA6RcurPxrarHz0wLjR
1a7qyn19etszzyZliUrSR2+VyU1MK27t/sPsqzxwBH7ioHBrhrS4opu4nB56j8KT
MYkHksseDvVeAikdUUPk1HiQ0I35FnGiqH3V3qkyJOhxDoYTawuN4WtsNSsK5iZy
eS+SvlN7BD5JAw089ZphIXFUxTj5C5z0rG1HXqjJxFkd42oDts5spCcQWRKRmCVd
xb2RNRpS7MXpBMzcTskzXCRMcEUfCMwPg2VtcALPgkmUv80cSVn9kEV2lYGdqLEG
hIO1Pn6UgWP9w7UP/3Rb8itSEczoeUZlMqXqm961pn2JnXz+aOWZaAIav6mDLYsL
faG9cT2agEjIMQLFNcfKtUeOLSe/IPox03vAvcNm0Rr6E83Wvn0bVZKuN23EfK1t
1CXS6JZ9LZutE5Ji/OxtK6cfNl6BJUM4q4XAjwZr+ITCs4z+b6qxnAjtRffWW/uI
fKiVkOvorhIdRJGiHK2Xwyh2adPFvKp/TMbhLF+RuHiPnlKZis24sjLppE3KmOYI
LlFTqBTXUNx8AJH7gbbHVlg8d3y+0nyPyLk84Tb42X3sUPqwTLLD2n5tCDRHxTY1
chnWJnIZ9m0ro0krsgXl/S9I16NymH6C91bWAK9LdjhMcZyQF7iZc1giiaPdf+DA
7FSDXwxX889idOO5mJ5aecxFEeH8EbIP2EYg7Cg75jh7O1TCJI6Amz3sGAlPu5WZ
qZ/WCLZpe9Gx3n8xBP2f5QepHKMytwAVU+nhRB1s/xJ0vOjvyZj5yQ7qunQng3OM
9+Uz+Qu6HcZYxyeAZHjfAv9FQOh3UtmA6xWCuApmpOvnXGEoPrRePVduo4fdcyMH
FDP4AboVoM313wOxCYB0B1pAhrYyIPSIWO0PhLAFGkAMN6OHXDtsucuAZtI9cIKn
C2hz1MHbD4IhTqeZMmEQthPz3dFDZyDp1ofXBXvtqYdH7u2StNGVKUBSjYodzBMf
ZAUJBx5r7ywNRJr1fgxBYPm7cwNq03egEoqImvRJ3mTvJv2x+9tfsudQci2pjmlD
UzLW7OOHLFiuN9K2saX65DyE4a6ArXqt0pB7G7csvkkV1vo/hSeFpb73IEZQFlCN
3eQU5+NEiVZxgCp9o5zG3DhFDJBKGDe+NEduPkvxTKRqub//ObFYiaaVtr6p5rrs
3Zs2pDj4d5pEHzPgGFa33Vw5F/JrQBdc4NUqw8XjjBs43fzzaeLEop2rsxSO94YQ
hy+OqF/kqv651tRtfZZOAhpOTQ2prAcBpYqwDzSNmMqX+uACbVvENR3wlnrqogvd
40bfI+BsAlmWqyatsYmbalhWErJvM7EPZEMahCcUGtnjhAOXTQUDKny87n5pogWV
7UgXpYoEy99RcWfT6mjaZ3Jx9pdEI9toVKksXtejuH6h7Ti7CT2YxSuDrgXCcrZy
4zqcD0k4mJBV+k9hKT242UWlMxlEav62URjmraHCUz+v9WM7g+7Ox8PXn8dFhrRM
zCEfo+OOHWKlk73q0hLJ58UW5vhvPXSAeQgVPn9qqVGaiqaUxHmmf2blx71lZWkI
48fmC2IB2eMWeC/zfgy0J3nXfw5ZUAJH/oozgISu24gmllI+3unbrx+ExKVXkHqe
o87hV1y9naB7gRAGYfg+dooClocTuE+5CQM7XC5tvtu/+pmReSIzlHHnw55yZr+m
u3iEYtrrC/7DhCu7V0dx6J5gXO/MbcN53/HFhFRaMX2/aWX9+bldRgIYD8ziz2j+
S8jpNVXVLO9L/gH2v/vgj0hiFRt0bUMsAs4bIUwC92vIuO72jG6SkZUVBlO7BRld
gQ0F62+JuDvSXU5eiCYZJSH40hRpI5UG84NY3YLYvlLv/CMvQb+vN8behdwwzgaW
xRYRcaTPXyMW09wfrkq1ekrHQiJAY6Tl2ZHqgiMZilKZE996OqdwBHzbo/Bfqdmf
w8j289zy8AaCJAXtlmlwim62AtuuQaRK4bZWcr6gneRmZyYSgk05jjl+5OTD2Ui7
0ycZR/wXiZ5hyxJNFBjG4ZQ7fR7x3RN/zOQ1dw3SodICwdOxQR9eYpc0OhELOBcs
yhyigdiN1ZjqtMKXakk4Npep1t/E5O0fZ2PEew8tQZRW7sOOi5ZhLZSayxqVKspZ
kwXDcjnmTD6Dways1hTLaV5FVrCi9bqq8JWo+GGKFV6XXSPgNKnKsxKC2tTO7gnN
pn5K6CsvWuoxCP1gU9AStphNtqCboCWezCnLINHuA7jsv+Aqd+VVA3qfF0c9Cpfi
lX9dicP5vD/PbSjtWXdjllwBpaoORLfK67XwttnDPGDspkdbSEyg1wazkoC1TPLG
gB1cwoXKJB0j40GapKqPwF58CiVQVOvAkFRZZ3WVLUIs14oLbl4nAdGrrpTsfPkz
mpcJUM1zeQ67BZqmOzE+yEwUagtcIKTZeK2CTVS/jdumXbIXiAQzx9OA7fUYCYGP
Q7cAKMUTpMFbmtFGmyGQPH9Xb2mz7CTrMrTbrMlrzd2fQqZw2x7FoVYE52Yuo2Tn
PLbwLWG89rCUOKMekCndMDUJEQ6FapXANgbXA8NX74INBGHVWTswjuNGqg7vlq14
CqxNKtkPTS3IOtMdjzGx29+AoW1a1pjz5n/dC7ZIXtW7VJ9tEMKjODZdLJP+6V9y
7qy6I8uShbcbhmazuQRfWLVmDdXb1FHKugGQ2kgp5ojwFyNlnOiPXdTl1fnmfSDq
Mpdvz0g0t///7fak9erccZ6kIJp5logN1cV3PsWlNRyDS7nK+bhpnfTcZQdrEjx+
nSL0C4rHTG4Qi7DwgB7VM0lbi6r+8HuwqhBsBw82xXc+tNsmQMVy8FREC/N8ddcv
tjecJ3RcT1c0ZIsPhy8roUXx7DM5RJeSpZ1E7bL1DFl9iGJbA/w1cMM8gX1uMdtm
qlk5fbTGM+A6SiXmsnAKYFfwPnk0ZqPEkxJOoYtbe2hJ09D3NUYaCnaUpJC53LEH
c+3EdntFZTm8i1yFo1onXZv6tRhUXrmoBxpwtMfqqk8GMOUXNfEHshRpPjXlZocL
mHeRWPcs66vP2uZ403iYwzwA05LO2eOPSWImfkKEilcHwKg6Bvxc2U1Fh8ZqvjSi
ww19KYtc6H72cFbf8K11TEWgVBsvztNvABY/JkAd7vj+MoZWCmQsB5BMHbtW5iV+
Ih1Z5m68sxZQi46jySYdJHc0OAQ6FjB6Pb4texUjR0fqOfscUfktKjnWGZ2iItkf
fwxr+sg4T3EdxxEPgrdbvBvrVogW19h6DkSgKD/z39Iav2vbVRwgGcaJEEVhwpz8
hhUxunMMsh73JRNRkW+92MkkMk/VYQ1gbZZONBPIpG+IjH7epZPpL3mg+VTIV9Nx
1lbgk62miwZf0+4M4Ktmar5KqdmkxKeZdzXMGlRiWzVIq7Qy5FE+7DgL8wKlZXuG
UIIHTDBk7aCjQnOYVgyKPqUCGarHlPIgQ5rwEEjLQXXZZqyJyuht3ZwQ5+7jLPHd
G2OFmRfX4TY+skcBqdzA2bojRL9GKav88WExJI3+hLVhqFisKFx/8x8cqK4xTZzx
H7K2MVsQVjgi8yp4SI5mgzUumueiGhIe7miWhEkdTi2bPDuOiKs/MMuyZcgF3svZ
d6MMmn+0L/oMJSiVqijAUhxgFaq/LFmjsMrewM5OpP3eDUklaNnrOty6P5V9UQvk
irQMRXZBlUF4b8rpwWxOhp0z52lwsqlvnMdk2aKdS/ONkIrWB7jnYLbfgIS6gLqq
5+5NGdZaK1peEKs6T1hqsg9GeewdUom15oDIzkrUYf8sZVxw6grEWovq9W5YCiTm
U3u0VCwZ9OsVfpBoTYkDU8Xd8/XeHc08J5XkrtGLxiy3SAAkrVsbFsl9zrTD2hab
Xxw02+5IUA1WP+MLl6yAS3bZrVwQLlEtVwwTr8dQO8HrNeceHumpXTdU8IKR4YqR
WvtmcCCeOZn2B+fso7/hU83e8U7WubdT8I4ofiDYBV9muBQ088g5wfyloKRh27fs
uFoGewM0E+FVEKbKKdmk+9vb7Jhhrh+vUhjMjub5T++E75sJTFFYGA2NNU58M3ZG
n5vyhqhdBsFKIkmDc7KpVBg1EC9n0nnzJUFdPixr0DeLhPV7StWL657v6NlubJKN
WkiK0b4zxJNN6lTHOE0BJCS0egCdMqV0/ots+HmLuNvzYEtotT9JX+KSLgEOBIf3
k0Mj8cCyZTCjovj36Mzef2aeNPut5vfBpu74FNP1iQrCtpxxOjOZ++rHUg+Nt6dg
STIKEalS/Rw4aa/hwQ53RzRWgZ6FDoGzSdDmidZfzDWMX5brmAK5pBu/NezXdVxC
SJ2ydN9sbp4FT8ovKR4fp/JHEKLZ451GH6UFW3kpMz0qQxR+toCssVIj8jCdQBvK
y7dY/MejpiAIKmH334lg8rTuc+SG06+5zssTg64Z/S0oGt9WAagKFTogStOOQ9/M
nycMkFMtTNfc7zx1pdiAl2SlSWRr+sadKtSNYDX8/uyFVQS9jqyhfwHORbyUWYgJ
DK80t6wFh+hvOQFVatVbIJml+gR9CJUHAQfHFmZnrSeGqVY1YpIMahiWp927bwEY
NlM75pNHt6vwbxWNBoFoOQ6JZWVmH6h7CItUYW0nJDmku5VfVQVT3BO6peJ6xGAj
CZuC8C4DqEMvRbASIietG8rQpbmTyvL/Gs5LbiT1N43aw1cjxEiNWmWbVp3KFBzI
EVoMCMQlMcz0zvPntSG7yN9tKN/vCtAjLPB7GgRimAXbBW1M/acgSA9kCPEE6MYF
1y5+2qhzHFJyHhea4R5poVafZGF8zSGUKOmQLlMbR7zDeIdDDw57RHwgZtrlpDif
3zj7UdQ2Sb1n4YbIFoTX0OGnb5SpoZwvahglgwxiqZY7rJ0+AVXewq30KVV6mFlj
PjXIh5TZgn44X72mAOLoy4V6QRlOzPsGh+UvmeGOGbelrx100CDWPTarvHr9OIh9
eMEuZolTPb1+ddvDmxmzzczO3TkO+EPujGZ117BA93tCGYjjNU1gtURiWLSdrEkM
b8SGuHF70aC4zL/4H/5VPanD0EQu5qXvnl7bpyrLaxliekpyz1MlHCVa+aaA5nRu
S1wDQ9W5Kck/b/dk628vqhoGzntV5GAXha6CllIL9xhLz0u2f4sgeHBzpOYSRQQP
xd7plf4ktdJhKBjG4clS/1YTjGgGl18ZvTLeAhjsHgrx+ZMPTMgknSYF/xZFsh/g
HOH7pSbu6JhzzfkHzjyBKFMJzw0QGaUX7kGpoWvQPyMesIm0cqUSCY3pFQmqbiu5
FMhYTBZvp1JBOsf48p11YOpka4MxSMrso1iM0+Hks2IpGgS6Kc4y0WRU8Y+oBsqh
8V81RjCnnshjM8xHJvclPITGnwZKCdo30jFLdbN83JmSHGaSwbtYLbn1/39Iw/qo
GPjCudvhqwb1uUVvAmsRoLpvH27Z52Zc3r64jmkCgM4ZAaWJBIgPwN3+sCbpufcD
1TBc7mq8xcZpGb5NQXcZYdyvSa5iNzpJXb+k2RS3Iov2iKbzjk5bDmXvHW35SMgk
G4W9aZ1sHUuGJ0SYNoLpOykD/ahneCsFh94mYMexTDF3l4roUZl2T3LDo8mKFzzU
Bewd1LsVGQEG6efFjS7mNVlLy41KxbyAvaK7gCHUeJpn4XshA+/1leg4Hhww00QV
Z9fdwdjNurDQQietUKavfRdhOyFyc7loiJCscjGq1fHrxsUN4FRX/PGzKR9EpxnK
FKgIaP0U30G/Lfjua51e2F/PRuFKfb6VwB5G5uv77e5vVr9ZOwqLRNEc+KUmGf8N
JVXCjPZhdT+fSHFg3wbsBQCbBLPJ/2KiYOu8oB8RdS1UjN2472a90B9nsUWG66iw
NgrujAEoPG28TxUZwSgOwz4KrZD6NvTEaO5Fda9mzoHDm/2hiQ5XAIsLVCPURjQh
m+LccHboHj7SUfQjuhDPvTgoPpQ2lCo2DSYCa2rJdR0+7bKpmCXJpQeTLj7SB1ep
pPud3cvUO6oh5bu1qb969IRcYuLnQ1MT/BX4bdY6p3eKHzwd2/eqkFzsAvUPZ2Jx
HczS7iACQQlisMxvBm0msaapUA8hpy3yKEc0os7P2baQANMa2voIrKUH3GyKSnqD
RwHdg1yLBgIPMs+/zDn1gI9qX7uF+QQX5Yu49Y0v2HdtwR36gqhbFHU0chiEpli5
Vf6Zlt3B69/cyysPiyQtiQLadt+YTdm7WomQDWkfGKReQROyDI0z1sQhO4rAtKWe
WrTWslWkojlAORY2fneEiMTulJU0Gs9bmaiisoc9S22KhxP90JgahC0MUk2NNlYF
pZDPqUcGKyJDba5BmR2If+yEapqIoAnJ/AIFKdmbte4NQ0SMxCz9cq+VxN0DUQ4j
JXMhlgnPLLk1ErIc0PTWFaFJM5GVccRhC2a9T7F3/SsU3rzEw6ZM81gZcvIdgKvY
IS1r+u9NRhO88uUv3fANLOOzzXXlsoHWZB94c2epukDtO5UOTZp2aVVtVqUoKFy4
6FSRbWLXKwFKZZT3+PPmON+ees3/4w1IWYBLxVwXQ5tvS9SeLqF43mvBWSKnHEfp
9QBV0/whelPgzjUiVcrNQvvoLUaygiKvLDsOlAWcH4ttGK/8VxIwcOLClW2ivtzo
qB2bt1EuI/d2LMrDTBYVVUnfUF+cgQau4qFKOq/ykwGENrccqA9jK1jLX9oKQ/yD
wSNxxss0Osndpp1kpHSZQ+eMx/apjJPm87L0tnzsGlkBLq7fLIxxAuUoR/Q51/+H
/JEPdd71MLAhrEVWBU9j0Iet+1mX03oA0Uvl7GtBuIDCqUKnIP5KGnTT7wB95itC
Vs0DX9NXkHmlj6em8PHl5+QAYLveQgIHdWkg6eWeXyFZ1ljvmH0n+EFztLH4L0Fq
iW4ARYZZmJRIRPUkW7hjVzSlKnn/A0bqa+/ME7brNIIuE/52VC/0FjWIQJz/0hEn
xPI6jTITNFrqGWzH3DH2VGAuelM2AdEKSes7YS2uzIJIbQp36OtCoJFkMywpmQ0A
Zj0TIUREiPLgOUCh9VmtCmIEURsUFpnEO94kJRbyjc/l8yR2nypX575i9OR468kD
WyGw8wasfRXxDyrmcTOMbZ8KBCidvbDf7FnTlWh/bIeiQGawo5n4KYPivUd1AoZV
mWDp8U/h3sl/BSTIV99/dNVnzZ4tUiASvy/Ml63H8TYUjYPaX0lnrsWVJSmHCgRQ
G0SIGDGtQlPgwccrHfOlZoGdq0f6FEpAVVbTde959bMGPdVs5i+EstFmh1cC5QYj
s0ARg9vo2647KC8BO1zMVVp/zi1qwoGi8J7Z2+Vn9zLWJoOq3NgCpjfAPthYVjfZ
VKCeiaXcWHbWkzwPVWvFX2ed6IY2h+b/5aDC4YmClBtCkAE2TGrtPk1ALXqvr/ZA
1wAkJpFvk5i58HVrYVRQzkYMz3Rlp5ozjW2XPcy0FH1Rz0qvc9n4ufF93DyCmHg1
1sRneTuRtUSEWSHf+yaETjB39XHFRyXKVgqtm6nqasQA2CUy1pRxlzpKOSBRvbQ/
Cxx1WMq4/RVsRkhFZEcu46lSJnw7n3X6H4zX/3TT0x4QSfOdzemDNfGpmM3CgLkM
F8JK16126eI8l2dYQLizssOh3Sa58lMPwK4+/S/4UdlkOWu/UixjMMhWISlChq8Y
ciksyfSPiU+M1yHUOQ50nty/UzewqyQTgjI4o8ml0xMTl9eK8KkFuHXubdSgc9td
cIc2tQo/GSRxwajsMGvOTKPoHx9DQ+y5UY63C9m8k0eNvRz0p3unkMtQ4movWtRe
nQz1brri7gEdjkKremkfFZz48gK8DlW/oISA2utORsAgW1lypiPXyErBgTf//YFL
CBjPxcVQYHkMHYexrv2qDZ8MhcUFKOdO0Ss0izMyAry6snQP86GR25wDhtNl+h15
9Q8cW2upMnCZnPSx0V3vlDhtoJxjiPl7N9ZqZ1R8SAqQhUAv18YeTcBSyE+kMD9Q
mEgEs2uMi6Te9XR15UnFZvGTFmNiS6po7CfA5/uda62X3My34AYuTwcl1JvDWwES
FssXEf6BE81f0AzFtQ3KsPeAjqmq0QRNjgWtt4MxsHkxH2cWUnNJ4hlQgUHOTkNR
JaBH81NwPHrUYu8xA0I/4z9TR8pkPd30MhKo4hc8d2F200Vl21iIpT7L8P6vXT1v
cTFAIqaYfJvKuebNop7I2+yqWvI+fyb5EFuKDeLDrZkmJcxih8cF6LWTRNJCSNRN
ginxX9X7PV8R7GBun64pDL3obXTZgINHz+6PW0F9FFdx7pMBz/Iiy1tYTa6HrCZT
Bk6NecVGYCcUR4Ot3VywzQbD982klnJwqJ6anIKTMn8E+Z2Yo34JhW7T9JKTP+J9
q6L337rQBAQikgz/Z/4NUrKFKfc8kHgMf9eIxstvd4Bk0MdcltqgjtdMY9O8gbOH
US0YP59IursbUtrg7qLYAvguz+rYVPWAOIhryap+4zVrLamoRkjBPpzkCQDCwaqO
dxWWb/AYtTxIQFxQ4O1MthbMuFFLwjzEHcquKTAm/vHrATX+gc7qf45GIHic+gSU
eCAbQuBgONSkfYoVgn8VsLGeb7uagEFzVvXyrshb/7UQFdNDKasZfoOI6wBocpDr
+QVOg58SLEXEJrgvCAPcn4H86zAr7OM6+OzvATFatzdiTfTAj5BRud21uN3F/bYt
OsVHsYAmE/5UIjxp/rIcD3exnUhEyYl0OTgaLNtsm9qea+Ago9kxY9Jf8JBjADgF
TlvZKkX/Rv8ZgP5zCDPjfaSqmDugcjiVvEtyXM2kbQZ7re5rGrDaBpEyXIWAcM5d
RmBQMgSpAs9cu1T89nMwbEBEtn+8hpHScgWHCpJ7t7BOtlx+9YkrwTNcv2SLXrGn
ID9P/P1k0kYyOYH4bZCSXF92gxGHdg+XqizyacNh1gvzoktYaVwDyPUFGYRo+KC+
magGC84PsDlKABVrJyB6+dk2urjayoL+VcQ4PWZgZ1HOtam5B8zyOA6BoM+QYFoR
CJup+NuyNh+s+MBd8t6I9u6flzvLYdQJ4vWlWOuNfFh7aIfnnvcPcvweF+cXfiXy
KhdEE4HgogykYB0lJonR134pL6cHq7T2vBg7I6xs01cPXftPboTliWSWXgZFsZoc
xVtF/hSSFfeudneLgVwtya+hpsCxFXj6r/Ffq56uCofjQwJYMZthANIR0+m76GKY
5rjPPUL6+a7no1yOzKvfaqoBYvoUc7QvrJvr4XbhXhxae8kF8+WOBK/cBjX1kF/+
I1JNXK22qUTJoU5qeqTku8b5y1Rug3txGvePWvNttevv/knyNXBhAWdSBagEMi4e
dghx8hquvYJh0iK/R3Q5tqZT39BDL2+uU2x35NN3dh0jJxCm8oybdIeIzZKE2nKX
TTUP3mNa92a5AfIyVS74bomun88p/72sarBzlAgEQOTNzQgHdKdL1QGkv9MUx/Wz
utfLud5Tm+Z2EIKCdC0ZM3X/RHYQVuAegv+wo5mRtoH9rqnYuqOIbcw2kaGUvRhV
01gZATnXOwcXUuUE8q7prMIvY7jKhkuBivh86LkltUK8q/YR/H5udf4eXkZoqfIr
0vSjjac3ggyf3+F+cMeF8t68wDD54v005ejwf2EldFl/xnPxwu0g/yPYbyydBZav
APih+JWI0qCx5VHIfZSjiSfdiXCdJlhes8FPMgKjbad0PEmulluUhEgMPaJ8Q4Nb
jSA1ahsULK2TfA351e1P4oMDhcHnmxcQfQxZNSSmaH/vtBcRddN6mjF41x279uoy
5xx5gpwwG7yGGglDYrGo4NMZUsYBtNKDM/5GxgF4mXpIb+BHoXwm/eHLFGXAUK6P
zhlEWntDs+mlJurk/2E0uJhOMasekJFZDmARlpRMW+oKe73TRcaoVdn3O8xD1U56
qN1R3uC71Hb+NKrGQ8v10wjRqyhunEczncoRSDCN+aLf/5wbqaAFgDEabRJZSvwr
K+vzvcOrlhtqSjxuT4+dlsqtyR1MrY87gmfdoksFUpP0QV6QkcNqX6VCKRfLiagD
fCfLXgXx6i/LsR22MRlWC9yqvz9xUEksE8qQS5SelUo1QrgLIGVlnb/RH79eyXTf
cTW3gRkN2GmgLoUxBtu7B/4Nd/Iz3oJTiDq6s0AjzEiOSWCPXM2prxupssAImBkr
5AQt/7UkRKYa43bvHkdimx3CsmBVciESY7iwlvjucpmADslFYXsi58F/7bK34TsZ
7CjZbCtdh+aLVzjTKhT58fnfxGkCxnVy6sQOJ+r0Psg5V3ubu1lD8MVgsNoXAzTr
fzGwBtzsgB2dn2lTHQWW5ppYvtvr9b7tJ8gRF6IUWq+LUikf14v8X57GZV6ykFTv
bspxsnuOCArzA661GMIwWH1+GhN28SvIO/JIWSBBJZPdeVYULmcIKoUG1gc8NLoq
mleayYPYNVI7+bty5UnJOLONkoC8JJHr8sMKw7hfY9w+4MgWqd8EWQuEljHsTsE7
TEOOkmGlJ/+U/tjTvJSAybq/nG3S71pic/QSuds3nsU8PXO/XGVab647FGCKyoOJ
vNFTMreNHWyiumlU/XADIV3svOwxPbfmM4PKa84C2LoH3wxma7XAkQt7eZ1z7jlH
0CeWrVaLt1katde6L0Zemg94y+cG7cwGF1CiyskrAKqIVYrSpzdjqaBsGQUcC/Ag
dmZlN38v9PneqCx5RoqpEft0wFe30sG6sIfrvEufs1J6oIGH48Hp9bymuVtzmgNY
TSaQIPr69Ljruhm2gFEZljZsdVahemeDi0cP8osRzyXbeqBVuBJDIJqIgCsBqhJz
wWKFzhhnbWIHkJDeUHMseLZ34XCM0QBq5rPKSn9OJI4ZBaWOcD5dY8s5E4B5JyI8
r8Tc+bSchXk4Z/oJNrrYYJ0WiD4VA5FaFDbxxeL7GrUvi5+50isHBYjcMu3WsVSP
zKQbZjTEHHveH+7I4LqRqy7PdE7Yd4+AHL3cAr6GjsRoEAFn2OH2YDz0C/g/Cc5o
pLtqCR9K+6utNcP8GPn5fqQ6CyKA27OTIrRmrh0qiUUv+iPerQAtZb4PfaSb0vom
xageueqH6pc8J3osJgjG6vvr0WyjfcSbvDyQKLWvPFfyHETWyBPbstErcJoVqZlz
G8dpoDks8i7Kt2Fgro7XHQ7WIptFDAOSBlCiTX8LEDNNzbazltaZN5FQRGa8Du6B
N8WBxuPnABbf/dNaWtQtc1Qo4e7mpPdTQT8j7lAXkJ5IZ042ZjAnvxKrW7txvabW
lpNiTGkOJoLidb2kvPZR+mIINv9qvOEhVclsqVtAAc6AMAMKMF7v2WHFkveAReAR
o+b0cz0g4enM5tuUIWr5Caozw+KvPCZpeS/56/REcsrsBclmlvzfPzzTl26ecE5F
FxAg+nM/myFGjgIopmiu88YToMy5yN+nTzC9pixJTj2YExNpzvQPQHkylVCxDg/n
494WuYGY1eFSMwT8ApT66p90ugxld0X3X+FZsa0IlXZuqXXlEb96n9fpZepdHbCK
1QxNyXpZW01jLpyGpwimfe/2iUAxn9J2KmKioC7g9pmU/ThMkUAWqBK3QDtIZYpU
JOy+CAYme24s+Ogdx8+2ZZB1rJKOp1K3Dr2Xzz3p1ubkB/NDZUbBvIPfdVqhMahV
+eFWOC0PYqTyMIlzSJAwS2KicBT5GlRbKjLWue/rjzmwCpSjc+e38yUd7FGfgsE5
grMf5tU+D3gEQmy+oqJ589wH02rhR+9GlmPMR3/PDLTlkJb5AUR9vNrcLFCZTwbf
eK+MhtLYP9qAXB3StZHARLyAMUpTh14qXrnuRJNtjwD5llbwWv28eJsO4r2uFg3a
0ReiMsjcdx0xQkhTj+d8HsKr01EUeJ6+IBQPat3nK4UYL3c8WzU6uocihn1djwQ6
Albxptga1cckUPaVKqTMiApiKXccBpTVBLieTShIOUJ6zLapz0HfIByT0uN3Zngf
8+qQWWMyE9v1eeBY1sKD8ufmSek9TUycvN/QHhh9NW5D5y1L64v+WAbrCWBBeXkA
WVi7RGqH3+ZR8PNzL9Z4ON/o+v3Y7rUpkd/bd48jpA3Bs7NjALw1U4WfHCNR5xh/
Yk8xeJzSmlivFGriMmFQ7w+6Ts9evJGHcbaJ7O6mcONiAgHgctc6AYwI2Ibpbcmm
rAHJE75tv+rVmWAGqnPKQAKoaG+Q81rbR9F8daNfjstH5nJLbElHb/YBEuOjsPh2
SY97dSQAmJML5u3saAIefBZkAzZ7skGHGXex4iQEEQNEWVKYkY9FF5GDskE/HUdT
LRmgE8NZ+9OD2CtKUzYAxryievi5K1ZpNu70HwpIG5odb0wbynKhNSDO+IJ3Os2M
wjDHkJKWK2aWgFTwL+fjl11fQORRLeX2MlLiAkFKkHQhV6/XfTbHRn6sigdcTqmE
olQ11STGnqJjLaTYX+wVnjf8M1EZQAN50HHy/Iws+JdL78WCvLJ6eSzzB1KCTKcn
j2Plr+dsA+gLOzcgbdD4vH/YDrZHAQOCHYkUQEEwabDVYMJGm7QCkC/Og3sRXOiB
48HqoRHmsicnVgVhO6OlVr06c9+ykj9MFq0pkprziisqlTiI4wqpGuoYbbaFiNOO
1BpYAyp4KmFjO8rSTyCU5dzP8jSSkNT8vGJjCQYoFd5woaKDy1PDN1wzv9AliRO3
dEs6TYQqYx0xMr6pQP6GLnDnITsnxPic/Y41vZ9yt59Snh6ys1XaVVnKZ5xzUQ/B
K4oeX+mq4yKFfuWRQEY0byNS/JnjFZigoTPSoqYgKd4aBNzNJ3qwDouSSwhQ4rk9
DixtL7F/EXI90F7RLWQwYIoqp4X1GUVGs0PTb9UjWsk1CYc0CvccDZlb4Kf58vmR
74dVT6hql5eFAyWf6M+euRXdKn1ByKIHnL5hXO0pw1XnDsBdgrYDsc9hruzgWGuc
MOWZlcC6dns1dBOkyQvn3eQFjyl0bj+DJtGyIlM5ZL4UGdnpZ/CgSVWFtDvKIPrK
y12PvuKoH4b7j/8gfx43ZTsjdWXPtHTUSAyZDZdHJu+bIlLpfutFXTSJu5e4PTKx
EV/lncTxFdxBqdlYUaKkvPCqFmZT8WaWTmLAwkjinftW/w2ChlnvHZK2yoD5PDRe
Djbl4OZX3DtDZfYTC6u2RKw8KsPsnVfx++27EOJ6z7fWImTxYbH8VJpsNXBimymZ
sG5PYRfFypLS86QN4OXDdPvndt8cHZx9CVvAuKzqTYzOuzeG+IC4xTKZ8AjmFxkY
ifi4NZEGbAFXwtexafL7Pw/uFQxpXof7LDvBE7y21zc1EvoVBBJAXFOnWKry1Oa7
gdkr9+kngeKWkQMi/yndQ2SnUG7eu5UGrYSO0zWmXeFVTobQQxNoDjTIlSDO/1fC
0URzoPg9gl/UToPrc3QFMl7xF3lMCDIVpUnBoZ1Ee1BBGvsSV8y1fTI4BVkhA1tE
DLbD9RnoZMLUXPuXgSNlkqd1mySfeTbdwoz6B3kg5GcZ7WazIXTJr8oS9wfLh5RH
rnJuQuRnH8AYueLa4WbkkBCLAirnAY4O7omcnkCKoTY3bFQKVKYoOAVv3579edIJ
Ri7PjHp/ajYXsgAUN6TY0eoA175YYleB01VND1PRPBr5yw/ETFW85rJ24bv7uYvh
nujADH4jKUiyUhJPEJMcAMI/1VHVGdRE6MMcDgB3njYOSF3ATlFDMW8OGnRtnwq7
mW8xjAUkVIr+9VIB3UxWwqIEECYeBbaB0hDFpDpfcgmcVTMz28fLbaGFJobAc8jL
7gEb5QnTNKjpiQ6CauPRJLalqq3WwUBzjmjJwZXpdxsp0R47c/0A8sZcASCrCySa
F/SSfvzAhYexmeIaejRjB6Nay7yGwXQ9pxUZnyTdZMqBpVoY1PO/rt7I+CqUOpaK
g6Gb0MCuHWg5N+ufY9LwCjKkSasLtsvlFJxUNx27oPZVyVVkBkOXvJ4k+Om9stA0
W6IN5aCCp++HVOO57lhoFTra9CrUTtkns6FCIT+IrBoy0IxJGGZAjCc6k86ooolP
i45JXval/cc4L2EaXJW5ja2goLpQ/qjvLS/RWj17ko4O8K/MqV7hG5mrcsHdrgKb
lDKyiq7lKUIviE8rx0wNn/nav2pBM8q8lOIfKOKYBkoI6KZQX6mw3ZewBsBYZJ7T
4EvlIdt7elzXYPG6qKWZ/akQr4I1O+VDXMcK/7mur2I/hvloKlgiZQzI5GwTIw2x
ptoQ4CuWXV/20n+8eYkKnVkwdpnkwdwW1YGogjISoU4+TOKdNgpG1Mq5++Qx44nj
OMPw8zgEBXM1Bfhgf0Q5Bsvqtm6ORiZURpQzj3CQs3CjoSDTWUBp+f8kpIF9MM7b
OTe3yKzucMMGhY1tIpLFHZFDR/aBnc7kmUSOPuckjXg8cIo1nJNksa/KeNNxkI/Q
znimvb9IvpWPq91J9gE9Yd7iWjmBrN4fsulS9BEL53i3zkOUzlMseL6ghKj0GM8r
55pq26Hub9Q2UQEadWwUTeK92emCwPzg/t16dwCwfTZdWnaBXxO+au0/X4297MSM
cip0CvldPc4esTMZVk0abMPm5F1Rc7eGlRHpa9d6YR4di0kL3Mw48sG3qRqJujY/
Q7ruAJ40bD8nF/Oy9yaLgkeU/6s20qKo/OJSm014XDBw0QGFI1IlZgCQtsthTcRj
U1u0CYhTwe33f2Wdms0XupbMGL+vonklKj5k8uin0QpFj1whdZoGP2l3pNpkaQis
lhE4TIUj5suhaxN0Xeu3LtFomkjp4G3UptzKet7IN79H5M5mgIBblgx6zBfEhbBu
2QTlQYE2afauVYeVcNC6gIlTDp6RgoFX9eBwWUU5bBrW7IrtusgfXONP9bXTJ4YM
3jMirWcxRxwhHshoWvBv0Mztl9DWco3oqlrT38UVoSWDUzKXvHpOmtrhkiObDQxo
uzfrQIs5LFf+uDAMspFzn0Ft1twojg216W0k62V111kyYm1BKoQUegXfNpa8wXJY
Mz6NetzhV9BJIJLgzsaqtdOPrwNdNL4/MDXZ/DUGtUuNk4nZr2BFI7s9Cpd1p6if
FQ1uGo7pBWILKytzWbS53LLo+/e5AA6nHEqwFWvJqJHLPSeVl04bicuGeqMDr9oF
Gs52c659RTvG+E2U0M0jxd8ma7dAhMrqUmHh1PERW0Ub4i75kdx8ibCeu0DLp25r
aiTuZMWoaptamFvHGC8cbJt0Xoy2k2pt22RfhjCg3/N4TaBAwMUTncwjHUglK+Gf
cBUK4U1SxOt+Y1DvLtsweF3biHGZj/zNpf3OjJFLhW3RnDkxU/SwssdsfLZ9Kn+l
HKBca9G7KdKFAwxLBr6SKUjQa/PUhSZSFTiv3jLsF86RTyl/YZBzW4hncP0IlG80
QlBJa2aaBcUIUlBskrgyOndNY2zDJgwr55nRzmtA3x8h93ZTJixZYOxJpDsJm6Ky
0+qKLdiMR3yeXbR1gj9iowm2JQbA0mAgILCseBX0j7ZG44c9fqZi0N08vAEgkmp4
bZKtHPI8Pq5uEQmAoraVVv+1fNuE9/lI6jTaSEZ2RZzGJhga/Cu18qfs70InO2EY
55nHrqEPtVq0+F+isBXnu4qDeSKrkiVVkOfzjZYj71WxLpO81YV437rqJ7pvcx2y
gSB7NzjAWrRAv+3QLWSdN8wmiVbhrKXSeQMcnSYQSGRxxA++UedQg/XdQS1FHHg2
AtzdiEpkTcDUe0DXB8fGyp/GapK4hMhT3Hwcqe3v0mG94mxl5S7TIeBWk0P4KS3A
MO/+MZXnIDK7dCr9oqAm3lAeD/y6AbKAUgBdL2KANwcuzdkBtvpUBcAkJStSSd+U
0d+1CVL0l9APRvl6BRTW2yYLRfcG0KBE0Ik119/NA61fE+UK2q7gkwkLbudYCWiC
w3oa+mvsS/YvPBMoJKhYC8FUqIkz1olaw3Rq02H9aY/oAQs6CmAyOj4HNoaH3jK9
00qAdneWoDZ9H//7askYGmDdFig6Y5BKTQkwdTu3nplBiY3Z48tH3ODOBkXrvbIC
1PyrfLQNC+DL4FWRa1XHkYnUdLju+OErD2edd7Q7Yfkg7A34cxbnkjOxOJ06szgk
SXaQnDVC+lItVbHEehzEBVWCJ4/Q1so1Xvmj2fh8PvB3mhKvR1HwJeFjNb/vYKEE
fTBu0S3HiRxbFs7PQoo5AV93aLuMjoe/UaKVRDkp8SwYGBYfwn9A8+vLEMUqkVLe
ee9/37t0VTK2UT4xRvjc4Y5hN7KzH1VMB/W6LoC2waTygNhlc84v8S8ycT+LXans
2L874XMPWiobCA+oRxojbLHcFz2+FBCI3CFWvs4v0M7wV2n+GoWy6Xzpp/EhIn9T
JG2O4Ao6lxgRlTZqd82ZE6bGOLN43nl7gPBBDzbGtFNFhKsjMK8eEB+TOqniYy52
d/rdkqlf42lp8lM3k6eTzvwbt+x586tuv2rVYk52iV/deVF8vGKpYnEDYVQwk58M
ivKe1vQWbxdQQxE6I7VSAPncONow8+Rdant18Zo2IcQGn41yVxrcZ+vOIaPBRLPK
Y/737ju/V9KPGNMltgcGiLDFkreagSh9wVlna+DYSFKfkziMjunNXSUpHnpQO7pT
conKZMo5CKLp+Bw+C96J/Lv+/n93VW2w82LMHVraXI3WZIuIt+cTWpXYjoAgz+K0
yjb+BBC7reUmAclEMDRTiWBD1vUbDB+N9iuLyHleJNBF0Zb/er1O/1PAGKm2RBuP
YdRIbBUXorby95aQy6aZUNUMSJEwjSnPBP3+VGLYHGNmNhxtNKMfk41N8Hr6Ey7/
XHllYr9vY0rNf9aDrrCeLUvakO4hQipkZ6dJAWqLCmsvx7KIbg+tWtRtK8U5rdW+
7AQcltR8aFvWL8wKHqJxRpSkFJJ08acVY4cVsW9cbByfzjekjMsUDGVqBvGwd22B
Og3rVNlgmY2kgkOB5HrcpUm+euErRzBGxZZPV6poGf4GY+d+FKCRjclTh/EXYIBA
OJPgMbDI91/egmRcYfdhU9hlEProwi2RVfyaiUMX3GlxagPgU3TH74KcG0VB2ynz
mydUu3SPigwJft9EbXUB/qxFiszbCGz4AK6o6fddn+qtXN0UhqCkM677ttKZpNZ2
1dCfyRVDPGYSVBIUGaDRdRijzBxmcnOIHB802UgHZQvkccVYeJWCgqg1fdEWIucD
TR8Hbr0dZSH+m9IR6vGqS4m748JV2xssE9F+BXpsZc8smY3tZBN6co57bFom6ZhC
pnp+P79PA8htf3s2AYUiRpI7aPItEe7+UJyhXIrbjnHdmkEbs8+jj+NbSC4ItGWa
nAXHzDFiSVYCEkHo0BAwC8euXp0OY4ozZzpYCSIzp8nY+NUWVfRNSmUWUWMXbqqf
8vk1kehGx8a4jlgXNhZ8j0mmrgnWOXNl6xp+oe6reUWqE1R4Srzx5SnxZcqUaLxf
+N/uhPx0yxpJvX7zRSvqUXTwbm/zMfCJhtI6hBI45bw5HqTbtJRgL1CErOBCidGE
qOmca9QLaz3SZcied47/1wbZ6QoxCE+ZQrvV8GUUlFa3qdliYqEJEaJZuli6My1r
80Yu0CfF4nRlKqbZbJJrCAgkzGugu+sBCWNxl8hCvD+WXgjEBppbR85OpWgbjVx6
bliCarz2BeVt+4R3gbEiLZeppWiVjqiTYjWfWog2meHKtb/rKZByzFrvD8sveXz6
TW9BWow3ylwku57neDwApCF9jyP81myX+Nv412vN1RsTYF/p/EByNf2MkoUmzixc
9U3lOosrUTJ0u4ixsF17IXDW4tjeLfN8hXHLFuTBryR4e8ZB7xbWwSje/CIVRvUM
gCZ165r3lR9xZEONOGrloBasPFq7Oyfw/YGUwwlnnUOj43rW00RYmZ6xzLdwEslA
DkkKSQFOj6lrtvbhvbZT4CZgq1cGxHL1XS4tFcDRyiV3PsGQBQfXJ9zihgnnY7nr
+XGf7vqA2wAsSZwE4xoDfDdZy9RE4XVe18U6Zg6GMqk7ONdyAjEPo5p/qnth5kko
CWZ+ZuIiae4+rMJtCTdb5F1G18nf+siBnYvKCarH9dyoMeMFzo4VXEJmbymRxiuk
F19qt0hyiVww2eZBPF10aQa6j+gVD3QFpEVl08nSBCmuL7YY9fPL+yMWVY7k++mS
Mm2UlABbWSbdHFHMayR71uThF/we3/mYWq9PhA2Saaxs4DJml6mDlNp1xTHXB1fA
JPJyXsLcCv93vDd4qQq+cI4FAAY4NZ/LqKAubLNanKDs8npM+7I9EjeCjcj2+8RY
k0DHJgKtLmz00wJuqcwwiNjzKUGcaD6zcD1BMLNvjqJiYtg1+j/Xkk305aIY2MLw
RTTW2PyCA2073RWstVRH4HWGA0UgNnP0XWI42nATakgKYHuArLt7TBzVBovepfRA
tK4lG+t/tLAQF+r7UMV/ZDDQf6L6URk8GRvpqx/H6Ww3b+w4CVsX6RUEet5C10di
XxDFRtWlVCcvtIs6y5h9SY+xQWT2mA7DbSNAND0+BYYtl8TWqKwTslqf+073nmJD
WnvupY6J2hhNV+UVWqEDaiFLV0QluFCcSCBgHTzui0daVh4sOpbSziiMh3WzVsIv
zEotKiJCHkpRwKvg6jrsTv3m1+/TP3DRaNBU710KeK036agbiOHgvz0+8uDJj7aj
hvbIOjtlET30k3T9QvRQHhqRD/p9dBRhmoyFVoXZiXViaUhNx2gFrsVy/7Qp+DNE
LJ2HjYXfe9ci6CyN3uNLJGosCMocqLs6YrRct0HWfK605aQKZ3xVMqTfOcn4/LdI
62fCsiOrI0MB7n5TIfTb9SBsynOpKSKGRTiie43k+6AiHYDT60ZxM2RbpHvnB8AH
368hpP8oZa1gZMrIyUp99RYJEkxb+VWBN+7Ixh+98hL3IoPtWTQSpDYHIRBRvlO9
xpDiFXiroBrpArYyAXCtUCQlOiYypbk9PCbGQjcWRHAqWnkKn6eNmFN6VcwpUD7T
gx9XRCzxobyvrN1pp+fKImWfHtqhCOu2ta/YCb6/k1fxM+KPkweHYa/t04Ghyepd
A1u04+dOx0NLOmh4pv6jnjHxxYGZpOCxwt6Px3FjKVsCYyfheGO2VFI21Y6jOeGP
tjerxrqrO9wH2pzF6gSfWoNeF6mxrvPA6jIrcH/GuAlOLTlKk02IK1eCrqSlT9ca
lztlhneIz5UEMhVcUMeKhTkdGsFAQKzEkbLxgRUONCw9mkrr7A+6Rlm4jjB8PXeM
+/oTWI0RAQelLwDU1DU20qytAR44N0tBkotaY0Ad+1uil9UEtrC0ViLoUqnu6THE
OS2MCCzO+USCyMzFuBO0gytqIllCMPsu3mS9nYO1GluYItZDhJFs9P/MThKJcxic
8fEw8c9nyi3aJigcwMgU7h9pJxG3yGjsItDpKLUDbwlDlf55N9uaMCLHCnQA0Qhp
Xuq3IIdfRhojmUHEeqYHDmGSzHKmSKywDqkIhL/W1UJU+RZaHUXZmvf12IEP80bG
hE0nrP1sXcgxL8cCTQ+3bOJyS+l6/C0FJDizpbs23BIJDMatHgn1nk9Zr+NHpUdV
+y8447CTR9LW8fcWKPOtpqM/9yhray9vgguPKjCSVOthef9U6U1wo6XXuuG2lNV3
NOgt1Aium2A+Djn4CUkA6ZanHlwTWxLfixaPBATM+o6rESnp4O7PT3TffJ1Czp24
GEZXvZpjzT2BstBYHGWfryrgDdQ2zddH8i+nzjQSbu3Vv8gwD/QQJBDm/fLd8p4K
nEPF/lGTQnatgdQC+OTjms3I8vi1jIXldBPKxDuVtwuNoO1uA+5LVv4E2ymGp9Lk
uxvphM3nQtgGzOf+GB50YwlyXJ/jLxr4ZLTKPBz+DxdDA10D+GqGT8VKKHH5Y5pW
pg4S9gnAY5yE0e5JIzI+C+5t2kSUpMM92FSv/8PYwIIhtagU3CiC+lbF9SzsoskP
n4M9PjvGNqbQsa3H4q6ujrs33/+bWz6S7WZf5cpvMI8SECGDU4IDtIDsVoNI4ECI
7dqGIWcLWCfElxWkdnte4CqPmL60uLlT8sZC8t28ocMamY3Qt2Y161qXjNANERMz
ZfMB1zE6cLfX5/r0qemIDnuG7doiRNnQiy/6FCd9Qm8XcY7WhI9NRqQ2Q3ffnc1q
gy/V2gx9ULqnXmVbLVRqAp+qOZoV3USZrpxD7BRdj0yjZVLp6JO8gLv7XFcsHogT
DLLXC3OwPATZagE2j8fRk4QhvhFXNrpD4XZkXY932/oN0d4cAv94Chd/FbnuDRKr
xLueMI+uBVBsZHFLE1RXU1l9daFbyVio93O05T82AhpY3eZ2Ox889Mbt6rC7B+rI
J2w2U5/9It+f56RzlPeMlnpSwxDbVmAW3JzZTRczRD3X+nNP4UlfvPu8kh4vxldG
YfqwXiWKmPvwJ/UzS8caCDI/xjwTTgLnZYDDJ+d2RZBUBTh5IW4jHigTWgD7P2z1
ab/poy/EK7Z6+IjO6YZ7K1S5RrHyeCiO+H6ucsXkonQ5if0k0k5lsYybcIo+9a6e
nnRWTVzugz6ZD7Q3Q+mnmOhwgHYstOxL1KDEelfedzFGLsEZbvMURB2nlmnW/KtB
IB+4xG83KEYpdvrBEJElCUIByVXmTsy1bKXz3nOL8wztEUrUFYoYB75uWW1KpIkl
+9v2KJtWI/GUXYq00Idq/leuFDCNA3uu1spEAjgf0CZ92HfByg9ewNWzYJhmT86t
SRs8rLVjghyd4RRqmOM4Ji50gtuZqbG49thMMNzTbSPxQrYFCHcBnToMBX+OXp5v
tr5LFOsaccGtmCaDtitERwiwT1gnXZnzlftnurfkm4Qk1axP5Ip123XQQBQvEy0h
u65Jex+t+6ziBi7J/6RVyRFTHH/ozekKqf5NtH1JGtImjyh+PL39dXXrqYN9H+g+
JWL8dmc7lVfZyxhfTb/cE6E4zWx5qJoPIBe5KclZIaKxYvaQXHvykD2WTHr3qNv3
fOcXDxh2Ffqo6PkNhAabtddUv3FCxseLmcwJzj6eSGcwzZLUiWK39c1LGFQmINMk
fHELCdtWYFP0h+cz5XBwiCo9T/rZ8RM7tqxvfgx4JQU0KpGfbTuhUBKIAFlUenn7
0dvFCUVHPNdPrK/7M4FFD24O6TDBCE7eGDRlnGtlcswzOlJ2suYa7ERK3caPFV1l
nisjP0bdAthPmoc/fzMr5GbP/HwvGkxZR9J5KinBjbAb73xy+BzYLqNt4MjxnDGI
jNQvfV9zIiGogFoXSe6jbwstgx2zxcqUvAji7KM8no1mvM0BxBj9sElbUJaYmj4T
+OH53D61y1kwmBp3iJf574AwIHAPPrOvq7R8ezJONv4FqnehSmD61uX0DLkxnP+o
NI2KdKcaTCKhKowu8FnDwTr5BRUVKH1XZBrbyfvZ1EeERWEmtPXboPZFipYURcsc
CT+tCXYkLyssChZC8Ii6bG/BZT3SEcMS76/ijDayDu7yBSWVtO1/x/7LAn4NN5O5
kW6jn46NoWbeGysZjebHfsnVjL40pb4SMzRAEW8scEKp3/rSh1e9n2UDdm0Ws1za
IcGIQ6A91r7TEXSKRdz5iYQ43woe58tpi3clBzLPrkSdgyAdvKPoKLUxFvkYo3zK
rW2UNOrGPVIA823bowfuTvMMciqD5IdAxaCEee7W1Vht3+WE30enaSQHpJnFaioO
5XS8Bl29vz2eUsujuxe/up8LM8AjwDAfll6EH0zdFsDD63TNzrgybDVpLvffTjYE
sOvwq+rpSEJBIETG+nn0yGVF2bwQXJw1/dGBLmGU72EMCzjNj5+hMKED5Hk4IOV7
8wcX7zobmHBJjkW9fvDftZslk8BapAMr14RMI+xznF4RbcLfXBASn3D93NN0U3gZ
0qF8qU73lNahA2hMddivwfSPpPZSyRRlUbIwTxfeK5fGWvg052G2JHsP4yFDZTl4
RXARFovMp7UFcSH9QrW5NlVcFbCw04ZOXpiDe35+ObAYT1f/2SoG7g5JKfX2K449
PlLgAKGIFdvRLwaGw9sz79CdxVV+K+sXPc8ilcvkwt0JPMUFHPymNnWZvw1hMVqw
cP6z7YZtX8llicapniZViFwpgV3zRTwbPgtCfEqTGHSscPnyss1UoiUxtJhfIeKy
8edYHfsL8xDANwrLZlFuLm8AAR/CVjTlXL+wWMLOk6TPKtqKXGwjFJaAciOGS/ca
LPaQ06tZSDlXHZMb79gY1+Tc+A3+LzmeUALMjOkq6ifEnOx102+CmaYTKJRt3qe7
PQUzuYiOHRWZujOCvHD9ukrBsbIt3UN4XOCGnw91Us8AVoEOTod3izE62ZeWsD6O
tVIL9h4vCv/+LWRFyliso0L5W76FeZrZN9+wexsTjGPWe8EYTkSesp+UKus/sQxQ
IDb5Dgk7JB10fGCdUgM0Amh3KBhIKNUkRbJKyw4XPgswFbzlR7T28OPbIDuHgwrx
/sxD+8Ad7GbDi4GDj6qItssV0jZlEUSE3WRGVzp72nf2dNXAoYcQG/lTc1pMgS7m
7S79SMEnXJqLLt0lGH2uUEaBOjEsIMwLELMrE61xwgzKctGh2mbkJwTVcTmk+qsN
OCXT1R2oltaEQiEFPWyNzjqD/kBaKfFE6sbrAl3T7PVg2lbWRPmVt3VlPYIrAR4v
rgAdbGg6Cnoi4jMnfAV7/jFvN5DN80V2vqUQUxz/e8eY6qyP1fJmVUt6HBjSNJR6
wbgCscaiBr1VIzxrdmIweC3NFMgDQx0XN1aemB8IxWM22FkmbB8HkqdiVl0AF8OZ
uWPNXpSdAzvzaVLACUhkno9DZB3cdhSn2Wx9cfdxpi5aGVpsk0+UJ8eK2jdOsH0l
wgg3Y+zDS/KRW77HcmMYu/BvQa51+pAlMcJELdpWM3FYmYozsB2bi7YG3lIxCptT
l69xTGvJl6gcIcuQs6he2/Nvw1kulgmGftbO9m7HUZqcdwOrdJj6WzFrFG3GMlS/
Xn6HOjY1r38ZVuN5NjU0DG7vntsxQNkOmmJaKBpmIqS/E7h2PLSfpGe4ln8Gtjmi
uLnMX3p/f3BMHe4/GvfTYvOOAuLoBHHIBsKyYfEA2zP50V7x1c6tR/RmRAgBtz3w
vup0RJkuTgMAeQ/B81xv9LPaC0YKmnpt5nTg1uXcK2y35cmu18Ax07RRA2DAooeu
zmq7W+YbvbQ5j6KqQcRDuzAc82m0NvmxQGSf+Da2pPgcRjXwCQsgKO2EbKSLAeX2
cRv9t43Q09B9ZiuxVt2NaVSnEw6U+IsSpbznSwJ59FAQ4uHprUGN54ceya17nrif
rW480uDyFPblyVNs+U913Xai9qmH+hI3dq2Vj7ctTEkxGlEk+Vt9YV/Gms9WbDqk
miJJ09Grys0Uj5a6p6rTnNdyMaotwQPD2D7lWCIeNFoab34Picx9pNuwN97+KcfL
jq84F+myHNOTJWq7iZ889DK+yo2aai0bnv+GOJvR6JdXJtpiO16pHDJNy9VX6AZh
dyjzXr8fHL0zYzso/w3fOsI7HF7i6+zkHTIwZPOToHsLhz4cfC4HN/YW0lfJDmK1
U7fjElo2OgYlEY21ypczMflhQZztHqhoZMkaEV8Sk9q5rIuD4KaZkoreZpe3ei6P
sjANdk0U6CiwzuCrevXqU5rZzvwVNwYq5zGGmcoOvR6HmE2EcyUfnvSmWe85ree/
ecvoA1UiIITURjDSkzj3YJNbbCUBnHsd+Fe4PwXvNg3lWiWjFbOZDz+Q2pdrdfla
3RSZGYdAvLSYmCrB8PkhzjhZdal6B05ppchrnm3HOm6/BDAf6OmnalkVsq3LLrY8
NTbJsc+Ci5mhWHKmGuLv4mLYNdopYkN6kgOPUjJgWyXgDHhLBqTBRXvHhKfHPoT4
kUECfDiEUQgHJCoa9UYS7/1an9PRQOr4fJvBAgXxi9meQLYYdaj5OAFMbMEC/M05
cM44NUIsVfoI/yjjOvYH6uca5Sjb9pNa8YTjgdJupNKxRYox72cNH4yZsE4wubh7
Kezw5JNdQdQ0yqOpYIHe8WBJ1aJTUghcnBpuyNpn5ILRB4bfJ4SKt8tyJaJoDfwk
z4r3IR91ijk8sAAlFnF2ROUbkW8NkPFxO+101FEZZKWsJkoSoDkMlauQ+zJ/xQjd
RauNPVhiU05dkKoH6qwu4hOblGQXStNZXVKjL9kpo7ZCrLaYoaHE+6RKd801D67F
vO+ugkRJ5BWOzHvxWfhiuZdcycurSAiWbrAANEGlsZ36g+HQvu7YXh2nK4qzUrlf
xS8k/Y9Jzj1WOJn8FWhq8Ds3XtmO1a0mnYr+G6t3kZtEwZ6jWidDqC0ADgo5BTOA
aYyAvPbiFz7apOpgMAhCIywIP/GE0UIzr1pxbYT7VZ1Ka3pusPUov5KWmgMcWt1I
9k+7AMnF0BSNOY6ivj+LjmZsFU9CYd2NK9mTL3oeYdhPabaJ2zrw3V0TiLQqUgYV
26IkzbIP2j5JKSn6PEBEIH4KAGS96PbVrLrz0FaH0cDCy9qBf2gbic0Likl367nu
GIffe8zMSYkcV2+2ArZp1Z2fzAo+Fwg33o+SL5qlBVYZ9yH/I1EDByCqQFUzn1Jq
IC5maO3LWOgJwz9sUgJnbAyr/MTtOm2GPTPw+uHVLX2C9o+80g/BBwiXAR3bQ7O9
KlzECDinYa7N2azGwEagwn0q6EHpJtgFNel5S/AR53t/nrX+uWEQt/ByLH5KvuwZ
h75UOINYatN0m8xIYj14HX5BEy8FkWrbhq4liRKA6tDLY+HTtosP42dKdHZLQknE
eHKzszhU66BGEUNK5cZH3za8/x4o6cIisayuTbciRZ78lYiS1iFixNmVkuFI4zEl
kdoy9Sm2hHplGUerIrAP3AE26LePxWna4pSmQd68aa/ghqBBmfDBdgYJ0hkMKhmn
Je+/n18DBI2cAy1/PtSB8Wz8PMZqw4vG0wp1skV5Gh07CTiTOCaNo/KH6JmVjHqM
scIkBCKvkLoJIJ40+2mBoMkl23deihPSAqTWFtMIXTf9MhO4KeLih6XujY+F3NiL
gYAEzNaZROoUAAgvwIRmOMDDb9Q3GtIW7+DPYwnCqHfG8S4L0CgA4kMx/iIW1fS5
SyMcsPQY6IrvT1lIM4yk5BeY3cGotbul8Q61kHDYsTqMk3tz1zNYn/sVoqlx8IHM
QgM6u5AZUv76/m18ZsftUSKsOg+VeKO1vXqgscI28GGh8dQ5HgmU33aqvSLFhDz4
iI0ie+LtKYPXknIznKE+EZp5mFPdqdmrUODnJrn6MH7zxtuEzfFd90CkB276Pir8
dxZmOKLajmyf236PWroYlYYuuHuF00lIqru8bTbh5x3UGAVZiMQLKH36CNusFvNa
pV3kJory8eI8O6LYf4drKlQaU8bPMZEyPZXfZTGf/IJvEtdoEJ+iVpYIVy6jheuR
ZTDDk1wIDys0IEyAxalRz6Zf6UXvX4LzCdBngN1+hx0QYSmtOQxwRExiO0830M5R
eQwVwoqCx8V2TMQ2dOwSqIBjQqqV68phYGO+pNDJNv1pIGN5kA9xQMjQVTqu5Sf+
nGA1mRwUC1l3LU1NajQIHLJgfkf4NyME9dnZ9y/Ul1Bi5dgmeYEUQTQJgubX36fA
t2VPD6P95w5S3vppQdmE9N8PPHdLtyBpkCqCqzRfvSOlMtHhXf79VZECzKPCVA68
vXr2v2PkD7/QIXMqv0rD1M0RAFi27aRi7gxRT3k2Mb1K4F/9h1/2jBB7SuS+KZf/
vYxYc8zCIf2jKmBVUiVHvmJfS1ozbIegal6bWES2JGhH+JVjqNW3008QtJspe1Uv
achQgPPpXgOKI7Smw6zRSZsEQpgYu4CIzeJLIllw2JgTe893t869EcZt8vjRWHWD
edOrwSt4c3ljY4ACzoJ1DHWm7xHzPwTI/ohmOrp7Wwrb3Fp4VjzZTxldjNK1D/e3
oUqzNAnhrF0aUXdKopWiR/zAZ4P05k26E5wCzfYtHobxsP4p6CR2LJ3LiQSVpIzl
5DE/zgMfnzTdlWzO4hQxedg9KOjV8jYT4MAaudUi5kuqFHJvA/qYhvCuS/AxHoII
oGC0ZXZv49ZyLndr6x0D0mO+VvRLN9UehwckA6dMSWVjxJMUy2OCOnYXBUgMHxrr
SHEgkbY3dNfhCzbfFPgzDzppgAjWb7tLvYsVDEAVGFUk7gA9jEvzcLuKobp9WwDn
w0x4QX2s+/D+zjT4H0uJinPIDGeprj3mE68SdeNqpp1IDRV9DNx8xXWzueNV2yvw
LcFpCBXYV6h/IvnRYUdo2Gobb72B+SNKvb8xBIrHD6rExNZMi9jZwcuEpOBF5I38
5ngmjIIkcF6O5AQ8Y+AAVx2MMQuDV1h/SB+g6WOQJyg3sQVwGuH5gGXHuH6pP349
aA7UK4WjPksdA3rEJqT3mGeR9M730Yz8KvyQ0IDVH4a/y73epKwOaiuRH9iTVaGM
h6yta0eF68lV/pVFwqD0QhgXQ2nnU1jTDp7ANY0WXDR/G//swue1eaSUBB1fJAS1
MHp1dIwKGLprx+ubqAHRE7JGu8iZpa7VOq44IMJTqhtWCdrm7prAJkRdwOQ5XvEl
LPe+iDt1hE+0tp2Ymj4Dq9R7mwYzx07GYeqeTiCm3KA3G5HY98WSa2aBVymhOgde
uPabePe9sJlTZ8JKrl3LbBEPI7Un4LA2OuPrDv+kNOp+k3mWau4rTkB4OQCqitoM
jdn8p9RvJgM7BCH/KBj+KaBgzw9bEYeUR0KHedwtfix3Hh/f0XI4YkLhfSxo7SPy
upkHPuHeI7X8kjSFDDTE/TJ+BMlKR9tqnbIpj4NinspJxwTf2+2UD8jC7H6W9CS6
VXcYKbEIjE+/nv3VhUxeNMqIBnauyR8SV0gdBBCSbl3E5/U/Ab5X2ATws0aqT7Dp
aRxOLTmQoAyszEQ5B7KNOgKye9PmVCJpZ3SKlsRl+aU7Z9F3T1rt72OUA677hMU4
BMy1gEfpP9sixLMJUPUDQksioY95ANoMS3hF8F7dlAdt/rwM/W1LIOKmKMbHzGEI
wePGnP6v/MfrxPQS7LMES1DfjcWAczm7nR6YzkFA6twHFOUmteHmBA9TIrFOFQZz
bzs4vwuXFoqwHkoBEuPNnnzIjwrnAsLlfd2Fbb2+aReKBcwdA5XlhOS6C/YTUhDl
pKfonx9pOwgNZbxD00+B4Rd2ATRps/ah9GFN3MzMOiRuNhgWSnEzy1OQyZrZxILJ
DVrl0+Y+9IGxQNH5aoN3oB47sFETAZ0rn3n/7g1FIdJgbUYw6YOrbBOpw8sh6ekg
dnt1ddvsOYZtV+YUit24H/klqqW9j8UbkAFqBRyCLa6cKQCf68Xg2NAWPHh/4oiL
HgfzjAbcDrEUjbPnPu9kyKwb1wVsJHQsOQcyGJAyBClMe2AMyzlVq739C3gptUmi
elltuU2DKbqCgFJgKvSsZE1aHwTmC/ncH8uEmvta13fNvE2lDYbGc4uMg2qAX8yN
dSN6cKu5iOlMUv3Dk59mkmjNGuifxvaMI866PqUy9bIitb7ls4ivkcs2jRzwiXkb
/yOXBuIr2vUstv3w1l/BD+LtQoj3qFRaNmGLDBGSOxpHNDF+AE9xdIkPyzAJUZ3u
vBNRAhvE/pobIBxxSmQ95fxkNbGgET3C6G/j2aaxa6TdbTA1j8w+4sQQzUjpE53Q
efgGuyiHxS9oKE6YnEO58kx9zG0ImOhUN8faSy2m/CU/gg2Dvn+isYosZiQeL38P
g3mI88BNcoFhKvx+uoEy5eNpxYQ1MCsiTegTLHHsnvep5Y9D539BtkFxPLI409Xd
HmkkoPnuWJk+Dn6oeGrqixk/BKpWyOHs2DHW3e5btQ3+3jJDqM9gadKARPrq+3Ts
1HU3bV7YYt/R7tApPTR/2Q5xRjowanMEMBMxESpDGYqv+HpBfZAvCmZDU9pWjFpL
H9AQdpbQbczm/MRzdBnp+rLc7WaSYBsxNdUN50ePWzPwkMdHi5VW4bBLslLhL2C/
jkFcXphfJZ3drJyYsMNOd9tP6uyboys2YAHku3mEQh5YDZsk9BEv5/kahrJABxTk
K+3xJRMSavfstnI0fCPT1fNbod0CAnj9DJAsf1AXpy/YtH34JKyQTwm2fC86PmcG
vVgZzMOCX/pVK5KJav3MHGh4p2abRPbgmGfHdf7iOSr+Vj3Cw0IWphJCPKEsNDNv
OtS5k/GPJvGeGvrPKuMJ7BMdRnRFuMmw+9YeYPMwNqQYShQOFRhsvjuyfjS1Gves
WmkxHKf6nh7RAd+ZZWRokDs+rv7tvX3EAfqbYaycBnQEQ9DLO9VKvuEXqikS0tXM
BEmEK53Ryjwg1T6xQl1o7M+0ZIi+FQYHhnvyoIfw4OEiL+uFnwaUtqF1TJ22nZJ3
NuAFhQwod46PGPYb1rKPlTvdcw3/OGKL8uoEm6WsDTReB9oQ/THRlF9iJgG2RKq5
pSStUlhJ6NAp124TYbCJss+o1xRM/OmKMjLOVkFKksM2wwanbjkIjxs/GKOkA5NK
DiWTxssp5KaIdPnSKg8nKTxrbJJiyENEWqyCTQvbDF0pSMEBWUyNJBEvaiIVLIHp
xq1CamqCVTnw6TJNx3nzCSCcmT0+6HPLcNwNCudvi8ZYUba5wYLA2zUHgnTmHSzi
qlOGfX2OK0sB1H34EOINPYHCXfm4J/SgPPmiCe29GwHcLg1jC06MqzYp8lGfdGND
wqPwVB36CJuKsaRZBqthKQL5UHP1XgTr1vFYqrkxmDezPGlyBLgMtuYZrooe+OlE
f/PxLeY5iCygJmI1CW6wLeeWevvhE0uU6gkQoQNrmDOybi1hogDb7KchcsRuw9Fa
UnsEGgTmbArQlOwNOGAygjfBnSVM0p8QrF7yFfiNs+x1CMgzo2i/O1dl9Sq0yHPc
hjKPz63uk4BSHQCmqMd8nAZ2AI935aYOHV0jntlubE2qV985MSc/sxUM8KWHnsqX
HuAXkQvZUTcj4h/KD/IzdCTKdMEBGSYTZlq/gNHdkXwxL7XgUiYEz8fHqX+phsw/
pluLNWG8vjAQuaN5R6usZk42RY32GWhYDrmWUAmA6iyGtiBfSCivn+hokxsycXR+
nb4WMcz3YIk/HZ/C+NqSa1sy0sWVpk0WYoUWlbeorwiN1Y4eNN6cOqCZLEaYMPw+
4jsiuYUSvvr8NpdS9/qZnWE3fI1wUHBn1HbViP2rYqgUUzehljgSXmDjcj6m9CeS
ZhFrvisCoi2srWhzqn4aDfjAKfc1QQTqBEiePbRS4JUxmzQTUvJ0YOrx53Gkjcdb
ePJACeLHK/a8o09nBb3pKzF4eOu2sqK028QzIaZlNyhHONTiOKdE6bgwrjjJhZpB
E2WDGtDDqrki49XsealvMouUee1abMDiLJtWFnyZwavnjlXfQkZCHrT4gEXomlMe
lepW/SD0ZalTTcWQKhbymgnVUQVyStkM8eQvrbmfi/jq2eq8G2DDQrZiA7b74zGn
D3WPTLNJbwAatCC6744hNN1FBxME44y7FYOThgWzz9Dt+utbGnjbZIN7mr8owMHT
gIv4F++Jcmlstn1ztuoLPGes5PxjVvSyRvcCpSCVvfGuqbtF3vmtYvqJa8HQu03c
KcCABXdy+oxIR9yrhTyMltXeoWkgvjrlRs9GaV2UykTrXmV1Ldo7UBw5o/YscNGW
vk1Hlg/x3IId4DrsR4q8lcp90jQcmjD/5L/2IwFIYFdVSLu0Uh47vxaB4fRIHXlT
6A8/yRR7WeMSd2YqHHdiqGAThX6LiMe0qf1JhIf4+awxNJ6xjQVlU/pBEgSm3lyf
8ycvBclVzeyVZ6cOh0nRK193mCCN58m+4qcjYhMRZT5FHs2xueg7NLjOPOaUK7eG
fh42L3wJL0Z7gc4U37Ewh4Jfhd+HebY/sQtepboAzrWhJo17hxfXGulR4GL0p6Tr
5z3Z2mtzAYYGST49P3rhGwmszpudR/TMUwagwlt0ld9GOzuHeWeJgy4zGFf0coaf
m699O43VhI9Cm51Acn1wQ3LyWcgAcwIwOR7bG5b2wGWirYqh03nm+VN2q1fS5q8+
OjaRce44cuRVp5fBWLTy6FiYlfsOrx4Quggg4uy2dn/u9QA88l+xZtfWfrFGYmkv
3SxqGcpLYJ0V610FyYFiIH74INaYq3/OoxImztPk4o7PQulUXRXOorLtmrBhWxzD
ptAFaZRTK/35SHPYJQKbC/pnu0dS1jqEqwfwmTPEYaT9cNUwEwQNNisg0ZH6Q81j
6gvL4ikPZh7inzYdQLQavyJhXpiH/abfqjLF7Dh1kfyaSRahMXr4HDGdY22iV8YG
t6d7PO0xsKTdlBse1tgbUmW1SmauDGwj6eP2pOQjKquvSVnj41JFdzH5FHKqBqe8
xNXgt0vQt0moIrp8n1vwgPZFgTL1iKQTWvvLGKZhca2ySDRDVLIs5wTpjSfNJXYy
MTpP5ZHrhY1rnbJxYpNZDNIPrnz2kyfkNWP4N0hBiTIRBp/SOVL7Zx9S5R4W4Grd
JwjypZHEkU25Q2EmZRI0Qt324bLN/Vlta1hKbVMCqBn18tBxEJ5yRbQsOMv7sxqE
yfV9AW2Iwsy6uzUVVuqqmiZ7sdwPARFAHKvrSY4Lif4/iMqBMMB7f95m7cZqFb5C
hsC/PzXuhq/AOGeTqWMtR7LBsgx4ZT4jGChL4R+I/muZykdDwWn9nk4a8sy0RbtY
ObO4HAOhdobzbVMjNOM2Qz//OHS7CC1vH2WcnQiYZa4ZPhSIWghPyOrdrj+tjjoC
q0ptRpChlI/+SRa9gJEsTrdqYur0Qr98s/TjR9fh4QVsfyrZPPG12DGgdLg7ZwMr
1YQv1HcToHKbmhIhKGMdSpF+JH+3KY8XvtrDHRrWYgPhmwi2ZeZlz86xyJrX5ons
HZVG9DsTKrEOGFdvKD/2/48rcl5kfLmnxRL2eirVQZXltzXFEOfWFBmQoKSbKgw0
tTD9IAGq3xpAgNnvunBwCFzKo+/kr7OJdcX+ryDEUSm5Ib/6t3ZQVftVH8JbcFBK
jc6rWDVmq2Ga091JoOfoegWcCWBrlk664ymGIxpbPHNOuenJj6o3+ifgrqP6Nv0Y
Kr9bl8ERdzg593j8OKiSzu0/XKjMJOBNSiCGVTldpmBHSaKTkkJMHPVSSqteHQhP
9oWBk5g2zEUM0PDt+N5iiXl6WqFiqGTnjJ7bCkVSkR0qizP65FBVx6QMc9wu8kEQ
X/L04FwjvN6f2H7k6NamHpRXfp12Wmflrz4Cn2Gx0ES7wGH4Ycop0U5Spjpd1fIv
4nqpUNOwZwuZerORiUVpIhfsSlWr3tz3DB3ntUh92qPWm4mGZUPLDkkPvxMwj235
pucvLtPhD8N1zFd5Vwh06Zu5WVB2mDWPX/Da75irkb3001qVK/YubEmSMVamiABy
nvB/0cNz4+bG++H5jhjS+laupME0eEg0o6/pWFZASs1QD5diIkKYs3R+v0jji75e
+QDOi5JvCwt2G+i6z+f/XEBlxRxE/lcQcLbHOi1YSaH2RIc4VD6sqRwMjT2lw9Mr
COe506LE//4NK/P8tDVdgDfksLCuSqEyENtzoMMna06f9dU64nqRBR9sNhnpPohw
7oJ5xguOHJdyw30xjT/xTgVsT9+6j7MxP72cQYHfEy+gzRqCyj6qUN9B/TAVI3V3
90N1ibTD5hAjApHVntuo13vlGmKLUT6AqT6+r7AdYV+DqLyhgpxrf6cHhs5y0S8Q
c5Spd2rVzDG6jNrR227zO2mUM7jpd0s6YJygbNOQYmUUb3sdLFWw9V9EuwBJffe6
kefe2k8q9+OldTeXzK8hI8Wpv8p+DV/llixGxsYe8ElgVrCKtXJRKZFO0mb0JwPX
l+ySHKVhYGeLBwaotanT2qo4218K4CeVHSg2rtPA1DIYfeRwgepuSiQGvPyq3LvZ
mv1VMserbriwhvYBTB7ab4f2N/6KrktsO2aaLBQyxY4duWxfiBnctMAOOc78IviW
9Ef0oozvxfqWzRsxBvusYbqugf05DvfhnopQ0MO+ibV4srktuH5CRyOlTFcuc1wq
+DIh/7f7kn0IU28KpzOiOyP7zffUEqrKuWY8udRYE0zYVC4LKRTNsvgi7zJe50Px
slvbUvu9igwfnRiJxqEpP/jRSbkXI6vIQdPSwapSZSduzS1HG4xJy6btbO56e/SD
7G9IhvEc/dRjLNQRComLwF0BCZhCZxFr+oz8O64/NiZeZOk0K4ZfdsZeBSzyvyEB
ir73h92acb32DZzr0IUJjuAEnumEL8nNGAC+ktOJJ3FdAwxr4YOYtii7ItCqYsoj
cQFV7GOq1nKtXUpPADuBffMP330as6dQIzwLp2aa5OTiMLKhE9Sy7/CQumNk6rtq
Ls2ZO8jPUVxv6hmBb71tgAv7PPa1t3+WWPsGeaS8076p/1uaSo8MQVsb/eMUAoSs
+73oSwjMI3saQb3w0Ao2Gud6V2yahlO58W2AU1LV0cBVCq0zi3Yv/LnaCzhjqkO1
qwnJF6c4rtWp7yiWlK25X0dIfFnh/YD9Z/SnHUUA/kdQIG25c6QwPwxCSwYjmuoj
0GxhnmSH+d4zE/VFTdpFCgKOyNaYR1e9mCTEU7rhh9bISnVRksJ47xJZBvSkFBsP
BDuD6D4uTLwEkWSiqhMa+2juax0KHR+6UDUdcYe4f85U0x/lZuz16X2JGyi/kl/U
VM6+kGYxYC3vOcLessANyf/b8ndwWF3iEhDLgbkUsmUa0ecHp7EVTDy+i2YRUWvT
gHwHPEPKZ/3co++S/5m9fJE3lCElPVGtVOgORZr5upBn9NOOoGSP3NCRidicqOzF
nnnqIbI8VmT0GQnB1ad+hIZZ2K3DHrVthjBQmXCcfo7+E3zeeGntycZzGGe5YofQ
T8qhnM8IHMqVPnpdlVJyqlAiq5iF2QiB4z9L7zcPyOFh2Qj1gdSgemPUfnHxZqV0
9OZkhEHh06tQ8OoLsy8y5rubjNSskQ/A7bI8zYKiKOE8E78ps1tA/61lyc5WmwLn
30N0hr4tMxz4URN8SwOpqpIL2zSBFrZRH3LTJWNzVON6+oHAERirYTfbOw3svGDF
1jswZqv1vEDkCFP+sGARGpRA0G3gJG7nl3S9WwV7QztfqxLJxMn8sqk06oUsPmiK
adND45xMC6eZ+nor+q864efvkrgWv+mZqK8acTHPDywj16jklpGMk4KfAEX1AsSN
drR6nDsE+iq4l2HGVjyD13qOx3QhByUPc/f9EAHr5P7g5Ea/se7uXVEBI5NZZn5W
J8Sw6JhCwYxUDdrsQy/PMee1zcjfw1IdGeSOXS5Vr48WBQ1l11XD1Qo1tRONH7Su
Gbes8SSTWNCUt6At+0ofW7ImO3xfaLKjrQXfhgOij9dApU3wRV7sL9nDiZZc9Lg6
4d8+fkNYozmWyFa97Dg3aiL0tc/LPGfDEJIuiCcVx+nbDwa+YuejzRlkuJdYEbEv
cC1a7jTZiJHz2R72DD7+zmeOXK9I0Iyatk396OniSNl8PA08ScWFQRIWKaI9QLrR
w+DyRkqvIw1hyIfdP4MPwnnPPvNlPaw0Ir5ACEc22jtIwBKDH2puDDxbZ5NGnr0g
8ZN2ssBjyFbZXxrmUynDO1vEMTeLb96rfXUdyREHWUTQEt4VV5vsjBFfQYBT1ZCW
nwbaNf1+QwItvE3pisOq0UsUERObuYyu0oUbY3ZBNih2uRXwi8qqNq8x+E+xVNV/
lAiOvtiZ6gJSO9G6Zd8Ytn4pfiV2vZPuvOxPjj1NbCZrZBso0wTlEsdVeWp2ow4F
QzIRHc+5JWG/hLE08MTipYz55Bl+VdTjM1FAEgeaEveChok395CIp4nAJKzPDvK2
ThP3Yy2vL3hzeFnzewUfZxI8WB1BRa2wtoHYEdzX3Q2Dq/Dm0Ysimh7bR9j1+4HW
JOBHaiFXQw0ibVXY7WZDfdbGUaOMOuGUWlV7vKndSSfeK1owmHf0TQYLC2MZWXUC
KiRpnoEXhsTt5VWIvS5NlY91sQF4gRFqMQ4/qboKRlq4m3ytFYEnJ7hFBqAUHOAJ
C2ilRiDXhTWGZECdRE23j8C6MhG2Z2iJaqVY3EKX3ox9UQS8Yc+kTkJav9nzJbVc
JKHMjqwUuwdZpHqSTv2Ehqg00noq+svcgIhKw9+ewOpMODD4/n+BVvkW2aBe8tFQ
9AW4PjxRhVaM9w9uE+lmQXLnF7DQyAJ/BSzE7su86xeaiGGWEB/bfi/SrUNNL3KA
tNOWlBVzaAndYpIONcLIl08W6ozMTyEvOjWs5vM40BZMLqKax01wV9Bn1tnLKzQL
gR6Ikc1WbWmQvJFdGBJbOCvRzBQ11hnKync3FKNH6XdGbSTsKod++sy8r0OM+o1+
MizgPpk991WEZINkBiJaArQ2A8skaUc0pUnNoDpp/V2i/BOXEqj5rx464d9l8ahW
vugplFu26GxDhxsx5dYa08Q9g3w7vTsoiy5rCdbNwDJJW5qk+K0Hbw2svx+SJvLq
V/n4C2ChpuLNXNWugnCmcjMhWCrzdTyY53w9/5agll52r6WOru1Rc3QGJa2JNajU
iKGIwiVqzCDujp4Uqw336HmgaRRCp+lKcJ/Ln5qiY8Y+MTVJApXkJDEBKGJQAvYa
BX1p1vDi7weQ8YgmMX2bMdjYPGk+igLOp0TbKErGh74YtO4JudpGTxPX4tdcdgMl
MQoZYDqqOSDJBGkJZiCr4+tYNQIOobgcpVY6Fmz5b6aiv9Cyst67xoZaQDAtviv9
CpuDp9Jkfx8nLgj7wuZ53+vzCdrUZjAX5db5Bx8XdYBmEd9q2ZLyK8jB5QeH34hH
o6EWCGbLru7vsG8fHV4DrBcGsQEJaWBoP2We/rbZm8xGkw8Bl2284t9z2DbmbYKc
dDzLyQriK02xD/kVLXKhD3K+wEtp+GHpmaFxv+uP159ok9qpMUw+WWNsuPNoH96+
IUeZcSUwddXfG05qpnHTyA3Fcg02nAs3nZtWW4GWZkK4PPjKPIo3QUZt2CfNVofh
vwB01sRgiFVyeLIZI/GYDQf4fIApDe2lP7dSyczHXmRfin8UooiuAtc4cft9tmTE
CC3hVRWfllkWxQtJTYkFXb87tVJXGEIcz5PI3AFPPl+Gi+D+raYPhWkvlXZN4nlA
o1A+f6pUI2I8WLZ4LqdE0BrPpuEX0+557rqv6fYLfxzCfaIjnelzj1ZpPjFF1NDX
fostsaY2Y0xS3bhxGrc7ATrmnP3YhrL+gU3EO82Qo05OeMycOq49gpJthKCjJnBt
EEqsmp9VillQb5CCAMzzajlF3/SABejjTIJjQJapr7RnpJkS/J7skiGZ7D5LjPxg
8Kdyw5IzRDUMTKEi/gtVLaD2qHrNR8HbiCewxsjE5uWqRc7SEXusoDlB6NlpvEjr
/sdZGcxBZIYtstWkV2TAyojUfS3hY10HR6eUTz4Muccsm0EA9lqpHnFOQPlmaoif
BumhqKk/+EXzEe6fQKhD8UjoINf/FmvIDZwDsCyjY9gh69ADxtPpAjXjHfbM5nHS
2OlS+gCXQbxWci2XITKBqp/dEbV1TBuS+EAA1yvwq1U3ZV5qqQ0SqYvND3dZajv/
HkXqOoY0QmcQ1V3njjGy0cNydIcE3iX1UGVv1INeb/TNgxr0bQxCie9h6MaHJLcI
Z5yTQMrnNhBMIJRFkyBeUI9YpzCaPZ099gchklxChIHWoaXcCzMOuSZLBEhkCpCI
xaw2/yN7+Zq6tyfeZhsH+dXDijXgbj/gKVmOWRwVtaa2Uxpgvgt8CHvX6sZG6MPj
A7x2DE5wBoTykADqtNrwXt81oiIDHYJumh+PZUbxh2h/VaEYxhMb1aMexZncFQL1
k1lx8haCe6/tUnJlZL45XDJghnIwF8/h0tn/r7hRjQgtf1unm5CZgfVRyC+br5aP
EY/Ly/fDAlikB5mpkQN25I4XWf194CSGOkxqsBzYxWlnaEr4gaJ6Y2IYwqGrHW1T
AV71b8dRpjupQIstFubUF7lUYnmmf6kPaQQum0PbFuPBa88iFKN9+py6AOQuJLim
BM2f58ZrRxHa2IDSTnntE+IYJbNjgsYKf5lx6HKMUY64cV7mxC98re+Rho1RubaG
HKxmrCP5LhQmAkpAp8jwZu0Bt01T2dHn4DnS2B0WuetA+4FfeVgJW8HB1Rwvt/lj
swbTqLAj2Hj02HMTssmxrZgoFCKtt/BnYTnJj1ojkH15xdlHAV0dlgVfzMHKaDMd
sJxbSA7jFaXGbDR8tQ/oXgKIUVQot33BqEWs9gk7zY/xVAmbdnWk1F4Fn8bVx2Qs
vUucN1u958jrjZ69KobSD+1D3Xv6M56fURYg1+HKMhFliodERiXuqbF0cE5Wz+ab
jn0vClkryHKcEKTk/r2nmIZCYquzsLdgfU8Xd8o2ZjdO7+pG1zHg/qB6+ccCgCdD
1uHPRSNRQwXUpttTcwNxyRU3Llp52zCqitqzCX7aFoj/p74qR1iwjkSwH/bnKTWk
fHkDQLXwXH5FZhi2xJRcIY9WlRoniEdyTDwIg3wPgqDh8uGNUq4gzpDUWUa2vMYh
pZ0Fo4Imgon9LhHOyC4gEm20qp4rXjixVWXLPZVj8bhawZTGALpsC/AQdGSg3xSh
SRvTPn9EANPqeH+LMY+ui9oUfWmdCSAmF1Ygk6JlWL9ajel1OCu3cVcTe1XmEV1A
im9DIcKeNSlsDhmU34ntKjtD2u3iRtju1jJgGU5ASFmbsqVbuLzwm4RBBB+aOiz4
u9JaP1E2f1sleITLUrV8xctwFrK7V0eE1P/lpjbVNkDOLeVpMHIr2CtPEk7UIaZN
ZBgUKkNSnwrOszAimiz2UMIlge0FUd+ontAEHx1p9JgKJ/+1ftuZ3p9bI0wK/dhq
xEiymen9BLi/vnqWUALyWoKWaTUj85qQBoiYfCJ3rlJDnShMK5LSqvpQGAN+EYEY
kXlN+WhqBPXk83puc/4Y3DWsaM/XMJ0XGPuTfHbCf226UF9EFp4Rw+Qw/SNFaela
zYzoT8AlMNOiBXWeJYDxVcCurTU4mtnMdw4ZXvS+frvYWsTqmEKUcjd6rtnLZVRX
iXrOqI/CH8fexFPq1rnCuPnqReTJjrs+cNQ2edOZ7qDSQIw2OW+jf7E09vJlADeh
NGY/YjzKD+2H017EVDMRYvu8TvZOkAMLdZRSXJDx3tbDIQxeeMNxYn7UsG5QIN9e
WU3YQbUk18SQ1GmsiG3FeZupfer7gPTyErhY/+5S4p+Egs0nPoftYHX+kQT9/KQa
7SvP1fs6I8jH0xnVsyb7BmbzpHh7or3STOflc0qWefmYNTzgpAFIbjA6HjTdmJOf
j+yDHAWXe1x3Jaby3f0PCmZK5AEueL0YWcK93D/6CkYuYHexOLAp98rZrOCZsgh9
LwLwOaJ/H4/uLhyvxtd1ETCw5rQPIAeZQ/GloHaB5EP/I5T+91q2lI8ft8mkeofR
Mw7f5fWxPU4nO3zMHvKS7W5TqkWxwasJWtJBLEweCrvqsxHUM5pys1RzumyroCvc
IIACYAutbzy46tXOMewFIvgKYk6rWWwO0qRD7R7fzVJyaNzFRRXSW9fL7AjJU+S8
z7laIRgnOeNhI2Vdc1yKdQaNoNrplsLob135A+zM4WRLn1ocCsLe0gESvccpYNw6
jezAhyD6I+OdafQlX7VFU3l2oiDzwrsh+YWL7VH1RFYNhdfm3obKelisfdg1MDm2
0iTg3lYmjUYbch99H3TvfdiHKXsPX2AATYjkwMGYWID2bAGsGCX8WENHI6dECQ8R
t5K8iu3wKajBgefLR+c5F8dq/21EP1a0YLywU2dUcGLe8ElaHMGHdS7u8mMt5+Qm
v4OTyv15GhMru6GgRzTJ6R2htTJsOJKgftq+5YN4tXmLK42FR1MIDeRR31vNxTqb
upcnjUJ1RtU7aNclNuoBbPcr9Khq0oHt4QlaLpeVOIAW4ehFGNurADj0e7vdZLrY
pwzndpma1rYFiwdHRBV6W5qj9fR9X3y14Sc9slYCta1tbZlTf7f72VHLOZjxhijZ
CemFXuXePTtQbBDERm54MaHLl1SKIlcO3qVOQ7bX26l6BD4srLR1VXs9bCxVIWjV
YKOPeMuaZ5LKNo5BzQwvUR+HhMVtaISu7QK3cdrCpYJKuOjWxHiyHDKxJ3nh073K
PSCtV+lSfWeCcCXhRMCYNqFEmWTrD2eKjJSi7MmfQ07/HOrGO4ww5JrWcC2yisAu
6hsrW1NDHJFMoKRdssLTjNuCGbKCovxGH3GnklfEKeCzjkQKSa0p+c2S2bkVrfi2
v6So4GldtztAHeNrG649oFgAtWQOnO8swoEtV/LS+7ygZeYFf8dTU+//7JzaX1kT
gowg1cURp83lHsZsq6trqLng5DYpVI5ylYjULcKJMrYjhX497YTK77Y+1hPAxMtC
bcOnCfNz9utfjAcHYrqPAk7cl1W8U/utHzoy9DFe719DI7h91/l1rmaOhigkV3NT
SYZLW1KHoi7xOPPCk7+to2bqBiQxnybszkhOSI54tclYGqxkOGjTN8xVDOJ+ArjI
7Nv3ul0BFM1VmpJHbWBxuIGMc3iD8vTAMiVdo0+0iTg3nBua0XKFJf//0qSPaCoo
NehHFNVbXegmdCF6YDHbZfEuqwGjnfTYUgiXK/Kci8Tsygfypx4FbZAgBpffSOmf
BbVOOfV8XKk1oItvFf2JiMKwqvcBd5Ewu6wLMf02WksA0zhX9xPROXuDsJCKbEyy
K1IqhxW1GSjl2GUA/UBUEay6rhCJ9l2Ff1jtUiQpaNx/QSZOCvo2I2o5ec+PvXEC
tQNxCF/HIc5rwsg+Eup+Yi56mj62pp2t1zsj9QFHq56n5kowCXZRywNL9EONPj6s
jtJaOwMUvrtXntthBmrGYtITSNFDDAbxTrDjg9pJSHAPeIp7nERBEPSh8Ik7YjVt
3QfMbIR60s3kgw69y6tUWUNE+gfC0TZkfXLIDDmyf53Jq1BYM6K4MtWASzUywyVp
J4ylKM/yuT8qd1eS0sZmrvA9u3NlwWeFgUtF9ofUDJTxpphEmawKa0qbbbH2/uIl
Hphau/bmmd8f5gej+Vje52t4vbTdUwBKRoXNu/MB0p/F1ZaL+kJ8yCERWq5TS1/v
ZHnnqPS0jIp/Kd9yovYRHSWtT1d9JryJD+oF+/EirCfNf1Gy0tUKUeVcBvPUyrXF
N9qP8AZ5B+fwWTa0G0qYhZ8kkn+oRWnTzpGTklqzy0F7fDTrP37eUwxRV19kb7Fw
8kgdyhXmhEtWbbiZDBv2yHWeVwN4dcET13i+ld6nyipP8LS3bfx11sPmraTVgoTq
w40eQkW1X5gDsFV0qq7bEN3uWiVC5Vk1Z8RMz+mqBTk7TvNQbGn3J+LmM0kfopEc
ASA3l28YExa2PATe65dkVZVMJwls/K7rgq8xMWL77rFe3dYdNotOTR3fFJQBpP8k
wJRIcMBg0hJCNkiIM7Z7xP2n4CekQl6y44pSNd0gyPcxM8G0i/IuhYhI9SvN7o9I
jjBakqX+4uvx8dCxNWPCZxFkk215CTBhRadJCvAmpKxY/flY0IQHdbFsmHKVJDul
OZDZ/P5eAM0zoqQxcRNgXJQic1CfvXbHN35qffRArMR1DLHVJH7HC8eD+se3JYh9
EQkhYm6cxqvOdxrpCmdJangaFAgELx4m1D45qUwMfbk4D6woTBsiOV6nlPKUiJ4S
lnYdFhw2y+yD4IlTMLqj5Uo1psL28a0TlmSRcLNOQapb1HqBTvg7DOxgS7Iy4xVL
ihXfYpsg+coNEKQHVxXUhwB2lVSPB+sVQG5fDu58LCEMsxMv9OUpf5PnayPB7ibV
JMXHY8g4I0+Ll1uDOfJDvvHaSiSPPNCXzCT7QcJd0a0Jy75Scq2Sc8aAkIEjcSMa
OfK6nKl3aDKAWKGo79rffiDDGrIzpEW+L4TNrJx2gaoSoKZ4EEkePl1emihdDdl1
eqOL6jrQlVCwma1q6LsSKDof0fjPHmHL/AIfLd1OToGvoGSKVghe1kWoy3TYrytE
dKdD6bdn04Vz/S+fY5ksM8l82bY0bgbN2IgCcCpA2RoI4GMMpFcQwIjctwpZxnLL
41RvMAQdIHYnEhv/+8VQVSiG9/pq/qOgPZ3dzynWbnsDNE9ZgYx2ihTMIpBhzPK5
24V+apaK6RkVnY269k/4B2eHBis9C8SUTDpFDnY3kRVQuyjB0/MDYykcdeUDLqKU
UYb6lvSyUpUtxzY5uX1gV5gRcQlYRpXYUo0toovcx+VwzzMYq1fgBRComoRDNCB6
AWYJEyYG87vXmduiHcbCKx/vbdEmSCX8L1pXK+Hes41eNNXvcUDmwCkGq/z5u6i1
61LD/qCVjocmW36X8Pzu4v7jYetJ2pqjPLQjUHXKFtGgPBgPgVeYxMVkcvFsUlko
gBgp9RsmcVEOJ26xDi2BU1R4qT8w4mx3YRXx/vHXfORueMsPJIRwrOXtCWRENpdg
KiKJneHM2tnh3JL5bNFe44SolAFj7y/+B/0VaFlL+y6KnaZraPZijZ4Uz8gES7In
C4tHQYcW8pBjTVe6DXPEM/pNkqgXaeyqykJoIxKDQLYYFz8FwLHoOh05J31uEe5k
T6Odw9uWB1NxNth46vb/c0G1QcHA+0hjfURjmL9729i4t1R+F0aeaOq8124v1us8
tFUVOv1JOFv6MQ+5Qj7l85GRbgbxUUY7RDEneLk8HpE6NGxq8vN47bEGl4FKwp/O
sBbw9gJPfLRDqU+UfQHFGvsbw+2tsqtcVlfAplrQbgibKVLxgWnJUy8iUNEIYyPj
u5eqgDyfyJRXIoE4WP7EErKxnHFRFUy8mNK1s9tGE/FjAmetxArhcDBWlD4XgoDJ
UGFsi69A6bhEifOBDrxF/wkrM3zbVqjqZ3UyO1LQz9KIfkK0DhN48FdcA6H4Tf1y
0Jxs2aLhnMduv/d/VNzoCqXs6u7a61KvDjCwPbCxzNSShTfGRfB2kkJvPAogfgpD
EVOywqTK4Uuvm1A8+bQTnSjIz03wIgmmL16ajrS96Y6HQWwsCrcydUdPEFrLDxIb
2/AIB9O4RMbL6rK67cz8d2mx0Bbx3aQRv4ISkBh4aGWdNF0mYuf0GhGZJ7ouK+SX
AnvrU/NNSs2NKyCQnD6UAlVooE9vYfdiZDLTDBFVEEUrLcHtYNTM3qAMvdtHGePr
s6GVkq9rmTq7yDTuGELF+gvz6fjNq9WLL/EvLC8ubStD0xhFuX+hs+xIqU888bls
bvSu0p86wuodZ6F+RoZ8QiTJHF3MbAx/41bvoWjPEz5tI9Wc8VinBXzi5a63UG/x
xEc53VeQlp91iMpK90m4UZo5JpHI+kdaF5e2yn48rWTvUJ+uvV9V+y9zV7z5+mwE
/Alg7uUljCuadyBOST1Ix1RKJvfEWCKRb5/cZjqIiwg4fkeKzhnjtzo9F70pPwdk
3qjpwlXQl78XmA1mXXkCJaJsCudKfgQD5H7VSgofDQqwrAEfHQ3P/Ng9TLrwjJz3
JX4pi6rmWPSxY3KAg4jdY46zjBH9PUserlPZ9K+WYwDgM/VPaSpmvwxeFW97rm+v
f5Qj7qfFBzzDMkkReaK34CV9i7aQpBQWedlmTKMPcy7BueWufTK6eV/HXfHsRGhc
wi4pdLmHex+vKJuEbozwXWJvSrQlYmwth/weICf1nuXXZZhjI/SVu2qcOlDPsVTq
Utuptmd+c1wSqo3TwLEpELt7lc2D/FaHhseLtMJk1bwUNkT86zd0UxZK9AeBQ+cf
3CCsEeTYcRO7umU2qdFfNXbe+nt2gwNNH8ItKilI8T4GDBB3GE03LF5/S+TBiSgx
Xz3Rt0ixl8q4JjXanFHZgfEVHih45iHcu0UzPBlAC4ofVkY8EDhJM9m41Kz9eGHA
F4ZSsIA0kF/RM3bQRR+nDC523vG1xS7zuhrN6w/fJUb0syHu6kHoGcABPh4HSfA+
ynHS/+jhgqATFgaK3zJtAdCJSWLnIQHZrP/jIsV2Xm1WfNeHF96nO0gku3w2//PJ
DvutGwUEzvRupR+scegOmZXn7G5SkqXWfSQbcSkEUidSOS3QvBjP/K79eXBikO62
dGTxQMYIq9dIoG8jPa2ORt0PwJkjCZYihpdcatZpdloXhevX0q9M6NA4qj4tnOdq
bywxK6ijwdIFs5CTDzxxI2os+IOFifjNiXqd7S5Y3AzhXutigEsKbiwQhigROs6S
zrwOEbsbh4m2hP9EFc7hevasTf/IbEFXpf+Ag8G5j0kT9/iuMfm5EJNkXyUJnGz9
72CLkPX5OUgNyOf9KJxG8gmU8szQ09uW/smcwuJCekDfMM4U1HIKJm9RDb/NV6Yp
rEAer3IoJbMi7gAYfVCn2k6OrzdN1hsk6wiNcArsQtcaZXPOKAmgGW3aGELed3Ef
5dcZMzkBsxVIV39NE20Aa42Erh32+JbRfULNVg5bVA3LBF/Dhc3Vum8sducJJNEm
TGr+zmIV3XL0eWffy/mMj88besdfeBJ6vzSr5HB8qUzB9xi8sWq784tx0LQSdq67
Fa3itEsdKdvxsW/koux6jNvbc91RUHZaubFUH9HozSHiTIyqRLQgnzu5ByLfR97O
TCMrXbeKn8Y6X75TsmPh5u19FipKdkVmR10vW44zGwUEmDgL7m6g69wYlClqG0/U
Jlv9p5YSrCUSCI/QULcrsRz1JOM89/F51jHKtWo+wXv3NG5vXhE4O4EVPrsedW1F
HdNFT9mu0BS4Bnv9Z01z1if58p2UvNpR6/8QnyhF3LhpCNJox37OPaw5Sacon2hZ
cnMsYrRmukScbof6VRjruw7ESNd+7BM5iBMLkL4UszXcSQpsk2z/GlSN49fq4fU6
8VOlfpyW14qsLbAZThOZChJqFu9wvMARg/v1KEBBvmUlyr+gNfwB/+m6TgvtREFt
3XX3QHtgnioRIZP+LLqK9KqgSev2sjfvttoi1Ra6UxiZyzTRgNHcsNhCzse0vPvw
ri3jpVqCehNGzALbF8jvxFu6T5th3qMFm019+7kL8CEOFG+pFWMeq/V0GJzNmiH3
JSZrxlVa4925CAtMH6ef3uR+YYp04ors9+J36sVEqQ7D0qz69wbpuRHoYzULhh7T
+0jp66ZBjN7QTC6n6vGoPcET9RETGLKu+3ramJDsxKFMl6HasihxqC/ABDZT1Ajp
Cj4H9sD3RYq7o+gbdHaUVVa0RRM/pmWAI9ZZuG1paGUzsYj8arJ8GcHyyxi81H/4
dya1ABjuwIupS6Hn6lrzUIxMbROVmRatOly7zqA6AQ387PNNIEnUQRBN01BRe95Y
4I89vPTphi9C44xfw6sqrKI7c9kkRtJQ3WS52OPq9R5AoJi3gWrASIwpbblQ2bpY
6EcCHQepB6DdRzKF9LrUSty4IiMy2mD4mowE5SDfv4DqqeCcQTlCc+kbv6ZVPO0f
1fvp2Ob1RmHTAhNJ+aA07RoPKqa2UVagaAXqPCiTfmY7sHqNKAEOlhxRCs++pY0b
HntNGGgE+KJDuqb08+V3mKwUdr0W2skmiHqA7PJop6Z8fzJLdVOi4oHDMwohn51P
/+lVBJfCQdcoIGmml2nn/H7cto+kZWTqCZt5kJ9uK0OXU3QdCGw5nOmYGO06In2w
pkBM+4YsE5LPo+D5mdDv9Lo5uqdJ53obqzL+krKa5SkEjN4fCmuP42LJ3WmhV3wb
TPFErv//dDIFx3oEoKv1f+G/bjY2wmoTyFudrTvYAr+gewSUm0JjTU5G/K+320j2
Nfdcf4rKE8l4MXUMtiHygbbNsen/ky/YkZgaiz5kWTNRLjKWt2JAnSidiu2s4Lkt
KITq4JdZ+msSYoxOksFoaAgT3E0ST7UzByZAgwtQ1b4gZGbvnDEUzizwWB6a+2ak
wOLqH2vxZFuOv7Wz1yr40kAh2NH/anaBbnhPEupt6BZTA9nNv5wo+6knihg1Q6QX
nheFmL0b5iIMautOKjekgOWDyicM3+tVaLPPRIGTVicmUn6vGi4ilo6gWpB3Cfty
EjrnZWhLDnePrJjTGE4nljc8CdAma3B30ahsza7sKrmOWvRdyRSchieJPzx08+Zg
5Gmts+BRKsmGsHh95nkVZSkg1Qs6D9jOn2mPVrJZmo7Gfp3jCj8CH3bm6cWgtzyK
cB1lrScbqBbH2/K4Hh4deR7iWUbB7lw9K5oYFPIRkUAuSplZaIiQBrQoiFs/UxKU
JDXC16XvaQ8SsAazapetgx1aw3Lbz6ZE+eNDihg9NrCvTpDWDQC9SyDUKjbnRrJf
lskFOE0ADl+HSyfahWQTWBkAP583IeVJpYvZZpRp9DmmbBUUTdwd/hENN1Zky1Yt
3kJQ3tXGf9f3KM3MGXuKmD1q4f5NvIvjw4mVpqUwj/2J+D5btDcBx9mzHGalmxUh
nHG/Bq++GhAJbC48KKbm7sFPZDEwjsm/H4JdYp0aWy7Ax8R3GYHODg9+VfoOi/as
eEivbPsLkFB/ev17t25x6rUdRG5kKd0etH+MnwJtHaGmCCllR1367P+rf/UlQtqR
XrIRbqcIH/xHxpaCjW8lufrve/1OVKOXGnsvjLc3QVnzfXpJXfwWGypkSkY6dfvE
WCOjTuTi/D6NPeWhS6HRJptwrZtHQbEBipAytRGMPFhn5GKgMb4QZvM+57+ITGJ5
hjDJ+JhH6dbRn22BqHIZFEI6+YXlvVPy/BjkZDmklg8VA+aQ71/vDzJNqoZsYP5x
CBKhJczoKJlauLGIs3H4CKY0enT0jH32+yUfy6W69KdaaEMI+5QanLSY8auInZ0A
Cc0Yh5AxtPPaVYjtsnPkUqG4PH0umpPa+Y9hoXgi0y7wIRxHIzLUw1UgzNPr4Jfb
Z3Ajb/WPmXFEYbwCEgTTYlG85rOFt7vBhe43ECV7pByU519M7kxEmvbmT0sVHzph
kcB/427qiyNlLIzYneGZU6QLeFNCxsij/N7X+Yk1rJ1vOg7b7k1Q7Z8uxTXRobAb
3V9yoseyidiu764Ge9IsLkV1cls6yPOPkHvAiluO1KfRGKP1y+/22/XTsQHrkp1P
JfPvZCHQlMGXLoxpFL3wJcIZDrL4gaYwEauGptClJPysKF24c5GnlXWPQ07YI+0x
+b/oJXLoj2c93x6cTaccSAalBsjZkHlymkPB6KWZ2FqtNAoOOF8rPgj0MP6Z959u
a2aycF5vE3tl0Vv5tU5AqjeaeoPxtg3W7vEe7ygzgb7OjspKrLdboYVDKOgSLfxp
N/DZMhanNOd72k7A4aF1L1aqJDh54aE4iN1j3JB/rGFNicLzTgHpFzmpJED48QAk
oiqpihGbIihzhSvKBeaRIRXloXkigELFBQnNxhWMc9mfz4wG40rc7R/Sl5gA3RG/
rzlSv21Pmhux/nDIsXXqfbIlVwzmdxWRgJ/51yhs8JdDjz3CfrlRucfPzJp5ntkg
E7qu2AraPYFVZBCDyXIVf/+ym+2qbKuvTeLUYN511PTXeswD3B8AUNgejdPHzOeC
8GuxPRUniJuIkYiJN2g0T3zEokqPl5fZwVg+UL/4QDHyBZ3l2bbUEGHrW8eD/ATs
m7G8Ck+cI/E61GyYraaSd32nSWOmsq7S3HA+dgD9IqFPXJe+6wALgJEbzaJNbcf/
/mFIAMN/xqa3QhSBCnXLaXA1FsPPp4zulX27wiMYWEvkk+xv1bpe+ZcRMF4sw9Jg
blUpaYTdY6vs7mRKEOpLC2oXZ7G/X+inNUw8MrT5Ow5P7rkf4J8QM7pg20KCmI6n
jncfeD6P3vLIcPXCsUtZR7J14XCqcwdwp46afGdLr2fvIef6vKFjOXkZZy/U/mAI
ef5IMPy+1FEXZHU6yna2IY2mKifXa1JHwmwdfOarkJF1HLA4FjK2n8XIHyJnKH2L
OXRHrBUDwN0UpkrKs6hTu51kH0lcckZLJGxJlgCAUAokYFfljLVcReNmqOCE9dmB
EB5NZtd5tWXqj/y70v3HMPRQWW00+FahjEX3XkkVKFxmncRMOseoP9vC2/NcQrLL
4FRoOsFtqL7tjjFh1HQUW4xEcajsXa9SkwLQlffh33JQv8bp5+954mdRjyGNVuWe
EozAmsPEHF9bgzFoNEQfT+U1HTeBq4SFTvfelCgedNs/5nYicao+eG+gsMyHY31k
3ofZCjwa1meXRmbnPYmpm0ubirL792MLtssf2StHE/N9pAHcjk8l2CtKDx6fbBc2
spa0zspTRRiOLw4Qhdp5HX5tF1OwCHg7+1tvAeE0NGUWc8cQitneyrUNqjDoaafr
lfY0fVea/lbUZhvlVF/8n1nnbHfC/BB0Sh9IVzyIT7EjK39k1nvz1HIj7LMon5Gv
AamrP7e+QOCsHX/4X0mnfhpXF+UMLZKA06XE855VYetahnVKDJ6Gi27OcysJM+z1
0Fi9T+o/Im+oIS8FisK/ZUyEMVmLxJIpD/k9Mai+Dx7VNiazcwsk4MeqCUjwFGFB
jm0F8ol/f2PX6qRZ0/4/EQ43eYg6tuBGCwnT/u2V4kZbFEUxbUz7sZo+i9KkIa5Y
OyETMdLxRxORxxbLvOQsMOZdaZ7NDuKlqxwJuhZ9mlnrZ08UXtjZ/HUx7Wz3ZF8F
cq3sB0IN6nu5+fnwJD48ZW7cTfio5SO5P0dlT7ZjD06yb8wtaJt1PamHMTAyEBZ0
EpVPaHtDeJLcSFwCh3+N/nz4onab8F7bPx3+LkpJ5rMkuNvfJvXs8HD+t5tgg/5z
kNFGUIurCqk4F6oYM9iJClZtr/3eBIMY3DE8L5UQsIVO70j7FCtuimhsuDpsHsg1
DQ9Xk2RD5wGVW7OSHS/FTC9+SV/XQVGLrOMhcJ8x0bOgB0xcdO//idxlF12u0XoI
El4F3tssYng2R259HdkC1GvjU0GjSDl09achmVQxWsSK0XVUzHw2K1aAAxUcp6D0
0oX+MepVsdJauTEca7mchjqvx6ub1NBVrgYee4ghnko49JQmcpBDPL925ig+fQYe
uRoiJPgnW4I2ypQcyCqKTgLO8U2rbXVVvrvMIT2eTfTtHZ6XlG+TLfCnFZXl8OSC
+2valIRcNMtNilkKp2DSqYf2EVWb2OaxrCwt5kwzGri14lYKn05tDX9pgwSqxHSb
Rv/FEa9ZuNhUewTY4S36SSsxsO9FBWorJui1r81/nPEbPBr1KGi50JeEBG1QNg/5
zLcxfZQx73dkBTaTxWLhZdQM5oMJB/07B4DVy6iC9rkTkwDUHJ+u3iS3MWmAl1Yk
lkq4wpH/mf/isPkkK7Ep8n9Sr045NVi12UXeg1tlh4CvJxOb7CH44rIPILVvQndv
ytpV1LVeuTgQLcm5CkD1n0I8xm7jJvZq5ncb5nykcdmBdRTcAtwQ8ZwiM+LbyrRf
wqDWNlQYKD7hZlhRUo3DIl2wdfSdNMb7ulddiRCsV3qWIJZct6xvOYZm/QPtxcp0
x25Sxboeyxsyx9gXM+K+hrv9Rz+EsWEcA5BvWEmHZPhVvy8/5U67D9mOyaIMzIS1
i2q/aYCCH16Wt2OgwVr4qqLrHq4hdbUoagxO3InIQd1W8NR75FZ9JFh5mqk09EKL
0wE0dflwLQtxZhlDYNURnktXhyJZLNprwp162EDepxWngNEoVwvnfJbR1u3LVT2K
hFagAh2gkEwNkd0ONQn588FivZy9q6zHWPsO9CQprixbdLZZ5P77DcsQxj2rCvDg
vKR5apY3XhEd+Ho2ZfbYohcfZKNbFeQBs0SKZtcGBUtBMeR2S2shErk0Gea960bZ
byI97a3IgcsTodNoY/s3pJCK/XqcsH5mY6RKGZ16Yt65rWCsTKMb8CUH6TaZFmsS
fiB4zOMLP8MaF6FHSY519l6SIcS9ojqS4Zxt7pXteOennbyr0z9j9K8luP/Z8+Ni
U3KzESk99MBxGniAdf85WTj2PumWZaPiri6ZSSBY1ULyh3P4CB8CdnigVqotyKOe
PJNnQcGmNVSFQ4XZxUh/A98Es09b9OFaRmDHE8s4zIubCLU8EZkKzuyDBIG+3kEz
+vH02QXCOfN5kNjZciI4w7puuHGSkA01bWHOnCrXzdssZfvfK1oovmZ3J9fz8c6P
55aQUmTsk0S9hz0fOFb+V3rVRjZXa+Y3dCAxjX4ESRsG/SprKnKpI/gasiYR+gTG
VvDX1+GpzM7HbaE+8cavayZ0IPSiWfbxxC/4SNcEyxyozpg0Au5/vEXETMarPB+R
kXeKqcMbsXFmlZiv1bGHC3I6O1aynptfTLB8fq7FDsA4dgApsNbw9l9G0hXml0RV
RHGfEVpbRjrs1EMlcBpX2w9y4szYLYFcwupzfbMZiOY62DxZE1eXE35Zpm3mIuA8
3/4Q1b0i7ZBV5VmCMQJQRuNdPxtS654CPugYwjy3FFSSieGfGV57m72eYdV9RlSQ
hB2WAapmWOybRRDYaRXzJnu8ydG0f8dWt9DNFRw3hl5ikOocWn6ey35lPFZANnJz
8nOK/FVDwgVDwhCEYM0xYTrLPDrMfp2C+lDe2gB/IfncyFHmL+HoxMLbeJRLYsMv
ayFkgx0jUqLS7K3rvzJA6zZSjPWzBDlsqH3VnucCYQUBaFd7m0805R0fQHP8v6JE
aMd2UXO4as3nLRBCGGcWlxLn5x7sY4jp7//IA50V9ON7KtUHcCExLU7rmUW+uf5n
Dp/UTocG6Vg+KjrwKKgtS6B4AkSVVaPtAOUlYuEPuQuQ4/kUVp8j+rtDs5Tx3RU2
ubKCpqt7XSTeCF0/ju9J5I052tMKI9bYUYtUegscSpYU/w1d5UrTWqf5uwZ2hR9p
tatMvJIEpsgzgwm3rLIJJjUTEG0SB3mFlRWVIxr7dcDDlCzEVB6vUN2VXK1fa5oP
bt9mr5A8wh7LnFEVzYThaP9P795u1z0HPrCpSBjaMoHjlP/yZrTPpkJIwUhMFgmU
ea4uJg83WqlTPskEck7uW+Upc/iDlfVsQY6sJ+CnoKfj8UjuvdlBQ7Uosd8hfwVZ
xZCKBw5WMQ1dUhmVKz3mCHXjSYIUbdJYeNUYLId78Q9eV87/UzGRd3yAQIqVz6kG
lveKyKJYSrW/Fca7KelW/G2mJs+3d2M8hs2smbja6NGsUCIIlVMLFlvbZfQ7VOsj
ocXrW1KUNSBOoHA8yFc5xAaEp0iltiALlPVUItJDlG4qdusvEGuIMHafRu/kijc9
8249N+sPgwpz0DuFqg3op3oBCo9LMgA4nCLv3Ktpzc7HqGM2x4+U4olfoV4aPqZG
Y7ZHVHLGkYB3DCvRe+zcA8x7JxSHNI6LcgG7om4VWruK9F81mDErBPEBozSfXgmI
rxXO0hBM7KIfXaWUtU7TsTpd/vtiVqCtuw7I0U6bbExJRbFrb/1ncX0GbpjmZPKt
XUeUQsENg4wV1AQ9c9hRjw0YNJgEW2+n8WuuA8NqaqZGemtfXytwULGnJjTj0ajj
B2ceumYP1DsVoWrwwckYWI4G9ALZXu2PQVGjoUluTf6o4gyErLUGf4ZBB9xbjBtB
4LCADXmpofvyUixwd8xxGVkVVTNH2M/Gnt01RMpRnmrSTTPvZQGpzZBJOpSLUP+t
zg7kKDAcCpph0K53zfaSiEOUUxCurqdojZjYRC3xFQXi3/rfWX0nfBFHSwzn3ZGY
Eav10d4RpT4186mzyxMnXQJg3VMhBOoMP2UlX5iJiB204t3CTeUinxnvy2gX5CL9
k0yNcyLtDapBXm0p6M8nuyG3wuNYy8Sy83Hd9SMbly3ihVb8e5JlG6TSZ9J4VUXL
M35bZZMd4daLuS8fjpgPs2tQGXg8MV2iikyrGQQytYG6GqZ0LrmX2gdmFuJ/oXlh
thouhu1+g33in6n1IWq9p1q7HWHeLfOtUCx8DXOKY5DuYP92xaCjRGGEdI124NSg
KnzZqWFu9VckBOM+2COXpSjjNcN/NLaiUqCFsjUi84pMGAN1mHjA5DrSuDobONe/
35K7cNQGR7U+yXEFYpxU7zW7///PfTALKjERYWH8ZyHxEtOro20OADg0T1562Pkf
QO9bp5SbfUVXlCoCsZ2Da83B+H2XauFHOO/e2+4WMGHkaQ3RbUf4tRtiWNcVZj0Z
ZCdfal5GX/0FwCkbuAo4eQQDdGK98mpTa+eVn/ZFJTNRV6STwWuBmFlmIkE8kgIR
wKkUy/rzhsnRJ0hZiErlPhyLSEQpm6ZFKZCRYQYotpwelE+TUcrYG8PBsI58TJBw
9c3Y7FXv0XRFj66ySfdSaGdF1Afz+A6ncz7zqx+EBMGMcinTiqyXwakODQ6bPZcO
SwSBB1Tbr+27jXxM/sKEZY7GzSEEc4hhYDKYlRUqJC0tARRSJ9j93Crn3frT7SEQ
fyMvZov5kpjvHTWezGXZ3l8MhmCbbBmaF3Mi1uycanqX/Xtw50h4G8M6YKbzsa5m
DVX94fLI1wOYod18gu5GON+HGR/Ys9QLkAb2tgwZXbPx5jiw7M5pwFtKJfnbxNWV
s6Q4E5h+UWYrbIFTxtg3GwegFn8e2oc67+36UnaLHrWiOJifx9MPE+OrVgR9Iqsw
i3vTq3ottIFmUpLXeKXB2ZLygEW7ejE8It8886wL70dBCX6kezQsDvRKSvVdULYo
SL7pvy0q01mDd+dwwfLpemyjry+07Lx3UjqwGO/U9MZk+spV2TBfUZSOwxdaZp32
9K8WeneRcJDoE+Mv6W0sIy3o2rlvvsjPYVdSKEUer025EnYQlVKnpi7xwE8Gecty
ieZP3KTNWOFm6feFmwMHZZk1d+ucoRuVb9fPhFsyBVTb6MFLoVOQzeeuLXfLSl07
GexEsknvgtDPT7IZEQHHohF/XTJcYSm5w9Rmbqyv098zHUNXyz1UmCZ7MYDgCdG2
JVilVW/TrNXTWxihhmjf6EC8UyEybU9qgRb7g0Wwl/PnqtQCSUB6MGD9pygdzKD9
4WXbGbqfulNf/TgwjlywFUFwVATe3MDp9oVWhrcqbJy4tw0pPs3jOEoiCoEJFvoj
uPDAHO2rPcAa/E2uFXlA6eCS8ONTp1uxQPLbLxsesr+lHPAKfmcY1Rh0f138+nqE
ZZ7W4+QkkufZlF8ew8aVUWgeaKZdPyngyHPEVLp36GbPv1yQwITx+WZrUK7wDYo4
1Uk43Bd4bJ3bsXiLLTORIub8U31DSLdIvvTsm6ERHtKTLJuw6JAixI3zKi9a+zO+
fNCyDpfhTa8IvBpdyC6l+acpcFfWDpEZMW1slmpoW3EVs2GEqDjPAMUJUsPTgNBh
Dscb3aBoUPv4JArLT9YIH1jOp/Xrow2KziLJVpLusw/ocFurT6ccVes+lQVMcctp
jIZUk5VbAWaxTFgTAJqN1V8xt4EPqJnwiJfg6ZX0xCzvw+4V3HNABcHdATZsJXXM
kuMhSerpZ+BF6Br3O63YaA1FXvnSm82cui/pYL5S42iKTG31kMkL4wDAM7EzcfRT
N4ag9yGp+gX8MzGnGF57rNKZYvw82bqS+2MruZAB8vjG9lJa6yzL+wPPH/ogwEUu
NIPiFDH5arfjXtS90V1LW59jiNujDq41eZYVjU0wQj+LXTM8o9hOLcC0IGNgkXKh
EIxraAh0wV6l2zPFZzp+k/T2rPn6kL8PYAGE5n9/yLAg0DZsCCOdX1biLNa1Sv7o
9lWcTNWAAHdtQQ1BAn4/nYfQokNsxH+EGxUXnJdUp1m0hYlijv8Fy9fiZLdsdWWl
8uQ0CHIrIgsDMELUHy0w43lkq3LokAHYvO5G1F4z31OQQlIb+DNzmEJUqV6++TDd
Aq4kf2KwJMeUtT62AfIqWeml/z4V6wF967X863H2bcoQaWF2eL9t89oCqRUZFzpN
Hl1RerhjqVLt2Oqk0XkzYmJRG5iJ63YIG7XAiY8+Zljis62p3qPLUUs831qOatsw
Zf9S63raAn5PoPsV8w+X2bmsedqY/mVzC3vYHE+KetEQ9jJkeX+1YN6oO7XveTv4
mP+NVLG/tF0W7SK4WbSjZ4YD8cNnOfNYlONTPl6bKEywZQTkWshno0Kce+4dHojw
3EB0kLvG1blRQnr/GPGNKRDw7H8i0/QQV5LkU36I1ECPal5BCbos0+e6ayS8I5BD
/OEB5XfLsf8QxZgCojCpIcRoY1ZBO533Fk12wIJkbWHRGEi1iXYsqvG6WQz77GjP
8TzU/jNsyvdltyFBdFH80TchN/M9b2o0OavV2D/1AC5+N8BTDqH/e/O+DJWGRTDB
qX0LpNogJqLvZfBL6unRoqCqtGh7TreRkK9Zhbsu0YEkGh0kkrm/Eix+KvEXYq5j
oYyLfrylJD2yi+GIcnbyZrPRsBvg3uYH4essBmCwFjsZMAFDaJsqeX9aXtxriV7H
EThm27kiAAcKlTZunU6JBZewEO75VLJ2nW70hWZsikGTVSelJq72vhkfzD8RKWGu
3uyIaQDaGLNQMW0DCfVs6rR3PWNl7jAyt8Kkp5T5HkiWkdo8O4hUuygeh9tbW0+w
UqZiUloLcRwcQtKLNGYbfLx4E1gxfNOMy4w8pRrn57qDxpcm9QzZZuyfiMlxknkO
/YfkEwfzF5aB9NayN8Iqj1/ZMPWRkJRVltpkps9eku/OkauK+Xh80FRfYeyCCBgo
MojAb3OdmGumJctoik2NaeMHZ+bmQeubroW/6dJebxGOBnrys6LMFsGMdUlY364O
W86DPEX5jBqKEA9MD+WRebCnBuzKDyIjBEdu+a7uHNvR2arL2fcuMcCp9IcRriKP
qBldkuKMFYXGuJICT8E0E2bN6G4P5akLC9aHHUSClgwMe7AxEljhzCyt5krCBULo
ewT6K+Q2vbEpnbolcm7QNrLP7Fe/cTBy+6ZM458uYJab2hlAobI//YfKzDAtpPTR
9F4yNHF5dfCdqokVI4qgGH/L81k8bnrStlYZOWzyMAdC3/EZkQAnVaAcHlNowMjD
35qtLmOUyN7v6sifQAgaHWKi0+p1Cqw41qPpJf3gCLs0esZxYtN0vAavqW6xmDL5
Hq5WMLCWCGj2fSTh3+TR6PQYp21bGuBjnboW/ISjxr/oCeFH31x0fzxsUke16U3J
p8nU9mt5XFFj4o+KFS0435Bqcdc9lBw1oup8E53crz56ZkFeUZdWkkGFLETooa3p
gDLPW3LuCzu+ohPJwe3sleRy0r7oRhhML9hL16zgLYVWqL2cDN/AhGtekXnov023
OrHeDtax20vacHTrGZqEYEPpBxfT0r1A8iTKhafv4f1bRx2JwHqBNf5dx9Vyt76G
4ZFAiHUkwSoYBSwa8grjibT95ki76FNkbdRprYp+MqC5MhOpQo7fHPWbE59ee0CD
G6vdx3ur7y8qeWlleFVM6+ZeKuG1dkb311RuLFY73OqtAdurQISY8ruAlpfU2dTr
Bdh/K/y3N/Tfd5Dev5hxWw90ZSj7gjVrBXsd69i4C2Bbe4s+DJfQXhVJaA659zXQ
o/kOZNMXNKpQEF5tmTvD6Hg4T8wuMtIRYbsxtWHBUnp9QInORJpnfyMzZpJMGyot
ElczF63H1fqJgwSslimtRK3LUSzuiovGJRUUNVGIhejDOJ/0yOXgzltdOfWPy+6m
PqMW4iQJhb1+M+JtLviG5aEb68oThzXsSTOZLPwFk96P8/e+DOiVPNi5pejq9tST
NSGphtjSHKfdOvPU1SPY6z7XrHVzgqZiuEZ16vQIOstigAIh1CSmxqa3RJ6pa3X/
fwsfZqq1ust9SRTdBBLVrwmrtm1sMeZLXQR9y6UTHxkT8s5ii3RFaVSVPpnjPn4e
cHTSFftxJmy1vtM0vzUbYZHNY96FJNtHEGlM03ZRrM5W8/DF+W/GIH/zFRS2GvhC
uDXoD7VSYqGdbOl2kSeyX+kQaY3W9AfGbLMb2ixRIUcjQPZ5E40VFiLO1iOZgDGd
tD2gXvSVaHJM+/oU8v7+CxpbrNvSuPpOliAbtwbyp7lkXh+jtiMAs5dbw4lIy2cS
cJ3uTHG3NUYYrIElPja8nfZUY0teWxYXbyrzTEOaWgwgmlYxNc8dtPkpOf5p7Rgw
6U+gqu2JTcV5lvKjVBUeYHYInQzCi+7UkZZ0s5g98lhtHvvjnahxyV4tBwlIj8wl
xJSnqBOBMaazNfP6/Omw0jRV1eAyY2KuKYKSJOJTAxr+D0hHgk9VIfOvUMh7ri7w
lWxz53BN2xJZUJORH+pEKTQ8fFfHuBMhr1jmsnbtHYF7b5/Apnbinlq4b47ykPXS
ocMqfNmPHdIaP9FQeTmtetoAHjEVMgNtUKsJuuPOHdk7ptVATMOWO0K+EpwI+jm9
8T3IHZEa1fA+qerlUoFQGZ+T61o4PPLu1gVIamsC3dbdTauofgEUl6+1GcZYbu/o
ANRLp2VvHGH6q0WiLrYYVzbiZ6mMJ3FFqF4cf5us4nHxlVgw5np6g1mqXl4Sr0JC
AUe05mWUE/y1Dr+ZZdYOVGwczXW2qiUkfl1t4Pz5iyXDuQabaYLi2pwf4EUFaoR6
bTjii8giB/IY1NhELpYibVM+KdwQ+KwKJd+WpCvSjZxAJC6izDLHAPeyceFSQDFd
Wz0KX/PnQepIkOOR5aCQqnKIRrBSSj98CQaBUanBL/klhZL9IOFvgluXPwTLa4xa
T0EYoLLl2vSNr0OCxoYwmV2rDJ6nMHJBkl6/GSEajA9OZp+bzZ64ovtjx6cnfl5F
dWmdvQ5qJvz0YqY2jkrqiPyRsRVcctCe6BmmKZwrcmiORjnSrtXVZwtHO2FhMBqy
NYSA6GZmoOT5/SfY7t997GqUqO/525FQOziRM6yQgu1ywtAZVBJH7EhN8tL+I9oM
0YD3Ar4UVF06Qe9z2+NyRc2y9mDNhf6/hyjo34vknTFjZgPPtoiVGkJn1mBVzQBG
ab6DBCM14BB3SmN//1NKqAVRu4QS4SEruavNVO3TdfDPAle5xyODiwdaLwEqmdsc
hzClk9A+1n5LOgbn3SA47Mev79bhKBmy21z7PwBW7TxcoPyeyQIrET0UKnd1d8VK
5HF7JjzZbNNwIC67WtDVlve5/uzjwACZ0ZrWhv0LvjM4UVdrGv2YZU4hVTsMNIZp
yA3dX7X2JCcQmRhEhEPJ47vP5p21/94BlpkkKfEd6ZJJ0HVq9yXewuPYZK+Pc5uL
YKBe0V1OqooHSCBsSFgwmrd/JzrSRPzJi0XPe2omsDZEqhpW5l6WkxcdO1cb4N7H
WQcn/maJ6mHOfadAfDR5kKH7yivhRnS0VTb5zBwiLKtLeeqdOpUmB6Cq22Wu1HNe
cYslXod6BfwptXWksKRPdXqVMs+Y6IQEgEA39psyn0hxNhEIqwqg+ZS08iMEc2+z
x8MziAGMhe1KeYFaGjYlafuGytbUqfOarK+EEbSKZMtt5NzEm+DLMuv36P24aYvK
MZGjZTZfIf0uVNhCfmI/syl18E57A2ZzzA86DBFmGwyMCWrDknYNCUINMzlkZMAw
a4XSkIqwhz8y5S2SLOCknMa81fDf7ZnZPXdHsuVuL0GoL1o1OQzdSeapnTpuvQB5
5qY8vmUDXJXT4PAMlFhUd2RHMDww2GTLmmgkKQAX0h7RU2em63wi/XQCC72Gwu8o
Ve53dQBcjy8Xc5VlyQOOhfiFnerMedsvrNfom/flY0Q9zsel3swT3R+iF6Db5RFG
vVYhovKcGiP3jyb3FG/EgQTS4TMKeKsrRyrSLc9+sw0q2NWWUMfb4vBuJ0P9l45G
WiDYcp/NfiRBnwngA1rFhQNMiiXLqoYzH4k90Bl4zFAvWCYswv31XS1R7nMGER6+
0rWPsbOnOeGkwT+osAvJ0NLxozZMIf32JDuzpEWddNorFIR7s4Sn7sTttkYTHEXe
LIPEanvCJLtlesggrmZnPtQv9PIkDLPhf2slQhc3rh+JnOBgMwhPmiI4gzuxnuU5
54w5MvB2DhEeWRZCybHebqkpONBrSi/LDSKl1UwIuynhu2nHeP1AotqqfHmtqBQ2
T7dflCOf6VEM629Xku7SAMOGcBOtiYbe82qbBgIgeWcVBmCDmnGFgQMIOyZ6h4s/
6xI6fG7Iw1gQb+1CRvKpvYfdi5TEXBmHJZdqur0ntVajveb9PHUa5mRIcGrDF+Sw
KUdAiHNfVY4g80hly2J6Z12vuucBxtoG3jlDfREBt1r+4shSQ5b/j7jlTUKW5hMi
qPm3wRxL82oktRQOL7uK2YuXuzd2c+TJmhiaimf+zEeMdPsHVoZY/3rCgUJU+np4
/w4Vwdai2dGyk7UbIEJgCCFdyan177qDO4T47fGCEBWYe2hEJFNTtqlQrFdSfndn
2BrICX4yYU1fUIFa+lq4Ete8eKH6AnonDqXfJH3QrsmuGjUhWWxKnKoHA8QD4bOt
xoJB/62THYXkRx67uEOrgGJGDcqBAxLtkPTEKpIkljfAfJ8mRldwIEQi0KpioOh/
UD7ZBx6jQv07zVwYMBgVRZ4IIeR4pF9gCCEVTIlf5o0yem33Pax9DTu0ikoNyvxq
vb2PyPNKPIHVHrsKFihmXiMe2+YFxrM+UcbRB3Cv3RB2Fjco+o5PPP/w/2V3kvlQ
jSwyUTLHhWii9sqrrmCstpM3hr9e5kIJLEAJauwkwEbxh9Ix0CrmI5Fz1soewuRt
o8NwzWyAmL5zR8nY0vl+OBbHip1Im6Ah8Nf9TWHEUeg0XXSFuN92LAXYh2ozh1EN
V52PLgxGda7Tog+0ILL1yXrDROqj+Ltkk8rwi+PK3BYYEb6jfaVYIstyheH78gWu
QsJzNlh9P3z1WN9y/+Zd2adP0jH8cBpzf0sPyg5fXUyGBx+zPma5Im9HoIpGX2lz
lcwXldb+RjAeUfwgoPdaHPlwKxnSrWLpdkSWw7/fj/G+UqNyoOG7WQys85RuG8Ba
3HCMztO0rEOIBqY15n6S1VquD/NecnwGh9Y+IdUI/1sWcFSfJJw24OMj4RSVzsii
zL/JyoP/HSbn0gn9fMwXG4aoyb9fD7LUdYLI0PBRF0v/ihGwjIRvpOCzHOIb7On7
ae5lSk15JeaO8x8mwkPzaZIFUFGqlwOwrJ3Q9OU0Wx94unhbdoXRQTKmCJdSQ9sG
VexmgCqNa4HYAs8iRXC3yG9ktCxGBBpLI5pdi1YydVnZT/12Is9y+IEbATCPgieO
xvUMZ7tTHNYA7/gFmzlKuezQ6IRgloEO6ihh5+j66Laho5eEPk7JKVsuiJag0Jbn
wG5TNQ/twogUwvjodYlZphaO7MZgtdYTDMXjctncQm8PrtK6a4YdX0x7YztrGddm
x5Eh30Hhnc8gC6L/nq1SksD1GtWtn4YRWh4lgHOdfVTye3Ub93vn0MB8DG15vWEe
ZT3twuK7WvErxyEh3xR9by9i8C9KbABI/OpLRt44iRG9Z0X+9ItThaHB653MPsOO
O3MrKMpo3m3ei+qYdT3GCb1VKK5NXBPTC7CkgaEd0393SDkERGx0U3NdYchd9GQ0
GE2Jfe9nFb5LFQ5y17U6jKcmZNUoO0erjYImNzmpsKUli24Z7Kq2jyU4jgvNwg4m
6d9LvRzs3WryO0UcDpq2WQRZzAj/zcjHDFCe/v90fPmCyq6QgrqTGdga7KoFYAoC
rpcoIltma/Ko9y6IBODcX7/tK8RMiOT9yCoizXuhOogBp/WfI6Uv2fvWU2vJ6epN
gJ3iyYFfC7eQYw+LEa145Bpta7pr508l05REPeGMd0TsBLFkhvM3ySU0DsPvXbKF
4KHriiZ0XZ7gj/Wmcbx02J/w8X0Sr0Tt0n9rlL7KbZkjO5rtVyK5d5Lq4eIwi3sy
TPWpj3bG4k4Niswo99EfB/1GehOzQyRDOE1xk/uXp4PNinzgvy9TSGsPPCMKO8Qz
zl7dl8o2t58JmjIHzzm5ig0eQ/zYPRu6YCIMWYP5YPfQOCM2136ZnzWk371C7DsN
X3uXYesbJ3scgH7bwD03a/B37ke/VbrRRy2N0EKw2xa3kpugd71w1f463EIRXDLU
BsArhU/bPHSbIXu7nzDd1YkajhKdQv1hNJ27gw71/qHNGcSRXhbr7oX7HOd3qd+p
PdMsTJiqmuZXgjfQdaLe2F+rlF7x9D84kbCSdLdZ9BJVxfFpFnM65j/l7I8DE7ei
V+Zi38HGwChvqiDqDcQ1MTPcym+d7FOL5sXX8l/VEcVXUdfCzicbflvH4cKq1HAE
dKIJP5HTT+ISTzY66vsIBAdO6Fi3JOoZmx4iokRi5q7QwVzr8CuDbz4zhIuiB6Wt
RYxLGDwGi0RaEFmzcaNP4qq/BDFnLDHw5uW8jOItS1/XrrhJQmMs0U0Xo1QjzrNx
TkdJaC2B5idG2OcRcOPITuIHO4DwQBA7ppc+UoHciGIOmWvloCoRELuGpmRGn0BX
lGGWyYb73e1deqbme+aflgR0E1oQqfMFo0SyEl8ZCxW4tZowzxsiZ4MGD7PBwBlO
XYptqopuTKHAg6vvcNRNoJsYm+Ao+w32SpPRGvgMbchdwdLKJCnApyfPghfZtP2Z
OyXsXmJKTkW2bpjxhuQAi/ab++B/doiNSU8TK2L//Nm9d+Oe2mI/fpTbfCDQCTTm
nskzFK12cGxViWpc46a2tsic8WxCzZ8Phwhdj6Sz4b7Cti7uvooSRob4ztb8MJO1
2lMSzXodzS0nNZOLm+ISrDSC9gNQVTKaX9zfCgZH/bJDr1/UOlufzjBXSQn83t2G
yZT7qaTG/7LR4qtfNlhQGEKF9tiA5ayvz+h9uNVgkSXqVlf1ysxOjNmmdG9K8gFh
lWDZJ+hdN0fE2/9ENT1KTPc+LtQUyZSBJOBJ4VAqahcL8vsnsThpbujQywX/WJYS
DC0BOUur0NOVIYMFh/nfyomZQMK9KOqSsq+kwjFBgLSrh1vQUlViQKOispNmHa32
8ybcnGaF/7r1LLwipBpAO2JesJdzYK/3bvgSXaN3xNxMabZ2OTIpleYNCmB8cYOu
IMsJpEWlHiUyeT1MsTU0QUYhYspL8aAghUg2pVNGtZKM4AfXoU+I1puR9eWkcoBx
YWxnoE4KyQZBv4e9WNQgDZOm4E10XycMy1b90KgUyE9odF0IXV3qFbYsVLPRIFLy
uCd7kitJMcZMNJPAMuzULShSIyaFBpSs5UwAUrut/zLlX4unJamPz1PObE57la+h
NMuhbI5fgs4ihM35xgzOjpSv+SAh3DQSELJCtCkqgLh37jGkUA97JNDSCDMoM644
FahCg6Cc9fJx+fDW18xKs+Xv2MMKrJqfDrnWtSL7I5vSQ3rNlr41R5ROVhM/FhNm
schsCwuWQnz9+oN4BlFQAc2Zmso7qik+UG8yF2b5Y6VsRin1Wz7K3k8gGhkQwwQh
W7e9rjW0rvX+2ZKWkPe0PnD3oVYr/1lAY/2M1DwJ4iM/eVXAPStZ4O3SkZua3GiU
09p+2joWXo8VvCF8/caW1HD6In7+4OjImaeelfinfl4RizrYPJrAi7IA7ZiFX7Pn
tSjM19SlK8yowpO8Z7tSQPbArtZzeOiyTtCW4nXIaAOT8RveQWmaDdIpoxeAHvCx
lP6s3pOIUYjYCINN+8zDlZ9FoxT+ugXEcLgtXEAetcrq7Qd1OsT/V+ps4oEOhXrx
2l/ID4tlhceR/EPBb+h5ohiWhUQiDsZrdVFHakqKbrTs12cDZgUphO/vWO/naCzH
8PVnfw58uC/4xJI1/ZNfs7ZuCnRY7e+RWH16ex889yWcNoLLACOpMD6GxaumEA7y
QDLJP5kxB8LbCX6k0JanCAsx/5DcrJ/QlQYTuu+c4h4+d6RJXXG2giMGZwJwK+0k
0b8PYyPaQtulPCItbq1vPTevEou1MBR6tBakkkacgcQK3+CJkgxqW1DVPw2nzVZN
m745CZLcxXALC/tC/RvMHORWk6xV+1w3ulNV6glV4z0GdZBxe8NrJOd1tLp4sG2T
vY1QFcqSwUofSpf0VStg5WVNl2zYBrLmLEmcdYrVcaSNqJSP+LY0hLrexNUBYyjT
XJGlPBbsnACIvne5Pz6A3QB/YLVL5WtsVMmOe54Kv+iv0gysXy+OiNa+HbIqE3Ez
pDZPMwCh4jrsNaDzxjEe0BbvnX5f3+W9oawxRzGdTCGZ9tTxzsWGZAH5xdbvFRDL
BseypnUHs8eQEQOJBaGL1qEO1PUHBZTdQqKUJ6VrtXxtFb7WtEht977gNpq7vYLc
/wfUUx+yS5N7zW3yc36Ui5wvHl3nn7lyoe8Km+HpMWerIglKG1xyQehPMyM8zIq5
T4LhTNHtAkBeMDpaPrPhC4oGLhBWBudvfzQai6xrY8Y8cWIIWGECKKkNvTaFOjrX
LPz4S6AxxU23ukXyepg5/Pr31XWklwCTZ3cjB66MWw9IJl3mmpdNbex1KHsLzOdO
zHjkeYcfzKhYLNsjQbKn8rycMKOLlhZPxiaVEP/ubanMnEvmAhtPCZWRy2KSzTgU
c+1SmbVWT+WNZhzbph0cSO+rQwBovhhhSf/9M5USbd6Axz+juFWN6hCSq63HPX1C
IetReRwIhu86MlosKkm/EHvNd02jMbWMMYGj/cZdY60FKgRm5KtNQzCLnQ9f37Dw
gmi5PrsITqDc/vCqrtg53HkD1jSy0L41enl6BJSyEpij1xZ+1d/FGKhPChavqfte
Ge9cmS3OqAmxCmhhj8rQ9M6V8rTXW1leLLf9c9Y4YdNITI8GlkEAnZnkYPdw+Ua9
5Wc6hNoIPK4VrYJYKgqLhmmrd/akWLOTNE27LVoxkBfx9LWzKMqBC4Lr1uyMdZQo
5jUnQTYBNuVB8ssW4eJ9wRZcfnCcXFBQr/ghO027DJjFKaGtdvaHFaL01j+d2vQO
VvHh4Dx6/GMwZTfYETGs3/DRV6Aj1HbNEVeiebGhiCRD2GL51Jg63MXUwgfXxTTF
gkvupqnuhfur4TwXsZL67ucGeZVEulRU8cJkBT4KhkjGCfGCmaDEHFwkzZ0X5Jwd
s67I6lizmqV4nBaZxpbTaPvlTPP6hpVgWTGcV6W73eKlwtRe3bB02RQATTRTOS6E
faoffpOc81q+k6hX5rIywE0869K00+/Vtc7ffhzCVDWLIcpwkSFaxnqak/JmU+BS
TkVdR4bxAOAuB1uuJyfpXu2Q5aN7flxfMBKn0l70ct7lj/sM6Pe0JFo4zwOQyznk
+R2SSeGdO9nvyYySdYVqIWuPoSAXXug1u1/Bgr2A8kBVGoskzXxBCtiWc/BEwBnj
yDwYazonvDKzbIYrMR+382mAcpa/Fv++LfMOVVAhDWooysl06G0cd5en3d4yVryl
/jWM2iu7CZ1LatGaQgKEdnI8ZoZDpJec+GIfZvvqJ6Kk7cPvbR4DT7JJ/dvQpKsZ
OVhyiL9kt89hv5jZAb4r2GjPWUN4Zt6UXM4xGY0Pe1NC4GhN4+T5+PwY5lbFYXGR
DJGY2pM/FZjxYKxJxqIxtzxfkdQ8bs1K9EJGkoIjuGxUj9eU9PctdgWVntbVF1C3
OZ5EbeZkUwO41VlVNW3Okrf5w8QIARV0lsuzV/OUWfm7zOBISuPlolylTVqJgZsI
ARLJdI1T83CqWEGlVRQiln0at5CdItOa8wOxGM0PJWklVATs76VrVYnfx+Wx7Y9X
40dga8Ysu66gj/Dws2pdWpHG10cSk437h3ukh44DqtIKpQJaiCcN9quLr1ddYRiK
+6u8RG05e+WFADYs3JdQDtpQkRE6I9HpyJd+35Gv7A3WmBYAcDLVAFgcaIxWdm3L
g2bDORuMElNaZuP+iKKAbBKEgvUbMQ0bJ4g/Md2BjJ7CU3YtcwRbewx8pNr0Gqad
nYtrCb9o6sx20Y2DHTRPOit/lSUJS2UXnRn9dgJbYt9WIaAyrEAGKdgH2g3AJhsl
ogbV+az6rcPqFEboLRimy8il9e+5yVmF3km/fMdJLZqBZdVZZ3s3/xb0xlGl29Ga
5q0nsKGc+GWSo3AZvu3FVMKkY0gSXJirMGbvqezsvcvgTI79AhHYZFZVjF3MWpGn
15T7aJPktUDWhJVBJLJ+mcbJAtXzOGxCb11aBo+H51Lz5u60OeSULRf6NEazx8Ab
ACO8ZBdf0i1iyTzwo/7OHKoN+TKUUwrH4/mi2tN3Ye7LJzCUG2kKe9ePvON+njc9
66VqlT4KonHlehT74vSeEM0eNVm8Wmnr83CjkpXUvjasrsh0UQBNpdyv2xCdTo2l
OV4bqTsgelHyO4hkkpWkqpucgixqtjCpuO/v6iuSF4dk2sKVKCEVZjsS6l1qyiLZ
UsaLgAsIjcR+u1vqIkYJNAUEB3EYJ1Cc6cJxa0bhxfhDqWkhEf/HuOCg25IeeJ7k
AxOIjWwnYEEweGkDcNXGczm5bOGQYDG9XzyqbNJfrE0SGUOGW/43hQhBfQucvmn/
QJL/YQRejOk1OHdqDqg6bRp0Fjk19nmiUNuzewQ5rWF6WdnEMd/qsL2xWat0t1Wa
2DC/5DmqGAOmR+ns4acT2KR+EdMWFh3dtBKALoHWl9fntbfudduZ9AqP3OAZ8T6u
Gkb5nkz12meTOK2IDL6ZIy1FHKa91Vp33ym7goEjWSm5FR3q+L5dlu/fLUeHaB0P
QW10eCA4rIucEvdBDnq7y5BSh4sArRuea7JmCnr1BEfrGNRAdtZU7klAZX2ioowt
5y7lv1cyV7MYOXGOGnEXiYBdBe629L4Mt9EflefnlOSOpK60QetgV33WS8WmDp9p
GUiJhqidNuO9wdaSi1nvTbxa9NASIeUnf4zmQt4uMUZQZGsrXaqUW/RXOUFlqwGH
RLuQW3xtRV6tKsPhdFpGbqn1tR871r06xJ2+oHGeki7PzJ65hraWxu4SRBgMjUrI
a4P07RTxnicSWOaNT3VAG4zPQpvlm2bxxk3x2LXEVgaHbgAJcB90i8HjxX3lJrcM
xA/0jp7sNMoy07dJCcBYyVi0gEx7rz4GvtvBFWKna7YFE1aTSw1gXkPkMilMfYzS
6GSGDLViRtU+8x8+zdqS11Y02uK72wPFUk4QMhKOkKqjh3toFGhyM+XSIvDsIFQ9
K8TJ2vvLBwTBTtchKx5UC+JSxtim5LuqIRiyL/RHAr/xKpa+bZcN46y6KRnavlQM
v5Q03GaJ+AI1cAAsnOVpQOVmZTcWf3ibi5c7uAhMyQOJPLFYMFkr1XGGzbjfxw1p
PQ9+qfSTeGzOOSUg6vEHzDgKAx20+sLdsNgilmuRz5SnP5fjbooF9PPHX3RMlGU4
s/kYC+O9mvmkeU9sNdpo8PqlH7lNLgxxtgpx0WGaR8NMjGPFQeKPmgxVD0aqZg4V
oFuzc/8Y3BrhZhrm/NEK65FS8bVMIeeW2dsmuYke5clvCov0LwkCCWpeS6Dtalxl
1cw0I3KI1uE8Waw5OKMn5aUfIszAjhUmRYtnm0r3hVIRsbqsQQbX39lldC1XVun5
oXHsq/aoyk2joPcaLuXV/Tsc5oAN4aEMgW2ESLCFIT4OKceQF4Cxy7mccXHwz5bc
TYLy26lXEuaA9i60mmZQrU8+KQ19HPa4lk2BbbL/kzb6zhGiZwv/SHprpbrSiOHC
Csa7TWiGGJtDccQdIwPDbBpYcOCxaVrG1QNjz/T0ItwWBF5CIC+f7vNCVY+Va3GU
RLNV3RehKga0EqzSqTG+XYdlhilG4fRHF8aHfp9QpmFJ2sDsoA1aG0j067Q5DMEu
KIr9Akzs7jism8b67wH5EYND4D9Q82cWOq2J3KDo+3llJ1alK+tJcVvcFIneRmIR
cns8n74FFHx5FNR+HEQFKjfKb2jvqexj06vwZImDtKwGG4x8PWMZOUI24xrOgwb3
lw4Xj6aFBWCCYqU50gAtjkeNvXNdseE/PHhzVVHYkbZC5PhV7PoY4D/lQR4R27r1
DcbFZaz1BBgcAKOKIZ1uMpuhCzmZ0pGDO+NxctvtMcZQTu24sKYlFg6ZHvf05Xnz
KlbO239MRMz4pqJKBle4i82d0Eiqrj0cxUPiY2ZOMPew9aQ4aVU7f4ihK+XPOPQZ
+FGbHalu+QNNoMgCLL1LYnCxK6e9W4QPJDt5Fm9DmIpwznr0xU1SBdEsqxl0RD4d
TVi90m/X6gL11pZssmP+ySYkL9f1LT7Y/G4VE0jdBUDDUmIgJiJ4cqOq6O46OgRq
83E8rTAJT/MZm+hKNhyjKovIdEZTxHsSPeNv9EvLzwokPFp6YbvXKCyTNQ62d/2m
bLIJuA5GOH+6Rc74F7dny3tnYk3Gh1PSNsaAwt9VkS7sPXFHYIuXBdC1gU/0bwZW
jNkSJS3Ividn910cUGweSrY+pgT+EkmjcSE85LwofzGpOkOIJqRE2NaQuW1tMsTY
7yLiUZXVhXyiOAYvWGqBzm8ww8RYF4829EK8Vi6iAnRX8sK+hOfzgeqoCYK8tNxM
60uWg1Y8MTyQHocYVUnUPjCADJh9M+Cggc0n2dVehnl6hLM+WpGYlLpgn8T8YKPw
inpfYvm8GJK0LCz3GYvjKn6c1j4rsDnmRT3GeqQQ3omAlhCwWQ+Ce4MKBDUS/bgC
CcBsBp2vZRzpA+nA3+0RSToq7vVQ9dmOLTf2sAfXF0HNkk8KC8v3gVDKF/b480mP
beY3+wwr94DkmOG6sGi4P+dqTxnqjkMLyyEHyQGMfSfkP1k8ZZ0zrcMlXf96281V
uWQuQTEx5T0gW3s3THBSGjGYCZyXVAQrUfP8wzaR1lKVjvetUMba7gcX2CNNxOzm
RunZrw9crGkDwmLvX3SStZyT3rlo9dDPT5iyOwPvlZVLCVa88K+HpHYVHCYbRD7p
RTEuxLMb+XMtVY8e9vkx8f0ihhAbQt0X6s4xIl6HJBcV+WNmGCGzwVCXvQHIZ5Hx
JsTNTE79u50UEgLcALlorg2gnZb+JOqCFTtcj1nP3DOzml0QwiwWeai5dc/a5Hkv
0uDtvAg3NH+bhir82xBQcVvGMC383RiBxrFZH6PnC2PFdoh2hVkcGUE24bJyoemK
7Nb3lNsF14woZQKPK7M4tZ49iwuHnb34RtSDBBzwCd5yaTEctMc1bJctNy1pmSAl
71RbBxk+qHyTxo1mv0E/pJ6eEzJSznHfY5GP9b2PhIVJ1CWjpgw+YtwVmB+dwfWX
4+A72XZoa6iLFIE+XFIZEllkmVkNlHXK27zJvNyfOm6taJfqRO6wYrIK0WAjJ7JK
2WGdGa1CCt9WEoaMwKxOMlyT2vpj9ArL1JaXiLMC+qK1R+ZVAFUly4Pnij/o2toz
3YFrGD0Gi6rESFv5Hgqs5mp/xLlrTG4FRp56LWTWdYdWkcSdVTU6Q1BC6biGrx0+
NgSv78Em0I8RG5qWMsnN4XG6rD+GX4efG6goSIY5w1oLr07+NK0QGm8qHY3Kj+pr
vBdg9J0eMLRO8C1T+EmbOLzletzzYuHHkDaRqhORlHPC1jEhPPTTZ8vYJFi6c2JO
bkzbydQMvLWCTNi4yk/FH8CsYKIqhVvM4wth9f51fwo/PAX6YKTsGCgjgLQZvHPn
ms1BKN81byzIPoPFYai/YKGemvg1vBYFx51eaHyjoKb0IjU5CSfk6IZGMhvQrZ/w
rZPi+P9+PI/W5fYMFoas76qMtJZzudszq122GSjyxfrb5zaJxnKCuTXr4TQi2A7n
3fLJ3lrLyNCLeDj86J7slAdtGcvV2AbDtojQPxI/1DVaEAhjQ195BeKJDYgYGTwV
svYMUn6JDO77aAHFVzdJl/NB/E0Pg0oGnZu76s0rQcBEQ4SV10Po8mCnqn1YqGsc
T9BxYgJMBmSLhBm0aEh1cH841v4gyCFsqZkqzFzz9k47C2/ku1F0P/BS7L7LcNDW
O+ffpw8jerhHh2VJwxt4SRiduluZ0NnPRnYJ8oBXKoj6Zj3eEecSb7hCO0F4QUu7
dSTOnAO8IjXawBa6qliHfksyWAkh2DO47Zn+J/Xw5CsgepxwthQTy4oXV1jb+KJn
71INI9uAUYHmh46FPWrXLNu3fzcf8DaEWyTa/JBMBKSvi1t+eH4V0efhKzJidxFX
/eCeMNpUD/sCIJ5Rczia5ZWqVYnKSEbInYu1/wDlt0+L1mOILkBA53ix5AJFUTK0
Q+x41bXXR8WX+SARtUmyyADmhIUAchCx96tTDZrfhbL38ZybTEycsT5+3y2TpRfZ
7otp62STKSLaFrB3UN6u4wyrIrV8OxBzPabj9GSJm90jtstslsFIo4e+FWZ0lD0o
o0089E+w7t04CCyfa1r9gbryQVO363sGa2vJz+OCwAGgjHTwSosngQNImU2EFUGu
3X5T01XNJkpj9WYNQ3SyOiB6HI1rGOg+hkkDTMiOmU1AksoGkGaQIyxrKOjVkXg3
S1g6Ee82I248v9B8Dup2rvSq+UwrpbdmqZTeGGeA28RSav3XQs0pNwuTTQ0yZXFJ
Jlzq5dh+VovmKv83R14yo+pbV/pVsA6Qkt9mQMX2M3WwU/7szd9FIC7pJI0QohR0
Pe8DkML1inarbXiIz1cswO7oNAq7kcdQSOoAYv9uC5zxczy2LJprgLYCPSF+LUUw
sbjiWVnKF5hsAPIR/n/D5shcnVThP7gC8TVqyh5eLxBdSX/cWgcKYlcW94q5rxM/
EKgtrir+RENdbZ9HVF/ihrESPxMR9NP9g0AsgRvuj8f9O0UyViKvrLIHyqjrPh4U
PmEOncGibCgSu1qE7hMg1oFY74J5RMeA4nci8UKPhxvex6tFz35SEYyNYC96Jy0b
bgByyam1aO/ylbwKSEzvWuGux/uwv21H+tnTi2mJ9rm2r3XYCfWpWJgOolqpPIZu
KMIV3yvZ6BFo4P3dPiBKWmtImx1g/L2K5JJZ9uKkFWtUn76gd/vIPFV/bqqsE0Yu
CGL0nJagDTY1lEjPMOdYNh4f2Bb5KRidStAENTDKWIUItTon7/FyJmw9TrOVR2vg
CI3ZxWjpoGcfuP9Mv6lEkH92iRNncSwJILfMLkEm7MzEfaeu5qiFKai2bim78RTm
eePHC+kt4SChb8N7uDYYGOur1j7kwKdqy4u3sdlQkkUHfaVxi7aFh35906jnJQJj
8p7I77pawQLqsqhnqdC2CkM/k36J3DMHhhZKMja3YzOUXuaOl6QXIevBP/JTdryn
CVYEqdWrM//WKdRXnEL5F9CuSw/kVOUwO1f+KymKufXJFFUVIbyYJinV4y8faOIU
rwZXPmkcVMhpzCsFi2Ar+ih2aLL8fCyiZUMJIhBCzPUoG1IiyQPtgdlbom61mHC6
k3CHJrsdQ3sNz91w36b8OcoPKzZeKXJVI8cRir5ewcS8IF3Gp1ZFXdPHS7n6hn+f
dWXP6Wy48zFaGVtXoAOhrjdCsrYbfhjEjpcCOJQioRi+CEpS3cSYayblB1pEBpMP
9aJYpqeYLi3hHBzh8X1v6UkwiL4EuECPu0jABig7CjEDhWb+wiXyRa7DF6TvhVaW
Ojze1+0dcPVR0is2dp+P+1vGl5KeyPLOcW4FYIQJiczzoesjL5BD5dOAWn41wy9G
/J8vJqeZFi5nRwUYkr3YyvKrlbd1dwbtp/UxEByz1OrH7/s9lgG2SVyMcPo1l3ty
q3ywDNiCpYB5GCe8fDmmkYT8gjMMDgay4rkE4cGJp2KCqJ7N9zGQld4C7MVcHijc
dyapetokSYJ6kd2E92VnPALzS4lUGN6wV9JofFPHmCevQlMPvUStOuFKiHr0ARDd
7xh59mn66cVx7WmWrwwxQXah/KPpmpqhG/mkG3ZzOK40UHT4ZpqVthERkAPjnufi
DSzl5SxEdyFuyvZckIixfqXnYkK5QSRqDN8nLMLlN3DcrAVagIovH6JrdPo3YFZU
ZLkWAOMEpV/gdlnmg8DjPcRUfD9xNZEnB3PwJ8LGi/T5pknJaMaaWrw1pBbhzUwU
ePSgMtxeDXUqQa6dSYERDjLfiQ0yN/sP1Eqwi8lkqQlR3kZ9RP8MSkZMw1THtOGm
IOTjXQgrfh8QTcQvh9rxxPAjzkarVUfOg8QdtNcy9FYznxZycyn72U/voDijh738
vXHq8KGLk5mwnqtkEEviTkC3ssddhKbGFkYVFoCWTiv8KPapSsXbpuG96XF/xW5f
20yoH96Z03Ncskc7KcTi4aw9w+38IHPcxTOJWcIqzOy+MxoJlwX9Y/rVP51hMLTj
MzUnXv4V+YkICDL+fBGtSAe/ILAJT7vfKhyq4o9mh5BsryEmWINMltyJ/RTHYSPf
MtnFMy2PADx+OjEmINZyq6+o6PQwikc8m+efo3j760aYmHezKfJc4qvCJdX+2cFC
k/TabBq9a9DpkHZBY0zmzKnpxSsvpoY2zt/XIfDKlZJWIDcjyKZ5iyjReM7RmZep
nB+KviwsfZmpZhpJcyVfxcBrR8xU9Odfm86jdg2b1gezJTyfEHIf7A6ouWZnDLx2
wbUa9nG9IlT7wfPulnCpDlCb1XsZd4imAmbEjp+xGLE4JvoCbfbTfYyMp9qwKO2K
IVOhFVBpcPd9BGFtmfzX7d1bAVQog6tpERdML9f5ZolFgHSqEPnPgQo9W/IXU236
FyDi++hDbXWYywsJgp6cU3UFByxnBkWgKpOxoRy8Yvt2EycXb3gjcLnHA1P9xPRk
NMBrCX2CNvVtrEQ6VZ6mywE3i5tgNEpWXyXdhKwrCuIwUgIAfep3gr6Jf4Wj5dyX
waYaE2TpO+QCWpqVNUKRhzGL77GRPhoCxjVzcGWmzymwOXPYk0LaEkECxFoc48R0
o5YuUpEthB7IeogB8ZXAUsDI021PxGt1Nrz+IgeuE8TheKZfygje+9VN1xzg5uSb
xNJHW0TRvNkvhdnJifz/M+OCz1uo3RSMctx6LTju2esfWI3WjbUFIIoBVii/QWtE
FlkkPPZfANMeJwPIXqwhtsRWAbOGmZD/Z3YTfSojgHufzAgmD0mD1wPHDvhK5QPa
fqzJeTsUC1Qw6TP2+yWQ8UG6Iie03G6qvmrCQ+nuqJopRSTkarXiBSolAQrHCWGf
qVHYJdgnXBLvSzBJ4bdTWOCvbcM5s1xZy8MMbiD5owi2BCZNj9DIc2JuOe9FxHEp
lv2aZGFeZIOFFSTBqXskSqrmhnT01yNVGZ6cABkCqC6qbXTmfN4TuMwev7XkVYNJ
jrOhe70KJ823djVe5k+NedjVXkG/U5/dGmw0xSVNmOm4B0PbspdHwfSsyzLZ+0LX
HX7SBeyCAvEaKopLJeMmNt0QGP8Pa5kSNxZXtZVc09XmFd2U4BcdoOgv1ZCHRQGK
PpDD/1IFtMDVkZrMD9/mie7e9iOGHn49Iu264EH+Cf7KAF93404QVenZRR/W/YJ7
mkKIPiLRIRALu9JTMW1y9+gCmezWftdMOADJpczvsagFoQ3m8KVgW9ZWNeR20HPG
1RmWlDbAClOie+r0V7wMItxHroJF7O3U0Kl4Lm58QdzrDygXL5q5b+zwqlHds8LU
Yy0WeJzsPrADPReCh1vKX9U83aSmCRIvEMfv8LBMahT3hCk1hIndOPJVzKcXv3om
39XeMs2lk1WQjvaNlE95PSaFETg9L/bdcGV4x2ZCOu3BsiesiYSbMk7L9Y7Dw4rZ
fkfdziN4gYD+N6XA6pbtH7NA8N4XM3cQDT9vfwXSp4igVVNj1gYucxJEYuUlxPBJ
6EdAl7rMJcAtJ4kFMtK6rRskKpQcQLUlmDBgR74cSQdOspLCCR7Z3tCHJyu/I9FT
zLmE7SpwKloUEshRt89IrIsfpNFBrfV2RqCRmhxj+s/6P4+qegSeNj6Yzk+hQEOH
km0Y3+V/M7QM78hUD7TGJTP+puIWVjadPDV3FBV9ry7PIoZ7SPLiRGkSK0HwHD7M
mMGmRTBOGB1yDopBAz4hJIoV2HIRRQSKfo1HG1uD5MklODaNSaH/fgjzfdwP4Ve6
rdIm+GgqV36DII6Z4mdPtG0aLNS5W1MKBEyie6yQWJnw0vDZ65GUZ5u881yVNYe+
RV0L/c28a1aVy1can2p+lRMsssr8G0ltrfnNQUPx2ATwc8Z0GsN3bc6H7yWPMIxF
FNs83wV27ipiA/mczC4Gbo7kkMW1bjLN2+4AK6xzH3Kp/H4GRCUro50g3Z5fgNQ9
xWFtarVn9FTJ5j1MBJ5ODakcyNkwBmRxB3fY2yXbJ9BZOLEBBXCKg1RLiJMhWOtU
kvrgHiIRE6BhtBDshqx5KNljva9Sjb0AseV7bowIl0EDvVY5keQaNb2zEjJqqmui
6MxBH6G04/qpllrJ6anQu9iavKMl4+iicJrMROmm2OHSAayoMOKMVE6cqBeP0VSL
PQbOKGbWrpbFWLO34KchXMPmATwYOv4OwfkOuTBhZ+lh+7yYVtKf9aJgkamHTsZW
oh88f7U/H5jFF2KuivPVSKd7GYcPWTaKwAT0W5flaXi6E2M0ldedm31JjuhYbYio
4boxQcjHKLJnKCBRBVa/mrzrsBl7w7gc4B5UYplIF1P4O8kEcnl1JCd652y/qMUN
5nxYbPGY+iTzDSB6DmS4k5jMpRaySI27CGVyA4GRQqLFqzJuX6vRKXm0v4nUE8iT
nMLfa3G04fI9lw+vkqK6AVAQ/aE1fDVZFhmnRu80IqHmJy2PM9WWVJMjKYvL8eZI
efGDdMDA3QYP50kgVfm8jZhQiRG4sJ5JCkZAoCawJ4eGZmd+oc/K5Tnw3jI6tqi5
Bk75DyU6hfUIXCA1TTKOnFaGtaKl8NdgMNNtxI9qNAIjJSILSUKGTKxAnxWfhNuM
7C/Y7+HWCtrJHf7jSneMfG8F7orxIwoeNp9vI9DcZ5jBzmLs9ZdgJgBk1PLeFy4M
VpZU22aWnlCi9rgQytZrPdR8LOKmYjSeDzNS2CXnE8xqZA3rOAPsGEv3BKSaZSK6
b0NGoFpb2+t6WJfCBNneWOLHZI5ILID7pCAhoJUA3Py33g38uZFvy7Qata7BZxEZ
hJLOhqY/J7+0lRBMCTs4/HIOMMV2exvrxov/4BGCa9tX5P8o9SxBT1ZKMQxL+kdp
WGIPlL3OkzjW6rbbbREBdqwQpWfI+DiIwWsunn+pD14m5+x4cvI4US0/9ufdxZPs
gcy7s725aos+cQ/VAA8+fzhhxgV62K1YGsaKg0BOXLD3VAXV8XRCoXcUZ+6NpeLa
shwgQlcTl5qMBwMw/LOMTevlqifefxYId9WlTWd/HrXI8jqlVduY2Kgu2pC5cvy8
O1kT12LppctyoWG890pZTlW0QYmPp20U3dW2qTG3rt+nL3WlBV7Uqv5pvQ/p6TLx
BZK9S3hRT965s5hJylBir0sIglUaPwMp5MxoXqO1YgGJEe0P0G2zHXRWxuW6GTCI
rw7neRcx3kYwdRia+rrK8qncweMgbAdaZTnoYA9NeYRUOFiaxhqhb2E2gbTjN75s
yMx8KpOXQZOkjc/HomYAeccIMTTTytX0i3oDmxNtkvZVgvkQX/pae/5dRjLGy0Wk
nZaeCsJJi1cYi9hVh20wQm6O7i1R2/X3s2U2DkXdOjjwxM7qxtAR3HW5sGglslAi
zIxIPqM/MELyqm6I7WUpUC3xStqbldYFUFkeWi+OnSrw5xCfhtmdfGYq8MQQ5UVm
6EWBCMgA46xQuQ2hBXebVT43nJWezD2gEFHOE8/VFAfSgM1FqpamWVVP0JuEQZJH
Fem0/7gkV/RKbvCxPMmWwOF2mBreH1qYK82oCEQBK/H1oI3+PVjERPtRVITPrttm
5uVHz1PwIAGTe6fH+t4jTT0QMCYIPBsPLRUDBwBMf27kzo/4jJWAS7zQfFDDla2k
2r+55ZN1/vbOhG5talmFTTfYVOpx6o7QQPmiRbfKWRmxAh8vVTJVb3H3sl1xotiY
MAcsw5s8XmtF8bYlRV4pWSCYdgzOYolZR+1nAuzoaMQHj0q66Nbc7kGuvjJ6tQJz
TSaJn7RuffdDh7f045D0eVhX9zyCmYYAkRNVHjo4GH3I4hVKHk8sMS2k98OOWjHQ
JoVQDNTlnpDKyH3zSlwIViQAu9AVde09kJIS/HJh6SuwwLUoqExIMUSrVNyYaLqG
fCSSRYFfER/fv46v+VxQjW4Re7oUSnBtnHfJQnzRdNGfKzeu5/rAdBW+Iwz84Ndi
pebFhynHT/5R14wC+HpDb/YBqUpXZQCfyli+sKFI9laCNLMLCr9XfLP+BOu8zkJZ
7IT5naBJrYZQDutjl0Un7TNjCQCDZR2wAa9+a40Lw+t5FnJSFB5bP+obYrEx9rSA
PG0OB3sWbmo2MQ56AtsjjHiSPRMntVIbLDpwYUauRJi0754EE3Zu5h4b6RWHhMtF
9/rYILFEXZTypk8vrlNZ0J1sgdf3NfI4ksgL/G3MZBvG+ubOnLBPnkdujo0eASu/
Ft0BMLyOFEKMAH4wMdYzgbQScHPoE+klArzhhNV+NlqVNXfqCQuYJwhTfy003yKL
5mSC8ewC0fnlbJNOx4stNjIudPeTHTwGH5F7zw5uyBm6DCHWvjD25RIISBTQ1fY9
ER+9adt3EfnZNBwI8aXHBBazPKE/vJYnN/LZt3/oj9BcDoX66RAT6yKR9DA326pC
p/HJvJ4QbvgBDoVfdQpN8iKhLQUGsgEVOBLX6y5ygKVp0TgCvS8kg0UWvLgkxz3M
erhjOAAhKO3ANUl8nTjJqs6RxQ3N4WIOahDJ+2jQxj1VFyYJiSmi2V5wqtI594e5
vqgA3eXRvWjFKTtktIW+HhXRSEXGky9C47oG0Q0DGcfrSlB/3zdxqvRjtcREq7qO
TObrhGfv0mvn1mTkLgcHxPY2lKtRsBLgrsAKNHZL5xpFq/laOURhLZFjBNmdsLSm
gaUg55sizzDJ47B7nAX+KFABTyxK94KbUtFRIdnfEsUnVKp6qur6oGhmQT5iSCSc
G45L9/NljCxV4BR34ie0w2G1r95S3+gvKOnMKTTBJfdJD/hC24T0RWYCjS48SIi2
cTu0ElQUazb+7fxVoNZeLkP2E2mvFlBnjf/9ROmXWxw8MsRn4eiMcVlI4+hVeReC
fsCm+bgwJhtOsnxBHGuMKOARVIh/ZcV+/f079sO5euOWN+17muI+Gfp9ty9ofit6
dadZw5eqkpVrpHt8F7f0SiGBFLMTAdTIODMoF2cQOPZxibvxs7uoDlhwiqO2POwD
TT7Mv0bU38RT/bn0BrQZsq392JujogJsnESSKPzdD44DG8JzdyWlerP7O10oxafV
WgaAfmWagNltFnR10xc8hjDTzMl1YCEhewvfgZ4AsulsT6YkmhRwWKq+PTgYs5/K
nIbTQknvF6DAF6Lr7PFJIZJAl6965h0TDI8YLQwnCiOVJV/UW64BB9sYo0/KBW2w
S4C2XxHT9DFbucMkRRvkXmB2EyggRmq5LJyBs59Grrw/VE98BZEOOEg4NxGrLOwL
IinbkBCgkghcXdifi/a3HWVzi0k1WWw3+X5CIH0VtUFttro3PHmmQiueacu76usP
AW2mQQ8cc/fIyDjNeHK5q3AHX5QeiOBkNVzaM/DWY50ZU0s4pEB9fpt7jkbKopi9
LY3aECQTqKulF6uPXIdzZ3nIqZGfjPTIL4o9H/hD7bmWJJuONZSOQv5690BIFyS0
AVLF+IDwAqDUqNteJdxfrm9IYAipgrZeh6K3lwO8bnGd3n5oDsSiYxFjo9r+zEA/
u68t4i1RVTIRy+boVil5+hG/f/23G4BIqh5yKoc7Q7Hvu239x9PQ74uQhsJyn9S4
Ydc3m1XATYeduNS2vtTIeOWrsk9ojyDw3h3u2+3wpxY8aXiHo2ac+HLNsxZiB9Rz
ANwYl5FqccMLGvq+wFTZrM39auI/lNHiFpf5sY/+jazlooih7/hkE2h2yMLQF7wK
JOKgzviINJsF60yBA9HdHTZoZk1rBGIRBPJHAL0vp59TzQVj/zCmDZW+JBRvpwbx
nL08Sgduknq7MSTnhugI7rr895Puu6IYR4ZsdUIHu42khwUI0dw3HjDjsZbyPrGC
Y8mL6/wC9WVIe9tzpaTb+Fcr4vHwtjC0mZDTP98onCA6zyQrxSzb7Z1qqIWtVrQB
sPTlPGaYbmbDPFb2WdIKsS2idsqYkUaX5erUW/axz9u0lEXEWYvKyktNXSv8R1QB
/UOLfvxZQZR8GHzGDpThEMf1xg8WM4L8usLsoOu2lwH9+L1oJKvp9W6zrxeWucIm
SvOePsKonSTHyvAI322ta/DYo+rODwjbhBuF02MW9lOWKltt5ZOkKJiG60BqaIAe
8PeBY4XLNVkPRaTpKum0PBiJP45CSJCxW1BJxfim2r8TkTcDkmb3j2BjwyaodcN5
51Jo+hEo+OnBAMqyg8zQfAQqco2hu1H/PbcpFwQkRoP48p6BGNX/ukPP7EoFkB43
tHv5Stx6GVTylKQ9RNQ0j0v+iKpVyS2JJMrcc1R7AVC3mH9dWJAxtKHnPbiLTRCJ
AnBJDDYggFaVnBT2b3DCZ0KgpRI6YjwuPCNQ512ZZULDTgxTcyK+CTbsY044mJ+R
fWUO771JnpWUGMqz1FkT8LieD+xCUXbx49X8mgrjcztosrVGDVQkk9ePENgKWZQT
I0IwvM79nlUp7a8zQgybR7Z6Tx3v5mlsCnNjt729e3Men7lBmxocIQnQ9/+iYXVZ
8h6jcfe8isy5k8VdOWwanT7rjuZRdxkw6RxeI4gDiqXhkcAXVF81dil//z8EnYwN
TS9Fx/kzW/ZI+Uus3BrWqXdqbeL8QxZ3+lXl/ZSWWx2G3p4pKR9p6IFjfwPAkgj3
eNwW4ZvJIk9PVhqbqmfUhd4gZqN8r9gAnAhUPtjRO8Ubcsqp8KBCj/mxNCThX9u4
ztM9JwQRbBj7nH1KcksEKSJoD/aeaB3d1EOiNSjb5vg6QLBOhRMyXU0+JAWDoW32
0lXvPb6psdQniidwuD+oq2PIsc2gxAB84P8b/v+A8TgDTXfoVCptmaV5UFrqK20d
8A2D3jw776vwgFx38iasm8CcCYSO8AWfp6J/SB6EK44thMu36+y4Cz7+MrkNPbBx
3DHMiAKMh02+EIzZIuqwF1IAVMPxJNYb2dqBWWRPeZySwiZOPmuGbNB15urwsRru
/bDVTS/aqsSluHqbRtc5ulBQZ5C5zU2mGchbk5dBK8ojDZem+I3HwUteu5L9FQJP
NpcMfCbgWW+8z+Yy8Ghz7zeTNeevlLsBgmxugVafu/lYXNBU+sNHNeBy3dyU3CIB
LdQfgsvDw/4eLmPOEQ3t4CEfiEn1RMNf1gXXDqE3vzJBTPaFAA1eWRUrFnRaysz0
9p/bkdoTnVHYtEL+AD8oFkU84XIcT1/HtlpXfII/JUteM2S5+p0gWcC5jCRGTpTc
DmgUlMVxn1OCzOcdRJXtMZ1UOI/a4EsvpWHkoB7vlEYAXLzDQpaCtDG5XqcyE7aL
2JML6TpX7V70TP/WLCL4FXTQZCy7IBg69SjWdVhngtFcfMRAgBxcW9HKgf0KV5dl
/LfCbzqh0UYZpPoAtPZQ140sY3L8c0en1c4TVQlzyuTp4l8zbCMdYkk9xDL6/M1P
Obg+30yVKUyv1RSvgiZZZe5ycnjc35AXCkFDTfpXkvfcGCjdnLWk5/ebk96AKiuw
w86wi1UR07wyWC0dwA9wI5uWHG5/zYam3oj2eGg62hd1tLSDCyxSQ52HxaAw5j9K
t4zSvlgVHA8eH49t4wBwiIwrfU5fa5DA2lRsbPdTX3h5C5x2YGCMPAO6i+DPcf2X
vIbZY1wpOaDjFYZEbsA1fKjCh0/v468bAgqIZ8kyfUnP9tFEHn+FCYcxZIUH2LvI
iZ1dLAptVpWwUkaRSPQin1xjX5gSpZGWfNggCJC4C+4noFT72PjEXlTJdusy/HdW
JW1t5hbFgNFkFE+2SsaYt2ojyedKmZF7re76FNFJSHqUE/JuI0XDuGpoXgT7vat5
d7bXbVikH3w+/eh/7EDKCw2oBg7IKrhGW/xl0YHp3N9N5zVgGvvCm/MNUN4VGYJ3
QMNACEc5sFS1JXZ2CWPitZ008Pm1xNC1jMRScRSVPlvqOCL74/XzJ0sPYOcakME5
u1TUaOATEsAj5aBBtJVKBis0EVCLSCYyoTCKEFTqgvMm4uiVJ8L+LFERyjH4KXQg
a5k9iCbnrlEMrHa+XLqvXn1jA0UYHoktTZjD/vuG1k5OdxIfiZjmlqNUXswUybSu
eScF7gTJXP+Ckx70LWIOilc7c4hKdAsswI1oNRnesV5IZqbv5t8/EFkh8RzcHc7e
gsvKVzCSmdAkTQaHBfLtyjl50iIiaYxICHwa3BJEUJhBlr7CD/S/F+rZXxigILCM
T3LG4itZ2EYeuAjNa+6Wcbx+vs2aOUP95D9KaF7rFuLMIR3wU0zzJ1hw30Um+nr2
0rZcgyy22IACdVZTq0IsMcEtnTej7s1udjVRNo1ZX8RiWvS3TkJFtrvLIp90+peS
n13dCr9D3Z8NFR1lkZ1PRcCG5D69Q+MtV2785e4mSU2U4wNBE1KqXyvJxmSQ8PB/
vy/+yTzNBl47i7Quy79KLdAlLAFKDOBJ5ZnKNn/HAXqdSiarTi8Z8zQGwfZPhMOL
+TxU2oYImIs14txKE0NfODFneo+94YTivvGL0yVqsvTMcbNeEueyOr9wjpu9AZ7V
4aq4iyU+Mv2aZdq6gNff3bi1aiCL7docdtti2cD9Q6FhMao/S/FZ0Z/MW0hycQ95
O68a4hO1yNXFPQTLwyNCwWv536eHbzxc8CNGQ1a5Ptu/DuOWizG9ofuWUndiWUJQ
wFwikR6GeX+ZKL7Q03232yd7NpZm90p0TKexzTQlw0nK0hw18mYJ1Cpr0lsaFSOA
g3ARghLo13r1xoRD2S+tQ7ZuAwbaiRVqshVLUaQF4qW3uH4OfYkIYB5T234T0of7
2l6Jx4lIA86E+2fNmQcYA0JClCdI0CaP4Vw2VUcjHNBUnWBMM+zicWbPVAIUTeG+
zPWLP0Pg75XGJJV+UShY409aW7bXANzLiWABno9+mSNx+zHbk217BzrXwk6FpXvs
7AxRTtcHQU1JoDGVu4K2qI4c6Uw6Hbjdjy+LJ8YzqbsRc+ES6fQe385Ay4USm7ux
ui5a7Hq/oROzdwK54kkgLayhsAY+i0aUBiyMsugH4zaWYp1O6N2q+hWvOYaUqbER
32dz2mmncuv8m8nydi0T3wfrINJ+rz7W4jagn0zw7cBuB9Ma4m2C/+deUz4ltENl
hGtFpxJk4GCeLwANp1hmUHhbQe9tL2BkYVvehwhCkXrHfrtSZmtTj7+1VapMA50G
Lp6o8+pk3UaXrqeK/5rLEEPIXIZw1nhlsy58J0gaM+gscvtMofxfqa4uFKo36bpS
GtLIm1ziwqg73wOe3/nuEB5zx/CzXcAXiXyihXPIvJVbun7FxF7cziJF1ZlrkD/j
DnT0Tb9Mqhn7kWR/cCSJV2hDzT5WnOlwHmFxQCanPa16SHZYoIXbLDp1+T6MBa4x
rd6nxTtajkjStzaK5mkyaYROQiO0/eXry7BfpYvjHfiCHdRqFr3pX8sP1TWr/rbm
OVx4LL7U+OOsVM+hJpERymJO+a7Gkm0rVb4HR9SyrzvXrnPzhKJmSkdxXOgwKn3/
1cmWp4giTUQWUY4uePaRg1xwE7ys0o1RLvkiNwMo+NkCxPrKXJZo0RjLIkcHgHrD
MoK1vp/BBO8luIhafhZvCFB7RUz0sOJTMmoz/JCma0K74lMHMk/nstkxZ4oKKO1r
VHP6BInQHHPNjXkLWesOCcMPmtNXcsKVVBUsHXpEim+y+UDUe/okaB/Je65IHpnO
28EYa/XbGua7HLxjJKa5s5dOJ8a+NBbyPiaXr6T3BCLopEMqSPyw5D0ksVHaove3
Eg5mdAeqlM/JQCEqK4Izjj5bLTr9nep5ZTH2kF6bjYRmEjg92N+Z6dzisqsSJ0jh
PdDVtBioKucDred61w+XbdqxQi1doOll2n40TpF0G5pMOHAKR/71/6ef1fXWR5JN
KXGXMQROgFzqKdlFRayn3CY7ukakVdfxfElQK9L2ibqyRVJhbl+LhgFU/MhZJypE
XM/UrEM8nSqNk2+9sJKkvrNrsqIApXy/Z83fvQLWn2BLoltsQWl6bRmyWYN0NCvY
MYMuqQHad6Bqp25WltCQ9YHHi5oZ6xKXHRLNa3wQRc8Xpf5QdFEBs2gNAPymgAvj
NIymrNyX06r4X14PJvE/fJuv5halJk6/Fmk5sQbcyn1GnUzwBT54arYAwF1d4uDC
ZaOVlsLA2NZQ8j0hTBFJy8BKfCvg++p2aS1mhSkeRKfWj+S7wdniu90SfhKcBpZn
OpVfZV8PwMiStm4SjR4lIuWc9UKwo115R0eyvnHOy6xahcbXiBhTKKM4JeaAcoEX
y/0+nX0WCG1uMeNHRV5wmptsu1Ql7wG+EMdJsg/Hc5QfhS/dNcJWkWwQNRogA5hw
7KQCqLjVko/ombSGNBLBiDvjyJsa/0KJJiTgkKj7V2W2Te677MnABi4nxzodRM0j
sQcvN9xKUm9hnfNk6VIPutqiCHScX+j9DlY0ygqw47XINnXaNwnDEJnUkS5H/Wkx
udLlkGj7/QMFkz3RspwvP+fEugJiZcTi1YM2+M0Me1cfW4dgaNekRCI7kXB2bylb
GAfT9AQO7SNpzXrBh/s8IhWnhVxfnMZ0L/UAPJraQanK7dmS4a9kiWRYpklqy+fl
wFoULr7ZOSk45qVYf1on/O9DM6tXCNIs5v4tClGQbzq+y/EZkrx8bho1gY+Jcpn3
ePym5xORq1eY4pL8bOA4Su2hIDXyrFFcREkXP6lwSJ/Uusr50Q7Qe3I+U5gSP0QI
kutv4Sje+WR4mov0/DHODGxwDN8xidDI9JEa4Rxb+F89MNtgfmRgLl5pp7aKnJBI
GWlfIhTok/0PNqDZspxor2Hdo7sXwEChdCAl7Tct3yEXclS0kHmqcaIleqMPseEY
wOiRLXE3wbk/e5+vQrS7CUoDDfkqTnjA1s7YkdqD2nTcB0S+LjtWbhoJxc4Lbz14
rRs2eOW1HCc8YZOqoLh64ovAfrtFdorgI79Z1cM6BOHbc4lXhJQa8xmFFWTQyJ89
zpkRSF0K9GJrmiEujJhsS6gA8xS79OlfvmvhGA72J8mA2w0WGd0i1kAWB/yoJZhg
UdyeVezpgTl687Xclgisnsai3+YKzl2dDLCKaR6RqRgKXWT7Zs5Kt0hOqOFhy8R6
4E7+6TBk3vQyk+Iu9XZhY45HlYekCeRzj879JppObKiQs1tlDuzDWfj6KUcvJ2jh
KYm85/u8q11sPsSOA7PexvqpkkIoRYtVcxir6gbRdi4mkrWefLHXKNRFZJZzDmHh
eX0lUe09/LuvsZ0O3Es2rUVnJMMY5eZbzKtD+cjIVO67vM0R+YHcvA05xRGiSI6J
aRpbGwj8uXtLMGSKGEb8/pCSNnrdivCTKvfmo/K2TguACd9cY/wvTbQ3hIIIM5Pf
2W0nssDX4WpuIWiTSbu2VulqxQFHb/ARJRtTpg4uMx6Gtdj4EqcnD6JkzcygwVIg
pSAtfu9i+C/XcvsZTC2qfp3tg1bJ3m7H/7w5p/86TdCzjjPL2fTRqzP3RR5/Fzw8
lRaZvsITG9FZkV6AoVTQpOdzRSeMn0lwI4PdqU6DgwJ4o9z+HeKacTW1K2rB9JZl
HuMcNtQaED9M7V3/sN4eYQWUsl4fwxo26kY3GkBEMOT8oYZa+CpJfwgSCYtxCs5L
z7BKKvJ7dzNBQww1EqRkAhXDKSku41hSKWZEhNpHDJ5D2MJEpuqLntHVs8RC5DBj
G2/foD4l6L77eU8hD5hRG3ki2t2euoiCh3gs7WebPmM9/ZC7Y909ICFVtNC4bDOv
VvYUU3JBW6kAXRgmiIFC3VPl1sKdTwMY/8dIVjMseRMOD2hvH3P4K9G/8KG+ZnD+
VwKvBSN/lJGzNGoi/3D9OsLXBUQR7IIuW/wIfw182OVWMh0vUuVNj4ymxXSmqTlq
eYVlXnfudeR0PHStL3SactXW7q5za8OaoHYIt6hVRkg+sZ/+Q1JnAb14dHqHkrJO
8AHk+u3zGkFtrEV3mhDPkDi0IYh3gynfHjBGB8laqOiuihxIQHbadb/mBFT1qhxG
gxWtQcs7F/RT0d1F7CeVbODmDZvH02PKDjUFbhUikYPEccLHDt2gyI/yVKQrMhwp
SKlxkwjyVbZBPHLLxzAjoiXsiw6lR80Cmcz8u4eWzERZuS5M4e3wgFpYTQZxdnS8
2NFJyqqdTP4W+6G1fBWWgNP55xIAXU94e91XC6DhIIjWwhMQZWBqSIJunmhutMrE
OHEh/7/3M8jofaxgTimIxCG4I68EjIm9ik3qhucvSha4iUmSGaxJ/ku5mIIuvbaK
MFOCj+R+pp8ReqYWYsmBU2CAj0f0rY8rsH5kTD01QjL9WhT/bet9fFvcsuZnFdto
zA5ArBIQcnc1gbflQsxHZeRTGA5JsSAF9IMo3vGvD86BKHsLkLMaW+cL015QJ/c4
/Tvax3hjDLnjCLkUeXehhuh0TUkboV+C+qp4h/McWDvOP9PiSRimgGDzRrSo5d24
Q9BmE9kmjmN8rbQnRjEeUPpUIaEkoW9DXkHtdadXBKUzL/Y2K20aSWu2Z1ItzUPU
TtrAyyWozZPp5sDY2+kI43j701L6+Jp7U3v45naO+0/2T1EJwLVv5yrDDaO9+Vp3
N1NqsBNW11rdOxBPmcBXmo2oPEEPGZqsl4L7boX6SduyeKz+9QoY3u8dfqslMd4L
rEtLmhjH8+DcO5LjOZjHe96jnjKQPBJiTz5fUITWdqJfmYrxvI7n1akp1dk6nTEr
8Ph9uaRs0hHn/vWeji1wF6sLYAzijJajpiS4r+Ivy0rHfvBK6hhtQdCCF6gjZwcl
QCidzJUB2YBA/pbPIkOYURnrabI06L9LYYWsJLzic1AxGx8P7WXgI9z6ebAUAItg
GmLIlN/jUe0LmQLPL6A/ZcMH95R6Jc+R3rwdC+Ar9yl2FtEjkKQUR0Y5K7Zxyxah
bRewDwcD6D3c9icaiguBvqyZ4iTN6gQ7VhhYEI87u/oIXQwKRqdQpixkTYQDKRA7
93LHW/JWQCylgcOjqSa2DJVga3ako0n13h1QC0wD5cr0gYlv52hoIvGchpIr79Og
HWzGZDmJ+1EBEAkHJp0J7OKCKwfzWlEdiDd8qSG1hGsBD7vuZK8Anp1/kdGkePOV
+dB6eAJnoYQvwvAx6CXQfSjbqXb2XAu1wHXK8wACpkcedcPb7rkwXBfZszf3rWM0
CJahswHfo1s6rVwlxNAjsBg8Nuf7SEstqDO77wdZkpO+Wkvr4c8HLuIC8FJEbpdM
IU4xOefC6D6ir7t7vebKYGCWqijHxU/77rT9j6xBBgHFDZmV5vz+QYCOlsSllvy6
eY1COYVn5QR4jhsMHq354lWTTLS0Byi3NtTpTBsAKIQEOgVpgduZgcYn1TVwqrox
yjq/exIyFBb2MBxDZHWOv529xOlsTyEKjFP8IU1gHfQ6LhxHIVYhyuTmDEAXqhEs
VsnHUEuommAVLTdZ9AfXTKOIFg+4OIFUfskcTk+bGJdI33hlDeWQNfsw/rtcXfcP
S/XBs3mzb8Sk+AaJgdkl9ownnpdDrlwyoTtUVuy6WKTpQ9AWofSPAarogFTkKrUI
AfF32XZ8RFmT4iA3wgv/Ik57N7BngCx1/vG3WvJaA+UUkz/ON2NoCLsJKFbgQXQt
tq4NxBmL4pURJMEfZPrND56il+oxWIZdfVNphpzgVGTj7hTMHaLF5yvhUT0aBKhw
QZLnnRXaFsDH8NAbkbC3rcUHUpnwVoYamYJ5o+5oWQo7TkmPemaNFtFm/AR5dBFx
fubytlsa21y0P8CJRohikeCzBLiBABIaah+AN3HXqhJ+AdCkuj+yZkVFmDQOJCp7
6hz3RaMvJBDzCEHPBLKwiOCHSYnbYhy6BPWdiBGfOxNgXiPa60/lZI5yE7DAqWmy
wEMHFyMLnfpOCsqvv7/YI9x+vUET+cyTFmWbScxDRw4UcTWHtKuVhRJdqET6LqJN
P+T0Zm/WuGa3Av9qFVKKs8/vSt2NivZbIzpXROpWV9pvXJOd8o9Sp/EKGDBKBjcA
YyuKcAjeNWSyh0set5dB9JWpen/Bm8Ao5RcKqIq4XWLvZ8X0v1MrMoTYOC7A+H0i
JZfSQ/vgJY+Ve13uLHthJJ6WGziMkhcBxFiJh1VcgJc1WtROnzH4fOHTE9ZBaQ+d
xJZT85h2FiJGL2CsXocefNXUHvaVcMd4Id0TNQEGaa9Rc/t4zgvbP5W31+qanTKJ
wuRSMI7exk6MDwZYjSpJV4y96FQisG8/yk5bw3poFsf36iiqybBpj/Vancsj0kmh
Gb6IoKM55JXCqYD2TF9yF1bvAgjMXIFT9q00Z2nLZhkyjzcVoqNNOGCYEFWf+gXl
cPGIPmjhDCjVSkpoId8GZViFSGMi5WbrdJgSKjWYZLiHtNGERUG9uk2SMQtx6f7a
GGdWQpEOqgyQrqQO8u6HUyH2zJpCflBrxb+cLu8ykXWBid3JLbFocEntT4JsC+ZD
bYNl4p9eaYxf8mDgbMJT/h8x2I/8/fg+nOxFk6a6UI0r3fnFs5o9JOSI/yxdgzsm
y6SZPrAC4sQcZVmAUFylbrtB5z2dYQdLiFna0BeSgBcMkIFUhimIoP+qnj7ruhyP
aNrimeNMeAneiOrk4IMEVyNk7hdzeK3IKx9WBgHg8ZVZ9Bi93tE5qtEXd2qPF9zK
lOaChY5oPHHdFnDM+s/FRLOrs/M/tOlct5J0+XX0D5Cp8ECAM/THRdqge7OmNzQg
Muw2OQVV8BlXqdDfDk0qV4zH0D0wkfoQ/HodQwK40UN4LArDeHWa2LRCCtjL6k0Y
6s8zyShmiMQjXi3OP42P1vxWOuh7h50/kNZfWJHiv0/XCPnIQHnJK2hBIiOctHYi
szj93D6Qkd7qDNBDhpFKoxw0Y+eZWdc3FgUGeG7G9qkQHfqx//RANX4hc+68ab6X
PqMBwTKrMZbJP59FpKviF1nSyIBB9FUG+lbsxhfGZ1TVMayU9IMs45fHMz0lX2qY
kYVU9ZN9t8cDJ04Pw7fdQ2sZtZ7qJn8h+tU/7bnayLefyV/6g3Gzlbl1cWb10wn5
3xB/3rnIIuyu64Xe78Ki41gpubYW7Rm+3gA9wGgsnhB0VCZ7JtBxC/bXFwHIU9lo
iTufaS8rRMZjjkn8I2CHr8kjmigYRmkcDM7NnksZ9LRHmkFV7U775WVvV3HeLrii
efPJMntcPDIsr2SuzbPgmki5RO8qm1FUJXBNgy73w2lLRVHuMM011/rflTeC+q3I
msshGoO3n2YarCMxpbCDhYpg9kuX8srVMyoDevVR2zpXbim/FyF1N47v7qK+DRSa
xk18to65HztUK0/+ZaiILh4gJQZUXQjhf+EEZcJYFlD6E/BiEG6U2FvCpoUv1zAa
4r8zhIlgr4K+q8hh/gHKSsnZeqX9QRh4FlY/Fla8/+yqxPo85karFicq9DcsCXVM
IN4tRhT6JuLsRAx5O6fEpD3A2PScFg9FPkaQtQ5lsHWfssWsrMe9rDsM+wS9wZng
BVtf2ugA+LSUjtFRavNcDeLHSrxB/oCyh0OFD1++lFC7tgW21mHJMfumgNjKEnOo
lCmdojCSklWrvcFJd/Y1Vkc7DEWg+FNJPl+8jGLWysD6THmhPLeiqg5aJyu3MLR4
dda+STNoNBTyBgX17cWg4dwWrKB5YZ858ods8OBSnBLOOkX7iW5bOnFWcy4nF/Uy
6TH86souyuvUnNwBhdeEKkwlCXdtzBlZHEz+Fk0LyFsyssyRKsPQoaNyo9NdAnF/
Z0+KVozx5VGSrze/5tXD/1cybperYnmfaQkBQHewjGNk6Jv62khJDTcMRKHGHouF
cNhbSkFv6PZzMsYrT1Mt2Gwvh1nvRlRH52czQ6nvDdOY5W++KmdzQ7wXWoRhXEkP
RbxNQKFgtDgj8ckRoqqGL94MD+0gMl6b3aOoH2RWons365AwRsEyr8d/C8YRoyIG
EBD71pA6VmsAJqZpC/0HYgBVY4DDupY/nRTiqGbWFjnknHctGbyDHrk7bLQufk6d
kn1XU6bQYG/0eH8Kdf3a4PLAQB3AUM+0Uix2vLeNtADF3S/Ph+HERrVy3618HEDk
R5idBHAxkFPqzUSg/YO9TKphPWfDu7xZcwRye09ySGktiZmuZZuyLQYg9UmzpkGS
KAuMiEQ85WjZIHHDsYZPpmNLnLBoqhbP4jqKqHkW7rwmK0x3/Li20BnsYnqafant
bbpeOA5HbJBx3NwldXFv5R/z8OSYmWa08PbWRTP7uNDh2ZsS4AyOgqUwubFjFjgX
sqq7jO6ox8DEkzbpVDxHO7QHE92sgc0tczRQTqbdmihLtPZEVbKEhdFcB9Z2WK6K
Og6voC+PAhiIZCWHwx+Sx6BoOgKsei2dzw6b4R6IgAfmocQI6+a8CY+zZN7R0ybt
MGI9eh+KHFNT9r2tZIsc1dZHpAUnHt8Esu3iA6TF6BUq2Yn0uZDYXRYpbKHYRFML
EYhOoYo+L6FTsRvqUd37Hcc0qIo9G9Yv4uZ+ZJddQ2CyVDJIrHEjkNQkudktabC9
+YYUQokvSLaJP5c6JCSQVwFKbLCu81dRkqYaZIOfbujYJ1cLj41qWL8DQAaJxvUf
JpdfmtPai/3Iup1I110ILBFSD8Y57jPtkssJzJ8vKwTMiIyBCzl2eiD958HbFM2K
JfvIVTOdlaLmMkjyJ+WWJJffdlzrt+8djx/yz3ySFL36/N01W4TJhjQk33LnauPL
6EtGK1xckC04VvqiCITkMJPxeOcZ1M2SdB5780SOPHYEIGVFSwWcNImeBGDndssK
Tib75n3PBHfKkcYHrt2JjukQweg1I8tD0CpVriW8fWOStYG3qX8anYXWQgqRiPFx
nRT8AfgfUM60BVdNLWyeLN4in7I5bdaCErWC85k3D3xgHbL9MB3US043fLdGC4y8
RfNQtDtsEpwF3zj9SKPWwn/W1gC07fVX+Bmecef5XDa0LCsQV2+Ba3bQizLP1iab
aioWd4VPvRoZvU19R2UmUx1ThicSUdPHJ9xAmJ1/TQ4kjYj9hiOEMA4O6QMZxYOI
WrMK3iutFwRjT/KQdhqU4ZCKJb/lpNflwONpawm5WD8GgRibck7qO7ofkmiaCrnj
hzeR1NIqx8aF5If1tgOGhGdJVfUIbDH5U7vkP0ej7fjvqyohrMaBl4hXVwtEm7OL
bh0bqRevW2hgDvAcUj8ojny8OwmJjZxnGJohbSQBa6EgTnQHREJUCytdo0KQbIK8
fNT0UkdYypr4VGAImsEXx2V1NJTEG+xPreH6xV7iuVrzAqiogxyOT2msw5k4cS3h
O+nX5+1+W3WBYbdQ9QcKXemRjRyTjdHVloO5aOJt8sq2wZS1y46+auMsgaAwR4UZ
BgGZwcUJGbRqGdtc+t9QkXL0rLGFMC+P4r4sxthpTaN0e8VuEsNWXk40ikhgdaCL
hSu6jRn4cn+AbcVWV+9kg3J35lvxg4Vehg5PWIFf1Qd4afrCrCpCS4NxSA4U4/n9
/7scraCkAmYl+Y5gO7IUUIbNLj82nJTw+f9/1mJy22mFdcpw639f6UJr4i0tcOgu
N+sY0u+ekDxEtCssJoXh0CtqNCaT6iRQKtxQwRhZrjlVXt3l0x9gpfwGcomKJFUr
DmI2kV3qam+jx1mEG0D6Tnigg5xowc8VabAC3RBaLAmDaVKOZPKCaREO93XFNgoi
TZY7fZwZPdoEI0ExKfa6cvMQ80tk7m/B55GOgKEvoiTz6+4n0R58dR8uApz3rWKL
r334WYtgIad9lEWWDSkx+gCjiBsQui6gZ90+jDBn6hWZIOVp7nzFyQiqpD1hZw7v
VpsxnJtwaNIfpv+B9vrAGt9iWyDGChYNGGdXfMCxwCeX1yvHlkok8enIr6dVy/3D
c0WTvNU06QoTrp9yWLil7cXV2cfqiJHNYuIppfRyrziBaoratcQIiWNCzpR5jp1+
df0IotRbpaublpGatHwYsqN3Tw8687jknsIZc9XVlrWAGIvZwO4ofM2NCbFT9jW8
4yp26TfHJ3fNtyzaBfm+aGRE9DiyvLfznGtYCoFWhQrKbuDtATz13XvaPMWin1K6
IjfdDFAM6DS3fT71ifo+/NJmlV+iN6rDSiEdhNxlY5q42efKl163kl77iIWcznz3
3qT+pctQASt3tzW5ozLtCPe8EHHAiScwVr9ayc62Qd/lROnthMyxjWHlCXoNJJXC
7L0F9qhP4dvsR7/4CGi/CfnaloHknm09GONZGsin88SJD1gw6gt1E3NR0avKoj/g
ljehvbQ/OdRjxrCyu1dGIwb18Cd3aDs07o+AajVytfA57TF35X2JcUvU+vBT9OuS
JpZWQ5Fi715iahpvF5ljoZ47jH07ArepjZTZwg9Vl4yCniWj4Med4cIHV0Ej+45v
mYtqUxJkudPYDhL0eF5mfJs1P0yjaXLGjHVFrGBVoKe0K78fbhmqWBOjYM1NEHbR
wF75THV+fpzD5d4F2U4VLC45h1/Tt6EGTXYL0OM2xdyaa/rQodkxeWjDyJXeqcBB
mqtEI5JUZKHtggreRg55glQXbYi8hC5n78R7B5S2iYVFxRfbvzVO9lKn2rZB7sqy
wMrgWs0hXl0dDZj+IUrjeSdZOGbHV8PxjkfWmFpLLX1VEudPurg7XENOXSadOzXf
m5Mak4tuO9jkUvl5dQj7dJQvJ+/EZtbAPZwL+w1/2Z2r+5UkmO6k6XqcK9foa2TZ
yN3SOR5jtUpDooDOLwD0tW7W6vCVQS2KSPrUVb7d98ZoIeUUyAUaxL7HNYpDYwFc
P+hK0qW0VzkdUeLmfMHfNaqQW8XJGfPdPV/HCSzqX7hRD3aLqvcyRF2BgZrY1Qct
KmJb4JxAOCKdTZto0oNVh+sCAiLY3uqT7CNzoOo9jIHigbHJVUHaldR8ng2c/GI/
ynLiwnd0emaxwzvSfwpk6nCk61HT10djiOx/LzkgzUsisNuOmVMLA8FfTypAK05J
LDDqWmePjrVnJbGQSFBLNwVn4GUreX/M2mjv7kJI1VyYSigNxM8Xiy4g3VBefSDd
KCMHIAv4hfypuntaeahplA9RfclMy2QikPgKHG1RQn5dCyfVYZ7FIc2uVlNNeV+y
KFrM2f6AqjwNaF0REK3U8rn7OSiDkSR6HCvfR1NjvJbQrQJFNmC/Y/VewzAmYfcU
tS+ZbcyBHs80jESUkwMu50LpjgGU4CKs7hJ8kvQ3V0DVKXhFDSvOk2VtcCpc450d
HbjeKfqT4Phw10QPxW8fhkMR1pxDyPRNmwHoXi+COP9razZgRMJ++gRHfJof9tdE
RgvIzKQNiszK4mBzQjpJ/vkI8caPaTe/7wm0UYl8rARgRjUNlgXNb1ei4KR8BSAd
JtkU9FQT27h5WFtqYqaNsYXFhzPgSYysyuOLkms44leBobIxnU3jg6ppEG8ThigJ
XLgzNWRCumsNpr/3lmqphXinyce2QXSii5cTdIxFyb6ATuLIFUU9fK8Nwc0D61mg
OFn/iZn/Hjw5jBbrmLypL50gM1WdOsIpYJTbDulhYxOR/jv/GGOG2jIXslCZiHWb
OwqVS/WTlFSwGZyZLaEHrpPi/lU/41mtdlyYBsvTAp70R4Q2JMTtvU+bGaaRZ6Ra
iUiL3n15Lfhdn4+fbmE6acgk+bT5n19IuFPyg+m51vSBsEsXAOUN8yZjPpiGNEpg
xtA1I+NwUhgxcvYyy0husef0etEZNw7qtVAWzS+K9jbo0lXL9clAND4GtssOQAXS
1KY9Gp5m4W1u1n//W4YUMtSDYpEStG9+KLjD0bK2WZLVs0MNgefDm+5YVCsWpQ9p
gXTyx8cp+DsjqIKJicnEWRjRM3y4We65S9/I3QAxzJNKnsvMwQwO7AHogeSyqatB
4zhoAUQ+qi6Lecpnest6qIJLbvnWhe9plfRE634w/QwPgw+GsSvtB3eXZalk6Qrk
mSudYWTb9/PzfFLZ/ZArp1s1aCw9qmwjIw+4JTi5+Sd8ilhp3jCYQnmIY4H4utoZ
q9T5RrRuMU1DxRpaqTb4t8oPch/Z+mYSPE1nEbDATrah37LzfIHQiLWS8V6hRSiu
ZcdNnmyins/XUKeM5z4pghk0HHTSSTJy3OKaj0oFeM+zsQG6TxSXI4uCJ6yFeFAn
9rMCQbotgjkyqgvjTKdA1yKZlwiFcm9dceEr3UcT89owySatiyIpY2B/lIlNNb/T
dGlhpcznLyxh+9FWrs8w97Sb61/1KwpwWEMTrzWJsfEKr9OhkRFwp5EUEl2/IEbh
7JCA5V1Hga8lObCudFpEoE3nH4rOGVyzA0Z7wMD8XmqhH2wfhJcd/VruxpguE3TI
bYxvnU/kw8F9qn9cn39UT9cjjWhytlxGzRCPJZbOBfdYBXNBQ9WAR37K7R4z2Gco
r5bZCaJd/vn5KVPNPFxAv3jEzwo1VrEAuQEmnum/AtpuGmfgVJ+wFKcIO/ooOusA
3lPmzcXYjk8OznTdO0aVaNpLBwgVLeQSGvZh5cOkpXcxOJ3ggIlacMfrm4qOL161
XwUfsmOWNlXOGLqdl+2bZRi3IDCxKHOHDiVey+ANS+Gb7yIpMsyWQAq/R5ePKowZ
kHAK0lMm0o+lIoYulirr4a3YM6WVDna3wz24+yELYRRxCHZODFhxqMFE2SblwGHj
8QztrbSoJtgDBURLUcYUjmBq8Q9GjV85+wlqaLEht8vUdApKc6fBAm/pNLx5xkKP
FDycXXWgVEBYSYD1/WkktAROhD+ttErEseMAv6zCTeq681TNQ3Ot/C+lmk65tQih
JlhAoKkwzAK7DlGXECDY6lAhsnwpA7Un9V13y5ur1O0CQK9Mm2YWkCtu2nWO4Hk+
/KSDoikfiSgiS8co7v9e5AJVJ4OjTKsz82tYqvBKpn0scSjN6oVjQ7pLHW3Z/Ik4
9lp70OBRyna866/tKht+kfW5o55/8a6lv+ePnkrrQA2SFqlPi95OkENX7P/yVoW6
fIfW7uUCkR6Be7kLItJlHGhxQyxMBFSboFNsR09iQQZWHXaLVmyKpjZuhtXlP/zA
M5qyMoqCI8yMJbFCW4ijRJ+r4BsqvPNnLGxSMaa6prmQCCywSxKS1xmumu+iobcA
dCubfuJ/+o2sYG4LdZ2JAoiPQIlndz63WnfIWt3vAErJ6niQM1t6GBoN+QtQ8uOP
aEmhzMPRVCbPFDirNMXMFf63hliPpNcDgnAqLIR9graT1LQ7FUvqYMN+X/sXwEJp
7CaynNwfVL6w8wnXnznEtFAH/kaaY8Gg5FThFNt8FuW+N5IoPM98OyVooVWfWGoh
vxkvPQivjFzIxk1v122JfqhBxhCdY2Xa/h73beI3RM1xaQLHFXEGSOxqlrvidUje
ipTLWam7ihGnMvataV3wbswVgQxxvLueaZCYCq11x4uJvOmDgOB329R32QzT4bRd
LHwS8ZV5IkckEYW//Ar5S2BDUZsHkrJK3xCPk/4Qi9R0vgOiFnKJfD1tv3s2l/Ko
znoZ8v6z2hdV0/+SzeArqiraybeh9R9LFlLAeZ09EnEWYq7HGGo3T1EesHDDI3lq
+LatQ/TrFc8Ue5/qunrNVEx643SCej2FhyOWaVeBEbyr4raE3fInl6s5q+XJEwU1
7+17ye9k8BojTv2G16w4y3uP8KB1CsSStp/K4t/ARCM3+Ts3DV8m01dn1xWyu4GU
EjzxHuUhJM91GCYrxqEvp76hl4ERV0Jku/Cr2bynyjJ8NQmPn92eGJoSMGScCjyP
ut83+Ft9yJh0Oc4WVgwW72ot00hoO7ecLG/hExEqY/cYLbhMTHL0tp9/8PVjee5d
jwQorXBXocDGG1J7P/DSR0PWcE1b3GpLmu/cz0jzTBs2MgQwq3lQxTBYeIH8xaZn
M0Bqy6pZ8DachflQpMZT+NZ/ufKP7MB/Mgd5HGHpqqSsYVQX4lY7PjGqiiBBmbtL
QNT2FgJiSKEx8FM5RAsonB7p1kQMMRGcn09totNCorZ0itlAp8bLwv+dZNlIEnQU
KOuMA/QRzzI+om6rmuu2UJMET+37c+jl1ypCuy4Tl4iHEYr+wqMVomVgLuuifj2y
3nz3MI2gbisH/T++zjed7+1ON/wPdwuhJLvSv7vXO6RR8dax5/ITnnFWHs6oWcdi
S5YXoY/sJHFrSWKIl/71h1dEswSLy7EfIs3fv65M293EqVQsfD8lhyPBY/+yIata
ZdZ1oidAwe0wGVWmDQDXbcBICvDHsVrtUFKzTfJtKIqw0wFjvSj+M9DcRoFegKcQ
yvv7PNVR6ePDZntF0eYWUl9IPI6rcYRBOTRWxDALLApqg7yVakj4Z7eQvfzSwftl
xVxtK/HUvy/n6xDCOC4LdBkAOtBcFX9IxO9RAJnCWHMUYQHVyBa4DMb8mErjyjSE
Q69rxkdqauR6+2u14Gt9cWRT2FrdbWhNwt8IgOHlLhpr8L8zRG9K039uUvKVzEkZ
2iyqdISffNbAFGkzdldKLDX1tLTuMsQOFo24E9Y8DipZaZho8H/vSZ2dmKdCXkfc
NUGcYKvcgm+1VyanqZQxSyqtmH7vnZ8koU87zpyMiUjvAlr7r3TCJu2tGPQjaNmp
rMMTNn03plrQuA4qT/ScnKzpJkZ01b2mwwkyI7Jeb3byAA8O5VOh2ZRe56VIMBpe
D7Q0+gHJAGvNT4sUfUTyK73n5j7L75xGZWOg6g1862iYw8u+XDFwjs9nExiwIa1t
S6gRBOKrOKvHldaJq1AfMmtNhUoTE2RuF+IicWHyqsYq7PMQCGMxojvsoEKU8znO
d6hZlurdoU58CiSUO0dvKRO2eVBomBGIiQrkG1Q9ZFBK9+qpuCF77RccBBpFcnNN
PlK1lDgx3n4+Efu4f0gSmtrRkUjLVKhuiqoJtEXccqWwW5gusdUCre+NousAMInI
8J3341yFeob7D1kCb2heAlYfcukNyRI9N0PDDiKZDfgkPbW+7MhIqMZJ9blht1/n
lMQV4kvpGW0nfZA7JsP578HbUJFdJ//FfyTV7jjHlOBZV2wiyXDIKUWP2/3lvq8c
QBipMvmqO216ixeoKe6XJtenVcV6+doE9bUWYdxF0VU7TFJvDA/qW2g27ZlftkaY
sllFMOup4f8aEoL+Vvc04+z6nRE8NuqIRTHfNeHk+oPgd3jiR7hTcbTPA9iqoNGd
dUO+PTmtrFrT8B+LWasNm8etuIwwY4fgzoBh+zQiry3WhlTpwzXCgNZWmay+okCy
Xh+eDxAMa5qUvcKpDnFiOPTDfzTP7Cu204rcK+2/FhA/QhJ6/wk2pGe2UF+qmGlo
VKQWTM1EhdTcdXvus98g5eujsHIpMaacHq7cKIVMZsoplt7FLINRLjAUITsSVLNe
+KXB51DP+pajcHhTjZUMTEG7gcEMFGR4SPWBDOTThh2zlxdTGaay8qnofAJySBwf
GtG9zaq90+OCnw6MAd2/ODM4kaMRaCu8s0WD5213LoQ5MHt4fj/aNF9Aes5fFJIT
m1+RcJlyohCSH/0l4Y6hO+IBfRLcGtYNH8siSqv5wm10Ad4rtI0KvIt/4VEFF5er
3flYt8EbfvnG2z1lTDJXwMvBawDIjYTx3D9FpS+z+LRmbMvt3ad0H/WGdPGh0d9k
qBwrLeoqabKytDqLcNxilmXDGCeBJt6XY6LMUyWqaZL0r2951gkka+zddcgNdboS
o9VSwD4VD+17a3wdlcsVYbC6sVKxJeVCAwS5u8dF/hpsevdz88CknFWTguxuO4Yv
aNE/uDmIn/mG5QbEh8ifCkFmryQQAiCLQRVD634rrKe7AbtgzJG+qquBpBDWNruU
irip2xnVY+MmdDmRAioDEKG76ViFzSCau4gNgsXnEbMPVxNr9FmjK4izgT8KlcY7
XGvFlmlIT/0p/nYzYNDCbj9dQtDuxUHzXcjl8o1A9sD1ugCUdN4XkcG10pu96r+1
zZLlbFxHyflMuDK2vBHP9lA2Bprca3eMRCbAt/ffszJt5YBiFrWbH0JekQFShhIP
agP7BVSrrjE7459A81VhTEr3ixFIYiFj4kB1phX6JuadyWqJW9oQcOm2r6YG1yZq
dit4uHggWNMcQAfcHi8gcV6c9b4ooI+W+vTIb3ils952oF2of38w+y6/ZG379ZLg
her787ngIih4lR1jqgK3txcegMRsVTsrQZmOHz4fxYh/INuknnob2b1lzWeW/2/0
qsbzGHOV4WKHDsf2OEhP/6YOIpSHOmY4z1e/6McdbfaukX45kWwzv4QM0RJwJJOo
Sm7RlGHUN9rZ+Kz+yc7nSeG8Pf2Y9HAcOAvSyyHD5Q7uLdJdATxUzkslak5p/8Ro
S69wdo2U22jw2Xqa+DgTQf15d62g8eDuNJ2nGJppPRJRXZbpEdewjTLoZvN8ylgO
JU+p/3+0E5GZQnmX1fcQrESk0/TK6HclSPskSjSG04wjknVAbcBSl1RTE8mG0hEL
Y2Zl1rUqc4S3BG4WuyLJ+Edj4/PgX3NdmtXfJ9XIioFrSW8NHugcuQr9lmHmyxIK
EgDixJYVMojH+CMYQmzTGOD1YW220yCVIR7+oPPfR3MATMaF9zR2ZGDnqZNaxWHU
SgcGw58s0BuUNyld/3/h/YaprmiqE1IArj0DqfUAn+k0l8clP9qC4L4htoC6USu4
D/Ore8af2G4nStKcDcfv+tYnTtIszlKQeB8sH0WqxoRmsa4raQuhsYXh+PeU4ruW
iTcEYpElYQx2DTzL1PpCvMC3YqDXc9NK5kZWDBd5aB4GBdA6s7HdC0fVIhUZ5DWZ
DSOJIXOUCIMtWnq05HVPtCC7sirjYEgW0BU90HNaTj48EtrB+imWOy4PkibAb3DI
Mwvf/04rJXzvGUHiIekDm9YRGnMQHTS50nn8I+dye0fGPgaylLZMpfuk+20GeY7w
gOLByTSUyM7wWzgZp+VYe0MUsoE1hN1l2ldRj4arAGjMG4Yw2W6Non8wKsVuslig
DoAE7ZjWpJJW7tCV0gJEBT4+ApGBoavqthjtycuybmgprSkXtPjXKgp5thJ0+IUf
SniOqoAFe2YS+/dDdRg3wAP8hIbLx9dFt2a7+fxAUAXNLJsvm9mcru/NmMXJJUkd
ezhhS69WiVikHAR+hntpSrUv7gX8fzwv8wZgzU5D+kr3cvESRMYp9cC/4n5pBTnC
v8qWD1L6pj+6Gmo/yq2ee6TisDbEAPRkXmdZwe3HsoVTCDmpgT4Wj2bZ4aasv28m
JAOPzpEDhATJFTDiuoP5/7EwuuPn3s5dqjnTdl8zdBwdEQJwrchteXXPE/5BFksQ
wEUiW+TIxM3ZvuiXkGiHeKjATTk0XU/6CYpR4poAWxeJ7tmI7Uam6JWo/aqXuuUP
rq5mfQ2N5jGdfZTAjWfgsyX9kyVdjBKEPBaBqid87DeBHf046tH1HZ/tNDNHpW1h
dgICP3IqR3tNIyQ+bcagGtwAGTaAKMehpt+PrL4qEbCADYRfjJMbQWBG6lxl62/F
3pZLBt9tTjfhb3eAncs7EmqGmKP9j/EJoY+1jaUoU1+UjghEkCnQdo86A6AVJQSF
KXX1iV5dBOtTG0K4ljliTr6jSaQm17qbx9PdNZeZrY2O1PVrJRn+rzbH8cyzsqBX
CkI1PmkwTPN0oGjZCQk3W+rBCvzVSvRAmF5MUIsoR6sP0pezROgM5w01WEna0Xdg
sFoIg1HqVhYzkQ36BZ4ZrUpnzHDEhMNPWAVOh2EJ/nmCgz5d+Ztf4HeSB+MqZLc5
rJWDIr6LxgdbQJ0ADm+j/sFxOWuKtFqzGZY6xqBkE1Vp2FCZjk6XiA1TgJIcLynE
bzs1jV476l2Zb2gvu+Qd0QtfqI9jtRMrSYhoGX5ALBl/EY0IwTZLq73Dkwqyv9/N
SP65FyR3nIcb2ddOcQ9xjYiaxZwxuD+TyKoJqUggrAr7gh5mDr4xg7/ZE5mcp/30
/SfCSclNOoHJe59tlBojy0h1yrb/PNIteLQ0JOnMEczmRaEH5TrdvtskJ3v7nZ/7
WmlOp7NL7n64bubO0xU+x5Lc4QTK7lhUQ+GX14in3WHIfjv7GUKpWtf9UrcjIv7w
V2QF28MY0maHFCjY/cLOhhMof3CMguG3sxURErOJ6KhkEbb8qdAeGFuS76CyEBsd
Ewgq4csjilIEqH6cijgK5oYMikZk/wFRjezvrC5nChhv0tTfueL16pBJ03IfaaNW
oshwGzB5w6IFD1iPAevTA2sL25tl/QeLp9L4ZatawoJCo/0YvXfouEIycHh/8g1k
3SlsGQlOrLPMbqr2D0lWt18r2Kmp3rI7qJYJ8H0Lklk66VxZdLzRj6iUjmJcmfwt
e47O82b1Gu5R0RVMXOPB3LYxTdHuH+rhuSiWy/JTAmq9GC27kcscRfOZZOP+B+Ad
0nJg2KaTZ3Fi++qvogdQ+IbUUfCSA4Mtz7t/PPSoR1y4nZyJlDqZgxsUbsMW3MNT
tukn4JTnKkI0nYmMSlM3pidwVKYCPzEIq0jYtyp1+f6TlUR+u9dQmpeVWfY5ZYBp
x3f9LE68U2MDMsiRsSb2TyzenbGr5DXhuok8nPSY2DHwk34pI+c26XqeQWwju8+R
8z/DAyerGOIQpPIsXExaYonwbivrCn3wfd1CPhYZyfoslDYwdE/NWo5Wt5qqAMhz
xPwYnxKS+ds+pHyx2oXrKQIVDCmfDC4J40N67TMR/3CFk30ToFSW6kg32Udwy0g4
WV3d7SA15lxngs4zjst/blllWf/0eJ2tL6TDYWUNtApqFy3OC17V8ybYMGy50z7h
1A/Dh749L0xgKnwOxJ1nBTutckgEBFNSlAgBfovgF33ttnmWe+j6Qm7eldFp2PrR
q7YNPm97QBo9nU1mrKfp8DpQ2vbTCHSVKmWCNbjxc2IfLmplvV6okrY6BnCklaOm
kcp5R8Co+Cynmn4kR1DiAXUX0Abv8Vho44vn8s1r4twDFNmKujsF5hxmOB7GXuua
9E6DctRY3gCmEJXUgavUmpaEZHT5S2EIZ0fPMAzSNQ8kbBW6bfIpPPPv1z6h/OyQ
MojSD7IH00CHqS++9OplVBFua69fyBLT2nZ9KOZ0/wgwKLpgz0T4hD39hIAydW8d
KztdTHpmDldkE/fOn6ggQ1n/MZstwivv0Z8U7EbbJ0+RHPk043v9fSPHBcc1oQxF
s59ctggnFCjPGzVPXqqRxj9rGKHmjKhNn2gkYa6UN9pU4xf5z8x6ZMKkNhXQB0Dk
rX62G/T+gfPeXxIWwqKaIJArGwLmdqCmpSEBp42iwCpfZN9TfrGfsX82D+X1H7DC
Aqq6NTu3mXFqnDgGWxwpAjkRTf0Nn34XAF/J/p2Rt1WPXffhPjKvzkIrIUSJKSBp
X3YuWQT7RY8IBuTg5+xr8BQl4HPOGjSbozcKugKi8F2s6DK7jHJMh2apBTN1awJK
bgVnlLqDW5n9OJeY+viYrUsOXbYaajufgZp9EBIiFxN//FQoN4QG3Z/8zLiknoJZ
O3xSx6S1F33O4IkNEseyxyLLsEskdQLQeuaje8EaddbQkZnquwEet+NHJrqPlkjB
F4VAnWGCi9VYXa75VVEjXCCOUoOeAm9xmEEXeCEKrimyQxwvRbAZI6BIO1GtJ0eP
ao/l6gWuBGxJx8ETDVwCDz9kQn6kNys8DbXO4TeVhR0sAsaRSldGQEP+DiuQc5fc
XllxuXMHXo2Rx0LCNKl2OXXWYhfHC+ijR8gOozKapXgUu23NRlOlKui6JIfDvlo/
IKcH8J0WchFGYqL1EoPoE0JQRNSOsO7fF1h72QDv88UUNMev42wU53AWsE8tnMG/
K8KHOSJAKdw2x9Fkn7liLGapdNp03uV3aOWS6mBhRAJjolwXNJHfoFAhubGFDXSn
larP45PGtlUpZzr2G6ypDpWGEwv8c/T1rR5a9oigS7nKFtcPmujMe/1c/h11bnB7
PxeCef7snhCUUV6NFUSxn+lIxutD+RQsiOpCPBbbdHoS4Fcb50CwtRjWwmufX3BL
HnLDwo+E9zOmpndoZeTpxAkQ6d3Wqsb74EgpwjHS5iCw2YLw4dtVdtGizYBQkA/5
S0pu1bzN+8NkLgcgesGEStGO+h3X+Z4/8rCqvFFsa2yiHl5EG1eS1kvr6yDB9qOZ
LizmThYAZ84krkTzxKRGHaacdwF1ZEMwoEf9gsOoWG5QqAlYFbmaf7L+3htuMAWs
WXZNEIY3IoiSlC2dNjcnsHvHUxvq++r2TC4inVUHQpPKOIBfc6qOwbN8GQzwiTzW
qA5SBYMxYslvY7PCsy3sMX4g3sbmcloM3P2Lqm8AGcmaNnQxgNrYmkzU1hMgArVo
01MDXMmjEbZA7FRCGOB+uTeCduHACVczEbkt6PlNN0kP1lWrd3hT6GiG7nTAyWNN
YMlp7U+iK0f+GB6MCNhcOOEW60viH705NBBXJl70kFwzIly0FRy16UtkLIwfL93J
57mJq8OIZEcU34NxItGdo19yZ+QlEdz3zWKbD34bQr56xh8o9XnrsR5ig7y3Li5y
kjOdJvbwu1+T8pu2Enf5geBCD+R2xxTDaJDP6VSEoy6YJv/SRP2jrpiMRImLugHw
DPf54gpm6yVEc93QYgd3HIsyM73x7Jz8t84aV6fe474sXxIrWkeYC1QW+e+PP5tT
w8+imNbBLlgTq04ZiLUJHtXJwT82ge+N2UJc7utuuCdSQQtg5IeTYl6arrzRq5F3
8zTTWPY66AqWzZwu2/InKHno9ovKt3JnbX+UYxmsEhc4w8bihjBbxnqmu70l09nn
F60FoGQmQXVbDGuQRSnWvkOnI0/yYyecPw1BEg2bU275T0axPG2sORu7EtkD9Jqp
IJeniZCFwn18UiH7lrXMthZVcIqz2meZRYFl4CX4uK5gbyK7v3qKUt1/7ceYdG3b
jru/uKoHZ3Oz+NsXeh8kteLZH26bhQ2+23wwoZT5Bj8Mgh2UupU+/VNCkNd4qgbf
aj/2ViLeLit4J/Y8WHp4wkEqFgJVSDfkB8GrHJcvC8ekyCKQzauKPvqfkODSxPnB
aO6ZhaWUMjX1bj8e3gIwP7LgY54hmChyR2/+cJ6tR/Fh+myaSSvQPxassASvX2C7
6LZAsq95UOKDbSWgtZMT2lZ0t2CL4Ew22LHV8dtD2mnHfewwDGjqxPLV98k03WdN
JjMJwZx886ZcOLQPHy7QSiDvfHwK19I3Ha5pp2lm09xgpIe65z4oRK3ZwbrN7KXU
UCALHk2SzYXrdtal5GLmRV5tjVfbxUBSxS7+EATCxqbrfZse+J4lYx2ZNrdJblb8
/d7iHKtDxHILtlvEacZPJuekvOgWbpdYvvecHeQPbnaOELKwT/70eoSAlllKrzpk
IRu9+nVnBBMJ7rDQhywXyMXViJ4VugLtljJDSx5SV0SWG41VMz6WlI7BclD6BhE3
SHwtW3fjwGmwWKl+f7S4hK32n9WjqEvTnUMVAd91hDJI2cQcWLkL9FwPSPJp7aPm
9xyfUnP91fNfMDuhy0q5eHUsnS5eSVEMSgFwh/ke4pN8EoN5xxjVgvMZCvmSHfwo
LiTmscnZjOnE+l3IRbkJrd7mqoJyu/2DwYqE5ZKxa+fJsBzFxzYwpl2qfbwW5Ox7
L5WFB7/yRJZE/gUSZCKXmt/fwJXzfqUddYuomVHOwqeT42A+OZIC+Y+4WyGa50U8
RPpjrnvs8gkt/4QlAdh8FrZBbCo6mxMIClKvXxHjUYYmzZdDxF7iWbn2n6p+p+gR
iVPxYFc+BqwKpU3qt/uawH066qcf7juf0ne9RB9rED1IkkryuUPRflyPi+jUKs7Y
4l+Z5FvMbfYSqQU1ZvlPfhYdSH7dN4F+I5yjo/bCBSGfYeOCBc97JUX9ygjvO//Y
QWxn0jKlOmE1fenM6vua18HHP3ri9kHlyCWOPpxGW79w1X3fFGYibookDY5lpKvz
5qLMRy3lZ7HgFpk+FlHe5fnA19HhFSQy9QwDYPmALo0+SEACfnyrvxnqJscc0QKF
BPZdiXhSjIgo6PqxUngCYBZ3o/0VtPc1Y459URSbNmXVmBy1yv8STfrT75bb05PS
p8feYnDHIBiwMrbgVLgs0pvQffaX15DhwYaoaJSPktVP0f4BznjOcNnRHJSJ6Olc
Q+/01llQ9iOh1ZrBOPStfWdlgH/+26P9tB0UbbyYs5VxOw6y8rckjT7Wl2IzoCpD
QUGaI1vxJKdon9MBw5BiuH7MZXUdAJRmuEJLXfMkG3kol1PazULwg06J3pb6L/FT
pzxiJKqzkkuEBKMJ4s9B6L9LJ836MH5D4th1A++ul6sTnhnI0ndJAQrMvfLJVgre
knJPxCwM1kkfupU92g3+q4N+JCHTAWEYqZGbZhNmnrkaawZqUa3UL4/usRA3Uw0Z
Yz0T5XpxWSYxWb2IxqUmYsieD3nl3lGa69Eam4+bUAk3eAwRjRbm3GkX49F+asuq
mX7TcRZHEYVBSANYaTFSJ+RdvoVSRjSOq5N+AqWHuaLpU/m/WYm0XdvINeGhzimY
1PBIJ6uDVb3Ixim6+yvlFNzIiGSVHfckBUlzeMKPX9sN8V/8T7Dn6YKo6SpH/jwK
4GL1nTiNdiMUghDgGauzqFxntmAP0FlZLUhukYVEzlU2LlhBQ+sQd7UxIcZt4P8Q
rqRDTPPoztZnyxvPmsVYyQ4KGECNMP+3z23t3B1sRInQa22bxXFNpAuwAABw4P5f
1A5XjmloXIZCQCPG4pvilNWBE9JmeB+wVnMDJa6XAuZ9tKRlXNXM1YU8gSi12y+8
uEpLihbW4vuuNuejGJ6UtCcrb1eJbn2VF8YCsaGl2bKogVPLpNug/8zmrMzGS9tQ
qn9HRFie+uFEO/gU6IY5uut1VW0pv1hKIKkwFHTmKqPQlBl1K0TuQ4pi4F1ywyAY
j412GG7/1MwLwODFilNYo/THtXXDaa1FwoqYjX3Cnmj+5NMPFqqHCcTuiiv2PClc
ta5bZAvGeqUfrfR2rWylbnQUmTGJ2e15nGa1QRXW6kByIUQ7hFFpp7/hZGgVWcYA
8nEFy5JFv0FqAfEyICM1+3ceeC8CB6WOQxQBqpHW3U3e79ytgTTWuv21AaWszZTB
4d7uK1hHlxKmBqMBEAaQ/5GRtQnFvfHYX2qjbzy35GzGNGJ5m4GPGlQmdGoKP6gY
qYxc5cCw/DDI4u3mWft7kR1C6neGTZK5zCqIhVLd9iHKG6KzEvGCUo7ohdL/0aWb
egzSj7btLh4BtExKgrbQDm1k/mseZmRi6KCEZUa+24zgbZfzxzuHYoezSmeHDe5m
kDVOB/4fAf+4nvUfRKmx7dZqDPrjG0N8IhM9CZFpzae2vwmuIGb+6cB3Dh8o3Bmx
WPS2K4OpytTwhrQtwlmpmBU+HIVGFTzuo9J2IY3Yg7VtPTkFyfDJNbwInm/sLYpa
eEp4WDD/lZiNjobmj+6dx9Cvh3qcvIpCnjmnj0SQVfkV8GzLLElSCqQaiuvu6wiO
cGUb5C8fjEtf6k4pHny2uhcOAL88bQoTmTl1PccQy2yDtk7FPk3BG9dBXGUshTqV
Wu5XqlRyMOdF8AVfIXwdu/MXSBDbfr/o0dY53IBKVBJCbHGi5duGhYXaOpIFZsOf
V0y4CeFHjb17THmyN4lgOaefiTbO/3e37pQQmD8g8M7mCclrJEyFu0dOgqMoqZ5C
PBPKqQW0AgEJCJMJ/EHFpXNGc2q4J4voXmEYlHha2EFwM8J4Eli3OhuoDLnlcts5
ljarc5DcU8lmS9vo87aP1TdB6uclUIqm3NPt16P5YKrHYiY1HUCaEnuJmalRRsoH
9rMRQToAI39sf1FyegNOGDidBb1UycyFacciiGb0wVbPREqBZQ3KMenr8T/Sdtk0
mFVB72Xa5n8CmbdJSTmcQCLo9I0Cy4RfW7/yzBKkmgKyFAFRSBIdZu7wLy7s5y0a
IrVaYdDRP2TnTSwKalCYV/p2Vq5vWl/JKenJGVWqs++LS1Cw1tYUOQxuG+g8gxpc
eDd9QJWZ07kz1GH2EGddOL5KlaCifaNBHt1Os7Xa9RcNf4xlganNfk4NUX37Ygge
i3ZATFBy+NupqMMGUO6EkWZJcp0e+idJjbRaQCstxFu7I1Axo33EdK5+X13wX4Yx
cSgJQZpgfavWmLLxNgdBDFL7zqBDo9fxmByx2du2q8ppw8IPG/wF9TKhK0ypUiD3
8A2jOdW4e56Cm7b/DEdEjHo2ZxE6wX7EXnw2ZI6e5gj2JaX9HWiQ1EF8BuaGenSS
u+IEJFIbRNG9GOJ69OukMdhgZBG1cZFDnC75HjkpP01Ukgwq23Ll3kpzB588MB/N
qi70gfqJmAjHpjHUIdFByElOsbBaG5e669qcKGnpK37VkfB3s9MvigAGcazCODkf
8VEBXZDAAGmfa+tlwutW/V87MKn6UxoLFadvOUuB9P4I4qUYrGUfuQHfuXv+NbHN
1qIylX9mR55b//p6IlxxilhGhXabful33K7qOu9lrPGJkY3cdBTHG2N2F5nPsC8a
0mj4CbAZXCiRJlV2r7NxzIjUf94jbW1HU/1MFqsjecW4Ld7IrKxuqtf87Rv5lje8
PmUqlSjtv/uspmJlKizzy3owOD2Dafrr8KRj6510sdF/40juwAQKTK6+xCB1h65s
OXGUNmltguXEmVz1PPRN5wzHTBqiZ2LXycphMfXOqZLFUVlRBaie608zl0p8djeo
zwnNajapKP7DujuAEZvPNUzzX459B52HFzng2L4zA8NSxdxL0LoKCPyw7yK+Wpon
JfB35Tkmt97RoBmn730lxK+pbD3P3sB3/aVNeXDx5ap3462DgF6aBDvee4g631yz
DMtOcOPAfvjWewuZZ+kzXZOyePtiTmLLCberNHtl8v2ja0edwaVk9pYleBB1gRbW
8Cph/9KCNXECofKFizxgJ228H1iQm7DlfS9nzAEGKlSysHlCGh6T9B/2r7bnIhaG
F/LstjyZdEoOVWh/6UPmRqTqI6OZdlET2onYqsMyj5CYEhE2a3IEpjPCaYsyXNL3
SmmznJQGhLwsmJW+uT2CSB5RpN1ba0uEzlpD/4kn9DeS8vvOSKhl13YBMKIl8e/u
uAqYHNRcGBVfQdXAWFdnuVqRrOMqG/ByHnLWMLkeitRzEmOEBdPqZLb+9ewkwJdk
uj5oJ4GBkqQP8oc2csGrn2i8fKQ8stbRL7/DP2uKyWy0C3YeedPn5qShEkIL3qeX
lUKbbJfM8N5jJTXHy/BaR3rjCmbImXVO1ZIHtXe8MLJaZjO7IsxkmJhUrDyhZh5V
+vpgcH0PJC+2mnXlFzu7SrUZc24W4HIUwhS7/fFYeEt54ALptqNfgV5Sia94tZoQ
bh0WBZ3OPp9nQdqTVK8AEprMry3wxUCxbryUL7x3DV1Sm6rVA3+K4mtpsU0m3Atv
2CU+/59g81ozl9scyxIlETOaY0+PH5V/fHKo3Qqh/nhzCy1b6+xH9O9Nne3fGG7S
qz0187xXEUfFiIOtoRnk0Y66rgHVB3lmyi1eU143zDlmpdeZIKVmXGZ3wGHXLMbS
2FpDIOnb7HBZN7WT77VXW92w7+m9FotCSqdIklO3RiZSrOPg8xs51JqfbJKyJ1oN
JlJCPd+hbcRLohyf6BCtOm4jCsarRiqWCPRlA8GpyZ7Kwp3zhbugBAJFEpgF0Btu
PbxuhKWtERNxkIz4KkpS728u1rGAZzPWqdbHiv1MEMAOtrFriI5tP5M1tFFpZMRY
Wrib6nR+SPGq8PJ4gto2Rha/lzEYYzPb9z/1zNm9c0p1w7mE3GHG/d4XKS2634aw
8x//NNkPhN6SMf7E9UmBqZTP7jaPl6hmxrgD4gjcP2QfvkYthhX2WGIR+8EwEQvy
IsXKRQVAYhqcvkwXA5DahURV85ieU81jZYIdyZ/KfknT+aDiGIAJzKpE1/iuszkR
pl2hvkPn9JfFL10RmZDkb2dvckljP8qOMNlSDtnjLol09uGP5+LCUFhcWRWWABjw
D8XMoNjvh3+HRL8klugnAVODoW0P+1sN4iqzZF7/Nkp4PcUBFkQoxt7VHdb/FB7g
OKsfZpITO2vUqQmTf1yCrnfEhxoYFY2HVqKLfDUXNPDetTheXnQKVuTrFhEnfgAg
SHbyoS+UU9FGhRAkALXbr57gcbSlO/8KRFavS7DXnZQQvGMh3O2qMb2uQborGPYl
mGPTieGsehJLRYdW0622hqVQNbHsI8rZdkfk9uJ86Xy4/PYONdpRhJbvJ1GvNiQn
7hILFsFW5vO641BQEUkYh9tnZYLjf5LQEYJHR1RSmYNdlz5RDGtMfj6jed4MfwZo
+AOO6QWYzswi4cJgfs9n7wBkKj0CRaEULYFFZs8d5AoOCmiJkNj/H4C+ldlP7HWq
CJzi7l9dCgsVm0lE8dgp+wRMTYbYutQ2CCwlpTh3DDcveV1fB3CNVPvO779Yi1r6
1zjyLveCjehkgHarJ05fdsro5CXpe+U3ThLp5osXzLM5eRNVA+OQiVKkHfjW7Ror
BqxHw1dRrJIvVihTs8E+myE4zOTzKfNJScGwmOL5CBQvWWwDsebwKorMvPeVLUx3
`protect END_PROTECTED