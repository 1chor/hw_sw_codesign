-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o/VZWE1nDCMTzD+MFVc2jzVccqW7qIlULla4YD3yWdjH+NxFJcDkWv+o8UJ4UY7zlxwD3PSQ4or7
rgHVf57HYHt3Fu/BlJ5MYXgAXHQr4ezhjf1Xl66WdW4WA3mRWdD7rJwoqkiywjlUMQZb4af7XJnE
dY5bviT2gVhIPilAN+/7U9b6q+jdn4s/OQkXyCPsDbcYM2kkuvAmyg9DZkAyTWPAS3lmT9Dad/5m
KmevEM/69zYxS7w+OnGKbC+yX3koEqeFhlg7kvQvweWAHTsgzsYnstKiP7X7MFgAWuEADhjzAkS+
5+BGaKd6+hVbNWhbZ5u0OcGxbe00DVkQMGuBiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
qme6d9g/xlC/SmoXBoKCaaMssHTX08ryDImxhWNiCM6E8gBaVNDY6hkYQlJ46JAEL4E5BDE8OPVX
jRlWspHlyAPnDTL8agjN8MBzsWNii+qLsgU3Oh1i1p5c0j7fCDAYceoCJsVXcJG+S/fkcmhEHk00
C94J6HM2/Y0zjXcxm1cCScp0XHmhbWE6NNm7goFii+gPzuUg+bUEvtIIVSmdsjSqdK5xu9xFAJhc
GzWH8WTDgjuiH4Pv2wwomGfwK4ghp3gFXDZvyFAEFDJj+wKEN6MSYzAGdeFurmtq/wuxn4JvX7rp
HHwQDpB3dPTJCA+kIuABfyoONpQZCWOVG6N/l4TgsMBtVlvYLFwK2pKcO/WijFC0+3jHu3KIqfzH
nOfRlnSJeY+MUe/tclR1D54zgmxthajvnUnQXbhRce5Ht69zXuILXyCsqvoB/Z/G+jOreQk2iPKY
zoZU1YD/C5ICeidYD9nsOZqTNnOLs3XJIY+6+yCgY3ZBBBGTXrmqoUKMXPCAmkrZm8FGSZcXqmUs
wd5jEPWn5oS1ZBSRNpihJ4xcFlECGSsFaz9r97pcDe6MDZbUGQNy8Mh8slcMURntekbQk+56Gu2I
UbWlLI8uKXH4j1AfHoTVNP3v4qvVAjrhvs+Jc6UsBPkiOwbtFtsUqrEXi/2PPeEp4ltmdptxidv+
BZEQdB9G+mp3/BVzV0KgojaQPXd7gkOpmZVpeFa129x6AqWnlitOcjwCTklABmNnrcEWWWJJbdDm
PbdMGwEfnW1hhwWu9iOH5bH9wlc2zHRfKGPz65NEkxRAhucKOR3CJNyCumtzY6KZRxIwdoCkLo/M
8frEChYdN1pLxZ/HWWhvnXJ3Hqy/IEB9zfvh461UpOk3eYFyhKoROqAQma8XnuQJzVoA4j4XbkgH
9m71W1rfeWkZyFb+sdBr+RhkPTzm4p01sMB6WTekOQPiHBs9B2CnAp4RnIq8PL2mhwcyxcw+Wsq+
kOcAbvo6tbcEYFl605pqCpQgdxOzG7kx7ZhLyx03AvKsz2rIuiFLk77XjC4Lt3ZABMFj7qXVEcUA
Le5U430zs3MbHnnjaL2k8PO0RxwnQeAnV2weL8mJQERxLSJ621mgYO43WJXLx70cDuoDIzqGW41u
N1pJcr8vka92K4BK+A6jU+WL+L/FlAhrdKhpRovT0Mih1XeKs4GWdsWvnoyoh+rXS8bkLSRmdOeU
GPHj4iS6R2ooDqI5lJbfam4gd7FOECnDu1IriwR8YtPI8S/vLROuag6z62vUvmha2oGilQ4emUZp
Gv7r/q1zdWVuwvvhNtXTjT9qA4B6O26hgVOOBV0EJS8qsvS8SATNJkLZyCKOvzBhgiAILfoXNUYo
z6OTHzSRseLYll0H25yX7xjNlBjqJ/Ywz8qZu/E/yIQCbX14s6KBkc/q0CyDdI9UCdqLx/gpVsFI
MEn0zm31sYOSvVdU8w5l7AOCrs8A7anYgybZTiEosKNeTGlgVFfxtd/Fe63FWXQvVf8O/to911xy
vbhgOri8grSKYzB6fw0Un119s11aZLKL34jZxvmH/vQesreir8C27RYkFPAituzXaG6PkGhZPgRb
sPakKRJuXln82xF4WGQcVKNfdy9zd4KUl1zFLnaSJ+pSyW8lRl3IeqX5nXx2C7ql3g90gTjagFCT
6z0dtSIDQtIr0umciWuSx2BOClscP07hrfYFDFLQf1tnUuZVz9MC6mZ9tONWJpOKzp0uuYCHIAMr
QKRm8tkDyEIM2l7g5095GOCctO8fk1seF3LC6JOJNZ3rGk/aqojRRw1D68cT8MxJntKnKozM2Oce
cxSjMfcP83lkKc3wN2J+ELiAQjG+aMaqBtf6bAyX0CjWbBc4MgQUqs23JpSL6pNco32Z4cO6rhIc
mZM0ngJZX6rWZJ2dmzfs5aSXIusO5NxAuoSEL4BQEgyd6x0zbx769iZoaPGcpEn+6jz3/ERk4JCW
YrfKL+VfYMg1JCXSTqg9yr4gh0DSEjQZES75wESSwyavbdkNyNIw90rILxMUBVGJN1k4HTW1p3QQ
RDmyyZ+woSwFm2KpqCqHzyBD0q9ZP36pTSQUTstvGMmRs5V28hZX3q2PF/zFJf4V7+0CLt4X7coa
qncghBIbOoiQ8h+LEI3NaCD8w/j75d3MxPUX+nA4ven1v1b2p5+jgtVN/icNhJ60XuAAyDfqHKfT
NUgQX8I2Wpn3k8i2yBYow2yyeySwZDumdK0PCzJ6g1867rVbaaGh0KXkus0g7AbqdJDJejs/MODO
+jla4BNwlrO008fqNuKIZ8OIhMbLrB6SfS5jrkWZkq/BlZ/MIOrrgk/nQRSjqI0M1xSU1THgB4B+
KIIPhJybMjE1U5lxoB2BoqI0tM8vlFZ5RmWJMblplB4Uc509nhBaOz6M8+feojIrmcSF1rDuZAD3
W/CrfQSYUNnYPDsFcWL4jtuLNw4eMgu1TUimXLCC5Qu0Nb+2JWxMksYH8QQqmnRL+HSxHYdShLiT
wCONVOqiTn2kpBHPf+gUWcUdKts3xImME3LbhvMG4b5yea14n94230u9/7Pz1epsNVpF6oQ7HqAy
sXCp5pN98hFlD+zbfJpECZlyIVuqS6f4FHWqshpcwPakzPpxvMABjogkoIVeZZE+xC24RO2EMlzm
DQ7iuj9rHokJ7TPwM1qCdbXmBfcRu0IdHjAFQiITnU8KQjWyKG96h51nSqx+c/QNNKMZoM+d8s9o
ybOWquAFpzI8ZHlYXBZI5qIiV8oavjCtGiY9LCbZamFz8o3Iijew4HIeBNC+Y/hwv+uVazkPHVOc
TKsbAyZ+IcVhTH/onBL7c49+FmRPE5oVQWe7Q5aqWMy9+8e4XU1SKWmjnsOWvx321obXc7ATMYd+
Dd3tk+xXsN2wIghy+abI6zMYK2D6ffcEwW7BMJmtwYMo4PV1PxQT2NH/8lNPZg0GxEPFb5ebN5Ww
x7Jjo46KY2rNVcqOgzEz7cOfGtn0UQN7ZQ5qemPxVHECaupseWGzJ5kICvS2Ihg/timPLcUkLGAV
UzMny62onUrbD96xYI13tZu5ZDyXD13WGHte42JErx6AtKFJ82mAKeh8f0ks1Y7vsf8ZvQGKeqMI
8dMAkpFu4i+qKTcaXidKgorJ9hBd7pLvm960/kh2J5K0UihC1YshWi/FH9H74KHAShWecy6XlrP9
t5XX40NesyOyVZQ9gz8FZsDC+xOPOA0GQr8ndAjFlVg1A0qlYivgrS/h+VqqfZ6Ty7emx+ZV7gZN
HUTM7h+4kyQ1vBHPUFaHwES1pFh889/3YI53T8yCcxYFvwfWayJgySkzUGEHyco82F+ttWwDW3r2
NJWMag2sXkpHYxant1xqlbx5yvXqxx78pB9XwjS5RAeE0oI2pNWmFt89Cez7JABI+F5xf4v4eF9k
jxlM1z3/N1zsjTk/wl7X9k+d9kLEycUCuO88UIPOG9YG77bsZm1igRp7zUo/ybCLtWrQ0ycSwixo
APykVw1dEBNF2w3P1pXWHQYTbQEQd/QJjcUPDhyDc/M2D35jl1uMECM2cxP0DOzXJe0MWnHBpbAa
aiJCnwO8i5tkd9SJMjl9w5jaxBOWDmT6Lgm0395hA0pmQpzKKyQqfoUvCavFKqVePKBGRqyKAAto
bGRcLPw9yHMyYFq635ZXHGxi0Nj8Fvvi6NJCGmJ+4RS8gM+Gx1ElXJp0XrDnysryafZVilssGn4z
gGQGZ6dm668dlRHqjwQPAIOqbNVpcfAe10N1jSNTsFMTUXnd11UxInmyudKnOsBP3LR0dt/dLHFW
5QjaA5gGd5viw0n+0SqoJ55kd9qNJ6eObtuulRsXeUNPIa8uiKbCM8Bfs4aTvMkHCreh+2Q+urtV
1ug4DK2jCzM5X3HidZIVhMEarSnIoRYp6CkUdqnDFGMTC6JlzD6j4sJrNAb92fTgLdKhE203MMTp
A1HhhuQFcHvMvHon4gHVPami/xrZ70AQ8WGKycRTHd1BIv9jx5pgwty6ND2ZfjfnrK9DNkiD6EdF
VJVx2JH+1CmGsntwKeH3dbV4rf8ZIHirbog6CL03/aTMGDh4p00urHxHmSXCWFqnUfVbv7+5NBTp
nsVFaOKJKwDR50B9JRsjytAOWlJVLKk6V6aAJff/ALU4I4Ky+W+WKOcoDIEW9lnTyqEsateU34ys
cfVYtaQ4Kmwa4sXtol7nlCi8w1o5ztPh70RbS4WsM8hiYu/8yk+cZLNlEoGX0zxYjbYA2ECvA+L/
FLJvDj2gbeeF7BER7KHrOhuoWliiVlKcx+TEl+tf1VUk5drO31qlByl7NqnRp9NpWdzTc3z3g5Pj
EZTycmRtGI9C6r9asI0iHPVHDH5kP0mUb13cg8Bkd8NMnVpZM8lqV7WvObYrAbS2QFZ3VrSKTB12
r1JmHkwjE/PCLQBovp61NuJYt0LY32NHkY2UP/GIUZJC6ElfI+gF08tsl/boJd7n4E49EqqbgKuZ
AwzGubyChsZKuskJvLUx9cF/UplOJfFqN6QYAHz3hza4hPLX5DDx3YcPlf2UVy97RvQ38A2f/zuE
S2xLHkr79VRVydpMNtS0+n/jaocAnDU4Saw66mMXPpolBEbu29ePYGERPCryRL6hqIVu17wjrurn
+PJv9bqvNynF008stwT8NsNONkCfROZxLCXmfmmXYV3KpRNCLp5Nj6LSef8/XjZm3c5UYrKERKwb
DOtUxhakKaLEyfC6LaSZGnFbRf26+F+AOfyi3tw5hY6jImzny4mAuStePr5ClD6gyXzRuSx0vcMC
5+4mzFDYSNO9Bjp+6g1X3N0pHEHLSu95yqs+frjutho1W5nq+SXAW/1f4orcRF9lYbFkfXKnU4hs
LKAjhmLFhwFG6B4aMp3cTru8yIH2NjDVkvR8C/9g5QsMJ/yjwB43fo4DK2jCzvDAyWHF4DT+Din+
g2l4lLSwg9jxtpdmxVNWmhehY8cFbIEDjO291PYzeVGfRJ29pKlHWwZTvzBG40BmD6/OzksQt03O
W9yLbqmbrUxof8ltjJvBez5pRn8qqHMgNwNHwGPe4kEBuYMTZTQ9XR5idjXOrokmq/MHncloLJes
0mYeEMfvN+iA2ezW8GpYWnzbGj2al1ESi95Zi8PgpQn3CM3VvoKftWM6NXxqx9OUXubHqgO22ZRu
FTwM/KPYn2SkxF2MFc6+FeJ2WyeRC5dhkYxQETk4/L86iRVX+0IeUUR6AQg7QFwGFlQ7M9c1WO9a
QSwmZoeF0FKJVsq3IK116VfonDDagEBMMjtlbXJRkxA2yKvvVUQf8hr3sTs02qG673QA4BZOCapR
cA8aIPNWfSU33agOV5Qim/qtNs8OUoInwQ7c9nqSPnUwF2rwAdu//7s1bFJf7J34FNzaBN3/9JOm
GbBW3ceaMDOanLyZFwIY0HERC6EKhCCeOonPNFLO7AGNn5/T/BhqK0z7i2w5rPxNav4R0n1ql1pj
xS58OxA99T56Dv/DDwUYXLT23gD7Upib84uQB5UAGqzoDK5Z7KuTT7f1r5h6bgBxjoq3xb18CnkP
xDLhRa88rJSWlrryO9uyfpCizahwB0nXQjUcKO2VA7QahGCrn9AOoci8lTMX55U946iJi7ilOJ8m
WK9rj4eACI8SOaXjpako3plBV4PdfAEwTSRR8e0r71Oh0+ARVbiGnS19JZeONVaHfCCglIIUWR62
G8FNVu4gcdTlRJp6q0RcYYnPW7m1oth0yjXr6LZvWD8TbPLp3GKa2jBBDRxdspvLPDHfCSteDR9g
sXLiFm9tb+CcLmqig0b3rklUxOWVhkt9+hTZ6/r8VXyOjiOVjiqsP4V/pX5f6KYOeiV7JvqHm2sa
4noLauXzmLVSqsjhHpDIVqhjckoVQtfyH+1zFoHuDwRnLimo9olpLhwgbp7qVUfEoc9afdyqgsTe
up9c3B/MKCWGWDB6hhZvOYaBAY4ah1KXdoCLnztJBwNGdQIEbU/mhrdqF0qHOdSuS7jXg+jjONSl
TC+00daVVGqnKwyOm6E5z+Rs0A5pyCDg1bYk01slhRMtBRyA/7djxGMkSNMfbjmd4zxJV6lWMz5p
dvBdPCjfnZzIYnrhxAcrnjTRqEPSrXHQ6LyiO8pLJPfpOWm7M5eQ5y84WuZpknvO45Wc3FH6d8rK
fccWZ1ODKpj7SwFUylF4MW+bXoqKOr3Z21gweS6nbgfbvy8l9BO6h1Rl4GGLa5zsAlxqmcEkzkuw
uD0v7oOoeuxtoYAQ6Pvhdg9fJlGQDcjn4qOU7zVGXsgdOjGV8nZakt1hIpBLTmd0F71L8lvb0MDa
obPkwXbsb5Y6qd6FZuEP8cyEdg+XyUNSzVNX2Fpx3qIqPVuwt7MpQrwfhGN8A8rR/6eh0jrHOgCZ
GghYgyuVet9JSct2yxkZYuMnP7DKLdbso3xGuvByD8wHvm1w0lW5m4S9cCXXUppnMkHvRyDHMIUq
SwBdYI3S563SVBu7R84Igqi/j8xK6XkS69falBP3VfnPNIItBZW+dppfAVA7vHJr9k+uNt4wSghK
ydRnU/t15LXc7GDCOsJH3ACw6jvyeXEDQgW15eQVXr3R1JDu9P8ZoEmL1jB3l0Gw0A6JDgSsx8jP
VUtI1JkXaHQ9qqHz9J9+tE+hnEokFSQqUPEP3BfuCra5vi4K+eaoDI7UFalUS+nZete62D2w1sGL
gHYg6ObXKk1X4zaZmDuMzxFtjRq20ebon/Ptm5I5KomJPRsw5nkv2/gxqgxrVgrs7jCuTc19X9bi
PQwviruy5kie6IgpHQJDGZAULfo2Y8FhUMa/ikpRvA9B9rBb3+J51qCj4kiAw8dL1k/r677p6p8v
vb/xwN5MNaaAdBgM7nm8q50m0BfHtv1j09ojSlldbeobts5a6BN1BMjcJewVMZ98NoVQxmBvEd5H
FbpdoIld3lkejtQhMzf1w5tFxM+vfoVWTnlz87LWsfBl0iCPeyR8I5Ps3w2C1vNGkU77Oz+7RTWa
S9EhV8Vq2GYA0sVGNL0q/ipVbtv/GcgCsjNMyFytX+XyQEsrV4ZCP0nwM00GK+t6J+g3l5tYq7hR
cOxJUEflDDRvq5uBGsuxPdgXtg2W7rcSuuVg4lH+vmCymx6ulVxyqHGrljwOhDt/UCq5ZN7ZkcBS
SxbU631T2bu1OMuFi8lgWI5RBJRZCYTbUo6yzfJ+9ZIrfSPf+djAg/6XMye39ihtFZ9V5R1yROTj
KcWK4Fw6m58wECI/6pm1PO+T1A/ZWEDJtr+3Mu8pqyYEI8m23UrnjcPYC57b0MsEuSSUZMmgC6ot
nrLjnQTYmewTyf5RAfrZJuclS80bRWSXfmClb9kT/Q8zlIURvV1hzXfZAbB8Vmoa3YCHA//+NcHj
vFq5jxemkaxbGDSW8OuXtoQH7MivPu3bG86rNaGGGsJJeMf1ThCUKQAbjGnKpwAxBR1vnxcqkXfW
Zlu4Rcv1FPFIFj0IoVg9zwAq8yJH8+NApoi6tWirBKJrECKbZBMpo5x4LgmUxy+RJ9R3etCcbTcC
lZ/vMx0HP3P6+IAsBdLGgaHMRwqLH4X+fJa16oBAp5BV/1+CMyd62nbb5hESArvxSeICQWd7sIDg
WAHUN6Ni5rhbZHB02QqblIq7lOcN8hCs8S90drpu1Y8smoKJJgiZ18LyYTC5/NvDV5sQEuw1bgmK
GbnDTqti1uHzupa+0QZRQtQmRjYnYD7XhMvu1tlsnovNBUBKyhxY1hW7C1qjbNYFZnG8AV2PPUA5
vOrs5VsvKFzEirrQB9fW1k5qcxMNbWloMxiwSQNB6WJvBGcnJJE41zk3HDiL7VntzcdP88hV+vqm
3DemD3fpVFDIq5LkRzLBpUxfuZLXps/DGZy0xxZXJ7G0TG+b9AbkLEStBTR/8JVvL2wmspD0yDak
GaocNbaYvNsP6s1/1U6bZppWZeGj7H6qDVWi2WzIjVLqPBNlp9tLscphQQun4CrFDcFdX5Us2H9y
KFA0pgbCPK8fppOuZJFJOB17J1cfWSnz7kz7qEf7sM57N42Lr9imBCtFBPQYZ23e0KOuSHJLcRrv
UNLqMOZAKiHWV5AUg27ab0T0r6I032G7GkivwgNTCsYoQJMMWguRZtB68opvJ36e+AnqMdBfX4Kd
u8BGLOvMZ9eRdo9mhsEI0E1j3ceTTZMqpOPISxK/xUKZza4NjZOq4MUroWZJFMymlcegCDdz9/US
UHwUTy6OBO3rDNvDBDUzqy1Atn6vJ4H9ExyzYEj5wfbcCd3KPIWf81+F55wdt6JPmQAdwzXvb/mV
eRx/JZafD0U1lZ4dpsd+dsWVy5dUvHpCVuHQfBiDuQFB+hbagmqHOqc0+aLzHK13yTIlP7b5da4/
1pLLi61yPMd/IPYZTyXhSYnWyfysZgAxm44CROoFAkFBF5ubm2N8Jsr5GES86oJ1Gq9RI7+SdHPs
aV2C6tllJa6sqolE32UtcfSWcNSotE6Fcz0VrnqZ1gBztP1JHpiOYzK5zcr0MtEfeRjlM85mGQer
a7SLr0FDIqmc3fyUKFqqx2iHCgphyamRwfEPc6bJcYAHU/0LenZytkjCyo7wiJlPkFCb9A18CsYc
zYQKNuAHbCUl5ZfmxecAgqcf10QCgEbUUpED1KrKhTNiyv58Ygl3EWnreCpzM5qhFtIKO3hh6/vF
A2GpUtNnJveb0o6hK7EHpkpcrAi+kP380EvilS7X2ZeeZK0mdJL/B+h4nrTuAQGZAyUlqXUJWzeM
UyBnMA7iXc5gU/NKVZNEo6rROMxTTu41rxQxeo3aSu3WdMTPI8qs4HctY5AnqofzLmOLpm5eSAs8
2SdOCuCl2YZAggOsHHB6vTZY5YuAIwy6SUfBI1EQd0PHN0vN55N0Ri7miLE35EQbH9Ou+K9lcdwK
BBrONj3c9Vgcbkx5GnhUUtc2qRmeB0zYC4x2B17ZxfPBf6AOchZ7AvEy3RSk6veP3UlYlf/V2HjK
RMtbZBU069UwZRwUmkNqAZr8okMJDZuEEFp1vRUzGnErlajkyd32i0n4GPIyynM8HLeN/yso/t5h
cnZEBQw/0497h+TusdJ4qq5j/Msu6DOtGUCzSo+ApJkVDClw0vmMMeColrDcXwMkkeCBKusCg2VC
l5qL0Y9QY1q8x1irIYDFM0FPZgWAuKSYBFX7EKWhAqmYItzIlXCouQe4I2E4/2Z34h4+98TglMkG
0xGNJ7lJ4o5hVQgzl+F6juaQd/L6lddFhAZWdcy21QHhwUwpGAIazJcFg/SN2UjCLNjRvppjvJ99
+WoGl/AWmhM8cedHzmXCm4FwU3F3rocMSgeU6q7BfNEqlcha71EgSYYYeK3FIaAQobAnrj+CVMjo
ANwPd9l/wfs4rmk8V3RyyIalpTmtRSh0ZelTus5zZ9rw9eSfNKLeF0xCvrfjiVIzwTDqKH3t2XuQ
3fB6of9Dlq0sNsfJFIouOLsB35rF3xFYU6jkwyrea9sTbxq7ywnGz8KcpmrvBbxVdmemUpnv8uKs
GF3wgN8HNalE6p4xtNEyuvQiqPkoDV/wJjQ8xr/v+9YHklvsDgGfVyNaYZ11FmSPJ/k+eom8zJgy
4nknPg9SKeWtMe0rQQb+D7F7Wwl82+kv9bB9JfHJXDakv9H7l2M6iGdGdJ55HBUXiFg7ZqisDlOb
Wmf3EzdKq+fO/N+eTQTBVQH+byhiv+JXdRspPRdjTjN6i53Bt7C712oFpycG/hExbBPN1FVNjjHJ
sralYkJRcjmyFSzX1jr9iSl3cFNcxcnbdaQnOvPsUH4ypl6/J+w46V8Boixs6TzQIj0QLrN539ET
Z9gLFseVElYFHj+P8nStUkTRGeXMrC3UKPikneVnsp7/S8LiJ0YmgycuptYG5vofO9lj/OLs7wCH
duxhFwdTczs2DoqGmmTIONi/g3oppPN0kxzb5FYuK+gQ39moJWthpxIsJpJrR68R7IpkmX7n79V9
Py1pJhOnZjYAuevPpF6rBW0mkF2VvAM/s8p7rLpR69y4WfKFr4hTeXWlKYX8JbDVqLkY9pqHwsRB
pDWAUyYEmHpDjEkE8SrpECirBAMe0MbBaEyvAbpdhxgR/4s53Ym4f0VG3OiTcfeCMk4nIAjEtGn5
LX+2+2Ds6PSB64qBwaD9DfyoIG9hfdfYRBuRpwysE8NBd2SAQ3iClZQ3cNS4Ps2bGLyD7DHJIcV8
/bmlK8g8IL0q8a+Z9DjQiTmav8tIVvvJEJ7YtDMNYmZmRwVfhwVskYGgmHoWGupkNhhfhoby0eju
I2Dbu05a9+9pHyiij8P+ies1/6gcGSjQ6GXTcdGazBtvqGJCK9SCUjbh2bIKd/PvCowOn1QfJoO8
kxbAzaDKZMS2jFJxX2hiWD7NNNOxlfP/36Qq/IzK5wMbioxyXc1pPbmF9fLtROxCOCPu6VpWJCuo
C6b2cKrXOpD/8MtqXEOvP/hlfBsUsrmT9Ip8NnzIhVIAAEAFYmyFIOWh3/+F2tkZdAEGMQU1XxV7
Ouj3B5qxYukXLkXubctJiAo7fHZ3Ze0uD5VruLXdDVjCT+SA865Cw71tQGvnj8i3KBdCvJjUHqel
Kur9tPBJ/OUkuIAA3SyKsHyeF9eNARfPXLZRpRcu4TXY6K+NRTtg6bzmXy3ntN61jHR22FDifd6B
eXyUAGp4+H0icXC6xbTwGIlw4pTaRuV8OqRTFGH4skBeOZlQxp5RekAG+kFXEwYEVFRiHqdWyv0L
yqN6MmRmWXzh/MPyHGg/qu3D+3Kfs5jTuzC86ju+FtEDwAYp7o+HLZ7DZdhLAmme5jGg66WgdlPn
OlrzSsdghg/PY74rn4AXo70zyB5d/8UxGUMsZwxwxOn3dF4Ra7k4wIJnLGbeFuqoqnUcFG/o7ntJ
TN4Ss7jaCoKGciCdpWXGR58Dw6G1GpYe0sAPF+6Kd15e62wnWkILhdDN2T35+yWK1zCgRjqNFF00
ioYvVYOEKsxcsuMLhNqis6k5F9Bpo/O+qZhfPHBjSiFJ5Z24AEh9Q8NldUUEGsZ0EIepwD6QfqXw
UXBY/4nS4KM0erpKaqK8ta2+e3SamgI/SBXkLeKt3jKPsqyr40qn7CtYd/0BAoPbSNdiDy9k+KIy
3Np1OMDD/jcXaObQVE85p5ZRgREvYYjG0Po5Gsfz
`protect end_protected
