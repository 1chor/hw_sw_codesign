-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
D+mHeyqmgv5Ei8qBgbvO/CpzuV4M9rkteuGyhQUF7YvDbY4/mzg59bu11zyWg083
16rm58fKu+wa5hnCsB04or3gHC5PlGBYNwrhOIbx5ZcK4WH250qwPoq4LfuFCPBv
FdOIAJ+vTts4hQhIqTckjHrrKoQgj1/zy4acJaoeQ1E=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 49392)
`protect data_block
TYx1rGWuVTBjcGmGuWGAtnFxIuLaH6kkxNMFG63eUT788Kv+9NFS8vFl94gLF9pr
d9TCI8K633/LFMGRVOd2dsXZeoE+OwYJ4LQCO/JTA0EBFEUVauIrorMeAr6kx65I
VUbTpIlnDkAospAyVtzWL97Nfu/A+QmajwxhhPYcjK314r435PO6dYg66QdHlW4W
fIpxfuxg0owOLDkwXX0oSGfN9FFppRMllf9ykVtR21UmICcJCz54YyPApOE95sAC
ItcqxvGoyonKDZ4xuwkiC4cm0YUnEu0WlO+etsNofdsgpQ/PNu+T0US+A1EwAci8
vhRoG/1qZ2N/LNavghT1sxDk9/aU0yuJRNAmq7bHhWMp+0Vb+RBiMCjwvmnJNBmQ
nojmRIojv4+TaQRuJTN+cZnSn10zYRlaEanYfdVZV0Ukt/kL4miwHkNo7E3BoIbP
sLM2HM5J27ypkLSPsltvCSSzrmhzULlfnO+Q0kXheXq9fTYqXrvAuYLli6QQqOfq
2+qdcOA+0oPHWsKXgxk5zGn5VP8YxEBV/ZAdcQKhfMYMOJqeqls1rYNpPboUq5OD
NAS8hjKoAvbc/7VU40fKc6U1IXORcI4RpQtcanXdJs24uH7W1nn1ZhN6Gm6vfsOD
wwAlpceyRiDJ3/VRuZoa0SaKn1DQggw/HnRSI7r1dMyDMcvV8EeZ3DZ7d/mLalvC
MrwmVSQOJKVySbdjg3yfeB+hQn0byZkidkeyifnUZHrtK1sGHG0HVJwMlg5NPG4A
sB8AOYf35nMkZTkv5SsqVVxEk4zcJJG96KJZlFsH/tNJ4Jxikf1PKlTCGP6jts2A
uTYCnT7R4o72zP2a8NjEFr8mrgih2DDsEIQQ9DDLKbFtaBkQW1ikHgd2lLbpOdiL
LvKtagHooXxN1nrKdt6sg6I9Ra6eBoZox/EQSnjFt1wxXOHZflfrGv5YK6qwRbj8
fthbDco0ZGsM9Z84cRHZR9EZEESb9ku74nDDCNKrE10QuKZQolHNSFiItmnm0yUK
YNozOk8RK42N1rpRwVpYIuzCYpMJuYrOcP4G+6lWgrb9cm7/ikQbmwiS0U+d1dnW
b9qfxuI50ZL9ouIeOhdSAU1qGbNCbu8bo7OkWk38Pt6N9jvHqg5E+8qpS0qLrSl9
w/v6R6/rk8PHe/265MDLI+7QJub9RwUj09brdvplNLRLGMBDeEZtWJIcnab6YUqL
SZAObAS6WI2gUbRk550j44CcwlNTb4tgpq4ROTOs7mYN8Zdr6stKDNFfeWPN6Tjo
WCGJ7hTkbFTrJItcwWUcdFm8hbFixl6310wuBwuklcid50bk6WevUmtA14++lTMA
sSeW2oBiqkH/AVKdfGWNL8JCzBhETpD8IF0dOve+09cVAvjMhS4+fVHT5nmeFEH9
AwJDlpplZNRbPuRBmwHqrOe9h6ODrJ/v2GZnvtjqOgtjKcBKA216LJGRQqAU8XjE
dIHxu+Hn0owNCWibBCLdgNaqzqqhau0oreR7/DGlNQWBIwPPRFXa7MhxsRrufp1P
hQ48MfzZLpV1gIw7DNSUOThzVr/nH6p3tzyIh2lag3pezZBEQvwIOzWMd5qEWOoI
0A8jX4VWFDC0AlS+9OBJsqTD207WS062EoDdjCTG8Vt8t/vN4D8icJ+B9NeUzK44
eylGmMLBIUuF9vPKjibgWAZYrFV6+Ux+Qn/dQjSDWP6p7lHGLsWCbOT8b6asBk8m
LOtXNUOWDAM+5TvY5WCQAndLhmENwyAIsOmCy2me3acHaVCLCeeXlnxNemUNBBoz
M/1jTWuZlGyc2CFRk8ahGmVeGL/eM2KhGe+n8FGYa9iNiY1oBp0t8dU1Znq+Ox2/
cBw6VQdaZT03sdnDJzLa4fRLLxuyycfT6sejhP3I2/v57/NDgIb7YBrMs1H1mOQ6
ZUkYQSjMYEjc3WLS85CGTcFSzPDcElAWMT3N65bbp9hncs9XXlHgqeGTKhYq34YN
5pnYSyNbFiw6hbrYegDCBh95dfrSrK1qE8hlg9PaXf95yn8WPe2cKrp195BHG2yk
/gixi4rFQEqd86Lomiq3o3+hUyeM/ZtYcbUs1ZCF+DDuKJ5kjAZSCeBWWRzs4QeO
GwKamIphqYWeyHU2CuN7IV8GDylmnK2PTahGnqjaB7aqIXdlASrz1zITIoV1UHtZ
c5xsKpzeRBvD9isktU5hmGSsS2W8wcCo9ALW35yvQFuPDcK0ISpBOoNwDcoKLlWS
MzeBp+rNjQxdVnNeWUj3a6sTtCIWDcGpt8qvCpsQWgsHcLD8uxWzV9mNjEiAsPQD
5f2tr/5NbdIe0jstl/fgvpVFAfOHFWh7FK0s9BzKyYplwUzHgKsUVQfvvKKE2iAW
0gT9NXWgYGQ4YpMu0NmQRByiaoOYX5phyRcC+Pp5tH/INW6gA7X+KvmNDNgNExrf
1YtiIJlhYprjacJ1ScMQjnEZw9qBtbzt9n4oGihwBO3iswRGOFTeMX7IZiayr6lA
0YyQYTbcTkvbl/B+2/fIERrySseuFBmNPg8zEtpqOrCAJX8Ff6jAloaGNhwQ5P4B
BAiU+7MA+tts2XsYoXR8tT7Pcb/jr5nFKr6yGfauk0lkt8foX/TCQ6QWH83kGAUV
pReD99dO2RwcHUV6o7kRswgy6w6uoPu93csVWg1M2qDPPQ6L7doRD53HHbIU8BHV
mG3SaZ0w31tGRVfg48DmJ8AgssoAG/GlD6CDoCT+fgbHd/Ez7ZmruE2Q3C+WzeO6
VYKMCBCpGoORYhlu00eA7OOlrXRD9VE2KTRIj4Y9YeMjgg8j1gm36OFt8NOfQ776
K/6QjiwUDNkHnZOpd/DkcZh+XXhUvMSW/RO0LbCHx3Ca5zFTXgBP4KJGkGgcJKne
KVZ8cKsGvUB18OUt8NpLTnFQtmFgZCG7K3UH8vytYf5ZTEAktoQcs54QiPjn4OMP
KKL6dSPyr9xtz9AsCz2UY3AndDwwSM9wDu8XQUwmmsZFM6WCrumxYyglmfFy8LZH
VAT2W2vyxbjFTSWRiBE58YO4XhRPCtXE+IH+SDNjJJGfCzefAZVJZl9JgKRlNt9A
raHBH3KBZKm3CRvv093IslXSBPIq+AgCybHotiSEg1f0O4ZLfvgIAn46ZvXLu2gk
flXcyVpc5QYAQBaI42+eFdpg2jBbKbklL5MmGRRMdJk6vr6WpU7frx/beKBvLwoY
j+TQbJCtEqyyILSCaX78KdEweLu2A6T2pbHiYaeT4UNrjuta94uQLW+pT0QdbNJR
tHaQhKXqCUBVjApQe/ovdqOKjxcldP2WWmt+mtueL/Zcha9oQwZBJ7Mao2YVUC7j
FRK10ixekTDCERPh6/W3NqCSt4Z4MlF55SYBRFX0YC2lRohG2aLcTf5XAFS+czpt
44tBDpUb+LwsLYkjoykFiB74dy/rzntyqPl47p7XYfmJ597TneqFuCGx5H/zjlQw
hNxUu1e73f2TlPSlHvo28vQ5cYS9kGhsIv3IhBROA2RF+hnYP8f85PuOICZC8FFI
G0ZkcAkqSD8PuFsnH/xfjyoibe5yTmOSN0b2Sgsk84Wi+wl6DPUeH0JpLn7eKWGZ
V5LVE0WqABpIlvFqpsCIC92myEUOITPbbO9lWxXqYmI4BN2Mni8IvMEzO2LOHDKX
mdtk9Cuaqj1vCW1W0ufJySbrNAGRbOd2fmUmgav+xV38OUyePZEZ2RNy11+4JoP/
Bgd6ABdsW/utxylp+LULgW+g/zkpa6cXUIBr4m7rxdoD3c00QxePN8Se5xvDFnLm
aG3XN/DgNnCwwHGJJIpzdVZiEv3tos13KkFlRqnfjvwtC97OCPkzucJTSi8ZBehL
b+BIrJWkYfF0D2lHNfzTuDt6GB83unDXr8xscjoYFdWp5tPGu1jCdtI78A9LlWf3
pNYQC6cQWjLVbVr1BahI8+vNJYrUOhuvkVT5b6F03j9Cjidn6Ap9kwyXojWFWmez
1I64NW3+4hAdDUDmESk3UAID4yQTMzVpGF39f+wbl10/P4nRHR3oHzumpTn87PD5
1BKxW0RG6r7rZ47nilA17QhnX+inl2z18UDRI4cuq5wOaVT2Kfj9FaAL/L2Dx9Fi
BHFbHiDOsHFn/UxU0yAZe2s7xajrYAf2lso9YHc+nRPIGCkyPhynDssM8McT5SNz
1rfzWFgiNaqstXV3HIBwxyjoM007I72otk960bZK++8hk8vgRcgJEfLYiBL91S2Q
gcZYmhgT3f0/UbW9ykVg7zAPJEz2fMTUusiiP14S1JGhGw5ULYs3zTdonvH41o6g
XwPPCmNWDpBuxzDNgopslnfo5VOrandYHQgDAWFdXwODQtvTI7Yt+0k75dEPUosy
tGvzozK09TMrUNpYCzrKHuTMDBq2zqmqLCD6k1kIloOxFkAp9IphFA3qXvQbNCQZ
emnF/5pAR+vXib32oVzBeZNtbcU4UPeJtZ0Npdg1aqJxJXXp1qpC6wPbAotUzrlb
r/o5QyzZ2d8rEakdHNR/GOKX2tVmkB1/V3vyFNRDs9BdJD1NpKfzD6MO3Qhb6shJ
sm5mNNFxBqmoiBrxj+0y1UNTiGOLhDXAgqlph949fyYKXyVhXVN8OJEdpgYyXFXm
ZBUPMw9Kth0kT5pNO3zxCBdRTWUXLACwmZVE06hnj+PmLFUcsdkwmsCJpUeYSyWL
+eIiUH7VdY9rbaYB481MehlIbsjN5xjTNJ8QWIUAY7lJfZ7r8mr7YagkFQ26Ly8q
w2/+ceoou2T1PI9FYqACGcbLPUTg8Rf7agi0Y4xp/ocpnXYuwr0GIRUSgxF2R78o
p30jYczOuHtWPnEr+ct+ruEINMsEv1cl5hmf+K/R7/2R0pByqnSTzcBQQ5aYSl41
gkq6R1BkT8AJDTKbze0wMc/8rqg95D2JnBp6TvKsgXCOaKEZXO04vXITPdVK5c6G
E3rHKRQBrhHeWZkKd1nUhNJKLRmU1aU9bO8iF8e2g4837dIiacvKSp4XjMi1aQdv
zeZ4367zuy3MDO7tFo+wPfwYKN5AflmIaGGns3DOYSNgl+ptDYe2ladiw8Zcq08M
0HVXycJlc6sBFdH2nCz82u6D83qUifq82z8sU4i/g+eW6TwZCz1kX9VnFHxhyWAI
0cU8ahHLNzebNRkacHFUaDJW01lXE9nMAvEXqHvdhtpmXWq6yM1BgFt5f6BJIAH8
/dJCMl6P5/SCSP3Wg87gY/nXmNqfQ7qzVZWFsLvwx8npGih8Z29gz2NprBVzBF0j
wmDPguQYMeEBLgTjqFkeTspRbvXC8taJb3fe7QVuJw0qwg4H7njqthis7MAMQlrV
wQHEdcbilLcSJj9Li8616yVOJS2NTALhlaBbkAgrqQw9JJKJhw5SAVCiS6Ojx+Dj
raqTaQp1mLVRF59rn/+nZFlq8SHTnm+EX/phkS1IGmeiAJoUYD5bY+uB2Mvpjkkj
B1W1ySZA3vf4+8heFCHD6LV72klBW6xcQaBFuUEqoy2G/wR8Co9ZCXMX5buwwK1Y
jy2HIE19P2IGpLqQ1Qo/1spSRGuJ6pIkWItmfchvi5rlr6wquK/BAmCav8hh+uhG
i7T2AjyrYd1vKNK5y3r/vYJ4AjKWt45qvCzue+d8Zixs2yImWeM842fM+7W6mJKh
bNAFpOgHtv6LB5dWpXVeqNydRLpKh1iOg3QXNFqZTJjFND+JtbS8VAlvyqXYnuQx
H71ZC3dd4YXacMYkdiSyLPemp+PuWwQsNe9GNvUnXQn45uosIMRttym/gRsUjpuK
SqReG9TjFEReOLBO7MvhaSWpWbU9TCbWvNY9uqp4YzwLfyRfGBdkxm13Y3d60+sx
EmidYZtQHNqGILqXKTi5DzAy0JMH/SElBelI7oDd32vbedZKkovHulxNeJPIoUQe
f/9vfwob+JxDZFzAfYaBBciMSGHAPGvpodxsZvhT4ZnudKC68/yORFxAhiPs604q
vUHA4dP8nOZ8PVPJnhRtluIr/h3dh45MoKuCJnUqyPiyRZuBsnXIDxuRl5wfp2tQ
VKYtO/s2li5eCReU8PA0hPzsAJ2DTF/awu6K/QfrulrXRaOI/PiYTsxuVTAi9ohS
g9N1q5E6WmYoIL2ZCPZy28GqOE5WYKEaeTbyHNEJrr1S6ULoEvzxg0FixrI86Sp6
oRX2pyVOGUudGF9+/sfPcgnhUdOyRpi2ZmxJ0p6iONKPNBmEAr1VMtd+omRRq77W
mPf82Vcv4G+xlSlDy0OARhC9aFoBPDcCQkMxOEOJKy17sQvQrxb0fvE8BAKiqJ0D
COypUjnFx4UMoUb8d/ELIWVHNC59cfVE8gd3RRVX0B+iXqdzY77FYHERnk42j0Aw
CFbts2J2vYgM61PwHcPsvACPVDIojFE5BS09hJu99YY1jfvBNibIbFzDhaxZ8mG5
L42jpT+Gv7UVqI+IDz5qO3DzLviNLBQnBT0YwwqKcYsbUwwbWeQwEnNvisfTpU1V
0lU2tFVowkXlVnammEsPc4cUroetLXeBvXuw+SKHe+SYpfv5331Velrz4AFoZNyd
UOKTL69IkVWcBs1cofA5/i4WhY3X9rYt6CjXpa2t4DFGs0Fs+b6Bjx5lxNOUmsKB
19KZYps7LXd2LscGE3FhG7wRLWmZjZ75k0pvNJ20oh6/RqFtgp/kqQWkmBDmHd06
v08H2S0pZhzaul7T6kcnmh4vUexVQK65O2oDPgbEQVYQH3eFh8wF3fLaKITzAG+q
IgRzxYaUxPT0yFdU8h4i84S2zLSkDpJAvgVF+RkAC1v2/Pox6Wg9rOEJsfURKJ5Y
MbWY6q2ShwyVhRaLourzhnFdHglVnpBy+VENsvrxH1VRA1XIFAjYlXIqbFlL4pEd
Acs6E/Eb994sel7w5/rJx4vH9zP/HYckswBlLoS1lMuiGgV5rSInOzTeZuUH5ndD
YMgjnaRlQZipppGZF7HCBcKbLjgD8VHKe+f6mKZYuy+mIECXQdX6/1d9431MWK51
byrs6mTUpeQwF2SFZcA1Ymez2nruS1bJnw1h5aYV5+SDd2bmx0x4A8AIhBRO1jW+
8iMN1bwrBgtrMMhBmWi3wjksl+YrI4e/IN8naRm0xKWm9Q7SEs7nie6KvFuZ3eBs
U3xH3sT9pmFBCedBjPsXKzFoe+CaO1MFoMkn2RzbCuc+SCo5ydx9hB2/40sS6dQu
Ap2yV7bHX4Eb4qY/HXg/9JmHkzYR6SH681sP5diQCxrFmtBMjh/nFTaQ7ZiHkEjM
UyvDwIaXhJDuy8sAa6t2TUGoJxvqvmyHhWTzrR0UPfVPq6D7Xx/ZKKWFNJSLX5OX
74UG9qVfWP1opVz0PgrkyLSKkgMAe0D8n1TmrucB54UzbZ/if+EbpjzJoUaG8+4m
zO47xTORW0aq6pXlK+oWXxpIFI+b+N+A4fFDNR4eVpm2fslHwFcCJknSFi9pgztA
6Z6WPwjb5ZVtpRtY5bJc20M5p8iWVxT0+bGRuBifrBAVivLO0e+Xc3QBQe+ilJvn
Pqp20A+KiY97Tb0o/KN+FrKOncuTZRvS6gL93A67aH3E0VsCHOUC2zLhQugkzhMy
+FOoDJHw7WFAwc7hpUEhp1reSh/idHMhkNr2VJ9NhbmarPKzpvaU3Zog9M0a3k+0
N5No6PYfejc/DzTnm/nMSL29Zv3bP2EAwqlWrLhr55AiKpy8Iuc834EzguEZBWnW
mgzlXUUHuBholz9jo+A7T4xbMtE7mJd4k+uu9VvTjj0pTiJbAbl2a/F/4bnN4aMg
9Odro7Y04rOxdqI2RTfyLiPA5Eug7yOThcnJxMjDu51IqKaNfyUIhgbIw+9LO0M7
oALe5Mf1F4dmcnX0cPGxEIOSPnFnGG7i03eNxWLdXG+evOJhtibf8XFL8WrsHSKJ
0d0sI+5rs+ZqME+OxoQvXc0exY/s7QEmjPWzcT2m6uHTIrEsS9CSc97DQwuv9zbG
ox4I/BsCYIJXAA0wvWHSq1uz1fAiNButqmbRdI6AZe/jeEUtfvhxpBzTmlDvVgJt
oNoNJzUj+kXjBbNt7V61hdb/sYqnWq841lrObaZqUlr9JmTUZsVKYU8Ge1DZ0eDo
ct5XbSL9LhwTUdkxtkEFkJOZ7bvOGqhgJJbdnLTHuH4gNlymxxGervJSdVuXxsXF
EhInBt6AR0M6t3IeYD4xWslqLkF5vCjMe6edYRBHED6UM3uuCAWFQuI+eSLitug7
C1YZ9kdlfXtVFvoc5UL8e7MKrJnmsPrVj35rlNcu0arGiCXer1I/8SYGxRKlJlnU
z6KsGMqJ5AQXoTnKdXyFE+yOYw4OoP4QhtrnONJer6kosSguMtDwUGx787frOZfl
JYca+5ox8JqHLsCwEz7qx9JsaJLsqpEBCzksOEgkhLzmyIqCC30mQwy86xelqWQN
kthXmkHZKWQc29ffM7SwdxC0J0UV0WPhrif0qcUZ7TK1nhC5faT8kHIx6jABLdHc
WTzktRimpmdW56yHublUIg/m3RptGU5xV5wRc4NWJZGRZIP1Dzdc4zKcPVgfHJB8
ZmsDiOZEdNuwakSqwqMKf3N5SO969gTM+wG5ai74aLGY0BZngYVcwpphMD3rhj5w
6K/SPdaQAJBuH3IqpTd3nFj7iF83SPrOtn04gcW1PocuPScVSSE/FPRu8Il83go1
jAJQhJlUBLUD9E3nFZWmemLsIQ2p+g541AoCeYjZFZaI2Q1vfiBDVhrhYciA5NFq
Kz4B2WezVuaPKARtSXuqtrPvR4JxuzZLU/w2wlI5qXQopMYQWw6QGHdxFp4Ofh3O
P7tEj47Z87dK6phDv9noliODvjwKIaz4M5xocuCh6X20TbbitfgZ+qoeAX/fCDrq
NP2spPzwWpVWQMEYE0pDZxQmdUsAOVzVbW5gnmua94zuSHAQFUa/kyxEja9pHFeq
Rfoa8Y1seBALmX+w9qqIE/BmXHr+6b72euSy1Z95Euc1mAQQdoEVjtadGajxjW0M
XYWOvxQesw0aHgd2mXoV3KmHG/j/G3/Hv2lKd7e7MVWcY1ZsUW1piwjpPTE65mMq
Bt5aO2u96DXNmAytopi5LNX9RoW8BBpRX1GKFUB8GqwsnPqvKYJFJCmiKGxILsbO
bnDFgock9ufuyb42ntGB6uW9GgzFeOjiFanoGFe2dlHv8d8v2+EbZddGuUhCjybC
85K9786RzrV3Ci3pusj2QbumSNCERpeHiSMBkrbp/pD3Fu0x7B3rbYi0YJghJAGK
XhQCCT6upHizQMrCBOTMpaIbq/trWfyHfy3PfTm8PG/TY9GOQZm5qdUl512gRm97
0d6sdsb5244vnWw1QIvg+qSKI2Zz+bRcLPMB4k4nynzP610tyHKSqKGWQjW/f10S
T92IwDpg8uGS1J9+efimoRqCT4WJd5hbTmNTNRGRW8yMoqxN6pNy0ITMhgSzNpzP
oHk4u5OWDBHFm9PTB5NKzLBjK5zZqlHLSOKvwvldnzmcZAseFjtBt4N76ZFma/lK
6E8uZOhcKLMsQegJ3Kax5zQOcjKwuQtZQ9/dE6YoCJx1efnHGPM2VBC/SPeFEFJQ
kZ6b7WuUejsU4zxST+grftPDgatykLPOodJvPp589b1A8pGwxMEWzlHQjGBVxOLB
nnBkIVIKemKP1raJELwiHLjXAFSIh7M+Q0cq8B+IiIeWfWlC1tAURz8m1mBQw1G9
rrtPLe/6lKoiwxDnb2NZNz9LwXGvcsjhRsfpbKzMDTZvVrRNtxKDy4XupAfD0ymg
GrnxJtiXD/Y9dxALdPICVSe6LLd/l/47uQh+dvTKS1ywZHs1RrOganMuRC+wUt9w
xVKVgHl05rD243v0NdiU9DfrbSbEB9ORaKEs9+MRPs45MBcPgui80GWrGzBcMsap
u5yBJQxRQdYxjtYSyizWBGDXuV62b4jvsoBJ4g32mdOEE0kHon+XWCgOT5T7OmHX
Hpt/8ylboA9pQ+GSpyD8CgdtmOGMe/7DLJQtItM+nY6d0Azj9JPW/UjdFGP1WII9
lWVSaUNf3FN1M+hXyrrhSnlZRz/sUlltAQ+CwRY0UwLt05J9JOCk7ZZNZ1pjFXsc
MgdgYuV4amCEJHkHjr6W4YGn5z0DdRqXvB4K9ob2sEY0QlTfImpqd2ueiXzEvs7d
KDi5NmAE6fRBZuP/b+IkeNgUiisHrMq3PCJpzsMRSp7bA3M7nquM6i2hp9P2za1y
5M2oG+GXzL3X08JBZOZ0ZvYY6f3ohiZKnFLV4xI5lji2lmYzBCqM6LUH54Wyyl71
S0KDNuf4IQdFVZDdpxM2KDIzxWP1vdm+QAajahfl/2NFCIfqmCG42pmSr1go+50O
7aQ/PLQz10vU3C6FN9fKVSxczOTIlXTavxuxcy5bSKUYMOsKitlKUBVpR535oGOE
7KfyCkNuqEfMFT4QByA0zNaao7PV0ZCEgxZT/j0eqCztjTTb1cRX3eFiCiOaue9+
RZtyUd9U9f8GOKolGtTd7OYkiMk5rav0rJUUFOr7Xb0jOCepCjeXBHOAGg5jGTNz
lzzI7ifAELjd/VjFCsoGvn3dBWGjuy20GWk+Oauev5VO4Ltmn+ttdmtQSodMJuvX
23AV6kOvzLGP2AZ2RaoX8s0jncNZU5oAERcZMldiDQV1AlsyHsHh/YAj5rug4pJ1
gm0nCLp+RwlkHOUNye8HhxyHQWhG/Fe56NJqE82bV6BOUQLo7Vt02WEcMf6Tr7Ul
TGMCd+MZS70RbB4Ha+e+vD5zE8BENmLk4ivDdLw3+Sm60kcoS0hkFbPlOFFnU3Ze
Gx/wkXuDk65cpfoII89b6UeiorFffVNAFfXsBNkPVHdA2Kjq17D0qlnP05puwMMm
2+8WPkH2gSE0NCcmH8RZA9CeTgfnIsXkWfCxlIKD8Qp91fJg9NYbuVKuA7xiDUWW
XVsmLUqXcC672WOeioOCbYw2KYlrlJys5mRe+22KyV7Fzj5jn0t9o84K5J/9XZLh
zRTnGR/B0ZPlXTiNda4z9wDopSX5wkzKO5Yu/xZ7zia7+THkmqMO6CCD2hi3WWAA
ZDeYwu6TzXcCM0HMsqr5WgN+y7lo6PAH2QAC9aNKJi3n8MBNqp6qiPKVF2YXQ5lH
x3ZkZnau10BABklUWmSJCSMKtIuYcA+p+USVdqakIC7mp6aCwlwD7On/6HbZyhQ+
ruLTQHwhLbcWJkps8Bq/E4CDy5vAv55S7JjwSUqxP6ajN9ah11feY4VqXAWvqjvZ
3d60F9FlIi6dbKcSXniLVQZKHtHuHvCQ1NK6xnlhRnSW3uwPILrX70wksMezRGiY
BPaAFPbdKZQdqBLrghtN+DV2uAmCTMMKbBvKPYNLZ716SbvhACesrKNqhJwApMFK
8qt2vRW7eB7Z5PNzSAE5GXyS2LkCF259ej910l+VADZJ2jn5B9qqfHGCPCD68Bcd
CgTvU8K8MzYIYtgOf3+RM6gPwYEuvicgsDe+ClAMDNIjzlUTMUWsZ6DkJQoL8ngP
6gZtKCaLDggRVZeP36RPthhjFIjUoIXNBSlL/tdbke4DRcfi9+G15dCtv+zPiUfn
YZceQs32WZJfPs1mO376gcLgc8gBwGb/Ko++yIpmZ2e5Yox61AurGusC9stJ5fB5
Jzx2IPUoAZfKv/pcuwN7fwhoBgzOSR+F8JeF9pk0SxuUhsLI0uA8n5V8NzlGapfW
DxH5RNgQyaeytg8CQngGJAlnxjUGjTmeKb5sUepdPsJehjLlBD0DFsAwyZl9Gr+x
X13Qlz1w6SbAxtCmhBJ3/p4x6TScg6s1ms8OIPdA4v0sUV5TVeQh6ynVFcSa40UA
PEPg7XravnThNIjc1/aEDt89Ev88spajOIALFOEvjNaGe22qvtWUWCUnASxuxZB+
HficQsg4ULwjl+3IGD5ruXlKJ8tokEj16YM0t2bmWIQYr7J6GhOreM/g0QtgIDxy
a8LODTv9Y3/H6nICzhkxb8d25pTp60F0khoLAIgDrXA+DWLpeK1HtujgawZzs4XM
byL8RfdDb8m87wSmJaKh5xWLdECGMgjPNcoKE1i7YpZaOn5ArpsaTxb94mDqPTvk
XeLXWAgI6YPRvan/ssfxfnX+DTrAl581xN6U738AIBtaM3SRz2FiORBaZ0koFfxp
UmxJNrmxSuZL8cuqJoeYScB88P3MjBb+aAAHtSOMBsau7bY6V4GdCLMU52lep4d5
yCfkcTdVGbjBpMZmvPxNuBV89IYu+C5IjLgUUnkUhNhgdh/+eZrH3sx1c6v+Hy0u
/G2iZ/tWxoLXveN/eluHYxV4briiycyL0W9oiUqqTp1ZK27aizp32vsgq9shJZ9/
AsJXm5z4dZqtK7v5ukIQ2X6Nlx0eqhnZYLeMiva3PO+cEi/2ibs5R3Eb1AyeFu6A
6ylWVKH+z/k3Ij8RCw/p1Rkk+OjWEoaFR4Am5LqN5RWpApZSZhmdcn3EvV7xpWPP
F/H23nWFsyr//aKKD62Jrde9w/+TS4bKjjfHgbJuJBIjmWpFRXf/kB4AdWB/75Dv
7syNpM+lrQp0b0GMRZ+6/GudKf/HUS2+7UCfUqyqWbFxnUvUol0AIx7tYXKnZVIR
LkEAahTQXWxm9qmbmgmjDUteCQWGgYgSxwJYzJNgYMkIfxRkjgdPAWoqg79pk0pU
nJVS1+ZuPpCvEcJP6lOPea/pJK6NA5WYsn3921mpo5Pc8y32jfzlNvumsM7Wfc68
rrnCVeuTOrm6c3TWpj+HzXGpR3zccQlckw+YW5viq4YbcHlRFu4nnxZ2gNP4JHZu
BqkSyoeYD9AhqTyhZIr4P41t1q4PAdg6XlCk+DadlQHGw+Dr9IhwnbaY8/1JVaNl
Yi9XDQBZRIeVpu6yu4rZjHwHv3umx2c1KrPcbpIF8sguk80sNVq00zsU6E3EpZXw
K3k0TNv2Y5C+pQWBvabPQjFy1J4/9YeVzTI0VD/kubDQCLNM1gD4p1tidnDdRAvk
NNC5UkAU8kUzvKM0F5+Q/QNJVeN+agPDzloGpDZZHbwldB7JijsXH94Ryc0UDVRX
Q8yRKQljnxombYWDgD34h8ItIzqiCg98cmJ/35bz0iQQzbkDHdVO0FCk8ZtYeS17
YqoYvhl2cCEpMZdIkfS09kUmbPI2HGktqexiB4QKEtvTtH2+D7gtlkYO//nPAqoj
WpqwcCAHNaHIvt9ij0g0QD3LmqJKe03UY5aDU5RM114IO7murca1ITd2NIeXL9uK
HKrsqdRnEkw71aIkfJxVpJN5UM1B/RoZxwy4kwHfEdiOizLmjgELjJJGulKIxpIY
cAx7//NFV/KI3ueLWZVQ3hMzw+DkQkMOKHzHEhxOyuCmtZq3oJTYUaSTkT3HKgq+
7wGa/X4nvx67oejWhgEXD5n1UL6RVzRHfmLwXWQmOZUBJRTdIn2PkGD1ZqVed7Df
3A1oiK+cY7dUcxEWyMxOWFs2+UociJ9qzGvrqFmh8JtkWfluH3eu/i9NZfSbsSc0
VDzAhYWxwDJVOWRF/gfh36xea/q7bnhlMhtXUnKHE1RV3n5R/jA3lL3IzmBZOVJ9
saNf5ufPIWe3/Pvy/mYCL88P0PLhMJUEPKYjk4+F/ecnhbNQa0OfpUsC7f5qXZua
vMPHxYb4ZcmZp0fsV7QdgO0IJ3vWc3TqfX1uhlbexzhvKJojTKxcjsyqJR2EJ4Bj
5rPviIFNQUAPmVJgYhW8RCvQnqUlX612yuCW0kwgRCnbs2uYnH9DRYQI4BptmC1F
39JrahkXw9l03A6GmBamsbsyReiY5pR2MAiTLKH1i5CNK4gmKncu4zgBbLcLurVp
gzfaMIRkNG+linGPyXM8UMh/9jHyImZasmJCPglsE0LFGo4pyjpAEGnB7sWBj5/y
e0iGUYMUR/Glzk4ImgOHHrA6N75FGHpotWPhFS7TwI8uHZK8wHjCoPNy63UrYo7k
GdIZDpzOQ2GkbMN5xmVnbgOp6Rh6ZTsp6mtvKYsKk8MqmeeX5EYzRz6bqkYOP+x/
tfbvOClaXYUGfReIKxhV3/MKTAHedQgP/28Zw7M/4XIXR/b4f+IG4gfP7bHsid/K
hq/W0Idg5iNm4ixkKxBI/tyvGO9z0idRJV3dxTBuzZlGG5mNkpu0MieSa0h2LAFH
VrKlfnAArI0lhfaLeBUmOXLb94qj5aYYndPlA0zf23BEChmvOqwUy//M3uSZ3NTI
F9RCbBH0LKwCtoAI/hUy9FhBRoJ57U5/5oaFUwEiUE4zdIvze2i0oBW3bMIYcu/1
+wXr3M4+9E/twL76fRmIsiIQQqLSvKH8MtcA81ddTlzqBWFMExG0N9bPQULG4Zg5
t7nfGE0526+rRkGvDpV6G2oxJzj71Ka8ikaKSkVVhlzqNt5r/DKIW6iuNKgFmFwR
78J6YQ0ZZcDWG5IdRbnBThXPUK4KMwFfWabrjDZ0YuHksYjrlk3zFTzBaVNINEcT
j8Hz0IR6TWPqVTQ23nHhaKR6tFmUzmmKMlBtYCHEZ7VLYoTu2BmUHlRn9VQRvFEJ
sb8jOYu/grHwU7ervtBqH2CS+4bB+20YBpQ99AuybQ7VRqI/WuT4OqusKKp064QN
bwzj9bGdYxjm0jeKKh4YNQIqaIIr0w2ZRqcURrlDEDSGQMLCp3mbdAfZT8uPBNIm
FlyQKd/RWhpMuxx41JMCbOwWXVmvg+5gb3qcH6CpvRGqf7HQYdIIDZb+EJAk9poy
cN9tx0ylk5HYEWvQMXdPpPO7/hcu/qtLyMPBPqy4CwLlNl1f/ThgWtFDwLHBblJM
NtwcAmUh81SHyOIJ30kCpjq+O0fl5EIY2rkuQ5+fMg9y3Encj2HyZ3vS88g8cAOp
JqIDpyb4UocLLTda2tOmi0z/+p0kQr9W9rETNnf85qC1X772Ad/qaAKzxl8URjix
P/6XxUYxupmZrSNLG9KhLhl5k4QndePvPXRR5HV3/s1WIMTOBFCb2/xi2QQfynHj
aUBhmzdzac/pn2eTJYNjKPVFYSYLCkXGOqhZM/p1+oQu06Goz1QFGXeYJpC0tXQq
3tiL4BCyWawiX1MetcCqbILDl9chfefwZWEQ77hc/JGkb/xw0FrsvBWDHQkcLIEF
UIpp22jB9ORMteXNItxRdNHPiCF7+joGZdO6RetbAX2FVxy6nTY1ozWMS4Tg2oU6
J+JQzC0+ojfU76jaHvzpScMsXJ6u4MusTN5bkpIKVncSg9lZrnFqkM5blErLAGdk
xZiiwVP3UMLn2+p9kaDqD+h7lmD0v87AeYHpMMA9JPlEZ9wUD1eanIjMJjVWUThA
6TVi2Rlz8vahkd6QqpG+k+plY04zbAJeAFYZhQSqCqkbkvcV88qhcnIi7vjG1Rex
2mh+BdDfjY3fQ2nWbNmZc1rUzKujvQVXclUihCrDnoZRmy2s1SboYhMDEOubW3GP
/GU+IPx1bO4QCjV6jgtjsgYyyCn+XZia2cIzjHeVrUeGb4M1el9VrGcm4jkgX+bI
UXckuXB9LcPs0b2H+Tqhv8EoYamUxF1i76bFX2SvH06LvPW64xcfkRCgp8/IiaKW
HCUwsrnaIMyd1+ra7+s/rOc4Xu9wu1R2mnAUWYBlzPJxFClA3NOGloGwF+OEufPA
/Y1GCIIcFi6DqdRgCXzisB2mxauOpxbiwZ/EHYkyWgVIim58eTH03k1tRTMNlTDz
yP2vePc72fUiTK79bPVbh0c/9soi4/BdRPfr/Io0QWRy2Cq31AEEifpoWKA0aWho
7plje3RBEBHabGVITz//h4IEwmiCZAtAg+hDFEbY9AptqJ0O/uu5ShuhdAGWObnn
FoGzk5nWaq398wOUyP1XJe/S01y6eU2nBxtIGMRqRPpg/7bHv47bAo688ylnmG/k
D+J762OQ6hgngHSG2ouLRqusDxDdBcOyU813jmZF7R22mNrH/QDt3RXeFhky8zFa
xeRiEI2IRoNa4sToVlJGmiUUzK6rOSFDMeHxCZ9LICZXJOgVa2U90dN1A/Z0sR30
8qUh7HBP5p8O4pzua8MNF4VjfCSX0ZozpF+x+2IBGuvDLyGuslKdTFL+9+eUyfqA
+y2q0wIt9I7q2wwWfS+Cws+e4DUeakzxKfBd2HCD4C+P7gu4mqbKCX3mOtSSzUe/
lHLJqM2fVXmLB6zBUvvOXxj+DlwfZ3Ft1KrCxWEQTyQ+EFp1pB5o644kE+5FbcCU
Z8NxeQjOP7+653aCeimdg6NyFjLhKGHUdsqGuzmXItHeCox6jE0izMggXjWVlrIi
ijhztZb4NnXte32OEVyAjDDYnhPQ7HFzSvusl42yJ0IihquJ5rr5foO2TjBYsvb0
ciAKBJ1AWAzvOieepLxIKKfmJoX89g6HdN5sjCdHALtWs7EGDR/FLv7/Xz5Osxi5
WTiTmycAAVMSlWiREj9M5NXZ+3Cyy/f8E8v+31I5fuyJhit9TBTq5Hrd5XGx0gSF
tWegzxFwT8szszE8JkUL9Q/iayM0aSziX/qXrFlOARUU/PSFF5jKrugWPH7GyRAM
EaBRtoMzUxMXK7gCAkZXsQdXHb8odxUfsvOMji+UYDjeTisFOPU/qM72qJ2ZafCK
Jad8peVPfJbofXe7SCllafaYZ+jcw99ozats0bxr/oQhaXf0LuLvvJIMGRRNlzKa
VMttViEG1zUSXFO0IdoXwmJu2pTJNhlrLwK9XbuGRF2T0PgGODsNVQVkGsakYqLy
/FFkz8uD3d1Ar5yb6dKzLPSEa2bfq5nR77PgXk74mOOKK4s/5+ejLa6429UVfK7K
/wxTA/hYNM5Q9dxWTDqw72qes7mUstMzgnOAzoEphsJeZIyLHb4DdmaVqRlgCi3A
GesFOBn75XRap3E/T8u5DTbGMHBjdNu4vVCR8j98+oiUeA6eWnpsRwXf4o8QAD5d
DHcM53CgThw6f/UfPllJamgLjjoNSMA+8jxCC0fm0CL7L7EuiAQPUfzFfVi2mTy+
P5HUpubHU+L5XR6x23QmPRvv90Vl9oT8liFcW2sDao7nATTPTu8YV11oM9zjse2Z
VKTRVzR3tMWVo23upkcmYCAnPR71b/Y435TdLbfsKFMQ3VCYtOLZ5Ee4WVTqcWv+
WIwKG/oX2bw7etaAK+ZMtMHuiyiw7g+KLUe/n8Wa67CKFg+lELZRfUM2mrEu8Sgn
PBcmxPo83KJUkdH2qWhMoP/TiUQEC1mp0E/DvufpBSaPBDV57S3KZ2CTJNMeMpQ9
9wR8gIirXR25Wy9G6kTJY/S0QFf2I24gw3Ju3onuHEPb0tIIGbQnH20bOeXyf1/A
mH6iW8CfF2H7erAuuD88xCllB8rcY/uGoz0/F4ZZZGwumHguVUeTBFFE2B/uUNrs
5l7XmRY4EZQKmLzQVeIVhyavv/1ocAaNWol2q4YAkPRaF6Nc9IoG9sj8cjbuVwcK
aLoWROvGWjgebvEh8I8AgTN0S2t5g2RloKXvEsFfefbxmJOhhVamNwdUvO4LlRHL
KP7RaT4sx/KA6SNkMS5KnzAGHe31r5aTDVG56G633i5UYZHlNXUu7UF6dsf0R52s
pJ1uZ1Gfgna2y82yStpfcPb1iK2+MYrIAldIu600Ecvj6FyX5EqOzQU/wu0HFOlZ
96MO53oqqhBvYs1JX/EW4llnU7+vZcTeqB1OPeSEZDapgYkLpgGbCNta3aj+s2NI
ZyX9X+MJz1b9Grtf6EkVIouoYKw1Phx1cPOO8e0Y2/aBcnbEVFiZwFRKYitUY+aj
uIVc2I8FqxhzIV0l24vCWLIluX2Y6px5Eq1SOEUWSI2oYK1uKvfHZJn1oBBmKUGw
1AS/EyxPe8hvm7ZhveNgRUIEjRPS08XEkk2HCwFwbA4eQQL1FZfiYvQLNIO8V4Si
/edEddhwXKNABUHZJFyruOJ32KsPO9pxlVGDL7j+Gw8quu2cZGXl0RF3er+NCSXn
6i1T+i1lb9nteyDFS25Or6KOMZBNmUAKaC8pp+UCUBluVtELNI3+NT9HdMd8gQFD
WgSUYlwoidUDjx1mEeB41vPWY+5kxWwN2jfGsChzfgfIv/Dnw/0+JBn1GwsbJwV0
Q86WQTaZm+H8PzRymSyvsg1o77FfCt//5U92atDxiX7UVw8Yplg5OV2VvHkgsgQa
sOeOKVAVX51ZqqcozvffqPhJZmHmoe32J8IIxDdKTaI+CyOFoJC+Zn4/EZeZmTi+
Y7xH70gl6vbyq1LStn2ALBZK3wYdcFk/3aFBhU1MFUk1gF+X2wfqcpBI+nHrATDY
2zAsIUpbI5VnBV2b34EGSOymRob4z5c91HSEYRWPdne8BIPDP8DlLUPUAsdrwPPf
yNz5od7hkLE3j7jPIY8emeQnyC6nsG504QLW0t8kixWik5ViaH/WXarWAEJb3rYe
6zjgQQqVpPRwMO+y1lAvroITo0VxDHi2AOPV+elVE3uWlj0mINQfzohpY51b6gjj
xkogjH9W3F22aI6d7rlcjF7qnOWxgAvuKi5z99bKR+biqXRW+jdKhFdyVmoWvog+
wwO8DMc+6x7cZSrKtNk6V5u0/B6W127kkKvp4306R6cG/HRao3nHqyKaGBXbz5yT
tzoCf1RAiKAWooSsBc5TlWjcRP4jePR1chC3b4EcRYuZmowD77TO7Pm+BcpRruym
2waZcOxfrG4A0xSm2XXuadTb9xk8EWJxmFvad+ak+85czbcdqPlq2hK3YO48iTwF
ryE9PDRefEKBKTmsdRGeiAQOaUwm547ngvS9woVrdmSmynCmS6YiK9yF0TEANyJb
3uB2JUynW11c5gG02+HKgFD+kdtaLf592YbPRZHlHv/qU7qmg3gjMv05Ku7t07OY
GS0DFAsrg29YH2rTUEMtU+vVDcPMKmUWdYDNXe95RNWYs+vWsERhafYGh3zReLfk
w89/dWWvdbbtPDpB3YfOFhEK2kFM2JulvvsD53frkPPGbyGAuot52T5vgd/pP8L5
Om+Q05bzQeZLYiKcvXFO49F3rYxUcCaIPIbcmk+47yCLEw4xMB6NcVzXdLznwIIw
mg227+1QYOm5vH4P5Zj/iSkgMLR57hW871EBzhyCC2AZ7A1TPj8hEgI10FhT+KHV
bfXfdR9oYTViFfJ+URJPN1Xcv53hU/Tz1ecPrbAd+Bu4qYHECOzLr3qAG2mdMg4J
sGStcOCImVGqDUW7fHRkqwJzjDK8DMAQpu3XpUEiNrBJFNo+4F/06OjZesaNzyyM
BkGCVP6wVVaqw4i5QgPc/7uRtG14cWzuncdMhMgcGoIn4yBCndJey1bHYtlzZ/15
6/7IkP5UKIznr27f/TOHrB1PfBvY5Y+tJy4OwccocXUQ9J60Q8rpVXAF92HmYDfd
Tg+iFscgeCSAAYVx8CkTf6FXph0mKKQO0OHgIXJweTE7inK2M/DLwb59DO6zdwMM
1ua2BS2tVvLm92xQvhMNy1gh9mZ+omHFds47TFEe6v1gyzSgsugnVttmNobufI6h
E8d4+djrDkis9ehlujeCkHDpOrsapzPAPhNBzg8XxZA0Pn1h7hWYBI9pfmIuv2/w
05RsP/aNwZvNQGR1MQlGqGjvwSW1IZMNCa7A2pWdItQlDIoFSUF9R+Y/EJiU0KTY
6y+7OHVVLK2hUm2Y3aB9Nbt8eQ5OowZeiQYTO6xTzewvSQ+uCCVMvj/P019b6qnO
TfZKfsiZtpjSuTQRcdg7aB5Dygow0MBlYrhECQs6kO4sv8ugmJlggaUu57evkAka
JDbhNrNmmFiolb+1uRVJaQ/HnS+cLGW00SobFwbkm9KnnISKlo27oZImD2Zou/m4
Tn2bQuaPG1pbw7juDfN1jL0PcwsZKcmR8qiwgaTJwjI/WX31r1F/5/YlIPG7xEMO
+i0cX8faVIrnvUmap/NZtqF4NjxTnrQFDfkkUKiunjwc9IVOgkKBK3bTu4vyGgXj
u2yYr7nBXjNqgJHQ3Q9PyNiAzjHvXQ3MsirqPg1GvhvtLQTqjIBz+ABNmjTDw11X
4RczFn4fGCspG8CPHOlYwQLB3cljij6qdb/ReOeAAlabEt2hNVeO9u46AnZMWECT
WU7frkO8Az+tCPCgZYbr9vfSEe1x93kNd1VRXhEUhcSUaTLcDSNGXOseY0rDK3q6
9rV1MS4gf+8diG9/MOOn8t9wfma1N1qemlR4r7QQKlbyatggJo4IuzYhMvsczetI
Vqd1WlG4R37IZL6rXoWWQgMRZlaFEuoEImGT8lxx6eIxploSPzP0rmPIMozfllEt
s1EEQzxLHzpKyC8mMARvyrjHbDloIpRXXpQibpDrLugyMY81GCjve54hLBFDM9wt
CTY+ssYh+JLMDRlL9nJlz6m8sIR5MZTMBow1E01Jp1bVezAR0/mFSModXaRJmIuk
//HXqJoPgMzbdkPXk1oMj6u0Uqzu3Gvx4DYBeDN9oKhfL5xYvNL2NRV0y0OeJeUj
4XJ2itpg3UOKKQN/NZgAK+87u3Wpk9zKJTZ3k/7kjVFeItzNIqmhZ4aFC0obP9Tw
sCgGk8nTPS/hEZpoJjqjt41FAsOwth0ja2mAgSNJBnW92LkeXrDXLF7D9lfs2ZuK
bZdXOher5P10STKkPmRZsv2lAx6hDtT7HHZb9vWC9AsKFklrPAqFOInw7lZxRHg3
s+KD/fBZbi55MlZE5XyR2UDIFd/mRv8HhFuKpOivMdWGTsNe4MtgLKN+FcZUG+pt
hTqXiuV1AjLKhQ0zFvEVWlfgJOEDqgF4nq45z/Yy1VFY75ZK6jvJxBlUQoASrVFO
1nY8PDqogdGKFZKNvhZn8tZ+ux8mHjtGrhJ2Wf+YtYrb1Prfziftf34wAFo38EH9
HQnC434ClweUc/duh5OPB+dWYqCf1jHNNaMqH+PzejiIxz54SmOFWaDEB78WpS6c
5/vXf/IpHFElDcakN73TmtJZ6qYLbX/0ywFkAMEyvHcXmj0MOfQ8VU1eC9wZBWS+
Bb7rYmiUVU5JESVAwgAXk5YOKljTeSVX+SaCJ5qeKIXG498PMPXXxiPS7BFcjql3
9SDFHyJZfMesrC0uUlVG+NoGcJcvkbA7rcUIYIf1Mp1gzn3BsRIGvt/8s/4Mwc/4
ZIv7xwH+Ea8rFzPPLuaVjiEyFtqWhjYctNsGCbBMz8Dimp3jQUf1DuCaoTSgI/Gk
byTlioEm+EnXhMgT9fmW98MZDbAClL/tiub9W9D8fZEpiOU0FyPOS+SZr2uz/FAD
QnJBTvNP4DYsWy9YIWrLkUua6+j/vy7ecTGIp5DLihCugVsRZK7uYg+MHDP2M9Cb
M0+pHW6i69fMU7Ie1zhGfDlzyfbxmW77yy2gDVrVlrSV1adtNHmlL9GVebhwPMv2
mRLdYlLFoQzEvUfzJ7NGlvKeFuhEslmN3Om2rPqeIxLJGvoZsUhCQwTGYCjwwNvR
VTpHKAyYdItx7Y4aGmrxVl/9vwvDxorfbzIznza5v4M6u5tKOc8yiKEAQ9svbGWg
uaYvDnVIGK7SLdqzBLWJOEsXqgxXkUmD29JlqraxZuASRV8kbzhNj8rTZ3NKaoJx
W0mY1pY/XjsIUDFjshAthVn4IQyZdowa76KVoZ6dNTZveiEpwyd9olCKvUaEHFax
dSKQHfyoiq34wQBIrHiyFYn7BO8VuGHO1UTbbcsHv29Nmy/4nfxhH462VeRWbzfD
mJlSmgxg7AJZiyiDd0KllaM86IxXipZx44SpD7nk+ciUhqvEpGq0ORK3Q2F+ZZZ9
WNU4FS5qQLWm8hnFzS69VbeMgf9pWPPqdkNTH6FDqiSj3WbCpgCs71MKn2IFE4N7
DwloUVGiOV1ijW4gs/pxoEynCgNPdbl1xaz6n7lBil1yXlZv0ep9BEfEv+i+Ayi4
ot19HhyIdfjCN1onh+Mw7cF2VxNmkYf2amTY+8Wxa6BuKMNxu9foxGzKmI+dcoj1
WIo2hRMJpRpYd3m0KrD0gJAa2Gckq7RnDaQvjbfi5m5C3T8sGS3h7z1R0GNPs4qh
dPSAaxULmFDEGxY5B9eFaRXBGNYRvBpFyf6cjz8oYDBiWzSB4lPUW1NCeS6uB39t
Tyeeb4k9H5Mrb6ocGWMHrzeHgy6FMF4U8OWBIZqGfI1r9pejjNxt8mfEXFN7t2hY
m8wisolb0IZ6IIeL3zhsKSYCu0wdzIpMrDv2dSDYbgGoeXnKAh3tkwuQQ4vtoPVN
MqLLDbQSw102yoLTi28VlF7KsASlfWA2E9Luk3vCKDH0+3lFJKXxXQC1aKr5qsY1
2dE/gUam/eGsCIc/wZyP8yE9xv05q0d0pg266QXr1OnKQPaBoCiX8CUR+qaTA07X
ZF9dHx8Rnc4+3dxxqvSBPu/bbGUmGSVFv7OFiV4mBw+Er/5PEHNCuvFGIz3oUhPy
R4p9Ou5r8xg1DcXk/ZCZmfH6idcifsfLHltY8gtiax7dFICA192d3f3mzTjmEKSC
tVO2+Hz3qgtbDbbXswtEG6sgj/AxX2fUsMvN4ylJaxkMNP53oPaj6Dqgk5iyT9Pw
lQtLu8Me30kLE8ef7kxZg0B1VLnd0/3wMV2s1oaSdif13IMU/C0HsLhwqNlHv9Wa
2BCO2zquEkiCaM4pd5L0Whot3kXPiyep1ftjwOQhKa6eXITwHsMNg4jikHE/mflv
UqsDjW7vdU0hL9e9MbgfNw+FgB5LVqkF/vB7vgxbDsyS2GUtp3UD/+kzkDgVzSmW
p3sCaHPMbCsmUkZPO7AmXXglUME6nL06fyi5qZinS8T52AudRnRsOPAh26DUoESg
+a+aUvqjWCJX4XKE2piT8J2qV1o1CSF49PnfbY/Nkq1vZvVRqBG+Hvla6jBJpkax
LcSxSqo9AlFf55upNy8VDeDVGYW6mOJPVyhNgDY1cZ7Rj+8EIo38yHxQGh3wSwx+
d97AmwgwfWQMQK7D++tbJwAGIKLQ/963TvKMzhTZP5A6Lbzyt+l3k9rJrgtPvq34
q7jx6OHQ2vEqF3N9gItNG43uhhUnW/2uFABj/Qsb8ZTNROX2spnN5wxPsyx/K0sz
sB+xdxGTujV3VWLzicWMtK2omgoESO6si/bO6y9Jf94gjuw9hx8pFHLbB8RgNOmf
nbRxtf/KD717ebsEZKKnnDTS3//bLs5c04q+Yb+cqMgilks/AA9/KGxHGRN8UeOb
vMy4XYErLywWBP2FHPi/UtTlyMTx48TgD36FDpwvzNVXtXy9R9CRHIBn8rStY017
gLPKejK5ulOQT33wxYXNwfpv5GL2kUmkRrJqKctXO8s2+txv9eQMXpqpxYUhTq64
GatgQXHZiu0ynSQaGIwE+DN3WTZh37oQB6Y+ONIRZXRq/NPVpFGYkYdNePqzrsLA
+BHVVU/Gj6Jd6m3IaIojHmehrUkAjuomkZ+b09O9FDF9t5FrUpR/MuVm52aVKTJK
mLjC4dVnGMjYmQlR7ClCjQaxLX0VUBB+hsjLXigji4Cm5g42VGgJHYFc38pdHhLV
D6wXy9CKKfwS+cE857r0IyRauACW8lFX3inygGGLru6QU442wrR9BWBXdUalKBQi
A1lMkDYG7ZpOalc62xOG0t1midMsIX8l9hj1PYqBbbAm05jthjooLFaYpgIX9DT5
hSljM/7Ui4WeY+sqSIw5R+E5uLKjUQiV+GDP1YSiPQfXYjytY4kxOGlzYEIKj7U5
Yq91nHC4nTJic+t7YxFoo3JGrDJV2ChGhsnBVLh/v7svDLEK6yJ879DkSgKJjFnO
Q4wfuEZxNDVdCzIOo3qURwwbjJS8hzK/wvZrzQa+5xaicTSWn4CbhWp5a0HFKMyQ
q6gyzItC5p6XuLn61s9IIM9ubjjHRvKmv8SRBZV6V8nRa72nad10mZa/t9/Jo460
Nmz8fJMaPooNJaw1Dht9w3dKCIw82e2VhadcDzzmKP9CX6PgldOQ+wubhTY8/yaD
ACcvhjQChuI62IiES6LZRhqUPxlADgGzvs+Sdl7dCJrcQntnAHcajnuVS7Rm4uMK
sv5w+chLBNaEjx3JrWSliXx4gtagq9mEhrSNfUB8U7UQ85jCuy8KXh/8sWy9Yom1
rie9Y0Or0YOmThjOke69GtSPTGKbcTqty8ylYy+ilMcrxKEhrAXbwAZkOQ6b7+jw
Tc/lVd7s05ldd+E1eZemJ4ktib0exegyL7TIkfQWyLrD076JEQj27j/NLq8zJMGT
wisWoIHDfsEKvNQJZhRVlP1CPkYcqcU/POm83OTTow9oQH2t9nq28jWHLcZFkgHQ
3SMcu+rxciGuT4cswcvZt8pECyJuIdsPzfdkwX1r2pr5OLZhceT20L/SKnJ2tyq8
UBMrZj8/oePkZtI2rLYMDm+Unx4hrYL9c1oZALGxCmvdgveDiTaQ4P6vpnfAD/BX
KRG3crwTI9rLcCAfro8YHaqV58JAqP7gacN05U5zafeg4bZkLe1W2wzo88xHOazJ
h5eN7Wpm20Asnn0FazvUR85fT2RBTCTX7Iy00cV9lFJAewAlCU6AHNTUbIMop8jl
4tes7mlgEV8pdcAZecBX3zk2XYMJlkIZrGL9o4ilmUGJUhnioHka17kWThyJdGoj
9qSb8oneaW1iXGThhEmgCL9ttBMtYMqYz97Pp3i9v1TlzOSRk4p8zWEgNM7+UYYF
oUGl21co3W2YrbNQb2hDas8zLqvpbuuTerJ90VyW9rPPn+cxqma8MSbuAicSMDGi
/0alaJPZt/rinGdgAWfvbYnvsYtzQF1N976fwDy2w6Zx8wjo+EhSIiGB54/XEnd4
+vhh9B1T14mBAcmEE8137+EK07Sqzr6o06l/HzVcGJLhdi7xGEkGwbCeU6oAiziH
A6lA+HCGN9LdZHGIdhnXqa3xkP1AmAqgh7kBZA8MUbB+AoCcD5zennCoorWjApwT
H/5VF+h34aZiFqCKNo9s/1vE5v0kAcoBqLws1HV4WuZCKUKDArGblQV7l0sQ5OSh
0oeS1XwedGhzifQnO3aAZ0qSrZ6jWnM9niTcINKPHG3ARqLQUI4iLItfZO34Bi5Z
dXQGOiIyNUEL/J9DuoTVahDljxxqsbbEoMU8Mp8f1TW8KmqoVIxbXWBNgHaT7LWO
Yr6eto3P0/Auf/mf9CRHSYkgbndGXdoEJQ9wvwy4pKrOZGAly7iKkRZbmWC0V9tG
BUYDZvePiUnegpbQZF8G/ehmxwX+pPqZu/e3nE8FQ2D4aQ+hyI6yYRVBkogFxn/c
wVLnTuvg3UdhcwXvWMa8ihIHcBcjAuEBXuk+BdR23jbl7AVcnWnpZhZYot72pXXX
7YjQtDC9oIyyQQV/+/i0LrmprZDDzoiSpIM0GkVB/EbiBnSYEz2KK3Efgho+5ClN
VPj49DpiPI9eALUY5K6SN13DIE316WwCvA50+UVdOqBb5/tl7ZldtqViKjfL3ugq
Mune18R/k80J3dy5AfHbaX22O+iVBfAum3vhmUwyO1RUjpQeGCYcK6jlz56uyasW
OdIuqnylvCqOx4tnZcaBh+bDqBotEmfv728SE/B0I3t08QTeJLyDQPGcYaxH3KJE
YFFj7YSGpNZjcGvEDTl657+cZr6uxH0vfEQuPuo0OAA1aLPomIbYWb4/Xl8b/4vS
LlmAudHtDpXvzootLyLYM9UVqGqw93An5mitEyQ4OHbqvN+8GIn81clh48JB1i4x
maCLvg4A4tFUsWUEByMpdlce3MSN7g/cqzcEs7MgEjxpc92vvI+79Aj2wpjU75V+
qoCHYUUx8T9ZkIKdn4lWiVOEjJQLbhmzlG4H6fQcmbSE79c+tZlzNc5s84xMcnjW
hYaMvrxkeubIjF1g8zK/lHBl6+ylOADUJBkooWWRKn9pBivauh741R7mdzq/Wl0p
ObFRFC2xVTGi1iGkPTADi4HDdsVF5eCOzqrnEamdPgd9pD/P2lbzlchSD+iXU6+b
yJ8u0ICsuFwusjwrexOUVL8O8jOHN1jcZSAYqMmeQ4tHVrUl0hcwsAnCAC9IBFTh
+asYATnps58QLueucwbZbqp7iakf2ECR26di1tRkDeJcWkREaYaMOOFilGIO17pB
hhi/YpTzEYGVLS4xiWtyPiMxdCHiUOf7a7Wg17GUrLVAy7+7rPZVkEVPiYseqOAg
0AB/c6bn0k3Trej/r1v7tUoAVVpKHHHgRnCk1LepGdiMZsAyIfOsQ/xH3ttHkdmI
giLGo/OgY8lt6mSEn90q1oCJ3VzOHQwgNKM3r30KqEoKScBvPCXr3QcCFTxXMKRS
GfzyNxEv8emMlpT2Mt/kmrVQykNYbsI51W36pzZ8GQL1uXULendfEpZ998EcLOgP
Y5tXB0OAAnhU+1uIpILll1xVedyY+zbfQo156cKroQxyAg7RmNuEcIBhRXNkDEte
N3I0CvspRna04dJr1T46TIE3CU4PAXc5J5smR63MdRWTbbDaR/R+Rulgp2JZK2q5
hH35tIkxln6x42X7g1j67K9UsILfYCZ9yv57j9AZ/UytT6C1ThpI/OeBHupXLdfS
P3gKUOOyUNWaViwhqDHXI1ErZoBW1TXrKcOlUZ/8cujfv6chC+zP2ToeDAQXIsH/
KjLqvSP+6cDVbmUhGtYkmNp+Jr+eXZvZZ1ed8qi1Xg/Amt2NImI1iU97nHngYZUp
TVBZclqNivSrThjD0d7W1JCxFLTQ1d7zJNdvwr2P5h9wElcjh7Ax1/XciGmSRXDA
MGDZqZCfQxcQXhuPq3TuNITFw6Dsa611O31gCj33MBEPQiY8s1I/y6t+lidJDCCP
WqenLoRA9MQ/+tqnA4Lz/XDVFCnBbO+JhzWs94ztn1CZq7b1UtZPqOyGXt5sFglW
C89f4GLZ6U43axNyNFEWCFVkF8jeDBMvBP+K0VhiD5GWshd8UGev9Ju5Jw25qcrZ
p6y2qu//lPAd4Ed+Q5OvCRkDBTWEGLS+q7+mKg00t6i0TiYh1ObeerIaSqU/rRSm
DRpqUbLhZqkF+PhPewR4hoUaKd3ht3Bz3lTDctmJl7JYZkEUOt8cKl19KPzHHwhC
V5mO8CcGm5NP0J9xpRczwJCF1u6/a+6DYVd+ApLFFi4sQxdHeNgxxFe6Wkp9NL5M
zwsHdo4BG6LcoV2soE67h4cm9TxnJAWs8ZHZV+A7/+41JxKJbdxGL596c1/oUEER
Sbxe9wOtFJUPorrsfDJMN7He+4bZGPeOD1kD6fnmMcfxCCsnqrmemzOoBecA0jsc
WGAVJ3zg1virZchTWIWMR7VHFXK48fFbLpNNkRcwcH7234WQ1RJuJDwFnjO/QebI
dQk4/Tt+Ols8xzVE45fezZp6u6VPTVpJmN5Dib7m94BipE9hCGCfmx7WhSAbQP9s
4b0dOtqzaj/BxcTbMLPhoKkf0uqbifL2mI5LlRbHJIvGTrTzv2qX0IySCcwIdfP5
Zu1dCnBg+KbdryrBj+43rLcNrZ89DZ5e/hErApY7VJpYzS6v3fEEmXVSzS89oPtU
dMJs6CqsNYotweC9rKn+O1QGq0A1ReThMjbWzx2g7Hnujpv0GOVFo9D9RjgtYL0h
9BYGaELNslyoXojm6ONJB6RBpq3LsNFNJsS/lpM5GlB8KpQXQPL/eh9lXDjb2aLy
8fFb22YcDbAPttbuM+IC9ag5ep/zH+If82ZRscP+5unX+w9cD+BE/N+BQSRJnzWM
8m922k7rXIUImafreE28IUUTaVF1SDLxfWafbqVzPOnFfum7nylIXcVGYyIkNBRn
tJYVJhoR/Yt3XGODUfwYDvwVwe7nZhyswYltfMYHZE0Fp7hHdxs/N12xZkN8lrgg
+inDh4ZnIXJrnZ5vJidEg3HPUobLqPAHDngJ6RBfh8zAIKtVZ618kNLH1RrpByOt
9DSbnK9UJziRStD8XY5pkDe9I5By0xTqdBe2o0inFGb7TMumIIi9WKtmqnHBeQNU
3r1yf+1DoCt+dMDjfvfLz4XFVW1WmOEWaWSuwAar1pZ62nhO/bmrz0085UlxQkSt
gV44D0lAmvXiSmKua//UIn/C4N0qMP9LPC9+dNnJEDqgooq1ekRWjHBM5gnZhZ6R
6hYXG7UQaaMV0/7NSf5AaWpVW12DQ8Ki2BryhpA1tHXGletXeLiMEalRoyb+1cfq
E65MuMSuo9JusY/tgGsZMW/qrbKsmIBayjBtZa0H2LMKamIEEbHuHE5hiY+F/oOh
2Fcq9uDpFy5DnOj6Pvyu4WpcP+gXEOikzz9H5wvLU6yr0gUZ6a7tXe2Fe+MLaQi6
OBGNmVb7UhUtE3K/iG3SMSDZxFjZvS5J2fOFUDllmKpmk9VG0xxykcTTGLVXKNAn
J3v2SZqDEvDaeMTRhClysh9IoNaaaMiYLiUugJE8ETGzPqDnKIy46LhRWmkRpvlg
v65mysOMGKyxpQ/cZuko5wRu5O6a6jX8mI7pKjB9mBf88IziraZO1r+n2qbnHQj2
2qGrtmansZc1YT+0cI2dgik7M6OVyDY6zLmvmj0x9vYzaPcp/FLj+RCo2wIo+0CB
s7YssHdeUL6JrvhHW4v2USkzTy5f5e7s6wNnpkcclaQfMvNirnOtNbUoFG9szalz
5wafza+fgoJp+7el5hu9gNbB8P4zrpujaNXUKh/uChahbVViDHfSYNkoa3DRIxks
54iK0woyAMsdnMtV+nvby/3jHiDl2Rv+ZMt5TAxNWarjAqG8LFNp9hHEalrw+syR
lhcjpGs1lsITnH583R7Qz3ey16sgzc6CUFul4W8jlqFVvgnUobi8vpui8FvSwt+M
AJr8BSqXND/rzBqZJQkdRyAGytlQd5HvxDvxNDJJoZDfTdkMiBE0aqcrzW88fMMD
tz1IY0g4kdp16kRA3RG7qJxjoEQx+pWSIXG7ZnggwzMDce/zHFY+tMFQUevdBI5g
u4X0u7ywf9BJezaBu+EmQt7z+PG3bAoXvzaMZZmCHnd37wHXaVVaEvZJGxsYml/s
gT8DepVrLR/70HKqQNQuDyvlBD3IYFQdD9u1KwShPYYH7FFR+7e0wvoCiD/0tvyY
uR2djxKxHNvnPVndNDbKtHJctQJ0qvOCqr/UMsm1c42lBdi3G4qdXEPZmCkM5rfD
tfBmRJNfKE0E7P9Im6mRe02vDJOHO6tHwhu1JBajDZcgltDTgNZkqsRPY88VCj7J
AEHz7xpMPzhZ/ZltqiVr5eIHjXeJUbOwI7PaGIpVnh777zgrtcNzbpD5kKORW0Sm
Uc2FLBNV46V24kt94GSs+Is30dfEsiuou3nFurm7AOyMQcw4+QZ3toAMRYulFola
VhT4Oq1b5xPickcS7sKDPwlGl2PvIxTiV3jr5OSYjemAeFbkDMWUzs25VL8EMrh3
wcvdQrwLDWQLxKssBVG5Xgb+VT1NnKWisaaTh8JSKJmJ97Ai0ircTde6L4jyUckJ
zo/3/NLPR/H/jh52IzupMZH9jGG9J6OxbIa6rhE5B01cT+e6PTOvZbyf9CvWJ9WI
Ms07oW6frE7ksK40MxLMFzzOYu1otlh3v9G3G76uPCLj5L2ljs3MjCb9FW120tUU
JODdtgnijk/TIYtA77Wb8+4Da8itret5d1gBTfF91Sch470NxemKiZsE3CRMSQAr
pA1ob/DoiIVT72kRkkdNjrIs874/CbtOyNn2ZyVkp0LcLxvzvuVXJJsT9OaabBGf
YU5FUSaVII/wxtjosyIDNgPS/otl6w1zLDtLRbp52r/vIboINSjQ8q8+dpwbLKwS
T1suAsjEnXsjb8bfzqFHeKEEWpXgxv2HP79FJ3CmUQTKHrylxertUET53XAekGZm
/Cn+HhuZOd6JJdgop5+9Fe+bRI++5DjrNIP7i7IOWYC3iLUBQWHiCBR4TIq0u8ej
l7EVQdbRChEyYYR3Gw9LLDfRDRHMY9U1Gl1/1Ln6/Qy0mhRLZXqIaP/rMJDVF5yK
lGcb81HfrKdkBW7NYJFtyGwNM2G8thGbqkZi2v6d/3obLd+v7HQWVTc8E3qHEWgP
Pu8+lk5aX2FrCtndZg537+k1JWkdHb1NXRzA1niAmGgeqnyt866ScBmY4Iuo+Ywt
95u3MyU6F9ZRqT2km9BJ9a8KsAYTrSVDxW+FCr+PxB1FyzxFMfl0NxbXLAiHBIv3
jSTRbgpQB6jS6K7VJ3AjugnssPCXTds06iiAVTU4zS+Nq3DB8X3EHZ2v8UVkoD1t
g5LsHvZpO4i717r3QCxNI7An56f9cFa+0JFBhy4llNpGk9NahTvUcFEJ1CeJiqIX
AWf84WIXQjU8PG+oGcqNiV0e3ef1JhUtuQ+D0S7wPUKdY5SrL5FyklOnheBGN93F
VJutCpMVWL/YglpWk/3htWj/x63nZ4SNqOk97nKrCOboKVZZCXDuhI13jFIZm57y
vuO+Xr39MXfHxpLxcWsf0DCneeWpsjqJY/MVBMwS6ZA9qpMqUdSebIVP/kuuJIyV
WKlX1dRsy+iGR0f2XntIrD1xeiIxW/z+4VwXtBGnnKfq0ck8QzT5uwTLyCLZWuQY
3E3F4CAuqLODC8sxlpwTC9//4f9+OJjm5j3ywjrE7ya0Kq05jerU883ra/blSk0d
VU1tM6gHqiVdsBdK81Y4/d3pfxBTzVJUW65qYtNvHX5AAfkZ/oZg5ltgfrAJxhcZ
8ypP5bioLUPr8Oyhucu1L3V7k4hBFjlcYaPydFYvOWkU2qmRyc2RPMvOf9WEBn4C
BT/HlCGIA9N8/dIwqckZCDUCnHIYOR/JqPsNJhgpVAXMqEU34s9u/tY353qzXTbc
6vpML2zrMKk+8Auy9HmLA+66j+AakoSimHMWcKG47egFgmc3Horal9u4d90QZCBF
MnsTKB8TfEDtyH4iUI1R9gwiblrxMADh5exn6G/XRkiBaQ0IU2IunjFFA5vmvD39
5hWwz57Oh9SPR+n5YQYi1VR/KDZT2rR305Z9KFRkDDtM1aJyBGd9dcJfhz2O1Yx3
BJA25iHieeh5XuqzH0WiQjBfRfA2uR/Kb2AvE/poYpb2dX7rMuXJz94Mry7xnVFs
xayTynwjgPRBsqHW6oHXA8ed8VkRnN4FSJPWcKtLaMAf34CcSiDV1OT3aMY7/KKZ
7YaBgzEJf3sQGMZp987RB+FwBSqgOUljKw2brfSl/8WJzr2ws6zqN8Ss+8H1zjF0
oEsWK92DcP9uBKWLxjdgCncxz2ISriLsH7SCJ788LZiobeNGJXMbHlzwZyCs/DZN
PQldePuUj0hVtAOCkoVavuDHf2UERs0eiSV3XTX2zdfxFXV6hHU0micssTxJQWo5
qi544hHVt5/oQVZkiLEHVFj+8IIeCTGAr7UskdVnsQjMWCRVFvVGKO5y1xyZKxiq
X3dR1WelnnDE/gdkCQ4XyHcpVxNQtgIyRuqYJltkeDyVpssWrjMlIz9VAVym8bem
ZWXuDsEpMc4XWKoonzbWVRvsHaNH1HpNlgSDq1qIr3oGDcp2SrTPI9Az6DqlaDPX
LGbu2YJal6TCIJDus7JdtjVUzzBCJ/q/G5Z/ABEIzWFeEOAoMju0F1iA5FXMCSO4
nZo2vq+mKJ42lKYD3Oi8Qtpj4sg0v3GlfTK1s2tSRKuhajLljdFMmFQ6tbbeLv/Q
55anI1KXrnbY4ga8NRc2EJRpmEtwFpYqxEsWRKvNQaNv+UUyGBjDTQxvRezNfeZq
34KD/Ys2H9DmLoG5tjmurYLbtIsVtUoaaUW2VfDsnJ52RJ5n1cTx1IWcU9nsMJ5O
X42RHbkxXtikez6kz+d3OWoABiJo+/ybxYepo0kL7eTtT7xQrykt6TfwARIxLLpu
A5tHCEHTySJKcxqr7l7Ki8lIsH8mWMwPrNLe/CPcNZtfl0JgJ2QSwMh+ar6givFZ
EA9OfCnXu3se094ZcD8fYsanba/3l9I+GB1Zra8sAUxqZh39ImGyBBsFOp0oM/bA
dLjSVIYp9Jfx2xiabZ40Q962XdtbOYkLheKdXiGG0eLcRacMXxXYkYXSoBO+NsJw
LZvqoGAAV4Vo7Znyl/4cZM8LPdwZ6TmFV2gXha+ZF5mNZsGhGL03Evs1I1j0sXqG
M9PTeOGTx8XrL5fo/Rj1SyJwHAAD0+QWpcfIwBw7r5IKKF5x0CQSAk3b3I5qdi/6
wvg5VqSaFRH6vc2gS6dkqOdcxyRXb8SClhH08E7+lJH9QbC1FWc3Q4Iksag7jK8w
kBht2hqhhsxCKieEHhOTnQSJk3zOBWrvrLYEw1NgCgJqTqcsVebrVhHi4teMwm6D
jSd6W4mmTlrknxSJd2EdA1FU3V7OHAHFzwk5si495j6vURQ2HDBeL1v+o/TPHyO7
8JMZL3pi0Pahff8H1MXJNIw50SjRCLimXwRCTa90v6p9aGtb7RazLoHGFhWc17dE
UF6w5BPH1rqgyMGlwubqPGv6ChtlgLTDw6ZUiJH00xUg71GsT+PTtpMFrU8fwwkO
s3Y0W/UC847QLuoICyBazIWUlvJZO2iBHORBYOC1NZxhUU9jCsSYlyQRpzSzZ/vl
XJKnbANrFDIfAQLcGHaDUWc28Uw3HVpT2fH28ahdgrWunlYT2/m8Iu2mwtj7ZY08
gYY7/EBR+jClaB4RoV4z4sOWSimClbkmSlVZG+tVfxINM7BCLjQp6jZTO2S57QPr
ZXduQJnhd29guwd/hjn/1kiuA1msWVIdS00kGW0MWCsrU0UqvpdWHacijtW7R9bA
Xc+iCj6VAiT5EdXGy14uy9yI2lGaf0Li47CgsByOZe5VpExYbMt4AnFvlqRdZMFM
sqz4EDJYv6+dOFPUdzPdyBXalN6/Re4E2vewJ3xGKI1gBZg2qnRTpG+ntPqMGSJq
V9SIWw8jnotjUQI7qSFHoWzagS62NTxJRqpGXmLN+ux0Cmnqf2mP/HNtSwJMNDNl
ulW0ziKui1Eg2IcD/Mh/3k8ooc7uoZSeeM3LtdVq9GQB26hwd8vdPk1omCoEq3BK
nC/Lp6ks4FCkRMJoNovkvLJ9+tNDITGolvUIiddpuGJcjQ/g5aP4g1Ebt/egtFCC
vwIm6MaDTHnwOnWo8ruM0xljj2npjJFlQXQL8781+od6a5klcTJFW5LQbJ/Pec8g
zd8qSp0xkXJWxFAnTGq9pt02beue5Tcz4NUp+2m2/q3eyWDXN9oSaCikIvs7p8m/
2txPg5JYSHxk+Axyz+u4U74bdkKtn9kC3Iy7hXKJanGoucgeT840Em6zF5asQBYt
SAB5bcusman7nExJr/tTfI+clZKaqYBrQEIMAxG9iGfsjR89g+gcrDeg38LSsWMG
3mJj09FCxSG+nJNRRr+8YwzYTaKvoSZodKZHIN861bb4GCA1Lx1bBTGJ2d5+0nAe
M+ww3YXckK1vgF5z4NKtRK7D9tZZQrqH8T9HFeuO5bAYqOKExt5i5afdxQM1sfXQ
6+fsOfzTwo12yiOezvUTVW3oOY73TyPRNQP4x6NHwEi/BBDPQYtxhjIChyyo7Sp4
w/TFLI7Q2xhG80PQfAIeBU+UDbziM7kGF+x0sfIOBfoj5opPkRuKzKYxJWEMfncG
JSucWEJY7gDHpV9Fxi1512ovE1EaTdxDCRcF3YNxlGLKFKq4Q5DtiHJvVNPMp9Ma
B9cUfCuae4aF+pzu+KKS7Oeb+Gdnvzkm4T2GFnEOKWwcr47IKsVLuB1zyPnDvPzo
me4nfhi+FhhFwjBqwb1xxiMJysy3TCTM24URgnNOIMUFsh8KlY7fR3RFbnL6vlpi
JY3jvYe9A4tj/y6PX4BxV4Iq2DmJ4XXd1fBYK93S/OwK0023FQ2rCquzonCSYdFO
/jw+iWznyb9WQz/sVgwKUXqniEGxarTXPp6ussxNWRmivfH6UFcvfzWn3rtiF+kt
7xzivfjAlwwbppkII2sPdE11GS5x3VTmPSu/DESzZi2KFAqTnmrAsRkWJym1Gz80
f6Mg/cRJsRHqjhPWB9BRxy/YB5mpDV6jJUZbdSLy1gf/p6Qi81qqwI97i5rEdoSj
r/EPImwsNLodC78zXtNN2XC0iwObEXn0R1GIY8SrHpPKUIi4j06mb1k6gp0mwVfP
1v+UMg22sQguVOHgrycnmOG9QKPhJBLWQ8Cw2w+6kyhR/8piq6rflcx+c7kI4Foq
OLkIeIxFmwNR2uZzN6jkKSyyexgRnP/S98ZO8JcCZ6N94Qy0fb7PAxwaMIqiwkiS
oqqZzT0Jru76i5WbGIOZCuME0Zc8hY6XOi8STwPf62WIsNHxCtzglkPaTevQCL8S
Bbhc0q42Pe51pGrkiWJZXvhtfJPrSvx/uAyYLyCk6/nLuaM+CLXv5gd8AFOjv4c0
nHwGH91Z5wIWhXp4HMeInqnEEfBFvOC2g3L7WffmTfr2JVPviLDXJBiZtRZz8y4y
a/s19uIuuviS6s92hEGq4vpE4IwUkMQt93Ne/yEntVRxoU/Ye40fOrtFwZY/Oo58
FhV2ceEvZ+TyslMS8vOpEVA97U5zjhOOkF6GCrXHH45ez+mvcVBFnyKe0DR0qVO4
8uzFfQWAyy5pTX4RJRpjhS2f+mFyO+znmO5sLtQhyV6NffC6hZGfLa8IZC0TDUig
KW3TZb4bB88lAXzJMejn5+Pxg9PiLVhgqaEuCoOgrcH2civt9+nBGO+bmV4Lqe6e
xSWswXSTyiVNJ6N3W7LNq8mwrzq6VNdcQilDxOfTPhmmm0+WKbQYubkocywTzqpy
OmkiVr5O7fL7M8wsSkw57NSBoXj4CAInbJFhYCOnindOTa3oSGXiZB56/ywdjxwF
naAX7Xk2tmhLv61+zmYJUS7Ad5yVPL33rIEhDGkOcpw/bnRwbhdIpA1m3XD2u+3T
0HqnaRoDJvSJU1uRsnurpWbyXZM8w9FD++yVH6X+tVNxo4Wf2CxY0d6ZsKdilzMZ
sGBhzvlOR5rx0Vok9zeub3GAfo83FqOwnRHJnPGEzxtalsZ5XQG9VXNDkLhp34L0
d/JznzlN14ny4Er4DMU2xs9DUT/7ejt8YQT7HMJXVk1rbMn3Rs8DAkn82ZPUnpoT
HQopt/3fqHOetXWbgBDrNlVzXphVMsS7mrlXDeI6wDj5UTvF8C6a3pqNfNlIqCCf
eoLjQyDrhLAcXqc6ISHwaMszWHuYegRqwdSBpXGSv/Np/BRmUgx0ZtzOsTL7sW4i
pOm6A7iy6vrXFVE1zroE/7yZMjh+5QxmaNObvTK9NidRBTWfcA2O9QzvouKFiXnU
I+wzMdGPwX3Er3uGszobPxv36Qx0Cf44rxPn7086Zf1SIwFNlKWzyV5hY108dmZz
LDBqkAl1pHGjp/US3e8PzY8E0mDTq3S2eIEVvhEEtfd8XTiu2hipxi5UQtA//4ug
xXffyb30H0JNIju4JfFDgEDKzcydLcVazKLIU1STruQPcBlKHeVtZwvMtTbgCGJp
pzrLB3FkD/P+5/osuzgfe2C60gGuCaTuIM6OZ16ZJytyT/u3WrNCw2Y4ZMiA1OCC
Gmc3WFEGDQ2xwoY/6WxMb/OZzGeXZoCj57Ax/tAh9eAAr7EXZGMNx55xrOMygD6n
c9d69lQoeNsnJwP8/t19dW6XFrJrS/K/K0kB5P4vNdwUrPQQZRjGVnbbS4rLlcUk
B6OignMcswOb+BnKarcX6OUGU40KloHUEnqi0rLpzDFsJHlYxP+rIZlb/wQAVXv4
HUI8C5NWV1V6/h9mmmenCWDEKpYlQfXHZj8an9yaPGlctwROi4bA8NPRVojncQXn
W0Co0iv+h/zmoxTNiypGWwGE2mnWLtlSep1H58FphmyDovKnjp12UOVQfwaoAH72
nikp5pRvuD7RYwKBLufAEm7pB2SBY6NjnFv/D9j++uANLgkLsDxzT3491eXMoieY
424Jka66i62wBhObPUOUXArCX29MID0PAp4iIg5bya0FfwMCUyRe9xnYhawP/mlo
7d9jKCjtMe9/a/89clLSGkCiS0ifqTPtOvfyY84ncgO0KjtUNLcjjCiAIfyJTGib
gnXbTiUXCBhRyRrnDgzPW23zcUegj0a1WhtenCb2x4b0njHGzTSRYUSiVyNAefVA
9htpuXcvdpFmHRAxugqCxXrrOFb6hvvjVw24yRdbqReFKlEi3Xmd4zjog5MUDNtF
xlIamR21e5IhvpugZaW3B6VyFQWToMa82Fufbj3/GF+T8IkXZvD90pKnRSNIOZ1e
3mX0E1cVwtl9jCwpks7V1v1TXi8wCgcThZRo6MGmmDEHbInR/8XQw1KmczLqducc
M2F6Bot2qt61f4CfA+/+xoNnUsfBFa0fLxmP2tfb1bgn1mbniSONC8lFqdFBueqt
1e2SJ4BPVEDmcxnD5ylihgwp6JCCeCv2ssPE9o9ilC0D0F7KVaeytloFafLDkoMW
I2If8DalAIiCCBYq6pkIYxddFON8q8ZoNo4+v1oO21DyEghBOuP8/bdzIZIBboE+
bEFQ4I/jLPTXx1Clx+lx22uKX6MvpiOq1UbzTY9uWjWlpuIL7Yw8GXf09gNlj7z/
4tMpk3+Z9ILdZsOJxCrNJjVyX/RCW59V2jszz3ttC95U/Ulrp0Tam5JwoElpbq+G
KAikmxmQ/C+OK1a2aqe60Kg1hPnI9X8BD0A1rP+yF+xwrvW74kOf8XKcPjyHHxFg
oD+IrAQP17S/nnG/KBXs0GfaYah966nW9dTBsPMe/qw3r5Wn9NBaaY/I1goCI5AK
DoljLbCu7424IwNcR6tYehfZcgtdJ2U5QcMipixjOKGWXSn5IsTSTUbqbUia/HoH
Ry+IJcohdhmeR5PQyC1vWFd02FjwF8iWX9xYeB1f4rkJCqAgFxOKbUV8rcYI5RSY
UwVzrJY76LQvEOXbSm0Niz6/SiDCsMWZ03xUiBasXH0zx3+9yQvIHBaTJZG/N/oP
VN+SHJhrAnOO8wa0xuer3yp/IFTAlYxXH67Q8jfZYg9BHlQomDr4B3uHLLqvCD6R
SsgRcjJDUAJxeNLibNk675t/apyGIdrR4r9pLH7tQIdUL64cvj2q/b8NOnP1mIPD
kVjYi8KRRDNd4Te9Eezohpoe4lL0XSGmLPMmZgFGFUH+RhC813kRXq5HNzbLOBfO
AbgaYpN78WdzqtfGwK6eLBVUqBPpwcDcSFKr7LhxlyqAhF1K8WnoqCMy+27sjYKx
Z41XN9TRp1XuaS++bb8SNkX9nsERd/KXWpDgHnmayjhOTCE28sK7w7pZrgUUXB2X
nH6rvELLAacK8P+mwtaHHckDn+jOy5J0zViJqciG8RkgkT3XyiLaZqS/26DqPa4L
GPJSE3v+Zunrp+fxew7Ja50TtUaJ7GhdE3ljbZxxmspZuWXpZbGMft3zhOOkV2aI
BWQpYcBKGjGQY/+ttrFWiEqLEWX0yBNL31TtxjRgI6FIGeHpeBy8lG8CiJOY214D
sveKYnu1rItAdCZ8LtOOmCVlYfts/2Xq0K69N7ZtsiF4MejbWj10X8awdVgu6Fy4
XrkHRhMVzWmdDZA3E6ELQLC/c3/hgu2KF92ujZoTb6MBFhecj3D4RbvukZbZ69Nr
CWfo4iXebo3maxBkZdvo3NXU6dlHKwn5zC20yAyDUTm/JaEifte/mJpNayTG8aBP
KcI1BRjlm7IO+9MrIeDscdo/thuDicF9vQ2+GgeMBWSneR8kI62Zo2QbC9ONpGbb
h59zopTptsZbBDb7d7V5vluOawtqZqLg51fY1PW0wXF5WV481vaSVZrUFRLllHwJ
mmJLlgHO6o4TpbWbrwBpZmc+fQ1cjmfCe4gL0TmjmTMnYaAcn1yRikXg9npSbnpo
l68XhIepCqhKtZmuVQu35+l/A0RE7R3ptKOSPbQ3VQnmZE7rwTuiKnIwfErKTV+E
Y+LX7FG+H/JY9svwqsrKFDmu9bQgc+iuML1O5lWRPkwah9lCzlSr/TXmlB00ec0H
c4datJoBlDFU53K5H7B/rTV3OhMLMy5xBh0i+tHkJP4KdPDn31ivwDPh3RJsbh6X
43+w/hC6nkw/6PuLjngIYT7vCQ2mvkv8s9xhiGhMXEW2TthUGMAE718hwvkFeyzK
8MuCmFw8VlufzO5bRKmT8nwqI6He2Gwxoud0paszALxYRTidpZlj1rU12GTK87Jm
s0w26Y2/8B+LiK/1tz2+k3gTNjpnGwEMkFR1xjMYurEf2catKEIPNzJv46+aelA0
VsNMhpYT2Bb3O7ncy5p39LMMSIMJ9Tc7GctiFqFlsEzkPaQQjMeDFwZAZuni7knY
XX/PxUMxzXsIFVY1vNCwZTlEf8m/m8DxMDiORtlO0BBzWfcnorECG+uWbbPNUALO
zRaR89NZTvQ7CnzzA8UJ/cQ24ufSBItR/ZKpEK5QFAShiWxVx0KR7xtx+LSKwAGA
QFg7RGIHHG4XCPte40ZW7mnccKmqzfjfgHswzE22s4NM0Q4q9vlDIoFvjiF1u3sp
3I+3hy0ub3oPQGOiPdpT86TzZRO6/ghaG68+/JGNmb8GXfaftc+QQtkkg8aH1rHD
GtYOWiwWLaxTUJc9ESiUFGyfpCDlTB9K2KnXr1GhG8oh34kxsyssJEWordPkZIWk
6N5fx9BDEHag/E2+/sHYrt0Pxu88qzfOwKzVSGTK+APVg5cCWqU8EW+8CHvsUT5x
tkYCPc9SceOQ1KMpGhbGcY7sQ569FZ3k5BW34PZhTC8/r/pk3hB1z22uFDf/F6zG
+GdSIw6fL9BUgLqonzYUemVnU0LcipJ3pxTwYDrbSmoaBCnye5z30HAhheVn2asD
7z+tvrVzMlaLfV8Q9d9EWLmreLdu9zXOB4QnUhhP/BlzUJgEdGZKF8glpcgNNft4
bsxoqNBn+Yut8q5njPGDQarFbEfEqe7bf/FecONh1BN+ji8mS8cAXbEH4VdjMgYz
TjtxCzfC31EDzNuyuTNs9CbP0+tv1Q5Aby/qkgcI/lts0bavmTgzLtAPhl4t5OY+
jzE5T1NMT52gPPbbu1MoEiM3X8P7bLPGNE5c6dcN+brWvHMmEkL9Lws1gKzvEEV5
N8ePxq8dx31o65cmOcd/lod9e8JXlh4xvw78q+iSInedqQ6YCn3Pn4GjXgzg/P+1
yOBvg61EoE/fn1BOLdUH8onEVLY6LGssvZF+gaqrtVbAPtt8IeCOlbaEenmAU7zd
NXKqyFooCErz517EJmHZLwmr8rbm66/6gX9edCicIJsfDkH7kaEtkwjJtDTE1aSy
JjNGV0j2RLDvlIF6DuA7xSS0OAmzLNhrcOg1dE5BR3M85bEcPbDTc2Z6+10rZOnx
P/ouCndNUveNSvSTo8k33wZMTl01eHefeB5amhVLY0qRgpaausB1FTLWYLSyqB9T
vd/5PGNNLa3tol+oSYndqiNxtINvHm3bM8FXk/Aj+hx1n29ZQeHXsX9BkSpYKG6w
8Q/JRtmJLqfyglPpp0rCZtBX/GkMI+PEMeUyQNLNpJwOJOR47J9v3YpIpYaqHLPt
8UfJ8gJFXVzffG719DdXTuRJ1xEwRiaFNRjI+U2Hu4R1kITqN4OehwtbjeHY2Rhm
ztX6qUb3yj5/KavpLM12azyu2UkyaZSQoX2hgsSNWvQ4Po8iasu7C7trkBVHEIkQ
bF2KM9DjvusgHfxzXObeUkNp7J6ZksREXDVubpxuAtj8F5Lsf1tcdNFaoglQeoDl
OSfpqFh3kXNl++8mC3SA7W6g2VQRA0Th7v0JjAMlbpcVJ8N13epd4vHnw/eELUme
d/Kfrugnwo5xv3HGYdsvHbj6F8D1u+6U4HEVEyT0fmQDHaiKjZZlwJ/QhSDOV4nj
lHovmSBiT7RLUDoy+4DTK01HQEvvj5F7mtCFWjmwxJojXZaPa9MJzRiGKPGiZYv4
7IAcjTH4bG41+lLkB/yqX4kGfM969aIEctB1zHNcDNUCdgNSfDcj6Jf04RUkzizt
ruKdD6TbXV/MEr7dTW3SjNFOhCjcKXfen5r8qsGDzxX5FICykyawLWkRc5WDmyy3
vdRPjPkY0AVvRJ6w7F0z/xkPpIpWk2bHkMjPLSeM+C52WYxzK95QpKiuzU2G9yO9
BFUQJCMkwALqrkEwp55Mr3KhL1VMKnsqWtCLL1wk4sGR1c/93yp14DWf3gLTNPFe
nTTLZXTZ9/b3GpU0Q5kMPnfUJYu4QBKQHFoEo0qCQuNBJyXlo6w2EDX1yhjgX5Cz
yASjxqtou0YeO8gzjvSEOpdL/1cJtVwbd71YpNECtGSpw1NKFL4wG8sYI1K1rKTx
r4hxxzzhqryvOUXi38EIZDSilVZkCRFBxEMDQFkdJPbFw9f8jIql1Ed7ZkNxSeh2
j1cSX/nYmrJdLQLbGGRCbomlXbTlqwDLaOCqmDyH2nE8JCd1Gww2StVZLnPsuiOO
2SFiBVNSYqUd30zR//ljRzLrr9bjb8FsPvBLWou6PGE383fbLKoqsZJ1+Byq8DTZ
0dTQXw/7YeyDQkhqamtkv95mjD+dGLUVx354cuWME3NFVMX957WVbR/rrHsuR5JL
cQ425LfCRODnRzSiLB7xncP3neSF5pIwvL5yjbIaFkm4uzCCA0k3l9jZ4sRNuT8k
8uC4Vh/Lu5UkqXME3Q44CCdQRW0jpE77e7/t7Y3NzgVaa7c7N/PJlqr22RKUVaez
RbGXWr+Aft7bxGw06bC2z7j/WWL04wr3WRAEmeNYyUurKG4v7pmEgMwYT4udj6sq
MAFXz2Wbv4KUKXSmxNZS3bgY3qOH+h+WKYcaLq4uYa4n/qV0oIcr0RPViLJx4VSI
XMyO/eMzOFhql0YsrkXXkgehSzuWo6M1xY0NmHbLFg6BGEThUfNGIeetWVj8ACW3
EQc4awM9mvOe18Ek4RMUfnU7L7znkXNYwNrMStPEYRs74jMxWIDMxIY34kFc3AXX
2HOOTMxLNviXfswFbpl8oHLX4t7BTl+AH/Mab3YsE67U9s9Hr8j3EXNuOkZkaVMJ
ahj5lWesVJmnb81eZJ/5xwOZnIsvzk0kjIqCtBUnVXLJUgi+iTPHmTjrT2sa8rGk
ChOcAmAocFfxgP8GvnIPNxQLsLCt5Qw9TiHVEp0Ddi5rTyeZSfM5benQ3D02tzLY
E6iBqC3M40xBKj78eDLyC6qphrrvIryKsbS836ed4FuPA0+R0GvvodR46ftgatUp
FBjZzNu3kuhoiXSpqy89k58vi1E7qe9prBHakyTKcfjYQG/8c4FkfUDhdtPL0Oty
ot5dWJBVhIy9mdvdQdijzYBLVW/gku1lRttkjXduxvkoqR+2FrZa97+5IvQBhvPs
2f9Bv1y20WP3xRHUt/MFJB9tzkKABZlx6oQ5itn4TBYMLGChQlAiIIMGizBof3/B
zvr9rNd5BYaSOSmWsS2OZ2ATyarcVR0RZjKY8sLVJTC/Cvi4+y58kh4k7t4drNq1
77IcmHSk+vayLkr6KdWnd+6PLeEV4+cwHpTzcOpzsxPpTgWy/70bIyHrRebCJv4a
yixT8ducSXAaDQjis77+NvY6UCeik/uOXZziv/xiBALecsaGb1uGLAgl67R2WFCa
WKmKgAk7pdX3kbpaEwi02uraeiOXhqvrXmfQ/JkUrb7gcmmw8VYWeF4wj6gPfh7K
0taL87zp6ZFoHH7Ny7jP4n2lJ1x13cGwnCiXXQl298lUdQigftbudUo1rheQegYx
0CvunUiW9erj0izLs8BuddA2fHKXz3UL8uqhptHwyl3QXjSXp5srPHSTEl+9ERkz
+pTWDbDNxjDNN93zyjPklLk3VrIOadDlfiiZjsfxeQ0rQVX8Vxg0zwUceWks9iWw
gYzyqXOA0bgZB/o4PbdCCtKbuA6JEVDIoxamAHi6VUUy80VP/xdrE+kdfDN9kyxn
9RM5attozt1xsjb9EzdGoeOkZl8STMYe1PQT5IRaxvnHXP6nkwRE2eoeC7aqQ/hW
hsNpm6EarMxOJkH1+ib6CjdQ4GCs+gj9c3jsSjtXHiKVUfcU7uYuBqjx+jJYbfp9
fjSHX4Z4d7kdYNxnodU7VxRw51U/s1tyrGfM2yXNhbiivFT77CK4NVGP7QeEOL3w
tIQ3mcfzO7vAKS0irN5QY4x9uyeRSlimMlPN7ET1st6N34nOP+HCXNufaqwdKE0T
Y3RH38sUCQavKLyCT/xKCIG1nXboaOLWsk2M2I8BdjUNjW5WPcvhfw62GSxu5Soz
5GbD3uG/6zAt4Tmd+9ZgWl5iXDkPOMJZ6ZZePF7rgcJa3YR5uNPqB6AFR7rjqMKN
IXUpI2LJX7YJKmGA7GaJHBLHyfq2oy97eHiM4tejS0jTmIecItUHf9l0gLz/eXLt
fPzfVO5PZlmSxn7usX7BNJSxZcWWFIdypFrUCd658ME7c+GQdecmouSbIjOWOHzL
cRqdW8YO1+vF8dpg7SVvgk0vIblazUdZGo7UkyVXHo0w8ldq0BtiQ3pjKgaKWX/X
IvAJFWJpYkTgo6V5KnEkH7QxgwG40kzXkjyLc1FYS4+H1Xd11WgHshK5TYG9koxF
7yKffXuw0bs2u861ZPJk4NnALEvIgfK+EY/18Hd1525nxm6t8cU7cycvxJ3bJs24
xXrLxXOKIbWwjvLfMqXXa7mxxiOcWUTSR9nsOpgaA0bYeJQW09A+ZqtdW17eDNUN
r4JNycSV5pPj55RxVbuECZ2Ebhn5vXSbLJaNoafQZfPSN4ExZ5DBhDZNnbpFFH9t
1jTLWvJUWzljfMy/J+nU08CCbYa4ugamWnScfb0XCe5OUyWtE81NIpp/hIe8NjII
hrsxlTSopvizMpk6GEgsW7EIXt+DxaRIb7vpaOjtWhBNlIMAXR+t/226HKunbvS4
OogHs4hQcGlanq1g7DHWQQCZqrwtynyJ/AY8lPmC4nU6iLxvuEHlqFdV1noiMNcR
NaGipafYS+Tq6j1U4G+0RYLr1eD4712M8DcTMbZlpbEFpHKm4arq+ILuxEJlxvfp
O/RcV5+hVgNNAl8HeQaZmiOBKHoVGcMgOlIvW0h85lbXbPe5x3jKYXNYVGJK/aMf
qr2arotmvmbbNL0oJ2umJRJK1RgEBvwuDUHuFFnarj3WgOr1VDJg0ze+oalsSccA
NNHfJf/uHAa8WPFEuAizDKhrZl35yYfdrf2QF6zBaxvfcQHlBElAURLFpAVvCSTD
iXGGcqlr03EC7UzF95PpyFcjz3iLYq4vCjYF3qSI/sUZGyXYQi9r17iZKL3MDFSp
WptCieh9paOaa4AKPVWE0lzoQr7xLIZqR76ITO3D/1aIjqS731zeOj6IolTYGu+P
W6wxE3/CtA6pSYxIdGmEdqIZ96Cn1SoDNPNmMbdg3ek0lRUegyhCMCJPIOwYlqQP
DmZcBV5FOMgV53QjFIviL0RFT/8rDsPGdIOJEidB7t4KFGaLRVDxE6H7/WMofD0d
P8T1GgJaOVN6wXfwX/QnWkr5ggJvfIhQLA62nIDP+qJ67DtZfDoHnjG5sDkJjoih
9KeMmYViXr8eScXRVMApgfaF+TzryOfHpvudhrtg43L4IUWF7jxnVabIMb4WwSGW
PkFDMm8SXGq7/8S56jpsJedENwAuI0/p82LlzAnxAzIHBBpF5lWS75fTqB49ouxI
1+Myw0lOCvACRVF3APejJ+hCRPe3LFpfxZ9hfONzr96WcQo4EbX/Xsmyp9L42V38
AvZuWiLS3LodF83WsiXMV0HwKPVR7kH++RGiVe2Wn6KB5kH4yhkwOYuYQY35IHu9
+rZqgbNOcH6hjFthn78NVJC8sXgWRJFSUD78+fUBxxGOFFdk5IRdvG0Ge4Ldrn1L
13DI50pJuPGgg/EBMU+ORpsTAZRKnDlQXpVQ7V0wkMARPUyeO1x3gr2wqc+xCyMY
NXbL2QhA8FJd8ShlKd/YSjk547yRBSlTa1xKPXcf1rzkCu6EfDl8Fmcg4OlvQJPK
/vYppuU8LT7KQ807uwT7W6GvPHuW8GUwlA1rhUKYEssLWvb6etklttTdozZCEe72
6vzqnk5B04gZOY2YfIvOu1T4Z8aEhF1r45rjosyqCw09Vcun5jhSJ+jOYFX0DaUY
+N+gw6dZOlNprCR+Q7IcNE5BZgcMiQa/2+hc9R2M1+MHlkRo1jTjtbc9Q5HQLi4l
VLgpiFT956DVbymAUW1O2n4NKlxS9cuzxPVdpqe+rISixx1hQRrWa7EO9XpG/yAy
RtJGfqDPZ47UgfKwGtRWb2e6ztwywi3GGl9nNHu9aT2lCsgL7EgDw2C/B3/TkASx
D1G55afz2yfZYzUw3a1B2XZTGF0evjWDKHCdgn41JgUX+mvUXO28I33hlW4It3gt
skopWR3g7pl6Jnip9vSgGe3hvfBAmWwur7lk2nFpIzf//kcnHfPLD1lmdN8fk+0R
Bgd8zET2aMJcKrkX7rTU2xH/tvoVK5WWWbYjm1kLib2JMxjKrjmOekPBAuHOWOwp
B7N5y6k/Hbfg261RwwCwTibNX6eX3CB/jbdIZaLOvyfiTdkstcsL+LrqvDenuQZE
gYX/Yp/2xGcbjplOid+FVCJM81FXfBjPQKSUAxjaETb4fNx6lQBGBONpI737Wt7j
VYggqtnIcEziKHcMlhhjbwlHUl88zFQYmhgaIkyEFGryXizH68a5VE+TqoG4N3QQ
PuTCFxQrntx3tY0VcrHW6NIAyIUaHf9JpfxXSpSlNpRjL3l8PH0zr0xQDzMR6CMc
rYkRGSWIizma2I8CukS1z8Wf6RZZYAyg1XEPHHm4TRyL+cJq6glpO40EEZ2FVwAt
BKW6sJsXVeqCgGRQ0OEgA5RmQgTsopO9tgxrNqGnYspbZrbr/bcxwfMDovlWVl0G
Y6vlKopafVOGKCfp/A4B3DWPpcb4BAqQqo1EXUiSIRTqvtOaMyMvHd3kQYj033sv
BY/gsmObJs2yZtuMy01GS8qDzkUru0H4syClo6dooFY7cNps7JMW1YrG9LLjl+B8
9gQhf8Shv6mNmt/IhNv78QSm3hRwagMrSyBtNPRUExcb57MygR9Bk5HjTh+2K3tj
WI8ViRVxz4iTuwJbCNDR8I1ubbbWr9IfVegCkOCAK0qEgl8SAMGGhp/u0S1RxWRb
HY+HEOqCLxkwy/zV6ber88jYCc+sWB+ykrHuBhrhBsrj+HfShcEbEHG5JoybZUf7
YGGxMKqcBl6yhW0sGLDg25SQHCPdc9PyI+Xo8kXnOPIa4ON9uPKKQQ6PD7LtVp0k
sIitR8MAvoG7uMw1/jBadsAnrRunwcnwBEwxQfo0hrgHyGJJR95K3/s7UhxPGG1O
/Xqr013V2xLDHfbvx7Xc6Z/0nEsca+ivuKhU/osWG9TAqEtfrEa559UkhmYeHF+y
EFn4QNhDrBDt5XKrqQotgNVtkJJUHc/P4SRMdO9VBsrOA0xshwERuox1IzIeRzZU
Yeq/mwkS5T+JqcT/jgH6PDjAVdpcR4ak2KpYyK4AzS2NUubtL4Lz7qHqxv78CEcG
S4sOKJnaCW+CmHEyWUx8F0h0s++EXmc2+zNRk1kj1Ho8zbqVRUtg4jAW6j6Kqv40
Jy1t5CXm90vS+qaK1VvaEbSFFPUvmS68kRceJ4PN+UMKhX4nZY+/E1M4uqFO2G+s
NSd2IGaqtgYvr3n4/PCHtSsNSIRGM16UFiB4BD4Ws2sclznhwcfZV9C7mC7TMzoF
Ez7xM6aprWgp8VLjMTxpZT1SnsNSIHQCFuVgpOkRwL1Eb+0zH7qll6jhK2x+YqZE
vpsavirXIytM8bi3s0TqVfHiXyz5YFSqR4B/0ES8q+FvNaTaJcIMujGG0fiAYndX
Qe0yjnagP85Uqkm8diTVL8NpWuzr4kgqH2QxLLsZuzjdcEBda4mAnWGD47nXrVC9
y0Jn6zxCuG9GXwEINshTlg3z9Yf7sWzxHbrxrxy0BR5e1+AT4UeuMiFDlEGnRdRX
/5N3XXIOjQS8zMy/hZiercZTdCbywc/2QAJm8GCl0eOsQA5y9Az6gsHPdtzFRjD9
fVabg8IO5Ud/t7JJphWqu2GdZE1b+ctk6tsxMQip/Nux9jr/Voi/PvfRAi9ZnM5x
ua6ZpBGjGafZKFnMN720a3TpLfBOutMgfsaHhe/4iS7vLvxcaD211QhC64aXNNha
nUhqCFn9pVkKo9E9AQPePfeXIKwHpz145Mu/rwmwoxIAeSp4ZrHm1KaROIn1QGmv
C+OJFgIxWqM5iw2IqApwiMTkgTZ6Aj1O9dxZbCKMeICvVPMoZaZ+9JQKig83ZmbG
0R51Niqj1TWCQJvxKtDAqlXAuaD0aeC7DnouY+Ql+bpObsdg2Z51BSE3xmzaKORf
n+r1LqdhTVDs7G//uJn6Glz1jKofL2r2KvUDnm8mTHXY7cZ4LJ6GXHi9CYzGYnHt
a7o3RhF4/pL51eGjBO2yIUknJeTNLsINnAtt9szyoPYq+MTBqNIbE8OiKam/25Df
AwICFeAUbdf++4xPc+PUESVkze/kVLQGWnK6rNPsKIcLmnPwofn5oGY4pUC539I2
FK7vdEKSMpVgWLKG9g1G0dVGLb2hmlZJGKP/AUBkgETyus3IJDmue4nOaY4Y+APs
VGYkOi33doagoUmkQb3gDT/IK9IIKmtqL+ZLXwroUaDvx6xSjzS97Ji6YMOMCfpL
YJW+3wsWsIlOzuzAwCQ/PUbo1NHn4U+9z4/6dmWPcCJS5t3JjtVncWnTmPIyzvjR
jjzn50OBbqjcN1b+sfchxR3qNmyKO5wQDQAnHykstGZO1GPaJHa/yMikC7hjzPPN
x/Mcgdn9kTFMBYPh6WQfWd1QcD46ZRsnyZq+pkn6Gea0+jJ21lpRwCydE+VI8+VM
/LE/L1ZM0U/k1RYxlIvaVqAxwyMHZdwA5FySMJHfIIs7OskFYDZjX7Tj7HzgqR2L
N3Vd14ijRGaD7GGpw9eeduQtasGi9XhmtPtRMh24ESd3PH1NdUJ6COViMXF7v0TZ
V0BjFcBFsLc4KC8+HKGSodGC2c8eOqM7D9qiKS1tOuFpsbU3JDhZl0nJEkzNxZm+
xCkMPCPVnrhhQSgw1Sv4q1XChcjUqgjCXTnKBLD/FnA7PAwK5x/VM9SLvCEXq0y3
fmWFzaonHPi1oP7mBbk6hCrd2Um29VtTe6FqfOxzLHADXES0F4MrQOybIXswEjTA
Y2T4zXJ0LMIk5bUWLudt6/eqIhsMdY4XOtbaIAT8Ixj6JrQoDlYupHsb194UAUHN
7fvby/E22yFLJEfhrWPA8QS/4Dk4pFUintZQlGBpdx7eg/EL1mvtJCPQJmWDZeIz
28VM78avdsxGceXPeCUi3H2GYKyKWXDDyro/i3CdyKxeRCNVE2YdVFRQU9L32EEx
C2CwWzoF6xNdOLyyJ8quXZMA1/Nl+Rij60zvndL03ATsmroj0mcPcXKrMSfj18pW
RI3uRb3Rzatq86Ynp8TxDa49o47/F37vmpQyh0e8arWJY7TiySNO/hmqIuXXmPU/
xAmehLs5PQ4rMJvfSnteUOqO1rcllQmyZYWiQEnm2Ubmx0Tq748b2Qw0KA2zanEv
oCeI8X7xyXiBSCgN72gfzIHwLDMsD9a5KYjdL3w8DJuovYXyLSnUWUmN4b0LJ4lF
el9VWeWCOEVpQkxg8ZVyLj+LrYU3v1P89IyLpD95ly9goIS1cijqMXsUgVlClEr0
sGCEH4pNnYNnrLkoFwTb//qLlf0SBvSOD1jwBZIsPPJOQbm8e0prZ0i2qXHDOrpi
5yZpq90A0gsVcHhbu1fYit5ZrlFnpi26zHHiwvf4RXDErR+vtzCBtV9kZtVh7xXy
LxV86pDA3iXnF2UzF9WNWwzJy8xNVbR+h7BFjbbFVoFIJldA7Wz2RPPwgi+2q/tP
Lff591cSQZOYhGtXTtWz+A2yQu1lfFsmg8eWzw/it+H6UAakeyT5M0YYBOZeXDAe
dIh3LOqypUA43+zwisoEg9ZfZCJ2yKrumH+SL/I07ZYyEtZDjUA6d+9cFmej7mdw
vIlTSDJFogu2i932BBZQcfQOTX+oa2yx5dNM7cPI2OOqK4UZF2Rf98dnR+x8PRLL
RMhBiYgG5mfsww6HjH1nBab6eePqolovM2p0l0OgXfN+mxO6Zp13iyTkKABseQA4
bK1zA4y6XMA51k82HcGLZbVJC/DJNEqY5jw7eXrmk9wzJyCWufhHhCDBdPUrWI0t
Ek+j0n4FgQYqxIQHKjglPOZy7MMa5w0hyP46xDBPGJYzwcX9D5okL8jbl1gbRBGX
GIsMB5yBXYQ8pCJpZfnCPMYp8NkM1/aFvUp2uZHApI5aYoEIUbm/FAjm6dOn6FIl
bStuUfkNHCNPmNsleX4q7E1+jRu8FDDtwK62bUPZwOk6uK18PgWJIj4dJsWBbvPa
5JCzOoxWNJUYNHL1ZGzmWr7hVPdS6+8A2T6aREHNiE7CpSJ4EtOl2jLgfGfU0LuX
ukWUfjQm+yC3C1mmuqqwD6J36XAXN3vfqYJ8z/5w48K47sQDeLOFlbi7QMYPkGml
uoQhNhY56RGcCE3RgwyUUAvvZeg9E0NpdoGX1h913vJ60tz+Pyp2MUO2xRJlMZdn
abpiMgpHw4/Gd2DxmUkJQleM772Tzzzfgm/jrZcUR67Gek2QIpSTEl6Q4JmIN5Ly
l/fhawWEmTpxMFu145GAE0426uoVl59rF9b+qxz+1FL7jFSOFs1MaveKj/UxU+zT
KJR4UNPx6uqpOCTKeI0FVmXIQJNLxxlwq6StB8twPDY/9RYJwj9j6yKAHwcOlqjC
MNBcHeMseyM+RNWIni+dS8WIK0uiIXiUk6XWqOPNIfauaTa7jMnZRCOh5h6rDF3Y
6XpjAWDHz2Fghpa8IN2ttF5ProEtg+cfuzlA/SiyyB2GbjpJpOjT/rDipw7ZpPDg
Enm/y877sSX89detqNNjypa4t2gVb8GYqB5qj5uTryCangZdDYS6etUBkBzp2N16
rtjIacWlem2X6+c94d/ss6PBHtFiX2DH9bRYolCwuf0cedrZ0OLZ73YkNp+THFuc
MfC6AUD4qA9nCx4SWsq9iGxzDQ5ZxKKkuPiaZBCFSkj6GjJmfYuejsUYhq67/cWW
PF6Ihy7K2+Og31yI5emx5N2aR/Kps9FsrgkNXSUrHILmOoScnrDsIyblNa9NXnsc
VjI4t/OfDHB+2hFCtGXMWa3AelVZEIdTdASzemWmapRih5ol6J/U1qj6EVfduzde
76JMV+B9BwcQtJb0MZp5v1dbsHILINlV2nn6BH/QMpPLg9eKMf/06l89teEpg9gY
mY7yNAI9KA2sdcWAvYCwjU2tjYBartMrtfIAdxJwwC8C5gF6YwO/CChEyFhRz8EH
nZj4W7s2GAnWjxvVVSY2wsPN/54J/B/5oeBYDVOykHYKQ0QoQf9SQ8NzpQxn/P08
CCQj7u2C7KX2ANbvoIpKxyGuFBt7UZsttbL3sOhLq91tNPKN2jspzG5Y50kZ3dyC
ZYsdjjYphTBx94P8IHVJocYlx5u4kCiVNI9xDOGbo5L396xVFHPx/hEhDH36hkKJ
s7KOdstvDocYNTlKjOU7EOx8iz0bMhleZTOPCRGQKCXXy8Sw5LkV9/+0JgwTDQeI
5uNSAskVmBFZhmNINWZSYfdEELvOTYqi0m95dPNFllGJtuQk2l6uS6Cd0JNgG0fq
o8w1doZqTm7cTM50hJCKptOR00vn0BO8SlD0ElucBZkPMm6dWUsK9tM3jAXHGFdH
o/r0GMvEoQEpzQ2uGw8og+k5pqKRKqdJmW3m/1H+xVldbr017/jqh++1UsVX5+yY
3S1djYGA8EPjR7G2HJ5alWqX9Vr4rHSIYrZrnsW/bQkakzPe42JkmGx4kbMlAliH
nZjk2EN2EAfHDC1aQAJDjXaCZEvLZjb9JK/DIC7wnRy2pppSQn88nA4X6i+p+Xlh
q31k9jBxXCo2NO9jvE010RYDa3jJzCiSDTbgcYEtARB6YRJLrtLpM4e0TWSxjWl1
dAJh4iJ/IXrnqpHursHjXw41YneKjLrqtl4BRvPBehl1yOVOmjYt3XsMy/HRwobp
gPgYk0W2UhmACN3gfXKQMlMLgZcrMlPS4G8j79tBlTSRp6YJXUJri89Zv8u+FQwv
aU4bkSVau3bVzWQexNyX4wtl3yCCjyZ0CqlWaWZJOiJIDunSmmFZhxwKriojbIU/
mJIdhTMkuqCqyNn6JtMN1DOjalBAEpFrtAaAZiHFp0hAFnF/dB8PzUfpdsnUV6pN
4lzPS48+sNKJvz6sgVWIccyhMYN9gvcs/5qTJWQgmKAXAg3cJa3RFrkeb36N/1CB
JuMbg2yrTKaf9nN5w/lW830PbGEuJJmr+s7weaatkvt4CmiWIRCz/m8ms0X2Slf4
Qw856vd2o9EWMIcEDJPO6bK5l0/yVEKvCE7nK36jToS6wAs1PszZPb/zFKuyq9a0
tX3C4lzN2xupKza2dFYkYGdx4XZ/mna0TwBzcQgHBoufBypkfV4glcEucMawhyA8
Ep5yuseASya3Hg2Qf+AJRSYazSh/GO1LnhGsJio/bHRry4wUACrpZTJwzMyhT5BB
BncUaBpO9kH4dBZHZdnxtsM7JEKAw/jqVC/nXFWSkLxJsXoHzUyGZT7C8TqxgD9Q
Y/0Fgku1a+ICAvH2kRVSEGkqS5YV/ietZQp9zZHyDS6oZxPuo1uOHowParQ6gaAV
Wzy6xJuA4EKd3sIGt9YpGpib0M4x/fya1d5KlHIGFktWiY5KQnMyHhyQ913UmLJ0
SDVklC1gVyXIcR7RWGDH40m2/n8H+sSdc/28u/EfPLJr2tghXbQ5LB7ZN/YJLyrA
xgYTOz5eFiI1yxQBTnz09MQg/6dy6gmyO2XgkMuRDC2u9IPvQ7zHNaOMHMh4i6FQ
ld/Tj3Y+6YYKlkBRp91Dw7UrbgyLvv6G62Qw03x1cdRJ3Tfbmk79RWiHJ3buCLzW
EfqohO+L1Wk6ZNsiGE44g5GI98AnmbYhG4vig5Rg6O31BTtMJzg/exJ/DPORbrHH
XtL2AcmPXeMFVGFDA5EKQSGPdS/cg+suq3gQ5IVlujx3Pwfw7KUQdkW3J5IKnvEH
0IniRK4Q1cRlwQG4VwboKw7juCxk15217rMzhVRfsYGQiAEpmCFKt3vRSJa80YKU
tNt1OZe1Dza3jkLahyeWymoIc0iGXsnPw3S6fcCplZeyhjewJy+x720N453EeYG6
0Q6VcvJc6guvMZ3Td66WLo5tAgh3PuBkOEFKHOHZxeehlT3fcBcyrU8MAfm8IWx3
hSFCnvR8u22A2OCmQxHoufhSElBWNdUtfyKMSWl+StbAAacNWppbCAsq4HGE6sWv
4vPg+lr8nAPt1qSI7YZIsX4d8soezBY+Rs3AibnxPO8djBsHRgkb//ogL5vmnka/
rNgoOOyQV40ReVpMh29SMFu42p/NUd71ilyz3+GpJe/iGSy+b6q1g6t0e7qeitFJ
AECsob/7n3T0XF3P0NBDs2Wd8nIHWCcW/4FnuJf4bhkvJMLUumLV1PFFMCZ0OhgK
+XPz55phblUR2prFMFRYly6g6yQOHu+h9R1zTFQsUAhumejI7muGWizjlWCZoZRc
fYImeaJuQxVPQKWckLlvQfvZtfsoln1c5o1EEHy8cBrPb1TzsWupXU4KB+cffz2G
73KHRUy0P00+sl4BXqJJKgxvC9zK6aIgKzQB6R2jLSNqMpx9s1YzR8tAAWDrZ71w
VWmq4dgA2xh6PfPQ/NgNS6QEk+ogbbCZErtSlWJSLnYQbNlnrbxLoyl+pY9Slebp
IRMPinciypDorpQnzLGWoZ0uofn5GXPoCWDAu5FC38yBPL9/Dbh1XcGVWTo3E5U7
y4BS0EOQ0mbnEQK47G0zagr9q/+hw2M86Nes2jbw3Dqi/ellPXtokUjVM723cOhu
Ha4ZKRfASm8nKq7Ksz1SIukrzSgTaXe/e91oHtUKQIkzy3rX8z0nAU5VqDK7Ez4V
PNZdA0Tuu3C2GxDcDzMkv4/GW+6YZxakO5519H/HcKK9aLYg56b66To1sIdxoPqE
T4W9r/nVM+rg8RoPtSqjaDEEEp26GL8f+36CGmTLTHCt7U+xjkAxe0G4GMbqRwUa
zbUGrKilY0+CBVfrE/OIkfkzj62EnIPQhYLZT8LfPIVTZ7s+X0r3LCLurqGIitOR
8kqA3uHLxoaOhBFQ0SEup9CdZtsW3g9tMmFwoJZSG9ktQQncCwIirj/v06gJT1uG
erdJnAQ7mVZFo5xR7gtIMUtcZna7fa9d+8fIW3y5R2Jk+sKsjmaGsBoxgvceSkI+
J9uEZRuIIkKqGr7EjoSuvgfVaJ6LkkWE4X9ezDKRXD1QF5rm+zgbRMXZOyJHvQ5u
AchYo2XRk5+K43ey/F0RUPgaidIyno377np1v//h3p751DBVOWg1IAXuwtR58ZVR
skGUo7itgYFvbyUCrsqKDs1kU1+37iietzGO7E2vOU18dPB2Ja/qA/9FKfe0RUrn
e8kOaAsIPVhrtbqwjAji7dofQnXntRhmdwWlYv8DLdmEUHg45z5SCCGM+sPZ/jBE
EaGgEbvANBEPZmSJ241YSkZc+ikSQl8snPbNMacggDJv2LETbGjwdhHIY10lYRaF
ttXiZK1uIdmWtuxMmX1w/u83aguY4WM60yoQJPCkEsaMHVWEHPnPEk0bR77fFVIq
2nhiGIfPZp3AdKQ3yTZLNRYfbuYMntGHB851K9xJlNCSiBlr24vxh5oq43AL2WJN
R4Er4fmclT9YnumLakMk3G04MHw/w0WLPl6cTqJ5zbEfEdbTkGiixqQ1MkJtM58R
6UiEW7wwpkXtS8IRTWpI9Yz+YcsmQM8jHd3fJVXNj5AJbZE8RQVlddW16VciVlJ9
phiFiLH7Za2aqEx6igvnXBcnPp/lD9EP0/O+t90OLGTUg5+aQPF4yhKMdbqDXRDU
8HP6eEsgz7lw3MJPrv3bQ0YWbyiOYO0fypbFABclGaS7kingPRnqf26snnD75RY7
ayvQwLgxwy4IIDPOTVQyK1Ib4tIEg9KtLwzEA6vz3jksAzBi25sgXmVan4n5FlYR
F3bhdrGliE+UhfBLAzVyyXXQIezJKA0Sw8wFzQsFB3oVqt4PR+09BFgbGp4HWokp
WkSbeYzlGm2nqgIru5w4TQ6Og1dSQG2jVp+CSclw9GkfWY1gDrIUJoOiLOXcApCG
mUz16yPwJiTgH1RLfTrUTLTeWPrQHbcFBaWOKennoSMTpdOsLQQnCo3nwGb72q1K
HjgZlG4RbrSdT588qvDNuDxir/R2oohNEKlTrTX7SZaZMNRLuLySJ3wyCA13wXp+
Lyz/yZB7qNLhB83bP0h57rKE3o4CzW1gC59ltn3L/okPRp6szzNOKm4ze7Ta5CKm
c3EPydeLYZug3vA+8j+D2C1SPITXfAHZaaI+lzu7KSoCPi/Pgnj6f5IftpwoAppe
7RN3jLfNrWTV+jLSJgY1MVNgA7UjaFoHk/+A5xqfrCC0li5L4mJRy+/uxofgAEaA
rzYnixyLVkX57YsglJOW1RcVUF6nEmvh/TUm5a5CINXRBK5/OdsYPLeiKaznXwyJ
kHmbsLKUm+KAVRJjRFQK2Ke/tLdzAIms2QoOSyrdcfYjsFHYL/j85wC8l+koyLIs
HaMTxBAxYz8Vvjg6mSVfptmsK4BVHD6470QnjVXtHgesiFBiXSS2rBw700GAE/CV
9B3ZeMu+Fv4iKQMtMkR0BVTZlB4yGfujIXrJeV8sEqlBBqRHOIysNr19HTSto0mE
p1FKo4Kb0kvRIL2KUeNCr5CKhoI8G42pddBhVY89GZwT4GDkbMuRpMBYPv625yUx
L/Sg4P5QVJjy4L6qTYcbsbU9qRpkP39hFSGiqZxMDSV632Mo8DduP6bGO9t3+zbt
YOm/u0ia6d9exye/A4XztHydkbuVFt+6W7kvxxcJY+zR4Kz7kyqG94FUl3+i2aIK
cEHr/dxO0l5nfmUU3oVwL2E6ueHUKoTk5QTP63Hhm/7kNcHRbc7dcCDqPrMWGvCk
+XBl6LCEIgDhE5AxcCL2RKnh8pPRwRNtdR0VPw6IEoQ7kdtGs9KNMNyB8hpRbDzN
q+WiolVzd6usWiVOVGMIadh9I6QVcjwiW5b4tFfWQuEc+eP1uFIVB+FwO3CUE8M/
j83Gp3wquC4+FqCc/IucinVFUW1NpsZqXT7JQhU8iFfYt1gG7puheduthoKgEUOU
5OgamQIPtGTJy2tbHuktpsYl6OKM1fRxQoEXwHsr4ABj7aujIIY7gGhVavUg3eFS
QGZFw3iI9fMP5LiTR1fggRAG3PI1/jy2ZKkAbTP1Sp28rTSsqDlU3bfaLVg/Ixz6
itf0KZu52sO6Lmz+oZObfFm0V5S8MkI5J12FYa1Wi+/gAba9PqUJ+F0ZMOFMVpim
cmuXkruel17hJWL2s3L+ZnkGYD/cWO41dxMBOZjPGOzq039K+ik+1sQlAn6DDshw
DvoBwbIaCRWGR1aJmvrl2Ftk/GDug4QSYOJmR0qxZ63/Wtgdo0UCQG5xD3N8kGTt
LJtyA/haBfWod0Re/b1YgWBVfgxWOs1PSx3PG3OfNfJDhUSd7D7H3RgldAUqyZb9
f7o4C8+A4GURLXV0fSXmKLljMwegYAG8KtImLoVCy34VRn768vDnGOWRBMXrjYbX
GL8M8AsWk8bo+T5JK/kVDJzmMzUfg2E5PoiRcOGLImH0a+2bvtxteRvSr/6u12JX
NrDnyTi1eArnTHr2yOaQFvSrTXWqJO+HcVuuBarYknxG7hteZYI1xlXa/oZhmMrX
2FITQ1YxE/sZbZrX6zSI5Z8ECDevAqPqAYfsNOcXGfyEccFFAbgjKFaYRfnajbwE
nmApUaRDzsq3sgh8NtwlMW1kFkB8ra6XC2Z6DUpn3CJ0GMNlV4+WbKNJKkSBXE0M
1R5jV7Egwx1Lb6OJlsRFGb1z1dgKGZ7/lCNwYss9EPQEBUbmluPwzdBF/vRT9b9b
wb0nKL48mLMqHJzemxfWLf3dM9rxTxM2LUDl0l9yayo2K7C9sBRgyrgk3nwcZFDf
ZozB+RvEpc9a654J2DOfA5syGGD/JE9xqJSZxYZMTz/4cam+LwEBOmFj5FXQPspb
QjVXWKOf40nqLz9ryDiivIntTr4sYXPpvRt5tFBSaxANp2Lg1eAMQrVT/t0iUxse
SpHJBwdif8CWUJ/5XIONi93pHO8+BEaeEH0uxjzgan9WpSYoI0sKmoUPsYIWgG8O
ys9KK0icJYNWA5MSyTGeKsBNB9ZI7rdQ07V3u5Kaar1mVIjF3MGebt5n7CgYT85n
fuTRxxTOhLG9e8m2sy3Nfu+6b+IONCDLRH4Vnad5ottG1iBO7qcxKZvUePq4+5I5
7QoN76u4HiNoGEb0fNlsbcDS4AmZ1qKXaodAbicXqviZ23Oa+oRO/audoYnmmZu4
Z3q/R0yekquJGGHVSJrmWXKOO8CXy5h2JxRfwnV1B3VWYWeHxsDNE6+qVgL62h6c
hyG4Ge1CDrmXbL8bOXY7Ou0AYsuCR+fSW9SYmbn537mf9UZDqz3N0yxr31IH9CAp
D568ckWI2vEOCi4UvlP2b9SLFC5lQqYuUbZwDg/N3KhGwGLvhFYIfwn6qCinBVsk
C2N/7udbZq49RYyOoXlg35n7wuYAfn8QzI3wYxTkLKdo76z8KpRRtzzGbQnwsGgk
h/M1VUWI6j8w2JleIdDSWo+amP/MBopHmg7ZSobjnJbPmgd6NI40ao1w7ajhi70i
jDE34LVk81wc4G123PWybflBvJ+/Ism8LobeJSmoMnLLS5saoOdZVii7nI5RgHKD
px0AoKNH8sKBy/kBMOM7LhdKh3POoeJmdkValqylzuGsRTz/TCpnttdFJbtqccJ1
YGPcWwpF8sUj5/VS4kRRVmZoW2q7o1sOAQ4vkXFw6mwKAQ5o6ojjmYqRzgpPkgcj
vnSvJuiHowh0L7oa0Io3RsN6yco2IsGKkvhQlDO+9rBHOBHMNg5NB/pvrEgqB/Iz
F2KmGMYouFYU05tUzAdsHJflWL5FyZLXUXYz1uQd2Ej2pCPYNXjZ60aAu76IgzzR
ixgBPBIck4sJf5Dzu36VknuFL7n6D7oxxD4B1KUIlmDZEL/NAfZPvAd1lk6MSs1d
FYGynStqNevRdEwt1Lp5CSknzdFiqSfVTBKWAfcn+nnDm764CQBAygw9vlbkGR6n
U2YF8SSFt441Lm5eufPrKQphe3JPDhTuScCEF+s0+VcIkdS8Lu6/vbqoAEixaMkN
0C+mn2SjxeDauBO8hSpZwzKe0yc3sz+rKUj09ERY7ZFDiCIWOR5VwuVDxcJDyRb4
IOG7DEpuQyGo15Ebie6bEPdxdeHV+Q/FOklSIt/hX9166VnobjGJEN1Y6AHwqLOD
H9e+TpgeDP1VJR7QTcrGCKahBXwi+Se/6IXmuGRC5KHJQtzhhEDWSDAuMnBJlgSx
RWwyuucdWZJg32j7mK5DSWB0rNB0RQ6RDU5AKhN5qMlaC5YA9iWSeHhFf/74oKoE
NaLPTwNJL6DGj+ez+HRIj/S1VG7xtvfDBnBZUIYVTJwuHAqiDWdEBuJs03F2oM8k
mGB+UW0HS0licxbiN8pT1/66NHMUfAi7lazXLNRYyuTWDzQ5Ly48z2EHvSPMBMve
jjPgGUqOl4l6mGbpHPRVoGHPdiB9Y0+T2RFQJ7sNCoZljleDnEWepeaHedS97QXZ
FbvdZqXl+Ar/ARaRl7OuHuHZ8mcu0s8k+HHGY1nvq6A1J6lgCVGem6yioS1cBoTb
GswUcbDldgP++c2267TCjkJQkQkC90n0rz6a6HRXuWlwxaqPK4s+R8DcjKO5HW93
wEixCTNOiyOvYfOpF/k/IrrSxUnT/LCt8ErkI4Ma0aYEUWbVUbL3my9MseEqFZVT
rl9oiULbeO8eHTs0DNgTRJbP69ff5vBe2Rt/mp3RoNiPsWOyGdauhHpM8+V4//PN
ILYi+z/NipAc3DmxwYIe5f+6zFZ/nh05B3wu8djLl60tdy76bVmau0kJHV75+45q
ajsY4GW2InhM+SX3ZNDlPBYR1crW1lo/p4xU9m/kBH3XzFk9TkMtsnk7ka8T25XB
A7l3s4gg7Qx9bmWx7okrzIF/vQHs2oBkSszevuHo66zsywDsahyXWU850RQ1/k/a
hOz+t2N0U0vRO9+8BE79XdNEA4tB1lTotfOgP5Eb5MG4k3PHXKkja3CdFuj0r7xa
0loXHlim9zUgIYLVzIwFNhmmWvyi+v9jR0nP4RwZZL4dOogScOAquk2+F31bvHc5
/8geXbanG4OXFaQbmL1J8TkLynun/GPaBXoxv3zKn1s47dhdxP+zx7pxB2ppYTXB
e1v65bMCxoFwbnXhK/skTfBJvcBOpwaBTrEckXsiQFZRq6gESOHY294J8gIBP+QB
5DbedTLJLES8dpnZe9+TML1ggeQlIWpW6/sZz9hzek+Uo59wpbMwF4BjZwF/cz5y
nj58CbRkZAwJ+CTZxdLYA58Jt82hz0KIjrYtUDxV3OlH4Drt8ukuCfZ4tGf0tRcb
YUrzK4NR6w0xfpkn6lzl/cbxMSgosg4iWRLxjLBtDGM6C+4szMQ+O18TTK4I5IKn
yeO2BlNnGj+Pc+fMmhqEFpx3Sb/YXhflPS4/y8iVFJGEj3DWc5FZjUFanJZ8D0rr
UU0TlpP4m2P8nr0K6A3FOZg++9dCf0YgimydAvXrMvBzuY8j1e+mB+XcrLfZvTg7
GzP+2zBj4umIAMSJn7J4d9ZU93PGSUVtBS8/kngmNbVqgwLhXODkFG/7Sweq4Q2m
ThsyduMZSdTymuHQvm1XXtOsuFo9ozdXeYpUX8xeezWJYKl+m0opWrR4HZEwLxZ3
DENH5wwL+bW4XK4qvXQcslBIgO4D1TCVRvtUr51aI/UMZM97yFTpGiOOXWbMTLPh
ryinOD1Dcg2p7RwT0SJbfdOOTWq95KmGVq2azRc/Y8nVy4sh2jNTuYYV+L86udBh
YZ8+cmEno7cPA58CRmdGEY11Fu2vYvG6ri7WnPBd3COqk/o4n3igQZmhbMZGyl2e
oWOMkywj0J/UPo31VjpA/a5nebvff3mDQoy+xNGimFj9Vs0EoF92k9XusdQX/AB+
dampuS3BzPomXwWFeb5QzGMMp8HAi9N6lpVzv4KRl27Q3Rkz43pTGR19LOiQxmAQ
6YYIKKYEHCKrQZus5nXyvzNTPo1nH9IutivzqvlT3cN+zVrA0BXj/JuEWBxpZm1K
iWtwloIeSkNWujnHPRzmRpM43QMOAopwLKGyk/E74hsj8HZlZlcJlZLguzwLA1Eu
hR5nbblL0jgAnu/JBbG8gPGu5+In/zw+aU4oc+s4NoD2rp7JHG/JTH0/mokqgSOq
jiAh/CMX99n8tkZ1S5kJKWOIqPfsFAkS0L8em533lWTt4sQlQvHIS4zXbYDSSqbJ
8aSaGwK3+7bHtncergs4t/ZKm+MFtd4Sj4Po1vImT+ia+HhK/BcnpziFKcSNEvLf
SGZNxYullbwbfDTgwxV1KJZbt8RT5EXTvPa5HpcmOKCK3gCg4c95bXUXrUBqbdTx
Ohh9rvnaXaE5f8uumlosWR/L9UR+Gn6b3KrofvFA4yDaEqD5KnauQCAuc1BY/gqi
RUVhB+jJIUiWpLiag5WJLEmfVSQiHqZ1bUGHtEd3mLUQ7tlsBm21HlPxKlre8T9/
XKYLv5u2A0A4J1OKN+CrWGuvgZaxaSrHptkRuyjZwUM3VyEJP8CoeWclgypY1SNH
eylu7z/AVLFb2klJgZcXGj0kohX+vuI0NM/FAn/ZHcvQkIAnpIpkEb6exaA/bpQe
iykHkuV5PSR+Inn+i0robrM0rtB8bgZwCXFbcFtbVxGez4qbNdOu+Fzu8E4ckRtG
JxmxRtO3/G4l+L9R//+vVqyskREVoahyKvQj6VHxnmVwxbOmWdeEFiOkN7mX9Ipt
3Xz3ixrChQkXEjTiubHw5DYdEikXhMJUcpEbhp7bVp8wxtEI6WO0Yc74PWU16Okj
5zAaE7gdWfG6/5NazZi56iC0vrNUo2mU7KNyElFpbFoVL4cAY+i4faYHDfGEyD4V
mmlrCbOpXqLUMJn4JIr8dRS0dmVTNWr94lyJYcSPj0rntWsZx61jyrxkFfJrEO0c
MdbiMPNh4+RrjeokryGRD6GNkHoc1aeoFmQKYN1EqI/NDsRwkLVv4Dc7xEiPxSZw
vF5aEb4Mfs8mogHIfU+tGcZg2rF9yd3aqJ2qnPPuk8s/1bHrzI5+LUc2+55ihhRS
78vG4ZAhnKE6HbdxHWZLPnbjFcGIxs9UkCBRS6+nKJ9j6d+ruvkfPmy61hxhOc30
7/eqsGO1dd2y1rtgKDP4qZ5B1SPdXPxk1LIBmSu+tyoIrF4yw3R3rtc4AwTRtiTc
6AZKXB6+i4m3LRdMFqkDtPL0ZEZWzjlJaeJ1qjf8itBPU9+i2+0oCieo2KUomZ5v
QH17d45x5FcQW5ysxvHxBuhIuqQ7UbpyeenaWKoUP1Kth0WLkpK6EPsPDR3ZJYT/
AW/XPqzRbFdixJ9TIJbxbjtXVORQoA9HwZaNs2H/dD7iWhchIOJowQLzaCV4EzmG
oxdxXnxDgk80oj6S9wshl66jvDi8d7gohQIkXIsXqArynXv0twK5OrZby77Kup4K
f/BcnwqhiX16JEfj7Q03wz6t+b6FQT009ny/TQDJq94YXkQ0C6aX15gaWgNcKDU5
xQjAWal3YIn3WUKEmPwcXMPhPmKvQRXfQw16DYwahLhAXlqmlznLKWyM02XO8QS7
yXis+lZQYQAHFB9ugjo3HPXebCsWAfmnOOYDTv8xAFnO8eqRlU9LLtLSThxIgSWH
3nsHzEV/wxsvGmpCtJnlwvj9lt9hBr32idvw6PMgfRwlk1NlPhhSjR+cJpLxyJnp
MwVvWRU7ZWzqjhjCZ5Q1HuNGHF7qJqvseDhSo6G+Pf47gsWw+X585hz/+VHwALFm
8i7m8QKm0qdWOyNM8QXer5Gw50GtvIXaSh13WkH18Pa4cbpN/bhVdziuITXXIv9O
HQvQLpGK2L0HS6rixgmPeuztkIJegLce0ebuxUwScAcLmuMmdJ2zTI7vox4xFj+s
ayLq1XsMGgP9rkZGZEaa4zuFU2cIVlJ9VGJoZ6bzVF+R+JDzxnBLL1c7We1VtN0G
OExG3p4yc80OcKPuOYJhKUajYjPlo1cEoysDYxOQUb5d4j2Wf4RCLHGeAqCS7vQP
p7FmCYaJAdALxmEP34COa/gv6BLoqTQfvyLWFz6PJsQsXA+0KTVTEi/gdJ419e/j
7znr4fBqNx8SWtxtw1zaqCoSIWy1jFh0x4Xy3qcFkRYFX/yYVXmsuARnw4O3JJC+
JE59QESMcINqaBx3V/qUapcamIRXiVEIdzZnc0rrCcryPYU8kKagpCsge9u9OCWv
7677S14VU5BOZw8m9u9ZZquYrDG8zkFTD8nlsxAw1EoWOTMhmax9UwfPadG3TQIq
UO2B2jcFrhTfRfMCRtDQvfboLu+070nN3d1Cc4oT70dADHfWK5VxtRiXYJgs7jGY
b8d+vlk7SArvQraZofVpAFAq2l5wIH1pO7D+inunN1hMIq6qwMnIyX5QYDe1gHmg
6n/5zowDQeDBspnF2x0o20vneGEz1JzeHam6Cb/zE985WaM8l+HcK16cjJ/m4U1M
9PJX4LmRaHbV1v3Y+BO1qPyJIc/la7FrNrd1xDZjyEnvtW5pcrIgxvPavhRnUuSC
ywtkjHHBBGNt/rQzJexne4x9mu9O2+t1tQ0MASM1HCjWEVR7pYyimNGCRuylZf+C
dBkEG4/mV4AhsbMkZdGy8CjBWR4EYCitlfjoYHWqUlvMkbWvCN2CPfp7M04viP2f
7dVy+rNzKVCaGzYSgL6HAOBWGigQ+3/bKJnvNBHILJQXWoTtUy2nTyD9mob2DV9Y
Wrja9qx/IQNgBoU1ibW5q8aVJL68o/eglSwFhbortyXte8dmKDpWte2v+l178iLH
DIiGQDYrFenOqSxpCWH6FU5aaCVj0MZejvLYCbjmgJxNB8peH5IVa6G1AE3M8epE
v/NGjje+m97aEKVQwi/y5fJwgJW7UWiDi5Vrh1YPIe8XmL+bunJN2Z4JvPDea4U+
StZ3i4R3Bdxd4C4jmmAVa3jzcnaOftFN6RNT6vNxwmV7NXPZf3zeY9XvlfWtxOpY
zeVe4ww9x+UAEjQsKYm/Tl/IZ84Q7tQ5g+XJE8jBJiI8nuGFiC2tc7GJV1EtLEyW
XlOQ5ZHXQKJv4tUET1zru54V4AfwzfzwnSFuuFXgf6tGvY9GCNJFxT7OYEv/aCFH
8gLnJw7LOiWaXBwDxc4d0mj72F154d9kNyoZIvyY1xJCcVb6qda2PbmAhp0cSTcH
3ytmDFgPTmrZw8nt1I71elmcfdNZO25nouU59nDDtUlkWO5QPdgchYEP8tnWtwJ7
9KT4uq6rUvQUz6drGluyChoBcO5ALmp3WAJ+G/hi0xvqqSDmHpHqgBqV5s6/Z3hh
5QUClF/RxwApPi4pV7fi3J35D59XEey82e7n7h0LJa8yCvuNw7CjwHC2QGy4YPpw
l05Py9XmJNTKDDp+fwLOcSVPq+fp5/41dDRNcMQRyNBQ50Z/2fR8nMTRYNQXSXIi
U8z0DL5Cwlq6t6//HphpXNDZw8f1+rdQkjYXDa0BNTZRi9qTrtudW5xTVKJzO7ir
fwzF7DyGRDQgVmU9iTJ/xKyIpn7oCMe4Ma+o17grGjoc+MwVnNme8EfdGhTlIKrj
F9Y0CeLDReB8lTSNx9m9zJ1QSPo0voQAo8lVz49d5EwDXZb3rYCzkeMX99bQKKBO
uqNnrnoJGrxo5L5Ic7j7crJEr07nV59yggIpHUkNWKoHInrfChrSPcvHYYEpnwoj
au8mH8aesaAZIvE7xeHQMqRyvXBFY41g5iB2PLNN41oJi0W4qdPNrJnYCgo1by4q
LqhCCiNylZ9P91GI6T/1jyH/+SrJ6gylJvhQgDxxiYWDmoz4Y2LRbD8kySKC1LZA
ZOwj2/m9lmqeC2BvAk++0od1XEKisntye56T8y0Zo3Lr1R4yWjMMbunKJoHKdKpL
jKr8W024E9KKakGyCU7Vw0rtVAF2pHJgV+RS05j3K8LR0b4IDnbUSPSD0V+LWDyB
UvgOc8ibght3gIN28GJdwYekDqhSh00m6/2Kkz7C2PuWBrkD6IlXl0epGV5hn6Ej
flN8KW3Xob7EUigRz2jtSTdstqb/O2fmcEEWb3BlishwtHuYqk+uAAAVx5X8478R
TWw7bgp48UsFNznICRfUulu+DzKOBID+8z6jvhdSXsMTk478FOb/r2cgdF3JGkL/
0wecVJET7D2cXszTIYDB6tI/REFYVyba8o07dAZXoi4BhEZR7QJeM8VvpOA3+cD8
uXdfdWPow4EjkEdWLnfB1NQhQxC5ltCztB6Q6iQide9YAxUmLHTCTPmvRrh+FeUj
FK6UajFM/xRfTUUsfq6oPrXHKnBfnZJAM4Z+kdggY9oFG0Dvg+YSlZ7twyZ5j/z7
jKkJYWgXv4Ca8529+4dVGcEMyl9rJqQVIt0kO7W4hqIIRGe/H2YIrvd/Kg9DtNvl
QN32I5s+ujJEPAdpGYHOotK8yUK6HyydQOGULY2iaZJmJPFQD/+YUv5k1l35KV5H
4vglV8eYeqgnmg1VPnMFlQlplbVhtciSeUVfEM3UFyd7otcKbVH11SCk9yvvvUAn
C+jIhclHZ9mFowM6ukWmxgQA4bC1bbfDrdzwgYqbdqr4SQUDdGt2YznqBLIlzL1t
OjAJW9fR+BJHVc5pPi32tdBn9xtkutLRemP3S2eRbzMcp1LyEdbgV3vv5TnXsw3K
QK4WPapCfaXEou2TaReB2ETeFRrnADiCq7gzNaZE7FyJ0qx9v73GBPVwIwJJjOp7
2roN7DGPkE342AcrInhefzWrJZ+gOcRcKNOEUdV/LkTHgQtsRn6lFAZIZ5nhcNzD
DiIDE1kpQW90yGr536hQiTWfa5YfjdqpMZI2lVkFgd5crioar4OL+GwUJmqho8Mw
Y0/UeSzoS0jcZ8R53jw2i4c8anUrs8ulaz81fb1yOfsuyaYPROCK12IVdtzKgCFM
BVYOM7m8Hzp2eP/BCXnlqsgXFZbmySlbSqzXwCFsX8jn6hcclnR/SVO9wjmn5Q9u
0aKIe9+ulOSVYSVRdFsqx1fIfmt9cXOnHegVG360eWedIfQ+X9ANTHMn+ZcoMyDG
TvCp38KC+qQbvi+we4QAdzRHnlmT7rgOhZprPqkHfPsvWm/h8UBqVr0tM8puGYi5
gpqTJIXEWvotV9+210eoY8gFtsluIxI8OYnWWZuJKwGsFKgpwKvQjzDny0HrtiWq
CPQW0ZkkexM4C7YbdulvLrKaUH3ZIe0utMzYcq2YG3bzJNu/SU5hoHmMC6B0yokm
24vc8CeNTIFeQG4OrxMuWSTDM76/vKHUxpttkFuYnIjXImgkHKGrvQC0/yJxECUs
SfKKuyBL4Nk0FSZSd2DWvxLmNKZFMfDVHNMbvGBChjPc7VuUqmDC4XCrw+a5wttz
U2Rx9NV4OjNC+zsj0djyatdngxcONaIQggpfKfWSPAbsFLi9G8DOkpxen+7Nn/PX
by2qH4U1Ye8k79dz4uucionF0FBQyp721csKxZZr4NuxNNRrU1TlH2CpPS1ybz+I
Geoe2yvC6q3BHJaCoRk5cUr3Z6alNlSzis3qVrh0O/2s2xCiW8KaY9pNb4U54Xbm
w+q6NA6eoZmp1ecTIJ+uTlp1PYcfdZ9U4KXfTwdhIRqEiTPK+W182UOeV3riFGIg
4MeAnwE0YNamoxhsq9FJ/3tmpGs/C9r4b2qtJ31Z8cZk5AZj3u3Cq07xwa7RoThZ
UqnN2BjB/XhJRK5/KaEAgNh4IJRVV+KnnFIFkEUVugbT7xFiM6JSoVD603le+Rzq
eIc5WIpsYGloSyB5rKJwU2A2yQl1R8BhOiNn28ZzPzv8OIEd/6CskQBiVIDlRXJk
2qQwprOiheVyfl7QaSIdwKxMak/GjWjULO3Yow3wkoaPyZbdFokkUbmM5D8Tgu6c
e82pcWgCnXCxfUDLNh7NUFUbg/BaZMAv/85xTEilBnu0w7lklER3ccpKcDhB0UTl
tOTufG84FtOFJWwlj98q2eaSYpvtw7ZF62TcmBeBm9zwSKp1wLSJJr1NdYbi6YiC
NL+7HLC+9hfMED844qxtF07e1Td3tBd1yJS+fouEkCZlRQS9IT/So0fRJap/XjWb
8jtTTs4aQTFGnF1hBY9BlsfSrJCwyYNp3KXWq3sBEadpM38oNHrkmG3/hDduxyNu
46cHBWWrYq+ewA63T+NKHZ6aqzc7pto/bJdk4UE+ZpJVF86MXiAGkO2G+yKi0mJN
UXXEStOZMrVlTk5TdO5zUh0VxGqVYXgi6qFQS0jOhNSK4+mRzjOdxwJscH5nPpiH
uHJWjA14jLguSNHzZp/xHAb27RWRooDG9P6uEWmNyam+Ei96ADCWEL3izuAaZ9R3
+Zag4265K6N/mm7IgigbFiYLeuKDhvAG3lorHjZpgf6OWgEWghgOWVFXkP5e7unM
ZVaot1x2IbzERSJw8tCngpzGpLo0iJk5ke2vCYoMXH8p7EW9zSI+lbfIiIgWRV5F
IQT2hk5/MzJaUwXES1XMbf5RgTrfwSyH45htdItPu6yjKB6vMkREoj+saT5Swu3Y
YERBXyM/I9NEyu9DkWmfMiiJFqxN2SjtAeJYCAtEnjlHCx++7fsQWWpPq7ZZapqw
wQjJIolDrM77aicmnS6M0apYPp3tr9Yfthjs83O4pCxVH2LSkbD2nWIplw5zmGOd
YYnNGK6WFfE6wPcIjzxg4DnHMGzFlkcNKrAB3dnAyRK/6tY6G6aIN+iuE3nROH7Y
INYaXJ2+l1pAYfENhTrSJKKffEUH83rouHLPh1j/c67TPZsHf/CDNRDckayzzNY7
jcDRpT4lE7HrfyaV5iGiHaFnzH5A/bZOS6oNsslnQmMz1VOOpEQ8MpzpdjUl9wyO
4v3bl1yi8qXCInZwSvBG1L0Mj/Ua6hZkqVbdtPZOH5bPOe0fCy82nP1jwiVWvk9L
let5HgtJzLWuCMIQWqsXXX+yB4uSYSCA4IcBZcXwxzCXEPhZxsTpipfXijQyKtPS
y4WfavnzJPluJIxIrq2f4aUdGRBMtFGE6Dgok4N46xoOmJD309okW2vuL1B3zx7k
xPzwpghcqoA9R8z3KuobMMAavMIoEI+QkUgRuDbkZgg0NiW6ozObraNTWY0N335z
yomdrsigQfkECGvHCjPXWz1zphs/z3+axKkPCSLbz42NtGydhnGAJPU9pagSUCVb
t5Q+vt3y1rc6tl3Zix5gdzq63wW3tLRb2cJtOuRHiv6cpWO74rqXvAF7b8hLJwjE
345D8f1wzEWGQdEfb57DabRdFqEcvi6vLiDxPEcbFM6N4vx0Xqep/ofQIc/isJ4L
tPpxhdbPvvcToZbgkTWECpxpKCVCYmIyBI4ZJ7I+9IpMikMAX0enoph4zSUJUUcS
/kaqEqeeZdgtMTzvyfRqEIYplewylXkl56oSy9WJnKacbFibZ/Oy9FwlbHAueoIe
iXNbrbdghVket2QFvBIGWZ9SOyEBKp9B8PEkEFS2ZuYwmpDfZjGouHjOwo2SJsPU
DHFBYLJx6+xDEqUx+UzGJQh+lAsQY7WkDNaFSvHMDfAvdqfwiypVJYjTcnI1xo9P
InlpEnfPyESFX2hFZ3KCGyCmR7Jb1LeLgsVFHEAAfY/V71V7/J8r9Ee+I4Q+NFzm
byXiNfGcMP3+Dyc/8KuKKVdvkg2WlBNGsXwhwSHg+bURKuaqJf+ZDyZG+TfR+9TX
v7SNG16kj1bUREjc98WkStpjoay5cTxMifqe8lPUyBxukBml1O4uhStKvZB6H8pU
EcdZvkXqpeqHjnL/8pHbvXZK5A9teNhlO1rhAsg1rnWsCnzx2fj46wfQbC5/474G
dAvpplWtLM+p827wPj11h77cS4wxYQH2ymedCpDrIx86n2Fp8mi+V0RLNcEqCANK
Ke1g/rizBu17AEThp6L8u4UMiUleFghnek0FJMbRzBU5R1ctnDutX944UaPVlbA1
pmwg8+75iTJQRmp5AwYSaZUD17RQ3dCyW2kY5cU7Vx93XWUA4QdUnpyZ8lC1zgSF
`protect end_protected
