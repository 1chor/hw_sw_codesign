-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
mNmY/vmsXCJpCfPc4ceEeAkKoDKDUFmH2vn4wKIqODb9BDC+MNdWZ577pGFBxVKC
tLEBLFYrj2dDtJR+NHIw8wnP1jrsUWiCtnbzdm/CyLfCX/gIwbrCo/Lg7EBABo+O
KPAc0l3u0DgGYXvpf5CkpODNl8KpiK+TXZyBJ5SJ6vs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 29232)
`protect data_block
6Ov+c+CxlQGjHHBP/VVyRdAs8bkhJgMM839Tt/WbL0SRUNmebsUtnJ9a1uCR8F9x
4l9MX9cpNOjf9RlLkRSGX8/szhoxMGSrU1nxGgVsTwPx726FQpihpxfwCgYP7wi+
MwtvE3i8GF0YmdSr0Q9pix9UbA1B5CxHS14LPig79LYQhr9gp9EEOZG/TUV4/pR3
yQ9Hv36amYYmbAaCDIAeGbPish9RyN050M0gAeC2XUZ28PQsoxEKcURMj1+r3vGt
2SH0dr2dvjlJicS/k6xTmVnDkQvJrGIU4M1TRhRYkxkZt/nhuKHa1Hv4PbMa9Y9G
OIs5Mb5P3yhZz7ruKg71vISlq/c3YRWRBaL8HF/WuQwzVuj0/gcQdyyS+rAr1ln8
qbntCkDCH/X+3hLXKN9/who3D+TiErDKsBM7Le4ZmR0qAfB8n3d9Bcvv2v9IgeAQ
4gKKH6mMLjnCt9i05PxfwLyAlysuUMNzydqvJaRF6+4dytFXLR/C4DsdBullBmVF
afjfOsnwP5yV8kgINOL8JUnEnwUbQjInpxA6PVx6xl8JPoDuXpT/pDRbXwo8j2rV
aaBtgl7+vBnzN1Tq8yzpKFxhgYB79iP6XdRf3AhvGFLb/3/OXFwyxKunw8IL1wM/
ITb/zS4ehhHynKLx6w0UOU2xIFc2wCtagRyFK7qHoaOpgyHRSWeZqvhq2hH0ZQZY
OYdQdtU9XeITYoapc1w9SBe9TvusW2uXai7s0//xYukgnZ35Im4vrDSHE6sPcHz9
gYRDXg4KpzJ3Rg513AtFyy9r6qdZ+AryXb0WbRFK3yUU7xRVGPqt8c29Zo9xKVNR
PwN4XpREwsSyaJ9B1AVzWo6wUvatzJMBql/Ar6nePPd17EeEU71FARMwAgeJwjhP
PI6CVcc4nWO28c7RPQ+Afe3Gfy7P5xQpHEaqV17k4dHHpShsCN8k/cQH/QpxSVtb
oNiF5Fp7Pp9EtORxKM4SMoiG69wRk/cOI0QSGf8uDLfbDOL518aHvppAIFGioysL
Nj6uqnOwhRZZF2uwKhNfppxKmDVZTo1dDHp/QsdFkwNV1XNpdg6JjX1SHCo+HSPs
F0rjqjaKur5OWPZq8NBoOobHUd76vEI6KZpCpCLU/78ipA2o/wHwrl27zW0OC3D/
vPltB8ly02KOqgR4Pdvf13EY3nw/g0pbWQU7ooz6bgN5wK1Zz9vv8Z5dgwf5X6vb
xpvCEtzl6LlebR4rmcdbbeFKRiBAeNLIJfRU8+9fgX5JQ0Z6/FXgDVNrE+50q5WI
jTR/LWxk8mdbQJ2taKPfiLfa7ycbMRp3fnVmd06xrKKnOdSthpK4ZFbT9VDUnuFQ
qDJmE97CeZiK/aRk169pFlQxwfeARiLm1zbiwGVqzi92mvr3lIQtWfPhGtXNVdvu
A9CD8k3xvvnjWVAk6vTrGtyGdQFCqFrvIsYdyiHGaa44r7U9v3ROqnDdpkJessLk
9l52svmW+fdXQ5Xg6toUtAwxZiLBLLBD28yGc8z0Nl79SP4LiEAxOHYfXun+yN5X
DiyuNJUQST7QIodnVNbj68J1mOh42kDTfKIZZRQ8GRuy39PsHyKhUmf7kuaqQPXL
hI49pK1U8rnBca7j3SlPUimD6YVO95A1UhhJtCQaYt9VtQvpfbkOhO97J3pISsGy
wbvfJFDyQwYHIemw8MnM3JMqtXFYR4Jn3hfp6w70u1kR/ZjlAvHAmvtz+EeIm9uM
AUv5NI+8gR4BJBDicTXKYp7sLzoorz3u1/gFJ4vHu37UMpwzn/P0JgyPrNdZYEMu
trN67DdzRRanPJ0XnE+FCkuVvIYEiN06xgCkrwyv6Zkv7H5f7rVKfbF1A6rm8tO5
ZIP53NU0OqdZ9rRJ0h+R7fWbAPt5iDoBfFFHqna1hGqkDA3Uj75KtbKVUF/vRPxV
mHlvwxwyUSb7/RlijZ9NM9CCz7hHvQH7mAKEeO9QtRoRj6BzCF3uJ1y3AEgFo+NZ
29RIvyX+O9yQMhqDPeXwK/fk0qyDaaEiyqkty64slPJYCAtxUjsQjOyrcA3cMCg0
hvAQXl3f+GZ1HGtKV4lc0bumgrFF67A1vSORnxyyUtwN2JlODZludOhq140D/T5R
sOEoyQLPG9WaMp/xjBoBDlA0XpGzkGIZGSWRYexqwr0JmuM8Kb1IrtFtSDulicAD
SmeUTevGd7VcltLx5HqEIz1ursgrCLPRVrT5IQ4orhnMIO6AIUB9coUFIB+3p+E/
NIw8vWwcqsjShS/kOoybUSFEcw60le/+PuKdiunxu4QZ0EAVtu8SXyzk6c2JznWE
VkL4eitdbscXittkYs5WXVWdh3Zk1RaPvun5uDqFjrx3B4xSSZv4/FeAp3tLkTRW
H/4Xk8X366NXPmaOa0WHrZaiTHN3W1J+26kNnA1yYX0Lt4SRIcZg93zgF4WoyYq4
GAI+1RoK1xvDuIuxyH4uzA+RdM8Pah6RJfs6iaornn7UPURidE9ps1lbF5hDDTMy
3N6H/0e/86TMDrtuVS/BRHOa5lEK8HL92fNAZMQppv7GzWHElzHlE7HFSH7JgIA+
/CYUBlg1iU2yRSuHr4SMIx3fTTf9CwpBNWyD8TfidlP2OXEhB3JOIPoTfRmFnXQ6
MCtR/H8PuAhddGD3eC8QAQIbOrUuFp1vafwPbHDXi2aaiOeWqGESgYRNrE2lh5So
AHEZLhjY/E2mkkomYvcOw/AseishbosDiA2BfbDsp7maNb9rkqz7XiTJHZEI6biK
WKFp8ysy7enz8HK4R8qowRU3WPus9t4B6qsE+Qgyj5/pdQfPJNAER7EDtlwTnJgx
t7VUgM3pKvG0ftOb2xKf+T2VyXRKBDw3K9xw16PFzAvYqM15/4NCVrN2EFZAyCOh
RD3ueHumU+i+9yfzmrgNQgEZrbkxcG/EwSMkDlt5VPN7lKzVz++u/mR4sAoZq1Iz
CK4cN59f/jP+He0Erg6BK1oD2NLRAkOs/8+PnUZOCu/AsOEnPl6Kac6zFvcxfrQB
l3aIdYzt2KtgsKvIA6NdDgkX65Of7hBtoyLZh/w+Apuk9mhrB7jEEgi7FqMjN4Bn
JBUoB8L9u8yWngnV/vbwmAMLzUEbZfAL9UMQm0SCFc6eaXJ7jZ/K54LhTDgsXaxy
W3ahgE9DqweWIVJ5Oc8PDGv9exIKnRTm7UelRso6xmFszMyr+DaIOXB4Yubgct8i
XU3ztW5gmvI1vpgtUa8GrOQSHTPPjPRlMx0W/SGxrIo5NydjDFQImTe2P0TJ+TJs
RRUAu6tMeS/eqsb9qEJXS3Gc3h3oJpDpWNaEgC+zWVbRwhKKdJxR6IRBDOFjJBo/
n6/kJryYaw1g229zYerD1eK7QzGW7GQniojFcw1MtS15hJYMFDrpqwCvTLNkPrzc
vEaVyWXIGeYMTBjcN95na3yvsOZ4f+FYnQbAS4sz5IxqhCNo8YmRL8XmpLY1hNjW
qaZN7wt4QwHqnkWbJCi3sBCxnDtXKBKDvd53nYNMw6/yw02C+JdHuvGZzfLgoP/s
O1HyVH4AHsJqsJuWtjcACUTN3dJD/ttm9/PZ5nwtr/fSmYi5xm7kwhNrTlkMBpBO
dpvgFI0d3L6euwbzj023nD5JtWN0UNfyeUQdqWCr/sB/6r8JJ6LtzfasryIHKcgs
EZJoV3Xz8CISwN55IDQCD7MQ5OHQrclX42BL1fCHysfmF7a9WVMrC2aW9Ij0p0lo
I38bMQKU4ztMYklhODRcOc3a97na7AtPZy6cf/zmv+0E8ByEx03Ew+arYSvqo2+J
iVM3ef8U4pKTUj9MnfUnjLjj1xRjSSx3sKA/Tp4a6d37R6ZUR3PCZb+oeHCfrt4T
QNEGqan1UeQX4fFP2KCRLS7gtjiKwshvI4TqoJak5pnVaVWfRqwa3HmMDy9NPFOF
N6q5QFXhBXOcqJeUyMZKGOUTHEkJG/wpFzJqjQwFrAv8g4T4Ih+BDOSeOPhShtGk
U0Y3920lkeImZFpHu4Hxk+DuoBJ6iVw5XP10f+9zoha37ngWGKyJPez/ZdyDPa6/
C31gqo9Jt1m0QuN54vjB4cEe0v5mk/8i4VLumTSG+uaxRGVp5zTFtz1HoRAE8WeO
bZ2Kpfp14kgb7Nz2YLfEJgT7i2VQ1Zy+t3+MkKXg1W7j6OwvW0bB36Ent5u1uWq4
lSWXq9VtYKyYVOz/yvSsnJcYeunTnGpaKjnDGUIHxrOb7b8egocIDn/zwqP//N5y
uma29RQ9RPyjZisX/oPvtJ7LdZoV1OpKAaFBk70kKSBJDJysj7cQCy7hk7/QKUG7
urHgY42O6Ac93ANqgOetv0lrxf515HG438RbmqduBF+qqGL3rCNETAve2E4styjH
8jop1sjj0BfPs6VxMlhhdRWaeK0G6qcHFzsPWjnfHrEFU3G/ZUTGjF6vQTak0y7m
ePsl81YtyugusfygJEtv3kp1qoPiszFpvVF7wWV55gXEusd0iLMlvSXD38TkLyVP
1MHN5YvcmQ+ZUe1JrGQBdo8uvJzDpzd0Qry4EqxGTZ73JZQNOYvibYIn3CwzGYmK
Kh7aMiLJdIRaLlIAma3ZhOIXrCoAysDl9haYUv0WltCKvcpXPhTxpWUcvL+yWyHq
nCVoJYE4QQ/rIev1colC7cIod4bTC3S7P+kzbWQpgZvSwecCSlt6e+/9FdmgXQ4i
JR/8NNtrI0aEMoN8CmtKy93lA57lpaA/AsTWNnpsuDgun4HZ4DGdw4GgeIsq8I1P
YpTRqnxJIeLl7RSe4so/qWI+o1ufrSQjicmnvgXSZvDcjIPWfTAnWjPFlmNb6VXt
xBAH5DGBGfq3pXMXWMoNjZaDLfyIN86046cMM/V5eE5MSA8Sxm0/kZb76QU1Zdy5
RKMHO1NlgVQH0EbMzWs27WM3NuZPqul8UGSoYRINb0GqYNPyTDuOIsbq0bRQgSf+
LHyPf/wtz21P6ST2k5NGOC7Y2GT71cCkPNZGvXB0QobagxNGPQF7uW8zyYw40Vya
lKbbu5fbD1JVyphz6bQA02GttP1yIVAWWzeP76R8TUAmJlaKj1/0Z+tdz6t3Ktub
drOQ8cEJwuFWo9VHWe9WcEbmf5RLEwpztaOXhRBtqq+dkK8SFir0DSsyBOwzpryh
fWzquR8wkUgbaqn4SaQd4UjhIP67aJmvIsgWHWsp3YjU3U6KDLmHAIf4d5B9US6n
a2++N7jxlYQgZx7mbuNl4wjJBEowuL3/FWPu07sYqNwNS+GTSpGCiVPJTEEvuRlv
xGPn9X/3PydoLCu2PuEa9s3TknoW1ZZOHtvt2nEkVB4B0uGBKV3mEe+y4n0oKLjK
o4growwX+2qscoZAIt7A3Q7vXq+C5HDvCxweHdchQJenQMzknuDkBFlk/HoD5gDO
6do4kc0oWByBBPXYDRyrCBW0Z54J8/bftb6NsFEtM9QIAzR7ACLHhjkAn2tfeThc
t9uQuEJKO79NNgKvDI27B8qdEDahxT1GAdDrYoOVm4X4nPSuBxc0M7QTUvIHmPOX
uhg9T4DQh7bA/gMemnuufxXp9SvRFZWmTruf1k2KH9RpX6v9ytugp3VWK/RIDzFq
bb8vI4qODH2n94qd0ZeSANu9WX2feMREO3hXIfIK9wXWrQ7DjAAU/LGbbNtGdSJM
qiqJICNIBkzDsBn1K5LaCIfpVk5tzgj7of/E7uNnMCe4BKsLtJnony2pdbKXIM6A
nbEvXgh97gQxE+V1iXQNMEs/djiLw6WTf1ESc+jex+jjo710vv/npfoT+5fyQbNR
Ypa+sHz5m0F8ITWjJgyIaN62/EPrv64Fq8k6JfmcUXZ+UXl2P0McJfvmpvES1a/X
1XvedtgQoDO2xW+Acp9dG+0erlmfN6EXLKiXmxePKP55yIS0h17se5jsJLwlKU5T
jS4XTJ+dMV/48Cdm3xTZL+IKXy0JwSAdjPCnCBnHcrBuzxOzUgM8+vSqrKhRAmtr
K++1cbR5/AH26rv/hJf/fljfB8RGJ+dW7gfrjD2+jxSepvFMC4bO41z1uP316XHy
4z/SXfKJO5DAlskdYjGOFB4zvaK4mOtzhsDLQiMsWAHBYrw56IXLIVvkYzpiNKmB
OEuSaTDRQcvu0eaigaYg0M067x6Mv3fIRyO5x8o5qRJ9JEjLFsFlFiKWsbzJRgR9
77YRtMf89UPChb9HYaBNwM5X+PLhXcDEJXrYDzCB52xteXi9T12/WbtAxkpLZwq6
G2MLCoCBybXLdCTrUO3nKDP7epJgKOTfZauHFKzGdyxZrQFgN0DIbchX4ebsNN2E
w4aXN+7fYJdJ3ngKic7oKSlYvVaT+xKI0O6n8bF2HjRtZemgd91EbBqVLBf+7HWL
ATECJJGd0duPdNiAOp4br4O3GsMo8MgFkqy/fWhtvA/2zupHyHlK5cpF55hK4d23
ZEbTmEVmT6e/Tbzh9QbFBMs0YwoARUQm+en7P7gpGcDuZOzpgKtcyUxYYrt0vmhH
r2RAaFfLlftcK8h8nJsiqnNP/1hJgQox8vOh5zbLZILDflJlSfsYvJhoUwCgtX3q
926FEW/+rYdkKoP8MraH7OD+ZcPdAq8f6UnVrMVU/0baGWULOxCSGKxejKh8PXsf
er7SlbQkSsE4mitLlofTZKYPwVGHjCFwJSwa1U6zTBfUwLh1vhX8mUd5TeUi3HIN
NhObt/CK664nojq0B4DE+RtQ+mq0EzpOCSwDLqwlH8SDhy8Xzn3eeLrIeiOEH81p
XTG2aPs2JaQJgxYSnA1CObxvot2UosycChEwln2qQJ22+xfRt8oE4OVji3pm7DDj
6Ki8rnk1iOjlqtGaf5/uRZaz4DCz1sMyFHOx7cy+QdEoMOowknsSMPI6wUwLwi15
310Xt4X7CbqqlpeEwAInmyQ9hu9zzzkNx4d5W9whCr/xdaRig2LwpBhYUp3vm772
eDeE8IBO4in2sXG4NxvOW7eJIGy6JP7GieR/GmyNlpm/KFU/AHLk7LDNZ/SRJS6a
Kf8BvflLclo1kjWrHoSOXai8uFsYvKsMVOYoh0ufdV9tJ/vuYGkO2UkFk3fXZuak
XHTLkCdhP4RzlpAniSbm+5AWrQI0FJlLEqbBreOcc0DrOubEYEv7PHBNe2pYY+MZ
P2jv4ob3/vYoAYOUHqXbKRpTeYLVJjq1cW5gmR/d8mY2KB82Mn5FeROZnaenvGcP
Jv7zm9r1S9WBmUI1KlZVnBKAlWyEKKWWT4KL4RBLphk+hz99egEuJ5GIvGNA751P
csdPuDca+pNGASUVpag+XGfWUEZ+w/gaTMuOn1TC5ZyqNOKUih4JDv9shARaUB9w
lomnu9BPXC8WD07s7L9bvkv+zsN8iqv5BAp1bD0Jd6fy4vL8/WIsBDDyALGBpQPt
/ih5uYH9JXPIMqFq/kW8dEgnv5xLDBCP7x8fxFwhHvsDmn3xoMaxQdEY8TreG9jb
aiikmTkk7ffeZpFtFviFtJX235QkYPAwxo49pfKkKy87NKCnLHUilQBMkSGJp0ad
OU37syoH0C9iH4rnfBtrEXZoj524z8t8eFfOgvZudfJ6gFYUkegNhlIGyaxiUIPA
0g0FtAmgHK+8/DQGYwG9XXMblo8LHQMn0/CodCfVN39J8sWM9Vh5gyNakLu2UDQC
Hu/zqMcv9JLWuiq29TuEcFwvAcEhZ/Bx9agKrzr2iMdJ08Sy+dki24h+hBDkLumH
n1cRSSgLsnrDlZH/biv73OX2FPhY18WJVhxyVLZjtLJdRjVxy/ikgIkpdntNVlS8
1E8ItkLGIuj54mc3w1uYL8JqppM+cI68siR1KRqQAew961eVTEBUnbbZrZNiWiMC
PC394d+m2MfqTXze63q+vPMs3cpMcYPezRJYWQbpxCs0Z3g7LSccooTqKpiodge6
edvSEE1QuRL2C5hViKJgiJlAPyRPAY6FeEk8x8WNTK9Ua73LBdMyyDrTdbq0bPrk
dvJKNrBWyV+ZQNoZfLrzBkUf2cATGxI8GxNI3sANHHhXHX4l8rIAit/GvJ1Zqo/W
nZ6I29ycKqos08eii23pEYxSfqsZ8ow7oifY4r5AW+mg3TMlT1vs4aHX1sP39WSb
e0f6G85703xf9HjXPMe79BqjKdsle1y95hbmS8GAYObXa4wrzfe3WyriRZ4ia71V
oKujiw76nBztSTsYMRd0SnMrRhgIY1EFm9Nm7Z7cODhX5rRPsENFOxAhI5dvZCOF
EawGyU8D4tQCFZ4ffZpp2FajEGo/nlLh4gZO9mVciGUgcwZGK7auvhGSrO/345V1
c0BaKnz4rd2wOfxWsrYDYlE9AVP4w2gXKuxtqXSJwucSyWPPQnCYkYxJaNzEZKPf
b/gAeslFWZmcQzuHaldBtwdtftk/ybIqKJ5F6P9lIanrv9M+p3VO8IjDSERA6A7e
/rHVm5Ef+2mcQBnqI7zrUqRU0mDZ6pJqh5T9k+iaRbb+nSxW/4/x0+daBOoXrIxA
rYy5Uqed0cSA3WIv0EYrqVlRcBKEA3uqNKI6Lz8wL+SWvQR2RStbOVSLtsohgVLC
ikTbZDSboyL06mcVFI/yw62UlUhHBMyq/Zhk7+p/9k/hVaNGINqn0KAUCknAWqUW
U9hjYw5wfKwADY6jXtkIe1TgAS0ohhQvwuxBQosgzIUDZ1HOQdNPLBtRsNmloFtt
Pljqk69aaQcicM+cTn0LkaEGjSsVn3eCdRJ+0Q153mhr7qwI8Z6zqUmBSN7tTo7j
+Ec82oANFHM8roPi9W9f4h0W1iIhKjczzqHE7g1lkUyyPJXoMm1kgZcHhj4UoXOB
awunfdojShBjrql2H+CWkGGG52YLpeT75frxR5E6L9Nso6oMGpJrrAbnc1s2gq+t
BZfrnXh9FfHiIWhaBEtvRBevDmnmEsfZLR9PpkgSW3GEGQ9SlMNR+Gt8BOICgUR/
Av+V1SOQavhPrPH+PwYFO3z6Pp1s1qlF0l2ipsBOqOvqwTL6NO/NnGpw5Ed1yaVU
b8BxTRdUIZCpAlamqVIlf/FpI8daODAyNOYN0ghVd2gUEh2zZYCA5qzxHrU5m3WO
IIdcY5HFWTS+Kt0JfNIQPvSQMATv3CBez4ogpdc/rV0tflSpW7UnMU0v+Oy0OYVM
AP76q4kkSaHF76Mi1Ero05fId5WiJYghvW+tb1zXqGS6Ef1v9EH6Gy0UgLMnETBm
AXXVorf9MrhCXknoaVAUx1pd2MdmNmf99001Saof7n8Ha/A6d4nD79Q4i/sie71k
0IRImgVjFpa7YqVZ1IrCnSZlLyxbn2JV1Cq1CvDij9KwCEelgP/YFXxxRuD17X43
1hpAHRUoNcrzQfDV6sETzEZt3zqA8sMZ/V8twNxd4YWbqfNRKPbSqkqP0fRu4wDU
MJBoKCuGgLzQGMgS1Za0fAKJt5MqgWilugpcAn2gCJjj12SYuL28TFJunD9rrx+h
6/y+5mCCbnQpIaW++IIjVOgr0iGYSJyu5xeRWWTPBcaPtumid86wu3UcZTxpHDBL
rpfgsyYKMHS5oHH9Xps2jyJbNmHFRFa1JGz+XLJ2+ikeMdIgmzCrnWfCowvZY4FJ
HGgJlXjDyGdLfkJ7iF9L0GAk5agc+8sAuooZSoSA+sHQUJBSgnyQ7pN3Wem3caHk
lxK69vipK1yYeuEFih/qDYy5a+Q9nymrO5ObS2XgMhf2BIdnh9kW/uaAZiLyAgaO
nyF77QdIXhypu+5rDgHntoPhmtt+kH0jK66OpxzedFg3pyiIF0TbzVhx/SsCP9K/
sROCtXSaJVLZJzBGx/bGO5t/tgcgyMIZPUO6Og8h/SuARWsuEA0PRVNOwQi9+dFE
JdCcvFDhECDJtmF9CxK/X6v+coObaP182r4Vkklqqval+3A1a+bA1oPmYgHc7v/d
eGD3GJ3ltQ7YZKUlbsLDGyatM7ZUlOlK1xNMGIPZPztPzkXdHBL/Rr+g0FyU1roQ
uuQPJYPl1QXnBMnkzVhGMktvLzCygnlbbBKQMQnBMp3AGrJYLxTgvq3P+jqXwx2w
u19cU8i09w+LvKoovnGteFz9DbaXpO2BRejNv028AiIoX77Ag48UyCksl3wHmlxU
N9rfPebXJP/Dc2REXBbVEwwSC+t58Z+h9GTkO8KRL5OCfP9YbF0Jwpy8XkQiO5ix
PM/gBvKfB+Fefh1ieW+SaQffMrTUrJWZhTK5LnJpD+s+Adx4TNFq/7uWduNsd362
efS08INIlvRBvea7ca4iY39uaUH9KclV5vbo1PdAAoCN00urqDeSMCOVfMYOjwmJ
uib0WXYM5xqTz3+0GqqydxZozX5cWBmcd4GCid4LjSwu0uNaBDpgpOCA0++iaCfx
Yjag66JB45KsHSFsdqu5QdSD+1+Fm3LLz9ylImtenqS5+cNco8FPnvY95feB6mwP
YDT2O4pkbWt7qLR1AuLKZEq2eR/1W569JdSwDiEfS/jB6tWerA2b3JtGtoGcCp4O
tp8m5hX9GaCkEGCx4BlOe5mt5k99woGOOSnxl7Wp6sCKWc3npdorRe9mCgDrEKPX
qa9wijuhamK+f1eWWxtdwyBdfYQKufuhmCuSC4r2HbmOxsapwNOEsysNtv01X8QD
8+Q3ya2zhZRDiV41KQzD0RKHHbCRwZP4Tni7tLPmo4jxM2FLtRHWreWno0j8nrqy
Ld2OnHZZRP6tRzAwPNgO9a5i2eul46evWL6RzvwKtSt6WX6U0uRP1WmRlUKBK173
sLdfjWEcwu1UrU1zzuBqe7OF5oa7YpFH3JZlTZpDUuC1B+5cP04Snq3kYVKDqxQ9
WQC1PFWDdxP/RffTsDI85aedyXbLvvFvq6LqrkU1m32XC4POpKmSTP74nZEk422o
0bTztfnCa1nWByeoIOTtrA472uyw5WPKcHtNsUunHyx+4cRkCH9IMuweqx+uEbLz
hdbmPcd1v50zxx4fZ23T8+8gajDPi4EThQKn8Rv++pbKpvni/M6Mxc8cpSxU+pZq
sWehTsQGICs4ScpUw5z2dlhO4O0UlCiD1sV520u3XGGPzJrGrEyyl5rsWW5DQ0tI
dxsJKrpZDazUkUM2WrwSODrz2JvFlJ3L1Ur6sG574gW6+42FUS18HBUW5rwBfqmE
PCgCi50OfRfsmH1rcoMz6A+S5b3syhKHmStx8FWgCw2rnUSlepoEPJue8615dP7H
++7ve5OOGyUQnvycw85eCpqaPyTLtWyGxorV2AQO0CeeA26qdDH4CXFCxyCG1D/D
Z6HRgjeuvlXdXHQiQ8VX0z1y4kwO12DlX/Jckx3QWM9j4eg7Fvxf5BJQM2PNS0pi
6Q88RVoycBMPsMvd4IV+ziJJ9br2Hta3abK7/RMgjMHcjm2WfKAWZ3ByQguZxyCv
r4GWf6taNiFMzlE6Fol9lGQ6hm2rnwxZ3d6cDaL6MZxB+0ZiWCN/iwCPYm2vHj6z
7ObLm2WInmes6aIYVdElZuUeqg/6UjvJFXPlCBwTMlb/6nrrNwZvro/cxqk20yx9
xnf8B9wYEAxm/LFQYIfTDguAFtC+AXMPv8Q438fjWoYJQl0m74WA49Ex0OR6hoQR
+xHP0/yAHQc2qxwt0QDDG6JkGw4URWXoNc6STNhldvQSK6u5QXpKUeE2FzVNNq3j
jEjAYn/oF+gTjdQ8EezU5yoIgCMUldSyrKYmMwJs3lSra6zRBj1E0R/nYhZmXi93
o+4GX1PEUs1Bl3JfVBDvpCUwJcfyEOVdfEWGW3fyu0F9pzxdBo+e7eR0vSb9304N
6tGd+152WqdG5zjfe0S7RWPLgyudJYYfswhllm++sNZyOk8ZrqPE6q8UBpa/00RC
sWIKJ499G1Udgjx4N9CaCxAMRC3GY5OM5bSHSMp42wIKpGVNHaS1ofRJWpTskaFZ
8wnLlyC+JIRq4R2II8JPqICWvyF6wjBSsKLpP79KOU8e9nT4ULdoA8p8odYn6qmF
9qmPylO9u6KlB8N88rlgd/3Otb6ldJV86qUyY9HhFUou+Z1F1MgnfCnZaJyUUzUB
j0Bimg50/WqyN1HxtMQ9PmS33iT0KVa0MjTOPOamlL72HCRAt22KeW/udNZCf4jx
fI1sfphKX0wCkRy1Sv5mJi+KsjTLu5hyp0VWZsLtnAaHw52nlMohGZCjg+exAp0R
Sv72mlt6GRnI0saQfn/cTB2Lz1Gyx/wj5LfGvZfeV89i/x0p+tbKK5QWbTP8FhpS
9l3o86+4oM30jBUSuSTrP8lac0Y30YfO8riwL/ihIcgx61nLU5vK6x/1slG+TlBf
obyzxdL170L2Xcofpnsa5QD0gBS+QpYABUFCttA4h4lpkO3Z/C2wFM4/BnMT0xvF
+TtvbCWhm+JeDeS1eAECpdIUcRqSv4Z4t5XfUTk+mochhlwG7ySJZ/BgJoESxvEP
zJxhPP1V+J5LltNyar8qPJlIIG9IQoOzG/mxywV6mCIF9WjN3kpLYew4JEU9h7K5
DTJKOxDOUbn6OI2zd3/mRbkqP1SPAzF0aZlhcWpZQ6XICV0V2D0kEg0ZMJcp/LvQ
HGrsqRlbIeOPTN+5OD/XWVmhiZ4+qIlzdB0PI0IdDZTgCCYPjxuAx2VlcgXk3vCq
aW74e4ALzUpxs0ViBPfICDPWLIsi85jDIt3PE7xRn2vEd5uXSzY3MUYLN7Mkc5JR
vo6kWvlD0O9wnXU/LNgp9A/BG/h3/C9bFaDR2RT03peFwDWIaioT255urV2Jrt1K
+aHqbHyv4CYer+G9LmX6LIzT9D2+obPWx9bsqynu+4woqOYiAwER9yCzqIL7JsGl
E9Ti2eoyZWwCTPJHn2vNGfmIo8tpWpWD3jDgVmK3104HuL3U+LnLVeBwLCRyRlz9
dUIrvq2duJuuh6IpYjWmrEOb44ZuOjhzZxpbr8NwnNyxkoxP1UnzrhG1EYoQlgh4
U2c9wTXZhhaQ77FWk+xKwI58T6xZgV9UzPwoBicX1pnvp4LOWiIUri32U2vbeGUc
jq4DS8Y63pGlLFl09bNzAP6O0qbdXXv5442PVEwA3ejqqSoJfbHA44K372fg1EiC
yxp5WIuXbRTVmWeA3imRjyGO17+9GeYpf0rB6LOMWXAAg5Tbt6WScXhbXQX0riDE
+lYc+YdkBa1EZ59H3WJ6b44rsOBkSp/05C8vYjZh+J2NgZhQJNWTVm/gDNSUIfWO
cw/yLIK2WbgyUnOeG4lMkw8Tld1fTfVO1MocAQfAm/pCFicnNBbOxy7g/wBJUyHP
AOq5JNz/0tour5yHuNGBgVKrRdb2zXakBDQzcm9ZIfHfxZT2PUTQhYR4JREvle+y
pAkI/UcMwME+fdAVk7DIgL73lqMxJHnFaxEEmVyif5cAQXW1GDtPuNSXWCJNMRgD
CRpxvENTeAtCIQ7I4mabRzz/Pu1Y9RE1JVUNs4FcZd4qVr3NgsXJrZLhoctExkX/
EMRID3VIVzLnKohPt7nYFRlz1Z2UcYSBcVtt+8hkd6muwkArLXpZjhiBkMlfLpNj
cynZibj2qfZEDmg1YvObEv5uJkmsoTJpaFYQz4Csx4RZmO/5w5+IO994eab4TCl3
ALhVr4K57U+CajMWVbFzDs7DcGu+IaBcgrarU0sQEbDFcP1QYCV9WK98UoTD1q78
0fVCR34ShNuIN1CcBsfEAtaFxb6Zb5GbBJp5dSJjoR1a9QakjWzSbzKWYIBBydOR
L5NzxyQ6j2QTK7tylUr3a9N1uyID4F0HmRH2aM5SACV6v3K9TELIRjrtm/ZhcIK9
yr06/ZaKmAy2aqMNAaZ5SxxwgB1nlTzSdaX5sZXrJLxBR1jNGr2x+PYK5agg5DYe
x8VZOq8nty18Pks2rVVpptQuDISPQDB2OzYfIvTN1o58Jb6GWw1GMBtQRy/XE9R5
wAfmnx3PRBdnT10e1BAKAGY+0Ct0qh/0T1N8SU9l+V6/OFOdVm7Slq5s7+5itPSn
FcWW98WRYKyfYAgicNU6+2S47nuBrS8P7eIBZQ2hmh9FZ+QCBHWVGt35ltA0bXCb
TOTHgz/HadojJ5bRSMv3sJGDAk3kqaF5AjlJBJ0EC+KDW6ACmTMii+tO3WAJ5iEp
pBF8qHZtgmLpVbpHmcjFnkWgXIy01EtkUvZV4ESB/xOsVJNXVK2XAMKzZEng9PZy
y3eyVn5KpD2DHVWVrpy+RQD8qKYoDqwSr+H+kJQTKgo9hAfu/OyAY1gqa5oCSfvf
5WrBHHC7oyfS/3K2NlYskPlWyduBEpSJkIaqtG84kjMV2vZwNRgE39tZ5EqlGPPH
dH/aV+uUgFXf0u4vUtUJ1lmm82vhNnv2OhFKvrDKkfsNlO7YYv6D9h10b/GhfKAa
0ZO880zIpXJ2UGjdm/8/n1fyA0W2AvbrIBW2szABNMWIi9l0e0ikT1tN/lIpzkMG
j/8Y9eIoevNJ7ZgDoe89atJhb0g3Vhw5havawgpeltDlrl56GwAqN4WnrfLPY79g
ptHAFUrWaNso95f73XSDW9NliWEcAYJt2fyRi8tVCrn1uqZcGOa0uaahZb7WT18j
9GRD8W82kxWyVVw0RkiMjFF3jB0dS1eTN8sT+ZmIM09AYwabjM5wlV4Bqol//Y10
OfwVJAIkP3d2yPEHgIQijs+YnNy8rGVRIseE9ixeunzHdJgS4cmpcivh/KtmY+m/
HrSJHeCM3Lj6yEc3EGakvBiEj+HUJoalNhH44Z2rT7LVBCRRmGU36SoKSdOFyv2+
UzpsFHmcK8LmUvYJXfdf3jjwp9Xt4ZDO5Ep6+msu4UJeqa4MrVQAa1gCwgYV6b80
F4hOokdJK5GB73/FhTHxneov6CtF4DXiCJtjIA5acFxavA0AzGW/kOl7WSsHCetz
tFyQbbU4gc15n1TO36HbcGHz17ShHf5odspBTehz7Ci+wcdbW6Q3BVwBGmx753Qj
CmItydU8tWnYf0+NA29qJ4bKIWiikB5nslOEdx0iluWi7IcpAer+5uEPMVbHmwsM
C5STN8r4a20Q9gRZGNXmE76eZB3XobIsD8xd765dn1YLB/GrETIXstgUwItUO/Rz
7EjEi4KDy+vgInCAzrhiC2iHJ06X7EDjOMOiA9GqiJssPVbB9yPvXnA/vPWCA6R5
szK/w+JTBdbe6Z1b7tcpOXDiSVddsN0cW5Umzrmch2bn8pxpVVBYVzFyYyHhX93Z
b15QIiQG8GGKn6S0OUnl9MymF50R+sl1vOKwxq9QS0cN/+CufSg8dT+iyWbuLZ7g
jhxcqOrtIcomx4gACYPg7NQqHIxk6MB3klQqOUstEqQt5xLbQqENWMYeQZuici3b
jaUL9F5NmA2dM4tD3AYQ0lEQVdjhqnlxMzOxpBVatOjTrOpI5Is/SzzPzVuXOQ5t
7CGvbbS3jV5lUpZBOIG2kc4KjK4A5q0tMHh7I78+s1xusdScvI5eoTgAFU8BfsjP
DsEiRqUwjHzDjElO5u5qSWCsmvcvECs9XXlXMNWqf0UmTi8O+y12zLSpJU4f81np
pdrZUoyH/9XYNIjMxPnhts6OZtlryk20wLDQeoh/kNOkjV5zyFdfPlwqY+bHGl5S
A9jvV4VdnIIumQDsFiFwjPJXEyvqlOEE0odDjsmYj7G3qq25DFePMHSroZ6+YGJe
VMF2N11E0X+hwPbwNkg3rZrVxOUcirD9kCDC0TmCGHVhphWkFL0IUJ9igZpmlytp
XKsHfmBSaDb7KlWuDdnfZhOFsi48lc37s36cdXjWHaE170qLHIYMkpRnUx29ZO4o
wCNkJEFEE6wwBzjsJkvVWwYexKY559OLsJ/ii33pNcZ2nsCK60OCLYa3BuDdytXr
ayASp/Wpvfo1fOHRJMYm6qUF8XDGjTjpLSajLGVEllU1c2QLgjW9sve2X+V19kI+
HQDf9DdiNd8GgK8RLgdkHdVklfzi0RYtUrqAgTQTHEqSIGij2PwtE5FPli0b6KZl
VDe3NWf0adCZuccvMFSfWjlnu0bNiEO7O2MHFoZc4XkzGxKMGM5pGWyEGAJhidoP
crO9H7e2uXl+9LKj6vF5Db6kMhuXKOtJqqI5Dsk5wJcjZ0qvXQTBWavKbbTlXibT
VxvNBZucr1qnSpX9wk5Lwl5pUCagSbwJR4bhKr6yKMB5Chx5KJ+/z849Qg9x/m3d
sDKA2N9i0X5R2brq/vaEJ1g6IFTlkvsKagtrq6gr5lIak7sRutmASX1L8JwLkF8z
b9pat66SpD5VS97jkY8vbiv3rU4uWkvvhBV9WFFImX0/pUXqrtZXDeoZ478CGrMH
W7IpGbxRKtoK9R3E+u/AchIB97Ot9mTrB+KCB3IfPO5/ErAud+sbQmBnQwaHi83W
hbq9Ec4cJQFuEHp9RyBivDEzaFTs12qfVJd8eqJGGoaiTH7807I+C8gYmKll0bql
JNrlmJ/AJFRDk2mubZ6/VHRqSrnZeYvX/FqP6236FAUiuNdFVFHZTsjixmxraFwH
xcLgiZsKeS1uegbF6ZSSsuJG8/6sOn6bXJNsQWXi6FDZngj14l5vzxRFeIQ2ml9Q
oIcZMX12xF/b4AmuA7+aA4FOgNkXuPUJwOmQU7ctCQ5eVIO5u8bUw/QfHINyvswQ
JoDYdp4FclGw1RwBFpNsgQ5ry/+mpjeIxdzMosK4sbqVMR7xgodLg0zHWKCxb8ik
oBSwC7wh95alxcrwqDUfBEoVoxhnAmuJFrzmriapvY4BXWPLrNoObcLXRfkKNqHD
rXctkOxDXqFxNWGIqPy5uNkNhzWhuSVfYtHJgIoggbQ8kpO/5q9IY+8yWbyRcSjW
3f3UZmULlG+gwezt8nyxYVTYtWt1Iftc9TUTxjdXVGbHZVSAyWPe7MJU2ReWfOLY
wNHozQMixhuv+KtxW6zSG1khmQY6BZBepfiBelwnXJSqJFGHtUiyITa/s61TnmsZ
p+FK5U7ajh5HfDTmIxIa8UOk3HdctjI8IAn9Ne4nVWRpq8ZH4mwZWIcoWSqFxdEr
vnFAwVGuNa1ewpKqhlXXoug0sKZmPoIcHWuXiZAxSWao5/OqPXj89dUxQIAJXvx3
zORGIS5yqs+IGfwct90Z8SMkeal6PQTpcpEVplodaF+ZDZXWF7hnRuAeWydiod2J
9q+qaIscTa+fqbYizLH+2uWIyMNKvdTnq2zzBM7bvZnfnJGeGCl47ksatEBL49tZ
EB7eH4dvoEYzoVjXQ0zIbxkfRgOSbAxE1yuS1dpyOtKIVs2Rxr4UYOc7lnRnwSSb
j1D9zpjBVue/VygF7brY+3wCblVNokbvMap+g+edE9F7D3ZyC+I7rAJHKvvBczw4
1lTcLBIADlGOxY+NwK+DC03PKLLeUT75Xve9mTRjqz9WiBIdli3OvqQ2I8JsNp9D
lYTqCuZ22tUwHqvjQOcEV4udM3xFfLBgLFJ2aq96Qx/r17vyeXf3i9RIBmeyfmaV
vOoGqD65RyDZ4Jc0sd0wD5MBT9CdXXgODbaLkCkBZHqcQ7TS5Gs024/4gRrydk93
J5hVZUXlAOw3rsXgp+5E2OYjD6jlP9LpmhGMqjV2YXPPqgpDsGfLayTs6U3rm6dQ
szy7pgV0at0IwvXZVnfhQK86e65qeIvFVJwetKaW5mUpC/SODowcP0XdP2LCD1GG
WdS8oCaHe+LlYWRralqYvYEkesLLw9VDVoZ34QZi3x8CjCQRk0POYvt6IdGjfPeJ
zmQBkBUe5hfPEx76omnH+rJjEeqWu7igT8vC1OX6HrbEcpoOhTYza096rKWazM3D
bxsConlVzNGoJcMhnZV0dZ8SZ5cUU+XNuFSk8/yr23BH/Yhl0Bf+qAIdbn5l8pv/
1IGPlGuw2Y4o6fiEcoNDaPSKAGXfIddpRPHx59Tm4L/ttAAe/qk5gnn8FAEgd5lO
4Y4fAp6nix9yFJGxKULrP1f1M2yGzpqDvckcCoHODbsVQfIZQrKXRbT5m1Q08J1r
rSpj0lEA3w3PbkpuCfAJa/rxj8868AhMiYwMU6alPSorR12+/Hnhg+Uq26lrQVgv
jecUCNtdM/pNxOrEej2duvIoOyUv6SactBrzTLrdid7cf4gAPMN9it4jwU1Pkl1I
f4VpHoQ8Uo2+aaqoNFAKFPjFy/sU4KJ5KMG7xs5udPsFyv7JFEwZoBrPP5FiIj7M
b4TIE1wYfe0T1Cv2YoKP4nGjZzs3xgGajSotxSOMoe+/HbgQZyB7YKCYHrWCErAF
vzR56JE7Di6fi1S6pmt1d+A+Vj0ZsyW+dPEE5E74C9Vg2pH1Nop2GRnkXUbN1pzk
bDG0psGUKCTt9JocRVzG5EjLYlNCxse7tYVinJErmAfNgQUbVzXTKklCxsr1ZGqA
XpXDzJkXQwWObY+1vMR7SKXWDwotDDyB28yUaxT6KPTZoKEvXPWIPeOnRAK+D3sh
OzmH6OJJVBH/lxI0lLQCfgJ27QfIF/XxGkObhDJjhs0DFYlrMg55gkU+YyCxE9X2
o40fD7r0ekRznRzDZFCg0kGJRPklPmJwjKubTEzir+oVQm4IYu1SWChgTKpIk7HY
O3du2n4ssqKdW62rXPs3zqyiNsykhoSXSFi8cABU3xok8vMtYX0Tb25HHyxJ7P4D
GnTS2G7hpljr3SCRxGodZIisxj4pGgeFFZpbVEDQuypolCIbwET8G7Sn5oyRwbhw
+GBDQQf58nMoFxGj2vOVX8NVUvY/DOV43FBpGJDyF9ecSnrXHLwfAnJ6SKQt5dCd
UnRLUBIK381oUtSQmUu4BaNatYb6NnTlXTkgLFxLSNhb9Cd66owAtfPO1BptiXO5
xalVvDM0vqAaVEwn+xxw9Dp6yvBDzClkhtpEHPFLWAhOiFIq3aAnQWzYYD9TMnUB
Yd+6dNTOSCgoL8a3jbsC6chzPp0sjW4h9FKICqrT8A2O7Cys70G2m7on5PxpRea9
jYXThTx2bIl3OLoVTEgyPdpdEV8+snEXf2HHU/Wx4krezVynxjdWBURcqzOpW1Cy
XqFwLT1I4JKHsqWDd2OAeXoyMCOSoG/SGr77Lw8fSVIp0Xkxh+HIjMOxRiK33Xdi
eXkSlA3Ff2cO7N+Ez9KMbex3TBN2QWXW583oGyvdrKoYZJODlQE4cuYYc8aXerkJ
yONFR/ELoEU5HpZepLwkQhlD35f+qTfQaoDXDm5jvEKzhC8mmw7fk/iIybRczlFH
C4mw0JpneO48jCs2fNsr7UyJsUDY4VVKXEEGXrBNFhSGZCfQT3+RBLw+wV89gMjp
jpVihbCCDT43i9Ln1KWhSiVeoiAyzPW22oCFoZRJ7iDU+TSDOszyjrdwQ+ku7VL+
s/uJXHdTNKuiUONienRzxXbv4o3LuN/Lu8vIVv7yY/scu/znZle+tSq3/782/oJh
VkHBWNxgFi2tKItTJ8iL19IvgxplD5NVk5IfsSgMgGslwezM4CLTYWox2xsH2neO
PH3jPoXm0JDb+MhaPnDWbAgyu4iHDybrkOdAYyPE3514UOGbbuClM16oXhj+RYv/
fst4njdPwbDh5ObD1ECAnBqkBOslC8VEKgMTDvpdYlb3vExP/kZ1Efqv/AJa4mzV
3iZbyk63ToQRN2wjNWaYL5aZ2Nzos60+lHdPCTH3zEz7mv757TXd+Ll0kQA1kwJy
YcsyxPppT7xa4KBYchMy7OwaSIQHTsLiL2FGEch/HXAEoWns96cZWebOUyzUDWWr
yQewNgkslERDBxE0TeHfuDxbH+7pT64QKyPc+qCxCzV+MCi712QK2dd56Ts1tcwS
VxlzCJgZBgtSK1G3pr1Cv0DBwpaOhUn2pjk/LAPPo+rhRfPKIe2HK2BgZsYoUJX5
M2kSg0h0g6Uv9x0iiKNDfxTndW8Kr9DQzohS7UayYeo4ictew3h8NoGj/JHY4uQ7
ZmqvQmq2wH66bzrORqv243kCB7OoVbf5h2fMTslg/NBHGNsVD1JDyyvazkZoWRnt
fKTjxWZTqpO62L8fjnt/YLlj6ZIB2o3xu3poZo2+iyX1LzPRfCPtAfnutmOS7ABU
46+yCa8QLMb44ioWMA8bXGix7bHvSmitVEVJg2NuHMY2ec00O9dnqx8ODE7AQvHi
1pe1P5R5FtQZKAVDR4iUleEoWDR0py7dzDeDB3KjLZKiBhCpnekB4qWY6vbUUATx
bfJptBp0KcNFB4Me6/AAqZMgGmF/X7xEcyvFpgyqOVI+2xtzQ3lIx88pIlgElxUp
uA5aPDPP+6mAxi07PXV9q1grRX4uXJhX6Uj6PA012XbobLgHxWTJvmXojY9aw3jN
vEK3By8jmM0z0eFElrjTXjLld5Nx1JJ9A5rBQSxX6pSOVu9Q/5+Y7KOEqfqBxDF7
C6FyuV/dA08wDc8AMq5Otpo8IzHoWfHNX1KCMBvarR1vj8XtuTi7KPE+ZQdwbTWV
vEan0c2CZhsmd3hKF8bq7b2j3Qr9tv/F8FjmEirKW4IA9Mb8FkCqyaSMFpgL92y2
4rvWTbVqU3Fss+jgRozPTisLD4gav5/MXLRCPfNYL/YoauLZwN63vNpAzvCV6Ld1
N8Y+bHvUYFVLJa+A54Xp3W8hDh235NuNt9vlycHmyvq+IlB8Vzt5Gd/7EX0aaEYr
tqu0aydxc0wMblXLua4rE+tDTDXVajrG8DVpZupjAtm1JgVAqho183QqKLutWE7F
7UBbq8aH9Pvwrv3Ftq4yFcf8TpOLhzXm+sjlNR29pfUa7cq+XJOQJNrVPNUf9Sfo
DxfrOpODD+/IbT48jqHwW5LgI1lU6Gu62XkKlRQd9ehinfNFitu4nYpE6AFqPGoN
VMWizrY73z497pn5B8nWCSHlkvUDpq1lkTCa6Q062DFip+bkndUub5pNcH/u9xSa
X0xYEu9+I4IoZZKVSdhwK+2+dqzgg+xuUHgKYtESbf8+fqhkLK97aBF8k+jAk/4t
vyWhh0wGVZjmAjCRSAFTMGLc6YMMAxzKxQ8Bvq4732q7GTQxSjDdXlaEwPV+uSfW
AUTjTT4SvPcn6cWaDGK6abh23Ca2nASOrfT/q6HlTr7d1eYTOn4nTNbGxneex5RY
B93jgoyvqnD6O8Fz6AdUVEdZV3NrFz0XiA39lvBDYncUEIfux4CGhGbSTdLR9yRL
8Ycnq8+wt4xHXQTV3EG4gdIuY8QFn1vRNo/LisAuQReXZjWXd4d+d10mENlZmP4Y
i18y0iaYBkX7Q4AiheWkf0CTPSKkWriA0N4iMYUA4TCOX5rLK3pSOOd6Ss3w4Z1/
00dxMQfeluEGEIUOBt4fukDJiQnZSWbgD96krw2PmSZo7kytOA3yy96lV8GNOoku
SNL7ImJPbUkYCOXVRuq8AujtQAhS+hoxzbGl/ooZVnJCLzK/xc4BCOTvfuaBgLro
69pojWsPm9POs7i6Y6r+EODAPRHDBgHdmNG811/loQyJCwb+uG8R8ntLpf9y4K5b
7V6nr+HLBwV+gKDpk3X251tKZx0PY2pZ3rFTHOYiN4NYJHjAmhKU5jQgUPIsApxn
xs/rWuO5gvi94Tbo8kYjJ7oR97t61hgwWm8ovijeMaI5U9iZdNnK2SV8rj5AmTo+
xpH/MzBZIkJ9VybcNP8Ty0uoj2SNcPa5pGN1swAPfdbPj1Hvl4PBcB/wyM3w3HEj
0nI17SjVuyDD8Gkb4aKap0A4TrEXdvWR8+6NBPd8s+CcDbYsc1VK/mG9OVkjqund
wanNQ8ctKdl+lBYpi4s2kfEszHRZrxrBimNds3LQESc/k6rGc5mqur2g02Wbvm3T
d9/rrEw4qe0zuiZb0WKSn97JO/0wajUd4CT9Z/TXhmZNa0D6gwWA3Xj9OVW7Co+W
8Jk/L0yjxhLkUonoTqEWSlZgNE9Dy87pbYqXqYMHWUml/9Wg28he2SxsMlE3ImtW
Klrf+erbB++heisjXX/ycEyfES+IM7BzhiEWHsWIsdTgmOFsTKYqkkSALslrm2Fm
zL3O/cXkXE04eIknYg3HzRD6z3QKX1rH3BLfvusHcR4iNj+r6jXd+v9uUTHsAWfP
NvlKZT7UuMq3ypNte2b0bmhvTjl/p/sRZQ1EK1/NEAx/M/dPFCZznRVsFW0+khe5
cX0pEwyQ7vD4zJ9okAGIZ4tC6vtlygqJ2IOs8UB+H97gRxhejZcBJgM6gCyNQpCR
JvLWoGMzePCEqiZLUWDexqxZDrOPE4vUq7sIMfN/nm0h9mAieozlNv1GaDxxLu99
Mf3mXSS+yJtRJiwAYz4pLq5vkYtqejIZztjcYS1aODU3AVo2y+89HnVZWDixQktG
K911tBFA8JSdVHiR7h4V/ur64ri84LkCkG7EqIBHQgfdu4PmuH59PVxf5c1VSsVV
il4PpxtTUNgh2wgtI+X+9cQZqZBaM1s5xWaLY8OAxM6pDoOBBv7UoSF4mA2LP9NK
cMaJgggxXaSI5xym3hs8/YHpG2FALLfgSE3qECPZVHKBcqY1dgAFkt26RKoAu8KL
B677nx6AR/gW9YUNixDh/Sf/8e2d5MDCpOnacZdFSarPMo2yjHucXtp/1oBVyKiM
RDM41vheHf5UaSThfNilwaOpvJEReFoU3E6uFDKsCIyb1vD2i9f3WHqxxZp32wht
6oOuiG917kFppUxMuEg4yO/nx7ZS34LKpbP7K02Lsxro8FOky5iwSH6mLhSiPz5E
G7uNZFf7QQmLnilGf8mP84hbYQAS13DbQnoFfC4lbKPbrKzxZp1S//5Se5eJxYqv
0LZVd9QVQTO8S7gSmDtvvXUAQyg5Sh3b1Ihz/QHwD7d6ciJNzNtx+z0xqu07oUlv
h5OwgWZRHTFlik9qsIXnQm3PB2l6e5j6GKa+2VPxsuspUaG9hm+vihSYmD0jjvV8
N0eIekA0x/aFSopcu3e7fYOry4kX8beeY58oSMCfn8kfOJEQLHlHVDErK8RmfjiH
e400KPawHmHSfBlz1sNsTQBFAOFhjyjmbvQMXzgcOlByfB0r5/OoxItVlii7HY7h
c7LPWzCvH6t/ObSM4f8R941g7eLqqBn7fCXfp6VGGPf5Dz3DzqvqDp4WbiYU86ov
lgpv1MDmzRIlPwyLVt1CWnY2UOBvQgTyE5ZJX72NS4oDEHkh7+8d+YhON0M5H35k
tfdRvA0ZF3FwtbI8U2+Fqej6JHUrIidONDr8gX5RkcDuqyXJMghc7z4/60nw5HD3
KGzA4CAW2pGUOGw8K4Hczv6EC69bsqABQm+/HeRV5dod9AUr7yMLHBniI0pF3JNS
wwVJJJgI+vuwQks3+/fJrWEwqtcr37eWlGHQmLCenGqHLEHYBMkY3GgRS2QJOXZN
PDQdTWUkftnnbLEEY2cKQCR8+Z7tjyvdSt8OELqEXLhTLSGlpZsBPLTDhUTtDsRE
eOiyIEvCk18RXIEThvIL/z/IhKwuOMT4zGID7LPnDHzVXiuuo3EZrw9SfCg4R+vz
tlDDvvIvSAX5YzRV9hWF92tpuKc5lPPG7ovaoQEpwlWzE8cmt5XAV28UDfbuaJEq
++K3Roqal0Bnw5FyyNmfYxpUOJXteE/lcbCgPvf0lWZnzu2fRnbaowClQNo7+60H
X6XetOK1Qi1Q5sivdoxH3KBiduX8dEJDpYmPsTm7gZXYRDAINWlNByAjxI/R0q9v
i1+M54RIwXXm0wY2t76YQ45e/AK4Jcl+4UzN1/vMDZ1MJtf7G9g+bnktY/8KYih7
yu7gUVpvh6n1WeSziIApKAO0YMA6dC4evOYEh3tmaTqp+avVnBl5PhEARzu524ZV
8haIDufp8ZROtqDpv6enF79lhEh6vOjxmO/ilIop3X4r9mqx137IURzECgT6dt5T
8Ki9bxWqRmt0xtkFq7UAraUQn8xR+SZ+ZnEr2aDWVnY4BN9mrw5335sSEN0YURAL
qJglL3uI65+ynT2JMmy0psTUJ1xQwMKEx6lxVxvo8e3FsTIVtyVdQMwOpuprxL49
ZdZRg+bAkxROxpo+GqSxrCsBsv8CaSTREx46ZRo6N8kDB5Fm+w4d037ygX8tA4bK
YP8AQyRbLPBX5UIvtA1robyJY4iQBqkUbwIscdlNz/Tume6sf+zfkNJJeqnYnCN7
Pxg0YyqtpYVu5f5IsrOhDqPwi0vT6I32ts0OvwLDPPGYPIvRPQZe4DprT01CmXUY
tbIUEfU1aBZd2GDDgzns7za0PdZwYn7NCgiulUwhXRbSblQLXzMY5ZIufNv78rVq
ozvUCS+an2zHX/ZCPyXHBmKN3u1ozoCgzWS8XoCRehko+7lYtSAg5lh9RE96CmS/
9u7S+uIi30njKowatJOhj2wLDXPH6EipHWPBYs5j7dWR7+xDF6jTpOuL6nfDuOXH
S7JEynu0OBFOUPyoJdKvP4eZ1wLRzypsoX6OzqXwZtt3IJCTIEsU0lhI+om7oB5w
45NQxw81P7BtRUwLOlXcwcbCTj/fzd6iPCSNcNwMH/lOYa2RIjB5Sw7OD6wXvkEq
MpnBewMovHjSsTthpKdlzCkygZs+qu+cp7ru3kTOuRJRvfdG5RuiAv2MEo3IaUL+
CZcDSfqD2vXpO5S6DC8uyNMY69xUI+snPgs0qPEEW4LnjIKOX7lkdh7TZkl7Y5z+
mmrQxv/yxXC1UXB4ZvWHumFCa1f0Bmkmsobwd8czJv2AwfM3Yfk4Mshp7XLOyUGj
rAd8P8LPnyVK14ZOwYlE406JVOX3vUqTxB00bYBhfWeNKD+Ux/uBeOpyGeyxM33B
IlmzsphLE4d0DZHETp0dh5yhGufjqtlGRFlKD1YAiPYUE79WdYQunDjDBeAVV7ej
CfbuBe2yqxJ06EAuLYmEmXgDE3Loi1LZVf5py6J7t6YrpsJh/2EtmHdJ5NukuMb+
acPjX2Er1Cc+Ft30b+7voJzLl9/FGcrqI4pgAmXYCaIviekCwt+7JQdK1l/ATGuk
c0tk+WcZ/TVANIYmq6i7wGhBi0B0YpeYJ1CYrhIottQXfhQTsfIgjc4RpoBKHHx0
UCdAb4uww5oll4kx/ZhmGrP1eOZrFTn/HTzdQ+ErIJbS5DrwdTme0itbIiM7FB04
Gapsoque0otAFJBVB82yK9IKcrUPJzN4fxCuklXDBYtvcMK9Kk/gkPQXOxp1WGNk
/PPediFr95/0U/PQjHEcs4hqfnt2FGTOJSEbo7GvbDH/GnFvYaPUbd00g/nPA5Xd
une6V33aOVNV79o7yhfgeZvkFTaCnrnUnLKOGwHP2ntJclmEeA3UCssV9iNxJYjZ
t0Fr5srvBKvVpzDJUKECibwUnye6dLV9h3AWjXJsPQnaZ94jphIgAoIpXLVoG7L5
hY/r7yg2b1ksu1X5H1u/Xv1XMEdY+tR48nuWNacZ0Tgh5WYrxloIx9ocxrjE01R1
SBWVpC84kyL3hnm7fMqDE0PYlv6nHOW7nTZqZLImK8xs/IorxVvejDF/YJSHg2Kg
GVw/xvRkByCkJNU5gR9UjzK0iOL+Vwcx7uuDGI/B8qj+LMRaPQLJV/uNpM+JauyI
dnhoYDk524E1Zcru+/TFzlASsSE1ZhB2oOo9HitSG891ljUU4ZkgyczMBmzis75V
zvKqgNZAxV4lk1AE2NvEXQenwOVbVL3P3zKnU2xzUpgEiEieEaMAp2GTqEMz5Xts
A0QB+oU8bLYQiksfCQZG2FlV3rIiX8Ukj7UY8xl7ajDXKtOFprCF44BuRnT9Tkye
5MsxRgFOkdJ+pDH73Ssie7zBbAAzcJ/eJbixo7EuDVtqvn7VroCAsI1tQ/7myhK+
ftVsxm3WOHELEMx6BNy+6y2TBEb1o4y8h+T3sF1Pxm3+sfgHmcWugVCSaTiUTyAa
pOwM/7lEyohseRekCdeZLM7pdvg+0vhfgAqdvzJm8z3ogZmwWlNXUG851RWSdpdS
kaYI0nq1Py4VbedId5tlwKe0kVHnDwdrW8Okn4NlaGJi7a81Pz9DwIc4g49GfMsi
/5/xEODi1AUQat5ycM1RuvOSHitTlGRAgY7p+bj6gZX3TJD0zHo3CqF868YdiNxg
Has8VrN/ekYSEydN4VHaUw+OO0IMg44Kt7Kr8Yt0QHKnL53nrI7rBuzhrwkeB8By
JOlqVahEmD8XlsuR1pUx2+4E31VMU9lyPn7gONmRhcEOBlednIXbzvu12/wyHPhm
jMJZL5o88xMM6aTYtjR3i8PVP2thT/mTtdiFk4C/sPFvlraeQXR4nySbIECysvaI
L1vhXjCWtBa1RrVasvEhT0+fVle8JpMMZW/91iW0BV/eBRaNRAvXMLtB3nWVtcF3
ovl86YPEKWzkMbfNSnlIg5zLlr7fviM6slxSzaNtJ2cXHtbRmJNMg+PrqzD+pc08
Z6YRPA+cFlsJ9oeEAvd++GbSQpOefPFrbN3wEIo6CoGUCl1+Q3e1V75UQ7rS6aAn
+PJXBU7BsSWTr57iOl/NVfEcsQurcXDgOXmXDnkf4qq7KbdEg+2PWa/j5iRTwchH
Nqa5f0ao7iDYmq6+MhIx61uWaSEV5QrS17q3wmEn2lyJBseeuGuSZZCrpUTObj2d
7k+mIZCTZceHT9gF1ugLy/ImtQ4uj3bmJCKxJONwRqj520tcAH6XLS2ESRGVEsLW
8tkgM8T3OBGO4XBipK21MiokxpGYB5uQZmp2lBb+A81TkjDWcYzheoNGcWT7QEb3
qMaSsULZoFK0pR1XyyQ/gl7s6Vo5TlVlTCsOWh2HgkwnCGaoAyndDShem8Hi12MJ
EE5fpSKYxwIuvxkpIaRYIyGZUXoVAtBiPbePxc+hF6Iqvuz823L717otEliYPRkw
ppEpwt7pDVFjWXt77U4x0QVargUWVmYU7zb3vJAoVx2VLtntRjTkK0d2moyq2VtH
g7LN3Iqtzh+GqeFItF+47JwYAxxgMkApppbXgpmVJlcNc9PzMFBu4HiOmo9rAFPA
oQHFtdoe324IRxDmBy9NMyuk1afLX8AJHq4qJkQGe9ali4dQr3HBOwwGZtAqnWCE
1r44HqEioWdgV6IinvFFG4cUwGU17kjSm7fjdEILDk3qcdAqwH5QlXzLskiXBHbB
c6ZsYlgAcNxqlwjmy2VP40ukXxHTYg60qxX7W5Q9PsmNBxmXZ+3zzn4ZjvsWTTfb
i+g6snux9yfuPvtKBRuaS9LzbxJn2E3KXIHhUbHOMYjYumREhLcKd7AH0K78+NaN
HIhD3ePdKoJkiiJp0E2huAzmbmRDuEakZ/FtrVneEaOlZPCzuXe7K4e2sWyGJ8qq
aSFEk8mfq0P67FO4FS0l/D+co8Xtto/ajaLUAoVX9LaicSpMq1G6vF3S5uZvLt9q
4o/GDaO8pL/0eQMkE9TUQaachqEec8H87LnY//V6kydU+1w4j+z6eECfc/BSaS7v
D8N/56599pUizZ0o2ChCmAFGDEwjoEudXrj4hXE+N/hziny1nwVimdubPXePw06L
AnclcO0vGDhPZiu5yMLdg6mioKhNuQq10abf/9naZG301XWo4UH67rAfGmXr1x9I
PCVnq0Gg1NHZ2r8WFnMcWxfQdlhkvgfmHn7KNq4GU7kPXU6cd0PECGY1SUbQ4s9E
Ud4QtDpj3SSqbfl8drWbI4e8RDtAOME8a49nw9qXwHXyyrZOT624I2bsBDlW8nI1
snEivXU4zNAB7GJfHEbiFYWxkpvcknH8nQ4pxZMdrEc1TMssy3ZIRpsHsZm/vRPX
Spf8WEN+copxJpQ9brAVBS6Jr0jofICNMqr0Z9wmXmp832n7lrFknQ4WCxuNCZ44
8o/RukjmaBM84wkF+gs6ZkanqEh9h/7RMhSdu+9Zsc0fqjQnURKpuS11Ap10ICLT
mZYx/kEw2fPTJo5JLy7G2J9CZcRzJj3m+3SNYsNLH9bYClhRORRiZ8Bofjt4EcRn
qOSmtY/cEK6dbNsiThluSM7fML3dhFQSax8oWO4KaHPZH1v+NR3/54DQnbL3+YsV
u9bNG03fLB9Zp9sbx+ae6DpYc8dsW05OOOuKzWzjVadHd41DkehSiQdyVawJ9INe
SMMxuwYCvZBMKJBjShtPz2iq2hnT9XrsvfTvR+aMBdM5YW3Qy4lqXIIPdg0GBves
lMMBpkIIi5vGkGdzfNlMZ5L4YUlXikR1DPJrAoFO9dNxlBYLq2JDNxyu8QpL3TpB
vQRCxE92zVw3axSbmIscd3RY5SximuhfGn9G+tiPVEDNaXWkG7+FKmXyt/GmOEQ3
67Uo5bqHYdH7jQJOvlA6eii5O4FJJJAUZnpefMLvXB6ADTIzL69OfFDacTFd4J9E
lzwkrKj2isdN3DTU2DwgNsEbTei3JzuEeg2odXKiiX4friHu4ZPaEPWDJUwbr1gZ
APTTBbcdWJA1JEvBU+YTF/ja3spoIZcncTtdjBxkplYRFiCZAJy13KSVnEn9lmdE
jsyO+psIv8bFVfOqKiD9m/+FFHlqNSNB2tliNyfE7o6hqxEsZH6laDK8HMVJTHHY
DORZTa9tgSeKMXrYT0r0jfv2sQf0bvjAXGs684aUiBPt9gcEueaHGBE9jAq+PPKU
U3HJ9paGXU4rtJB7fxhI1HXejfMJEyzoeAVRJGUpaFB6rVKLbwAdT5tGcFWf2Q7c
2TwxX+4kQAE3b6l/3jXe0Zg14FsfYXM9oe2oPPPYUsPs07hi5M/AT3gPC4Rqk0fL
a4rmyrmj/VdZvS9oQfLLwr6Q5XrWBneR4+11cLZlExltMrPVorWI59lR7TWRrfPO
FfPhsDh5tF1ZwBahQQbnq9h//7qVdCQDi1ScOwRsIP+okaOiLIaA138h0BzTZ7Sj
3sEuFMgqmHhi3fW4GmwFd4Md2A6tzTUtMtQAIDhwhvRVc5IQlUOvITJljJeFV4Vo
v+/h+qFXs4HXIvRoY5YtKkGPPR1T4N1FspAQeU1SuiA7aPYtTd7pGA6pTxImfw3F
yjrJLIoOP099slfaBsjsGy9LpLukoP9wqKXZ0wJH6B35DIWbcINbWyTDwv9Mbx40
hvAc2/FBgyRoKqRmdgfLhZwkNrQuC+mQRsmkeNFbW+klX/D3Zv0PjkAje7Kc2VO6
su6w8hjExcqHGHjqaiVr+nNs5Ycj1H93C6n3Uj8KchiH3pYxPeC/rP6QPE6NVb0k
3sAXineKBmlI3xxUQIPDvHqpBqzGtJoc+fL7tsEUyEMuP/sKUPkDsDyXU9pKmYTH
JHmin8PXoGcWVHao9vArpi9FrR9+LSb2I+Bs5I7cHBrDTOO7g++qNVM73NJTnz57
Lp2amw5Jz8+C00PvTuNiYBkZgek39OJxRLin/Jn9iCf/QO0+8k1qAr6rfgh9llvo
ifqfWE6hLIRnB1JdoLDj0QKitMcYVqSnNmWJ/To18pxOriju/N55E8qAGiR1Dpu/
uVVH2lXIHhgBvho8uLu9aA+emreUmfXsi8wR1St0h229NQH+UIb8c2ihF6J2SKgB
JjSs7X2lTJG+TE00O5+Ev4CLUNQgJL2qRMkwtH/AiPtXSAJK8K9KbyspTv1BRXIk
eQZGSbHJBHMNsHJkNE9/obEd6Oi1EaaXaA4/JAa9MJMIloqLkdPxN6D4NDethv9w
1zW3W2cDfIDdj5eNXl6cjVgC+p0p5oTtQHxI6vAbHaej8KuxYMyvxEsUCaB1mu4U
xQrWeQ1d0bALtVUozdOwR1S+fPXug+gSGFeaxcFHGoV6aG4NxPimMxfyC98A22KW
+dpK38c4onZFXFznUsB9KAMwHichH9t/0aGXWz9eTj4pf3inuhFK2Y+w78ibwpwb
7ggbZenM7RNiXz6pVZxOa7uHMcaaW/YEajuochmvHJyjNU72v1mwfcXQtYJ/Ncjz
BYQPk4TaJFYjR+kIv9epCxt1jKO3HuS2CC5CzzMFTo2/AOdiRPNUuLZYuh4AXUPG
ugb9xuqFM3axiNfq5JhXSyZyuAbSIBDmkXvo4TdWEGGF37GGdHCSkzujnU0ekqEU
5DSm3BMAwIauGq/cJ00Jtz//eP7Mzdb0ul09Y1TXy2oiZYy1iCAGwM2180eQh/KN
xrpKgOeoB9s/u+9NvMTuZaGe6JBzHrz6KliQpWuuPOm8wbdY2NHzC2iyn/ZmJRFx
wCc0ctP9r2X4CVUgQDnO4fw35HVsBZpBi0DHsNDTZ74jluvnSSTFF9i6B53m54vR
1bsQd0Pq+I7rN1w0LtfW2spZ9H9Dw/TDC0X0LdvD7qLm8P0mt7YTUphix4BOqPuq
AFZYULNPU/R6owas8TCtUJ74eKDz/rTIfiQAdjIWXtwXD/MJ0LV6ZcLNqmXXxRQN
0eY3bxqHXCm9Dojhmzkk2CIXIi6VmTo9RYJesCQg3KcB7ujoOae4FJHqF3+QEOa1
kBc6E26S9cX+zwU1onL6iFyonZM1Ec2Fy+XCy7hmSf2ywnxZV25Occ/hw+YLbToR
u7yBU+s19mNrCCXIfNE/R0b/MaA4xgunGjZhTINI2+2E7rTVg6HLe1eoC2cII3LU
NdfnjOxFNGED1mAe2LTPnnxzh1nDoY0T5R6jDPnczCtRSLlv9SiAN4vspn8PEQFk
w6zKLwB9EWT9wYb91LBZ9es09zHkrOGAlQNkwBFFTIexTyLhRUva1cO8Pkb8evoU
QbUvR/TueE6L5haf9lRc6GC2kTSZXDt6AiFzv+QK4pDiHp8111W635U8aE9gQJs1
SPNGKmxq9g1Mpw87pihZaSuYHL7bVBo1hWljqLPErMpCCT32kC+WjWsMlugUVTXG
Dlf20zFkW7PD7eaW/9GXVFdi0fn5oxGuiz4noCNEHa3NVae+CqwXtfaTVWpvUFJG
0/pw/ik9qC0uJlfJUbdfKU/3nWIfX3JPdrLioCZerzXaTJdc1eyw9xpaScTZsEdj
tVBKWw1oEqqNYQRcaXpZSyh11Fclz7Bk3ZhVpoWv5SZ9YUHEp3d02s+X1ovduaTG
Rph3UXal8aAZApbLC78vMcJEltVIcUGC+OGuo3XckIj5vE2rGIhOKqxeikWLNerI
Vx0zdcCMrb/14J+vwn22FzTKokOs4ZEZaCQhvgZMcJLGYPQ0A1UgX9K5bCKtGjho
EYyj740mHMcqHzSZIyG2fTo94dRNFdYcKpSVyznhbQrsddw53b5ruBUciG6PjcBh
V0Qj6cavNPTl3sHzGvT/X/uKeP5XLomPzE5MPob6rvORmFB0mb+DccWlfv6rZWo1
wHSYisWUh9SPGdf/UsjYY/zK1MefXf2Mc8X/1UaEAslsU3ctY8EAzHHacK/Kzbjt
hohlIOFYWcmxQWfb+yK2clniVSXVapA7PWXma5c0a47ratL4myKLoC+/Xa7wg5DM
5YOmwHNxUi1XH5A2tJq46f/pIJKXrpmiMgDzThuJpl+/r/ckcaq4E2BBFDv+b8Lk
aMP/SRj6TA4P1SUnm4gZFXAVzibURzsnQ/yvydNiy+ofUSENsXRN7jJPht0kyh8s
UgS+RoAAdbl3/ByUw/Cio6ZqrlxAqt+ZwSbAskUrjv2N6jIdHXHkVBVKnAczAHHS
fwO357g7/I75XgQXEkWr9CGj9toUBC3LJ/rs0Kj3rPVGLysHzfDGV9kTlg0DfmOO
MNkD5tXHenTQ/VoJU/1f8lOhx4+6kNe/qkklgVVPyTcTBBFWu7BpRP+wdUiA/wu8
hrR/6taiE5HEJgkZ4H0N1hFvWcHhlFMZvC4sRXiFYCy+ngyv3mUgA926+fx5/cOX
MGNu7s39HObobliANvd5rW8fe8rpNQK84BDgoKCZDqvY3iopX642KIXM78x48g5V
w4bo4LwnxheGfCMCbMF9oUy6ma4PxJUf1cSse2s3ixFDV5Ea7dfu54Dj/l/0pkFp
wdjTgfNtKH4oCNiGSKQy0AtgJA6TMApAIo3uDfZj5yHq89gVqBMM7d3+vZIQoxYX
Xs1JbbXIrDPHY7RegjPqGWYoTvrMVYZNDzw6kykEa0wlpy7ryJ3FfDz5tTTKVCNP
jevRDywt6nUsL+IWFpfIZ/9vjJ1AhnSdFVz9LIwTFGkKreU8VCA+nQ9PPBb1xe14
8XLOJJqTauaqWd69/4icfCu6zFlYzAcHbJg/8+MspajaPjxxPmvCQHqtZ3U934lJ
yyBIEFoqgr4K1HoXcchH9glv3aYp/M0dI0Jo5RK2J1SWCpYQrDVcE/PtKvthk7LH
lIon9vtKHr3/R/p580j/KaFbBvlz8fPsJYLkidovyfoinVjiRArdFoVmhJ4hK7cX
Oxnr+v/H/Z4mIXUwWqFitLQo2N+ohM7Q4HlMDY5L45IvXoBVEFECoWLE5sfJogyT
ZhzPU+Y4kZnZbAMK2Ej8wJmO9FmhV0b5KxnSPQWugVy7Aw396ZV5OBztEN5OFK94
HySKaLqS4RTRlULUXJGTO+gbK4yjJTo+cPLKEsIS62u6LO5hfJPi8eI3SfBe2tgs
AAW80RwjsvAxyeuCPjfZ2jgt084/FI7xUmCVX6eB1lEOxXvxOMftU/tEer+QobXn
F5KWz0Vpi1DYM8Kmrwcc/qzZuqPN+uM8qJ0FbjKta4ujJpBgtCAdbsNw/2vjT6Yb
oDUqYGj09Z5IWVbOI+QRgzB8dBDLxGuZlVY47P5JMu81eYF0FNccoHL78eLOFpYq
Zn9CS8qB7wtxNqGAsoNbLadiw5GjbPLCckbdAZiSp+1BkdxcxAdV21U6Nr2xqN1J
B15NOYtWKvxIyJYiOdlIgCUlMIc7v75iiRAJXvnFAyCnF87IRtijTnxbpJuDfzZt
en/Db4tk/ehF3z5I0iNAdcwuBUF6yaHAFbdL6sZvM6qqlqUU4l24Lz5WEPm+s43n
6CknG9uTGzkXvhEPRFmX84L/SKeD/OW2MUmi+Ji+TiYn4c4AfOsL9trWZz0P01iD
E2X7QBIKSUyiFDYLLmeyN4nr7KiWiO/7lP/4OQ4Fwddd+SatiQQrOr2ew/vf+fdp
xhk+c5ZkQdIHagH3jDG+yNRj9qGkEcCUB3LVbsUp3Xf0gJ0Qf63nZPHnwOiL9+PE
2F45afXCVacZG4BJj3GhXsyYP3o8+rfT2vYuwWow1uTjk1n1bY+AAk0J7iImC3hV
rq6aPYqzYY35RktgrBjD9YPAYCwGlb6aH8IFX5a2MooYZjaTMaBkqIgTtOKGVoVN
oLzs9u0N73pDzKfCQJuIcdlkw/3GEfayJ+mYHTaVY7ZUM8yPNNM3e7daLEMFCg4n
cJYYNgGlGGbJTl5R4YcOm2UmYGygVQratWgKb2s194fip9fR82KmDlXBRJHenyou
Kn1jsBPuDYDnciKdAVz4GIMwGTHlv5WJG7qoICpdTXRtDHZfxfHk9kRMUWeT+Mkm
A1tq+rHbrmsjh2FzrOHLNNan7Bh/6QZIu+RU1IDziQagiYXW6t2L/lmSHfz0Dbnm
CgtdFqRx07BI0VEekkaaxygZfPKD/tBNVBLuTnhgIC5ww9Hg3brL/bA9A0hxkbkW
EqGXFCCwzPFtJGPZFBWTV6tDLKZTLBuVxMDi/YwGZIA906mIjBgPbfJiWxECAe6z
T0GZL7vJIhX+lZ0FamUwwBoLIlZzzSN0WJNR9150cdGWOgQkX3n6LvajZP5oz0e0
72ta6o2uxoXpJT7tlcyvVVRST5r4r7MFh55AI49hDl1P/ST2E4PVltw9sNthq5/q
dj1JpNc1S0xmOTm3XW5gwgZegNUqfy+P/1eyGSLboqQ2LV1arU77wl77taAg+rCa
HPs0/XJ9E9u2Ak8pnPH9HGTnqlWCfwNsf33Wz/aEH57rKraVwTCZUgeBM9MWGkBr
iw6GZilG1IcEkfSz3Yl2b+tOdmj3QvUPqBfBmWIvOfse0AkTMi3pDXi3WXw5kyU5
Fm7fMwg8gvAXR1QAOPcN1X3Ov5vLd38ELg2JnDUukorNlm0zS4HzR0SYvK0pcIpm
Jax55Hg0ZkregsaPAic64fGsWyOVa8uTBitGL0G1iZ8qgJuwZrLbxdgU3kpYAooX
KElDaBgzARxuhDuXM8tS4P6CNdYZtMh8rTqEpNrgaEK9Az3n/QbMVHoQfbV/ZHa9
kU9qeVw50QyoVxwFGonedME/Y4fE/bQUJpDDgt7nd6dIgi16+jMWvK4ZBCA64MMG
alk3Ue9NDPWgfQG3iLcxGIgydGGkE/Zfqnptyu/GixDj9/W3/RNgtkjcrNkIz7qF
wIR8VruZMBIhARkk3QH5Lwc2VSvpW21H3+1+iP2+qD6bD+q1Z1/JhrxSerMtii2a
JyDiFN1T2jCNpcciGYm4otm6ikOxd6Sym6HGjRQcWNLa+nbuwRJo83F+EIb71B18
8AOfo0dcnt94gPrjvpFv14BDqMAjo2bR58msMMS1tYXUj0S3kZX5x2ANr7f7losb
rGZsxzo2k4mw7iGkrlnm9pR5BMQ4ku5A4Z2u6jb8tnOUEFyKl7kFz131UignRJS1
fYxMr0M29VJhlJKrj8MROvaHKO7mJLdnsSjkV1NwtmOnejFKvcYtIkFrKx2JtqDO
XAr3kYLOfRZlIyP5muk4Uu6cK0toj/mP8yDglwhziox0lCWMvZr5/w+2UI5oU15E
xQeeC4/j/bFDSUPfclTpSBx7KUloFp9kkFbKsyCw/eFaZ+7d9KRl+7/rz8hJdeUs
qd/FAyimEx3ePcmMVS+LpSdvLQwx2Y0Jf5xKYZruHO5W8mr+WKNj/mYHxxIC2+Ro
Opr9TlG1RYGQX1P7OLs7PxuoNN0IHq7s597SdhMWQ+fRj2h/5zkYQWjRWw7QvtL+
LQ8Z4+gti/Ue6b256EZDwqrFVxo43vI26rZlnonBA7foEksoGpAmkXV2RTotq6qA
tN1VzMdoNzSdSnL9tUi146eL+hTGXHFlvDj36wltUoYoQ4MpSL7Re8IGO/esggzz
eZFjJDspxGm4MiaiUuOnE2VWyOGFPwztE5hiSUJwlevSXF1cSJ8jM+4aLgUPFanm
bWnNXGeXZqrkTPa1fWzjFTn2zaBDP4iVZInUc2YlgnWt2zycSW/28RD77czQKlGq
UhrbF107jVN9Q0alBHeLlwV3+hLFHzkiYPuigPloxnBRsIJ3MP8wfIuM9yuxutVe
Crxno4aLDaTkvsh4ZWq/oytbos8LEXzCbH+MV3KvFYADmKuAvue2JTkdRvVlhagY
Xace3+2jQD+Le/EuzVyLY1ZlvbEENp5RbXI1UqH3vsr+GBDmlKjMg+jDboK6DUCP
kyYIUZ3CYbWnWqf3TXTeerBKJlZfWFg+jdR1RPUb9XyNbQMZbhmhw76CazA41d58
X1tIF1cQMoyD7ptR75D7CpxLlsA7WiTMuH4TIYohyViD1izvpzBboNYiebnapUTf
9hIzsy9CiypEPpHpW6fgQVU1/LyLih5bU2cfJdXGNrdnJiN7EvRqKnX7Tdb6bL3T
jBAZV+Ik1mc2YzV6WsAONu3rzrxvHpoNCw/Qs4BKwVBaVd9tGBf75cw88446j4/a
yfZKtdvNML4EYe6pvK1B64jIrXQlkD9Y1FRl2/RMueci37DQ5kji0vTLbg2k2Gco
S+Xz1S1rfxuplZoNU7Hog/unIu4kI9gtqaj2HBliiKXAe7c5zUA5aL/UJU2vSkDm
mD/DUCsmvsIkJet9Ry2JfjbYZOfntHx/aUyIuqh1xrIp234gGVBqC9Yovmgo3dxU
1rl9o7MRKlYLdfHtft1nxqFE50thwhh9QHjI+AbqWBXls9CFpB6tykc8dExl6shC
NUktuJ5wNfOO2hJ83xgOtrCGQs6+m2wCxVKEA2hl1SVqwj9MW3oBC71KhDRragOF
9RLMk8GkQEgqJOEOPP2KIR/cGGAX0D11F0guOQWj8Tz8wXGgFxAAb8WPhA0PpAto
BQyokxo9TGtwtDPy41blxryJ1wkN3heW/bskRFylbJkZgrGlgiJWJWn0M+GnlvB9
E369OMVczmkerXF1ugfTdQFgBi6q2mOAuRQVqWqffn5aEaAhEDZhJauRztm1MaNw
1k4UZBUsUgAFWB9rMB5lqlN2i4xhCgrfVVA9t3S841lu4I/6oDI1bgHStG8mmFBU
HctD8KBgc0SpTlcKmcenRLYLI4LhwD3fs0EFJvkt1LooPlTxH99x5q9O8iCf4rPk
SBHbEBk/586DWZc3e193OtehbXJmTl62TY1ojbHXR4PpRBB3oddMnZkni8EjIhqu
HZtKhvFAskp+6rDd+vvGxoiEb6fid+cHj8xJUWFieuK5XejwFPVVlQO82P6Lug1N
vbI175AUIxm70guUIL1kIJGtQeymaVjt4pG5X5kVNsgpSjy1SPx9WG1uSlQ5dAHB
9ZFogWgV6ySMPKBS6Bwgd99u/39iumObgrnm//yY3/MV/G3OJVn+1jouPxqPt7Fq
2HG0otuKftqxDf9EPJ87OcxjJqtrGBvejdo1GZp5U9bMrXzPxpLmuDUzfJ7xnhz5
Utdb0I+OhZAwlUuLGMoClyvad1jQvBh3/Py/2K7dOXAP16bzIUFlq029jgcvXyPi
6eM2RYeixMCeT4mh8jAF7H5lGDTQ+5qW+fZCts9ptZvlk4AwymIOxu+WNZc0bDxN
DjldO6nfruH5bV4s5GiHfgeAFWTJPmw50QuJWts3W6JKSCYz0dT2+YiSy8PPdJig
s2ns936Z+76Cd+2ZYcUXAl8yIHQb4fa/ulEzkGGYauOw/b5+56neU7DezNDC5aXr
pKBswj1P/vESGniXbnlD5JYICxgXRSmPfNV7uW8eba8yuewgRnOqNDg8OdYFAKdE
tdSjS2XWrTbMbU9opqy+365LYKV7WageeLr63WiyDyElGCkUwCuQYNrwTczumw1y
37thNelsdiZBDRT7GaIlgmrr1lguBR4b0wtdnKV97oAFPN1HKHFBrndy7MOU985D
FN2Qpp1rUphXE38ody3eMl6ts1B0gSutM+ThFoWHby2QOhHfCWTTNAYpsu+1AJzp
eFTp6FCNK3j6OFEsIAcvAku/hkpnRMz+157acFwhJolEO8+JNKOSIifW/McSxmLx
W1hiW2Me88Wn0sy2oduU60VOaRKTVPXYAbuEP8x1axqkxG2MgsOhznsGi2LYWfO6
y7CjozTY8UMLn7Z9yzqX1tHBlfNl3pMbCdiUUZspBb9qAvd0IFiJ77eKWo7xY1Y7
Maz11WAtJl3Oz9SeB13QpJ/iwOCe3FnbW+NcDjvS44MagiUWKBxEJgsg5E26iirI
AFhmmw5NkZo9HhSdFdS/8DBySL7zUifod0uKEkjFzb/ILLNsBkexuvuO8N8TEjk3
AFWC7BSjXk6adGG9Opo/7NpKgmqlnqd8T6PrgpnohLdeeb3/F6a/i3XGEDGBjnRb
d2lCIOHIjGwISWuwEBd79cuUFXAMeE11k3+A4dOU3XceoF/q1opfnNHVqVnIgDa2
lbhWa/uUH95mFfHsxQ5ytYm7DpoKIyhysieGurkcoSZKjebrFCuzqdFO2blJDH0b
K1oQthxZ6ylQPMWcRS4cNlu5qe1lT3EVwfKCGjXB3wwSyKmgz5SJTJq8eG6jIddm
aqvegYwp2E2ATuNJ3abKVoX2kqGjGM6EEYARxyfkCSTYNxT0gZs8zwiYg5QMWOwI
VO3lPVQV0KB4qjJL3f+XXnKXjAOUVCL0qmu6uWWtWS4+vP6lBbgQ8/89DjnMMqUL
s9QG10s/SUfzeA9+eVJX6HU4Z1hrJUCaB37onARyXa23aLrHmgvfBjD+zVTblBJv
n4v3gRuYLXXy6uSzf2n2Prdv9LLUmULrAODql6bu5FsB8y1c6MdfD5IlKJ2YlfXp
YxjkLd2exF3fjONEWDG4huhNqZe5EYKi7s1xR1lZrcB3Kyve7srv35hlAoSvkHk4
FcHGr8sVjAv58wZCi1V7DruIXKJglttA0iV5ZZjcmgrguNpRaZkD7J3N5xr48O/o
EVHjjFQGkHNHRA5xJISICu0uL3DOncOoGB3rqe3yyt6Lr57KylqVAWvRgeeGzqae
oTTGytgKGUMezBm8a8jIbvFEmFXNE5kmKqb0Fy2sazMFM13BMsTs8KfTfloYtpAi
Rj5XPoZe/KdUS3Huf+u6uw5f5DzIHdggg1qmGL79Y7UH0e9NEfYXwzXisrELZ6mh
zd/VAC5SVuO0DpQPiSEkVZR3hKG+tgZQpyUf415cthWAlBH/XkO+YsrfGvrZMH+0
f3mHwZrWMV7D9/4Aq7KxfbGbjxkzTWUdWfAaKsuNe0Sehu3vpmYuRbAq8bpn23tL
rjPjluYt0lWBtUiwLr/JhPyaUTYfVcPRz1zDJXfAXFINQ1My/5FToDyz+O8Ga5Ca
/FSyzJt5GHYW+RDmnF/QCByBfU7s8dmJurMHepwuxRQdkwgDeAjPZRKLyG1pEBg/
77kimfgJO2V54lZ/pT5pOwW1ohIKesDYVPI3yzTIJ6aQjO3rkRsaYhV1JlJTPz6w
4pFrfJIZUQ7iBRiritz1dPnpQV0ED/ua1UCOizLJOP3X1FsPoRdKb263+PgTp5l5
wo1O9/lF7HW5+LZbReOACJGtmNq0wMRAEwfMd6ahRyvfo+c0uO910oyuicihQb4q
Rx9Osd/EDzvIjRPhTY/0Bar5Av9S6TgnF2nmBRaIvpi6KIvMiQE48/s4CuGPNy+Q
BFI2ePSIxoGxtUxO2Vvxw/a5UUMDBvnim3vYfHkOquWvKRs8rL0HJDVqkReKukVh
8GhXGDLDJSDkjhDS9uDx3kIN8KoMYwP+DbcabbsoNcEyzaDO+ZW5bb8jM4MbXEkt
u9jIxjR7wRJ6rA/AsYbAXCVTau381R7gDJxrKGnVaExNWY+wDfTqgd4dxuvWaGzI
65D5eKpFrnjQKLhxZUMzQpMS/WMeq2EMMDfW39uopNYNr+t2wsCyfdoSpz1gwvHo
BurLEWinXRtoWSpcgj/iPKXu28GTPeTb+klNJyVoBxYRoOaJrIRfmZuViIgDb/lH
qOWJ0LfaUjlpV5gDNrYS9xhftC1uwGWJDBcxJuAdtaQHS7VAGWD3ctWDsV+WtnEU
YsQrXZ/TOUxRFmHTGqzmXplapWhseFLfyBEqu3OMyyEz4emdaGNSpqqn/JRPJTEQ
79s9zsUMIgaQvuPTawCS6YmCE0YVlqwRICeYZ7o2+yKlOnL67MvgQ2QVZpn04QRm
lDoHJLnhB/dX50ZudHQMNW8yUlDa3v/lEvqZZVPZPPRLXOjHbfWoi3fX5SFeBrTT
L+LjAUzbvZCp0016oJiXyCBP1grU6qKjf5Aol6baFDGIYwVH0eFRa/fM5zVj9FKS
`protect end_protected
