-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
0UADS54FswngcWUu6anUD5IrVCiiJIQFfWEZnKmIYKRiS6P5TkP/zyzQPZ/npJuB
aXyJogYTIqQGu4rjLnaxpCu959AF0p5RwNMIGsTG1PqlkmhTEw5ZPP8oHfF9Ra8O
4kvxIWwUOWEmubjWhNovrZ6Ydibq2lkY3wJYGt93Jao=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 98352)
`protect data_block
6yBOr6sFrhXMsRw0r6maZNMNlYytZ4l05aJ57ME0r4olFuI2Qot3FD/930ZQYCbG
D15vQxZ8se2hzHyKcB82DCfnHsRUepcHq6QjTiszShtmyPLkm/BM+x6kJtUs2jyL
VU+cLc8Tb9tjLLqDJLP7aJYMVepSBWkje1bTVQV7PGl3rNWM6oeDgjrlB5uNP7M5
45GGVqwNBqOGP/Xif5luHx1jN+K884tygEyNFWbH8LB0E+eBODBHCsN2kDUD8vgg
sCH4KhdFnRhuFE2ohNoxF6g9BIBtEjsw41QkG0H6Jc+y2vBjuslqJjBi9gP/b80X
n8kUiVwOCo0d6jbMHyu7YNAFJAh02lzuo8GrKazN4a2v6DBBL3QEP4M39tnju05l
KzVGoKXZls/CR/nNqnacF/ey987Z7vZ4CUumLBE/eMj7toLMKNAZmyNodyo20sK7
yfPIzJKp4hNvjYkjmfesrV6HWrdo6kUXxNMdot0noy+S2qGgx7DN61Rn2A8u7nE1
xvF9Fciis7CvWc7dFn+nAv3O5efk2pg5Z6f82JLCSpJP8bHP8ZGI2OomW0Tak43F
BxU8L8UZwz9O7wxVVjBIAnnPdijU1Ssb49AjJTjOrW8Pye0rw+cfNeiqjpq11/F9
I4Zy1PAGvE31rlGhANkoQp4X4o9PbJe0cGF0bddRoncT9LcCjIm1+fSJm9gD9AqH
ktYbOZSiYmS9NsCg6/BFZ/H7KdSoIPgbt61ig2y7RXuHq4qoTEnCcf0qxQakCil+
E/TSEV6MB6ibF22FT4N/U5sOoBCgZkW5JvzE8yauzV/JNboDVE2NLKJd6exHvV/J
g1qV1O/8T7VA2yqIb6/MCUZDCrrdMsoV9zfWZI68nwGAggx4AAcN7ZdEkJt53tNa
xh4IU74mqCd3SoARisKJXlCnlAuzu/7zbQfsVD8z0S4zt+MVfoxWz4M1Sy75Jtsg
RuHgb+mPox0HTZo5AdNsP0Mq7ckz8gw7r6achQAVCekvETUpOTYMzgo6EB5naGMm
Atyixff5YErC61S8QA52GD98KIeM7M7rKHGeFDPToB2kzgCs1QKqBeiIDIUjQ03C
1JFLU88TcfcaYohXRc5qk1Wl/fi+yW/ijR0k8Vztcd5esvHGf784tUglo2jSpM1T
q/UYXYiW6AfPQu5srvDtMqmMJz2S9dugVJ8HYbTq9jmCRu6kmpH6RS9OCG8YON8z
fyQeNwrrelExOOTKj7vXF+N0bIkV/r6q2Bk+B1+/Or6Q78wLgaepgRJuRB7P8CYY
NFwry82i16kFt4yvS445znXIprsjSwg2U2PgI00kz/bjkwJ2IRfQAZk2pyolbJpe
3fMJqVlsBukuzK4tGHZoudA4yqM02qoI6duaXCq86CK4DZpSRSVMjo/j632PBs2b
NY0Iz5YEcgHnQDZcq/v/4u9pc9RZTjrDQgcLZtEepTSG0TduG58p0eidhod/XKwP
0i6wo4lbH52Q1dxcQ1LjAKtNSpyayLerGWGkb+Qpw6KmVt6kdShCgrXBajB3L0pX
H7jwpaGYfzjz4W/BhzEjQypdc8W/2A7lFltgLOM1h62OsuvbU1uti1UNT/zIO1UT
xw/cxeTKLCzZxoSUtczDCTtFreJXGk88fxolLv6698KprzCszcI5ZGQ7kZVwuXsE
uZm+nwYoFYhkCofjVC77Ru/eWIKekjqeeynSEyBiZxittb2EUSp0A6yeRrCf/3Yo
yHBY6iyTcjKB/NZl1M9dWUfbZ1BM8BWXK0XahQ7cCX0ctYlXjS1MwU81PtSTrhBs
WmgGxOtHZl1NALMqnrOObPKZfG39n+fC9RqaPDpRYzGRFlbhCAPKuDPKoQu34ikP
4uZenIsNeCkwJLg0jH+VBKqNZqdG9L3V0KwpdgIB62/T8VUSY+r8nAU2yTxJCZnL
jpX8rvf7kvzSxcyRJC6jXO39hN9MfiFMUCLLmw3srIzKYCXJqQwC+zxfW1ebAIeS
R4NUCOFLG3QMdG5zOt37D1GBD8twxUzOeqS/1hlQe1rO8tOFJHj8t66/x9dHLRuG
aMeHh7xva6vTegM3LNfZQY4ZP4XsIlSdqfeWLHV8MkqFya6MRZGNVGlycTV24wwp
79wAF8tzJ+sAirxb2dej3uMlAYSw/dCuMxuV6exPI+9ZNd1qR/OrJZbeRnjRzs5f
NqT6fM7O0L0lWx+3mrfxAt9mEuLUwmOUnI0bPmPrllh+Gc7Vu/vbYnWaVPQK+6/1
x7q8tvoFgK8HqoPV1/Kvk+TXR0NbSjfT7REUqKhI5/lI5ZINVFN3bT1imZUeRG0/
8v3PxnInzkBKnyLqhTu6NhdUFjfDIHerarLNe59AB8jyAhiRngUeVUevRwSIgTj8
fF84wcFdGc0zvZdjZrxpdCy3Vv7AsvagcqOnptrdAVRduBEyO0mzyYIYeHUViutf
kzKELKwIYbno3Qo6B2kace4HNJ4oH7Q95oxzUAUS59+d2WIBoEKOBcM+WHpQxneZ
E2gqPyk5n9WZxLnEan9Utk2BLh3dz5afMKtuVyxKZzSm0fhcPQk44TfInVLv1uyV
/I9IJtxeFm6MDDTccaE7F1fagvKCk436ahsLtshO0NWIQgq/Q2V2qhDsRPVSUvXW
8EwL235ib5RCNJ1ipANBG9214OxfhFkJ+oojfwO2dRjDr7o5aSaZPgTxBsFRO1Uk
N+s9nlmaLs+f3tawJq4wMnrMpmW/qj8dNDx/TvJTIbMyCGYJuC4vw6KslibtG0xW
0knzN8cBaD3Y0j/zntLpIQvkoUMr/E5JjdwGxE31vnHfTeWRPUFPwKxkXvCk2gc1
5FblcnFXOf87Ol4AMD5bWyt3g5ivbLdNSzGqVyYU63wnhMj+xpjhMkYAeQiqdlOc
lGckzE1EThx4iDCrNXqkDnNvYrxhwxTspVHWm6yKdxC3NsUjaRFE84lHd1hi5YMh
5R3Q5VEG/Je2sSKijH1PWtVgmua6k16yXHz5orcSOTeJ7b07TF2QWZVPZejAG+AS
DcZTSQClVePQVuRw9ZC/vp+9lSIYLDd5/gL/9sog2LIiMtFg9qa/5umiS890Hg+N
ujfQcVReZYRbPwfixZlkHiBnip5Xtk8YdHJt5spza0x9BnwQs+c3CoxoxI9iagbx
Xoev6hQtNFLs21rqUbo5Z8ChEMS5Hc/aca2WqMGqzlcoNiBbtoppSgbu9tZZ3Mfd
YadDOzoATAS6WNgjAPLNkMg+BjGp0Xh3cH+oHOLv7MxpiOo+Mtq02mMz9lI6F4i+
hcn3tYvscahnDZ0M6edVHZlSCMww9oa3p2ZYbhQ2l5IWqnvbzKHz8DnPHe0h+xtj
jLg4astROkOt5HkJEfju5WO7Q/qB0I3P20eAV/Fi1+TYi4Qz0vN43FRBxFv2yxmr
vMdxXtOkV/RSESqVUrZwvylvT5NZNvhdTMHMt4e6RHlvtJBACWVw41m8BLSaz38D
lqXzFSgGCJI2OSHKLP8ieA5nqSRJM4MG3N8DWgYdZFxxLJdbODJwRghzs+BsRRtA
xvvZSDUorzcdZ4Q1aJfTbnW9BUiUxCgnWl+NQlMVsnNOblEXEJRXFub6XujOaV1O
pexN50gNluACpyqE4f8Uof2I008aQ/iiCcqREAf/Idkbat42yqY/sinWjy4Oh96W
gJXGINS1aaI/m8QiGV3PgFKUqz+wtQuefBou8a+aKpjN1Iddu0MgxBPi/z9wIzng
AUWJiGLEJp1VusH+ImSZC3vHl49s+iNsgO5ttpzcaaY1My+pIpJ4ChwP0k+TMGD3
cm5HuQM4vcGRHvJfhu5G9NEh01h5jTjrq+OCdObRKp2MI/FS72FFQi2H5hO4m+1F
DiAH66tQ5qejuqB3ed+XHHCxbJOqiNa4zCrn1adgkbNHBTc9JbXaMOByL36G2vY5
nxPcc3Dwiq10ign8KBjWQgd3IF35Rw1Z1hHg9dJKcWebJMaTc0+czJ6BLhLBJgKg
ywRqk3fKgXM6ubh8MDLM6n7bCtXpO88RV1HDUFRfWb+x62e8lcjnjHMf5vnjYOwh
aDIq9DsAcWixw/jVv2AZ53Gna+18d+U4Dxe/DkUo5e4YDHar8rWWk/GsifgFi/Bb
51avIj36l1gNb3y8JPnh3vzDK9KEgMeqlc9gPCZMuI474oSCICaP917T68kWGxTZ
RuXdNPDOPlBqCTUbW3ZekP/ALMX6dpX86d+QHUFl16G++QpgCzra4rzEy0bC+Mcr
RDLUjVk0RcU+BPz0DfeDmvx+Qcu6i74nl6cctEJcMhyBlhFHlJcQ5ANz9zxKMC17
fbEQNsyuYebi1XNo4k+VWoyGNz14vjP+Z/PXdmYKV4l/CgDWSBEToOb7pu1+LZW5
qDIdMQheFExKOA6rGvSaeFCqeH/860TndnK9EkxK4Re1ltKSJwWVsnFyUjXMh7jO
it1ye2GoVvUEJEtuIwWXba1ZVECSvKUyZY/gdNXd1SY6ZFJ0iCmsfe9xgdp/89SX
dVwlZxCrFipphgmh9oR66bxJ0nwRsJuHRCKkPQvblKQGECDXDDgHfhfl65KdAozl
ed8qBrB6IQbWIBhnjPHuPnP2woU8CPvV32d39YNhGKgglfs/FGER8Rm6yxHwAxFm
LyHbimW+f/P/GKEz8shPNUEFKUtlWuUNQvTer3PKVDwu33Vk2I5urSwdk37l01IR
LItFhdPkmczIGMJcyntZOGkm++T3yfQEBQAATruOZsHM2wOHxZpj/CGh6QYawNxd
6Iz2hPRa3NnZ13DPUGLgQGH1uXm8SIIRrE5mBIsbi3Vx4ZpEagpLQ7Dh8bUrc3bc
7un91kU4AsokIJMGbNf6te/LlFvv1v+YFM2JEDkvxzX9h95iQ2sh1SinLYCcjzNo
jfCvRaoEuqlfRjnNK08OSDU1aan6h7PyQ5tQDOYLpbNEEgvwVBoTnG4pTbAi0MMS
YkARaDDPlSKdsGDGGMn+4PIK2Wby1c3fa/EI2zYZwUsLvjUeGdb+wCQTczuWV2hz
Ee8tw4N9yQBOndZVgYfPfqrNCyXGy9N4r/AaPME506vt9JtPVKYVKKszg88xEAe/
L+JBFWshzCcGePI8bDqgkNy+0oGW0b6qrYcRLIQzrE7yq3aNHUa3bqdK0A/XXW/m
zeLZMYFOMZHv27KwGbPAJwzzSmxMpg9rc+BQ+dfA6kbRtO/oNjJdkIdYTB4u23AS
xV7Zb0jpvGX/Z96hN9Dt8qVgCqPA/JzYcRNhheR98+oHUlGgZpHsrg40C5QOLC/i
hHbHjAJjySUjh3XBo38/60mokAxIh/Yg5Ma0u6RkiQmTQLKxfiWoECE663Euk3s2
6Fyby6iWauDGUBC/tvOklGMw/MF4Xf1P6EHRhcWj6h1RQ/gdU+gg6/eNR5ujHm/1
NLg1qqBqwKqLnnOkNeEgW5X6LZR3YwL/B8glGUIkJFKQnwz7C7dAlDsUTgsfXyZ5
n/k+8ugd5yL9L0ICKiqkWvmPyRdB5qDsmkXya1fSlARd9g7VgtDOrovltKlFoiFu
+QQILhbJYH1fZ7Q16w2PUU5qZaSA/5/7wZFfg3sSSZBtWuH9roYsFKwTPG5EnKuD
RDFZVkoebTdedfKk9qKvsbIv33a9XeYPMyivXhLOga5v5Pd6R/v3tXJPZVn8UGh0
qwnO6NTIUytdP6j+DB/krEjmBJkSiTqP06J2lzqaHOTET5n0Mz8reNneK6UbBuxI
0Sbv6lpEZqWB5HgLE429xk1XDaUwKsIkutwyyIz1aYPxc6xvFAPzfBYlqvE7Rvbc
v5YwgjgMOEkV60yyQZ9dZUYxtOT4oJwPk4SikI/8GpgFJSg6rFPfiHsJ8O9F8DZy
WcJBI3dKJ6Td/jmnadXtrCYgaI9cEwYqX9cIuVgeAXXQkmqs1wZdVJxN5n6hzJNH
VLBTo02qEJkteqWBCBm1GCzB1uFUYOI0l1l7BcYyBKAVB4kNgXnWPegJ5shcReyd
p/P6Lp7plnKEupUV38SeAkKRob9FrXajazyeQox9lKssQTOHd6zrc8yzGrb3Ee50
pLqlUlAsyg0On8ZuUPQeZO+h4GUXUj4hFR3H5Nq6zxqerS46D6WpTEMdAXuNO2ls
eeDSZu9GgDc5jmR/F5ftQw68ZNxektZ35B/UoKC1yWJq0Bs4SFCFD3vOVTXUO2c0
ayHfzeyZe+88sJmJjxphCMV35iV8NHadeuCpFEWQCj92QydxGvXF00pEYJcS77cF
erKB4XwJMqBN6vMW80i64TURSVW3cxi2jevQoWL8wgcyQULh0bkBsXaaYxLJTB+0
4bytEllWaeREBgWM9oAUChHEHXkzeIIeCsDoo3ePbUZu7sMBuZNTR0cW3hzNmZpT
S458Su+q/sv7zCddWfhH1qPts0LsmALX9p3XdC/rMoVgz7xAxTG3auQMCEX1owcu
nKy1Oaiyw2oayTxtfqCT0u/oHWhugiLt1o1GEKgtvY0UZn9E+X7MHotPrNoKXkuo
I/cPMngkzgHcWo0G26x+OC11Cdl8CS/NLRr9CgAHa8DnMaFJ/93+IvwSLxJkx60J
bJybO3edAwMKk5ZX68rjWL7Zc8E//sZZzsbw4NIvKb/PQQrucIvgTD5C0Cew23pf
DRwaDloAftuLBJYzj7sixkVonstibe232P1a026F/H5illwbGRh2oW8hC/KdE1nw
SxEKeQ+T+n+KHfkK6nMjupb6fTOxxHYjNeP+EKExlrwvghbL9lXLbzJFAcfVS/DY
7EQtyQCjS0ndHZq1svx5mK4mtiB5OWeWj5TKn6GzvlUpt+CkVCwnUmFsBLG1X9CD
xwNFRA+xhlh+4Zqg7XCrx9IsHg5/I1zAFO9d4td4h7o/Ty5zoA+m8wzolN6ZVxC8
T2fjNaGtw9NXt85A5B2vRP+Vn9ZPgsBdw7805jn27Wqu2S48zm2X3xIZUPbjU+2a
84sGnW1nFvXRYL2lTsSPyvJK4DHLih/KOw2l5+ShtE0/HffXEnIV9LSpD+xPI3m4
MW6Mod2/2IDouGUJdvvbNV0x3LABFk73NRFbZo1a7KIWqegdB2F51THw71IGT020
tEo6rzgKckgXAUVTqjRGnrwO2yXIgUAV1kaYo55RWMQ6DBB4u0RXwNyrWCkQk+Fq
tqPj/KwBtYleost6UKXgk4HH33i3QFk/8gqtrkIF8Bd3Y9qLtPJioktRwdbzoRVA
auvYiB+iVSS0Yq2gpM/I8LMf0lFgF7PEI+X5+2H7n6Ekd34tpjGCkjLfre6rQKZY
ojvzztnkI1AWXwv7gi8VGqdJFUhy2PuP3n9yak4Mj0phnCwSEqI+bQHCFmEwNLO8
KkFmi1A5wB/pdw63edyibpTthzbrsYh7Xv6vaAZBx3K1rqgoNLvp6+0eQnKqimVg
c0na4/b4qled5aSBm8BMOujWViNOAlp/wRVco6QLnEaYohiwJORx3Gl+oCCorcgS
KVGzfYExwBKZ8Bj8v1me6pkiylYaZShbeW94VQphcRtAxEDbm3aXH7vwl8/n9isq
EStG6Z/3q0FxLOxTPmqgR5PycFOYc0+t2EOgAoHdLqD7pXOeeX8f6tUSYxZugNdg
7SDKa8VgMViQIklVdNpEyPX2X05OHlu5AIckJyOCgV2zgBlRD/wk2rI0GmjWlWSO
iQYdCmP9dlGUvApV9SIuwPuYp5LHIfbokO9BCOQzdfGdjeFQXWuK+oS4SpcuTimo
EUXgOeqhdUbQ/sgdqn2/bwqtkY7UOSByYv6XRI+TphUZAmjzcUrLFDBppmnL8Sdx
UI9gSffGdHC+CgF+juHNupave+/4LuybOum2JbqasYPD9aoQn4QKWVkbFp98tgz2
zoJcDGUO7RuU+pmbvIVvI9nlrbf6wOa61iGtkDhKnumOsHv9X13eQYwEZPuqSupb
4uKahndrXIr4YJvwt9X07Gtb9nCkXknOPqK0tPQh+hav084h00AUY1vzspnGWp3W
kIi3sP/dCNzzt3lZ6iKABXRjgZut+sgbglDAwEmndvIM1yAM1YvzaD3654ZUkew0
d1Ptw8is+SsD5sQyLoT/S8Xnh+9A5PE8gi6w5p3XYVJDfEFwZdMhoHQQazKwATFW
0tSYBvSQJEOQoi931GFHn/nSC8Wn1S6OCvj/EFARglp0trcXa1srGGwLio0irw3i
1cr7ENtoFnuXos/ZX65pLOWsUPyNYYolt1+ZIR4j76yxt3ZBH/nH4Lxw71WRptlg
Il2EV/2bcOREyKwHEGoSK9ph7CICX1+NT//p0UfUGjXaJa3Tyl4pm+r57Z5DuPeT
reuH7BEDJ6AYaK55hq4stDshrf7JkZyp8jri8oSswRvUELmC66BhLrdWQ2LZbw5K
6V92QQA3UTBuEUgO+hgWct0IRJJjinp1szOXr40BkK5nJlBh9abjL46iPILKIFE2
RFJ7+p6rZ1OZAOoHlG/gVpj++vndEoNZgzEYtl8lev7ivHeXw6U7IJync+DUGdOQ
EkrbMQApU9Q0DxgOgVpJC15UsBc/PSqTKYp3qDLkbF7iFd0lxPVT0xHaSIuGOGLV
FyLS0e60Ks0ZCXumMwL17kqYGnO7+CeSFe49Ss9xpgDMG7ugfoCO5O6592dkfH3M
uwPPrDGrZ7CgkrwkhoUB8fV+aigaIzsqGgSYzXuFZb0CY2upTIyy1oZF0elHRSD/
TkFFtJcM0xyUPU1GW4NAu7aqR3z73GP+Rj7uU8ju5GLaAhhJj077T6kp/LBr4Kxw
f/rPv+x9S9xuF0HVMGQUdvHmAey+QIvrwQ644nWMLf2Sh0IoIDe1dt6bTX3ikwbt
kUZeATMkqXH1D4rGDHVAe3nGDuhGTKwTvWbbhPpQ8mJPKavP81/DWtOC8FnWsbdR
yG0/NtUTNNEGQJydY0sNYOsgwlPW3TyRaVZF2jKekBnZiyWCcNzJxmDu9F2jC+LB
oQ7CLdc68lfvpylSXE/ZlqztJ71b1esQUGL2DkNo8si+sGKdvLpG1Zlw7yUoKUDo
nCe+lnd4YGalCg5qQBQoo8CLnty7TjVNl6l3B/wYMsJI8ibLmT68L+41UzdqbTMh
8CdSQNORrUcHIVeRfD0kISDo9ZMXUj6TcnjtWTsCwOtqdQIgbJEAJ68F8qxMwyL3
FleDiROqktDGC1StUJ+pGXKTPLfVywp3cATtymKRjj1lqUuPZBfAjFaWMGV9vWbS
VeyI4fySpXOrqcZHveGcpNrgfSjO73T5FLniktNqrRZkL86qZlAvpGdvxhxhjn4T
ZeYA3QIysK7WMRaplsGanKdDIGaVBRpOvzOMKrOYvB2yZQ1I+ryPOyWLk1wlpV5z
huKc04GjtXpDskgElVC8Km26qMwJoDsJE7dvsjV4o0TSH9BMO7vrMWJ4unquNp+O
qSftR6iIqxRce90oLQHhf+ZqSaCByrkT88mcFnTfAwtLs/wXFGrY64PH8LN2AQ+i
qu3ECqDYL4OkKsoFVUECi3KonqWE+h61RyHVhPPSAU0nTyw/bk+jB7Cj2e+Meprf
Ay4HaSyQ8KSFPqWWcQRXEQATGt7Rd8tMibWElfdBN4neWQCTxscbeGAZmNnL2blp
XYoA1bTLC4NZfmaeEWxFHtZrFGuzeqCFMc76sx+LwF/RDXVnnIZ/aP7tZgInwJ0z
P0pWG+xIMDP1yjIhMDnOpBjgog1ezcSiTXiMKdYfFxUsLPofO8BtRHftBfLsIPo0
N/7xQmBW1koW80ET0r4atagvIEP5ExYvCbSLQaTAliEYBkWEKvQhkZ7wE7mPH6Kd
dUU10EYiy/pczBtxJVM0S7ehzV5FU6y/ZUBn+dSLf457mEvmAKQcj5AsO9s4y9iz
ybMgONTFNOtXJc12egM4H/mvn/OD6IfyK2phYGg/5zyv05zYVoCOnKWzgZPfUXSC
jmaeEr5C2mL0lP2SV5eV5zD23mcCI1jVKZVvjq54GMS69XJgk+puSC47LB1XhKae
xsaYEjMF9Z4igtbDQWXBwhlI0htJnXFU7bdDB8J7D3isB8zw3hwgr6f02dv8kz9f
YqP7mbRlmjRsqcYOwS+TovsXS/UWmsUAzRHjZIYOqRv7p/BgC1BC+vG+dvlfM2vs
TonjU8ynoETKukdLWdzrcFeRz9nPUl4sQhUA5cMmEe83iKtFwc3I0rqjWG1oUedk
/kneVpfIuBAhuhz1YLVboJCBORhbABXSioNhtheEwRuN7yoenldp0zD/hcMdPUC/
ZU91aUWpJi3IAu/u+m8hFv/oFuP4slmEW/yLmFJg/cCaYm55RZXGOtJL921Zevgw
TGAn8S0kr8f5gTzzcrP5iLMV3PU/dlwKnVKSb1fVZqh32AKDrUsdMU50PnEsmZtC
9LuNbtq50Nw7qaaqTh3TuqEfY3n76/mUxDqY/LbTl9rSyY2FyGAxk+p4+YFWH3hT
5ST7Cic611ZHwuRVUeHHqO2mBSFJl91wLg6orHPiF/CG75pmYOTX0Sh78yr0CLY8
s8WJlkBsvAoc1r1g17uVA/UYeg3HnOU8VquJmnqOFhRUo3X9X2aR9KF5td/fIvjq
Qs/7jRjaPsfAwVfUXgz8WqjIEY+y71Z1RHQvn97ea/rnqVoV3dZ6aHiRx1fnud+O
grwxjVqYDmf9hmUE176dHpEqZZtNE/i9bfx4+33/uNW+/3g3QqP64glimvofRTc2
3gqPfRwGVbV6WlGdYJQI328FioEM+dYa08aOgQG6tJnztMB7SS20HYJ6Nr5Dhite
sNHSA0sBlUrTVrnqRfTHBb+yn1T4zsVoU8i6l2Cbzj4aQMlnIlpdJ54ekVKFTf+H
UEaR22YV/MJtaIFcDSKcmwW22Oj9WV03tpwdExqiYtnmBPC1RvrSSPkl3C7n6K66
w5LUCwZ+sEbPYNISaGrVE5X99wvcK0CdqtEpuQzOjrAVJequkZWToPlkwa+3tbtT
DjoOTb7Ri6i2GC5DlnoxgVu0K6tqyk14r2aHx5vFeQeo67HQ4jdp2BL3VpBAW3C0
DJ8Ks9lgMuZhnpXt3kqp7f+c0rrQJTxby0cCnaSce9sxryfZFaVTjFt5eJxeztiw
Z3dP258JxlLgOelff7kc6v1zZplyUvUhx/k7gWtJkM1aCtecorCiGwTqvOE+DJpP
IvW+b6SMv+nuEWwDwICs3skkFwHXBPM96+oVRRYHqRpIH5r6imPEh1CnWOavd3CL
w0clf1P485FYSBMTWs8a3VaZRgTd9hU5AVLf+dq4r5rK7Vu6oseub1b1qIynOOHG
Yml6ast9aAcrHjjWYI+ypHz7J/4x2vcOlZLny8BKEk+Z5p8cr8oqWomquujH71P2
0dEQOon+LR5qDN/JnqyKj+BXebqLaTb6oHmeZxD1qfcDv24v5oqGDa3SvRTYTnFy
2RJ4tiAXxPA3ajvoZi+phs4zywvIOmOJpCi6R8paX4pAPArb6R7yz6Ud8p3l8Q66
rBe+Z1SWR85p7RB3w2XbeiJIzGkLDmKC4pErxA8sSqZX/58dQvodVpiXqpwfZ0YU
wOSgd1Ctz2aJWWhWEzqrHlZQxWiifK5oXtdv82efIS1hlOoinUd3+2GyqYtY4LSJ
uJM0yEZNOA5rB5ADyxLgxsVPjsu5rr9QvfVFVRBXQRn+Ae3RYSu0QDXJa8rpg0/k
Oc95ru1IZco+ojNsumRKPU6ZQnhTE7DhF3aYbKN8RqpfMlk7PiAdW30+A88gNDsm
2BmfvfcO7ODNSBkUSxhXof26dU7e6cTakfpza0dSHxTB9J3swvRmuHkZRq3NLYqV
2ksmEGcwIaeFtrJKi2Semmf4URD13rnazaF17Suno4nuUpWiVfH7+oaSdsra8ZqK
nbo87nIr+pvz2BUAXsPuFUiA7TtmOJL6eCwpLlTbb2yW6iSgy6EZ9R/Wj0NoI+Wo
lQbW9ji0rczYYOhJZNZ0vNAugimDpsBY7fokKVHbHtwIF1WdcwQN0lYnAYp5pu5X
QcBkIxkOh5FtUtgQ/7+Bx5VbjVAJTSixl+R8wTjjbf8r1+nG8/kqYJNOx+4UD3vf
120LlvO+lxRPeKbzBCGG1l+jZdUzdE9lq+61TO9WRIpB6b4+OxP8/vykT0SmWTD/
ny0GIP4ru57fPktXDR5veOP7a2c7wdY+hwG5SuuWDo7wHfPyZ7Pibr5nRTrCdlqz
rTqpOaI10tO9EtYagQooCuEVROc43wspidz+rFgThU2eFhkTgu4+xzmUDhRH1Ofb
hHGCiceSRhqjzKJgNDzIkfFIx9egZIvwGP0ZPYH25UOefe5Nyly81rIQXxT1q1Ii
k1dNei4dyW3Bf1Rj2Mj7VmjGlz7RcHcmyfVyr/85ueizBCZN4Om+aAf4f7UINfl2
NIfWDZx1kN8pv7t7zbXbZh/u0VBKIwMvBtIUOUSmMx6FzlkGPpjorUdl+qtGMoLd
7BdFM00VLT1pDOvp0SzbE+IAG/dajuNihuOWV3qWQdm/V2np74QVidI9SEnuwLcl
zNMbiGqyL+zBsZ8mQKvScGNY2L+F2KfOwK+4ruMZHJxiL8QMQGBGt0z0D/yoON/i
P/UlGYdp8+YtfPhN9uD/+zEhVQOQntOMQUgeNzbn54llOBLxjeEjD/mdjq3Ug0a7
3RSDik1OP9oQHQAJOOWw8+AF5pYdZOg1omcjoVJBdRDBLDYfZZjKVCfzrO82a8pw
65EyEgIoFLd3aw+cO6NA2PIo8mFj9lcie6huHMv0MEoZzwZX5/Xk5seqiM7hWExH
Hm0/biQ1JJ6SoYaNVJH7Y3GFvvqlpLnFe/zpm/pbUkLaApPxncUeQP77T5IfPZYZ
SOSRvN96+iZ+Se3bV6zKXFdq9oHPK0tQmNscLwGEeBYiwWl/9IesU6L9GSF8IFam
K4sxqWp3ysDiKhWKV5DaTluE4UE3lgxaOaMiEoD+2tJ3+xQtZzv5bJIeN8WPkjCV
VSPB6CnWOlFH5XEptmf1ADMCAh5nGYb+ApAnnDGF0FSuVpHLFga7JG44pXHus6/f
NHBrhb9y5YilUFSjPnipr2/+clNHv5VW1GenORHO1LjsvL2yhKuBP6K8GrZpqU5Z
xJ5fGRSGjzsanOGzwJwNSoBc1NSnwYk4vEc8UD7tcsA4TQgKlqJvIfp7Yc5t4uvR
lE2Y3wQr9iyEx59f891BgpN2/2q1JUS0V09/4bRG9nmsWHDcHUMGnf9vwLBkcTQn
qLvEhZ19QuP/PlnVSYDyRHodXC/QYO0gI7fkH/YAEpROZ7hzUx01CqLcTTZLRtCU
SA1rKIAwjZG0cTJcRTh8V+lqljKXKORX8kflx933BdqPK2zcQ4FCszSD3QKWB1rL
NfaEW7lbVM07vsKsMqN1s1WHYcbxWBcWJO8o8KGYD1Rnqsn5ekPua0d8BpshVkUi
ruUjX91B4QJIEqzC7MDttUr/lFZxe3Z/jIX+SAZskhdku3moBFnngOIwVLz0Qr2d
2un6bKkVStk3aqIXQnNwkTSKNyarjrHezODxPOiKvmTbyWJV1mMWWzwjgm+Uf5Dn
pJ+SpksNG9v4ZOHuZexzAZDmiw9qRDgZ+HndiSzUGyv04kyM3w+FL4aAJJKKm4Sy
+Nh4fhd/Chf48rCHZh5jdnPygmwiogSyuo2EcX6NEQCmvSLF7ec2cgPTZLvb3QR4
8sok/keLTh1t27d2VNn2D3pzYJzVw7wXqdX3eYEeg/JBj1EEpGGxLSKzgfbdKSto
FrYkeK0NXyXfePON3C8ZIMxatyzHlk7dDmSXV65PCK/0eTo1JEg3RT8w0ldmi7Lq
wDo/Pvpip+M3pYnQiYhasomO0KcnCt4XUwmlDuT83FJdUV+oW3aO+J/JLjajVTt5
+b6xDixyuRTwb8UE+xpUDBfkk0X6UDrpcZIOU6Sb9euc5OP/3mSrfjNrRe7rwA93
d8aV+7viq8Gik2UROo3RMfvO2s4/FhwcJBEfqe04TsV1bm30zsIyIWOP87UhjQ2N
rzr/Hfmjxkapo0nOQgTWgCoMgLR68t+ScGWvEN2SQsO26JeQVdG/2wwc15C7WpyE
6JhskClW6xCjQKZL2i8odM66Yj6CwJQqIDSoM3OaqYST2M6y4bILTNKqN7eJeTM3
pigXtU36HpxBOg9FsZjwhX53WFkdNtXXTlbzfiXCH05MPfdNa0kqB/31QqdGemKA
y85p/tpBVGlq9bOagN+uTAOExEfFSWcuuuuyHBotH6qMDgVFoQbyBU2eRiIiEoxE
W07adyh5ItIjrpNM4l60Yg2bPfHQh23zc43RM9p7MI+yypNfAkny03t7IN8NDRf/
TJA+7oeS50Hsk3vUl5/Zoe/kpq3azNFJ42PH+vcp7EbdORy9qPL0M+i07X0jdLyt
5CIgex6DIzRoGM9YdpwhzaEkkJODh6cgAqlZ53GRV73qbQ7lvTxuw+q3SJxG0AI6
Wjs3ZV47dUlKk+MzEts7Wql5SXt3Iss9agzoJkD3wIuAUdny+j7d9ujM9Z0XhTtA
RaG5D52gnSVGuIzmZPku6xB/rfGlemV3mkxi5iZD+f9TMO1e6xHWR9kksNBnZhcv
SlJQ9xrtzmRoxOrxDYuKnKQ5NZVIsmw6yYZJo02OFqyorFO9UuEiKGq52vc1ic0U
ieiRfNs2V3aA22JePKvaYdcfYLtVLPn3aRq5U3qtETpxagmkvejFKc/MMjk3sAUT
I5elqVRDhqpc0G3Ih/xf9jjXFYCR0tgaGVmwXfsKsPE1cTzvAYR2c1OnSI05ZY9T
f+PK14AXBYSYCIaylHkg0hDuxzS5qRPJihpauzYV9xEmw0GAsq76mjlRGWKevHFt
yFdHJKOfd1zIzZglK/Y3dn0gpI1krVgIWbPIApdNbBmA4wz6Y6bd6+UZBMeWsS54
Q/FG/BCSZYSPb1n24XoP0Hd8fTjMQANCXx7VCBMj37+RmBr9BZIaW6qMdVCzQTd5
wn3zS/uqbhkQ5RYODJdwK2SMxwsD9qrHSK7YsKNLXvm3daCwMdyaFbwOru8khuzT
QNuZSBqPuK/gEnnih5U34KC/ZLQqje+gaIMO5xNar+D2AUyPj+6bj8n59T7/clIP
309/fIPJ8bASfJg+9PkQz5zH7pVTPftkxtHAQHhN2vhJud8SBYIPACW/oj+XyLIE
Nrq4cLE0Bl2Q2EXphHtO8U1Hj9DvStxKPsIcKK7auoBrem6dVgN/7ggl3gGbcFt/
0Ra6S+gwois+aAltR4Hc7GWgiIk7+WFT4PG0TxUjFumsKFIKfVdRIxMuRX2iDKJn
v6Sb0LRwiVsgWgUb3K1b/zwh3pDPrRPkA3flv6PdpYZHLQ1lmVLyL5RKdyzJTvDL
q3P1i1KoOvhznIDzfEX5Q9n7aEYQ60Dxh9PLtLtCs1o+wQgdIqZwa3/Y6soysrLk
i0boomNoO5eUvVoFM8/5xHGwPiG3VzIahNA8ApcewbcjR7Dq52NneDfaROO0yk/S
dTUc7X1ANy3J26HqTNmNd0pjD0iY2UaZ2eOQQlFaplXwnB1kAobweWnnfj8KUZqq
6WiRmk52z1+eEQgKcJDfVv9yHlPpAw/0cM1Q5aOk47M3z6XBf7e5kHP1CcD1i6dw
YrwaK8+e8dTZQKtCqcQVwHeufo0VrvxfBc56URPFpSTQAEKbjl77rvAPh0nIePTs
lKdRh4zvkuWWf9hkhetmkMY8HwsHZsnKVcU9yLAt1/4NgySJ+SSXp7rQ1N4xsDbN
NrCXxCXJHtURfUrEtq4h3UPQC2nu9y3vEdtBXyEQKWAmZH0cB+LIADRGa9QsQh60
mV0Pq3/sP/3eYOpy0qt6Qq5s+XUKyeRI2mkoTOxrwZ1LtVFTb68POz3xQDfXt82c
HyAERzXPM5Qs6/ynBkI9Jh9zLC3coOHjolCQoSe7MztpNamb9R3ZO8+j357jTL8E
9RoZsDylOZkdteeeSZ4oob4NJ00aog9R2HuMXpEJRJs+0p0/V6HtzdQhZttYYS1d
OeOhx5sbyHZC46RMfWLzVbGp/GTznFZCge+xHbvqcVSG/QodU/e4ngnaKk73QGM6
SMAQdFJXXmTbM+NIPISpAYQB5wU+1QQVt/GtETMO6AE5eGwTz+9H842sL6KUpyJ9
YV34dY5AhU+QXN4s7m0yhJkiMMPJCAX3Ycu6S0wDqV0QzHWoCoqpRI69m1RKk0Ja
rlq3bwEc9LJu6nRbYeXgbE3URExo1qALrhkujdkymlHnrz4Qsaf9PYX1qNpsVCqq
zN4Is+E//tkW89cIbB25UjfGJHKvy0tCPN0lYKWaJUuJkyrD+X/xG87jb05uQcfi
Khs5Nc/ElJeag9KDn1PhQgDWseius1zdd16gsFzAVYLR+IdD0BX8UXCaHHt4JeWx
sTp2l9/wBTyvDY0JWlf7Kw9YydcFFqlKi54BDeHjQYyBsRjcFSgma+9OAVezvhDa
WcK97LuN446rHZx6PxkHaCXCfA0BbMa8mgkw/vF9sSPQza3J4OeUBueN6e+8Sgmp
/Ozr6lTvkJywXq6oiHMNSWpyo7OBvJzJOYo93RJE0oFx76FK4HrF1KqPXW0FPlva
ip5uGGT7p6uwrkRzWylmZFL7WA59gionSqoD65FVsRpUjCeuPsuoUIG/gvXzlyJy
/esvAbrcJ4ikT3gSglYWOJt1NcOxKCWAgz4wHWgeKjTU7Crzp+TWAaYIJmoxp3B0
WIrD2Ef1giU6gfPL3A0q5xwnWVn7Vt6iFT7M1I7L32qg1Vc4MMU8L5kCtWGdDetE
3KViNZFb9GAa12i6/qiaZPleER2DJTpeiSyPPQsuH/NUFlpYz4IUh8XYw3k9+Dmy
hSjC/iqtux+bb7xeiLVGZQzNPWUya4H6BCpduIWYRPKt21W6VwnKyfjRKWriG9zn
XHoJCxlg8obBZU2fN+bSsaXYlYfXpLqp9UlCT/T1rsEWrc8Du3GbbwvE/zY0uukp
v4ttRW1msJQV5KqC3bnR49GNtDJszDprcri45hx7pW2WYoTwP8IksY3X6WGZji6v
ep+dzV0V4Tt5OAEWiMh2Tsi+48i5BCOPZD42r4aA1sjdvHWJR5DgJ09CDZaFutzX
lAEhkg6eSp3GHQrzpV273Dcuf9IWFyml8V71fA2OFIk2KTObweAQ2jsDFqFj1ngi
KsDszda3aFBi8BgEPjHjrfKcAC+U5ZEEzQSHbROlvtIOUqBrKtLWOZEyjMk5dLEA
vsRxEo1KCsT9EvB2Ah29t7CTPtE/qbBxBi+aA1Rcj7F5onm3uXTDU50JI5Ejwk6L
5lcL2Wyy3PCjmvejgtjFOHG/QCI8fP+77gxQ5HpM75SGIGvCXuZxs5lstvY+TMbs
srsSS8czrEKHfrIRMNgqLWJIZDrBzhU9FyPMqX0rvKVDLLHN9Aie1E60nG+HbLMA
jV7RUg91Oo1/+msrr0Ml0ZJI9GkDHJAcEd/RjVgp8EMFpYWWzzcBje4EjCtkUd8g
mbWE/ukCrZIfbOWgvCltieS5ELWhWcWumECKljZbLNi+YIuDRch7OT58yqb8oj/C
ZnYW+ZUEiLOab1sojEU52uwMv9bb6q5AjICmpm8lQKYVhuMxks+X7fjF9me9cRKK
BTrnGc5zyRONc+naMwT/I6T78ymKzjtnZ8U2ckK55WK0NV0yJtESYnqg02EBDjnx
ueLkgBDoIl2lK0Q9mLoFlPU5BD5pbRnmZhtopA372aLaxtd7oWVTUURz4MGZuuoO
IVx7BwhCHTsla3ZBxAl11w5xx3rjdOX9a/X0qAZZSBLPwkmXoMhUz/4T6SXTxosI
WR/dUCn+ZeqpAuTb9w1mRZr/lmt7n1/EkCvf2XPQyecfb/aWyNzilpszDDHLwUEF
ah6PoUvV1+NR0mEA5Z1Jnt1eetVrURafBtGqdnK0WAIyXdQ270SUdmemAEeX/Hjg
qy1DRFfNCp0O98d9yM3RYvM0eaXl4kSRoLG/fk+4Jkokrmr33AdpVbF1xMjzCRb/
DLE5ZQLpfRaFji4sfDDuoZ8J45aCd+46SPe5iM4oH023VcCco8NQhWc3eUUQmABf
yrw6E3PWCCM9oiyJpuR6Ml/ltVDtZs+uQvTotFa4cO5i3wXldcA2xMyDffuP4N6H
WEz7KHdVtE+/aKoVD//hL2wVRH/X0Z5UjLzqAgrq82+lkcOIly1oIdFpAaJIqxH9
UnngPnNylstkm5+rdh5jj34LwyZhQqthsV+pmHyc4VxRQ7nUJlM/V3jiV8SrlgBF
mFquwmSS3kkdXlrJRoFWiJE6L5cmozRz7VSdoFACtnIiocPjqsNM7QQk8u71Uai2
CD8PIJllzUY47ejUCTal1xsz+DxonsS/Uvh5UqSRDzk4Gv16g7kso9JKxfIkCMVG
xTdsRjPzw9fgwisy6KVbGA0D56eq+8kfKj479WxULjW9t+We5BTBIDWG10X/c6dP
PGiR6vMml5ovOacpm8fjNZdcgZPLTARpQALN/qJ0IvUztr7qBR1RPfUeKJz4RK3U
X/CGpwgQwIN+A1vw0xCYh5/aXWkK/0V2EFPoK81RGFpg5OsciS9LlOXnSt/mdQUQ
A1fXQ6ooZJ9YFcEMy2K+ZzZ078SjAaBfOe6J+O7l0eoRO+aSC/OY1zm0n2ID2n3M
+4PUPBvlWhB4Bp34i/RtZB72kUYV3RPQAn3q4Kv0QQyY07vR7sXXKAUkWzCOuu6j
7zQrrMP6+TKbur8RydAoHQfhsBXhR2CQZZ22XsXJNoTWlxzh4aBMmBtv/S7O7sh6
Z2ijOevt2Sc+7a6+l1T2HdRZQkKeWzBKbBqL4K1+nO7Zf5ZefivTP0OvlFKdhRqn
hwEkF41en7cVFYCtHmu8iqfhBlu2IooBSE6ccjKzLjdT36Q+7WjQ+szpIAKTWLpL
4bdVZco7cruNGKwaGW0y09LdLDwCdACvMoh38l0o5tcMChZ51TmAfwIOV1OfBgTO
zSe6/qWByZ5/kMgOfI2jn9a5xcVjKoOgl5yn9sDIMHDk5lmagv2Ru6D6rPzPsojB
UF/Uvj30ix3Uu7aWYblRPirNhAgZnMAxa7T0L8n0yv0JZAUV+bYSPzj9pVWLeB26
RXs/jtXyVuentzZ2jacuNee0DTw1Hl2KRKyczd5dB89cTlX6f3INkRobQwxsrBgl
hhV7cc4mMOKmuGJbabMFLD3CqPCR2e2gRthEJIqhHw7DcX6BQBFwTLb6YXU+Th1e
zIFcxfc22j/W9YGffgsGpapcGX4Egza3mPAhl88FQRnWhwvtGUEF0u6M+jgsF0r0
olpy1Lkay8S3YSfoufCEhvPovmFj4hGusaQv8KcjvH3XzmS9uzDG+y4EZRZ2+XUe
CTCuJoO7l+aBhIRLDxB/QTA4Tq2pd0dLAp1fx3dNWqnY4AiBGAlxdYkOAoPQoqCZ
dD1cVQ/huqTzgm1y4HrMi6E3phiJ/xqZzFMfD0XamPUMp5PcYJnxJb9YXNXcXJih
K4VgsfPe06tzIp6GIP5VAdQTjFiqK5oK1rgT+LSUrP/5tAJsVnC3ymxONrbx3HJW
z2oyI0+2QTOEng1oyioYxMLAbZ8/P5q2dPM06+7nn/xLCdc6YleWw6JhXjxqTiIA
mrrx8i+b/X/4gnMSpFRulmz/dFnS0Ue1oosTYM8W8uI3TQEsV5zjr7bI+S2OxIHa
k9SxkTi+9KnP9WQQ5A6VUJ1283n0noUEiTI8AYpXoffNAMDJ8JUqe5g2rGBP7L1J
Us3LWICUUl1Aw8F29McDT6sBHIg6Axa37DtY+ax3jsuK8J7l3S01yAoDnouhcVO+
oV/Ly4XrtEqSde6TLCwLom3jgHGOYYr+8IhGhzyADsxa9QlhFQI/fFoF0eu8CXab
h4VhwIfIbgj0oD24fU2GtTmC1ZkpP5FN3c7Zf1S6+fvkQq/nB8Obpb68zongRWFu
XqoFnbT/KSmuFcyNHwoEe3Nb8yxqj6qdmDx1KcAhM1GQNVcV2q9cKZ1YK5z4YByG
Fal+vX/8gtjXsLCQQGyeddyITRvUYpteqnGMdOgAim26vWOFS1k5SWQLRHqGZpSE
mPZ1Kp9vgQwsfSypWOROlRDrs0YKfUGLouTU+ZELamxfxOf/xWOXVltdGjke+DFn
5Zxioh13gIso0WxdpVC0yZ6ZjLOzWe+Hn5JDCFVz77kgfyNsRDmeJvU3Dbsn8Xi0
4zZXdfs1J7EZSO4wz2kmPgdAiACtMojKPV2Jhe+J+aPXgnS5e2y2G+s7K8GpukQG
kD2u5FCe7uW5/5Kbx9RiQQcDrJsEk1UmkaDHiPyOun5FWzWT3BmhqBW9rlKqP83E
YKLn0epCBkKfzzJJcZzrDX46ecEjOmYesxI6eF+AgRr7+25DyljGPoZ0S3D7QXyy
THZL+pcEHalJnsakJfOYC7VTmNOEkM7y960JAsNl2Z+s0ClPGkgc4GJCIOY8sUtp
wBsfydG7iDvCQNRHwgp5jr6Ap7xKHO2J05greS+giWXko+4Zcf3Xd9p2VFvVlnO1
JOn04pNbvuGZWh+XXrEnBTYRRK+SESzq9wRjEbYu9817DR/vcq85H/3eyKw7Ya06
/qNz3F8b4qmESoxfOAvny9dEx7Hpoh4k5mZcBy3yDljQABVcsUJdYgzS7lgbDmXE
TxQBlKc43lZa2DgS/UR0Dovpn2ANa/4dd0EM/m5ngv+T3VFE8POLYNW4+sx1qQZv
PciMDSfjVmqkN4GKq5z4BlUVdVlq753eQ7nUs0g7NYe3F9j2QyjQMl4ok58Wefhy
RLN5ifLkfMI7Ob5s/HRhIMzXm3VC+mgPxAR75EO6PWD1HPbliOy67RTIMjnIeatR
38CHsOaBcjnFycNxRGNx8giN2hunr4EAtf6hpRVa8GZUL+lwdELvYVSU+dPNYFHm
Xog5Q2xcP+E9f2o2Ms3jNRYDwVu8dpW/K7Rjb6RTjcAC0MF/ZwlZqs72lOtomukl
VGkhjeto7jdfR0vsMVmh4DcYjbDoUUQauEmZU4ankzwh+x6iskEFkc2Fpn8I2Rzy
+z4qMkULUxb6zjgi1ks5xvKydtHFXJ9RVQT8PpCanWZSqzaCGVzPEDRaTW7e3xmK
Yc01KdmxEUZa4oe1Hau6p0vgiKGN/uE4JzwEXztNqJR4rGf8+n6xaYkDJbQ/CD65
wR84bRv6yJt9Umgj643lSSCoDhDgGZPyqYIDomHtQ4wixjtrbiC39VKguqLp7BSO
6lxQkryvWxaBEGccqD+z8bB/9uY0yRxDFL5V9d4sfvIFiOvrom2HH1Mc56+n4vkg
en4p8rgCuwD7q53mjiHZSfTxptaSb9AFfmzg1+Wa4KFqAHV5Sj7Gm3pLm8BSqYs6
tdB2TZv40yF3KJXZBO8qmGwlCOwp9ik27xXIgZAg/L0dVjryHaeC4mqFvmqLBXXA
BOTfT2TwN5QaDRWRZQ/3Sg55VaLLo+dVv8eI1Yj7aT10pkidcMbrBtWhHZSmmQ4m
TrU1FuvTWeahcZ78Hi8DrCAXmYWw2gXYmZfbO2mOR/VQ+oIXGh3fJm2wRX7DPGc1
RM+L8e1gGYd4mbjZ66uk2zJwK02jW/RmBAGtxAZEudDbiUdSa0EuctaYxT4omZds
z3qTZ76e8ODLf8kukyOUoJyBl5iRYO/piZQjRHSVAI+U3hukijHvamioY8NrcNTW
yhIj7HAMIBzwhjqUKPlqQ5VA1JtUfVSrOg3OGXVT7xDZfwJ95nwhahoet86eU0gb
FclwGE5eBMAgPEposmQTp79lXQDgxN8MzDR2gDNXB+jQrNxFnU+eORPiEiTdtKcR
CiuWD9lp061g1tJAMmF5tTh+/oqBlnh3BBLfDk9tFiky6FBFHUZ3AglX2N0KdoQy
JcTbW0ZW1D31Tdr3s4C56KKANEd2KtSTSGxvhFQmO828FujfwiKzkpZeJCF6/HFz
l6lmfVj6RvFsaM3dkfVLhTrzE7Fti9hKR4Z21Uw/FOvlyDOzp+gjtvJ25y9LLRxV
KMz0DchXYsbHqfwM2EAcrRFANtDm1fbh95bkW9uFCREXDIIY2LZQWc7si4LbIu+6
BxmbzLY1vs2t5U3GztCB3SrOOYHhc6Hgum3T9D+wrhKmbUvNpYbjyCxqZJjnoxz3
bOvvD0WuKvD/1ZWqeEQJLkx2w+RHY1TU/gaYLRUAIbEhJDc6JRYZZVWFR/YQB9Ve
0+ImFw+dGNn0bFVKbXuDcuRssgjvtcmeRMRA9RTj0vq6PNefK8iaRyNWcTzz/Lk4
L8vWixgwGZvLhnb4mgvoxOKK6NCg+vQ6HvASQwaaqiVWzyHtTcQA1suP9Gx9P3k3
wYCRx6/udHU76k5Q7Hl2Fv/8byW6W1SD6lsFIJyuvfiuE9VR0TB8bMJSLOu2Jc7K
ntCWXYixyb8sunJVkqt5LvO4R8hDQnbPZ2DxCGF6sADuwlQb4k93gY9zTS5DglSI
wn2ZtgJvi+CzrHRDHW+vsZiRyOHta58vlb7trHC8Z/TMPJAtEizj1wdO8uCnpohg
f0zmWSoFcCiW1ytwE39RAOXkHTL3wQ24QPJ0oIKXS4becipZuYJG3cJ0VULoG0jD
i7QcVp1OfvEzWe/Gfi9ujZkXH97a9gpN6RJ4q+UKOS+s5EUm75hz0KwsvMioHsNI
PDqnYMUKfYd6pFtZkMIdhJ6sj3IdVWXIany37FRnHIy1zBHjjee66gWtKVdHma1L
xCrRqiIm866WDhMUAQXjF/Bi4wUxLrswvU6bwo6wdY8D/NSJ7JBoPy4e59WV3RYs
AVcoHNA3YTH5V+VH5S5F9OINIqg9OEr+B8Hy2/JvAQZI2Fm9eEgjGHe0wjoYTJNM
9tCaWE1EaZpI2b3pAZaAT6hBo4XVszuDH63GJ+zGEPp+ESeixoOrFD/TXJkRhBjw
6qLTnJwWPLm7losyrelexy1iDyGhrJTR6nQx6i0X28TeFFUJg1BPbDVAHmTbY99f
MR9cv6L2SbF0Vgo/FKvHGlUy36Ky8BYVNYxmJTc9+47NmynD3UqxXMcAdsmUpyzU
Z2jCfeBjbgFAQmqPI7OaxdQEr30qQ7gtrvi2aA+LzFKfoajyb55NW2WJ9V17ej1T
5BfRnomWryZ4U1S9DPbn9TpIgPyP08ddYPjXVCXfoYXOg73UCiVoVeQUY/RJ8LPc
CGX6q2ZEB7Uj9PH8C9MxdfVuXCcIMzVtjeCz7ni615uRL+MtQSYmPb/mAMGkKB6i
7DUrhuklw5/laeG/QHOiB271K8kltYc5/mS81XyL1PgBZNG0OkmfDd7a6Bxtel/f
GFzPBmI6CkNtKdO4VDSRr/F6yJGMm4CSCUI9cNkjZsrBfMgwd5FxM8QnxulQz5IJ
Mb0dNVwQ4K5ehE2gPLAxkXdqCDdw5Sqi4fYbprwS2NXZBpBxIBJptmLmP0NlEIcm
QYU1eq2y44W5vd7yZPJSWbqMIVb/fzByE2JKJY0DBffd/U9CylGtOLg1ZVLXs6xa
S+iZ5nLjExmV2P+BNweAjRnAMQ4pVnXCPT9RPpq/rF4Xk8/AsMcjl28tj26eU+pC
Dt2IkvgusV4LpnpH+dCW2EFh+ZKHtCqSpAJyXvvkwora9aZXw6FmmOrZNUfo4yNc
buHuI47IBOXKa2zZbM+pwuDoYtghLAezDI6xKC8qW+Milu2hgkFXb6g/Q04Crm11
cZEj8CQvBP7yg5ojDXz+SvrehYwLNDYcyt3pkVmV1PNmkIx5u48l+RoRNyw7PQee
EhIOLsk1oG6eyfEZDa0bZ/44jbRndgWo9bRKX86g7P6tmuhWg/xd0ACpV2hU1lp/
SkWUhCJMMY/XHcZduBJIgWe0KI+VDha8aQQ4Jmky/KPN4x+pFi+eZ+PMkD6HeVXJ
sI2PiO1gFbrARrb4PrsHmtJLCfWQCyk6Q2hf+I5VUY5q/YO6P5FFUR0PayDj34Qv
vgV8nBlOGUFGSL28HxxHFhK+cWZh8iw4QASXAsd6w8mkhZ0pDRhaTAMVMDEtCgb+
OcHMa+eZ44z8DfffEWz7IXzznUKRL7Zg7rIs2Ns5rWJE43IMa3R+zrzqS/Ge9WeR
tT4IbWvkir91dZp4nZ7S+bb0lvrUmtSwGbdg8iwxD+tzBiyBPkAEsEzj1DZgjLLT
nbZRi3ccN0sXM98KUWy2fTEzptk0h4/MOMfSlmI8Pg5OnKSID+2Yo3A+JNq8upk+
dVJQJAT3aH0a/W83JxZGH/lRBSZZpvdXhR8syRuCE57cfrVJynce6BO+jfUQiyAI
MlpmhpU/HWlZcCb7oiFQzkyTRtYFhbCHGKCm7q1FFop3G090pAVYdX5rCmCeWCa6
6HTZgNpG1qmtzKqq/mjA/TqFxxAWRP98fgzBCHucSrHhv6bSHjiYxZgRykG3YYKE
tmblo3Dku70pYWMYkP+x7J5WDBjwqyj6/niQzK16nnED1L6NxQtybl5Qg+RRlyy9
OBYGOHq4K0fE1M9psklgGU1NuCASBXGX3cpej10iOH8tNQXCgRazOx7Oan2hcIeb
SZ5K1l49JLQrzOSbPnWBC3kg2cYGurW5BAiYVFH+a9SBcQTzhWb/+aCQmC2evNvL
Bu7fjyPnUoUjKaf1i2bSmWrHCW4ht28zI1H/qPWWW+RaiRpTxDT2uA31uu6weOyM
DKzIMp//YBWWiWFd4AGPABg0XONGCik95E+h60eqT5qG9XOlsUQAF16fFrcQxaz2
VNjc2s3vfgBLtNo6eiGzTWuQaduwy+yJ6NF45uRwxi38D+B5eXx6U2tYCzgxZS2F
oqs8VTgBIcVlAKckpItmuKaK97SkWz0GFJOan9AenIwP5QVMmsklitt9LTK87iBF
khoKx5Q4UN1nbQRlPdifAl+TOxM1phWKAvV03xZ6TiSFZd1a49x1R3bwD6821895
kBa+6/NBQ9SOygPTISiKKEJzKfyRXurN+zh1eiUfL0vrYPL4u1+bgpvs62YhO4zL
WhanrHSi6QUCYYoNpqBsV8hhgEIZw5MyYJ+bkOW7PleUMx5HwzGv0DIbehq6i6PC
GumtpwraML4k2i2XPC5Ghb8361ExunzTw3lzDCNC0xKakEaw69oWeh/8PwLRUEd/
tSD3q5wqvap93ILKKBGIwJQF8YxGvREqlU8qUeIQLrMAMOEU+7o92Pf5R9qAPCgA
a9lX4myGMncswIadft6yBTtg4ZMtZJGlcbXjHszy2Y2QEEkTV0Alpxg7UfJMayGv
N8NpKhryaGOgZAuDODSU0CIIfMzm9TzaX74TeeXtxcBZNeXTZ3PIbRBYgnTBkyal
N4A+YHFrT2AO5r9BM7PZbN8tML03Ch1X2f934nJ1eiR42XNPJWS6Ww1QByboRMq6
c38IkPxbyHGbDvchjs+EHK+TSmKa7up+eJuAfmIJ/1zM750BUomdnja0SncwjD/T
j12varo8g6UGYd4+EiiLIkBYhHqaWFhKhiJkWypMv1x4zO3Le0hRAxRz8ZacH3LE
QIT6VCKj00BOPLvuwiQ3D3/IYNaBfrG16DtY0RjBR2t+hOKFHJSC5K023K0/EXqr
zXZXltd+vP/0XBawHrMpiZ5gYipx8HNMsRMuf8KL8BztVOm6/fyn6T8mD08HFDS4
VgbaeKMDzJm1u2EfvyWSCxmdY9AbzqoQjy5NHQgZS3v81DaJe8zcyTOstsYIfSfG
lavKTTvdfKaARCGBzIIgW8f03EAaub+PPo0R/XOwhKAxT2e6gr5mMwqfySSqRhVX
3hxJcVhTcdHota0OiUgNFZpGo2icfE/krc7zeEKqdOSfULQXGNU7s6C+jtdqgDPP
7aQTLgUt7IVF+mkWfhSgH296/JkntMHPNJdIBi54WTCKWLweZsVWH2gmKSFLp7iC
WmTtQfiy0j7O6XRtfj2tfq5E4DdWQIGZM5FfGDFEfXXKpVh0/aXh+wPjXo/Hsjxz
QmvYlLRLXLIjGBki5Ro4FM50tWgGRt04Fm7bTrBnD0LZALii014NlnRTzr+r0pgv
Pf4MeqP1AXiv6sToqRb48G1/00SgYiOfCnC2iEGBBg6K+1znrgXnWFTJx1wFBBPx
CSF0CO5E1B1jPG8CFAimmfDebFFkINn+kReIBQD7TMWZPN+f/h2UckuzH8s+OYfR
4vLqlEoUh5SYetpaxQ2kDxgwPuvZChGOfJcAef/qdRNrRA/N9QopFaveeOaRfxP9
yU8Dpuu39MZvDr+VTlLiu3wtK48ydTZf2ARyDSTsYWOhb1ja0Re5eIGJLW510V8n
8YRp5GLKdjvGDH87gNYQ7Kcm9tQgpbFa7gtwZBXWi2Qg0ayNSCGC6Y98lUOWbPuD
Rjmx8yPW4SaW6yxahCjdDC+fGkUbn+lqdo8EBtNgOHAHHtLVGpdvqMZ3gpwQ9QHb
KeVNOiM5azbTQTimDeJrAKbuHsUIZP/sZMYoS8S2gc6n32ndkRGXr7VOcDrtcS6F
Z7D9Sl/1VTtJNaefN25SYAwS88A+o2UPoh0hrz43E4wPuPxNbEgk4FR1w3bLt5QT
fzlUULAKBJzQRNN3Cg3RNIxGSJCbivfCTPQ5eES1eRcyIRJDnXErui13e6vTIyNd
EeyHsSNKm6f5zNRV4Iywgk4AWJsBzQMovePFRdnmo11keRb6vVhSFu+dlte9Pyk8
F5WbI4CitpNsn//OUFhha7y4329NDCROv3cmf/xfQEkdFyHjkUeq/QY0c+AXIxdd
wVvIzWcjcfSho4H8BA5KGqNL6j07V9hE98rygzDz5CSqYrd/esJ/tlGnMAnxC9ot
4N9rQPeMwgAjco/R4DPBrjqHcVa0vpNTsnLqkqwNPxfBu6CpNBV4EqaJh3j+/BjB
CmDp6GudHeC+aulqd4Xc5lsXqNPm8hAS5smzHDmIej/it8J0Nq33Gf4DuEfheYcB
Hkpyeb9Ny0ca4uQT41c27PVgGoBt0tMvUEFvukkuuOyKWV6zMRlZP80mOzgHJhdO
XgBSTnfpP3V80NomFaZv2GSfi1pT6jv4b22C53SMuhsETjCjwaTl7opTSTiJAd8M
881Kh7biMjgOyUGDUZ1e0WaE8If4ritcIWCgwSYhjHduDvFvziVDInbtVBe5KmVW
F6WhWUKQd5Bu2r6/C4q7KMZUytqEGzI8Z4CXbBZeYA+BYKwZDLgl5euvX8KoXg3z
x6fs9mhRyig7PGzv0JS7dd/1TF2n+5//ZoygKeijdjxgfou6csS7+/j/5qemmUkf
JgB9MfHeVobGwju9TtsHLWai4ZEFREbNAqpXXAW3By4Loq4BbN0xOKfyE+bnY8OB
P4pPZKk5E9yqmzDXJ96LRDPNTsuoXmcyUr7VPoyin8CNXK3r4gAvOYvsZXS8CJpa
+LFyx7P/GEC5MptGmBlEGEDDMJ+IpcSZPLdfCmKWx4YKP5854s/k5TFfg2oETfW4
M2iDtnI2Na/Zk2+/227Wtay37AYwBxEqe4fD2Ws6Lj+64DrVcf8+bxEjA2XgCTrF
u4bhtIeDv0WB1zvwen3YMx1k96eJ6rVhgTReuRcQEFRtMZQcVWlLd0saO0JS9p21
H8matg+rxyxG7wHoaHlki9TJT4T4wJvK6Q+en+/UoxFhklnJ8qWerJLBWv+lJTeX
TYE4d0GLZLazxU7WP9SqpJ+G/wP9WVA3y7GKGdfgN1A8G33537l22hRMTcHMrCfK
RP0uX7tPa2xfYJS5U+ihBHPlKxS1EBrm+/JC3lqBfWI9MDFcHY5C+Rsguw9ppG5u
598+lYZUvqF1lPSWGh8dc6ne4MvtERPqb7D0rUFWC/Zk1Nfi7SplHGI+i8SwZFtT
euHEusmuNmHComiz40csi/bQQAciSc6Am8ct3LTr32oopUbOaTs4mMYZzE5IV5aS
EjuklMchmQkt0qlb4ZWJ0WcZHL8BZL+O5Nlxi0pqW7zrFkPMTPG8UExxWt1scIZT
XW6kVwmowkhnrXHHzNhFyyz/KFC1KYC244lIERA51nv9Vj4TXa0CXHmbuC9h+dYP
owhmEcAwgULkLF2ziajZjyz95SSiH5dxs2I4XS9Y3wm3MT5eE/Oqe+N+urs7nn2o
Es7R//dAP7a+t23K6LvW3rgMLql7DDAOnctvaOsfEObUaqN5QrDWxMpPB2ys/MaN
XsofvzbfASm3QJADL/WlPxL/7OEzyZFQvHtU21nu5ACIutCr2BvcVygPR0l6GM7D
5+Yq7gtju4uiOR3F/eBllAO921AscvZfT0xwqin2Awir1VpLnoeuRQlEVDS7U4t3
diibFPDe+v1XBCKwG714ElSAyDzqCOoaa6vPgyOFsRA70FYpqsUoiZaliKKVvOph
Ldx1p2lR9XFLAH2GrcLdy952ZAnIkUKpFGmXHbYgaKwYCLhfSlgn3/QTBMcXlhvT
BHFo5OPpd0Ti1+oFUUm+zklv9RKdd1WgAhTj5iC0SUV1Qkj0y7y44XC99t60OR3W
nK/23YgcowkfdOA1qV5Z7RWznQ3Z0nxqYbPymy8/933ej+16j1Hnw+Z2sIUESMWM
1xJUWivCvGA945AIMNXyrldPhk2eoCcQhfwecpMB1c80mTeWVSkdAbHEv9gSJvNl
hEle/IhSIBtY4W5VYZpVXBccgmN8+QWuFLYHubUFAWn1TDBuxNmTDfoHgiwwYh/2
/i2EAdbI6WBDHD/LfLwWh+aqoDtnsLOJJYVcew85rjhTf7x4MnaxxSWnte+Gq2P8
VC1TTAkPBPXQgZZsNQmrpGSDZuCsJC9YvwUzdJ2WJKF3eYXp956peWcryEXUXidh
z/hPoJGBsu/RQZVGN3Jaxh/IkYIoBSNeyoEThwkCJ+208iprKDP9jlpgtpIWS4pW
y42EbFuKVAhVQZBj4Nd8a2MG0iCdA5J+ftLKfwb2flqX5yBpeXQi6FA6HsuKsXn4
jq83Fg0MC3P/KnbSCHhLRJwwPAjGzbjBLUBU0mXjR7jp5vUb2YM4P6S2XX9Cz01U
sUF/Xr9TsDjOElmerCy1BlUIGIErMQxvM1Lt4+m5yJX50o+hlOopDdL52C7mcyoX
tbVSCz7Z/RATXoNzuSfICD0iam7r5y70Mfl1PljKszDk/wR6Ua9l8y7UUAMuatv1
PHltYkD9iSeTxc2lLRjJgLHt5zXtlbmWfqAAsMU7UFeSfdqUvOfOhI0pKBzonwcA
xcx6bS1JDCcBGsVUXMRPLSMWYIaHFPso4unSTtSMOdbucOZRNrxt/z6gsNUHcBs5
4vhMktiCWJEFIEELvZPFHJvObG4a+bnnyuBQii3wVLH42EqHtRtiXheJB2ycB3UV
J3JvX/+IkPXa0J6wJrNtDK5su1PSZ8LvtNE9xY6TGKXnxJwALXvjhAuHollGuBUx
xF3r7lT+ihq9kkklb2TMJYsgBvw6SZ+gvteBrioocIplIBjzLA3g5yZB+LmnnjxT
gq2V61EQJ8/t6i3F/QXMzmT9VR08wegOXbUl7sKkaFyFYN3dq1smjB457vX5GwIn
mZXrGNXjXq/a5dPaYy9UNhQvKO++kRGmUc7dR9vtxnFnrUaz6ibYr1HU1Sz+BFZD
8ymtg+B1I7am7PY0Bk1jdWNfxgPl88o2xPfVSapyIReQbrqbXztNjpLkxP1Czz3J
p36qvthGQ6XpEP/uJDmUaDr7lkj5baB4hHrxIYvXu1rNsIKI+IJdKyAdOJzRxJQb
S4Zypx+6ueJtk6F6H4I1NubmQZyCL7mzTl8whrHBgDTap5XkS2ztBgakG3JNZpei
G3tw7egTt+WQQn7GdAtyvfYfQw98u5SERflkGz7qfsmb3OU+CqEqurypXVeF7sNa
d09zJyBb4oSV8ObNP1K1v9+VpA7XONWGH+5a+Bi25UiQJgrsQ8OIKWzbXzjS54vR
+xYDdyaJuT6I3Rrlg8wlhLM1OE5rva8++htq6VgO/DdfsL8NA2JIXRua1q8uAB8e
i2vltG7vSrYv0AISDOE/ND6BDrhzefCpqnnU2VmAedGhwrkIGAx9ylWRrHNXNlRT
dFJw447PaVo0llIBm0W2SBvuiiGgGeuQ66M7dYFVkVViQ/LdAh1NX6KhpGKo7nit
B2aLteNMAcfWnmYDUjlAbgozml/xWFnXr1PSgvmxImt8dSRm3pv1Io0hIAu/p836
OuPrFcQbpMQNHOlGUVYp/kAlXusacJ2TsFfaHL0kQUR55TTbr1KEQLeaRtuahC0/
SAd24VYkCWD2LCrJ+rgGoJzqYxiIvQlQ20xmeXACK88qRFtFqZciWVg7CxX6jVZg
bzYb0e27qrY+YWT/wxieTlNs3vuo3Y3ce5eaRNioGw8qODt0jz2BZsptvjXU2Ksd
egMxth/eidER5EyjPREIP7wQ4QQwkXDTLAsOzZMOjT2FxpuQK562/vbcnzdMwu4M
0wR16pS6Z1uIqHzj1s8//rB4DKP8e0UkT+LjU6Hf3Fd4wXWGgoi0n4qDEMtOzraZ
qneQydNf+zZO3l5dF3szcio2BhfzXtUMNqdH395ltCLWVI93dTDLJ7xGqEB5dTku
Pd5FE4FZ47DwB5BQgYtto248IcQxJKrvnlmTwGn5OJ2NE7dJnp9fp7NmLXv6zzit
leVpJQyXHRJWE6W182b+WFdxNlxIWI/WAE3RNUhMl4PE52Uhua4N8uaUVsHUUFjb
HZLBWIy5UmrRo/BVx5tQAfA2S53tu0GlUqRIUYq9XJvfXtD5GvVMzwFpUgvbbZ3V
QJxcWAPwp3s+bz/pMj/sHoMbuVEJF9FoCD3xs+DOLEtmv8Oo2mYSDTxO1SJnkyGf
AN5KZ8a2p+KEMBknzOehjH95VdaVlqDJanUaXlYvWTCoqCp2Pwgw/VMQaxG1Qt8f
MGOEnfu6QPXFlnfdpq3kkyeCaFsqSfbyI6fRRCRAXF66kuzfwQYGvypGcTYtlUvq
K5R3msyXVfJFH/HYuiP0tICR32Z4pCL9pVObwXBY1hB3EuCdfKFLrHx66zoyOvhX
r08K58HI+/b9uVwOwwyVg8QWmGsuzmzQkArPMsqJNYT1x3YCH71QN9MEeQB3eK5g
ga4X2QTa6g3087lg59RORFJpbE0IZWBhEcYj+6bfG1gchc2LPHliw6J5453SZb4w
lLzwt/yzvY/pdJVj5ykXdEnUwA96NQmesaxhN97yuNqS3eEgwSu6XpgKwv7nL5bw
KEDM++RAudmBqMaz7AHGWYJvbzmYdMtl1vBoz8b16QG5E0J93pAh2qevGeAKRwsl
7Ex3TGC6P5xS/Qy4oEGPxXJTtbTdIrmTsoVBBewXEk+enux1oLPOQ781GWmShjEm
4eoS2hUvvFN0X7DXIn/XuqJhlMd7J8DzACNZ88YzqDUgUTJCmCmc2LWZuc48SkrR
fdD4VvIPxES29GijHKmUci9M5F9SmiDCU1QYjpAgip49JT9tBOUUO9Ick80LbAh6
R5X2V1fMhMuLPKH0+Qqrorh/OU7tkte2ZJm9DTplur+HJiYmvFn95Wyxth17F+7H
vNsGW09ktLY6Bsnj0PuhKoMcDBOqz5sFYD4v84zDCXGFG9zyOI05EYW0/x9iDbXj
IHGkr8d94oHP/huitJPvES6pbtButqKawPXih6K8bZVv6HKOi9sCrYIBcB2aN6Op
Neq6kmr+D3E7erGsXcFc/cOWkguuGnkKveevW+q3AGTDezj/bpkwreH1DrdEvgJI
o+6VN3OGPh4mrArqUNtKGU6cOJvokCUkF6x4pXWG1KrOoUSnysLJe2d8qjjV2O0W
pyZS3AZ1Fu35VSXIaj+0fBYEt5l2KViIb2JBeJG7qwTkOF9BUNLd+LsVb+Nf/Mtn
vCChNLepvGh76he4iNb9OvreKNxEGMTkk6C3wHjRSvx0SXEiEwcDOMRnMCqydPIt
ECLTEI0w8RmbrLkvUMxy6ZCzWImFV0eMcX4PPPUw3EfH0irN9qJBktQ6v3Iys/69
cWv7BRjtTKBvw51Dy7ms8fi6XOWffhxbSGoVhLAppTYW30nmfBrGCn8nj21xCbyg
DVhgpucZ836OWAd19o47+Nf+eRDQ4kctSSadyH0qdQA/FcBK6pH1Hgilc2eRr4Xk
mW7U0hpwC0eXcblt1sjgE2wCWAMS8Ibpd9bp6px4uIt8LVSGfYfLTyr+L/C1g+z4
1rIMo1660TIh+q7p2vMzKMt4rqUa6LW2m7bcqiKpQDRB5CYogCwnTd5PCwBOeFeO
nG69vTOdQmEEFH4Q7Gxy4VEnE2yNWHlG/cCyK2yZ/wqLxzVxG5vAeRJdMvV89S6I
p/XMpDFG1bJZ9DtErQGfbUQSqJ2rphDOdM0DZT0xUTX7VqqcCjfYQ6tOtEVjnC3W
xpPTT3TOhvd5wAcjO2e53YHUs0fUWjLQys9/7PJ6Qf6ceTj66jUkkA0WGOb/N5WG
AvwgpFvlnToI2TF0YauJ4GHeuSfDlMZUDMlcTbuzy7F1JolGs1UB4nhHJzu3aBf+
leOeoUEajpKbP4tcdYRDRy4bmuSh6MnZUmCsUQWKnJs9kmCFZciwMFqKAadw4ptl
MZZ3kIUxYbnZXBTa9tARY8so7Z4m7mVVzTyxN8ZqEn2HIP60lYc3IDrCndqeRbzX
Ko7B1AqLAJhFgulScU7SEdO6tlsQMomIFDnxBmrb7Mjmags4/j+zIMN70ztQyf19
jMAFIzaywWNpxFqd6E1HYK1Z7l/zV72n6ETa6jsaHIgpi0mrFtR9e9nOKIlVQjYv
CwXjk5+1e5mLdEgOBljwlGIQPxtAz5zKCYspxMLFHqlfqiOgOnSuqOD2hJrhEGNw
1rwTWwgBh7ZiBXLcxXc/R1u5Bfv6fNhVBt/j89FTRK2kxEoEyCC0tMidwYJHdYR5
xhY+N+j2TVgwBE0KbADqYtfJpkpWd5jlRWcNh6Q3txWvJH0/ecbnyYuJazT24FUT
PlzJFQIuPcRB2tQlAAglfL0GrOkPsbtSgKSDuPNZBvBaD6YHrCMMhpl/71/DZS2X
Bi7cbY38PKn7m7TbumHjQmAj5MN+wfAJ0Qc4o4wbIB5SzfAjFNasLk/41M6fLJ+T
PnRm2/6oTUgb0wOacUVn7GxYtuexPUNQcXHv+/5mcu4U5fY4Vnd0tHvZzAX7thAO
xLDN7d3soIITZmoNwHjfB87wofGfMEErC8QvmSjzy67ED4Zb+pXRb9GOu/lm9AdU
Zia4vfcjN/G8mfgXtFAAlhrsLFTu9OL0q3E+rfF0bRnOzOui3Ib+8W1GDBsK88sD
L2ZeSptlH7tozce0fWAFCpwWdpip04saz77MnBeboRxReon5PleOmcbM4amfboZY
E5jTh2TqZeIebmZcVdi6llpaw6wJqh7riDyU8UvFKkxRwl89zD4a1imj07D79ZeE
7DhgN5XfzN/GtyqEUYzkCuMQbopVE+CdZXZ2r8JtRq74fQhn+fKaQC0xHf2cF+bs
o15tJ63GNzHBom2FK1C014kelw2YzTBjD0nLL3/eIB6Sa/vqHBKISEkEwcfxF4vO
xKAkk4Ml+lpn33r/tF13YQ8rOskXFL7omG6gayfpABcUd7JSpi+EqN/5WdTrV0pB
Nk1XuQw6KAK9B7gQnYml3CrBF8dYI7siiXCtQxrBs9GAhq3Gfawi/01BPQVQ83J+
YEdyeGD7ucPoBAmS0npNOlKVkqUg2M6SL2T1ws49IxjljmTuDl8VI8ydzHgk1C7r
hF3hcwWYKl+b77lb6XVFpgpA/yGbSa7nxv2EEaSfYO3SoNmDb3J5+w1Es78zeAWC
RjX1Ege1yJhX6XGe1DgGXvrqPbr/ww4OaEBoUG6sHJrWhKZmivhjGy7PtSk+Ifh3
f9OsIKjMpkw5OHtpr/riscSXvWVqCCRwidHR3TGBqTex/Fp5gV8Z9kX6o40tDSbR
hgQ+ALEe3sxNUAdWMVs5Ng/S9EN2W0Ei6FoAQ5iFecTTomYbu3raBu1T4uU2i6lR
TZlNH/8PmtWc4S5Au+Tx2fBGDgpBEpF74OOz0doHedV9utLTUh1qu6t38CoMR7mo
XOFy3mh0VzMmgWbeIEsFJsYwuViJgVtfBE1Y42ipwiPZbSt+p9c/qBW+seYfBhID
pMui/gmjh0cl2UjTCEn0kW3d9gPTjJ8Ie00mTzzqibgbKJItJ5rnC+fBD3+Uxk6d
C093GsATAZBxOa0L/FJHI6Et1lM3yL8Vd8h1ieSq66+OMH0s8s8h+jt2va3+5isk
R1LeYczuuLtBUxGO9dZKUvHm9IiP2jhbWeVHoczHbsmrgnPevS752/KirMXo1B2c
H9BiNEGQi/xQOxpXU9k8q5CBQ6sPX1KnlYIEHwzhNylCAQ35mP9qhPP/71fAYPL9
YuSa69oUlPK3BCRNlQkKbyV+ZhHPbfuJFa6f9VdRjULUxoaYq1n+nRyqD+fUHLC7
jJry2ALiFpoHfp1heuzuF9eQi0HaAFhPI+4+1jZNpeyVtOS+nFZjz9wwX95KjME1
gRTbqOde8R3/WeOalpdMFBmYVfn1lZieTjKetml8rGehBeyhpA24osAcFGERzreI
fO19u5B0wQTQYsjAa4m99g/F5PpjM6cinr/Y1UBYcoF04tYPmsRwJ/M2StF7YxJz
riaS8gB2O+9JMf3CoLhEXXAgs/OkQJpoG6U3uh526Rn5rTrFFBnH0DXM13OZ52oW
uA2YI+vYqB+vSmg1C2wqftgMhydgJktUPvunQzXccMMlxc4WmKS+ngmbeXia7iyT
AmUSyLi2DovDFYCdPVOc9BlrIF5WNDIOiGWDMwB9SNE61SwH+6zB0FUn0g+pOY+w
UUSLvUTNyXD3UNVZn2xIV7Pdalicrp5P0GhLts5vzBBhorjZzxyMPsy7RridNg11
8XRLoGGqGruO7t36CVFgdqDWeEJqsuoVj1OHdis5788PbhrwYGwFmHeNFF6zV7Id
WF/a0Xi/eRQRjrA1kkvH9z2JD3HD8zYLCMUfSQ7dzt44rDUyPIp9AbpZX0fIufdu
oTCYunmVdYJsmuw/2kMUgzXvqiYt7UhuKjMeIw6HUiAYknPZp1dJ8d3s9FR/Llet
p5iyKP/OOUMdrZmeRSbM25TfafDuFoRsmuFBScJNN2JL2ODwNsSleVMf3ybWB7PI
1wwzMR0Wcqrtphh/BkTecMkvYGzM8WYiGgoJ0/pyrh9y4p9auFuTZ3b0wCecMl6r
xUbGNxFcTcGImpzMa1NWJv59kOWg5N3SPxizIBXB7Nnms1OWKNbTqR0UZrkc6Jiv
3B8ROE421afwgNvin6pcFNVYtloz6eZs/S9X2A1PQGmKNHSRAJRHvOmNG/ML5nv6
e2+D0w1zJGt+xHi9WfjI17J1FPo+XYVjt9mXTUQp/bbVU5Xt3COrGJT9w+EFCxFZ
yawCMU61pXzmKE7XvB0njj67Z5f3ZY4LcRKSAqHmQ5W0T6KeQ92JAX77RfOdE+fF
JvZHy5+rebrz5/NMVgPl+4LBIo6YvQmHxE9TfihOaiQAy3lBKEsML4B0VYoryF2W
jYQY/zpJh0CLq1haSNsNjJBwockXIScfUidJf2ntRnQoqZNcpRKvEHJHC7M72l7b
StQy/Vl63AhyPhZGCJsaxqHNBCB/JP8ztTza7mdA34gosWgWhNE9btyT7brnEjfN
5Qp0/ReCZsG0szJ/+Z7M8ETlfi2Yp0/PMgwqNLUd/aC6SAIoxL6AtyawSaI0tbOR
NNTGwCOSWs7fzYhmTIg+leT9hes5m5hm7uDYnuPYinITV6mCjoxhLZpiQtc8lxLo
PGzw01OEgt5u4pqp2/LvcEDCFpT2FXRojpi/C7BiCumAxfxuGJIc0JfzZrqyhL3L
3pH2WkLD0GppB+/vHDHKVbqZK61xWgMBRXE9cGP+6qxNbo+BDS152IlRwLwc+D/C
eGIc4b/aq7rJhwqLvw2rWPxHr0UHmkfbkwa2fsyapp3tS3toh2KJa38wXHxDdDvB
NTbOofVvz9JNuOEJpZ14+E72HKKL0+Kh8VS+tbl8/uuqsBaN4KKrRnwhwO5wmbuz
2vBsqckHUyZ9/5kxaIhAFET0GKgZB4aYIU1hjbw94IfYDblcucdPlVd7V/LtCxby
2Bkm5F/wp+M8vtWqOh6Za/FWBMUyXaUtTx7H/MWNDIou3JKuFNEoArrbCR7cbKpc
wkYunr7cxvx3avGJFAcpr+JqnKIg5SmdmCfaIzBniiNOLNUsXEkeUxpITQYiQ0I8
HFrMSeoNXfw3KxSEZiEI+i509J4PBSyhr0ghwrslqihJin/u0+1oM0eiqfPQzbOO
D98PrZ333tXvFW3HIj2w6Ng1KA/GA/P7G3PclpvJCygye3ed5vyHdrCEtkYazkk1
8iw5VDqnCCKxUGaNq+HoSUcp3cG1ELPWgEQPDsj8Sy4lKWxd2cQhadlvvjgKdI5V
Gj0OSepzaNpG/4UfQJfTR8kgtwaFCKE01zW5kkzpi+lzUi3LfKwV4ykKOof0on95
YojBxRBzCHcnNrF6eHWSSUY0HcWEgfS3pl0Jba4WoHxyVPcigk21Mlv6aFJ7Uus4
hdL+88W8NTcsVf5Of6xm/lnXDiLNKuF8vB/1LSg1s0xMyVmRovYh6sKa1iYnZ6N8
KZKkN3ozWVmKcNIylMaorPPqpTmoeStB7F/hUG47yEuBr8C/K84K8WSt929Vd0TS
Oy06H3jmosLqE4tzguu3bu2e8Yk1one41Bq9lj4TOGVuC6G/GSt6mcPeA+rPInjs
lwRFKs8G9Ua8bFOhFS5BHSwk9qVdtEQOUuxLIUkNEpE3yZh5GfTAxbEwfqNI1MxH
iG297p8qNdIG+8s2qBMtk7Ktzu1v6d37+0rfUU89T8vB5omT1k6iT7t4B4SGsLjR
/p+mYDomVxVesFVUVN4uuqEvNB7n/pwUG+PjnPsLD26w7V5kh56Fr/hxjMT7pJ4b
phdLTuDARhMviqTUfifYkohlTRgbOw1viyPfaLMkwO+qMmWsm6rJEkWRTd/uaj5V
wqYo/HXGR9QCsqjT3QSDuXkwvmkjR30GBzdoku4A0pbUbHvY/7vXffpG6o99QTDe
RKHtNE8H0ibgXaojSSkDwJsX4zGJ8az08WSGPLJWL/RDCV8nEqnUoDIUc8M0FsQf
nsbXDOd/Dl86oJl2d/Y8Br03Lr4hX9gb+WC8+sX+lhtbILUOST+hjDaltQjmTUls
4nU2GZ7n7sJV3LVxFj/oV6CbjQjbI0nJ9SHXea9BQe3EGb6QGk1ooGcMKg6CJ0gC
GWxg0qrlvM+PTI/MixY6I1OQaAmvnvVh/jqhXp3OnG5oVkXgieQTrQw8mKeWay6F
VTViCpxWnHgB6KxRMftlR4aqh1JXUyHnCKc3vpjRpBiD0ZG+JL6CEYt/0/KfyDh9
mHEQId3HeJ3mAg/SdVhiYXTHCFi8xqMFe5hIfiezv+B1h3HLYZHgyMrU4aVeGBrk
a8psJ/DQrQnNyutTwSgbNl8smh52zVonUYN6piE+Mf1vO/VqM4LfTgQfurH5pXs5
4BbCYXsodAvMeycmYF0xjz/faLMmal/TH8qMRIY31rMPpGvxpwEyhNAGbn2G8I9W
L8DfMvoQveNqs3yOWjKXzeSRdW7dhJo4pFTk7/KYRuvGtwGKzrTrW/CV04YbSprh
kpZCGxqETB7VxAk0uS1Yehpe1Tg2qet87gwU2F/+vNU1RhidTavQVC26Qx+9X+KS
qW5Fqyj4sJxnfWT4MSgqL1YrXlOV5OhEnEDUsypns+SRtWCjp/cN4GSDk1KS1e85
LAHJ/xK9W9gydT0O3cEqSeKg8xlbSCxeLjXTR7Bw631jMSDtXkIGKootIJQGnK+V
ZicJVCBvjrfEWB9Bv6ilY4xuxBGV0+Vz70RZrKEz1ldBi4+6ctbwGG+HYIFTBcl8
6AEptZ9OiaIztuJL4nzdQ3ogKfsUQAKWmQWxZZu0B+jJpqhsl74MzD33MTdB9GfA
z2cy8xfXCUmXsFkY9y7yPqSma10QTUHZK8NQKu/CwEVqiDzRmzFYw51Qxa8eSGJ/
lHnVExeuDaVvVO+G3wqQXiaGLXrKaWKe/LVe7yiT2fFlwTTt+7hoa13AaC/IuWXs
ojekJXfg58gMAzQ8c7uer3dM380HqdlOSqWX9Xu/0unWGQMIY5TrRM1HqTb70oD5
P37rFyRzvTFYd0b4KbVIuYa/qyry/o6Zmg6YnhgfWFCMWM84B+wlg4GAThHa+QaP
OM071kysa39oryfs5lzBe97k1cKC87ZFLhxyRg53e7xWfgVJARlly21sOQ+pGgY6
ZUdRa20MDrVCxdvcaaTRNOMiw8y4SFMbtt1SdLopS0kpGWlCWyvfEjRaD/Ge1+Yd
ropXoP8Ut0tYHGnPs6fph0GkDj50ORfjtPNr8r6sSG/oxjMo2pumqDXRwtfThD1d
dYqraYjIg8DXEEintbuUVef8m02QP7P2v83f7uVVBil5PH3KPg23IhPbnTehdRmT
JFRymG5SJoTO6/dnadKhIfEvFJyqmD31Q0u2vQnXxKPU5lX5E9rPopUB3pZLR4AR
FNrbSgEkML7Y+9viZwCxnHxrv15JHhjBnEziHph2PtEZev8XNUKx5wS2ufxTr/2Z
oH7oyNWh0KDdx7xupyJz25Cd98H4HeojZXq7ysSo4hwRuadprwSv+JxYjnbzZK3V
Snb0ABx9IPW4VwA3y0jHIpB/o15tMSqLTv5QC9L8qfV5McY48AJM173F3+HoSlBi
1OxmUN5dgC0BXFa2VU+gGVPlWDIAkzyZt4r1+rRSUbgNO5w0ALFDRX5c7Xxigqgo
I7L6shAJqEMxkk7FzsmgmvAtj5UmKV0aAz1zUiH1BNwr06RB2MJ0xvN3Re395hxE
svBfzMANiJRe34TjZuFKm5d3bpC3s6aSxpnw5uiMcrjOvJAUzMVe3V8KxXSGY99V
r9r/TH4yrKnTAuAiwi6KiLlYNDZVZHOz2Y0IvzOe9t4PBEQv9gnK5wvbO080H/ng
x3OOqV8wHVTMs/+j033OtqoFgt7Xrkz/Vd6gGd7qRAGogNz1hYDU+2sS5RZnV8lP
W9Y9Eq/zHvT0fuBnr4As7r94i38dH6mOeEhnr+N9swgfxrbSSm0uiwDtnrUZEoJN
LkPzoXEtUyiXQ86Btf/tVXoYwjn8eaZdPZTbhZqvuDAgQrSoSlzFtlyUrq+ChMSu
k6dZTWR7kCFw6NR++RzJ7+sF/Ck1HbELrswq7TWjEBoD/o1NPt20yK31V8hb5R8P
BRcXVZ/M8g/87u0AkTv61oSqfM008EwxucD30NuBgnayNceSyYi9gXeHMeI/wLBe
tKbNQHLnv6ZlHWuZcoUeNSJH8512durho2Qg+6syxBod0eSXBcpCpbvqgrz+SMmM
Tcs5f/GLFwcdTiB1yJ9aobsmUj+Qp7gk4zClBhrEo8M4JW8SaMLXf95Y69s3xO31
YAZ8r7lEs04zw6Ae4q2n/qy2/n5ZZiYHyg86uu88/s+E9Kd5WDF9kzdRNiynak7e
xqdSsHLHyX9cGQ74u/SJrz9BL5YcyLdXaBsZUl0DipGH4UKAcCbGtEuuzDRHYXfh
K7L5J1/Aavf3FLN352KljXzjRBVhIyE5L7FAoQbrU+GsLafIXdtLuEtCCrJLrMzP
BDXJ4e38TT/TXhAF8SUPoMh0TlTDtuK0kURMybK51Vd8PxnbOtwgmVCZ6PHDieKO
Oi09owhJf1LY6OGDAgS5aZWZfJzJD+Dr2DEz/jx6nxoILIfckJtQYvKigqXaGdxf
TjwFIaivykIll//NntJi/hu8nC2e1mnk1aof+bgcdlwQ5xomTTO9/2VJIwsKeX1D
xdRxzOJsNVE30CTMTBHvEsHk/ZZ79xCf+/aALsocboYZ6jp7zLkK2i6WWFUo4Idn
VZGX9Sj9l3iGoVjyrfx5RdPgZ3a0IECugdZRZruWsP7cwMzfslE09XFzS1WN2bLM
ZC5yNwhoRsuYPyVaCD0MBWSjcMDtgnESTZEVRducK9fwHZvOwetax+DtsiYyYSC6
jvBkGQbzCLP77SCqTRC74JyAdpgFRPHGu+DvRdZuPALE0VC+y8pGifbv4nLUhdz2
1Pgg0H4e38wZgAV49yNTI9U3/jH/OK9eozYbY0NDkULaT2Sjo5SwtUhMgX8bmASx
+sn31mb494o5DSMI4bzYsKP9+Of341uczF5dTUxzehX70A4hkKFJgBn9Tibib6PC
TaW0lEmM4AqUhnSjufsdYov4/LgFTUkgZxChhIWlyzvi4mz8TsY9HT91B27r7KCg
03KraFZ56CxMxbPJUhOCqFSy3ccXqz+bzl+UTFiX1Xo2NNrszaD1Xt3RYGmb3Xxs
OTxK041MOI4nkKvEtX7Dp//1E6XQ7CWZJEkkD7yBG/1wGJCE5BMi9DPYzGX+HISX
VG3DcXOAwNyCIMpM6TvDNSXJVz/qptJM43pNctiknxjepnPppp4uhWdnpWrt/YhM
TWlFUAb5RrnBk4aQ5ITGwuSWs02eypLBZ0BGBeFfNI5n6nbkwbWL5BTXkxQpf9DF
y6z0XPbV1HFcUUWXyQbmv/YULMMfxF5eOfH8Eyt/92B2x5bbu22QNtrGpZAgX2Du
6NRtuwc3sBuCXb1/Isn23freS3xaapC7n/WmTONfHQdwmw3Mv2I5r+Iw2YC8T5QP
lQoKtwe0tGECzOXYvubA1ot3PPGkwQYa/j98ni0wXkmj6hYnurwHUs3WT5QyYosb
M4wdjAwo8M3WR1IgOURfhmLMNCvUkVQXE95BEOZauSA6tN7jdw0cDUDn7mmOmAdv
BcK9sfjwmtnGoJq9Eym0o5asZV622zSo/kH0lE9HjndmpCgMDm7KBVcxyjp1uuja
rFXDbCwV3jNqL3e0lQ7CPJw7+yes6DKfz4cTElPAj88KgyhJmQcLB6Bg/qxPn858
EP6xBPv1w4NFmQxwne1kzSds54OhXaDeyXxQQAbRzIID6veXvIVehBfbX9ofGwe3
XRhKslRN0ouNQkLFJx5ChaiY3BQxjwzYKyjVvJaTEgUat71EA1VMYHR+v7yTXU95
8/3h6bbluMfB/e9lD8evnJxzk7veOlvRliBnbE+VCwe1YjDBUPkhQTaOnlztjMlM
MvHj6WF4QRcPAyAnm0YRRdGVEyjVorARBCYSvZTnNWI/GG/HLcAzchQ3cDlwEI48
bzCTd9YMaS6GavDr2xl1u8OomHPtaQRzt4VloKUy5rTG/c7bK/Uq7uxpL3C6GHfs
YjkZVLl/iQxCLjLiKatWQvqKS2Rwt9XDrHL46OMhGmUzJOvusEm5LYB5N1rnC7yV
hRDsL5VXDXanNjcVRed6Wgs7VJZeIrmQ3iULDKR00hqpKY/wpAy8t2UK/PC1RXh0
Kc4S7elYf8aCGY/djp5NDcXagfTYR5Cmlq2o4dtA/sid/qrPrh/2UixO0oyLQjSx
9kyzSKR2aX9bJFaAVjVMxpwruKNaYBEB4ZteoD/FXEb5Kesop5xyBaY/uyhNPBW4
XtHugwlA8lAyy171j7f0yofo4vDNGcxGj+dw2wUkAVWpRkK336tbS9Gb2Jy0Qev7
VecECtgiqWKdWZ5Ymtd90zQAVYG7j2qqYY0FbxuWp2jBdLFHdvDD/KvQKvtg2aZk
LIp6GH3vm6+CYC8C2JgsyzNllS2MtAcjR0AwRhzKFKoThrgDOOE5+NUFu7z4L2m/
YBcohHc9a7zlWf0cityHx/h8qwGNZ2s0Lz9y3r9cVRoUqgxxWx3xKHt6zWRQiDSX
d7RLfXPA2UpCd6WB4RA6NU8fqJIkBEgAhv2rHDZI1y+chMv8fnvo1KJpGpMP0MzF
lCd4oh0GJiCj0jQKnqfVESooPuLHZZjSk4XZ7Cbr8NKoPW+o40ceIayS7CXSyqS0
Uq/KPAgj7aHZw0SN53wGBcUOSYMxOQRjDYPIphhsS778eaPb4CRYndZ7ae+RAQC+
v6bmmppvvVWG46nZZ+CaBZvRCjWWUeEM5ApA/6N3vE523KLrL3PfsdgR5zOhXq1T
p0m3oSvhl0TitbpE7g9ZgXymNwyHqdh/8CvkM2CX6lrwB0gDZRBwOED6/ZH7+aTT
PK/xkR1gcgnH3Rt8/w7pelBqgwRgaPaWZglbZerl+k4IKz3UMExQ7Q9jF7k5H8P/
hM94UXw5xJMHoSyqXzDvTx+nhgENMC1lHuIXxsVogo7kzTMMaVvuzLEkLznNLwpG
ARfDaF92/9LH8WWBbIcxHbiKWaKdRvtKbj4EB7YePbgwCtNQlpHJhEr8Rk8ctCfb
sUaJKYejjHF6oO+cRAmI4FQPJ404rgJO1hmU3ZKJXaZL+kof661nD9vhiFf8yt2h
GQAW0I5VOwTTYZaB8TAN5mqtxJEMAaqUhZKcqfolg2sr5tRIUftmX/2BIT/eQPZp
fVsu+TFLQ3Wo+8RRcrtdujmzXUq+wC3vdp4mss98lKvObpNMk2+f0ZsU79+0+Yuz
Jq6cc7lqyiL2DRYwSJ64E4k76+NKmGGCgDqZD02R2roZpfTIzzroXXbRw2Lzss3i
acS4kMTaDH09JCF/WmQQVciGragd76jSbVDrvSaVbaDsgRiiHkAbTIYoIaacvjAc
95iMChisS0UqdwzfbIaIfKmm5tMBWMxUGtwGKHtYg5UFKWzM/IjXx0vqx6/k+ZhD
Qvw7cYF/h1sdIeq2Xr6LAsnr6LTaxn7G0QYKmxx6gXOOvClodpqvjKf/5CWu5mq2
CJgaAjbp+T4yi2UMZEBioRGGdmqQIsHUWLa1r6CwFuB+BAHmkEy1cE5DOmqdhuQ/
2iuZv+31Qy0I02uCWr7h60QgLBrPcShUkuBRDctb85ZlV3J/IhCp8gV3J40XKWBV
qvrKlqfr8MNK/upMekvtlAGOdDGDPal7uERaHdh+eImTE6ANOAxSiYAglHoLWg4w
ZLFBsykYfbsLecRHpLxzbI2eHWq1P4WFC2jkWwk6zoeMKigBkFubFEQGK2Ij5aQ1
BqidobmQjPD7UXMAnGrvHwuC1IeF1GaG7F0MTvwpc+JUxB/tDrTUaGsV+icNCWF7
bL3gO1jsPDuYpUgUT0tpnWBrROcjUIzV96dNkREi9SHM6hcg7fb3XAJidnzkTgZc
LNkTw8SC+c1xxz+lsHMh998F9CTKBYddUi8tb+TE5/kr4cRcC3SDwzqHKDKQEobd
VEhJIukVKCUmYpdYnH73jNjm+I4uFNjlAnQUjbSBAL4Ux2Zs1VxqQxtXMaS8tvaM
StT8Ny2aBSmypH1CgbWvuZDtJdElvdjTJqMKPRrX0A0VqwIwUR8rCc+Cd2URKPDH
q+xNkaA6k1KeZcFT31gHI9jJJBfmOwFcQWn4q7IUhz4rEhuf03yUPGGqM955CCOF
yxEyjGrihEhP3kiiq06WNt1O/NodUehTr5eQ4JC/0GU9HCbvHIYzMHHTCRHGXy9E
HJT/fTrVTbCAoKet1c2VGULc9QOxYHN4fAHygGshH4I37/JdvTySofmLPtK6DtsZ
H0kXcZGD6us7wfXBZJd3cOPNTH/P3u+7ddemrXID5sWrxi/fgkqDRKWNjhBw9SLB
pTfyWxV+l+KUQ9ZQHDfVP7ChkEmN/QBRGPsyPSAq7A4G+dpzYaYv3vqoeqPAv1FT
kXa8lp4IuwCieV8Egm/K15IAQNTuWxKmBtsglW24B44aMLRox1U5I8jBvR7dM/Ep
sFfBzr8I5wDgEaIHnPdV0eaMDr6LO7p6bcq2P7wq4ADdOVF47gTi9ivmQMbD/a6M
bv1w0a/CZ9YdIWryabQFjrlRGKhJnq98dqwdUOMFsM1whOLVasMDclnHjoeMBWkn
FPcDKc4sKmUwgQO7FkuJZDThsNW96FFpCPlYZ2lMaX7yEMqEr6mZtXmhqW7Ygf9g
btpyI/OYUmN3hP0P+86qISuSZ4tfzXCgXWWgsobd9Xq9lK0Nrbh9I6RcYdO+Jq40
9btB/GOtqZcmdmOYi77OevfDiuXWiyXBmvl5+1NvQ4dy2gCGpEEDQmzQ9tNfig1q
8hgpQpr2iwxxNam2CJqr6kKd6utPtQpajGI4L9yGah8idU3pgp+ldfzCwEmAy3Fx
gBxXOGSvhKm2Eb2jepo6NluoKHUUPTRKjpOvks1WEU9s4c1K6crAq37NuwQdHhco
ZOi5NLBGuA35GXAx3jbgm0h71+8Zq8bFfZUjK/r/SyRXTx6XX2GlZuR99mbmVfKO
AyqAKBqWJr1xEihsCxUoX0EF7RHA6twzCW/BW1br9cWgupz7oLTbkV9XkB4cOCYk
7OP4X4MKmQhTqPLZM8LaIHBsYR78wOHNBPyr9aTU2d/xqJJXIXcjHMqHL6Eo/5Wk
U310R218+bvF28VTI9EGO/9MBzr2aJ4ABJQogJrw7PQjsHdPGiynW+1QI1CGo6cY
Ionsgwb9fVCH8oEgWzb6nuKgQcQgMrNk9rAjewp0MH0lnFOXZYzg0+teuy2wpZzz
ln3Yg3B8TM7vzS69JQmJb/pterBjF7uu8n3yKFAPQWeSpjhPaJLTmXfWFuazpdV/
SGjEJcXfm+C8UjEyfY/1E31e4/rguuQM8BTlRwwa6SoTRBIgKgpC5THupDg8y7X7
/6Lzx5OfnIuZf+b8zFy0yR8BvCM1K8hzwtZrs5GwV0B/wWeNuXv2W3TDdAPXXD1q
kZfCQ7sHLQs9rBkgLVGUAIDUA/Sgqkjl81VsoxsKFu3OXDbyoz3O1e8cEf2G7xvJ
pZjKvphJwJ6ml7GxAitJU8RQc1sKUs/nBDsRTa67SkliX3bV4B/kmtFIinQSyiba
6w97mo6SGrGHedYLPOMtuRMHB/WdJpH4osB2RQb08wVtooJKm8l+LHt4YAjkJA8c
Ci/34prXK2sjauxy0401K55/jPZJI/vgPJTHLTkZOdpD7qCDsrkwRCaip1wPQKu2
tyn1fVLBJLHlSTbPM+6X+AtMSaZdny2TWvxf3mLJPAQUPEfinx/4ibjIKh67a7UO
MsKmsYtxJtFoHCV5qfOuf6Odx0Qzc90W4qbBt060P7khI69S7qOjAwzQNXOHYhnT
cRHnEKDllSAsTeTqbfFwqqYizj0D+l1GDPyNLh866nZHUbMPJGJgpsvTaPpOiUCZ
S7eoVjodCNTNnJ60Bfc+100moSM0GmKeuIIDTd4aaZXS3A7GlcI/47HZ01Ug3rK8
kCmYAoRSe5dwDqq0igEO2JbmTlfmZY2xewbJSIhhtM1gZE3b9Vmk9WlU4eNCtvLV
T5L+MzooeEqFWGMaMnu5yJrT8rSRbTpX4/G0GRt2jWpkJuDMKpogDanUeOhJD9g2
wfW3D3N/2QkO9a9C6W8pJvFw8XChTbaig2cExl+gL8e0i2KI1nKiPLEt6H0RSA6x
uLjS8ACM4Q8Ef3KzxnHyPcfW0gVTKpJEOlzwOI2T7WIPRf40T4w+G9HhaQdKNgKy
kqBYy5YY/sy08RfHlS8qRfd9Ob0YWjXlqlXX7PBCFEVuBdLNixU3eeS9eIZ6ldJ2
PwWsqEwgWzqEt1SftRUQLE91DoWUvnorxX9sqIHBCoj6MOYCDyX/MWG9PDu5IXHy
hD66QbbHxOU7aFsyMhFZ4s9AicDTcbl/FAswgAjHdEryI4kITCLbDlZCpb1HHv2z
CSTkQxkEjH3DORadMJjZH7JniWEGfbKlEfRSWMYBnw/iQgJCa3U2HirReVlewqAh
RGf6G3Wl4nx4UXr/FyopGUsB3eke4aa5aEpVF4RT18jYg6ElZcaad+Av3H7f11Qt
IlknAPkSYkLlcxjKDikYR0lNUmHcGEYz8W4NRZ0ZHK+Jx70utLGs7ILG8TBlJvKs
HEV3g3favl5EZKy+aolBC7SjPcb/5V0OlJLJ4y2KZkpVoh2zEMbmUvJwlY4UI0sk
xC8LPIt/mHauXFOmNr6wX0vIrYYoIT5sUKKVr0N0OabfLoL2lZw2uoO3AyTsXQuh
FqNVbZsanYy5wD0uP/LtJgEU/4joXLZQBvuCbg4Q7xUhRj4dYbx46GtQOGNjyWb6
BMyMWrqZN9JCL17IMqAeme9ivVAwpbMBZjov3RRgeqild+2Yb9xsm9bVs+dnSAR1
alWulxUwY+QDijACs9hGHPBnNdHuH9UaK1IW0JanWlMfkcyNBLRFX1QCFmN2GTh6
IVlkAAopRYWdqTl0OXjeorrnbyjaNPToB9vRQ2VnZ/22KzQw/gA4hEoRIS+cU+HS
xnHxOS8WKV9pFh7C5QkrGnJvQ3E2T4ToGhPUeeJtsug+fr+r2m13XDmNPtKkLh8X
C64nYCACeBEiDbMST3mYF8+YxJlPaM5UmuUlZYbkE4EGpaln+tDcfnHqGwsBUPXc
muQb+PXAa4BNuDU3WjXEkMNWYylz7XJKLc4swEzdQ61od2Ajtk0SirqEs7KdjuQU
OZmNiLAcDgIxePL6whzqRWguAf2V8jQ+6xd71xWixy57iNYUWQnUZVviEsOP6XPc
PwPcLW6WuQYmElCK4Xz+j9Xfm8xk7uzC5Nn5HSMurS8+wqsP3ReksrZJt7jkIZkP
pVSz0cSOWHD3FX1kojBEL9oUGA4C+lEI7ciTJxZDHVNBHeMhx80ppniH4fNX0b2F
aV+DLE07zQUePGEfJiSDCjCQRKZnZX/ZDUd+dPreMcMRPPaL3PrI1Rkq8PqBJlhH
SFtJq7u/zOpWVBl3EHUofxRqaLmCvW+GgEF18aFAsVihsuIHepnqntpGm1C0ynai
8FXdkc7Z0QMWYoY8FAhgmY7eyZ7z6FDdUC/HjIdwxHJjBZtt16xnxZKW1En7+Ybr
TrBJZhJWiPngGK5CjzMWaTekiupVM9orTh4bBFulAnblQC//OjDGFG1e2EZhjDlv
XN8EAsd6/SbmXdghSEJIQtVoabjAMdZVvoxAq7I+9aCc4nUYCeX/S/AmTsNNzX7y
AMMg/OycdcS0yZdjpK3c66FLciVY+gVfkfB4S9hUD4lmWurqETqDxYNdXe80RLvd
AL66SnFqUzQVeszAPYHoxaD8KsLdsF17j/MpagBP4kMgWN3vJAaGQ91s2xe7FEW/
AOHz1i3x6Om25axv9VW3KyrwLAWu5VMCefw56ik/62Csxsms5CSVZT/CaR22q+zS
Y5yWY8pmGZJV3Uytb9pVOXWBWqTCyfwA79wDgE9bS/mPWV9XR2d6TSGHQcqGSR2H
G6D1ytLziA+Y9W05ixVi/1T8s0wxM7Gv9tDiRJ14IOvrc2Kxv5d+s4mfoDTvJKvA
7h41N7OOHTsXOlFA9JZPgVH2gnZsAXPgcPTvxTkzxLcugRIAvwfNYCWX+oP1rTMN
PlAtU5UbZ/lVImmDoXRx4MmJU30O/KawFV0KNpcc/hApi7CrJBCTBFuEOl8GF54o
EpsygdIjhb7gotlk9s2sIXuivRyge7n81AZMKfA89YSXV4+eQ+UFvb4VOaLRSyON
Dz71wdR8fNmmurlo+Xko5I6innpZnifWTsdG7RxH0tppnjQTKNW94ZJsF6z5riVJ
ZSe+d2h7/9a+UIAuXvYm/8NZppjNgz+0CRH3eNS8EUtHOKLP8k/gIGj2hAe8vZFL
UgdZAXrYnflWo9LJQ2mpXGtgLWS38IE4V7Pt0PwBZfSAFWyPL5bFena/gSbspfa5
1MZEEAFxhyaOGEPr4hz9lOt4He4HI9cM+A0Q7/deZGY9SL2ZSuhFD2eF8EmY2OXP
blUfl+HanK/nOfMoIFJ+EB28trA6Hs3sth1sFiN0OH/v86MhhdYcm7+cObEq4Xal
Sw9dQ+QsJ9kdjQFNk0rIyIJl7UN2grVLU5Blye+eHp3+WbIJ7mCUkQp0F1m2Bggr
zeOgZsmxRgmfgQh5xX+KCuJ5021NM9HKE1i2a+ICXeYqbxmCu1JRLhtD1ZcsTah6
sbnTF+o3wg9+LQeBA+jAfop9pirZc94m9oj6B2LzvN5Is/9MT9l6tr1RPvQLHEGa
nHgnIJdPCeK35pAdfTQmGBVg0dN0LT8mDQU37SetI4kW3x8uflb9st619o70Jstk
QKPGdixMbdYA1wzqihPg6BUlDR8gY+2RY9klLXO39wfJmozKV+9kesglVWOF8Ab5
+XkWuCnJOF4ju7IV8LbuEhwvKR3VeOOYqQobUPAPp0TU2lG60OwkDvTPKyDPezia
Ayb+xcp/PKDpvGQX2wJwdBt0m+hPw1j44Kfp9cGUQ8oeyTOHl54N6+SVjUBD6SLt
StywNjgQgQQhhaS7I1I5onpITKRwAFAqPBJLz9F05oMHjXCq13mERYLkB4E6KPGX
m2UuxgaRiskMBHamec7EwAWwnOmPMHcoP0TeN6LdaDztp6e8naFyqRC8Z24pM3s9
lqJE1jBolHIuHpAvNaxU//M9gvINjb82x4k0SxbXkkA/XW5N12jwlf76Lt+uoFR8
mYMZoQVRl5LdpGuHeOg4e0Ghp1ZlIFYIa+ee+1RWDcxl2ixGLQv3wkYVQC138Ps8
vsmRLqVnya+4rsDdcRS120hYz7JvyzN8YNUNQUVu59t35/OTl5yRJo52XeY3PIeX
7JJKy6HFbdh3HPQQm4gq7CguAOlkbR0ei7OhP1KRFKjlGt9U6DS1JzQNfLasNn8k
kyGgoIqNON0/ShcmH6ISJXXiSDYCjrX8W/mdGyAgbc854xc5hEJjHQPrvDLRlwIr
RHZayFxpwSX6jttQnPIoPW0F4VPLWq1EQ8v4I8Xq3Hv2In/zyCCGU2ChlKM+c9ll
GRXYtFAPAyp1IE59MMWo5+q3mBsRu/gHiE39zTLpjR4IQj6cN42lyQNFLQKfNdbJ
pNbuucdSHPWV0iM5/xI1W/m9DUKKDKa6JetD/h2pS0AWyfdStpFtch/Kj9n+Vcq7
wD6JGGz2QL59jFzesrj9ZXAnBs90+An3zxPkrL59wc/h15NdE72PaEIcVHqjOq2v
VgZclSYfqXF3EtHD7KAfvhR7LqBcNiYh0zXF+z2Ym5jZ8+7+26Gq+Q+klEyPdaLD
aBAKqYK9o72SR2lXdIDhwALtTJwui/dF2uJVDQdMYiDvcGKeKSn7B448PxqqNS94
0uNgfyICu+JWMQJOwRTO67iwGhOd2aSrID2y29nJzPxzH/bZOcxBNOwfdxeihYcG
JlqCXY6wvLxKVbH+t9KYjjgT+efaOy7RFEkNVSZdOmxjruRvcsgWwXXOrMsmx3t2
ns04T/6m7DR9vwV4NI79W9FCo1cyUoF1AJiPOTnw5AHL5cYR/6txea/XdF9+rEeQ
6lqK+7ZbynyrSkMrPW3JWzm9eQmdZ6jeIn+xhuCl7DvxwZz2eBJi2j+X7wKLSbaH
arwwxxbX+hh4mPGQgDfnXzuPfNyeg0dPSxJVMlNjW88QAHjhEBRf57RpRBUS9I48
32I5zFEEnIhY1H61ASocWUita8vLj9eqJkD3IidOzZ4hs+E9RzCZDJGgqmMpsG+P
+7yIa3Os58jK8CC6TmCXQf2g5zUIxbvIgdIFSy5Pw/II0a5G5YPluDHvK0MWus3M
M+YsRuWqYgsMepQoIwlRL1pr3YV2ZXKD3I/iKVZwqZ4qs5TSFZ3+SctcduypCs+0
/OMSeTwYhWkL10E3cE9yzwfixzLaNozbtY6oogPM8zSuYGwnwBe5+Epqcr0yHqJJ
2+ytbkYGsn145vGwJHialFJcSbnMvV41n9hv8X7SocoD1k+ll59PVhI6LREMTrFz
UerUoIHwSSGsmcvIPQcbE1I5V07sWvaj4jif+TfeRr1+c2jJW1JrbfjFotf1PXDa
WRPMO2Ij4GTy1bo6XPMuKNpvRQc8gntk3Mtjb9sdSXw+MtOoH6C/pb+RMaBRAX1K
e64q7anIboE7Hla9JhwxC6vg9eo7LaWt1pEuMbhrAVBpBwWLccj3cGxI04o+KNZy
6WLnMWWza9VIukTGL3VxUUdPfZlPfCeRisHYvBBqdNCX4S7CsBx3ZtBhRhCeRfvN
/FL/O2qfyxikDhgfY9kEU7e+Qkt4g1yS1IRFB+XF4b8YhCgo/IYTHbWtHDa3zqaR
6bMPhs8+jw6wVrWf00iUuQzqa6+gRM9XxonE97Hjjke3kU+RyzBPqnXkXXZB2k3U
W+Y8oRairnAxFL8usFGAKQiUnYz6REuhqmegIWp6OwklE79T1FZAHAWYZL+8DFCf
8xFXmAzaQnbV0YBtJU0r+Lm4UuiXra17E0j1fSkUiumwhqbhnBNRJdkYSYD76qqx
iveYFmH0iiVP90IT/LvgJKm9AmDtW+vINFu+y+QcirfhBHfByOg7V6LTp4gAjV4k
eMBvCQPbXhtL1fTLdS6/3YH7nH84QJ/7powjS/A+aMXf+z7cbi3tIDe9w0zRAk1l
6OUk0UKeCvp9dB5ZJep4MciaFQLjPZ6G/YZXQHN3DJpLg9FA0PrRdNp3g4snyDP6
0iD9emKztFzGXpT1q+AvkI6crNicj7w7isS+iGEWEj8EMUo7wHP6sW1mk3vKp+GO
qxTYplV7/tGjptXOB6jRAbZ4ckh4TkSbVkR/rG8A+umBZEWmVfAeObnJlDrjYyHS
kLV8ZufnNLalEHh5X0uRED8ILd5jp3vboSwPdFeBOW60s9d2GNgFovkcSuVu+sxL
Q2AKMtbt+f04hVB7BF5npHOWMBz3gs66JJ9xGTEgY8NA6obVu6LqRnl6LXM+biMJ
nJ5kw3sozfm90czvdx/bPvRKqUR6lllHOgblHaZMKqj2c2mXh8OJWNnRXfv/pfTx
saVg1RZ/LTH/HfHdYaN2bL6l6TSuSJ8jEIqiG4ZIt9goShEI4CV86ktKnOqsaqVy
gU6QbXRPVJ4Yd8TYAnEUsEcnP+K2W8OLlkkA0KMlOMCtB3d27k4HTUwCZO+XKw1+
8gy7NiyMecupLWT3IrFSr5UAKY/JMv53jewNrq4e5TC78zNpCbzUJyagoSwnxzUF
LCtzOscbjqBcyL7XYiPRI9ecOLiPzU/xB1fpBdv66khiK8xLCnYbUhvwPm47nooe
n+3XI9w//U5OIYOPX52gK2hhCAOrtQpnRXbBGPXk7wy2g1hlxu+iOFJsf03vlg81
RiDwX0Y2GSSG1FGo1uIY0tcoUh8AyoMGy30GAlYlHf7sY9jz/7Gt+h9zlupnc3bu
QKQt8nnGw55K/s1yU+++Vc6T8rHP3lUldo/x5SMrCt2IY7TcKjlebqO0E8kghkS+
Xw2aUh3rMlI8ti/h2mn9Qss40Yh0yk/MvHGG/NQ9MFMFFjJRQrpWOoVBtwngDIF3
GR5+tcQPfu0dQvoY7nBs2I7arKGuG2iOYG1uWLlnwY5MiRUk6snKFWcjuYWxVOCW
uuNfy0hFc8ZaMoC5RlQip1QkTFqk1s9jc+zEZ6yo+5BDgSxFE8VORFllb8U08TZ5
PwfDvQmUh88v1IXR+f+lcmqKdIQrCzuVhBfaVc3ESzk8Ma7oQ5tjgWhFpyGdo8Bw
Azf7w6YS53YZJgajaukW1VUAV2L6A2Kcb5FgyUa/cwqerpdMTvagfNHHG8I+l3/N
28e+9JfwMYUIQZIP3M49vdbwL5vr1fGEqwnit+4DKDPBePKyl0CJmSpD18ioPsEo
Sq0L6WWZLZgpUVsUP07ZJfPPXA9gouvfJEtMg3Y7qN/oSVVVWYnM8vIGt37r3ZFc
muziKxEwG234PXGsLhHy5T81WqsQtzb53/8U7eFUf+4ui1u62+akxlRVA8B9z0XQ
yOuJ0kv8QljQx1dB0d4KDcCtac/9Bf81On2VhcRxrpn8JngZe9621UaGU2ElrAil
PbpKvk/OPqkR95hx6VKGm0PyCzMHWY+98C/PaogH4d6f9aePHMjA2wUwUTr1j2Vs
DriK4aIr/BOKMAoMQyBAoieBWhIqmxyZpcoha60RPVognXIJ0OHffwhTdMTNrPZD
WKdBTiyq3n+xjQncPHhUNCQPnKSOnOGmZQ97igcHx/x2SMChHH44sEeLTrc/ysFv
0utSg3vn7vgpeBECgsi8G+WwaFokOPcwuVZjzpMlsKpTUMnVuzCJ+rs4cx6/Xo/q
yT0ySZCgfx3jnlnFhbbA07zzf6uYtM1leRzL1p2GkQQbnVqMSdcP2oaRQ17M4FBW
k8G/wmNw/6NYpAhJ/QQQo3HWz4PRT+YNNYIwUKhUkGirVE7l7+XqDNPwgYsGFgUY
DzdYBAWQiZ5zCgvp2AeYLsgKHlE8XLZLRL+5dt0ZcGziWUwOBwzt/NFurdUbXZd1
4MdZ6pjQQZxaSayqTgfmlBQnsGmpqHxX3U0tfByAgn9dj5zrZe35+TCvx9bHrPte
5wqSsygBMipwwLAzQkegPVkIJxi624MPrxbOLk4aMmNgxLOh5V6Qqbd0RDZ8l9lg
NxzJwMASFaKAGnTDUtoZuWbSM3IGHpu6Xs5TzV01u7NZbFG1nBAWaO0ryFAfkx3y
kOUS+2R3Kpa6f2BwTb/za0h0r3Y5FMMHW2MHlZHnk9S0Dfrqdry/bZfx2LgyDmqo
ggu7CIJb2sLOfbQu7LtYK5wwOaRsCYGGAgDy1kakVrDaTzzU4ASnlsPf1yOOsXaL
CPRtEqZW2tzvUY0EZnhJTTKbZp+5YQ7IcFLh0d4m1n6OouztFKTznnn+OaIbH7wl
EsHXUCD/fuvNDWqEZLlPAXaDtZlCvZ/QtiQLay58yY3VeIEKPh/CUkxlre6t2Cd0
/B9eMBrdR2XnYpLUIUhfrgKHUSel8UZ0v2pcYlFE4z7QrqGHWtqmvbkDDBluCp5c
j6h6vf0ljEg8AuzPnUV2VqdsGQsqsucWT72Cuj5vdi+a/JQyIFioI8Ujh4X5pk54
eiI6AmQzs5KOumt6hSv423MaGVhzc5qKDuwHdzx2hzHPTuYwq0c8UuiwSIAxVUtZ
2OMp1Kh8Njbsa/wGc4iZVA0oI7QjysvCypo+M8Yb96M0nXNG1K2Grchv9HOp3nW+
YY1byGD9XWJnKrDVfMi3ADjTCnOiJFRDOsqKHeMN7Mpiuwc/pxE6Pxbylxmfs/b3
+ZUrggC5wYh0uKnS8/qibMvrII24wREz8/x65wjmbARijh7WiNTVgmmo/UdT6MGL
q8Cr2D6xwzQJLzXPmJRBjrx6C/3gbjAxXFoEap4GBsRVhUZL6YczBrhHD8XNkk/u
NXL9VQ3rFpEhaZ5pwlwS6ozF7V8G16JEImh38cprtegg88Jhc9kNsHLDJyOK6G1u
aX9rISi27OXtOXLDTFBk8ojG7rZaUw7OLeusrLGOJ5YIe3m8ZvP/ISSRjcCM1tUM
BOhFy5eqj6LTNbOUAE1ontmPw3XbwokZT7dHK7iQ2vhvRan8QN0c1GFLmms6UjQl
4d8vbSFaa9nbZrOrbGwFW/y5rIl1kNKeBcHKNaBVvkkro3auswmW3kP24M2BEqiD
vpP6R1g3+9JiVoQzADWVL6DPQC4cxPSMt8fgcaJB+RKIDtCh0htmE/IwQYqNux4T
CBLCo8tnZZxe6f5TeadDMwrqa7INPTRYPt5MUjIFvHk0KqEI4gDv2hfHXgoPAVQo
ojrYu4H8h5K2beWClsKZyAiBoFmL7LpgwzNMCq4mEXUYojRkJRAFYw8qsYJDX517
ORpyj+zYUfYfsmYgtVxWwYmhRUE9gzU+Dh+gR4UILh3+p4fxRIyxQI18+UBgDp/1
LcsRr2pAx8h5QSqcAtQgzShs5KG19YXfC3RH7BZx1XnjDfLWL8a5Kq8EqxtDRg7v
EkojHHJHx3JTHPVKDA4ZaXPxaFCDPvNtXWJCY4K5AHZk2pnPMC/wpXkt3Ja8cGPx
3PZUbg5F0N53h3ms8lQOhabBFh0Xt0sQkm/sgCn6jfzghi0O7mFVNi/jzvnLlHn9
WyPCnCSGOvgHitCNVl+ZUdrKVOXENHBqjL0XgUXZw0H8VA+Pxkp8xdS0OrFdhvS4
55Kjz+5PdKB4Q4JvwSXF8qGczaaxmbODXNiZ3Q8V9yOxHcFDj4F1sB8bD/5+eFeH
fNc/4HVoguLpJyTHHU9zBynoxEDa7LQImiNjyrcr0OcHai5iFSxI2qs9phBDPxpV
V1CB/U/fK3CxKMp3KDOR/1coQGLuoq+RCO6ql+t1f9/LW/1ZO+6dC29xYDe88i2p
OimXLDr5Fb19ea0yP7xayaD2BMYmvbjkf/DznvnjtkTCKojzkwN0qSyY8AvE39Ot
bG3OyjW5X6UAlR7d42JAcZS+u/CkijmBg0xXWwc/xprUsoKOlOD27INsrQ3ZUb2z
Ta2ZRGb8nNoqEyLS+Q6zmFDB9FSXg0TQzf6YoaXu6gh9ztl3zbEAMJLwfAWNrbaa
PZ+IGh7oMY5JgOkf9WaDpVemxWP40yjaWWZS6d2gW/baxKNJuZ8Aaf9Hyth8kh1J
O80LTpVtYW+aUUtOfC8vSmnHBS20WYT4hVimi9Y9vTn8M9bd80uSMLI59Hcipfm0
IyyTQIsW/h8JyTJVceNkxy9jKxt7fBFrCDbFEMDFGgPiwAvy8uIoCmYib2C4VJiG
UwTRozCv2e45ZT1xGAEioZ+EHUfwu8ONhlmszkIq1eN7lCURpRZEQkNa4Pj5I2CB
1wmH6N18owBfRtd5DVL+8is2l7rTl8TIAv/SLvDhZLktLG5IuAfuDpP/L4NkOLvg
nfUtteQDCmibl2DUraeFZuYXiR9+0PdmPOI6fsIusUULQ0eJIkLhFw16EAm7VOof
qf6ebiju1BQwUCfkkuNgtRCJkRi+tyzsaYxYPHFJeEU9vKSmN+lPPX3u+oW/3jnC
vb5XRLn0TJjTWOO9tBcgnd5TjCKr7IktDzlNYSGro2eB3Qz4U+3m5uouUWBEqn3d
ve3Baz9kDY5iQpT6JDeGaL/60fswwrrd5Evvg4FhUO5Rta9PDrLHwcfRIh5CJQ4Y
PQGxxIYN9ICOjoZ7bLKHQCOV233PZvm9TzQoS1+HUdbZJO6cleUHsUTBbg3lM2d/
k2RDYmcL8afRucK8pTuvpqYvY74EggL9coYRQtzTk3MEfBz9ZuvN403xHqqrb/eg
z3BFsVmSEpIeGJXpJwhIOKDuHwiLcnax1On+3m3C5XeeoKpBK5iCeFsrtF/q9xvk
tipVnZ7xIVE5BqFTJmBdtqCYoPCxADcQEmjVy/iOggmkXDgOml4Pj6ypFoCbC2Np
Snsv4uzXj/IqZ/mIphFMiPdPHLFwv2Ez/Rz410C7y6hYKW3yzxVypbyFehD0MclK
i5lfk/fi8nrOmKXmFjveRaR18kcushfCbbTO+RvC/mu2kxDJujzY1W/9oJLyREW8
WNQYabFuilZjqgHkkTj/osUsbvaayLXWTuS3fMVQ0XbHP3OxiHGtb6eazYgDAh8l
vZ/HBjZ1wSokiOyt+YKRvK1s6Fl9kKSSuOeXSmhUHVJBsyotdXrlpjsiwcgjogoJ
EwQ5fV7NpqqXTMSC031A8XA+RGpWhuPXqhFtLtWzt4GKn5W9Ocr1GfHHrAnBLFJE
/suThu6aE/sMNfrwwKpLC2369xoQR9XwJmGyXCFDXBsM68atvAxW1sQb0lhWaS+t
2hOXW6CMFQWr2Oh+V3LmbmmBifVVlhrS25xzUr5YLKHkuZJPEGbN4UkUj4ftomPJ
1RkPts7zPU8iwH6GOsJBOlWNhpDFyjhfuTF5NBIZ+U6s6Z1p0nMTjYSoun2LtN4N
3s0m4DqauZ61cGPN3PW/l9tC1Ho1ZBvJvF9/9pOR/BMLh+/52etNzfH+L+SYRmE7
E/pQQ5M8PMCQuDbdf7R9LJ7hcjDOYf37Y+28TtbtEpr2ivSQ9yM9Fdp+bypBUZ7A
8rjbWf0GTOcsy9Xl66lyVZq09XWss9SB9Lo++kCBgC8W6JaJgt4OlKsKkbloDkP1
rkP4Q6EQiDR7hQmWnljOvjQCTS9cTQZnG4DzGiU5cRJVX72SX/gJ7ikfr6wGLu92
LROiiHBDa55uMRyoaiWZdVg4B6HuM2Tpu6wjkYbWCAkbh9Blpm2if5LfLlytKm9a
qzZNRwQ/xKk/pMFk/oFrAR7GJeJiQEh5b+azhFuBYfUzMMh88xcNxQvngQeSs5u5
tqLEbHojGIvPLIAoTYz84YMSYtPTKGGmAShy5j1L2n9p0DGmteb7ExyE/5ScSNvX
ge+mqzEOaxw4zrlszVpKylyNk880pEKmzgpYX+iHmrMcJbJL5nrzsKxYVcaURXtb
ijiS2I3umZktbRk+pw8BrxS6Pm6FzW6V6b1OFQ+6T2ufN92Cvvm+Hq63VPxgKG73
AsJVGbOYzzqW8MR52A5wRsf6xNMFnzraWfC6EBco+Hk83X1O0HUXuV8Dphj78UlV
KNUio01mQhwXAxaVjiXUeE/jf0mjMCSpyOXCYUODZ9As1RuJClQcYdhIzHIwy4Ge
iqE/+f2D2/edlfvczi/Ljqs0trxH/tT9UbSXU/7l4BnhO2ErFAJPBPOKD65eV522
LHom6VTjzI0UMqsuM32jTSTDTYOfX6ESVrAVzc3PmLYJ2R2xMhyu2Mcp2iOGUuTK
YhJ6XsuaEX/uTA7/41bnwd2fUd6Nt1PODH9JswVQSLMq52//feagX7tXG9qWpymf
I1PcCfRR6Y8CXGUFyn2tMFLrpr1r830OD0j2gP0ZFSRO/5tg0MQLXL6mBqqap5TK
7NBlS3IjUPWGEJ4xlaM2gHNmlVWseBZhvbchgUgovPoIiEU1Ozbibegir+LO4dMV
ZUfIX+5yTctaqtMKo0p7ktu9tk0Or0BzZmq01912/zsMWS8phkNAGIli34gG+9bn
YbHQBiRVlMfOMXPRDWiSVdTP/Yubltu3WunypWmDb2xwtdBnGR38ASx3BN5pmaX+
p1rDaf71o/5qf+KhnIRtncCTyhdG09yjGHEq1F9jAUGsZc9FQ3lUfHkxyl1wAdB0
wptT3mKzPgDJFu2Pc7Mnk3HKQ6HkJAGxXf2Rero8pcJNGPYj+hR6o46Ra5usJbzO
Ue8HoTPxK/0AnLgXxsNzQktjlGeN2wqfmmu9xBf71CBzTVpYuuirmzCRI4tTdaqY
B2JphMor7OnLj/zfRtWtpxjyF9n2w5pFLUw8j6jr7en+dlaSy8iqn/T5/qcWC++o
dNTCxa1lDz5OYXFpwKciACzyWgJQJi4i9+ThtO7Y4f32RtnTwKnGSa1VdaadBCfl
3JQ14qBn3N7EOflpF+YN8xUAIxquLuk8mpXrzQxccVyUxoXgWyTPffE9MSiockQ2
0eIrsS950mrHId5Oqi6jgQRq+xdpCDXcFTiT6h/1xLglgL/Xuc+43t1yqla1Fj5K
JpJdMiqcT/HlvpoHeAkpaTfx3mYUfGBEqJinONUT5MaO2zx9o7jcDkTQEZtx//Bc
X15EsLDxfXK4/6Zjt3FohfOzN4VfAy3co4ykEnEql9ZYENCEhUXnA/SU6HS2f0x+
HLEEWFSxxKZF/qE5Vctm7O1vswymv1QQQHeHTK8UK/762CUgbqgeeSSzqbjbBCRH
AdEU5aoxQRJSt/ynCTQdx8IW+nvk+5BFa4feQH90Z7yTDIZKV6dmjUqFLHaurDlP
T59qfrnkAXSMRKGvduTkDBNyv42VZ0RawICLYAgHZJ7clUlqads/A6pim6vnzxmH
ar/MpUz8Vrpr4EJEe4iK7IZXkTLZIoOl/uf7BlyFCPK2eaPh/MoWZKIkn+ItpySI
QNE81BcqS2mOkwHaU2SLv+ibraiv0BQ88y24Dda46moqzmU9mxhq+JV8tlSr+H+q
+RkR71gIyH19lLRgyyyKDBAxSkD2Bqs3EcY/fERszg8suhkAb7CNyxBVNObeRKGU
Ei7I26tTieImfQLkWFyG0hKxX+OMc/C6EbVQhT0UbX8EmljpNR5qrWus2uKLAcig
tS5GVIRkcljx3kG/LTvoEUZ2H6tlyUs0dE0w8qv6yty5AgwhiNfYIDZSm/C3Cku7
I0+BXeIcJRVA9ANmbltClE6JHdZRCJ0IeilizSRCtGMKa9IEXVVpkyZkPDHtMZig
u0kjkg0ga5C9f56XsizwAGIcEXLTMi3pVnsjO/4wmYVcV5DeVMx0tQ/BlCqEXhit
auSMVEtqCJvvptTOjeXcDpMU+vskHNbtwutY/KbSgpTuUKvIQdOf4wLHd+uBAAjO
baIOdPgIDvo+c6zSa8HuZB1ut/NkAuO3pLuosXJ1ktc0VwYQ0wAWif3wst+MFoC5
X/9O4FC8hDe8m/0LVPvgoKQfnIhSTrH2XM7rKzjSLnYbYX4s9BipWk6Pdmjzhmfj
121a374xEbAiERC5a0+94FPIogYpA+gpPLyAAJ4mty2hFl6gvQdrErAOIDZ1Z90J
bGIb+YGR38bsocnfY157aoZddMLjBWoeb932ZK6vQTAj2rQZgKTJC8m8BIWA6Cqe
ie4RhJUN9CSuu8oi5Yrn7uSOzqf8FxGAHLBKhHU1jbDRT0bD6IlV6iqpfz/xHbSd
uYpyDwRYXHthF3YAMCHSvupJQp4qQEkmJP86H0AmytsBMRAkL258bMDB3rOPLT94
jN0QedN2SaFZmiCpNfhpb81EfKt7PvdRQ4PyO14w4y0SMaYOara/EdvvrLFoDXMW
d/oDhr3TjItYnY6B2ahNCjyUyrt+QJTMjhPX3B5mhA5R8scA63EQ6iu5OSIeIYjs
WmCDXZcKNwkoEXnARpCT4UcW3cxCO4XZohbR6oFaiexzcp4yXpT2dvbKckzzRLdC
N5IaKmzJ1TM2RClY1eXMaFdRsdRX8QN7EaQQAZhCOovTZBwB+gviskd8g+INsQoH
Ou9EM3sTzxKzENK9931+R2hepllYc1vtN+eQpS87gLH4lwZc9hzak30b9IAb6qe9
bl1ommvkMB+2cbPGiLbxK4CAye049aVUFvOBnM5Vho8q3gc0pMr5p6KGbRz/Xbne
L4xB8LK396RaI5pMJ+kVmRWm3b7XYcEEmAyWdMBR8sOhu4hBcubGbW1h0VUslwQv
ADaU5zfdav6Rdu3BV2K/tlzbjIelFUDeANyru1R0P1YkHTAjxMI8HHhiw0QPX0Ow
0P6oZDcCR4MYgTcmat1xaLZ6ZDU9at3crt0wN2FHNBRjcUTGD1dGGYJ8cVAA3HVd
Y667pRNHynl6VmdF2ilf9q0pnzM60ldS3mmmD+axkq8y6Ch/BH8SsaVZfXvZYTF+
0JDOvHG7WOKQwrktJ662ZoVK/OuUTVfJxSw/m+uzScbOiJhk1uJ1phXQK/vpkwEP
2VZEfb44Iop8uKyKf7JS9zJg9QOWSXMnu1W2MZILIyF5s/+q6c1Abaz1wRG1AoXS
6PNsM/EfcNwK5OUOZWTsVoLILZ/l9KtQppUG7FtbLH5ZPF4qzUMFJhA9OFImkS/P
Y+ZDpAnKbd5JPGZxAn/50XGEuw6wCnic5nFMfZ/4GPu4c8AyqMmXJWTzr1TEnOl2
3rsG0F3awUhbF/QFWCsRz6zQ0ZVa+YyIDFoSCg0D8PIKNlph7wvMGoFaa6kms2sI
Q1aIVjzzr3sh9Ffn3IET23eZpZUqJCrLQjF3siX9QLsAbrIRtMiN8bHYzCILyFKt
3+4C6pBWY46iUAiUR5HWTva5WnkkUueGDB1je92B1jmTGQxDA3ORLlASLlUp3yoZ
HMLwnovI5yzbxfY8DhUVPZbhlLRHTk3NtHv9betI1rgptuoz31JcEx1UpxeAMJEU
ImJ+qALTn6x03bemc67L5VdWeZTDNrvE3iql0kovkYSRf8Ne6G9VWU+dpsxjR4QX
vqRCroETBW/BS4BdsA+u2KdkPUTIiv9honW2OlocI7aKhRDz5R9uPGjUU0m1Xs4U
AaCLjMQo2eQeomgOMlQ+QZMXWSWpcP+F1cgtbv6YKBNH7pH36CtVg/onbYaIZ2mD
cE/65T5pEpLe1wUAGFRTQawpht81DtlXsBBQ3hskPPh5wpAlrOJaHk1Yw6k4Yi+p
bDU7SvYLwMkf0dGklZq04dTzsRDjOiyzadzImumHKiORb1Xb6Qn3s0YOCQ2KeIkX
BAAK0Gu1goYZzeR589oLyWOuZD4xZ1DliWVZSnXWUK2meX6eDLwetVEamaE7HvKG
YeMhYZBc26I4rysrAsgYxQ0gHawP25nGvaWTUhwpJMOj0cfX6dXGMyUq9RRLULXC
QOkHNrJCca2puvHaHFAGMONaQegKZjBjVeTArOu8Q1z9Nt4Df6Zu1sO2X25j3DF2
pyML8hLs7czTDJmZqNxUJgl4ODG9aAzTfY6tqnH2nN0/BXHdasClp9kinHBcCy7T
LXMFMQW2ggI5QtMhNk31sGwiYVYwmninQMHJ/5Mf4Xry2RxpR8xG+axTkDFDRzm4
T2oWu4sLHhI4m6QEX/7jF+Hg6euVLFA+SedWzzk1rxa1sVI/Bx4D96CAWNfBYrex
Smz/77asZtZfYJ4izgbRBFKmWzZ7wvJj4Y5AcsIYcovPtr/MXzSPVTt8AqbF3jAJ
GSahXhmkbEcznQvScDdyeSS7i1bQ/ASKuKAW9h2EQZYoJ8TbakmAOV+z9+onGdVY
s1I29KQaN3S+yYMIqfePnh1fNh7DJfYIKp1508sn/fHl53X/1mI+i6J48ZEZtvoY
k0xfpCRa73gkRcHi2FSmt3dLtRKz5A42UyH5zA4Z+at3qCPyfO0lL/ivac/ykCpL
dJpZeJlE+uqSBQIJQtqIQoidGmw0OMUJKyLyEmg3fznrlybcUECHo2tJu3rYwqwV
gRJFA3hayFFFvR3QXF8utoPbrmb+D1N+Q3r8n/PVzo6Qxhz4PhZv2BJBjNgjlwdU
/8k/HDAg0+9H9FAPmh5frqG7K0WS1xxRy0bFWJwjrxad0dMhfUFZuCyZDJxVFEnF
77+bqPuL3cMrhJ5nNYoKSDkqjIEJ/WuRTPjQFqRPdGy8mCPHxSyaXGnTRWvQcWrg
sOYitvH/CfIvbdAIY+hQ9v1xf9sn9Ayl6Zq+XsDZlJr3ufycr3beqcD0DUH5m8Jp
R/8KDBuhHhqbrKlREAmSPyrbhQRgbjnbSwAZUamqHdzDaujavaD1uUQMQA93byPF
PWpKBvL44iDuZkkKZYxEro1W/Qgc+YYJXTAYG5XeeClNbQYXoVXLddHGpWasV+ni
SYb34F9Ci3a/R+iJE3KegFaVZFC744KtN4GcZDC6Q4ovxtQAObctvHcZDy7N/FRl
JWIPFUnjDgJ6CAxb3i7lB0YCyun7gk6vd+YQR9hQvv3dqQkgEgj9E+0Qy8f8yGzq
3HvovKcXwpUjB624tMoVbimAyvUZCZmGAbdeA8pmvVVCpN7B0a6xNFitzvgY+7re
KJaBc5l8qGj0Xg+aF0XkGdPtB8HX0fveaWVYCiR+01fyWTSmBr7IPgNtiltwRjSP
fmjO3IAvMqCHrh1UAXOlbgDSuWo8NfLLDVTUEPAUO7d9EeRbtk6uRcEJueO1GCYB
turtgMgwEoOknSGulppliktBLj5b090bJ8+HkWSesvr5F0euQmzPqDTkLiBEmopC
qtmwamnnIJGC/bapnb6yS/IJpdr+4LUXjfmzSQmzvWhjb03ww4pioIioVUG0tWwO
STUjExIx4S9wpGu1fW7pF4QAYwwZcABKhpJ/1WRjM1Vgg176PNLnzXgPzjwyWxoa
YuIyt0EWGTiZJqVQok5Jno2IBFfsHAFBNXftrIdo/Pe7m6RVhgHTJDCVFZXNuAyP
or7YT73/6FD61GcIJ5pAbgEqQ0IcUfjHJecMzgN4uI/l+QUdBeYGtmvSCfDuD53U
K4WgbXjtND1udPYiKyFDEnyyZGFRoODyjZwp4EuxiXunr3atQoRJa9ZLCPYtLGfX
1ez826FP1pKne61pfNQHnhfzTfKlrACTNl0fhfTkuXH2MTe+CECaGe5VhLiqFesd
58zqn6DBKyqkYeCYazD7W7JJdf2vjlJjZi/L9xTfA1MJv7aB8r1/0PX+RIoau3Mq
7Jh06G5gg6BVJrzSminjCbvzg/DGPISuPk7Pqb+DBgcfdVhtEsWx2N2h2BhEDgap
l0fTYRXjufgs1uC1qaavbCS8D58SJ6cg1ktqM1I73uxL/IOCZgZHgF7VH0kFWKox
9kL0ColgVvRbQ9DAxi/Vsx4xM0WPYk+aHnRk6MqqUTum4gx1xQ3s0brzULSy/ute
I6FXBePMDMy+2x93VQgmljsyG7FuGIezsiy/Ys2UGh2IV7ERZmkMDeES38v/ycyJ
7+2sGfMd7//jgX4lSG8dUOiEM/PYSNljLjBE6U2nmEHqzwXHfb5PdN7d2oNE8DO+
uSVYhNx/B59uUUhuE9QXAA1AEI0bU9oZF/Wa+dCFcLoy60Ul9RfHmrSc5bYOQ91t
Me4VjF4Eo2IscEZnziwVP6o7qEzDfykwufkN36P5cWCYQR1Rkm2ES4QdRhd3/Nhl
YGlySOcry6w4r+yC9Liaqzi3idmMzBIH10yfxGC6DtLVpESslgFWkw8Lmb/atGiX
5ZzvZLUTKUx7E9/3MkXX2rhSBWtc5Oexj2wjJWLsmOsbPqkxm6V/JRCdI2uMygIJ
SPjTv+6+pAybSBEfWdWGR7smRxXzfkbVjeumocti/i3hfxslqDcJLlpOgjCibdic
cchP+2QXfh/ge9vl/l3wcKOHrclUhezVwV8yJstSZVDHqVbOwa0CLlTawI0p3rU+
7vfKoZocCwC8mmDg1ais60On7cHfvB1ZVzuwVUC9zKCoYyY/iy1EvjUMiy+Y44b9
cZF4R1J6RiEdj6akyTyZLBlxDKXbBiLh8WV3kRXrIkc5vIVwtpoWnLEJa1iOz+ar
bCr5GaehSgkYZ7pTl95jqP94zHD1RaRcrYJXx1fBnBQKK84n0fI4hjVzaDGhnBfO
kyS7V0sGRPdNn70AvRzfqjZ85i29nhVpE2D0y8k7AZeDT5jWeV+uRTaF1hD7GSk+
+wXn+LmtXQnCSwAjH/5EuydqF7JkXbxnk9DhgcjJw3Hv2wgjMokmsn2HHE50RYX5
UekGXkruk3TGHLH1vB1mtDQ6saCk/T0Uk26fSui1L6qeVirPvYrWmgAPVQ44jzXq
an8B+X2cZQ7+TPgzMdy7m+P41RnwwFw+obKpwU25cvk8lsFNYNFwHGJeqmVoXYkQ
VHnT3AYd0ATDAGqdOfis6E43RKMXX8IcOL3LJIOpt/niRbPhvNKmf2lXlQDYsy7b
djivQyJqe/Ii8H9qJJc7zQbWwt/tx26GoI0BVv7IhBzrZT1Me/qEH+D/+wsHmKSe
RTQm8JhPtRQ43e6OGIW8HZ9I22kqgRE+qSiEJjHbQTnHNmbl7SK8UO5KSiMTZ1rK
MRukFbToNA7yWPPCIenWjhVoKKq7/thnoY5CEgmFCNblDIxrJGnkRb/wG3RLbH14
ZTvzviXqRjwCmptL633v+vblS1jPqmId0ISzb+3JG78GC315Aq0TNYa9er3p12qc
z+sLFojAY+1163CwZeona91oWHYC74Zk1mF5GIrtW4CutQrIm3UxA5L7a+8i4FT6
QhDge9p9wg3KK4rju/phOrmMb8a/zPuLZ1Vcxlv80KUbbJW/J1UbC9kuexVREfDO
FMZOfut5WaKn0RncPErjxuuc8R4GqkPYo065sgioNHm45gm7GkRa5cGQkHXdT7MS
AcYHqLHwFKboFrU3mNEwLPJO4ddfos5PehaYLa4dKOp20Q3vygZNAhWXpbpbbOhV
7LReipwAo2JlWVCCSvvQzGhvaQ/BW8H9El85YpNmM/E/iLLT60pQFk7m8YASS5G8
RfzcTGKnGcq+1WQsFRFJRtHs4smq0K0OITBhP+EDqRSwgkmoBMt+Iesod8mPKGIb
fCMZ5DIMUgPIuQ9EfVRmAZqXxsIDKFkr9xiHJClrdd68ugfm+XtlPBAKhMURoWAi
l8TQkGByh/MHWkxnnO+W2t/25BOZYZdXp2ytNLoVKH20Dh0g9A0igDayxBa1hDAW
QoWM0m7V/giti/q8fTWs23vdqpEgyYdWp/efu6PXP6oU7EBGv+hqoeSD25fEz0N3
qAaHi68kfLDcNd2zsRHf3F7OQbvfcuhumsfuIG4PiN4WpL+YTXJd0LzrDFU1iU4q
FC5o+2O5YkATNp/gjTTi0G/A9zlZBuA11oHriVYrMzq4ng1SQFMijdZtRZoiT9LN
mARhjkyz7cIqHhvkBJvYIifv1Xamxs98ICswCHAJH9Zzo1ByRtsvNCwFtXFxVUh9
2SM9XxXuuam2p5Z4NuAMb0W1HIcVuimwJAN2kYWb/rk3mAOezCQdVgkKaAWEhkH4
TX/6rrE8LplBwJ2incCQnQocUui9UVKp49RSs6TQhoQwNQa8uuBzFQ+dRJm0tVkl
SMpmPd0zQBopbnxkN/B8CdrWFnAOQ8xPwsRNnRFkQ+MSHB4c/W38gtZgMyS/f7hT
4mqA3rjaMNtFZOfJkeL4v5GEMyZLq6vjdjnWA95W65chBjP2c3J+SrTV6SudcXIG
iTsKpOWvCxvTETrWnio+E4RFVFecQjfL2U1zr8BaewhnEWCrplJe1G146UKELIP7
WkSrOGjACjXoZ9FMFkq4U/e5iSvGe/58x4UstaAN5LLgUwKbz49Ziy4FsYFyGRQk
9a9N3RsC91xW+WELdUwxopcLZ0vxeoLkfSbW+XxgZHliDjPkPd8eKVCNx48oYnRJ
qXzgYe/G4OnKXeVQ/TBi0TqH57y/9EEhFsRrrygGyhwfDYHNZAD/T9KHhr17X2py
3dTlWcr5sOFDA2/RQAwk0/m02p++Kc2BGYu4kASDVxSflPQdhmkd0OXg688Gvftp
zHX5Ym2sqRy9yMg9WZsTAVA6uCSbyLRFFol+WDTSjTWCM3NOUtFPDfmi1N6I7hHq
TtlNgQswFEDnD1w9Qpw3ArhwPtGVCv9F+Igrsq6lEcsX5zE8RNn7Q2YSHkd4xgbM
VjlX6ElYnYBorkzhoVUnMhQ4exAXuDIGlBdx8r4P3tQHc3f/MJ8U1FayBMcl3M27
TC180j60F4Eat+WmXXsIY7QE+JOyoR2uHOocTSVstZ+pNj9TZdMgejJBLilSCNHG
0P96iQ6JXvdTts4hM4hdX82xzAKlyxtQxGBbPevID/ZX04/f7CWq3jk/9kzgGRe/
5Tx30V9dkcoahMQJ+DdeVHCBNcyzeJUDMeVRQUrLKTjoWXA/8MdZ2uA8cL9T3uB7
PSZEgBJ2oj9/NNBCW5F9ny/+ZjQGFK5cDrNxQ+NMuVylaOIVjnt3mIeuSjHJ8W+T
M0wZn+k27PM7BbA0AqA0jh3CVdt+3xWdVjHaPwePX0ivmFq2Yw6HjRbBgaUqU4p1
85tDlwkp96lVXGnWPlP1iOBKd/dOFAKfELv4QiYkHiBNvXzX0TN748dvUFMwz2Ct
SGBW9EeEKj6TfYJtRGlFY2r+RTMi/EAtXmOUbQCsRyi/kcOg098n9EMPk6QSRgfd
EqCo9r0ZWBf8kA1gWED9H0Q18oeR1X/B2inXzEd0eBr/R6849+QYDpvBHHeCI0xv
RW0i3YMCK5AjpJCybIvnt37OefHrjslCftn5WKTzWFIy6dGSkieDTTYOTZR+cqzI
m/e/Dv+9IzpwBRb+h8UjLAmous+BYis1YIgtqQZyTdW5/ph6XImn8MlBGbhnjJxt
CRFbe9E2PEUBbIfqI7y8xKqTDER/i/JkD9RouSDR0J9ksrCejXV6qBFpMUUxzA6L
K7C4WmLE8bp9riGw3QeJl6HdezMEWeAQfqT5eSHK8EFqMLdPTfQnOhMolcnFndzm
7npjCVoGw40gV5d04kQkoZZoDPXYlZOgJUVonOd+g3AQiAml3LR67UdWzelI8z58
ygvRPPOYMnO2iIoyAqrtXzVhxEfHVQdIX0EpuQ1JqtXSr57EbPRA6IOZ3oPPCr+f
awfpHfcPWbtmVbv6pircLJ05nVaD1MO1Ih4kmGGtXIOfYWbwxIAuTdDRqlRx7NxC
RuqsT3m2fpqzjCwoYrYlsE462phyXRF1c2WpvLXHjDIbn8q1KU8NhGoAhtOxVvIR
tH2KeWvVXt9TV4Rcy0XqEpx5/ARp3/W5BGde6KzmGNOt72w8sBi6ekQth4Ju9cVu
l8aQu+1ObpSs5uZk1859mDPxVR/KtVnfzteLYcvfftu62POMRRT/sjdd6gNlueQq
e5mhwF+VCONHprpB+4x3duF8gjY6AW4uRlcmK6M1u0/uHHic7gFj3w94EIUXPull
93ykeYCUwhwK/a76LNDzqURb4GyN6u6orYq0l4dMszqQ2GM4FH+3kSRWsjMSmXtd
bK3Pv/Ic2rAuxZoiCDxHxIyCePdnLF3nE3/m/9jOHVP7ij/5qr8aDQbNPc/dUynp
smw1s7Sc6mVTemQYErkfXsNH5Lgr9jVRpuZ1Yr1y5jQy7xEgF8T5niH1HhwUNNTc
oHoI81PImO0fPPbaLa0ur9v1Rqgjmrxq8BMDZLLll86wGm9mz7bdlplUupxkZZhs
vHTVL/MdhP3cY4xXlcqrKNZtjobhUzEwN6ItLTvXQM7NH33N7AmatA4PeiQ9E+LQ
/NDMwrV98MNzZp/aE2E2GlOukMDJugWCiuCFawSQSolcOsioPu7Ri2rRRV0WSCF1
5O5g+F4atVL8L5zF2dpqoZb0Q1pyUGYygU5YPVCa4Uj6BpdjDuUN9fBjVjIie03r
PETne3JSv3DWq3nRHTfQjpi4EVLujqet6ISbJa+5uvC8xwxVwoE8DgggGEDheN18
/QCorWj9I2mcW8OQSypxnqT7bYF1mfk+oONWqNIQON51Klh0g3QUvQTappqJsrbl
ecHDujKduKFHmoHejINNqH+IpDheCu20QKzwJvvH1tJuU5L+wrg88rhUXt584nyC
Pv95rB50recSNahBAojJ6gBycq2eCLjWSx8X6dga9QlTuZF3oyIFU833dwa85HfJ
bPbuDdM5hLT1Bawjvkp88wGtj3dtvYqaBqwXJ3fsqU2IwUtK+ja/mCydGylZN1oK
a6s5M6A5oxAb2QfcvZwZFNJ9yC2TMdKyvYuAollbYGX/i7CMCy2V3eyZRk9p2uu4
4qJNAZnoPN37fkFxyRBBFQ7xhXfGfVv8sJx6Kt/AYxbyRFIrGnonL5GtjbdmgoFY
93TPTsR/HBjarazYOnReSuKfBTXsDnTxkmSqqbP4CeWWqKkc6AKIW61kzqsRQQK6
wPqlFpwVqMSUwgcY36EdDZBA8oWPo0xVq5D7sPD/4pC3u7qJcBrdGBsC5Bs4TASX
e05H+wkCUvNL3d7xRPLwhn3Cuf5e/ZNb80SsZsvZfFUultdKK6vQF4kdmyxYH5U+
eiAUNJZ3JQLewsl0fvBbvzflOr18jwn1zLu6MOGIDmAeTCWQj2VhtWS8jEOtzPmi
z+F10gwSkQ+HpR1HSZ6wK9l/wndGUzu6F/psacN3FuhLZknWWICW5Uhfcv49QaPi
AFlqM8aGiWF5UiwEmXcO5S1YU6qt0FsUTY2Lfh7+hZcDXMgMPHP9swk6VIfsTtZw
BZrD5U5S/KbBuUJd44bcTdB9DZ/I1ytCnx7sqCehAaNjWw2CYWFgQc99PS1EGNqo
ypeJMNYwkYn+Iw9kZis7YiQANqlKblE1z9iPXBJvnFYUjtoa1GoiD6shsUzMcY9N
ixfsGfreuS4PzItMJ0Y4C9p82LORJoSxI/0qiviPZuHJFGu9cigQFnm2AEZ/rWO3
JcqL8v6SRk1xcbdAS9Ua535kNhLM29gPDk1E1rXNNMOUCyh5bIfDYST4vSA4BUGt
0i0OQEElXiVvH/MadAT/csRek2lW4okAmZeXNY+zlWK0dm4HQ69dfU9Bg4VegOVj
aasSFaonfmGZmlJxuYDM4W6TyfUAc6VHyl/dR4H3yaHY66EvSAX9/yXzRYViBZQX
VCY4WXZ2PiGirLOazd20D8yn8ACdNyd7oUNH8/66ioj9QQ+2EclL6VTid6FA8Ek2
RW+KBAc+6TM40oho9aJXxMEV5Xp8+2Pl+Eq9Fd6VmL1emRWvm//bAe7mbbv4bbzw
P+CwFrnfLfBPAXtRbD0lYJCSvipVurVGRUmFvl5B6R6sYzSOxHik0o6YhJsR7IyM
v9WeYq0EF6A7/33tWquzFpYx95C8qG/CIFdNyLKTPP2de+kMK2lFWXEznbZ6Soc6
lnlYHWdIP59J/bi2MtxlotWW5456U4fag76LC2lQ9V508Dlya/9YgrSfQc5PerXT
SGjU9V4YClbf73oQHeDYIK4HUXpwO3FohSx0Jh+mRwFWaBQgtjkz6oUhB8Qe+f3E
fOTiMkvg3LlECWGMwv/BNEGB5KD+2u93czpXdkao39c1DhPTVPGqaQ5UfwV0b0hU
/MgRrOkV0Cj6hCPEh0MDtWOEvTOcZmZuWbeJgI8qw7V3F9lobkj4PfyUscW5dgb9
5KUBZNhHRUItd8tWTMvDZyggmvtDT+U3Byvtc6jbbVnRYxaCM1WEaIRKgSjisjsC
Uj1NVQNzExWtzwt2ICC4QFBFqyyzHlTJM/3OrjaceFglXRUWKRfxe5hjQ2Fe1TN3
izac7FD6WiML3ZaSJJMExzrbT0veb9Nv/tTN5bvNwbmxZ4/F0ErxGP0smrDGu7Pd
NnXwUCCwRdiLHzHBxgD0fqu9aHF19weggUWONQNOo6Ven13d51Lptwd6mwMytYS6
Mh1vRxhnb8oJ9BP86TWuBFeU4LnGufJbFryhspP98W+EG0/KRhG0x0Y1w+ODjekW
26h73S1cmJ92J7dm57SOM8xd9YucduKSBHn9RyKuKgQ5URIcS3ZqQrhorV1TJeBg
k6AvVEjXmuppcQVWONOzYMmWuzZkzgl2ooCPoFCPW8P5yTUwMV2dYCqr1GIOKUxq
69OWn7nHsP65tnoxQ3oGu3o/tykf/+e8/CZdxRFZVuGWmQEM3WFcLXZmXy4gkOaj
BPNS/r/qAmjadqykrTHCbjQpJAFHt9SQVWk2x4w7gESY2nWaJUxBG/TtHF+0Fjjz
nwdR6ncRjEUfCLSo7izZE66m95nuQeXgD5M+REmbPxl1RIzv/JcpVYPxG+BuxKKy
RsANHZ/eXSbMgNevfFxh6DW3x9bC18/pYEieqlmnaJH1yTG+o+DMERkr/Y6MQV/+
895j8KkAHvIkZJTRDNgCSF7KvjgA4fu/hxrUcaTRJ12CN1/nB69qqCmMG7oZuP7E
Y5djfTRNjUhXdKwj0SLxSBgjOBLsHwD+c/sqTY+zeVOLjfsULi/bOsFql/wUCU7D
tkTurjrYZsq0x75ufKVV3wBzytzVc34zMf/cUeedVfuljB6+7BCgDD1wilNVWQf3
9OQN585vjMEdbIYQFbX4wkpDxyLWQOTR4hlTiyl+xFk2O113bJk/d63yFhvAqHap
JjJL1dNv+6b0517gg4UEnGWG0K5+LJV0X8OVgEPvljGw7FWMY0/35LKtoTTf+vav
dCCCuDEiAXCuAJYxrtcwWkaQJUlBrvXbNhXAm4qRewVMrtQ/k1UFRk751kpcRbwc
1ZEkdTr2KwW0hm7ykmMsPRSgrXPshHeBR4JvgXsTX8eJUPZ7EJK95dzUFUCGFjWT
oBFH+SR39Bsf7iTMxUZXn6sHFm5zgAA+cM/a6F6jidj2WUowiZHLITkMlSn+p0WM
HBPaud1WfPd2QRt06jrFM6W6FX/O2vRziV/PpvQObrOksjSU7U9Gctz+B2v7mPoc
62Jd8JTwHQ0SHMeF5z3IaXKCLMLCtF3J3vKm7mUqwCaFdmX6/BX3BKsum0i3vIsL
MB5WBVtba5MUO0PQr/nR53FljE4jPC4LJEqF6zTJKNjrh3mIlzRKJDAk9H1/Wr3/
sdxWRz0gsSLVdRx208fNk2EVB7y3uedZeVuuHlUAr70nEdEGLRup/9trS9luhnUo
36xdPmRfdVujMkix828ANgsje4vh1hZFXm02O8XfEfuFLc6CJJvHk9Ky35L8K9xj
6WfcX0GcFhkAvC2Xc6o6ViKISIDsNu91WyMFSgr0SdqVaHon9nEKinu3M2oZLo8m
wuQbcyT5jpqulNXrzWqkF6VHC/+7v+zzilsN4DApJLnVCI8697Y27GHXRPsR2gxp
AVNDb6nQos2q9yjpCs9/BRre1n3gLOJ0cvcHUfEJ7tt3POnEJGVLiwCRY8w4wcy7
rPScWXoOfozKVLP2AZ9kozb70hOjsb/6rXnAc4QvokTKh45aKhEH96GaPBvAQk7G
cCxhFYtKpdJozCHBAtCcwy+tjp+UEuJFPA7iAJKn+16JAGXw4uOLaSPaP8HBEUfO
lHVzQ5z2KBGbfMYxggfUJDDGqSZ1jkIsG8LB8rcgemDgc81VUw9WfT9Q1CpSPTc4
UZZhTd1xXCiHltxWM1bPuID6ZPgHU9imT7rdJ+qisorNzBSVFZm9Y1Uy3EfV/TOk
qRAnCfYFig2sXb+EtXdVCFp9IiXIfQLYSGMxikYX/18oC5cB9bHGypBZ4SFgO+ew
2ckOCorh1VNsh/OuWBMisibhKxS9WEgFsPTBeDYQLdg0obfzx30IC5P2XW3mZ2Oo
Yw2n0AnUDrEqIwA9pOQMHnfm50rDWxFdfSYxPhbawT8cUejphu4y2y4Gi3r6MS24
J0tqsQEIBXOnJ8HuKvFeb3ATLIyzBfLbCxlNYNryJdnsWZNDGO9EhpBL4inRl+8Z
oTqaqfB7d8ZID4o/macfxQF9PwiXIaEsoqici4vg2PmlmI3k+XjD/1sM1tPV1vX7
goiuPu3xuM3gwY0Rv5coEOu91VGeGiRXzN/eJh/wTYEO8u5Cglu4H5R9XhUTQXzy
JMcqLZt19L2LgxQDbzm16OjL/T88blKNfQtzmzHps0YKxXyoomUHYMHQESUiND3n
ejZgBINqU7MK6x6j/W9VolTNXXP1Foqdq/0scEWzPaqCNi/WqQ9fG16iVYl3yz46
EUFQmqVS+pr497KOzl/gJ/hfDK5f90rJx2u7z3putCnJJ9ZFslbqO4i5MXDphWE8
lqyOh1tX+E/0ypn2i8GpaioPeHAEXjMpfLr5LhKPumzupjoB+5pHD0PWaIScDEUm
JA1s4STBeEVXf/TFQIuxHMIfh71cThHfuK+u3nnE3SPrCM6VgZjr0zOyk0pmXnFp
N8B9mCIhtta5qHP6XHHD59S3IdcfJRPiGD4Cmj5xnbraP2zy6zcw5dN59Kgr5Kht
AKRRfzibK4bqLhd06GxP/RHu3lW6ZajYAag1bSTM6C/Sgo8eSyyuS4tP2aGuD1ln
J7tX1RVO+7+ke6tucKiEfmdn7BzdfCxAL+xVxaqb9RjAnevorfsNaMA3Yk9Q0JzV
nOtshkjbrVx/yFFYE0dUsbr7X6ksuZik7jgGz9FVQT4oi4a3wCYlmBH3YRnUIEvK
Hy0/LAJiEnoS42e8SpuOF2WcmqRQAwTxO5rBA1veXyZlDW0s/bPgEPKYozjr+E3I
32rq08NEOW+N1syv2MNq0nh8gFLuLUUenR2h2IQLGlSb9iQL8Yu9l6NL4XA6h/rY
Gtr3hsU5c23a3ltt053/J5L5YIwzKnxj0Z3IAnz5erkBwSNgJijadzuD7ZWFQ/fW
ca7y+IKFSlN55kuLWHMEnQKVLksRysz1aCGDJhWZ/EdG8pzuq0b+UrrGiGayAlYM
Pgcg1Qm9GO/pj6M0n6gqs7hGJOuMORSNGBGR3qhXjo50rltCaAgslooLd2ktH307
z6pKw3QWi9bQzBY2HYk6Xxtiw2u5UPC2dsK/jttVeesFv9xjY6JqVMGdp6SlkXNd
Jr8vNqO4ulZF2Btg6pPlXkrys2E67IVhfzJ6DYRc7HFLcdHX+vfbBDPdrIfG8Y+l
YtG5ctEWHwk2uJ4lUH1FD4aQmkwi+bwj4wamdyQRNFikq1vgyjHty6z69qsi6JUu
SD4whovPf7hO6gciH7fRzXosbW0hsuucdQGdv+9Jm0Bb8UHXk7S2xfOyfCjISJh0
u8B+IroDr7ya6MHDyAY+X9vM33gdhdfV2hFFCC3WGBVLkWki5mCY0UWsYtNRLRYN
4ivT79t92q2D80r5tLoe27PllPWo7u+EUYToFaGuk5z2w3E1VbdpKh71YMWAcL9T
u0TWTSRIjdNbpb99zCOXQeyHlDPhHeyehx707lIcPaa69NMwNo1psh3/rbf4a+Pg
EcRxNrGRi30/lHLiRKgG1UdYQeMtSWjuJzaBQt9kEZXOsvlwY+WJ8+fJ1aCgbx6n
nU754WoKvf3GKlBS8OFEOHoPTlCFVEbjDepeEyNEsAocg/oyCssaOt30i9WK7CVb
Y3iVqdizYafbbihipUjwRGFsUZkfdlieZTdVFHXzWoj2cG/yH9gfCy5F5+1KlpcL
VgSIexqUo7DThO8oIc3a6qDo5w6dNhyoELkxcEEnovzeozpkiMnMpgjD+Ke3cKOJ
iKy3GCSO2dxjTazNIgGcZ77SxBaop3jjJ8fK2aUf6zZRycvHw46P0P6yxvYfALGe
NlgNHjad9+RDZRTR4Wu0z0A1u6vwVbxltUBxNOTgkaAAodAo4tRXmeUivpP98ox8
69vkFBlwH7zyyz9HxveRec9Sog8IRbwl3o4nLDqQxJ1mD0V9QpfyHUFSa/Bh3wao
dT5mm65XKkPDglKSe8pP393K1HoJbjxQvxmanLNFl9ZwqXNtA8KMaSGDUVCvIDuw
lPfiHxhxOn6fmFMNjJJ2QxGUAvbqESswcakt+6dfZAvLpt9Y+gxPA1VspAy3pHJt
eRvQ5QPZlCmF76ucaBxGzd5WuUbTpPE4K/V+jN6D8XHgaWGcjQQaRm95B1bYPA4o
6UTi4c0KmtR7dHj8Z4JXCGFYwGEuPDrcPhTpy29tY01Tx0+ufbb9ycy4am1BzR2m
s0nhaJj9XZ0RBOiIFOUXz6W31/Zz2DvFGix5/MLH+G6Sjj5VuGi4NeFX/I0a5ncy
LyCUUoY6cZXX3FWmYij1Mph1579XFSFVz7jLxsCqhZdDh9CXI30sfSGdeF3Rrq2a
aeoPKR5el0DXBTB3BCY4+2gwUjye2iYR4yljL5t/CUDSwjUujljbXGjSb/mneJuC
XSFfLZdHhmUWTRuD6YcOWsCrj/MZ280+6MdhmREeQISJgXkVXvbdqaS4CzCwkisv
LQhq2tP9WRooUjg8Qq0hOGAQDe/r0Bta17jTCX5rnOU+GDuzjiqMJChADeuYwx3w
8i7EicbwZFjOw0I/QSlAdYZ5Fd9RqupnU0UCeij5/cdQXVo+DZgoR8lzVRw8nFn1
G6w8L1fC0DYv403Ub6/R+pvRHUSPGXclls4D2G8UX8Cg6Jk6C15bM58JBmyM+79N
1A4nXgt6XdW8T9KJtcJxXFb4OcnpxifnfJjJSm8q1hHwTXOEq441b3v8uQiiKZdp
fxleMK5uErOxiKWX6uoeSLB0BrVQy8fN3Kl0wr575FlAxZoRjAugmsFn0ZzHY6M+
IN50+t/TdWDWPBIueNEtY8p4l/BeZlCorBQ6IHDVk/z3CFWi9ipnzdECOM3PJ4er
jZcoEXDcnniURBWDbHmdW1Q2wA3UMGV72dKjUizqKh6bIprDXt+F4TdKF3zt+Xk7
06nGXENMgzHYD/y/FScLe/k0OJGWgvEaRp7XjUeilovQtggAFeFbvyCkJnYkrAFQ
xN9uA7hG3mUvuUG41osFz+mBWmXgx/WFoNqISMXQnA+3niEcIiVI2xJ7eYk000rQ
bKDN5svuolVnHul6XyNM1SN1fmPb2PicAeTQneeDuXOro7C6I+wX9MT/tjiazDgr
uw6AG5UIoqtuVqhcXdEKJ1IgALAH9EfG9I3c1f+ER64sqgQ/mMgrZIa4LctPMvhr
KRUk04TdB86MeqLkMlMy0ZEBJSUWTRZ4PPheSlQkDpXy+vIM0Jx+SWALheRLrqpa
Jb6zpsEFl086CVK4vMI5aZNni0eVGC/P0HcChhZAFpVNpnWb3k6HGBaRAS3ReL+B
jUBXqrZfzhkfdMTC9NevBqEyT6guWtJ8/D/lLWSI3baYiaw5eO9qmb9ZTkCA4XBi
5yDO7TPUNG5wr0zkOY71gA5YfFMcxb5xxJXM1j3/GCryzp2TzvkLOX18HOI3j1vy
qkkdKDFGzm4f6Dp1ueixSr8q/aJ+y/nSbQDZR44HdxRbWeZlJg8O+QcyLqn2TNwO
e4G9CrWL7fe4rYJfqzuCYfB9S71qMOq9iqkzG6Nvma6gxVvf274WuAYzb2Su8djp
FO6id3HEHQzen6Q5B1Mqae4NNNbjXiIwmwFoNEV6k0pFGUiHBp+KJMvvh8y2MUk/
0VkqEIxFSFnY16nPFYGVq+WZbbH+Q8OYXIEakHwIBq5mdy1GyHIHXqQOB/yLs3si
8RTkCY5GyeztszpoLFQOuFRaOe2FSFMM5F0QtZnLBaMJH627RgDFdAuELfs/ZRFN
C0+ruRj+8DNfS0TwKGTWn5WT5IJ2Y+0rnHiG6BC7rv3bfEbIFIsUO6W7bpHEqbiV
1GZ0LIUgKw3qXAZ4278uYCEb0+WldBt8ORGE1ib5wZHtAsAxkp7bnOhOwdPrjglX
xYDPW8ZjwgcLKb0HDyGvTRs3P3PFVeKldU/azcPT1b6WqQNNdQLikOrLQtHNI7wq
c+bkPwrkosFH/HBuf/sfzfwt2xr5KQkwdcM1KnLV5DTXzbCWS3+zI6m1BCe5kPv/
sePh1Y7YOgs6+6aCpGvMhbuTZqLH+RvHirtCAjWIzo0l0o52/qcRXm0CAiSTSgHL
KbnkGgHPwaCxz4NQmWMEo1DCMxln0eu7/3D0Gh89XxCrOJciFBfwcvCtmqegSrcX
eO3Z3qdipsySPqLcp6sQwtGMFdBXIdrHRA7PS/kqmQu3dz1UEMKyDpBGDmVkMI83
U8Qp7jGNZMzNZisfwupHcv24D9MAJZ12ACurL66UoQc4NlmSoIqe5LShs8LxWJei
HaA3pXgfYEeAGkMz0QHsShM2ZiwfAOz+112epO/fuKMkGoIJO74ygwLBobMbU927
jfNgMvYBw8XJa7bRfOJJ2zF+lsAWY0ihW+ePozdALTb+OhOAbjSeshzmUKWWQ/J6
EMYFpSpNddmVhRZVNm2TlTmhr8/yBvxs3dh8AX2KsYZnVo/yKCoM0vUNBDI33V5m
s9E5zluWoJvmuYbXZDYCz5YPRxAn4qK4S5UMRufpFPnblr/eymAhylIcVDRQhXAs
7UMT+9X3Frrl9Cgnp2m1zt+puxWYbM4HScaE14y/oeVxyZDVQBNsM1XhOYisgKJ2
mSmhGd8VaejcgB6Vq0ercoMWTI7j7yl385FTEX+71UG073UinBVssODHe/c4TzQ9
UgfsEZDVpFpbBJCmL69k9oFMGd69tbPTng9jp0cv1UoLr2di8hmLbL/LEzkj1nTn
jcaCQtLJ6iEPt0pmCkuGEo1FYwgRhh68WsmWTo34NbQvRTYfA71g9v+4LFldLzzL
i3cQ0YOGSL50Uo3HgURdCYCaPXZ2jvvmzHznNa6Dr4s6Bfo/f0NhocEClVnxJ9zr
/G0EbXEzqUFveWdwv73jn1k5mnQLn7QjbI8O9KXQomIQadKCpKxJR2H9XuzngGRz
9O68yv1wjSr5PHv1ilCSOVFVE7LZ10k6Dq32hDLxYtu0YzaU+PUIX4feBKu+V60E
gMki0koMjVA2NMDKFAj9mty1qzkJN44mmIyLR+kxuoZEGTz7xI36wZ3YDi88+7j7
RBphgQxbI8MsWFBc9o842yAsL0QvuV1uuMJ3XJ+5eR0oZ3kohuX9PGmfDKJ8F3fC
4IecdjLqVpTFLLFFcdQY1COYJAJ55FRci17d9BG/SUHq8ywJ+9mbtUk2nL8/ui17
q31SB5SoeCrpdP4IZrbhwDJEndsKb+561MKp6U4dpuFL/y7ahH5XHvDlsOksYhUt
cyDFYCoadFva+ezLmiK30sf+ANVXqrKn9X2dznWJU8Ii9M52D0ISgh4sZ9Y8ZY58
eiDYt8x8Rh5oQNBPaZ5tUeDlw7PxytgHxMd9B9DZYREiquoSG7+y5CRcOy5b+AxF
J0KWY074JZr+ROW29rZBVoFaaxeFnIh1p7LtTrt/iDwCsQIFdwLdCGsPaF1qYHww
rnm3Bge4SLsU0G/4xBMYQP79hKyvhqT6mWlYTWwU5WFweYeHrg/Hbd94Dwf67PCd
VdMZ34BfydyJ1SToCUvG4h5RKykgaTNX260WVkSPHPHcmS602onJ4zWkO3opyjE5
HFEUk1ozliJK4uXxQwSFilqVmCLxcLwXoFRTPBxtvxaRnMePn4b1DgYbZ+xvORqV
1vSJMc9R6xH7RXvg/AqLa7kv5kRquXiy8MNMsdZsBRgPYiE9l62bosEomOpLSfSb
z+IqMweIuiROGrCR6aR8WWJBWuYrst69YyMVHkuAviNVQ7ajWmw4c7Gomb2FcBRp
g0AOtQiZXaP1tjlvuhVUj5zsb/gi5HDAreYP/9eRElAlbP787mBSCr1ojif2aAkF
yMwCU14AQIJpMrit1k2ZZQ07wZrB3AoYA7NzM1GNg2Vix5ltOpyZzFHtpNtPpbgi
B6KT/L+x3i2BukU6w7j0ZHdUgawylqeOf9PbsYZD54/o9tuDpfkU//TtCTZRxUX+
k1B6qbPxaolSIyXrAACV64iHgty5Aw5plbjTrdoMPmN7A4RATi1LwuActcp21HfC
lqd85iTNSorTZ0GS4Ub/Uhij7zKip73ce35GWOie2xEm4OCSg4qfFk63BSEmwHJn
dMQjRag3F7HGOU4h/QjnJmrkZuDgiKDAbqhJxau4AB2zKtGOlxTAZAPmfnTYWpO+
fnSYbILjWvIh+gloCGnmvX/6LcZ7Szayz/YT8NMvvgdVEmcY+3S8PwSbdkgeakaa
xBJ/z/Gd5H9aVemkRZ4IXphQrpT9p9JoCoj+yNX1uo+by+4GsbOaoJn6+zjc7YUh
wQrOxN3Gjz7aosUbeB7jieR3Rub8Y3cAZxmQhED6IgAH65SS3uR48A7gFsdMwwli
SSwhl9JW9B8rSGTfdMkNp1lnIDg+k5+psn/T50ycS1Q6+zCE4aC2HbjxFLufYVPK
WA5pj12seMdvQVIrNMy2lIVwkq/UStqMl3cWYFj1n11WII2O8+HLJvL6a3gZdjiY
VyV69wUWYFEjdJfz6xl/DKwQY2oCA6NBKY/jyIThB/aQ2BAvsNOu8eLQJXPhNSqc
xMVB74I0+37Uxj3H2QLMvs6U6CnE3kO8LndcmSMQYYb21FmNlZwSKJfHG7hvCTvu
+sR2uf2VLGL5Jsc6CH1bGNeSDWSqlRqxMmKPYC++lVVZdVG1SO1ZYdWg3cISDS2k
X7x+xinxfi+gU418tRbQHPvywNqXlNUcetVmQBNx0qceCL/6zUXaZ60uKZ1BSW8b
1qQ5WUnj8YBm2KaDSLYcCB9bmq4SxrQK/VUdbVLSet6YVT9LDWwyvG36IkAKmpTw
B9lVpmSzPUWNkBb25wGD+6s3nVZF1iD1NHA3J7YJD7hUsFGH9foSoGWJf4En1rxV
BfVcRd+jBCIdN9wVbGfadB8b8EWDThV3axhSTfv/swIjyS3u6zJDjms7h06runZD
4cKj+X8Ky9Q0y/w+QqLU9U/TkdT1Z8lYBW+ZFqFlzDO86zobJm8FzqadyRRFWSKp
yEs+ScR1R9AA1EGz9oBuNgDlStut6GePTKlPNumhLuv0J+t4Df5q8H4YCjKNLrNG
4PyNuyXzav4EvxnkDbXHr9NWKWRuZjXu4oinBLpyfST1fgXpQuBuyjMZin1Z8rIB
UkWCtp+MoeWtrKJujqJ7G0EkroqGZWslSOgvbP1lCdvjc4DayM/JcqqGlzB9Bv+V
Bo6NJQ8IoBfKpWxgP9PAYzbElWHRQYWT3cbe1rulWMbnUj01mRH9Zw9v2tpZ+rD4
z2DusSjjiSujB7JXlsaSROpgpRziJaiOKZ1Dzl7PI9MvXsMXAj2UP2YNs8hJWYct
KOEIBNbO3t2BP9Xm/sdhy+IT10LFFGTLzjalN4LB6nJ9b9i9nG5wxMhEOPvDIyCy
RzHO/fTJpA6gWQKx00Q2iYMBvfH6oECHTQRfyAMOoar5dX9kZF1pzocAQEOcHg8C
p54ib5M2Int9MIYqCCHFp7G96AqiuqbGbSqtplAPWNxlTgfozGqXrWgrySC7V0tT
hn5QgDhS55fQfBdUFp3AfJH8H3MFvwT88xKxdAVVJYTYoKzrAjzSzlSFDzBOhWCw
rNEJfWpLrtYa+nSBQsHB6z06HXq+AwjgJboLnaJHHP+vorIIe9MaFGhuA1wHYw1/
uxgYF6R+nZHHCYHHShFUge0x6iLbdY2zgZHJnET+ces439IJeDp0BJwA71jiOTfL
Rt1tmvsT05Ct445Ydl3ggryC9uImyf2DH2Dlp4NnR5n6Zq10t4fdfe5umy1B1JKp
+xuc9wIdScKocCRDf06sNO5t1SkN2m3rsxMy4P9SRbWiNrMcRLbMQUbvvuqmyHDf
fBkMnEb6y8tacEAvvUhsNP/h/Hwpfxub/wO9IhTdIkABY4vdoafxZ/ARHhiePXWq
igayoGdO0kw6SHn+1awgp3Zasi1Ddq4xdyt5A98IdXejH3LxTkczHJMLYl3yQUSd
cj0LMthrBP5Ow3A5qyBRAwzycO15lomyMe59jvOM6nYwox6UfNcADGlkaOg4O0nE
DzGg3wiMHY9ZDe77xzyJL3TMTx03Lc9ErZmwblR9H6J+MH7JPxr9Maq+8WU6G24T
eorKYPoqtL9aNntG9M4Xlr+XFAI/nzgCdLDZJUTR7k7L12WE+XlOXHa5jqydqJAz
26HLI7/7olwksQHjMTPSZMVwX0yZcKOfR+0Vz1LQrNNri+zrRwGIcsvIYQo62+WN
+ZpjEQZs3tw43mlkugUO6ZT4Z4ZdVr+oFHTkY019NzAojhSUT6llIyyGRiH4FnDp
MJ0qFfU3VLURw93kUw4crr44ZTYbuAgumbReWhkC328v4x5tzh34EtCvUk9mqkjO
+QB5fQSQckyxHDPTwNLczb925JMCcCuXR3LVqzrA3nHweBPKLf74nv2YCufqvi33
xAhOvf9tZt/fkqkHEmfJ0vZXJBKi9xzfI39hEaUyl/A6lFVktkDcY/n12tJpJT17
yzGG8XNtfTlBE2jtTlTYxDe/lHY4BjtolC/bMWbE0AHNRBhnbWXgpKGMhEHvNuC3
zo1XvqYnwzgbx5kx0ZMIjEFFa9t0JtYo8cRfW8P2y45F3oM3EGmk9BqZFtS+s0MY
DaVBeC/Fzm69aSZ7h0dC/O2wUt2tLOLrqpZ6ppg/VHj7sZI+88WpORLj6veqR702
6ELUSPaQPuafyjOYaajnOxp4P7tSguFxCx8xeI1BY23rwkCgqEg1GPCGe3tNazpb
dIXg0Rw5Fl8Pa3HeByQR2zpqUOui8PwgX0KBsmRxeJMDqWzOuKKP/QHCKpeKm51x
v3QBs7DjRD+6fb+3GxoGDsECgQhAMHo2Z0xiRkS/XENc1tod8j21PyAplVoWF8Vi
yP8tRa2Onav+uXYRe7cIzNRVv33GgqEKdpi632nVETgcfDvqaboopNafvco8u5lv
jcjB26RI4EsZSqZV6Y9q2BFFPx3auVk7Hf3g98TX2VUYChNMqsG7d2eOKZwCity1
Liju27BCBt/TatvukWKNtw8IYFhkA+7ux4UaGgdMs8yc9xNgrTgOnO/z+Huh3Ih7
DZD51mip576OjeZvSGBt+A0+yZAqF783O/yFc7bOErLaPuU7MEZR3ud/3Gij9fGb
y6djDdRXzpzNwrUyoPqXEbdzZLZd3XtLHIeuJcqjwwSHe9N4in9A9q57aKIDAjQt
hCQzpH5Soa56bxEGgctlpjRSrWf3UMRu9K2ZnjREZEXJ2jTG+FDylAdQADPdtxp1
xMpsBOtSEN1+SJZiLDlVWNiXBCfknWKTmZGbppThbM3UxpqQTs6oqIPBFN6X5rdi
XglNcK+SDjqjumOqjMyQzX0vZV3T7/mo8HsZxhHegOkB063T+3WEXTGEYH/OrDej
nEoakmZsf1pn2uJp6abZRPJTzetcdmA54PaVnw4rsjrWdYvuwV5jMsRXnmCYbA/b
7apzAwFcR/TYdGgB1Wm6ArdoOUbOtapXqQ/tyyjQbUNw+08vvNStYsi1fXliMMdF
8Xt3ljBD9jLcs1GUxPOmew3ffsf19P1UHu/CbK4mKM3mgdZI7LPfApGkbLfatdoz
gaKw/zqTeK1q4AgFTI8kFBZtFz5sGjIZ4i3LagO0Crwa/XUHXdYwmjP7ffs8eBzW
/y8IVDanAXY3shyHXSaCQlUJbQmDutYNACx5EkhhpcTXeWj8diQVUBCsh2l/5xuX
0ke3UlnweW+FTRX/S5n3IYIfrPufhmq0jELRwn5ceK+dEksTXm/XaoxrOaIoPKvU
QrxflXCVlX66l6CzT5QokEQ4unobtSmVrqMdX1t16zBKWo77QxWw3FFQLN7hLIyq
ztYotPLNf0QAMr8hCP4dzsZltWARfByR+ibXV5hNx+6rj3s6R1haaonlOOAoDjv7
WzXRjAZqWBU2Ecc4HVRew0UMFIYs3AjQFxRpvdUFuXxIigyENDSlWwyNcKbT5tc/
NtOQYW7LG3IvIJj8XF7fd8sc+AiigqU0ycWmZSqj+1dULnMACkTPH7WjoquBkXil
EbXmhfmH6ZhSEACb0tcJ1OVvKUeHCj8IhBMrhfNO7XTAkHxJMD/hNaWzMzPay3Qe
78wYHMKW/43bjNpPS9k6ciqYtzvHPstUMV9C+U9/cdWmLH+cqW9jX2veYXx+tUH6
Y2xkuuckyQivYFeVDAZqC6jEKWHVkDCIR+KTl1NFkBRoShBabdsNjFJXGSvJjoj+
ot6YlYcYcfMpwcR817xsDSCx2cfAc6tllgqAYLYuueahK31/y8dnoDNbGudUVLXk
iNh5mH1ynr9zM6boRG7oMJgm+0HOtCGdiTs1b3qkiDTE442nZByPPPilAv25iRRC
GfWg+Egx2zjXxCKJq0+3XwulIPa97BEJ9EviKvHfPJQ4/MXPfzLC6/r1LZyozJZa
56M4ixWiIV7J5E7WmPbUFj6VQsyhjjTiMQF+dc2B1OPikxzu7BdeeCmE0euxORNJ
7josQDgRhwBDodscsY2N0AMoz15VYmvJYdCVWMs8zQMdbVXecAb3Q1eNb2uSGy3F
3QP47uCQcNNpRi0GXySNs/qo+MIWi5Vj6rKLYH+/zrPxqHxFqUEFsvusyiqNEJwe
Eyv+sTywzxNGIFzeRMcE2JsoQeTP545DNzxh5FJ9ruuU3N30+LEXN/KFJsb+onhC
Q+Lx9XY5orDHQ6+/yo2K/an5GAk0mVjkSHf7DA/X0bx/BTsVNZib7RbSWe+hMb9/
QZz/6ivqZmYwO1bVDQi5iJhR5ppchv6Sfa2SUZYFs9DGPB39nKiCEsWgnEqaeMDq
R4zPXrNOO3tcP3VzbAlm7Y6MurZHnPDWcOhMPkgtRzRx5AxGvwKYUwhxJyFHZBVy
We3yWliVxupmr0T2Jf9OIz183iOw4hRuLNq2an4zivOZNbSlcS6Uf/aGqi3XIEBd
6NdM1ki6Fd7xiXTEHek2WuBG7j8CxTmbwY7SG/uike1O4MR/08PHawDHKmFCq9Lq
/3z6/sRTsseB42IMNtNJkCTTPTImKrlqPbMcJ7g/1PnLpdbFhxDOUIkE/1woxCf/
1LNTmmBJWObcDI3t7YtoGHbRJl+jFvVzm0xVKJ7adOdNboJTwtiW5t69BYD1qRZs
aoiKPH3G/fOgiI3phUnbm3vXcRoMKAgxgJLWCw2nZAf67zJ9GQi1xXo0KFM2gapO
Xsm/w1FfUAJx/y59JNLhvKPBbm/CetB28PV7Hb9XtZhWwAOSME3B3EbP/Zjcr7r9
Z6cphza5zvy3RCY8mZbTh2E4ypVmfV+mxu2s/Ob8D1fcz3uR6pcJu5s242d6Mdps
4hr4tLYPOndMlUHSYtD1ECmaWGUKue73Xtvua0enDGQp2z0XzkdX6AvQRGDhLKj9
hsm27uhXifRYiwEELMoHsM/D3E2k4COkrxcTA9kHCQR7bnmF/7m0Ze7RWKeKe1ju
Hxrhtwjk2I2Xgi9QVfGK5A8E5Cm6Fjgb+/eQTRX5+5uahVb1KVsFX3dTwsC2BF0/
A0zoQE823HrmgfzvytlWYh+VwBiUmZ0Np5NnW+lhTxa73/NAp+S+qREi0f6ExQl3
CFjAjmZav+WWB9TPdV4+iIIPxUuGuTYmtzIbkHRn0QNftIKTSArG+pNcJNWxZtks
73fwv/SedudpArXsLibrxizBm4uNxjoke0iyZQueRQMp3pic7yThHdkA0nSuaNnc
EqFT/icEUbIb5fS6qgl5zrpReP05z4GW9wMF2ticnsnY5TUZpZoJp6wGTNsZCcWf
UXLMrMQcm6Y6C3zOggI7yAFrJ1tdA/y0a7+2b2nImB6btm0TkezYqqyg1RSjvoR+
AA3nYV/JNOmdGjjgNeGbX7yrDPp8r4eZ5cy5R+6xzsTCHVjdDhZrjDkpgpDBY470
aM6JZ4VaKJ8Sx65cPRJLJ/lmwz2/R2eCLmGvsoVbOG+nW4pg0Tg7AxvlQKSqFlHl
4HDu3va5+WHDxoW0mddUtmtewjYKEBPYB96OOeeb/Hy43OSaYXNg+0PfklX2GQp+
D/ZYREQNZ9BrZsAZi/Lwqp65qndKy+zT18TACZO6+NtmGRi6W8ZaoTLVI4EKt9oV
VAWaDfP0nOQf3tE48EgIzlJ1f5miBNaNVGEycnHvjSY7K0gZA6FgLNddla7I7Be3
zD87yNtNPSeYC3/XiR52nsAHs7/Oauu19Ekb1cmQbiv4dYCgzX+xstKHknTJCoho
y0K6k9ouWbLyoOcX5eS78UPc2l+oOt61YsfWqzqoB+CCVUbyaAtnx4vo1H0bBB0z
p65uanSs4zmWGu14MtCk/TZ9NEyZOmcM4b/M/aGKpaZ2Fpi53l08+lfpq/SwllMk
NAOUbvVJW0R5foWbVjsfVLZdsj/JLVAU6myX4zo31op+NW/F9ZSD5EegBqg/1CpT
id4FgWAmZ2bqzhmt3YWhQqr49E9f5qJXAa3K/3yJ2u9ogoEKEfHi8XKqLGdcV/4p
WXvJS+9MkTJsYzYooNQp3mh+ANBTl+1ud9kJpJG4DhakoldWwtJmUVnlSySBoFZw
R78aV64Qi08AMS8+iYiklqBcv33NGw/06/WjNWWdapqc9V2YQKRHrBN9PptNUdvp
kAhexUplQiFcLhaBdcpE370gslw8PiuM1tTIPUx/d9Fyx0qIt3p/jJh706/K8G6a
wx3mjgNFClESEm+YyfvAX3JbhDIfpkRhYykgk7bhkc9haBvdgQmMiGoXdViBoCSa
Hm3xae+bC/R2Uio+FIEMxluc1u7CnqMe/JPww60v7LVwBOBj4lbyXjVnPi4RZR/f
RccY9kt44Pu319xUKun0brw1jttgLv9v0WqOyd5gXu0V2ZpZf7xWGQ0ce9nJBhTy
zcRZDLpO2FbEgAuHn2TAEWc4dq86yU8eZv01gjRW8cXuPL3kx5kkQ9RSfzeImEbK
K3NFEAJeTxdK9VlB+gTlqJ3roX6DfYDL3fzjCWtoXM/RmgIwj6vwpCZE2WcE3gZB
xv1g/ONj81jlBhFY3Mit6D6xVgUgPI3gt85wp4aJW603ObgUsk4fjP1Y/1a+W0wy
bm7eof2zvrVu9fcHN7iATkSuewkHzibR9pDnJcoknR3e/oHhjmnxWN9EHOE9LD+6
/3r+wkBP6v9hFZvmv/Wh/G6ouWIHz2XrQYwgtZwCsWl6XsGvilIPnz7gzWWKxYko
rGo31B3GaErYtVFBSYUosmti5gQVtvd8ywoejYR4foaFLThyGth5PRok3FlV5nFM
g11q8I5ff1ZwUnH1d4kAsLZ9rG0SvqTxV8rgMZPOzJgG68QZJdOS0CC/ve/AR/e1
Gj3kYutgKWJVn5AgnHA92eNLBhJu7LzL8E6ImqB7Z3T4Pqaa2m9TOIY7QxmXSLz/
0U1gk3fgmKjqb0gIg4aGIhT9eHlvvrVV3bHWmxTh3/0igCeu9Z/9M70D0bzxKBry
0SDD4EjKth4fDCgILHxpHjFuiEM3ZbWt1tkdWbvZLvE3DYckSJV3iaoS3BmasWpD
4Al2x+U8gfRmt4x4btdfK5QP7bASAfjbaJTsCBZTX/go1ggRL+ZVPZL+pMfBJsWD
oLQ5EqUpKXkDwDLTt2jy6O2VaDeaQJdkS4bNo/56Btff8Aectl/IXg0HrcDLXQnO
w+mlPnh7Amz9lOja2uEUS9NVrzpFV1bkM9avPQSnc1YLFy/zjfSo0tHoutoxJWhb
h72iPNmxYXNOoqtZuKgrDhfQBw5IiPmGx1W5Aci9gpe2xOiVCyejch1cjNtUQ19Q
IzxJw5QtmyQPgPelZiRcYeApDp6svJ9AvTms0Ruh/LzTy5g0LDmqgV7Oi4hWhr0y
w7nokAhifL4lc8HKFE3k4pWBdxobN2ajp7W/nSdsoIDz7007kvuNv4RAaHoHCEum
tOS5EQ1xeWI6gtvL+opxswQIr2GlpmOsqUNQM+NvuItCdVT2URgce8qzRhKL29kh
MSmK7070TCohz2RLDqI1lEz9l8+LlW2yaTWBXJlgOzJyT4b7yUL0mtD03O/UCVKD
2DkW2yQ9bbFcJC+/KEgVcRyL3UgoA4YOGjvp4LhaGEI3aI0IDGAEjUPwo0/8z1t+
9S0HaKFOySlzi6jeYZKXQEDXFIbSlEDCXRp9DDCI0H0OJNWk2RQZ5lcIvx2zh5OS
dUiG39uumv0Aggz+fiJzxFl2Xj544qWD9WPzmalvtr5jUVl9qlIhbSF7aM9Pvc1Q
sFmBd1eoqEKakyu3RvLN8X/8CfAlohl6I0v2vMmb6J7VV2S7c3iwwAp5kYuU7YAT
ICsGtPXMEPOj1jhv4tJlwx05OLVGwLUI7pNsRpYN9E4cf/9orhjiVLLorSfCQbDN
iD9zM2EOOzauaHYHtFY8wMvKR5XkUWaS22TlUDx0V/vUkVpCMO7X5oUEEXLcCDkA
RbVe3jQCefPDqMss7vBFdLsobSRVnmGYQwTjgT2fJQGCVbcr9feBx98yHfXCyPPn
5UjqRVtykXvrAgM3gukRhdV7n5SXf1LxlXr7xnGX1hgau1uiyA01hhINF9wloNtv
9BVYgRw1BIo8DU24IAWMZ3sqYd2OYQSTXqGU8oXIosdDOV/HFBkfgx16rlT+S0S4
luPmN6dfpZGc44/HhGP4WuP9h/I7gX8cbWqwjqNMFJMDqFcSFD4OE7nT7cYevhGr
m9IPplqBe9JqoWJyNeO0A5kzCHzW9Y9Q3XoVz5OWo1wI3mrpH5pYIXjDbDBqQ943
o4CsLHlFgTYmA8vcRbZ4ApC5x4RkgmnlvdGrr6SHpeXcnweKmsZ+TeH8AjcUk7aR
6MJh06liEdL4AzXj2SSfR7PSnEQnTBqwBVjHtgpgdyjmrnSRkIlJ+V7mPxZcWxP9
kK56VPRA9OFoo2c51NlAR/FCXHm4Fc0ICOOznfIwqIokHT+1KCXJKn5JsN8PIsjb
Nn29uF2itsCuiTcg9h5zFcW1ptX3gbxAxUcooILxAajfqoQG2DZFpOfURMqB4PGl
7p89wnYIDOMtaJ/8IugJF5l5rd2qkDrXHm1VYgYxK7IaF1YgOoDgbZByHsA8dnY2
EuYg9wc6wGEQA5Nbn0PWvaObo1GseZO/QpK82Mlov+doIGzjCAJKF50J0GScEXCl
e29IdZd0BjiRzgSX1WubIIgxIqHNi7opwmTLFtkFQPHEbnxxoLYPqWpCCBWSyKeS
C+3Ypa22sI9lEe5wQ6pQ/fsdcGmPZC3b45E01oQEG1S8JZn5/xe5Z4FvBXFRWa0M
ts9VYBe4wj3Oo2zBhi1i5pWCYXJrobQFRLMRnDttXDcR9z+QuYN1qBWBYSl/8rG6
Y3UBB6opHBW1K8lnxdDFy85TghipLsaTlw9euq58JAwznVHRpGu2S/UIAruLxSt+
FT9ldyLasZoOqM8cR46nOTOKHt41w4ejGY/DWFkhba2MnUKCB19zZmooy3Zb4xxL
3+57sVjl/0Y3q/qBeOaqGJpNNvASbrgmXAPYXud99v6gZ9sjrLYwCzuq+D7q7Ll9
WDw3Uh4l2zmN8NOC6fzW3mWQr4n/3fbf4j1GsypUmfVVOYcGQBBD2X/rb5DD6yv/
2bon7ajsAzwWDSwqQAxKzAOcBM9sWC3YZO8ufvULiAUQAvS7zztK9bCZuni/OnrH
nTWzWAiMYH50GtoN1e35EdZs4Yk5zeRwX51zAyCih/yfA3cM1ikaWhXyyUtDMmD+
gNdrxyd6Fg8Xzr+gRHvvV+H1+kK3qMqPEoKWQAaSyzhEWijxvoEwV0GVaycZoW5N
E43x4EBQixBOShCit8TesoPsAVcMUzzZpp33XUxHKrC3LO5F/HS+7cz2lh0slPI8
u+BOBBLeasQWtT1818D/tkKnGwT5mzY+wUlA27cdqfJE9tlM8LHjni9Z4Ubcg5WV
/F4oUbR0ak+9/0oypBBqXRYynE7nT2eaNhVxH2J4WjMl6tHPeusH38yRDpTOKsfc
ewp0xW6bhoyPPJbUPe7GB/7mAw7Mtwe4p0TfHMk1G/Np8/h4ro0p4/6IfbRNFbwR
c78jWIFHnOtopVm5BxY7e6pgQOqJx5+7cyF4GwEGk+Wo8ddmqHfQlzl/FzKvZ/GB
neU9RfVZ0OjA1J7ERzCNMqL8IQnOMcIhs8+NEwB4bPdoWUcjQy8NhMvr5k6CT0ZL
89oVkuh2U6/251XWFX5T3nhmj4GYTmHPJOo6SvQtk0vSuGaa7ayDJ3Bkdf/J170H
zIcoGH541ywUdLN36e7h7tKSozetuVdhWdM4PBITWdDWg269ADpFkNx+Km5w1r6n
UR4VXO96GIdodJrYIQQ4QXcqFflcB0FmKBsFQlEh/XdFKUa54ApNz1pvk8snu01q
Usck+ugut2jx5ijcfWrq1LPW0S+aDgyfTMoIdb6b1LgWYISdpB5JlyhBY68kluRg
0m/T57YCsWUQBFX3smEcl15RXzUQkx7rZ9mu8M69+TSO/ozFLd1vDuHj6kGDER8j
WtgFiiJIe0Ck/SuKMvwzvIjYlwM4eebz0SmEb0Q1+BAtDATQoflt56E+VCG8M8Be
R94rc8wdnuViq9dbdhBV0FFzDe5/2wuwUq8VbNPLKNqLALMPl+b4WJjvzN2WXl2L
YSMlC4IggotKfEGrFd5rorkz8m6SRspAb9fHNPOmM0ORap13+pDOKM7a52TJVvjT
BjbW1qNMRG6o3tnBKdmcTzlvwD1PqmYZCRaYn66x/H04IgF+R7mlrdZ4HMZ+sR+Z
XkmZRGDDSzh9Tw0aladWhG8+xPoXuPvhYI0afrfXks3QcHwFcaj429ahhLWJq/is
KeXf/FXvZoeSRzNGMcuXIZ/7x3I8q5CdvDTqHA2wSPVTBDqXl8rI7JkrFxPVBBRu
rrjOG4SX1pJ3ldRcEow6+CkYlJtxwN6M6ezA0fnNTqKGfV8nyhJH6nIIKzFHMqeY
BWqjPQjX8HxEyhTNRj4A1TR/HqgiNk4pdbp0vsL5KOuAfddxeZinv9uJeWabTUgn
R9wDDliBwYYAEJTxFVkRB/jsg86n6bgl5iBtPy6EOGgDWjoCD0do8F56SMuxgn48
hs/kx0aK6JLWeKKV0S+VRcVsywhZVbb8b6jafhjrD/uHitIO9dJd/AcWKyhTRzvQ
5OBLaG1WgSqbSzEyAcg3JfY9ycHGoFIixok27OzaRCe5FFlFTkscc73D30p46qo3
NsmKTdHjhcaahUWCh28T/DJjIFfK0yM7aZx3RlNPhJ9ed0SaG2oX40U+PqgyVU8m
cCxkAC7CtI19Ku1nSZwzZ3Svw9U7nRQ5A9KR/pgnkA7HIqkzleLXMei+fgpTHxX4
pwnSC2O1pmkJ3gByld4RXo70x3odkF4mrcIgEl/XCtC+dSNJ3nyYtx8G3AX/AAaL
4wpVwPULCr2bQwQFtUxEkVW7UPVEzswyxkJzASQ4gc1zlsEVzHYHKrkyzPERzszq
oyFUOXsLo5lP+dSbyAmNTX7cc3cOqm18LgV4cewAW20EG7GC9KI+ORPbBCwH3dGR
SpY22Ax0Xk5SqlzAaZEQuBQwyJj7KndS9DL1tLaxxpei5Xgrf/3xWbjZkgb5ea/x
njhYYOIE6MzyYcipRK5a98Am6fXkwYUVhnps07E9eE+utbGVq8wkE4ieIRGTVhoM
Ul/XKbmUtPLmfh15xkLcoz0OnvQu8RuOIjP/+YyaEQ0Gj24Hno2W69vFPZQVyJ1Q
AW0obJUGPTN1pPUf1RHKcd6ysDjxBZobl642y1i8WlrD03RVhvPHX2T/7+aPHN7v
G3yQkJEsAAGQexzsaRXk6eTnA/d0IHfq9ChNEnpTn4kFVsbUr4ePCO7smhSGo21J
xncnWTTxw8S4b4aLXrQtZaCbYnnX07WNfNmTvQKeBQcDlU2ssL/+cre0B6nBeUFS
24tcuPgHG0qS2EyQdc38QfrIRDsAOCrOJdFcUTiVkmwbn+oALxbTvtDu/XspyiZd
6Fv1HXnVe0Y8Oqq+dN4JedWWddIE7PdSPqCQGcnHJkyVSJqGAFK6FKlEO9ORf29D
38TNWnaC0a8h+yJvyDxmz/40MjJiuTEvQyahTitkMQOAwfO4R/0T/MDDezXLsaFV
vr+ti4O0BAvKbUQK0rVxq8c4xlLUTr0iGQCZQQiQX5U6nTdD9AuCuh4teChHI4ZR
faNTSTmn43jbPMLKThaJhSsVTPlVIbWeLX9Fuwe/uIxnqt0YZEHqh+UPpyAm/lsY
aety4ry1EWD5hSJqQ7yVNIKM7EZXOqwha68EuvAm5bIAKLELwyyclFYYQLQpgG5c
FnqRDX2v6Bh8vAx8p+JCeFhBHsnkR44AwCmyrqf+StEKRTMFX9wuHoXYFAi5YPzI
gC2YVAAOlRExl3QHN0ZfbYZ8I6aRR5dXG/bCBvrxShSAYFxMdLZ7jwBfp2bf/R9O
m2AuctgnUdMoSJw+vhByuWkvv5jV7T7d8FP/cK5WhT4nkrUFUMyqovkb82PUlGNW
liHtTLzPv4yAdqSqh9X2GXTyeCT+LISQHXV4CuWjPl1Qz0bztbZc/cjzbQq3YgWX
d6uVI8s3wK03h3YlZhcUV4Otw0c+AT8KeHkX97qZIYEvfActMUAFtwDjNUhx1/eN
vdtiUY3B9/ZQgsbJYbNTJiCkRN/blLDbRyH2O60Q5VkwFWKNmdWNM+Xtj1/A9cPg
QSNJlhN/lozmHYvNASjLACAIK6Bl+E6Y1qtFuxv3zuSqRU5sJuCdB/TcCNKNXXgK
WNMiSlmPWurmb5X99u6I17gXqGKhOZhwRB+OYuDEIN2mNSCHLr0hDh5hzWyqY+cZ
SlsvYC+qc4EoMAngdYvrYdF3cDKy/CO5vUROucqA0Hrwt8Xl1YheiapjkZYGYAsc
ED6nawl8VewRVhwdIb/yVWhynD7FpxAzXYk9U2FHmcdoGdIPHlfvfEJhNo4KApmS
PgKsZt3yAFwV2FSI7ZkugmpH/sXcDnK5qSGTff5t/hV/KmXkJkEgSia1iDzOXIvm
uVgUf+pU8ETjkoZxxwloPNCphKnOXLUp9C6j4HSsooby2JAqur5xvf3mK1WobvJF
lBMc1vS4OVB7PWm5DKpufA7HgzYAZOifcwTtvGlO0DTY7MdEe/dYutd9zyorQLYc
32apkbaQyIzpld30vcauLRSEw4pSm13vqazKGkodAgEZH3rQ7YFXaCORoNgU1cVe
os9+12ots1ItmOGGLUcFvgefyt67TJt3bdW1iUsvarD6XNKvCPJenow5upaSDLCp
LOr4PnETS15T0tCV9qbCq5VySCzqngKhDkPgshUfjUuYK0uW+f45h7Rtwb3yhZ6K
3WZqtoDfjRgZUl5n16CAdWeSFAOU2sbtyBRrKoJ8bf7gLY+jnETVTWt4twnycLl7
0Np1Frel14JxsWrx0I7bPueihzfkdCcAN+dLK5LrEn4rHuQvWt2FrU5zJDfsqLUA
YCmSsbbtYmOHSwoyndR5hFvG1KiIgc1VrSfUPyX/J+EA1Jjhmg1+nJiPFg5Dl8tt
5+cT/LmjLmMO7zqVvaY7FOtAZCApr6X0NabzPwC7X2nQQoX5UEhW6DiRpYi2me2H
X8skBx5auv7/676W3LhOIPv7mMm/UkJ6Er+dG8nNgM19nWvUDqBQFNsiPeWbube+
v6tc3GjXie79Ncd3IKSO7W2/2hGmmpf4hnGIQHmkHIK70T/JBeWD7dQzVelGGoyk
9kYaaFZHoW6RyAjyjHhADB/CisU6wmCA0HE92aBMvoYyz3L1xE2x3czqn3LfY+Ss
6Olq9WMtSfCHSxDX0OOHo08/U5FAXqB3EgGnUOraTT9rLURAfj117Gs4aWZ5Q7XH
dh3HUR5zlKTucBeEL58wLHX7lGdYwdFIctU/ux5U7PZoXMZ8X1Fek8Qig3dQis3k
E+QcNg90psvuqsPgi547P/ytUkuYJKya9XpdoBZjQ/XAETfhw24RROheVY10N/uS
71NoItP+ejdq+lkzC6AsskQii8TgV+Cs539AGP+2Ixigy72Jnl9zB8fvwbcdjobo
ac8UOUbSBufEL6akYNQkWIy0NZIOTyK8cQdT8+Sxr2W4PrQIcggm2+KO6gU4HWqP
XOcwdeARyl0Y4GRYXTOsAy+kQkyqX7YkXd8vg+G9JSeRQTJikESTTXEvrmDM3kCw
63DgVDbBarPC96H7JRepBowu9kUNT4NBkENYvHaS+xxp20ZYsZOqX9Edk2+fPEOh
qGBKnorCEQfs8lnEHOlbgFuaVuHo+cBGonq4mKUYiOx3PBXQFelsFWaOlcIkppeC
pQowOk3zFmdDSSBuGN+Yg7MRyPjahYKmfqVwf/L+MhQCrU6mx/9yhu8seHsBDKZL
69CDrE7YyU7tn42naFwoWWDEIxfc3DsagrIb1YOp31zuMzYT7g1r6jcAfhBJlbTk
bbVx6Q/JyqA+HqUs+SZeorplpEk3qB+3lwuKAI3BxsyLenTzrb+C8M75O2C0SgIi
GKJohYsSzrFquVk1p2sQY9DbWPS/ctNdSjTMBc3CTINnXJStVPUfiOKxbxN7rKvk
xWe+vuUT6vIYKNX3tnZekjYKVBa4yBanSuIEeaVw5qS257BIP3eBDNbgpjjMzqBy
SGyWZOfE2Jr86KZXql7tVPvt6ZMNSyaJ6XUyXC/DB9fwo+bj56V/xTzrPpf4VSLT
U924d58Ow0Tkj3tSAlKm/nKVcKjnx+m1+eYknAngBNat5QZwNl7Pl12/gi8OuE5T
qaikeAFWlqv2tg5A+4lMPgvswLEs72HsKQxBQtLkQ4g7nSpRA7JDBAxkIHghUJKv
2mYH3ZB5lcmpdkhTI7dtxv907snHkvQ6g1nmEYFIB8kBSAn2spyk4Zret4DKKmtq
ZLoXKKUN7VpQGqORPtitCru3O/eOp6cDwdTW+SeAFZwISMReRM3yLM+ggNrzhaqc
L8W5d70dgHjYbsdSk0z9JTr2uqKaUuE8ZoR8PHMiVIfBJg1ilGQIZ/kl+VBiFmRj
YgTBN0h+4n3qid3QxILIbOudFEPQkHbyHDqFUveMoQxJwht4dDZCCS/1+StxK5o1
XKfj4XXBgG4TD6wis3ZHsGweXlraSeySUBP2PD+ALpPcUNy4sx03IdTALFQi00ah
OaT5idCTLhtQnOrLj0QJaijKpaZXbhB8qrRsDqshRkSvWOYmPmlyJpNqVSB15gW9
gbeYRabbLarCWzWavYtUxT5faRIFxyJVOGVjcb6psDBl0QrjiRDwQo6hvKwCaNT2
joSAIWjm5VP+3yu6+Qfaur+Aq+7N35Chd+um2Zlhj4thbge/Cktcq1PRHdbl3Dwg
IyUQkWnFsUCeR/+vk2/Rj3s0YD20ehMNpp7HlHAUqh3JPACrIcRp6Q9mcfYrWzJY
Q7N4aWgSnEihpmi4VMbDfPQU1iCPYR2E51+lU2iQraE3+H1WcLSk1YLfYBaTlsYu
HKMe/SnQ015zKT0e7mTRh4nrcSpSOQhp+x4Ky/GTaPcp7oO7fnKV5hHD0w46AQbh
MPPGiPROnadZfO1jbZPK5ojxECnLdwAX7/2Cawv8h1h63arx3BdxmQ+o/zq5Sqwa
BK5oG1qhKBWJNLPutEWP7eRN1Y2bnuvmh22lhC+hEogJHwNayHYqb0IYz0N+8JeF
7UJNyaHdWiKe2n2UmYOWFIeolv+PMWQbXhgF+heyuzKCM31cRC2lskf+8ovakvJz
4f/Ly4x6q2GaAU+A5Ju0fJ2goC4HHi0IzCYgoYJjhhJKjX8K4js9SfwQScvII2Fz
HQfxdDtEjVwtytLv8FG+5uOCZzRuWTTLY+eE8XGUrOTpUE92PkGhcWe8ccDL9jqK
/8gzifIIyU2HYmUjLi5r3z9iTUQD7rdUQiClVQv68lN6gDUsNfbJZssc7MY/ss1F
kt7WoxEjPKkyN3fiWESsGIFyhDo/DlZi7mGoVy6tgTDWQOpYdhY4CGZByCkw7/gC
pqberOZVkB3AJgJ5a8JJbIEwhD0zm+xoCoeDdMZyiJQzlVygfLj4zJeRGJQdsdht
wBolm+Ma5dV93nCaxKJP+vlUgcPhufCw7jgZaIs10oXftmLeeqj1HoeZPDsMkLkF
MQOtAg9JDG50Mtt+SNqiCaOqye1imXnFfcxlpJNvH0Llu+Xi+W7ce1xAe58211oZ
6g64+4HsBQnHn31u248VtTSp6ocr9wzwQWuWlofuNwtu1Pzns4WDaLj46szTubKa
o2LQcgVUQMoRKwZHcqf2GDQoC9BOkeuNpheoLT8Iw7KuqXPOlxft0OsvGMAbgdms
Jv/WuZbnkKPK+nvC8rsnan/2ssINOTNvglAgNA5URI0BUjIy3RqHP8iiBc0Wsjnz
sftnaCG120yJ8GDI18FuUyq81PLNX2kJZhFb1Xo6HIR9J5avmLOerrylScdlxCdS
rdU8lCCDKGyaTctIbrxjkGddT9qitk59W1rSzz6GxNOv4w+duZvSGgBMQ8BQmAj+
RP6DEikiW5NgB4Dc7WBr31oIvQl94VsuVaX2YSwW2opOMTedmQL8Lvdk3LWslflB
ILxcTQ+DJjgRs5D3f0sQbPVVJzCtd5Dro3S5CD7dXfLQqKgbgzO37awmDz4BK6b5
0dFgCSJmABeWimlCZfQPhqb1Tw9JOyGmGaWDcjvBATZAk0XO84RNcxnIXqLy2r4m
LqrzoncMvOA2MwwaY5U28il3ejOU3w7znhglIGSkztRb3qE4ckY686LARRdiysUB
q715IAkqDkI8tfFElN6nsIrmVmxwHJN4ynOSWPo74bB7KFm2CdivCUAzak85pUMb
xHjk/K6VU0fV7yDWvayKgYSAYUBfS7ZYq3b3sYc28W3sKS767nTCpZoyP79azHdC
aEk3TODlsaKYrjcQ7D0pa70gRy8cqo5YEfyTi+C9wvI4dXcmArLb2kiv5CjHLwS8
7kr0zceNboOm2hm6hRuz0+HpQprtYGtArgOSLfjR8xnZetnEhdFSLTDS6RYTv3pO
PDwzbLfj1AcGTDdmUQ+oCRKfWaf8xGO6VoN4NXcq9C69/bWEmIyEg6HvLRj75wj6
nCtV24bJpSpVUHTJZIQVpfncjOIRGvp2Po6yYIR+5JLUk39m6oNevZ81Jfbl9b9j
jeEtRTX4sYf+YSgJlSjVNiT9N8cS16iy35se7k2Ts+g0khbW01T57iiTe1q6HqTL
YhzlaRgiG7SSUii+L7xn3cL7KkhBcmPkoquZCvm4457e/hS+wfyQMBNKFSXlMSkf
KXHJ47y81KiS9E/lpn/45+x+1mIgWCxkVGgc01JTJgEGhXO/j8MAbvlHdXXeA31I
pfouIoKjGH6OLSfBnG8btb5lB/yleDXKVvT9yVaFwi9JRuqOUypIs1Xo00qU6gpA
9cRJ8ES9vnXGhUSSSGlXP84R1UfbQSR/TCYH9S9essonxnrQ0uuP1fvbtUCJnmpX
GrlFmE1o7jIY4+lMbKqGUh2oF90aaJpRLiEudfObzqN6ZbpYHdZ2Z51ve6648/g7
sWzy0asiRZfnSqa+aaYasn9IeMq4DEqiRIhsd1fXGSyb31PmqMAU9/M43kE0IDcm
zmKFuxUYBPiqSzXJG3nXY95MvqYzvBRARiLzzUBoCxjnMI06VxoocuwnF0hrTxBY
rKNc5I53oof/vj0v/JhQVztCcwStRclZR4GjvrukH6utl927xBDUAdHQBw/H4ty/
iDpaMDcFfzrj/2WDatNiVSLsf74jv61mdbWfq8Sr4Qh/N41VkZBd7j7O2TZmaURu
rouwGhoE65+/dCZ7bhXSBiBdC1GmTsSMK6TsMrTU2ar8GznOax5EDBH4hAIwxi6C
iYQO9WLFOc4Dbf5QNus12Ia3yA0eGvkhdHgHgoiVeJDzEtEBmel2C1ttLHbhLzb0
+EJJyxmGBHZ2JNI88qaGJnbc0R7A6T6+LPM4yIxupO/3Lt/31ppZR+IiTm2wnHH/
AQ7jtuDkcH59uAGjdLZbxlaNjyn638oMWpgKyOShT2YvhqUxV9k8M0JxFnwdMK/F
ErCMgXatO5MKvfJLDJukXNaCsggE0sMbTq/2h2VnC2f6yJ7p7KeHzMPRJqGU+8+N
GKNd6o7QTJL8xpWKTBHUvOl6xEbHiBskb04UfLzQwoHseNqCcBSp80j7Un3fPjaJ
Puxu5B07Xw2dYRbU7ADZvMg+WFhu6JXG+aApCziEpwSBGTNOgenzdz3D4WuJNOLy
989WJTyr8JAXEdwqltXKaArEoMnvCe5AX96U0iAzsyun5FEmyrYDG0z8Gn6ugAmQ
dtg0wj6pktdarlEs/4ANnXqJ705fCM1sASDK74mDNlFoL/6XhrxYTa/cjsGkmygx
EcbWMqJNQXPC+jxZNbx3EcKiRBohHNuZxqdxPtx2QjkQytxbxG/tJjdpKjctLLhU
vNEQYdfFVZg4lVloP+25yoSuKsTTxISmQMMv9jMmO87kmrckN/IpFjWj+vH+OChn
rMiXzzZlizsRgV0Bu4S0eN4ZjLgmDpq8OF68MBvzCLhPUVR8O1tUwj0VkOtvMUyI
2hRiHqxucxN58U6x7jLs4cOq+7z2GtgQX5pJ1VuVfehrcdOOPSr2OtCSWTg7Nv7l
29IkOvkoUhpbLCr+zLjP9vAofjGZ3H+5TGM3+aEcCEsEDtBl7XqtbkICUGmYCFPb
DBDO/RLmvg56gSQBxmUr5bAa0sg8tb4FhZrDtkzINmpvxU4zkWI2Q9emIxnXjN00
3I7V++dgxqjPUssHOl7uNbGBkvj6sXjtfYtPg4kCaw/gVLHJzOtQfU5kBx7NRnvM
e7hcM00qJZe2d3Q87ZmJcaCXMiDDg1t3/6MnqzPjb0gzaJSt9/m4ZJ29OTF+Zg2B
Dr2PkFaYYJ4ptDkeDkxGgWmjYamb/5a+b6JJ6ucx7aEYQHpI1ktzV5xcY7bLtPiW
ls7J5BOt7DcH/cxbMISLQWxdBW9tleMJSmKz/1B8cyKGX4NRnssUpGBnWZbIuygT
KNh3wnGe79az/6U883zOdTZBOvX/q4vfRt+DjNK3oxNiGhw0Ib5mpF8Ds/zKvFcL
om6Db8Y6cMAtF3PNB+itdbz1cOFB5OYDI4ebDC+YxNWlNhSClEwKIjUeMLYWoMkS
FEHmOuQ9T6AiWODFKtu6IFd/B1evN6kUf3MCeJpVszRqYurDN+mx5aoJQxeCbK/l
lxSk6y0HZKgwCHx1/g+85xzpAhucYBcl2ooIbiXlRbalN0+75Q4TJCdR9vuWLL81
/jvukRSk2CwSResD3hpqY87SKX2HE9SCrQwhkwtneDu73OJ7ZrwKL18HZ13HCDau
ggyvc4MmaC6XvXpoJGDcjBbO0Def8wOIXywmW51960rYfzNux1I/Txpd7wTw2yqs
ZXI+/mmrbmerKjnp/foE4vTOj3S5QDwQ9R8RL4rxx3JyTtk58va8TvotVPloxviM
RhWbS2+PDHs6mZcy83E8AlHcBpOl3Ybb8qQunywh99E1MsPcvZoRgY8/THbEUquy
aNya3jZy8csgDxcIUfCpMmnsBIOt9pSsfrFXmCMIZECM4ssHpoB9ehpSCvq/9kpY
1p5Wgza14CW++Ew3jAvN/jSw9ca4iVzXcTLtIWn4gT3zTH/TJL36M1LiNhXjkSz5
hn5ICIEoAgVhErLUytnnx3NvkTqTUNtca5VSqYk7Soj7exH6OXRFEj6UhX77tJTN
Snlf0lF1DHnco6ab1jPxBdkttFvwPuKXIKxKp9039kKyRN/+J8RtEB44JicdQ9T/
BPca9XBNQC+gAUBK3GhEz82EI/fcosHYayuRpQdRQkeOE4KrbyprUarc37CGXYsu
LrXqY0UODmPvteQLpXT53L8Yu+NiouRWGxCfry5r4fGX8caW56v8FErp2AOBNk4m
8gzIE1c/9PY1C3NZLwRKlfFXYqJ3NwJdvfkyqhr2OF1KAfMXuoW0/qndkEi8OGmJ
+N1+GYlih4ZQ27H+blF611dQ6YPlx7uZHZVDp/cp15XclIvJbkIi3p6/r4cXp41P
gmEc1d/zFAl/uEzfhprUDGvv02P4lKENrT8mB0+cF8N/wIfnXX1XPRkk7SaPN1l5
1D7iMlIVDXYCrTIYQ0pFQAkc19+NRbeikhgnBktzr+d9Afo3b2Rv34LfSSHchc8e
vNB7517qCQ8PVh8fn5RM/9Jm9mugpe/6q1l1bUqde4jRqGcL3pt7+1Gcflu/GRv+
2JMBOz94lxvBE9zIO38700GUPVb/Qvs4PcMgBdVi1GxiyPVHQJrsDtJbkrHgtczd
GbVA3DFo1iySmBCgkbf2SX4lmmTvOaIEORfCyXWkXrTHwgS6qvxcoDAi2SLHe81p
seMrc/Q3DlC9ecy7LkqARXeECnVNvd6tCeerA63d1kewYps/8JXdpq3dMXaf426+
zw04iRfuebQiKQ1uxNo4yr7Kx/vGaE6R+3kIowgNodJvCSRnP3qiiIJAkzzXfTKy
D+XITQbi8GXbIcR9EZwhF4E78IlHM14iRleYuL9qAAKKENSbkMyO8p4qVK+D56RS
78zAwFt6WPgGSYevuU4pg9UenPTG3wtaho4UNyXjUEwC5U/Dt1bluh5ZPcSzosgD
bHNXp5tBdnUr+kMB99SZ/BfP3lBmlmOPAnXZ1Xj/XqQBXNUqI5CRkBW7aU/uNkMu
6ONAOqdnSMeg6LJni/SXtxI1u40exobUrzYZK9r9RQgTuplQEomp5bNGfum9+BGB
qeqmrEbvGm+hRe3TuNgohqFHUAK7ImWKrqsm61tnJZ0zXEzPQRkflew+7QK+Zewt
2/UjuD6Ev3OG3Ocm0eRe4UEzwpnOyLKaLai8BLUcSh0yOcLXkEiesajEXNnIzKGN
ddTzCB2WZOdI1MT4IWyEQ+8ssxNWbLXX9+qbqOQTQH/UJPao8qWe6qJK5EhciALg
2zFhTTxjU7r9yM0Y3vcIW/PQx7uhoZ1hlKL+/HEkyw5QiGq4xgpZt07eCYi3csnU
VdT12ThhjpAjms3OvthvT+GhBOiDHMhQARAX3qxJaiLdH/UHQwRmtB5USTWNmVL7
3NtzX+P0nHYkkIUtiuwcSE8ocE5pBd40yJITgGyG9Q4c+S3ycCxEECITJYdYhfQQ
KWM9lrN1OSXq14NGitX1mS8c1NAQM9ugJ/TAaY8QlXXmxyi1CPScFAcOMx45DNLR
B6meHTxP41+ghpPGbLj3fOqKH44H4D7zhi7785b41xV3Mpzn+zjRNK4/3yeZhI8a
qPXMPMHM6ZW99lWuH7eSC2WVL9Ofmp25JT18xVd8b82f3+G/PnQqcuWOcAcJVj4i
qgVjRD+pH+BUThXvM8KmWOA+zkTeA9W0onk5pCuqUPPxxi0h3PU+CG8csO4lZ/Bq
8zMEptS6izBcts2InFcvpf0kSif4YupK5pk6cPsyNcD8uLmT+e3/TMLid2N2rfvP
TKM/xd+gJaSV+lnH5eMB0mn6R1tSGg/oLBNqFUYn1DssfIQr1EI7Awv6+kQo79MD
01PMtbVZ1d8xqJ3ZYNtBcSSVUcUzrSirBc/wU+9FuJySi10T8kNo7YFEJ73N0Zqo
V2E7vVxCu7UozcFIdXwI0yg11xTjd8cyxXfNe6NzrJanlFIKc3JpnoYvxzAjGg/y
agtq4GkH2aqtV9wEY2ONx0C0ANvCgo9Rapu6vM+Xa65NU63A5g09ljUuIJRDeLXP
+sJivlP8qZGXT5GzHH424rIydr8hHFZD4IyB0RVMiDv+pL0xmki7RT1O194zHjXn
Wg2lScjHnGWNFe5DxKvMav/nnkBw9RrvU5xSqNCZ6CM7RKWK8EJbhbOYKU0t2l9f
OOkmU2cf7yaOIhWPUC111y/icHxxrn79ZNGTm78E1MBlAbFHGvcU1nU0/PSWg2Sb
B6TzgCxBIsBgrzhF1oHFHVU+8LXXPV6E3fRuR5Zjr7GjvJg3viDg42M180EDC0Fn
IgKaBJhmSu41UcZ0s1ShUQ6UeIaEAClZLyEmCfdcIcLBJUerWj3KTZmnEIA7AQUa
vhNY4Z5CstLexM8nap4QqabOU9ib6gOfv2CoCJSiDO2zps4auyDpxOk3GkL3+Jqb
zCrsIcPx4ey65HJoKrUfLZ5Dk7+4TffgX/Vn2apoaIk9cGUMTBj9flVJtPeVZ6RT
S6YVUCnMMSVGLaXf+QwKyaU4lB2uLwl1MkyeeJrriLbYS0SSP/ZOeswLd0HP7VyE
fAsL1cWBcCF0jsen8lQeqzq6NrLkm1s75I+gApGsIX7t/Yda5dw8kXNyNp9kELZC
Zrrz+9fHIVr7eaapKqofNO6sNiriUb2/d/QNHFIHZjS7pT/dtH4OWqVwILM8z2ez
Ut35AuqBj5UfQYTOt74lNBW7fY0B7R3sDsoYvsgCl02e+2Yu6uCdyfPrYCjwUfSv
XAR+P0oEDWG9absIx0fOEy4N99f2wVrIlP0JyTaxXPPHLDGLKCpoCqJ5dv/sqAWj
TeH+Ytna+cRVc5dLWtROwgjAe7l92Lm3BVainVACV4GeF2oEayg4ZCGTCq5MD1WG
MBIdGLTSH7O4/1io1nn2tm8Bz1Ty3zm/NGZkua0wLkVHYm2/5PwTjtj0p961H5SC
73S7AMpHxvtYouTcO/lGUhxB+eUv91qd0SiEIdeer/EzwuQ1Hxv61FvB3IRkRRWH
kHV4ZtGrtcX6XASCwIeOxCCRMSuAVFJEw+jaeXzdbAudprHN+UGH0/6I9MbcHlfK
6lFpLe0KdmrT+q4aqrWU3VBoTW0VU6cA64BdyOIAjIzhqYmMzoJSDh/hxotZ3o9Y
x5Mrcvv+sYRbGZQLYGp05Lyje/MiKW6oPiblSOwP+Ay1QYJFsCwEFuW9exUFPmCs
foqwx09RRtjjc24uGirOravcpWGoXXxCknVXHaET6d8rlqFdB0c6WJEA+uorHCgs
q7+pfD/uoCfVkr7mpNYcxwr7Wc96A3n5RAjrzZmOED+qSdFJV92iTYjAsEyZEn9N
G7At03bKKBHRLIyhrKiG+VvsAv/7IUBiTopnB8W2ru+ziFsR0GXoyG+gxQA+6G4x
VgJqmcs85Zmyi5FaecInQqx4AIqOXajYrbt1h5iZqBw3asWuCSEA4cSsUib/7TIJ
KWHYdapthrwUpWetdYOBxeqiwOFXAkqD+4JMSy3WQr6L7wy+LDQ5jbqV2Pd8z1cm
DNSdkAWGw9LSg5XZ+AjWBhQDRc91xag7mShYnz7f4YF/1RWrx2Yd7Ft/gD2DGi40
plQ2+40C43Gw9Pgbz5O/BTLoSvlDts+wZ0zAv9a94FujBD0VyNx7WfDnawSWgjAq
0Rg1dxF2MmpkgXbiNX95Q9bNyVi+DHPcyFuPLUWly+5bV+DCXhPCa2xSpMi+55Uq
fcsQ+juS4fNteVxk9Xe9EHlJ1Hb3TyTJruPFpNeKRBLPEwdA2NsWUKTGjKYhVBkF
mnDDiiuGZa4c8yO7qmE6F+F2hEtwdOzbRn63yLCzcfCjHCXf/3/08oLH3c0zNBAn
+2/WS+IcX/1L53uWa6Zwg1R8RQgFNhy88ngOvh7/IrR/3zDyTDQpuVdwz/zlyfJs
b3UuydA6CKxnImXw2C4/UHVT5/KiWE1oFP1tiOdZ21q5WAerfA2hez4mAREiyUtT
ljBh8u2+g+tqVQpAjiV7uFimLU0eog9dLqBvx9swkdB4auLd1ZH67IjJ5bRAEjO5
fhZcQZhc0pPB+cwxv2AoNBH1SbZu7zy/cV7RnZTHl52vtVunIkz6cgASARJmYMaa
XahXvA5ZyrQOeKmSYjWSgJS4qQpLgP5KCgO/K/8LHfsZ7TX8uLfVfLJMmuIH/XsL
RqDHlAB8YyBQwTPHHFcgtoHyyh1Abth6GpVtQu0yXqbHZJQTzIiHwx5MgUZQmHD5
oKXtndNEDmFDzfjrWHU3qkVwnJ7aOR6H86ualaNPMUp2fHH1eigea7liDqjnNZA7
OfLW0dWmL2rOTgHrqvGndF5LKg3JMoCeLTW2U44VCZmwaQkOkafbg3RrdJDyst5e
twq8VL6DNt5evqwZZtte5AeAEvxPJDZAhdCzx1y0aFT3BtkJBfGRw+QCU5UT+mO0
g2KindNrJ1qHlYMXEnTca65TbKquaUeV2vULrkzJUVwPRKrEZbr2BcAyR0ruxBVr
GEF7x2nxylzpxO4KON1uUi/XwbWOgNo9r+aHAnwf/k3e16Ashu67FO2Nrj6NyQhB
R0z60JhTSUKOktU4LSeGU7i+KvLFzFBXav2CLv0eAp4vf2e6thGB8ntz6cdSZ0A8
K/k5jVGwPGhTWfuU8L4CKWaqLdoWvt4ebgBnbJADMdgz0GDscWSYRHAM36BRsOu7
JOM9MowPuHrE7KO+9CBseuDO9+7BGNGEYi6WcJ/4jslW5Z0FtiazaYSlDsc+2S2w
r26Et7KaX+BX1xH3HhE4sbc5PBs32flwMvflU10zEucRe1aRTIT/7zTGaRwSDvsT
H7hPlkueFfF06z9qGCbGQPCXvdFVcA2BFrD9uWvI/381a4BdDDhmnVmBcROyQ5e0
Y2lVK3UKn5cmtBt4wPM1P2mOGIe8KPC+n9US9tjw8Eyl7j4heXZy0vrchCiD0Ptg
RkPXwA5hPWBBrNlMRi1laFMSlLYgoZTbRN3taqAdUYhbKDcqNwv2KRI38sthIr1p
unFsS7jUiSmKpfnuxDRsuwfFKau2BaKjFJr02DlCQttSc1MGCr/ZJFAsrwONiq8Y
oAT+RCfyhH4e8Bn6mWfff7trtN0cLd90oi8fLIqI+gODU4jWsW6VKH+WE/RPOYGX
O0VnHDPZMYM/zvdiLCv/sqTGqom1VPENng+8D9dBQVi2O0ZP54j8hKPuW+nS26Ni
TQ9/mwkD6QK1ypgT/OqEcqjYoK5roBVAK0vGKyo9YKxo08LQFZhugmyVrOQi2dwT
E0QQf4xJGXSXC7aydpDZEl//tRnw/ZhsxNXJOb5D0fRO8nknGs/dSjiBmGDzxPrP
lUDRJAosKCpOiKMOU14i0XkPO6NFn+wg2PWzMG13mdi715bOjepjr++W8KMw+3PE
fTcf/FRHhGiIXYm/gVp7p1xd/C360PZcNt/ZzKKVBGiofKnOjqlUXgFlNr12IF2C
8xTxIWHMBJOL2RF7ANZn+W5b/BoL5rRx8Er2ihlt/LeJjPBI8+MrCMudtGDCsluG
UJ9zYhBIkXIQE1LyBP/PwjTe+6hhFdAvWtPEvlR+TGI4Javf+D9vlIHeoyGd3qZe
THTbWUALbNk9MnuI4qU4Fm6FcR7ncQ+louxiJwnxFf5uep8QMA7xugnDH8j2RGW3
z/g4OEd3uJVwGkA1QNuWnZIafkxLme2q0xs/jIdjwobiDipGkleXca6Pz3FERiQB
yobCbqtrJIwsBWnXErP8DC32YtSGvRdyFU62matJ185NqqpWmrQJ4hf4DGK0L7rd
SAVi+gM6Z/Q2qSUwwOyl2Jnm1SsAuikh75UlSsC/pHk8OJO5aC2fyEPfb83ap3to
0uN32voB0m0hrHdTOMwZWynUlHgsBcIM6j+jzZfFO0mXYkFIdHCOZsIanP9B9YFk
l4DGCe1tZXFn4Fdc6/2uHS+/+UtI81nOUlWzWM7/Abm9UXTW4kcs8z/lYS7t+9t3
3FcpPA+/DpXAo/i9Hx4arHR1QzBaavo3Oez0dfpCzQZN2H+pCkabUqkdJgqCwrEv
JzxAlAmBy6neG8f2Rm1ElHTmd9cWc03642OewHmMm2erWw+4xOKsKdYf+Oc/d0Cz
tob24V9zBjx5Gfd/cgeEE6vAxl0iOgBJTMpZKaILlS2c/Hg62FI3ALmUd1E/G7E7
Y68NnrnpeiWQEVlQeGbVhPxkBiLBST7Vj87ix1iGOwUOyEzvEs/nbEVA2KIk1lxo
Xnh0KZO6GvnyN+p4/2qDos8V3OM2AMzabEL/cDqR1HwtMB+9l8rwaUjsZg8mwULZ
9BtqajTewlJUyNKn6eC7YmFRtrikrck6cWdyl6G3Dp32lr2aDqLXSzfRoYMr76r6
Tc+yX0TNfKE9aHIC19RIsiNuqqGw8gw+vLgXtN6N60E2w8YsVZewUGwIgyO8E04C
ct8o4FVfroh1smJ8Ya+kXOF6E2aFm6DjdQugLZEm6rfRSJm3bOZoeMuY+b6fhQye
SvIo7AF1Iri7ap4IQeWNOQ9wObNm4sFcLnxLmOC8LViA03PK1WlzDRYI5uycF0ET
86Fw0PluNFKk3OsoMxJsS4J5sZqgCg80xzsStsHLJYxTNTcIK9Es+g53NNkqsJ/s
rqJs8xePIFp1Pb650o0KEe1FJO5Oi19Y+xsNp2zbU4K7nLGGtwhLUDzs8V/rcJsP
NJtGfbk2bs7Zw0YVgXoSFrgZmf3elerNlakS1tVESbnMAh/r5z0ZIHEFf156c0vl
vwZ1Fwn9nz+B7QhyHZS58eJoB+ssA+DGWB9szKcVzMuoMLJYY/afKCTDFRApZXTX
ftVdepx7gi/Uf1hdALB2wehVQttVPEOgpAJp9YXkD/lh/CxPd2r3KzT7gdW/ouHs
jdlqm4tHmhANUbBHO9k7rxIXmyB9YT8dLyY+xUcVHMO8WIlesxVEp5D9jxqKx/2c
XhuiaWAqh6Wjq6i5MYPdyd13Mj7j7mWi6qkhXOUc6e5y29dwHemB9UcNPBtUbc+9
iuC0TNY9c9a3a/kKPtWmaO2YNHOFkbf0+QpBAF5kPj87KOe9KUTt5veSE7PRd4Zs
8wfXMJp/IuDjqMmZyUZ6yKUa9q8iRaTAd80Wiga2/To9YY5fyjGOeXfuiuJvYcEp
eG0hAxvrlQ83aHZ22luOqadFJmcSBFnTLz1QxnQNNNLHL/a1iH4vRS5V8fYlI2mY
hdzsAqOt7KIBrJa1xMqMFD0oDiIrNB4q9KCgCI3VgnGZuDpBJEmtQxvrGeukIcLU
veKg5jAx3yN6xdsH8ne7w3ARHbXYxzP+VKTNdKRCay+TrckRnX8Im8033mZQ6ZpP
iJV5y0+0NLyXj14Oh49WEyRnOHilOynGich7jhX2E1vueMHdnQUYosJteWJYEs1J
oCDgJXDHlQ6IAvIK0cr4daOffl6alrPEPjfKDd02rpCotgaz3fKzafpLaxFCkP38
f9SXukEfKuPUDSTXgadfZNtzBiI4GHGIlEFFUg2MwAuMfhxAXK/iVYCMej/I/dbm
2gOZDN2PZy3kZ+Z/DpyBLMqOnI9RtNHY7WXZ8bCF+sa7Io4O8WAOeT3F3UlVhdPg
9xiyi9Z4jOTBL4fDROu1u+VPngNPCHvnUrmgtP6EcfhfpeVJsFOpl9o/8eC+EbaZ
PpRqFOrbZ6S6gtfShZrDpUgzDctWqQB9+Z6Jy2/1nIry4JwYwL7iES292YUpsQtJ
HOuiqgbd3SERCMMloCLNMB+TVqvbudguWjSiOcxV98qSvgqqN2G8CEffDgu4x/zy
PYqE8dSMqKzxO8YBIbCOYtSujorLtEj7mdG6Yn61Q73fefonRFv8xEHrh3cxpMxd
c5mmtObTg2VQDccbhITStjia/UifGYjQapaSjTqe4xqBNWTikD0Xr7DwOXyXntoS
mcRvrYk3syubZiH5VPUlD6rAlUKnQvK0aFbjqBaRMrK6HJFYln5WhsXiSCP+iQLy
33H8D3v4mm3efHv9hn1k7H5a9rDi9QVYR48ehKaS/5izhKL6Fwvr8bdKC3QkV0cT
2W6C5P7NyhrmW6dIlvVIutLVlW4Yk40y3nAC5v6yJ/SyNrfmKzFLvEa+w+SGwaUa
KcOagS63fuI9yHK5Eldhr3XAkT43Ru9L2S1c6jhh/M+WG1CRrXF+oF5jGtm5K1hF
a6v60yTyGUB+pdVmaSwvGVh38gTNA3+gx8aK59683+GJh/nS0cqAyNvfPVqz6LLy
VAVKzsUA66otxY0hXnrba+ZF1SVOM1ZgiDVmFbWcs2zoT+DKAYJ/5YlQaVs2er1f
hrPwkEVwi+SkKMwfHh11ss8R76qySilQ4JQO50nFmRKqb+KxbgQRbEdm9JW4YRn3
a/Z1bU5ATTmTakhUkfnHlrpGeCRQ3phN7UWUQxuX/+zk/Qm0bwneZSR5pWjvDzuA
TFvzVvcaHI/qLc3+9ur+NLcO4CpZ2dXwr81Jq+9fOgOpsdduviu7i2MBUIuW2UaP
U5htpMPSXN8l5VymRvlnnRGyTsHV22C6sRpqtddPP5OWSY+XyUF1AhgY0ksy8UKo
DCdPJWviBnWQQElM9GaKvpDXUt+UClnNJMWPDvrWl2U3inGJX5gTccP/giR/uxQ+
v9hrzH7ke2GREo1VK8BMg9xUDfVR2MBN/SVZr9QNodBK8rMIF2agq2ecC6FSTR/v
cwwJ2LcXgoVyPQLhn0wHpGK/6laZpYjLkrZU5XncFwIBKU3X0A77BEGqxlV/7FhQ
e3RyTMSrkHyWU3b64+OFgqHx0Qcb8gveq9v/jOcSLoUKFB1gxLNzKhbgaCp522JW
CorrtLyc4fuJQSsxTKiLSAtRUSZg5wgUrWzXfkCtNlabqVgB87HvAYqr5PKR/XGj
gZmjJeBFxVR0urq4Zyes6OqAISw4ljIxVgVZtxWcDAJcdBQY7ezfzOtHN64kZ0HQ
f7svplHcCkM2LLj7rtTlzHMx5EAt5iuS+rZD/JKlHXBU+yVheY2bS/90frQ/wCo4
16Zk7uEEC8nrqwe/UzWM1Px7MpYP+MEb/V1NC+iJK1vEmB7Hb/3MsEzhmHodsdeS
Z2P1oVR9nPhNHYUE4I3rqiM87E3kD6Ai/KJFR5Ozt+zfEOiHlIxD23JMNIET/UUj
7z7eskTmOpbRilk2xyiIiDmkVxZAMkygFVSbRkiNoBD7RT5xyWBcszMfJSoMRALF
gscz0JxJSaiP6v6lRtEBDhatSzDWTj2oFY/dyeOv3gWxh8ZI7i399dbhIs9m4N2J
YB+sbvQ068CISZmalt+tKsJD7BEyzwo+RLVCY1yOM5wCSr+wY9vqVHm/THQUjdNo
RmGYFpgK3M9SBYEbWEGIdSfV3Ko5bDwGgQYW9h3oRBYYccclYjJtkOhzRSblMz1+
EWgGoMk4IhGWKKTc441+iPTq2etd0QwQe9Q2FmuzrcttgLHOMkxNEp4sbvpdIyot
spyoRG4GV0QRZZ5wKN3zDpOn9V+wZYP4+g6L1Lcg0smDEzs+kFamPDP3VUdIt1jz
24+xwGiHdIbgOCn5dRKWoTdVdh1B53Q+92TYbBJw5rH6Xh8qCbp0WtqFM8gctIeC
KYLGOmCC04BZYLAvmmO0wcjZfp6d6s0CxIJi2EM/J5UNinVDlA8uUd8LWJVJXhjx
y6IRpXBhU6dnPE2hJuOcUhhS3VkmVOQODcFW/f2EeG+8kmCfqaZThp3zDaGNSWuP
DJW3FcyMaEgcnjd3Qo+gB2bhFWI4htHXVJ8AJPzpvXWLJlJ02/fpcKMFw1v3dz4q
z7wsAwjtSDRtj3CiOOry2oj2xAmlcnglgN5XzjUhpmjpH/yCWP9z4U3ICVr4WSa1
thx8Y6KeVXUOKkTvOTgqZX8YFhRKMlNhlBpKwBoMlJfYtNc3R0ZQ1r7Pgj4IRcbT
h1SFGwB9SzH9nFFRqOgKhK6mBukwzXsE2dFZoqonSPMAN/H4iYjwlEp4RYy/RWIQ
2h1KHoSv0N+e7iPCCD/fhmWHV34UdSbv0Zus5vsw3ZVKvQC3rIJJQqKUgpObu/p+
Hy5sOyR49JTA9hJVwYfd4F9+LxdT6ciYk+PEwc0fF/TdwoB37Znoqb1uJb70RraT
weMBiX3zIYdeOOy1qLHU8YcHVL3AE3aZUaHmYUZ93JZHwmgO36ufDP7pyPFELzK+
1j/OgEwrlBGhMOPas3++xUmtdluQafG8ToBjsyTosCFBkitkiiUEjvbTcKiO1RWd
AtURzTwljmt4rO30G/UjAo8kG3TdZBorSNQ2k4cTMnLZ6TtFTAIPuY2xni4BmCr/
btSIQDzSgRPwna85Ep1rA/bo+J71K5dLY7kqHu6/PmHgIYHJd1nBvs23sK8vmT1u
dOfXpvya4vARSHCRXyknWhQKBkG6F8aRz6xhx7fjDCwWBhiN58yoqoVAmNMImMWx
TPU0fORR6ahrRA5WgMEofnEXwu/RyV2f3P9+4iwC4Q+DnAdQPz+gsZK6OdROlzAz
LCg+QkKmdASiTBhg54OSTIpgSF8ssBRzr2MammllhYiBE6hljtKt4RY0oNhwnkB2
bVmwMYxs1yXqlCSr9yJD1pGK3tPTEFVgb5B2CZ85P42t9ylO1xEJu2pF9jHKODZ1
M0XXEaLKGRI9PnryYx+JYFA+B1P4hiS8H7w0CKGR0ker5vSFPWJ/ppbj0a6bR0Om
bdtoc35jhXKDkVLeXWVyQiOCDdngKdwH4ccVY6j+T6Jap1SxkB3XseQZCiGhzZb+
MaNSB7AeIwFaePvwTEsnWUWDAToXOB57DswLZiMIWZrO0PEWG38v8ZuA9aFxO2Rs
h9kCV+m++WuDuJ39r5deZiI67XbjCBhgnMDebB7tsSzx0T3b5/kbxNJYG4TIOge4
+lIsHkuzlNVU6lzSBByDZlhuH3b6JkE4wwMdK/BScrZatKLykiJbk5tDIVqMEvg/
QLcqFbrKq2MYtRLC8+dI989SdP4Nki6sJV09tOBkjxTbBHHF7R4LeoMbd07K+7HC
te0iPlAYGx3ZxDhSoL25cwu0zNCI/MbRDGZm90O/ldcYdU/5tAP9hXiXa+9TfSAl
5r5CpBB0IdBmzhXIlDrH2l2yPAKiZTEMhV2lg60o5I9MHwzIkbBJTWkSaJUVncmP
2tZk4Xe2LXA04485inp+z+LoKQXBdfezf7XgjgoJntTK0RQF754bREMUURdogfC9
a+G6CgDSxMh4f4m/PVGEmGVXWnG9gDwVdJ2pzm6H/DQDKU4FXHnx7jYjteOGDSfm
cb/hxtOZSbkUTFF7Fz2NWfUBgslYxRscofTmPXkclbGcsYLuo56aWB98z7UIjHCl
rvRs+k+jc+nSXgnNZC5QnMfZfTzSUBhkcO9oXE5zrlQVqwSkGfrgYOkFkdDY0eCu
5bSOU5zj3hSX+WOlT7dD8VqnBmi5SN53q2ImoWDx29QTmMUI4q88cJHNb/QJZuE8
xqwgGOV4/QAghAgeFMG92fAGh7eRM6Aip/PJXY+EI+Z7Zr6jF/FLZT6nh1CLTYY/
kNiK762c5zY7mu120QcEl8DTxgSpaBgHeiq1Mqu3zKXB7urE3IdWQkDm3jnV/rwO
MP0FGSX3UbsMCGXbSZuO4ClYcgYxc52zA7FSWUnv13iTOoGCFAm3kdP4RFxLaN2L
BGshYM9t47nKcSGIoRuGewxECIg84sdgXAacDDuq3W78/Vy7zn122R7D3bEnaslB
PgSovWru2RuRfPOIVAXoASpRfgwy6pUOZNcIAVUD6qmWF0jvibFrSKwh6Q1dCpS9
CKuEB+0MqftRBqTFD/D8wF9b6RJNwQ2aaMn9H+i/Ud0yhVXXKBmW96dmyITmkY+Y
Jfj24Lz9NJkA4+n76wfFEvT1msAtbPvxHIwNYnvq9km9hmD7ALnVmwBtOYCuxBzK
ceGBcHvDARbFAHKFR2v1Hp12jsBWUXF1vX833Kvx8HV1BhrnL9+koQrHc1ry8vU8
TOonwhGsiWRNqfhV1H3eG/Ts9ulzHWiLkW9G8aI76lvYo6cCJ28CSl0pvbYi2lAp
km3AENGGvB2Sk/ZQpIKKlEFPjEMhSvIpCyBfpYuXsB5HcJLf5Hqc3dqmBkWBcM7c
3QXVHcYyECC+NoRBlYRYfrRb6pO2QSyF7f3n8pBUPR/3Ol1kXSZD8aBeeXpqI2Kr
kaS1QDN2VHZqyHqF0pN3tBErAl9afzxZvPhg6JgEJ+uvEZHJtrRVD1WzndpXD5fU
jBuo8dcZ20YIECHrdJBn58AOl06PhT8R59IZYZ3zYG9p9iLB24Du3Kfr7FGlgjF6
DQUCmDvJlnmegYvvMHfZ+T47pZpwuU71FrIVaezXXtHebC/Ug0LhI+wDFVqjYcdz
DtxQT7VM11VYHXjw/MoBSX8pM4OeJj6quKuLEVJAk6VKBwVXgZPhourO3F0IeUpW
sIFicV0SkxqRHfbQrpo5vJ0zN7V5BipXTKnodKpoR02W7ef89llvfVowua0ZXbMw
hzYAOZjIVY3B0nJn4i9f7Qk+puMccnTIV7m/nuwto14JN6f7XSyolz+tlSudbfQP
A7CYugMncFy2Msoi+M3jLwU1jnkfnkTG0ZFfgV3prcMOWUa7aW9rtk0sPvdzPh1/
zCT2JK/vcmn5q9fjyD1rMb8xhSGZQX2PvNvKenUvYNt5zA20jP/HVgHCYL27eNSA
QwgvML/BSCiZ7hoGmjNFHU7C0qX7AtyYkxNReXySEDccu72v2FXl4wQ6WCwUpFO4
pkCSrUm5YBZsNqKCqFAdGrEfDKkP7WgffTTw7R7Fl20a8RiD5ihWD+AKsIYEKhDU
G71dR4dMyyXwnslYSI6Bz4m2/YhGIHbftd3zvqP0jrJmofr1kcjXlMswB95M+QsR
xL6/Vv9t2xcy6mvSAKQI77VOji8BBbZNm+ywM/OgWEXQa/qeCEoEVSv+mCDda2rW
iNWcoa4PMazEbUbT9sbRIViMk9+W2GZg1fN8lbUGKXLOPG2H2QGgZNkIQBphtA9n
wCnp9sM27xvv3yoFOSCldr/esmAMK9d5H0HAR2u28M8bIqFO1PEaygwgyAoeyR0a
BBlYLHW9BFyzROcT8cV7KsCsQoF5TgGR+vj4u50PLAJl08XR9y9EC2q0hq5AJSaX
Zp7XVoLi5DNbFyQGr85v8LsL+UXsLOCfhkhbLYBSm9v/w+PRCKxzsZRNu/xEmrW4
XD8/QSDTdk12t3Y10a22VR2lVtysE8BzRsmV0rBcPODVAXUkaH3KHP95r4Aw2uDQ
ceSPTNuknuZo9rfHvQ7sL4cgFPB5geQw6+QM10bKnqKKW4cB+QvbA5vdWpjhZpAm
A1JYd3tbV27x2AIGX0CKgsrnGlhXvAnhAeU7A3FMgyJDPCPCNNoorZzX7W9slV34
WWTY6AtWQDHI/tqOp6MpJV9+OuYX2cqF2TzajDs+ohSwBJSdxJ5UsB1nhHv+TE2S
5W9N0vv1xCQCjRHXGofmePlsfEmqu0wf41wEz0L92seXGDkSom3IOD9jG+9SXKql
+G1GJ0L3hv3NyAx4Mkkrtq6AhXnS2jOp/qfgAWX0JlcbgtO+yj8BFx3yV07PG85W
MJae/PZgqx+ZaxtWwfVGIrHoTkeU7o0NdJcIlSjfem8+BPkZEosue1yS1Pg0ltSa
NlFd4I9RRF6N4xw95olF/m7PbMpsCXCOlxUclZJOErI7Fa7riqOS317vTwHeDrDk
xDblIWxg84/7LEMuE73xONglUOgzbZzC5LNpQTqS88meND3NcFVWI7XSXjGEH9mo
BIOqFFjXlCD8SMCj3xHJ5Yve0A6vzYHQfJyquDOyhonKRNDGzE7njbD2kh4YorXy
wIK8FpKHyveb3pNe3hD+VQUKf5VyV1pTqGPpu/lxFwUqYEidgjaB0K8R4apkAEiB
0Q1j5Ln+P2Kg1BGBYnnTNcuUQR/9ORxG3JpblIuzGWNl0hkCdnvu2jEhxPnDX7iU
AGXwOPt5iFYfEPmfBu3KlDvrlQfIxBZJYsB/1w+p1FYQEMlD+l2HNdTCdmZO09Nj
Z1eIHz45Qm7DvpIoTIKAIOnkBjYRpZyY0SOQbDvURddCwfBLuBHVQEwTxGZeqIZm
WVYsUfF6kNIYTe+q7pTxDDpB1oIvqiqItRk4BcnKTQXjWrm8b55u4u0Qzjhmt/0/
811ZfkZ2MIAmLWEzre4h8rHXpjjrOFOhc3WKlCpanvoMMcJH0pkZAfImEikgPbns
kUiMrqS+L7OKzKoS7ko91gMQwcm0X7U5s0UsuhoEIaFRwMTBbOSMoz2wmC49yXHj
znimmPKA8IyIYrwV++PGXAaxRWOQt6ws7gfyclcK8vFAQb9nPpT7TZNE/81cXk8Y
sGbLNbwSHh5T52gpxhW+GhislUrzm8Tk+jdjpwx/Jnd+raVwC9n8mQgotegyJYZF
X+7NvcfAa1bcyH628g2hok7AsnFtfLu7UQroXfXnTR+XzStTvIgMCHTqPv2MSOkA
UgWDhezlOl6yJwcm2/K2OTFcebhJ6CsmnKzXppBCRH3QaxRhORF5MQqd6V7eqHs5
J+6z3PmmOgm1tcXSuRETzL/DgiyZG+7iorRTqQ2Y7AVkdurv9ZlZ+3WXq5TGVHqF
ecDS52fUdd/B5FFHHJFZ/y4N8AXIQkjK6aFGHAIWqWXNJbWhCbvxsv8rxFIC2YJ+
jl9J9nonKpYXcobybG1Kw5XTh2nMJ3FDtDUKagMa4INEkmdxOPKzzWrN7w+n9ctK
MgCF+7wJp2D1B/QvT1nJLuoeZpz6gt66Iu0/1AKtcmzgd+vCcfc0EZn5NQqim91i
nEbGSYfLSWTVkEs1ZBMuVoSdKjo3GgcuL6eWM7rB5Kgay4Q0P/IXQmA81TOK1AZh
9hIYyTOGNNaAeT6FKkjs+cN3slhXH3Hv/GH+6cdeoPzgglDaHIYBBpER/sJM3YiF
VA21V378HMCDKiDSFhIncxHdn0GQ7nZNk3dgeHizg60YuqsmZhcs/dfYaEQ6fBpB
3DItiBZoTH/IcuVp5L5XVGiQZ4Z2IIantpKByGJKSTWA7tbUIujs7aI2P8H334zv
3d+XDTX1kzevP6kRl7iDcOiUB4hD+j9zPx2eevkT4OtSKp3tvmPQU8seb+Vqr0pS
KzXBKaaTCFM0KfW01KYWlh3MOzlR74NanTYK5GuHyx3ElvDrZ7ZeTpBOXkqeqr2A
sL5B2R0VOBmwubD8tn93lOk3xLXSqpOEJ+4hswdsYh6xHhfqCmldlwf0WbaEWFE9
oUYh5HxBrfygTCaQWIDZ6h3k133YTqPoKhQaxVpX3tUF6sI88Vmn2kD6xjkM/eqP
/EuL0I7tdgI7VAlFlkp3U+iv89ix/hlNUH3s1IyQGkZQPvC1flOV5ujfNPKDtRS3
XmTLsbXNRszi/+IgTSQ4wQ3s0aUpyW9sWHXMp1+BbrwkIIS7OPyawZAVnExM2M2a
GNePWyv0fJPWeEJ3y6PeeciX4ech6NTpg8E2opxA+6CArcb/MVVeSdBGCa6DC5qA
4ABE/dTtUUooVRcP1fEd6I6oT9ui8wTCFzVeh1zb3d+D3tJP/TzrjGX0PqnwzN74
grG4XxqP9tX+tV8fMfNkfth4qHbUpDmaX383Pj1QMQR5z6Yg0eDJCM3dz1QycLXX
w+42l9PupYUWNOmW0PAtwVdLvq0tFyz46W1XC64z7SDyDhyrgmh/LqHTBwknFUiB
h+X+BZIEkf6YG7vfW1LUkam4doV211rOZ2y6WM+TepGd3wrcsKXnmtxMQWjbuFha
D2qaKiPbaeCERC2e74HoUZcbLenM2/0C5jdE/58OJPTcp06D+InMa/4SN8cdv/p4
QeUce5TQQfA3td3Q9cLH95aYoSYyS2r8u1+pckCFoS3himtgQoR0xtZ43eMELJYW
wPrq2wus4PtPriF1erA+JkvNQUXb3AQJEEL+RXbvZG4v5SsCq0ULXibXK95rA338
8VYp3HB+09/OhY/LB5bMKBZ3gH0HoSCTpRBmALXo8isUqNX35dNk71rdc+sBSuyT
IC7/n3+N/hVV2jMsDgjHXIoYHg8rmEjPy8ptheveWLx7NOQXiJXg4mPDJV3zcRt3
kYQK3SRyIfATxkON1KOmB0PcpXtQpvT2l8gA6cqQAvK+qF4cBGoAprIRpm+AfB8p
jK+dRanCo1v2G+dH+rd0ZgE3OlPkScvqRpOeoYCtE5McPuOnK0B4nRVjk4OmBjhW
V9eQgqc5cSfarHke5tsANp4ASCJUdgc7TwWRM5/TFguXAt/+RHLDSV6w2Yv+XJJY
dk1fyPhmhP8NtenIR+cdjt/UIu0hZUnon74/BC8UyqFFWkEsZa0Tw2yNAiQKjjmM
8VzArNjBXY1nyOY6c8pEqj1i/zAWITt1BYJkEBS+F0bqMMt3p+F/6Zm2r9BcCJL0
xu7K5a0JqXBLUJYY2Py8oBhVdaUxOdfcyzaqLmQ7oUzPxGB5Og4Vtw0zapA8oh0t
Rxf+4+ZM6UBaIjlU+ZdxMFLQ86bLg0DMCFgDbe6qpOP3Fg7d9wg2tGL87lSSUJA8
zBfQZM0SMe/j6yhS3gsdNhfeRtgNgBLMf8GZW+9JkU7AUm929ez9tDAqXkLjFMc4
DMIOJKi/Xg0ZT6GEoX4/jbjqAUCGv7lL3t691cTT6lTf5JARXX4nHELQJ35GbVmh
dK2d8ay9olsEEYw0+4aA6xd91pzI7aCU1NW0e8Xg9xcYRmPOu4gsxoMMrze4N5LM
wWdWcqE7HTcLnvN6nt3gPrEby7619iARS7GUpofYEu34zli0syyJR8+Lr0cfensm
ZiOaIrYNgJ0mqY00HAPCVyqcvxCTFC/slKiFv6TdggCxCknxvJ/9CCPKEl9F0UhJ
/D5vM3ZmfMWO6wP2LjJXBQAi9yeytHm/rKWk8QtKnQxT+/BzdtvuAEp6F+OJToYf
ZzipF4nsHC8M9+PLZVDbrN1VLnidQ2cZ3HgPz/MVanHhV36Nv7JaouxHrERztHUT
hqt+9KGocUeMTwwoDXMZm0xi1aGcrgOzv02BqXMarKhRsYhBzjSy558RCRVerEWE
9RDTQkvWHtv8Wzc5KRyIkIXLM1P5XK9Gkh9w3h9lHsZcf9YQZqZx2AWx/8kOAn1s
8KUEUvk01TfqxdbaaON4qYDzWYJMd7yOWzsl3gdviUqAqUC6kNm+gayE2U1pXL9L
+UaMUwTVxTEd87bkHJ0BgNIww8uc+cXBb0a5ipYeMlgXu/IHzXAykDLJqxbJTavV
ObuGYqPLHyabdbgQztBA0Xk+1cw/FR+F28CYVCFDGiboWPl2AhkCle7tZ2JCBvns
9ciA6dh978JMUqpQkAEy3BMRt1uAEF7OuaES+0r6TQ5jI+M55/zewd63mz/HY98B
IzyW9bJB9W3owo8cqNkXLibfN8szl90o8cb0C2K1VOudko0t/E0MeErGkeqKnugg
2Ac9X+mYAPkq5uZ8CGcRj9D/ThazbF9P1WwaQGiBYEJ9FYnVmAO7QHwD5zSgBDiE
wmtkablFExirMQoOtX3JQ7ef+EGRTn9MuHRqMreJ7PwszZYd0qNiwix/dEkFSUDn
35ej4z3FxTuVSNzmRsITRHJVnkwPYNIgPighA9TeXyLQCq5VfpyZzTJBGf2VKFM7
gtkvKmjZ7pR2JLaDNK4TTwef02qMV3kfs4a1YuPT3q0P/I15r08WRXjRI8K316r3
x5/ogt9lQwrNB4GlTEqT3na3K29mnLRBXj/105P8CneMaPE2MdtiHX9SS3SZzeXv
v5nilTojd3i1c935vYn0h84k0CfU4rTrJmoBw9q6bw+UA6xfpuZdU3tKDM/DlPgp
v3bJYhzQGVyJmq6ishdjybWVeOTqzaIan2nAvIcp+xB1N2SbdVfBoQyg+rUBvJDV
YE1Na1+hMZ3pzRorKc+Q20cYr4q5fyum/STgPO1C6KWlaHwPaWbDiaglKDzOidAd
XiOcA+IKE7Ek6Y9MAS4SU5mNJdUPW45FKIuqE/PwNPBwHyrNrIHnqkzFrNIicnZT
7mPa2TDlyh9Jt5Sdl0PX71bkBA39CN07NOZrBV1VVCbXwimKna4y/roSP33Lix+f
HmS7IfxYRDtwhXsuA+we4Ccg48/Xc0VkzTO+Y6uF5qV1QG97FtIXBstZ4oorDlEY
i1k/qCbOYfZWpLOXcZ7R52c9j3ynys3k4I5sWD43+MGkMtzMPbqvSozXMNgZIPFt
dcaHUGlgqGGaaFfzg9QMTIdZyFvcohuEPczx2d9nOeguLvka9CvKFmE0zLLLV2yK
yIIWZ3HqYm9+bNwvbJtQjGeRG+9TJwxfsCJCHXZ5OPx0dnRg3Z3KJP7NJ58MNL9J
VoV8tKrJ5Tm5aanzzh5CTFIWLOEPqXbOm/4MfpxeAyaXFK05UkYWtzeDf/qQxTzi
+yenm8QqnOm+yc6QmyVH7845y+iDK24fMphP17wnI6KFopJrKyjzG44gU5n5woSF
nZSiwr8kTXtPYgV3S9i/qFZUHNv6gkYy3pybcZubTwLQEaspiCViCtoqXvpV6abO
Oui5Ohjzx2cdN0jmMX5Rq+GSSCQc3PiDvO+LfDCZakQtXjBybVd5OrBGwXBjyuF2
3RXfq3hBW+AEMfw+eNyqaINuVXh7ECFSK1saGAAHZRcaKAO4d6y6Gs/Oe5Ku2z1P
BRWPagalzf6uhwEaJD41+WuAXGp8afGqC6/hmZ0QsntIePo/TPNUZuK6A1IeyTN3
91THa4TPTbCsmg1S5qZPyc0i4KSXjl2T64NCGcPIQoQyEPiNtuKYqe78WD7+Rvkq
M99yzqhQ0mL/aJ7Tg3seNHN3i2k7rHi23Nj/IDuNn1J7hvmRTssiM9rzqbsPeHWe
uTIGw90da+nDUT6juVQv/hkyngIQ3STl80cyKOXfAyTK2nGBZNe3PHWWLfS7dEBY
yFfzEq5iHVfZkixYejtCLFYoUmJ0YlAKX8T8tz3j9MmAR5AlsXnAVSo7EggqOwls
gSj6luWzSGwdgVEWWsYij1ZUSYgML+OCsw8gcBPzjMCr8bDtMgW4fHr00mKt6eRL
oao253FBs9LjmdKkr9LL8Y2I3OejEPkXVD2R7kXd6tPJgq9yvRhvDOlOGSyLQgQh
lDw/nxFPxqe0LSeRMN102HjqfWCUqAOJCpBAKliWZQvdpPXT6XI46OCSoyldbcMn
yTN0kHSQYeuMtu6SpK8fGq/aBiR2HBZDi1NKSFcSAT2IgYXyuQepbMnl3YA1tvVE
kWXf/26EHsS0uLeB2947tJu0pF5OAeSZ/KdBa4lzqEirVf7oxn8gVsqg4qNIErWl
5zV/Ix7YZzHDE8P0o57s4xovzLKqrsMgbQ/fCHSUJxdLi6Y4geennadnAQ2IfCDz
MF1oerpLqUXyW0i5jfXLMAGz4EZV3msgW50OtyYhfYckp9ktd7Amo9gGyQ1P/hbL
/3+WCHZdksHz2JyuVDVIqFJgFk7I+3LN/rCi6tQLnDyNlcG9aDACIQhlB3rQtdIC
hv13pkVLpgsecxmHJdQbeq2NOIJYOm4KHkDWOoHlIRaguhh3eE07CFx8N7Tydr9e
bwaVG52p57+3CIgMDaCbSQt/sdzl7WeoTfXwH0WltlVw+lBqBkVlru+htFeztooT
ZrKKCFlntr11JEQKDcpslXB2ZxlqkgdpOG8O9UmD4bucZ79jpvTpSYO3L5N1fpiw
l5EWNjuWYRRlbI1ermm3JW3qNlKE8Zd5B0M1pSNswLwmP5LJssGVB4nqbueDVEDq
czvAe/+qxSfUmQbO8OWOr6Ojf74r/uizhYtAg3CSmjhXKZcsYOLCVo5LySVPRYxf
wC+hTYaPqd3P04GBMGF/XydD+w9p0ohjlzWffuDLn81xI2jqiArcILtFh0RSIryW
9WaGSA27UQl8X84T9PXOV/4nAMe7iirOYfEIOJk18Gy+thjOCIBKDm2mOh1OVoXF
yohJM2wEgNxYd1yPAA3Pxmlu2z+J6VQo0K84jdXZJC7/HYx8iSQ0zTnuwTUT77qG
/qi1EGq2sG0tqbkG+lZOR2IL+eJi0omz4XvwYyhDQLiveMHD9bQjrNsaHDovuKbZ
1Wt6H3jwSa90yhZTIDY+0wX3d1OoiCow8U6E/H5sxozD91cH9H2rmGsPgacP6hzF
fbj8WgrD6NVFuU9fcoM9XYmb/aP7e9g+uRxh+AKZzNfA/SBKa/cTJUV8KHEZnDX6
hGONwaHtCrd/GyBfumwSNpCNcI9EwVtCfKlSoF2DfkfTdk3ET9kGukFokytgASJm
bXNUBtjOcLmMYLWMcQJ1YYR1yAp7EXlDDrwzOPQlgnV6GODyl4SjVD+oGLQdibSD
4CC+LAWCupkp8lu0Do/5Pr0XB+u1jZIqwSeUwa88ymuYjyGl+C5YSVoVfEy2Yqpc
r63rpkp4cmxq7EvFlFZQdKIfRZguvOHyiIU1Jevkld21pCvE8KDtfyYzEa6SKRXL
G96U8+W55aHdgjY89e5mifavOji6wm12n3OESdb5f74tYB5v10+1MvNGh8xX/zKD
4NOQK+uc5Kph246g1+LxG/BsYDlxWeyCZ+VJdn1ji3+IZ9RP/Mh6DgMtmsWmE292
w9QsCoo7nBBVuXr7/i6DnnrGeMzlmsE8jQVhgafP4wZ5FCRWoHRNCPsqS3/AUTiK
s1/ZbzjWgCGXsEUBBiH1HbNH7FfiJ5YS7fU6SAKFf/M//c0sFHwI+cqFMWYBUS0j
IHyGlwgFjkLjYEAvbVUtL/bHyFxApPAtnwIpqgMVgHvhKIOLjtOZtWkcKQmicHqr
Re5I4drt0C7fBh1BqPo4z9aJVsDEbcrvRUdaeUuZpEvyf7mcgpwlb9PGYS8ZFIz6
wQO1milEZDAZkmBlaLCu7wTW+lBtyJCjRsUs5PU4SlwRQFbKH0GdjYLPodhC2d/R
I5jUYWMuCpWPWhdDQ+axCrTQDC89iL6XMoGbA9cAKNmzuzgl4wQlYIQkt28Aalvs
sIIdqWiRO+gSTF/b42ncEdBOb431/Bl/SWALO2GATQoruaIUsFE2+X/Cr3Dq9SWC
sX7DGuMNbu9KrlORRg3gxMyZxgGE+pjLrYJWgXZJH+Ku8lge4Jpv+13OCFGcjpDA
t5PJWVY6v9dWVzK1Xk7LfE2+bKbyc6DHyJXCn6UpMY3Htn2p3qYJHV0bFS0jUtvy
ZikgYPx3arogZbizYQ9BBiTAFRjC3FJ83v4a02DgOYmP6NXJGonzkP0yJZ4+t64h
StC9rzDWD82yUpHNAGaZ7SDH/9R7vj38G+JXenqBzrgAq5sXS0RSAugtdNrAzaxH
j7b0rtXCusUaBkzPOysHyIhUJCjIHh+CxHb+lbAMafW9rnePQ8Z8vJvOCiaPuE9g
x6z1ntLioMO3CbyAPUpr/qU7iIX91YG+XjzeJznR1RBZbXKvNenHBjGW+Wk3u3LS
EKngTrW27JlzNjIvC8G2tFYxJJMWg8UQ5IEZvmYrWpDhlTnk8ctoS9yKpo7061Jr
+RRc2pV23/x4wogwHdH3WovsM3o5pcaREcgs5AbUB5/dl1zIBDECy/5TQLVZTpi/
TR3xKsbNifD3SccRDIGuX4/c4kQNRkfe5UNQlbq6SCUE9YK+1Hdqa3Gqv8HO+ArH
wMGLfm6Byg/Y4RYvVr2BngtdViNTr8OklMH/XVAM0TR361HVZgJR5NTJT9wdawJ0
dYTWbRr9cA7vh+x6mMfrPwBEVpstmTnhvbbbeygdfFs1pjGUPdiUNt1cQ32DbGbH
N2+immnwf0uUuFBW9XQv6hopl8a0OJmwJ0Pa+/UBtdfKM/m/WiokSYGrm0sr5Tip
/zOsZ8e5YwWV1PRwo+zUA7UrAU4YlxxJjvXmL97Vx/hM4IgVip/hKVOfy+oFUOSf
uNJ+4dYAVaVuRk8yJxHajQKmsd3M4ddaVsrfVMEseK3ZJDVgYShRV2gLXVqUyJxj
ljHr54250MAxbaVCbRuvcsj1/08HSWhbGobDR8QGLxP51O7fg/Wh1yK9ZhwmiQEw
pTF/Qv/j6bI61HxqLo4TPN+njFV1GEJO35I2ta7IVga5fCorgDzjH4sauwoVVteE
UhxIDy3VurJFeJ/Gl9PnT+23dK6PIeTbBJksSrOTTwkOVTg1yiLwULBElu8xEsxf
LVceu8hLqg4wX6OB6VSHDlhAMcY3iSz9mkkBI671TkzF0WPwwoqZmaJRfi5ptY1N
qbFvH0lNER9dEBD+iC4+Bi4rCtlUp2+qZj2ZZWV5RX0FQd/UXRk9DJkwnDoAoKBY
redS6ihVFhRrrFEf/zgbD5jeVpTOH+7v+4uGKSYvPEZ/wyVXgzwp1INjI+gOfZoq
r0K3fp9siRIQe4mImLHUOV8cwy+dOg3J2L5gkxYgoXFPm/mMxEZj3AaO6qAxVfPU
zBqwjnEsRIr+mhwdhiFoPc0F9fO+DwvfRB4bA9jFPt7BGMaYANloL0hDWYVHQpFw
+rQU8mtquzvnuYsWG1GBEX7zlu1zVJrqncQv0Du/9jt1z3qF1/a3bT3GNwwNKyZQ
bw4qFrmGCrV07++u6WqpdyfWGoDDnexwX452WRAIVi2diawROBgvA7dnUw1bUPp9
9gOfJw22EfFfOXyLvZMzPSFtBOSQdBBPY0WN4Txa0+MZu56X94vlxoe1YVi1zAX8
jHObT/jvQMfqs+n9m3oedyg9XoEKDCEwScL7zrx3xYdbSzXpbLIIHpEnnuU4Z0rk
y4hWbH8p3P/vaODPRC4DqDITsyU53l/tl2PjZlZtClpV8r3n6djERdlOTTuII6rY
V4HiH/7r9oR7QDIv9wZFay6cx0mna4kzdBWVua5FXV33m+a9CB2pNRCwbLXmyimm
gGOXilUCD7W+dwNkNfdGhhi1jF6AmuawUY7/WN4u3if/cEQSx3j0XBYbzGi4ceIk
EW/58GY+RlaDvSEc4Oef3Hv1EwcZ2yy0LOb7XTh+rVqJRhiw87nvVsCovnkkqHwY
tvMCRzDiO6ZWbPz0m9PjgO7gldrOp4nsB+RedIRM2vbpj3MgaPKm/372LMD7IWIm
Izs31VlvgX3MNQtSe5H70TH7p7Pe4rhUCXcPOEmdABVXesWkXw5lXurhDKqmintf
ROJ6RJyc0OyGu7jy195kdVTSsSANp6DT7Kn8dnqgIOI05t2IPLURwgfLq+6EJ7ta
SYXBGzCz5avDMx0gaF4C+uXyncM2nTSaBosN26nLs0kq9R3NceO8O4e9IRpAOkr9
fGzfhZWZGE+WwngILRJ9AWLhZ7H9JHoBsgMOLFlMzkBNcu2KkXJYB31xWpydRq2B
i8gQjlL5NDXveXFQc74Pw49nTGZELd9pfX/5XjCK1rEdSIjDWgUny9/U5D+GcLIK
tfAabxntNZuDJl+Ek6NN+bYYXsVvqcMPUw68UCfCc4IBx9fqn2/RvLE0sUQt3wPt
srfIehVE89msXgUoWFLjF2RtLpJnf/sJmA80fnck/mT2nvUNQjYw0evF6g/IUYkW
E8502Tln1fOHsi0/t3xoCDcQXsnrE890OdkuY/kwxDhFQ7P7BbGMFpXXHeg9oZ2V
Hz4xqQxC+fdR3ejCQpXjbVeUOrj2Eu1nxOI2keF3ZseiQMq3GoaGx+o2OjvwmtqP
JVnOXJBSZ3eM2eAM0AEQDnBGken/byXLfObVOtCnEETpbIgMwvyamcgq7KOVQRr6
riY0zOQITQWkfUjxqplpH3O5+zS8hEFYQGNWFDp+WCRlNlANcGlLj+Ak1SrfSml6
VOMdqO8dwTm56vv0r1Y535CiSeLyUuoBk2lbgCATkJYQWisKAvIFpS3Sf92A+XZk
vhCxtmNHwpQFCFEHbTi+8BGd3ZAAg+HhwqX5ICabGKSlkkW6yhWmpNTrjB1j1YTh
/GgTHWu9qLDl5ZPB6H1eUBrdXvvXTjogZOzSaxtn5fHkKkz4BpTDgJlpxUwe9Zla
Z3SOzKu9BV9aMbRRvda+Ef9GYpNcDa0K6ttEp0W9niGtYBoIrHCKdCkNELLPZSqz
P/GmxqvjD3ZFwS9Mr0dsd84gHGSfVWlqdOn6IER87vXDV8MOGrFXfqmxZdi1C0/Q
aFeGUobwlDtaIaTE+tGTFE1ogwk8pPaFFqmLymFhohiXDqCUgfCmM/1zC3cidmWj
ckZMCcsk+snp3cL6XPQaR1GZ2B+lFN/CTb/dPhsb5XYWjocm2LwiZoAmslJsyE0C
86GWDbn4I5cFx0Oc+10Vdn0KzyL30cm6zCwHsJeqIgMZqm4kVlizHPTeX9ajrx+X
kZgeE53a1VOusyM5CDQAouOgKrAB59Jolic8Oo9XjCVoxUEISyBNcxjTMplnJqti
Ky1Bo+tiQd6si1FBGcApFufFB2/o54RrFmyfZK/Tg7zR3v/8LLm9gatZ1EUQUTv1
WqrziNf3277ikrDyg6RVIKcDqME3q6YRFkdGmXr0URQQMBPS64BpipSXiXdYfTkG
pSad+dh4+J/T9VFhzjR3P9S6aWtqO9qMpPE6OXwQlkXIEMFQ2ee2YGUqwDGzHmaC
peCuS2BBVFXA7WXyJ2mFFSSuUie3xw+nv6sEFfWIig4r5//kJ5WkVHUvZK+zJdjf
0b0FLnGN1QZjmCQFSf/LGP6E9efLXlc606uFl0gzJ75vSGAyYr9WBT7G3feuY3NG
vi7ZRcLY6cDDlo6gf0eH71YCspJF4PKnHYybOuv7WQGDxYlQ/Cd0/tuniQ7QZmS9
Ia86odvEIhLWBNcb+iwT0aBu6M59j2ZNI/xGGK5mZ0VVWO9iEbBd/oERBcKZklhl
TjZ+avwj0Y5hdcTGNRQ9BpQebsHtA8DN9oWIB57WiYga9XpHlRN0FojNquMqckk5
H88Ozrm1A6W2V7QPzgP4DJaUFdYtpohfgpGuiMdFerniJbNBJ/OtDGbHGud6NteB
H6hpCAH/aVfpwtwkbj4i3V8BQXgL10ecck5pomzWPF7YOgst4KO4KOM9SkHICJGy
muFj+wPfIBqvo5PxudvQrUGL4kHTMt8THALeTF/XpvB2nhHu0dlWUxC7FVOrxf5A
frZ0ZCv/bQQ7po0C6AD4SVUm7Zao7DG3eGn+IITOhsfQOoq0j27mCRM1IlzELY5T
IYAFc36ZaFYgns6XPCp5x5uZHOlABCBv9fto1VhE3aycGwKm1rfdYfvDrpzlFjOV
ONMrA1gPxPVgaaHlLXaLcfZ5SKmSyw1d4IN4ZfLY+3FcM9UPTlCpF0+cQn8jFRbc
Z8C9rqqfC3Vn7xMDalspbD0zvYRuLBWpe9ssplBwswUDI0yk+ThrNiJcW0CQ0xti
XVUoq01HlYrCLDMVhelig39dvfiLRti9wYqdTe0U/6vJvaPdaqK3audcArfg789Z
UHWJsEdv/ojVei82BK6NhCsMdgIylGURpgy2f0nM7SNFBJ95IIvvVOexdv2WmQdi
X73mBPV8JXfZETfX9rBrR6a65IAGA/L5tjT45lHX6p+tS1FQaveb0XqJbyCIMTcg
xgYF3vZ9O6FG5fZEZvtrkA6ky1znbHKqthttaU/hpRyFsx2wNlRVbuBftlt+8h3n
SD2ZmOIiadVRr2u3i2LTO37pvj3QzX57G/VFRfDxHKoaDTbpAlVttD5GOgYDGg/q
0T5DufoWEiPSsP/kqbtssd1zoWiucCL50ZRaGEFL5ptzXLuVPVI6XQdsCPDEeKsi
dv7l+emMHg+KFM+tuqxz+cCXJRM10uXRqE60ObrVu+cd8ptcH4kX0g+22eDvPDD5
1qULrOdUqyXjoRWJeQurZziPJk7C7zVID/OYsdFMSv8wMIW2BKClCsAVwV2fI4rR
mF6HqKXeZtRhX4Xr7vYaUakqnY/nELk5JVlEmmA7qVdVaZIN8x7hlddQUGK03Glz
I+RLR8cIwsTnu6h9X0zKweTnIEfLXUpxCkuA+SZp9T+vV1FKnjTGz7kCP+Ni4OOl
lX0HGY6+oT+gQRPkdCtaiYS0EnomutD7Bgi83oR0kbNABIeXqsky/RZqUAcnoFdu
SgXStMMjsAnvNgpmj4PUlVPw64x+z8BmgOtAFH4TzdtDs7biRxl4T6YCKucYvHcE
Fn3G0RGDy+dN86uek1v1cp/D3OgPhnzXY5UL2kvzeqOnADvuPA+nmB6wdFcn4JB4
Ecj/kUudfaY7ALVqd0R0TQNLrsL20rg2qe6WacPxYVbjsLxm18tlaNLZqyhreaHX
rT4Em3ZS3TAObeWHrEwg5sMGvjdGwjKTjGN3DEWNBR6TgwX5pW2H//maW2I2ORh/
lO++8qKHO9Vgqq5WXJWMp9HPL+dBuPmHOa6EUSAwnHeLETiafz3mbyN37zzzQF06
sW+aKVSyguP6L9rjNVhj4hx1FpUmojzPcArHBubPZTsSsvlotc1RXJSE2lhJ+pAg
+ZSDwu5HE64AFqwC0Z+xeQdJyk/t8MMbEwdhdbQKb8meTSAtfO3kSFLXlRPFJhkf
Lpl6QiZhmk+sbTNq7b5Jl6GmRlE2tbw9i1qN+lt01WThzCCG8DWw/6Y4gx5Ceoz9
o/mYnGG2CMj/Km0QdjsLLa6zRbfEFyY/X0igQbXPk4j+7lwKzLoYnjrviPjrcMAJ
d/fPx9LfPp+NtXIrqnlJheozT3RP0v88oeHupYWuS2uon+WIrccD6fH+BV4D3S8O
2FiWqzXge2/nJf7WKx8MMRuAdZj8NK5fH1/Vco96CRmoBAXsr25PaeiNMhA7LkhC
OYoaIvYGW3FSGZe85xfftRSAEXJ4iZJMiGfytt81W++LqJqcTkeizfMvpvIWer71
caeTiDtmo51t8HaGZCvi5s473a0sBu4kx/9cu14b4j6bzsCKFwTWtgtZbInSNgea
nUYzYbgymcDsDjjPAUXnGI1NlojStaw0km2qnhV+ELBzIJSOMZYQUTQvfcqNBZf6
Dq3fenokVWVSodfX7LI7sLnKahzcI51nEw5b7OiDL6PzjBpXuaiVacwQxPfFweOH
QqtJqZeU2pRO0UUlo9W/7apmnhoxNeSbOhBfG1HqF+QX4mUfEUbpq7MCrkjiH+6w
rYnrPltzBpuyRks3xxyBkmizS9gWH+lZhf5ReNTyepewS0KQKPvRfrMp3io3ReC5
n4NlvyM8QtL0rxZ/3vZtv8mTLHrPpZncoO9S+oFMqmaZbJinew9zRzChl1+MTABm
kp950Hp85MLr/sLEx5LME8/nNaocAn4f+XeHmAWDuN/3LDknPfSj8/v+CmRdDdyf
pKusPtucJbi9z5SNTyTd7Zn3Rl4MaWjOPrXwQlP6kSqIZ79Q81vm++UesxtFCMiW
q0XhLDbrShwX4kkZuUrQpeJ8tvmEuG8hkmcQPS2E/L/Te1nH5Z4rtxxrwo2S4TnH
3P3ps1fETp0DqVnLBSkq40Swu/10ryv1qCQCxQWIvSMitWXREeuIhlUTe1UznU/W
HJNI85xvsY7QlPec1p0VY4/svKg3/o1yjJGhPBzsEKQJFf6QHBxpeOD5Mt2lWhQp
zEi8FKSHXrqi1tjUtEcPZJmArxlIX6zdyQh36Y4kAJtAnW0LAApROHAjOqEM96h4
XlbfC9doCL6OEXP8lQhQK/yVnVQbtUMvu6xTTkBnB2CfI306AZv5zlCFoiv1RBmV
OHE7hHlHYQJ0sHkyMxzrKt42DfG1SXWFgOOeohWZc5Fju3rM+WJ1e0+NnbPPndOM
v/alhniAzOVrEob3E33Ga+BfHqJfFhbl8R2w4PSlDIigmqrJbbstndSTzRBbqerm
SQS9szfy1Fr+rytBdJUIqLfmsV1pNeeUTObiiOYvPHDatzuymNc7R6feLkjN2Xb3
HO2wdE9I3+X173MIg72NasvIbxmvL9dMPiOjWzFgaXKMD3TnixBv/xNGaxugMrO1
p6wdg/b2NV238nw4uZlYdWxKrfCiECCO8f+kA2Rg6u27CoHt8BhSQ35K5rIH3g1l
UKj05pzslBJYna1vzYL90dNAgrRn24RUqXDArllzmfja9PqJB0E+g7MIpjOM4ON1
XMDUYSUgi+Zsl5v+ww7DPKpMMCFojRKauDng9sSz2AKo89M/GREUx9Gi8LN6GhG9
xXHEAyppjIG9EDlvaHyUhloN9eb5nsFSbuL3tsd5mYHyEWtF9OkWZDjSAsSCN4+i
MxrFaDfJqE77UywCpdVOWCWDzMFUeB7cb2UmVQZiQVnzDGvd+F6xR8YuVrrJHZOV
BCme4GU1Fjc4/5+SY72CQf47Tuk24sCxOlh/rLRMJY7rOTuRW8RPfkbFdt59Lm5C
9S4xx/Idz34EJXWv+Dv0F/+qZ40dSxShxl4w/3HFUMXK5yMSSMWiWMWVw42Ln4HF
Fk7L8cQZtMXVxnL+UDk2xtRwdQwI6g0DQWttcOCoQ51Rw15dEQ0+GTMA8JKpay+n
i9Dt0KX+FdvZoSUeNLm49ukPNQZXoxIlk47x6XVcT8177MdGt+HbZAbBFfo1c+Ua
JjMZlcHtIUSFNYbaHLeODQQp27Uaw2G3Fs8LRPyhoYWGD9R28SfAYNq+O4zv4RDW
ywp+kM5krtHPCsxdRvrdfYX7rUrNkK8JWa0+VC/vbE1zX0KT2GVi0LSgMlr2ahGi
SBPmVh3hhu99B82yH0nxvcvSZVkA3CQEwKWHuUWZU50YyRAry6z/T0w7n/OIktXO
rtmjbKtcHqFP+z7AtpgdMp0dio3ScezOkX7D9aw2TUsWWdfV4HOvOKTWvKVeFjzM
5tt9FsdI43kQ7bWTuAyLjGlKkmpp8ywAaNdp+xeC9eFdoeZj/NLbimOBiPkr3JBw
2F1ZwT6XQKeuq4DfNG8MqXUf4YggK365mUSF1vzTmx7nwKaQn9b7AnTih4Xv38gL
cfRJauGOd1GVkR3MkYvZPa2TtWmDycgEdPQWbTBn3S4SRRvNlQutaVH0WZevyDOy
HMlGEwbJAXOTWOTBlmM5e7Kdm+Ssoa+LpYJmeOvxw35axlTcoouSjd0IJFLL49j7
6G93QSv5xfdRBOg7GQA1Ef0Ml2bT/P4zi3JS0dwXy/Tic8SWZqLjn3CdSVF6C9U7
EOFELNA4DfyDjHLD4HnuESvpfL9dpmI4L8k/ai34RZ9rzcYviX0QaYaW+KLmKZt1
Q0c7CfDUv73PcfgNo0V5WO9/qDRi9kVT9/zMMeVbwdspV+Lus4oUbZmvE4y87zkV
kkpBuRFGurr9XzmwRpk0fnojNkVVPaC02iSU/XN0U5POpCFogs4THRu0hmk4xXMo
aYBAd4loxwR0znQ7EkbseO0n1X2COHLZTnZCAjx3dnx/VMo2xuKZfxNhYm2r4GTA
BTNdi+7ibI1hUKHt7g/JpM8TJ/CoHffrN2nO0xIwPbvgSLqTyLmCjDMyKfs8YYk5
yks+FJVONajuDncGk/YOxYjMoPvPIK5mERJ+UAFDNnKnFR+A1P6jKPNuU36PqhBa
sT0jSm+5bVCxhl0BYPdpbxhTzZwgskAyB8NkJGEI+X5ReWkX0D2/CPHb2UnHSwDh
DdNOtvtZLHX5G17mt9a4hjHh9s2EzAT0Q2f24+Gt9Uf2K4a4N/5QOIvnZ/f3ls4F
lQxt8UVs2t3O5d+hjcyk5xevH1dioROjeva9/cq1b4itQrIaA9IAq4VGV5vGq59X
BFR/LKBpAh/+eHSIL//aROLuPxiDHHcjrVq5sC76UiWiO7cQ0Pa4asVQ2v9DHsqH
wyOnyRMEt9k4ZqJqUEBe1klBT+3YAmEOwOlHJm4U3bBlZZbYa26lAqaKySo31G7t
YtQ9VXFcmeDVH3PMaoZhSumJayPAdw6VCJ0Ck2pU3bkaTgJaPwnr9mTmq/nH+YU+
jFRNxteAhiEM61HxbuUbk2siwfM6RLwttcWJ30f7uZPnwofPM/9RptdI0096d6Uf
jIguIOwPOgEAv0cbMGLywdP5EtyDyNOW1BcioIxEUV6D1/EGFI2aGKE0JARyVF0K
NoWLwTeGqsXOVjTTdSRF6Y9YCn8k0O+O6JwfJokcqVIN+EZvgfnVOY9OjD5n/NDU
ZRD78fyCb5lZAv85PlkhKbEuTje6Ycs92hT6WbWbxxs5ezFBR3moRSPW/ZSfwMH2
cy8ZL/CUCl0/BvUQ8B431x85jUbuXGowyO5smh8fyuoSYkQX40CbFz6B3innSpEA
9D0u6s1uMddIealY3u0ZnhdSJKxis1kPKEVyBPvkC8W2WJXzxNQIz6enInPnzU7F
lrK5kOeM163KAlh5nOOhGmtK5bsVicThGIUAx/erhP8ecFTY/+aDGM/QnOrBOOCb
cuqQCHmBmCGrZlw66lYD3bId4C5tYh/6tqaVXA+NiOhZkqhodH5t/JdImm8VWMMH
zXSddQ2/iTBgOUTEdv+50shx/H6nzkWhHUI9R7mH7H+rIMgIZxU27KHL5/Nh55VT
FYA5N/WsoDWgJTZIS3wz8GsJj/fnUdAPxKBffkP3/7IhdSLhtE0KtxPKLn+IAC7l
++0eddAMvmeat1Tb4cKZZhPmz7MLjpFTECbzMKS3ENWbHaxrpOvvO1BCKM+sZrY9
XvLiahp5pK41gizjMnSnJ6KM+EG0NdskSl8x1RVVm+PsKpZ529/hlgdiWxLoZzGk
2xB3K2YxFnMyEdfklLtfqxnJe0svIuqkW2pLszh0P9uy6H/XZ5SQmc9dV33S5aff
0eJabMRR/Aq9siWajmQlOrwPrkiCTR4YGDvQzfdzYEJNCGC3e9s8bKqZYERZE53f
SJcudtLheIirIl13OlNbrjv4uBy+qCIgZl0/ZtYh3aUTIQQEQK+YpRnc7MNaP1LZ
Qg0Bl+Qv7K9APJbaczjwCgEbDDEY9CvhVfegYfvgjJtRg67LxuIXGmGJxBnn6PKg
sYejBfw5YkjWvfzYjFM7/oDfDSa6ir0y0x7PDhZYH3WDMo00GhtzF/ze629EynGl
G6kQZT41iBcIoect6lIWMxj5UFhyC+PNKQcyFb4q+cg7Prh0B3c9UqiR4N6QhYfU
clngmeJedyC/m6KdrqQo6uNxkSjHTpDp/jA0JjTSiBsAzIbW8B9oa5sAlfq8/KOs
C7xQ4Yzx4V6utHcUo01KJIGGI9iMxng9rqvLMwIZG+CIj7UI1uf4Gnf7+Ac+Ijma
8X0HFj85LQx1uB/wF0lVSMpMfNGYfvxqR/qbar8hqgX495qc0KzYjDTKCCGR4eZk
DIDV1W0ur7ivePwWhA/UDO4Ar+xKpLhDS5CMNfney/LeUtXESsAhqXpbRkRmaKtk
9oWawPeCn8EAmrGO8wYonq9chX7qN/exwW9y/zmX8ZLHqDpgnolBLLPKnOhrZLOr
iHTX4kLgAULCVTBT6j0y7Bl2JRThg/OzKmO72mr1wh+gSDckSYj0+7Mdocs4filg
H/L2MVkoL5ZUr7MxoXGezZQ+nMxnRm7N1EDBeIpS9caV2fPKrcGPS1/15S2mmZxm
TtZmM9U5AhmZrmN1+v2RIQ2yh7mBJ1eVAmL3mmy269sFE3qgjHdS6GbZowNwb5ew
Dm5Jqjj1BY+5nOcfyD12xvkUNLglp0frZWQRIr7aQhLT/5KQdvPar7teuQ94xvmq
XEOc7PvEb2duDGVSc38/TEgy/+QTh3VsiP28hz+hweP/PBgfatl+Es5mSLxlGs5A
2Df1F5oK9G7FtwLitVuVupYhm+vkd+7eXAdgGYiFUrmzy7iVySeCmV/SuFaCxVHn
gCIZ1gwQvyspa7rxaGIv5GCXm8zy3AXdaPz0qBrWB/MQTLMUiCGOmkYwDmArdli4
qDmbHJS4/Yy1sd2uUlVogIdluwY7Dahf+AILkHW+dKkS0F0slgMw3OJqgp8WIbb5
rJSeN6yEbKaCfPFPb26fq/8G6ZABV6iX6YhukNx7rqyPaMb9/XpKriaMCplevBsv
fqm69dm5q7W3MZvolh9cF3F4CpCd9C5J+5EKSeLbdvn72/gTfRhytTB1COa1u3Ge
1B+jc/fbl1HO7L2SsCxrC+Qje9/h71PpwsruB9D5zH3an4+aPcDP0Ou8136Qccnq
FCk7VrdR9RSgtJc+eDmyD2o45hbQs6uzxIog7GBTKJP71DCJvGdbb4urLnLa+KnK
LhBvGq/VCd/nLpeXC0My1DksLiuX/rZCAEsfjBg/Knu6euY1pqVPIn8PEzg9Axhd
DPAIZf89sDxrsh1puqnEyivHqZccyXVbLJ1FzCnRHcmRDjf+D1pShojOr8OMLRgh
FbY265sC3kWIX/vIPIcpCXNCburnKHxcX2L5/v5zpi4jBmP4TOdrNhyY1INawXjD
cNlsP4MBhUz9qhyzw7/XakZQ2cnm5CLU3P1oMg6cuQu/f/h4jU/NXhiezIIBuejV
YQJ4i6ilK15kaCpqe7+XUll2CYLmKCoKWgXlV1u/F1EFlkiaK5q/mL0GR+v4xfgA
QCRTMv9FiVTcg+gWXqI5A+1ToXyYnnZ/a5clfuPPmubWhe1/AZhBwDEtVtvvoUTj
X+DJdWnnMyeksHlW2JxS16jTsD6TjcYbS2DnWHIvUxVk7o7Z8ntINWWIgP9WbfEL
5UFGoo40efpZNbLTfWiCk1iqp/SxEr9KHkQTGAyT4qySheDL8gp15TMkiZn7pkmw
cs+iHHthe36YB6iNIabS6OtbWvmzdba/rBYrFBdDsXiHAvDn94lFNMDLWCUoCQ9t
aRrgNxAqVaQ1o/pRJG3q5LKNfN8zHpwi9jnZrchWxbGaHh7IyAkc9u3M9oFwwglE
+n1SvMpZJK5XjQ+27YWjDswgAz2Szlr+UeYwpJB1WEdG6943rJrhjQFfQJaXnwan
rkuCKUVBUxSlJ6JyNJkrq3X49jFSOcf9eUm66lricO3SiBshrfFzuhTopwjDN7pG
0uwJ7GmzwZRmR/JjalX/9yZ8iBTwE0V6UNJYQVYMc1+HqrkD0yz1YEHW13fdEdvs
TAgown4hP5RKDSw5EUexEE5IDQ9HnzkIIH9BjFqZMTaD9gIabXMj/+/5E6w8Aflq
K8CsgH1iROF7rDuTSp5xekQkySBzDyxkMgCz8RZnKwOkaQf4vUEpN+So47h5OCvm
AqJiPCKPp0XdJDqvrR7fs7cz+N8PEjj/jE6jxGgyCtGP+/zEinDwrLiDQTvwMEE7
PJ5kzLqWI4+D9vUcaMBjyWF6OOGonxn8r+rog0jcKfDY2vhIzg7X0+/2hqVrY8W+
Iv8wdgzDlFRTyKFF0sPWba4R57RFFTtyC1ZanTZstZ4vRp9a4u8EcSFY3tLxjBAZ
Ewd+5YvHm9mCLN3u/adIl1nMsgy4Vbo8XGK8kKy17oJhORW7qOK6QbEEJdAArwjh
tM/O2cDRP/v2ptxHfqisxRtWSZM7y8tmZxRvM1BEbPr7QyTC75G/pCAQsJtvpTh3
SIkhTtQOxOUGxiud4xfICcvI6OxdpVTolJHXVJTU5gNf+4nHi+E0PAB/v92JCcbk
RNO80dAg3Rhj0UAIvwK4Uy8PbK9z8WhC54G8DP9e6ifsfwACrsnNsJnkizA09FeW
Fk5Ed3ayo8LYjFy68NFi5PEVx9TCYGbsyc24du7d7RwRMNi3z5XjfsHXEWf0AFkI
4TSlO7e1TxRf8Gjbd0W4ql+ctAPt671HGzph8pmAMpiMLH/tDHvwWBqJ1A7LM/+i
GHb0kPv83WA6Przr8QTIVRu1Q60gZAE7WUOWpB5Q9a5eEZ03AOvh5vM6A063ZQIg
+JXTJ0aiVIDNioNYD0yOXWFM7hYf6ySZYNv4q3tPNXU2JpbuO5/B8fgssgq3o6Fi
yG1IIVgjFYL7fo4WN31JdaeDcpiehNy0VS3mxNDT8WMg5O26rDCS4VcbJfMs+EKB
QM4RD+vQC2ivgPx+Ch5hNgsTRIMFRdX3hYhML3PZVZqLmsFqJYAQy1/8k336GUQ6
PDVtly4xNZ5bqAQj0OwrTAZKqjDXuKlN0gNeaSCkAAC7wHYguXEhuQ5c+Bl2fNGf
nbGi1U6eZnmpF1PsZX6Er4d+ZpLV6cujIzcjWA2FV0BTVPG60g77kxcsQPkGcba0
dC/PYYKVgDddnfJM89Zy8CWnJj5W5v1TQqg+7QsWLFTIYEEzqlva6QRjpMhMMPoc
9+LTuFAd1Hk9F/RvnhFgSAJqX/TOeC4zS4m6iR1VN46kX4nB2eI0yp7iReaOo9qk
tUCDh6IX6ZN7fewjcZE92Zvy8GWNtcUb9RdwDKDzBzlABimt3KCqsyeonqkSEeKE
yKK6bE7unlqjR5Fw8MgJf8MgSLHiNt5u9rsAuFUTLBBFC8m0AP3wpQ4vuKZ3eAml
0TDUIhW5MpOz5M5v1jTv12PJhJvpCzcdVvbpML4wfm9L4K4/BeLyZA6pSdfS7rcI
iPb6RMzVuJ7+DhvKbWgD0xBLBy0ddieqAixjBlu7SJxuTNmCIphVYcA2BiYZeFh5
5nld7WONpRxOfUKcgSoo8JO9FmRWkkfQqLn4UyhFu0+fK8zB4xIa+4nsttjT7qlt
hN6g9I7ypoOEbxSb4IwofmcAlQ/T89iy9WUL6TRPibNHbgmVfULPm8ulpU0j9LHl
QKbPvyWi/0hFq8fnlTBM9emp2UTnWnW9qyoNyMJb9NESumdPKWnYOjvaiv/MJUoE
MVvVs+zoIQHfgyoU3Fbad+TcDbBbUT3TlM+mqgLSOIQxVK0nKOolu22bEz/o36yq
LAQfcRGY1hR/RXCEempFWuRSiKW6lrJ/nd2OZGdU++0URqWAqxa8GYo8OFCdlR0J
SAWbU0umhA47ArzjPWHi/HEr9zajKCAOFEP4NEfDlksIZ7kR8fskImcAUc0IqAMk
hxH66dLt+IDWAnf3mr2f0giZ+5fhmENRuy/maEM/uFL30MLFyrjY/h530VbONssw
K5dZm9T9Al2jsrXW+VuC9/fsc/oHh6iwgiBCoY29ab/A1YOtmP6/1GCOXjtS+a94
uc5oKS2oxMRMJZH8tu4k163BszYqv2XzSkLruHzixxkcYgmIS84PUMijEDB7dywq
Qza9iUb/Uf3AjgE8oV2oTQA1QDuuyISj9gGk5G/w35zPsqvfSFTXJVSiM9l7DjeC
gbVodFO+bD3sqlNggnpWAArQWUwa4UabWDf2oqa0AXHFxLWrE6M+st/laxEKYXIV
VOrdCUMP9gqlHIJ9A5pIDqZwfHmcspfYRcPB4zgYcvL6Q7lYeugSBsqMw3eckMh3
f2QkZc2S5HE+BZiQm/dFQ1pYVNayJaJc4nAoVmg9Hqf1Q6h/zfpmAGrd1UeQrwv0
TEs8FkNB2zPs4cTkjFUg2iwey+Y/jrU/Lp7TTu9yFHVBNvO2ryv2AfravR8QSFpg
9pGGrGzpqN55efkRZKmfPrVC5Dj2h0mU2kSaOF9YAZSNLLAtdgqRVsatbU0yN1Zi
DMWHyImrUZGZNJ188zRfbGQl7P7SJoqtzmG8XkVZFq8W/2fsNLEgyd8tdnXMos6K
9oOxou2/YnShnSgLKxE+WYAECf82AXnC7cU2Pw5VCf2PKSUr5rPPAt4yLPKlxPxC
1lTNngOlR3M0N/Laa080cjcbu+lSAphELnlIVbIgDkQh52HGscgE+QmFKpjaSyV4
1B3wIYLNyu5YEwJmZGKAr3RwsjCRi5+/ZRO3zUimHQZ7AlSRCMjfO+DK/9Mf3g0c
A9rZWruZZe6J0BZaMoZehzKEAl8TCDW5xc4HcEpGZLPrrXCDtQQR4CWQ8x19kGSM
GwUIw+WeEcsERFzuB81CVgOgbzDSE3pave2HC6lyfiGMuLKduIya8P3uOG2mN/t/
nY6XhIn8t6b3HiA0GxYKH3bunQZj5SbcL+eqXP3s9P1Gx/YoNzneF/m6LfajG6Mt
gkOCFMwp9+ChpwHlVsnCDAdefqCXo+HDvuqfm9gLuvHEERj4Pl8Qy4xXbT7zgtWi
mHwjzP3f/L1NCMHma12BC5uTBokhgjWyJSAOojPiwKn5wiHVZQMZoe3ftPJHCf6a
`protect end_protected
