-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Ndp+A7DXevohMLk6sH2VspWNLCggoiAzQy65S6sBJY2NCZWQhF7xylm4zXEhnw8s
yWCxD51EsrEd1ijv2D3vTz5nH9/ssXWvmnb9NsNZQynH1hYVCox0WM0OadFLy6Mq
Tgmn/ISqg+LyzFwULKrXtig4UbNbmk+ZEEI+xL9RMsk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 14311)

`protect DATA_BLOCK
1xsvvWp9y7V6cVX2rWLx7vgsByUD+6+5EWwt5e3EuttrPWkdbOU5edFnWkE9286j
GCs0LoTvcURvqStCyFpgClWAZtqyDA/nY909cl2qmeMFDpDxwlkvxwXgDQcBZwzo
PtmODakG4sMXMew4GiMaOHIbmtass6vKWXLHA/a9T6qV/JO65vrMdcWlJjYaW8Qp
ITQnTyQ3jxdkfknezrB0xnH0OUicUS3/41R5bZRsEVv8mCSxLBN1UJaI4uPbOaf0
D/vkbtjMoZKLQ2eTwIOoYGoWcDlVMnPytnXZFDftvOSuD9eWlFXCYz18XcnAXZch
XIcSeZ0uYg4rGP2QACZiz99d3Y+YO6W6tNWYfMi21b4YDyPz1QNaObBi9J1U8nce
G6njW2pYCOey2KJnIPGbNQDkCGfTbPPRHrsa6Sz3iFivziK3HBHfuXmwrOVbbWXe
eBQsczPAr53cTQW1jpMN7E0EHJS4u0RbG1uPYN/Xy3vt3aGdNdIcw4wLO8ReO4x6
BMxWUvrJs6wl44g6XpA2Cqg2ef1ALzMKdjNgilCUy+wUBVWT9tXVKNTSy+AXp3Hn
oSClMchDevmFLwD01NsxmCSsTuA0+mcdrwkfIo1b3lEG+wSEdsk1gGT/Cfbx6+PN
uZDL6lLtSAslDZ8Ad+VXbm7gGLDTK0lp+3EcW6CUYEGEJ3xODdTp3qRlBADWFq+j
B2IW2vugec/S8It0jnyrL1XT7LUVYsNPYIbs3bsVRkaxrZ9CHwFkcKgxaukgHCzy
3sJoqxJfdMc0tuBYRpeaC7fjwcubmbu4XZjag9JYQFcF0YIq9cbXRonZD4lUtjE7
f5bx8WhlMdksxfuWayhpr8oVAAzoFN2rDRc+Xr6zOPrH/3pgC9sJ/SaQq0UyUYhG
u9L4nUHCrw9UPEBieR7qhKMBE+b5F1G9lCvGj4KG91VHgjtY9CsVPgrJYh+ESJk5
YLbPZA3Vf+sVIXc5TO7c5KlRJ6vXenEBDb/OuUqb4jgfiZATSNp2sWxh8aUSVCcl
uV5tLXJd4WroiAhCyz+6pLbZdvthcj91zjUnJjkt8kGjnlJTfkRdB4eJlzBIOARL
KOIQOBTVaDVy3PBH8+COItecNQJgIrwWWkyPSSCVEkRKKCsHvFncliT7palRBwDS
ClbM9jQBCussZGyGaL6eSBCedsm4l7L77IalsDbvdWg/ijobU8SS5GEIgIRgQbvl
pBVXxEtwCRfZk4T3IMx8/6qRm7aoPXpNyckobubf9khbOQiTW3C4m5+ryLwOXuSY
SQhEl6iTtlkLuR5tXr/is2yOmqT0Lb5GH9ej3kfNclk9tJq8nT/uRSeE63/dAfvo
z/F8cbIb9LvWGYZ2idCZwDtZQdb9WHMLXBLqShuNd8tqShnRgrAaldnoIzSH5tX0
MxsP1WB9TlIBU70yAhmL9tSeG5GOFm4OdMKxRbdgabnHwWpDdERJRYw+mNZzKis7
n5L8rNboyDhMUZsExO/wQXfB8u1vCx9ohsJgl6szY2qR9e67s5Ml4FcWtgAGC/k3
vPW3iCYAmjxcJrFvORlRbo55R+L+1RyWhCoZY28BFOmeyBm5/SrfnMiVFsmO04Vv
O9qXIJgjphE3GCH72S+rYMo2zOBq0+flXhVW65YXYLf+7zY/GOYf4dZBkxCEfa8Z
NkxjFCrEDzr4g7XniDhse1xHSeSXHu1ukwoj+Snuo9IZ6vAruFcWmpdaoDN5sU2I
6r1fAndOgxtRHZk+ltVs5kArYisDuuXQiCToY7Pl6UnVf57TbPNUlG8YQjUahSTS
y9bCn3eGtnP+aMCIFa7eKloySKja6XFtmmgrgLRDpdSev3h2J8CtOcDo/zLYIgr9
Q2RW/vT0COIo79oHsqHN74Yc6zdDFcsf6FUVoNNwHeExBgf+AfxwISnGjJljZDXQ
Oj4OjSwXU76e48b49diKXA2h7BJ7Nl0tDudRsXu4H3eBppUAIwv9jFo//8wzcRAs
+oTvrQiSh1nlgTyhuGHxyXkGi+Ycbe+Og59lro3JF0AnorbpzpaSLuvIoE48XG6K
RkIY1dXPM7g2gzx1BQb5IXIvXSlz3cMoFq71K5pqzrE81oaYCzz+GGAUqlJID1N+
MamrPSyBj7pydkj2vOzMYV5uqiFjKsevnXATGuFWl494hbkjRLBfIFfEEaDisbZ/
5GfgbNzGw7ZzPiqugZDLanuPZCZL8NU3kPp9l/FQfsYal/E5N7dxV3RgCFfPP6Ca
zXfR/Aa2RYvjb5L3xKlrOaq71K4YDa/6KBHasNywmHEBdlwOmq7Q4OqZCzPCWiu/
DFKfstWbIHE4/N5G91PSJOiepwaI6WFuRUOyvD5B2Rp8oDJk3W0GH5xflMWxP3Yi
jeiNpZEuiaAWK/DQjvxTVWWKKbszN0OkafYTc58MC8uQ1zYUGi4JTE1XTb4pUHCI
w3modWnVu8RKVM5/ISPwGkYtlXZKlPpcU5CILDrcnDGsmsNEEDduw4LUm8cXRzYd
Xyitbsd2hxCvNEwf6nANvsj/7O0F9ecBQ67fmHlBnFSKfbJqPZn7Da1+vZht5RJD
/2P/ScgCcnOiVhFukJQmR6VOZxMt+gbvhaVZghZ4msdXEw4CWGvnZ58hQA2745k1
j0jkx5yvfN8PBY4djkcfgtfgdZxnklKFgQN82jWkNemzDPZTs8Dge30cL7gOAhcR
+A5sJtTY+psw1enzY4VqGQObP4UNUMrm5xczCD+ICVpcy/dcUinSymS1FPBLFXOk
mGcKuV/o80C4lLuNjjRtEiq8KVMba75g6lZQmR9pFMS1i6Go1krDh4WbZ0/boLlw
gv6cKJqdUM6K8bRXeR+lsZopArhl7UAz6j2uGHivjJiKtyaCqG3+SZtFlZsdNsWc
2zPT1Anl7uTsKD+CUkik2CkP0Le5Mq1oygO0dpBDhXPlWXm5pSC6cWwEgcOlhLHV
3QFB2LSzQ6Ffo9Aj5nS29Y4woU9wDSnljgqZJMo7LYZJ03bakwR8tC4fKRfq5vCL
9djokOuyPiQDTU6nty8eewoLLVdwqUBA6AF4xNJtW0f46EX9/7ff2TQfGuP6KAzN
SspeRtwBwlFAiCb+lMY6WxVKMDLf18leMB6JKSxan30cSH1F2F1gndiSJQprraYr
+tizSFk71Cu0LUZKwtvQEeUhCyVzyqkZOkKTIcbbagP6k1TLbrHbDCeV/rBI3yjg
jObDHoP+yg0CqOFt1pQw9iaMoM3xIvHj8+hhooyKoOBLiAJ3o/ls4O1TwQvGqR4v
nM1FmWkkB/R0xf9l8bQos8md6iAR0GJIDwrkOstHhPiCWvZ2yriAsWPWVjWJs+Fx
8EWzC5OmNDzoXZy1KGyWRHSQREYHoIwku+0zoqVeRWmfUHMeXyXCsYAW6WQKTtdc
WH4shWLzG3evXP7cfGntmKnCwvWVsMB9R1G7wqWcaj9ET2Y/YsrbSRDVk6q+ZKCx
eG47thMq0h5WBDVVHs+CYg7UF6dQAHnm72wCIwTy75/u1IDctMGHmb7j0+mNbZaH
vZFF+0bknoobjvmb7l5JaOsaUGltxgO/2eOm5Hz1102xSEUvFm/7ngTy/FdaF5Iy
XNBhbwVFXa0KA4rCuvr7MzWcfeqzbbjlxlrzNJPZd7+T5mgyq0uvFQxOY0wWaw07
CVPQsRxJMI6Rf/7tMr0BJkChbTtrMpftmNOJM88gTIf0I7a5wea4yfLMvHGdCZs0
NfXI7HsUoffbSHcuzSJ4fl4gpNbTBJqocuXg/pp4+fUPVpT8o7Ueqc+RDGb62PSs
M7hgLPw8plwpnif3rJ8HXH/F0uRRksRCKlJiSqCWJjJR605ynbU6Y4PH6lC5i2S9
ivAufrfnT0mE+Mfg0Z/dxj9gG1mqnDcsdn03av1+kdps0sdWzbK+GqR6t5gSSKpL
BrPHpM8U3iRngp/vMIQnwwQxRx0V4E/C8SW/mlUhVeRsS8ss8vS5SF57CUcISXMJ
DFe7aU/1VHBgn1JbsNQDutrUCFlhi3ZEqSzoLwToSbAJdlwXfSeBszL9/R5PQnoc
J7189oCDzAwPPBX34udcRAY6PMAP+Kz9wZgCvNXdxoh9bxVvkYUMfTzT9D+inEaj
XHcnDXo7NxSUJH2NdW+2ZgRpaRujDi6qsucqNkTuD/NN0w0bbVMg5Nyj0Fq+lD82
nyybBuae1DHmNcmgQZq8isHhRFrnEd+HKTFCYLuAjK7D23hG09+o/9Xz91W3gLZc
FXkqYKgGJmlc5Q0KOIHLfsbhg6BI36KOsK5038ZEy64oE060oWzHavhn9quc6OtZ
+ecFRI7z7l6mks9byBn7rXqo7gq6IBuH+LgJOhVQctLOTQ5CtWjQMw22Qq0YIvTK
DjLqsFfo3K1XNySvEa93HrTlAZ68b3dSKDpz5+X/wUQ+XrDSPxdUS/KVeZCRI0Lr
GxR5UyTO8rZtm+Nri/DVyyWCJl/PrKJpT8xQViPbhfu7xGIVy2gP0iM1nYeJ2OYQ
nyL5yXdsJkDkkfXAuxYdzKj0gru/p+lAsCekMDktJO558o2h2u83/q8NT2wm9iVN
Wwjdx7gBELqxmmoQcL8GhA/CBe5LhNthQXgwOE6iesGmjKaO8iWr21+wMvSW3/ob
dWA56Mq1E0d/cJhAD88L8kSX8/pF0q01zbhX4i5syzCQ9ebcHSLo6sReeNI9WDwL
Kd4vlCpiA+p+oE5DQ7fKqFf/EF0485nn5nN3e6pXIEg2pt7BUfbQzEFCnWHmlNAR
OpVL2UZ4ByzFuFIW+Gzs68Tpt0x27N/UWsLYc4jLPEhlEMpo9ixwGvLidHBZu9jt
EnRqVoINmtbO8IMQyqwo5/942LJ6oeM9gH60/d+ri/eg4bF/x5qfEdJ3mAJ0Hbqr
VvWbZKQH0to1206L8bAMHnzJh1I3sNiuFkr6D6BiEC+u1limZ6DCRSaO7GsFeh8I
jmi76aGIc+s/ZjF/PNDBV5RVy8cjnUqv1aw9712CH1tSVDMM3BrFrvc6uOXicX8x
6brkLib7vsmU8ofjb5iq2sM+133Q7laFwrVwX1KqwAUoJosteaDIMYRkSjJc/iHP
aN+Hg7HvACkwaUDoYqfhdYfKk0H2nEPGGhsIXKwGvuY5t2T30qKV3kBrw1EEhI0X
JhXSkDMtZyNB2wleN4L7yISUdhwULuEsWn6vwxTTWzrrdlTiOb1pMGIAK3dpwhqi
Lh+0/gw0q2BlX2R2dIIMzHuRGdZF2/iRfcWsEb6AG144KOC+8cXInaVEtC/zkMyt
qHllNEFyUtRhVGCVuOu8EQbE6qrU8f0XSWowquK/8hS40rwJkhQoq+8EqZUXfG3n
hTb57rqDuNULTg2EhwjeW4Rih/aqN6kW2OFH1dFx4AjpAk4Da7BWF7aovDKtOY9J
RhFk3NenkNVZNmXtkmV/pklGQM3QrhioWrnKeulvoDRaBXvvFXBlG5lj7fIpzos5
7D74ubRHRyqH2VkLeV9imd4sD3xfWHCS3OYi86SxT5bKtHOAxknFC2pCwmYephkx
pmfPC7nvBSn7mKS7bxl2n1Xy0mxodVESxp5CBu2/msmlWjsWzyg/aBv3AVaiTjBM
XJdXhOhuz1v+vx3aLYPI/gm2h5RsHdb/WgFon+Cj24fLxBCfNANTzD3a3lvL0C7W
wvTNpqtVRncHv4hyrJ0YzbHrQkywGhYdc4iDgwoAw/IJVsIlaVVO2fhCbnASTqsS
uA6DLMjySpQxWnv5AMgTSoUINbDVyEKA2hKdY5j2iHqvvEy24OSgwN8PCZfJTCp4
W2SDandYdUn9pL+qH7WjiDukgO0T3vCH4g1WIYLAYoIUEP4B8XaAr6s/03s+1cM5
3+OOw7fLBxgpLOt4xO8/bOMX4MwiyiM8LtZrVbOECYpVD6fABxNCbUK0ZoMp4V+X
F1lcdA7Q2OtiveOCc5RbvdZ5lzkcHxyKa3FxobyToZ7qf+HjMEIAH7K03r83EvPY
+gYXQkz3La/gzyK5LYN/o1lCOZtzjUaYkhX9KddEh7hlWyn3OFILZC7UTmz2oTgw
1YUO/f2U88wc77/NtRcEbn6eABW72gLhQoDlXvYQTrPoxCGxpdF/7SxI/ycK4Nv0
05UZjU0INSB5cAm8yEoDgRIV5sA86VGpvfop8G3LkROHjr205TCpaN5hKJyO99kV
jARBWW+PBzCzG07a0S8Akeh2M4NZEQfmuNysM9P4koZf+yUkptQOUXzNAFZddfa8
fVocxcoUlt93rHVQwlCmY55qmv5yFm9DAzbr3FwzvW1afx3mdwINpGjvNMSiHdYD
j6XtQjcqrCpsiP1aq9ABzJOD1Bn4lLQ3fCx59CD2b4kToZiQOJwdQQ/XKtrfZ+j2
qWcLJC4d4RocXaxB6Ph3D8z4Hhl5doRCKa3fltejvbBUpAf3sKtYVRuuDLGTMSEw
sDPS6fGzfX+/kcYBzbECrN21MrE1Awz9krx+qctDWMchYoXnBEmLYbUO9Oxg/N4t
tk1BQAur530mV1Pxp+DyZqhjtvveyfEzqq3shhm8Fxla+B3paRwxbmVv4lzEzfR6
ulpUwp0wVtB2+czUjEbZf1LMQqxwgT7QYPDyW/6k4CmbeYlLruKJxE9ep9vR76zj
ExRZXfyOQgeR8xp93DUj4Q49wZ3rd/usJrzCUvq/dXU6MQmFeXNoKp4iC4Y9DgR2
DkPUyUd1hHaniRhliqvflSrVtqo4S38aafgFV4IR+wFjAo91mgTP7xvzffafrHNm
0MIegIWvzuUhWXtsfJKo1RIS1Q4d0Hiass0ox32ukUQf+WfG12Td+q1dAB5sFNHI
+vs4PXfAu26gEgJb7bDNfRanlNFeDKfbSZ2TnCSJF332GdXjt1kQaRPwYTgoZcIE
n7kRWo0UaKjt+VLYZ0cb7KVJWacsh3C8fDrQZDH543OR1UEcazSqP+baMEMYiZP1
Be7rDX7XMCuUZFUp+DuyUqBQqwl2RzxYqY0+DJI/WJV9QSNJoMgQuPPCOYiZNSRo
BFb6hXo+7Ip0Ngqwxb4EwBo9ws/HLXgs6b+PNFF/jSYETM5WsK59t8MbV8KeG72s
VGkWUoR0EOBu4wJSG1pSo+M02Ytyohjc7/Jt1heziTSshzoZHyq/d+5YcfF7cttc
s6hnN5M+Qr25TmXd7+5In2lNicRGwdjJruVJCyZrXDI9q6TPijFC5ciUh8Pdc7oG
r55qxUywe5rucLMgCrXYdVDLWlCifA0Lx9tMESJDMriVEwWKC4DLv4Fmk/H1/nfv
YZhsAxvXYHoe64A/802azPMcx/j7aT2BXFqGjwb7sCj8oLMMDc/Id5VsVxPJcezi
+yArAYzkTZhOeqj2KARjow5UcPtARpYZZ2F4aJi71Fx7k7qIfvCbm5iwypdrLlK6
PXeHe9pIzKopgGCsYNiY4KmTviB3+OeOZLnqbMePF8LADjpfh7xifmCrl0tG82KU
rri9yXIuyxsXeXMb+R3Q9Si4XEoZ9QwWfZWcpafiBVWObizXqaebR+K3XTnI9gEH
Xcgwl6YsUM0ME28MUZAc9NiJlkaCLXQmhE5tMAxM1FJHscH2hYMsq9Ry6m+uVz6s
DBwWZeT21KysfE9YlBewDV2vfNJh17HXHFR9VvhhqN1F6LX5HyxXk4PWFmRaOWV9
6En1Qe7LYDZy1e6g+antGf4/iMdjQaSQ4+kpyAez9Lc6cdpMx9rzFMEcW/hLcWYI
Y1Ww/dJqpc01eKZiDmOnJw0BhvJX0s/jVM9lOD8cKb+fpUhc3Jbh56RdeEgqJs+b
WJEj1Nqyfu3QQ2PNKq5HWCgncmBxHzScZY4ezGjCh9UnYJMDRShJrET1jSjFJJbQ
umkJtU8yuNBGG6j82pVzxoCXUBLEhulWaaHUzWZhQ97F6TCw8q4pbJsgGvSIU5IE
ajDFUNo1oMpZrGENEUK5lLviFunF3oYe7RlsnKuZJ+brQ2UcfvKFRGIWKUWBvnGj
jnudVzxcjveSRZrrXfEnYvcHxsMShnn9l1DBFxkDHYo/HXXACY/+pHe8+7jsWAAj
BVaEKEPSiUad7GpdZT0xIjLBoyL5LrY/apSFek99esOuhccnu7klrXAafH8w/MAI
G/YSjbaLOUf8/THck3WVhbAsvCCJ/ZPuM2Ub8fZ8QP6o+N2OJY3QFOG7EFEPVquJ
eMuhqLX+NrXehatXreJUjzFrytyz08zUB0O1UojydU2raQRMaIGyyCog2K4dN0aU
7QOxabML0J6sNV9zNThmn3q7mKYVNVhriZU9ADBO7WSsuP87V7DFft3sBaX0DE6r
JT5A1mrOyc2xJ2hlUw3iosBy0SD5W4dgkNUc3PfW0HVPEwXU2d0xLIAbca7zjbQb
t9Ux/V44bCYerx2CDQwudqJakqETfOiL0TJUPanvbLOl1i0R0Xbt1TzU/NgXnk9j
7ZMzw3zzvx12tEnEHwXU19KLA6zcmErRyaPBAfD/rPlCEVQV3glT/+TFjobEmgl6
QezxPtcteHsNsnRyZJPf2lJ4qWUuJOtfeR5bhY46p04D7faNqMVFmQEfNVTqQj7r
vlGUNc7H9Dm2nSPBblh4Srfy1C/Xsv08lhgv3lAjVt9qmv8SzCqOBI00Y5EiTICB
CgCAD4agAg4T4M+4M2nA9Ie5XcehgDu/DBMQhJ6V6RLx+QDfBnRw9/F27FSx19/U
nRA73l19R+J7xykBuQod2sg0+8YO/+eldsbXv+7PXFsdpoXZ5fvhqlUJOJWo4/KY
mwtyp1ggQJXQcv1BoIb8cRk7gLVFKEk+QnalawiyKsxOLCoBqygpMhgs6az7R7Gm
vmqw3fDpjTuo7e3Oj0eT9bcjXN9eZqCmyeKVnvai42zXtkZOfSwrS0lGqQhXvzts
fpsAlhvKL0YSXzjiapOFCrD8FcZqnPUqIDCenOFZ4iIM91TjoVyX0JQE+gHxGPwk
L83VgRtHFklJwhOQTsC2YfeAeINWMLyvGOWW4gkaQNtGMAzUzGy8UoJyTlTy+NLV
BITNkhoZNW5v5JQU0Hxwp1xgCFEftW7AMKPe5Uj1haffP0KbI69i5SMS6rEphqEz
/0sKsbstSBmk/QrwTXr4Oej6qhXmOSGBkwzGcEg5btm8iQsfS78Z4KopTxHJCcET
XqGawFoFs3SCbhy+yztkDVahpkKzSNPidu3y+xjqBhERSmF6eMNDtA1bJjY4R/Vt
8KtngWOJYZnvxrpK0JWZKBjkDvLU1R4IW+fYLN+SxsoIiYwn9DERRhuqGSE8D5ak
f4ELDm/zPP/8iXrAccBjagZeIM/XhFMcMzlFavjIVSOyIpoh8zDUQ5qHs1/tt8Uo
IdnsDH6jn5QEEXsQ1nAcMrlclrDljV1ticF0OuXNMtvxXflZVwW3EBiNWA9cY+aA
ZVKOwCvartXxUPgm+SogYCQdtu6H3dzhuB4A8yxQ3/QviSGrMjpM/sAM+xJx0ocA
gTS/tD79C48wCXFXRPwkZTKhVviKJczeiirl1yOXM3npuv+DxGuvwwwW/aKtAJ91
oB9pOFkJ/B8JOP3Lnki+bFZ74Lm0t7uODbLsAXbYqizl+zQKqq13Ft2ROp1NZwBs
YrLFBPBQAzCEN2mRYcSc7+Mdddi3LFh7aMK09RLabRnvZve5rI2hWfAsUefbsEQJ
1+M/+B4/DBKte7alJZuR/Jbwix8VkKPHRW0ZnBoxzDC9gte/acu5NL4BZOZNvliC
hxMg/X9JhWy4ZmX4ymX9ZfPmAH8MsnIdrtm7SBms4OhVKtIX6peMaCv9SzXny0+o
fdVS089XRL4hLuYPOB0soqt0zgHUzgK9RdIettOyWW6ajInB1/gdhCsw+eWo1vKV
Yky37zHOTvo7MMTIuJnSOFsG/8Pca6onkoqUHyQsajjzt++iCf5pWRJYVXQ256Li
dbKDDX2KEnja2JH5Juc7I/00pwXfw0TZ9flPPgLbj1xoUaCwEkaX/VH39HfvcB5c
WZl0RXJET2vODd0lCEUZJr07xMbD8FOKdphL5pMrrIG/44VX+ssi98Is5YxxoeOV
/kgiDZD+J2OV7hcF42V8osSBqSv5iejorCJFjOFoUO3lPHDRo/jsPPyxGsTQmCQ7
bw3IUBavoneDktk24KTNJDsCwtZ3AUkMLg3cCXWwAcDm1Xt37GJhmDU9XyOV10nd
HzBzORfq8EN2KY+TTd8bk6jUvmVyerLgq4uU+t+xSoGh+Yi/ggMIO2QbnGbnOMOu
vYUgkzLkCzLstiuDa7P/FRl5L8kbiG2RKmBmNwVY3YbfPSwyaJ2a4wvnWClZKGbf
fFXJLs/r9YqMI0P3zsUKaSWNAnmYMa81Q5mN3+FhvN7JHWgQZ4z0HB5C5UPvIkvi
J48hywbVpPun+mmSFZzlIfmcbeKAYTSDMwUewBcQ3uR0geSwha0AcBn/VPrdipIh
cQlu0PwrYHB+InaHPAb3eWmnkxVw9gz96tVD7an2RHFq45UrI85GUnHyYYiNQthV
YJ121RMjT8lAwuCMoNJGRfrrJWrpqFEfAz5B9T0wtIIhIPnd6NP4LlBiRI5ZACLO
dqBC++A6VufaQLekmGnfJbD2fRpazUIQmzrxwgWEYXeveYDFkX44a70ybvhSyZg9
efs8IwzbZxUekdtDeS9f9m2w7Z7YxOX6rd2VuZZf5H4KYaOSaU4DM6QAEIOZtykp
uxiqagt+UYIIZclVPYVrSyUl1B6AruwHcdQeRHlMH73cTb+kzj2KYtotGY0Idb84
PsTNpJqDhZd8o+SWZ6Ero6Ja8DAqvI79piVZfRgsqIabj3CxFhlgf1+JhvbB6YS9
PYq06wxtX3+LrEIg4MhmLJVnAKWxjDl4XMEbE0OXX+mqrHLCzRAfxx0WJkvj0DZC
kDu5e4Qc6o3vxe3iPU30CJ/EKdt2GkracYZ+ghqS2hl/U6Akh+ilhyalWoOmh6XM
BEQnoPq63n87JjcN1kPsIoZe+AcSdd/LeglCOwDtaH6+cGCNJ+zxGgP4rqlJWvaF
f6sVCFXayQEzYg8sN3G3y1iIQLlDYCod1iCNdt/avebLa6AxWO9tB7LJO21Jsujy
jKFe3vruiyQYKjBr8n0T9s68RbcBC6BofovnrZvOAbJ2esAAT9pMbeg5hE2zujou
aO3N80OdGUh2crAZtWyLrJuTQ9bJIc5A7tNxNZrlGwIbj5u/6PsdIXiF2fdvy3qL
zmQKwKpbwjNv5dqSX1k2hf1FPhcNeoQzG44gJcb355gK7ZT2JOOqWGRZtcnaJtuS
rnx7T6mR+YVFe+X6CJfV/zxUWltw4zZqBt/Pmhw0SdWlVvXEHTCauJhmf6qHUIh+
00OodQc7dzLUKhmnLAh/y48nYXUqNkqv3cocMhptPymJRYyyKvbJbf9ONcFulPjx
zqs4ODy6EKg7mlfAXre0vhLYK8v55JWGz9kmqxwpz5pfbUzo4NzA3dqfJYhaGzeJ
kO8DM7YepNhnqegszIdZtgTyx39DrKtx6V+zO65JMNEApTKWbp7zliITJnFx6JD8
Nw1OygeDk7YPSPT0vgMG4LOk/rB88fV3wULMpnGGIBRR/MlSbgRGtmnil8meN8rr
UZXgwWRqw+6mewkT50GFocMOW86ZDSOqBT84pfvwHHGtzDwACeLNhThD6V5JFBn3
0S5DDATgdfm83qaqkzUcNfHKScB5WBxSnAcPt1P8pHAUEP3FdDzkGE2IFoy/jTM6
8mJiTEjL43ZUxtdYpxMowYxBPvjImUW08ME6eX7IwqW7+/RZNXihq7V/NT7f9Wy5
lJXKYhuZB0337BAtlzqBBuPvnIdV3U6N3jgn0Q31J3LSopcgHkFiHWo7UeaDVspk
xnXSlD2ign0zX9gAXNHY0IMiLb++pVisL7aO85Ud2gmFC/9qB9RqROA70rC+pgC/
m4tIeM1kWKOjWLbzRoeTWy6w37ngKdFFTAjNDy/OkDFVLdknxgJlM1UGNEDJIEYB
lfUEPQcCRBUMCnkQp3uXoNKYBeoHjaHav+8mtEcsXHRpCyiqaWnZX4IVs+v/K6Vm
gTJZAQTEIemtn/7FYzxFGaWGGLjj52J9BlJfjuOX9bV1i/iQ5ZXKS2p+RKOkLyMQ
0Oeid5nr2SSPEksBnwtfjWiLDizAm/4CX7eZLGhSbje6K0biVI+XiJNHbBWSAiEK
AMk2romcn0KMD7hDD+jAtzAL0G/OvHEiAsW9cKrA1CudPb05teDqXMn6qzA3FQOS
yYU0LdKOyuxEb+FCcWc+9toYlIm4FtY+x/Mmj1Uy48vi/LFeglyZeWhhrLchWLWF
jGT+0PvOPjPO/0nDnEKs1HsTw+hfGen8rIhJK/HkCeLBdPwpTCoSaiW6BNn0vgTg
/MvORY0CtJ6Kn9+yjej12+ZmE+Rkc7BUjp9R+LPTHAm62BUTVddLsxtrkWpu1zA5
aSTanrL1zSPhtHqwCpoSf2fGVIJfnqH9odehIWWLv7AN/1Fk9u5Jii6u7XS0o0PE
6zUHAyv2FxwYfCdqJn3Tw7EqC0szwxL+Jqhm/9QjUeFscOgtEGcfY6iB/li/gGaY
V3/oD+jeO3Xo49gOIrqzrE1yFpD+nQ+Z15WF6ljHJy3QKQiaLN7nb9zQspZ3Rhyr
tcA9u8P9dWxYh3+wHcU6Dc7OrCMOqmQaAivJTTmVhyfXx+zYM4eJRu8Dwky5Htlc
HbUghvHMjLpWHlY93zlqDR0HByQLzBtNDAICqiFuV/xO/T/lI9GIhKz9ogduh4z1
8yhtiZQTbzbu2Uo8qk/3GdKsSE+foZKRZUF9d3+dCCvs5O4ZPoJwEfFlN/HjWlxw
OA+OCbYYei6yYTJCz0WynkoJRjuEhTH5sz/F+7q5oqa8BEMJgBl94cA1gI0HrDKm
dHLCyG1KUeiY64+ze/hYTESD7YOI3LO3F3QBz87Va0AW6qtbqA74BXt3s0jHwiaB
IJTaXDrHkfJBr5yqSmQhetbFr8smWgb6vnhUcM+ZTApKvjxTI9/pjJVuG6aVOw4t
BCv7vHj00pLVdb5AJOB+p2grZXwFv3hlOYtLESg7TbNrR+soeiKoWX4g1OWhoY5G
l3Ec8MN4FmAePm4j4Zo42NUWJvjdJaHjwZrjREgUNuXp4R3hBeN93gtSgrjA+cJv
s1G0Nvjb19h7rWEXdne22IzikO51zXg5potFJEoljJPn8h/0ouvCwnkzAI5cyA0M
Y+CTsD85ldXllgM8NQykpwC2agIHWMiurPuyaG7LQTW2hDYoMxbIpaL5NW0nYrU9
GRE+ffvHOH/T4Bd+wJwKgZxHFZwRhRrWoTslhLTZ4sht0KFz9Be/j1+GGOXLXvf8
rBviBASi5Pwfo0Gmun9m7Q43WluaJ4yUCwX3Z8LQvTwkSUw+4ic0kCgMtgCR8tvd
nlw6oq7T5Ul/RE20ycJHT6rizYjy8+/Fhuw6AHqFC+pOl8G+jqpRagAjABlE4xbk
wmSpWDVKi5mwp4XeDYOUJXcibMZTRsLuJmgZpu/zuXXYP4DpyBEdZpBbr4AWDE7f
zwllq/kCVUnGWV10DP1s6YDODrvWbOlj1UYuECgWPA/BavCfGb+Oi+VeWIUbD9r5
FhcImt+JJeVXA/ORMS0LyuGlXb6Y5zmeONnsLbT0SsIru90qPVTGBgBZwOl+xdY6
MzOpK5F9xEaGKdD8XkWjWW34TCEGBXSwE4DD0S0CJ+ByfWc5xQzDqe8W3i/REes2
bSCzyq45D07MBFveFB9QZ7GJpN8RkHSBnoW9na0nfeqg1evqJXVY3o5u3tWARUJq
32Tnjj2Pryq2kTpkP1pb5uXC8Db0Vpr9khC228SzGQp1gdVe3EDXM6ai3UULG7dk
Zxmi99j85OVD4Fx0kk/DfrHqZErjqX2shZdhYagx/sJjv5lLFWbL6qEUUjGsraTo
9y5iZ54MS6c2sxC7huWz++Yqvgq0RISsAYd4MHLt4GeSSO+Qtg8eK6a7hCn2edn+
Aycf+MLU8TAldbfKzAv72v0tzwMiiDIU382MTvGn+rG3hvke/u0N2gcM1AS6po7J
2qqFnQeieEkel3065MDOVS/iH/wKtSiOGWOMVSveIvm5bATB87uFKFXzfaFVV4AW
LeBwwSxQfVaI7oSFNKeGZ8MDHUverC1r8HzIrMdoxvXKNsD24nAKrxDZ1Rup3kRt
hRrZQ5Y5I+d1i+KyeGlMq4m9tFW03x+l8SGuGzn6mgSRgrxeggmwkAA6peLk3CIW
emtBDyBmeZ06cmR2BlNtd+QkJegJoigaO3jHYGdtO5fK+bHUothKzsrjEwbqADY4
mnQ10wjEDnifV3bdPXvhweUzZr+ldF3cdFQPbGZZfWwziu6OgCjetYQ+r02iDKdP
/WndwAzBbU6P0ntNsqk1T15wJuTaqxSOXfSBcl1Ixo/vzJYq3BhGUJ+QT1kZpYzQ
UWmC2JQ6dhvlBeK/NsTkzkmn0t/XnxdxOryD6W4J8bYpEOyU0khUG7rePK+ZIvw2
knF7M5CwQ+t8qNPdoAtFpA+4iQ2JQPAL8ZH+dIZ2/iDKjtzYhP45ZVV0a4GfiYXQ
SQczPIn9JgEwh7l9Jv+WbLVmGq8MKDPtWcT3mLSftp+ndQhYwAgmCuAMzoSvcnxx
y4SKKrm3dhi9hlJwUWcSZQs+qsmiRUdzh+GK4XriD9dp6KLqRx3yyJ/tYXxWm+57
xUJsFKTu6yxkTEv1BO5o0PPibGVYi48Sy4fQ9nceGdrlTFylsSdbjSzcbkjzsfFi
+pKIouhFEKJE1X8fbsm06h6N+AUTw8luSFK/90nIOqhas7Lgg7DNWslxnfjKgr+E
VTkVuAfoOfV8aY1w4Nbid3nlskkySW971aSK69Z8oJdXbbkH57XLyihKsjU6wJNU
LVphoxUJb8behvTIt79/YRFdc6LCiEbRBzQfpC8jeUwbt+oZ+/gSq4LY4PXIFcz6
E2c1zt92dFDbjZyiavGifSd/wwJ57+hJzMMwRYGMOyDSavIFKatm/ZBMwN/ZS4uE
WOJBK658IrC15prikZXggbdem5wl8/ouZELa3RBk1GA6BnfjtRo9LDYUY8fY4T8h
hGs5sZJ69TU6VKKOVprrmHIL84SgYWhq+WH1H8l2/FTY6WlUszCWuyQTcgae5lds
/otVeJrncZ6bLv5E8UZtm3QXch+Fkpm7yjEkdMksI2VZRN7uewGovHJfjINr0ciC
Yt6ZSxTYgc19p86392AGbEagi0Aylu/I0J6M4vk3KvfI3QQLA4aClJFifNslOGv6
6yo/QsXxM7PpSyOEloo+qudsT0jjA/ezzPptUmrVEAcOFYN/qS3bIM79rw0kcpi3
1ABjVBnv/2XGYsGw7WPA7Me100PDvxVjJ5PHVuQNXw4L7bfsvNXld4CwjKwIBHzl
VVC1+SBxG6ziutOXqKZA2t7YY6zFZwaOdORG/FFPx5ggNK/400w8QcavqlSVdpjt
KF1TQW0t0H8qT21hVHl2/TNq5xc5m5H2EJ6cO7KdB+3OA+4HkAlj7osBKQnikAiA
8SQLmVGR6Q4Nqxl3RojjkrWVENZtLyT/f90S4vT+sZPwvJUd45HFAgGlajPU6Mqw
kgKVq6tGL9yxb/ok+1zZMJ+OnOGjfZGTlOBZAGuPoAe875Tkec+qE9bgLyFTCTcm
LMBydLdcXqwrIRBrKpBkzIPLy1proJ/Le0rpTdqwfgWNAoZIOoE/ZwXO+8Ekm99T
mFXuleQOIrfnnpuwjCBjVbqN3LcX6kWeP/L2B17QAVXVF9pfvzI7VZ28dthvON8E
meBwye6FrKJNeB4wWDd/F74Z3XlTXdApXj0XQe+VilUP9/zXs4bAwKWxHAuKPYD7
t6pj5eb40/ixzGnGpTkWQ0FdCKXv2uyhZkm3zZCpGe6f3xbyLfHzewXlQrW3LZ/1
03NmiX/Yza8yR0b6ekKkX5wjwm2IveXetK8VMEHSATvqY1RVHz1r24fF4omimJXT
WXImN+r2G+bFK8UPjcSREcJodIw6dESEGfIeZpzz+qnofBo19NBf4NV5BU79XKWB
aJmOel9PW7VanuAngeewmwmP1a8gg+JJLsOU8qaKUdyYyW0Rgz1+oZzM4n/vzC2m
8Z5Jb1dovPf+t4KRneBhlNPadkys3PyjfsfcXhTJFioaQY8wXbqEsWdxnnEIDGTK
a1NXU3kb6AXfP0XTtXeHVrpEYuUVGnMvhu7LV6KP6ek1pIMM5pJjD14GyxlCGTpB
fzhUAJ3Dc+0ahaSaxZfaQGrrRpgE2E+SGvQwg/5WRcGSIengaUrJSoYtLOpCmnCL
JqeO8Sbx8pN59XvoTs3/H+lA/+VOq4xc6YhTrWTnhuSmMKIHeo/5ziL23KwVsphz
2WMQ85rMLIvoaJXl8t7MM28jwLbr9cbpfCdKtijxsO3GFTc0uhOYeYYj/m/rLL/a
SbWXIUh9OwMCQO78NmUCIv9Y4UKuv1pU7GNINDv6bZThEFRB8lm+DrCsx1T9FZf5
KslxTqqF3OJAqm0e8+eviqbOBlzJIYfqIiSjJP+ulzTpyd07WIe3GF3uUouWv6E+
ipdYjFyCWEQELkEoeny9Dc2w7V1xK6hlZoxNQP2JkkWBf6CTsfB2jbVdLJ9Sq3gy
fAjc5YUgO2QaM0JHREsDihAbP/bNfi+UE7OlSTkX1jqjI/bgXY3wTWjT/VyxyROj
aTh+kfvVfbCjaoHmWXiI8Mfsb1IxizB7P3iv0KbhVjRH/JJ5kFhSAkl5SQmzWpbo
FgXersid54U132bQsuMmohIiMBPge8vYEWf2LBFvyjEMjCwfO0HhEi+R1p1A2aVe
UBUMd8njKrqr7qG1lXAzuiGzkbAChyCl4y6FKnGvVNwdBDEqXcPEn0j6ShZYfu9y
kJ7YR6J3rz3Jd8O7ZvRiNFJOhO7Ga5JuY//zxdimxNlLIQRx/qpdre35qKFYDW4+
I+Sam3VJe+U95ehwVHkv1BbyOnj1NfwB+KjggwSA9EfFTDJJuYO7U3pbNQTjep2Y
J77AKLtZF3aTKL9unyyrZOKDz5lkFAx8/tHgQxhHpThMXgANEy14qUsjsISDBBWj
1K/ysoFdNnu6RNNnqUaLrg6s1hOYFfSqxixmVQ4qLEIzjKJpekapXYGp/DCbsPxR
1rOWBpguFKyU9HVKYEdtxD/KxVY5zHBa3e+2Z/0ndxoYCDeme9vv3727E9/lLLcC
BeOZIFHjjW0rpqMZ789cWf0k/Nu2bVG3htsa3BQAKt7UqGyiE2XLnRwCmuA0tQC5
m87M28fMf/QUFYOD6iAQVtoEHdcjp574et09mkXkETkSU3QQ7ykv+XwfziUSgoyL
eI6lNEnfm8H8GBuNTI6xvUj/+vzCyVT99v0av8+CXMjA8WVY9WvCIgrcajiP19jz
7cutTVFXCmzsefi16hA5nhFLm+N00MT2/NjklvJGLYW2BtZOesBVh0k2b6sPrUAz
7yuhRRwi7HHRxbLv8iOpznanDhnUZx/QHR3j8zk+raJViAo65o2a1yzUW9oSHAh1
JkhgcxB8rwPigQ22pDVBBKG4p+B4IlM/n+OkxoIEa36SSLv5PeQ9UxE6q2Y09TJh
cx0S7ZxeA/h9NinT83jQGj6UgIjtDd0LoLaOR+CxGY/1n4iXb2cS0Hne2U5ULuHV
b0tBPM4yKtlVnQAfZo4EKSmk+d5H1b+w4AlbVVPUMYYWP2np4CJkSXaq9viZ5w2v
oYhkbW4fURt8rVtxw9eRA/aBd7SMmK8vZn6TD4laNPwd4dEC8OLUzEYaaw9BvhbO
/aLXg6D4ejC4KHeD1Eqn7InmLxyomE7MzoSZCuyK9EjWKxrXHhGL/ptEGf3Lq1OP
qj5GcFaow6e9vtCdeGOzaThiWlhAm4cUz3oGv0NsumYsMJ7N0jhfgv/FoEV1Jq1i
Me0qeXDqR4F+5BwzmZ45KL/JIhBr3Bj4K6RRUYwdJEo9OgHYm46EDbBX2NWvCX5j
DmhrTzFfYBbLVNOhrVp0lKDUPzqaoRQ0qfUoaJ/n8dp6juNMtC41jn9NoylvOf4F
+Wx6GWR3KLJfak7umIAHdnrcbW7aCH2QCOESHCMtoyL8cFrCQ/4zOxOZMDPjNxXj
9GTzcuEvomMM/q2NBm+cYRsvm/WAowg7BaHnHl4+GdIyxamvTLnpDjfThaQV/EU0
qeCAEfEXKiqxoV/x5z9ryHgsWKdTvrEty9w3ik9EYnB8KHb/2O8PPODxdly2evmA
88BIGbWMLxMw/1erxmMLWVNw7TWg5AyKYXKN0SN9cR0XF79yMw+qur6EDrykH39N
xOK8qtj2IQvXmNgIeZsUTzVoX64rx9BlvgZ06Y0VjhwYCAy6JB18GfOuQBBCAhU3
ZclbLgj9fYTnoAHHg8K8BDVOIvCu3YGqjsraeJG4z/O23UPJSZbGcreVB+Pd3eq0
lrFLQYE0i6MhRqbfb8xv4bWvqNAi9EkYP0Xf344L8sn1hjNCA6WHG5Eieu5nHcv3
dERqeuOtXICR7V1xGpp8aYgR/L7Kf/eN2gHb0dP7K6cr87IWIDbbslSvlii23rAH
TYC9inRSMHIC7II7eSyORvKWdZztFQOEXzmAgjg0+Fjl/fZImkFeW5Iktv1C+odF
oDWhPqVydjGKQgzjxTHZu99ObQ5Oe6OmzSzWp4XLodjdzMS9e6lg/TGvyU72Wbqc
1rgyA15Ye7zRJ5mfXwz6MHn/W2jiDedhzvTUofB6ItlBD6SeXSmtgCYACA9wyB4f
kFxYJekLxDuNVxTGOxribCUKhcUeFPZgUsfKaL+Ei8DXlCass7j1jOIu21MnLOzL
Goi6O6vf2/fy8WxP6gDOU4Ywxems+dcghB9MTzqkUyhachnhIP8G25R8sN06KTCl
XlEICZPXIWvOGFocXtBCs7wEqMXGshEygqj0aOV22cSAC1II5oVOaKDi1dUYmZvB
oX1UVtFhIM9tN64NrgZ4QZd1/XwFvM8y5kMtNiNmA3PHuLFehZMzuU1veP4xqAdK
WtpSYktrd1ZCpDD9XKiYE7mLQWl2B1/349/WopXh40fpP/Naco8qaCm2/gXajGWR
TVmNjqIKvxkP2i7Sy8/ipkdE9/cMfb7X7dcz/3Gj492+D1het4mAxoqZ01zH/taT
bmX3qW62DHhuO0cXM598MsfYSED++8i8ZiLT6aGBfdzL38AlB6t+8QziVEHaPzeT
x5KRqTaoC0CXb0W9QSxw6yg5rO2dy5AUXVYFkWy3PTQ=
`protect END_PROTECTED