-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Bn+e188ZPK8lZ5wyzn1QPw8v8v6rW2Tdn+dou/KCkMcwVxx0CRh43+k9REx/cjJz
cX7kVze8ykMTTLDOiBJCce02cjtN06mV4j5m1m2KM3JuTijsu/4fORwrPUyH7U9d
MQmjMwkYfoCt6ZdyNMeNAAsfhKhB6pjhCWPmDxQwJpg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 190085)

`protect DATA_BLOCK
7KwiwLtSD5LQ6qlFYrBT5gAKMylbnlL1iFauj9SqmS6wUzO5ki3NULqedYgMeG7w
L9/m++PINRT+vx9chnKNPljFBRABA6nlJ5ZB3GAttx4cUBEYRvlYj4bxLApHbuEc
5/LSiVhKnIpui+xVc5UYu8Q3wg3NsGR+fUrNfDvzICmdQn6IGN2bbJjTHMt2d1my
06A1vToXwKBntmFRmdbpg271i3s0maCgPH/Fue5DtYazYcVQz/pf+7K6kaM7CUlU
vU7m1d8i7bj5n8CgZ9wjdAeYDEWurTACM2aHh4THW6CAnJKp/HwjZOskVSjT8EHZ
kqGpBaYhwVTQTiT/eaYeroDLEMog+M6D3ESk/CbaPSA4PucJTZI3T9d8kjqF7b++
LJYTnXQ7b2vNc0oXhOBcaU6yI0AyksXsOSDZsuYM8LLPsA3WLzWLBE/OhPu3SNdR
EFkdm4efNTlrrhlvJq6rucpsZj2ULYM7W8aPxTtpikdOU8kZrnjMG6vbFAQJHSH3
i4OdIzDzt3BJ/1GJiOl1dNfFB6OMg6xx3gAplX6u+ETrYurM7lS2sFeq+zbP0l8C
XlAdI/JWomeZF2k/f4jgJb8XJtBrzNTZfdTyEcS32bucfBw6FJNzd2D9D7abX5Vt
72UqSYVeligrMxJWxTuoVp5C/+dtXyN1fGxlrAyCvDN+xnCjNjv4LTWzne+rOWHW
3pGfJNNVHSjupKIgigDub5YjNRdasROj8ztfTE7C2+MQ/BJx0hDmEO4kEd+GE30o
e91A+/jNRB+CqcArATf9Zqn0u8CWx4hFEO6s/0JYfnAeRDEXrYGWbNe9TQapwZ13
qeFyRQ2RjW7YFBDxAo4jL3XE19TJZZtg4BDL97GJ1wjRpeh5TkoR+1kJpQg9Jn5H
6dSfRshT9BP+b/WwbTbOtFRwCb1lnYvpTwIEt01PIFIMPWeYVKR1FtuxQQNVHh/A
zng1dQKerFSZiBhm/KCCGd+bWHdQt3vnGjvA199DApn6EswQU9tPnRM0dAGX5XF6
w9uvnpPH+lq61MnN3wytA4cjv859M4AnVN2mIjAJ5mh67e1Su+6FSxEb/c4R2C92
au8jvlp/M8YvDWnCmAOCiAEYfD5+eS69zi4lnftGvgXWoG5EtQ/bOjrYwyT4AXWQ
J5IWcdkLXpqUyCmGUkQKa6uIgXPPRvK3t5p/G1ykGwWu8LCcxhMQ5UVekJ3vTmti
SdohDZq6YMluPL41IrLceBkf86W/0Svjc7gH6l0gKl6dY2MWmMG1Y8iAyvDLIcu8
0B6J2fnOz5hY4wsTrTtUofVr8VMJJ7/O4SLrJkgwYBhf1/+ifVX88yiIfv1zJ9wI
wiaB2JjnNXdkyhjjkuO25SPnl17/bI6v/3IR6b0A65gI/9e/Ih9i298YnYAxwFN4
lPnfvqL4emxSOx+kPrr8OG2F5mgTdBsnvlQG3/Pe5wvyBH0vZeVU7RKdx+F1RYGW
Olf5KbXAGEolqXCK2D5Gd5s7UoGZmS38CE+mHtuHH9fItPI1G+yuqHrEbaOKjDlH
5XSSo8nkecQasNF82W98OUOjeAO1L27gyYHwhH2YRef5iwDZ//YYX5LZzKZzIeDd
AcQ7otds+J882g8x66IF4Gql6/vWXawPZhW2bF4soanYMC5ki/HQ61qju0bl8JTx
XDUCfNFd8qStTNiadfKw8pHSssBWQC2tv4N6IcN8dAOh4OzobuHIeXtR12PKLTh2
KT6QuPKcBacjiN0LX45bIK6OrT5qWNDbznqHS+BrpYbsaFnTb6wsJf/yIreZHxCw
vnQsy/9ao1VvBdWrPBfk654C1uwzjEoZq9j+Fo6cIrNB6ecAP3ABKbyaKlKBFQ2T
DuJoeXlf8yQMxKDeOt+M/ceWPRtGy6EcLup12346JxqMcDfijO0r1ktBGWgvfWNf
cs/s+hAcgaQs9sNUO2wXMCLIbNtdVRiOtahywAT4uJJQPvpLpdpQsrnPuszyVFjU
1gO8Cn9nCdoeS1pTJ+YY3IfeAAmktYitDADbVQKXzhsIllD6CgKALL8JfDg/lk8T
tIAev1ARQCe9ukCESn7shnA+sDKRRP4hsEO2WlAZFE3l3weYpLMYlVwJfIYs7QkI
5H2m3YPT+kdwaq1OUP/+VgPbB059WPy236k5jzNb0N5cyAiPdFq0FJH4DI9Rhtkn
P8f6+L02uAIspbtm2kuluLy4Nx4u1NaAfD9SDlfMypPJp8lx+3EkrUtnhFi4aKrP
aZ4QfeccMKjWrvXGwJo21n1eJIbq/dsD7Ng2R9viSjN5vcJDuz7vG/ONni2KIygx
TKQ6PaGDdtcno7FIVBt/3CRUlq28XA0vVrX63pLromw3isoW0J89Do86F56fEtaB
yjzo3E78i442uT7UCBAl0PLI0GFiccs7ernL0GwC5r0CBEs1qKwi+EAfiTuGykJl
6X114qYzj7LcSiIP6E1hjerAX5NwYasDUxR0CUri/9DeOQDPy4if09rzYIMS2llE
wIoRv3L5N1P+meqbgPmNONJMLgSJhjJWuhnDCfoHGQkqvxKAM5VC/vZlr+yD6dDn
zdsUA49LEEZmMy2QOWgPsT7Ggr+di9derj9lYFTC8QSKlPdq1Uwv6u8arPhYbiTx
RVYf9J6CoAY4qB9DKzb8UYN20+s86xHwuHolDyq7k+QpTWKRfUzCRw32Eoi6Ur0t
4gm5Dn94LDTozlFAH8HryHw/NQAvV5H22k7gfoNGAdHph7F/B1hsunlcCpeOEuF6
Xfl0CbDuhaXwbOIOlMY5bvIkBaUy+nJ9VJph4/VcWDtg3x2f9b1wkVvoVGAgwJKu
tB6p9tLAnBB+Mlxv2TVYWmB1GjNDlcdk0k1R2OTUV4NbT0j/y5EAHvpTjVonfBc+
xgDlrURPTmBfPZKRW499A59GCLkqJf8EZgg8y5vTSW8fHz9QsMd5L5jVSZS49qBb
hzHyLCe0JzgaryvCMs54f6hoYTHgZFIz5uwRvH23B3PPjpmyZ+O1psRVmOh6Th4L
HxuIOYalDL9jHCrqjKiMdxD0jmd20F2014KLavhsNKnhoMyGwdAT/TqWLHNVAbVa
lvu8cXsH4rPlsrvB2WtP6kSxQE/W1bHKhv7K5lneZaSSWIt1BIB1ZlV54TukVMaF
DImFiBigKwpDAuPNnXLqTQMDaWukyxpyYah9pHYiVJR1s9GEIttK5CA+a+PQoBij
dkxR11MQs4E+pTYtMG2LpciQv86/yTuBqFqC2l5tz1DxeHGAR+hNwnJlWt6+hU2w
4X0d/97gOfd2G5Xw/030E1yiiBVXZYh+vfj6miJvNTw4uQrm+LGpjOg6tzj+yYOI
jMtHYtOXdIHmYrloIJYxq+CUhPCBJhC2JcPW2zOhOBc/ylAsPMgdaNB00t1vBscv
35CPQAdfUSwO50qQpOaRJApMOu1y0RFHALbh/D4zNsMrxcBC4K3TluNDuvvJvkSM
WSMe1XysuUn6RMAetS/UDubuCeljxFG2VZ2lY9nbuxCTrJOGdULAvh9IgTE+TlGm
dAoqULj1NPBk4ZiCqr0EQ1jSLVaeVrhEamLp5zIQgzJOHFL+VAE0Lll2QJHJ8xXO
kceIM3rlwwhFU5WH3iyvL/iuPN/FYrcvHz3C6wtJunV2mLvnRVzXpo8dLtVZ/0b6
QR4qXcOCKDj/0YKnRbQtrd0S4R7CKVB2e2v3ifNul2owp7OIT1CjNW3NCqBEqUnh
7BTWe7L6VdX3mQ8/H/PS+HnZPQmaShnLASiXQJUcoZghHaRndiqIZfLsJBzl+jh4
jAQPR2tKBHkMhWDOkypbYnCtoCzSkUqYKktEhXTiNwmK7uNbpeFv6nd4t+KX1i5w
vt6glU/bbE7iwgch2tNwsFL79qRW2X0Ki3oCEO2WrDffu24BgACzQY+AO77rNNic
YpplQw4niUsbPAuHaYdgPYd1akshpdBRc/re2gEN3EFZghdQSxfJERgitYRkLhik
Mr+nLX7uSqM+l25qacewcIggsy/D5+Zv1ZTlKyF1C2lgIoL2XJx6NPznt82afm81
GugQQWZz0N4yL77AdQYxYJvQ/Q0sOKGPZozmdXK17P7muC7krHeDeeNKcaKyO0gp
vS5knLl/SsveBKHlaViTZJ7BlXsbompcz7NtfwRIJrGengAW92szYBY0rhnecfIs
caBMfDA8CcU9AP7791KJAiEjhORKTIZX1QWWt6qKML8yP4rNlHUwBA8erR/lpjLS
+HZpMkpCpI/RSWUFyjGcF827zlXnw4d7p6CskynLncz4k9aCbZxUol+ISX1rr53v
DcmcYls7Hw20Fa77Mgix6GF4TnReIUfhsSFAcLVtQ3XuYJOHYVD1C/k/a8gfqO4S
XlKdBXkyKKKw6Isp8vFpno2LTz/AtFa4US2xWQM7wJkhzonVS87zLMv4NOkK5tTV
aLJnGgOvYM90ns+XDDRA0ppis2hn1YvtyMiCDlFJEgCE/Rbvu023oqq9U3oUqQP1
a37PxxkhmChLQTjkp9bq9PMQi+aBPWfF69ps2ssQ/K0DPgYJaR/Az9LX9yJw2EKe
jw4a6dZA6Q6OaSiX3r+ye8Fid4wVDm73QXU0Vgmr4LPlsJrVHZhgQVMxijZdlbQc
+b6GjGfbhNfbu0lnvHREq252QIlec9DY5p9ABfoYse2qFYceHFehqx5wl7iN7o+z
KkEYpo3yyIQ0bT9ISlx3YFqoMv/JvkVV8BaTKEWricomq/s98vqgknbYIR9NLtKZ
b3vGizTXBnQz+H59nMMkPCJW7NHkln4TUhty8x91t1KJ1ZkmQcdxtK1TwTPUNVtU
WxVAsFae0bXcAE7jC3S/23D82kfFOnRXWtJRwR/7fQlz6JPeN+TX7QhoNHpzyRia
j27Y4SqquUOFAtuxbTMAC3XoRH8IpmPE4lmhPnYAJ2JFAvAlNvvGXttow2MVQqrT
HvxdxXP4Jjo1H0Wnju9m5L4d+EaCGhVktDxzolUC3uuAMtEoTcwDix4ZptfQrh3E
D0bcVlvYNV8BuktVO0SeEbsNxpJtu7b6oQLV5y+N7RZm8rtYJxWvBMJ0oHrqRLGe
ZWtDWiBL+uOOoDskoxw3OYIJvRe6lE2DIOT3pcmt3nPiCh+OBqOovbNGZ2r4ZGH2
+pht8L7GX5dVSO+MyN5FfwNPtEafe1yflOlTbPRF/WTCagG6mgKCE7pbuzobXd91
UJg8BxxDzQTjnLDEFLJ+MgulfYt+Vz8nq3n6nZY7VX5DaVLzAo+yTMmj2i6ADFg/
Vjl2iqYLJUGxDKApJEzLLkPdVUW8Jkl6uHWPqM/H55ZUEiQu9BymICkjp+vlHvGw
rnGwcORjnSMgc0WM6SHTQY2BJvcjuamcND5CIJ8we4JXIJikfi4KQdA2PCTlCKHr
LBEJzPalAGDVxk5umgZSTlEqVFakwAeu+8NUhNy6lRI0myCi+CAPyBXURVQEUmOq
AbAdz//tReilc4BY/cQk+uipUKV+amAhDI88DvAl9JOL3bupBMK2B93GQ/54Lk8I
WeEY/YRWDq75et8YGtzDSmWS9FqAR+EyCpIjwxl0q7Srrvs9w1zOzCN/ue22Eh72
Ej0AwyDs/NcpOcaOz9DqZCJvrxijNBR6ptj/40OiG3qZHdwMI83u48H3FVE2Dfko
CLks8xoJMQYDxRJJnzx/PmoUwZVRwCl+0nLNIg4SueFtrMjIG2Vh/zEBve/kagte
gkDU5iachY5Yw/bHxDHBp6p2mod458IisTg/6L0iWVB4GZ1EoVTVZCmASqUwZGXO
zVHzT7eh2r0GW2aFDThwxv2rost8NnwZKgi6daOtgczmF5wdICEcrMxuO9oufmH0
q7WJmI+mDDvQLH+Z2VIZ3r3y1OUzMqbKcMqpRdAHfG89olBcHEXSs7dwFM/cDH1d
z8FZ1F2Ni8O6eAg0pnycxS+kKVMlpVMKGIQiWqI4g734wAnvT/7VOwO0WYInohjg
AIqPweZpZH4TaL4RWCroMXKAR/O2eNxb3t5HfNVl7GWW09RbOa/8YuiFb9J66ytA
dlFm07WjMw9xYzdg+qyWFmHEJ7j2M+SZ9RtkYD86xL6jic6HWh1uwSgwS4OB7QRi
v88G3Ko6IQjigguxgXm5TkD469DiaxHJtrEo90C/2lGgk46cwybu9sbzns15ZmX2
qLgRrAXBlfH0TARYY0Jle5L8ijw2ehxYqfh+BsVR+UD3yp5k8wzU82pIu75MlpHX
fuA5h27avRbfrqRUEcBRBpJRtKIiLfCeNgUmcp9Q/9doNZ8QlPvAg2G5UJDIPKGv
jQyqC+3UOvU5LAXNpl6I40DZ2BfifFEDaFcfHzEuepRrzfItp3VdBGIjYX/RyGDf
0udEbgwSdoEiK0rOMINRMLpUaRmr5p6pay6g58PLq8+H6a+gQUp9+B9a58gP1i/u
YXCvoOR9lUP5rjFZzUNbbonbOG8OhK6jzrwkg5nztchvOvup5WgnAvYegSd9JV76
pDAj0wvbWGVwSttBPZNzn/L2a63tbgf3dNmHeOXkESTxBtEs5hN2ZBQyq9ZtUcLF
6SALay0GyCoFlyf6pkNVfxUHvq7T8hUmxG1lWDlxcGc87vpQp7ZAP8E9fVa55Ihk
AAERpjv2l+lajk4sit0G6hcHjG9JHgjf85qKWAFWme3kBSf61yyXSqIecVcCON7w
U4yc26mvotg2Jr5mDixV/IfjvE26ggFkpEcaWRFn5VSsOmq1EshJE5Slf40vJKAm
+YrjQMU0EolDCdpdByQezguD1crbNc8P/UDCuIDFhlAm/og6MPskUwmNEjdTB5xK
gM8gOs3LA5dAkktgXR5W+XI91PKnozSOOGQuVWam9KdazKhRvXV56aLN20uvSABI
MszNqpVHxkAB81sYiY6/ZhkHr2YckTGZGaKSkm0v0rGHt7aJSQBI520QQZXv7Hyt
lHUK3K10Cse1jS8YJRLeZnAfNLjTfrEmpfI4qjVUs0sqvvg1NvOidg2yxjOudRxh
aS0MY+O37oT4P87cafaYMb6XyLxUrp9ByyX71FldAaE3wRlEOhrjucyLaOpvoc/b
frzr76FPmmw1gaRQz/Ux1hCJAvbtArkc0fgwwU4RNkZ2cxHPj/F8RMl8Voxl6tsH
0hwawuxyNotb4+7utLZHY6OBEtLSGWgtFnZ9iW6V4ocqiUSMlyG0tfo97hAwOq/I
dYwbieKAISmUUspdhfYk4Hf8Y3JGHIml8eYYkEcMXRU8jEMYSqEuWuzWQ80cmuRb
fn3ORf5sQ6q6C1JNQytv2PybXgPAqLoTS499RdGfBZgPF9VRW3tDQDkcrEFV0+uX
RlBntECwL+Eu9wpJJiqsgB5fQ2i5gOVhTReLUYmfcg9PYjT16yYxBUT6svc0mtU5
9fI7h6CswTCer0/b61THAjtQbgz3dxSJr5dfn7h4dKNToOB+hsET/ktl/tJkAx2s
7J60sbmYinPTT6DlLIUCzKa4DW/MANlH6VuHGx7UKhAS7lK7VRnlKLx80UK1OHZn
IDNlCAFx2qbC+vrDtlK8m4rWJ0e4sNuj3YZ5mX3z4ROZY6h3HeXeSvKlhnAwTTx5
UwQUqXpg+KG9gsN/5Xp0lPmImGCPdZFJyVG7BaOOAKg6bgtIoPDDyaC5G7l1l63e
UdczDYF25sg5EjzgfItnnXMpbY/wQ6tf2hKOuXNLhQrMaPA05qD8tSiGyIQIrOND
c4lZZe3en/1ewh/lXc1f8k2ErY+cVoObj3rg+o//D/8XnUYMoa0YdkuyH1h2Rer6
SA5tkx1fHmkJU3HVRbZc5I+o5IbK94BNMXQ9R+YR/ss0PMWlv7bv00quhsuCQGDr
CBAXKoKSonC69UfwB40r8ZUN3a1eWAwRUoATtAAqtX6+QOxqwX8irVBXUtp+0YVZ
A7TMNW2YSiSKXOIhkbgECTRNhDY/YPrBh+AgtMlgnQlSCappJ4jUxvuja4Bq7z40
YmQQQ9YS3AIN/s8OycMLIHVVX0JxFCmhM20YJFf2aENAPe7PCwkVxgBUWF0FblpD
90lzSrG5XriLqYt8zD43o8KlX3xkEuloYB9FCIkC+U+XT37e4acslBV4T4ryshxT
pls1klQw86/8CkjbwfKR36wyHdszQpv1j+KZzoIOksjQBNs46A/0kamkBXMK5zBf
Jk2A/HDKLDxZr3jqDjgfx1xBJPtzS6ExbHIVNI2OHjOOfXMY3Dq5ZlM0EWyTqILP
hIRae+7Soou5NSIXvsOP4F+L7Sq2fLIx5RlX9sRveHZ9ZqWA2Y/gjc2M8DLLGZmQ
QDF2uTFlQFD3JqVCELBre/lKACcJeRfTbq2X4qF0KQJNIc6xkkBUm6J9Y8ueRBqW
PoNTx/Xy4tX2J9bf1NtXSVF4Frri3QHAQ6wNRyQZLfhCzhJpF9Lp+1Pnxi+M+uJO
9akNGps6vM/Nw87I2I8jR0vKt+AVD97XHgibPLleTE4LfaoaQMdwUUEIr3QBIBeY
YSqYdUPTtSwNxChGkCkUQq5aqePmS8NtBmO35YOt1ZTTuRwpIxDNFVKKF+LC4PKZ
+UIf/0F6Wm8BI+G8Otled/vqJi2VTngM1zN9JFKF8NGnleHmsr6893jKhy7+Z3ER
frCalnR6DKXOVxkffSDMWJNAaMLEDssJwWz5VRqAf86GnE/+uqt6BU1U/9ke5rrt
poS8KIJdFjMtl84YjxqCp5Hcl1mZRZfd/nQ2WVoFrcRcyiAQE1Ct0SLUCDemq/QU
JzoVPCkmmNGFwr+pEHBKvkFgGgz0djrhtfAhqFnt1t+DprPvu6spyb7uFVl52OBO
5QmqyxLMP+FxoZftmF1ZdC/kQEIOLGEyRKoymq+5sa6kzgAQhnLJMsjTvtZ3FDWB
zrz8G2IfcpukFEaFoHnROo1uIneV2y6QkHCOSoLxW5lV8cgqffOvu1a3x2zXxzvF
ayYepc+PcP15X01wQwfkotrvyb/v9HZ6+KC1natiMgTUCxmPkCbxd2rvI3dMQfH6
+pluj6pVFNjMm+o2NckUBjd9zvMA3FFDT6F/1MDfj+0FHBQxFZYnio/l6upb03is
gXwhWTun3/n0g88PTTmhLYk43M64EM9ROJ/XcbIkbos1xxEl2X0XNkIIChEOWjIh
xM/GiUUIQHOILAczYjusrsgN/e9aLHkkW0sk8VoJkZM7k1TFDp+Sn9WewZ/veRd0
ihvnKgkM4EcGYSB1l/a/0XpP3dSfdSfYp2RdTfAoXF3eSlg0IQWKhX2kzjz8T3BX
Xtz9zb7Tzwpxi8LO/LDV0cNDgomTDR1rbOw27fUW3Xi4wxnA1TJqVJ+hYDr60zZa
jXqWEnzioBTLDWZ3tQO8CjrqRuoLrP4dPb3HXynzXbU3EA4J/bvFRrGdXJnqmOH0
TuKHmsKUzX6DVfBY0ZAk2vCtAnR+Fo9DnvivUJMf4Wnka0Bl1ScCnqx/5YpId9pt
STe+l/7qWUgNW1dqyZPWRmBmF/XfgXJbaTILTdS8EwcqiuygI1lSHEiFDwVvutQk
QASBbTj5Y1VFu1BubayywCToY90Gzvs8hjPHKDWQilGPoRjd7hoFx1yeem/I/dMQ
6L4Q76x8CioYKClkGbKVfzIss4ZzcpcsudyOVxogK8GxEO8T7N1eHzPHltcplWwi
M6COUjRwq2s9NF6P6HqdtTRhyE0CE5En/qk/b2CShoSiWimqDmd7ViDxCG1voAyb
theqBgvqSWZ1x6z4dtyhEP++Sxd/ZBfzf07bZuCC+9OihpIP6U0iobFrScwuMuof
5aIFntQFz0R+Uh0S97cpEu7zbgj0SeuUpV8BfcqzfeH2NHa0uR2tr60wJsNwvDHe
V/MoXM1C9aozTnj1giPpNIqX7aY8HdIkzWGaR8PpMNSIeZ72wPGEj8EvDKQy870S
5J3ox8Cr6kn5rW1WZqIHFhgE3qADJtYasq5E9zR6PqoSicpMd7IA1aPQvLGD7h1u
way8XUuTj98N61KR1qAkQXpQIwAXRWgfs97TqIH9OominsXDzYjfAzvr8bZW17Nc
zHQGO1W5MnWpd0rFyf6FZNEHaBxw2efI1ITr6OvQVTVKLDFWIfZSRxy40ucskQVf
VgJGQki4DdSjQhH6Ks82c3Scs89R49fsRzvlsGxis99GzRynSIQtBW00zuJ6H7+R
7VsuPHcFobgmGRmuVHqI/kmQtMaSMnIP/LuSewbf7NdHcgap5HebQPaQJIA3zJQE
fDrlS7d6RMHLSWc3iyHNTNenCUmOQ5uIUrFsMtrgCxTWiz9N3S2d6r6gR2gUw9K3
ZXq/WlfPcckw11GEnS1iv+4g4zqDT4HYmQDO3eFK/LomnKOkySwfkZiBXqiKxGKb
xSNZBBuiMxFPMdAyda70NxIYFKR16qid3ijLkQOgVNuSGv26EgtmrIdaegRu0BJx
OmF5vbCYo4Vc/8QomDMzQZMvOXEBgbJOL2AI+EXpNnn736EoY/ztm5dl+bdIsmCM
21v4+3RcqddB3D8HoPHIG4wK0oLAeyV433bj9oZfXtaiWxT3m15Rqz1gZ9HdfbKE
Rd/KIhQNObW30PR0pmjaZT0aUXo/+Y7nbM+L8YfUsgXduRRHW+QUDb6Dpf+0nKLY
6tg0YUlx7uV+Y9SPuo13ynkBzO5+sp2HUvcy0yhDXmoWJq9X+qNNujZPxUYoC+9A
qet0NKZOuSZZvKtB1qOI5pPECgooVBJSkl/hwIcZA641GmlPewRH2hWzuqZelFMW
MUtZAJ9p9SrrLGXiRzzxk6w9EzBUt0vQ8JcMnPdacgwXRMTpEafyTG3vduQ7Cn2H
bnm6h+CZee5cB6A+Dbr1mos8XTv9lFzyUEBkBcBXbETSbr6bJnVuxY5HT8sObPpr
Zczme8wwyMRmt/+7m9rFwXfdBvwz+jIrAr64egbaKl83w1ZTGy6L6voCt1mYYPVt
fOaJ4IZntmfkf3Vy3RX8B2ZlTL0ZbFxtykm2djSWjFC8UdAeUksrEiLkzBNNY3zJ
4Z3bEHUByGUys0AGhnl2QuC1Tb8zCIMDn+yph5NJ14trYM1W1JUoYsK4zI1X0Q+f
om4yHKuDTElFKyWtZy6566YUWalhXY1EnE+/sPfdPZJzHafoCUKWhtXxjA1QxKDG
QBgxnMVwq5aotMcBM1Dygbbasyg7gWGnQX9ni6QSWjoOAe8NlUF0Tge/JHc4SbZH
NF/TIVzomcaK7rRBrmwito323xf6IKwC8v8QBahqHWiJVKCtAvSXTcNMcV0aG1XY
P5JXhBiBquRoYLNXAeumsnBSXYj19D2y1DBKUORGa43FK4RCDXWN1tbO4MbbARX3
1cH+fFk/67FXliLJVQKMTAwfn2TPQB9PoxuJlIyd4wZd8yVPEry9LyLLq/MpAlVi
XJVcSGVWaYxZ4wnAhZ47oGezbEo7WDdJr0mMCwZsTcNaPTm6OWJOz++crAYHXxH2
2bF3zAvyAdAbllV6io4IcfDHhFmGFbPWNobDcBsL5oZZ4RUbhmM4D9Z5Tg3WDrm5
M/nWKxW6N1lbR+erA9I7GSy0JgM155wbM6/r+Fe8GmJ/hV1ECSeOoum4QzijJhe6
aRweSqW1+PsK+EAS4N2rxQUTZ5OWZxUfgpgIGeH6hAnmeaEit9Qg8MuvhN/BOw6M
H83kkM9uU+JNdHs/bohP9afajRkkIzPWGh4moqZz5uKUfBsLCi2a5A7hYw2E9ZpF
MCzdlShrr7DeHOjMJo6N9JjeA2X/bRp0ei6UTeIGw2nbyP+gN18K1orLIijKv7bn
5ktHECqsIYi08UTNImrVciiMNZ+bbQl5l6cJdkhNXVcqydx3rdomf6zOuzM2nMWw
ddx5XAwC0cVzb4sZ85gX8tyjH1mXZ3LkyId5JiHH7eD+evM1kuBZAxIBHrhe+7Iy
zN4SfP1yM0t4VKNoj+retSU1uZN92UrcRDofmZDenF4I/PMPn7guLfX9N2kQis4r
GhI4VsVuweUUmleDnQxsSV1LJxtKajxQjnzKRRz6G461Fu5ut4R92oLt7zQsPh4J
CVmD+ZwCDGPqtdLP7MfM0c8aeEN2PY1OBd4hBiYxjrHdTZyA5NHg77TX6VDxqCjM
jLGDYF0c2RuVvo3Wd7PYOP1OaP5jdnxkANHRaXrTEtUq6beKKbhZ2Z2Q12y8o65J
j1ypSYupxiBjP5dw3LUAbNgAjVH92UfCsW1bzafBbl1c25p89sxpqmH98p7t5sIJ
9HYpQ+jDOkwKA9zQX4EVhG0Z7OmP5w8jlKdK95cedxUWPD5ixW7ms0oLn3LxyDvA
NUaWIozJstRlFrD+QeyWl8/tbRHn95gQNvg0TiVkvb1TuOzlEAkGtzlceL9iYyV+
JII1/Ac2L7KHbxOYCTgUItjJoisZyR5qkJdnGkdomV+5PFrCM2ABZALPLpOT41pe
nKy+uFmEsBC01eTy4SuF72yKqTWajaP1wAJXi5VcyZLmmUWviM+AsgfwqgHIXmB8
5LUZmJHQNM2sUi4RpV3Oc1wqWC4/KvMbALApNQl3k8coVxCd6K3YRJsSTxmaEW9B
3MrJ/bo+bCtBcZOG0kKDKRcOYSCXDKihQ43xBczcnIiH87YkaFyDbIKJYGe6a/dC
JihHTtn7mBKpmm4XOLGlUke61jHakmeLZuqV/3gcA/XPUcgLiuPU4th/YezEw0Ot
2xZ4CZbh8D8GBvbVhyVdFIWFspXKC6mQkGDbc7RG9K2atthLmsKRRuyIlxSzPn4X
/b4yk3xAVOvVdsvWC+BQTeKjV0lY9RRoZoVovxhRrb9p9wWSUSt2nMyzy1hGGKF5
oEZGEshKETY3XKTZKdNfg2YUopSdFAM0FPGYjwEBUXCH+UMkcOBN0FW77uPSQDOJ
HbqbG2GLpDiy2OKzLzjIozmdZqDfwNFv8kRu6WGUMitQ2xoZK/YcCaleCh9pB/bt
b13E1c0Rm6UN4rOiKSIbe8TghEWNR5btxBe0Q3JPjOZN1wZmuQpCP0VsQ5Gofftq
HGhE92bqEyhbZTkCExEiXdcOaGzMggmfmVEGoqn3VtZ5OZbngZ9FSK0295eX47PK
qLzd0rhjFzNGEiR2xy4lMKsySTwRi0ITn/nDMuYgPXmSNANSah76D6uwdOMI0vgk
+JrPaMiVhtcIq/Of+0DE7lxK12P/1BPHZ3CC2i30jlEbK5/57PIkZK2kLRSpu9yi
ie6bCKTGPSnlTT1EB6d8ntJ2uO7/f7m5uECPrjCFeHEl+ARXC1yiVk5nLn96Ohcq
TQlH0rPhpxmehgWuRX1AD9ZylmBBvdxUr/mbNhqeLyrV1obO/Y7JnoOMwH6hF2cr
L9wNpOxwlyflwIRQfuxmjsAeGo9nonHymqYFPnuMwqg3nd5TQOkcOaUsKwj5ZtmD
/J1xAakox8nL6cM4c/bwfccp4W8pitxYypmJGFTR+Q22x5iAm1geNPXVZEs8ugEi
n+ijcYbf/rwSc4dleSnTNjvoQoTxfYy1IvF9OBwVNaDfi2bBUVOAtWpjOGpnSsBB
8Olw5/3oPbTewVX0CVkw0Ft3+3e2krkr9c9kIm8tJYZ7tYPu3yo64XfNRbYNIeNQ
rB1+y2nQN4um6jpWw9eZ0cnFfEpqxN6SbLNkX48ymgHNKWpQ4aTFo9urXOVYb4A5
83Me9/YYyk1WGB5n033On2oMr+IuixlKR9Eh9jzy9E92VPUEDYDKGu0EZTrGgd/I
y3IGH65dQT2sRnVHyX9MoKoge67ji4fRPdGQwYmvJpZgnbeSlqawaiNF4HY205HZ
+gq03E45nGGS9zR+sqaM8QCiE8hFGYf5e6WG40yI6AXd7J13MJgwlWRBV+oSHPEk
nrBN6oNpgZYUe20tTgSEGuvJpqtMnkyEDXzx9A3//3qA20JWhCSbZF3xs0fYkeU2
LfeaZW8EAfUQLBjuDx3kGS2b1g0V+HJmWUF9QsNE6s8oLDtnJCQ6HBHKQOkGFwhE
ANTUnnIa8ZaH34YBTNs+lt6+nyfWcIBCCRhlI7TyvlLJjfAVeoAKV3QWAriAvDdj
3DURfJXBAQO3OrB9uh7mQa5XqNIJNRS+dRjqmHg1okaOzZ2syoWFDaTvyr1prUbF
kPHWxMwnwsXjKHLA8SaZVOXx8K89kDin2ypjnLLSK0ZAz5b6nnEHp2l4KTu1PpWo
vvkT0gGsGFSyZDnR7NkxkGxuI5TAQoKsszVc12G65dAZ0raedI45c8CzBA44Xc1m
tZPo4FwnJEoL7e2MxuxMfEfjs9wNkgmQqAB8dIJfA/PQtUUiNldCe0ZcaATLpQ/I
exp3wJ3h8zv648phUEnmB9RU/9/qwSR5PAqPDUR8Rf3scashMwkH+D4y1oKnYziQ
FqMockP7Y/OdPZDehMfQC7yk9W+rbXWcZoESYlEOmE/hu4Kz7STety15BIXqTsLb
9hKwDi1KQsKy3Fhj2hRijjnf8s2Iy/5X1KGUCYu42kMWEBIciChbGPbjBPv+FNWx
ssNQXiJaAdEl1hpslE4i8CB9yqgnG5HY7XKZlEU5bo3U0HzqfCsQR63Sw5mjxeZY
HWb5WUnC2XxwdTu55bukUntlJeQog3jX6MrRTsZwnCLfcX0ebhLqYfJHet45T1R0
0EdPgdN7ymnJ5E3iCu0mbdTJA/GRJJ9cjOwaPKdbcoFwN49xf5kHIeA4rKd7Cvov
lBZibiN33KlsumgF+RqdU8Fp5O6KmuJkrW6WBZJGSUdFTCo41gh2L1X/z9a1MeeY
eFZTwmLrNWNz9aPm1wJ6Y8Tu9VCcwd2BVPxW/vDAmupXTPFjMz5NS+PtYaKNBT7w
xN54K62GTO23XrVnHL8tKmK63AwlZ+UUfSL6gTCYMSbCEQP2hZBCMWr7onzvYrsQ
sEcwwt1/YoXiLw+rUrGrv8rs6ODdwySxHmJ0dXi6P8lPq/nmukfgsVz5axehkmOF
M9FIlSyuf8Le97HBS2f0BPKEJXq9971YUKWRZJJhpnBav/GrgQGwM2KUMxTjk8zL
yJStfJ2D2xkREtf/LGH+JVNLRxF/FTeacdq7K3F8HtsZMF9TNwDjMbXotn/nfKOa
UvrF13GjMaGgBXxm6iq27TiQ3e0aNmSyvx7LrvPQiLURxQarCG19aR1K8wHhy4Iv
u5FD9/EEaEF/vPnepFYYrNrHnELR9UykRD7ajv4cuY/KgzOyZDefiefgCmwbaFLl
WiZ+J7od6q6IIxcLtTn2KMi1p6MJLvF9QBrCcBU027bdExzlkBXOwwP3xEgPAM2d
Ph39HuNoPWD7eNPAZyLw25IA/llwNVElD9KF6xLTiSNuQE/9w9mwIoBiiIeRoH5Z
wtck7Q/HTvxc0nbE+m6gbpFK9E8wnf0riO2KaQVc8eGzIgMLOOqt1BYcEmG0YLZ5
H384IgM1mHw+NMx63oiegZpbEzBiTMZ/70J+UUvfw14XHCz64O52CY5sSQUXdGbm
7533wVcNg9sbfFAkN0eACNSD+rB7zId14nv24jWujTQq0HHZEBhx90bTiaS0t2po
11KvsglOJXTtVntlmodsLptU2zWdRAVlK0OJRWhSE0NtWe3WhsIUd2EIf7RZtMfo
sdysBdqrezAB2QU3VwYrQ5tVempBeCCw+Io7MLIWz4JRQI0/jX2ZqPVqqANfAAS7
SkUXsPRitFqIGuYg3nEFgvMUgLq1rrG67STLoy4pcrnS2nFXwPEIRoBMDuA0LY4U
Ghlwtlq7SSPND0YUeaP/1Cx8/Y2lgSzNZNtPzp/Wg7tH99Re+9xkugLoqNDjvWZf
JLVGIman/zyOSwjBPM02NIOdBmv2SjOm92K2XaYDNJ/+9wgYHS7gPfBM0pGgJfcE
AuzrhV7JSArU0Wk3ItSCYMlRpuBScKGZcEXaNfm+zuVqG05FTfdfClTFhE7q0Mld
7eYjFvQDxP+ne7wchEuOSj4Xaahq+v7tE2gTH7n5UG6tYg52rA9aP4GAw5eUy9P6
c1sZSjzlTDl4AU1OgWCsxmloaGlArxbVyAucGW1wt+5rZ4QRGiFTIIns7g1VOT0T
F53nlCaNDf9UxeCJsSNmS5BlyEUMjLQ+HI2AuVfQHYCrwhNh4HgOKLuESPQEBpps
lzXVRK1vClmxTdd6xJ2Ak+wQ0kYyYsVEZ3MQmbN9V4Nz/mJC0cxPb8vUmkZ/d0C7
GqUvIZGdM837meSP+AzUF37XUHwNM0axYgDQYYHRezp2rt0eyWpys46FcQI97qEJ
zlq2NwOvR8L40HYFu++2x1qbVSU5moWa4QLv/k+hUAWNLOPlSpe1b8edXQk776SI
rkpDUw1IobFDr7tG79AzsMB0YADOrBsVeDETBGOyeICadskXLN0oEWjwGUdzvvhg
nWlV1TlmdTSBRKXMmwdk2KMk9sKT1WuaID0oNZ3TyZQaJTk6bCUadgafJgRhesUR
iov86WEgicvpYiMUgduq1zUjGdH3Jf/CRttjU5OP0l7/5JMXn6DRfcr9xcgHyvzo
GKjXV1IzRVz2xETCDSiS0Hrw9HTkzpP6BiDUH/LVWuRayqeP6E7YjXa/RiQbqB1v
cd3dXSFv5UGMTFhvx6TfXcOwfjBa/sf7lPvKt2kT3yS9ci18kFABFZh09X6IfRQC
kkYvAhbDScvevhF8Lu/zj+IbnBSYWU13gLrF19xdgKPmKa+vZRV/YeJdGhWthNLh
DhsM379750g3AYnK2ENSK+y2E63CUXoTmUxDbEUIfQgJlgosI7b+o7zIltZtw4oJ
L9LYZWk6vEJ4dOZkKSLJaRGZwHMaXB+k/E44lOcIkPkkWkzKwqWkhbDXkT3ME2H7
+D06R4tnXQZP03v391UvwV9nab/q2qhx58nTg/dw5OWbQMhw6bsBU5ydwqsl0mKn
AKjCzSRJFQPaL7fLqlOdhGdNj0nf536nE/3qw3moAHtAabnoqdRkvLVfXJw20lOu
rao52a4RWSA9CVZA8zdImGjXnZDvyJgtwfVPPLYfSkzsoQ2x2tQ0H27tce26lGC6
onxs1Lx+QdxzGPYsRptgBtzyUMLqHRV/SHfltFl4BVNZBw7G21huk2o6Um5PeqT4
3PXmIiVd/mzAOkwg+q5AQEHiERpnX7UXvbZXU7Xkb1qRmtvsbIUYEXnN5A5uwgYP
rogtVyvR3eVnia56I/CUUzkddvRIymFgtjULjCtkCw05EX31wRfIvyO49jl9F4k2
Q484jE6exif7ZFO24G/VXzK39xKLCvy85xw8IqkACV8GONMEEDUVFstxZaL0Gk6n
4YxFke3DvGkmLem+rLfLMDdF7R+z0J2ndRCUEBSjv1XGp9T1j2oY2t2VHxpnQBni
NovpJwf1gCk0JDjYL+IhDk3ePP84IaC7XSP+CvU3cy3/Qr5d82vr84OZoCaivkiA
d6vb6tn/3dp2kyUvhMkmdoKUMVuRB/metHK1qdSoGtqjEyOKIESD0hjK0KftH8Og
b39d12sYwKVbOYeR9M4QJXpkKTw3bx/Oyr6TAzBnsSf5TWtF+WSfhtIun3CwTTKs
OVsoqWcyizorm2UzNY0jCQHL4TcPdyq5iT1IMkGrGsuRYM1B0YEQnBYEvI901cmv
hl5nEA2U09J8yVozhYb8BPbwWU5ZgMHOEaP9Uzf7stWkFo0/6U7x94g0FlEddGjO
xybjNdkQIGcrMjRvf+36/Uziq9Ndk7CWNQC1PJT3HithcqzAFtnw1uFnB0kYZ/h8
NGQ3gbH9vtwII16kCtdTG6yobnVWsCRxKjZdeobzWt+1WCtg8lfXdny/6kdtHoci
I+nR1fyYUtavnN7rzXAJv6EFEn4riKcsHSjAz0veHJyMOHR4hHIikh4iMCT2qSOq
dftU/977V2dxYrHn/9ewRi/2zfV24WYfFx4UwiiD0zuduX7jjj6zGjJzHIRc8DOk
mh0YrvZYBG7gpv/SCbZA3rD53qmsdGZHtiD+EPMqGITc+VbvgIH8B2upp6uR0go/
YR6rYQBtcibLdSaxAE+s1XHq7QIMibImP5sQb3Be0c3pyntmLWskDr4qZho2m8de
L4SovZbjFMjXJSgUkwd2OZf+SgYQLwIpHZzRxMUh+vsTURnfFJgJWf3tCUl/CS/Q
zZkwNHYI6aysXrRzhW1hfZfMm7wuEyk1amj2kurSCpIAoOEcs/gvWUc5dKu1xo8+
CCtRU+ialDUuQgHGZyxCM2c0MqjIVonGq+29v0IKD6VGXQlQbPI2geExeaOc7jhP
ylpgeqvzjionHTXw9AKlobSfp9CvTfwlqH8ylsq9PE9wlHevPLU4NGHTxeLbJvZ8
EJJF5wE27FAqHFoq3uxsFSQO3F4XpfLyXAJD1CoxLe/jDME1l02m1qhlK2IcTBsM
1F6zzwtqwpKCL4CSDKwz+1zeVYWjBrbe7aHYYoc2QLRV652/PhOS1/wcfNW5xCVw
QNrArQqQdxVVKhgLZFrT6aSp7V2ACOc+rOPY4e4mo/R1zco0G0Z1DoBr6wJNHwBt
0uiNwBaNr0H4okvRXKY/7b6qrgAMBLO6FcegJdveLflVOmPg4hDJMaRJXTo2lM+u
r5HZc533edDnismSM4IwkHcTuV/N9vRVLZYgEh2BlHREO6YfjUGEtNk9i76i+Awz
8CASJPdeiWc4mCa/8W7JzpMCP+xLXKQ9NLqIuYRbuYzFqvFxBdGhJhV9tTcdMhks
7Ugafu6fYEC6XtJA25a0E+xxPsm4lScO20oAsYH2xqOPjSBrkWD4I+IsQfGmrnkm
Dneprqft/Z3XFSapUUYn5bPv4nb/pPnFgUgIEgLdn2GKAzBzbEZuI3BbAncjnK1V
0lwGedtMybYDt08ZuqyaffXm9X/wDNQFyC4xOuzgGQaHKp6gDTqyX2zG/QpTjhsF
xQn8pLa9mylToBozOUiV52ETp6nnieQIFO9bq8973Jq4y/sZqwXYVl5KZ5bXdNeZ
WXlv20lXqwlE6LU8IIJFswdfBWLj6jarqcEEKZaFtG3Nw72z+rxdz+76OFvWK23G
B37He9ELmJDajP+lM7Qndsy9WhCTcfFUDuGw4FNU0zQVMJXeOcGY+pGxtflhUU1Y
kRezv9IRVH+d8zK4/OL3lDsm6sixYmceRhcVfIuhAbTEVTFjwoDSv88RwsDElHa8
Fz3ClDcr+6P8OyxIQj2a6/jfSDe4BR57Ezxya8KL2tStOg6HHEMXPQdySo8hR29K
/L47oJJ6qwJXcDJArwKWYkjW4lCDvRmgvqPRzvpyS3162sEu6q5EZeV4rWJCw2xh
pItoLLM0I55FUFQQO+3TBt7SBDGN3wZHJoT0VwT9j/EbM+e89GRntf9e2pa8wpyd
/eB/KXZ+WzkdGsGUyxtR7+wNgLh8sqVftuY0wXAbEyHPrcXkfU+IXD0pvw1FrXxy
+uJr6yXnWJXQlxoykNQba0gbMH7o2ojfNOLcpqKUDXVNp3oarM5I1hKxzHq0897i
cYkdA6Ze4A3DqD+HKNcsLMDsHCcJzM3emwiURdrK1TU+HLW5wnEFqBqsUgLx1eOn
PyXZTPet5TxEEpeNgHPOSxiCPEP+N2VGrkSAghcqAEqR4GY2Epc1cgQiaHwUGGD7
cb3pYtbOq2jcPhADIoblN2+e3IyIETmQHWDYo6Q+WzYqyIFXI16VHeWS/cvnkC9s
TY7/Gj7/AXQ1bbi4KFuulJK+tn9JAetdE4uh/UcsulXOICwWOr87cSGou3mUmYmV
WzVq3MtIScwEul9PI7Vr/Z297XZ7nGkgOLNk375u+8ENeJQ6RG3Fi904QlF0IcO/
umOp9UdxPwZiGW83erst9i2RS4vLMezTUgUJF+3kpLWGE9y/dFTEEVLTmXop3YdA
uILnMAHyoL2V7fnDvyOHUBPJvQGb4GpoxuszV+QLy6B1O0728glHKVPVnZSXwFRB
EoFK4FYnYosXPl49fOdTK11SUVMV6K6pc9Y8hNPftz3+0f7JbafgvHrEPVDJdgCp
r6Ff2U+DhdJbzzfZkkdSIw2lgkS/YmtR7R7oVdyFcRIyTcjHOP+SDQ+4EaijEaZ/
R1fzRzjm3BDgPYLigilqNqDEDs/PIYmi9WdzzwD3JkeThRRYSe+q9H6kbHGv82EU
q6y8WOfDSjNxEFwiaajX1wotnOc68vmRQ35kwlrS80uAkExag70mqP2UHPjh4Uj4
6JWgQNYuBU5zCmHvfs2w6skNmF2SkJhyyQuVqWgYBjYM2jRptm+cSi7Xq6h/dgmF
HmRk70gXG1S6GU0QaCynNUc/D6KrbsNTzmR29e2GplUQym1hFuGll21cZnfDIjGZ
0Uoli9EDG+i3gS+4hLXpBd/Je9zg/Sa3IetruODd547LLGgmco+wOGTyHS+HyxRF
T73kF7l6qfPvuzlmaqF7L5+VG98Y93nH7Dk/WEgaLCzxGwbYWRPdRkMGI9pSYrO+
oEYipT/GelIC6RPgUbaXxR0cbEkMqrJDUOs3Rpz+xT2x8LIdmqNhXV8XuOx8Hccu
B6OWGK3zkHNizfSMyQGzqnyLMtBRcUHMlNAS8qMMaDf9qkQdOKQRdLWcvdXKiQhq
8uqAed6K8GPmMBU5Tqh7ibA53VQeDig0B3thu+u4B9tBIEVw8DqKc6mrwEqAuOho
ayIOfqPAYcaiVpd0TWTJbeaRVBdC+hxYY6lQkZxoQnK1W6xMWIdd4FIfgbIuD8XB
t3p1U3r2PHJMHDxVOyvp0XqXAmUD0mtzSeXTdfEfRR+z1Gut2nQcqY8hJOb+y2oq
3RRDx2ECn/ImLlGSreq/5t2+G84/VgER2oO0R1DOV8bIzbfinWF2+Vg5GVt42nw8
Gd56O9TkQR/q1lrBWGorxGfEnrrDvuv93fduF8eDk4DSLe3wm552zoH6nr5uImP4
NfK+LqLPFo8M2FhduBVUJRetbSfEpltT1hTfbf1kE9236XwrZeciWChUr7x59SOk
seF5qUs5+Iif8U/KZGv0qcbm+03lLG1BB+qvO1CoMQKSZi3lnPPAeCcRKJKFKVnj
lKfmNBtAw9/yq83Sn8ryc4Q9ZFWNnp4I2vypxWt24EWJb0CYrKVWUBEl6wUMGiYI
qvRjiAUD1U0yvB9P5DNzDCUHiGjSP7/cOHuiko/cLl4gbdAhVqMNYk4xZUynTmw0
+Uyy0qE5NiNeg8kInVLumgKWbjq2w0Bfy67ld0ehlKHNYVBd9S70zXuTUwrZeB8O
JnJAeirBZKHqblkanzS3Cj2rfJkxEAcIxq+QAznNW1KWNhh6V1HshtHb0Kc3y56V
3r1o75hABSjd3QSL+7iStwfFtDj5adErMH0EAHE6dyJaiz5FpOdUd+Jc1nvEEphI
LbAKVFE4tnX3uhdEafijtKL38N4JM2uNvf+zg8EL7Bxe5mKI5lTC9id56DEuElcA
frxNFTprr5DvXs6uFilDTL9ctwFVOU1XLu73grAEIyGkVdU8aEKjHSt052+cyBj+
n+XKBuzPlLDO2tNWzJy62rw+Hk/0mcaWwHnEHq+RWMy5oZJ5mP4yhKcDeRr+TxHC
wwb1S5i2ZIX2o3BC/xUvOYjccKnqOX/7e4Zq0e5E+DxEml71asVqzIocED1uhMGi
VairIKx/Aj2LPaCUPdCviTNPLzRd06do4HdKJH2GyMmosoxRINjeQVYIsm5chzGA
yEknCoGk7cO5Y8pmpa+FZScoH5KqXCrNERFdYEEKnSzz270bSPGn8h0zpuqceD6b
sULMjH1T3t6audhGfVU7gfW4qbIE549hWVLBsun3rviQiqW2P4W/iU11v1I5YGGd
Qh/ZCZV3WSD/C6PouX81VmZQ72VNIkazeaqEl/FZT2xwo7C0CHH+Apr6pnyfav5T
L4xPMiWacBYWfEKxHgMHvStjQmNPmux9ViAQvDDZAgQ4XrM5yq4xG5Z3IUqaXANb
w5uSw/1dw2ubvH794THz4V4rs/uFRzWzKbV0vAOaWmA6deF7iIyJL6HIvWQPFj1z
Lkw6rd1dZxe8ROHb4vDHMiw4PirkMsamBdR26zYHn8SU65YhLlp5CAt9Ka4AjCIH
CIh0GJcWrm8ROlsZenBE+1wnDYAUcekSwzxan+BzHH+eddonUqkGWlBxVEtL8Qb5
Q9Yk0V5aMi/H6ml9xtVRO1vnzCBgd5Xlrzhe0Afswem84hIrx5vedegaQ4LS93K/
TA5po08B7mAdXtrl8czJRZrHhDkzYsH3rWSXAmj3lUJU6Pys4fyVs4jDrRdH4Bii
YwdP8VtLHDRp0a8IiBnfpagflL8YIb5l9G8MEWagGj1a9HYYDN+3o8FWDBfNHvYl
CgtuPgJItQwZUKKmDCBdXPUaLqQc5S9ItfCUgA2xC5CWEgopzxQETKkTO6z8cOlP
wwu5sLouNkbcX2c7z6Nt8n1DRSX3JaQLwypag6sVIQuvOqqfoMZ9bxRkBcmYPOcU
+h60xMTM7kAEEoWk6fYZBzp6OlUCqcbD/6o0R5e+hbOJeF1aD5JaXNklZPNz2xBz
zx5nKcGQI4/h7asPJXjgqrG9ljCdrYLsLq47VTQ4wISSgZqblbO73KE9UltZss1J
UfNV+xuvutpI1/Jnm2pXCSO/vEurVDtC9KzswMjV7q41RLgE07ae+kiqeveRxrsL
qphm2TPrMyEfX3gy/4KNMYfqSN81dQUpiqCf7Gdm4keRPL+kgmFHI1phZ8/q9eU3
p+AcimM9WVy7/WXnlODd8pdXW1HuCARImaJnUDgTZrH/CVQC2b2zk0nAR6uiibYD
XME0WE+ycpGz7ulhclhUhBeJwd4LeA15Iua8UazrztOGqWi2tCT5ANinqnOgRgVc
0hBkKcaQZ+fABAH6Xc+wdLvZD2ldsub7eGa0OBmXzM8Dd3swFFEvIwbt1OlgPw/w
iAj/xKn3XaYO+MyIJpbAQzhGvOsiO7WZJ5jG/Cv/vCPUhMgU1W6+q9SRQrYMcxdQ
lFAhaX42MGDkUNfn7qo+1W2iQ94BgkwXz5AxhnAVaKRu1XSQG7TbYbS3yQqMQn0s
6kPsCRWB/LbO9/LKjwu4DIlTcvWx5DVhhBLr/wYdgkUr9lrRm4bYnCLL+bxC1Oi6
JoR4hE5ddDcUk5tTtaM+bI0GbxUc+KEkV6c8kdhmrQw6LYHcKy5WzhuguzlVUao6
G8QNpmmeTg3SDqqJLHL8tWG5P3Q1WLr9BoWmPOWoTPnViPbyurLkxH45AoBivE0K
kj2reXhds2o4Zx84JRWdQ/k6avIas0kU1wYU3yblA6Rahl4vvfMCVoz2Kjy8Rl3W
0kTxrQm+LUdrchHvJZdyGrw9QTnSbDu2TGigQIOpggtq3LSu13bClu7tXh7JixjU
eV5U1gjP9NugES3pF6anE4CaffnJPrIYd3ae/nXwOfOiiBj2OBVubKl8rcj/yxQA
NgePjAXROwhY6NUUM0HTSJHj5F4AM+PZqJ7eHgYzIOd7xUN3gvrTPGMeR4tU3l9Q
Looz1buUmtN76m2lrawCWMJF8xhngsdpevGYgP9J4lxtp0zgohsvP5eytKaaHSJn
FnudhlFEtZHXpNXO/G3UHbeZBddW/mtOTRDCyvcpWlI6E1h4E4/7zHt7QT5ob+vc
OCE6tbWrszG9a7aBNgewYvdBF2wV689on14gpibvjn5T03UoSJoibXM6KMmiVRxb
fEPXYkZnW6MGualwHJoMRNEzZLVd6/w8xMvxl0a0QApUXT1bW7h8OVXaAp6DK/7S
SkqoH5ljg/ePBL6b8FVTWRqZWb2b+lm6fNqAKRrSHCbZJYrTSQalper7uJZmpUBJ
XrZTWyy4vpSzike9F6O8dLnhPaXyYOqs9petB0kvBlcp3aRwOeAmL4lZU/61nYvU
Z1sjhEeWNrDdLNpKQWo200gcXLYIqig12XDZ35pnhVmw7Jsu4VnldioeFZshmNkV
ykuI/I7IakFgewNZQGruyV8Q3HfD7FRs9Y+zc6jjwfczOPxbYl1pVGLz/0pw8cUG
PAYCNPTMSXzsb6zvpUb/9MertUXAJJ7ihIVkA3k5oINDolXF4KR9hd8OE4byaOTv
h21I90sU78d9Ry4w+j5uYvt+57KQTh579VUduwXOgkTXUzl33Bpf3l5cOPfOyau1
6fsakpZTCO9Q+/AJvhY9TtHoI5SDahy/ecQq1ojQNWnMGZdA6mHJtWAqqnuza9Kq
518d74ok1W96C9NStIee5oN3xOtqMMD/8vhhcY644aaUYuBWsfeAzlp68n3sAHdf
aI70MEr6VVc+Bt0JuKeBz8QrGXVlQ88z9sngYVB4sSFYFalxTEG7duCamGJvBUl6
1cFI/szWf/0g6EgvamMdWBhjtLsCXqHnRdzBqncTrstk6y5KlbSUsuWSiZez4CE/
s6DAM2hmnyiK61/PkA7YnKPf2w80rhymQBQJr3eS7FqsOZaIIzTDn1nOEIqe2y8f
XinHS87J3kL6ahBWGzwa9axVuuTVG8PQoxgDF0HauoYUsRmXHY2adZht1p6JEzVA
WeYMQIifUPVDUhl6VQv2TYEeICYVBtQ8U6cJhRR1/vl7zzYIN9U7bN6XRmp6Xf58
FxlPD63PeQut8YpXDoeZPYOTJzivEBByZgh6q3XWyX1mvl3GqXezQ+NXm3okNGSX
pBidaFqtgWjUZGv9gCQ51a7RY0djYLFqZks9iVU8fVm4OWJgc1rAkGc6RLk00ghJ
XF86fqrY4hQoZcR8gT2wpOJ2wvEyz8ajN5x5Polyw4mm/KOjX43B1kIWQTMR2cZY
DDP4nOucN67YlQHyuUrSIIJjL64qFKw0XLV4KQUqzDsZ+4DYx99qLg7+Al+ADZlv
fRk/r/gYcCRTW4h1OM0phMaKmvzjQEJ7kcBxjbhdkOvlyVHNJcGOiMjEG7g/OzdU
rZhOt31mHkrvZYtafNhWt6dYgoOYQHNZy9ce2EarYRrLH3hsaSu1gyt5CXv7WYHF
XjcgWyC0mLvthQd9Py0RqRGEs/Jr/j/V//WAhGYkBD+WJVqSYaz0Btki5cxFaPrr
c2Q4YxF1Pz3OHf8HMdYQkZCiDaUicHIaHDGzCXlMGnHNc+tIPZVo9rjkC8nf0YEb
TuwWBb76dQkLDU6GzHXtVlZFDGu58ns94bTN65ncIaM1FBOvQE2Q+I0Flf+e35Eb
tpM2XmqjrBD7ZI88lhWx3TEjgqy07OmV0+ox2Kq0j+lAcgpYYMq41nx7zQ4OfV0s
dnPUF7+9ZFAVUespRGIZV1Il+ZuIW8Jrm6X4wkMmMgn9qPJl0L45DBq55YgIJk6s
R1SLVFgMZwxu856QFRaJ2xYEcav9xb0kgT/wcZMf1yR1vclcdGey02AmPriea7BI
lrRXW7GwxQfyQaWCqtFE8MWmTKP/yM7cFpxgQNtWHgj6WmKjiRC0+p+GUHRl/ArG
GZDCBgUJ4adR1cD7WnTDmWAbf0Rx+KGhP0u6G7CJZAamELHqrxDKECyDyhsSizRR
CgF9NsNiobM7VFS0vbRzNMuD5SYHLpgXGdi2z8AroCMmllqVJUKUeixt2aAsBsWu
gXPnHLN77AEU98YSMUT7Z6dp+BC4QVCVsTyDkL9orl+Dom4xpJttqUGDPe+um7DJ
Zjp7ZGPT/GKGZqCUpa/OMSaCfFv4pW2Zzwe/HbZCR/IJPILfdgM1iQtOz9mVY9iE
2ZTUpOo+j6UFNAYsBkpzcOFJusIVJlxZHZ5Rwp/z6kPxn7FZBZ9RW2Cb2lQiJ59U
THVtYjlIUQ7bfI0gE/KrWb5F0YNR6BuaZQdCBtqHIwJCXbw5zbxOdPO/skzQt8hO
O69Bs8ZIbIi8bkWCMcttxNtHYyEHBmqgmmPQIW7Z/EFCYWFWTAXizzARG6QRqIxp
ALuB563pnLLXkk0T6DSgWEUHl9WyZXfjbEV6s+Hgb7VXmqmUSZK5uGd9qhifs3Xm
Awgfml2+Ah9TfVBTfnm+UaFyimuvcIcLIkGNDm1/UOiJJjhw2N2UTwjhAnhVgngf
3/gOw/5MAKq4tU3NuOmy49bc43TMyBFysAysit7ApUv1Bud/jLQ6OqoNdeb200Ys
4SjmvxXaUyVuWuwbKC34cPZBmluwFawZ29J7/VxvoqppgUNpYXhfe3IHViTec16A
Ds/wZsJdbxY0pJc1zE1lMZM5tz6TPDotNLwZKLaGNX2shTTbCFvB3JOehq7O4YFL
HZxuJ1wDGLVhBG4QZ+3Gkjq+7lIUfoWYwqgSIvfrL1ADlxD2ubtx4WSWY+QhIN9p
SxASU8Kg2PoRy+X/K8s+x4ebjovgt+8yH5Kznuu9IZ5Oi9nzpnMW+P7QY0co2LTy
qXuVwxbd/rocc1MGWKhNRyykAf8vricO4JTSBeUEGbDGQfpjIa6CQDvargqF2hvx
DLcncvit3zOvlIT+kPmfpiFBa+MIHpDQyFwJUZQ7rWUtf6AxocPvwcwSZ000XF3q
OY+jzTwm9dx88arvqqXI9eFGZ2ZI/DTY3926QzkBO26pGg90F8nr2itUJuld0leP
G2EDI6kHIGS9eTLjoSrNwjK9JyOSIwat4kj316MxgCITLlsWjyqkietDY81cf9M+
vG2CEaTY+u9TaV4Ot1/3sx1pwiDl8npraIoEydp3x3EDSQFbPt/kqiNtTonvk9bR
/0nAwNzJh9eLjEQtonJpY0fw5xI4AU/Cl8jQ67Rm7tsdqayjPuPE0NDJjm9n1zAR
VYUUoFP17gTrQNibhBB1fZqjS47UINem70NWhCpKEbqeo/FDcGBfzhVCyJyDnf06
IeN52WStkpXu9RZaMrECxdDPYzNDP8Dcc2YwBu/1bV5cl39RWYXsfz8Txa/1/phO
iRHK4ElcQYbplN+bDxwP4hsNsTzE4zTVPCbbtDfEodMIVavhmtuwZFp4FL+SurOg
8WbfxXFwNrmqYL/KgKH9Fjlp35qZGgZ6IgvdcOFp3CSVz6q9x5m3a9L+vGCCFt1t
/IYL4AUjieP8qW5s/EMBxL2RciiXiy5BZQJYEnj0M6OWYahiMNq6SieUPavvI8bF
ipinDrsY51IyNgX8pmKoSV31xhqgEFxUa1Z8Kmb3mG+e1LYxMXifnACwOofQqYDW
0vz4Yp7bSxHf/w2ItsZlIdJ2yPCHCyhQPlUtZRWLGRkjyYL47n2BFG9j+bgTZ/mR
SCJLBPGFpNV2fqvy5JokSz6re47MitylCyULgvul1fruGS/cZbyZUnBlGgscwD99
gZThW8FCw57LLmK2UB4oFk4ldnXp4QsE0viCqZ8NawhfdbCb0fhf+l6nBfpuYADS
p5scvIqRgWOT8D0doa3ijbvOlwEltQS6pN+HbD7EcDRtUcWnns/tHju1H3A5UxD5
sfz7+f/2xX2IgkdDUHQ7o4wowYQwix4rFGmWSSuljeT9TnMYIPV/VnbtHGMzZLjx
6GX7IQ/npmw4g73cp/jGSNC8lgnCv6+aZmmdkIaJLt10vTK1eHWZrEksS+2S5ig2
AsBYNt/1tJg+28W6mK29S7jfPPhClqnUAsgZtUTdtjQJiastRFNgg1ZQxgZbjKPF
Pw27Ub2VnMEgLeVoP/UBk0HC6o4GMxG+yqBhhoVFunWwL/iE/aDWtdKB4gEqpsJo
uAsTYPr27WLm7u1NRrPsc1g4wubow4S7yhZOSahS8qza3eGwI0vxSWLJQJcMf3IX
/Wtv9Y2cHkVoTx/1DfSECiicXfdGOc0orSWeA2JdxjHQ1gbf7JeoXJmNpVvjQDZY
LEwm/KpOkNlhQ4qbro00lpNEsrdM/7HgFvgexqdMYX1UACyk1XoWLrizLyCi9Rgb
4htwUlrh3Zhno2MhFPmsilgjo0gIVVzwKbHT2gyn3kce5hzlDp1oS4RjEf2yVapN
Ys6g3D7p9p2kR1Fi27pQTGYlqTcezsOa7ZUwotDp6ak5H84a5c3T+82/D+QRiVjk
ObKgnkmRWuDawTL1USvQprZGLUOx4dJfFEHpeBV6SQHkT/7rFmitRYolVDavmQV7
sOwCEa3A9YNixibTihybgSUXIku/fHhuhvcFEb8WkQrlFTlctTbPc1bgMkuuPzLm
SPVV13vPHQ6p0AssCwrtYGFAqJNUBEiJD2Y2+8PPcA4iomFbVZKeaiToU/qnHEbg
Ceyu/XtDxohpaEKnKxp5cHOApuMHqk+6fQ7AaV2ydHW2LhU1/Yii8mkFnocjaJ+E
1Z9HOBUqXwHKT5TmbZbnfewaPlmb0D04Y5r9NICQ/pb+gKPiOb4bXg58Z7J0Eco4
dnfFNAeLnRSLPS31JZ44Vuc0Qak9cODgaP2dzoTb/aDN/tdjUYBBbmWZnyiEYphH
zVPg6asY1h1O9wGZKx8LKnjiER8DmFk7d4HA188n9C9uLK4PaNTl+XZcIo0Yy+OP
NFH4V/NMSiAqT5GYTrWLzkLwZlpfBS0tTB254xUiml6s3EOuELXQmeIfBLLDnmCE
0sUKpIB1NxMO4IClkX9LDayWc4xpDL/VcIkX5O18fSDHBcZ9X7MHG/50r7BgazPJ
0MJIB7+iAOOhhFzmOwDKPYP/0BZEjsrBIujLCfzb0lhJgepBEJ+9bB7mWkBvmUE/
G7sgLJ4K7LHq26b5Hua0qvvS5RHtjRWGFeB9rwkwYHdOMEFWQaRJZKKQ5LAYFVin
DbTlhRxCGRvksMHiXdRFKO2oxEFQQeGQemXZTdVna6ku3HJB/aGdXoKmedRYmb0A
8ISuN27VmkIxeUxufVhdPypaCMgX+Rz17ZhBXkn4qWmXbbcOtCLnKOIU7uD3rxzd
IqzuTnVUOnkolgHyTPpfthlbcxX+4EQmugtctkaSBjFUQbYl3o/zdgsFFD1DMDGB
gP+Ao87kzsY/wx83YFniNkJHvyvNVUXFZlc27mt98JSAlhaYV624ISHYlfPpiBEe
PVPQcALlYg4WMyPbApqrt1GPR8Ohq3BdybuvMPOih+RCOR8NZMGEikW0XuQ11COG
qZiEHt5RnOf7pawui9qXW2iwHpDHhZpqGsgalFja4RBgADtCXRW0K5kVP/ldS7Hg
x67eQXUXGsJKjvLxovPiSJB3gY/nnvYWBs1pKzAa2aLStXB0vHShhlKfVLu9HCcX
qlE31WHFuhw0hoM6MSxlWLeGyU7zFcqzQ0AIfDQ0lVLWIOFWE0qIMm+loOa59OGC
OEAi8b7JI/33tndvVP6y8BU/9Skq62Zo/Ow6/gJw7syaoPKprVBE3Z2iyMEexUJc
qy/cHEsinjeGauR9qLRvrcQGnxQYe/lNLXENzf9EPXrr2Pstp/mrK2rNnLHXN1I4
0px5cAAQTKbmGIv2tRnDv5LoPfwTXp8nim+0E0Wc8i7xTIgGtiPVZ94M/GxAFn7k
f1i/XiBcya/RgP9sb9cD4tm8WCr2dZKaodkawbYKmyARfvuiDQY+FXmpeTWn1Gip
JdY1gy1RCB7sowCeDLJEYkjbTxjFPzQHjO6uN4g2VDIjDPeFmAZ5z5I0J+2Uba+u
Oor5A7S+Rqk+H0QgdcEfr9L6JoIxIpGib5OeyCVK6zUfB6GAbIEmHtxHpA3EMUYE
0tBhP5sB9jMjiuzKNBTi6RktpRZ0qpMZD3HXvaAlWMlmMDm45cHj6rhxq7sh0GJP
XaNpgwE/q6aLXD3HyJ7jB9SlkVM3bAJIwJOU3i2HYwwrOVhceAV8GGPKDvMu4iBF
cZhUXaJs+GREXnHpc2ZrOL0Cr1sQmnr64shBq5FqjWCphZywIotIpN+GviF9nVfu
KpabTgSfFlIbKyUByhnLunqXrkZLRklKzRsiGnnwE6eIP4HeUx3zxVAxXj0IAiYc
V76gJGzuLI6RnHXFkdleeIqFq1u/URK9TZ5w5hkbpPnyajk5Sa5ZidcQeLfyRsWK
Ds6TUnCitLEQzj7XTEIr65hhFFr6XUV58FTYz8g466Z19GRopHMjRK99maEIyBi0
I4dR4DCt8Z8/UFsrPnBLpGqg3xJ8okyAvPxGiCdFXHFe2m9B3bG87sDiIN5+9Axt
/HXBUnFfnrz5SrkkOg9e2u37VefZ5IiSii5Tl9vJzHNlDfXFxQjIY1SHyJjQDYxH
rr02tHfDhQ7G5IbTU7cTEB0lAEexhfhPZQ2m0XPoIiorTgkaTTkPDpLm/GUJgvbw
7+KYXxOoL+1uGOCs3IiuF8yOUWToavj+TQ54Wa8A53jPk95glP1vSd3NF3dlAJnA
CBt2tXhzzREDuCeKDCFX+Tsns8xD0wLhYIgy6kc9Q41UXzJ+6p2gY8Fwi6HDBar6
iihQ7nDHaBZiwk3JFL73oWZu1teLdnOeVRm41G/3qRijtxN/0THkh0A/779AHCGg
+DEQD+e0xEvfXiIU4sOsvW8hy8yFJjm5p81j2fDkEDq70Am0NYOmO2HnkFTzWYVN
y4GLCOb1kXEBxc5PYGLQCbP39y5bwcEdxYNlzpr2JzAnAbCDlvvb6JT6fVD2vHaJ
OSXmP1nGbmop+LqsK4QKQpSvx0mSa6kpQjWRdFcNVSTVQCz8KBo3kFRU4gdfH0Av
Ud32+tids+pB6z1TB2hCwRXWWq4hh5i8x6qr7l4cQfwYn5GEfvaHJfP4vRvmQcda
uXwfj3s7GSnC9iEvwIFPWmqxNmPxT2x2rpqVbbsOOIMQgQWd5dQMpVCBehOxwWuX
RhEdGBPbLuCweRagAwXybG81/0iqoXteHclmPy8DxIMPkGjaPlUyRf4bpWJ/PehZ
R9epg1ctL9kTMBUN6g1pkvi8oendsT+hn295ZSWdZH/e+WmyXH/ovR3I5xIvHWfg
OY9l777TG1P51UwvdnLT8P09fCiFd9L00ycSAM5G/Q6RhaDR9iM3uYMSOIM3Q4aM
gtYkzR/wn5npn0ZPYejF4Qj94Mp2HuC4pXvbY47K4k1ln/4syEYH8eoELrjXsDUy
VxqOPLAmNfy9Kc9LQ/kiI9LWXv1Ts/AngJlPllSt3oop3DxNxJWwD47ypcoGIcJn
BvKh4qclpluEVtEDN2F0yM2vuT9YR9xcE8HN6LM55FNx5EgHy6SYDajRz1ssDcas
XTEwTs2MgTqSgzCyubZUvoZUgy/0jtiRWb6HpLefR2Kc2lkV64LQ6T45aJmqj6j/
idAo3YkrVpez383iJIQgy9+j6IhScYeQbPRJJ4al4xbJRGCrgIP0IrxEWPncrMG7
lX0YDyf7TWX+ANlGJtV64cYzFln/2F2JoB2Vl80Sm+enZmEiljbBdkJutKUWBHof
j8amRxUG1OhE4fYQkgYRxa+wYNSn6T4GORP9FNBrDrKEWDl4RuedjoLjF+/0iFX3
H1sf6T/IXa9ZxL6ZoHdhvbBor3ygyXxRaZw+bR9dkryDyCE+mvEr2fiK/qlOvsa4
NGMgH2yEClr0owQYSvWAcSaRZJz83eVZRK3sjLMSrFHMn/lwW66iPUoWCTrwnfBF
o9wPR230eSAJmC8ac2NmPx8v7/UWEjhmTCoteO96f/g+Jplfxc99CmVcbdLPZrOe
vm6qpIKCalSkp7+HbuFlcEX9NnYPafndPKpsG+x+jjgxbxHrgcWxg7njeE3d6sHW
qGWwc2ND1d1YHz2PQ11dO2iAWiePVqiHZOQcTNop5xrxVdxuVIPNqxWgQq0VtMqX
jwrh5Q0jPaRSdbcsOYf/DA3z44x0cNI0CVBD7vW9Zo8/GpZ03HF1OOYxnt0iPmiB
mcTaza+u+jYr6j1EtGFt7o31BDmjZNznjJTypu2N+9eWiELaetNOh1rNSHmUUytq
ammbKMiMLgAH60+5zuxxSYAHLj29xonIuFCdiPQkT9Mz+RrUAN5bcugLUJI2zRU+
FmBCcztqFQKjxqWugrSjhigJI43HIYnRdeLXJYzcreqrKHgzDGYqrzoDMi5IrIlM
891dp8sww5k51cWvt2rvmmiLYwEwxXpp0rLA79q2ybbzfopKBCgh0CULGirtqhYm
THCYXK4JPSoalOtfZi4l+Ns9PHP8tV5OBHgVrmmyGJiAaLgj/JlYtZkv6JoQVKC3
SFO8jTRR8v88JzS6K2vh8irKlV8jWbfIzyxP8VLqtN+XixvaeWO4f2z+X6h+jzQ5
BhcN7DZUwdVYT2Si6DN7dEo+VkEvBS0LNSfIR5pX8x6+8+cKfE6YK0/iSwuwPOuP
CJMQ74ysm26GBbKzHgynXZNgWz0zZqATuna+CKOcUZzogVPyhYfcu08vQsH6PYsc
JPgv3RbR0ZZbVxnK+1mq5dhyjWlxB2ADvYvbMQ8ZY+SZEVkjxzsxu3u4acDG5TZ2
jdb3+h21aI6K/feJ/9biCr/1rM9lswJmaEnhkHPAPQ3Zf6dgA2/mCjCUnV0T/NTv
9jpabNbaa3QU8hYqi5n4zPOmAcqdNw4WYFR2E+nh8F/GXdehZ3CkVdzHRMXJADcM
juN7mQDHzWhZrUxthN6w2XPz9uWsGKLy75dfSmahoXJ/ciGBp9tNWZZQx7eYuUwG
jLRVOd+EHjYzk+WJ6JjuDsBg3ErNgA0xPUinCm/uAWszoIZ3XLY+5AAlNr0+DnHn
V5fvMzL082mKwvd2MdRjC1YNW/c9MJabXHJrsmjaE3ui+30mhtfZmw9nANU4wRFd
zHrcuUADPKkGt1BaRB5r8rCnN3jvY3+MvFyT2KCZtogLpErsdLcSg9GzbbKV78yq
FGC4WskCq6aF/hgmy0nFwJ/K9lUVeO+zagQXXvKSQnzkE/0Biwlg62Amv+XHnsWS
L1vrf1hjVB3q4C0eCdZN4+iJ9QNdi21I3yAi+nujGWFVmk58JwYHl8+ffmtEv0sR
4krk53dP8pJUB68Kozx1nEvA2niOfXJXmACJj0qWdTfR3VjZBWjLUpjrnIyAyQqF
QbCBH4dBkoCAKXNSgDo59z0Upd1GpEYUgEOHdc8H0krYWHuQUgvdz24Dj39/R5TC
EKf378Y8i/B/1b5FzgRUJzwLI7kUAZ4S2ZyoURWqhxxUQbk6XxgpRzz3UUavGKcV
U+iTVo8UDovAg7/VQEUDgwoFCWn5IfNy1KcQnDtr06HyJcpW0pc4Y3hr5ft9bKZA
4IzfpCi/gO2nwmThISqSnpeztMo2S2oUlq4j++PS/BnpgvsHG/8ElBixwzYgjKYA
L2q+adwOeqyHK02KYlvqwkbDHatVlxDSM0dAL7g0xWwkSeh2iyqLCg9wKGXLspHk
Surs75g0j+Kwu7Y37nRhHqv1InSY9pE3oT7kwrMjeLYFPUD0/aPEOIWr/6SIPDwC
9sqqhlpt/emnrWaMZATMf1m3m5hC4PB0fiVJgKgJS2FqpQ81bDHjfRSM+uoY8ej+
+OSEd+FBihSws4/6pkAda60KfWGm8FLZDtoTO1230eE2bDIkr+8CJbEeyMFQ865G
elyoGEV2gKMYzbp0ttIS/flRtD1aXm04IPKjHxyMTViblU+zfEjTDYxzUdJPhJmU
ZL8cb836c03Fx6+qR/epRSo/be9UJS9ONxJZSGzNZ1DJ5AaMRGu+6xlfm/xL2uxi
RmPW4rvBwVTEC8YlIulty9Nzurbf28JnmCq0UgLT7PMDqYgvFRjq7fMwvwKenX2V
2kuIbOzfBr5CBdnREmsrqAboIGcAUsvMoj+2UiiPhMF1yidg8T88NeE2QYq4/U/v
U4ev3GjU+PKk6KANpPuZCG9yRueS+FT2BCVhJVMyI0QD5cv4ZBzUJ9T/9ptlZ5ZK
/T7V+C4jdvVNrEXCs3Suhz05DU4MeLgNWEIC3duw2DrI6eUgqUird5H3KkD2Shvr
6aACt0wMjkHBAdRjqmZuO1hQLlA0zJzhukseZD/BJh+6h06ORTFGuzd+Ru5Vni3A
aZO2FhrTeF4Z79OXE8uS15yoSF3yT1hM4p2vq2yPSwLN+Sn5yykAp3u2GzjBV6Bm
fmyvlZ0KWMwJuJ+WKF+XB4CKQGuLgSOPxREzC3ULDl0XwPt8JjxCcnMhQY6hECc/
/WZvUHh0PDxR4e8ZclkSa2RslG6FFZKlAr7ZxdaLXIr0JfrMlu5ndjkltGI8fW33
V30X8PzQwU0wN6jhGxl1x1sPWOcrL8205iF/ZDIbUhxSAQfOMXsO33gjf7AJTMo3
8BFAP/9MmaQSS5hQtbqEkaqyqjOFOwMKismRVEAnxZbg/juvmAnyHMjpC0wHZZxn
ZZ0r7KRia7P9HwGIcm4YIpnwZsjLJTDWzJccTnFud5z/VcOmpW2x/+y3AAkVRLzP
8/ocbpruJHVuWQweYAHGQvwJeIXYNDlHJxLeE347lyuy6CH8pAUi5c2U7DCbSBB1
31MgXRwigql8b0u+FtKL/Q3Vk4nw83Fs6srjXpv0j8fEylEE8hjiCjYIKIBWCcmu
HKip3hm76HZznEg8On0/gziH/tJlzFdRlNonLh92DjuTfz7lk7NCRZvk5cDYGkHk
Rew7KzzgVRRYeqpMJTB/ytntElLGfkq01H17afvylIxb4S82cxvNNZW9y1u6pWUj
IMDj4MilrpPk5b39g3RMX7U2YApbXCRYL8RuQUVotTp3W28OvdeE2XXdUnAJj61W
Rz2Hr7YGXBQ7u5tXKi2aHAAndFmbDp9mBcNXc+NanioJJ//lXHnDXsaKn+XgEUpx
bTOHxUFemIUOzRgIXQcUjmtqSUZZauILlFm3PQK6vD6IcLUM3vasnH2Hzbam6Cm3
tyLyQHWnX5h3j9XELlP+RIFXoGYqXIcSx7SothodkuIY88rcRwZXnJbFZXGC59Pl
m4oduyB+bW41K4CvHfEy8WkZuwgbdscrF8awRf1tldlUvbG9gKsaJM5I4zM1UoKa
+HT9UrFOC0cXExi59o8FiE4zbUSjYXoa7KgnOV9QXwD3Da31XdvOFTl9ZKkpsUMF
YQ6HVa/iIN8f+J3KuHRlNzqyxpAnVO9gERWQgxFz3bAjgHycbRy2rgVctE+EmYDN
SHpW90GzQ0nLh6DaVVw1qo2R3kcR3JGli5Cv3hkr0CYB+oIbIp8xR4+5ME7m4Hta
LhssS0XkDwMgJHqWVSjQbh9iJ12hco2bI7R1dZeZUnSOKx8EEaOpME/xbnQDILwC
evLla/H3OAMymWyL7HX2d8lwvo1s2u5xN1Fe/7fd8HuJjGk2N2h9mSBgY9nELqYP
M2yJg6/twtk+oV/DEOUwhAzQ8MWd01jqfoIkT3ZI0U/m8mF9GED8DxsPjDnEYnBO
NRoFl1gdlBZtGGT+zl4WFu5ipXyfGyjqaoaOzYKb04bnwtk5JBT7tvxvJ2DMDt+9
OUQmfou/05iJ12+0LpCtikfdywF2EjprdEdocnMOMbvszTQ3ea2CBtqax2CGniNW
OYvuNA4H9rrPsd29y62CQ/9JjS3wXiVt6Vmr7Geq4Dw6bn6K0xYVnabk8tax9kj2
v98IiFImXO1awWjV24pid8MaaQNYWYs1FQF4kIJo5BBAB60h5XAIHSHGCwQnQYxC
ugISfXsyrmnz3AqqIVaon0mz/58rgLa1TaFW/fjgsGP8OOZj+kn1WngjHYtkXv8b
rt4zz/xTNY8dvjckTq1q1S4BDMZg/gVyF8rbrg4hXXv3CRnBwZCCSOW5pLxUygKj
NO702l+3f5TMwHHUdqsfu0aVR8cSyjqlq7zNJG/SmCgaiOSjX750LK4pfKmjzMoA
NI5lfFuSAMGScz6bVxA/DrksZBeJzIyMszd7ZQeVJfF8HyGzKKa8xnyrirJw5jR2
KGGUqiicb1mxpOHe1V4H429xqL6H7WjuY/5IFM7y6l754qEoehikWEPq5AGu0D/K
Crpc/tPtWHQqccpilivYmfUGQtHsVZccY+k73LMimmvQAR8Ex6IEe6h/odUywlBQ
zIZKALmb9yHfIiRs7NHEqTpnpHWYkOzSvNpR1X3gxZASwu8sO4wstNjrFizTBkux
o6+edacAL3yeeWCzoOy4LIvdHwK/63xMR1TRtRZ8m6iAHorrEPWTwPGb0mbssQwS
4zvLMrZM9WO9fL/Q0FpfybKjT7ENWmP0cZdaxxOAJJ8GwRlDFMJBnuBdPSA+Lap/
XQtiIOVsniozN7K13KWYSwxb1qu89uQh6j1q9oQf3OzOXRtNkTedVOusAGGJ5uVV
4gJ4+oLx8/eoPHIf/PXuk8kpqxg6rnFYXuYih6x/Xv6nQmCyUK+Sbnt/fvidpMcE
e2yKwPyBOfyConSRaSw4OgZ+6c2aolpTUa74HxtfQVt1Rvsw6GsphxLTgqGKISAg
StNNugy0Qd8+YulxT4E18tkrt+mNDujoCIORXqa1ks70/DMpArRZtGGeujhwcFvi
5RbsPicAeX7Gh8ccaSIqwAE8Cfc//miet88yfKs3H0kRL1zONbMwKzCu5FV1BAtV
tPIOslx8XQ4OWMQN9Ui/mO0ItNjadF3aoiWsPtnsjtV9Jf36A8VyV3n1dt6ai88Z
2F9H5vwtNTGCF60jJZf5IU1gHh3MpHCn46sRkNnWSdKH944VaqYfESbHlm9DGPFb
gi73L2GKytCSadnftJAAz/eoZtRySaHkBrQKszUeGfCJpVMDafNVYpJ6csIiQIAi
CeKaDzg0Bfmzw0hJEPNc0jjLwmwS3XMtP5nsQ8+a4zCsCz1nyP93fHiAcWLtG434
UyCrvMPk01AzptGIpbCa1g83ku5IYdmVIRA8ccnsW/F34QUf4iTgjvZSmsbhLNNP
aixdJUhrwEW8PGOPRyO5zVFMLWcYFzfBIyuifoVnj0JL6Z0x7PK0LE7PLV+Kb4q5
4rlV1W69NZ/UhyUCgbyw6sb63sOESYVAEo7bMQPSYW8UXCLAXBaCdxFYTy08W2vg
JFlYlG3QAX5DUgUbcvbrLUJ4G8oUCuQ6aUoRSp/05WjQq3Jxyx7DBNFz8/4QFjOY
wPTYuuhxOSb2y7ARqgMiQBVCUTeEdNSgSrDheEbvg7d5NuMbGuh8AWE6N+R6Qjcq
iJOPPdbnUdW+iKI7Czyn9CpqCRi5sI8KhusnCJe9BYm0Dd2GuMh6CZd/pAYgYHfg
Mm+6rts6mKBqD77VMCNjxgARIVI19Z7zaw2s9D06nUMrrkq9W2FhrZ4283DYvmIs
3nKkOymeGoj283/4P6nr3hAKnSn6tUpiTgHFbgTLlE9EWX7c1AJjY8xOodLy8wDU
IjH7y2RUdTYguw7PV+wWAtoeJFjarwODW2s5qC4NYWxuXHY6WTyMw67q08XhU1qY
7e3EtcH3MkiIUKa3yLG18WzD/SsRpKCUbMQ8Ag2NefD22O8ZZgqDGi5G/k4+y7pP
axEnZCUwjQrPoYNoFDRNEwlL1wJwGQ1px4v6OYyCrDxTxlfOENFftJx1QrVZ0DZI
9snug9+28dyQleIICyzVbz/DnpQc4r9hjj24l34GsQTbLwk6AFUsV2/+J/fOWJ5h
OtBUYwZsEkZwQaALpVC+URas2+wqEu5sSlLb02jQ9i6YQr9XMJzzGfk38dZrXtcj
Khq4lIYVa/xGtuZI8iX/ZUS06mlmtZeKsFITUZqHQdosHa4XgWD1/K8NHjfFrFXB
x4HswYPS64TLJrlNpUvkt0fjyGcS3qSDoblusx6e8Ec99pihctkc82PuzCmEVXAn
3jiCtgCxgBywN4fbBDUrg0b05rTbykKIRe9KAwuZ78TDR+c++eMgxhpd0zL4Aysq
mH6RCyFn1yg5r6cYfVlRxSPIKA7G7niwEa4VHLH7OEIHDP3SIoVn36nvsaBo0TGx
N3e4S1OZ3vRAAKDqzSnGmFU6iXDeRul26VvF/pYHOpWJYlUv/ciJbnv2qtIUXm3T
n0G+PQTz2ep/XlbTCHvthNDdNksl2vLVWQYWaQUW8gsl8i1FB+V89B0tHUUoJFvm
0HTfdbEEYxryo7fzt94JyreVpskKGa0zsYWQLEXNcSrAPFPzpYkxDTHm0OpvrDUZ
+Rbz9DAqP6QEauDUSx++oPeoDOQI5SRLAZlhWBJdFcog3aiqftCRsuHmT1Blpm+b
YybkJgzL+Tq3a5soh2nOlonN5AWSkZ7T2WV4YQqktuN2LdmlCjO8h6CsY7TuaYAn
hXT1BP9w1Av9E9RJ/d9hlkOe60vvlrZROAwtQVAyLUXmXdEmbL3ljc68Uvv4LtKN
eqym4uAZKd+GpY8EqTTbGv7q/ZD92/VOZp1or55RQZTl+KTmyxMFaJpy4IWHEjAb
fbJAAcRwEoVMRrZYq+beVrBO2WYC1OhCsYnqUGpIinSkiBLZp7x6bega/ewAmOnh
NvlCGLnunVK+7sX2nVYK2BaHjQW9ptdcANjW0fF02KjZOlZXC9doY1MlExldF2HZ
72KJUvgGTuAE7Jyk3cKnIt/Z/ghbz02y9Fsm6E3N/587qsOo3MTOfC+KkDnALwgO
mCmi9G4EGQ5yeRoZ/RQY/21jdIwuCjFez75wklxbJ737CvNfpsBDIrquL4ihLCoT
+NYx/rPD3hze+M0a7TX+q5w/SdGS0TQ/YQJqniLoy+B0JyTp3AJgfnwVZ5mbtnIF
/yjJVu0SA4vninDJg0mkZUk9QtcS3yYp4GtipuM9nDnBP7LtbOu0PWWFsXUGcW/X
RxOUYeOg9+h131cro7hkWfQa0QPuknuqHeoOhGt9y3fOj3Zs9RVk5YaQUJC0LllV
c7S+UC7Ta8ebsXxj8Qf+Sqf8zVz4bYSV1tnQ1Iexajj+nWhNLRWVfOmTuCKCxdU4
mawr+qXbDefKWoNa3nPcbhRt9uCiLIfKKevvx7FYd5heJm6H9OksIHdQHLtrP9Fr
1q1b/3V8a6CiXf5fIaVqfp6J+FWJxOY+0btsfLghv/+ESsbLkGM44UKqknyaNvHY
/W4pQOW7mLngHOp5RABtHTXCQytkJnttiNLgJ74I4ilzxvKiasKiya0zhg9PyLG8
ezY9CtVPfV7xcm2n8CIYZaefJSHd9Mh8K95E5yYsi1pCs3LAlNvVPy0Pa+f8IxyP
TfI6v5hU3buQ8puhL+BPgi2FPEMQzyDZ/y/cc31/9+KLdVn3iFdFuCqj/bzHNwX7
fhu5u4OABMoRsGrh3M8XNENphfUVX6FSnscPaPiLf44cdwV+cRpNvvJdJBXu25OX
sMbm/kysb7Td/dlh1Z0vbbJLiVYsgx1LwWyeVn8aV3JwjdCwfw0uNvLD0rd+C/0e
hNggdZqyX5Ymxh/9QlS9ATRP8yvl6OT7tzK7KTd7enqVU1K+g8udUI6To0tGLbjd
3n3cErScZU3hOaNAuhnZIrkllmC/2n+KwyCLBOIUv/aJ6WXcu7cBObvD58G3O5Fw
fcNTbkAkBCymgf1Cpgz1w+NiiRZe8uuZCuIIukCK3bpr+qrPkzmTNJwBsX84Ekwa
URFn2fCfxsjBDAxGXPn8dmwZSQT5cMOCRfNxWLmT/dGFzk1RA0lap2Uh7IVL6VEI
xs1xifaq6zmX5j/w4bEzmwYqfhBLQbqcTp7gHW5WbP1KF8qT3m2BtZizU+Uk1+zr
f1kLGr8+h4flPZEVi/hHdH1+90ytj3C7ShnhA7DEOX3WFO3/y2e5BICufAfb0mqk
TVOPH32B31+kLCB+yMZL2FFvJNVVPMZ3KVHV7i7WgNQE4f73edtly77R13dZUNfE
cpqRNr9txzRObl2dgyE6/6lkauouia9+oS8vJYP8wEC/B3j5QHRO0ALs2rxdKaBq
4VaNNbgJJJexoa9wv9wfQV3KjKzF+49oAtReCQE97Rdp/CnxsffOdGuY41pRJHlB
Dwo+1TiAwjVY9aW7hivrh5JnfnVxBJtTZW+Q8UZrEKLdF4I9ZsljPFu0zVg3MXQJ
CjqtFxn63NX9iV8CiNTuhMr2rrNEViFBgLykKqintUbs05xOsfLPp9e0T5UlT24v
/8b3XrOLNmQxlWRNofc+zQ+JpttQEzEqQDDAr0k/sR7sNhtdDhn6Utpb0GDbPYu2
yX3bn/oF/7odCS5bqTkTOPRajmNp42LR1DTojF5EVvfQjkijwrgNBvLU4b5Hi6kb
c6c1BwrI0zAvvUG6f1rFUyRiwGVx/W7YzijNGR80T31tTvx21Ht0ivgZP7m9HsVE
m8UJn2nJVVVe/YaA1ASBWLjFLIOx8G1nvfz0LQ+wcro3NaOajhr6F16zSNGDgKyC
jAuF0Up5+BGb5abDg/7OTdGSJWX5jZhNb8EYTxaDhAx9nWN3z9J4gBJ4m8bCKpsk
IY8OGN8dUxOFpUfExAmSxXIcrHyHDPxUzP/XThvLmktSS23gVe030fPo1iVsNqTl
bp7TdC6DpuVe8STJk7atE3EAkqOXqP80yX8NElxw8Rr2hFBC07CvVcK8dZMUB21M
UhZXUTjNOEnqn+cI9BXR8oklesdVxgT+wUjDgDMxNBdr8mciecESuQ++7sPTVkuj
YDGdXxLeQy6JOvCDgcoLM/RbczCNQ8eCAhHGXa2/YZqtJ9oBU48GelVAB1V8vDl4
s39r8jN1j0fcaK9fmNzc5GMF1V5yW8k/cHQzkLj5bdjy3siSFfO3E2v8VdnaC7Tp
QFB3r8pXBtAbw8geRuDOEyJMYxaWOCN5w2rZD/f2/IHIYajpY4aKlXCQR1CLx9NX
Is759nCQueWZNRCFv0QH2nA13VJXzLqg6oOuIroawOb8Q7jnPzvy6KUyf8aNj8Vc
cenzmpEsqTEMyCTie3lAlE3Kd2cNybkYZb4gywHoQEScMHDsHE3vPnolb0Ewx262
ep8BrhmpCDFwGbOqbTj/bu6q4yXxISeGVKpwitwkaZZju8sRtVmrW7jsn6GZRh78
5LpD8JLcYSD9IKhb1vjikN+HIjMqnA7ai8vBwg/irkFqbBjDYX72Ad04Mks7OccZ
zZxi33C4umz0IwxuC5Mey/zylIiCtAZmpeiGg1H/8GrhTZBQmi1kiEKZyymLAK5X
0aCfWQUypYIEqeGIwi/xE2yyazXBBzPx2NBlwKWEmbVm3FcYUrebA3yQdMrpn6Pb
i40r2UP8HjOXHUrIkkL9Jo/osd+6OvmkXwBsgcrQwXqEsklcXWanVJxeOS4rVtib
zdVAIQ4KVP1tYvDVU1oEnvBssVQA8l7m1SS2iAaEag5jINZaaUNW5OCXDQvY6v+u
gqAD5lc8S0eigFdjRSJRFP5hsEBZ/QbcsjXHvKw80AjpedaGOWkMDUTX8L2sStY2
yrQsFm9JPagv1ZojYVSmeomsQEmzQBpmGBp/0mL7xXeOe47lmC2fCsVEHUWbyGPT
+hVoozn6BOfIm4Xyfsr/g6UovQ8V0vZIza9i3F7UQBZF3JBr0mGDYDMhlI5DmwVc
jhTlzS5piNXVxax4XG2skCAyRIJ8WHk+dxBaK+QNWBPdfQN0lAnm0XnV/103Pz9u
kYekaZd6On8iIJy37bstZll9Ftvf4M3nJYt2LiF7CCb3Un2OO3MAN+uCFmtg0JJP
MPMHNt+A/MRmQcDLHa5KuPw9e6zkJvTy4jd4rgvm98G13AsuYuEURLI0Q/wQrqcW
0iFcmaU7KFXcnNrbgALGpZ1bsJ4yY0Erv5WOHI1M4VOxmDkeDtwurKFL3NzOkD29
G/h3fQ1UCDk30wRhi5QPGNtwyWWvSE/5TacJlU/wX92f/48F8Ilx36hz485kMQ3h
UN4LPPlP3gO83jIzwP/B2FUSGx9w4oWlG8YxL+RrNhBSlSk4HhQMJ2Aui9SDVynt
hN1W3KaCpf51a2MPhTSwe2ja84KmgPrcWvI8ay2H2JTJtyyALAzxk28aBEYELib7
ZngsjmTDlH+2DjYVBuw9njVKx6SN8tInxhSzONYb+uWo1zeZ4iUGNRlXhtwTgYc3
CvZ9N9frBkuH+ewba7miX6ktQ4v51gXZyPo/ruD4pB3BIuEmmI1YlCdbFpeJ8L2Y
MAp95zcCQcDAOh/Vodl0bSuHL1Q1IfwOPSPEn91HpmMaSHhDw5DXWRltzqk1BeYf
9aoNZ5W9M2fyNVTM5XJQ46v7L05FWblh2J9XAhr9YHCSifmD+Sz8o+AT2N3JsAN0
8lJ6gA41EmVUTNLdkArnXf4fl4Ftq0VJfWQMBOAY1WcI9wgu/SvVTCgs3Y3IJD9m
p9ZiIv5YBH24ZywKDUjbeCCZpNGwVXgxDLX9xc7G3h6dOl5KehQgye/HXWdPMI7k
4sMhiAn8IlvT51HlN5Not7o1fAv7lb1teUoQIuFcID+5RWlKtYUkcqypXgaAfkei
NZzyb1e4wmIbAaR3TuWwXBoBSf++irD9ETeI19v84/lP9YYBJ6MSHE1C7Q29558e
an8Uj3Ru8/cw43RZT/Eg1E0lXrhbvwk3J3qzVn52FMxlyfoPtbzbdmDmZuc5I3bb
+wyPN/wHN27vsjRKSE2NsJtjhnpDEjbO0l7RQ/6coY1QzNe+TbsjqvnMPaqh02Aw
jFvBE9i1F0DT49Fkds43jxVvUSIVM+NgJRLahuTtvY2T6zCakyy7KlcI0cskcVg7
aShmrQ3crA3wQh4Tas/Bz7AFLAX1vHPL24O8+6UZ3jMi+aEc/+XG4wW1W+23Vejr
Mp3s2BQ4VpGgIshbkHwflNwvlnA43vveAWzxFanklf0IBtC37JIEj4gG2mMBfNx2
eGYVQEcy45fjpoaTwvHXXt23aWyBCpO8ISoMuNGzBIFMsWTUwuXD0cksnt8vC62b
5g0XkpA8/4d67aP8R6dFjI9KvaUKaDpVSqT7SGKTnhqIaWDJKRazfPlfGztFFKq4
TQsUdSjAS0Oa/uI0c+/i1Cogct4KClnenufoo1GSwDTawFwgAbN8IJQvFpV0yRhP
+NKqU3aiJefbD8J9ImnkrqPbLmnS2HQZftmnzkD6dXdP0I397RZTEjJWMwB/weBL
cN3S+MYBVWkTmZYlZDPTqbfQBFHtLxX4jqGLz/0BW/NWb2PNZYnipy0ZrPUSSf0N
VCoxucWUFCMh9YA5XSE0zW3i7/JYTSWAY0NySKy0JmNUjWEnV0PaAsfocUF/a6gd
FzQGA31FMgLRdTmBb0W8QVhjqZ62bXFJRo3rjSzRK1b4PefE8ChvjKes0payPjpV
lg9PKkqVjRhIafPGNsusFky6cPeMa2paLx5PPRLYFBtUmxTjSV3QGMRAFtglyqhH
CCxgS6AY5EjH5L/dY5eL7rZ1kXqvEsTZyXy/gaA4ja/5lijNAyHbiA419rbXJjYX
tSoGCo3Pb0ryHMMoBEGK2AI8KFFfY10JZhgi+BKP8ZJdUNkkm2eGwU6JydTDZGqA
ILL/P02UEYtSZLW7PSTLl2VI7vTnBM93IiOgTmvFwmj7uo9fqPMHfUaf7uXs6SM6
EsuCcNt88JF1by7BhwcMcplqEkvrhzba5KGDK9DLszc+PJpmvxu5D+t0/oG4M3k7
Ur2jDB/O53Nx4HRcZABgfRsE214SRx2BU6OlNl9FoCUgQ2YkxLv6thBte4/8JHDF
bs3YQNceSTAosuJCvUbGxVhGTlopOFA9BHzeHOWxh/6RmJixjFFmdu/dE8yfn/OX
UIjL0MaQK65nBjHjjwtuwzu0trBONFSMM9gNbgMF4PWU8bZdc2x+GW3SU9E+kGig
CSjkNL09Jd4KVdr9Y5DjzBiHkD6hTsXUUZM++4XeRUQLqcZTZCxOTzqxCQPWPFcq
ldqkbPiFPQIH+d6g3K9X8IY6B3aRnsrgHpmZZZjS4AyNPe6802wgWH21SYtC/rSi
YlgbBS5kqI2F7G3n6QYXqhFHb2KApo83oEEz8bto/MpPGLwFuFK72hNBugzvuXVp
bwHaxEujMftY9k3eGgFBTNRH6IUOnGsGXRWmQRgQF1myAZm2YZORRRhyNmzylK0F
AXPWXaoiadsY8St/sdVC9VXMJHrhm6T6DW1OQTT8qUFdrGU7gKNqwdLGZVG+EJkf
nNqXLKIQMuVjwUy0AfTVWm+Lh5A3D8D2y7XyZSlOhCqYPbzHEnxLp6hexP6ROrAK
ZxLSajiAvifQ2UNBY2P0dDalcBVNM4nffWjcVkM7zrbDJYU3/wyg6nE79rwdxQIU
r1BabaPxAipsjTgoQMx/sDDtd4LmjEKzuavDRBG9qZkHN+pylw5zZYGGlrcemEzO
qMShmx9YfHB3avR5VoZvmg5acq7JDjYWslj7Rls+puXCot/6Y3vh+cyqXnpZHj+b
eYbq4/Ktvo7OiiVEZeu5t1PxAtdwcOW9937xYM/EZyZQAUbnRWcIHN0DUFNlyg6j
e/Ow8He/fXsh28lFf2nZyCzWDw36bmyjbfNFJrlPR76j07d/RKWTxQIM5GVM0Oob
s1FhmAFQgCPXii7aHRMFkVC1hRPRGfyNGtNnrpyZgzzv61cuiqDiV8LFnDf3l/NM
GcELn1U40S/75L+uaUr5Wn/7BnVXmCYB19TfA+PhzoJOq2qltGJYJktd6i20J3HB
0tvi8zq6xxeuS609qNuNqdHPW9IHkb5mo3pLhDVt4XWu7z2YcbCx4b7Ujfvj4Yl3
Z78y55j7DGnY6Qf5AX+VFJu31/QeyJQeAfiN3RNOOwaXBJekLXvfoAEeP4/qritP
E1YvnnfUskLKjR/zAbxAr2C2qHys5+zeAnIqsXJNvD5zIiOOn4Bqso11LARwSTjq
aAqc4keioS2Fc5jxfg1jlVenTCZIU3wqSZW/wIt21vFCgt3j696SW1/4CDOtpzeO
bK5TlGrTR5N9e/Ceewsf8A8kv6AyBzBt1fEJMs/rYipdw8sqohLgUUbfzBnfZOnq
mFgXLnJGyGKC8Bvz3tyo0pDxUw7a83ILFl/7V1jUybP+05eb4KVXaaMlmtxLoxwS
A96qDdrOhTT9k97IEs4B3WSJ8pMcKLw8a0wbJJGsUAXXeQYzRMbSKCPwUqybRUVH
rK4aJfSIe0XAQ1Tb5Bzba4OFO6zoJT9SkmsVDJwHGrNEGADCHh0FThtQI8iXNM9L
RBW7q2kw97gVZswHMTlrteQx2DxZSjERWk/Tgz1A4wxPIHBqb0+Rsi7T6/vF+1iY
P1jfjp1q/+zU6VlBBiJuwodSZPr3OLl7rETZjqz7QzaUEmquKIb2t68B0CanZA1g
7WlooWRFPIfG3KFHlbLCPAaGzacjeczL+LT540TRhIYWJLHsxOW1W7R/eUx4t6jM
inDIp6EDJqe2SoEfqQcZTvz+q8njj8Saq0oOT4Fo2Su7Ijm8Jh524pwYq/V0VVA4
9oZTKFl0Wg7Dy04bK8daI7eJHTIqUufp39WPHuAjUILsJkboYVePIKsnfBBvcu8/
dnMTwmUVask2o2lqqX2MUXW4UUeWZHFg3kIo7pOBlZmcZzgCKjPdzxnwhfcRMXKZ
MD8cIK/t2CVJTOjfOtDBQtPEJHaC4fyTBflRSeapuheuLII5fw9vKMSjM2Fi07j6
XArTi0ruEONGuy8VjsdU54AqOosk11KqWJMcIIntdsi7aVDWAlwuD1/C6kCfbGnl
16CPpgcFLiOIjjTuMKHYfj3Mof2ZBWZyGnuxgbaMk7IzRzArDYmVqLJE+SBB+5br
n6k3CtsXAVA86s/sV0aRqHUQy0/T0q7QE0I0o8wIJJ77o09oeacNMn8LLM1mIlh7
dksBNSt7vyPv23YMGznWx3UhTHZ2m6ZSemI/M/XE4HVJ4TRwDi92oF+H1f5VKT7L
UEefHue4mM1vw5teYWdCQEaWC2HnOlIdqBmL9vBlCO1GtIuzmLOipceODBcxbO+W
LORDtMzqATtVCaCtR5iPKW0WFf0sNQTS6ogDpsEm1LISEJvtmD+MBKNiA9IgJ/Oi
u4NDf3iomJV9/B01x6m6AOiSUIzv0MQUPUNQREHCGJQFGYmpWRk1/CPT87JV9hTH
XpYSlwrLb5vTUh1mgrtIJcZqrPWXlaOJRjk41AmQx490pCd5nPtawVNIbsaPeI2a
2XdXPBSPCKa6LSGUonMIyJvjOS3Nh0E5xlWy8v2rj4PV5CKICxzQMPpKi6G0unxU
cC2QPbAnJFCuWhb6vIF0BIv7BClpo9iQK/x38XTBDUTwc8pruEMxTALT9z2N0GII
Z3jkUAGncWPIA4tCzVORW8rJkNBU4R3PfX8EBzr7KUVVxjHQygnZt+VClclaFEAc
Awe2WWAAkk5MjPbZUzy83ty4dOFUMD84J+tF0IlR4j5WwCYjFqD26kdc4Ro4VT3u
oCQNh0VkRPiqcJXRXRAFen77fdfvK1ayjw0E0xWChrjOJIzxWTz0dgt3O3Ne1PKQ
nNvTN8hEaw/hYPFiCSIGK/IQ9U8BA1ausIWZo+3Qx8PW3qsPDd6yxhgMuOBTbD80
YjMobM1D7C8sXavGNUh4GmBcyH4naaDM9wWSQWXHoquYojAog5wpIwafCHlsf6DW
QRDXItFIBCDebNcvDjGx3YpngaBpm3VhSrWizb+qYv4oJ9rxxWrHpLjAnCpff17o
ZDbNOX2us5JruyPfp0zhWWDIredVATc0UVLIbw/9iE1nKHCi9XS0H6Dh/ZRgbgF7
etCkqy74psFJ/VHNOPyLIYZD0GmVWjHkFrQxNr+filcmcwHoG/AdueLHicUnWm6p
WwmGQyJveZarPP2s+bznLBlKSIAKTd5XkeVU2+WijirIa3nj5t2KhNfbSw6JNOKz
Il6lEQan7qML6VNzn71O00LRWOCNSiZ6X1fBK5PgvFxEMtk6ejq7Za40ATqDXM8w
4sVEIbk5UoOFBkdmzOyTfCUIem2rmhIYoUDvT58x+H8IcUUPhozxApy6OXJTOFR/
SYB+39MhfFAjcmZNGZS9mzXnVaulYNZxVuVvInR8wpJiHdHHZlWAqFMTNrc9RmiX
WNET9egaoBtZ+aKEOyA1h0jIDUNZI20FrkxcmlMQ0urbPsWquac3ZcBTJQ3iDUnA
CEv+B1oM/YgirpW0jTr4NarAYylFwx8l+akkW1s2pSKkAYf+6eKk4pZCfhvsRat4
SwQ+75hLE2McgYUQ8+fnPH8LxvNFP4SlvUWk8X8hg1j4m8Nhrdli8CBCFKYpy0WI
nNNQ2mRDFmswEP9Ftg5fWr0EM/o4SfH6rW9zlcjSoVCbcjKrc0oq8sJHy5fRm+QX
B8s9eYZqXL5He5MZAM3eH7zWMT2chPkPz4/EzswQ9r+gQTq9DmBFZTZK739UlWOI
y+RkGB2JSyRCD9DNnu6rdMRrY5iDKfhvsVXZTtzdRs7YCEpQ4hC7KrjMBSXdW8mS
vnqZvxMqup99dF2M5bDOqcAuLDqNCGY37tRw34ZS2Dtu40QWmZI1LrEW+zTT7YWy
A6gysDAOnpG9Jel9asiIgsYijM0NaHMQI3D2wojfiUflC4Jd9L8LpaF3SHOUS3/i
Ww1IBc40MwdYNkiy6lHZ7buapWrNIJSldZuTFjvxmWLvbSX3FjfHnW3LtwwxPuNh
ufVBC0MdlY0TpMLXq7FPxLR/YPr2Drft+hPXcubu2R91HwXF7USTPVe4IBSqk1hM
Wqw85feKvAmMm+aau9ISxCuNkNxWU2TFtDBiyw177mNnJ3pAHoOHTK8jTpY6AMHF
aABjPHjr4ZWHtJBlkjrbClVR+qAHaQ45lNpkflNgw5v4FU+xmVbexgtq+hJQSbPt
m906lDISpHuzvAYQbZKAPlBO4OVzmxl8UXpC+zLFr3crkTZl7ibEeIRqJ8b9j6aN
dwWxqCau2ybz3hKwNC4L0dOWGgKliHBenxnLmJL+drTrh/FbA76pOMll0ov5y/Bb
He/T2jbRmLd2Ovsgpx4DpWbiZilYzXss1jCmhBsFIGBriGuIBm2EEGae4EVaqGK7
x+YG9s01lhd67gXBhJQ8BtyzNWTQtNK3rli1BGda8ceWCbxwuSpl3/UZR+uyxTg2
Y7Lko8Ng5/K+UJTQkgW0j9N81mXs/Y5Z6e7BIITsOq0blZSsOxnO3c4moE8NJoVo
5rulgEmdwFhGLNbZ2zQPf1o/tNNugYr/NwoqhhwHgxCOAtvPDzylfuCzMZgjnT8K
Z576fev5Hl/75/KMmD3skI3W6kgEJzE3K4t2bzYEHkd6BsfL/M5H/vL7Gd5Ek1R2
qZsudInw/hfleXpAYPFze3arUUZQzL/WEKeG5JEDCJPJLRo1Uo4MiliO31K57133
zh7iY7XoGs741RNnM59kwndbebOnkAVgTFIYZuY3h1ELjkWx0khGQomhYWxZs3zU
xijkDzdDuVKDc+qK2uj3ePCD2may0vxXyws4+1dBp4PWNs+S++sMJxQNo72cvsqF
p/tO+i8BQ1J8w570VxpU7nfr4Dn8jE7s34SiESO4Pcv3zraCknIYnprpsEKJrcWg
iMrle5aj06gHzGIXdLf3W6Ad1RHzMqq1Wu8TI5I0SaY1vSbR2IDdnH/5+kJ/cj7+
wuFhhz4sPXnD/izDKgJNTeJBblB92TtCFMNvQgsgVVoDyhjAL7/8a+v0L3WKy1St
yzMpvAJhM0606OB1TLnX6ZdQE1B7MuXWyCYyN4fpHSigYuKC+ns5UpvKeYbMP5Ot
L8QsNxVMzSEJu2cCdGfOWRehmiP4gkFnjTASv0Jv53o2jijBT8YTByhPQdRTQNUS
OD1chrrCEAV3mnNC9INqCY9aeVikswxF1+knjpYqrwoEvdp1vjVz4UhwJi4gW1pF
ELjtDmk4zqXzrK/GZcHuYzIOojlFHF66iHVQTDI5UwSGnOeb2zj+R21u7FMR5fkV
K316GwKWgRCjO+UmBqQZwjkNESdK89oq6icCOCrZ4Gwhod7ZnKW2YIwiSsc2NmNO
I931eWapparJ2Spwrt91FLew9rqPYyc1lsWj09PPmecSAfivfvzEqjBxGn2fN+Nm
kiTLzBaovZXbc69QvckaLtcJnALh1jeD7hSL3Ty4RfSJZPVOavlF/yqPfbhaXYfr
30pigx3DBBkesiAfLIv6pC+PDaCGRA1Vjm9wDN+xaWjbLOv2bWSlv0d0CNZOivqQ
r1z4+DWkIHLvgM5Ov49qNkiRx5lsujqiKbLatat8pZUxqY2bRoJog5Yb/vr8zPv+
a20d25Y0qcASspRarTYfETMoHHmo1Ixh96E+nECUKztYmh31m4zlL/ZVbNk8E1Cm
4/eQcru6Zm7W746hM7BmlUzPgvglv9GQ9Np7L3iVxwx6OlppmzFaV7s2/LAYH/rP
ezlIoxsicd7uMXYwTn/DHghnHYB9oCFsGDWcz98FSGCLGf01GKbsO4kdTfMTBV7e
NNypEIV8f2hpPQPlaTK7yeGJM9fDKUA7S+vGju3zcdULvlDrtLYh9UbdcunPzEvK
F6DRh9y8vZJkIQoPA+Z0Lf06HbU+KjfMu0qdZjZpRWpIMvJjnn6QJwYSp253kvR5
aRFHkRJ5H0UJJMciD5bp8FI5l9hwJzqmlp4f0vNVU/YMJF2WCk+BdKtd1yuHtIVy
EkwxQtZYtUeeIv+jg4VSN6IZlFa+fnrBjrCdlVFgJFaIQA4Q8JJRlwvRmMTeCyP8
kpyqmUwBOuCrodIcolwBLZF1dG8KiA3iKD+cahdFGkPDeMG3fj19V+1ChaCulaT/
m12THk9jcpzP4bSlaw6YHp0Ka+uMs9rtayjh7OtmAGIBtIYb05qWyCF9JaXwxUOx
ywkv9gA+xzL2A1Fuu56/iZ3MZFy3rgdmobdjxQZWWhICrlMDqyMIILjFIxZsgeK6
p63wAtT+IscMc/nvD/O2vr6GwB8ehuSQcbQulscb0Z2mrksFDM/Bcf6bl27ofHY0
hFsG+FdIuYnyZIiiSBdKvGBqnHGqSIoQv3pp3ns3GuzfeXK5/vQ3p7hkUOpPA7WX
qhe9saFjTfvk+tawByQ+0PjPazU3gatJYwYgPR9N3Y8+TxoM4kxSBwaZ3BqgbohC
fN60zPQG1DkM/YljYDqO876o43AjYZBfvdF+wy9+2Kh7veFs2yNrDSFgWKuyG1s2
yvV74msFQH/E3mFjQCyb5lbiTbxHLV21hR0n/z+Q9+1mI1zxiozt3jj1AEtollRi
3DH9en6tCDan/shpvecW01KCM64PsmGjf47HhiuSohh7obmGDGT0qc67yPqGaya4
vkehHbwBclzbu2NJAUl69TPnZMFOfK4zjYpMxcrasJpgEqBxoyJDl1a1qxq8w0oH
yVRuiKGu3Ta/7YSI6fSc3ftuGvKqZvOEZMuGCrbWApurZvaRAjCaQ/IXxDfqBfQB
Tds2LL6NOpq5U3fI56b3njGMI2wLu5HNdpzFZkdJz/BlnpJiNvknUtN56Mr/c5a/
rID5qMqeg3fW+a9Q7QYrlaJcOR/U4hyZr+2uxaVa4e99WCzAvZbK4cNQigsS5wFI
BSkKBIneNvUG1w9TyAFl3GLXrDrrx3mJUkL79kjXquufxYTSLIJYKV7PRT7TyOSv
npnbfSIkil4fopc+61UBLpv8XVlKpbeBRefmVmJP5gHYsBDMRie9CIDd3c8UKAXz
Q/3+5lFS/ERviywXwP6PyCBDW58WPJxYPLiG8ftIoloiByehNM05xkxmiWuUwkUF
EGEDBcPD5ni0a647rQkBF40OnQ6v76MoAkxDCKqTVvNN7GsF+vFlGxGMTsmcFncQ
FtRdhXO9ArI90oOlW3Hf04QY9HJnFC/TLst8xE3DhsKOI7uAJWeSoZ27SaXowxiT
hRxz3JwlAq9QDVlNmsg145gn+l/QwV1WfjZggt1jriHcKNHgBz1dhyUlFsBzWIkD
090mUvsyNibxLFBJUms48y/Ld8r1/5bwt2/haOPdz/e2nDlILR+lpHTaKnEvFqjW
dCHBIsNbdQYG6Th/EYPGZvXT1jwMXD3d3EswbEgcWfPOMwdbTdd4CC5TxvuLNd/8
s686UbKNifE04ROMYW3Ziu+1VyKkXgzv/PN1TS4WMle84/NZxID6KhB57cqkaWwn
R30giZenhwmzSsSQ7XuKk4B2ORgguxGsaO0IjOk3KR22ZuHW2bBUvwgOSfMUUMRQ
EuTKuPwcw1dD6k6Zh9xQ7ZKDo8mexp7JrJcKv7pVVYYxeAXGTAAY7XxK3v4yqGKh
jZ1PN34E6nUENMxPYVJTWyvnpp7N5G5fnSHdPdUBYvpCIECn10sg5n49x5Gcvn/D
Wc7/rarVNe1udZsv9rCdDqB7TTHucGzH9zwRUIBWw1hf1os44RUk3g52yGw63ED2
4f+qIiyd3mjglrzNmA4oH2wkV2u2LrD89wyB2tykePXvVgey4QD04KIbUfQ6jd1U
4ZkblJIUg8iyhUh9kqFb+w1AsxvUymVbtQchztJYUL3oKMTcQ4EdVSN6y9MOg5sn
BL/5mODifXpdvm4xmq8It4bFeeD9rktmISm6hVJ9nN9kH/sCZkBKa8jPvqBmt99W
VUf3R9jS2+w1mkRAfVOfzPgjLsEtxC+wWdrAwxtUj4DxHfCDXp10fAuNl5d4AbHm
JyHiIPH2DKzNIlArRqSaVW+pbfO90J7M94EnKK7r5TyEzqoxLNo5N3Rm73WIsfwJ
9s0/P1MuYh1MUcVeQ28gEkPmMjuquNeo4JaMs3CSeOd9S05bisaRVS1Zkkwi9iWc
/QlhZ/tbOpUu60uQWMrC8opKvNgPraatU/G2CyTNHkrbKM4Cf5mvdy5aAreTpviL
DCdE73ZjkuTCKYp+cs3faVL8KCYrpU3NcYfAY8R/QUUa3eNBRHp7+xWy4IDcuVQe
VyriLgfz6odxIz/WXFNwhWnpEdbs6crUc1LFPEExOsVXL2eO7Fcu45qfW7NLxZRy
0ajodmpFSUV9Ru4GRgYWzrdEjlKjhx5CyLS3guY3jvoe76aEUjQfwYqjPiaVxsjt
GEwiv4010X2mtHpC75UheZ8Jm6bTTBwqsj0dzn+K4/Jwui2Wpf3S/APkV5lvhQzD
zm2ki02lvZNnyRKN3EPRBTv21thB8MuBlqam3GEemZKIgxO2kRWdBWG784ElVfP2
Kklz3B09L2dUYTdcDXRT5L3M5YI1+ApdJFgEPxO3ATgvTcTzfdgvp1dctpN/gyNK
/R3coBbyUE0nLglW4NhmFk6A6ToBBtuHPH2pruh6kIdeVJ8LX3m3yARevzyNUp5F
+WCWpQ8vIP6GebK4yxT8n/GMUbPNXByMrpchvuPZdWiWzqRmOPsYbAfGMRs6kLaN
DclWp+64wApWnaSyF1h6kdK4KT7g+QrpTG21w0fQ8YSnD6K0LQg/r398HqiGOo7P
urrMK5mT07vA8kn/dkS3950rNU70tTkPcoY61qXW0RlQTvQTbYHmXy/aqawDfJSz
YU29mXlQRVvpSWXelCo9jv+UMwXRDGEDFxAyXUQpP36Sq+pArvLW2QSHC1dfdpop
eGhCfea08ZbeVm/MCPjZLjI7sh4vTUtvWfxB0a9RyVhCMYNU4ZoqsJcekr8C0Yyy
Bf5+xZZdHTFMbvyCOPq2cBVh5W8r5Gu2ru9SDT/MFaoIXBBx5JTdF8lvGoCySoKj
Hi/yoFNaNhr6oYwU7qA8ybVogq6PnAMe0syNbXnqVPvaZGmi174MGnMUyzZC2b0i
kwoGu7nvfbNTuwpi8Gzg5YXL0wcGrNE/w6rEAF642Je7b5V9GpG+ETel6d3Zz3vD
lUvrGyYr/QKrMO0WDhZ05Exb7fAG2TX/E6eXXOtyNtXbABRKgBUED8PYu/lG8ulg
cn7BZahEF5WpIMfvjvGWjZfYJXk07W9lMEerU3kTNP3guuhY9C2UIf7i8S8iqwmQ
bZJSkRPbU+407h9nQv/tVunnFRPKsp9wrtr6qlnewBhsDS5fEVZOCo3ChNNAmYPJ
22Gn569apik4K8l1HkyH3ADmDi6HnI83qRJ1RXjY+XTWV2j1pWG/wNc5nrgkkq8J
nveLy7Y8iMi8EdA+zhbEhjzVOBNptBFdbo9Ho0np1xcV1Xm5c5w49aczPjsMKvLy
mvVLx/bSsfncnZt46LSv5LbV5iWBdkS2kmcNvD61OzY5YV4xd9nzpQmwlKtWThB9
HC2laOJ46+rch57gqXMiQTMpqoCf/FLXI1JhRnNw+jTXmCarFAXC8EErVbl8JbW/
L4F9zemqO6byUxDppleEwrAMZiOJdE0Lme3d9LmQREcbJWAQuxtZ/TAmVUe4wlny
mTB3q6IJDj8S6oaAUiQEs3EVF3trruARR1wYN5oJcPTdKSdC9jmNTG2o6M+OEf+x
23hEGu06HxSUO2ckwimieX8xnXZ+m17dh8ot+nbMuDcc66jH/65LBsXvXYXL9PZs
QG1srJexUpIYK1XWa/wsK/248MJ9cSA3tccqTFOT+Tl6METXpja0gOCJPuCwlGpX
ydc54QiV4ENOau957QoQwinVfSwp/47GTzkUH6IdmDSVDLQfsLqAnvCkHFuZ9Kzq
vi3saMoaFL4tDmfsdOaq3wTfan5VidesDVKiOoYQIG8v6HFgocXozym5OJRXKk6P
65g5qCc12jYvnDxtvvs+4zXijgCAX7d8NSTGDD9HjHmIk7Ld5i5jW+X2V9AXN0cR
JWCjQmCtZVWPHEVj5PI+8HdNTawsw2PNbVopOjGpepXVYUhT2hKqLlRViSproGgH
FtSP1U9bJkD+r5M0vXE23VAnQmBZqGr4Bgb2ReeX6/+O/KvISNHodD2RB7FSCgSQ
LzPZgt8l1j/VBNsKaUAs5nAFvvbv5l/Wf5gF6Ug2I34qL+UbExokEWmJ7v3wZY49
99YBBRLa8eoWVrVNuY5/VS76xOb5mig0WUKPXpt2vCdhadSdD/OLTHebncIivSmw
xn+2h2js+02/b2quCB9LdWxoy2OmWc2PJ3J++3NPAZHDwMvBNFnHL1osJbx8ZRMg
dexuNflMiqRb0A+PY6+cuJ8AXlvpqrmFROBNcEVvSqx3iBiObSdRWwrRVhO2XR41
hMvUSZoVYH2vbtsQqBkxZ6EEzAXzMtCrC4d94n11kbCU5SHyUI3UnZwWrbLr+PHV
J5lFiaf6Ie3wDz63STGUbr0PUlKBo0xkFVZwQrRluhppzM+MJR7/bJqZ7ooIU+NA
fhkBzCPdsZL1No2oDjQAR0hJeXHSctJkTKhXV8OWUNl0BnkR+LJAbIJOz/eBzfOQ
4AFiw1zKESWfO0M1I8kxECAx5ZIEClRAfuY56UEqrnh9LvrqtDCAKZ5313CFoT6b
T21JQeiM9+nn6t5+6dmJNS4tU0MGqpZ+EOA8Dz48+W4xwk+xrGXjIhJsN7QNHLLO
AJWCSYhvFkg7Umr/UabMuA8vgpCxNcmL8n8LSNHCd733NWnVrZMrGDBVz0/HxyTO
HGol2m/42FDn0Yut6wiV6CMgsCKeoHr9KOAgE7T9Bf5ZGENFaodJ78NzZIv6P1ge
OiwcpNcC9Dre1kTXwv/8NyWREgfaCLtj5iXThd83BINwsdYirvP/Usw3ybeIQZLC
GcFRzKzr/FvbX5owGoHCUSfJ0iVz4Oo0xr0tAdAAV4B2GOYGi7MMScmyBapG+i6y
3le14AAFAfLDUcX8WZmu1ZNf9Wbz8RfeGIyF9Nao2Lgb2h/kH42BNNApBtlpilza
SBWGovKSannf+VGFE+u1JLBZnvT+rmfVkDN3GkgMTsKeXA3KtD6goa5gLNj4TTBG
wc7c0paXVPc93HJZVHky6aYvq1XvD7SqrbPJdXn3Tfvzp9hh1xUL5bs2VxRz37Ky
1eOqy+2UnabLlnUIUo0+FPDKfvAZ1unIzug8gDZ8oqndhQoPny2z1hYeYSZusquY
9p0UIuJpNXculU7IR0Ff+9UoWDDzTuLjNCbdARFAYiBiE/vAiRK8y7tw1pKjL5wJ
3qtPPI1NZfmuNiXR1b1BMSElfrDTlIuxwwJdaUXHd5DN25juMay9uuuHji+67Zys
06BuUYqo6Kb7uSbOPeCMp2+jOXulbFLvYSp6oI1mC1o/oFlbGroMDEhKgZnHt4wt
bbW7Iz8Nxx5UGWPT55463THNLjcgTuDEKXl2ULncJHIr69PHuMxXtQAJPhTBz/KB
1zUC/mYXsSRlhw4nT42OJ5h0//XeeZcsqTpL0DwP2T2dxQkjnJCo8hVAxPOxGHPQ
XOCNce6RjHqLMf/cSzz/21eRMv7Hf16WjLqGbw0zM7kZDzzYaFn54bJy/9WwAnim
eTkYp8xhJlCcvrkNr/8MuQdl0njMKU6SQtbxe80iY7xLZABgHUbO+Ck5V9909J86
d8RrL5Lr4ECqDhrZrjOEU2QHCo8Io0iV+UIA+WX9MiroA3xP/YDRuFzaCn0EMvEF
QhQkJ8l4J09ew1cz6cwl4FbonerUWwqYrEyMqgUGBn0iaNpQFWbxgKHJY37w+9zk
P/GKV7bec5ymLE//d3l/Uvdt7mxi83H3/AypN55UBXigpfI1b7ZhSRcRiZBBiMqL
2JgVQM3lQOUlRHY3Rz+8MioOfG83/8NvEPlBKdRbRgDHMvD8kWWXQO80xnyUwYGw
4aTKtQQxJMpahi0ubeYpRtWZ+irbfKjM9IMAKYmH/gn+rmRAmI/pkk2enU5W3BPg
E+WDnT5DK0tp7+XD5o2b1fHlzxsnm+c8sU0FRw6LOl0240YG/uqrlzeWJOvM/ljD
ODwtMwXWHngVctsbkhtrvHT5gSMBoOJ253K4hApnNBTy1GJrrJRX4JCFjWFyPq8C
YwbUBaR45gEAV8u3xkouIZqjN0S5ztO1P7ax0V3r1JRHg2Otw3zysI7XpAHGPlvj
O1DjRE+TxI5uF0eK0JoN3+yRq4lSogIVH6N0831kbeYtL+LglBziDgkbLhtWmzsG
yAfwyLfOAT6R+SxAdP1sLlKDxbdhIalXZ+Yca+MuySHXSAOiXXMa+lVJ8lXrCoQ8
irHyklCiAH2qLah/NK6KqFHdN3o69whCcz5OhUt+Z2Mj2zsp0eQkASIQ98zs8G+g
oJUy3TSh0e9zsYZCbrhwKgTv0yEeRE4i0S1arOWN4KDTLrkEDdDID+qvgU4ScBby
HC8WhWcOUECRnrzwmuDAkSSYzlFk9vlsF6ToYOnFHqkLT9gmHMjAmRsl/cPuJg92
jt3d2/Ui0xtjD09N1io+7KGc5t4Bu4QSA04NjrvpAOFsbqDOqDjus/1fTapQLYHT
kb96Bhn05yYT821AgfvaZTTeBUsbqO38nktXGbxsw5rLYYXWZnkgFGSasDEdIsjl
Uop8vkiZG10fzq+78g8wExzXlDERl7D53xNkvvswy6+eF3MmJqFSS0dLVyfZqLxc
HkSjaec5jrvT4kibReDt5KRxIucJVhKPT1iS3NsEgaeRzdL0bUfKfIQtVUyaF0JX
FBIKd5Ows/OMVRAmHJgVqOCzkx4LP6yyP9ilOPHv7HrZU+bM4j0PGAXCx7Ews9+L
fnoKtl6x928XS6nEXkKmI5qeQlu9VlxUuA17iMjXOGW/fg507cHA8Tq0kYOCTBx/
fV7qh0ffdJrxFF7v69qHHpttSbHFGgz5qr619vDE0vjl8fsRn/6pJ9hm0L2jYIWj
Z1ueaZPPLdMMsQGLauTh3nFLURQMBuTEtjShgbNCnh2ZiTNd5X26edqr8mOVXFF5
ZDw8+Q4LzndJZ3bINY3Yf5/18nsiBIG9eFK+DXtjZ+1SC92easTOZhrM9vNWKYr1
GowRARBJTizKUIWyVr1qTNBHu9mJPoCOLiCNBmjMc1Nh3B9uNV2Y8ZI/gqMvUkQ+
BAbNbnRi8/sLvDKquUKpQINFCt4WFXw6qTHhNvTVO6dTN9iU7qQYKcp8WlAhI5MA
bTB3jhoGqEJetcMYCx31cz0n+jZqDV7+EtzBMJrakCRrZZ/KzQdaiIrBxuC8P5KS
NEPpIUKdvLdETOUovDx3uSRjCSJ+XeMZflCwR5yHL+4rA0knfU+K2orSprxDlVYu
uy7AIP51Sh0ThEPlXILOELFzfAAumYTitrGL0CEf9fx+Jr/TpACjTWYwhgPnvUvS
/ZsZYQkSmBuoaSVbqwVYp5kPm9eqDVjxMKedKr/2Kz4OyF3jsRp4chMgrI1JCCDy
fvSpR4NHaruUVjVw404cB9MkGblSc9GJZRjzMhfNu0is6EvfYSdv9p5IBYLdbCSd
l7S72OEwKQ/vXmJE0uskkpbrXGy8zF6PVHqziw+5loOnruxWblsR5xS7iRxVmQLx
fddhG4T0KwzTg/QgjRICkSPF/kd4Y0+tK4U/bh/5NltAgGSYrGtzCz1zrmeiRLmx
RXEvZWbwvFfXaEBf7qkkEULtAQQKK6LSRk5TPYFz6SbCSLudAofPWdOyQiFp+5h/
IIuK//MJ5HbV8ecBRvbS1Yib98t0BU2HOl84vMfkVUFIl3FGSoeMIxMGYauhVk3d
gDqaWVgiWwmlXPJn2x5iqwCANGC0xyRf5A79V215+MKPXYZ00rMPr8QgHrasoQOm
BEqI9fsdK589AwXE3amNKiYvsXXtnBvLUmCWKxfe4T1+62eI3F2IMGvDcHTf0LXR
qfDHKAc83osAPibqyx5Wmb8X/IWDpBmFNtidp6131fpG4NPX+ZnWV54LVpcylBqa
wyWsbXltM9bkzyzWnDDXSxcQD227O4iJ2weapmVWahT2GB1tv4oCWU6VLZhsG+Yl
Z0KLtyfVfvuX+YnpoVnMa121uhV3FEH68Lyr9o+coe2rrB9o9478laTdR3Xfa1fm
2u2NSiOcSinHNonXMvKZjynCEF2gGA3FnEy8GLUpgeKD5ouMTjz+mzZ0ncRS5uxX
amsyArpTtntYva2a8AY4RF2dX2kD44TliXB5W+HEF/n3RWyqNwBT4cd1TqeaIrw3
PZY0zp+ip2ZXzs4GT9wQlC+YhoXX/cRWv8LlbZTfeWS0DY4jeBFRlSXZzTUFD2jA
HwKarnBRE0qV6bF+E7mngU6xNj6gJQQ+EGsGDPmq56VTtxdr+TxJ1dFCBtAHW+s6
LbN/YbNeDRlIaJIGE9LnxldBHysdNRYZHA67HSv/theJjwwrI+wDHf6kKmRzRuNW
QcBDHP7wRZJNWgOojm1ZFEAcaaOVLhuvJJndSPJldEdprOl3bSrKqjVPM+24zW//
y9u3wZuRRUKqm0ZxhhgihtK5t+yTHwCkI+wJoVFBV8OERh7vMVhE1bVtNaNvcgQ/
GWXLf4hpbDOw5HPFj4MjWVORFEObB6B0iXcCASJuZTeCh8GC4loVNZkCYwyc7tg4
fNwCkoWmAMFAMJE8LKBXtFuHt4xPSzWAMIK4DqrCwhXgN0LydOuV7cgtPChR4SRR
1c9duP+Atpvf2HI1CHSRgIcUmW7PPrLa0nyYGyeigkoLDDzw+EsGdnzDvEcIoZfZ
L3Fj9YTm5W4mmZlaKZw7d1jOpyaoy3uYMh1Syx8JPyQvHGq+BIgs8yPpBP1hlX/a
nLwcVciH8s/F5apiBm2u1EQUp5JO3YqBYjJRjGsMaJTFQHsPFXnDZtB4lL0Q2QeF
SaWZzPi/VIUEFzY+1xfpAhR6v+atExIBiDiS0p9L5TzJJPEhZPHcwwIKgt1sYVSb
5+3E4vhXujhw9/8viix5xawBZ1BPrzfCbGEp+Pd4ivdJbeRkoBz7HHjPEY76ldXU
AsTdVr8WKinXuXSIVLJNlukf0MGn75swJKsjEFoV/VnTnI1tIYeNaj60Ap++y5Fn
qX5EObd6g8LNP62ucxUj8klvKQqWfN8RaNuLiRhnoAywsaMxbusPvl7o95c6+lHz
ceYku3R8Z8/s4l9jCqFRLN30Qqg4+jWfmFgSGM7oXGIOtLYRUsDWP/yBHZFv1lKt
nVQ1UclyoBLXNh7JH0tliOjwzCOse72hqXClT78/3DXOzL3MEgyjKSmHTE0URuhY
5FlbJyN3LH8qfbAa0mjR+X6zZV8JPkB6S2gYQ8jcEj+wqrqZUILskU1UPcVMl3LA
wenvymOkdt7q5JxLR8FfFSZ4d4M7th0nkgEVanwebwyjpRekRt04x6zfb4fRVr3P
LDVDEhPsmxVp4icnzoP7JVhl3bGyjJk4gvQaKYc5dgcurLDR56Z9nOt2EWWxrIYu
/KDfzfiBEerjzCEnSt9t1/luKDPvWD9JjmP8FDHNoeMpj312/uBsoF4x2gnyXFyI
86Bojxj8jZhRfIkVQlIw/FNVJ6HSaIpC/T1T+48hT00tJ0NMdN3EkrLVirv9rI3u
hx7f9ZkwgkOYTMYRd3NfxH9EpMJ6l9xgE3Po40U6VTXgA3jdg9qq1l1vU94Gnd07
GHQQAHtDdz7C2gHf1q/p4D7KXkcEsUTTxQoSe0KRJD8Uu7/4DOIIcgNkkpKyTBeF
CoptvSl8wVYWE6gku5ibNykjkFcGYObCwkta6HyRncnAh/X6+j2EZNTIGkgIy8D7
fYF1CLD4VorcCecjSOK4tDmfyFRroaiQ/ZCErGaDyfGu8TpufLrHNn5msMix4zJ1
bh+6RKgQ4X51toefAbapR6jPlOCKi2O7xJQ1RvgDM/cnE3x9n2SRl/23ro2IujIL
qYuoF3+Rl8Fiz147QJqPZjB6L9wCUPlWslvDXTXCxx4348feCYC7jQn38DdsZIuE
NoOw4fOk1DVpfE0Q18KSabt6Cr4/2uJle6q+eXYXTt19vtwC4xW4pMHd+3MDScyo
PUNePZjr8c1heIVadYcnIHC5lN/uEhy2px56RzeB/QMEW41Pr4J7kZavh+LleWS5
3ZOb+3cn1yNyU0t/XnIzoJWRLqdLaLIunhDxiaz2Pf9tvSQFJHNIZ0mWOLTnesRD
Lx8qyeV3kOtDqbGN/PHlVt80YTM+r3nkLqiiL3mtkijMYSW0rYnUY2aerDyrL9BX
BsVl1X5h4KuIDnrv+WseZH/cmRoLJF2giwRlvvv6QOslW78DycyzjYb1w50/2VnC
8bt3CPuC7ZHEPzEkO2KDHozDAqdw9HFnClTrT+VsdwIb/+uZD4XkWO9xvb5AVuM8
oP9ZsUsom2eCJqcUoxVSp2zmKB06/BI2Pi2M0cG5yrcL0FerCsQIMq6++bXT6w2q
d2nxUHLI7/GN7W2GMViJ/MHpEAoi65lq2pDVBFCIKOhz9DWOvShqQjvcpv0HxK9G
PrjrUykOalbvzzDECnfGr39dZQYdP1Nw88NXAGbUIlK+f5+d/sXJcow5itOB10cc
ftF2VHjMqk227wit+vpH7EgOYkugmh1L6VOGKG3wpbudgzoT4yXw+ZIX92hfDRxF
Nn2GEXL1bZW5UAEqmCI0YB4jAxtX0dKOd0MhDt1g0zS7zBFcEW5vXftIpEO/WbEv
54xyEQ5mCc+aOizvRDBbDM5/DQ/SBr01G8fn9PQ5B7bB9Lxsg0CFPzbEnJZhnvHk
2IaANkzVWArPLG5ob675NTYp3KOJblH04ygt7GfLdrfQCrbIgl3Qy15HQzIy6NQm
wXQLGo0FvuOcfhOzA9iIWBQpqXxKzRsvosEAAJwVsL8hMBYrVT0YrXiMIkMqp1xZ
rzqOZJmUmBbpDsOdJ0aqlnFHjgyJyjmYWzZn+UuRkw1GlFf3mWoJ6CiNliKC7zyc
6Skn7lGMbCcPg5MmOf2FiacGtcr/CezKkPNKu1frpfr75foeYh43U146FeCmCojW
w+aZ8NGE/TGZLXU4ioKVt2AKaPiIQcqDMyK1MlRVfqGwOtjkZcl37tZQJbdtIkVF
Calpft/7vDHfjZO1WOMT2/feiYuGxEy6lr40kd55oAZDZLUV4b/gXPssd0yGj0y4
GHR1J6wmRJZJygJA0xOWiHqSsWp/+8y3HQ0pQjd1xjpOio0pYbqajnEpBVHE+IIs
12rZn4XozXcDis9oDOexlL6wcg/sQ1KHQInn8Trp6fcuYAaDrx1TVtN2QX3xo2YB
wi6w98lp/quch68UgR1WMMrRvcrgcDC7drWWAorcnZTO+ludIEAwtDGjsFfpICXR
7bWNLg+SnPN3GywxKqfdfS1KUt1kJ7GBnIs/fx9tUFe8bHMZmp+1OY2kGa8Crp1Y
varPB96o8PfNcljMYnGiBrRy9kRhC5zBVzO5h7U/qAAo8DWtqDRif0ifHFuF1Kr/
S3Zw9gppKgeaVWWoovdFUzaaOolCYykPMOSrX0anCNYk6qhER6gwhUERSTCyOfEE
d3q+fSL6AMuJci+rZUsACvVbv29au5sOoM3FYADW28VtY1BYFl6M5PPK/MPXDrX0
8mwoT/rPiJ8blcN6+pKTCid2gIj3h2255CfL0Hw7M7kVrqwyPXQ6Ee/PCs6C0mwr
NvjyCmlH6J0qdcnatbm/fNEOy55e3yHURixG5s8+0I138QpsAc5WeiTudXJzlnHY
kCHFkuStHXVKyQSlg9ioWmIudHfe9SKTRl8atRDrCRJTY8wUEUlwjwA7awOnmIHV
9ntKC78rpsBGPNdJnImRjYLPiNisxPlduS4QD0/ahQyAoYxAe9+qI1h5tZCaWSgz
h21kY22p1zBJ+DHhuxZCX5J6IYTOnqOHhqya0DTLo8BgH6ITrkAJ6+38TCLG4JgA
9QjrcdKPOw9YDKFWVEZOnRB7ntlRweGeOZ7wrFGdT+pn/yT5SzLHfl8coRG4kT5M
oN8h8zIbehuMzCOyx4mCrlkQNTMIWGpAOdVjyIDpy8W+vX2tw7I8oK3bNekld1QZ
BdT4/wgdWk34g9cel07+WRBIMJb+gmIfoAGKkg6K9Llhah9Nb1fKGHZ2Yc+BFG4E
Gx42U8GyjBgcuYnrtB0ui/wgDyGF7nQVLG+NfDS6GLXRSaHcA+opMbNSgREebf6l
T4F8LQ/PeN/KUR080OfPNQZ/WHBhXKK8hKimAeooJaIbss8+5DVhK7w3iPboI9dr
pn0Y7YunB69XFHCRaIjUqZPZvzwEIpsn9afGEPW8793fMc2kKiqG9RBLzpSdYl4V
jOtBxdEn71fGovzBK9rkgCx060dAGpza6E1pk/5+CMgQ2rXe+i327fCUTsLJdDbK
SkmeOZCP9HW1wyLMWmV/bRKAGM/+bILNnRsiLvNvLZmMNFjjN/j7nlTqjBlYPcpL
JwmdWkUxHEiiWqB2DensFlMOjezaQmvXFxoxWbDCdcXMK8RBKqlWzotlJMvr7er3
9ZEctSE+KxfGNts2oxJsVDyT4436UJUDg6i7XCfNWTb3Y+ojifyIeogizcMu32vo
TlnuegC4L2QV8BXHSQH1xZ6WGkGD3vKV5izj6/giQs86gzBl2dikO/1FN/skF0Yp
HCXS0Gak6vUh4iGoHhDzi+PADGIrx1s0nPmT/2ODjINVBKzylUWibfgCLGTxaHH8
+8tjMLX3VcvUEhCsmTzdx+GEt9XwOML/IqPYMbxxasWqKWRnx1YouMAAYWhH3T6h
KUWmHNgYUaPPehhB/Idew2AiUF9n/4Briyepkjg9pVwT1Rgbu/ZPRHE3YteC7tQd
4xt6MXl/fApBlNIvQJ7WRBihfY/EjtyZCL9V/wjQXETWHO0G8K4KZUC00WDCpEpJ
ub6hlcBZeiZlqznxIKRGPGAyMUlTf4KVsRf/EHEwjciBmk4Qw4WUieKyDu6uZgaG
t1Qkva3puWm/hLzbR8CajMlyWGvQ377yPGmdZdJ/b6QLWKYtkfM0zDRf3RV53T1t
7VBtfCtoz1C/v5en8B8E0YWRvlcPhuN9rDuxpUxS1eJQ3S8l3KOZm+AYqMbU7frv
9CzJ9tutVx8dE/hf3W8f2OMC+/LKHap1TaIvtSzgmnKK/5cJ1XCLMRHdGnpiyujs
JsPlKd4PiMJxxsdxG8/f+oWD5S+VsNlaae1P9v4ewkW/H4TXdBuqFa0emlVHe696
gK6+DKkSDlGZXspYxGW6f8Pddsh+EnamdczYdqxIMdy6YWZW2MVTZ3SGsTELFv95
mtLsDpSnOGiqiWhLnpFfyM4qqxzBAkBrEQSIkoDnq/KqRjDuW1Cj6iH8WvTt8eaW
Vf4Fsh6yESX2gZ7Gd9Lls93XncdtFN4EyGdLASvS7tdeWni6P1hikWbuYZ3K9IYk
9z66YWnEbrARkCl5umqzSlbhhjpOY+51h1AQo2ZWn0akbk4BLbY9jhqBbU9xKNu6
KM0RQuDXHRkkJWAuS6lLCToz/NHpM1r/IWRKir1kPMg4XW6fosXUJoaSHMcWrRWB
fPLg0VTCjMUPnSWU5TLXh4PzPU4lgLB4B5xwdk86R+9QCt5/6OnL+UhIK3tf5Blk
D2ZJT4/gT49XyvoqtJQEQJQKvFMmcETclSdGP82P5Dybim3oP7gMuwSnhDRPAe+Z
Kue0iITDcaVT0iSjJbjevBgF9mmo2f6oP5g3BeC60G7unJFeAsiGj0hKNjqvkbyq
ogmuAqi42aCPTIHM43cgT1boO4NorUoeBFNpj1Fx3ct+zMiKe8xBcFEZ/sx0X92n
bNWF8RIKAVpSmc7MubTkaJI9jKwly7feB4zUH24TAxAxJQam2aq+bKuWmWBljqRI
hbcjEYbolc1EuTTZGKzBqmk3+eEi47lPQNubv8m5vSkHpQl+uUpfqHrateLFI8SD
cnLDEy/nnG7JMyKo9yEzjQ3nyt+BomP0J6ldkosQqSj77aXv2YknwI5gLUIecmsz
sOvtE/Ri9mXZDUTwBLMO6z8DWv6ew+EMcoAUPh0wcx6QE7iYXLkei8PWEYTn7EY/
77dM7kbnRjnp/Rw58pFROOptGEnUbIMRzPXE9ny9nEVkBv9Nw++OnOt8QHwNrpgW
OhybQmoVsuejmLDBTaOhUQDsqiAyJFrZIIytBMOClw26juwjNSoUZrmWpHH1flnH
B0Hm34QKuZMv1lVNYlHMZSsWy/H+79im2LOw2JNiOa89Jv1XsqE9CclDkGKYGRtP
bOx4F6B0v1R9sZfpBoFbnhJEWBJ5tHle0KMFmO3/CfZ9yh3SN7Z8vWxuzWLICZAn
mg/o8/xZC4UsAXzc4Gz/zek3ekAtKQ4Ze7+TarK96tL4g0SxGThgugAtWgUa7UyV
uqj4+4kCcYho8sw2pu+B2GGzpFVZzovdAzdO0LtiwGYv+AITLqXOcKn7g64V1VMG
9ytSmfC6jrnjqH9lGtbIX8kE+UJNydjuAfGCKb+COrxDPJVgpjIigVbAPMQ5KiLs
+AKCn9te2W/8mjvOBJOPvV+clakC7f+dHbE6/sn0nGbosYypt9CcEdAmumYXTvOB
vPE2/N601+ftL35cVg0EbZC6T/qxiDuw+uYuROikbsKbpd8lJUz719KNs/r6cGdK
u4+X1FOpS9ghMyWvjaaaUy6rHEH9pg0cUTTjITaNkf7wvd1C9MHniUBKO4PG+hHh
Bli6S4uJQQ3JawFw42c8V7t0tyJwe3zt9ImYdQG702JNki4LtWoN2emYFjelGF3A
JQd1nCCbZorA0f98gzbppSYnmzkPn2UUSAM5nZuyAFMoBbIl9TDlveptftd4HQ+L
6TpL4nkgZ1NdpaKrdDVGNbQeNqwcIgIT8lOp109vt9xxcdq79kiHaBjRk+HuKQ2k
DT7jcExdwHeiq4aOFv7csjQbkVIisKmHNjAbYVfm/q1h/D0Ou4PEFAYV9XFX+JAt
oUnZsqmBJ0ZWnYvprWQKXD1t8MuZyjKcq5aDAgEsVXzEy3z1eTseJuN0Hz7khBD+
QbCCMbtYgnZ1IwWs7MFQRM72TxsvctTY9Fcz8oIFzFg5SnS9KDXavaxfRp+AyFq3
fCrUjhArCLjKCvbMJ9VTWSjxneXiqP/220+1UkR8vO2/5e+KlmwuPcWPDLDREi2y
pTF1dd4di3EGrjjxPqnPdCax1/ZwhNaLN875NJ09CGFlWr6LVhLKmZaUnV9za2Ph
rce0oPr77TAZI+bk9U0l4nHNpMDcfh+3M5thE6N3LjSeZf5h42WfKj6hy71Yu2DX
7EhETs+prEOPscWIduKITiiUIKFyfXzH3Bkrt59FHMsDlzC/oK0uOHhAxwgehEt5
W3eTO4yN7mwrd893XqPdCwhfX+8SAEcwCnyoa+2cPN+S/sTGtMjHivCAbS2mxe7d
blQIkuFg65sp7QUITtwp5ZVUAPhhZGLqqmoJlDN8DmcG7WhDDkiLwvl7E9fNNQK7
JPVz8jm74KKWLq1Rhwet3f2UqIGYr4OAc/k3F66uVaWXIa3sL7lk7bfStA2e7qMh
wGdiEZzI0xgJEFI4tBhD00myY01D42JijBHpMiO1q8l1znXQtD7zNV+JmrXa12QS
95q+6Xe03/U4TSKDQ/BU0MPp8ReENHcs8Tlvr9qIat6rMTeJoDP1VTsDA9ip2y4t
iTM/IydPtb9/bcHBq+W7xZTQeOX28gV14A8jrLRGylVMdU4yPlDNmlMd3oy7orkK
dl2cFT/BPx+L5IQoVWpzt7Fd9L9B0axvyzIAfL0gjPBA9dLEak+OBRgrhVehuJIe
F6h6bEA7qhuPmrrHFjBAwmx46NiXv5VU9ZQyGmGlS4uASvh554qPaU0zNtVXEnFt
2yBXa3lgMU/MdjZ1s/vNuqlAmXUGHpWdzuBTPZ2Wt7oqJuBwE9DPmXRdz+PKKjtP
BWRm3qL/GOzBVOdPcxRwB5HoUoRFeIafcwX3/UsHqCImv/sgere30l0tqPiEvyEM
c0UlksS0otw4iZJIzuN9k+9oLmi9yf3p2J95wcXKHcNNUVRLhf/fWQgghNOTKEp1
iBq5ZLo9+qrpda8wWtI/JRw0qAZJc6mqD6q1BwfwD8trexElcDYf/gQ2i9kCswS3
i6mJo1q9alVnjH7ICoa4eBNajOjn0SjVJv7b8MhTjknul182afaaFkdKvl37hHkE
B+ab5VGuOJpli8mRU5LpgmOIGO7jKeE+GMiUL9c1aYCKUoEUUgD/14lzM8lh4Vus
Q/sqD0dERvgRFpU2qBH71lqpT9euBKxipw7mLAiYUhwy7Lr6k7jQxjw1WScMvL6p
Zj9C3Va65FY1qxvTVwmH7Xjx6ZTSjv7wKdEsJu1vNHB01bNfWAEvEPu0lWmwVAYS
3Jxiqrug8kX+wq6bPPfSVqckFcYw9j2vxjYjAa1UNZUrq/VhYXSFOp6BXUnZviDv
dL/YB7pSkquPat/BHMpzcdW+qahheUsIykbb23Y62Wyj4Vk7RNCh9E1YdGN0U2r3
tjIMqo6ibFczbbQmdenhztPkLDSBH5zdyGCsz6S8nnAon1NBiGyJsT/j4XQi/63j
65FGq94fKXLk9aQMNP3Q3udNSTw28Qm+OUju0HyCcRtQeFd9BXu2DhuoNfmAjkk4
PLFFv7Eth4D6QyRv5Q8Ajo6ZuxeD2dnokZCznezE5m6ZhzIHjdYlvY4mL2cJaUfM
jj0VI0QmEMiSUvH6swIL1axq2bgK1ti7GasVOYvEE6Ec08J5o8UUBAJFnZktf9yR
+MsIH5k+gRXSmT258B9TgpYNmMJFeEG2XxgHytG9BCyYs/Ntc8tVApDTN6kHK43Q
UGEElYMq9DphLTXnoMS+u2qqV9GWpPacFwCmXUMyDgGz07mys44rX9qD64Th6qYz
brI7K/PjvLIrqgUI4wQ4uDFQ+2n0WVY2E5qFuPO7huhnBvf9Yynsh8NwcqNaI/do
AVvmfuMD48MCKpinvWgR6Zpw+wWaIkHdxkdNbUwWuvcG0dZGcPlv9R201gIChK46
2cZXsumHIX+paHIzfGkUCWXOU5bM9ZMC5/8ECz5YzVZgSTpkKaJd2ilwNFBpE8zK
v9+Ls08Vaf8GQHHN7ilUptERigEIuIOUUrRZ4Auw2oc3XqFh/x13JDXXG5t226Cb
2kHDM493z6Hi9VsnoFIRNDcOpc2XLKOHzanIqYUSibB3qP1dyjFHCaZ+5Kg5Y+hW
S05mkJz8sOXwkUme/KSljhyqTH7M+GYuUmUc462hYbZfftHORvsPlT/+P8friNzX
jRb0VHu6gRw4SUDOl1uLEDTZUiwKoogjJMnVe3ZDg0JqEyS6WtjUmXuvXpip6wjG
Os/PeENxtK20Tj2OPjdnyIGafGgQwgrBHcZJZ16wKTFttZVvjb1toemEIiFLfqFH
YGBQ4x79C+66fb8IJSnAa7f7kFweJ6GZnybRv2W0YsjlRi7yRil2sviMNEElD5jy
VzgyooeKC1YMFfDBkcyUezv3So9EA7T1YnBpOJFSwxwb1jQ2g+mFb4cRaKXpJJDe
KZarFKiEkaRXtIv3TK2Nq41RK7fy5AzUG2D5Jr1D7r7mrFE99RwELKEHUDqnAKdl
Lfdbrlf3ky5Ni+LMM/Nc1/PSI33ar5wtJ2a1W/KsZGVZCghY6+M+YOk4QhZ+e4cQ
qZt3d0nglD46mc8Vxi5ixAogChHJVkLsyLdgHqqg5VrONSfPkmkHKNLXeOjeZfSY
fVqiEFrOANK3dMhk0V6X6b2dYp05NwIhMIytkYQOKfcFWBqCHxBQvmKfMdxr7+iR
MSFA8MibWBQY80ACKgAdIwCpdsry9z1p7TplT14ccLr2i7j2l9ijQcF2Pf8ebb/+
ts2U3G5Zkw+z24rzTYp763zSovtmq38uMu0aiC5JljmJgJpnAaJn31soVTx+i0zW
TnTpVnz78oAZH3qrvv3GBNd7vUF5ZPUN/8IFQ3dt1CAPU0GiGjvJdGi97V6Wgl5g
qbDNW+VdOXD2LGkiqQ1odfwM8tfDNyZUuhML1mal30BJZekmV0gIJzxOJZoeR84b
zmFbktC7MfwcuqpmExloQ1vN3j9BEghqEQ9PcKwGMiEWiQX7VspGgcXBXjuIT4Ic
rB6L6H1jF/ZIMW/2ww5epe0tA7FP5vzNPZ9/urFdI/vE/3yfcWQGITv4XA68feAb
NVJoUb4OUySFrFjyewAgnRe76OuHVBWMyXZZ3djBlSKuqq7ZEgTV1yKigtBeHLIR
vazz7yGAY5/aqOZS34j665gc0jBw4wbMob4Y72Nq6qdVajM6WjErWdpQ90pBiZNQ
Gli89URUEbO1HdTDZd0DOax0sE8LuI/PJivzhKyQn8RHAWsYNrF29ULYHxc15PaF
/FRcOmjA6ovsDuSMax2pQAkpQJ9KKWQzrnEEPrWZW+VdPfrUNr/cZ2iFvzwhWokW
QEKjF1bxSUp3rCvKJc4kFZjErme2fhM/TcURzUB1AwDQs4CM0DEZoem5iRRx7OeB
xB+qXWKcuiiw2gMsL6LGIm9yoThP4za0jKN2VoLiqF77xSY1AN9+rLvdy6QQQ8qW
hNEP1N/DlOQfM+DOWjhVPcYRenxzCFsZvayWJADAgSipKntKb1bjT8WKPCm8D+rW
i7C7yz+5Hjt7woU5xQVr8pfXv4Vh2APX3S+2RvPGWGcmzMeq5fCS1s6DkNDtn+9m
RNnkFgvfmxFiSBiFmUPZMy0MjwnpPozIm3fUrmQmC8O4VsgB2MDt0chAN9Rccurl
FkmhoVudiVWA7abarVzajexEz7oNXwAQAY0cNUVqXbc0wIY4te7DPSs0khgx5T4v
y/xPKgF40LLJIkyZmmxggDRRNALZ4aEmAM6oyOUMAcOsdAMGSCVZ0mR5ynpaebVo
SBw79Sv+mom3Z8OQr/gLX8YQlNPPsrNbofDZNd0mzONxvWAdq31n9ywYZY+kFCLb
fIWqzBQYwV2+JnAachr+cezs6gAGbIk5F0++fN0dUfJiERAQMGb1N5W8uOqhOO+o
DtNLKJSmZJCQok0w7Ur2/nuplguoUUss9qbYph1h0nGkQguumN38Yj6Ud4NhE8k7
3didq30IQS0m7e4cW9WSqiErxfLd2O8LAV5TmI85DI2V6CtFO/oIOtt99ZlqV9W1
02hPZ1kG/HP6nUZ4xfFBu/9BiWVHerXEJQ8a2JXJadUeQ3u8v0urqeUAaw+vDfGz
XxVYPTRJedRtwGeEMRBN3CpW8JUpBQhXS3dActxdzazyMzxnKYz/VXNA0gX8ZuaA
r/y7PvCrwURPxa3WqwyZdrAx/kqQCnjvJvP8Zx0lJWcOGATDOt4dNd2d5Odbx5qZ
Fn5imUVb27Zk3+qTBV9m5y8UMvYU7NidmQp4KcTIgNuIvtTaVfQ3QGbpPMxEyidG
kjeZIEUNIc9XfV/JFlCfX5NnVz2Jqjvd3T0aUkBDa/IWl6/EhFUx6Oc3YqR/V000
ZOC2EOcqR/KlhWcnp+3SsgAcIZ6WjzUg0UI1tI9C47mC4Gtd4MrboHug23a+61KU
p6rLHOu8uUf0e4ZTH/CtAYhyhR/zU0t4Yxz8Awl5dOOwSr8svR7zsit0YYsxqwij
tlzJf3rA+puOfDw+JMyGf4EFp+q7NzvRZR1szWyM0HFv7Cfr1hJyquj/qv1xrDfF
RJG3rPeQy/2UYFJ1DIo7x1we5Dv2lIXvpw6bB2s5wGj/9DPKKF6Z8NiP+4x45soX
VGAJq9JnguwcA/kbiI4HUiAL/D2SBzRSrw4+Hh3Ot7DC1JZaE79DVfQfIZ5PKhUJ
8IVtvLUQQMYBVoCndPufE78yQjaGQBdF2X8MXYCEjtSQyY4uviTuta73z046/O5U
vf+rmSRPuzjpmMFlhuoDEbuYvnVFjYTguZ9f9ZWr7UGCpF3UzM514SAtLhw7/rzF
faHCT3sQAQdK2rbJYXnMp7K/uZFQAnQv75KxFisOf5CiXnHK+pskmu3hEIGQzIgK
zEU4s9pMPAeG8XO9PC8swa/IvHr/7QAD7bKOQUYZ17K6enQRo+urpWQpx4cYBIXo
ILRhgMdyxn+FA91rdtZADdQd89txwk2YuaCi5tORHYTbB0veDZnHyVBOUNpGEP48
PeVpw5nOzBAQ8yPuDE5vnAfPlvrNNqavk+Aa9FYNaar9nhPVzHdibkv4O6NlicMg
eLNaioCdJyDqamyGVcY00L+yC7GPoXdDd0uiqI9p7H0LkjtbQ2YX1nJxPMLGdbFM
veDIamEpLvd0hy/65eQm7AbxlM/sBTdv0WLWbFysJE6/Sz5K7RCfhWbTvnAvusmo
o5q8lbqhfA34EPW31ylbGh8R+zrHAO95OrfhgcgeGV6JS4FVLxOwmLV01qyX/iY8
yepasNdGyRE8lnKBIogY7vx9v+L1NZnOfgd1oWDCL+o7OLBr/YFs5YE0/QttjDMK
TKen8Z14T07BC6FAZZq3DOo+ntpNKQhDw+UUsalBnbHKdr8yzuKXM02EzMNQXWBx
W1IsU1qO3151H/s+TWJWbN//9L+yEa5YD+4UpJO/TC3eprSIl5ju4FMu628YIwYp
m6ZEbUA5W3L+Wg8mpNAHvvOjJ5a2NpKN1Cc258inMbuWwhV7vTz1g/ZrluISCyvk
1IqYDqPb4wExV5Z0Z7q5LUTWZkbDWbLNUzrJ4PxFrhAWEVudUg7qSSqzc6Gio3K7
VajQEUP/d9BsVimqOCbX7eIJs+P10vjc3N6d7jqzIJqtrMm6PhszTzrgPuN8eaKV
MiBycuURXg+I2uafZWgGXxMudE64h0/x6sYje5Nz9isO+tQPn86+7XXOvPQf59U/
lPq5B02i5MgyuEt4kn0KZVWghVjhbrYCiRRrTSEBB5Et5BR7rkFjP846ssAfI9Hh
C1a9QjazCMykRdp8KtrUkAc0DJkc7KjVe1J30tkMlYOcGxhpbp0Fzmy0Yt3mfmwi
q58UuPYwDkYCewPYY0BETt8HoChoo2poap80TkBvt+NxTP4fWXCXfPWki8a15RAJ
V02ITfTtboQCfaHQ2CM9tlWbN0rZl2AePkpX42m23cTXdvcTuXfH1PKbweyU/tHg
S/w1zfoAnpTjd5aHM+J/VYzpTDdImwU142ejhIV2zJyh062IeglRS1C4lO9f7juK
qSlKSFK9o6TTBbOl+8W4lmnLF2Kw6+NdhDXXik+lV1fy7P4HDBos0EAwg6Su4Kwu
Da79nWr92ZS/WDQRebIp+TC2KAx7wGlktxrMsKYASnoQbb3qUc6qs95ACDKrrft7
wPmeAKMnQ1cKPBsQAn/q7FG9F1saPt9lmON771hDNEjBRXb6FUE2LkbWM8USc0fC
PvECTSLXbZhyoz9X8jimFM9WvkFwJ6/lXyEzYZ6p6eICb1D1p0P1OOzw4ruc43h2
xx5rv5/k7RXr8Irx1sehcXUyZvGvKruTSAlkMJmTO1kQQ5ZGWxp6pfmN6xypj0rQ
dQSwcUoapY0+G9Z04Plz2An10sKDwoOwVIUNCMmsIpRMSVvFfcP8ReaKXwgQd738
xHcTpSUyzB7h4M5sP4P7V2QjAldbUxQHSKnDmUbwJlhUvcmun0451eC1nWANmAKQ
uhB1AMvdvBgWVsEJUGAorPHwHs2xV1BKxo5x9X8BhzAw50iVLPT3I5MdCx1o/Eol
biBWZSwTWByPJlWrX2JjO25V0iPmc2e+3uttc1BTXLev8SmmShyIK+Nyon4DdwKj
+P0vaIX3FaFmr982jh6Ct1ghUNFrk/n1gQUvfAcMwnisATZVkODOk/0JahcXi8RF
7eMBMSE6DZtvD/0ILmGl9WNQLib+2N91b6qLlUQhocf0ZRAovzqr8KbGq5+Ehry0
ncZdbOUzqPksg3Px4/TTb6sotN793bJZqSb8BTiMbTOfEdpVFBkBi2Tc/c5yP2o3
342xayF6QD+6AV4NbmY0LTdtWHSc278RNV+SdN07Ei05X98wIS4OMaStWh61NfMP
LkTor6y/WPbF2rybKIUchbQ9tfaqCiTKcDtZQXWH5qio4aQcq/xddM6zH1trt9ic
mXy4SNKftmHyd1vAmKjRPPJq33A55A1zEDtMPQw3LT2ePU9yXdbE5pBQ/sejIEhE
6VZYZ6FDFEaMgTUt8rRvbkRYW/1CGe/ejdyyLAF0cPp2jbS7jPI6cvvnHEqvfaF7
s4hAT5QnIae1GKcZv1p9IOaG8k+H96GFpKCyBqBidIvQpEX9bHkYkHurRPyEUKyp
ct8niKDeJAQQ/qQx3KyPHwLylJAUBq+gTBJ0BZIlTegZS4R7XaJSYLr10gEA6b77
YldYiJjqlxJW+WPOxe0RFGk3rOlx2p9jibKMJnzANipfKRBpYFShIQ9QX1JZZaHJ
EJlvlJfV//Y8LeEJ64IbDbKnr+RqOiPrORDkcJYfR+T9QjpmH/uhgLcPRRkS0NEj
rFClgRUTmcJ3cn0736SyNguOdOqwp43VskPa6ACzQHmiNBWhg2eMCJ7tITclx+2J
TKvZ3DSGPlQNxl3Mb6XH1nZFcUtiq/IyE4GECtiK+Xv1JbBFxc5WdOC4mLrPXriG
C4ubg7aFOtmu3CyddQEyqkbM4wc5hqcGwzrhdZ1XCwlJcjY1ZewRm8VUOFkt8xpI
tK219Q9ru4fiUN75LizH7vLqx3/BhzusmcJBa1uBwbjkIUuyowEEhq/6lgRdtUtQ
n0dbmELb4243q09bq7UkD9huWPFcMfpgENP35Z8U7F8GaFvDtCXeu0pknIRAyia1
EFS+wUG58vj9NI6sTIxzrz+1eHLfGi3HxfCXnInMtoYFktn3ujOONJdvjnBv4O6y
ZlnO54/L0xT1LMSJq9WkKHSLXdVSQvu8YWtoFI2iYTdnIRuD4oEW1016PWH1qGBx
7nSaXmnsAaRg4VuQtLyRRUaeCoQs3cAngcctR1Mg7aDxmYmjl6BsduMnC6/DSY6+
qRdbK3mMkgl5HSV6+DX6VEnimu57RKEerdERbwITPY1wYURXI+NzWCtJC0X0U65C
4erebhJ+n6mcT4SAM+Mt97AbCPzDOKYMvmBxXGVddUS0S9e4ZxM3KTGXykGDTV5A
iXYnFNptUmb6AHB8H4uvxJ5HpyAvbUmm6ihPUr6dtBedhH+Jvay5cqThc9ibHoK/
8n95Bomsk3khbkhVtPYYvy3iW7YuzPTcFzdZsKgxrnXrjJLKU6VdJ1qLKkU1u2Iv
7xkcehJq7+l8jlB1+ib5RB86VDoL6xHjGJlMt9vzPRbWW6xzuBhBpqu3aWTVwxZY
7gvhe0bFbRJehRX9/lJ64W/Cne0EEnET9XgQ3iUewOwxTtchoydZvXonwPTWb2V5
bs7LYHW2Ikk9vmiibdeisXxnU5FXc4len0ULu/g+VvSP1rale6qheLIQ0MRAQuQK
hQvTJITKijyNFbDkAbAhDKH3l2Jmpioy4xjgdxoJP+cjaVSiBDE/1A9Oqm8CZBn4
BkR72vF0prVMVoJ+BGBrDAD5KFG01NMhph2hCStea76GQdXdV4xpmZzZ2R0DPnGJ
U5zRRqMHs3a1wytCjgswiBoomwG5dRA0jeCRYhXkrZeY5yRxzT+zEnDJOxHcw3XC
WCd/oBlMIjc+jJPlwgbCf4WDBC+zsJ2ksssIVji9/+29cCn4phNmvoQ8OK6LXpTK
PnS+A4HlOZvqK2YJluM5SlZ0hTGY1l3mo/K249cxXRz713lnUVTqKswHP1lQ/YSU
vAhDFeUbpckAMpOlR1eMd2QmIxB8Ug6m4ABxAVWTST3zDt8ixQ2Mbs03axVRiPOx
n8oMiG/kzWIE2jiEItREz6J5br0bXOvUV7SJi6NSBnyniIKxRxXdIJk+one5RBOe
pxlbbkH7DI3U0W611JLV5XwRhCyBBBvRWoSY8LeZjQjEPVSBJpk4QrYrZvSIPHZM
vfRk73k4eGW8cEgMgRWf98fv0f1LPC/Dy2r7lj3InEjAarDYLmlHL1BBu55FWX6F
fV24VS5cXt96tAx6KeEgIwT22AVsDaxFrE2lqY8BaFqRqwkSONRzve1v8S4OA9Yx
JLDE2eMhoffIQzppkzCe1SPVGOjofMvPyLnXhNhsXIRgAyCFHTN3DUKYCsUmRYUT
MvYFtVoxXv4iCNlD8iD7RG3LlWY4KWytiCf2KCvVNRX3OvzGQ0uUa/1FdbwqEvuJ
1qzHGJvF1qCmWm2ciLcDocPHSOlo6H3JPaCCcUTqktQk53jGS/rC4G/x+C6+0bYt
oqb988sMIOrCkfX+k53xjoy9HwYheHTmjzJcLwThrJuDK4tgPTNcYZt2YbuRNvN4
qBiSGGfjehycKp4Ep2f9hBPH3rBN4UsyvXeGOi+T3eLYY14kzwBudHKda1qzTS0i
EcaENFP9gDne4rJ7hBc7CbPI+0jqIHbx4DthzU4cxyTHDKLCY6EXgSWiFiwhWkoO
uO2IiPGkHxCwRrgSsL9C3nHq9HWk90B5yo/Xl4XNKHwlNDhe4VA0lB5aECZxNvkc
19SaTdC0hRCUgI2gDYbE5elN53iOlS1KtIfaeeAXAi0ANDYJ6BHZMmlFFWjdcCF+
EwBNAW+MFFlHvYGviftD+ttUtf8LC1pZa+V5fc0SDw8N3LpXB4gcG5MvkZgSF+tr
md7rlrv30rCqZafJpC95bAsP3kU3wv4h3ipoUcUPjbiYP/qPwf7FMXTp8662xHWZ
gUqEWEEiyi27JjEP5eYaSd3t3AKHANn3K9oYEG93nma6r4RyG6j0EoX3qJJbT5L4
E/22lqhz/1azg7BF+H/3mGPAC0nolxqBfndUD2uMAlffeULf6kyYs8NASyH++taH
m0J9eeRr7XqrY+ZvxbGk4Z5Nn+mKcPVDpexvyvI0B/eXiycJhLgy2Ywx/efnFn8h
cRUHCaaIrTDr7gWkpb8vDNFc/oFk2k5XZawq2a4mEwdsJ2AneBVH8Z3GIcEyd0Mi
r8597b/LCOsJFjPtaIen8REYE2CVkxXmJGz4J24/MJeTEMfuWlqDnJd0tSWuv+Ms
UReX8e+ETtXvR3jey29zNCPNBuu61BgPxxbVVx8FNu8YxtQPQJS/TqXfK+ippgYS
m5Y1NgC/qVz7ArnxfbXmJQqBK9HMtHBWsafGj1f7Wr0AoWyrkvzJ3DXEDewadxDb
mO/0p7486xAkC+M3X5Y1gcHp78oNs8sBnFZgrHWj/uVzg2Je7aZjiKe4+ZESTT5a
KfjaEyPJ50Z+ErlFc5UxILuQByYSKFkntZItF1xy8xUAKhTxvLy6BT1PDlb0v/rj
q9QJBNwc8d+caNDPk+iuVfBTnosZX2EHeZUOI/UTjfSBZZEMC0F9MGwfYRjih6tR
eUDp816ybFced+1G66ipkgbsRubzzH72ZZlfUYeDQ/cOyjKlcQbDoMwKoP2p3U/X
F4aZTMvpTa+e4bk7bnzWeemOwlXd5QuJ3QYItpAltQZ7+6OhuCjK4TrumnT4W760
XaD5L4ZmWruwTsf5TF/H3tvKf1re4sbbbW0ZhphUrS+/W87Z67NdbmpAL3IqHijO
mmzVyW990I7Zjxv4ad/xXGMazO2JjpO8pjwgbj3lWlGjc/ULmj+j5ov4BIYQwjgM
CRg6z5aEJU/0Gr0dKw3WJYWG2g4yZ5ZJrbd85B0W36gk2hCFy4X5OKPKrwvuRSY3
LjERDRQc4xJ4RDF+9bIDvEvyCavFLuFUZBanZV0E0Pf9jl1u4z8qxY+Uhh2HsYtp
d7g+HANKx/QFLIlY22PpZsQuqvErnUx1W4POEt2KymsK3ULvm6XxLF5a4g1IE01E
eI9EMx0S/J1HbaY84Bh/IJvjcC4HKwEHVELfDzD8Ss6J3UBd3oC4KqZrX/D+DsAJ
sj8MiP05PJSZ/bFk5Ieo98HY2gHvP7ckEnFyr7cY2fAITTlf95SGtxexxwIwoDlA
d6NHnbYovFr4Ayc3JonQiDD5F+Ojpt+C8W+ZVWonmz4vF+973Pap0Pa81jlDlBfm
JL5DR5tchWFXpvlUMgi9YSGjFYNKpu5zLoOgVVQclkZq7PHqoxVszPCtdjjyfUC8
vs4oo8aPxRDfzKjDY28qgPKWRoecuqVcT0NyIAM3VrcHtrj7iOmbSk2Mhwz+2wUb
06lphyKSYhBopwTAfMEE2w9A/sfQToCWG3Hp+v6oIk8acpFbRF3qvQlfqGjOqvGs
pVCsuIzs1rnUHtz4+JeSIB1+UNvgL1BmV4AgV1N3euLZY+71n9sStLzo3nXl1tt2
wlOe8O+lgyRTNcpUK/f5+9ncyEywqhemaC+tih64sdU2V6zJn32coRR+VschesM4
ecZdfl+3ss9M0AKumJhJd2JZ6AiobTpcZp7kk/C00RVkKRwMU/mAgxQWUKB9ooy7
TTVd1kNZB60ynG1JTVI9TCTa4guq5cSB0UBoyWAe57i9TmoKM6a2lZmHbSYdUtk+
nv57bdFO9Rv2DR9z028Cgr/ODk7sWGiUyt4K0h1NTCGRHt0245x7Nt6t09h/Ko95
DcPzlsBI6XI7VSOQt2vbwwnzn2UwNhZkSUprpOAAZcsBnwS2dPa8Mc3YBWN2lztM
25rRSXLFtHvGyLUtQHMXxVmsn0kgLxj4v56HPJBgV/gyP8yvXQOSKObzgAsNnU+g
INV/1Izm2qfXCF5InAENhoLGBoYgfnDF5T9mdcO51gBVGCvJ/P9KQD2+bmPCX78H
0lpxWtJtOSr9lLbpdiKQpiMDUV3qCW9b24MT2F2QLSZ+FIrwKvngue2kBtuwXPSE
KdRYdJN1E/ATGcdcqXtot4XSOFyc31OzQS9UZyIsRMgxQfwwYnJje/mVNCfkI/1s
YWTc/bVAvnlE6Oyxr3m3o5+ObdzKcy9NjqQdQQ27wvZ8Bn2huqvQrRg6yn6JZwdr
VUp7Ek+emuB2PGI+QTAbsyQ+4f06z5mD+BCprpC8j0SoCMgndB3Dx+6jKc+m8G7c
fP/51gEYJeXfofgwlfeAzozjMV5INdM/HYPmFXmho+kspqQtxgIyEsdCaTMVTq8Y
yc4y3Xes3DdjTx8IfG5OAA8BGNQA90y1qdwaACNyEftYvnVzC/CHYiOPm5yu7y8e
rnpAo7ZbzlAZgu9GNSXHHpN+Kr2v572w/IfazaIydmpDTYwHqMfVZjzB+shmVCMD
byPtHq4vzUg90U/gTY8TL7Z52D8jypiF9XlIYzxnOelcZfd/YdU21Y9KH3ipyare
aLwmbNxEMLeoNckaiyvSMOiJWIkca9h5X/qokmxxITViDF1P0L04APMEdyB+P2+q
wATtYU03FZVnNalW7il93skeXcnOUA4BL6JEuiHZGmKdgaeRD/JppgskJuJqGMIk
37rtdfM4+vsDvg4TrKpwalhVLsLdx7gDinLg5uuUUhYsC2ZNY6uqzisa97sZ0yJF
CyyJk8jtw2+IBrebMkR7aQ6CnNHNChYhAxjwKR7yS6GJ1/Keihpo/UnwX3RISCo8
OZmG7UeB3PoQOdvupB5xrEEYD4B9BocKb7EsCrZf5ZYg0AZNLg618a1dVjafkD2N
jD9OzYa9IPtTZRil8swCVvKtM86xf3kRaZgunZxPZAvdh4NmngP8bXJeYrXwXPkH
gJa7GDRz7ettX8MeN2ORPVmgB3eLf3gY6EcCNBrkbimtkYWCGoLX3GclJ1fyZZts
or47c9vtyRtIv9aShbKVku6jWZDgA9YHI2xwko4KDOl0ppcL7q7RoaxItYnGJvd1
6FwN1Gz+OPutEY2FdHtAVc77atFSi7kwT1pSYVwBuTw22i+bZWjXxppPgrL/sDjg
COrsbpNiShooMKeH3kMIJi+Zdgf/qlghoAzoVmNmvdpECbXn+Qb+OGO/ctSyIVYt
jFm+ECxNWRFHRkl+jGT4qutxKTRCUnE/cYSmchjpv+0VkUw24KWHcFPqohBG4mX9
UjhWEwq1oj82Y+0mUGAGz8xC7F1dj9J1/dW7181lIIez3B4po8Lrdcpf7+bkcJRh
2IyqWby2Mf1sKIkThsUx4cEqiyGv0f8m5y7y+FFcPq4mITOxNKsFnOXnGY9YE/t1
WK1s8kaKZBA6ZQTbzu+anTBdWoBfKxrGrIV4RC7dtoPcvImzS5Lg+gTER2wv3jRR
jlxovLS49CYYXT4djFUR2SSXDqk90v86E1vXHMsnM672700IQ69tM8TjXP6WHf8V
Qz6W9clpskHeDkfPaNEBnBNp9UOiOuhe51xxNoWq9zcMp/rYgwuV+YpXxicgYjL8
5waNtoQwHznIo+22+umDdmsAGvmFqdBokdIBwWu1RSJjOqp783kshYJ29WKlVDLi
Fp1GqCDcWMz8Y4FHrlHHJKG66nh3ncqrgx0NdR8gpbk3pFdTeqeBiLr0uFoxgu0D
g486SeEkEo2UquCipo6iebsyZtUR95zq62Eh0faNf1b/KgG28KcVE1HSCAhzFcAa
T681n94ZQCzQHi5zM/v6nExhqgW8iAhiJg7OURhfnlftHVPdYjjP4Pm8l2tDcsV4
V8ljV7XYHsLMNMU+P6hVF7mJjkXUlO3yHRHha3dbpuekwjzEBAW7WTeUoWSdYm41
rlGgAYU7KWmxCapFECssV/A4bwPrqiRd/Rnpd3bGEVlUX7tQxIYeOfff8Os7bW84
4pqU7x9aXCN5MphGOHafeykAx9iyEfRENLNMAAXIIm8zZmi/F6YT+REYhgmlw5mT
lMIF5YTnDVfATIGSFEQueb5L18oWTvA74XGDEy877e/9p9c3RFvjmzcOIBL59U2a
3hbhb7AXf3r0uSaNdPt65mR3afH2svYb1bd9rutrKC/cNqQ+RQ0Xby5cf8fgM8bY
VXNVEmUNCKg02VyqU+3HTzQQ09aAYe8S2kvk2FO6L5+lk17tGhC2+ZWf/sjYx5iY
kIgfV7ttcwN8v8D7DwA+AcHMAVCtBg9fds9A1MmnQYSofm/xFRvkkWgyOCFqudZ5
DEDovgjnxPD/u7DvKZP/uW+wFSTnOf2ZeC5q+c6Lv8h8fjUpeGJ98Y6Xr/rRZFFQ
lSTHCNCx9nYMhXluXOQ/T/6AlzJZT78Z8HcNH8zzoLmfbF/penZBWNOoz9umBU1Y
rp/DgHSreGAZU7y+jIY3W/HctJsVpMA8Pb9AiMdAXLu8IdUtjJZg3HmxFGSkwCxx
YnAaTTJ7npPrCU5rlddpZgXFUo2u2OTkyO4WJCZqkkfuky30Zgiebj3fVQxiTB/L
Rw3bgNV1oxMVd3xDUGkDRU5IFL+NiMPg56+wcys6xB63KB+9zK7yWB+VeH+7P2LW
y8By0Ajg1ZQ7xBMIus3VXrSfFk/moHyWDtN2kHUzsqfAn8/KaCkunQucPrQB7xhI
fWw4+Dg/FsVLvlo2VC5tQIa97bGNgARQX6Rjl1+Wc1PCSjVtigyMQIR1mg/GfYp+
jmEcdv4ZbtZ/pSHjUrNg7dLT0IkpXsP+hRLbhj5J5gG9lGvqUhBwqZjw+5PfJ9aM
U/PAUR6KN2PuJjSNejvRrsTzfnm+4owSFp4tad+ZIM00PmlQOzH4AyIDTfq1k0ph
lU4WqEWDxHO/HWrFUVAEbzyBQvSHtgGDVAkDx4lqg9MJb1eAtBMOyzx99kS+XAwT
Pv5Mi70EOQREMtt8+ZqIKzC8JcarQ+lSxlCHckYOdrNTzDWyN/BjUw6DPaHWjG+A
rAc0VzWihIVXrfaWmFrz4/Omsa716J/iYcHWvi5Jb6R8vFBcNewGGVoHzs0KLY47
TxGw4nQ3HryH6POV0uotZ1uqDiKBjPVBHShFPVhc6YGOo0mZImVgaMLvpk8nr4zq
o8G7ErHPJMFJHgQIfWwWn5J0geY4JbYhPzG1rQTcUpfXWSKEmaV7ck3LLCFtbvMc
0vmcmEkMakhqYC27fu+BNAJXAd0iXUAgtZtmP5tuOwfkWHcuvA9NWiLnQUapERDj
W6WIR05sWXQKcuQzRqnXkTPGXV2TfAb9t5QPIas1Hz+RKNZ4CgFhTU+fcl9ShHxV
BCabEKi9AzhudMoY56Mc50JkuIPGzgBJ/Hxxy4SHq2prLvq37fJR1hASusVNhx/v
t7uI/7iXUVtQ1NSoWugLcbOaOxDzA2yoeQzNPBeDnd84zonjjaa8eHglASQwQ8QD
qMX0Xq+nK7Q4FxsV+rnh3pwFz9sI9gm/Xx1ezFQ2LFUCOAsM1ueT2d2ywJGQ/gAz
NSm8gkoSwJhgYw5iMJFDXmJ7xxWjDF2dfjRZYzR6iQ4ozwyW3jcnHq/qDH/l98AT
f4ZJ9FqBJQ/PRzlDRmLIgxy4V+WPaW3vVDth6AhUWhLoEI0tMluiCLDhrjLDJ2rb
t/iWpSRuOvb0p5iH/nHBQL69wyYbev0tFtGa8P+MBMs7mzv9DSOQnB1FLyWyU2nY
rN3MlPUfHiSLUDpI4+DO9pJkA76WjK3Oq9Ag+Coml9snFpuluBfrAxrGiY2tmtvS
lXoz8CO2+m+OQVpzKqUNj1qKIqmBH53dc0oj6uiszimKB/1g5DkHDfd8YRMHSJUU
5rmcdNsL4R4Zpe0Q1xlNViNGR9DXUYuWWB4TBfd5WQ65ujO61OdlkAv4jNRMCiOM
LAoJ1WNb8GRJVVXkoCkx5YWjq4aLz1FEeUqzry4wwJ9g6ehe30UxQ9L2vrrcTQC3
60icvD0gIpaM7MsZS2DTuoqhpTV2AqD+4U4CkL0Z0bccA/RPF2qMPwu/1dpCFB13
Cqg2EM0WJ2qcG23AIN3aGR9Ww7QRfKX61b+CrEJ5akDCSeN0rcWmDr1eFLDNK6+j
6AIOZRE5UeJm1FpaqGjeMf3IGuX+uuLLK1U8ULlkrYx6o54mBkkf13iuviy5GOWs
p7wLc5N0fM4bl0WHDzuuWGaEoJKWcaIMcN4jRddldE1CvmsCULyLHA/XmoGyrVqE
sDCzK230nA0pNNIpGpwcOjHfIf48DZbaVcI8VrpQefmtdUMDJ2Z9ONRHNVALIGIq
rplbYel1gOk4wYbaduXyv626YmZGj9jDJQnpV3e7Qnsuam+EazBMGTF462n+k95M
zwoMflz6tXAFHaRNGP2sWEjQ1i8JFcfIps/1H/4w8QCKSagf3iI3Vx7sovcmy3kt
Hz5IZ9lEJy+goQiSAspOUKRH6u+BYsvujtU4caueEF1Z9LqWaZccVKc2bkTfNEq5
va0aIPJK1v0KqNHhs4pNV81SM6DR5avJD54pGKXY6Wt2rll5hoUsF/pc5BwAgvXL
tWVo/hngq1J5+XzoxwJEnXpGrfx21P3Z2gGK4QFgGKdO6+pqITAgNcIU1yEK2XQ5
iFnA1Bwv5Fh5TR7wyGYKzt5ES35nD2ud4MHTBenUbTvPfQX/qaTz5sTRhyL5Pv/M
H4V5ITAqY9YG1EsPVlOBJWUaE8Vvpp5UyOM9QvIKdQd5La2PgLSr895++EW3wHUH
yp/pjRxCQMq1/+xFEOKQimWSQtDNfqhFU6F7PECb/uKXaUoILxN17bnQKJBpze8C
tQh3Zf747JxbuTHafSAqWrjOg3vjNJiJfg/GMzVm71fbke15fK8b1LVJ/m20Zjgh
o/sscY0KG1GqA81zl9/VOdy3u0srfPYYlWUO+893Ykk8j87PWs7DDOFjLAmHOhsg
5+0GSgUppT9SuRM33bSih5+k0r00NrXculfrN+e2fW+ggNHrt1J01BqqEiuWtCp7
6IDFnFBaAJasqC8DbGP2zKbfThigwkjniRWWSVSHOVqqW3+kxKNe+sKmnJavHT35
RPFLl/L819jOr7T3eeTOqAlGWzPaYlzqgxCj88wCrtNGAyHEMjysGAfXopzxnUkQ
FxQEJP/TMnibVNNGHAiGkRCcWEuTgyY/+i+lW+sdCncbjwVMdD+NLd0eBC05J4BZ
tesZ/qZVXm1ml3rler02m/HiyS9eBujxx2r4tgOKxTRXmELrxL3y7l9R5tFfe1bC
mtt9D8Lb+lavofNFzJcaOwYp9CsRlEmWx9h1l5PGZ65RX8aEha1W5dbBBIHXRwxM
subqEKHowdmljx9yd+ZhjLZhfPHL/P+n+pELlO4G7+5OnHnKWiHSmSuVfctOu1on
QBwg09x5JIts1y4g4N2/Zzx40BpwAHNuoH+20Iede+Gac//dgrMsrDxgHU5XsrIu
OdQO7OR+UHSXI8ZQmJxxv5ObcpYYWOVo01AsMTslTBkbsp/SLf4y81f1Zp15ob/n
5KcJkEKdxLwx8YnI+phE+a54bSr0CGPywYe8hw+gmc/MsC+r7V0HS/jG37/YWvJM
H6VZLrRKlbvwx8Ct/KscaEsLtOgFw0O/utyakX2IfHRnporXnrZwrDSy1N5Eu+jA
d1dYXy2AwEJSVBCgNtmRSQffEa0Ta/C02xWFjR28bNEBOgDcuWlP09NmZMp9qCm8
j1QF1VcsO62gEYhTHj3aL1QGiMRPOJyn9PgQ/V4cm+0KVcwkixoG+AjqDcFtEZl2
Evio6UAXhBD6bLhv/EYPQQGiJvxdBWECAeU69nfebRCxD/t6SLYeH3977uQT4wyM
XQlz9rcQ/0Xym5Q9QyZ3gNUTPzRVNxrFh7bvYAVAp5fZ0tnL06vpdWU0X4b3x/Yk
BLZvFIWI2EeNop+A+eS8UMSbqlMJzF/NyrIV4GFK0x4fnzCY8pm+ALAYh6uxX7WM
9wkhwAMq33rPn/ALeo9Tx4eB12KpqVyNoy7wyTBWamMCqLFAQQmvW8TNvBmENE1k
MxKQ+QtTQWRS/R1OBZBXb/U3RM8TW69E0badx/Fnv9twT+YRait1GNuZ6GMxQDVH
+glpBiBBS7WSb35SBEsiqtKbHmK+ar3WookyHnl0xyqcEzSLaLPQ9FlmeQUlnImp
3NZcoIVjz6raFqR8WF1udB5DhDEZMNceG1JyJD5Ou53dG0kHTYms0vGF6Yt+8d6T
NfK42slfQSpy1u9FkJfZQ7ofPA5UzggxXl9LS+Op84Go0dyM2GpJ8wa0PHlio8km
hXEpf/bJ0hBA0oYrCIey0en4Xr1sfzvrnMIR24xpmeedFo9sIxxwJDQF1uSsunw4
HH6jpjHU6wJ6M/D2DOz3edjS6i6xwhpKDim065Es8EfKsn30NZ3jIRRdOeZBMQV+
U9hFXrKa/SYHv+QzZTueLY/yW4xG7SzaUB1hdcd/fypkfqso1gYGQiHw9AIa7adZ
fixz4l76UAtvtYniAn2Y4LKeEbAYL1H5fk9zAuWX5jV16eZw0LeFBXwt2Y03eKG0
JymZ2AUMM628k0hebsFLLKOjkr6Q50TkjNiPZqJ/0HbUpdyAjtW2U6413Jf+9lYY
UMSGY6exgh51jbTIDAffc0NAWnNHJ74Tv+rtaaWpem6kTmlWVTNkyso55MO5hEqT
7Y4YVeHdPxWEo0CRFkIA5WD6UsbcnZIx7R9n+fU9FdTnELy0xHhCdiSQ1J7/6ggr
kSUlbqeuKQHkIXheGpPy4nR+UZwCZulB4ba1eaSyzIoav8fWdYFp/f5V5ziyHAqD
5LP+Pd/+7XWrzqxZdnuB1aHxYuPxw0Z6JLCXVEbquCPh3OZ401eUvZ5ib6/gmHHU
tv1JKvcLub0IhG9b4ZQsUCIVFxtbTVo4syzVaiDJDQZhJLcC1NLY7Q7YParsHRGe
e4OBKaVM+b2Fs9BJvrz54ATXq54uFK+0zgi4X/jy9R6PE1mGfYLCLiSKKNY8ECuj
y83om59pI2fWvg7M7ZA7QR52p/l8buo+Zfp+Ttwtt5+9i8q4Nqt5+75A2HFTKJZ2
0AsHODqQM/+pVjvsMGihkCC0maZlFtwunSoDadONx48LvTrRwmzS0as3/YrU8mqw
BjHZz8ORPh1iT8ig0zB/vncCgqba3Yt3ocL/6f4G5VtxlOCayg3HcW0jpGZ0+VXb
zjLvYFgU0rdru/kbgcc6rseShJDiqgyZS2Ym4aGh9tiSKmATvjPHhJbKrHg/GypB
sLKyIZa1monHapnLKCPB7sWzUMkHqwMAgpQgx138HVasnaG7CdfZxVRGWJnCPO6l
TRNGggwnelCuPWdkPelHtW/dIy4L7iXq66t1i8X0FviTAUWAZaVhDhR1IdILNY2R
2qjHArLw/GVzZrzyQApPwFl/LT28HTT8HYRke4+3u5ZnGHf+tcOypkhB5Ooln1zE
6vaqf0BQoR7AsQYbPMlSgdx9kQ+9gDrFmnsooObU90wqcimI0lnDcq8pGFTq5nDw
2PPNjgey7OLlKxU3v1bkbTP63iXvyoXLmN5avSaCKsA5tOiyWbXQv6YYZw6HTKee
YBvsqkkjr7uwPoS19QqSaUDCKW4LC/4tycUs9b50LJVmeoJPn200t4eRUkAA5bV7
ADBJ4sUZAfANDM9sftNZ78ymAoBq0DaOcy5ryjn4LMNGlo4kaDTnAXYlqgS0BcxZ
h1wgNAKG3zag1OiMpwe19laDLzSPOTtikJN3m4spN60X1dJgmmMbsXldCLFJ7NDS
qr1qi/9CTAewysLb17g7vkn74E28lLsxFR+2xdnNz9mMwV2Vd1176eVg+HLH1TfQ
I32Xo8Ri4LfUn+eMOPAM+6aCX624gP0RGhzWQVui9p2uMgaXA6iPY0zYE9dm2jcp
9BYGNk/hWu6XX7G+FQDe9OLvaeQGLg6M0afQmpoTFSOhq7KSBujcWMxEroMx52Me
tKSR0N2JwQbmHXQMgY7hdfCDObvt4ot3AHPn2slbTD3JzZ81o7FvMJt1gR0bI3Jh
qRVeGw6QrpqnpI66ftxTlQ7czVYUkRqiu3w+OzoI2eB+AdQ+YZifVv4oi9jc4k+V
uUIhVQhFnj8rtOeir7uzSI/MXxBHuy4QajaagOmIcKVswVyEr3IUYuc8wOKbqV0f
EQxpnNdcekJn5IiEj7k6nPCqo+L0V9h/1tR7SDL9xUVb6MxMiBUAeipB5+/SzyAQ
wSU6ClEGo5FSNedkia8ia9bwiknrLlYbDjyxJBzWmHOfw5dDrkM7uIY7iSWurquT
XVUpgm1xoL2YN4TIrvehyn4zn8FFZ4tVpva3Pi47mukOpd+wZPEuRqYpT4f0ORtF
CAMYbC7ks+kk4ufCkUnH8haEa0JYQYqzXvygajPy50Y8wBAjtTDB/G+bCgdf6iES
liugSFe0xDfWdOomIvIoCW7j3h5IlpdNjiR8V55iLLLIVfqGwCL/FqZQs57kk8vg
xWcL9j0szkMACXYiQ/I+VLr5F60PBZZqStpS6KQQ6unQxL7o+knMk8l70qquxgMP
iLGRHCu8MQB9VT5c27r/OELgoFtjXxh0fp5lpmNPFx5RhHH9Rf3xeWVkT4BQNzV9
OIbREfxBPe7XzpLJWJFZoGqvzv+ivJnPBoGI4yjzGuEQDZS+xamhyq7EVjRpkEz7
e6J7y3UMWfaJqNF0D7FYh6+5fAPiqcOsTSpuE6puuAMTKLxXLZCXKm6OpOH5PZcn
ePD2os7GI0lm2jSf/MER7xdOtUvFnxXhAtuu9j9aUHxdFvTYlufmOYnsDQFHWuDT
VSigqclOLiUeFIj+Teqtcx/89qGlAGKUsmuWRs47NNwMjErGhS+J6P38FvWxHlz8
iCfoSmOa3KKF5eoObYFgeQ0fuqzpUmN0dE2Vj/tGu619zq2W/A9ZCNuTuOi4KkF/
NaoCVEfDx1fAeMa37vvu/NrAbiJ7rYqIAPa7vjeXJsj9RnM4WsRlNDMGUwPj3wJd
1Ui35k8NOoPQf516zp4T8/ytU6hutU3KW4QTBeAZfj1trkeak/dt4V4BHb0j6GAw
2XpFZMx1ZJfGjN+VoBdm3hh9ig3MQUMIUD2A+QQ/qlfvTS+5+uCW4MtWa/5CpzZh
3axku3a1wb1Qh61G5gnVd5/ks5Jd7X57iObVsD+1Z5ngWEcv/f6tBwqFvZUYiT/J
m7y5biY7bcNmM2xNSKxf00VblBlxVABAoBI8Mu/0CvM7Yit+wMMp00upsbBxeA6b
cIktfrz0CfuAaPfenTNd52L+hs/k8KBgi2jdYUOI7Tk0hP2h5EWqQ3f86uYBnkix
+PApAp0XinblRX10dBaO2met/zNpI4Wvjxc7CNL3ilKgF0mAZMiRZTUZWtN1y7AL
WCGOwgK/rupcjf/LIzjlrHn0Pu+zWiA5GiJSnOCJUV7ycjgw7ulZRcACK4hErEXq
NWxggBXpWxYQJscNn4+a5dMNC+qsmCEDhaMgMyTDvtu6tkR6SrwvXgtaibhH8idd
mNl/ijzqKfl0zfKuwVl0pWtPuD48DYP3JSeiI6z8ri8dmkpkP52RYEq5hhigSZEK
WfhNqbOCasA/Yma8TE6FFFlJ3mNn1SAJkN7GWb0n5UYv0m1Y5rRah4wx3Z6uShwz
PAQ3/uJN8K6oZhqHDfyjwJ52bxSEWdrX6WasJFfRfpgXD8oGV2zXWaf4ftxLeuSY
ydCXUdkeV6mfLxg9aFscJYKO8oDBJunfvgUaai2FaF0L0rDKIdIRsY3zOcTeB3k6
kL3In/2+qyMi9vitzE198Y253vQdpYTyq7Ujifm6zmzJfCkNUWSuColg+5TWMO+o
G5xhBS4UbSpxWji/7k9UnBehlEFhp0ivu2tFusY6DRP7ATQqDksB+64qFNmNjrO2
4MR3VSUPEwOSftjboXF7jv0uXYqllmioxs/IfbKcwejP7ZC/+c4oz7gZBzmnhax3
WCBu6i1bJAg9Igr0DKwedarvsENq0vqHr14C/kZIU9+zV0gTT8ddQTLGuARYbrk/
JI63fNFQphh/SZgRfT+MZgPixUu7RKZwypUl0cOsGHDq3CY6y4gNMfO4n5ekrC+u
9pt7/VLQ/Fl8mm+vTiPdZwaUE3hqXSL76XJAZRf6Mlj8KnYVYM27wqsDWyi+70WM
OnyJgXsxsKU4Ad38CMFJ89PS96YMSYCKoHXZLMUUJj6cN2tYLGNSippCGifNgfWB
gCN4kk+omwde/MHnHWrQuKBnEmWhXzvqEfQvyquMNTJixt8HPl4hePuBHDUZt74k
oBwalT7eO1cZ1gSbrVFckOKPAe5RvH+YSdt/0MShbX1VAM0TFFIdqRJgSvqsTZOU
0m83M9ZLAnVYDy6PRGCUJh9Ll7YGAOQF+1fiEJ5MZNau3eFnhAxsXUd+aciCHMjh
opkrhw/NUHuCoutWCIDnkyvApEPDgJ36I+q0pKKMSdM09oLnf6g4CKxFr6BJJa1U
BSVjjj7mU/grimA9T+3FEV8pDpdBxhRsligFcXgBBENzzGY5As8eR8YBwZ7pafdO
hpu2Jj+S9who0FcXjb39M+d+/Q0r1VjgpLwPSwkLpWgNvOKepIeg+ygkeSSlQrpY
zxS6YqTV9/9k3FjYeIO4pqvFllh7/Ji1LUHmflOnSw4gWiHLZoYXj0eevEi7Hl+c
/WxzX6JEVOeJx+zfA72CR7tUmoznrXcK/2M8NLUv1md9TL2oHnpxH8G3m+/l7bKw
Kug3P4hOV6QLKdzix+pdFpd8T1pdIIZChrOEJAxZNox7O2jnJpcp4tk0/JS/Qcdl
jWYAVH8KlJdqRzFIxxznB9OfbuuZRW7KJWsLRx+OeNmKrnFHcGXSz+g/GhfTwrqP
ofrV1++DE+/Elvma1UfNtJnhD3INib46DAMyIAHO11pYQQeaYd9BWbJgF0Ljv7Hk
S4FnerMfdGMPnq2iy0/4hRMudjE0YMNsIj1pQlmq3QObCeU/pJAebtSKiXtR0nRf
NGL9INgAxMAUIrpnlNxQkoi7TBIZ3TfGnWNu3IeDI46aAq8XmkTCir8VqnJxOmJu
davcpVaSgOn5AIJwTgFGxLNIF8ox+PUkIg5kc6mBGDr6HCA+N5anK13WCUilmxxh
V/emFNcmAPztVfluAaToM33Fmqv6ANTWyXuiwbkY4DDYXVoBZMucws6gVja4Q64Y
nQKaAed88Ah1fLqjJm/sFauh4JVUu0R5eE9x+CJxgIBwaG+v6yE3iP9MtHeTrGQg
n5FFM/EMMNrspqXYsb0QNe4wG+wMMYHoYEyvhn/IYyUx3q+uhVYkfNTMkbHDesn2
jd5rGWiuUJIZqFg5iB0aY7AYK67t8xw866XPXpAkTdIpF/NpsNjJxpY2PfLvey/o
ivTM3sEzL2cV7hyvlNokhjXsOr4XIpnQ/QDF3eF5osMQCQg5rdqHvo7GyPqkrHt2
9Yy8wVxqgONvyL9MT+pyO54NCpm6U7/PnRaZ6reUOxP7GW7H0GZg/dVdJE/6HLV2
CC0mQeAs9xAdSmPDo0ibfkiGthsCSkVfaSykTx3deZ+3i8ghD8dDHQBJAghr8Gph
ZYiGdHblKUoWbB2eNdqwmVTNtGqS16CI07ge7NIlmlzd/XGjtAW9CesOQ/Yx/fKJ
bzcgimnWL5XCyn9SdG6CFekXVCOoIbiPRNQkp1k4Dsr/lX8L5Zu+hSOh4pgwOiSD
cHdiBmV7QtVr7Ulaho6/WCqqYYcwY9KjI85POe8eba6QlgE9I7Sagngf4QECXBG2
nkLaZeAPcVCQZ5mVenFXCB8immEtsVtV6zk1QilgmEBe+JFXrIGOoEpNHNA7eHCd
D9rwA8RcQal4Ir8H4YeVNCpf7IgHutF+I1VVtXA7GvBhd+8/VYueWAIlvSI0APC7
Ph/WQTzZLTiiMvG7FsNfE8Tsa17qvz7pN1E/y1ZFl0kpukJ0M4UN8PUqqlsuU0ek
v5bhLIFYpt5iSE/i2xZQevr/cwrYoFFUDhyzt840/9l28o7myoa5pLIHqpq612mk
8T4Dg0sUCc7kkVoumED0unWuLmP1G1rBQPxvgcOj+VcTeZW+l+4CK0Wk4vdBmO6q
H6HwL9I8MHCcFwWX2LyCRWwKvlbJ2SRC6cuuBoOw8RfHnRI+E6ZSSzUWwCPRKYVF
kPUJP5gmfNWM0oMkTvLroVQMDfSfVJFWlUNuexfVhmBkWNoURVnc2ffuYhKNLqFp
pw5MI3O8uilFLxs4jL48a4S8XEWR+cluSiJHDGNhfYc++JR3c40GZyXJV2qCJpF2
Rb1JrWpTYCjO/7RMmFlhQTJ1LRLHQBOWS0XulGDh+F964DLMFnHcWLeNxmdBZTw3
TMp9IZVEd1MUI/rrZNElLJ7x3bcRO13Ggkm2dMFmQS6Genwmzs6qninoqnYtE+u0
XOvkaC19EDK3PeGMuLh3CB8FUuEvf9dLsnaQv9O+HnJjzyDEZ0UWTCYM8aCH6Q6s
xZwsnmBjAfn0YR2JTHr/0QCLiCLp9EgFG8KqRQtt6zV1R2TqCpBeXohzCQmu+UDC
UBpKHsgE9jUwIhpyKsWpreGbRA+oxBcuyeiy+FWHaFUCckXNvciCCB6wX3bOSecW
nADAmR+yQSnDFuw7dSL6i8hjSVHecVg19n0KcXYqmk5uFx6sFkdBcKHN87YW89Gn
LGRe/Rb4yAZnUqwYVy4vr98TEknKiXMHmVX627aCkj6ENYcCDNF32oBTEgUm1TnN
HS+RBMOAl5oqS20NAn6fRroICRB3FWGadd8StcPimr/QWUS9QKmMpiDS5O7hib8r
IodcHCD6dYr9AKM0rDXXzrQHrXJLX3r0L/Y7sWzGZZ+pEcO67gHD/LjMBZ0hnBX0
NGiynXYACo5duGgrrkaEiOgDdMY7N9oth6Wji0xEypAP0yIwKRAKcyesSAOqr1+d
JHy7VEzqdJ2SfUCFQNJrLblpQppWtmrkqEzpul6n1Ee/uUWWBy8HksJ7TF4c3whA
daRvJwFimT504z5an6EG1fk8t2r5rygSuFGJ8ulS27h+Jjz/GhJKrOsbVvWM7duJ
9OYTJZNVYIHYOzVncCGvjcVlbn3zD+6VI33Y84DHJNcWsNU22Qtghadf2+RdquyH
wDd+4xUixYUKWnVR2Hw2AhxNXhqSI5CI7XuqRqqAlCJ/a+98xu4cJ1esH43DQ5Yp
LeAH10AgImM7RkqTEKcnpZMJfloVm91fz24dF4+WEezFVtYzuqsMSNlj/pB0qQuA
QxZ322PN1m392WX3VsQuAv3NJsWO/PKrTOd1eiso2nvRZRRx8HHU5zk8DuikU8/f
KSsiWsY4QLlhrI8EbdNq9quq5r2EIG/GUkFeySnYZCq6HEMUCAGJUebK0P2pDJZm
douYigN0UT+fzoltkvhZh051ISYxDKokYkb2VgRGLEiRtuVkElRKnE7nuIZzHz+O
vLqyycpGw7zAYvdzTLjPH34brUVTmFPl+/iO/+48d3nQRmUsE76VMM3mz6PNFmH1
2fuL0Rlv7+WYEPEOCHw2pfoKa/wp7pcUWuZYAQv31EDJsx+UXCPdedYkxia4o4ib
5V234EMXenQeGEhYIwh6hgD2SjhMAaY3/y5vzLO70R9C32uPyOyn1M/gmKFzKGDh
LoRHfO6L74d7B7If9lDJ8/2DPamEufvozEPwmS6cZ6FnZszmX4MsA204wEo2QYFI
jVxPnLwLXtf5218vIu/mi+4YkKZDrw4QMqGaGjfip9HrsZoh/j9kGcQePynBkyqX
+T0kJUmtfFRR2SGwpzH6xLlJ+pIKau4u8zxTlobQI7OkyRgDz6HqwIcnJ/iYotyC
yZamI7Ta7JeangE6C/ccELZhsilx6ljqPO2sL4DMy9FS0X4Bh5OlOMItmgC89UdD
sFML5AaTZsJ18Dlk9sFLw96RANms/ei0jErgc9KU9cW2TEERmvbNHZRzCOwiKliG
E8etilfanEpRcQq2z7dkRuQgQZdt6m7KnjQExlTZ74/R+n8pIm4ExL7kjmhv1Ab2
haHp8r0zXSVYWbCD2ZHw2xqtCbXWLHI6XHhS+SWPqkubs43/vE9fW/ilCImWojHZ
KmbbtAy4W5Uoy2LJ52Q+o+6KDwdz6RL007/lyEmo64FT0Mqe+SpQSYF73BlMHTfW
IOSS9L9hcadPlMR814BzRXOBWQjQsuPzeqMTMOquZ+absQFEB4oyTZocpfdo+8Gj
mfSwF/puFYlHkR8q67Zy4dmEgEj8UsRf8imocSr215itFxP3V0NLDWdn04rFejFk
573FbbXGQn0F70hMV2B+8BgoUbOxkahymPPx3cOf+iXt7TwYisJFBqepgu0x1gpV
Lf9DsSvO+dPaHz0p1Ol5L19RyAmuF2FgXHUfT6o+oHVn4lT3vM1u6XobsaRvcuzO
Ep7LSWQRAp8OCPzPLcguFSTeXSUac/b8bKiGkzMpomv2AZ34BldGxTYLLBGouGno
Ct9MdLfyJE7UaKGTMHS8dA2kFu7NsMexfdw2wXxlpk9+Vo25ZVKtIsveSHF2EP1m
Aps96CVZpIUCEuGmBUpkPfWbvHnrin0j0FwpupzmK+Wz8h+6wpd6zuu9l4Cz/wQ3
SHrtRoE76VvX2XDyLyAXsoO4Qv2OYNZsRBgSgQL+9X6DDWKhge7dtM9mGeTCRtL1
hwP93wGPbLmFsEnVdmJCASkmyp7sPM2P3U/+zoU94XP5s4tzRWRrzD90H9YPuMOv
3lIPZ7cZSahuMGbb+36fx1+EE8avJD1x+XmNs9/l2yzp49Yya/t5Dp8bDdFTLjI4
WzYICY1G/BcPVyRBSeh2y8HI338yWDsiBl16ZbsDAIFEL9CJLyJmNr7jpqpax3no
VoCKKwGzfAto0Wx6HkMRlRs8rPi8ODhIc3iC6qV+X2nwMtgKuf74FzQc+lXfwHug
vYSxY74eqWURWEraqR79EWnBjhixfxkz1XQ1BCmQ9Nq6R81BfeoxbczZdK7xBWFA
h7thYYkeKTvPVP+P9A1xTL3vAUEXK5PtNkH3KDRFH1+pzUimdBBg8n4f3UuH2Egf
si8pnH75pT5KjB8EaKU5cV3xAEh3mPYNdjgyh7hDusGJvtjjZ47LZzFG+P5BbR1s
IDtcrbRAGR66IR5sx1t9nJBxFkWeHUMBh+7GtjVC2C1s+d0Dq568gWeDIUNk8zTl
kG/twf0tB8HF2fypi7zmic1yCJ3ILz4S4nEgIRXtxcKJ9WVXGzcyS2hIRD1d2Hxb
A67QqEi0Mkt2oiTCIY/OK9EU4PVEA9g/wL/Bo6twJmEl7v0lSbI/ahYy/BoTzyBX
ZvVXlsDJok/kOSEgzveGua3YKIY6Nhhe9MP+B/9Y5BgrWlw1j5oAO3x3csC0AuBb
m4fUSp3FLCVVWJKl+CsHiY3DKHTFLGB7Pq08Epvx8HEK5ZucqljAUkTRRaYlYsWm
semH8g6PfSLLdiv2MDCSr1uLHcdVN17Y4gQOrLxRt/28tgZyw55Ta81DoCXry7uV
H2QxmaPYaXPlUs9fUkkm+2fjB6bjGS3/EhF7U+0IT3bYrWCMKOv/FqtDQlBxQFlE
r8jVaZDyksQKj3Jhi/Vq4DIdlUmAwL6SDcO3qgGepCsuTOFYYedgX2275F+FzVYX
suvbgihNkIQoG0xASN6ryL6bYSrsdLQOaqGLs1v7M0FgAMBmyh/CJpfzwUtOPwLp
/VvkVTU3r9OLpTjzEvlBjzqghkauD2u96noHO0/SIvvajJozM5NWpOmDl+/xv9g+
48eEsl2AOxMxRpge214+S5/WyLCOdkMvQVvhxkKCCp9kLf8XFsNf0NGSpQUojkH0
pPW41qYTXnM1dG1LK8L71ot/7J18Sep5Gocxd8hI6HlS9yPbQDGggLqoN7nErf3k
gAMFmrnZXgFTj6jMD+8qXa156xe2icJ7qCddn2vYrCHXqSMXYFR2iaMIxCwG8rO0
926j6gSEJZwsORiR9gVZcRPEY9H3N8DHhS9L+Y9xpTIiT7/YyemGk99wyc2mh66K
xht5FO8zhV/xYexgffSLnwEP0kvAeH9LDjyk8pMnBpLeTcGTI45dQ7KRNLxCkOAe
9iS19McPdjN2hJSZuSMVMmhmd1jtR7AxAxBysx9R+jLHwGpcX+NOXync9g8CzF0Q
GnrZcScnWshYw9Bg6bWuwYKasNLZZ/aeep08fi4raTVA+4En9+Go41fiAfk+NBFm
oT/Hz919dvdN2s951VVQo93SjDtbKKhH6EyBSf1Qwo7pRpP9W1SMr23+ZB37z3YK
K79p6lj8WDapbL/x3NxzKcvS0D5pud01t/nASWujB4RZeaoATgOfcSC3jk8ybkG5
g6vvUw96XIHsXk3Z8OQVLJaimIUyW9e+eF7gIn+Rm60CH82OecHXlvr1ku25Ebub
BuYFHB+ClHAqj7Wi5Lx0ADLuR/BRrnLZgUnGye7ke3GoBZVnvKF5vAF3zpCYlplU
MhCAwd6Ine+WCjD5aRfR1wY4GVBzDo8p6moXkRWly4EpJhOSTxmB2VSLqZUjytMK
/QjXs5mnic1agvSNWGN2QSHWa4lgyBRCZNWI7c/wnBy8Be55Lc8ahKpg40yiS6V5
xg58p0H9zUDxXG5QAAAIPmml1SRsdRqXJNwi6fcx5hytwKl1QCYUcQ6pEAEwvgy9
HHLdfhoBLzzQKyBUgGNN3KP77O7uFPnyo0Fag5Axr+rJw5EQgan1/JVIF4xtrB5C
kGX3taFkqYaF69TxyB9JEpel749u7qwvHNhfjMl923qNQ45EA2KNQ/anOY0pI4q3
EcFSnz1BvZa6hdbE6rHNCA8esBmSXhggeFkw9wMGCGDBqMh7QJn0id92lA+TMNmF
ICKGNaNbfRfZ3tQujN9XV7Ap3MSAEByqPTDckBMTIo6m22RAR3KELgICdPsqtm2O
/960Ydek9ok02cuUuevjuYjXA2R1RMRwyPEN0E9oWrEQ0DLQu3YTPu+90yqdTvUt
qHLxWNn9wfDq/b5GBGvm8hZKIp6T9luduRKptELl3q0wNrYLtWvHc8Ydyr/rStBr
YUDmSG0pXHSxD/fWOm91rKlq4ZxTj5A1aeNDo7ors2Y10QjpM5YgbQAcSA8G4c2l
ELy4FtKlbTzS+B9XGM4wzQ+N9WttUUgISFbIF2OFK2G7c03n2Qm3CDA/YTogOvxm
mA/f9XQUV0bUQ7G9GHUZIzfCxb5OR15SeZVXiTZFCS5eHe5uONeGgtKHB5dYKVID
5NbB8/e3bcxaQIm41bRVI+kdn7ty/VdagFr/PxzJ1VJbqECs3P54Uyi6u4+9KWQy
7NYCXGb2yeM87BzRLk9Rq2y2hjdLfG0T62CF9bjyv0FWORx1F9QC+hdVnLbdmr5m
A+C8D8tCcI4dSgfXCGu0rrRKDEwtUA0f13OWtMViS+8S6CAt/0FIASFvDygU3MR8
CdytT4ilQcvGkNu7R1pR1gsXiFd/YVhdiG2xGKgcLbDUAO0CpJjysJw/Z+QIMgPr
5TRIi6XIe8+JGJIKZcrK+pb4rf6NZui8HU22hq6ski+wC/Eb2ld+nmwsUq4gfeGG
VbyV4wW/15TxshHK8+jBWhIyXnDMCh+Lf6KZdvZkxljt1OvrTyG3YqA118JOGS71
d2oyxjNp7gRaTjVNMJXIhCKv++JPwInWn0YVlyDlfkt9c94FsRVxH5YgdQS6u5Qs
y5wv8fqGS5bjlqE9vN+stVEjD06SD3v5UN52d8f2jUx6pW88G4DYtXIMSobWNN1W
MP3YRcFDuCVxsl8snXpXvglS6G8OcrnLTy5yZRcIYPi+smbyEq51tFmGX2+Ry7ZZ
4sfy6iAoJ8Ge6sW6lkmOsxunQtKkv51lZpQmiH4cfzkMQA7uYJ+NGUuYbbKSTmXX
8A2ffALkXkhhf1yPOvyAUIgJeYpBQRhvo2dO26zlbRmUDH8uYSXqxptqwXTCYcF7
LPbaulgHITjct9aUEJ03h6jp24NSmjc/4Ny5R01rotaHwNg5y2P0AMhIQ9HkRwCx
3W/HWGy5lmx/mZPxy+mWh/Hj2LjMEfxyx/EpIjhulkcTpgjwFdWLCy6N2Qp+87XU
aDO1MqBGGvnVAsWssuuzm3IoheRmhPaM1b3dzuDm8Q/u2v3ymlM79FULgAeIRPeY
pIH2tSQY20O56uZODgoIwYtwveNaDG5EfveB5EhjtDBhrWiCoHdKMOIliG2cCnEb
pZoKV53ND8s8+BRVZJyhHVEWRHXmJJaQPHfEQTUODaPdDAfwYlPyiAJTo8BIhp01
2YNcVROCoBFDvHMIgp27R1e1GXMdr4drikBDW0TAvqzZTCqgxf/kPhh62LazEaQc
HsCiOVSYZLBsEiCn9dLuW11NKfLGOMv3vU3WG7czSP9don+/UDuC+xfrPS8vyL9q
2QabshQJ0JB3QtligjAzCIJIcdWxBd7SDTjM+KnlGkvwK+yksetifTAQC3BIMykC
E04j1um7u3EHsAY4+uXVhYzFYY78U6TjyG7uA4x7IpVj8kvXeeHI4xqfxnPve5Yi
J+b6BZUvbt2fEKG4tDHYAhVNSveori898vWMKdwHJ0S/+7iL4yUKb4A9Zjz1unky
AQD7qptJ64tSzUvN6nyjLO0mmlVI2THus17DqEC09Zer/T7snS/P4lhIK85lZFsr
M+mxnlaHCqXBeAbEs2gUTP/qjALEl2tpdN792q8CQPl7T2yu7+d7YoYiaxDc9uTZ
GPjVV1l+V0a3dVaZXbyVJbcwull6d0NMW0GdlblXRQIzx35GkaB/XJxENHnFYnfx
Tlzr1wpJ/9o+ErKlkwJOO5mXRbeJTmuSgEmh5uiiCXMvGZFJ5xq3rSblX3sLmK9Z
+qbUMqIJD7Z7m/6Nga41tcjM/WJSBdBF81yho7A375mn5sWl5m8yFO77P+GGfjts
l9EqRcDsfn3GLO+7dh+rvNK+UNvDM7hg6vrzTF+PqVRhFzMs6B+lUUSd7+sK+68W
qCu3n/yCqfOcVgp+Rjx4JsAprsDEVxL95GxCUsD7n1ZQWmO+4vJcEjrIZjdg88Al
XsWb7kyDelX7kyFHkdG/Y4Vf2u/2YHnKPTPgw7cbish38dXc8KLVAX7jrDn8r1g7
ZDx0iorUm/HxNaTEOX/eYY1wLnGRXxXWhnmJrdurQHHg52vDNQnLGLXEreABcnaW
tB56Dlo49M+5Vau4B21lKTW5TGnjly2jNu4zwUJ87g+NVvljK3qPfpUYdyG39+KX
/ieo6PBhmOxc1E1zUCgrhWrC3YaRaV349hp0w76g+VTaBH7tcaIbd23egofhQnMJ
N/rROZwCvhRNUHj3+NYd0Z6LvBxyY0bMPJTaFeeUz14Tz6OTM5fM0HvR152GZRX3
q6LEgLzfPwzHcALRkkO3d4iq9dwBi7koH9fSkwS21ARr9X3byoegtPSKoOgEFyUj
Jk/WNDFmC5nQhbBiPf4vu44H6sbigbzdV7YTCsOAgem2NtZSFb7nMrWk59ssXWev
sk0g5vGWapgQD1LDKzBFxOPmnJUwDB0N6bCcvTHm7uSlG9ZWM3f9E/aIZSHWip+q
d4BmOd8U1Vx+zsxPgAYe+Dfku7mC9d8u0W1edB9T3dESuhWQq/MjnPwhm/2p6hje
4ygaAlV2+7i15d0xf7AjWeDA2ivQGuBUZ8rTbwKnpemUH3Ti1s5NjM9iOICsoC3F
qNRt4co+m/Ixur4kkNiaJ1wBG3wPEwtDmM/xl9LtmculNHVoMqbmo0a9bkf8hu+b
f2AP0geJEZslF9QjwXS16tlajY6bIMkJbUHrtRAxfWguN3n5c2CEqU/8K7F8odDq
KfqMQXB89ze58HIqNYtcbWCvHc5I+708yYvB/qJygED2zP+rreqNVXFsaVzaDwgD
OLAvn2SlQpxAq4zQEY+7rvAv+guyaghH7s9OEEL7yb+mlzbUbDMTN3yuaTj6EpdC
FIdQAtaVA0n1T8t8zwOe0+2PUgYh382DDkcG0rziui0Bbmbm8Jdy95Nhy7QILvhp
qqoVVNoLMeXfLrBbbECmP/nkCcTiFjmOk6cLWQ3VdwMP0lspGNM9WHXcknRdGIpA
ILFIsQTQMHGFzcAeLZ8u2/CJGAPtV/TJQBcVhRmHjamTuU71lE+aH9YnEPld5bar
IZiuTd51Bms/ks/UmEEOBFMrO6PZDpRQejHQUITWBXhOfcxFGtFi8M9sPi6W+ER2
Lx64W+EFslNRU0ZUcOTfcB9rYr230MhytAxWt80t0yQHx5yyfa6zLeQrEQ4n5Oxp
FRPcBCaI+ylF3md2lafGOjt6HYK1tVsiApE3jWzdonqzJ2kDoJ2sCnTbmyXBu5gq
u8CBPkr3rhmzaPBokO6rVxd8jEmggTgNoVdHTgUD/SOGMTigMelS0Y0KNo6WbZQe
vpCfDRKAgb5eL9wn9rnt4mXzIs/KzCg1jyNKNO3PGQ5wYCmRHUc2/YdkCJZjETkV
73xbBD1rx8FhqeXNPSaa94E0piSzwwRa+EwSbs3EM2qy5p7Ey1YY30uCxX/SqT+r
ulcKMTZh3uSy8+szY52N8VlID4JJv1/Z81VRtc6hGk+DUJNylT2uZ7aCCCw1qw0J
tjgRbuSh4jJ+xFdXkxvFhawZ7WInBPUyXBr6sdtoZEUzWmRC5dY4xR18CaGeHiuI
WwwZXt5/QP1MEk88jyGNyQBQEjEKRJ5C128Zfck7r5csrKDfbUjG6n255jeqkw8b
ln01ZH1Jeveq4RbZHJo2bLjRtBXTGc87lvmL/yMfPppMfrwWa2fhPg32yusPT36+
m2C9E+407SLZ6XSs1hJfvBVQxhbkS3wsZ6SHcsXiqlompN4HL/EG+pJ66H0rjv6F
6GP5Jd6aHsbS+9i7LR1xeRa6NEcrsJweG6mIms4y8T/XFxzLUZXFJjAAkywnYa6c
IxYerK9B+HjPV4DJ+bxZWe+jIAPD0kI7scCgJcfF4GO9W+Jd7pIF3eYdMyqhD68W
ggDKbPAQnIzjVCHKHtBQf3GGa/sLvzzPgAUI7NcmVxPjPfrH61wbvzowwkC11d4N
8jS/4Y676j9T/ULjHNEHGKtxXafDIiZBxagzdplLF8h3N6inpuowTJapvS/mv/Jj
JXY4uqJQZE788Vn+yyw6jiPDiP7LDfHAXuJ9tE7YxCsKPPhsSIXeumzncxiNziJA
HNQmCf7idhqNazIty2+eiaBsiYpjlsRgD2zM7JTq5VAe5DHvapiN2ihcttooUtt7
0X+q4OQakx3VBGprEdzm7bO5R1bVQprX8vacW/nxhW1QxyO9O4FaXKXNGDJE/vsC
WzlcFqkPHbrgYSqjLs/kPNWYCpdnaxxI2HZDIIFeUBSwPDWIahXhg9iHiHr0T8qk
OIgjSVppY9AFVgWXXm3qflrxAgL2A+g3heDMcapRBCyCqcS+cGSCmoPjcZq5pbEs
vabGyIWOFHVUSW7tkoIR0MZGCEzj8ptNc/yAi1Ydex8oVTAbdG+JZY8Znxafy7aa
ajihEJY5aPbzu1hQDngfc4PCeDUZfQ9hXQoex/euvFOMBVMI+5XnHLypYll71/tE
A3SRPtcoJ3NO1wfleIFtaGQPsHudaAWOd0038hQuqgodUJwI9jbIy5kytJMqFIBs
f7gEdL97avixMyEi2p7ZyIBGp9SobxMohMJ8yGFwGMZwwp6E0k+My8mZnVuoe+Ub
TE92kdDvjAghKjWDljqXsQLPuUh1MqYTMMVmWgksWMjQUZCtBaxgKqvIa9f+P7X7
4S7CVZrnIbNBtdMZkxk3rJTAj4z/915aBuL6r3vIIj/dLbRMN5y6HRnK3MxXy7Za
Mv6apvJcQHzmHsbUtOtNP5jBCqjyYVWRJaLE2Lw0ulJ6uqog9whyZ3P2XVdj6weD
7/5C2PyTTsRpSFAnglvwOJs1RfBGdQmlx4Q7mfmKwjWTaYJwzpxux33Mj554bVX6
VZa3IjBFcPzeLh2IkLzemPrv3UYYrbzsEEMN4PXpaeiRXfS3djr5P3f6v6e9PyxA
FZQmGac7eB00PvXqiU2VfBxasugzv/TVXBDI0c3MoOXI/EPEkE1IyBYNRd1AY9O2
GDa6pfXCrwZR0ydeVjhYheIEFNVCjiAiv4c1qXlrbsuz78Co8zQOwMIZ7Bexixk5
hX4Kk23fgnjZXuREDouNiziR5Xoo6FlmTglOORxhiaY/ITG/rIAFfqjravSL4zhu
V4w5qkceySWhFQT2Rp+T6hi1sankHWeZ2u6T4qhvu2bcwMkHss5qb9gPxNaCNkzd
NqLaXwLJwSdMytv+EFXi7Bt7oLLPqQm05mKVDU/JS8jMOXrKdFXj/GFpktHnDb6m
7DOtEt+y3gpY64AL3IVTX5Vjo8PePnqMzpwRAtMTURqjREpfGgWqrxM+Zyf1hYtt
Bx7Tg75DnfsfDVT0zMYxnsfi4iAuu7c2zV5YZLaihlflYrkPEQQbbjyGJlfovmPR
eHc99s7pMg/7WB2/Y6lA/FCVAcizF0EGRf7+JxDxHwmsYX10wSQv8+e5EcQXq0XH
x0yMArDp56TWUcLlPvc10qxGjxL3/u2DnF66dPM7ZR2oEU5Owung9FQMPOy+6t62
zwJoib3+Uj7m9aPkzA6GfwgH8B9kx0z8woXfTiBgMoajF17mm6xglxmsqpq6OGRP
fF9NjUl84o9EGLAzWoomHMF1ynPtExTHgdGQIYZfff2lCo4KjE7t/7Ha2mgmMQgh
2SGB/T1ENCmY44RPRivPCgEpAbmLHKgw+rIqP9MkkOkSHeeysvsraUHUghGgD6i7
zy2LnWUyH1NM7OKsfcMf5jGGVvLCbPaSbYmeB6/d6k34itxzAeZd7k6K/4wWBZ5a
5NNggieSm6xfQvrUNcHRhNceYeSJJ0r4vJ4O/wmaAVaihsy9/8+qf3fXhJ19OpER
RADxHp2FsJNetc2ZhwOvgTq2dzChuxzCuVx8hm2zUoVQ4gctmb6Hk521Lq0OKrx5
R1AsVzEMhiSE/SLfJ/ZyWiEIBb+9qLUn0mNEmxiSjCjYPpDkwhK7dHTzXse4/fYL
PMNuhgiIzmFFxlmGdiikcPOyXm8UdCZDRyQMCYjj42ytoshJblSq1imLhKUcDTm+
Vh3x7XTiMtfWyb/ANNjz8hLrV07efGV/UKxwh4CMjFpJafY316gOVZvUa99NPD5F
Ro71liTD79UGic3tWVuBbAoWy50Mpot6TynvHNzGxgeWz3Qbjd5+2EW+gppytYC0
tL77ftCu+ipGJMZaYpPJTwhErwasVjOlJUHsOskZ7sis59QeG0kuZYBEqnWWbBre
s3QWfCv1o7yhdWu2cqZkdzj3omAZ6kSYg05DP8HSQqCGl5Wk7rv7nrxplGyUG1Qe
+vutxeNKmntSUCoguObxFZJdlvDG+ktSGwjAWiIOiIqvmASIRhtl0qpuLYXqS8Mg
Z824DhWTXkxH+cbO33SxxKXjfgt6IWT3jfiZdZgzZtcJj1GJ+n9Xo0O0hQk95PRf
3fM4u/fByFty1yubXhd2Hmy1QZjjQjh/zWpC0xaV577lqRyZcwJkZ2Kzqrw2caKT
a1IUwjTjxI9pikIUy54/vrZWAZovaHjJlIpBw2uQDlPP9tX1AE9A+lwKU0zeIBf3
G5dTHrgvdK+R88b9DAk4z0At0U8kssBbejMVJJ6oPWXWNqOBDzq3uZYm7woS0a5/
i7FgrfRM9aG+rjocg0SULx3z3yo8AjXprX3q3IZfGUeb8UcMpTOmSWpEDER1J6od
XBj7xA7L0sAGsnkkqnte6Bp74A9MpyaBG7SPd1cR0KwlPjhWdRv3/WCq4HvHe+JK
cv+bFDevVlKddy7nryMcsDOPN8vyWxwZx5qN/0sRgr7bTUVs2QmYydghWVCTDGnu
aH2rdKVf4LrmoN9DcDUqrDaJjis8UR5m0+pV89yP7p+VmzhTsFaN5BAY+ub2uhKF
4z9BDBMQ5ROP7HbjP1FWBzPJaiish4uzJ7sx4NNXJkXe9XenKjelkyAk4Gxlr9Ym
pLXDvODhqkvBccK2cvSj73Z2F74jMEOhwLwvjMv0Olwjct/8GfT1RAZ1dGpbcI/3
kQpFUPANQ2O/w+F69004qcCgLc99KsJtm8tI2NrwLsi0QjNX6JTfTf/cEdk/e0C8
+9xeyzK/2agE8kbkldsd9mOwfLsosMhSON5j0vaVNhsUbK1+/4LAB3qBKpkYZL5R
sRNG3nw00+s2cizWbCMhA4zRtTWrrYqhKMhrkWjKG5+JBZamExG0xERGH8t0RI5O
0RwM9BzUdTixPprzyyy39K/k2YNVCUljM8bk7BxUBNCIrWc28//cjc+qfdGXdjqO
zdlIfuh+nIesWvay8eH/MU4gR1hQTJ84HfslOfFjqjO7r5hqcu36GwOkaGlhn7at
0pDi+/YjoVTqpFWXD4d3An19UWHupVEUGe8w1kkxExWuwOLx/bPeyNQe6Cc9O8C0
1ZntrcV/iOs/nxgFrrnI24MSaZHSmmR2rHtszfj0+h9sCouufrHe3QoyRixBGbe/
RMea2hPIYEpCdjRn1NcaPicAVzir2Jzjw+EYNS2kkjHrnzp0ie+gt7OYCVaq1Rsj
h7fiTIv2h0+HcFWFaWuc8rWdiLDczRqJdZqLxn4n+qakWTySvd0XXWPyFdefuWGP
qX2pQdCtg1Hil8NcteWl/9L+uk2T6shTPATtZo/MPAj2jUSYMN7Y00M7KjICcY/d
8n+uGCrgPNhZb2MjQwWBSf1xO6cSt00Gj1UmYRyXxBYgVKx/Rrm3APISlO8HadDH
GETtrKfTAMuwgoKKbxw78f5eOLfs718AImFOltM5U6FWpsZOpv+t71+UfYsGLj4C
wpYnCWh9XeUTv4VR8CHSJy3csfK6K6lKOYeNZAfSUgO5C3VCiQ6NjZoZq4cqWLxL
4btoZyzEU6OdpoH0bnKI3SvdwaKGJGC3VuubKAJN0lXPuvNqfSTY5GBxa6weUR7R
XX4UfAexceNX2t+YInyUVsjLpAVHz9m03B0nimSEJKkQARlT9Ze35wwjifzTF0lW
X3X4u5seRlt2GekthZDU9Q2SCyAYr28+hJCmpJ6XwcIt/mEBjZ27i7ZWR4o6Cfjh
a+tWcWBhtsKfD0eOZbukChXIavDzQOsxPR/q6/Pd50tyV+hUTkiXFqkL3m3xSC4o
LnOaZZbPgg8t8DdCVIlctwq98c/gy9PkM5lsGyyEpgKshRhLE77iO+XdXVs4A8Ey
F7YXOSVK+W9mSZA0L7HhTTyvm4+ER7Jw3HVb2Egyx+cRVYJ0aAjW/ROm05VvlXr0
LtZliKUxcc6RYH9FRSOzC8axp5pv6n/m7JAM5d2qq0pxHuPXcJZI2rqJK/2oue6H
e3vJNifDjZqNx1eacbCXSjeCAJcLNFaIhKc3CBHn5OkYyiKPkauEkQJ1dr460MBL
ubrrD5rTUlgkS7TWsUMCi8vJRxmCrMXRrhVvZMa4rbpCmh6LzwNGcH2pTvkCH7EH
kmETmqpP7Hb/830nJh2ppZbbg/i8qHtM1HJgwiJn7DcVTJPKt44annYuxAKIgnhJ
C7c5PGC1zdBs/F9TXY4xejKnywxeUcpgGz4FjeZhPK3STK6qJr8+gXfeCyscocE7
3rFmqB7A3HTZ7tFUgvleL0eP2ZDMIvVWVpb+FmuiTTVJ/v672DyZAAyWEh95hQEd
Sx9Na00NQkeQBm58DPo/L6DeTO06DskepSm37dU2Hnr/DID/rindixQ0V5xqkNzj
q8FsmY0iP2u3jX7Xk57TjugCslkeIwSfbr5rmDvNzlHsB/h5XvqbhauYqrGK9lwV
dG0weQUSFuw1B11rPw5stOuoZYh2r9XNCfrtidsFauN/OxhY6Mr3BRsF6Og0PXDu
Qri4TWfAXOPdi0hW4Ye07Sm8O2nYQRkTWL7cxDAEpLhVCAoRjtjG/WtUvyBnfxZB
Ha1CHzSOtkyy53o8///XWLGLpBla/x+08aEDIEIdzG1MFplB6JPE4VcvrNJKwTYk
0/jkLHj2k6Cp7ShSSDGp+SXE7YLiHvcxHjqIMjnWy+XsQxyYgWQelXUVRjCBol0I
HNwhsdrk8gQbazGj00Q5upjcXSzMQouf+japCjsbmX/UpPII+mzBaZ5VcI847XcO
1PHirMgUzoIt7aKUwAje2XxNjasFUmtg/xXfL2Ftq3Hzm09JlDi+KOgFFiuPXMru
omOZHdN3HWZ6+ndSxaXYgeTsYLWorst6M3lg5kj1R5FFRg+teR1p+3tLr/x3gG0a
xdRHakqh0tLJrjWlWY6sIiYhmjx/nArTv5HpsVnIEYy6U8SPmir78S2v0oVOnM6b
Z5VPZTaSG8QHEdJ/igSdK6DIjRg+6oOgqDHRBkk+9tsDhr6M7Y5bVSv0/09CZLSh
5vprvvCuKyEDoZcnxKJBkWpo/RjIc0H9wkY6eXCHOnDnDYbp1F5b9dRLE0FyJpHW
HTj3brWnDIDVb9KkjCK2DUbvQjU76i6Ak6jPw5BFfceLfTcgANnqntIvgSeW0N7F
JaCnPO2gZ5jDKgmF6vWw8sXg2rZyyUs5r4UOoAbJC39l34tn2uPzsSh2D4fgCcu4
GhKtb5wpchSnkI9VfWHF1FjWnhvDucXNQQNiwRSOLiRDFE78mXdoZwwYbBXZkWbc
RLUEOqmrOqVRY3iVPydWFsEkUw26GA9ceo6uwgye0UAI5SJnkxYGvuyHr90HXxbT
tzrm9wR2IopJVB+t4IOVxvZ8/WQvQFpydhE1ihY17cF4ompCKt3T+C9X2HPtbk+1
kR7I211qI5mN15uS/s90e2ZmGogEH72aT6ElP7NNXRrIgEbN4BI8PUa6bWT4yyaj
0oMg3ioeZqX1t6WfUpPtUlgO+oRHhREcwovXt4Xp3Y53oCbMIcT7P8Av3FS8Zeks
o8PjQ53Ezj1wMO+HSH/u/J2JO6g+4DGAslErb7vM+EzOEoAI9iYUmtEUG5gQpWos
tl4ZmpgbJQ0wivxDrFgs3i+J81pKvHtsDTa6tlCszXrBb7IBl+5Zgo517B3oP4bS
qaDQ6FCMGIdKw2VZ/G4TPWwtzR9I39fByl+06hwMdYIEu8vNkq1fpAPCd5V1hYMJ
LcG8SovKjdcLDjT7g/Br4gZhizEXS1szJYv0m1VxcecsRjNJFo1BX1yB4Pw8Jr+X
4dvuKF14gkUFKLeQ3Yz9aoKBqNzyVD90B2DVGMxgyPdVMQv4NmkrBkZEKfF3oeRe
xsM124XSRcc9ZkkE3r0THHfGKHoQFZuzmTZOXNnkRQThmeoUPZMUzinlbKOXhetc
rx9DkNHDHS6AJ2I649vhyCO9tbzBiRJLNJJnyATHpVW+3kbvbxRA0x9pLHwlObx5
bjnxK+OZsy5YBkW8fEZTPxGWmRJPXiJkEowrmpKEcDEIonlcACCx5yBBBZUaCg6T
V9RyGb2xwvYRwJOGuCioLi2l/3GV75B53jwdQnOcsefR9Sbu9AXQCTujQW/K5672
RTXIJxcvDzcrL10z/5D0g1XDmU8JqNeTJNsB6mTIzXRX0v1T0TiiXETvRobYFUWS
3mVCJU41ly7OaOpFUKJnigFR8adkEmMREB8VHAvnmva5gicRyGhqEs4Wv4MiC0qK
tl/vbh7BRUhovfG6JdI45T16BOwmyvVha3ltOvty3f/9Ce6F1NuUWhb8gkQHFmW3
+FI9vp/umKjP34xPRPzBA6zX8I3rtcBXCScWKTIAWHEHhza+B0RhbTQWiiv1pAAs
42XquMS+WBp3HJPA8WhzPtVdr7dbuwzbkmsfZOHsSNzrpmk+EwflykEQonYBG/le
xqnZlOGLmSZKi9VdAh3+2c2qLmdVJZi0beku8chT+xdQ9h3geGciu/IbIvcKSvme
UHGTrPRBDal5Nx+aZfR2557oBsVKGCwh98I9AHnnh10ifOGgpFsiH9UIuyqDN5wW
uOcqAknoOaGAHu4q1iFn4x5oMACCzwaqdpuGAJEGIbWqq0wy3WToB+AepcMQU+Lh
Ut5DgZ9x9dejMEAAmd8DOmR+XOUi6afpQIdDl69nfmKygN0KbldkEZ7mpupixWU4
8wzvzA34fpy1UxjjRyj4TxmsDt5UtBtsdT6papxXaICX+EN8iF32duVZ+JxAGD6R
6uDRM/+NSaddqPbKgLxL7BhfQ1MM0me4wNtq2kL9ibsrd9AfsVt3/G33X/pCxEiE
V+5QNM0DocFpr0Qg5aQnTNPaRUEj4d1wGnjUrXeU3T0FN4plIxPAdVA46TfdfSLx
Xi77yD8llxOcTTqqaBebt0M6oVDqxnMyxnv2zIIk6W/pIferdfv3W4f1uEsk2BD8
I8vEiXhiXL5lz8vdZ1olJUPU+mRu/b2DPUkceX90eQqGZkwK1n4DdAm1koJzhkQl
W7K8FZE+RNMEJpUyhCUWlfghpKnd/WyzEClgzlVMBxBLZQy2a8uZ4O8BCkh+pg90
Qb5CjpdOkCJAxUNR128z4fVbO5A/a6EH8BcfRIuGrKswdvSL27iBg9X2pEHwUIAj
/HGH1E5SgJn4sxbSanjz/L+2s91ip19tPmHGjd4qEp1rLJ/ohtxer0rv/EsYdO00
mgUT2qzWjAuCyAPVRegU1w88veZYxq2/N/nM9vsd07jERImy4L8AiAIotcHaII91
yRb41BaYRjwqHVxqkOyvrX/rzjjQfuQKwOiM5RDWjLmZLWx4LjwJlhtzVNZDG2WJ
BV3cCMxnG7LhCUCCwipMmLY3X2TOl5nVFvHW5Vrr25ZHV/CKngMzzTVy2MEpIaRu
4QqXDkbslPUxGFKgo4pqHB1UO2QhkowBLRPG8zNwnUjvLEhIVDCP3EkXEVtDirHV
G7DHJ8jW0Xtf5hJET3hvmrcggJ2caIKhOYo8694csdI5cjERh4TpRwnsFtBWf+YK
e7ENQcHdBmxU+7RT/vRCdLi7ViqJ7d2+ygIDAW24k20FhC1KUsU60tf0tQcDpUME
70jgI+idyNIHcmQPjMPM4M4gI1qe4SUMiGXxGEtTR47A7eoiURGisbeC5kPrLSLR
/fvOJHSy9GFxQYv5bmnZpKASCoHa6nOmObkVDHuL/c1LPOM/cGa8q1siVMeGUtnH
hJs5mWlvtgUbuLsyPsySryudDJA0/poyhB/OhsideRbpexlTdFZ6O/QnoemRdqNs
1T5OuZ/eXRqsPVB51JXRnXEKe+hRGz6SHBaoHBegyuERAzkicskPlw5ABYJDOUpl
qxigfDIgW7iplG7cXgUM/QYTfGPmnVnUok5Y/kHIV0ABSAGya8AKoEGtM7TUytFh
4lHoNm8EgM8n1Te/lflFlBQocNWSRQFAcg9LnN2CG4K2IC6WHKZ58UKlT2W/zc1S
oiQAC11TJe32nrnhFeLDHncIJo5M7RPG9B6kH512LcDmvfl2KxuMI/V3DoJsxTYB
PrfNBMeFSb5AUaG4my0SAX1K9ZcxlsjyoWGE5MECYx2v/t3bE0aJhaI9B+uoZMHV
AqPJlB6GnfarVAcnrwus2kVNUsHkY4KMVHyoz94MxJmH4shmSLnYv2BRcm0yIGzZ
bk8/03DLd7c4lIhcYuF988FevZBOSL04X4mnDGw7gMhc/rwwh+kAFgQ/jOYvWl5o
2zCsw4K7PVPKGgtpsOpNgcadUDqtQO+fw20Ztad6UogrhpNFJ4NUbLx4+0VK9mSo
kr4FG8dUxDtXrPgrENI+N1zBH+baC+VPNKKuZu9l5zm3GeHVjSQHL1mRYYdTbycR
uN6kBTd1iBDD6pdDXapsysfOw7b5vQmb3HZuGUSGuJovptTYHeh28PN6Rd6YXGc7
UHP5m+p8LPZ74S6oAsjMvbh0s2ZL5cKhd5nPlkM34XwTTKGmu1CakgD7z09qb8Jd
i5eVlNqFxXOmIxz+FnJCR8Sb5ZO61UbiVn4D4jXWnT429IDT/aRMR/YS9Dy4tYXQ
jtI4UxdsYH1D9pkvTz+mKhqs2L7jVWD78YS31OGf1xIoWT9e/MNSPEMBnHKEOLbK
mdqfQRFVZ5z0+TUr1XQF4F1k8sIwZhHaZXiNElVxRt0UGbRAldESCk8cqqUf/sIt
lMv1m5ehMK5MDlTwwvh9ylA+Tz+oEJEi9Y16z03hVSKLrUqYxyQ+R30wtL/rZdRO
Ue1lhCD6Gn1ai9AhigwY/2oGifESfHLmISeEsbziWjA0nbuWp+wFZ8dBKtLpMLQQ
EQ6zfopgt2C5KVZ5BmWtvqrRcwQevYE2hBrHCECLqV2ArC+45HQeqBFQNjWojy06
Wm2HDk8obGo7NlrqBuF3h0stEv3tV5R58Y+tbEnaMKUqX3fAjeOMEp5eH8t060m6
fxR2tMYKHNJbwMt1+x+RA8ENUUDTtUIIkrTkb/a/dZ/VGXxWmYZXCgcdWKaGbN9g
n0BP2PMzxRRlux6CB+cKG61wfWCVwk+ol7l/IxCzh09i4Zn8jtbgU2kW5jEj+DAY
s6n6SfBL2oss9csE67Ab5sDQmCeIpEkUD5iXihRj5PiKUj60CbfK3288uxXoOxos
dW80wgKTbfXtSo4L4K8hc5WDwzAgSMsHcJCc05RHI9nTBwlf8jyHVMMwYJScSB25
elmaxcmMiHEdJ4sWT25kiyWSFgTe8wX+t3Yp0grmmAMnhBOFQGlpgQKgl4yOwZ+S
St05XojjiPHdP8zyQ/x2pEsfEe97CWqknONDL1QoYGe11+3rIrkh0tIFNp+hBFBF
ZpNEb2gS7KlLU/qOcdNS5aWUvaExQJ8Z4OOwRn1CcfoP9B3e9zNYu6Z5zIa3mktG
q3HaoHVfT6MjIJ0P4mxr1QvJPHYbn2ZDQrcIVp+wbOPXynBNS3U7N1+3XhlLw8jG
aXSfjlKVv+/ZoJfA+0rdEZ+QZ1GvlzPg6Z8IHJTEDXYZ5BN48Y+riAWPt+5eix4D
O+UydKpMY8+AXFeDZu82hSJIqn9V6eI7jSHFgaMMcTq4nUCR3MPoxJsEOMrnoirY
rj2b/FjSKAsYTg0TRmlk1jJlnHNfCFSU/yiELAwCH7BGUALuuE0FmmNhWpcQjwKv
MaiIdkHrFdQS0XdGdNPmvhN1Vx6Hr8COCbcDurkq7AJCnN+A2bhJbCe4MTJuxqqH
voYxEu9Hjn5082eKR34hQuFaAxKG4HsA+2T/M84uZWcJAK/VRMagsyugMzJVsncy
BwOUSxWb+kKHV0bZxU3nVZLGJXQzpypRrxF93Dr1jiVsovFHpIEifhS6iBq/j0jC
akCuh72RIqgRqBRKXDZ5bixBHrLCid0AH3BR2PKQGhdTUlMgw6husSBG2GhPTF7e
Cl2/d01ErWKrpsC/EoOLlCoe4mVTGyHChGeEr7MpYptw5eypBm+Ut6EIWM5SfGNg
mcAqReoRm6CFMftlaX5l/5je1cq+Tx+qQ5ebECcv1oJ+ud5O+zgjEoAX/+YB9BPi
hZPukRHsd8yRCB5vd08kSIkfXqfwyp7K0TrcruIhZvZsiFaQ2C0q8r90ewdFxfnk
fd2m5x9+NjyEa0h+gMQkEhrfM2Thf/5Xh+dDf74xHirpkx4yFyixrg6ZA5Pw15GF
QqsFOyvLqXbaP6CuO34nPwvziANN7L5M+L1Q1MykiLBMmjm3TkiNm7Hwlg4piD9W
wWG6WZdQ6Rp1iH9tIexfZk1gtVpgFNHte00MCyddP+Ilqa8GWQVRxpdYVqVJmXCa
0MtrVgM4CYVZ4KpkO5AMez0JuToeZai3yPm6CdnGhTkPmfGgwIYVB8W5hltL35O9
bDhWdjbV1eWp4F58835IvcOLv+8IFsMKVv/gfKLnX0kHzxqJunWmadrQryzz0Xjb
4B5HTLugqRqpjlr75Rw10ZMl9QO67diD1DeJkKuhPBlIsAJd6/TZDluze824GKs3
KjZUsO+OP4OSk7exwoMnNsL0NF0tcESEX+MDTVB26SIA9mC2nS4deyf7A4uNmFY9
6qLWIalx0WUn+KAtbQ3Ar7M0bS3eh2RcyXEws7KfMjRqB4IlPGMSyPl94BlAeAEW
oaPNb8vxt/xFHnc7x82S/XG3ZktuTyCJlq4Q5y1dXXD6nudhJLRUCJ1sjZphxMfX
IpKSjxsvHnUnc7IZ45kzNCVjCTukG8MgIrV/+HUhsQb6dKy/vIQQTXsAS9dEC8aX
gQM0HFVb9QOtDCnpnegieOwiN1M+tMyVNYzqwOPzOxPqQUiOqu4l8P0MF9zRI3Wn
1XPJ+4Lrz4yHBppart87o4z8KLWup+PQnN3iTCnqroYrQ5PMzcVUJ83YEeRJrXDq
0fP4FoBqvx39kwAtSnBSKkNap09ogfn1t+C0RRknp7NoaBOCALMDnMJ2re1ywf9o
e0CnP1t0kTFSjY/C+elg1XBcSkld+r1Ohj+V/4TWEADaJ37Bfma0aAUGGIWTlHsR
xMJJTyYpBUym4naqn7FF+Mbc4DMNGYip/0TjsiHC4s6cdjDvARJwgHzshFslADAM
sGnTZ9X4nMtW3dB7fqA6eRpPyXdljT2xg/4/sjlMNa0ZD/JeR9A934uyGPUF2FHu
fWZw4FwN9P4/clI/F0AR2uoMFan0Ww+Km2HSldWdyMtLM8LFyA9cj4v7VCp79efk
T8p/HoePytQAuRQobILlmJOvJmT3/GPlqWh9B8Y4Zhdg8HseSUNLDiy5q88cfjfG
bcEdOAfx96J3oVIEkH187l1PC3tVXbGvOnorH3g+3k//WylgY0/EfOKPHwkreq5X
BNyfNgprb7eZRfICtBwKmjHlA5inGaCIl+F9FJyh3GXxAJ+tCmcHzswKfeUj4lND
HKA3J0peB5HyHj5oVMgnz5iCyWw+W5QG4TmIwGtZY/3J3TpTY/d0tQFJTtolzJZ5
FXayORNjue3SG/vGD80ubJ+5po0YNrrIAViwdOGiVb/qMTok+0bPhG/R+8vJs21A
36y0ptOfEf+3b7W+7CVhSIKeXoAeHAFoI9RVllfK6AAAJLgBE9LE95QFq2bJk2O3
qNkuM0LzKj1FAtKkkYwA0PO95O34sKkmmPHtAi9rZd5qWkdN1BYuPgBEJS+5vaHG
uiTC4lryRiNUP4OoeaYX5814yQnDysyDeD/jacph5B30wM7nX9Rzfa6jNxp9uoQ1
/K/hTFlJQ1kQWzlrZgbxZMpvJWkiQ5lRGwiLC9YyZjEbPyWFDae6ZW6SPaxsTu9X
NxObdjIKKza6ndxDzeshsT2DsrTjl6uXCl/K2RpSapXycIsXn2RuYD1+hag+AmFE
s020Vrygw4dGO9BvZ4ylyQS85aFx3/aKah2Yx1IrkD1mdhQB699u6h5kWCfwiE2k
BrnfH1YCYz5dX8gKjDrt7cf5TMTqZwW36IA/kv6SknBUo1kxt+O8Y3NvTGqZcjtM
wSsckhv8YgPglPfp9qq9COhotkzZf/fIKQFaAjRwx9aV2VmPZgfzVRatmZMtzSAg
XXxdfFpdyN7HwZVMISS6NdrCkz20fJnaN9Q0XRRqjs7EkaAOikqlQTFjxToQLrKn
0XOsJlR2cofQtxI/GAgfgQPO32VS0NKBE5KWi0/ZdL+wrBFTeMNhAcD6sWL3Brdw
Oo645V1l8buID6mTfUHkJ9lfZ4CF6TgcCMNlsHqQWPDSHndmBcplZYMg3kQool/p
5JovN4SF++pZ1nXQ0/ymLAQHVxCAQe2KgHEvidfHW501fwGZ4FzWGjyGOMRAVIQw
88m3xneIilIwyaTbYiUJhLmoRr+ptm410DwDk8wp7Z5BZdyCJZGba73qRekNE3fa
hGcCTWXe5oQLEdBsOB2zeqvqRRLzYsgxzq/NvA8Fb+CSb6S7ZW5JOu/5unS0F5tH
qCRmt3ydIhPTWzA6NHDRkVxNm7ImISP0vVddqqv5jFMwRYZeUMuHGuqhA6dct/0s
tFNvBeEEFDQv5yxFfoGtqQ+yWEJFPC3s1ib74wz/tUzwls4N9LEmnHItS5RZtC/c
+RE3IWzI/7uZin9hWPHDJQDgy0n4fdih37+uEakzHE0ji6ZlsvijkpujJjXkO/9Z
wIS6pR4nIvjlFVFTvbqYkuvt7bhL3d6baDbrZacyVnXRvjmnCA5/ltcjHgg+Q+dP
Mewk/uzg2hSo5z2NreWHLVbqxNzqn34MijoCsnwH57SS+cXC2DkmrxaTxXrshgMK
3QHcKvxsqVzrKLJQZzmWgVSP+7mZvdNL2ABGHnLOEayvSiQ+nrbWjRUukL8nbck0
HJ2ESSl/Ez8EP+4HwCprQ7T7HoEDWhBYwueFVkBQ9YpBPLsn8RYVXMB2DP+qfgA8
UrcUwO6DVV8oHmbvCL1jGhEI/YJtKG9Ska/vYKLrn+eMwkn4r1KbXa1A3CaByhCw
t4KR8+Gb8Sxf/ODxt+NTU4P9+uDRUb24z/W3MTsOtW7ndp6I3Bxn73qUCyXdCats
z4y94OBO9CJR9Lj3zZ2wK4R8VXpopKRGevRypy2XTXJwg6A/yqXlPfNUl0D5Ca+W
ilCkHtYzquVd3bgNHbwEZjTQmNyhwwc431qyQ5ZP68d1axRUZj8bBXnJq7lWjpGS
ZRPy6+AGSwfUszI78w7pc8e9SvAdyvhNR70YJM/LugTjedxwYKb/i506FbzSP0OW
5TCKzAnPnAlXFnzJSNT9VQC/q2p07N9OBQh/Lci1y+SjDUw7ciXQGUvm1PEw222H
gKqKz/mobmXOS21oRvwOTaRc3MzTuP0U5PnqcBi+JoXDSXN67rsN6r0XimvlJTSF
rIhzx4DsE6V2WZFVqjSSGoIH+HuqFegR8JAhx/j1Y41XZasesMDcWNbPNTrZ4d2b
ftuFP+gnGX+0ViYV7/YDVXSMarfXr2ULhnSpB8ZAc0zmFpLpg3sQJVlzCXNZe9/t
/InRqeRcqybtdF40vQn4hr2IlU2fRtnHNZXAasPbqSGXjqpTPdbHhpFN6PJz62Ao
79yyJPFMwWx6HRzLFNOWEbsEPr6e4sBlk2I3LT8tQl/5mL3Za6saGeqQKTVvTNfu
wIUiAx+6waYEmOH9JenNx2+FCUqDnLdfzpcq/I/PJCBbDZ15txKT0cCb8wtvAVgl
5OPxa4rQlfOKj4i+vMUzzo1NvKb9lfT8lL5i5nO3kFqbWBo0PrrWOKzXBaHvKZo+
IyY2xuJEGSDxi63VnJqYZkXsK5QGLMrYWiKY9cQPiVNtW9pzHy74JxeQXO3KzuuJ
t/JV7Nu2zlvFuzlIsGjs4/ovcFqg76bktbALs7AdlSQMPzxPFKR4blhzvABZewRL
GZSVKx0enT5B9QYnA5azIvnh4zV0255aX08xPQVcDbduDxEWMb4ZuadqzaeUf//U
ok0PBVqYX3xc9fV1suRGoXK2JMLc/vPw3Dmo52YgXrHp9oK6YkafN7RLLVymrdIl
pCGW/NS8FBnSFBG2qKcuJgoWTrv/OI2aJUlxRk11dvGoskeUmYBsSWE/CD/WT0Lu
7zhqfN0JFTE62BIwzC8JsPj/hCSVBU4ibs/MpkzhJISKsIL+mUxsWs2RI92z5YCR
/v6tnFhpc2o+1re1xyNIcjp1LULogvQ5Fg3jJR6lXMTuxAaIISv/p2p572E7cyet
/QzSOXoFzISo2s03EFcD7hkTHB+4vtFVgBJmvDN4jPTHfHttDpHdFZChfd+b1QEH
ZMWJEwNGD2sHTJAzE2JYvnEYdfMQ/kJmRnRLjESmkBStehHHaYgSphrJ42P0ldeP
nIfbmHcMbWTScL5fyGTKCyuRn69UJnGKVW8X9RLO+AY7LkUQmq63GL7trxi29Qva
j2SnwnyCxqZvyyEnwiL14m3ZWPsRunHiPM5Nq3QbKrhqqWJjo8CLR4yjsZ5vj24h
RJ4I97jLDlcI8o+LRFNEQ3en/C8rtusj3zkOmSj+0UchxuXuMYCM2F2mZa5OZufA
l2IyBIrXvo5/M0aPJ5GxgIi9l/fTXPQY731sHtccmGtLCo3UWuN++9510S01uFnN
Gsbtg7ec661hjvC5rOtp7qKBWYwAWCDfJY/PICeeSLCxnXlI9AFQt0xRcx034qAO
Ibjy5VVfjItV7tpwXHIRzwQJJ+KuYSfInjknfqE45tw8qz1nERZt0XVmMTNyEDIX
1gb3gy78aSoixBnLKNJSy7CJk865JP/t/wZOohA5YqZu1o8Pdbnw8UQXgTWc6qMY
9EcXj4lI47g15BqbAOeNqCI2rY6APwOzwwU9LXmPxQyt50x8AvWHNch42RgjDH0x
5XY95ZB/BIpk8iAIvovnf+8uCxV5p1b9DilYcxht3LawpDBbsLWBAsy/xMoJ9RK5
dn5t13J/tYlJlYfXBqNjB4AXyCusJLLVYhZKvQPNruFmQfPG65rR/meLdJ70vTdX
z7c57MlUwDJvEybDqOBM4IMcHeLYonza25djZL4/5aBDXdhu0XG9U+WMkuGvGQsA
soE4dcYoYZcPB39+PqODA+/qw+0oTAiu3rNuc+zrxjt/xeCl6NBIbnY+YqmVkXqs
2vp40Zl6Xa8yK1pujQvR6DmakeIczgajqkxJJFrZMiGKfhdWzFrseRo96iKBNh2y
X3zszdX4wZjyey+DjNHaSZYqrd5jTNl/OF75Q7LqvGHiKsowmld9UKQN4J/lJdXK
aB7KoXwNfXhYMbSijROJWFdlyec7ZZj3qHu3+ho/dlfJw8qotWMhNpaaEQGuH3M7
4Q8fuHaDLmwurZ+PixzrZdlfFAepgN3bpWpN8vCfIE9M+1b9RQ1I/ISG1H6JmMgL
O4Mw83ioSQDFvfbja13kMGy+kCKeHLL56OfbrqJVNW3JQ8+DLJjmOOGSdr1N+UQy
99Uov+opXeaftk9J5vVdeceaBI0bTIepxTxX/R20mDrvY3sB47BXYclJudRu6pBm
JSr5/woVsFrkw/VmeE61UIuiH6zZgdbe8ZHcT9+y6wiqnBixUfhRSLM0sYM4EoXn
/Saye4iKFq7eUq1YADmWsh6C3gzkDVMFRzFp0e5MfKJaDY/DjDKyxTykLHbwVKMM
evBAHDwNd6m9Mvr9oTBmQi0y4W9jIKHS7hgxUPzPO0SOYt9LyNPdgQV0697sUfNX
yyabItu46BofPDJoMa/1lO/P2jJyfLAGpvS0+z8x+Jy8fTVpgndWrooFpF0s+kGM
9Y85OWyK6QfzSeFCBDk/DgwHkGtrmo/eM94nrBimK0QkFsKFOcB25hKYtAfCiu3r
uTVcBU0ANbP/4rXsZfKy1UmGfpo7xPxcRwj9np1EywltKBcNk99AROOtjrzLF41D
HvAZtMdqAWDa4jE3hCF7C6L7yv9MI2NzesytQWiLbAodwF/T0g6XbxKYm8ecS+oO
UzSYA90TjVJvDhvRWKkgjWDqgiJdAcSzGOoPdVLXpQLxpvpZBgzf5U5DIMZOqZ9q
B0TqjK1D8bwlcqpaBRtX+hC2gKy5u7Q8yrpGuv7ClsMb/d6Z8cdaw9XJ9vUWwIM4
YwJ+I3R8aAXWyGp13C8hSO4yRFU7xxPxcTMUzVeSC3df+MUorrAyj2TEXIohwF5I
MYCatw/KSN1kUbdLPC3CoTb5plq5e7nrMvs65loFBbQdVd2aelCuZ6tTHTnEUbAf
HX57dT7qZqIjCmZQaFn5At93P67xBp92+LtDEknu0XqGUH+NXJKP1vsJ/FzsgzdY
IWiFEWEOm3z25sABvTKc+LvFrXYQ58QMYlALXjrVyLVjGO7S3HGkWaC7m2YbsaU4
MWZMTM9mvUMdrmKXjEJE/BfneMFyWFuzH/6iPsG8bHbPLzvzGZM9pP04YQTHus/j
jTp8nbUpWvJCvw02F7OnPkaVm4k4A0QjblmtEHQziBN7JQPW3+aDH8AukFnLIrUu
27Nhhl0oLvNOwCVgkXsynxGfW2eofXNb/DSAt9T1W4zL8dBbVAqSTBoeRiTrLBXL
ezDWPgAsuOuJpq1ZebQFcU9B/nqgEJ5I3GxytsDYEUJ65OflfhqZ47ArOHOHbV4z
B4yCUdGuEdNgeMRVMSRfo60CGa4dcfFqB7Uc7AYAnvuzSH+wckLRp8d97bqhdhyE
oPAaGs7gIFenuDqf+IV8uMpD6quOKLc99jxXKB4SLxbt194M7vdPIQP+NUM6BK/G
ynaKzww1pBhgZKCnyhb1Fezee+nO2demSWbxFT7yJCrRjoTshIG35FCoavZnjaXC
67g9F0UlG2PR++VSXjrXToAXReg6X/pt/oWUo3hww/3cXhxCh8dG/ex5MWJoBDVB
AtIDMSzYZi8peSThQdKud4bPAHTIdo7inUCxXmmW/mNy0j5PeyYV30PVii2qSEm+
ZV3f11FXUsNaW758lEfQ+voNHhcoOUfR9V9ICORiaSHU44SVp61g7AUPC6Bx65Px
lCBbnLZcfiG4jtounGLRq2Xvhq25dZAi+Zp+CNIyssacblYnvsO65KJReeWv4WHK
UAfKW6GmTXH9b+Hxuf0RJmx7STucQmffuXpjJ2A2HFh8EqMxdYAbN+cTEfZc8ewe
ueWs12d4w2TUkPbSSi/SQ+dd7a9hWT74k3J3yDl7GQMfcTcjk5O2E7AwLIn943Yf
z0Ir3qJ1S8Adg9r9J2XUSHLVoEajZv+gEMkdIQHK9qPC0oAEMHlMCFFIbV/qm1vF
E3XRgJDesCohKRrBsdcu2ywm86v8EO45MhgIPr28+cGlLhJYzJgKj+ZekH066Bd9
TZx36lpetkjS1GKBfCHtvYtbIm9LFSsOEk0amupS0sA3qaK4X22lMcz1Jan72oV4
2UBV++9FD8FyN24p0l43G5orQW1KUZaep0qTGxgp3nrtQDc78GG0hShK7C+QtM2w
kBuPqPyKTwN/+hnGjYktm2p62bfo2omJ/8cziAIPvYuLbFB4NfHPwWG/7rXJ8sA8
vA8JTtzNRbLZ89NULxGlSjY1q4UOVTl2/bIjvlWxead1CCO0x6mxQLFNeWFI4OpA
NSDQ0s54FOA6uGcYkYP2ugnhbtSt6BjF/+bjUWHwGN9LzTuYKLmVRjKAXNFs+USW
RXn9HdQ9GZdOfnGmRzZ8beTS8Lad2iFOiA3OpIB1BR4W8UuEfG2/BwQRLw5sAM5y
rju6rHIrRqqTwbM7jWSXZNlK1GmqSIUxAImtde+bTnEEEw/nsKk5ZcOBlv5PmQlU
3QZWciQgDP/JiB6t2WRrJXRLtoH+fqF77FWiidAUva4jTMBEq5kbp7GojChQvO/Y
kssYqPcNqjNUTNfjjOpJUsaEOMaxGyQvzV7lrbCscxODmkEdO7Al4VKxXcrvvgzF
Et9wvrlmjcsARW5VxtjBEMDJj6wbW+qek/StC9WPmmsj7gOfqVtaA9CSWGxcwlsB
J0V20YC1ucDIrvVjaHj90hOoZgM2Potej+NZ171BHfJWlhyZBkIDTEbpnZiW4VhJ
lFM8bfACz+6g8nDNvNvlDXxORSdUcrQ89fUOpBzhmLqi6YEAGIkr7F0GL+7VLi7A
W/eMDg0TKK3KZDTBXy+gNTHF+B1u/RfD04V14Z8a4dyY+L9P1xJRXgMZT0ET+Hli
8UPmswkKE8mOOPG6+8Wmwzcq5dWLvqUgfpPr3NKNz3LXqDkYFdR1rcICjIaFDZdA
+nbB1AX+SBmGdRAsHUkTzCe4Ap/Oq04wYVTl6qwTEdoib41WxEP5Sthr2VQRHtJ5
eD9DX4vSvn5Dl2re9/5XeZjn05ZNk7IEaTM+l/KaIBGwyJGWecp/Rdbb63WR0/dZ
N5S/h0Rulq2iAUfqYkr/knHLZKfvNNiQAGPJhjo9fqaEMgoSepX21XlKq6ZXYruO
gwUr6ZyCsNBna8vwohv9a8XW/wF27+cIQty7eVBjulOSsGy/hyqLdB5s4DSE28/U
hWDtDND9QiEavOaeYrsx3SMRdmw87OKUK5Z/J+jHlV8Au2bAF46GtX66N1SRY+lW
B7bDZfzL1PC85KVt8LJDPnzC2HTTZ1aGO3GE/ATmNA+/9n2MSXprScEMHQxJmFSS
vGMI361+k0nTGPff9fvUrjOLDfbndj9iLO8K1BNbprPMuDEXU2rTQGVnPTbc/oiE
94hf64o+Glecb71adXf1qk38Qnw+2+Z4FIxfREl+mlIRHB0DG8DxIspz+qlFRFOq
fqX2+ME6KyfSNMDldN1yCDa6M9wT2GiAF2NVuDPB90xfIAlsjQwMGy3hWf6QxJwq
O1qcTYCPLDCZ1OcfQSBlDpNK+4+ai2jDQzZ3gSJPhD6wObAD7LKSX2j/8ietpJQB
Hab4Bs40SdmKz4Gnaczix8nNDbNDqZxNyXUSEC22r3qjoSyBGCkHh8lzmxKhibXA
SLmre2KG+bQ13vujq+pjK4Os8hDkY6apweNjNDDPt3DvlzAmnD23S7V/W95HWSLg
rVgMSmiRffiVBWz5FPSXxUGUcR1esvopIDypVuJzPtK4J7joCqCTnlH/9WSZeOzX
24DPzIqmHNWjEAvl+L8vd920Lbwl3wkE/VIMg/l0BiwbDLC1Im/yEuDeFdroub0j
831JJ6F36TGj/f83WBnHkX5OEfR5r6He+NDCpUgawZYtAIcFJU1fOTv/Wma55tNF
Z8ht8dmVsJV8EDraL8Qd9C1Yrd105GDeFeCwFUr0xZph+z4lxXWmdHKDf//vUqAT
AqS47EgTMfU5m7Em2zQZ6rr9Glb+PYF6gdasRrPu1oNMt5wjSnSGCTpYFe1BDXs/
bRu3IZ1MmYh2NG8LGVqVvXbj30l8iBN8EYPGC54vzadrW8zE3fTzHum5PewtlReB
fUovdLJLKRIcuUATpVxqdToAXo/0m62DgH84MpAiFZDCD9AjhnJ1rRmogNwsoRhr
6mqWDCuwXB2QBXSLsjP139yvH23xZs9o5gn0qqaK58+E9c9+u+fTPn4gLOqhz5v+
BvJWh6XYKmO2Q5OT+EJ6GjMOj0GKvN0kyw9VFlMmj2nuXu3Tmx129Mo0lXiMihEg
NZa0hK2dCBA3hayzpr9b0hTVQvcd3aXIttg8BnLmOpOuOzWpKd6Ub0a61pi5nSCK
aL/P0TuQUP4vFWpsrndFUBhLPQTmyKIkkMGyvFyad/Z0X+JuYVmU+hem+dzu+cOo
QzGHP1K0UH121wvLmNgN6vuhHG/xzJupitDsAmZ4aHblwIDvSADAkMN3YzwJgCgX
qjzsiUEJMiiND6qhhHUq+UVR1uQQ28KtoktpjEXg3CxqwJ2DIM/SxKFNsN2tlHRn
FkEH+J3pE2eB0g8x+nKJYYoeGXdvXsIdXHlVjFeSbhvYv6DPN/4T3rC2qmuAeuwM
pf05sufD1WAzAl+2KUGLdV6p430HoyzeqGA00OoUuLJX73y0thxgunRHJbeiRdwZ
5jO553GS49KLNT5jey66SzDhbI+77UmK9zhGIHP/243sqtYtAemQr4QSlUZQRpDc
ab9mDSZ0Z7Ya6jkA52gsoEI2ruMvq5eawJWBtXLReGUrvmhITmnrUci8AntgmgJX
HAiz2QKW4GoLBNY9QrcNv1jW20t7y492Hz49vZvDJcuPi7Tl2X1+xti8N4xyTj6J
X//Acvbc1wYYBJ3IlIR14NZQobGedMZQvmWdFqxH/hpgMJQiD264jG0Xi9hAhw20
lUFXqXRu+JSBICZ/NYoC2rtYyLBjnT9vasi1l/sn87vpv+2h4LtF7Xx4qyejYtSV
v7r4jod/RuAMgA2mrfZ6xBvMlJg1qdpN0T3NxpDcfZEYvlsr5ceHMiDfHkjFk/zs
ODy/FdEeDDEa6KBGQDpadmyb7u7PU4Ou/wSuo+zdHiKj5hsVoC+FNwYz9T9lhu0q
2BdLcwfAIKc3UjF1bsvxAwLauvosTVFccTE0tZmoevB0naCnMA/2CpHM3awectfl
SgGXfVNAdFhdlh60nZS52JKBdAkReHYEuIKio/20kdczbcIHEwYNp13jGbYPjxBz
kXF2WMSxEEmX7SeGF6qJSI3zocjIwFe0Rjzr2pK0fTqykDning3tmFG6kb1+v/bM
vTtjW2C2B9KPOqWKcrEhdKNd73OHfVGuLQVnFmO9YydNvnYHlSabuVpMqQFleGmW
MNOiYp3mYLcsiTeunReg6Y8wwIJXCh666jQUF6FtkEYDXKVqzI+nMa+yczDzaDkM
C/BHF5Sa8kYwkDYmiN9mlvswSG1Gqe4apYpaWsZm+leuO0KQMlh+GWNd5AY7+iWu
P5I967q+4sOChOqHv10NPdmmxLdtt0TsdAGW0TiM4xn8dHzs2TS4RYiSIYhHYB6V
rzaSrBrI6X8IiSVjqsc0zkYZP0gp7W1GUMp0Qcii6XQVN1UAfLfdBx1NLJIJmHAS
tFt0vqZUBxE7EbAo0doWCein45nGihsHSxosZoDj0rNj1gKXUaIbSXGg15/Fst/I
vqOYbkO84LIdiWv2Kyf7GvgZFkBvw/y2Be5lWVGDJMt3WcYf7LHVDDADriybh0jv
APGoq00+R+Zqr7oY2hbTfoj3Rf9h7ghzta2AGb1xQruK+IQuzVhklB87jScO77Ax
ASHwEvuR683v9g0Mdnh/MVnGu002nuytDgE7lbKAOeteDjoePwxyfn7qYZJOlQKS
WWEoDeLo2dww1fbpjyRWLp2oMYwSM/yPnSiOYczoPxwGsar+WCaBxl13igXvRxsr
nz8MX8BmEbM+l0JyzSg6kOAztlKwxHAsjmUwlr+l2whjRSj31WLhHrACLlJAtjQu
6M1lL7D2QERKgIe+Pi9lvEAMy9IKhYeKjNoK3EIbEQlS2Teb5NsXBafwrLGmSMJe
paNuiVZOI6TYRTlQhu/Z2OWrFIcd2zvHMqcZBDKeMZze+h9YVgMrDwP8A0j8Qai0
oruNpzkyYi2MsP4SUVBHzqVZshoDi2lRBS7nsJJPSekJTKc7lX8byA1w1JvLGvRd
OIv1FsWsW9pPXg2KoKulquhUBv09MQLRzZ/L/pRCedn7N5tpqw6g3olohljRBSox
Swm9lDfm9HkCwn5CcUPMtAeu1U5uV+M8WOfB7CtDucowZ9mJFG3p5K0pgKZKS53d
yugX8n+463bwZDM9ktJJmiQwzs9zY8kyNA/xuvNsVNeQxFBvl3rpm32PJKNI5adm
P6XspClJDJGuF0p6GiFmcPuswtzwSTopGXWRDcd+/7LqJJmIaDrbs3LGCc19tP0H
IaPWPYj+55RXaBcNw8HNT9WkiIwAKHd7TNWUbwqAKw3c9woedQnzc1ldmfy3tin6
z6zWHsMgWSHTN4KwRIBAw2p4uiOdivt+UVS14llVjjtguS6xuAKCgb43gJZN8BNI
Mm+B7qOBr5ifr3SUxmX+3hp+vVrR/sKAv5itZvCcXJqu0HoFHDiJyM2ncey2+36q
cyoO9Vc0aXJZUR2EF27f4RxP7rw+nidlQi+qpQlCsezrDliQaH7G/XAjhsRwX+pP
4CGnzTbFX1SgLjj7k+Sz/WZNrAoYiVPxsxwMAhDQpmBNp6dQV2O5MTgJ+DJpZXwv
/pCCbe+zYgBubdepFLQFvlBkDuxoFT90TaAV3pNSBOGqZTiURQMct+zb0WIAELqp
6ndsqvi8bujUAyfmjvcHkzzoNlvFJpDibh+2Rp9RsmSrrHDo9jNEdp9AlLNgw6bb
PcVlsi/zZg3P9pxKn6hHE9B4wQcbvAGHVB3u/5/Gn025PVliG/luwfm6tFHa7U3N
dVmODIZjHfLfewMv9bh3hhan/ViAT2ZXGEcXcxDcSj8ju/6azm/d/nT4V4xbaaJy
zKonQmzE5b/mJtXiNzpM2psYeMXHDKXM/Ydwbc1psIHKdF7yNi3SX5GyTge7vs/A
YA3vaOIcLYw9FxdxAdPiiyrtxOtaQerOmXY2Hn9M6keYHLVwD8FyMSNEp9U8e+sj
M6xRca3sIBJ5MY2w34ou17L5c5oIGZ/8OOfsAYKA9N3M+okRau8ejT/crYEr1uqz
dRjG2x7tJ26lTgmsdQwi+mRJUqcXODgKvobaqQqod9SnoD3lpxd7XwmMMkFOrIGv
d6xq3JyRxSS9aQeO2xywhWUz0PpMYHreKwZT7aneZKnwYBhCRWZh8KItzhLRV8cO
Q580/GHZZoXDRfZBgMc1fCkw29655ENo/gucX1xj1OepJojpGsiWUx9K3/axB8qk
oMowqwkjk3VIh4ji61IxYmxiuEULZzblzCsVolK0TiuGN4dBgWb24jbJiXw34QD3
DuEFTnEwaqkbs6ql9UXDkn2SX7MmdxXmuQwE31E8ri8OuNOrAEGNwsYVbwMifEye
3LbAWL8VZf8Nxz2+b/NtdgmGsr8tWM544nH8V2XiH2ZOTfTeU0oTZUzwRCfA77Mk
9p05gO3rRTOgVzT7dkgcX8MWXBBUOOCWFjMmLVko0qIpiLM32FQ0avjWmUJsc3zt
gHaEibQ9nRlS+ScYtw9SxE7+GgZJ3dZfDN9qtvuPKWEINpObK+ZG4hxEwE9hnBWF
1iU4SXeBlPJdsiT6CHlxzfzEMNoLux9t4ANs3EUMJmyzPZVcLVjmZyQFBgLIkA90
RtWl2ubcWQv6gcfjg7evNmZbvv4hrlpwnDn6HoOrYWeJRTSFLLl5PgGnWS9W4rk7
XR2AoNswCT6+cak0JkQ/ZDRIVGLSEfikXZfD0X8k8Rn9yyb41ySScNRYnwYvlVV3
0veYbWVkiAGEcEsNTYNZvmk0G/waJnZ3V47MRyin0Yn453m4LRm7vJwy13NNbIXG
6YPzqnR8TM6/5GdiwyLPyARnaf56WOdS3cm/rErMkMGeZbyTexrww5A8ZRLhIIDM
miaGsWaYdXJiXBUAubFhu/aoStJS6A9IWwmEt9oGn5H6FibQFlGfkjK88Ql7b0+a
jTTRPMohzeDq4nACumaeLbrDjKuJr2M1OVoea1pNO00jT8T8egS7mdsyje3bHCy4
oTHuJaSstW/9aSZBbcUaixnSiaaoyXmziGyhhfD+dJRfjU4/yX5gUxqpmyGx32te
6bbD2y5cE5kk17uge4RF5RqTBbLFLERevJ1vWM4oTVNLEPe64SF80jG9+UGRvlWV
C3UGeMmJItvl5ToyFiaGEEyX6voQHA7P9sjNdZX06va/klMlxiNUSrdmeA0VJm+3
w09VSw4vhMTw6ShK2bfEoIr2DEEu8w09CMel/FXHky0YRms5vGvUvQ/jC4v6E9C3
bYlvKbFtRs/NBLvBCQ4BeyE/EZROVvDhLfv2qiEHatmHdrX6vEQWLoVdxUP+Yvxx
b+zMJr9YaKCPdr0XCEdtarPcyYa+o5LerlJ6ZArMNOob0l3UnpgvwTzrTYY1176G
EnyLyDszTXD+BV9byBuS0JU6PSb8Hsa1+Msyx3rXGAZ7UtdgrXtlvAmCkxBr498b
bC7UPQTZ5GLfCoZr4RpIxSDEYb7k0/zJJPzKytCydj8+Ru9ydNIKZYsXZuqGtsE5
WAT8jy0y48HpBjYvRO4QEAAJZSSNnuWnUssr+dvW6QQA6sFyaeeBsfo81YaEAi5E
sOPIewm1yLaHcjtrOg/ZgBNH3SveKaP3g+HzkGUUHXvGof+2B9DRPq1cTZYc5Iha
x5fjDKAf6i6IUJ5yj4LLmL6KDL/nhWhdn6CZBoziU1R7godpeMnGvrCNOfqFQTzz
Dp99wyd0qyOTzMElqWVU2gJhhL/EYf/q7/YGkE8PRbKilO7xqKRl4rxieyTIXsnS
StWXWDZHnhMoyjpJAyWpcZQHJAgaT+7aQh7DO/fZM8KB4xCiOpWG1f9WiI4MjNcm
Um3c1mNM6J1uosJ8lb+xKO8xDtNIqfhJncgr20RybltfbEHLGuaUKVeNpL040/n8
AbG8+ffntVcmh4+km6KCvWsJswiLBKUcwcXWVsfZtL/5Oo+owdTpx3gCbB2oYo0Z
xz/xWlX2t+4xnva6zFFbRpTGWXeLGOieYv/DJGF7dFrJ39/tQmBgZx43mLSpCrGC
/nycxO9fvLwM2S5QI1sIGRdwW2mn2G68PNpysWDxpVUhjim+HqhWcS9h9d5xGKD6
wP+6jpMONGczXF6l7zPjR1v2Ikl6LgDr8pTE4no/jWChkd3kjmArZ6yXTPVJjdjV
JfFMIBrbMmd8CE6iESX6fnyXF7/xfBGv0ZZN3UlKjMXQU7YyYN5VMRxClidGVson
NhRRycs7xV0NjwyMTjeTJt+ShHDZxQt82JLVwe762txKuVX9KPggDqCw/Y+rmfdl
Oaik9M8HnJRgTNn3sPPVJTyAR1E1tRZVZr9aedDmS6fQJ4muHAbB0E7mB1jWI0Gw
DY7FYSvBdPLw2r9mxqjVT69NAvnTx1LMO3rcuIuCh6cORATAul7IanxZ/uOLkA1U
IyDKQScw3GchPT/8o7UJCIJkC7/4yrteBq7gYAA+bm2JghWoA0HTKIkoW2P7aFhq
GnldkEwq1l4Pv+dTqpQhnaDTWLATAhd1yaAZht1Q9RqEqPVgZ/imH9Fwv71HB5g1
HbmVkwc+Ru71sh3XLQAfUyj4Z29AzzruCz2nSCZ8+FH0xYz/V/ALB5YKNTlScNsL
SHpa8iAjFzFp8k8/iZ8O9sW6BM8btW8QnzkJir34xbsIYe/+OsH0ZNNpG+EQAAwt
cmNXHlb3BYtkKN3Ehq2nIvSpTHOj8VDTJY0e+6WW9C/GEbykimTJ+DjbAscGVjDA
6WkC8gjS6cwmv4+lsmeZ1c+/oO3+FtqlLw1F7K3Y6TOXY8xOU6c+mG0+8HL2N5O+
HcFPSV0HEAO4goZywH1yMln/MiNAQ7/fYShIIUCey7bE2DTeqkHjGa3BRK4Y8npM
N4G4YxgwUYpRC4z2kJBuZrMVvqhsJyh0SviDX4y0e5zuHtaNaQr9FDby8MHIYBj0
n8bsjdC9XWqQex1ludsVitydgf+/1pkmB/8JzWhS65XbJqSGJ/ssFDKPJ5jxLwCh
nU8NBAuJH5pZobsQv5O4Mh4Z+vkpU6loPDsAmCBIJbhLmUTOuV7OYLfisjglrYie
Ef16I3MCUS0c2MX7A8FJy++tFED4/EhvTpiqHkYgFN/nHvFxMQf6Fav0Nvn6iGlY
40n45gtcfpcPo5JCb0NBMbfF7M0SEdJ/CVQPDWWrQ7D96B70V69ai4m1aiZRZej6
1Rg7Yy9pvM8KBsH9F6CINpJuG1rp6Xng3sBmvPYq5EUG/l9d0xhFiZBFkzwg6uCa
94JJP1Hsi/bJWEDJphGCbYKKPOacv3FR+h3zAfc7+SjILdsCgfgrzSZ42UouXg20
iArw3O74KB6EtrXCwxuxhdJclGz0efzz2NTrD1mvxLn3zwX2vsokgsD78xeZIj57
xOG3EwbJOYGHPex/DxK9Nt0UvbOMhbN5WreobiU4abmkg44u2/j4kVOWiS4gkczJ
23TQLpHt6S4pnRMKBakqNKHtlpFxVqzf47LZw2jrFIgAHwEXiKjpSh0VSoeHBXif
WqLK+cGLLYOo6XM2KNuYhUZRRD+dryZRJlel+LViB5F+XY8QdV5Bo5MgWuEuBpNw
yDXBcMjPasvEpW/VRIzm8KNj+JhqvuESipGPq+Z6LR+i1yDG9QIl7L//tZ7PT8nP
nbo+82KksZL0GYaX5PymxINQXyKxks6qcujh5GHH6wFm6BZRfGep4H2Jac8aYvo8
GkP6n8HkI9pLOBhze1HjBpyW7jIm0DMO9p/FhtlrV5AAsm++/o149srUDGt5WQJs
uNqqzF//txkOqCyJDyIZ8VuvNiSyFUBuenPOdW/YacQLNWnIzJuIhQjAAB6pmb78
mHeOEWEYFPD1vDEY+RIpsxbMmiRq1LlAlpoaba8XcH59H9/35jddvslI6Y31kzsL
JQv0qOmdlqMeU5+Kab7UnZTXUXucpjiZ58/wZLlqaMJqUFx1tsiRPlg+ya6oEhZi
aR+mqhzUb7tZ5LUdaADsqDCZYS0TK+PH+85IOggctHDzft3AxcY0badYqgAjqmTb
cc/J0wb6N4ufPcBuDo63PLowpQVPpDUTuagEfExYwjwcU2Hf3besfUaYIBD94txI
gy3X24HcBCsVvit0sFGvlrYaITtnpg+YMFX/hIiFu3lFz1hqRPkLmFT/G7/MZgy4
cQO8jFOWZjxuMEyJ/YvuuX9K4Thpz31kWpDC4qp2q30qhGJdINq+DlSeOfbhZjeI
Ps0njJ3l3yw4oahVLhqPMDwWe8QVQgCKcgdj8w0POYEM/avWnidLuXxAWxfNDsYp
Mp82NnMNgVGvPvJ+qo4iFhQ076+wYpOVVFj1pMbfQb4Qn/Clz1YVJq14eHq8ObtO
P9EJzkabNsKFjkPQW6psaihEXyHUCxSvCAMqTvtj0zzLsyJTOOOOuEvEzt/z+t24
KJa5Hqru/d7lhNxvvf7bQ5V1MbAM9nMaNQbbihHqljB2kof2s6XbK+P5XpbTPo0c
634HbjtvpvETkdPAvI/we/aTWEHn1W0fuw4THMBVrUnWb840Akml6t9Tc0sEYPmf
ly2ZVEsCqZ8SVno8jN4yInPcqD5tzVjpel30PbNxqKvMELEURi/me8sNMGHOYBE1
/N4wlGYPdSvxqSx9Cb011UVXtaq0t0R1hmETlahgA6IwlD21EOtlBc1CGrcSJBK9
aHRkVCIJjNGzjjcp/0NJqZpB12zi2E6+BsuHjGBw7sEZZFgewrLSP/H6cuErDkVZ
Vehn1fgV5i0fPye62XZIewx5jV1MsUWKkYdysrvZOEQHfYqkEyr3Cf/zF4alHQSl
3dxQGxDiDUY8ywQYc6JbgeOTEYtD/CTpvfNKssAtIlsL09PpcCyMvn6GEwncYEcn
jDdELhfZFJabmqtLXakrwGpRyMqiofSmjpa7S48UNEyJ6ZwAU0mc3sEgjMiVcSn3
SsC2bSYlI5OHm+tP/Jd61GcevnWabtapm5qTOkYD//PsxEyQ8CM9mM90FajURWGE
lMw3S4DmV0XnP731x55PF8mZ4LtF6T4eNOQGKVbdzyYgBPdLJ7yv9k/ZnuXgW22z
fxqIUk3nYs6BhXwgFFq3OYhsdds08BkrhHbwh5Lw/DfgCkXB3atNMpbneRxqP698
/DJKBI/xZUobCfkp+tchwnvwIF4GBSpAQo+k03hMAjXYmzOkT/wGrNUka8RUWHNn
VxrQWzFoZkuO5FTVz57IRkfpdiA93uUat6BItDNvJLhlALaByWFxDeEu8XyweWY3
BBeIapMqaXH7tiCUg7ZGX3/24ZGi86e6CHGYeHl2jWNM55XPTQGZm8+P0UespxLp
84ANZQXt1fBHJBrNG+Hs4A6imGb6fJuOrN1MloXi599ViOJpO/6XVf1RPWbEDTYH
8a9OOw70HqFXpXoZDNpM4NldhuPzBaLlEsKepdpUXFq/vCHQMCLKdTWHNZNhyJ2+
DaDnR3eFi58uayJDJGDVmfKW61agSn17yuU7vp6UWeVVN+svQWyFIsC4jOZ9c5LI
XPi89y23IMWMuGDSiwMTIhQYW9AFTm28Pv38VvqF6ANlEnQlEukG6gFHF7RcttFV
epWOHh1jvtf6VN6zKKEWq/Xr7aZi6tnB0qHaFHPK4Dr8WIK3yIKDJk3k8PFDLWMW
1+HDDf4ezBqqjC8a0e5cg2vVRWcEyGA1pXpDwRX76vfcZQJNmA96586Y9SBPicCf
bWJ+4VP0aeU/x9uR8gpBC82actrnOJrFyHCz+K8dt9Q/lT2RXMzouA0dki8CmpYL
M/VR4A4xxOxt+tSnT4n6C344+j8jkiuqku7JosLQMVq0jLV181Sp+IEYsAOfhBav
yM7kX76dK8E82ZmuiclIkqv5EQ7PM3hVryzPhAv6wQYTdF42FnrCDPWjhqLylk+I
jR0iB1cSXo9oK2IOBHC+QKFhdKwfkI93+b96io8S2fYWDCZ0nl/8pQjS2wr86T9k
xjXyJ2fYCEbWtat0vzTBEbcbgY4I6LuyfxrLscouDyHFDqT7mAB0xA0or8Z1gaZG
H+P/3YY1c9/YDvbopwQleDFK3nubf7HifXrli5cP8pn+gJ8ZdHTHWFP+3K7QJ3yf
ChSE+LMbtRk196fHMAsUoJcRBEl4PbSwYaf/5JIfHJfT6USxO2fe08cTheIW1+T+
L42IOvsblePzkWDtyAEQdaiO3dKzCTcn+UAi0Ceghd3dlF8R2FYPg7o8fwTPkVBi
ZCx9vv8OsOoogIzEAzf4QMpPDOfRlykR9xNNsgpgbKiM+ZFjBiJoQ+xbXCQXmbN/
Idg3a9UP6RM+qR/U0RLGuwrSbwg2emDDKuX+igakXO8p2JEzq6fHg8dRpFcfAbOn
fP4oV4KKUCj7Z7sbVsuSh9713vn9Qkd+yEOsRQ0tXTzznFwdIUWYQzEYzcsl74qM
/Lr4bU0Z800CKO6A0dPB8KivzDMbt8mC2COtX1DfCG4+1GZHgQ8pfAmjq3+WluFQ
S0lODsywFCreNm9K7AXbkzYEcUNABSIG2TMoJZUuTNtBABwIpQU9NW5EKcGiQheL
N2U8m6tcXYD9j2cGBM3HBSee8UAS36uTdsfwYE2htXLXpOuVK4TmvjJlsYihsN+L
50y5JhxIwiMCKvPLpzttX2RE7A+EzAOTCxl2uTPnHnDCbHgjCjqMTxsLhdjbm6JM
qtCXUjL3XyO7H2VDwCcwWB0aU3bGQNE/hTOt2LRVGCHlEGEde8xnAxymq46beyH3
fkKOpXcDcfy2G2dI07E24BidUmLuMWo4lzanjRrUGDi8wXkcdfuKzzhkOTdod+fC
AwzliqtzoptT4VmBf3meFYzabGRkJuCrTzpXkzP2QqT+iheyBheP+5k2xYH3fGCq
suTY9igB8gnQ4w4XMPUeSFIk6Mj1QpJOG2DLkO8MQlxLcrjAhXVaGX+iD6/BnkPc
oDHPtSdsCYRQNLINpIO7gtksKRHL5o3UNl5cSTnGrxjsFvfMCY/grbdpZ+1Vf1v0
kgq/amIWlArg4IB83zeCbvlowYIkEAJBfEXA8iz8keECUgyHv+v5vl4fXx4C8k5N
amKVdMNAyXioW52vweuDHyYmWSaYAJQ3kErMt1q1coPL4tCeJj1OpO/wIklHBA4n
YiZqkV4ySA9Yqsu14322Ot3pmVvi42LD81xrjFReVnaiKMb1UzjS/TLC12Aqntj/
hM5CbYnFv0QcKj2UVT36bjugWKTZyr0J5Ga2Vi9fL1J81MOO1/vXh3DEwUuyTQNR
o7Wfqrx5S2J536fbg4HwK5J/T7kCOkjJmj+1K2YjGonkH8ExHnBZ0gC1Vqsl2AyV
tNMoNrG6Inlin1m7X7O1M6Tk+dPWYegsubIDkrhbAtBXYm28tu4cqHE4Z/Rgb3Ql
ieit8ErkFkRlwqGhdcqm9YY9vYA5Zlf50Jrrv3OcibtxH8UDriK+7bITqIOHJOZy
fu0j5JcKoXZLwZzzy/MfqqqbxoGOaBvu9AaBarsmf2yas7W3K6EA94QhPD0uxBLp
5Ol0W3lgjd8JKKgp/BBjvuE+IEvab/NsvJtmyL3i2X/3lEBz+ZzP80ki2IFLkTll
6utde9GTgzkjQBISiLGkkpd+NZ6iVbAjh65Z3Yz2zvyp0IlxzUOKwp+jzUdSSLsZ
lJfzPYGoyfoR0ePZoebEWux5DClT1C1x27reoL0C6KOG32j2Z808D7AJG6SpHK5X
F5xag7wyEF5mb/8ZGfMKNoWDmNX1+BfsgIdoc0KpqzGUkIICGpc+JfDe+3RLXUmR
Pc8x5IW+8QGoPUD9xGQ5B1fsFmpHh45OAhs91ggqM9UXBjfZwgpHdzxu2b3Wcy7f
zPR0cmMiKchry8YSl8YFhHgHuYX3rwYcu9GC9lF3MWNVK2pf+hgKd6Tz0envtZqj
ZnpWQIQQzUxzFfBX0rjEMCBKSdDkn1NGkV6l37kL+KcR5pxu8hckCTg+JeJpESkS
2LcQAZx5l/AvhxZ14IfkkGnmPG1+a82DHZ7Z7QDzcigt5O3XlbRhLAGLIPA0DyNf
WBAnG4LhaGEx/OYGTDtf/pQGS4XgQiOq9P3P2w3zGmeI36lmTlsljD9SCj4fm/Dx
m8HOSY1h8eC3btrbVHvbxXdPR43ucK1jPdBkqArLkropRmR7JD5XoPkCYqV8BGay
S4eFB98/iLy7Xzr2vhMngCoPvEnv0dVFs1XLgaCAyFu6c3Wo6iUPfXsOHPoZ/2J1
w1PZVoO5biPps22nO27ZBEmpyImPiTm0VNtINUNrqmnqQOshZEsXpRqg7ICeQDhj
ga/+JC6OqgUy7fN8AiD76WJezCxdXvuyGBjfrEVgySjfEIHc0CBxXEhI2EP6b6fX
9b6arLbRDGBFwadW1xzBr/Pnqgv5Y75kdeIvx9CoM7A7jm3h9Rwk5iJ44bkTb3up
mIdwmF94f4NptgeP4QrY/UEJgsKJ19ahaxjp2SjC7yqEMBPvpxuzEgdSgYxOV1V9
OzsZSNQYDqo3A5BnnB15BRfot4HmHrMFBBS1iKOrcow8dBPXc2JaXSlpfUvKtZvO
xfvihugHVKVi6NJDtiWEnZBDTbwmH/nDy08kCyl3fZN1oBalZzNN8TYmpOzWyLgk
hfhY13gCVI5luiWZEoN5q5nOc/PWWxPcyNTMQpalUnXG2mXZpKiOCLWO7Cyqgh3J
727etsUJJvzYUCvlPj5PMts5yjpmVE32KegAgxkQKzxyH42OFOMU6e3PxcF2K3zR
CleJ9XKcm26AKmNFs9HiI5IHgPrn+TTvKazqxQ/ialWj3r1J8HAO/xRRdVUvPOxa
uUM6XHc7wWQ+/63KF6cnGV2HpLKsD4IIIQQFtFLebdd2FO/ekQpFSw8mVyBigXNl
/LguY+nIpOmqsclSv1x/SEeIo2RINogSFosz+Zy4vNkoPmno/9r4azKO7K9iCCpU
NqGTQC/aU+X2Sy0zmFdy/IXD5XTYhmWQLucm/L89I6QNkVojN2T1UrSySoPCAjnB
brFQXMUR0rhlcUYauQDVpZkLfJc01eDMmaqyIgKXRe/EpYJPAgGd1BWChedtSp3x
oNZp7of7CGuPpI8XDXWXWWx2BG8QBROvCEt73TaBsa8/64fkdkipxbK2Tu5tTsv8
i0mhHuNvuFkIgujmU7B+EeIMAdjDjyEe2CZ52Ap97skXE0BGuJEO8Skocq1woOv3
+tNPE4gtlgxpggKgMBGPEt56ugAIqYKjuUENogxlrBhJEbP5zyKzwlDxktSLt/yd
rzpcsoVaNwpyyWLKox1SDIK5CAdfPFyTl6CtzsWrnosCg1yB/eWAURTIZzbkxLJk
zwILEk7ZRy357X05ZaGoskUBFK1XXPkgF6vCruNhPVWJLSBcgZmIZ7jK+8GWLVj1
K9ispOXif1F5uZhVIe1V2dC/ATuNVL8LkWOKcUhrKxw9VvyTGjLfy/jMCSwNZj05
Udq/dlo5L2agcuL01NmvIgcibFXcGyXsLYQf4QrpqPq/wyPylFKkC6uQuU8HRZ+0
1LGiUTMgCCxSU7lWIMe3v4Wjdc82Kh2P1okpRydvr0tkKTFM5shdG30C7AfH7aXG
eixoR2beCgfGRu+P4L6mFkBOEUI09Xun2mqhVLB761UiMX9oVVbuFFkX4ZtF+NIk
iD7DTP/t65LtuWsAnMDtKObUBOpmgWBSKajUa5iyhHOR36TJAAn5FazAU3Roce2x
cSvIlRixJrXw3ZQ0HhyEnBUVY4qYDFcWbCMAR01RCDPiEVhyZxir5TuP1rIBJmIT
TW0qUxaGI6lZFbuZKYtFmyoZJ3xWRgBzRYSO+TInUbfJ4dIG3cxLArHG+X5ebHOP
PBlwJgA3GrAgfJEenHuF7rhcTdsMOLbSdQ9WYu6dZZKt0yBMQ34+nK2eK65K8tt6
llC53givhXZUXf1aYLc/CQmEaUSrAau2HypawCctTQj78I39Tn0Hw9SeGg2VVV/7
5kevK/2y6kD8q2j7XqGogOPBlXG8a6dKJ9mE2P0MyDWmWK4V3Z5GgNuA9+lAdsmP
oTrAlkJWFKe47uVdjeTEjgfUn+FYb1ycJ9OpyEN3YIVwIHKX8PTDoLidXW5OH1jS
fQ6nP/f2E+IDWasxz7+U2P24abO5wJpt3WdZ+GWqe78PEX235yqGbNpJhGpG+5P0
OPpw+cxxUaucp6x+HpnRxQD14aQXdcWqmNzYKd+L7/ONZsRUpcmB507xlHsQdMCm
LkjsBD1h/b+CyBf7XnInnehaQYXEWIPBMUJ3v73QYnidTSxDyDHmO2rOlXEI+lUN
qj7TjhGqUFe05aVS4ckDmqbq+Sc4519aLgHZL+nPAK+juqzbRt0xDzXWvCYBlFB/
MdpzFSEmMACMFZ/PP1PSGgbOp2Te5ty5VFBSzvbS40SbWRKRL2GBWDSlWqwLdiqW
65Bi0Ql4+vVG9jHvU6wnCRjUIif0FCavc9MAU9i4kDA3DBCZMMzBm8ftXJUcYFrq
X/lJYt+JAwbmu18Jk50PXZTOKbNK+Y94pLTXoAv8sRUJe+2+QUbqOf3gi532lTLF
HxxLRtTiFLiSPJH8ZE1vmI6RVYJD3WNP760SlCUl89LzKt+KLMNxgh9iB0Zz42Tb
8YFSxVMq1TopU5mrQLAC3Q372yezBmzE1PcVjVlj0X5F+GUqMGl9Hkwfsg02FbgB
NINe+UzcsN1P4Dts13B+HcRYhuiS2ata0PKCOQhiuuOYi4TZDbW88+IqS7mDZUg5
hLpxbYwoKFwzPyYwi7xmnJwoFkbWVYfo7r9BibH8bY0pKlFSeJr2mZL+9mU1PQ2r
XjtZw384PWreCxvUnxxrKoy1Ej8+9V8O5zGhtbU6O5xkzZXbkYbRMcshfPtusiX3
NsXOrccIwPyK/tSTXRTnKrKuIJKh1OJGnazF9hZWa7IMnBv8cbxIoLmyOa6N1A/3
ZhlDAGOoNVl7xI3n9ft0sAYwDdRJdkcoJozENyxBl0MJbOs5eXpxEkRy93kwfdd6
jr9yhweVHWNmp6Z4A4+nxPX/weJzSWG4orWsLFgVUE2RjupyAKn7w5FgUTmYIhmV
4ZJ8rJyFRpS7pY8YH5b8WILAjQa4b613plEx1ifDXRQY/X69f0fZE4qE0jUmgEgl
AmIRgoL/NJn4zo5gTfRmr988Z4rQmuSPzU+n2fbU+4Rs1OCha57l5xf5ARFJC5MK
uiRLMkwWbSHjqQO+9EhL3rw0Oj+JrbBH3fgvH06ZmZvL6f/URnqPJEIeqsR09VKw
hAOpdAxp78LuSwLggpQzalJTTOOabLWmjRp+zC+AF5g8J2jtQngQm78bOU2xTT/j
RWH5FxLEDjNDHAbhnB4npk531MoBpLIy/XWrqOPeslE3YCNI+9Ijg7X03SqsDhtt
gWdiz8/tKH5z7ANWcfydzJAVzViVtdqPuwCNmnRAMODEeJuedtl+u3wmZzuWyOL3
w0D3wvuzsyt7RLhp7ZfK2YtIODG3JJWX0gpzqPsThuoFmv/WA51LoiXXoFgixmpL
W9WETK8l/eYTde628t46SVoptnW7W18XA7xIrtFYwMi5hGVNz85JsyT2IDEW5Zac
p+AQTuJ5cjGzl/5hmNaGPiAN3xq1Ai5leZDpqgRV0AUZnXYR5dFTZQCqc1S7qVaH
otoDg/QvFHlYxu8KvRKIOPkzOfMRwnqSWoXv7Hs1Wnb7ymhD+yaNcI083SBYa1Oe
3uF/Ws4a4phR8dnSJ/KHVx3hSwvdSWZJ92QieXdmTseMOzYTbsnVDhEHf7E22KHh
8CZTSbSPKI+321b0tZwRXPexRi7KCRsi5s2iWkuM8WjrGh6epkzxR/jqyk79SUA+
70iQRArpaf5Qf5rhE+Pj+RAUOtZd58WMPsbafHcgyKAPTOIRJyaYzW3zPA7SbfGJ
+MmjPE5X2Glqy3YVRMMc9iUiwMXrkk40uFlC3RaRrsbfap9pR5acW8VGuJrzN9i2
jQ2SA7QlfxIoOxtrJVddESm5Zo3Ihfz5mbAsFp6Ay4KbxNK4LGqRHeNTcSXJnMGL
ekp9r1zUxlpoYJ1bcevHoIfmDPwFJHoLViNMIUKirNq4Vtwd/1eSwNAgmpmMpDT+
m6S+2tHLVSRJ6mjBpEA1zUpQWCnrDY8ycjwdDNklyLBIVgCcx7cv0UHctt4hQuzb
Tm/AzV1bDaiWHUZeVa+j/d14kenaPoKp3nyM27ji4dzePYSaI4BFF28IjgcDjpIO
aqdm89ga+4mIicTN3a0ioYCQlAlPjcWqgBQRhk7Un5YYkvRb+VMwH0sJ5sX5iY8b
zny4+AVhJXSV4lcrAGX+P8dFoXJPRE2YsXWKnA/9jfD9h1A82XCQQ9E8r6JNq6AI
qp3nxDYY3EY2I9uuiGANO1wsWllaVWC3XOVdaoDfqtKYuENO4do0Zr5PN6aTNYaF
rNjswxIAJlr4aXN4C9vVgCaxnKZlJ2tQEsDZpRC5xoHb14W81lb/NPDShDrxaBKO
qy8+XSx5xn3cML2bRHs71hN84VeuGG5uI8lgsHN/QRb+41kBbum5d7SOzGbZJxR4
xtkxl59N0kuZXzzdN9u6PKSCyL2aioQ9gwxL2EIfTYT5dIRvUeYJSN8FXs5rehj0
i9tk2IqVsgArPDa2LehGaOeGbCcXXgWB1S6ZjO9OlZCdSVJJ1jLNdZJQBC+fzGiY
+VU9xO7eg5cc0BtBLMqrmtcoQLDn3gXMyzQBN5Ptvl29zEW45pWTS8CoFZhHFCwv
BAtSn/XEJr4Webvi9ba3wVxfqSk/qpMa6suy+frdJ3gPTm4mYRliG9x8TIRE2pSC
c783pKv8FRwbPcdWYGNfupL+N0DgIeMAkizbcEm7WJcP7igKu7n0AMNvhyAz810T
Z88jfHJs0KfPov9xJMO05xvVxK/WCLp6LN5BtJWwu2t+5Oyk1B9SKGsvfk5gXq8Y
f7s1GQR+BdvuIcmHn7WT0mvRcviF2L7k/o+XfMARov2zf/FOKRdgE2uHqQyeJTEZ
9gQGTsuUddd8V5lyY8iCnKg/EpqM2BWKLXB6MS6CL+OQTPwPhqf9TTmXZITbSyVt
Q+m+wctC6hZeXeEVnYCIAAGpGJiGOvzuJE3Vdf6U3sgKe7ftg4Xu7OpYAfKXygs9
qZcCfQ5hdoQkclfLixWVTGz+L8PN+z/x62aw6dlxLuXhd6LOLjpw/4dZF80lXdmc
8mCNXA0xUtKpSISnAuLPs2zN7ys8mpuja0/8Pd6fG3kWeiv+Duv/R9BD/zdHgZaT
57LXeVf4RO4YeNezpzq1BnW60IizoqWa4x3j5NZCowr24F1tqzCLnRxtGmOAVah8
vaLHbM5TruqPZ4i5y/sWLWQ8RSDMT0v0VSvLOOAnSZwa4p4eJvy0G5H/1XECumPw
YtxNfwq+o5G9U4otLAeFOI5lOzoIe3hxz1aINMDCCIb89q+hHQRlC1HDa8QEjbPv
0LiuBIdMyNHIrGau7YMo11UUNyogJQLVEiQ0FPsC8XKbpdVNIXU8TjMe4gsrPeAV
fxMDmpLtbCRUhKySfRBP4xmjk4wwBRQ2s6OW84VKO5dx+xZ7FohZdYGRagS1sA8k
juzKM+XiwT7sTD/CP7Mqi+fRVPdGTEABGMP8amrBzPANLEjfM3BKFjnOS0lHO3ET
myzycxut4Ma2zXfdWMfhZWf0x4R/8LXE7uqRUR+J9QavH4+vPMRYfUZ7GxOu6Osq
cND66/tfIObLITOmaYW6F8hzwFw3IfeASMKdQSWkWfU/bNcdxl3zyVV5vSgyEmxQ
iI4u6sdak6yI2aUckQjT2TlVSLWKKgXBGAT4gBC8nCxPfbbqdUcL35coZHMaTAGK
pHEV4BtWCtKIGPQRn+8DHoOi0HhwG2Euk3/hYeFVL6B1YTySQsd+3mvqEUG3CYTO
xGdldlLr7miIO1U0EIkHM7G22HIODdo5FPEOQSdFgujb1RGJWW0GflkIKZP/Hjm0
mJ8MBnouxb036+BnUu2O8O1lmfsLaZbHjBfPWWM7OSxiLDS1wyUPxAt6UQlKsLhf
aM7nH7wchYIpAqfpQuKNhN6UBKJX9kc1rp35WbdYLvvWszjTEUOdOA0PTSZj7L+T
yyPZKJFDENQQnRiV5iFJmJp7S5clCCsvZFsvEdLvLRP8TP8BWjiqx11Lm8jAISau
Vh7LZDhKk6Fr2gNs9GgEM4XguXRUbFrcCdIWrtHU0+qcAwKD3fCKU2mAvk41eyXg
s7rewkp4GaFBpfLAUPw+iwx/baNrFOa1gohox1rGA63Jj7QMhm7B2lHgWkUzBSXt
JsnRN3OMG9MhK9sP7vk0kmoolffSPKdW2RivlCSCCqUwIiMMyAwZ6frolzw6brG0
DB2StpvsWrEV8Aji7C0Bamwtsjk3BtDNDsfHrma7bhWploVXxjN6gIEtp3FnDi3c
r5Fh4+5DMsPXpS3Sus//uCevFUYM63NPjhiueTDdfjRmWhm0L14qE6CcKwYX2IPE
/OHzNg7TJrM7ih0Il+Ectyfybifhbmi8VOPGXoJsZy+wZ0gVz5RO4FvZNN7PbS8e
XCXXJrhjIe554AYvQFBIeKlSnIszTFzPdV4ILRTed9WrHzIyZgX7N/jNM8yYD+Oc
+hgsD97Rwh4d2CooH33gjSqJssWH4ooW7j+mzDzEyr+kT5DuzA9N+GiQS1mI8ryQ
VIlt44eV+mxXFiVtVuqfznjV1FrIYmazCzq/z8viVRNPQJ41HRYF16qof28Rl66s
FBMvomLFWSydAui//55J2FePB9Ulp8HC2r9BHblL/9b9iQX9YOUdWufsrH9kPOok
oZGmwOjOJ0FADkYte5vOQx5n/AVRCQlXB6aRUMRetNvdyfsHHTWf/2ILBeWbOTrQ
lSnire3LiijqMklrUEEcS9wAerpOQrrli/BtpA6M8QFnHgbOUMQpIZyq8Gd4bX0Y
QF+nFznTI71/Cl5MnQo+dsGIP5ORF3GJoMpGS2mx17ubdVE1IBtXwDtxXb7rbYHz
10GnsCxCq66Q8nIrT07SdwiOwVqrPwaEACDhulQyjFfv7oNonx9D0cIkoNJEJMV1
ziYq+rc6/HyRJQBea7B8Xz+fv0GTnAGFH5YxyAiaKNhcqFv4pcpmhAUNMhla6M0H
3SH6oQxcXWKKYtxEJF4YYDMX3clemFlERx99VCUphRroRmbzzX3qoTZo84IVwejP
BK0XL3HZ9LK78m0biaTGUmVTj6zL/IQtsP3Th6+umRq/hhrHV9krGPFZVsQotbeH
ui2vTVyO0mZ5onObcZ4VoTGfsrlD2G+OEZXh7JxxElHvAn7FOlOstetfCaIoE7Jx
jVq4YKbXPElaNWqRJivUrFdYAzbVykzohP95ZeE2XpaHvPkhtr1Q7XSnJutzaZu8
5UiqMCfXXkESmLlzOtRyqjgZJ43eLFM1HILM71aCk6SQCoOII5PSMrtjmQOnZMso
KvidFS02K4inZgC29VAPo/46uIKCFVJ/DBo62QuSaH4QVZO1EaX1zBy04vkRVgke
eeRvQTgK9NRkOWaYQXswFzgXRZWz2qIsDI4baJHkkclKJKTgru2j8YB2KAjNrzVq
gVOBgkgbbm0xiRav3D54EABEaNL8cWiVnJeKKR6SqVEOGgCvXmjPpfaxnP7NNVby
5KxDweRX6ZoLNH+nqwGiOq65uWTnwagUIGWZ67ZJd6DtRKCImX+4NiANXhd0kUK+
7jkFhFOftzc2APNkBj3l+Ebmwp05NB2bYeSPapP4AFcIPmPgXq6+c7zTzaJ5pGXE
W+LK8hIaXON4FM99JOTBPvG6rONvkaBU2chalo90YYnq967bwMPYDA4B4+vu3l7B
+QScq8WDvsrhwPjBfKzwa1LpWEYT0HF2Fw05VhVCK8DA4zbPFZjixnPs7vwLujDg
DGPv0oh13oxrcVP6Q+vMnUtwzMoUoXoBESIhcfgqOdm8hkX1SOKXBmfGLGIZjUtY
uwbqLr/kpGRtny9BCZiqYFq69Y9A9Pdc4oLYYvVhnpCcozGMxs4xLLkiL/TYeOCG
cT4RDSrAkfTbAH9w1Wj4HzUWrX1GT16vQu8VDyGi+bXv5SrWVBFT/KW6vqpnj5k/
YNVEytcG3G94V652hdaAQU8MihrXnhmUq89QDFB0u7nEDBfu1FnP/5IQrabvwKPR
dyE1+KJgHnEslQHW6/23Ofput5hMgpfS5V+teyKUO4yzZUg5KwwBpOr6JXO1wZov
nvGHZjXrgTDCIiCmxCqOyaVbaVbu+xKq3kCqAAYrebAAQ8r71GCpn32/HyycDg78
sS7z91t0EWLrhN/cKKIhehHI6abL9DFPD3bM/xx4qqQmpaSnHWXQpSDozKFEfTu0
Kem+iu/gSQD8NN6FK5qpMXwriuBosvtvE/W8J6vYAjbz5zu34R/PUwSSvhbGHFp2
uWV1o7pduYtVkZEXjkwO7L+cZndVI17bjLyNV9cP2GekP3F2BYxjXXyElc1SBYCa
PIbf+QQy7axQS0VGDekmcUWDXVpzzQwIzPWmP5VSnZNcQ+GBehKr+YhQnok/TFpr
8fI8Z7kLpB78a2ftKF+zDyfFhBhqGo2Ea7hya5IVQtd3FVdSpn3NcSRk3s2WaV4R
tsi7hbLULAsa+njdCO3Odj71RH0cQf/pnx1bvpNLzobKD+Lmr/LMN1tX4lFG5O7V
ci6tpopx27mShqy4WE6fiSMmIx8or77mEXR9tk4d5uMHTZMpqC2ge7yhOyH6IKEG
z+6U66v8+DfMY8jMEQ64+RxMbzPEh1TWCcwbhzrDwF23nytISFlu98H9cH+WLQ8L
xYs5XuH0xZfRrMNAXj/fCl5oUgiDURjURihIG45FBk6Gj78fEcAEwaSnKEEMwvZW
3uwHaMhbwSU22cYt/y951xFQULsTGI3OraxNKz5C7EURo13SLG04TnPECDSaxtP4
cNp3n1Q8IUE3wNm98OKQpuL6lMbVEjqcilaTzP2Dle02R4IxRr4OSg7MhUxbELV6
0GXWHWV6vRq8pfeGWRjFAzmvZR+eqQfWZS+94m25blHgg7arI1jvth+C7zwMRZ22
ExRdHvh8Cllch8m9XTagZJJPQAYjAu/XzwvQmEpWN+TM2Dz2sbkbb2jVTsoIf+wU
21Sq84ksa3/I6LcFvKxiDvTg+8ODRKcWhr1gOEyoaD9fHAy2Ir5EkdWsiLJfpJ2z
ZHU8alqDol5wy9feEQkgTyYbclv2SklysL80eca5e0ALnmXy1319j8zsmEko2aQQ
hbwSjgokQ3HBK/aGnZngOFU+ZHLRWs6bk5Bv77QmmLADT4jvvceUiENLOFSJWpTX
WRvhv7ey9KULFFFiThCPgIomEi0rLdfAXDTOwhmVpZN4DKoKNKzo20MO21O9DBIT
qUe/iVh8Wfl/DuE+XFpErIiITuyAepam3kxkNytFmTJ0xVDCIDwQv+eG1GP/AFuY
+lmnPSZ6wqqKP7TXjvQPDcfUtFnyghe5k2PxgPv5qhy2zoyq2I8O+tRDuYflhZxQ
dS5qzUQA4QJTj0k7kzLZXAWtdCjMghFHGWJECff8HoSbN/skmH1d6EX9RMwZe92n
A+oXMG2aHCESGtqHZeoUrVKCCDa5ubaXTNbU6oYWGgEqHShmWfG2RfwFhmF/8yq3
Y58duqO3y496/4EX/ftzyWsA5rtpqWIA6guWwQast9TvakWYCsie77QdG1orHDjN
trmNwTUt24WnA74VP0FxSvdDliRblTD5aFgqKwJI/fZcf9zZDD4co5QeEcFINZP1
t1q5gWGeSiZQomIJPeVSxRFVE78j20WS2tWhxuWnSZa8u6kZBNyfUDeRIL+/jkD/
i9f2P8e9VNfbYabgOUCKXGPCNgUDd9JxBfeuixLhfe/eOa4YkY/JurUcPtCghbNV
U51E3Zq3ZQFVIg31NV1x8ynm4zdMregOnEj16tPF1YZCJKBAP72c5JdBDU2BbER0
WYrULbNSvlSJxF99aTqKobqdSJYuBvRzN7QlXpqqUr/VSCcPJf0BZNEnsrdLnxp4
zKpFoFsPQLKAjb9N264gd+Q6jK2iuAQ2mS5MRO+XjGy6J3nht9RyuC4YzDlxmXyV
lCHmj0FAmU/tozphqNpZzs4xkJHbVoB6850aWmJCy+ZgIYA2ednKYbonUM3KRwab
AoOIdCKdX4up38iQRhxj1OAgwRt5vEvZLsWOvL/DsEERhTdWZw+jKN2NVpyke5Jz
C4IYzliynPVN/4QE9yc+Db8rLVdobGCy4hQoNVAbYLcX2KJoM246xttQhxfEc25W
BRRdkJdybkARdfQKnrMkCoS4+8cUY5hvImA+RUMhal49M3UxLah2rS1G6UT9g0IO
uDoZvD7UO+qJW0efWP+7YXbb/GREe6IlrcuX7+LQzaVPojw6zomjCUwU4pobC8MC
YJ+BCDVHTVDfn0a/5AD7fPqomZm4NzfgyLqM7jl1c3aXrI3ZD8lnn3y91KvKH4Z3
m2kcRDtJfcYWcLA6/Jc7AiyG9G/YAbcjJebesS3i8XSQvyIKzOdirVuC6m/l4lV6
DJh+uheuEBB6zX21diyyspA3jSgWxLEwyfM9A7brha8XQ0+hopo/TDpFWymkDLw6
Iok/0UFbYsyzYjchGEuuEFb31N1XcsxK0HRs7rYXwDOYN87pnVjnxYHh/+Hu3aoP
iqT2pZw0CwQ0fUDD8Taxu6+vapDQST278JZFHkGC1mzJWp+2O/3YTgVkagCInNze
WanYwibiF4GwNW3oQANZUfGkxWYRQRpc1pTbkygzUksNAu2fl0akKgQ4ypSzZzBI
Z6FJfH9o8h05oqVMlDcrJz7AEZjlGRpXn6su53IplyAbaOluHnUNwTHkoofe8FIj
fDqjLv44PTNbdsR5rm1jVl4fo8fZR6mNcSFylI29QgghAIyBVwpNv2GwYaWbeRMj
rPKsOCa3Y0pGGe/Yf7af9pH4qSZout155eu06rZaAT5xIDv4dJxskj/JittigS7v
HO/6Gor58Yy1UHND9dK2UPG1SWh+7Z6qBXSoU6UArywTB1Wf1ZLqYp0ITaLb1Stt
4qL0QPAZKHm4yEC7VX4vg/BZnREuFcitC7BtfryQOSlo7sFvUZq0DMsWqyjSuhgX
eqDKYkndzMuIzhAPQ2llIXU7gukVASKi8CwJzdHE+WX3pNa3wqzhCGuYYRDgwcsb
40vIBJ0M7Q39M4cklWMBcYkrSo/34LKwr+X/bFqZWc0TMAmhR0uVyA8iSOi4QvA9
rDsXw979zxLrpwGvsomRUjmFJCVUSixYsCBhqDGyh6Hrms5eBqpgufXvyX4T+3/V
LMJWtah+i7yP1B/cgAowh+LIIVNTxDw2hrjtBUSVF/bVVaNIfKv2/xVL9cyj7Gql
69KAtuZnQw/2dL0Ch3Q6fXM1HbFTSf4p/DbTlUKhHM8fhK2u2smXceMAEU0T2QEC
8t/5kPVfv+cngG1ns9tww9Ul1bYOBr7bpQ5ewZBhSl6705dQTW9sk5AtMlyjB+6l
ujn0HeivTSq5DY27PdUhxZTpOrh+TkMew+VxX6s9aC8geYhWzdFxzH+ftf3aDi7f
Fhem7yFBHXOKFmOLR9jGDVvs1i+uYIZiLHN5DO3f38U7kJaLtJcgo5rUFfjGa6GF
j4pegtYYUpjTMsyW5P6NdF+g1f5qPa7Bey0pULNBS3PUb9TZmGoGzac6zlcl9XIb
3Epw98XF0EHLAgGKF4OB7zmNHMK9Gg/UB52par4Y6WuE1Qvhb8IwrbYkegDedCwD
54R0ljm7INYxLB0hOHsZfS4SnArRYitEJFkSTCQPWKfehCuGa70IaLXoXBtUWENR
v/Hva4Fs5jl1djEzUmy57qumVBRp1H3xu6l35OmVELQ4/Z+WgSNPhSfKDt2rQHS8
lsE5ai57EpcOTKWPJtczuOqVUzHZW0QN4IJctRJjJTQQPe078LIPG0FNoHc75p53
5GtGTE/4vE+HxqNN/HLr0fcE6FhZGkTgEfvkwFIwuPyjMPF4jyuwnDCEfo/A9qOg
mw4zeHuVbHfH3D28Ci5zmInhkF0nftQBdh5Yykkzilfs9lAFdBooA8Q/RalKljRI
jmO0TPKY0a9hZmN//AAWD4rpGmI3Kndf/75+Z51Q1XDfjEuHJaCJtvBHIZY9htL9
YH/d2Sz33Sjq/uRs77DgOZoEGnDmMfGTaedMR9Nl5lVdk6jDNwTyv6o67NKITTMs
y7sRExVQ7Or8jP/lRXzZQmX26am89NsFoar/+wC9rs0dd9hmfhPitDqHgZvJXFTc
2qfOaC3EMWlrstu6l+AMnMtv4uYoSIDeV+Ul7TL/79PansF2dg5gx6gH2tSF9jjd
x7GBxISqPOHKn+1mJ1Iw4r4NMtsCGnT0eg9eK3I5grkfd1jON7g3fKAcIyLar+ay
Vznq+Wvc+gd7U/yO9OrhBSBxfcvJYr1zJFWAcR0Obk3ZN33e1Sz4sU0vPbO8/NTa
K7YjGbN6lTIZVF8012kQyz+cYVffw2o8wVA65q3dcFFzml3tywNKjFPK1ZTY5RVA
/35sSEO7DhLU0BOcQ5PXaHH4xcHs9t5nsBFDdrElCpyKB716XZKoThn0EyNn2X3W
3+aFwzrqKYRW0tIkNsTvHiqLY47eRA1eYo3QhSs+R03ausThEDXeeVbsSGyDTPJ4
q49gjdnzubH2LXYfXvImIrkShbi6+UDOlKRenQeMzuRbAGEj8h7VZcijEz1pP+Z2
ruZVLnvdsCwMofbBLXfM73bAD9UOlSmZmdJbYh83YhpzBnorYu0XVKops5TTh5z8
CV6hBge/b4x6UjWnQkqiffb52kDb6HXxopZaWsIEjut/fBwa4DX7juOuMP/X2aNg
dxlCsjFJvXeDvZHeecvqAjRtjM344HFXml2o9nj7ogZ+BZWPPqnhK67MmSTbGEP+
VpR8jian+qmov88rlaUUIza5RgRTw213lVbKJFZKJKM2T9/t0IIsFFTiSPSxLFtp
mlLPVSfFE4rmIB5IE01/dRGGts8n9LTQolSWsqymuSMTIQClbadIFIxkJa2QhYAM
NocKyQR1eXt1aF3MW+IdH3Dkwtudqh1LT4aAEcSc+SDuzZ1Lpq4UrdF+zzMtSqXP
Urw66vghKQOSpvRBbPRT884wSoCx6E2SL34nO+q3XOhHYJgizUBNWcY7iysiUssU
cNGtyqa0mBgOv/QUGc4Tr3WzDjtxpMb94ABuylsfLzfjB/qNb1afhuBB6zGmDXJh
NdOgi791XcPI4a33e2gzxj/7VjhSsPGiS1E9AbVwyEIoSZ5YxpMmEX6wIx+3jJbF
ZFTcyRolmmBr/VxkJe4/3jX0GaRUFCxHINqxb/9qhGMl37epuTari/HiIJRkjOP+
94oz46V7KZKkgpw1lXfvSBpDwLCRXLQ7ddNmi6VJXIJStN3lRepcz0+0Wqg939L3
MZP3hgCypH41uhFDxFjkVP7iba/NMM8kIitEMUh5DaIcjouVaXTmoKft0U3wcH93
p+CeJfj5JmKymCJy7FmlJQnm7qmGf87u88f/hnWavDSAEwMVwxUWoV3ChriLk1Xa
dCd02tD8o93ohEwujZ8n73uParOZTt396w4c5mDk8INdMUFwuaV8OzxVx+nx5jF5
ymi0xcu7wZXgPy1sHdtA6ODEE7cOZjzwmfpR1eCotFEuWG9MYqm8i31kwbARkq+L
hZv/mASyllqRb3rbkKBfXKjs67YBji64242BM+ZM1tyeG9XGlxBPGEbkS6a/6vpx
NiAxLF17fjNCFhOClhZYDfj+5eGTTsa4nohykFRiultlCr2xXGHxoxkvtR6vhq/C
WynlJaacuDpi+ix0EfamkA0e5huKkGtwHVNLl7/GfQAzUk+7c8sCEyHl09fDsUKo
lQfNEUdDyZrX34l0exsaQNv3o1LnhEHajNM0v51VRL4h9/ew0YFynztuQzHYk6Z4
/m1VurAwLQ9ct/HVbfzomSGe3nfTSEkCgqhCSJhZq7dbJR6RxsLFuQ6dOrW4pQ9h
SflFdl6wuDWhFLDoEgjzcCg/SCEETxAq4wVme6PSDuDkhl9815D9GEQJUslU9Bux
5rh3r+dXTqB59puPQX1LKH2E28PjMmTy9jI6bpVVbezYa80lqHE72/OCGpi8F+nL
ZAFjlxBBuMrA8uZIe+v1suLsIa+5Kpc/Fqfp+AGLK4PjeFkU+v/ymevZaEU2+DfL
nehWCuCRNPMiW9KSeCO/PwqnggaGF7iDnSvNkuzq4zNVNT29G3N5dTGM/aqDfPqZ
ov7lZCoPlZmlgcfp1BOWNu8KT60Jr05RMiRAvDOH+8w4PSn3eX3W8cxuqd44u+pq
Jxr+TtEt090uBh6ltmjYRZZf4FyWu9S7d7Fw6wnTDATnXRANNQix84SB0QycrDEg
6bYeDaCwMZ5RDhEK2XCUXj3BorNlnBNVNYvVmvVnhYzIodRbryqEa/xPwYdD91kV
BW0yCtXwnqb4C+sWFEgxtHQb9gEE6BSamMJJtBSa5ms5cJt5G+jB4rX7ZCwzTrjk
nEYXJpMqq1tmMEYI9ql3eHT4ycKIAts9e0/Jpm2Qv7h6PIr7hNXJXRUn7YmAq/3p
iZ5uRLYz4gOjqb2LTtFHEm721mR7xEPb0Q5ZgbsNEb18arFKoiNYLsC01RWipsrL
JM/gAae0HXQn4VrVwxYM289FSaVkZSgPfFi99aKpp33dB5u+Yhggt/CZCRgsfXV2
hqN0Uv16US0BQpkXNyBhQKFC+gOzYv5omj7EJ27IBBUEOHYhKdZKTz5dd1eMyPh6
zg7ukuWhRT4q55XbN/TGsFTVYG8Yr75EjTV9AkgsyCfeGmiJ7UYLWOsCfbp+8/9R
gz6Tt9SOOSEb98UlbrW2CbmMPgwG8vkz8ebUoFv8m7X5OjiH7DmCpvlBhlr5I3Rr
WIRcHfJz7ZJAd9urGoG2Bc9XmQlRNo9E5qykMvKM+eAB8HwKh+UGQEO+9uTizVGb
ex+0b/sZo7lO9FwqRZ99a3jDjL+gHz/UfYyPjTFoqUM+FSdrl1Bdr7pAhZiu+kIq
caKKCcFfm0TTJ9krhMewqc+6J05QZeFCR0ERgl6cytT73E6ewj9eSoWrF04y+Ysv
W1JTnUoUSV2QxhgkbOO3vhHUXjrAU2HejJhjinL9ZiQcA0DWnHBmoKMAkDamydlc
N4IUUVo2FED7bMV8b3EhPtnCzopQlRLyjs/HhUoCsdFQeD1jSP1HKjT3rYQa/kNx
XvoQlEkJwUAw5diOtAtbidBZXA1mshOEocC85scxONSo0zr2e7zKkDhaX5KpycJS
dKb0Ipkkr4+w+qNQUcbhki9lOMfNGLw5ta4AbQlx5jlD2WvnfMeUElW9A0VdzLyF
Kxs9YD5BM1Tr+fwTMcHkSXI0KhN0nfmYXPvV4TsrpTsGgJ1A0u71HjQ9zts+z0WM
80JNvdbViqkOTMQvgJXjimYirKyx6SFut+15OCcUg2QQYshgUkkhZez17ZW5F6q4
J6ydsd9svqxf3sPbObYoM12t8aL9F8XKTRMxEXEiSge7vYIeRl6zNrtWqb84zlzY
GFAG8iqdz3r8cF7/9oId5gI0cgAgiGy3sLPkAsM73yqG8rH/wwQw7QEe6UjgSNC0
S4cF1/mUuVVdgCSlKKCn+jIuzyPlJgeIBb1wULl0/RGMZqhcBaNCkjOhBA8+SAbg
CKnagbeFDdZBsVbTZOpUMDK5Qtlf0M3gqSGxr9sIhw31gPVjRWwYeNLMaq+wzOFN
oKQ0TGyrmKyA8Csu89AIG+lofXA4mnMU5ANPcv1BIWkEFvkbNxxB8Z6IW2tU7X28
/QuIF6lZkRR7/h4ljZt3COmx8dxG8Vr3qcd4nZ7dbiG7+gQ9E7XjCR9iOrlnagEq
gk7b3Xqk1XldOLh6ExZmue9sYYiKM8EHcR1A5Tja0NdjY7H9bR+6ztLZhSLpR78Y
9u3r+59gv1zYkJBZqfsX+cgtjDOqtJT9PA0MkSF0CeZ7J0yDdCDylaAxC3tzDPmM
p82k/p+i4/mwaul4w0mA1cMGpMwrtgN8/gk76Lm2/d328gc1tiZNnTEud69mX48N
CYTb9ifXx29gz4EXHgyeuWmPzcMWGfCqBj5jt54OGy+5oOXmgGLnv3AXQqa8lYeB
nE9hOUf1/eWHzyg15O52Op1erPVgXPBOfwrCYGqJCVshgGc2VBvy30sLGBPYtTL4
OUeMSY9Nc5p3ZTfyjP0/EoxNQxjyLMJF+7w69S2uERc0+L9134KN0vYQvwOp9TeB
Ih2Az3X7/qIv6JQbkfgMdO3tARb9MeErtP6P0RwQmxsGKSuPrQCg/dvQpWEk+irD
9uJ6YC8y7M7pwf6hBN8Vr1ChykEYh4wPEdQpfc+V3DuNg9D+4s46RJqHlT7FJL5C
9uOPKduc92oRMEFjoOtRMfptXCIGbO44IFnKZAQHkLFrv0ibMM15UfGpl1UYPZsM
W9HbXuo4c0pGG/RPCQ7238jAL2KZjvWdquLFTfb3cLkQfg4QUDmCaa/lQFbo5Np1
z0N1YXqkY36pG3ebc2JJi0ZaBZMU9xNKpDTRad4d/SCYfJ/3ZCZxUiNgf/8OpfR4
4+XHf8hI27sruSNP29pkyvVUBeXuzLj9dzdmjWuSBkafSiiXpOB47xqUTEqg29dS
TzxvNHvfqxxyslYvUG9vBGpeaW0oFkn8GIGH4mX0rJQ0imIswi5OA98GTa8Yib5u
+R2oIHs0BawMUYvzJt3QD5ar1h0v7xG8jqsoF3eixR2FQL/SsSr/7q+nswPT0fo0
wcw6u0YVtkVoqYBN9WiiorNikv2Ynj8Cpe6xiTc77oM9N2JS67w30OfDcA59sdNQ
ug/7wa7HFlFWlj/VtiYSqwR3mdBNZAbLGxedzkkbIy85qFn6XzNqjpd9bsqh37R9
msCTJtztgxFcgynpjB2pqc0Cw7gc0+GeI2NtM3Z/ek3fFfdSHnCboJxt9kWoPUWc
mW7dmW0jIV8HDBrKAwjoaTGmRtbI2kHbyJ2IlUTBklRBiLpJ/qXq1mOxZm8gMjsn
nE6t2QLEluhJ2RI87Rveu9A5Qvi0jZrKw19+4qwNCmhGA4o03SPLG+C1SC0JnDDc
jgIakRE0n+3T6aE9F+cm9v3cQQ0qZpzQ4jkUeuKgMjKcPIMvtYMcES2nEwX58V3E
fWiGja9bwSJ1iOXS+ztZV9qFjdkMXBby4AcxseoC3r/HAIO8lm2TwsBwqJwELUTq
C5z9+EHWnTWnflX1TycKivQnI/7r26EKhb20AT4yCK0GUCInu8nYTqlB58UqPdpJ
Hqzx17cMZal1sQX5IgwjmYQDwJCSSPZ/8R+dsqFBRKeQBzDyffoWxbRVIcDfk6bu
9i0LVmxYInf9NIkVfaGFEpiWdA44fCupt9cKxqYunFy2CKDq6gI4RmeJrg7VomdM
d5/6B9Lg97Wf/L5E/AJ8Ld4288g8l+aLpHXl1m7xMsgnAsPeiNJuwn3knBYRy3DQ
fp8SIg/zfGWP4pTAof8l7dlzxCl95By+zhKPDr/Y2f+OXqu7srayacmc+qXalxzl
yY/gTeNiI37D88OWD1BI0zbcso0iGbT/zPe9LIvdraPNrYCEoBRKqP5jzQvFgPw1
5G8GBJBbeICkn/pYrOOFOKyhWEfL1TpP3rPKTdBa9Pr93eYFRCthA/KJ6qbWVs+9
4Tfv7i6koti2ceXc9sP+kP/egya3SFYrPEMU2+j14VjBc6aS8Tx5JCnyv01bZmkp
W/BJ17GjyrAK450c4TlwHT0Ul5BP2jxT8GAGNd7eykbXD/aNkVBn239oigTw7gzv
+44cz8hfZwyfwQDJJNZw4DRqKDTEHvpg5Umqn0k973d8BTFj1Mc/8ix/RTZ1gYS4
kmwjQ2vej3YFQtpcDXNVQWlYpmGUYKGw6OHXzc7qP3BLwnA0SZzvksIrLazsQpMQ
5eFW5dCGrzS8AJtNtlEZoXCt7MYuU1Lm7I3F1FpRtEvv6bhBUruA4lbniw2j5oRO
LKiRHf5Y7LWlUDK4Sgm9CEt7iZi7MyvsQW8IQ9j8N5C670LQC/Eh4InDAZyhUXcA
l3zcYmx9JcP/fyA/CR+Ft9y5pJ+CeKsSoi0oLKhgFXDae8eEKmWC87LB99JecOsE
b2LQWo6eR0F6gam9WcaBzjG15vBJk5M6eKjuDlQBTYsj8WBbgQ1lFeK0rRBkWRPV
VvI/74+nGKsnIFLUqtRlR4Y/v+DKYQBDQsifKAP/ylXta7bb8crY+dV38qAgzhac
4QTJ6e6Zah+w5bhgmM47O5bBgrXj8cOhuSP7hcWKvvjhFlT26/M2MzLxg20CHBGk
5A1ZlerlU/s2+2bMjxPI02LIr66B35rBM5ynh4W2NZ5aCncHjXfA/Arb1Hj7tlxr
HlfsH76/ZIeEZRf9MSTUqHgKkxiDIOnZNg/88h0K6dKValYZX0msF68j9DxzQ6sq
emRPoQVoGdCueRG+JoyeB9DWgv2o2XdBNJXdphEcn6V8jjKWL892BIQ6L7WI1hyS
LaT0KaMqvkEeYdzIc+uuvVq1oNSyvMBwLKE340N8qQZr2xXc3ZoWXwKR1w2Ig+eR
sCSkICWTCmppDNCtL6MEGbMj+tug3A9xBgjYqYjqpKlp0qXjZm8ND9O+N3FeQ10T
9KpZbAkPMdXHgEctozowgllT3WTMD6DuV67sAV7ATuhnR2EbF+BFfnystm3v/Yq/
yWpBJk7sbUJJaxTt/e8plsRLNL6k2b5Uxf6+NKZRyplWRo9M38lySTXV8+VLd/WV
0rOUZX+YGg8PQpS1p62BzVvOIcLhpKl+iVGZxDJZ00mmQ8MtjewRuMQAiXBm7vCo
5Bg/2yWsNunRNL2nepGh/KjcOX/6clFePpIWG6pexqIQnNGI+tOB82nQ3MLgVXcp
j3MBwS7BR/7P4dmdK4rnhhz35Pb1gBqTFfjgoQWx6JylYPA7Mx7CMs+6Ijn9yOOL
Svisj0rc1oXz4BiIoNY5ocl3/qb2eo6mRyUbOUhKn29Q3Ds532rgA0w/y3Qv0y0d
SfaaQMPyfoVnHv4z5r/vQobtJQsePNeC3W/srigk1beZkbMiIigHWp/7+j+nmlxz
6wf9prnHzMGPJhx0865uCN1+5anQsrSY/VakgRgSvRWHHX0GmQe0OllOnvonLK6p
ljET7WQMSDlKoSMfiUgWM/mZ6w6YVJ/TiK4jae+cnRGsAL4HCHbaYe/Mx4tM2+t4
hNkHjFCU1eq6Us2aycZVLwOUGqMZp7XyHY/phm7r3vM+felflm5DuEav+ez97Q7b
vk0cqp+poxZyKeQPyWIdoHSR67V9zaaEpITDUCCJwUMqKC/G2OJ+xjpNKo9ehnIR
JPWMP58INpHcgehViTbqEhjKpZqB64IOLitm9l3044mrD9b22/TaTGuEMat/LKlT
LZ5anIMwID0wjHtII+YFFrriIxq0Gh4d+V7pR3ZDNMohz5PUoxWGGJv4o5kPUjcg
MLGhLHuXu7e722IyFKEhDktnHjx3ad2lbisj7WmTn+pxGzaNnwb8yDVg2XUr8LYM
DiMdbP/obV4WiJj8Q2j6NE1rV2RNbqjC8p8zOpiLAYGfEHRSVc+w05vCIMqI5qKV
081LhS2T4H/WRCZOEeYhJBpDU4c87c1lcnmV26EdpwlWgnIKFsoBJIL+uoFftv8D
RtuPj0FbrP+ts8GTTnpBOy76I9gJabkYhcgmUK+xdPtt3QM/arlxGy2bvGkZACky
DQNPK8lGVSRQ4s3ZNIF/Kg9ogo6CbvPh4qv/TdCZWskcdj9NiuDj8rRdcCM6OQiF
rIHLN9pzTRwc4qQhF5toN1WNWxvf/MbVsfd+jw/WMnJ3pNf+a4PE8LZEd6T8nsHD
w89Sgaz1w/gprg5eT2eO6piTDTya4dl2FAmP3zRLZZ7cmIsnBgmBeZkFltxu8mTA
/EzP+PGAtFl0st+iryyqfH8Fcntuc+dHu7CMul/juS1+OM37oQFQFdX/brQFwbVh
U0KWZV9hek8Rxy7MOA03bua0tpOhwrL8lDKEzBIl0hsmnHgB9GJ/MCQaCFNv8G6y
ZTuN2w0CxrWOE+c0ZcRghvL7aCVZgWtqvTWW9+a+ND95y4EWJvvGcDdIDBKhlsyq
ZmUIZu9clSDd242HGcNQbZeLn3RWC/yAdI3F3QcR/dYfzHVEy9ZyjElo1eNTeWrl
JoH5eEFy1yO8xp/l/5vEZ0USZYjSEKa6n1miGrXVC47gcbT+EuXEau7qJpnolgqa
LzIdeQuEofAn87Nhq3/+hpG3TVixIQ3cMXJTs/beLmA2HNjv3dJtD5FwhPP3QqzD
mRxSrzCJP7aMWqS/TNg+mFypmBX1QL/i12aYE58zhn/pen7OSEa6/87zXIx0zOe2
4Va8tHDfT/zUOzGuFIQA43FDXGXu+v5bdM6Femeb+dd8XQF9KqlhuSyUlluBIL3B
LRc99FA6MqLarsf0omjFSBvQrWl71Ef686pqH6y8ev/vvTUXQjQpQsVFIKPgF7Mo
pEfSdQm9epfJgzPjpA5Lj4aqrPNq7NsV66L2XZhayqr960G94/UkJTXa8bI+mFao
Eh80R1EzAWaX2UZJcGwpxybxaqfoImSeEliHhGP0e2YTvsL9ZUvrQs9+0HBNME7g
aBerhNF0Fr3LS5o0VUqO5LQqs8wn4ZemC7GyjPaOs+qz3zSzIjCJiq1MQHvNzrIo
+nMwV4SPQCRymVPhOgV2rqxzhQ8NPFMDHax8FhkoJ6l/5SzbA53YYcWDUMRk+BZu
appJfRhi4nywCv/yWvf6OPePda7qCI8pzgYanwbGC8EKJ9QhW3k+4O4HBrCdAg96
FIDMSCQS1voNEcpjeKBSLmrauqaRYf0mlGW1jcZI1Z78BqPmphYCwjgXqzijDxqw
wgr3v1TecGt/kHS7P+VV4WicCkmKtWeYi8kx2+rZCd1n5xxvnEFjgTbOBkLcNW8w
C19z2Is0TooZ7CnR+4rx4KO5LyUw4NYsPz5aNX+0NJp45H7gQU8g47n5/JYCwcgK
nTJNj6HTVXdGtFXH+3IaKdnjF7cg4cwDhLpfeoM48YqIx5TkD/zW0hGdphl0QEBC
o1esfHRYCwftNaTWBHA7NXxPErOo0ourm2589zLw88rkgPSBMTtTcpGHzYCT9WHd
gEn79FvO5FO++0cDcN65hVdXkZF3+yzTtzII6x3bgnoJn4IKBEqDoKYj5TC4ab5x
Sxo6ws40EYQVHulRBlmPHAxof6mKW382BOcwd3Bblo32gVEE5zplmwZ1nm9gRSOi
yB0lAra1z5Ke1qbP+KaQWM7cDEtPDgjDWn2y7nKAzrXUlZHSIE/7Ojj9wkrpeBM3
K1NUxw0N27zymnowjhYpXVnifuEEGCZedeTW72BADDw2qR6mHtPi7kv6hBXJcA+s
EODRUH4taGiM5YOugFJvhik8m70ev3S/AN5QZS7227MNzu2cLRTjkCoiGLCp4sA2
7vM3lZ5uELYJLLlqDQyDiJ4GK50mbnN3ZUdmptJ/bA6bvlZpDAs55qEIZmxYckoX
57vDr4F6164EBVRuiJhlDZCgWS94vx/a2UAS6RcFxtW7J4OFgISJ6zMgiqxAlSlx
ZclDTCmFySlApgc46p7xRLvbujatEL2ighkp0x+a1uxlRJU2ipBCVCiEGp65jWuS
WBuqDwrK01jF/mJIlG13vKnwQXn2YauDdk/OGKRRX65/wFEi1/6TKkk7jnzM36um
S1RxzGVWjzuEix8++0F7lymA2gZwbCdNafTGt4rHP0oPkQ3WjmSDCp79/sdHLaaA
nqFicxCjUZ0Tic1j8KLCf7pC1rlb8hKZtRFyfnvaVBvX/kfpb59Vl9EgnKcRy45u
5HhyPl0UnCUzOp6aRh9Ar/ZZLvzYjQG2D82wFyRpD1BA31OTAyTnOftxv78+OuEq
3RkpWmqcves1T1xQdtL946YxFp+W4volyI9HHCzy8FtV0vZUPZBJGC7EA/QHYUT8
XFu+aKOkRxqylMSqRp6V/+Gb0LBZ9z86+oJiSZMDV5UyMLzul+w21JlmH9CueoIg
JBDbm0TH5vhMgzMG87EW5B4RGil450nKOXYtRr3bP1XPdiUA/aMbm/qvQdnOq81m
dnYJIri8ZKrcibFJ6v+wpf6Wp5XaN3pahUTD8mGO72pAKLNOPxxJMF6vsRZfNv4+
RnZfD2VZD4zserxxHOStUC4kO5bLa4utulu/pCH4ItEgkPDNYKmYYYLuJkqSwLDr
uVQQ4vaBWJB7//V2AkzG0F3eNuBzDHF/BTuC1kEXfViDJEps+75dC0qPAsuPzjpQ
2UBvztlB9JnuisUcIps9Kr8OmGFWhFgmJxqGnpRPb/GS0403LYrv/B9Y2gnuBLs1
ct+gF0/lgiquc6CLpZHYrU0jkirjBWIh2pM0KbN1KEk3gnA3WALqeu0RAhpSNG0Q
3fHi2yftreCm1++eR0XVDfo8XAmxNDOUys3YsFcGW9/e/vcI5Bv9FdPkc1DRqYax
z8TnFkqbZwFpN98j84SsPVNF3foS6WvF4dS0Boi5quhBFBWsZqYZcEdyiEf1ivWt
tAxUrknx5JZh3HXKkmyFhPEWAqFHX1w7TRqdnQk+eQH0R/3Co0k7Nu0vxhH5wAMx
xF5Mv0atDV8/6v2Q9fIRHM+tXNxdLjgSZqJF3LR3Ja6JVqYDtA/tSidqQe6u7z31
RQRHriHwWO9D/e1+QBdtOsGFRDLR6wzlsCTlxO8eujow2PjsF8GTCgxRvH9cfXP4
bdNefIL1zjlgRxrDqlyB/3jYR99Nua/ahd6Qvd8UBDWvkhqPC3lU6Ohmmp3z9Oza
SM3yIRX4BaMaI6AT1KA+QC82E6OWXZuosHxgx8vAcdtCVBX3g7D9NXqhU8zbhQAU
zk2uQYdHpt/xLa7DJ0wVPDyIliYMhovRZ/S9Pv4Di0kgLf7OsrF/Wa9Kdet5XoFO
nuDpPcw86FUutsGy9RDW8TH30HCUXvlqSXIWFp8w2o7eNiZQyTxu1gGHUdiKuiTC
aE6e6K3P/7hJ/tUvRB/gJw4bbUh6gDv7+ZE64D+0TkdStZSNkRMSnfnw96DXEzZQ
jXPDZETJYBSybGfQze+8gRxF/SaWPlYunyMsWy0UGW1kPhLm9uHrVHP4tYiOnlM9
lLjDZITasI6EQyz9Jpzd4xHVFSlotun/h5ZdJSoBjlIO/YUP+dZiTBWUQ9AjJ9XS
8z09bXOg+IZ9rLGYo35IQCtnGsa69cZ6cx4ekWa2OHTog6wLoKHwFG6VHlPweNvc
R6L4okJ7dWnHdY4zMo5Px8L6m3r93hnploXyqQDAlsC7Xaw72XVp+jeTUlVxUeIk
h4UNhvKhReEp3zIovAJrYBnuvtjJANymi8FNgPs7CDUJYkk1kO8sm32OCi3lPCmW
mKB4uK1vwJcVzYhyygf8K/wf994SHQglB4pkhn55X3uxywI4/ikfHoJdnHvyaDtj
yGB1TYV+LF4UFJ89Q0j7dP7+/YUy7Zz+qlidmHsIqiw7kRphBbnQxB0bS88WJpSG
TH/v2NkcUNpYEQ0uZMJhM8KiWmg8dwlvnwCyi7H9MH15RknGPt17fZpfH7wdiWj6
k4dNjVkraBLViysd7n8b19J1ZN1D7zDy5IAFax5kHpzVzctONxiqVVGAH1wyOEaG
GPTipMRJbSiaZSfdiRDnQ5ZNwQ4vjGkTPK1f2oRqLLBqi+sWeYEsNlFfp8ZFYn8l
fUSHFT0GxvIVwPhM+JfDLYyE1VSgjuRM2QpDwIId2F5qGyGFLRZR35cPcQ9YnsM8
1+IDvxeLfN8OSXKoGilCbUjqRIXwV9p5ut/ZvXXMAX+JVkIAf59t7+uafzCiiQ0h
odC3On+zpJ0CcIJra+HwYajaw+/9bT3veqmOtQtT7nSPWlug20zRJknpeJJOiDto
S96raAjLbTojvWj8vJKkmNyCRsxIOAie0D1+GFubyqw7FPQyPDR/y6LhWqmPofGI
oVVzfFL9FnR1rrjZBsg1ZZ6ss//XqJzt6Fm5j9rMujgJSuFZnb0QSiLNEp9p6Ye5
XZzSuey1qQrt/Z032cqaL1FdrfVdtS8tSH8ZXKEYrxmVFCp5T0LSEmktmEXGhZQW
MQGazl218YORLum8vPdNfpFQdqZeWr06aXo3dGreXWtnUGeYSS3rx9gCrdyQDnU4
OSlYtXVd96AiGsgi2RJxLheFOGIDo77+evSRZo5Q4LAaj+78vTH5Iafo2EvyDG19
V8gTdhEBqKYEkDKHGUEfRRwJKUWiW1TecX1n7zKssRQizNAi2HfR88fvG/+lfcDQ
7Gnb5dU3JZ2dl//osAA2oNVZ8jjCxqZjTqhnIX6eITvV83bENExijB8l65qp+DQM
qiIBJacZXYa1hgeeJvrpWtKCVfUL04RN8aab4zE4gbIMvWf14q/772cAfzj+XyzQ
mwLylZtJt+RcY7aoXwP+/BOGZ+8cIiu4928vWr4QnGwMXtxlGrIgzfP+SPbbwBdp
9qCitwVRHAz+M+QAOHU0BEv/oyzlJgBW6ygaUWct7blIVha4MDnxHVi24kWvo3x5
KD8theW35mMjK8X1MEZIC08cdoT1E2AqYyng22qHfAUMaWkko8EYP4G0o1L2Fz9u
YKSszkhtpUvv+S5RkDnDLo0W5MUlqyHWeXoWUnG/9gRYZ41ZkZrGnWRKOxq2uoLv
JOmbT6IJW35mNDaU/OKvN6QPE5qAGM7nw1ZpOrEIEhu3cd0/O6r43W/nas1FMZQq
QKRoe8Y2XWOSX78757csKAe/Rehv2NYnL2XvyrGh3pqNUvHKPiOuC1gSBn/yDLPA
NykajwhDBMBwXXbEQacwb0TgfYg8Y8R3kxYVvpH6P3Ess4JWGa/6DLXhXgQjAFBp
k251Q0SnID04wqezdsg4mOdtziuiaig4vwN57EI+ZG6HGh0gf43g8hUDUmiOKCss
9cIVwNp5Y+lsSJIzPpB2zNGLFKzq/QQXJFthgQRNGzPe3XJb3LdHf+3jMRYgRLDw
iLZUh/n2wP3+MQTzDh7pU2xxmSMcXnSet0awNsW5u5pie3ZCMjRbasNQmlv6msIA
W2o1Ssr9uX9hJ9Sig48du//Vu0mcl/7SexDQULKDTT165A0PxLgQrug6Eqbjau/b
WUiKfcyxg1H5SkyEj9HhfQuEtfHuh7+bQujjYftzi33w5+FeyBkN98/gz1nEs0rf
Pbuw5JY/XoK2jVfpVsTZ3flhkcYvVbthMjRcL+n43lxcMSnGS1pnc6ykScNcRuDJ
jUWSKdjkXxMs8ziMK1HBpdp0zFu5lUpMZJ0AeXA4p5yX+DQR97uAnEn4beGqpGJW
iLlLchQQ7BCN1jSfjDRah1TGzna9nvROmHPSg5XwpVXWAgWFazp1O24uJooi/XDn
zuaX2S43DNpdhXaqs8ZGSVOq5mj6WHWYHh0P4stiExrH7ll3+xHmowBTPpIuKpGO
RmyfZCNAThWu3YikrkL3/U4KmZQ+uS8cHpRPANzvasL2aQoVFznZq8Rw8GXXVnVw
c8fj5htH73pKAEJvPJ8PCFTlnWV1M+BgkqbxRe/7N6Lqs07MQfvQOyZVmRZiR5di
Q3NSSTCJ4M6eEM+1bJ5QgMWc2whoykhRmCZZV/5lL1JTItfYs8ZkLhibOWmtl4oC
Ky27tO548smxOI9xMREBdMjWeljJqcwXZU+fvyKqUx3thFX53P9LTcEk2g7i0h4+
eGoP8kjkp09tg4CH1L4dvSkjI3X8GWsvBC2MGnaCuUjQ5SNZRs367tC6KSo8EU6i
N7+Y4hjauWgm51COUGBL6i1hvPZ4A7Br+oOWZRGCVHNuF9ijUk/31b9tQLEOoplX
pE8XNSD285niWRNcRgcrrJ8INn8s0IMXxKsiOyrJLEAfHY6g93ZWhsDlPqAQRDDD
ndizfBcUcOXY0JB2qZUKZ7qEnQNfPcd/kNZ+NBlaAo4vdZtyOZmQgjE/KmudxZ5Q
lfQNrK75xXGZkZPXI8qbi76pWUmDn2+/QqkOsqJyzvSzBUqeytCayM9mqWiMuHC0
5aj5sX+OV1HIm/c4mUH7echJZnPcPzCxQxsCOhBSoCdIh/Gk+j618ZRf//9sOL3g
tWM+p7eEtmKUuw5n1OJkhWu5JppDiPwTuJUAtmVQhwZ/CQvO+25O+F3FYsb7O7wL
CYygfLQcAH+KD667fxmsosOm+pfFl/t8s99FZJf/UT2lTx44+apCfOizl3WK91Qg
3hZx4fAFo5a/d2tiJXnvZ76FbZebkoYpKuvvh3yYiP8RvCMcyb+MCDByv2LU4Iz2
QpmyIKOM1rxAQKaLFoX3MgXfAcTngHjvSMaeSuK5xF0Fc+0qBalyQsQvIfLuoEmT
n7bRiaDLdnoUcLqkFBoIQnbLM1g1grEpTBkPZjUczzIbCkZSpqj0rgYZ9fwiDBXt
nGy6Q2dxdUX6euRbvzG99r1VZL9gLKbB+9rlm2SfvehuWbcLbS3WMcQT79SVHWCc
1ggbXu1yabrgPdXZ/hfVe9dJasLl/DQsFbADggjnYcwd08WcT96gwNHC/4n0HChR
NNMnHGhDFP4S5zdEAJn9WI6wuJFJWFvzjoQdZrlKjZXQ7mTxEHOOnVgrv3xWNkTw
URB5xPQ4udjgB9miayZMrLrFaMsxRRCUgXZ3ErRXhVCQ1mNePwA7YPPpx5pkKjTI
U9pFQqPaOju2dZlVXK+TuDry92MJnILL0UEof6GVLzPjkgYNOXhTqmZRXuOB5cLw
zEkQHHwtCLH86W3bFsnxNCqJ5zh9V45sP8y1dZ/8cJZVCyIEAVTBgrTdsj5YvUSZ
210z7OAhgi65QgZm27K1QoRJnVwxyW0N5kOGGastbzo9bWriF74GeoLKp3FgIqLP
FgA+vsUTjBXpMUga2SpZY5CsFvInLR0pXMmukMsA2KWmlRp9eZ65Pfi9VQHov3eS
GbbxdjRaLrGa5B7vtw8D3ZdkbbDxCtXFNBaI6PMx05KPH4gLwFjY0Un4e/6ZE/gN
S/nZ/vg/cMzd2fPt3zz6h2OXP+gAqUV33qNR+3kgkMHds1ElJqyUVhNHuJoE8IJK
OYQzQAaXD6uTaF1FFCusBYuC+rjt6Ry2nQQm8wKy729091QTEQbDy1cO0DDZUitv
DWCFBmQ4A6Rbjm9PgeaV+zgMd7DVoJNtuUuSYJBk93iCarQtlSMAX5zgokKzCdeK
VuctOhyzgwv0BN9AIcMDlX0TRU6VXmEJDFmHLr47d36vldDONSJSOiWBU24cazct
zjDm8XyVxYSW0jSn9ddJ9lreKhfnIRCeaNC16rX9RYlF82WZTvCKVK5OykeHe1Ct
LTwfYhj07o3jkYhBh/oXyCg2DEMaBhSEaVs4rgLgCLpB2MtFVfL+n1svfn3SDreQ
MbUKGMiClbg2DsGQ86pHSjqs99KjN8+PZyYMl0ODwcRoYrIvwUwqd7OBfaBQvEEc
NFCgA69HV/TN+/jRmFQW6NLINmQkNtwq7pER8+0n2/0w9m6NGsxsbWYFjwn4AB9E
4hOQiQRQDBT0rE3GZK4CqgXtmy8Kx1Cx1F6N5GK6Kz6MsldutReyiC8BB9/rsZmQ
B/6Dka+pVrG/ZSAvLMK8XqG3qbptlCJGsQNjl6yEtmY7rGB9M+8wPec63KxH5nW3
UIF+cpAMROSsZZRKW61hThjClD/2NLLfoeqldulZg5WG+xDQBs/FMeYlrFPyQPKI
8RmzCnrnRI/oltpGVAmImS/hmtDbf/ywdVf02RBRV21ncBXWKxiAHggFbpPJQMCj
kRqSERvfEqyay95UpJhrGs6Xb9CK+jKFtf8O5029V78d/qRTDzeHpzFj4xHwctBn
BDer8aBlYJVtLLtuqqQD+LjPD/k9ifid5bOA7TGi4lXcFtO0Uu438PJsrQ1FDAuc
qw01anbPE0JHyI40JLwkyu41b+kUqTqFZ8BECcZ7LHnl7NHn2+qNP8Mxzz+S6Up0
A6mwrH/aoWhIGzEUiOiZaIuTv4IhU1k2PGTl31nM8okxEqu7cOfD8P89/uSX9cvv
hJb+8Uzt+6sjPpSgg8R26TuoW/AeaG7baLu1yJvtFBLey8qIerKfrMB1Dk/bmlqN
fvQtTgGQIS9AoKfgiybs14Yt5ox/CrbLhttY6xDPWTunw5dCcorKiaviSA9wjTKV
zAPB2qamuLhefoU+WiXivTZGQnRBi+KxHdt1Bg6oDEQHzAjd9/5wOPy0d/Q9MYYP
F8ySLE2oMDcZJxdTG+tvfXn7+Got0cZj3xvbXBnH/3rnutoXU4joa3ksMlTX9p7E
qqgT7UtY+D668LBG3wYDI+jl6Wm798HamM947rTfaUoSDk7GAE8JiH+uvW52KzId
0DPdBRV36EKM+xS+CTbd9YR8boC1i9sCcgaXbS3aivVb4P97Tpmuj3ijlFp1ZpzE
5vInoLEHoVZqOIBdkqbhnd37RhPvqU9mR7B5F14HirSLqpWtk3tav5g4z9eDQBvm
ISMKL9VXhJeWd6HLFuxE1K/FfhThBzZFmaHFhSzeuR2b2AnCTSSW5XVqk9KP4qiC
L1yNhFLd12UHog4C2N5MjeYO2F1LpVLkXCG+d7ENrSchvLlln72bvJWOCA0sbPm1
jgVf9Oc2ER/z6D96562w6LD8+BTmkxmltENqpWcGFkWIUS/YRlUGyfocj5en+4dV
29137Qf24oVYOmqmRq7OcF3v5GrzgFSMgtKkJvAbWYZW88VrZ4LkoOc7pjFTCfK0
rr+CJBvQn6mVkC4AlucGt62QrWO8J0EFsu9v6C6QplXAk4twibedNZhdpnTps1Vc
xyagnoH9jRmAAI5cchbq5HY5Zfmqh7DLxyGYly9qk1uvXdGHMtMapqwDa2PTwp+y
IjdXROWpZaqBjIHFmjkh6FKxL6PkLruPuYmnWZrdJ8URNSEqiNBmJtXjlxbgqQCF
OX1plsihKNbyCsiAQ9Dkn1yZfCkHivaqK9WkjD1/Jhv+tBBOzFNA9nF7BRUtL0eQ
7rJ7LYR1omQ4maXRa7lALaOoQbix4TXBcQ8AXRE0OC1PJlcJqwPwg6btHP/Zs74q
MZrJS66r8fsWUM/MtkkGnfgk2NETTkTJmPSDxU1MBO5lVfUj5/2ZLn9Ms1z4ujxA
49eBBiWOWBCcj+Xp6SFkIkav0G03hEex7LyabRB0b/iBgMH0qTvhtzbB4lAglbdf
3c8rkam7ZIn3F0khAxWba8l2V76oJI8mjiD7PZL1F6PH8cTEMa0kC0Q9yCJNSMSc
pHtkLn820HxoQy6KjhuRlhbnYpe1nxy7IHAXn6zDXcmtIqQCzT1ae6rfT9fmCZ12
Km1XsA7CsMXaasocAzo6AcAex4LOeFZkptdf2ezHfkauNU+as5aAloXZP+8rcBxW
tYTua1oGExzCZ5lmERa/zjbIg6MJ5Z5LofiJO9J6Xy7Pa26qHNoMCfhpjD9eZPVQ
fq++srF9jfpTdnLNb2N8fKamdpb3iLYVK0o46Ji9IdLUSGMhhpPPjtLO8lraeuvW
29lthWAxuIUeuS16pHvykP5FYLzuwOZrAsfhidsYTwyCD4uL99iy7eigbIt/hgdV
poG7B1nvPZdNfyv674NCSwI7wkdbezAX/JkuDyGLIpnqTr/fzNjVmCCzl3Mg7oZn
qGMkVii9VxHw+gj3C47HiZBwZEXOQaiuD05uz9rYKSQLCtfBF/a6FxWGjEcDSlCZ
bUgnLEveXHhtpMb/VibigO0ltYMXIHynRJGf3GD3kn2rJfXhpdioEr9r2GUGvY66
sVzkK9tZaXQriUYZVkj9L55CVWe3hy9efRhqa8a9zRx9jH73GO1jkHcTZygWZc5r
JxPEQYUBCNysBWI2l50MMUI9wXIE6u+CgHn5ae+SXSegLmmb9BXcXhl8LMvqgvsr
t8vszFhMzd554IHNdfQRc7/BtjMJNpFo+WCuGDEUp3BWR4jXTJB3Vk0c+mRMGEyA
4OqwWHngTMZ3tkdoRyL27cU1TWwDEE49HHGvmhN7o3t8Tgp+j4qNoT4JzMerS7O4
J+DBD7cfsfm5EuPPmyx1GG7HbRCWi7SlXZVBBG0/dX+Amp1Nn1Fr2ky8kHFNC4TG
zP7IrwNMlG2Rcb+1N5Oa9NehPaPBD/iq7vPa3WuYHeCzRJ1VWuJoNlypwMK+nYPP
/wTqnzGh92KJmMEWuyZskIxyIE21q4tGPOzFBtdRlX+1x58N6FuxkFcpC4xdF9qY
VTpXPGpdXUx8Sb4lZWNcmEV6d7gC5xPHC26F1xFZRawua5dFUS/XOG/jVs408/OA
BQdQ7tyTH0FlDT2rNf/I09OvuOddUHLVODueR5FQ9xoKjwcO+oZrFzFMtM993MKO
Z1j+QF+kNMaynv3F+NssQGigt8ixR2r7YtC+irHHQlQPIp8hExurdfA3kDqXwdHz
bExrRxPC5DqE9tbkQOslwBaWu/WZeGYYYkNpOykL/3yxZ0LH5UvwIFe/01g78Hzi
9dbv+JVwPrJAL4GJLEZmQNFrtU4BYjOswBKi40z54qhExiPQcguC2gnQdrq8Vlc7
CEmmT9PIXrRFmWKBjWavI+kVLM2Cr3+pPEA4MGIMJmL7Q7RDI9vDAfff86bNYy/3
HjG1IYNDakJZeqa5IU6nS/T5mejyN5W7iz+K5SWs6i7+mrX6ilKpNlkLg4hRQ4zu
+3JInj6XeFPPO8LO7i99BXkwSI4Eskmj4U/uJZ37FJpPeAwH2d6VIJ3Gf8uIQgkj
sS5KFLmypmzeq4gM7KKcv06BrYmvF1GFBpiZbpietfO/94WBT8tgBuCWfjaWsU9V
esTsQofGH7vBBw4555hlz4d8WT+vVKAK9FNqdb6aaPqOTh723cdpurRMO4U1oJWx
72xNQxJ0H+IsqkomRxwzgQI34cRQSqYIVtQ6NYjZu1OkLQmYy37PvqCzYu3PYzbs
Qoo/plIDnlyKt4Yow+gF6a2UbnLnHHl5fCfCr/5XYcPlZBgrB4Df+c2xvuObdS6o
zGEhrkcYGQhwfnTeDd7cgL2QH7Am+GzRX5mGi1CCQq1go9po6rj/VAguwgd4O6kM
2Z5NJwhca5UrCuPL3aWDp9DKWG3D3B2oM5ZXqQuUfSFyqphel6U4racjLHx7dQEd
svfA46tRYQNNHsylICxu3ghalCU7MUMe4OLWKY+lr7kwDwTPtebGTdn0f8N1apHj
eJZw9Qbo/xchi4zGpmjJFna3yYch5sVmUfQihoqlhEF16bGtu8kRfvzTM2fL4eMa
ONv8wEAm4bgsIsEZRZ0DIfg3ngjQwCbPy/S/aQGcSpXxBJ+drsVJLxXxf3pagQFl
VaL0ppqkbG0g1N0WN/fZlKq9A8uhjugx/QEVNln0+tmVbd6afnkY925xa2YY7Zf8
zp8xUDeoOkA9qlR4p0diwf4g9gbHR9rUDf4D7vWSDXWNZ4Crb47wex1qnb+kS8Pt
0gszgap7bfCXl1wC3AoU3mtnMzUG2dJqnKVg/VFThDsiC6n6FG7XWbfA3URg0b3z
xynbsW+f8V3pfH2ji7ntw8HekUWaoej7ha5435giu94A/yInmYTIMNlTLj57TfyT
RSGwttASU7h6x3YFLI5VTuHpcB0GMR4quyxibxmtxUAtFGF0PLYY9nsgVGZ7gOKg
N+9OjN3H709pphN+Qj0XbduMSpp4A/87i4XxxEycFmp6O1p9voecesjAfFydAmd4
ZXK11Is0/WjhpbmNIr7RgPv89uSZKZ8V3XJNk4C16NcBgFeBsidxiqg/GEfimMwa
rpR1AE1ZUdlM6Y8kK66gNiovVYFJitxxupOuiHfsZ5yS2BJb2VUrf/hZmTifsBv3
Ds2eA7zQn33SXR/8GUQUxG96TY8EYVI69JJk6eY+WRBTXg6lgJSegwc9bjrDyNlQ
hhg0w2cJ8qAZpq+7RYb43Dinc7wS+dQorW+9oNARNycMTr7BiJwIgxjcGnyqXDV8
SyiKPz7bowVU/tpY+ZoExq96rGoHMxUC9ZhUylz6e/8uGq5YOjRhMexEBKI5bQX1
I3PH6T9AHqKc5oKJYM6DvEsTrllcEKUd9+0IFgRjmik4uflzThvUuRJl3dO5Qz9u
HhD4pv70sfWjESpLCbkxWH2WQmdBFp3y2fV0aNZOlo28BYsDIZI4oRet548KIkU9
BCL148I7HNTprgg1HbDRoBYXyJ5PypKdwKtEvYqDlMK93bGEk+iRer1nLVBkvICZ
Gr6FRSUsqeGB+90ZhZ9kgzTGLuPXPdH2+IL9xAgvCmqMHtO0yJOIrSv0fQ4oxxtr
mLadIUfIqKkU80I31ZZjZIR+kpFZvZa4Zw7AWYlxYABeZ2wHJoRh2xDif6MbB1tX
k5uUYvEE/633hmITh9DqO+97WBty8bYE4xPqTT/jF9NprWFIONKNXAW/jbRJr5hX
0C7qbtHmghgt+1O+eHBCgQNXCK9GAFnex/KqA+GwPeOvWLT2zfk1GXWzf7CLxlxB
esG9TtFMdIkDshjhVXeq7jnm5b8khjQD+Kxl/q+0gV+IeW2DNWNElddgulc7BQJ1
1L6sh/7h0PVTn6VhYS62w1jSsd3l2bCZlN/2djTs2Z5kYMMgybb1ndB0wRvLtc1w
8f5w8ig6SPWhHKqdOg2trJVUnut33Gu9VgWr5yiGqCPC83Fvi3eHEnRqiXOdgKLY
ombEq1vvbqjkspN/QuG6zr0DrFc3cICSDlze+DFb04M9uxbkkvCE5kVNEbtxpdgM
bN071SrYEyWbAiq4AeipaLX7b514w5oV5cq77NyOh91Es4kkJLcrqIfbf7QBC1n1
QnR7xLRc2Z4/svbkHE6QyvhmVVh0rSeXi9Pfx5BvrP3DGJaTwSQP5Y72dMXSQ1KT
uZnFzfXVFi9BXBWcW5P8fu+ILC+czqV92tv4z+94nMTeOAS7Az+lMyFtmIDjecNo
GaNHEM9N/+g6B6wgjesXyNnMMjF9vAcCi7YZM3rJbb42zTGFJUsF6VlfJ/6Br9bX
TZASNRETtXqvlvx2WhfH0CJTVcpyOchbS6rOKpbrIHHPuf0gkDFI7eaZPbl8W8vw
FW/Qg2eoo42ldmvdINRVpB/Fic10iRoZ0LLIffkNj20MDXWzk+xl2PDbXzNoYFIs
B9zExzENp11YuUg0mRN6RU6nQM/E+zTKCNP6HMR5VZU7enSFA/BVwBKqZf8vKn7a
nWojXkAxO6jGP5oN+mWwskkrMALCMlW0CAJWYb0hnTzI7mTrk2FVw3h1u2yQg/zh
ketV2+XE7jUd0Pt2A2BqKEwrHOnB6AB2OHgA90+6pFsvxjYlwx2a6MiZaey2F8cn
ojrP4jLSdsxBq4cS+3P0LdTadHQ7a3RVsUjIuT3Jj4EYqZh8wTDbgu50aokIQpRN
xGkMrH63yP9UpwgeqCOJS8zi392P4q5mgqVS54XYTR/mlpr7atBrsMl9lJ9F4dHP
T0hbitmBesoYOVIocIFKWDB1jLnTM23I5V9bD+4WCe6LUu60rPOP2MNxpT+Zqvvv
24dBTAgJ/0EmFHCil2fOK5MzrkkN2vnvSb86H1qiYQY0eR5FlX8FemrikCqEX29u
Epy2tIThg/X05gYGz0xQWKsIexUObRx+hcVFCJKT8Yv0whCUg/YpSZSPFCJ1FNqb
4KCM9tZCGjG70ZkvA/X3c9KGZ4coL3qpAyX5m9qrl7BM+64NxoCjQAddvwRqcfwF
ITJK4V1LeWP9gh1UyoeqszIy1+SlUtU/zdGTCYEQJtZcOmIIYR6dV7gve5vpp1Ib
U91MkjTbIPOSC35OpzlllBtmUUD9sehM7aAptmyHzTtpS8Ya4PWL0QC4R2kzRc0Q
p0SviRR5BSEjQtm92qvh4/Vvuh1/ELwDNofu71pr4Y1uig+w+XYIkwDFuxR/6KHk
vfUQqhX87v0qMdjvbKfrmvHWv+yYS4wfApDPIivFFQCOvoe2uqf6c+mF0VXjgzhJ
7DWpRNvcqFV35uVGUw85c3vGB3JcIFYyCS8ccJjiTdIxKWD9jG4zXOnffjkNqvQG
aSfWvIsfHX+IbGa9+MmeP3S6Urfb8doEfzTVlm8dNAWizX24vioqBKUKfoOS6z0Q
rLnEpzRZN1gfdvjAs8ioQWwLZksaAwqPj6hETpv1sVhfff3nLpWCChevDzGqwnww
3bxBAgiIjVLo+NMwIpN8y/mOw12tCoIC/aUf1o9lRL0zW84Ymj8iGy3yHdugL6AH
aHVcZ8GsYk++pIr88OWufQsg17m5TsntZEKFP7mwNmARJnqPx33AuY4P3+/6PcL4
FO/mNPus6LQ2cZxlEfjVkSra9+cJkC8XnWNieh8OmYWs4jr9j4CZikq2hHWlGvKd
8n9AwUA7yXc7/5S6ZGUZBXfTl9V6o9IBmLa1Gv5l21bernXs7uEdvQoaxA6GTJol
SRSR0kdG7luU5bGwCa6LETlooO1sZf9iV4pwFFSiFo7X+l8H4bbQiGWYHEUd2+1p
lmm2kyJzA+HdCejcPh8poSE/m+FIPR+AOqsp1g6vQCN3Oe0y7Hnrak65aU0qtY74
YbjHwmYnzhzhi7Dslz9+op5NP7Ym62PuVWG+hzmlcJZwwK8ZX7Er8bKYDIz4p4dH
fkshSTfWZPxNN1t74pnXNnuXCPKixBQZA4AtX8QGMZpmIAOWI/SVCE+jntWmYb6p
XUN33reLbeHbQFga7/Fc0+xI8jaQEQbU0tSQdUhhrUxOefjYa1r2rRlTBWCdiaSv
Aiy2vJ5pS3KDnoZkFJhNFkqX2h9oGp3+948StR/6zkKbgp60pXsH2auaKAZ6mUPt
gSX4DFndQn+LeDsVrnXbSzZPTA/ZpjWm/0+FVqloPdqZoBp4lkHHHlkmjwm1O7Ey
IOAgkaBQBOirZsZLX5WrsusbAoWRTbGZBukKTKzO3WqivNSl9EcveYJx66oxQAkh
gtLPqObBw4pdqmIYJTYLQd0IayfTvInZM5IxuyrAJjZ3hwTaUb4nYicpayCice7r
pks3GGmAITdhCp4o9fJV7Enrpdux01/QQ3kV/7NwnM6v5COtgqi5QlGnnxA+Es3V
WsetxKwBQFn/e5sqxMNR1WCDeYwZf3xqMDLGdezHNlU72EGGss1YIMES/ycReD06
XCNEqQmAwXk8tgNaOWhw0b4RdLdiA+y5evnE19YVP07sK2TcFvOSUFqYxDx4mGVN
KHSw0DUbtSNubZ/Xv9qN5QnBiN4Q101fRuVDLvV3xLxKC5wXQQyK+ryyZte6D9/i
tKch0ug6maD3D2AWv79A43MPIUHl+Vd0REjPJvqIPY9KsEPBS15LA2N1lNtAeTy/
ZyUDc7aabk+yiy2NLbeTB4YTGhqJBBKbVNwBobZxuP2azaA35F64pa6q4b/VNNO4
R0dEyCLy1HS8soWD9gyNebtK1RBaO727Sa8jF1sSwAdYm71E7wE61X8vbeoiwk6c
yI+JgSDe++g+TyvrUW9ix6xIktVQkkPAsI7LvRrqRsVNdcA9OH3eGikWQaNSBDHL
zViKdPoMwwmjQUJ+pyEgxQHeAHDP7dLeUX3+aotH3KScEkBDM2xH5SQ9gFm+VGmv
Skb6xM9YSu82gDR1o13jZX9/J/AwIIEOz0sywSleSD4/5oPwbqQvMVx/Fp5QeWED
dYxlmV7mXYm+A7oLgE7C4Vc7o7y565qpTAoHp7yYpd2stIJpvFlCuFk4h83bvKwy
q5eXW8IC1OQAcZVDX8SweNnQdmJLgCQ3fphFbztkP43z2aCXP4bwF44SYMVT4q9I
KwjGsOpRfChDTqD61gY8vneYMAFoBN2fKzvq1L6UEUGdFv836PUmJ2fRdwUWtpWk
WJ+mEHmpw0ZroNDuf1Kjq/HxaRkYtw4b2Yzdkmx4ktRepoDAR+fYj/JcByx6VntX
zqSxIJnSOttZlbZhOVAedClqUBrp+BSmFpjav+UIb8ARVGUiRh1ZR+LU/K05QEAm
ET2FB4r0iyJvBNV8apVDrO2kxlNXzrqvDKrrhRPT6tV+Z+uzWUs0gHJmak95RemT
mkpIcenBhbCwOSYLtz1wCBJVeiZmfiTjixuUu/mBBOTei5cB9i1LkK1h/Kbp+0FG
erSrq7dezUnbvx+ZefEKCUDOu8SDIiwYpKHAGC3ozSGpl+x6te5mA1ym9sgcAGJI
0jQKmd9SD2QoAm+iHrrKjmL43Rg7KCbATxiu3/QcsCEPufWLwn3tlRWyTUIB+JMS
5nxgNV54V1Pva1RimIhWmRKWGIBxe5dVeizzAt2icA8rXufkpyyGHgQMANgS26Sa
WMY+a0E4u+sEiOh6uc1GMP8TF4nDAFU1//SCAyCcklSnTBA94+jc13AYYp3CGhRv
UVEumwQWom45bYQLdGhXEn0HnGyW/3Cx2U/88qHRdDZDSxhb9Hgxn49/CV2Sv0Ck
oQiN6NBvXM0A6E3sZVcbuhHW0ZrZYdHoihGnquT0JHWNfb8ugdoIAtfGa9KVhsOL
qWtykY40I4zpmNcDhwZ4WeLvNF0OvizTJWSeOT2zy8Mtt70X2awGErHb19jdXQDd
oA5pb8+BwTJrdgbzCZovzT7IGQIxeEc2mQshwUt+7H/6q+9cSiEcp//fO5fGLdP5
VK89Wl+KcqsZpMSDY/2ktP5wYrv3fVdQFL3FjOeGAkeH37Dp/7uqEExydpWfQEId
dDVhaJBojcKIuRSYttYfUueBuNHYkRK/5MXuW2ngUtxjn/OjEZWzkQxJuoY5Gs9+
kNpvddMTpfanXLstx3dgH1yRiptLWaJIrqpf6YNiDLKebgSXUi0wyGrDO4WafBVV
4aM5AO4eRmG3L9n/7HSsnFBcGwySYs+EDlhYeqiSOukixtaG8nNhmPHo7nPVfhSF
gkQhgpScbh3Od/KGy8RuXXqyfZaxprJAiAGTbjNBupZbi4olieH2MAQ+5YUiFspx
yenY7n6a9+/ERX2eOKIoZOU6XrAS/IqcM68VWB4GxS0ZXQispILpOb9zEqp5ghKu
dY3wVDWNT5boilzazghGuqcoFEJ1KTW8lxnCgUaSbjWLcQLutJZNiLi05f2wB97V
0Ceax8aJ4ZBVo8hQXsZmYw/9NT+ta34DzlwStadKQTSYSqU6Q5L1moNrGw2IF/FV
yfKu700W8rTh8sRlI2XT6ADNSxi2VsWPN//1KnzUR/9S1DawgulZCBZVKLiNJgqv
hnkdFVp0yxugQ1xwxrJj+M1TtLKcQk0o0zgQkdDFWWU3A1QgXWW7u7p1yXsEzHAt
fuasU9OJfRxKsO1Bc/EW1Cboj4uQUbdAbsm80uAyiAolpj9Lihg8iCG60c3oQTaQ
DwzrNoAj+VKl/GWQZqIHvMWloIenMd0fk+0d6rla/sRc+JGbLB2LhSLu8tLgR2k1
Hdkj5PynlN/AAjOhnohX8K7EcAZhMchzfPYaZ5PGJRFY1hcQJgwYFE1CPz3RSnlk
5FE6YFnwUFcC3eAS+W+xIcdkAL/S+O8Rx/R3VA+8TYAe1xvMk+pPg+GEeDcTSTae
hxy1JJMhruRXF1VgUVI+CbTmnZMTXfXPo7FzBQxqoSzD8SzwJphT+uUD/r4ZJu0J
R6Sfvyc4HqSAAL2XyNrNDjE6Ou+4d0qjU/Eay+xnjO3QHFADqyldKvVHinoLfDm+
aWIEpR5lNBPObbxJQcJNb7E0WEZJnKHb+J6LjPQONxtumYD1UB1BQMBLrwniovpM
K5bvbu5Ejz1LYn9b+JBZbJCtyXplwm0Wb3WbUYsv4WLNZ7QfMpQ0Tl7mLnNqdHOz
pCWW+az/9wGnvBcWQJuqYa7WbEwJkOC44Gw1ua97PHbclIcIxTApDNxuG9HAGBlv
SaleSTBOwU4cdMoKCnVwmJzeydyMxuV9cJ/RPfm9w449LHEzsqH4lA659APl8mNB
fVwLvhG82cPbqcnBrwFV6RurSDLpljIEIkW3H8no6DSa7aUsEMMUsdizrYk17Txc
kg5NZF+Fr1EvTdaL4bTEfXY6ym2oMMjVsfQHtOzHtRbN7yw8OsjCc+xNQ14yq0JA
uHxYh+lKedVXTakKRC7XLPuVflQxI8yaxsPoEKED6vRgai5hZWtsvvuHAazQL2cI
l5c8zVo8OefnQq1d/flXiYr1/LRjb/n7T4LtzBZ8RNqykvAsNWvpcvRsBDulG5JH
M9clQElLb1pJiDDQuwgPxOm9xjPyFM06f4ftfqd0UDJ0bF2GrvYIUNkfp7s+9q3u
BmF696CmSFttU+vNuvDdKgJqXfJTgfWwC6TwPAfCycXMJRSDHejyGE2uUTzv8LcG
XIKAg7AVKh5OsVVsALVaMpUw2csb6uyPy2dRo2qj85XUfTSygD7dM4arrpBuFuUN
SDTloZSDLYUhuepwM9+gt3oZGatFJZTjp39s4dXaxd2OkDn+nKBth4fEw3kLJiUD
NhS4VuuQJ6SgfNeVDM5WCRZ6bQfpG0IOLsGghUbln5gV3BJ0DzY4MlleJVm7sngE
jUSpCKinYhc7YV7HPhfAUQ4jPvliIdZa3E5DwcJPUiu3yIuslnmP0qfZv3Fgh3AB
mKfdR8YRGdB99jWXg441MfIUlCTL/KBKoBrvp+PuS9b+v8YRcDkJIf3AV47vO9eG
TmhYA3s/wPMZDxvVX1ygmPrg/nvdEbZICL3WhBU4BUeSOwn7pWeaj//XbnCwVMDQ
v1VVjd77xfnea/j12vbGpqyNTAn5ZrpNoNykMvshHYM5MTplHj5Mgh2ZfDaPKX8z
CecpfSl5oN0nfMmxYmsRXXFEeC5z6HzWjlcX+wViQEjR6azDCl5E0Z1ys19YmHzc
qCMWaL0WchYsMKFjL0fc1v9OgBU4Gwu53xotOBoX7GPIbrVegtp06RxuFpE47jmU
oGGmVc0B4SfKHmK04wt2vngnfIB+/6uoFXwgtXG91RZ5eCsRsoAIolTFrbd1d7PM
55VZEJdOCyGRHI2YI/itOQL/H1n5AU9FmRj/6DRZMXH2WzjBm2HplVxRBQ1xW9Dc
7BqD+jtNlN1PliwGEOK0ysJOHF082gviEMDx2m6q3q1NJxk28K46cpW/1HE7I139
cNzP5qhaSM6VanIyxx3UCyLD67ABJQYtdQ5GqeQm9cYbDZTmFND+NMDEqTLlkQox
I5OKTSJb/4uuFLh1Ftkv9K+uyORTKpIvi6iopRCuxPnmdjLaxU8nVtWEiZSbBCi/
AGCSTheKRgvkk3SXCXCCrBAQKmevsYoWl1OsJOG/mICtMU1BabV12/21TURM8hzF
esgCmqPfpAy2JAvY6PlbIZPs8x6dVC1LJa3w6sKOR3a5d6+MP4GiXmfUcrmMptq3
OHmRlAQoaYeYATjNIxphZjgcEA3Bt70NcouWx1NTLiT4vjLOKsLcEcEZHYq6rmhE
DgILQVloYBsjDXyt6efDiVcCZWzojQ4booLsTsURSUE/PCITsj2rBVEBX9OCLpuI
zyZiE56umAsWLVD0c7axQjJxKVptXD4heqKg7nfW2sjgIIMABum0+3KGYiMUGiCE
gjKO+UAiWUW2+VZXmNScAuJ5LNXWzdipKWX5PVEHfYDc2sDSTuKIbnVfUZCIGXyu
CLAyEtYxihMrSZa6SWP/x0svedoKPdFFykg1qlItt41kmHcMfPMyD9YcIoQOBqcE
ha9uEEqKWjR6gkiSJoKyG9EpGszOy0jWSc0VIQLELNI82Nej8sldimOKXLog720T
6ZGMgJ3VxQiaResVhtXD9QwsWF1cifS/wG3pDbwybYJosJAOmZx2aFMu/8WxZmtD
PchsxWCCYsARYEf85sSwm8vYjf6XmAkM9AISgX05uKxVRUkAc04xScox0/ucxZWC
0ph45/S7d7RvNDUIC+o+v73vzGh5Rwqc1N66TMPoCazbyZGNU5Rp3NUwShIEaUWR
TlMVPNhnNDtZYOn9giogWFu/0VI5M8KgSAlQi6iQ0pGAooAjfbzbQk+i4FCHy/eX
4RoSdQ5IIQPsBCPSCoAX7Nn/jx3tRZB3h89CalgG4z8C4nsTeByZ1RJ81Bl2AEc8
VwR0ArP8tFB943PrroyiJtL4pn9gPL2OFZ2ekj2AZ7hGfxwpljFszu03N5bk+ls6
C6bHpou/dhQQk5vxWB5PVd/cH3AOCKLnp7IE1WujQB8Xd8eKHmTT2Xok8Vaw8iA4
tep322KMFjMxQ0KzN/AYb+0qHxMgrcDrY38qPSEgE496v+bvYNqnUoCAJLi7mjxt
+VkOmsF8d+KuYQ9TUsVjEr2sP/qyenQpFtAr7fJXz7UXbFtROxCgzghmwZ+H97J6
b4bXmkl0ktGMaVjU40vNZZVUOk86/WJu+tUKdzO+jEEqEuvSSjxqO4790wiHi2M3
nMzUfcjCX8VIpgS7H9OGRZztNFdB2U2Sw75nO1/RX222aUDFXMNq7k1LTjEWB0cl
T/duXnYUISzFr6WivwqHNsxMnu4wIOpiK89cfm5Avye0+jyTSZ7tf80nca4N4H+8
cXmpn9Aoifc5G28Vhb9qWJb/ZN4CfVZOKJOsPGykVGwskDq2CfPsDDPd/ruAbhBy
bcbrzlkPIJd0An4QHTHuJukm4QrulOya6hNMHP1DjNKh8ZZxHBN9Zx+foV3B5Dw8
ocCETZy0i6uMA6CS75AxR/kIE/KbVN2NCj4/6Wfy8f9R6UOJoPmtphPDloJAS/hQ
9qKGUifsPBg+T7Fa1xfF65FFlsXuwZfr+wzFL9XBbdmD9opyb3WxQAFWkW2fJ5O7
lnZuSQMZCuzHciJvkmrVedyw2KjRX5KWhozWPuRN5irQ+VyJtaVDQDOaGapuNF4j
m/x8W0+lIpGUjQe8dgpFiUl+ziexuCu0fEXvm+wIChBueAWOvpse1yXdfhxDYnhC
zyQT0dOrbQ6C38pQyhMFjVSAhlKPVMRjFzHg4fIxe0aEslhPRI0Vzyx2r7hMhDav
7zhXlo5MDy9wUbIXKaE5gdcU1zREN9SzXpj77cDcu3bRqc4oF9QXNwa7m//lQ+L/
QJURpOP+qmw9zIk8+ENoJgy+uVjCchEebPzsqOR8uTZk2MIpwey6X7ZxBP7ybt1q
vhJntjY60HdmE7ReJy/AWvhBTGH51yUVPvclFFYWwmXA89/6F1Hk0f4yWBzwuIvQ
agBEbqXj3ix1tlNMJOhYWbRcMAW+OBGqy8YSX9CLY5DA7RbNScruPT895ZZh34Fq
01pLzZJJs050VzmG9SQsW+zrI55XR1FZ4LE3cHTRbIw/nbD+KS2TFKBIgaDEcl+w
ytvkpoTYB+huQOW/0PmG7hqdgEjOh1grb7r55l+68sSU6+HqXUy+lvu3EAEnBMPP
cBMc+VaVTRsrPvnLgj7tTqopmBTx01gZhTa1XBfL3oITY5DWohxuUnx3J8ES96F7
2W8zQOr+3GugjelFmt8vPq1G/reQe0F+5ANLrX6fSYSct4jXDiC2WLEb5ueZDeL5
+9s051n6KcYGq4dgiFMUAg+zXopvqVOty3MmYO7nKvwcLCajEyeycU4xqUPW8nfX
UuCi4pLF0cCs3ivKQ08XUOcUf1aw6vGTtBdWB05b/9ecosk03uMS4OY10YYO+G+q
kXxAFEcL3Niru7Lwqn55ZscrAlD5dSo+bHe8sudstn75+3pCRBRbomjak9tp8XLK
e8s61tN7Lm19TH1UgyuC7dvgWiEoHH/QUxXYfmh/zBoaoV6DYFWhR+3Ktw8lvOrK
ek44JKBpFt8lQy6Quf9tJxV5BCG3aQ3Gwlj9ETYGCkTkqjNV3vwU4STgw0qpwAxd
Pv6R4VBoNgDaGJpnccz+blac+BiPMm7UEoc59gjAsIwQ8EF+U0kvTCTeTEO5EToe
R5VAf/rs1xh9/0aortt9E97OEmyWLIQPXxY9ODPJMCR+WTowNovUGBkeX/yVkB30
cJd204ETo/6YspBD437lCJgrUKBdePKl+UcWeiXWQI2I0M5gI2EK/3aQ4BhlhCVm
4dZADIehvjsObG3ogRxA+aOqB3adSVKAFDlwgIyTFQQfM4GPKhoI/A8V6pQDekn7
SDsuLdd34YZw3uE3O5vPp5tybRjIWtBgfYEHh15xCcTbpIzrIs+V/USLabOjE1LZ
Pj+hOb5jUAoG8F9o2jPhiSPkJq5SDIuJeZybIJKVRFOmM1WWFiDT54YpphEPzOgR
uaLwY/p6/rftPmlPa65gvnqXa0gT82TJAm0puYLn1jdLg313bXGHGDpX9ld5IyfU
Sn2vg4RswbxkqbmYtAGJx5YhqcloP95SI52MUiaiH5xIASLjUxrZ4+PGO8HEmE7l
/mgGDTCir9VihFFeGyPr07z04aZgeArSI4RLkQvmNCcumXLsp8wj695aNCDmOY1g
LbSOml4YmPO9HjE3znFDqwJiuUlxDeJ2gdQ0DUAgC38HXM/u3vNzZfAxiItaz088
zVVyaHhPMFRrKbWF8GS9IyJbB8qKjjAAvQTMiB+VGQMhHSCYiffbmzXNFPxCpfR3
ELhS3TZ3QTDOBOHuyB58+N+8Kejjsbx5hf0mjApD54RrMHAdeFjJYu01t7SQzpY2
fpbwh6x6zERqLwhGRBoTNRQM37ecRklm/c9OKfhBW3M49Ntzt7dGN0n4Cxnk7YEC
yk7bNg7aTmcDURXh2apU6aYkXyIGoRAfur5UIeLjKZ3BKsNQWOCfaLD6QgmqNDp1
Wq47ghcAu7+5qKK9bTHWxBPEG1eopYJn93O+ee9a6R8mGcLq0RRrJmO6JgBkr3PX
4GMDQLlcP8x21T7H94y9KQGvjZ9uzPWwj1GeVYoMtURdsf/jjSiWRiSewZT/ezvJ
FlzhVqrcb6I7gh1BfCcyON3fFCO9rrDRUQYYFBeoTl06vbqa4oJYj2D7zano+DXq
1w4GYihHVUxk6+OrUrWrk80glT55HR3csQGH8PBOn+0qzdpbIlrYNk0vqyBItaPu
/RWnRncf+v0O5bNCAsX++fFrhbS7xutfDdd48NSBcoIQm7TqjPKrp8qjkDlC17wT
sf2PWMwy2HAhFvnK3k0mCwcprOC6V6wHC9PGbjxW5fQzcDZq62mvIamIH6E5OfMh
RqbxeF/lkMp+2IaUNUrKJXGHW75F5fLcPFHGWGTh8hWHVRtJaUNJ/qkwUBgx38M0
1Cak5v2y4srbh/1fKyzW5V9B3LqH6iulHyAxt66O6gAEYlNJucoUvKQDV3o1mKsI
cX4UWAB+ogD5S96Uw6ogXxf9XSfGQkaaUL+RsAlnE5CRMmuqXAyMKZEtwpLKQo+h
ayCHPk+0uHjX92BsOLxO0VbxVC/BjRTs0dYQqV+F1rwMdpC7oydZKylPdIcHlkUU
CfdXabZr1e7N17NhnpEaiO6nZw31mdenFIwDy15DDt0L0K2XFhCmTK6OJ9+04/pw
hLa9dwJl6MwM/Jad7PwLj8hpkIACDjMMIGj3euW+q5q4WfKBadpIvfR7sABqqQ9+
ny8LUUfPpg9U+cgUKKB5gs6lr7Fx4gz5841qlfRhPNuA7gcwqZVEaMN/3uJm9vId
Eqcj4zHOR1nccELw+ApWzN+zxQPa4Ett9aELqHHDPOU+PIVjOTv/hEzhnXhZP0mP
5fqEYmnrtS2I8EJCJgQaWtFMxPq+tCsf09OIR3OMPyNtDc0jgvAH9YHIdr6Of2Qa
SQPmxtQuO2hI5yCkiBSOHdqJihU4w3auVIneiZsIRAlwabND5rFJ3NWgrZ/G4suS
fKz7iOaErAeDS+oLpjPZQggDhQGntZ2QfeWm9cz0ral5g+dySdTrL8hI8IJTTkuU
yETIl/BctSq8M6Ll0CoHpsoNlPQswFC05b9jiZJxxiTv8GrIJUJswWWCd2UGnFb2
JBuFpQfQsi82hQs+wXK+xIqjDi2s+BOtouvKvJy2hugEvqC927HERdd/3Bh2XT+O
fnY1kTdv5QdErk/6xPWRxKSFBXmCPMLJmPnaZKDBjOyjxwkPtNmItcnk7DFl74lL
aK9MW5RgQRcqALHGL5V0nfDOUpzouCc1DCFM30jbg3LGLf8vr8MPbcJ7Fe8zlTN2
vs02cM/agBa9YH9m/SAjlRPxioliFYLFEibodFn9VMlEuWjIb7/Qmf8JwMaCVtfX
1HvrhT9DX+IxA9XdF47aXUKi9y6M204hRjp5rt3sUeaCLy1/wNTIqc6E11AytNQI
CXCMbbsQUTrZgbJ6PiaMtmcEXh64LHFGOZBLxxXfQNcnW0g+Pv+763Tz99eBUzA1
4et9xRTe+2zyx9IK5uABE56PGbraxFRP64onGdbdn4Q8XVj+vQgLYAh+AFPEdmph
Oup6p+Sw2EZNZRfQgPudGyslKGR5Vxjh6RmD4QRN+tHsXilYytuKQlx0ksku2wwW
e+8D9U/BLjJDQimqxnmQWRXVkao4Vq4jrCIAjSLwnxvDmuJFykvvCg2Pu77bik9H
lCsjxQVAK2sriyh/Zz0Y+Xx6qWWOvv6a7TTrLoESfdcS4eS0Z4Vyrmxx6vkwaHfe
MBqpaAoM95Zn8RfPn9shGWfW57g2AgJhp0rXC0ABo9RWE6OimmHtAj4lrC5+/9Ct
EE6u4m4pHZeZlX+VuaTD0uNf1Br1W7BzSAw0+K8PEXn+gl+EB3Yq2Mnep3TGRBAo
BfnDVWdv/yZWhkL9hvIaZDILGG4jlXXvaWHl+GoLlxw5KovLt/xA2YkUqFFdjiIM
omdj+EtWkFK8uL0AoUii0jmwx58zqTLACr6MQeUuLyHycmyRjULS1n2ocHd9MVXn
abFgoqKMrZQ/AE2nz/FhosJINqRsE/DlL2+kpfK1Vbvp3zYvxsyrEJObyUEQmV6L
vxoRO3PSUQYtil/dTe/eyFftErYD+wekznDMr75g4WblK1KScaiCjlkJeUdR/Lwo
SraBOdEmraZwD72+2G12UU8GzDGvGB0YfkXVvTmoRaTn5RTA0MmScQjfq2BNndWx
iI6g6Uu4shsbVs6rPK29LA6FdOtSYpkDYjobEI3QjXzFCUWu+nAi6Gth7zzLE17n
L+N4rwQfTFpj01o8XZGSkh4r7HjOAbUQrjC/7RSgvuKtNjRqj+GrYXs6BlpiFKgQ
NuQic6WTjHmxd1xHDHxa1fLZkslAcnYF7M2Bfv3mum2DmJotXXYV5lgcsoBVNCVm
4ubfh0ytpR1FTCoyzVbaa4DvMt4osre60S+3nHsGwFIAJUJNJwXLKxnd1z2YungL
73NiQ+wHrk4mcpVd3RyBexGaJo/t4W2aKArghPxNA7G+yh0/W58oYT4o6QxsHlmM
55D6Bt0d7q7YrWRda0q1PDDpbZsHylCDPUjZbH1UoLIC0bt3CZeDurHB0383vbot
DWH44C8zjHYAXJXN3dApXGoLy5WO0Z1j90XflQo76rw/5lzWEm0lYm1XkC64HASb
s61l/Td5qsXnExloINuz3t11JGExzuYAbsmQkcxwzjKATym2rG7oCzCYye7d+s2C
j79bEQDn8j2snt7sQHtZgGD1kHCJMYgXF/xGkqQ+PMzHH5hsPoWOPcJNNjxnvwZ5
Rp9YfCczfQ/a7jRX4I4jrs05ER6zE22yEBkkDZkLvzEzm/AWVLuStMpERfx5sRyY
yTNs/xPtLdGr0hYY528dP0YNr7bd0tRglLpXRmpR8TyWnacLSetSfoyqJZUR7EB/
wKpFsjtYwyx2WbtHx/x4BlMv5d3f3rYPfrMbT8WBvMvodwhL6yGEwvgwPg/z2hwM
Sd3jW8oVifhIMB+oTd7kOsJ7feu9/+R+OJTyKqM8YUapRqZ0vok2Wi8yULFKzIaR
XBvdNIuMjp60EIo9T54zZoXJWSSvNy8E+p446Qih586PPrNKVj0kvGKWI3CP95Nz
4sQ3KskI5y3w+E8ncXKqcQL+LcSm65sf3xB/ypeFVHICeUk8j32UQEXUd9URLCA4
L2ATjG7Zv76EJpVPnYfHthktLZZuabc3U2PSDxWn5ihtPD6pz2Tc6SNlIEMTrA5t
r56L+ObbQbR9lqUveR58s5PigiQJuzHd91aKU0WmC/w/4EGig8LPUFHRFd9E3ZXw
SRde7dp1nPvaroPXccK50BcS8LKVj2JC+yi+igmDEeHjVp/wtv+e47yqc6zaek/q
BustZ9CvMQJdvyoj2VC7wuxBH6LoADLnuZJw+4PriHLIgjSE5IC9Baa5PQNhUJD0
5sxEbxUIKxa4pnmyW/NT5ENZdXCABY/4RwxkhpflAGILEgWNueJuOt7dwOzdyO0x
HOqrEeOPRURvmF6MOHG63BPRNksfcwxHXeWD5s+H9lKB5uw11OgCkELLY1ISN8sD
dHZ9Q7VUCUxpjF9g6W1IA7BV85/QJ39OY20ROLtkVpePIj6SLb88RVmg5NcV3N02
YDQWrJfukuk/Unicfpj1ARtm8Xk/1IIV5kaRfY2OllftEC6pPC3B9m1YSJ9jX4nt
ufIaK86lYG49rRHH9CjJ5/NOmSv4dQohnfXZmPUmr3lES2TAHp4EfhLdbpRG71l3
jD2JScrd/6O0XS7ZR/v/rUlE6P7ncas2aknia5RKOqrq6gogmZpL+HdSDE+e3Q4m
Rpgv9Lik7NbwMYzojaZlDWGV95zLahPa28/WGx9VjBlGPtYqOUcLwO86uphNKjAj
x7NxpD5LU0tXl+34qMApKKCfQNYTD2Dpj5aRsWqc1KYzHHsYFxiMvqWFyLFx4AZO
3+miKmAfiEhQQpnwIQ6qZPabS/SiBSlNGcF0lIcb1ihS9ZLh38ylU9I+VUvugR1f
EbN9pVDAFrSio2wZHZBYXk5D71sY8rxCX0+XbWchJExQ9NWEt9ke6OYj9BVRxXEn
XzHG68fCW4J3SKOUbsuMjKa31VD6L0vIQj4gR59MLa/ZnDf/vESXD/jkFnXRFNoY
BnmSxvylD/MpVz8Afm7k/V0TU8BM5dn7r/qwgTD71a5QCvIxKb577buv3sn4qSYJ
R81Qmm8W0M/FOFg7go7ote2jXBbVqfMSDsmHM5wqAMQ0y3oBFfPt2RNKHUHobnNZ
LKJfKsz1VywW3FCRBEPxrVN/rY+/ZJQ9ry7i7rwFhMLm6ChlsVy6Om8hJ1dMPWFe
k6MdWvQk2wt6zZvnHRU3Cpu4nS7UKFnY6MpQqIyNtRBdK+Tnz6YYOrAjTq47VYN1
jycHM0rGpCSIZIf3mayl+USdqEvsWhgi91XNpzsZZOsevJ+xRXMvzKAPWy0+YhRK
+VMsLVaoTqNQ6kT8vHGP/MBYbgyzf6UCv6dSIt+IYbqJr3wqYRdbh7hk8NQNueQ1
GeGw/eclkHNko2mKsPkq63hbR4h+Fuywudg6RJe8+Od03YucSLIy24SDesbx1JxM
J1iRp1Fu5qhsHxx6ADPGTnd/xkfMj5ibhS/GDPppqwUNncbrl1Wo35jl3hLUGqEk
3AT43cYL1SgqXfWFZiRVHQ3XW8hbFVJ6KmyOAGPVU4TThWJ/Vnw7yC8BXSTZ2rXl
KnzLsR4acDSAkD6g0ISXVmaWZRPVt5I+fxMRskA0ETCrDNM8JON5YycC67rIkkUx
1ZRdNqDDPuEIpeysvL7X8Eh5Rsc+tTCCzyO/U2lH65uTIA8RpknpRn9jZFooBZ76
FqUxfNoisBS3g6Hs6ZTJffs20Dpg4obAAmX/v3HeKNlRz64bLt7w5QmKSz6nhn6P
q2ulGSXsCj3Rm3RJ0Kta5//YLVppvieA/8nVHylhdBw7sG3TFYI8ms41l5UFpLCJ
1wqvkWPeJ4TKhoeSc3UdI0G9GCdiWAvJoItoANsKqpyj0C93y1X/P0G1+/u5SAja
tqsTwT1mSMso2ertC3Cu+VXQ/F8gLo5ljl6r9NynTY/NpWgroTevi9C+aRuwGu6w
JcAF7irnXB33vC45T1Rs3daEGRdFRzgMWjo9/jwLLbOCsRiZGR3AkPlwsNbLSy9t
KY5eLhFkzvvJXpX8Hpufvl0m83JV1xq8qt42B+kJbmb2ELNcnCUipiP+rkJsAOY5
AQOB9bqxHexj6xLmkqXF3WPthYTPcGaASCji3v2h31eXtjCXX7cs+Tadp7a0QbvG
hVcOPkHzxgVxJWCbCmovzEsU2EWkprR4JmKCu2cjxtxdkmyNPJWAheWK0aT+vV3H
kulWm57G9E5GTumSwzjfj9SfRsM1ah9T34s9NbbqsiH2uPYvkp1+E8Q9DcK68J3R
ts87XZmMZBRBg9613NTeb56WJpqISoaE2I/hSCdA5j0miOJTF/TOWLGTXY9fjVdX
Sz3U9c1D05lzXw7LOgFGzvbBzF0eZXhbznWR9ZikkAVtKqmK2qICZRWekqZ8l5po
sgKYKwFPuvMCWafjTzYCP7Jxy0BdgVBze68VMtKH0L5/htQW1TlG/hc8B7/kfccH
xE/JmzPkHYlJp4NPi93JDb+RLEC2MiyF2FLNrgfBz5zQ2DszrBGoG0eAGUbwcG0B
kGYSJUBsDFd4SjXwN4RAKBTDpkQaJXhtuB32abfhX00NH/Mzs9DKtO7c3WhETt3J
l9RwNK3VmV1mAitn/xdZusnvh2Z1kF46KYWVqZYfTDHLCRLxz/rjf33CXBySDFJ0
7uVPfRvjpg5f3zc7fma0/3m224GqIzhPg5Eh6pNrpOy3s1Jx2J6zljIZbDzjlusN
ICqW0qjXwzg/ySCnZbQwqdPsbrzAVqlrtDMaNyU/LFYr2qbYNppSL4TiiMgJr2lZ
U3KQR5FOcAGCJxBXZQmZrAP6Uh/6enN4h1jRfN22YosvAFPL2JYV1McET+m6QJrn
iu8WR22AmfrqK9N81qaoW12qsmNVWPMySC9McZu+Yz4EkuhSSDrtkADMQn0W8XLv
qBroCTK89r6AScgLCBSJIjGLoggu3R5/snp6KyhAp/XNwApRuw28du6qfWni7KK2
xUUEJk7Ff6S/rcMv68rcYWytmT8tRZVy3WdyNDB8mfQ3Gde1VmP9LnkbMWmVLFtv
O1Opu0vaJg0uC6pBk/24q8GzW+bZ2FPc0bNV5DPar0SrqWt2oRO1CI1VT1UuyxY8
KkPsuQtaRg7UBOAZA3cP5zzxZ34CXTodMgbJGh/Vn1Od6Wr7UpHQ3YV6P8uaqUIE
G8swsqqjECdL4mLg3Dg3Alr8Q3xYKCRoJ5ZeuIWOW8F7sHPtdE7V3I9I+Cn+lW0z
nGtBFCkAqjktFgsQUWFHoN9jtyjGS0TDh2+yz+3Cn72nExWYXQBXd5zS3KcCkq7x
jwLuZrEWNfPXg1k5A3vuPjnBiEyoK5I/jjWFfuH/LKoBJgqrNKHkEEjp0zVG+hTU
04yY21sCHU61ovjZZ+LHN92kQjHD2np47OUoJce6Fr2L5gI4PWtOHyulFp+gD5Ea
swNrgnI71adXPCcOoE0n5HMTZrvbS0BICRdz5bGq90ZpSGCM/Uy9jRNFkMUxDKTt
OhmZrQT6DRjWhtSHvYvGhoEGNby72nZdXvtpNP6PdHbNP6XLaPp9GG9Bu4qUJQGP
mzmx1Pup+yktsMcZ9mas+WV5dGU36RWN/nsHhdsenTPA8k7JW1Gyaes2AqXympVc
aFXIx7gterYf56nZoCBtzoWcfguH/x1q/KOiTYKl8rKEI0JIVN2GQz31a1PgsYn+
XHGtJVZo/9vrGFlXcV5kZpYnPR2Z/OzeT/8RPBvZBXhPZ43+GWIlcQnAdstzid29
PbQldcdjPnwoMNeKcEuJfeQGcZWxMg5adVWx/tnPYYmc0a25Nme6qN58Gz+scppM
1TedZ0UfXPM4bC5Jlzs635hYp/T7kBVA4CYuOBgFuJ7Yxfnj43W4p/DQtGLwqQo5
HkqMAVfkw1kP3UqfqjRK/NmGVz70Pqk9loJsLEBFq1Ny3scO/1/0ibZDMagRGW/V
tdqzVMG+AThnhB0m+xsKVA+OBWi0S2LOVkenCI6piLNv+d+vZmYxsjwuW4/dNpbP
HkI00yKTAXJkpZ5FLaLUmOyfx298jtn0fHVhfwHrgDFE7v57IANoSF97erj+VKAQ
vJGZAyuaXFVSgbWtjTSVZK8PJzatI5Noq8KUjEyQdu0Ftfa2sjYIGKomH0tXgjR4
0ZbP7cbRKMs07K9OgzQT02e85KM2CAdIPCwxSN0STZhbZxpJo0U5nS6GsoQBl9gc
Oz9L4EQDY690Slc+RQ8V90TEfkiRnZ02RTDPq3Dm/zCrH2aQKFOFqDhHTu0/A+si
jpJPfpZ6jPe2EdhxsLyzrv9Anxm9WhKDCqoPs5yIEJpcpamr/NHI7QupzgpdaUH5
/iAmbj47sP9oG69hHTBhMjdRX4SEVntL0nuf2jUx6cldSa/ERuktti5ZGpBZvd8i
BGcheuJhOYx+Vn2cbMsR3PLORW0/zbVmK2Q6aGTUTIs2Eg0Fm5aJbOu/B5ZJpkHZ
fD4wCmz4haOe6/a4IvmnfvHb5qQ2zFhXOIBAf2r1bsxmEUZ5pOSiW+Q6PYh/Rzhs
qScgqDEjUrbrOVevLy/PNDxbWMdNc2J+OgsH2XisWR2YCsHXwF98l+ROuXHKiAdR
PowqEI5y40y8NP7ufN3EH8zwyYi61N/+OnRX0WTJ2VqLOAIkMNVTI8wgk5SXewIg
8d1wuOGtbJVyu3jdN2oQOb33rk/jF6xwpYp1BwSldeQrCGQq+sslq6Hf8b1eL773
JvO5dnyaIYoNsgbpLcmKEXnUidxSz1thRxOv4u2iuDKxZsqS7v0NWQ3W7urgQzEA
gRRuPQ7aibL9JSyPzERE9l6NqJZddVzd2s+CUZXBDoyZOYSvT7/yKfdAJyCSZ9LD
Q/ecIi0KPb4plTNtuDe+anWPBQ/fn23e0tg/xtTrfUtk0jICa0wt5xloAWIJ9R8v
fVFpcTcduAIjUNiQKtNGbp9KBahdbkrYXBIsIRs+nTouPtLdif3yUJ0+GV6epKif
iyY2pJAhmIPLrkmPWfXIZfGE+miOTo/8jzy7qVaNjwLrofsn5QO2xlfbV/7MeIF9
wne/QyAbu72F40nBrFf9YrtTTpKzGTBHlkV+8vXquit0xN+henS6si+cXfJVeZkt
E8YQUBPyrK+/3+0qdTy3G3+KqdZ3fcEZvgj6hFxsevkw9mhBIQZlJOncNXmMxgPD
q+HZxZ/6jomcGHtQ18pt74yJ7uRdtJBzYXrrZVfIoM4R4K9btVS8fXtn1kmDsagK
HyT5TNdMExi8v9v3WJkhG3w88CmBqBfo03/fgs+hhm4DytejdbdKsUjVtCAX0RQy
0HDInBxo39R4ZQQ3fIBWcqqeTtkoHs550teM9jEpu5dpjJkGxGMDMNxK3wAqyktC
gVaisZ9KcXXcSkKbAR9sSOSh1atyFcDWgJUC/NE4XVHqpfQ9wFq+ybIsAs299SRh
AKo1sVmiLwlsG7VXo/q1xybtQaIukHpY88fwnqZOZFGQ2vGKmVSaBgGKo3GvB1bi
LXwnyN0/wS+jGgxp/mR519XQaN/sg9BeofXSTN3brpHaV/iWx/fAkV6Wm/QDIOws
mUDkaiDyAK3Zv4yiGu3f++z7fH7W/UpOCkD7WQJbcLmLRddk4x7j7dFPajE6RcGN
KKQSSwEZ00ALb65StHxPCJoD99SDbfJy3jcaSpUFJVVVvJVVvo6g3fv8FKW8cpX+
3/cIxrvXs+kAjkm7qjoIIlq8x4/a9dJ0SZeMoHD5DH4KC1nEHrujLEf60blYnGxA
qcqXpJRslx/7q+3aNAGCo3EbMM23uHCvC76xyiTORf5cEmpJVBvMLs19vx12fOFr
ri9pnWN2Gj9D1FHdC378p13dURxN65/xB4uFIZfGFp5jBfmRod3QikNz/ckMwR3R
DWtiH2AB+XkntzfTK3mhtluB9kSMts0Ab62naC9zloRYEKqjPyAUOoHVavmivEKa
iMl1/nA0su1wYhJTCrQ14pdp9Msba/XFzXBCJOcvHUWtuMdFXcQht5peTP4KtWJy
9FmPEh/1NpkgtLsPnEEeEpufPEd2GWgLmWLx0d9VEL4Ed2fBGzYiQBUyFxXfAMF8
rRSAtkFvrU09DGIohUWZ5W/tR5F8AxpTSf5QHpgPhwZ6juYDA9NElZq9O/hQ1MqJ
JcgmZvoJ/w4HCS/Ng8C2VJcM88qXMUltrCFjwDZse5Bv3nE+fnkPCH/iYzKw8mmk
i5IXahJCGkiSDBIbSw4t78YxHLb8DUwkq1ts5pg5tk3u9LtnGdU7OhiA49Ebp+Im
cDA2XX/42h+stB3Rx8dIskznPb2DekYz8wocDBq0aO7LAgfTjVJ+X02DtrCp/6Se
S8RBBndSaLCRPhwVOlEtcDMiWTHXg8QXM6/ucsM4IwPtda6wqsRgUfWRAQVqr2L7
VyB4NJVoViPaPDOnF0iDWW7xHASIQtnBRfvb87nJNDVfR4HWR5hcYArygdfsmhpV
/kWsiz2GOgJ3PeSMf7KlVSf10uEnA1YWMH4UP7TMlkN8RfNkBCYB0WYKhjUfAivT
1WED4UHE95WM5t/BQcKH79Am22EXe3MTwCFoQ2TiOU9PWz5k0ITI6nhAf/6t3M/W
NJsZmdQjZfeSd5AxYIufvAT3WSYJIl01t5TZ8RzFGJWBMuOvVKaBWHHLAcKuIbd0
6Cpnp9qM+fVrvrJKXhdAfDqKXr0BSzGK6YggHvteiU6wD+DCb1UNsUuLKBe1PZaX
Zvo1+mhNc1MxDOkOlOdh3/tcgwwXOzM1QJvavD3dcD5e7Uaq71u41N27IqIojtL9
xL5VsfaYtCmhpGx4Z2bloiAmlzjnrXxLtMqzqG/ORa9WNaXWsm5fExaErvvY0+0i
bNWbRTn/JxfwwxCg3gdtLl9qQI2CrWG9y0Jlqv+53hAPwQB1z5fPyn358gK2/Tdv
WYpY6yXiZBdNv1A2u05NTPneenWFsD7r2k/FwMbWkdbs9iPquAfyv73cu3RajC01
6bWuUUEWUEeRQ0UeGLYZTp8gG8PveB8nuKIlHQRsHTNbnODZRjg6CkfWuV4dRw4x
qefE98g4jhBX2nXmI3LCqU540VqG4NxBMA+LezLH+b7EkDyMSi8ALzWmSaQjtv+a
Wnvn1/m3XfF/pK5d4jUPSWGU7Q8NJQ9zG00f/eIJwKITxN+cu4c/MGjlGXZh5d/b
TaSgXP+fye7OMd3BjU3RdoS6a1hoJtuISytc9jK+Alv8L1Jn8SSzPGmDxeT5gNfG
zHTvzUS2KRqLDoi/M07suUltu12LYLcnCwDlipsUIi4pn5L9T5eiGonq6Ukb+d7n
WNey2QGGF3CYSxaKxncnzhbANyXsmkrYIGzSw1x1d0Vs2ogfBts61QA5KuiWAS7w
V+s9O7lLJs3pgAE4zvF0qtCExRfGp1NIYMvEdEVc/1Eb/bjuW93a9P2y5bp5708m
KO0zhpskOoqmf8X+iXP3ZuthxJL2xV0cLgrtamABQVCwbDPhKH9E22fMLkDz0REc
7UarVQmVKKi8HotqV8uaHTzzImuye5/OEe3n4pab+xdO1rXdQ57ZN0HFzE+KvGz3
ERbRQZ1cIqSYHBwfQLU03R6SJv3Tzqu9D4IYyfC/7aniwV3zhNbOcIOg5CK6v5rh
JkWHYPmTYCcyYRYj9cWgJ4g+aSpYrZEv+QzGQiwpZiOe0eBBaCgtJFm/M6Z3o+66
1yylUkrI5lbjVZmVR2nUk51Nwwz1DfDLkCWXvFI7D7i28yBraKGbsvvnRFuPWXsH
BGR9NFjlBrZP5imrYCwdvLR41+WeQ2X12RVNd7Xq1pwPWAiA18aVCp897sRRAW32
dv938oS066Ecq6RqyN+9jYwZq5tpspHuN9SmJKSr/ZfbHs7VHaZcXG6hNEBZQu8G
Decb/JZ/1MNh+cw0GzLlUJGDae/HXbFNmxTi15IsZZVCPg20WOP7BrB0sTL11sMc
bN2+wFRepibB6+dlzOHHofltJZC4+LiAnmaMvt6db8p/dN/QkOaylYVKHKOgfUPB
ANWe22gbZdj6H1LUmTY0aPM9k1jOsQcYvwjNxrGrq9gtsLwkG4QJHYH4/z/5iPcT
Qr3HrlzMujYtZA9J+TPVaJGxy1dSOXKhXTIX/00ydUB52js4CvrhVL3x1JUMgg4W
mNmXE1oXEPSSAVfgWNn+LJ0l3d45hpr0OsHfsXoC+RqKqmq41E83DANRnWTXYQtb
CEQsfgBvP+6kAVxIOXJdeO1xPG1W7EcqopASVaxIcvL88kaEaWTxQ0bMVGAVX5YQ
osj9TMNVfawfPnWsZB6eXSS0frTSPZ//31QaKcokjaLq6JlX1z3QoaiAWbLfZJkG
oSvqrrYBAL+DfqPaPvU34qzDAP35zwcr0PJlv1NxcYZg2ZLNjxo2qdQDRoGlyBWt
v3EfIKjDHOTUY+8j5Uj1KtLII7KtuZ/g0oJdESQc3Pl1uGQL0u5RHUmVU4oOJfA5
DLUKSBV4W2os9QL+qsyKuq5YJInBQGIQOQS2WW6YxJN+LLPK9K5akDaHC6o3lpqQ
lafaag7gRqbuscvzShDh8gER3uL/HMRkWKJ3MEtumHdkLozkbtjdFWOd07c7vGvs
xnuXXjDhdWJ/E41lnMQ+rcFZZzu4G6EbijXMiYbJqRkKuyrRnCmm1kfE7xAATCCE
V/ne5WS52VhEkfMQGS67MTTxlv9NOs1o0kjhzwgxIRxvSY7Z8je9zXDIsClVUMlg
ADthHyK2zed/nsMtsHVewcWL6L1/J5CV43fNAyxE2ujA4duBBDyAJmMVj8WRxtCn
Qrjf0lvVy5DBsqU6jsLxDiOE/1d06poIWIqU5FBbFbukWR+Pym0foXKJJBBRBKA2
xBFdoTCDJNzYJPlvg8lN5c8yj3qJ+vif4zTyKNb0ggYSEdc41Cav6inseEUqcqFw
WZKjGtWFu8e6rE3xKoYHBnrSuNjVlrzHeqZR/ux5mtpzkGeT2C3ymtKU+1tqdPBZ
g/ZyLBkNGuLaWEJeQGBbKvk8ubIOPGm4qD15/UH8wZ2otdNnCYvsACIa/PLXJKB6
Ml9hX0Xqpz+8zdTxiBMHAtZ4i1UfIgSN0QZ2xv2wW6yTPvzscgTygeuXC6Exs+M1
K2GOL/RN/R/g+NQFidPSlk26yqekzfoPFZiTWqCfu0P8gbHuaXzCoRKXmpQtj5Qk
v1EfIdaSFSUQPhXIG7BudavwJIa0xaV0xpzBCYI5STaFU8TgueeFloyjSjeiqOnw
vgZY89a0AA8CrSli8kNf/cSmvRaLvzZMDH1kGU5b63tPoaDeYScdpxyQb3CcyRMS
Wl0e/BAxT03J7EaBmxmoJmu8Vl4ltOVw5JfR5g9LGa6ZLG0ke9Fz7n7h/epBF5Ee
ktqmBCA6apQrdhnqTzi7cdrsXEnCbeTO388HJbOPOI6QvmAoqVd7VzU4RPJHJkC+
L7HRGRKBYN/hd7cJIv2h5Ve6/UQpYYf5cN/T9RlkkzV3WO9qy1cyRt9ZWa/7qDaa
MF4Rp800/bOGbtUvs99oTwEImadUBy/QuhpPzmy8P7rk+D5zMQ4E3dxUCIjAF0/+
ZfSTA/XQf9q6gxkTr/4rUQZJzRFoHBe2UrsHhXDbW9fp6Y3unAt4rDNaxpWqF0X/
3uE+yjSec5IRzCb0HeonNgPC67YivI0Up5aQqK5h/7VV1EvfkSpwnnBKOlkwVKG0
qmjAzosOKyCz2XD95B76NTMH0BogzO9n+m9+lYbLXtROsbHfVZoHQRJx+oqffeN3
Ak6e3UzgkRbU355F8BtVRHMQhX3dE4l017TIRKxM0EFfwAUqVXYZqp/0rHX4rbli
CnReqcbKpLBvpwRSslJf3mBrsk89IHDLN5xgj75PS14eOwG7xhfp2hdTK1hW+Eyx
cgsIWGc+aX04xGu1xbUeSI+L1LlZqq2EoGXlt3pQxn118lTDYWGyFFQLzkpR8f3Y
xIcl5ZYo6GZ1VEAOHsExzVZz0r4RQJJxHNZUItEpd7+zb0tSBZsPPvhnNfXIC9lN
yqcra0g5P3jweLTSefYgOAFPAWITXGFv++iCos/SHzNNaGw3Y5aPd429SK7EKjuA
aJKvAQPjzkEXDKarqaw/MBcaqvQi2XTJOViYhRiGzofygZwAApV32oHqWqZSnnRy
V20WFWB480A495Ih+DVWdq6+5qM2H/4fKD5EYKs9P7JJgD7v+XTaVgXkcQ/VEIBJ
z9s5m5kWCFuUOugblFXTYiy7H5GOKwBpODY9u4J0E302SVNWcjMa4FWMF4DBuBKa
Fsdnpfl3gE3zb9U4FTrXoG1cEhyqJxKHaT8tZ4M1gh+80Bhguvm6/01TwQKsJ1v2
CV4M8DLHZ5SozAHqP0PpYNkwgG+CiyLwfixZD26CyBp6HiLzN+2ajYN1JkdTAxJk
ixi1F1JrnDiB5RmnXOsUzpdbqft8SKL+NO5TVhlTkarBA0kLia4GZmq7nNGkk0aq
E7SuVaYV4qNpOX0km8R/OmPX0CMP33BMQSrCZfM0TjCrLAYl+blYgZuSQhSQscGb
WpoSKI/H1HKFGon8QGC/CIyekMtj6pWVWnPcH7DJ6PZRZSzWZKLfWeGZdaF8bimC
E+CuX4ozKkjuNGnJqIMNSn/I8yiepicJ2k+R0kRg5Kn720tY8q9YQTQqDyH4Wcew
nyy+K/E9c5CkrwLnGEdr+U1zw1FFGFyHQsbyEz817dY2/hCKWc3p/o4EhEnBWHfC
GpFlWMU8uCvWEkyky40Vo/GrskfcLZPlCrWwj/4snaA+XNygkZCGXD2fxqDp1qJZ
2H5yctjqA5IO22jZoE8h3W99lReiuSOKgtMJAPAWG9el6bX2JYcXxB/jshhTTr7I
U53mTTAcQGWvxOQTt2ebJmNZG4BERFa6lXI421idi1ZCw4bH0WUxBWMNp2r7SGc4
fkLJeLaqQqeqRkhzHtq3kkLCbShbuhmb6XJUvY0FC+vz/gHMA7TVHmX0aeY4GP6B
KDrCZPUanu0mP6Jr3bQvG6uS23M5OkU+YDEExhjSrOlueTiNurwXK1xtI/Umk0KF
aMbnpoW6cOqtsVk6Oga/LNxcDOPdeqQqSqnIobKwoubOYO4OuhvJrWR8OpkwCC+i
MHlt0DocQ4jqtavV8UKFT8y1aP7V0GJn0ILB28ACGHGmI6tXv+FOwacJfjUN352q
MQSXvgDLx8zWivQiE+meB4lhpj6bJYakY3FZ5a4S0rKCUj692isi2zaZ2//YkXP4
o9HunNq+2eudHIeMNHsx3b1Wda7HQ8WKhMurw1yjeEK4wj1MVxhRsfYQGXijD8qS
nGvO8K6uK0CGVfXghzsUqPaD6Y7qa5sHR9Gxg+C98qWPU8HRocRJhwiLWuGKa907
qpfTRswALt4DMkvqhqhkhTrBZMF20wh8mWyKELHxoAUMO4tT3O1FhYsezMRC9EqD
DoXEvq2uDZqYZYSp3mb0zNbKt+yr/qhSEozq3T8L3PJUC77+4Ep/D9igS+fAxoA2
wwlFT+yNWGTWba1HRIxtaJWCxvTRhvNY2ZJAVoYv6dOK+IevNk2DxNFrJAM1C8rL
4o/eqSZOG3hogaxb8y6NqijhRRLpU8CkCD7SnZrutLg+Eu0SFxC27FhA15lNOv/a
hpF5JoSKeVxUv9ZjS2DJcQ620PVyOm7T2C7W9SwbFhcP5a519pJBlfUsQSe1Eubx
JCnaJDa3cAkZemYA3/nsicoCxdUEArkEWAEkEnNlarSXJGbFP4lhUx9j8caAyHFc
u2/H24JX2Wz+7L28HviqeHP8BfMvXO/N8LnQuS/grYZAFjmWLHqw60wyiNnIChu1
zn4rGuX4l5xaR3AqAJRSpJyXOADWZ5mNq9m+hCgfuVS1gxnTAKUb7jxmxO/tO1g3
AhJxI5JXvrFQl7jYZCL1FcUlon3NszTcWP9bDiZ3di6F3K94XV0y5rTLDBGPo9sq
h/i1uBBEYBUsv45FCoPEqB5dZWhepBFPRdZYvJWjkqHU6UM3LZKEVZGyj1BB/k1B
5Pc9VssE6dCEUeSP1i8RosJ6i5KeIpDjSOsLf0Rq+hflxQbwqx9lczfiXmJt7b9r
gzecJP2+eDqpgHvUEdmc8KGkQG+5Ee1jEvr7QhFl1e4kVD0AUTYh63TR5n4cATPo
4nU6C+yvRYK+i46P72XIrhGKHaVZAL7lP8L3DLshRYrLqdVJ+2h6I68bqWsTcWNg
Z1TEhCgAkiPP+oNNMQsheyk8hbcCFqztLCdwvF9Y97UixViss8Uxp+b2gLDmH6SI
TY8GFlHL6halow8Uzs5Xwf0krbANQScRa8KhZ6Upipd6cp6VFh+BK8EhUBjNTcYO
xNJr+5Iuy5dd0+powUu8LI+9OUPxuud129o6OnrhwAeKfXtp5pz04Lmgulu8nDp0
Hbfmd9hzh4fEef0AFM2KQRqnWhM5XP2d28NgyueMaeaOXqTOlMnx1Dby6zr4CK1m
sl5q4RS+HPrpxiABP4KysqA/xv5srE9IjARLsvy5e8W2MvmOmYL6ZW4lchH/mv6l
HON1j/0mi14qquPEw5tucSHeeU9rqyHAvnj3RPLkzt2fHrIdG8f91TM1t306lB6N
tI4e1NftWG5ruqSLLGdz4DfZLwC5o0tbOX6lQJtxoV0RMP4pZagtcDCG0cWDWZjb
vnhAj0IsRkmKIsZKyaZ0EMVE9ou612tatLTHgd22L/1G9PnBXWjuGGBSC/9p68z2
kWmUGd06ect8DyIkq9NqbQilNp8ytr+UxE6ZHzx4M4mi2rMcSvDfWIOAcO6+fJmT
gyZwNI6AR6JPU6xIZPhP5Mmn9YY1ZHve73sHKjaUkjFhRxvc4wpGDXmmt963TQSN
bdOaa9+RWMSNIjgz/J6ItlLfiTelaop/cwKdpVpxJ/bvg4fK5OJ583qVClmvpSFx
Y2CjZm8ABJpNyZgRBkZxbLmy061OZHYlILG5WDl4EQGc3j41aZUg/jjjd2D3J9jB
wr4qAX9211o81EF41SR3E5AuRahHxAQRwxtn/bqO9X0VgpzCNwh8SayJ+HUddHrO
8RUr9HuCCYcYduMLbQUlqshnHzCsXXUxKdjUy1BaTP/+EJbpCEost6OtWsrDEBQZ
eJlc26oe83pWp7TkyCbcnezmi0IzzVqNKpRohViQ+Q0TeX2Gj8GakWlmVX9EqU9r
NnaX9cXU0w6x0eotxHmCf5naS57zQAgPbum0j5Bk141F7dQrc+mPH6qd9jaxd7tz
6g3Oy/2/Dm4IKo+2kJtKv+tsIczUcQSJG9up4vCWIXgkq95eRctuNsUlr3GnqVfP
C8a84kkobTX2/XTm0huKYl5ptmYrMLYU6V7/LAXCS/rpryWLX+cs9Pe9AlSUYXJX
WrHHv6oxXi77dNdur3bF0mDhMwmn1zcoNSdRHsoJsdrPuZgKnYR1ib+JXz8n0bAM
ZQ1xKOwISvyk/hmeG/nfz1LGsdgSpzViiWfPnf0ruHP3PSU1qZkLIDPXxo6mrSfc
u4mwIKTzJzr+3FZ5Ue2MG0XiiJOcKxrts59a4pLZ57gTz8bxSvCQ/HqQDeEvwp3R
JvcHqMNZYbj+GfayNJd2caU/B0xBv2Il7MwnpJ+HOIHwDRQOwPHHluez4pqAArbF
0Jya58I3ve8xVYtMc0uWn33+uwJFFsye8+cfrJ5jmIYcrbowgihoShoZHh629WXL
GSZJ01qROfAxXKmGXzg6Aa/DKZoifhpS24atrFIZEGHJLpmaHSxuQcSWi/VD5K6L
xWXxQZMhvhQoEWfrEFSuUMxbNJnGL7IC7A1r34jbpsK7oVWemB+hE9HGj+jmTCW6
9Eu7W33xUq+YX0nfzZblDcezZXHrFhYGEI4DshJ6aBD79zF3EHcgKgVxwYnF8iQn
STydQrdUckjdbk2NFP1P9hdT1aDMc3gGs7kMRIv/RsYRXjOfmYj2vhqYjN1FoT2J
OloNLZlP7VejbnxU/vccaPKJjGTiLvN7W9s37TDWTk91e6ZdmGuBToi48PM9CHSA
eBZ988YCt8pKUCu32eRf7e8XbwO0MklmfY1OyLItmW5/5yZSnuYZTkxqDd6poDgX
0leQZsKgjbN+vTmTcV4jgVYhTNmmuWWST/c6A6XMCLZNMOcB9vazHi3kQ8lrI8nU
wZYAO8oUym9CU3z5/AihQYX02glKSGBDwyJtuHhRA7bm/O2gjhrcVwzetpz2pk2R
gUwYpqksyelHh43mGCmYKEOb8vUPr4XYXSguCpGNMygBL8BYlt4FrTq8qbuZdYmX
pL5y1k+8kuZj/9yfPNAH5KiVqIAuDgZjKBcHB8k6fBEqCxM4/Oy/uxerGll/J9Km
ksSR0axFaHwR+QMw2TaBhl0HWvThvIxrP6Pawre7LDbY7JtU8x/eA0gb9b9QZgd0
3eyOSCvcRW5tcf6yAIRC51Y2Vd6BC474zXPfiu7QpyykJdgmglosZqFLXWjCnGtK
jvkdZ8b+UE5c+R56tYWuN4LPGr6rMZXlvvoD2IWZNqvhGx2N4V4lTrFh/06dIRPj
wi8BxSD1ZkPw4kuXVLQJ9FBwyHR1cqpGiL4Kj4Qep5OAo35+UxNrFHvDdZ8Rl27n
DJ8NEYAGcZXc8XtCvcHHiWSGaGKGRvrm69DQ0+h8etx+j7qvZMyepkmshxHzz5nL
VQKoSrCHG0Eaqu0r9N7e7jDtqV0R7cslVJkvjt5lgqKlhV9nCRqeT532oDiAweK4
VeATliLMxBs1sbsh8hUY66prR0kci6JHa2wgYESmKQFdATj+xuk0dD3ckME4zSGy
vkRt2dvdMDSOn4MNJDV/UOkYMBYWvskz9yK9LQssZdv+ABMF/NKz+lg4MzzGgqE7
NlKEBEVEqYRnbpDDWluVeZg2eRhHEdE9rNkOWikMP3C7jASv1vX7Wo91hAnK+gxg
2AXfSFwfCUvZp4ffcu/xkwTWsI1nNcGiDDlDkF1P/y9sX9EkoAu1PjzKw+HUU9YT
FS/joR7tVx20pn0d7QJFSRlyl+AyQGZcAQqJHUbcstnJVwLMI5O/uR4z+SaTo8Bn
9yVkGZ53cF+8aUbdlnFR2FR3gQgf7qLWpDgbxeQLyQRjVCT9yozlXLbCHzj4JObm
9wvgve9B+qAEPE5jdUDVT9DBkz8T6+QijUIrKlAtgQkiU5wc+tkagMuSNR/AUGjF
zNQn+5+qGqHr6YB8B+B5g8WMf90fyY1x/5lSD+EB8dPzkP/1+q8hgouNBC5tZqtY
e6LD5y2yrIuLknUkQ3wcbRSoWZRWxpUvpccj/VpNdadmu2nlVgHxCnmR6DWdcesq
TAF/iBHyJ/f+KUQba957RwRks6bRngrRE5fkuY3SM2ZNvx0vJRmee6cywL3l6W33
hVnaeLIUH4/Km0DdQI/eol3uyfpt0SRyQ5vJ+wjp8hPXjn2w+ILlgOIkuOfg4qA8
Ov5K6FccLaeydjVkYQTdj6UwP2g5GXZFL87hilzdGHkBCcdR+sTkBCZZGdMaTuWS
y2DIi1BunxkwIIhucrbepad4NJ2tWPwZl8dmwcnLhx1mwGmtE2gqmoslcw6xKu8d
o1r6qdKv9Zq9byfNaEwbjdtjvzj5d9/ch6yha1lX7ga0abZ2r9gWOvBztPATC9po
560DVs4vEal/pxUKUoP7bNgAu0mVIW+ZvQhpf3iIvBzaRkbfcRAnP+Jzrq/+ZB6w
slCIhuCl6U+P6QmKhOJexpA8LYpVRBDkxP4Xlgkj1Y1dxhisyUG/NArElbNHSJnt
Yv8uryTjSC+aXNgbG3B1QAjGDyOPZ2/vuLzRsJ47y8fBu1rr9rfF2590OAIZ56lE
BicJqW6p75Fz5xDSN9JodauDLIab+5o97IQrEl45G+8WJL6RuXPPpnEuSYcCJlzN
LfTGGEb1fB6pX05pKFY2exh0TFFRm3lG7VjkLXsbspgvoQ5EZGa6XTJo32p1N7V8
bI+mOf0t1D2mhDwj9ifP4lJT+vkA4mkPg18ZpE583kXjCVunxKqVBIfskJMOPe+s
InD/0543NsB1VfSXRYsTI5U6+AGK6w7TUD0lAUDha8LiH0jyoEoW9tar7P/X4Nn3
s59ujH4f0CqXEIc+dYwaI0aS7UmXMLVQdSg7yTw7/kZefvyLF4PZcZitrTmrHBNS
3TC5OmXi6Z+oSteL0jJgVIxA4e50hAnQtTHi3coyVnjY7sMA1eDEb49gqdqh8lmP
AXLIaehaVUJMSlXxvFgiReX8qM6wat8iwrU5DrHt07Gu7nqQjGq7H6BuH4srW4J/
t6Wd6eQnVgQXQ/HWaoID1XN31chPcMHP98Yg4VyePNgFCzdfJCp7lxNuh+eYiVoC
uV7qpQ2ATVxQDp+FFt0T0yK8JSnhkMbfygFLzmLEo61KOoa+ATi6m1p3klxxo9wT
ueoA9yZARFsf/7AiojkRAFA+Uz5U0TDB5/cIuzIw3434VsbdUu9mNZUMSb/ewE8d
58P1EX3f+DDgwVZ4lCj7FCuoIDYVAZVZFgMXfD1CVIlGrQc8yAYLQwNV88NOtQmO
lmoIGfSShJ4/9bbnh/c+fuI9qG6VYaFItNQjPLA8pBjGYHw3AB50TZFlv0nE7KF9
X1nAVne7TiVIw800mTepEQcBK7ESLBz8sC6TspGyYR4FQM2S0w7WTRGoQQy9473W
N0atij3Z11CavYb7JHZZbjZXAcldbvhy48DXwS157iWJ5ScZVHV0arHuFkgguCd0
B345TvtNs5uhM45KeeCSCpNyNpx09BTPigCK+qH+d680UETSvmxdjajdrPMtrYMN
phxGj9O6HhlY/f1+pw2nceJzZ4cGXqGuIdsSSvRgw0NvgM71T96VNn0Ipj2zI+5t
WxlFZlsxcnQFK3tbMKJGj/no2Lc0djzYmuBK57u91kjd3xmqI9UdH5bzn/zoJEXx
cBbW2qTFApnMOiwBAJYpyEVpks0KMgh+Da0NkFmjHD4RKroTN1cY0Q6Fq7ZEA9Mg
wj908zvDv4XnV4GHWzWB2RhPawF3mI0fcjBVaMuyT8BR4GAtR8/vXKBwy5WiyrAc
jk3gBKmbRXO0XsGjeYVqSiL7iT+Hz4j6aX2hUeY+1Ngl01cnzInMIoAyRVUlWf2X
e3bejkXMRa+nMSX93T99FV6+l+ZrC3qLmwLoMEBsks9ZDbAb/SN+PfGH0OShZ4Bp
+NzwD6h/mEZeqaZgCzJg01qoT0PZa1BCrblMtd6V68KX5+5eeY9Q3pmKAgJJRLWw
r05QyqqI1P7gBAxeWmnGN0savS0/HAFpskULtcd+jKqkHkq1m4ozmODimVYogcKo
8CQY80je9dXdY3CH79B2Rj5eVGc1MmmZnDNSbwMGUUTqAZrFqxoRl4kEozLI5+qE
pfjqjf1vcxMTcFHd+acJY7GsYNe8fTZa+8pSejDbzW5BKFk2/vNWrrszqyd6zy5B
AhQgRmtH55Itv4MhsG6jNX/F8Cz/kRrFc5/AL23Mwe9uYnjIfGfjXjCl3IxoiJxI
OlQr3wcY3sLch05RgcCc4lesE1G5LVvV69jGExKZvVP1PHdiZmdCbu0q+DTDbPGk
6mjxWPaD4Ybt3pLOS6Bk1mdf2xJdb487hq2Qfx/JP8hFN1xgPvM6Dm9SaPeZsOg5
vPEEoPlEwafFJve6SVPsWFdHn7M+AyuILmzUZcAahjv1fpuUkI7RzAhy7fK+hIxi
sr25u7qCp9Qb0if1sfKsr4z+GvkLO/e1VLE8YHRBvrxPhmAWX36bEoTWzithFj2a
by7BknHeYB/wigTYe3auoehY6U0RRYfnsKJ9xPB1RaET7KXEbXgvgvZVIYDCuQ5r
ydMOKFbQ3/FMMFrJFle/eEiDXd3ZG+BC6Zalzmj3vuTYFgIUnBE59gXNkXLJQ/90
K9MdBr2T7+lugaqkPX44AnrNEgw/sy3/xeeg4gulnUAOUI5OwVzct0r03GlyueQ4
O2jyda8Z0CpTbpBdmhJL+NKQnDDH+oSfzUtemhcT8HLqvIbKuG0SLl6SdE5yeF98
c0R41DMoTDnNzbJqimo7Ga1zPVBd6CNglMNeX8qDPUpQ3Qqs/Bh9QYdGg/hq8dVy
DjDcQIpu+yHEV7YZsNtnQp8ivb4ODlyL8GYIerlijnWVchwbbDKyTyXx4ed4jIQL
y5ebxNEJOaLbcJ7ESo0zZ7QoHmGbUiGfhTGJbFr1WBqYb+MTM5yUtuxWlX6CpJrY
wo4lpf1v9b9hMhg6RRIM2JhgicO8qFXRIAMy3tZ5r6oTKBzbHiRi6I5t50QdBC3C
hNNKqscaPtVRMSc9k3SKSkhl9ilCn5xKOszFa6HscbMfVScL1X+QTPgz9qUf49OT
8D6Jk23FDZTHqGFQYXjFM2xo5CpMsknk0HnvWegJqhyFUFg7I3O3GwVhKI/zAuzd
8W6g8cjSyZ5Ofie+xv5FeHrByyV/6aNKMvANarQzsi5hqV6D1hUOlDY6INAYfOvm
GZlCEmdGcGNEBjGnxpTyn+qXvDJQrPI/fmrgxnlcXtr7fvHXdnXOvyxm9n8X52he
TsBiWhIg714XC4D6NaNncu2MG3lCtW4RfZV6k22egqFUpnoOVAK3C/0/IsJzc/LB
ouWTXic9hyA+vv/t5wevxL9T6LtZrLWvq7NPn6cHTDmsxRpJUJN3iR30aFzuw28Y
qYoRAgbQKqJEPkexTFUPq3q2Et7GbhLfO56teAdEV85XRN5J9Ko5hoN7tEqmwu6w
dXP6kXdN5wuTLHAyiAhD0IyrnzH1eezyAw3secoyYf6z2fAD+NME2vPtYVdRSGDc
gQP5zA/ipiZ8hqqiLirhaMfprgVgg1gSUtEoDFwGNE6hqzGMyAQqyjXfICgmnPjC
DwZNpniRIQfrw9gnqeNYnDeFNa/b7xNYOBUdOpRTT/3HoUEbidU6DWJ81UaHEjcQ
40iP24200JtcvNTurMLl7USTcczE87mBSxAILr0K3YsB3bw05vgU89WDzBOVUD/p
1xmjWXW9sBBj3BHV/c7UHbIgBS0d3bkjtm1PlGlQohYZ59J0V/T8IGA04NL2it4z
8ut7klTXThyPLsdIfAiZkndTid2tL1bjS3oq5l3nf5E2H6E8+l4sjsv/WAddyL/3
e89umEhio1g5v7ixd1iD5hBYtzUMYfzyrmffLN3Kn59IAE1tFbpvE2b6/T4XahN1
PuLqQGqNrz81up1VAe3Joc9mkkYbJi9THk70gfvI/dYVM77KU1pPEowZUJGW5R5K
jDKFsV+YOFiAjBQn3bx1ES3hPIkGIrhfsQjR7dgAUgB+oorlpWKltR1DuiSEnwfB
o88C0ToFOrB0u+unuEfahND1LB6eUAvXFcIqJgTIjX5uY8Ur7RYvLg/G91ql/Vmd
5Z/K1mfLyen86JE657N5ODtTmM3/wrHKrV2IsV8hVmGfp30UavII9HFHOJ+ENgsv
fd1OmjQjiGQvL3ou0/t67iaiYAaxAjfwMHNYalQaVw3nqScW/HilvVvriFHP3aBj
ubHg1BM6kLcqPXVjEy/3JIXiXYQMqWTusaQE30GcppuuaQu6J+LjDriQR9vGNY8b
CWYCj75dZqy7y6wQf2ooZNuJ9HAu/1n5kpEwMXawGYjthdW2CSi+oDKjaqlxNYYv
ZJsi5LK+a+P569Sjbky5kDXPOAzvB5EuSU5jDOKqyhXcvvNOvfizBzqzmjkDCiwh
iuBZfK1NLOR2K3vbKjHvGGTQ/6pFSyP4ypWK7PKU2mpWwXnNqkMxdSrjtWjNL3a1
/2v/0d2Okx7iS7/HTOM6A5Ene7Rsj/SlvV2H/qJuuduI/qRAOBvdpaTv4+WTClCj
GnUjXpFz+5WefahRJO9pLaD1KCZgrrfCiZnND+svqhrDexSrEmBj3uVE/oLyF74m
JYf2Mz/az2mlAFrSI2RCNsOHx0RPsiDj26s9000RXfvmoU1MdSIiD0cL+YWr8+eh
LsRJxPFpBTTUNkmIC3gzvFlf48SfR0X0FEDGD0WurWJMSw0IcJnlvyL9o1q/qqNP
FRnle7aLU2C5ztboWriXJUCwDBJz4l0gybUrOORB/sKxaXJL95FafYDXJC54ZTym
JU/FrA4GLASGd2hKQx0HmEXZm4zeqXsZZCTFDa9XxZTmVwnkWrUu6IPOdfMqlafu
haSRlsgKAL3BwtAPrVRbBb9IuVrYGXk2EQhH3RJd70+w8NZ/JW5mCVhyUGhQiMN7
7KuGanIeC/XO5hr/clBHBE8f5ndLU3C5NmSOkaKHH/wGxqBlG1TX64VcUPDjEVl4
P0KImICCdMY3hEffxkKbdi80qJrhRYps7nqLQ5LAaQzRqSqTxrO/AgItR27H28jO
Jh4z0h64c6CaALsQmbZKTVwtHi+G97t+arn+6y9pvZnAeWAkksosIssaFdTovTXb
xlpID3awAgsQrfF5owuNZwtkLKpfLVAAkylv1wHxF5dEIXBu7n1o/+ellwLtgkgm
+RSLcSXLwciumL5t24L6pSgLPiHQmWuwWY/yh0u5yQB38vvzRo/Yia5IJWE6ThJA
0hnkhS8XzRlgG+CByTnJpHRMBl4Fodv9yLo8KUfsSqOBPQY0gzvM+vD1oH/7NbqM
my3que1P1nw7skKi1777yFt/shKQKsPoudfjClc1oVFcspehQG/usREX+tIt3llT
s6aTo6pMdRDkk4zNXoZqvPyr1CIY5kX5rZm0BzGSiAH/U2wOOjuSfoxUkrjl8k6W
4QT04U5yIwPKxLIO2P6V7k+AaxRkHYDAzQ5hWqPozS4eloZLGq+o/gsiO9QcRs8i
MWaE4+s07GW+rafKcmJYH0HhBLyNC3kGKhuME7WJ2gYqQsYl2CSxd0Z/UXHPD4+F
3oZXH/n6V28d17DAgk01MHf9RyMKorN8ude8hXRrtcuoOtCSZr+qA7YkKrcaqRYV
2DE6b4fRR3GGbRqbODUuwGXGz6uhi1kT1u+glwgCdKelxkGFnBCqsaLtZMYYFZJY
8QwscaSts7ae7CzM/rnACfAwePsONEtbrOeEJfX5P7I6RWirTkXAx0oANaurxzRP
ZiMYLi9qobZ+bnoLoSbuq2WSLSMMP/ZsooMofacynoPTiQB9Eb0VOfLy+wwnySlb
IU4EdA7QkT93vMqelRJNkp5pTMVLTMSamUvX6tLqREuMYl6QAVzMemKvBQC5Bxpd
g8QDyzYQh0eBkFehSH9X5dMCInfUXGxJwa8Fpk1Q7OBLpzTStSwdk52YNpLBYyz8
mgrk/Ig5oVSPRQfDHqOEdmVMX9WWZaBCG5VOOE1FDVuf3npzj6dKqB8jHF8obwws
Ulle3ePSTVSTqO6HJENzEP6nSOQ6BUgDkVmyUZuPVOwmfIXEbC6wnfI11m7XPf/b
2iGjAnLCUow7wzawISGlsAcscvqPU1dK+2iSuSvN1/5/ge6modKj0rDCmXZ3Kyim
rdWw9RMjGSMeRZEm3Wyq02Lwo/zZpVFsLIAhlQpg1xp2+o3u6qardj7Qo1nqUa/n
ZMpOPG3Dse/uEgw67vGIrDLxHdBC0TtAdy+1BESoc7cu4L04bFFaDeiO3QSU7Akv
9qz7Cc3jltPXcbpnZba69YRQ0cl+yk+tJ710gL0LDn/KDB1ASTbVt23xnanxbmdr
s9oQs0vc7SLDjz6D38LlIRnZn3ba1kNpjLvaGURMOn8mw+pE28HoYm+Vgg7t2MZo
dS5HD/j3nwq5fsQn6JV5LUJcX0zXAskmS0H5INuLvZc/fjTuDwQdV3QbjHpv9kf8
J0gAkimPGZF83qk43AcAUd21aMc61KuECUtffCRI12hQiJnMQC5PEeGZkc/0TuFn
ZTVvtYnEUrxv7t8JItEuSBv70I4NNg5WJBxiwGCxdl6/80mbRV7ifN90lmgxS4tC
tGDsA0MrWm1+9/KTX2+UDwNgeO3ASe8jTxlbupUk5p9BYbtT8JolqCUOjfXS9vlk
vb76Zq8ycN6gdIqW3aswYi1/sFP0VjyXjkVesPV/KrFrx4o/+XMjzQ3Pa2puPrtC
ALc97Z0SffJn4AHIDBaWeZb1bMvnBXCj2WX9Qlailw4/NI7PEdguTyserhzIVgSk
LYjSiaCwsJ5qWcdACOpkEXidkol5KgVUI5jpb7BC7/FwlQT3duj7NeCdzNIW41sM
4BlIxkQLh+NWeVBlyVgyfjw5ywdMhvFCWFXL/3I5sCeUXika6389br2Ca7WujPoV
hVtL840j3b2+s6ep5F2CfWMEqNMbTVM2jMUqyiy/6hyENm4MDMDdtHT2wxsWrMQC
LMc48zHwduDpuN9KGJBwdUr1pXEcKqVLFB78mnq+MvMXP4NgE/Z6hapPLkXIBRY0
XclsRojfinzPhmSxsmS0l2od2S7eP2cON9C/kdjyf34lzs++XqShL01GeLIFGfCA
aSERxRd28elb4N8zL5kAa9s+R46PhltM9b2e6oraoRqfn07qj78Mq5kl7CZTmKlk
o0ToRXebrP7tspWKijgVH3K4b1ReXbbFZOzN1qUDZxovWJGmh6txGThV5lLQSxSI
hqYqGBLf8MPGH0SBkxxoXOJuTFmZ7NmQvPjVmk+aV0MrqfX6e31YxE/u3nHc1dVs
sxClNWYemECh5aXlIs/bglIZt0zeca3mAMkviSUYboJTJc86qD+5hmkuzMfR/aL3
bizM46dndnSgEiaQ4AnP1DhK8t+y+A7NgSmJSirXnEpM3vYw6ahXZWDgZMvoWY8t
shdkRhKD+60bSmSyj5ZRtaYYRsHmS4G7u4DKJNwFSDxQotkdpIutkbtfVXQIbSQy
TDU/uwQ6Z/cPLNFkoDVjIQ8JRIlSfeYP8ryIU5fdTJIa//ajVun4YexA+u0inofM
uAEF9RRSkJYafx+87aQt7keY1k9qwOnALuQP9G7IgiyPKrMakR7BJfitWKSTAQB0
EH9AgZWSzAmbGl3WETO+9pll+t/klJDYCOVscf1dtsoVXD6gmmlKkoAogvqc7aqv
xVBaExPF4HH8BYx+VmQbKMXSPteGgbO33Qc0/Y6OFkMgUu52CM4tMsOrcdT+9aie
4hpschA8Yt6ZdiH+rgTvHpCpRTWgV+n9mOMIpkuIgaXDqPgCcK8+Ee+7jQ1Hdp0x
4NzK/zkJEAXk6YqER7plKhrfe18v7J1B1DgnS+RJ+vp0QFXExXY3ScWRtkRTASUm
SFdrH1GVV/Z86bmU1RWcrR3J9XuqjOJPX04UM4oKK1Sqw7agcFV0DR3H1Y3vvLJz
b2oI6e11/n0O9+PFkDfRXcnnkkcrekBBjB/TB40xUXw8Tu2+VyQUAl00YaYBbRdS
f7Zs0GvrBIzxN2CHOlikW8KHXwJj6FsH5Zg3Id4+5QL0n8VbDhK6i2uorkqshsm+
qKOpdO/9oMjipRuhf2cEoAFA4hE3P9+4tGZh+YdfRX0nGMTQ9iXxQuU8wLosxcla
N6QlZ0wFW+W4jxounAhz2Apc5Cdtd93tNmwDZtUwKO02HKX5M4z7T2SyXKD1LsWv
8weMZeTTQRskn8nqcwVjFEkEcDVn4MFLzG833I0eX7UQjgkGoINGZaivsIB9Ry7j
uEdqOovsMYVaWAD61Oh9QFhOZNfCeOWKLbtMzpWm2p2CDw+loBc4vhXK4UHH1BD/
cP8EhRSPuvMi8jMQTcxw+fsU+krJjERzTq61q0UAj2Vw77FglyupG0M5E/FS8fql
gPJP73V+TaCrGs/9TbqvS+4bviK4w26AowrTHfQV1vJAmUmv/b5SI71tKNYw9BLE
oeGuYkBomy1BiOeN4zZ/0Cg9VcMiVw7rfItPStYXTwMkrCTZnYoIlONSBuSGn/Ei
DK5qMPSSdS767KwHbRTWCI0PGccIoX5GvhwZQd3Wem4uUmA4uZitwevz+tBIpaEX
PPD2iIqRWqblfigeeUsycFzc04FNbazXpcJemy11X2gvU93KJFdvmA4oF4hAf5uk
lVI13bajhp3whwZr14IQs6WVz+HtSwQe4EYBp1deSYqkC+Y4NBJiWLU9gX9V3jb6
ffWb3mPVbs74OmIKnE+bwLVJKkA3+S+IFjIKDTrN/zTf0OCbPgsXOFzhPB/Dy1Aa
hKlFvt7cB4M1J64knbOdn8d6jp4f8Xe63MAI0q8EfiKkRJILchpGMT0Sqv/kCAB7
XfiC1uIuvZomdNOO9IbrZu8TbpPTxR6Vq6bUFtctdeU9qJi0tnca63BzwUyf/K8Y
7YFa56R3W/JJsD7sR8Je+GPd+vaJxqDaJ6yrvXjY28b1UOR+ZRyFfcO+RDD+gWN/
5V2nGAI0MXRLwY4Vyu6XZhzwGXP4Vb3P75cosdPpJBAU8czEvST60lOYGUhnp6+W
2DCvCQs1EdTCv7oZ3wcRYUebi6oT2HVL/683eugosImtzQZqowEErDzy63A+w4BZ
bkMgVwI0+INoHog8ELYcG5vogJHXOR4kT9RFNJGTt2to7RQMzVBQj9BrEU4w9UA9
6R/cBfABnL6aWmWJ9DtKjbFMgCHuZjP7fMMR6CcregnIMTXJPWUb9uYE2lqinPei
dDXEq0reSbrPH4v/PIZ8V54hcCfN+L5XWsAfXRvVbRsCeRiXnszOl4VmlvorbQkz
lFSdvUYlo8LfXB6oirS38RDQ0zlGUp3s/tLkzt0xEju4wsQTztdamNGtm3NTZQ8m
jTgq5B3y4ogXs9xQWMbqY2xEnO3523dwRW0nuOjXFFSFIps9U7jPPGpD87L31bIf
9TfASjxxDNLrhKGox9Hn74feHhUyV4zHhUFsbdwYlzBZem3R/tfej2EaeAuRy80a
e/WNh+MC83NvJAxHleps09wzwxvq8F7x6MY09dUOnaEgMlCVv5atsnBNevvYeKFz
Pdb+8ukEL4TTtZjhu5i+uNOdq6/KSmsS2MN19SuvYagehqrk3e042SoGhOBKmZ9E
7lnG3RPV34sjSWserR0zsNJatlFqH+vMejPNVAMD/A23c+P+o8eFiLKe3fg4Z/Qv
TtDnGDbd0xKVWY9Ks9D3NMwvpTepRbWQtRiI/W3qyUgTIeg8GhbZEijuObkVIhXm
iZ9KMZMEWdIIcwxuyEReZj6kY46qN0fYnu7yl45Heu91et577K5g1vSlUCm4I6sJ
f9Uq2zrC737P2j5D5h27acqFrEBGShTxz3X5qKuO/oJuQkWfNZjiB9KnLO0N02vR
1ObKUuWi4Cpcru2R8iVc/jX6thxfk+l3bpRWsh1YANb018CZzWt1FN3gQ1R4GkQr
z8P2zy/QWiFZZK4zEj7IXTaAuveI/lSBnfmW1bXEcmiCrpNCtNdihnvUGh5hpvlF
cX9IUzojKW8bJAQxpVwC+ZpOGSLOUmpPrBLqVUiiweMpJI+I8JvkrBB2oZmwJHNX
t5kk8mUWIXaNMZchdVbVmTkXnWjJZCGXltwDzXX32gtZd2t7q4waTrYBpTdTdnPY
CD9yHUqULYtlJdMSf/ZrVTDVIZiHnMq3BW0mkJOBWfWkw62XwHpA0q1vozXdFUDP
vJrAneACOdzr2F5tEkD5VflcpgY9MgU3gFuKXpyQap2bBYunPz5OhtzzTjJ3pRYx
xenu+vwovPWKE9mRckaIVQVcIU6NXnNH3uxLJIzXMzW4/rmMb7/DfDr+D/6THnnS
iHaXNQb0CqdeBpRM2HdWkbIgJg98MgDx7lLs2mhYcouNFIJuhAPC0clP8OUbEqR6
mHTkJiZszNdf0y+C5YhEbfPENhNcedpPqq0bsgVoS3q7yoFK09erfz514PB+ZU0v
KRx8z8fN0OtDtTCHK2By7Oe8kQb1U5CQqcr29sm+hZUYHVcDZQpsQsvTQv6H5/56
/+cG6Eie7o42fUAQ8cEkCm466rjPkELu5BC19tu9FRkV/5I0yoEXkiLnrhprscnh
qx+ArXrvA5AdHUjrs2E60YDP8UeLTEiTDCFo2aGFs6awcE7WwyBagGbMGGF5BB40
TTlpOxxRg+8G0eid+GL00C6BCawjWf8V3LcdiGMBOUG7pGfKERns9df3XDUDvczJ
55K1v+YRkYpn6HWXrxXlBfC4dkkpr9bkvAUhdn9ibEQOEF6J7hfQ/uxga1dsApW8
7eKKD38vOOdVrr/W3eWPWyMmgezxRFC4jHWXbXkelQd3JhhJatqDw26yLWTCd4hY
dvb1Q57sRGPNJYZgWVmNzUt4qKEEmFaQGryh1Pa1+vQ0SvNcupOG8EMgRdLNrxsR
hZOHiOGarU57esjMyFnSzW1gUI8prdhTnz9zHTOeeLqx1Kqp7aHaS1vq2BNhYTb7
wmx5DTWY4nWVNTH1YnDUjlwZdKP6W9R2GJrPX9z8yYxDvO064+9w/A7dBCBZlMKL
hxmj+BMFWpVspGMwROLU/F+hzfbCY7iqs1LdHFksOq0OIgefM49TqGeTGDqDxEeP
L1lO3vAKY/I7xtK/h8mG1/9mSRGIAc3N2G4nTh8hSHH5asto5eMdc1nSwXPT9MwL
pyqtvDnE/fcmTZHp1UXyr1euPK0so+Qa6bzSafto1PcDRc4IIHfkSlDIHxe6dLBt
J7UxHg1Ysaau49TbvbPBLloaec9VUR3Ndb6YtsIUNPGsUTR05E4BVB4n6dGtB1dn
wSYXaOD7sycPOr/5cs/tcfjXea6qXgNi49jH5uHnMKN5BBR1Q+goKzsfIeJxtILQ
o0s7Wqx9UnS82ljQX5TVnmH3Ysjo8SY7nQRG4oKvyOQJ9ICM58pQl90BAsT3HQPn
6uBD5ZDn3Sr9dJxShq48+KOq9eKCIEHz6fSlB6Ds/hKejpVNtel06L9jPI9nrnSG
rnn2YCoJ5nSA7+6XZoSFSpjeEmq6WpScKYfxKDYq0H/qOTa0Ni2V6w1Gv5XEB2C1
SOIRs6OmUzQAk7V/rXHPN+hOgFDrlIgHXx5HzB5qz2SfSDXZ+hOWpLihnlU3IIJ5
PaYhNVYC2Y3/ywWmHUUZweZjgX7vcKk99ILBB/uedtSFyr+AFWvAYIAzhuLVHTZU
HECYoUxRO/e46G1WDN/FUdrijBMKZ+KBQraP0R3G3NpnilWMiYTk4hdWo0WwGKkr
0LX7zPLO8WjCNICeC20kg3X1j2yco9Bn8sPw5jmjXQs0SEB+NimmBKnqDgY1brmQ
a0N/PkS0A7nG6LhXox/edEistbj+p914JzZ5gikhd/EA8aAuw3+dmu9P7ibhuC1S
kpnq9JLT4sThua/660STCWwMiTyS4WIlcG1bwbzUOKlgKiORkRZuJWY8gP7G+XsD
+K28Rx7NTgA4SxR/o3uY9uMOd4e+51rwkXx++sTNf7fhjRdzzaI+3KtbttcVDHuJ
fCrwk8jzxftLRguugxfKotjPj8bwBNOwtl6OaB/COyea3T1UO7p98QDCyK698gcZ
mU9DoQKLD56xW7ibHtSfdKLEzVXlS5y1nAx8D2/tw2uArRBq5wi9wVcagmzM3edU
PDUOgTYTg3EH+zpprM2r9VlS1InItA9M4G19WpsQz0fKEJlRmxLnLbDTd8Q6rCG6
mYFlELwBNXlsaknEO6SWVnMyky0711LACCVkaJlYJI8WU6rcLrZvW7g3YUvY7l6B
lKDNEMy2orpIGi1DuOVftPSVZVnkEcrEG7MfHgbqKivW0R9GiNKi03DC+0B84tV6
6s5/36Qqr2zJnuEA8jVDzWqorBcGVVQeTJC7Jk73IwC01N8Ze9twR+CFEnMa7hae
M0e9fu6GXeKXfLtfZiJTbM0eKe1bYc5a6Zri6EyXYmGCny2DEviDTf9/QnAlLi7x
U5HhOjxnkSAQllFuXcIBnavO6ukhWC4n9wQ7n0y+uAWWhdajv8EhjAmq5qK1gRjJ
Cxe9uQC3nmhqgkmrUoVB0V0J6+kKVydxIj5HwqdQLMIQPZxj8EQFX5/Od1ljhb5r
5YNnHQ+jU7J0jFNKsmKOJ4WKIlUv2OxDYF8FuM6X/Bz4hIjn9nSl/cG+vrHOrAhD
FfyYCiBfMUOfN86riA8JS6tG3vbZp3sVOFbKB3f0lwb85qOkcgqdOX3vPcAAGCkx
PTH9YxT9XkmXJVdKbBHXMePu12Pc3HPkav0AZWLNkLMngwgdEbPEHmw6Eg78EwUx
nHFZItHBgWekKYGnUn0L1TfdrqQhogp8kWmLY/llV0oZgR+YI4uXDvKqy2aRzkXr
JIQuuifyfPzCWvezz8Ml7b0scMj2llDEFNtCkD4aMZxB3A3fqYJFQaSEdZiAVlYJ
E96vNg4IwOgMLt2QQW1MyiDqN5uWHz4crSSgxeX9YoJAhAkG8FxRu53xVuvjWLD5
pXftZ+CM317GddIlLswKfQn7m9WFK3yh5eTaWKkkiGcNUZtyNiCWiMEAD0a+AhZE
ZF3t7fmC0SXWHB4qqp9Rdd3hL7Q0o0D5k81htBgsg19kWQI+YkwF2fTtTHDNmiGR
TXkKH+uK3/LM2cGtHkCYeCZVQUXByDGs4N636Bv9Gr1rP0RSO7xoHUx8CSxgCmAD
RDqsk5RBJBS7j1QgNMhdXWnwTQQt6V6I/gRPvWFnsxoqwFgZ3Ijk4Xyq37j1pDxw
UpGRuFwno64aRzYd84q/awHyZpYQdRNBc1qfYt4BhLdp2CM5EI+6jl5OYBuRjr99
c1LvJ2/093TUEOnFU4lGc23rPqNaRlaGojPNUILDpQ3PDseq3HBvjjJTIEICqh7h
TSkiqofZB4/TdbhZq0znssxNftEE3hFFHhLUoUfUN7fX2/IuczZUFcJ+XpcQ9iZR
Pk8ijO6aUEQvUpOLg9Zt3G8BJ63UM6Ucj7SBpRbP2PSNjNzRIeM6bar+8grNnIXp
3ivJg1NPQqPNvIIMOZ+y8YkJLAt22WI4jT8yoCMpamRzwX/LV4s00MeoRPKOR8tK
RlewM8p0XOoIWsRkCi3ZvzzvNQwewhcDeJV65F1yQMg6vYcLwS7kIAzzkY9uDL6I
yJuoN2RpFrVZXHPCqHPPfY5iuMY9IyAzs9Hkx/FZ785T/bx11WzE5PIC0+OBAB8y
8fAoViH2GMq7Tbd840+tsBhfiDi+dDuqxNWnq5yfYCnhIZIlOV4uBRszxus3m0PN
LI9gMhi7OH4ihqZ8aAck3CwYxkyJtWmf9OxCvcJ92W6/eF8OV0Ze/szwfEXXZvxJ
qGa3atcWY9HqAcUcjEhQsrVU7HpK7Z3c73OhZYD+vSXkRSXaMTiftnwwLrE2e02N
GoUXOO4GQ9Dw4ky+ediaJbArRt49N/BNoWa0d+8s5nZy4zLXfcguLX3x9aIwIBJd
jWyKU0UZKJ2vU+wfAiMSnQBuN4Efs1KfIaeZzue4PyaChjrgV+FwJ/Z6pnl0/8iK
TvT6sXgwetkdE0pPRO+HbjrtG5DYZyXTqqSttGoMN53EB8BYbP3KSW97CgEJkxHa
uVfHgd1VaMeYujjAUvinj+xeTBYEE74N0ozpQ/Y2hhqGXjAZAg7pDXl3DFORO9WU
BRqcCo48NPY/gjgrO8aNgdYvS9sl4KKfQEgJQd1RhvBr5nC61AL/1DenZZxTN7NX
+jXahNfoo4kOw3i4K7PLLBiXN+4H9JOisRaR3d6JU3ak54QEKuPsYmCa9twmU0+j
lEkoxb7PGmvj/bSuImJEHdpGw+JWBypTWnRK0ud1UTgzhIQ4cHEq1G88IJx6Hqtf
al1ihERTtd3qnEcJV5b4bQMA3TfyYAKD8PxtFrN8mio3tjLmsxCp66E7N12rVXa+
4rQEJmfV/9lmXQd0OqIRw8x8vuu1dWK0zLO+CukyuhGjyDYU7KUlsHeyvhdp0FaT
Uwy4vIxY/ADOLsEK4EZZXgsP9UP3Fxknvbw5zr77PoJpcCfzCpTvor2hjcSVOzDG
NUW+ZDBhiOCUpP9mZm2ecaRQoNQLUqfrv7nIbHmy9XrjevUdKT36Yn10dViDNw9Q
+C7L9xBHPvFlSyxcxjke7/yBFx5IhYJe1e2BpHTpi4GIVJRbF2+qs1E2ToTyuH2u
HDzG5v5U2oB/2e16PCaolCE5hKloaEOmXG22LmDSstm+lvDfsmG5l+i19QbgV4+5
fQXooeXA3AfjEW2cIiLzCQcSnEhQ3stRisJR0ZMCFvjlYRfBHilTpMkFYsxuHWbC
P5G3oH+ZNBflUKJXYhZaY6fovS1Y7LPKgUOe3NWwrp9IYhrI9UFpaejjp/ur3cjd
gEi9k9PYyX3q+sKn4BdqW+py71D1Nk8t5ZrkJcp+JQvxnq5WnfqZ1VzYHxoKtVwe
FYd44Z2HvmRr6J8dbBjsHlogH00jlBPEFccPiUUsXiW5KXfhzBhHmog3zaIMTLJ3
SzqeLeTS4EqSFrWcIwFS8sC/xWPTh7WM64jHZTLONM/g4vjoKIJjsFAfzdv6qJzr
UydKd1FCQa30EBjlT+3OJswldqGiAs7MuK48tM8rnRbPHQXxiM0UxWCG3FolOqw8
wg8Qnf5VxYzS7SJX+qtuAG46la95bR64xTjYS8GaJSmU/5gKhBLuLdp40SruFo5E
yord946JqoEhHwS3kS9YObMwE+FS6XhR4QAlouuLrSYLBT8JlGFKo3t9l4Tb+x8n
WJ+pgUDGAekOlLXCvVEOmplaMa6B/dcb9u21rAQb00imTZcRMkkikCr5XxH2Xn8l
gP/u5AoOn/Lh52UOtekE1n4NjPEkll3oFFOARjU7815EEvGpGV9uk8l5TI97XJy1
EDDABFriwKEB2i/JMxbQHHkLt+QfWO/jEheoUBFfmLtoKP6bHyoDHGBUR11mBAg4
eKwQiqCkUt3vtONP/e9/hdLnmKl6DodzB1qQy/9hF7WqDVydx5FXAnai37JcXEqg
Mp9ArKUoLz1B/I1bxi0gnu8IJ9Cqi+JV1+ihtISnhZ7blxFyxQUagLJZxtECHXBq
dL+FECLbXjQaRcUaEbeM2laJ1ZnWwUzdU/O6c5LDH/Hov04Q7md1hlJiRQ5VNYWc
oh8F7HKfRYGrPylfdFW481zi9kVvgzRiYWUq/9d+bGMgTkJLs/Doe4lNAeQo8rJw
8RGGRpvUm3i0AT4I4UPAwCpFAhVr08lCkbbZkKTMoR+pvjX3i7kyeMyvfF6Q3IRb
Hg59yso6bnT9lywQkK6aRpzKR4z9xCWi/5X3+jmTXN7y2RD8lOIStjdmd16ekDHA
myYYoPzoUhtrjmxRMaTLNhr++uhhuHTezh0mfMd2K4ALCSl06Gbo3m4wicOt9ru6
jZttOOb62XZQhHrNEXx+LN35DE+rk7VeJ8MKkxG7k/scrF7QSslJcxw/oP5/AYWV
TQA3cfRdEQqqmqFxKmUdgenAyqCvdE/Uq7S8x+FaUBv2K/fp/iosOI4AleprbgNv
iaRfsiFpPW7JFX6zGzIh+196UGm6vUDyWUli9YFH4doykuQ6GfCLzA/gXUQTo29m
WJ7cbtIfkXg8zEc53+MV4rbJOjQnN5Cs+cKlHe4U3ecTaomZ86izudYHrbDHRYR3
cONKOWm22UV+0D2DnrYne5HlkmgS50Bx52NWsf9ijr57YfZFVkMP0YXomT6PHGyN
RXI5Qxg4I+l4XQ8V2zkt27jZ2Q19AW4vj0ktGsCu46PaJN5rk5nfJSFjOzCJu0+D
2wzz5ndxAkVpOD5p3G/nOC1rkxUqrzVD9g6KCccAni0+vJhNPNfxRJwa0ed6Jk6C
aZ2ltGOCE9S5YcLw2xLqk00nKkhyNpZnfUKMi8J2FGjUtlnVg8okhYRxVtb5sYMV
BQ4jIGt1kUFGIs+UhZ2Pcde2blGnyNH0uYoi4g4GUqykNsxnUy9sPtqpK6VWu6t2
VEyqcFqggwIHFLd+spao24XggwSUt8iXdDECHTDGW+1DOIRnHPDt++Khso1SAj8n
A23gh7mOUhHxC9PDngqy6fzV6dVHHdIu6+FBx5/Cx83cWhOK92C8MrIoaH63v9iJ
4ac2mx0qkMIk4KvDjgPmQRlTvLLcNmbD0ZDZaCmNK7xfbq8nNgsozviyASz2uQ7O
po8ASuas1o2nOR+3Uk4yzPMKk292yL6bbUUwrW/rolUQfY6d4xu1CieI27OOeB/q
5c401m++j507J4ce3rNYqIKOaGevX2KDERLBQ/7Aisi8di4lYGisu06alA5LW3sD
//2bZh+GLSLjMTmTfALVmsNmXDG0WGqWPIWEp0UuBPyE76rSuhl8JwdtNCPAlwAy
uwi6CsYHh2uCHIvgVs6QSUyMDrrWWX4JneM1I/uIgyczWD4SXEc8LmpzbuCVb6mC
ti6/Pg/AqIcFKRS+ztOEh6Mk1vH2rH1c4L7SREDYOr/AmiNllvCODauaQoFwmAMG
vuTymuDptn9ovqBPAOyQFQpaxNVh51VLD66AOJ1mMiKjsAnJM+kipvlNtJS9oKRG
IOSFs4RTrGAo/s0nsWQCxcQ8mOHHUEw0ehtPbiTlvI0+jBr4SnZ621CpZYo5Eq8P
cIiJSgk+hT77i2LTk/99Rlb6slphY/ayZPiFTybA7kBg8QSUEmCTXG0F3xlqHs1O
zzlpIzWzaMiaqxDFE1phBhv3FN8Unupk5CPLGFQTitG0u0p6k/ibCeYQeSrdgC/Q
u2kOcytoJPGnJH79TQXHkoLZ9l9NGn3qGvwW8kI74jCnQrQxYJ/gmhWkCw4q0wHx
R5E9ZVLB+I4fNKqOCffzZdvSH8TPPp5qK645N+GCrgZrRHVy4X7rnLdqb/fiv8gm
ckeMMifoqr8yUwf9jskKFQo4mzOXprIghYFBAYI69lF7RYrvyd2Xf9veHZZuz76n
Sdis5GEqYNvI99q/UWhSIGcDNhAVEBrgAfTHlUVjWA0Hbfjz76mX+q68gnjPMlGy
EZ1mDDtV3qGbYMI5FJEpZwP7hSzMed7eQXB/IBQf/dSbDR8QoYqpsIF6j3NlKWuU
+Zdwru2s+byyBEhVahNNyDDY/K2r4QT8SejQXnDVFp2jUO3dOhyspAhAKwL5GL7k
m7NeAK9wtYD1Wk2nnuizoNkOUQ1qfuISU/bIjI1V0rPL6rbe7vpGk7Xo5m5HPLyw
7/6CkGgW51Ng9CqX3z64NcLUaM6M4jBhpz1tKQJFj2Csa4y2YHLhPzpJXYUSsLZh
seklp/8W9AVS5sITa2vLAvonXWPbqM3AOdmYiTCOjSZeDSlo8hb3mxN0f4HNHpCd
lyqaTMjzh8nZEwmI7rq1wqwEuMdl8Q9/S60jMa4J8HWlP2aDf9zohsoGZMNAN0Rr
lA454/Nle2Ue0g4CAjVhrCO4cSF17AJAqmKOQEXH3iyYp9K6l/OoCCdvukX7tQyo
spCC9ro2k77G1rlZFQ18XWVmxJvR4gfaatb5cX/IbdI01L2zzjIsnazPGgmfCDMZ
KnyrWgXI/BTs8cifaR3f7ny1n/0OhpgC8VjoTv/DMC2fsqTxauqkv76ftAdRlNC0
U+LnxA+Sv54y1y+WCFzmf3gj5gMOUlyyMQhKs24RqlxQd1+AtR7/MKfALnAtPUG8
al3X/qMJm1EqJrnQIRqQkoKSbrssJ1CTNl2S3PkxOF4QkA+zzpUv1Z7xVYTSiJw5
UtXOwSoH8eG7s9L6FJ166z2pfDtrhnwimf0451PL4h8LHj0dBC7nKMgMe89mG0XJ
xIw7xuMu7fGirAlOFqVaJ2Xsa4r7k05R6qtZmy3k5qMwF81Gh8kUZ+4AFhBqVv+F
hkEUx0pLF4D/OD5atOAF/4RVUj5pb+t2iet4IXQ7oAYfxzzzzQwsKMMCbCanWMQT
M70RfVwq0j5EUGfHXPfTaFXbf+kpwFeSj7OFRfsrn8OILjv/bCAxs0keBZ03ItTU
dulhbpFxk2xgI1heYpJl2ua7bW0q8dEi6ngkOYucGohO4pkHVIBFtq+tR7vht0K/
ADwG7eOvYuO2Pr+O++S2OuXv1mxcaAQzp1IV7KM4Wuym/zRwLNQh0CTrqPB6+C7b
zlajESxVF5rDZB5sNNwgdrlRKB9W9Shl5qTa8WTT7IbJgchdjxVhp3/KlL4GB/Wa
UOB16RyiSmaGPZgkB7rKR8utlznvcD2Zjpxqy5RgvuWWuMMIBy0veNWLjk7b10qe
ShXOvWhLoMymSy5EaMeVK3hztueppv/02CQaIskTJ33kvv50S2cGRrL2M+VgUZ/w
4VLbzLTyHG11hVis7WRZZEOVH3Zg41j1+4L08RS5pFfa1iCv6clBXMRLmWRH7/kW
gep0IqPuyPZUlZAOxAPC7vwaukFUw4ZP/jxUzAj5CSLBfjs/V3Rqpnd9frnsrPzt
xPbGm6idexA/mlnLzuxDX+/RHjBSsTXK/wZ+PmVAa3hYFlCylxUr8e+iynIcI7MG
8v2UwII3N9N/J6H40l+4Jzq1oQfmixA3G2Ihcbum2Rf+PhdHOkV2gI30JwYrAhWi
j4dSuQLuORZk6KJCpbc3Sx9dFzn7pWZefK7e+JjVF4Oq1ACwMjHJOJHtSEBDfKpl
Jg3eG+ZX/IPegRm57yTaGXvnfHWEMGzdUmCTFjQbE5eyz9vLw49PeSe1Ugal5MdO
1uYQAAUVgD9xfxBajEsd1lJ4XhA/dJRJP+F9iv7q/NmyO87hvssUIkfrHbhjxyea
A4wB1FCyYFachGXD9K8n/3uFhA1+6AIOpp39IJaVtSsYstU0XArN/gdl4x45JWY9
BgXqTi0WF63c03TRkeVU3u5MKwAzkfeGGpOxS11zRFAIePas3UGASIdueO6HcRjL
IkNLLtrlmie6QEft3vg7J8DX79WPd+VWsLUiTmnIquJXHPN1fAqYJT6yQeUpOUrp
n71JbaZQ5EhsK2RUstD8Jb0Ui9mE+2yg5EIEKGLu9yL50Mcs8yhjo4gTvgWfvp6U
70SYyWXMwUCC3hjXnUWBTahf1pPl8Ew5KGrh20se0Ui6V9XKOiUzNGuDz5LpQBGa
6pUZ1bzBvCKEQVN7WL8EqfZiZ+oOvD5mJ10eMoMFLRdseLOwBx05tuWwyiOdy648
HWnroXh1idTTN4wW/9+EGPp3NPVkZngLHGVBnKxFYbbja59dTJy6KNfAFqhED8Yc
V9OLXI1Zu7a0IJdBsdQpy3kYrGf7Av2EpTBEutxIb/3wShHwJxK+Th0fuOl/I5fo
qttRLVgbNVK/YBi8clb0K4zN8Mie/i+/oD7GRC8H+Pwd6UZRf7X9SAzAVV8t3K+y
wZhWXbiSyiwk08+fT5DpIk+/Eax7INAAYPeLiW/rmtOsOfEJujf8oy01eENe/G2v
WG3fWP6hKjmYz2lgrxgsmHiMFz2MP8AdkBQ4qB/w3KWndmuMiUFSN1wK8276b7R8
0lPLUd6+aHZtDGMVwt7XXYtvc3rAuT7bVh+LKOzHgg1d6l1sLBADqbhe02GAa4Ud
vNJMx01yfublrPweSdzHf3DjVeo/PIpjFyIL7NxZKno+kjXy+da/yAUOOdDk+OEj
hBQ85/goJXNM3R3EwutkgKi19h583y0XRMIQ1vIXR9Cd6aPgas6INiymng3vJ9jI
340mRx1Cy+uqcCqYMA7dfwDamheOs+TPQkc1P+SPYWN12k+lSQWdN2lUGaVrWkop
6SI0sAmRTYyFJQbKjAEoBiePLzu6/ziNPhaNQD5gZ0Pzh3COCye4VZ9qb5i0ypDT
0Sk3EJkE7ijUJiMwpWgOWKkR8UPYdVh8P+OcHST4R1Hrgf37wklq03KIsCATJPkB
jtltfL5rreUJGcMC+loz89JgFLbg1Szto2jvdY4pfOhnW7QNCgLFkLRRk3MhUzep
KMC7hIpIAUIikgd1toIH20ssToMDrSo29LYcEYe1j49rzsc4naajvdcz3WkKHcQ7
cy67n/QwCloJ0b7N85jw77eW7sAc+tbkpe54doo0yBCOzgUgOyDc2HFiDdb//YbD
bk7YfmaMwgPxtf6glH+153Cu5ik3rDAnB7BPWuDTefNuCjM8vgErOP/eKe0cE9Bu
9HRSe6mIb7uQ3rhfy+txhMXUb1fGotZ1VTao4xDHNJileXo3nvQzcl6jwmNXIbqS
QUdKufuMKM63xJMcQ4nmYoZ/LSzdICzUrJZxhA7dmtHYFmIyaylKjBhJX6Y/ajmi
uEswNfQCuOVq1VJ8KLx58yOJgpLxMPrsa8sN8TvZYS615rQ7l/V9LfJG4KMtJACa
OUva2a4xyhDoq2uf0DI88NPbz1BvpMZE+JsC0kDeVMI5XwFmgm3QZyHcEX8BHcEY
F4zGss6u+/uZ1Ry/g3ZxH9onWR5oIKE1LmUNs3t7X26lYSn6IRLuS2ppsLeKzwSu
L9ShsPu3Kzio9iF8rCj8JKprKe+y7oCcvjsD/FleEeYgZzbiZESd8oakQbvKZi+i
iO4qFSu22FLaaATQSotyxIvpIqXiooxam3LgriBTAfw46stloKW99SWy+S75f4wW
eRQ5suoLPWoUvNrZboF2O40jvqdlSOB5qXkKnOXmAVTXjrhQGWxqWlSNR7HSznCr
lra1GM10lOYjJC5eNxRt3LpgNfkb6AC3aJtmzOHI1Ubx4hNnrd4WxoljkParmDZY
Ak5IT1cmgACrlMamn2QyRaj3+zrtahf5a3oAD6QKl256tP8lwILgmL3OdYyLZ7fG
MQl/nD4r4Z5v4bH0wVPt1X8/2TBDNyAjn1Cjzza3u5F/Ax7kJCP/LtKeM6iJ8PHB
tZQmbz8dwOleRo/K5kPuemroYLu1VzfWs4iv+mAwdVsTJD3PyKNJygsTYmO1TYxQ
l5C7bUQNHkQgFOafD3AmhDuaU08BKmbroP777CVx0hE6PRTztiNg3EgssNLcScM+
dh8OZAXuiWch+R4USC1ZKYj7wEj4Vw6wlWJElRg77unt5dA1P8Pp748qbKUfvq7J
Hx2wSKt5kaOZu2tfZ+bEUgx3zHmg9R6Q9ouEiLL7ywIIp9lYkllEb9j65M0Xk/sZ
HW733p7uS7eB9/Oq001nDntHPBRoZRBHDOKztIfZOtRIaAYnEGr6FzRDtWwXtl/0
O/dJZLcYTXHMzV8TDb8Ap8rgZPNSmR0nIEeTyrQ6A5oAkJLxtiRBruEQdJv5QQ5p
trhKWxD56DGFxWrFkUYa1wNjTS5SUxjx+j4/th9lP4L2ubDdCX7C7U4NBzpOGwGi
jOfqRsIppA9uokIbg9aXMJl0IGSLpX0oauXn4j/GPAnBIIYyNp07WM6+Y5isNkC2
PpjNq+J1abBUCALmDqmL1/6jo4+4gLHH2t4CIIVBbSYfI3YXlA9lrd5DbkvpWg8R
GTtJI8qYgd61Jkrh89gPRzlEbkN3A9ZsqWlSDn8IiKZxcUhvDtQgIKgz1KBkvShd
4BPU/H+nch+xFgIyH8LH80D4DTXQ+W7sAjkFQndRkAtWSKGboKZ34c4JbjZiEU/T
ETNAJojZm2r/uW7UJL5yfhpHACwwTXLdJE7Rhv1wUetPilGgxbjlaEbnjnMmAYK6
amATZXhHWeRXsNNuID5WQUnXpUWb5RMbPUj/9+dCLPxm09YXhmfs/qthsy8maRxL
UQYpaCzRVkP/R/rPp03iW6hwubpjsJgEAmChS4MvXCP1FHM5ZQpjuj4fm0UFg1r5
4iv6KnSkOL/hvtz4wiACaw3QDN2ch5Jn1+gcKiIveYtcHz+JbmN//sF1N3tEqO8C
Iq3LHjV8N008b52rQqjRAkWk9aOxZOQy4GKiwlX3QyXb4WjAwnjPcXCljBJ6wKNi
TnSUBgtlhHrtb40K/7GUd37+anrP4BBKTD1x4D6fN/jB6gvGVFL99TwBSizTSkF+
Q2np4EgCYn4JOrS+uJHeT1MCqQfA5Tp9AKsLtv3mtX92myhRuQ/Z5cNhACLIBSJX
iFQ3llE20zyK24zkqEeab6PG0+gjZ8E6t+8QAKUwMfh6Jq4P+EbCStQdca9rr7Ee
0skNVn5eJq2iZU1ZC9t7n0/OsK+LYZLjYJ02jNXQwyKXwikKlV9qzFGl3xg4v60p
wSPSVv8JFD+4cAm4iZ8Rv7fQEgixYq9GNvLmbduSAf9QlHgC0LD//pG8zkvPyRHq
5KVT0vS2ojMQVSUNYHWOJFjCw58/XmMPNOk9O+rSor/AYrYz/3bCI92pW0XaNZrb
j/6maXRF479ED0Kjr9zYgzF+m5krrNIkZvX3XKoQz2VYuoWlF/2x7K+3Wnv8b1aV
eODv4YbxkmAewGSJ3QAryHX4VTRVN2sP2m+pGLlu7ExA+kFzHdSS212I+bHgDai2
KJqwKencr20rF3VA5KeSwL5goscJo3uQ/FXXYSmU/fRpWD6mnP1sDH/ZgMndkJQW
w7L6knP+r3azDlggMtr4MSbW6PYS7GS8wdVjYxXTAbxPar3IzPdXDINUTLPVPdl1
8e/swwYCjyRbPTqVYcJNTmmZRCzOp3MMmzYRrOz3hARFFwjjS1xjUQGJYbQ7c/nd
8ZOYZy1/IEGZqOC+MEvVNUQdCO1MRPAzgws+sCCPfWKUV9yykT+lbkTuOyG+o75s
zTStVLQwfoE7M9EiBkB9vpPmv/bv7WcvQcTokNlv8CpFCNF1bHQ0eRYf2Ca1xSi8
P1VHixlGTQjrF1tUGeQNmZ4b4TkPL1MBpvqdrSxkm2YoNLx6j3badxVLamGEi6eg
l0WaDh39iQN6SA+CcjKvPczRKY6I3Rds8SIrODu0LrD+ppDyNVeC+b/N69VKCjZs
tvkO8GfiCXJUiY3wJFMh8rEtP+gCwI/aw5HTDEg379RaD+QAFFWeSI1L7LDvgRur
HiDEiFNuRtV72S+fAT92MW53yeMnywl3PrmEtekLZPs9SvgRdndAjIYXd2OcawPh
OhFUjEGatMmidE5nO0f40enzvCChFGa/FmgOJUhtzRh/VWy6Hnjkp6bU63LDZjl8
CW4WUxpAHDIEH1zMTlhYedN7vi82+UuDcHDC61GzYKosKeyI6XcOY/qWqaDT7xRB
O1YC5bJ00+v+JKxBNCOis6oeje6fbp3UOhdkeIAwisd9JG/rc3IKQHWC4bh7xboU
3OkQKQbFichlBC9QAyyDZpnD2n7n1xHRqJ3gfivNRkrIRE8vbdVaBoL/a0EURowd
ObTOFIPRfEz8x4q6QhiXSsenm+5bfSBthVG6cKWiWNHLriTReDPNGGos0A972B2z
XXPG9XQ1EY7vm5k41V6AjX+LE1gzaahnvdntf74AUEzdorV5+SEizoI0ieLVtF4x
QUrWscH9TKZvAA4f9zZaWHEvadAlp8LYJfV1aApetcAGYfxJlMHtGNvARND29zvh
y3KVZa3VZ53ry8tigVcvfPsYZhOGz1AYQFsrD3VRKREp+1n+I3i7pGaz9LR8yRoO
iWOejIYkQhRWxsrFm5Es3BWnycSYfrXBmvKJZl1X44C4/Squ9zR5SxIwhx0RV+MY
voFjCDvJ42dPQdR90GMklhRKMjRvbkutznA5Zp1c3KZSwMSeTO7R5ify2KnqWqsX
F4dKGPwYyw/0e3qrkeVaRCjySoP+OdjVcq3BsNnqrq41yB7KCkUXe81dKNBZfJhj
VSsxPRfkTF0izH2GQ/9Cv8JjOKXrffvb20IG5OLrZ2omXCN9YAYgHGUdlXUt1+qX
1/CjQC2rlgxlCOJcW0c1H9hfx9CfXO7YxLrZ0RJEN5J51+943zVVDDn9lhLcNU2p
czF5K7WqDzztiElozpfRbrDQ4Wl/4XTUSEiGqy5O8tCUxfv3wm5/h2M/2hP36ZeI
OOm+pzzn6GtEgAEB6pb0P42LL15qHNGQc3MuUhzmNtk6QilxOktLOEIUbuhziFgC
bn35cA4WIKQ0vR/SrAXX58aewbzgnNx6kPGBFqxBiJbKaoWZr62Ui3RuFw0TvlEz
MBVDyiVemlJEriq+WQEaVgtE+OqivYz57eJtiBHUT0UCCOQQYVf7j1r6PxglYye5
1UXdIEUVYVOIeKab1W9mJsf6l+M5bTdCdxFiz1GMv17GAIwGfoEsb6Ux15Ts98Fv
YeukJL6eEeN4/Ghf/PZVZVKNgw4DshbnE9aeTM1l2TtAVdFWTh7EXiiP+bJOnYbe
9PoVRXm+IuPUN8+yKGFEUfdncR/kZM51CjTElvAisGfvIGdNZL4QijrWBtzycb2X
qZFkUEMSiM1Q2h+iexPrus8PpOkZxPDbHPrkECsoaRfR8vyrh1uJSOoiWERgWtqr
9+fg11k0kiLVsw05kLnQuD04Xi+qXm588G2tP7UdZlsaAgE8DRs8Dak6waraETMB
V4qC9ObHp0/ZC97G33cU1u83lqtS3qLI8FBh9LY8kLU/pWYzRaBskRNej3nggvPT
rwjD7NdJSHN1mC+8EIrMTfEIwgTCuuZTyT5y8Mg0kPwDQJ3SYepV/9DJqO2ZMFo0
avdUAa0QsC97CsCVex8u65QrnQlMhkH1f+Ef+o/60z2Vh/uHLPaJHMyOaVeZxKq2
KQ8uySuUsoNGMw3Qt/2mPfy7BacsOCGPkpDyajiLxqED9t9VW15cEM7fD1sOFNuD
chRUn0zuPZtRonWzAI82x7gvFCg1SBsLVGKTbFMEZRQLu8kcneMKY4YZrlSV0uOz
7i/EPwM1pmGSvxsSWHoIp7+PFWTBg0ot2Hr7qbrchKgNjVXxPxDN7HGpOnZRaozr
gC3BWG6D7jkssnKTFK5JwQ5LNkPCftZKYjEdcATrxp+HYfXNSZVaAeCdCNBFNz9r
pWEb22yH+QKEBKrLByLjXVQPjyzntbUCcCLnzGl0zifQWSDP04W3AXbdCTeCahG5
tEc7hoBV6QABeNAW4fyVjFnhzfgrO+BEePXKOEHC3rU4xZY6bQ7OklxEbk5sg1ml
gfXOI2l3XTRNE4CmgEUhwlJ7IMmLDKewVBeMeV2ETOoIfH/fgYaOc6Ru6aopg3LZ
55Eq1oMPffv9r/woHxhJQJJquC8xYpdJjTQRBxUVoQ1jo1lOUtxl76Z3wE1aiYqV
v0gvSO1VSDzlWfj0DuU4GYmBNl7GxhYIKsYboYuM7QnIBiMwQq0vbZ4xSvU/BcxL
48aPJ4nn0xUZadnEZblfhIsuqVJj4Mov5lz0my3x8mrGQ2Na7kDXkE1ix0juXDMP
xksC0+K4DeA0Jq4NM+DkCOBrFE3VVwx677tp/GucvI/3KUlFBQD+IjXi+4rpORi5
N63eKDVAnSbiFs1Jb/vTHtWmXeoMLSKF5D+jeMxP0JnBgs0PGTEAG/936F92MeEE
jpioTxcG3d30Vt/K0SqANldn6K90EHMgoyzWx6+sgOCyP4Twik1W5Jm7gAeaCm6X
jJk3oTO2CLF2DIFfEcDGNMoz2g+ofH5K4RAU1pIxILfj11GGQ2J6O3flLa9v6IX7
hhAyA+0Lhrpa29vr2z8NaiZf/NkhXxZc9nvY9WNguCF9Sy5ZiiFPlsKL88OgqZPS
6xmVyM2z/B7ihHQWvVlyWu1OMNS7p3xIcr72aD/tvX+w8dXl8La91yn/iOsAhVSs
oM8WKQBLXJewbnXxbPLEMw8IFwE1xLX+My7ZrIxwWBiMTv9YbVQAcEzBE95II/sJ
cRUN7f/HeBVovRK2oo085er0E7sYKj11ujCnSP2ZRtOkbpNawlbq5Dd6TXr//nBS
NIIknDkNUMv3FUHOmVhtum2qhDCZee+oCKe5PcdX4ONooz4ifQ+Ppkwv++2xElQJ
+cqH1kOSvps6/fL+/z2OJ7kJYUJX3NsJ3+e83aCKinHoVTzdo7NAi3pBmZyzGFNh
+NISpwJTBf85IPQsrG+RhZqKWXFwCV0qF4vR57PKQhMSvJFDEqw10sPwuYKeO47k
l0kToLztlNL+Ql6kZGZl8v/d//qzIUBzM0WT7e3EBXVq4hBpIfjcXY79kG1kgdYk
kN1hiLlewhOYFTvIrm520cy6EWovurRvH+AtWcQS7CYjH5BwULXrsNhsJeK1OC5X
rcAyIXuT7RbRjBLjVnvUeNwjo4IICmR1mAN5i2n1/2nfckVKU3fuIAm092ClI4NM
VKQpFyRNNI4dDuzBKqLa0nkGbIUB4j56WOOzuh1u5xjbavbCNIUlPPyxpWneywda
RNa6YlgZCCAcjJKav0S4pExV6hByKbhmfrML95b9TE56+FS444QToNc/K3Vh2rGu
1NWqNoBq4YaeKFLeF5GKNLyMvpsM6uLwtPHML+Mi7O/DSLrTxbGv52OQ1uBoz27c
exwFkR8zezwhTW7Mjxqb5C7u/8BoOQWWnZR+msSAXwjgKFyqTZ8Gvs0nLCeyLDKY
22bOtlBN+d3wogRYQ0t/iRCaZJHXnnHcV2NZ1Prwt6wpFczI0Oals3eGYHN2DNFC
0S5ms53C54adlVnHheggeuSe6q339sBVA0LhgX5d+1uvuqyvnoKAzQzKZqGR1VdA
jpHeTvgs1Zc7b/izYgRcLjrHHlXWj8/V7gkJzszxekFpEDaXCGpc0TbIpvCM9mjU
z7BHwjTxpiJTB8pevY0jRqdlsKy7t/IbV2oPFjJg+Yv6rb3xb8lmv5eMN9MjsHoh
J94M0kYX+FNrxlDdWBPO6ZBcmBKXM2zWNfa1qha4wQxIKoo5hGAWoXLEL3UrTb11
OCgeTyjpAWHlREELIjPHpSq5Hr+4eTcmkjrWGR0ZEZBYzBHDmk5xfNPMma8gbtRi
Li8kacNMMudHSYemav6sj2KCSKvXafWTHyIMqCKcbW1mXs+F2DjFZHh32YhAowra
gCHjEAwwQ8QGile0L8oXhCyDSMf2vhj8btR7RGU2sAdzvcyh1dF7YUMOIf6oibof
ksV53EM7cPeVi8nunM4zKqsIWomZnd1mJo36d1v5hRqSx7cIeW1Z2wgXDhjwke6i
WRmEtxnwGgK9WjRInWdP4T08qvZCHnFcwLJg5EgUk5G8LVE+TJVPRJ+KnrwhRqC0
+t7P1rE2fFZgrdyGp+M0dNyv2SK1CkqHVfeuLS8kEYPXERU8zBbFR1RHu98Alp8H
VuFXjJQ9GRTPqwleAwaSgVS6zJoF799OW8znPF2DO9bZK+RBurtl92jWsztG6Hg0
aZQszr/HWquFOWM9heB7deIsoFluzpJR1G3KgyqXE61rAiwuw4yx+XyqL+fMTEUS
1uI3va1nfyZmMnnsGbyMwzvGv0XqTNNAkziKLYYIy+dV3mG6HBOGaXDWBJW8Z0jY
RQ8yMgbWgj3RBitc8zA4Gcm9eov/fr0E0U3zAcH/6VliUE6jzvbYG4JjzHGKQb2J
blegILZsYJM52aK5qNIfUtpd5Bfa8ANZGGl3L4fj9rTtPYrUtTwZaPAHC5R2nY5D
dPsOJgqOaysPMl6q5wUItdi6weWqjghnFXQk4BUBplpqIS918UHzb7xE7hipQGtF
hsI7Zph37B5t/y3MWrtokSqQW4NamaXQWF+jvPW736KMcKArB7ZERDL/s3eK1T5b
RcJq6zJzoLCWnVvK6OkYGqKnPB9u/f3ZBILR1Z2g3/ZVE4fVzgadRoWFpN3M2ywE
I+pi6/edReHY1VAT6nDX4fupuVCZBDiylMtfxwSiELO+i9cdQyFJGk2YQAHcIIQZ
Gtp7Pqh2Te3tYjvn717UGgxpmHucnqY74KAotumOmuERRXJrt6+Brt8kmJzwY0t8
TCrhkd+a0Qn7hI5H/FGDTV7cLYQQ4gQL6rNbK5w1beWwAWOcbD2syVfRANw9IFn9
JbQOBYa2nmk2uZ2iMVMdU7fxgRYwolKOctIlKDFyKYiuqL/jX3wBBzzXk7oZKK7l
d06KGMZ+hhhacA36O91Mw1c8Ja4tj2p/6zn0NsamxIMoH0oH3+EALEWgG43SHPbj
XmZcnTPyIltvO0Cs6yWU5c4RMEUU9Z0pej2Egq90lBhgg8i1o9kV0eNAC/W9xU/V
MTkJ47d7ip053Hlc/uL0K7hBi+h4mDLPKGNdXdqt11xp3evWlHbngvCEhQeYMRml
g9DAltuXvDbe4ev7wclZNMr+F4t1Q1Ca6Fmc8lJ09R7NAyVW4Gv0cCwpfp5WofIp
svsCZo7vAUCRYaACUZAEjmbCnlApv9qQT3N2tDlc7t1WD/ffRXSK6CwIPSGYMbxF
J+mgWkfB0KuoQ6D7Z9/t14N7GZ9CR6d5Pq9kGS1I6Ks3vUHl5IyA1Pi6uLlxAp6Y
z5a4WKU8f5v6HpFf6sBHwVQ9jEOxAd4fYJIA0ddSz9cFeYtetvXBpqxuADhsXiwq
YamiI+zVxQwKAVRxuBDaejHwBzCBy/srEtBhCMFA0MZZ+IPjpY+k8gu9elXY6qKH
xU4UOaAOZ5qaLmlJYHqN4VjDeMSYwMc/H9y4/wGw6ywGJIh4mcHtvMQC2zRA4WPY
h/MzO1KbmKQeG7gg8m33+/YkPJRIt2XWf9sPbA/ASe3eXtVz/JGh4HCyLIJLym8e
oPR15KlT+CWbHM2v+SYW6FqC2UIt4VxHzfPCFCBqwdV2fcuS16bli9X1ai84sr4o
sm9iW8Ls7nS3jT3OaX+BSFQWLXkvZAR0yzBR/Hakbx0IH0XKMlurp4NC8TvKqzl+
m3ui+825rVOUhW127wwW76drXj7HVGb6oeSuVGihdeoT8cIjkjWXjL3wfQ80RkQy
7DynlSr3YXBZYWviCZzTACYwWuFmQTB2jnc7FmSamxWXoxiy+fUpNLugl1d9qRrX
5Qunsa0FBfaM3uKGhFNFvZMTkRVseobtlYY+dZNSuG418nJUszkdvwFEJkR1hnIP
g84r1CHsu73thpBo5h4x2Sg/CtiVnzN8FE7TU7RKFD5HYbqftmONlgx8nV/pdRt3
GQDDAF7iFVWv1AYNKWPupwpwtbRDUG/IgZfmqqOE9xZBsaPmuomtT8C49eSLP05o
oBCJrrWT6a0aO3UyZErbdG+kX//XOQXqmLXDIqxptoGViWVOZX1mmxvKQj370dnh
FXNHSJtYNX9/4rS+Kkp3nifhUxW3U48SvyUlO9uHKh6gg2qAnDissJ4+547Z5QFt
zTEYW9uh49Yh2N4GDfBfk9ORU4pxVAJ32aoFg7pcvju7APvjLN36EMxOMvkuBFdA
bf2PUFlfbp+ywbKWN5vYyHFmcMQ1YPPnOM0zjwVBDqNI8ef8F6/eJK5Rg7Kzbm4y
30TA5kUNWqrSGgsAv6Q1rJah1V4JuBtE2TqpPw3qx2haDR4NrEEyKmZB+hTJuEJc
Px2Yxb8SH3RCtF4euafTX1eRY4jvLo/Tkef1opQeYujgWJ7X+6ywswxr8jm7Dhvq
RJcCVT1sb/OgPfzXslBbp2jekaYZhbwAgKG46BAMTEgj+GgiTEhv1ENhc7wMIB6g
XzBpHRo7+03hdmA8pRqajqdoqzczDSr8ZUfie/KgnUlJAW+FsO7JzqjHWfOYsMY4
CUBG0rtoz4UPGRSUFrMm5BBVbSavQO2QtuTZVWQZ5n+sViknawQAm4+sHaBSXqi1
nDY9vhKrZrHDR7gWvtu+0kk2UUA8t4rBCvNIFsA8XbyOP9LYbGTo9q0EWz6qQT5f
lDpEdlSXQXLFgCAiTDw4/fH8Bl9+E/odJviZM37Tq1hAbQPwJFZhZ4EKUckDD/w+
chlpod9HNSWad9ZJ+V6I63R7Htu22spQGacc12KQ8mWj8BlqFPcSHIeIXN6dz8Ii
cinSGZdhiPUu6SPkcu9dn6g88WN+SCvcFdfHlle3Dh3cl9QYo+7FkSvEIBI0DQX+
xHHAGyTNoOTflP5Q1FNyeB5wV6r+D90h6iLlhwzVUgBJ3L/RDwTZArhtd8E04BcR
5fRO/6e7d8X6VHZw7J/RZ9EJ7nigjwE/VcMqr3qaEpEtqTi0yuE+wNHtwUMBwOPJ
pR4vlRYoK1Qe5dBqa6Zsec729pk2eijJ/7S5ar+9JePU5rhyK4AyXbfrZHGWG7kr
rlNSxctD0zIZ8zpF4UCvbi/bUPgaZT8GxR4uOcw9+7YbNwsxf5p0GPPs22Kso1nC
DKw581dRI+F3uC2px8vGSF4C/p9Z05eOmOZ82cM1Ge3EZEO6U05yKXn5ne5ZoSEU
upn6COcqHJbFTSD058qzvdFNNG/fWJtMW1LUK4hx5wbCw2PXAxfg7xYVe8COkK4g
x3qvN+Z77jQ4wy0CXHbpZKAEwrCflzJcLOFYZ8FWNLEsCwhoDI/ZJmQdxFfzVcVe
6Irqp0DEyv1i15LGvQxOsm0IE4mfv7RkexlALXR/xW/UZxS+dPYJ650WiNqepb4p
pOCJmZbRiVkQVSsRmGimDRc2jcIQ4Dggt0dgOB38yjMpvVyIZd/UpKEELGqTDeRd
g+kP1xnSd3QiyfX4h4Z0ufdU6p4RW9CupuCic71Oyrc0IPnvQ1dMaZohGkzu2tPT
ZsTZ1V12IUKR+YfbbOwO+iBoqyZK94YlYVX8nFDwCTgw0DC4hEeqlZMsz1Jq1XlP
PygwG44VSdvwlYuPmecyaNra+9w+YT1ftC8c4YDD6Kq5MXBynwxeMA+12S8HF6gm
k8nILF1BSYLBe8bj5euQmy2Omvy0A25VFpbfFZYYbJbOQBEPpmfYy2rSeG3Qzhvg
KIZDOGzOI9cbTwFmIcpTCddp7qcGlHpMqesQWcITa7mNS+nYbHNrBlFentUvfLX9
HQeQdz79gPJgR3HPWPbyaCnEt9/x87eDcQf0kClp9erp1xUU93bgzKUMLHQNYU7x
NDz+HV+xbxNYQLXfGi5SayDkrJy7JnQAnbOGa/HpJTrFCLVQ7npLAJKko5bY2jF8
9j3X0zem7lJ89+i54NYkspZPYzFGi9N8qn+fuBqY/hKGMwSgtYygZ9KMTYmtwcAh
ISJ31U+vv9BspRqF0p3XEa6UcAwiOMP+dXnSyd0qj5fgln+vtXRGR90y+O2lmLPr
iYYmKbXi9/iYpEAL5nmeqDCToX9BLQ7Jnbjq24nfB+9W9rx3EYFo0HsW+wyBEa2o
0tk0yDHtPPqtIXFD6AfCHDXP0GAFpUNPyyvJrXD7RrL6EShWKPbRruBD6p5Gdxve
a5e2oHqNL0N+ZzECiR/0xZtQ0jZdNoDhyn+d32bKlP+vgPCIxXqkjHvpZKjWIpLk
WEZStNs56yvdUpiR4jCfu420I9xm7XDrR06/BXaGTsJ47zGMkC9c78+is2XL6lKa
xh+6ePyZaPqqh7R2ETJvlZlKt4a0MI6hJGrnv8RwFGha25KpnYxeGZWWDfqeZcCp
q1qAT+D+uVWKerxlZf2tU3/bgAXs80UCPwqDuYGazAaHPltMxZRD4675oWoiZYpf
kN0dZniyfL7zpDaJbes1TqQeyFEHAmhniyt4gLD7BnY5H9lBrKuAySHY6RgZPv6Z
sTW8lI+qvRTV/jOyBvB/r+m2xGM2m/+49lUt3lMv5oBGpoHhs1be9E5Qzb80NVU5
MQsJSTcc7avIEBgngshlKTYElkBZwEshxgyH55eMN9Uk7oaHiFfNFFJyHm6UaXg6
fz0JdSHmPde05ZyshIPcWid8XEBQ1fOMHJjAweMkD/r1wZO64r63k6LFIW8A7Shm
y0oC2wvC566xNiMKp3SXQSLdlanoHFazOXOY/sfwdXl32Z/FqWq2yQCLeNTDs2eu
S1kyqzl7OYQD+NRsJc8VBFsWpAfzsz0XvPKmlmTgwqytalb0w1zlOjjyEbzPQW5H
Wep4o+EOeh83lhgkSFCZULvqzom0MGddtGcPV3X93dLtHgl6GtTP9R3qGxtAfyEV
JXGRw/qodK6gLpHgZB7XE2AmNzwa6qPOGKJyaHfrEw+UYnrYFL0L4osh/3OUhjJb
wjKaImrurAfhQg2UTioWhG84MkGYMvavnbLFTAzcaw+1HoHOOqGwWiKxnhidZ95r
yt+PBtGAaZyOgMok83lzsUnTVrC0ZLQASSg/lh7pOFDLHgCrjA8RnkiXxnoPlnIE
saCKuGaTzyk8KojCLc40fu6UCD+C12vDw+tZFPpx2Z2DNaK1DChDk01DNHQWLM2R
bBL5n/ks6wTP4o/nSynSjg9zZG/mABbDY4MNY9ZvvpEfO05x33yWNoGNhP2nxwxd
pmz64gGDfE2PLOAJZjBVdYcxVmbq2O/xonOaW6/V0SgHHDueUpiVAduDbO8qNY+D
ba/OuQzKBurCjYYbQtKr2wSPcTAATeaAKjncZFAzsdo1gSdcpZsWCUJ/2QhnWf3p
XL92ymeshlotPCrhitQKYAATCBh2WSbbxyaJaPuyo6ySvAhIYQ1LY8JLKiZhaOLt
0KGMZnMOewxIp+WYki0Niswe5CROAlvUY4W/fPkgPSvDjh1XS6Xa9eyucTXgBaE1
2saaVKzHhWjHWu/9Dj2FOgFBdZcC7YPm3hVK9aXTTzjh34POmwoxNT1ZndOB/DJc
XkDyOxgRC8dUrAuFJPzFrbXNv5wwoymzWUHzD3azF4yrEzvXSfKQ/YIeEKfSO5GJ
0caV1i53TyT74Ftj5Ud02nLq177BLJTsUKepDXiXiFEX4jxg3P+96UyKlOR1Kanv
EkzwtCPNgBCsZX+UTEYmhuync6Kmsd+r9HTz6CqCN/S4Vrrzw31iWi5G68yparWa
KD6cjJvKB5OGondY2XcLo7tKhJKcwu42kjqtSjwgieYBq9aJpNSaFbOZjLoOlSD4
FeD7Lokhz7Jk490n2KYwH2Fedv075rkcTNDmqXqrWt8LFxH251A0iJSj3GY5kJaV
MNiJ6lEOd6th2fhwuW+uEe5cTknW6AVY6HBPoWWpNIyy90s0cQijllBnNar2RARU
P7QdEMckxU6ehKFLK79WptcrXfFJ8xjl8tMmBieS9gLqddppIQwxRKCQnAphZ5gH
T8QobMpY/T7s+18vE9Y9BXzHICQv8ntwQ00lRr+ZlJxITgWdJz3k33e0u7nyQRqu
tzB8cPsN/2MV31ICzyFsmcjlOS95x8EV4/HR6E1HAZJbZqWrhI9hHgySDRjOWKma
ktToQ8aiXU0bjO0YML/dQpd3btmZgjdLRNa4VeZomT6q33WSR6T0wtXquSty3/XT
NLX42vY1sXPAaypMaxXmq5xqbhkPMdosV8sqgznpy8N871N5zHY9uhhLDzDVnSOG
OR4wzVCMD4+xrq2o2ZG923WQxs8BqZGow4X90Rg01gv17UZev0eddUXSuGiPPt7l
vZWZidMXL3bmU4oyx31Xv6R8GGdWrKeOERIMNl9kWDifq2CVXT6UUV5Lr5I89Mbn
R2Lka2VnGpWT17rlAT8zBtdwBf+T6jX+qhsHRTM+roIoC9fACt3kiaWmcWCjXbaH
4jTj2A/DBZWwUnt8PyJZJjzasXrBj4urZt0hyds+STm2xR+Is3FOPZKB8eUzxrSU
NLNB3lsDs9Ei1iwIeCbBJ4cwZ1JviqpbErK0hTSjkt236ZX+gTCsvPvKNgkGLxOH
r0m0JehaPYzvO5kZf7VgoEa6fOlFDE0OAUIhZ9gAHPXk5SQrrLHOrZ6xW/bg9Fh3
KmrJMl1r2ZG1wJ9yM8taSvwZEl3t9Y7sh8KmXWKshZqw+aF7xmJgo4TzcxWnymUn
RomSBU/C4LG6LYNwIymgvySZsaqc49doIswNDh2lMgiyZVsRFH7E3WYtGh0DlE98
4A68mT6OyEkjFWnQIZnTyW8Vlxm0OgvG88PCCUbWfqab+SIYd1oJLz6Nii8j8UZb
kMxYZfv8aY21iyvUzoM/qv8ObYueEmTwoDDjiJQf8+FAvQfrgmSrg/glX1IjWlvM
7jLRFUexQ9WuJ/0I7kVunLtr1MSueqsy9qzfXYHxcQxvQB95Cr4t9+8f+TnUCr3G
henYq7w1uqgqS/pl8jNFCqO/4gVw8acCvQy/SUTREzFAaIvUkTlIOm0TOxodU88X
4ZQ3Zz3+JMgN3r8nNwQXR91Vxqp9+4/meTUdx57Z2JuCUX5OE3hbevOU5Rp16D2A
BL1nKAtmsmcuFc0lDl4OPCrnSCG+po9MGFu+M4dRoywOH2WsyxpywNRE5XW2+w6J
FVBVDGOfIANAojw/SiVWqR5Y+IId+K5pWma27Phcnjeqf3HzdDZq8AIB+wwVj5vG
yug/A6Nu54LgRm/qcRTiAGESZb1IFhSaf/7g6CAvS+at1iwE+QF4BWIc0oEazuLw
3SODkN56edU1VEnWIkhfGOlHGAskaL7MCA6KYcbhjN3ge/XaLAUnYQAhCNxuNHz0
5XoyZrm2Hr4CDdwARZf8XjCxsEfX+v90PfWjHRV9wDc1/PQx6lmV7SDxIgUvkx3K
MoUFtBPfBdv+i/BPkxGE/JH2ISYSyylM6uqa2nWDDOenri1b+qz/wWta1J6RGIC5
8B/99tLksr54Zkh22mFnicU8K2l6NIeOLM9q7hjb95c7WUTVjDrslBQJKahZysgy
TcKKZT39cL2lHBcaQzXFm3yhddR2RlWENKZXwk4jbF/QD0jr7g+QfiYrTn+Tyvaw
BGlug/OJ+tZJ9zRyig6LCIHHpCAP8Q2NfX6QXaaQZ2/peT6xJ550BgKtkIJNDYt+
eSMN/C2Nf4mIuAPSwzYrhmNE4j2fX/rsIBgJhUTaBc95e6zJN+d6D8AKpTmad7bV
Ay7c41m+geDbQOw9cMsLrnOlnR+UdPNlhJiSc8AGpQz7xyqEJniM9pO4xO/lhzM/
fRx/GSLRpZMX1GsRNFGnvzuzU9/aYP9dADMKiGxdx82ml+X5SKGnD5YuUwMHIhsX
vmCmAiZ+XW3Ugp+0l6/viqNEs4uFwCdVxQf6UQYCLhiYzxGTWlzM0Ujj6MWc/bqb
flvqaHWxHcQOA4iEZLEIsTwFAOxciRZ1tV+1AUceHfvVcTBzpvq83Q/peam/nuAd
ENFbKoxnMGsr7KB9TDbq6znWAe7s9VbpWv1eK+E4mV6TjfJU3PPeOVzUnCkIkjMQ
iGrrn4jogeRlKgK2WWZ8mXfO7UeZXACaWunPPxCUKqZNdeErUCBWuHYvhgReGKTU
7xEaKqyraDM5KV0n2TtqByE0e7D/GYIhfS6jLiwu6STjC2fg/7KuZfqnRL1p1DSA
GAqmlFUTBLyxl9fqEQtRMrZA/S7yrfpcC1yCP7y+RLuGPYwEW1os0pYlhX1g1bAf
R9BbLp5VfRpzunjq30wmJBvkwc9lMC1QZpjQCTVxhelCGrtq2O+3is83RvP1QQfn
ZtIJAjUHOji1yezaq04pnVoMUZhKHcq1kjuch/S6KlAXdcu3yAxjYAflfibCHQm0
evgfm2w3ZJFgKLKcIo1YAIe2IyT9M4BWd3xqDnD1gp6FBNBrrdL/IbxNuds9u2us
Wc07KrV5G/XpXzLbHKMjIPl9AJtNWLUfVdGNaTjv3m0X84lHSYatZC5jECS0s5Kp
SYL6obR4g/GqdZa+C5NocbyzQfr6e7IsvP+BUwIPIwoQXCOGAaunZCD1QfV8bX4I
uiQYLhzGFKeqm2o4JsrrR9zl9FBfvkFW92oQy1ewDAhyt1wVppo52GcMw2oKXAuu
IKn2qNExXoEqbRe2H7yvqaGO64xmDiuzN/uwr/mZ+zihO/YjvCVAIBycWEmN2eQn
f2Jg51tWfqmLO2axWrowAc7EmEz6Hg8FF9w4VmGGeroZDtjBrmZQzkTriHNNbCZn
mYR1SR4LCLB4ZvImwFD0IAix6DwkVXVnN9KFoSW41tA3vBSN0JfxuqGVw0cx1sQN
5Xvf1jxpSVGBTx4m6MWRHXxk0L6ugrjIFc31fJGNgl8mShhn1GsKExxVTrIPhKTk
asDpvZPlbDKuW64UBWdMTzVSuEcIRaGco/7OaLVEpQNZG/ef85G/qyRy3Oj7Ogwr
CpTZ4m3wXwb2EBcnchgLmX8bJnGMgzTTpxENykb2OICc5NfjCBy05KWH32dDeCdm
nDDdIquSfgvQkaAYKqs/65PyQNLZMFMzTqw/FZ/CEcu2pWxEkkBXhk56k0ZPVs7j
AofF1Nf5LxjOwIfFPpQLPz+ad680d67aTOnSpJUGSK/SZJzqpSvPtACCqoG9gWSS
K4Am9re79WOEDRYcqUPsHYXmfGT/WHEjTckI67DTBf5nYl8Z4/VLFtmbvLap1zpC
Djw52/oxm6E2fjNAxGfMcg+8iXIbwvqg2xaytcna6NYegPxft/fRhQh+d04d+xWo
0p5Y08gAjVlUtJK/n6sW9lKOz4jikmNL2XLHbl129OJ+mzpueDBIQg3cxblMAgR/
YYdFdvdaFfRc9Jh6zI+KZPezQ0jDeF4ztvsGJFjSmRWnuKjhQmLcBz/1vi7MCUqP
ucd3rcWdxu7YG8HQytPYvmWjLZ3Jz1SOnO8UTs5xGppcod7Z2estSJfm1zTVJbmh
zLLwMYnRnsiuDjSShrd/hqpsdYsaBVqwAQJVpI9ybmbYmIvtVThcw+Wb4tLpf49W
QKmnLWmXTvujQJ/Jhvr8on37WTP6W+kMetyRDFlNwj2wI9A6WMpvYqV9Yxjn5RkC
JQlsj3+Dp0j42gr5D+rWcWZDhnA9CPFLoj8N8RqnEJc3lYwoXGkKwEhFM9trSAEu
/BCu83yzoJaCsuEmljW9BWsTbJoIsyugvAl0dK4VfgI98GGbendr4nUK+HQ384mP
rgitimUsVbhFO7csmA1w7fQ4kOwgNT2DW5K9OKVqn4z1tIKeAOEv9QVbd77pHHlS
0CFBc0jZI7R/l6qTYNXThpebmgxC3OrZrEomJe5bBDvOzBRd4yA9ik6OcjcVC7Q/
/99zfJkyVysGUFETjR5o6zsaqVgGKy5DylC4mYj8A5t42X2LF8lnkgOcMmQAKR3I
b6PQy56Urp4uRlEdurfNJU2V3k/FSsXDma8AWIuX9pp8Ckh013QTYiI+sAMc306S
DE35XTLceOp7xydX//OXQ1CFWoBbGVWeF5c4N9e5XHE0kS6Kior/uk6Gw4cn1z40
nUwLH8b0zRBCO+1QxyW2Q78m2+z+oLYuJmsJLK6q22hhcDnDFmTmvkvbf3eYm5iU
mFX7JuWiS0uHmv5f4h1iXEdbk8jEmNVJ2d7ERJfmGQrb3uCtZk70Fd2/5eegF1Ba
HD5Yij9bLkWA5qdjVpwUyQPDllMBKuGb2rjQhM7SdScHnoaTTGGAAwguDOy0SZLv
qCwTz2VmZicWeNGzyZ2gqoBo/uudbAtv7khHqKMzA5prpi9aZ0MX6xAm+sF9raSd
nR0pwhEFjnLRb9hEYT0rI0CJp1flhrFCGnbAkw7RmMZAXg5nkZPCkuGoKmUt3tIG
qKPbBmFGMhDsdqmCsIHLnBCoyoFvg6389yLojwoBxy9sac78MdY1FSXq1woUijIS
b8rhMZAeFSGWr41MWAGMdhIK353CsRgT3fahvdNAg5PmJQHnmeMvktcV2edWAVNz
0aaLjOZwyiXeqWUBmfRzrfQx+epNtTAr/SorM82iehLJpXIy1FxxBgj37KD+TAYD
m5QrM/OC+KQAaF0YKoBtT21D0XDL9XY/VH1uFrIwudJ8vJdSCynDBD/WrUwozWjD
nSELWMPPK96XOXmiEynB9pXtpQ4kk1z2E2mhcuDx1yD0LoCS9auYqHv35FhbXz+5
A56UPVAK7eR51x59cIC8HSY9CneAPOVL8qHKq8AfMoF2eTDOdg8zrDpV1isU2jEn
x4/MYkW6pbAAKjinmFpBL+6p+pq3u57oSLEf+Zb4SuqVYSbXrm+aT6uEsU7fjpSm
dKYJkdMzSf2WYana1iwAch3zjb+W913ii2hlkow0/MqMQpFPmf8iMy0VWbmdHms5
HHHaLrM6kyQJtVR/tnYLI/zO30Sm/ZiFnmbMEAbJ2MJrXzI7wwtA7mXXqN13Qe1X
AnXzpDJ5virCzM8b+gzqV+J2hvxdeSNIJ1lXOha7wm/EGmf9Bn2OymnL6EP6QLNT
YBDthXEvxOPFQ/npwDv4VmBtBlCPTShXBk2x9qS+Uu2aTH3VoqPNg3D7pekfcIhW
3PYobMZ1jZawrmyjJL8LOjN/fwW0PtprGbX6eD+cRCxNj+FD5UvRwtrXR2cpEQ6L
Yy5vDGXG4cQ3hoHPFE0G2axh1U8V+Hlu4hFOGd3b7mAJG1m++miy2GBcVf3ttxmE
G0Q6pzHg76WAQOuuDNC/CMS6rmZjW92uXl8HzavAmULYqMEuykxnLgG8Hzludaub
q16F9T1nwfcojnEf2f+MOi84U7FfX/bUYGGSibgSQU4SVaBkvzaEIoFe4o+BoJXl
kPuMy8kZ6quG5ontaDcS3wEhidIlwF46aFgRwiH8ESBFLRvBgkdc4covSUSlD7Pe
0zCqaDuVMr4Wg3ksCB7gzGHMa5N9s0WO35MXjlo5GtV6qTCRz1x2cFXvhlRs5p6z
yPQwZLw4QHQM8xvFEOqJB3bea7crnu/U5f5Rhq9a3tNib39orMCUtepZ97M2wA/h
VYeLxUxpojLk4qwU3FKLqdCB+dRtFPXtuITOygI4u9LAa7pl1/YqKkuqPROMho13
3HVQQKSETzUEJlDn8aJ5NpYqgJzPTefGG/OHLxCZ946ZlvvMG1Bk49cYjpTFtp38
asGEkB+mIteimLTLyBl/sMZCjMNjjLHiOa5SUrfe/ZBI8fg+koJTNZjWFYK6Aj4V
C4XwH8sh4UzJdCtR31JUE6HUkFXQtt4HXMNoLFYbNS8Ru+QRuV5eVsqPhL2aXJYm
BS14npiIYDDkYmnhY8tPohsEhT0oVCOTK2hqQBoMnPiRbwx1Ov+SXwIj89fauWtd
x92Kpjm0jGkGo7/QDNLVRq1DbCs+eg6+snDWb1B4cqps2wZfyBAGdH/MHa9ibPw4
CiNbdmeBqcUnFTHnm5KLhx9BcyxRNHFsl4CDCoDvg+us83whhM4QgSvexCA1B0sT
AznOp5IiIRHiaiHqmTmBQuyyyN1vS3OrrEPT/PkFcTg7efN9K0Aux2Kn9jfuyubD
sBW7gol7xFtRJd8Hj9oGhgOkm5Z324ES1J+qYFJknlKZKc9rzyy99LROTgyRshD1
PFzb8oyaD9+dIXeMw3I6DXRqbYnQIls4bPJo7fq1adh+kVzMm2coBtFaI/Vyv+iF
b3NijmPO+PTym/gcbVOmkD8XkqWc1PqJ0HquoQEGk3NS8/KJWvP8bgvzk345scAJ
vs8SgXI1ZQokIezHQG1lYBT3z6pWvdbe3+8tFon0phW1b9xvUODAe9QJ9hq1LRmI
mNCAAnkGVHzPC50ae1wgCdTMIwWMEKvNWIhHx7cYcem7BYYqd21M4teROMn+r0kz
YsZaZA8JyLEnEWBhkK8WsMJC7Eco5FBoNRLWRRoesbebELTkMtHaFmx7qc6Y7ebZ
gYFhpFXh5YLx0Zobm/kjgGaOlfAwbHMd17pP1zdUispcm7MKaOusGW9TQo9BQQUI
l6c2lH7iYuMJ1z5mfEYGvNEle8XiOQFkFS8ueZ1nQQtSu6wRFPP+oGkVnPrfiMIC
3Thk1rL5OAQ4S1JTfVtw16IbQpaNxTvnA0mMumFKjK8DTI/IQuUepBMNJVXng/Pn
5yNWizheYRP1kGfpd4CiX7c1/zDNPshztKKNEikIKTawnux64pwGcnPLqOkvDQ7j
mgHTlQdumuClASNmH29vnDXaKbIuRS4PGhWU5q9ZjaHaOj8mNaXLLiNmaNlTnNdQ
QX7wvtXhDQ/olFLqB1OuGv7ut3DH0L+zF1pvB0okrsjIdfvzUbkctKjgLYts1Nah
jHt4kA+vtmpYtd5oSmmVwZ5dds4meteuX8h7rXNvdXLMyX5/7JqS6HAOHBcJzaBp
fXfa7GlUkDoyRfjJGQFTvE/LEVpOnht29NnTRTQt5KjVJZcuVkCocMsTyFo8zuka
wFNNF3ZYW1bzJYloysirIsIiLhtFCoHSBsn+konAvC+oILa0/7PSlkmDOJbrQ7YX
1qZRGeWA4WAEPB+x1iIOHjZey6VEy/jfwcm5WtFHl9EIUcCZ5PRz9Em+1B3l7tJN
q4+O+bKKViquvlnW2YPs9ZCVaf4WWHPGn7tnXktyEoYDdqXZRoCBaFdxBD53aPhK
LAB7E6AiVZrRaMDkDFpO69EHPp2maXkSMupLFjWZcNG7fzkH+/pPm4sLRz4u+Sq+
80yOTBb+HpAY8Jh1xNC0u2ffMhSyyQRxp1yR5g6UX+vm7D5xxXndssJ7BkxPIH/2
nOaTl/ZhQc9IzEinJUt1o3g6NnfwdXdujKUKs1vvAKDBX90FlK3II8Tl7swyKx5M
JY7NM3iptk4OUT2P9k6Q0ZQvES31tNZE3DY28FV6AKzvaNeZ6pI9MFQqg2wDS8sv
xLCFK5RleMvTl897wHPePpm2bu3SD7vJet6m5voOjXk3BV/bYQOkVdULlL5Hf3MX
h8QYRwWRY+BRtv/By9Fz/wczcJ9OhzD1d1sEDKQknS4R7gdLOBRUHhVH7/jluzCU
KlGNlxfXMbJKmgcC0ZBOU3DqFykMyxpXvYX2PxORVQ0/mtib+Nv/avHiRcWwTYA3
FSSzj/nDT5j+0CDpIYCEu5pMbmAT/O5wZ9lgZeNFurVIbCqw3dOXhSMs+kx5EaWF
CXS5JehO+XLCRWM6PZllC2PnW5eC6TDTQVACKlwxTRO19+d99KLeDAg+dHx4LJ+J
Uw0iF/3oJmNhYi7wR67q5+0BUmmbFAcQlACjyEMtQuR5/PpPrlfObdeQ4nu9vGx9
wgDOQZNT2HW85W+5E8rFWtlTbmnFsg+W8eGn8f416+R2t0NqNdpqHqltHQYMsPTf
kHqkKcX4VuqaXzF0TPSsTOhdfcFHCH24jZeDY08PSJzAvt1Odd2H/0Ozmz90llGw
ckl2iVkwQ7dg7DWfGAE3EmxDCnppa8TLx3XFKY4UTKolYQOh25dYbaH0qIyQ0yjL
OIFfhhJ6mIYG81y6G/BUWGTnTuF+hDGLs0MrQdIDPil4PprFazTUPldiGjOHGEX6
GvoV42T6GzEpApilgujPrLNrwbMChOLUY4IKzaPC0ugrQ0PkJHgYUOSrAabInURJ
KsTmJoGGts7Y5kwF3o0q+mS2frGm8OHe9aHtzY30JlBitiXcClBH3Iw/bvXRGghD
NTQI19hJocBN0vy4I1HmnjX03/4JR2ra6+EGU4sFykGevrVvb34JMcfPtMqu2YhO
y/VH6Csa9RrRhJKSiDO8KXyA/MKyuRYyQHI6DJ+TokPVitNnlYkXPFg5sudztEpj
+YP+axvTnnWXDt2TXTaWx/bb711K+9MS3LDQYL6E7ihS4WZ/5X+asbEeiJJs0zWN
c4L0GyWohC/3M28ghHgn40ZrFmumrBUQrlQfE3KqYPBjNfOgICyERXB7bMVta2tH
G0xg0RGHUybMJlVQ1ahyVxd2gFMaO+5bIKub7JpYMXdKF/HOXJ0g2wNOVQFGZWcL
nmAA54EfuDgJYyB0TJNqNW9MDM2kyYhZhBruF7tFD/yrFavF1lDnyytAsBbS4JCJ
B1QxABRNxsPkAb7HkiBOzUG9D2bm6AgSOmt+1RS/8no2EAqFJjEHj5xHQBYjhJym
8knWvPRepJUFAPaE2iKSa/RNqaOw9O/SB0DlK6JI23qJSj6fO44LdCP2AgBMr1xO
LcCXk8Qbqdk/411WXV5VaEhs/6/buid4koHimuGBATkOlx+G56jlleWPzVV/waUM
yoHDmcB731YDs+JQMGUgDMaQ0fU+MTYxexhbe+v6V8r4RrP1gzUpFTfwoeH7BePr
Ib46uR+yaG2WGrrius29eOICN/G2qVJiTfy0a/bZvEF0m3Tji55Up60oVAsvXrhk
oGhooKS8tGNN51XmnP+l0B9CBAt2rkpXlDKa1H9c+YjIFZN/t2RHqA4GDhhZQ8Ia
iguB/thWG3xOFzMLc2a4yurfmQDzMXuwhzyWM2vDuA66wZpKmTovCG1gUWu4WqL9
jotok5sRvtDAH5s7c+xeQthgHbz+R4ETcOwncGu7lhgQxoYlQqqTGtCb8u3g/Se6
hXf38KcWCRdZE8I+aJ6coTXp0vQrfPtHVJixKFm4snXXrzrKadnYhkNxODzuRLnK
z2umBqL8wXe62WmnkjCEzYM668bwVvXtAGAr+t/euYinAPNT0QOQ76RRBE+3CBOc
wiQbKJIASWqN/g8x3eauuDeXjOhV60p5N61UgT1eueEN/5XzT+x+9d0c3vREKch1
+dK1BvIYHai8Ks17uIC8eqXbFmnLp5vWQq5yIcN1dEaiHbE+tDD5vs8xf68HgCY3
J8AhzoZFQ1Yi6vKb6yPbg7fRQb2BRqrA2A4omnwlZufzHzm91ShL9PV1N0fO74cS
ZBIP5dEye+jPTKiALtItvLT900/MXwMd3ENw6uZVAwWfHOBXmwnqpZbCGYLSrzhw
b3EnACpzpy/VIp73YmdllqwduW67PUM5O97DjT6AOa5XCTeoCQmH3612fi+925lL
n6pe9rLUr3Peiw1vuazzV1TSTBT5bAHK+1YCM2pUCbLJRY/GYHX3vT0IURl0wsyu
n1WrhKb0jEjDJuwimqY6cYL4qObvIoq3NPVmJAobmeZMPDHzACocy0GrEXx1gIdX
3a0U2nd8MKoiF0AcEnrO7uVQvUTle/6WL/02eOPfaPZmsvHD+xgUNzduTLwxxYQX
7ar3tub8oipRYRYwgR+7JwdtSa9vvFE2HDLW7WE89PjXS9cMIBixfqzOGr3QVf12
HBlV9rBEJABKBZJXnaeUrIMnzyZ1wJ+chi7JDU+pnZ8wfdC+i6ZFvetyk/xKFg5F
T0v19aDlxzucjj3s3h/iqWbiZlGNkH0No3SanoIpNUq0+fPVbYcYl20QQLdzLN+a
volSqubCc/TvGd+qSqpj1BDwSB9nuIzpqkhSX5y5UpmlQJrz6GMg36wtfhuKeuXe
3QlSeNusga8K23GZdEVeMVQOinvJw6B/4ZNG7Wn1JgfFCL5vMkhHqiovf4Zojfvl
Horxh3njUu+ojvz2TXdDk9fcbrd96dOIk20xt9RWFqYxS/veDAqTbv7hlqsypypP
ZGn2m8DHgiuiucFVnXfiMHl5Mh+gF6FpomtffyDzJHY/HRtkX+0oiGmjXINa97ib
6fpUqTtBLVOZHiApCCz4V2C/ZYbeebcC6WDoW++LFORi27njwQ3cuK3wNt8pvSZ1
tNXyAciEQMq2/W69bMI0uxWUgy5FXI+UaIZWTPTLZwokbyBxZs8JH5HauY1FiXnh
u72QUq6+YjynlknA2WWNK+MSKwqrycgDzANM7eEYVov97XJHMtAsUGZES6cv7Gq8
01CpHKDw5PmCyaJkEzbvxlvSsgEwYDUNWQBFHddaFMSKUrHp2FD+9DHOwT8Y0ZQ5
KYcBJ6tmSnCn1wTbLq1vrVhh3GYeblY+UMWMaQGwYBNmYyVN/h43NoEPYyeoK4L6
YMsa5ktWuvYX47zJdxX3bva0Yy3sxMEFnkTC1E0iUMT+CVlKYbDfzwy4nsoIrNCw
/q3cY/Ex036mr7adU5SL2UXe6XR/RO74Gnornb9dxE3clHA+EsLJqjTDLl8UZMV3
j4T9EGxdxgRkelenXB6Pi1jvOQKY3STiv4RHLmpZ7fXv2mR++st+4nDCB56yL5Rp
vFjwbcsCb1aAqYldZvVUF9ddReEMZE/+tWmDIKyJDrTSP6r2lk7Q/4I/vqse2F/j
twmvcT1elP1Yi6IhYL/Ag7F4gkP57RdFje8O7o3LG4JcZDesVVwloYZcXEACasVZ
u5EXSEFHjm6i8r9+RQEQMn3mOaXlbZhx7tVj+a02ben8lkwu5cGJDGlhS1C42t1m
YXdC9FZrlTc28TNhIQ/JROjDYvkCsq+M+ik4omVLJgMDmP2QIdRa5MlAsXcUEOCd
VODxzR+8LY2tXmnYbAek3WUlINRNf27uL5wPGHwA1WgXMKM2bTCfb2h0BOX0Blyv
Fa6WXM8m+3d6wK2Rz5FqQLLWAe0fpHaphlLdXMqSHDLm2LqqxmNQBIsPvTlYBe1X
JxeKRLjFR1ud7BRGIvnLN8Rg61yTZeitpVVPYDohhOUh5nJuD/+7+oF+sQ2VvcqY
unlBS+tO+bZTrd4PPBRpXy8TThVqsB4wwn3kABwayybvq/JmceLXgx07VX3pYoeM
NBlgOtujLhMs87tyU1fo3oKdUlOZm2svj2qyHaC6K3OixocVht3cRAnWe8KkmOif
frp+5/GG5uCzZLBRl2yCfDto+xbva1l+OpNkEoB3L2bA6ujSXXPikQaCsPE4QbFp
+VtSHOaJ1VggaVknn2K/AiVJdZvhBgCeI6R6/Q/lpx/I+bsbuXCLnRCPGdAcVvd1
boEgTDWJohGSUpenFxQfabtRqE2uScYZsxQObM3MAjiGgcfKuZI/AlyUA2Xt77P7
6ITlnAGOgCxZbkG7RKBpBU/q5Oh0pcmEMgBuIANdAzs4D0Kbr5JZpohF/IXxlu7/
Llt6VQIA3R0imB8Inocm81BJBwCEHhpga3OcmhyhfnGGf9KfYtLX8E/O3nYrUX97
M9l05rjqzwI7TO7WscF8tI18ScXAXAbkyrEkpnKDPgMBw1E7u1mRjVkIG/IL5SKj
lU5npq4/kkq5n4Ero5G8Uuv6SgUYwYEV1ylTV2Ex5TT4V0m3H4h6zC5BjyHPr2Uy
qB6c/btRFUQN94IgPcgbSD+fvVY0WvQLC2H/uqX7fYHLhkKt+ngkxDY2eDbiaVPo
kn6TXq4ZKJEVyLtE7gfJqeqryIArX60tC05LYgZJLVdaBSBMhlSzeeGM+6l0NNI/
DAqBh81zwqlbR19HCzsizZOsjQdVhEhJ4LFseSHsH5u2vqkBW3+VqUf7PphJ/H5c
FWGh78GBl5rfFJQ/DFL7U/JjeQSvvdaHYgM71I2mzqJ+i+1XFC+BMQ2TlCv4EAv9
esy/96y5q+olFEe1ZQkK+rg1ykC5P9zszLw0wE9aaWst8YT44c1yJNwQc1x8p9Vd
QWnTGrzdOecWL2VxiDPCFEov3gSgjnT2fYlwbl4f//de+sIzLRphhlqzyjDKirV1
NyXUCfAk6AxbI/DfJ/er3a5f0gdxQ411y4URoC9zKP60VD05ooeU1AmIasESOPO4
6kQoV/c94aD6n6rIMWrG25r2K3q065kRkqlDtgv0w/H3Hau1kTn3jwRFUFMkgjv4
01Ydg3xKwSLG4KIK9Sg5+AmdnY/L1mTBqnTkjaKz/P54b3/4gN6U3h1CzsuyAPX3
Ly4g3nN1iLcGebEK4UJM2xU+I7CW0sD2IdrzzowmB3B3a+C8mQWAQBYyJld8xElr
2WI2MYOCiRR0/Gs2DmEejV7IpEiQqz6DbKCBUcHV4g4Y3emlfM9L1ELnHmnYO86K
y8S3Ry9IuMABa5XPwtzZFm7WDGepTD8yUuieHr1edVxUEXLA/TgyBsGESlYGneJ8
NiAzaNjLH1Rz3a8KibSvFU/uoahu7e9fYAruK/+a+J6jANtR/ahrI0PuHqM47mRX
BD/nKRIa6WkxqIOtfphcZ6JNBPg2D/JNU/oVI6HfCI3zilGP5HMuOp7NptSWhZHZ
Is6j1HRSm1RsRfvrIioxFAOoFvYHGqx1ZWKzlrjdbErR2zRquNwebBbiAPEl8I+c
wdrZ3M249rvYG6fjivEkGC7iQtbIe+BFHcmFl6dn6V9c2Eg+hUheEZPeW4KNRFlP
ONH+eSTdpZy/vkSpiCyP2fUHzGkg8Ji0yEfTvEWZBMjZz/OTPOTSNrY7I+m5KAxy
n+E5Hc0YhlQZAOO3s9j8YZywieIzXKnZnuxr/Btvl3mV8aOZ5JwDOKSMBAjgGvLM
skOqfahxdZ8+I+1IiuRMyThiPHqjIktLT0TiB8fNJ5y8VBOyIpv9swDXatQu/wxh
fSAKov/WQdibtqBXI3Rqz0wRP4zxNBkt4zQDRTDcuHJSX+5oUKvE14+JNBEope42
bD3BfRSSbvo5+01vx8nQVxXEvhvuReRdglyvatMbVFA0tk1w84EnWYe12sraTMxC
T2C+lYi/EQn4yhd5jII+e7eMHlhIgfaLLYO9baEbDl8+wAnwAv7xGVtRZ51kqQNN
Ocl0q+7qNNNPQFD4IbsuALAgY2cEffw5j0IcdvAmxaD8N9hmWBI8PDmbmyVid8OR
xU4psfqmmP6LwO6pp806PNlxlHYe+b+cSvGlQieIqJWCBfNIRV9VOQHiSOWfTbci
ZtqkIYWDZUybrpWIKTdSbvS7LeaXp88x+XlVjK4lx7VVbbOxMRIaHrY0uHDT5viV
1fq571E/EAKyYnTf2OFAMoWmHZ9mLzvAUCwYdwX0dj9FvwY9/o3hQ+SlfDHB87e2
3uAJJTAYnixhROFpyJNYq/1FFIrvEePEcRObFZygi1hangitsYQ3ZyeJwUwku1bh
TeDbrhYFRolbmWISZD1hqugF3LrQeO7arFPsyjANYtZ9AiAyNbnc/2aijB/p2yeS
Er14TvpxJBUJQk+sL9s55Zww86dV8k01gN+oufEA7yWyUmmDPC9BBC+TKnyAxWf+
ThxFaMX1BfKT9qUVMn5sT1lRfBnJTmQkAcr2CnK2f5HGt5Lqp1kTzWLPE23kOCp0
zWMqn671bet6p3p9ZoHJDJujY20l5qQSEA6y24touGOditKBbH3lpzo4JgoqONnA
pl6pdUiv/A1WVBv1pT/3SeZdWKiQ7l+D2ELQhJ2HNY7nMObjKPP9Vy3u4WWhRqU2
85vTZa/C9muv7iERiV04YanfA+o4KxhT52Y3+n7nzbuW5ZfdOVXT/KNKJTaIaWX7
eSysjGT6aVEMi+Dex2rOzeUmCVGLyGp0NdQePLYhUfMLZuXHgXLQmBDu6YXmVDG0
C9YwcpQJIXecofd7GrzzggiCLb1fJ4JcPmAUbiwds/V190Yw7b5DBzi5fMlTdURV
earP5u3+ijTotHf1cpqQ1rmVpLFyDAKP/4k2M3GB/LbX+RGAF5xjZtqaUCYEebRE
vhZK797Pq2/rpAVSpUk+KY0XvZ0/qASY7L8ytQkZiaKecvxRIOLYHMQIOAnyUiuD
mjeu5+obcf0JFty2JKNRj8PKIrUARa87FhKlHcHiNNj63IkhmRv8jxZGWGtxkT+N
ZAuwMC3Fek4J7VDrshGG+Pp1oKCRadzcLgr0BH4PS3byi1hQNqykJnBdyets4Eyv
H5du3YXoEH/s7lDDD5kyMdIjqW63uvmDRGCPvi/Ad84MZyQ1tPRb9herFU0ZLvHq
5uuoxVaznatbHFrO5qLOzZ1rtBWsLw8woNpXkr6nqbUL7J9viT19OoV0qJ2rpsgl
OmZ+FWMsWrTxofb27QV4gFLwCH9w4Ymx9cTwvVnanbi6EKegAnwaKy0YvCNrjF6n
z7X1pwdI7wfpxGesrD2nfnuATnnIhyqSZKsIOpRI70byJ6ryUO2uHaavKROlRWB5
BzOt1J0n8zBbAPkZa2QdvDYyZzvoidpXM6bHwuJmGZ4B1lfeFU2Qcld3HDgh9eGu
PteVHizd2QYbkPfnxnU0q42MfL21jJBAIRr/YtMzMaczOZ06JbyAX5wtV2CkAz1B
QMpPhjt0r9QNy7ElnKGF8rtOLSt/6uPfNm0R26CY4n7N7prkTYN7Ye0fPc9ieQ6w
Mddr0W5yZ2JMmO9TWNt1yDVSfqH8tRy7kF3BqkX4UXHrfG0v3Y6f5tLo6v2uUvLU
+wvfKNflBjpJjUZGrgqVrgrRDDGKPotIQrH8PYSIvHgKeigvm54XeXZT6iO0s1Uz
GXcr08TSlu1+mBq2j+Y9ysq8Ys912gIeNLXtCgSiUY9vM6K1Qwy1MXvRxpc16ZSo
sS6TfbMgyOFdogC6WKkL0LC265N9VmFJH34HIEvqp8GbfFt38S3gFZ9SDzEevgpd
MTXIftiZDi2mYxSEsIcgD+bQOqgFHVBC60yJZ1Hi1RMM35MRz0cO6eEpTUhrCxai
pEWuqMay8/sNxq6Kfa8QyWGcGTyLdKu8Hov65BoWs/1qoCw4MVu6uyWsH2DHA4kr
CCUvBuzp32KvUPuK7SXLt9NtzpWSjELDjkHdVWxCtpybWKvdzSGwLgMyDXQJDwTl
Xw288BvtiYivAE112Ehk8MRj9BrN1FWDTU0uzkJb8avMjrONaTR7LL4kNgdcSDnb
H+Ew07hKy5EmnMTdLM/+IxSHuhRH1qWyDrlv3FMusLS9JLjyEuhI82Vnf8SmtW34
dxAeSFiVgPZ35TV0scLEpsoQL0gkesY0cRVWqYNE+yBUJPrFyXu7hKc9ahCO2K8t
bUJ4y1GS37fDnHAMKKgA2ik6qYedK+35LCmFQAqaq5zs4wZs0Qi+5WCGqfvxql3c
l9hVShSs+6c6nBJ75veHPL7yeW1U/dibTqjRtTFWRAaXj3RW76U3WmfuIgFGl3Fl
jgefS3ez5Ce92k2VOlToW88Mj2aZJL7XtqVDQehEbmc2lCw2HKKiRqGPHXCW7m1H
KyQsBAIKfE3xsUEB8CWf99La2eRafqwVBvXdr/BP60CMFCD4/iHWteRQNyCl7Q+U
tpMToXl88Pgjh5WQMTJdXOMf0B9TVxLTzMiLhqK+Znx2kqyjqFf7e2mHKURF2EaN
quJaKXoXsWX0xFAVdDXCiCnIIl8xuPrSvDr1jawo/NXfIX0b3y9s2Tn5McHGPIHP
iAPxpFjPJai/c5RR30CpqPR5GDWz+U7usaI4cfHUUIsiK1D4qliCxTM7gkkUandV
Hvbz7AZbwIiH5KR8vBP3yF1aj6Font9/CS7DwLleyc5wTe2HI5u1+wURk+5zKof5
TOG2LGmxdN1i98OfvOVGWtsk258lbO2FkTvme1fP1HNxXJdt+GQY7PFNaxeGYz73
2HIhwJrk0U4hMc0mvQHQQzjoQoKOSX9/A9hAPCskqkvubJl/AXZq9QLhYOtr19k3
ZRFlwoixoy20K6yPsp4tZzCyKOJ5iQYAbAAr1sirLVw/QAHLVOJkTUznAs8U7lIX
uYSUGSYJjyvmFlYDR/5/bwDVs1ANa+TBTsp28e9bUpZD0Y+YrMZj2EzA0XTuCUdq
4JbkYkbswOacUiRbkjDYlp2JJ8ZgNyWcqvyAtFEAaRl0t1ZCJNC+AmqiJeY/ovD0
pgAF/lm1tAja6e50Yc0rrTcdMrOM27olLhCIGWSqiO4P3URSHitGccyQHI/Zb9Mg
Gl0nfB48X6pedAeCzrTXf+Fsg13/CGrl1rNB+LDRg3TAMgdj4TG2iCw1EBiBOwaM
jOOMSlGRSQ9TwMeA65qUzu6rApvmMsuM2qngd5rtj8CyIL5Hs2e5pD6lrpwI68VG
hjuHMBxpcMud5TFZOtw9GP9DYWOjYKvnO4LuoDQRxVGuoC4MCrvpptSjWNn1IdN3
0Q2kM2eAkPRBF4Cc5dcqodLWRzOyzL1Fx6llYsw7HaAX7buUyuapv6bnCDkJAfeK
lzllYWjArfHyTV7nLccIp2I1vHXxVguhWFIj7PKZ451eeklDdQ5eKpVVfHs/ri/h
Hw8pqXkzNirXAa5/i9QbuC/OIK6spWgIuiX6f6JRYLHB7p4bUTu/sVtgoBSvXUnY
NbXWCzgskwJ8TT0twVgy3xrwanR0D15lZn1kr+m4yTyY8jMc+4FtkbIelFTMbhqh
iXwkXo4HEdGjRU+HGFPh4SNbFmJ50rTCGgOMf2ndwJgGLIAz/6XydQewpQEPUmcm
VFMzpzN0T9bDlkTCEPvZm9gZk2t7wBVhDIOqQFFqcsEclnZG5726HPnrY9X+MYI9
iLdD5yhLiqo08WgWIl5hYL16v1xCrPbnWI/APF4B4K24Dsvo7QiE9+T5wIJ6njno
DAtkZBjc8hXIUPO2Syo2wWrgV3tKgh24qHfIYPJgkExXcGbhbxNHi9+mQz96J3dr
h5JScqGHhjkdP/cl7XJZV/fUeXMhuDtwsYg9W8As6k6/09qo+84YY/GtE8dZdHmh
xDeKquq5CXNPBAahw+EpC8ECeSIEfIMNPwbNZWd/X/y1SDOF6/NAa9NjnnYbX1m0
zSERiXxRfgs2H+d0NzEj0Vdj7paPrTOx4sObExTpyypbEs90pWPWi3nDVQSNf0Nr
sO7DthEmC23b588DRHR5MkaaPkredn4OPqctw83Rr7a6XB79y5MHqVuFW+9bAvG9
UnpYQhzh42BhtQKi8OfJvEMGKs2A9LpL7zwK/XQKCSLhs1mqB6zMs7AasUoybfws
Xi/ANMkh87SZKUVeuvys1+5X1kTecAEiC3fVKYeCdS/9zULOV49n26idknRA7Th9
oqAyZrR3aQxnEuzoAoYA+r+uSv1Ix0JSrm9C5oadMTFCTY5l2RFm7gCz4zKHL28r
r4vbeD2AZHFyXLMxHKOXAkENgxDpMLLL/tYoVScwzg+paHE8oBn/vMc7YzxmSuGj
pr1bwLdmC//WNHVqV80P2SsFFXZc/+8N7Ti7kEckIEefxigCqZ8IeVFvULWIUO44
j6lsoj8CDoQpgR9eDfg8hBLgONNuJb8Whf57TGkcf4tketSnorB2GOeeABTD3lrb
l40UeYb6uLJ1HLXBUZVuEArHk+THWAQ3JlggqSLrOHLBR1ee5S2SMxbeW2Gk6lyP
PpjcUgxLxRWm+Yomfqf+2vOghj8NSZXkZ7QaJt69jxIfnfVlPkgAGUeD/wYLRk9N
gZZOZmxzVp3cJ4FjIGn1CD9mHkCOpmjwueHz+4ncC+a32/hxw5JpZinQcjM+o37Q
WhhK/EqZwgCqMCJfeEMx1g76ZozQyikEQBcjOsMt9Ns8S79ie6pkU9PgpJNmKwYS
mhmqEsFrrGg9KcGxj1oqVPLWX1raqlMVNvfupQGfD+fbWS+yniR4sLMd1hM2WnVE
OPplvGJqNn7x6B6gJtRo9ATaqrW0sBhp8Rb9mDIcr1bnEEHMHvq4dhaGAGAbYKmM
HjPHf8QBSfneH+r4GZak+WnKzfKAVnkTVJ9jX8/mw4QyA1awL7ZlEfGrnqquGZgu
gTIMdzKiqRytVTF/9stkN1AwamCzO7aIrj2tXKzSAucD64CsCkp23LQ3snABFl+E
c44DSPYv1IRhO8Z5LJ6uti8jzI36/VyBiC/XNCCj17Ov2lLKmfwTmOm6v3p3U1om
koM+iCFhkDqRUFmeghyGY0b3qXnbegmVcGJYAL9BX6k3xH4cvDIX69sXm8WPZ7Mc
Q+QXfKMrAuz8XJO1s8adbyYjvIQV+IQAHhb26kIjTAGRgEa73La6HklmPjcPkmq1
VDm08ZZcMmB1z9C01sBdollXSYOfGXOrzQZA0iQHKv4u0zT6yYbZkZZ0vYuAmUAj
F+5PXsCX9AAg8ODZE91JrN3iH4ZFrYetl9tWiztkGapbcomyjrgY+ZfCRigbFTAa
Dni2r+OSOsa2HvKNYz6hgK0HiwNvtkKUDSi3Q38qIkYa53TlZQ49DaVsfGhas0Zm
sdLGOwF31g+sY8GtEiM/CCe6AOIbYRvbt7vBwlo1cUn685mysyl0uuEhnXdVtIAW
KyKJiRGeGRumsir5l3x4wcI5gyXrR2ASBHjF5KtqsW7Tqt9jLAIfvYUI/GWho74T
lkgw/qRyiGZek2USDHelBD1LpIKgf1NS0ORoWclDUvbn/glxJJAfGGFTefTbP8yK
IWjV2o87oYIuAjhuZ50zWRMFOhS/rPy+zHBW9jhPHGWqLl/1rWVEEoWeIlt1+qJm
KG8q3bEZvG5aVMFz7li/qKTWTcPQ+88mukb2al5X5IHHYOXrZe//Sgahg7FjQZdU
2vOeT/tzqWgbkBcWgCHFQ6fjlw5XSstJymBbMTGNZnUvec++NuTc5yg+BSlaJZqN
9jxATgtKlHz/BWHIOPOD/jS7jQXNzwIndPhusIVL9Jfm6L0USH8BbYIaPi4O7o7K
hmb3/4JVLfhgLiAlc4Yvh17dqqfRA+/NdriKz0C5IoR0R++Hu6PF/2kFhvCoYyaM
k1AJt5E3EWuZXQE5J8RHIaY0xVcQR0022UgdBvc/f5Z3HU0//saGskt6ErytSw6M
HEF+WFAju165lG3amKQv0iN3LXMZSn+plPNBVkCOPTOC5Fha+S9AYN6w5PkULIq+
8gnG276nPk1udbJF1Db8TrUC+Y4LVjW3XjyP4OhTaDD+YJ3U2nKwFMzpMjL7IJ5L
7OgFevn40f5asX+7kyhM+5U7kq81MRcyUIAX96l6hC2B1ufPkXVtSjl2JRNo4n6T
SUxf//UzHsJ/7JbOYpTrNGfORip1ca3LRbNM3b8UPVqzI52WjJ3bVQ61Z0EBBh/Y
o+x2+YQiCRbAEP5XAY8zIJWf4CKpBV922X8Wz+kbh0Gbg6M9/PIdXthulWW26c8g
HV/cNYDKIYx340VfEk+4dbtxtnhp+G6sFNqODEQOOCECPjoDrVn5liYACKSQVvw3
s8MxWHJGuxaEKkNMWjpEz7hsxDw/yGmXGk+/mYzOuadz2V9gzxguOUazZxEW2pCO
ccVaZPC2ShqhFZlU1ovk59IHos88VpEDtmoxh6rvs8E+/b+PBHXc8ZWCDksWHNMP
LDf8o3w0/WxNG4Aaw5QOmczyU4vPYYMY/KiKxQkDTd0HHVtIkhXZr9UaCydqrXzf
N8UpWBwGVfYePnCNQR5MWyCjKmJSURr2RaExEb2pPdo1HQcLJhvOSUI8HOmoqz2X
VrZA6d52lxGQBJYZyGELgr2kT/3rkLmhjgjMkCRqYsjdFctvLLRYwuOhyFveEUow
9se20MqXo16zAwfnnTMP2I+aixNt8jPJeGOvUIR2CAK/hGxcWrUl8I4UatsURFWx
ESKCuvkqh3BV0rcf2wjL8WJPCHq/nU7+pc4bf2esvZvle5FFSGWRMIpncUPIiHoE
H+3jX/z+B5rPIK8DjZl1ek07/9RO6Gtr+RKyD2lOf2Cp1mN0Ple/JrpJw0ar16c0
XTUMnoooLD311cldgIwhImOQnKdIoNZfm46NCbTFr4PegfXXkrjI/lCFylqrt5Vw
MHqy3x8QOlFpHQxqEcfiq8iLE8hQm6IVs843AjuJnZ/YsXZ7VVU+J4PWh2n21g+V
yDAb7AXXfi1GwVbSePuj6N7fXV4wCFiShk+6oLDf+l3VYiCTkb276lA0GrVNvZGs
ceTgAYEA0ohHOuBMeEI0OfJakSTS2cV2AF0wNY9/TS3pecbXYVGC/VZLx5U4BogX
Dz6XP6ate3uxMG8k9IUd0hlVjQe1/ON2NlU4/6gUsSkWb7bgNBscULohNSkLYq/+
upjyvahlH3gIWfl2SsEHuzqZcfECAUUFg64z3EuoIKlKzudl58Az96TInQUR/dbq
nxJaGBfjZTDIQ68TA+Dho4x/ZGQ809n3XGwfl0KNJXd9oTHqKHXjc2BMFjlu8FuJ
cHl0jCtjNOSZmbisFc0GpZmO8vgv4emyNdpOjMQojB5qADcQ904Sze+qHPI8hC5B
UXqqtyRLUQ3Q3C8w5OAWhcp7EFv62nVPesDCWEHf1e20CvzoYuq/0uI01OP90TeB
8I6pWQL5RU3HjbuBSr3elMOB1TOB7li0QpKGmxpvAdOlK/TwR85A1hnLAVdzqzoh
IYuXMhxz4R2V4OASBPexzd+je2gI6R9QtSr4Zpj8bRQLJkcFl0oydczg+4f3kIte
K0k4R7AJtUre9ie1aua98QFWatXRm4kyrIDVB2s4U/QtjqzLkGxZQxiDLUd6zig9
UYX8WP/C12uJYQSG4AwQj5O44OcrRudIskV3Vh+cPALNBGeUA4XILyavjjwN5FN6
Epfpct6St+bqsvGiSslxHXs9CJxKJmJk3Ejji1HQTJDT0SmXxsu/+8H5lr3pOdqL
ti53GcIbbdb8udLNYkI4sR6HPOD0b0U2IpjyaKESaPRIy2PV4fh6Yh/DY1eAsQZy
CxijmRZxmVddy4ruTN5Avi1C415q0IPaUZiALrSKU2qP/Cwo8M083U5QIroeSbnD
B3DGva5aX91ArFna3st+bwfH0anskPeeurRWPIr8RCyC9aOYij98Elo0HbitvDRs
IIRjZ5RvsUrd8ADmEEiGd4fn6bYEb4ggaeB3UT3y36qXZHMMAOYk8xsASv7pf50B
Br5sJ5j29MWo327NyQvUnVCkbmUEpTFIsokSFXOoBzA/qye1ARim7J+1l/LIJMEm
kWaxuDqWuQbr5TWHFdY78hnlZDl3j75Pw9aSv/z//bA+HgyKLorOpX8MSM8OYroj
FS5dz3JNILIB0Nfm4M3vR9z9RYYLT1hW/kNbHcrbNHMbPuBN3KY6v2Da7HfyH9Sm
QUMaiCeCXoSGlJxulJFZ7wyD4c5edTl8JxLydUmU4kVoxWtpG+BanW+8/4a/NqTB
91QcMHiwzuQyBn8hWCqi6VL7YAjtcnOLH8LLbH8kP5wqe0vOerqZBgQcLCBMDJIu
T6tEaN4TXM8d5Ev9jkuwLXv/VZC67MchYCunELlIiwgkRLm4EAMEQgP4BR7LHjMe
KytNVPfrLNcjoskz2ics5VMZkF+ajSQTDec08WVrUT2LN1oMAsOc+Us0lYFIi6t2
Z5CoPV45b5Q0/CiMl6cLqMQFjXfs3wrjIYmdPjTBkydNscKo3c2bi0GOjH6rub0n
hoaRAj+DgWjsh0E17YnbU+EqquRx/QBYTUPobYDadwDx/3gKsYk+HdyfZjV28VJh
L5oxDv8wAFfSJK/mygcpuV85uarg3b8XuO+pB1YZ7ZVkcfpiySFF3/G+bWtiv/+6
5fnDtb6DnyG+FuK7n2me1RiTi1CNNd55q7IT1Nhw7j8Xoib1MWdTQljasl8ZgVTe
t+EfbKDMLpCMnOkprWivhidPwX6yF3h+jXS+5HdGVAa9FoesSWjywHBAhpe2Z3hx
eSmINbe+nP0a68gDsKOMd4b+7HYTJd5Dqqt9jA7dM2+ZTZjnRzoyFa0IXyVG6VKZ
amJtMnnSwa0useMpezecPnKrh0uXzcuLUOO087bGcmR3V6TfonS5JNJ7O2u2bNS2
MiqrhE6hkWYewHi3ByimwEJeY4JaMs5IhmxRik/9PYR/eSYkbowOMBN/XwenEjk8
lGWBWe7ulD0rbGP8h0YqlDk8RTEL6URbwlXZJHHYC5gM303npHZi326Un4VvdEQy
kWdT9Yk6sWj9n6uyvzcMNEZSa//mUvCv03DKkkp+Zg6bHOe9dVTf2QIqIi74Ibuh
KwWdcQ7sjLWd3rlZoMxelnrwmc/wOi4QZU6M/M8HvWx4QBjGhpTuj2ic+vOaIrYZ
THApkRaoKVQc+KC2ZpQnXzCnoTZ+7aQx9JOUlG0F/9wE00NE1KnfgukeOCS0W34N
Dyujs47mu6dSxbraQkG9WQJg1okaByxG97iDe63RUpM5D0ruKRf/n/tIqbT1ACxR
URpJXoMtM5HIgcLwbwIuRjKGxbYPeJRuNRVY6BRmkYFZWbdpbh9kNlatbF4Xik7S
5RfOeM1JU61z4Ubo1UMWSpGNkmXij5HHUDACp/pBbJ3kL85y0G63TmjkRI2lGfOF
4IxSLNV/Uq2eceQOVnewYJbnQqnZICjdbqcFTUXBLAfxG78HlSzRkvf7GJhvQD4B
CdHk7n7K8ySxIMlq6MsTQVq7obchhVKfVrDgO/sYRCF+1KuFPC3PwL6Ojgwghsew
NU2Tq4QGZh2CKHIZxrrMBxGM1KGZUc7LHeNHN7je3cxJ3H9CL29ATY154Zy1rpIM
0qet5U7/FlNG2LvX6px7yV/lOq4GlBOIl9UMdJ0DQjrFpHXepe9jM9+ZWahv3VD6
1xW7HaOHca1AKq0vltiDi1so1JITCWCJoIhSollPFY/fHpluElXGl0e0WAR+fXdA
M2f6kJrXURTdUDnvCfQJfikxDL9EFwtzrqrRaLlSZ3VozwtPFEwiAzpwF5Rhy7FU
LozcvssOlNYpwAmZq/xrAAJh6iI/pJFPYZz0EsE99+u2vEFQs4A7Cqqa3p2E0pYj
rooLgK66V2cRgQXs4InVIzwcgYLxAm/5BpSjArntfgr7dUDPbM9L1mZAbgoeK1Rt
Uo7ZvE+/4/zq3Mk2XrN7siviPvktR/iTQ8yIhAnff7Iu9/fACMpGIHIEQm9Tqymi
/lFdVlzbIwYuLNxitOe5XQii6/XameqPOoYAb/utddxhxjlQjsS8j0QAIJNejPP3
T/y2FjHl47I+5yN7CxD7XJTZH13iqzW3CQ5o5AEsxvX1hTfqC89yZT/MjtpPaSID
a3NYmfVYryAIWOlAJhSdAXjt64mA2fSrTAIO66Z/fGg6Y/2JPybj/m98B/1gZgE9
NqrOo4hqO190VuNgeyllDkRofcPYGL8KYknGiE1/kg0qY/96W7J+ckmFQ0SZtoUm
YYdeimeQHxpt7IIy9DJ4WD/iRWCppfOKHKHsYXxZRp3OoayHhYMS3kzuOC1Fzd4a
W2AtQfE8NyTNMyT4jNBSvbmlNKBW2+ozjUDazK3zwXMQYgZVsx5TckqtKS3OLL6f
Ie2U+mCrJjnRq+IGnthH2z3PHq31QxvSj4IdCPqwKvB5iLzkLGMw8iHegjhnvwyx
9lOcyv0hHztFlzliTjALrvNPeungaCu9Zyzu8vyThOK3QaOkB3Ot9uKRdE83zTXT
0yHdgfdFjEtbKmhBYpRlfqHclxNFanKLGtdUvvlhoZL70pLiJVUB1KFLgGRzvwDC
hMRTbTRzmeJbNfFDqUkRzMsd/uQkOwIMFdWymbl0qy34ewTgY3o5aKeLHQkI2zNk
JjXROiNZ0JMPZo2Q/UOLjYIeVU+zSv0PbzZ+l2TKlIxumY522oH91v+yrL5DL81l
9qvjUO7M77dG98FIJ9teDU3XE3cTy/f7kBiz5SMMvzHW+1MN8v2LjAEyuE+DQPyL
yM7z9nrkmHsBDE96gUhcLh3H9xoR5xBJGIo4nFJukUCbHFOqUHuePkCUj9AWxao5
l72RcxbIrAcw0tqZQmxktNCs2zYWmGj9EdoyeLEnwgywx1QKZUKXDHaTn6/WNNBv
mNh3d3JHC8HgOUH4ZBBIQyPpcnFg5BoZ6w5XH7hNsyf+dwbeg3uc1Pfr/Rmt12C2
FyTXQyjIgnK+PQGvoIJ4EBHanWJZeLwO8Nh6A707xklzKMBUrPG3mdVFcHqEfaxp
jFg4BIv3l8+9OJj3FLxxRnJl3NObe6WV9zavddGiDjXlTFDKIyI7MYmra0O2Imx3
vGtOdas2Fpecywk3taWzmOZ/eDd5IU97RnLLVw1twUUQ3lmoC4jSmsNxegHAUM/e
7a+HsKJLXR4ZqhELRgaj7OXAs/sOX54DAECtERZXJqIfjBQ7QVso6V8jOVCYSd6C
lfRwIvWL84ezTvtU7/8O9n2jlFBnG+f8k7IpCvLXQMAXGxwAS3365eXXB64q8di1
Dq90tP+19VlaZhdM/esR67T+Xb3zNf20DFNK45A6Wmc7t8XhSFSiLYhFD4qQ1U2r
15R9z9PYurUzOAPYp9PO8gAx7EqeT0IXa4dM9Iq5amtTB/RJcMs8/FWYS1yzpHfP
Z8I53/ADTS45EgphS0a/rlT+GnrSVsBihwUaztD6O751F1KQJZY+OVBQZTZaiJ8P
1uAMPs4mIkKlAZemO+me9CmuRmB8CjBkJyRdifzpDduonBa8AYIiT2Qie5nG7203
caCILhD/f68aN7EWcOl1zaMbNDho+txvQdkHh+3BLL5g5Q0rcpPrAjd4ikA0/d9t
zgVuabwdV88YlHxWV764MTyb8I5w8hWxM5VbOUCFbP2730Py19uTpEv4jyEZQ3w+
1A11SxBTMeN+iWn1OKoJcb0QXAH5b3leq6mobMuF9qgVWfMF95lLDmUpuWpbrYxA
EYgdOlqMkyalNhhlIFboU4+R2K6W5il1Ky77dtggPrFgxaqRtnRY8//bcVwkjiOF
wXxz/raYPEcPlwS6Ky2gV7u7mkea8mfcX7rxQ240/EZsNP3COHw2EoroqclCjDPJ
n3EdbyKHOX94d7wbY1yy3WfvKeqJq2cJ12K3OTedTCt0DYab5yEIbN0rjou0iG53
5rt/YoJf3VtrwxsCLiTlgxfdQqRWVNyHgOmBfNnfYtrERjWQs+lzP/EDiDKDcoeA
hkkAp+UigLh2fwzew5fC0ncmpAC0m21JhUZzcczQ+9hfyKWQ2JZx2mXberAl79Tz
c3sNm+/xHoAb1abjmtHla0qfEHP4fYu0EO/wJRkRWAIXbLF72cup4AjAkM4Jxans
FtcbX+zKV24FocqFxjpI6FwkSrnNeJszxBJDqYX3FAZOaZU6OlOlHdk3QOwZCql1
1vXgH6GaynoGNwbHRczTPD8/U69c5V+jgD9niz+4WH+vCvxCC6bFbFzlTuLAdfcx
82ew+HWhnzclqfRjFKMp4utZWeGYbmH1Prrk/ya6pQQIlbcvF4wZ7THhE9uX5h/6
9CrGp9/5RTkYJyYpAh59Ag6Z6+Zp66lkaf5F/rU/KAoJsYla6ifCh/SYCbXO0P8t
mUvbUUZuXNNOTZ32PplMSQW9tZ8r5TBlQf2wPAnEkJeAokH9YxnjFcLfJoRC+pl0
w2z9hLJJ9BEP7PhZOliE0uPZfr9sq1f0CLaKHN8zKXWrIO5wNwUaSxcamCEcNpT0
S65aVzwiu9vmTupmK3pZ1hjtuGG2St+z8aiNSNdmaGrb2ac9bWayQAduDohJzcA1
iBm0tgk+bX1yGzjbgCEuLrvqumiH2ukVckycfqPqEt8sNapnwNiBqkSwOv2ZhcP3
u4SqYOTJnmW4GKMMBura1nP8bJDTJz3/HYXfUPKJsaNNuQCaxgoUceaHCHDaqiVQ
Cw81SYutlikz33MgNFEB+VltnTETKsImjbW6UHzk+n5GBXDkdGng+5VWusufr6LO
gn7npznQhi8HsCJICfIkC0R/drGeLZehcY+UJPGqfyx3uqqXQTRajmxg9ICHvSB6
DuZ1zMdxrQep2mmls0+u87pcxE0A34UjFkL4gRJ8SW9szJCWSkJEdF9cs7M6eS4F
MdMaPehLHZBmiz8qNJUU7AFepwIke0u/Iedq+r4UcNpffPlncsziBdz/yeKaLhYE
NLLpx/wAmdoXcCtwPSTowc+jNGkUjfQ4JZKJLrzds+RQIq25/CMuwUcCRWnqTMs9
wtEfP4ROafkWQve6g3g110YBi6zRL2YD86HrysFLnjQeEothsTAXo+XThpJLNZRu
N9qP4RjvHThfQlErvzuErOSUGvRBVwWidsun7pYbA0Mw2tExYSzsYDEf26pkRKQw
o5dshvIOBRcwtQranRXfaDnUFTyF+lbtu6eOKA310FLfc8Nyiwl24Xfj+gZMMSIe
YSt7yHc3nPFxPvnNoGsRCKJwwmXdt4Hw6GcozlTOHky44ZnYP0PUuv6k+9M6sTwA
uPzFiSsUuVQum9cMw+aMfBqvGzXtFpGfNJzYgCoCGLWJPh56B6Q2X0fXTxd8qfol
P6Xm6RXNrkWDOaFj3DuNVtGau6rxuHBJWovkRsXaJdmfUGGPMSs3abwC+Xl72kA1
6A+DlyBNWoG7aB3/RQy/uJFjcptq+E7GpoedTqPKGHeqHGhYD5OU2aYkLZ2SvuCw
a2YY3Sk72F4EpNxL8S75/GNFwjYs62FMEaZYWl0jjicJVtA23qkqwqD2q8ne702A
VO3eGoa+ySgfEm1AOffVLjP1q60mwNK3zDBJmL9CQAl47EghCoTNE0DPiTWJYDsF
EWu2sucfma7OxVUhE7KAOP3ABfNnlwFpzP6ofvQlfSSPNdZ0p0ck0qfNoPrG3TfR
KYTIkKqMVjO6HCmULItiiAHGV8MGzz/IpjtGduB5YEeX/ShMA4HCUuiUj+/gcDCK
L5TYo94up/R/ZOPase5Zgd3WoS/XI+H06ddWbD+64iwr+vsOTx5ko4CxziIXX4he
k3njUJ0QlZGmZmMCPbOfGEH0Dqpd60q+X/YmJjHVhkG+y5Kl+J4CxMFVqjK5mWFG
3Wy63FtoKGwRcYJyuZphvLrCd7sk2EcwqFC1ctTKTEfpjFeW0kc0HjJpMLObGj0a
YS+aeRttUUGbNxl9KL4ux/Us7+Zk48nIc99cXsaRL5y/AxZ4cxF9Tsyu3VBlIKNA
cTY1fmSjtuBpqjGVBj0G5s1I0ZzfU27p4Dym4NGVHfmznAfYnAzMoz0bATXIFVlN
8i1ySx6GPfoEwEzDvxofOLbMHU2KQgbB5Yhn+VY0lFflCI5gJCDwJ/VxZtiESa6R
0BFNvXxa1hgEjfd2/Gxmy3Gej9DlnJxjvDAc8T+AtFzPTmYfiFQPLItoKT8CJ9ZI
rXITextJxNu7z/s6myLQlj7/7ER/NllarKPGXsz9r+xSaOefpMcIbtwn3cA5mCsp
w/Caw5GpqtgF610cpok598dCHtxHyrU7GhSKffSsDDEIvAKZTlvOM1akBJ/sNA5r
puyrap6z6OyVorh/ErE+sLp95NjiyXRIHSxcVvzAUclIzfnWmrNQTsWQAeMGMwdZ
beN2Ya7KvpzgGkENfn4fLV2GfpsGoChklUcYHWeCyTVVpDN0hEBEE0pj6jGASZNU
5pStmi0ufr3e8xm1HBbt2aax2+kEstmLNCjDzBdZXVlhiSVQhu2zYgoEZPvByA0S
vtcIFfzdcoHW6lnlDuEi6WvdD42PQ4LUq6xYe85mbkNAx5N5xQBbCikkg/Q7V2ov
NFMkA6vTM4Ld8a0e/tYocagVTakk/aHAkkhutpwJGjOkz4y605GgcMIBGwqXT9av
lJWtYaIeAqizZ0DUlSTlhu0ncIWrFFfSLKlrJ34ff249ej/BoOZ2UbwaINQ1TNNo
QuKOJg0Cd/YebZQyeSMqAnQ+A8Hqg0R0Fs7ngcnsblE1pP/MV1tZHzzfyttdLgVt
2HlyW5ce4WEznCpVcwPECA0pacRLFXk/WvHBuLT25F74hA/cjvlKLt29KOxYAB//
npcHYkxN9EV2QP4oaPdG4a2HUSeS0wx9Pg3fB/3G6EcCY8hyqE8KS9uHEKaem96q
ZNdk+2skJarlMMkgg435BlifvKZVCfhZhTBCgjB0hyXFDUWy9bxgILRHLdaP9xSe
QVqvGjPjiIlp2BiaKVzSjJYHBcnYlaYK+HxJWFZu2Oyc+/2l+Re+Z8QjWWPtqutw
EeKNMn/LFrjsVJ6iddPrb5V7+aVQzdAniL/Wxa0n2n062L97bR0rQqS+FNAaxVAj
D2YhUeCYJnF0jpMSLwb7t71lKRo8vM4N1R0HerKYdhzJIE5yw3w34fr7mJ6tYAZL
xbFKgWgIZzj+Xb7VnVzDryMR9Yp8Tdh+E59A74oT8BeweiiTVgF+j/4qhQQyaT0A
KUWEB3QmJWtb4OqSyehtidMlGrQqQ+/fKKfxj4Zc454Y2/vwXaYaTH3WmN8HtrT+
SekHtk8Ym9dKBbFeZfuDG+wV3YRCniJ+iApqsM+rEbs8L1NSCTpZpBZ+mO2Dx+ol
0IGQaPl+P3HLOgIbG9ak+sh1mzhqm0x9U6Vi33rOGE/KL/2yv2FSSPijuzpRAbps
CN/2oUWLrW40eAnWvTty1bf/4w0dd50TFSJHR4+KykMiR5+/FRbZ29emAbSwkssL
veuUx7Rcl3E02CdmQ6HUBpqJcxY2GWaRjt4gy99Jfpjt9zp8557quqJgkOG/Gb1B
vVaVrBS1xVye3f+UzuwL/qotK/BOLJ96NV6P/F+WGN5uISPOxGO1ab7Qv0sLz94C
Ht1LN7Gyn61T9bTD6r2lvgY+Ur3+zBWemkfzLdABAiesildbE7ZhmRp+1YuoyuIL
0uPUnP7Wnqr660ccA3N1Jc+nrd4jpMnCurCNpctDGlI8l8E3miLtvWL5XRSa8T5h
YUJscXASqsd3RdVruwU9ii26A7sZbXO+nTY+bkG03HkoKczfeVK2hR7Ptae7LNtV
Q9DptQyWG1xlc9SB8Rua4AwjwtvelMcomX6/We7S6Cdv1Stgl/O9NDrpKvdAIhf4
KY6Sjh5LZyvQsdmGoHJSJ8qRGzqo/WObScXksYIRcFc3LH+2sAJN2fQazp1R8MV6
3g8u7nVRdd67EaUCeh1cpZ8ydiUY0M+CMTiyb2Qn0p1urWsLvJb9OXv2IQDVLjiU
NH06fy5ljEiPqZkMh064hxNoRx5K3RX7qve/ADWoaWkRDJJkqi+LromG3hsUmJPq
EetRdXEt7fDr/ulEpKaeGSKPBCGG+zo+gg27mYo8MuQgduSk6HPEgGKNhdcgOWYa
L7hqM1Gil2++EBE7UGAq0wyYtXJwNbZSR5L6Q7FY8fNwxZOmmK9vM4CZQflngqFh
LcgZw9ZMTATgMo9rqARwdX8dGoiUqS6t7hjwBQemJqnYl81fgd6hpSxQ0Lho59yr
kLtW44CMiR3zv/qhu0lljtO2S+6sC6PjGjQChlH2EtEDxFvjYEEKoOijgYZ+Przz
TF21HOZcpsUZlzqQkem7gxDOmbVNIXpHnZYfktf9sN6ukTAzSQ+/a5xr9AFgImBd
SgE7zez2mgZdTW+4HPqiWGQ6XT183ZRW5LZRCtGeFWFZVuOtaqH/IJj4EhCHXfud
vOeBYl7snnxn5MyurpdpaKjHSx22q0/nS/Qr5LKCwGEtY3zyq6wC2Bd13HSblsF9
+kRpzejr17oFhhVIjFHB0RIcc3MOdFi5mlFBBt14/KRlBo5lYOpIlfyVYS+knokm
qAGWJ0YVvKoaBlKz3liC/LQFfxOE477hRe0yTXKiLN7iIjGequpoRMbdgf1qj8lF
4W0XfA2QKQI1K0dQZVjB1HJSPPxR4lywaXnmFJPJgP9J2j+0DkreZZCzCGKOVECw
6cYQhhNdfNtqPPiDI3cPp7MQxroRK878ob6MZgG4/NHWU80bRFcixXXXFN/gusVR
EYqBT0JGuj5y+Mg/ynnVa2aj8xgDxnBzynkXdkhvx0OoCkkIwKhnA6EtGWe/Jdw4
mLMZs9sVuZkDH9O/jGzYbwEKxIAeM14LaH6O52G/ZRpkgyzVnGyGHk5t/qZRwz1K
fGirCaEfPCSBha/iMlgv5yTd3PGH/gUWk8GgZMqLFyxKmI0KwCnO0QMeVwQgHl0O
baxC5Lf67QvfQWR4/LWZ7Zg12Bw/OqbkLDUpvekaWdiT90rmaoaKK+i8bmOs6wGC
MwzzNYzTcBm4MWSSWX04MVX//YTH6IoK/HEU3AdbMArJqRfwEFR77NCiGNhc2F4H
Vuba5Kcrebeellagmp3niZkEPevdm38FJpFV31RAfd3vigLwU5kaJpDQ0Uvf3MNZ
j5/owKftOqYaPZBTaicdxJUfWffufCTgV2DmXLFh/GammMLUVpEUzF1ehhmbRes4
jWZ32v7jrwWxWTQx02kXtAH8yD6r3/bsWcZE/4yFwHUuQFL16wVr+tHReA9Gw6n+
V+5SFqBEWeE2vk8ovYuAUJgdGYU5fVc1NDclPuP7n1tLQgcTytWnJKuCYBX2kOGi
tGOVsh0HgbHQ6IWpf+Txueif/hdIP12ZtDeb90ZNm3aNUEeVJIX6m7J0vjvyUyIx
fEVt2tQAo3WORfDoaCnuY+a9L+g0eH+HKVdali24c+I6tOdyaBySdJI9Chd0+ZQX
5Xej3Nf6RT+70QwigGz020eJU+kpfRYxBYNCJI79/DXkvztpF0cCEkCZhnw2H9xZ
0oh6gthlcbVd6L0FdfhOMnrW5AewwwDvu+/t2KBb8ZzrS0mZe6QwK64QAfRSLG/h
OwwdKLIhtiAAsK7AATQxZtVQW85t8CAUTyuwntjqrXoG+4NFh3p+uVT7Itc24QqB
uC6DfnL1FswzlXdIlO5aoSHUf/+UwwfagG+tkc/JO+bGGR667OpTnJtLqfl5kEbL
x2Hbgq8r8VhDs/22/Bc9bnAku+3Z0rp9dR6mVyDurfMOm3geONrUGUy8bMfa1yI/
LKCJYKBgLXzzJNknoUO4TRDq5weV9hyTBzKueByEQQKjRAKk71PWSSoOZ8R0WEQh
3cV2NRvWsrK9AMXaSvRZcI5gswfZwGJ8HjMn8WKtVT+M3FF7g2aaceFec7Zcd96v
cqXwLwcVkKqmYvT9oh6s2buUM6JpQwvnjdkyHXHg16+UmpepGRvyTizTOyHqh17A
NOYZxHX/Dm4K0MaFFQgBC2cbRKUyqm3+Ux8/9c39yT8LrbHHPaceZKC32887E3ws
gKjFME4+8wbcom65Re6G5iC4sUxY4+1JbbuRabqhXTmLMIyVNP5A6vln935US6Z+
hUWhNWsipdOub5gatQyg/PYUt65ZIzpAmjoy+aMTycg/60aR/jKAM6VBC8Ejuml4
ZQMba5LJ+L2o0iNlaRQJl74rkmCNWlRtZN33L1pafOtT0syvN9i7MfqcN2Dbq0uE
YsCBKaIWDYnTGWo8SjXVceeftTmCJikopgkfke5nTiApXLt4pTztyLgO1couu0Lf
2/k8zfJHIu3ehc6YgvAplkRYO+Zq2WW4qB1fY7VwLliJo+TjHz1T7e9fKjF1BjvK
CoPxVcVSLaOOpCFf6PVitGG3a/b4KNj4JGg9PoYWiHVYjDDG2TDHbfL7RgS2WWr/
QFel/IVAHhhRr3v/Ik4OcyQQNJkELR+8JV/WNBujOLlQWmnsxzogOmdMAR9vCAqB
sn3Ag30Rp43t3tHH800kUbOKbFhCfpsnVv2c6UlRYCqMZawqaV+hSkey7i9FwlZH
myiCD3gCwR6xc4kzbgZkam1RcirMBxST+m3CheVOsNlIiqjiwTMTqCEfrEoTGJ+6
zZBwyThxz3SCXdB7uLhGn7mifezjQwDMQDnS7OQUH8T7QqVyCTz/jCgyQogrh0gh
S5WtmgZyE+BVRHqdmeSnVYLpU+74jUDSEIRVaBeIpwxQ13wYcpeaiRer8yEFOowM
ZU21EgRem6LhDw1lyUy+mcm7Vc4NL1HZOGZKx+fnSCQpMjOeI1l8lynKOKVDW9ka
UrwmsALmlcwNf3X3nZ2D/eKn615AWElbba8TnAP1XVx2BJFZdnyGwrpGkZSNgnDR
EfrrlRmcR1Z0G60g9ZqUAw79cl0KGm+YkCjGzY5Fqf3mQDzBtiul+R879wo+J6Ao
tuTN7ljFrjwpfvF56h1Od2NCGYESs0pMg13m4ed54KRAz96S29LatFKxqzbM9H/n
/X8JJtfWwP62ZIms8BlGSsffpJPWXg2uqIqKhS+k+x58bn0rsk2lQ8dGvorBY7bh
fzjfAefb0pBg5TRrec8H+ZdwTwSdHPg3iNrRTzgnzBQsotUQ4eQORgfD15QMTm7U
uk8P1mh4k07a/9MhT85h9aXt82aV6XCwUlT83AzJPkceg0OSaryfHTxQ9rUgzrOZ
EIZ/ldf13OfrK8Q7796z2lk2E2zI7cGUoMhLeJTQXAGvuFT2dmFblpNEuKftbe2N
Zpurh9+vPixYjIrOBzLgW5QHwauFEfv0h6r2odadIBQz5vrE0cIF7JDBhE3yKGrn
ZAkObQyV67eOl4zKtGhd1cXI1YmWxBthaM/4ZB8IqzY1ENlHSUWGApLSAW/IbGFU
wwO5F2yBpo9HM7hVMyo+Iouw1Cj3T1pTB3S4yj+w2cuYbch+O4/Z/HhLwsN2eSjO
wlVGwkI4/F4pHQGkfA+Hkxymt3cUGOuZ8YKpsRfcST0RhsU1GuC322dU7nuudABG
pWZUgC136w3V810c774tvnA5YwodzTyak76kbBi0PSNSKjDIBXeSSFXTsL2YnVN2
whuNamMGWjo0xEOHADjfQ5GQOMNWYDgEHkbNsTk1hKmCXYBFB7BPLNUpwfxvF3F0
t0DwRZUN5KG6o7TN1pVOXACQlXULW3MtGZPUAJUEsZEwErMKC4a0NOeXjgJlRQcc
G9dgJ2hrjFtFgiwkyLnLSFL7VB+gkO4hXP4sNPWGaYabJUhlJWFEg12J4wTT7IBg
5GJt4meEbhFzOqtQjMZ4yIzalDhV/Jc+rILgK9GKrbk=
`protect END_PROTECTED