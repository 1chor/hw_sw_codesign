-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QGf2IA1kd6ZYUeYTwIIQuJPC8JBcbfv1qnEHyoXupan+xabHL9s89I8rZ77OREmt
8YozSjfkdCZWF24spIvxwfbpnR8GA49tK1DLp+N9FPycgmARC4/nTBs/Pj9gL6JU
aqJIjwhMtYiO3kSbPUWojKNQculNvWcpReBuMk23IDY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8667)

`protect DATA_BLOCK
j3xTS+9vRCPKm8oOcOGpswfX8jKBLI9q7jkBvyxr9Ij7Sk/xzoovkR9DMeio7j1z
ozFyhVU6cLUaVCdcDfp6WK7WrNAwBtYUPdz2FrK6uy8/PDKsgyLCSouV60xVGMHR
hFvpi5InT2w5b6h/sO7pyEX9NZPJCOd3bpUcs0hrO033wsn4OikStfu9lLU3eV6e
yGMmZkeuUSE5pXxkEyjDSZUc2/RUpTE5E2wACiHomjQsG+LfcHMxH5s8dNF3a0fD
yi26V2ivArsrBMjCfGRRGqaY5BnYkjiMKjSM0en8OIbb3USyYmHc73ygP7sbx95a
i89VIyQsTreNCsDpyfm7PvLu83LHcq35giVvdNSNLvL1jMggrzvo4aB6Nek4RDlr
6EcNijbFMccAGrIESQanE85DqkIqes6lXHjC3O1DEdK530t/24HR/kB4Kte1ax7q
qgQwvCCltRW3dFLC8AkkDWZrZR8xv7uM9+m9qUJAIxehY5WfZw6Kl34MMMZxbe/x
ZioP39FBQERavvDqtKB4pbn6n2j29WKIeDTYo7l9ByFvlank7uQs16SvpN3sVHfg
kXJrxRnJ0lAFm91hkqWGu5r2CuzioDAFWQ8W4R1za6zoA22B+LjdXOtCj+d8YvCh
2IJ/MrgiG8Oc2j5dS4USV7PXbHheoeNwkxoDnoV4k1/gb/5H5VHh7AcyP3iPTK7i
493YwTPppZCVIMGb7XWuw/UMXAtAEFBXxhwjFxLVwNVr9XS6lciYPv/AVymvUHOM
iN+ecVje12BYwFXlUBEFWyd4emGjwoR5ZPoUH1u3RJDWSbSN3qx8LAiiWHISKIrO
mavNA+um2GvWBFHWw45H6BbIp6zcrJQ8yrNFSlUkceJa40Pts1n2jCVxJRtNxmmr
0fxP4ErQ5hqtvGGm2q2YE1aThD+cTVaUA9YBtMDdjRfE4xzLRedjRAJrPTCn+FGZ
QFr3nmeqgDAkXVcJF2TjIg+j5tzyxGfs9x+FBtDIAnY5vw4+4DpLA/p8pL6oYW1B
HEiS6B5Q9BBRkkX20p8+9bxWoAlwnC+UfKgaLn0mYaIudbm0ZzbisRc/xz4z+cWB
4Tu5zix8uL2JySaCM4E9mLQtbZdGO2QkH6kLZGAQaaH3oAXOLsLBQi/0bkskpFmA
SCnrdipFjfRe+2ZfQGyiipIFOjDrlWLWC1F0ZvKxUK2gUooHpZxgrIggpJp9p92A
yux0gDhL7ts1rFEpt6CAXKKnSpXFXyAU3XVfqhtEthTWGzW6GEHOUE7D9rJHmpcD
/mRb+GW1hy22Hx6Wtb6wT0wil+RyIOLQjKXOTRqxGlFo5qbmwq2uGKj6rxKFyKhy
awDDQCtcJcMWhftgtwFzjV9+ktpVAiHqC/l40NzlkY99LRJONqordtv2Lb8SRnx8
y2127ivh+qmpVH1D9MIRmjO0mtfr7ZDqrxWioAj7BcSV0uboHAgUNF3SRn8aXPWU
p0d78ZIcMTJ249TM97EAl3Zbc2VmIuBdIFb9PWl57srCBof6tA5qXCfxCXXHX32T
d19YAd23HtsmDvuB1/7JFzfJ2e5Y8XOCrfEjsDdVVcukZd3VN72EfdaJ/QenATNw
tQuQx8MvnsZVbD1Q+j3YzpTX1zm6kKgLwGZl7o+rijcaqoQojlB1QG2AicA5DXtG
YZW68gS6VBz8ty3WWcsYx9VpoaD7LB96fgVS0BxxBCLkXXxyg9CON/r6p9a7mAHa
cOGIWlhnnrw+kgmlYhxh2tKmqV0jygBZRG4kIE0+cyB02uR0SwnsiWvudQSpAqhj
0OAKEd/Wbs/H48Ov8kmOV0SIC3iarAPEV5nUD8+w2tgSfyQVvLnnCVV6WI4mdKQa
Elkoi28DXDaUvOI9RzmcIh97Fx40h36pJ8pppHA/AVg4YCJHSJl7c0ZeomYscRtB
rD6Y9lw7Ud3cfpNj1RdjkG8muQmox9OjsRh5xFC4OmS9kks20cjH4XhVf4gyTIEg
SEDiqYMQAaZE9jrytcrO30dN09tOl4n45HHFxwniMX95G5vvQb6C5Pm6BZOo3C7/
1Vnfk6iIcC+ukCyCgHXCpcY8B2MJFOB60NJicXfRhONWwrcAL47WriG3f0rQhmST
sgLmQ7XxdUM5S3V3EqL10icTyQ45OjXZiHpKCu9xYVdJWYjrKRhyo+P8DE74jNiV
DrZdT5iRoVrjOG/GM4kXy9yRN6icetZHEPUYSglrG/+2zJozhxNDDrN+ekTXLgW3
ClDswExdrv0dtmGGRvIKJ6R3/BBjSA26gi2pRVvGcaXQC9kGux8XJ6WQDYPdELsQ
HygVt3YLauJJjoZb9l00SGPrfKPCNdX4tOp/UAklvE1EOTlQ05KBxIYN8MVZDqWk
jx1Jivev4K5BQ6F7rKxV+UWzC77ww7G58Vfhaep71T4KbRyHxpr5QiWSIX1tHIhU
rjkq6Ym2u8cAKTnV0PVRcHriW1nO9/sfpBr42vNpAmNGCWMriD/zHuf8viP5fGEa
9Q+PJhE1q9z8PMTw47wIRIKKTLJWu3f/JFI8fp8soYJGKyIJ6zX7pcurSYbR2j+t
Sn1NgctP2yEODGCa8fsbNwBwxQmlBbagEAb0FwdvZN1mxsiTkFWgxMGc4eIBpwsK
eU4J+JwPMiyrcSw0hUqNZfRFjMYZrcxQ08YtiD3T1RmIfZnt+dG3zOq4/gaA5KTK
cBZcwgsXOB5HSFC01RDgRATUQC2rXYxAM3FExAyWkLR/tsLwI0sy37n3Du9eycc3
3C0p+b3amtRVmTBZrO+MiTf49VERvMyJ/5ItubJzpfAPJJ3GSKo5emLmldyWGzyS
AJL54fnEL5LSFx5MbRvp7UYZrUb9NIVgFBExiDXSP2dhP/SXSZtbUXDkdug1IHas
wmUPRrz2SETSVoO81+wk2+Wlor5qh/7gH1UZNttid20SCJCMXVaCFTSGUgF9IKR5
GU8y/uH+xZcnyMGnkiRcjtWujLli9yipRMHaH38eGsKZm2qv+yuiA0wV2B74mmZ8
i0kFPQdqjbDtB6uJlKCuyrI80oouutA7ClrIRw2aH5ZsgBQUNmORu4Ogw6ao/4cZ
5E3Y3qRcEOSv+/UyCQxnoLK4c86ydH553hjVV4HJyeUoUHmg5lX5CiR+9UKcDioe
7xLxQKR5+Ke7O8NFD3YdP+E+5xyRQ0GMCH+90XWN7wvDb7ytBbF67vdX3PIEk8a4
jKFxooIEJ5siCBMGFB1YpRWpj97QUa1LzQC6oJOJVCqMaCeZho5g+ZM/iFhy0Kon
sB8DM4XqKduLA/51DCjDL2Ss1Jif6/6NVcRu8nnCfKUlT42VOn1vooHklOCQmXEs
7AcjxIkEBfhoMQ+yPOG8nx3ZpQNb4wiKPrXZ2U7Wd+s0ARSAydXx0qTjswG70nLl
LqIMeHebZ5ph0fUSZtnciFMnN7ffIDiQnGMVUHQfbOJEstmT49iAD15fQJaGZFwk
jNuUA7eIfp645Oyqos7q7I1FXkGdVngYpO4dWLeekt5wNOZcIBnMf9rOZLSFTE5g
v3JDrH3VMgVx9LFJ0VRoPI9v01TcbuX2EvqqKS2OwNnPqR4pXVkg8fuMeQOqRFl7
dELfvS95QfhoPR4mHv/T2uzpTSNf8Y9W+Q1KmLRdRIQ5rHRR9tO5a2j+O5YDotZ+
JDwwUKt0XftDdEEhOOjIV2xwIM3nIVQsYdmhMBcP/TzCY/ggvm6aiZipHADFEW+c
XijnUbvmKCW8VtxZ+dPq0RM6mvdmffrAzQDziSFPyQKJ8DUgSHmNT3YrRBM6R1O+
lOXP5SGoWyta83oAiw7HLJwXVdXnpgUk0tjWOcBx4uySb9PaYNTedDfq+gtm/umR
fsUWJ9ZFDE3/iLThgRdiFrH6ho8gZ79T5eKDle3BcgV+hDrABqLF00L+CbuozBdd
EwINT+J3E2Mitjv2aWPdb4MKsgh91EB/x4Xg/GGLQmTetvMYuGlhY1vQrA5izoaV
pk/FvBxaW5HmE+mIn//IKmw7wxc6Z5EWs6ob2MyW26/cz0y/QK0YN7Rf/k8W9xrk
zdYwxNAmH7dedOsbkcmh4Nh0HY3XOGiL6ck+Qf4cUVwYVsLBiRjsZW59t3RiS7eE
FTbpeO8W4ohceAiWm0VEhLtyyooUUOZYcy1+dE2BAnBSQYI0uXO8l538Y6fpV9qR
l5XPocJEc8l6T4cO9AfCZRlb6gfPQcSxC0I2rhIVgLebFGRSbPV6aNypZdUJA3JY
AMt2IHEaPzCQgz6IEHj708Y+LbKMwhCyVCBGVlwDe1eQZdbo6s94bMOFxA8W3TV0
8iue70OihnU9tQwTFXvEjzn6tSNugeJHKm2SLN8hu6njLnX5VHZ5jDV9cVAvs3/x
2x9nKSEKtLRPvsm3miPOH+rOHhV3NDYn27nIvL01iCPjm62ZdS36nnKD4Uep/NIk
g4KkmwjTdGbY//JJpyGJFx3c1MNQ/QvwcyVGiImXOh/Hs/9qPCFTvBW2rPZS2uyQ
lurwZPQ8FO201ccZPgK4ugCH4QsmaAU/6LomfVPfMIPmJweUO+tl038NYCNm0V8V
cfynDFnRCo0u79wpGcnEpngZeb0NXKsXjGyYUyBDbJBzQkFejvUF5gce2Hpl0riT
RqKUh4Cujg3V+Xl34nn3/mCaUrQJHIwdPnhe1vCx1PAE98OYTwYammFDAfbpjvhL
BWkRjgFeXv5FdOoW2NvoPkhl2iBTaHLwcgow06tWYo/COCBgq7Jbs1fBtV2xGguD
TKRWF/CN/Mne1F1cenUdvipA5V9ise4dDoglQ99Plc5FbueMkzReN0CMAIPJ76UQ
dgFekD3Ppgn4602h7t35CCoxAJiAX+ujRlQMoZ2RnNGuFgW7cIQRaozzLGfdunDC
QDUPJOmCHVMtOGchue4hGqz2H/9sLo+q2BimAeg1DvZ0D2oGstsnJ/Jl0i7T8tiM
XxE2P7TMnj2PP489W00dgrNSXvelXFjQC+MxGw6SbVtALmDAjQIVo+dgn9Kf/cJs
RzdNw05bTiKJMTHS1pGLTbc6k9dedOBQ/ee2BbycmN5FtwSbTwgghaU9Uby2W1i+
0m+dbgJFnBkFyZvxDgwCF/hjLtCxghRRrwJiP01/m7o96UhnQPIj/a6m+sDB6U0x
dRrE+bj+xEpuzLXiBVFLHsgQI1ItyTzVBUsfC+DbzSWyv2nF5YKnUYTleGtCJz0F
Ofd8OQV8RPZqEMny3R7Iui4Z51lmWG9FKgaFaPOy0NDURKQPAQGw6EdN+dkjVABx
0AqdBVKOuB9qNPTcxQjeTYV74tovla+AQee3CIyu2q7y9HNlvpXVXK8RMKB/uuTZ
iA8B01VlgB74DKlhpfB4+JZ5GfNT3C2r3QMCkTGBHDvuTpuT8gaL1Tp+/IemKs6Y
6uOD4yc259obhR44d4rdiuH7OZS9NfFqsKa7DwDi6z89fkvbTq6YqsVpfq7yMAZ9
2aNjNrXsCapObQ/fXJnqNsBuAFmqKNjUHXovDg1Sycs1oX0GN6EL3TRA5Jt+iCS2
RLtBHscyu2zdr9ANkE/MJSeyW1qejw840FifBQW2cBG0hw3xFMsAEpBBqjowOL76
IIjGtkBu5t07nIKZKTQbE3fJChZlvNsSEuk0PhLI6leL0GmWqE/4SJUVhNPH+NbC
fLfuuv0Y2VpeiKZDlYohHJtIYnzxtfLhyGYixdeRwvBJf+7r/+ehSlk0sMy/IDiq
ffMW7gz7dsoKNYRUp7W7JtXFb6z5fZTFljwEwpZJs37KCvNsJq7O83UFLkwT22cp
K6CMnOK4O3lv4dLaR1538niSL4X/3u1nap9D6y1muKoMint0aVIiOAEzq0bERAZD
AXkgiMsd+DWliayQiOPh7FSF7B+RsiqyG6xQViF8rH2/31yRB9zUn4Kybs6eFreT
peoZewrfoGvm07qcWSDFu9cefOEdqsBCGmBbBgsMCm9i6/TSVmx36mHNTRmyEqKC
Yp18jkbNGjpVDb2mqE2KqNNp+8JiIdAC3JZdVaLAz9fRxT+iQdbZ/k5s+zFrhC17
AUO59sB+zlrmdO6lhkssnqWaQo6mqX58fnqEjeKXY1puIjyfwENsxI964Tf732up
FrFsxYUnr14CS13alaIZxK9VvthV1IAuavB50cDHrgEsvOsvoCdS03wCYfaq4MCY
o061MQ06q2MF4/s7uktFzCvVePkupA1nIn/cjeN7acWrXbYFMl6otgMjaZt/U98o
/eg0cs045Yosuu9WJ2iRQnhOAQyC2cCyYwbWxMiCPQ+kT+QQoODjB2iYCq0hbetw
Fto3eSrKj3/uoDXmllIqYTRUQ/lZoBGhtke205BF3fXZ+q5Qa6kc5Qhj8AKaE1pC
ZJ8BHLpkiOo+PAFhf1VO+APeplWaEPl393L6Zth8KfcyARfmQjVgLYbbJ2mf11PV
qIC4VO/WOUKFaeU/Qmoco+9Kc43fARsagmMYnGAvE1nXaBhbzU34li+PpqISintC
x/DYeIztV833EEkng1y+qEaype428I/aOfJIrrx+rUXb5jju97tmpdyK1KTvQiju
Z+ODXh3XHhLWt9mCczr+fZ38URChDqKpyPEoQgonUJiC7I4uf5f6EpvYf1MkxYSc
IuqWDpyE4XdJ89MO2grbtBlNRBGw5e+cBGH4aISqT6HVPkmbwkeXn3HNlG6sH/VS
+uD9PDDqxsDZ6wVCCsvN5OOqf6iKnBfqpp+hGwdidw+EcnH0fa1Ti2BXawot5E7T
sEnA+w+MNHo1kwvC6oHXh2bkf0pvG0rYCOBJTaUcfJPXLjYKl7/8mr97QsfLNlsV
IFeyDeftr9Z8y3eyRJpRiTLqRi91flmTP2X2SBU83BUQO++D58ZjhTjCL+U21NLc
LffK59SbmmnLFyT9fR8C5PooOSCyIAJa5iY6A6pUeZqX2cxLolESnUL/0wG410kK
4RZVWnGEl/u34tM6NXqQ7kuon6n5HzM4fBkHg1+xlujNEETvZ8rHIe03hDlwWcbu
4IHMVVopBdi9ATmba7LGdIIm8hMQ/MjvVbJQIrjstya46IhJZQ5/oVXwNNHH8uPI
eU6KbRnfMGMaIvbHKOE+EwAXNL5Hd68E6M7X15YOI5Ez9CgB5riBikbwc+52Z8XO
ZHKNFnpjCI9VK3/1XrU8Z1UTb9TBX7y68lhukkSDA+/5rAZJoZi9yxw4cXlQtlI4
073UQMfjM8/npJ4MJju/f5ACEKyFXpbFAvbGuASz9j03d0HGHO4w7P99ks1diFxR
vqFSPotsOt59RCQ1ojZ9MJQwTqrORi7a+58i5PDjhTYnmQBylZ2ghBVNxw1QjCDl
67CG8UYOftTnryikuWz3R6dMz83N5ZnpIl5erNtSU+/iMtmPa8Il9mJBBNKclz+/
cSjitX28EN5GLmIRwJX24elsgtpu1XxoPGT1EIeYJRaa5o8drN8LuyLcYViyVdI4
xoSAy3rTSA2VMxrUIIr8EBgB4zrhyXUrNfIuQz7Aq88bfG0b2BTMuDxT08nVagwT
i41/3zz1nSDBU3+DcqAsm6RdKXbFq0un/qnkgdevx7ewA6dx8aKfSx4NrSm397N0
dx1zUMTfiTadCYH3UhKg/UIVLAXc6Dvd/QwwY4ypvEyWwEP4mEHij6ZbNCSU/F6K
T2xT4DU0iSraseqIPa5AoHTzOa8PmYmsPv+EfVoRmlVjgz1XJJelyl1RJs5QPoNJ
+2fEP4oCcrP8ObhFr8TKgaXr8yHgQeJI64eW0DUv5jXF4EWLUsU0hGsf8MjreFmt
2x6WyiJ3QBsRHPh8An1ln6g1rfS0PoOi4IUTTSOtpAtukt8x47EA+v3vRhZS0dP2
q8dx67iTGVNU2zyTQ13/IMHknF0q3Nh+S/0DoGXj30jDjWGnXWe9hVudOiQqjcB3
uG4qu57tSkwHk1SlCVhE/VWg+UCMOK51umfyGKE32N7WJui9YoFJDrdct8a1yvth
jCiAQX2rQm+N0rhxJDxJLOe9BiqRa/vK0sbmwasasEv4O+89gZYu/c5jf/ntEaor
Qy0dduc6Zy7m/U8HSPi4xxQUv/5j96mbFro9/oelk+XcYYsEMFzkHs3wdgl9dDgL
mGG5cC0+10dXkg4gnwELCOjKtSWaDPeRFNrGnosM78kPlMxtPd9+reINVOXJ4l6V
FCQtkQQGzSM75Pgt/6h5gNFKnWYemLJ3l/ff8nGbsTpoJaestCX/OEB4nRTOeZf1
3l4glogb6CbF7XjkYVdoXZ0GGDQrv9O1/s0qCxE08irTKyQb3Xpzm6Dg5jCzLCOg
QrQuWjlqRcm1gtCZ0AGYFzuZQ52fy89FC5lYXdR6zUBK6Pbc6RtmJ87kcxcq8i6d
Hywt6sex8G7Z46zbYtDHx40fBfLLNP6bNPI4IaCgfXfRl3qjjAeCrAIYewbj/074
nyVNsTvyZvqU1iARGdXIH7sJcP5dLaNgpJTcPAMcE05YDcKSf9l6gmiPzjE+ofOF
sRaWCSPHy6ZRB4VGGwYABg0egoKT/yKdceI3M15yWwgM9gWolhrznE8wIs7EexPz
u02okhBwL3npD6HxVFav/vJk+KO3+ngDil4U8vwx5zak5dkd7H5HeIjGMBMK+ZNy
gil2kWERTa42zfRUDsokIBn19y9SsPMIQ96TLtG8ofg3V7VL6QvZg6xatJSJCDai
tebFjEOEZM6WY5MaKmUPXS1mvOreDXkXjqWaZNSf769kSkJ5F/Zb7VQuzEQtSN9E
UcASAxjQBVLUp1/rSOk5WRFEtppsyinrcdr2uAZBXN0DHVdip6NgHTPcKB0ONkK2
WLxlkkwuLQBMynoBVwRHXhzD+9N2JIAy7RPPjVQDB0FgdNwUPTynafcBO/bShUKP
PJmShoUB98leIyR/NNUnQ0gR6Z5LHpoBOQTMWCzbj+Q+iNKAV/uBfuGNaNrzC8nO
zkl23UluSQ0wyjVEH4KwV8rXP+n45a1KiZarYpRRQPff4MVJRc0FDoYELSrGBeHT
2x3VLmGY3+L79Mfu47ohJCopRCGoY8WGDzpyArbjc5jzV6DJ2oV4jvYstmJdhksa
7u9ZGQOo2nsFJaucSrPBwNLEDohP/VLgKMgQUQutyNrHQDam/OynQOMto0g8mA80
7EnpOSedb0bVRGazczytlH82+9hRb+97kSsGBY8KWgohHgOUKns3/FBUd9MnvUYn
BezNd7uM409cGziQRVmerz46mQN99uz6W7Pnz0vO1nAXH787qYrto8Br44VaM81g
nadLcybhNZom9gDkaDMG44FkM+KCcL4LvdVI4/u7j3mmveUjwWE2lWlRx7U87x9/
J89FUQoTuTg21dfrMJhQm8eLXzm7kbZPhaMnpwu1U++q0MANFTyvBDC80cDBidIt
d0vJakII4DiWpwXV0VwP5wYMxlFtNo3uSEEwJtRvFxTg7PyGHkrEsNomgOZ+Wxp/
jFeLTglYpYJyU/3kyxE+eFzV78Ay3sCVpMR6j038nNJwhyGoo0iUh9zGaELu9kd3
f/lU7kEQVWUwgQTqf3HkPcuYmF4vnDcwn6AgLHOX4NLZ6vArNAGZ38mGOlqY4Lj0
WzGvSkBAPb85r1YvNdBvYPGXrITa4Vpu7wvy0sdGfK3Qdz3NXNXYsJmI8PPokCIp
oyoGV5pR1BClzuZP0NVTcy3Epb0WBohdlI01EtcCQ+iZKhbyKFqcWytBWjkjqeG3
D2dqINbIkiZZIvmSWMjoqOk5qnA2T+jx5JnJTZgz7D1F6LLx6bdHozer3FFr+Rym
EJmiFxROg1MpvCjsYbPRk2BNwA8IfnjGePRlnUsNCn2UTwWvnkQV8hp+vHqDRhpX
GtFv96Yvd232RJzW4jBNWjn/1HSKeMfodObvKgi1X2Vwt4ZVC6U/Iv3DXO8AJKCw
pgikxWjM4vzPA71jYyX/HJKPJ6HwzPJ5qDoy0UxK3jqEwCrfWG88UN9vqyluYozQ
rL0TJBBnHD6mBh4CgSIJ6noA6sgaFqwMAihn06PtfVFIVy4j9eO51ssGOmz0ZUN8
b377bmYSYGBCJJpk9IMPly25YIKp7iasfDYSAOkOGbT/qr4LUQcY0CN4mUNqX42R
HSFrBQiPe9GEq8/lQZr7Ze4rEOlFgf7FOSOaVchlCB0LW/5U5XsBzbQJgyhsZT5y
FbrcjlrukC0JPhYuARf//xH5hRxfTXDmzr/20tokaCT8eh2ZFMe030oKCgnLdqEs
X67zUiF9IBqj6ZFanRiawkGAkhbv7Rt/vYMUE2paMp+hGUhIwhftJXTg7wJWko0w
8TlUl5BbV2RdBPZUIS3aSgzOvoagXsyUhHSc4M2CxvOCJr6OyRL9uH0uVxePs34u
gg2uwuV7qMWXwU2Cz/+CqfooLB87SPu1UYv/Kzs7vsgcaf3eWyX5JPNNdwRMVZx4
2xYITHiB4KUidzCIbDRe0oBLrIbknC0u78+eHiyibkXj+9LaYSsaJgTZes/m6eL5
qIn4VgQaHRPW0/t/5Iea2hC2FmFFMMbOb23rPq67kFonOT72iAIF2ssJ8U1tnRwm
Ryf1KDCVV/36s1hvvMp4UPJRVG7gbKnYqOYWmCe1sLSi+Uxh2XzT75OhlGDu/N/Y
5DbF3SPVEtNcfKmQBUZoG2swbJgOG57ynqqc+leQncdxMDi7DW2/778LWWq/9xir
rv8GnHl5xWb01tvwbqGmWJ+pVXxUNVkw9XVQx8ltfS/YxJ0hJDSkeGTUPbPL4DTK
2e7ltgUov1ioMbIMu9Ish+s6TjcOI8kG98GHQ4TGs+W50AXlrtRyirMjsRsWgNoA
jMgkdlGxE0/4VIPf1+5LzWj90OUAPjrZkYSIbrLH1RlmJe8y0I4ZMhYl/zy/O2MI
h/ejlshbL6csH676faiJBvCj9hOK6g8Yqf8Okp1b5Gy5EYh24DacRk4zK0/p/LQJ
ISav1nMYoDNShA3w98uQbSSXxkoJ2pqGngTqtd3I6MUugM8+Kg0ev7Le/AHIWERF
xjFyuO7JYY/gZn+G6C3NXHwnOcN9Gdmql7VYO5ZSTRi0gO2evIlAwHp/9VQ82vux
zk4OVuy7MthMY7kuwaILhrYiB2dbl5SVtCDQzx3HMUW3gRtQuegc1LibG8vTyOoC
ECqUm2kDAYks6BKi0PZKAkKvw5Qc3AJVKehtuKk0FE/9XPUAFsp8Pyrdwnx/Okke
CoeA6BL+8X9a73O5ax/VklJI6ss3A4b/tDg+lPBZHu4dD7SbvzWNYGyeQEZHCxnm
v3knqJ0M+CheXlPIjVO74tfv/cpzaelkbheh6zfmE/P7bERRIKOA5JRlFn81TQHE
lg+6ewwu3Zrrfo7S9hKlZSB2ml62Gwxc5g2OCX3yGUsQjpYLp0qH3QXBksefJw6v
pbkOzf5SAPAlwfafCfLtegsgDQrnwLLyamKR27DHTvuQcybBsp8IspSbH39cgjv0
BDmV/n8YmyvAGg81aYg0UhcAEMpRq/rnFnuUCEJpy7uADX8873f/dVOH1YxH9C8N
Spbl2IMknm39EOrt/pKmceGkJcRHNqIXmRyyZ6QYKy9jdHK2mLWJY6ZiqOANa2qj
K6X+t4KZLBuGp9xhAa0XwBhkLQ3q1P/MuQMCtamD/+sQ/Pfi+LIt5foPl8myn9RK
`protect END_PROTECTED