-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bOSFOl9ZJsKWeJ8d2h0FW1wfs/wt4EGzhmoO8lni67DwEnaDXMlDoo09gvAgxV0L8945KWiMIr5z
tJbUL95fbJuI0NHjv51/toFNDdPKDS4qjUWNyg/8D+5JHtK1CG8jUSx81Z/fmQ6psmCBYar18/9Z
NgD8Je3yN1cRzsoAGFE0f/9iXQeW5mgO32smDSO6v9P/gBJkpoURh/mxWzhVbcFEjWmtGujUIkfV
IhRJQcWCD1Qv195OgLBcT0NQKQqo7VUd9+SbhEKZkm+klLfY8Dm9QnasMvVLc3iv8Ew2Ud2WF/UN
tmMVPJsVczBMm+IiuJh3KhMuuXfifbkvRKXAhA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 88416)
`protect data_block
+KqtbMjF6kxrmg9YfNwnLCGphsKDhXXQB0BeegKbERdw46bZ1PoqUU0Jp+QbM9ulO0webdEuuzfZ
aLbQfet9wrK2rOQyjGfe5IkfSSspjSl++V9EhFd2+HEnYvQQyJgnq/up3DOssWn3KoAdxFyO7EJ9
q9SaFFrsGguna3ZDWI0jqDLbEOU7A+C/vIvOvgxBU8bvRDu5lVkT8TpxXP3uiMIr2u09tAge/Z/w
gTDbYQ9lWnUcowN/FcKQ5z2V5t2s3fMs2IOhLvkPQAavcUaTA9K04A6Bsy2n8ocuDVmt9/LuFQN2
+gVfaXh+i59Li+la2i9QvccZCFGgsJzgX5GYq/KYSsJKpoJWY5tfj7hKAZkn1/P8+2ctIX7EofBi
dAF372E6sqkqcmTXceD2WRLIW7ga5WlWeXop38R88j8GN7j34Wfx45I8jbiVvbqKIq8e7yLPAxir
v3kt/D1a6aqGXdFzEyUGhy8qCXzx4bZUeVIPaBdPTQbcgBOZWWo+l+Lf7gKkyHBV4iFiz/yPBGXa
t75jCsUgVgTCOtnwutNV8nE0634le8TixoS0Kx7N57N/gGnn9+MPD/NCaQZc+f6YWmQSS2gHOg4a
0/oAWZQa4fzIHLoNVexukuQyT3BHpirNKvsCFKXId4yvNI6hZaY2rhlwY3ggbEDdpEzB/5nzvm9+
YK5p4YE4rpDMjG1FO/wat43lStx8NaOU5J6k45uXLmMzM7XBhMaek8PVMfJtDc9+E/lg4RJxlFge
AN9swRXoouIAfX1N/jyDu1CKm7AxGM4mdkQvXmxwUuZntj6Dq3rjI2GaC7FOOc5TTHcE8qNku9Z2
txdNHoG2bnaHPO3GK1gNf8p7UfYTrJuZ3lZc7/7Pw9XD8WiHEPKxRyuFDN+w0Pk3illYvtOeCPJD
BQV3yLdqcSBjKpxDbMDJi9M6R7X+1nnt77JPr/DOSVVX8p+77KoW9zIoP+Bkbkhk29tVEoETBpLJ
2x2WLsQyhU2wDFGv9FtJ0IJhQrxFaX4kMrlrg+iUOnDrA3CeFWCIMfugTVFO9brsJeCNAlOIKTH2
fojpZnKWpLhU7X/1APQWDr6J4qIBtutF9uHa+qBc+LXNKrHIsQpE/jSzpnaHwFrSe/wdVfFH9+m4
ExXYypJjzyEN902MhqgOGtpdy4Yeilq2yfXrGAd+E46Q7zoXmEoanm/H13Vtrk28ZHJM9pAsQTHj
5u3gkk30jnkFSqhhZcqRci+j21w6vqtKH6e7wAucfEAMIhtuhS4MkI7JtQgwAjGQHi8AMHHBQ7hW
FrfJwC8/8gc3v/byCYxWfbhg/S/1AF2ki/L3+9xWRSvXQUu/canAK/BTKs+FoAro3jS1wJ/fM84U
/wE3zmBx7aR7yR0QFCKNSiM/g3n19pZrH4UTHVLA3/VKDv1PXvlz/jdWXlOP7UrPowmWipvp8XIT
w5q9bsm0/qu3name3WPY7WkkLSFc+X/JeTir/nWYx/WNz/MhhP2jQStEcVj+9Ldh/tHPYFdpnFp+
NoekQs0gM33aUleMpt3nq3oVuPGmwRS130K0Yu12+zTSzQfRxAlMOqqXIEsYHML8deqkTM5ve9R2
Xaai8Y6F1OW4/yIUhtb4GEqdboWsMW4osMrQBrh/CVg9SoWqch2XNmr4iNoF0ljfx5cd74XYoJkR
5gg0TCySqtiFUZJDoYHigm51JrZgrGfAmRn6He9UAg7aL0U+zMgvXcZPKbwLCQnqxEonSa1jRIvR
q8zoLaThhnIkafsVLaZjwaHR6M9cHiT2Z6FrDtzjeJT3UonFxC40W+MFEDq/lVXOL399PFy5S+ZP
LSVM696Iw9KXAyt6+So6cw2QbKMdhkOGmNyJr9G6gYpP0+jwW6phwMq0gRStg6EML4Eu+QWZZLBa
KdOKNVu7Dzrs0UBX0VPb20ByjOpSSyCzBojjtiWkxw4Xy3f724QSLxXtDQJF5AK+mt69NsS76XCi
++BZso4Z2i5MfBXSVukI0u9TzaxFNUxPMPzF2wAKPLbmrGMhNuoFKoD1B/vPtyTqHg4Om98wCiks
VDYCcIWDtU/a5movXL4coneKl9ZAjgWF+ZLqbyisy6RxgTOBwmtSFVTDXSmVFUD3CMAjjhNPsH+O
/8kXRsl9BL8d9Z8s7MaDwxb6baaRz/Wzki7gfme0E4Ft5J0Y7sb5f5jCkHReK2AaGqldbinEVHCL
neWxgoh2X3N2i3r0CT82Ki3vJ7L3DXm50bGHdrxBVOLcsSjr+1CZUZkhbRGb4iaS0tWR1dVQ0KoR
mzNLlqJmBRZEjYCXZTTywnAmaK82KD40o52tU2gye8iWiXMq9R04F2X1k9vo+Fmq9rsAVLTfN+Vn
mCV5d6q0qdfO+5K8JzZjNaNHVEeYi/hjMhPW9Wd8vAEn0iJQqRs1y48tcn+XV807sjiVVfh2pnFw
RfoHIW3aaFNXMQajJGyJVtjIktWDvXe+MQCcZAqAGHoUppgh6zA3ZDwtB5MjffZe+MOLbxdOptkx
dyTDlKtr+mjSntct22GfmcQ5y3TF1OArSfeXxmZufaf7qNYz8QD5ue8oT66eCvLj3DK6Zc2XipGm
er4pWA6ItsJV2kCB4iklwjExYEPWGH++7IJenmZAAQv14IUjod98xDEOlrd62FBitg1QRagcfLiA
IxHZRpye6hn8xiGc/DoAFFtFi8GefT0kbi28o6MXzkilF1BWM+ccSqx4CtH5fhtuSDcJf0fohPK+
3z7U9MlfHHU3wweJpFMz6ileNfC5IEZjdrnAcuj5MBsbBqXiq9kew+T6owclpmF11h8A4kHFo1cr
TnUHbDMopJnq/6H4LT9OZC2by+LLHB08UbEj19sRHAbmA/eOuQXi6OMEKLZ3nVvE09uWzyJA5UCp
2R62un+e2iRFLDQwF/GN4mCGaeHEBe7ic8yJ+ulB7sxNy/TQnQD2jwhLnOl3l8xSBqsJ7g108Z7n
TjmEGejd1tTqMHEktzfkNyUc06WSSxvLl22yOtHXhCp+fjWEs+6ZSfmBUTys9BPbcK4ksgPv1Hbq
3RtZvcyNpWobIUsKALnVfqlLkrCQAlrIGpFsag6Ihcx0DwJxs2kt7YDxZ1g0yxtkr39R4Li4MdGX
otFXuKYeescPWXfYSxIM+gQyX1Bbu/CTnvHFXJl0o0QmF0DK9+zUUr3qMUWKQuQ1nNJoHbTeAkVD
UlJYl2LSeRqadvTvwiZejQGxAVZ0Ko6AHciHcHICqgVfrL5t45WB1B7oefNXPPfT+nw/myP7EF3+
CmxUBhK2urS3ysBz1y8Q8LJx5+jQmGokheo5e6opnZueM+YwkhBBlhVPXYJ/vwCErMqOcbcaACdT
jDFx7u8xdDoKH6nMvJymiHf0UgEpn8x5cZmUwdognKcBYRqPYiNRRYq4hNkW3uWQL0Iq/y+wP32r
HkiZqTy6h+43037V0HmK92Tc+Z4ETu9fte4HAgqf1zmplaFrJX9EBajwldIjreIKKXZVfxasxzt3
g1h+2BWthUGkSfzPE6QA/qBlBIDhZZdIyV8HgcRtJA0UevVSU0m2xC549xuBXoF2oHr+mBfWRtXx
zn4oghgW3halUI+++VJdQFOU7AZ9x8l4W7imu8TwXpSCBvet1wT64pldr+gvSc7Xl0dIhX4M73ka
RJ5zCdU+al8rnRnUQIoTuGqykSnFISL0NDGcam9N8tBkEHdx0UTRIyp2Nhkvvlir/KQj8PItF5Zd
HSRn/+GnXECvzac9D+HCHcsuLe0JMsqMmj1od/YwTwkOhse9MAs+zlsnrWu7XHdbgXqyQFUr7aLw
QyUAwA8xqctosYo3kXccdOArzj3tYW7zAHhcwx8Ct9aucfE+PbgNKvOLEQOyzm4YnE/5NZsBoF1i
e9fXBCcmDkS/xUVftPY5XDXUNyuBm9KTIb4aM/THClqaPmt3c+0en5q82y3Qbi1OCwaso3qx/P21
qKuZDtohCj+Y+8A2z4Iotvb3z4BhOzJ6fYDllj8ZO+mJj1H64ssAi6OPfK4OjW5//rakdN+je9u/
DRA/mPsn24QG5ZP1pUY3i4RZk0+MmqCGNstvV/G0/YBDR9r3yRrlMTSBEg8IDduhaBaSa+fh/+fT
BvmgtUksVCIGMDUgg0EW6gZvrVDUV4IGpZLdGV8tXxG80jDid+B3ERnrUMxsd8TIJf2+gB3rH2oc
6aLA++WqIg6ur/XzYvFxh4ucXIYhOtbWtD/nDhU99eiCKsaAzT7V0m76qUoRawJimBdHVPslbJrX
egm3hb6UcBv6jRQSzkJ95Ydd2K3dKiMbGtdnKc4073wdi9fJeYgXKt7IPchDljbekjalyJRWeWZL
MBLMNGHedxD2wg08b65qt3LsMtFNr7cYKrn2/j4skTqVP3SiY8EH1c3iXkPXZLw5Mhjf1IfXvf0U
22WnB5DD8azfqQiN9vsAkRfhDBAKHS6H9Df3Al4KugYgH87knirLUwsHPAISXIdG9fGuwR3J6HHc
kH+ZAB44L7FZ7/fAMqAilUsIsieXyanRS3RtkcvrfQBTbbakH9ubYKerubU5Y0b46ON9UGgTQQ6d
qAB8Sucy/u86R/ZO2fb29eRb6xRxSi8kkLjgr9gyTbw1a8KOt6gWnb1SS0ye+HvHYA0I2NnzetcS
c/t70RghMz9YfWrWanFRq1wvT6I+FVwW7yR/MU7ffZ7Kbhjrki9eajyW8YL38E9KDnRae4A8smcD
CAYGKeVKdM13xyLjBskS9+XagmvNMJH/4v2Aw+2Rlg90AYO90X/xpfjg6BPU1XpsGDvzhI5lUVwC
CUZDCa/7KToTkQRFCjkfogtsVz4Lk0cuvEe5cgXK6j/S2hIGsrOpiUvUOtpKwN65Y3BuTYKr8BiN
38bhTBWExXtmvHbVFr7xQ8TYvchexWZHOwQ26+3HvnKb0tTks3JJdT4IZlzYaBQYNbgWxslzfdPV
A88El+khhkysP4FvKsS7HJOc0r3vg8eZm0af4TuWAwvN9Wx40E27WeAqqdbEEXp5gFzYhQFG2vXP
Sw51gng2r8fLzxsQWD6btOV4wyS4PnuB8yg7A/Ae6PVTiI5cssLeBKS/eSg+MmORn62KzQM0BffD
acBy5nIA+2qbauObSPnx/rVuYO0Yl6zQCzxMuLnCt3qh6DTNmv4tnteJCAaw7k99WpU4Z+PRrDbv
UuBhdnEq0gUKnRz46x4oAKQHORQ1ZPH7IM4AUAHtck+Z5eWNWZ/z5HDoXm2j2RvuilWCNQaluiGG
JCub261aUyGvx8M/HU+6jwWGkLq9DrTrTNvgHw/SO0gwgTYCruMUv16jAY0VrgTmmvtUqRO7NeuK
/0XJZAdGLtzieVA0kPMoRXJUOtB1J/UnTknbH1iZ4gDPVLzI4H/LVnY4u6WfYXYHYl+ycwz4fP9g
U1fHTfKux2xx/PWhD+JquymyfHolxcAFjNLKsJXI4JIxqNRcwhNjedVPMw+TW0xq5Ahx6VvvySEt
cOhhXAoqBJOtXOUs82TgWDuSk2j1fvjrqlqALLD4yYaUNGNBs7KbXZz8Sw/RRqKFHlJmPuHR+pUs
OcH9mgmW9w8iGLUAzaIGo+gmrkCfq4vYraZ3IouzFAUjj20+CPqH/62rkJk1e3MZfRwpQGyYiyEp
E6ydPD7YDLBq/UOkj4bRZsBizAQFYo4KaAPtryw593wkFiwm8layoW3cH7vzK+yIdhwRIv+j103L
uTJQfLBrSoMRtw4zV2q5D4Elp/362DRIYe11GQNGReE91jAhtxcXYS3jqh26kO0Po4WwjctRm41I
spp8rZZE0XZy0IOIBSRW/4M05f6/ofiwVY69tkO7f4We1UVMWzkgBfoeyuwZ3vMNhW5BA31fm8B0
U1shhEyp/WlKVUu2OWS9FghZrI/p72UQszqghxmgeDdO+gz3VUzmOLJZLN77K70NWU9necHKB2mZ
GQscjguv2wbarmYshk9B2N6cBbBvtGAg8v5B1pkM1Ia3ZetqtXCGGoJIIXtJXWQBet5eLBVSIHzW
5B6CuFCudi83ANP/ITB3SlwhYojW01x2oaGmqPkJD6jWOUhl7YO7gzbGD2vuq94/OcmlqWpY5zp7
F582lBpJbxgEx4GTC20pA/XWw3fII/yhrnVZQePrOsh8DvMu8BYEPbbkcVvC6uUxEM63/6cLFuX0
J4E/LJHMepWUHsN3XJvws79OnB8aax8ZuXYs8GtfGWG2wQOmFm1Ypu0qZYr07EjKhVTXHOD4rS0Z
s91GUJ938P/YMgSwfQ2K1Vsl8m0RAHG+UoHoIth7i9V1EeczuSKr0/QKeIU8edchhdYxD6fOVA0F
4zwRkbgTGDPSpKsXVYkCEdyeofZTnTTrbO/GJv6S3ASX41aKjUIw5Hox4dHZ9DiFQ5ZRMBlN+nPe
G6tVSz7wQicuZN646VfDcsAt4MJBtbPiVYMf2gir9pTGJK44+GZ5qqV9bbc1BHIVIcXizH7pU/ML
lBr4hg4k3CBt6Ku9DO+mdH8U9qnyvse8JJ8K1FrAOEZlQfPcZYQ0ULjfeQuWOgu//3zk6KnWEyux
nGQZeMVo9tUFAKGZ0jzOTDC5PZhm3qOt+S6VpqGNpZiIo6i9kR5BiHjkUwGGpNOnwrczqZ5DAuHJ
2WXAA05qgrgRVZiRPnj3/uTxb8238kketf1wmvXANr5AJvy+WpHpbDdjBpfiDrD5TVdh/QZOdpwc
aNjJudBkxKp8zZ3vVCGd0EB41E0zKAYxCwNgmst2zVBq12QaqpIlvtrAFvZmm2R4ersWduIfo7D2
f+DtGBz8AR6Y88Jp/caT/wsUrjQGi+ULQ744gC9o7HcmvxFRuUpiprvRvIT2rmWcnX0E4aQWraCP
YL09J0LrO4vbzBASvKNF+dSHgwQsF73TBo8aPEhXUBIlnuw7re1EAp05oYeb0asbw7TGkY8dtdX/
x8kjMrqq1SUHp9+h1E58JUAUI7obGnNrPA7CFqRejT3SUMx8o8LUMmEUW2M59S4QsnPqaqRZAfXO
G/Oh+fl7KbyIVS27856hKPlB0jDaL4NNCw2V156DmbQeWPRewcny2cyi1tGB4PZMUo5oakUJQ9vF
8fQSSNjX5dgUhNy/K17mK6K44xLm+09BnejVw52GNRYC1MlVNyXchPSKo79WzCGKy8a41VP7xrmC
+Jy1sJnSKqD0jXcI8VeJAlMEzy8qWtjRf6zImHEuYf6r0f0uLycBkSLwNbkrf4XkHiQWcI9IoaN5
pPiRqdZkJaUjrAdnlatJggpyiJ5+P8YV4O0LQCGcF9u0ev0fIFlazDKDy8Y4hcQZEEDBk+RRbPi2
Cv8xUXp6ZSZcnyHgW6dERtqAZIuBzru2Thw1LDP4B49V1RaXsuFitfqu5fpr91EsQ1ba0Z89dSxb
COhOBodZ9wIk2ELudd+F6dE/JNnqUz2+kPf0bZc50jlmmvfOS4suCxfqpirtfbqXm0oVEUIgO+rh
ECnUB+xE2YgENIJ2Ey44zJ5PbgdAZ5nmqiljoqiSouOvgE3aIu0pnEnjw7J5yRl966Av08ofuBus
BQHoWMKIblJUR581rsN3R4BYrQ7QaO3u7uA66O19ttoTDrqRnd0rQvNSpYkvO9HiWSRWOK7YmBZO
9MFJEGoOYju3F9rI8Nlw9p14rpKsb1jzsucywVL0gXsJdO7h3LTCk5/DoxnZa4rJP7HKr1DSPumZ
QC8rI/zYFiDqb0TK5cX5c3anmelKT089DrQmoaeCl+tMVr7Vd2kmNsifQGbGkWvI62Gy9p5PXyzn
q3EUKKeuuYJRSRGTbkEFY9fQFUK8akVyg+dkGA2wMv3fQPNzPoRK/ll+S5qffV2dTkXH4dHS/XFQ
JG8PRqMU+fprKFfVEgtKclx22bYkUAXgLR4OuJt9K3vpBHGo71VRNwufNq1KpPnf1v1n9Yno9LwV
Tv6nUBXXAFQCFuToBI54qyPbhy17FtdqmSH6cOU1hyHFwKEp47N6tqxns8dhDghZ5e8U3s7ALClh
iXoAMszKxlnujV1rEP5ax7mQkD2IDnK3hGCt7zFHtLizF6hXbMoMxpelcJ+ADJ2c55EVK1oJ9U/d
0/QlYLF/yt3UvAvnF5L2ZG4D8SLih8mv5lkhEoSkK2EImy05CbbgW/tyaCKP4ibksE6QsWvhWtXy
ItuYyJyC2tgB+HoOyCIgGl+iPIqz5I2HiDXGazTuOLi5/1xB2VWsbXdLIEpN88QjV26BS5h+JZ5s
HYyz66hp1hr/EDawYzwqUVQLIhqI39ziJ3Eu2WYiL2wxCvCya5bVbxjKI3FMzVZBTPozGOuPmlyw
tt/flFf17E9whym7wMEz+NRD5OkYwd0kOZhMkTmtiyiOHk3roGX3oqOLc66r5vA/uWQRqmk2F6Uv
Gs0tgOjxZyqTFgfGSZZkPEuPVeDO6zAp4LeHCRjF4LqAFNLBxmIE9BO6rasBth1FnE7lcAacQ9Ii
uVikUNIcS+4KMEp98TLOwgPu4P9O+gwghHwAgUWwoQ+88RpGWicH9VfwXnGHMJ1MuI8c/hHvbAz7
Gh7qLzD1T9srCH1Z7KfdSjkv8ysJzNJDMKo1NILouDGSbPDWpkWlF1WBKhVXch6JppElQAQH1s6e
pk6ndt0lhuk6qECGxfzImO4pyiSLge8pnG2VDQAsLTDbfFoUJTS1/CkwwtTGoRjtLYPpm8x0FurH
tEENeyhZBfL0O6pQrlE+TKRdgYbXt4l26G+no/uKo0JgY4lO8fpOvLokpTHVQVsS2J345Fu6F9id
UzFUhbTb7DSneVHFcDV4maaiBQK/vgadhTP4KrfF398T8lkGecbnkFaKQECH2Mt1NJGSW62gtjpB
oTBrXklHHRvO4DE/6djfJdvpjyKlnT1krjjdZ7vzrzNk9mFgw25rOtYVt+qT9zXh4jVtNy9NdCGk
f0zEX091SLbpAxorx9l1aZI777HnRjVUtXAF9LqOYj1wKQL8sbEqGBqXWeicqiRJky7b3F6cZKT3
Q6ZHpTgXIOCwveJnv/JfcY1qOjrpWo33bDtkDnUobzQUv9xPuEmeAz4cjl7dHlRD7S9PAWwZ/LPj
7jJkI3rfgNClwr9umhOkRM14IukQCJRXKRNB27ZFYGLYxwKSaX1kc4IzTgn36Ojc3rheLfuVj9SL
n/cv7q8SQSZ8O3nOuY0Q1JoTver3pmYu9fPQElE+1ssLdMESMqwoKuLxT1TZ5dwU+KaN4CMtftf7
VVL35GuslYtePxALOlrUc4FYuM9SCMeusp9w9qenmuHyJPatlB5wJXm19amcG7bVudJabhigA/3G
4NK/JJmD7Fz635jLx1cz/W1M+O49XR7rcMMucZ6RUQaqR2HSmXBcvFywpCGfvKXi9XxxuMoifR/j
+4IIPUUgk8A1a0xXLxoBgKsQ+WbBcaCkTwU/XUW9rwa1rBQZ4JDtK9ZOK8rgIWK2hAR2U7qyUDoI
jG9Q+CbSDyL05ZAxyurTX5gV/+uib/dncG22SijqFlf+N5eBQFuX87fYTyD1/bwH+QGT8QmhjcOq
pvlEMx4/2Y5Hz+CeGrs+9jx5TPBK6evedmjTQgX6YeyW8SpYano6NQRJBzUwAZ/xDiMYafxxiqlR
jGu5CXfc+yyElzChzy+yGWpdwtf4G85RNwIvt3Ab/BdcUH2P68CW8zDcVbdbItl4UqtAB1+MZBNq
XXUjeEVK1TFRxJkJwVZf2wROYkZPaqdUdn3df8KbmUfoaOMxiT/wjMI20yEVWjoian4rjmJ5l6bI
NEF7dmA3/qPFUqFh2AGjiF0l1ftPRKbkD4of5bU4H12/B1R78C4wv5eHG/F+2vveO6TFtgJSHoLL
YCzxPRQuy2IJMajwUa1qS3xXoqDJ9sjMxavwZJfYJ1ysQAxnY9mABR226QqmqIlJe9Fwe072FdiR
/lzyj6Fks/zVibfwXPCNeJt9xoRF5hjeR+PNBb/7cZJDDc8GKZ7bnUIQcnOUt5IWBG/kduLNI4Nr
bFBocXi+RPhuawS1a0jbh8rCVVEYYvgXE7SnWe6nOpheni135bOhw3a1bwKWspCaJh/U+h1E3a0m
XmZ0SDHnturg9an5yFw3ArOVdGNpqWR7gKA+OZJlNXePHGwWU9jxtW4GX2SMLg00dKcLWoBTpZ8V
oqPtxH+WpweQQeOPGgqjI23iFv3h0wlKiMhMdGTN/KEbDYl9VM6tkT0i+NW4SkgrPl/HoPxfwvUm
QLm1qYAuKVZTDnvMbVEuQ33vjgWa/VnQ7zZxGReaUoXRQcBwkPmluqJyp9d/S2LQsGQSYFomBx5j
Nxd0xyj9OM6DGT/0lOT4IBOiO2ERCEpIClumtdbbEW+ViLG/OCLdSEYZp5fdKnBqEsJjs4lmvTC0
WkbjOE34UwB7T7VCGoefQbD4LLwRXaEVZZKopo3vv5r+AC7ScwxUBrvrJWF6RKRxtsZNzq7qKR6O
bSBHFrFqzLlOqirwQlBKnoFK+2DWM+zdk5DsSuYfk7Yww3FlakNg6u3nOPHhrpuJyGUcSwgdEW6Y
M7Yj5D5V9NJnFA1dtuBbQMoNppIIINmgN7wA2elAfpD5eHxJFdS5/x3WqbDjaj3v9ayazgGWoXti
1ug4Q1avyhGZ+SlYIr89LrH+3F72qs048ApsET53zthB5FdjEny+jEUm80/0wdhcKmk/TYDX4Mh7
uR5MEmXxJo6sqN67y573WpHCzCwWcaZ5F+c1kC4XNwmdge22MVd42G9IE2q8yKPwLU11/ejyrCdK
Lq4Q+esf9Onh3vKAz3zBS8qYv4ZLTgpiUojK4sjRjsYCekM9A02y/lPKKic53ZDA6Gk/z/Sg22U5
SoGj0t1qB3cnHbO9lVxwU+GPajzDmgliKiVy7dpKauew+PiTnos80ihCKoF3WfQBAZ674i/9V7Sh
ppCjVG6aTMjWVwBdT5mxjU4usMEiUEXAUV1JITCCw4f5TdbbAfWwpWGnwfWdSaAlhfgsOG/fGO9O
X4Jq5WdcPeQqvY8cQjg0Vos7Bo6BEBM56aOn6VZoJnXfI3XWMjanKfjGOAhFjIoK8eEEaCp/6PhL
cVf9S2saawPVmFbwFJFD/K2XqR5iudkFzRrcn5rfUP8GacSHBoaU21KsTkY7tkckAQktqoInFMz6
v/fALAcXg6cERKImOa5M7da7fy5lpajbVHhSXIikmmpGwRB1/7W+ubxy2XaKQ4h1/dlXBeAGvJgl
V6YRZsKtWxm/LVqziJGeen0HE8zqZOb+Tcn3utFwpNL+bsmycSVE4jf02nyXm94maz8QWh2v6reV
YFLn9LGheVo4zEEFdgoF4ZbK94Y2DLYcslTkS6FyQvTORu7Hrk8wL6BJXpzb6WTxR8p05CepMc+V
EmRtKwgEUu5NyOFf/Rl9QAEgd5oy8hGU/f8dNBp9v9g53B0bCqM4yIvsl/aMQN4XRd8x5aeYTVRF
f+0L77yQBo/HUWpbqj3uz2A1kXwIe8Mjz24Itiukh44Gjd+snIHMi+2kJMVy9bg0WDz7zlybLFLg
/7xpGhZfo5PMHPaCmImDmdZ46G4xTEZFwxhsHs7TPX3XrKoQ8KnIlx4h/eBRkQHRvK1ZbZx43QQ5
VTOatLMAGW3c6NWquXGy3GUoinaqoroGK4CskTA2eyIlV23GgX9z89VWBn9Xvbnb6n0KceQhH4HJ
OcyDi7U89Vg5hvQ+PL36NjbPtRuaLhvPwDjYsrIQjpjzqxFCsvC1IxnTTlI2/aMF00T26OGPGzGs
GMwzFZ0RphT46GhShmXW0bkbCCKqz7WmOBrdaXJWI0fd8S+eptL097tMFKRSjeGVgASHMNsmsqE3
cXXeuYSwoU2z2YQYYzIXPchRfj5DvBv3o1lnTU8ZfNZMJi/EbL0Mex0D6tOjZP+q967+era7y+Y9
ZSbbE5m3CbbzkGKLx1eYwPRXbKFaLjdDM/4n0dBAyOyIv1GH4GsIzq8dv3uc+1irf9CRYKUgdFNv
ag1qE6QQx9Hes/gHdWuuLsmV9ktCOVrGyjnm8Ti6dDKV6ngVpAWV3X1PZV7Zx+/UNcYyvPobWdnK
+j6PEADc2oKxptB6pa4OcF3YQHtjKw5oGZq9J1okHLQ+461nsrcLMZc6UfA5SFwaBw3vm2O4qV/v
mCYcyiW1QUKkJO5gs4pezjeUQKBs3kL4YhI1FRpqCvCIsFbkEtz6tNfByLsqvdCS/yI7oPUPEn1R
T6elyrFMfHaWist9sMQXccznw8BukTwfBoOtBoGczTZ3gd+rNVrTDyYSKJIuPtUrMEVxGTrqyVSn
Ke+Xyd+1SQpefW4GNFf8EsMvuZM7OahDcPn9M1dSCgG/HYINP6yN4ohd2pSjLrcfSi4o0trv+CXC
MgO3vhuNUnUQVXWqt8fWYFMYn1yAZzptfnAGnYocA90QZFub3MnKiV/qEVgHBzVvjRIdKcLcOYVS
CoyKqvEsDUji+jrHOLXLPLBmKsCKTiuP30KBkwbQm36/v4nomFn04jpAStqV83YqJuCVf8ChgC5g
9B/E7GAxZ2MWvmjL0Stntks4u0aK75u38RjWD9WyFiFQ1kQ26CdIy0/Soa+tMQCqYQeFOw2Xmju8
jm5jG4dL+wjaOfgf3eina8nUVLtcTd9Ai9YrSaH1XHGCreURNmkmAhwa78UE5oaOX5yDpVsEYmfo
9JOLQDgMKo9mo5CgQbnuu6qR80dOQ4++TA1O/SsFE+XmKM7zoU0Afz4d1TbQdgQ5VEW/x5l6vHL1
himFi3DLBnFtJtOsyrAx+rnED+GUFydxQMyXVZ1m4CKCwU+/6wzGhSZfAdn/lBSTUijRTlSAFQEm
8EMgN8vWVdSNWULJNrR1+6gduMla7zxs02Ez+YPutIpgTYuV/6uGUlb7/u/gZPFFg7SovauMpDkG
un+oAeJ8eeuGF5MpigyH8elx4eES265bhzmp7nCmGCFDk7xZSeZkQTw6VSmxxRN5n3o/ZRQUOGn5
VttAAN01zWVncWl+mS5t1SgEA0PNP4NgAII+Pf09qIidxYc3npSdwE60iRu6G54IQWxQ28s/3XIK
oaPOPdJKlK+hPFUHHSRIRG3B3qkCh7qEfa4Fmkfzt9el6UE9cnXVuLmUfRB3xEpGMGZplA0Y2qma
JFeIiozxLeTLkS/fZVjsyvqxQ4PsisHw08jFnIZaoc1jVwgOm6/1BjTpFKjTyZGNT3VEGOmWugrN
yeeZq1qFDd4jQPGuX8SWR0Ggm70ExrnkHKzM/bOA0ulcAUln9KyfS/ZMKL5WxXiggMsu0Lc7wHSI
g4mq+2eEy+wf26F1p9xBFQSxsv1H0JKjiKM2WuhJyDFYGbFH/gCfNMmOhSxnJY6/XgtZlbA02AP0
e4NmVpi9JTXMiLtPGcKoHU/hev4yFhwWVk706p3EzdiyxkdyJIlE0vTsSntdwXkAv5CPe1M6UtJs
eOtRaXjNnqSS0eHKbR383Ox/Jd3WrYD6IK+z5jNXxvRdcgIXtAQpCHZotCUsn/CrECCABDeAiaq4
2XIn4jGWbhskFpxSwtq4YGD1siljz8Vnq8iaKZo9QJ9+dDPotHOvEWO8++0TwepW9mJ2M+mHq5J6
WJ9tIh+jQtUr21xw8QXWhl8FfSBK2fILtc+N5c9+2McNeEekgA6Ym2tw72Qz0AKXro40iyeZU47d
gMdhXIdzlUONjl1rEpNqO2uBd6P/F0pv3/o3ZmkoqCNa05nINDH6fkz9BXh9LVOeqj/yy+EZ2wZB
OcC5d71cxJbGoedKRkBSS3yVp/FdqDh26h8jl4a0PzSBCtwbZkqeanXAbpfOu+MY8I/sJLY9Ty3w
gstxrm/hj0HQhnOCHPfNx2iABjOFrAK0ClakdBD6q11XJiv1JBSw7g1rB+QHiXHfTE7L18HlCvYp
JpvJxjL6Q/lciqYrSjZLXmV2WXfqfwW00TitHpyaLVWFm8zuwV5/EGC0fHrR+ydWmS6TWbI0piqU
y5yw04LAEOIFka4jRWn7cQt0IknQz//8jjyQQm+5Lc4dXTwQz7VrZ/vmnvEMhC8hbKWtRcqPwZ0p
anS0YlFPKUDOdRSxyNWXLZfBBhjTwmTW83WDE6IbGGcDYd60WvX/UbgHWCwZsNourpFWN5AzHpec
yG+GKTzwKRUEwvOD3uhi6GY5Jp2X3JNwGk65+YvTyZJ1cOtauu1RVTVV3AFeQlFSS5aVZ+MbVFDC
E57dgHzMP/t/QF893EFfMoZY3v2mMw3wD52bVEBfhPUvYM4/avmiUFihXQ0jK41RDmNokX4Jh1SL
5rlg0pWMp8watSY+PV09xTXBEVQGSwr9ITWv32NmYD+8arJeAHLQPspvoEwpwb8GBzXgrU8SMcRE
ZXhKgCP/wrxl60n9IZLiPFE9qw88JFz31Jmwn09SNNMcGSsPVctcoytejcAuiWfyZtz9N1Rm3r/O
+t0Cq73uburpQKXd9vsBUnSC04KsKlayYUhM9ezQsM+ZNk1+QjbMSsRVxqoJmZIiDLPGHKOuWikp
zmjn17qjJBT5TyNPGDqkAwXitwobCsmbKpYGTfwnG3TtIZ3mjz3Z/rgImgV7QGNo4ILOCC919h6b
U4THjsoCcZhOu1nIiEUxTRTLdxg1spkM1SNejmAT1GuaPSIutcI6hIYN4GUGRh8nqJgMxd3XddkF
911P2isEcWv88QMjOHvGh8yNM5lw24CGdByz01HRFvpxx7dpi3LEJXt7yeqSgKS1Xdgp6yws7NgD
UeeNfEkqxHkZhfZRSGQZRG9/0MwBqcD+L/1P5h/7RQyCsSSAqQ/Axc/bcmwrf9s8mQUPMUrc31Bc
c7nLRM0HFwB6aAD0q5AoJkBoEjMFsUjRiGKDsJ42T9MS7azvVG0xOJhOWq04zyYAe9AyUKLBjDQO
rETRq6VgoenRo30fX36aDiZDANMddILWtO75tN/GqMfu6MGkzwcAC/bP4BDvex9e5vU7xBCVbxXM
bpwFU/lJbYA5oHib51KNSnMcYQcz4EkEfZ7N1L/BLQTWOhkQwL8LI8SLBPi5Xuxt/6OwV6I7Ijj0
bZeVmzTvHp66/CsiJslDA1q2jUrcoh2MHc71PNZQS48GnENgGO9hEJOEbIwSJBr4tjgoRoC3Fla2
8tIGsRqvDTc5BPHEJpbLs2ASnvnHA91GERfkmvs7Wa80IgNQzyZGMn73d19Ijj7kbjetrJCo9BFb
jZDgV6KYn7RQXDvM+DUALjQEIV2MW3twarptxxZ2riFqNHeka+z1ji3n7vZKdKDb2sEE06YsV074
WLgR38/Inu5mQn8b5TGOoEFrp5Sx8z4kO10YpUd1qdbh2Y+CYyO8r5+Wh+CGjxXJNkEGbwbP7Kvs
dAuihqtQbRUjldVhO+sFntM4InXjDFfIGhrPzZQszadFl7W6u1AMXRC0kY1x55SU7g1axlVEIi7A
MdRBNRsMHH+/G1LffCKCKfkNr9SsujWB0itTFN39Sz8bc9eoaxQOmhbni3YGxlStI4qlbVAx8Vv7
Xzs8Q+d8LMlQxRfxyAVh/enEbuMtk05m1+xP+Z//B2cBtFhjShfzvx1ic+p1bUC72+6o06U2NFE9
w9YtchTRlz87QNFJZJTPDG3G7c+EfUbvDNwoMLd5zhKlvEhbSdFg5WogbT4mT0tQGoOwbQcAhMo7
DvUz/XfYAZ1w/iquaAXc0RhwxAxxKGhKurMNisKzqwhE/VLOnYbl07HN/YIDG2woYlyddWF9/MxD
JqZmu9DI9yJJV1G1JP56neCnyrAgn0s2D1UJEnFb4pbG36wbMhQ9BYkDdphJfaHfq97bLgTxpEgC
PM/n4NLCmtmAChB+sRX+b81GZfNqORMFVO6JPaj6pHsyIxsTItO6NxkzVpvQjoazBzBibfVWT8/A
eASlcMOqrP02OvhnMUuYzlKS256w/gk80nDsuRnFjxGeGjErWSvGSyE2g0uKOI0aO6rqNqNhu/xt
K4mPECfYOf+CfKCZmsVwruXKVCQzQWeLAnwMS9K1ZkdylfTiNUMZoo7uGi404hgaupLift4iMo9b
H4httTbDDyGvCCKZCHF4tmNrNl0X9I7UlpstPeegxyLRHr7HU6hQBMhMrYRgv6autD5jD+pbQDgz
VK+07BgKWK3rxUbRCmu0Un5PJZiCKmHBXiEUc1x+FF6wFteTPZbFy7UUX07wkFZVTiU1L5VKagmm
cNTE3s53ExpBvE15bO6pp3APiMwTT7vpAeB/6/dy7xzCR6zomCqolR08XL9zckkMp1VTF8oSZS1j
yzKqP5WTnftxmLNr6abPPSk0VaGa9LZeT7UNQHYBshixTzpSqMaVcEI27m7BCPVLb3gl0VXjdatw
cpIIKRkZ+CnEer6o+5apQWlFcyEBRkMtLqIvznqFEFnWWC0W7AIgpaws7oLDG0p6scfZFBU8K0Cy
Y9OImWIG1ooZlmG2VSwPnM7Oe/k8f5WJO2NX5g/a6LAkzyQz8+zW15uC/wVmugVDBUl9UZktulgJ
Y5FHyWbH1Ed7hnFQDvmQuiGg7016sDrrDo+ZoDm5+tJuXgbDBUYouNl3TAMwxW00vxYXJ+LHleot
oPqUmLqLlD1bbOhE9KTSDf6U4vVJ7ca1JEo+G6SK1zbjQ5fe4p2jr2zkfnWrwE4tQ2iB6ZNpPqWO
bsWeOqpSb65yZ0EUnGynlK6TJZwcUXYB6DVcOaybwwCPgM1OLHzOyJtNf0xzmgA9kVXWJ0/NqN2w
2aLWUBxik0z9vqWuNSfPgfR690yqqA9pj8OqNdxF5wSJUs9onsSP2YBbRha95AohWF/wPWt6ieKY
Jbc6yLC8ISYdu2rZghklmWxlcUbMRdkGL4gYTQaxYS/SyxZZJK9qD++6sehkotNF37ZQCJbNLJgM
BtFY4dyfQhvAJd2FtS3g8hFBirIqFHbtbZdwsY9B7n6oURiBET26dg5XS84wjdJH6A3nmQxa+c0Z
rrGwoXoHrWhhN7p2ojmYipcrI6ibjLqvKpDJxr1LRsCjdPO3Ch4f7WRflGpD5ij15e+uSaZeKn8E
GmwsA5aThBTvKepQNHrp6i+gS4F9J0M5ikb0AwW6r2TP6buh1oHcOLKpacgn8QdtaUp56f1Z3bHc
/GQckTByfruyYcBQIqkthnyS8Ev/aKu8qEVWMxOILeIFX0w1HUgQ+WZqwxdDyRYsEZg/YgTE57Qf
GhXjp9tDz3WSqgJ4LWgTm4xiXVYmIaR1BLFcVehbimP8aXKFY8My7+Or2d57rsaRuaYWypX5GM5q
sdEsDfUa58nx82oNrkFZ/y+KSDR2fj03U58gExcQ4Sf4Gn9ZEcb10bH912x0Pl36hRFqdmXTJXCX
k9xwBK7wxaBLfLx+JJj05H71d7ZljoS+wIxBgxgQLGQlSpGJvddKYZiVh+QgS231NvDmQGGcEd6H
0kxTXgeyvWlk7+2zPN+1AzELQ6ssMEvywjHMPwOCizjaHRCnDCEu8TvnRx7ammxyFWMxnqdKJlV7
HDkMK++wwlnJndiX6zbWs9AebRiXmyBO0mWs6/H4nEHjgvUks+4T3Q95QFY5OXYAxkdXzD+x3X3g
J6V7398Z2A8gENsH92XalpLDokmJHvWdFkQg2xkmikfk2bVCUESAyzoJwMjZtT6uzEEnXvlRa5D5
qcEjQeMn+At8tqXJWDbTOIxyNGyLlOXaaIODgdC5FWCS598EGwcGtppYknkIfAO1z5uoZjn5nQb9
zklP6ZTHt0SjSvewFmwoWHd9piPhXsfJJqAV/+3phJsK2TQower3cg0qUIWn1b09doKwk866vWW+
cZvJR2D19nq9w+QPLxI7khU/ErQpG0EXJ/JSM6EHJAGUXwxGBxza3IN8fyeYR5P71XJuTaJzMixc
yXX9NseoxZMy5CCWoFWULbPf25/0bM4k1LWyM+oZj8Ft4kOdzXYBR7b0t12RHNR1+0BR/QZyvy6H
5yY7VOM4JBG+P8eWt9bdeTthKlxopw+hlTVjve7CbhhKcketXhGZfWPqiAy6BHIy3qZ4t3WbU95R
6ndUlW2Ptv1sDHUWyUYtCyf6RDcMuc+abDUzyedooMZka+rgNAKxMtacXVNligXpd+Fh+bgiZgIL
hqTkh0Z9HaqGpfdcvVjPu1n6B5rSFsNqM0rwKeH1F/duHyxv1zbdjrULvqVyouU8e+v8L4LF+4hb
zFRu2XMTY8jsnwQu3iPBq/Um238H+BASBtvJecefSH9IHDRijxbvRAaaHufxfIdf9AloyIOqt44Y
y3q+BCIGXpocruyIksZ9iaqwfCLwMR3GN2iNL2ijNdQsjumjSh01Dydjwa3piRwgZ6JVH+Ndu49g
3hDNMYawC/Fz/BUXE+Ao2k/C36UnrwuQMUXRfX48+8Ah3/e7/vA+utge+rAj5Jcu1mxTR9x5gUkc
66D/T90DreT2K5mTK1cpI9o5izN+a3Od1ZCiTGzQhzcD5KWX8dbDyJstHIokck2O9Kmu0TcADDJZ
aYL3P/Kls3saa7I5qBx6+D/eINZcgSbzyEzuv199vSUunRSRnZ3sWHJzWTmfxX+/BKLJOg0SY4V/
fcSrkNBIMcWKM4vbodnaqUwE1BZEzLK4tyXFmQOngiCqn7bX4ms29jVUnRUzY3qoCfnGwa/OdYfy
LFO1CFy6I6LG5BT6qWDj8nAhwYY4umzp6OqQUQyh4hY1gjXDWB0V2gaPAXffeakzfkKEaSMC2xIm
N6KDNLwB58HDVOR8lV7EcQep+h52HMDnwhmWLvy432iT7dGTLORTfAalgSj71LEUOQE03tj+gmQw
swWWP4nGUJKcwjP19n7q3PjHH7Iwe4EO7qSo8kwUQ3UzJhJxSTQYh4QLcYZM6lciPeMjO5d5Uk7q
OGJashvj/VPnAGxJo1cI9z7+tTKhtx1S/ypifIJsqfN9FoHn2GyqU4S7x7I8HpigY3klVja0HvED
HWFpeF31ffnghqRYvfzZelKX3RqzTrD3c981IMmHVEcRXqSpNUBv6MB9uB2bYq9N2ije17R64nw5
h571cz+2bTTiuCBMBCnB1DOK8HPzex+Wafqjct3SNYb83OKXlm8kOCcsTzT69hkuREWqcYmsBDJT
uPxf1aexBil8fOMde69iWoWRmtoaXcoQ7PqsG/JHSys7fjI2oxZNCPM4LmYflXC8X7spKq8vrF7v
x7HrsEBJihNxIsdYLaZ3bvbY7nABPTzx4ZahzGIVq9Ap/yCAHJwGfBdkVbka9XijcfrDnWh1Tds0
lMMtcYpbNhfbv3PIz9jrr2EYdlN9sCKMcPgBj7pR0WsiVLCnS5RKppHvhRhAxGMpZzXWUeUBgliW
yA6m1CULiIqEmRw10ToXLKqiZge6CUNXeyrmX21BDiRnRgpoJ/81N6uC1kv22ooq04kN04xPvJcy
DV4QGdbv8MO6xjpai4rhkKoX79ZGVAHxHYUm1LQP6tO7n2lEN2Uy3jf5gZasBYwvRfPJAiUThnt5
jbt293kuJWtPeG0Dd5TENE7GWZl7oDxyKsQX56mtYQjhh4xjOrL1bFvU3dCrf6ypLp/Vv2LOrEcB
v4wyb2ShUUxKhEJLYGHj4LOJiofE37hiJHwLAXiwDujnnvb33Uysx7A4molURlAB6xRTrEJrGwu+
DuIIByCY9rNYz8Dxb7uDJfn1HPgHXPjwjT/vUN8hTwUrui0h+s2Ey4i/waP5QjU9Ki7b0tQbAxth
yelIUQpnriO6VGH7x2MHVplNbAkqx50Eg7KuNQsOHZSgx+tXscO/fWFYPDc9LX4MEB+rhvP8u0Uq
BbJbmIcl1DXMUSi5sV80ALIT2PTnqdra/jEjGw3QlpNE92IW2OqkTbFNoIxOBGQPE+vznj/2Pwyt
OaP4bRQMGBiysDy/bno02h9hjZGyqdrjUeEONvn1YxskiTKHBT0RrucSrBUZuxiXa30UwppLg7Vj
wivPCsqBQXySWDa/d/oJotjoGUN/m8WTKcudfE7VxBl199buUuxRWaHpCyKBcDnPqS3TYDjQ3UC6
q/KbgroVykku1+vTwRYgKMNMaA8HUM+9GrCaCXQVHWs8JKpFsW36mdcs98ItuPGqQPO14YAXcPDf
A8ENlrBb4hzq+Kip7GTX9nW6iEgg7xkzG7gZl7uzzZ7igCFCjgR3WOa5U8xa1A1tbro7QEdzclp+
aZ0HnDuEcEiNN67hN1b8v5eqZY0GXS8dvJXsrlPCecunMRvOYCVk88QUjkucI0GTRAZMWoNWWm5U
UXonUZmh360xcygBW7mMkvXI1a2iOM3/NZo1PcU4lmzg4aoYaPd30NjkhdjhjAsGmuLnue35nOcc
GiopMBT+iFcw/pSQZnd3IBA+bl+g8uLKXlOTngKhEOKYJM3bgHnv8lblWm4ZLeZ0lZ6YbmWIjsAo
1HbtegFkL1Bm5yLTE5XmB46pi1kqm4DwH0ncIdyJnVEDZFAmalY9KNQLj44E4+TPfugga8eDU+n5
XD1rnUYXPa4jDBEj7yW9/IM+ItSUUbihK4zZvKZ1+/s3VfxJHWp2eUJ9HyP8O111XvT57tjaDB3W
V68XtBcIj8Th+VfLh3nlcoZSHd/rDwo4elk4l/okk37DzxeYkQ2+pctR1FUrBdNWMwHsY31iNQpO
yzTkihJlHXdzme/iv8J9jZAA+7YzvlJCDRNHRKxziVkkX2yuSVTXxCaqXR1wb4ZYDGIIqL+IbhVi
E190v/XIcU65eMkLr9dVSlrdevMDnGV/J68O7TJ4BPWD2iHcwIkq/yi7zOrYYmZuBOyTUlSqTggN
3cYg7BiopEAP6/km6uI+tyPhkq666GMZEnDITCtNEVPC6/MWE+Q0libc523CV2K6jSkLGipyoiPx
4bLTa0gtNK4Kzui4NdCHdUYUBL/7ydQKXFKGqhpNCBNMn1G0ODXxu3bC4XhBef7WLJi+aQy7ZKp2
hybwA/C1q0ZbOsHGcUqiQfxhQJgjIwXPTgoPHv3RizEU4lBLs6UrjJHNjsCHcOo2hpqBbM/Nkv3N
9Ox0Z1pum3T4dtVbRtfgVc04Zr/Vv4owlKOTplf2MWR5+U3uI6VmzYy2GIf4obJvjrY4zAD7iFpP
TE9S0Lue53F/U4YiXnp/iaH1KLXFnbFa82gbIQkF3XjUj91VV8UU5afzwf1lusXpv1zSJnQfHj/x
3Zt6ehD9KZCfg1+ZsaV6lcJwU7iXR2frPvcrnKgOi0I+Nfh+9f7W8Igxz4hRwhmKTUpoNfrKDhKY
EhmO2BS8H8EQcuDuV+8/1Ao+qztN9b1FLDBr+NNVikIpiUuKWmp9u2hJIr3tw0byW14IwCcMatbg
7jVRmQo1My6x0Z5LI5hk+Rcj8h7yahr/jkxIBQQUcwmjrMqqAy9BJgcI2jepykg3wINDX6MFxmso
KjoNolIOHn6G46WwcEDtn/dRhjVR8r5OiIC30RngOMedzQuf1YDtqokAqRDK5o06LOXUVn7iIDMd
kWHv6qsgN5KV9mkpMRNdcLJiFtBw+xxehqI8K1GUpttfc5ZVNRag4Lku+brY/4Nn9h/CWWl5H5HO
fgymuZsqVknvQn36pkm59o4tcpnxYO/Zus5Q5+kfARkKtaQwfpUmmk4S4B84xDTfml2a4WVQKj5J
oF8Q0Rptla6Cf6fSCnOQcj0JuQe8nUnPkx1Odn5GAESW30eToCU7FzYy7DKXzYjPGKpqKod19Fec
QLKfumjYYcQ6DZ0p4gf81TpaKbdBI+nlj6tlYZTt5zfDcV4z9zR3lZVeRe6NVA1F9J2i3m9seXZM
Nhu5+P3XZTp+ykMTjnUdkwXKfe7RMfRPfGBN0N5L0WnyD2pyc67Or6X2ESLhPgNdCrUGMPe1X6D7
kHpm15Rd3pKFAvW1XTDC9Aigx0HQmBNl4kHnhtFGkDEDelIbLc7J283oEBm26N16WFAbUHddp0Hf
xmZykOLw4cPpNyLXYta+IOX4tyjIDT3X2dqpDohIjBEB/JyGMcwim2bzY4/wiOtu3JQXSPHRdc1Y
dD5H4kfIGvkjSBG36eTvnNaG1vOoAtkv/cokHa8i1gH5xIYauVlhF8MGWldis7q9SR6h8WEW9Na6
AP16zQbI7qcQpwoizGlTBJgLveoPvgihsbl7n/T5jXhFJ8JrUN3tQYJQDYDeENFj8ngUPNamI/ZT
39+fV6wRlvpu/x4Z5uT8E3x/j5YfHtBCJt5s47kNFmGRT1cgmgOYxXhj494s0aKU83ScT9MQw4Ui
m1BropWxnDoOJqRkf4QCGP086IpYEMpt9p4OAjoJfh7KxDOW0xbrjPclPftWITXdh5EDJYBZy714
wJwK62ZMhZrxLC6cwDbcb8lWwtJWy3BuYdGmxsGlVfbN0bYB0flOdoP7+vAcEUph5xvnZmPL4s5r
UJnrURlo5Eo0L5VOdRtPIiax2uEOfrcj6RNaSrB7zd/uS+VDKKj8FyBOrEIye4rU8xsAJ8YdnjJm
KxDhvLZvjj+AJGMbg/wBbYclG4SISsEwAQGGRqt0jcaxPiPiHqnQG4xy2C9Dh/xHpPZLoiar47Vg
kDEvJvHZq6CJvNxP5xGeSCihBLIqyozdTGPV5J262JSkNDJIwcATWpx49PuN2N3nTjOOxhdj5BPU
Phe7tViggIsks6RPiiVTTkNmGM2LflWP+jwqop7m7kFrRnfT+f+E+zOpLbVphyWBipii/VDsp9Ix
PTzHa6cI/CB0hJJx85H6phHQFT56Z2dSxCAlVdEH0IZA8SIVJDJIApaQuzJmtVKdKsPpVXwnj8Ok
9fU5ITuIMIz8wueqRSQ5C4FeK44c34oVwyfwDRrdHPDhgAuaabIjlyIcZ/irbihfg8vIPXcXqx2c
cCzt/C3ZSF9+RwEXrvmhr3yXAzJC40BLTQiWzPT1WGJpLym2rrdu9BBYQExXWZYaPVbaOc+aVT10
1CcWE0L4DOI51db7MAgNz5hpgrdZR/lGIqaxgUq7AgL+OYkJx5ny8xlPJ23dBFHzip/CS4uGW6+6
Qi4xBGFNqXo6jd8notGuemMedR+qW02fOTlcVaS3Ry5wD+oXbkkj9f+698uD7+LPmAFWSfXCQBvI
Xa+O4kZbpM9hSdiRhT8znOJZInNPt0EJuJzHmfBQJEHNin7fZCb14qOtuyxMmdTwBxI2fEfyiOkF
UmHUGyqh7C0gF/l1B4Mxrkb7gnQk44bRHsJNK/1GpHVEyoqbEYe1OUfILB4TPaiJRrpMBRRJqvRG
9WWfKIemUMBnyi3v7CktjagRIpoR6SvrXBdwkqqNPo9DOYHoXjKxuRkw48WV3MqAYZNV8N12P61+
n5FcUK/kPPRgZHkfXcQ9K+hXBSWbOVo6lNoClYhM9zPpz6aXsGg4VdFWWNYgjRfVZ3DezP5zNEVW
1scAdU+owKImJekh+b0LRXXq3u5FxZ5BQsVm3d+nHVUEOwACw9mL5I/OumAC0P2m9mwaRuFvh/dA
8T7BXrmCV6L8n1KcrND+3O1uM3aRIkoWnHR+lR5hdjSKknahrxiZT7R++uZu6qcQrYwPTbcHujX/
lB+qQE2mNGrLG+OHbCx7Higp7qlhc1oOO20+1F0zl7xmArI8KLCZ4ZsQeUxDVtPV5Z5rJMtdQoij
th29aOFN05XXJrtvwz0uFYTjmOUsKzs3voCOSzqXdReDcOte66Pkw0CkwESJcq2iSTCoUBOfShJ7
d/b5MHZ452CUJGAkNPqIJceKHed8KUHYaPHHhkbJhmR9qyDgUWJq9dQZlbcCtWv3fhLzO2i7pTqD
v4kNHQkEA1c3WofSVQ62avDH53uFfTWpUcmk/E74KJXUM3L6sUPGH39smWeDcp6FDdRMHMrMUE6v
rIAIrBdOsXvcaH5L9lxzpEXihxOiuD4qCtfxrwnERtM8/b+KCkkkIPwQs4qJ0lxajfy6xjMBSloY
lPzJdkh/FdulE1PBsq2m6fAB1nWTn4w/i4KtzBFKAgt+4N2MWnJGHEMzWhAZFAse23mrf53BV726
71mmt6BD91Orvd45/oGxWpsdLnVbOqfuuPkaetBLKCABzSH11LPlSFRNXr4/MMfsNLPXeF84Lrqk
pZL4JIwk8fnqftrr4GDWjmAjyOyX6uYk2+RZv1vH/OCJmikJMuTujTzBPRx0rYlpdJ9M+GTyhwF0
O25nCqapSY9BuL3GRhgHBXYlpnWTuq6BFwJuKv8ap2pTBqvcj7x89SwdLGYEFgZNx1bOD6HZQgNn
WuX9IeIciL61FmVxHCxX8Idn/XrEeFkND/o9IcSlKHmFzA1diP+82CS8ykbgRZr50HOBhOQXkKBF
jHWLR5slS0APbtmSd60uQcTr2C1nB/AzJ8voi3psPiF7KGLoVEPiz+yseK8HyC1n/NXO8A952lqb
NC0pnPiV5g4+S5K9Mwae+x1NZFP2rGxG9ldxBP2BrN0bt9KGQJw5qsDvKn5KIdNZTp1yuqmAriKr
6aOe9lNccVXydSTanZ3xCqV7NJBG9vAUeX0aXcpGhOnNggLWwfCL7n8QC/JAlqYgVmP0UDOcnsPE
paPH4ytu03+knwd9JoiHhjI6ApYe/dEIJcqkRc1DPckjroyfAVDpf1y6z1zVeZu+cUzG+TL2tngo
P7YAGSGwC97KDqsMmIRabMRL959ALTznJuRM1zZazsQcrVT9mqXsOC3t7Pbkh5mkZAySmzC3DqcA
k/PfGyV8GvJb6ex+b8Mscb9zvlbjpKjqAT5Zl30jpBAksR1xq4m6Z5ahScqQs+ITVgbDV7JrVOrG
fZ/wL+sWfXYqB9ysbFG+qye8sNg5RHXFV9Z4emTBplc9bE8qwMdXX0w5Ws1JPibNCGBI9JHZmqbS
ubkQ339LY2FUI4gt1zGKR8NM/q+a/Rort/1asQHm36uY16RK1+e4pKB8lywgl7R0Qw4mLyWHJuhU
sfusrS+/fJt2gqxhqTWL3PaL9iGTDmSWPrvMp8tciXOb8MxBH3Fzg7IApbW4yuao39f0x6PenJpe
1TSHvs5UubUh0s4IqApSNwL1prXvPpHkWSfT/Mo+S3TBzW02JcL9II+nloJtZEobGCBYlpevn0UE
uHk/9lUQF/+79kl9cJ8E5OvjLv3xvXcoXnIlH5n4PQw8kWx7dPKdk+dLh8aPSGwhcOuywCbrTIUU
AYKRNVeaV3HIZZWtgNJdLvxMe8Zt5IWuksKTzHqP6Uqsehpr5gjsL2mLGvA9rHZwzV2JRpOLM6DU
ldVPd/zKTziWWHKzAWUbiG2+Y6u9TcDfM6dGz0/3+QtVd3pNPaZeclCkRBs3qMhtKltWHnErO0me
vfsfunU4bdCcLyzpYhFOgefyalMjyT4PiqrpqIQykDeof4E/ZHNsX6TuZ2OUcdN5KVCPOI/FFbWH
wO43TTPI6pZWaVZlxqmYnlQJNgyTwEnMessUj7JYbGtuyv6E8hp4Vio/4JcMNf/ziX9ILGNA/vtv
vHhe9MehLI8VdWz/W93UZeaZmls2qGirQzmrBz6pQvp8QhqMcRau5A1d0AThy0UWxHfgMnHAVRuW
FBO7bqwtfVHfzqz9V2Y+eS8RshkG7dzgBgbbL5FXMwDqmn4B/1gLxwBWjr6CTjPk20XgzVW08UWZ
SO1YlKHcTKEaXUloRlYRXkOplZNspBK7z08dv2lCgniCI2vJScgAcAZ1OC0xDyO568fh8CxWEqH8
kvj/fbYwmeHULhh7Ac8hyWf4CWd9uo3hV92vjiG2lUNeh8qmTYGkEy7aU331hpV8zwsL5Po5ojOC
Zt9mS+tksxTwmqZKjg6xbFDpO/PixSgmfXzkfFaGuG71jHis9G1ubxB7F9nK5Mw2J0Ntb+uCrH6o
SdzTGRkYdArlwdGVgqonCWfsw/n0LUZfm+Oq4owhEJ3ObI+8eKycK9bTKlzycJQZTMpg9R6amU/W
wuiKFzuNDinv0ekhk14jsWsTCyQeg/PPisB5j4Y+0P8F6pPCl0VBECqtPXSEbar6WOmeRhZct/21
lKh5GZwSn8hxUwRT9PAgcs0O3wS0tSeENfSoMh5T/EEKbUSKHiuCYdHFo1B5GqkYBHn00TAbCaTI
Texbya3PVQKMh/ZJHmdHQiPjcdt8y9FYRUqKWfnOebBBLT+BDzwRf/0gXTQsr3Gi8dVNSfUF4KOA
5YBC23QQ5niKkpq8WtfWUCIA7+EG0qVxlCrLO9VXU2mvv/G5JX5mxhflv7rKINrZqGRZz+KeIGb/
LHBjB1MlmjZ1Qo2w7jsUwwyG6lM7x5edPHlX5KkZ2eaUX01ywLnK8AXQekXXqhYFNoh3vV5lSnLY
NvcQB9Rmsn2sbVLn27FJ6Ur0xDPnLiJ6neC9Xuw1/2UbUjqgL1Fa2pl4ekiEQQxiLgbcPadcZJt6
Fy1kmBdpLYbJ7+KI/ezC8sXhctjMRELASjQFfI9sTA3usibFcA8Ny9dZrxkHjomqPGhHVGnc3nNY
kSnYfPa5OYuMkxPhUpjLvaxsO0X6glKcD1aexhVQ4knc/lUe7+FFCIv7z8BsnrWPVuiJ0sXkGjhZ
DgFFV8CbdkBueoCpM9Kx2378jZz67xI0wTRb9KSlXao6xLHOP74XxCIv/UdDrdysGC0XIZXJwmED
AFVFrAQ12cgtsqTS5vVhDXX7qv8NV6Ya2y2E/iKDDclR7H6rrmCITEL0m+5tnNZSubZEEasifRcc
1NZNf5TSf53CEpzbHrhx7cd6y9V/JbeZP3ADcSzyL1gSkYvk+9O7PZqALs+thHpfWHojarUhID8E
vaehpY3JHkP50VnqK5ltTG3bHva8h349aE6GtwoTaOicQASQzrcFHd3HlIq6unvT3VzsRTzXGbRR
rPTh9Dy7H+XmIljOK0AVYIjZRaymbUwtyQNTQ1bf7sK/vT0LV0+hr3T1AaJTS7yPC6rEUXCmwqfk
2N1Z28ka0l4K/VSGXlwwY/RSPPL7XBt0mfkDLBUCn5tT0l3dFjR+D0skVtDEbs9a9x7a+7Jk0JQW
/W2CvoDpIzACkjp3vi43Zskh+cTZ6OjkJEGf3DiAAVwXCohczyTtMhMVLbl6dZeqzwQe0FZqR4kf
lKADP0kmTMB+MKbANPmZtjdhqZzPvcyeKYOg2xe2ho77iD9Mm071HNqrBfMDr3XuiW/QAAm8FnqG
Ii/FV9RFeh3LQQoUeapOvsQqFCQt6wsOavsSpYlhJPVI48R5nHRi2f19F1E5+9d5MY5q9g1e1O0G
/0uwm8FYjR3NxtwlBgaucBWXq9vwHE1fmNcS5y3k/KwkLzE6Vy2ezG0zrIXkyrFpKFwwvNmGrbYt
I5dia/5uWw5SQChuU1P2KyxkgU22CjdnkIU43pF+knNOUofR5fjEbwMbE3b0Upw/i1tmMJ2t/zbT
D1VcmPAsKfro+sof6HmgCFTrfmN7ldvc/cxpJdxYzJ0H0hCg3KecTPc+cv0JNcxESHT6SaUoje7n
zK2cPU2NJht+IoGwz3ynJQ/GIxSoP8o/S7nyAgCCiEMO65zOQL7YNZ6K945Mc1qnozBp2mqHopJK
vxUNnV/1S7PcHZf9qN3NQrOLWOddKTLmUTEgzAAyy+Cj3upLXEy/KvOf2RHVNhp/pKcTBuD1FOjN
defjc/EgIUDc28AtcyNbx8zf/TMS9hdXELBZrwOaGufHx4V4959eg+TQ3o/fvfkJ1CDn9euYC4h8
BFCmOhza8tsHjXRft6oCF3VzbKao9ZNrK3W8ahYS/ZOp4JFKgsqlWGTnR+1eFUHOARRXdn2B6Bh1
QL2c1eKMvQsSmBLOCu0T++35wZLRgMdpZcmxwFsKxiUEBmk7EfE73smfkYP2Kho2ocaY55HyCvv8
2weAPCcZeMV7OP3tSxCknWyUj3IeCUWXD0qtev1lPJUNIGdhFKBq8rAzQVEVGJ9xcc7bvzA7b1u1
vVAJ7XQWw4IxWsskgK58PysDNeY1/dIV/+Sgt3Kuw0IMl9RZ9uDs//4o3cqgd49IUkspKXs7EREA
61k+KoGZPdzUKAbUQM2BEpTq+ZL8swkIpSSXhpi0VXPGEZxglaB92DQUpzdENJJF4YMZ593CJuuP
pvZELHS5NCpPGGPxP1GXxFmHl/B2nf1y0CsmBOZO37dIrToAhnSRQ7/5LHhYMIWRjTpKoPnjmwxg
eq12vo/opZwmE5CLB4jA+a7+1O0vp/luRoxZ+6z8IdnsT3RVKyihbdgVGJdXQgLcVNDp2xaa7i4g
reuml04Msxp8NpA5ZjNKu+ni6pQagGwTzUqA6tKWiCQ1bENEVTPz4CtO6Br/sIavIpPV//iumkRw
7cvtzsYuLCFQWwjKig0x3Q1WaBc636YMCt/RJVYOVFBjbwW5mzlDZSgR8OZob7UaYB5nOEhQCUy6
XWgyuCUOWW/2BQHJyGlTZYbg1fekJ4w6xmRp4Ftfel6RMNsW4Xkozd+I2WGd63kn8VLWT3f3M6XD
0LzYnzM+sBICJpn+vOtVNnp4UDGkXzxq8KvQwQ7daHFNNLSajifPa+XRizdLTBmhBnDdaiPW+vfX
bsgFzdUGXLde8s9pDAyQr+N3p5Whn00aralwTmXZRH7NhZtAuA2Bcbi3ibH0iD7n1WwmoCNAIvhZ
GRNAN6y/HccS+JHNcy6Y7UByeIbOrHnU5GTgmZk2gNNBQ8gVM4uPL0zAXfWqijjvuaMs28QUCRaa
VaIehiy4XnktXMKaDcgmWPbC2pCz3+1SIAXebAJD7bJpNraZCbI1ZGiZm/3cGWzwQxWbNFeHks6x
ENHTLxaKRGQJBQgX5k6m7G30z0YtlQTRiRCXbOVBKeVbFE4yhzZHenvhijW70bQKL7uKqz9rjHFb
BS2ivQSKmzKHNnc0s4OYbAP4ZZlg18ry4R4GwPGLfKKdejuAJ/9XFXMebRAzwFa+BdDBb+6hEPRY
d+MVgxmzLHAdyt2lYeGH6OL3hDeVY0tj4EBNeb5O4PeQzkJ84iYcBy3ePedSvBPkTE1jEgXzjTvz
XJJKYyrWeFs64zUTMqBaQ3/lSl36TxOfkI1TGDUNFxKrroKjMsXlrlFv3/Zt48bYI9BpApz2VQji
qIpvZvSAaWjek4vYAmXnP02qlJHJFQaftA/u4xzdd/NNvZdh6GaDDoGlgfhW6PrB/6++8oIvJTqt
kwBkd5T6KJ40kcA5mpkcI67W+zNVNi65w0Kfd9nrTB5RdNh0jrKJ8fmDl0gBRx4QG/NCMAqi0Hw8
/gJe0CRpgerEaYzJUarTU3eTIVWZcfskmbBYHAJcDMlTQid2NcIjhBev/icYYoSk+sSjAhh/FHKK
OCkczknVoXO9BJ9eWkLq8v6YCw5weWldtykyW1nCk3+y2JVP5pQs6q59SCLicCK/LtydhZSJIzte
anaE11F0OFYlgCwZD41ICM0WCB+Fgvzko2X86n6s0sWFNtUrQd/6khpJdvRN2JtMCn6pcgz9XuXZ
oAyme6rgQN65yG+DdKQHzgDt1m5lQn6gLwmGOS45sbwcTWnTtdCiBIcXz32A4eCrolbGd5F9S/yb
gn++KMm4FX4mmxk4yinqUJro9UkwfNmFT8kHrkFOndad86sXkQbMgC0YmDd3gtTtqT9wDGd3ONb1
SnXvJfvJ9qY2uFIWvFVUQFRI89F9XORfwcChWYsK01NVNEWc+d6kbdqtYq5EgGgIHDYd1Tx0iW+6
Wfr28fkAxZnrwIZze77AOPN0YCfTSdjVtBNVDuJQ2s7KyvGSBLom50W1TsQ+qcqhZGWOQ0AIP+I9
OEVWRyNiyBDIL6E83w1GZtIharJHMzdTKCytoTG+/Azs52sWYICQDBe8qg/81c8kYC1d+hwIW69o
jBMu136Dj8GqnE3/Ev8q6dO3wUIZ5b7Klat1vYF3my3pN65Bd98+3B/r8hOTorb1MYczRmJ7Yuu/
ADVzSvKO3rwMCn+vcvpZfHPG4kmozM/8G+cFW7PbumYBx4i5q5C8NGkiA/G5uSViveLaFyt1GOvR
wpEr5kWY9bqeNHErbFcE5EGmFCEyJUoLzko7mIT9ms7s1gVgDpi417sqE0v8VMI7jR98tIUsOcEQ
+BzFhVds/DV+R9Nvcx6kE1cIvPsaKz2WctT4wSbp7qYncLJg14lbVSDq8HCzSJ7GcyFFNO7KXOrv
KY285O5n+kpkapZPSBg36KwjQK/zetsvkO0q2yFv5d1godZoFYlvr3kY7cnsKCFY9eWsApnLiadl
V64JjQIMae34AzIansXTUB2t8k0l1aqlw++RU2WORT7ZFTGUheYLnd1Q2pQcddItLyezrKSclcyp
SkIGShaVq9Q5itIScIiUC+YNdThLciur9srUHFhexYOhjkBoaFMpEtZDPpJ9TIKAUSZiLJH7IboR
tc2bA3MrE8TrbgVjTdsrYRcAR3MP+LXvJlly/m1tmbQe0KCKqgMF6K17jjdFjWCHIjlVkml8GhW2
AqftLAEyXtI9YEsmM1ac/k6M3LexYByd3oKvmth7tCsmWT1W03RAZscMXUgpvgDbKTZPeZQdqs3W
sgHvM9TxwPvYJ734zpnbdp/ssuIdHtjHwwQoDJIaFfOZI4kTn64rOUyLCE2TbC8tv1xVO/SCjukT
bLGLfDjmphGsfJ9bxo9Pi6VPOn+uynKB39kV8mxaKvY+nWSXZVUdHAgbvveBn5l7V9nO//c6CKw9
CBwf5HhbIH4Cssfo0TGRn+e2i2seHiQtIh1m6pAabJfyYM9H3C2CApBPlHeC8u2GSDJzWkaKOinn
O7rFmgab+K5jxx3eMDOAeNGrpMdS5VDvyFVHyiQTtC7A1iAthH9k43qlGv3s+57qK0q8XejUjyOJ
r+3Yi+ZPRLj7xQX5OawQc3q41pRpkz++7yUZvwSv0n/LsBzXPpNrhIarBu4fQo+1BDEB5zrLopwU
ovW8sql7YnR036W0lJA452jwKELadsaN4z1IcLVZJ5LRhyjtNdO9nCFsQSmi+Om8y+iHkBkCmqaU
7d0gTdkINBIkT2V/iXwbl5J/tn0feUANzwIhF2hM+A/JHLNCdlUVOihthaEXZXOTGUT1Vncap7eD
EWPSMPCv03XugGV+Iw3AP70gtqY7MN2QvIUB0FroMeqL/pcGTnDUs1UXMv9rNvAcbp6A/LXtl5vS
0Nd2LoOsORCVy4Ooc92GzKI0Ovw0qx+zG97iSuWV9kfErbOlQl36NuwXOVxCv04HCK7oi9j5G91n
OqvZhE3OCfRtG3r3f7baywY7XWbh3cBfLpPGpAk4uzEaU9Lu/OyKEoh7vIskxFZjqOVCjIQotha6
4/zuGyY+g5oog+CGNp2MqAavIevyC4aysUgAOEXmzbE2zfvWSt4HQgTVP1yPvaHuZxU88/mrOro4
ecRzZ/lo0rvXQ2fQa39leo5FRXFs9dyUsjKpigXyDSEWZMKkffam/NqS4q+ECf2y3x/i0vUgDy/s
8ooO5WpTnxnWzM8jJMQC1tDh6/qACauu8zukOdN/z8DzgJp7OLwwnI2k8M3a7sH7g0xS2lUR7+ud
mtN3hp+hinNTTbWV1KsxTsTisUsj30dgYOzj+SpvaLsRcHSt57zN/M4YqTM1nN6iPDtW0J5PQSZx
hD4f9Ry07InVwohLBFvMXHmgKnGtHaLNFTQGoE+BQ8mZ/rP0iPekNOKcnrzmh5+dQ/SfRmlfIso6
QdHsffOZT68sIUWaRGiZo9RoXHq6QZBZExh47OeCxYDFvWf8STWORr0KF/47Mjfh4WxbZLzPHj4E
728qBSwZv6DNZFn7Isv1IwQ7uSAegmtg9T4trJh8dHCZlIon/ZPO+qjvfwDmNW4YwQkpPHr8Wil2
lbADtVTpHXX8FsQBA22QC02/RD1dEmaT9xkqC9mAc6FwZXfIeUbla92rg/q8CQZcI2uC4cTf7KEE
T4jB9nZV4hBChTSpp78Ja8v8VRFZ8r2Sk2tVDm0fWu+msHwIqJfmNcKuL/ync8Idxt1pcdBhT/2Q
gS+5pzXJTB/SHS8g30yNrlJCzczcpAJMPkfbbgdRrFRWDgaWjaFbPH5S0w7LmWMOIXbiApCi0kdI
2hkj3PF59flCRizkZEQjQlCWb9lRTA/q00bd8XLJClD1em9tNBpunAt0H+gyuJ9oPtg1AeLhgFd4
S4monUskh+ErwlurepR3+mNhvVMsd0g73vtBybnOSjnVRxfBN1sL/0Ad9dau+WRaEkpE/pKsewDV
76I7qYKJYLq9pObRd99QVoko10o8iRYu2UT/wRCEfnJV+BF2lwo7mPqP9tW2ypx5XmuvSmDbIkAf
EfNz13Zmsm0en21gWZqExDNHNOZQeEC/16sU7IBRBasVn5KWSXLAlakuht6TQ/WYNRuunWsWMrRP
QSaZwN1mJvzBPn0D+7hclLhNkn8l7oMvmrinugXj9mCkMPVP2MBK0JiSG7dXDp2uQBtNdpQRooJw
Fd6Jyv33APO1xbt/dpL2TxY1KHoESiCk3HJKB/ySHiIYfARe586+1fYW1Ti5FbbSStKIfBGb9Dax
VXRVPmJKK65CM8TwlBazS9EAF+U/3ANMfa6tpBC5czfb4gmHE5CPAZ/ZZXcyTytysYOMpYA+vW/T
zUeGvdZv5rhTD5kHxEb67ddECAFUP+7tndWx7OXK71WKwJyRR6xOUhbvIfZyteuSeAzEMWzWf/Mj
64JVa4ctfNlrtG4FqSAEvpd5TAbGVDdC3/DoVsTq7khXTU9jC/MAWtxouSEh9uIZ4lFpPT5LgE8j
yVebUUeOx6GF+uHKFJFm60dd8wHEjpS+OXHZfxJ16r2Z6RA+7Qkg9NhqqWfC5R/8FEfvPz6aFOLb
x7od+lU47XtmisUu6u4nCmFt88DEFAqqsaFeAuQefr1wMJQc8fpLdtl7p+IG3hlWo0vYVj9yF86+
YBZS6a4XPL5kgjd+wT/CKrlJYN0nzQjbKxl8wIjy8QgETup5e1xBCz9zywO0tru4246c9wcr8fbX
zo8ugTExTdtq4r08c6ieRqBIcmYWSe4xXnftuHAT8XJRU6LJ4acxs9WQsnoz/33WAVFNbN8UsaaN
t6gyyUQtd79LhX2z5bPYftBaqRxvWia4axt5Y8Eg3/wid8JyCWuIVISSuankMQ1ncw5U/ESd7+IK
7VNTFIn0rmDF3WZB/4Watny9pQHZFbOZ0dcA/Ug74y6KSo65roB9w/Rvb17pF9RbnVa0/rJ7Vt0C
h9ZJhVs7zX38xA1jKn6kVBealPTLFtXY2T1VCSZr0PYoO5JQmv9dO0Ks7Mw2kd5fsmBHd2bqwQSx
vpYD7NB+jkqobmprLyg67yijkW5A+30N6TuvHAd9n8u3CA5oTciPS0YhZp7j/Wz1kpk87HjxOWke
uoD7TpuQGmwEb0ZszUNiCwfyuonvGV4Bcushifz9WSZk/2F65jnZuARgogzw4yKH0FIDz8W6f9sL
wb0kH6kG8JS7hKw8zaDBh1qBk8Xz+t4yPRtl5g0ymOxIP0XszebTnpqnGDkiDmgnAdkUApkPmhu/
bfmdLuozOkw0w9TzQ1MQHdwAguaeUvAb9t2Fi336hBayVLiD6aAKbX5Q8BSzbXPT6cpO38xW0xOA
mTPisfFwE5XhuP/tGYjqgLxnebnfPhqdLs54CL3MClHPUtqkwviHxFs2O/LhxC42dHvyVWvam2uA
xGZNf/Ecx+PJ98QQfmEOogQKZppSpktJlwY6bVJLY+uJimL2J9/pn0xPLU/xgnDz712WfExd+qEN
41ytUo0PpSvZLNrf3c2JNsg9R936wV6rf1GhYsj8cBsGyuqOFOepM+TLsOwWYDXkTZYrl0oqw19U
NaLzGD2o8LuGamYQmUOgD6uOoutZKudHBed+Y2zjrUa4wZYIe+fMZPR3r0H5q2uF8UMayKF8Kon2
4WfVUPixVVOIK+hpYh8tIxUwdLnQlzsTXLHgE1yxF7b3YdBvBu2RzTN6ijS+TtM8mmJTgINOjqYy
bkLnMA+QLZDEzBtuhC0PQ5FZYq5Q0DWiEbjTjJYjOqvqKS1ZI+XXfIIL25kDx2jHIy4aEZPkSnzS
iknRjiWKR1VJEVY1/zdKuBI7ITA6GvH7Ymq9iTxnYfZAyy12Nu17E9HV9Oc980JnZVjih2G8WBOL
PfRku9XnincyD1UHBE/9+d2LGdzpLbHd2XXYvxWwtEcGGIfWlun3HtYf32l6FPN4eXo1Vf5bZ1FB
hZS/+EuErBXJ2NA2TIpx3eVx8fDzGt/GCivRPtdg0vO0PoFFhTu1JpHDBNMgb5ENo41NywgsuHUB
EnLK3AQyMLGVlg7+hy0sDEWIOAfH6gNwT3Leb0lqPhZjE3BlL2vTeG7oYxYG7AWKzAxmw9WkIzya
GZMIF4IehHEee+bmzgP6K5yY8hb8MKqLgnTfNnVSOHa4Alv8oRHKoEKamccX8NtjLpsLhP+oFbTj
fA6ULuKtkDWVkKwIQz/0eLYOCe3DWqtVO93co5cTq2EIdKaDcLNPfYvx2G/WvtNk4+Bmkc0R1/f2
QoVsOsg/FJXOW1PW8ZElpwWehgJpmdbxbafRLh5prwxV/N6tpsAs543uI8+Gnj91VjNkLTH7nOBS
arGxWmEtuw4LUCcoEXEw+CnN6JW81u4mSnxSUE3+okfSm6ox8LOgL4SYc6til/D0AfJO7DNSUqsd
WxWOBKg3ruxjC3gjCwWg1KKbKxH0vTkE7esG37Z86fJeaPgaJtwosCC1rQTjtf6cHzi80ZdcDDRi
Fyyhz73464PN6jTGN5I6hWYASyoRv+qmsaQ+CeIUogYi0qHl5Q/7la0aKh8HXjwv48RrpnZJzfDJ
ULYZGGKJvsuPdIXKDgDvmUm85K8NTdNbzDPodERbaTMNKMstcHfT6gsLzYPl2D5hZkvh6rkmWXat
VJNYrb722QmpC8ZNc+uYJa86FVZNh5O/KQkd1wI/gZBlVHazjcs8JfRfmNea9pd+ksdnbPyzGOg3
QKFU6xbdzLh3tt6VB/wMoKHHoJjZuc4ejTBJvKaXXkTOZqWw4Stbaii2d0e8/q8BCGVnkdg/UIlR
p6oxAHtoRJmnFuJV4dy5UCIvO+PfmUgMXzzG9oX91Tu8sLxvKgz9WTvPP9MBidpspoNu1yZEHbF7
Qm63nRT8TeFMQkwvKM//njylR9U5BlTnGkavbwMEhgJS8KAT4Roty1CtX+cmmFJhrMmfeB17PhOR
l9PFXCy21akQQ0Ab344hh/Zx/j4Z8+J9qTOURcfRmdhQuNah2gch5Oslx7q5pKWBi+WyL/TwqjcO
vcoRUin7h4HggXMRVrUZk1eGErEStTzajxanPTZJUsVOtSGAPLH3KzmZ60FMAHKsGB9IfLN3tYLm
NzbTkc7yVcIWlSofiiUnJ0b6okLdo1+ch9qMEzWM9wu+egnCFFvc8MtXD13mUoXo/DbCpyoYxqGs
K8JN94xiEmyxORC8GYu00h40i2gXQ2Nw/lSkJ93h+tKmrK2PhD44MP+DFKhAUqQI5W9oQ1jiXzsh
0dR1uzVa+ITvJbZO1B9W2Z4dAaQG24k+XsXisPznNpwncCQjedbcs+vQALYumaoiNH0uqze1RG7N
AIBD5EUDnI2xV3Kb9Xbge7eij+ZOUXFCbjO+9VEHN3+G7Ay0humcauNQRCFVvlgq7P+ucHYOiCbg
Hlmyh8uyn6NB+ItZ1DQ2oAxY7tm4qDTif2QpwIcKlxyekhia+h7FAITOk7ZN3GelRTuFObQO7pV7
Z+lPdCYkL0AFKiP+LnN5dcC943/eJAuFR45vko5oPnceOI4fNKkAluZ2ZmNtk9fCImaRDNUhQbhk
MvoKLBUUuCWCANVI6+GCTztkT7IkuZGJaomuciTmsxl+pES4EZrECJ0jdsQIDjlI31sxfuSlQzw8
5XLtRqXBZOix10fUyWOsRRXxyUWtuFhcaRTrwjXmJVLFOzhuTi37G+UaqfWbqw81kfG1bJCAqwSF
zEoQxv1e0DEXMAR7fz1mmBcxItm/OB+/wB3hyqTeu7pbG4d+PRRyudsfB61HEM3ZiEzYBeSTmhWq
syh4WYQ0audfhBY2Tykn9qpMHMHhUYVYunn5LNEwyiNvx9+H+C22SBHfTPnaV7b5J+KUwIwNK84g
60b8z156Thoe+m2BfPhdQOC++uCylN939YeFQixPVMYswabMaubYWO8mHOSRkAKCTFBkSK3Gzqy+
EafQe1RgFXgBVogKS0Os1S+kptGKvXdiYpAshKwZC4rxlvF9U4+5IfqxWBGmqvlbdXy/vFnBN7Bq
jBdSerngcHEYnSi37bEkCMCsncExzmpnaQhBUg7lnWv4bP2Ut4lRjMLp5+RHgqoJTcs3eITiaHWM
puI88zHIsHLYLs+RXeMnWABjTUsQSPONTEO2wt2ICo47J6YOW2ouRQuGvOHvrvgxvKdhQfknpUeK
z5GATiy78Ho7F5jz/85g4tSk70aOO8yo5BnlD47pz+2VbcLXPIVuHpxdU+IxNdW7frPGIM1X47St
Kg7TYDg6zuKQlGvUjyzZAdGvXF0akzB9lqpTmPsgkgG/9OrqwDD8xlSfy6HspmInwUee2ACwjm+d
w5ZyAvd1amAk3OKbhBPrqXhuPTLjcGvHZhbKY67ZW7mf+COAfrLlYUQoz4hUPsWBNXRUwFlFM7Oy
LCv0WGKyhS34IrhdEiEB6A3b1/2Gx0wz9c5lU+kXH40jogTpTK1qnXnSbDE2f/qRyadU76qkdrXp
E5u/OSqhb726JGSND+9EZc9t+3beUAYCX5/Jtu8xhIhWKQAeoYzuYfU2nPTuVR6+nVmoHr+VpInq
q+zLKc2+tepp0C0ZKnKnsZthgIZSm+BwphMYJkBA9HfKWnNd6nifUA3QC4yLqfLT8mFZ2ylhpYoM
nm1Ao4hwe5A6fxZgc6w/iAgbh7IBdTz85Caj+o1eLqEAhHDs6/xF8fALmLFSJDqPFRe99FuGXCa9
cHGvaodj/iL0kTgsx9Uzlw6Jy+OTNKAHLgnZ6e1F8wDSGMnjDe3/2F5WZ+UuIl6O0Uj7Vdqdk7kv
UZsyRDa+jdy4i32yISetFVBo2IvmQAL03kRlaBZh1vUOYKveHWCVyFM60/38OCf7F4T3hfFOROeP
kWaTBstZuUJb2JWm33D1VfghJ2Kuwsr/e9OgItl15q1zdf0wMp2uV3tWa95dH3QPXvEwaO2/M9P3
1l4XKSp/7K/WEpFDBfMqXPj0coPub5E2odef8BzNRtK+1RAYjjIoMnPV2Qwf+uA4lyogD4DewHbk
JkITAPo7g8YvBWuv/Zdk+EskzKWqfuXFabPXHqIyzWBS6YymQira7E+JCSpD3IbaFsTWJOnInmvW
scBuUBYSrp6ZrSv8iAcNrXPzxAwYxpYc6Zn8fAsBXwHECzpA5wOdbVMhi06StsC7/YSBcPK71yyg
Lchp7t8SW31wdONuIRHruGwkDVe/zM00qK4uDYagZUz7hYv7jGjxScoJrU0B8tnLkREtm+IRfHr5
+VdRzNtc8Z65fhhV9Cx2hIr1qryRKTSMN4WLXR757QZ1H3fSOzNTaGvylFHICeprxhDI3ZuUWAJf
WRu5RBopolliERpCvAL/5r5AnLOODGP43iYDbGgrASML/lIQID4+Ra9ZVnfAtM4BNmjZPxzth/mW
+zmjmLE/ol6VDu0qzEDL/e+3xef/iUZaLBA8r3ruJI9FEUMNQzRQ9yeQk2NXhT5TVYY4UsZzVcWW
e3a0bli/BCqG3EDFeYWyFhH9qhb4RtJV59UkpoPHzHKcpK4IKktQLrNZ/APkVjrDs5ansQhDfTSI
VnuNAi3qdzGAfK4tLBvTKzRscJ9GojKkJF3femw+xrajSmU8I0/VNYGwhIf7iN3wvXze655SxFnb
gN78/88DUc6jDNtLeevVmn4QASvMWfxw1wV92w2LnpqEg1Fl4cAY2Qx0ecOI58to64pHuhWBynme
IthbR6J1hExi2y+tvjFN4u4rxTbuIk/IYhS6NF0ieKRChO99nmtE2NovFe3o6khnCosgBCiRxQPl
L+0+SqzKeEOaLHE4qX8/U0M/ctjEFV0o/Y1ogIx2qkVsSObzJ/OQRvR8h+DoCPdwOLvNMV/L98dY
Ae60Ni617BzeSiRM9bYj+kGSmtxZ3O7sez9MhZZTCYktAVcBntA7qN8uQ7Eo/wffAvgEZ/YZZPrQ
kkTL7EGtjhfHxRaq20rZlZ7QGaNvBQNAlyCIgfWB3R3+2kuz5Cn1BmSwDCXqwQbGz4uILqEgI6VZ
MUwjPhK87/dRLQbZkztBOIAfNge7c+64ns1Aind4OjTzuUio5P7bgrVCeeglPfzu2ootktfAsDdv
V3Y+ldmDcFg0/wF3dAMRciqIzKkSG6vVN5yURDNcwIk1biGypSzaZCL9ZwoBY0NnbsTpZ63ADTXl
nWPHQqp27jE7Bh55g3qAjCLjWbQSsEGA06SDKDR2PvQTxsyex7PFM/t1EL8AFY8SPU4YHiicfBl1
FvMZ8FNVnwWSBVTuImagAZcrcPk/GOO7Rqf4B+2wI9XMaTLlnQ8xve3KGQRGggywEOEZePNFGej/
EcJUpOqex+K2F7zpF6PI/3r4FMJLKmOGJScO3jIOcUvoEnACBcFl8WkhXIX1oYAYC/NsLe67FH9j
NDq7hJML8BRlHkr6RB5pAxP7oNFqi94ZBrRNethrIdvkrYJRxdkJuF0Td4hWt+5qYzko2eI91D0F
9cRuRtu1V7vroWDQfImXXGIV/iD6GuD5/yAfwYRZHzniNx1bDbewnOjFIItQ6Fvub+q2d5u4PvCD
Ke21+KTJPXYvtOUACzqoJ56hQsdrptfvyT8W6oPZvMXO2jYbg/qmA7DoAglZRJWAh7GPSPbbH3Q2
47dV8wTBCdtMzgJOc31DGMyK8Rir0iAWleRGbnhctTXii57cByNpMJ0+nh7lJO8NPYB62eFXbB3c
j9kNBzojzH8hREnblj52ZUOtpA44B0DWQSQ9Qwb1KjnEajeZQsEA71oC44OBrT/TyD0RDZDnj9Ju
6hyFcMrcIJkSBR4Ttcr13g/ATRgTtWN30n7qFkBHcfGDcP9Kc0oHKbx9KnystE49nSFnQLknvvmq
m/Zn7Oj8WgGwldRWke7Y2JMGUevxk7eRLs8fN+eP7HPmOtQfHOXBraVBCkJ5hP2B+w7OSfoG8h2A
+yqKDnXDNC4xp34EEYj+ugw27edqd7sBg2zH2hgBBm5V+oea09VTBPFBMveIV40TmuPN4omO+568
bQMGSBGO6qNd1N3RVrF+g5b/hUdUprewPsxJueNNgrLjJRIBzJk/zvQrKmIt13RJA16PFTMLB5Tm
0K+4opca4Gy7kmqt3lwbLYpZuiDkN2ldYIEoZ5YK4tEiej+Z59gpaMDCja497P3yDyELAFRGdCAR
GUXPU3JDskdIMhsvgztr6xMxLP/EyUZYFFv2egjcJT3dPu+u7dSytBSfiq0YGq9f+mfN9QFW7b8C
jrxfCvRChvAhMJcPqxHE1Gy+vhipB4j8pznbvaH1SYEI8JkcO4Q7m+SJc4/nfIgnxYDqrI4yZrlR
dBppvhv6obSHj0ml96orK3/kbmTJ2W8RLm80hUS7D8JVl1JirfR2intRiCPg1MaCFPGlrYcntnOu
gRwW2ilMxSq2yQtW/URTtnV02BBAJrWqxqlqpbhzqfUBVyCjRECUbO7grY2UvCvDvH/F4UEtTyht
yM88MbMsXhRpz9ezePa7VjGwyDrIivKLX+BZdc+K1/RgJcib2KxRW1lVO/UsCOYtxxlopAxNF8dF
96FH65VG+iHVxwAF0No2W24YPAh9fYpauEhSSv+fAybSmQjyTqc6iedWpr2GL+H6hUDTqcil+pqw
fNpozojc/VGRQrwDcHbr3tPJUgU8ieesmaWuPgpxP+mD+GrglGZPRTgyOg81uCW7lvGzuuCDnpka
xzL/bUSfGrwNbYkx6eCShYLdhXvlycMAlimkGIokhnKY1xU1tfGp88DNqDswHWCT28cEU8SfYiyz
dSAc03JixYPv1Nd+rt84Q2VXHxDREtRa41HagFxFDo95PVKpP5Qb9GmD+4DVyTag/nmzcZOxmnzl
3t8So3KXSo4qStOuBHcf+gNUUM4ItmhydNxi255BW12T+OSBrAvOK+UiuGkZP9bbcIoCMRwl6oJB
P5Du1nr1aG9u4fguFh1tecAvx3BLin4S3OcsiLyGnD16Z7tYr+SKcJyiU5NPPr4U9M3GEJNAsHi4
9Lnno9WDysdEXGgF6MyrBWfsEqusmePg7gy7vQcyu9BNAohQopBTGjvJeIz8gytp/pAvKXau4aSB
Mv8t+pzGg9+qubSqoRa0LSRurFR0NjHgmIKlzK1NpwY94VZ7znez8jXmyB3/VLwCIDwSB+pcP6GY
xCsstlwKK0QaR6ttr7N6+Mmolkr3EskRGUlw5fhYzN6f4SRcJL25Q1lAZFAlGjUxRlprXFRbXXA4
5lGxaUyCvcCG34YxC/R2sXcHW4Gy57Z6Q/tqcPRvsIrL22RCptOgPluHkQcj931W/8mchdxWX5Hi
9cvMdv1edmA93pjXxLGQt9CLFRaUXQST05eSBe2Wm9XNqcjZMggRJpp/YwOXJoMlcehGFZvV1ThZ
jaLZZ6lTgSAHryDY1vNPufoxinvb4qp7WzZqXiEwcA+vLbJFjUTV4szja6q3Lvk4nQdVNUyuVxdn
Dx4dHf4t2KA9Kb6yEukpVwgw0rHqlKUfq1iP9tXJU1YLjHqjIuOqQGxXi+zs4feq4uJtockArJpv
xexNFoa0DHzGScVkvM3qgiLZgymJccrlqATHnOaTB/iuSfleN1nzpJTaG/o4fQoeOGSzOiwzyG/J
dE8HMuhkbl1bCJBl0qw3n5nMMIf7CPJs0zQvtxUnJGO2iBcXlg9U1HJ3NbLEtW7QNSholG44EYA+
ok6TzblzbBCne6MJnWRNYERr5KJqAXiIY4QRRgrpsga3zckLMZfuMQ0udQnA/nc47dAWeveJi/GN
s3R6ZpG7LzpxN4zlo3jutQuI1UFiIH3opRndUoyE8HJJqT/BrWu2Sl2YV1FmNA6HvNBt/ZIp0TWg
uLb6B526nA+DYPXRSi9ZEz4x8EXIXmuq4CpDbNtoPoU4J/cpYI2M5IR0tlP4Wn5qA7u32whNK66b
SIcfIbvvIRxRebQ6sgAJU91F/waTaMU0h1yjx7T1zcX1icWILn5HldikUtEDWpCS58upbqNkM4Ne
DJPwRp2KMVBZkDTfiYdpmogX6bduNjkYts1k/QQq3LUlJ6PGQFgANj5llFfOuxgeOdfw0aSlDx0y
I1g7kD1gJIIlm3IDujRzNzjDBglh8TiGWzyIGzlIfmeZi2mqhyOQQOVyd9+bDLCUuNJX7G3XRZJn
b5znA0SMVhunATaFJUujatdu349kgLNKhZcS68p61JFjNzpiEXnPNAIZ1dRm5PX1mLRPqntvNChg
ZbRj5hM9gA9djxAGKMezLIU9gtGK47Qa3a35X8WYajqRTzT6h2OYzPjDvkfkrrUvmmy/g6gl2KC5
yWgoXPviH7XkAxfOKVxArFr9qc1NOpeP+32You65sbsxaW0I8g87nKT6Zi3PzWodTAQi5DpUf6eT
IuWYNjwukjinjVBl5AxVKurWizwWgXtOQ7Wp0lI6VEcJk6ar2bW0lWjmpqekPfGhu+VjDQcnZqq7
bT/8tExkY3x9y+wkIHjsUdkdJDw65OkbTFOqx7CGMTr/yDvtcLU1t11sbpt1rDFaKIDVrrggcTtv
rLlP7zTTwZGkJg90ouDQckjdVgcZBqFrtrxGUwn4/uy+CIQ99eDQuZXvJiUKjOXw44lEMv/JnWXj
JTvlR/ytzeehegtQgdKhp93QZRCYI3unQSBJHMHXImrDFKYvhTCk/WgvXzTxGz8U9rbVfqBB9n/D
WWYRU/IWBRtiBJX6Mkc94AzMFznhspueX1h2EoFBf+mVKXy6gvKttWhBAEDC0aaJ0JcRoLbicZta
+Vmi2Qd0bNQNmoxLs9g+Hb/OQQ8C0BRd2V228KmkA9QYXwkHpKvVbNdizTGYkXjxlWTZPhq6B4he
KGd6NIBXQFj5nIv79JxHclD7xUmyYlbfnfJMv6ebLEbs5CvQbGq3Li1b1w0NtV6xcKkSxgusWmEx
mtcRvg6K7GifS/eGeUjkC+yeo8YArEYiNBqcHAoLbKo6pTDR/xqSluBKau2SR+q8EEOm9AJULiJs
uegm7XeK/ImvmBp38Gz1W1Hcmzieb8Qczm2APEPKcmWO/93FN3jPjzKeNHh12r/2cKO4SXtg8Xb7
SZ+N/Fjgp0eS0cfnKlFdIRJZMTLzrfhy9MYo7GrrFvVIEJ03kPLoaEYFNa93LopJFBRIugWvTMrJ
QgbE9CrgqF2CNLOPNGw4crND4mlJjQTqTY0HpG2+9S8DS+vs2BMbhbo+necsOklc2K8aUde3lGjk
M5JBzkk+AzBsWkKIT+KFiYx4ye9GPIDn3HphKTaFAyyiHXgGBqq2MehiKmqp9Rj3mqgL8ZtuUSRU
zen7cFFiHUrd1AuhmfOQTXusj3yboYMaO9yGitGOR0SWIkrqj8/s48QeypAUjoNu8peHzcbVBAoM
B1jRHT3rBcKlJ0KxISHvgn3KI95tjyCnfgj4YaVFHqMp2fD9vHXa7zA2wdFpWUzhLHBcPmjDhqj0
fpN+mqn3VOJ431GINbC2UCgAbQMvgdiM9cK4ujzQ9yRak1ObIRG5SM5Cq5C+5tb3xuVs1PLFjTL8
eLhX1gYCvkoc/htXyhbOCOFmWIY/Tkim9woiPry1NQncy11vInKhQtRFBzXVinQPk3s6oR/YmJVB
3Cw2ZwJllIEfH/z7L8tPR3PZy6PBnFSOhi9DMa1RbC8NWakRelcgHyvfASea9XuMocEt+oJm/rjk
RBjkDCn7saI6WkvCUoNsONOLJBZpTRP8j9UwwGmQGEybz7K7aWAIaY24u5wYwlZYQxbDs9J3U0kB
XC2WuosTrvuqOGCHW/Ah3f4/PwHJBPtQpG+CTdMZ9letpD7V63XEtITKBh2C3cGxA8FphlXjIiOa
TB2lDOU8F++2rcyeKqEzOmT2VxUmBvKe6jyV0xSbjf+1tGLBgssvHj+WWjgQUeHc2ozc7CBclVmy
00ehBRF9ZlLSfEE77XVRkghhutPSPL0z51LZKVmbyt1wVxrR2bkhnkFIVBhyoMuYBJnH/4M7oVpT
YZ+szc38zH6dRUElkTIOgV24jkBBpXbJXkthvImvDGKwgn2deVvKzaNZfXic0hZga0Dpw+jbQQVU
raNAeme9IJO9/lVvxFuvRnACPe7KoJjUccLJNHu6K9Wsb2ZkYfDnQCHNT6l7P4MFML/kADcyCfzh
PtOEtWWePtuaEZvvEx+kgyBm/LxLtaF9IjBgVclQMNG5nS+OfD+uM1BJ5awIjyWt+cFtD13JPvuG
QAYkyYy2zZNOviSvEinDp6hG5DN6Il0C0BQDNtdUzOBMCmH8oV2d/0UCKIzdk7MH9wdL+10lg5WV
n4TpZhizJdYJeUJZrsjrgrBuQWZmJjWQaDOQL0xMhgrQWVGSJX5SZA7C4207s2ynaZk+4JcE/bXV
yfCYv6DnIcWANKew8W/6DFLPFWWMC77K+OnAcO2xK2zZPBvzAD/vWPCxIlfnj+ydQfsDLECFkwiQ
MmBfATTQiZuh065j/ScQWYdmYlqlsYOV6diwFSL+PhD6ViFRLQV7lpvW1bKJSegvGUnU4pQBbBW1
gqtkO/Vgx9OCeN+d9mUKAzkJS6W38e159EgejCo1eNB7matL79ZWhPszAyZEkSVwbUHPtSbBaAiL
tK6KlqcqNhkxOt6lux2iPuaJCtypL4XlMParjnFY9DueN9TZ9yildNFPm2m6QFsKDLhn5gyhGMD1
jSR9V4o3jyYrfB/rlqu4Srz2ZJUZCnDLDTW75NGL4ZYu4ax6b0D2C6MG57RITciAuuQK9maChRSp
MNHZUdAuvgBDROxXzpA/90Yw0FYm7niGIdm1gQLliYnqob1hUivq7eRVP5JYGRt9yQ+a8jQUhe2l
B+R/T9Ow9D6k5en8Tb5eNQ4oRtB19Zz5zYUo/rRh1nZHTY0hD92GAx8opi5SvgwxTHpfSr+CqXEO
35RbFKaNJPmoYCVK3mzzakwogb4ZtOGdsN8XGpvhzNWWOtS7YolFzWF9vR2PuC9e+5swIO0Mtpop
QQygX2IiCi3AmIgKbdGnAnkqbJJMHFzV3w8HWu6Q6gC6f12ohZveaCu3F8RNK6mmGP7bDcn2a+0c
zhnFTAxDrPwb/sK5sc5sE78di7LaZhuljUyiZUpsXD7/X1lPnFrvfpu9A6BcujtVUh6KJR+gYUbT
bzCI9G/CFA85gc6H93Ka6abe5hJPlB/sgU3aEZOjAu0enZqWxRG13GjuSgvp/lVvDgcqMCmcxL9E
hqC4ZbpCd8PVPz/ECuU7vruMdnVsQEAZSBt1vQhOD7NxaNu84cbobGUPw+rTI+h4DXzpGnQom2F3
1F7OuXLzWFujLA6P13efVvA1PVHueGCIYuXcm3a2FHmWAWGsNks9ogPfmohxjZRSDfjF1DBzJBWb
qOHVk0HeUd6IWdSqBYe0yQ9NSaQ7MfrkgkxEjt1IlXfQCS4bdR0a+mQu9scnlhoLMNAHL4jJCEU7
sQryC3WhTbUzf2lGMpvUapcB5mIasOA3FjiabHMYEYn4Kq6JR4au+7+23OTAkv+7PZScGLW6MTZB
SToAkfhIw9l+P2jjFvfmu0kcCfbHsy9FlvexUyupQWUIYKQD7RyXm+N91iGCyee+K9cGYIu+9wAo
rbh9k13ZOnJjAlRaT1oFftrvpB7oJjWPcuj9sK3oDKqL+ADvQD9sO1A3aZ7DbYSAlX9yDIgC/Rds
T3q09t16s0e5CCK7Uq4rFdqd/j8LrVtJ961ohi03bXBhCz9cSUmSD/l0RioJAmTCTfQA1XQTwmZv
C/Oa9f+jBL8lHo5hpyoUN6s2pD00jbRrPYyY5BEC8PRxVf9KcvG/uQUx9PUDMm4UgVbOOzwTtNJq
gWj1YBX0gyQJTeky4ntnYg58dNblI+ABqk8TSGpCEeSjNi6Hw8Pm4qpnEbNbMojadOs1/7a0d3js
hv1ZOYHFVBxiOoqxtp0ZqPs7qkB1/bNWxkx6TM7GxiAe86oH1nlziOax6LKDU9KjgLdNOTVPzzBL
7dxspFvDxnvCMR9wRqpumYgMUImjoha0yfNfaOAdbD0S2Hz5kKZwgNHFEIP3FvztVqsamTH7Y10w
se4SCQwqtQFGisj2PrHotCjyTU+mSnJHXOQvvJ3u7GCgfDYSubWDn8M8c7GwkCLg5Qmicd3htHxt
veuOOpDDfxL9k/2jYPiqzM3qYG9G4hX4nnSZJ/oJIQ7BPzW3Oo9QcLV70n7X92CbmAd23CGKvN2T
BiyYC37u9M28R8Bxx5+BoIfN8bU7x8Y84xI+HVkSU/HDuH8KjtUpmU5EZpvtwa05CEituKmaClsq
Co5vQTTfWNO1ElbPik2Tb6+zLckeHBaBZgyLhSTWGmhThZktT4ccfnX4sk9fc/7dapCRUQbvDUsp
6IQtZog0ibGnhDWBfWQcrH0HBAykDdXxtmw+QXwBfaORI5FxsaX5jV+I/PRRXNvnzicmlD/gY73c
oFl5dNSCgl4lYcz4lK+65QYeVwxD7ZJGpAGy0dQWoBDuJDVJL/OohVUMVOrrM3GkfQXv8zxLBgMq
019C7tPQiPpT+zfbDRhhQ9jUe62Y9GKc3UyBskd+jJoQ+c04vpjgnvUrCffBP7BbfBdzowEUJOFA
cY2mrwo5iEM5ItfecKOSd5ndlimc2wNWa4vwamD52SG8qyFv//0PJUEGTLzZRdOZ9gWDWgT+ha7d
pwNzJNdMgsNQMFC+WlRDv8qh9iZLsOnQD02b+wI5o50I5x+V96TWqSL8oAzNBAXmJrxDFmZ9ZXUQ
R4ZhbD3VkhqRBrurb/CdOV5eiXT1pTVcM6YfIXrs6PDKqU3Cz39WbTO8fQNKR/k7Xz76ER7ApfCP
a1vFFAXqw3boqThuG9dcpAH9tAX7UuPLu2312BrvnS3WsMoK5yLol/MnG8CsH5B77ddHl0puT+z0
76jb/yA44a9FzKhxUvRec6mHbQfNU9R1Epe6BADX3GlhpDIva8+dlDifleKFHgsZR1lJDnW9NVdA
cIVKvrLOhUL94ubMylZRCWZ6pWjynqqbZdCRjV4DezLMhboHNvCpkO4MGEtFG8xm6i0Yo543yAs8
JtX+0FT7dpIjX/VIiSlFcBYi3/msfs/kNFGbKTXAadO2lAA0VwG642M8wQiNYjHu1qCtLa4Ml4ae
0MiNkjw1ahwLlbpkJ9GTFlONLjN1VRzh0HrhUsoHLRZQ+JZyNbY8R+PXFpCLk2u0My5x3q6jjSOe
JC31j80NO+6582dtnzZ2QiFdKSgI+OZ1ZuJl6gbrMalTwMjisFr3Wk4+ZzaYBRbfB6VexBWDdu35
inPsNz6ELE0tul6UZdH0ISzfDE7tcHq9oZ0pdUn+cC3dQiiqjvjFFFQg0cYcv/gplZRxO8u2b495
WfrP80wqzb+gedXMlT3DSk6Vq6yeU5H06pH4PmV+Rw4i28N9pgr0R4qdkUZxei38b7l5v5xqzVsu
RU2IejeRVNAYOmjKgAtSlOblSU29VU6BA1OsEFg/zJsbKH1eyfTZ3FjUnLiKVoJJ7vo3ek4+9VWB
jdofM0bmxd0EqnHgUkqTAO/YONpgXGQFFg6smMQ3jW+BQNkeXuu35XPFZwg1dtG9yMe/ShWjM8Xz
NO2KSET8I92K4nUDrBHLbHVOCEmC6kLWP2iwXFKL96UjxohTwGqgLyAhkZq1BHiPf28i2bCBqgGg
vnT69Rli+RBagHOQJ7k1MeUyNPDnDoRGLpe581h4hGXoxL+UbOIoF3SHMKiUzXv2S97oXSCf5fMu
Uz+yFr2KQYUD8wS1feZJ4FKsGteGrC6RFtb0YDHW8pXS9g45EHYAB5+F3uFfAwnJeHXfSdXyAqWU
zBLtW+J0sQ0q1zov5ogKHqDPgEWW3BY2Dp0CAJiOiPSFLIPPmnak5i8Hbj4wrFMncRKsdE8h/bmO
KEj2Lmc6nOChSXGC5iHGijwiEvYQDclaoMrykQN0JIi1G16ztoaWS1OJZln5xivAeRIUueE/GZCe
t6t9FLhRFSyQ3luSLWoIA3HPMjMR+rAgCTpXzTsKaPWoxSmirtmronLxVZW8/IhOSL6XdVENDEZB
yM+B4mrZhZ3173prxN+6k4QUUPOSj+kjlA7w1cavRad6q3fQ0CpsXdps1YTm8t5hJlLcWaqm4lLm
wir4A910KyS9e83UFLs8YzTnztMoQFT5Zwp/kzp6MvUjg08enWti7nhePW6sGl0jUc0puf/rB0YT
N3WarxorEZ9zDU1ZszqnTHP4fXbVr0tYrS0erU0Q22h4nMJdEtiZZvXHkorKSNSqTWcgyWvLMclt
/1KKWKQQ/awLF99FG3z3Kbjn2mCkV8xc4WCQjq08IXB1lchC+VGZtIIit8BiEAx/DCZydYcjVI2J
Zta3+gV+UaM2zGRTKQB/8L9z8xhN48D+1Vkkw69RneovrgICxWAdGzSN4VTZvn/BdHsvynupsQbx
OP28iMxR1Fk1h+44r0OyKzmQHWaZIPQZJUI2fJXd2b00A9jbsvf8WsKLf4QnAcdRjOhaP0INw/OE
yMtCPh2+DvJAsIbuEP9ieRt7XyMSzMFnBCzCJjzKlEIIR2g9DnuNFbzJBkUrdB3WinQatE3DYA4k
yIi6EYd1BgKSDfkNBHeex588KoD17SWGN3CxcVBtI+dskjrbGHSwHSox9+8EduOnS1FNfPKp4Sw7
oCsh7v0i8nV5CQ5EahMo0HyLB34my82pYQ+8swwsBkWiRHf3tD1cbGCA+v2tRzHpg7Ker9HDFjYy
8NoBjBLATl9vdZ4PmwItzmmyepIpzQmsB+WkWni+ZECDtRojsv7dA/Tyq/FPeJFYDThB+QKV6EFF
D3XOyW6T70vQeFn5eOoYptWh/iujnVf+qTHNMyPe8F9yUUe1mF27wfTct4bQ4qWhcYx5Ux6yOgwb
2gxv5jgum+8kJlCFcwWHAA7o8+ZoA/j0F0xwLnXv4mhKW6YzlyUYSabPu1llW7Sg5eYORLBSV7Zr
URINPpcWqF806ZgTg4PF8zau2Y41SE4QEEdZzVfQuD/i+fnBlRHGob1xqco0F1J4GY2czLSUZxgW
q9QmqT62vLuqVmqadjqZgw+n/r30SKgWnsq+bVSiPAp3QaSxO5KATvu8Zqnq6LLkM1Ro3cGbP5Wv
Z0YZrefntEc1+KQd0aYeGyFi9J7RSWJol3c+2duzJc9tKkMDbL5KMq8GSq1YV5mIAkBz0bJEnrQN
bxJikKLpFiIKKGQRzdxQwfKdCzgsLZN0gG8VMacmUosY35bmKiYRkcl5jEiq3CtlOOUjWfLQ8miU
RHkgfH4IJUXzE5UdQImAx6tzqGa+GGoBA9bT+5SBqHhoOL28JSBS79a6m0ycvW5UO166X6i0YbTb
AkvpHZsLQfvvPFZ7xwHA+xmysW3Jcv+ZuKMMK67GfgwGWfTg6MSnW26i5xdNPmyCfuMRGYnwiFYV
kXIerZtr+S0sL3Yp3+uFsPCcMKp+Gsa3WO8C79kf1QCNjlcVehDxPycXiK77R+sTm6XHoh8QaxNc
T0f6VX/6yvtNrpeW0QtF6JKmKWjt708it6MXlj3CDCqd4RYDEAcJrE+6LQBLwdz3c1E0CqH+pmgq
r6D5JKMzFr+GJyy/AtXyptSIaWVdT9kHZ2ysKADN+VPB58gCIo9me6M3EkvIIXjcs3E9p2vjhky1
28JHTlLcIWINECMjvfbCwju+RTajQVSwRcpVjAR3IgsxFwgd1JMQcJ7VJuXeS2nihxa1CMLf6dbI
5YvrE9vlStbKX24Ugzl/L5B/FpQjaGr365lxPzreTITUCa/XSvtrnvo9P6eHty21EnO1k87phqCz
2K4VL6ZssyMwFLT2o84/LVMRbqug0t3wP6vKVBeiwvsx+3DNBlXmr8woQc+kIRdrDrj9RNSPAoze
Vu+iy5nbEdSHdlIPom0fPcXDHeK7TJ1IR/uz6rOjbxF+JUoBYpRgbE/V2wXMcBVDDEYjyb7lJJCj
qy2kR9jKn1NgyUQz8fj/zeH/2BrX7+HKEhdlDIoEoavdhxhqLN7ZCRX4NjQdHg/keZ77NGncCDEO
xFObnLhzC4mvcmRJgXd97oAXDvveRK/by7HSO9SFU2qSuYZ8a4X6qyBC1XhAvlMXrhAuKjnNufde
kJQKCx+PyB6VuI2mo4RJctn5x44ve+dAXMlcQxROecQX8kWtb7tp+JzLN4JZu5XLUd/j+lxybztU
pVWkghiYeccENBWpB0y2ip0ljpw9OVvOlAODt82qE46UztLQR9gtwYxYC6/eVYRDR0bb2+NkYHnq
Md7b84mVFamSrswpEJHmipjGJ4UPXl+kw9e6P2XJCHi1iyKUERZ96xk5RTW/uFoi7dyrdZ4fbnO9
+INWxHaR9EP/YUGyqQMBhmF9bXBbde0pBzo2u8I3odQV1/fQMrGzenybb7jgI92OPeN7XCFxEd9Z
Xw21lTe1TwRZB0H98zSatGqiMIccN46KHtYobUCpiAYQJvkJBqZ0ACqvRKxktCZtxhdex56rpYT1
0mmEjC81qXuCzEyhMeaI76XkdISuUfBDlr7X+bx9yocDm0krwEal4WGxvmApGCHjwxHtAymXinKF
MNSEr3p8ZJlm6yW5wj+kHKrnTlLL2kDCOxmSsDH6osb91j/7YytyspOgKfJ1qOQbmGebpYIQnmMd
Lcpc8jYa4cMGAgzH1OuEqGZBVaYV+kqi0wBLIA8qrcvj3xtfSjC2uDgQoiiC6OIVT0oXBItRvveU
HhbjGneNM4a6W8b/XKHl9fb3PeJtFU/d/nnWquOdCUMSiwWfuUdHYz3gnbMjnJ+vUuMOclyyeMqT
gFcamDXRuyGDjHs/U6zxX0tMM6HBYGHHFvVaabn3GgCK5yBzLpedOWiEjiA+zlUrJBcITvYvXu16
bjlv9txBEb2qWM6Ke6ffyp0SdKI003VyWEQXzxUSxYM/xJmXE8uWmRwwuP+2P4dD/0Yevte12tHj
0+Q+H1Zelqlu7eLPYWJIXgtBuqX/VRDba5WHSKqrD4x9UKdo5jkSahUFw2odnXLtqYzIzkBg8lEN
JlAXC1gaSatnMH2IEjm551rig35K1oAtYuyLlT+EYInJ59qlgkp2IY+xwCwJ6wFD9dZVcWXfryRF
swRqM2VobhKODGnr70lQfPGFqhZShP6nfZy6St++fmPliFM5htFwcQ5eiv9l+tZG5LRCH8zXMrOz
TZ5qmigU/9Or8HhrR+fO8M87k28M4EMSwUa9Hzwf90XO5fu8DxrKZqGR5Z8ZuRW0LLR9dsrcnNP6
Oj85eavXEVvJVhseoBut0MXX3AnuL05A0e+kSdT4Le2VvTezY8wVUEljPmTQqtrvz9tazTRJh+mn
DFnX+TbYp2EPLeLeYCB82Nzfe9E8ZA3lBDXgW05oxd5FguHORvCUHX/50QWlgPRC2e1xH9RsHWK9
PZ5LCsJHliBpOY7QGlSzjpuZIRNum+f4KFBotQbJsxVmy2nhYIuNg3D/vuGe0ZyZz7XrEg8g1cx3
9VxselZ60Ew6lrnM0DJk7HRNONLYFz+ZQ8G2PfJP/Ggf8iQXoPLj44lA6rdi8m/A7IcG+c2Wu6EM
FjjicIJLYt7BkxuoHTA3wNBdnuOznDuTaMmVTyjRBY0epStte7wu/77FaIlgy4Gh1auF64cB8epM
qqGghT4vYCvAIduj0nZdVqrXgQL68pBGJVUPfOFhkIK67NRPEvSTJKEtiLYQywktd7sKEx8yi0Pz
3GgmNYbnDKARhzuHdqBDpw6zAHcy+V3hfNhxLjE43sb95Fh2l9/wvN2c/NlwT+6M1hhhQlxtGiWH
4Az5dSpkkYaU8j3K+mvg25d6QTw5g6jhNe1NH+/GWn4c/LlTW3jkmkGFSu8vHi+mcx0/3gXZEcFT
TICzPXm0yIKGRzsu1ZhqylxOq+R4/+7PtzcVd/5cm1FAGn7Lx3pjL+So26zELS/S14RCL1WwBlIG
FcbzY9+7HBsDvOdwchqY/FzkbAKspn7HkyUGYove1GUnAjdaCaSYMlY+JjhQCdZq1QVwVDF7SmgG
t14z+97cdJufKkRZdHKTHp35Qbu1degJiEV4zGKypxvw/JmIWLo1WopWVsE3wrNB7p0UhdZ0Mblb
BmTdYO9SIbuAxgHQd2PTGkQ6fE1EZsW0XUjMlNS8sAwjvpPHdtHXzPMNx5K56n85oZG8ExZaTOTb
TWfEcZKzt1eF110KFBvCOmj4/fyTMK5SpJ5xuQSDIwx+jAbA4p4IB48dIPfCdkh4Xtum4kVWYCsM
dsqVEO2fUkvuNbjORq7O34wSA8P8jTtOkb4rt2b6wYZEBB5IH+6rthKswp+ELG5PwYkb864sBzqJ
VcGRgerIwb/noSWVSaGhiIxQDUVqRDxhCrmBvXyCBuX6zma5r6rEndivXF8YPhCULg9K9yI5H4N0
XTfa3yrNfbexH94p0zYSWTtgSreXs2B4h09P1bsrVGDe8Jw3HpF8LqtmrEOiZ0qYOdX+CV2F/A7g
CYjTO21PeXcBwXYVGWj280Mos7yUHHqIzfc/OHLIfHh+KoBGQnWzGpA7kZo++TmpxPvaK3R1n5/g
TGNLgk/qAtP4gg/Rgs2LJ9RJ4HiLyUnoXa76pa8m04Iv1iEpkQXYMYXqekUtGr0MUn8vutqyGyWY
g/Wf8zIyL5KNLaDOrA/5t+BZmU8OrYGP+g6E8TrzlvkAeYZQQCoFMVHekuPKR5XAF1SFnOoJoIJu
W2PVD0IVxo74tXHYks+chv7ItxuCRzxVP0NNZGSIKT4nUgNYLJPda8H/DJ9Y1zsSCjpw66u5TEHv
wMLqWnoysaEvko3qzYSJlYEuRQ1sk7wZ5lz5TEMyi3Bl9TOQQ5GqLUKk3ZMQSciBlx2RcLcNTwVx
iHqVvcIVQMWgya+ZvMjlAkGyQhy/LD8TE37We/fhqfE5OSqpoLCbsQmqm6bX4bycRG2GI2P0JG0F
ZRPX/S6raHZnmzQmFiTItgeeC9nG1WJZgb4LD5sFhUlVcRWXrLvplBtu8d7u1MPHOiet1Cov+jeT
SoTtBsxTETr0eOBWlaZ72Q6E2kzMchyLRWeup1D4lz2UiyhTBkNamuNN5cWI//JwElOGjnL5qIF4
5A1Ax3czv4S24ZaUdYhUlWKwM4BwFW2yLJbuC2KH/vu+wApYPmGCrmL+aQ9WFivOpUWkMQmg6Q0H
eUDIfmFOaXX0wozK/6ZY30zav9WVFftrgLIX9xKXNSiD4letQgh/+vourCCmDsrtCKguy388GzQe
J4KtAemJQC2aUquKASIS5dmBImVaADw8EDZqG1iaqEvvWW+CS4i5zQyCava4hrB9YmnFJTnL7z8w
JEkV7VhFYD+Azo115sbFVxultGly5cv8XOj0kmIM3X9BxbDMksbmH86JSPgMEHhO35lZQUuqnLMn
TBzCmTGB+UiLDoRsTWl+GPy1UGomVH4FMcVKs2L/Ijc0henfCVlwATdCU+NG9XKkgS+ogiiNQ0DT
z/txVyn2ZFsWfQHSVCj3cPhLCVzzlBv2tqvAvXz8YJWeEjr5RHTvRkyF85pwpGFX456nu3AOoRWt
8UvAUbL2xd7aVhPDh0r1gBt5WDhzMNPqRvdVXobS1CjBCgMNfh893IcwN5Chz3FJif8247EWBF1r
SoC7G1zAXFTi2gT42dBg1e82B2Qhk/dsuz2/Eb/FsOKCKLAo6HoIOg3Ta2XjpgvkuKt4QhHYc+ip
uBIGnlyIDjki1l5NK/aQlv7csa/W/Gh6UEqQzhi3kj96r5Eumlv8gbDTeSDadrUv32Xg0wZNEQw3
c+dVUjyQ8cAlKz5exnVTZxPg4ZEbC3YizKGRbfrgp6B6xy8BSdo/uIvuzMNEsv7jCmrd4gwSTbgb
OxAygnsOLVN35j4prG8+mDF1vFVncK9OhJCe3H9Yu/58MZO3pzBqviqYru10RhBR4/SgXR7POyn6
4ZaedjQRWHLhS6UOCW9mlVXkSTsbybV3oz/b5vpNO1JV4J5D9bTbvN879inDpvxw+MQ0XC3VKWYb
DDi53F33LpOZUBNwxJpEXbq7Yq+FWaEuG50cFZTY5h+X7ZmXGWc4VZe0+flV8uXJ0C/V6khwioIw
uTwOkopRwY/KcqRpzTv/KLk9zHDtFfNJDZ1dSEWXAJ5MIRHzqxZorR5x7wKxkRkSG4+mBaWL4z0n
X0rZxfbSgr32TQANt4CtTo8P3ipq/TX8ZHu3MIFjs8Mr66FWhR0t1A5VZs38OIRvwnUomcGehnkW
H/EW5pvpdTBAWBQWPO331t6IazqOCHotmgSzYsokSYKfASwTVpynEgUDr44U4GtH+Yh1QogE+EAq
mMDcNeHPTjYgSuSLYgwUZ/XF9KtIgaAVqZvIu6MjxCmQJgYwfbA8OB0WeQIsPn9dmNYrr7gcKnng
RFm+pW7lWffbLd04MsDlH0/ScviGfXT/hVhHxHklRatcZtP39NUUgvSnetNYOdFwbqd112TPC0Aw
a/H1EO6/mFWVc4jQTiYWo9j30JyyfQkpa+Hy1G0dw8cPySeGPKfBxz48wVg5VdjIkJ0ff5LploXk
wbSFfZ8v41O+uY+OwlGuV2uHDxaGUzMgVMNwwnSdHPNLo+MsTbrfvP1u+dm2VZ6afu/WWpEo5isW
3HzfjWCx/Fn+c6vcEm4eVrWnjE8xC6vHq2eWjRtsYaMmL7Hb7g37R+oeDxwdyZWbQGH2tq7/p0ym
JLGMLjBMxLbPB7GRO4V37byaJVj14nhNDHDJx4MjJwMpV1DxFCCSksAI7ieHTlfUD1fyYd4MgwrJ
AXjPMck/NjufwMufqNRhXMIJFgBkGZ3OTfDF3FdPBhl5SJCaRSLCL1P2KZne53UHIiPa9NgfrIGS
1NiVEDoYe0RzY53ER7mmoRY9e4c9Kk/URo5usmjkhz/hO79jhVz2S2MRm72OYYw1HbcwwmIiEZ2E
QZBPoU4JmW4x3NhHh/UktNj+zzeOUEZiu6cwIzBG45Bv5u38QBUWmNP4ooSVBDeCvRGKtAk3F9BF
h2iVN/Qv1eJoqyGMOoLoR/kC9sVqh7LUPwwdat+cdNY9JSaMos55qCQ6SskeCS1uZt7Jl9KMb1Ss
fqzqivcHEa77QbY3rjo0y3eqVS5rmKExNsB+TISkS4Im5WXqu0e1ptaLHzooobIAdr/MPxSK9Ybm
uIp4KBoe5gjOAhr4gpknUx5jUJMYsj+XhAP0Yexw0R/7VqtzKWINe3egkFbigv0GZV5joKC66WSs
tBHse845hKYtHNmOzQnNzIf+75iR48D9nhpAgqSRlgJ1xkLo6Vc/wZTv8caT77/yh56sLAylu8yc
fu+VkzqfBlei1ba41Oegy8LJvPO6LoKBMiPB/vEcHX6k1B3PlNaABO9rUtB2Vtv1DXJkZTKyL409
wFFXM0DZJrNFsTCSGSLAOnuKxS33XlJdk5JP++c+ndzCmawIBEK0czxiOY1esFLgb/K2ML3bgV2y
Mht6dLE9FvujiY3cd/EgjX/aZBF00sUjxHfx+sDGPEt9e9LLPfxTyxxRmof2276Xj1U28nGHcNOS
bW4Qw3i5CqwpfVuXiqW2MzcVKKftB3v5PVAmjbfN2vTd3UFXFlmxQXxejBTF2qQGHjni6kcckWzy
nZt9ihmk3jTQAiaiNZDbdyTPGbFyzQ9DAd63xgEDdKJeIZULZ3vRRFSgZqcdPKddEH7Lj/2tkvwb
7CYy6ubBu4c5BcPBywZJBcmXIe/OI0AVgJI+aBR5a5OgoN+SMKUFPWnqu9NcHFJSiLzZTLQ3yubP
H4szsorajZQNy297Iv0s3Kkln12tBZrOrh8epajfqMKmjMogKIxA3OYtyOcu/DL5Pso1iZXmNn8Y
f7rjPhVvUHjIrPmESLAH/npSZ1YI5Gohl/ZU7EggLwGxuMm1rmFcMHzzL9M/sc5clceCuK0Mrkcn
GfPG63cBWV5S6pp5SHYbsWy4p4UuvaUD3YqoW0Gvj20nWr/9Eic2avr7A5NluBgTX0r2wxIgRsxi
tI2kDfEbPTcRhs8Ro0zOodEji0AtCR0VoY/Gn7zNliNf89hR/WLvS9anGnpQsB9XBU5aydDshHYf
skcLhKTR3PT9B4dIlDzn4/01/cwNBdhIUM1qFSX4ZvBv+X70JZZ8+XGask28g6nTv+CRQj9C9LDS
JnxZyKHEVx17fprypPr25DckHHHuD/5aO+En8ynglHI2PYMVtd4aB2ok6lkoO9YscUoRYSkCEgz+
CHBVXlJLqHJl3LvbjOxtr9N9pfs2Z5eYnC+GFq5zxr5LNO78kTkhWx6Vw5AVBD/bfZNTZJ+gjC6a
SXgnBjeTWhPi3Jmb0P+X6dtRCXz8AwtcE6hhx83b7vmnkpSZ2qpUMHN/aHwuFe9ajkW6ivNihGUb
E/Vmx83xIoRLAbpeczkmoSNmWQXii+1jfsP/dzP6eaFrh9oXRuL4+fgonuH1b5hyr5w5yi8f2FZ3
qNhLKZEP3Din2L2zhbKzR/Qzti+gjoKdD5TLQydt315qQ0vg0aIAgCITTqLmQjCn1bFJaeMaJ8Be
bH2sRfJ+JWOiIxguUSue6EyBGKazk+HmePnzmE2v/jsDn0SfSkK6IrKNT74JOJzxNSMS921nBgGK
9FV3pME3y4hxLrNIQLYy8hppvYvonM4MOWTRIVJr8qN96yecAn27ze3Qs3kAXUaSOTxd1DY794FC
XdSoHNG34WC1zxpVY2ZbsBNy6wxuLcXgiBt+WgJAGLsj+IfQ1L/Wkn5gBpvE5svMM3svIBiyW1Rz
7G5equx00ZaEsV4aF8XTXjHytu0uz98OA/vTrjoUDrK9TDUcWOvDp5Ek3Iq10QqzLc8AUkIir0Mu
gIKLcywtSdgOHIOWpxgWQqF8vr+oD+RP+PnnbnzFS6fgEu6zJ/UowqW+uXGjwmGgEgRtcbwzLI0I
nfcxlwjE3IFelYkVEGcv5u2wwet3iGHV87Vg8dQ+Yn1S8Ugy4sc3EEJKjW4m39Tg+uCgWceHJSNV
LhIMY8U3fdSPvBorjjCW32wJPUbl6jQk1sXV7ljQw/4YRp5nluuV0qq/6YSq9OysdcsLrlmm2vzH
2R2ZJAcRs22lFSLP8EW3dCJMaFTwgmrdzaw8Ebf41M1ByCYgo1pZ+BBgbYla8r25hmIAu3Rj9r3a
BLiGUw03OuM2cMhkbsfjifefqPDfwOYjrSi6Avn8hvv5eYGBnShmBDZNVol3ag1MrZSlYshjYuTV
PmVVmCHaoxM55CrB/BUEZT3k/4DdomT8Hw/uf6Hn0UDEZ3SxOH4as6M3rDmkRj8fNXow6x4c4Cip
w8sN0AfNdwiTR/FYo3b16kZ06QlcClOqww5jPo9uekcH6LEcAeDv7NjyG2CSaJy2tz51wmpnXbCp
UqfZMZ7hIv6RCkFZgr3g7TOFoHAx7Alwv9zeAKkdAtxFp+yT5roYAdKwHSUx81OP09/s5k/F6Bp3
Kjl4eUwhxqXu4l7o4tX4Hy82QIuEyWv1ylXWdSsgRVRtgB0dsyzt58vCKxs1P4CZokeRfQmcQmyZ
iiOgq3PDHiiLQAW9aWlim7/1o3NeYbMmK1+3DRfXEp96lshMliVRDycFN0GY/yzs/CuWZJnhk0aw
QPgQKi8hhO3+liJuou/fe5YAg6XFUqOR+AjXxNN+ZQPPDbKrUI4or2nzjCE3SZVQveqJiMf6a0pO
ilCTyzOFI5DswnZakSW6angUlfwMNeHRTWj7nKfMRlpswpxwlVg/PMoWUbdT/fZs7MnJX3IlxnUb
b44tuVOzIZap+U6H+UNgYe8IW8l2ozSG1rxX79iVBN91fKzyqL55AZ+5duNT6yxuqM2W2f56Mpqw
79yoNbkAiu0iyp+0pTVNNbndVPK59pRsTjNzuL87xSCkqgx3Lu+HHRLb17/P/KTSjKUmptUGl0Qm
RvARO8InjAV0DFquq7k5OuaS1si7LJFj5bkZfXT/xgTw+Vmxp5ZINcKatwUfNaA4EL4I5ELLa/yv
0AMYZUz1vLjnPSJB5RCLkPTodamJ7muACp/J7EY/s06dNMe7SYogY8w+TgWFH/o6cMUm6w1Ki64O
j+onch/G7MpBcZKvVn79OqqirrLKmDp0+4SAJ4tSTxt5PwoFUpw8mJKKalkpjvuJETbJbWo/xueY
+wJYwrdi+BS6pMnxrMinfbS3hX5SgcJdUD3IqCfmfS/q2dlT9sB5YBWnVWi4VZTHgZeljBTfY+di
8VPxQqjRFvgVnQtXrmVVvk2DLH1ebrUUU8cLUTgRg83/UpP7dqWfMq+MfevUELaFFoegWEJDBwkf
dmdiB2E32zqhXPi/sEGdP4lTCVTi+ztE1ei+fVeR2bkCYOKRF32149wK/arIkE04np9yTNyA8Hux
sPTXZK5clTfn/VAVTelpd8yiR4PjwwlTcvyvdkAKw0aNwKua1GCMb7HFkaxrqVcjs9f5dOqvxeVE
7ndth8L0XeILzynD68rmC3CPNNtktsqASlkMqxaot/e5qdTeslECa1v12vNR2OCEwESyyMo/C0VE
/4XBIfSnMhQiBfIwJz7yqv9cslGF9eZsnLPQQ85OhWLKIA+bw86WSBZLQVllL7zXaV0Zu7zyYGts
FXAGH19d0bybsHXZkKFhizLucnbaWm1EoEIX2jczR48GHiueg8rO7zUlLMGzLU8J8nY1KxR5LAdv
jFUG49zQWq0qguwJWOwlHWaIs+AURcqAL+Hkt/CuHhdTC6/VlmOEwAO1jY9pU+0k5vglpNejNA0M
MX59LKaa6/q1wUW+QdoPQHH35JFAE9S72TyDPRVqdGIgDMnGOuVzFjnht+IECuhoTheB9WABzpMK
TdOed0uRzFnkO6Dwu99ZXemNGU4AnLPKsDNfI/mWVE93eMcEJlpqf2FT07W6/qYcq9nChU/EtmwD
jgATCNj5pylavniujbIGcj36cCSlvrMaWWLg14x5yoF6skOazueF1o+ongRR9BDqoCWUejcIpF8T
i0/aeoBE8tQ2ub325H1rD+Hs3TEiAOKwvAMn7E+m8bm04y1nL4HYuNVFpMUkajYtEd9i8R8C/fto
p301fF1Vu9LkeqkG1xFsA8GbQOU9sJdBfBh5Jr4RAj9uHqQDH3KsLM7qtxigi0tPFv+0biZ6YDml
3nuY4KAyezg7bFyoqV0ySZfKTsexKVCGMvq+24kRvbToh5yZml4TVpdeOq1BKsS/6nQk9jkSUfZo
CIQsHO4j9OZEYe+uUHqgb5TzQpPih4oNu9exff9eY5nh9xMyp1W27ru+28C5Yw9dXDVXlPdW9DL7
bhfht6UZxREeEnRfLmmi1wFmeMXxs3gAC1Cht39eGVjMkWU26clYduCkdlgEnD0o27WmNGGDTwzp
TIiYXNEHLVq47UxfB37Wzwvc8ei0mhE4zcHiWP4fRkOYE0rs633Uqq60w7GqUslq9H71wHyC0UHv
AaVxVdbGEEme7ZSvj5nLVFbxxxaUaHyZ+4na2gTFoCqXR6qBt1Dzsv5V+HgS3/MIQ4uvYRjnligh
NKwn7LA3KibBzOQ+jmhQZeus0lu8vE1tJ2i4ZirB3eEUD0IuVEVHz0veHMzeMX3wsf9R1svir8At
hmzIaJTZ3v+DaomTPKWSN0Tl1DYh7VR45GdOe6oqPKUM5I5tgZwhW/Is9FBCd48EqjpUJ7myYwfu
JKgaUyJ6Zs2EwJur+ur6zxUFag5fu832ddXxTAdGaoIkDbhthK1Zj212d1Wgvi2bj1n1K+6LQViB
cprxugsw9SmramQBCnKU/QJD4b2Afu6I6UiYtbdojonFzGtip7qPKAgZ8DejKeR+RI4z/qGhQDDi
Y8cOphDJNgDzpwdXfozoSJnEzgBqJwWTMIP7XrbrECutBG7PZg1kQ+5BTHheLPmXQnj+fOnGXv8t
8v9PkMvGU3flKkR+7mSzqQo27v6n5UQSAwWGy5N1hZaS45GXJKhcXUt9pDS5F3hdqzHmtu7zel+t
k4+K+E9NlSqZkAGGjfLAXMLIS7v0iqhJ50BD+9QAOUjXMZtLJQeuukXdSDI2LSmGQUfSB0REKkEy
7JNIV+c1XKheJTjk7vOZkdGhRTSjWaoZLMA5NCIJ+SG1s6JZbB03KwOatvN2RmSbsP25rEU7hOe2
aa6OmEbIue3BgfvILDVhf7AZT20mY0MYjDODL74EFu/iMAwHAPJEHh/bY5p8L07OTDblzmZ8UMDB
N/ztax3mPiQY1fcg8g50w2z6ATfF4gQM10JRbgwZsNke8DMlsZtdvWRD0UCFeV4cUuFZlxzg460P
fBNPLLkMgXxzwWuxY0j/qWyV70+Nw7soxsh2f1z94EWXgPIkQ/aqaRWRLbJNX2smFvvJQ0IX5IGX
O32Uw1oAaQlTCirer3m4bHFK27U/r1moQwd2HnGKk1qoVhdZOzAUzzt5pkCUdJSHquvcSv6gwWqG
Xyvu6dAq7Odk7AyI/bXQUpC7AKv9tzK2V9iXK+Tk3MNeLykgQWwgE4TnsC2XtfGnkxcE9ITFVCNQ
+TKNDHEKASwYwF6l44ayOUT6QQS0hfUrjhyx3hjsxuhnwXxAmjRGazkN+nIqRPJzuj2/bfJZM031
rhUTZHgxolMWGIBQkUZyibrAaqHlGBJiXNgAJC6I/KkzJp1lNbcZt+yeYnYG0RX/tO/hY/TilSql
CAaOy7NNBJwJRF9bX6MwncLaE4FWZLmgJu7OgSeLVVPpwoyFi7lTGz8DKim6ChPdsGscTJqyfOje
FFFsR3w9MG/1zIj+O5oMMvjdN0yGwnIRRobhW9vvGHPZ9fEXkyd4EVrzsIrqwThe/7Qmf/nxlxea
iGNGdHgYEUD56YxpXVNsY6KGZAELsnSqguh6Ma2U+ueAguP9eTCXLjfdrWoKy/+mQi2xr792+rrN
uyiRcCOZ6xFGoCzr5WfYHPbkB6G3O5Sha63vWgr3twh74KRQrjUN7cXQhZO/XUlSVSZHashSj3hz
P4FG2qOJiqnHs/bZTLUG/a2cFIaM4SEpr3iXLlslTJ0ixNvDrI5RnMeuYVgs0pIIvhs3hLhOIe4H
/cMD+zEAdrbCdeOpY+O7xE/hTK6g+Jx3f7u/Jd8kGmSgxvkShq9V2W1PNi40M8KZu5rUZzNi+QT/
2c+cDMsf8ICfa54bgomaa6+jor0BhwtKy6+fMlu/l7DPsTf6YpZjN0OVnXt+POLXEi6wWO/GtYSH
YTn2m0eREJ8Cn46mjV4iK87f4XqIu6zHGXaXPN5rt6k3RRqgPc2u+jJjEpfQg7wNgoPXxQ6Pr2Nc
5OYlMldchdnx8QLLId1F4gZbkKXVJzXjVwW2Q0Cs9bfvW9JfmIF6c1qaqUzDgOniU2wFHalxhkSB
Ymg79QyuWwlgYMd2USnUnaLz7q9S9PPiw+POa4l4oU05HWtjN+OvGqhFEejLya2ZoNNnCOZ365kS
mA9HdvrNYoaeCQXpaFUjg699AQvoErPg732mGhb62PE5bxnhGrhFAMc/jSQ9JM1SqKA7l6ZnmEsQ
ad2q8wwpMYWcHfHKpjcF0tfkULn2qUKtwAWXZCUCVPbaCoZ4Gx0tidsPTk9Ac8sh/1GTIyrAVSwr
xG2raAxjW+wsM2Lw6LUSJFsMBKa9TrtsHuu+y+mOBeOfmvTEhII7KHRvZFzm1YD0VRW68f+E2hL0
h05giAd3KwPU6M6RkfSSIWsfWXiB4GiIUcsPhn4kEhhAmBo2+wkg89rWrr2MYSLSMngiKLdduN7Y
d/tfqWLD70w9qXKMM/fUozqMWBeAq2Ys7PWttQty9hCHQDkXphwvgv+FDBsuMrEm8vNp8EhtH9Ye
t5jyggMKdxeFrG3imvKiKF3Dq0HyoI2/APc7o8EwmzvqMx5jfCnX3jLQwUjqXPgWS1Th9N0uTtig
jVt/jg22kSLsxwntKggl0YN83kEhy8u8BqjKHy0a2K7O+K0L18A1uX+y073md5+UHintMkC94hxv
ccGAy2US1nDuCyXy/m1Kj4/eSNZTZHa2cCxQZ5kIDYCH+KWYMKs8FRf19ikMT1hn+YwAp1BM0pR2
yKOR/5StbuvnAL+9ZlTVXvQFPi/UCG0zv7DLplS86LIMd1jE7VNUbZmUyw2QcMREXrSugVFrQlu2
k1Ym6LMGyQC74VezCEvZ/CMMgKEWHM6fVs/jCLBakcthytoNbWtb7rRWv5mVnA9wLZrZOamlm53O
8tPMnmatg9inPkX1fBqxCs+cLmjp1KK3sFrFIFd8GVf1ld1EKrJGtB6bcP84RORTsT3lxvJJBunl
yCs0zDyltNbr8YxkN4AQrZOo/DHsbkXPVtAtY07YzFbWEGtboW1spagoiRgpb12+dcyrVMQEyqTy
HNfvUUxPrvYqH6gxovBfk5+NFbMU+C4/tKbYTqVUqTVV4mrUa44HBGzqHuaO9iYfHagEJ7PunG96
ZtD3neyR6GUpWcHpJvYFu71YGxgAy7plpX9Vqfssc1U97dXrghwbbndOvQSNy4L8RS8zkz4qD1oR
xvG3lvUm3Ngj9PcqwTlgDsd47hPZm6Z4squ/E7h1+8tm3yrMclR9efwaIe4MK1uX4abOmlvTNRxc
U1rCL1He8kT1C5foWCBahE8oxPf3tCxpZzIaUtnElM0wgCWsg7cKSyW6896/Mto/W2LAKkv2OybL
Re8et6mWsdc3v4gWPUiQm9rL+HRmVZc7mZXo5eYjcTaGN/qfUxwnVE8h/5Gb66g3/aNzVTL2PiS5
CU+lgLGVU9glK0EEMqEcpAK17vqzPK07QAVTeOZKcH4IByTkjK8FY+Ceypxux4WC5sLRrQ30yRIT
9de/C3NH7wApb6T82F8ZfLGBy8/tFnQG6BJwt5HR/iw1IqwFAAFpaV7mLvkT61cYLzo8hPXuDWOL
jQqTprGbWhdgBC/LJvoFjlzgHcu3/j+McSd1l73HMAae6+Pi/xVMeCsLxeTSu+fHcnGNXXMWREND
XgkdmuDesoCL1XE8MjZs8O49JoU40o+Z2ISeATFx5dK1c0Pebqqae+7B3kfB6aIP+iU72g77A59F
o6lBnxHflwt1hEpqyofo/vgnLfYVZvzrCq0vvO3lj+tOQ3JCk5XAGXqxS+zKgSTOW+2ZZPN0rIJX
saN7ZcNyZXp1uhK2D7gISQH5vWdX6emVv+oPbxTTFxXEX7H5C5t6t7VLjmYHuKUcH7Uv65KzunHL
i4QqDk+Y/76hLIh/pIN+C0X5oVb6f8Aku8Iyn3Hrg6al0IjEKjWjy1CMtBANGRWsmO/IJTRKjgCN
ypCN9xJ7Qpg/oN/KOuVeQ/cAJMGAyXBwJA1l5pZa8oWVLpCpR827l5qfOqJVAXcG19z75t9W9fg3
pCfKv15meOCzZBIsb6iqPCB0mN9luWMHDCey5IoApoDEZ9PUABTqiorra+6TeoKygRi2woPPflaf
fXLOVTZEe+zZWcI4kv0UJv7+lQ31fdNHrG+nhxZxsiogkhSmiip7d7j9/cVkuU6l3lTFoKqYhcgE
Vaqlj0QIYYNVa/NzFwm1RkTLLiKq1hNSwhHWMUpLjj4kzQpVZnLIzOJcScg6kGWkkvFJmlCLNve9
O6fVkKfZsxMya/etm0+FHR+fF1Qu7QPHQeKMB+zxTn1m5n1Fy/S3Sid9pX5U77YNwfUzWWs7zApo
SD9LdD6Q5ZlFfLu8a6hGl4nngmIoZ7xR1Nk1wsSKv5RXJxJggu0D3Vp/BakzE9JCA2nVkrmVANkb
KWLWGX2jcWyacFpGUjpTJl/Evm1LFZr53PmGFmrFuLpn/TIU3Vy+QdSulp3fwli139rsIeC6L4XT
W6OBNA5IdjxbnfXucjBJeCktX9Lkty2zjuCw82chZZssCElud7QV5H8vzLfAFQYtLXsZNV+yBxkW
tN6UeClxO/yFpO86zkLiQDcD3EWnVsxNiw/U9Dr+FdnRoAqkTjhuEZe38R5t7n+UAql6bMqZjYFE
SsPMFleGcj4mezLrsZgTDzIQpZ3X0E2h65SUIbT00EFUaSxoPFSLPju3P3y6B4m2maHRoYQE8yq8
5VnlOYkfTMjui7Kv7nsN+hSMkD0Di1Pzbh0PuSZW8Vl2A+hZRgEFSiOn4m23RwD81kOomiW2NyQJ
JYXJGUy7qix8b9wwxGlVbMPblBV+kii7LDL3C8FnkTbQv+WeMeOfKRKiJN2HHjc8YJ+9xLVV97Rp
+q/eRmtmG2ib1V/MkBiTFlH+TmaNimxiRhqDbXv4GkvG17ZjFfsrhqqId4PlnnzMLycGGWOkk559
f9EGX38n9fyNV9EQ2gLEMwOcpJ9VJU05omZVoYCgTkLAQ1XdwDEz/ea3kZHvcEpXrrSPXfcStbR/
z1/n/9FFqmKg0z503Tc0txKYkkpTMdjhhVMZmeVpHbSPPygqZgXNRhDDcL/D3wUqil/6BQMezBjC
Av+ly6zm0GWjGmJh5V/G5rftP6yOLBR3sC2kjOyecbUWwFTmDL/II76nQqlH7baBS0T6f1y07ICj
HJ15u0RsAiV8PnHqV3on6ajyS2ioaEaNxim8XP0cfyL1kh1nQ7dE3tQ5KaDRWDly3acUdZu4O/9L
rWGJ5pnDQyk2PDy202Bi0TW1gIwkiLGRGfJC7ZGjtPV5NtTYYguFeUVwrHjRApwxRtOUWz7LTDVZ
QrelgfSwl7d36qKgl1EuAhD9KGdL1KEGP329FYEt7lYH6bHPMlqX9grdlanSrjcEu9F0Pi1Rxo5S
vvonXLilOwfyDrlwIA+mKkfXOrpdO+4uJZLqxlRX+T/An7LabhyiUG6zRwTFeD9WRxlJ9Vw7YAYq
ucuwissoZ9M4zKhvNBn1f3scQeLNa+tooaQIba83FFc8wDuQ4RAQ0kL2Q4XPoawJtvfGrNfLk7QZ
LIU3Lq3VoQdURHp4CZRgWNjZO+mgIYbi+k32q0N2xc5HcW59Fr89bE7xhFgXD5XAGHhIB3pBaT+f
q1zCLturuSKM4Bzm31buon6NhmcY8Mb/beObdZ7HH/K5gEYeusAZeGKn2UVW8APSD+jtH5B/Wrf0
eP7M7v0xp6fsUoVBcp8YznD2pShOYha1XOtrjYQZKhCKUCdGl+DH43MXtVlvomHm2NVO5M3Zcb3O
nCvyhsjgJwfAY5wmGLkntfHGWgDaN0zJpZdo257g5YxgIFoWM83YNEz6ueVR1f2D1wripF6V1PpI
FQlK7xe22ZIC3rNVfwKFIQMOp5RqWkt4YCI5W0WDGnarZcB1KXUE6cnPk8s07B5/SF1iEKTGAtxy
xj3OFnQcwUnMBNknNfyzhX1Gy1cimgX9yVAyIH+fb/eE2OQL2xCA+sDek2mnFgI3//CW4iU/8j9C
rOG37rv+gnKqYBczcKbdyMkbuWTLyCL4W/lrIYxtUsZeATwHMStbFsegV2cXz6/JoeKsoaYiqHW6
Gii7uIU7GUzuTZoZsf6Ev7eBXTUUr1lGp17a/A0ovoGu8AsWNjcHgDgAuJ4v6XpoxrzRbJE3DtRk
5ysOj0YrFD4d+lbO9u0cApk9QeQjfIIYulPS0Z/9Cgxm9GrAkP9K8dFCMo+IOkJK0noCuCXYLKOv
V4ksS2+rdX335OHme02HGpsNi/syqA7a9BpNbujsBcLKQ1Pcc5CKIfU7Z3Q7y6J3YBpwSheiThM+
j9e5PxjtHDlXp0z/5XZGJuGLERTwNOg/pGw1hD+wQfYWzg1SxkaaPRaTYTAnaYFV/SKchWRXI/79
kdl5VNw/96Hop1D6Mi0dvoBN1Lr2EGFn7KmgBnBLqFjQ9DzQQxgy9hkY9yCgqUoEpLYWvP8Jpkk8
Iu1xYcBBjd7unq3EhvP+SXMNTk4LXU0jbLdfgUwwzy9TUdLA9C1yKtzMFHzYApoJdn7bwgyszzXU
wmYmm3vqJM8Gr4b8LpXIAgEbuClbRO7zihtSVTWbNWElNNGlu96ADupAbBMLIblexCqzlm3hmMJa
xLtndk0pmrVrvUfeROhjHZEH7IJRJ/MpWYscp4hG9qlNamK0SVHL84EYk6CAZnNCkTtJ/pA+8KpC
YiFiRgthRtWvxMpdxtQtXk2JWvpuhPAqs4CxYnjfuw9Y/m/qYQoo/O1ZJ96UbigUfgUQuXsBpCA2
Re4NK/LWr3Ccq42EYzC2eayAIcJcZV8OliK0y9AZd0hZEE3AqTRxLw+xyUMTMGjATPrH8SDaos1B
FfRNU1KUGl8M/Ubx/S9H+EvquVDnyF0XtfxAKJib0iEwPw2egidreCX3slPf7DiQgUpqHQzvMARB
qSWorRE5n9TztNMi943XA41NkcsRupO8emBa9NaOHHO1reLjq15SSjTrtiF7Y9qagKg55IhLprKx
xo2653+iVHgZ7/eo3eZv4TnduwU45iGh39CxNIUjT7wQtjGkN2WoFuZsNVIBxrTjNPjHmtYX9qNw
1iX8TvLDNd4DLgJNcdvvhv4/OQ7Xh2Vnb2rjaLIZVSAZ/KhOd925OuljFIRdVTskVTyukdyY+SYe
i0O8oorYdtPzJC/RlR8S2ywLdOe1pV3pWGmLBXDY0QtgH2vFz7ht14iDhB3FJgCcape2LqZlQPjr
RT+cJsfDUrpuJ3y8hBxNsEW9vg00KZ0UKid1Dv4ugM+ErXQrgh0c6037ioaJCZuO+eyZFnDqM4e3
Y549EdmjFJwITuyons9MqfcdlteO4IBHZ17Q6x9w+7yzdNgRWyAhmm2bzyVOX8TkeQgSRsjG2hgD
/iXtkOR0dRgm4hjDECaoj/eOkn+/0rOX2REE8pI2SXHtrZF+K9L6aKOstvt+kyZvk1cMSSFtWgU6
8xtwDwQbnWSgTYkD8HIFiRa/W3cgu1msGud0mgBLiVPuSYK54m95yP8uVFBlWvNcTZ/3amJtI+32
zDAnXh9CCrzMImggkb8Va+oQOd3UVuQYNvcWOEjxLjotMhf0nwQuc9PB7iBSg0aFFAJnf/10pqPF
f5WWVFEZcD/cngbSI6AsTh1UAiUPg50KEOf0LcUj0qm61DxTTK8E0+8HrAK/TOeFuhbQqSTP16ho
hLmDO2YjscvSFWMelIksMVsNTQMj1/lYH/a8sXNR8WlHxW+tUwAq/EkSDEdhGBQZiGWKfM/lRvI9
A3Ax/wGdYpSm7LAA4g4EE9mjFRiKBtsqC5aZMdE73pDc6eccN2knSG6QS3NYbs/GU36/H71ubqeX
nJam0VBEImSHDv8qimp20ESCZvGYx4Y0DvMmtnzLzidPXs84kVlG4YvjwoVR7AT7S3q4LhktZZx+
SLYD2vEOihAlYER+6VRw5kqWcT4SJxfBN4LDk4V71NkDiEn6PCJHCuC8/8vmiW1xfwNnIo/A2L6s
ookqCo+QDnnjraDlRDvhpWzP2Ice6CruP1JUga03aRHBCZtJKL8LMmeqRQDFCZLa1KnwSNppVUlD
khNRHAdZO9j2BUOcm40MSnYTsQa36xiKQri77+3u58B48+GR4pzNcROA2lnUr80NmcFKxu7Dbhy2
YqSCA0m+Lwy9l+mMeVi2PAOPnpdK5afvl3lrrc/hFjVRU0MPldxDXQolfHNh7Rafcg76/x4r5Zdc
rWXSGXaKObAl5FIzVuHHJRRJf2jSRWd128+Pdr4X2apN3Kgy2qdkx63k3N9eNYDmzWITvc/3WoRv
QRaUYVS/FKc5kA+cZPQhUN5EvQuMCjahj4Ch1YpYxHqNXRwzKvW8CXgUNASbbmf8Va+zCFEwL+Wk
F5KWXylu+a5zKLIhmeIFMQ3KT8eJqJPGG4hBWurQepm00talb8meI2qpiwI7faZ81PJ7TP5FfSmy
FHsoVXzLG3d5cpBtDgPhdJqTepoj/tjE+pTl647bvJIKovPKGHeS5XA8uU0Tmuo1N5Me7VwNSjRI
mK0t0S4/NpX+EvVD2f/fr7BUDtHtQqehDWuklYsDcrg17JmC2c3t61T1EU20HpOOmVQU3YZx+RdQ
NqgXMSQ1EZ3etGnK2PLdufyE4Nhkpc8GOz1+ICVFnuCg0aDbvUCOpG7Xhitr3xfskiLX9W7IT8Al
T6mGmDW0Zs/relq84+SVYAB/ISrf2/0tp2GfoHEQ5GVGkPpbXc2RRGkFWKu0SDNlKJp6lvGWCyby
g5/XWF+PokNcGxhOBJv7TAgbj8D4+Kh2ZsH9914Pux64s+GYZ/+Z81IVG9HM4qy9UGljJFr/q5sN
K90oIon/6jscIdlQ2E88kgO514EXrMlmtoleax0PHxlfNEp+53806lLRNIvbLGAk1MSAp2ChzVqE
Ph14dfQhZsYXJuHUUHmE3kWjR3JkgJwg3W0pMD1hhkW7dimlhzsWZDaKq+YtijFbX8cEVAtbJIlu
p08mAFN8Jirr0mZ6+BBNym6Z2heYdJkVi89yHlWL17uyGdfV1lqQFcqe4Vk/jyG81GgK7DgjJ0+0
JKU+M1gwzla/hh1KXOMJlucyA7ldCsvD+F1q1hL+dABG/Q68T/O9gQdKkvo5lBLvK6ra1bf4oN/k
9cyZLZzMMmAB147lnz7a2Fv2u6wIrLGW1FORVq7o+ZEZN6lWaTWXRpgNHxpthpd68lT7Sk7+9uix
Zr5V5GhgstGwKjDIiveljlL80jbPfqNB9g2QelDciSFOOxbbpNll9vaXKTm9WRKteemas8zdZrDX
Elkz067KeveFO1ET6WTXPfMZY7ifxJPCt28LZUy1FoGb6+a3M1BaeYOsIxzEi+ydVHZflNK32oVL
bBOdgATSDMLUxMaA8MnBToJl5MRFlWpHurt80Oncgedov+BSPdEguuOyHq1RJRmX8qNdpkrAPqJp
hRWFLFvNLR8v6UKtnTp1VoK9Btd3XysZx7UiWVjLT4o/sqRVvlLdXokE1GT+AP3LadvRS/tAcgvq
KSD9cCtrSgGtjooamH8VBR0yxAr3n9yJBEsObrqyRkImntZ87MzHUGB8Z9izsDUBeDOlagMFB9H+
c314ybU8QoieYmqvnisT32/Wqg5ceJbBVvikmig8xlhFa5gLOJ8YyU3GY6MJdPE1ZOLU4S5szfv+
SvsD9KyLE3XiU+qr2iaYIX8rT0kTsMXw6hp+S2bD08LTDiIWn58HrArTh3oaXdN110cQxLrp4MNm
2zpMrD6vuT3x1vikW5lbXNvEkVWzk35mSjYCDRGmriMezKaZKIhmp2gfnOdlnZVIvxbVrcVOsBKV
JtcB4ERFVx8ChyXG505klLOS1kzVTq1qq3IrV5O8Zvh87sI82VR8IOYBgIpjAcmMapYlF79MIWYU
VcyYrAo0x6C6d6n1jJwq1YcLzcQY8NzHc1JDk55jaG23hxq6JXONn0a5/STwo9oXph1OMG7zeRSj
q6DPOD83gaFA/AfQVqNZNsZ5K0x6Mbuu7TjTJoEnZd6pipCpTNH5IZsQV/EjMBxN6rrfmeLpUItw
5KSB5lnG1RNNx4ZGSEX4xcWqNn2myoR0b8DrC2N/er2FIdzr3D+dM7Ya7UxPTj0Zvhy/aU5Z3stG
Krep4BAfYlt29QPNxxzTRJPL4Nn/+SxEBuDtb+rrQ3Sc4pi6EfMGEiVmXxE+38LBoSW1mZwNl7p7
Y0Hp/ecY+DZHfTepUIBdftTL7K/1aPJbk3U2O0KKuMLFsvJLymrp4ybqVSlxysz81EvDllNLYfSH
tLoPBlCFYKyeYiZ1RfXqt5ZAvpnKD49+Hk71Ae71irs2yx634/z47GKHeQlrKAdV/co3dFddbHEc
BWyVasS4sHE38F7nTGtcOv66hv3cP/YL0YkaOYF2iStGrGehEqdziL4ymNPlLt/37dzuGBIU0zXO
+M3kxHMNt0Tqy8iXALCKx7OdQ1jIPYUpqRmWx8DaaWTikN3TQYJeEHKhtq/n9rWt9wrxUQcemM0S
d/6p+IHewRRjPQCYmbEAzFWu6TAhxkVrTiDtSLbEmmoExa8y7mcCtmQcdKtvc/rzhbALZthfKtI+
/9ItGUXKe61bRHz6uvHmDCQJoDD+GxmTNC0j95hF1sGUDIniSfpV+a7MhDW18/P8yvqd2Fkxl+b2
AzXgA+21sr/1aYd1YjGy6RnFgWXUSvdOsD6tFnxoPzVm7r6k+R15bHwzWCxBh5ZldlC0MpS3JJ3X
/brWd6km0TGlqHSqI/LNrfNtinayoYSkPkXJn0McrnpqkJmW5B50GnWhHV/tXYcNXetzbcA1CKWv
Ufy+hBLTaI29v352VqdoSgYRDsQxRqLlySGpHzQ5r8iykn4p9dH4PWDZd+PX6AvhUq1kQ3Vdq2Aj
B7nkVNYwp9EgyJVGbiazjhb0ypK+6JPknYHDpmzSY0neWES9CTh0W5CJOiwcw0c+FUS8d3n63zaE
mm9ydd+vvEmri77l3fQd5wCMpGhaeOR9RCct778rN3DLVTYo4gWihanOU2rx3r270LPy8NO+S9r8
yYF54OdEs/D+DK9NhRxMaja5KaXrACey4FHRNYeqGHvIfRFKqn7W01xe0G33L3lUJh7licVup7TX
QDUsBbrO8tgnseEVlFKm/uTyyGj5oUlC8Tdj6vcKeyYrXGIExRl1ykHYIwQAitq/M81IBHPKqtKT
DiuGLWD49T0wM3jo/8ODy8mQCFIm15o0IHd83hs9D/UBNwbcF/xtyDryE/SpS3EBSIee+M0/mWMz
qjCLqIID5cWXeIb8DQrbXd6DL15IROVMMzpvIjN0y/FGNimq59XSBb7Rvhrwl/VwmylKOyq2TCR9
fXbyyce0uA+uBr/AEMZ9dClrj28iCrTFpS4aSU9ELZZ2WJNG2NaOzjUe/Xt5pcMHVMcrCRAfYP4+
2VFqq6cub5ndDas7nZgaGhaXfWIIeEMf2ydZL7nogbZtziUNbjusFW5QQnp9Fcrg2u5L6MzpxHdl
Q/+i0wQe4VC0BOvlPHn3bqT+mky8S3PZkDKJUVyNypudyLdCg/cgERx6SoFM2NNhQGUyvj8MIU/4
j3S7Ee738HCQ9oe05XGV6R1UBAAZYUhIn49AXMRmlZxQ86xyNle0AAl4c73lPR966VBZswQP72n0
TDb3noqAJBTBl965/yEnJAAAMZWJSWxeW7NsySUmaS6+GdqWdkkyT2v3+0C7v+MwsqkYNt48FmUc
bnIggv6SHn7PW2EkOKWZzrVJ+yKSTU3CUjmtDmwqYMM/K6pPfPG5P1JtUYx29cob0N42jJ08x3O9
mAS8urvLHZzJTysOvXUWLpJxYYy4vc+a8+cRvhi6jjqwiIUe/IDksTZ9i5HYiRbVjwHygVL6MPUC
GZFxHwlaMMmPfD/D0okJjcd5i+FFBuBuoJMql9duUrxv4qyWy7qBRTs7b7h5JxnVvR3ymkMKWS8Y
3FB5nwb3fjbL7fromzFqe6CAyS2u3AlZ65M4q+ep3N9cOa+GziZ9gbs83M7o9SWuu4GQMnPOZnYg
LHLahvFqVroUPLTcCjyXTB6WbO9SWPcYUG4ZIOiHgVsffQzKM4jXHyxyxaiticOWE1+DujXz07nX
+GO5+Yi3Z8nHufE2mJ5y57W3bg1FQVFaPzjXPohWbIxZydiX1j8QdhDeM6tLkJvfioend2JIMec+
TxOB5yngu0Uv3Do4x/lM8Roz68WhJKt450k8KvCoRo95OrLVO3Sy31nhth4s214Z2yTHWoYwjUPv
41PmdBZZ2Pqv/WkG9/EKc66pIAU92ytAY6OTMZzh8kARmZseytkx7vaYZtnM0hPPKBQA91oKNi5t
YLL6veNUw+JOKUy8wITXbAoo0GueTJSGkuqvKZ8ze5LLDCgGsU5GCXZnZSxidqH1KBLtcH5KGAtP
UritZpyd9VBKeQSgFUUla0gGTAKrV95GMHQi6hsP5OZ3buJ0lOlGm+jphWBcsnP9GF0GxkAxvWRK
7JEpf1YC71bLRRj4zFG5YGeuJdmbtR0u96AayTdQDuU7scwAsWdvRdWUBSNhqOFl/xikr5XSpkkh
CtRhF4IQey7/OPVoSAZ1jMMaAExkLnySAB5syUeFdsxUt7rudI29kpnC9NbiSRiyEyESu/h1p+OH
moLAc/J5VbOUoCJdGF/iROVCbz97BkfPcxjLl/F8Bg18npb9hDkdyvzbsse4+E4c062rB+lcfh2k
wwr4INsV7iEzkE6BEY90UtDhNFqLh41ygA77OsHDqpQq8nh41Y21HXBnMMJoaeMLBudnpWEccn4k
iHeilsbIPQhngxNlkRAYRjCxBeIQ57UykXVwa61JZw+MoehG0wYTRFHuiI4F1c1o1hlhzThTtPAG
sOTYfiu31XMU2L17lMq8V1eNuC07GE6ts8P3wqtGdnHUe/iu9JLhDSQ3c2ph42ql4EWh4oFJQTRa
/1Zy/zv289NNfF9cpolfjtJ7YLJQPYBYtTxSRSJDaFQQG3YYVzMwcuM857npwV336TKQGlaKvlmV
tqijslDXX21H97dkJhl3jelxIfKdgdX/BC34rHwl9ObS5adlxVyVKI/snHfumbz/q8WvXYwtV6q7
vjHBKP2bXxR3NM1pBg7uwsDZdX/DkLm+O9vx0+mAQDNqGDpM24lRyqniOGDG9LDspf3JI5GhoR7c
AstYLUItzapwL5JHbb2ufL66Hg8X29EInzZJ2mdUFTduC2GbKCfmCf08Irpr0XHIDTSgcmO+9IEw
H10Hw2/zU3iSEA/gOn1wDsa7AjUgZcBSOSykWrhO32q0Z3hN089S4N5F5KaZU0+4EB+vTiEwgoK/
lg4e4v3vQoeZgo+4EcqrYSc89bETtDn/7dvUpBJGyW1/CUSfRAMJi4j83lyydoiz9tTpDP6whfZG
8FPh5b2hYJn5ykLahG5EbwspvqPTX3wPQD7in4JwOBYr/R2ocQbaxT18cPSQo/zc2mSjsXGczOtJ
IMZjIKRLERQ1/yx65ConTUo/iQ0JL1d8TJvjy61dcnaU3ztWHIdQNfcUREcLEjFQkBfkSgxnbOHp
r3uPAFIuToiuuTbfzFDMSLkkJxH1xyBPUIBbOwhJhZuzlDJVq6s39Xe+sXbo/1dD8VTDi6LcdA08
3ENMe7OqsZ5EM2LfIbRoZU3bSscxQxG7u40qJdooBYszRWnR81SpL/vWevMkyNpirI4QfxVAzIYo
N6/Z6mCbA70cvNNpJyD/FRr3ONtWWYkYV7gT1X0MrGMYrKNUEkbs4X5ur7iDr/+FHgkDGV+vOpz6
YPxrzsx1lIHNP9MhWfUwyTk95SLTEgXYE8DMPowQMoWemSuyTMrZmnAfgnEdtFmSdu8pfqKpLW0/
mzyPjKUKBd0PbcjK2VnVpkHhw3PJLByf6ZUiiTtv7v+DSnvHsrn/Xz/jGnPlHdJDVp6ncvnfLIqx
1TuZ10xL/SHcecCNWoWoJ0XCSJ8M7WMk4NI/v5Bna/JQBuqui/BF2z8emM9fXyy2GnkkY15r1eS3
zasmrjUyCcSZNt1jpNwOi0YlMfENvudixSMGhxPmlB5nEMWe76vtyBlti4as9cmt2OMosq6wS/yj
7lRKNm5K01ESoY2pqK634nJZdmV6vZpIftAGKPSFF69Az0VLm/6f2Jhs4U97pqtKWE0Mhm6KxBRz
7NCcBfNS0c5LI0T/AHJXq0S73cQTPE3r916uUt+AX1IcahmUjBMcHX35O+EWEFItePhr1Flg23EL
Cycron5nYRbTJ91CnlCkO4zQGJTrBwmR9enSSGrB8OdkWyP5Q1sxduD2xg5xpR+KUdO3OiDFTZdU
Wv3glNw3GrZQaPf/zvwhUfgRHmmqS9HkftXyj+bLoSHk6s2IDoFeOwRKdDb7WdpqlpNXY3hPqJ2f
q2vuQ9n9QE1NllK06R12Wr5VPyBhTkJXoCZWf0GvHYh3EZ76j8JwpL4nZcQvq5aoDUJGU+Y7yJNK
SHzLol5ypY6BC4k6fSRvPRgLNV8g5Pyo70slhM5pahHcs616huy1Jf04zlZ6s3B5gwH4DubojPVE
RpdZPl0T4PyTwQVz7VTijfmMQvxMUur+Eto1NgPbgZG9YG/+FbgKgNWVaeN3c+VhcC8mFz8LNMW6
D2dQa0ZF4jtsmqShoYjL9gFp5quZSbNYDk0Uv+3k+8FR56h3DrICFJYhUX5vmIgwddPjFq3zpqux
STC6zIGXuTcn6hwxtNrTUtYaR4Dt3iOVa8T4iwm6z8xDfYCodOPQER+UIjkExrt1vK9MRoK4CxW9
TRTHguCrsRhbhEgCg5aIOszS/nyElcavyLyb+Lk4aI9QVj/Q8gp6IE1iKjp7/kYYz5cAA1JqaBtb
SNx4SBEfsv3HyXpOzSgw+tbGiOU6gqlKF9/I0hSIpgLFZT2TDUVNCizEqdNwFBohDoJhIgeLYdtK
a/I3v61szHke2G0mYC2RxNDrYIvImCWe1WPYNqic8N6Jr+2XgTK/gsttvzw1VwFQ+YGDS5kS4r0X
DIMeOhMJSRX+xphv24uLXIFjVMP2MCUXNBC0/2mXGr38c1hN6lRBeb5OZuAluOZ7NtU88QwJHVRL
pmV1Udhlsh86MmHKMTa/NWkstEmQLQWPSlPRQMiH1qegXfUAHd8Baq+AXBigN6uxIfuvQ59va+XR
awzBVVVXjw7WK8zji+bIM3FxEBm0bS7MiCsHCneCjg0/xQ0Aa7mbYK4Punp/JL9P1yUOpSimYrzi
fpbSSLYJSZPa2Q5pPts1h/6lwuvbiuprCNSc5ZGJd+kOHp55DX3vnJzKQNbgPVBNX0G4twQX+aif
ZXbRXAQNfHsVim32adaKpCl5NfbwV8yK7cOR7QOUmnjPywg3ElsA7vjJJlvj/PYQQ6nGkvtAGOCd
VnwCSI7UTYaGeoTLCkYmMUbhMx1blUZtYBWh4vo+Xq0JXF8kAFFbWLPYhEbDkI2OgW6r5VP++f0b
YbYRYPh7g7v1GZHp0wQeQoXu0zxEtW2kLzZIDso3AAe2frpLXOeVECDmAOG7rkjaIzltN3C0kyCX
QdNydhzh/bqs0eG/d4HKZQpr4mEHO5mo4zWPeYRpV4DaksLCksZo7OVBi/RCLVxYMZCaUH3QWw7X
nIET1ijbzcpzP8O5Uf81JTAvbYEdFtfxDENuAhBjFh+aJ6Dlc/7s7y5UPDOynNBEMITr4eA5pHIg
TpPfEhmvFRTf78r2DwgozuW5nqDUJ126TaokAQRtsLl4+BMkhcCwwP4JLtUrU1JuGooODKYr1WNp
K7uwhiQPFG4xx3obCuLWuCnuJKRg2lybYOu23/oSnaagc5cvekY9w1UrYpYXoY7/JNLLV6Mw+LqF
VZuHFq2n2j4ZujNzBgiJw9YADzkiHPJNaxsGcT4WE7WTmuUBypsT0A0VTovlGRVr+D81ivoegdxS
bVwKnsjCfgfGdpiDBzQOZb2Zg+tUr8DRbyPXVBwnI4zrJ7GUlupL2vKVj4Qkd435qsRVP3W2D2rw
K5fziIDXmhxoiue0yEze3lNoe851Yj+bAUf48JwDnInqCcGajGlryL93MKEtZ7Cr2WjEFU58pFGE
yWzN9JLr2IQqIfkInyY4KPMZZGG/bJp7Jl6DQuynKFBK+gUT5F8Vok4oyEn/Tk4N2e63vvmfUYUr
IOJEh0zrdcrdHwXKHd+F6WZ498AnsVbbLY6hiB0Z1vCLpaZO0EWaXXCHDvlOiyaP8ROv5DtzmKja
Q1DJpW7hQIlwzk7dj/CEkM5PGFwuE0IVut1wX3nXb6UmXr14hc0CoaZb+3fo7AnBQ8iFpT6VCSJz
YY71g2xhssMSvK2VyoOdqZT0+3RV7uh9QDB60k6tim8SX0dljHPgLBCvmddwj8DqZN8axJ9OKPmd
Rg18L+pppEiQgOO9m0kJFPbRDL2xTWKse9MOOHMutN9J2PwGuD8YDjrDyvFQwVpOe8hT/Qw6/qvk
I5nou4aAw15QEWDO+RzAOrJO93kOUbXcTqZeVv7k3iTNKWVtoSSqxWaBfCgXaVJHzNhuM7MeK0bP
nAIZ8G9YU/KNZpUacWjJtzyvUCVVegdqp/sn5Pa1fqlS/Up9QhzsJeeVsfIiQ/W5lPD4j2zalAUF
YuR4SGJ0PR2qi1am4vJJkZ1gYanJ24urqIyQkb3UoEkDLcTFNYE54ROM4X9+WkT9OsFu+wQG9J36
P5HfJdmMu7Yx4bx9WgH33+dh4bhlSI/2tUAXWR9ycP5w+EVe19Ti5OawHqCumc6z/+fvLHZe+U7o
QdK/Q2acpjeKp0u/vn0MP0vz8M1A3x1Fnj+iWL8dGN9sejdRPqt3/8GaxiiP2vwIa3TGFYJnvBta
TDT7bssgGPa2h88qRQ1VRCcnDTx+GUeaX5dvzk6S/jljkvfVYW/hBmDu+CWVcSG3YzeFKIlt5mh6
KeGZg0tsPQCGx+Y5uBhtUyjqMkxGiRWw7ZRfIZRAFWvYR9n7N12a3NA0GxMdDe6YlMgZiCi02pmI
CFeXlXoz/Ip1yVAe50xSsdeqbyQcj2zMJLtoZtFylyf3kWzA40ok81sMU5mTNYQoUpJekReiL/aA
pQJ0gkMxeLbSuw1D3TX3A3uyZJFAmfA9KOm3E7QiT3wVKgQq8jXdLwUgP4A9Qh0ShlF6gPazqXC+
aeE94ZXRyo5yoZ7DP1OOnh0Y/1GB6vhTjNyKQ8jEa8rvA8BDv5bCXsiINPLpNksjTjRVLNvYkkL1
2aHc9ferN+WFt8IQjfJ8eCys4z8xxCWcr42MDtcgmXW/QiJujbUJakLdjfaoZT92wlyAOvyNARJ4
ZeIpueb1MbrNkCZIy2Sznj/q+QRKwK55925aFwNU8qB/i9krHcJ5mfSa+boQ217vzzsVo96vAt2P
VLABUlUmTyvoam9O2OErFLnIhYXGy5SPjoTKx48Jib3B09Z7zyZYp/GCGXH6flxROKQakkJmUdcm
+Ua9Z10oHoZgQtDnikT6ZDwkeMKPqt5Tv0y4208DvbKnTJmmu7SNEoygxCIaqqIuLSl5E6Vk1Wm5
0EuAriCmhpBsd2aChJYeC+1MsjKAFt90ozHCKg/xs/rv5pVpvcTRQuoVkAK9ZX/AEoJ0SnjMiOyg
1oqXrdQavMyqM/GD3lJA+xbQAnEFmwW4Oix5pTrZA9YdOBhPvEU1fuWs4PlT3ZOtA5CqmJsiS4X+
iWXP6nFtwtQC043ihDXzVuAqNA8Vrh4NClwrLDSgc6MKqM5GRaXGj4u/Bz7/fYdUDmidVeU+2WCM
2a4TpUOAMrDH4QKcphAQO2Fes22UcpuZfv/sYYg3fDD2MzFuxPT4pmzX46zCZEU8uG6WN/hD9xdx
xpXezf/jZ8PHpyemm3Y7q7t7dhl9DZ7rGUzghwSTgxYTGJDsuNBc6njU/c07ydK0tmdJOD4DSxJ+
NERkCnCby1LpX7P/awcIDvrzU2kQh4f5ltu68SFjEequ4XhZZicaBYLosA7aqxuJvsYOfZdGut/t
gnDGyy8BLvrYJYuR/bE+H0Q685EkgQhKkmk2y8rpnXBhnCkVW8n8wrYJMe2TBmu+8yrroUpa5x4/
3KOVsD/2V3s75y89BtSYRA8HVHHOv7/d+yOIR1o5T7GgJN2UFDlajAwETf1vbeN/+X0DATGazBui
LIRxYATjlilHBjEq//ujtJwD9DNOHISIDPKmV5r/IbyhdRPg14BX86DXEn6r3WVWP9cuaDtg/aqW
z6AJfwUSkmaaVz4NxB5CenU0NT4GcYLvxEZbBFcZlETUY+uuiNDYCq4lGVDPch7LQQPZqpXzhrGh
kgT3a6LoyUiuhWtYLsf0m0zSjlYajYHevdhIV6KR8wpNms8F2sPvsXROoNHq48mgoG3dEe9WcHWY
TBIX96PrZMWoUbf5PpB+BzwQrHVDr6uLJUWgSbUA7tS8tlDEVbr/E2byzkW1MlGXs5cNSgO7NrfA
EG0HluG5q4IkRgRRAxeezq5L7yHVaAgvFFP26hwRwqLQmb8viNRSDHym52SDn+nZUqbob4O5EsbV
tfPSQ6iaBRZvUT/kaVWh8j/0SYIRG6i9sdGGQVnXIApsN5df+Uv45s5ofDkfAo6zIklb3g+pbiZf
fcg2dqoK7CkBTQNB+fDD28APJrAuF/MKOrXbQ3UZE7pnSJnHmh8o/W7AzeZITPBTQKhhRsk2rZ80
ZLUR4Mh67ruMd6HLlOg5pMoevBdOI67JYTrQT15AZHeMZ0kMfeeSJ9d0Dd/STxZ0YO5TNcstOw6M
07i4tSrMZwtHYtzm695bK0QxlU0H1XZaAq4kB/97ikhKgFop6gMCem1bl+pZDF8XcgxI68E/HkxJ
WvFh/FRFU+P6QGu8GoUD9u2+npRw32+gjrbkwSIcgpWxrnic/bttrLOlMvDoH+Dgz52lyGsltF2p
wrX62Kxsx+wTBLMlcXiYCuZWo2ECyGOZxlCP4eI2TGkC/Lr/x/cI9REnM2Zn6oQ8d1+UsIOi9KNF
eUYAZYEIFTm86Yb2gk8tzywXSeTIS8tkvgrk4dyuQ65ra0s8h2VHYhI94HW7Xp3OQDPcgdP4FfYX
P8JeUwr09ZOqSuG9L2q25upTHxHI/rTE1pJeIx3bA0uEwMyVSj4ZLJcS++xv4mXontpmt4gs/ZkM
NtmHyM85MjhsSO57/6chjm9EgP3fzj1WpBMRojU/YeJfcYumh1da4Aqq7ohfQZCMBOllowlRUF4M
GaQ7rFTWTgW5TDCxmcO7eS1Ab1tBOZOQydTOHmvZiIyqotg6YcxzL3yGJ4E2FgH8FjU5JaM4wfKf
OvrCxP+fS9Dux7g331LmgNGWZFcHB6GIzqZdKLvceP0WUInb3KGZfp05y/NtVmn6u6Y3YUR+KfZz
BWjuZ5IYlgvWkX3WQZHlzNlmmSrVEwTG5rrxL7sZWSZa2HsapR5Hab4+XMwOWTQCvFPjSMtVnLIN
TvGu1TgJCHcjMq4+hwYr3HmYTBmSEFiGj+utmiXcNcdHOZZ4AaybDxN2xQUsds3WFNk0kQOGXymG
BLlGTRmvEw+ofPcCpyrfdAnK3gsi98nSHXLrdbZ/44/jj4AdhMer1e31runrKRP2F7V3MEyJySzP
fWEV0AT1kl1HBIDr6LTQGhKWFbXYM7+KtL39LfSGFLBWDEtk0tcWyTJHr/LinrkHQ/zsfNOauPvS
Bl1kbJPNP5IiZ3Pxva+bXqBYRj/jFwhnlsTKcgKSBFlkSLwX9CsVXMTHGPgyUAWxWp/AuvhDufaR
cywDE6/OPFYrH2oySRqZFBd1FcXEau9JnznEIKf/TWnUQa9ZJ4yeOWSMQmM8ZIITI8ttnoyfUhgf
EUOECUd+6xQR9EgNcHnttakdeZHdAvd1GXU//tC9UVadWay7hCScbCFl8yU7fBBYVStoYcRL8LEh
SF7m7m7eACb6L/HH8Ncu/IJN5KhxHs9YQfeIX7R2TCW17qsXmnz3GNdc/weWOhr+iAiF5aziAKVC
KEswrZhk+NXdzUQxcasDRJNOzNhveZLuNU2zGZsxR8sQCf0evg9Xe9WZT1XduBzjsKNdwrmDroc7
4k28sIyXcMHtfXmPKprAnbT6Ygv+O+IQGRkAC3Y2SZ8Xrs9hwwNcJJU7a6ygp0R5mTV9JLF+n2l2
1xrpUlO0eLiKJvMzSwAOWIlK2LyWVsnqshH24UOOdOnVAxuv+jxC9UhAxxlT8KBsM3FjIFG94dDU
xVEmWzoMjucDdECajKALsAFM5ItWWyLsJ0SDRzE4zfhIUejBXywcV2pwCtegyxhsex5m8e1NF+1O
YluwCeZhUAY6Bys2A7UlJmjDu416yJBl/x+eIvKcxcc+EvFZsxgFa+GKw7d6uzBN2xxMULXnLgTc
w/tcl/9EhKCOqluA+VFnxaYl1qQhtKdFLdVvp5UkftexPAbHppN5oz/NgMZK4UxIwsQ6QlzoIWT6
3giwrIDBdOnfBhH1Q99aqn/OMIRsYGt/IQahSDDoHVwakjWl4sZmqGro+YmOuk42XUSZeJ+3m9C/
vPvlr06f3BmS16a33y3mdTOmzQbFF4J9GiB8mH/+eUBssRC2G3UinpBtOPnOqJtFYHfhKgYN7Y0m
6Y/zrDevxvl5Tr7y1+VAHuGfwTKCD5ofs5B1mPmHTfgNN4Llfgt6/CDmYfqK1eoUxKsyjDSmKaK3
fwymsjliinc794+qdu8nwv6sDtD/KzDBhCrZ49SDQ+J729GoVs/ix4TAcRPfKuo20isF1pJJUVKk
5JbHlo6IMt93ndW2vvouDb1OIcxzv8XWLzn2nQB10hfaw1cmpqDz57I4zssagqruyR1ygWLWcvHh
pAaUg8JKr844P6efNNzOKWpK0kIESXXp0X7DkGiuAxvAGl7wLDcSatvWe7+u8G2MhBgkIMqHGPNc
LqzctDwWXDlgoWBWFSn1WYHKIv7YZUqGMpSxaJCjrn5d/enfREMWE/NpZRijqj0omOgF9WZ2IjZ3
ZmpcsvHStAqfLs7wigHAcrGmXUOLmJUAqM55YBza+aEO7tU3MKkkWlwHIkpFQjgozAo81eT2uxOE
dSLBky94zGWiwfTq5LsdJHhsvxl54BxuCalsTFEJCJxVgqAf0r1NTLirzGySlGca5IuJPzfmho+i
HUseU+XDHLYNbIOoFm92+2+IrGVMQ56tCCNun+/TN3Oe+G77jNfBKuW7N+05U7P8b4LOlYgBgR3R
8+FfYABab0D0Y0LJchYXP9e7NnYgevsNX9ZN7bpTQnpPBrd25AjCyaqaiz8c1r8tN5LMsV1z+I3p
dTeHQ1AeVPuh/mY9Nna+eF5l60eYxvcxw0fdZ5LXvisF4OzCWeMXwdkEd9JwOuLEmSY4ZxK/YU6d
XMSS87sOULYv4YhL126GsrNy968V3JyQmsPvhmDj8echXcFfs8vV0Zhu51BNMauJDrMhZYEAB012
XgxV4bTMLH6O4OJXO/8Xk7ZSg8/ej0YOM147/99tiImKNbThAjtL6RkIfysPCUcLHa00/A5TZKod
G/Wo3Rc8wzPYRuC54tGcTrrATOumv8xKQ+LUWsd7LGvJmsMziCkUttQgEKzprDdu5nEP/PxAVCeI
Yqhb1soLucRc4LXHyfvcLATaA1Po37hYUlnj2cZNouBsSgLXYX+D3nMJuGNQnI7sZYtbhmZ2NPac
vX/qz9ZjazKVUjiPcwMnTIyWwQlAcA2HbYsVNysk4LYXGk1TCPlhqz/iI5XlrAdDRc7W0rukdVIs
ZPZEqfsTJEF0/12vixvYl5PHPWfUNblMd2oA2xnA8QR/0BMcU4bTNm8Zijy2NXNlDSbcxQJGKP4R
xdOll9d9pxzLpb6jGhihIvW3vY4+4ktVnCPocTrEQFD1aaGtlwGpoj9vxJW4K+QhBwZDCW270B5K
H1tFibl9sqsObeJpXN/rilPLYrZxuLOtB7tecUWD6FNJToze1YXAkwsfvAiuBfHDTElTRrKiz16T
X46bly0450va/lpa7tX0ZHASRyx+yHRvrh5avVJmKjYX1DwZrVFGmKlDgjk3IU6gOgfQxpSDLGMu
fvzkoG67XEetkEXDqoStk+X6lYlH0f45pbfaZjXaCajTx3e6fQAbqsWN/bMAP0deYQ74k+BPlKts
8kRKmjk51q7yUmjOPwAlwxJOQRx+0mRMm55Ltddsim2Ilwtba0rz8Tga350tqUf2hOMUTH+N4mbu
k8h3j8EE+jjYrqCb/R0MpefLJo4h6MlS8bZTcgeLVm6dB1zmUb+B4tks+hcOTo5SO8YSbBFPKHGl
sap5b6qsdcp7F6blSsXfuwA9RjUxlfeLhoNq3JcqmoOXRU1F5Wub4ImWE2RXLV10AKrgG3PNtGQi
/2/nqbb6DrAWg1hSUKIF5KCIVK/bUeHsi39PIU4pJsbbhJn2Bgc4lVz0z38R1A/+EG3iUW+tmZdv
QuIiO0VyPzwFYbB/6cxxtoWbzfpQYNp48FzHckaSz9kTF6Ti7lv4CxmLTxSAZMsz376YNRDO6VJf
MK3cqavYFPHYXrpo2xrXvFgXC7KPLBlFPXiAqs8/RMi49MBMqxuqni1z3akVCV+4rnQnMRdi3Fw7
GFBWGE19sXM276/J7LY6h5JvaK47l3Ta5zNJI7e63Gff7OUOhIfU8jg7rFDu88lphXxNqKTHcY5A
7FLtvSHCRhgEYOYfOiVnSXHhf7+dwPl1C23svQ3fIoGahmMRgzzxXrx/ZuY5BfeIR/iw69gbHHBE
gw8WXNx++CdAwmWDeLA76OT7wozp7IQoiM7+u5xst6H2n1+zmGzJREL4neE5JIOW/yZ2EQgA1bKF
RtzunUamyCwpT5yiAfep30UKzi3BTiW+JXmlLdBzrTz6VGrUivsMiB5T31Kh9IsQOt08WIrlFhXd
q4Jl1iTxD7KqDdx269bdB/TKldqnm5wWJQF6GnJYb4S0cskMo7fUtJqNkMxbLOXb5arKinhn84mk
6Ybf6K+6pV8cRP5oJuowQg3U6OeDUIIKmPmg9HTs9yvbK7nulHojJLLnqB+UuCPBy+dFqY9ejuIv
Yt4IiH8lMCMWtVXuGqHG1ZhfI1oXr3HmSLTS44tR6hwQAIYh5TbMNrImsYl3Gc1FbhV2ugz3pL6c
1YBqAAIkQlc79sM0W2Pu188UgSlpRXi3ynkA+XD1Bd4DFOAGcsU8J44RZXiJ8kp53QHhwFPxrSKh
Nnph2nAENq95vZXfcylxN16fp47dTOdQf7QMPHPwnba+o+8myg+rI8xlTRfI3qjVqOXsE26argji
FH96m7d4P29eZECJmL4OqJvVpSSLBJkN9vXgC37Y2NFqHAqHkwar3+11eovPmcNou3syKpcVKifN
GE3ttjf7flV0CnPJNcN5xcHTHL5rgvq2gkYy385NekX36XKiEJiTdo+S1mTZFJe6iwSGd0FJAnov
sUJJ7j6TDjcvOUsLcIbMFVcfu/dSqB3x6nzkRu4tDBsLkOSnj9TMYlozcVhyqk02Nj3KglOpFnKR
ryRFdQJpLDTdKq8IVFMbt85mLXwkS4E4pDgh1PnzUQmRr2KbcmjX7jeilTG80EbmXuE1h4uk/IvR
G+6yphuhsZ4k/+Ppfk1alLrN8r8hQnXeWpq1fq5WATvmiRvXpi1vskSpxzcPZ9B4AJs4Lr8cYoKZ
XKv9OKtRTbVTTePEeDdJkvwpCP9u2ShRGNTNKTmoWGYoFjiRW1lqEd2fWlnhJdByEpsHBjo/CRvJ
iRM+WfXybpXwQ8OsuQOHGg+be07y/FGGdvAT2TOsKRXYRw12bh9L3LyarzUSZT5xxcILmQg9YEjl
SHHEnBN94YFxXyhFIz/SiM/OOqKNw0XtE1vdCAQHcaBSc/or3s2uzj1maPx4wtl4Ejp0Yz09TE8L
sw6RiP7Cb8wBeNvxLf10nYg4WoeaCaP6UJVupo4OEGhrhV3jO4YLTv+P2MzPrYrhim4fo5Hdbp+1
sUR+98BvjDK9A83DL9iFcWK/bUytiOyKPgWS2135DF8xGjtFJtSQXNhrydixFam31gHpfTm9MHiQ
3D0qiM2mpQ/1Ffa5ZQuQfnkQN90HrNT3ZlBRWHE78UGkr82hUr3OoUgaFsOy8SOqd5PXkp6rUjhD
v8NxnaN0A5D7KaTvtkmZdVDlJpuxqk3pY610m6BFHAqshduQ7DfZBSkFuKpphvpNvxAvrTU82Y3Q
f2C1rZnOeBrzkU5h0ioGVMcKe/cNvOveyGiUFVGbiCu5vK9axXFIA6XB4s/oWI1D23O/sR3WSZde
7kZAxDvDqWcJKLPafbFUybLLjPRlTj8dISvgTXNxpm7+nq4uFcif2m6bxU9bFt5yrgmtik02bThJ
ya5psnnZja8Gu7COfPeZIQtrA3oi0YWsvZSWHFlSmT4t6jHpuh+OI3RyJtASFlRiY7dWv/yFuPvi
4kSsMuwhweew0Nk5h4tVUOiaQUC6jud1lJUh2KFKA2htzb6Kp6tG+FGMpiZRO8Dyn7r3IfeuRvjw
4+u/zVsRvoQGU8gCwYPfhurUlptASMFT355fzqrEDjg6GM/NC4ssf4oVbG45RcdQClDCviCdk9Jx
EMuP2VSs5lnFYCq6xznCUMtnxunogXbdLCLBFym5vUu27qfTjvBD9FQAtrHnMW7SP4wj8CHcOOQh
7bAiEPRRCpTDndOb9fuTDZsac5oSxMjC6OAYcC0nbBUTg0EseQHhT4Tbt0ySS7iY8jRGMkJuoUv2
E01Ba7xc131nNSW9v6sJuOw8Ywi0VDkJiD8HbcGJOpMY7YlC9plWe5h8sKj0XGxyquBROK6DCCQC
qlFy5PQzSBHHCGYNsYOvweEb3JXZ08McibeUJchAfHekNpP5yu9PxCo5S5gYOKrRSTp+NLqmmfBh
PjDGD323vkRUBqbTyoPpCO6k8fuvGlghI0bXV9WCqmGK5w9udkH4BmYIhM+tUAerbl3dOQiCedKs
Gksr2zlCLF5SxJ2WtRl/dWBbTMTQvNoDEKQ/WHHHrxUeUruK7+LaeCyF3dIjHmC5Dd5iQOLvhfrT
BELCq4TGNjOODSdYag8eIO5wkaC2Q0i7fnmUzjNW5RkoL+5rN3y7jdAkzYdJYzlcnvWwVRM0LN4c
fDBqWPn7Ymenv6220FgTIHn57MpIWFbH/P2i8U/mFyW13ge79LRNnpY1AggiEVor19X3ORmR7dKc
xxnLj+aat/7CG9GxMmKu/R4nP24HUCwiy4mjtQg8QBA24g5M5lw+sayCscSPl10UfFFL8dKiDHtH
7v5S8JjJyNqi/YT/HXVOQL7h/S4MF9cvPHVqV3zzqtx3glyWsNbk0mTlwGa9cY0FY4qsj5vtjosK
GMkueoWeTtiBYiUw02n68qjBzizSYz3DtPN+9/7FELBxZnWJBdf9nluAZNn4vgC1KFepWzbc7bmY
J/Uts2YRcgUtEdOP/NGU0d8bFJepqiz6GWAYYPeC2GDMgFoMvj+GkwSqNEWYGuTuPQtNu6O5ofTa
hOwGvzBxtj+PsPAL7V54hkb8dxBiPjXNKl+rjixQ0b5UEBykMiZ57gysSHcyz4P57jVy3xbYfsXs
Uo58Qffchg2doJPP7a9gmvmn80oRtJATT1i4v+ZCshmmCJr1KQ+bwWj424dGdlmcDxfJh0YaSj6b
oHxr1JcKDFfeoRaRsAH6QQlyIvEQIk665NHSm/3Mh/XKcx/nUOniuZmJHf8IXcPyrvD+M7RFlH2F
a7jQOZHWHalsnjhZr8/6DePjpDMea0mNAvTlnXNonsXE0BqW4NZD2DrvamkZrqSOrqUfHVHOnc7h
FKeFg6tXE4SJqnPc6ZCup5NRf0OxP5hLbM48k1DB0peRz8HIYTvTz4L6Nsyk9yH1BJkY2JBbzAAL
Ezf0HlLoUlFurSxn8orzPLektmILD3mOHdRoeB2f8EKMvDbPc3IyKBnmCXxBiCc/rFG6kaVRFZKg
AamYn0FLxI14waSS16z7+R/UrY8ri+g5DAICSk7QdBg7QwMOsTJa1VlAak2eXIGr5fgWzO6pndBd
rygbha4liuFJKLnWbYJli4LhXBWlsoGtYulx/qNcbMYHlvULgkeLENBWUhLS+b4slIUucRnbqIfh
lSU/f+Zsapon7WKM7w/xPxSK/ArSFRbWh2kZapdJrDE/hJzrEvoEuXwW1MyPW5IqZ6zwHM3xNsQK
V5Ys9bIqsJKJGJvzumMK7VDf10HYkBKlkTK0T4xvt8pf05xBLyr6IkWDx/lPSWT3Eg8lS5w0IzSg
28uUve4pl6oV/5CzWqZ5NewpWPJjhSRtmy7eBsJQn58OcQas1qXCDfUt3kHnkMX+7TNNXJwrjAxV
gnAo+bFYLTiNO18cQYPeiJZmwXCeQmdEhZv4P6F0iKnuXKXFZoJXC5xDQX6831TF+7F85qgRkHye
oa/NN1s8oPVxTXV1a/bSTu4sal18W0+L4IHSrkeJx4CAyE27jU7NmD+ro74MxTeCQUkoRijYQnWY
/un6w7F9QrKZmlLdmGYfw1voKud5T6NnCuY1Qzk/0sfnn68h9UDHTEDQgyHH14zcUkdp+bt6XYSQ
aPbil9UoaEoFFUavPGwndsFHWeSmd6TdhDMtIc9PXBg8s82Mk4MyPnWw/uswurKeCMs4M01QYUzG
Fa9taMvda+aiL3yPmJu/MCvm8CftpHmMJp4PZZjqaD/WmlRqe/HekAtv+KI94UcP70D6YDG+EzWD
70StMCAdU+StL4b1eSA8zVrnouhv7ezkHr9Juq2QqRGD0bNSOIcvzHD0CJjnzt8bmkq8DyKguhLi
W0oRRnSmuXwzYe9apidmpNAFWlm6BwLWnlokzrmU0IVpw1xThZ4rVvMM8krBBGKJ66c5LX81WTQc
CPBdtVIkfeRL8og1DHw16axZeiZQE+Z/os303PsRSYb0ZogMvbmfmtPcvrA9JRxa+9cdfyQ2IVP3
ZqZN0XRQ3xrxftORpENCWUgHrhjHG1Jl9Pr5WhS2ppWQQDhPl3l+Mb7waiIzNUvYNzl+GHO4UKIy
qkEG7B4r90A47LfDzBofTwBvjEbpH7jlVwAcxV1vzK6TMSSjTsc2jt01RmzJvtjHlnMSHwSztrxH
raBrdZrIylZ4VIceJI0AfHPA6Fb1y72z03ZxRqyBNzTwZ9NjB957lzz0NvH/v1Q/qDG54mIQPbim
2Bzf4rKETQ6QM5HWjBhqNBdYnk1S1oNhXv/aEj2Yc0meSKrguebCc7iZKG5VNL/mvcri0QouvjV1
BDHfvNAbmk5LeySszX35wDY5eKy8DMtlGW5wkCdpEIK/A26l6gtdzzgw8/EfravdX7A0ureeD38C
Fcwzvk5oIJDzqeIuavXlhdX5isXpC9CeEAF88CYQhBQZJHCm1/CJyZTfD6Fg0SiLbBWoZ3QZ88QF
8L/dz+ewPl7YXsMdvdwvkQ8S/ZDEbVv/9+C3dnEbGq/bFZft6fK98p6WdlEcs1O3FZSbhiKuGHoB
p6RL/mpaze8ILrUmO+2RqJ++ueqiM7Fx3pCyq1BRZ2ZTgoyjEyOkmMPPeMfE5tzKpZb3WUx97kdx
RSXk0rH1FPlqFZvoX0M5bNsTuPgBVvbcQpLLpBauuqasyUzEK3vnHmM8Li4o05j1N7gKBZp2402s
cjdhvRXozxbvme1uvfP1wiyPr23Cj+9mspT9o29x5eW6/sGtLeWrv0CnZy2vIST1HozD0DahtUM5
Br7aMSF0FVFtbY4K73CqqxN74VGrOxm/VeU5hEW+r4Jz38qAQuPg+EYOzAH0kFF91G1qN2rVcl+0
V9poSjURuj9tpoHOl8Hic0lYYh9xbgM2S0hfMnCmv1oQjDRSkIKTd5FDoL9ID3fTM1eMyoegpuZl
0Ml6frTRBFvhrNkB7qdJd5Cx5lIPZWIgfIbmo5tY++LkPIuSNdHQojlab8kSycek6E+eTRyyqoaQ
VWcuTFz4sWeKyS42XT9Wb7qdBfbNvs+H5n+Sfc8zD+kkUdWO7/4zLCP+2SSvh4ndfAwMcCAxFXhg
hR5GGpKwZAfjvCHUWupuk04VIDjsBjUHEBu4oDptY4WqK9kTtcCZSawEiX4Ae02wjXZRpDE6Zgrm
xnNw3tewKK0PBRMeYY/lkCRMmxp/vS7z+47SWsFUWD1FFLG9WvK76Tg/gIqR/2Ktao90cqAwFHez
nLMKLY/rQlWHLSkK1s1Ln7O0KYu5leMyq0EyNLglq5CFkFXUfGiFhbR12G3WtyOAPVhlZo+rhxte
htp9AdF7sq92/XMZacDgbRIMrX89rL47CTTHlVDBjW8EON5YlD8aTC/lUhNZ37K/rh4vNO9QuKc8
f8cL+hut8F153JUqXeH0vWrnX6nbsBAjmmUd85q5drZdbVF110/5PrYmSLaQYVDI3fFOEXUhOn4+
/EOfxQR2MmGzXYST/uERxpbVVtTutCoFMoGjR3EbrvA8Eorunm879QYvCQ1RWyI+zAgkPHagcRKk
8JI+MyzUdLR0GAivlA9Mm47khh1teI4OxOJ4yMTjH5+Sq6nY2XDpPJsnNQkq3GkJKMoCM5i4N8Uy
Fat8MCCqNatQ2zpYNhmvLhuJDETPoyig2fcIHK/Ri2QrjHtzmlenpmqZAAjPdl15hHyc97F4eap+
laMhd5P65ESup269qlAE/0orVfmi9R5N0GecWoeMcicWX34zSzEccx0zXDXC/yjVnA5lgvBySzQu
cnhF4kkOr99WhR8gBuyPiQVpIM4CwJgEfqVMHsBnx9ySu3IpX97gIm13Nyd50QWskHpSgaL2QRcQ
N5Q1CtbJpdaWNxelzZPGhbaT9ho4DzUhnccXYHrOUoANrK5+08p9eMh7icUsRkxv/lLIdDAWFMdp
ATtGs/+itectLkVuAuk3Xzc7iZyf2NKwOqbROBJwvpWL/EYiWq81X+OlOgB00OkuuppVRNluikIa
KUFrsbXEVG69cePiA8qTOFk4FclME+Vu8AU+mOnbRtHIRsQC4SLd6nqvN1g9tOcRcy3S1/mrTOju
R754VvxmroQKYAvO5gVSEI2hSjAlatwkofBoaJgqyKQibOqMh0Xun7/ijEfTtdiDeXwGvdUD9V76
Ut/7aLhFvPIMdKg3ENignm0IGjHk/KcJpDvrbnZHRgGdNMzx3NTsqnyjRZm+TVDpQb2FFtnGwYr5
u/9iZLBVeqas1h5Yusmfsp+NEvsLKej5bS/z+QpeCEaOC9mm7lIS3xVBJZ8e/0wXc53B97oIOFU+
uRxtUvkIdXQT9c0Dgdb0AlxqVPj8Xcfs2UPbyZpVcF2ZOqvY9zlILPqkdkDuDkLLVX5vYzm1R9xQ
/UhKMbRMveYEDZPSkeZ/f3PO0xjdmPzVQ2Ymtx2oCLESKsA7YM7L3y/wyKmHBHcQvzl33qMBYBgw
3WpQTHmx8Dfqv/QKX37tyBcDeUCgTm1NHvZc69uUDdsw13rfx2A5/DllAh3JCUAMCsRDxNcKBkvi
yDIbfRcVai/F2ZmcycAZiZaO+dUjJgHvdRnlyACnf1nZ3q631Exk/1RK9dExcZZDXHUQx0Ut3mOV
UW0RA8m64a8bUvIoaj1SU53SUuooG1DzB5YVSyXwsTf50ODACQruDFwUtf7K8szU9IS57Ouz1cjy
edta5mP1rI5ipUJhylItGfEYKM/+teHsBvG8bR4Fh3Y4ncHwh3aZCoXmMAgZl4wU9tiMbv+d5Wyh
4G0kUCykBsHK72Q32dOJfzegfX2I6yRp7xlkZruT+N5hk71eA/HBgZ0MptYhw0GoGJbNr2XhgaWr
ZWqrN1tkzPoYuldSLnp77nDqNdu9RvJ9QLEcQA6MFouY/ubIdVQ/cvwEBCebZYKD+jZavRybVF0x
KGwVeX9G2+SRce9hGcBWCIskdDdnDq/Rjp9hRXykboldZ/eZAPRwwMosdIAdCWGAfk4r4H0QxzDh
N/wYTTs0+RRtQdJDhdkqDzwJWAAHrsBTVpsySz3U8QLxmVfxLAZoJ800nXR/Sf8PiOzwdpKvG9xQ
fc6pqKYQSs+2Il+hD1jx1Qsq8uVZ521a6ek697kBQ9OiNE/FJNqIjeYmlHws9afpN+T+qKeOrMXY
WuliLHjmK46vQ9v1RzyrO1dXozjPFiWzVxFmDMk9JcHITnrdEtLXoV/P3g9LSx7Ji7DmjoVMiB3a
5voWzGgghGmzKEaxs5zwwMzemt7XIPOUr5mvtnz6xC9/bzsBpjiIFn2vFORqYtHrJRwmK0dfncFq
VGBqOTc2X5h3i+DAOfNfKuKQVUQt9KLkhl0ZTS3rPNythEK2sGliN1NZyLUezAqQN78hzRNnN0Xb
P+ZsVKnL1OQyHn9Cqj6lRP2fQPmKnyVUc4YufUZSHXurL4ng5qZBh4QnyFp0iFrsDp/cQoWHqXkG
Bh+J2FDkyFU+9alVIVHdhGkj253L3WoPUV5i9AM8QXjPcYKemjXC93BNSgW8wf9TqV97YrqURkut
1JjTPibJigcY285xmy1eTLOvGM5GGb9ySt8GczMeMlxBRA/cHj0UbFdq3HX7KsP5eC9vABlMM9Q8
8hKQFVuk0gBDK7ttX3sVbaEyUHYnOMoIEyro2eSgOTrRDYq+BJlA9pQShyAJwSoHXTg8KaFnUqo/
dOqybnXEkzy04CKMrpd7kf+HlODZyQqKdoPKtBlkVjB4eGZdEctIF1g8kTUQbwAVdj/HxDw5UlDM
1+pI8CdSUxgcYgz4M8w9tdDIiOzXx9kfaPmbX5UcEFcV6+ucSe9l3ihomE5vzcRuEhWbBM1UR7xm
rqrzD0Fs5Lz+i1dtjkbaRx0Qgj+FqkFyarGc0OcBv9nE7vIB+3A7DaN2hiIXTxG+9ROcOnxpNBP/
bwgAIBSyC2wrRdHE83i+BB8CvTBGPk5X75iZS/gXcx/qGw0YOxUJnLKn2ANUzzMDP1gYraBAZEgm
32TTW6txMoOSKXg+A41nE5S4R6ObDUnMJXsPbPUMMWOl8SHSmGFXfgg5MZqpalcpKHkpvqiRTHK3
Hv6XQmVU246NvvXw3UGHeyTUcyhGVszUQBduTTOLyjv1CVN8jL65TuskMAXZtqJ8VRNQq7D5zU8H
9JXn3LrhlBcaQUEU74Memuj/e8QBP0t6AOMZXVcMZD08VvlpmtYhC0kETeURFffNJeBLW9nrwN0W
14AA/h5g160hQMimxWA7Xuq/USSuKFKHmrNk03Bx4qf2ckz3HktYaDZhEXQSweSOlAIhC3rCbXlP
fE+oKrQ4WcyTR/gBQj9Q909hm2fsEy8Ej/SJx4dvp307+460Z8l8bByZsjZ5bIjlYZe7ZNOPPXyK
PrOqEP+SzwwUBCVV43XuSor9S3DhPpdvIFTe4q6pa5vsRU1/GKGDtmHqd1HTyA0Oj3jzbcmhVmOR
NXm/M1nhYGvt0ByCe9VWYXQf59II4ZJ0QLYqbvprAqR3/beebk6+D9otVDKIOOi/ydh3EC3Bw3CJ
fssj4X6w++Mglqxnar75y63LMiJKO+d5B2FNj0TNtiDjV8Z+i3HW5e+fk2Ev906l8esisW641aJX
9eyGsoSmXju8jjQ+ghWWNgoD6zjwAiIRyKQAZflBSQW27D7RYFl8bIDRDlcC3EU8pHUin4cGvPxS
MXauBvRfNtRns+pJ7i1EfdVNefg/RQHxOAeOieARq2AWk2MiK3bTl5HhtVDEejgdTtsrKj78S9mr
IVBNSszWF/EH/Yg4ZjAreQuSP44Lazh9+RGvLUzRIJfqwvRHWovcrw86xZnWprjE65UDS3gsq3hq
zzGcUW1ogdgY/KjK+TlxiysKNnzLXjzNP09N3vzJUYlMyFTOrQQli2oJcdlxUhvJPlSoqu5Q6BNp
rQ0T2OSWnh2XRjQqNewuMd09klaNboI0cENAG6p57aTfpw3jZuqt0C2T2rwkG65qg2Y8eH36hVqO
/DEnruR2OR4lMzsGJSoc8tQ+cL2ARKQXE28tFT/MH4GS6hfWhLhQIch/sNZFiAP2XhoPFJEjJ0P7
7qg1D0/cChUhFGUexTEM7flJtyauv+ZEqevBqxowbTCz119jR3n7OEFHilEQ4Ty4yG+Mexiljlqq
DHXaUskJ2EoRufuROHRAUkHPLT2SQVFDKr5teIZDBf+tHu8c2tqG+dhgkV3iuYt0GB3F07XC9AFe
8NFbFGdAizLNsyuPOP2hipAilG7xEKjexJigfjTajDmVqEqXmyj1sCnNdTxwKIaxAgxnZohCl91D
l61ksEqAn4vC0qPUwWpLnwhm3o2SYyuNm34lh3OSOMWqvbmKY1xpGJDkAx/5ldBiOmlRQbB6kFCr
qZ7c7aNoL35mOg2Ue07MMR6i+sRnMmKGLoTgXBmcH0ijoEWux5C/zx3gqZYoOnKHuqBpb3cuGluq
3GzzrDomzI1MRPHm4soIjIvYdc3aDiVjdFaXFfFmdUhaaMq4f5TYUM6t3OvE77XBPbc/YfZwUftu
iMQrF6MuMS6PBMRIXbRXPcCmRgnaH1H9x3lUkd5cwodvAZI8vMIblaptZ77PADRdAQMgFbxsUepe
K95YF+zOKxibbpmxk5NS1BkZ27devn3/fu9AJnjMIyoBXPnhjT22Usc0WQoWbwTSfOakyYb3mwJv
4Ns4SqDTocrOs/bxTCO46Egr0MUKdriWXZmx4tFRx9B6x0ZkgVC52R9Y8YYHlu8WQqnu4TbiLbe9
VAvfZrIHyg0pRlW9QBntixBW4FBlNi5+ahMGjbCTvmRvUnnpALoiVyY590HyTftUzLJfImURimfq
x4IyQniPc/xEz0Qm+j9NCSm8UIXry5EiG744JyX1g7HB08Czxbx8CLbB1J0/cMsDUSjoCJIV9QrE
oF3830WG5EaY0cFJPp3e3EbiExeAKRODsZ/Abgie12L1QCXnKqEY3cMFM3KgMLTEi+z0xUV0d19R
MoeTJWn+aWBza40M0ZGTGY3q6S2VKk/fq22eG6FAFaY7AwxtlvBwhZaGRkX3I9jlRrSwgytRVjxQ
8piyK5VyjT7gcAVD58/eF94REoqjWmXoFkMaVE0HrLiuWEZ1dL3PCA+kw+fOId6pygFJiaJQSVfe
CdG4YAozvzer47aAfslbJ581Wk7TQdxyBpumu7UcJmIuxepGBMci6LItU8ojziztToq7KKVH2vD7
NR3UjldNn37c8Qmu9beCzL0c7YpJwK8oPYWP0RX6Q/xChQsqgYRdwJ8RFcpqAUl6Ku1cG6Kab0rx
mSOyd05TPd/MhQMcnMQhRPKBRNf81BrYbsf6o3ItDwCB2P/JudlJn16e/+M72BWmWcg3qwz8q0xF
USGDZNuKLeoP3pjKT6T3V8OMZ2AaKLWBVPngNA6TMOAIEKzeeCPH/kaE8IvAfHM7GA5TKmD12mrO
dsFj7jFj3ITMeR09WpDkoUy7PFUMRJxGSEit40Uo97b4g26h7tH72bnNsOfdFmLjhLMzk2Jtv6ry
TNo9SeU1tMkvPVCx6JWXXtOj/NLiMBAsY4hfk5xJqBXVlotzZl1fSuvLUjj+BrH7C+qdZeB9BYwb
FqsSSzNzA0JdDMDPnC2rtlNGyDi0eQHjrcaKod25nQkJUBXozZjbAB29lOrUImZQ1EHJr2FMpIyQ
DIzP/PQaDlH0L3DOm+oIuJmkSd7QUgfX6i232EMS5V2b6Bcfd/aXi1514XdfbpKaAPuBJNr0vEev
KAC4H6I4vVQrRyhqZIYKyspP/2ONc556FcH7rcGYHk8vhBy09H3cKGLRgu1CydTsWLvBZyRy1+TR
g1wKFF1jcgdLxrcLFEAPS/jZJwE/OsntgAbTNzaqNUkCMQweahZqC+c7YxTmFbm5EwItT4xoBVhd
Aqk2kABp8pLB0Jnpj/R3yGCtH7kN59Kk+9dzVkN5v0UYFVSYYLms5CJ+o31TFsrnKWR0qiNfiNWe
qPKxxW3Gjxo6unyyKowJjDBC9qpsqevjCjWzt1ZRKt9Nl3KYOHB6u10ZXfB7Qe+qdJUjkdfu/dmH
c8W0spaIBt19CiwE31IhIRAQMUrWYdJniMuECnueeaCNOqpLhrI97tvuSCKgT4/oZxT9eO87/zkx
jm0C2rTsS6QhhzT1lD4sDmyHdOBmO9uVAtYGFBI1r+Ag4jvBkwpwJ8Q0VmxihWhNzrPlhgfJydvy
6y8NJLDn1GkQa8Tjv7SXHD5kCNHNC5MfG4otXEex4PGxh/yuR8Y8a6T5LDUuVYQ3fVak78QrRwJk
cr0ygSTYMeg1z0NqM+wyN/nNzMT7bRQKOMIgoK2cIRwr790Y1hRx2mEiAkGxlQwKp/amq5GOAn4z
ofKtMp27y9W81XyFo6DVxALSIAIYcrU71Laa/fdW9GSjmNra6CBwGwWptkWbvSyQoauBfHC5JawO
ptxDtlXnG8sn7cZwKz941icSLk+UjluVn5TxmIOiElmREySR2JiW91WSombYN5IkrZ1i8dKn+HNH
XHFAHJd0mKbST4WcO6eW0Csjht5fWWLMI6BtnVTkhQmq53+dHkXeMJOTR77ux2J5R1Y7Lef1XVI0
N1NainsZVPQM96TuxlwuR0fvJdIvNYcdwhPq/ehOdyoWnFX48zLcIjnd0c8HTmvxj+v/s+tz66Du
OgMi4JcZEmdF4FlLwrDoGxoUROC4RJR5c9QCugGBYGhkU89pHPa+b3eLY6tiulMz8lFcy7S6JoWr
oofsXKEGEap0B3qW3VlI/dWRqx+GmRpQ8Zw04NvJFraFnLL2a/5n4HoqyWb2FD1tbKwfs9ZhpPf8
H6iZtW0OA84deg78d5s4AhfT/EPt9t4oFCVFofU71LidF+abOLLun+zsQ+/uhvrFgbXqvQCCcqOY
5oCzoQhKYRuxQbciCTDmgvkufUpLhsD62xKfsLr3aVtFN31hY4c1yxJk7VRtJOppObXvDziic2L0
msrMhUpd9Vo5O9+AlZYjMbu1PpwoqlCl4lj76ticDeziYew5/TbeObpizd+8/S/5tz8KKmcXUYth
k/OI9comGx2DcMHvy/RU3YQZBScgJkw9j5YhR/T035AwR5MlyCfZRsw0ayCgOFKWD2V9jdo27aeD
eIdwEuESHsvdRPX4i/jMUYyBhC1UYY80V/Raq6K8zCoZy9fEjhNvco2KhsJWRmQR8LqK9HUiWVcT
zKiK1il8ESnjinoIjisf9MnLPR8hA4JOHTGAFtwXprL4xl3XCllzT1UPgSsjsdHXPAsUg8h8WokU
9t6WXPlDXe2P+PVgTeXUDPuaNeAn/FI3miqxSma5cmcIztqfkwP8aAbCVjGpAMJMPS9Iz2gTrSd2
LGQNL+CUfFVUHfusc8xlk3xYuONKkIyvmzwb/ZqV9SXHR/g1ZdifZ4NIb3gGADHlSV0cJ/firNjm
4CgXJRnEzw+uklLYxhri78V8FWnmfUsW9VSY/qZnzEcfbD+V0Z87LEVR4Jx0LNvhQhKGuaX/G1G9
HBvnOuHpo1HDVDSUPF4cTyQjRDyi0530hR8/JbuLubj9lsJA8C/lX5SAD+E0JYaHEBES/Cm/nVX+
1EkdNcy0omKTsXseOq/QqjBJpzdAdSAas4A18cZ1AS7hj6iz/UHFkU09Lr434dBpW92aVEItHfXo
l0tEyLpreMeU5ek9l/Aa7tE9Ic+P5eAiNS/Pzb7clijg3OZsesqCWo+EMtH7rw5FO8N5xHfxQ3I9
+f+Ue7ZjuKv0nIghIh42KrGwtDyJ+2+lnObw8Np7ANshjouBhIFJ3yqR4rOS6WaoO/pgJrSAgwfw
vUIc8xOSFgs3nhVFaUxiraeLYx0AspJIer3w8n+tPMqsUP1v3I7olQpRmoEMjwWq/UWLh4/1Gi2d
93ihBTzeJWBy6JElHNEWdhEUC6TI/UY1UYuvP8j/ARu1iRv0soWpgXXA+WXE0kTGOF5xrfWLea1O
nWh0gxydDf5EFhz9xqIz002OHNW/lRT3F2rM0eeQNUBJ6IJ4KUdernct5L2Orf1P8elj+sWoqb9a
7rNp/gemB/LnNXuMF5rzWj4IJ+devEtibQ5obO3vB9puiX9g6u9WEB8b4eAkFyEkKvk3HJGUZLIG
o9HRrCGk+Q7BhubByTchZ/8yg1zg6nmcqZefxsOSqpqqf3BP/ENrBc4s/TqH8EUSLMrKlb3YSeBf
bCOu9r5xhXI13i5Dvavrzjd4acnQ33H77pXV99uvxFU+xoQMz186swKCknTa2Mhzme+dkgYK2vb1
P7WbzeV4OAxzipALmMlJYAZXqMh4uvlnCWyU5XEAjovdiMpyiS+8V6d1LSFpaDTyME+r0X1SJWNd
kae09RriQOs0AuN2o6rBkHu5wLn6jZeeiqnIYT4bNpsmLscR4HENpiiiv3G5QR6S7p+G1BdgvtM2
/LspC6uezFe+AvYEUaRILNDXUOQwf/xvdk04eE1+OjvQl4ECDLeYOgfgkQBXOzb3yszKA0vjm1Pa
vZVnGbin3x+NCnltr3A2zuDS6VlFGf9Ew8n3uZFLLDRyGxK43WB6qmG4Qvu/S/e+2Dj5cFQsp+Ya
PrXHyezZuCZfZjRViSodY/roZ77MCoUT2ONonDhxgM5YXwFA0esAeF3T8TX6owvpJIGnrnmN/LDW
5iZZRCg9qPpX6006tM/n0S5xTIxpfMzNneTdUEIU/CtK6pf8cP6gGks3tdJ7vOw9Lo8Jy2Mq5KaT
3UXQRINOi+PU+govy2cgHnztlrHu5k11tHaTUvyfpwrfC/yCAQwsvrBZFY0yLMset3EkQrveQbMb
SsQN40xa1+pjUovnxf7jniEYbA7/Q2AL0NvU/7/r3bWH3DDylZ+dBXjjHyfec9VBufm0rgiAb+CU
/icRhQ87gu8Cu+vrzMloLOvTYSkBLvgERX0U4QzIWgwKtwHOd5Ik6WRvUFZA5x+oMyKmCiuMps7B
SOeOA3HuDOZy/rJfdMCO9sjNnxoUxn8gthebjfo3xg1PTv1t1Qty2MJHB+KMcInux8qfLpS8Lx1k
xP84PE75lec4z4a5VMnIZ56hAq0B0qTE8CBgTp+7PtgKC94WA0sO0gi5qQ13Wz/yHD6rA8t/Yi8s
Bj8102ky30uqwp9DgxJRXJKYcnf0NMsY/wK8dx91KtXj/x7sL3M9y1fwX5VDmNf/t+QYIOEMMcQN
0r8MzQarF9oqnzmgbB7tWcK1PZaz1weLXDlHcsK4Kuvwn2bgzLPlz2JxwZhMIZdXtq1FrDN6k4ov
hmmZ7QoEQnbeSWGV//dd806pd3k0WQw2zPd6c+aGay0A35wz1t92wfkuBy+QItyKtZekoG/R1pLS
gI5GrLYSxZ3Pb+hJeBh0Kv8QAvww0qNXoeVWYFQCh0aPw8wH1sUqSVsGQI506flyaBuEnNtleTtO
lbW4FuJNT9zrwmYVYOLvNEkzAGB/bgSUfX6n4xQ92rhvL1ZOMfyZ+w2lut/xuHN9YkgeIgGTVCzZ
kqaPzH1lwpIO/Qx/CKzLFQ60sBkmI/vTFT43ENJyxNxHwGJ9zTS8w7S/Of03HzQWAx7fBgKrLhuK
CFd0ig8rXn44vfBq2yfKDJhcqOufzSk9IGJbKTpHA+nii5dDoZJxS5Y3l/IDYfNcPEZeFJ8l9a+m
HqMcofdxvOoTBbGA2hA/jf+Tcw/GD9VhsW1s8D+IEFpj1E1Yj4fjk1omYg7XEMHoLGlGga/tCrQQ
pnCTOO86zZxHHp9FnDe429JlAR+r92FyAusc0wkWVFmdbIWvg2CSrUMsJpWlPL4b65MurkauSMM7
rz1zqZuWwjnp1iGfaCJosHKirYnddXezXMP7J+U1MESasGG/gQnRxRJx1nkcjkJVi3kP2O8Ujw54
tODyohhhmPCSCWO8wQmJlckM50J14MKYOHeDO0KuaXfLA/6Ce0imxRr4lWOoKgV82xq3pe96/jzx
Ge5gC7AbgB4LBHZOEyi/q+gO6oWoxNbEioTnSyci20j+/WSwDnIDFiVtJHDp7zyFjUm4HyH+Zcrq
GCv3WvreahfdOtq/IFMnbobcuMgcrBd8YcbckwojVmmnvOZ4mVWQfPO2qkUBOa+LvrwybpUNeURk
wzhrOe++12viwB7+x8GlsqS+Q3qx89d4Q4EadAKqSEPuJ/GH8ci5L2InmSqntfXcJaCNsSSxYknj
XOdy7g2Hc2+DUe/oOZCT6UikjIZScklyymYEduY+iT0xYmqryYZdTcsWKtQLL+ep8i817VxcB8V4
CI/QiPRrp9QLnMiQY2uXkvqd7R6jCyzespTpmsiFn94Sz3SnC3MGIZZa3uAbB4r3vwW8pDUI4gSh
hQqo0gYdrltziUDX9tC7G3VYouZanmbCIB+j7LwtsHST/3GrHKS+HIN64tw2dqv36+5PFZvD61Of
zEUUyliD2x97qo460sOSAbCf5b2xX3+wMJJVvEUdZ55dtkDQ2j9Ik6N5uvsOej8Tg3ABfOT893Pa
qbmzHRddBF/bt8/pfbjkm4BXALQMqTyt1VUSbEMkx1FEGUDIBvJCTAvCyX7zDra8pM600FGQW4QM
sEuw0WR3yhmnynHm2LhFmgY7CrnTmJiArN3eo2nMi3Waq5RXM3ed6z3pp1ISICO/Uuar6J3F+fJV
1psD/Igg5EPE0BUx3r7T/JDcyQsutkMC4tFjQjjK+Pn4M6TizLswRC3ADjp3cQn1L6Iu/A6ccFfm
979N1IYJcq/uP88HQytjtaAVMnA89A0BzKjck2IRx43GtJA8Mscu3ncZXXbFEF7/RCFxsdjrIoFd
+iBHeiuggJ/X0A2aHp8cFXQlGfO98CmROe0F8bYFevjeUDr0HxRiwnsC7fsxP1zpJqAokXYFpBJV
o74rJx9NnDxhN5wjZqxXE784qRmxSKmZbuSx/qoSeDsuXOETpT8RVRjE8ynmd2aen3vPKQBzY2yh
iIqv4E0CeKfIyaw4spZfUQY9B5X6eFrNI92m5Azj2/ZRZgDiNYxEjpft3rbKqd5Uz9/Z3pUk5y53
a8D4wasyQR+J24cGGx/2eQj2GuYr/llr23cpeCC/QLx5buBRC6SQSe7FT3keisKMo2CdvmqOIIWQ
tbnyXkiahJf9Y/02is/gsSOgOQfWZbB3HOUvupVQLhmKYLL1+M9KVx1K4pKVThjyxbpPCJJdwOy9
c8H0HzmGPrxEA7t92HG9isKiVr6dEcKknESDTuo5fcnrpXUfnMHX8RJCgtH8GrjAk0emCQPmwCst
Igg4uqEv5pdXl/QtXirmAu9rG12X7Hc6TTdp9mYQWAeGeAUnGFOQnQgIlqULaO0ezyJgRIIcjVtZ
BsiYLcrYmbpRzg4dEyLA2fITy482oE78N6JzL8ZZP4DqQ+MRIup7tNhxKWzaioaXZ3XqCYoS/F1+
nPb11mRSRmzzJE8dXBKaDdeUoVw83B4D1APkZimH+wpEzjLBJ8brtf67f2+BNXgJx0jg78r05V6v
fSzFfD7QpYF2QBOOILLYDU8ParqHFbuu3Qk1i/Pc/FKa6mQ07QHTZlFc3Eb0PFjZJsjqxzMd4ltt
m2jnsLQPPXYvwsBgdSqJwci7+FbBq3kDtJvWuoNEwEDGoSjdFIjwtgAUe+R9qxLI1VHt4U5iqioM
aEjOGyOy+gDyhkfa8hj14fS631tLrvFu5ZutluQHjNPR9E6WPEH6WOgzTdzfzF5/c1rAuDhkET12
I/s7XCnX8MVbCHoCS+ul4qckNdVZ+SAcq8SH+4nMYMxOy44Ebegzu3Z7iKy33ALBOQoxEumD2h5H
JDD2ueOGZZp8rZ5yWN5gGuKoVCp2TNbjai8t1uo9+L5FrUUs41CGTyOkrbwM2fEMIdUyL0XFeeEH
nmQPOQCpzn6zt+SRPxhrYkBWLeZ9Xc2oTuTTI/iUNjwbea/OvsgVutHtgy70m4+o694K0etDj1FG
xv0vCt7ahqAb/IbKMc5UpjlD4iuGeMjy0kMJB8a8l8uM3mV53jLT6IbKIqX8Xu4aHAT2ecQTXcvG
lL8+q9+Og0+zcUDD53WRiyDAzreZD1E6mVx09Ypqz5f95+3MxPcNj2FQ+4am1X3Xg4bV9gvRJdmp
F7kBKA0Ij8UuHt38TNBm4AD9M29B9dfTwNtL/wdnOGJRU6adcVbXjN4y6kI7nGsr8AYPAtq+ktFP
YrCSCX7mZ2YpIiIJaSEJvtw5mi+NZkdNEiC9OJVZdudYLj5xDTVQxz0140+jsvCye6pt53LAc06V
ocht8lInTK/9vINyFCPxn1Bo+DOMvkh/7IyYdKh3N5aahP+FvzXQ1TqHu4sobnafEmPtzZojdJE7
esPC/rga5AlhQkCqsgpVzAONzeUjAg68LMjjadQiOpD1PS6Srowbb0BxIknojqhSZlTaCiR2Wa7N
YgJ7iXX0eO3XeHP7xvj/imZHbvtcfm74lbFGtHuLECLt67yEJkPMsqpe1Msms81SDNQS6KD5CIj8
e/9LEVs8PdsjES6pYqIYeiSg75zu0INvORBXyr2XgBS1fnhSQVqQk1ABu9176kyeLEI3sM6OYWf5
P+cJjNaSNdS0dRs7cf6Qmy1qzwk468/DAQlciHJIdRx2ABk3OR1W3P3xnEMLaX4s+jzRFp8kAz13
h2GRp/8fLEcE6M/HD7d3k+XbEDW3wrAy2Lb2jrPxdrSqQBWgoE8JZE1KMzfeKjnX51p91/IcRUZk
cmrxU00dAKyWp9uX7T6BzE82nugcG0MJRHdDS90xV8MBKnasvvqemddAjZUv7noll4nbGnI3HzOt
ly/Lv+SBw3Osz2GXt5k9pbl8T9oiRaQZqbfTPjK6bFIqj6LUGUyCWO9YGlfp82AMcf+7aljiJUKs
57PnYDQ0vF7OIGHVzJtLCsP8q004hYBv2aNd4FnvXyPAP7EqOCH6vZK31Xa+Ijiq752PVLUB0ln4
W0RfY7vgdhtzlCTpc41jgxMy8YB7f5Pdk46g5QQ245KS+mXc0XvYTTdlVtseDeNhrg+HA+IVo4Vg
z5KxawWDktPtJ1ljK+1eJZCkruD2DJOyqxF49E0A2WaaGzB4goDP5gq0dbyM0FSQ6y/G+3SxknMn
2bBZQcTnsxClMzleYASA0CPUhzRd/nK0HG74aNivlWzvIQ2S9mwcLYUHZsvf+sacIJ6OCrqFifcR
x/9fdrB0xO5BtUwdi0V0msuWGsn5GDi2zhyWiv2ODwAN/mrW6A5DfHA7+jMBhU9YNk0H19VmYjLG
rHlbL4VrFTK3JAjux0pdhV9jZO0lVt0J3Aawx/ejDoJbjMnq9qBmLndywXT0XP87ylBWfUBxAt/r
hqwiXwYaKz6cGbox96VQBR3OC7XIC16X0nb59gfVd41Jaz1BgLfqjrPgO5b5qFePgLnASqlQlbZk
ce+Yr5lRjzVjRTfPhneyFF0+7hTXA1s373q6CiEF7qpThe8LvQL9kmG07hdWInjeyHupeB/tzAk1
LzY3CeZbo/4ZO5uEKuaBpJ5krCB3G3A/rg5ewWQYKJNGO2G6D424o+Cf1UWbpoOtqCR4L4q4+0To
K6W5KUf4rlC0cpGBujoRhKahVav0qIq3J03HBKvr4KDLxAU8kIaH5AQq+cUFeLoldOxO1IEDAylT
mGGyAUsQsJqfmyzQoDJwDp2fBBXw1j2GglCdVSAShxl2l9a7xYbVoGBPuj51jJgpjTYtpIpmp7UE
oYhFGn40ZpB/8rEjIcGSoNcZn5mEBPq20v3cT9cUEtcUDGNwtVbtaCv56A4kN4gkSx3HT1UhKsz5
TQ1BC+UI21Ds4EnX6yaJdlAXSS1E/WrtqkWPsziikTd+NPpWQwilW7OBV2yUZzW9dL/N7lm2pVBo
MCNYQlMqa5D13GlrIwRpfq/1LvSl5lMHJX6jv0isDuYpWimxL7RIGu5whp3vqiwSoZYdZ821qxHc
SyeZtwJta8I/+qIKFwWsFgicFi9dlHIExLjz3fQR1j1JZkhH+m70Jf50us4ljtw6v9Qe79XPAzw6
vKJgIXziJMJgy7zRVmPcOUPz6QrSi1qD2aH7FlqPQkjEogeTlkujBRtDsioXWYZJ37aPV5RM1m7z
r9Z3IpY1tZxwgqdU4R+DiLJBefXE+NRjQ7Ts0wvDvJ2lE/PYgPaTyFJRKQM/Ixh6FAqxHitmQgMj
9WQhpB1K7alEoA2hZCaQsFJWOwlwnA9sLAU0KJpau7TEVCP8wrIWS7rHWGO9OmIBagRFabTj9jXJ
LYSfKRAMZImb9LbtXmlptpY7IphHgf5FDNNs1n/5TPTqk6Ug23lGqsQH8XJcs+JOT2CwVl9yLLJ2
YJzJx8XVpP+Ui0rQTXsaM4AeFVjIcBGzdQZFBDpzZUT3AMeyQB6i0p3lh/vRQ1b2Gu63ar5ln6GA
Mfg6psFHFYEMniZTTiY2ngnw33pNA/9Si8OTpSpO6H9uvQ/2x1rphjJ/DL/TbtADIZK4jJoPHcm3
VcKAdksCINh/p/mjVpQdKPegh62uJURj/9ecLgbKMX947cdnfIlhQhmKFzXlD2dghprWQUmFhNI5
HDeAcCkv7xkq8qzxIddXKrgOsnfkBIgmQTSJWEVEau88LtO68SrljQ1AFikGM+TUHIOJVhPQJaf/
Ic3O6qn2I2XBWyWzKps2foh3I9ikx7t4LrlALk1jmvBWhg7CgnooW3D9OJHK3Q2HR94YNYTjBris
4QZsyevyJl+tH7+mqMmkzwl/3hwcSYrXnlQs6LxeDfUNbfgZC2bldHwkIOW6d2kLce3ffO4HYKJ2
v8/y/GPTK/oT35VZJtOTSpRKKpyGiViVYYLuia/RUS5PRR3m91iqYRYVo2hZr7axIlYJJO936/DZ
MK0QQ5INMLEmde1Sfl9cTRNtJ5DeRl4e/fUUcaMbWg/920IP4KynslldVIKSafHE58APaGj9xREZ
xhSYLt1mBCEGg2EyE9mIT3fArcT6O26dWDLIjm2pk/k+ZdSlmf6hWOjF8HqZl18FtjC38+IoMCj1
gJaUW13HVJD+oAM8kMY+AmSloJPHMEmRugdYDxL4VogXq4+rcs2gAeOEz0eJniNhehwjm44lGuiY
og5WuXhaoUFrgywI2ZW7UWQVN71iXwLj1zMcqdWldBEuJ5YQPBx0wF1Q1EGMAICGCRV8czN7VPjD
xaKCeSqrxFzznw3K8nqyAckvZ4zvymhbLywEkQN0q4pxZg7VLZP/5QAFpWREaJiBKzgLkhBmCMUD
0/tiXhGgcUV83rgG4imgu85WvgcJ8jkZqokcJUjFyOJBXnb2z7fb/eJyjbTmCoJ94qvEaNZXh6Cv
ZJIwn92J8OgPHzhae/Txoo/hHd6b6v6l1n5gce3DQfhPgyfC1eegEebFBlBw7ixB0i/iDgOooa2x
7QkeGFEtBtjTt3bByIcqOaYdcWnB0CNUnvSS/uZc3OaDhMCIBhjks76SxL1xpXKSjQk61F+TOcWw
e38ckRD33joQf3Kx/ZlP14IGzaleY5zYVsafzdgIOuSYdYilRito/W+Nb8Cjjjhvz+VMEK5jOz9Y
5nvJHwWLJUdfOnyi58ea6MKgi66ZD3JBP0k222dIDCMIyPKK/k8+Y5a6/BxmY9Dw0xSh05x90igg
YPHM+kW7oEsFnmfGaqA/AKO1nqUA2Re1tFkUIEeQn96QHWZ8cGAVzL6sAZU3QYOsWU3c6JEb6192
IwlVC3I3wfM4VdGra27HTb2S+CO/kVX2du/dAvd8XKuJEWAmPbj5o3HEQObddvKWeJFxPRKBuSP5
UIISwD/4E8BucVPc8GCApp4Td/7ZA7AalPNfVATB9VbYWrWqAXJeiOY86G+xUczhWS1o3Jf80APL
9rMdbtwRjebtktHfCHJxC2eEyJRMSx8glIKdKTmhLK0KmPPOZAvqlwmSxAAP2CFtsE+EM1iMVrjQ
eEePK48ItjfmhGUuwzmPJnj0j51kvX9MJV4c5AUl3yPrtG8Idwy4sqJldvkILJp2vm5eULF+Y9uX
ir4nmkoAbWx4HAjJFMp3exneXIPJ/zKqiNh0bBkYH0C/PR+DboGx8OZj0EVWBDO4Ku5nyH5i3mq/
omVRUQJAMQgbhVfb6utheTbcfAzVR2bJXoR0QAqBAGbRPE3vu/a2ZCtSMw3CMeWsEb/x897/73K6
n/VaneBivTuq0oQ4da4H7IBciaJ3x7ZckhnN3ZHjW899n95LYsOP6xLtuzxan/j3zK4MQ//rEq8Y
xxo4YZ2g98asimCOzrBr00XVX/4k+6Q2lhNmcRXgQmQCopKqkukdM6mvBCGjMOY2AcbMrrMbkHWq
OJNBnZ0Plu2zvb2KjwL2HV2Hg2rsTO4wb46wHcN7v5bnxwaOw1shX2HHR+plBVuiLRdEwsYl6bLA
KOBLTAdLuVTG/hsMs9HPfFAoaid2ilLe0OUaSh4Kl4w14Zrt06yFF5Y4hXUMuOg2+FSu9ovBRLin
W6GD/eMd8Ltf4vy7+CqcKRR3Mk3Sl30XX2Mrxa/lzXryXMUP76U9DpmseVZvE0kbVOjMj/MBJSG/
AJNpMlpB1BzHOo05hWmkimW1n8Y3Ws9PMI1u+/qf30D94bg/SoGXyKBdhvVKVjVkmxGBYkvSRRgb
7guXSMQ6TO5j5FxXRvuS/agbc63l6nWBr3fArRgNgzN50hDuIYVmatHycVP9kMSeqfMbcMm/dqi2
wzixSIXktnbXYNTh6+Utqv4vL0Ib2YLJzMm2HPz6/nB1kA+YfUeBIScY+BP+TGFk6OqRYU2LSt2f
WDVgDb0gn9MwT7Acdh970DaOnhVj7x9+UblIburG9x7VkL6t9qPoUIMJYOsvBAsd606q6GTVwAD4
Ubupgl7zrgtFfxvcOLEAfWXFMIqKLWr4pbWgbw+JHQWPqYClnK9sGLXAeJF3qSyzNl+oYb1BRnFo
/EOzzSIfIzpTi0vk4rzhYbB561XrwX5VT/X9MDEeywNyXLnJ0Uxq2VipdY7fyc2vkbfQh4F3/jbw
nCGyMcswAqxeEIYRIbrlvvGnmgqGNP6t+0VSXur5ZinRaxXmYCeCwHqsd7Pjud/4c9l6namMNgHb
HwXd2sMTyLCD2PJaWHMkJh1BzObfLHZ1QWqR5ItDFuyUIy+UNse+JWLKANw6LnvWQv2Kne/csyWa
WPK2e4o3IQoBXU/P8W4iCbVjtHo0s7FKCmAWg/qhTR9AUD4frph134qy0eXQzwIHlCfZn882Uafw
5kPS/JTr810akeYOZ/SW0c3u+fZf4fxlO+NDhfQ8aAVqX/qEMb8GIPuj1GcciZVe+EM6vsur6tty
ZtWH4yefuhcOfCo+K2qVJy47IqYIWy4xY3g8lUuBiOiiSmptBNqpX+sIjZU5a+NN4FejKIkkyTD5
umD2Oo/6SC+e8/+/p5AFORUV0Gj925RLSCgE/EZCvILVwP0am7un9BZ//17EFYtOq2m8NBAJr2yx
TGZZqPIhmoJDdscEHKw7aLt7o4s29jxrbA11/R4DM5Ym03sI6uVX/TbcJBbzcrCcIoZjYVw9gzo+
N6Z0Clzj72Iivhxq2ASxoTZ72yJCobc97ygih5quskIGGx9AH31MtCDCK5JNq9tLH6BUbIlN5AmS
9fDeA0NOewqc0V/1QlFkk6rBngUQMGsp9Ap9yH3PSr3DnPnxnSV9q4VSp6v4evoZ/b2sjY0pVqXc
yr7O2ObAjbjxxx2leeACcC3/Imk9Jc2kYCwvanQI61N4oPwn6XcVtdhCkmeLIG8Tn2QyPuKhGKN2
vlwC/06qSR0cEOc885qlBIxq/wGEEsMmN3H4KCH67QTs2z3vbZXkGnHxzIcAjmUUqkhNbEoCU4U8
JU4ryOxBGjmh9bBRzvkrGhbmrgCO0FHfQfG/RsQ2/0KzR3lqV8wuDdGtQujNXJ23NGVnhM8Zmigg
55TEdY/U+22mpMQLSsQu2iLgB9AYO7s6KOARlLgcwMJymRiGYzzmYwc2MKXmUKCOXmXwnYk0AfLr
8DRq0d6l3SzCr+IstLIGWsi4ryrsfDyq2HY1/eVUhoXaSJJyxSwSXs5JHaxuwIJ4ZyG9vEeQUh+i
7Cfh9IGgyA7/jKpbVogP8cVmIM720lwS3h3MFU4xT2tqj30Lpp/7oKAhb874wuPcmoZBYbcjvxce
W7NK7foue2YR7UXCcqAkON96iWd3SPLzsX4eaQGPtKsF8Iv4dtNOkq9vW+bXHj0zB9Q9Leo6ER+s
O71kB68MVUumDqtanQcdmgA3ZIFhfLc74OINDE4wC8LFpli0EXjcwHdjTd0F64cAfer0UNfKPx/d
LKeZyndnJBEOa8Fb3DYOlVvzJwL7LsRdHEdMi7mGtNv2HgSL/RIsYKsM5yDmCriAY6g4/OIasPWP
z12Nbknc81/nZScbPu4nwKys7MXGh7oem9NSBSDd6FqMfM0epX8WK8yrpvRZ517L43D4150JSyPc
LcFDgZeFz4g7Z31yaOibv3qUH4MEEHExnpvRLIuXHRLnfbZX5glGrDPKS1PHHUL3VWQBWIhE74gb
B12+w0es1htKtscEnmkXyF9UmToH3sqxBYiE3aIN97HtvV3tWPDjdVlJWxmG4Z5dOdLQXqYmEiCM
han2zmVNoVwoi30UbIX8XFYApTPtdS/5GnmLCjqYE/2ZT5e9jNSlvviOfv54z+kaUVtiGcUX6YFV
lnJwzqXIQjSxe2kE4RM6D5qbZOIWiqXQF/NpUOEIQszk3c7C+L3atW6rtvcs17BQ8cMn/ZKNRHLD
cPHk/IbzTzv4htxCvzf3JOnqw74dIezBQ0VUs9CMCK7pjVpkONDXwkBlNqiqY0JPcpm+A6nFh0Ak
Emy5AIzM37wzMAqVgIJNOE+p5/JLYn+7OrZ0ZVeufZkgYOx5Lx8i5lojcxCyB314pKQn+7cg2MX1
Hz16MkLOt+H+T3JRNOR2vSTL9h+4PTO9YWvalpl8oFmJ4p3JxhocPdMgPRr1kaeOmBSj8FH2kIS/
/PhaHVHdSVI1VvUpZ6SECOiBZnSu+4ZXVIiCoQcyLasFaq7bQSAlb4XLasbpdxjPPL0p7a5MLkB+
/jIa9pR/sWd4zyX2ohc2Ybavv+CPWfMJnNXUZ/+CY7daNlvX6hxxhGBqfqnCtli5VajZLBTdxRD0
RxC0cg602tofktswsZbtG9R9HiUBbx/JdsJBOJhdCd86RnEzsvGUR0UIFpsDpelhwiFFWXPdkMb3
34iQz2Lds+Alykt9fM2tgpD75SbdiVKmXXcRxICHf+TFq2K+3e1wJPSrcHRUBOo/IR5LIJtlI4l4
N2qxLvcsf6UwSDyIqwd5Mq/A0FBnguc3bC5kpj8VP8XXpF6cjX6jWpCcFgi89VFi3hDlo1LIrOOQ
+wWJDdibKmpodqEBaCm1Le3DBNDdidJElyNTXV6+vwRagaMwrprrMDh3zM46jMqp0thfqApByvxp
OIhPmAS9+NYh6Kv1ZMJM26McPtwcxFW3Q9oIOiXQ6+f8Xtdnr7DHcfl4/7QAp8deP16QWYofeEbv
E0R2CQt8Zny35ahKOyRJwah+RTXmHJTtHVETP4ayQlnjoat5dWEcd3jKxBvUzmIM/NBF5aepK+F7
95kqBNHQMzICt0Bp5ZWuYDHiGpZEE5Y4LH1/0jbd0Hrk8wwyZgFAzmiJ2Ob//j9aYYqa9Vgi5JcQ
6SZQxsCYqOsbHIhyf9StV37w5W4kvdyrs4UvpOdE1r6gTyeAxfL5Pk0yxa5tq4+lFHQkxE6znLDi
r0ocKEXaIqa2Mc4VKt8GbWaRE15SLMoALtx0nkq4s8F57LjTTCBi50UdjAjfkZ07IxLVW0H7iFWR
b47IAufxssXyEbF7p5LnNCQue+XiVYNSxc7bp6Iq8fMEj4FDz/zcBZVNw1ohipDVxfnaNdgw6KXY
mFmuHzTZPdcdX4+aGTAWR9cXqT7RTIiO6HCYo5j/wqpuNDGUABV4g4mC9XhVKEtIzAQm1WrnhOGG
ZROonQ6bzaqs9pYZb2+aYWVK4qw+Zpfcv9J5c2+l03ZaNyaeQl/Coz/heuq+BTBAGI7pnzzFJ1wW
nu4CUcD9afq0lDPYm781nTozPFjrdscm70sJZ2Z67t7sgComg254f1Ywdyvg/iP08MmRCwFyLbsa
8jakgMRC+walIe5aEJU5d35i2jMah7BjYfpeBybcUoJkiJDzCmEMEMfvt3jQ7Zzpn80QI4C8zeyr
WU70ZJmmWnh8f2JkIz0LnFRfI3ccDxpMdz6+DL1+YiRU9FIdqMu4j68TmYQOfQzI4KaO7FYKnZKY
m21rkg/YO0t3eT2bBDKVdE7xy2ah+f5IwsdJhi8D/NNelgKNXKRDEUl54EoIFkzr26e4+87mW3uA
rJdeXW3wPysYaIrW/S/isZyNM5fXNn/AXG+t+Sb29YnabR+VR6p2kZdgNoBufGxOBoHYC0hB3pLt
D/fkkCIXAWgHs/6bEIBj5wSEGi9hpGsXpyDaF525kWPLPOkTdrBLrKOxjGY0iAcuZL/E5whuhXxa
SfSYq30gOtJY+TQGBTcZL0d4yjuyJV5xtDy8qLqDpgzj6G/iJYMNnprF5QdEDiwgiQGy4rQRlc8c
QC1VgLI2s/HOqgk4in+Wiu506Q1tpj+ASgxE5AGC3rsvSO15GeevwSr9xoHmE8/Hm7BVWVaoWwWD
jy2iM4KLVXvLNnHwCgY3R4xAd0YMpE1K7g1Ufk5ImUzBiqZm7Pk/+/Psk/r3FaiTBbhKLDJ2qLHe
mfaesATjpfhlpfxLRPDAW83I/L4c+HJtGKgXDCY39yHkf4Hg6qmNxfDSouDX5aj6ih2xzeLyxExq
OdT2Nv349JlwFa6XXHozv/neUKlpnVN868d4dAl8KLHKniSP3itikk9n0jnaVXRNbR68vjrV5rH6
gyMeh2L8KSxdGkqGDfwpZSK905P7YVqBYZaTacnoYi3GGMuPAaMppVQoYrU+SY4rfe54/dr17tjk
QXCZulYyJlz2AriScWzU3nHs4eCX4Y5XZ1P0eQc0pn0k07fUtdwrvPL7J0gL+Kl05YA5RD+65IF+
O293sM6QKPv4RAjvuVFk0CVdfyCzbVCHhVgYW+a8bZxKEBeGqOlli0I4FwA+fKuY+eP7UmHR2fFa
GTkXiFCoC+YM3ATRnriHwyNNRu9AEGSTOhwBnEgVvT/LHj7XHp3vwRXbLfExeo3+aeLvy9NujNbF
aRNWsHn5ZwOY7qQQ9vMvOaOVmHAInkNfOR3RGSh9dM3yIg8MA9bP8EDqghotJZKi5g/CaLaQMrDY
2n3sr1sCLfeYmlphw6VN5mYjYf3BMIxFUbBEd2I28mzfKryHZ4hShN0Xz4PcGdYIzl5mRHvm7zh5
Bv9g8DqEhGyrhNQgTqOHzDYTKql1FVUkbI7fUV1Vh+f44KhE9Inc3s4X+SPgnUYPHABE71c1qXqU
3y8azwBHWQC0zJXp3b91RH/8+4pB72aecmy80hYZwdK3Ip0ikVM7QXhPahXg6pB6kKP2HrQiVWf9
p+c8szUaA1IyF5I3QJegwyfmp/vKK9KBAw4gSXoHgtmqw0FiN07qPKDO43NOA4O+Mfpd6jbk09MI
o4+sFWlIZ63rstsLC00kyqQkQe3kNqw0dEIvh/TdtvBCJLoEPXqJGwPM6dpFJpF1hoY/mRC/ionT
guwo7Ti7Lnclf+cuGJRHzAEtEYiFDior2xUB8/HqkImvaVuEVvMCBTjFIbkhyo+YXet7pOXUfUvm
HRyMBFZ52DKOFaFNIAb3hasuzPlOZZnVpmXi4So3TkYPVUrhosu8mGxGXLug39SWp2wMYFDAJ/Zg
9m8uCbZ3PwqeA9I8Ln1GNaCGN325ElleRrJZS2sjAnW85DtW8f2zpA1hQ8AcL9OfuHhARAxniycg
LVfn4/rbBYhXEclJ5IKvoyj4c9M+t2IuIt5Hxe2gA2s1tPbISJEz1iad7UB7Hw8gklegxT4jI4sT
wBqgO9vUANYfzMpn+yNbnPxriaSmJ8YOFXR3+WQ3SNpqqaIy1gyj186zx+lRiCyxN5JFRtflA04b
Y+NXNtNm39Od9HUvpVsHCb6rNO+c4rMH8pqPUJKGu9E1csovbyczPNwhgZAAUdA/ZxCL7DxVZnoq
60/Ag0LSq/0sQghSFH0CANfJEIqMPdM0zehLDsPPpPlDMrB64VmJJLXRolB0d8gJdLWiedWIdZYb
8ad94zr1DPdAsdnn11Qcvvt7k+Ems6qHXpI7toO2HsgcHLw0QZndUqVlDWuS4F3nwNIrK7rp2dv/
KduvCnDC6qNfrs1BYK8zR1pqAUsPgVDDzWPN+bKaNj6AoL8Flwy4MVQZifenHtsyU8qVYyV2rA9x
0Kpw1uIr/vVW/tyQkpB3oLIRVZymTmbhj9QX6Gk2SCQKlA2ZkV11ZHmPBPkRZhUvIQziIszX+5lP
Dt0AmXMxsil2GAc181O+YSOS8kAr4GmokYVo7HsBzu5eSYIWfGIY2fACP4EDageGEPPaGcSPrBg/
58ghlobt+q+pi76N1VHT6L3SbT9bvuPVcWps8EnGjdOOaONGeMudl3Il1zM+m43oXq1rYSe1aDKk
8MTXavRrvmWICcBL/9sC0V968fMEZKGfMDYVeU/+rmnfW3S9XmAyQGhe1m0NB9qPmMaG2SZrwjuw
Baq/ba9fBSZ7RY4/CQ4awpfBtV6+Tk31UZEXDvR3pgw28e8TYqBrFfMwO0Rp3SSnvpMEsW+0M7De
+iAqfa2EHCvdIsri4T+gyhu7XPPFPCyBPMRm2Ii4GPxTXV/rp/4r1urGYnsXnkEq4OTQNJ3hvPEN
a7TGxlRbhv8Sj536h8T9Dt+WtarkkaEs90niUqjZ8IhDr+D0X8oIF6RLJk0kSNsdWWFbHLTL2QSI
KcU+Xf0LsMBhbRC+O2fz23RhOkUTZ1O6dxUkeCZHte6Et0wB5cVXwO1JyMvu16RhvU18QaEf24Ma
bhHtrv3ZYXZc+ms8OSw/qrHlOHVBfo7phy04sUtECmLAK5OpURHDcbxbwffuWwET21X//Rt8iLCD
7JsLd13CrT2j2foAo5m1NXrX7W30tOy2E6kVcP8F9NZwZQOHUBJC2M6l/7UwisRqPU2WWL5iEo8u
6EiyvBwb3sZU5JIWvsfBLcU7YkDM63I1zAp2k677aUkUleeCDYJc8fJ3aLsDyZeEiQc3HP+AJRux
dqOMNhtUPDPssgGBIEcenx9l/oaOtBNhGQIZw3GQJMcEXhQYjZAhAJeaTmMCOMbpe7Zgsyt2TK4r
vYlxIe0KHeO+8I6Y/gLQycs/6+AqZqsiV0gMPQTEHAKt3OaBgjXpj6+dGlArFm/sCZDQWjrb4ByF
nJO2CkQ5Vsxdtj2fGYr4T9Kxv8eSMGVVdwHGQpAqVPgYi/Sa6h+rTi6zn1TnRPnrmMTy70KRAgfA
sKDiM3st5/EV5SkoO1kJPOI+Gnd5yDhlUk183+AwhmbtgCBZWTMoClQ+ukhbFRrtfRjn691qe8yv
5zs0oPSjqE8v1srj3HfDDUyf+v4eoB3E4IK+BI6i3RJlGVdoUMG6wmUlQnK23YmguqeY+YX98LRP
sOxuo9AE7lNP1srxXAW+lydqk6pVHRaLYrTTNS7YYpHP06nXldtrvjOpClD25j7uYg57yMCFFhXX
yLkWM4anKfiyEeW8c+9MH8d3C+4sGDoSj3RQCs+MKpkNYkCwkQ+joH0R5nsnP7+BKKVVOAhQv56I
PhG4PyZ5CLDzzLynFWwFN9LCgVqNehOHqS8qga5e+WBjQHKq7amYoVWDmCVVeF1YC/4CvBUDGGN4
sbd/57GlN1EeM5fTgCmHQwk/u45H66pqCXd5VuRD3/PG8sgZBRGVwS92vo4UnWZ2e0ucMbxh1HrD
eE+kMZ8TwgIDp+LL9bFTAMk83cchjB9T48H2HlTrfrhx4kabqWuixIHv/U9AccXKVzjS7+exTKgr
noPMECfJpH3nh5FmUzvYv2dfbSGXQMC7fk9vUoiwfq9rmSZrMsDitcSPeaYaA45tCMr9Fpf5T/kP
23xWj5z20t/B6jTLq322emte7woS9gb91ZcZq74L8+qhHhju5OfZojknJ5AmroGlLlHqd0uusYpy
HV9hDM0suVt+WokY74+QUSK0NYdt16nrt5K95vPj63Sfv7Di3c3mqNUcAWDDvBXB23cwpxNAXXGe
zhjaJdb64iJ4eGvC/DTvI+uNyDOdHTL7i3pqfGv0K6FuuTv7E9f8ob1YuJGtNNpX9bSKJgKpOrpP
+liGgvoZoZbrxv2JoMTSdZ4VC2osjpo2lIOLzAjhB8fJwL3lO/9RjfPhdXK5dEHCa2SNsYkqZMbc
2bFqf1J1SU9JXHeyPboIxOXCoVOsCBzCvV1sHDrlf59MYn1oNAVKwJqxhuwW9acIYk6mtXsD9CVa
dAVpPEOCE//oFewvM41/JR9Cpv3nq5eY8anbD/W1Psm+2bE8yi24w6UQlSGfNXaFRuJbc2xBf5yW
lNfxPcLv/3P72r0NPj22K6oluLFwfwo+gG9TIVeUICS38m7EPoOuQ2MIGSg+jdwlGJ/hqKuN/bOj
kJgW4el5Wr0/u1l+4Cw9S6j8/VYigy0rtWOL0keJpwJUN4tb287E5VE3TN8hCMU0QTr1wE3xDMzW
Lf3x2q4ZwIgXA00TQlBtXNxnqK6x4lOakMBqnHraHXRMNrYaNvJwNQswIMx9nStEMgKuyFgjT43b
FyGmyGSI7fTz2YPqOo8VvOvzfB7wt7PeSlvqs6BB16y0fL3ENXyqSqEgCQmPOsfx7Fo1aRymz5Se
MJSGUnJv/c2H6JZf1xp3YpPEQKctieZCTM18fG2pDOVBmDR6WbnipqsjDsqE8CEz26V2ewpbUyHs
Yb7ptfqfIFfEBaFMzTtZYBaYL/Xro+8jBcHNFV1hh7Sa86hP6iUrKq4Qm4TbKG/HQqHPdvVNdXwi
BSwCQPj0o3HEOuEsZyCObRPSAD4bHnNlqg/vV5Caw/SXJNU93xAbsDas70aOsGN56k44uJhH4Avm
YQYfYA4fctGDTFwVEkhhYfYFORAPnYY4ijYcdfN7ppxm5/5I5lnqSLa3+t0Snc1IhfWy9k0GGeLb
a2s3XyZcYEgzITTRR7f7yRRBISsrGrozADSTUHfO/e841D4BSVkiLs3ME02b2OIBygo3mcjFaFLu
xCs9yctHK0ogrTzmTzHWdwOz034EDui3vYhxUkex0YCt1FYTLH/fKg6YU1rAcCUasciYBC92ASGm
8xNMRDzELwKGmW7ec4al0yAiHjXxYK3EWKcUXE8/RASLbO6Js1hQE2yNS/63nd1MSlSfgoet3Y3Y
T0RRKVwPQnStnyJtIJPHrOzFlQcctd2TZBwlTAvZ6Bmu+H14g/XgbfgRw5XSIOoLHzLzd0/eRiqI
Glo1sl6Iw1cZorWQGlEga5Ri2QVVE58HGeoIPAZ9dbqTc7FJqeQzGuoymc9uVeClxG7TVug6A/F0
9eIir4YItAWX0NoUiupfvJTA4SnL8BsXhOnrlJIjjaPHxeiERtNJMYrAEfV5f/7QMhRa/moO6dyx
XNV6s2Ph3hsRbclKB1vGw5zQFiSABRoOx9ez/2JivVL01yKiz+T3BsUUofJSqw2VDYV3PURSK08+
FVt5X6HGKNYXcGzNCCxpqrXnlB7CI5bYTV1p42m1gNm2IYUXeEGYy3ipEhA10a5WCLDuGTFPMSxU
Y8KKAi3hoHQpA3ke4deuOE0zgySIENyEab9Vx67217ZYsvA/s60HttdflEykWT9ZGgIrU0F/0KCo
zIw6nC4ymjyxuCqHJ1pSSGCHbUf9FNECWkcQB5fB/scozGGYAzogCW6sdWCe9yMeJ3BHlpJSDlR+
NqglXmq91N4EiqMM03K3uMtO2aXHt0Xy3dCtJEMPjlR0sCA2vqYQvxeVQNmiijFM+22aG4ttsdgK
5m5GjhZgR/ElfvJ1X9AOJhmh38dnxSDfCs9kA2j8sHC1yq1sCjbpfgg6z1eC81ealvHXJ++OUQqy
xxJdeqTK2s5wTMbSfoNEoi6Fx5S9FCffdKu8JL7XFyITjua2OWO9Lq71iMywFYLThD9Kdh1syK15
DALlDmTmREnzXDZLFrcD0iNcbnbF2zuC1bzoES6Ysb5YDQVswD3FLq/RFI1iHEfD+GVu3vJ4+1Kn
76VTGayohtHfi3bqinTHKTWYwZn1YCTAvMq64R7uoYoX+cMHeQkm7tGt/FzBeTgXYTYS5xQO2MuT
ipqVXQS7gsJzkPhZuZ5f9bmwrO4GLWOMOWHaFo2xDXt+5Pmao+MiKeH+xAv7BtSU4bviLIaL8Cr9
jV1Bzt2yMdQkoozzVK6B11WljLDetb3OtOF9GNv7dSk2c43H80n+E/WkCv3Ri165BTWlXEZXccqf
sidIx4s68qT5/YKXPEkTKQ4k5I0OlQybQWQavAgqv9RJZu2D0XLlJ/BagZndbXFhnk16wsMt0VQ6
lv33WL8xSIffJp/9wTgyCi9zyxlfEVn48K/efdiJJcWad+vsF8lKSn5YClyt/DkAQ2SPYOHVDJvA
VThizXWATzuZS2lwoWozRoBzgR+VcaJOoF7fr+jbY/XPaJwQ6AwxF4iQ2uzcgfqWlXWhOl0JzWBk
nYqwSy4pUR0PdUjuxdF0oBQz+tHgLT9xOqKjdtPc/VldksPupMkNxm4OSEej1D09Tnz8lmZzirTP
gfr8LmRiGycMMsIgMzWFCw2DGMo63paFnSV+dKlMRV/1k3bycMsdbVLOPXwD0U6Z7UxzEt+HKi25
vkKOYHwTicgWoltjpzrT1gtxh1Xw8oKUjY4nsqhc3AkdSuinnYwbYfZNpqqCY9sAmSX9Hnzjg/6w
mFMTWD5NUir8Rtq21BW+oebKms7T0yTucldllfpHOs5wXxNvp/Mait3DPSl7ec937szKhslKA1pI
xfviRdlfzUYm415dFYIa6g88oL7N3TsptLegNDZwMxKP24k9MO5ia+Xj7Sw0R65Lah9TSjSnjIu1
UN5BBfW8oifnxgJNd1YTjGh/+x0eV9FjR530ikGzmMYzcZbi3vMgSVSK7c70IiaBpdFLjaz23IAF
SxcwsPv+AKDKHvymZMSOjiUZXrNyzJvEkiKhdoX47RBI9hfNjJ42NLlseXhaGfkosEwsnfvY9lPW
mmMqfiJ6vNAD9dHrnu2t6Z2V0TCmYg6pgkcbcpAtDexMEqK1mS/+hmYJ85j6xADpYaJcuC479YCo
Vm76TxUJt4fylIGpt2WFAtEqNFTFm4WMTJtjK5mZBnsbTxNvUBNhXZeshlWf7naTCHhw6zFUrdcR
WCgIfwLcdi+x+U9tZ+Kvi1CG3iYw8qpJLfIkM6a/sZaevyPMjKuUeNv5oMpgUC3BuEOgekNSdwzX
HmhkZi/+XWCLdsnAD7R0TUHwrEB24hntRKkLSZ8F0ruqcObQ2lAYoH2h8XPvIgZ1+9F2IK1+YVSS
ZNQu5kUnqnTCHd7s0eq517wQdxreVd8rpqgbJ2OxKAaUQSeQw83CuwHnvK71lZPeNSfSfxBip9n2
18peQyEyeDsb1QGFe2/7Iz2asIpfHyFYgrN0FC9rFd8HIZqOB68qrkNIqELhJgIisoeGrCKHqbqQ
WoCOOBvbwgltWiJRbUuGCzwI6UU86QPazkmeNIb0W1b0Qq5YJOnZZ74EXqZFYD+YtZkO76rgBfKO
/GozOrO+3RC0x3G7FkHZoxj5VzQIyJdhTMIfBLvzxUsuw+++B6+5Tn6EHeRrqqiG6PjEToogNnMH
/1CNtRg+4uzpu2X2RfpCbxQmW/ottqg4T7Ak9iq5yE5BZJ7FG/kV3B3JMh0bj3LFxt7pmnP+vmLY
Nssen7SuguEb6TQb+WU6iU9gBHElaLcy1UhxidxywNDu9xchkIuW2BZhGQvwT/Z9ELr2E9fHpbgQ
rTR0mjUXyI3HCvsxhqSU8KLTftrtVqs2APAXPWvOsEJX3T7ifYTQuK1KOFBpvg3rdYtWH0Yjxvi/
hFhCgGwCyCmgeCXT18vvGGJrG9C9u8Toya+QPeyDK7MqZ6wxl0IGAfz2/uiti9c9r+Xlm7YcSmuq
yXtAapEhWejWNiZngYwles/aNQYqnY8D22FN8t0kdqLN7vUvk8YWkwW+j8VoUKB6THdv37w8hSv0
RvoAbCHXY4GWmum8nqC7cjN5Ph5u4eKLW5LLLmC4EHJckF15O9rxRhzze+F+RAQMvf/yNul/dv+w
SLGZUQmJzABLPnqq9tsCdsnGXxHGVDoJ0WJSNTRjqDn9s2GIYPf0QUu9i6EPEqBnqY0sUw+wI91V
p54b1yAJMytmH3O0kaHAU2ucon3xJovRnScWBk9AkgCCbq8XbIv965X5VTqxgLRi6O5rl7V2MDFS
KZRYu4L5yr3+WpFNuYahnMPAHtHGkKLEbZzAuWQegVbDlGIGzZoXbl+n/ho8ffzL1rPzcvhI8dTV
Hxw8RtDLXwDs3MAqsB5L+0cgKidxOd5SIQrc4H9jqSr3eTXdFl5iKr+5fryg8Xz32vg0hyiMmQFV
a2Qn1aO9cWgyD9rORZ5whC6RWIyh3qG5+MgPAiSzM6k8hSp+PAl4+UEWuOjJxLi05xMV3B2HgQbp
H6lObFHs5PSpfj0qOagdEFdKUbgH6adE4osbMPdMEEoXYdCEZuK/I4Vaa/jRtfaX0k5IxqZwI2GR
LKD6ubBYw36TsfX48fgIqv7ylUvf9z5iu1fmDdfGgFhV1U+kYlwx6WbTRzCH3d8oEdarD/RUYTdh
4/f/Ccs5Ti/CXvZXcpaetj7STqRMFda2oSBz1kMAn0O4hoZUbAfG71V6Pet8dOHjcvH9y26cuyf3
5ypPfNjYt6gLuHm2ZUYfTlxWCsaabzpzE0e2EmtaGwGoD+CNNfOwIZvIp8fBX6NpmBvUr2MAzE6o
9Qrs+ECRQeOu6SMrLI158UWV0gXTHcPEM5tYI9oZN3fvUS7z+mwVoqcg/TeV99DVxjyvYVsHNVXe
OzWAo5AxGtRaZwGYXhuZCr7G6uivJj1v0iFUhOpns8HcJlUf//ONRfAPIFeVz04OUWIg2GtLDhOC
iLxNjF/rnHLslhP74Qa2vucm9MfjjaRVux+OAGEyPubOpVDA+bsX/f5Uhs4FShcwwhaoKQkciedd
Y+v3xtDFys4nsBS/qNbkG5AJ9pWCOtjyq+vPwcbLFq5W+oQQA2IUqRayUrYYEEAUeXXdro0XWLhI
Pb4s11qDbRttjy95IAxk3MeIgRs0hsE5EORg8rBdKrfz/XdFOzq5ryxWA5FSYBSchke/ZZEy5SqG
V6QBf0peyAl5JyfLlObZddVfOSFWTqN4ba9NxsOX0o1CP6pNx0ANVPKPWTeA10fSiXVOI5NGhevN
UB7Piv5iBTGCCzHMx69knuKK8CZpYbVavS2Z0Q+2XWDM7ZD+24Ba+Q3zQFZhCphqdlWZc7kiVBxr
hR2Yuiw/jKm+0KtG1ead35uG03bNpMWKmGfzJ3YAcgEy/gXlZQdpzS0dPKdLMCpdBsotZI8z6IHP
zLHGOW71z8TDnbDYtAtDseHvmCZTJ0189szXeWR07MMdXCZAFFv7ZFRylpuq0D5gEPuBX8h6JT71
g+/PeHzY6SfsojHZZeZtSFXApuuywJeYvdb/nhUDmP3t0StPdI6CNt9kWW+Ol/xPr1SALySNuG9a
38i8S5rCsTXiYdzOxhvwmwnLZX75AvhiOZsBFeCZeIwGC03b1X5Llk2DP/Dv74a/z3kEtJf0xd2T
q9ijLWy4HlYZgTWdG1ijWbz8nWW8vZOo8vfBpeA4JEWiXJkAcL+Tx3+JFoykfHp3qtT/yIqvs9Gi
oLaWa/3MEP1RF/F3erXPcCLdmcwlRHV5vbZCP7Ha7WidJ05zzSzRbvWGyzTcqDygGsEU5ftiEeIz
8LyQC3qWPTSFyAChkAK//wjO6l4F2eheYee4evble6IhzGh2qhmDJYJh32RZh4d9cowrCQx/PVcn
H+qzDhoo3E7pAhGG20ZuGgfJ9NErhHC7wrIvTb3M+7QF7NbSBZntSO/PndMZENtxABYvdHtkHRAR
ue0dBGoPSHOuyb6LiKjqfX476tpNulT9Eqe27exz35TVxv/DbCUxDObDJzxmJNDVFlA98ODb2lHP
Lm2dbPWiVEpVGTEXwU9EWPTdaSq3Y3ap5o8+XqDajrZjIJiK8nABEYwLP5N5gx+oqtN22XT+vX8Z
/S4VYuW83TnXuXOIIicqgF5Djcng7FNBCeUd9i2h1FxrIm7QP1/qkYcKcxJTQ1I1iFiaCo44vD21
WXI/icISg71n+1sPkWMPbM9HpjBTLkVE3R3EgS4APgB5oWT52MXtRIlCdVEpxG+fSeoF4a28R4Xk
qE4F2JVHTkHw/Exqbqq/uzpwij4DVwDcw1JprxFuRsLmDeUXarT5EMSdbm6D3kG57gu1UMwzltA/
r1Au/USramRLyNDeeXm5tTtq1wezkXA0xamZQER12c9jGLLY5A+BchGN2/nGP7w3gpuOsxQ225Dp
TSmMVdmqNyQ9QgbvSh1NBaTNn6lC2nxLwfrHOL7bIJVeEfexYiUhRO/6bvz0vxnfpLwqllxd6fd+
X87t8PyXFOCKl1pswH/3KuUdXOH6A0vhcB6l1hDN8SzhZct0P569fmjle6BUPOKpMLmWpsgcGMUe
7bFVBXmLN+ZeXtYPZKbe725sziZwfC+ejgvuw8mqieobfkg1g2PfeSvJc6ERPN8WXPB4i79kBrDE
icPk9/TWsjwZzlpeDwCGvqq9rrV9Zikl/HmlhBCQIrc741s/VSmV2IAuq3sDulQmOXRs/mBDkutT
JtRHMr00w5o6mcDm8zb4wvfI+q76wDrHym7VVM8I+ytQNQ0qDuP52EoODZDbu8d/zHfBdpHfOiQN
yrYbwLRY7KsgG9svawUk4R5cb+c0QqPvbUtQvgW1vpI3Pm7emz1lGHJNC/V0YRe4WNMupDYIgiIF
Yw8hj7j9xrmIudNBVD5Kw+Bj8ZHQNcd06cFaeTFXRjvIY1jr5vdSvGw6ecrjfVdZADT5x0KkKDUK
5pvzvRSGWGhgnW/IrzdWlFL+hlBYzdEqb2K71CI0CPfnqH2dEiZ03cCSe1DCI2K6/bBgWgZUbqKd
fLmiVLw59HfvxPpivXDFnZjyB0Q4alKfYyiHtDU+Irf0xerAaa3O1JgWftaklMnBS1sq5St51l0z
Ml/b3s7Ip+8zQHPWO6W8W8Z93DQW02LlgiQCEN+TkgKj/JY0uKpZxQwoxZzK5myTy56RU4iN4a5A
m6FnRV5OtCE/N9AqObCtU+pgU5Ovg6hyy60A5JmNKJeWH5sTlIVqsNLj8gljXPNzEx1BPZJX41GH
AhkLcOYri7wHe4AMrnppX/aeZdc41jc3nJXI9kOoBTy8h+Ve5kiDZKYTRmjfml06pIwLqSiey64S
snrLrJ+qaTa21EYjOFzbSMLWV0n2v8yxk3wamIkHGlV520jsmc83XemTGYcS1fUTZbqurCj16TTv
9sl1V9EVGr0LVmueiFSefQQOR00HkM2XIxRDbab87MEeuFN+kTfV2HVr3PojDSNrhPcGrEtlcjnT
9X2fM8qakMsWUDo5fegRD2J/ORmccl3xJy76Nt7ovPp0keUIVXxeOLgpfCZuEkAvqKoTKU+V6fa4
MnBXU+oTezhvFUUgijke8x++YZLM+YY15C9wcs2dO7a5tmnsBR8ZHR8v27aLN6EatwFoBSgIqv1p
dIUbPQEt29Zi2l9q68NDzvBz3vs55B8ZNtkfPHIm5vHpzF8a4hW7t+z9l4YY8cFqy23I9xO+QtFv
Pz9SeJwNYRH8s/odyolTgknam0KKFCPHWwyKVBuxNTRJ1ae7m5V9RnqJ3pbVgB3EmskeyKZArDRL
swhhnGBKQa408HMQy8EEP2S0r8cC5dEWSQbvQnPxsYGeXtItn6D1a5fA1kxN0GxkQyrAnIi3S5hi
gTtVNkTxOGDTWamAFYN6K1C+9mLAC+KRVNtalzMdETN1r/2aVFgWgYflMQh21tHIKALSTi0NJSHr
M972O2MciOoxLAWYQS8S7AWcfG0C7pqUel3fPey4wuujLZTbowj8upy7sEfRtXoTtp54pBPH8jHw
Pt85zhjE38EN
`protect end_protected
