-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
gWhg+YIc9pWspFtw7ej4CPljpIe2/GjKOIeGbRXu69xX5AGMyJSRkHudIkb2DUMD
KXofWUvZ7ULyhh4kSfd1SfPmiakxWG9E77yrPrlDURAri8h1oN5JocQdsF7MvAhi
Kp4A9jWad+fnZIF0VF6ovVt7PhNsqI19jkjgME3Vtt0Pfui6RG5w3Q==
--pragma protect end_key_block
--pragma protect digest_block
lC3EpVIW3ae0mZPGE4ccfmWki+o=
--pragma protect end_digest_block
--pragma protect data_block
rP+A/tcvASZN/erYrj8EUxVZcKipBKRJIjJE8CezoBd6sV+HmhDdWEyMs+xWmWpP
8b6M21QftLV/ABs1oV99GBHhfcGx3bg80R1KN04veQo5zHYuesM2qQ12LgBNHyHI
X9zAg1wjFGM03pYaXZzUZo4vsvswUKapls2bWhUhO71ojPWSCDszuHkltSvyhfB3
himC4BzQ7XQu7y47qc83Qo/fsZdaGX4gqSjUZOjixqSk269qpx3gnldHVaxUnD2T
biIPT7AcQ0CAaeLT9SZnOjgtSDk8RixIYKTG9wuegT10OVGWF4MfgVqaCXF6bvVf
DUuG1bcQ1rt79swtIDxj+uEaR2pasWeE2+gIZzNTQBho/lipUuGgPkn8U0ux+9Wi
jQ5n8i2QNQbqLySkcQiC2g+0OsuS9fY5Sio5hMbVf8BNG5q8go2JifRp0tiiCOZj
8ItOQfpCdOEzl38IAPRuFfxS7spnoIbUnMEhfiJRI1OALKbAjEXoRt1HnnP45eJ5
DRCCdc16SBPWqVZnMB8XKBg6KRJzcg+As7N67qMPfPjBhBFT2hptHhU7UNy6Bp+b
OH0H/cUFfFT9t9ykhIIjP1kWmlNDvRyFv7sPeKQSPk3jrEWo6JUI9F083hVWXU64
RU7LrKR9KvrE38Z4zcBH8Bo8e5HS/hFTrpYwtrhu6yd8lzSFNbpOeeoY2wpfbq1O
MZSvAuFbeXBJibvigYWyOK2FtVPE/vaonTbKo+4I/ph9u3iKuPgeRiND0KlIlXle
6+MkQ0VVv+/v/IeYI7fqnL5eqE5pVOtYga7AlSWTkss0NOUYConSpmajp3sDVw2I
bBII6lPGhCqZfR6ck7PrSzB9gE/RR4uD0RbZs/2DrhbBz4WuoR3y8iLQ8Q/onTcv
XS5dRi5igvHMAPaaV60wLVzaTykaKB6BlIg9RiOfqtgYMDQuu/3798TtIijpHKVF
o6iCtkFYbLBWJowaSJ3z9aCZq36I2gRtvKbFk5v04F7U5d/bEkzVw78L95G3Nxn7
dU8n0Iq4VVjxU5z4G4Gjrrg3HSjkhMkhy97ugRoptxLlNdbqXi9tL6bt1AKzGUJg
GOg9nfnDIzNo1DHhcTid0/AZQjsTYCx/AUlJwd4ZnRK700yPXY7n3ptOwhwIdiB1
nZ53OCeI2EQ9BVKyAbVJFUcrLyVXFWq32X64QIkERNvIzKT2+sv3Ne1EcvBKsnFz
+WEoBbQkVouQlqbTdb53ybKa7ihHCehblKVED4MW+LdlXyAQyNOCjv0yLA8NyY9y
ps/5smhxm8Vo9Uq161ctU3BbXpMytQZzBKeJdvhN+dsiOm9oTebjlK1Ex8aRbMuQ
tykO6qC8E9SXL4dVwpMCZAWuuCUZ9LPyZHJXrdD2yPwfOj5aNJpZN4dG74Qsuage
QxqSGRg4n8ogZ590rKnPLpSmy4zsNjgFOlMVESTGW+F1YzK3a/xMG3URtpl0GDmW
mC3dPSRN8PZjfeHNh7SVWeCxVFNq5hJfVmXYqPszAKmeJBCl8uAlUsG5L3k5kR0t
Kx+ERFhYKmb4pV96pXBR/vAYcXo4/W0c/2mbTYbZsnigBft1DEu/cPwyzwQctb0L
I/x4AW3nEgz/wTmqRYkiFCN1C2gf7KssOrpEDRhnlnYgdhjsod8w/sDY9KZiIBrq
85tU5t0bDEU18d3+MGfY+dqucGxnPgcLgp4FpKKU72yFQnmBCx5vr08s3/wRwk6d
juYrHZtNkq1QIYA76ztpgKwsaaZIl/dgpsD3LA5yDyJ6atKApszY5/mQdewm6lSh
ImnxEfZUEplDEwb5g3+gdMnDi6Kt4bS/QNBIk4kUkJ22RxPsNW+rtC4/EqMmLXJF
N++sIkUX+/ivVIzIOUyc/ICulFgO5FBUIKDI5/EXY54399boQ6H7Cy+WkuQlGBQ5
HiuCqR2Xfpo9VXrhX7BgBOadDBRXY/iQgFCHiTR/EjfnPrcU0mYM7txmF+cYblwK
4RXJ5Fb/PImUbkOWPleY/13cOseKt5zhM+vwDEMvpeEXhg0JknEcjfIxzTo/rlF8
zr59N2r8iO21r9aLln1tG52cfdZAhBhVKP5a/yPgZQ3SNlwak2N3ZYkDgRf+CTsH
s2LMdvzIE6pOzMvu+1chEjOo31M67YkQNDuc9h2UNnjfDtNozVSmOrz22IPersl0
ns3G1CVbMhGeO8QQy2CRMozXwhoX9+97qHwi687qDlfDcwy9m9kmUpD5AWltOFHP
NjN7om7Byl0zHJq8NphqNnOW+9Jk2mJH0oGtX3G/NG6eByt/kIgSS36JRN2GJM5e
S3ZU4rn6r53Wmza/AHKPcVvwJ8tKoXXNCtsgF3+QUcowD4PXckG7rrKtefX12Prc
APVJLumifgHJYWePlswYfDI2FYMDpaj8MHAPzftr3ckbDgg9WrcnI2UZzJKHSZ6E
+fXf9WMHvaaI8OumZfcmWmYbEg1Uu76GNzQaXnP9M1BvGXjhWB8Nj/EJuckHdJl0
OhAAR/m6orq/9+pIYs4jAjSuX3ewmhIaOxf3PDFHqwLQnaJWhicoX8iNcd6LsLKO
lA97KKaSpSI/FtKGJFnWz4TGYwJJvuSOmf4ClTfD0utWVqPTSwyAvw6nFp6dHq23
JJXwk/NVv9SwKZ5Mmi1RzVAbhGLWRIMVDThvh7TNGtJFZkMPM6N3N0mfl7mFPl2v
ktA5DZY7faMOkn14LVqbc0gsNQNM3HsS+NxAfVzwIznpSuqczkqtMw3yEkg8Z1o6
EybE9nrLgoWNiYyzuFGPbEbQEPY0ogzwC3gvUZbSYkKyQIByR8oFkX1/tVdoz+8k
vUJed1iD9b3BEumAtzFR5XSgPo2BzoLst+NTFAxflncLuMEZNARmrksRdlDMtfen
bRc4D6wki6DPzxvorEdoHsazEM+gyU3MyrtSKowFlhQU13YoWeT6hl4eI8HoOihO
roSsnzWPh8gX2tMn0a925bGsw9WEiVo7E7+PxgeXLL7W41PWirx02cCbj9ZEQqET
hR0c66mi7DH3Wr+hWyxTI33X0OKIEG4UZTIwqVnTWTfWQie1XH0hvJiTgMz1vu18
QsDZ1txsOdlZr7RAO7eGBHGWXpsuhp2vLRK+WLP0IKtpObzw1Viv+RNUtfukw62K
Qx0jyYCihE8LjcunwDZTrqVibBQ7Fj8XrrhThFg16QodvuPkAPC2F86lP/TgmCls
IqxlaPu5JAep3yJbaQ+RyCD+sxRAtCoI8dB58MB+/OBmuJWgyDums0QvjU6yh6ev
1HilsjEPFQ59TvIjp4aojbg74IzbQdjQqpeuKf0+qzbqrq44F3aHhup+tnGNb37U
QAxdmF+fvHr69GFXk5Ny/3peYWcP3/Jfgdf1fBp2xKKu4d1U6KDS3mdKqg+AR32h
HfrBzs53x92O8fczFjdftiEh6powE2dyiifO9ShBKkFQiEYXamp9lihfqdpyrJaF
lltisfftadmX3VclDi8XHxxf9eMxf6ue3vQe1+EA9hDGCE6CXguhYDR6hI/tCnYH
7b7yMqlGhqSGQPMPn/WgWCz9azzNptEMAWwGEPX8lZhSJx+q9uEw2Mtk5JvLd4lJ
+Ht2YlbEJbNawk+6f10nGspxiQuOEvgPyhjK6ANLjUPYrNiYXhDXugk/bpf6LCbT
ke12hzw71P7I7d2H2KFIU20FzZ3qN8aQH51sXG21aLJ3a2JX9iYCdd+qb+5QL7CW
LgUPvz7zCstftKSgAKiQjL4A/99xcAtd9+dl/gWPNKHjl1weKuF1TQvW/gv57+XP
14rIYQV6odEHfdMCyIqse370+Bzcls7tAIiAaehyhyKpMGmhy+8UzCmCd//9oMm+
zRIl1OdWrKh39qQG+kmrZPJKJ5MQuiHoOsc52IS/8fk5N6OVlNdMyrIN4TsgghyC
i9xdihps+DyJ9TOhbv/f1Kz2msDoAT2axGGwoMKEYNuEcvtoyI1OpqEgegWT5bms
W1rpIK5/57HKRrU6OVM2IJF+386fItHa6Ay+9JdkBXYoVlKHfjW5gf9i17FjamEp
Of1InD+mE346QlP7RrNOTxY0oEQn1lItTIIntnO00M7WavhSq/tdB6laDeRE8l6D
B/U/cVgml9a+7o+J7B2toJq8UVirYP0sJT+CDUrGokJufTYTGpGfn8edwuCFthvZ
HzerTDyOyKZ9FZk4kv7ZNDAfYTKh6wjpyHMDdMzwnfhI7cQtVfZWumrxv6Zg8qLm
9BnAJ5a6x6yoK2YtDXZfHpQ4vP7e7FWOhKZJ49NRgbnM/Lo8JZBYL4lFlTgGYcQq
xnyF+YKb1UphTS0SxVbhKdBRdOGxZYoJzGAtAanGlPE4UYFyNfLBgQXlD4jZXgzm
0w4XYAMqZwSKeUJTWbhZNcuWUjzBfUj2pAJKSL0XxG39croSQqpg7l3jc4zQh0SF
pwpytr6bdcPzXw+eOseuLn+GSHaMtFiGT4fzBvDuZzyw6pf+XWAwgTmzOA2LxDeT
o7MdAelf5PI7jAoOknkIaM3dFwb3ZGKPtn/MyhSGxLk8xRwbt+EacpPuBnaJLSZ6
Eivp+x5C9T6L1cy9mF5Ccn2ZLgbH7MNhfdIRcrzy1LewOzgB4ljiIUYvT64fwJ9w
JCD4SirTFYUCiv9kx8wkAaInegjDQWjLjiPqforTOSeOt8pRj+r46Au5Q8STDQDM
CZ2S+TcC6M4ichsLMPRa4TuGLjtNl+5yZzuXlAI1CmQMO8zArhEWeH1mOUIfXlNH
NV6TfJ8Q4uW43zDrgqUd7zFsxFv+wXNVTuNJgRXk1od/KotQ1gg+s77RtzPiUyMR
CWHqYadKCd/ZJanVZbl3/RK5bv9YPL5W/sQsmWcE1RgsrVihvYFPl3d5zwZ51RmO
CvgfB5iQ9BwgKNyq0++0MwABbN+tD644N4lN/gaAOdfmW40se4jwcMeZDZ2gmXxp
EciDDOGCljqQ+sThmNqBNFXqighrK6J5jYYrAMyp9/FQPW6Y1xoZ4nHojDagb3G3
/YVUTVJXhN6jF5cWfDE6/qEPmWA+q7271hQLpbVrORX/c5SsEAyewKSnSjMI/10Q
IE9XudSBkYNeabZzr1xbe++FQhu33VBKD7jirjfPkUQ3dk6PShTVb/XdKBvnWsPt
fBk/4JjkWrytoIKVZxo/eFmpyiQcMekKrCO39KARK/43QISJ1w5QxSDumDUlPpcJ
rtMQ1nbkzHUB+LepfmPeSLiMvweX9V7fLqx9HeA3vU4htvyB6SP5Tbf0dGz1Zxkq
eLnMEyHw1+oB+KtQkul6hZuzfQKuMJsy3co+GsJHaif+ceqODERVHF/qt5Frpr0c
3AN/cuWOqPJHYEprpNP1N2DxMRJI2W4HQBO/NboGFwU5S0szFwHd2QTvH8GNrFv+
4xjtlyLhxqvkYdQ57AG1aQxAL1kkgzdgniY9cL6Pyzxhun31U7tbOtx8JThw47GU
LX2kMLSHUsX2QeFOR4TM6BgI7I8YVrX+2Z073gNtxJoWUBC8MJ9iHvUP0E898RTL
RpVZMM7YWsw7jd59FcOu8RluMYNKr1qvsPkjNNvz/Ucgc9a+h8JImYzMeb/OWpao
3zBhr9DV/4fdaCxPE/bt32bpBWziw1OW3N6QeOl5bhuNXVzIynA+ab1o2IMEOgER
VJpd70CO8MQvYXTeA51RUdj6nsSDKXF4iTfdj0Axs76tD/cSfmpEfc6ul3BwT/5W
vIjL1dsFrMqxrdIwGfEhADQIF/PCZMRoM7Wr3e+mKtwWn0WuAzDNxg51qy9KFsVN
5RAp+GCLuPtyJ54K85ZWebUVe4EBZFjiVxNyIjyT/hBV3kqSXhxLQg33ddSeGpG+
zkwpXV8rp9mgRKS044+gdXB9PBuXnTvvk9C44/14OYy9qZ4LHPWOv2KDOvjKoauF
N94GJEpNHpSImlJcZtBGmaLnexp3mNN7ZYkekwK5lY8Fx5ui5rRSIocbAHXg70Yk
p5lXYqsRMIHW/kkNh6sRHGmBZHfYfEDijJmQTutJex7HGec16m5Z3lZSATRczgpg
eigIyZMPms4VMhKYDAfsOz9ZVQBSmdNAieu5tFBQFtwQABQqq7DSATUuNMlQF95v
DZh0NgY0Ry3P2oV4akPhhYLlDhuQEA1BKJmBznmF2PngCZwC4yXCVAbBQvKTbTCE
n6Ix2lXSGfmjEETxTs2b+WyFt7ObVN3WiPplWXVwb5+P42cfjHrHSPgg4pcqF1MD
7ZO5aoCBV4vYx8lFz4Rkne4u30httEoljQSgImtUbKJdN1nqvyaLN29VhlakREYR
GmdkFMpVzCU562qBCT7TCkDj5i5v2LRCyEZ3BG9uizgFf2IPZbznjw6Wj2+6IXMw
YPKQtNMQJTyawgpQEVTZsboqMsvABa23FNFBt4A8oAXE7AxMRwdLQ/NQLXnJ2QAT
a0pVR7WTLVrlNuiOI6S/YLlzyTBTM7WuXqgZRoZ/0IwOQmwX13LqxcqbxlMjVzri
W2KbX6U9sf+UEQDOGvghxl15iaifaXngCkjiugQbdIiodyGJhkoKO2/oL+NcfrcT
XOH/99FcXOCi++EHN7YmutO3Kwpr7Z2FW9GBcbIZTWxVDPjHNZWCCoUwEsErLoPQ
j79JCTReC4O0qEwnKNjLUN5VFHz1+CUcDXGxtwkRRuZpJMu82Yt4SPLGYUgZIz41
JkvI8SPwStOBLGfEjNvUJ54aSOBv1jCeZTVtiDs/8I6A9HjSQ/xPlkbZgHwjXl9n
tWLp99pd5q4oE67fp0kxC+fK8jkenxu0eVygY8HFM5NDY5wEl/r16wbcK/QfRRK1
Ta0rOl6o0QhfKSu/upPoD7eEKHL8053ks298Oy1vzms0WHKcoW3W3xsfuHOSPG6F
ujvgfMxMSyvnped9E3+pEzpQW53TTfq5s9Ah1337smsMkFZcynH0f8WV1f3ZUYS0
JyyLYl7TAsMN1N+eJ9uJ4l8WTKrdBMwphTzWOencgrlLjBYaygiT6ssZE0l9+HLo
do5Dv4JPjQ2yCzEg6jlwhW3z9giVBl/O8BK4FFvIN4GXRP0MiEf0/WUOgPscN6Be
k+OWWWeSbJoCmT3ETfo2EkrAD2o7kXPEweXXsOqlNg3+NAE7b8dNiRvWnU4PGO14

--pragma protect end_data_block
--pragma protect digest_block
H744mxdCrl3HfsIoSoRLIpb4cbw=
--pragma protect end_digest_block
--pragma protect end_protected
