-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
FsOYWurIbeVbr3ezmJDTIL6+XpcQMAh+apqPBD0teuZTm/Ds8mY5xgw56HtvNrQr
vLiXYP3I9acG6hy/SV4lQFlEoxYIeHy999MxlRhe/q6HmTNR6ylJ56APJ/wtTzrR
0w1IVqCkE8uECuPFOx2UmfWuaQ/6uc4BZSGQvjXFEewCqSwPiSS0cA==
--pragma protect end_key_block
--pragma protect digest_block
AeleejO6+3DniS+9YUx+gjYrne8=
--pragma protect end_digest_block
--pragma protect data_block
vhNyBRWkFUdh/zwFJez6uRo6zZxM5UHS7vXhiwCZPzpi94h8CYwnFS1yjW+fOdJ7
AziAHernZwUTU519n3nuIPClFN/jx80OzliJonD1vv7PC10Bn5HVr0QbQ8x72bFd
kDV2nNbZdlTp2RL64f2hpGVqDurDU8bNabucV9OWECu0JBfVEng46ja39091a5y0
cUMdVHoDPAWERxRuMEWxhP45K+6Bb/xPltJQDqZTEnxlu+XV3P99fLVWL4GyJpc+
UDgOh3OVFpkZpgl896UowZybQhDPluhITLb6i/7tCXaAtQKv+PhF5VscF904zsEW
vZGO5FAYvVAiKl5A/pttPtbGpP4ZJlhsxsvF92/XySjPX7irbsuguOg2YmQYgJle
cu/KOZwXFCri+xtYrQBgMj3gx9DXd5DWlC37Ufe9zCD8A3K6Wj1VjofDAVYxkOUD
So3xXE628mqvib8YlHEuQ3e8y87AUIONA2SDnxQ82wPZR1V1ye669EIwtO0BX4EN
4yoRt+iv7/lCpbDOn6wbyWW8/x1ANzzR2i/XmwY1BAwo+wMIWycSPahazL00S2hE
lKw+kNQT8zoo7DsiG4S1KauA7wcNYmFGAzTTyqqCAjQMd1Jx0h24f1Bj13DaKAX1
5YqrIiuwWQn5K329LvO+QmmhXrmTfFkL4JOv2oLKBKQvlMNbljz7jm2cgN2xhaPi
IvoxSyRqgoNkREg7DEqaZvcjC/7RU1agOIQqYGLwXIDiXjiLsXTfbS2486G27wxO
Ums2GYElQawk6MaVF0kBCEcssLQP/TuBjzuM2B7BbtnDbPPUurLAVI8GAluYsbXa
z7BXpYOIx+mt5Btw+KPmvzS7y0LX3w01MJYOX4BQvystcLPEBoiv7PgboBN62g0+
wvyom++7WqsOGQ5Gz1hupScqp8wZKqRRAW7FiZqRVbVskle6MKka6crEC0SWKy/e
5mjzGphjyRNaUdIeqD6VIJ9eFo4ETtdnvx1scLdtzQG488+4N6UP00gSKgLSGLJ9
fqOSuoYah4bLBq4tGb+P/vCd3jYNS6pXFfG+In2KcdBEprJAUW7ELx+V25DP8loK
8j/2mpdOO1MXfbvLIL/tvI0nYnU1NlCVfqF+j669lnV0N3FbcbfsB5/SBtrbvJSz
Gti9m3mQFyt5EV6JPfWnP57+WQBPixMsgt/AX5wLHbxEdYm2PaZQlS5K0bGZ+rLN
MwmjbjFfKseJHrT5ZTJIifWtlXQzlJymU9OM6dKOxES+7fZGx13VcFlwwy4VNTUo
vvKOCfvAzYb4G1MN7Kq13B8VwfJwUgspi+n0F2ilugob8Fn4i0jY66j/se7+t/fW
wziKiqK8RPzbCePcc/UxQHSQPmbWrwxj6+xEcOdhqdP80PcAt9R0xX2gQ9xs6BGP
tkrpLGkz+/18BGEMrOM7hGh7X0boacatbAMNaKbZmjMfEl5awM3OyZ9PfJGbMg3G
7vH78AStsqnJRwvqHsnH3BgLZu6AnVu+BJeWc/I7atSUCNPbIsDBUXM6ht3pGQsr
tEtVIoH7w9dvKGuNha0eReUycaSU9R7+oU+nlPgQnree+vxxCaFkX3SiZpRCeweD
DH/KtvR2d3bt4O8Rh3/u7+6durxM2JeqcALidZJ8hXa/oZwv+jHnF5+0cHp6v7cW
ZPqUrim1GPC/K5qRTLRhjPbDthdxwryXYtU26vf5BAbZTEM2R9VQTLQK/gyxt3gy
l7JK1tTjLmKaaU0p2ZWajoRSt6J97/mLYHKsADU9HopchI6sZzh7WMbYEdjgbsZC
2r4QLNQ1Hde8EsCJb/FqfFyob3A3LW8AvJvihLYpQWEZq844iifAhx9k+9hSI0GF
SxLGzkKYLv4GuETxmf7F5+FPj/MOPFoS6lEs5xFMn1hOI6Ir5X33fVILOJ+8CFbZ
537izYymF0BH0V/dzNB1eXY0+jN/AybgKA4abW9Xf9EWeKiHPzjVy2niu39Nf0US
RW4skFGLab8YTISB7OywzD23Q6FyYrQMDHNGTmUsYbKwYLroOWACXyylUUhYqNGf
/gQfEUuIEgRrFM+bgzka/VcB9gw5t4WFBjt6rQhNmiAoj2Uo5lMXZ6c/Hopf+hok
WsgqDsG8HiXK3OLncMcr323+yyVXcy9Fkea2b+jagIu8nfIIxeuulHYBEEfRee8T
+Fg595smjA67oOCQeWx+GC9sn750wvAgeNOCmUXgvFcdbpHycQ+rj1JlirzxgQlw
GO+MHxiyIVOvqOnwNx0Hoojc9RZ8Fy+wm7NDSU7psNHxRoPh1bp5ny7xHZRnn3iE
2VQWWpx4CE2pyELG98A6q2+D2bTugU16Y8sK308XVWN83qrFkEWJRvU1yVpL+3Ab
lgh9TUGpSFCOGoSpVMFORuGDeBhJYc98JI5thFNI4tQruCZrx5F7RV0cx2mnGXFH
DnL/hSY2l7qlATj3Mse1VCe7z8gVShfIWcO7uRQzAIgUIk3h4glBdXRlqY3RDsCe
4FzBYC491CcJBKhXuuM/5/ccOKBbG0tVmpZL9Bxn4y+YUfOMKNr6ENILcxylrEVR
uZr1slp2iyVooCHWAPFA0gyljaLOEiz69yAoqFF/OFOVOrZu7J6jPVGAr5iqyQPR
4n/OAJyhAvrk97qHgSnHdCtZ870yJp0GNzqhbFjQs0DyQk6cxufjuJLl/JJYNgeO
WMpHeAQLCttZ5MUkuuQDeWVv6d5LLQ02PvfysHWWcv9aVO9YjaSeNfXWQ0B8Z/Ls
rrZXL8eSlo3LBEgW1QdDamosZK++7EEWkQXwgGXnHWWPBsVjtzhGMmczy4+8SKdA
MRlDhTm97oi/0muMhquDiB9BfXVJo9o9hCKq1BOcvszr7uckmUSIPmKZEyqQJhel
eBA7apH9e6T03m1PMTEhRLBtc2wVA/OkLCyxrdwAeZWXlJTBaSu4Nb+nIsupJ6vf
xex5U7jxjaJ067Y864lS8KSpHWzqhsrAHZCeEnooS8pJ1Jqg0qupU5c0whho+kln
oUIzk1sOlBNHaqfbm+FWcbwhO3e5cMUhCLu6nxyJb06FgHcgHHYtgse8LdTXLvq9
xS62La8q3gH/pUPV3Z8x6dVnfB2FWNL99ng8VX1ZeCZLAgaxTMcc78CdYeRJhf6J
bL+77Ry2FmzqIBn5EZj+zm5QfiWqyOp52ifxKi2IMy8VRMDlf5JntNrMB2TPzkPu
i+EpeCsbEAutQKcPBk8Ze9/WmRf7VIkg5H3i/EPF9ovQhgfkdTnjFoTZp4vLzfr0
I8WX7C1K6DZEkml/zvr9bShQ+/ZsMJUOPvwWgV0miLaywIufYBjVP9flVFzWL2IV
xLpAH9KqZpfzIVwdotNIoDVQsA8/wv6n9MsO21btmLK25qVDzyc+XiLEw4QxhJSv
8XlR4sOpODT4FDS4/2eHmXnDidwZgXggDjtHOfWrc9fiMFoI5wJCUOocMwZ6RewL
Jpoyvyn9dg9nrYu5IcddaoVjHB79xE+AzAAH642wY8Y1EjQ5mTvOANJ8wWAeJtYu
2B51s4vIo9YpOc1kL1NWgF8us57jKTTEs1neWh5ypt9HUBML60BcymqnZ/iQ+HWq
I7wqTxZyvn4R2dUyEOCkNeipZIoKlsD/9czHrT0PyT/7SbY9UBVWqSh+R7xFAhRv
rd0fAhy/pE3Xf6pb9AtsRheAQXzO73r8eGw90J6Iyrqs0FfOqRCPzBfxkqTXyiS8
wQqlEFaMKYPAObnH10gXKRSQCiHiXYn+FGc7o/6dniRm5WGA1j7WjYWuJgZbt2Uw
TgwSud8HxRP0xgx4PS4ty61PJRBOxgy2WCPxkAGKGFsh0oi+1TRbjPKhIIRZUkSH
Lw7dzC6zIdv9TUkmTHvbbeFh+7HSrPGhWlbeO2yrJ3rOhBMRakTQTpflwC2HjSFZ
Upvcxc08z4+AVOTemO9iw8cgct4U3sgb6DJ4xLRn1G4IF98EqqnO1n2+4ZvawoDO
VSX3pAyBZHxgeI22QHSTs3ye6RaFdII1D1Hmmdk3imTAE/7Bb9VuR6OShKLPQa+g
43Wm9asL2HWqCPV0eokZfUg6GiTywiV+Ij4pAegnUs+iXVOP5sTOgBBlXEYr7y+k
8/qRkokalPWFBCZ7ucmTBrwf4zYsqf03sHtJh8oOpHpvDgxTp1V/nqWHiDQyjcHN
xzxH3JxleyrowUu/CW7gKpyeVYhk0cYOJAbdE0iGicywtoFkE+1n97v85rhvUAKO
WWaVLhfH2Jk4ri7CcNxrikjhOF7MGse/59z8fmoqPX08pG/MEeCWJmsqsmUng5+I
jBb6KwlUMDY/igonYW9Hsot/P2uQUbauYS5X6k6gfh9a+M/G+ZNQqKx+wlH6Vvs3
tDhiTG9n44LSawu/90HVNEAGUXcS7PncJ5sMlTKDsHqPPvDcX+woT6DfouWMX5y1
Rgafk/wGzlzsUeYQuqhBMIw56o/yAmAuzPdgo8yJwIPzw3WxmBZO3rqkQh4nfYMQ
dVG2kZGHSdpyURdKrLq8Bb/GriTZiI1/PGQmfbuucTji3Wo8hDMxrZvNqKIKPo1u
q9otsARcxZSNyxuupfrsQGCQcIwjCmSN4UMIhRmIPAEBZHiDYamvBP/inu/oeUd7
kx0IfrEHXl5ak40vGOcOJROBb7I72TydTtjcQ/ArgkeJsV/YjCDigERQwvA9qJoI
9eq/k1QWnTmxF+V9cy+WglxPkq2rMK+g0ZzbcbSPFmyrtjdMl9kAxl/UyWKo3ZlA
l8xI+ZzEZ6YLpQjW02JxugrVtPbhJ1KonROLOgdXbNjaSYJ2eBKAaP1VP42dcj5B
+TXYV5zEdmUSpSsKM/H+62J9HOqCk0+k6XQWO3j7SLiBsMOtbNUNKO0kuLRfgTKU
nDXala6idDTAWW6fVB1KEku+rnYAJlv8J0W+3nF4GOeet4Wb90ZokgmYE261fJcI
nrajf8hPlc6Evk/S7LotqJPnJyq2GEmcVM43x0InS+DN53qxk/2AUIIXhVasVHPq
/+bA/QXN+E6U/dbnZ93307UCVBmMz8vMHKkFmT1JLX7z9z0RZ04ePcASjMsIakjX
Gtm3EKXp4aMKJaUq0YLUwVhy52/qpLxGbdaFkXAASlpXuhGCUS9biBuCZk4BZDUB
qyVTFcTEVqlXO9/7YQkZCrjkcaSgDXGSyhL6bmaiLbeW+2Nzzoan6b54XPpX7HgZ
RUQDiUFwFmeChZLOYRTzKtRzjWpAVUqud0hcW7v50Gki2OrS8m64N2J4wXfMk6y9
1WNI90pjHJNoc+UN0XO3dIUnNdGq2pUaFKM8iDQkJs98TYfbpuHgcGgjp0iuzy1U
+jfWHKZ+WlFJQmdQmaAIxml5Clw2aypfLbi7qLOzWCNxAFrCODS2ugkwl2Wzb2Vg
oD3J9Y3tX6TWpqJHp+7zU/TfwYcur4CxAQMcbQ+W4YRlbM88MGnFt+uB7CeA8l9o
HHohVzpCQp1Gb2mKfASK9TLFWUhpN22IzS7PaAkdLGRVyHnTK5FcRrhAqOFASgUM
9S/cmsa+dh09rIE9YU4VxUp9AipUtn3daA9UINE39gN2qxhfsHup0Hu/nS3D1uqf
WLXA9DnxuC6WUTfnOq0niVg/7tnz0FNFVXKHl5Eqa5vbqwaoTKa2fglT96Os5drr
GtSn5tqHxsuhYXqvF3Fu3GjDlB6fSGCLxXyvtv/eEatNbogJq5I1EDJscqeCkJX3
cExnQLK12XYbxt3MCDYe6Km0b3cr1QVeQB1tBUx7Po8T8JWLR/Itcs4fomM+uWB5
cAXWzQUwGTXtfIcuB9rT2qcxfIvUMrZ12dt9NK0by+b6PR/aI3bx46CVqK9t3jmp
eu/s0g/cFSC2VeQkva/6cg2DMVOs/Afi0kYB0oy850x8O/ZBC6WkxTVE+AJpW4rG
w5x19+lDDrfZGio1Vb0c+/QjQwe70WyagqswvL4Hpw8VXR0Tc7ilStYT4dv2juuY
eZklIQ75/lFdmb1rZJk4jj0PE13/fNBEI39oTFrYX6kBWG+iBAiAC388FDA2YGAS
dlBt6dnwUXiy63Z8zb/KFnE7S/xf45BKilWyLGgohYvJM7V4WZeKfZfBf+ifmq0z
oOfRvUFTlRWnma9Uq6l9+epWx6clfwXYWjyuMD4xLsbw1C+GT8ZFjnbt9vl4e2kD
6wdYakjevZIcn+aTx0/hv7zMoZl07/E6Rd4tmZY4AeVsOsJo9GDXUhvc+ef/WGyI
OTp4SFVznTL4OcmxDL9zDE7BkseCtB03kYhtjahliRV53bU2Kod5InQotCWE6SYj
w6qOkgQ+8rUD9/UA2puWMtmAJPbwoDi9Kzen78bj4vwo4pVw1oiAcJuCpb/JOS2K
/D56xTlS1FNkOMD/mSAJ05K3TzgmRYeIkgC74gV4FQEatc+CgdZoiGuz5cyLGsS7
Adko6Sb/kdicnCe3ppWiNHXELMhfDUqv2NiwpHo3lLMzVr8ZUyOP/ntsNVjI4x5V
5VBz2GzYhWC/mbK4xFcAxlL0YU/2X+sN/wHkLlWk5xT3vK/HV2KHeDBzZenY+JRy
LL42bs+o6RtyjISQAoTkx0hRmJ2+4RvZE3ZoHKRwUfTsxYi8e99ozmBfmiL8EYR1
OaWWE/yqRvHwa4hwwsq7SiAb5tlaYBxg42vKty6xf8wwRr5WWG14Ry0gVeEFRkBW
j7b3D+KgqQaPsd06jiRTVw4usJb8coxk5PMG30bIIyHGPt54zzMm2rkiNHzxIUto
xoQXBE/IvOewxsSDpWO50zuza8+A4TD2wUtbBpaOSxbLBFVQO9bu0fOyVElFZmXq
j5o4CIiWkpdgTYYRD0qJKah7fy0M/sswRZKhRSn0tFjxY5hxaWJ/MXRCOMISUCEe
TwobSxjhvUX10O22ZE4R87oOuHvFTnFJQIl7NMGd0PPx46pRtXRQLJlcfBiwdDrv
peSYAhJMvd+Xt0E+YcZ/z/k6LCnAO4ootrVvmqzxJQjS51GP/2y7f2cU2fRwvJEi
1xf8IbKpjmqPwucxmfA+FZySySTS6l97CmRHRUCfmfkrPiSlN5sSgvYDxSHZljWj
A3SzEeSnusHHc6yeTa15KDnPeawiWDLjbhub4mhbyF4EEGtqjtN80QaFwamPxyhk
MckWT7u0TXpWBH+fM0m9YCtNuWYv9VmaZu5/8lv65YuUUvSPWTgWbLwZu1p4D6lr
RdlrAD1PzE0J0XiXvIkdvG+ohmxX17YQepYVD+zpxZjWOMqucIUBw6cAG2XHFPHJ
+3/Wtufi68Powan+TFt0psMDz5btBDrvdd8bjxC6g/KEFdZ+S3QZIJ3INPp9dpta
cTpcUPF/oOhgio9Po3ffeBspf9TLy/DpL/NmQL8paJoBiS1cCOYENFrDzfNFfYvL
69H+2GUinUhTEfb215T1PxTIUgFMT+SFYemm+0Cc4tCFKgkPLGDfZ6S4WyE13v3J
QerUsrs2qvmZqIG4FbGJDGaeAs4/Wz+vzUgOSNplOr5ps+IkwqxZPGxlv5fIyJHz
77GGoETX26hAZgJp8Nkvj1RA7kyDcFwU9R2Kd7RCE02o7yvfCoLgkCHyouushBER
jg/7PUWrJnlZB308gqY4iaB6kCPndsYpDZTpyv8XcChSPQbZYWcZvkDVEY9n01Ei
RTYa6UnTSc6oQCP4FofiQvyVr9hkmzTig2a4nxtVJINSrK4fyh8lZK1npyHigpH+
7RrPBysbPV3DsQC5aqoFQQZmy6lCynoNOXATxML+6kgI1Al3ZgQG45QIjO7hI6xt
GWuYC4Vdpa2YX8ixkRSEQh4q6E85e0t/vg2JCrw/Px0r6tVzG5B0B4DgFe3uI2tT
kYfLFzsgn4nJC+cSec7+387DCL/S2FPuc94TLynjQ+fKTsY0t/dq99p9SpVafyc2
JZZklzY+lj2fkJL4/8+P33T6PEF8+3mNp5N1+KPFwSEeYHl2cXIG2otCJk3fzfb7
dB6WR2kkzi5HTNLDphWojIvkpoUI1Ox4yE80rscDPU/NxB+RbpYd7mRuXCQDssZ/
pxSAr6aj+T2onsNUGainMRBByeze5rGrLU4JETl3WOVPleh9TprQ9YXbZlxhrdLG
2KV9di3secdr0uWj/CHKsb05S6JrxFM3kuiXEt75oNRswYJ3A4ox/o/sdY0NFKY7
IG7KvCrNy+NaT1bt7mMGpUYuskLh0Fd3n8l1OhrNUeTbhHnBMg0fMrqJgxxOPLwP
AhkRcxh3FjFi5Jz1NvKInMVEqk5HMAmpQKSMMPWLedZ7jw51JB4WkTpptvHT6yOp
AjuSk+tlNcydIlh/G+JdzaEw+HIxMYQsZGRxi1MPcA7VbqycYq2YpvGQly5afpqj
WEzRJRoxoMCgZfWeDtZQ6rrox9StLD9VucL5VeahNu3XXUAaucdoqmdByLNB9n1c
5/WFGG3TZdWClW7s5pQ8Z6a8blVjfNFQ15Mienk06GWV+XGKyeA9dviIHnJbMxDR
jRtMpOSQ02Jzu2FHfPaYgaJm31xUHJarZvbFRiPJT/7TrP0SnCoCWZzB2EDq4/uJ
cO/OtfSKju3HceQ6b9Co9Cp8SBG+7z4OukM98qqSi3a0Hd+9RKf7ozFfz5W1A/mK
va9FYNwlR+VwkGox8VjHtoPpuEe8QGw/CSuZDfbpfvstBzqt7O3MsTeMHOVA8+1V
5bfl1HgYbP/q6Z3zhtdpsG7HQHaHKNY7jgc/PsKkeFq6H3QdB/pIY/1FCg0o9KlJ
C1wG+FYcWHyCKbmHC8x10B/xbBYiRdR/PD74ZCpTQI26Drs1acI7jkLHUStz3+UU
z/eZySifHrDUTD9KOaLaYyz/WmeVl77STtOXkhB3BmvlFEMruynTN7Ze/gYvVA1X
Ml3KZidK4lFq2lFkpV2Sa8fi7updvTv4klR3fofl3dVtyCQcU5a6+dvoh9aaLyC3
JUNCSyigIDFqou2rpY5fbXkU3VYFNb9TIY2t4fZ1Yx4Pr4/h8SM49v+wbwExn67T
fLIdEsTGhwnNEjjyl79txj42DETWAngbs3UMAvXKAjfbwPd30mMupdf/LBREGUO9
ZqtG30RPFhwhApq1qjruJEoUY/QQtaMmI4NVKRXHTmkZk6qh6r2DapCt5mqo1guB
6ackX1abG7i/ZBYXpysa5mj5GmCMnkpXEUOcw+fB5vAB/BltFpWLSSOmqCd+L2id
9XJhObRCwQHh+T/GZgJGgJkiJDsn/RUPj61jO44hfi6kea3R3VKHMi9CcG7AwDm2
0I4s5XkoiY/nsMtiqcxupOoER4hlZxVZPxu0lfbgw0opJmb0xS3MBSjSk608Zk9Z
w43ekQoi2BUX77kOUJ4B/dO+0yQtdxzOELcIE7Kj4qv1m63v9s6v4P7riDxeDnl/
89RkEfD3oUhjda12tWD3VVaJrcoqXbe90CU/MstD5VkyRFhM2Jhr6KlT6BPw2v9G
s/gzNw1Z122QMbO8zlFOAPowtP0U9Pfm3gPYZAN4D5MmnafKT3oUYCykbIP5TVXq
53QaSD6joOAzDIMPLgJGZ0XQrK1rFNjtjSt1n5XsSNgiFGQrNx553nf1FbFY94Dz
Dw7Z++DFC6h0lHsGtxIC0X1d2fyDeUF5P/F+vmmYwHkX+lo2wdqODVHqzy1sqZVZ
6LWxaKS57zDxSeGAos/HXaBRUKl39YcfSNL/zFDH+sw6Q9twHhsrPTzsZ8Xuf+1B
Gyk/c8O6rjbXLxMTrD/I/BIFX/GKca6zx78xHFmcgoieBbM+XNUDduHxNkWpFY2x
0S8d8Yp9kMd+zt9ehGwlOGETGaSaIi4i+iFpxYeTDFpBMg6d7922kSWa6ZhJFm5l
CC2OPWtaAgdCujTPEV6oBtXOtLb+BIwZlIPJjoIwqFgxdf9Q3Qg4WU4dmI7vBOHa
niaNIwRvB9JXVVXho4g/UZLgpcaOL7HL5IM4taSrpHCrVSd27tM/zKrey+Zm9OZS
jlS+/adYnfHAIn3gzZ8RI4lba1ZKMetcaAy/oU1ZYeHQ3v0d6PA1uvqvgrNvfYo5
hMe/Rm/eluoDuvTuoz4M1mrXIyGWqQ5yXGt1eVM0Bt4WpoQe+qUBuT37J4vR2cdI
zZQyqILiMyD7SCwpP+MutDHaRJuY0ld40PFpNwP7J3Uhz9M8HrJJIz2ip31jwOiI
MANJ0eNSvoTFeAXrOJXV58/mmn7oIQjLuQfPgrnXcw72oTFAMMn5fSxVODs+sqim
C7IGlHD8Us55MuYU+5NKRcE4uGc46HrxcKhNHPuWSnGWHVTDIREy46Q96wOJx5/T
ZBbChNsJbNQtezR78mKzPl4SfazTCgrpYHShOnjqbA1Rch0B6xQ/VjefD+P3qzFX
9cFbgRcfebDkJPJ18x+tsWktZ6UGzz/sRdnfOE/+/tqbd6GtXxTiqGW/FMnlJuRr
S6dFwgnXmHvPgGgBpb1EnScLadp1bb632ADNbQPWtFuLbMdsojHd8nO4bBJ8kk2a
WM5pKQQDRr/g9vd4MtWTF3UZJCTar6fshbzw36XTuTZTVDrZx7BBpngYxYLpKfgx
dMs4LRTiVKqWSBcS5nH1L251U1B3MLGSfrOSw5dARz3dRLW07sBSvcS8gHP/pffR
Rcr0ksQoj4JUxyjcTdKzxZjJkCnfWdFdFoLogXrXw5GKNr9pc/kUiJchvhTcFX2n
Av4PXRxeGdXfIZtGdxJ/jYmPGYv7NrBxFVvZga0NjgJvDWuLSGw57Xb7xxo/ecss
SG//RH2ZlV8BTXAcEAdrwptlaoYLxxX/7uBzT+rTtoDdZ7j9k+sdU6Zy1AYaueUm
v3q3BZ6RyUYxzy0rpl15kBGZ+I3/N/VazbS1pyi3K9JWjDR6chT8KXLv2zzAcAO7
a8vQRUb9Ta2EqIqWKPgnGN6KavzOX8uOhv+AhWVC6AfHk7HDVIikiLBiK2bw0VGT
DieZj+bhPd1I+anowltNkSqqxiPJSjXmGo/gyPKr5siNHpYuqPbKO1jFPjAk0MhR
cPZw1gmNaHaAupj2ZLMQ7dcVb90a0lkBZlT/keAJk4kyTx8WxOiIjjMJXWSYepoZ
88NlVjiBO37c8QvBXQgxTeNyF+p7a4scYonHZS2Jmy/ugM/3GGYIFTkp1prZa7X8
tzetnTxwVHU7vMsGfK1fjK2RrfdTf/M2yKPvqLlM8s/stHbPA2iuukpH5R8gmNBb
/l5MKUizqQFzBTZ7W4xWkvqJrsU0XDebc86Xhmf3VrRTvVOmSM/DwUyPYHLHzbx0
/oyuU8tDcEpKAa0XG4Q97BApEKoFib5x3lcgYfs1dhua09C7Wxc+lz0lZi8H8SCa
8RGgw/q8iirbDlIrgB9VWBtQj1efryReY5mqrNsEh3R2PoZoHLvjF8Jr7gpA+jPe
gEJKaxfMcpkYyQ85bCjja/g4ui8OTDgcxWNu6hzh/b5Gul4SA/Kd3TBYOrDrqIO0
5kW5B5L9fRaO+gwioVAjKx9acxPa+/l0OIaZJKF5J/Q8g2sdQ5ZrwajBOpGT/imW
3Mj6gGrpS1213vMiYAV8+D7Yeh9ju17Q4mDdL74iX+O34fqu5H+GMdFUe1rnRgJF
wD6HVObt8Ir78tRSU78aurLLLWZyK0lyeqI7axc23lRGwzVIHYIaIxQKDHpXhNsw
RYmj688zt4f/95BpgfRKOurx6d2FK201+d54jd5WZRop2MUMu8x9DfiG76o5K28t
9dSef+YzO++95LgqxAV1yBhPuGHB9er4tIbwogItXg2prAcmP4NoyJBu96GiZgiV
YFZc2YLMmWcLljtQc4LcI7YaO0ekr2sYIZwNsWaTHOoOFM6EDvAPXJA7Z8RwxkZp
EnqzEGpcu3qltdTEJFoON2mEQTaa6be9KqzuqmIgyP1ToYxmrtXeR5QW/2yMEsW1
NavFG4rv3US1Wptg3YNeUenArrS6Bs6etLV7qS7sup6v/uUvW3KS0bfDoJwm21/y
sDGctz0x7Wwm3E2dhmQ8u0EZpJbwiHJfNgj4FE9MI5y70kPSwDRV2wpXcdpUwBZk
uTEZPzDGLOrMneGcFjwrWAD2tsxLzUiiPcLftgHPxIA5xFGEToY/MtZZCKUqEMmW
YW079TztwDK7mSihUuYIPy450HIWiGgHg9yeFKK7NOpykHq0z/gxpXALiD8Bh+7E
9D/b0L6lgRrd7N4C4Liq6sLZIxm4ORzUTmunXgH8himrk0gsITrwOFzle2TrZ+CE
WqAcc0Dwo6ZfO1maJhnoxLCR1lMreo3p5eVNJDo0doThVimPrfi2utwIGUaprXPh
RNmq1WKAulU5WjBb2aTp2HUU6/0bwyXrAPnWLUHk3TbjNjEOwvVEzIRgEwkZl4xL
0eLHqRVMOyS8wrSj8gKqH34+AsII4y6ftD2//9cRmwynHBY9wVK3u88FpzsoC2Ct
kkddwwiIaQWEm3275BFvE7kQjanq7ckJT2KgdG6jKeXklo+MWtZtYPNxVyV+Pn63
THJiXIhFuDfRZvMlfL9BO8nOCkvPEaJuDnQTQFOO2+e7ZVPhv50Df1OuMy25lc0x
bdLLHImefSS+p44i/orQqjk03PHDnabOt/U3U2OK92njAOSEXvE8VbkskvuQzqHg
bdAMN1g+wEMmS3fwtsw3q1KW793a1jxlPztkCEPoAbXte9votreBtMBwqGeM4WdS
E8u8inMc3qbnpPRZt5dg6CAyVQEFYCcEe9NHmEJKzhKhGv1s0cAdO88zu8aRM9eL
n3wak26sOJCoxeAdDeuc21BPa2kckdWZ8PHT039KTBIZTtzoYm+dgLmapW27Gfyj
AxX2WdSxGOIkBwlMb7PkuX7ChV+C0DzK5fr8xNbQr6U2yJJnqafjAO/DYfM17swA
Ul4pr1ML1JIFlKUqMlgChw7fml9GqHWA1QyMt3x79sr7jOHEHGCMx1ZjxEV1KdzU
f0AFFLk6QU1yvf0SToFuVTQVSaBJS8ruLH0ZapfNjI3trk3I9hRY1UNDhF/4D5oM
JrbWiDuV6AmkStd6g7sxNZNoLlrZOKj4PYzXA/B9NCz0eCFxp+SKAjIGiget48QZ
Iwozptkqd/fzqQolmpiS0I6LhGlV5FGCWSLcE14XtZqPXVdVfR/Q7Loxj0GtURU2
BB5X5lca+cavvXLz0pvYsSCOl5TJoYFPAvHlUligfeo7RUwkPNOlkz6w/dhqgeio
l5RG2JePpGUydHIja5sJKBHpgZKQmVTkK/dIRuyVGD2imIbYnksAU5Zlq5ngbQIn
bD1RPs+h94fYLPM8D/mZO/bNvP3VbMic6t1m75qK7DXHYxOpoL1Fervx8wv9xWTZ
RYCz6dnel1ZQ1RR7ivwgGv3KpePTcjdS5/XgF/Tszt8w5gMMo4b8sy9bPMSstBBt
fV2otkXILJGikPrCt/Lsg1cYTRL8Gl/lInyIGPmDqeI5wWJKmh+XvG7Rv8kuKxl9
oEPDVbtpbsYxD9MPnqzU6xCLT5xf0X4QMtwqfUDZwYTQvGsZqEVz0UQ9t7Sq255v
FX/DCD2SguBSnFm+OP6Ts2pFyukweOi75MLaSgnOGe4PYYehefRUc6tqusL3RSRC
B2Hx9302KQYoZWsnuT3QBXu9+1WtDidoZ0R2efkwnBbbGqAyH0mCicpAO2oiRe9J
v7IfBCYkqi8L4YjSfUvyOA1Estw9OM2q+S+oEXy6mwUmhMaNE3TaQ7dhJ1Lf6UBa
tDM+i/60SDLgsCuXcVsqmPOlL8wUbElio5DLpampkpy18I6icV1FN4V1jGEAAZ03
CV5ZCtMTiY50gyvf9beIWkC1arXxnCYylskNRqXhAUNX3RkQodm5n2VLQfN7Oxoj
KQhR8Z8QbLdqMME43Mrzdo20o9wON03O6PYNSjKvJ4x9uLv+oHJ2Ud/ghZ8fK/bE
4sBMlwd45aXw1SPi3SXHVvRrGFQJoNn+18gU2OoKwMTbQv1PKb4mi2IaCI8h5NvS
AZL3G+zI6i4W8zDh+tkmySCQUz1xO5wWLUiLXoKp51pg7zaGRWeZwoMbzafp3sD+
AEzWNVbGUeAUnHJzyd5V0lzeZ2bYnFaPLFbbvnjUFc76iDOPwKNsVOk+MHKL0PRs
OHL2UTYQ53r/sBXlPiozZZl0zABINad6p3Y3YiW7BX+LcxZ3FoMyP2hVRDrKcg6t
JPF4nBuqnkk8TQ486NWo7HEtYehPSnE0CytNO6gEc82Prp/15exK7tVT29X6qyHa
2fMJg6gRyjlZ2VNIbF0UxKhgE4MlUovhfOuYRiddpw2NVV6t90BDtVW30EvL1PiQ
WNICbQZp/1YUBFPdDTLFRcglwF3S7ZMGnH/304cRqykPYWAysCHuWae4S2RxIYFv
9wnBtYF2KO2AncfasaLj2/Sia6CpTlMnuAH9/ury0wQCgvB/3FiMw2aFuStBAFa6
rg/DWoj3U5PmvWpzs0TcWaVw9Id27ZEz+ym9+Akluqx8IUcR8FIrdOtC7D/X9G3D
pLq50EPzKb5cs/0FwC6/D8WcHSc5otM5hT+D8ojDqNZNu4ua1/XuPRek/uzj1RNh
zFIE38f2VPjG/x0YpVywdFNzmnSAEOyf2pCtCzBRKMjLeZI+n//Q1MlEcPeNAQH6
Vi/lOAC7hUH1IssPkJEQsZwkiPY48GnJiAfJBc+X0xv6XI0IjAYfNW+0JGIfQsvM
j5Pyfs+Bh57k6CCprTkaDSSJww0O2NT4TprN6ueOR6AvBdoH3jNSDwnhBsGidq1+
XuyXdpELvCy8pv6juaMxCK/6JhUt+8GSIbUrhU/RzIQSCPdWc4kQ5fM6y+rPhxuA
mEjD/SANa3xQS/8m6apfrO01AVouas3Hy03rRvkL9uQ8tpAujJyYxtUSIiysH7xh
PPmr28vPJMzsCjF0LnX4E0kqOAQia4HjHZd+6udbJa6z0TnVQaWfLQ3p+CYXVek7
Anegc107XLPKW0c40XBhXVMfBT/fWOKe3j/ip3TxsrpIBsmYEw+aJgWo9wIs4IDJ
+Qz8XmqORwsSHJK4tt1mv8L37JVL7bvP2kIxPeQo30Y3WAs3TUcl7FxmDAH5dXiq
LSycO4WRYi6vMur1SEaOvsAVavm/phMgsiyq4Sc5RtGQ7C1FPd8folh+hpSOlw93
27+SB5aQCSsW076vcU9gYWEBV7vrT6EVGczpSp4AsFZp2tYagLdD9vHDFS1EM/1w
VPMl7jfUsIPI5QCWV20CxH+A0RoD9if/abnb9joNZwDa4LvzEuFwxxwPhW7Ub5vH
D0TjIyWPrxKs444ytEbZFwLk49iRnRQhaOdjk429wbdA/BYBzolX+Akw260FlSxC
6qOI3FLxIXVSd5nPuCk8c/VuHGNiy9l0q69ZcTIC+5ZSrixwjxWmn0YDM34e2vcO
JrNpj15t+Lh81RRSntP06OpzY1vjQl6M7SLRnrDf3f7gAiuEZ9FOmT+Oz3yLznQE
1RsPGOQNoRz2R+MIZ4J0WhsAtMJr6u/7Vge7hKXQ0bc2w9Wka2UoCyJgZNDBncev
EeYQJX30MLEdbq8Zq4Agbjy2R0FXGFCjxqThfNaz5w4P3sYqXqFk+VqVdV/3Blm6
T3qHoPlj2ZBL9dhULrcAvIJXTSbSuELhKZKPu50sVteWCV5a14unDXNP63ESpBvS
n212WR2Ac7TROgBov+xMNOjVNnmICEh5fQAOoKU3DvhZkuvksJqZpMpT6T9Tv4xZ
21WEoJcy2GXnEOaA/2MSViBw4YgE7yGQgyBb0LvVAv0fAlf6X4IahfLfKilWpStT
BohkPnY5yhotOfuGDVESFeV/OFSH8AryqIi/s0bodMXTdIge9xhdB8RhIfyJjpTh
E45bEzbJ1ULBBN0vL5G9FXPFdS8vuDuOTl8Z9nb3n8jQzY0a9QQmqLeryHbimcrI
9ege4X8UrEUKL2sacWmeOAnH/mi9LzNNyLrXxzGRJsIhPuO42mSRbEi1pnnkMn6l
ejBRtlsTrwJCqjajTMapGXmZ9Ri3x4mFV2/D37NahYrzN6Q79uG6qd2dJWPzVMCq
BwKTXCLGFq2dR9a5CX5Fk9fFVxUzDZMpH6vhJSieCxWr216N6E6fOQGeGZuURwpH
qIGzE1zwBKiKR15WRh56FDVlxZuiNVfvo45BN1x6ZCzMw0Wpaq/AD2DoiZhB/Udm
df5bk3aT3Bgq3QH9zLiwj9ebDQcAccn1L6++3rdB2BBwl4WEX9LgU1hYgu6zNJQ5
JnYM/1Cln6lUBo5eS47DSLfDtRDQtzTT/vzlNt1ExaiDcsbwwWc0dFs26pUmAhEz
si5R1kdhxvTGP4aUyirzalbBbv7hCgi4SxPdrFvbluQwf2S70Z2rHttSP2pLfOch
SCJ8fFshvzKfdASNQ6gboJmhbSgEu9fLgX7EwXEabwcCXCcCmbczXR8D84gP+PQU
sEK7uZM7UF5s5k7EV2RqBrf/htxL0GDx+kzDvxuqsctNuS644DYworyzrWyQAGxO
NwV+scSIEb1Nu+scvq7vsSGSlVff2H+Lp5MMRdEdGTjV8A2JL59A69L8qUvTSBlJ
i2e0v7rSt1VBUX9/Zj4cojyanfsalUncpnfZ8vSd/FAXd/T+dt9fF9/7ivZvUP5h
1WtiqBlXggBlFrV82OVH1V11O97L+D6XG2ZK3SfZEezpUeSYUboLVDE1N2kgpAng
c5N8nPhf+Xo0HkjoAnB7EQTHSdtbrQdJGN9fmLYewPtf9GcbyciA6B/Wu1prFgxl
wNoUUzW2/0KZyTZqV9CBNEK3id2GgFcZdBbK8Z9XmWBzyNc/IDyRgTr+OpeipXyr
CLiWCJ/etUkPzLrv+dNAWl6zJe6PgQE0avCqm2sJ13FIgIbmaEirkOaByONWE6pC
OBzkQyihlCGHAWtXuvXXuB0TQjl1BwfAsuGldIyHke3cj0eaXsZ0SVAp85l4bQWQ
A0sFXKti8KQ90HzObxeTU6CeMM285quOJwBt4UnuM90mJOYqO2MDKNdKKZYaNd9Q
GIQ7CgEiDTogEaxYF9CSUozZg5MD3PA7Pdombn0csqGSk23A1kx7WxaCH5c8Xl1Y
cA4h2Z0PRUTgKQlVT0eEsXbLhGlV663hrsXU5ayUcqzpPXpCwMRtTxJC1J9Egcs1
gEAWLOExG4TvLow047uNWz/gjNNYVX6UCxQdV2RCibTx5jQXlw2cuGRYfsIVZguw
jOxTcNJwo+tYLbZl43k6xZqYaNyRkL8UgnMKZ7b+7f5IatfWSbejT2s8D7WsIPnj
kuWG80a39T+02B4g6wZIYLnEi+XcBkeLg9hvOax2YZLeoVZI5IqIMAi3u3INakgt
qGwA10MsqiJNKgEQBExCMWrSOIYWLiAMoNYmKR0PDW4VZ3KQvEnu2bKhI4qSMZv7
yF74q6Z6tcOl9SHLwdN6lTN4kX5y9GBN+7secCPjO8F7qA1DKZUkyfxb/hGYmKZt
nJU4OGOaNUyRhvBQ88l7uLOY/9lyhf+JP5GYVmagxqwblCNBemsxpsRFSjuqA9Lh
/qYR8aKr0iJVZeSBr5ZUU0pmHP2qgM1EZ3cayANjf4tTgAev4cvcXq1stQoctffg
EB8m6jaU+WHa4CwPpMsRWctPl2aW7cOezpKl9mvy7kE54mfkyHjDBAZxvOJejyjz
mPtQOkD21zraJb+sSQ1wjJDkwIZJQ/qvR6nUPXQrqnb+FZC4gTSJqzXI6xR8QoJ3
iO3pPUEy/KXGut33B/Mgp5sP2LW9nnFxLJJHgZxyOHNu7uIiZCgZT+x8xcPsiVNy
+LMSlPxSYK6E161R0EbWUc3eHY5dElGau6NhRArye8VljTAnzDm6okhOm9f47yhr
NhE/I8pYlzD8G2zcoRfp3HMAgyBasF1ABHwx9y+xCXynNgOUWdQU8tMTAwk1a0XH
opN0Ol7WlG5mszmmgvwvssTjNL+GVO3j8uJV5uLc9ZjeBEeVfIMdIvInOginJfbw
dWMHjO5WHYKN9pLAIToQ8dxu2Ad8IsycOcorbvR1En4tt0uwd+AYMuvOAUuTfNVf
7jt4ZfLAUbheBUdDWD3l4/vjfmHb2rO7vkBmkHnxE0S2ERtY2FNaqClk1a0gCVxl
6Qmg7LN5McQUTiPmSu/TFkVlcg2xT0KbPtiO/VPtE0IQM4HUVNV/BmBJOwVGQ+Ff
Iq233ow1GahmasVQVGEBSVgSZtEEF30Zt2f/C7G99LE9QF2dkRg0S+XB/nB71KVN
VzMbd8sOhfCX1pt4CCRFn142aWia9vt2ZoDDc9qbc90UWxzFw9dD6neMdvJ5FU5q
mUSHVh9CNFJS+UbkRa+9CR4yrMItTj1kZ8r+pkNgp1KmiZs23xucOX5L5rM6THlw
OuaXxNthJi3kF8FH1iKDAEnyjg+AaVET8pubMJ6dLoPXO/oT2C0/ufWvh6iqHNm+
1bTjRPLzdaiEpul3/j9JZGVoZB8MSld8YP5Ww3kF7uzpM/GDRO+o7bsb0m12aHte
z7YRvQoeBlKWMmCd5Uoe07+28uRBtrNFCSbHPlDP2SQgMVt8xwe4A/wIvXG2/wib
nMyA8fTLXDRzS0UN60dA2nXTLkPIMAs+MH9My2ooAwvPjuEm/zmXHLtLlEMGgt6r
RHUzWZbFfSZ96N3gmnrpAhum5JQh2Ch7hYaYh/0gpyqPHLaiineDCoEZMCBY/vfV
X9dQrU31oqgVp8J7cWipmX+HWLTTFTPlRet/+i+I3VHOP6zlR++5E7Yanh0bG/+x
j7Rn6Z39mwV2c1BJG9txfV1zPKHigpDirstanz6X571/5ckTo46FIgFuEeb3TC/l
A9J7O7p97cq1UOn1fqTNvPM3rmdYU+DupjNiDVZInT4g1BoPSHk82wtDjFPXxcd4
JYncUlV3slMf8ec9hEY/sHXyNShYB7VpBNZ8PFiIEg6sQBjLjsKPgb9zAx5SL2Es
MB0xGFcWrFOEs46w094w9rXPcRGIyDI/sqRfsg8UYQoKa9l/JZnmMHO39Zo9NKOr
eoNyfFB09N7+3fJ18rlReNcFVz5gGcJ0X2xw4QYoFuNHa1CY7tCaDJ4tNdL86baR
+xJZ2mJDY4BkEK3ZacxGpTZycaLl+/TMLOv4x8eEB54K7E8sWfxsfNVxyTn8gB+r
QVMhip+MgwqvBUuFv5hgTtEzQ7uNQ4hiNV1/7R1AyRy9xXRtcA4Nf5I3iPhzpSt2
bX1f29PnnPYB/K68OVUVt3L5u0NUdYzg1UXF14XTnLl4eklTpoEtZTpe8lcoHMm4
oeT+G58NUg4yerE0/6eUbgTXfZ52kGeNyrqCjWI7HMYhcuJCGewIYRL2D8pXREj/
1q1d/cEBrARaCgJr0s4Ed035oh5kPg5zItKQBQO2TBtUZ+8lVAFmNtUruULDukWW
lPc08lPqDrAsntMJ3W7jsn9KPyk/VFNvEbDuaQQzuB9Awv9r5px83CMTPzj828RU
DRIylz4serZbo9xZNaai4yYD2qdn1Aqy5/c/x2H7MaXzDDqYE0cLss9OsGsRys74
Oj2xn04IazCAC7DcAH1u2g==
--pragma protect end_data_block
--pragma protect digest_block
DdPccPGPmcvaFlrvO4BOivSxcgg=
--pragma protect end_digest_block
--pragma protect end_protected
