-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
5GC3vAQA546x/mttimu684Td5oSHOtCS8s8DnTNrVurreJ8m7F0oIVXBwexkn6nA
fk3E9rAXjCreo63ILj3WTLFtYnuqCSXLtktoTogeRn+QZ0EXU56+TGn/9zGpKid3
Qm3BUsV8gT4oQFNzObOEMywJwlAg41kGHZJ8hk7JohT62v1sx3Mmmw==
--pragma protect end_key_block
--pragma protect digest_block
NtYZLIzwkCuHbUXYsVnBLc2J1Q8=
--pragma protect end_digest_block
--pragma protect data_block
cKSCMz1z8U/b7c1Y+M6X9jxXF+T5S0+C39ccoohaExEKHbKwJfZmiEX47Ha/Zeje
5CYYgi+5bT/X79+1Dv/0vuX43mB9hl/PaNKYAivgOU9mm5K0DZa4glVN7NR9nnWm
3RwZ91EeyNu8EwFguw1M9cAs1zf/gDMcFSMTK2hEUqZVX6lQGlk8z4E1VrjnzD43
B9rKPAynEE8/0AePDTOwucrwFRMkQfG7XNX7qXsojfCHY45pcqH1XIqaQxxeYg2K
gJ1Zpf7/SggFfkxuKXbVZxCSP+vQJGKbYpc3ar06O2o8sk/pBo2EpyjCAGmC6uJb
41ioN8oxYELBGDwaVwsTSGW7BCT3wWLV2yLKEql6UQY/WzE+/0hROjCBv4ozaqlJ
h1ml4IeiNxLbCq0UcdkGBqrKea/7DSAIVC65EYKNlBNY8P9qaw8negHBS5oz5wMr
gONXxv0W5g/glOmXX79x94UD/KK96rRqDUr+GUk1kISqr71V7iDxgFCPX08fVGdQ
Fz7Pz3omxuB2Cjkn3V4pDFti/+nNVF3UZKpMs7DtMrwn+v04sukEezDvQCwqecKM
Lt99MZs/wPwy5V3AEwZNwoyDdS1PgYlwH26Q7rU1+UPIrbJQI6Ls5/wET/muwYpY
8Xn9DjNJ9yjSLGIJBKt/tGmcr1tZN3PJyOOobFxV/jvO+7nPzmQRpjKd+VKIlCdM
uJcIJKZMSckjtXpeQG1f6M5+gzPE9KdJT2WwtQiefYkKrrEn4hFfGlfjbHEiVmlj
cNTb4w4VcyJXZpC6RjlbtF5E4Qbobcxt92b5amZOJ7op8vFbZTsxc/xB/DCPSKqJ
6g1NeGs0bZswBj1VOcaJHZDS6mN6gFoaP5AiZYorlCFv0lFjQ2/YxOmWK5efPEoz
wfLLm17tu64mBI1zJW0/dZMLcEILePknJvVpZi5yOjzQU9QeHdgTD6+z86aoPdZh
yyxGt3Jk7Z2GZ9oOOp3CT+i6vGzqYCiXAASVUBt5ePr2dMNSOTj27SNHxUxF9PDe
4ExNdO5W1/Kdvw7CX5TckAD+zDtfuhVDA06B0EVtC1N71ZmkulRyQyrHrp/4RhD+
FM409/TeFH+703Ccr8PGqmXmwCLOQt4Y8PeZC5Rph8XZanKgHKlmMTWSVTQGtnmw
+Y8cYw2nxNAdz2YbVvzCgZrLFcOZ6waqA0vnNsEPWIII2+f+DDBfv1kxRRHt7FtF
GGoHJLmmZegUJlNHCJwddLVhycydm+tTxGOketjwmFnBj/EP9u0Tk6JupBBEz0UL
20dw+vPCFw8dy/fqdaI3R7QEOiVurPQ76ft1zYYnEn441FqEJ9gGxhgCdX7ouljx
1UWfqgU8mxCXdAWHVEbgA2tiO1zO1swn1ax4qrVA2at75AXzLDgKmw4dRlzAhvY/
0UNYvDLqP6/ScI5hrwEsrYHC8eaLn8hMA0Q5VRAMsTRzPRFybIqfB6wDv+kRwI+n
72MRo68JVTCzUMTRUPf9Vdd2fiH1nw3UuPA8gL/OR35SCy822EIhxG99ok1YkPTh
bf8JH3JTVCok44hNfEb8hx3F32+hHEs8gKq662ZqOJ7vHNxrD9gAzIiRAXNO8RhF
wBPK1hyKOtDr8HEFHpu7SUItQCvLmKNZXplMesuWxXx9PuPjRl2QL+AVhAeWgrFJ
7CdSt1XWZF2JD+ste8NxL4STAJzb3b1AbsDabYcYl9bUFRVvZ0pK2NTy7QHfdA2A
OKnZb+varrFFK6A6qCY4hvADb+gS8UBiHLTVm65JhczQx9UaXlnTc0d1/oev2zgT
pmrKdg8DKXoQAUn6iZEPj9HI2tSL+cTClao+ePqFPHqANxsTQnSjmd3W66Nu39MI
Tc1jYcLiLFAV81PtitTZ4xMrCAiJJblr8+vH1HA1eHMS0rrwFe5c7XrpndfxaKMZ
L+zSP/Ap7rPABw0yqVtW0Qvqy+LVepyaJTzZkkg6S3YT4Gnn3RDX0nqkEnsC2btd
+L0KvDEfhPziHHmAsBt9vBQK6iUDE5cmaxWFX2W7dXrWVwz1K43fmfJESM4k5Vhy
kUEnsZ+dMNAVcmx5f8ipeblgNZc9DJ88xyWXuqWp1XGLKV/CB+F863tO6z8TI5Mf
M6r5MSSUwn47Rn9kpv15YqUrThDXgxyCNnY4k77CRVYK0PKw9suAYTv7lNIv6N9x
yj3Q817b5I9ETADn/3l6sffk1BGWMwdYudMRtPZP22W1WAsYAajn1SYu0lQz9lYJ
GPq3dxF+Fa3MurqlgXMntOOoGxjAs3hg2qS7Wk8hxyb5vIBbdwIlQ8Cgrf0MySJT
JYZssDV9bDmJaAga7k8NlN4WZwmMGeKS6t72L+hlNnPn6mPosxQVW4YZF1MFLc/T
PpUSWtsPmnNonYDwrxTL4rp/c3v3vqq4pHHO/udEJexMtGW9W7NLNFTTJng+e/dF
dcv4mmkQX3i/KNHOEJVk6ZUtYV7rlc/rjRcop4IcT2b31TcMHFKC2tBPX6q/lCLp
5JbOJVrUpI/nknGwxmKFYDv+gc2q8WYVKc4inc3zjnh5kO2TrQ5cTzI4/uXlCGro
Ii2tVDInfE4Ty8NFHEeWix9gkN/xAkqcV/HkHP0CxwyVKw2kiJFYCNdFzBxzo6bM
TEfNG1yuDAPUqC1icJOGYxlOHX880HSvB0pRTD36o/p5d9TuX7a/8u/47uu8CY9V
fZd1+05ruYzuILvri8Y4llWxBbEOO2KhETcdR69iDLLouMJ/0Yh685qGWVZz0PDs
OKO0vbOGCVY4Rbc/aJECV/P7y9qxhFfFsGlGlaD6BBwotncH3af1X2K3maEWx8H9
KzTR+CA1rc8Cp+LFTho8NGFCcr3ho/iA+2Irkj+n3CUfhdZd1DCeTfSxMXejX5b8
i8ZVEpGLaeYXk+QDqmsxYa9KvBBwWf6/jZFRdO24ei868TDCRaTVGh9VgFvhQF7X
qA3cvV1GKHoAjiRxlqpCZjmTgmGaQ75r7M9sCzvfY/N8La47t2aHnMWg6yYA3iAx
Q/8Vn1r4fKn6/4fzAJ5NqIfIJ3lcjAhGzcrwM2jSiM1zwZTjrzH5KanvtuhzkKYo
d3R0SpmzCz9lyv6O6cbI+52vB9GUXfj2gmQNkNGfgu8OMxzXCPYmgV05YBfCx2lG
vvC2wUlFu8HnbqWJ4QK9wW6Ee73CEoIop0fcbQ2SCMHlhTvpN5XdI0kCd1ePFG0g
rP5FjH+OFkKoclCvKu2wtLFV3IxUIZBrTFddEs9dK7TgECrz2ishItAC1I3GW9Gj
JUHRUnczM3RgbAt0ceO0hczFMb7wzwZG8pkSmfcxMM/qom5X7BVNBlSxkPnoFHfF
HloiZC6JmBWdHmnl1I9CSO+4riw04DUUppBeykQboVPZWxO5JDVqFixUHNDmw7SN
+MPoQA8pQdiTGVWTuDV9sxtiGpQxFXhxaGkG1qgdjOOOZ1etfGI5z5C6V8t2m+/O
kRb8UbZA/hnJY5V10uRH1mqpNguOLTwLuxedNvvwNWcErNUqEu3O3PvMggZ+hCbo
WB7m2desGarkGUJlK3xyQcOfXljtGhqGES3HMHnv8N8zU4bfuL5dlCXZj6x2awYO
MGs4fXnYE/4lI5Pusf6FNpvxtFdS/f0rotV9wZ6GQwlK/DDJgMJavGWCR8IYxXCN
hMgCAmR7/4MY6SWZFPr7YhIbQKiy7dVHlXcgpicdm02xYHfy6chVfsOP0J6IbICs
h6pl2tZXZZyYfF+U6dbh8bU97eei6H4su0gmScfwI89yxWVS1RLStN5kt3n0vUT4
FUkBUJrCe33nb7SzE1clm1x3XkN/+TsiYAsmOL1uY8g8l/bjnmEodUN1IC/J+Xut
vFXVijvnVH2n1UtDUxg4rH2kuExoKiceqMdOqT6/Gk7/nx5qMYnOhmWtWjoLGQBn
DoMsO10D/rBekxCBeAXhsIizwJ3kKX6Xj/by2j78cRDsszEuzQ6aUvvcsM+HFf3F
ZRef1Z00FbzMiF5r6xp5B9vDDrTTaUddGHavVrZhLrrL0rTT3bwch6jSKMRMs9Kq
0QaGSXRvU1d+3CNVIW7u+5i6I1bnUEwBwxKxy/RXlpjtxIx47G5OCpHofUVqgRiE
hgcpAktQ3URF+2pmUH5kE6Mb4loiul/xaVr1Uvh2UlG9ouYjMB8zOZizlPs9Nhz6
tQCpHv9hLpUjl0z6lEMSbZCOLVRi8JHuQuzEdfY6YVRWKEYDizOUBcGW11Hr9uxw
8l0c/4SAvUcQSvtfRhcHQiPvgnUoqQyq2rxPZhiouxOOBXnvTJ/zlIUTu8r7OTFM
muwnlQIPNMtD63MkJg+g9h9ksTvQlI09ZeGEVqNdWu+xiEJXwEDfbdVnDDl9BKdX
ypiM5ZMtTBjjQQjq30LwJs2M8PpwC9yt/9oWmQpFqisxY3bvSquN83NvR+vH3Kw2
CRbjSgMadUiTweUPRHhlboqDCoHt37WSv1jcXx5yurhBl/3oY5pHZRObC6LNsIbn
OUQ9mBVNTTlTroQAhiUhzpG81vczfYhwWKrxj7lEZ3ZUzF08U36AIjSfqEvwt6uo
v8izrDNoHp3nEKXr2d2062kfjkYQliBvAmTqQWPqeKCBaVu+S3VffM5z+yN0L1GH
0exq3+Q+nim62k5AbVU2s8esiPwy/8qVZK0Nls7OBmKE1tcL1ch9UHn6uS+xsv3D
CHM9EkwCMOiAJ8H8OGJIeVhcrRwrA0K2qASsAiaIB7MLpLdT9dIdECw9hsNzCD2d
wROR3tarZBpNTjCicHv/qdV9z5ofpIAFCq4t/GYAOh0Va4UAfE50ooxrkLQpbf1K
7TqyF7OsxtTWnIoeQagejGqjKxNoQN4/oe+RHv9zKvsYlLIzSW6XKd4/xxcZ9Eau
idVtYsePLtdpVfZNJL71BZZHIfRPFmgOczxukNsrSom26aTniNyuoi9sGm61nszb
FtuVZRox9TB12njySO0kdN/Q7SlP+H49SAjCoGRNpzo/BsJnWMr2jzAUUpTMj/VN
L524iisApGdC6PL3LnhRmJJ1yQd3iv+kWzyGLlxwf+Hx8Y2l1BAWbqvp2eW8uX8R
YoyPysOpp/cgM6UAHmGUEw3ch27uYOCcQP8pt6AT8zHCgJUVAWHQFqJAgrxv+uQs
gRYwL8WzKb6Obitxus1fuZNo5XEgWwhwlcObJKqxN6h9UmzKBoa5bXKOvL0UYIt2
sy9CH/8zIQIBzLwAtMp9sXZ/95WNdS1mobs4aU8iTExdpVyOznydh8GIl4ItY0PA
PDlC7CY2VF3ctiQ0U1x9iJth4Gy+Npzt6F4ZSTPMzc314zO11/AiCiPIi1UTBuSG
sjympM1tPBNklX9lgGe1uerK1Oe955NdPJRDhAkTnlVELu2fkFQ7vayVo6m79kJc
vYgwViPg+XyAYPDZNyk7/wMakGIcY6E6UJy4Bet6XyV1MUg1oycXVqFSKyBcnhFa
m5tysv+2PgBZQGMfol3mK4uLpsbYLh2ZN3+KQ6EC+dK/XC+4+Babxt/Sso/5zWUl
Bzx+yd53a/L0j0kleyz/CI+nbeus1Ww26/nOHBVV548spimR9jhhRH/EfroaVYyr
1bLx9WkKh2uTEd5o4aRLhSHlsufybF7J73HrF2YCUHJmmC88igsGsAXRYl5klIa4
mJFMtN92lxKSGkeRgYX629GhqOvlmHqwmM4u6rIl8IvPFnMK/BcZDirUq8FX1UEB
hQrTWy8qnVk52x19KyL2/lOD8l9XUZT0rpagraozrlGw7QiKY1ohl2dzH/n6PX6b
BcBoJ5MEdfBLiu0n5KF0ww27T5x+iiIcGofABQwSaoGy0IGxW+wMHj8ozjNHe2Ww
k5SWiHvCGAV991FvQy+DVhXK7/WOUISiR4EwyXiU8oFth/Va1GUtMiCn9IxQw6qO
SohcYUhYb75ZdelckVyjUhWd1IKG4pf7ZMYuMnJNmTCZwudzfUwP5cHF/P+hdt9m
5Bf2OZB3q85M/mjdtJ94UhDEwcH6WIfJdFGBi0T3yJFmVqbgJrU/vFOtXuIqgCVR
oD5uTnkg5jiGo3XYwya2fIYN15NgiNwPetnMAYyXjFQIUZSmgtFqtCV1zftmkThr
/5Em4In15bolW2nODiSkyZtZ15BXXoJxqX06Vxj4d+OgFMBnIv0hahgESrfCjvM3
v+MlhLqBJsCBzEVCp70SyAfGPUG+0O/msTSYAXif9cNUEiSm+Kiye657BWO2XFSF
jlwrx1V0fovGrlSATCHgmNbxFp0Os3/eN0Snb+s3FQeTnvbRnjfPx+LKJa4PCM0p
GuSymak75rz09eTEWQvwL8/XSJbndwFyNYzxUAyWfBvbPm/LO/qKaOdfqrXqHFeq
E1PUwfPGmHvljEYD71hb3F16J7NbhLwP4DmFS8MdSjyf5ZAN71LniQX8TbepZ6qK
Jz7KHj1uY7kK0ULXeQJSRT6Ni+2V0tCCtrY8DUCyqrYgfe5TobXgzm0/Pz04S60y
oHMx3ApG87EeOPCyGZmTot/AXQiU/cRGhQHnPiGJvxOXn6n0gIJWFqPVwS8cZkiF
c7ZyuCFHCouAq81CN9BbeyGtIoFedhblWDUCazOtBDrWGm6LwBscXmI4Ai0k81B5
uh5e+UKLpah0b4mXPxmguIibSAx0ur7+YVcPj8HLCf+ofjsDjQZirezr+dQrL7xY
M+kx6KX4peNnclCfBWqP92LYgvjnzgqSVG+R2pcVw5K3h5LJvr0FTipj0zVgPRZ/
CYwmwAK0VaxDhiOsCvVOYLLTaEmpzhLeDKjDRBvxrPLadM+Hp34vWrN9s8+FKNYg
kvzW6qHaxbHaAhg5gwyL69udswP9CtTl/32T+2/ndal12SzdtzM/YOedwfYjC42R
CLdMuXhqPFty+jZPlsp+2SS7+Twyq+aJ0pxEcIiFSW4RqgRxJkkUC5XrZpG1ShQF
RF6utgPfkXSzzb5ITISG+oelaQHoYWSJBsSLeS+oKXRlO/v/iHzWyIXTgUrjceqb
d9tiJ+1zrtb9NId4N9Crc8OoBCsnJLC7Q/tIXEUBJr4uNxHejr0VUYUrlqzfJfWM
sezvf7rmfHOMFvEwEtKOMq+x0oTGeRRZlCM6XSficiqrUoW2uRmmvCaO7nRXDxLe
VVb9Oem6icSvqgnknNqS5KVwUIdj3b/iL2jk564YTPuCosiH/5v7fcWIjJhmk/az
4GsuFrJDAa5Gr3nFkIh0qJtW7SxZisYJSrSjpYFuXjE118/DrO7CrbSqX+n2TMyr
KLiNLdxfitQyW0MHTacEVPUjGdEwDatVkYUg+FpAJJFx6ZZv4gN/f4j8JTKbGhVg
5of3PCa0Neu9XQxJEk76GOwYl+6VXzSEeffD2T8rr0lIRJPjac5zZnJRZcoo7QTv
FUZ3iRTbWuPN4F7x3TonmPRg3d+g8OJPjxqnHihdzy3PUX0oL0gBv31R7utbvGnf
zqK9bL8820DQtWMtaRHssdlmA+ql/K+7ZGa6ZKDC1WkTd1uWTLpj5XhHNfhkBc/O
RgSWywNduTiCotofMiupTBEN1RJg64i3LCnSSMM8WLq8/yBTWQ5cLhGkrMlYnMTU
n/AQApmCdI25/xKaV62hrxNWwgP/uAvk72rcWa6m2gL4slmpgNQ79B3bhn1bTrA/
x4R382iaRiw2o+1I2RRRvbH3vhjsPUlP7TjQF/XP2q1IG9I7ruFwWHE98nHcJ9kJ
oxSD73e6FbCjQxQhuaped+g0hlT5ng+pAA6NEcS+Yyj6+w7PU5QHoSRkmzHtH1Hx
1RidrN42Pc4UXwauEeE1a2nzkd4/7eAlcrU3GCfIFO5tlyJnzDLx2In+jQtAvu96
PPSpbcP4aoPa1L98mCK6aCfoiaOgyevFynWMQ9iTHbcRHvgcE7kXGBTutXd7F2D9
M9kqZ319kENAHvqOOwaA+UW3dTCnqVDIX3ueGxwKRa38Bq1icwDeuNviss0S1iEI
2GFjFVIg1D/mg0lHq/ZZOSIE8bN2hC8b9vTZhCY5BEnRRbtWG9bjY5N6XbAPbDhL
CmNh5AO2q05W/vngVv/mOPmNpaVXSmpEHSfVBJ2E5UOEHEQLinYuAIq0oxveB/qA
M88aYq2s3seApa2+mjoq3K1Z3/NdpWZC7NRsLg7aVlCJcLp9eJNXsmqjjDhlbSVk
MRp3jp9c/jfjxhprahjKHG6hVXtGkRZ8mP3qvMDoOvCwXlnbDH0w3ICyzVopI3eW
JML8C0ioxfcerV363NSTIa1uZbSJqyKW7fFzcwwUChu/jjcANFmBXay8rSO9be6x
YtsDuUtV1n1rKUXMcNJ3muhyXuAmPPmkdWqwTtf75KliXjYbh3+NuuSnSoYLblkd
zRVRS17xMvd+6IgHDN3sqGeA5Vp3L7yubwirRhZa1puhYffUDQJyudPc8Fn4jBC7
tX7UuDuYGLwsBzxDiqvrlu+gpnfOLlIxfveXmoVgQUsHeMllaAMNvixEuuJiDnEw
ZJmDhbd39u83+rW4ns++N4rl9C/vhv8Zo8mPxMH53+6LeUT33qT4XmjVxyBRkGWo
q5IuiwtQ6hFUET+SSW/MmK4WClwQLtXnljOt8eyoV38vrDVgX+Cpen9BvZ61lbq2
YUxd0nwzLXbPwoOjzAcW1LOp8A9kuv9/h2/5bKfN9fZH4nJQrWg6tS00gPDjyK6M
Z4HuRxUiUC5BqTx/sPw909Cu4VE+e6pTBIOFtYUa/x8LWyLBp7SVf6OOp3GGFWTl
ZNpDFwYobZjTa/7F0ACEzH+7O5CGYVZdu36Nl3lKGVsTfes37xO1qchoVWRumGqC
LTxo3iiapIOmf4VWjhuGgKQtVTxRzJGs4VZSB5ExLlZEZ7IZpGCBD4Z+XoFWEwba
tu/k1s9sRt7mVw3+ReIZeXn7XRWvirfkp1P6sNaTZnfxsaxBpX02UFRdKWeIVDs0
RyZcYDcHfzrRQ1yIgYbzCDCr4S8jqDxcGto+e+LgXLOX9Rt6xjoQhmvb7352P/mW
f2UgU7ywKA+icrWBYP/Nd+vEas+GGaAojlMPvAYqqCWnaWGNO9F6d1tzebRuEvpR
7xrIcNQ7SaN5Z52Wug2jjBhXjhRJK2+WQIDxdqPFyWrj0y7j1RrrdJfwnJpNZmBX
Sf79dOXpj3U6Y11T8wgDtAMlbwbGWkM0TcVoMp5BUYq1VOVjZB5QdWniVsynlsqZ
xDf55itaPREFvzhGEiY1GYgzsKMP1/og3OhJYt/OwE4ZGYoiV+uTMUUO5p7fZ/tw
nBiIgu1bwYuU87ahR+wW/MIs0U7rfRKqVqoGmRkfdESqaY58i8qpvpaisbOycpZz
kVrROIIbWbKw0bUkpFkuRTwgkI2Bhd8rEdS/msBJKc7kg9xJXmg/lp0p6LgCaVHP
e12NVmjYoyjaLe8tYWdCz8Gbkzx2dBcK3qkpEs1JEUkQ5988bPGArSSw9BLlErGu
Sji2vzYgV/MsM3XPq/GQh43PE7KFCuH/p3J2LdLbMK8tv5+n2IBwYmW5GYxsMlFA
ehh9BPMagdlC4fvkFjP0w0fo9T1dNnQ2i14L4I4WkJ6Iqjmtet9k9OmIPdfnQTep
23qJEKwqnrgNjEYFNCeQxfT3fj6a0j7HJxhiBDDhACcifXPZuug2DUFzHsQh0E8s
D6sMjq9lH7xJAX431FnaDleNG6tE+MCoQpKhjEqD1eZWcYvjf0OqiwOUrxx9Mz0H
qX4ggNfwHWC4jXkZDBLxZW2Nx5pGWlcKBD2zfOL805U7f8W72YdHAc+QvneBs8xv
a+OkBif3qcMfhgw3XCcKHBAMpWZMvEzrZI5Ja+nYO/O55X5diHmAXQcu1z9eNAvX
H0yVTAdq3nSsJll9ihZ99ocuIhGyDvxjR9lIMugPkSmTA5zAXf+bv7U90WjIRnEd
BSmzPM6YNXFCakvirB8sXOr2YeJQ5G5aGbRquAOyFtLj90JSJxh+BQaXm+PI/47b
K9SNhfufhx6u5jgUsOzCK3GrIg/zOHLRsTp/+QZAT4PBrH4uUAbt8pcnO08b3I0G
KISJ+rhGAyjjv3fWdzK9skz39uKrWLyJSsRXM2fqIskiLVrb3H/eWXUdfh5G7Utr
Uh5f01U4h+OKUbPcEXomlxSeL34fquMgwa+rEesloLlrwg8CwibQMyx8B2/Yl6q+
r92ZmrjiY4KxIdx6UnDFzkOlXC9GrJFA7T3aMm18cFEWNnl5kC2pe4wSH678AG34
onkPxoueWLLCd63uUhZIKSE4x1BdxgNZv6HlbhFj/7yp1ktdepzPaywGuKVgYEdB
RcUjyU2tQoE110q1OIU3pty5bk7Tm/QgllajQt1fUlIZyOHFgmEHeWWGoS/wNbiD
lMHKi/0IunbS+gwvUyTdEznM2JZZrFcxM/48CJvmY+SrCgcQvUi/Jsic5tJiwDM1
CnHmL0sv6JWg+B5a5sH6v/OnbWb8wLW44lDTei3kuqGcKn7m48IdqaTiBkEj/v8k
kJEVAztrNuNaVYOBmlGw/TZh2YuXEXkdmimKHnQ4bED8x4HZGyLAKfnL/Cdir+NR
fEpAeN43Xu7iiVWx2NF8rRUEjUwFqApsof6EWcfabUT7Bo4AIDdRDpTIivmKehqf
j78KWzYlSk/Q3KKkO7+lxAA570ypiQpMw1Etd3cbQ5mjZt1KfaiSS24dIPE5Z6eZ
91sEceXAaDo5Z7V3XMK9HM7UbdybB8kqm1g6HHt92Xy9NInAoArfi6/LEyHarwJm
vHtGk38nvbP79nZeXkWhFKsbW/NPUfN8yIdPpE0vcNPwpQoZDmoAOeTHdwAbGSQ/
XgXSGjAzzQOQmjk50nJ0tzNG/JOHSn6vgvNbceXgLolNQPeEAjtM8c7cWTW0qqTj
mvHb+VIT/F/T+YdySqt+ArDGLeRng4et1PhjoM8g8vzB9Hc91CPn/0dmu1JU3TCB
xZuVaykIVbGzfHXF/gvTDSIjVn5NX8o3Ty234oQMcU7NmRF7RbRIGX4dNJsu7vpC
TlMc3h+s/ChvdXjHhZmUvr6mfyB+OANTBshOCCjA24mA0DjUPAHbstDaOn24qNwU
Y6lLoNXg5QKii4YRt0oKHoToSZPbmAyoOMllIXQhZcZfTDTi5LwH8zoECti/L1Ub
vYHQ46S20hXJYDdKNvvAulyu4c36SXhb9QqkFcKx8XBSJ8SfTvGspmT5Woz/4ag8
CKS8sXnxbMR8JJjy+muNF9eywGhMs+j8FfGnPDWsx7SfcAfhsTtC6XyGwaDfNPij
dWgbnjNj9BPPiSRzKoExEsHe65D7lCAolx+EabZLNgjYE11wt95WYXudq4lpjutA
8WSCvaOyDYs/CGCgjqzVBu9Q4VmnIG8ihXpSSCVn08fwWnHMH8/+ztlPRk7FkLdW
uZYAEeSCFMzNB57typGCw1lPJj3YEp1ngbIixQGccRpU75MZzLu/cfiBmwbuaYKi
uMxSK5+0NByZQPY2OlajM5c6QmSUEzifFv7mFiXdjj1bbKbie05ygP3+wVjOTEHE
se6hg0kDgJf/NWgjXkBpJc/1lgWtyuDJvhW8qOIIAt/UbWbgidJ6gEkzpYEnwRb4
yG7+LX8x1GKJsfRhCMtwWk8JkV40qBmKYjCJBDdv9oeNSGnXYHc4jS+0+qzwBPI0
jrTEczrZy/ksFghdgc4pwK59xrRen2FvIWBXy+Sv45Zt77o7/kehiHdlvIcdVuJ3
8r4xotPzySp0EC81487r/CAVxRiatG3gy3rLSP10BV1v/3e9qsW9YOopwM5gD2Zq
4ZS2aVy/XRrbh3bEL6e/UWt7TGGvOgzwl6Kfx3cDrg6S/9VIi7uv7MAZ0ORbAfkB
dNv61QtlwmPJv1C02sezVh9bD0VEwuQuOIb1O3TfrXhcme/YGpNxGW39Ni0R3op/
YXmJO9wMK4bNwDq9vKg96sZh+BHSqDobVrZ1EMpzdnOWbXhwGBz2bso6oxTjZMSg
pNH1+XV2oziZoq85S8uc+n5/YEuj5/6EL1SGQ82OT4YaA7SZLhpq1sKkQp35gDu8
ES8ulcOrUmUpSPj6jPyD0Hfc+YWsCBWro1uZbrAQ6mHwC8jJq+6baAhUnmRdCFZG
oY2RalI2ZqDq49bMDXJQhZBONokPzWqMfwbANjes8WMW3dblXF2F+1xfbiJs53uS
qEsjM8CbU69tLGG4vTqEkHePxuoWIZ9BkVry33fJga7x2mXeQ9o6u3Pz4wyRQce3
KiCCRUNzY0terEz0NTyvizmhhxKPk1g1QvIr4RNdDZuoBZmQ9PmD4q09rrH5On/B
eUz0EG9wTL6oajePuaf8hXo69HL8ESZwns1lJyMrnZul5dI3hyh3BrQFF9dWY/mh
AdjjZKYSRiv2sylWLZw70PAOEIBRylYzCiZEi+ydwx4aZsyCKKVNZ0sI2BrP8z65
DtIm4sMXmaA9sO0MlXe3i7bYNP9w7NU0C2n/utNEQ3BjlNhj4nmqDaFP2d0l/h2F
M8T5p3iIhXtdirzHgLhJhPCjuWqzorF0H2CilZ2y+t0B5eyPmEcpx40tjw/eOVoc
zoZkYWExr6an6mPdfPyNfeOePoPpmaDVg9Wu1jXm4OVtz6+qVU3TlwSkn2Uex4bn
tR28zenMZNd7eWmbAwVU6bksTfw85zHTHGKyzwkc1oxS5HXNs1MSIdPOpRaJPanS
sy+z6lkaN2zR7f3vEBjzrlBPbhFJEmuVKoqlw9piCDzv5wwkgaEdSYm3HffCw+M/
4K7blij5bfDOTLxfqboDUiYNlIYhytNqKsx1kRr3dRERiMC2qlUfKZhZ9rsJPJoD
K8EiGnzLCtiidinp7ucexe0CKIzGJr+Ag4UpzPKpVersABWQkHPXy/bgbxz9U2br
GT8I3MitJHgwi50LdU5r9TUIRA887CjJwqpzw7ldw5duF0jLMxPd7BAfaIZVJQwa
UijidVY8+uH8avos+VkwCxqaXrs0C2nJ5kaUsTQ4a/+keMmmEgxJ2tuhE9SG+FVY
4ZeexHjI0d8cyg6c3u4AwDOatfc68IRe3CrvVmLquLAwuWuoOPbc2o86PBhLCioq
bV6ns+O2Yc7K8cW0IK9ONlRwJcnK9M45d5scRapmYD4nqTBnvUs0zacZwCICKAlT
1AVFYtBX/uOM+IYVdKFX4XrrUVvqVU73yuxG5swERcA+S0usoHVmCwI0C222iAHG
uFtg3IaL9sM/g03O3/GiJ63CFurELg6hzsTxOXYr2gslf+9YDOfxK9OxKdx8kIAv
BzOcEI0At6pPVKT0sBsx9LtJ2mr9KIOhOWm7ZPSS0Lbn774+A7rxro5pibvIkwEP
k7mVksAxQOHw+3KnSnYGy4sYrFBfiGtaR7fxWM3R4Uvi5VqwQnBQC+A9bv+2Z91y
4JtFDOs5NOEGabI4HK/SmtZBy/EwEdSkYvrkMtwGgWHltTVhOGCdMEW9EUOPldWG
zVJk1EVWCvV3NCttMzb0+Z+ZtpoKyYqp+2Zn8TgzIqF6hxTtOsDy+LJnTOkR1TPI
21DwoQJuVVgZyTnVQGhmcNtCXNxHLWWjgAx+GmM8xtNADxFR7GW60G3FcSkOxWO6
jVeUTstIwZW9VKYi52FrifDnR93YmfmxC6NrS98FhEUJVis7Y4Ta8SOfVMuW+jf0
UpE6uzumPKcZFEycvyDCyhcSRZZafiYB6zbZ8Rqqr/tjKgTOz7ZsipVKchW3dTDd
6vNhzw0eV6uHDU6nTFt6qcD/5oqwvvBYMiiBcbYzW92ufl5HLmGP8vEt19zwCVXs
44iSOWYgbuPkkcPM3OQcLfw34ofHtZxSm/eLAvcsCtHaejL7O1fXQymopN1/1cQK
7nZAq7RgQBL7IZY5EBGlewB1vwwqPCwXkK5gtqhKqg4P8joxbxLd/5YJuHxhe2Pl
TQmSzAhpiHYZwuGvk10T7xm84wFQ0h9yhWb9fe5jTMJhiHgseEFxHjaEwzYWKYWE
tvi9gCeqTxcaCpV7HgFXJgoM3g2bXHQxvviDC5CP+BVxqGJBgviv0UkoKPL1yzWZ
jsJ7IjKpur8X1r21FonQTIndeqp292c6Gr3I4wDVmP8nkbiRFkUxhwulD8MZu6yw
oNisjMORlwYM3EQfxGp2reG/ByhmktVdiv9yVa4rdyCfsKoIjjd+mzv5Y6Ko+tUf

--pragma protect end_data_block
--pragma protect digest_block
aGSCpK0BU0CixGM2XHMxoSApEZQ=
--pragma protect end_digest_block
--pragma protect end_protected
