-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
mCNlofd8PyTBMOszLYx5zJm+77sheoNsxIcI7rIlZ5mBAifPVoUze0qdQCEDCCYB
OFoTUJBIT1pkCAObW2DDGBEox/opwa5ZjIHKZ0GyofLLxHzgWxeKtWzUkdjqaRfP
Nso5Bvcpo1RK7hkeP/Sd+nYfEXhmAOSshFY+xsFHmYWXUmtOOa/yCA==
--pragma protect end_key_block
--pragma protect digest_block
XBcv9uvfHXA0bjbbetKpLChNZA0=
--pragma protect end_digest_block
--pragma protect data_block
lx/29nGqbhI7ztS8cq1MS5awqyoRBxVphf5neU6i7plnRgeWZtP2I9GohpMz9Q79
m1ZVDkZSxyW4V5qzO1hAjJz22THLimorIARrq7LVT/BTgR0AVO253d+esT+jiVdA
zRQxPvBR6IpQjQdOJgkZSbv3Z+vieCH8t9PQeOdo4UqpiaJjXIzlhx1KpXrC15Ax
duQRV4FMFlntR6R3dCeBB2kDye/T4vu6+FTz9mCwsqDYDlEe6muxxOlrI9kSQJel
XQGXdf/SQeNjGJt9PP6yoJJ20nc2sgGj7CjgwrqnQawn16uDYH3u8xDK3rLkbB5N
3uwLaEiqlu7fOvzlz8l662lAccEeAABvBl2PP7l5NZPGDSHx7kF9rcjDRsMlQSxX
B1v/wOiST99rVIKTDTl9HydW4LiN8WxBcYwiVIBV/h2gDJEW73eKLR0Hl/ERlEjw
Sa7MH+H5TyR8AQppL1v/6kkAIRZG1B4zMAwZn+iVva1wFWkKstn7+twW+gSlmLiU
uewYIJiqKty9WXAazUkApOQu9AW451XInbG58uAc4XhuCgg7x5S4CCW1nyCsYRuU
SXr4XEBgScqmfLUShMDpw47z34jQTX9dF0Xja94Pvx4m8rtC53ZbA9eXJbR6OlFu
BO6Inv85Hi65MnTJ7BLsMrg4GT/GhAVqZA+grLNqOT3fJkYy+tCFqhSGc5vs4TtS
ISrmZoqpUL7bEAAO97ZMZ5WK4fU0jvXEl5v3WN1O1ffRWWJhan41B/9/M0GFtcRz
myr+DCCk9no7PRVHYQ5Diw8AfWVh07Mcgloj+9IXEekkGzuuPB7Pd1AwcvFNVAIb
m2SXTQllO3Nz1Vu7VjysRKJmg1dMGxRI6+MoGyWx2wx2SFleR0RD5ZdkKU5fy9SX
QDUaki/vyPraszrHr+amAX/8G43w05b1KUmtBqy2/QDMfMbvOQBR85UWyWH0pjQc
KkhIpmI6C/x4zNWCYmu9X0DTTYTCzBTXIu0OB8NU18l6+5xBQM2am7SO+wJ3nAEf
HU24JhcolCRaTtQ7VKBZyYWgPQSwufRDAVPx6eSvkyARG9Uh8z69QFff6NeLrXuk
lMyWC3GvBUxTcGiZJactRJ63A0w1w2ixy9wBhLGolwZpMihhKRdbQYesD1aZ7aLB
TUALSrovxCAsCLlTevtW60Mn7xmZZsEcQuzHVUMYU4c5f0enaJrdLytO/yW8jV+m
RCT9722q26+/WyhbM6NjifLpuzkrj83VtLJcO4kosfWX+ZPZtk5CCj5Hk7uqm/XV
YajoY7wayM2LnFcbFquYg6RrQqsmGh/o76CzvqLxAUB53dcfb5kMw+WqCnaaKgFm
46BSScJOiR8PJDye1di4mCGYOL33TViXGvBEBp64ZxfI8MCXWwHLaabl+67oYBB6
kKIOUY/diixRljKNn4o1e6Zt4+VT3n2zEPtzLnr+UR8Sk3w6kQdhou0VkmFVgmno
vnwbZK9xlUyfx/tkQpwcamf4+q4FuHieKMDqiyDHFzpWKAnwvkpqpH2gr4O6X6h2
FUWUDgHuHyeYlWH9bdwetLLgP6TU92CE6dB1nYdKimriqdsq3Lcb1UmYwfuJdcgD
fhh3TJfta6TFhZ5a7HszWDDh0vrghN9LJZscQfwKHyIn2xUxUTRHiiymfM+sbpH2
7+aL1Ito6SrRXB1rjaVfE46KUY3ptOyq00lWVak/DHHxZ/jbJCxlAi9xPENZpbeh
OyQ4PSv0x41Z5Uh8FbdIAF1YofbrHNNgc33tl3F8Fsqzr50plRAxZLQyfnRjtiUw
32obkjWhTKAVrvXrwyTR1gvvzhTfhK88cskZaLWdP7Ur5LGl+0Ol6ipv+kUmTaIM
Jbzx8BNnNoUnoETu3b5kGT/i1RE1fMwirpBnkkBHbbqohi3rye2loXZV8OEoFW1b
5ev1SXOXw8cToxQhkSum7jlb8txQmDR5ZdCovpc2JxG0iAO2WbfB7iMZ1RiC8WSU
A6X2Qo22uvvmb5AV4FaUhPJS8q/54qMAmO69WeEq3sSUBppDnGdGo8poVEN6WRAg
7cDs6/JXULF0RF2BRwPIa8TMacOCex92lECabLS+v15AXc/VT46od4mhOXpJlynX
2RzLx3KHMiowiEqjEeo4G3Q6n6fukNRvMUW70yIINa/8Sr+thba+xEY24KwkOEF7
AeOfa23Dcb826W5NGH3XAE8BneV1aYr000WarY5B/6AK7ZmoRXv152tbQPw13uUg
09dHzKgZYbgLpz1AvWarw05zFfdMuQ0oVFZVOCOQoMGY1aD8TA0oPPP1mzZN10f4
rbXfD3VutU5O8sDQ4kqfaEpj6kzuFbLioZNtm+bNZaQBjkOmYTxRXDUnbNnrXIrP
9o31lr0/7fXvh2GoC9tZJYeMNC1Ykg/CNv4MoQJ6Mb2TCJ47ZePZa2V6WSWCg744
5bw2McnMZsl4U/eNeHquYHoOck0BGixG1XkgeIDlGu8H385BqP9PbtbmoASF7FgY
2fp1KNv13eiekcdwtd21TmEYn56H5OZgdkMR8DVhIQGGujqSNv0OeZZDqPfT38xl
cJpEdijb/d+dMcWiKVMTb5TWUhvHvThdGR2LEPPsRAZeSAZA5YfFyO4dXuGhkDkq
uDxFwwz/yiru1yKR9sN2Hh+OZNirtZUPKsqU52e9w77GWy6l58C7es5nH0fnCKfg
KkmMPUITr5PmV27UqFwnMntIrqpMVnPy2MQ3/kFT5yY75IcZshnfdGSwtboF32YT
n1FYfN7vkPraRNmINm7cQUpATcsy8b+Md8J/xmkDlBw6hE3H1oSvK0Isy3An8mfJ
an8c4bK4X6STGwM2FSuq11xLMZQ0P/rhyhsWuGutHC3pmniDrwovvS2WVmk1QTGr
xxI6A3g0strBpX81W8ceZpOc8QlGVkUJiFwAgVog8JYkpR7WAvJFkHsCV+dfmuO/
orFMPztEcQANsVZ7QPqWiK9Rls+BDVLdoc2BICBwpKnvm4ZO+mLvpC4oKrDdJpDe
XP3D4I2kF1Qzb/g7Vj67dGhe0L1KXdjlH8OGBPEUk0Wjqz5VpUIl+NUWttz7Okvz
oliPPIZ8eTOh96p7GYHs6zWorBYdjk6iGHVG38qCYMW8OXmvSHgWsbmHZGUsZrs8
j29He1YdA5DOvwkeK8kyPjBn8PEXG9HE/nVEjRIdwa8K5kGtD0dz3qpT9zNg7600
SF9Esl8DJzhPp6B61iIQc6NrTC/GbW7jbvwSGFRJF3BLhmsRutiiKbODVkUic2M3
RYK3wHGzxpNoM+bVphy3Bj6GjZ+iliETCLzMMGWQnv8zDfYVLkwGx29g1+esWk6F
r/07nQ9ChTQSQ4OmVz5zlO2ZZEz2IcPmX1ln8hh0NEzgA8Zm1Q8VYvriPX5xt0ph
vT/jThaJf8XQYoSCeNAng2zTMigcUgJWouYnprF8IYn2NTnVAPA/EuFiQIpUqzPg
Fvm4WXnFAv1MdAyEfpZ9CMrj2IRg/ahUCSKhc08g+ncThk/Vo4tAX+Tx0VJlLMP6
SfGRKaseh9/vwwhIOXuLEKg2abV+70Bhc1qJu3BRhcVRFOZ710U0IXogpKYW3itf
Z9JIatqd+zeIIiYvlIC+9axuMF2br15wrGkG/GPMuJ9+crka6O90HSBOwDN8470Q
w1s3TCHI6s3GGmXvZQ5s2qzwbdmnOoCEQuANdNEKOQwglt7fRrE0WS+x0emyDwyi
zILXH1U+SQmc3JUEkJN6EYODZjXzrWmO1n+OSir6l3RmlaD5CODPW91wYvTTylPj
Yyx1Pg+sHbnVjyx9deJXwj7AnUTHBZsLMK4oS11tuWhVtWkRNx6w+u6a9J6sB9CX
R52PxFFf1XxKOBj3dRrmxifYkuw2Fqv0s10sce7733xEeNCokrg+q4f6x3ZNzKcc
d8e0cQ1HJBvOBalWVzoVCF3fC74/Tcy7/JOoQQ8gzthUf/8hoYRxReEvqmTczy6f
X4E6vubCAz4no7FcZAVbx425i4IhWU/6gvfCq9doOwndzMEnO2iiASLf4z5YZjAY
vXSSzcwiy6+ACFdaQ+ktg3rGecuvSZOjqZxdINQz+ZMKMkaFXkCy7AXL6H981KRt
FbTMp/ZP6Us8zVrshm1h9PyGUXLjdKF9qNR7FnfPueq+Xq2GRAPR3bckwk9scb/d
GkjGqNUEZeHji3PLh5F9dwJ4Uwd8ixyE49/lQoWnFQpIPULyqRl26qegtzmyRpJX
ubGMPGujnjQhEb0f3WSEzUst/QBzANTbLyQGy2QZkE5gCSQ/RNkjPqIyjB90743J
r2DkazEPx1MI6Cx+CM+pp11sgh4WepaleGveXuLzUUxdt05EUNSnhqx0DDDdH7Tb
LZ/rbPUBXHPsGmhYi6Ilif7Z7t2CRab4th2YTgiR73yBYQV9P/LsO36b8kA4oTKM
KsF9W4Og8a9ycYel05yUy9Usedmdk29jCLhCDOCIZDu5N1UtczyZmufnCmVjh4zd
9JOzQKVgRF4cO6WTLCVyqiK2lP4S4Y/5Ng+TKsIxlrm4UyaThyWDWpS0YuFVjL5e
YBOCwmB2wm6w0gB/0wupvR0gpcHsALmgUyx7tvpKwpEJJEyBS32jASf5p5j79aZ1
v4tFrbhwovrkhDJsyVaDS89SERT3lcUaEk0qf2Cffe8JitxISvYHjazftIm64xPZ
wuQfv85vqj/uBv4Ez0rl9Af6Clu7RUCY8/XjwhxFJcxtqDoOMuPFroGVp1qFig+w
lfM8lNZcpnU6n57iAsj+8NxHp/5PBteiZwAOWyBBYDzyUgHmBUuFVV7QSlbCdASu
5KS28uDZHkom6kkeuDAy9KAwpKk+KfsbBwCkh4Xgl0t8xyl3ZbcsC0yJ/yQOR6xm
UlpbFqzXGHa75CL6794J7dwnrvOmQIzOrTtSRUqi169zRs8vjFodpiRap1BV8aT5
o9EDAj/bGcqGty0ejXK//j0ZSfT9gWd49ul9KSMb0uTG/JXWFnxr843CGjXWS1Ex
1DboIMcMpCGZhIjO5F7Isyj1fho+/OnP9e1FLTvoOZfkXVRHhQlQxgvVJv39I2sM
5M/lHVDUc0aqdT12t0ie0jtfHRuiKuqLatuvRFVptr7uA0psOS43QSQ22cIh/Agi
2a1HFveBgqAc/20UjjpCumNxGB26t0wjqJw1S1/ULtZI2SUffK/2marPInzjyEGU
UxUNCLAdOIXDs5UQyaBek9C3tX0Utzeu/W5x1QnOTCglab7hqHjNK3m+LMglXLbl
OBdRnBdKk/3OF4UVxFI8xxuzPf7xeIIdb+zHss593bqjUBt3hXwxIP2ksMmCupAm
T4VaiTUDKLKIFrCQa0vhDLYkCk+Fyl6fLqlKQrT+992iRkDuYrXjOI4FdoKIioLo
rlSn8lzuYwIWIoadl0QnZ6WC8S2r5Z6hKtOVOdBn6KfNvCm20AG72ZFkoRuLKgbT
V1ZlQ/m/ohA4DKGceR3VWfUEnIl3uVlswuDZXEbQdxx31NfJ86+nhqaE/KjXLpi1
P56XnHbE6Mhi6ug6PZZFKc2JbVBH4psnvHXpSf41+dOribpqhjFd4ZnvBFrVZjLF
jb/ALjsET+PEYYSQIPv7leIRq+99BTSLIDhiVoPlbVaVigJLKSPGMFp2+WsvFYJM
/WSuM3Bluy1JInxLA/QtJMIoW2rjqMTCNWwwuK2WGYxStYSTef7ADwpRFRsGfyIL
YBXft4nxtZy2W61ZygoBO/0ie2JbJMgUhFbSMB2elCUgmti5bVHoEcT9afqmm8Ja
aBiBRjD/KWy75LyJRcC4RYqt4GT9am6falhMX0nedGIekeLoNqBcd54EFKSvc2O2
/lraEp4ARPtKOZ2sZAi6l3iRvY6Vfxi5kj2ivTqphEIVB4YeOqA029H+F1XW9dI5
gm0UYlkbevE1d0/6V4kRfSOeyeiismMCFJNsEBpZAbKQFDiiGMy79PqZyRoobIy7
87HlRjs66zFnBjhtxWmCjPJbstwC8j1WYrJutNfvT8eQ92oYBws8llNZIxX8EiOB
YwJuEmq/PXYTf/2ceIx3IiSNwqwUA+COVdUM6A/7kWBiusRJMPZFHTMkny/n0DEE
Rxl3vLzZzBC6NyUU9M97MHG8EXuJEBYYRej8ckKgg+MRyTOrauXyMVi1sY7vNpUj
C/8BNHDB7h0/gdEcmHfQA4RCe8UaE2uuJ3X5CoKM3OCu+pDWNTDsnW5TY7gFAp+1
7Hg3Oamdb3lzk7YB9y/36yiXA5ScJxwQhGvlC2X1a3gHkxQ+fnCOXK1s7bozjF2Y
BhjFKsljUJQHmgds+Sgi7g7gF3pIxSjkL2ozeoy5edmvw3AYgXsSJw2CX0TcInK0
exYuUhFGPG0P8KB1XVpfYNlSuZlU0omIM0Gw2QyErL2UR64dbbf//GGoNYhg0bZb
IFV3FeHMV01EyHaITd21m3mUue3ANvE8plR2yHTxvG3pcuAxJHO7aHzsc8eX1a2Q
EWw64QlIfnvmp+awZpC7LjTFs4retuj2PlFyvokOMaBMqH7i7t5sxJMadqqLqu+Q
Gj9BqFZQ/9YCkEEedyGKu4Nf2NZtWzS4X4Ya8meE8XGJ3nyZRfgKZK+fpkZ2xR7G
J4OAnIHWYMW6Tpcqg3eC7jZ4zXQh9JztGNpYqQvam/UCF/G1cZ4KLEP7kuFTquaJ
sKhxFWiGpHTDydbZiCdSpy2i+wZCxonjTdKI6QsZVyLm9yC7I2oIJHi1ylibNxcE
upYSeSCxeYvffVgYSrC/HI9yUiORjYN1GudMOxPBgXtaUawL+n0ZpYUiLQjIoySI
8Tqg3Wj5rLfBGakX6IhCThu5X2kFgxeL72WfXYKd9oZn/9MTFauIG2LG5wByJ0sC
vCvaRLuMOk1QtSNk1rgSznE4N+thtN+eSTkFwSazP24ev6N3Rx5wawWSAA4i59l1
otgjERflkojpVc0eJmWcX5OsZe7JSQhsEMuxGUHcmLZDvjWC3+/ntTEVTGzC8SCr
GO1/Cyja/vpob4yLHNUn3ILtw+iUOnGhg/QX1dNnQQlrITtrdD2zwp0RzDdX49RS
gjY54AE8orUm5RtDSC0fJTbxCP+soFAY7Hwxp8XhM6ai+JCo8F6fibGbgM0hvQHg
2PIWPmJO7FQcjrf378YuGG+fvgCjLas4gmIm+u/3YFK/A5OgXyAyXpRB1X9ji67j
0WsYEltwIwNPfAyQJOXgAWWfMKWLEW5BKuwui3UGBK6DryilgwiZMZ5sCYBOkk/7
p13PQUNUVX8r94BHMkaVMHyOMBosic8zi76umxjjG+Xo4H49MNkz3zDKin9vf2Iy
9t9JW5c+Qo2LlKEmoiwUfMurJHFTJO3Dhl3mLUsq6S/hoickq704Y54fr1nSfdVo
e1M0H8DnCTmnLZSfjbF4uCUPrRQSmBGMBT3zEeB2wMfxKrqfW9KXJmG5TJrtC4OC
DaiWTqbzfPcDfL3pAnj87h+yAyokAnWfAnOIaqzx7TriCPO1EWybNZLGUu9YKmDG
e7UCeo4yw/28xL1B/jqQg21JrBwU7N+KgJVyd6RTR9xACrGnBa4xj9JuSBEWr7sh
/gWskKyXPRTaTV8jpzGgS8+0qQYqJplE7t0U6mRWIK5XMG9zPxtUWBVnp/rmKncL
bYxsEiubZvpNc6zTD3AnYIUH7iQ63gKkfHMva+h7LvSSfOY2uu+FF6cgCOc9grVR
W3pCdRdEWLWrfjMMdv0cdgYiCwlsKvCqGjhT8yf0Llr6YbihTFEpSpfZM6AHVe9l
X0CyvGObBhdpVOmRih8OQaDuOpPMLTNoIa8X2+kvTO2q0jTnaxLQhLItTZUURaNj
32BrGSlZGULrDOXX5gWDOMsY70ErFfurwb1lJbCvxsNQXI3eQfCW2HGBg9yAI3EP
LGuhqr5WFiW9IVIM/oMcOnzETwErVEkBi6D3eDW7POYO/ulujSeL/m9gyWA5A2wS
3W6Mdy1YUm/1KFqAmfIsrTnEhIf5ZEaVwFtNnyWVmH6B3aA2VcZYLTb8cCVHUmW8
xBlccJfA2uFcVQCYrz6N3UUHsGx8+K0c4R3fG0d0SEBo1Kb+m5M86zeMJR5ngLDK
UQKKR4wUf6nCMRTl1H4iYd0ce0JyRXCKDhQrn3Th6QP/l4r2e1WBIvc8DEAeYGza
qNnBTpWLASygm/qH7iBWpB0QtKZ940FsFnJHzF1pBQKsubVytTB90cjLyTFVzCXK
SdG0TVg4yPFCoCMpJlUQRVeK8oxr+I1Rw/h8NIfZpYzbfGEXpKOLQGr4AerzeVXO
Vs5kPDWjSySQo+Ig/vfDuo+9L7bnHzF2COrD8XZ3OaYZ6I1OOz+S+/N74O7FmZLt
tASJgg6R9lBAuoaeOjpgtbzzPSyZGxtbxWpvnFdFIklIqGeeDJmDdPA+LWwGwdFJ
6g0NvLcjEsWCqzq38IzLWdOZGhTQQbX9ILTYBHs+AOuRnD2W2hD3m0XnPUdJ4UYy
coqGs4nVvYjYNFaP0AG6/lPyHyIQrEO+TSqxdzSa5rzqw/iKTDtlF80lRImmpCWT
02s/HJUjY48puIdwj8OHYGVltGI5fOmmnRMt70h/l0N3JtoC4GtlwQhAuKApmeN+
RNakT70+TyPjaqxTLN2zHIC9ao6YN/xLSBH8BHuAPQde1xiO5v+WBH4XCCAQP88d
Ihkjgl8sdosmJaKvpoyhrP6en+DfIaYv3TxJiAje5BPHINB320dqW1cLiwCe4g7W
UDCp2QtttfTGquDkGBPrumM+Bs2RAJ8tqfnsuNEiOPTqHqqCs5K6Y5fo0cG8TUE3
FXof/6j8FGbCGM/BAx0uGfwDM+BpRyeguZjIOI/QnHiXgQCLebqmigdkLPpg1Yay
rgj/0JK/8CWFkxKqku8joRceHlSRVTQ7K67uMk5aHi7nGIKuaSJtuDwBVQLCqc+0
c5QBMMPv9urFwRs9exMoIEJnH7ZsCOJ+ucgVQIkmTpNRL2DtKikhS2FZ/xgvX/KU
5VtMa4JTU9tDED49ghaJhRNTtvthIMowaDnUc7Cv8ZD3PKO5IBTt1y+Gj+I2gE0e
2kWPRR4pevbbab7SVjAPa7KpDF6soNI7TN20L34Au0mxcABHdeHxm2rID7RXUf5T
rX0K9mXkpHmexM3leECPnDpGvQrCcLjX/JW0uI45VH4BAZzpmdX67jUjUQiHT255
WS/dvSkPezQFPtj5KD9JRh28wMlGCWrwOijYm6g/1nbHli0MH2D0QzwEr7gQbn6B
sshOpVsphLKOpuTOdRfzgTIGKdIhY5cgbyMLzlNKFeOJuf7eeN7lPwnGjGI691u7
0Y5BB24MFAUQHeabyt11nfVBEEFF47lKKK0K1jvSn3S7THkSlYs9EDeeW9buSMRB
I/r1ubrRCq9Q1M0r0lU8CcIf2gUNIs1i4NDWxXx7iB7quSQnc/do7rweu08Cl91E
xqYiOBPmoM+W9cTNBO9huJ6hOH5qLPPM+4caka/zqbFue7McaHbxFH9hjUrW52lg
d0M1OFyC2dRKvNRaGzFGA23bXickqhu3B9NIE0ipz+IafpgH5QXw4RWRJqEjw4gX
yWrya8lAZyIX2OkAD7KyrFHrfKCgkAgHZfxQDAmG5bDidWz6txX+IqIXUnfy4INE
tCTnDzys12beyGum7ADCW8mFWOZvTv1mOFYJ1N8K4WAHzuDguMsiFBC6Tfr3+d23
779UGrWMKCWllGkTxzNpQ8APju1c4fWYJSIcSKegJOzBa+Vr1M3PjvUnvLk4rwQS
iSbTfVt8vRGtWO4THSBuKzw11k7CXN11WJUtBmFL8aJrw+47AnzLEKyE35pInEKc
qM8jycevx7g1onGonjvVKrDoWHJXrgpQsbLYgIVUIzFpcvCDyoHT3alsE0uhtYeO
GSxEpvVz/eHDPGvFBoVKNllP6UQiR2rG5mvH6/rtBuZ0GO+7acyNi2dSlx/BB5qk
dANmOfSBUmcvYydN7Mp52q7Q/yZxmfG4Ont5DrUKV9ctAexD0zuc4yQ9n/FnHKDv
qecmyXecgWHq9pyy99znJqGZ1hOL3lRL4d3E7W5Ikhp776FQL5A4vB7buTQL7O1r
NuzOLw/zJUBl0IkUNYyos/CoY3yx71vp58ktZu21u8i5ndQuhAEOO5mKGSPLUmrE
6YWF7AwMx2AyuIX6AFi4/QUuU+8yqKZ2RQYj46y6VbyROeBPKhgvCmwn3sUWVB6L
Fz+BSa8K8t3RnP7pf0rQpI+Cl8gUudfmiPTnkBK/MpqnwTQ3ggvRhwosz9gkHwhI
1AJih5NQgrh0PzarE+i20meNjXQRxbmFKFaYiGW//v1U74z++etCmo753AnNGwMa
xRiC5vLu0FOpZlYz3aywFQUFtpc0QRhlDl7YXN/F1dueo36VGf1JdekPO0Eg4EZ+
dQaDLPKCF3tIuFEAZTibXDS6FYHynGg/Qj8Hlit24HuJ04S985qrQq5BlvhWQOBu
DFE0joiYeBfHK4kHBYouy78b33x5QkjOb5RBqMea5zXoVtjojqTdh7UzZdOMg27y
Y78gP5TXETWpbT61+hidb2MfOJWB92MGmcOy0d59Dv3kr1LQFAhpVGvzsPGb2XNi
A5zT8rCbFx4VBcI5WsPlfLxgFV236pejmi+FWLyCAOkovMw5kJaHZuUei7oovNhp
GjcPYdm1m648XF0WhROSmJcLMP/V11BEK2s4JTysYdimSm8ZyzTEZ/CgrALGn7c9
OwLpvzJJQYTKyE2f51kujkWIaM4UOqTlaSnW9p2VGkuhzenhfwQkCGfUgFoxuaQT
EvTNyjVdsRHo7yTJ9ULSg4b/iH4D0QCuwq4ugxTLL63F+6Lp27lLPlbWfhDsiZfn
ScYxcBZlcy182WP3TJ3BkJl2oUfJ9jEjOoeKsqo+PNRZ17NA9C8Y1caI2FNDXDeL
atx0ff8uDKNZ04vnPGjNnsJ/YKwJTT6ol8Zkjw+gTPxskXOuw4ibqPxjT73MR1km
BNIdJL0iht4DCoj9zxJDeRh55v03ghQPOxkqmJyz+/38g3deJ8ldAmxVjor14PUR
FJdMbDf9SRDCAP4+bn8A52+Jze6n6n8KOJJeoqPjLhSiWfqpaJv0xXhXSkS/lYqN
X0hIIKFXT6g3uUUkH3coXGhkp9DjlwRpODHRa+ZRnJBOuNjuwlMpCR1WVZG8bQ1U
WHKhCM6pTlGmtklAV57gXjcFbn84ckdCsh550j5pmZGiL3CczQSnf5gSA4t2B9z1
GnwX+cDzCJp/N75uba1bRERmq/kAtQzZQa2a92spB0FSdHuyapdZim6LI4stDFJa
Th7BWuFPNIJD40gG1Ke00fxp+TdZZR7ryIHwBpnmvvi1Bu2CJAkxcR2v4if5kqln
7Ii5HdWOTE2Vts5Cn+vCvKLnj7LVyntN8vhl5imiTxQ5MYNXiX5HM/XWXRPq8kGf
0q2Ocm4UX0c8oE2qHRALXhLcj+G0Jt72dA4PYX/UYftPItptzkrqBRGPbrHbMkYG
gIFjI/JXAtBEsjza8VTCksRHpIp+NxXdMxsBzH9OsfCMQ70ZYxYw/hXN2g1+OX2F
k7eUWUuzvHy0/R8wu8DM75q/E2cwldfmzhBfBv6qwAIZIFVecX37Ode+R5Bk/apc
6/nAFnNrAe/a+5gbIkGR9a3edGnC37NL8c1e2r1cywPtWqom+kQinwZimGE9MGH1
cxmRTikWyVcoK5mmuGAxsa5ckwCMIH8D1yGijBC/BXZv8WcnmKnLUCPuHevet+oH
Fr3Jt43k+kkMYGhbiG5wbWRgT1egKAkAezKZLfZXwGZVIttOtQFjq7kR8UYd8h+M
5JbRauHOG8xLDCIHdLwIpvMjzI1XUec397t5vKpa2WdCH151H5lQE2WltiyuzNav
oTnPvAia/p44d3gQcCnxTlJYZacouKPnQhhNXJFVsid/171UH7rBvAp00Ql2NucI
RKHya7drkN5PPwlFqvgfQ5rPMzoqlPZoiBsvOeJ6Q8tEvOjOEiLVIgaCwGp+Glpd
2c2Z6yM8NdYkltb8su4eqk3hTxxsjDuhfCb6a7NGdWZy3yWV3CzR3ihLUvvTPRa1
cNDKxYVlTWHtMpltmldnB3EywgIc6YKtA5YqJNIKUm01k4Dq5I9Ia2fid64EmPjo
7I8V5/1gbCfufWEndcIJEo6JgCMdKqB3A+LZfRojVyp3VB/XdGwq9tVwZZ+pD/3+
QRAq2q54TyeR+qO5PJdkM5eKfsjzRYQNz3TJlLAyMXpWlq+f5kMfHHBweWghmu8v
2gOV4YAQpykUq9BGvjwE8GDjibDzcC+ZIrNkWAZYggHyWkfotICfo47pXIcyUO0S
Z9YjoZIMSQO1VtVT6Ldw3rR/AAcGhv/SGfwudSmrC1MuAH+ONURSaPhwNSpTVe/n
vmCR8dHwnXf8lYl7UHGx3Vvu0Ft1KZz4jmxbT7H92oo3MTGLGcVAd+93O0G3Ci7F
7ctOgU0d/phCRxe1PhYcvuyW8dgTikWbhZPYAP1Qkc8hhHbcdIGuPBAcMkR0UZeD
rb8+/AIECqRk52U/uW0+6bb4S0Sf83pkn1tEBj6BZsMatz6MWlkw3oOp4ss8pupt
h/zAM24EnnK321f7EPi/2QHGkdj+hByCRb3qeaLvxx2JKcXO9qQi8hrwxiorqK7S
a/8RSbkw46wfgW+61iomH5nz6B7VFT9lFvKckGuMT2I3HPfdPnMMqRsWG1TW1wlx
grOJRA8RTutkYvCYFRfbnSCZ1sxgOi2SNl7AqYSyNXlu7hsBsVymMYFjJn2JTa2w
e4zJ+cM+w0Bzusi6ROJcf23gFhPbvgA6z54G+cMrOIWcIW1A0SP10NBKcVoJDDSB
5IFZL39q8+aWepbJag9P7yZzjBPxW9Z602rpLp++Vr+VDawgzZlCARhdsZzwSyj7
0TyAIZc+3TyGQZhZ7iRbdJa73WT2OUXCgQtGkHZhuPKvhJcRSX5yTZy1N3R6rVpp
liD6S1ehbTrOp9JARhpYsQogbzW5QbWwrkuF9vi9OhPGGFWfGCPCtCZs+657C/X2
zDrUXa6vf2ZY1MUJvcBV12xI6IEv8VIIryo90XhIgyX6kOsadI5H9oXK+sz0uBPP
nUuYoqTG058xC3GB+3GSBtfESFEcjmUnILiDPC6r6W5cCoLr6aaid4Sb70qjqYHT
hiVieu5pMyxD7ON12y+M0poYdRHhc4opycy4Hct7xFzA/rNyPdIG0aylh+Agf/I3
phIT6ndXc4nfcdRuuoLPm/eXTbSI5iR14bLi7/SAtvkHf/W1FzR77T1p/yVe2fti
aT0iI/Zj67dnMwbvRa09n9VVsbXVYSCTKsXDX19TJJjwsHN5QbqaGldMxVN99emD
LfiqBRQ7zAkv+v0/jWtlQ4/WOiqntEYnLbTZRTA5q6VdzObJs7H8onCPPi55UuCQ
zlFH+l8FPYhSsZhuwkohe/47guzXTyQshOWL2l4ec19Ni/+sNA8UvXnicjG8ZfFj
jc7bsdvy9UUPbB6IRAldx3YBToAxx6ZKblJSxpep9UCUb6suSQTQJetYx+ibbB81
of/U49RCtC7Zm4JGx9lcb0ob7V/LeUCx4Av6IKELmplc7eO2z6TzVxrnMqteF/si
7nWe7RZrDBD+aImKYwTEUREJu4MwaWouRpx8MPup3hHDAw7SNm9hD9DHifp3QaLF
3zEjUNYDeJzGWPsJW8jYGdlS7wVQphl+4SaWlNbEv5w6JqVgP/mh+jj9X5CVbz76
J+HXPzteskTZmU5PL97s94anO4/3sObJSMh6PmW+ph/jYZG2b7E3sv9HLIVeZVvk
7YGE8t46xKWY+XzmlHkrwsJLBWs14QdHNtfJRB8ewluPFMf/a6OSpmT0fYa4xOlP
sDrJnS4l1WyBtjUgyK+9G5kQ9pN5ZrLJ1ZesdmOqa3BS3zlczAQ9uvALQ9oS1GDW
AGlnYyQRDsG6EcROfPjqtfKXzs9+Lu6x8CJ2GJSTNF5wZSDS2hVBDdvUtkqO5HxP
5bqLd5WTTWmzA1sDiHe2u/kDt0RHFOy1Bes41N2ADGN3ziIuPuRNejwPu+1jew9e
h4t1KnRaulDwysIuX72iqmTONgpyWzlavKNT5GZxC7f1oGqpnDGnkkGjx7pfanxN
r5/u/fCnCnjt2VU1RWG1stcymC4aJASqmGvuqR9UmIf0NyYYZb0zKDIrUOjO8CtV
l+GBNj8g5Ar1WwAoNW4CUp22wd2qrOlMwBIZMVFjS2O7e7NEu18XkTHNGiFMwlrO
QG3flE1FU6r27kAGXt+lR4bZxd4VL+HOkMXRfevj//13kT0HyqpxvSbLVw2yn7wn
TgiCIe3LuwGz89hn+kMOjnCYIgJ4B+01xAyZDRuwPRaktz/HLeZeXu9T6N5Febn1
TLOA2P3JJVEAJ4Hr2vVHOtqRJ0l2oerLXY/IKAk6xafn0QkP6b826qj4NGmHmQuw
gr6ooSu5gdaRJc3zwijCcfMEiaYal6ON1nuMVvv69tqEvkHt3fBoHda6bWh04I22
pqFWFThIK66dC9Fb/J2xjjoU+S9PzTYXXgak0ONt7Ge20o2G2sh+8eg1QRxbcRaM
/D5fZb5UyYvoIjccNDLgQ2wguKicYduSP0msh0PBt78ofEmX7nAHy6ryh8QvmFl5
vM02HmrgTgoofJgsxnGbq8j7zSyxMWgAjwQjn760J/qgcGbSASxnwkZADkLzLX4U
V+ds5fVl+TyElFZ2kMINiyRcL6qI82ipN3SvC7QvQCCcy5nRc7Xwx921l3kL3YRj
CEKYw/f1oMISgxkYTowvzVcWqeeSmHk7RmH6qVka2D7TbHUX4iRNNxvWdkYmNQ70
kPQn5IwnCsL3WeMuWzRa9fiDi3HIFpHawSJHgqn3dn0R8K1R5ZCvBDykKrabTUQR
ySTNQo8g5ckjy1H6ykchnmdQu1JNfOl7D8lIm6VViwefTg0rADgBTScRV9cdeklm
Hmp79vQWCwhFKB/8wFbv8ilz5Nbpv4iQ0LIWb5/5TFKRYNmxK95ihbKF6FSRDlG4
b/MSNjIHJFApjoyQRfpojBLp4Crexkrxf17yjbHaW+RJ2jtafRVOVNGp9UcsPCzS
f+TbNwhqebhjyiOiQ/l0s+J5qRhevMKExJ7Ja11lYOuYGaIcqpXNP+nUxHDiNAvZ
cJJkWzXbas01T8AvePVRazCU+SHfbkRZsMU/MjTneYQantesQ1gkH4U+ezCWK2QG
rm0Hxc8yyBISoIO9GIbBN3lZy3MqGNxoLrdKHin/vSxWfBe2YiTWFbt/uwZdFTOp
BKuGJr6RommYZDQO5TDyEhwm6XhpAZKICdCVVsDBbkJAzlLjrPEOgWdYMoDJOaL9
l1YihzXdi+1KXRbDfFrfufB42jQWcUhwlGiWf0A+nZSdFuUAJwNgaUxrsd+NHD+H
Dbab70cmw3c+gqqodSb/hKzlLdP6Kk83lPRf4hC1SLddaUUcEwj58TWcqwofKOR6
XvjGAve8rJEOJnnCDAOpF9bTClATWL+zz+SyfQ5TN2X2LRP6TYDKAQwYJDyHIhDz
c+EhzvPXG7KOIeMxMuYuJLQp6zbjL+aBbAjdGspMQnJKHC2dSqlFI0PAbraKlhQE
TrfV6PEOLgW+0Aee7ah1BROKGqSXafUcCihu3qjeE4uzmtOPyGQu3KDYl7D8D6Yy
qmvRdG0mpZpa3CNSqmlA+UuDfsrm0+5rVeCqQSpI8w6FbrbXMDQQpQWL1BWeRx2b
w65z4BHvPEox9gZOMXhvhlOUKnZMFqh0X4xL6FFBK/8SkyweCGzBfBOPSRZQvlNm
ze+2ji11GH8r1DyyEbNsa8Il26VYrHOobwP25slPy09bgl9CsSnxBse4iSUZBRp0
/F5TE9yA8zqlDtHHFgUZBTCX7Ec6pZlXxqjfeczTPZWQJGcodEHIzd7fj1EG0Idx
BzJKJ6J1XOz/MoORJ+SnsfbtQhI7FB6TIiwl8b0oJN1scraaHoFyaODj6Q3kZlY7
lVhn31ukQ+nK4yxaYBZt2ZOFJUKvhOgoWrljVCCDls+/kFm2H3AzlRfLCCY2hJy7
iht+p0rZ9FeYC2lC8sE+3xTmsYRo37IcebDTyJAU8J8QkwD0MkWtztLuiRhNplfy
BkJssxCPAG2oKgcqfrF93gOMvhFFfT0ZW2QCqMmTHUuMQk8Ot2kqKZCLYOIx7Pgm
eGkx7zN/X4DO6AuC6utM+TUCvK1aoP5zIJCWyNtXjndPPueHqaqx6me0XhwYSjcG
03PrzxoZW/COnpDqOgAz52YmqYKXiE/gFYjnyfkBUhilf1XkcuyLAubqjgTS4NuS
s3D+oOz7SQLrBnPDfUUgg27GZm2rNID7xjIUiiSZqpoA4sS9shNNPiVNXf8zIJFZ
QcZMPAu9LpnKybgAHW75vzrzUMW5oYeblfhPVfp04e6cdR2QMiXmosg1DvL/Wj9y
6l0vkXATaSls31CVZ+2Nd4ENBu4aUkF06LJgu2Aj18TYSY9d4mpRNUi1g9dYWm5S
sSV/pzbnNTe5OAUVKuAOcqERHwZSM5JRLVYgO8ph/0M9vmAtNOpH5KNuKd63R7Nt
z9S6fuBsKJMJL0k6thDUiyoGmNR066YSfE03z+grug6Im048NGOZgvHcuQHDvlSD
f90VrVq8GPdDCU/mXxRKrgaZkjJ2vwuHvcebqSCpNCfmsNSnT4OIMPRnP+CvUvHR
2DV2uVSlGDYx0lht7C/c2x/WPDcDVrTlWooBI2kYyz5Ne4MThzfl+gIRSMrjVvEK
BAl6Fv1u8wwNQw7VZof475Op6m12GFEKa5GO51K3Jn65rJqujFdkAFRoERGEdjIh
e/vu5mqiiY4t0G7t24gjhxAeRF4SD++y969nTu8I8Bk7ZRLBc2uIrBVcQM03CrwI
5OFEx7jATaAgnI/eXkWBN117qH2amlG4CiXO3bAZgQvjMUYZEYJzYkezKFDDhIgW
b+MdGOIyEeuGPrrlDQFQF32ErcRv7i9a9XygVtGmTXn1Rk7jHPlgd0+D2dGVyKo4

--pragma protect end_data_block
--pragma protect digest_block
1yAtBxCQn50dSiZQGW0Ve9U2Fi0=
--pragma protect end_digest_block
--pragma protect end_protected
