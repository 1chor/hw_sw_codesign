-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
JctXR8OLhcKxlEUt8HMYNJY7axKoIRdRb58GseFTShk0RSericoR/1iLbNTtitEp
unIj5B6HYzlliHdtcpqR3fcLaSVVha7KT2OS7DuTELqBldEsFfAdxN8CrwJbglwP
PjW8XJ8p0+hnEj/2K+O15NtOjIvS6M5MoL3metU7DGM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 29739)

`protect DATA_BLOCK
KiZn5Vmn8WRj77Q4YAzZs3cnTHRDTXD6llAbsqUvsgzNkcTRWLYQOdgCaKQM/Bkz
BH4BzH3CoZZc7ZlQoK32PCawZGdpfXDoWVs/0B3uOBDLEkbI5EH7mac+S3P1bTra
h6h0YDwbZZhXghNL9PZW76laGet58y/FrI9k+LXS2pas/WonyLxaznH6Yah/B214
tUVEYI2cZ0AOzuRcFKsky2PmcEuQ23lv1+YokIhi8+nL36395dsw2fKByamsteXx
1AfF0cGJW8Ze9jBdfHN1Sk4mAweK7Kwn6Ad/9b7E1zpX0LCM6lYC5KruOtlScFs7
dTv/CyEuJuUavWGOn0XsxrrZdR0/WQvaXzsMuZtJSQ5X1rvPLd44bj14RlWanOHs
QDSoiJinZ2jpOnHBcUM6QfLlrmY6R/mkX3Jnu0lBzwsvbm/cdVY4tmxU0xY6CPBf
85dmqKTNFdxOo0cCbJ3lnyJAnO4sxmmcjLhc4PAnBsLUCM3xcunAuKzQHD5X7sYX
gmMZRBVrhl0hYSfb7tHrokjiLCDJvV8MAnLqgoKsJqgI+yhYWHV+OuK7RQIzYUFi
aJZXLvit0xqN8q0P83A/WioN9TyFEcsNj6LCjNSKvrmlzh0MWIx01RScDgNNGpT/
VpxuvpOilmHW7+OipZ7cU4C+RLXvyVNtKCMCtSz5khOrshxhrlRO94FpWwnqGgOG
adf3g9zT7jqtF7aiLYEHwV+z07J1nU7I3EGOr+C+J4NDKuqNxvl5MRMn0oQrKd1O
NWYusSzkgpDwq6lqlbUKLL43MTnZLAvpI5vkKJB4YJiB/4GZOZSPk/UwJ83aW8gy
tpxY+ybvdLxljOahIUNGITLVn9EwCezFb53k9Hyt5Y8VmXogNHMWprouchPSmO8b
Wx3KvyLaZSWzboCKIPR7+jC3M7k38874o1KnJ0r51f9qqNkzUNQ8HfvrvPlCMaU9
UCh4PA6WhIjWYQ/7vgv6FAYftaO6Tz36C/9Xy8mBw96rztRfA/fKrCXMZtxVQjd5
jQ/9SGedINsS+sk5lu0WMICO4yObzDp+7xBuSXgD3pQ0scYTigOAW7gnuY3imaFz
HPxDQgp0WbmOEdxYYcxEZs9XKxxn1n3LwAcRiAON1h+j3ryD2dP78n3wprXcTRJ5
XRrCZnW/ViC7wgdN/otA7R5ud8a1p0WJs8ITAkMmCbOoYJQcA04CM0nAQvTzRlkY
3xp2WhuS9P3hKFfRARAyK79xw3a7YJQYLfQYo0pt2R7yqDTkrFaIJ46CKNf6Qs0j
vNRwPf2OwFIDUtPjhpnVCTbEiyRxRtGLgDkWH5SVYbrsVpKS9/rabqcYEJ+liZlX
oprn4pU1kR4SuiBWP4+6JDHYK1/1Hz8U+/86/XkPlaQqvB6+vVxyGC3ASlfbH9qx
lGcgoiKO8KE5BKHu2F1gb8RzhoMUXcIAxCAzpkopyscjDj/L5WnXyCJGCmd2m6YK
SAN+0EULxB5jS8soVVf9/2ZqF6V1af1tmPwJ+H4HEPc4jRS/hwSwHnwA9jQJ49uk
2RlKjw/dqLGNSfH6QlIB3KZ/0B4ywnwr1BmyLyeBNLloJioL5+4qQXw4hhQTUr5b
pBXgf8gCrvZNjK3QENcLeueYAZMPDMj1iObbvAiboNWLXtM+py0qvzZCTZQufkGV
u84tvfhMpra2lknW0kApPac3D7/WjT4zbXF4JvsCOdUef3LBsw+2bEqVqceBCb2m
71esQPuAKAxH159lmLiBUQa9GA08k1Rf/4h5wUfQeMwyZVNxs8OhNA5mxNs5HreU
NW9SlkFIXrJIAbAXKN02PnzJ3kpk2ieKyFK7JNgvsgGjrf/+ZB0FN0qvaHlywmi8
2LJNn62KHUOcmmY3QXxjfRSOTpB0xeVvsuB19ZqkdnY3zp/WmloDn4JXh/+TCxOx
jZliFfnTmUD+BrxotBbLcZK7YwZyuA0QC03F5h3CUov1y0x+ezKEOJfwoQ8ns717
oJEIb+3j+7MdFJaH+6wRvSHxsemGSjxTX1r5tRzpqpwIwsaIdq/eeiOyXa5FJKQr
ZELq5lqk8vIXTWjzy+tzosY1GTJ1i146p4oIC5mSte+VhOKZkFrvx/HIr4dENJJX
aBiNtQHSDlDoe0w46k8RZ27SiktC9QNc4Zlj/vXK3XzsPMihgqsrHQ38N4gZt+dK
D5jRnCnGqY5JCx7+emZ0ASsyI8OlpCCh2jlKJB60r08yU7/S9UeTm6QXkWreqVQT
5jqgMr8nGMMdN9D5YFJRcYCIAuIkk+9dOusVLpE8WLFQUXPbUZAxcGKjMrm1jHC2
VxebOZc8SD111Iv4Xh9qh/L4zy7qZttbdyNUfGIjp4CF20dU8Nv3qKMzxJ/znhyA
NW75ZdFvV2kRDmfYqrUjwxVlqyE+kYyfinBgDGdhSyE7VZXoD+yU+gIug4eUyhen
G4YxcQQrtliZVzk7bEhXekGwmMSjI7TJU8/CMDrfbH+hCgTtWABNpqa2sz9Kddx6
M0L1aL+tUMNqma73+0FKwYgx8Td6/nc/amPR/KAc71zxz4Lb/FveySQRb/e3/m/o
iP0t2Pi5w5+w5pb0QD7ePAZmkU6As1DEOC5DW9aIK57kJkZho3QwyBTLqWZI/0qc
I0e0Na2OYEtHhpsySDsxt1PVYcJaEsjTcYhno/3nuIimF1XW3VGNURMpPyMjDwON
YFpZSyEgCQyMGuKwxFFsyHSjwEwUE2a3b1JBvyoUAAEPXpog+cWiYs4deG7sCaKs
xxh8FxULNsMFr0BJ8gEgSxDQcuKC3bbUPArMZ01OZ3cZH3u8GIIxiBlnecVOibHN
+d+9eHorI+4+5VrHzhJTmxdJOokJmZ77v5SURI35D9OS5bRYmc96H/UnjZWBtbhu
8zyO2+6wfuzNw+qcewpCpQFuWWAgZoiNBJQTxXBPopfyW5ZT4ZxpTkeGgrvIt4fb
5jXt2zfcWDpH3/8u9GB73M7/KnCemri646lGYtnLG+F8KylIsdTw1KfkkERK1lb5
iMGqvN6rYJFEFFIuaakqr8AtD16aDDZr5P+fsBPnAIWhZl8KsO9BYFvgz4o0mku3
6bKitE3KAUbbmuFHwi8rDm9u0DS7A6H7NNN5Iie9Ak4zCHFvie+qgt9boVoSDhfj
9QBi6jvsWoeiFFYFydlKYUFbGsZvFUdfXOJR/toQwnjvyfRz+FfcrSbJLMRF27EQ
siFNGq8V8PQZvrryZ5ThCs+uwj9LZnR2Ul7EAYGAUuMqzIe1J5U6kSCPsBzVkcGi
FVjiFsIpJxX0L7rLqz6rHUKFo+1MLl3h/Cl1I7EGofPRN4WmCpE3sGRg2ThE9t/f
49gd2pZIP2zOpAnl9dNzdmAvau2dITcn+ARpHWWyR/W8afQKty+W/eYAkbPcckEO
9xwRjvvuyh9NivuBBjf1TaN2LQgZ1K4YvACPirnQGsh6H1zaCh36Ee2D8F4bOaZl
YhIGjTB2i7Mywrf37zO28ltV+vWhklxszuTd7165Cfs2CyedCcM3sZl3alNgxxCy
OG88HlP6GEbCt3MTt/tYzwbygaCv6AtEVbSsip4qBTQx/SGo0LgGXu9LHyYY2PA2
ufBfiiA1g2O6W22roZBW3RjEp63teZfWs1N2T99zvLS71Thmzq8AvGuI3AaRlT9M
RPl6HKSJ4Jl2q0zunz89PYF1n8tFVIANfsF64OU9f9wfrJ/GlrXRqfPqRXQt+9ac
nvoA2/OWInhdFI+ad/tRqidPk15It14CZfiltMS0x+XoeCRoS1wGau9h0G7ar2yA
KNexK7NFuWt0yhkJXej0d20sWkh7+zu0KxUVBqj+2zwcuGiSItWHwzc+TIIq2z4Z
I2v4udXT+er/nqtOKzk+wU/Hx6wYS0Kzyjp0yWko5fnMmgfpBz9zfWo/28pRZMKF
rl9zD02aGl3hb9Apqppfr3mIAvwIp9qTcj8ftKtzWeWATxS7b0/fBZ3NHF5bkgV1
dFFl+J+NBmx5cXgZC/9TSwi0dq9oHlUlElyvR+HX/fiTN4h14pIccm9VNeeTPRxo
PNHSQUjnAFIlSIrGKFso7vcpSFkoWtyBo/cqDnMhWOjnmiyAz+0wFjjVxewaJsh8
jgtAt6YX4QgH4aXyn6QH2jIbipqThE0LiRBe3Nvd5VaiWYlpBpxCchJ8dWNun14c
Wz+xI3vrKE47rYoZb73FFDHvb+1Av6SplixjqWZ7SALr3YUk/iUhPI4GJNLd3GNd
T76TT2S4OszH2giJ0/jKEr/ISuc98s3gDR6LS+02dPK5P1ploB0PtNkxhzDwyMzU
J/jyW9IptZ0o4J2l5GrLYf0dSt7gITDnJCam4hbqiXW7NK9MTTsWWKNznFzw6ema
U7P4oNvdfeXdhnqtKoTgXq7X/PaFzZnQPukG/hmP3P3yIm1dwHprHDFLKgZ5SCsy
WmlZFBvuxyBlgcPqTVZXGRmPcS8TmNzzz/WC4zXYlatULCcNMrxlwzvhwU0zvqzR
DbV1iqMtKHlywY+pgAzM9fMD94JyceP72TtQKDczHJIaxsq8qzqma9QfKwUgNcWg
q0YYUFqV64YCStOohkN/EnW0flD/KitM6FsIWiVAcveDCWT7ufAWpAKbjxnGbaPD
kkZIDuHE8+PfXihv+lyvjHKJDeJs1fZHuh4bH7AvXrQWhaOPT1e9H9s7Njzu9jBb
U3jlFyBXgkvc1HVJiKVD9GOacC5Ipo46/meDHlRm1Ww04/R8N6nsgtHmWgJxWc9i
C484oalww5k1LAR3M9y3q7JLrE6rukYgmr5KAiauCLKU3UNQ8bdD/qQmF7ZOj1Mq
nNkBobvpgI0lcklAzzYebtAhFt5W6Bl8zmnAoVPKXL8kOY8hVGgOcNrTukcz2Cw+
qJ76a2eM4gaHedo5L0dzQ3jBLGH7Y9z+Ag96d84bsqiJAlwkW9+OuznCZVFqtbQd
Qv9oSs5rbVRACvQbPnRIR7WYMAWqlap2krNR1beqr8EFBeO8C0Fq+IaK8jKMAx6q
8hij4VO47V7FLuyLDX2ToKPtRRJNa579raQMehSMElvUNYpx+LPMndZCNYm8zpl1
mGtu6TxtI3l53YZvNh+y9AoZiDtnjR5NJkZVgNpm/0QDYlC0ZWI0sT1M/Gcu2gN8
vbPR4+e38MyD5/GN5xyDRuS7TUivZKz2p+eSRxVNzMzyZm5L3v77qE5x8reDjERW
9hiYzI5jiWYOcOa9wT6wpA0yn+pI1UPJ6CfueHL997AVxInpKxOlFcoCZ1HVF7ng
D6flpsnwM+0OT9scRxEQORb9qbgR3ZbV3moYmPhavCTVZPu5yktrW9Xo6aYtr4qn
kOok/Xstja0DBxha2OaFnQXOYwAqsoh6eltVV8lTVOBLqiJavZNdEoqfhoULsLJl
SRzqHW5lQCaymWVnj+EbYefgYK9+MLGO5FyphWnf6xaae/AsVA4K1ymHYyrzQ9T5
2BBeHdOVv/y6404B6GTVikM/farBAyvWpsRskuPgP132T1VXVcI0Kg4qn+LeHvkJ
nknLCBtlwm+NdrQL7xpjkzq5UU4+jw7jjKg0bKedgxkInD91jXqJLMmcjc3rXLeq
i3ujdqCNQoxXE+ieavlVU5gDTV+XqyLDPkOwI1+IW0wAJSrr8mbL0j8xM31Sk8+N
bxQvFtX59vhymL1DncrKDEwh25FZ5qZ7vEs8SBHaTcj6V4I8/OgsycD5GLVdkcLs
vMgoe94o94Zng44R20hI6UF5NxXPKNlzX1c2lDJS2P3gZs6OMM3SkxSZtJhMtSeC
4PiNNVvYvyTCFlbFENfvY1RW4K6JD+Glh4z3qbZHmOIr0fUD4lBaY/QmeXYqPEMr
phphJT1DIP09kGNkH7AhYSGof17Hr8PwQSqrvtS8xyPVWi0fWmNtlvmZyk/W9ddP
Fxz+QAXVb2DN7Jh+xLcrHjbtyunVZhF3gmkozTdUBNngKlUKZNNXEYO4gHPHnUwj
hI+nOs6mG8Ixh5jXAJK+LqNQoaqoLyHHgLlm/S76tXQb6KiHTxHEuHNnMVivkPMT
pAi6xHFEBwtjp5/zZAE66KywBHzTvpmjrhOb6E39B2n2NT1+x4Gens45ZALdQJdj
NqUuL3w/Z/eqSvfqRv81FUUvLWRHUMNgpNGHCzBq00rWpkdgrB4UU/P10N02l8f8
5XIKTxETsRtKUlSAApOjQVGKhrHqonl4LPfj5Ke2H7N70zi1MJqxcU3SD3xQXOBY
pRseuKJfExz3qmmshKPLRiRef8lH9XU2bsPuwCKOSYaL63ulQjLPLNC0dQPQg3H/
zHj2iC6hsYIykyd7lexZrZknKjiEB+fKM8NrE6DzsJPiTKcJeK9PgNWJeaE38Qy7
duUeGbKG5eXO4oPge5qguvngO3a5FuNcfHQMZ5ZdN7T1jOiOln09Y6ZKvhFWLLjm
F6Xlyagvk9cTgz5UmOMNVVoHCId/h6PEmhJl2SDAHIw55PCyZ6ZoY/HryM1xK60b
QXvoEQoplJa1g2jy0E9PJw8nwsSphgk0Zhi+cg4YNypw+RL3xQOoQtSn6dVWgLKL
/HMe9BBk/PnrHist5V3wpwcpbSpDSSWoJ3Ue1mbrg3r5/dXXHwTk/H/n1NNjD0nW
18myP5mCXTpmW5egFBav0F76UXBbmTb+cNyKj16EIq0qvfdLaG6T3XBOjt70IEna
bMGWTO5S8FuoshECHJSUI0rR1KX1h6tfrEsQUeTY6j7U3plap5svxg49hluRiJoN
OU3kfEtl3+9oDOZ+NQsLiAdv51nW6P19sPxrWHqwGiX2XZjwUx7k+u0RnkgdiQmg
gyHWejsufRf4fsqzNzkav5XVm9F8DjTEJMy0m47vTFrhL8v1qSW0iI5gD0EUvVe5
PcboxuBKb1nfM6Lpe1/G61EWxKnayXQgSjebfyc00Z8XRTCr7w9rAJ42ZkSdu033
QXIFbq+MwKA5A4PkeFhG9/KBoFLNYcIQP7PNNV0W7Mldk/UtbmijDPVGp4kcj5w+
cEQmLdD9KDcTh8AYxPhYoXZzoqQ7Hv+Nejho/lCKFCKfDnzW1oyG/rNXHtvGF4dI
pd5jPnaHKRpGPJkrMyvetngggCIV3aNxaOZMLtnXGzS1AZDzs8ZJ6KIi3bUs74lF
TzeHv2/mGjP8niYrV6xJCWi4aPko8Bs+Zfjy9ZdQdvPiLtdisj58N8zHjVKAkQUu
bCgUno0o20LiOstZRE+xzy5bqegU/HUrCGAIpJtCTcVaMpKWZ1E2zd/cqIlr+IPA
iWx1LmfPEtznZSymr6BTiLGVMwf2jBTfcp66vo7Q40Go7G74/TPGD23TFhxIao+Q
5ktptTFxr0iJUr9gQoYlh611H7Syx1Ceslznk4PXhQlK7RMorGEy/nTf6uLJcy6I
uq0mhbyvj2Kz3XP7C8og+YY8BJEIVSIH+zrqC64nmH8mc/S7BW4djw1Hl7C/Fkxh
56r7fyaDYrPtAJirS1L1y8kvhLMQFx9yG8G2I4JvV+3lmXIf5liWBdLmVV3DXgzF
988ce6oD5OMLxVE6/cErkjWQasJLltfVUpYgi4613u+5bAa3ng+IYv1XY37amuMM
ILkWnIuJbARFyvsB7IKtKy56he8D9MbPkyFOa2Czt7Qaxj3xgRx0e8XtobRqNAWA
HNfggBZBuU3fh7j9u/ma8R+9q52PKL9wup5bRfJB+GhXajkeIYsIye9fEmw/CZVC
Fz6JLz3iajZGj9IEGK9hc59FbIff3SBnBlXG5a9eTHmxX+dWjDXOAu+gcvq5ncdk
LlqmAXhagpjyVuy7//EeYomoo+bsCxlGgRCD3h3udpCPbGmuSpdRED1OzUbhEYvo
QLjA0Xs4WpWptvtMO+DxKiJJw0ycZlsZywUHeeurhBAfkQMyayCsitNMuDcxhxa6
axOP3mRH9hMFzf5D79OLS3Gqf3I4gObbd6AeKD8pHDjDmM9Qf9eLV+4rQ+nIYOLR
bQTR6jhWG3I6MAhQ7T++tsU7o/UCNJ6S2ml9xpFzDrnqLRhFOs6g7yAW7a1rjOdp
6LR0UnKe2Dhn5BN9GJBgjcFt2AbMRt56na3A09PfGu8F+MmuTantndFKPvLPIXoi
SjZ64qipopPNTAf5Fdfod1XeNDX3RmkBZjjyvJUFk1adkbVUyXGfw51YaUwnRUXa
YQm6JjZy/2IDS4ZTWdF/hSs78q/2FZDN7MZrRU3J5TDBsHFdfyOmej8qfnY0Ryaf
w19shSsFaetkmIOC0TeRCydPEGKKKJSiP8BpHuhBLn0KaXyYjFPuWDveYoYKx9eg
yHwcteK8zEgcNvbFUwqDr6BXMGU+JrfpkPvScXRmD702o9A6GZgKPIUUGxtLJylg
9L4fdGLckggTvu1b/q3ljnLVfCY6hwnJZZdntVpYmktPNgMspFg09JAafsLI6qfQ
pxmqQin253McfzyNsXEWioPsXH7c6Hwn+3LGgQbbM+bzczxuyeaDDNAHeP9wnFI2
lIv+t48gdtLJX/gVfJAFwtcXmz4kk2oceNat5y4k9rUuOrWomlAI4tDVoatNi7hE
FcBmeoKFBbjeLwzruR0QaAfJgxXviJtvg3nJJpry4mcfRUtdFj0aYqlkjynFz6WH
1LuCeyZC1L4DCw2pJ4AyMciqnIRu3q6T/O997XIWDqu5CLC6NeueNW13nHoP7XoF
+1YWvrrWba0ub6q4MduyNSkMAUSnm7E4HN6pkJKrcbPKmYnL1lYS/lFYoPoG2tKD
wsqTWUz2I9YWYJOPA65klysEkmOkXMl1107f/m+2LhqMNXv4gNXzZpZcNN2N0E1g
HpchvBzqXqtPQufYQRTisKHvxq2PjC289xinY8yMdiZxmqUhAKcUnNvIpX98Pkpb
z1uhUVH1xcrGA8VqJMjNkxBiWUvyoj1q6FlX3H5fJAPCBgCv7WMahuwFYwkWqq4G
+MN8OTZ7fS1WpheAYI+DVdmHwQuSdNHK1+cjxYGBj/9gzoa2ZfDm1RzwKhRckhVz
EGXhddWjZS4hxq2ZFkLt1+7z+nvDv0tZ2XoTQk7/411XgC+oNARtkFBdPEKM6Tdh
rPD40q4376YY79quimrhT4JuOVaqqxsUZ8jOaswjBSg+81dHzPQbfe9qimtVdvXu
cNLCvN/85vJzKHuDU/Jk8bqnLOaRv7qh8mblQxfP+sGzmAbJqTD+PxCovI2s+Ji8
6SMPI2gLgLOYM99+iUxM91BknZG8JNO3YeKafLoa0ATwh8/1ncR2cPqmtl9mt04Q
dlKCKyFd7ro+PN4Z1FMeWjqcP+zrhziXlrjRFBrsvVtp9wzkPiHo3End9BsfGYIn
5iAs/syuKvYBwbYDQ0M0Iw3yBj5zrcg9dI3uA0opGmLqybDkwDtBSgyDEOlntruN
7Q+kpW7W6oU/7UDTlgEdzQ0sUhPHAWvRJ418Nl3YHRJQ+kwwAJvQaX0UCV1D3Wg4
T1/8fSE9lVV2Ok23pzMW0PXZpHCFer+QnE2ho0njjSkkczscN40Fkwd6hIxIZgmi
srXisSBR2irekYX26zCSpdwYWV6Aa35kU9rdeGlDfqlYVLEvgZHghRvXGGoHsLQ4
zD+wk779rI/qlEtspnieP2JgP+7l3V6JRTOvwy06TUCjVafV+JjjhaTgU7kvKWYx
Epz+vwAAZGOvQ6VTloiyuGOm43j5UDWJXcAGKF1lckot6UDqsQGIOjIQP64qOJN7
oQwoZIJock8D/heIMHg72/16wiM27e61AJxK8WfDA/gciUpGh8ZOxVRseH5Ehqyg
ifo8wu+atKCPqQkVGh32pbiCKwk7t3zFuoiqGXMuK25kKYLcWBOZ39Hy05Tm8BH9
wwUj11Zd/fojjMIIU9yRRoOOcB0xZEvy5vD88F2jOjvamb2fJ03cpRgh8c/zRldk
XR0UpBUFevcaBn4kmaljTLJLYnwAmWsvNFUNFRblbtkyUqE8IUuC2mMoQvxWmD8N
ZETVLNgUAB1NSJt91nr2ot0QZQrI42gyecxx6mY4WufkAwwPkORMePG8Sr1vyFaE
JLhWKg8hUyizC2xBbTvLhX99B62fedYE3f1xXl7mDRzaqNlgfdmomdzdyEjaF2Ao
yLN2JfpontsM5GraSRiDTOvmlap+kOK8yLvUSZ3ps3pNrFr42zK9uIYOwLVJGukl
q8i5X5W5JOKDnfMwu9QgKi/bh4BduHjlfrz9sSJCjYID8pkkAr6c6gVI7mvEaXDV
stLRUzTwD1H/lYWMB/9hJTV9vrCPz8vg2SvUB95L7BnsJMomoskv8UBBI7euzZ80
0ASjbghqzHwgteDaqKhxUqrB+wEraV/hB058qD89HyVYqgLENo7vPyDJzIxhfhlM
pPQ0rksXqSxaAIIC2Q4wjCyV+2Z9yTqijY9jWniidynvm9IKipsxivksunHBpJft
Ad9KK2+UuTh/s+2XBKcFqIjbnoBfFKofH8JyA6rwAJbl0hiI0Q/0elSihmIN+Pbp
NBxn0Uc47OPdpPSFZpjBkQbi0uNyk9QdBIWj8l0gy5YLHC1vnyzBHv1KhYjIUFGE
9r2x+HtGz3Uso4/UON+cDccbMQVbVGQNVfUSbosyHyN0ODLubC8jwfewLIQj3vES
CD55stcPD5kh2c8kJQFKQhrc7Ye1VL6T+QvO4+1Mv+SSnPdw+26YhdOMgVbAx2re
kE+LdAOy7pxwpSmZUkoFIOxiXzuDm41vPKCIkxFQy5y4zG87FXnXZT8aHQQVQ59g
lu9sDI0ctkYRfhozEB8B2M9udnKHi6kxiw8YBl3gyh2dMbnE/981uhPzWLd3/Bnx
OWtBPoxA7RfMDSZqRDAjlSGbNrROUdsevyYMHwkew5j4eL8X5emIB3tbwrF3nEmK
gVV5mnuWnN2tsXyhIKIgQAey4xjc1odIi2GiPFiSH/M4yMI6Q8pLA3c/mxk4XIdt
YuJAZWlWLzNUn3z0J6WtosDa17SkQt7QV8yzz1P1RF0mX1eX/ejVmG2PWeHfKjmJ
t2eX3PRbhT1wxkhYYXBuXqi0scQWQ++3/Ne/3z1pyKdx0kaOXF5LCsURz6kAEbwx
f+UapBu1m83SuAo24pFDy+Ysp45k6pDnvOCnYfnHgp+c7ycYbeoLGPx86VfqGiyO
1sUTzSAeN3FfIpUeG00U5qDjuWy4lSlMxdZxhmjQtXfB0wjz1gxvg5KgKscFQmtF
IaQ1kEFcmbiRIlb9uQQRY/h2MmgWk/6A5T8JeGusnqaXQsTcxpFqeEGeAcY21sT+
lDebvEgi192pB/GH+gsrdV1qOw3m1Bpt3K82Kbr456CavEY2Ileh+dSx89Liobur
czO456/YYhpXND25Z4x7b8XYV+HcMG9vy+JerNPD7iDz2jaMP5wOqr/uc9MIg/62
6VeTZuLsbUW8/wwfFh3zNy/me8orQ1A3+Tl5p2jGjsk+wj3TmRViwj+dV+gUg1ab
kZl3UHYuAEWjFCtERRfEOCzYToNg53HmI7vhxZ7WZD0daY/ZxHZp7Khn8PMAJiBy
jfncJEboa7wM9WHn6wujwKMVH7+NjxRJqzdn/Lask21F4B7FpRnPLMyPzWBoZMZ6
B8svk5MnEyrUrGtT6v9kV6dvJUW+bMl0U6u1otCmu63UwcA3NjHrOXtUmUa/j1ha
2WLygQuEhSzOk+lZ+e4Nbqvl58Rp1kI4X1474DEvjOSR7vRxe2LoPwG3URnIifqe
SflMhlUHof9Qe8bM7sS9qW1S1pHlkemWZ5M2rLMEBqkyPnwP/WDVPCJi0qtkOtsm
EIe8asjBh7ZIp6gIpyr04PzmKDdVjSdkPqqIo3nQlssHMzpWuHyOiE84uD0kMPNB
Bm4gTmYpjx/fQYHX25xiJcwQd9QPnl6HC6Ir7fsCYpbKBnJEM3xVCEDzDfUWVmaV
1LaB3Xj6oEW9gjms9B4qN0PrATpVbzUwxxTybYIMmYiRV1shRP07z+FXLQy15mBM
k4TgHOmM2rG2CR93Zx/e+VaxV2euRCIrPTNqg4ykoHEVFREpMu/CawBeaQfpT2em
NXls18kddvHYodWsirugSCxrn1amVty6Q+Qwmt2F9T3nub4PsNG1RtnLzXAYRD54
3pSbpZooMsnsBgSc5Y92hAkPwqUJ3Fh9VKtd+LJwELi/1ODB2MDf1afXtxo1SxZ+
aSAyvljEjW9zz84fRBqNs8hltdXMikqdAICfrRS15vC0uF11clnPv9Y2fsZcfFMk
3PdWVu+Cp/c3nv7PvnXiV2J/lPCipVJAUhRXg4WQCTsjE7vbIrdoaYy+1VHL/80s
X9jF0IRMpz8PeNfM2Las0018z7f0smS7YDPk31/TLvFIls28AqHmuO9ArEhfQ/7M
5QGnherSz2GyLkW85TApWEAvAR47OSIh/EG0jAEg48LG7+wQ9bdvFTqBlNTTKftH
vcYkvX+wbzYRYZghDluiGObn7CgjXFmgGoENQ+xx3lxhqJ/wPryTFFPD3jnWFPnF
ZJigizmKUQGggBwDpIn6EXYay1oBiNmdj3CT47LkO1yyh4F3gkbDSYZARWEoFXFP
ixQDM1XTuNOfHQFywzi8sde9dl53IwGmFABFQ8mDDa1PmlFI1TQMr8RA9qJFbq+3
eN3Y0gS7QII2WP8AQ7i3VrC6QHd7mk/zVZ29sq4n+eyEiYbiz4m1Y2T7jgG/Trfy
h23JH+Yzp8uy4aVEcjjJIQxo3JaQBbKnjXhRSMouKIbTxeIMA5Dl8uk749BFYBhB
Sy0Y22+qFrIz5WmhRRPgn7i7cpeknbh1eVQxqsKVwlxrkwBVeBF07QtXLkX/fc6V
UoQiZwfgX/aETMzBWqkU47GcEjNqfkOH4gFWijWrLh+DUl2saTukhQ9reI9hOj4A
HbcEDDcgB8yLBaGkuUyJFsHfQsXGAeQalwGUTZpTkbi7ZNvJH7C+Yyiv6GnGWpAU
ZmBt4j93B/w66FQ6W1oNMVaTbWOgls8iCvvbcN6TFKx5TEkZStvOJsXVExU0yYLP
wQJOUr4hkPNk94Qjm3j+SGG3/rAY9yeesPL0QO3pId5A/z7gbiSLlRBix5X3k0Yr
0UBxFfhfrjyLrDWEhmb+gHgcb9oNenaratpmvx08ESl0UZOZMERnlbJeTTyePWiP
SAhQhRbt4U99kMOuEutbcIiBB8R/3rSfldcv2M3wYs5gI7zSW7H37bblWYGNMeHD
QXnVLCsuQY/F5dxFvOU27wyYdRc5tYRQ6DAdVAaLtIAO8IJOrR3HrQuPpFhs5Wbo
RXYop4SRy9yTg7hczj6XBFA/1k6lF2UOJPfe5yN4ZlTzGbZLwW89hhaaPog76quK
SETYhdiLasnOw2d/h2aOJKkAD198zRZloQycKW+n1lNezv6oMBx0B251+8+R+ab1
CE4tWHU1VnZNcudmCNmOHMHrCTEIqba901S5ITe/QdDx/4Ef7IopyPEvcOZU2EV7
zEV7dytcUknQgPMN0cdDl3l4yM1952s1YcYX6cuLZ1xwGUt5ups4BZCGmOF0Hxqt
SdpoGkuK6ZJob6cOYqTwstV5O/KZnkPvrpE8L7LMHNgchmhYFdQjzDG9CsxiLzxP
oSCuIrJZoA+IZ76xFY87DGeQr/vhyri4d/MysZJOukDsJPU0Fs5ulih2BewLos4w
dGP45EUI63bzwMv813DXTzH14Jevd7ZC/rCH/VweeMlTN5i+M27c7KAbs/JH/oeE
px5Qvlj4YbFK97Oh8uJGVnn4tuAxLoBn0zn1F40dvs700fle2AACG3nx6cHycEOv
+4vv1gIUAnFeHxkNPFe1WqIHkkmcTOh3CThpO/EfNj0ew+tQx55o/bCO7xoeiCAO
jEuq3KYSwY2ktNH9BL5Dpu6sWBJc06W151RaE4RHIOqXNGc1ZV3wMO13Ne1nYOh3
nMRuLfpTvv35WZ6x0g2Q/w5wy//D3qp3FH1wOw+wVto0m4j0NhdAe/aiXEYWhgD+
PqATeGpjf6ukZIO35/IWEusiA3QF4KfDJ8u7VkO4lTYr+RUI1vfAt4ZoVbpMQmYc
jrrPsWpTwpZtI0MaBNgCsCD2DJ0XU6d21ojAuLkd3wblJyurxvFDmJmIGzgkCsJo
HZc9nWxuUSrLqCL+A178LuiDQDJf3p+yyzuLSUP4jUQVLDNfouahYxYAq3hupORX
RvmF8ESHpIlA3GejSUKPX9TE6wzN4JGjDJg6P91D31g5ZgssR2TwKrIMPVEC1uB6
sbGnwYBiaEQNmyhEmC2LvJMsLaZaxaMLIYr6Z03VzsEK3gmEd+F+POOS4qC8wfEU
hvsAslYlZukL33aUpXFVJ9cI1xd6VOrIy6/5RAtYY/tJ5cDBc3ksWv7sMqG/8keX
mcXnw4KYSmDsy0YgVTozkJyimD5k/89raU8Zq0tX598jhog0EgMH2Jh4T708bDqk
BWhfvsb86TPeDgDPsD0DJQk6n+iGjTn3akf07lGBfxjzwcJ1heWZZbD6EJ6iehEL
01hAXYoTWaQyf+By0ERpLLNfna/BJ111fXABOzBlSvEGnW1XltIo2kOXl5gvdCqY
XVk+2UXFoUbnRK5GTebYBBnhKirOJzIJNJFvY0L/AXp5N5zm+SJalDIoW2iM4CQP
hTP2ZseKT5TC0uK2XoH8fs2O79gEH9FyLHO/xRBiwwXz62hBROI8DFlXkcFV2KdF
GLKsjBOIV23/LbRfDSaUUCjV1XigrFpYOvkXHHaT70PD1SkwxcKQhKxDYo3JfIRP
KZf6+4nm3lLNmF5taYDOQD4Fs3x2usYbNucZmICxrTsFjUpU34bLse+GGn9Dol7e
VNZpy64nb0Nwko5u73VZ91xFV40ANw6cOTZ9+ZBZyVYjtXTdPCvApDwvjPnAILG8
tJsalwxs7nyj27E1euibBu9sUs/0aRJZVRlc5jEaPEniii8IntI5iIExbvxycxTy
/1Z5YW+lAlVWEvlPnOFPHAW9FyECBboFOJ5+uKqlUJNykZrjdcl1hLquVIx41nPu
3neKl+kw1ckm3w/0QTymSt1P0+rK7PoDj5XFnDM9KhNKm5VSoT9wlG0jihtHzUR9
sNbP+x1wD36mjg9I7MSk/k7kBiVZPtVIWfNmPp4RiVpZGh2G8dRLO/cfiaeHLxl2
nohGDUeDf0Fiqrskvvw0c/wbac3tp249Y7PxPH3bdZ84ymNKPrC1g8pbNNCnJheb
5gnD2Y+E+96ouWLf+nRr9L30bQqH1vnR9NE4SGL0dpgq4Gzhpd4asOk367wJPTdU
DyyAZGxRnxgYkjQyHWOV2JR6S0E0rTgxZD6/gEn8zyen5m16M9xhYEM+k4KTFn9t
QqpDY+sR150G3BDGppXqQ0NdhwhtgKf9te0W7oU3mDJNYlFZrR9X6IHH9QgYKSBB
1xXwMVIQZNjAixOcRg2qCxuSviobp5XBE/1eNoSIY0E5fG23UfBhWOt39BrTvMoJ
aENJzT059QLA3eIM/Q2/2cWDq8Y1rPiq5v3vqkRwPd8N50l91LaCpRPLlY3IrKMR
ClSm5RDSf/N/9kAOusLJ6LX5HvgkcWKk6aCg7mvfNrl6oQhXwCcFsq+nUGu0MdST
U4cmusqwZeEvrXeglBWaPZ6j/c2H5kWtDR3WNxULLku6mES39K33n+u+D7ljmVRx
K4fF5VfzIi/8YD/FHcdxHcMmVQEEeqQRksSmUloruu6fwUWD3LjvP15UEIIkxOu8
16z2Fa4/5AeIRCbDwRn6VdUrfzpeBun5cSGdC+dF/H7oRLu4V0hq4nhMeatLlqdT
7KrNnSsfdNs/GK3QXnjH9CDLT63XlV57TA6XWDp3mOpHSaZJ79RgFdg9MEP+UTvG
vgR62XH1oPC9G9ia+XTeRLrV4T62DsmPK9fjato0NUv5VoNANLydOjr06bVBkszx
6RP8+INCtX4jI1UCur1WNwfEBG8l9VAqlDjCOQ0TuD80aLQb18llIRiJcJ351dUK
zs3X6HXPXh+SpGRH9LRmFbkP1l0R+beLS8W0ubsCpM/uwu5ULw2e4s4YnOXJT5rU
C7bRFWkeySH5hDflSfGKPW0KKhFmCnL0BhMTfwzu/ktwyV/6fIdnvi+LvdH9m6f6
faqCyeCSRNbJGJBkJt8ccf8xuA8AdRE5vjfjA+p9+Cf9OcwO2QePb1sqjZ4YpOKz
5cMMjG4ckD9F00VWvh9yqtYHERZz5LBDGycaFDJiZiiVHObLhGsSBwvn9G8U7MXn
pv+qbmxi6Yn5C/3LnmW9CULUQbsr899wHP2oa+zvCRHA9vhjzra9gTJh+7qfW9ZP
ofsgShco/Wlki4fvDBY1/Iw4WVfFiM3CDwBXzF3Z7a/9yb5a/ZHe8in56mpKjZW+
PB/F6tQyxwE2T/p6VVp+Hva1Wg0z71H4HvOpNdUBABv1aLqNQAtyFq/q/ve9yUvU
Uf5AXwSzAS7t+3QwAYYxk1a7jMlb/5+eJ1sMErillfGlx0w/V1L/G0dx+4e1Ycan
/Oxnv0Xs3z77w2uQyCtJmaqFCH5xdNVWcDhMcF4wgGuzqf3nMz7v7i/v1+Tvp/eT
P5Ois46ch7bFGdWFrhhcXa0hiLGQmDNi2L1RbLf5lGke1oLy68Pwh6DeDWUozLI7
e0jAsmSdDpur3LQL2va4XSiHL309qDi9ViyU7S1tHQef/+63AkP7dgV0C6ptgvMZ
QdetqOpRimWZ6SP5AgLvRMZS6pSM7JtvnsO7nQU1Ar5oopE1NKYF3vbqIXvILYR9
Yly4Y2FJGQjSfeBGk5k4Yk8VmckXcs64k5dzIPJUbiRUYj8rnVSmXHafjYxYszvA
9KJMMzWemFEYBmhNG7abgHC6lcnoSP37XUaWnUKjwsMtrTztoc1e3PxjmxxS5FiV
t5gznR4w1rNF7GTL+I4lh6dJ5a2u8M+QUseD6uIluAiyzCTq3B/nY466WKGpJ1hy
FWnWvpgpzxWDsB03jSOWf662fajRdQrfSECdL5QjM8AVxhADIIzM93/SDVAGjixP
G6l4WU0c8O3GVx909bfEbJVqyBI9PJGVv0EVqJsw2YOv1jzq6yEy9dqXkoFRCX5Q
MEfMXVGK+5TUO3KHuIkvd9nwpUl5FErRKvkaUNR8taBsh5TvwrbCVO5jamGSECqY
ykE8HueOIBw1AUjlhqY1X6PewS0XhMsvSz/P4BJf9eJkL27czcyMWdEGhVz5POmt
CBJQWOg7BwmUYFntKFdr+Q9+Is6HotIy1BUW8ce3AP/GxhRkQKqxi8Lx+gIbDScW
qj1aNRjaT8m6ChblaJIynupLEKC9ba+emWLrW2Ktii3pMZHE+oqTDZeLFSIuUxuy
u2bsUDTrzUyaVTNQ3v9oRWxERfUMQ4vu3ikiG8WeghfTwYbQMv6xMAY7z6D09V3u
XEo86WSQNlxtlk0EGnvs3LPE7/EZV0uxYC83MztGQ91T73JhaoUsLrIBaxMD4soN
4xJL5tDhtDDK07ucszj2tfJgEhLTXDJOAvTpmB3rODTmvriJdux7Z89I53q8uJ0C
7GiiAX8iE3iOKq8ECZDv8CPtxBqAnhnkLSFV78i/CksWOkjCuXiwk9/jldixtRM0
3ec09jkSTpQ4kQj1boTrE9SxGG7k495y0rRpExdTQks7wd8tkzX2ah0pbMsiz6Yw
f4WP2YNZC1VYHURVAQTcO9aaoWjrl8UPEcv2lIN3RyBc71ULXWVjlibIUoS1sB/6
TnoLnstIEdjtdt8XZH4L3Jv9srmSm+Sp382QUl9VaVbUN8D1NzJSXXU1sjdLBI9s
y+OllXLusb6G+Fth7xrF2QwL8Tp5YuI/2uMC3FBYZRJBLpJYuiiIXIomh7LAbZYK
HM6uPDUNrGw+4CymRSjm+edDCQqxvslSafYFpgjA5kR6mT71fj3nt/9Pontqvwb5
kxU/JEyGNPs6UfxzsTFloJ5fgnvKaRaaGcm1yhxFsZo3gLub55jToiLSSEwGfDvp
+6p9n7zuV+nepj68QEywUxf3wO/7YYPoKX9AB2U7hoeaPXI+WLHx9CdUVoEoe+BT
LEH6tMueg7m+1pWehUy3lvIXVZZI//Hq3VCLUJNM9eSRVD8GKgplg+f5LS4qSvhf
yfBVu71nQv88pxvwG8HnOsWkCj9BN1mWwP1aHAyKX0zqNWFe9tHYIJxmHpepEm5O
dNIDi3GWORm6TdJP4dVHtLr5t/3UbBu/bNjo8lO6/0/Q8BIIWDDii6Pzb9aj9UVD
xEYU0S9hSRMZBy+ihkAJOCTcnaJa/QpTsM11wiUuUs7Kwhyn/zs3Eq3s+K6VtFME
ylBFOg1bEy8Jzz3AEVg0e1+DwKXvJOq+Zobk89AbBZ5X1awMz63KuV2kOgKanM35
dDxdzbGgkEe1ncxgJ7Hy2x3hfYQ4pCNBN4SeJFNM4c+SuzmF3erjE6OFssJZATG5
URbc1rEEIJv4UQXHAT/roWEWIMRa1izky4UlKtVam/OEKCETxQy+5fQmNtWi/u0y
y+h7ZKDa5f/DvH3ibWMVvqX4qJNJj0kzEah9RW/lYx+q9xsIJH6vCQjUA/jfP3AX
ELO3CFpPQFd5MD0WrZbcPe9COdDUPlzJJOmXR8/SDler2djbuZNjWxiEci1bLgFl
syWwk8olvrE8iKprLCrJeKxMePfHHvDH28/nhieNvGSgvLwNwIxsXLOTfZYL34Ie
v2+TpY7BcfhCxkD316VvJ7WVuinW+t7x7AiJUcldUprpaQFod4X6RWHLEuj51MSM
50vHWru/rgWfJ7E4lk2jzZH7+FFVZryqE++4G9cBwBN5DYvf4TH/9eGat6RulATS
xl0fsiJ6XBwUMkPldCjUfd40ZUueTOcV+tovA3idbtvsBRtlddLBHl7B5fveRTVI
owFg1Iv4pWVzEkTa9zfOOqlSgFXjomSHiN9lL3YwDjIvQ0rTPOetVSeQZLjTVwrG
wTm0h4MfcA7JMdT40kfsfp10bMyTeQWZ3+x21eYXz2UgKBwDc1+BDnkeHia0fJq6
WMlXaeXI7MMWmGyB69OTz+s4ZyOib9M+EP/icOuO0uGUMFAIH4utCQ+9gxPYTHF2
J/4OOBu55WB7NtVSZta9tbcsk7/7Vffzp36bWCiWiQnQqu/XQFtdwhnWNZi1CIYV
k88bE/r1kr8fd7MMNTgR3qan+yRnPsJYCmsZkR/KsIr5ze5GlexVf86leLNv3MvF
QMgplBBg7XI8rzmLJNa3EatPmaEdCMfLQkSokqIhp6E99sDEk+dPaH8zhCjST7vw
kPEDGOBucYV3aM7vAX/nvZ2nVsnSmj1wvVgjPv3wnkn9ZQ4v8LPPWiIwM5VsgU4K
5vy/nGAxfowTJJRmxJj2jMKNVJ5o29ojpwP0AahipLGmiW9wjFWjDkQTiskHYD+e
j8zlcAfkmLKSIHTH5hF3brgKmtZZgfjtx+dvVpf1feo0qQmLnUUds8z0iSv/F0dV
k9hjbV0cVSeAIMOorsRHEgTFB8W0SkU5Nbxr6k5pNxJObnunqgD9IuKO+NaP5QvW
1ie20Uo0gKjJbPzYK5IEcTUNsgq+ThzWiY71p798AYLcN7tO1NS8XDamewaqkfcJ
LkHDXlraG01Lg3SaA37gaXJ/ABaX7WKHgQW3fM6nz/2rf2IS17n/6vniKiB1OyCA
eZ4B0Z+0zf5PE6ItutXOIJSfJugDp7Y5Ivw8NigxjrKDCssEH+vVVDbO4p8bTFuB
Vetz2THlJ4W9GO5hUCznE0jXUnhPyW7e6+RaD2xrPJiBCyfqW+cks/xmlFHofcC7
8lDaHL4Y00ANTWInciEvsyq1rEdAnEptNIUA9oGmSuQ7JbLgOl/BC5bZkYV+JRkB
rDFmhM5kyc9A7SRGkgOOYckDIEh+5rizsk//DZ0w9hSj6gAESUnVAWYhzI1cxwxR
rpCcZs2d+g70ZxcAdEYqEmc8UkhNEJpFicgMM47ANBdMbQKeDoFy/A/vHU7dRDrw
TP44K/+aWatX4FdMvw6/eWj53cCBiJTAonQ+sb34s9p5nNHFgzcsk/NeJUDCkF56
8u2WCNzQCPTpOza/be7+Ng8aG7pUQ3qq/X0mFg23uVnyb56VZdpneRWmBXNXu37w
T+q5Zo7+T5XopO0yIRoiz+AP+wq4UKDY598BxDP8PweQM8eZTJt3pua0EJFz3Hlj
UdAKEtIluuHpQmoAnPWxyOGwREYDeIw8jkKRBfor00ObCEfxi5tTBzLCXDAPSo6z
Cv5aAhtdz6Ikd5+8Z+DqpT1GJ3gSQn6rseZv8Gx3Tl++kSll8KozhGVGhYR+fyHb
pQaycE7g4uQTt6op/oK4kUm6q/Zsoi74+y/G2s1v6XWIt5/d9RxeH3OvKATHIodv
DgvnQaVvEEzwGE6jkHDRjemVhsJwJoMKnqUcF4cJHyFChqhQmFoKIPDHyIAicnve
8w8i1i60nuONfxplFBVpEzeySme3Voei12uTkMwn/K+GfCjf4FGWrevFWRL+WLo7
IOwPG8cn3z7/BIG1iS8e3/3nvU2D4BBmxZudXDyKmO/hX7mh9SN6rK9ug70sGCXz
RD5xLcFjjr6fFJP6Pq4tX91Ytbn25owqfw9gyJSd349mxzCkctXMt/YvHcxk8tFC
7Cr2VSovYNMRN24NZZlDX8dBxPLQi4AoOzphbANAtZiuvnoPM64tchtlQLCCFt49
SO8JoKfpzwB9YjY8yHIi9dNtthY+8En6Y3I6WojeRC/HiC5QyUgVQ597PlMzoVA+
+GkE+wv+SdKQdOhOqwS2wegCjb8pOyz+lK+TeQSJMmfJTUQSK56j7vqbsX9t5cIs
OeltEy7PMLAjdCD2DaxAo7Hk3q4onn2LMnlVeGyBMpc+6Rw0FKFv1qb68nyKxxb9
a/NRvi3qhWhVOZbvBylIhchTimaKTxAHwMaJ4zBpa6BhjaIKCOlPWf2OLyFSe0nO
TOma336YeD47UAb2thpTWOwwry+zMKtx1A8f5A51O3C6Yj6ZfqB61UulqcjbSgDg
R8hYRA3sFKhnAGmhSF26+SDeTACs0SG46Cm6/e8xjgQAlO8KpmMjtdpjD1tbjpKT
JRTh+D02cpWrPFunyU8r7sO4doHGsn9B3N4sbcos61l321AxbcaG13JqwIApqlCP
RpZAHXErW52QgTNLcsN32Aw84ZxeolmqlPEgdWypt2iHJn8piLG+Wp7BWRnUskgn
Ikh0AuGso1+PUC++3mgAHuNXQiWOar+QO4or2NvnW1/9M7jiV1EJtMHSZnCL0ept
sNLWeLxyLWhcBdKAAmP+cT/1Ke84KcZ4eIR96/k8X4m7S2KNlsEOC1yAFFTe4A2V
1SBKGKxENmNU9R+cpFXeJuf+zwXaT6TrjiBM2LmIys7Q9wC1EyqzpZwgx+TYF1yk
0AiaKUGf9PMU4csSbExmvx4tM27Stsp4tcMl4wy815T7cWVNculY2U9QMPtXeLQs
cqB3yn7zsnzTvzlKJJYoo8QK1ejWMfrMFe29xq9sWkrAu1G0bc3jiPievLRl7bk5
1ypY2dD1GTg7RvSGOhTBEyXYvNK4ov/8EaHeEMUNEqO0/CeMNSYqQs74j5uopfs6
Zkx09iTxoIWaZvIGtoY86AlPpJhFgKaJybw/N9FbFFym/EGkHgGgkxdT1bqd8WCi
VfMtO7VdFi7H/zm9OD+qExem2AyM51+5LhT1MqNB6wPwElLTfKPiJPB6JiNrQw7A
6JhEvssytDQlqGs1fKhIfV0gHhXDJwRAixJD53yS0x5NCUJCOTCCNUnb5odKHn/k
nordybW/mzlLK2xy61jvAOOwvePwId7ijjzRmrFeZ5SYt9QZyVrkh/wP4xDIPX+U
IexFRS+wflVav1mzPymkwFf0+a7NRIO/AGzrsSlECaa4hqHhFUGyiOEuz8Ueel5P
QcIYjZRa2hTg5gojv32tk4ly7qso4CUXRyQXsvS4i87axyZVYcvQcVVD2I/g3sky
RyoVVw1bwjrtM6Yyx1F6gHWlmQ9GeYZO3T8ghsjwFQ+f43FcB6W+gXuKmvzr3SvU
PANSjLr6tOcqWhLR6mXZPY0kxMGAIASueRryqsPczp/ukDQjRmFuV9ExRkW6Hkh5
AES969dwQXNv5bCepxgjBaqYzJikMkWPy2GAcXW5926Yfdo/UvIQLwbIhzMpHwCY
YydDFHuhoztpwHt7yGT5nq+iVeqUKRpZPV9XwcEn+zkn2Uwbv9ex0YpmbHvV+mDX
HoskxNPXr6f7PfBz5N+BUuZkHLM/HwFaN3n1wVeNmMiVRXZeyRsWND2XwqysvKp6
1jQP5zD2nKjQaIVPqmA9OiPCNbGjvkuxv4WRwdKefgaHM7KWxh2ClO9zFkASCf6y
VIhe56PrNiQCjouwJw0Yhwue7/hJrwoLnL3c1KzVO4izbUlTjSAGhtf/to9297et
XAkQ/jx21mm92J+XEYGxU7d+enceEqGe5HFgV1yvk5lb/lvLLEZAdCZZ30WLuM91
DXFG4igSe7C3PpDc+oFAmVWaGny5sv4UiJlFZ0muKuDO7NQvXnBN37PSYABbRkZU
XFXQ5MZawqVylxd11HcFdiLh3KqENeF7jCR+iJsNmNU/NdMy1jZ/2bLY9yu1hafr
bf0TaRCVD1bTG7mAjtrSH51ZfEyudgkFO48mFn81wbgAhkJ9BeMEx14hytklFANg
SdWJghsPq0s3MAC8naVDroTlnXxICLsH+39oA/ypAd3lZF5THZpmJU2bIv75TwEk
tlYPQGleDFfwWZmHREc0VwdHiuSw3FMbR7sd/2wnveRcxeEdTBgKhYUogThc935K
1JgUgPtd9cZTcJffO2VIaBBMrVTbiDeigdQMgzKJRtibf+1sXRUZ6TqD0Pok/HgY
0piddIO2pzlNKW5qOn40Rky5hMQ2p0nYvZlUvhNGu0uftY5xhYJQFGNQdHEQCKKS
QzL4jyISNHBhdRoZroJYFak1FyxXdvF96u0odJJiQfhKWXjDLQnEuAECPmuvyOXr
G/IK7Ywcm1SxmdDNsCjCkWHlmEsNxtn1sZNtRZVQrQX2lCDAFxkHczkM7wpVYn1f
SxbScT21gS7rfHnMOzIVC0+MNjC7nZe+TCyDZH7ybzYfeQzioYKGAlJJaAktcWkU
SX+ysrH0GbDbUKyDob9PR7XOL9c0vb/T/WEP5kICR4OatEILshNqXlZYzHRJVeKs
1FmoLU8IzMSbEArVoprZinGdl7d9UO0EkJ55IzsWIoW0DTfo5e8JGCvMJAVIl2qf
i11jHTWdktR/hFP5DYdfokWaUDB2MQHTbVKEfFTgnQUeCM+MsCL64r/mWxu6/uir
EkxIpKd/YDErn5KknjRKoJJr450gkn940NjqZXYdzxVPCsCjoBTOm3TeqVKO3fjR
2OBRufh0PUuS8AHBjuDUfku/xkZJVTzh3BpCmj6R7uU2Kf7dn69lHNN52+DGDj3O
Sl/E0/Ae1HFZ1KmaVmxbQcRNQGgyPpbp5PFXBb2oCBKuRbYfFDvNTSwxIElhKmZI
dDzxCuz4YeXpvfJ1dsuVZZECdccMvdBnuTZXBJqtKDxsMnZEQy4Bn3t2JTuv4Ej3
CeEkZufJ1ylVfvJS9NnZ+dn42dLXEBkdwT8mJuzN69Jz9mc1YfwYYt6f+2y9lSK9
xUlLRz0X9z56/5YU49Wj+v/YEX3WqGTOdJ5jgwzioqWFUlyDsjraQv2GuNIlnFka
1+5MOpW1HYvfNtl7UyeSaAjQglUsZE1wKMyGlPrfjMb1Vv6f/pNJ/zJr8sWb4TKM
n9Xe0Mu9psBqaqFpXtA7e+/qqS0E8UPl6pplaoaVau7Rcc0x2i+uE2J80hitBH2X
D2tuJM4cJC/s6wjPfrha7V5H6DNy7abdURI1eCsqq7MIflZWFGwruSff6+DqR2M6
2Vm7rePg2uDoKbkUjLrtjHZkueL6HtZ1gb6xb7im46rtLnMH9QWiVL7IrX4QQGSB
jP608r9du92ePLsQhs5WWLDLYngSmbWugjEFJ0zAvhHmV6u6TkMucJETOURMR23V
C0XVnm57ntqm04EhT9kHtPoGHaUn7YTxkQ+sRYGHBRvZHCV1Mq6PR1wwNGZEqEhP
QX7f6KHu7AWHEuJJewFD7Lq+EkUIgpQNsorA0s0h1ES0VTkL81vBJr92I5HpEh8R
0U7IaMFyi6WHd4MTe5W+jL3dHVNLpXAEEDn7rjCEU6dDNOlmp0YzcoZU2rO9XhCA
Hcx5WftU6vwTdySfiwYI4+knY5XSpvQjMbediPdkl3tca4hLt5PnukXgr2nk9HvE
PmmEeb3BFJ1UHppitWotxjwhexIR7y8G8v1dPxfem62fZGl8L6fgFp3cZfH1A9Zb
LrH7ciqTIzEUn9nKBOcyNeytckVDAN/u9hItizbXpR5bFjvVKEFnt7xGEtWSCkfn
9Z9Vpx6O+FbTbpjtiiHSsUM18okdY+yRhzPAeBWfaoI11uj6MWIfLpcNWQ0F4Yv1
6W9gQxpbFmfC9LzuIeO60RYgbUEC/FNqT9laUh/x+iYeXKCH3s0nmPFjyVc1oP4C
3K/mY/t5tTbftnhzR0UEs+CUwT1K8ZB+LUxjWn6TnkAye5mLsvctPmtoXVKJDlF0
mgEgtExuJYAljquJKbdqy8UYB71KVzIhCgiOj5EtJq0lOyhhT+CjYYB4nC/fEff2
W2ElFnIgqwA+fUNvH/0WdsKAaLS1eMahp8eo7r0WvqsoisuBFuRV12BhW3l6ZZ9B
KVYdkxGvxsAGEVLgmrd1BOaFwi0iNJqpZAJn1G6bWZJcEW9aCyZm2nJmtIBzkzyj
k5aZm1iigfYwZbh68xM+YEVsF0TEHzq5XyPW9WIjOSpgKUjopNW6dNGFR4uraQKj
uGZmJo+0Iszg50+qgTmcc2bWae5aiGC70V0HYdVCUrxZbAmZdQOX/fcJ/TJgeUAb
n9JU5iql+dPL5uHiTkL9KInZ/pH60tgUSarU5JgRQipp6pbzE/yN5QsOOwKJHZgP
trj4vydvqB0WzVDjs3CtuiLibVaP/+B1GS6YssgrdJQjVEMd+Q1WNCUSS4TjAwSi
W70zXTkwxqpUG9yXeI0ct5MazDmZWVWcSlI03fbzf6Wt8O1Kn0Ti70wjuZHumzc6
7Ss4MJ5IjSahAXxxNtWkZB9Z1mdodSmmEYi63v24bexzhSC2Z1lixrTbeR+bldGe
q7iuEIrA8LSoXUJZLJtfnyx8uVgcS4KOC5QnHxBJ6osHJqdcIPaCod9H+GrRuLYA
qWIWXVNuMEP5j7RREeJ41CR0H9Et+7EXWeqqkfeQOQPNIbJ22/zLdFEoRi0mxOE/
qMIHfF5wYRrj4sOq2QoL5cpIZX0YQ4XgVqURGqpP9441LbjRtq1eYTMN5yg+cMc8
xe0cFMEpWBLR323CjdqoltniNim4BlUULtBgU5dsZ3XiQ1aQhfwr95eYLiwlAL/w
3w691qD4CrLATZtvM/4dUs7Nb8b7Y4iyqClKMfM4GGToNZl3E4v7HJ1pocrZpGu1
dM3X3IEd4qACZD4A069iAVuJb/ANQZCeD7+bLvIsaQecwwJcQhu9EJOQ5vsf/LD0
tt5GcRrw4k531E7dzpDiSUng+v9oEhiXXRB7K+rFoKv8BTDPyfB1uAVL+bRhqKMf
+P8BiGoiKe3+4A1ackcZRyHxxIyTcI/qsurK6iK+xRHnxRgkir4D7b3+Yb4hmJ+0
Do9jEK2Vd1iPmtjNl/qOa2cv73CASCHm0CN7pwVU5LL1dBemNvtOtGlkKfOToQ5Y
zkjheY6+t7xevDoBIjynbCR3rbJnbFWyLscWwJ4u/t/1Mk/o+qf7HE151fU7Y9P2
oo7OUjKnR7/mxBE04qCL0U4LJbL0JD6hPhpwYnEGbjm/g4CzQzvBbmTddk1BX7tE
mDn9wKvaa/cxKK49+fMHZvUJh20b58hvJJzlHWYZXdI11DtUbWMZVuIhS1sD+pJr
gtBoggT5WTEwVk7OvzkTCwJ6eePNHeM3ktdpw1AvhPTWXRx0Bfz+XO1N5HvtGDGi
E/64RgRneoP1kpZesuV+gL7S/nUOkQPHS0ZYgnafmwerwaTE4k/QeYkaK+dDXMqR
2dshOG36FULuW87HuaxEWlVqmurgvtPNSJm/ulZuXIei36hH7I3zkRgALrfFDaF/
P4PNMBxI//FtFjAKTic1NUiklWJnbks4NC3VSEyPGPCDPSgKmint9dTjb8xEhpUa
pz0kd1JkDXG/85Lj5nIaT2bM3OjEFMCauKhnuoihG/jqREWvugZkbonHQojXx6yZ
d60clNyOxfhMJXYNSRFCqWfexqSIHLYwaOlYJp1o7DRgAoNOKqJlbkeA8N9OnCFE
ZREqSrfWczbOiIJuHJ+QxXRJ9pNYSDqXfiP/CyJF6Ix1BcguoVC/EmfH/yU/Nscd
jaOXRRlNBTWUy9+N4is2qZOgHgAYja1XKK6LwdJLk9PeC90QCXrY8okEJdrDGIag
67RBG1sFrPf4rXtLwaktp79N1thmkgwnGddvox4bU7t0qicSAmFVlG/okKRauWZ6
qe7E2Xow4FQxhy161NmU23x8JxELjbOZ7TQkUgExo4aAdA4IoTjCT/qYYLHV4XVA
cQJ+BBxjy2gvbjavkgias4F2Smae76WiLyYTv8DB4WNyoCw8e6M15mFLDjulcpn7
DgoqHXptv64hblNOUE8WCcoMKglBqNynurinjGD7uQ1s6juUKCN8lyFoJt8QYbBS
d+R/IGDS4AciIsi4bFdM2aGE4h9HM9a2OE2NzFfHQkVtV7KjgDDCjUWJMkuo0GuZ
Tu79wU1J0gk6oo6Pb/24lfDItMYJ8bRLud9rSqF9cKLUUuRQlM7Z0Cn4UUA9pzCR
v6Z5LnPOcHa8nyu0NjaTNhJpRx17t+t+o22eGbHK7HtQGubZ86pp6OwBPh/5DU4V
L3BiwzqDqXddkCJgRweCx4RCIAqDNLW5Fjb+PRQkR+P6YNmxayxR6ds1AxnMp+2G
L2gESJ61BROvgTfkocHLfY45XKzzFmxo7rWsYCnjgLRODqF2i9z3TgHoMlmWW5jk
8vR5KlM1dsgMYqD3Uggska4XJu3pNOZiCAI0uBJVUXobFcKAuSnePpn73E4rGSgi
O4Hg7vWoWZ+VMjzPUfuMHqLqD2YWapuN6+QLSS2htnwcsUG27L0/i54GgWkW9jOG
iQ+NxcuvDYps10bfyBVYeYB+cpYUyYXdnBfL+cxX+k9I9wO3sOAFBnYdVODvXkGt
1lx/8tjUJ9XzQrT1YXwsak1V5hW5BqZBxML+woiHMFyTmKGgyUdtoaP17jmfvddU
0VPGZ1V9qeqbnl5xvNw0O4Ew5gM3qKnuwGz2HHFYaXmbXfKoQOXUguCKdEVJ2kk0
Dt9l9dnNpa0m2rYuhvBRPEEVXF0eO8BQgsGzcPRW9eJgbOIcES14CPUmfCOXLpBF
9nok8Dew2wIMejqIQxrwappW9Pjmeys3qAOvUKDgLeNL7zPLAb04VFibc5BvA2g2
PKOLWkrtouyddP/A3rrOoY/bqhfsL0kMJsGv3kCrStV9zuiHg55wu+XiidE/+mvo
0BCjK2Zro8u9HM9rMP0W/4E6773SU6SIraoxU5kPTi7tAOfN3iGpUGjQosntwl7j
RkAfta42F3Hu/LaW73xf2aLOWgwQ8CNpxwoHiJf+fuaYzMKct6+KMjrbz9h6v0sQ
43unMUQpMtz+kHiWxRxex/BiZus70QTUECg9pe7u6Jz7ERwia/xcjMn/8vRY0F4+
Jj9ChvjNvf1eTMDULsYV2J6NUSeBdz9rHpkxzZByRYz/CWXAkE3hFyeEtuGRHooa
2r/qloeKoJb/XRFx9vrAQOQP0PCRtNAy+a5/Z0Db/pm1zbeBo0GjiBwjYbAW8hBj
E6wRjXiyAjsgjcTYWZx7+PGOXNk1HCQuR+pNmek60WJuVot6yGFt4qhne/wjSpi/
8xevKkH5jtrTLfOJYtBsNEEax7lyKm1JrM+uRMLCMDrBzY2WLNQFEOuQYaCRwMFt
f73dGFWf+P+ZSudlNkjc3oxeLSWzuhdjnfyEF6L04+fUgRyW0iavIM2o4gFUKaMC
XMtMewzbqwb5+u9p0h1VWm9n2PHurSt7KiWVbGu4Js9l52GyJg0te9dyPHWso0Qw
PmB6XMT9/JhAJHeLjpteHlt6OWS8ca9HcblG5eRrIIjmhK9Ihv+7PShjjJfaBTqw
TWjEk0tWjA5BqdQ8/380Yd2yQBX2Tv4IsjcbSCPk4rW71Gav3l73TePe3pk1Gsrw
aenEPswRdPiH590zs25GT+kj5ui2qTvHALQC5L9AP+v183/TLitpTPeOWqWNVW/E
q0OvNn4wdfgNxHeeLz5HXXgi22hq4gOB6lOEy400kA2Jn8tmRAqFvmp4sedPHR8e
IYBY3eh38QaMCOucteVbVjO8KCpameRRlOM+fKBlbsbdVttJ/ExNRbN0hOjHgUYt
jlVwLAPk/Kn79p9ZyvELSaaStuJ7nQQmwtIi5VDEswHfXmBzmQ59Bi/42uc6znSE
5odRYbH7LfY2d+VvHtUKDvsnbQJJzaw1A/bwZ2aKGSwhYZgtDjqy0tLxrjq0MwA6
ycTsdH2ilE9gTxgUBnIrVHDwK/DtedOCgDE+Pk2INrcsWS0HOxJMHtebzLTg1WZk
BtAhWl0wllw9DSIfAxKcSIc1+lvX+/mCz1ICj0PheyeaLKnL5QNijd3m/CupL15B
yYC1uFjC5bpMuDarqEZSU9bWmoWboDlmV/hEpRpyQW0sogoaUBrBdiMVgdLjvEne
xl3o1MWuNiuoqSXnvgNsm7KSe5wIfcC9PxYgGkFm7cVwZaISZ5IDoxT6cqt1wmTC
Bwjp8nKOu/R3pRC0EYrv8aK2oe9hh+U2y7q1SnB7q8NPRQc1t5Pbkv9/zHzEFIk7
1QSy5RamGolAP/E6erceIcmLL+lDPlAz7WzSA/QV7/bt2+YmWWS1bmJuLBCX4sAG
eGVljK77nxN9Ej9crdBEP24ouHoOYNwGARVeYfx54lg3EZaEmK6O38wkEkgUU/lA
z3fuGMxdi85t5JYe9/jHXsTkYtTjddCjprakHN84PQJ+8I3Zsf9TwEb2ZSuLHpwD
OxvZkeejmwu0O4z5AP6uA8NpnROZ3cLL5BsdC5r/N9Z6ZjBzAsy8ZIQuwfw9ztuO
KKphrofFN250CTAbCHV0DMrkBKO6R/1zSamW3rRLaSnoj6kLNiVnLlwn0Xzjxv44
YRAK+et3+J99FDw3XCLKv1TvdQKTv4NIRlgZrevDB3Qsuw7bHYuttxioWlqLefbH
dZe5x87JLlvuVQXGbXvkXuTgmGJyUaqDilJjV2IHmrpC4OSfN/CEdBhtul+KELbP
Cd0AUOiSrkdX75neZyWBS8pbiHJsjo5IXosxicpvF4WzZPre6beNYLJgB+2Ex3fa
GfUxRPuMypYFd/Wzn3P5+YroM1WSaF5egaN6+OgLTZgYxFXhOJsfEqL1bqOyqMBK
GwdwHRHC57ngRKWrU3E1yGMqlWruoYcVZZfQcF35ixd0BYtmdM15yPDiMPqYHG8F
WKuETCxiAVF220duVKMwu1yf7F2URSqrGeJEOVcheSIIGMGbLPdv59u/3DBc06xR
R7oI8p8qqfMXK178CxfK0F5DIU6QpRK8gxqvmnsnY3G86idQYtvoIned6j1d8GHL
aXMDnPMgJur8PvLhpsl+GNTOkDn0/WvdlUhDB+K7lT/IB2N2k4ZK46hq2H7FOJ2V
36bX428wGd8rWCMppeKrxnTxDv22X1FNHCj8VtovnpwNKgJN8r31GZg2IV14jhhI
pWpJXZ6iVkCsapgNisixuNnbDNQUWZqSuIKmbGwvRPhY+uejKQVGzeCM5PWxNI8U
LwHfd4pdy/uXZYSOliUjXj9oc8xgLbDX+yP1ZxtwHrl6IyEEsMa1/NqfbgAMjDqO
uU9v6ZbUJPNEUUl57sxrIyoqvVbsmosYWFx8suAlu4VUym6pv/LGCbOXrA0REatA
9MfoRFJk5jG5K1UzLmYx24o4KX9HCBqUIW+OLVeFL1nJNKNTj1fMavrypc6zT4hv
4FERCeppQ4FFlKrJBdYGLkW0QVzKzQ1sp55STxliw0C4nomp9ifELyV84ZUbFywk
b8xzRv6wndGN7uRddA+gJb+uT+4sMfWHyrwfu8BVKppmVsvtyj5KovJzgNmkfU4Z
6iuP17qmhh12NdKbJP7ZnauvQOHNnTVu/VxdUigv7kMG5tPJz1hDfPvIYbwk2xPK
O8wG8TIzrhDpD8ovuPeb4hATw//MNanQKpwJ9XfSlkz5NbiZdlbHNfK1fZlwPkPG
A8DQISVy3evyTbdt921IKBmgwwxjEcFbfKR9v5TXW2bXlJ+hkhnUkzpoX/Uy+hv7
83GTP4j4oGhHKqSBOCc40mLigyh/TQQ01VF6yHowP2jkylNb2DBlhB5BodWMk5WA
8PYjnTzfmCk+STD1/gViwQyPSkyS6YTEjH+J7Kb9W2HuBZfeR0pTMfY/OLpm8Lze
4TWc2xVIHmpKU1e0YpQ+oTmo6MnHYLKcnRj+QD/ebJtpN2GBXO/+ETVb35oizwPd
y+S7loK898+JuWX7k/La5d1fMKQ3CwFrBLgsu3C2H0XkMonbtedlBgfeffM7CHHj
/0JavtbiZ9LB0Mg9Ke+tIv/dmQV9m2RyTNaehhhZY/AssYsSFhsMZezE3yd87SP2
YAQEd8K0gQBcqZgWAqm8thrIo6hllVvcd2JyO0CDXGTp+aV+b0J8W1Pgve8s7LJS
1cdFBZ9QHItpdmE/KDMPzG3jrFpFPh5ak0x5uk1eVoXt+t9wwFITpwnOQSN7Z4ez
5DfL97Mcwmj+A/OjjJPft5HEFf0eMp4j2aJwiTgQnTjH5DIQ1KklXKj8WsqcQIrN
pqcK3UyyN8Kjz41+aHZp5mhHTBFD30Lh12pTaWnrq9Jr2BlB+Kd4xHKMo9h/PAGg
Z683rbVDuSMzkMGHKwqzy+sJztMp1YALj4AbFjRJV3NVNzl0rakaMdxA3NfJocVN
y8bbb4xDMyHtm7SsWiLqt0iXqkMxIlh9+xh48MV8/x3Dl2XjOBaWemGXLAWLjBVv
fwZB0zAji9eCuDwRz3CBrQ5mkiAxHLbo9N7sK++sKEdYuygxH3pUX8ErVmV55HXz
CMDPoyrvb3v9l071qMJiZxK4BvzkItL/S7fiqvLuwul67TX8Mna4yKmXBLfZ21sk
f2FeusHe5nisna5QDXVKKXdvTtW0YBOzgXy4xG0acS7tUnJ56KtR9si+wS50eR/B
IIMLJaJZVWbE1igu5Xqxk1IlxcQhbVdp6sadT0YY0Vb0PDHwmJbSxuBx93no1VGc
fgcE+RiJRDixdutU56PXqltTeDFZWOHdjJXoAoeCes+v0raw3D5AsOhGF4Wb+BH4
29QnRSznKALUYmqm2nrlgR+IRQnQsS1XEfp94wMTjue1/6Bnv1Lz3hwuHwu0OpzZ
SB+ZYBLFWFSeUl9TWtalPcSGmA8RFWKTsvznXWGoZWUIiz8Kaaiz6IXrVX+qw0+7
9sN+O67EaO73TAHKsNJGEO6xCOATYv3fRMEu05XYQYmxnu8uUZ8D0Mo5dkv4IkDH
6b0oukttO3fxc7JSMmLhdm65VohsYmXS6apHmaFHSJZE3eRA+rZ8WYUrtfLdvi7+
HpZnPisTcgTiulAj+MKhK4dopfRNz6hLz5dw60hQFg0GMg55xFSDqvWUoJNIACwr
6022a+dHIfQsi8SzMcW9YdzlZvJsLtTVrEUsD1tIiZU0j6HSca5m1eTqTL0jLIhg
ETR/CvuE8t1CStAOzt3Ve6cHeIRRAJ4KZqk1ZneJgl+dVV8xU+twFmERyhNFLlKh
gaJONMz6R/VWe8dFLgHq5x/KsbUTflwX/i3gbfZyNofh+00gAFI6AkbsayW4U4Z/
ljqQsAeQ0YXZsDCHw+MO6EuuPfAXOxIwtbX4CmtN9iT7DrdFbZn9QNbrs1G4fufp
MNv6m1v5XECiez8bmQ40D2+fAABYSfMuYd/mpot0z0RbBJIwuLTde09zBNPgb0Ko
oiuW5BPZI2h4t3hkS6jRfyeW/d9CMRcWV9UhEMFLnoF/2n2orZdI7lv+zcR8pbBY
7hNapSnPwk+QFx8gfQkafPYNOPvTLRzLgB6CObupxBbjAFp9iS/PRpKzCD+pt5OP
U3XYFFORALJXSMReSa3UQK6sN3u/c8y9gDNC1f5g6Yv9tZhbplHKW07JKhrI+OUb
r458le+mtP3HNqn+cjmOIPJIqc7B95qZXm5PX61gM/2I/CN9wXnPFLVw6K12XXer
fGYDvixl2jSqECPFzWo4X5jMYlhMUVg79X9Cb1gudKTYKds+zYCf9pq7a2QcL9BO
QHFaMk9hvg1jlAuqGKe0/u76yjFbAtRLJIRWkp1p7hEfkUQ4/P1vf44CEVCwd6Vh
BJg2r8TJhkVcGQ0t8wzbOwSIRTBaj64O/in9VdVxDdQqHdY/G+nZbiJ15h+HcbFt
wi2mUPw4E0zTHz6VNDtAt0R1+V2kNwGG3ndhk1X+aQd1lzsReBlf8WLPTQKURHu7
55p9LdaCozeqH/TNw/oquqBDuAEqs1xW4EhtEC8SzCiUyd3/NHIL3UQOcgapLwiL
WH1a0+CiHQhtt92/SMc6nKgqjhlQTou1afcwMDPHoSdwKFxDtzaEvpJHJI/9zrur
3iG+7rHH+Gy1COend52FYeHydt0QGjj9mf9cJWS1oS+FdlY4covJEtcwvh3WscC9
P4kouX/p+j5/pJKjBq1MnC0l4s3ftTDLvHOMPdsh9TI2u/I3zitDuNbnWJYz9U9S
+/wp4NWHhZ+geJCHYqKROUkeCeSoqb6yNaFju1WItt8POGDIUFdBdBeO+boUHcBO
7S35TGrbzlH+5FY0BPA2OTIZ02uqGkGs4GiYv57/4V4Bp5g8SxJOOAIfvqfNlU5g
dvmM8bIPbDQaBuTd8mSeD9EhmHM/y/f8s/dyB24yO5NZnkT4pI3/tBiRuPXfqlM4
dZgZaScCLwnYetPPTppAjGjG7Srno51GO/3ZBMdgZuTQNerMNAaQ5TsOAcZ8yLF6
oPfyjJcy1TxT7tr4PFjs3DnNGWwq7aGishO+GNQb9O3jo6BAk6BY949WkrJH+CAq
J+opHqsb9C2fv126/l3tklT981mvn6h2o3AUYRbnovYAUSss18dJviJLFLhiyJod
CbazK+9lG2SMuEJ9M0Sgo0tksirTXZpPUejrDh5yS9KXRGD2/feY7fNWB950ZWjG
r2W6jqctDBws/PYmF7wWkSoN8Mtzldxr+72iRmvAV6AEx/xgK3N/c3kAoATYr51F
wvE7JrNhr6p8mJNpllXOA2gH7mN+kVQTQX6ID75tOJGjTnMB+C+HV9jTDzgWBNxM
qOK7nPs7FjbEPHZa0ZAYV4B6ysRHWnORO6FXSRJ1ijMfZ3EAPzz4+cRgDLWZl5+N
XSFM/H3fHAENzuAhyuYz5a02GrfBw3SBCBhZGpCov+g6LTy2g7CcNblL5nvfGVmy
uyxCzeMNMjCDNeFWwUFh6RzOVPSR2MiBOb+3MOeORwT7c6UvBvlXKN4D++8H3MxW
RhjgTKhqBNfTqPGssuSSI+s4MkDjNbS6RCNx28jWUfPeAgm5phfoLjjpDyAivvOJ
VqnQOZYEVrPctcFjmkdVlW8JMnLMtQGrugtllNFi1AMw4PTQ00SrQmgLxc5HRv4B
A5C/7c12Q+TrJRnGoyMWP9wpsVU0+ml5cqYs0ge7Py+qlOuOq50L9fV7tYMNC50Q
jUl68Nv/NwoX9nhZpqa3hCUCWz9pOQTClV6znye6Uh6E+8gzRcnX2dXmbgd9kVpi
nwk8rodEiyLdiVr2A8/b7rZMfzJQM2z4VBbLLuX9gb0DqLTX2e238uSsXm66pazx
dcs9N61+U2+NhglnmLgHf2oJphoGhUQo7rjh/EPiknAZfJRFBVdVmqttbOCBtL8e
XH//oRdKF3hJZaA4ISmMrW6NxzAJAfDlcT1O3/ajIYeZ/woqJEjJJN7gWgpUZ+xa
K/Il7YiHdqPHZYLtLl1SRugUDRgtxfynSVZDavY9CD06Y4ckd7T9R99/qynBWkOr
/tEz2mOcOBifYYH3nu5BWfKaqL5sgQL+gJLz/0P88lCMvmDCkWTEyIBcpwpFZSWN
p72tm4074ujp0ttVL6FlmiQE5ocjQ6Ifss/ZJMsFo+VAB9Lh6DkQhdXDrAgYivkT
HVmdR7rmaoHv6lgHyzxCWoxKtSbHQ1pV6abQxhOt+WU3TY6Ftg9Q7BOMWuH1dX93
Bj3iPleJrZxZGNbm1B7HH/nOOVRpVFKJZSYAVQvdruAwaUHG5mVc8Q8t92TLuTgi
l/Xt6zVpB2v2WGBDyKUvVHPe3VdS6IxJg0Li8irb2FvQWtdYM1IvASfbcA6tsdV1
yfxApm6oVxxsYdCydKzQIFwH1rxep81JWzwwAoEia3K1fDDpQ19OSmkKYHr+Hie3
y5PxM5fdOj1O4znLLFNFnJIef68g9i6cj1F7lkDO+qfNlwINwHF3lSIICOR99pQl
1bWFY37TVgMzK2W+DVesof4RNXDa3kmPsK4p4NQhzP4o2dWZRlu/A4exdKO6GRQM
Ng2ONsoyvkj+BNulvx67O+BuIN0poxO27hMWxlk8C+DEHJF4Xl90Bbz7wiZxgilX
hruqjc89BHB9nfE7eCbKwk6Rd0TibWPPgosyxS32b2XRFUpyYN4qHi5hh+XIl3O5
X9WJr3CbP1XkEq86TIoznPijZoNl34PZewW4JPDwNMX+WogoTnlJhbb5Ma07uol1
1lr8knRNE3o+4t3oC6hmILciSPoedvjIP2R0iNUNqFGPYlJsVZ8zmqUz6xhwsN3g
XmW8QVb1Uokl4I02yqTZbLmjUxUMHpM4sdB3yZRt6OGLsi/O85xVrBWKkIkB5ggj
zfy2UOtzn3k3U9vnijgsdbBxr/wR0WNJNjEaY9CiIp4SYGr82AO2BDdmONizl4YV
lv6z8bvRHVJ4DJ8Nkgk+PzT0Stcy8V0ZADgNGc4Sjz9FBIQN8zjzSHJGp6el1WC8
CpjZ8sMfzr+Z1ALpya9ubY3qaxeWq+U5OjaY8LzHODCQDVVcrJ4QyZwNCwYaVaJF
5n1hJeVa1xuAOXI3d+Wm6JrB2+QTagNT4kjr18Pe8fPpEIOHmBtR/FycW2w409Zz
7yA2TFy453DzsNuKD9M/AllaSochkMlPg0QVS5NcCEIf/mKEAPCpwvN1kXHq8slH
zpmTHyDd8DK96BaQ7eelcnDq3GlUb3b7lxP1DcGu3Jr9jAf2GMySSw0Ca1HEtHdS
GRfE5IE0pwLO64GNm5ywhLJIcaxL/yyDd+G8Eo1t0JMqeOpZNjQCY3g/sWmI5eUr
6uvas2reB+pSpk4r3zj4BpCwdpfY5NNnZ1y4vxWyJrvDdBV/t0dhCLaMP7OR/xet
Nqy6RwiVEhop2XgRrzoo438aWfRZiVhAo0IlDYBmYawM8ut09ytYnIvy0ypKNd/e
gzgnDmuE9DRrn8ODv4uMQ3E4/1VZWEDVuQCcZSq6WlE1aJkVk/RqPHj+Hgj84oj1
819tKc/3jHROHpHhsO0wtdxcKgJGdfm65A92Itw5LVUiADtLofFAAw0jSgr5Uwd0
prPb0rYxYTpJKBS6rOfSsMqBWwkCI7upAKc4a5whpKLoWkoGiEBKdkk9Mnv+B/6P
uUFTCWTw2zTvYdmB4UcNetUrRDu5NNUh+j02VLe7ay56CuOgPdK59qVLOxdXqNdV
2pjDZAwmScLgBG9mQSSG/k8zjqVQOlye+2ppIiYQIMhwf7NJD0B1yRK0LXdkFgv3
S9c9FHdN/vNYQddqF2m1UHWVFcZcQgEqXkDfDvJ1rTTO3GVp7+ur10FSm9eiXJxF
f3nK3xz4mOU6u5sjBMY199UZapDfFWLBkiUus5DIy56kTvCVL7gYJFSdN6u9Ajan
IVULVml1LGIAmTuuACrTe0/FiGftO2ls4PfDAM2wWLFKrN6+xHesz5xYDZjeR7wo
nAblJgd89GGnOFkGPUYgK+J5ZexqfHRZz4p6E9MQzEPF2bB+MdChAEu4wg10GtFy
NUD52VwOfwEV5lZbSU+hY+AO4satCuh0XgacFfLQmOUL/KRtLFNtOLw+C9RmWtmg
gCwebR0xqE6Axjw7cL64uOjgVTBreHq2Dc3LxHmIYjAYXvDDtyyRpVbkDHsdZs6V
H8hMQZANMbzo7LrliCnsLqGYgMk1+9+/PvvkSxiqUNEyUpED7hEhXMMd+49efeOg
1vR2A2d2DMyURsDNt9+Wepg50phvvCErV8fFKWXJ32b8yq3gj8IGj66mFOAhyRUX
TKOy1y2Dgstil9nEyuB79HZvgkjJuo8ZkMG5R+s7jz1HcgknWBBvF4eBF1vEK+yd
F2WqytOIXeb+vTJlCxE7E16taktjIkH8UIic2HkX+wYJjHwi+f1Oa5PuBD7WJUAv
MOrvj7WSSj0hv+7awikMxTn7H6jbXuOMW+pJTPsBTf1K7nBcMNzXXu2efKkVnmva
3uIj8Srcf6AsqMf7XFoHSR/UzYdXYN5Ve0XPtL2xsuFdelR2XGhCsyaViUFNxKFg
YCL2TV1vQs8YjHx+3nrBkDrdkkLgAw2JV2rTCz8UGwYz/SzXwtln+xg7pcXGPWMr
TR/tq8vHm5H9MvOjWBRdqGjtFjicMUGAN2d9RvG+eMwdoTki6PhxORjEQO4hq0Wd
obrj1j7+0sbaLGyZGYcBOenhKXNmjAXv4iPfIcsYkBbofObtUuhOMjPB4E4AW9Ca
ufGfyrd9y5bq8hJ0lOSKCgr8oHlshseIyD8guGdGy+dGlgppGV/PeQ0AUK2V9fJ9
ZcKJkhh+V3/8d+bt5LjKsmLy6zbSf2+py9DktExCpq04IidK4jreThbj7KfW5HbK
0dUB2TK6muQ+ZseLU82Bpw5A5VZu4YUlJFzJV00QLJKYWF7apZOrfcpaz4pI6qZY
cRujBHeer7rsbM84YEzgfygcAf5kbXwvNf+5fUSbhX6W7wep7qlTasCjfS/DkGTD
3b4qG61+ftJYuoWg5HrzmxIvHoumUa+9YUwVpLq+fDtiBx9N2amKjJO3qM2+Cbm2
/sJgnVOZiWl7VmPUriVqEqEqt9U5P76FITiozKXpAHQqhxIjvZNfCVschr3JDONw
YHgWfwH+rzbkSTvjDpoY7MmlvR9Yh1JJCer5wqWLij9Z0LSyUg2M+RnsIqitKHna
9zrzYbAfXT5gD6akl9P/yo6RjmeLmGlvLtJXK7D6Br4OVMfn38n7vTpI6NgeamBp
M8MMQCD6IjdyMh0vhSTUoYhLbStkmSXh7unx5yFUYdbIEp2r4rhIpx4Nl1V1xJ7T
t6/TIVlgmMP0ZWnGBf32KZ11ZrfFSeQQOUTtK+DM/gBlXxHxh+XIDugSkNng5JaA
TNAfDtzYgv+q2Pk3LCcfAEGLUmIox880naIoDsfz+zln6AiUuB9FTlAd6BefAq/9
jxLrqIP5nJnhZA351UzKQnnyCU1PjWK2PmafOzs6btSIxTRaQDVpfZh2PuCl7nvG
dD06BfkDRzQFSo24i5zxdGZEDEO9bRzsLP0xH12MsFV0syiLkvgeuLwHlh//Ty5s
5TfZQ8YI9ZWg3F8N+sIYUw6BwwVVLgaEG3kHRxZHPzHLc/pveafhLkxXzD4IKMkw
+0m/ZPgWgyrvTRFfULfu9WaGUf4KhtnI2/3tIaIR393MiRPiB2qSF+RzhAlqNNEN
E2obTbbde11W6s+LhwllWDDJ4XW/QOfx6DiFFboXuada3tl3oDFtCoZ8jk477j+p
B40N6wq99Pd/aQRcO9TrkW+QEuHw9GxkEh7gXTGRNZilPRJnnRQQ4cWL6C6BVMV5
4CdDO4Q4aUnIAS2q/5vekKg6UQ1j351FvymOiz/+do7Ic8Il5WR5DPDr5nSqLMSi
vnb6TTdk29bOlFt+oIU958ctQILGsa1R1CLGEvPIlX1J7qIMhPifxQF2/BaFlaZq
l6HzB7ovVLPP9QPvpRaIpXMttrHpnPdXCb9RV+g6AzWixel+s4a2DBajKXTzNZ/L
/849LOKP+6Z+BTPiWyqpocQJDftVjNzYHER+geFMT1njPUFtkoNxxdZVdSFttGvG
LmoiezQKsjeJnk+gdK36zwVCoEwtLQlyysLs3tKkMAY3cWbW9PxjFXwK36u44cXt
AVKh+IGjCLLwsOMmiLOKRHQXw+lwrU3gz1NcqqOY+2p7bdDErpT0tnrnyQzSahH1
Stee0TnWE64JqINX/Dt+JTyP3u90IjVATR9mXeYbVQLsw57iQPRKSGqv+Bk0gOIP
biKFE2d/7eCKn07vMedClm+GqIektHbnF3UmaaS7qXP1bZxgj/1H9GJSi2m3fEcQ
F9mb+yEYA5RsMZxgtc22Ei0Z+qwJj278ED9jLEXapRVSzoYY2pqRtPyVw12eTTTN
5qRlhoXXEliS3KqbGGVKf9ydmrcB6p2Q1i6RN2pxZE8Fh0eS6NqPhkKGwYXVFspm
KqvIjEmlsA+n0B+aT/DiIDEYuyKt5jPot6nbSrDbdQOjki2eyhpAKxc0Nrak7YOJ
bjyaSaizwR3V2L6eeUEygyyZL/tE5ha9VQJxx2CUc2htRF7X5/PJTQzNLXHU4Dj5
HCFOxI0xGkzi7486A5V77WCrgMNENqJzZNV3hixGkTMIXjLaPgtVmKpNHx4a+93E
X8iQkE9rTSKeLvY58Dj5ZU8INmTlCIMd86ZQgQJIP/OkOLMBXymOQbuiCcSPmsbm
/v8yQD2NbWctegLaCazpRlXTlPcui37jctJgKOldxbWXOa86AmrjicYq4JO1IrJ3
cC/i6ay9mwpNgNrTd8KxpfefzQcgU4JcufBX/e8SqN1Eetj5xAn0A40Q0+B52tKB
K9sE+HsIKI4GS2uh/TEPUAvbYP1rklQuEaomu1B8B0pueenRgIg6v4i2Ft3Uloke
WpYuy0RGv9VadT5LnJVb9uI0dHULkWqVw4lQFRJPBmuPOU2NAKZOKy+tDi+/wTgm
6KaS6om6zFpBsm4KGHRSBTjOL/W1QMzqHj8fh4C4Nopn6dPGcWqmO9YuKfyoZ7vE
01pDayqXnwLYEcXi/sd+RQgFxMYh0JOSSY5hb0eDJ9uMTeYGSdk4WduCI2Ql8b9O
nyse3g7bWAULM4Q67V1FLnH+crsAyvI8yZjvkdn4MuecTbz1/+mspL9RC5ztT8QJ
yozKOXJdlJ90Fvb1am0J0rcc/NBAfnePmjTZThdJH/lfvda2bsprhMwa/vCc8U3I
v22Wg26SPgViqT1SJZJSB96ASWHN0xhb8BEO6hGaRifq0m5+h1z0wRTw+1bT/PCL
tTZlWs2HBu3KxNwYMGt4AMpDpVWWAwmoUE77ksmbZZVsW7hi85/FTa4mDh2yQbgT
qW+jqMzIrBfC9/llbk6/ng18Lb1uXrMi3oRJTJzTVwGetW8wY4NIArnzYaSKObVy
bKTrv3CC2/9TVlTXFJPA7Z9jfoy6obavo+viFGk/rSY3TFKPOciAaJqcYW55N5Wz
f+Gmfpo3dyhhdYOOw+8Udn0xyDzrFTvFp7/Wf2psvH08uiBt9qZS+8FxDl0+1xPG
BWle0Vz7CHqA0kUN3SvTMTAtFSizLp/lTtj31leFV6QSwDxcEXpdVxUuhDOVubTb
4lZm93ab9h4qQYlpXhMviYsrdrZrIjVbd//6ykpek6gJsG8s0nTMPNyJNX+dFiI2
6uiNHEV4526pjaBfvaswWTFw/6Adt+bQADxMBNQcEfHieLjWiRvPmdudD35qtLwy
e8duMYTZL/Zrb3NWod57zJh8CAs6s1O1tbb6HM4ght0vumRbj6o3Pn/l5dUj6z5M
`protect END_PROTECTED