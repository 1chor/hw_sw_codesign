-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
SJBSfWEJJcw6jRpZRzvY1GzNjawyHl9OagYDU5i3dAo8aITE15HvtUmUsbbuUxo2
f/BbJg4Ge7loaUmYwt947OxhBEX6NBqax+UGZ7xZjFYBWNDllhXiJraxS3DBWyax
m2A3ydhIzFbVmXcpjFknvkBqh236S1MoIcAtFYIV4Ho=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 26384)
`protect data_block
dxCtgbZfpZ2b0hsuMbMllnwyy1aYDmLkvADsLl/Mid85BvQLf20i6qihUrH7zTaG
SYBY9FyJHsRwRJfx05LQ/FcvENecMOPse5QqOY+cX3IwmTEPPdVU5DChA+d7sOHx
fNdeyzaZ1oMnRtWBhlibVC0AImGFcIPNjBiGFrnUDD2eONXVBnadKvGgL4PJVwkK
eJpD8cSUPPWUG+pEAcKTNswn9kDtFAXSjoh7rgAHVlsNmJbESglPJtmZbRIzrN32
eBDVaxVfUjkdMaqjAmhwYPhkvniOGV0p5/oRZSGxZj8XS/7WHACGe/bALRvQRHFz
+RW7ntUO5s4eqCNshvnBP8bw7Lt37SLtkpKpSzNdRMMjufgcIlQKjtz42AAcEWhm
wHzbJbUd8l/dNPp1uFtnp+HcAykv8A1yKHUL9hDVFtUkbO94raruWJR5x4hQR40C
IHxCkxRlVuMRiI/KLWFaxhddGUr6bVUOfVeZxC8BMW4ATBp+HHVI6KwqNfPecP6k
ugmbJzZxxPAgQnRpgvQXNHh9Wd5bpkSTUoM28N30oIHcJOSfuZfbN9SQC/YWDzHr
Z7iYurqR1J9VqYG+4Xjo/qujA+5q0PdLWQIWpy3UkMRmAjHz2Fujgicn2BvONc5+
UrBRq5/P4o3FOAC0tQPLePmBlyt5u5hcpFQXzi9LJSyr+gwQIbnfxOeBvt0YElCP
69+/MYWxzUJDZTs8ucVcr65QXj73iuG4IPGq1n/HRZ2e01aefWPy7Cp5ymKA+omC
5C4dw/TJO5ghLT90pwyrBXgiYu3b/8TrVBtg5Oi0EcpYXt1syc+zovaJbIKsQ5r6
IqTgttdaMxNq3Nkoh6sYPYhM36rVIFzti1KXWQuTXsoglhU7gT7mLmle1ljpcgUx
Gm2reAs533jJ62f4h4B5Ebj0AwyeNLSSwTnSHHZ79NIwsDpv7zJ/FoPS1DNwnway
aKjNzbJNyCyURjUoF7EdeRyiDFnCEivvXPVxFdLfx+BQB38c1nJ1F2BZhaCuUzSQ
no90pfZ2qP9ixV5GC0nQicsOxqESDFKkNDCTRD+xW8z8RiJ3XwBx4mmrC6NKRKNy
evXVqexbPUbeycP79Yxjv9v/TCjEkEw1ZS8kEEFf34WNbF4KWcJxbYhlRTKtD4v1
o+rvksx1A2vLs/RmvQdHHpWaaCcIc/ATaEZpckpDV5Y5nf/4dSMLLW5vO6ZYV4tv
I/n7Os7zHcYpqtLR73ZotrNU3dvV5zVN781vHFEFs/vHYov3T6lmjAYAR2o0JYr3
/nEpbSfFvh8gHZD8WE0ZsKZWkL9q0C76JJ3C4aCYofKRbm9Q9pxMm+7XB92OWAds
EbfoMg4N39aHK8P2qnaoYJFSWYMyS4HwJcbyxcuos7sSyCFv87ZAzhRZxjdzOp/I
EjyI9MsjuQ0JRgtxzm72mkq6TD4RB1p8D3XKAeNEwuOtSAQbcAYx9KY7M+Gf/D4+
UAGuZkU/S9trGjmpssUmotSMlsLjwJusWupzAx9v2C5GYZMONviRmSpKByMAm2WT
ZfBpwqh84uoXvOsRgape+pD1p7tzadod63ZUs8ia3O672ruJcPfiu/wAnjYqA+4I
t22ZR4U05Ya4K7hZz1r8QBrYGB/PFL6IuOgJiczSCwYfOJpjuMJ8rg7emx4pJ/ze
gu30ykPmr8eXF+bGpD4ZDi8/LRyYXrPSWGBIxVLboLmp+vd41U20S32fAKVaefyw
C1dksebZF7Hej0Dbww1LIGuz+LKMh5AITOtbdnVFPcdkc+FEIasZOA0sq1dJfVgS
9nCVuv/nrHdihh4cTurjaLOtOANvr4lRxHk5YmM5u/GFOHCxxlgxzgB9vj8QzQrF
w5ri9y3iL/yTYCE1XiUMHEwYJ/81xDL7Rsd2f4ozp0N7h7Kxt2JYC0Bw2LPZ9IXb
ozx6+hFR14z08/8aQiLNNEXrl0fJe5I0e+YhnsNxdN4X0z45iL8B55Up4CKfiFxl
4jIZIHGhXohk9RXWmWsdq5OPt34gqwQY1hn2KLHN4gu1WXREfz1jCkMQeZID65sS
6rH4IStMU1TzNQIKzHQ2mR9JtdnqfqLZDf9mr+rRRMnJRIvq2SpuNt2MuWmgKWBg
FWtYKonK6yCjEKbiVcVL+cFUZc/X8qOWuwtTN4aLM9Wo6UL46yOT5rd4Fd6ubjnj
nfPDDKXl0hYG/hdviclJah6TjQVYgo1WoJ9e1NSCdX9k61GBmHbKo2rTQzI4YCkz
zoP6Qlaqh1PENLOQAWT1OZ0B45F0UwTBjk0aJc9dhpeAHEZQYrXncGfdnttLQnGT
+kHGbqgVZ0pyS7Bt/91NXOhQ6SAOqvJkBN66NUWYX6cpFMGU74U5TozCvxqnAh5d
D2O3a6bMd9ZD9Kohpe6reWlkgQeu78Vho2d/kl67ONXPovf1VIX+JhhuFOcuo7XO
67nbjC+MVoly7nSohlyJEnwgqodDsBhRRwt7ZWCmM4jdglvIgJPDZlszl4lyMkXF
8MMNTbkhWEDHs7jDs819p5pitX6+D+3ANBfRc2ljWdxGQOZGlWhT/5PfcO21vVoq
h2HrGB4xBeRt2HX5Z0twez70mesr+q8Of7c1W89kT4wZC0cEMYSurpX1KqhXVeTg
2EAQ8brIPLkRqVxfbyIKjv7lRxZKvAFoGy3mUxHlm9T1M1QKB5fdcvXulKqUEyWY
Hvou4plWJP4Qwrv9LJBG6MI1F6Md2kl/cBCCOKQluYtebHAdkGjJ4osEg4cC2C+A
5TK+exWjpBJ6AlJ7t9mCjihuz72P+peX6QNKss3+YvnuosTkHLzie4U2gYSP6DUd
6goSi4YZWjshZrXyqAAoGH5L06iDzLISg14QZQKi+v2FzbPH7muLxvkOvDRKca//
WwhdoMFNp/Rl8aJSFC2LG7VIUhkx3ZwuBTgFP+n9I9gZQh4Yl7bxz4Ng24N0kooe
mq06Px77lT4xpTKqjDdRGWtB4TYJrMmHcwn+FescaETwF+IFIhgPlptRDakZU35P
Au/oO03gjGpdNgK3Lnk21V8PzQfeicne/dKH1jUiPDK6DL95/jY3Mq8dIbAfq9fg
EcTs/QKOlJrrX0IAZ6HxR3YHzjyQ1YLCxhSdqW8DeNEe/qtKDS1mzkXBRz+m0M8t
CS3bqFSbj117MElXSalU5T9gceSClyFVVnD/QwdQ21EQanwa0MFADWD3OR5VQSc+
0DvWbO0RXQAGp6jHV5nrD34frA6rajGCKq1TzyRzWeWhrlxN8k7pYCU9GwGnrtL3
amHcl47gy/QAdMcPblALJdWv37RRMs4A5AHoHva9I5uWmOCAbA29JwqgC3pgEIXC
3oX2694S74Wf0FjSITFhF9eOLChmasl+LLN9PKRWRbgIIQhEfBe0RR1dqGyNIinz
REQ8DIpMBqxH2SF5CIvMY+k6kGR/1EmI06pJ+ywlLLhhfLIxLVxEAnY6p2jXNPNQ
24QBpTgmcJJSyUr2spU/TzWMM1aVNMhBgkbQsNR+J2pX0OTm0I/RcOTGlweBs34P
MyEE/Qjtm/hnB492LtujaKW9Au5aozUFE4p5UJmuW/7ZfEykJATS7YKfD8i437E1
KPlT6GT4UryqFyxCuIFAGxwrQR+3xgxs6N2/KBXG7Dqc8nsiPjjrPsENuWk+eKOy
KrOczURFWClwnRNs+WI8L0cxPz3vMjZq/+zfcWGoSXcvasXMMJW6Gd4Rj86SF4vj
xpwO7EfcpPdnRgfUEUd3iob9A9LlIjzFrLc0vE6lD6J+lywcN8Ox/V1D7L/fWPm6
NPUcaLqK/IVs8WWC88Npdk7nsQyMPeD3NAe2jUE4FZhZT5L1nvZU7H7cC9W6yPvO
XapjeK9w4zY7syJwxhD7aA0CaNBaStqkyJe/2BTH8qqJkbfWsJI9R1pLpH7qI/Ak
d3c2ssG/mkZAf8SJBH7+CNxFcnTS2Ps7QVG3CbdNdXvcK6L6fRH5bCYqzIHfb8gn
mQLh9gIZL8cWH9EmfXxLkDUsYnJ2Wm2WuTTRYdKgyrurEoI01k1tLlbqTnV5KLFt
LTFABB3SYZvukhcHJfg5K8hPXxpvWtUZl0bBk5+NEKpYs4WFEDN8U/SIuxbimdIx
Bd/voe7QNJ0M16Vc3OCVE/xymM6shMmUV7pC7+yV0l7mlx7rcJXPagwSA83A6ODX
okKdJriyVMH0yCsEteTmxFobJF+5AYBISAz51OoHkoDO5i6z5bnz3pFjtrPDS1rD
O3bfheAlfAi7sfBEUpXq2D+kVmjNloDHOzMdcPwFe0uM/RHLRSl8dSAWb8Qeh1PT
96tai32CRx/Gvo0E5STo6wBOy2Fe2UrjaJZ+9VyzOCeq1/KiBe9uV5DyVd76UW/u
qZB1P4tCW3EzKuemI8IDlNuxnw8iGuN8oHUp69NECf8pL2zuO3qk7FXxbbjLSmxZ
/2QqnKDaTFoK8Z32IvSXeOMnj2vjY1XBW4zwjz8E002epXrATyhkfiTzknK+cq8R
UskFn0I25uUb87ufs0n1keS4/T7lsGb/FXC2myH18gfTedJ6SPWt+fVMLNXy9fvy
yjPIyWgjS7vpejCOTEhH1LE8UTGxmSuHBalN0SltLlL1JYWMO06iFQeS1E/BRVb3
prLJYAedxoCFnaG3w9bxgSAce6jdld89j8x6SpB+PfTnzrN7G8xtv+dySi93Ic5y
xq/2LmukspePMhoqajzAmFxY7ofZBCZAK/OLKVaHUCmTgXRgxDyDDUHRGPmfWHnX
anJUNvRripkobA/RCTUJUnDXf8cmd/WZZmP33ZhSF3tK/x427lA8rdH4aR4OBlFI
XmzOPp3Q6bqkn+jxMXV6gbNxph0MVelWJ2fuWW6FBWR6LXK109VrAxu3EgBfBFsG
4vhG6Hh34OqqVYPLFhNFJ9u1jzTr/uAvgZ/MRzbst6fubflnkj/v/OwQx91tEygs
+5x/M2v40eNs8vDPRELeHhlJhGNrjYxmH1uKBoSeWFNicHXUR9I1feM2uRasTCxx
2TQmyw14bvOTV5EGQghu2+5bYPSnD3MJNQrXmSMjjSzHOFipRih8YEuAIXZQCD5w
344UH+GNqw80JKNlK3wxI8Sk42lpsyIdlVuxza7LRW2r7AkTo4fmIehFCwjKwbAo
S4lUrRf8HEmr7TzlPDSm6j27Hnulxs7pqzeYQ6RN3eVEbiM290ozZyT3nPQWPLSk
S+mhmg1jwdTJwWNaQJt6JZezpnDAjL0bRodLd1lO2dKKsrlwUqniuRX3pqm8Bws5
M5fb6jCzBaJFya2eviXOjCm+Ghdbp2t//Q4lh26QVzs9yjfLTYMm1cVT56kwGNBT
7e5x18TDG94fqvFK/zdEon7slMqohEDylzX8ILWpAOQPdQz0AyonAhOXXBU7Wssm
LKO2Jzlq8klybHH7FwpsQ6IzQXdvFHbFcL4KPnXa+/P0H30HwGjXXuNGpP4kf++a
578kss9+90w0Jis2Kbh822/3/aGPDfBU60llIz6Fpd66M1PBgh++8eVNQlFYOQgJ
/121axpC6wKn7oEdyYCt/d2UuMowKlULwPBxj+Fo5P9oKTQ/e/IpzRBzsWlDb+Rf
1P+PgtBedA77t4V8uOgTJ9vw5ZFMkENzH6RBAN+JqkRQp4JHdMigAPezSWejkoUS
bHJ25vnKEuCCAT2WE/cJPEhnOrxKsuiZ/WfqITLp9phCy7eoBcyDenzEMkj1iQLi
RpUYhRuk4BIr7nTrEz+d84007Hl36FixjQv6tMRndwFgn+kh67/AUDx0KwlblUto
h5ikL31f7fA+pA8tNdabsYPzxEzc6jL0OR4vmTixYdRlO8iv1EwMpp0U1LTwAltJ
3xA+/kmMsrf3aq0ik3s3XMtklBflnovBn0s1jcy9RYh+ooKpD3Asc6vXLeroWTuB
TYsrOGTiE9s0Xfeordkq6b9SUJy3AmD3BW2JVNGBwCjqathO8YTSG9PeaRuUM35R
c2+PY8F+BbcyMV9U4+NF/PYP5MUhJU+1ezwDvr5AILQYej5H5Txc7jZy/veKCPGe
gh7ROcJEfz9OYvO1hz1EJZShaD5jQorWmhNwUV+9pgrafD/x41jnyYYU27oiWCZY
A/E1viYSkMVgPmVxWV/Jy1bdgYXV2w3kCHEDLFMYudXTQRMYX6sgm304g/7VZk4A
k6hKcKfbB9s95fff29LDeKFrSkV/7RbI+ukRtahmiaQQ9nRxRFV+t7GzQqVounw1
O8fR9d5I387DavFAn5Rl/jM7//1FenGFtzF+Wvh9If2aed4Wcv1eG+5oOcHMNuxY
8mA7sFh06G+8Y/kskHBqExfmxQNKpM8h54SeNzapvoPCIN6/q/S+meclam4yzKlc
TUNWrx3dbsykFhsfvcRPjy+Z/uVtIuiT++I7mvLIjlcDhJB0dMy901U3GxKCi//m
TY8Bbn0FO+gKeFRLD3SHr93dMKudOoEZr6ITXsZnjnYBEmQnPcKcEV+wdKKHRmES
7HfH2BfJu2ZEQN7Z3h7eiJv3p7V2vikwfdpWWaxA36UVCjguyMPJqbseuIlD2KTw
CX80lhBA0vVhXA3eB/fh6NRbP3RJoxPpqdoOc92Vr9QOg1oyBKzA07tUCphEnekk
yFwawr3rKDubd5fK+oHK8wy7GDBer4uuqSrABeEtjSRXKm2TDVAMghlMcvWCtCXy
FIT1Hc7lyozERV0gJvLSz/8Hb5+bpjsLm+P72Mh88kfW5qOGMZfBbkR8RP38tfu/
Gq1knS6FfhBKpdfnrWWU92EK3ZISy1UKTMrqNiB1o0dtN1EZpI08AGQ7WGd3cM1b
2IRda3OFEUswllqur+kWLrzuidPsIPRhi+kK78g27wNvUI3xLO1Ma9YOf5b82X0M
35s5gzEdEeNFYZlNsjKSFb0cnOGcs+6nZrewM7Nu2lhLU2pE3sFbpetAW5P+ZlFj
JVfS7JxxX5QopuLd4b3UY38sxu6YQmebQSMEWRTlOHFFTMok/gkMxOdaCXOgatQU
HVD5bFxu/80lCkeLk78dj3HaajAyBKJ6ABkMiiN/zw72w8Yd9O4syldTp6TjlLI8
UaiDV9S+LbzKQJDDc7xwrvI6EeOOO14Ue9gh5iFCi+OCco/eSAm1Y0cEVIbDw+J2
OJv3x32/FHK+ctx/0z82Ok2R2YuTXlJw/QHVSwz7AaxTwQjlP/SNk7NUpYcZq9Uh
2cspYmW9VkdWt8YXzMYrluCH/Q/4nGmFRo/pE7x4wEtPzZAK7C4Z5O6vNB3rc+7k
Kxr+Bd1+1KiVhHTGMlN1Vy1LmshHm6pUl2y9Jdr0SiT/FBF1V33NwGUeJYL6flcz
Gw7gI8o4BSyXF1FEDP/wkJmXEiNn2gQL6RiYLQGyD33CN6DyO9xDJ10A91sZwEXQ
5GiqEdLp3P5fGp9KdUoHG35kjUaz/XlmsbrCZGhjs4YCCCrOQ35iHAaXNaVU7sZs
/3hMrBcNAwnC6Unq6P62YwZwX8ASEZkemgMSNAceMUv4NHAUnducoP50RPMgcDFd
zoKVjitwlilryznRlMqZTyYtKfVqwAhnzFUYrO0MPU6g/3T+HL31vC5KXiX26N+j
VEQ5EhmM5vmQxzRpDVpoEZoyixprk3SKvO38QsVBzeFtIITIVP2QlCybFKcPIGfp
BCm4nbA6CZK1jGTi2Xtm2QZqLt/mhb/kWADwt8wgYk2I3uDksxeDI8AvWZKQDfI4
dK2oz/27dVY86GEQS/TM6jmyVKBTmCcVn3p0PgO4O4+/ZS5hVdW9k9uQsnouTDxk
eWGapJjF1rcEQP9bmNQ38Ir4+VcsUYeV3q4y2ULeDeGx3V1q80pOvN6AGKqvzwHC
PXIlRTz4gUhfEdbB8Q9zGDGYehFNdVUnswI4U697VIEpvP2QL24EqmAExmnRPLhL
xOuKH5Aaz1vbuEjlvqjd14+07nhsBPM9ff5DbHpXcdtEa/M46jESNehJ3GlOJFto
m6ARqFWDFhrLfbEAHxdFqj6SDMAQ39VF63XZbGtl6DVWv5IEtL3aBHPrbFc6xqVh
H/zEKXWQGC1fG6I3NeAw5MES9SCZ6b9HlaOZJnQenBdNvWDEzn2wMmBVn1N+rClB
YRQZB7Ix79TCUnThQ2ySTRTEy9u0uoYhn4rtjLNNG5Bx3xY3dGr6q6ft9/46kuBB
OhczZSGxRuRhJN06IFa+Immx5R1b9pi5889ecVT36KjPKWSxETviJwxjFstKr+MJ
zWRXYBoXLCUBssgDWnlz3vMlISGcT5WRk1AnVth5svng8qpEJUgBnw+BrK/VxGvn
y1uIgxXhNTSeRSeU0kSmdlqiMrW/sopC4N3ldsc3ZrvDLnjbj3OvcdypLLOnsd+y
EWH2FzxmSBrGgvDWZA9r0S7x2O71CXhxXzqomUZIm48iTK3pvAgY/Q6AyLcMcpKj
k85Tc/ipvDyfIgcrXoQipi/lOus3CxQTkZ9E2w/2rYXfUnpRShMEgLQn1YPSlaam
2A15L+ZJgEm16bvgetlEg+fWgEwkCgG2cX38Ok6x3wFk5ejPU0OHikIdxQLI9Jr9
hr+K75GpB93tr0V/YyVdtuWu1QhwyHfaqhKOWvShTkJIftjPQGdm9dO8mxf2rhCl
zqDyJ7e1K5+dusdJcOS83JkogOEh6MXvBzWyGyA0NIUIlNBDo1v7GcPnYB+0Zl/p
VhCBb3yRH3SrTMsnoIEBLSISBan9XndmhZ2xyug7RaBseKECN0ReMzhUY8lg+hDd
D2cLou6/aKy7qQSnmeyGwo2RGe8xPe6CZC1r8BWDJ4eSPb/t95xGQ6a+xoIRUOyC
DgfvjV+s4qnCk7pXioqdKoI0NkKHC9RFCJXP10mlwSqiPTs+kBL+qOY2j+cj5Yv1
YFE2BOdIkTZGjV6wwa2Tilcz8N/im0qMMs24OtHuv59owtcVkPMC4M2TowgnRv8H
dczfQw2SrmggK1e2uqd9hcfrZTaIurqlWVPRRTI+kkyGI2OHrsT4jjbYFDXJYanW
TDrKSo9vRWUxLY91qnD0KpJDdkFPtT1GZWhorDA8fpY/GXB97WzLGBI3D2UGsMvx
Cgw0M521b/sLPu8HjDke5CTquBKviK9PS0zOIIND5ChmtwN8MNZuotHeReWEBi5t
xMvVy5y8Xgm+2AZKit/XKn16WEAI+9im0YMyhawZlh7POAgRuMFA2haqilsgrf4c
BIbcrWfA4xrE7wAOB7nQW7uNgpu2tRg3noRMwaz9EXVUlBfCXEF89EH1lkaRUUzP
k0Fn/WsIrBQSfnDEix4nfjMolVCzErbh1pYnLq1xe+BQWRgJjWR7uryNocx79gf0
Trtb6RtFB/vpQ7ZbjjoRPPFMhgV45UITnVywjT6BVqS/Ur++HdlZ/hb/PM1S27UP
uV4tRMX7iL7N/BG8fDVwelrzWpYSYtsvSuUFQVaUDw+Ypet69bZ7fRErk9t4uN1e
EDPYbxJC/asAr9EghxA3c5+CrPTzUWqLvhgH4BM9TKEMNoI5DcxbMkMIk5YmffPo
1qKAZ+K+HgPB+Ry7mHnoGlyKiL/AvntA/CIX7Rg4mlxak6UAH9ZoD+tZIxaY0/gZ
3UWEUKwQNn+EE2M7OLxHsW7UKti/VGAOqgacIUI27WtnxJq2o7QHJdF2Mvlwy75T
3VkVlfve5aELCROOQv5go+3EgIKR9H3D5uldbTY+C117FDKEhlVwB14oKE/L0EYF
zeVRfA8htgTItgRKCmjnkJpd99WJaJ77nmXTDldEQajpuMyLjo/UCT2TMCBNM7o0
FD9x3GLyjP9WY1VJU5zh2sdv203YOube3jcFsiXQl7EiSbHZy7AZObkd5haqbEPJ
X5AJvy7e+NRithAmmBOFksQDbKHLMeSExO4/SLM+WlD6lfKZXm5YGSTeCXyne02E
OJG+wL+GSUx/wmXV83QyxlXVJ1f9/BSvNNU8AYng971MeY1Us5c2PFb0rGLrSCVv
cmVPDtHQrppheXFQ5fONO9tRPox00dLJ8jhWHbGXPgxoPkjFnAOZROZDpAQn24/4
jT57hbIGjjI7+OZulBVXAJzt8VwfRQLEi0LzziHXhS2fwlykH6pZWjAtaMZ2A5rJ
0RYlaoVGC+qOKncans4omcXqIyUEWXjzPXn2JysBHGdnpXYgt/uS9Ww0b1FHuVPS
LvxZOibPApGc35spVkrNeTjF0MOcs4PEEKfgEA70HT6xN+Lag/xRoTCnfaFSLOao
kI05VbTsNhPGnI+S06YO25isX9H/1IL3RZ2L3+dX2QtPy4vKNFYY4ov2Ngxag7qi
j1BWo4/rp0IHiFjyFAVzn/yIHfWAd+Iq2mWDGgBPTxLqnuVz+YsplSWqkoVMUc8J
jGaMj3GXY59sQ4RkWIe/MNKn9Kfq1HnZpRHAFuz2MtZ7TuT+9EfRacGVudVf+MAw
gVHGh0sFes4h0JehNDVtr/qFiVH/TR0hDHB53SN6P0vysnS6jb7FFLZFRrei3e9m
hv5WYV14iClmWCj3LzQfOAj6Xyx+22EHzb81v7jSbKy0PmcOIZNoqnJgCkHrNO2y
zuoyGbMnpSUJzp+wekqZ5mfMXNuewQm6d8i3suTdxpQBBWle279R5+Mjhu288AlG
OwXvWJSN0ZkCAuf65wK2c6jPP35qKKPVSsCy7zLhcyhzL/wfSMNzCmU4d609lC9L
WtJ23tnhkpueivaEEuGbXEZ0bS00DF5wynbouqilwflm5+iqzsEpkKjMI8xwm2J/
RZqyoFYIss9mWJmSoM8e5/0BwzPLDluEMbWWsZFdGCWYL0Rpxa7skwgqspOvL4zp
qNPu84oRyzinxwPuSLkyzxgWq0J7uE8DsRAiS8gAURVByWWm4MEXcL2UqskfS6t0
Jv4ANhNPpQ5fwoWdj/1bLRYXQzS4YOH/iKii/R8BzYHiwuO0qwnFfIaRfFjoJTpD
dDxp295G56UuMAKtXk3wilGbfThtQsJoT8RAHoGx7xwRpv5AjK10wL8WSDlCfaem
+7pnypv3iR8Yzv6EI6zGb0OmFWI0Uzw/fPuTHL+TXzpZa/fU66Fq+SxHWN9BVLXY
D5EJbAEcN+pxRwSsdswL+lxSj7zURbmP0okpxHxUlCsD24xqo2pa8NZO9L8ndnf7
t/3wV8z/KOy4v59miZ/oHu5rv6MJYLA/K4s57YkB1r90IXZ0PCrJXPQ4eVj4wFIM
2CmlZga+DjQLwL09o+DXAUut2qeA9hHPp1pzZBwBLs5HIHv7iZ3990T0lmKZK1nY
YL9nmwHQKPxovRXCWgREEGeLx2E5oGeQgEAbNkaMa1m4u3GtumLWJK59NuXERzHp
Zvp8dacqq7+tE8qldhRZNVTX+7C4SsEK41SVlsolyGWvEv89HbsN54O4rMImO9lg
ZZ8BXWR8vh+RWj0qMfpyB3fBCgrH2FcuFHWBFMr/Ngki4PT7TLXVDrQ4FabwoazT
N8aRPm3CeumAQF5TyW6p3k8djb7MNnW+o2Vdf6MNAtWTA06sFqqt4UZhkyeEk9lj
sw4TgZAJzvJS4Xfdp5iGYLoTdCucnlLXibDagkAdxNblsVwEgkSYrFpUOem2oZHQ
RWDSRGH3c0isxGi0N6u5qscllS8EQ7+BuZ0wP9o4bGxisXCIoCDR9X05PPtuGBFh
1EQOnTkDZqCaTltinXi0p7hEw1uAExd3H6iNAefpMghkOES8eQE9R/78Ys6IpFf9
bQWwX+djmckHb52O19gUq6Fi0Mh61p8AmlIt+GdhmB7Q9r2NTZg21GObIWeGyghw
rfv9UydsLUKVH6U01zzEpNxpHZT5VGbeJLl81ktJfbDYT9vspnrSMCtFFaOhm3WN
piT7PGYSWovj1V90i4WXixtZMrUH5/oF981lpv02LeF96NGdbf642yXXnjvZQRCJ
1b2n8q4j+8jxdOhJWAoDElQirba6Gm9aqAJJxgZjpIOUTzz3MHzyZKcTa73Li7VO
vt2zqqeetgRPY4lx58M0vZUbkatoHZFYlX8T6o6dB/r6lHagRI7HQuPJISyWyW2s
QdKTRNUYTBQE/RvaBlTEd06nCvsirrz+ZiRxO02XVhU07Hw06hZ5Hv5qsY7B7mEp
NgWbdMZFYDtj+lqmWyZUqLzfsSLAmRsKnaX6hJ6kVhlH0hUiNUf716bhJzJY8+hI
D7Bsuzk22WQtrgvIhoxrOoGEvq62fwz+XhL4Q8Ef/7u4GIXynvD0hhHh96jJA/8N
BTVU2miRfOaquYs46ctNwGLpezh6He/b9YgktS7CzZtf6g/owPxD0GAtpbFALtE7
xmbgVgdwUb82C7twCrOOjJ7O0Xrrk9YjvJUZDgIyBDJKiPiiIFLVJqhqDRLPpdOm
A+jmoiGLzn8ZsM2yh1lZIpSQ6h0wdZGlPXcydj3AnTnFflh7mncg0wNIODXCTHXN
vo9/JKThBNY03XTvcwx9DPlN/Hm6U2zmcq9LDXyIY7aWxnHZs0jM1QWNkQP7BsA5
JipiFZdsR3wOZfa8bVPlovywoMpVYoHp/qikukSO+uegY1lAKT65Dp9gZ8++M2JS
CDR2sVhbqoH/hdYcBmhYhZm6ho2qWXGF3x72fIEk7iSqBpR+qY0XdcLZTSIMsPu3
0oflsOuAL9XrF6XzN5wxvDuG9UGyPcYYo+dZYiy8QGDGzRGgQOGH2yN0PJtEWoEy
2x02A+vp4YUjLHSLw1Y5BIbOTmRBdKo0M7jwphFxJWcm68Iq1pLXzs72ccdpNz6y
oU9UZX/B4p868XEVHZro01m3SWG20YisTjdtj8xwpIzG/Uh5cPelLJ8CvCm9XcDG
6A8kvnATqKKKj+sWQUzRw0Ha9VILvjaf0E0h7d/zXoVFIjPEl/2AkKiiip/S8a7U
zBW/EFjYs9qB4KhLbmMgs6hIdPPaZ1tQcJe7j8cJzRRQJGhW/4ScYy40I8f6Xt4f
mraVB0DOMKD9e87S55tYU94hGXq4pjT21UymkHEuxx8LjO/aUHek9BayB8oX4umT
nmLSgtOBONbq6gcECT/w6fa6V4CW3utyFZZ2mmq+Ye3yphr7A0b2/fzOFCzeRwJb
Er+NCYBv5sHRukDbMQD/+YscOmzibefI09HwhbQLuKyGkwNqEBdaQNEIjfK0ME0h
48ut2Xm9lr1Oed6/FpL2B0o6WvyrEtJFG0MYmR15Y+BD/e991IRSJHMlGlLIqPZo
gv1H1Busf9aG/spkHHdVthkkvXpc806p/nfUinnsFHXbQQwjtoU1Fw4+7mNKfsK2
7+pjM1479sa6PqduCt2hDbLd7ZlVGXx0dN1O/EpHbuGXWvE+bJcreWT0fgHLgszE
yFrfYRolHLyLcq+Xhr31leMUYFztVBSo+4DcYknBiU6JTV2XCY/Afb9UwFOuOszC
JHfkzcMuVWHoSltQWWMVAfHwjlbX5Fet0iE6bpyoVhiQvS2zCvV7H3+11im/4MGm
XufkLlL/jnYx0pIo27BGRZ3Li99GnQ6BVfLx8TwyxM1aHXYwn1I218tcwmzl/xb3
I+N2MgG9q7NJ0o0b/W7Pmznrks8ZFWqKr0ncdKn5lzus0SS2RqsKhsbRLi0MhgHA
VStAo9MW7zMSoaH7E39s+rYUKtnrL4kUeBPVGgJh1Vjswq98p25N1Cxj+nEzLHpW
yVyF3gIdaNbkpS0A2OvnLmSklYXJkU2PFtHx5MH+KwiLgIUHeUeAz9rdJVE5EUbk
BuosxWzrPsd9pCBou1WyAiY0h/P/sPNeg64dISqPWy0CMrBGDA4JSsT/Ud+bfeBC
VrQCCAfklGoPS/dh3f/QHVdcAlFpNjmYorMGaefpZIEJtfIbxW7l168ZOh/ZdF3N
uqSrQZLdj+EEHM72M3dOOyH6+C++c0DUtFi32GtdVf0+wyLsaoSw45l2ciC674dh
5lHvEtMIlzMG18VUWUNtHD8LhWXMmVzJRwhD+pQ6Gtf0LzotK05HsXMog5jTQQga
wFquHesiY6upZQ+plpA19U7MMB0atCR7L84M6xKN5nTlLEjQBplWMzrgIWztpeU6
a78w0Nf9oJ1ibI6CDLDT9nlEM1Vg6shDV8huUJYzW9guHDmXfEvCWrn86jS+TWpl
U5ifTlQkaDpKgECJuAdF88xkpOm/7OoOm5ks/Dyjs6mzkdbFwxdOrz3tatGwd2ic
T+gdUFQGygD9j6ovISOcE1Qx4aArKbdeCN9P32v0LNaMiETA+3zPb5c7mv81t/Dl
zQNmoQtnBXXGj394abK3leOSPP92AqXpW0b78OuwtfqsdlvK55cMzTcgZaD4XrtP
4OygoyXEFoDXI4oqt5I6IGIRUsyoXww+1pqr6XXzNWqh6nYLUMy2rBKsvtmC9HMs
xju8aZ+zyZ/mTAmZ4yEcH1LwOVAax4OwJsnFuWC6jeq5rpKLmIzQrNnVz+kZ1/TU
UNff0NsZ1oJ19T9xWgbgo9LS6DSU5dq59WMKFAfwxRBKS7A7qUiVrGTlVln0wdM0
Q5HqUjmutMgcIX+jH1tLxI8EPPtLMKKlWi/QdTbhVsRK2aVmuZC1eFQkkmkKtl6B
6lN9Q/sKHVx/3UovoVoKe44MpUCcC6rUhsFmMrVqrphU347s1IgKjAFUySfO8FWj
fTb1esDBBQRTh1fI9OngdT1kyFaRvl+yeTNhoLTVw0iGj+sQfVrECb3nFj/m3e8A
p/uoEP9zDh1eezAd1sLlk7aWCU8Pe/hNukevngj4nE4+QsYA2Oum7jMoO9VMHgDu
XbYhNImEryfxQPfsrr7Nl9mkTMljvMmFb7m1+PG7gk/pEFNUEHVd+CXbPiGQ37GD
8eh78bM5wQRmhkN5GPpnYosYaPiR5TEDTTtKDT6SVuLb4YixxW/8kk518FH92Ded
6LTOA6CxZcn49d4T5Yz+8PpOLdkrIRx8P4zW/1FPvU8F2Om+y2vXp8X7+F5pbYm/
800QWwo5DcF5HKlom3QObOdoIsnIAB3DJNv/kXFC1ygvAIV7/dnbGObg2UhN/7hW
4nRmqxGDtgwYOJCr/mnOmSd9I5MFk3zOE9s0Zhmr4W7yB9lmCfyVG1HQ2sYcZLpQ
MZFZ/y5CDgrMC2iGasXVFglPkEAai/5ossB3xpmSRthqY7eK0VkuikAIm4vtnYRF
P3WwryNXFKiBCFJvAQRnr+/0JgcEiy3W9wweaTay22F2OW7AJVny1CWup8o4vebh
znlPiwNCjYjRteeZlKvit6qGqAbusEUUeUI+s2Q7kMS1Eb/aRxQvzjGKu+SxSDmn
Gh3ykZbiIanN80fFaf9WZI+FT6cO+IdQmOL9wgQDl3aWCGQd2/l2K7vmVkd03nDr
BMvNe9F5TrvXCrGRQ46ry6cZUV03mz51kjYq1PMmK4WBPUeodkolM39jtAvtxWRF
2He5d2V9Dk0cyjSGHzeOAt27IrRw189/STOBt+iWdGwCmpbkbhl24RNRJLOaK3F9
FZlqMvG009sbj1rjNFw2HDn2LKU0PdxQl5hmmJGtyBQHnxJtMdYUiaWvwLUiMEl+
sj+HEMYQpeiqrIbx4MGImTWcLjSAp5No100IyYUxpkVKAFVngZ5WXLE5CrI+eNfc
iiMipctfhGqPDCaNzh7ESsl1v08p9KviPqQLI7RQprv9fAgIOaEKv+K0koLeAsvc
00Q0QZA6ITOJlvwrrXElwQQZZ/CoOWi69/sIIRJA9y/i04lrVsnxhj2t1k76nLSl
sCayYLAkWk7+y4LNI/kqXwPDqong6SD+OiMkf9W/f9Kww00v5D3aR5WKoFomtcTj
SWDJs235i5dQlNLwTHo5fheuoJS++zLxUpQUxhR607loIXluC/PWlLXZcKgJDGiU
psJS5/8YwTVMSazxreu6h5aU6hLEuwGybiDq08WBbbVeZI/CIzueSGh85WapMyl5
xhhl17PdqnmHwpetJYi5+J/6xQBZivuOGKLIhOxxiGuXW+MXHyDq0HWLZkPayElT
eRjoeLfFFiw8UNDvqQIK7kBDwxScCcHTP0PVxOqzJEpHMCgzipH2jGuQ7Gqj9ubn
kMNmrS8/soDAWG2JGnWvNDUJaJXyLiMfNhYMiROeudtew1VJ3jyL22DpTdz3iYqb
cFuPzhVkx/GTS7wb2Cu718uhKLCNu1K+64ayFCSwJtXBiCr3gYcLYH4yiFJeOaFq
J8bHcJZgbPRbqVikcs+DYh0OOd5VBdUF22Y1tiIU635ZLi3i5jDvrd5Vg4WiPOrn
LEfhhl+UtT74Wtf9t7hzMmMztGzHM+6nPTQNUdV/cWvsZL92I7kG+g8HlLuQHw7b
6eTHJXXnZtJc6DX5QZeifVQMB5L3N1G1oaoOud/esfmRoaarJu6r3hD6aMTvJORH
s9EbNZsxU2zd4c7mIN2c/ym0HOYluKc2LGOhcQapxR5qCJRwPGsvSvg4nrEr67zx
SX+EJY1iJv691nsR5ADwqz9bJkyTRt+t6+xOzqPJ9v08hUZNUrBT4oHMH4kZQQf+
TgZ+mBlbzT8M1kmrul4e8TlkAdN5kRzhuYq8G155qd+u1cxshnmh+vWMwHAIxIuJ
ihLdqKchjH7WvAvVcoRhLETPzM2TaR5CV8FglvD6Aw76wQBWplY+dsZa8j4xX9Jd
zcU63k1eA/EHU9eZ/aY9JCOVg1rgkpQx90ODwk4cj9OcR+y8AsW/Wurc/dAVu/Z8
zUzSgJd/1Id8kOnGddXgy8RAHxP0IF8cNGWmta0YFFnqR9HPQBARSfA8dZH01nJl
572+QTe3yQNfaQ5KGmsF1NFDvxZ3o62i94cRcOXCC8G9TycruesrWksILstVFxUa
u1Zmigf+KUaZz+25uTksRcjd+J4QQXJAOsT2ywCfE9iCREGn+yz1SgolXAX0zJj/
qU1tasFJtHIQh+vSM6sLAfH4RYD7fDjkegBPOZ7F7/IBKWXzwl9wnBJRGTDQjTdg
4yKYizBAeM4t5+mimRwn4ScrFFijK2rV5S4g7MO5LBuGc76HLPO07E/bd9oKJvwy
tDbv1TdXqupSvthLOr/W7QBmP9kl3UGP8wwGHGdNdp6lXzmJXDGIObqbrZmHqDSW
Ft0/idbNWBYWAyCCkHJGwedEx2IpzLXxW85eeCY8+4U6skdh2lg/9FG77/5iKUmu
Yd7eRBewxqGaWLC5wvY9KqDwyJfNIV25PeP9nrpSV8cJWct5ZM6mpkBXAn7QiTiP
iDI5+DYnY9Kh+RdI9iJ/hf423yB+LYj6MkoftAY/qBMNR38JnW2iq80WK0Uv5Esl
HdEoTkvxSn/yhp8Ej4cThhQq6/Ks5d7q0pqIsOSO8XCTYP43GP/S4pvsmFpjYllz
1whcgTiZHtJ57kHcPtXmwfODatUPRecyMBsB5oy8Cob5nteVup8bmASFIbSxsqxO
6uRQWRuOYhK/0KpxnvgNMoLcGwcSc8gW8joVM+XXJBsWGhUU/ZPvjU3CWDgyBXPj
+DHaQ8gBVvlDHpjde9bFhtzUYydyM21dj5r+lTdlTEK5QfG/8AP1WoCqtLdDnha6
9CObb/EFIdigSYdPG0pWr/8qsc+urdgEHEYE9Z9KzB04Y6E5W6YM6vohIDhIjfHg
IYl7ihPI6vUGaP6NuFHprsO6xycT6LSG9cHhF5J0qVXGDa/gydY2Ro1ZjH3EMZIK
YFitgQDliP3cSR2QbFUR8nRhNfT1E0fBAclUPmW4DGVUq5aetQVpkkBjKE6DVt18
8pNSstN8eSeLRobGoVqwy/qKQrWz3MW9s0kf4+0TghWJuBmLqFTNsNdHqOwHNaPa
SftJbUqGy1YW/3ThFIgvWswiE+AyAhGWIk3rkGPmCiPZ/+OrUVAYX+XGP4C9vLDc
s9qHIEZfazIsSUoEFUhvfj7PB8ZaxlKwRy0Yh7Hf0/1Cf8tTwm9KC1/oPpPGZl43
0Kcd5Lmsgc0bG8A6UIXeBwcQFeUP0+Fx3iZCdw/pzVtaOST9vmlaRYHgaMT2XSJo
lSWKMyg8WuDIPdeG9v3B5BxHFH4K88nq4EjYORNgZUdKbOXFlg7WSRHrc2V2f6ka
mcRqaeSUW4pC+QqS0F0MlAwwtex9RByV4nlLRJeR0WBFGNX6kPFKIYYgFkk7PKAQ
tiZB2hAm9AIsEjtxRroqklOcTzwLyT5uk2X2006EXnB1xYf1FeKovpdJ1Oopr/Ta
3CLyCAXer7LDKDGy9iS+qOV9lozKSQnLPhp2p6YdGyqlS7x/IxOCWshTFkt5dlBE
utT85L9STaG9zEHPVlg7sXvh3bvNcpeWXVbknCZv7aaSn1AKfX0y2nQjX87wtNGg
4dNqJuiWcLtYTQQZgVb/m+1ocl5LC3gIOk+Nmnij0qJy59zEVK65bgnqY2+sQFeL
hAAOKUzIou0rHsRMI2CVP/KsMwYhO+xrFME0abcHZIzH6vHykTj+2nVph98kctUg
yAO76Vv4e63XFtbMzt8ghbgE8/NntZPh0ykUKltqjm9+0UuF/cwsiixY5bbjuv5D
br4jAMW/6Xg9vBwAA5Bzlc+TG4CSAM2LpvUjp7czdNPcMpt+wzhpWHgSEVVqElaX
B+Rs7O9Bvz1v3g1ajNIoQTiIEzlSJH2o5oDn4zz4NTfNiLT0kOYWQcJ+A0vDKMbP
ZQQKToMjx9t5+JfCOfZNixN6jTKTB6L5O4B8lk1IwzoVlbn7WtK/DLLHaDu27CKH
y49VJd8+dlARH6y7tzh5+lvy3ha1j1BQjFKbNbMFLWQpZu0j4MyRus4G6K2+rOZA
MgmEnfx/v+tVFKmzZZBfN4bfJSEBUfyPWHx027cXR3WYJaKWO1TB0QHtkACqdrkn
aL5S2ggAABJ+Tz7tFAgVwBDwxu78FrPOd201kEi4IT/OXt/sW3D3M2zoc0xIAP+H
Of7V1x34EzEtEqtOr1wJI7bmuDZQtutKZ83ankkkRi7M5MZC7/X88+0qqwbq8rIj
Y13LjUGm1O8B3GdRPSmYegd7jbxlJ3HSLAbgIaIhYdUYfHHH1YZJGeDv1cB/w3py
2RVwsKgqayTWhgxd7EbPuAWCWdzY5dbQT3t8BhkvS4uq6LQGTU/qME5Utg2EyKM3
xtcoLD5E49sdGxwZ5zvj3yo4uBFtH9E+fik23vE/isinq5ESQuzHO3LtUOQTaHsX
cW1m49Y8fQfxnGZYjHcq2P7tGyNa9rlNckpN5ojRUBgLiBy/4Eb7Bt102JGx4lok
YE+H6Jga+4xq5o9foz+IHY4RGY+nUBx9Djx+Zgzv0wmuOr2zTDgfIbhmp4il9F51
QhRZAMyMR/+0EzujblIRjq1/akzTE4kEiyhr75RtsuHhsXq/LNI3Ld/mrHP2DWUD
BMDWlRmn3oZXRBMH2EdF5HHtRsDFcC5Rj4BI6NuqA6MyKom/7Qezp9BI2MemkukD
1kl1Of2hzZpWuONp3YJL/b8KLknMhrR+u9Wy+B4Z+NdLu/aMLDzIqLTMmIsk+d1B
fGXi/rYT8pbt/0WTJ2kISXxoStwz4aQ5duJB3LcqvYj3PlLhtY3dAMwgd0BSzqmU
JsZO8mioMBYCOzHRzfkH6h8GyYsMYw6mELoevIkOG4fESUuxA1p9vZaQ7QovcLhD
ANyajNg9JIRp6mzceJfpnRKgUlD1qPi8mfmHFPQZz8SGyyW2DKiaIdUJrXBvRWlJ
fky/6dmMl57+Bh5TGfsCgrwpFYcMa/uctUdYfbBLTe+xYyahzI0kU7iCJT74sV/k
tKAWr+dKeX0n7XhxPi89EUGfJpgnNVVRDie0mISqI6D7qZCxjC7QPtmyY/OxWERE
1EjqkL73SwiiyKKecpR7OkuhOs7oy4YSv1DmbHBcMV615HjQUt4m1Bo/QVhDuOXw
4NjgrF9OG76G9kBSvLLwbVe+Ka3Wab3jQmb1w2XoLqPt02dmVRmJ6U7hexc8hTko
oUkCq6bTLL2ydYluOdSaNv+ze9pJJ7CFiZoG3612RbWQgcUFFq0icBAvfcBzC8YA
AQ95buBYtHG5T7pZxaYqxnzO3WzrKMGIbslR36ehWeeaLONlubtWuAtY0uP0SBqx
vyKm5oW9fJBJuzBfeg9cHUen4z9jDecTa/IaulQpW3lgpTkqjBhMqBsu2C4ybZgY
LggZWjEVp8+JX58FgXszCVQ+Q9Fx2iYxNIkuBu4sq1FYCGV/tJnZ7QfXQ6Fx8J7z
GugjhlNqah96Er1m6Cr4U6j5kx1jts8e8kss845gwtpvfG2TOTtQNsquf4g4NpGu
gVKHvl3b59vM+yd7hh7tKGGTnEH74KGfxjM+yKAxK152wdroMcqjzjcUHculMdJr
YafrTYHXXx4In2e3epa+zmAZ1On4o7gwSTB/HW0KH2/9tz0ujBIrnbAibuytu+Fs
ZvuQo/gswcBrMw+vh5SqP6Obd8omOhx/xGYDTCjt6Twu8kJM+riYche5dU1gFpht
vWvXcp4Pf8M/2BO1CIQ2GxSPWeGZoevSEfuugF+rWpAAg5Ibkid4gFU9cFMRUvoh
192y/s0UXsmy+cCT1wFXk3kf5wkpAuvGL1INow3XS4tj6Zyf6f8mawLvuYRTADmM
1oPo+M7WW+eMD/ZBIEyzXhLHwea851tIwY6axVr07/8A2SIvXaxDO+zHglec6a7y
zoDqbWE5fzbN7Kmo4DKSrd9aihME1AzyEBHdLfis7tdA4AEQCMrzg+txnbbHD7Ns
dH+nX5tw0rRjyje6C/v3pW4btXRGvnzj03YUV3Tw5aUjozmQsUBV/9Oexhvj4Kpw
F4ubd2d8rKFXCYHTlvkRMw4n4kwMvZWatV3aIVV4QX7SjpLAdgWa9kR6upwJ6U09
cnyla6BRDJGmRoxvULWgCZtPIuW80dAm1RipUcbwyy6VAOJj7DIBIKnQ20kq2xLA
vbQTB5NpyWv7ElZv0tTD1GF9CW7ffRgTEvuYhBHgzACUFZIZMuAVWB4UBNnyvlHU
Nx0z1lQrRTAAW7BZKDHUf2y2Bakl7SO7tic9M1UUGcqFES/SV/mu03uVGpbUyHbR
ONVNNtdpkLrlsH3mHqnIfakcOB7Wh8elb6Da3oAgv5flI1R/RbnI16WaNhLnIRsZ
JDLoaC3pPqYE1Ir2lKp2sp0GpJX+fHa2NJUkmNfWWILWvnyX/6n/WaP31TUrgjxn
mKVkdW9gTzIlaA5NudrssMZ2EsmqxJqKPBUAm9M1r2U/ITMLrgHwBmVe6k6Sskm8
2CooasAOzEVbS4IptK4PdL49/wUbkzS28X2jqpSZsy7lHYCcN4BdRdnlDxXuKbTw
3V34RfUelv+NwUOLT2PKfDJ8I7SDVn0Gf9FV9B9+l8oCFEK7P+/Fkek5gSqNKaEP
3Km3fcjquo8drWbht0cAVexIzWKFictplimJoi57H3Bw9nEwg7iIMEMMH2GDHN7N
tjTKM2wWWe8aaFjbAnpyb9AtfK+Z67u1Hew3kqc2emhtFC84HrjCsFLdoptVNQeP
VcAwGlKRyLoAFSO+xW5lO6rDqcc1q+1dUzUIWZjmbvt95CDh9buYaQRW6tOjndLR
xIPmo7d3tbioPIXqOroNyYmB7Kum+SMwr9FMSW97TrhJqOyuSEi6DmCqtwJnH81f
u8r9w08hCIQZgWOGPP08x9alFAtrfAP/uthyqL6Oup7Zjlzlr9wmmhIF+b2eMtLX
3QbGIumPY61ssciN6zvH+eb8ELgb0qd/x6K28tNClVp4HxqYY+K5sldB+snPu6uy
9e+hAdnwsm/K6lhNbMQ90TDZrnFkd/gKtGnbePqSynGLyXripO/G9AlGCe9YvYSn
ZYEgyytkH215GYHiEuTDaL2uhtuOeIN45s3ElY0pfhUnQwWPYSPA43E0Bx151TjK
56HZ1Jn+bZ1zFg1rhLBqPlzdJla7uYCXdPhupRR6UGrm0rPoNvdSWpGJ8l8QRKqj
9Rossw4sqmdnUaKuc0JfxGdQOHem7kGjPP/u4TnehDSd1vY2+SuopDmMShsxua+7
W88bKLEetwTX9cB+x/bcikZPtmUug6AzMzbaIjnf1ctwdP3PkMxb/G7txlAKrUoH
M5RYelaOI4o/BHUblEbGev5NxVDs4PpH2zMpq+JOsXygb5fygFOm/zzS44QfIl6I
ucZd6VCVkOL+A4BttlhVXKQjEzMEZciJGCpAa+JGS2lmFSOSQcgdedNs/NyitL2O
AqqvPVrtGOx0IYYYUmuM7TrHd+rbArDyUGYnv5ywyJg0ro5qqY5koCgtfSLueCAJ
G4DCDv8b2kfGoqwcz4RLJXirJ0NUMy2/GW+ucBcvuDiqrVC9msvXSGutzJGWlN6F
6Fgexs8s+JbPnA4/jzV/KXpPyqKULHr3oeIDHwqs0QI1Kk3xLkecdbo4QnnEe/Y3
bfASJaiDhLDw2JNroSmeJS8evLVzJONIVu9hSRtr3UNNBCfC5FdWUd366DuRGW/V
6fVjUERoQnX4MMYwEoaqEqakRrPzQ2dAoboTqm1mWrT0EyXKzU8SAkBB93cM4X/N
FW6yf0KStQETw4wCW25v/BwNXdBEUZXMefF/y3MHV5SU5IbqleWsUCd5RmvMP5PH
2Jpu3y+ZIIe7jg9P/jv/8/Fs+ratSUTK7j72nkYQoPllLQ1vbsgaLmz52mDvZr6j
i4ETQWpT/yCBh+ZeQGzgWTdmQpOF7mJU8wrVG7UG2uv2J2cjnndcDWI8LKAW6f3E
nku/riXjOEnzEzXHsApPBuO++eU8APqXbzZhjKnQZ+Tl8yzNtMpAZMGSSxTyhLLu
SU7P7m/powXtYIhpSvDjVOezrIP4pPdLCl+6urFXj0M9QEXlxbDnFJ55gtTdLzHD
iohMjybn4MJPLx4dJCFOHjtNaWmy66kLvZx8mKlbZ6YESGNcXsNIhy6eOK95AYWS
wD0ZZFbHo9kSoMxoOy5jtxRckqX8HBamkBnw8+GVaNDwyeWGo/G4ODGpUTL5PGgr
SkPqT9o9cumuQc8KV7UdrNlEeTxAwXgAizXaNtNNpw7piP9zl3Y0Pk0+pBV92QQ2
xijyJLU5/8ja18VMGwGbKCdyXCIE6K7dFxmNU2ikdgsnB6fxIbZIr0WXsEQaXIri
1kHPD98YZMtwJgoYGW2JgC7JgNkNHUZ1qrQaKfIw4Jq2c88QGXZlh97G/+h8t90v
MNdF9ic8E3dXkrlYfIjKWSBKpFBMbtE7zv08n5B7Dgpcrq9PbGJq7rL+g8wh/FLe
mxFrDS/A2wO0e3ahsGiI+hYgQun63xxnAAix3DgLIfOexer+oImdY7J+z296h6n+
S2ojvc71pNCuroZQXpXF0UbkaupsEuROUMx/9k3dLNBd8u+FkROQgkpYle1I2jr9
cHrW1VOqHgZPSIf1eTrY5Q9dfYAXS1paDX+O618Y/YymbMX/df7UD4YugrVuWj3P
b9fxUKKeCy7DJfonn5oMP3M6SCZQpjXn7Sk4hqbuBPf3xc/+g19rO4a+m0ltoJzV
3ZDCTx34YqOG/rjEoU+NuOFva4X9WEakEgdmXABqD39JRPC1s2159csCo4aOjR27
BJG2aEglT3FEh2ywXH6qyTHfYyK8+udNiseRXA3PxzyfKb/Y58BW9+MD6SaiY8p7
67lmTbz6SGDIKq1KG5vQGD0vokfaAS78eVPSbr+Hx051g2HBwdr5Bc6fWAssLw/Z
GOTDHU6qFQtvQLtfAvywnX/xP5n2mACf6ibS8XLwt4BKzLP9oLs4bYxHZOnFydFk
l0TcsYTVsMOS9mGDnV9b/caa3h+bn/DmgY4VQLYvQ3vwQ7D4HYGnP6IW5Sql61+V
H2SR5+dWc6gz18is2G05QS1N0my9+0kYnB45hXO7LyLFf1Nh8AgpuMM6aD5OUbp7
fTSlS4sAaJBfxQKIQdptc+DUWprGYNPsnpFXfkkezn4o3HmBXNomZPujDIFAZZCr
W+ISIh5SjVE42FY0uaBpsSOLAMxhqINAA29R3HSFd2eAQpYquYprIPaCCliYOlJS
Gy0d/FR5eOThwiHTJCTR4b/Q/ZvBRieNPVVPKMPp14Wok/BbajCO90IhRL2JLJoV
ZHOC1wL/vYdhZ904QAeOH+TvAWKFSkRPzSMJiCjgLtWcJxApMk6XLJTi2hcPsHca
Pe2cNIO4w3xIogB9WjvL8Ee8ezeMY7AkjPIfvlVP8E+aKK5AnjKabv5A+yYvI1kk
KcIPqMqeIHu2bmLTPuNnJLspMaZ4vIvvudptpuWIajDxSKIP5iSE5p2/V15qiXaH
OsgnwOhbZG8LEGMh6N6Vail0StxkqxFVQTscveYJ06NTyIDdyZXfMQEXryu8yshf
sPy6Fa5OYY4H6jsKj13974QuHB/KYCP5Mj1b9tsols5m7evGG9icrqoOIllYm9u/
ELfHilrr+BMHH6dvyYJBBg6vmMOSs5ZMIjI2VUXEAoni0yiEeULpdSMr1Bd2Fzdn
MfnXofKNMcVKv9bpZc2MGvaEtyV6Qoeals4fh6zLJjdvCey38vsE8f3KEzG0aA2k
mPg/8zbMFCKkKrDbA4v06rknwaL0WOq2JROgqEPeA1K/R45LjJdu2Ft4aVsuuunK
rtDupu4E7dc8yioZ0JBp1CCw12V9c6hI1/sdxy/Tyjrf7rPF2QP2h8E/nRUCl49d
EWdUSUS8EbBN5ng3W4jRy18SrtMPJVM0dIjA5B4FsAnnOd+4OJWzn3SA+zgsGYOh
36rQ79jgPwmeDHWFjeOc4SdN5vOwGfqgM5v6VjXjHkhEJdBnyeJOGbcvikoCD4tR
JpDjcET/PVvT/eOH010Jy2vsVTaMeo39LgBwFPoXUFojjnb0y5iejWsv8dhy22OQ
kEcZ3UURcn6JA95je417pbB0SNYLpCBf/mEG8TCdjUTHYPV2T8kKALJ1Jlf7a96E
elNwWIVaEMsDq62aoKlZDHbQsZ0zG4fTm+QJIWiTrxOvYLRL3vXlqPecFXybL9M/
IOz+PXwVU83jDNyRooUlAoP+p1Z7fsy8b0sZGryYxLENnO4C4Fd1q18+EPWDxEj6
VcRTcmAymobNO+Afc2zkrRx3PTpb3lMQzVNGeO8rCFcI6Iwz/GRd8261Vf95OYKp
3xpSrthOzqSSRTct/9feEWsiZDohJggwYkNJqY5fTrvWSKaJLy8KUthubetze4ih
W6y355sJV9eakFFzIzRrhX6S+X8P22+P+8ohLClsxLa2ftxdMkgP4yWTl8uwHYpq
pnub9bI3T5PDAkmP2439YsiY2ndGzyUn43MqjYOqdd1vmCEVLZwJwlrYoWpry05S
wRT4xpmefmTpzq42JVPsQZM8nVWjr2QXRvMZxrWtzUuLg3z7291gM4PcOVxsb0qw
V3Dz9fk0WLzVNIr6R0QmH1QrfmgKvK6+u5kP0Ez/SXmU0vkQrmpVfAyUZDugFoVR
wuFhqKS+5gj9Ja7vw6xqXT9AjT+UJ5S3E7CaOPDpB/76LYMoxU8z6jo3Z8sfocVP
FGJE0LpuMHrpAD8EsYhOhGYqvHaU0eelL1g1pF4RPJkW9ZMIRrCiDq3UwK4ccvIJ
gRVwL9mB3/pTJT8Tvii0msmKpSwQVE6B42zUVQOYvNP/rSImKnh+Mxt0vTUHn6WX
udI9Z6oNuy9pRvo6OSm5/Hv/kUOAXf94W/Zpo2Wq/ntbuA9MVvnX+sT3f3ypLyp8
/d2CYp2idu+9HV25RfRjkNVCEG7IFll5+h3L3WrhYpFvJMn84ZcUtUB+VNtxRiB0
l89DMKgfLd7mxxRyOH4GiPC7pKMQDAl29AzB22jfItpw84YBIFee9ShO6hkU3rzp
ywE5mFQrr9a7w4lqtd5Gt4Fd5corS13IfCH6oJ8K/MByegGKrgdqFDyyRPZEKLsp
d2u5Y5D+4u7Du94IM08F48AMCXtm6stOdGUHBkL25MAd30BGt8qurgetKcsphpy4
qljeSeJKysFatnmm/4yhK1MNdC/sV1AwY4Hfw4e7S94KBICY2n70w811aR1ByzcI
JY60Nd48vo6FHxb8GeDQPDFjuK208pogxY50yZ5AXIC9ld5bHBAzNlEtmcjZzPut
LDShiLMXqkFQl2sw/CxmfEcerajw/7c89Pm8Ze5G1AZa8SDFB2Jd4rhKeF0hA/bJ
NZlwflXu0isDuFSAfq5y5c//NyYhKe7vrjTTrDl2OiAoA4ccMXB0zFL5kD4uVbGC
FWvL0iBs/m3UbEiUWjrPGpQlyQ8HzRHXNw7A7vRU5f4DZCedgM/F0ZeSP731ki1O
+2yJO3fulxirFqfhF/lBeDBHlUd9i+67pU6RmRDO67JuARohIF6SOX8NeRAjMeBV
b8ZnHlKsNVQKQps7qZHJB3NFG2B+xyDQ0/IIFX0dqYVZ1nm6+/n4yvBhSFROXA5Q
3uzPB2m4wbC7Q02AKM6nt/uj+TPhlIofjeyxolpVzRZhAr1Kl0ThxFIhZi1RwkOx
W0SlXQtLoaOYPButVHUY/6qAIRWiBGFTnyu0DL3/SzJEaPcRLdJvLge5IGJiIkmR
DVUQoomlpWyDqo8pqsCuLzIQWgmfuo3CLnJ3aeyi4OndOhGkvqAVdLFpfsX612Ae
gBYD/WB+Aozmbonl0CVh/KsRl1xPT8E8bEGSqCGqRqM09Y8sAB2vjSDUzKXZ4aXL
nVq0I4vGqsgZRaqjOeiQlvxRG8N40/b3tf3/+h1BxFaFrnro2M2pTuxiPoKIjxmv
z3GNk6ur+zmqBCWfobyqf8pOG0MITRgR/o50vMimPFBE5o1GuVGUFYE2FNBSMz2k
I7KvaT3T0nodBuk4gG3HpofP9OXLUc4m9CSeSv5yiwvwC25HmZkUMHVtkMgqNPOm
tu+5WCcFRsR7KDHtTqVqsQyuM0ymEPDAiZ6TUBQ5uo2VYR/8zfxfI9vxx2d4v/LE
1cW2kNh6uYT2Zm515k6+ngN4DL6Q2kCMoLwUfCUxe/LWjzJeFpjKccnIWiOOUILK
178KBCXRkkE9jUpalW0tgrg860ycnQrwjnaVbzlsHJMgcsMRsftp1agWcSfcTXLC
kM11hOqLIUBqM8TPxVxaHUxY62y/MY6PNE3QmPwkfyfIn0hyV/ji5o+sOcbn6MV0
9HwDd43oUP0gCffPcIeYHiaaN0LnAWI7lL1dWSmCdGtlF2tg9L7nBvm6CO/GkNB3
1pxFl64afy+8VZnCshTVLCFJF4mQZEV/KibP9jMK0BpTqV1r1e+iWZ8uhL7EpFuh
hRMRR+aWGqIlE0vqjVgzcorDwOYSXY2yCTgIK90XbSzanPUFhBj0aWgqgJAk+UjL
c65BgAmRVcCEw7gMDMTG+q12cIeU7i3BkSiCAb7pPDFzXCNdXsc//5hg/rMBgFNg
I/p7RR15dnOWqWwWX6x3v+WfIfBwAtJw2AZ4svXGLXtICojWet0/FSz/orofK9uz
2HqWEA1GNTDNypXB3uFLmcC1Jev8WCKto5DDGec9nDH1Rkuwb+QKtaWJlwKKhXnc
n6+AHfKD/5kugyWp/sbhdGlriHbzn/WUZ5fMyLlqzNtUzhQ0+u42+aQ4igSzEDsM
bFii1znTMDQbk6SWYvYYzGwEpTrg+ZRSa4qL+LW2qtuhJnSvyA1RUbKA7mVvQCrD
/C01pAQUzxO9x/y6Hp6tQbUEfTRT1uu0vpti+/4Yi2VCEOfwzIr/0WMnbfHoLvwB
wAYlDnU+9ETwxmXre39yj6QGxuqmv4BW0slFYlanQAW08tTvEU+ewcKkA6VzUXnv
9++6/d+qExdOXD2eO+Q2Idf20bkHCuCNY7/N3apA+jMxarPKmr/e0lk0JgTXjQ53
UBuAlhjtZgqIVjMvTT4+zr2lWNGPPXkWQvflFjtiXG61e7wNFa2vVGjc7nr/EIxM
OszzTAlIcLkf4Ltc+bPBd3Zka8y2X2oHSIowCzCvWLSF0zMVGKvqJK6ExyQojSSU
EhU+zBEWh55ulAxsgx2xaiYhn+oECDbOen4I+Rl5dDufTCXjygr5BO7BGFbEmB3p
kkc4B9thhjk44aL1AZGTmCSnVESH7/9Yu/NZjFJ5TOq14gGqb54Ad9SaB5HieRUn
EGZYqNEXc96NRudSWqL49VwZYz0LmesMpH5njB74mUcbIG2XlZjojexIobN7XYr4
2dHjOF1kyct2V5WYaEgauVzG6YB+Dvq2uZG2dG8uLOsE0YU7rxRRlSyzdK6nrYif
5E923Be+zd11t9sEt9PzLPiWS+QzqIMJLaMYp3PT2mXwVX5kzsI2Cnu89/AGBzXI
my7eeFwDT5J/CY6r048aQpmE3UgiKc6q1rEy/vx5zC46gOMZYv3hTlg5LcHvGYHB
KllEgMuxFF/0PlFFKuEs6xfQCiuIHzbKAgLsvsZsUdWc1miiu9UyV1yDHWvSsFHX
AqdMMfsDZTya1ytdhdY8qAYrAfBhsesHzM1VQcXL5COTtrwZPnK2XKDQHFmIciwo
1oRyMTElEc/6RXXUoyTP4Zbe0MVLDAAKnPLHvu5gLOau1AHBwLTf/QhMsi4GZ6QX
mG/9Zuc6JvtdG5exBe9ZBFqCqfmnttUeb0+QCEtuNoGxo1iJKpk8WC1/hflQK/7Y
19yZhYLS7bnTT9BjsQGMcz1dxZTR+QN9O5oyRzHwUIQ4Fu/DKnZQVlFBYdsDcIdk
+gUprKk7lMqlXMqeFVrsAyCRGYw9fQxpL6DC7HJwJZXsutZMnVr0fdmguFhe/6zQ
nya993Rcp2k8uHfk1/xrhcNGm5IMrlu6NBvEuSvvZsVG63Y3xOt4nf7y9rmSrhhd
9lwE2OxGIpPd3i2nu8VpDCTJWvwSmNcaztq4vhVpz81jX3QayC+Y0M6h4iM73NpT
jDc0Xoqnt85OfLU9MMN3DQCE6ssOA1QCDKz2H5gIP2bYqB+9nv5HPDPWCunOLDRe
XHMxH2kHXVtzRcNj64CeXuvuKxVhvmktAWOFL2u2zeQrEnnB4QA0nMbzXGRhoyWC
f/XAbffQepDtKdNAnWr5N2wf+KMWpSrU7ghu8u1shk3xLatrjydFWQTkjIHR9lPV
jcOyGmHfu6LdrKsT98sic9PuPZKIBPCsmAFbC+VRHu9ufZgcnvEjcuz89raSy9DZ
XqsDMMXBUGcg0x78TkubUd1TLrO5UhXYzEevhLqLU/3keuJgbyCkPU+k4JkYwLm5
/QEDxjijsJqw2ydfwrGXW2wz2gChs8Yfy3uTAi+U1BSH8kLkgmnv28LOoXwEWkob
zBfQKQqjWKSj/OEAGaF7ENzjRAZG618d52u1wDJ3Z+95gM3p5mmbjYIxl7krJb7B
1xSKJxR27l/9Si1T4ELcfV1e/rAZxmdI1hquugcOXAx+78boYZUAHpbXwslF5uTY
Q6shB7kRw965zrQaxOGqPeTwSJ8LNu5BZHnoH6OlxrmbihxXiSQFEtWOF1Qtu70r
jEDCxtWuoZ3xKvNViGdLc5NLdNo1sK6ZZ3NtQUxtfgicUgSGkeI3H0krky0IV5O9
hacPB9WQ5yihIZ8A8veQ6nSwOUvDW3i47EpGE73TMRuvEW/+KBJQ5Y6ojXocj4Tk
6LsJ4iOKpPlnufOW/OlWaS+whUPG63sQE/dnlm0C990B9SVVhRjrSeDstvIO2qCm
/7a4ldu7t/GemuStUS2tB7mgnAOfS+8ITRcGHFmNUiWAGuTLLbD/WwIUut6P8rw7
uUAYgFW589dKzGt/vmrK6A9XyCPx6kS1DBiDMmIhQHg+E4mEntomFsYuhXk+LhiT
OBACxkrkWhl3Ni1+deRbPSmEpgXVAL2n959keWSsMuP5lbxLbEyNEbQVKt7aHX74
OHtGfLtJL6ZlXUjJ66tps3wSRBFT2L9vHJO3MUzuAB9KBu01MxTzmm9kNKW8pGW0
ImvAVXy9QLB4SFfDx1k6JfYWs+YDbbXxD8w6s72qSFL5HQHisX09/xMNdT6xh0Rz
KLMz4u4SSw0LsSQFoIcMmW5Aeim/hK6H3g4BivUynUnzJWjSD1wHJ2T9vL/cBncK
cEkZrbsXm2TJ5DfRDRuwnqwNWe1nHm7kOse2qX1WBm74ctGc7dPowM2jjfQSkw+p
86T5yMU2TrjjsNBnTHWUgXBDj0NkETC/Tns9sSAds+nl1Eu9NvFgwydjXVoQjjs8
IVaJ+6bx0WDVAuCG/bXFnkQMW2NSC+qoOO52CuAkZ92NhXj0AEyAW6a66+PfHKHL
QaDqguFCrJF/qlSfPzLLdxY9eZjl0iC9jh7YEmyuXUY70qO9W8F+BO9CHmWXqPqr
8HvS7WlHRSp3X4vMpP+0OJUauzpFeOWz7x9EEcwi+r0i3hXBU6a7KUWk2ya3vnFC
WAnJZHjZpMJMrakA4bv+fKuc35KU+m0gyqh98oPngaldtghl+DV1OfcwpxlX6e1t
dC5sv4yP/5M5ebwAq913lDbHeJpGdkxH/27d0k1/EKP+ThRBtCIQOmqfk2jQCIv0
7GijH0JNGAgQiSRtUs+2OvJ+imEBPKG6zqm+YAwSfDJ6N9hWsmEgM+u4qkrC3IzB
GdLQ/t2cLIMIOWCynGmRRhKhJjCyfROjwmLhE1ZYTf4ymfcIc79+ZsPyOA10AM+2
d6MRjxVtBvulrvptp09UDuBP+miIAX9v2lQDV97GxQgslw9tj4b71JlxYZM/lUeL
hYiFoqv/La6/1c9YiSoqgdHF1QA18cKwaouNIjpMNlc1JC77rECLpQyBr+VJpzsE
/DZuna7mmHrBbTi61ChF8MRbXPLIpUq+yUzBqC2Pgxbbkjn0pwejkaoppjqrsv84
D3Wr5H9gOR9h1gMCMFSL017lpcFzbcMm2lZAQPVaoP1wNd4qGNpqBlsK4xsei0eg
YFAQ58fCt3khwJUfNvBwWGqyx8dNgva4mdq94z2fMEE8VrtD+c54Icy9dsrL+20/
Kv5bJj2Ob4FdvkmANzJYGpQdnZb8DXRJDqGIfPBLVQnfwU/VtnEsuMQ8BjcnR76p
zPBsfm//1rvNdRjo1E9Gy6wlvS6u1cYBujbV5+AxcogcTHmGhpDIZPeYDqTMjPXX
rnIFSp9qt/Ckgv4FAX4hxj/czbFfJi4NUAQ4k7ldetacKXtj7NOqo/z4r0/J7sIp
tPxCGiOpaO5RCmD6GrGQ/QaqcGfzuaJPhb+JpfFO5INHWV7brWK/rQI7skLHn03F
n1P0EPar5kAdyAvwqW5V0qbMxNXMW8OPWXW3jD5bQEcuycA39/kiSHG1y5VyIc3m
Mrh4WzslIggt3BhuQllC62EWjgSCPWSuJ5ugZdsERQBwPM2/FJoCp2BcL+bbG5On
rgMdM+VYW1tVvIDcE/r857nmjSjKurBVfWiWX6QkdbiqAfVvLkrDtmXdSlMopCat
OdK2TlqILI5IJGpFCsR09Htwbx0Ijx51I0eZeZTiS2G2Rd9ZR/kj/uGMZQuUeByb
0CpGamxlAvUIEjnNlTTSfiJvdscLcu4IsLxA2JmiTgJ/IDz8RYvuIlh37uAzN5pq
mKsV1iZQCP90yZmd3axrLrSEJTIXE7gCyGy/hwb+HoM2Vzk4158O/KQYuZAqHcv9
BJ+GRnsP2XnEMYAqP7rK3Fx2vB93EhB/1FVm/me9VpZtRVG/lOwm3qndXkO9+yNX
VSBMDg2/bmZ/1KQJpb903yqKGs7/xzDJcqDniXqXu2GSakM1VidZFo0IRZUVWyad
Ad4cRq5DhuqqFFAuM7rCQPMDB2bgA9rxV7IZw8L5Qet7nuLqDNxvXREnVm1Q9/GK
3g6bQsPrgK5jkYyEdJ8qFrtuvM76wtWzx4nAMVsyCs9qlwTpXlwkCxUA7NoawElx
1x5V41zbaRN9Fmxk96uf8w/Nptq4L37ZiurNvypWUqZ2YRX5vBox8sRO5D5Ql4WP
aDoAH7XF9TqbwELegkaY9q6ACbhYjBpdMNjcJJ21UK9bBgsq766+U2GYnjg8fErD
/1k5dLJ/Qs2pHCYRyjwgPOftsk2sfFirGs/By9VIbi3eLB5xMRXBxhrIsYNHaw+v
likpNtSLuoAmK0hFhsA+74ZhqIkBlp1gN9yR1LXEqYnhCKrsJeeNcUh5IPmYQCRF
WHGOpenTK1jTjtGlJxLugSg4+HUua8+1ef3+Z8N1hvjA+ZEZCzz3GOYkrOzcb2wk
asPUda4jox45ed6SNmh0nn0fgU9Cs0GaOcGCg/AgIiW1jatz+Lb1uKbKJI+YiUWq
S0so2a9sO1wAvNfqnUSOCLsoB3v8jBH1280v1K+FIpGUj9tPYOYXnBQA8uJ0IqWx
IHWu9TUJCf685ZhVvbny7RdTjtxrK/1j+Qy36+fCKAbZX4F+EbAhGo+llhA+YXut
J7a4XdR0oc4HDEIa0peGcHzLTrzGdCvD2R6wTrS9gp4FDnDm+5UShByQKgCyWvux
jz9hcPPi2Zpxrna4i9tD9jH8N/uGalji5g2BlMB3vsKzYlSz6797/Ax0V5J9qARz
s4pVOkl5nah2XKa8qCYQVKcOK7KBrzeWkrz10SNSBBppgCkDnE8hDtfNUAe4xjJ6
Z6VpfDQYi8dev6BWSonxItW5HCWKhw7VJm5tBAIg31roKAk6iIPtifrFsDlgqU6n
EqzQcp6znlT/dQDkFXXjsTGdI8SoxtXVMs2cRC/896wHTOnv4N8G0+qjiv8WGP4f
qiKH8wMYzdoYrnYE07RFtqOO2JZ7urO/tAgWrRvU1gzhunfidvZXn7q5e5AUcqXo
+q4w+SLTqDYZWPtjsBjNuK3VoG5J6fqdetrPY0KLAyUPBjnr1bbdi/FACqBcYQdS
7ZiEMf23vqrJpntyxzXr40SPMSCS0R4bbfajiUOlG37ws2ivdXzMd056jqEc/rFX
cMZ6aagfYhmfWZkluCOu5oj4n7T9LEyhzwTvh1zzzmCXqBVDyhI9duoS3nlricwj
bnbehv/6WPKYP7vcImFLxm7v7dvw0xP+Y53RcxS42kjzepXvU/HlfZqZGcm9CoiY
KX8Kg8Snj47BbfQjzEoK7vUUo9B7XOKtBtfK99ueukNNJiEln6Fk0f/rXugH0iiC
fZ+5aI0TgFuyhW1FN0J6LfHeNUtv37n6MFVPHkJgQuGCVKQJzDHKnVehFuLbxdk9
+aNDHGK8oQwugjpXmvOAPIWB2z/q+8Rk0vvmM3h4RrHT/ylR6RZ0Ewt0PUMGYl10
APDSize7eii2LnoNIr7n+9gJ5wVRkby7dqeBR5gVakxnn1epn+gso2OJGqFR27Xq
GAtjBLp1GCxgCUi4jF5uTzGsctY2EOv0wAa8qo9l6uNR9gDrfuTUSKhGhJevA/Go
ZWyd4/jhsuwLIZqt39Shhrx7t1jJ35abuwtrX/MLXZZdqZkVtJRHa5k7Y63qLQZ5
N152l8jb4celsQgTXZPJK74JaoK9YxyrtFdJQsQVm2ryPyQ64tGlTOd+eTUd7Tz3
fcPmdNzaJP+g2IHVkyyiSywWc2JkfC6QiP+DW7AMfGTRqxPycXvXZHgmn6M4KxBM
it5eOdQWbng3yyPhnrG/Iec7qu4KRNm4k+c/Kfx/mC/XXWHLFpQNg0/w4nj2/sz1
HeH0ARyladO+IH7PF5CYif9k3zV56bghApudwIJNuff008dycDjTsu0li3OalL5q
RNFhbftT3thbC8hOVVEdK3mw/sa3X0gOuUIEViSyN33zFBTiuPib5ClBcxm5QyQe
VKjzvvYWybdCYe+urPW7eqmQE+2VgisRrxL4CuMYc6AlM3hTYtqXQlLmzBCZaMLA
4AoIVps+yIBHA/Ubjyf5KN2/gQl1pSr7cmls9wA8TKS1VS/0L70XTRdPkdbb6b4r
5BuwbFDuzSJcUCSEWXV+rZnZnReaDWQdv2Xk2Do29XWaRGt8PpKI0Ws7nDpelX+e
079BGKAoTluYWBJFl6y17bA+h6sxtiOHiHJH6lEACWlGtbi+PawSxm9ZXxdgP5nb
PtZdRy5FGqd0C4S/u8BKzUWxwdh3HMHuvD7SvOiWHfyjuhXVqRPP3Y97uaEgcqz5
7xb7KKnpwFRBFvhaGgGIyc4ewz1CGt+PvgxY849D/l43ZwCXwl1THV8MhP9rDI5i
uGAwGUzJzQyOgHL21WjBqqbhjGvizRblAw5CbXvWbhlx+8jREopxp6V51sBOxB1M
GUU/Sg/HNnNRrR8NcDJdaYHRk3l3h0WtnNFNz2Fcb52Gmy+88g5Ds1/E7je1Zj5l
EO8OV+L8hLX4xG2Qr3zW7pLt63ajoMLoI+a4EvWCgYmTg2SMlmzU8FGYo45bZ+4T
q9bFr27M2rhJh3HNvYmjIpsYJndT5qsH/GUa/f2VSygG2DQ/5lWIbnMlKzKgi6l5
/6vSwSiJjJxWsVB/CCeGU932SJw6VzrVvM/dMmyjgD595ikrmVc2Qw/iaimtVq9w
Sz4qEsr6pok4Qqt5zx6CMBDTzVO7Zwmt6jtfiurn8IyQIkSjlLQpwmpatYlH2vw9
ulFCumqDJNNiDzemLC61MjzIvlvQ7rZpF/rEwQxk/O8WJJgY6jPdj3hls3psisB7
CU/pUwwKEGGzDgzySh/sQzR8OZv6E1yjFcN2tXf0bPLiYNei+Yp0LCoUrC00B8pj
UzQIspOiTdk9IjP2Ras0WFDU7apnuasw9MZ+N5kHaJLHTnYeqvnNoGdTyI+w6p+y
nbvXdqlrGQArQdndYdfoCpF+Jf24WGoVFpZNdYaBHMrWJlWJM6h27SvL515/HMIZ
NyB1OSw1gA1MqPBl+ndIVWvTex89NbG0Fxtcfu3n9FDTi7YJE/z4yJkMok3+DSz3
g9JQVXARf46ftLUW8nT8cmF8tHXAbPcgkYE4WN5R7qwAmVipchm/POrJ/3zDWRm2
tUuj++AZ6e7l+gCPHjGpLsA5Kyzs08x5v23UVyEkipKxkGjefEOxeK74UHOXXEF/
FOVmbjpRzXNi1bNWEGEYUxPiJhmAXgWYmJ09pd+hy6UgrERh+EFa1UFNnzaRWnP/
OVyPt4/Fvi4Aoro1WBG/IQucy+LGO9rYsauG7PRpTmXZwVlILaZBqcSLkp/bt6Fn
of+BcOlZxKffsVmFpuk+rI9E2OsaO/92gK6E+th/fw4hXELixBVN3ZcIJ7tu1hDJ
6YHmmapd47wA2oliw6Xr+z1KZgc6fA9p2KdCjaFoBsuZM3h40RTj9JC6Xq1ZabHO
D6UntFBTFb5Z8rPUErvkGxQNkNHpivWzXCweq2zwzEPW10/K05x1O2N3bZRp9G7t
pU6G17/tDtjkhhyRP8IrrVVa8pll3GL0oVkl+foAhmqkcmUQcsq5vlzzMljRxA0V
lg3R0KmWseB+SGhWpoENYm56O1ApPMcUSrGa2s6FRTgq2tYS+1ufcWRNzMGXuZ9z
juuMekHL7JfvCOl98oI9xxYV32hAKLEhWhB8eBpHUqPm2py6KLSmuHLkx2QMaKlt
RLAjShdL3G6oaQRmkxVAtTnFuZ7W+YFg4Ux6i6l5SZc=
`protect end_protected
