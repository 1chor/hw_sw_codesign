-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
G+/ocfr5WJynD9a5b7YntGmCZ6tWPBBaZnCjW0ofcrXmAABi9VL9nPxCjQjZS5wef0KiIcv3JR9b
Y95r/HdPnbSXO3Sjm1aJc9L6TYjBY4/dLDjHi+1AGmG0s7Rj3MMzMvQpbyYIe3Zwwdsk0bJSS1AU
HlcCej5e3OxnqhzbSSyr1b8SGPiksJWQgQPgEgSF8phaeA5jGkbDx2uVphp82GpflJEfPtubOnw7
4EQbAD+2lvkEApvh1UHrCQi3Co3BLcHiyDZYs3tDPW0iwDU32fy76YdXS+Xdj53FFmU2JlJqfjXK
tky85VA1il+5sc+h1xZE9E9mziAT1sXJfx4TzA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4544)
`protect data_block
2ZpOoww1e/iwYIV26+f3ooUEu3k4Z12xa9GRIcxwllGpM336jkB6SFbFBJJ6U/gYqg/18jH3+W8U
GocAld7qsCIf1G50d3Akj4ztOniCsi0W/SAh0DxFcvNscvp6LCah/uRaGnwN9LryippoLviIoeQy
q3rXeYxupqR6tQRc5g5wVsj88gomk6q/SV7RISgfzSrtueXj7T/DCjOnlzAc3roT49+EO3QwYr46
uZN/k34lTxlk4EuOKeNlhvOBw9LfNP9i61BV46ImR/8txXmjorN9jtSIMC+JAuxNxklwGTQflOfV
1EnF1eX0qfCFo2JXb1hvsz1IzmKG56Lc9B+DIG58iWFJNB0orn3OsVctJKcWKAxQRTyqBYljfom0
3iaMZZR3LK0+I5YFUknYK0VfVdlEWFRXZxXuftDK5vX5Yi+YMg49JUfXk6KsbMhGb2uywBGuYDIL
6yeyyKVw2l0ig6Vbrr1HmOFXu7IWjEJfRYCL0QL1nJP7xSnArIo+Nc7DpFFADYo3iklZwEgrxQiQ
Mrm26021jzATLQMkhScz5PEi7wkayYOZobKIVRKO+uD4axi2GjpurJbrtBRsCdmYgXJY2gboJEpL
nxLoZDGBijZ2YvfHN265bjjMVYk2Oa7/3DEdWoZrUClhq4dhrcsomWs90UGNkxPf4nJCVtHia9wY
kAMjHG6UiScm5Ek/bPxXZQimHy5BUv0UEWVs8A7+OpO2W16fwD0x1vKFI70qHa9Z4chtnhgOBkyF
6jrRjq6FFKjoqoozDCNsHurcQwRzL0QNCVIg0G+qG0GVCmBa2tjerjwz51HP5wybVfSl5J+Zr54x
cYHS44v9twtKpb+wMXSugXx+N59wF0Fbrka7ct0cT23UihHdi8to7Ns9RP2QL9HIQQM2zGpdrhDO
zW9klMfMEROH5SzZvdryFZ0Jl1jpRNN+oRIS8To/8rHxic2f73apWcAdf3PIqm2a750aimcbZhwY
A7Hgexq2pDrAglE+DCZpitNP0wlYj3XQ7AW57xvJAhz8M4CTO3Lz2087mw4cW8auuOf0tCRLnlpw
imXOEHrNyOmseniJzfH1m+nsZluuYPZ2ZxuO0kGdkxvDkorS/qDNXJf6WZfZgf3dGxn6zTVq1lOr
xfFtbGYuGES0Co9p3GqhcTI3NdP1bVg7nAWaCZZn52JtZ5gsE27jpcrCQBH0vqHZF5YTnV72QNDL
tc0nM08YR5HRJUet1nd6UiVf0pAJtUy3LoBtD1bniB/WBiLGjVONO65vxkugIAmQ+a/7olPHMIsc
yW5sHSFbhUPbTEQcwPTUrOpYCNZEQsfbZzMTpjSQN7k2q929v2VF8RmP01XRRfRWemgTuaDU4Q5U
4T63/eI25JWiEbmmPGYrm8DvGYyyGAK+Pgqew3fI+DNo3P4bD9zPocEfoewgj7Krt+ZdSsyEypz8
HMFgqViVimskJPZ7XEnS+eALd31+hmLUHO3KrtVrkHqhg2bmFoV/4TtvZ+9/YA8EHa1RQWbYQL8R
YTt2nsINoE2j9sTuG+/jtuFtjL2djUEZYdLz8m/i4mlHqRzJjDWr/+r9LivtLqbHgthc6/snmaBk
w3RP9BHPUI7GsFnOvto5TTXGqYV2d3VBkROh7XOtmUmal7yaAZXRX93OIwsC3Yrv9Z6ZZoJs9xMA
EsrsCi6Gg4Ds7wwPHg3AOWyzgKNfgdZyTC3TwQFbDB35WeydcBg/DMT55o1rLbBxlwYMyTKubTpy
2gRptlwaG5EdpJFDRZG0M8IXXbQFrqWEXmd+xKVV0/dJSOqUMNqNWWQ4tAS+hTrebjUBrW9La8LN
QBaRTcxW2A43SORIFu2Dsnz211MpnoWFReiLlbARf1ZBpOv/slkIBg3h2ouIGE+HiQH0JqGu8r0D
4HSFCm+dFZR4pVSwiYG6UPgARSLCrWIg8ulVpFYZRsczgkEZIj5rW/wXSdG0BXllRdCS5GL4+P/n
YY2pJegmtYx5+RsmcRuFCityHbJbBDIIUv45JbK+7zClpgZCOSM2vcgfNkRYx0jH4L/3ozfgvUq9
PmjJIlV9xx2jo6PIx0JkITDn9EOOh1VPQtSkpHD7kDmDB/PuATjiA/2OfCHRl8gxx3fnHucJyroP
U9eBrYccXM3hIX7wDCNj38LJ7Zz00ybP4EPS2/riSP/7kbeTRTmUCqOplba+9/HPdAgjUJ2suteR
hILeYkHlWAv9Hw7/JN8wlawKs1fIzFmbR4semzzTmK9tVROIZ+BwThSl+oF9thEYM0jeJIaFap72
O87skvDgRJCgftOqN8QeuQEBvzN4RUYWxUAGIgk0OY0HW+3xFPg1q5z5yAB1M0sx2LrIdiaGOGp7
GjkQ0/QSvr3b6J50j1ZFCl83+n+9wOTWBJ1pG1/qJSowpzE/HKGwxpZtE/q77puU+z6cV7Wv1QcK
5I67PadvgMwRkchAXbfF14MPdYllksU7OCVcbG2emtnfCI4yw0QjWJKhXMH65rQs9RuStVP74P71
N8Sr/+kxN2Jh/HqpomdkP5pkwln8OhjN7eJofPa0SYzcnttNR/VqvZfZH35MYqKRPWzKrySI2aSA
uOOHk/Kd1EVOyWs+10KV6ottgIp8n63PDuBbE4rzUuC6TmScMlfXc/bWGPRoPH76DA6lhRqt3w00
KzJ8INnB54F3O8DFdq38yWy5fPHwmnqPaH3ZB7hnj/H5X/wjkSCsMv6Q7uPSzlBKxiKjhbAKDGDX
19SGNk+I+28MCt09CfdTnC/j/0XhQjYOMg8mPtwtA10+pzlQdlTKOJXyCFhP6jfqn4t7lkotA46P
4KWeVy/WaZujjSgd4ZyY9thEO6Y425V91sPkY7LWxi+NYoPJ3ROhLMilEdk19qyM/Lyq6fxo4fXG
wVvkZrXIs+DbXcLp8lTXkomK7VQJmTYJ8+nASyuRKgy/W7h2HoUUJmyJ603CuoPv55OyXt+zzA2x
yDKr2KYg64KQgKZFY/GMoHy0zkJfzJYGqazqZlD+NoLq78XJtUY47DafJt8FXSD1nzYD7T0P6J1U
ZwNkRpeRXTmd/dvpI63VvOchdU7h7jw96ULTK9PaQfuDgqJFEYufoylKzD64mPdB1glnt9S/Y/Wi
Dsv9K0b5/44ATYu/oH7zjU1ClQfqFDfqM3RxfIUsmpEY1myIIxf/jCvlcgNUIym9WWa+G9kI20wV
7MHuEKipwY5TxUIIEI0g40shUptgV4E91uylVnvZSTnY7QhJkGm20l9FH22x2NB0haHvpuhEY+Wu
R8iFizTOBytkWZbvAnI3Uchz6pusVxap33bkQaLqJdEGEpLdBc71yPfGGNwQvrQzhCZGh8c7usyM
WhvqTMw+NemtGg3cf5+KBQSpLNdVwsbTrAtq+kmBns93llaDKqAhRqVn+OWjYVqpoiCyOAUuLX9N
8RXcRoCsZokt1ug1WLXr0oIsJR9XtOf0oRFCe7c+a98XHA27G9tmMd4uD8PdjZa2W44OUQnKkM28
TEsUT85bP380v1yW4l2NKnrCLWrWmF0CDDzD/Izl1e+QD1jtlcAVtwwGdQrukv0OVGEFH5vyFHQ4
bhW53fEmeYAw5QWUz5GZQMuNBVfA1R7y50aX4QZssOb8z8Aus62Wq8dQSMNK2KTAFyfmGGHjBguV
Gy83nEhyOsRBObK5lb7ZV0DeiBFYJ88DcuCxzR1yx+KUaYNJ1HqehojcmQTk9wcPOdwPm1vXkP3k
Eqo64CIFA3eS2qEgJXS78JKS9/8+Q+s1FqxCHMtsB8cvRp8bPr67LjBPc1hOzJQvqU0sS+UJeIrj
g61hS+wuRV28IINeoRUlk8BL/Tt5N3zEPfIoUSipfMiaItTnYbE8X0F5ilSuKfxqKZrfuvPwDgE2
CzBV+pJabZ+L2vtOyVxZJwRUHq8g+ojYLmLeDl4YB9EomyVyYSTg9/xug1fPr5gEvoPl3pbEt5Cx
VfUxQzVQzeqMtOKqflLoqdV8rHIqV35NcAAcJMWoEYwxTFgr40RuAZjAEHGgVroh0ntPenta95js
X5VFpLt8nrZy3Of5CVqR8XU3rHLYJ/RnXfNzjck39Gc61zhg9jLvgANAJSoX7RihsUJcbvsmet1k
1MKRUfWU5ayyp7c+QZA24qkgjKL0uTTb+WuaNWwpolgH7U4VQjwe4tLN9JX9oLlrTzG4tzl/2His
5w4vq8ocmoiTQfk2VapdZ00I8BMpNKbtdiKLhJPodKhLa1nCGqaIRMZSUhiLLPJqMwJhYAyzHli3
q1lmkWgZ6bvu8s6KXCVLog+qoA52Mw+Zd7JhfLZsahK3QLi+PYktb5H8KB2w5M/KEZBiP3kHFEYt
8RZYFjiL+B6K6wY0z195jv51T3v8vv7NBdhMNndqYTRAJYKFuHNSG6T7IBttQtMYpMhmnfvoGI5H
sdEfzSr/f4Y0X6piOTWrK69/gRMbqBK+0NP7JPIxi03Ru0L6f/xn3JEKnTTFfPeoGp62hApl78Nz
UDDfRhViPNc86GTXc5yYQ0nsTu7Jz92oCSqhlynoLQVIRBww/9lDRywC/1Mm2yzFtcW8dF2ROEdF
rmTYN/y2TfXBpNIf39qdanlB2vUqhhWVJYdZICk6OEtSNfWEEwNh7pb1wQeHnJFIQsBHDiyad6WV
5/el0uwdBZkMLzWk1tkPq0OZQopCTvhNAwwjp5ZUTs9Vsi6gm0jAA+s3eoHifBSVK4FxHnIxSMSm
dwjWNBgaUNaJbQ2TOjuBRnQhK0yer/gUknrazu1WOBlZehh+LeVehwBQYIrS9NgUonUDANFu9Oxc
NBrG72rsVKCgrr5/CIehqQiKnJ5jMUkDu1IOdFA+TnX2ulW0Sr6bfl5xUnvSJNyy6yrSGGaI35NF
XZeI2sPXMj6L929tqCgxjhhTQATwXcZiOxlN5lPjXkjd/X0CUYgGzkjhJIEkCubQtWFNHiRS5dBD
zvgH+RfaJhoT7SVR+WxHRe8wf1ezZ9196mEwilgdwMMJHTVfkFfszF3e3NuJRdF7ANUh2lrg6X+C
pstrUjQ0uKhnx2xIc9Tq4Iv/Lo7tuguWwGGwejAXr5zz2IshFVWPtVyZMerTNSCQvhx0Ho/83d0u
DtidoA6j9lsZLACnodWbnYojtoZSoiDoD4z9tSiRRZrnaZRwWQJlrcC0nN5mLu5XGmH81vhT3biz
MYffrwaRuZlL8gCZObdnfJC6CGEgVgitj/9SNiNjK8yzoweRnh8vuKCM2yU1dinITFEqV1qiO+CL
ugWhp78Y4elxscWHMJBgM/qOIkQBBL4t/gafwy0ydEhK52mMG7732xtgysA+sF2PwWLg7GZXK7I0
Cy5t/zMvTVYtwV1HWCSdbwtwSqq3BQqVwUqzrRD0eoAU8rZt2lPluaxDb3BR8gdeYGbyVZY0IW+X
eWa6mXacFAFmARRX9VJUWPs/YhbJ4Q5FcINa9GdE4Vct1FmCX0wym7f2aANlshwRaV+FmyMLb8uO
dkeiIKfk8SsptTOpxorU5KTQ3jl4CiwA2k6mL/7QOqjNjI0mI3jquwWNMJo7Lhu6M4fsI96sRlIk
A/6RWWwqQzs8RpcfQjTyKDV2QfGFA8hawLv4QhHes/JSNyyyWuGPhp0DD+bNdq2dcFwu5n0NMTpi
eRwuhw65NWerM+CG97qXNBiDQP/ECtN8qZ3FibEeW0KixvpZEXf9WBVL0C/m8sNNCBBV5v4hkwwe
rpUCMcKZFuizFHnpownzLdk2uADPAfomEIBHkL3EKcceQ7+L1+vmbRWrbD9QOePrbMHpyFgm+8L7
wMoR3ELmyNIpB/7Xgu/XPP1cCWcLYqxHufONja1eeGu9EMe/s9ZFAHVee/Gbhn1OxKuzyZkKzq6o
BWn11gxbOPLG85+JuQv3b0sxeVTY274WD+fuyAomrbX59s2y4m1j+zHH4xp9nIVxAuUpu9sQ2BdN
QD4CtmakQHg219mscr/CF/1YjN1CLSjUX7DSvBAmlTtNY+ZGAsjNbPGUTy+eWtJe2XNcqJ3ZaqzL
LYnkDgwfHBdlHf1O2xzDWcn/LOtVjpBG9bH4Z885PADJkYNuyQ1zepw=
`protect end_protected
