-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
KSQB6jvMavxsUngPi57Lfsk366B/Pb+NSzsus2UCgfKQZaIV74etdxDLJukJDOfR
vQ0CrZzUFUKH4L+0O+6UjtK8ftKg2/O5Bk6KyQ2Z8k+HAwQt6WuxQaLpGimgCzja
8d8eY+uUag6Ssn3Jwli9vjfolxLXSngKNxQB+/Ed9/4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10064)
`protect data_block
Rlb1hHcJNclV/AL1twFrZ1x5sc6SeThf6BMohuMRxSPdx1y8X4i/W0h1VKLCg/Va
R86haT+Ds06f5KVKqJ5Rn2ENdd+UnUCENPt2wfAFmOQZ8y+5mxdODvcKsj0Mgy2c
njoRB54lnxmpUE3Wi09NH5OnkvLqro/ED80G9PjE73NLTHNrathLwIeKJqW6EC0r
w7mMvHO7IfrtU95YA4X0rugPChxyoPnvLLgiSjv5HU5V31+1G4zXvpqRDg3Gp5Wr
kzUT6fbERe3rLQjbtvDVIkryRdf+jwHmgH0ehvrVRcRh7pC/evpToWu2YSsaMley
R564ZS+nlg69NFRmkQp9wo0ETBLdiNW+bgJ89WFoOak+milmOdhOh+WDlUXFNdPu
63LQbXy4KGDVbcns7eVyhfhQGNvIeAyBACqZbLPKM5Iz0dNDusz/Lz2ppn1r8k3J
0Sz0ydATKyyFnGRT3zBI0uNAIcNdDeVE/NR+4fhbpKKzMqOVYuXJWsVBUK3wmsJC
7F43RGMai2Vous2rVVYghQoWXp+PWEdr7UyJvVaiXH7RoiNM2o0kWpDQl7WYehjE
PqXvauU4/vlRQ67sktzSyliEL0wDXNCAYv7xVdz/i9x3P34GmLmGR0vMh7JmB3mQ
pKsKNrnyHIq1CgFDneagqeSZm1c8prBi3nKHntm9shfyyl7oc5iwgdpSSuDQm4b2
x6oGSeHrNtYIiSJik6/kJ3foaSGV3DBTB9lrbxeJdBgVRBWwH4kBctA12IyAg397
IoGX85XVKxIrKBWTx1xS+AlfGeA6E8DJJg3U4VGywvtl/cWOOuFCNWCJkL3gCVQZ
5St/7PL7BmdrLiyCZg7EU8Pos5cGdVg9OHv7wgQJD8+Xelqlk3TbIzidUKL5IGAn
imnQwUMtQDd7Qt0veLVcnGPHakuLgn90RJiT7t6bHos4hbBfIzc34iqbtYsAdXVQ
0aUXI4B0rXIadS6H9X9vp+dsSIsku6ZzTsqApfDMYbZGtvZn1j/CHdW44KuH7WAC
gzO04x5OqfgXndWyE+WELFIjd2GXMKfnL4WggDGazuGQ4JG88jprAZc+k4jo+7Hj
AFkvgjNbjS3xHXZecCEp1wjFvXryv/Kta3Dx0a++wk13QaO1EYJCMmHidd/2n7Z6
ze/xjlCgUY/xTcat7wFle6n/d5NeglouIglMDQlEuQMmOuCXTyOdX5adAg7PLAh1
lvba+1xTFS49xtaieWp8V8xaExA0hXd8rkqWmRu7jABfABE0x5CX8LGrqjlgykNR
Sfje/4pDpOgVNnZRB+FZqzQpHze1yrueBMakG4TmtScMCIwQ30t76bozfr1j7rCB
4UdAlj1vtHxe3Qz0jnpPQ6KSyVxABdzBRK/Q3tsw5kSKFVcqmg6VKNGfwD6rNz6l
a/dmTOPeHV0czEeMjGiUL/eYheGA5Ml2EKjfkuEKo2GHqZ7fSTDC5UWjxV0GZWMw
aSEsPZrTlGZICQWOTOvvWeTW4PvDKbuQCi+Wx73MAGqmxHE3pZ3blnVuzh+dD2Uh
PKtOQfECtyjIOeNo648k4CnF1haMLbwZKdR1ovo3IstII4vr4CvL7w39/XVcvNTf
TP5TWZNF6Y1jkvwL1ymWbJsMGsYifFadXPMvRzXxrAtGagpWo8TFg7Gs8OGasQHb
D1XSEZ3RApvm3DGk2XxPjElLhTuigeOlgEOFwH5Q2a4JBOOFnSjAebdVwdKkgaeO
l7HcY3Hz3r695yWDoHy/BByHmCG8tae0tEEpnh3UIoCdGp2LcBvi//yBcSIR/XNR
4gSnlmkYHS5sjwM6StZctNivTZEAnGSxttUOKROOYI3YiJTWgXk+sbbhVdsxdzmx
OeUshNYp6V4Lsc7kj78/A1zawYyLMumjk2hOVCn65t/yw2NJHWbjvCisjfkR1kuP
xTN17LTxQNzsFC9yuZiqY0JczaarSpXXzsadk64IEeThl9PKrMTSEveoDK3WCpOj
oxL+CqJdC8gIh9Zhcy7Qq7bA1BuO2DFnSgBp88fOIO9An0v7rKCm/XSSfyJ4Izhk
ed/cN7EPcyYphqYqegYl7Af4Vq65F9rKOK+yo1eQu3atlgD5BI5ASYSgKnAux0HX
U4RmXxbT/sMtz/QMLQl4Qp3ITTyjr97JJrmdsnfoF+L1cDdI6deXLxabpXsqmpJx
McAvcYE6pwJV2Uufd04t8k6TPVwueQPaBHa0dHAN4Z2IkFndFPp1V1Z6wGbXPwhn
NbvTqVBzdI4Fiqy7BkkLKN/wfhIgo+DTm9Sx/fBglfiSs56U3rwLaquIcKRX7ZiG
8Si3qBaf3DgTTnHRrH/MAYxsOj7jUd5JaqxG5f3Obx9bvuodW9015CJmu2yKZe9H
Q+YRivdobF9iXv1ipWWUhUDac+hczTrpxrNIpVmAt7uLIHR9ryJewCP8b8ib6TUF
9Uol1KtJCuUd0RzwHOQjCD457p+thDTPKSPW47hEhEPS+qke2YOtbj7yG8QEU5mk
PhhEbXZ8GEp3h4DOUK4hOqa8Oa7ugSlu+TTD/Al/9Z1SNsJUmUi7awBg4RqvzGDG
TJzi15XIA4i2MfiwN2U020/i+CfNe/yxejbj2kYHFlKgkVKwIYBQWOqawtcvSVdq
ywA8Piba1YjcxSOFaQMyTt/mOS3K0wJrEHrk0xxotKREmat+99/AqJfUW4cueqa8
cLpGNnT0NJF0CZNc1h26V78nkBD3PyGMBEv6TY/ah2pkz2S7+NaWw7ry81LrYKEF
r6CzJr27cyGH/qdX3EdP8Kcgfli3Skc8242heFOXMdbjCFHSsgQp/kO80vlpNPa4
IQtDupaHs/MvGipvfA8qC0b6UsGK5TVadcHt/3x7nqrAG+xHAybkJYrqYrubsxlg
vQlc86sIhvo5kz1bvzZIua2kVuBBqrQhDCtpnT/yD58Dud5z9xcy4qqnea7jnXaL
jW7isEkkwprGWF7i4l1BX6cP5JqoX+YNmBBxtQ0xmOnz4Z/YBsdHtctT8MeStTrB
rwDKq/I9ENFfuSQfRnkHpQL4pt/k0hsfaF1S6i3hDxnKYP5EnFkSkOTs2wJ8rb7j
Ibo0DxtiPuSjaV7jO0dD7CJdUwbsDNY9pkO9KizrDRmXHKjj2mBLXNmN7aZbXq0I
/zYIOM1b8nEykkCrBYtSxI0yeiseH1enLeqaKu6LZi7OWYfpM7/1NGqAMMvyOV6i
ePziOYsUMKXZ5OoLSwlGK5zdvJjJzxeiCqyLukxHEvaLUuOW0TisJAsgZ3K4GAVq
QT1wQxGWSXqXbUEcwQ5VsLlg1y7S9nCk/B79JbG/oaGnLJnGHLyDIDCEZj9CnYzB
KbYhFJ6vuJIntVTgXExBHIWqnGGEEAd/1dwqCunXBZ7YksfYh8yfHukGQfCaCNp9
wg6TwKjhPeDPUakiow73QR0raEFJukF5So0q5lCxNXVGsYpwKFHUDW7BJl1zJu+I
CMsBvIUM6OtSFaUzvd+aFyvGllL3vk0gy9XhAwxZ7Fsv83rZUrdyJE3XYcuilqZa
AQsJG2kcKH+4iRdIBJ/grq/WBP2aZGdrEwVnuPIrGXK0ADcUkWhC7aX1ABGLbXI1
4qTF/KsThnwl+W4WqHqJ68XTQK1k6VXCAQJHLJrr+TvZvslqoHdhiwMhcR4gg2r+
Vsa28srAR+VgAUOII4Etf0XkQ+c/zDaPwODso97h1oCAdcA353hs5OftnFE7zLyB
xU+OJLKnD7sjCx5l/8DFn55Ekjk8kTfRW4CX9VGAMyWrJqzM9+eepXQtn24B0J//
oGoBQtFprTggqdguPCsqyRbwejKNpNZSSNeBht6FUoXkzC4KO2SsTI3POs+KQNbN
IdQaep2x/uaaDailq29SiM0vzUAiLRkFMUOe8XJZqycDLR3Y+wzKvagzFPzEascW
O1+HbBIq0xX7lX4kve5ZUjrhRmkwzH5m8nHiLI8va8682TndY91rjBY6kpfJCbJy
G2K4quMxlTZ3eNf/TRerIh17GSIcOoU7x+3zNsu+t+s//RhXDuCexdVP+YgfWInA
2ZM91UM/bYi+KLCDV4rOzDqEzb+/3mGUVxC2e3FTnA4Zx7DVUfcDafIew4O/qjxR
h7thtZr4ae7+O7jz9nS8XgWof/iFGtQ+l8UW32/OO3LG6PPw1me5Vu5yLSJMR8CD
3Eq4mU8pgIPwS9GQy3LRyxXk+fEW2cfjDeJpJniIlqWKDUnw+Ce3MU6s+Ur9SqCt
RtHEWrRcwlVZgHzdwmuBtWp3uNKQ3f0y/NE3hZcax0H8l9VXXTUjU7f3wS+N7hcx
Gfd5lZ+ql56lBu8U7uivlp0vndqBvooHLdqXfdAuqIY5kZIqWCfSVjBJIu3xKmcn
6ghv1SRWfj3LjsIPF7qOzMGOeyL63kA1JInyP+Cherh0QmU9gagRtCMnVzLJLef4
8ohm/BrA80cMwQpl3wgcMtfl9MjmkxcnmZdAv/EggNAY7kAOfsCJncCFuoiLT+Ti
2Q7alUeJmCkJpFzRywESazH05coJ23QMpHAGU7dOmnck5Hj6Twybd0ZmkAFJ1IvJ
V6TG+ZUnTYZStdzMUCNhcoGwRbptF7Ov8Awt4Q0sBeNtjPJXZOJWMdvGU2+cYOyo
oro9kvk30kt9nmd8Fd1BxmsvhVh109gsRGZIIoBBpqs2rKDK1LC+57HLBKhH9dK1
lwIwdzS8YjXmiSqGhP2DvTnfcLJ7uQWaRQUWYF6JxfUADTKOFFj4uRiY++r4l7qQ
/a8As+DQ+5vKGhVvWCqfLH98TSJi8sHpkMgIO3cHM7z05rqXe+gg9VXVrcHL4X85
lb2O8RWxV45a/tAwG3Y/54p6goI2hhowc8K40aC2ctqb2oyINHYjY5SrfuNxBXsS
1jR5k/9v970GxJzcrcG+R9wMsfWPI5WZww+1D0Y1mScawLSFeNhezu9DbAW0/2RJ
TTALVNwS0p+8R53Or3oDxTyIyzPhRY6xNyssqB59WPOyfpIm9H35Ct76k7SbbbiB
7rTQXBzmyQDm+hb3rzWmG8U8WYeNH0cc8nhIpIvAqlFB6pkNDrDflca9RqOpOLul
+OdJEP9ZXhqGJM2LEmZvVEOBKWtK3qqPDSLw8MHdAd5XJmpwlSoro/+DAUSkW0Fj
6ZPSzNHZMEp+JDi7Vb8diwfdPTbJWyNKxIXB7+cqmzU2MwVAEZo0xXmOzEpq44zp
13MsJ6dx468+zihMBHHd+3kSdo3GnAFrHBy9bXsygqF/CbPaL0cflYkZ0nHBlpq2
YWXRRkQ9V8aE6mmW8VSjHOIbU2lbochQk40vYb8Zm4JVuTZMFlz51f/N4n2anS6I
Z7rGzrtGckZjvXyM1sdJ+1ZQS0WhQfosUNvVdU9A0RcQvMV/qSc4qAPohJbfeDGZ
1TQXSZyzxOLSEYY8FggJqx8CRGEBDYmxWl07QHqCnlLPeSx+A2EaBvG56wXnQgzJ
CcWJ0l89KFZjZ/YjTuap+aPctctc0TkEiXZvoVMXuOGD+ZYovZUr8bd4czKTWLGN
jPOa0SmMPlfw18+pMWxbHNFbmSUac+xykzwKAwKcDXgZfnAlP2XbUxOxLMEG0sAJ
JxcRkS/Q9iuwYl2jofsR5V0II/8QgzmR1kFPFmvuke7bOlfArZNfvcgcw9n7dyW1
IY3QrXp1NeYeHrHEmJHnquiHkBwbLavAJ1fd10xHQ+9D1ENnAvs9mgaxuSCrtgEn
F8SIGGz1EFfuaLotd9zksoqlFwTzvUkGTXFu88ZmxvFBlmZGVgPepsam83SaNU6B
F+F412l+s2BAzHOSrO6LPsdOy+XlR/e7DMi089gQbtvZQpMU4uAy6zk/+equtxPF
cbLleB1Yifonr/2K8ZPkPnAtJMWgp5vfAN87QnsJ9LN/dblD86wRWXFJwHBCJOKy
y23OFYET9/xLz4IWXA4s1Bfl4qKXrmXeCGU7JHz+/hyVNBp2b0XO3uDiRnsb5hvb
p7G8kpAHRFgtdg31Umded7BMp6mmVr/hW/mvKnoo9s3h9tgmAHIeOkQsYYuGk1WN
9snM6TjkDcyuNWEYmxshBpPpHJx6kWHTMdHPtArwJK7EzkBIEcH2M2Fsigvvov1x
wCFsyq77txy1th5Oy/nnKEHS9Wxa5jEs9ZU+ZcnrJIcOnAwdYihx8NERboWJxdMc
Pyo4bbUAXD0s5Ok4FXcS7u38ZMRkx0T/FbjOfcqluaBfzLb+Dw/KtHMpS+Mq6HnL
QSlvdxDdvT05//681Ey6EqxXgafq9wHtrj8/a68DhplBM7GHgWk0K6kOoCPJGnGS
8TaClUx6SfelKMNDVHeiY7mn+z/ATMV25ErXsECfK9l6k0EnyChUSQahZw+0xGqD
/ZU5+5LWDrqfiyodGMME8epmdkUfIhbHhgrjLW03x5ATaXY9sQ17OoNVDb2a9bxk
HQ8jjqjq9vqsgeVKzQqnY+lbePGzLHI2hmy+Z16/ocvN1qTP05C/GGF1hzRoJWZB
y6C069iPYRnBKknoN+kZs39GSa6wUMssCSLOTZ5X4eT7Hqd4wRLqSps5cDIyOi0E
06xlkGL7YPgxbE9xPq7ZcWTHm7IOLlE3V7AlgH72jJhsdWps1YhuqvwwoUmW4xhz
H11FxTC68al9B/L29lwXuHuz0cUEpOJ4OmFR+TF0Uh0S/p5YU828hCc9VxKjstx2
jKu9KW0xKpXzcKCX8zwDpuq7cUKjrNL2l2wlp0ABTxYPov50afnzfQxGDSBX/8vl
/7CzeHqsEaBB67KjLE1tfPfM9m4tMAAc5R0lnqeNJ4N02ud7KQgcd7IyJxXCVu8y
s+vGtBL7rgwH8LkH4qxHkRWv+Ktp+4LiyttYpbgukFxN4V2qRcskG4ZOlCyRsK9z
Zkho/g0VuDwrr0wTYYjyJ2fIj9OCCxIQuUQX37UQdRazo0djBakwgnsKenSw2V6Q
2CReKLPGjJGaDoLQnA2V7sWXFETnlFNGF0VPHP6OSEwjGKdgIKzunv7EKNrwiLVH
7BvNDZ91B53C/RDxzXGr803wdYtz2eUNw98KehNOS/wByaDjpxXAMpdBPatnpwxT
XVePhdzku/apysVwq6GDquv7aEOWsxUqCSUEHubB3Uj3EmSDEHUSRBTVEjyvEYS+
mOt8yyshKRtQq5NjyIHpcEy+ZCaFUjuD1XoD9cOpzyYDDuyCd/GgMxPF9d2IMjE+
NMGA7nGmH/l3AKgqIfCGUH0q4e+TsRM6uaJqShsQAh/y/GsDIqNnS8ceOZSE9ePi
+gBaQnY7AjGX4JAm3o5ejFqQ4UXb5HHW8QLtPqRHaU1qXd+MxW++Kk/WVMyrGmxK
83Yrwi+B1COGjUJ7iuKcxY83uMp9YDYyc0xPkWsikl27qrdGvyosy1CmG47cCZb/
do9bvSXfoyt7liDkZ7Aj2V+38mATS6LrYe8kN+0SB6/vNpw9h6kcnDKV4ooI0Pv2
Kb/zUSNsjA5Pvub8HFLVlxsrAwB5Mg7zp/3eTfO5iuGKaiUibEUWu8DLZhAjjoFu
PugtUjhA+RzbIJjzW6k/R5efB1/uAmqImQrbcfCSzA1TZChQWRT5PyGizfoEAwlk
6Mmp3huK7Ilk70CGiwu/7GhBxkUuZKoG/twZpdx1WvA4DYocct3zwW1KWjqNeQiY
+InN1FAu5g7LQ0LvjGWULTfztKE/x7gUyEt0XSiPEuW8wHg4yg+0L06qLzkayK4K
Qa9cJDwgo3Hu4zJ1eCbMKDPS+t1/NwUjf3wBDmtJkIIEGDhbzspf3U2JoCP8XSB5
Ja/vbYtteQyKafZ7In5xY6arMB2iV5bQRjFD1QZjq0uiKWSWAp61MXm6z1LY4l/O
zu+zPHAn3aPTl+Ck3gHB4Otp3Mzuouy7jaW7KgYw0kzCWlPeLWCaDZoYeW4rV1XD
xDmp50LebOFMW6zrK8O2nZAIHO9kik4+q7Bqej7FcrCFvT6E0w5sRAffPd2+MAoi
5jiOYDKVChOIcENM2RpswM744q9OjQFCP6vy2wsGBDzMJ2liwg8CQ0+/HSwWnwAL
sm1SQP4SA4VhCjywqtgUjVD1aYMMv5oxgWmGnDtGeFhsZ2HSTYJr0YcYYLgxEE8z
H1hXbkYLlIBx4Fx/BlLO2WQe1QRFNKOBqiHHbuXXPke8v2VtbwN1lDjZuDiFzYLe
Hc9mIErLO3P6+RXPPUTc6A4qTM76rLl82QlcRiTvYpVNsHIW7c9TisbKq717Pqpt
08rnYx7/HRBLMba72eAgfnxqi+mzEY5Zc0YMuxUcjSXNGD08wE7oL6UhrtFEG8Vn
uCBgP2d7yT/iqOEINBmZZcYQWp53dPo91f0WtuANMhGjLUnVwnaFFcQzSB24s74R
UKzNVaWuHJSnzHIgL5HMkVBS9Ov7Z6dAOK5KCRL6YMr8jBzQM+SYNy/4C+2yRfKN
9LoP+RdRIDTFXHtyPlo5BvnHtGKbbD5BE6qSaX1KgxML0p/OJy3QjOHA7RNlmBm+
ihCgz5Yvlhv0hlEEXFns9jgbiMX8owMWHni7wptLpETfSqdfrmDFOiKEzfBNkTg/
nZmZkcgd4nN0kywiV+f9jEbhjiR7k188eeHaDVF1PrxuOLr4U+l9ZsCheZop6yjv
uBoSdRP98yScootzaPmNxQZg2qYERkNttTsZ1b6v4aniS1laBrAqXdpn/TlhaOEo
Bp+Jdnl6omhMvojistfC2Fimjb7s3TVJJ0qpH95dq14qDH+bghM3NiU52wPNzTyR
XnqdPsXLJBfq6D7tAsfarHA71Ccauacy7nmAc5q45uH2VMoh+SAa/m/6hlPf2dlv
hskBgWvU3dIeP1uIoXVyVI3LAQvR84ybDmdiR12O+bknq0ikrMVsnhhPjdgFvbYA
iXjW70JiEW+xnHx/nIxFeBsbg5qIeueRftzgfS/dulzK9x8C2l8ocVMUrKWg8y8n
hFEVZUOsFksYmlSnqizYdD6LDg/HRAcAXXBSgqRj0R8QgQkdC3hrVhf3lMmh37LZ
tD65txv5oZ+KWc0p2IhqyHK4n0S8/1mavGdfX7+c1ELIVy49a28dssM+dMoDUbHv
ImkYC5Q7SPkOOVeuGgUVZXcQcdkmT2v/8t4WrkKy4z0SMXulTsE3VodsalaIxh4h
FLLOdWpQ7c777qas/uTcWBFpWunvT1kBe2cMQUA5JwEzxqVb1tjGjBPCWzuagM+W
uPxFF9ldaarohkRg5XKTRb7YleGlkQ40wptB+NfCh54vIP9Mu1HvMrrk85McqZbf
zdgyRvrGa4lod0D54onKY2F/H3uj+50PiuOtOoVOhQuEYu+5+YLGMSATjzul0hMH
3P7VRY3RWZ4J/lNSKJnF6lrUCE9g4JXNFAP8HmKHV9TrDZpVd/klu24iway9B+68
EChkY9Oy9ZTMMeFtNtm9WE4zzWRbTluG2CQbHkbtu6PsV5MiQL7xIMF7mk1Lsc9s
SjCJyf8Gcnt7L8JhlErs3bnjOd4zZQtuUH4PaARfBSr4gwBdu50fO3EDuCr8/g/w
+2hOCA0/jW31RUUVnTVb2gkR8i1H7MFGEdo1zqVOSsvicuXpBbG0SgXgGtcs62HM
fUtfaB+yvoRp4YuSI1nPWnEstda5naNIfAv8Zg4CWa4xPZP7Y2jJSnO1lpAmiCxJ
loFeB0295WOr5PhTllJ60v9yG2kizpsiwxldhJw6240/utS0F5+qt606j7DkH0vJ
OUE4UcaBFsaJvDRFjQATraPyhzqUvRYB5CzAiGSINifZInitoS+6Why0TJxx5csa
w1X2WtrllAeABpD4CRzVAI3J+pVfUDjtosC8bZoMlqco9PNFlVwLyyKTYU0Bb/IS
rSPehEGQul9loQ4HTop8ohd/V6dwV0HZX1tZxNqYDxXpBg2HoSoWkifAMA9cgB4Y
nex9lgljLnpv4oE9uSeYN33enJC0XiN6k+kJnme0Nm4X5kgVs6MCmb1VC2aYTdqd
XhaSHEb/+Rcd1T9gH5R5MdslVQw0ufFaf/Pws5nSpOTvrP1eD7eqMph4EaPGJsQN
doyj5ZMXxGS3zXTffydEvImFmbNex1sWI0puCqfWbb/0QV+OHYBfVY6wLKUriGVV
660uN/PPLZBpuhYZx9FDzYLT8OkBjUE40TEmVz8ndYulju2cuUcTmtt6BeNSGAI7
tHBmdXbtwY4s2AefeUPhRz/bEthAi1UnzqCIfIXAMvYV2nmf4jR/RJc3/rwUEyhn
xpiygbG59DKhHSVYGIWMtHeB+zdu8lbjiUYkdj0hDDrmKz/hTjdC1nCRIxzi6kHD
ltXw40twrls4Ee5kHxi7QrP0U0rB7a8TBnem1UKMH4TuUOzAkdSpmlO+NccV0H0T
5Yc/kGX2KPDb4EqLsM7t6BN+kMYMm19lE4B7/nApU9ZJ3emij2cRStCwweTWg9Gx
VJlQ6IIoZwiG7ucXqONr/1z2GbjjvveaCiRnEnPpqzLslMtXHu/zwwfVTMteyvCP
wDYQTKb20SDJnOjsz4J8mV+tM+5mHsPheNR3lLSlE0kHdTYjqqUuE96LRWMpLF0x
1SfZHcP0PFlMXn7GxFz4Hh8hNWJpVt4uSnfKCL35TCyIrRu9p59n/LMg+k5AjZgl
mchOrVvGiVYcKG3FdYzGdSwFFAZC+2Kg1O4J3QMVQiILo5fYTXQMvj4vN4X+0/OO
2E2mhzj3J4+ZcQRc8TQzfpOujjurzcg/GXlAeAfgV87Jd0LGL9jR1j0QoxMx6t7n
REZXvguGl/8VYw+ceSeQ+WjpAnbHQDHRrNYeox+wZ/xaVGwQvVD5GKvErb/9jT4k
X96pZfN66rJ5TzELWwk21EohFoUbLpD6h8Cv3alozTqiX8/u2ciN8copbh6zQbB/
O3BPnZcF9GE6e3fpmo1OztmenTzBzmtkXfZdhFiKLKjUmanyTnctG3eW54ozmLb8
ULcnLHcgqHLCV+BUayobiG8ABmMrHxz6dEqFZjI3Kt/dkiH2WcJZkfA8XwrEu2wC
jZ7f/QRxu8zPlyYYhZpUgkMaspYFc0CduDm3OoEwu5awzr5sL9LiECG8ETrSOJKE
B/BhVKDQBPaypqqHfwCpUtwpTWUl0PsVpT0VXoc+to0MusGV4Og5aU2drTh0CPhK
/K5/xFEtuWV0g51g3yBrR/UdIXiN181yqr4uVFqUUvWslm4c4evmAky3mir7NPfj
y2YR1u75XehwWAt/HKhFcPET+XebziAoCoPDR50SjH1KGwacJwbM65JVcC2dcSv4
VEl4YSFqaV58jNfKFxoi1LGfMcdXYevWwYwuXEf12mXygrg4VA9BYMhdwQPil1Sk
1NSYIoQupWzp5sDQEdJrOfT5Fu0WAuMgNdn0flwmtEVkHGCGglILTi+xrWfMACN3
pYo4KIEcxcjIdWDJEokDEXzE3vQ7tUOhZVuLpOo+LZNe+K2DsTEMMpwUlmXr/Sr6
LuUT/vPxXqWDbqrkwdcUykTlzMsYbGFbkABW2doHC9eGGwPjPkS6pEiicr46zme6
CwM2ha9c5rD8HKW4qjf5MNPZvkR4aTwJetJIUnfTtRxxajl2SjXEx9FkcGwzvI8P
fDeZYUr3WwUCMotaPbOOVnqCMLfkkUdHtttYeycmRjrzRUJuKV8OHhAumjTTrZuw
LBMjOljpotJhoS9EZ/ioVXzKJEp5gVqL4j50avCnmKKq+FUL8ZqhdVvPUnsRus29
mGGBXUnkxwyiAPuaHa+ahXwH+B/M2sp1eJrTG1zPbgjNh19a67Pse+l7mPnl0taY
fCD64V6ERoCQG4wdKInEyBeN2AMyju1zWElPRZQS8tAjX9pevayky48TVYAsZ+vd
TV1hHjubYAStb8otLb2rXiTe5zMvjLECMotZH5UmihDpuQoQUsLpBEifiMvMqvZf
taQ0WKJLJPMqpmnRvP4efgHMLwWsDp/hxXpYEm5ZGtoHo4dvqPVSoae8jYz77qm0
ZxpuYdw8N8vERy47nhHDppY9BQS1xUdpCeHNVwth7PaR4iAKXqMsHFD3r1bbM/+J
G+DR3fvzNQkWcdBdVvCd7tRmbKxAu12DAjvlCvW9qjqdsAOAg4Z2cVidngAiZ6Oc
e8F6Wlvq0xDXHYPqyPkwkI4POv06/dkF9wftPnUuhkDwXB0FpmZ+MsWU6KtZsW5t
pErxUi//rBAEDZLCKm1FLKPN6k/VQW285VgPRrlZAMPzYh3SK/3WAGiqZB/JKMKp
vjkvXU1qRQqanhJLd+km07a/XkZPfO/niHxt4pWVWYJpmkVXB452ztQ+Abs8k6Kn
hltHbZxG+JdCRVod2QPe7auOCBc036t4Y7GzhRGpiQnH+6P7ujlQ5f9HRz8IFYFo
4yFAfZEQZscuwK1GAAhDepvBGPXodFhI6/8C6t+M+bw1l9akbJb6inyQpoGwzMo0
LhLZc+4FHAY4feefpQZCV4CzfNCIwcqqxeHiRd+Wj/D83cQiScxHawTu3s05Q18x
ka5u/hQF37F9dRy8jPhEBMizJ4kjto1J3m8C8vyH1WifAG3f42hfBB9CSZSfNCph
LsxxLr+DzbHlughP4CTDNcF3S1Y3wjzGMXsezH3nG+QpAflRfR3kMxefBMGDC6iQ
DPVZIDNA3TI8srncED04AXTNVJOp9VZaviTvbnNOStetkCds2SggV0DOIeKYlbel
bd0pikvRUOYp4n959MtNX/J1xp7/03tiHYVzqQypHrzHN3+UX4ipqF+48zqI3wMv
qRHFiF1dSErRh4usTBXjijSrM2CIEzqBGuzEmEaaOTRwkDyXXoSzFoVK9GacElTY
+OI8JaXDTEaaNPSdDDIqj3RUyl0bpBGiI+sXqU8TZKFRHI2qMvtAAwkY7DUlIF5h
DsbJwrB5jGDecys+uNuvt8ZgV9chNvhT6GCrWGiCalGzma7TtsK2qmUUSVY3yAV9
/wSQPgjvFLgJKjMSBljOsz1xyx0X0C87KlK3sWHBuKOt799gntCMEtzufHQSlVwY
XZBD4sTcprbueFnRzcu8e3WYzuWaIDEhctVhrONg0fbYW0XKHI/D/7hfZuaVD7dG
RfFpr3iyEUt5ciBWZ5xqxm6qrJ8kk/HKel9Tfs+ZyQaw1XCPMC0P31Hsxz2Qg84W
eSPTF3yHlG10Gf0xBiu/RHNWiSC6o34NIfbuxY4guxgyKR8DQYL2zJwm3r2Dam4H
5XTfJAZzgt/nFL4iVVvnSsRBuwCtn9+ADgo7SlMA92B31xT47d0kefg5M8p8D4/X
KHy/9zq1szQTFuRzyzimOIHwAHMLCcke2jqWAvGdy/cfdA0Yz1NjblL64fi5BHBB
qi23k1jfhPffIPM/Jc9ibj7Rxvonrgawl/2wXDa9DgLZLxDJpRS6jhiHW+0BMJ1/
+1WCuKX/7hkFRTuRxZxtgxNCVpdL3q8/b345t1WLmd1AYRLKHHyU3fL7wjy407rK
Y+JmdTt6c6M1k4OvxHMIV0cMdCi1NpkYmvljJLi5at0=
`protect end_protected
