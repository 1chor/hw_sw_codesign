-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
LinwWHje4pD83UHa3KsMpB4YMNiMe0ZSloK/37im68ZFaYBKG2wOM8kh8ypQ5u7D
avqgalTH7kIeyh8u8RBruFZwttfZt2lhHgBo3GTop7QAu75gRyn4yU6ZkxCWXvVL
rVbtl5DhUbbmUld0HJ3XQ0AiaZUd0qpgSdVyElSWcxk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8160)
`protect data_block
Rc5psn4MeJdfwLGIdrxENnL/9z/9P9RQdhqvy73Z2nKK7W79TbkbzjFDOMQTWQls
px3aI4nhU1qBlCVkqhk2cjxN/5Ky7bQLn+j5MP07CzyAqK3BToRSV8fVWoTBsZNk
Amil92aNV0A6ghDtUYM6DrerJ/gow50ENLvm0MCS6ez1u0i7wWSTUmc+aPIug/+c
NFOpN0lXgaDdxOIdcnhEwOykuKUpcqXVZjJG+W+Yv3Zgdc9v9I9M/Z0XfXbnR5b0
QZ/ZyAayjJB4be7XiyuIqGn0Tw0Owij0YusK++1NkGfMssBhMp5DLzS1zGBBQ/fG
yV0k8m5tQOK28CUCaNDDKKn7Ys9UHEfBLDUXdLfs7mwR9lm39q90zwc33R+9OFL/
gA5vhl3NIgOMMo0t8cWUSZfskNyXDlyOWGsCJEQ4Eg3KwVmflJHZfS3AXTbsGp7X
1jb7PEX775sbIiY2vB3coVV1XgAyirxB8uWqBhH+a9lfNbrm5OkWAKnRim3ZyYYI
l0fKaKWVyJrUeDe/xdcm5oxVh7zLIJdvzDG9r1x9xHuS4Pyuf0we8iCAj0c8YF6P
qHy/jGURbBz1hpNNwF81pP2zUaT3WS9WbPyldY77XE+J20NV3qxdfOj51uODmyhC
d9zywL5gvZcuaPFQz79ZhccUFrQi53h6Fju+N4WRYoddIcIBd1yS/RsO5EkDFB1S
6h+UV4+xlqoLySBJxHm0ji2pJGTo37ntmuhNWDPgEpzOBlIu2OwEsHOfiTj38JwQ
K8hNsBkgDmynf56LA+di3HysYURqQhMEsGXvRZmFoblI6Ne2ECsM3XSUFC8eVUcC
sxqwk/aBE7wjfMLvtBLtojIiT9RvyCHCE/hzLMT2o3mjl+Jflf3NUiqoWuSoUyxl
wMDoCX7XNfReA51o0ZzT01B+wTluMtumKE0buOu0FlDgfpHqAdZefc3b8O15mEI0
9FLGBNIfJGKFMwNT9gjz56N+R6f+wIB2llXg/OGjl3tyLTCiVGzhgD7uqRhdua2L
datPpPd2J6qhYypmZtpOzjvGX78GZcOO37Za5+jEhMHyrzQxGNWD45IzpdeQ0PvT
S8NgcKPODPzPDx/K5tJUFBxSvJL2VtYmxwYMUsPbCw1rErLYcHnfQHRvxZ+gQtGg
N9K7X/+id0V4dnqMsQkrj6oUMqjqIWHtPFt/KtElaKtwgjjzSCMy4eQSzyIe+Dn2
g5nuSE9eI3WQDGoFYpnfqAnF8f4ogKC7vQ+wDiqTdfX0usvsxk4KLJJiWW0M6DUC
Yy33d4iqs+y2HH4xa9uOL4TnPScBr+7BuETGr4xYu3uqDGJozFwzVAeTzYRLT7aq
gW/AKg8AWwP+Lfp4TvfaTKynYJP8cOJtVd64QDJZuK0BZTLdUhu/IojCHLUKYETQ
3mSqgCnlkQRy7F7eo3JIlPJvCJw+42yHzf7MzXQurk7J5VaiIUxmh4dWfuVEZUPv
BlWLaXkYv+2CaANtJnMZ9cSCtowGtqpwXU3qZkMP/26w3o4ZKNG0vFDa8nTLI2bL
F+NBbUO6LhkEX9eE3FjEqayR2IxrLFWM80y+51UPb2JyABfyoLtXFGUNrtolutg9
8u6ZyQy6fta8RlyZxPY9ha4omy+6U9EgLrUGQXoVok1Rjee1dBUMHTyevv79pcLm
JT9hP75XcuED4YwGY3b9nIRUwOG5OzYosZwyCQKu7Ld5Up0Y+ecEct3B/JHpJeBV
iR8CIhOwEoamqZJgz5GP/dJ+65mOuQFIrDoqbU15Zp4F8KosW36NqbilfEu7Ryew
HOX20kl3UNXic93No1tYabWX8F76AWCAqOBpCcQbrb6b7dQNwuGjMvK5YW39Fi3y
LuHB3SzCHrkOZBSJYOm5s9tIb/BTYOGGbHXkX6qJsaGgZZLKypDkiDwW6T/vF9S6
yWXL0QaLBhpXo+WYgDTF4f+OqW3P6AAQgsjXVQE5L9iC0fc5VeyLXfiPMte1Iv9S
L2tN8FIrv0UkE0Q3haR3J2Hy3jf/dfKE8sIJ5MmQJl4V0SnHEdK+jK7l74ja2Kf3
9q8zJuZwav13s6nkGS9hejtU2jmOTVbBj4xtzT6A1WLFPbmHaEHecragJb/+9AtD
TlzPRRw/YJzNuSBjlk25MRG9dkhjgDy4G2nqZqPxen8pNioga9L87ZBj9N6tCQyW
XEbSb++n4ZoXYh1MRpkIeP+AWQSXRiXouYeJO9YsUd1h0FhAGYOyJ2VMLrWX12bJ
W37fqQDLvveuA5Y90AeIcww7dtKta+hWk3QOyQY/410nTGyM+9qm6MCyVumNC7jQ
jSitVTYQrwJ/LfAFtezUzG/VlW8v1chgJHa7YgMVLAz+Ifr2fi4SqPyuZl+PuEGQ
0TclBdtqdkY8/zNib9UQuzvSdR7ogoDvccvk74UToWBPK4CoQF9tQ84SetnACgzT
Gzaysn+JjPTbREi508I0hWQYA8jfm9c0F2AcC29dQ9baR706PxTisElD11eIf/Vp
tJf/C7EYMCM/6YyXOxwhOn21s4AdZwFxrTLHhRKBWiA8x4zkAxefTyksjWHTY9Qs
SoFtWpE+7B+On00K+UuBCIm7p4lSAwfjIFda4fPKFdac7dlOwwmE2t4NUyss+HYj
kwonftRCXAt5phjF2AFJAvKG2AEp5F6cMnXIDm/VAfG7TSGQcjOgd1d4wf4n4QD6
DmpKCAoToXqZ5B9A1clDqELUY344GQ/vI9gIOrrJdiiqIEE4+iCwu2cGQ80nDrtU
BbskHE4DZvmY86jhP93M746tyA9IW1cXJfw4EIAaJTJLeOgyJKxKo1+zBMAIMfE6
qOClsm50HCWzXSAuCue6eJRCTJf9zeWWheQvmi3G2zlPIlCSawoarPb1YQzwYZy8
5A0fN0wctQKc4l0f/jTFU5dQSZZA/r8Sq/5+B8tsIXZNmfNaf0osN6gwGb1mcz3K
j4EalVWOJu+zOg8yPorWQ9OlMEBHqjAYr3DTMA7pvRk095C3gjRvIzWiOWNUkNKT
UxCVnX5akMRX6pQvEmbVcJNtMCPm/KXE1O/zLpRte6pNPEDWezQQazwJauEBJ9Xc
QOc21qoRLaWc9Gsw9tsmkPe0oNP13q9cdreJKUgPsmjhBb6nmkfka/fzogJD2FL9
ynOOMmZoGCwcK9iMV0XAQL2lKJni+n30HvzsmMyYD2YwFxz7wl9kKsWZsdTsoxPK
a4AUs8egl7cgv15BtvVFcjQZW0JvCG0MQsREviDoPzMHQoyEztuBVqIVwiBb/FYn
mT7uScpUZsprw1yJ7DsDxHWY7u56xqVMV7wiafV5ylakc9YbhiNpmC0q2xk6Sewu
avK69402cXZkdW9/PgLQD2UfXz10FzgeR3j/0452nXTumvQQB8qFKQx6tT2A2nlC
t+Wb6L/2ikoofjhTchmE42XXJUlLpANnGGSwAWkCdfKHEDraMwrtx0uda3pfgghC
ime7NGWfQ+HxxH8AgZlMVA+e7Yht8XHul1p9ZTUiaDyCktyNjl3XQyuppreWqB6g
DjmFeKapqZk+OOgjjdERLQYq9QwetnDDw8eBU44ktR2w4y7656YCWi3j4ZssVzD/
+VdgvXjXai/MS/YuGKHnRd8wFkr1op1XaTLWfc8XMfVxv9wHWcgFB6lvibtxdVo0
YXqEiSwALSwnKk+EtlEhX+lkqqcoHauiuJYC6SSKTwPbdtazDZUPY2HiBj4VlVP+
7l9v8PHXkf6VdElCBPSeJDR7I6cnICMbqbR7X6vL1FmbVnkhuN2GxJEXGV+S3i/Q
w7TGKwgYq0BFw6B5MmTXT1YnKJZigw+WPsJHW7zhU9nl/w0E0RfTGxeNiepnA9r6
G/CWnjg7rE1/Jn8jTRpjoV5WhI+YKRW+noJcm0x0TXHOTCP6oZJQ0MhqAo3Wtvbz
sRwH5F3x54zudZa9gOaSZf50XPmcISTqAOvc2jUN/VDCQzYXiOCgDykaMsZaVjsi
W/s+t9k2B5DP50rldg8NXmH2OTz0qeR9Kp2hqRnLLrkg9sevFhh5BUWXMeN24upd
Vh/4J0bj2lJRaIGCmvvmzkQH9Vgr6cewEvxXBkGfA1F97Gpfa0FTRpuiQ3gNcc0h
7H1q85RiBoyoRC1GPsPTdGAMsg2r4nygBbJhWf4dNQrrAcFEoU7rpQTzdNBPvDdE
74NuIg3Swr+hqIvwj38K/PGf5H+4kBvedgapoVTGxV/TqzZhM0B57MxjtS/KN9JE
TZdethYuELE6ZZ5fuzGfO9jM0i9mcduGZBQOVYW64kv79dRRBRyfKU2LmpxKOjSt
HinK0Erxo1Nfdfwe36eiub1bBBsyc1ZtG7h+j0tKhxmDhRYT2VrblQxoKAFvq4iX
pfQYBs31RVAOHw4hwII3c19qHEFo3O8EpoHGbUgPYcrTSRNZnK65MHb6iu9hsEZk
yjWOkOLYeC2vmSW7f9YvA2AxZGH+Si0HKhqXX1WLHpmguYf1CPdW+LiFQrz4z2AH
6f/AyUm+Gi25SvoVUnPlvvKRWGHQpSjI+78o5ezJGCnKqGehqppnw++/ProNp6yg
BIAy6mQ1l4srgx0E3RcObl9UsdUIEgXF01HBFiYH/XO1sx+aZOKuifLRNK0AImrU
WGnbB9OGLbTlajYhxarXFIyfIvOLb37NvQjv438wiXoWNPADHCbkPb0aSFoGDfMs
MzwPe5rhOPspGfkf0S0OPVnbY7lGjATMdaiO5fQZliq/dhK1IxmhyWqYh9ZMFwKN
aE6MBbCqPmWoBJnomoSFKb4ru3iKn2o4hSv6kCBoG/8GsORF/ZoEtTXl4PovQDsQ
RORryYCtDHHhxF8alom7k1z1E+Gy+ksKz6Znmx9cfJieby/kCxqv7qeZJ5Ad898C
+KyX3uwWXXtzx0r8Svrmzal68ZZpZowoQn68NkwSJiBZYJWiUl6DwA7GFuy3YbK0
hWl7qQuaPkUmzWHuDsj2CfiOs6dREr0nWXMuQ1/t5tgMc80u/0eNBftkGXeOR7za
D8uePpOfNOyZ5BpUZH7slRKeCzDUl0lA5jdytPOs+sO0JZ+V8+sFIDbFj6ANnJ4Q
YTxehVZQ5scO9AmoIC2CtYiFaycxRAHLbXCf9QcgU/0PxU9kFyOzrzeWYTUDrmEx
61uRwT0QluxcTa1MZSSQCdTywCH+G4QnL8xTMB53pL9PGkUMye1vCsXUvptfnwTq
6/R5IZn+dGtG+8L3mnjQk4dxqDDAmWPzZss7CB6sCLTIs/OeO15HR1Gg077q9k5L
lyRLCgJH+BOVw0p2kBGyC3PTOk2MuWSzEpRZFGowL235sApi8UK0nWGm3qy8BoEb
/iLt0UkuZi+1wx/FownyfG/NW/i5gmfHYWIp6MgyTifVALjMFaeZtSF3g927XQ9K
ubriQyceRf9qaGhTVDbGHRWPQtQcZXUnO7WHfYmVkbEEEyVtKxM/cVaorueJby8G
8qRnen9P796twWxhum/TLo38NRCgGvZGgt/h5uzggIAXapWny5IK3eX3QDEsyc7q
A1I3guerko7u0etDArL9GXTXAuQfYVkU50vEqwRCHwhlSv5exXgZvaai2eP+ft9o
1XXwTHqr5zsHbO6tseSkin4kvSXhuCd7sAzG/8CKVyIGgyItQWMWMSJTh9L5Dvmt
BclEIyXMcsFzbtZpEYLYKqpnqpnDUHDuIBZV51oB6YPGxh8SNuj7XQSpvpf7ggNq
dgsxAYDZmtN2sroT8YS/EKfzB4UzXJOPJBCa3vEPh2Rkew6deCvX9EFHbNLwMQay
VKfUjL3fIS7T27bKNGKPF8ivm2u6ORIxzyxM4sSq9qI/agFWwCs8lHCbVUFVYZnd
FuUHcteT72yfJzibMXtBIIIn/wGdem6TRqoVrzjDagUXJlx93YduBnxOIdEqCsAY
1CRaiLrQKiA0aaSsYnz1oPeD+waRl901BspNXcxnghiTSW2Gqj9Gvh8ilvPO3LTC
7WTpUs46sZbqL+GkqSPcuhUA4os7WJw4nmcVl1piHhxtU1jegCq3t3sYqln4+Ant
Mw71NDZyIyIMFCg9S6JDEB3E2VlFxfYwoMV5h6DYLW6hcADNVP2eP1hGw8oZlgj5
WPR+Yrg6jQW3wt2pSoYUa94OQvS1aTLPp+5kOmyjA4yJfj4jp0/cxFEDi2vPuv/t
yoYMCK/quMpbtJWt6xfFsebqvQrxW3FZ8Qt7ezJMAR4gu7vd2PqlvjzN1pCxeggR
Pz869SnHVhP48vWIf96hi4pFQJ4tJvL9apnUdvffdYqMK2Y1IGqosST9BJ7jwztM
37Zbkv3ZezbSgjjMNL2ROr4rWCxM9e41N/WvclVILrPHMPAeperKW0qk81z8AqBX
6dwJ89XoiXIyunulcLygguXKsACsECDeP9k1SyISQ18VKV/hqdxv7yv3Sewrc+ge
kYCJrZ6D+FKp+NAMZSaY3o7Cu2jSjiMX3UPIuYIMwdlD1WJSsX87Ay7v7cWBPTKq
+O5JBfNg8apLkgM2i5b36eCsGCGH2+7NOcZXq3fzq+XxlTD8cJn+bBXG6xQFd0JK
OhLpzusT1nlCHXatuiexeCN87XutIW4Thll0PD7vGMuHFhwE+7TwFaUi1cs8Gtfm
n4IR3/1M2WAQ+FPX9GkR6Nj+Kyo8/FvfTo8icps1psYHWUMz1KQeHXLQndJ1G6It
7bC6HW7Hh35zXPWW/NPRLQmrxf3AsM6xVqz2SEtqX39g+XRO5vfgqofkXV2TmZp5
mX+y3ip+xOljjILg7CaHqR7BYRMdqjMbmlEXI8yUcVPH0YjUh/JHNWYqVWgsL/K/
TdG0vFNFrqsL1lnyFW4WxW+hMV/MpppHHx4BPh4FChtNX/soUlcPtMYOATGJ7pVf
N+AYEgoya+ppDuzWD8OPZoZRhdDBObq7GBLiAv6UT5e1ydlueVtrh6l9icKFWACj
ZEVPIfFN05jSbAqE6NleGh+vXZTFBGgj/pKY613deV1CH/elftm/jiR7ro9TL3M5
+uZj00avZ4WaHpdMpbqqaUaQ1D2mIKMu+WL+MekbIiaNtXXYx4s9RF8gj26UFplW
GNap3Ym9D8MwrwQyOBj/86ul3cdcWbL0XCjmk/gTPh3wo7d7WjgA1Lbr8ezt2KMV
GDT2JCJ6+ROqxyDMH9fUMPBI+Srskd/7VShmmU03TOQfEtBmJ5sF9gDhVJkMQmx6
0tXGLlDua40XvnLv+9wpYSEZ5GgQ8N5A9jg8L5eHEKSqQro2SzZUNrGAVRSO6gYi
d7I3q1m38h0CbeDIzVb/+F1+qkhxt9Rk2V9s/5IVYV/mgW9k7fYP88yQCEoy5tt1
znyjn8jXZgR8wL5i2jLxfDW4nz/5c6Yg5wVcpsqWeyMJxgJ4ONXP2lcP8XI8msWH
L+fJ4OXKB7Eqk6T9bYqyBroqSFLimt5oCiHE/V81FpznGK/C53FJ+LoIZrlDHFEq
u53uimxUOxFlCd5iywxzFCYoQz6zKUAOFf6UQqiY+yo+UuROkT1hene4Z406L+zk
7WwEbTTA5uatKe46EohfTJaJpzKQ3IcZ9WmTIsfKn/fJMY87hIstV5c1eI8lY95Z
878dR4QHACR4PbeKoGQop8PlcPD6GsgsPH+pRJxum0oAX8CAsbIb2fvRHreIRkmK
BXdszVqzZ1b6UPQ+CNOczeJtyKUQUuEvutkAo82YsGrSLUySm6gEVhOdw3RaXkO/
nQdMSkMaXcZx+KTMZf+9gaXlyhqVZJlJ+redxNKUdUbr0SKVobQqFzmTlM/+Wtjt
rKUQjRiCXijuKmvE9xlQ9VgjIfdwbJp6uD7iYDZlE2h0CRTD6EpcW9PF2O1cYr4e
ZumF4I3RSMFqH1F3igacvAIi29wrtovZ4PEeGv2ZuBgf4tsU1TrpRLB5Ptm0gnHF
we7kZifx4fote2mzHmVz3CcI/e1/vTbcpLzgQiD7ECw6DbOdab6gdHViTu/mbluj
9aS5dUsN80NU49tY+3VoMBl4vWNHVvsBfwIZ3P6nyNcRtjbi+MDRofuE/+QWGDkb
UyaOLx1wzPO/IUTIOQuu3hIBTcnWEOEMv0EMPGBteWXTMYVm3W7xcNA1TzdMLsNH
SzKUa4jRPzyDqIIQNi7hFekvsq17Tn1gq80eDfhIc0S/FiNEIVW20JCXfNtC4vy0
SBfshx/2RWJrbxMcV/fE2h21/GsCVWUfU0CrGWqu5hTj242oNiFrFIBM9JFUS2gp
MdMBbSyqH+NXOwfymULeYh0vLblNshIdFWJ+Fw62O6molYdRWUD0FtManzO34Q30
9ngmCldc9REvN/Mq9EnJ5XhfPX+WLlIOAzHWCv7dW8OA1OqNGdBEsnl4QPhDrrtk
QZxX+hqnfjW0KBmFGxWrP4Pp2GnzXIhRqfldwIcwXw0D5pxCB4s9gs78FX26peUN
03zQP/CyXHJCQKXc57/bjxC5aAVVqNPzBzTYSVLrqGRbnoKv8qdjRgfu9JKLnfBd
rI8tERneMKV8aL6dEgr1dktCVJXtIboGAJpQsRTLGL2gZoyXACRHX671ffrX5STK
peRmAT4/viCMsuTAJJuBaazaoldppleuY63+HesIPlrzmLwpZmJH2pq3JpXqeU8R
+YPHvi11hGxD9i3t6HL2BKmpHbpPc9n+/3IfmgqpdQr1xg9SgCg4Qdslzez4USPr
GXJo/JRwdJhccrkYuP+jKH5ee0+Iz12P7kYLtk833ii8L8grgJyXOs3QagmrknJy
jXEMvrm7eoI2sLxCfQCdqAQVlpR3gZgyoUyNrmKgpGbm908nLqWIAvzzKRLnc7tx
CnjVgq4TdTygAMhoxXKfOAssvaAUo61HNwDQaKeziC0gbjNyKHXSd+vCN98tFnct
JzzQ3OFaU8W5n2O0b+VHaAz27dzLM+7dMDp28Y/2rRC9dNLGsPdpv9ZSQZWPTlsQ
EWHY+tWOwfjws91PPO2qPZh3Qx521dI7mVFJKIqygUp0+x8aIrUZ//S8/Kpv84ry
T72PUnyRiwUMUZcNA4tZsgHFP8r+98vzJ/fVaRHWhhHAL1aUPQIJcvBURHgZls7N
jlFUiCSE4x+K+NXir385lZ3eZ/2Jnlv+8WAG3eKGk/sHq1/a9/LyJGhR8TzJ8FWK
CvRJnb9xiVfoLSAVbhA5BGBF1/lWz+Y4b99w8XEmnxlCzJpqk7RQ/CbMidSfwj7b
fi+6lJGlZXY1e8rBWqE04bEbLO04kbkwKiiqkKHT602RcXz3klQxtyOy839E5jO2
jD20ya6xlNjj4j3WxBK824hsnhhBcdMNOLtLtNdbFkcDC5hXXfBbYGPitQ1YYI6u
fIUP6HY0Nh9djWEdU1USPTtoSRyN53mU386YyTFjiDCQ+llxaEtY6z8yQ8fWsCEg
cPvKirCxMpTVIX8J9Tb4REgM7oxUxHX84JSwMvkzNOBce06qDsMPv5Maz+Pachql
wfygfTKI9e7Kc2iRP3woTiG5snfGU5NVg6WqPDAkwpbelwQHOD4lsQWqV/E1S14W
GHKjfKzjXsFf737FASqozMgnHu2DKjtJ/YbnzecsiqRzJ67shRDRSaTdQoHusL2r
rQpgYnqeSVU4KoM9J3B83yKGWl2u0gdfbYIFs/xVa+h/qxxIO2zeMnqfUKeN/kH/
TzQZe3SdmO+/7rahx+sz+4DeyvK+8Fz8Z6vWV/qtYFBbezBfO6BibSQ46lLUYywX
FjTobheGLCFXy6CaK+Phi80wiGsdTYjN7vGxcRymX1TJ6AnelayeYoyCeydixdsD
vv6pdTw/1KeXJGEf2P5aanLo5qW/a7ayi+IMv4F5A9lNe8FxOldq+5VrphjymD5l
PsJV7E58OPuBxCvppM6DTJZ8WYVAFsPr92N/TyiwZLRUSw+TSoLE1m/OkVUW880F
MZ2iMW6kOoOMyFV3ak59hSOeBzMSSk8tNavV/4VdUE2GOCzyq8NZ6lGc/h7Ntaau
BE5cq9KFSc02BHMRAJHL+jOnhTlfhs6mAGA0oWs+nHFcwaBxq4aWsJnfhPTXYkTJ
gqu/tHf+LJqcZ1NSZXM8KzNcZojvL0r/r7to1T0lOddCxQUtsfYnT/npE4LrrBxa
Suzmh6H3iThMkwafkw7OPx+QRGde9RApKQMe/+buUCbPttYL5bsjgK057dl0HwXa
51p7XGvzkUQA8wqHMNqP9qIVDwlj7P5SEurXyRCMfQX9t24xqDGf2JgK/dobM82L
i+VdJtpGA+EXPFg1q3nE8OK8yloZtud+hT10FLjS7WyN2XbWuYw4MaSjhEA1CLJJ
x9L3YejuySeTiTlIhVGKEiY2FTIEYgd3OKa5mjyIj1HsNUbSz6wL731jqWPCrde3
cXBtmSMSCqhiYJ72iNbBUJMMjKt/E4xeJ3PQv7PXvdcnUoBSz8bn7yH7dhYoxZ99
QnsNILf2bQNQhJN1O3XcFWSY9kQkon8wdJjAxk3L53E/vtAMFqt/LA0mYOyfzBF+
1gkew1C1OHYB86CFTxak4L6IFSgpqr9qzC/jcdihDtRewQCxoz8QzBaTzhzHtIYe
tJJjVsvBv3ismbgm7cURARRbdhvNQ9859HGPxYCO8MR+FtoAYAsBP3TQnbzQwxMf
bqSROAaZjfwVXEeXZzlhbpb3D69tBceyycow6LaDqTxoJHZ8nkMREjsr92j5dAKY
St9GtjE1Tsla1+5cBWobOVMtQrDOVB+DdJdZdOecIgXbD1rPD2PWBlmAYucNhf8x
O1oznq0Vfv/XZ6BNo/egPAp9P/Phart9XB4GsnbURRqfTqrV8wTBzfppx9MlV7up
oyps2LMorWoq8rdagup3+Pb5Xpr8gfVja6pV1ISqBQUI+1Xq4xvH2XbFvl55Usn1
rNOptfPKjOUHJyOoNWEE88j0jpZHq5iFtKup2jw4lZmsFi5TKlFN5bbnXE42uXTe
`protect end_protected
