-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ipr/yiVAMMm5+kABrs80fqeERK7Ee1NtkP7+FYc6ybkDrmu2imGtSpZ8esquNpdl
sClG0BRhTKMZHPmCZsDlZZlufRiozXa8/NeD+6Ey4wS9QaChID5rVx2ZmQpoeWmY
dIJLapFQQTNGjL6R6yAVJ11R3ePEDDlv0nc3qZrfCf0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 34416)
`protect data_block
jUurnXbvZ/ZvKo+lq3YBUdfwNwG9pNQCjooAgOgW7VP1EnU5n8tYc+fstG7VD0MW
6WFfi02CTVXXWDSZqTu81pgPm3PxSa18k07yOwL5izfEfJ3WsxQWHlZYYuBmFTgp
L+4LLDdhqL8ZbTh6FWR6ddOb8+bsGnhsNMCzgljNCcWIt8syIJXIynY7wFvbqO1q
SkPQf7OTAuq/o85uDwZjA2gOOD6nUSRjeenCg0AfshARczYGceVYftMcAtridyBV
hTu2QM36lMHf+Gw9R1pHrgAyC1Ra45Hzn07QRDIMaVzYmmuGIr7fkLXRS2etMTlF
ZOQgmYITm8yUhZOMn0bH2xv6cvbkaxiWQyHHv3VqiD2DSf6EcqgGw0gYyvCrYHKD
2hlERCRfT+97+4xois0J+t4KKbvW1ErQocTV0xaYflBygDV3kvUw+59EvHN+LO4b
KJBXK2UGsKipHim/bp+/c6shXzR397+G3eum/ojXISRoX0UyAya1RQG/ZgiPhnyv
BOjaFyhD1+C4awau0eS+pwstz0zv0NBzg4+1A7fyPXdyfTNbXdK6/09vxlasz0qI
oQfimW9xQQ4NhWh/r/xTqeoqXHS4TY6HPy3Oa/S6tJM1MH/c4nVcez/DSvviLAJA
A0S+vIZvdiws+v5B7ftaVGGggJiao4dycG9rhB66DdpZo/gyzjyp9Ovy6Dm001R9
ZrcHNxj04t84ZmVg0HvEUZKsIdDeIhcbMUwTjg6lDzr1BGOqgaAZUL1qxX7+GZfM
dfa8v8+5/526IAPkv0azkRwZKH3pn5AxHngOKxcNNJGuzaQFZaODNbXUccU4+a3q
3zjHbIRgW1CieT8N+87ZWN6PQp1HhzF0mvqX3UOOclB3nHOUlwkIC3b2nPk7AJ7a
DytBsYo7V9cdcWeB4WUPCa3RXeyzKlc0t8I1ynk+958u46qIxSG1WKc/CQtafmaY
qxh/IveLDcuto9ldqnXscvTRemC0dmceueXLRHj+TUISlrV9DS4+epHqH0CS3LAi
ANaFSnUAoKAVzxN8u9uV//LWEV3BhlxSel+0aCrMo+IZOCaMTkx3Nv3KeIyV1veC
xhvjhnUHsIPPeLDYpPQRCFkDI01t5j+69vkMHtGzGj40I+cVIHm8OmYhufJTlO7h
OOrrrFV9AzxYsYTR1ZJrKyXMnZqKjWzq55nNAzXHqDrfPlj7yBk74jfgth4Q0gop
8Hwi7kik6PgTHdfhOGwfbmow0T3YSXAeHaZJsh1Qo5zCw+TFet3zMIol0zlBDI6A
zCmtTr2EmAGtgJZ44Ua6bM+SMNFhJ8/3UsEuDd8WG12lEeANIMuF+FJSYDntHcBQ
e/kZtswXNnViGBJKPA5RAemKA7MEHvEQt5NSvz4aLEOULbOitxnFLtz1ebFE6eZk
+pBOB/MnUf75/g10ltgBeZJXzmYTTFD6KpLvsjLgDBfTtaHnZJ9fhjovrx4mCklT
UvYXgTQwQTvJA5Se9PguUUsOydyozLzmsbuivMqtD1iXnvCtGLvCSR34YhE1lI2O
qcUC/pNQ7s6b6HivEP6AAoT9DPgcHLfNKfpXHpUCSKTTCxPt3d64dC7bYGMuyTIj
YSB4aodnw/Lb/3V5pjuohVukpnzOJQ2UQNhYRb9nDcZN7K5it3IPfkhaPs6Rx4fu
6qyYrZB36j2BCXoMPd5QkPYxKf6Vd7k0tt4m2ZzoP13bY2jxo8u4H5YN0+Oxm2Dg
miTLW5NNEBkNFfWooo3EH2UWbFcnSBAi9e5+SWWJiRz0sIttzpgHnKEaAEFMtk/P
A/8NFZulWF6gdo5oo3sBZhhw6oF6QYe/yQDTWvimNAOeFtPZQssEilP+z2zp5o9E
992ZejAlxYkcoUoBtqOLANboDDP00vPoA1O2WdY0Dp0j5dPcCZP97BrREkpw4OWb
GUWB42MdiVjc/ax8n1o6W/YtK2GJEK6Jw4zwSm0gJuaailHHN8WfxHyJ6maP4P+9
+PHM2w22jW7bd4HzHoau3l7dwlIIXqCiLBeMHwMRigjsyHl7Le7aeCaZRgseji8k
GpyTPsdWcLAxAhhBXe32TxFNLLD+OUxumGB0kRmBHdpPapomPpRCcY0QEq96HZi4
z0U0qOMNeXrj67mt6q7+BcaLAcEFq0HeVKilZUnW0iPZiVpsPOFJqoFr4I3sKkWt
k3mmSdpbjJjsAwEYNrpvVD/uThfq/y2ITFULZmq9rg6mfyQ+Pb7e05oQ+ocIc7SE
FNG4UvQGKFgivSWa+5gIPxJ3mVttSpSVF6v6UCDWlUGPfLBdtFT1HHsADJ8pCrc1
+tI2yvBRgW/IIXTwTaZ0c0REu+Q/Ff66f327jGbFDuSyaX5nlXrZo9KHxYaXOqR8
AjU1lhISPsSyErSdlhE1bR5PvHOd6VBUBNCZhVl0PSiPa8brD9OWLFTveZ7L4Cm/
170dAD7E8GZwnnu92ghDrFd6wfXG5Olh0XIHCN8bxlUF0N8UngDK6vImIksTkbve
7qtLqryq93kkAlTHJGjwOPlImDz3M8lM84WLnD8qzziNo0tam+ojXrNJqwiQh1Aw
qP9p6X1rnOTbAyJEYktp5K/nlLtvxz5GTy+a2NcxAYaQ25SC9Cm0QEsBnt6RROAH
D7jUKNiTWekbblC0M7xYHM8++UWm5W05VzJ1I1yXaP20/VWM5EvrnYqIeUnUXdyu
ERRDLWIYAlj1u770PxjNksETByAZjEjT5GdYwMXKtAfK9PIfvQlxksAR2jkGlz6c
apKoV0U4a+/bdbT8URSRR5sug1csJ36MnjvZXcxMutv7aj9WoAsGMn5fZnpDfqWi
/IOW6NQWoVgDBnapjMDEcQkgdOngHi/iR511qxUz0V2bbniJJFVkz7sBKIg2NLus
AK03NOzOdZm7Pze+xLhWda6nVRYETdCCO9GeoSq5UPuqZRKJ+tcei9LKWdHB/NJN
iJFLnRqzI12ZQaOUgVvIIZfVUsEcXeVTvwd8SPpBt/1I+rr6IIR4G5Xy5PpvSF91
nqV6bMgLa6mWKoU2B3FXSlm7yjMmYv4PAUNOWlG0J8oRBOiVRrqOXcaDqImDCIp5
qX5gRE3SNRWfjRI9scM8AjdsoL1fToeZ2xCz8jkOLzhO4PnVRjxRn/WlNN9pEjZh
TSsAajRXsYYOxETRck2mu1JxEm3TlK6VXmmI2yLMLZWlC8ia9znLqzZUhWgi4n6q
UGfQw7gV97MH7HWv1cdKxoTWS0lD8M/aiM9N79gta5ews7vaKDOAJfuXU9rclO/a
LtSBxCszWekXi3tGRIblXJCrDGV878wLgmIMwMwIi1aA9SLSLtfn2MpxCx+JqTR5
d60xOKdY4VkhBQkmbXBnOjnial53q2CTfWPPCwzqOSp9aZtT2c4nfhyku2s+iMnM
LW7jFZeFATtLemEwc7I09ixLp4RwxO9OVcF2SHf7nuFYpbiXEExg21r+WUxLVFdQ
zlfrIQVLH81crubr6k9A7v7lpCLvz6FgVtVWgh7TEPDMki21n7Pwx31iwEl4YItn
K62KWUPh/56x0y23hhscSocYVGscSGYbD7JRA4dbyqJmfHjFj+uTCZC8LZcbZ1FN
8py/PvU/1cJjHalu7PyJvBNfAidQUThuyEfK1oKjDx5Vf/RybnET2aXS71TLuR86
R3xgQ3fCcNvfjNeIsUJldhL2NMka5aKtjYHmoxuU98YcFZx0ulsjHCz5ZTA3mqWj
JyV0sPcC2uSqmMlEMAccYnU9ynWtInn6t2UH9hNmwko6cHuRTTFHbArJy5zkYy54
KRaGn4ILh4QYOjgd/m3rnM9tG0TA8uYdqETwPji2ysuj2s4zZjBkQegJKLgGBTfw
VSVV3MVL+lhUfYTg5ToVdow1FYOXYl0KYtisTEdW86BN+sEvYxHhyokedRQFLWYT
fLQOcBGYcpajMcxFF2vJNzjcJvarpEcoTfBFsE2QuvOBFFY2tdRD2kffVM1VYVCe
UnmuwydJo8K3jhHY3FhL2SnktTr3zK7SLdHpUvaXT6k4RjeBiXQjuZHZq7cso3JG
OU4W7OuJEY0a2qurtWBMgcShw7t8vebrxmY7Y0o/U48sTELJk8TnxQyWRBzXnMcI
gTd2AA2hbVWMFsJgpCqnPJIZwvhbzPxyDnpT5mwgK6ZfbGYDHtv36N6sdR1w1H2N
w4E7jziCf4dnGt/F0ZRWuwdGy8r8HR1zjJAIjrcj/dW11TTJ7PldqpybxXZocCOl
3XsENstA+znnM6b4KoYTg0i6k3+VQyrA9V6DJmjbQn+SQgIBoKBZyztBkxXsPDo0
7vE8m9gddJMeU7W5cnRf5M9l5OCYKhWpZkNzZQvO7A0ZvAmugWV/UEGwdNWfzplv
dhdT26pmx0ywO6maxvDhPVNBK3vkhU0CSnW5/6LVSMIB511w7IWmkvvZkR1cAXcu
NGBdVowvwkAqyVhcfy+1yEFc1FOq1tWXnOozzN2iXsUQUiKP35D3TBE3br5Hd99C
NjTGuO5kEsYE4pYNVFhxKb7I8hLy9gImGiivNAW5o8USmfBj3+uFYEJEM+cMXVnc
dwoUIeh9LWE2lQsA6jxq6tUS+8yDch6gtb/hu1pt0R3bNRvVFOdrnPVQ3c+iWmVt
iVP1b3kV+uuYRfiOpfM0vVlN5PXHvX6AEC8eQQvgAGMW36WlU4x5jNtKololkcSt
EFNUue2wECKmG09qapay6sLS5jKlJlX8PqOHEa7wcTk/rMrv7xHk/BjGIU5vwFLA
BmspIYkuzxtnaYormzHdqEt0B2NDDCm2OYnhnSNkVRkNlUZfsoTTtti+y7J0Ed2Y
KkxgBIpcsX3qhODhKtMWbMdxlCj6FjYZc6A9/oVjuPx5h3iOuLraA+lZLcZX5XmI
NOUJuteosIuVxDW3g5fdBXhuB6KH9c2lTq7pwP5nVX7x/EVl+brPGh+u5mAmdR6L
62qnPIZw3BDAgglvlQZcUG2Le0x5u3xzgmolWsSnGho82TJxpum6DbTT8Vdq7aB4
lMjAdXX4Gft+Uu0LZ4Id4G8DEurMWbUx4ampcccA2CRVVGl0mcPfkCg69ISAq1P7
lIq4FY4qqDsaBQ92D0m4G31a6ne0n3dusO9qaatEV2hFTrolEBO+gxxZHY/MwwBI
Yhr2BBrp0wwrSJnnoCsEBWKvSWh+oO7566gF1hfaGTbL+isgMJTaIQPGfZbWqP+I
T3zQOhYEpU96iHeDM86R/vHAFEdknKsR0qiu8XUNvraqNgG1Y9O18REn15vxt7kK
FClZ/QCmeXT0b4HWQKwT8lz4U8gawZj/vTRUzKvqMeEKANPVgGND1DZnlBLTIMXR
iWILB5xGWtyonyG8cOgaW/Tqv9C/YflRk6+2lOhHdi5mZS6QUoBzmMPI0FJiGTM5
1syHTog2piLW3qcJPTXMNioQ5Xxb7U28qO1TfQlIXy7BGtUWrM6j5+3NnSL9Sjfb
JYPnZZz8XsfVLTbOCaSseiJpFhAfo/4VbK9bOB4glVKJKOn4GyXoq3HTCbmq8QVK
+Hg6+0hBj0JJSuPYrIOIDVKE7ohVkBWwnA6dp4Fbx7yEMA1iOgYDHmixmXS0AZjh
asSpTCtt+Dbx17v267pIPHKwOzblgpMTTyUA9WpN485405LuHF37qF/1BF6m1IZU
WJJnN/W2fT40f0MGt4hueLYgOw5OKvkCidzyIn2s4pvHhT6iMjG4YnEYb4zNg/nw
QTlywtKoz9Oju8N6beXv9r8cn+kkYuXjVbhUav49bI96mkvIxrqpNu2A62frR2i1
rlavbZEXNgbkhE8PzoUzs/EOR7WY5o88B8XzicJFelWO2a0p/t8OPl+QMV42h5sw
6zsq/yChO4mGBQeM73Tf9WK0yX+iIn6ktqZBS0anXZdwWNLpJcbn2UKxNqn63ce3
Ei6p5QcEQFTwx7rJ4+QZiOyRSeSwTLN8GqA+EXvpHSLr9/ZT1tBcAekpNV9RLW9B
XCEeNgh4dpXJ7Cgbe/eg61Ehw7AjQQBvn4+ijbAhFsz2SuQFC9/89Tavm2k0HmZU
+j4SMt/dtT7plcvmTUVuWIWvsneb3dzpVXhrz7dSmzAVz1KSRkJp0V3dt/phkk00
fbelEU0rhv3BOIIWph+aiG/VQvJwUaT2kAW9b15N9Rrp28DopBn9RAvvp5mU0LQV
xyyXmLSye3SVobezTtppt7vphwNxcvRpZaoIdd8mlqzdqYIabilQSDLDifDnOES1
0LpBa6geAlEkKxrAixQCQbBCT2Zmzv3V2reUeRHf9EUbbaXh6eyxV0nF+QVUXRXm
yctuELg+imGROSCn/WbQ+0yp+zehUT19+ZD8v9nkXNSgJFlwdkPZEzGiDnZC38hy
p2e7t34LoaYf9o7M++EYKmZX/+nF38gKgRMD1FIxLxTVcP/v3CX52irwT+4lgBp+
PcXtqVIaAkGISNOGFwGzOGPtB2HpchiVdgYAIh0KYkDiSfk+KLaeuNhNzErl7suV
Xk92uraIE842ANwdK0LmCw3UZ7dGirhm/cZoYwVWKdnz/n9Q/Y1HIFBeTM/QtQmy
LnwbHVHuWIE7G38UfhTq8Hj2iF8BxcKqtXbUNDQOlHDGi38/JKFrvpRDkjsZbEmQ
eYxemXzdepIYY22kdEJvquFCpQM9JLkhV6djZmGT8HHy0PmabqVTXu9kBoa+kpzU
uoezgp5JwhQkesxlQszl78P/bfGdHOWwJTuo5/9F5y7eBKolFJ06Iohn+P6MTHCH
s1HG9NNmgqiq7EG0chp8NiICjBw1F+RXFjVJTa5fYFH789x/3U+0XKNfZ9MrJd8P
rv6hrjdr5aNa+iyoYzfs6uX+izXS43R2SXI0pmoCuQs+Z4fgdgktbn0/7brdNc1H
yetpsbopJTs+CARkXU0cUPd+qSsGu4YWTEp7D9m4shqEYabT4QZHAkYNsTREw1oN
AFjIJ0PDcNQuWgSIrNG8QHds9pZHXh6vytcYVBGLNKbr56QSk5ELHYKapijvjtiJ
5v5g9BUU8ip87FLyT0hdZKvkpr/np8lksZmpn6J3Ic/wDogcf1/YvtHVp8TpRzrT
m8lUssRacfVXPbzZJ8OdG/9VjOJANli7q3wIrXbPk7853T4K594K/4chTmpOC+1n
cEW4A507pEy1HHgkvRPCJkeIONwsiN6XEtqJDJAFSxA0O9hyI7thr3KM9TbyAiKc
pxOk9MdBQ6jys0gOPU0WHj/XI6qfapcIUD9vjfgY12/318/6PwLsPW3eTRRgPyaG
qkm4dgofzw3Wrbk1WXiJ7BNGspCNpBk4YhEKD9kxj14mc5Ool/HHMh+e0laNIK91
Rq532QiHXkQf7ugsE+tk/Olj/1zaUUyIbDa8yVkIMkmmrKnVSPWMJlKp/bXU8yql
u56XsfVNlT9RfjOurUIltezmdWE5P6938LHrxYD7fnGrfADbtrSvjAKWnd3xvvEw
G2Clv3EEJOeJuf/dI3FW0ANBdUSvUoirz5rUTGoVo8I5gBKPoJkzVeDmqR7iGjf6
Vio6AJuU1J4+3Sj5D0rmkoTqfe2MGG8YTuZAumbETvCdjY2smbH7b2fBHTlkj4wK
OzYgkjTzstJaXQBt65YOJMNcbKRaXjAcLZFIdevFT20wQzHSEN6eO46/yxcSKVNq
Cz/nt9FhhomwDvVXRW199Wi7TZJNSHqB94l24GH4xaN9/5xmIkQFl+DfWHfnSDfF
ljF0HpAIKlyQBnzocDt4oFhrnnN3CIsgxQpiB+bNA6QyqK2VqhpCu49rMaKm4PN9
s6VH0xZ7J0x+Ugw5qSOaZKwRiB+fTGMpIrsFuSH4FoJMEGII/bki0WQl9/rajBOf
UczxHhxpuHsz8f0M9b2mWvYZNogbiA9vfpDhRCEbvy4B1+f2GWoYN+U+vQzzvwuY
jVWNRSI/xbTbAHmcMxzQLHMB1Lcgrl2Brvsu4cWGS5GTKZAxYV4a6ByNplwMUIxh
BEn6Op5ZkUmFNmKib1G8xHIpIGXF/AAzqA496M4ulGGCC51W+3kjjatm1eVk7rXH
wIPMAJHXhaESB4vxDL5j6r5C0p+qBScta7d+6qy9hAB1Qfxqzk0KPxeu0jRjOn7P
PE/sFdd0Kkf7S50dmwyJpTmt9NIAieawBAn/erI9WbSw3IfJAktNnbi/StGMpbWY
aKO8C/SP+o2Ns2IEqCe8UJYvKuWP1Kp2mIb8AqOXzKsS7/IieVoB4eyHkBixAcHN
1v+YzkWrWA7mMpvMjJyOKAaWHGwB0SGoJ52TSmGJPAbIcaOIdl5vFZdVQwoQ51uk
mVuvUr0sq/xjPGcpKwfkgaiQ4n/o752DZVKnNDvqXAp1/W6FtARVtHKciZA/ptEU
9MN4t3hFoLnPXRFNx3Xx/Hr9SD8KKZpJDMKtdSlFjxG9Hix2YtQQdcUPxJpc0xZZ
ukwiC0su4O+BHfWvBaqWeI82RsGshZd19g4cAzsyz/Sud1taCcmLSUtX69iQM9AU
9K13kqbwx+7umuti68kZ3a1x0Mi58OIJ5wUU6r+6oS6dpkDNNq4vO0r3gmok1oJF
9yhPYQmXMGdPYd/nSnPxosChYdOuTLqZrYhd4e39E2mphaYNl72SANqQDQhP8vE4
91jXqe07uude2NfIGdujSYOgazlLQDLIcgzwO9ga8sayEAIRwI3OxRBroxWh7yhu
udx+9Tbz3uPL5nXNaqXdI4EpCb2DBfGAeBGXaC9jneP0kSCLIPJMAH068k3wHXcp
cA86WJUahASNaUzcwuNxgj7Hcsqkv9n2Rjx4OtYrznFopl9CQrUYSFOyLrItiZ/k
9F3mrSTULgHER7HGZZ2bwpNKw6RvAzxkY4YQzIu5+d4h0vrxdsRkPnLVCK/b7xVL
w7o99mIVvm4L6T3gWtOwjRXnCwr0aczQR7FG8bkrGR1MaKrpHRkDuHxFZdwEh1yn
YOoHPdgCeBqp5YogQejvw8PfaVz10U1CjBmRXr/1MY+eKM4DupMz3enY3vdM7rEv
GvVhD9wIB9h+Bu3ubPTsPns/2vdhG/VVN97NM+/iAQ9tjFDm4ywhLx7vhvk+EMxm
/WVo0pzU7Ogx9gKqt5rEpT+GPsaXkGhpfrxINcDS8ortFQaFBWvn93wh21plZYKU
QnSD056WzMLBbTAkXAUo16LrPTuzy0vDRzj8x5UPZ+WyvbXwsj9wn4w3okfQX8aN
xg//rv/cT+onPc2dWKe4ahMqd19qeiwYVWTbFUCTc8VX+KWod5XMMScucfP9awYJ
1jsIGjfQ5E95Kj2Z5Z53O8zmKv9RP3QAJd/6GC9scM7YWBOK/AgdoiS4MQc6uK7A
3eg3BdvaUHXF/cFKILm41dCaL6eSjhr59WcqSVBGZVPIGHFQ4QzlHuIGMryaCvIW
UAROgU/IzWEGscsZSVUeK6tUiKhsvIJRcAeQi7QZ1jHgtey4kPfSba23eKzjhEnQ
zgVy3Av1QToW9In36TZzglvU1+B74nPDNBkYVL/73oR4fppnWBFMXR61dGuAKdQ7
r9URPvmgRxyhv4Gr8JQcYfMIFg7WnOinwQvwTwRWhCM5JGb8aazgXUzHDpXQx2P9
ache3yBmN357ukuepmPyPsT0LoV5/7Vuus0QOhtfK/18v4iBl1dV7GPnfDu0Y7ap
f5GOQ3pj2udMHGXDgS8A/vUYlVHXxutZyh+zzGRAsPew9IEkKjAoeIGe62rqWMCD
XEoJwe985Zm7xG6P4LRlunZjGq4iUhURxEkxuzCqXwz6pDIa7kc7u36irBOkvt8t
+2NIrS/6yEHQaMHO8ADipeqjp2tvy/J9l9yC+tfkcfpS6yNR3pUsk9iDqI0m4Nqd
LAt/qBD5Q1LBHSefUlFOhm3p6AaZbPfcc/xJ8WzV6NbWQI/XH626aFvlvrfb1IKK
vUMEt1DhajwixykmxH2//XRV/DjgvM+yYs11nRXzu3Pyp81p162to1m4eXgSes81
2ge0VQKE5/HFmvybjOY4Vt2YuC+hpbj/D8IxeqbwpADmc7+O5RzNpZOx12Zctb0Z
J7UfSMdfb2QLsfKHMPfAsqSZH3CHWCgl21xQyFtwhmWfPftVfjdWX8no/uVrlcFk
qMa2bz54l0FH6Hjdio69sDted3t64HSPxF3AYHWGjSuJpb2bmdnFNFtKwfvHmzzN
hGLNKLuyvUEH+e2uCx8E1kVi3sAinpfdjiTSG0acqAVpUrlYoPKxxUfzuhVx3ubi
aXqIVCdtq8zW2ibqFdgN+f5rdPGPC7n7FmZwyEzjJeBU65YJbUsphAH1WnOeRAoJ
Zzt8QWmI5nmyyc2EsvJg/1ichAbZg/555Ob8voiwz9Z1oTUqOr8gMhXqYaIqff2E
4TJmmvrIUhrpydaythtYfMkhj8C2e81X0aXgiWQH25DdmIh1OsTlnIyTBofblrUg
DKokHm0BK9ywidcnEHkMtZ8eJF/E3zXvAAm9e8ihtdTkSDfA7O2r03SAUMkQrA3p
bOGCzXLhLpUU8g+M72JyFoqlFMxzSJoM5Q8NNJqbwdD1pcsWLrrheFEiX6MGYjYb
/XhkBRDeNzXbFVqoBWV20C+oCRer04jFT4YC/FMBnGuzyEFLm5TjEmR/TdMFmF19
EEmH4qF7Pz+FfRIL2+g6srE8adrfVHy7SFsR7GWkVKpJt+6ZMPrcRWhROFLasPBb
bOyzwB343n8ly6UsBHdMlQS9pNVsrZ04jz11Grws6ENchMOZB67cnTCHPykVjytI
QpoAJY8PxIn6iCTEM9fnT27BQ6RLMLN8muEBskw0IuMlZZpAjr229yKSRXoD9wSb
Csz9EvJmYZ5TDHOvdTTRtEPEY+7oiTROsYJkyU6Q4luM8SZJMcQVkvjJ9i8Ect2r
m+ych8JZh44bWGbfH23ygifPqbaQutZ3clxWZ/Ts8QIyMWjFG3sOblpwtXS7rL33
kYyWsWxr4HLjzmVTSsaJWxnq8M0IHbmHugYgYs7jlN3D3ns4d5wu9buIxGk1DVbi
rLi+H93my/HyAr0z6RXN4aCbBFJ0hkanZ+w2okrQZ3TEqGJrkPI/GDGtBpClGXbz
ElAhLGWUS0m5FeJt7tm+IguN0Hqr7SUwlZZtJNBmVob229jIDzAAWZBUjEymWteS
VMivygPUQaR5Qynf+EOjapVrA62jSbCAsrTKZJ5xpFvVQ40/fDMe2rE2UEhXkvH0
pWX9yVZdjhu1ayqb51uqyUVLJN4sVvyA/xbSK4Z3XPv1mQ6BNYt5D+f0ZkY67Ckz
2LLWMZBV9AhlGn4wBQY0Bo8N5sYz6AwQjhZVQz4WkuQP4drztVygyEtpE6x5VsfG
SaFD0YQTfutbaNnGnwXJqr4ELCQTMBs9aDyQkhutl61hNO4lSR3H2suCYVcdjNfR
z+NwNwJ+86tLsV3s7GL6A3TfEn8DGs8bLJXwiskBTUAIuS/u9yY0zJKpiKIT5riJ
utPaTzkTDCSvN3GU3xRMNUorqgwEVXJqG4dJ1Nsmy33WbYP+NlBuVsOMPfg8RuNp
neSUv8i1XzcAcZsy5+4ozPN9weReXVFTAylmowGFXguvkbO6k1Cr3JnEd0XyEVmM
H/Sp3XqP6z14gHORUUpiI+ThGqw6fgXDyg6b5ljVmQrX3+i19sI5PGFMRgzy6kQ6
9ILyjFoFvJSTBNxAumA/uSB9eBI3rGZML1QeaKU3GmDdp3H74CLSAgvji5FinK+F
bO/rtGQwlhIEMSmYM6lu0Q+Y/1srlXO0fp5OChv1Vezwf62ANmy0jh/WdUKe3whb
haIXB6UEr6iW9vJk8/LQN/pNaYmkbmFav8hZJ6aXMmTQHz5FdI6xsb0IEvJUqSUz
bPLULT/dHZ4Wt736Vzlacz5oGLSNFLjlImiHR7CEQx5f4lnwbTNh/RIGuyrWuXNm
0GWBo2Qoc4Huw/Jwt2jC7aNz0/FToljaJbHVaKLbuSxOZTGf5EFP/cw3fOCyykVO
4dw7X9doGv3fCfAsKfOiOVs6BaQPgrVKOhTX16OVlH9RUSqA6UJS4wT5A9V00woU
YctAsg5l74N1FV+ayA/Sm/kTQTxZVUY1kL01oe5Y6Km2DdcQiEg2UvcjsC7f51jP
OFNZdoQiAWmzQJsJLFptGJmOtMm/cu8EKENhKDfn+L/ghaPbZpZfBnTiwxs/XXzI
rMzfX+O816FpNqzLH3Kv+B+AGfU1O9nVptgCYb7P4pkCw+NMWgccEm2Jq8G6gCdL
y4Oq6uXETq0GEiNusC3JpjcpiWG8OLwG2Uyt4VUFuKL3icwDnVewAwBtborWa9u+
DTS33v7/iJhvwCKiF35E9AKmRfRChxQ866GDbk+OE1NGCT665SISDCY7nc90CwYK
otjXSUbc+SV8T7h+st3kb8skXPD/OYZ8R8Dz6l7HhCQ9mDeuwErcXrHQdevqmI00
umSZ2JmNRFVMBwENSYYyKshb7DfBq1MiAS5URymgVreNYmPgu/wGDKj0MVCVYzS2
onxr2DF5dNG4heIc7GO1z4spKxMmL0gHa4UetbF1OLk+W6txh+yGK9h9jcqqZPA3
5gqJn5B0thuls75NxQqIlJMIkY81vZLYl0h0FC0ENt0wrnpQh16bfS4mRkeyiOYg
ICplSieADWZJQ1hlQIi4D8elEFdjggzcCnGB9UcB6KZ+K2grFm78Maos7cLti1tZ
t0mjLeU66ZOXQ4K52nP7++NKve5fezUWLvOrIC4UBHIvQQkfEhmxpGR8wYlpyfmS
dp9KA0ttdw4oVMMzmodax/qxhyBxai5TsGZVs76g9K2jpj4Cob9CX27to/TUVXHI
XbTORj5PfVL+Vg3UhP9yOTAmeKZkQzkEv7eRi6Yy0ld7Zkw4MJbt7PDw1indQxgg
R6EA1u0l2O0VRCM1PSeJbI1VZIhJwupMEsTXk+t6OADrt4Zt3g3kzsioQB1imlPz
lAgcyNZhnlEqqbHTxUcw3vpfIOYiOCvvicth9bdMVC5ZWcwQo3P+kVfT/A9D1mlh
rCg4ODOlQFhsScDoTpqJMqCKcmCUzJHrm0pAqqmxhm1v2Vw7YVmHl7idk/4MXOkn
KVrK1Upzh/6/VY7J/di38QoF6XFLwZfGL7RKTwIoOHcsffLAro13Ce7MzjswN6Q+
lJJAt7tw0OMmoVXqvbfr3oC8GiEiP4V9rS1Dkf96jrz3ym5WlYNChkwGbKsOG9M1
aUm1awWLn/Ap6a4u7W09C8JasgJjgMLjnw5vG3ku862McyDjGfEoaHqQE2+Nw4fA
GYgm0wW2nPWR2DwtLkXliWaBhJThllVO8ntJErL5UI03V2Ji5XMbUnM3wgZqPmWu
wzklhb1PIC0+Iiz56M886+9t85KNBtNjZ7wg7MAxcaqdnnuCinDhBACx5ugrnDcp
PRdZFd4Jjy+9wjygWWroa4TAhVz0OBqaOaio7/hQU3F2Q5xtbdLYKa+YZRkvLJnR
BP8JwMXIKCsBSInOZ+ohXAVsZ//Xn0n4P74ez01m8x48a1pVGAxA7S+jwR4yUy3Z
zEZtTb+PAHiGTZkmH5Gx3TNDqvdu1Sfe/uSrpLmNGPhPrg6ZjbOxH5Wfq1rV4srk
dn8jITcxHI2e76ALsCXHdA9Hr4cWZgAkYbwxCg7lRjyCO7oEQm1e6nFkC6j3UsY5
AcqVJilIOYbE1umdiEdhwZck1/qkzTxQfbPFwqKXqMV5DZTZDwqlFj1/5+Styl6B
OgH8NcGu3XohQJ6zmvzgeBEiEa5KEszX1UXK8AtmG8oQ9LXV2c2Dy0HD1oOflios
qQswU/Lg8xPNrBwOALcmWro8EeZQ1Nmma0xGq67EvNC1zdhUGTO8Svo35D4NqaOe
mydzrOH4ZAAqZ3+RN6KF9JZzQTARowB5aFxJ3RCiJaOxN3MN+fkpeayy48NPQScN
QsOJCnzZotVKzU4dg00WZpxqhPD+R77PJBN+R6NKA+Tlq4LGSA8jbHEGbTygw5wX
ZIZZoGkHkcyLxPGzi70CFA/y5eQjTiiGxitKkeLGgkuf+53iA6iHVWUrYJVgliie
aOzDE5xSLR/NU4GAiRhb1W4yRpCDMmEwHMycAi7zMT/MCy3C++qOT3rWp0xmsjPU
SRnUir8lzQgpkvUCeu897Ly1kXdCrPpL9k53Xugr4mnzJBARSvzhG8WiSXQwA3e1
aAxXWmUGgCc2vFXQQ9dWPDAfpIXo3zjYBYgHynq/m+kUaNHNRbrW4eUXqUu+kXbK
wAzPmVOjbsUI90mxcNPWYxk6VQm6U5Pg41UG7YWvq80GCUGyn6uansedpP29u42B
30wNBFBnjdscLC+1Ckg4QS56iD3M8ggu4LAq0TmnNUA7e1dAp2e6go7bDXJQ9WAN
HlELHx81aGMqW6xG2+gc6arlMOux745c4NCVGAI/3h4/IbQW8dGG6VVuM7juKG+h
SuzxlcGT6rQWAzB8W22Sd7DlFt3AjZQ9PG+zFOvF0cYY6UIFIXqEGp6kyqkjKo5z
g8Sia7fDdtYIuC9Z/giGnXqlHnszVrr1z1Z4sBQIpXfkiXLHc322NNbVX+v7VzXJ
uui7aKYtboXJnd4tzKvoVovKqEJiNQ2XtGNr6aXSKUaE+ad1Bp8ffJXxDxypr9d8
2WV1KFny5oW2RrqjFRoLOURPqeTodHg7m9pYMnTypuIyU/8/UUDP4exQtUY6bvr8
UbiG2ruUlPRNVYvLJ+yBxJ0MK8K3FbdW2G4ZGlYBvfMee7qgtTx3PXR7qV8dHWVh
hJKcnjlFcBmwvCIalh864rW0jhgE9LTvC6cBBRv+qRvilfli3+LLVadn+7oLpz7C
IDPOk1hAogyn0lfUf1irW7JjAQzhftc26MS6EMb1zCVxl2J7Vjl7MUQIhf894NaO
pYyeoyrDHRnnt5N52jqwQUrV/njgimQAov5CBxX1dO1P9CgNOwhLaCuoAKtB2ewz
cZPpAqGtZNuCF4ZBYBJ/n4PzcmT+o6t2zTXsQrOPQQX+ZgoyRjHFOhwqmLfiB4tD
5BD2vw7QKYZ9S5z11V6GcGljetu9FWcfSMhyadROkbTf1FRp8Rjsk+lhNkvqOfsN
mCWWWoYcAtVgiv1AMmv2BQZwAWtQ9ywKJEUpwgZN4nBULTEPwlPD8W6H/9ivhyvL
PPxu6nG5f5bOyQmktVtsYBk0sBr+UdX/Z98GtoYFPiDvD84Uszw9nT440h+lxhAh
pOJ1HWhafv8ynV/2pSZ0gJG4FZvEyC4j7ZAYs2W2UsX5AgYLby0B8jHVTD+Roduf
3hQsQQY4hRfwk5g3J2F+ZPYMmfrjl4QHgNJ6f+axdhqRwRpd1WndhCtFoZAo9dpu
cj5+bCPypSDIAUXoz91OtegJkpFU+5Mb2cTTBQjc15LpJmv5Nntk8ndnMSuby2aE
O0G5kqgT6SIFIyiMl5ML0+N4iovuRHD8QvrvWs31CLZQK5BbzJmTRv7/J7YK0MfM
4lt5/KPeEHGWNFcSSKV175G/mF5R05Dxuswrfq2xwrhEhzvEgZ3slmsa5tqqfkoY
4NrCOa4KWXwTaGLuSg75XfcScoRnM/fM3UbI4vPnWaeGJ7TnGNjKrUEa5nV2FsbG
/abKNc6aYC//Aepht8lnqgziMzfTsP7ryqkMMpqAXbLuxVjHf/yzZ9fWMtjoiw+K
d76Z13OzuNTimKRh7/8dwADQdT50DRXlV73mevC4qO882NgLsDYBxMNwVF5MeXQw
QkF0ezZVTewxd+i8ldDWZrNAjecpGzlF0YSZfQ0vhZNr2UySoIDIMZz4rcfpUpoF
Hb+fvWrW42X046XPtd5YCSOYMDbNehgEjtt+1zvunWYSeV5uo5k1ZVGdyO2pYgJa
to1pUcLtwFEQdDxmVBnXm4IZZFsswKQTVFvUfGytXgGoutiTVz7hR7zDs/o1yr97
JePjtlCH9WV4ozbuJD6uK0OWCbgCRd805LvSooSPc6uWZMRZcQ5KH66pCYLOUJcO
x8ldFrXGkG3M0r4X/+/xgqWPmFVoM2IIT/9lFUjuqanFtIhpIvMjA52iwcoqq3rr
xR+Ntbf4mdxepuxHB4OFeQWBlPWmStb87jjgGKC5dkh+YjjOygvXYy5H2faX+YvQ
URH4twbgOjbMkbpWHJX6wRmf03+iJYUxP89E6cALAqaNWEdRu4RMpeLy32HW0eLX
/cjzeeh+ujJHnNNq1ifIxulTfKPwjqyjJrUuiVKeNRQj68Atx6MVSrnPpdnRz6Ao
3OU0t+FjR0bmYRDIYO/r8olvw9LgVlWWTvbK9edY+Z0+hZ2ttQPKtgsa681lZbBX
zRziYV6PaPBppkBAl2FS9o/8HetRj6suun3wqakPomk4pPHR3vmNn3XLtssmL2xR
o1bxZ9XclwtcR8dMjX0XrsErRAccj3ALJf4GLx9dmYdTcaZNUBQXC2sL1yf6B3si
B7uhLusNewfZDUuAabnDYu//rNvBw9AFOOTpiWFAGTsU4Az399MD+mHwsRQF+su8
nMO/yDdfzpoGmxVUMNlJ5TN98ja+dhQYP/6t4NwKPm0fwTVxt2QPs2ZcyfPS2/Nh
PM2hTJmtYNkCX2JdeZwAsHEF8spdoyJuvgjxSi8lP/Q3kfqLrkxu4rNH4UVDnD5Q
ngLFtefQJzfHwkqrY3THTlIPv1ezR4COX6qwZ1pXsJA91eH6KKEOnh8EyGyCnKQ2
fa/Prlsyy+zP9a+cpAMKchcQCf6RkvwbZj0vWYGf5BGCzq8b8lbxdhGMw+dtX2Df
wg36Xbesx/PvsSwSllnOAfN1dDgosm3hpK+J2MebYpDULex4+wL4bObyPf4ys0k/
heeNTESp/WGMcSHgtFCemLcqsxo8MpcspnszIoSKMiqCj6bBuiu2pakhz1tHTdBa
1xxUzKoYM7A4KuL9vwr91l1WXV1NMCBHq5KAlsVOuipTR+bVR5vYsEtyypwRaOTj
kz3scMMlMpvb2fVYMh+gTfEW8WHZrbMBYDbPQ6yBtPTSHF8Yh3wvk8BTLtdeKM2g
oPAbdSNd71kWLgSXuRziPIzLurv5chhmpb6iF6YLwyZfPFYH1wnopylYC5JQi3Oh
aDECB1Yf9yqSaBQerPlNN5qTeu/oRqhrf3UI/1t+FlL0mxx9AZ/xqMRAWMgNzTEo
wqXZiq7L7FwgYy2qG08l3o3WOF/At1aKELMxJUz6i9zbfhTDMV9TCRIWy7pG4eg8
z3mKL77l5Liutgtn8BLq+wPLh0V8Ic8sKh1s6b9ap97dnFp3dmPJnGgn0fc1kI+V
uXbksrfBbSSiX0NGRsWkXO2lNCouIb2WDcr+l0nK1Ft2oJbvunp8Y0CQTLnxnPcV
OvZv1oVQPDyiOTj//7i8+kLUCr6CgkYRWOcgwGd2RsLdpDgZTSFUBOv629QIfwqN
Dktdo7imEFyJHhEsqbB4Gu09hCnHU6TqBLBF8PrpMmBO1dcAbJilhP7tZJuIizEj
3zWVmYS0TRFowneRkBVRzSZGS3mG6uuDUS/PpI4H9lrymtKrhGvd1zQHCrmDQ5CB
alf2qmhLIACaxMB9tkHyahdLx93Cf+g/APt/NZk/IiazozRIxSuWPKm0wUYzU2fB
B3qOnw+TQIA/b14D1qXpXyjZRtlT5CohujuC5XSVx3gPSBjfpI1hN5T5ny8taBb8
MWespj++CwPxNjZSxHTmVA6ZRUAU7RC1fj6Dp1friy8i+5x8g6gJgixCUyZSXSTg
lAwozraPIS05f7k1Wvv8G1fIE5NSKTHJCQFRe/XK+L0SdT2eUD//5bkG9strcF/f
3U9c/pe/N1ZeGzoIeg9QtJx/ggpDBZHeNt4wjQaefFlmsRQQXVaQC/ADWublm9gi
aTZqdiagcGonH4MspuI4AkW2eeV+uGQAmUUWujvtSpboQ9KD3r9KeiAKFnxRG7u7
XyaPM2rjfk+GJALTpYlIn+c3jgURqGmVHgEoXutz++4luyB1MCYEnvqDpKw1aLP+
ba2PDbzh5hDbZajguPwjnCjcwvkEAzOkW6Ek8CiZHo7AiWaXQc0NDTVJQP5jgX+Z
boHUGAk+oHuj/5aep5wvGcgKEmGpJaCaVpCjk8kqlaU0UfD2P2l40SRZTqaFGVCa
NUA3rIRDDpZqPlO2E43RYExZHT/e54n0Kh1xK07aLQsrYtJI4ElZXiMSgQ555OZA
8FoBsoXqc950SudsIVd5ogm2n1l6iS+U+lo00fudimo3sktO2CuJ8iyAp7IKEoJY
ZsZ8X8H+nUFG/4G4PQ3YZoP+qtqhQ4yNlVlvdKC3Jn3UiEgC7/sNniD3fiu5HTFp
+auqzlpqngKbyfArLOoCxkN0cbIcU/lp/DGyGPI+B3HerOyHbFBDEPw3Yzr+d9wp
1XLKorsgM3Eo4b3yK9pcj64yZl6wEAyGT2AtWIkMzXdX/FD9DFKk6JNupcgIaMqO
gwrBiedFwfaTncoZY9iDVuw7jvnSBLin6TYAwgK3lr45B5SreZoMW12f8FpYcPEC
mGYPrRDqHreRBaOQpzwa7D0IOeOXhkiBDHeVkORSZ9b94ItGy1AmA6jiTae0uYeb
hhq4MMsRcqSs+Q9TfO/HDfKMkeOfIUzyBR3sunlNfVU23mSPrNL1gOACjccf7Olt
7OikUVHiZ1FNGZR9hY22vYGyrpYwRxW0hVzFe6ks/GHl7P2Xoz6+JeP22VOynleQ
HlyY2Gn/+VJxF7F3W/iaowAkSCuEWFu4J2BxV0Mrd3xk1uIs0ShhSusEgBYPiQX+
Cmg8udXy0ttnj12uphdv1o5wp9V69YGXuUDEuzNJWmgUZS/PByhiTum0DeVspuSc
8nxfSXEFPDX+5XfhwsFLeqB2il6TtbczRPpac3HCcX1gbUwIajnArbXVsST1UEUa
D6WENuzK13vqLZes45a+0abP6muIklOpby1IeAW5LlyaGKYg65r5yd46EjnofW41
+gKZqEbHN93XqqzbPDIrUzVpfY2ktLRCG1ksYbcQ5uXnoCcGuteZthsMnH9+06du
0Atig9UAQH+rEJ7ZpwVu9G5M/5IHbA/BQkur2/e8PdNV5+hpP1jjeHbRIt9VCc0y
5MsdThkAKSShiXExyzFulQh0oBBusgF6UzsvIbllZNTU9oAeYKhRE512XyD+gh55
MdMhCkTnBjeInXbDHaFJfIrKTMQwoGijvJEQM+Ye9HOnwobgkXTeZKDHOv1k7KS8
Z3A6pJc7Slpy0k/x1irhR0fCWCktLWbQNP5QImmMRH+N95r0So4usEFWVZK2NEOE
N44HH3ZorROX2aFgz2Yw0W/izxBmM4ZEg915+LBtATNetMRa72ZzTlmK+T63mDH8
eUz3X/nXfvYkZF/imQeM+Uhj8zuMyj0Hhul0pxmS+qSjIq9CYcVlu7M/5DBugmcw
wnWe6k3liS2aUqplWveJPKMSR/Bua+YowIcZxnNGiwNLXVA7gn2QtTRm18KXsLTi
44ThYq38wENNjp9j/zpLt+KWv/zsMOQxIXOR6cOyz0oJe8AdHIZnAsrfEmAjxG8X
BffAbybMOg9pIkofTLFnevYItd7T3JqYDiwKg75srVfO449Rd//YqH6SUEiBhkRd
Hf5QwLFX9GtfhFdgi93onTQGt+3n41wENyjT0WzpPl2FoTZ8Q4ppeXEJL6VMJef/
o7/eS2e4Zzh6MBcLJeF74A3MEe4L27NMdODaXVa+jmab0uh4TNIej7HGLqYkQkXw
STJh+UiFOvFgXgh1CMx+OI0cpHIQU3Vj9VIb8FIt8fTGuz1uTuQGfLmseU3B1/Z+
Cs96/SEUdrZ40eC1wiiCHQei2yvGquFYTarXGThgNLLemOUElpM5GS6tkU4SxdG+
r3llB3VSbVq6YVz2zz6t3qmpuqAOgF68YxQk+S/iy4W0aXrEvQUqfBzoBO4yyUsL
H2D/Lfi5ov6cNXsL+kfdG4E6XzvgfXIEO5M03V2XCeVgsJFS04lQktWihQqsuNiY
upgJtontaTsxdqPgpK7pjM57KATP9BswsUSSgbEX1om3QB8KOfvvStbx/pFDYu+f
9kYDag12MCsn3ZpMNXgyfcl69gzlVXFj7IeBOPDiKMSeamYjGrmeTHpXxcNAQQHF
Xcgnon82senjmB0eHm+/6iBA6wr5OxeAsB2yHSQUzOadI8jY5SAaGpqv+NBZZnGQ
6xAL9ZBukhcOXqkZuwXwAiQJEpa29rl01KwluX0fMXX1I3ohrSKNzwbNLphdtFT3
dPyBs9zpHjheF+F2l5fJnFzhvfKd13aNMZbbCtUagXrkhPOkhG9c+TdouTmdtsxD
7q4LV16iVTSuM4VTICWuUqWwpLp4+vkXxOGY43KGpPpLd0K6FV6mPjwRJoZqf6E/
g3lANxZS1C80BKKNjEG8hqYPVmMQxYbm5rvZ8jcKpuGcHovCteLclwRgDaqtIoKX
LC4EF0evGkV/5VDJGLczQbgw96/zSyqLkZj85hRC11tZKLCID6uJW3d2Nbfant2Y
+/jwarHheXUD0nUq9YbSdvHBnLetSZO5KCiFxLrSe3P3qn+aATdk2bEDZTHKw5+r
48PxMnhnS+jd4xKTPWtXnSDLmobYYharijscmnKztCzFQo2VssmTTrS8mVJq0j/o
QwnIhMgSWFbovwHlbfr6qc8pqs/wl1vc/dTHcffb+95MWN7Hrb+PMchHaiN7BDf7
oZPSbcVX2ZjSV3YZzCr2VIdJVtx7qvenf6nGeNMnr0SeCrnfitbDtqlwavQPhh3n
ScztAhkKqFfQrH6mDBhzIQp7FO0qAyIyCXw9tPhkhYrwoXoKCDFxd4aS2oInrQkB
l9YMr+YuGal11yUuX5VnDWKkyL2PuqznQJM+islBqGV9MLXalg1F/eNnzztV2GcF
tr7kEXF6nTiaWQjTT6Jr4vhw/eAsK2onLNTRRY5G0cupDjUa50IuZsd9gd9dUKD/
IpmI0/wCvW4xxw7rKaJJ8YadAFL5u0QAF0twxpXus+weZsStkjIBtMbDGE4Z7Vd+
8/CeJP2GXnGedBEBViKxb+21XafsfT2E1FbywPhbzSnpY71e9zTv9gmVWsMBcm8y
7PIwAl7f69FeUSAKYnJjNZMTy2b6TpVY+LrruYH6I9Vhl6sjUN3hc8aVfmwr0en/
U+/qlJ0FgqTMxk+gTsF0+puA8BwEc2TZpwIaL4TA9SGnYr1BwFe0EJIKgNk70ZqP
s1U2bgsgopoHzt+l5/oydsD0FpJvGjjBaUDrPoaS2XsCBiohBp463ndijFBfKQ0K
MzXx/2otNvYmA9Gc62GjEkvN8n7hiitB0ocQ4oXrFA/YinNwv6yYGNdDca1xvRXz
E1rzhEdcy1tdyh8SpcYM4Ej1hJ6YCaLS6PLPsugI2Jtx8i9qVwEfyt6Lzzpmw4Gk
qQ16kpV7zuFWenNgIthgcx0BCTpEbM1v1YmW/KeJFxeBrQi6v/F9v6KxURDlr5MQ
lC3GOa4MO51fOk3c7dZhmyjO4hQsMOoREmKZL91g7inNGn2riWnRmieV8hnSPWpD
mDvcFDf66STqh3dAeO93hiETlHkI+m3UMPXoYV7tLxDW4EOdbMR7U2AGcn1qOM/W
Jb/pW+lyjhnOdc5eU25D7zIVHRO+GJ4Fz7wwwFYy09ZP510kGFjamL3FNOJnF4Sz
3PeDlnclpQ5yOzjE9fb5xIW4h39u1Jj4/orVlS1wP5JHAp695lsNGXwDcoJKA0JN
0+2yK6zO+VDG/W3kdIWvAPDIejbpaSRNtdRE/RBoxq5rNQRQZNim7pjU1ZKaGCHE
3dJX0YGp+cIOhRPTduhCAz5aZJI0r/8LI8QPcdTCEaHUu3LOzMwMSA4aVO7ECdX3
qhU9f+y0BjeKENurMM75X7DNL8dho5oCm5af51oXUijuR719we/YxNxtDlystQds
veQAoL48XFfWvUB7NhRqatc0CIibS245SjEk6le2KDAMqPGzkCH7cbZR1EUnFx6X
jjr0w5avuYaL2vmG+1mplr9inNuwyWGSV1XewLz5lAddlewZbPHc7YcfJXPpfkUJ
M8OIagunBrgASXht3VTMd0iU2Si3FozUPPApRHRTITPqJqcqTAnKwSw/rG45fpOR
SQ1EOfWVKDTManz68NJNd/pRIlfYhxO987JA9c1L+0F6Kd13wfTjsa4m27kF05tb
oPBEP5IcMWXfBpp2G4qrNKE93cIJ5Iqj6SYVTgOunM4Fi0S41qa64MhRABE9eucP
8lDBg45RjQgeKoNSOfhCjgimBnup5Qwvv+dZodmb09se75jkU0TQkoHdGYiSqpGA
UGq+dtsKGU7D0RLFjjUAInoVnP8K2CUW7gVFjlQ4w4D2GK2CZFCMKFE/Fayc+G+n
9/LrGzISE8ROEnHquXaj6eJgr1W0huWxCO72Huswsb86HDS1bLFGI8nhyMeXfxCK
aHgwOs/hmteoCQxzBHyT/1SI+mpnFdm27yuhzd2Mybnz/Kj+0GPWf+2csQjQ46Vy
z7UvPWXKUi5L5meiWOtCDPEWdhA0FZk9nIWl8nK2opm4EXAuFB6Yh5Dn89yodAId
1XLAS6qUKn6RNFM8c744wxJNhpZdeHaCESXUfBiI0upQl9P0TedOy7Drvv8uXs40
E7DqN1DTP2tS0UYa7KUHs3gOtEFxBpRbgqX5w9dE/XNE8eIUXJMggd/NbeiEsF/y
jRgoe7t9fAdoTaOiPth8eDFDqyAgdATfTLzLl7/NsWEEbP/VBopPiYTrpAGwdZeV
PF0KRfwr6UhwA9kaed2xA0HfmSwM3T69j+qdv/aKOaFTaliBakJFaYN5VpVB80Ao
ans2LGuCOxlRc4B10KL5w+hLPk+QHV4sXEuPvH5G/GJQDf5fRTkrAuPjF99NZjcn
uX0jJtD2jfBOXSdZ40/EuODaaqU5yC8+UKSpf4M+jSTIBFPtNbAbWHA86mj5rJRY
jfrD9vaHDP+XahOyyxnqJSgad9F1ua4LsGuHMnXmBKuMytPGucQsgzg+tBDMdQFQ
Po5yu6ak+NYrWY72I2mXzdGXiJaKD5A5qTwLxWtWSD/KFiJ9y15eWIE+M52QNvyh
FuC3Bi0a7ekx61kLJf9g7FDTL192Y0wa5U4ywEu5aogUBPcSXB0DLSwzudhi+IJp
wD9YPAtS9eCED889xIUViBoyFOxwEi8htzYwji+XplDysB0nE3viv+PlM5omM8Yx
TmAsWF0aWTcvuYzbMY9RYSmRA/HbQzG54jZWubgrxAvZxQo0aFzOMp0cO6YgFBWL
M49xsBbsrN6EqJ8qjFCyDf7TmQfe4Dhx2kuu0NUW++i6dub/PT2OVs6NgPqtDcE0
pVDqpPo0NMwtWAs5ipKr0ABkl/YTQ2Ungvm6dG0Pg2FpwB75j+D7RbN85nGXylJ5
DmF7XIygJRDloYuTKHiSqa1sSeyRR4BujOz8mIATiuz7dWQKHokr0SkPL+buaM2y
YIwdyciQlFEYuOOpYL1mtQQP+GnA/QmZX6sj8wTG8H348C0xSGSJV0fi/Bim9SeB
QVSMVZ3h8pOT+e5X0Ks/80JZ5UZXyVbwH2tp6vDExN06Eb/m90IWZcSxhZV7UsQ8
ia0JRqOK494LIdf78+UzNhWMFZg6Dhb0GTrsWHZ7WD0kHv71/0hz0a9KJwugSeS2
4LuhML8QOFTWeM/jkoYh27GihXrv8BbzfCiMtKe+6V/TH1TtGoFgXesavwfEEKr3
OPcJr8i9ddP7KFVDI4e6z4R5Q12ZOifkn/55y+HuS6q/0gMBk+4f95WxBTwbUC21
ZUVnMvnMtbwA6Os717K3P/3BS4aTMV/yI+JnBA5ttIaJeul1p5rQG8VD4Amuy4Ah
PF7Ydp3R9Bhs6LnNiXhWj/4bST9fdN9wWfr6AF7VEYuXhRykJqWM65I0ElCr/x7q
heR+oqg+Pvu2zryLsF0hOQ3vG6kMoLOdDi2QkHF9hr33oZcM7BPWMxyeJb8M/0E9
xASCvArcGN5Ky2cCbE29SLijO7RGoIs//blUCEM5/70zWVR3cVcZGVbee+n9EOjn
SfDSTewFXUs37iTRx83wCIzanV1fKAd5+paqfC3MVkxT7E62QPJHBtsQ72InO8KE
NPdUQ4aJFE+sZYx8wrFM9jT3w+06ZATmkH3omeMzBzdBLBmkZ5DTVF7fP+Fkw2eB
OXqSDZFU9N10DVlwVlCQ13BdjcfSRfwjXjx4SBs9fbF+GwNq9tl2mDJnw37iOxAd
Yn7Qn+HpdJ7bQuEkordtdTWiHtUQStSmBFWAKdOynrERd+0cJJb3yiifmhLvhE2F
zwBhK/+URtdEadzr/15YLZTFoXxBhxjYPTBJ7a+GEEGdOjWYFcEyQ4acfWzIDO57
8bE7eT+oxjhq9NrbKzM+II64lXxDrxUMYH72Pft6wx6GncCt6Q3waQgFL4XFNSkq
/95n9GWqX+tggd4jGtE8ru/Aeu+ybqT1qUTGapp7p+rPxc41ZBsv4ix7qIzR9U8X
lpjr8RrTmvYglcTD504UyHdowR1Tg8rZanILjHqXjuptNcRPD/VZxSJrpiGzwTAi
YJn4EFc/Sqw20nbGh/xpHehEt1vTECaR3Xze/B/QTiMotwo5YWxxL6Y1sq9Z3I5K
TSz8Lv15PWozyK0zgP45P8ICyfj3GIFnT28zWBO36uibCavYeD1Uixf8R903uT6g
+bI3z6/Z6WCLpq5wXr54nvqR0/pjQw1TMk1MdgLZHrj/6b8K3e5eWNpOVfkbtCcU
/Bd5K/LGFyEcnB0Gd1FP2sRhjJbeMUpkp6P7Rk2Wv1LuYfF7js1kVELbvb6A+icq
Uw3yYZ7ytgvDbJ7R4nMfDfCI9K/QwFUJ0MH+O8nRnHfMA6/m83VgOC/zLx1UQ3F+
WgdYJIa6eMGtBxnVO5MagOY3icvf2XcvB9TuJL7YWldu/OVcBWBuEnshduwXi5/Z
bMSyotzVfOycqghHvJ0oFy4E7NxeP6FI3QGFaEKYBFAe1mqdARXKyPBarMOeiGwB
igdsv3qeKOAwZ3KL/PM6VXSkAFDriz+9AQ+05sRnBPKrkPz2VXR9kDn3Cv9jyQ5H
FaxkAWpSCYMxYXUHcDWORTMH/MTqYrLNmmCysLwnLkNNbWtdfA8zckR+Zrwf4MOg
e9xthIkfE/J6OJtmxvkZZHel+lA/nZc344DiAWmNToeJSm2/upB/6wPKjmPRiXIS
UzqPfY9eBQ87xDXQfjTezeqdZmeuVfjeSC8WOB4etjLLVOO5ZDDIWWA/7jyA8HPH
tIzdLPlX2mpPWNHLl5w97dZTXiRNor5F7WTeLHmB8kC+kvxyNsg88hhT0F8uw7i7
HC4oKhu3fBjTUXQMnRcb38CRPAmvZzDYGn95IlAjZz5+EY7KUXMTpnilZNxeGxQS
mlN7A4uTeeH8TnXGoMk9TfSTPZ07WxcYTUJJgBH0AZrH6TaIBVb0o1OATP0Y28U5
YrCbafcmPPsiN58KGPxZwT6OD/jOGEmr5q7rLvxjk3U5BTOTNtCJOQf8ObzBJzYF
2o6e6QzZjTChXYm2lTs5Px/zFr+fXdSSCskvZLmmL4Byq+38pXfYTs4w5RgyXZqK
A9sGDb3uATgLszMcmfvM9v8iWwiLmLEF/zfhsz48UTKvZK6aWJxjJtTNNIBgXqst
8Ok60tusMvsDUDYx+Df5atOlUelkB0H6xP6Qa1UkbH4xpL5qyZiylKyKhIuy4nEm
3PZZyx2wyaKCLFhNzhWJD2O5mEPxH7TxCoc1XrP0aYLZzRLTv1ZO2y0MlaXr9GF3
sqhNQa19J9un2A7lofNbN5Z9J9auI0fJZv+zDqBiZZ00IXvRjZtv596zQQkrlJR6
Qn2d7pyv+ETgdhDQicorqzvrkepF59vBQX6IFOWsxFXY3Iuyo6rqhfHchLJTQ9oI
XlEWh/calpcuWa8yHkJw/cr/GocdtwTvwuXh40GxAXO4xi9tZ3rxtWBG1ImINeU5
ki3HffXtPinsC1xAC1vm+qX8AcCWjmiJRrcrKSFpy7olSuVZaafubaNR9SgqIz/V
GABi08c00Enxv/TLFp0cnfrAFdHFEb6KNVrDLwhHVCpPGKX3VpM2twJDTnloAGSk
O2TGfFcwhx1zWul7pX+F/YDUv2u+OUuC23IHwVyG9Z0dZbLDZztJMCr8cgO3Rgmn
DA6YRwMXz2cA9pgWPcWALIJ8g+3Pa4r47WhGqhQyUv00TC8oJJVp8toi/y0OmF3T
T1dDe+eeHLKGrzHFEByvoqoC2AE7qLf50deMBrIHbXwNvwMPEvLjbMoXUrJKhLOV
zOfotMxy/ZCiFxGAjTL4XDyKj7PvDhG3c9e0yUdCjAjrgniHtce8zVm2azoGpY7l
gMjd6dG63xvTOnN6PVXyWaPVLOlj000WYOqod2Ue2BBTG+xZYA1+sqQLj4qhrrrZ
NMxYxiCFaKEFyE5Sqh6Y3626rCQb3ypPDSPnhKkYXkMG1OG0KWJhnPxgsAXWlxcK
gzbAWSujlx0MXEk35yYnzCNYhQolCYRlWIO9l+s4/e/rUUIBedqWCIXROh0D8/2D
juwHeZ6J76crMCke1FEdwpTziWMGxVu9S9BmMtW8XpuXj47FAz9BptkhUq69TsVr
hKCYKxGGPzt+33T0fni931jUr+RhoxR6OTCGCbzHET2IpXMqsdBfDVIxupkl3t96
1MWvl8Wi6aanjp9Mxu7MRqdTjFVcEBX5/aJIdf/kioxEdI+9RVvsYH+WmWPTUJtJ
5EfzEJc5oA+WJUetBrxLCg8ipEvycedF7yZW6eJp+ztwegiZuXiDaQfP9j1NdUGe
doTjXnXH/81JVVh0qMdvmvR59r1lkSwmpjFzSTzp993khFf38FkJxiMN5een3k+m
WrKFAAbhofdLP28GK6gZGYFUiWuY6aSJS9TBSZN58AEmeJloJ1EUyz4E3/DapRwE
WG1Pq+GkEm5jW9cyrvs2aQ26/AsRsv9RlG8i3njP9LCgf2tc/HSsd3kTx3FlDZix
s9Una8+9QgnCfZlsYe2JLos8/ZV7dIKxgpf9Wbs6Z0Omtdly6d7QSdV49gFxFNE5
nCWjfeNpVonFhpgZulCDYnV33M2wfnzhWQYuYkosgtp64DdI6u4MlPqwZ7cBF2HC
vnmLSpg/MdICN5e0F6mU6eGua6MnHs0ZNpjUF2Xul56VkmdWJksxLK9M3x0YKmwe
p3YYxQxZUsUi1BkjuhsCDXmWpB+IQDFoSe5epsBakDsd5LeeCjTtCxBw4j+lEK2y
MCpRw1SsBLk7NNk/pVwb8FdaWKRQE1s3GeGfLrM+w7Qtc/+t1ydtPLFGZWYBKAT2
JGGkkf+Dv41uajiusMUtys1NpLnSQBAGBAMNoMum5tguePlze4jELtlR8ATQ8PBd
XQQ9S4Cn4CjeSEtYGGJlbGZxk5V5JbuwSsVfOo7C0MaGbfN/2O+fn70pKY6BTpDG
MJ0hRe4+I29gqJo+52w3X1Ch310R2t6azF+JNSZPEkWoU3b9fDWcV7i2Q8jZaapR
WY0a17zZcmmvOYjylNNF0FPNGFG/JRp/xVSb7VUH1sGdGyXMeaEMq90sdIwOMLT/
oglDcqujvN1vllWxHiVWKMwFIYVlFJpT7cNmeFSehOMdxeEEZoFSV9cwr9KBsUx7
wQ1hqbX7lkz9iAjJrl1azyQCC3jokjy01BK1muaF/BKI06eSSJtYWnzQxAX3CKJf
1ijr1U10FitwPDD37nqSxxVR8AkennXlhIJuQC++r7ilPamCjF5ZJQRwtvHyjNSL
n0SlD/RCsfduEZUGkAdffGZiw0yEjLnpG0P3aWHSsFE5YUs6l5Tyao1veYMA1BQi
Hv6kpGrHLpNBx81wbHNZ/j1x5SUQGj0HIjqJ9kSb8QsOqFKJGXNaurkI+jbTK1zq
SK6H+amrxFwk9FBhXxFoINLw9XrmxO7A5QR42kq+0nrbB8FCwDXL00ENiRStEUcD
HQJpl4JBsUzAdp1Ea2n1zYxvvD9hEPkVOzkTPOD8xgdEloQ6Dd+sOPgz4QMZaxGU
8iPRLzZYabYva5RJy/uBl1Ki/TzHUZ4+UIA5dIuupHaB93xFLuXm6cpSGQCa6opg
0O9SRw+SYwxg+fqteuH935EGLvlnzKn1Ccnxs36kq2DFF8AEslUS+xHfWZmd5Eqc
oS5VRbM4KfFiPcfDr+JrX8xNIbW5FJHV2nlwS3gg+w4asrCL7XYcgAE9iEQBQjoo
NuOJOqNajYJy9k1rNL7SrAhmbNe5M1CKTS7qoFN56B8FY+ueOR5A4a5Qz/w2WjTJ
AwbNOhrToN2XJc5LyrlDuD1/Fns9V4l2WomZrrqe50x+0EYzIipqPPu/1GPl9O7d
S421IZbN1tY8AMdtw2hivIbTcZK2t1ep/S4chodPu2WgywB6xkjmF6TkEG2PZVmW
ne7ABOuCrqsEcx/vH1/zpC+RJXjmBA+sDLBGpCNJybE9mbOkKy7fNOBuVoW1D8VR
3e0C6xClgnK4bAul8/MrJsnLV8qmkUUAUtgUf0cdd8tW+CrMgTbOVwtx7+K59MqY
nTC7XANhfdGVNj/5E8bj02HPmpkH0tXTE5wT3eDkRwR4yrISzcVMnRpRz/ky5Z0x
c7Ut5vswkkEwoJXCXkNT21RCsT8rdxXGWqdAolYhhpgZv53xzpkwysZU7V2ZAv2K
EqiNsFPPPMTWY7hxfn6c2JRKVMFOXvtIDT7Qry1IrBocV4mRsC0SAkgjj45pXZKf
dSQXAOFN4IOdoj3c1n80xXhnyBtgwIJLspdhUZy9cqLMH8MmAAAO3bZjIpzbmWEm
FeddyI7wM/pNqznrAuJelF/zLr2PBVwDuGZZGpJapwojulj6nQFvQDwQJA6srg0g
MypmoHjjTi+uqkQnhqLy3xDKH3kwa4Ez7QdyU8zup/o08MnQE+/4a14jgz7uiA8D
SdmRbOfDaE4OzYdNBvGlULm7/86Fe3lYQMuhC3AARiaUsEMl+J0bVnRoU3dlEwQV
P6Q+Cjd0BScYXDsd/chQw3jZhcuIbna0/YgvLCKcSD8meGUD12HV84rQMXa5g644
vNtNuhjQTIynI2tkUOAbAmJWkqFxvdjs3S4kfbew71ViBn/jJdqCXy+qhFATomCP
KKhsFbb/KTknZwanR2n8EY/k3dGcyHGFZKN9xG0ONyz0WeEyng4GUSRLnim4wnFS
WmGY/0GVq1lAx53OVv9tGjBuRRcolgExXUBxIRdlzSKKHCOz0fDmrQVdJ8vSmF1U
2tHsjATDN5wRARPjGgC6RxRPHxt88eaR/+3eUVHQ6QfBAPHZ4Ioa5TzjSllLofgL
GgbNMmQy1nNzydw1hRM/Stlm8/h50jp6O1PLAwwW4hWFjsIdHjI9b8evrOI0Or3z
SlsbH97zA9xb9/Koo/Mo4QPdYbYdmvgCWxtNoOsz5QEB+0DIVo0Anym0ThzGg3T1
GzvJ4rk2wP+eb492bUXw6Ff4K60YrEL7HtkSfhKtPhC8FvQcwoFhlQ6D+jJS3lky
p60dGPwpA+oQ9QNZfmpy0vcGQp5aduHDk/x9tNPXptNOWdK8yTQdtDr6vDSzWAIb
s2/4iRjA2f35xNE2nywQ9iSbVXg8Sps3xxTnXdfYDk+L5awDAY0LYHOKbXEPcX8Z
WP8hvBkvmcOwHekllOEb9uNRCzZtrFQs+jNmkKqPfIOiDQrJEYqHllZ2f1B04UzP
iDalhmfBjG//GTQv/mR9VJO9/fYL20mf1MT+IPtHjmM/r9buBBkKdSwUJbHnV/df
o+tcvispEltNmns0ja4W7obDZt4j24m/Ke8irWgiTic5OGcjzWc8rzkeT0mehkvf
n8GFCxwzAYD1AcGT2LoCADUF2BZe9n8tAfeOMQrphhw+WmW9xXKc6O8V6zY/txiy
rlS0T+Q+r0UQJuawk9JHYkl0VyExKTdj5EOvAKq73uBIKUkfwa2EtaH2WGv5Y+TA
C5oVkd9ehZvQ0U/ViwLSJDSC+BhzHyKBQS0WjPW7iWw44hxpFRLvyS0zXyGAxETn
VFTXZZD44K73QErIkkbChgrHls96MzbHaKHZ+/cPsXY2Z1A6fjuCI7U2zzxouLj0
9X9LKI7VHV/dbtakiTR81360xn43JSsCnUFX+nJJ30SiK5vOga5INOgGerdVVWlm
77B929VP7k4W68pDSIKYVNY/OuFGWPAeuVPdJnk7/AAVC2jdhV0UVtCxxzgVvvpF
gcv4B3DCYPInmy0xJI6rmA1w3G/ewrpKHc/ZwL5osZDBP3XFXxAja25x9aGVAmeG
PAgKOX34x/vL2DSYRbeK5yuDb1HtM+zaeLwnV5dXLb+hfv8R+k+r7iXnYFWiCxp8
wwxgIx52tb/vVttElhnOoVoXnLqOYdtjXipnHcbCzfEh7BcK79mkfQ8oDRLKGgNO
EH4OGs7UuxHoceBxMrCDk8f3S2G+W5p/3jdIPb3s2hlR4xpwln9aVab10EM1fc44
HnVkk0XFo+PWy+aNeqH71ShT7YKTXzF9Pikl3lShq6BqZq1eBOL1XUAOjJnc/Cq4
OMbzny40zZtyen36oSua4sG8E4MTAcwC+yf0QhbVUYrY/q2hHyJwVGECS5MSfHfW
DUtO5oBeJjiIcT998nAMcONEeCEvCAVViewJkTCqgOpm3K0Pi5ZXteEMpu8Zfy46
ZUZEO5G4qUIC+EsqMQt/myn30/t8qi4OsgAj6FVAd830Ml9mPUzloKOQtjip5y5C
IqQmE6WwKEg4IB6IWGDeF96quXTcT+penZZ+20E+B8TicxIHFU1mm2KIHnC3Q7cC
nVGrw8nECPmap5v+Cg+WN1mqVSH7DSxtfN5VSwuNZaG1Os6aCTbKRpjFTQj3ChMs
A5exfk5c91Ge6st5zDjoVc3fzv+tMmczJkNdKUyxD1DMe++HVyZVgf2S/pqh3uHS
8OQ0zps8UZtivtgxtGDeqBNyfQld1sxzlKLr2orwGX8ByXI5eQAaOQltliYgrket
0rz4a5hNy0wus2nEBi9V9X7TI8lYCSWIV0/kNCSvyva1rs3Evn2yH3caLEbM65Uw
z7DHPTR5aV+bMBceBdWYS3BqRslJPzL5ITbLFveCVDuNo1os4u82wYSPIgY70GRU
8BOr1AqH5DYw6d36ziCjvtxjrKIvb2OJfMGrFw7ciODuzXAfoTbQdpQSVRWsT4/J
51uxoifCMKHyBiOjHNdkO7CeeG3s36pHvBJXOPSsMDAIXWCk/xQjavNPQ2lhIk/k
8hP1y8KlBoqKYgdv7ZSDS03u4znrbeMKIHFV1dqYaMBU2/RUpIkW/E/6ChKhFOHE
F2Bx2MCg1V1ARZLda5U+g+3IG/W1W4cX8u6wpo340fv7ygP3VEByi8YzYFI3z99g
IEUMouERNeZmJ2JNC1PmglAp7jb+bk49tZen2MZFKYv6DdhTiKHslO7p4CnI4Zgc
If1532LBDMln5rq7uyq+T63DZLbnJDfom54pRE2oLSPW//1DPdwfYiGZ8oHxEAFx
aV8ePsqX7RMfsQ5ow9bnyviHLwqVos1nss48zCEwcmPEwfazSpR5dedtflAgtgjD
YguAd/A2wKid+PUxtxn4ND+hZJFti1u3vAlt5GUU22ubztx/e5ObnY6RLE3QSgU8
YMCQrvsSgXef20xZcEeRL8u+pMecdT4XM01ZG5f/x0iuIAg7YzbkPHZ4yVDqb/Rz
3xc5Zk5/447e6NhybF4IAjvuxUHXubU9hW3ZiyXGr1rZXzwaGYcSTwMudGmhvw5H
hEddqvDORNRDTIMWDhNAE9kfTwpYcL3b2adFO6OhLVyUahJHFS95FLuUItxPgW7M
0Emq+1EuPFELnBnDHtw4qJSPJ6xRKxRqigY+W+yY4MQqPzonELn64u4uHPcpYx/I
CpJE0CcHhlAHJlqSUcl/I6erO3xpUyFIujN2EtgVBxGNsS7LRvOOmQlTQuCE5O1J
iHldVHKAyrFM600enaPbmyQMyfQaAdWOVdDufo8+e0g0Ys1hmAh1fwlt4MKf6BA2
JO+BHaQ/er+vmd52we6Tj6dQDNM7xGqTzNk1MqE0TYclmUDGy9rVMRW4B8jkkVci
9cts+yHdgU/PSKDA9f3vEta6nQrRaV2qZAlbBnkhw3oqgkSVUyey6RgSZuwinWqq
YVJlRKsNRFVcLnXsh0/Vz/XUozHKDOW93AmN0x6SVaIZIFSunMuMxfE97FnIuPcZ
pLDpz5U5FW2TB2IXAX+GistBhquTqlTUltquFSvPqyjNGWtNcXSGO/rNe5f1X3aN
dCRxfs3sc1T5WHtAeClRfhKyhfOj+IIbg2Zi9eqANT4cyu6M0HDZ6Kbnu4waViRf
zJViENrSt667hAGxC0ZPP2dB5+S75SLHBh32Nd+51wAPuazNqAAmS8Ozedq4T+WW
J1pn2mOSS1eMBmo9arKLhAkKSOK62ah2BUyZYOSrMRyMJzKH5LsKaQgMRbxTUFKT
N5mdIkczoLGvo3BlBs+WOrA4ZWwxX5WeeB4C+JMkeWWNqewRwa5Yny6v1T7NPx6t
RlchtxyoSznvt8JwmVYxnxJlWc+0UZrpxzb8MgT0KHlbFyXDZox5WMRRNtu+YE+w
c+3whqGrADIz9kjGlUvQ0Sdhj4VW4PfVOpChxqVmFdWNLYHW2bn9TGdoqCY1EcIX
w4RBw9ZPYsXv8aSBI5lRI62QdMBsX2PPtgmB0WehMotUVKabbqVS3mBVdQdJrqUj
yZt6uDRO3LQ8RLMytVkMWpBh3nadowPqRIUvPUBATeUrcwNj4kC0RKMLNcg6sAiu
8pMOhoGJOlRAaOTKthiaxlJRv9Ll/CnUVggLf21b6PwNO/jPEMtrbWM9F8L/kcSJ
MUoiMvKVQWolC244J9p+DNgStHGGU+56zXcFAPrJIVIN82yLInoooLdcNlB1ojLf
C9DWGYZNCNBPUNLX4XhYI9bEYJZVTULSh7/AjMrzR2zcsCdZw8R4niPwjbOkOgT4
jtbvxgaIoxUBQzNOd1oIBr40gbzLij4qiZl0RtXHYuBMqgrBorLA1QODRCnfE4d9
hv6qCo1mgmvtyqa0VThke+X7AMRDvnhFpbVeRt1utKPUjSBKFXTNXz5HdpH1PQSm
lnKcVREtPpG4Q6H2C4GP29IsHtAHtcGoNamSBmbrZq4ZVX9jB7wx34Z7X0oI9WqX
p1P9M5KtJi19XmYafYOGcUo44DDv/9dhsaL3AWAt9PsBdTmhfVxNC30TC1GCeHJJ
qlMYXyKk+QKLPDrzuIgJ1/FtYVMr6Cir1V7PkXxmTKhUQ8bqADSpoHBgthjjZr51
HswQ3uOBQAwv+GXn6uOMKdYvJmbAZ0EVurv0f0AZtsQc/IviwPxdCe5u1rHA6jYb
9tYJo8dnYAScKf/BYhB8eSpl/hBTjjN99fPeQvYajYnFsgys7S0E96nZXjq2BhMM
za1iBZ71c6TN5+tNpHQvwMlIje97GQv86Ift/FD6eawovjGpyXUXxqoXU7SIPxR7
QFFIJ+mFnLRFJpDiBRgrvEYYUhATzw0c9lcbox+a8hlwNeWXirzcjuG8ksSyZ2GW
Rr/MpGAm8Epuzjbm577u47bJo7LvNfG4vv5edJ+ksl7ZkkL/96VwVUMGJpZt7tSW
h9jznU1PLQrmk5kG/cDDyqvOatZsAh9acrqirK/IRedyv1AP3KNow+/3F1UtdFkK
mB9xiYd6C2x6WpIdYEBA0XkXkBYPdvIngeCg69v2hDrMwRO+TvVtePQ7IKnhAMqg
VS5wd7H0vG42iZQcSPprT/tMdPY1xl1BQi6Pj2l07tOHvB+g9kO/bmDo5zW42gzr
dXAsO9Csss72G9h9qAMf6sGok7u8FSC2bLq/VhRKwYJ/yBQeegQ32pgCXObSCtH0
9sS7afa0gztOtHWk4/0io89vLcOPJMf7MP1FZaUtWQI4vbVNa1Y4L3YLFya5ZzID
PLvls+b3LTjLI3YPR0WDE5gbZ+7pysbXmaQBw8hWndUs2D95IWno/jWdimFDvPsM
Im01x/LRbEky9fBVgaQI+glRMsel31nVG8/J1LUGepU1NtsW9t/dC/sOVt6bvrXO
PeTu/9XBRgWgUEZmkLwqZYO160DSnnImIMb7UKtMetfh9IIWs+lLYRW/1duMJlmD
QABaZ/XSwc43em/fFIk33P1pVuZJzGBeS/QQxfpTa7g1OgnK+aHc2YvjZnvj6iV9
er4iGveYsgia83eGSpewWIWvCv3YX2+LsjDtdOyY3r/NiaMD5yuvkYq7oiOOytAd
z1YiitqLhtdvl82AimxkeDpESbC/X9fYV4/vNjt5CJ6TJPc0r4jZc6G+XqlQyecl
Wonghtz1QddquJyNyPURxN1yDSmrucqmfMMXglf+wxWoo6IikxwBrtfGg+3DIAQA
JI8abB1lzjXwGfdbSjD27wViXJxhoJGRysnAr15WqEUJJ8E9TwsMd4HpsNaowMAd
DtPxe8OxLGJHKPxcNzTEHa9S7s3p2eVkBwqgIDhpxkVjwjLN2qLB8Y6m++oWdwq1
qbBW1u9mcX6Z9jAPjXeogJqBOg8HuTFspmcFSjYgql+206Yeu+hVIXlbgyRpj7u0
omVnI6PJJe+HZ5cZLAkavaKB8MKzqlWC7eds/pcj/14eyfakJd14BmYn2Inb1RbB
kBC43bcnC73miM3rA7H+d02qTthOMosxdCjUVmXDv9impP9IPPup4m6kMktQEjMu
e1Ukgr3GYCbsjRHKL2AO7L/pU2cJvbQFkhX1337bFqjFBk+U9OB11mMzAtsIM5Db
GxSdiq/ZDlEC3gDBA3Cbq4ihkYLE8UAUv0t7GMmnOIaOtkJkKvB86u5Fta/Qx3Bj
lA87p+kDUK/om08JpqcUUlR3S2D2cegfdqTDuju0CSTvp4KI5Y2UROADpErWHM5y
1tHIk8d4g55wD8cwa9nq+345oVL8yss6yyMI4hywOboyi2cHXxrXaK4ziSBwpP/z
ppCN+o2CA5YykawVkOJUXQf9bmDL+ITLFmmdvkj5Ap5CCXaS/uLw1bc/J18dGfX8
UPoqYM/wC2u1XPplkgEk/LUx6c/WdELPuw9bCrBGrtfuJh0xvTgdQLP+u0U1/qbU
JD/YM/tKa84qNGmdYJeUS3QA5CkGcyfmO7VTejjLcXOZsVRX/AQUoODGynlm35np
LGhacKSPwTDY0TIN/FoDJhJ15FretuTjD1+alk8yEnszSNZFqkV5dn2RJTrmDsqm
sJWaHiREMTZL27LDmcmWZ4XYWhxwp1YG3OxDAbpPCmzJrlyKRS9f9/+pD0swlA7z
TLjj3i0DgKDREPFmGDHROGRWsoZOO5/2pz/T4J+25HKqQEzbIsmkPplafd9vxdDL
thUnp7Uzg74brPRWpl9LRgDG+B8icVS69ex5yfvLfIYl0Fm1ed4YqLu3ksDjVRvH
H2NvYIqPtuQ7+kLvJFL16mmMqHuqz6Tq/p5fn4LO1KUbOn5fjfnH7M/MZjYqb30z
JMY7tnz16cjVdJTH+glUCZYtDPENJ8Z8jaRULCjs1H3ibwWbPvuv/Oniu1osFc6z
1n+XGdr6MVHSEifXVN1NjYB9dlaUp93chsb0T++OzrsjTmCi7Bdr4+tvmrPrEcQO
nKENgWtCL8x7cF+6K/6pCjUs6ovES/3+Kd2jWw6a7rcxYUlyS7S7wY5cc6G/Xejn
1CCjVHKsNh4QzIlIhJml8UQ5aKtkBVlBUeXenLVAcLBK3wO21afa+Y7b36t74+N8
OpROeIxB9iU/VeKU8q7DcISI92ZTjBP88BQ+10ijfybINr8KLQXBeHjyiaff5kDD
hLg64tHbQDHIpvoQ0fAiczOY+EP/3v8hkcy+YaAZ6Rd+KtXR8v7XV0sjEKU1ovV1
S+hb+6onkRbpKaY81dfaAA5uWOmoQ//XUHhWFelEPB8pkRpgxojgQpooTL6zjc/Y
Wxbuk089heetnoi86hzGYJjyHpyzrgf/xiVNYwcvWtssNsVehYMXrZXn/NENb1Jr
0n+27sLjCe4KGZus7nPExQjgGrY5GftU9DIeueZnpaG0m3Bedc2sQy3tzFi1qCqT
1dR2iUbcexsZqa+mSTsL9V0fSSFxaIZ370jZXRVYOER3wpPH8S0BmFghE98Igv2Z
hVRScqY2ZqHCoPIzIZxf0wXlAqSZbB/w+Bj/267T1vQYMEHOBFXbMzYuCWmuDjI+
RcGnqKF+Z4EnvTYaOq39gTgmtCVYh51I+a1piOKLDmyXKvsq9LfERn2bfzfTACO9
owJ5FnLaVNMh7G+v7YarM7l7oaXT1BIjgpJYMyHfRLF2fzWTieNHG90h5va3rHQj
cW7EFrjTtU67OmNS4zKtRSqfTsry9EJTy8U4aMMzcyzx9TeM3C27wd/M7NWrF+Rw
TbdCg5US6PQoSX01+g2XFpJFtbDyjE2AiBEOPWJfEao7flBMHmAj3s7zWejtQNqx
qVWEV+ldAMWqMWTNHro0PpS4+eJBPegXzJXQmpkjbtewoOZaSO6fmSJ3w0NfOgeb
YQSQtzuBVU3nS6hrBSamg6TOi6mu878UhtkzSFLB8gHuJuW+l2sfuCKFU7nENnEK
MlNc106Orb5xJ3Ce+uinDh7KryHrtieQFkYZoISbIxZC5NE9jyaXlCJ5qC+Zezje
jvxAoVPDunoX1GZUUAIPabkdOXic3KIsOZyJiqaFLfVAWL2pi9NwG7Nq8Ui9Z0ZO
zytxYerNUtXGPo2JIfTLamxBg0FKfaE2CtRsS1Nlajsa++8pTtV7DOkw4JKn0JaW
gvtW93wt2ErowcWlBJMAKb1hNk3OvbGdXl1NG24OYsgJawCc8zLYG+eXsCnbi2+X
vkPbEtCKNCqdruXX/b/7//68qR285bAcWf8vgqudlixPFaAMmv3dqVb999EKC30t
CRg4Q/aaZjoGAkCuLtTXahp5isyqBbrB3/yd4AeU1q7neff/Ro1oasbBxvTtNKLG
2zlyrnXIWB7mGaAdB1uOb2SBiHTi7UND7o84zc4oF+8h1fZ+9i11fnBYifIWbT83
lTbuRdLrkfGj6QlNccOmddIWH+tY1bwt1L+kNP4CNTIjO7exm3MemXdgEtdzoaLe
hUkMSxBhGwlN4u1Fz9NMExVMhgNl/xbKi1CLd1+JqFKUyEWBY3Ezbd8XGJCIcFf6
IQCDP4r5Y5LhKCZVP0KHsCEqDScBwBudk+MEaftnIvFG23GBz5kt4hIyATaSi6wO
jrXe5E0MnG0ib7enWPpjhqS6w4H8FDtLYiLoyeQfXdV7clvD6vPgSK0VhmoUU1Cn
xPY9zvkqSNFS+HzLyIjgQLMMUpdUgYT6EvAIgkwr6dVq4WzuAhXCreJwMKMZIhgN
ohrGB/+IRO5mAgs1smm8C8BhUNZBWEW1BJZsq/V8HaT9rQy/H1rSrkO76ggwM9oV
L+NRxtEbru1OHg8y/AKFKhgfILpNYWdPWeFOBupclZrBcpG1su5DL+aXqbw79Ibi
956Hzfz42dTzK3+iC3lX++9ILdbYR6plOysP9Jjv5vJWyamSOWZwCc0lpRivJAme
OSzPiu6vddcV6gS2b08ePsddMSf3c1VsPAxVymFpxQvOk82cIFIKI111KgDQVphj
yeL5swLDpH1JV32q28OHM1VkLSmBoyKIWaCaJfVujS0s1xuCtS0gdyzfCLJzqSx9
jETD9kh3uU3IWt5O+e3WulW4wC7c+M+gRpKi25VYlaRnF2kUcpWQX/5YkQCo8gN6
IA7FBZWXds42KQ90hQoWUCfPpA4lnkm7deXTJQxFzDlSwwQBv7gjvorbblnYGnQS
5r6c6K3Sb74ugLbKQzQjYwI7FFIeknHaHol3vSJzWr+M7kQRaqS7nwivcgpFnKlc
ALLpd2U9am2VqIX9GpY8uDrzuZzqunfS0rl/xlcTL+oDhSkgQnLWHhPmF0cvWSa+
uqAG17V898ozeL2RvpHzI1uhcpz6n7v44fky1ZmG1vxPEwONGh+VA5TgczEx++GI
buCGa2WpQket95f4ntQMWuCZ9ajYtHWspeKXUoX7j+pwr27yBffxOHAOJPNWel2H
QFItdk2SyWxXv0771ZGJQVol8F16kcHsF99JNtbFX6u5YUpd6NbeUxAeoOEMdB49
HaySkSmwIPfytcdVqjE5Akq7evGbEJBAfuPHTNCX/VziX0EfELrxQJUgCNIb6nxD
jtbXpWCy3AW1zr2QYXCIvz1lLc7/kV5VH3g3vhcVWfL10yO6dO5ZguEr8IdJhO67
scezXtdKn2h49JuvCO2hmSzAn4ChLsasVBMeISKlGkyzXFgrm6uBw7qNd/DM94YV
QcONEy1Mj5+imz9X3pILaz6/4/37ACb5TMNcx8+ntVhrIZm1+sgA4bp9wOyGosgB
s6k6qJC6R2l50/Y0c10fHFQEb1b4m+Pq3n1TpGwcwUnPaDlMkvXEG3p6WrCEVYJK
OqnBXmCRmwR5ryEt2RIZ+9LIkohviJXBplxs9+y1jqcrjgGYczWB3F0CXvpQGuQC
4T+eYPtwGZPdsYymWAT6xJ/DpuPw+5qraT64R4GYmVsEbCUMq5dShqdVL9JDmOQw
+1tfd+it1ME2bxbZ1xFwDPzLFYVZjVRG8id0mMYqvB/MGwmUxy8aHWkglGY5gqcb
x2OJ20gIKlF3PjMMTE2chHORanMfCBfjSmRY6aMbjiNnHPcayW4xsTEgvgobT+1c
2G29r06/BGrdunzbvBgMbBYH4UHc07Fnd2MKWZCuMe84RnwTSskC7kW3qrVVZKw9
ERG7Ih2A6xVCbl/4Z/fcwuMaxnDGS2Nd6fLeLLlaxdwvWnFJOJVK1TDE/0YgV8HW
p7ke3yNSG7T5IAje2lmRP8U6sWLo+tlJqhz5Wmr9VCZatDWEup+U/veguD+yz/cF
A/6dNL3DwmvULHjGxMJYdpe40rHZBXszgc2aN4jChpUu9k3d7k1mSUxoeiJayKEb
Tu6z2FWdav6Sm3+KYDyMB4kPpaPC/TQpf6iw19RxTjK6Y8U36+THTteLzj+vQvuK
g+Ca2nTHVHS7xbh2QpkmXFZx0FIqFCvfcB26ZAqOrUeyC3iOx/rTc5/4abOdt19T
VtfLdLhy2jAEiZclr0ZdOeDT/FbAQYk08JZRsxHCLNnkRj2VSmPaWNqF6V2jKDHT
rfnezqKwuCPtfrG6nMQlRp34RJkUA/q1Et71ZA2Dm+QhMxYuvLFNv4My0N306ibZ
uYiLp8AX7KPqAUsRi8PgjtUpb51cJL5dbj+zBuGkuNWZIBjKyp/WvfyYVQrrc4tL
KhCszTBofNjwOCjG3coD75t4/ypH7/pjOhblquFjU6Pblv2mgdewoi6omqmJ+ovG
NA4ViV9+aSNAyD3E3QOofAh4fP0iThyHy3eHaYbG+Y0vk5kA2LpvBT3hxKJoygsD
W/Rbs8U9khEmD1drToOfYIg9QsuG7E/RDqLDE3o1lYZV2R1Q2IGRAlYA1Qk74Eaa
lW536pZA5Y7OU3h7HXnTo4vMMDud9sAynOrUC87WagqhYGakVxPmuWy83qAl8z+K
C66UVF9tm1/WEbvP0jjllF3uFxfgBU3/4vtsMRFn93zAQfIKaXRjvmCsrK7bzOo3
n+URKwtXvnVTlcb2XevrNPIWh+FNeImI0UTf4eC/xmk8f8wkRWLCdfOFEZMhCLGj
Kno/qmREfGPzn6YTNhoNgV1HUEl5RO8zRrO0OY9/rKQZ4asxdzalbyU2UGX7S6Vh
fZC8UydeXgbpIYXgprbunQCTKzz15VSdmb7Vv2r0Q2I4ECCjKCNuu16iubOWm4up
ivrdu0vM6Nu6TfbAg1tD5VK/PKN9tzpxnD8OT65tNZk0pg2wij8LCjeNtlQZPYBT
9btTH7UtrJaAvk9T89G4MJW4k+sPEscLe7EloSJMDp56sCJxF9+LAJyGBP5HOxo4
GEBowFdEYBVigPXII9Qi11X96hx6P5R6et6lQzAE9AWwWxWYhw7wwowPkBH0eqAR
TrCkNkM8lRF4KDidaH+khFzr6WfE7KQHMYcm4CVXGia8wMUTRQ26DclTp6ffJR6h
y9vGhB1InPhLEo/Cs62mkvDiJdgVhkJ6caQyt16iu7rjHL2axGA1gkIOU4GIkp/F
kloOcedmKblzdXjuXY88B5tiiBKp82bUr2kizUBbTMNaEMTQIMoQfAT4L3e0ye5w
o9GVFuIfD9QlVPjR8WwhcwK9kSrmIB+BsldtXp0uUn86dIczovf6nufkXpxANquu
RAw4jJCOs13WyXeYfGJ9TXoGz0TKZ2VfKGfr9kqSte+1Tx3gCERQPAZqoALJcrFK
IgOqPq2dTmQ2QbtRhMqXPqoeWC5QQwzQTR+Mn1gJp/jjlG4HqrEysYlv8EpJuwoT
CRaM8GI6b6QmjdcNTa1BRybDB80JNpO/GvusBjem7cIjG2qxjEbm83B5JiqjB7pk
7iWreNXI3cEHdO2AsZFFudaOssxMxXXkaJ0fvNuYHTZ5ONE6AmnAj/x5BUgJvwP6
E7ta9P9ixEEQu570mt9TEIHEJ2mktxJbiJnYPFWTDL7IW/5lxWnNfkneGWkqhvrf
3KHyQ63D7K7/HZyj9cM7uI6AUBhqZtUOkDqSWS5w+lHAIKcWIGwUSWLFNHc85gvG
Oj/WTH9uZ6CSHMtRbXkMpzJKZ5G5HZhSWCSBl4AYNziIGgAyIQos9mg+jJv6PvWo
jV8Oh+4sEb+IbTANAK4++GbPSepWDzSN6V3SIj52O7eXOUfi2KOPrxrpBqyYET6d
MceM6r94KbYwkL3sKZB0s6mm16VHMC2GM+4hCFmstvV7w4p1jULQKw8mhqYKDBKQ
GIFONpPBvLQSh3rf9FeoOARAqBz8Kuu8mrYvz0hcmMipk2BX7ARHZ92DTE7BaYoz
ZyN2SNknfJx4jlC8qfDcRi5r//Zrvo4Fh5cgBvZb0rtMVz+A8YPkA+Uf1Fp/fHNr
o2hOp+5yQAtvt5TVqhQgAM2a4OK6w9GJo1VPbV46NhK4Zcn1sz6STodoTIIuTxMF
B2yh8Z1HycdgnhXzApvvYKrVRFW2Cz68ub+7RFEgpYeIY6AzBRlX6OaiIO6xhclL
roC5dltLqTZH3DjPdb1VUZema5wVPHco2B+joGPJPl1SEaLA6yU1yG3WbTt4lPZ5
/IFijm4KOrmODHkwgXpM93wN6j93mOO9U5eZofNSC2bR+iqjIFrwVOyk5DjqQkuw
UTJEd3CN/fGefhfEEgvspUP9WP8rH9C49HdbyoFToha79CbBwObjdvfp6VocYlZ1
uk/nbhU1VTx7ajcomJ0qU1cJm3c/2nVlPjkVYx/XN6m7BCJyE3XfEnL3MGdHeJh9
gRZsB8YE96kexDyrfoJ4OcrIU2wZV2BJOrjRbEoLPLXPiUFWAsPfsx4ojjT0hw8m
8uBZrBf8QWBQnX0TPmiYpADhb0kPqmtv3grMBr6yghTnG0b3j3Frx9+O/CvwlZ9B
Y4LPVIcpYIXIDUMvnu8y0grkfSQkEQ8/cxetmeUh92oZdmJxw3ctkCCfnqYK2bQ4
0lGOE2gnUAeK3+B9WaCNsAv7KLN9o1ArDjVPDap7eKTBkOmR4qNBkL+cuFu6nQwa
T2PfNyz4fuB550bsJwA/q225nzkQgTsascuJJ5zCzvN1K/93u7oaTuu9as5A0NIN
Z4kTV+/+5wB28JZN8XBYQbDyU7zqCOKFVHOlAvY9PiX50AhgY/HZUUm6giPbBmbq
bdoke5x9zvOLTfGxaH/wH+jtIlJtHji9pP0a72EH2uvN/LPKNpYNzW0fz9OmuVor
dJrWFyITpw20+KIzkYg0G++8SGv1wv62egA+eX84DAr0ga3FcM9nPsGS087lyD1o
A3l7T+4H5li2Qn9jFqIPZwHybrg/uLd8c3/qwSAsfA5FzLG/IF65W58fl+SmiGeQ
yKyWj0NCXTKqfWYg84ZaYmhpH7ohEiaJjpiqHRIoGuzKENjS/ZQnj5hb6wWdIMYX
Qva+SjsJg7vFPfPJmi6rAjp6ZTNHyuWG4qwxgF2qBMDxfREhKRwh/d3zud6Y5cP2
SptdbztQHnB8ZtWZY9okPV+ie43jio/Yo5wgMiJXPCMqzVLecL12aC2OWa1OCrdv
puloAdRcPAV4NLg6YhOCdkUlK+lkJxvaRVaucoWjuZ5dGTt0krSF5WkgzZFN9tRE
tP1/9eE1VKTNrVAm1EIQVQkRM8gRyil2pGm2YEATZFrvW+kK53jogGYPcKrQ2ECN
Phbio0xmgAuB1OOr6/3RpEnLiP8depztcAykuJMP1m/oTAkH/sCa53jSUS9aQP3l
9y+k+nalxq5ckTXVPxscbpE8pqnRTp7SBrygJppo4kSD9quzefvgs6lXXD7Yy2a3
CgkpoYDt7XpUrX6Oidp9S74GsQ5qsCwQDJOp7IpFG5tiQNcKR0kOsiZ5iwdQ/ySW
VhMV/TAh8S3G3Aca77Sz+M1bhLU5a0lithScR3DjDuIifD0vaBzIgij1XQAI3+Qr
2ARgBTKlvbIXRu0jc7uIxlV7ZK8yKvoi4eHJVT0HZvYCsWt/nh/KYLWFVpJq995m
tN+YvMNt0xMVN/MzuqInDHNG8fkZKnU+bN2dllSh+APbNDbS8S4QbLQqThmclFOU
5l0DAWFOWXHK3815bTHFUkYue/l5BoetsnjTmmGD1fYcZaJF46wPS0bBNLN2x3No
tHaT37ORYYOY7fqIaAqEcDVJYkHvUrWFGbLQGyMbLk37qI/XuetMs4gHHIuEw2I3
QuRa8OKIENWQ28Hu1q7mzxkANt2h6nQfEVqpW2OUmHiyAAdoEJbKsWvuCiPKZyf8
OJUZBS5BWTJFTjlN+IlZntf1EEvHJyx2El+Ql94Ilr1eR3IfPanb+9HbfXxPcJLl
aJuefoCBed8O/8cr4OvfGKhNoxm15IAYq1FwZ5ap2WVUNLAregDgH058P2kQgv8n
L0mt1aAdwf6zS9pbNaIb3hgpEpqfbfGn7IewTpIt5kQh1ijvE6yLM6NEYBWAq6IR
TvVtUyZHkh49BYwted/c1mnGsfXfudqw9134UYct43hl7UUl9vMSoPdsZ0sS9XLu
dL3E+4W7a0GksSb0ELHWJf/o530m4WPflR3kOWaNrUJ+NwLvKwXGTRX3f5tp1q5/
q8etQRZ6Kr5wj/BrPPr6Xq59Y89Bk6CmMtOxVrwjK6AUb+a5EHnkhM6NzIDgGyh3
iyUqMLMzvhm6f8PaJvVj9ImcWhrE4SDnwNEitVtuBGKXdZK//v/DnL0FuzZTp7eN
BgCoA4jUmdSn4+6H4xvGwIsLHE0Br9869T8ObzOrH6ilkLmODqTKfcPwCq/bXygh
pZKYcqQvLmsg4abC4eIhDck0Zp1qwRzb6IEMoKNXtRlEAM2H3F+rUqYo/lJy71u2
GFWlnWoc0bYCkvTGJVWj+96gkEmvZJblJ5d9dv/Mh+6POtG80N8RRbNe7/roGwuy
kyEXdIZruQ5oOh2JMJw5tUCW0+6GX/X4ydmt1KULVbGXDuRaNPbHy5OCv2ND0ESl
UBL33CNKRgLNg10vsfc3bmJMJzKPUUj4eU2ubpUVaJz4b3hNnXSa6hEEkMHzVWPn
FmNW5tNZNN6lKcDwtDuz0ajP0fqUYQnOOvMO5w5xZv9Ylg/uvji6ZmpOpgKsEtOJ
mb2XFea8t5gL3KxCclikx1Jvhr5UggE2cxvYyTR3ygtj4x6QDzwHQqQJAQe2+X/t
3seM89KwBG0M74Mhb+KJIERzEiC6m5xqN31ov6bc+2YmGtyI8gKuvIGoIlqVxQND
ok77Rd/wRLcdKFOXOj+NiYFFIuR3zj3+Go1xub2t3RGTwX9uLbl8xeQvWG+WHaT4
GhjKW2Ox7sKpSeVAR0t77CbEFoQ7Ut/hhC1gqFV0jV7l1QRWoR3VryWWbb5JLNOt
W3r43CY+oDxQYHUjD9jhRU4FLb7CoM7rLZexv0jpoctFa0W+Wamj1WHQlyAR+Qkf
EVlvJsB3udObkDvt6/zXfZ0rHFumnl75hgLop54UOAph8xYkBGAwXzLCgGmp/gNJ
m3v8dbS0Uu36kzr049mPlObch/gdKg4jD362WdR6S/7FIJmCRs1ZFDi5ikK08RAh
6l44ij+XDtqRDB0Lb31WLSRA958Rm15PzunbRY2gEpFdgU5LPB1fdfOQt6mSZF1u
QyyqYr64l4RKGLZ+5L+vcD4Y71ydqncoR21cFoxbCMKKTqIeyUNm6/WZvwKKqsMu
ml7FWVeUw69fEMbFJvwf3E/ZbPwSZAbPuPeCGSSXX5orwoU4DoHXbLzHuGfZ8Spx
vuRJQbezY+VzMgGY06Me7ljFOu8tsRPG/1qqSK6BWmfBKQo86h6R+6wljeX9fPXB
mRtxES4ZaBQgNKUdziI5jVcGEpNaXjMwV63ILmJqtokKPmfYmrSjeD5qwT+WgPwr
oA7KZCmLT/YiTH8NfZtwG6AZelsZ14IcB8voZ2jXBjmQe8KPRa+QcfVRfvM1B6JZ
mZmXGjKvRAxissDQt5GaLm3sO0yCuqb6RhI4mXJ0x4Lyse/aV5DQYnHJCf+h29cS
ZqWrjCi++HWfjv3aKR9duYxRHrSuHaOnwlYqpFOcQxMJxiFyn2caolNG1xCFN3ob
BmIjPskGh92Ob8GqMO6uGDRI3cz1VpJo0Qv4junETnPFAx6fHfAli0geRJEmt8eS
FVIJR7ZhIjUEFw/AiMZgP73eiuY6btHMxk4V+tQLvbuthf01Nz2pp0dIUL4Adeve
Qsx90EA1wV9nP/qXeooRvCt0M8MYLJ8t2qo6WzVAR3nUxJ7BCsZTvfWYzvEhkqfA
S3uK9v/4WTD1tnqRLpILEod25HVNjOFitno2S8IshT/mO1qU3i1womu9oo53l7yn
SuNRMqsYBT9MToTiIfsowSoGyRUoQ+rY+dLMcTT8puLeXZrXdcwyGVUQ9JjS5aNq
5A83LFymN6Xku4Lggm/HinGWNctK7iq9zsONwhrBZOht4lIVQzNzXhqZSZQTJgdJ
gts1QTpnYRGZ7brZk5F0X2Nrzk3feoKnPu6SpdVfBhl6jHC+snHahaEdN2JmdsTY
qppn41kFs4ls70tXX/yXsjYhuu3KYzbKMgC7y6R5SU4ZK58v3Wz1IYOqH2bxU2Bk
e+KrQwHlCrjEhu9VCRpgZM9CeNhVilTltr39wD5JcsacM65WWpMhwqsqS+8YsCLR
lrp7tjGRM94YhuTFtOj5X4PhLKnuXTPRzIzbZwj/yOzkDc4OCJUvaxgOEnUj7NLY
p1EsHqGloP2TheZgSFtSOXwX7ldcg9wGcYYzlT82KMuReJsQhnZH6aEs/Kk4abvJ
65Nbo1Ht6N8r616Ne7EWBaoPaZvSiDMjuEG7AmVE5SnYrlOeYHGeWgbB2mEtyIj+
4a6z7NFsKDV5mDwMnHK9JrT7ZlvCwgNDFrCcI+t8GloghFIaX31nzWmbubuaSCGX
GPn93aynGMvCCbPOho0i86gIMNtmg4dmwpUKIA97KPdMyZuc/KTsFeXvqJHMIyFf
/DEhF3bBPWA9GPhU8j3s48HLKkWDFsTIWpP3FbT8vpo3FYVlYqORwtRPh+kS2oFb
Hk7ESJqfHBM7E18jOROVYpIv4yGn3aWkPgPaP1TV519MToCKlk8amKpQSDfnXJly
H0nbYFSWub/M/7dkCre4mTZKQklCFRg5XReSi4cbHL5LBpgjQ+3mMIR0lhSIy7IE
5bldxJBLECeQyYtoZ1cS8fNKAunZzXVOZe+owdQuExoXh1NJBAFIr8aFCn5PlCIB
jp3r3lvljGaaoTJgCOqTgAByZZAx+QI89lNyWhIJKdHZy2i8OwvEyG5dI2nThuKI
ZKxyC9Da2H7YmcJtttmbF5BxGn67arFLHhs2LYVMlVS2MBgLK3R8tk/mVEHKUuBP
bwwj3oevYMnNfr5QR8gvfsb2Zc6yKJPJM1bqPXgMsr0iB4vydYMCq1zSUnOunyoW
879Rnq04sskDDSPb/ILPOsM+jeeEgOnP3W+NDcmiDhm+TCSDbnJCOoPzA3GJhlmg
t0xgtBhmkRnviyveXbWGlvF3UdKWCUjuhf5e5lffkMX3I+mSK7vO7F4I5ME9HjjF
cDmXDsME5kCjiTNnmULoH5rAlADJphhCxXxENloGKfTdn80UZ/GAn8n6f7jcIFwG
`protect end_protected
