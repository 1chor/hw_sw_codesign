-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
LUZxUX8cgmoKqx1NrGX2mvC6cHtn7bLIi/2KulynXEGQhUIvNi9k+Y1thl679v9K
KWqvPMeJSQtf+PqT2+QBkzqbUxoeXW/sdh5jOZTejWB72eXNPmWjgK3bmPu4XESC
O/JvxWl7dhzxdA3I3cHWEyeEc3bmkyE0uN9TfhgD8D4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11614)

`protect DATA_BLOCK
GEVfnNk/56Py83RHsS0ZqLZmBO5IQgcaiOY3UliG8b1DeLXVPDKAUVae3x835f0B
W/MZNYTf3yHNRScMo4qJ43j9hh7J5SO0X/to6ZOtPyi+hzF4cL69GK2MrKaRTFGc
cfPpobAh06KfvKXq/CCijgIH625ik1nt+Vzo4Jk6PsUNhK3HNJahcF+yqITESEcB
YxHwv4irLbJ8iSxl/YtUdGGKgnCm73lyXfiuHlMJ4dg58wpg3dhMIYFnhjvGo6og
YuXUoTLYhB/9zb/McfGKbKN+pN1SbSdGC5yQZPsiOmv6eMEmz6iGc8g/OGAjH+wl
zD2lMBGKYLk9jAb87a4FmvdHulsr6yH6ZxSG/MHHmqZ6Rw7VSRAzyNzZJUvo1oc6
0C01Zzuu7sbglLVk9ZpJCDMb2jWS807teLzZ1UKVY7ynCXxX8ePZacYYKtKY/3LV
ss9oZx0RzZERCw/bKrG4BZ4T3xw5ahWo26UlX/Qkiv7z2SNUR/GqWL4bW2UG3PDU
0bM371HN4pzXUEJwOOVyp8iSxJbuTJn/KgukomCPSJMVQnpWC1uDo89wOpE2Ja1+
R4b6bZqUSKGWcxapLX+Zj/3TGaOqTlIh+bL8dC+iVo/eeCdqq76k/42M87SSPrR2
8Nh37HSsF1j7oqYUbj7ogzdpSDAiraxOTHKRZ4lOXrEXEuDPPWnVXCSPyqqDAkfZ
catGjFYKxvCF05HsDpciAHm0dynWRLOWNMKeMfF/YFhpX/FIujWxbFd+aJcWeIoL
GHS3gBCZbSrCZ0iaMsP0TVl5aZZeMzJmLSlIrPvPO5FhoGZsb3Y6ab+Fp2dsYcCL
kUKz/rpSNNQ1KdtCVNC7GByhQrmLaQVhvipH4V//m0ujNNsg92IFPviXaWmymEZE
+MynS7tuAYkmAVpVPH4EzYNBesguCfPwXxQUlCQpTenf93ypq0l9IMghRz7NNVcq
zX/HL9o1+WZjb425QmEUjOKxFKu1uhJASGCdsuc68/NGMHOdFNYi8TAQix6pDc4n
fu7q6JcOE4L3IkGpMwY1i7x9HVs3aO7S0AXbCl6454j/sMBamYcaY95p1jq50gDK
+l8LXejc7uwDC0ciOP5fUFGGc44YO41IoOl7yuJ4V+QhYGILpgeRpG7UxODCISxV
Hdr9O9v4vI6mnEeBtXoQPERnIyqhRacsu5ZgJZ/Uw2J4ULkyCk44zh+6M477HBsz
ffJK9H86juwBy50v3YyCz1DBIK/Krjn4+sKoWK6NmvLR3txM1TtUwuT/EoIZfE6B
EiB3elsF1er67j0Vf/c21ISJTTkG+MRPwiQK7kW5Nw/rjZIqgpQPGitsNCmZNOgr
ifecmZ4cneoUdi/LxxUF93Es7v2pIRWSx9bHGsxXqGqsVR5UfGzgXosJOmp+rO/s
T5d/LqdQKqhBP+BLAtcY6JXP//HfYNdWP1WltoEtjwEIEnPcfDSG3P2vygHIZ0MH
Ejpzwe34CVbl3RGZ2SU+IvHwOxyWqX4YzU910FE15+vgA0VUOQCA4uyiT6fivWQh
tSTEYuRizOd1epVEWAnvZ/cZlL6HvkrAqzkQYja8QsaAPNcB+hEKp/WHMSgCRINH
VNGPX53/4YWWBJnuld9gDxs6dvg5xI9EABiBYEcYdDEpdfbXtVg1nBt3J2NIjC+h
ArChfJrvm0FHLqNHl7PXCcPcDdDC1by6S7NTTtmKJS8Cy+wrokbkOnTHQoT84B4U
TKmc+KyYnMNrysFWlcZQiCBqQTYNCpyMmepEyfGUuike2lmuB9Ou6jaK4Ia6lZ7u
sEB4vR8z8er+mydzTfjioOv6EPV82aY7fYCdy9AJWzpLHlgpPut+zLaKNp0uQacx
xh2X/Z6Oavb6GI5uIP3qAlQBMomCicgTova8SzIdVpUxzqTedgMsup+Fmrz1lwlg
KlWaKANCUh7pQIKcbv89i6ChuFCn6LQi2hZBEPQSOaDg9ztTDwY4pqJqGjOe/adi
q0WYsEBjDA/XEGKJ9PsIjEZLjFQahh5O/xTWJLszc1d7D2hOaHO1ciBjVpRXEQNc
EYjpV6raz/YvyWejnoreFoRMDcSeDj8jNzQTWvvrCJZAiJCXz+6IDm0ay1GHnDLW
6czb0uPo6TypqbM6Lj1sszWmIrpoXxsJrZvHP8ser1kN8udFj81/slQC56WABv/f
O0cHMNI3zKzhq9O60uvQZutUWdt1582RciQonjlCc5Eq9TpSHHATtBM51TXVG1se
0RgAP7MoTmuTDtxw58XRfv6kkRQUqq47gNScLZKRJ71ptoPbfaQOwQq6ccPePOoF
r/w7Mv5NzPruYugLoUHnx88gT/BUUsMZvspCaQ4BJ7h/AE02HK2/XLsoKahA56FD
tNnNNB48ywRnbaJnTxd+Ihk9a2sHsRh9gRIrAwKwedxAeNBulvmc3ZHEQ+MuBuO0
MmDGUakgzbFCR8aX7PAtTEQytkqzJGiKEnwF4hct0/UP3CdKc5lwmXknkgDuDTBM
LaxJsJuSsV8ZvZC0w+hr3CRqDGihngYOMfsklQiOsp1KQwdPxeIgDeL7Ah1a1qBv
6TakM20va6Y5USKTGrQU/jiZ4CxCNEexEVNver8Sm2yQIYKCIvJRYS9+NcpZFFu6
0DbXdKaoQNXFxKpZNij1uyyxOGVawZPy2H9ab6q7b3+GthfqqtPc7eFp5iBb8zrP
xFmM++Yn2hGrNWpsqil37z1UvWr0qorP0ntr4clu/bsgTSsOIO8IWDsZnuU7u0ON
Cjc3w4m0FhFSL97O2GbVK0d5J86EY18N7bPoSxYdbFxe07ulpQFFJFTnr0dS4pzB
Z3AB6jhpBRFExkjgBYFDx8spmIfKDrMMA+nWwzzYHv3Ir+wGib52bqv6PqcrCH0w
EhHz3O8xFNb8SVohdzHtMLoq/e5FJc9XxG4kBCCBesBksNqWLvtX/OrAbRF1FFJ+
eXY3T/LWmaSUMOTWFQwxJaTZQoD8YSLK9UJy4sFZ9Vb3pipgd3C+BOUq5kneOBTp
Q20prTKUqO2KiRmF1IfMYBk1Aw4R0mxH/QKuK7pFVuEeqo1L43OLa0UM6xA/31gh
D+vrRKswq5Zf2FJN+bR41up41dC5U9lzLY2mguxXiV3OeDwR96EWQRxC3ep6GbcO
piL0U/K0mhDnRaRh5+Oljuf4V9lare1vs7ofu4u46h4t1QeN17XTFyzodD+Nvjq8
MvGQUjeE7HcLdXJE9Ol0eaYDkch4jqAms7pv3naXMmmy6uXcUK/NGrl87g4zpm6p
bLSgs/1n9zStjFPGuLzap88ZglxWl5LefhQJJydYhre4o8jSYWIkyfTCFSif1TQD
QRamg/1ahgX1+/UsUo0zzdQi0+d0mMWCsWokerwaI7BWFDm/apzA4pXz7qs9p8Ki
jfBuGFoir/7AUsUctvjsc+r6H8kgfrrJ3FpfR/prfDWUjMGUuh2fAjSfqvNPwg8b
1JC4IKaYqlS2zJBmThIbzqD0ITtALpFpFaALjA1U4wLg2/iXDBFZCPCRL6NiCGvm
pQml94XHXz3/CZ1QHXBgRHISTiYUrDFxtFEElcM/88mp3IfKcyN6Y6wpQo370xBD
ESuFXLLNB+q6/LMWRimeguhzWs4IXgs5K7buyi9XTLEv/Xn2Nf/FTgDrUwVpjW/h
NIMooYIqtkjYIIY7Cy0B+pkJujKR+IqU/G2Jd/cvia2flrYI83WnVt6BRnO5k6dw
dscXCDWNxdKbQIQi3pOmz/iWOX47HQ784VyAb5JAKY4Tg7eGcrQ3j4D/AzBeNkVJ
q+sHIA/zVW3tjp/ZzYYEnaRPrkum5Fu3k2An7gG1jCSql1ReBJMXUbl5G9SjNPFq
Gz4Gpn9UBZEO2Q4PNx6dtWyAUwZbOWzbdoRRRfUSshNORUGyD/vqlZEnZ893RRPd
b7583kleVlrXT+SsAG9xQip0/f7waAyFPDzfueHy0rQR/cmzm2T+VJwCPNIrTzJD
00M4QyvTUwaPbV1t3nKgM7mOiOP7AJ0qoorBWojHDN1m/CdVwm3fmd4wGCTo0o/J
4V9BbOqePGZAorR/RUCViP4t9YX7t/HjCnGo/8rIqZFQNUV4Y21Rxyxl2dIvdNjn
Yttn+pf4GrPOOBmUEakikn4ARy0rs3uOkKnem2JpxAKD+c1P7dGkZuqvPPYCVwza
Y4wXWa94jJ05H0rQ/422UZKXu4DXrECizY/bXKS9CQ8RmJgsDYWY4kLCK4XsopJt
Vd0n+DZxhjI+jXvgAdz1XA8Tn3RW9cJ274fVyt4pbD7Mm458NHa6gn1oKrIxuAkL
8HL97604jd7j12Ty436XXrsDAWQlT3E2GNvO+On37eHilZyACHFipeWuRPenZgGL
HSg/zh1N3ae1DldEUIEO94hvY2rd01OpSKSPnIzcOe3nUKSNDdZUf9pDJPAQKjU3
uygnQ59Hjg/qw0JnlL9d9d4L5VnVum2M5DaL/uSGjTkbd9iP6hDksdVKRprvkG6c
VcKQXbH/XYdgS6kp/LB5hLj6Y4PNTRjxmXDSDNwNS62deIe/wc9L3+AReQBahOOI
Y+RlNgLaJMXkqnXUO04/9QYCRU8qOj2IqfzEfuJ7CdglfgR9zY78ZnT2+qBeVIwR
9mdpM7/+N9TVl8YusX5qgKPAM4XjNMp4vDBP3Kn93h0IK72TN0Jhog7XaDBEDquf
7xiLzJyU39b+KBU8X7kdcDOoP3qqutc4E5H6vPHRJ3JdrLL7pszl6h5jKG/Oydtk
cdb8BPVfloMS6CtN8n+5bP1y04BctHXlrQR8QP04/NMdmZEfNtHH2u44GNFiIfPR
wMEvEfx9f1fCcmDERXKWx6BBjHnrK5cMoU5IJpdVSJQJX+EaTotaa43SuCsjzHkQ
wD3FGzB6RIcclcDFzEP57/TgDuPI3dB/MFuFiL12tJ21L27TtAqSmn0ZKBaWnj6p
xLxrd6oaxYHZRSMJ7N4137WFkJ3N+mUPVeNaaJIqEtNrT6WjLef+GqxJB2JSC9Fg
ncqfOlqkyoglRb2OsXAN75PyP2Mnfd7mSLTSZLlNa8BWxerKVuvgCFoVmA/158FY
saK4pZ5sYxZ/51aAAITtrVwSK8s8aYC+bnkuiNvi+xH8tsXC7kJ2JIwYljaYyehv
L8UyNxBYlLADFCtuy5LnIIYB9UDYxfnL1/7V2iOHQ7I7we18nVfuxORzQQQutzIi
j5EiXlpWNCH/ZzctW+3W0dBc4MVzAZ1nCxAMjhp0TK8b8NW8f923AspmneboeP+z
itKMDrOvcZ/GT/vkqsKGLKcRbM8wx4auKN7IbO1nBzcBC3D4E+ISKE/kFgq/cMtb
TlNWUwN0JaONopohkupACkI0INtHFEUNk4Cuqa6n5Cznv2BUDZmPVAjMNtqgVeXQ
fyVJnxatS5expwQEOAObXHjXJkbV50UtybLeK5m98irc33Y5hKb3Zr3M1QZJQQwS
O8as93T7Hy1VLdiK8XkMtSkvWNlOfB9QToqO3FEncqC4EzAtzLC/L/VDILcg8O67
UIKbNfavPQ2Ibwy4IFRTtK1MS+MC5VaHUI6it8hMZ7Hy7eEuTLkMl393pNBW5UHG
uVX3lG+ORyhhF37cLQMRZpolT0c3/RS/7OqALMfdpYj54EQq22QffehbXA4RxqQq
9iNdr2KjM9wOdx9LmSZ59HLtrkF/02AFrLvXC8w7ArwPOovPR3ZtFhxIW3OlPcLB
dJSorxDmZFvgZ1Rqor1E3BSsTV0HaqH6lxgdCmubdMhZx3P4q2bi0/Z4R6WltZaF
o8TVuX5W9ZJLDGTwyRH6sIpPvquP+JxTPRbzVbeqotuNNfWVeOhodtHd+y+JCvYp
5VkkoxMeatRJM6In1Nsz/u2Ge/YKE8uaAE7PQC4rdpjA44An6VG9BfGAt0Q1f5ck
dyqZZldT3lq6U3TMqdXJk3PhXAm5ZDIStI38nuoDFgMjkc4wpuH4dTV3d96nDij9
izkOcE7gpUHWPUgUjc3OoxzJtifxhsKlMEu2tqMt0Bmc9PmCzRLFuPbfY7y7J5On
kGsW7HT4qr5trXBeKkdU396tOafl6Wr30enYIh3Pojq4JRxCpZJYY71Qvqy43SVG
Tazdo4MS4jHamPSInWfTvk4iZz+55XtpvyXdClFBvD4IXeqQJAMvvTFkQb/FeTTt
/FN1COUNqG6Awq6g5yx3Ny3oHFVPuJoP+NTD9+hCG2nc/TvNdk2KLaEp+xxxv270
wJ/8OUR4GTcVxnkrPz5U6MDMoVs2ZGpjt8eKB7o0wm+Y63WYWICXpwxT6+jm5CAd
njwJN1Xso3a5KJh/iWMuxs2TxRCfPrrh8FjQmBrds/zNXImWUB6uroUG47t/qXck
kxkx0mr6UVuP93DwpJ4w0fx8RBzcYx8A10w80t4Os5ublqj+qjHbpTRr+q5HOQJP
Mv8vVI82KnyPUTnZ1/he++P9rhnVEPevUnyyBLrkV/48opZKLLIN111cSZZZec2G
NpqgQvnvZfdPCzntUg7b+9nZ9oJOn0jaUejPBMmidbcyfRlkWHrXNSLTXJ6W7CbE
veQAxjrC2QpnPmADkDUXSDWfs9fiu6YcWVfuPIDzzVFpGjDd/fmj+RKfq9XM5xtH
YQgaLXQsXHynmBFch7W5AdadEqCU/x2ToKQrJ14MLrZemoumZMDHQwWAX7KlSTYG
E3pc43Qa56soecyfedeD3nwUksrMg70tSS3I/LBgz7DfWHcuEYLjyrtkIUnQDG5n
rl3R6t7FLQZkBI10k/wBBSNNS6kW9CXXFoiflER4RlO3OXFxpv9euxGfwr0solc9
YpbutashN8GY2yZN4gpSzsLZN3zT3We0TorwzzQYCEWMBalfvjrAsdzRnPOIFMUz
VQzF6eYI/oTz4ha59mg5n0S7iV18Cb6mjNAia0sLbJBPvCXO264QrDtvd/uzmgsl
AHzE5ay+4AbPe1Fr5GtGUHtnoVIq8ORnJ83D8XeIt4MYGXFty4zaTpDzfZXvigTq
LbnwVH7dB80wb+YWYHKu7sPyztfx+VIyyVIsEDyTBxJhtYCkrcsZkBGOxunSkf+U
Z5tbNGIt1NZ/6CrksRzkWPVAE+SfnGzyzsnO4avA0EH2XhpKdfmCT51YiOyqk1gj
dnNLDn/qK5dIjk2T2jWtRRXPrOehxDqBsZvTVdVA5Ja6I4vhMFy5STh1xi2DH3vS
uNZmUOiHcr6fHg1p0tFjXr+wtDWzRgW6MfKRt/YDSxyuSSupbyiQcbyOVTocjEFB
PdnYlk9YFbvT8uyx+0CrkpiVPyxtT1/X93eN7hldIM7Ar5eZdIXHfeS26Fgl1WLm
aRgF2TCFozEOO1VQPgPXAkx9OxhY3gfLgBRu1rzjt4+bOTloPJy0c2AxV/OXpIe/
pIzSHDa5Smqa03PWuJjUWbuf7tRtDtsDB2gtTdaSQqtbskvzlOBRKUm43ZHCetGn
g0pMN9BHSI9GdjKr5+c4P/kLj/ps05EpCR3ePhtL0dWqjCxBkXTANLBofPqSWCOl
E3n4nC1G6aVEb3lm1eEvytr5iW62/aMNE4AMfMe+av7iACqh+/RScryxyejbKDZX
bDpsNgbzcJCEsvObdK+7/ZHl8sGGS96QAydttKXkMztyqkxaZXGASlZaaQ/U2eB/
thvDbtzVLLsg/SdLfklpe0CbNO7Kvv82gMOwhsSNmKsfHEzoUwzrMIBaqRZte/Ii
HkSGtuKdywsZPXj6W/q/Xf0DzuUG4+qEpiXhXjfM6ogjjiNUFR8n9fXMYl23oKgF
WihfCHyBOT5b6mF78iqfsNt2tfYBl3WLgWbWR+70sl0c9bsq45s/Lr9RDMOcaZEN
I7l9nkm2zODpCGhTYOmB+AOXaSb3KSZbYtLsR47OIzSOMBBzKOZHF4BIIpQij8k1
zT1Pxq+xkT+J8+zVKqSBc3MmyiFdQ20Rs1jkRC0XNVstO1MHpftjZWDLjy4hpAcw
9BL2neUUiO1Cv7P7oldbIkXFQ7KC3+lQkcphQthIRH3FsSGa9cW0Ek5Xjk/ZZy68
YBN4z+MFUo6xSInPdNaJF6CQbn8dk+ZwTPHsg+RCz20GiekUDxp/Fv9TCxnf/+UC
BMg/ftOe7anHYRYPKfZS/oaya3aVfJUnLlER6KLy3lMFZHGv6VTgDALjLFQ8umdN
9JtlqsJ4+7ZwwPLEXpyy7gcZOOSGv7yzTnFGXCs8oOQsclcbcv6xqsNkb/sTftf8
pxna+BB1YcIqBBpiqvxi+orS8j85s7Frn2ZqhyM+RLdWCoD5MJLlARhKFenG5Fxz
5gEn6XChV4Ufw+nmqzwIxuTpMoPmhNDicQIlZ4qLVwUNXbXlQevofHE6/s5gFi2a
qDFjQZ7wdgWZTTZoKr3F3eXrK1NVwKmCIHi5jCs/HAr5wakrTVByAaVimAq7agXJ
GdbLy5zSToz1mmy2vpIW6sosig03Wza2KAeio6f44fA2kAvu19hv/dw8MAd6wywR
YTzmEIFwRIca9U+BaZgBvqCXg65E6yuMGv1YgoI4wSRVhN8AsTXl95Ya3LZ/B5ga
8od5oE6JKVX/g6uqiaHcsdbZdD/VCXWFWPXL+NXnPX6GjIP8H+YVOt2VyIjCys3S
mzj42Zcttc4sjyvE0lBS0DvE8v/g77Da1GA/1qnCYXK27uiW0iphcIY77aHOcaH3
TBfS+EFK7KJXPJD6eu4efr+Qb29l+kzEdbPIOjMOJ710vIsRU1nUSvrOYZsexNnn
Pf7NHxjxHe3Vllz138AJ+yyuAMRj2ds9Vr6P1nXfl2QjO3Ch2mvymuoM6NmPYJwG
5sBEUAnlpTRRJAahhpt4WikCsRmPZp4uz9+A0cQxEtnun4GKh9iDNhNayqEFS3wE
W8UfUp19fkOLet+jzubCWqDmJ8XBxpxU39harsqJsRh6r+DufpnofA0dYM3YvxAd
IXMnTXiFiSvrV+l9qRdndEl8ty7z9754gImB0TcY9Eb6bLCXNDhHo9NdCYrnFOvC
HLZyeisFfJRgn7uIX9p7yrU7xldZxIA+waUcwJ09eI9N7cVludC70QjYod06kBQb
pM3G2khLeBkHXczJA29uiBWdl5o3wmxFp4HDwM4PAIYPBLd7RecS1HMlg2SW0RpY
hQA3/pj+rXqWr6eh0DZ5bdmsNmKUOqxrt0KjfhoU/m8OUtzPja+RnTl6KzPXK7sM
KMuwlXPA/rdUUgh2fyT/52Jhzz5sNsU/GjBdhtlsJmFUhPX4jvXJKK66sFuqLDFT
Aj8hpLkmPGlbEjP/msZsilnvceQw+TaIKZrqpJlVicIT+quTGaf9LqcmYzWHYrp/
KdGiCX6gDN2VIQITtrSsE3FsT0i6+xvUN8nY2riYnVPh9pDTTJTNZLavH5ArSUuZ
+fXbFJsSKccs0mpXVdh9VRrNEWbdwP5bMwrchU4W6LFULR8Agey70ohFbtKGktQE
4IvwIgDj3kFNJoCa5Zj452qVbdbXzc7AlAONvsJDJQYHEXlwi5dj80hTHMxeRCca
8A3pG3HPXXhSR6WZPkDmRmNqivaZM1MamxHs4IQ4rfXm8HZ1qRn+oMvgqOqHwScL
NShe/OG9F1wSGT8QdKbNLNtwMopuU4pxPvW+YQewWUC/osQ+h3iOGjmGJ42ZtBHD
dL34cAf4bZZ6E84j0e/Yp7kOYwLRj0CbFxyKcdWmNEf/zTcYwg5W16qHLToYs6xu
/5IxOhOZpEJl0RM/4rIxhE78LdjjAZh5kD+eaQC9WegT5Z0kVLZt4+wFW2Cdza9X
LWrWbNYFxfGyT+co4xS4WjI4pbrWf75OKzlwx1ssswqplpRZw1G0Ac1bVBbVvchx
f7f59msDwgPHZTojo+mbBsxjfJmgxv1u4hwwJyFX8ceIswG6EnHjF+J/TpwfQxrV
fbPfV+WTaRnKmpSwZdU9CBbVuzJaZ1JJBnCnV7+a4hkSE4x08NNQ+QVb8yN0T3gm
uW17zKWeD2qxSHl7cH9Pqye0lu15FXMjny4NrXEWpoCQMt0+jNNR9MjebhY4MH/+
SU/m0vEtyqX8exGXLVz1IlFMZHGB2kMobdk6Ept34u1Em7IGSl5bip5NCyprEQxz
qcAgdJrjlbso0pcvMwXpKOGpO4hhyof9tWictXcTQ0+CH1mYo1DBoIol+yeDsvLM
PoAV1jsb+Zl51OjsA9avN6bQXaCyihBabv8CdqeP0/rTtHEzNCL3qGpTkA1hRJta
roMV0DJ6QZC9n8tQxERn8lFnOHvCM4gr8AYQRf9EVnXOXbf5LbTBxjtp+gZhqnpw
tukevC2bJ99EzeaPa2Oen5FxCZrYVu0SdoUTS23uzt1edyNDyTgDOQi/oGKS2Lro
hAzkmzs1abzxoPpWjXuui1BjXb3Ah/RGVivTdnM9RaP9+5QPxlUV1oTHcF7q+DEF
SS464wQkUqCAAlBSA+nV+au/03yLF034SdY96TXypJMaF9gLyMVp9EOUU9MNnnVz
456tB6cQYHdwqCwWhV+w1gBVDm7hyo552RghKlMM5PygYt0ip5i8lbpe5g6FYogG
A2wUcEHKCaQ3qLOtmKPNyeH46jDwZdUmfYKpmbqbqSKUefL6+zIlVf1mbXb8w2ps
baD0U60t5B6oDROgk8qV5OK5gXNGBctmZ/9FmAwTdL/o6O+tyl3Mlls1ysbU7XtD
R5LNM/2M7wJbzOWL8WzQByzuXH7Kcfhs/KklQ19P3e+ob3kmfLvq+gg7DyE+TGBW
KUrY2LiNGPkiJ7PIpu6rO9zq2le6C5CrlBEbyvs20gqDQtn3XWME9oEcQR8oRsGY
VumTurwIxOnvbmbVeK4i5YeqwFNXI6F5p5xj088POysAILz9WrNKKSwQUJshjHXH
yAWphXsVraOZGW2HrRhjCVW8xpowXtTVofWino6hopwV+L4tqNNqa4/tgLPEps4j
bBjXC85xSz24PW8AHrX0WCP0A+4gr+0PE36lWAHMinsyGj0DTotGa9lFkzelBs2z
a9sgoRjKGnrXJH8EtNsZ90QySE62ZamrQLMEJodlVDJ66p1sqZqddxdbDcCX16TC
+5jis0jUElB68/Z3ddoGml+MExB+RrSDMPjkNRlPd34ZBNlABHg0icmPZSw3MuQ7
OaW3DiU6MB55raqVxj9sOJSQ00OTWl1o3e+6EwdU1WFCq1hkctLApW1kwFprcFs6
jipBLuphfyBSa6YK8auw8klMltnur/YmJm4z9JbrCLeS53mUgHzlqX4qZYW7I1By
OjBMPRmoUhkD/B2m2svDtKzV2pC/j2EXBq1Yz858+XdVwOkfO8Jb18hxeX834nYJ
J99HcqWLs866GM5AVDUZWEkcguuB9hIy2I+ykDB4cQWUmG26/QQ4hYapgDbhazDL
2aTWsbhz5oz2Q6PBtO4jJogj+lxfERY/1vyt6Pp731vGy8ZO2yctxTutfj7EH0ks
NtEOeeJaRsUaKkVFpCLSGyfJdohhKujb1h2PS1WQRgYn8LcfrIWFP0k5myUJmQDm
PFtmRnUv7NdlmdzsZNJxvXnrW6IHLpu7SRhiySmcNkJCSDivDLqSNd8YOxy3veZV
0HJdkr1AAmTVggk3eL5zK75dritm98XxYbyW3pEuVYgscb4N1irqwP0YD9oSTYLj
AeSG0m3wJcHoMgJknebC5g/bYjdSZ3Z49z/i7BKNNqJ/i8xPSW+In0GniU4+NWbp
QRNi06Zh5HkTGbK8yJPVQrCOx2t0LEm/cCGSqj6Ae9TtKbrFzGfWumx97t8K0mFt
7Sbu4/ofI/JqHPf46dnr4n0ZHA+wt4X+aRCdp3XseT/qkhliIZQ1ogHKh3aq45/x
RW9eLv9kdNOhfKj7NbcSWS7BFmy7zS96CmUWptth4iO3ALLBiJPAceQe1F4R884y
Mekpzfw8XhH9912YlLalbNfmFr8yLePOmpJDHm6igUi0mjU9mH1zW/wmw/oGN2y1
R24fQumXEJhIwbueLwJhz7Uvi9Ka2YRyCwBFoIoumEAG8iCVEI6EQBWFyxWuVWZt
emUMlmAfyVmxeV8wZSG6DLABKfK+Oh4xVjAmbUlh8R+pGBjmrncAj9LinajTacrQ
rPYL2p5tLMQaCbxSH88SR1y+SXBJSbgrBo+AdP+Lx3tlINTocbmS/ERP/E6z4jTq
6pl1eGGbJJSz8/llC0caYgS2LWI+R6ketUJaG6Tsrr8r9SyjxSEH149v++BkSmzW
4dabXN5S6K7WU4+meXDhm4/lSvXndUj2eUZ60/8Vn7yujKr1JmMHumnQaeO6vQWK
POSZQTpcl5jzsXfwWLg7HMjQRsSe96bOUk84oR7pUBIO2ZNqL0eZHI8NWeGYo+R4
6BjO2+DMlJ8KTASl24lhf187tPmDgonLaHY/2G0w0I4GRaJjnxEgYCSxbH7BUua0
VKXwu0VR7C1AA+h9Y6ZBjg9+e+fd+gGOBZ9zSbAHyxJ/nPcVeD69uj7Gj7smZmAU
7IQTEoLQU4HyjGx0Oj1dFzDph3ZI+Uwa9u76JwmLQuPK+TrIv8p5JkUEGxzlb5bZ
h0cOPIGIc4uxBOZhKZTdnMJV8r7rplG+bXW8OIn3oSJV97PygoDuoEue2IHKINr/
mrtEBGv+DPNzxHAfgTs/XGAhVvwNZlZqSDadMyDadBxJTKYTy/PHLeHsobyj3p9/
uUPYiR55oX6NuFiri3UKYsfBHjZO/NxKyLOw0uBPvIH6+0l2wbEmFv6tB9r5Skgc
yam+B1E+TXkruKxG2xTsOeRrXSioUvzaUooYU8/oo1CmmIWYo1bSWaInUZKvVFAd
rg5nFvBbAcPP7ZaZUUhWCY7eYVp8JMj2m8sTn5yJ25B/8lWI+mlFixfIVXhCc4qu
0g5kgj1Bfk+u9JNgCP6cA480XKdTICMD7dYtiD0AEexJN1Aslv0dE93GShB5+4Ic
GgOf8vzahAimuaf2q4amJNLTetS8+JxiLZv8PdAfTKbxhkVqPA3qvHwjUncUBEP0
1bBv+9GPyu7gSF0lt4n60pQiEs0qfwzfVWpH6qJEce6+Hwo7o6opV5jEMr9p48Gw
eup47cd750LWFl/aQEtk3X1HKJ47MFFyNKSl1vvf54MAaZJsahFzJ2R4v9RTtNRt
S/J8scYJ3dySBMvAv+ECUZ1hAAYR5Cgk5AuuhFHpvxSgxE2keiIW3H3yqD6MAarv
HW7nUchTXyxryEL+WvMoin6243HdNLa5Jr66pNjEUSRul3C9VoKGO364AXnM+fhT
mZPxlsHMOejSTdaGsUmSmcsqq2mUbyyHRlfBTg/JrB3AXElKTs4cmBOzF7NEf4xw
23IPhADXMUNXVbwUmfgUqYVi3rSzdB8BWe/yDEPSMqwVaoK/nKXgQDlm+ppQ9ZJs
+WZp08fbuxkpTTvCfNjVM5nt1CgcD0JQqhpfu3J15A3InFsnwfRBXjr1jW0xrZOr
PUj/lV4DDBRnIDHChC22C0VFTEeFAI19kRSOyZm/sMmtyJVwsu/VsQmtWaDW8DG3
nSdiOV+i1kUVC9gHtuAxKv8OWdpPA1ME2kZeWhf08Hxm/u1Yikq8XGOX1tGMcEJ5
P318XsgKjyrkscXnu/RXJ1KxW0jOVMiPzinKIJSp2xv7C0XyDZjkyaFY88hWl3YF
kbfG0PyGL32/Q8pCih4VhMkgv1XtYc2PY8jcb/zAVj7BRkkaMWTSzMoU/d4LQzqr
arCDPejLl0ozWsGFs38cjvqDBpyL23iad1zIBRW9JwjJ2XLao0o4O9MsaCY2eOc8
2jZPAP1jOz36r/dOWPP3zESx+QMJ7V1+Pfm6I0B9pEMuzPl7mRv87+f5lINl2FJ/
cHngTn6UeDkmR2wr6/yGyHCFvBEOyPY7CUE7WF4y6BGP5J5XaR4er0acxH5600k4
BsoXii367e6RgXrthoqW/JItbc9l/ldwsiqOil/eGOTYD7EmXPFTibz4iE/6NKol
LJX3ZIR68hU3tSsq8noYmGoOjXRc7LI3z6rLiUNh7HalnyDKsAlI7QqPrUUMvHnl
TwJwaIeZZQt4SkHuoOzvhW+h4xTpkduTBL/lRjBrwjFGDbqESACf7dGaARpl7Fzx
avfafCZwyCpxdX+WDjnXHTNArKqMW4bFN8w7bhS8YBAwbl9V7bOYDnWsNbgiE8h7
E7het7GGp7Lcp9IC1XJz+aCIP9DGqoCoFCy/VUrBWec5LPOw/r61p6rlrtVmXfX4
Q/s42zSyw7ksNnerr8KEpTBJO2ZVKKCjBgY8e0UOlKzv8zfvnYxGmQMgPR+9H6jb
Mfu94xyL04zHdaNeOGZW0jcjxk/iT+XipHPb7c85baQaAUQ8X9VrMyvr4cuvCB2z
vOC3F43cD9crGPEix/oQbp42vuodOut8mBJs+BPAhhd7XYPEv8jub7/w7xCPj68s
EZqhUU66Ebvo0d35/rMVn57fArl52Tzz/esGbY5e1tgtEugkUHeTlj0ik4MItFQw
ZJswf7xfQPHatW4lwwbXNbaNP783ZG7YboPXZpvuyw5VPGq4LG9r2UXD+PatdgK3
/7oMHOdqY3Ba4VgXRtKfXZKzScHOrAygF6S0fVKkLmX8oEJMdk2+ydRb4ZIaR0RW
l4no9azQph6rgwZK3+NbS9gpujNFvq0Bn7ekDdxnVL6fSS+6whU3jEyfvKinAdN0
CorXcCTsrAEKqE/K+HgMel6lhNPQRamIn0uGvAeaaKi1vHSeYPlVmsNcUckBJoRf
7T3934alNEYJ7n9kb1usr6TWAtvuuqrbhiufA4wZtTzeSh3+58xj9MmsSput8gPV
xZgQRUgp0yAhTtzPBh2cVeCGxm7NzILpm8A681DrS8rQ4p6i3QlgPZIsW65mMb+D
0/nRcC6zeROA5myZvs/csGuQxa/u2jfM4w4P317JLfjIMu5K8gdvcpEVjyPEYL1o
eZQtvfh+7wjd4BjhTzCsEDfjJ7mrc9y8n9Lq9YX1E26J+GwM0IcBZ09NRg6cqKVc
trSLPh3YO9Yq2NKUBdMl+vi2jZQYwbdrwVv65OcsSiLZ7lD5daEH7L/mo6VarGN1
5tY1gMQtZnLUFotD9thIh/xM+ECBLV+/fj0arA+kLzb/6E9sz4HAfqfnXMGoMa3X
2xCtrMGNwgmRAFbxYSelrbsdNp+LuqfXIUsBQQeykuyBqVKwvML7B8NF0uDh1chP
5f23kz6kOLTQLUDAQInoWflFiI+W/EoyZPLc/3r+5jCpqj0WjKH/NcjGZtih7S3f
RoYct8WOah1gYHupF0u4plIHTRQvAzLixkuoWv6/60VN/rAjsvAwh36McDChBStT
JAPSkryki2rpkEdIK8VNaXn6LJngNnpRPsWYwDl9l7janCSSJDoO4ZVvTcHbo1W5
633ngVX3nvdw8nHZSyc8LXe3R3e0C0pjPbutKLYn7jQKAQ4Jpl9JkzPJ/FsaVxak
L6FxWvR7cqRlJapAAoMW0YdKFNyo5wVvO1qEWNjwTBPzuHsqD3yRBf3AZL6sZIur
QACsSp0egDypxiXzXblNwpjd26xIdCzeLQPyGufP3kBWEoNz5udpJ1h3woug5va7
u49rnvtDgurazMMv5mjxOA==
`protect END_PROTECTED