-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
TYgk07HCKefwTCWjzewLkhKfW4FaBYiIrp290IZxkHN76zHleCWR9VpTZi6sEHN+
Ytdl7fGxvgXZKKWUezZfd7bVaDfH4mCCZrRfd8P2hqCosLPhCAVX+1P89q1ZerYZ
xJSRM9vA9+zIYXXgBpDTL2Gp1DkMT9k/Bsukkjr0UBQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9777)

`protect DATA_BLOCK
M1Y22FTilZ8KzS0JmFo192tCK8rnP6FCjK/uqvZFFFG0MZcWAE7LoERueEgElOuJ
QiFe6ROTijzWsbGKKNmv9skbmLak3X512M5QRPI59rFCSG1ZlQmUjYJiJpc7N1Tw
KBkMefRpERkBMdNz5KFJv281zoa5XtzSk98Kkasdd21aN2R2KE6+bkLBjXUNeT4c
NedfNqLaeUNuNbVMgHbKaCSlelXQNrJouHpAN1EyhveBaXnoGYQVrKs3qsWvCHCy
Wzu7humgA/5CwsEBAncPbt5U0Vp/bF0N/g5jfH53/GITO+gT3rTwMeoYqVxlrBCd
C44ZISLRMdJodICL5PjXAsxwf9k92RUUEzaRHs5a9ByGJDtQ1OWMDtrjNKT6Fp4Q
nmAeC8BwfxXf9f31ntjbsh9ste2lFllM8kKUkgWWAWsW56s0N/hHQKb19zi+xuFT
wwtim1bd7fgRN9zzEPFx+S+gj2cwgIt6NQfgOh24t1RC4xyv2kN/6qMgyZJexGbA
xWS/gDNN5zkrtDq63dd52uyVn56K+Cd3oYdryGQ1ABU2EBw9OodRtBp2miBXfYH+
WmKu3mcNvQKyt+53cm+FOrswrQFT+xaHKmTbh4HFyys0QtrD+MbWOHAnfDjW8bnE
9RJ1fItyEh5Fjdqhh5wsgsLDd0OG6CprVl95rZDfm8PCeITbtFWhZHystuWKJN2E
HR/3ED7Mg6ykVJZZMnTH2fCKYfThAdyQ+OyTlwEW16Cj987NYQP5lIMkhhV9lp31
GGU7e3dGboHNsZAYIZHh3CNzBtQgnZ2HSTuI4vLyRFlHtU/GcXRiFJtalq6D4ZmX
osdFAS8Z2GRkUg0bdjmXK/q/aNhCjzG3hmOZG3SMW23ENU9gIQrxw0mfWoFMtF0W
bSNY60/7qtNaQU73LilpyW0XHc+uMYQEHDxMTGHfGsd5n2HoZCZG2lpYaFLRN4i7
aTn7uTJrQ7ydv8H7o7DRh8Vh5tfuG8nl/rdS3/qdqkIKmS52lZOpOX1ah/D3swZK
+nV3TqvYWCiC22rYH+lQJyyIWiPNoWQORpTHdqawj90M3GwDqX7x13jgpEOVeOeM
0cmLmnb1FRaY2bkUp/wtD14cOzF+6321imEj7FnT54Yj+R9oX9+l8jivrWqxdG61
mtQFZcg0TGVoPavEzRuvVwOQTNL6fwPWN9Ww2zrBccywDIoYRza2CLIgsFUJ5yvv
XURLTxIboPHHFkEXoXHreJGMeFF5H0nXLwWefC3sU4JpOUb7V/DKIgKgavklOs1X
ZvNosZmwnfchfIEtL3oj8it/mF/H8WLktmsx64G14XUhMzhvRc6PiGfxcYawuRWb
+4gxLeq8/4hlNgdGwOFqhgNzIwN9H7RDzjST9poQRzJTkZb1Mwj30vCPvtTnidVw
lnFxxBqUmtlvGLpDA/DrFQtkRXZCW7IF1w+8rDooh3C6yX6Ia9SU20KolsPkDPYQ
bXSWUMzyLIyJVTEvF8LlKS2y36NmSAQrzlgz30M4VHRKFLhjargvo/vAHZ7KR/bk
DmWpVrHAB2QpvqctgTjDVu7HLjkz3vhsxUTJtm+vlhZKvo1wgOhbWm1d8efLru6D
oRictmsSVWlwZUWxERh44lqVnHfspFcHaye7LIMRkyxOz+DjIWycgwJsqXG0SNWP
SF+90W0EwgEL+bQNi68rDtXP40tqAPX6TRl930d0FHgTFDm0OAIPLzb81/Q5Gx1m
WniUjsQks2UAN/5i0MlirV3y33SwPCRcmg41SNPIfDmWrNZ1A4lLUk2/Bfz4PJAc
UN1l9Ww/8VqshRyyUIi9Trrt+mE7EwBzb79Kh4OS7YufeYkJpmwwVs9h7Ou64ETd
lUQXfqgnELms4wMCd/cEsXUOnSCnS1XdxuUzGPHeyTkU1okx55J1vLBlhEW50HC2
ftZOmb1XfmspwXEohKjNMYP6YvBYYKJouqpo67WwcNk+VjkqHJkFM7+6V167k2xw
RGTldcFkwJAek4qpAxoLN5+rkr0MImkDNFbYLVQ2oVLe6xu2jziXsbUewRr8g5n8
wGL0aNLZ0WppI1adhl1VehMy3lWK8owzBkj5Zn+rCX89ksHHh2WbvSjWNyTvsK3Y
SckyfxlvHeuO4bbDbYXQhfzVBN8fG/3wvaJD/NonAQCNDXbZpagM/5db0DaKbRsc
vAZKVhd3bgLWCpaP9yTfyBRa/hWuEY0tNeB0UY/TOsXfAc6z61ExFxGNQXzP2g6u
2Y5mk3iCevYt4vi5tJrhBgkZvnLt+tXTjnDKmRdNE6tWxjGGtfhPtRleA3PiITCe
qXfN77vTKF8IKMpc/b29bdhsIlsfwzxdx+DPMIbTSeK8gFs9L39ZJQiYj8tEPZLK
w0V2QNJ/shL9xYl1TyQFbFrXcqPEhHFrS8onEbnqI7Y8yqTtzSjnRC97trrAd4AO
o72B+d/KwK8jk1XTQ6rKJc2B1QJ5X+jlHYKkPRtIQrOcV274czNmcoCoqA3O5U/g
d8xfvzqqhOeeRo7TqVZ3BvBio6sJT3elWvJcBywpTpJaGvutR9y8TEDZ0YbXu9a+
3MKa9rQ07c661DFlWIfQi/gCwmMOXg6tl0/o4XTy8yZPFc/iRMBJNxXTnO5eK2zl
oEucpIfkYoFKcZ2kHwX2tm5QdrNQE+oV7Q9AWtB4kqv9gl14y7dN+s8AteMJiXoa
QbiR4cILcVYbu+yGGQVNXmwhWukOrDU4Wlh7JAZgCDmu5x7gnGmfnFWmAaPGI3hT
e/hJbuIuSBI2T4ukg5RtAiMQoe3e4OnX3xzcBkGHP9AQgDmuB992QiZs7gF9Yiir
b0Z3A1O07w3qNkwIm09urUG2w8iO1MYL4N64WO4o9CFh/8ZyadDnavx2yxvWrDV8
ZZzzmDZ29ArfICujcl81QQG1pdQlk6/AFi2wDNLXiT7lS2OXFFTgzDF0VCwThBXV
8PI7/v0YDfeCZfZeLY+j8j7qE+ZEMW+F9izgSujxB1GUkvTR5n0vY1YfAE+z6Lp6
QuDhmbnlpe1ueLBpKDt11EZ8ClIHEREV9Uo8wAbg9GOfodvVtfjEX2E35zCJ3gi/
wYFOzqC8+JHFz/Shu6vbptagC2bAxjHPkrARtVeChYEGBjQQAegGMNbSk5VMqfY6
CwMwBO0NnnOueNVvJuKzxFKqytCoTnmKYmVRszVyeHtNv0FxS2TyjaDu/wdhB4aj
IcZtWwLesEM5j4NLVDpOOsSRa22jod72G+7z4lBv+obEnkY2EwJlCZi7MGrckB+c
5O0WyL8naXA0zhbBBA7XSoL+sbo+SJaoZ0eHLaBG5i0HdKaraAkPTVmtWHqoI7+i
uaHo9d7UaplAjfHFu9hTRo7wBJfQwa03oi+o909SElwiQUwUAcRSDFoOMYvCR5gA
bIrf05of9FOZ9HNbz9aW95ze7lfJqLtCx7BoTTL3QsNHaYnPPjghYXOYXtAfKSDv
U6g61Uj74kZljw9DXJDeorNI/JtNymFD7X/q7C5FrJOr426s3KX0CsQ/azHpxrKq
AhwWO8yIoQa9dU9D7RK6RiacphAsE8qYVJN5aXSynEdU9Oy6cZqt6CaclfUFdwqn
LwV87nmgdUXWswicS2sC8wqHE0m9ELqxwrPWd+Q9nFazshHg6+x2A8tQ20C9x9Vj
kFMFEwb1pFCkTgv6dnd4vVlqhMUfvpZUPLTaHVQSMeuewTDShKfmX5PFt56pfwWR
fA8wYYk3bbZPr3kcnpJEarFjk3eoDcy0JKJB06ETxkl4ljhf+gBflhd0wDkNPaO3
2ZGijuH2CDls1erPpjnnZ1Oob9Xw2chSNLhFeD+9uuRc+7ISc39NxJTDtfpI/duD
oKuGDic/pI1+5p1SwWniQpiWVI9P7Y5CFNikG8MIPGzPMtWXU4YCWEYHL4O1Jda3
xPquGgXTQ475E4dPGffCd3DXVPak79TppsVGSFHLAhAhYt1I7y1nrWm1nxcF216G
eeYYNcRMVQXQSzCJuSjDe9b8/glDR/nbo+wkVqRoHOn7cGQlCNOQK5NBf6g7+YF6
VJ4/6vbWnBd5g4RlLmQh/3pliWEUrI3Sxj2m6YUWWlrr4QZLpgD/rnX0Q2gchjEd
7eb/4U+oAesARYNJKNxPfz1ocIMoSqhilVdbzkaKRdScVJpWUesE7MP7Ergr7vrl
k6IcClbbBUJndC+joICCAil620v/xJ3Zel3ms1Tt40KbJC22EM8uvOnEhXTXjhoz
NO4DjCc9qQJ0PVj8GTvVmY3sFozIOMdQuENPZK9fvUuTHwMYlzkzYb8g7L8kXq5w
9sw/d2f2rzvgZSbLKOLVmpYUkKnXUD/wscs6z8KzxgsRZr1JmfGhnCaxtjwtj7o4
gU4vf84c2y3E0PQfVG+GmXjXRGo7zcgemZKlR2A7efmJ2MgPX+2VUyS2dHEoNgRV
l7dbLf5TQVsASaXnFN1eAm2IoUywUwG/jumETF2CEA9/jpfG8oMpDVV1CgkcVMC1
0Kpupe8U97ZfS7G/2gHMSAw7T633bCbY8Zs7vjuMB9diRgiKrHkz3U4IgoZJJ1M5
IVJpV3KfxRyMCe9WUEqmPbD4x3xfD/24/NzEBsXH2k8XN/pde+GqHdq4ECYZMjrr
EIoFojiNRiwIbMPiNkLiyBL3uYpz5jJ6ZAO5odlq5ifsifuWm+2O24Zxlut9e8Gv
dZG2f947VmYDpweyJ3T8LrmIY9YtmU2tj/NsHBLrT5v6R8KAmeR7Te9OoSUr1hTq
pSVVSHd+KbuonFWlD5fQXVof0SfeloU0IzO4jD03+y9gGYOI28Ve9VEz0o0icP1D
QOzXcTSUpycXBEDgr5v+fv0PJqz2R1Vk+LsZAzuJ/alkQewg7oUSxG9fuejTVhPV
68pIMEy9csIzaHBD3hsuQ/lTRgydaM/sTXGgujAWUpE05vSbhJ3HXasR877z2VpC
S2ud3ilKC042S98IDTU8HVIMUolkDiUOvNrj21FVP6+FzwyaiaeTCZ+M6sjirWe9
rlo5XHDy4jgXcR1OXJALUr5350eZv6oLKuge1nMhtCj6cbXmglr0fLciZDSBBw3U
6YdGW0rs4CUEpCrjY//FjZlaaAPSQuuknjj26CsEueYKjfmEqxTe4Q67M6a3nec6
90WQ4X4o5ItGxbTm2bftinJ3WC4Pisg81ErTdvzfUsNaJo7yDe59gDJ4Ef1kp6+l
32COMFFpeczRp3BZ6rRE6xgSdD+yCFneTvK0X+t+gOM736IDsjB3/3fWpJHWeO5C
sesKnRDgS5I69R/fe3ZLAxZv3qoeTYxK4isAGaxz9h8+geWtZ4LTvlAliSTbvozL
cNTuo09bIzhud2Z61mnNu8ikQKtr2j1k5mvjqpNz27VD23AXdTtlydwpnkiDoNAx
+ZfiTX8Fa8k3kmBboS3K0k9/ivVAuu8thEiM8ybtPt1FvrRDTvyfBh0WNtgSB5ha
ins6nr1zTmGVS9VjhWpSNWpEKUdqgsOSlvJ9owU6BzrybHdWj8yuNWoc9T5LjOBN
R+WHWL2vUAg38CYABi6qn2/x3qAzQDjzE5jWU6U46yUnXHAlh8jRLwaNl34CQlAH
krD4CB3RxDu/7Vua+uQ9GdUsURR0NgYbhUWbCd58rxD5iHkiuLQG7Kv8uMkMansN
GOhds2hjtRPY6jVs0uHMMVwDeJqRGB6ixkOXo4rF7P9lC4XKXNHBo3A7hlKp6hat
wNlnv+a91M1ntP3yvRM8bpshV5eaC+O9yVPFsU6n5908fppSpchc8ZhAN7+iStY1
PCGnIgaIG+qlpWa94qMSO381RrOCi2YWYN0yaeoLguEjwjMKOMjMUu8ZLR9vy/ko
CWVwrYkNZQvv3JVAaCUN64alJ1MQT0OYx3ppZv0BdfwDA1mjiPVogIQ/eJCmLrH2
Ut6soMqMS0wsVXKvbnn+YAYb8gJp6fIcl+bpuasg8XjfrospoQRb/oEsGtGVN1Io
/4Cp3qT7uHbsT+57sKY02PhOagcQkwh13cJgZiIt3//IolHQDQEMvSqrtNmWxVg/
WUAMEdRxGDVEXVEwzyORdW986Ovb/oRzTkoHkMcPrDCC6B2plSOMkrkgK6JVT1Wx
e1FofEZsEMh9sYxnRR56s8H/gsbUR82vV1sivKODeNHUaF+qnFAwE8x/KnPAz86A
BaS9FcpHCTp0AtRsQ3sLN1G4f64zUknnJSkllfb6CeZD5rr6nKD3FDTBveXv2qbc
bdPUPMRS7UiropVgvOVEo0ii9GPwyUj0HJjgvNFjzfI6/eqMZhckzUO2MLDK4o/n
K81A6lryTu+JtdIgbrIuSdF9WsXhDubWXXCkF3K7CQxURbiN47JExqh3neY3r7w4
dOAW653Q7M2ZSme4r8c6X3Fge5++rDwgEg3qPVb2harD9tFfH5SQBgpCawJ5/No+
L9UDGT5kXeyQEGKgKCNnPOsFxGBXnfDZtnTetehIOp/j0J45fK+WzCe03chzMv83
MDSAe8ynP6MsGwKIMQI6W1hLRuYaXk7EcsT4N2Zh3tKRc7zVxl30yMKD3jPAL+LP
SHY8fSiMAc9rcp4UL/fx1TkiQNFgJRitq9FohDrLuo5+fNlAfABDjiiDxTycwXii
2fFvh79eW+PcPvVpNMVCs4IycrlCKMoOvr+G5L+YYclRbpbp/5c7ikO3opyStPhk
Fy4zq8uwYclFPP3xdFuuPiLYngf2hRd1yVxk3/cEM8Ex2qxmoddZAp57XHLe9BFh
8nc0hGTcE9ZReW/PI+ky3cbERcq8u3elfgI2/v/LrYvsjPMZHQRNjelj+fxJzGE/
UtjxUfdUSajyYbC1sTdHamsQo9aRgBZ90sfvf6XkNrG1qtTDdENMBL445ykZtCrT
zi8AC4bXyOIPmH0eGkIhyfbzKsFL7pZxYBact1k553eX6yiTgVNJMiOTMC/ok9S+
oN5LLlmG+2eg634sQLge6P/cYss1cPjN7kqzUgy9M3DsabEgjqZmA+NT4TpJJEvd
mfMMDz8Kxi8OzU1PtLxOQTbVwSD2mvsx6IViKwEqp9iVLrOusJFHK9594vI3nd3I
6s0dqgZ1iSFeBYPRGuBnnFrrZse++M1b7ikvlcpvl2DptoZyEnRm7u4ecjODWNsg
6Z4LhexP1/zjqA2a/5soe1mxDprjVFGdMMqGrJIuf5afXdRLSUWlzqS/osSdU8W9
tA/lw5qca+LziA9iVMtNE3PeSrKJgs7pYhZHkio98RXMLiHWtIApco8Hj83I9ZDO
7t6TL5P0BpTlAqTCFz33xyYjQApllgw6QuYnYPWDJryUbvQp6e/ffaBChReDGvTL
wZEpZlg40dmlQ8N2TMl3VdGkoBihPeruoQoqbhPh+sn7qMQGGjQ4Hy3hJF+Va86l
3WrCadc8UfvM7dmblUSjPyRlgqWs1WP+oi39zAVUk1ZFpO4nMuTrX9aa/KEf4v4X
aS9vJC8eQveeUM2VJQzSgCFJsmN21d9ZpOKvlucQ+uuesRpa6NOicVYAh0BIeRHz
DmVa7plyxu00nSDKzMqDJLu/tev3etLWNQvo5BmJ2DiTW/eVkc9zy5+QOtDLpPth
qWiUVKcJMMOmIX3hrSZzlDSj7wWTIzNsavctTpBakOgfFLPbCB0QYxpsTRRCMe9N
LAbqq80qnPVWRnKgaKESbqaHQGF4D4Nvs1Rc2eICQxptCMCbxdsMAZCZA5HZW8kk
t167J54aJPHYAl2hexHXi0TPnKWunQNwT7p+A+hDFo7HKI8IUL0ARz3yfR6SLLlD
82D7ZmJnqm4hRgIsdewwTeN9bEfAhzwBpwbxHPGs5THgVyDk2xV9E3xq6K9BCEFf
dCOy/kSHeSw8ZLSTkv/XW2Y6HZnbufic538qbEYOG1VlTf9Y4v8nKVBOQncfknba
MgT4Zos64vzJcSubJMYVWL6hqJVxvnBgNxzIjICJWhGMr3y/b++/1Yjr/8XCUlnM
e9t6u80tApXQFd+6zT2kKdPCux5pEAkd6etJPUoUv2Hq+pIWtNi+xeCQoTdbwNWw
p8ob7e5M3CsCD2BBf/VxrGHduiqSW+Fm4wyMd5bPW/Et0UkF1vZb1ipjdBkOWUCg
v0/yzH65Y593NeBmUesQl5Hp3jRUicoR5ZuD7y4XDvIWYyDDS40PVI1GMgav39k7
w7qYrpadmn1XM/1NzPTNtW8zuqxLGS7a/3cEQdG69eOMKlNMZ/0kNEUxLFpJAsK5
J0c33L2QOjZUcEk3fOTSI//6Iopw3gsoJGXAdgoRDiVUxXUa0K/SlYQjGA2/uCw8
s1OTT/7OxPYcdyX6YquzmUnBRdLWRRyDLEF7aQZhNuKELoL5oDy7WTvnylpvl4Bl
Ux89OCvL6iSdPOwTN+Y8kcXrvKpKkJiCyfpNtGWm3ZeTdPW9HF/uj0Dd7aIPzCX6
KY0Ljy6BP2cPdsTbF5NS80aKd8IOIikGdsscdaUHxDOnlpcVVeJ0LWZ75Rv5WMgT
izsKZ4zekdMy9l710EKv+DJBIRmxIib4hTPSi0YpXiFYdkSHuOfE47fjgICP5Qro
956c+2vmh1lcsAKeVaRzBCvi6s9yIaqSpyAEa9cRWb70ViNOE993ckzt8in3cMet
Y2veHuEnp2z8rH4u76npP3jz9WFKsEmwF8RTNfJhOK5TtZ1NAyf2lW1YBcku2gwB
03qUAtRr/k0foRiPyRhz4j2qtHzbM5C6TkycNOh+W6wldeeFrQCbsivaQiduvHHL
RXRkkp9fQge3VHBdbqK+0ahQyUkeilBJgs3D6pHqhCk0jaDjOznWycwrD0XP7Ezc
biwK9XGlYX5ZmkG9E8PocBE/O5HjUdA5EUTNDX+zQdnFJmaIwuZIeQdzVLyBOb5g
Gk9LZYR46luMszPprgPAm0rGKNuIg/ZFjrIHbi72I7ma2mVLQqR48nBDq8KzMxxc
Od1Ck/cT9d7UF7CqgtGIw99RGyrTemtzNs4wwMfDyrkZY/R7PPNBzP3CSy6hh8jS
k3Fzy7f0ptsaPXKLUC70ChFBS4dmeCabE6tPcDWSx3KmWJ2BEoGTtc148/IPRvkY
1rA8dEvgl6odc3sl8kAQpk8UNgvILtuzGC0iolOoQLQYCQLlk/CQ31SC62WaMM2V
cTScd8cewlwGXgQiNmw4gZhpY/F9O1zM6H9KnZqlwtFPo52JBl5wMQ80kQ7TCbMa
wAmA5MvN4ujq5lWfal9Bgr3jiZ71g4rP4cGbUgmUcCIqnUfCfulHixFkedNLpmjz
Ta8T1TQwmERlBMY6m9cvYxsVxEcG/04dpCBBIcqQSpsYeJPh1tLCbWl7U9TCeUzi
LX1DgtsMz89NkDJOJ7ZHoXHpKbyu68WXGgM8bFPVTH6GMSyH0NX1PotBryUIt+XG
E6450gVGyxNqvCse7HIpE8V0b2uCDBuONFnBVn2Xljk/E5sO8mJLBuP1MpPnJTY8
FYyRsKrd1Dt8LRFeoqVhzP6e8e2egruKd/9EpX2qHJNGIWkhrCTuKgKwlj8z0ykv
X5lQvIMXsE11WS8dV3wu655iO2RJ/icgOdFghF3KMWoHZ+hrbabjv+/d9xQo7qej
6gW3vDmQ/zcFys3HVa6K9SLXpWZhciDhvmie8AFOuaw9v7/GwDIcM2Eks7dtFpYV
RLQgvwOhFH0+WJEP2HleaaeiN3jiiu9bqfgcc68DsxjulNQcclC3XfygfvYjD3bK
68aySGUOByz9P5OKSARORFaw/4iYfQXVEat6yaiIV5u/L946iZZPUe/Vegna5UUm
gmyN4XyGh+kLuvj68zawjQO5ECTLxCI4Ydc9ytyXVC+URYkgTSdQy7reflliueDd
5huECZmhm1NtAWk0GFBiAudnxeOff/9OX6Ns6jOmz/QXUbmGhP4yzYu9A6NZEwcS
k9R1aI+YYr10L9h5m/0BttWpxE44rEWXQWiujc9px6Fd6sU/OJfdnQMF/kGOY0Li
AMKMEMe15ozZ1vGYP+AcgIEaPnzR+yl4EUbBUqDpVz9XxJmXSv9JUIo2wjdKXHw7
2Bjgki6EZsBnuADxd3vEfrnPSn55Z80iLw/2AmmlRXOdjLlW+yS2KcOufIGGU5N8
vq4IaK1YVbrYaLDjes4nYqHuGRGKJhOZDNgTPtDikUqwCRovgBQJYL2+j00SFvLE
qVXF+MBvcS1J43TAHGSnF8D6mkC5pyq2ieykvLnyyZMR2qc+jJyiU116DZJWfspS
0RAo67mW6AefwX2L9zjSe9IeLgD0DKqvqiSucLtCO8hK78wVkq49nBPdm1b7Idi9
mFWLBotSd4rLBLxKWZFwj0VuOAoaNah19qGFg9pMHpeVFYjHPVNe9p0Q6inXXG01
AwvMVmMNCKGyJKjcxJkIo9JF2lOOAW2ANSgmQHAf9GzdTn7lC3M0Dw26JgPN54c0
SAYG+NVYSOdGvqwwcB+2Lac2EdNehmFKXeADzvnifRtPP9rjzkBHQvO00RfOTdqr
S7xZQqMcHodzwmVjnDGjz/dIF2qhNVaU12kiQFtPuslUeBxB6mhOvCniOm0ltKeQ
E2YNWvjRFZKGLmMgbu5xiyh2iA8ZSjot2ZSBHCWV31sJY0b8QOU7/cEeBzjJhzM3
/lOt0PPkMDEmrQynlWG15qGl1DqxZgDM4703GvzHP43XC7B1PPg1yER+fDD2kJet
nZw4rNtmIZcnAAd8Qvh4kmbrYsX9P/6uj3W2JRDNJCShSq6BzwZAct4HUHlD8YkD
KI/n8QcvYpiZU+7B1PEApyt4DD6rZBT1tOmCO2Q82Z70PLytVGyJ6soiPXMLCiVA
KFNQPViy6TGHYJiM5l317+JRgFmXVHS2Vn5Y3i7wmg1tqgA8X5xMGRXMQixjIOWu
KZEDS46cmbWAoq4xbgcNQJuXD+4i/8+WZbW8gzcCtvdPHsFtNl1/oB0Bldi3YyK0
aGkuLdBv+0fnVu3C96T3v9aCHFpTlGirgWAq1BN7N1TzcWzIlBS91ii9VHbMjWHa
3lF0ZMviCYKUYB0f90ONzTuqrXgXyuDXPR2qdMh538GTRyeqPmojP3Y5eJmcy7j1
fGG8EjwB+PsTITbpYtH0s69xE57uzV4k6koRiYsnFFd4bOtIZR1rgQ2Dl31MdMh3
kNN7qDO02KShtanSn+4bHLHAuSoIzHcjbdyzEUgo/eXtT80NtUmEhdapq8BeZHwo
MYolgCVX+Lvpvka/ILRJj79C6ZIohSjJ4g3nNsP0BbpPW/J8WtznMb/3YQUTXOhB
kheIIcC03A+a39d4cBpst05aZDnEh2yQ/3/DvG22q/mpcJZ+s5fglgSfPwsnArBa
RldRd3k7S7e+9TpYTwQyRhvT+rJALOq+nvrpDNFoy+QGb5kqZMWkY3UYgTaYeVn1
C9jLlq+DPDkGRw2vLtL0XXm7Ocgm7jSqhZetsdmYWwosoVPVyknf6gxcEz3PIeeW
wzQTll61F7qdWdInejki/BCxoUhU7W6TJX/w5M0sp9S2EusmE2ZIumzI7HF9nP9G
0qoZc+HtsZtmGVfw1IL68L41WjPUdP7hG0LhHYDqSk6hX1fos1MXiyWjvEAgf4mf
KWO5HN80aSjNHLVUXoXi3cFplZP8m04c97AQcAVX39Eg0cjPeUv+n/3eCP4mqc9H
FKYeqvQMOEbQGgF4d1f8oEyLIoSRC/muK5/kMSAMio4L6Vo+5iWlDP59Uzw7aRdE
tPaQEgx8dz8yf09HKZrT9L7zlZ6AnLDbQG6CK0CPEIq6mGcpA+pUlOi4nkBkkmuh
7JNdSaXbEXIsqEcN8sS/unk6isBTNabkRRjka+2Ah5CS08U8HBZuLqUsDnHmexa0
TxlBvTCSBwhTrNhhHSvvsq4lg/RZ9O4+RnG/Bxho/2i4jnG8WOsXdOl47wPp5Gwi
Z3CMTv0m/mTw1nxQLQlmMGta3s29vj0tbwTPlynUD5wMWXPI4/qJW7hHYL+XSrBd
0ji2sE9LV7ar2FdVIRJyadC+MpgxqOfLda1jP1DvdCeXe0q+jWn7+60JztwkQdZL
ezFZD+HysiFi9rbfoedZIeBotZ87BlWWuevbDIVWnQ72lB7QD+NRaLxoz08aOwTt
v3IrXuM/w4voX6cChe4geMHMQWwtBvldeT5WagcIN6hgGB9C3iCSns5wQrBefKoh
3F4cba9HyCAC6tOFeeO2udSg91azrcQnY2WExNYd2o/TWnA9KqB9+3A8BY28KCLR
PL0SSiXitampk7y38kj4j0Pyt2+vROwjzHdWaev7Ezrwly/nWF+ijHz9yKlupwGT
i0wScCiPK9m1SvTVjClekGc0bXl1eyVSKx99BuP/J87j3gsPAOhnNfh9ogORAff3
cMd5gMORWvRCl14Hv1qF2nzEO1PJagYNsTOEHotm/9UPnEBLCBQI+tj9ZE+y1J8Z
GElSsH5eFQG0luln9p9Zm3Se5EruYzBDRNWwdq3S9gwD5Bwe3xgTqR/v70DxOVgb
1fTI8WMfAdPgoCekaVPlX+V9rmweLiJr9QhpLW4DRCCI4FA2Fl5xNVBk6IN7UBy+
UB0Z1y21Ep2JjmaC2RR/oIRdMHa4/nFxjhRheh8gDgBk7+ZHCL9G+AxrZPAWYhzL
GdzvU6vnhtvR7Sf1eptYl/7LDEgqw4gbiy/fODds2K1Miw2SR7IeBU31omNteYV6
sdNg/ZJ0t3somgFUUtxvA90P/4kqlBpRKdAtr0jTvLWUbziR36dgO5PxkhdA5aZR
DzP4RLlcBM3sVJOSHBEltRw3pyvn4DoKWiwePzxhd3bmYoDcewIcWRBjPgK9UvTy
1iQzA6FAyn2OAHthk95B/oA3KnLWP76WDDDwDH01XeU+oWjtoltAM0NkGPIoFJiI
Rm9p5sGLdHYdwRNA8tbQZoToW2RXauLoMAbfhmMvSyEVD8hS77lB6aCA3AV/tspk
wuoMa1HTbp7OGpdsfLr40B/M5EZMe7PjmklB2GOPwZGCTpbFzy8pilvC/nfU3hpL
xCoahcCtrqHxX8POhvNwrDRjGtFzuxlKGWKQf9Lr9lwru3nkWPq5h2vEwl1qwY0Q
2PGJdi2fnxi1OqFqgTQ9hKI+2BGpd2MsyredgcODuPzewbqH7UwS8gFeGrkm0Dyg
rakB/+07VCJWW1ad9uAqGw==
`protect END_PROTECTED