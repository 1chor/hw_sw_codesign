-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
S2SQIrb4VnAQVX4OI01yJHN2tY2h5IcpeuSb3sXJfIjGGUSN1ZqhGojwHuikZUBo
gfTgLzzUgEqs/7V42wXMPR5EZWhoF3Nzy6FixzRXMRWKlq8ZtkeCIo+fFJERrjaI
AMFQ5ARbLNbae1V748OLvktuJwuo9dqViyIiMEMKKZo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 99888)
`protect data_block
+5cgXcs5r6WgudofmEAHrdVTHOD7JPkuEW2c6WXdd149jTV7+qpMIqxQG3pTso7x
QfOpb8n4Rc/zL+dUzunAR0wm3lb3a171te2uBG1JnSst4XCfh7pPx/vSYL7hXemx
nejbn+PT4rLDF02deSaRu7HtJhCTaWtZq3z8O8prPgwT1u12MPKUpAoF8mW4TSyo
i1z4nvaIKcVRXAevUvuWeIoQYObg/IqLdxhRwCDTS7mf79mOfa+kG1eb06nvgv5/
y/56tRd3A3FEhHyQ8NXEITYBWubff72P4YrhcahzRm5eTCNVwq2fCxwfLTXSCMQT
Z1xf9bLVx7Q2HeD7Yv/9gt1fDKbjEeR7Jer+yXKFTAUnnfNAXJ69CL0n98YIbDzZ
OIXkdFWSuY9VEWC6qrEG5X+gTdgF3HMMne/8jVa59p+6LrH6DYG31RVcA0ZeYW6+
zNFufDhGbja7JkJFJYAUNVtW54XOeStzZGW6tWAepWWlIY7ZxqwW3ElNrWq3yrmK
LYeAuYhcsb/up2U840UE3d08n3j6xwdFTHJZ5ZfEoXCD4dkuggDGH02q2TxBfDe0
+TIa6drtMJcZBGxisAFXu3095QflLXmvqAVFldJt4E+vo2DDi3J6QeesE9nRj6XB
X6HrAtysbVcq4xAopPLu/AWygmQvsjngPXOaOch0y0G42/UZ88TKjn8UjroWqYoR
JmpAMT2qVtT+r+Vhx8EpWPCbEsiAGbVBHxuWVAc0e7EasGbDAnK9cRFNE5AEBHbc
2Yj93UHvUvUEJKIHHam9hdIgtm28HB88xVlkj0TqGvjAfLwdZBsJJuMAxrL8ury3
4wI3fhy5HKTI9oCQGqCDBRTjR5jlfA/7ZU2wvgIc5aPayyGpDSDQGvAZefwSvngo
4noKYGXfJ4WR4goh/5KZnay3yK5qA0w3FBP/ZUpZiBzrpN4RMGsnrGVp+SK3gAlx
g8+VnwUizu4yAPVY7BbD0YcK6X5BDozHbTg3x62QVkrbOh2Wn6yCfXjD4YVyC8Uu
NsOtTi93QmgDko66G2lQ06MsJnWQtj1J0+E04suZSYaQI+McYB2qA60XdBfhUPiS
L9puAs9sqZRhct+A+XzHCOiLZ1rpfwCg7aAWAb6jaPnbNlPwasp0A7ADdsRDO4nr
NBIvP3zCd74A30ZX8cGqcsjmhMecX0Q6AwEctlAYqP1ilvKV23Mj2cnw2AQXZNmW
04zLbtF2ipAdeegVdUewGUvpyiic4M9kfLT+UWqQpTv6SwtKJikdDeeTYFZGthRx
X4cdLtnoJLpkpJ4lxQBrZccSvvofayVqbfw4O89/MntUkAFYZWaiJG1r1C7MIRSe
qGJC9uxepT1F/MaoucqQyHv0Givejr9XIdetF+leiixI82AVtiIb2bqByZ/5Zf+U
cQpVzeTz5BKdiM14f1QYR73Xp1mB6J8j8LewSKGFXzPSMVhjIcP52imEmzx4CuCb
LYKQ5YNqP/0tq/GiDmrGlePTpR9OPQdteltz75Ry3zXi/mt3Y/u/WJIMLeLT6XP7
qo5k4F45cqbOaLl81V2iZLpVjwH6r/DDpy+P2emHMIMkfkf7axNFT4/m7FKXvLtC
RvHpEOELrq9l2IBxRgPdbWlNSuCRUteQd41a68xAEjdPUpFP9UD05gHm6NMiLKKE
oepOt6G76xaskMyotzMUfLED6qRW7CydCPUqPx+DQLRB7LF75Q9ZYpPzZsYHGPzT
8RuqtnqG8oiIDlZBI1YJ9vCNUO39CZV9FhJyeMhLYgXVtuMLTjC/B7ebKMCWIK//
0WlIrJHeYjbi6lkrLKVw0RX7FEfmT3hBYMCwG+1dnNxtGhLi6aLibrXROytPji6w
O4PicZfVqHtRBzQE8OUUBIxloSmzGKdzT089OCtzuyHPLW0wo785UvzAONAcpNQH
o3Vv0/bo1fuf4NJx+wfOsNqWWnae0kuve1fO+iz+dfiOWVzj04h9GIXvlSXMcX7d
SpCyP7EC4hV+fYtwCg7KBNxGeI2WAVg5eNS0tXcLVXeEJKRzfVIt5vWp5VW9arpV
bdw98yY22vamNnAZ1b4rcs+QJxXIl4UeYXlXtBY6E7Xyoc3Io3vt3n8jN6eJGAhA
+PtqKO5bR76ls5al0f28EBXvKGVh1ooFo/Z1Mj4gR9jU6LMfCmnrmKfRFr4BM62q
/AADnA64FMJK8gaAIarNr2Phm4JijKt45mtPLxvB6mWVS+IBB3SYPTvrQ0P5Vykb
NedSomMPb6eV29B3VP1jsQyRg1sP+OMbDA/1oRKDoA0/06scR6HOll1Z3Nhg8EI2
14WPMfLIbHDk0G3T1j9hjFRHLZQDqUCJDeItUrX/UuDiZ19obN20ISib04UIxnny
GvmA6gnMDAgWvlIEu95GxVW8MQPCf2tp7UrQnEA3RIkVIEVeFxJMtL7gWt5UXOTd
Kkzs4Lx81ZjKD7gxlKmIe3i4nW/Qgjbq2ggAImVHKj0zZ8pMtnNTSPcP6/SNeYLK
0mFGHa53+bJ5qthKXHao5/t+GR6f1/BrUYqBqmZZw8VAdsKd/efK74MVX1eJ5T8S
oNUnQTLmpWvucRa9opvj2XY2EmDsiyeCSSQyab3BYKn+/TAP/0hq8sv7q62BNThr
JTDuAKaUdyXnCRfnMTB8PYIwTCrENZ6l3W8PB9DK8WwxuysUBfZhID/F6Z8R1DLa
YYcOlGs6ugxzbEsCUkNnPPqJ84m72T1EU/FS2Yh09xuHWvx4pET3xWvjsOLjsvpb
F/ivZ/zFhy5905vs/S5fYMFK9DilYs6odSg3CkpxHxOuDwchFIYkht5M6Ue7INsE
lx6MNjhfFNxqqbs6lr0eg3mZP3NRNU5fgp3E2r49TKkQWVlV8C5A7dtDDfysZznR
uTyt5p8gH1Fgx5yrG8ZJtrwKUu0twVjSyBTC4wvEzC/FH+Zr4tvM9u3dze/H+hfh
VYPNYr6ZrKxI2vDaMqQUaYwx7qVGva3jkFWLvmoL1ahZJRRayVxlRWwq/t7gV6ab
tetKDrozSOe0uYtrI7KJgGvEglFQkmp5U42wlv6ajORFeuEiIFd1o5c3mtJWrL2I
ZwfLw8mSKYGlQL8Jrcbh+K24S0yj993SVTmZoVV+WdSnSsUl2ng3k592JC51Fw/m
i3YRbnzSEB64jxnyNgy/aMjTu+3Af3E/0EFlXe1++FxC6xKrT78VnQtvOBJzMJCx
mcAtfKPKO1/cCYrrVbfVvWRA7EWWgZLdHMsyteAPV1cjpgg4isL1atMS5foCle64
R3OJQGrTaGQh6vCk1orrLT+EJTbfA7ztmHKhGM0ivUcU0381+lMPDrOvNDpojPYO
2+pp6gmJTrmxqYZa0tJmubNIgYt2xlVhdTeiPchm/OjcpkiZ4cPk/qnbSRhZ77oX
FsbroGAwQev5T98ASlBJaGjuCh5sIB5mfPufiDt4+v83ifj8uhxndU++9zt9XdG3
okkB31p+gek/7qlRwSYh+pYdkQYT0RB2oNuG6MlF/8VJ7DUPswbBHn/q16vVUbWm
bem2kYHsMLU1oIBy8oPNkMstkAhz69LowvKxUOdnulEScNrtgYpAua2E9jxVV2+p
q9oEVOxugLBmFHsVVyDB254G3iHEfVz0BZD8EoWTx2JaxlM5ijZMk3zaxHwHnrLJ
ndsCHFe6UgMYOgYHGOqKhUc3dpwBf7zs4AojklXzu7wERegPBWxjfezEyUKZerTw
EH5Q5KF93PyHCdPU3tUlGzg/eZXDf0WKtPqojq5m6//d4DikDyuwxJWwtLbUzM8m
CyBX/QTqCBKSJnwOJbYIOBrM3OUJZJzWuj9AD8NQfUwbSpnNvzJ/Wncc/RZxzlsz
/p2RwofKomoi244CVkebyw0v+SFkHPkZaIQNkW9IddDWUfcGUNd1tzxKgTTs/FLJ
rE8SE6Sq4XYjs0EUyxUCnXgOoqmoc/dC2ICLlIC8MDBP0m724KFtbLBtK4XCVcHh
w3XzRmzSanStc2d4RBSejOnKq52ZhzPnnj+dTnUHJ8sCIs1MeS/fgTIVox3nRKNR
RkE4z94nMHQ1llMOwvmshIDp38S4J88/dOKn03DwGlnuOGbpUDaikr8Dl32j9cMJ
zSrHA71RsUxSAUnTASSf45T8AAZH99tL3eNCv3ERKPRvyCjyW0BkaGFnqlssE7H9
UDikLjzXPPw5Ir8qxjn4uHmlT1BjGroFco9OfAMNf060ZjE9hHU9RO18Bh4zGqsg
IePo3u2qXVqAje34ieir4TVkpcDEQ+q8OGF+ZfmQiSk0FgD78e8ykkVClKr833Lq
7eF3OViGGkFm85Xx2YOWt/v17NrmNAoH2Me55UOVNEEtf5tS9sjkkJoMu3+8ECDK
zlnHrtcI+riOU+7106/AZbLHbao8Xg/63/7kgTTdQ9kmNxKGgSTJCWVHhwsaMRzc
yxuV3pV5IXsV04PerGWsU6z6L0if2KSbEcpMaBLFMQevUUDNkUhPugjM6i4fCXgH
h58lmntPXHr6xe/BKXj0RjYzz3wtKgsxIVF9f6PP8V4sixRWdWyVr5d+D1WR0Pdt
La1rpMgC3xjIumtFEQiiCFvmwGh1tR91P4bl8WC4HFYcK+oghf6G9sDGmZYqUEi5
gS4aUtFnfdeNOfQU7AE1gIuqX6qWa0IquSu/3Ppvgx8m2PbBaCtUDzbnpAnu5eNG
cenonZbDMafvEhni9JIOV4FUug0L5dgwaUqJDzAUPYHhAZDeziZ3pfxFgYNUgewL
6GmQxINNlTz8kj+7gn5CXr0n6FkQMuK1zFK/xSr4jdJpjk4/v0X4ZBGL8zBJpu8D
qKArtCH4nEWEhlwcvCCznFGdTi/EqENuVelvOTES3+PEf9dtg+N5qHBWO1YyMiww
OfgIdVp0tXGD6ufXiE1cNW3Sh8/j9/vRga0cFmEjQq9J4yVFByvG/7jDWKdl10Iw
RSWBGH0GGLC1UNNq9oh7zR2OF7rrlf+EnOzjenPahPXDf/O9FllQkM1UI+eMzLhJ
QKZ1dHzRhyd/4HykVulUXE7gGLIAArLTVm173Ro6/W4N/elbcoNJQwixgkQvLFjS
e6MaRIuzjHrv3FxiTU/czHivhMeiptsnuIiGbu3moKmKhzL79cz5g9R1mt1DEaHw
lU6/6xgo7XPy4ATEVxPo00oEFaKPdQPofImGxRYhIfPqc+QDub/oy06ToQMHD+UW
5zs9pbeo/DOHGNpq25XGihXd0uC3tML58s8TTtdBR9VkzZ4pDeG9YTGo0tImkZJ/
VD9sYYvulmCcrvDqGGTNUjqWoayL8xOHS1I7hKCy/DY0vc11LaTxA0wxceyv8IaS
pgRd+WuvP9bqxFoKOLSXqEPI2da+55gmj7OYw9KvnD0W2OJHU1vwQpFIXQMSkV5Y
uAxqKkDaQfF4IGWWHZa7juT5wVYK0RIm3/jbkVzhKZ8NY9eqBWedFy/DKS9GDaUg
k/bTCIMOnRfPQAfwHhS758HFThM6gAiT+R+b5HTM7HHTkVSxDZ5eQ1jM2n4e9Ojt
qUf7TQaEQBsT4uAjSW/XSHgJy1W/bL4amOs4rK8Qe0T3fKBk25hwbY8trnBuU4TH
HxDuVv/5EhXyDD1AT+DNMmtKayDITzep/1rAJQYSeg9ky5oyxtpYD6gXr+B4ql5U
RoHJqeimZDWCYU4yLg3n8JJqi/2Em4j35LKRRwZ9fKQxDJZZSFcCOIBWlMnRGeWO
ivMgo8LtG+bpS1y/Ss1/8XOipDTHkDdQNg5q07I7nUsdJzEiT3MlrdlDQuDW6LnY
Tt420VDTr7ayGtPLQfjM4fZhyoWXlgDJlZv46ysbBieRFZmsdqqky7WbDNOwl8Aw
cqY8Nfh5o/Yk15Ww1kMA27GDZSk5oEPZCF/uGOGYtxehi0rJmg6g2an6L3qJUjDy
kruow2vWZSv+ZN4Zo0Rzu/tOhO0jLPudSKE5jwgGvRng+V++hAC+eW+RRc91iV7v
/k8hNEalF/eMdUdTq/x+g8BczoRoXuucJU0Ax5FHhVS8cUiV6SJE1L+L6ZsC51+/
kbeDxdt5nyg1lTmfv+eBGxU9/Q+tng6yNtmTYxXH42IeRXXu1wrR75uvfq3tJZYE
0CKAjVxzPM9vypwQgE8Wv6/Mg/kvdB+9fhVJh+/Af4bEOYinqUIq1pQKTpzzbN/A
doLuHg83mUX/LeP5qK8uxf1nv88zcHfbZgVitGaMqZpfYgX9P35mgEKB3rkL1+0L
wa4mrF5i6AKYRVN1QcseQG1FJA3Xf2NG+0jm20kNKUTeZhTjqEBfTycQYZ2NX6PL
dbKqQhLtjwHLKCQIpUyTw2DG2dmjh5RZu636rUU8sEPZyOZQvhSAixG68v4iBxw+
/SYKD4AnbQ01gsjhW9iAS0i8s2PMBV9MHkaafnf5bo33M5x57L/KQmwQayjOL+oc
cvozKMe3wi7/d6GgI4t2GLY+Y3PMlNtESvDrToX+9OPcwubYE8Ei09uFpt0KI4+F
4EpYoKg0JjkZDDixF/i6xtm5yLo0dfrqdIWpBrjkdYgXnQXqAEyhBp/Mb1hmSovW
HbYm0ypg8x7FmaKBqXmym/xwVwXfkQ4fL6CBxOJXBQtpiepMzrO+YS6PX2vV0+q7
ZvZOFUIP1NlbOsbSlhB1iwcm8bbsMumjKWaJqc5qamdn4fexafWQKrdbE+g5Kp/k
si1ZDVQp4ZVeZdMS0Ov0witmgk4ridWunY3S7wv+L61Uz84hHguOcQ/MnL7ycVvf
6hPjbGJZv4WiyJpEHvpQP9TFOmcTGVjtSOJHpW4z3Fntjta9ebIzuKriRfKsZ+lw
Erlz6WYTTbhBRpIyctgGgaBYVqZLtNtq3iMsD+B5kVSQvnbo4Htxz24I4vM11o7C
RZu6T9CXIvpduHjZfTJwCMUo1RiWZS5T1afONZVP6ZuiXDZ301tBpjDmldDQPUjd
o83fvmCpdFQQIkNArxI6sNNjBLBZc8qE0FiXQxBWKCH0fgIEJajuczLR4dKfQZkt
3sUObxZJX2cPG9wDjRBtUlt3cIK6PGaERDUHnVkRZGPJ5HjSSlcO4eTSh2eWn0Lb
YP9YLzqOgrB7pIy+Rodzj/wHHmozAM/qXm+/az91FcIeIw215oTWuxUArBiY/uJB
m72zfXBF8xoFuYfaIag+mODzunRAVoL1LiZ5kPwO6YTbCXOv8lgLGMwbO4oRhWHi
15ztVJ0dIQJIPFkUbBnkoa0rpzeQ+y5tZzYfTv7JwZ98cefIg1zPJFNduczMHU6I
Lg58PVv7APSpY14aMPWrmaNONPk57/MC+PBNCoYBYoN+dpYhFoJhwDnIUdT2Cl8i
1ZrE82LRtrizFtz7ZMHOCy6q/9VeDK/HFzWSYpQo6igqdgBMx1+eVK6a17qWq681
FC0lNdoXTPH+Qa9MXwAEkp0We0umuO+xrrs/A+Q5VOInXsQm1MFEUm/uDFtsktOJ
lz6V0DxKpQMjs9lnvsCrwvPkUeNsQIh/BneV2UJL1U8OMB8uSxO+ASRm3USU6UP6
r8pYpGFnP3MFb89TVFBITpuC9wggpSslITFvt3UYznO48CbSlTTNiF28ls5GzVxs
v6LahBhppsuwvl6p1IudGlHEbpONtvX27nqMXQdwrOgDlLoMbmdKX1YPqcpKSqIk
5gLkvN6Ag+pAWQ/9MgvFGKe+0VcRTVwsp/HDGExIpqtBHmEC7kHd9nxCdONPvuYs
i2K/xACy5i9tXxYenW2CU0K9dJPuxFrkF27qGLIIPbE3WZ8M3sChsQHy/VF68g91
1kz6Z3Y3wFo203teWyXHcr2fexKsFwopEP1EOF4TN61qL22vuxuSABFKGIorFrqZ
YTsCOC2UHnIlGYVopuPj2sRxrZr5FCFzcMe1G+GNP8J6GSSfGmz+aViN/xM7tt5j
aVal+6OWvsmdY8kGoS58p+6+sa/IeteQkxhPQ4N2MNlRD+Q77KRxMHL9j376mCZg
Tkfgpxka2CkoqOEzn8IkQvgTLpavY0w0p7AbMJAQLnf6DhPhbUdJnv1CuVwt0h8N
2EwBL/0E7tJIYOTe/KnKrEof9O8gqsVSSN41gmrl1PUScTsJk1zgeC2L1XeAyKL2
K9Nzz3bYqd7XhHpQ1p/gPfVjcwaMV7MSjGVoAroqXCmBIqthqQCtORcuXY96Q761
TeNtswIq1lHVRZ6vD9urX5KorICKDvhM2RljNX0uwdlKAgC2KU/WETb/ItuzYl0R
5r5a4D4oOz6/mKbuKsI7Mcq4m28+RnRq/z8C/oavmB/9as4ji1R+j4MQCYbghsXx
y/FTgadBY/Y3VBhwNTl+HgDiCZC6i4TuqK3LNNuMB19ocbW2alrLa2YoXmbQUkuM
5JoPjZE41xVEEDqAE1N6O21gD2mLqozo0W4pylmZ5ewiBga3GjCXcD3XKmQ98me8
XHXdTp1/BJl2YF9ZQbjKlvsamdxZWzZmHJ5Ov+U++6tFeFJ7T0+f5IChEDB+9o8w
IOUmlI0LwEEqL/L5HMd6J00oicYgk9EfUL09SFPitlif73w+5E/lNA4vSmQZMnBR
oFbDh/Pq2rvyF6yvDB5QW2Hbf+0h1aUiKTa8+HiMQas9wYfDPfSWA7YXV62RoV5Q
8MwSc1ZdQGnfACexTvwNmL5qFCXsAwKkaz3TyWB7hgIpfsLaQaanbX+q5ptgv6dV
WfYqJRQcbL3xzfwXU4mj2a8v4rswIODNUMflvtOsf+VIvZnnnlvbqj4Erq5Kq7Xj
/jgt7jhf1SJXtMWy6YaZGUQJPelu2qIkSpKAASjlWBUbxRYBUgFUQd11mmy91Wk7
SEtILEa2qOIQa76DlJDpa1GsHg+wey4huZ5aK7SEm2duXCXQBgqDcsDJi3Xo41mx
5gKBdxSQiIbltwNcPJh4ceQzOvnAFTFdvKePZiL3awGbvUYVf/lz1XkbjgwDKhHK
9SFoCBhifq/g2lHzOO0gYw9JYQVSA3wd2vCnKtEKimowzNdPDHV1wjMWZXI2daFu
A9ShuBTlHrCH8fhe8aqgjeSFdXTCKkow20TZ/tKBgayiK7twCQr6Bp9Z4OWFM/vI
7L4zk1jZbb3933FMXM/f2Ae1hpSMlFPtOQjEPoASsiq82/4nRsY6MWIksiQWswOK
GKG+Pigm5IXG2Kb/mJKxiPAqdNsgYmv1jpwXkYtfHtRsAuL5hnVsa+QGkyscY4ra
AZeSPWDV/314V+X9bVeimEYI0jbeEFESWTpfTRm2SOxk3NEmPYI3efpQxT4bFC3V
fZ8D/wTe32SR4L34KzYD2RN7KizSvjMCjXsS/s5nysmmRkgL7IyZaxRbkPYE2j++
d9pV0PhGTCWOpVdTbSYITPiJErTgoZBpmD6GQtv469IQB8H4kp8yEYzBy1GSJifj
6a6JBGDV/Tq8DyXj5f9rvvI2EDz0Fp4ykdcIX7imihQQqPEXDyFYNkz3gcRQDY8g
0TBA9P+qYytf/DpcdUMltRodL6IWursQtVWvC4LwdxIAdKHD8InrxY5I24zENoG2
FlE+BY0p77Zy7x0RBOSCYOM6kUcan1YPKmvIGAeLomZg4XYO2ai6aRPQtw9SnQ8E
PN2/ujd4aPlpjiVHwBeh8HCJw3gDq5pN8R0GDqN140uYTORqwcKS2lxsXWW3x4+9
tz9GeVUVSGyIDKm9hCmjsglezCGp+t+cRm3f4NPazhTfEmoyTufPxrfKyypkW4rC
diJUCAUySr8dVqafD6FrOQYn9zqhKMw5la2ql35IW+f5Vwe3ue9NJdLj/yQiLe+u
dEhrmjSLuhoDc1v2FfGnp/A4jE63ocKRQLeyiVfJmluAnO3L6WGZSZe3kJW5LQ7m
jUNc9hxDInmMHvt0aRGCNS3g5HoL7xNeJrEMUsKo7LRPJfnZWJRZhNT51mh2mYYB
QumomHC7Keg5aiqR33DVndKkIzPUE8E60e9XHUYtCsl0FXEYzHvkh1tzw/iaiec8
zq4xBQ28AEUuyXa1kOYSZ5+1xRsykEL+fNba7TBfywrYVHks97GOoNqKSc7hquYa
oA9G5f6NQgv9m66sMw2Yc+BnN8g5bHoNhLdOkxgS8C9UwsfeZoAGCHpjcOZVPL6Y
tIisL5TCY2H7N2kMw4RnKsMCHmtGyYN471SbPziLbhYl+JF/fCKwrUN/dDgQxhUg
h93amY5wvPPsQAaUiH8OzzFP3S04jZvsq7da1dg4IBkElI+ZCHilcIWQsXLKLwif
55fjHTwTG7DHup69+9irqsPReZKyIaJLlP3BfCYbh63RuGJrJyb4SSsfocNbING7
nZMuxqEbYKGpLhdSWxUorMj3ChPJJW7207NzcgPHRfwtaMau/x0tSioCXuIJXwNm
lyt9YW6S7C3J8SF4WovKv0qXpxaay1/ULscwxHf2xtnjppWrVx4vX9vlWHDGcY+7
+QgzZ+hO+OCM1mw3U7/qqcNZEArmeKNFEgVinobTZvfEbU2B//CS5UxQsazj90Y0
LZ2/4Td60J2PfA+vW/i6aD7SaDDe6BcCp49jzl4a4ZjLopl5mPLPZn+29W1GMl9m
Urf/2NnnqMk1pFTkBTlNu88n+rvMlO668P3UVxU3eL4/oZhXVRetHtWRz+NIpum+
S/nEZJrdzTOkltIr4UP/RGDkReCpYXFjttPo9MxqhB+/P7/cgjnMg/u45ofto1d5
ah5Hydqq5cOsl3IusBl5HV/i8TTaqjTT1/TIdm0daxup23YXuw7kD5nB2IDXHHQj
LQlA+ZIWlUc/Xqk2/WoSmPx9NKMcDsB5iywK98eL5jv01nMRTwOanZ3g4f3jtVaj
oKaZDR+yGYZbWlSQs2fpxiSaHvgrIIMP8M1ZyyRXiTEL7MdeVrT4A/Rh71VdWGE8
FI94VpCJw2DS+F3kGkZ3aS5JXbGNoQms1NA/QJyPO0iHtnt5WaVM0HwU9gH6otdY
am2pzwmUCNKIP8Fm7kwrGggysrFygDLKVE+WH4eutCE7sSvnbDbshD77aYILYV+6
0m1zwlKOL0KTrGCVpzoHQ+9xAL+g6WwEPqafFaQBm0dNNsUQCEelKVBXDG6V0CtO
7g7cSXK8/Bw+s0YEjBM/4I+1yRLTGY385oDVysu/UXj1n1UThfQcA6eVR0ZOrc2H
Xgc9of3mTvathAgrcS9YqZS7yKTtvNmXDV4dxidFprSNzoIrMLL/jD4P4aX7B5QO
1JyI71J3Epbf1ZlU7C9XtgzHT9HSonwA0tkZiHVzksqv2c1tyEN+Ui85vQPGu3S5
D5B9wYJ+x9KPDa4ESgjrPhiJ5+HfGngiIyrJKrkYbzSUrbQ5dpvGgbrlUCSeHwTi
4j7sDzoWpIjWQCheihwHrRapQ07jknzBPwQ0t1ZxjJ9HN8B5Ff6EwSiIntRPIo4j
lKgWCV8nYVsluvrzpGInsrB79bvm/6RVe49rj/MPNWmcCE/kQXgsUDl3VmwcNYpB
Nvs+a5ixfkdI6EcFxgBWDt36k25ohxhXr4+UBHtRPi635Q3Ly/dAD7Z3h1w31Ipr
e+YDRnGwVyv97RXaVb0VDCfeC+MQ6LBK+l+WqlO++jCnxiOHOEJJfV+zfeuX699j
bYWQ87ZuicXlCLLBlqhzT3yGZRDWE8+rCGNrcqhXR81MQ6dyodsdp4tIdsiC3U2y
uNKODKCPSp19MvnFHizO16NnCzuqOLJmyCrrvo9cHDg2rPYDxmCPcM/ask3QO98R
LAKoKq8YsrneWGFuiu6FPdmhzPQ0UqR3FPk2bpPEVhjAkxqRJ0bE7dbhadPYf6rr
dYigBWk0cC1s3JXClGr1ksBcqAeoQa6s7VKzmPU1by4RoUpM1kZkvlR4KNI2p8gc
FTCgwpmG3efJJsrCMg/DU2ZintgVNolhZtSz87kL3O3Xjo3MzEXNqYrxunGMGLQb
fOAUPhaotUShK5UFF5ouu8B72xpkOmlFyBLqwfAOEahdvJp0hcP30+wjcz9GLOJ7
L8k+3a6egTWoEZQZKJs8+4oN8XgOELq15NU7g+EhLn8Wlwkvj+A1MSWIkCQv1JCg
ZuX4D8dADzlTJEC8WhLWLiwUGyHyu+k47vbFjnG9Ek8J+dYuqseP/vQFgHH0uzLM
J4gLIPe+IyO8lynlzp2xrD9uPBm0y/WHpf8B/oc8i3LYBGzQzmk19jBHTrTn1Ce1
YX/1YviFZxQiJ9oG+MLenEgsQmtHVnBc/pWQB6OxdBUMc4en1VIgBRGpsRBINqRB
hQ+ZNVz4KOnr5xW4d3gHogYe9OxbBTXumZsGI8HkypufqBXrRAKFQ+jP5Hwol7nI
7bPs57f8QtHGmDLkera1vevScCgOXxCpnUptvj7uQqVraH9VAbgv8mueOoyDS5/i
3wO6fymHIqu3Vu0y95wamCVRnY//NxV1yBifKJ/aWHRmNTr0yo8Vjk2GAoBKkbCg
2J0idgXd8LKr1ku+fh6qwvBXe9SGi1IfcbqfT5ywVP2F+QHpWDTyOKa2pMtnKPMK
mWmvAFT8F0nFVhruyepst+h1zLtjxVwJpZGo2OHLrzJx0+3dtSI4x1ePDhM0+nI4
8oSAKjThPWaj23uO6z+d+f2MbcSZP99HHtoLF/TSjiZk/oOF/jYiI9xtQhazfcWg
KuoY+8X1FrF4uVjGiTvaDZ7J/L5wvMSkxXQodWYThm0xcUUksbbOyxaX7urzsq64
VnQvYG921JOAN3Itl+S+K6cKBkdY5laI/sGZFxJ8r1XENEJNTXjvzB1WAR4eWzvM
CPy+8bBLXs6bvnbr0r7BRWmC9RgQGUkR/79CYD8Rja9oL9ITKda20kqHFk06gDmj
2BEUMDXJojFhmKLmE3hDtspjiqxAQ8eSsaetCbytSCA4nt1v4YNmPDDWMrKWCYnp
1KWkFKkCJ23nNMIwct+pxCqm2pH4+1219z98FanoFh+ngITrdz8rS7ZnfnayN8LX
v1G9vv8MiAgluP9IfWji4gzdwSgvykK14B+QqanTAdl2rQZO+qpq0/q1IhHdMYof
fZMnrcLaJEiKdHXJCG7hcliCBk61RYmL9m4e0PnE2b22pb4t5cumGROYaRNuzdov
Ew7ejO1M9gHsCJll5cP7dy5IkIz381KKJ+RhaNe9LOgVjhGhkODrKM+FNO0hN04d
ECXEzqFujleG+8CwO8N/y+ww4l2hy9s+LvJcDPo1B00MCp3tpyvILJxpk159rNMd
xPoQ6O1BCmLoUYqSSXSRqx5boWlNF1inUquTRk4vd9xdpt8JryomJc0BdQIyZIZZ
lPtMH2ruc1wHieJUSYeNIHGu6GggrBoSRV69lmGKM8jluin9sLCQSaInXNXLkDv0
4gB4AGF4Whw5KjNYixrZjzuaNLsr6gpfTm719vHu0xqeQZvsKd4/2XE4ueHgXTdd
6bHgFvWXl/LfotIDeNNHC+2aEw8EcMIHLpKkKpUwQ4b+Y+qoPXwr/iKr8Cd2jfCv
z3ZdcM1dVmxBk4Eq72D7niZ+dzAPGVRNn0On75+BX6PFMaCcBiQwcGQr/4oTHMsZ
cR+NzL8YOHnr0ifrIE/Lzaw7X611Ru+teqH/z3iO6xEUBmuR4cEh+NXIHJl1ppXO
kbpWCYyq4MGi8ABKmXcN2A2WZUGocy2eB0A5mEhJN1UxK8wQsVn2riwJzBcRKO6C
EdH0QVIKUhKODnxtasOuTBWvIcUHyjj0XxNK1XPlEya7r1oBT8/hj5uOQfUKjaQm
RizprSwYtyGzLPCbcbn0HGTWqaSES5BuLR0LZEuydOUzkP6TKc1fSSqyh0/iBE7e
e7MASnYnOiZypefg+nqmZlPD38HUA4RulAMkcBvkY3B9GR7zBc6sBsUVAInNie8q
4TsmIKeQzNWxMjk7OpnnpktgnfYDRvk/JavBZAqvu699pKPETaYZ6Ol7hjt+Y5cp
89LZHv7rFfeTm24C/RoAnjwaTwVIFat4xTBCcfyn3vbgVIWJkl/nQK4gpNsU/nqv
oWM0hOoVZT22is4y0QNRYT3mU9k+2xGMMLlbYxdO5m/5p72aBCf2Qn89JUen6u9H
XQow+hxTvI7f8WniZyZWebEVq//A1AhFuS8fSyVW18/uLrs2/nk7B8mTA80kqMEX
zNE2r2YGo4U1lh0YME7WOdVTl94smJVLQ4Yg5cZzTMZjUD9b0uXKsD4uExVPF/xP
Zx5fefb28ZHHUI9fr4z41e6VGOIwsqeUbu1JjanafVj9hcUeyExmdPqE+41WKXuH
48C9hWufvmlLMm7V4NdCx38c3OJuQMDgDpzii1q//Hkh2OlxohJ+mmHfMnUUbRhS
g3L/EYZKjr0uSbRJQltNVF3yvJBjSanqlifFarO3VDHYesYNsjZ5edQ7P/a8bdri
3PD4ykNHqDKghAY4zSUoFKPmhH+JyQ+o8Nf6aHEo6XHGUjy4xQ0EdjbpMi5qW0YQ
cNn729wkOKuANsg7BLGvJ114fZw1rvun0daBNjfUa3TjRrBnZGrhG+DlzDOelU/e
gaD+DrQmjNK9NC4eXlbFmpmJvfIZ+q2GecQjAFJCiFoqgwf8JU1dsSspOcwiiWtN
JgKnups+17T+msNVDoSNHyJkG4frXukbTaNLvjiYn25RvUY9k6xassBHqdfbnYy5
BWHDAOa/VG+g2dQQT8dQXHMksTHvOCP1DsEGUIpFnml3p9qt2qMaCn2dzVSORkWG
uknn3KIYTPOcsTvFCMm0880Q//CKubsgdyVsgNhfUdHRlxCS7CdNbf+XQ+DT+gnf
Ky158xHeAXtTTwd8za0PJU/uVmydR8WFBTzjVFLDWeAa+fLbsK0UAJizAJw+qcpc
6sD/ukibgSH+FYgND0QUew0CKxtt5vUxpvpwKzYLMOqGCwuKvde6kh983nbTiHOs
VRVhcFP8knZVPhvC1xPhfCw7Y/ylAZVCadTHStWKseLbj7eKQ2H9h43+YMUHM7NX
+kyWXpUqgU6qKgGR3uVms4DhwN9XWpq9cxxOMxImrQlbz8aMkG4/xtPhpbU7W+4s
JurDYhWy/olj3qXoKsHwwpnI5XNigSlbqDd6PL0tzeZJUS2yIToUSO5ErTXigG5G
vaulE1LUVa3eB53YDM3EiXNSJq7PbORUIz1i5ayyqlw6iTSiq6LF7L4R+vnHea8x
KBMFXUjT+MmQad37OUapZbvZKA9ySN3999RHsJWX9gxlfe6pfL1eD3OXHJYTkDYl
D3EVy982rKaf3xVUw48mBWPk8+lU6LCqWhxrvnpwHkMYwc8yJZ39NiiTV69gTb/J
pf8eKTGefPU8p/JzjtRmPdf6Zm56LUM6oQEM9aCuyVGC1SI7D9OK1TwwkCcZBipm
+e9u4DfZaO2ORvj+1aVbHP7vUp4U0J6BW9JICcUyhxJMoBVfePcIUo8s4RoyZbaT
OT0CZJKs1qrlLd+bHOnZf/WHg7KkVH3QwGrOWTkMXAqr+Ig1gAY7AfF8rK930/Bm
1uduqtkkHkay/EbMRKNGaEJH3CTuAUDe0ZIGlDsT4DO5k2sOF8tLKamSEJmCTx1X
apauvArYz4dvIP0acoEoOtYKkykhI/XuLFLXMOHrC4LTkGO9AMMBfvFEHvnwwTIS
iy4dKVJyycdMSO1aZ+CLQT6vdGm/19UOEzQ6aNYz+Tloi5zKF4EyLx6EqlfMWTbt
unQI0OgbQcKJncaAS3kfKe4BXulHl2GC9ce3e03ERWPqDLOYF+OygG2cTWZwJNkC
o5OpPwolLf/LjYVlZKRCvivpTotvxTOO6cukdHN27iWz4u5/HjTZDVePinEPNFpb
5qjRTiPTlYMMdJxqmyGTHRNwG1wf8N9++4U6z5d4bvFlk2jr7DkYvYWk+gPIQkwH
UzHEEDSRVBEbkzT1waMpXarY3Zw2By/JSjBJPBFWQYwl9ptsoAKQhDSMMtF6nBlE
Qz9tjiUeT4lNmBFEBE/8nNZij9gZuHNt8XR3CUG5z+6wYsuh6OQyseBufah3bBOy
KMfAsFrrTOpIMBlNYCYSoAthFmfZHef2KWrykk6uFiBFzEMemQiDx2UDacPSpgtm
ETMRQB+S+hdquf1xwyA9MzBgtTusNy9Z7PqER97EPso0AWiIK4KZihYwn0MhvHPq
w/10MGMI8hwkHINrQ52LmY0hNRM15jYOIj8b9p6tSYzb4Z+FkwDDZyXKmX+4y6Xa
WBwOgJedcgQ+w25EjIP8EzSG3KIA5zfTimSi4sZIalq/f9Bdv9f4Yz3P5QNtsL9T
oTgE67i4xnZkVnvRKRecwC4OQ4QTcJXz/SxgikPahnFU8wBZnX2Bqr7K4LOcfPiC
3ttRzSM5gqLajzpvFS8PThZOc1l0+/DfFfIGcuOBgj6h78BefR6ao/J9peV9Ussn
B6cMDcYglhwimFxl0HtJA6xnZE7y8GmunhqvKbqyFjI7MtrXGI7DDspF35DZb2iu
m+vmGTOBHyXRczPArU7IkoR8ZtQazwpD83V7359mLd9Ai0CvsRyZW5F/JP6L+Tq1
U97Lho1Yy7CIJLa3zaalN8jRAf/ao+5zLyRNQzlBom30c4RdV3w0vI2BT4ffPH4B
Di437+38NrfK/+YcZ/KXUjC/JGbL+g4nxxz6LTkAgaOwUOX+xPzpeWCvyFkfnD90
ybR2pUHBEcqnKXH9ealgG4kejngW6WqMvqZuVNaFxc3fMAqOBReQdDBmgTm8rO5p
CXkFGfpQc57pdOCs3y859kzFIp9tFd1WkYEn560+Jzib3+mhHQJnmdoGD8ljo+kc
uqwXcUDyHE0JOJBwcDl2Fsh8sJEefczIoYcRzzcPPMrEMJiLKgCJ0vFwMbhG1/pI
ou3M5OnGhO9FqcNs0uVnD9ZGOqY0JJdT5xkraSjvzrr7eCR0cOliweFgCIBKz1hF
mEpJ4ZYM2ZUzNdZUOxHR+nV3DFs6tJRwoIN3mQVUVGEqLl1lsuLGvESOa4TQU+rl
cQB/fZHAr5PmF9KVKnqv6MqVF4EmqGWCuji0MBZ6gSOd/+OcWtZLXm7zPd6JC1Vb
7nJ+dDXz8bz0YUBQisFTrSLbWmjh63UqQQ5+FS/QaCPFVp2ImEuXZ6lbBobKKub0
+ES6z3RlP00U8y7Pyg75LoKoZieRUbPFxdMNnqJ3OBQ/XnIJEbsHsJmu2advoWjb
p7+R/FvdRnwMm9DldZx3jebzKv5rdIOTl+IlN1uzHpej+q6K2Dlnc4SpY6sfCUzc
pLVs3jNsg112CbwUJL3CdaKfsHzjL9GIl1Ymo4pDGTj4So3xK3H0zFPZJqoOg50D
7tJ5ZdRZCkTUNogXzfh8lMAtakdOeKx7j+Ou+VF6pi1sldbmRpfCODueJOVtbhu+
x0qaKBCDtHYokdaKjVi3TGeuA4WznrwoHbpB0EWmTnzTcDUB9aw8iDoRYpfTAFf+
wwcSWw44CHY+KUrPHuuaI3wHNGfS0GtpAYXjDZ9XJVDzAdShCEtFkNrt0JHUhKgW
+sc4aZZW06euAdAl2pXLEkfBeMAocryEJBslFiYrGNfvof/peLC6LvWYbDETDbJN
Vkmxnd+u7JjZD1FJNHzBOxqxTI8oCEKbG4mVSXQNRtrnBAZtn2GVfWJ+9a3qmfrb
mtv50Tk9OMJpZNZFg8af789I4Sbv7tja5G7BeG+LFuYzP0ypSnibbiy0W2wviJOP
K49AyuxNQjUsCbmT7JcI3q6eYKRRt34Ga3miq6jNYyRPp4H/aRh2dstmn8mXLnwt
mNDIpvlnQvw9CwWwLir0CNUdZqN7D91y7VS5EfSu2Urw/KF/Oc28LHETKUtwMrBq
wuw1apmb71IfKvRM/3bxCHDwe/ridQrprJdeyhX2nmtWVafAc9o+VlSQ2rHcPMrq
rDAUybbMOXSx370lGC1ZWsQ9q6uqa6GHEX2H9afpzF14wduuOM6aDkpJouQkXZ6v
yD9lH5qADk+zbkdRREiJWScMS5a7rYEzzza5eHTA1p13xb5FOA22br7x3fI26rCr
/Icq1O01CUqcVGwQ0DTtr0m9k+MSbnR68WpbVKRBVgeTKisjjQjnP2IdcVK8i8zV
qd8uL74oMl4/7Kq7V1ORh6CWDRo4aIWIBPeyWile7C/7qnwvafnaakiUvhlcV/9R
ujobMomrmyonMJGNLrFiXvUp519JMF++BJSVTA+Z5PkY9dY8/RNZghCm3gUdDerz
4oJFpDJRkGNURGTVmbpByAzQzOBZ+yATDbBqUrOQIH/1l9fmar/jDSUr05wtJ0BG
NgPsxvDbmLN2+jXIwMrHYRC/VMlDCDo1T3Pmh3QNRSERp2nGgZwqbqlXjMjFq8Yx
FI8YdIgsWf9/ofB9TSVGXxxpONPVWxZQB5VbrIxbC5p5rHMUNp1EeLynP4MV5Unq
imRKPbkYJ3oWK27AGihdFJvPXgazfNMI0B9zFxIZMl2O+uK2WuK0USTb56IoyNkk
MDgcgEqM09sbzy7mw7E3YBSqyPjdOP8ReyMCTuq/DS84Q+cbUbwUMrU8nrxboObg
CHfHijqRfXq1B3Z8duSWTMGRR8834Xig1EA60sr0t/mqwoeTVsVjfnmAgfp5WF1W
4bFY9LXQx6vudjJp+bz+NyBYlk11n6q5/ME07F5guznK5m0R4AVqkHo2Y3CK1OE5
0+OVn9I3yYvDL/4pFeMbkMJ0VxW3oTKzrxO5VV04xBis09dvabCGCZm70yz5u3s3
ZyhrjJjqrQVHozHYS2EmtKIlWVW0U5XLMF5XV9Dp+r4XFzqJCheMQUgRA5TlVvSI
UansTiG9wZBfnU4s4gZgOgfKI7kpa3M5t9ZazeSXZUwSK1DkqTEiMArvwl6M783s
+eywj/u+B/+J2ErwYUW0WM7HvZ5NDokOiop4iAqjwRL3oa4k19YRkVXrQdpiBXaE
HEPZe3BzA+XsQpY7H4Jrw5/3y89IbonBtbZ5BP6yxRpY41Sla5kNKxcdDhHSvwAo
acHClPPqi2yrOQj9KMTATxGe6LG3ECB3kJE9Bn/uGUG9Pf1EJZ27/sElbekgP/Bi
4szdnb6OmP8+AsAcFqxHR6EtSsCg8Z5blIec+oKz5LXM0HlElxlQTsxgt3KS92ST
XmZPI1kXCOjcMqMJpncSgP/zId74Md8ToMt0d0COUpM9vCb2JPX9rBEhRuu/KOQb
sJIWvt6N7URnPgnzyQaWBDLegTDgSKf/m3yQU4E2BPbLg7xc3bbj0qtvxddEfGk3
y7bDD0mfpqVs4DOIlI1yNvfBclhS1n8cQP45mkoancE6YFkUqkcVvsEx6zFyNdJa
Zcmzim5TiSAfMUFB/dOhz30RsoUPcks6abw2cX6NSFVc7aybgHjZBdo+xSxkUEMJ
rUhqQZrW4afFs+Ji2U7TF78ykSIeErlKp+yasiatDGrIu2+Edc3XpDKAOZsJCq8E
cHeyqdUs4Ql11k0FyLscZuBBHnPz2mhpWa9PkSp5j4jY49JR4lwrA10hDztVrPFf
YmLbE6jp7CT2GFqui4PlMtKKteJ3qlmE3RH7eiJZHZyigiKw7xAJg2a/iU0Q5VYD
mSglQvklQ2hjjo5Fnp03jX7B9c5NqNFTqWQZpCGOBYvt8pww33inX1T0yz6fa0oo
VdrE47Tpgd/lEl0E6txZ8+SJCpbbaG8JmCYDKWBHxM6mhZVe2l7tlg6YJeEKkLZF
HJzidf0w/YUxgpAadQbSoR+f53+4ceoZs3Eg0P1Ju1DN8pco8ANmCpuEZmRTDnuW
lKEydGd1GJlLpOMntjxYhDcPUXLrIxbQnGm8W1KdG0OQTlhhv7IAioNOK7/eoDSb
OuTBsc88AMwbAvL5OLWLH84FCJuK4WWfncLSjZmxoR+dnllXi1eNaBpCC4UQbe3/
4RXpOZa2iV+rqq0ShFf6vEhyAy8rVj3x6GNkIONB1AO9CyVNwYCrD19qZMpwEBZw
L4yfdm1XUsZqk3FsSoIZ7Xmyp1EAycAkJDUMx+1C0Uh+d1ZVfqLfn3TVwx9V70VR
SPXWxt+aW1w/5A623c7pCfktQ/FpCsf14wWH1wHtHUXmAwwz8vHAWLo8U07CmIN8
WPLZ2ZQxLzNYIMcsMKFMAlDD9SZVeDl1FTOn75k80x7jAiYjXUUB1zq0ZtlwBohy
bKsOSJeHRRnwm3Vq9mXqPRJaOwhumCWg6/bjtde9htfCuTe6J9a7iAcvMSH2z2+s
xYnuMCAdxNP7f3hA6fTuIqGSld+Nj7PRT+MKfrDaMO4gvszakk5gq5hyLuaojbvq
x47PCDzREw9ZbT9Vjs2HqNv4JI1Buu88Hf5P9JhfwLjg+HCfj9+pSZsZlj5qC5Ba
6g8Qfl/6D01ZW9EEVBdr4pCAlTaQ74JB4uIhEAw3TlJSUx8jVRbqBaE1cFrJOwqj
Ebv9SXjAGFgeal7+dO8jNvx0/Gkl1cMxMRO9IdGMSgPUR7NkEsKCBKheDjMeUNQ0
lFsrN3tXzWMcZ1u3vhLpGn/fmmrwripA+/PDy2iSpQ4CzalPir/X7z7MVdzfA5tE
A0Kg7uHJZBFicqFSht3yvgHQhl4jbT0M4/lFqMQT+JdRjOGjAbKljZRXKc7LNDs/
fg8/79m64lLzAVoRIbMRuKSRp/Dm/fqjx2xB853wkquvu5P/hwfnFEGeAIqv6+HJ
WSdu3smY9oiRZROpnLPtZztP1EnLB3gPpq50nc1bVJadh37BzYecunIF5hRcxp7+
5FWwXCXqX7e/3Vn+taz026Y6nPjnHXzfnBFWF52jwbL5thvuuLnsvmE8LRPO3RHE
kxc1E3XFt6QZCssOgvmwPacxi61OB66Qa2u+vtUTErW0CXUk2ZuQJyvvPOYvNvOl
zMrU0GchsnU4YCzNn8IANm4pTccV/fwDxgQLPzkzMx0IFjFGJ2eP+TRMtZ1As8QV
Cvjju6Xo2QKr54k9iqZl10tbe18QGu9zOvLiKi2CVulDwjQnp9XVkXYAs/caAz6A
v+shSNGAXpO3/wqW5sEFtB7qxeYfzSDhnq1H2grxzkdgMedfQxpUuJGlEsU2NCu4
SGPuO41BXB4YvHgE8mxB+mxvuJbASbHZAkEBLaVFcwf2cRvTw6cO//Cn651G/b+z
L+vV1vCk+BFxcxXIWvMPQUd/0Eoxgoy3FsTBiwzXJ1T3oiDH7a10mCWOb7K+Lp4M
s4UsfQexjBPIPR0llJXEaUg3oEhRwVPx6UyqWF3YApLlygM1/32/jfhRlr6C0YJR
KkSsR3rM0X1TUKQpKfrvjPpg+YczYDVUYSO7oEAeXf641rQQeaOxdfp/eWk6Jd7Y
E2LY1WSFO8GXjr+S4l39qwdheOHOoKn7cKt8v0m66UMLr9m3WepzGqlL1hX0V9i8
E78769qb38DUYR6XLILwQg8sjsH0mHouY87DHSSqXzTJLVKHfwjwZHp9Z559JDjC
VLjqJqk5p3Hrvq/BCLIW0w7na6DPGyZCdJlVN5huSLvjy2qPA/wd7qpco1V/BMVI
8b5HLg6C4XOMjsnSHFW9FP9LJFZXgPkOo1whmS+tgf5gsuoWVqykYER0bzFXQ4gK
w/tdIHJAb4EYeheiSrWRT4SzJl9DF+38WFHkZPabe/+mCJfySX9buai/v9Yt1MoQ
Bx1V6WtkEx9UcHMfw4G5XfNX+8wD9lJqr2VY40rDNYjLjsVala0LeuTsMgUSd5OI
zPakuSlqlHRD6Vn2EGfy29SKuesF5QxZxdZgJ0H2vcNCT/e72mrRTMsIjPyXnGnQ
nSi0ivxK9kPwtbSYGcusGLDLv57MvDQ3uiWF56iR5clY0CrSHiE+Lc/QdB1Q8Dpy
cO07gzH5a0xRCTjEsLy9/Ssos2mU1XmGleLakgPS02QKDGqtXoiwgNuxeucYZC/9
/mcqnGXa7y2XvZfSM2NLBLgye92svxFxa0NbT9TUvj6cjHe0pk5bDpD057qyVsbi
vSNZfg2flI/YxLjkehRYbJ0hpLs+D2I0lb9e4tGSjoOFfhiiqyLTvFZ5+vfCeNFS
oHLdGMojTgdXz5MtAVMpHVniU4TW/OPdpuCSmcdFXVX5b+qCnVEFO9DTmbk7fcZb
VWW2sQKMGpWOFX533YLGFLoEjlbM9yv3BbTEyUvaVPMpSLhd8bqr7i4Ey7COANpo
jUMYfv7a4M1KROprYp9GV9iltYCzAyASXvVPTpn8fk23zU2iBVg9PKlAU/xqZHgQ
QKjNesEqnfxDbljSqQMXr8pvmvM598ChePkBaBInfhiOcpHbIzlRUGHLk+q7rHEp
7oWrQpzgvODfX0Ao7EPP/TzYXZ3JiC+Ftf/BaVu6TGSbXZISj9ZPK+D5pgXvL8N7
o9E8iCar1Az6TGOPwX2jjscGoZO3FuUhujxInkpj1KOkeT9pTmerGIrloC5+ivc6
fbicKL79cmWVHEyhGQx1nnulHKXwhBwSOnsesS6TwtaiurLELvTP++qID5irIoEv
dTnKlLZFv85QpEkCOHNsDAkkfUis9fOXCPs7IaFEEVZcNDgaB/Rpe1/qiMwSMfa8
jX3BOUOe1vlRfCf57KFpHU71S6jdgAxdRWgwguyuMFdFQ9A8HYzCR5tbR0HrcmQX
30tXCrCFmW/zJDT7R/RC5ss+M6ACp1zaxf7RP9spUTj+CYOVCGcFhXN+ci6Zg7br
uVUYkZV38+cWiamJlnfmeIGNxV7XD12QlsPbSRhkjA7BSS44v3MHk0GI3YdUGOOf
MXY+DNt8C+ZjWRYTHzYcwiLgknVKK+o1Bj4tirAGebx7v+3nuCCacB2sPtKljrWc
A6H2lBvQ6JDbeRXtue9wb0ei55kZPo2cCrHJ98CTvK0ztU4yozOj3aJH7f7TFYAM
F9fJVaBX5x1cKqY1iJUlXMhqqurGnND878WSW2xU17tO62KoNYdw0pMMfxPHDppe
Y7S32HwVxVysmj10r+4Q8ydXSHmBbV9csfTyHWGd3J7REMhKi6VizxcvOZu8wTWX
vbz46glPdZv4/ZTpJC+D0YI4CtGupYcEguyS8Q5eHNsYJbAB330lbzjJDuuGS2UR
mglpqltwnYaxdg0udjdbs1gRRnFamOx9fOGWpbmeurR+xG3VpnZT7dHhgBRDr45I
jQLm89zEl+cVwqP0vncdz0MpSG3e3nLoxg+XLUzW+lDVL+w5G/HCtWp4+eUilr6a
jgWLwEHc2/37pZIhCTJDzmjHoHFapTYX6YkhKQ2jzzcU5zL01yxqZJi/F5Q7IyL5
aRRhBwRiE1w1bXEHQbq4IQgxQIYYhCkmkGgUt13eUE62z4ihvN6RSlwk/uKP0+V1
14SsWydmbS/7VgIbCUqlb42DMgI/DTEyBVGzMf9VC3zQ8SC3MPFJkomu3+ElKYiJ
owWxkKlAU3XMkgEsw56zqSKoo3mAV5zx8XRW+uZWOQgH1bQPXb0SU9nOxuv87a8a
gb+tuOWcS3yLehGBqqtzyHYz6T/O11KCMDDz92sLV+Ry5LnNuBroYKJ9pPqpHs4W
wyFv2DC6PUTCi4S7bVQ1+L8ft8+qpDh2ZZ7mZKvJhHYoeyIzt25qPAMc4j9wNS3u
18ytInRj2N/h97Tv3P+nTWHQ6/RTJDNQrLULsYjipjRnlB91PL8TSOiVLDYUFJYp
hf+mYyABXU6I6sj/kNONv6OX7l76HgZO1en2TQz+PnKxmt/x9pePNaQ/AT02LAnM
C1kZKzPbbTS9XTle9Z0nEP1pl+icKwYwnfMolRIP9AYgE/WC9luK8ChM782mQ7rh
pJOah6KTgJbo6BEM+IvZLjz157yQ0h6xPKn4HuWiqlvf8MRd3UwdVlcscxPaVxCo
YgWfUk67gfOT7ERBeLYL0k69RmhYD8+7/3glaxH9Y6tcsqso98Ges7fDhZhoTDbP
1NHUgzPW73S4w52bD92+emBZic0n07pPW4dC/Cj6aC6uaSUwDOOyE8nUhGU0Jiwx
yufK6dBdAo6Bz5n1Gn6/6RLUEINGGcYLO+WaPq0fd047vbkyqFYSq+ZEWjaNt+Q8
PJ0uGOo+/iwAdcFaEJC6Ac9kTU2FAxPIjOf80r78weFx+e1v6SitDfWSXqsVH6T2
yyc5KaQkpAEIqdjbh/U/YTXl4hh4AYTRx+mGVkgYzN8vRdOAe4ulx1vhdGuxDTte
wtmfhACeYzYIyc8HeJn6rTo7KbCEMJxQXsAzR8aO/BE9fvPLkihryhWqBfc/oF9b
eXvAeGHI6kskgsCvtKlnxrRkIupQBj3OsSL1COB67RKb2Io+rXvfCGvVNxV7nCn+
1jhzwHDA21xvdZCWUr9PRqn8vrkCLwBDPreow2/5be5lBn9aDW6BS/yuBJTMTgUQ
07ufgZ2t9dgrB5huPQX72h6aJeZZLpH2xRAtk6n8zwMpzTv4T8Q6mqa3B5w46IY2
kKHWhRWGoRot2MH6Jgw+0x+VPfpzZvXKXjwW1HlZEBaH8JtKZ9zxfYEZxMDOzL2V
mAvmSAt0s7UtPETBQEvDgB7x8NZYEM9sMAb5+Shcfc1A46UOEUiUgOlCvgEd3GyO
q0cxtkvqGwKl/nFbHJMbdJKK08mWSQZSJ4iefT6nP+c7u+zuw2zXS3vBIdsRO9ge
a2rmX4riFt5RToHWy1SCcIKfrou/jppeWr182vxW690wb1j0BGUbFcT57UrO0s8T
DTsDIgAKiGWtAGiijYWTIhDvEal4wjgp9luFll2BqS4EDFL7Vrnqj+mSy3bryfUv
S60ug7Et7VM5pQl0nF8Nz6YEaJ4odGDdRu/7M5N1NH67nfirZVuwPtIdS8CpRBpL
IoW7ZO5Gc2wTLgU4OX9crSNPOU7lAopPf8RsjP7IfoAIq0QKjFRRrTWoh5pGTT8j
LHtVijsw6xoRUC2nDt7hlBStDP5W+fpJm4r53cUVeEN5OgPcBtbz7zUwjP38xwbM
jgm16bjAs7KRgIcZepTZzCV7oe1bDppjzwBGClCKpInf8AwPa3Fd7g0YIrUPj1Nc
BTf12A57qAyDWiXuV4QcqyIqiPCEHisOXxrl60SyUX0jAlEzTw9QWxZbtvX3G6iD
UvazD/3G3UTPx5cgXYme9IB+6z/sIAQs+AoJsdrfn1Bt3d+Ju9W6IL4lnTv5C7v3
KqcZHdGjANvkDU870m64JS6/2LLZCJu4iReadVDnLjA9ds5YLwUDbYHrMIufFDLS
PxgC+wimBLaYI7k1e8SA7d/gJYAg2VMhXwSlLfxnwyMNLE45qkwoWF9rkkScGxb2
k7XozvUQOWpTrPmRmP/hpxHTonbBK3l9z4rJVKib+97rT1/xc2Y0549EzOgMk5vr
ZzgrjusxlOKfgwfr3eI5PNaRQ4DyRGv6TosUJA/7iUT4PGx+1F+htBqbUeDWyr9l
wwvXBO/B0EDFy031ZfpJJyaYi5TUxRtznkCe7aoGB3qfGHhhbTzE46bGTh/Ph+x6
YFHPd1yijvfFCLxdq/C+A1nbhKIysumzt5ADjceIrBcaXZzXibjJLQSy1/wd/IOF
ndNUmTL9mYZ2f9mbmRwwBHoD64v/+wHePtqotRlF7OKnxrc36y3lC+2EGLyblr1S
Ao2bwwh9KVYDEXwFSv7Ymg//X2pStvdFyIbnyQkh7ms4osuRo3u8gitXxZaUwjEw
0tFv0C+laRKvAMERLIy5wCT27pTblFG5SMVkvHp9r/a8Tq3Vp6Q/0JblQPgpEuFK
TmuPrPnBfqMlwurkr214GYTTo8mPYPh2nHyds8vHpSVQB4PUArOrFbNYdXzQIFH7
JVecm2ijdLd2Aw/lBiQMajDiI2mJuw+YYD7LIxwQD4ED0TQGZlWu/QvWbW6levLg
ohwIdy9Ch/cdJELO6/n65YUfHWz1OGqAXMfZc6mLhn/QTbljdRTTAhWLGWQ7RDXm
FhIGgUjJM0LAa1uhyjakrBcyGZQBACgO1Y523uzTJeNgOeFwnWcI5eCwzp9r94gG
I6LY9t5sJHuIc2QAFkWDriEhnGJYZKcu5k59eyKNjUX21dwV8x/0jpdgjOd1l6B7
lt95TDn+sbJ+p60BpVJCf3lp/HxauHOsw91f8a9tiAGe7GBjJcEK93mbbr4b857b
WiAfBa3hhJyqb+0aiqPr02KswTvLCpEYG0L+jehO4Q76ajLFSJBPXYA7/AhX/z2P
ZvVUxBFMaH7/30txiBYfIUeLNiOHOfoYEGnlTy+Lw9V9dTSRnR6J1hfAvVHRmi2T
aZxlo0kuURcxgaLx0YueuUUfF1bDIC2Jj9XZEmUyvC/J0BJdqNGjzp4P+lUW8Z3d
gHpbYBH5nJAMIiG/eAkw4yJHB7wYvOYfFJlgkKbdqixvPS8Yj4xYliZpLqmt632M
iPHQGCwbxVkgfKJaK8KfCChZIztJoWlXGTJSrJH9UXZySJ5eU0NojN6cskBeBHA9
PEDyAOS1TlsjoQJpRutnTVSvwO6nQ5jOESZ3oC+BeeatDdABCnZF0mZVCA9jZbbT
hLV4j62MCb/0pgdjwMvXJyyKmDQnCcVQuL2BWRnxtcyGFnRVjSyWz9WxCNkpR7jB
8Nv1VHGB/saEJC9a0SkvF2DZZBcsfD0S9c1FiI65PBN34SQ0ESITsBYm1aaUAZXz
Amgmv/o8EI8rCSczG3iyzO80Ex080FtP3+/SKeou+mn8LXKSP5cDjosvz8/trs+P
nL4lqHBVw5GKxWCuTMBQGFY4RQEgKGtJdpJ6GcuBCDtke6uqYtTXKOkgHX76sq0D
ioQa/0IMe7jowS1uI/tcu1RvxkYki9MZiyIN1GWUBO8X43wAwYGoWoH4EdxD2fP0
ZzFMVoxNwYaf4enJcYcpNbUcaOkAee16hHhNsH3OUAIN1uAr9pHbLEoAJtVsCJBh
UZR3n725/oAk6sFuJORNuwEUqnekRlNUNWi4x8AVGXgwl8MVYHKzK/SIfhRDGwPM
2P3DXJocY9lanXweEBVNdxbhKcRHcXSCmydWuTVoj+F2kcHnirrc4+66oH9R0pZK
3H00blIp7/Fno6BpHDfmNWiNQspvatqRiKKnsoY2GxXJTN4swq/Y6vJ45ezCNmcS
zC/XU2GBMdbFZhKCqNEWwdvqdn1Gj2Z9YUJq7ondiwuC4I2WskgwVXQsz/Iic6tt
anY5DUtCvlNFypfweML1khEyvVVDQm5+Mzo9TjvhHRoMt/omhCBPbfRGGmU0dwli
5XKTSueeF+VQMOQ2SpwRsnke7uYt0skvu/Ck7x6sKR5JWTDtWZmfvy4SucU4bo6h
9Lzs27ffysJgzesqWN+24bZB3fM1DL9DI1jOR644fjM8xtiVQqE+6ULTooiycZtS
ylUU/mGap4zgipFwzYsib7KgivKNY5pQEGiYVG5KFh9lTa40/tCy9XytaIi5/r+S
i7IOOgLcyWDQxltwDsquZzUzARHSpYi2toCr5UlYdmG0y0eMGIzQmxfMV4DkTzKG
GGf/KNv9umFjTdcViQ1nizaJlFHsZh5Q6tUi/PthxhtP+aLcQkSnDV1ZhojetdqA
z8GE99hpxgXPBG+Q0BRTgql5ASshxywI/fU6IIZYJB9HP72kun3IojMhCT2qskNy
5z9lMYXCmANcYZlc39h46kLgTKrOWQEN3JofhF/yifu5bvSjNBo6C5rMqpbTSo7v
1kkzuzBgApJB0YyB0B8kxgtY1uU3feFhFt6Y81KABOJaEaw5rHSmy3hEcm4LG/h+
Vun7fyvbepi7iCUbjD7wC2jfgXMBd8CxMCPGAcvS8ZdL79XDCVaKKXHcw/zFDIFj
Qf6yncFT0lDVxhmlM0vcLsPoDo6AZNnKWmPPfaxddDKc+g5A42yl/xajnKz4A8OF
Vm/PfqSOJNDRIROYZR/hNCqGrT0st3SrneBuSFE/q6ev8lUcj5AItW5jDTH6BRxp
Qn4Cesv3UnLb28odYiloxb/ZJouG6r3Z51oOIAa8GlnitVBbNrjPW4RrKoIc7yG+
RYNL7ocgmaG94VH1iLmZYhLOJXVvCsl+0Kxmk2ZhW4fJKL9YhyFud5TBHnzW8cz6
G1KEPx/2oCA+rJMJSzo+kfNURvkJGsIEq5BaWaC9i2XdjriXLU5S3M+97kNseNJV
i242I+ir2KvYqXLPjgNXSszsP6Tv0QyYqQYSlQxDoJqcJFTKrilhfrY047+M6060
D9ZXr4+431z9Te+lC/ltl7DMJRhIeLaKbjrs6PubVyfSiovHOrQiYD98OdRoEKWz
ymXFX/B8W1HcrPJmWG4jBCQVrlJR5/HoGvK8SCu1dVs1BQvL86dNSdXqlbeoutL2
stvxBmX1fmK8/J+iTldtaA4ZXMgHyjkjmu6/BmEEraiyuHtC3LWLg+Dk2BF3qlOP
dh0V5Pu0J+RV9XLvJxvZLbvHgrQqYdQ+1nEMgoGSlnwxfKPwuYeOuL+Sa5qMJZso
I/TRivQhcDy2MrR04nePT7QEUZE8eruocoaeSDC0Qfa6K/qjAVA5jA+kjT8njfh0
s7wSfZ2Rj0FcZYtsPsV25h2KSosMVaTViVLRxIQNuHYYwDhGwdEltuTRMSaqbCJq
m9bYnwftWSd6WLzR7YGMQuRzV2wpUgo5cVkENGCpQo1UtSJpAOfYjNznU/GlOmNZ
oH8D+o/kvQOyyWdn5xECGrAJe1DXslhnEDxiTZggjv0j9QKeeHV32yhSPH6slFt7
1l1PPIKIyF5/A2kQepcW74DlbURB81oDxazivDXTOesQe1fHZtEMWta1BOcw1qNh
H7SSdGF3rR2dYglyAZWy6Ca80z2Sx3bptX5cmOCf2NaOwHh6bk1vVup6re9u3/ZF
kyaJETqayJ6nLAi9SnjHRsKbpwcgJADAc0h1/Adf+Eg53jHnudNoGLA92orVKuID
VOaf23sOwFkH0rt+9ZlSEA6P67Bl4hBpC3mG4Ow0NJvzTCk8EN7+ysVknxm2uMtP
bXcXgYGuD8o1t7aa9Y/02DjiIJGaN5pZWdHeW5XwxLg47KM5bNpZ+TKlOIJHnXsj
oTFz+SIbhWV8WgMH8qBb6F/Cnjw/3EmsE6xyaOaLyhbDMZ5nHT/UakiqbMaNZEzt
F0YJQm37+yqhKC9Wp0Pu3YIwxGpEKINwupannXI4fnsPlcc9QMroWZ7dna1L3qyK
u/NPlUAir7ZhNcfgbs4X8E47g3GdYRemxXkv8/H4VEA/HyDyX1QDlV+IpIG393w/
M9pL62DyzqWEhj3TJhFVqQQjPhz11jUeIukua2kH/pDb4V01QBbyifrouPbeQUtl
5YPWzKOg+YnqbQVN/jZUr60xNT78IB+VpRrfylKzdn1aVeSrZ4tQWFBz/rrSqFvU
/z/8PLCaDcuPje9J8CqmRl8oPT8UhNcLjcYSq0QMpx501eUv+vl4DkZJMwf0mVZD
//dRLjYVGV1muq1zWu8iwNWFYEgkiomBtfQ6RkkXknKF5T2Zb8p4kj24rnLDIu/u
8nsbdFyd0exbAMBq4MQ8D6iOrtltRXIxhVS6zu42U01ElugjucNW+mKrl4JFe4fB
2I1e1BRdK+Aq98RM3m74MeEZTQxeJem9rP9OuKHNg8GHd9plxwlD0UKul6wQoDxL
bag59JslKKy9LyU3VOHwLZ23pxvftZ+kj+13uOZG37mO/XmyrBN6Y+TORlzk2fB1
4PUIhI42c9ZcGtglYmtJncPFpi8nv78VcngfQs6ohuR2KCMYy1xSTPDwPtOHnRot
rKDew/IWxsOzZgcu+VvEm5bn7E8uyO55TOfz5rYmSFYoyCySKNBbOQmn/RY5ON9s
5Yg6dh46eZ3wmZ9zAhF5bptYVBKJb1W2bwzytC1pG3pBC4E9FdaK9TeLX1mY9/5w
/SBknh+AN/HQZu+VajQ/s9RZGm0uLUUb4RulQnPHBWE8spC1LgQyQs3NGYrMYoW+
nxQtm4gBKYkspjAFKttuvDN4bRk9o6o2vn+x7FOggLiNpG+ZuBPPNFOXb7RRR9LB
GfmtFwJYOHUt9WFxUDFdPqTrsDP+TsCjpW17mSs+/cb2/rKmyxK2hWmXEkhZa9k0
m/KMgJaFne16LUVvg5Dd+s78OnAGT9oy3I8qemBKLAw78AcqFURCuDDBLonl1Eio
4JFmphL+7NmVMcwhEzcJXAuAuevR900kXj4UqXazSANuEAzwlp6fVJULT9V+ORW/
QQNBK+j8r3H2VjeKO2wZqwe746bvScHuSL9SQ9A60oFjwJAb/XEE7C7ZWFQXU/Qp
RnRF0Tk7aiMV9NBti3r0RbbmYxAGINLh7EGOtH71iI8XQOOTNPWDtwagW4hBXn88
y2lKB+xy7W49x15Br7Z8zBXbvbxpeRKdTh1iFmI27PrDYcRooXgfMpasg8+8mCSX
tgTesJrwcprj+NCN/5Nz0avIcYTfSnaV0t7pUnl97HvHD/puolpxFUuxajj5TJzT
he+6CUQPyBG4kzOsdAnBWz/cXznLGR5xgFas6kjiQXGshI8q1wKysMv2TMkyK8yh
AcANyFZTjrDDmAiJwN2pF+lVnANX3Y+Y4xM/pza83QmGU38JjMDej8NSu9D4LxuZ
KU5Hx2/hB4Ux6qbv3CmAe5lzN0ibHyrcsR50r4Jl+GTTZ5o0i0kDpyNfFEfXh6gk
ZntTEeWHEDM7MW8h11ByeAjRLtgjWEU4hQblimtnK+hZXPqXhtvTeH+aPqe5Tcwp
ulQgxSF5Yu1fSPmpu+YClzBygM1nVWSK8nm7Yrwl5IowZYFyqeo+DK4KS67/G1aP
N/e4BfAqVbgjgoCztbBGc8SCOFST51qX95FZ3aa5kYbMKUkhlNmjsCWfm884BtQV
U0bsmWiw4hUDnnWslkwovCMPoKCizceDQzAFHHC0BsUBcYqV6ZY7nrJAhs38MSe1
EKTji9i0HL46lu4rsqL3I8xkLRaGvoOobmbenWb+FANVhlmQEAIN1HrmyjVOakyK
BL6yEPIHpqaQ0psTCli+360K3Gi8/Di0A3PPira3QJDwoiT5Qc3YYOvy+winxmXV
ArtTRv89GZa6XPSykhFNchPNzbLbzB5BbgZ66zSp7+u+mlgt05t9dS8p8qaOkn73
G4Zzh54O1sgCDOLzcON7156QWFrRfj+vaE+Pv2ZWqqQR7YBhvKtK3YmBVuwsrDLN
icDY8w+rHEyqwdWOnNwHU8x3DO0Q0SDo0NJtW1PCviOAJuLnaPwbUXZFfhYnZs2m
2i/XNd0YDp2x/Olttv+leCFlsu7lE4popihobzOTzDFs6QjLLAMLJqPcjiUb17j7
NK9+FS7eGUl/tt4OCxXbTYU6CpojHiwWYtR+dngLxwlb0lIKfI+qSZ1C5akhdRot
yPA2apHMmanH0bjz1AptI3VoYmYugx7d9FxBiahELRC6OkT/NdQ+V8t95FwrE+ig
2rUZ4dXooYryhZYxL6nD6qR56JIs90Y+KjFKMl/mbS/HgQNo9JqUTrlbVsOiAzHY
c8oW23kPEZrwKHsn5U+WjfDinTLZ5wjAxkqtwVLxDgoyVp82VmT6Qc9YsHa7cXKC
b/e3genP0OC0A6oQCOg6d4SLABznN4vR70UOIrCJLEhWCjxU4BDxSRGTHwRGpp3M
oIDz0Lz+z8aRsxrqwDm03T47a4mcBSiMMDRDHo9av6oeehva3KJ3WuvZq/5JSPSL
y6ws56lszgduNeWrzoh1VuQkcm5AGCv+DnNkvICwVEYBLoeCKyJxDwgSlS4WeOwg
PSR4TOEDiBc3PFXR/SOG9zjj6P6kqveH8S42X3Wff2c+wXgqK9sBIx94VJYtP4HW
wxWEXTt4KzywMrEmvR4sA4JsTBXV2D2zpOSTJLikaYStfNPUT6qtqM91ohDJKHIl
hEtpz84hw2fM3tegLrKSJmOxjvq+eYWHEcM8jLhRaySF5w1qFmRZzYoN4RDYB2Dh
ZpEd40HuPgC55L5VHsdjhqEw4/ZqXhomf0vY+nQ0N1j1c7MGGmJZ8be4OLT7Qpqn
STWIB4fJqssTr9zQcXoUxorrStCNNMmdEVuOTwizmr0IC8Uze0EyWwv9mcmX7XCV
TUM74WtZuexUrfH8WyZHuSNkyzGWpNrhKDnGGKLVjfB8/9Cvryb1CknU6mKNB3GZ
jB1orio7IQ0Qxy8xn4BQnFJ4A0Zyn84OQHYZ02XKx/OB+Ml4Zze8nptjPvtOxQec
IWlhBsrT2/3SkN1QdmcEu69FS1IS01dAvBOdgsre7/V6FzjDw+22H3Hy2gBQcjvW
7MMzS0+1d3fBntihPQr9ETAne35SXt52PYQVXYsPdvatntVSN08VtUrUFY8zOv/T
lEJhM7Mh507uHASzfptjHeOfniC1zIcQOYMxTNZchk6XjXmMnw0F1LOKuWaIB+Rp
fnjOpf3VVZck3bwQrM8xfriFi454KEqKFJDNIDpFSr0SIEqs1q4U07B9itWwBVeN
EHJ+pR3pR4CF01yHXHKRWFMUXYCrl4xb+k0Sasw4aGma7VVZwLxAhHQ4Kjy5CH5s
CcTG+l67XeG2fRRFMeYA6nPCUWky2PSljgbyluEDwMyL7BAuqRvE/1WkJOH17fJX
lPySrZ33XWcRUKQteChHNahzzPa8iA+O94FwPMkauIO6hmqajtkk5S9i1AfZZwU/
OAKfCTPBqXq0FAgwce0RH8nIzbovH7XZU/B5QliAHLMK+NsdVVBh/wxSOdkZoqLF
21wKvNNFhvNLILRMnaYQvwu/xsUWc6zBKAAUyh7SUVtb5QIwodnL+1MpESYz0Y4s
h4rx1i71K6yLR0CdiAPViY/bKkCdAIlE2hLT0sNqwA58V6haFrppJmivxpHRl8Yn
wZmg1drsqUIVc/cq061ke3Ye4CxZg7JFtGnBDS98wr5TtRbpdDmSCh/RPXhkgUs8
hJTmwr0JK0Myb0MTfWk/F9b4vqyNsHRibxn6dmSulvEWHetC5R0BuJHaiuGDpI7Y
MUHVjMyBiuunIMYjVryaV1PWxBhWp938UTzkKX8wS2qzO2/elvGYTL8DlZHfXMzj
txohwt1lIJcZbNkpmN3JsXZHRbEI/ANbXtTdeQvu6exAhP/GakHiDpIDYXmPczTb
qhyBzeCCcUVQKN5FOHe/4HpdVfFJTfmUeC03YwrctTC5EWxC3/uCBg5m7ace6fCV
r1i4xCFuXLLCtim701+rrPyzMqmQm+fSbr2Fz6GI4RT6wK0kRYrRiiS87dAxrA6j
aGgeyzn1ogAna2Ltzwx6fFW8IXPjWUL4KzQGqsTzyreZKfrpx9r3n9pGK0tKDp62
iSoGL0yrdwqYHLAGNPCpxCUp8vnODfKMmxYc0jteJ/Avy9iRFaHM0ZUaLMzBtyDe
V5QjKte32w8B4D1eTLfEyAXCng59CoHOOOvjoeFbZBERUkNTOe9hkcBsYwLyesNW
fDDTm1wtofTQckgVDWl9yNXmkXZJtCI8SBsAo/dlNTEuWeuu+anEpUFQjL/km1v1
UrwTouU0iXf+8US2TYaSBGm2G3lwmbO95Qr2e7AfFkqM1asjJXAK5hWpneE1CZ81
RlEAD9XmDEe8QFvLqZtCZLuHFIji29psykh61QAuJkgqp/W3gNtfHir67xHY1nfi
d3ii7dVROjJEmeKRYoBNXoLaM81J4HxpXPz5lRhyw0ZE9vGDJBVc01URRRI8O4vW
DWKXJX4C9n6YxbWc+mmg4GOIi7tDAH8Mx22dZO+ier1IRV/zG5aonnQGPV2qeqth
uusJlQMv2PMoo9QcqNaLlh/yFJfnA6UyU0FnmU9dLsfmXL1eRqg+Hjydts5e/EHR
7o1aG7TmwekZJ03R7WqhshYNKPFQT/hqUvjFshNotzDI8mHo7YU9y6IklWH+U0i5
cnpks9pL4/emSDBvoWywoLKvz357WTelq9udbAp2+HDBQ/Y1po1+z+unTYMqjwdf
1NrxPi9pd2F+r4dXZt36QlNgp9+Dg74MSXz8Nncwc5JrH1ACS+cnQOUmymIoYwaZ
BII0RFNqiTRJwexU4hMk5QKRUN34XasHWLkRCYAYewdEgEK3mRaajcn0kZtX6zBw
swlHaF/uFkB5bLRfPg9ai/RYoEb5Xr0qvkBljjtxCfHi+9CcNiXMcBiBMLS6I7yX
3FZKhkmVX/gait1DhUkm+LezkZYJsZd+eUiwyif5oKVpaQfd8IMiYnNS4wMDfdmn
Nt2wgRZD0Y5YKxmAtxbJPaaRdMwOuxw4Bbyd83MG96op8WkuSe+v7uyecaMSIcZL
V/5hyimAYaa11cvBhWt2nxfAtIosk+fJcbyNPL4BBQO2ou+matchODGaACZc9S4L
c61R9EASk1mgrJs9PjZR/3+adcHLRQB59z6bvG5IehAHr+yJhQeodxZVBBJy+9zi
z/6ZKjlgg3JrSSEDD9tSidZqhrDHK8/cRRNcqQx2RqpLu9+76rJ2GqMp3SIuONDP
fe64mJPjV6K4F8jKwzgihTV+y6eV392W2ZL7LmX2zzRPGZJn1xSolO2qH9hyzVV7
T/sm0wxXfa4RLp7+MLsjz0BnoKb7cr5DmLUJF5zIm2Uh1MRasNENl2nmyMGsoDxw
1S7NLglsy1qihb++eIsdMvZqBGAwL1onzhjqKYu1dgu3u9I+HQc7XjOUfq1uPcWb
gnhVuSdIRyxBH+u44HZAQuOWCoHrIlSFtHjDsM9s2IiKdfTjtSmrGopPTjYKuY08
bWlYzmkmBD+SmitNVCEKrainRtNNsC9RlNdP0HhkhZ0aq+h2v6APHYjHk7ZSTO4h
GSaU8l4NTYDnbh/kauyIey/IswkuYUbNYJDqunR1BJnzo1fqzoC5Tvkg7wOZKCkN
jWaeNTJMYFFxJZy+zEAthbuc5vJ4KbeDIXQM3G7n+Yb+1YbSf+wfw2lHNRaFV9Zg
zfkeyKwLUUiXMkjjmggbLkE8spJ1LqB5+0U2z1ETHCAX0LWarOfLzjaQ1N0i+Um8
Gbc/eo5F2M5nGAKf/Hwu6VoxJhJhVv4rYPAkSaMASMNjj0gz6vJLp51j9R57hIpw
+zaDYQFTZ6gbwTTF48ltQ+HVAa1Eq3gkNnuZVXCmV9g6Uq0omJQ2pofgCzvf8B11
F+OIRB8YrrspyP4kivh+h33ReYBn2EMPOmN08uvmivji3gc1lZjXojCeAR2ilt1A
UnOtxquJSI9WW55YS6p0n8k+3mTBd5qkprxhc/dmS5E6Sw3e/72Lejz4lG12gHQo
G8KYs9PggaEYWxCoe5T3eU5SKx/gqMrAevY4l4VOmM1pHYgmV4OB8hUk0i/DCXI4
iy/90jp8l9K7PnnPYrn2xfh2NiUUITy6/g8FUpsvKUpUuIll26fCt9lUQWyBUoB+
EqrFAyg2QILX//TsQme5vLw3pPLe0Q/EjOAdSQdmG/Q+xEFs2M2P2Jm69JPi00wq
mx4QVxhUytl69OFB3DGrevMRWIH7r8ndG1hWkHrlEcmWlEE8W6owxVtqouqFFS3j
1tMg7lWp8XX7E1nnTBLGGEIzhVdcVbLNXgp42GY3jhWOxekzrxznDJ+75w8Moi7l
lIHDMd1UnuNQ+EKX8uYFuXnSL/ZfWHDKoUD6WWubjzR8xZQYLb/yIyG8edArxk6B
JbaeZzBrJW7Mzk3t/p1jZ8BtEl4wzpPNajEi7+INAbxKXjgQqDMUYEtaV7Hm8i0+
x8ovD51iCfGXT26NHPXNFcChB5xFtSjW7GQ5SaFc60os70ID2/kjKxSU3YOJ1p3b
a2LC/V0n0EmtRXiesbCSvO9EkZPB5wrEFuCNxoP6ybPwtuGwDtiCGsOOwLIpwLIy
te/WWMwxomZBPNDAi0TmsGMsCByy3RjsW1kG+nhr+1uVtK6vNvnM5evKUDOcyWSL
g0uJsuupuaDCNB5eIjvMu4o4yXMyAKI6F6gkhP9BQ4N6RPSujg33gOY388MWWHcM
2lEMDFdvO2RIlOkNx87sCfKtYOMj1JbCs0WRzR5pOomzx/iIQc1ZKeCp7nKbpgXe
+3MSI5zwur9/LRPhMCOUGAITc94Wr3Y5+DKV7DY2Pf3mhS6VBnJHRWNDF+77ZkW7
yhT8/nT64z/0f45o2+TGiTVIy0fs0L7xjGNdO8bKvSxiw9677IW/rmy5gAzcGgYW
SpsTWQ3EWX0WRNbQSQi05G9WfMc1vj0CBmt9iQqOAu2GQlBCkGd9N4mfRBKCiM7c
nTwNwLxwlpe9eSzc0vPJ8xokAaUA3K3Gjqs+HHHyeCBPEYeKcRyjGYzT5NR9eKzX
WCo+LlqCBzGacPyNdD6VTJ4N+DG+3yQfK146bUb4LzbcYtIG0aSoGzNOaUgNUYkl
vPVi5jamwCXo1WeVlcOkyOBsyy/NVnGuM9q/MJKV5RsjAanh4GQrmuwfGLOYYmH0
fQ0ELaxclPkOfh3G9GgD9cAIwXvL1EXkUWmUy9Hu0fvSZZ8HCS+vyIa26R5x0uH6
4Luw4bSlW+SlurAgwVEsWelC1+1oSrFpAqg7LgogQxEELV5txu39+nINZHazykOQ
3pc9FCa5qm5xoKpx7A6PiRhTSZolEiSZbryEnapGd4ZXdiK83+Awl7UYHHloaGWt
bKYhDfErytS49rVBSwutsJJIqVzGDn17WnkG7QHrLzTn5cWd8PjociwIZ1ocUfZW
d7iQZbpdMX01/a/N4vD2iwZfaAprPqRuMo8kijAOiyOdQfG239DuQ06D+oGwwZ9Z
zN0Rs9/kayuZA/oEtEmHqq8ALCxncad8Tq77rBg14Ff2FuqzIxvzImsD62epZUTG
AnT/WUx3AVuUdmrolJChrdPVTWwacoyy2GwRjL3yaMJdDNs8KLxKUkZ75yKtYFpg
bqqpUNbEoRgxwBgu9eVHkuoSFvFan3R4dymB6jQv2DMf0RHWmyyrMrI2twma6ssE
nSbGDr/bwRkh7+D1AKWJ1SVBxd906HKEGJ3M9115A8Co2qvfJdpRWKMfwG+u8mCo
QfGwYb7qkzN4jNrh36iBL/tv4ScDsjKE2lashoWte27clLx9MHEuw9kyaRaMNIA6
Ml3TAMyFR61riIzj92dnMvN3EC5ZTtdh1T7LsqrKSP5D69ieZehGuMtrvMWEyAFx
GuXyetdtFOeft9PNA9fSqgPa6vTsaL1313SFFBt0WmGn8PQ5vDNcJZTgWPjYEIoH
AGugnG/fWUO+txYDCyOIr+eXac3OCaMNcOZByXyIfadpSTVVbRQuV6W9VD/rlZ9Z
KtoZntZHrfhnIImduDv9ngsrDb2kzrZXXpE1RnFTMS7a+94gJAPvmm+MzSZGgmb4
JNHgKAT1iIfEWdP0BN2U8q3LYS5OSedeigZeU/k2PmcQ1LL8OQLpZ4pTqZd+1UK7
0elYEj3d9HpFYfqYUAaTGuV/KGUWZjx6F7ZwSDujKZcb8CGGWbPTcRh8aXD9mnLi
YNFcsAZuYq1y0JT+iwC+aUQoXhtufjndkkZ7Zk1thM4tFg11YFCFi1FvpkjzUEej
m82dPQ4XaDtRlCbI8TLtKXt6AVhOFJuvujd+NN0GsLm+Rm5D+Tcpzb6dSCFWOSIi
KWnfP/W8PQGEX+495LhozPYg7AO3uQON2D29Q2z0Riq8XQQOFct7EmXQu8/2Jms9
ozVQDZktUor8j/FrbdZm33qjqfpk5M1sFR58h0I6i9FYMnWNGUmyFa1aJu+lcs0y
XyXqsEVDzQMv9JBZB2l771w9VGQEcf/L45Yyme8X7Gtcgo1dBgiwr5rzifFeMKl2
9b3jQQ74fmbkg1w0T3pWsgDZod1zRZpxDeiiYvUsP8xAUEDfH1xxwDTURbBSRLLL
+OmYbBjPBNRZrPVNCIeuBZiOdmnM4/A6LMabwFXDkzvqeS5t8g+JLyd+RVQRr8+s
F5mesW8XlEPUz6tUrngYNjd7+UCleOSDUEUtcGkZTPEhmC1eJSq+DbUbVCUcUSTz
W2364aDFPg/ynYLvaTVcdloxw5700tgZSCysxyORgSFpngWvqctoKioXYVdx3fcE
IuYqgT/m1rmZ7lcZapsNaDyCoOLaxvqctHrJ4jz5Dk1r0+fwmryQ+RaQVG+iRj+1
z9lBLsb9Fu41+CXb2wmlwjmnIb3BHiWSdGoWBR7uxrjB6FNgUNMW3ssmqNeWa1H7
CbMVdvonSEiGZfaRfT1yzRLfZEbtIWjNMcNdDl14myKFMKM4V6xQu7PU11SLcv2n
/OZtPzYq0TFO8BwDhz66kVivtfbOcWCwOICQPvgYqs81YyjnoPCHjfU5KOmp75ao
GgfYqLZgEIUY3D2o0SXTl5ePpaIUWAIoRblXGhbtUignq5dqNkDMvE1NhY1EzEC7
JLbGknTRkqA/zokPKYtzHQ3LuWPNP0bsmH93JWAPio1nIdDggPNg6xp+eYT1tqwP
gTLJ4PrpFROKCsCKdEVKhDLMEG9ILQIlxPhQh/y9Jmy4Aj8cfpsQWbrVSB3dWR4x
6DUTFiwEQoa0GdRvnsMJD0x3DFGSTchjgbL67Vwbp8/RHYNQl/H8al1pi12PggUS
66zF0JweIK1thGNp5EMHGbrTspsITI87OpvVomAKtqGSXrrB3FZSrXL5s1ORkAvB
hNGBXMsC0Yc8+EGHFqmkyDshd9Aw2gAzC+iQIE6M29ok2RVRRSDYnpaEhqScAgX3
0tNYtJHIVfwYSrrFmPO8K29bTGsXVfFGmVZQMPXcjQpE5TCnoX/K8/NTcwsshXtQ
05e3vhPDWfJGR2mCiZNPWHw5UVPPQB/6kCqchundPTg58mQ4041Khb/q6AItkftE
1twaBdNC52QBTzXq02h357K69kE9L9HnnhPnBsICLvdfTn2A3FxUdGZ0SzU1Z2UV
08QgI6r4G5TtVstUgaRCse0nzT88CaHSv9NXFOJCOXD79AqpQ+sUDJQHF9OZtCQC
Vr3qgInktNVhXoZNGUIJyjHSd0mqizxDgT2J+Uxa23tau5nFXqmtsApgDRr+zgt3
ICRx6p4/6WZ+DzA5i6qdB2HC4nAV1TcJXeJ5KWa/JdUznF0IDsa5hxn2agWO8vb0
4WT1vT0ibS8miM+fWQF2ReLOLG2KsnsV+NtX9/nPqOB8jBpajY12fPTFSqnmUuWm
7uqRjSWXB+OipxrgJCMSM3HJNYht/l3jCL2+lHYQ8C7/iR6qFVmZFnvqpAcsq/3K
6RPtPJSGLKtcqhJckEsB4XCumm0qNN/r4m84Iew1kk31dxuBbQo6+iXzdxJZW/Cj
4SV0VZI67DOmuQzsjQrW584q1HWu4/GzYyAvvT+IWufmUZcFA5T6x25R56qsAoPB
lGdi8fmN70m3o8Xu102IxlY928nrvIhoEKevooKSSqh7T79r1TmJ2HAN96iHcipW
3lNZG3BeiUnwe7XpISpMGG1E9aDF32T+VUzffwZDre0a0aB61ljthdG3eNQc2G2p
z+60pM1bw6k+ecbLZkJhVp0rPHoq618GyJo/QyjiYQIg3/p3gxpgCBDDC9yMp6cC
XX82gKRdmGD4MI/yuKLz/4xBFXtWozdukHcbWrGYr805mgqipeVs+7b+jC1skINA
9aTLtkfaIEZDodltXHpUiniLkDbvR6d4g9a1UIYhNbio6+t46DahQxjzPP5GwCMi
wJkpSEsXUpr4LPTduk7ChGOAHf8kQq4cCMYNH8hqJpgHUcbDnn0NsKZZqoZijrBA
lcPivCwL9H/b6nm9GMLLGrfg45WWQWfz/PwMHJtbaQpHCpDR6KXT/tAfRW/Qmx2j
y+85P73edn1I4QwRWcQrRhcDHmvonNLwPyt1XMykqKx9uiCVgjE+2LkzOtRB0ZlN
sgolNU0dNtINnYisUBLgHpmQdiIU/OdvrcSuJfzY1GaOQ+rU4hdWT8mGStS8aE+S
5UG66sHCkZT70NjiDvz5Fkf+zQ1A1Nz5AAuSlhCkl1xtrnVuRgN0GjEZuWAxKxq+
kwcrDiadP+oCpyBxi+FOYd+YgFi62fLUJmZFAM1lDyZy25KTNKihcgGOSnYKegXv
dIghu6OLVPTRdeOWmF3FdMCYK5U+m2IIG4nvQ7/QRc2gyPmcSOAA4UZrWItaDV+H
CUhy6Td22CFQcK1yisWrGrlQaTIK18/sPKvplbTHC0nkXxtpADYHQ5oHanNj9sot
8ARhSY/WIr/l/KP7wtuYbayVmlED4AQjCHczkT2rLRgRoOA9/79tzgm2VLQq9dDw
VDmhwpVmSc4/ca2um7RUyVtovMrNKY84tz96Zkhm40u5rY6eaJgACBRrqKb2Mtst
fkSM0AT3SPatl2j4lsgtHljppUHhl6kF7SkYQ3WAoENBMzunaut2rwVBqMn210zp
NbFD3TJ5/Hb5yxDO5Vtf4q9VsLq57X+FErhN9zLpliURYmlQu/XjZ5d5QnzjpvkD
v9pD4NDv5u58CqKfKHAmrkMcpcAOycv4Tlvg0ToPf8//0mn+YmUXmocI8kK2FDpd
5ciU437RyTCd/N5TpsrbGLUIRHL6LYjlaSLdtAei2L1oOoIf0tB4RNYNg9V37KFB
G90xblyVgspefwwJmmiALUH1YUt2m1pInX50415mN4n6uNwF9OCI4LD/2AW0K87V
sBdZwdFSkRiEc5C3k+X2fPp0YZA4Z0oJQ7RKaAn1311jSMDE8uWa9y5FKyeTQraF
1pHA2NPsr/ZJoAuON0kA57I3nQTyVVI2lKgV84J9dH90ir+HxSIE2Bc7IRC/xaa5
jisQGha816jhFJKTZmXqGY1Hs0gRqEBnR7SrHgOz9Pgf4LmvYX+G2nwjl6isRMX8
CMiqXtc7ANIO8oMe+tt+ydzxzrsVulEWA3USUyVMY+vPXiD9Pk6wjkbkqeIopJP9
f1rx73YUtJSJR5u+uMv8UQYvLI/G0weVJE8RTmlPdgSa0SDjRLmqe4sZgKiKYM5E
D8yRk1kQz/dcREjguQaDy/CS3GtKfsZsTEp6WdNOCP3Md3caQCwImVz86TCyXGgu
/FZ1bhClmHHbPPq06eW9SORfyJhu/zgXZupRje8rIDe7JuehiXB8qOlH6qcybYpm
T7NCJXAoZbBJQIXYcFSyD9MIGfAYcDBLaBQN0217vlVjKaV7tquOpvezY6NNE3NZ
HCXW4DRrIhTO7UKsWET1wn2v5tJdSX8h3lDMOOgspFz61bv+CZbg9aNli6Y16Dg5
Pl5yxCbR2tB+Nu7H1sCgwL6UuzwmZcqpMXz4Z8ofj/iss/kzHhSIAxbGc/tAV7yH
CZV51cxo8K/hu39hXrJm+o9ID3dwsnr46A9ht6wn7lInedhRY8hkQqVpwzX9P3I0
81hYo7OtWJqVWc7+5p2EPZVfOM/TSXvKoZLhmrAEl9zjWzuFJuuUvs7yZgWDCUy4
WB9LXlu7VYfYn30RJ1o8ARvcBb/i9bkYdIaDHi+daLI+lvLiBkNJGrjljMMLlAzO
c7g02DVzJU5WVTNper6uncHiiFEOos40yAHNVEqRwNYpOBLzSDxWQLzfwmZhSBoq
t1ecLzNMPviBXPw3AZIfDeFi6Nirmd7i7rwWcIk2NaqK+r83TCAQ0Mfqtvd/7O5M
9xXykSAQ7LTgqI8qLUpMenkBcx0Jfaca8mpCZ4ipUE0OdFxdCurdw3AlRaot0ZiH
a+OWCGslZz+JxRgangGzHDAiS5fOGssnKNgWz3OAsMf5ve7EK3CcIT0hMIm1SDPz
slN2Vk85Q16x6uXdd8SjT4Dnfw+Nf0ZwG6hgCDdADjyh0ONtldMJNa95MJFajBBE
0M7L4BD72fQrT0hPMTrrma11tBaDT4yNFcCLeBMyDU2+hnwYF3fSkIJmhrJBJ6Iu
7dxw100JQ+5UC4JuMaCT1lR4sqqrbu28vWNccvMPnD/KT6dgP+G1hbIIDk4/WyX4
hh9IQWGsGuzp26NZyTNIkpIyV3ZDNs3cNeSEs1iaicSoXgUO5UzXDQP8fgz+yjgG
b6seuje1RnOgMiyI5p1KONivZAqilhk3Po4oDAmZOsOK0hn3yMN5Go6Mht1zGnMF
oa688hXNYgd8uLNTgoaLl7rEYsJCIQEOsKsOkN4njgPHZtIG6rTfTNxKsuTCyykC
NDyTIwm/u5dVgWVlV9kForjCGvqj40vIqvAp/BMUiSPqjSmnNskwI1GODZsKxt27
4X3/pmiaiDVoYG7ixesycMNsL8e/R3xg7V+aiM/M9XJ96770Z5ONm47tKKEtqXNR
kobh0Skb0zmfTmrIKN9airk+8Rp4ucLp/Fc9eQkMBpUwTisGc1P9arB+SSyIwHcc
pGFsZMNiTor6yrfgmhM4DP7NHnJoJkD9JpZLMgt9fV1VXjI6/nBBG3wSGiAMV37W
MUnnpuRC/LtyY8AhTI6miV7W0/2pkjcEWrM4NTPMKNiaOZsJoSXkXGawhKOzlOQ9
MN3sMg1gZznkL/Ki1kKDcfPsBsx5uFM/k7f5uN+I9sX9bo0BLyqLPdCAMCYxEoas
JpmSuzhNHXfmIRpggxESpna+9psNqHqnQJasyzWBGg2xNX36ye5R3p9KWl2IrsYu
1EKLgNc30AWkC5wkVKZuwwX2Xkje4o9R2yyWJsHY6AvrqHABAc6YPp8FWcHDw3sk
xd2bJnGSVAE/eOS4ctU2gbq09bLSZFgc46/iEUPmG0ACYtVlNICC7qwkeFedcebx
f1GoMk/wE0E2qDuIlp9LeCNg1xMDZlLYR7Xl8wkhOPLUydOOBCb9FKIjuMfu3NJk
v4CtsCRE2Alaj+1xBPUdvOo0+j8i25wEHI7WBYGG8OSlGdJJxJDBJ09MVlag0lUj
mZp2k4waa6kmcpPhvj295JEaua8xCRmJ54e1rfT4QbfcQgd2RSC6FDG8sQ1+GMG9
1tKOaBILT2uw/HR8p37phHte48/jBy+37644lDKNNvz9HsM6dz9BfXS7Qv4n9UPe
q79msI6dSguQj6yEQHpIlE81NCzkWcphjUfn7n7tT/aUFdNMJqvBGWqLcX5zeVfa
zswk/sXdhULvA1U/eTl6FAHNBwJ0vVe4qHnAUFawaFNWR2RCwY04DALBI2Hvuuo7
kjPK/KiYl4e8fA/vfn80ly9nr6veqI3dgDd5BwNM/mA41Ivbc0lsQ7sm3oChiyw5
vrJDzWmwPTqYXBkvg+ppNXUm4Pkz8q6T/N1Z54yWfuz0KxfuYgqcU1K7M5EWJ1jg
VMJD9Dg5LP34n5RaDwWcHRD1Cf+z8djWcd+S5ozPulmP18hRFzBrWT8wSBQtMyda
gmt21j1VFuoTiilfoOz4uUq8nISmeYpd2VjoQ05epNfoLynBjVoOLNWfjw7o8/d3
NYgHaId0p0lPzeocC8qHDuvZaYficFVTRsYwZ5AE4NCUw5MURF7TM9Gbnr6M6Tgf
fiZc2EKcAfgASITp8n0/e7eeYxiDSmR5aP+Y2P2U0z23SJBXJ0Miz+2JvR2s1ko7
UzX1ckKirocMtBbkPrKG5V0ZiwhZTKrGAWyXKQixnpbBRBoaBlR5T/klFlL9WF8w
7oPptRGpzQ0/Tzkavo+VbfwudAiInkHgks3tGfX+p1KzJZ9n3/TMybegwsjKS8v0
mesbS2m1jXEY5BSlPL/rjTmbfJlnVM5VYpG/7cSCd3Gl+dLvTzQvH/JX6iATiP3R
inrCcXVac06pZ0rw1y31heWeWo5mll17fgwoGRn+7hR0Clg4z5+5B2SHLiF0t5aM
OBvXHfrnTHODpYV/L4qCE6yBbDc/ro/+/6gATwia27Q43UzAOYvUrKcaiEJdZdiC
UNRBf/r2GMMMuFS0bQMqrn8FUtkshgiPTDia3vQ1go78VWF9sMV6oCUbWcjEQkq3
p3+Alb4N3L8beM7FoSkgbl8fIlLHp+b+xU2xHffw+pnavdXG11qoQQzbhV83wIMy
zc2oScfo8hqrGvLrrt7FxrwnjZ8tW/xb+/mOfWRpHjNo5YckJYV5OpBvuW6T1h7H
cHVBSXSmDk/DlWqKRgppZYN8CSWzxJgUQGJvK+l8g/hKkUwNlehBTYYfArURdqhA
7CGWT9v7qeJ68BOvd1hQmoiCJeG2hgmj1L8jJQKFTRgTdGQZkxJ0MSOkQZTvsj6d
sGlkNeDNwSkQRDkVX8oYk9aKDDkL67//FDjq0j9GnSNIzvb1Ht/qpGLJhchnv6Wk
jQ6I4Ilq2wPun01eHi3XIpWB3svw0HmO602wV3b1BzrEcgxYv1Jid5lPPbP+GgaK
d2b7grsDoTTCgOPAncVCuQTyPeCvyFkX/s2wZTg8MLIPA/Di1GuTl70+SV1Jlgfl
pWHTeyVzBeJpad5bi161jd9UbIJOffwOKBK+BJtvtX6T+s08yEy3ke9UGGaZWC3I
v1t3ZgKuBPencQQz8+CNfPeGdLQZ0v/56eg7SDJuzoe2+JRoa0yAPsnol+l+LcRE
XxiUN3XEYDcsyF/+O3JhhqDX8eui0RdxsUviPguCwbimU0LFTN+hooUCfQM7hprc
3lmKoJgp+q06FvGQgK9Tp+WTy8ILm8WD+rQL+dPNc+0BjHwFV5SsJGldz8xE3B5k
QY3DtcdHhqX/pQF5JakUtfxXV0vm4WNr/eqU3v2vqt1fepvcWCLh+H8zoQmBCcBO
pQSC86a5y6sGvWSNHEZUyrYJAvSXXXImpDAPtzAwWt1bomlN0VljMq/Hu9ouPq/G
dhD8+lCV1WAZtEKzvB7l729apsdEOn6LyV78Ypjs6HD0vUN0cPWpHKHOnDcB3pmm
NT8qEzQpscsFP7qPu7K6DnjbnlQnbJsF0E/f+CUDOoP5bYT0fVfZNL79+Y1eWvGr
4sw5lqFkYN+7gI5lpAzs4TPn8z4+pK+RHgTa4c/rgyYkZsqFH9Sz7gPKA44yoqOW
jZMnkHZw0q367nUwrfdgYidAXhN0FPIlv4BRaYKiIEgb7uR9O/HcCuw8OzOTrNZz
RLN2G6i7PgO+m0y5xz/iVudU4EbF/TTDuyI1iGW62ZaB/YFBoGWHDyOOkaflVDhK
fs8M/IykpaHwBhIqSgcVhXiKicbAJES/2SpsjQs4joEGRg1ObRuSL8cHBh4m1xQe
W1O0MNbQeXbtcBU1HWtGbGzqv6OsCWFfq8SYwtIxkLz3DQ1ARz9BSHOTThzsStWB
pKsV0bxKyYewDivPTOTtjqtokHs6dLygPcRMWolADvX290Iy9RCp7qqP6xoHXLQN
gBIv2KpJ0dHHgD6+i5eDH4VJ3iW2bA/cXQ986w6NfDmoHDQqR+prcP9EGF9CtkmJ
TboGRjvVZriZC5/XWfgEW4KNwjYRX/cCVZlH+nZGyJuj+DZJdkQgX/xbDVy+tPAz
bg/EMFczTyWc5Gw5ZJs6dFAlc/fwW4MBBNEknyWFpVFT/OQz9nbBrtCpW+pVx67w
RWHoUxFXYTMd3AL1L/24JoBjZ3I998L8fZEvy6PSHsVmoY6v6dLH9mA5BsHdOQal
ORhIYPBY9zm2qOYBD8sdjzVltXKRxpBdTSFSgfVVCbOSkGKE2ng3rfDHYYO9DXEv
lbTIvEVfUk/Aa8djlk8G+VWamZbikQL/RFHFB/GUg1Kqe2lylKwRcTbEO6soRDdD
I9ZdgHL3RopeGRYzmyHq6jT3iw08LlmzQyBCqB+66negciwVnzohSBNIhbUoROfS
IPQYhd0f8IBjRDmHQk23Poxg80MPFtj+/8tIYiGygvQjckmclQDRT9SR6UCKx8BC
iPl3d+s7G7xiKGUVMMVZWLIeMqEEmxqx3k4/o5x43RK1qhFmEu02d6a21AhQEsPP
nsPH5SMm+8d/Y+UlpS80urRLwS1AgKisq5cQqYxcXLmcyq9MT9H8m6nerQBuHPhE
NwjiFMNGA/91bmMO/T5bVW+zJGq7bWM3hDTaMn74tvG7Yoix1qQvQAYAWIVwi+om
lJNA5PEuHBSBss6+2h8bFxRao4w9XjLQGWBWEr+dRirDXN13MlXBKpZyH7Sug0kV
u2+pLGcLvm8hz50bdU5YxaZYsMpR2JAk5PRqSmpD3aQjTPLNK6GUkZ5O8irdQNSC
LguT8mB8xmX5JfYG46mcknOznLVC9WdX7Opp7w4bSswbQ11FJWtxoJdCWPYmr633
4CdEsau8sQwPVL0bFTOnKcosUB0l0CozrbN6T1HnIXnufngUsAP47JKm/I5eAE6m
yngliAvol8Mxn4ZDa4cmmsxm7JLOu6kn/dryVMUtT95Jp6tTmndPFiydZwDFAwIR
x/MpCogvdfCEcV/akv999BuWbe8gj/ucHiIXaE+Ikj9HJvt8BrvmGO/JwZ0pSGhd
k3HXd9AW+nsh+cA+xITWqqPaIRtnVbWddPDHDKjpTpHaqu3UEGo2Oksi0Q6EgULO
9R+1Pw2hHIC9CXjtLLbhK5oI5H+Kl0xDYGY+SrRU1w8RUewCjiN7SX9ASjufVToI
HK0+Gth+1dz9QZJxFRlPZu2eSOwiz3nSVG4jqqNuh0BcNmLXPBr1OxnBOULYVfO4
uYofThK6/nRUD0LsWzbDzrlufr0Ob7HjKdw0J0UTfIGB8hOTsxROlkl+lXqEITES
cOFzj2/LcviWxOXGJkT04J/uM49dBTsEs+AcXawl0mL5Id8PIsXKcyJu7sXPsR7R
3HlmS04D0MdNLAsMJEC97Nla+Rh1hZBZXG0/YrYAj1FPwFjrHlq7rBQD1AXdpKu8
gn5Q55B2lZOiUjXjzPrTud5iUXLFc3xKgHmgr9EWuPgmQCfIqOUtDOE+TSi0nCJL
fV7ISwwM/d8U2NehL3uiCwOpBvMJOzSFH7cGlKd5sRysD0FCmrlMR4QXdiVHoJ70
Oq0fiiX75DuzyJj2bQqxRpn46ePz4Q5t0SHjKMzKeak2LkAncEmCEYS0AdDZTKd2
tND2oNjg7oMcCjq41ULQ7ASFDalnzdn3cohPZZ7tzd43mK9vVXEPfBd5cJwyijDY
yrCLvE21NaJlazbihsHzXR4LkYeXEn/1gb86DxnIVdVbku0sqLYh4S3+468nE50A
G9p2pJP1xYltfixQ/PevrBpU8wRHvzdc8ND+SMYZJG02CMl9+TjiyViK/H4DNmrN
YhgFeoPdNs5GqbWoeD9Fykuq4MhbAMWHin20peM5MqM5twe6nxs7ArI6ykjNfBn+
TX2gtvnLjj/Y8Ri1E5pPqNSRr+bofZiYiJj2t28c0rbQhDfkJAtNrJf16zrTJS52
ABdp2+trWXryVTu3c51xWJNpanaXWCEHuNBAYp0KP1GL9yBpucU1Fa5tLSeFO7/p
QewZMtHKrVuncnwDUZ38PRmHL1Me9ERMzj1wwkor5x/ZrzMfm/3HCYwqeAMewyMl
PmeKl57mk0CbY/198LDzUd3sRIHz11007GN/jrgta7JjlvcpQ9v5ktVh2miOBzx2
Rx9AVeLGtay+ItnXFwtUgCtQiRVVbDx46LjytrrZ36yB6uvqGI20w0q0WDzpaR8p
WnX1RVhOzuSMMR3u0u65lAtzKBIS0SyBS6SMPKOU5cG4u3N8FP7QZDvMpxFZvaJG
5CVQ5ZgHKPhbY93rxZoMbZcGEh9luamOH972uTMd7cghRBs/TY5u695KpvP6JQv+
XPDc07mjF5C2hEpo5PZhUTT+zCXU23IhmRNOPlpikYq+bJrq68r2AjzSR1syqOKZ
lr5ppOD6l2VyUl/l4LTYK+UDFSqp+RjxCZsnQlUQGS7RiCgR2NvU4JRBfq/Fe+uI
6g37ak61tby2CtpyII1aA3rtPiflbOx+o4EDCzTkExQF1wQjdEJ3xOrwwT5gU0jV
Wbt1lLcz2eZ1GVz6DtRw/p5UYhHQB6PnnkD8dGs14aQvV3QR1QvuS8BTO0ReQOkc
sCM4YxrEdXm9wSdZpkxjRXi8bEisbbLVyr0RcsoserhnvxcZ0EXQk9Q879ijMx9F
oeiMqbjK/A/6XN1KrpUco1bY05747dyuAMlt2Ij2BhAfxcU+Ikew16mDUqihqr5i
NP1M+44ake17NY+z61RkbCFyN8BxJFXj8YmFfysgtLSQwJVn+5rzRwg9tvYdwMPm
tKtwtjkPumcVZiW6gpAbAxxBC1YGZAWfOXwb6wDBstXyPWM6PMh3mC5ssZGBjA0s
Mx9pAFlbbyaS5oAPkmYxQ8SwLZYzjdHnyYkaZ5zrGbrFjnAsqZc1eIUZyyhvs+Nx
dsVo546/QG21Cy0mYtMK9hM1yIL3ct/IkX0bZ96fxrBKhQNogTqHrVHviUl2qwSV
xQ0HHwATScOD9BihrdUngsWd42onBLK+b0EbmdWvxWgzYMjlaDlm3oFyS8Jb2yYz
E5nZKK4qVd0Ik6qrSW6jOVe55ZeJshhj+cR/H3KiCBFeusjKFUfteYUVnkogkMcd
oKvl72EbEmp3kDdWiGZ1x2x9Cr49n1M4uthGO+FanucCV3EtHuUaBAyzJNhvNslO
lvAMXXjV36a+RTlMD6hQRMKBwThlJXvikkVj0QWBpPTwoE0Lxi1WIUquBJHQzAyw
dG4xf6l16a9XnAUNFb/p6w+zRX+oFDFcpwIhiuenmzU2B+CQM4ulkFR7Z0NzSxpe
HUpULjQDH6tomQ3Z/oWXLQmvOrF+uoxtFMWJOnQW4bSIkW7MUavvfgqKgdnS1D7+
BzTn0Dv3pKf/ltDbVRZlyXzg6LUOau83aROucgHNHTDfBOX92FH9xerYJCUHJb5v
shQfzqMJadNuek21qxN/r3yYCOK63+OLXgu2ZXvP/clD1eawbG1yRT+uaMDTvANW
S5fBL1tj5S9zr3tT3jqEY+al0Ast2J5MJFEOo3BLN06+G0Uyfn6CfskOHZECRb4h
doJiP408Un98rqgMlF1vxovLJ3rhKecb4je3vaIXlM+/NU0mV42tmf7fsY3eSgpO
/bH1JdV7SXy39I6loq2/Srk3wlLYHU9ShCDiH9gxfe+LWHC/8lbQMf3ep+pTI68C
kXcF0oeEJMbpuYwn3bBPGKzEBCePyWiIrTfBh0PR2fR0oyZb0Vf/yUBjNZv3ieZP
Xug3AuMrh6yp6Db18KUSGZnPkg8jFtRpNs8IvwVYD8BwI/1uipZU6FkGGdPWqszR
4mGuS2bkuXqJ7A31UZ3cO3H9WKm13YfsDmOoPUDMFE0JqqxpggSLOGhKIDDQcIK/
zC9pAHOI0FL2TAyO6Cshgwt0505bKdVlEuPNV545xRM/wa9TfWCMpnCkcwB/Z4Ab
aaL6YoWarZ6wn/ZN+tzHDGrMAy1nel0gzdqVkb8KhmtrlLNTC3sYJqUFo1kgy3fZ
fDp/lMninCBKAZO116IeYpw1nGzShHjq2Uz9EfmXJie+N7NI1XyTXzQjB8E0diEy
Jx6ZBDV80+Hbpsif///sYUTgxGhPDUh3KvGf03s1jCGMOu3JGPQtUushc3iD1tem
enoZsWZrr4NUvmH/p1kwjLPlTqEXhqWzhnCDP9ROAhV05mF5y6qZBivWONzJjfl7
A1PMHMh+eMO2bfpu+DMYvAfaO/7G176qJE1dUBCs1aKmCudAvdr51MUUIPdHXSmt
sl0ec7VgE7sjuBQLat9ln+OCE0sAo0Kg8MQWk6lBNvr81bSANQKxUqwgE4UnjiWp
JaQbLZkTyhHpFCZbW3EYG9XDhcD/Ld6ZSHnJkciny+/Vh12ZuMvBpCoU1NyVNFbo
HbbBsEWYkbFZBB+s57iikYBEtEv4Vv8xFWmpfa0pa4uF7YurENoM2Ni6OW3fOJQd
2MonqpNUDU6nSzmJ5pWk02elGDWwPRn4q6p2fb/cbcMbX+tiy+gYv4l+uFtJtdAU
ghb2ANR4tOvV0nwVHY/BHfQTxifpBX0oC0kHrwZ0t3o5TUN4/EbCbADqOdKhIZZD
xsDtL9+FXtF/P7WdT18mLhhA7tTlZGV1sEzh3/rwkxisE5DX8mneSfFAGpQFk11k
l6b3g7FhkxNylrpd/ioskNtOLZVsl3DeRKPdF7Wtyjswmxymrw6l5tFw6dVlKwW/
gf66AwnwnZ8IU1MPrves7ysKvPcKzEGzwM1ek/7RmM/bj6BQJke4iNhkDziBA5Xa
CfZWQBJ0b+sJB+Ei2p1hBm7St0BCBykSoGYN9lgWdBTZB13E/RpktubkrU3cMpx7
GxkmmfyjhOJTS8fvcKkBfVTp1GbG99nm0n0timq/F0+GFFyUWKPCywpUVvp6ya82
J0ATl8muVeq066B2D55bTBRFxgXJGKAAjtwmoVb3kl2RUPCxgAKTmtlkDuqbhsxa
qn5avFUw02MNq7L8E+oChvV2UbSggWvm/WcpAau6YBaMzyIhxVTcg5U0g58Iw+R7
yhmOaa9sFGXKidGADgBWggvcDNp0ZMaiqWRqPCVMtotJIdNQgo09Sgr7nxwv4ESY
zf/B1H2a+t4gFtqkSzY+L5mckYE+tbVOc9mGa2mSl4B/PWapFnoVxgqk2iHQbTfH
l62i09ltK5bcpFM+K8sGF+5YR35KM0/0tsGLSVqqUQFyPri3bG5yb72E4hw8N8zD
N6DmUjnTSC4BU9ayFsBi2iwC7EIX3moK3DSNUiSmYYcVGWtWrLS933jZI8/F7X+N
9a631XFoOGWMH2gccLtupES2pxbpNXzFi9TBkahcilHRMZ/drC8k4PFjamKBO2HN
2nt5dBRc1WF5GG/rbG9QZlYWnlDPNrwtFgIg7QeHiuG8ML1AsFrJLDsWY3D8Vvao
gKpTZ/A1dTcJ+rzvQSQzRQ1uklvhvMfIfLI01RqxcfXgno2NyuHq7wRwhhNP9piV
BX4bWJX0wdWBiE/e1JeD2o1QKmdatW92duSpDIaeeh3KEcGZ4BewyaW+hAnPQYet
3+vhtRIEQG3MsT0x+r2w0PqCvX3btX2y6opHDNFK4ux7KDEFDXbMplregjONFfcr
bNJUwkX1ZALIyp8BJEB5tX6yyCD3KfxAP+3mFQEhDBK37w1hnSBMFV4NDrOIfwAo
/28s0dpLcyS1FOoc8HYHRrvNTFCDQ7xf6I6SnxJvXKHz7b3MfaPcW4HOxLE0gPTc
nWXDlGxJiY3RyNtAoJbHTFNm5Urse+1sRDJcUpfwSJ1UJglomXP/NfCfD4pZVexd
wtfaFEEjaCA4ymdayNobX3x7wak+B3ZHgG0E8zMonr1oy1rHFiaKP2Ipd6bKEe9m
0Cg/9SU4c+qbEfcwDtWUiHMWl4j8IY9M9EQkVYMhWWK3N6obWMDK5Tn1l+aGpnzC
O32hhwarLIjIF3ZN6xwKfa1CvgCOyhUQI++pwWubpGTJ1D29XUY+p4LeukZCs+Ds
Ly61azN251OfDTNaRfy3L6NOqjA3VMteXnBvJhctDsxs8eY2YmeWFbrgIyYDZjwv
8XPsrpjtWNgS+WilrmqtUJw/HH0syTk2394vFPHEjk8haqyiEWBsXUNpa3eMca6g
vu8PiwbM8OY8DuvDuB2oGNRUFmA1wQ685sad4pPH7rimVLzCL+mCoytquvNW9+E4
l79E5Zl8JeZHj0lnNtrG4Jgd/UMFhrmuZe74TWplz4BuQA9OkMfR+TkaK4ZJSggM
Lep6f4McOJuq0bVsl3R+Gc9kihBFvjP0ZSMpW15yRIX5/vH4R1Btzxe6iJcdN8mn
XqN2cXBW6BIkTa924NbZWGQ8hejkd//LxaVND/s9HkYUnA3/VcVFYYf2hGU0JPai
JjfCHEDZ5NTfQeVsazhiJuFbCWeJ2EynXl+Vt8NhBpaswZnL/e4WqnfbWll07ALw
LEMKrMkKiu4yH0gcKl7yW8s70ocTm8ZuW+ZScMG2VMzlLSj1XJozs+Fv2CZ8ZWTt
MdtZmGzfBN3FPUYLh4yjnGrc4dArFmw5uVoupM7OpFDPCut7pakYTvWjPOuu5Oxh
JVCx9LHNtUwCUrUVYOM16RBc9kezG+ODx5HgmYoym8X89Dn/lmBJzICKedqEMboo
Nj1q+ynBzCHhAITESMtPLrWt9/SEyC6QuyMj0Y5pmEzbJC/BFpOtT+L2XFymhemg
Hvt1uoLM4pIjN6gEnFjVK+JuMjGdR5fR1h9V5eNP+8XGl+eGhJvNsOin5fkTPGuU
n2DxlDqFCFZWQxS1yFvbPbrqbcdLE5u/wGclEB10GZdQZkC9eNQbr4ISv6rCyq+5
vgwN9CEYsLZs4bmN6/FOGVg6vdAC44B7Brq6xuXfsaZI+CEMkoTZjY10uHviMwDh
lYJyRpV3VtLSv8H61dPz1feGdUQ7zu8ulv/SlbDITZqUvlfam5/Ygcp8Tg5tnZ8X
XnDw3hU/PtQkc1WXIPg9wNimaIerO6yUrOjNnD5kEjx7HrzNiYOV/plQxi1LHDoJ
iP1NO0hEovKArWMo1CvOKgS6MSKw+EAVfIQbG5I70YvP8rTFMGg4jaFDHbhGzlhC
HnGI8+UGUiliR4tcxO1qiqGCDZsCRvZj/P14KJoCUmtgllzBWj3Crnsm6q2gEprV
cKC1u+UA38hdF7MEYnU3DzECcy0NBJev2emGCEK064NxczKz7cqLawQeKLStImb6
2zozjIjkHsQu4x0ItVXeQwIo2vOKxU0qVOTOtmZhmhz4juRiYZn3TTPpB1TLtF4k
Ryek4TPgXIvQPcYGNI9OMVn8dK7K9l4A/nhMk8Fg7uDobyd73UnFxm0bF3JdRgh7
IufESrmak2Tp9ju6SDXv3+W9rT9zzTu1gs30oMQcy89YWCGMfyNVyXdkYOcb2k7U
viIsziv9UPsM7HG4eXFdbSa9B2EBZaLYn0SYtlI05UxavNfZZ8ClbQ5WA8tbaflF
KgFQ3S5u07L63M11/fipiKjtVCl6QP4ZM9o81qBtD1tixJGniYzFMba1qhFlH34A
oiP3OkCVaZZxpms/4RHb43jHZY/lLx7OOwZTZB59QqL1l0yHA9zzGBrGhgluIqdK
Bspt16qZYdcC7haCrGq2jISZqC9lDlAg2o0YI+eG3rbdK7N0AgnraRw9S0slIPrC
jrJZfU+nV0+b/r+a56VfbjKRpMOO/z0NlET/8Owx0dYGwJYM9ls/VONx/1oMFuMy
fYIJ9DVAOCMsCUCmUKRrN7mjXTfDYYCon4bGbei9bw+e8FpuaO93pisNUt0J3QDN
bcGbJsd6wGhrCCmowSrtUzGg7vGMAgbXcUmwT+506/YGHB5KVi/qkPw+LGc580G4
HnyYqfk6exYIyRSJhW/mA1IAD8cg0hyUZHtMMl8WTjJDGDFmeKRDI4O8dqtLuYaH
iHxTiCtKrfGiEnNsW4uqnvuuqUyv0DDn1i+dMgzpaQ1MkK+Ko8PgGUqMgfkub9iC
xceRXisjzKOloSx8LPnDUoL0rMSW4smDXyehbZODS+IUHDuXIe2lEgkMeR/dF4bk
e6NNhFFKhYYpzasiHOQf45OLxQcEOGga1z7Kt6Lxm+YCZYCauYb234KXqeCFYJuS
oAty/1ozFbgCUtF/G6ne0+uNEY45uF0qG7Bm2yvhiVzKlU43S4+f1+AtF9BnA40D
nq+PR7Ey/DYm0phjEaeqieq8bAKQASx35htSVH9NVzHmCT9hT2+XuzebAujtS5A6
1YXEHXng4DPoEWQCu8zYeJD3AsvraNbZFPPPyfWNHC+mHDjrLRiHngMotwbEiizz
4ApX3MpkcFAacE1pbf9tv0xcksc/Pvp9xBglivjptKMeCkAnW4+fMjsLOLtf51kX
QmphMIKTxr4wZwMLVBupA/mc3SoObSlxvGDELvWwjTt6lYRR6uPgyauQMkrEfG5G
GWQ4XFpCZpIXPXeYHcGz48GcWb1lOr4rZSFazaqgPrjST/W+N+SkIDShe9GuISCA
NtgmEGycrk1VQk1jjlJKVkHawrqHWJ3cZ+lfa1Lu+wFJ77NXAJhMJVyDt/HLO7aj
8YjZuHry3bjT7lnPEsCFVg3o3kpeAzwy3ccw/qeFpmMF+l23GYtF3P8NFJjlg36A
LxCltLPAUK4vKxLQhuB4InEWhvc8XkB3m0Av9/ZWSTWvOwpk3peBn75GjN+5xfgu
Vlb6aAr+Nu3HPmeCKj0SvD36LveTt8kceVVJ4SG60TiZPv+Z4BOPSw4EpYAtCq/B
k3MRRhW7dNdtjKyZoYIIsblxnPOBXkdwCctrcjcgs88U0K/bdQf6Af1rqhvLp4Wg
GLrlZq2YJAYy/Y7oCcr416tYk2P7ZOsIK4Mp2jgkFfjnsyjFQKQyWSMNaGqUDDxU
8tq33IxXiEbIo9C9MxMloxKgHyliJz+kzSfGFBlHJwSO/TUl5N0Yz529j1B/Ryqc
HuNy8QZ/8E8LkXLbUCNMDDG5vf9cQRVZ8WRVqtvKhLUxM0yonLB1u718m/i4g1jV
7hUot6dkqq6Vyzh3iOx94pmj8bdW79E/KmcBo5YSyk4105uNjJOCta0M3zyzLymW
C8Xjuq4SV+/6Kcc34WgU8PGBdPoJLYycZyPySHYaPG866HZOitQGtCQXDx1QrD5L
Ce/hOsBNpkzFoQwQ5fM5Uh6UbCTNevMaKQC0v55bSRFsKjSDAlTAB/yJY/LSwPoP
ohkC4P8GKHgmGHYP0gW2rGLvVFAgh+Ihj3QNKBp73uzOZ7zw6MnNItyPFTSN3Nue
zdIzeuTr0wwnrGmBrtfGiiEwDgvUEIjwSdTInnlddBM9dH9w0GU31dgkIR47d/ef
XDRYveyRRxLq7IAwfSDsqszMnSOQM6pBtikBfcL8/apYYg3WLZEIrouiHMYyD7ew
QMyRAlhNOZmuUXfhL2n9XAKZybba2yAM4mgp5r/BoENGwCcb5QxRMbKUTIirDsPU
/yd8zk3keuLXK1eAz6UVy1AZ/2SwTRYTnI5fouxh7JnfoPP8sHM8gFeNtPLJNzWq
ixaNVhblTymvyDVLtiCZHMRSn3ccCckKBFWbf+abLzpTygqOrd7wbVc+T0LJx+0y
AvbNDJIrf4S86ZEJ/MleH2GYQcMgqxUJXudFUDSw5i8C1ad/wXodfc0LZyNq8Sx/
JdWiEWQfh+1hQ96j/ndZvEk23u7ZQautrwCgVm5w5c5SgdN9pf8vNTdyY9eM1zZZ
t1DgpzMqkOEpPW3xN/AZ6lTTzOv1DDVdfmslfKZB8JmRUSpCf0/ZzXJnam0+Qxnu
ZtnHOwy7Xd0a1f1OPkWv1W8yRDl3H9kCpBMu3WuetiJp3teJDgkF/1H7i4KiNfXj
rH811qvUn+w+RRy9G+EJpDdTjMq9XcfM1Bs5T0HVS8R4DW0A/voSmDyw/8KELeQC
VJ3UlkRiAWfVNz8zo0bSvLsTTXqB7gor676v69c/D6VSx5HVAaqnEt5oZ5N3QfUF
OB5/s20050F+KIKXA6irJU8YrfjvmlFSV1jrqlYwDSaVkHpfhhGvlKDWtlKWJYLd
rNNWek4i/1xbv8GRmrLicXiI3aAhze2lVsZVIfFo6pYjQRUY4BppbVL16ohYXSoT
DdX0oddD5mU/cI7yU2t4lsHjBunTTVhNq4H/09JgRgd3MzSOM1FCKlyIYZTS6fAA
J9LTYF827dttgo1z9wImH/beKHMrd0pYYiqih/rRnU83IqIRCpyhuivvX/FP26wV
h82KLNJrVOZSzyJ9O2AM3hJMKQlaMddBJScgAptpLhZ+lYiZIIEh13SIclYL407x
LzdfLelGFadQorjuUFhnjEGBxN0Z8mCW9cv4d9IcJNd4ZKWy6R+uMDezt9kS65x0
Tj4pwdg5bxVncJwWJieJ+W+cVrnjKB+BqlAZlAxxsje5xbuccvWoAZMhYqd/LI1H
0blkGwQ3b/ncABG0rKNtdY2Viz8vCQsGCQEnxJXlj3XFefxgRsm+okmU3IprI+dH
JA88jaD1s4ZbR+Y+451wW6UEdW+LvAyQ9GpVTehko5ZkfQKIOowV/nZhXfd/iUcI
heXS6vcm2XHuPWzxcarKwjIoI1P7ahOh+Lp8A8BHIzk0yStBG/bFzc53VpkAWIQD
rpdjKzVCJmfqErby8NKIuvuyU75AHkRRhF/NSnN3k0wTSK1dQ00w+DgKp1H/a694
qhJutksl+Nn4B/O6pm5DcoS1ao5fB4ZPMHug1xnUjYxjEOc4y0/vXL9Y3y7zUxx6
h4651Tks6hJi20vaG324dsfv/UI3prtHULo0dk7CYcMsEb3XN3DIIFLx4XvM9eef
fKXOLqPwZmxKIYE5GTsE7i3gw2QNSZZr+dU7vC3OvRp2UC9LGJd85d/IomU+WM/2
YhJKcGNB+hVb2RlYoW2kgqhVVDHz8Nw8AhE7fFaIBKPJykhn5yd4wN59kR51+Nrp
nsppujJek+O9PREp/i1+YH6epGt/+cVZyfqyox1fSlmZDTV0l2Z8Cxa5qygusYFG
bDD9L3eYtYHuNv5SP2a3jRVsEii999xm8CqltFch5M6ExcNCMepXZbjFS8QTI+1P
cWsoYFwEa1pvut0w9vR50B+XB6OKZyfmEK8UNFoh4kreOYMHvPZVUjFLU7NTzFY0
60GerlJyNEt1tzWPTMbJjzShCFq4avrnXBU3198xiTGptN/7uP2pPFaFNaaNVxme
0q8yaDxxmzrFsyQr3wd2Vq4GmC+GXG2eNeg2GFV+J6ezuXCPNRjGCqR7LPCVHaJv
I0zpzqD7Qk5EJNS/4TWMhdmLdZWBV+yC33fOj6W5a+SH9HkoQADs38DoMYKZAy9D
b78YUkoSyn085ogCp5hK/r5p08byqELyIoxjHRo3SADDpMfJU9UqCQR4aD/sUzv9
/uT7FVWAD0xH2cPqUbBJ0oxKO00swvoUWv5cadVU5wNfQ4EYPYatd/8t015xKrOM
JazBDXOFlQNuzaZkBTFB3eXAQpXgFzASj0mF+9Y7Ct7GqSd/tlspw1bNXM42QHK1
zDGKlLXqqJCxPosDOYu2dzNl2jhWDFVzSygF8LHGII2TR/IHSq76mx7XYZAhyTjU
0w9NjiCKBub+6ariD+pTHQ7ONCdNGxIiotxnr7jWY7jpkxdWLr8g4uKZ2FGT7NUP
YaloaZ+h39yYbLiQ7hioyugH5yUe68yddvH7v3+kZKEAY73rmXnB5VSVNeozdosp
vwTk8QURXOxh5AY+ywtDU4t31go2Y3KJD/WgRInUNa15jesb/9tKOkYHYFwpOXoE
fo1cmEWfM9bUpPBxEsiPZMcw6EFWSFgp6RTlARm8PRWbSsbIno9Uu2TmxzhqY8nK
FnnFiySNc+23ouS5jIQqyJQIWjaj1nTKdkagFOYuomGyJaPFP7o8kynbFV8SEsmu
e36XF1e+UQSJUBAw4fuZnlWLGycwMbZ2RWIqDjBIfz7kfsyxT/wnBj2rVa7kiow9
J5bHBAFycZj3QSSKZM9FoPCJ2Z+PJRQJPSCxcfxeR639e+aGVosAWW+xmRNHmBo2
d1H5dc3JGV6oNPQO2qYkHvG5oHv+De3PKqRYc2w70itqAgqU2Ho7uQsqFNPiDUcV
fVtmXKzs9xfhd9f/Y8AW9rsGpFuOSt8k8hWwcfRJ4MztavGW5I2w6G7fmoFfH2So
Tc2IxaVxGW5FAKrHLAcYEfNBNyaaZ4+qSNwWQ3tHcj0U869MDHc/dS0QKN1pw2r6
EZULS7NzVponIfcAwJzwRA9HpUUsHFneeN08dD6d38w69jNd/vJbvH0HgB/pvPg4
kL2S6OF89h0oKpTmOtiIzOu1532iUseOXUAtxcGzXLfuPWlil9bgx5IgvCyRHak0
6vWRv7AQx8SgoNzoDwLSSRgddmjjWWWY+XQGPIOOp+Ep++dDnKVxoWB7V7gvEv6v
0fnxzbN2P8We34Onekd9w8yxwnvlLXc2QeoOVrkpCSiLkhhLJLbduJ9ORYuShY3s
0HOdzPY55WnbxxMLPgK7CF2TeppYqKIpHfq9C8jPvrGiVdvLdVTsf55DNI28TANZ
aqwoDn6YxVRxJuz+3Gfm5jd/NkBUO0jQfbrFyY7VCdMu9t5X0zkKV2aV9iA1SRtb
hGdCGC0rjGZ48PwPVihVinEdXKX7c6wm4cEawBpqc2s/k4mT3+0zKugnmgj3Lf1p
ab+hf/sc3HZgSTtcofQ4cGO8e63L4VkgRrmM1c/3lU7a2UkFT2bxGxrErDwS7U7i
MdzWcqAJKi6xrN9PqO2+vUbZACh2Mg8iRMxK67FitZwRPUku/CHsmzx7XlR4qDsp
1c+CWNasHA62MARmG+FSk+rqQZv1wu9dVKkfPFzQLu7Xj4giAKU3ngjtuf91t8Ck
j/x3NmglUYisD5TBdiUSle26XLst0Gd5qbpGph1ZAqNacX1CGQNCYU63YIPDiY6M
5C8iYTGRwkv3YHlIWTfPkvE1f73sV4DG7X4d1O5LTHjFdwTPT1FFEgfneyP/HIDL
yMn+JtGYJwoEEBnJ39TwZLXqR8wCFcycLS9BQRp0MWGDKj+0Dd28vFCBgLZP4Zhf
heRD8oGDwMkuLdCOvphElDIfa3hjdexat2PFFLBsKQywKxdn8zh+CGni9HizENlQ
eqg1fxUQhQhdrZDluPv9R7cC3zp8F11QVE0tvFxnvnU3Cs9uxvAEKXyfGVdRoYwQ
eRyX0J3JB42UBZzkiW3emftoPdgv9uUtSJOIaXl5fFBBFvk+Q05Po5oFI/GTXscy
BWP38bjsoBJMbzuoqBVJPTMXTi5FuTik0LNUAFne45j2fn3zq5TKV/6xxxUvbnnF
GOUXZO1MK1/L+dxVb9hGC90EVK95Vr7xwr1ID77OK6XqcSXpV39cGQXs+tveIh76
mYokZ2c+5h/M92cVmig9npMLxgkXMI/86PW3/yyKOR6mPrvCVYmM2x/goEqF2w2b
Tk8as125lcuvVQa2Yu+EjCMAnoU/6HqGCYXNcZOml9fKR1p3rmC3KiswxLyngiNK
KF/PjFRIzcGp4P3Xr2DZ7XfBh2tBZT+K9qocnyEB2ED3kj29fIsnN7trAZ2b8M+M
p1VF1+91ygQ2o6jOy2NKOfBR84EyYCY+ajYOh5QRfbch2Cm/oPA/hn4/q7fxUNap
e8PZEr7nBu0HTgVIUYqHh/x3ilS8mXC6c+8eL7DHnwFbliFbKJvlEQbIUsHFOqe1
anM19ujkSbozMxJk5AjZHtOYJL0oCioeZn6QpSAVyEn+hOe4x4vBmrIbEnbQ3Dy6
gsvy29YWCqZ4WhDOR4MKMMp5Qxq9NyJGhAZg3FyDqkmaAULhYl4ffHHtMDrs7O2U
fMggpi5HbfFmGpohdSkpdM1PE85i7y0q0ZSmBOlrfLR1uzq99YrmagcXFKcb4lk2
Xcp9LFhMCBsKHVTziKKvOos8iuAAHE1+5sV5RPAG5QzdgBYbZRl5QPEZU/LOgycJ
WyTBr/kAsCRcZ9zHhXXidOiwohLyiqdlJmMq/m8umFh+rYwK51ofx0TDk/d8fkEi
+lwt7K+RMBsCEPBpI37x/hRKWZFDByMuikLCAJRMFst/BBdiH6QWkHU+iGR8sR5s
pyJ+I5M+nup14jxjz0MrfcjadpcfKghGtWAMpJFINyBluPmbVx8us0H/uuLFfP4d
VnipE2VVfqse4GbQbZZyhVlzoR6MuyST4tUzx8crfjO1ZKZ7jxNtiBmCxM12Uaj+
Zqmh4+qewFQztAWkLjG2vsD93lTej3h+sNGntJPvWWHYKcvBEWbKGHErQ2CB2yAy
KPp1Mcyzvcu8dCpit2N0/JcRbVoIfkzQhqQkdXPCtXek/veDFmFWxoncLcbV3QhL
lW9meZvdA8+PkFYkWilC7ceXeL9+BsIL5cvCGqz14Rsw2poZtoso+3YltKKEFJO/
35YbiBnOOGZ54izg2lsz1anBxqeGS2yaNmF9j88HmaL1UWviMNWQeL4+/UToo++P
HOybxXjognaVHqrc9vmdit9XCDqS+dvnvFty/wFs+lhhg6565XkpmDeLVOivSVrf
bJACb3NHExZCMb8iXZGEETqhJRc2RDXIPFWMpUFzwwX6SROd37OO8sXe6wvRdRLj
KgoEACbbIN+yr7ctb86loClR7cNm0ChoAYBzNl32RBGjyjr1xcPtt0WwPwiFdKuZ
oartlYj432qkj5/Q5DG7BDU2Jd5jV25EHuri9rBPQbn/vpRpQRJEdubrXeugafev
2wuE8g90rrZr8Y9XvIUPCUHeWxjvx+9IV34/ed/xceVmdGssWjcZc7gezKYSUL6v
MuptV7MvFueTEex6Ul8aDMIGLlnytbLhApV+2Yspte1VH1oGWR6qrMrCBrS8UuWJ
k5O77S83tqnDzzL39Xm1YQenJd9ggb1wPEPl/ppng60Oqcv8UnBuRXH7RIrgcXIh
e+1aciqMxx2wO52j9CGEeeoxvw/GhGynTIWDqTXvkVDvq0PH1UJIMDjBOvuTGJL8
DEIe8tGiIkIwbsArINL/CUFHH429eih3vh0coLiE+R40QKMStkqUW8RqfffwPWWk
gTIFr+6yuopUvlMN1gVJKKhKg3+OAFppCXTOwY+r/DSW8So6DliydWemKB4EUqUu
416oHVl8wmtKQAd0v5PFbZfh4pP+aPqyN/cG0swfAnBywTk0ip2Tt8KDlLZnl3Hn
UWa/KRtJfkY+GzSikmaoHr+5uGVt0Dk4CV2upA/BFlfyQmkbDgxTojrA2E28dnFv
SXCHcAlGsY2/vGvRQBxJZOEIZ54/ZTayJ9+JPjw/kdoFSjrhHn9C8J3yjRQzH+jn
JeCcQTTChD+uA3x1PR5IxxZMDLq0FUXeWJnEMgZKCNKrcvjOqhkdnodKp4HoVDQ7
I8HijSiOSaEaHl1CJkDzZVIKyIi+ElVvnRDffMwbKCH39ObeVDtpljiDqJ1f22F5
Aa9tC9A0pDxyFgCSgB+CN2kMBvM/CLL2qJe259EYx9tntr5hCvhhCnWauPkzL6S9
qJZjThxScdu9CcoXt/zaYZMjWbkXFKcTE7p4uF8DbpE54O34Xn1VyqsBvULhS3Zr
GY5qJC6QVt0YXW0lETfWRIxDFeEyODXRu/8svbrKxuU73wowipDLG58DUXTj4NX+
b7UgovLABlbxVCWvuRHsgYyBjV8r5dLkWFPVVWezcrZ7d3MfUng+hhunxfNDOtFv
7xhJKZtw6gk1j6Czi+7ZVWGnbFhmqz22VTnGWoWSk/cYX9MoYxLNSm5rkwBRDams
ZDiQpkhjcQgTkCjgSsfmZqoPEQdtmsS021ItfSN0jqNK4DbiazUTU+Phr/jwmwyj
SldhwhdCyIhuV842oiGZFQE6UMMZtAf+951hrUYvxL71EBpPfD8yPZ4tFj312ohn
5LkJ7i3vezH/3BFV7qlr8ah52aSlR6gFahmUiIvsInnI6BHGMqV9Z2w6sGo3wWXx
tKBTboRMtcIrnXjjdFZsWszDEEIGSiYeZEQ0c4x1EteEnJlrZyQ/kZNP21okkZV6
gAI82aCzvNXFiwxOZfHWivzar+onMd+sGe/EBsFgznBEYRjfAPDZeSSoUzdqUkX6
XmLRjPxEAjlMlm4TtJ+oYiPRUU7XNvUNosWgYhNgcihv4GsXQcikASq1CHCBXcrT
WOIwaWlllXwrDZJVLoYaQqRcM4q0ClpOF/LUuY8yLW053GyohgrFJU1QFbCSXrp9
JmEhY7aapUArjcxyzzir340GpJJObK306xuy4/FQhMdu/kd19SV2C1ULli3ck6Hg
H/n2Q4j340LvapXoLdvBhpqgNWOBB2IvEbgVk+tv3Yfp+LSxQ9nBD7QY+GqoqgnQ
vQ1+qNrASpQJ1h6b16gwdCcEz+nzQYu7Jxn06lmVJyELczYB6dH3Iv8mZyDFrz9C
qtjEYdAj6ZBMgOd56B3RgimTEJfyvS63XqlH23+jALANqRYL8MqjSZFnQoUGUZH9
MuTiwfcUv3114eUBff/5BZEaZbea3V3tWj1rsggwyDCZjTdtK2PdmbkEk8KWW07L
7mKqgoMw2c9HL63BtU+khWE1sFclYmaxaBdunXaL4+Gpd3WKMGBkrYyKh/Yo2D7b
24IF7UdTiFjmmGS3/ViPYfGiLnLxNnh0R2c8RaFLuBg/txS1I4JVKimAZ3/9gyzg
aUqMKRYnFF8MSmOzhrINLi1bItxdOVGLUVddgpagQOUvOW5Akq7lpZFLbL3fQ2tc
HjWI+czkDNun4iIVaCvAX0wmDpiBIUMRuzPqbGmGoorkxuFZIqQvVgW4HmtSuC3G
Kad1j5WWIkpr3Ld3/mIuU7JS2QHzjWCdoKmaqMqMYGDNoTvux48NVG87eHWGFs3n
r27EjhuB7t33NJcJitg2uWnEse4gkLy+RMPHB8l9HKVLJV1inr033pHgJDZDdjwY
BNiWjbAM2r358uqzvEzCp7MznB2+PCaJd/oKCN2Rhvh6GpvhC9b7walzugFyym/M
+NS8y4IBpSlN3eYhAYHOfajcQjCLQe8Xy7qKFnUpIZX3snbfyUFHf7sbxN7UBtZa
e0cdoHrQFOnq96eZ3B58eXu3FYvLdfbfH+D9AFnT+B/UloIpy7NG11OZn2Gva5yI
13kUpFn7AHSuUHIPE8laUavZQDnfdaRAxWVY/K/jCotB+hlTscNXIgFI2UfUojX9
70vrHg3zvKaZ+hdpNsEb5U3U7R58KoO9qIStHVERl00U2W1GElCDQa+fbUzyVOKj
nlLWQNiV+EhbZ2sIoBOwhGX688mR4dwjdR2caVDqm8cUTGerUwowL0eCdr7GEENq
D34bDtKhzFFWNLFwTih1tncGB+8K362vxDbIITZhyiaABexvOXYNvhFNfo66ziaI
8n2u3fsoF2C4XnL0JIbgMptgw4az8RavYEaAmBL92Tc7hNM6QIJwQFSXaLMb73UN
VuKWPLAJI0414+a7beEPc6rNe2DzSKneRP0/IvYzd6/s67k10RkkCGr04bnfhfco
kLSVK2CvJ94ZyPYh4X0YgaT4R8L8RNns/Ht4/bnfn23oF2TXqhYQW4auoZ5PxO/1
ufvFsdKmOxTgVHgzVXSe50qPhKvtsibNzD8DbROtyjQr3Vb7KGX6H/QNUA7wkCA4
0WM1XO674HPPd/sjCD7kXk/C0jkRqvT318OqqGAuA1EHdf3LSi0U5zrXSaZDDV7O
1wO+aD/CySz1HSP2pP5q2IGN4sEdeCjUW9zYelx53rC5SAtPHi54gMY1CLNp86mS
uX8BDuoFVEh9qxVu2hC7W4aC6eiXEL1V9Q4thAMlFIXsNitv4zqr8q449xPd5xa6
eJdhxB/ggsEcP3mphF4tPQEBmooooz2h9SJHWlKJHnM7zFhrnPHojgFd6Tak+U0j
xUdWg+9xYI3f49uuIrBIyasdWWh8sR2hgYAmdH70ubQqAM6o70+tXjRQ4R06Xmq5
ImVe9Jlcaq3n0s9zVMqy/d78dBf5Vcp458Y4WgaJ42pUKHBKup/hdBroO2xKdM/2
Y0j7bOHdwYueNr9VFU7XzS4Y04DmIAmSVgmi0/RBWfxnSozO1vdnircWe5W4z7eV
JkMVijQCx01KdvkWo7XiiukKzz9JQn7BgO65Ef6W14iL1JBsfjietR8I8AODqloQ
zFzF1BNZ+CxGzQlBknvNEmnVD2ZbteIPAakZOZcxidw10nlSc1zTEvxePsvZimQl
OTdy/CiM7+kNJZaj2TJUB/mLUSa8sA5XUsTa4JVwJMcqQ/5PcT5Sh4ancW/gzZME
Z0O7gzxq3G5BAcMaQNm6CW/vqRzN1h8XBbP2FY1Dqtgm4i9QX+3FUrLjEEhFPDgI
leCy2CejLG2YskS5bcjTKyA4ZjhKvJ3O+7ptB1NzrE6mOccrMU9j7nDbpEsFn8DX
/qJGt1hfiEUiqDAwip2pdAXFOC3T37+MoYLYD/mEi51fIKdyM1C3aFmtDbKl02VR
PoTSmKl02fqsfho8hSQeT5/2fGMC2NbNpwYrP4HPKlsOtoTUakhAfnztq8urBdgY
uyyLQ+Kz4j/+k/AtEDQZ1lVmoZAaE1pNBQOyKTj1EO+giAEOlrZs2YJ1w6INDZs9
i/UoSCwEZhV37jmKalczWK4Kg5mrIxHJ9UVUVFapnUwvcW1jrH77x7ed/ymdgIcp
Wp6Br6s0ETqBMK9rnclPl7yx+8qnXQje1AiSB0S6UnefpQ01pfEAvJxmcGMexH86
9jAMpUMyDUntEI1HsRLJYHGRrzm9n/djOdAdRugTKa/HO86etzyAWjFzyXNcSANt
xno0gxDPqBQOzm+YV2VaEqT9APHisAkLCQGl/ZDKJ+7gQGEA+jSbhVRHGkn0J5Ly
hBjRl8PFBZARXebLfMREwPbgLNGeXJClL592Ce5VGTTNIAAfCdx1j9SawFamJmQ0
Jxgyp1tMhESjJjEIzXHFoS5RVTfu4S4dFeZexaQXdChYZ6dNyqpHdu+vNmqMxprC
YxiI77lCADD0bVwRDZG6axjUwxwCwZUAUucsgatnmc6NAIDPcuS4mHpBIb6piWuc
US8kiRMbLVbQclUpAm1B5o4B554YmYReaads+oDxRdQMjQgcgF4I4B92UNvuY1tg
yr1tBiq0e6g212sgvDxLrGKj9WbMzdnpNs3Wka7A1oF+Us/vHKd91NckwfgbBSp+
5F0z3HxNH9C6nXsSqMBWVpEHO1Bhaylb2MX7oQvZ0JQYBuV/LEcXTUZSb1baoOzW
bwbU6sT8B04O41O/mJcNFymI8BG2jgX3fnDGTbfaFwtoNTmxbOjQ1v2bRYdYsas+
/2t4drbUJhsLE4D87SRL75NFrBO1tMsVl72uCHeSAOKgc0DmaLR/hV/LUc6hNwTk
PmoFfP2ID4C1lPovBvqVR3HKziPXq75f5QrQxM2kwjBlurufxwaEqahkssJAgDwx
eSvQ1vYtcEk84p1dB91DW9lnRVYihTnqf0h2B6WE9l+qUqLGasq3bD5qZ0xqdPZS
n9/uaC5O9dw+Q8s9+WgpkQedCNH2NlN1tP+ztUD+36tPVJtbFfcd0f7YAGQnh67D
xE2rGTOHZ6X/cyGuS6oTSHQcZn/QLLfIocsiQVgvI0Bzivqgw8HixVjKOJyaC1FD
NhCuKWBRGVD9S7Yi1zl27HwOlhvJQct1HNXlNgAHgZWQ7etiEyUJ6KD4rFEizwnN
9tVz3ltMcitq3rMln0Jt01P9S/+P2NpsmC1ZlOww8BdwRhMQVr+Lz96k6+OxJZTR
vo2GcrExjSelfqWDaGng/oLeVOCmO+lr1caE8p7MoaAv7PhlUza98zntlw3b+SyW
GJBfnyMQYEZARAXPv3Ru9e9MoYcSaRupdnnyeboVWm05Kfm91OqfCsCke10TNgCn
cT9zo3u+Xe9mwZSzrH6A9nT+BubvUIRz/meN/eq2HYnrjsChcmt6fSe4BaTGN7vH
6XqWP8XpbWXE5nyrrvHEdQmjFDHwFMQZ9KcHOuB/rZlqV+zfDK9Q7nDMWR1qFG0Y
4PcfU3odik5uFbWvHyuUuaSq0rBZmnYd4xWb9Sgsg9F+hOk4QOfVLeYJsoEWFgp2
LwVLVLpZgFS1GByR7qR1C1+FIXS7aGLYOc8TvqbvvbBJPvHsgdx5krb5PWBVmro7
lMzFVSN+RpiLgYfBsf+5Q5x+2icsfykkPBjKOq5EhhhlpM6d83RGTSMBRoLnNGOh
GSY28GzFrH+eFIY3mjJ+yvwlMg+vqYD1JGcFXxSnh+fmrmVho/dmRye938Ojc+e3
4zzbebQDs4Gqiw6kto4yR6qfbgTHMeP9X0J3K4qf89UVZ/TofW63d6XFnG05XDa2
uIij7mMEtxLqCVRLs7x8ImWzIybTmkr0xscmqSCx0yXjXZDRJCmtF5iRO2CvMUyt
Lh+JjV5C3BKLw8bZXFumI6se3EE8m5r1pPtQZoLonlf7qJ8opNYb2DWN9EJqE5lj
aaxvOgFX3pvwSaiWJrAk2+98+eC2sJ/5ZmEdeKmChEr1EZr64M/SwBFbQEt+rC+R
z+ovqrQt9Em8AAalrIUanye2A4gD1KoUT+S2kVaStLSJO/TmQnIIK/8MpPqUW8+E
EqRKjzR4XZXn7fpu+XNCUwYRoyDituK3FoTnp8/mdeF2olpWqVHKYN1ULZZkVKAc
8LMhkKoZwVqycHZMC/BBqmK6KTyyaEIDhxc//3V9M/DwrZxEoXDGV1/2AEY6edPV
WsF96EQhYeoI5cPeRrk85Qj5biVYItQ9h1O7UGMhYYiT1ozvr1nPWEU3knsV5B4z
9jpIv4IvxpNWVnjUHXJJvKMNESip0a65vOuuWPe06yT5wmgPOMwVWeqvll0h1VRr
nPavbnT5s1g9y37egcU5nI4HqUigZXdrhYHU/EGDYchvP+Qe4mKy+pNNbw5OB8SR
KZTbSqe47xX+C92VnPahGfy0E+XHM+7dA82L1Y4J+14AuephQI8ffWI6dL8B+759
vcdrY3HT4rdtwVwjMFF3jdxNBHrP56bd/O6i7H71ps27EIpl/OR83m89VIk0uvcs
BRxRo/HcrkHodm8loPux77MRJj3pgHbEOGEbhAIXdvjw/yl7ZrIRDNTjOvai8kt+
JmkCaBvNOETzuuEHTPE36DekZ0DCf6p01A4lHwo4moTyHzOd2tSTltlFfjgKxCI9
OuozPsivZBJP6MMK+bE8Nsoiy7pEfTUUFaWuycBgXvCWzK7Az0a1O2IZespvUerU
bcfiZKH6lWNrDCQXS1oUj7u/eu4HR/yuqVpMgdjpaE0g5CASt6teaAN9NB3mfp9/
sxG9NVmoEPFHRtaIduDgptoTzhWHDmSSYPt3BQ00r5psk78mPjEqNwoJozPo4jkW
k9O15LUvhOvGbw48kn+BhDOehujgkXBptKbf6hV09g7LTu1kyL6ILzmxmANq4NEn
4llipFgiMvX4qUNZ6yClPZPyY0n3oI8OmRy3t4ZO1DDRtB1umBdknuBPv7ePzg9C
RwlFfhJj+xpiQpXik/YQoyVqZVSL8vzA3Wq5Wb91XUSxHu5cVo5DMuRv2QpSDKtz
JtYWpPYRqdWCJsBJlGy27FnU8u+f0/kTa23g3ZmFK0A3Sl0RfDkHzi6/0x82aLxt
Sb0JvchXzMxL+SQZLHRjC+I1WHls8LLAckgZqNc7nR/KO1TPPHW6G8bKQpVBm+yH
iiyqvLeawTURAUaQck4+EYYfTDfsi1rISdo2Aot5Q/vR+9yhaQLNnYOOH4XQ4Bib
pST0O0IBG40xXwmt/ddz01mODyXKBCpol6EDfQjHYVNGMSqf/iI2HwHSJiCQ9u91
jIdi6wanRWrmtqA4Fxwhywk2+t9GggPIM7ylWZCbaAt4csCnLN4MFBGWc/pdIR5I
S1sXoJCqKoQ4yxp3ZYR7kYEfA7gT6m2bEKJgWd7UBHHtiP44SeQMdNnYZkAw/prj
li2lQBrMo2QrwuoAGmE3vI0cMU8NMeOvxfmpx7VmdwaLLVVuKPHuxGZAEOQqmjZj
oxn5dbRq3N32BaX/wlBvBWSnM67iysLR2tSbw9/7p+XC5kBnzFcMOhr0efkVBNgQ
wQFfr86vddgXvrvFG3U6g2ZkQaZwIe8pDz3niyQlZ4DPsPGW9iwz/EbHMcvz2+f7
9a63hLmS7o5O2DC8eIYs9TKIfhJTeQc0QkZ4Dh+OZT3NMs/5gbmGbGDSgcJrHLd9
6/xZxqwmPNAwIjvydIHiIk9qxlU6/KEQO5aJqP3J8PxZxnfKFGipJ499yoQq4U+c
0GtZejn5K8d6buVltGaBKDH2dA0XgPyjntHcXeEUXKkC3qjW4VA5KyZkYYRkENG6
hP+qmsuipmhQ1o1betMvqX+1tgDwtaEyr0fNUrpldlJ8vQOy8wU2fX/vaeHLPjav
HeYL4aL2l3XUS5DILB8cIcJyFAKxnQ4zkDSjt4ZvmcJT70jbz/NFxK3xZU3izn+Z
HDx+JbK3nQuYdRbDMt2BCydN3E1ns1n22xRx64Hv11LgQ9sRS+xt0Wf8n629O7FV
VBFj45H6wrFMKDz1jmdsYakPRV7XhfglfDfdnoH4X8SOb9k1bfPPLnfdEIUqQm9s
n62C3TKTYpDsXxmORVlPxHLRRk06iC1or3xbwWd2HV1WdM2FPWbjSOlWNXbXk84D
3Nun6LMVG+pR4zeEF9Yor3qy7+iWfiYDufIiDWXp0c6pLkgqvOCE1Se1Gs4eWSOf
JSUGYWFtb8UGiwcg2QcoorNwRK2MTn3BN5mWNVdUF4nekXL9+dKxPHWfXqTUJtUV
xDxTM+i8m8lD8sMn0LwcBd72cmaZH0WtdD3iMNh1tLzt6xBFLpzF2owfU6PzaY6r
rZMEnSrONQ9+ciomiAk7VwKsyW+ZzsIjb9521vQt8EkBN0tE6D09M0KdIyX1Cq/F
6VjqCR4QZQLccIroVKi++ck0H1suRP1ndm4ZlGMdT4UmtIxXA6yOc4zGZBY0bIov
Wjq0w7H1ZX4hqMdP0bCl7LTWqcPAqC2FgagQrBzs58r0SSu6+7SqaEhFZZmFc8v5
KTQXEAPahPR4/F08O+MoZL1PnFn5l833OXG+ZcGMgA0z9MZh6Je5mdF+LasD/X89
/TF6+sTPwTySX8etB2dJjyofghhJavGfeNkQktOMsUBPIgETLMppWDCyiCwZjL1I
+NxrWvE4xjWeRosOMRghqK21/dXgb6cxuA0kIXTlc1ZllL6XMtc71uM562say5nj
mRE2DXHrAioRrFmaZDdKLp0Z9blyuGFU+egX3JGwul5Mqr2GFxGJ89RMrFOAvEB/
MtA+lzXxsyMEPKcw9LZ9IyjvLsqsqJgQzgWKEJPBi0jJO5FvJHB2OXEgU3KrQ6RI
qiZK/mkOmEPBoVx/xtQqOO6OWpqFKFoR3d+xA4iWjRFEm6WeOit38GmzgnvT0agp
432HHi1RUGCS6XE+gTloJZLUnJG0YuJAcylpOIS7usQM/Q7Be9yXqBghR4kFU74E
4uXKjA4xqN6JT780W/EuWv0DQ+PQxTr8szN81KBwv1LYWqpJQLUh+SMr1XLbzGQN
xjmjAcTQj5gpFGBJlYMnEl9Z4n6WfCfKQp58ePYdWSbu3GLQUyjLmjrMRY4oxBjE
JZjlrmrHaGpxW+wOn8Dn+fmCu01Byz8Gp/tIeMQmrsFy2LtfiRGUjt15jlHkm+eK
XHiRPYgdOUmvWQ8QRPXrjwGLxtFwqDAFi9UCXQTKZdpjPIgIN2vPmYYViOxDBXxi
NT3V5+nhl5MmgO9/CXLgnICJkidfy0kU9oTWPdin46fsswuB8JRHhU7a5yQ//4nc
HaxxYSj1nO8VHECJMeiWR4WFdqU8a7MqLXLYBVEW1EcK0E/+1fK0j8DnAf/uiUmD
/ZpDCYD8PbPrtUiGu116PeuFbP4kLm9+Bqkl9lF/dadvq8nkF4NNo9G2nRqOaNy1
yhafGMaZ7YQpeXUKpik251YG1e/5q9OMx9+ssVFBVzPyHvk3VkCCD9qn/mBx3Qgq
F4eOhkVjozlL+lfiNMk7Nc/u+JGFDRWWdcb9ZhrzOxi1L9up2m30vxT/xSVSLGQd
BEOFIHb6KfLkRYwU7PYOkp79lYX002xuvuPr/RHV2/Lk7rWVGrXh8eaEJWjYeR44
GEIEhx4E9fxTXkCtPdHwlsbPmv82TL9M6XiqpMUgcGrLhMIuL0NVZbcap60xmsb7
NeGvPJopuW4UFhwBIzckGSgo6xKFM6yhqTQqmS0emRQLlg544z5Wy7QjcpbucYoX
XsukHdqtiFGm0ofM7E7bv6Zq3zbk0tAHVSHZDd5i3Nd1zzdU98B1HOna8lqxDe3A
Vxmbdb2jTYFxANUf7p8pDIynEzgYK2tn+Ci8TmyER5fKuq4sFt4gfF3hZ1DYthdo
F9zdJSTq5scTZmBPZxDplBWxY90fvVACVBP9fJ4e944T6vDW0H1EvvxQfls++91C
qW5V2Msi5IKbp35UQKaooZMVUYwiF/32ZefMP+ie9MLkAi0PBBMch+gpG6SCTRmV
pcgzHEA/g0Fqp4q4Q2Xfkp3Ua50vocXm9HjpjbArhBzBP+a5scXyh5fP2PJIri/g
wvUxyGmHwJs6A8Cfu7PhGNQPZ2WqmxsgtLDP1gQ9aYLaRtom/XlydiTR8sqHrTFt
3V1HYKr3hgyb2z7RXL6HTgnystoZ3QiFHviIji+LKZAFrTbw6QCd/RAKVeza3EiQ
VQBClTdsB4rhsYfYfALCMVirCRKTHDs9Ufei/BhoPc1u7RE/tuPEOsgX+tYDyBkp
QpZR8q+E0rXEF/oabUsesT1hY9mUvMGaOvI4sbxOUsUfmaWX5U+w12T6SKpyhi5m
v6Reh0CLIYmkeKTWt3qTz2OCN4w6YfoU1mCZqKK3DKJWJPEKpKXGHIOsFbUvXIZu
MPZa33CtNSg1Oqvc1OVnJNsqhm6FQo8T3prfoaiyjAlax/eu+EBR9aJdkBuJWmuL
51goIDgd7DaF3fzDd3isK/HFgd52X9Oob/dMoWoBMj/LB23IOFvSGf8rmGo3JvkH
AKjvep1krdSmj6p2A+QozeN+L46YivDJ7RD1sbh2YgUjIQAfVNG7yBr0FzHkBBMo
j3Z2+vwXIYxu8zlT7SNr1jVH1jtpJkinYZzt0CD5XzDV1dHZ2Kwre5JieNcv4tpN
yV9z7wJoUM0EmFfrNsWJCzckp1ppjjoYj6/dIYiw8NCv0SZYLzo99CHsDTUaSkGo
3eA2gV077sQnSm3v+EV1oikO3Z9Iy/Swa5KxQdKlY7eadxR/EZ72lzjk6hU3vwE3
ymjZQfEbPdhAHpW+mvdnWWJ8koweoOvKxGMRY22w99JcQUAXvaZpXb9K43VYT4jY
1YP9vMreqODSLNjUBgR5S0iipzMjE8Sl2fSvPAb13CBoHueCJqcy59sjT8MCt3Qn
TwUKire9Y3/ldm/IGpVzi2qFcVCUOrUEduyX9wEseSYm8dNH23W9FggPlUUOLszN
8ZRTAzhOQaiSU5Iir4wkRfpPtsAI+m8PlTNtKrJFT+CMpcxFouOyhOXGkg5Ct/Es
VZN3t8VWfzCS+9+rJkFQzOTcjCuWiO2i0CTxaw6nLlPrqUPFbzRsTCousa33Zhfg
N9bCrMB1SOLcSppGGR+RHK/LPZbWdtgD1NvhaljZl/Si/b6UkkTlig2RgOvCQKJd
gGUtwqUp25CbYP+I5SGgg2xyz8mup7bNL2Idv5A1Q26eDd250kC+BDF41+2U+gzB
dj0Q0uoJnCtQBwZPakBdv/c87QcJmLphr9exk+cKW0Yta666j9AiQ3FHhM1ul+Pp
sDVgNS/7DiKBS2+EJu6qlGF0Bxc+n3bX04U84BUCIqCloKa8gzUhJhRFQRrWhhb+
CLcA5A07Ft9SNNhypPe/S6nIocv08x79GDd4MnGIvtOO/QiGIdoipAR81zzUx/5m
Wk2HqOd8plgp84n6tgWU/IqxyCqrj8ZI25oYomdQ2TtGyynXI7TzfXQkLvyLOc27
IvOrcYXm0GBl28ATi8UNqmQkdyQrdYX8khAXF7CjBJqEOYC8OYtLkYwJMxKyb4cP
97ndThW/vQbrOAGckIzsFBZkrzoVxcl/h0K66Ddkh4jVwsGvFwo2TrhYW10v+ssQ
q8B7S7MTs2AX+SpfEgewyObpzXd5kFAunHspwDMHqMug49d4vsI0M0b/WCquEW0J
PveLMiDXYWjZbnoZWz4KRxmvOfQWwLAMWx+cpdq1K/OEVsuTqPIukx5Qx5GEhnf6
rtNY7Zzt9BMt2nklHAIUCoxVDS1A4VRsa3Xl8RbGFnLpuTVsCixBRS5aAQfobP7i
HwnVPc4ChRk7ZVvnG/ELOf7CQfEE+5oyBMf4oskjGQ66pSU9TxbPoMP4ds251z5h
t6+borjGHL7D52FzvUXsn/XD9Gqx9UISQhkOHpx9M1dBu9I8ojn2xDATGuYc7HMQ
+UxA1+r7hhg7I6SjVsZTEcn+B42Ao+srYP35u9Rq8aSGkvf2cCVcZUoRP0CY4Pj/
UGdMlWfLhsedPE0EuA8+GXLiT02p8LxD2c8BijDRZ3/M2NMJlDmBIbeyT0bQ2Vn9
x/Yrm88Vk83LaLG41uJte1VTC+4bH6hN2bH9Uma/225Utyqyqhh88ssXEo5f0Azm
GnuBJNXw3S2qiCLtDXzDT+eoeJC6LOmvMl2Y6mOrr2Ft6uv7441N9IAay0UZcnG3
dCzZItd9vBGp3ps3iqyyAchNMlBJR4pdxaCyCt89/B8M1nn77pQlLGoC5/ukR2f0
miD6wEhipck0KFUn1u0uPRsiogy7F7fJ0l2LsDGTST0VAQVXi+lnjx8lT0g459rq
uS3+8EC8pxa/nRfqwLk9gWktjvglnRdElaYS87NnYn9yeEBuxgq/J7EZXO382ecJ
so9DgcnjCXaFNsSC2JNdoZr2knPAGwspgNjkUAIjriL0L/kO4nvaG3BALz//flBT
ezms+dx9jwOlQghEW8+paTdy95sGvScyRC25hNeXX2/L034PvJr44ouZatH9o1H1
jkxfSXeCSfY1FPomQGz5JBszBLa0A63e2RXC+G1zSZJ6th6JMxQkD5N19drVXX4U
DeblDJe1qdD8kIJ6hsswqNyIyoCjuPiYIiE0mFlHz0bCYMbGkzOrEtYUaMyVrytq
p/l+77Pi7hEAUZYejaiotPEMWWlHB1ZVgEeAzef3hl+LjBwPtUYxCZM6JFzN0lI2
v+u3OZSJBXh2uW6LVhXlYOFmfJmfUxKjo2pQIjg9dCLbdz8OmRq18pGbfCoWwNVu
xUp+Js8Nykdb/rBM2c0YFe5qiX1rH2sqPk5lEpwSCAuYULRRwYK0M0BhuvSJcI69
yPOkaPi3iLosDegvs1Dt4ySm/Pjha5G+3U0s8Y73nzSCKg89fERqCz7QdNd1NqIR
37L9bqcRRtN5KrM4I6wFNd8IRT64Z+xK8IrJNMIjeggC5dIdJbZ/o3uE3GPhUzIz
tEP/O+velAYeiHMWxXuXOg83fSfQYFzY9HJayo2XjVfZtSB+pFD/Kv5U/Whcd8jr
VOCCZQFRuXvDlgyK8r2oJ8lEc8JTKG1gubcms7kDBpuwwpCg56+oVDzDlc5mnqkv
0z8K8OJNLATjQr3ZxFjOIeloWMzApcuoSn1mpBl1H8wx3tvHPreRky0+XlAEmCCl
OXMPpC7tCT79Yo9sIkl+CB/jYBKhojh/hv6fyvq2LIk//oPIdbyNl0n19G8q5jhm
WEgljknjxbn9cTguz/b20m7geEtq5sb9AGsB7+SJwdziL9G2QKZ8g3zikqECsOeR
smkjPBUR/jpH6LsRKARWMupMa4hla3pF4slw0SaFE1YReuOlMqBFtZCG2FL/37SQ
teQuV3QV8Op8I0Ypz9y/yn2ONOjVf7Qywvdaq6LmLV5HLsBa37RQfGM/+Ir6Ik5K
kQH0hY294Mgc77BF95BIQ/mr0ab3Va467SaOcT20uvSle29CTVPnh1poP+hPhC2m
73yINPGom1YUCV8IZ4qppsr2YpyxmIbdL8Uh1dKdpWOnecADhTsfptpvltBFlfog
MZwsqHllyjI4HlyIzuqMNanxekZ4/wxDrFTaf4nOSqMxXRPc0uPjWo45YK11WS+4
N5gxlrhLc5yEVSufInbi5F2oQW/TD+4H7YlYA19I0eRcNkyf4giei7PG9mVm+ybn
YPBMBNXIWFLSU06D1v8C8dej+Vv8QHTGjgY2ZWAy79c7N/BdpWjWTejY4aNfWgRm
wk9LlBVnUoZqrz8WDhDXvVRam5yvXHRB58m2UmUiqXiFhwOL1vMYoxAnzNEWFAnW
/BQLsMMy7V7yfDHAwF/fleJCCIn+smfJ4cKPD5pLn+ET+E/avahjKmsRJde/yiHm
hjiE/y2XODnQv8ACNiSJjsdYqljLQNQi9jfyjXgLci7X1u2QYavnUQxEfEJAezpf
mpOysOT+eOM48bI7uzaFm+I3ComItSzelTnqKs6jlAm8V2E3e4lrz3EgbfKrhXI2
7aRYvYstoKComuHhKuAIb2UNe/yLezWcVTlZEbpsbYXV99pVZekQzDmp5FN2o1y2
OejXlJqdJbTn+8jEhRdpT2AHJHEFS4N1L3joknouJKKgmiLIspA9aVOOaMqlX862
NI68CqE7d5fBd2LnaFImFGa/AZ6aVGMP2h/u1lH5u44Uh8B/Z8l6rKGT/qn5d45e
rzqj3wL8ippRm81ocFALyPFiuvoJuFGIfXqMYjcMerLPQrwBnLynzz8CAAEtwT8w
DZIkZBAHgWXnyn9kLg+XhZW40MVC5Rh/ok0JyohYq9HXhGYxdE0Ggdbe/lBkhwWq
OSA9JhJPdXBAFy2xyiYbpyNUU0AoWkvQc2/a1TJpZH2XrP4MQ9UXPJpRED0OfZa+
oEpSzWLIbvS4lhP7TujKNe91RU1VZG33A8H26MCe9scXQkBSz4YgVjTB9cdv59+J
J9X/+PvimWEDNatgKUNaomSyobuRrm7LilVKXnBzsm9hUxsDPMbNWlm7ljL5FsGz
jwj1bVU+Svs3dVlLjYAcFE7HnzO0Dvtysw7VA+R9kDcNSLX4//Ids3fLzDgRvMPy
KhQF1qLXBdDnUg+urIJcxMS9A8jd/7+ryfz2FgtGP2oSJLsQa39sF2DVLEPnWL8F
dtwDUFRTvOXIS8yWCHib1SJCi1jIk4XY0sLHSEnp4HODmVmCqUCXPlEjrxTyimc2
v5AWyt+VqGFLvznAghjabnakVOu2HicvChylerSpimdDZtQQaMzz0saiXrYJjI5u
q1pGO0crGbdLNBG0f7QNSe6Sj72JtTTxIN2OaDRLol5IQvP3a7oVj37Gg/r/imzG
RNRoP3owH1EyiSHWFs4TPfSXerq5waKedNWyZv/cns5KKA2RY/txuDRgjzQOC6fD
VtucXCc2zvgfILOXQa8L7hMYDU6z+MuFM5tBRp3Y4G6mTUDL3MjlfXtlqRG2ppjF
2iFPFhfBVnMIGUpA/PepwgT5RQzH03yWTmkP1Qt+ru4P4LN3ZECikrYgK+0qocGU
u48OutssrKqYkmS1GJAZlngeIgU8zsWGmtpx1t0SO7zz/BWxBDOpl3A5doBM4jw1
BAHFzfvjSVi2tweRQ7QgdwyIQrB6NQoKx7z6/5XTdLLOZAi8XOMyAfSo0ieQSlKL
oT+6sAETnydw6uZDNexPSGeHCLvTnRU/uHEIsLZsXfAcrGjR8qOnfUJFZ2An+RKK
RtZms8Ey8VFJ7rU6RwHc+QkT8cZ7gu1G8y66txnYjeaTXetx27PtITo8Gol8xOgK
QrhOj6EmpZbnjlkf9E/AKtYA/BoMZxk8lHGsgrb0eiXi7Wf4BAQHOdDppydkOsVy
dIyW7Kmib0QUvj/TmEH79ya3rtGvzWl2mNOgFZ4L3AfT5lngGAJoGbWEN1CvE48M
PrHjsmjtH0LL/lmCkf7Jb4oCc6Jx/jr3k0KaF4ADYf7++Jl+LObWtkjIPvZj3J1M
sqY3ZS2xv0HrxRys0R40nPy1iSYPcs8cNetpLqU5iGqiH+ScB8yoqFyZaTVKa/F+
bOgspjuLirVH2YkEznQngjzU9HXnAM+VerCKZH+eDRj+D3O+t6VZS6uX3gx94MF+
PQvIS+rQj4p8lS3DWQuFCM34i2ufpVMXSJhMxy64e0qva/V6Tb3o0r7MKdBrMs4i
Wld27INIGedLIJb001ued3J+uvvlssIEdSGUKG4ePzFAYxmUG5BfKSYwNomrI5q3
ngfOWRRHrkEfmuPBXyZIjgsngoBRW2s4QXcsNkMa/9DSMlcfaAVbfjNnbBPdT2NB
XupnLrs1GtWPxyBBmHZlF3mDzbk2k3P8KHZu7+8MzRchr6U1RoFT8Yx6w8G/vdPW
1/V+mathXQcaQm2cNtklEbwYAZzRIn5ms3ZyOFG0Y2C3IGOIb68ipdlQaI/te3Sn
zAuBOIG+WhHmiQdQ1EnyeV8NqNPNBmQzpOcDUv67ErvO9ZajTMTD6kdPh7EyrgSs
UG+SBNE7tW42qyDGR+uFP6P++9gxcEW/0P7Etr1NGZALkHvRkVKtO4ey6dnx1+pG
OykaaXYZuc1jM7kYyGBuqY8FLcGJppJCIIayT/xtYMl1oN2rthQQkd+RyLpgIi5r
hlrAAshklmG+8ZnzOkEMuY/QVHKgJ3k6NvqSD7xn9V1ocSsvKJS/V+3o9Q2M3shy
aNEokp0TJ4sho49Mb/NzjsZBn5eFbvChJ3i2RvMtcDvf2FBIov7VfBotU5UbdR5F
b2PIAC4R/r6VfaCoEt2nXcoU5vuQe/6Gq6fCExGubeOoox4TOAvO1Gq1JJSqoAUB
hXGYvAWJuBkSm5JyLyhzhdeBBxT/INynHLGLbdFtrpzFuv5axZT997umnI69d3w3
gAlYjkUGexTbfXB4Qp5yvaEk8ESplQ8iFupTuxbcLKrtpE94NBhGUH5S1lLWJH2A
tFFM+ISeiQYoSBAFfMMzftLLnws4FkCj1n6BxP3mBKoAkJBnlG5zXXZhJBc89BA2
ByG9tnz6MBrNltXp5B5WnQ243tHiKx1NZeNRxh93LRImfMWdtICYbKiRI04GhhNp
cIdJ3b5mvY8uCC5Xt6XFQaJa4Zmd+gvJ8+1WOXQMmUcYJHqglLrpMfTjbRdSXINu
PZ/59jZ6+aXAZa4FQ0bOdHpvrq9YPSraOpNoWovhWRIFeWQb9oJ+f9qEWgasFBL3
Pd0bdRuvWvLrtYHY6R+loOXctV5lSc8dxcgV93AswFyTcYS1B0jCs0ohm/k4FZUQ
3MWkkT3CL5N609my9M79kjpLcJ5lxZq7r8anwPJ5NMctpfCh95fpWqrRRpnRHUbJ
GXX3g/F1SyfYZIOu9NO29057VpKWecTlIoo5PEULIld6nEm6VbD6m0ob2VA/85Vn
3pyWOO/Hl+txLTS2lKnG+HGMFJyzt6wuk4rqP8EwVy5NUFtXTQ9FfjaBS4EgE7qG
vWtKDLOzoFDCiGucU2lFxk5+fd3qey+wspISd/zrp1df947bgPSvm/B2m5WXglJ9
efqgTPuxDJwMyg5ykPLByuKFJL/Hzb4WjkqWu1x0wwrvwroDe92+eu36YJLJ1hZ9
Lk3Ml8lwAUpAICVVBS43bsmnzT/OqEXy0P5p+J/U6RCCPAbQQ3uoV2+Z7exMfYtx
NqrI4O0FDlgLLkl0z82fgaIlaDJOFI7Vw/VrNd58Yt4NvjD7HTcJY5d+BQewiZZE
S0HbImy/qmj+/TF0TSeJ9EyZYGijTCJMrbTOlHIICZ8h/wBEo9npvj6g7ydOBNX9
yswOAirUL9fOnzuWZ4WY/nqv+SWByAUUMDjpbm8WqYuytblIlVPdU6CpSgV49C00
s0Cy4sfO6ZyUwCKfFtIvgAgC7BF6okVJvqQTa9cZaVCnRBN+M5pC+Z+RpK/vqURf
PNKT1x2mt0pNNyY2e6s8+8BYoSnwV0W4Y55CMf1Y8QtpYpDIBg0lmu+vJ+VtoSDg
tQHDg7n5OIOBOoh4708SgCwB2QN2+M057+9uPDM7SEtcqXDDFB84iMTJbm+Xwq3v
NPINLuulDHFBfnP933N9935MM+pLdGIdS+0muZuSVMrWG7F6+4D5Z1k/0w3NjFJe
Ym6RvUd2eHyBqm2YqkcFT50zOFuhvx4ui5BPQLsOQrYGnM73ER4+8pi8OaYCOHHE
IYo6dW3dp3lF8PHDnpa76Vsh5/YCdYeQ0rrPp9ngWZYDyixrGUS8Sb6huKH6wy54
TMEEMPRxH5Q7ovrJwCuCloLZXY/A9TSIBiYaeX1Nljyk7y4OijSSA09LElOObzT5
2BSZ8NQSVEd54EgTTsM24HVC97odYYM8GLwxRTCDgJhn/aDhZ3uj7uZeNj1F/QZq
cBUL6BmNNOdXGEIbJOft+5B7GDyf4aHIsNCzlFoYuLK/eGjc7CadbuzO0upZhe5o
XT0q1CEOi3Ep74z4ttMDXWh0xm9VfrR8tpBel/A1GV182/VYhliqa3HrxnUO3bci
Egor3uMEiqunj6KDamM5TPUyoTOvplr8L4YyDVMAmLVegQq0yqi8s2YaGGoZw/1C
ge+EJoxlVrjvUArk/vGiHQzYSswL57IysAFqYx6njpnPuJEJaDhfQT2vVQ4Vo9zg
SsyG6+ShaCU1FY3XBH2B5lG3zw+eu0y2jLrJmEVSzqMB/7U01TqxQKgWpFnoTpXy
vsK+8LvrnYqrn4SkuKZeMcC02+NGpu3PuTU9ya/1fCzH9fJlduOyBwXVYzaob47a
mcxd4SBoOUBBxcDnEns3XSuIBF2P5gZrwjSFjNernXkefwcXn2ZKCmNJahzFfzcT
4R5Tno4LOm3n1DkC5A/0Gxb6yws56nXCudx0Q01PA4JcfW+uwrpzOBBTVkQJyVoY
2sOpbZ360PVFNlTLRKsiA7O2oMP/HQd6Ut3mxjsn0uMf2uF1IRuDc8wN6B6ZCKYb
YnSoJb4L08DS5RJ58pI86SsP8us5ugqe8wIJZL8gE80Cdc4ce2YUjAdoaaljE2V1
t0WLnYtJsVMwLGlmldgsDtqERsIEe76nxNBVcR+h5FabvmE0X/8jFzSJISvX4Rw5
dH50t2j7MMIqjgKNmEY6EfOvIPgp2ubEdV3I1IDIOdbo+/8wYuNAwT+YQZrvb8bu
AbmqgJd8LboZ4284bWxpVpcgSzJtqxttNItbxiHHprrNkbWu29Ch/JXjgZ6lmENS
Fu3UxfLloNNZbW57cFOXCsMBXl/1CCenqKB7Cj7kto36DCqPUuDl7lLmBW2OuNiQ
NEjdIihEyJTWzP1wNpxa5BDXPu2l3N3CsmGrZSZ0Mfnpk46gS8xzpSJVCJl0pckU
n/V+2AHhEBBgdJGgpWOZ+OHNZ2RNhcKy/G/RpOEhv6/rxsoXaCpNY7M720cKjsR7
5wsSif8EtqI/7GJNoHIgOXFezsWuqhkwSHtQLD32YwgDs6HF+i4GGUNL1J3VC2pO
4NUEu0NQCqjxLntOtwyKwEiufKMQm0SGHfdW77PydRTfNA4iLB0T3dovyzQe4WCE
gbWrvqG9/DaTH0uzAFK31zTS72hhLJDTqsZflwE6qxO07KW2ICBQzNN+J9yU7T6p
6iuzfKxP4Ku1v7J5aHEHjE9rvepa/uawWf5r3nAkIHbQFhFN08yaurCtdBSjem9h
O9nnLTbU5dOzZNHjQIHCJUo+CB/PeoHog9mg4uF5LAZemKZ4N+1cfZCuNHE59gg7
Vt7d3Tbsme/2xtvaZexFoKn0Pq0UXAn++Opn3eEF9jUzzSPO5IeSnItwXV7kpHbh
oUrXgkKsuXd4z0Xc0HE8omdIUQYDtoqBlakWbLgryljoNL8c551R2JaUnHa3gEfH
uamNDmIC5bUS/N/lQ4XgFk/lqUjBQTn8fkaCz397M5jpDehvgLSVIF0uH9fyCRI+
Cmxujk43PeoTgEjkNBoCbnntS8bsKPMpvTwGtPJPxqbSgyMaAN0JQpIygYfFnpZz
dUEPdsup3dCNeYJIZ8mRXTA28fAJmQSe2NJO4KBxPMbSmRvFQU08hEJ8GMvWU9gb
+luXWeERqKpyjbIfirECIUJUv+OHHKjv7BvYNSwareeqX5yKkV9+WvbgoysfCx3r
qurY99kKeqBGo33DBXoLjrNaKt4vL5YPOUAtbgK0VrqKyDAFd1eATdtKIGoQyI0d
RJHctcNXeI/G3Ly3dNjo4jkJToNgkDpJiaWceGVI6Vh5X8PKb8setqMR118i+0Z+
xlKjFgVgOMPJaTav/w5J3xIagR30y1QFdLU17SFF+5a3JeIk7BNhF2Q9m0lZAMHZ
zarUMZAnk/LMb60Oi12bbRpvsWB2wK/yt8ZMI0H3lfmdOe6DDhhthTZDPYftSgvI
rFXyw/ZFkmyYqkX4MSLy7y7iBB1XLL7seyliwxQDmnoa0Ve6WuoGp9TWov0/UCma
R9p2JnXskrANkVz7rDC5xBGaxfl7yhZfl/+sXpsZ10q0en7JPNLu3FPp+9M4oMIU
hwdd27NTfa6FC5HYjK7T5AaRU2HMU0uP3TdOZGjWsz9muVZMVX9V6AJ8ymEjuOOL
Ca7t2CUdn/5naZ2OgjLlxqqTkUXV99biZxBOUl5+OfpRKLWwmztPsaHH0n7WOOvb
YW1+BtYUU+OPTNw1ZJx1d01Qvua7sg5EONq/FhuZgXGbturFOAX9f7fpOJ/i6Ma2
5o4lLlr7L5uYG1aikUmOcULwkLdXjkvvnPPqELxIbiIekJEeI7LkTLw0v7TGPp0i
fF/umurxLAO6aNrRYqnbUs6JZX2OELlHfTcgKSRyLLFBcFa6PIoF4iKS7CdbPQIQ
6xxKB7yBg8NC5Q3nsPGD/w9WuTRApqygAVCBu5rLR4wYrkb5ChlNlRaCT+KmV93F
Tqa4JWQMYj8LROfUklF/j+wYPrs2Axcy9GNS2Wp1va+1rMHX9C6GqXE5OyvDBoB8
XeYOw/d/YR5KqmyQ0rjE+QuEYow8sw0NcRWDvfy1c7DjWCCKjG/GYb73gue/Zoat
JlH7sbhOdDsknqmZJGiYzooxIlSTNcfBJX1HAHMgN82yW+1F7tbEVfLJRbM14A6F
mDSsT7c2kHGcZco3D+lwlxHyTntS7ZwD1HOnJBT9P2vdYUuAyE+o1wrs2htKVxDz
kGd3qFHDDPS/CrEJKwpZQRJSrYS2lg68zC1GB/4F8nhW4JHdvsWKl0Wh9//S7B+x
GwwzZFnhV+PNVx3BEYhnDeVyN68VuIKRYtJINcVt0LoZl3s6WLJDR3OLtmi6Mx5o
NtNVyDL3+VUV6KtXAC0uIWGuy1bGv5ssvG5G/IBWWMFv7ok03HrI3LeqRMH1jVA2
CtqoyTfcwBmjBVUw5S71Qjwn2PwMIxhzewvMl7nyrhcd/+nGlxfN4h75KAnOZpnW
D84nx8YeVEvkySFJFr4BVtz8d+iACfQhE8T+6X9F/7tw+96MRBQ8nNazXCFpA+f8
dllEwzBs5itYNZAKkXJS9QFKBBeSVbuL5LjFakSMhl02bNPLgq3jAtvTjU2Z9MG+
Ei45nezg3bVairuaQUC/BOkfTtJzQ8JTgAQoJ/HJetK+y0w3XM4QkS2HcTtL9v7h
1PtupIPaLEllEdVH2ZFHvAJulelhYWgBKXVQ9PWgdHlJlZu5mW8q0Z1ivaPspjNc
Zh4uPn4DRpzxhpigF2Xi6Djq7YXztQu6oxOzcsjdkA9aXJTKXLz8mqfqEmuJARv/
VB5ZGrLA1fwKwbJm4SUWVIGEoOmiUw+LHuq1c6gNwmGl+QZeH8+OcrOOg/Cp6Alp
5J+zdFT71HNTcbXKbplAx2KUDb3nHltnbDZObphcytaNPvthFzZ//5O2XIg1pUqo
34fIGKUuRUggbYcJbZ5R+yjKBj7JAJwu1EtIkIvvM8B0NbdjkEKneh9cUt7zLHrU
tRiRTFRm5Mp4VDRErcju/+4UY3zivXdy7AKUsJSDEv+HNlM+lGRnAKmdxdupmkEL
+00kjh+UEhm+4ocHUVJ/E6BFHvzURucx1TKQKfqBQVkWcyayXxoX4cxnRkuzi99H
ogRwlBFwBGsiFn8a2kSWytijcL7aSiIyhE4cqG1aKSu9+mkZf4f9KhewpG2uoss0
Err2g1To6+pPpoKiXp+vF5geF2V2nW4kW+rX6p71diZw0O4hLBWcBFO1LyhGcOaz
gefLz9erHbnFotfO9p9VC4Ap0sLdhlBG7Uf1G2sWIm0X6MeW/ahtQnKfxUzRufG1
1tP/JVqd0uIepResekMiX/coydyrmjIDb/feMNVyzZ+5lw6p5Mh/DPDtiVeG5bLu
iqZ8cAVZKScXkQAaKI8igcTIIWDDH1v21kFxNysAtQXYKGcWBX0fsWqJ9HJauguN
8ht+JIVouUNJVy2umzLolXx85uBYRrRpj/0ScVksoQefxGCTXusF/UKbHoGEzwrE
D44xwlRUhIK78dXUKGGGpaJZ66EAOrbqQEn+5plgPmr7Xo7rhQU/hEa/P31aAQcK
XLwMS+NBI8+yVIsB6PU1gQgZsra0FZbprSAF8t29izgV/ZVcfXoxhlVQZ+opCAom
pPqF6xiVAibB3WNZTqyPplS3Z6RsxN21nkWdB1jPCKYTRaQVuxSKO3AG5tzbBoKt
3ANI1YLxdtxokiV6Vwfi09T76P4yN9erzLsgtonR5IfK+fMVFqTfRfA6pYlqzv+7
+dSzBvTZ3+Q0pbwleFV2UfbOXt5sJzmmMAmHrWb10b24hYXKW/NTyhCxVOCapGrt
D1odaYBQt+tSyGUvAJpsQZvQk7N1hlQQC5acD85K74TgHWxEY/Db0C56tnQr/yJW
G9ShizzMg91KBTv4H/MQ4GcagV13gXXTCIZNLuOXt0txIP2eOV/BQ033Dka0hPGh
nUabP9KVljGcLgH0SqnI/EnyLYK7A6bSzcRf/YTwedALwJXvlmirC5uajw+aqGUo
Ie5H7IzRipE4/Fxnk/12ZVt4JmB/lLJaA/0v1x+q9s/WapAeg3Q7Y558D3EmmYjb
4c1sRyf1UpdrP4MqjSf+Do/+jajpzwPsfCRtzuU/6kim/kpOiPdPZewhfcjr0f34
Y51hrOA6mkw0rD+Tx6XBx0BDgxcKFYifbX1UdxqfCJci+84zb7hKNVkyQnY0zadk
Rs9olziwb5hhy/l+L8Di0k7eYW75nu1EXtm74tN1iHoDXQLvpvVtxjlx/PV1UAV2
XUEwkKOjZnzUEFbZLMAPpaBz8LTnYVFpQhn4V/DIOlHXyPFgXkegMu9QeQwRh6od
tkDdRGnQ7I4qBpkmTWpaNto4hwaBiyssWTGq27Ae8d0ZohRZvd4jityngLmjUscG
rCRIIGhtALplY4M8wm7AQf847DsQ6S+LjSdAOi7miUl3mBaz2RjShvZR78G4L7yp
79DPvs1jovtEeksypEUyljDy6hT60JbSBKBi3sGI41rk80c4WnuvTc56kqrlQ0K6
NIdVyq/QOh1Z92m5VZA+dJXoLWx+SdWeH4AyGMsQaBV9U9UPTOWOHdX5BNrCe9qX
qdIzjNURMp/ooG0z4Ex+zgMsFY19QwqgpkLf0Mje5Qbq8OlZoRqS6wgVFGFCbdWr
wg+VWuT4DaJNzdq12oZ71i7+NxaKiHSOrBML6PZxnE47B4Ys7h+/M/zGp+r8q2ic
uDgQhe9AP4+7wDbkwErvKqgtIXssoYW1mxLPci9h7CsZYxn+dzMdRWTW1/cINCmJ
nfoyozs+lh9XrQ8ahKbKeqgBfqDj1F1wvrKAZ68m4/yBRS+2S2FJej+FsPQJyUOa
vBYlOz0f7xVpqyXcmBeY5kakAA1kgQaZO6DhvnpkJPpfNiSiKqPL74rPdID/o/A3
SumCfEi8Nso7vYKL9zxebOUk1FHdxdW+De+6O/rZKw/2qMqmUfl6RINkjqTJiuGU
3Cy7hWTOToZs+O027x/2bfwVXaTO9v0Q4PWr5DmFB2txR1P2HmgJnByFYcUB+znH
Xau0CtPePBoZaZvNMdeeipYGpi0WaqDF7ebbY0/LR1CzV0/lanyfkSjMG66p+GGd
7adVvvXjjfewjMO/4ZCBh5AJmOXYMkl7ccgIh4dtRddKaJeayLvptX9E1H1ps9C3
P4G252YgZunXrfLA7iTVNdoQEzc051m+1cjTROxtz/6X+LtvxKBSIBCxt9f/YcDY
UbXCsTbbC0whsoo7igPKE0k0iNi2Z4zyLY4VvMZ6IGXyE14Q5ANjobAtY/r3v/ll
LDx9EeoZIV+wSkLVdBZyZLqDTNUdhNJbC5BjMWJY1ojr9JXLC7uGOEDLZH9MdP0x
ira3RriHQAlKwFU82Vv7Qw8bRAvYCDOXfifLCKdsq5zce3NO0siHUcH5LEZ9ypzQ
rv9p3EQr/A6SjGWgFtzQvxWKjcEYVY4Crv643o7H6QZ/9yfVjyY7KKl3gRLdu+UF
E4aPnfOwNxLorcPjLGCc4qjYuZ8how53xrgVbKATCF6o6rUML6+xTKsangtY4KVp
UEH5alAx0RmbVe9WHbfKZ3m0mTmR8zBgUanUkWalDJ+fkk1pvKvHVq8qsyvLzzUw
pTVecJwvD1upoQUnF+SWwjXUX4vHm+Lroo+SMuxBA+/1i9HT9MfGfksUQJpKWORm
mJr9bSTq+FaDGfUb8GIAcV1sFsxl2IU3lLnfVQZrXcytOFuSMjneLQ1LigZ3c3T1
iOBxyPrC69hJ1r/IiJU2zPrtcBB2ipTazW4AAcUHtdwMYe2WjKciDHswdxxrynz2
mLX9EZtAZBaHlntQMgeF+Td2VgWvbNJxCYcNhIvURwQF33W7z8MeaPkUS5cD/fzF
k0C9Vd1nX0NoImFWF3Bm0IR76AHBTi7O7Uce/ogzh0IsoTCTucTeRJydDEjm7H28
GEd3GNE59QqqhJG/KlQBlrXtCFACMm9QSH1FhRCxC4fSW6el+U34wGcamh4SIpDb
EakuJChrDsODcPpCOZlpJNYAv+gvGZFe+ZI2M1T5T62K4bGCU63MIDUV2VV3Nh+F
J5oaBKpL/6/6BVFkvTBFlHCPS/G3ykAFL6+qf/0b13jEQoeUHR6MNdpOKbISFk1x
R03xp3TxBSHpazLu1cAb7cdIY7mKjLxKI0QLNjOGE7rq3/hZ4QwwtbkiEktkLA9L
6CKXPfInoF79n/3LAtDlld42MjVhtsamw74IGTwdrJznOW08NwVfgjUi+hOj2cLg
vXlXdrjs9SMRIMUZO8x+YRCI1UTzOT68SC9vf632/pRMvHwd+V5JFAsI2j8nrk4k
C3lwd6F1XzuJVScf3GCwTKda9E247zh/stz83tR25k2O2Cr6gpsurN1egqukn9yU
/+8C/NS2cFc5S7CVEkuCcRSIdKRuYb3mXd+o8GEPGmz6n3frHkNjMT6Cz/ITGi3b
NgYpj6XsJxSHBgL+cD088ST5BVYzTGXUI5bKqIpc6WKnLn7xlkczvBlESMTOUXY1
Qo7Pa4XXUY6kJm7hOpbdUwOMmH7glLI2P5lDAtvVGIjYiwdcsgP3gV7GYxDXyjTd
Nd69jNisVwHuFMMY+j+poka/ics8+XoYwP3DRDZUFvC4mfAsrGDpVMzpcmDAmB8B
CuwCEjqO1l+1DsM5vDkVtycJ3pgE4D70OcPt8G2CtmNuOD8zKeUgqMc+S4lJjCCf
p4IeJaontDjWYGLgLruK4rGH7gZ8zCcZTZA6wn2Qrq0qp7l+PUzc+EWLLP7vSkBj
5uT52N4+RpgCrdAVlv3e7VRHZjSa+PaAh3qjrpn8UMlzYwpMqnkhM4BMnUojvaT1
BFlaSq76Fi6Ch3/CmK+D4od6NK/8zrpcv636Q/rAuTU9G1TCISiUG4XBT5toAdf6
Ea3D3rqiMq/VhzOvA73da/QKm9jXwGeC7RBFw7HaiMU7HWfWGMeKua5Uzkalwvhj
Wf8l6mCLAxNw/aXVELmXXq0pFX6q3tWwZ2A4KqnIEuXZaEWcUREP96fl4CKeCDcD
qeXyvlZVMWcfNDs3Qk4qLS+0eR2X+xczILhMjjARCjTH3B4Pw4E4jdEOar381MmB
osIKE5cw1SoH78clK9pRNrPVdc3pJblYRHtjea/rvS6sdGrhIzHZV3ZfZB1HMCvZ
hOmaGsx0mIEC+hk41eGmD0p4NK89ETHUc63poAPCWr/0mDLS2Mjvoyzziela4snA
WxXuFQKZy3XAFReJ06GVMeKMqymsDvTUXNP4rV6tvNQxR2ngO55Nn+5bb2PyQPw6
iWDsIUsTfhm1JqANlEsSwZFK7T2I6WFPG42jLdJ6s1vxnAznQ8bAQnwENq6J5nBD
ovgDz6qX+O+G1CB1DfsoT/6lLLW73zP2Q4H1aGlMESXIS2AgWFJdmKLxhKmTTZBA
rUUomTXWMeqBB47Q+OUxNjSCqLvMmfz+treYZJvH5Eq0RRbKRo7r2k/59v5HOZsy
1HtsYqjDLTZdUpMSmx/OpACjfEJcevOd702tz0+RreF3wyTA/RL2dqOt9A8xPOb2
Lwo4G2Iuf548eXV0v0aNtIlDDc+hvVZRKFaeI/5rRvt/rev6jxoRHTs883fYEfu8
aoIA9IuaKnrfcPePtcsEsvok7avfs/iLnaBFkNyJNqZVj0IWG32Xar9OHVVmY5CD
had74ZcxcOQPYXadVSfe6ICbA1iP2i/DRY/aMuMuzcZSc9tkkA9qOKd0CfiJwkvX
RDF4esgO4Jx7kXrp4LJ7X1X1pFhOT4QAcH49zGwIt9+tGRrCn+262erxoQcU+nt+
ONzPyU0fRvixF5xG9a0L92UgH3rULZEjZmtKiLRVHwnwpCDWKTwLwNS1hGYcZ5iL
xBnH9oQm2byFC35xZz8rw61OiOsYpq/8kPuykrU2Vp1i5NoxvsmXZeLtzwIgup+K
Pw9nstRQH7UBOusClx5BdBWFBEuaL58TWbdwj2Wst++Yve2sAEmtLkrxdH8d89Xg
Z0OG4bNbeIgmO2CaxGo0XWGmNcr1h2153qKuELog8JwK5aAWAPl+PNsaqolhuJhM
+s33CN2ISI+A0TObj0ww0g2VPAZn3LmTbSGCjg6kPZsyv6a/WlrwBH5JNrM0fvrb
3d5N2l8FAoam0OzyqDEYIBTHdojMFvW2ycFJwbluV8+PwleITVwbltSaEbvAU1EW
xR4yuvRReXXoGjJUe0E+NE8EPjVmO/pZMXLmXXvbeMk0IkKpTM+b2kZ420HhHIAk
qZHU8Lz+3ssMOAVIdOllIo+/y1Qvi9h9ux4C+yqdFgHc19Ciio1WYEI2NnmO7fHF
PmOvA5wtVJrB16hfi1wE2cncjdgFDMVNc3YF1rN7KFoH1zthL4ocxvFpzDCXScbF
rzelQ98xRyM+qTTgWujpgp55IjsxhE/X9CheR3BPe8dDB0it00WwTtz51Cgn/xmj
ocIReccdAsnwYvbQjznIGdUn4+QrWjnQSK2JuLCFI8KF5rJ/p5VfGJZAPTWAqN4Z
Prnf//G1Q+dzIwTZbrnJ6dZ3upMkYKnmCM2RQ2M4u1UBh5PS/oCVYUc76cTTHmCC
8hAbxMU2IVutObXBWBLHXLtWy85/9Q4k5Tr/MCiBKtiEf86rL9eBlsdeXZevaQFo
nvsp8oeU6nZqfJi0voE2EoUr3j90rruGXj+/t3LlYiwTlMYBQs9TIYG97osWnk3z
TGD0GU/NGgCCca/SL9WtD59YCvh98E/WMlH2uGBmcr1B5/csMwvehXM3djNe/mQP
SHG/lMaLWy8QrVob/2MxHWVK4IqsXYvSbhYKsGByVG+y4XLgkzMFWd9zhXgEDVVt
tOmmoPIb5E6PMGaGacAOnHVR/cOKT35Pbv4NCUb+urw17Nh7b8USAQA5mvsKSg4/
BIp1c7udqzCGSTgVQZ7WBScH7N5Nu1Hr74k5DQ2nsbf5aeKi2UCkpt7QJhfxNAAw
4TdJ+9LiHp6cLAlhARCPVCbcR3L6iOKSsZWX7j1X1NFAz0doucRGvvtDj2dPO7YG
NhniabbFwW2pbUFsaKMB0PUnpLnF3k6EFxhbycwtCZRStMgEObu9l9lbtpKZKv5V
hBZv+3ZBiKuJcuYcZDGj4OM0YqSCXDOX0+B/j628GrdEwS6YvlnIDipAUWORjKJt
c7vRlsReas5rgwnStp3/4+vfs7380hBwXGzUVSp65SqXOJtjCS19MW5X3kedU0QE
7ZEC+UG7lz+VI/Y+NuDrx3CZ2NxALMxuZ6QxNXsrcLUZkiTQe48iiMPv4oCngX/u
lXSS4PWslEm1NkhpJ4w33Ojy8dB/iX7lPdMQEMxsq/aCqPLrVRzvjBAE6DHv0m5N
bskZgmsO8ALIMcx31+mjHhZgdBa/lQ4zHMShuZ5Mv5n4RIgfrV9IA56ueI7oG57A
ivbNxQfpVXXJqO5PKg58wz5ApXTZugdms4CUl67hbgejvgfELJ2aQxy1jTJPj/Jx
B6AbVmyE0p75mssHACz3a0XXzpdCWbJenUuimzgZNZUlC4LK8z6NmsAJC3m6e1DK
+VCQdnTo5SfJ8ew3C5pEyztTJ7YXmRAMLWOrSx+F9cU6RXgF+5RrFHqgW4DUZsvN
HnsJxsMYzMepeF1fGbtGLIVTn+m3Z5eAvpLgGJoy7PlWwjcaQb7spT1csy2dmzOo
yRhqJAlrt7RuKmmwZXrJKc5yt8hS33tPMS1JEwz/987hPeU4Mr3RKJf+uD9cmMnO
XRd5zUFe8CybLeinGeZs7KoirdCSTJUkRHIpdKtMqKZUeJYx6MdkoaChU950Xi0Z
vbFuaN1fl2jSVA9oAWDlrxNmN+Euru1APd7f8ptyZ9nmwQ8Sw7PX3Zr2cwN+tcet
feRUoHxSjLRfkMLOsSXV7qFkeVO/it2odEhSwC3PS9hmKEVV87V2i9LNCm1pkiq+
+3BBEfLMOGGsNEhyewQ8ttHrycbcmLcVc2d6j9q2yUpbtC2ula2kh/4jPmdg2T86
+QGy8dh/yBAWQZyHuXHQKTxojHzUBfNze1riGksE3QYMG3Bk+g7wvy2DCnoHEXQ7
Qy92GXrDWumEMN0ITNImMTFULFt8pYt4IOfs4+qAVup+1r+Hrc+5tR687jvRAElh
KaHyG706RFlsRpYub5tcZuu1tZGO2UxPKlvLQqFDOko6WuxrjWD3pwOSpRrQjkql
gH/ICGtUgOheKhng5drsoGbBHHn6QwCXhxD14uuxgicoiyQdSR4ZwtSBQEG0ciz1
XTGPZl1A1jqPjtnM8X6SmF0Y13WmmM8gRtHV+Wj9LKLUwfkC9+4XwfRd4DqIAMHV
qxfLQjPOSWc99RkYiNqGlqrDKlqCdlm3I8/Dx4xXmj5+orNbWKUGzxAwnJU0EP8H
H+kg3e2mIm1/Pa3EmRREuOAt4eDvBoXMcfab8MXsmJNsfTv71ibu4T20Cz/1hCCN
RpVwpQOiNHgbkY8m8nHPg65x/FDyqaXQxprB9/vuvyYdx36uRuJCtjoFf+t852CI
tFvBj+ceA4PQvOyRalfagU6pDQXYvshsCggMIhzo2ra0pAmp5Re2STZtet950whr
yCckHgFU1DczEuG2KglHI7plQ1KQGWxANHG1g9z0QxFCJ5JiDC71HHmTKkDRFVwf
awE4fxV95A6WHtzfPIWKehVeay8f5BU7VnapwuZtlAQ0gX644KScuQjPpF9M3GjC
ngHnIYkY0M7d/DpauKfKGzAVGDSZCiJS2KiFdLp20I0HVMFQ/eaUGSlDayuilyPv
q1pxxqAG9AI8MaZ3FnJOe3bW/jvUDVBOyWVMY07djpYpWKJ4EPAS7LwI0l2eunxd
uEqTCIhiRS3j4X1ltYvQ+YV5zZI6kumhlll03555WnIr7+1smHPnsiTGSc7abtfl
+0j8fg+2GVJJN9/2KFiD3JmUq13AT9VjPfA6XfZxSGYtafDkiLDxwZUXEZmr1BV0
KV//jNS9kr1T4ltRiyPyvF/w7ARyjXu21cOXq3PRJ19H/m2uA7I+IZeVJcR2mShC
pBWOyu6jWLf3JTQdu0FVInafNrJNTajVJhEDiWQCwrvTLal8YVDjCVz/PvpD0qxZ
WMSLLRePehyCrKCk4qZey8/HzLFD4h7+iNKmdExdqXCsyQ8QrMQB3B8LBH4vsval
3TbDas//kNF+hQ1UYZBSkmbrxA9hv3PdsezQ2kmrIXk90LV5uF3zR+1SewZ9wuSC
DqoquDNAQRzNrZ/u8fwRpprsJet3CbXRJ2Mdfyon50xyzog2KYoEmPemVC4SEpPt
hmnatF2KeBPMlV1SzfZRD3Ad9JD9fQQj/XoLRTVU2cHtPvvsnwI+H+9ze9LhlbCY
1VGY7LwLqBvQ/Gi9Yv0i/mh6+4zUAk2lo1cYthoOXdyqP6L1p3yEV8cFY0U8kY2t
WOQTYFJNtzXCWkDEc2kCvVTSy7EysWvhXwN4ZEuzotNi08lIa7N+U8ZjV2NXirMR
sEL176cuumMKoMWuTY2fJSfncoHQALFHMyNqJkumbXnRkkcza4Yt4fc4YKtOF39V
TXIEQAQ/4f1mN3gLCck+zMPCVOi1YX3+/mQTyDcWqgs5rQdwuQTYW4PtLENck3VF
gUT7J7ALV5m7ZnHruVJXfL/LUpk7358RWUoVKbQE2Jk66slSVCp3uq/QW4wSYeml
8b+k7s/6HSkpypjhI5nL8pmsp7805/zug4YEsfPO8WAD5wwA48I7RQdzdbe3/Cmw
HFmJfPiKYNwNnVq6yeXpxKd4wLV/gio1zj+PA0cdWg0fsw61+wJln7g6WkvpEU+C
xc0PBI/oWL826z1NV+j7/dlIviiXHkuOucQE9E4Qz60dIhYS31QwhMXtvQQazSyI
Q1g5XRG3hQPQQzgplhLz/Ma5zFVYH7H8L5XTYsAhoDzcF6pF3sKqMXt7TVcIVlG/
eQgT/cbrMsxw2sWlXedwaRVIFmeW0SN76W6rax7wR5Kk0bIh2LQfhA0Tu9iOz67z
WvN9LNwzhKKqnrnC3SNewy/cluyYnQQHmmRlKSeHIa82mzx+CYd0i5bhOtTTu35n
obva9eIuB7V5nOZedllpynXi7ixJSFIwiKR+nBBNmnN+s2dO6q4ezS96cSngx/2w
rSlAkDekNBFCeGqJ4/VanLS+9+UXzsKRHAkS2+cM+z717svRtD9bvXcUbxu3y8Dt
hfgnai4qcYAJ4vIwJ+uw/chp2nb+AXQwV+MqQ+1VUXFvzR3PhkPovsCAAgufqw7/
3yybB3A8frsto3cPQV1VGl3RrDkb1TcO19AFxVDyMTcCRP2MDYBXVU9tZYWjtge5
3NTC+slILtiyX7J83LMNDOD6rM6DQgv4jzjeC6N6vNEA5Uoq/NlZmzI/B/THEnpK
j3wz3yWk4Mk01U5sKotOrwy6r+rrD6yJWlEXDsfgEmWKNf4OWf6ua4Cmh/RcGtyZ
RxkR1L1w/hqTluy+9hgeOEy4x0jSLGw0ifzXgIYXrwwQB+bUgqORqiKFbNY9zD8w
UCEfKNbHY9wL+M3BY+34b4iwyJttx1mgIg7EgegAOsTrz5WWL1lvj/e2dWU8gM+s
FEihhZEFO/P1gJt9bfjiK91JjKcQbZJAKbnl+Qo+Rxog7xq3p/woI/tjCZWHuzrI
SxCE3KufdlXKH6jUdJnt1HnGr/FmIy6YqU03Ms7zQ8ijRyBCmRae+HF2yjMXwoaM
ptNyuLKKAkUmF56eou8qIr7xmCzzNyyZpGulDyZ0CshrjTQQoeg9bkasm4+yApD3
Ml9GZS94CBgqb4yKDasHB+QQ80eBzLpeGnlDVEje5Gpe5+MFwmkWodZ+3samaaYk
2Dt1AKLITQohvPCpua4qkIu/pKod4unKriHJx0cM8whJd+ZJ4K+CLuqowvFjB0/e
X2uICe8L722nRbGUtREvJsHbGQANsiZRcjwt3ddFXbLoCoNPcmzraTui3S/STtMx
nX2ViTaL2Tj3sAbPqHQo3Kevv9RC0CgUTAFGtJ0+kn27/c9pSORMcCl7YKvCK1Qm
n5YQ8OW5XZJYAePa4R0+HIDqujs0VrxVW7PKvsxVMJKcLygL8Kem3RniKTicwkbe
JFolF1hK/AK5aFh3NjK1dww71LomFim/nvRmVew55dAH11P48IL2GZ4veQUZ9IIN
zLIFa9xLB4vuMXI+S0HsFcF1rvKLHKgLH3ZODFWcL0UbXTiZ59HuP43dOB2dIns5
yJq498Tyf+oQEmEyiKBomWM+zkasrrf66gtlZMDflIaJyeYxJE1SnudqgGtBB+BY
wM/iYeVcMdh8YtEXKuRcw2mlAU4df7gDfo5D+lCfPc8aR8HTn8Hj98BU7kT5Z0Bm
aaBjKh6YUOkxT9TN7k3wWzPiWEr4QRJruE28qr+zHeKsvILTqkoScyDqbrrVisYf
CJt+70gYZItC8eK6cnIUzSXQ+UtE9gWwcEdDHavNQVzqyGa+Ae9RZhMVjQCubo5J
dzUMu9i4eP6M2NFOkF+d6XOUzVpBNFECxb0OxpmN7FnLuyHu6k+seF47bDnq2g0c
d32xCxesUpT7eTAkZPL7sLHmZEq/ycoOD/BCkZqJUodV3JFf+78EtXJPt/eAXLdi
hOH5CUMqCSdlXGZo309F7+/ELeilObodnxXov3CpnI1H7lHy1MoeEp4/lK2DRJC+
3/GKstE/z7DP7zETFQ7oIyTq1CUPp1eYnu/cQPhJte7sDy6avO8/RpVpxrd1COVf
fzgzNgtmLN+rraVXwjVw90rTiUdOYVbOq8PUlpeQNFSbJRDzVDjGIAtAgLDsKD1o
wbWM6bOJCuTOIWAEA0czARsi0CMrNerT+8IbEDfdai2xYpk1v8G/TJBQyLDTFAU3
QX6+02OQTB5lTKjP7Eu1L8ke3qm89EoNt3XAgJbyakkj59nXJO7sizrdl5De3JbF
aEeE5L9pTaxoMRqk0j5ozIyKiiX3O4xw3LqMjt5zD7lysypP6GUcK+RaSFHvP8r6
nWZiJBFWvQeafkwLrqwgQF9Py+TkYb+7Ptgyuc3RwYJZpWpP3vF8mUHkURYVw3Rf
UHeKci9D2w8owLhJ6Ek8J2NAuP1GyDUDjiske6ZFRjqQVQV44LeYQ1fwURYztH7N
t6WaDN5AheupXHG7YxRkwY5VYMuQyXzq1s/+lY8Va3IVtZNB+erOJrd7Hkfhcm2r
UvT+PSyUUVkFp2e7BPFymktyjPdo7Z6s4F2Oc8S1MPqE3t8/MRS6O5sEQzJu2uTw
rmmN2t0ArwSQ0B56b3qc89sXowBUuta155qsQ/HbsRP1xN3hVAFdJIPhgXau7gfY
uZlv9czyKNPzyXD6GYYor5ueNMneJjocy75l+7oLTe8+EbJWjdSPQXQFJmX+63Q6
ulFsxQ6lUS6/cMUMY8eO/26VTPoEeaeOQ7Fs/4PTh2eqTY7+GwrWnemDi8+gxVn4
dwVaMaVeksfHxnLrXR/VPb9jRhKez2kETkHv1XtdhFYewmsLyIQJ4+Jmti94giu5
9lDpurRXosWWkyLI1eWk9zdO89MF8KfI6cCopwp3aVtDy7q09SSVeQYJpQgCQjrr
dINcW9dwFeoyF/uCE07/W8M0fbX3H01TuAUjK3bAS8swmg1I1VAxLMj7OLTxZCdy
oo98OriS2B5sbNS7b2nQ0RFumaKpCWY/gaObBQu83JBvL0hw2hBZq8MVXZdbM0Nj
wRhyVqrnH+JneylEylC+eqpEMGbGh3aD6sdk3roTMK1JS9HiPd3K5w8vMVl4T0K6
LwI3XXznh7KfF2fYe6tjxbiRAJhSZ1pF+oq3Gdwfw3Slreqg86W8trMkC4flUIEq
ln1CdAYDGvnRKGm5MVy1GOhDPWuiSXM9zWZwzhrJoAp4Fr7UUo9eOEwWUvDXjP0x
8MYiuxaS2ELCCsK/4tWQHNuSzKIMaworiyv7gsmThzzjzY3178MML08PMOH3qGZU
k/fIHyHmPGm66SyUm/CR/60Mshmxxc39a5q3GWw936ALOTHYA5kFndOiCos0ml+p
oyyaA0FHvG1ZXfR4Q7nd8ilUcrDjHFXv3/Z48HvoIoIQhlwHQ3RB2PtbtU/tSWJn
TBRo/RgouCYsghce9Ins1pgwsd/NR18UdYrR3q00FYT479icb+VEtrWwFzfn7DDR
gHLAkk88T4/neIuwqbaiXXJxkfqL+q4qP3F0XS0Os0QEtzkOVOu2b5nlHBG//3m/
ESkGYB8/1nIj7dvpCARmcFTZtrhYiIlo6kwMKZeA/lVBrmreYJVDq4UcGKJSTHHq
pkWZRAOpfGVRLaqs2/KFxTGG1qPOL4eALwdsr3g0z8e9dX2pSjO5l8zFr1P8yNGO
3ivp5koKhg9HoYzraLnj8p/uhm8HmBc8rX9MUF9llOlQ31u+MHVSKVt6v8adxoHB
5UlC1dtOimfsnAhqfYPflN2oND/lvFRziTG8acpTSjp8x88mbDRCBcPTjQ5MNdMX
KW4TFprQ2CTDPabdgkB/gjTxVKbDG9sbAe/Z1g74ydely+QFyzD8fz+WGwU+IxRy
4sBCfPB2t7FbpwCBmlxxe8aa4muy4dZ7r4mGpJ7sVFc64NGoOv9whiIswnNeMTT4
pYeVIGHwxcR3eBY8sOmWKgGFDQoNRgaLHz4mcqSLHxE5HbPIdPw5V9zYdpiRhpvj
j2UdzDcNpmbpbeKTBMTj3DPz3uzfBme1KUo3NF9QAkRTGEenbBXbG0I9EXvVwJfD
3MyLxGLizlc57MYqwFubJRiyHPSJGuMyIXXU4+u/K3EYBDRJp7qoGKbgiKiRLjAZ
DxzAmde0Uq8P9xV/m4oYEKEpakcl3EE7s5llyYUjcdEPsW+z0vDIqV3p4j+tyqqf
6XWmBJEEJ4pyvHLwB0pg/oXCZWx1CuMM3eCAOEz3NBRo5YbcVZ/YInIMo5S56+27
bYMjNRwWdWYLnxvAOF8JhG5Fsj6cRB9gkiC3HTFwHZxD/p3HZOqWiNoNhKyq2yRw
hhq46W2rWXUpDvSOSNrWPJOHpjVCwT9gcPJYDDjeJYoovzp7RglL53kEYjTbuYkJ
+Vpw0VavVUYK3OBTRjBQ6jdxx1t0orRH6BZQBqQiwTLc+jTEBdB/X+jy5EqX1aJT
sqRRCAgPll90USxDwkw7gUZNB+2znoGd5hTXJ6onE/2ni6E2fj6JxFhcwe0jsMYv
ec3sfacktTmGIU8zb84JiVqlez4kJFmXJbiIJ4peqj7g2zChEzcQ5U2r53SLPeI5
AZTMjLdrHguxEkOM3JRpZcE09jlieUc0CsAwqLstEED1g6bq2T5nB5dfi7NdTygl
FfYs2+1gPAE+nRNdniQ/I936HrQSC8pQnjKFcvLqlESsRLZEzi6GBi+nPeaWkzo0
pNZrsb6Lweccu9x1CynIOUGijVbLZVVZnW3z1UKu63uOMDv/5dyg2DfAp4OB1x2Q
RGjvdSyn3sxKhwssMtfMYWdu4pWvDkRbhj3aJqikvf2ykqSV+CqTPsqVyosneFqY
l6JZih9bB2T68tHQOm1ZCAnkGF9oqnlaR/K94K07E2QLelMglwFGhjFQD8yufPWP
oV6JhYFxu1A4n4EKN2oOAvRM0kLtGWFImkh2iDxqqtpU7B26x6xBf4MwbsYuiXnM
OtEfH7WrViIg0++TM/Mn7IgKks6747jB5s2clsQURsMuXLnFOGYAsxFM5zY310DM
X6BktKBlZoxinfV1CL8++/Rdy2o2RDMpqx3sdWTphcIGXUtMQYIMqg0T14BmBl+L
0qdRULcRgSb91Od5ecSBwFw/GQvVdJ6H7NMd140GyrWOOtcw+6FZiPs5FOB9Capb
lRYvWxegvIRc00xyulxHVDKAP8BnXzKoTl1s6b3hmSZ5o+PnSI1fPE3Ud3tCu+Rp
l817128Lrnn3wZeEL5v+V4un9WHLZF2uQiRqBxyh0l8ahqxJQiXsTpL/1g14Kwk4
PCIqHkpxEoGUghf86+Z21vperIQdkU5QwLRhbJMwNgc3llv1V3a7I0+GVwESmuwc
b1FeCYlbv1f8JESCvo3OT9qguhx9ISTND3r2anobPsvklw344DnfWddW8idMaTtH
d8P25GgVe086qdHD/QzKIJARy4XJ82X9kfDcZhH8KIzFL26dQJWLr6RA6KQNn2hn
Fn5C1Rc+1wD1rj+NaaX27t0yl/glUqytBn1SpE58Yu3XEVUn5qvmNN3+u1oD8kdD
ugbzt4yDa5pFDpZTJi0EKIRKbXk2b1GxuzoQI+O6FW0wfYrZeSjsm4tE0XF7apdu
HziupydhEKTonGx0c6IgBCTP/Qesh3u2qUP5dtRXD1XWyP1pypPmi/RD3gTfbESM
PIn5gA02cD9EA6OYbGHaAj0GXzpPjH4WaOQr6Iv+lahfkS9CK7eMgn14HXfdX5Iy
YZPDmuxfmHfsISapQBO/gNqUMEDFk8Gnh5tomi0jPkEyTLzo5D/tnV8UBlbqMU8K
H7P8aROwTTEBwVY0JeE1xtjR4hXblWX55bB6CXP6PjyMZPW+NvmpRUQFvdGO32zA
6uUVytBQxth0NgtKe5MitC3iMA8LB4DuWD7SjG60f0CxZ+Wd3b5ipve8s6/Blf9E
UAggBo+N2Mr8OjDOCO9PBhrbEh0G++X6r8P3e5jGfVlpvVqpMqJYkTwCVE62db8/
C0a6alg2LtII9VGDWzJ7DYnfwc3hgXZxCFMYMpJbEvDPKAAiEHih3hZinzItv9GH
cmi88iQVx08UhjbZjzqOronQyfKmbySjWM31tn++aj6lyQ/4qKPmvD3Dsq0Ezpel
mo+am5oAJ9BW9tuUKPUbiO+JSp7b3qjgFRu8VEqV7jo7qiNNmBLSLXJtMKn8G9K3
CgH/z7tBSvtG//sXoh7SlGEGZKtSxwp8rbjGZpExko/JSDHIpUPJ4esi/rj4ej5D
tG6rqpIMc5afuYLxUan5r7mbkDMT9/rY8Vb4/lC6HeWSQGJNpWSO+cM4JAjtby6j
WVT8RJAVe1pQysjtC2l81/vMx0bA0pDt7nzEI6aWOGuTKbT4vWVuE759iCbEYEfX
oSYGWtjuPEOq/ynohE+n8+HpZlMcWg74aYFeNCD/vtNwXPoP7ipq5Uc9ppIUWlK+
33apdiRdnh3voRuxSFXGGSCHOXaSwT6xf/QzbhB1eDnHuTRhZgmWxDr84D0VaETB
W80bNnFX4vS4KkFUpHN5IQKDSoGmeRsDDz1QyGblCpG4IUnuuBGIGDF6vNT4+LnG
jTeTqf0qnECmeIYL7W/A5G9+TP7UBOr6wPixHLeVY1H7j3V65hpi6nOz4+GzJpG6
3KKhptRAfMfPEpeSUOULIjWHqkrG2n0M5S3rpqu7dVJpdQk3GGMj5Nb5uY5DwQN6
VyfsQ6F4Sg+otVB/wXKSdsJVeVNL7CEVF9Y2wq+6zzCAooCtBdCcaFJGg50Ua+99
c+ifOogtQfz2tqZXQ/qrJH9PS2zmPiOywzrH2cf2O6iQHKr0HEaSaBlDGBtJ1lEE
A1lLbyJWj8eHF+W9FFSkUWN4RVijUq9e3sAPA2Qwt9IgPqU2A2kNmo9RmIXbdBrk
9cb8O2K7bdNJh3Gc30WmIorw6Zg7ePSxACn7AIVNvPVDX0g69fg8jjQPXqtf2Mns
A4D2SuA5V7s7jVPyHf73kaDaGHnEGrwcwDYc1+nJQKilyb4Y6JoGTguMCpCRBkO8
XyacEp9IsHi+4ROGWAku2/GBCHrpmnSKYDkATJ//zycX/kLvlsPvWJkizdw5sWff
b1KaNCKwSI9yKPnT6R4jytVBYHdM3fYvj+l+GaY6hzoXprHl11GAUb8J2KfAk9wj
zmop4rSZWKHUDDKZ4b2XqDtvvFmtd6yzBjOz2ySAw9xX/cu71dVHexk6+S0fX71x
rObvbsIA4nf1Lqk7laFWb2kSRSSjAnbXxQmAlLOEn2BHKw6+/fRVzrnqtEk2yzYA
oUr8+IMTbQr9Ck/wmWX7f35pqWnbK2sj6n0tBiQIVYbSeJOFwUUup08IizC2xDnD
zG3SiirFRwG3JGE0cBdKK24x5SH4OeVLQyoqQ2bO+E4C5mi67UkITKrEf2q7/eVo
hP+v5SyFANGA/4UZewyhVJwTvuAHWyb862kUAVjxnkUr9LaNBtTkMkcVF17aA3nC
P1/dZLN2BGxK4zcB4Ar13wA7AQ507aLOQ46Ccqy1W2XKk+HlYPV2+P/zaRMRWi/6
6L94NxQz44uG4HFyEmo5n0F8HgMinVm9GLpfWpocVh7Bs+380HjxIAmZgxrM+7XD
gtbAQrQx5KnnrCVPBKqnf+LenVGC2C66rsy+VlBmIz+wcbqQqnB/VFJORvTqBomA
vbsciUgWKDg8i4TjhsfFRI0XCTNmqSuwfrj4Kd72YjY7RtTI+Kd3fEoGluhdMmIR
4dMxgMKiRG8KH3hEUzMG3ngQ2W0lke82NJPcrF39U9Eu3NG6oSytGHFvn9vZftdB
mILxj3JtJyuahtNPS+2Ssu9TQbw6zjhiFgh+MwGBvHdBt1uadf3IK5EXuPbOOTIC
tUoXNJjFdXLg7nVMQIoKE4/IZbUW/hWY4NSimYYKMnOYo2jus2TwdBGkAR5cnHgM
id9frilVe5l1OzJMohJ7sfKAx9+RCMYisC7FOGsL4djIVHEgaNadg6cLDgfC8QA7
zf3T6dVsf8ySYEqfoQpMoVmVlRtzH2AJd8sSB+5mhSDKyoFblCojdTtUHtlkZgQr
/RW+qoukaRymDsBIo0zlNHyZnmjV5eyq0sSqo1TgrhXoEFOyDM6tUBL3WAyMo0fa
d18+JQH8Q9v1a/hOSYjhs1wjVav/LNnutr7uCoflfaTX1K0M7B7N1JZeHt4tyDCu
+L1LC/k47k8e9Jo4P4rFvDcPK1j5zE0SRxO2wJhp4BVw0UZJA49J9b05Z8BiS/RU
/RzCneVGCWPbijK6laPALi4N9BGQkVmA0Cp3yeumHUFf0WBSrlO2lH+ZCVczXjMW
os2QQbX1FpOjVQQCa1LOFmbR+fA7w7lPl3NI/Cm5y0mlrIo8oXAIt9wFzTJ1K5ct
MznT0n0rJ7yKK8YUlE+wOA8hLA+Bh5lHenDSrMR4zws16OLxpqH/Lv200ZssggE+
w3eZ5cb3I4nI7axhiiuR043MNAYLdmrkN2gjiU0hysz3G3zFVBGW5jtxour/Lec5
NfXiyNbwZ+S94m/ieum45zzlt2Lej99lNARpjKOqCo5jt46L8gKSIZndYtthyXmU
5aTI8QIauTwgS7Ci/koRCAGbmxXEq/6ueLdvuYCVtXSxm9zjIizg+Ptrp154MFw1
Bv9oPhqUwneHPw7grZ9tD6OWDPCAfB4VgSeFWWCCdZ+2DPs/B/LC8cHmmpuJXerN
0kIFGduvphLwUZb25CrlRt8609t7ZUcO7d2Wtqg/X1QKy1/bwYpyJu28hK8cfB2j
weWOAQDOiewfAux54RUdFfa5HVrnD/8C+x0PxseF+TNgOBUz5gqQJRKeGaGt5jVl
sRJWahqCcr/df3sbfOngkM0hKF3GtRf/zpYxOBaw6LOQddStCR6OGEbRQ/YZmUts
cwHZOXNnolv/TKwIL3yr3eHY2fY8QAB0j1aHR06iYJltGajUhnYhTJ7yBLEmgG4i
G2bMPT86IbL+AfZxwMG7stG95kccVO+QiG9F9KkxXi1qNwoRmu53dI2hfbT81SmZ
qgLNeXGVSB8gxBlSHcB7PfDg9QBxo2Uq14+RKKvH1i111yYnKPnTjQDHIicbefFE
ygHQPZpBuHl3zwwsdCi+Fn6HqkVg83L28++mJyuO0bC1y/lx7PKUSkD38L5NCNnt
bc/WmGJDgE9rPHPLz2CQcTbT1Qzz6bTjmLXiqCLVUEdZosGUOfCicGHNgVdSHnB6
7VVdjoYDA9OI1kpx13iPOEGbhIUY5UamszS98/W9aFEoOCS/3IUvAdwQ1JF/Pa9W
XqbIciwQVc6s3sKQNFsGmaIZrL0iuW2bzfVo0AXRRw9b+h4wSvQWmYS8Jk9hhhkG
3/os1cRuZoa98xE7paa2WVkAExTrJvR4ieprHuifo28Uf2OPdYv0p0ZByOCmfmOQ
XUdmq/wDhnBWrtgTyxZNkPz+dksrwR/SJavzdKSESvpWdotUrxHp0wLA5rWqxzEP
7O6slaHdfZQiLeYZXOdrQNLnBPdhzJVBO4CXi0UL9ZsUAMrsr0u46viBExypNPgA
s9iZPe6C4kY9Hr+fpvV583hyI04gEhDMtDoc91V/AKnWFtTkq+G1QYcsNmeHJPPr
yixNG2jWf+gD/gMwPwOgvddKpUCODQyP3u15IDYE9Tk992oRkisRCt+egZk8bNka
xDpRRvctv3HtMurtfJN6uOyqVEGTJevUeY+mKqYGZ9nZAJqze3yd88sKBCU4WWmV
VFrB8XLo4sYqUbPUAKqRuhZWigSmd3vp59hAbLhygrCTN4yf2lxusFotBun2Vq0N
vQVeHbpsJ2R+IFnfWULhshX8p0qtVdHcOz4MK9Z+IvXlflE2f40bGAmumtftiwRR
R0mF5HL8baiG0/3pMgyas28iVL8PJkkzPJzcUchpLdtStvUnSO+1kRO335yBJL26
A80+foV+9Au8vwCTsJLC8bzxZbf75QhTOayYG5XFW7OmUjitNhKwZeukJHo3NbNJ
4Ay6ocNMc11xXR3OyXzd801Bp4iHrjBLLRc8JgfKtmxViwLCpdrMsW07nlevwhWD
Yz38xtg8akzWRQ/SdWp43tVoKJxzdCydIbttuU5B5Bp4NW+wy62SkfrUwEOYOVYc
ueQh5SaB0PBraCRoo3YmegrZQg6HGoiHJ7N50G/suwjzLkxguoe8uaPz7G29OrwY
8hBXBD1sSUdajS/MsnhsRXBgDW+tKYR/ejLOV++kl3oRo2W7OaGKH0Mx6ehNS2lp
jeCgRhDbV6e/wuYJu3/mZwvWeswlDn8okdKdzQlToCf1HrIoAhSTXwHNRFvBtcsl
qy8X7SfCktA13sjkhde1k76jdWpI9t/hrHffe44Z0u4enhy0uum5553UIOJPX+C/
wwNg6WtqPdtlRKAAZweEHoAo0GiIvkoMGQfc251WqU5msGv9EnjdTDL9/t2IJST3
/ZJdILl+0AbVUvpCK3+5zVs+NBWl4oqtLLBqv3Vwh4NwVihx7WCCcyLquHntPrS6
G0QW+ohYp8dcvbkDBPxbiOGNC0wT4cVW3/8brkL+haXVW92MO5qbPBm7Q4lw2UdM
0DHfRi6Vfj0CymEW21jD3VFqYnWFp8+LQX9B+SW6eCGePMV/sRyg/BurX2pvPOx2
/BWD8cqekt/lfJnTaxswc9A+pO02t0XUskzwTDXJ7/0UaIV6VpbpUYximwF/n75u
uWHsQBXQ1rv3ngHfMrr7qLDF233TKT1s1PEzEvJ+Fl5P0XzNEWCBrGEcoWDtqeZf
0Uqwk8avoYisE4i4TC6IQbzNcJeVD4BOH43rtX4n3cveSIyyBdRbty2ohGZLC4JJ
rsLjKPHO1gu8vyyZZGlrlRVEEo6D3Hc7Tr3T5EJGhIs9kqsxhDl3NmuW7l9CMHGQ
eJTkSjViV4W/mPCoaAMvOmcgVRKEiUVoXZo5nOgUqwVpRXRrObGmr7zs8lOddJFh
bhsIA7XRgWuzpQy45DA6zpsSo6lZbVVdevFlfhV2c4+oYfVeZY3CocqX7Zs6AG5x
w72gp/IxyvcDZ38wjcy/SdYpM4XlyiSCIce5CMw8LOCeQElH2irHALYgI/Zif71s
4DSf5q617kSmLzStTReZfNgeIKPyd5vyOqKgx2sUWFZxK5habFcLswJZBWFPUtSe
slk93h5R6yLK12PlcJio/dRCK8EZNzNBqW4+gWD2J7IpnYe1Z97KJIYAxKVA7yzj
WHCJKCicLxj/lptww+2ZpBJ/Dd7MSx6V9eK1L8zCkIzf7jVhM4IwkUT3sNHZfSxs
inFHGmPDNI/xgI+G2EyKUP+10hnhQ/oPbSfr6mywBQdqtOn94PVZU7M1I3P658X/
xUZxPP8vY55OTlxByUArNrbcFw9xdqv5BtujbG6BRY1YIuTPvvDD8ZlhhjmFHW7X
Kw7svfyU6AItyAN9uYSiZWFWBJXOHhF6Nx6x1dwxaU6V2ttcPkoQm56CZNAY4MbB
SPHp9Cam7pu7roGp0rLGsIAzwCFQc8rAw7j8PyvZdiVkiHNIPfV8/3HPW9nrXMSs
J/wGTzCBt4n3NVNzgpUHM1REqNVNaOvI52rKfnEe3pGfWtW8Tn0cJpEAvlwNi+l6
f+zHFSsVJlqgDzWNooKMzVXsuDZKJlBVv9MDNzjv7rvMOplBVnpQ9Yy+9u7vvEig
pXsz05tRm2+yQZl5C+gZ+jYWCfXDlKingeEKE0ubvXQXtIRMnurYSwL87eyEQYqS
zM3BbbczBI9agKfKUEtSPCQgYeUrQZpoJ1UNKy6ZOMmyVYO0mehdDFPFuyWdeH33
8iSFO1rZMNVFEi962nnBoaeyirvcMz+tUJRnrL61B5Na9IL9YJduYraNFwstMZbj
I5TOZ9XzK3RD22Z1TEYw/TaUZ5hB7Sh/Db7J52q5VFcRmH6mAIfNq03JhEvzvZj3
7uDB2C+xji4vDrccr4kBn1evNfRYinp3I4rmEuyckpQtkcdLYhH5U0OGpv0BVfnc
RH9qWV2yWEcdtfstEGkIlUGZREupty6Nd2YHbSzJuylSnpKqpNQe208XSIaN4Hfk
rbEDlcPOHhi7Ed///zbioV8fnXgINtaseH9ii+pm3Sp6rml+JXCQVS6xk0mwt/4z
tvibWxewBVi2F7GB9/TO59o6RcX/CyoPlpxUFfC+o3uBnxH8yeRjhKvUCJKuB7iJ
NaJKl9AetISJ4Y3ok8uzn34lGxsPRl0lMx3XM1qR69TBjN8cKG0yx+DTv1D/8DKE
aQq4TtPEnFY00P4vp0oy2MaAWo/6HyCGaDqCvCDmmmSZPzYJEMuAnVl+a5uh0S+F
3NBR64BMbKwayKPKsXnxI0y/EKhD0FAkiuqRrvBtVeKH7vyv3JVDtoNySYvy6wR/
+Aw2y/5LJdfit6tDRFEm9xU55hw7xd2oPt5T2JPvUYibkMTg4kejDSz8jXDP/Mw4
mDqvQaM5dx9LYiIOYZU645iu6EWFIfSW3m27+dkfKE//ZrA8E10aCmF9KEaIt+yx
5ltwg/z4x4shw79D0EUCtFaLx1tC7Oipr8oml77DITHQNYPTbe4oEK1h0ruyLbIZ
ga4CrdTb4wJtYN/315yBih1xy137Hk+bSbOcuSpMjaoxRISl6IVf/cwXx2sQShnv
G20sGKb8zQVUHB6nr4LSyIU0kx5HRzqw3AvXX9WHe5hwlGdBvwDWUyvuRZ3ldWz9
rLbHt+D35h3aiU0qs2Xgr3GQoTOFqaKmmeZhVCJgKFAT5jj5WTMwiSrJhwDlWg1F
oaIKvYAykMWwzGTL34d1tonkm2GPKviWaIKHcVQ7FWcTwMzcGc91X8SLDqf3Mm/C
SafK/01pbdMx+M0ul8seQ+X4H9j7EHs48OTAbTXuzdm+rd54vpuKmsPE7B9CS1RB
v4L/FkOIJLLDEh42OqsjMh5HRsycZ+/O/fcM3zHA/PZxXCMUfS3/auD6wcAFCORq
M0IQp1KymDSGrZ4PQztwwt4bpzZ6MMW6ek+KMgD75J7/XdHHUWDBiO9Zg+6r3VrL
+8BJOe33nikpGj1dAS5OCBbwFzhpHWcrp6JO61sCTKmEBHE5F9gbSbdS+22dX8Ae
7PkwIzpiZuQAMgZizCT/M/0zPDlJLLHfohYNh+FToj52phhphoiNTjD9MsM6XHqj
So02l8d9WzBcX1417enejT/pKHifpsnZiP8xefvB3Y7rLu+ZtR5N22RsJrgFoH0L
zzBsBdieKYrhLgYz+hZThtmR9cE4SmBcnQAip0xziwg63/g0EhSq03XkSRPNxo3e
1nHH5GbA3p+EwiuUQKld/d4Cxl0+le0Ow32jncH9EPyH5sdvkJ5VQWo/HnisK8SB
YXd/iyZDHc9KTkyQKnT7xlzzbOScTkbqL3TJD2JiT7ejmf53sakvaNmA/bdxmsBB
t6BSgG08nxaJJIUqY0iR+5Z5q+UGntigsPNI9coBGL5HxEMxzgWPgLiOlsr+OiBE
Nx8hp9jOwuoiOw3mNZzyvcL6qD2Ej6keMLsB0XexGSLHLCa9ozrBqMEMj/O5BAyG
IwWur828O/Jn8zOSralKexxCSDvRVop+gFeqg2woIOo5N3FM8bexirO9xoBBk6iX
dOMvpTMRWLZYl6f9oYQqwMYyPq/TZOZH9jPi+sswWtNDUAeMv7FqtpJ211Xj79Pv
Jx670d0eHDL8CWplmvBeAK4MbkptIjGnPJtb4EY3P/EEFzZoVjuNZd4NZGTKMKjo
OdoUhvSj6RxpeeU7gz3S1mg/kYeGL8mEV5T8j5cK5kidCRsBjjUhgun9aIKx7yP1
sK+h73Aq2EsLEGNfRWkRrlE+8Jwo+Xp8YNCipRnEEfcTVS0VUUIT3wlaiV4K95lw
jYcEPtRxZyeKs2DJ0cK6Bu1NUaDjr4Qb/K+EkmWy9YtINJ/vjs1qdcqHvJwcXexn
4Jj0RHFALiMDs9WnJamNSl7D2+EP4lYDm5FW+JZfDf4lGAHqC65OMgjIsyKV3h87
bklHEPqEsysHwlvAs/l47Ek1tWaC59GfoHKt5pEZNdWrxJYodyZugkE5+fgB66ly
taCJAOVpBtZi75RBdrA/H/N7hCEIvcXdtVcRP0y54Kv3N4B6V/9ymGE/5wmgZqef
JT/FpEO7/ZkwUGuLH0QjldYSVleDuLHgzzbm6aDWE00y3qe5ih0h9FGD6XcOLJdS
RMu6bEsBwvCiFbQ+lP2QbuQX/kdWP2zC6u6PgsFKAmF4eVmck2PpQmOBgaiTyeJd
9n0SholksHDIUIGE9qMCZQrUVXgITCCOAXahBBi5721GPxuHSSBrriioaXKDBMxP
6X4R0bXKlxV2oBsHOtOZUsOhVbgn2HRhiBUQ8aRY4SVdh7YzCappKge1lDoP4yfb
MbdMo1+nCjYESHOK7ZwEZKqEC9qgJ/6aFWHRxAKugAP2phrroTcJRyfzYHu1aBqF
cULPCGjJGtYNFhThuvAIXVJwiCMtnKD2oArZfKHZUM4qVG5HZe0QkpVn/M29230t
16wtXYzEg9j4GGFFDxFrijMxFvCYzCNyCdNeNgDcqCQJpWSD+oWqBI+Bjw2CbXcS
jCGimgcRP5mxHZkWFlAg/Tme2GNL/2rko2KqtawdpsgHb3EEh678Dpm7DrAXVwax
771PqEic7UGFVdKcRD1a+rK+USiYQvmJwdYJz67TOpbb/r8GrnuF3ChmIjHZOXNw
2mdF9BVXkUjTGLCyLto5x+3PnJcUeIbnq7o/Lk2ggzIgCtsm8xWsd7HZFKUQgRxx
o5w2Dc3k1YodmxgCrr1kNd3AsO3cD1pOuKVCN4HciOk/tkCW11cWbnKS0sUCdwIJ
9uUk45QlB1Zd/RHKUkgnB8vpx3XuTMuJkLXsTs5IYqCiAzi3s2x8FuxfA1f87ULG
2Mi/wJ7awBaxeKpNKMOAAgqh3ia0jx1glYh+dgt9c5mSL2qxc1hfWH03rKdmVO4g
u9nfgkcIMe9plA49DGaa3PP8MFv911HJG9ZQEgHaESME3b5KAET/S5zVd1Z5xqb/
/NywexJ3lbsku6JerMH4XcB4wKCYj7mHR43JYchcHR3VRcVZIxqNtNK9wbCKI6Mh
mSA1D2ycioby3eBJGgfrUIyNJVCUNBBxiKsBDMCp9wWBHz2Ddd39VQRXsWBSVLq8
1krhT8Q6l6fHkdYt34Zb3yZt5puICs3h3V0l60mmWAWtGFZHuInaZzDqKCzfruu7
R31699IWI73ibsvQKpijXdz4xW+S5JkXk5WxD7+KRbQGjFGOgfEKJXTEUraZM8e6
RU4ReZVemWipoRPqP6rVTt0W8iEWBECR7xxq+HcXyuEQcLCb7/GK81EBoBglx84C
IBH9IydCEJDilSI0Qi/iusWbvwzuBl3B0QpeJ3tG6viDdc3FebAC+37Z6XKB1GPX
VScqUMkVZaZIo+Dbr2I3uMvFc/95s0gvrvxBEIu6VmMrNbx675KbD1uqREWSYmjm
IhQJ6AzRKCp/bbB//oM24qWLfTLudqxK7fzUfs6kHa8EYsopla21eGZq02KyierY
O2QsHmOBw94L36slQ0TmAcC+vZMfalQDJEtDzV8RBWwyzgpbqujhsDPjeghETIj6
kKlB5MIVk+mTQERTHqihGFToRKJcYdefJgcp8gAjLYMfyw1m0RpaZg1Ssb+eob48
IeRSDHFsc+vJdLrY7mzOOJr5imCs5zsvk6uidJEv5dDPuHIPKoMBE2bSloH59GvG
Grco5NzHUTwizM7DBXBI5H75IXJemIiuPCvZywAP3qQIXpHBM+z6i68r3Q07v6nR
OjlnwnmAt7h8s+Q9yjwkAXmLKuxrIDJvXsB/9fS2fGeH5Q1is3n7MIdSXEUqM7El
BdJyDYi1E8PVh1gs2wM+yBwIOsCDpbK1eZ/TedRqvT4PMPByA9eitrBDc9BTpERx
YtEmV3ilCgSYv/lUP4ds5oLa2+2Kox7ERjB8YJPFcE5v7NU2nJ5RJEGg/09p86QU
j3vOPaF8n/A5Iy4/Xdi5eFcmbc+lepcAnf9uO5lOL8T7JjHME/Vsyf+7li3YnpDn
afJ2qVPI2bx/iMZHLvfieLGf0vcOnjd1jYBRT9ltkf7JRYayVg+PQs4r2veotv3M
s31zfnMNgyWVW7V+90bBvvOITwuTREu9bOLuPiCDudSpikaOypqWZ/ffK7UxWzAU
wMcj53Fb9O6T4kknsmi2oX1votjxQAskiaWa8w7gLPzX/YRxHs/turyt/CRPVdDR
QIEDksyC4jdi1A0N8BB1SoSPV+/o3dDE386d7tOsGT8wXkJL9CCf5xFzToLk0NCi
kPVI7+la82MDZ8mCbKLkBcNaPwXYm9rG2hrbgvYWcIsWUF+FRmSpQ++atl+y1wQf
g8XudXLR+56Wg8KI4JonC48gE+VWwx1LU5o+pq47cs8m4DLu3xS34C3hNYRdyYx3
WSv+LNyUa4r5HWQLzXJI9CoeeLrNXJZbB8R2csVbOYEYarTipk8PstGcZmBQMNDA
uQeVzzx+UY1Mf4paF4ZiiFYYfiZO61lP5ac53QswgmaiQN2I0jymnnSurys9uSwL
xQUt8YwDrZIFl41OBA17KMW1bCQ3W/R8EZjZA1mnPE6hW9ZAGBq7zGcWXny0Vvsh
ub48yrnxbsxCQPIn/369CzaYK5tMrcH4WCZvJ5LlbU9EBVB42p//YJlNQG2lBYPW
RR/YudEiLC4xDjcAIExnM/3hHLl21KkwR+cizwmRGhq0tI4Wz5Xm/7K0YbOfmNPI
Rq9A7883Yt2dhmFRW7h+HEMypBeRSoGkd/lcwT9J7gAA6oX5CVn03PNZ/L14Ay0m
VPiUw52FCIks5vdbsAqeWDPeBArSq65+GVEJMb0VMHAfCYNQ61p9xbjKYLwwhing
FBOnoZ8IwSJN/DFgmxfp3ZfRWZY2kaRsTqged6LNZC6FiIEe82QJAtD4vSdWB6+E
RXFYfdaFkS0qiLkIpneMMZVluC3TDktL8sHtowJCeVp5PdVKjA7chUWRxuKZNWS0
cdog7SjVhNiIDWo3Gfm1qrco2RVQuyo7Wv012gxjLdobh20x24sCQr3MLmx0DIBb
nHe7lQNrefRHv6AHzftml3uRmGFudPKVV0LqQWpmjI7+rxKFo8AbBPUhQh9T/Gqv
f06HzDLD3K4Brw3r7MxNrmhCbYj9ADgWx1xF2NXD7jzA08rBYUiYnjEqpFJAinnj
dnTiuWV1L3nH/O/+0SQ7pRZjQRLlTCNsP7yRYL3kDePLGM0X1JfwSW0TsgCeGFo5
h6Bi6u0K/MCy7+gwkcPX6sbqTF1G2zjtZZBSj9CRPTUku2CKRDrps/gzr5WBZGva
nj9P1h5PQaGctVzGW1+UTSuRBJIR38bKrnljgg4l4bsrP2rr7xRI/qPFHjw+Y3W2
cM+yRygzvUr/hlCVnJv2mG/SmX89vbAuuYJMk7EtdctezcUO9zcbrmP58Kwdd9kn
8BOV1X6Uo6xaJ97CAZS8oFC+uqeTYBipt7Q8JuqbNY6byMHznSyOLLs092FHiR9k
0sSvJMvtnFg1nTodOY8tpjEpXKN1o4kMl0a+Rh34qIK5V2A0CQ4nJDHb1CfyXFiH
Eq2+bAhFi46sW8z7w0geVuzw3z7Jk93ngxL3FU3FqFpTEiEdA6oip5iO5DFgKQD7
fu+uMXlG6wIo0Y9VW2RJDB/WzYgqtzyhwf+1LKW3/PK5ZlMjbZnLNKTMtSFSEZ+p
t8uF04fhtDPoPFTJINZULOZGFVqlJygYWIJWtEhMu7nfoIxFNJI8OSJBAYZ3ImOd
4y0bpTY+WBExGRj32LyaP6IKJCNP2DcPNv6gX0+YotYQXEG+IhpQCPaB7ngNYnrN
VFpUDksXBayLpcN+fKNv5ExlBzJYnJfIqzeWlr4IrSLNwD0WZV4Y5c3E+9Vo3uNn
GsWXX+YwVQxmm/Q6bgxV1Q70tDzxpEFDUpBCCqM5SPvsQ7GTchcgJc/C/enI9uAC
F3nH8kVr1Q7lQUImGV0qcQlJIaB9gm8AsHT7EwTIAvJ5vo7ps81Z1D0Ll3HCVOoP
a+cuQuZ03SsQHk8/lrwLub9qPv38EXkne02D1CuaNfUdpZelGmoOCENnf/A5SmRp
xAWVWG524CtQQpZ/TsidsUKqS82LZw8UilDroa0Vje5PeqDLUzGrZZeMLmNIlLUL
Sv25ueVXRUXARM0XOXSrpu/flr2fCFsqvDU6+iIt+Jit8Rug0f3I7UbePpVOKAEM
Mms5dA9EvHWw/K3/6x1ToQx3HQUcvMkqEJIskJUkUv9HRaT4cEYLBChM0+p90cpV
/KL+pqrl4V3iGkibzqWwGDETwfFfhHe3tTQI/O8+d8P7wR68FXEVoPFCj/rL8Y7a
ssMZpKNxsFjfapZzNRmMFV9cz9c8L4H1YpLKP8u3FBkdPNfRN7snrzIZmKsGv38b
tk1XLctmzJJ7SKqnOAPCzf12bZBUGuExZGtKsEERq4jN6+Qka/3WM6xg6hDLUmBN
EtPvVjDL55sWCcjCE9InTOmSazPIuiuQNl9HH0Uqe6g837cB9X1Wx1JpD6TrfgNt
TlalMsojC+lYbVcPrzTZHAucVfJWGtW9bEhzCwhZLsJWe9RiYuGY8pnimt1lyWyO
lGT/YACBSz3UW36NBJa0ZCrLODWE5DG442wFOxLvnAc0jz75Ca8qAiDwbdFfHqI9
AbNsl1hJSobAZr+R4SDz+UNWVE0g1pAggVX/Upow6SyNdZTEh4v8PBBSdSg+byA3
Uw4y97Hh9/O0SXmpbmTVws7hZEPhPDTJfUChqCOLLcAOIKNyU3nFJ1fs7AjRjTXa
CfWKKuCkV2MDLeZZthRV0um5G7bgFTveFOlYFe+yauApLUYchSmIvaXl1Wy1MW2E
lvNgcwWm9qAFW75ppIENxLGNXLJ1RasVNgJPP1WDqHInX7oOkNT611eJTzG66MRq
HGDphXilm/IsVEEt/BA5HIOHp/o53BJMXDgB7y4E3MoBYRwIABrZseSoeF/CTJSp
FzPJBvsfjWb7tKwve6xLjnhfzlsU/SyOSTPHS+IXGvVTbVVQOWXEGRnX3d3+RFDu
g5lW44CDxN2kNUHmmq4G/7C2lsDfXAjV6xDzWoOfRVjAElYXfzSprL96ryPv+pOe
uxaOFOCIT+BdORdkuC83iGpIip9IPnpzyY7PCXD8RzBmOjzCp9XrmZYpUvnkAWTx
/mF/V8gpI2SbkSYaSIxvm9iqydIGzQw6cRxeTEt25zNJQRGBFACNLXFwrHCCg1Jt
z6K66LtYBzvBp60K/BkuaxeH76/VsOiaGft0xjosKlHLWo1U0gAA+tJ9xlWIwSeg
X+a5ZLg7ocbSheCrF921mXjg8xKnvyfEgnCPs4URE9tKaXQKgDF1XIrRapSehkpj
XaS8x849+8yn1+NqwWtC1f4cq0tzTtgtSflsV7zAP6nuNf0UyLP0dGh32vZpH0Rw
xNmKr1CuNVFyXaTlbDrI4u9ch4rnDdPN3NWRNseExK4E6Z3qmraSRAi+737lpxPh
tCqcO1LaGsrqp/nGWLea5BY4tb2YrmsO6koBdsWz1WrFMqw1QO9/27s7LRPND7b7
O6pRzAdyUon/yeTS1xuOGs7V6Bh5mwZ0zeUCkvnnQJ0O7BPzjGz8ABe0bGBu5HrG
ayeqI029gzu3UpZVxKdZlS6ng2wla/+tRDX3jAmAQgm0469LceP+TlwiE7+Ub001
yxCEq/RrrF0mlfd6jXTNSb7hW4mV2OIRYx7mZU/cY7OUIxQKl24zHkJ/bG6Sus8z
jzRN8RqYY/AP7Eyo0aB7DqINDxStGr9HT9S1z5S22/hR6N5EpEz9qdTV6c2/RT26
HU0DMMfLA7yvflbb3ZvrCNSGtERRVSi/ZacZ/L7JEP/quXRI7WJwpLV3PO9j3c3n
fai0AnhGyzu92LTvnCPxSomNb9t5oDNHw5JbPpyknZB2Pqde/prt7xV3ATKbxLoA
SXndN90Su7wCk+GZzRGMcrSG54PTEI9QGqxboJKgnspdWvm3BU8lVzmZlz1WIkk7
taicJ8CROayGCCsZ3Dh8gt9uk00M9oJhOmHYFTu1qen7VNOA4I29PAM9/RzXAyrV
XONd/febkQjXGoPL1Ss3LJd4uDzKobnixXkiFkRvbgX9tUWIRaMI63ofPPDM7/e1
799LJcTX8x5pvktv3r7l9k1zRCHODVHCjFTwxlng8YrQmuiO0B4clr6LkOcC+6mI
lHE8PChGfHfXU0yuDjft98zvvb2QgI7CyRb9AA0l8e+C3VQEH+aKn5znStVWtWdi
LcFyH1RTpOm5YYX6lXO8ULDSvu5o5zXAomHt/7s5pBOW1W2PreyEchjGDtX55eI5
woAUn68hZAOtQS8lfgL/Z/5LGobpo7tUZHTGVJRT24Sv+gzFoIerbKwS6sVxYfpU
8TO9znEwXn2b6wJYSmCNDyGy7tcPx/aU1a29pVZi1V2mUShH6UGLANK0no+DXi1Z
yuS8j6e2pZwoNppX24nRsEXZ8P4NM3noStPa0RcuTuKkswOIhsi5eU+Q/r4Dnexb
AZq6tnSooJm4nV27sDzVY1YqB2wxe9Hjsdnj6/dIvGNJNKGWYsdVjETJFQR7Ztec
vkma9IXRHjPIanxlY5hQJEu6vJTF//H4x/fCkXTnxu0Yv85OpXVMEZ1TtHzpvKWq
tYWFThshPxWe1I+lUKG7S3dyZsldPpCDTByyKmyH0NxEz+TBS5I88CMxRDcx6QTq
MxPymabR6ZqiBSB7evRpbIXQm4c9qSbHB0vSIth7C1KudQRPsiNM09Qshp6ujhZU
QjDViSpo1hefSi7cPa05plVuOgFYgVYfIrk94DSCNthutXE6E7P0l3ixAjdgkSca
8fopoJ9IWi7HQ5e+UGpxmzwv7ZPyLhzvsINh5iWIUsF6UzlMCVcb9y/b/RF+1qfd
4xYVz+zWrUFgScoNVx1BFPL/0Aah8HDtAWP5YyTXDsFTdBrrOkofdXxc7wifsLo0
cdFiq7++BfVX3YmoTTtMl6XY3hI4+NT4WHCPUQt2FzjNUxpTCKVhzb2QSJcY4iMI
G6xxOaLobdmvohx37DU9g81ssJqjTa9Bw3Pooqq6gx73l1SvN96nma1HYoEjiWJN
Jxx9c9duOiCmgQhs+7Mf1ctMgynzBXNKoTscMy31wr3r8PkOY1J4kcx5YEArOi0B
XT2rCaPIJu0AQXFHfDl2WSFXnPdKsK/69JX9k4FnfKiI9NpKL1V0W32JX04DqnTB
Bl/Ho3vctCtPdAfNe1nbX4cZ0+v8RKm63vIBc+gpSCMZk41fmTJ4Qd9sXuwUhvt/
9i1+7koGzmS/1PLoSWeL4hEczffudwvW1zwCnF7ekdHP2tTeUes+fprzSY9VuEcf
j2QrflW3VJl2C6YQZkcpSY8PyQnb5xYqGJYSwnM9cz1+16I5w+l2z3NQlYvzpKQ1
6OTyATCR9RvZHNKmraM3kgwUgdFyLCDKyo0OUqyKRCiRtvgdSa3b2rV1pIu5siHv
FJ1i7t7hYxSoI/udGc3Ynt8Xt04Jpy3zA0676/EXCrtnnGOl+nO/5+aZ3MjuVInr
iQ0Fst8RPJr/yXw/26tntTUQnks52dw6yCw7xg1nglHTYSqW1dE2I3q3cI6nL/CJ
hOuiKdLO/1Y76claxDvW/4x6JYh904jt7C5UuIYrqLpCf4CeF6skQNgUt/wuFy+W
eQx/2SekadouxTJwfQ3iA6QG0Ee+g9uoItUOAKaKSMD9E6Yezix/WOr+mj4A0Uuq
FglVF9+8dLNuoRrgwRfElwiMiNeWjSqf29yQ6SjqG7L+q7rFag333fp1YMaI6Jyu
aP4VJhrRZ1AVJZ07M3NsEX0lnUneQ81AWPC1LBkrF0mFYIufeQpnnUKNnAwmgAbG
QPIEjNOaUtyMZLQf1LfC47wGpjkkZBxtOduQyR1iUxluxmnd4ZgZdaJ5BGjZbqY8
OpNTVC+BxZHPz3JfnimA9jcvmUhi15Zh5BJODnDgu+6gWChKaOCrtyZOGptQx2eX
N9yGGAiS485KUJxkJOMM3XJN3GCrcwKc7A0tp0Dl/D0bAKm7uZHujzOTT+RNwK6s
5TaAh3rs7QG3Bh8Uk2Z5wU0iYtLNY9fCagPTs/fz+L6dTIM/ibkq1uL1rdIIiXlW
6fNd9wzouZFWdoD5gFkdnfoR1cgV29TcA+GYukvATko9jBaLVsfZC/MeC03L6Ywu
rH+ZlQVMxe5cbqBAXZLr8K3JvBCKrjI+H7QL8QjFC0td6rjNYKqYC+rbSR40RQ8n
d1AvMqY+RsmrIhjCOjBor9eiQ+Csu0JxrDfw3t6Q6OfoyyvNP/V0+ODWoSFgsuf7
PdKfSW76iN0b3QfKjFFQz5LwWjVJLOi2VBrd1jfytNrwz401foZVrEUa8BoFnHLd
ezThETNlT6DAIbiBf6S5/zBMh8bv8OZdXh+cfUfCHLX9EQls/9nQjtoShvzxzygk
K/nfmpPGxQtmDxebCUA5y4KuiO7WoXEXF5yu9VP5Sz/OxmBO0Mp8Xg77+aqM93Pr
VEUk5sD8z1FEkDfpssBxEchfQ9YhDhTSRM7f1tVOP5EZK+stlxdC4AV1yxYewjAm
JdoBk+jkx5Xni2tNy3HWAjC4/5SDup6JAVAFr0pFHbLnXDOY2kPFcqwKJc8YsrUR
dChaKO4IHZ8n19P8o7CWhbbGNxJgunGI/DqEpUmhnOyfwncwP8lIyKK1Tzz7VNtX
7Dz5I2PY2P5NRnIdtrFqHGADb5xGLXrRrcF/2LJK0oHcyOLt3oo2JFTOG4C2V3/z
PAQ7XS+hee5DQMnf38I+FZ0ziFLGk7V/bAFefe6kmWXDxFDE5zz1rXzFeVTaqWBw
t3hqcrewJVfpyQACeMeUV+TR9L15TFXMOz83/yTxubcFD42DYV8Tk9UsEicJyA0b
r1xD5yGAQpn1X6OnDqeVfwDtIrp30XTBiSxN6bHoDU7q64BXW+CY0ACwYp31igGa
jZ3oD2Ro5uotcw6o4/bzEAE/FarsIvcgC7uTQBi5hBBahxg/I6eT/jiFJ8lNlwYt
z3ztthHEBv51C2+HDuIodrt6EFPwlpMjVgr0tuPoKC0w+XQY1pE8h9buY09UeqwD
1z3i9IJCvJEvUOrWJ43rQLl+Qpo8QjdK2u0qqGBa2stVdK0owCXbJurAbUFfJ/yF
Oa8c/cl+q2Yw69vsl74zYcB6HiPsnknqMZITciui9xhc5o9n/tGWskOShtlZLF4Y
CkIYkLctDudN5qTvxUAYpOQFl+fh42bqtoMn4AwiJr9eSiGovZafqLffiShIzFyH
qwr7J2XjrCcryN+GDFk/lhlGd9wM+zTbw6hnMIFMNI3J6B+0t0hyT7dPjG8UgDvP
u2XUh5ahtmNhUlGTOYeyR/n8/sIy/jp2LuoRuZfxPQMip7A+9KIfJGnkJEPaXGnu
0l+PG1ZJNDUmPxAffecBvP98b9JLM5YrhoYi9i+cUE6WGgAOIoWRLLlhKzdIZ3J2
ou85BcY1BPo1gFCGU7umvlWvBwTUfz3ToIBwwSZ4aBtqFMJl1ieJjcxpmqwMad7q
YKXaY1Pj4WV8i22EeAoR/wF8z7rgi1yA+/Woevt933bqSTTiIqba0d/rv1Unc5lx
2rjBfQl1cipb3Zqi+Xi0/goSSwx077VMSgMpLPaG//84Pgezh8eI135lhW2qj1vH
Sx+CPwjQQaw9GAXz6j27Ie1x1954oOq3eTb5JF2G3ya8+jVCgJvEA1u5nFAZaA72
z1LGY9UCFUHinIxke/FonJkElEk4BypotRGY7Mi79psbg3w4TvIPQB+bFqTaEMfc
uoegdpMkxw+CYBotw1ebz4nkCWzHqydBQkVhccqYMbiODSTZmhA/nqaQBOCUnM6/
6Yp0pnoEc6l7ydeIlil7MMTctaIkezmwMNTuF2seS2ebdvMWPp+koCSVMtXQM8H/
YgarOQIlan+D/1qzJvRDcgMAFwwmtZzLPcYpHw5M+EDVawQK1d76bnhZa+TErSwI
GRY6Bae315BTljAgVlhXx9B6tOJ52HKIRcoDpGeGlsGu0RtwzEO1KHfFoRihdWLi
fOByjmhGciRyY/3lH+Q0iPTGWFIeixhaR0hbTaoIkI6dg8nl/sG58jjUtkxCi50s
OU8IC6JozCoZ5+nQd+d1BssRbRN3O4JifeshSqsHirvfiXujVT+u22k9jdnX2dAX
j7TzJ2G7sDezctNNyES9cg+nc1sI47y29HKPmCU2NwNOsMesVLK8JwZqDoV4GZJJ
B7HbNzG5PWglnToF6vBZq4nLNe3tzwL8p6QHetBJsVSwoYzMOcanKqYpcIMh6vrP
Kjdg2OwRg2XKZwOezTUnuo4POwrrWzdhEvyFUhsx8CT5wWjTRaOhDrCFJRfN1YNs
J+bEEOTBeE8qQ2CHYMnST+Wj/R9JYCsKj3UDPCyBbYhbi7Vy56ahc7rkHWQPHvpL
fGmVVrpXrnRWwVepf0EsQPoZvJyaBAxxIas3sr1UL67SD2XzoHvKreIgklKCKy9i
SJ9Znn7er5e9dUw+B3zJAUkvVJrHHcm/SxrC3DP/rzlJoj9w6eM2ICDveC4PrpmL
KczFlPz4k4erXM4XHAdy+njXWswF0vHGSRNjIY59Vc37X561GeoQqjpWk0Zp3Xen
Fcq5A0FBr+DzNP1tQ/YYbCkL8eBvlgvkYrGUt2m1BMMdWIt58iE0K/LO7XOZPZyM
xjGU1vuGBlMG2x8zRaCpVbcxiUk6jAP7te8025X31TwETsq8xwu0Q6vVvemzSfPX
ZNSSr8HNDkZcYfTFYDVxqefX0A9atfWiGcFsm9zQRM3/SATY6Vu/zNMtHfqsZiRD
UtJNLZEV2TScw48ZQquvbxHsNOUTQA9JhbYkatUUmSskiNCsmehTDuwnIYec0DqC
ZsLcr22NLAkYa9Pe+sWcU8B8zkaRLo8YFPb/Zvyh8Fz/U0JGyUG2FwO/N3kP03y7
h7gUpEtJKKSPfvd8NDEkGLnrdvNWd91q8DxZZOzqPPBYi8wnxtttRK3Ombx3UrBs
V1PWbrStvsBuoaVUSY6TQ13XCk/3ISRvJp3NGyjHgJNanA0wpG12oWH5PnqiThUd
UUawnpty3sfgIKcrzBhDQPVUYI4gkGs2qABRVYcuHsm7UKlHAAPtm3jOsaQMwtu3
R5EI8D6bhcnCY4TVRalUtOH++hp6vkH59b6KJPRGIDTz99ETf80a4rFqPB7wR+LU
jkiCz0iKcjf+T2KbjDPnxqeHSGrRzLBEApcSSMsS90Mmea/SCw0mRpjrgxWMYJ2F
8h4UKixgs5u4+nIWMNTX32zZzPQy7SQVW46KKUMmvL0DQVcSb72B+Ql4egnHQ0jt
TFEH/cPmjlUtVxZnm89LwDjS7OcThbzSveni+FqqGEaok9vr7mSoaIMqlQduCDs4
8eQoc7jPuAZdSycYydIEFcjw/JzyHhMhYB5sn9Jk8crN7tlpeEYxbPNe4XtdOKZJ
uYcAxH3CSTGzUcGEB9SSBGScIRB9jSmjFSoYS3u38OakPMA2Nblt+ZQhI/mWMaPt
zrr7rHgjnb6DIFkeztAikoiJuCfJrnfZjTnbwqNz5Uxif09DWLcRHQ20npVNpYAc
hCzpESWq0qp0SBX2x7ykZE3HMOdYaPSe+jhtEZfo/6GIKlIEmQKuMk3BqVIV30Fk
VKOIsiO3vXLAwTz0hW5uerz98jxcYF+bxh+3ouNZnWXHon49hMiFJz8q6SksU6hs
ygTkWTeD9LAe8Cws3mG3Qrb7pWVUoGOm/UvFzA74Byla5cI8KYP4Zr97Fm1n7suJ
XKQSgSqqvZqeUkcoBnpqOi6JliCoICbSO0+jFj9x8fZVOemwIaFYfdvdDk/4l3Ol
fIH0yK0eis4TDrZkFvygKjsodSCnR6QZczR0MOOd26mCp1ntZ/5ilXG3xF+OIO3J
77goQmsFD1cRyRmmfsljuXg1IbI79/n6g9mZhwc34ck0KvXwgstk8UYeKFEaDj+/
SWCbSPNQHkhTMtF2OEgb+Yp1H1ZieLdXNnHLO04U4J28iXa3V9nViLVOKIdP8GQa
LxR+UIYT8pyJLPcewztoJVe2mL03lEC8wFox7SQxl6kLbA+XB3Kq80R0PrDAhmPa
OdRUoQqXJNVcp783yh7lBhXvdDs1rWS5grKMWNXalf6WK03ypBfnLTRGJwx8ng+w
sa48t4lxEze26HIONFlDtqdJZ8viYREB4HxpeQ6mbgin+guGXm6gn4ZFHpPWwnp5
6lhg1XAOnBmv99DxjNwRDEK+pO/kGNNkFl2EbqwLwqJSCWfBynNZCEDdhFv8pbET
4o1XBK5psFqBM2XkkXZcE1BmDVJLeRGNvZrB4K7n3ZxAKxWCzDY9kBhX8XEbgc4Q
7beKvMApUZk9PkQyp/v5apMgYbz+Rmc+hV8oD3aslcmDmO72Zu23WPrOEzU/+oVD
iC8OReYw8Jt8GfAqd4ACUXW3jiWWiDE86Ae44PfDNkf/UBVIUAZYbTkQi5r30M55
R34F9A/qdFwHyQPo+I+ZXY6I3MgXDEn+FRbW917WRsLtZ+QjS2zT8ZnKGvJ+wj6l
YsJ73Q3XBXVC8Kp1CVZ5EeqaX4o8QMx7qHNaE1T0GkHM57i2y6osvaCHf1kVLyZP
9QobGke2+jYKzdZMhUaxvI5eyoQhLNl8wrJdev78EnEUtUOfUl1BrK1RGymEMgsq
bNeUpxRQGLUgOv8EiLbvlmKK7e2t0SdpRAYslJnqsUKvedny5cFsyTIz4Sd8esJc
G+4OoW4o6v7x1xIEl2yJJ5FgkA3KYyuVCZD1mHbWBHxO0khO7gSSxTwg+eBcSh6m
1i7XMAzK+At3ru2NEFu7VFDd7jqRHrAWeJRnIp9ounKatCUg8aaRQ981ukHhZQ4V
/kK6Z//qXQvGdaqtk0DNekeaV9Lrsm3OYOE20mi5TBUvOjRifjtgsYStiQD1BKVw
JLUEwd09lHXgaZEeRTIZ9aA2ausXHHyoy4umFVIiYi4fLj+TOzROGyVCmHt8RdgZ
alZCJ8EB/oJvyrCMmwCVMz6xvweg+da4Jow3ZrWdLYtL+rta3EZohMMA9QDv8Snl
7/hu5A2LnT+g9hRN2IdH1NC70b/tUOFHulqq+QjLbh+JJByA6zJCF8QYCSWmYXdE
g48ZELpvEvHZgGxYQMYx640B3UUt5o7wBrd6B7wk+H1pdKf/xFk953h2lTJaILln
DThe/AkedZ04hHN1dZVnfa7TnGWL7CVxqXO0WKdq2jVnXBYzjhqkSLh9drRrF4kP
5DC/lpiJSF3uM1ucJjZ82QKdKAQOvgytpm2tjci9TEymy6Q9fHEEHW0lRHvWK0qD
RiFkbLdKVwWmf15u5Uq3V1NCIWQeSLqaK5ho/1v6tqNvw2iwSxxKkYXNyfYA64BP
8XU3+ich7vpcpS+EFO4ca0gzEGldp4ad1DuDKvcPCuBxBVW4vfhnxbVBahZdDpLi
uB+YEKzeW5CEGj82v3t+xZeqaTYt6/P0T8bVz/xraylbCpnS/modNOhm6M1Au5Wr
bc31RtONKFVQxuzC7Qd0UrP/5mj42/MNLkT8PGjOY4C8MABwMNps8fbViM0wVlhg
wvS3GxZEWH2Ejl/y1IYW+5RZCGyePWm9BH3OFWM3JoZbWx2qb1UXcZUNxX0rHRZq
GnpcZn/GJ8KOiOj4pBjpjwFV8TDa9E3sY4iIKp+qGYnc3IVvzvS4g9PUJfxdtK/S
I7WuEpuXyGhLR0m555CpNzDWURwJyj1p0YiR+FYPb10Pruuej6nuambuf+/VNkCM
Mzg80IKk3IfVw5phhAiTPft9xgMYRJsogBJ1rJOkP03xhgEC6BqiKrQ9btTa2dFj
ZIcK+ueQYhgED8J6Thtfyya/Y/8fuKcZZH5uGQ8PExKJpgM+Y+8k+HEUhqaTNkju
Djk6Jka7j4F3qNiFNhpUySQlTuBJ/pvfWmBkrgtttKG4mKFs73E3lyFIlvnT/lwP
2Nr+RwhRXNoIbCGZsde/uNaXGAWp/hYQGU1XhKa1EDOiwBWoKWsQyeDBxC7WZwWe
pGM15LHasn4fpT//mxO/2A9E8F8yZ2QcO1XLqPF2VDgIGa8oFrPzcdJl762XOS45
hEUlLvVWDMMBMzTh/cGEoci1Ys4AxPL65i72gsP7tmZplC4kpBng55suVOpqzVjD
gmJcQTp1gHB7z1uRTq8SYLhCYUMnkh4zif/ANOD5rN7EKnsRIzqrrNlvuT/gpDQF
XHNnfDQkjALGWGXvJQr6O1QvbNnHcv6X35GazcqmGpFpnVsltWzaqFa/JjOlU0M/
Cr9b+kDn+JJ+qEMWB3TcE9bREVpityj3pyolpplY0aSvSmDlVdAGBBWnEhvtYX84
dnGjonk2Pb5Z5G0LI8BBrEXyv/F9u9ovzGMZ1C9t4FY7ZPlFRAcnoxfE+MQMRGij
L0N3MDsc100ILXeA8jfZC0Gim1BYGvVCfe5yfirZ52949ih+1w8T8kbIGqo5wyaM
mfRaEVJRq27RcAB2wVlMj5+q/c2hkxVzdxQtq7EXpvi1zYqIluoZbR9f23MdwGtQ
SmsA50WPgrdWgRikzboxI+A1vAh8yz3GJQmDh7dfQFlyHpYn5Fe2SBCdsEjxpzXD
QZp5zOtkMiIqkFMmeKSUfwdVN+5L7tfXROcF3VmH7Q+cz/6sTuY6rXkOvLkoyrnM
2XfUWv24x7MVlVWv6ihnuO+bb/RmPMmenJyXQvPdc6uBOBTSYJkhWKpBQ2Ln+Z6Q
BEzuWS32eQX8QfUqpJslfGQ+TfwdvRorYLEMD8/hBNIwDOci9lNCGHFq6t43LD/w
WFyGKZBkVpBEvV69r1jfksTsOzshRA5jrMfkRexL1Mdmfh8pVJA21X07fcukB3u1
daXM0TFygU4R65DpgiDecimECKB3yj/L2yjyRwGYP7JDqG/DuH3sfBZHgNLGPuaR
aElFvaiVzR7Ph3CN4DRN9JwCeIRidfEjsjGRShhEFamLS4srCgnvjeU8/Voy5CrU
20vWbXGs4mSrDU7e9Sm+58ee5hICsZ9RNz3Oqq/HwLNi8lSmfkQDsyk1/M8yPv6s
e1MiTuUmfmgoRHPwqXcmlQPcZTZX0RQgC+sk4zyjZ1tBcCggO15DDefk7Nfk9lp3
jBDRe/AxfDj2yp+HqpmMKsseQEYBxRoq3vT/wbaG9N/lYg5uC8Tb5Da5pavm2dAR
KV4diLMrgOyZO6ulFDt6H0OuMp4XM5dGXu0+V4xSH6MH50mChomCGfkOc0pB5z3C
TmA4T9qPHItzW7hySq7KOuigYuGdXhIttbYhjzhWWBcma6NGXuJa+rACNFOa4Tgw
tFANSbTtGYd8sLiQjG5ZIYvYe29XLmady2Cy2zSUI+8t76oct1XiSh9gOlrNTOAU
H4yPmIkETfAG65YqBk7jBiNpMRQ2X5URiqpU+gZFx3/VzBIeIWFO/wC17UpcBL09
iy2DieXoWly7FZuejIDSFi4EHrWnt1EJ/Lv1K9Un25pZdbYZGIfz2ggfJPs5Begy
/6ibLlzcDcDqHkkKn0AySHS5Ylw5/ZGfeIWYcO2WvwmCcHgiZr16zBPqK4NDocIA
o2JVTf6S8sEoPrvj2kUxRtOrmHB8eP6WPq6X5BW5u92mMysiY1VohDB0qwcZ9RgQ
vzBo3jKIsEciIK+9xOce+olRHo53tH0j5eOtGkX2RsyZNKVELLYAYYR+PmPxq7dp
/xcJOPnX/LQYVYjEaWyd9tbZRSChOrRUVBnG1LAxTP2UqDhIy3c9vh4XVB6ttrTe
WGeIxQUAhbI1LaNOwaiCgzyzp+DODiumwIueZg+zqWB8yj9eAzNRk4n1wUw0NGmq
CcPBvNsBTxc9kaKsy+FD3grHM2HUunXt9SJXxrDe1JCFaQOn7UiUGSD0T40IGNBU
8nbvG8WGfBf9zCBQgARZCpOTXKfsgpL0lJom0LUcm3F9r0nmoAgOtxatPk7TfiiX
O7o0zADRTqCD27PJb5ElD525G3CfOAs39RnjZJPPVpcOxRW7R544zJznfdFch3nd
Bq6FA2pwaDV0sayYT361dLpXlYmm762bEQ6Pv1f7Dr3FPenMXeO8vGHrlzSvRqxi
2n9poPAAFbfIZrQI0PwYNcTqsVseA5nTUsGcJHtK6O5CDIu0WmVxWqqnfqiuooUW
3pTRwGChOf07jSiCfyfDXnvDcFblsyyj1CdBk3Obi0TA4phgbTt9TVCJTeQ68sW8
UOaPgBWCANDcZT6YcgftD2xsatIYgBpavNjLx5MkmVL2Wy6aBR+yKylFe6IRO7g0
Wm6Z4AFSYS2LMYpg1Sa+cULiDLhkcYs8ZcacaPuseBWKaaguET3+JKE/K+79yO4D
T+/36ANQEyMRziUQdDGZ/4aJpxsANiyghS8cXusaUalxdWajCXKmqhn0gClfR6Y+
9yL6IvpbEaBWCm4Dm9U6HXYe5HqHhK2zD2JE6UOyClhnZsTohXOCQsCaWA9PhVOu
RAEfIEsv4gcg0XIb/3VnrraSRwanz5gtZUQg9AELrsM0zJ53hXb7/vAgHTQ6tVyA
UWrnM/k+Dt5rf27c2JFH5n4EkKnpbVLLLIsI12UFwmoiPUGgiCV/Rj0NLn2p1+Yg
+BUN68kGGgbaGTrqDxvc5T7Z/hkjP76XCy/bWzfq21SAdG2OMC/E3x9C640MzTus
JYdiXOKU4k+JYlFDHXC5s7j78cInpg+OU5RFUp6sii+Iokk440NhsUaWW4U2qVPK
tORxYHi+EmZvD/Yp+ecAd3w0dyIqIr0jgRxvSBuougtXC7AvS4HoN2PIrOP+4LPC
2NxdIGXWxQ2oUs2hn51arv3Yk/xu9QpBA455AT6HD57U5VvxGYec+RxR59OIL9gp
RwbiTPjs4/Ww/JadsaGoe5vWAU6dpmdPLOPwrXNYzXBmvEyqKXXlQUVDQSt5fUfj
D63lFy6Ha8n1wMWuSkVNFuPkX6+qJ5GddClnhUFWL009Mq3jCg4/yHX3n676fa/u
L0ltSO5KV1t4BeQ9Gu7OeSZpzFz2EW/ClCXGhhsCAawpy465b8jUvLFEjkls2njV
EnCbfO+BnpZKbfioaw5tniL6kZJrCT06skdX7XL0hyv01kDpzfrGWABKqFbj3FCo
T+SjFI2lH35f/AWw6HIAUnRI5l7PYJn0Ps+rRmnwfeavOQUyuWF1CWGmSPFcN2+z
HmT5mBEuAGRaTmlzJ3qKQKTaHuyf3oBcaJwN91ADfYM8G9cDuigOTeuskpvGWdlX
KFFJqci8IZkKg8XOcu/ItNe1SfNC89lzFaJyUJDPmGxHjeuoa7FGszecQ8RaoaTm
zhI+PVcYdr1EBarymZiEAyEI8d106WIgyDZwVVG2b9fl4/DBwB7AbPzLQH/gH+Z9
eJ3VTGs6Tj9gKb3E2bli4gxP063Tc/XWYbm4yGxhmRVJG2MGvlSoD72InSqCghMu
bFI+Z3Cz9t6kN0GtdWro9MBssh9hs89OUU3UNQIB/KUj5AxbAF1NJO+C0r6KaL1L
WAq4/gfa8i9hVQwCj5E0LDojbHCJS4Ws01AEJ4sMsoyvliJ/InohzF8/eqFukcDd
l7GVd2UqlvLrK3cV43q4gvjxKiI1B85UVZVhBXRnyxP0Jvf1ZQzseNeSIgWFM/Lc
EDAqd6b+HoHTqn1W4gH4rfzjOAZ6iVMWEZpNzyMNhapA+GSLwZ6FHCGjy9VNnk48
lpht1FggiJfBv1Pdvu7ksJI8K7H3r3EOco6Cf0f0HeuqiVyTgac30JJtwB2iDbn8
VSNCDmlFtAWmxVBK6hOFQ9Ja0l0XT5cSJ7EmjJt+1b+XAPvfP9j4sxaohr7hgXbL
BPwW2ERjHn4goyGlHoJEtWvXU2vDXr6nLCuMAiqFpYmMHk26Z177XjmYaSZl5QgC
Xo6b+9GKaUibhXv/MOMnMM/SJ/EecYtu/nYnJykfDWrA5deww8AF+xk/xv6Vd9aW
r+PcXpxUu9E7XN+m1RmPGlcL2ouOpPNqrQy/QgXF+W1V/opCm4XRoqep9yOp4zbY
S/3Nuzjb7ZXCQ8iSfQZ6IphXwp6Rmxu9cpoMLc1OoJzqKT9cgMTaz5ccS/REONAs
Wg/ozP4xzrOlyGOo1Znu4GzsW0OCvjF9coWLOLH+Cpg553yz8W8ZttpUK59omsQo
HQoiBquT0tiWFQzYJz7obVstUyZPPqhvOkZNNA8N2ovByXNzmdfj3i/cZsj4ajp9
6rQdP7N71DQkTev8FHKCISqfRicZO1H6qoB8KmmQYq5A/FOqgaqKKpTzexeaTsUC
HAATTjJ/dvr/fi3GsCoBy/X515yEzmJbJeo1GuyDvPDjmWta5zpm34wPHcyduRio
Ewh8FOJt9sCdAwKSw2rce6s0tkirDbSv2AoxPOiYsME7JO8xNbZps6+lN9EhRMZ3
UZ++W/W89ypGUANDBHh5H/czbIzpE0fHSIVaZC1OZmt9tblrOlXXTEPeBiyP/rA7
4U1uWd+3o1MQokW7wyvEcyllgqVuPr0S++wRioVNoBcMI37AiO0iMwTDV0p4BJPC
PyFXiQCXOAJi7UIkutbWuo7Hz2F8Jnaj1N+zHdt69F1KD2kCGT+JUPiMelJkilcA
waivwxbvgRO1l7+BCI8yPZPH5qIs647y4K5UZV/t46I7LVAER0XoNDjRT/78l3Mi
pebtUwffpscuKIv9XRG+8rl4hAosMTOEhrpRFmGqV/iG/e+sWv3F1Bv3hgw2BjEH
aivLzMaJ2hwMWE9vr7+zHHTntK9DB8x8khbZHzPtXPkZual1ho1A0hyFPkPaNt8j
C5d1bI5kL5Yy5JKEws1wmJyK2H/R/s/fq/B7K79VJKMjWTSCSbDtI9Prsw9rwIa8
hCrAjJL08URsy2Jg6gV0+fZdq+xc7hXOmT6eApgDS5gX3OoxCrcULWpo4sEkyfGz
VUa9Wxom3w86gM5O720vR6cHpTuX6jIihmvMYb+p0vWY2wv9CiSmnkKSUrbah/8O
aVTnYvESVwCiwGETios6WMBCWJ2dkpFwkR9WV1KPzZktdXTlAylNhCvVHjEujSmy
WlmLwvZfLltv30m04E30qdRrsqhcPVXj4G//afe7OcY7JKM2u/X1dEHgsFAL3XLT
yhC18a4RlgLOTm9j+3wFhYOsZ6fRmJpGHhNkQfAgb/wZqTSUxT/fSXkSnzHb8WtV
kUyYCucZto0aKoRdzhUIOz7Sxuu3sDQ2BlQt3DH+h7gvkM6dGyfjqGdy0rh/w8Xu
JnqouF62j83npOIWDdYwevYYnRbJ6axHvxXA9TZGzBIuDPnCAmlQ3yfvMTvYXkKL
wX8NVSjAuL65Z0k4Fbi37x/lQdAj1jIO/aY9mVcAgNSyYwwoLxqOLXM3Re8qn0KR
MYMlP7QagZdvewi54Q3IZZuqoQRk3QPgcwo01njasBRkViz8jQy5f3x3hPf7U75U
8T8Mu+qIZnJ8psQAqjAySu6L6hdQEQfo+A/dccrB19+NgmsOZE6Mmche7p3Y66TK
d9u+BQUvtcxPIbWC5vTkC+57Oi88LB8Dk1xNYsHv8Yta1/YDUviYCl0Vshc2Wwh+
uZAty0ML06ulvjDJbtJEpQrYoogF0letd2zWVeDGSgotSWxDmqpLxQGqty+yNPj9
0dwpe950s5lIcStnxWCsKrT6D3twd0JSf+07ka9fbXjMPbHZQhq9OBoUqxsNSShO
PoISeZYxcjQBR6SDnIapgkq4mkqZ1gSvCLv8NThGoiCLaL7OvZVNvOpQesWmLEuI
/LewgMvCndYqFFWBa1I7kEFjk+OfjL6RbPnrCi6w3a2/wEg95+EV4zJH3fmtpYbE
oOZD6C4EnWzprwdTTEGYkwXN9ZMCD973IVliCo6heDqty8HihTL5SsptsW+8Nru7
ZI9O2YF9uCNAzsCSqXNaU6cEaWmjqrkki3Ml6risGRAfGwjpAYdZHKBo2B4MPoH8
W1p1npNGOxGa6PAFw207j0aXYsdBUxho3Jbk3Vj6s+vtl/B8RaaNlv5BjDDj4h8Y
UrYy149rhpxHmZq5ZRl5ee3nV+oeaS4UxKYIe1Q0u96sE1C9xnQxg+2kpmYA50Uq
vymfTyNCirBjlAgFnkDPRR55/DXXF7YuAOUvEeixJpMiZ29deaFHHCv5MilL2O4T
NRt7d4i8GruHvlL/c0oPHHL6fzBx/tHnC0rdEpjD8nr6TvzMCWLQb67V60jCoKuO
wLOtXDf8O9bDvFoQyrqBzh37b647wiOddadDardZwSNUiPN0cNUO15HFj0ocLOPN
xkA025GH77NzEcINdQgYOFpw4vBblgC6WVmYgbOgBSHFqHr3F5MNn8wOU0OLYYEq
SBKyBzWC3tNTIUGTVX0ODJOzCBGTwt6dLGan6LvXAqepbd6bRga0hkKNl453Lwv2
BrNZo+5IHhseA40M0Y+fzSJvXgRIZi5I1YCWzHxwNVc3z2cDzARH7zY+/jmz1CO1
tfkECEUTQZlpNw0ioq9rAn5vr44Kml4sD6EQTBlMYqEho+Knf2OpbOU4Z2TMGeur
SpDpQ7FiZ3j40vhb5oa2ypPN8W2SeB7HN63UgYDbEfI+fnrf3bdrBeJqyqKF2Oi8
F6KxfRv4dMq20WvHXBtg9ZxaPnIy+NTYd6i9EaT9jhlgb8MlPdHi4TmM9OFaW1Nl
i08zMoys/iytOqLktelLTOkTBMDfNAcA5eRhvaFBPoDGeqIs7e0YiesC6IUMP5Rs
AyelTHf/xMnskY3NJZJDw6BlmSA8xQ6xfqyWm0pYQ+SOI7EVQh6cKu+CjbFz1iaZ
foyq/de7tYIKa/nIB3jr1FsiaK8ibOtPkSda7kcVrefgMk38Cq/pup20849XdYug
fhaRJIlERdf9kI7AmuF9EJdqfe9SjQD953g7Ge6A9J7XlFxHN6b7HX54x3jegyCD
+45QHWEwI2K8488c51IFtjt1mBDeIXxg3sZLGl2/JlXIw4AYbFDERvvhzPN1Zx22
d/aU/uMSOy6hfE2WjUtVxG5DasI27QR3QL+2EBYKGrnfq2sPDLrlZbD83tZtRff6
qiKfm8LkgiWsPrZnzJ7jHxQIKeCmFOm1Fb5FX9GrQGVhGjdh2jOvCSPjESmCBxbs
AcQgoA/rwHuxR5JETZuhdCKQjue07j1hASLFMGtxAP+aOyBUFVJvQd78OEv8KT/2
Syk7gaseIX2/Frsv6u2BtjA4O7qQ0KCIfUwrZgJviPlUhn5zQdzRqgRrciH1Mvb7
FyF6hL/TvZPAtqH4GhPt9yirJe9JV6QUpW4WwQnAPyYUuPCsO8+wTl9momoBvQhK
b8oXv4WA3J26/2iPH3KjBCCFXDvKEwY7jRCI39pP35r8gUshQTsCvGAXFxW9op8L
wwlves3vVWzecIYo+a2IwYxkvKQJTV7vkGnjSzVCfdg/A5dbyw2PqNW4VVA8ACiF
2KnEVaTTjFxIJ+Zm8MzfuvpAzrLLY0tIp6/enAZ+IVCI5YUCQnZmpr913QFdQH4x
6ToTMb7UuKUdcC87BVWUgBy3EQFs5ZW20DZ2gKeX90087NGEFCandplXQAZeygxo
4Zl7sP4IVSbIp12pt4Dre7UpGpBiRydpA1sEDeHqW2qDOJPjQdZHQmYTQoC4H2KN
EIFiT5689VoG4Xa6IkCLtK1TuuYv84HpkhsSHMoZQLXfTyU+pi18E5KnLZGelony
JnXH5E6HT3cY9qyKYAanDBZNHPBJ33DcNBiAvEd24giUs3RGYIbccKpfZaMJrmJQ
BOO6iAmhUXdASmekLCBpgGq2MhJvZdm9CZJC5cB1uk2ZyViijTUAOWiHpKvDsC1C
+pSV8VxPcA6lgs+uLaqfY9RxhX+Lk4unpiss0bt6PGTkqUTzGTguUZ2DPRO6Wk4Z
T1KNff6KAerV0s1E4f2BhzKwHwIbwWyZSBqpqovkWHx6c+JS+V0Iym3ryJCBJQGz
MSvJ8WQ8J0dsyKSpmtKqlRdkJmvkAXpTuMjHL0nSWRcBkTXMEcnTHfAg5vJcK9iV
DlfwtirskJreL35QEFRA/n3C3XeATcpj03qNAohKrCjioJj4NpwBqsUP7b8mS7C7
Kxl7tt/Lpy4rJz/di474JHBE/QUiCtokbJVIK2CLETC0cPcS13ZAuSo41h0TfqCc
RZZTgL7StT8gkQXSCTSUWB8nObYuMYa04lieuOtEB/9o9MiDMQ7fuxZslNy7Qd+n
Wxw1ZUc2pCpo+ImGUAH40BEw3Xb1QFgBqhQ8TUeECZkd9AmGepEv/L9yIfxTZ3L4
A2DSyZIiV9feft+pkuu8+GBWTn29khcT6Hibe3s7e8KqEfihbu3n4hxFUGnA/luU
3wjW1wmlBfG3Gv6AshpoLdV54Ys3l9GpHpxtD34iYSDpgVsuT02I5PIuA/jBVKlG
gKaycWVmri4QiSDUksPLsMdEpxG3lIJW6YKP70xNPusigOZbBFDuKRXUUV1BD1O6
a1wnQMsU3gSbt7hI3iIVxQ7W4HMyIE7+mSc++5rMd7q5PWlQLG0j9TWpJqbC100U
R9q5FWwIfXtyGfN9Y/qMVGhrKSl5LabZtuzZM8K2TQx0Ph2RH7vsFuTe6KuGtZ/e
1JE/MSYeyPYBEXP2KviXQwE1FwrHBdTahL9jDZYq3S5GaEshLPpLeIWH9dyFaVjj
fyUX3t6jFRJzVlHAmBuS9nILvl5DnSm8df6MarWUdm8C2es+kqAB6xWBfXvLt0mv
ISdHGV76vxLOA6Rsid+8qAXFg1cGIX7WPrgQXe/B8vkrejeHhrELQemBOE50+TfF
KxR4HSr9tqsjNNjnpfjlYicR6/qMfTuFqOVe3TcGmxpUBRxvMoR5UzZGRjpyLiP/
rALkeUVCEH2Ld2XzcDLkigrP8D4SNaFWF25v5wjriQCOBN7MwYdAQYcu0xa8Znzz
AACb+mNoRW8xZ29SfnfOqi7YG6WwCpybrBAmgGPWgBLhdaEzhxlcUBqsGzKkhoD4
Z2mfhHOcao3nxNP4xR90oLuw7EJuh9dVc+nW/eqFZRa/WnrsUWSVToRBRj31lPsc
FGdFoD7xV9HBMSRTVnpf6iD78uTOLBU6H8fbliWLIFiaaR5AJl5ehFXcn5SMmZA9
u7ZQvRT0kDZ+I7fzndqkhZ6VJrWjUe7bPzUOV8zjLxSFfZrVLNfBlLc6oTPXHHTE
j6dO5aPQyR3V/LFs/B3eH+NNbWTmvXOM/WgfyTh5alrIXYUQzJd3d734GCX4M0VJ
jndjunWk7ewT9xgqjyPbczEt+a2jhblTHGNXHIa9l48ES5t4YeljzfTMzWCoROQF
aOyow7wx4HfhxosHWFuVZHbjv+Gy5Cuy0gTaQQBNbLfFVTy6ZYF9Y4pQGz1FZtGn
45UJnUgfpfwCFadKoLT5vDbZUgttKYA4KH4nSwlNW+PVhQtfRCNmU87BVCYn9quA
E/f+XsBZ4aAweXcgq7ZqbQjupJkgZiyGL4/X4LckH9spfg9zDlTHY74M+Ge16Ccu
cohkHGhlgLyrs2tGazOAMUT7Nx8ZxxdKqQksJKmR/vnFclBboiDJvSQbhEL4Yk0a
lhAeoAoyuA+cLuaKtsA9EGkLl3kbmwUdX4M/G7Hz7704lmicIPELVqRi0qOq9E2q
5RQExSxblsp9dR0d0u0pO7/fTU8u4drrXxWfqcfKxOlDRpKjg459DsYhcHD8tQE6
s8G3J97swVrGSQrqgV0XJ6NTemYoj3YwJv6W/CxjfGGRreIM8aEPVM3Tynma6M7m
E3C73RucwUiyOyv/RWV+o9yzgAuxlpdoCXHjXCsDhWdy7JsPg5ZEPN7aGlFaIA51
pEYIb/IH5xuXO/LW8JywdK4UVI8Rpdkwj8Gf7doNA9rBfkWOSqqk3DxqvakHkBIW
qYJlEO5k1GVxbAtt8L151Px9bituItEgOonNtRWi8mjTODTrC9z35m9g0rCJZzWS
9TR6ZQJT+r4GMCD49jzeJzlKcjxToG2/6liATcdb7lwyJD56fA5Nhvz2UpA8arou
8majyQW2tsmKiQFXcxyqFy83AXISNWKTR9Ws2pEuM6swGzsNNn3h81wGbQt5sLVs
Uv6KrY7/7Cr+1OL2C5lhEWhZXSv7YXsvjdJ2bOPK2uhfmVZCrF5KKcb2Lp04bfju
WC2JN6xLlN1G8+MHa6MKGDMkBI+WR2v6oXRrzBywwGQKLxdlT9DDfVf4wu4plNT7
hrvCdtJT3mxO2GQq+AQnCKQbH3zlGtXdNwmDsDe/c5VNeUa63+faGLeqvrTS+vbn
eX/8Pwu2G5/AMO8GA0wyBcuUcQOPcclNHZ3AJxByzaUVzIhMUIq9c9V6FfGxd2dJ
kAb26zSzKcW27bAk6pr5Olp4jVLQ69my+Rgg+khZ31o6jgtY4XKj4nDT9OCsc2QO
wPHZjCexerdlgUe3y7O2/+nasK+6b3IioOl8N72VALQBq+HtH7QcDy+goI/4N81c
pGdU6WINHC7u6G2MHhqqDrW/SgcbUyoblhpxAhsnqJsG0cbZIlje1fAIfF6qF6Gq
r0bVS2qjB+00QL/hJhVLm/XCv1L1xkagvsB6focrvsj2rZa6N2Eso64khFrGKxA1
dRMM/vUB3AHUWCUi9TRs7+iFKkqAW6u5UFm13aSgmgT7yku7ONB7e8urBKPRBQUz
QBpF5x4z1ZPwAvULj3XEja0UB0//h7G5alYtRIx3H5pnWZ0bjcJHSexqjLEXes0w
aELXDknZk2bV2FCTzlihoU24gcW/0AfHrw4xImfhn4uamIS14ijJ2PpSfWfOiMy9
dznUt2D/5Va1jJkAo0DH0JchzKRGFvhDuWWSWg8ceO6u0P4ZGw0ShQKxv/H5QZ8x
frKdzXgMkvgitNWnsKPAqmKAUhapztKbGMdDnMpqcdO24ktJA7N6giF3Dv7ItEre
lj2m8BWj9cN+M7qpBB++kbOEYzBSxXH/jIaW07ZVSPL/dEK7aYR4/pdTbKtxblsi
cz2TVdG42VQx1CjW8h8lBWVKsyV1MW1wZSlEzRfqfy7ngWKs+WmNVD0yNGfgRN6e
s66HayAiBBZoMrYye/OhvlFGVDeAbLXZfUqoAaWGuvFsKwZCXbQ3jJyk5JXl3jkI
l7a0VPUlD0RWbwwGImFtk6e76VfqY/A2WbYPdmkOAYsoCwyKD2tM09lpS9s8WgA/
Q8AmUIkxdS9omfelZbRo7I18ApLctnxHSwUfvXT/4OFMU+cepaQQoh+TsPMGmb8Q
0hUG07PBrtTBhL5e1bm/i8eVVGG4529swwp/uy0afOgzNTYW8+MOZKfDW8DiVBe3
eVxmx3UlRMxMAfv7xQk6acVqjCwVRu3Tb7oKJOoRofAzjB6ig5oE4fl9IY6o+1O5
dgYocfzuuTucG9bewBA9AG1o3BXWDUhBDlGEJhIX6Cl1rLY8X93Zqtw+2M1WeBk7
zV5dMPdjRE6X3fnvZfj7x+LKZ3QGr6HHcdDcA1JkrNXMA5mASvX26DcoUvndtaxe
JCYCI//fEc5rWOEBMRl9xUotFwCG5rXA091eRTyxBz/cINRIypGiICL1ESZJioMf
x1QjxyAHleO1ay/emwvyYPhcCmV9VEOrA/uEjA3FS03RMe8Qa8VD6rpeWrMaaloU
kWPSZ/5+VgnFTprTDsNZaNVDbUob+SiVocjfYcV1zvUtY5v1ff+ZSTMtANrRg3mb
tyCmpnjyExuJuNqYZ4twXwo8zxshD8SdSMD8IzabIbvVstPyRKeFatcCedO4lfE0
3slFAP02bnhfTi2IAT49HHZMqQgoDXg5goMqhXb6b8DCoo3wW34GdqR4Rvfdafl9
wCspG87FtizcyCTLS2kMNH3e/VTQhVDvrBPzQ9LBQMlk1HwhHXjFl84609YCSEpU
JQjvwCF7fRrRK2ETBQrjqlQak9+uqJi80P5WjXKNQylgs/L/YgV/3lwB2Yd1URzz
UtYOLxJ4Y69ao57BE00iUTQxAsoDx6ePliqPcKHjjfP800/V8UaYr85KKH+/c33Z
kQvxbu3kk5PGm84R7ReHC5h0WPs/rh01nZ1jRxKfKSQ3zN7dFTWD9WFeh8RrdFbC
p/LmI4SBTzAiikZWLbVFsGqPID4U2w+McWDxP7o4/ZFn5/vg68B0va9lVcVMW4I+
oNWZSYroNqfWUDviPYI6/faVOUXvP5eaHYuPurqYGdb6ovyYJhTg0eQwXFa0K4um
hlmXRFVOZe2PqKaoeHWvSjU5uEsp/P38rrIbMglQSmU0YmeQBQPTTQtUvbKkP1LC
dtEFclgUe/PclZnSpf+4poK8Z2hfUa6vD4rEPA1JB7smKyDl8mnlO+i9eJC4nLNP
QfoSfklvYzN+dDkQ4Rw/HrmfOR1K0CcEear6xRnn1VVjLdAL+/efIGd6mosxE30t
qXeYPRC5uwKMMdbihrinxgfskIbHunmPMD4TR7jxO1pIkuJrGE61Yqj8QA9c+1aV
5RZnmDGn3u66dx6O9t1wKXDf5vZ9TjiX/6qFdCS7UgYDn+RGGmRA2hp+K7o79KbO
tTk04c1N2j8tZ6Lmcp4FbtBTQf+LPe5MHojesvPs1eVUhkd2RIkJ8D32VxeY2DR8
M0gCsMGoYT0bU6lrLLT3fTr2UPydYaIstdmOtL3CbZMUkkoJcgRxjiN1KisMiFz9
gtEx4OxZJ4SQDfhVAcrVhNl4hHQLDeGEEnhKA1hVozWXkqFU5t5LVMgleLpwO40O
73QdPPY0kl5UqAukjMBoM+oRqVX/RehpoeSk/v7L1njuNX18/i3kep5hUIvzg5vY
kpIkKhDcYYWS7ohkxi7tN6BPWIsTZ1ZATCFmZkaBJpYhMjvJlMQOYNyOIiPbU2tu
RlrxBkNLAkiLn/pngsUMUmxthDBs8jIZTrc2b28WSTQwQRpYPHEabIeA4fd8nvRz
kDX88zT0GjZ0UDLpAnjn1QChVal7K7mvLNpSyn4L7l6daiMR7TdOOhLjpNWkcNYy
DpZ/ZrKMHCPSSA5qEo3VpOkaV0NOqpauqY3kptyNTuA4R/gs73XOiiL4q+Uz31OG
rcZXBmhAK22P8Oq9JYH5qt9gPu96j3qmVsSsrjcBEkpNXLYUXOOHGtJRSfturLyG
LslKBKjIiMKdOcDTtcNUKSuzIKT7tQdZAZYdXR+ddoz8sV4p2OkbI8U1J8XGPwSP
T82ZUlpUjbs7y91IQupk5Lny3LkfyemcMmeb9JcBP+f1ov0+mc0SnfimXdQhbnLm
PovNEaKhGB7HwFfizGA4MpcweEn3hawNQe0qvFFcFqHS5/gkgs7JU4nAkXUvM0HC
6tzieCGVFlXu4SYQYKuRfJI7CiveOYDibE5Ovj059jFPO9tW3jL/XtLRcxghZ6G6
vS1JQ6/13NpLZWqSx9Jd2TgS1aNp8Vf1MmyRbo0RGIYyKtEdKYBPSyjVnb/SvbYC
8nWEFGujngT9KRkgeORcWIqVzw4IFUqN97GYsgvWQzwJIpzOHxC4lF9BQdwZGrs1
pblLsMuUBXx39FV8MGxTpR0xofvMNKB9ZRkVJX4jNqzde2Pq1o4WRgrbdOvqHby1
YbvnbHhPxsWW2UMoqgAkn85FKHrOwTcUd9O61oyvGtFG+rECeeNdWiG5Hra3NGUd
G13KjbYzU9DBQbGdlYh3uym1FcAu7epLub/xhAJ/wsM6WoQEkpUhwB0bGs5HqJet
a4bAIS3pl9VA8TsUVHvvmmuFYKCeolOLNss2LBa5w1hGyN8vHvNFbZ09yeC+e/On
bg11W/y+OvjqUdt5bmPv9MooLrGIPbUL+OehdLlS8ZC2PPygMvtO0FYnnP/p+rk8
FU/ZiaggGOPheRzpncpH31ygpril93ow/TIoZSRug5ublUb5rEfDZ0t1PSHIBsoc
osfGhCG58CrSaI3p4Yn3nzRxbO6z5VUgv/Xmi4FwZW0rHnoOdbzIO0/3mkEKtj3E
+VzTS2T4HCmJMkWmIZhR64GU0RzKrS/b97kgDqm3Z6JtnNmkK4+BDa4o/xo7afQ5
b7BGMx80oP8eWRtkIiw2oVkLM44XHwBeqMqwIA++hY0J5y7EWEGNAPfBJYHx9XEJ
IQrs/ytO/LMzBmTZEOSDml55ci2Jigk4v9dlujY3wFxH/yNPgVkNZMOxl+CqWPQl
RnpXNYXBs+M9Lzy+gm4XvbAaFJIixf59OtcnSM4qNK7yU9vcBYArRoe3a8GEKPZf
5d1G9F1hdJ6MRONAHYatkEN2jHXZDMntKigLf8M1xaCvkdYPrPD5K/0F4WLknJ3i
qcvrHz7TqWdZj3Tpl1wCdVVT57WY98mqBY0gEQ85OgVzP7qNA81V1iuRaR7Q5p8C
AAyhx/zO1MjujlJvZ4TOeRD40no/20uqGx6h5JDPJov3makCTFFXlrJc8+6tQ7CM
v9OJ3UGMRUJo95VYOlbeUkCf5l2nJlR64shYvL0Ew9xppEomBHiMzUyMR0nPzHKI
xNRHjM6NmwnkH2Tw8zdZHtXTWtq4fkjX8R5fMTwwlg633r3aEAYXVCx/r0/XWAq7
WYPQwQ1TfZfP3RpN3EGjoK8UXVY8+cg3D6nA6OrAgwyc5/gVT829XFMDk8WdIRQt
fuNtYidNeCzTNh2QCjjgZqpRr454gs2at1DRWuwGi7Bb72/SH3PEp4E16ng/G/vL
ge03tztE2DoQfiisGt+KOwZzUzdcETPzE22TLq1o2Wy7VwcBls6p0NLQHQJCxnAy
2qgart0YuYbzxy70sgR9OzsRMJQauI939LT1bozMMIQi6RjjX+5CotqdGXJegaVD
bUvuryzFszDVTaEQqhJ97tLR8wUsWsxFjxE488XLl7Kxx8AysCosm7yXsvPx1QLD
XLUhJJmbm4poZbrRoUiMMfhL10ZlSz7wD8sLCuYLfrd2dnqiKoc0JctFrYPdkgow
sXKa1kPsXKjIxI7Sq1+9SAjDet9V+619wdboZ3Ac01QJN4lxWEKbBs50DtskWtNL
s8MpeXCvfmhKkKJMIXyBTAzW3oIdxzwOEGbieeGcLcb/Z6mStsx9nVgrb71UF+ik
8jLsYykNZfXeZmNhbDmwWtpwevOsyY6TqasaaEmfY5hY97K6YEg53kllJg9VbTY8
IZTS5zvv1wYlQfmaC6vJaf5gMHhurHOBEHSdcujA1KzAfg9rmH5Xi0vjIyo/qFQS
RX3GWeTzIVNPQGdVkXTIkqBnHk/rmresW+dLmqVd4dBEYVXy0K4QE6MrOSUyLEuq
e+IUXYrY4ejhSIfB48a9thBMNAkJHMxSuwRu+5Dzd5iE2hcWYhqI463LJytXinxE
Th8R88VDpQXtTd5ObQNcLi6JpgFMzbrpcgxOg3VUklHgtcYdNC8Sq9WDWemurzGp
fTJFPtUER+dLEAo+Bwmfc/x+GmcY3FuVZ6sO7Ve1ittSIhptN89a6yDMTYfuaWqI
l27NZ4z7qopcZE2wvGHJrzEGX20N/mq7MHy1yfQEIN3IkyE3ahF00BNVB7F1DhpZ
bYoKDJYcawwTA+XhWheZFWVNrdlUFvhijHNsJsFX5Ek3rRoVfCp83B7r3QkLKqcO
xTpGq1+WjbNzhDZYoPEI4U00J/lDvvHaTToRtZU9uoGsqEwVeMA2gUKabFSFuk9q
UwTQDjN2vUfnP55mUEXl7QYOHybhniLJq5zmy21/JE21sgIOuLzcXc9Z8vk4Z2/Y
V0Ekiwg3mtkMecuXFrfqixsXzMt+aviDRj4CuC+QKpI05XqJjiCnQc4G7IgBYXwM
oyis/mc9gJY7Xe/EIZnwB1gk2KjInS6Iu8asNFZ/FYEO8I9zA9ZjIbVOCVxnlyom
P77fii9vRNaT1UziZPpKsUdD8JwJn1A7qqb5pNo/tW22dPBrPrDKd3YgZCg4ojY9
A4GmVbzu8vhVO7Z599jH1OQYsAEMFN65B4R464ZUzkoY1bgsPW8+lZnuKpbKQGzh
ah6siPTYCMhutKD9rlBs4DbQ3KvOVfXMojWulMPda572sT74NNcYSANJx/YjALQf
tVXJkmO/zSDz3GiNQ/yVPcXSi4vIJhD7A8oj4mCMXgE9CG1M1FqQoq3su5I345zu
iYmV1/XPI4OvJZ+j9Hj4+e7l1m/JY5suY4ntv0FMM5p2+f3etd42uQxsYn+yhcv7
OCZ57bjBjkhCzPGWN5v6Da8lio43eHOE5DN8iLr37nxGr+7axs2YuFY3souAtmOg
4DPzSH+MknQjNoi67629UPOm6wFY4OMJxUkJMmBEmthcIpr/WCalB8F+amvBSqs4
`protect end_protected
