-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
9EVjwMOgRc/9jfeH/eFDt3Zre8tBBs/3/G7EgKWQ0EkQHZ93Kz4tyLNURcdDOPfa
xmcCmViYlDRvTzoIYBTHgmo3Rb4cljIK3tqWxduYFp47tUzQQN9ZB5rK6gkgEm2B
UhUb6PyuG4d3V7BB0cYzFnXgef3TkuIK9Msp+v6rjWVxu/GRlLOu5w==
--pragma protect end_key_block
--pragma protect digest_block
jDBMr33YafvaLRry86u4twj2sTU=
--pragma protect end_digest_block
--pragma protect data_block
NMeFZyCBRl0otHlwAFGuvh5bJkTjm3ESrIf3OHgTWBm5YzskNE9xad97qZZnexfe
b44dVkiSQoHf4p4jZ4LT7jmnQOL/1isV/usa29EKshGiJPNpKhz5hFnW0HdpTijO
kk5miM97Q9OIzaTpVzoFg4FeBdFY9Xw5ujjfbgiqvmHOrTrwEHTdzf3k6qyeSCm8
Xd9T1Eq/TWNw9YgaqutE4rXkNPpzxNh3yw6y9jqj9WJ+SwHiFe2455xyOS9g+fdf
Gd/FTye/I8/tu9igYgudee5pe+lKXfHygQKr4v671lA5D43i7XWBnEsrbJ/CSEHA
JhROXGHJYl/TY9R6mOjOso9w5RCzebYZbnxwizur9mtR7hp5/jB77g7gEaqiCzJZ
PMTw4SG7DJ5I3kJjljmf4H8s9eZO1MMlQ6KU8rAqaljLRZqhzt7aO5z9ObVSTgSe
2vJz62Dhu2468ylZMpvHP6mDwCV40tt9SPMn2pIyuFBFPM0eh6xUehzupMEngpiq
76Q/tjG7OsJS1WiAoJgI1rhMRIrY8h8KljEhFciiym8QJCEw6LO+eOTkz6asrpf7
sDEyvCNC6JETInDWJQvOf539YJVZiNgXwhZYXyb0kl6IsR+4rTNX0yd4gBTPI4h5
0cbZCSXcVyTljm9+jfHZ7h0bf+1zO9lOWnnTDis8UwsV42MuVj9dRSF3wzitgoUl
scT0pXkRWcJ1o8AZNfvytXxlcD/YTHw+Twdj1I//2GgmR1Ber+3x3qdF5a0BJAX4
hlm9zzQTAPcNShxBSfQTkNqZmizlm7iZqE4gFnaaMZNQ2SWS+rzbXVRI1UUlt5jg
lBGQ63CX7Pu84M5K7ZXxeDDlRZWsfpKT2SHSW89g7mEYJ+mXsz1yQZZ1+WdMulc3
QPwzqfYYSUD6qiNQHRMxErqi7LsEQ433NTSiIZy4xGNjlwbvrSC6EWT0Kr0mhz/s
XvdoVic7EzI+IuqBurIOB0/90vpDwVlNyvDo2xgJ8Nx4Ar9DsFaGP/AwWPJztWCd
ju+vZfm456G+8aZPVBLMi7wIGS8t4U9Tm7OSAjdphklqNONGTwyMF7R30Gx83Lhr
qu2fOJ7Ri1gF+NGARBPXelysnzO+Tdh1sCLqBHfidN+ElkoJl9LA7mBjji7XMISx
220DVjhRW88Syq7AZMgvGls/hLym07MvUV8pUniP0JRZTifKPwpIktHJkyWfFWs7
tJRdYxETZy2oykH51L39Wc0iCGBZ3gG1FRanSJr5gvqhZMUVos1PGyOEHS9U86DB
ZMYKr1/j0E+p7ea/zY1GjAR7OKJBZILznmkMrDjUYDIR9QI7GgTvMprH7Cf6RIIk
fsFMNZeGiUcVls802AT+kJ5aN3slvWEo3+SyvaOQ4/W7155XYq0aoaaTRIc5KAUd
HYOPXwY94a6hkPBgUaCZj4ut2vika6fM0VHR8hV3u++nUjCc4ADCHm/EHJ94JgUh
gJgbpQALvyHApNDiKZuiuMyZMQae57286Ai0hodFpK7l5zbTKEubh47vZICV0DtY
DB88icX+na55XcdjkaFOLNUXyUsvmu/OEQEmPpR/+0FlYufeheKn88jWesmCTqut
Z9rOAVzyzgjFdSC9Md4bWL+O23q92xLpa1WkkgLSLNEUq3FjBg+Liq/SH1zsUrn0
nO3D9InhVmSPQSXRkOEUoVJ+BsuC/SANl00zcYOspzNYz4CEof4mrp53fCP+v9a+
nPSNVbO7fHTJxqhlybiwIYd9tIeoD43TYJG1mWkEXylZdB9aNpo0RNHp0eSUczAJ
ZXoS8ChO5OK5/mx/nmthxpFF9/3SLzMP1x5WR/degbQDktbiVffYekUzvSi3n4gh
pjSicZPqYDLG0iOuA/s29pdt3dxtMG7vL/gKVlrPGWkD8IUlAnuWiOybX5eyig7l
iTxXkzy/YRc7id7ihI2/TCJK7OUK6HIWPeHLEmQVLK3rpgEOOFqFWdHX3js49eXD
LcQ2ctsiNL1uqy4dzlI+v8QE7I6+61hz6e4IS725eJj65TEt4OuuY3mD4jB03EIM
1QJ+x432tZGa2bvYpqZtTD2X/BrUcnac3WuLi/OHN0FeFNIvBe0lWBFdoCEhITPj
bUDmO00a2fQ8mEw7t44wgg4c7CTMol35G9+B8F4wpdbwAKbGFdPmNmM/lbq/lGZM
KITRNAjFurKagrHtXCk/v+5H4FdCEvW++5ijNa6KMrlfteYfgp5jxMnv6Fao036O
sZ4EMxhvasm/4z06NnvIBlHENTTqwvCUlaPZYoskBaq5gNgEbQpU7817RCuSSjH5
iC4+eoBV+d5oBIg2gtYQ56ha9kdnj7a+MxSxxzk9/vj0sm8K08NcfC10mZQCSvGC
xU6jrsqxtIKyZ90ZvA8Q7D4omSuEIKCazrmvi9GxN6DtolubSPGja3KTahFPvq2h
XSCxKSZwYB5fXGCMaszgMlgv7ZHXsx1iF1FscagIcsytDNA5qE5RoRkCY49HOOi0
krvO06rVCNBuDvvWj6eXGBxB+E7bBrNTfc2EkJjtnJo656En1/q9td3UY27vJCkL
IKxscIMj5WmygrOA8SqP1xktfCKPBgFMF/F7Wo3G76z/LLqjmcHVlQSoO1ucCp7h
q9SuonryP7nOIsz2cBtEa8XxV7vBwD0M1qP95bFyc2yxv07yu1uc4Ef4Dt1uWtw9
J9na3znMKveKpq8RAFIVqHUN91XhIwaLG074z21l9UxB5zBwUoy98JjmXnEP1J1j
5TB4rtH63Y5+eleyvLRe2uBdL601Fxfi6Mnhea63UTzYrwAJWjWoCwv9ar/1feBf
paiQS8zXzKJ/ogNYcl4jCyY9GkIaaUTmSbmCsPyEihmLZvLJoIQ9JxHVfzfI4WFC
CNjRhmKEVXPlI86o/afcQOBEJCcrB+ewWG/B9sURQC+pQPiO+Cay1Vsx5OE01Uvh
y2rf0jR4ZAclvZeBU2f8ORka1GK1gLbyaiUeNDL6IqM/U0m4rjESl+tPFtYDjJae
cFv6qx4CIbqhyMHpsL4i3CLWjc9VLtSc+xeqkpYvIXmX0UryxTXOGCeBY56eIWbp
0lfpdmsclCRdBNaVsqaU2iZQ9GiocmeHudQKicLO60nTACd9XHUZ9ZjCJuSd0fBR
Zk2PrHP0qcHgHIqFpco+0mYEsEr+4lvwKIB8LeTyvL75APAOqmliAFtYkIUHCp4c
Nn3Fsh5/WHLQdlXKh80SjSiNVY7G16lvjfi9c3Y32le5v6lFPAIaC+lVL7koNRBi
mJNWYj0JQlLg0axnWTprmZcNEjkHeKHPjeqqVP3VMR4QjT5sA+E75pKvgzEzAbRN
qK1Q2Grj9wmohe9C/CFE7VxRFQ0U1i1NFsw3PJD+wDWvqemxmEVxyS2OLW0Uy32b
gf31roKMs66pVOSM9HAubGbseORM2sPL4EWlZsldLZCq3jQnndbQOADbaS53JvKn
1VKuY0ZUJNIREdQITJX3mSIzInkNtPTSP7ngD3JnkE/XZjUnkrQpj42YwyNSIwLn
fyYZXUX31cuYJ4pXzHLxFeYZQgHXbZA6DKTuj8FIOMP2Eb+2M04dL4PSxLjzI0o9
ELmerGgpQpTpxU7iyMHLrw69hDnroAb/0wo9FPCwSfVMUmwefEn1moGH7LpHV4Zv
ZnHAq0rIgifHTG4hlp/CKElms3bIND6saS4srOFpsy+eys6dfK2g1e0y/+7/RQlD
v6nfvUjGkIdgjki8xm6v0XHqLM2BGjmYCGi9JAfVJdzevIk7voPBKF/ZIyBfq0kt
8JENLNCJS/gHJjG92wizpN2D3kAAi94GciKQGMp+okw6UtxirW9fXqR1bfIG/LWf
QbWhu3G+f1B/1ww+Z0pUyCcEHcBTIVIW7x9gWswSlBywaQC+9CjusJ1NcGD8YbeE
cUO22+jAu2664bzTgdb7LciBTE892cliwpKsX2RzhVA6ePKVxDyXI82NUuV/KmpK
mfdJGLjS8J9AGyijBU/DlG45b7F9eZbNI3nSSrNTUDaEbLqAD58CXqBEfwtxIU4s
OIka1vLpps6uY+IG1a7dRl7cE9TTqsNm/lt432ju5AynRdFehRrIU4bKcnp2zdj6
tgKXdqEE75t9m4MrVTcEgPM7Mi1WxXZB7BRgxRV+yBeX/CsUKiWB13ugBdb+IKMJ
5B2//tTqgNbk9Fdo7Vj7vsUIWEJwllSS57NHfLMOi7P643/+SrhoplkEJcj0dWjg
fzQB3tuIADT3gmLItY4qVxkHhtgXQt0nIjXgJBx4KRvgDCq5vI8E4InoDEZ0yfRQ
YweOH8K0bByMSyEB1SmwPxUNSPcSmjaoFIQhiWzRdAez6N7J+beVFSE/V3RMZa1h
z1U62OkytlgvjBB3V/Oasj5f4X8qz6pGPU63FvPATi+2TKJv40bxxzojw32BJCVt
3aV0Ra9AE05/keGPu76RhEhCMqkOUyPE4hkaXjDey06zIrgJFLCwgAmIhPVy1Jgp
iQ3K29m3iievxrHKe+bwGhOpCO5Br/3H2jFGfCVwGwTST22quQ8+vRB3BbGQEohR
4CetJmeL4KEhmqjI+wi1HivyGwWPAL0fs9YeVUi//5/w0f0WZDEDwbQwDpUE0Dza
UUJ5v4kngIQMScccvFo+aZIC83Avi5V8aMoiV2Hm/RXXUFyFVDtREWnueG5iADr0
emqkxSKRsrFvmZNlF2icDT0neYfAvZN2MVaFvkR+ihOJZkjiUEyxWDyM1EeJAJqu
R1iVJKJ2kvt+ER+EFX3B3QdHo742OaQYJ4rnIIYIgsWo70a5yi/21G4yuGpZCB/x
5O5w32rP4s4VPLcahHZ/oGYC682W9K6ZbuH5tDoXwJ2LkTFbl06mIbe6+BVWU1+p
rx+C8IsUgdHfwk5hQGDoEp+EzYy0UKi/h5u5vvejiaQKjRVj5kNVzA/wuSYzGfJx
YmqCCKpbFpoRXFv55Fv1vjRsNAY+9MYpJZaTsUEXlBG46q8bbUQNYsPC+b/kon7G
VcoxDow7ZJAkK+o9okfI96dTe5wb+uEDNvOfvvkVRAsta7ZLpl2Iptc94cXg0YMr
SAnK7gdjDLZTFw/dRdNM6R/rKazK2Pegfss+VWXjQYK8TNNq1FVNGArE4bfEgmd5
2YfsDOiOiB0y0i93a+9VpD2QyYyTVBDZT+OCqlVn6Oe2bK1bzfjmyCm12kSP9sIa
GgEL1KQuYdKz6MbdgxrWzhC9buI4OkHHajbQe9hwDFxAhI0mLAgnSofmwP2F4yA9
rszpUD2SIDjiHnwndvKQLOTiSXhRtb2TnXCF+02KclWXsL8SZsq3GwxQJXAnwECG
STi4aYhoHthUPT5xQ+Ww523E0NKOYzIq5cfQ4gWojEAvn90/vE8dRx1mzKullmAI
eyOFB8HrAs3YdnV25eQZn8Vqy627wJSBkpkS1UrWKIcImPWRCt6+KI4dX7iSxPiP
WAnCKb4Q3coaXGizIoQ6+c85R4YUh/aD4Q9a628qHRlUxLOKcouNNhsvotH2zBwQ
b7RJfU81UTZ2S7S/uunDxm4caqev4S2CS7FGRLMjWVKzebVstVWHc/yrf5WkIapq
XKlbOjqBug2rbzTwMnMU6F/PdO/FOF1hjb9HR5C5C5FRfNmvNU4sl3KtrQlkSgPz
nzSBh6AbsQYM2APDnILl69PSjG8QrTbvRZjZpDXRih4JTq/oM1cxpJb8xFIDmdc9
aGUbtSdM5p8h2BQ1FbJAgvot2jLGbr89C9lDtiqSCZG7QkjXqGf52ceW9GMaF7pH
O0RDXx5x4Iv9U6vyvlyBgCZWWTJyj0KotRqtaZawTOTCdq4M6kUqHmQh06UwPR/G
oR5mS9KkW/qTn6WEN90iBN8Jx8pLBjIHg+VddFQNlOlKdmCzcqYQOxYEiJWS6Yek
SC5ToPQfW7VX73GHIEy6rf2M+LkE009kdc3+D7fE35powjAKwnY0UOk+j1TK/3lQ
TaTsGiGbcZPU2/pq2Z0mwvWlGcUE8Vdc9Qcut6C1jEj+6xqPIOrTjPsmkMLweRT9
UD2DZe+70EJ8rZN7bj4tzbjFn6CkjZcP4CFSYFWvg7E1IjOBHbv/aG1GfKV+NOnV
Hg7wICxpZFbEQoVU9CRLfMYLoa4WNdlOAR4Tp0GVjYlw9+rMHMP52DJ2a12p1QcU
4kngW5iQoHjPrRHcgUw2CGJ/X6gJPD86xE3eGKmBi5xymlRJpvPHEOO3xm6xJ7DK
JLrpqWLiV95WBwsvyYu3AbWeuTNwGy8TxPYQVWQHxYOHkbmeY/DZd7MsUXHgk0jR
xjzRvoVVKVr5roHr/fsyQnYJOS17tWwwKMerutsVQ/tNkL7hwHyunH/Z+uVXIWlX
721ABKbDzGSTwXJfMluh7TH6pJluFBdDE+exRkYi4TNB/LeRGYsnk4/3QVgdx8NC
AtqCYmlV7M0fm6D8OVbuNQ7m27jn+0W8/hhVW4HhzKNu221QkYl/f4pWbwJiuBmd
NtaVEzLVROTSVpxHt+GxZZTqV86Si08Nnlq59hiMcuhnu8rzKp170o6cMSHZu6f2
e0XX8F2+ABmJfbGj7nCZTpB4H2qjroPeAeOmY41N5h3MAxMkwIazc31ynYA1++HZ
WS3xifBi47qR1i9rN3SCzG4PcDLelIC94XgtPqJKXl/+EjewO4RVxBujDi5VSWPE
kzU33wrnCWztfRzRmHp51Nqlvi9Ne13g0t+n37PWnc3JwbwdoVjJccgwP1XKkMOg
SmI5C2+mlFkGiMHTKBiR5WMqQQmI/W97jMiPrk7hxPx+IjDExL294aQ2KuKfi+Ef
HpPPtmk8jH9LAwevN9yecYOdzvCd0O2PlhoWVDJqwSXKeDwcenKKUQRiPyV/noCO
fONi5piPbhkFVVzKls8qK2sQVYEYBkhoVsiw76LnKiM3YpTcngF/oiN7COCNBkNg
U28XpY8A07TIOeAwfinfxZnIFganHCC+jgsKMUec9GiOC+tKj7Yifc6NrOCsGHSk
D69uojjuaXPM5GpAEmp/mnFTMiKXl5Kl2od4LatTE0YaWiNW6qLMXQmnnoihntWQ
6Lb1a8To3SLf96eccUayPf6BPJZLpRUJAEUnjssZz7OJmxD/TsEXz/QyhX/oiJ7q
Iqlj/F+KjuN4DiPvS8lGlPfTq5aM06Q/Cwbicj6BpQRxyIWvuYd7C8qCOwD9saXX
77qvynnYmAHIkkzhmDJFQJq2BPzIaLufK4/iC6iReZ+mAISnMyY3Jq++DobPoyav
x3QmuQYPim1Q8m0G0sv+xSVzrePKydqjYMuAb6LmyyWkvHoaNP7SA8bkDGFwlJU2
tY8IXG1hUo1VLaO2/mMIyU36nWsofocuQ+F1KEAypHz5Z7/R6/AVi4LAs6cGYe+D
KNVecW7cUiOH+eUwf7BXRjr7yxrXJCo+JpzwadT5nFlor6v6leMLjNLJXZxNCLkg
M80oscuAjswkCCbzw30ZeDrOs4m6vYrl+H498gHQuqlp1W2XJWUagrw/SCkFawrX
7qXV8MS2EYhEvcZXMn36opFVbShQIK7ChKhXigFLcvG5STGy+6L66X6jbNnCOLsU
uGMPNOEgkk+7xaHFHm1p+OqJnZMpsyhPO0iAqDIu7nVoLYnYEM8XozYQLZeGrTy6
JPleNuP989yX7o5YW1+2zNpy5hxkP1REAIJ2Fh5CNI71JW5yqUg2w5+zYXT2Oaop
4yOKr1EzON2AztnYou2CyavrUlhovsLbYXZ2TncMMYvXvjWNR5DXMozOM3JwgLCF
00iSdV39ZUP56dKaB8VV5Cdr41aiSTyOoa9Kyf0Zednlb8J84PzL0b2q+fGR5QMK
Tn/KFUIZYcoPZZ7Ofedhl9FStBIsJRYieG7MGkVS2PWMFl2glZLjMADTWUomfIBS
JvznZWhPYHDJfIDvEi9uH5bWamSgOtTDkeNQkjbC3vRW1AZgTF2s6aGKfmUOO8c6
12DBDrVYyNECkzT2JfBY0a/osMJ6WUoccCMSf507W0o2T4CK/r9LA/ZfUeVSCJb2
gDLfetw+oLuLarZs3eraWVYvC5DHjr5+sM0Iqqpal3jOFTtJUVeB/2a2B8L+Xp6p
WaDSMwhAQdi75W6ROd5kSmMiYHoA8jlco05+LHozg/3JecsQsfvo7DA7+mZbqYWr
/di1amzBozD1lA29S5IdmYG4psXrl+fWm3UpSuedZrlNuAFpWMH4VyqYT5bMQy0L
fRucBhaV81df0tjwP8b4sAqmSgPMVxr8cvLYaV8mTQTeqABsfL/OepOQj0vH/41z
qfWr/8DVL9n1DAnS65zOZC2Xoo0NJnGIhJGkoPp0PZpke3uEPt4zlpbjLAVI1w6J
sjY8vrxN0cuvJAN4uEj0v8n+KZ79JY5VD8/02RQtL104n17/cp1ChW2//guBi/1D
h3CVTQFCoVNynGTW16Ub4lRWrkLc0ZD81E9yC9ZRUwhO6qyvC2nZng58QRR1S8B9
T/7EUjqicrmvVaFnzTOwTE3yRs/B/L8UNiV8B3PuHD7Bn3W/dxcvyRGOzpUYoQ9v
ihd5jiA7fvcHUFX6ShdORXleyQttojpfTGBKGlQ/pFZ14coCpl0F6FfUkY/3TW7l
mW+1bOHx5tlrJTR41P4j6A9SZYA32GaBmJ6EKCjr+ozbP9w7Wn9dsqkDqjCJLs/A
SBNoHOW4/2Q6chcoNh2+28QwO4tB6z8vAWXzA6HCON3yu1kax7f3fy9Ph64qR2hy
8mkw7d2VezzJRMzhBKvTtlyVpWKuxJ8saMqMPq10+JxXJWwRqCY/hgt2EtEKX/CU
xwOsb9MVT0FtsAV6HQKEBYKvkY1XxQyWkIUKsaqxgZ8DpZrI+0XJ4N0gauTuNHJz
XTkhN/S50YifLqg5vryOqQtI+Y2uJ9XnmE+6x02qHzUAKrFXoZa5tWTlPA/pLeiH
xvZWg9QJitKmVA0xdHKAd9J/L4eR18jOiTahs+4WAuwVsldLkKpSmgwmAa/nGsj6
qWCKJ2J3+79uzvJ3b+95o2NjZGywI3pCPUQdiUA0yGrU9cNWsjtKqq7w6mZ9v+Q7
aZKtTHraBrJiTwIQ20d+BDFGzTXDzL8qHfsxIaUPossx1s8LfTfpXNRm2JVmCbeQ
jkrVi4kPmSV6cURAidKSg/A6ue/3qxSZCF5ecQqWVol1AoRzG0KYcIeOS373QwFw
KuXcfTytZDKAzqH6W9AqGXQ5hh4yvBDmKb0yVi+wIvkY/BrCtPXNkWOYEJe8AkiD
8D06b30iqoXiPq+zRUzB+otwgN22HRG3DiZkU4bqQ48n4nAywvZxjb15Q+owppAw
734XWU4J8dzmeRwj9aSEwFsoztqyFu6Sy0bMNzhBpJ8UDzDGELwx9JM+GUfspaLI
9jq0lRFm+669DG+rZQzo2pZuUb/GkXUOOeIP+kFeLafVsBG6HAGUj1ZWuH+qjhZ4
AG6QS5/xyOACzdoN0Q54oIeXQwCIUKiUUO+oKO8yoIbW1VfIHFpJi1pnbQYPtCeb
rmcS1TPS8cw7T33DPov1Z+V6pqaLT/VjqYtiyBPt2/E8Umb8f96XVxrk6aGfdhNi
xSVkL77+Q4qg1YcbCOKF9xyAefZDDNcPnTwNWFwjYx46oxmza1y9oJuDiPKP76Kq
UuwiYehjIBjEU73hRETfm3haEL/YzFaWGSLYzJFLymKFgN4GVprH7raTNBijpeVA
xuQ9AcOJYLknFt3nfHPFxRiQiOxGfa2U6q/LYIyFKmeKXDufw9V93p3PNe7unpcx
comQZMJBcVHne+lGGbYg+2wyKaV7gSPpWI7RfMLS+9QPrfWyWPBkZHTH0kfTX7zk
atYwCSF9I0TJtfmxJp8zmZIyprCfWZ8Md7JbeSr6QRPAUkcOSO52UDZnvKmAAJHP
MVO4QX/H/S97nsfM/tzeAuMTk1CzBxF4j6AD6/bmNGtFg5lQH8F5cui6E/CNLuZy
Cx4mvN7PlJfU7feKU5po5QrFRLrCOqCbfIskPEab9DhWqtNEY6oJUuYLiGO6cZIq
OxEg+4Y3q9HSbsuIFUlYjsvfVghJcZYbbAy7DKZbdXDUbANsHNzYzE/eyxsvjKUd
R8L/6v2JElKy//FzTxK/yHSnErhrRf1jhIVv4+n5PR7YuNaA2iNlDtGNy15jAuY2
Py7YCGu0b7h1l+hPwvvHI7ErUmAR+zymgnGNnoybJvWvMouETHM0Kkf9WtBSa7ct
BTIqBBgbSfsYO5wcnRqVLUjfE44AFfyoNXevfY2c1jO1/DIJ3IZbItNxqSfylQ9V
OGN9sjI0bDzHy4stJs8cJVv0IZ5a0mCwtq28jaafNDVMt1DPCEtZ1b8q8lSKsun5
0UQSTx6GbHSNZzMRUv5JbSM3cjiBXlQWL+f0MfdJ6uDiq+PgCgMStLrelrtJBt8K
mK2zEnImyHYdz2QdRhN79QaEWYgwP1nvpSyoXw8/KKR2BD+2Z7KIqfF4Uos3lrlx
PJx1vH8BV6tTFqeYjpTMh0ku2VIz9ozYD7ML7kAxerVrNsEAnFOBVYLSlunh2wbM
/KyY74Ydwr47tUOXzdGx5gNJaxvKimjK/xhZvBC6U7mGvMpUceC/rjNc0+4XrZ1H
vMx5GXk+5TLpOhwwWhmB+iCQdk6AnPcx7LKMxPCM0Nhvr2IHaGz/KeeK8PvAVnn9
UF6vp6tasQJZMXNq5u5qY06TVrJmPB4Ako0bTgRQcq913aZpyKnXdhZlH8fq3bVF
kKZJYARQtny8r/F+/sVWUcFYhzA4PYi+w5JV3+9+Hg0Fkd+nPfQWwOwazoch0eSd
LhHTm0DwoTWvfzjYEwu8a7lcrXIVxcpE12734toSdj3WMn3XflyTkLOjcxpAevNG
doqYQaujqGxr8T24ds7KWfXXJnDL8Jy1Yhai6y0OlcbKAytqvB7aSykjLKjTN+Mw
1sfG3/kC4Na+Ii3o31TmRQIUs33BTjDCqoz0ohBzPxosL5hDO3+wbfvzE6v3xWku
cEy6X29Ep7HypDLiwYAtt281SqH/y53DyixRW7vi+1uUu1QYnNaizQnvNYMqJBrS
5IR5ohFcNXUopck4MCtGnh3RYYc8HUGxnqRfMUnGi7zcf12TwZHCo1xOgJw5Ry0k
flUAADo1Yjtz0rMlfXYwYb0KT3mrb8BvmHZuukzDKVxSZqulH4ViSVrFuHTaM6ds
kFU9eYVtToKKZuOm8zNbh7A9mwpLtCP9TL9WcJ9ICK2NlsxgHn1uOMk23EbIhWqW
KxpLC8EQknfNzkzGWmGY+tdw7x4llrFgT6rWvD4SPJQe5augwUgycs45LKXujrrH
dCSJuBn5SGPoUfWYuDzyUvA9bgs7Tc6VqAorHE7y/LKHcvvfpozmsdrWiBmI97gi
IfaijF7/aQ7J02ssuXSBs8CmbyQpIjZXm19iDh4Ey4kN/zhIzSTGan7xwqDRsMz/
pcewxQE9u7W72kmJu2USBrOUjSeHUH+CXV4k7eUvAwzScQnakYwss5VAjpuyM0v9
Uxw0HqhfbbpCQfeIU9klO/w3gHe0QlYm3ecJkeyQQP3KiI6fHlCdUES76UbjbqaZ
oyC5iLaGi+Uc1AY+iqGNOEECmQD/aITorsOplXHP6EUszR14GrPqSlsYPXMNMusL
qcoqWHPCg/3hnVTpwfhPNw34xm4C2ODb6uEgDNcuvMOpFM0s1gYIJxxjEKy70JGd
cTQ2Jg2xanBsdHmOS9jlWnqv2Qnn75ITReS8QMtQ3Uk3qybb1dKq8xTQbJysSgCc
XyDlV+0uD/RrxNoCQAmHMfJEk4pS+NW6NwaZxSszPQsvtnpAR9gzWQx9Rzme9A8v
vjnAwBi0w8Jhp+MjRfuibo3+3QoARASMst83t0JmocfBJevegcuKo7DzteE+Luea
sX40/tVzjBAhlX90FrlINra6uBdk8ZCjRa0THV2JIpBGRr6M87UTH8izw+rxQNxh
u1hxMCX3knpxtq4AW1fUKhYzwM4VR/sAfTizoWXz1DWImhxlZLBKr2kKYCTdG4a7
lKpjrxGuUpZrvbq9jYXE4UL07esO6L3fJ4Q3+AJhTEFFSaDOgXHCuuKMF7PJdtFr
4LHGivt7wtjz+IXUtcGqAYEKw7KZjkncANZiaKCxdFIoZbrZiQ9aL518AI6D4QTW
f1FwUGTnhA/FcDtQ3u91Mpeq8ydCU6G/Q5BZAfGI73sDCRQHAedQQ8fWdxtqNm3G
IbLGZuhPXB5DkKxg0FSXsuCw4gItTfkoQJTIEIMp63YmTDLYkjWChzsSRMWl57E2
DG1YzJX7cRLcTVJ7kNNH/XotZ55oQEWR3XtcQV0BkmHP5xOjQE0iXAhTLkd1tVwq
pkCuB8a7KWFx1Z2r4ZqIKhF1Dt6RMi8zA5Nn8V13ByHcREGIDCHW3kmeZrcuuwgx
Z8Cql4VuI2Fi9nJt5bFraWZRahqGUU8LU8v8fyEjBjqWFCScFzHp/pTzmRCxV5lF
XYSF9vdCbNmDDJQA7o1uyXZS6us04t6vPRWHWUYT22+GnCXRwFybVUa8EiHyHkOC
iDsnJEvLITk9GtprEKSEptdap5+TCxOzWbIZ0eA+0eZ1EzZuvKsL+X0tgdfAvPkJ
X42MEg7vigspcNzqQFo+KGsDkZLBUsq8+YDV9gHK8oKHp2fLNa9iCYJVy2GhPOQI
SVVqVhLM3BT0NX5MnhD57fV3KfVURMlk5GfV/D7HpynPWhrWjDaixvB+0gMCJ20Y
UzU7LBygFemPkUKs67TdW7/ega7v3bXpyWvabuCLYJBN4v+rJj3KswLKYut2xAzg
m4I7P3XyYdaVaRl768TjVFz1hQ59vE97i3VEPgKUBHVpItoP75lANfz9IPYdRAhe
HkZID/w68pOoH89PXKad4PhS6ALEpRzJnJcTwJCjXu9Mo0Xcon7d95TzktxioX65
83URUhoIwu53n3sXten/by0WSjFtAr8qFEWF79nNOEUHHJuVcaaNyhr0xjWdGp+f
qaD3jQc5oJ49dEKqacgPZOQPa8nJGLCh2oJSep3HnBOOHh7n32Y2rTUeL1hw7p0q
L1FODQ9YRzrjsDzZHcevAi3Sal0bxIEZKv4WI61fLhqA6W9qUHoBWGG/OpgoaByJ
3tr5SmHHJbLKJf8LpPqAZR/7ZpXzE/gX1tLraiV9HTLYYHPhgc/kjFkggtK1I8vA
76/dP4PZDqZTU57hbohbAF0IFtEjIQpypEe9HP/aReQUP2M481A4CvV6ZvouYDpU
FnPz4tdnogGgtwyvcBm0w0QGB5mjDyaBEpCMoOIj/f+3M4//q7q+wEhEzabO93qF
xaaMf7yZZ8M9wSs5RE8Kq2624GGOPY9iqu6z5EaKJpw3NhPK6rGXG/IiGxlA+JpM
IWCiVTrVBMGDUd4tosqpCNMz5YjOjs1LtdiUvyOMW6EaqgQn4j0ApEPzS/a9B0S/
TFbZiHlIuLSp39J90ITDqtbfgzStBmjnIOjIipD7XeTgCE4fTY7Xikgop4D8fx6c
x8XRbHrgiI0mWq8cbvJopSOtNJzFwDQ/fgsk1s1RcbF5nVkanUKMDq5NBsmYNMsW
wkL7ejv+oF9+aAzKu5YfTM1avBHTxOs28JO2UlA2veqqnZbv5nluylNTnjmpLMdF
Gcwsd5OEjFkSCs4mEn3evj5ZszqJHuK/KW8tAys8jlnVO3YGSeHapQJitahsSnNm
zB5+PeYzsnR8c6vGzDkWWPBj2FppsH6bvla9JfiQQaMyXQ/jQcz0CX4okDJGLQmT
kzEqzd+0jUdWwwhmRiPBT4uXW4JN3alXivZAn+m5AyWRHzJ15Imp55DNrUTHbJgw
TaCEwIXw5+dSrGY3ZZgf4QWweADmWLTH4ft/xDDRHqrf/2cSexQyVrIpBr3hR/+A
qyBUdj6RWNwWA0DVJKPMdxz4Uq36Be6n4OpdQk4+iWrOLpWC3+FXWoBWPsoUvAtH
KPOP1XlzqLHae5GFbiXLnqrqrCNikDc/NWIXiEcmJVTr80uiXq9kgE9jo6uYuBjx
QyOwvMkS01OeQTjnxqE7BLivL/+AX1AgXsQbPoLKNNNQeqIw90JgnOIfb57NlR5U
LhQIoKtd56mUZfN7r5nc1NLUrorXs1dCQc0wQWIznEhDC7zVqJ1aJilhMUD6XN+P
Axb1wFlt4vGjV+G7zTRo/vyBfdgCGLWc6TgxU7RqNx5yFBRIqQMSZiMtWG1+dtx5
DEPV6QnmoInGq6wXJQ8ALP59tssk+u+S3wWUsl9RRJIjs/SLYy3tvalOyoCuZzmO
YF7WixRKwPh0o9PN+XAaa1HfLSFCra3ZTgzl8zTJ8y53rWGvl3JpWJbIE9Wm5jRu
bcNiXjIOvHwqYWE5VSsDIR6S49cM1Q+1/Ylds5hPXiXA1cLLdvjR5zxNv2bevM/a
drFRi+F+X+ByK3AjQrfvFBwHfum0nSWXoH66w7veKqsnxgZU7BHq4qr0oXZ6fRcx
adZxAaFexeROWamQiwOM7XDO/N8ACpfKQsIaME6tkLvWcVOgDwkKuiqWAIUgX1G+
uZXHsFwT2My1ofkb3SkxeQUAXyaItXs2SNH5RmqQZXGdm1DFsDa9tJJ4SLO+oC8z
hYz4j0EC1n6vjlVROidof2YHZTdQjrmvIEKThbEXtN/Rjkt1pJjwa8LEAPkTTxwg
oAqmQ9PWuqa5lFn/n9KAMz+HLLrXW+TmGDElwNFVU2Cq13AnCFOXdaScnQL1f0+a
QByvS+43ie//I1eonylezKuXh09o7xIvpEyCb7t+ShkmcQ5Ei0GGl970IVPTPIPM
bMTYl6Ia5IplmWuIBMqPZb7DqutCSOTcKXhvyXDfelf6WjWKpJvlCF/dER+g4As0
6jZBTckvNpBfsG8MaaN+VwC/yjrJgbxsI4BGdZbXZe7sg+Um4yos+2MzNe+VbeS1
pPDcu6V/Apff8tVBR+ZPizgzrVqgJxPodyfFIYra4eMxj3oI+HBdxZFs39I9Q1Y2
V24b/cn/pyZEjhqhPZWdPA1SKrx4+VxGWeFw+6uoe8jmG1qiQlpEjPLtKt/05BMi
h4fB0ha72r+kgU6uiHc770o21Iwkt3GJLAImB1GFGIeq9CTosugG+l2r+9SFyU/P
yB2urpqg1dHb3iifho/cUAPn2IHe62x5QOUO4X1ta9V48XIy47us8IvkmZlZuPqv
CpDvSZIaJGx0QpxHYT/JSy9QNOfSdlmoweid04pFx2VcsKg4OgYpYxXGhMOM0vhj
P2mgeITohTaUjNyurlbRmlzLqZIJn+hH2PyXp1RhkdrlidHIuRU80OvvX6Af7Nii
BtPtPk1/SoGTSqzEQz8ZEM/pm0hRPyNbWgi44AY7Nfn1xtwjLnfN3gA8xyXP7t1J
u+yKtpPPHtDMREY2v/XH2+m2s3tFYEwvIxHb9gDNl+u88mT+4boKzgYemY2F40Yb
NWI7Nkpqi9emceSrxu2znKyX7Eobu27rFP8KRDl45q8AwWF2uhtaxPY7e75aYqrf
1bFqhIIh+k57c5wCdjrBAj9h95tbek+0tTmGDchUNmYkDxdFHFnLz+pPmLF5gFDx
0+gKe8rJIJsEa1eJStPzT6NHlE2Z5Xe3kUVY7P8XuzPHvwdJ4L1iosM7RKZYm4UL
ep/HiPyQSM30wv9d3WtAPN3TBFvEoh7zfn7PTnSgTr38u7E5oOIzWAihNiCLKOa/
H+fNBfIG/4fHdj6hQ9wwUHdi6ULVhCq83jsAp/ttOV7nv3aYNw/DlCC9FLV9XS2d
M1K4ExVqGhHncF5Qef7tEYx8gWRCvaJQ5BtYkYa/3PlL9qmf1hGH2i6sp1nUbMTz
1zUe0woKXpjdfaLK2nZMNPE03AT2B/Ejf2aHlvqgZoAjQOykyi4i5OFvrHgrUiMD
R3+44nFsunxu6eFy+EqDWYpfyhxXOscuTHEHHgH6Xv1yaT4ALJNG0PMTvyoD7Zkr
GvJmCxKuKQj3gYK8DRoGTwZsPkTlR8Y4tMbeg0biNEABcGQDq8Aqg/ChKqqMCAGz
qQUYRSRZueTHP2UjOmfgYZ7nMmw5Nv/HAYhARUmOBxZDPPaH0eGG3BvUNpGUH6cS
g0vI1pSy7axdSAXR7aJiLHaSH5SCbEPRtUuXN7VZINT+dFev4VR+vRh3V/hVDsqQ
cvg79rT8JPQajt4NkAR4MH7q6VVpAJ3zQD6HH1dWfg1Osg1fFYmgfcFDynP5jNCt
Pxt9m7jDefBO1x7432JzC7kM8PqWbFKnGds65yydO3SI7VcgYJidXNZuvVvuQyPd
K255tIhs083jjZWZzA9vATRHUCqyMIMWssoM8IBZZtw8ncka3xRhfDFiyAZN3Rb2
7ldD9XLvD/05vbdz9RtscO+uR1TkJUgz1ajrFJn1MM6mSVaPB2o3oBzgVDBlBSYk
wKZqGiCOe05f/mPQ6hmr+4ePtyu/5ZybOBCDAGbHx10EtMbowTTyoRd7Xx32cTtb
fiFbfUTkWVQw2AC4gsoXSd/SGBmQVBlUFDHC0RxovCUKgPd8rP5uM2aSyCfEZ3yr
8V4sET2BMPTsEaKDDUB7re3MUhU9wognn81yNtTyXroFGw6jhkYcxhv+SCHvq+0J
ykzTjLAgJEdn6yGVNcUCCTYsyk76cS/MVluG4PHvxG4POjX1WXnTJMIdaRUZ6em/
hsa+oUmLwqRL/ehEuDSimHwOG4KaVuevQlYeH+1l3KVzas4awf4ruP47p2pBbQ4D
gkPKIa4uHvyP4vslJDxdaNBpNfc7+uYkWPQ8/FLLslYn9Xlc/VElMkgaEv3rDjx9
RYGaKbjOLu5e92RQj/49hzUqZwJL/yGNzT+oUlYeN8ymn5QMC89NXSduhnCnKac3
wJ7iXyfZUPhcxUQh0dPwauaQYbJ1N0uQYGqiUywsIZJKmqoz5s6OwI9K88+176EG
9TqBrJdhgzNjWzzmCpabmtU3bOQ/IOVIAcFmy3n2hi6tPbe9ekK2CrLuhaHkWdfv
WbyT+yDZGEHm8kEMijKrN8VnasfaDaKr6Fyw8QBbAt9KIE6FtYppL2OjpU5w90ut
DXqLsG40G6n/zDxPRAUSMiQQme6r+iGk1OqcUUo8pRglPnYk99eIUWQRpfgG3mpm
Aft9fBdig5Q3KU2fsRtxkuw8VTeea/+v3++vlzC+PlZ4nH5NdBifTqXLdSdvlmSG
amR0jbl9hCXioStDFCYJVYPLGFMPa1S4d9vIzVrZq6NMrszYsLmsod3VOO1ldMHv
w4rZhh1crvQjO7Ny1Rcy0B+WDNnQQVXilmb4mXUXzIwdWLgyJInpiW1XvIZL8piZ
akYYnG/TWdGyk3llR9kewB7aa/LZrE1meKiAJpdDHITM9V6w41FqLf7ZHsuZkghi
qp7aTJxiTIAHyf+xP75Ey/hSacHn2D2TAEtriQZFh6XgnFK+aB/AfNQpvXT/unWr
t+lwhwaBRl8+9ZtE04Os7OZqu+GKY3mjRui+pzhZfS4KMuqLCbdLUcxYb9z54eq0
RtyS6SSODJCHTytaST16tvLcs/lDM1u8VxzSvkZlE7nY7NGGVNPtNEcJaeJIXkvO
Zm72FWaVm/QnqgcAnjaHVD4uWz9IXgZxbJs+1nSUoYeZZfkNExEOEnHzpEX7xyEC
QvXjyBCJpbd4AaUd68tRvPhTLyRlE2a4nr3bhxQ0V7flJuwJ23+pp1nojC+MvfsR
hZbq6TBWcfCAHkJobIFS/RJ+/zLipIiH6EI30X5zyqbJQwsCHVXAeoFK6CQi5Heh
uxfWMO9QhMt+xxqLGFIZG3dkuBSL3sPcTpTgJ8jcXKZpgjQdQzWdaaUj3wpY/Cnb
cRbN2EpzXEkm+vJ987n5v297I+4uGB2BEzco5jQ/N6EmCzqvriV2mfFv2SolNDf3
ZgFfU8WjJnh+y8MJpQ/0fx1a4rJzlhmxgM2CHyNwBG1bH5q/AZIS8hg0uZdkuZms
eQkxQqQmW4mRnwXX+piyWZStbnRHhjwn8GZixG84XPZX+yfRLzMNJEiv1gGjmtWM
Ewgeg6sSsWjDiIttfekPJxHoxqc94uybNqGCIGvvqE5SFdR0XlUg1Kv00Oyx0rBA
Fc8eTEpcv7GsOkXrVBoj3VMQjRFjkOFY2DNmacDDL4FTAKLxHbkmDVdPw7QkqIJ2
3tKfAk0XMLGZDZx/p8Vc2SEtbsufRWqQ5hGGYmD0GE3gYkokQEEdIhYS8wYBTo+O
fBR/rmfHBlnzu5KdgeecTjAMt+J6Jok03hZSi1FV5TCMWUb3dtaUaSmCcPzvzUi+
HCV+OP29aFpkA6T3kZWnX9K8we8nAdpwEDaIwhRKKIsCykgFHsCWvZwtXaINrF6u
l4D2+cMvAS6Ae4+CApa60sILxj9rt6J3w7cxLC6wbfDKU7mGtq4YloHcO5UgHjxs
iOPuBi6NIO42N1pYXxaAFRGtlT2Vhcss0EMjeCz731LZUXr1nZ9bb6vF/n5L9H4e
6BMCseXYTe6cqn8jyDi85bnH3oVqEjboXjkzRBDG59Bh6YBsYb9UgV1z64xGHIZW
zOpjvmH153L/E6s/lHnjtU1RWUGnCf1x97KMNJjZMU7I75tVxqcpHcfHoY0pT9NT
m36nprX+JtKZ6Tm0tl4TWROX3nde2Gwb6F7nf9s2EWyNFDbz62gBzhtMyOajJvHj
OWC3VXFnbuWrizTnR1B0sGa60zapzljl8sN0yqMK3DoqwrDINp8RGZi1kTFMqcMa
s8yAZuzZ8AAx8S6ew6kRC1WAiYCFkG0MozRcbV9Z605wWX6IFkNZvajvHwQveOAY
z1R/p6+uczdQ3a52PVVfK550WjG16zsRzm3khZxhHEIFxxG9IYPbB84MKRf+/k3A
qyQIcogh9CixDtoM/R8LlykJhvd/wPREgmk5BrZyl3Rqx3UYxL61fuB3zCncNlrw
phloLzwFUtp/1utoEw4srQT6E/Nx3eLzWd6r+YWa2mqK9EMasWOX6NvTCD8jN+n7
OvzjVEphG5Wa+4b9ji5gkE6SbHlNoom4QstRHeQtQKt7rWMzhLdvD6W+s5It3tRf
tNJySH2nNSqiVPfVn2QvIYTAGU/+yhr6iQE8/wWhQBdMn8jeupW+UAICvS1k8Nl0
W2PdpXRhSSfKzkcS7RkylMEnmFGOFun3pMddw5a3JDLsprCJnLo0UCA+Xs+v6SGZ
RALCWlAl+xdQvDN+eUKi5NlGiY91S808rULZCMotYvfRarX+9nV6B75CKFwqur3M
0w2gZVUWNfy0Nq/ZbLZxtUaqxB6arB3QLZguKg/ZVJfvTkI3Q0YTfQkDG6wW98qh
Yy+YJ5+UPpQ+unne6c59SeZs953/DyA7Lbcb2P/kPw2Dd8XlB+nRKi/34YHYYe3H
wDJwyZODt9uRDhy9dbaofQBlifnQ3MUQQVlD6SgukUXSoY3SdPF8BpR+9b8IMNsZ
8OHZ3zp3DcWTm2Q0yVIX1Ur2G8UkOyUiDWYc0R+iE8OEE9TBW5zImOmynTSLEuiF
3kZmzcRsDefyNEzl+Fq9rfK/UnpNlF70OrFTm56gS9WP2g3lsbOT0HhkIfwXyWSs
maG0wpWtIoF1KJl8O1mu4XbKvh/+3mS9aK6nIyWy2goCEZ7mRDvqPtKGpKeOpUHa
OftPnRyu4FD798/qKdKNdRLjtiV3Zcnp3IZj8/z8OX2owb1egboc2xScb+Di36WV
fK7IKZR3r95SawyasmJk+BsxDlYdJBYa5zfxKvlK4h38Rf2NrS41alyYB5J9AplV
wXwZQ16MPvgVOyc10Gn8aA9T1DcSb87mKpFUzPQIzf5Iam3ZBwL50LwJCnH62d32
REtOlJ3JxcGgCqvk2J2wm6uQFMAQqsiizu54DM7vZOyaUwe5O4IsY+wtSEoZ6lBv
/Tbyy2iAtgh/c0puVM+7G3D6Q8CEV8CzphXFVSwF681Ee8KywppOkkPXK9htzePr
jKBNwC//7vElF8BoYO/gLE6JtmftzjEETTK/FUHWCx9TSuHDLzbplq3L3Q7ytytc
ZBb6nvN8pYOsmUyHYmxKg3dgXgVY0+NVzlERR62ZxWsZD0TfVHGPbvqHrLii2lT7
w15nTUbrhAD9H4fFzYbeXgmD0mXRsQfMXuhHMz9JwssOZSHI2XQtSxYowNIOmIWF
msMICjrtAVVZx/C+rB383TCdtDvaVOrni37Im3YcJUM2tCEyLYAMI3XqtLWYhuhh
iqJRe3VLayiAq037yN/4trdpfKpB4eiHWWOU7N5YAIUY7qNKg9H15Gx7z9t68rlx
9QujNfgX6RrAggIcZToD8ALBg6Zv627o+0rzrpAJl922E4WEEac8XZrhLREEAq6+
ubb+cd42OM0c4KId4dV+SCz3otxDCac4ofvScjmJijO8N2QzWf0bZiLLqQcTkQyy
tbOxpqkPR0d5oRUM7SiAUSYMA9OBAN6aNKtF3CtwgwRTOrO6sarszmiuMqGAGJlP
Yhqg90oTQDxjYn7tgeTxEV9gSXZ8M+oRkJp7N/Iwq8hPbJxIq6/PjPSlGvF3LrQx
RGOKG2R2PUfm/a1IxJhQP6oCQ4tzDG2tCHvf1PWFCKHMWlf+hFilqi+JmM66XLR2
CxbpRtc7o4KB8/R2rbLH+NArjfEiMkkWX0LVT8p/YGg7DuDOAGr/XuPNo8wfxTWz
GQSqxHjiIcI5/7vNjfiK7z/TgXSIok2yNWOtwXWakTHfy2wEDaEO0h7AmCuveh6o
L9sX2MIRUn27vYJ/C6maPhrCCWZXNZgu/KjYAkuco0GREyV4t+CqAz4iP6B3AGrI
qIPI/Rc64wctelLNALLyertn0VqX87EHUXxXmMu2ZGdw97id6mTS3HSo8BpdgAO7
MapobYpCeJQb/ZYSl1OTxaCgN7u0/TA3FVW9gaoCBxdYtLXWdjpsQ/yWELUOcOf6
Hweq7WyP1UqF4XZUl8kqwtWeBWag64QkyjjsXukv64a+sg+xxdblEiUPQnfMlz/b
Mcq+9r17ZO831pUFiIouaYR0u7EqOAMy/MtYjjfoHTykYNpN7nxIiRoROUQS9Qvw
CM15mIm1+zSsZTB4Yi5cy/jculHecZk/EowgOtgcn8N83no8mFjVSPffIlZJkxAF
1aCu4ZjdqAkZMeMAz/pAvM1lALBg4AWyBTEtoadMtLG3dhBvnIQI6gi3ZQLFclWF
JuVk1IpRoH1ItiHaoOecujG6iuK2lwZNV0ZbjuTpNd/dbelZ++7WsYc2bP/OHQfQ
X1h0ZQgLATObF/4SLnTbI3F8FiQAjR4Ie09WmbAO8u8NB8iuGXUC70tVQWnMWgrS
0USD6vu4eYqAGr/ToysoYJxjT0TqSq2JaKn10jSvbmVqOVd5uo5WIVwmK9Qb6yME
ecF262jvq1OXOkw3IYtMkxzU3OptVfEHhmIJUYZ6Ny6HSaMkpe3fbIcGpievR/7m
GpC6CGRcXDjQNLU1DP+aa1xWa2nxsONWb2E+C4vfC4H74BS4FXowrXVaus9sZ5q8
DM0EljG/J+T7lAcm2LwVyQYgFAl30MfEnNmVuFtMdsBnfKjetz0rT1Cn2G74Hr/j
6Y/OaO8fYCHf0LG9siSQNttxGr+6fjCQMaIOlAGEz+qTzfnAWQpWT6g7r3CQrhON
k3eYfP3eLKqeNLW+Y9n+k1hVGJKekTDPEUg1aUqOlcqwMfKR4ZtcBmMWUY3Sh/NG
uWw7uOjEq7ufrM7OMnGUM0D5ME29VCfj9vZsQGQ//c7mhI4I5M0rLeE/FWsDdw7y
lciHlFcHxylAfT3JscLL4E+1RqdVgJm2tUVg5W5DcT1Ak0ZROx+gxIMN2Tw81NQ/
f2r2s8z1DHtc7GdUHx96Q9BIOVfWtdxXmgcHaOj3eAZiDIEmAMJM4OguKtTTikAS
gThOgpxOOlUusnvcm8Vob047qDwYQJS1W399vM4sOcu+eRIcwdpaCJBRa2nXjoik
Z0AHmXFDFLTSq9ySQUFbi1w+dfvVkfEYHn+dLmbALetUvgjm0AJKO93vr/4CowtL
ZBxwvSCac1m6xy2vjZ2vd958dJuJ2cQ03Q+LrcdJz8TZH9KroI4cb7Wyoo2E3nf6
Ewtb7/jyIxoUiFHkrRPGSBalhpVo4rFxGIxztsoEVUFmDDB+lCGEARYDMA0ku86u
Z17oWETZngDnrTIEzzfpxXmKh+hpPOEGvQavzWbVIKIWht5DQC5X6hxDaezIWSMo
VBPJ85zj7csIlF2Yyokd9o3d6jSiICIqg23JCBuhMwQBbthnQgBmJPjtgh2ewsgd
Hvr+myhGq8cDjqWYZHQvZ6naQXgGbrU4dwUL3eplEZzuPWz9QaxBa7JDd07a1q8x
pxtC55vGoBx2raFy5ROorzIXytv8xccbgF4C2VjOCaiIK4ucNxJ9Vs60J/upzGse
Pwntuh2uiANrOThg4xx2K+ULKmH15XUePn/wi6c3eRnDwNVprfl+beJ6v6YM1bJu
jbs7CE88hWltkLAk5KSN001AWyFgaQMxuxbcdGz4goFNhm+jzGSND6ta1oRULLJ/
IsopvRjHzu7SoLJGCfGnihVyck10tOTNW4mVwhIjuGWNIcJq8BXUtZJi3bIEgjQH
Y/TToZ8myJGurT/IAQsCNU6akwLTyRGHtFU7NwAXa1RFq7LVQbBMMDSmjmTDuLeY
7510utq0hFgquX3kx8iL7wGClnxk0KzcHUCjXxzw4wYQ6jCTriukYCT5GGglHgtR
Jtms2btoKJUvpw93KWfhophlCA+dyHEpfGeZhJbrjGBAPy3tI+EXSDx6Y/KTodt/
iAB+sDeHR75Vd7ds3rZCpFRXUr403xJsAgWub1SPTvI/MWEdTSHjnPPCTvxm2sFE
r0e0xvHsaRYqb6Sb19Ndz0ohJSlO2uPgxXKmmiIxFAAEPsDFOV9/5WFEAQV7fMi4
rNHVL3WA79v0NvhXiXx3+MtW/JJ8+Z6iV+yjL6W/i6xnlbJsF40ytIUwzsY3WXPw
JbIvB/PPVROBUxCmFZOP7VlCC64zyiwp0FD6PAOGV2FF5hqEGa3QH0qj2c42oaH0
x/4aN/eJ6C9PXbZvqSo58yr811/XnrBAJ6kaDpRmFsy5+CGCj1mHBQGjVNW/lHQA
2nUrcWb2NZHlbMdSosKnxoseTpfZQy5cSXbPOG6nzkRWdznp0cnnSJ3gmGAE09Ee
/oVVeeJP+3qwd8C4pNK0LCOUI2Nrq3GTHVVqqy7OoEtJaA/1F7hj6KZsmARnHsMt
vaKpCRPpEGlgG0KQ+pzcBBV96gPscplZPlCH2uxEE86RzwMMGE/VyhjwVkb4/CwJ
+0cNCzyv8YQ6oTrfbPI4UPlc2unfa5/CmQt/Z/nzK/lb6Z2CLuTmlDckw7U/8YE7
a1xwr14t1BPQDY7REDasUfxIVUvQqpBJIzzON170RgSnSxsR5a8UXCIz31tbQZYr
nBkSXSCPA3l1jRaeVnR9jcm1dEEjcj75LM/IsG2p59FFjGBy8ylzTEPO3Lq0iFF6
f6AxoXXTkd/rB/TDaoeqH33jYEJYVHVuJr/UVn2CfXMxZ++3rrKER5ytXB6uv5VR
4k+bDYIr+8L4E0JJEu3hMhCRMAj2OLOM0Lnz4zYwcXPBfK8CgD64EyuxF3/mjcPF
h3daXxux904dVcEMwBQXnb+WnxXydzN6EbqDVqEVZsAa5MElJ36Q4oAmAy8JeCRX
u0t+U13x7yYzPmTY2l3gZJhLKQgocxhMxjMC84m80Kz4R1Mb+YrTZmxvNCwxzj6j
Jriy59QZg3WDgkeLBIBOag0VLi8toThb2ohD9N71uflwBxDYKPS4qdBROhHL52GI
lx6CMYSxnijXPtTacVVrMnr+xV6u57vJIqDjJ8EtiRjkC5VpUka3Jy9mEdYdnSpY
4BGegH7QmZBB+lcwpfryNbWKOn1NzDzbh5NSmNH9DdLnAp6wLcV9ovVtge+VmvkU
WNZU+DysDwIul+zsH0oAE18LYbaANFIIoaXFJNhTX9mb1L78J2bXU7f/U8MRoVah
5BWnZSPQkw9whZPJCNiVH5po1ms1r7vbiDux3RoMN1im9SjWsD0ePOcXZVeBVM+p
ODeCRGJ914+FiFrb3KIuwfDCcbds0R848QMkvlH/GAozWHWykb4Bf6XxAJqUV9Ks
30BL5xWLmL17kSt8hI8mqbuT6UFmUzdp0FUn1/kxoQc5/S4VO2eL9r6Y05f3H6RK
8E24SP/HmVckH1woR5pFEVUSQ90jJxfzC3UvCUKNwD0qy489m0LaUkwiUrSiJFTK
4X2M4tCrlf+BVQlDLg7xs0S97pMd02u/m27tPh7ODw2HBeZrGCg2VCHX+ksFLQm8
RIFWZuzF/7YUrAPYU4oNyZFA4KOmtV7cJAS1uWzEQIZzdZJTF6xgR0UfEB3uNasG
sqRvwZ+ABmIilM4g/kstbC4NJuWVyX/Z0XVGaaMXLj4IbNOt+mdF1NTS8ry4JiCT
sf1bUNVaoKf7N74+ZA4hchdvFEQsqDmLnall+rz6tWTyvqlVgVyXOd4R+pCg1Rfz
uzoOYByI4LSxKhtJd2WW9pOqqYKrFl75/d+RrKm40uF0llkWvPbbpKze8KX8I7Ed
hCky3UBqt2mo0IRLutzbJ4sKpPGWgcKMLSEAJT+ocaciR+3IVLWiDeQseLbmF9xc
LD3tcIXZOxuB4xBnQ3UyumzTnL/Vv3g0CMgEYbxuyHnjxrRCAipiL/Vzd71tFk/5
xdENNOwBvKpJEfVZdt1zv+8lVPgY1b1L7NmE/LYRgRBiTstp6o2PbsU7V9/5k4nn
SuV9UJl7cke+2FrxTPpSwIY8WmXtA7QujrRYiLEcZMuWOZSizM2vsdrMehPjUUwz
VjRFnK+dR975EtFqa9uPQKBBjDptgB6fdtp14QJBk1KunznwMOhQZvAHw7/TXOup
GvgXPA3LVeQNRwg//CMdkZ2KOBM/WzNrzCJdiFYLnVQZzHzS66L2kP+qY8HsxSnB
q8OmSVgnKvzgLmnzPf1ah/A+3mU0aJAbtKciBn/JFs325gzCux9gSTLqCWfl13Z+
1vRMRTPn0lIkWsmUOog9s8uuP/8vrNNXbRSr1HJoTztX0jQr5PnOL39I/soQd/XK
ZLoKHP96f5TQxL+l8S8IUZj548zhs8hbXq2yOF4X0QtzXiB0EoyndN8xR7KF5Fnx
Qacv+fO0AoQxH1fZ1icb+hjs2tFZhl5AIVCuP/JuNis2d/38s0LWjs0hExSWeuUd
BUL70HmGpUq1qKTn/VJnu0aDSa5d5ssd7Obtf0bcUCS3WXIJGcPvuRWRh4SYBMMl
w51eL4ssId/KT9ssKRckguIwgdrIh2VDgLFBesQJpKPijs7bPHKk7+aMB1D/Ekd0
iWGkGDZMNg9qG+agpGNnYd58tgzKqqrswG/Xx6cBV2PAUBcJ0DfwZwaf/PuL/NBf
+n2i+GVJqt3X3SuMDMa1elKTLjvB+ClZi5z4O42M69rF8WOxHoTpeDwjxqYkCdfs
oSng6zOb5PV7P/2Ln+n1oHr9tlu2blNyF2hux61T7HBIMuGXLTUQgDLyeDwy/of0
kxswm3028NzhtCYbILzJK+MCN+p8VdTVcHEoAffxehxN7HEiVWelcYOdWBxyupZa
k8uFImzQBH5f1vZLYWwzCPkarv+IEidEHt7GAx1PolgtKUt39w+oN3uZynmt47rp
kEcSQvW96xw1IHiswRieXqgFb4AeR1w8T3IiOmurJmVV1cFDCMMud/xEFaiG9vXM
JloJk14vVibzbGaKBoiYFXYKhtGaba39z/+6B48npCMMIoCpgmMtJATf+C9M/rKc
2CrMaP+fmjyZtxEHfse3XEJiyv/brEUmonbXGgmuUmcuGEiVirvp+FEQys691Oie
m5u4zVK2/JXWjbhvbeUY2a9+dpGnWFqKgjRc5ba1+jYyDLZMHq15tQyBBGYR4PKz
YWlKh/eyvYDcpOqW+VjZJtP7OyGaM0jfdpQPBvWLX58mpiS0s7lQLoSU1/G76OSm
HPHsSg67bfholFI5BCgn3TToupXDnC9AMBlvJs2DTsgUrt3KXzFnR7JN1FCmdm/T
J47Xo54lDD/KjQUUdt9wN1g3P++0U/oDdRMA8tCufJOaJbAqoK6UBHMXJ0/WzBaW
PV+RWmSLLdh3uqqjA6XijUU4KzbWu2VdLSD2N/M7dRVf9Q50fn4zMjdSN4xgqG4S
yZXuIGsoyBkh63SQ2GuBbZWtumaCFIBBomiuXkWjyL2sEPjc4nD20qPX8DmulnEU
8YpbhfP/TbpQo3W0B8+yXnf6WBAc7xmXzrBiQFdZXQ3uPQcp9pn9a+d2uVZI0sdL
VLbk9p+jXrEmrLll9duqu/0bW7R6ED0kHMOWgpvxLFo2EWJKPla3joMRixLFLSav
cIrC51y5heg9/ZqUn93ESFco/AO41bElcAjojkj5dkKs9LRzJq4A2oQRSFuIlB+a
eJ1lJexPt1clkPbRteA0bMJ3CZFJ7wEQWXHhTUmrfXx64gHZcuRzsp4GDVblJ1kF
ZHQ3g8fxATnuz2m5w21BLZs0sN0h04dX0ArwWVfSNQv15Sql47+s/N6PK7719sLu
uwNHlLuyFLazrB+iQBtYLwF1yu88MaerYb+rFLGvpyvvtEhMEzc3c3m0Xe/9aWWy
C9c8G8dik950C0HZJ+v+V3HvLWGKYrTQVgDIcPWRgGmIal6f3Mot6ye0/tQ6nkG4
VGF5S/o81qGKvJo9uEqOCgTqFpnN19g5gG+HEiwM55CZRMhTvUo1u4inJAsgPU18
hAh2Jz9vR4cTPBAofPemjTo0OAmFrC/tiDEbYfCfxBvAeunuN/28a/yUrSLMBIy2
LyunP3Ykfd39BNuQF0LLHKxQVTgmDxtTzrLQ8Q5AwZekVaHtRch4jcZ1nY4dbqnP
3fxgzK5I0NVTZaVpI46ZVLByIt3aAX328u3iLvJTBnKIeJXjgo9K3343RUZF57Bh
w/uoe29siU17Q+oJ5OW2CqQ+QlE969UBDFTXxF/yZ36TxKVh1kmjQsxL13TqatHg
ZVW49TjUpwAhMPoMAhaW27f6UlQiyZVR5XfhUWAZHvDWuz77qoTKcV3d0zGQvFQS
7V1dgkjdB5rm6x32ONALjTWrXUAb8UEc6iLt3DY7srEy5Sb1+c+sNGMFR3gV+Zt2
bY9vRKxHwk5iFhG33MRMQXSulvJcNL+PRMaJnvt1R3VRtZ35CXYNHBClCxo9HoN9
X5nzE7PcmgD+iypnbpPlckbNOBk3pWJ93fqOEIoXNq1/ulyONveBLJKHpwsPbO0H
fQeXdZfFd3XdJnVjXVHdEOSP6HkdUe9UKpipUHgOLwEQMn+Q4Q+zh5WJ8ejuwrWI
0QubnB3htbDKYVxJsESver3eFkYNaCfvk5QaKDzoWngscYojQFmC7qbv3Eruv6tk
YeRVVKjIakbrZuJc3UdllFREdh0fhVvf4AkUta3uNZzGfZIszokG0fDNVyuZcKcN
iawwGqJYf0Gh9ORN+UPdKEyTX/xshphK2oNpqityIVxQ13MMyzQm7BpnEzgHo5A8
Ic3FdW0I3fqWPyves1DqplLoecDllV3zKDbTEb2cnm3p3IqLickHXl57Nx3NU9PO
507YJ5poLsqZ2aG7MXDWydzWhNH2gXGK5sZU1hPNOZH0HmpEOAY8bk2UmV46kNRe
efitb0Z3qyrNGkw6U4XfVto1Nl572yqLVGzOoy3iuEsrXPPulZwg9O8TBvFJVvHk
0HSuJH16qEd2WvebKkfET5cDZlFe8v6ikJDjhVXXfrgeVcxGDvpWLxaioP40hURH
brFzb8orZ7PZtl3gn1fV5YzI+zZq1GTjPA5xhJgpMPl2Chz/1aNytYLNfXjrJDmx
2R1sLpXJ6UxkWbNByUPaC0tbals9DWiOBcphjg+C0z+xBumNfA46pE4JWfYVKTIP
nDzTn74uypJN++VucS3W82mErU1ZoByUVY59I/c8w0MzXN4j1qBqXfXyV2yeHgCO
YvVPIabTUu7/qnc/bs5O/ZFfq2bvSVFajIi24L+x+IhFW+8SdFkFcdMqkniAJzen
ZtiQgiT2ZTHhGgWkYvockgZaSM3T7KWBGxyNq3fZ8T6aLyByeJ19XPtzWUhnw1aQ
Yh4PX5c3/Yf/hN1dNNbHrRJKs35ChWqYKUcszcdd4uSqs+04rgEk1nwsQCMVap4D
bRibboJb7BfZH8GPudp0FhMpCZX2SewYOiA4M3Ci2RvtqQ6pzr4xkH/PItn4cbvi
f+ACS/3V0PtRnDPfVVlMHWm9LzfSCAHdeevGKLVfo3q/YaQQBHi/xaKM+0rceufn
EU47WjqydUWxBXujRr2wVfm/8y8HdkXSlNPqcQbFEQQi/GZ939TQngl+M4OV1I2V
y13VWGaRkSqjOgo2ARfHtlClaxZpdJyeRKR5j9oV1+z+xZ30VV9Hg6T3ljLSUUyP
09wjBSw0hWPCNydrq8Rcv1q3Zk7rCoFWp7tS/p5emCU7lf7wPQ9lIMWeWNHsq+6m
zGIhTxvBCb7EI+px39/2N2pj77UfarfpxcQkE4zy/wmWqVUAWo+6uOhxprS4lBzo
eaOtHD0eYn4Pindhib9K1U0V72+oIjjWRUaMLZKTV7ktUVcwOStFLrg8yJEtbtTJ
15avXC1M6Yq2yeu8F8Y+JRy8iepHR52vZ7Zx7C/lbUb0HjHbmOR/X6WcEhXKWo5m
NOkOftiy6FpSPc6p8CV77AGBArQ9JFkg5Q80BGpJjmrpDseW3/UnRcc5M/h8NFv9
85BFkgJw+bKHb/MtR2Qtiubt0085uUwrISNiMZS4hTPE4pIDRKiASaMnnFNjUmak
+eDessKIR7xKWnf9p4CAKtXhxgH+kQBRkiJ7RSjifoxwv2zcEgDQ9N5YH58KcitM
4x4I6wpDrIV1ZlXKrfb3P8k3Fxem2lsas+kqJ/bzfG2Hj5vwQ/YGGb2yPHkGRTdn
Gi2+qADefQuWnKG8xQ7/vFQNQaXxN3VQWTnFrKG1lKwyao/WQYOxNrYDDBgBXiyI
cYYgYV2couHq4F4AeAS2nbyO5Utunsk5vAyFpgZUdKv8J5jZ1Ck9N57H2Mh7ojJ3
Rmz5oY/dqe11ix8m3FcbQjhFu3fvYaDzpVCtQ6OxXbkqbE4PbBwWbv4huA/TjDJU
5kf+wnQ/uJCOF32FchrAZQJiQ7m9ASRD2elvUqzScnHvvXCAAo2OxKYXZj4Ems3n
xUMu3hqIc/WxH9q/IJY/3L0wieHW2RUiU3g0oeODfL2YZXlN0pDcs+TVEvKH3Me6
Nm8jUs0Niu95gR7RV8wLoJKIB12hP2p3yJaEXzMPMVN4Lr7V607mzUuOkjel9YD7
P/edgkAsP2Xh8HCGA3R9TZH/QCEksC3/3fpEVYkxHkqBFB6UqA4KCQ7db/OZPLjL
nZaUQi1zSgVnG9QfAL2wKrtu2sHIEG52E0TtVR27Bw5bUmygmDLmEQ2pIZ5e42U5
jpiRf2mubNu4Im0kn6tSmgtq0UuZLRwN99+myeBJb1zxZOPUv3FhtcvsnNgc6ubf
ftLvfbkozfsGEhwGyi0skjinIno1B+dWmPq1lOASe5QESXYMoWrdCgvXWhqsQJC+
d5X5Hmak2iBloKnGZIHTS9gAW/bXWmIqC/K3whjabeHhOsf4dNi7j4vQfqMc6LVg
R1oTnUPYrYQFMAU29dyqPT+PoAK0MgoY5vE7iZhOOLuf3yDgxzzBxhwa3rthZxYg
QD4TJg0TBbV5TAEOaM35aczow7Ps5o8qAo8/rdV1eCTaqavgZTQ6hlSE83/z4HxM
+yCn0tJ/stmKiAN3wk7Lf/XXp0t8BQMX79memqCr8+XCetitDSiB3U7lW9B5bLQ6
YrQTP0sgzdL0jn3xiG2Ga6j+irpxLVbizk+BvCGK3eFMvykL2J4N/9/lRmq9aPb7
PdMp5QW7rXbX1lkWZ5IyTV9zzd4RKLoA2SoSAcIKimHJOi5QdvPyMDvNJ6qujcDZ
AvXkXyoYYOvEzydRL7qXMVM57I9QBTEK0gGu50rByhX1XQNVhPExBUrWVRCCKMU+
UJnH7Faeqleamt61U6D19cCsp3cwC1IeDpbiuW7ZljpMA+sNpZaCJ4djiSSpA9v6
1LlRX7e6oS3zAPVz4dpn64FgXIi62TlUaVmDNzuNAI3Y+XqKTUkk9rXG4yj8qv4H
8XFkgEc4cWfpMPzfnhKXVOLJD7ixXdhb9IQ4sCvjMHtbQpeuBs0/O2vUOC8qK9XV
W1gJX0Av8qju5/qPm64aqxIwnsjyYn+8r6vSPVfxT90WCVNsbo8KNw7PAQfOGpFu
skotxMjVP/ihQlz4q7iu/tqQuO4I2iUglQgw7rRYJdFcfCRafUAIutjgDIxdD2Fl
DlvttJHPQZU0MuxXqBtrZCgypNW2LUdL2OOMoW0AL8mvvYGunvgx+JcwI1WA9i1O
4NYoIqA55ow1+btWV8VerZvwH2niOLzqvpRL/HN4RHZY9f4WOX/eymVtoW4Uk1gh
Arw4GnuuCRSfST+JqcFsWxl+UJppUODEDyZadx4QtydKLZt3kYBbMop1/A+D98XO
zT3Pm8+2BnyDhYA6xByyHe6tubbWEXaG9yg6qBpW19rERaMeWYNxMonikLp1hh6Z
mVyXPPRXXCriAxcP2/csqRGrN2oN1BKwmSW0QwaC4CWj+69/sSP0+8DfT6nF867B
d+E00g1dddPSn5017lCOcedHVanj77LJJT/FbmoNUxzj/EPfq4KikJFcCGLCnXdI
7MaoJ1eT8rtOmKIQ5ykfhtXvunMCVTOLz39scY8i17HOmTVzjeFoGHlZmQ2nhhFx
dSxXxNLD2MAI179UVGPLAkwwO3iLRPHEN0sKxfyISK3ZH2LWU6eBRl1Km0b80b1I
4vi9rkIkabZX4U/1Ra8pqVP8gTu++ujBcFd7hK4r06hjP8+/9R0B0Xf3EQakkJ+7
YqMKN7uXYRqkrPHInoR1Edox5cnAvpm4B03msF5ciEDbS65jrHQ6y3D9AcICYjJA
tnnJv+y4LOrw26HeTLHK8wh/tIuVSueEKBplgG6JZn0jo8f3KaUk7uepqrHgdkop
x6Bw/fcOeHxRQ3YHBUPmCuKU3fQL5WmHRsHpUwTEOBXhDU3RI1VvoMFa+Hg4ujzv
DpnjUs14lZ7Fc9QcB49tuCRs63CnjVWWZiiUdPRoyUGFeJPt6yzLue83lzX6kRet
dLmHUOpfF6+5QmS6REEuU/spntzfQuRHD96JI4yN3acbBUJhLMc6aPuGpAQm30eS
HrFGWtDXLFrNeuhh/2hmMfyKGwxnTq/XtC96337Ee+sqTXn2Xul1Jeahrg+dfWeN
Zlxr3+S8HCAGZcNKWi9RioAiRo4ZknQ4C2kulZK63pmn4ecs7KcZ6Qc36cYD18Wa
4Su45KIhQXarUAqMRQ/Q+lo5yD47wpwFLwyYqsuFTTGn2ivQWnVSNvaUsenHhFVq
clt/1/Y41ZIoOABs3PwQk8XhyUz9E30QvjKGGpAFV56h0jXV5JBHTkD/hfN+pPtE
wIpLdiTdXS/1DyI11GeRxQTWVakcEqXggUaBlE4BDpPo5gcU4/KT22+87O62Rv5V
ibD8851vTdtM4Wo453KJmEYynfbfOeKTo+AEVsJtbWs5RQka5zOv1/WLqeXt6kUx
26qW1KHzVvolW4SL7Lmtf/p6bBMMCkobMGncDwnXkVC5RfNLMQkEGzcfwyxvv/dK
ds/RXEzuUdzOYKwoaHvs/NNUSfydxIfeO3NXsJleHdQ/0aBMy+g/GjWvepqxFAIl
djIEKZEoBQDi7gnayywpXb1dDPs+K15hxDX6oPr2gFwzfGvqa3iQCgrvifoQ12tY
UyCrlwnMPLUdFjJlQVcF1dfSGRYMVkUPx/r91glAyO+UbYn2XYu6pbpDW3GNIyj5
VlRkHvQ0qeTos0JGBzJ7vvfRnzaubGX6aW69/nWu0UrEEFQ/3DTpcAHFiGNXJAN1
MBZ12lk+chDGI/hYTyiZ86lPC7gMOg8likntDZ5gq9bTzJ2i5Ir8L5GLd75PN7CO
FaPIXcYN8NdGxGJ73ydLcqms3X9BqPQZWPk2VNc0WORHKAhMMMrizBeXGxV7dW5J
k6NjwFHQCL9pyrLMjeSYXxh6DfP4YuQVlARXYQ6h3/vVaYRB0GepaVIeI7yFnuvy
5jS3efZ154HWzkEFFo4+ubisqyWuJqYkbupEPxw0Op/Hr7z+Ddz/mft50S5FdzKD
scM1s1xrCD/pO/G6yODVYv89/PVg7UwdOSe1i9fFPLtpOJ0NettB0+Yh0LSKQhTS
ZREDaKf0jfF1g/C6MRbf/txWM5HXQZbd+MvKSZrUWkJnpZETeWwNw1jm8+hagcoq
v2qUtA3b8mg6sc0Vq5o2cQWyuL3y6E6Sccd2PKq0hNkeFic3IGqfbW52SWLJxa+z
unsnwfXWX40irH7qvSVaVlKRo4po9CpD8M1HE1EzeL/nRFn1ZA8syYsTbHVkT7uK
HmT53hYIQthG6DUQS8kLculqKBVtVwX4d9Bmj6mp9x4U1YryvxX3wn/QlG+c9Chr
NGv27PvyLdKZikke3UyGf/Igkzw4S3E5LJBDpwG8w2Z1ElxtqdKWmyw9wdD2wMrD
OUlwYQ1BTMcWP2Jc8q7Ot9gBzxTJ8NQO+XCzKzwJws0PbehQ8Bcf9QCeaHf9APjk
pXJdvPU5b+UhVSflnbvqd4lJT/Ljaglw7Vev9hYKunmNL2PifznMb6fV5VH9KYHY
1MNUSgFnTtcWn0zmK2G4YntFPt9u/O+yr7tWxhTAEQ7Q60JgHGcNZ5P6jp8Jxr7A
doAeyUjmFxCjkoZXVMYuohD7QBjTegdMjX486T5dTBRHakL+O6P6IWcaJiiLb4A6
7uswGWKjqi9hTr0Go9pS+bHdG8pXOZZO6hsdIYtwBYrhEO0UvOQmvTlaSxShiRTj
3FrJJnTTHjB3x5/hHAvrSjYivYMrPPTlF8twSHl9gdKszuCFWYilU7IXP3QIdrmR
4uFWFxMNc92bsdOY2QYPpsNSDuOkZIAgSiT8iEU1JSFpwjl8O2Tmyq9vg2v6HWiD
LAkpDbJPdWwXiK0Hdzdzlexg3rUhr2jguoskLHqUAUKtWGXBfB5oaYY8beGr7l4l
3iAGdCRwebu2l4diF3TEGtvLls84xjssP4XFWDzCJ1sErSoVlUnVUacbG69hqX4/
EV5MP1PFRlhgs0sEvsizA8Wa0i9LClPqBIYMFqbvr8YI3T7bmTxaNSWqtDzMM6oX
OQYmpB40loIbwuRQMbsVaqhqcHVhavNv1FG0YFeBgJw/ewwy+2W9Fh2Z00kgR0TE
X2y1IlQMD2p7ufRfFHI/qtWOFac80a1llUuMqoe5an5YiTk2QZB2ag5cLJCk6g58
s9o/poskabVeNBGjtKzKnkCTLvjpLCYUMc3luxvOEu+VrYqAs6JBuvpvIr5d3LyU
lGOdzkRrCbIaD6Y7l7BaWdsP6F4kC22tb3eAVzNjOlwGDgx9MEfP959CpsRwWiBD
B1FiY+SoRwIUX5XEi5/ml2KFhf/QKjfloM9AqcIKkX8Ubj691uIjn/u0z4gfzI8g
SVmcBWJyj/aq9/I+m0ByUr/4T3cE79FSprVhLzESVdQOv0Fil0/5YSKCV/hbEj02
MM6PiMWuP2/oSRgq2bZ5zQzkzJAGH/kBxMrWQpNaje0lmiI7nxFzHdrdXnl48kK+
BYFg/DuQqqSCA4iiKTbb7IQTlxfckF5g/DeqMS6qfIBRUasyCBGsTUttsBuHNtUv
kCfze1SVrf0oiSvUYtBt4OZd7MLqGF9Bl1XH64oN6chw3OxaQ87uzhfG7tujWT96
eHs3a5LJmVOjepYndgAf67GZ16e4fOzn8KDsSC+40zU73GYuJKqiupuJQRS7ZH9C
tIogqlgsAov82G6zV+hOKFy880mmTdw4eEXY3lnYL/NyhmePIn2v3ICb0EX5lchb
ZLc8FU9pevBuh5UDxIwuTDZRdip+vz/2ZJI/vrhD/nhZgQzSFFvQD3QuI1fyQaWR
dtHJsp2Yz6tKXklBL7oZudyemhewpdL4wLhoK2rjmySWp6ltSkr9Z6ZqhvFTSo/s
xutuIHZ1/TzlpOFAqOCJYMAi6Rlsl7tgo8cgM3G7GGjly4SivAU9+2W2Dj6ueOL5
YSX2DNb6EzG8zD3u3+2zoqRyiQYlyrDWDTQsIINQW4ohP/z0rE9xcKW9wjOlkySI
MXo/ko76hLozlDkwe9FnZBFMcjrZEzBvlVExtQQiYCtbbsC8NMfbcNbSXF7uuDgv
7rrT1oz9Sv7+jVNS2LBnM20GHPO3LW49JR4eFJe9q8ZvVAnbWJ/EkGFibR0JxYK+
4jx6+z6JTkPYFlcpIxvBgc6NsOaJ68fIzX+S2zyeBWrzkM9In+SLU9+0K8TNKRaB
2v/fTxl2Jbidb4lpavzkIjoXJ0JBn6h8IpTQwcD5Q2Q3C6BThTJIgLSbAd423T8U
P42tJOGNF4nlYTfqIaNgNqXQkmi4PxihuB3wDgep+pthNxHRn0XdKeHbjP65R3Bh
9YkwEjJF0CqpalKn5HfoThI+ZIrx/+ncFZMJ+YkcogcsPOuOIo05Jn5fjW7a2B9Q
1skVe/oKfux+lUcv10VG9xGpMxDke5DusPvUUtSspfImVrUUiUtySmwuOkO1GBAh
7jfOXhDcXCdvBw6Kxl4pCWkv7EgRv//rHZ8l8tkA48Ulw+MElJkB0WwxC5KS24UW
eT+mpv0OlPumf0okbz3O7V7wkTYFgoR2V1I+uI4/cTrG0tE38ZD7yaqzAQi+A58W
tuj8EOYNbpQZAmudrIjNpCOyNrey9YL3bkfvuCqSet7Y4ZvawPvWzk7ZPrfS2kQ2
f28CwoE63LUkS8lVHUVKz4b43XROOE46xwKWxcfOxN+MOSKK8ZKh66N66hBi7Xut
cGlx6ce1ME4/oJsCyKbKJqRA2iNaPhrI9c7EeKWIYKRolbec3p84MAbxrYpSe+io
3F3HGnh2nu3f3LZLe3POhddBlRwbkA7iJvf7S+8h0JTqtyA2dnNe2eMxD9Xdx3gQ
y8UNG6nVNPUA7zNRc0B1rcg6tHetcJIRekgxcVdUpH/U3FT0uu9DHCDS6FS12CC5
bqOnH2gSaZvJ+KAW1VBrOtlA4IyXFSOX6Uiyfcd+jQFSI2RG7IZVWJdppHWW24Nf
RjaLJbs3cuBefmNBhBLZ9zF2TPkJnUggwxhZCaB3Tq4M6JblQaX5JeSMSk7K0m4Y
/zxlY0jAZY2JnxVK0xmuFZbFM20YzRbHw4eKqaQkmz9827PUUQEv2tOC2zOvqAI9
sOrNh5AuLFV90VvD2ucfT/SPCZheZDMJpSX57ZvlAanWu3WI7TaR6I/2WbUWoagT
Jx2e/h+hdr99NF7Qy60vFOxt5/JOVU9C9hseu0SZUBq+wVRQ1AdjUziE0+8oM+nk
qCz+Vr8LCyXsWaRieIonKCyZJLKM3NmcdXAMBD8SP5OAvA0bCzXrewftK+EEdpe1
9vPB3+kjfs/LRV6FZvwua1StJI3+pE2Y6HtMu+e3EmHwyfDIQffq28JEkr+O5MCl
iq8vmDMXCMPwvr/JwiCuaJP4zYxP0VscHNrODxi3uGtevUG4mZY9xE+PW5Fg8r7h
yQU22cT/F4yd8aWd+pZ2yT05/Nhh2T0Yg7S18hufdW+gKeHl6lp/GWkiGs5rdHgN
CRwwVMZhse7OGWetHCxa2pWrGQfDb26hcScY1jbsO9OQUjYMgiLKptvgd3Pso8zp
OXAVtWqcDN1dIauKUMQce1R50j3fBl6/U6nUIla5Fu0SMUKcheZqJjVAfvvhthmX
o3IocFwe62UTKRVXNRXtIfj5bd+Wp5XWNtCHmEl6NmnLWWApsH9uXHOfjTbWahem
GRwC7SxAiojKYTKeK9TySsfTWbjWpxoCxX1jPG95+IU3ol8rFlqtDV5oLKpmv9tw
X9fzY+IOajtttu6eNslTFfB9iFoLxf+CN0k9mII4yHrU4DO8lMWLH14SY7TgfNbx
QAHMYamuqS7TJd1j75uakJJprLbuS1+cWU0ZjFPSrxfPIGBvNM1+WayZjy8dtvIh
FGrkaAiQEaNo/8wKveKstV4ja/92FFcxH9Wvjikn1aGH4dR1TDZaSH/Nt7YMJjp3
+QtYbuywKhhilOeoYfiRvNQv2WPVSLrX+mgWYqAjaFjWJ8LE8MzazYnDfr4uay03
ucY9AQlKiewmTeEyX/SHmIdx5SdKA/8KtdGp9rSwr4EOWFipMSkw3xQOqSgWHU6X
H45Wtt2bEntQptGC7JYQT6EpriJpMuk9peWhWAUqi6PXFYFjjCdTeHMgKoS6t03o
FCBoZXWiGXKjFZ1+RKRhPRAVZo0Q/xX3Gr81ZxMznXPg3alYFE17N1ly5UID7F5o
PSSpiLaN2bPGD1Ez8vBNU3tpJB4G4q3CVI759zhisylMRIXPbEOW7XjBFoaBXB6p
qQocuVbtNVsxiCOTUeZMgzPyT/0WXuUT8WuNXMlu8qNb92W8qXGjRFw1RwW0BioP
TYWhzFNChuzD+sbEopIb8HIfRJoVetrIcqQyxA8lsYrKTOQNRUQkgglhFMz08+4Z
J7z+DkBKzUOGae5BCQ0MH5j8wgKoQtjSW/Sg/rDPIhMj4YkutZIMMY4HkJPOXHrM
uXL5B5hVERZBdzubvkCK0RmahkgVEwVo1W1WSOYMS08M6fF8y29iQn0QWOcmwhg+
G+A76HpApq9XYTvJJeKKVcC6lwUU6WJgRjS8f9+Z2fd3wAv9xPI44qHsSSuMdh/d
NELXIIXpxJY3wuwitbwHWvkueKxjrhEVBoA4i/wgcGL1RNS3Y3bvFXQV5jgX9cYM
iV88SfQEMmzRyMFHqt/i2BJpDPnftJPo0+KHYTZpLpqJueKPQOCxbgqeEIGuweDx
/ksmX7JfjS2HKCpOURnOvn4o0MgiKqKQP93YeuavppWnKadx1zljnfoyCb51j7Nt
Pa/mYa906HPFHwa2zlM2nAghQDBEIdD8nLq/9d2bPDbz1ruJZxIPsp7gkjYbFuKh
30vfSAORrHprhyusO/1WiCOGBIavxqH5JksXSdr2cvzYElVOpAkNUOFuFtzMn4N6
7CUg/vGfeFeUqfpVlRSb8XX5lmZMYx4aDfC8SJLlbeUPLgwW2xImdOI8mM+nkmoS
VoA7ZMPpzy5PpYP/n2YB2E5rLpb6Q/z5D9X/7ZZ/330R2mT8GbwoJfh7xUCxJF7e
XTv9S6mQCpDVPgW8RGfep66SbtPP61GNeuin+4HZPqWX5RE9goo0URoQua0bYB71
mfX+Nki3OXr6eo1Ga1TbWROlo3/yIBIn8CLxG87FUpJ3Q2TGrWzLV2mfzb4oAQnf
9tNjYDTuJRk1QHzvuO80ijYdU7qFXlPG2l8NEfZn2EJfMr5AjhlbOSnflijdFBzl
2ZJLe1K8Tq83aJok+lqfRRrRFHFgVh7s+UCq2ISgji4A2/TfT9BYVCl1+9brPOcU
r/CZ95RT4ff5biVAuXBI/Se+47X53g09xe8nHPh6YkN6fTfuAOMdmFG9BDaIutpz
u3dvMc6ec3htobrbCjCY/xlp39XgdPrlSqQS0uGugIanluu/hBExAOpvEWgFX1Ed
fj1paCoYb4NlnEjq1rRJ4qhyhmNe0b5sS3ywVuBS3MMQu6fizmSlUcNyYVhTaqMO
6UumyjsoJMmweChDtWKN5YQfeZvE3M/z3SeduoydWCtQqIYRyTskrB56m6f8S1c1
zLDSl/ftwIeZg+ADEEHaLOkuahiqUixqG0sIMuQ5I154bFlZHqpyQ8+Ys64ak1qU
5qPKzBF+Q/iBWmijEVfQ3PKXyppxtbem7Qk1IH1GMgb1++GlzPdz309DgXgPX2sv
0BvWNwwisNC1czRjFELCjycppcf9iX2B9aeh6R1Nm8+aaqcCKVpm4oTjDNcDy9Hz
XvE3V2pawiJhl3VTn1K0DSNaPtYql6vmEEccIYkZf9Vs6WYC2eNgLrCo28NwG39O
8RVOm/WFsorPDQ6tUh0I8ZZbG36zX1fKHwFHA6VYGJMGwVhnGRiBzvKt81n9/Bmt
1RuW7t5dftUAxF0dUR8yeCabFdVTEAEmGxnKn7BBZki7n6XVKTa+VBWL24Vz4JHg
dib6ILc3kIsUhQsgewtUVRcov3Nzn1vlUlbLRH+BWUE1/UqHjXsSxZxHp1mG4H9L
Gw0E561Ia+NBwGE6WYQo07pinz771z0pEYabzQPMqbdVp6IAjog7WhPTRKdAFiZ/
kOcsgZPtUwiby1y6mFwhoYelETU11jHKYQcafmPzFEgFlTmlMcipPFnAAGRxwyUE
c+3KH4DFW8QYib5B/4bARv9HGzgy9eimhqDqdefAdHhTLA9DKYPngK6FRLGlUAME
ecxckaKhkaLnHGjaL1OVuF18n/Ma0Z/cDGsOhuYCHnsQGi2dFllth1vS3nCLdkJt
T7E12iGgRGqp24rlWxDroAIJBp/p7XaDngTLhWh59BPN53USQX97hbH8e1trYqK0
+vkpJpVJiKIGi6QDF4xMHSIfg1BnvHnxTBAtinOk56m2xycCsjjpPbGqZ58/xvW3
EWrgTZo6Jk+rOn5YNnoFQbLyKXuw/PjgU8teNNXxDGLtcaHwAoWbDCcj1zkG1zhO
A8meI6gVLQY0/LrT8YMSruGS8novP3ZQ91QT6oL7WeIj7JyZHEQuXqvjdIdrShkM
tn8HoeNhVwKD2P5gMnMtsp//B4GzeUjEcn4F8dBHY3c3v7UJF7Jy/dkEn7LcUFfh
xTMuo84U04WOuMnobMVsbALIE7Udnz+mLj//c3Mpm2C6uQgZmKftKQiWWki+PHe9
HAuHgUPes5ymOuSj7CWLFKKIw5pVegbj1tNDO0b16EyN3Sfh5LAoYUEfsFwtwT4O
7clx+3URaDX61zLsTvdmSosbFYE/k8b3Jy7nDDwINxcByGs5K5Z3ylVBiG6CD+ZH
xgArjmkBbl47e8dkAy475qzua55coSSfJUIOXz28/m252Q0FM9/uruoyLaXmBwqW
/Nujxpyvf0kOYB9C0rGKbYrmXJR8gxlVr5y2mKWV+sN+fP5bknKkf9AmvW76j/bl
zIQx7oxWYHCsnYZC9SaZtLmz/HWFWUdWuajwZLJ+m8Bdwq97XORCBiTMhgNKX7vR
WhZNcgoyv0ZwA7HjN6AeIQLQ6Q4IyL8Co7sNipjjRhVJZyKeDJduLB7nqU57GM/S
G3bh1GtvU758CNahj9qbPfJ/8iFzGJoSeHuSNMn6cOw9Vmj2hrGwUxDBYN298w66
eBCA5umfET2Ojvo+EdC5jezT5RUTzTlTPjmOE2DhdnRXUeHXzEszjaz/ppa1FMgS
tZEb45feWel9fiaI5PEMOeWbkg2az34yQHDaZNY2dVdu5Xx9KPmZZaV6KxPbuhdC
1oXzjE2mK28Q0C6QTUXi347S5tF1bFm5zGdlgk4TrIUEPnKT6I2fuZSZb0V3E+6n
FNUzMOE6Pehd9eKLGYseqfqQRFmvN1l6A2RNukrUWDuwS8KmvXQQ4wUqQ9ve5exR
hR1mK2Tjmh7Vt6tdT77WbUqnPs61KpGnOW149BAoRqXdlDt/ObiaI7+6FwN9Jmt2
67GhxOfo3/hjBK6okgj0g2d4x2YmXXZbj+Fx4eqGbgqCahfHVdDHVOQSAZcAjefd
U1p0467/wXIknvVMPcBOvTrlBxbV8qdPXCvS/M98++R9jyfNEijdgcPP+4Tvbe9u
wb9ajRZjKJ7T7mx1XV7nTEM5020eyibS25g+tBUtH5VUlW9KiOo+EZqnU+JuE1o1
rbI1j4RhTPmVUIOd23b15BqFf6SKTzDBT+eVwLQAsfnh2TrtbzRU0z2Ns6dLiEx8
diuHAGfoH37cMH4tVjGhNDVzjVNGI24KkxRSaa7RbDo/++KTosCUtdo3cJCJB9eu
8swuiLyh5Hw3uSdXPzc3Q885wZDUU+EYclkqFc0sRCCYuB/kpWzuDtdeGr62izix
Ga6nQhJXD1oDO+xHkIBqtUKkANH9+gTLYmy+BxUzqWpDUuNj8YnB5TqhSTEzZU27
LDsGhcQLHe8e95wunJSFXKbzvPgTMHm5Ca4PTfJqnNjteMKLIfGgXmAjrIgpG2so
SfdfZjlT2hfs32IB1wL/x61mK7QQgTawdwmTve/FfydG+00pHP8PADEptYr4Oa9q
eE6zbElVP6BoKYBhsEVUCjBsQRULJxjVv8CC26F2MR7AfdC6J/5SCi5jNj8TmNBH
ML5mgZ+Plsga1f8ARr6hOaa1Yx4L+f5D4R4I9jHu0lrGcshsdWcd9jpyAH0HPgKh
5i529iHDn26I1JzqUKGGZb471nPq0Wb15+VQQauM1yKIKkA4jGIFGwaV5HxFamPW
rqMTZXBgfyr6lPG/4lyPPHf1rrEPcjAvOq+vUT9ojBConVOrqqREINzhu9L9+JoG
1SyWGmnZ+hGXNNlsmqGK5ihLqublRplv/bvHkCtm4HMny8ltsfy1YErMjU6SBQTx
YQpoXif7EfjP5ein6lATbKmdMjT1jw2ojPuniTO+EmvqxC+3r8ZZzjW/1rYz98IK
BXcLelT8+1no5jyhSBDkxiWTbX6sVm6WV+5ircYZFDObHHTia85QskIF3vwO47tN
8UblIq4tmNyRjKCpBwjBosznrYu6cogqfljf4h+QSfGrYbU0eqb2WSYD8Wg3LrUW
b2REzb+WeKeh7YkzPFOLJZRf2YUlenRquFskMfSY0Nfx4vFJqDkf8VEPRoFoHURp
AR2TdqsTvvUvOzTzKoXJEJG4yHp7jbypT4UxbmeSlqagZHfn8FjIkKxszQzYL8JW
MskENUqobs4iu73Yr5FiAR2kdJ3l420tQbIj5FkWf9rtTkMhGv/tBv/6cZs8m517
lx2KkGfiSTzjDcjjEMffrc/bb8SWfLkU3kGX3iAQaRpZa/EDOirE0/q6zEnyhlFO
NKiEQfvGvdXzZ/yXQoh48DKBj6+zchstAlB2xHQ4v9uT81XzLvXMPRmxmZ+zeoqG
eZ5020ZZZc9bwNGalz6rkjY0ioWNNTgT3eEVvRs/zeu9TeptqKPO+QNnq1wkzl/X
fvvKrUBzqwB4Cx659UXSX1W3MCj6kNLivMi3QJHdB07WopyMhD0G6+DgwzuyvT7E
RiaV8QwcCgMTwFtXRBktK1ZJcHBpmYY+g82V2EOd2J8hdJdhqpLg/s3bjX/+34U6
motKdCqMFPA6XIDuoy8Aw6D2wbM1dOW1Amak4kNtFWwo6hJ3hZ1qljbcpNjms6qo
DSkluc7hJ/4lb5Nr9uJk18S0DOD17SLRHtP7nIP9X3nFDMhWDKqoS0JAf1YQiL83
n9+VKE+PXWPOyHvZsBC6xo9qWGrK7suzzRgE96KHMMdC7KnaplrKKilPm6B6HZDa
VJPkfAV5AyPeDSegr+30iaEoV/UUOUrvC1W3pFzWHUJlawDbalRCy7wIe/Z6svyK
eznWBKbslN50itWY9A4UN1Vf+zO1hskDmD4s2aoLJXdpZhjDh2eAAghieQWS8WGc
n98cz48Tt9qTtlrXiLXwLQRW01BKiZIl8VAazoqASNEwJBvy5nLPy5C9BxB3x3nc
LL21ycHtnSCOmnhZ8RCgck1Od/bAKqjEONjntEhkQiyNFlP30yw7RchJQccmvBY0
G6Hd7LkV0SoBCVsu1EVWLt+2Y/BHlsfo29cVPCbSJuSgOtK+yJ06BTYa27Vonfk1
X2SdPUNwtwGmDAJaFOTow2xVjm8N0I06DzIqup7aQF+tiUiDWmZxTSWFhmkkMvTd
AuuF6aR7gx73pb/JeYyU4i3CASHmcgMC/CL1tFuJjDLhZGYJgn8Dc7XxnZrDbqc4
wqx9kW/QV4bpALIKcANDKU1r43LtnTeBjv/6R1WskJIdssiddBaxpI/98hP168AW
v2j6UgcXw/p6P+arjo1o4LinJFxs7QE2I4fdJ/4DN4ojUt6JdQCFIotCNCj+dJu/
ZMuDV37yiM+0mIdax8/wfp5qvDnDS/MuKHwMx+GGvKXUSNuaCm/uZ2W55uTrYdjU
P2hyInA+pbzh8GSEnHWcgPanLX/ClM/YeaKHm+scyNajpzjGr+RUSHppxE+5laMG
UQUMg/fuEwwJnL9etyDGEKzOcSCj6z0Qvfh74fJ74hEgWbgn6GF9xZTrB7j3ozMX
uB5BgAmjXi2RyuXGQZDOCIATr7nY107/Aeh3Wt4summETdHxo9lmdPNPUDhGtkYm
HV6jgGVnY5AXkXBi/sHd+WCkF38AcFwVqL8tvBWgIoMgTgOdBBRrVAxbVnuQgPQq
D1wzWLbPdsQ1+/3iqV1/aOanJnzDrCkRoo1VC8EkMdvSIyhRiZ5wchsHxYnjREjD
rSbMAC0Uo2mMimVlmGAI8diWq0CKSwZp1o3Afpj3AgpI3syJ8yOMbegDwGtYswfe
KO8MHwV0w59f8wqTRUZ6zLBkfZBJl1P47OxmqLJ01e4vnrFJhA3HkvcIgJzZlQtH
c5GMRs8Q9Bc9VWYlRlTQ6Nxh1uUUd2vfyIXeL/hS2MFSxFpcfz2oa1iK1KNhlt7k
GF4mBC+sCELyT4abyyBpPe1wVIq5GsBoL/xQSlC1rukH0XbjSE9L/6KbmSyaOYI7
Rpn+bGW/iXgAHUN5ku9UVOJ0iH6HOLffroqMWTOaHdsN5ajCmoImU7lkzdtSQCZt
o/D9KKvjQGI4LlFrAOEv8eJNEo+LRyiH219fN2RckV31Vtm+pc1jvZAX8XleM14Q
1PMYrxJ2fgPf4G45CLe/UJe8YwjYPtF1gK/+xAS3A9MJd/ke3EA33UFLTgDaVMfG
uARUqrVimlaMu9mnYCS0hy2TTheyUcqJNaJcbVGGI46VGMjZghTejdmIhy2A8vVK
L8+Gl1P0emn5om8BbCWZXUH4RUzWV7TK3qUOrLggHW0EvzU/F09zqULQOUW5NXO5
YR7lM9eH1BNz3uWpEaRHVBxIxWC4RMzflHL0/pLuSdDWjYrD/yDDmxnIiFYNK0jz
LL9XW5Gg+8eQWGq6M1Vno9CXXjOK57S850fEEhNAf3gljJ2Krcc/ZuK11iFA+Rfe
Gr+YaRLCWwcD4dKJfchSxdiWmUHRQjwJONvwfi1SxvEPOeJPd3ISu13dStveFpxr
mErAZEbTM3tPn5sHhaJqJrYI/QhISuxUfcdfl9TBmmPoLC1SY4nIwyh7RHlOt6CN
XMKnmzCwQZP91fsEgrahocTFPk0Olhn6whNc5MMcdHxdzOByVDohDGG/yowtFkm2
tiWaAp+1YNuz9z3dnQ91MfaXUt0rnulAXN1c9Fqw+/6KbnSt4Vt5NIKwmBE6GlbV
Zlxw3j2CnU0+XDmsh+xw259OzCoTAkMLgl0oSqPzZ8JwvQR/gCUF8GEw3//nIT20
I3NYqnosI0khmdQICbSrPooe9Ao8FG2q8noCWT5DHedMdV4AcVqIA5nrReOUtp0H
T70kIEf1OFOjHkLRTuIdcwP8Msuqb0kfLeaH0HOa5+2h7gLwYuS8ghBxmOx45A8q
fh/MvCJwFIBGQVS73u1Ath8N2V4Z5vFwVWx1Vd2EnMH/ITygCtij3+yeaKtZUidZ
2Q/M6XcuXinerHzmTYRRghx0qzOlspp3pPf/hwbVOnhDBBU9ATyx06OAs5NonkDp
FXwT5s0v9NYyNcARofyC9YVe0lqcnG/iiJ7lvnWCSaNl/H0D9IjLKgZ3KbUzromv
/bAetmEylD0Bytpy+gW2bITTH8Ar5TEX1x8WXFCV741M3HNKk3ncYtxrQ4eQ9v7q
zhePwmzKLgClky3282Ws8KWfylnSHUX47QhJrQ6hD6Tr+Oz3OXaTDX+J3jA2dPUa
K9e0DLqYxPVkvnuX+m/CDfn2JWd4E+3cryC3OtEMnlQHsjHb0JjfFETmoR0BPonF
yjGgA0s6gk36Mw0leIc5Q19n765e/1uZqtvwToTCUWXDFSoYeXlN7hBn7mn4AVQj
NJ1691g5++UaE+g4uI9GY6tcGAaAp1HA5a0gBS1Aa6o4aeBBcxkpksBfuenUMi3B
8PiSfmS64ewokgEEaIm5NFZKwGq/QS8gCH35CpAR7hSqSNh7G0nyQ1F0Q5qJDH7b
Hos9kow+jHs5KZVPnZM18Lm05QLpMGhDBLV/4NrKt/hOsROr95TlzEMKcHw8T+p3
0UxNVrMzRO6hUdQ/QkGqTH5NFxpOYtgQJenbjui4ceN6OVwn4aL0ruIHlOniLyFY
nadIObcSwYYt5Qr6+RoYCOareHSQ1yANZ0hq4NAKK9WMaN4FsgcWXv8SBQ3F8FxN
mjOzZFeAIhKyyTHZcm8JM+1lkUkBHPyjPbjRSt5ZtFK00j8EhoV0qrLgX7e3OcZ6
g3uRrZX6kN09KsW4TFLTCTFBgWSONRJdHfTg/Tc69sXOYf4dj7ORR4lDPoYQlstO
HWwtpJXq55zt9gUB2uZaohvyrNyB0rCGoZhB+3QtjLeBaJT4ULOA7AjvbFHkD1Lt
J+yoGvfiy0U9g4KSadRoVv+F2hpHc4opUZjP3AC0Y+c4QrmsY59CzTOWyS9VwUdK
Lu4TxNuYpa8i+hOYqyqHQeTbNYoj9zeCWnX8xA/SwiwC8YUCXx1QRsRZjAwK3T7d
EZ82QgDQ4As+PYMyGTr1b3Dbx7jAhJ5xVjd+9Ad9nDHDaCRokyhIeZvUBR2kSNLL
dZlY1JFxdGEglReZdamW6WjADPETGIKTQlhoakFmPkDCQp8Vch+kzPtbBMPGSGEE
0CEQT+CD0zIIQpP0D0vmmiK69JA17sDBPNwOTl3Rd/YZ86v/9ubvHX03bjRSyZG0
gEy8yrEdBK9xlC1r2zQ+q19f4JsgXLQxWEDaddfZwkr3hhy2pGVZhog85FNtrs3R
U/NWRFDdBmrM3lXVuc8BvX10nSgX2TozXTtib+2T8ZIuIkWd58Ya7yhSebRlrd8/
CFuwyJCtLT2VuJCwmbvQD4iRIrqqvK/eHXbUbMghc5NqidVxngJXHs8rLpyDj1Nd
10yJecRd6t/TjXm2Tfed/3vY3JFhIpzGMUzxzn3Rxzp87Z8Suq0u4frpiXc2prDE
Jv/GEJU1EDhUkI3QD8ozmyRvaUHMuTL9ip2DYzfqH2W3ts3PELN/fQ0aJvH8sAyj
vJkhAQtTrVskYcUaJtIQMM7GHZ92TwUchbWNguUC8Inya6yY0AjGxGndOmS/q3Di
DJaNFoFqWhXdBYaNhCz9XASj6cmn0XB/XYbb1oCoZHNLmHHyjOMOZzVbKiwdAu25
Rj0nNVzX8p89E8nbUYRF4goUJfNNL3bIZBJeqz2H2zPLGe+hHiPRJ9AO/5mtYYQW
CujuYI7NUE5jHCxb8PeSaxTDt2310876OYshGXhsE9hoqR8rvmDIKUrbA0VtJogE
vFOfhx4sPBF3JBWnj9Gc8RrJxVHJZd0Qbss1n5LaXeDPCwM0zJr/zCWHiHWOpGkm
D/VHSafpfC0kZnitI2IlZyqDZyxtVP6NMUQ1dAu6w6PfHRx01Kt+p85KGtjsOKMw
uZyO9L69CyEvMRBAZ4DQj++Bp8sI7bKxs7jQkdatYcm5Axb2hU8txJ6mvR5dK5SU
fFGCz5ucwzYytmveyHt91al5YxGW0kqWJnQulYBM9qmza6cDQtyf+Rc5/Ct0tPJL
S8ZewH1QaqxYHwJ3DgeoPkTjIedVBS7tJHmEyNeruB6xhQ2VWbLgUPT2mHWD67h8
wokKKthVE5cIRgdKhSne2Npf7kZcU2pGcxhj2s7V4+NUVeQqXD31W/qp3TzyYKgw
hP1fKN71ouQRZrpkVXPpCC1iirLv72rMCLUnVnZXezByuRSvUD1ne96K/VTBSdBI
4OFyu2Ke/lFKordMUOljDyw94uqp2/iNbYO/QfbuQymHE0SyOdPHKVN+VAL7vXk7
9Ok3O7ddbVgKXgMXOzJVL/0/i3AelPCGySgE1bBvguSWY75u1rnK7C9FyZW6mCYc
/5osbzmzcO7ZxOommx+wX5mlsJ/C8aP3t95Hpwg/5rmzk3S6GhxYGB078kHi/5Xi
lNuupAX+YhhUF2k4//AFb4kofbSOclxiVGuVn0a7hQyoS227/iM0oQrWA2QeFork
a9HUBTKGyHA/J48iz93vCRLdijWdgob7p5n3Qd0rWD5ob+rj78rywdkDsxgfqIVg
ATa61IaIgyDVfdcZp0/4WlQhmwcq/j3J19nEIexZPXpKY/hZbJcWp6qMRyriI836
BBAJGA5EJzgnAGYfgmFAmIi6eEnlKHu/c9/9cADqu5WsNezV37goRTdS82y5DVR7
iVlIc8XxWS4bKYYF3bJw1NPek8PS1HoF8HY6fMI6nNA27lj9dCxTXapzsoqZj8HR
Y2PhEDnbuJukIzpwpAY8A51cMzZpBQ/mMkh/hDXCuIjATKn3BwGOm3MA8BaCDJab
ZBHUHnKBPvT6+7WPXjfRY+OSDtCkY5VNYbYI3SomMrw8gvq4n0z3p6Wmb+nswtTF
cTivY7EpB4vY7be+ElnxF/m4UXDxS7DQnU7FD3oFct/+DXlxiyIZPmqz3BX2g7MP
fOAPsfBKBp1oSR3pHJSHnewLzR8suyV4QbPl8I3i5O9t8imn4UoNOGlD+XO3SLKO
4aNDaOVnNuuyQuox/V1brxjRy1O7fCMCFHvT7t36Hv0aZkwmK5I0FtQzj9LcP/c/
QgcJ9Wyy2On4DQu472VfZD6y7S2G44wQen8wa+GSii0SKYlVKD94QUj60edyyyFq
6vGRe0krUW9cgukEtTcRCW1uT1KpGeplgGnIjxwVARdo3bRsu4xbuAeHSjbIcMmO
EgKjLfmh1mUpHz6Dv8bwl+E07qecmM+JBZ+2ZczOq45RCiCM6tpcTWT9ovJedUvD
nIe9tXis5YMYPc3nbF/4Aa/uF4Cgwk3KKCHzSWUbOEvJNerJDqloWX3cKOVgjkmG
JAtt0OHvkvMv41Rp5J2XsZ3wFMvyr1fgzR9ylPl3FP+9m5dOakc6Fe6M/a5+yZjR
pdbCnEiDiYdANBEPa1YmGOVLXD0hrRK6cmR1wRr3yrSalO6WOQa0XuJn6IHJUgrx
1P9aKliDecJhLxb2zi4PMPuvVG1/kwXnffWmT4NqEioY+jmijXQJhQe51iph3Pv6
xe+MwEeq42YoK8XYDsMqmHOfNsIhUQwfubicUkw2Nrn2eo8anPUiFx5ruIqenDhF
TEE9SJDuc3Yn//D+GK56+siMmnlcJRVAe9hqzyQYY2PDCJUx+XKq/XSue7WYUCKP
Oei1YgEQ6xKBuJTkfERtFC8aQpcqfLTDu2OHgeqqVUe4yej4CDvDVFXqSU/mOhSs
MKXKx7AzK2Gs1HWFuF8zR6DckqF1BtSTUmckjPDvys1+HoPb3zUffkIc2Hsy5GmI
OwJAP5gmPsLouFMxtJqKPvNMUlQki56Rg4XdIkvEAb4A0C+JEOTiN2LIk8N6e7wb
iyo2pMGLs5miFuaGPwliANzhjAAZQEdncq5kOXTYb1bpMsj05R5PnURzgKdAvxiv
v7WJcQkD8DalGbl+/xTfoq//66QSUltCqSlqtXKQyilCPMldeDVxbBYEMTzxA6kP
5ZTBfewsH21hKzNJOhqH8E1p4fwMclEXgwLOf6Vd8L1pNkzt9GPYR8tMveMCGqXq
Nj9L32XqBgETfOiwFe4WdZYu/bAqlMaeCd8HiTk+54PgUxS0jpIsWJ0tbLNs369x
4QPGA59wTUXBTqgjdD3QVEG1kRAo4QuVF+m9pCGtKKx0Ni48JKVidSgdIWZUKtfF
lfulEnUwj/22AO2YqyQ+Pe70sMDa68ZLTqlhNLD8ifQvV6j382nbQXImUuA/2xsC
CQ94SgSKJpEuVrGTu8n17ZonhOq/FHfH2MZdjzm/6LEzRgEdfLvziP/THGjJ01g7
ahXrJFWM/574Qi1etLhhJYufv7E7b99DC2TGJ1VdyKVSFsyg1ZS4tVcMz7mIK+wM
cxXr6Y2S2Xr3uzbj1YZZD92YNVhOqE6EsObxy7JxdClwBWl03LQHDa/aKXLEw1kB
+vvMCm0X+cDPOSgKuMwtIJzOFS+9VZbY7o75ztl1kqqdikq1zNUXyw6nteoc5YvA
CIr9e5M+wvxZEFuAsHmEc5gwRZMeDCYbt3/0SI3nsBOmXHLISBfrGPx1XniEwdHu
oFS9ePcJ8Zznf4G2sr5Z/N5ajVEMamkTtoDVIXMS6j9etlnr/26avTQ7uyFVaRIp
AXhVieDmwEt4QQagQK98K3w+OPTPBFbxaTXUdY4nXwh4hsA1cxb9jBJRfl7RO4nC
9xnON0husBvn6tuDSpXU7Z+eSJxJUsEuP3rb67M5tIQa87NvW7QZCBHxW6Qijozp
vXigRTkKms36tTPq2MPnWO4JPeosPcF+pPt8XZ02gl+64xFJ+F72NV1sVBEwA+vE
zUXUwS1iwjFxc9Er3aACVzWY6cUP2lapOID5agZ97p89WY+ssENZyvNtZg43ppR2
kl9lPyZdBUgjDk/mOX6NVlbhfBnBAiBcweRqaisZQUOTCRDuJfrmEkhCo4bkVL1D
3Velyn0V0BZ2U8V07UlbOmfGnIBhCNaBt3C1mNcsNaqPztLxslnQqkzj1FlZn6dL
4GKSFz6JopC4Kf4Nv+RUQRubANuP2YfIFhAiWXUYUcLoiOtsPVQB7YtY9OYet9I7
zjpzzllGXF+gl5k65obcB5V1DeJXq3DmFKlmrlkZfsOIs/zVIyB2iBeb0H5lHxs8
6mUWBXvH6hbif6XxVQcgsOGiySB5EppWyDqYn1IlDo2Xs5bsHlBlVvYAlf97MLsL
j72uIXcGEr6HipWsfiGPbke4nsQuBkyOLg//moro0En16Gsnl6KEmV/RhD1lV/Y9
8KvinXzB6gEnPrttgyJ6RpChqjZFh92NxooiRAdcuxZY2iC6hpnN9aaJ4cWBxbom
b9YwqIqhfMP38Knp5F/vSInDz4NTHK/RH45+IYM9EsJK2dALv9cFj4/H4pz3LsFa
2ciFRF78ndkjtkxwffW3aYwDtdymPiK4OzGb0qJX/4MI8HRVJREF53uR6QgE0FUl
vk/TYpH3tF+Sugjx/2IBq8z/x261hGrxaN906Yj/iPXRtcN7vQE4vkOWjVE5VKOt
GncBJ5y++TSB5YcM0zVW0EZWL7ZodPAUEigpzvraLrFlGoADqfEJVZ7/9cPLfDmy
rqxTLqnNqRysFGPLb9ON1XW+tQh0o6CnJQSI7rKQaOhG5mLcnFRduyMZPRcyCYEF
/cHQuquVTOsbH6NHNpQsEJ7J1zXwuZUAgV2GJv2cEqnVh7rJCWOTlkl7zqDAN+It
N10FPU9updRtGN84MR8aur5ojXlWL8vAoIUiY+o7Zmw4jhWZNTT+JOS0jToWmfb+
s5bOKdDROX7XxzwpxtD5anGUU/0GpAgMVnYokVbvQTGh+3kseHn9T7VpXgCyVjp2
6vSFJKwl07U/pZ52en/cV4MapYvU4pS/9Rdef7ZUd+tsHAxnBEFovVnHIrCcCMoC
Ozfw+j7j1kUvikL3CYM1J/Ejl59V2O5eKs5HEZg6X0lLQPO55jdlEODOkLjztGn9
Ux6QlZOrLlm8ie7XTnqMt4qZfpd0tHLujr0nFmb1sNdgH42aDYAVgZAibEBhTdDg
sXff9BOwn1IU/GUVcYZkweaeWyZ6BEDJ1tXqs8tP/Gp2ALSDHAH8FOTtkX5VO/W8
88FWIRDmcUORBZE/+pU7ulctWAAjDjdu3xF//wxYvrscnKHSz4KvdZ+ChyiEP+88
L2XOFbQBJVEBZZPuuyQdS+aMw8hQvU+gDHD2bIy2EmfSozDohW7VEC02X0SRCH7D
IY10dNe4mA2NbM2bnxWjv7RqQhniJODHFIYG5cNdrfZZSFKxqI9hzmzEpdvHyg1B
FEnCz+ZAgCNhxaCviGMFZ9W+Crh6FYuhvyIJv8TbzXjbM67gX7n1blVHj1uZ/YIC
zsoZ/xrnHyT6NGFNmqr9qExE//r5NS294pMxJZY229ugMcCt5lINyC9SsDzhwKf+
yatil4yLlQzAfeE8Icxh05Rs+wrAIODJbWYfHTXff2FQIVwejMWxndHplTR7dsrE
mjQ5/PwPu0YtrzRsIMy2ICTZDEMXQEZk8N8rVLuVQaJubi/mlBBNtD30zxLmS1xI
yhRwnX7JllxHlTEgAVK40fnnU8h+Tcq+X9cacpf9Mo5imesBQFPUzAIc3JoRdAgO
XwKB25GCfzUQEfi5M+GN1wqO/8z8dnmAHNlCmxjtLI/byHzNlpzVY6gYPSr12kqn
EwSKIOmA2aKLXRufexApSdHnG3RtuMMod5KMgOlrmc+vnxDo+hOJ3ekGCjhE6/4I
dlkNRWIOtozJXGzthmym3dHYIugw9aLjGk0ghXh+FiOYyQMjGB6px8mjEy3MBVGJ
q3iMWYTgeU4Y80TWrS9q92GsO+Dxptugw9X8/5mRf+kNNQydI7XxK6o6yZ86Fv7z
PzXMIefPFByhiPDMk5X9DL4oCJeKSPUfEk7i+z/MH+itJdJjpvfRidJfJ5zKG3g3
j40uxjgteBsj4SEBfXNdyuqH1MhiZd0PRnOqjhuQtwaA2DB1vnhAiYJtaStxJO9F
hhXAn3dX1lBn6qAIv5x1H8hnPhXj5IJek7Wxpb8TAKqISn4FEjQhXDvrui66GCQf
+1VoFQ9AdG3yGACoOxquX4oVbOvwOlCb2sFidwojNmy8fDpXnxj+b+3zB57Vaz3B
u7tgPn2rw4LTcQ/cWazQfsHr06fubPbWZonnP2fZGu2/Ciun7Sy1dGVm13iO64ft
E7H2tY8B6/oqwC42AYj5X0Uqu6KJ6DPc4/TX8UpcCFhQX/F1D9uzgckYxwN7PVJB
rnZ39bOkPDHUtyna2DYpoickTXeOiFsa4CqCLVQN0cN8sRuCqGWTYUMWkQCEi/Xz
H33eus56ZoJ6nfYNVjtS4BTjdx2Xd2YIoTIN3+8qAhqhJ7smxcGRUUXFxPsZ2gRD
LdbLh0dVuYRPhdsppdEGcgDsp6ZBl7u3B8pbkl+6J442JMDr7zPg4lKyhGaAs4Tu
XxcqxKgqhhT2DnjzANJKdKoDgWvik8PyEOtRGWg/qJ8yaPqMi8bSgF6eASFTV3Ga
UJzXuRJ0eUFzzhKhJaSRwCQ7scsCcbMRAQn/IL5ziyOc2pwkzMyvTNTr2a1XlFMO
YI3ajUaBOW9Vh3ZRpsK72Ch79fTah4e/iodFICCWUIdZQa66KJ6C9Y8Gaixt0WnS
JP2BDRGy2LMi+As2yc2Xz/AKlibU41eawz73eQKnKh0/L0p1ext9wdOAc28ve8ue
R/yZO22gUbcqqJXCuMtzprDQco0xWqKiLZ6Umz0U4OOYtkIEa3QjNa7PrHvNWEBa
Cfm9GjzhRiAHDHn0DvHJ35W+aYtu3uguI2rWuOVz9UmaZrC/obgaQYiIB2T0zEwA
Y1E7wdpiiP4Q02Eob6imQ0FwBFhBsr0Gxe+DHBwG2AWcAo07WmjyO7AVRL/MrEsY
LtXiUblYW/d/u5U1Dl2yFIdXgG5Pdu/P+0PmJLJCND4eUkrgxhs432FhqV2PEl2j
HufhXP+jj8tEKe1EjQ7NTRXYspX7XkxRYgSbSY9aC7f49Tm64FWHc+ipkhDbksGz
0N5Ye2bBfmqAhNS2XiBKSD22KCzmZM1p/aw53xz1mkUBgKWaBvUjrQkm2njAOeYL
tQ7muN4grYM9ZFgHHsciTkJWsihVR7Aw9MPcdyEuRqpeyGxDImhI7OUrLC93gyfK
eoofWvCarPIr54P6pAwmDan6WvVJ4Cdy2F6WhPnW7ddB4S3e3MzSreMsIsane3IH
mk54s/th01pu3VODRfY3mxvFlvzSzP62QWHbj4nUWWJulobrZh4qNYgBhpfVzg++
tkWvjVNjOtFqusOzLlldSw+r0/lyE6EYEY+bH1iKUFInrzoPk/VvIhzeMXHG67TM
5HP4q7Rl7DNNSzCn9uKDSHv+zNekINcoxyNgHsJ/5L5P9UfQHLu0Np6KdTv5xa91
Di7jWD503VmHtwJs6dYYQYErLwU6NXEsVGa2stP6KmS/p/Lme+L2+MDYCy2SQPZm
47dJDWUIiR0W497cGBMlZzzSZzEcWPDC4fLkWWWxBB1Guzu6PYdgjEvBymCn85sj
/7iqtfoPXxVHyiAUFRqR63WNcAUsA+Pj/BS/31meIDNVL9i1yXtXAGWsamPoEB1o
0oRdO3kNWBHGbTKaV24GkqaCkCVMtDrY60IhHln0F4VcEAlUfyVvLVpwlKk8Qr6q
I4wxonJTEO/ZFV7F7LoBPc7/tZ01bL+GXhpcZmeu1FDT/p+OndYuNlnMlb8k37mv
DR7bSnanIpAGb69Rhs8b457P+wDlTo82EdMOsq3xSgd9rQ5r3kP1+zPKWICgpVV7
Iuxj//3OLPy/VsqM6VO+DTT0bs2bLOoGRovJ9minWBUTPUZG1DI7IpbmzBFDt8M7
FkWuEzRCNpuuZkD7bNCkCFsD4SbUU7n8gJnohRJoVRDP4JpJvsF1fdVSZZq3jBNE
hELDx8LYUlxvdbxkcRbL08DRTSdI7+Qvr1zHrt8zFcgRPAKZM89BZws2wwIkWE/n
AOnT0UNR5RA7evbT7WxHv4kf+vvgGWkbctkXaNRJns3L4QIQ1SZ0ALEwutNKqDLg
KgIGMdrRV3E8vjta9TAeA8wJzt84uQxJk9FATdnLt+pwL56vCj9+cIxrpfoP6c8i
jfSKbTBsJizc4kGe2PK01LNLeI6v2ElNiSKxdaRWsMMWitcWdmeR/GDeyzWQlGEb
6Rs1J1dBRohyuTBgmZzAaWSFXcTxhQCuegTS1b7nhHA6dod9LgyatyzuXl0gN5T4
hAKKenjauSo7QX27t47rzUQxg5+D9Tz4asW/7TLtc5sPnhBX/NgRujQXqOLPxgbP
NZnLm/QAnpKg6GiZzSINqa39GEXW76NQpQhmuuuwKBEZ7HtZ74DdwKtd94uqC3Pt
WXh3die6blgRr8A4hDDSXIBLmXGZW2+PcxIkMLL0p9RZHH4xVbI3NmssRANQ98u1
n1eue5fEUx5uAoy2sThbz0M3icCiNWjWXpXXQTw/xBLtBScUYbknnd/jC0ARVGSv
CD5rkH8IDXPmsDnYppFRiCLw/TbO8CJynYYMBtzLe+BcPxnOny5MIxGd65SevgeN
qaGBq1HHdTA1cpbNK25uN0O81ZGZiPHQWG0qwH3vs1oXq//KaVQ1153VZyUOiHpx
0mHw44dg8A2MYBeIHnJiosIVnVCHwN+oJL313wwI1vmf2iPl31ZPsdy0KSvuuwUO
xGcqyeZTqnxKbLpTI4Mg8YeZyMsHQhncGIlnVltcJ3RokrO81QwQNt1WrPBtBkmM
LzXoVf3e0CCHzjKeV7IAZoXaJB25zeT4zAK8GAn02cXnMcm8dIdIJ41hiSok0tEP
rduOVp2j7fWeExeGdtd36c1VBJbE0kRCWqC+RmMrTeF4S0/MSE+dxxvtPGX1JDNT
rrmXflVx9rsFQuC244dWvHl+A2pVIiNlCFQtkqMDRBGAmgpMFyKF5hS0YkbjxEXw
B4wh6e1KtXrDoCvUKr0PJapYM/PzFs5Q/Eyi2owjii+KxgYCjwJmXRQC1+vMpUGJ
NJnxPzj2HwDM95JjKDrskDfkcDX0AdmT9ED853MwGCS82F4wRmDjnRARGP3xmoq6
gqEDxb3OyIycn+AqgZDAUbN3FEwSKuVKKPvBeFsKbqZq7XU4NFCpS8hB4X5yGjgr
yAj1s0/eROlASPmcEzcgrmE/Rn/bBwW0Uv6n3fIO6ZugsPImFAS1MZhDnGNfSB6H
dHgmPJU9ZR6sjjL/IIdKjQT5A58iLxwCbnNGzi5ppqi/YV8PtqlTuLlBMpw/vJDe
+1wDMqK6nPUa/gcc8jqGwvWU7RCkfKJVFDv42055BGv2H9rfqksTOG1P3KB+jkPX
jFgwsdhfSruqsmRkCkyKmRoa3/j6oYAReQhhBHaJCIIHo9gP/KIxHF0HNXSEBPEN
pzaqpmw0g8pRDHYCnv0yF1MBbF3qEz9R+HXo2T1zI2xR9g/rXPODcqwMXwbCCvws
M6oNb0QJnYCj0wXtSaYUDZOQ3xKPK7tVd7kpC5ukqcZ7QGH1IJC+/hyX2V3ciJRJ
UOptkjjo5E3HFYHzzPmrrmr7klIwcZHnHloW7GTegD8qb9nNb3BeNdI4aWr4n/Nw
ntkko4BjKAYX+LymJ6Fcv1SLMqPJSMaagGKZNw1kIh1Eez2gge24qxyqapvFHmmG
tsRKjD6W4prs+eXjwzKgYKBTU0833xRb5xaN9N8tCieULvobVD2zJ9U5HBisO+x9
VdgrzVNdgnATiM3Sh8jcgJWxISMyBUUp2QqjMPq9H2A0ZIxOTGQ0AWHq9KiHZh4B
5O2djVmRQr2eW7VJUcY3Sbx8pYqQe4yxSfMCwe8zbuy90o9XWVKp1pOvs0BxxDqI
tLDDvVU1tgofbJ53rm5uYbWcgoiBn5z2YKVnxkuC19Q8O1pNvPE3xee9Wxah5XEf
An0MD/aLluLp6u6DCbmB9uQZ9nxdlgNix6m/D4OwbWqx89nYOlKWn7tKHpEKL49f
lAe792Lh8vrZErKdW2fzMGSmnvva4+vRCemqwbr36W7m78J82mvnnPscwv16IzKG
NSBRqULPb5MUQQvw/deM8dpqj5ElpjR19vX5ShjCAZ7nw1udEUhSB07/yjqLJ6Ax
bYvHnQHBngU7RSVsuZxL/7xG63qOGD4u2xs5V8RxfHIfCVYbj5sYzzdNVN9b6l6f
DrOp58kOo0PRCn3Qr4Y+Mxf+54z9NDyFyOPZsCMan1T9Rsi/syQSwqy7REfpnYdW
gxkVEVYYAKx5u8UeP/xVwRW4Te01Ow6YV18X6eSS8mSLGcazlBmnoXndedk0aD8M
ouVfJhEpTdu9cjyv7xlxJiFqgqodoXtRxDJCNPfD5y08gmxSp70T755EemqJMP/o
/U4I5jWS1/virNDbXXFvVhJUKXRpCOOMESYQkwj7tpn5XRAOEFnAxnazAvIdAg2/
NcOZazL5Jm5pM527mymSJ5yGnMGEb2CuygFjsuPpRQhW8MvaGwabCwvvRLeVCBBb
umGCLRmsXHeTWqkRt703Kmj24sIuHqS/ozjeIPB5f9N2Hec/5W5fSq13dT9wYesL
3Vz5FCLvOMoO0TmoAa/D+49k1i0YKTKTtZn9h7TFQ9rIpagngBTMo7ZEra63w1db
qEXozY4OSBV1wMST+TcxFLC35GW3Uk8VEQhnErn6c5+W80skcu8UO+0i/g4m5Pjp
pNwkbBzsZ3e7Ii31pdiFSZttGVO8MfPdDX/9DypIEji0AigJfjJvRtVFVd0OGSdU
XwaYrfhlFVFIaszbCPLCJ8jlvGRaqEvfKkXjLBdcK4xiV/ALh5Cp/qIbDydxzeuJ
+IkKYunLbxa+9Ir/aMJKiGdFnNeMsIYdLALbTWy2WYQ9/jinSNlapJm0aXV/Eyug
78G9SnNmKvLPcW/+Nrzo3yBPvzx990ZbQx9fflnc3hkAb+vhyobxQKGSH1cXIuKo
71nxwv9ZH72Su/sSgg85llyXAccwloLLqroAgn5lG5NY608LCkagWnTL56mOx+C4
kk39BhQFBTZCcYh8cmPvz1NhTLJ8OV7vEjGIOnJMFJ2b8PBVWkdnW6eze9mizRqs
1Pm+xmy2SMa1HGZbm5xCVHX037Pth8G8tR5XMP59wne4g4S3OgvpT4wbL2DGjuty
CsN0e5yFH4pxvWniRoyUIsc+rTxOqY1vQAESHuAcST1zFUt6p2mXD6AStAQeKoho
q12dJYSPiOMwW44oBHGx8sDG0DaILNRhjfoRaTqwPBIccn7yYzsPGJjkVf15LuY9
ufYchYKIS87t7x7a0XgJgVXJSCWVSeN8yQDfTcmzexeNghjAu8x8hUy+O1DEKSYX
6u/PF7B+vtpr485dJQX8eSvstqu38IDTSbkMI8KjSabeymuW5833l3kNQNKxia27
Y6FKNT/VTWdo0mK0yrL6v+TUp3DiGvbsJhbcx0Pa9SdSZXBTeaszn7ZsddXiZw5Z
H8ymdhCLIcCAKynZL4l1KVv8BRPn6QzTbEfaySBVllcOa9HEt+34FK8ZNn4ddOmz
Xv8/IIIFWypo7azqCong2yuwsc8pd7xUVQlF8oAARuqgwbkfRYsWxqBz2s81Yi9F
24pvTVlsm8BhoXToJ1aRo/MEpvt7QdvqRF86509ZyV1cSjB0ZfGZ2I5TDZRRqpRf
NrkAFzjY/p7sXug0NGu2PvBhD+eHKeyeOVIU4MM3vtmUgKMOntWhq4zj5f9kVTEG
wDB4/1iyo40TVNZ0pjkxGqT5QmaHEiZ1fSAJXyC2QaAtMpDSwlx39u6wo6mDsrBS
Idb3JEnXxqF/MJhwDdTnOuLYT1YVyg+FhrNuvdiJkrmdY2Mh8u1wEA6B51rklzTN
oMIK/e+BJPaHKNqUjMWS1NT4UAl958H0xgxHWCJvN9xXTV7Qv4MtE2uit/p/oZ7k
tGTCrrIaqLWXjdMj5ojJ6qklK6WCXeHD1YSbLTgd0DPa0QEY1J/oU03baINKa/Kh
Pd4OLdHnko5sLehXv7V9vXkAPRE8VenA4Byti3W97kUbdEvKhd/nINquwVAn5xUf
jf/c3z9bNCZiwHcLkc9DL1nHxi/ec73vjWxec1FcyAPansh9QA5edHBKPEBUgsbr
6CxRZqFtpyscMwIjnV+Qe+UlUp4tUO95vQ7ePKlyw40MIl1ws0dJPTv5VZe4nn9g
vtkpS4smBw4OrD4ZJcaBYq6nMiKqo4a7Pbyv02D6IUdgXHJE43StW22wfQEyHreS
alMVMxmQ/jz+RD6rMFQqVfUzR0+cU+03uTDJUzm+dO6+dqmCI7Iri+3fV/iLUsYM
1jOGIDriRaHaU7fExqEvPabx794HS2k4eT3F4E3yckYIiFbnHmVf4jj8//CPwAeY
0MQfcsnia6WqVn+mtCm3wCTUq1ixkv3VYK1JxidGkrozpxI4NYSMbUuvUJsVs3w1
QTGomuNiVHdypGe6fIp6wkl8OC1vn39Z4uW42TuP7EsbyvK1PGEh5JPjAzyuJyc8
xf4oFzI2n+uheY5AqfnoeRSL71vGgp/NETsz0JSP5UyWtGWAN6ldIJWpOuemBrNn
8arrhVfafaWLWrtIJWouRBhuD9NOP0E5mok8/hcDX6hVkB8e3l7fqm+YvfCvBvn5
9Y6zBB4Gn0DTe4imFeRFDhEMVMHYlGFSPSljoMslVValxFzsElS34/fO92pbTeYb
6fB3kpOW7Jnik2oApZPleWneOEV5wDem/2o9R9sH1qYCNE1uGPVinlXwTM1TFDek
C0SAzBpCqzQ5kM+lgryrzK+bcb/0SzMgMHwTnhZ0IOkDRUQQLXfA9SRFGa/XiaX8
Q3WgEBOvRcHcnRgu9TUxOaveYi5UzcJUWkYf86rGTxrCL+Y0ebN6mcO2gHZ5nUL0
SXAn6eCnNPQW0Xi/SKZzylB58+5mp597xoV0w80V6f+n+GtaqVwWk9CdBUjbmGD0
o7VSEjaiz4JdnVR+PNbbqma3TpNO6Bt/g2pHnQ9Z9yZdyQSY22IXQO5EqecFUeW0
YcrE7SZtWnlC9y+W+/YpRb7u3i/s2dPtWmt9+sZvNBmkKoJ21K8fV+6oo3ksdrwn
AhB8nwtXl1MdZvys/NsdtocbcLyFEExCrXjmO/mVRsryCfeOb5g/m88CCV754ioX
J2hNJRh5ho8LZSdxyAxhYL7yqtDX/IY+I27m3c2UQl5tualEVlGANN40GUgPhZTA
qfgWghi9CAD2Nay+TLckFPGw7zIr0OGdZ4GPkLKrFnV6xBR/jshGw0TmCjylSjn8
3ORShdBUWcEQGgc5Tt/gOnEf/WETDNRJfovAbndJiROA/IpcAVNpYrsJ9YzUe+oF
3Bn17zFhOPisANQuAZyBdDOAOd83zQNZOZdQeen4bu/+JtF4bkwErtcDGhZFxRfF
euEUiCPOAjy3DR/s2tmHkH1d4aFVvCWb07kInDy8KCI4WafXhncs8CyO43KhZ8Nw
z1JJTVmMDtzmEGPimjMwkzL/pBaBKLVpyg+SzPsNXrZvHx5IEY72riPvMczRKaHn
1DTW4XYjAGzdm5nqd1vjJJdjuY0kDDvRNweK+i2pS6fedXOLoNFwJGfUJg1xJgVf
e6b0px+vFZKYRb1sW/hKnahzMZAHBwVKpOEid2HuglT+BV8hAzrYrOaMNYhg+n4i
gNU6abaQviaX47d6jCmH5YlaY7Udt8eTwKJ1s6NRLQUyyl5Wlp+p+8VyuBXQkHNa
ix3wwUUCiV6WGLDQbT3Ia69hTkAoIX2YNqna1j/Lt5bjiIz3X0a5rAAdWIJWJOxg
nAP7wjrt+6DKRtQ01ePC1Ec8Ps5+V7hEbZW29qOHVu9/EHcSkoHiz0YHeI/IEb0u
xo13V9TcWykekCS0n1iP1oRyr4bOZTaPyiJkl1+S5dz7+QywpU5Je4QMFcDiaqMS
4RZA/EWkMpR4hi7YMifO2O/UKBkDZ09brytdLlv9odej6HIBTv9xJIh/axi80jV3
RRfWwbNGkTK154y90Es5Qkhw7kp1XFgLjuboXVxYZITl8rZ+o+Vq5np1sq3KY8Xt
uZs6bfa0WYRq8eFYi782Yq7cfy5svK7rtLhiXCjcaFOfpTrejPgkTARFtRXLtWbY
4foA89rDAcIs88cD1fwWuzNr4+pS9gr97EmXJ1zalUJBO+/MG7OLhNO784uBIOYy
HQ94EpIcp2S6rfmv1+EUZ+XhAS+JdFC3rjWh6YCVvdJKSRp+kyM9Mx4+hZ25lhmj
gMWjLm8KHVd4Uyk7MIoBUCsdnKPh6waYcHPkmasnpevl+CC4o/Wltr9Sn0Hwe3TJ
rn5V5qP7EYPVNJRjB2yMsv8W+EPbxqwq4Rn6ivMAL1s0gMhet0deT3tbjR1DX+zm
u6xb+bai5oGVftxkb8ubvmIyhWFsNfPYIyfUXHNq6TTzoN8CC12WFJWYduJyYKRr
4kgzsc+MWANCgFPafbOhR9H/k05c4PSK99JfGqoiTZWSTd9uGNNrmocvBohxEV4X
aV9FVleixVKAXSWrgX4VuBYnyUorR+sylXQXCeLLBDE4eF09MJey/3vH+Iuxo6+y
LJeyhEPVEAmM4MymjEdtDWu8VD7VQlnDRDpXcyqpOVVjALz5Ku00oPhzKaqQPkVq
sdkNiUjPdbXp0ZcmwA2wz08/5EIYMCGYmdKYWbFYJS0tiznzIYfWhHsY6/X4rsbJ
6iNXFmcNRG4jQirFbA/LO8A/W2jB2J9CR6JhxMzNcV/t7JoOAj97GXP7DxvQSjtM
bGCkwI6wsMnepEgAv2rmmjaniVU9KsK0db+Bf1ybgm0idb9AgPamrCwXu3R9rMYo
tLzfLt2ULgJ9cUOMCJUC9dHCO5VUh/gGys/KnRwYDzEX/bzPFWMu1Jaqry7GtSHG
Xm4MzzOa8fG6sFHfmBCX6nbc2lZVsB+bwTWbgghGgrP/RUMPLNGB9RtjXCNNUl+O
itffIqJsE5Tm25rGlEqHnw3cbOlAa8Nf6EyiG6A9AqeIkq4Br7+Gd67Lp4b6uJwi
FxZup79rfQYmCNU4OtfNeAu+PamNc1+HbI6rbmLCKHyfzIAZXp7fXmQiUFzPDaww
1sLmHZnZa6kd2I6UrJyVjiNSU4slyc8CSda+TOmLcCcDUJwNGB+Q77ehUolSwBQu
1QQpFqibFc5geKlgqP81HbhTvAgZimbLIR+tu9Tx4NSVzDg75SyVBRSeS/Um1+/R
hI2zq3RNHHd6sQgfT5JjUK6WDAcRjdV2fJYvqEhLJU5zTuwLLWlesml0iQvWYswc
7BbxAKWw0bZCF0/q28xlOt4J8mZqUS12q+i46E3kLRpgT2Ykp6fO4NyNcvH3CsAl
vtyXulcKEhPjqshzed9Jzi1AoOVPP7UGGX5gLZmtGtz5ewaPx0nVtHRXIlXXjWw/
PSgdZQos+LTDfmO8NCBLO2Ai2tDArYKVEYr3Z7rh92HjNHVMndr0FDQq2Eeo0h3T
IL8loWwhuizUiUbJEfUA5RaIFNiM96Jd5LkZ8ILqOaHZJyHt5TZlhZEKaDcZLzv5
Tq19Cu+64YEL7Zr777ep5iwgO6rrpOelmT4lgXRj0yOiU6Irb2cu85D862iMr+Gn
xi1YFFtXyNR4UMM7BMTV301b3BkCrYS6ZivmsZs7V1oHEROzFAzSu8gY4fVhQJh8
yAsxCdQ8dqAYhWXZzHEyKreNDWFhulWVtnDYRoihOhMWbJjkJSUVmFNAI6UqYGgi
+zBErj4+SvVP6Udx0LIkts7alnHMnXY3IOu7VMtc+/L6kxhkhO5C88X7Z5HZh8MV
QEntOU4/lLPZxso5uBJNYl6SqAvQtLPe2S0mh560eBoTI/MEue9mgRc080MYWh2n
WRWYBNLUJHvgyOPXFWgwYZDp2tf86QxbPjKOOwfvtTP1OOrJkrYSEwy7IQOCSseD
toAEJgcUjJHEmRgzVbjF4uVZ3gw7WgsUJy3HXoRs+DNZQ3AuxykcTrzWtAfCBIf1
iPSalGoo8uO8QhW6LTAiDegzcamV8Aeev0rcNR178HldPeyX8chnpBJqwF8/PZwo
9x0klgUIA/xl5H/mKo7nkpSXmLWcZKb0A5uIilYwBWO5pjU4IVSuNrzoZEC9DiJf
A+QGwhtfSB8om9Dgu5XS34CnjGAUyZBDvEijN23YdNw3jk2GO/obWDarwbk4JHuz
CvekNp2pbP4pYUfYQ+a4uWJyXJS2mVv79OekDOt6vFIGDF9k5NPM1yVYUYZbeLzm
O1AX/g7JSMTWVAKDaZD+Zz0G05qHNcKC+QjaXYX6GLV3QtbVATAYOJdKsLX8uNva
rbzhXAjrp8P18QN2GFYf7WGHiWJFNzs2h33Ct1hABQEi2v+RjNKVYn2tg6D5yreM
ya8d+rue4ELwx3MxOYdSNpHGZEC53FD0ORrs3qnH7kQhZjrwkVEbgBRIekZ3YhhS
RDntdi7/qhV16vXaDgMaYnDRjm14JZ4LEGCy3ehD7bvADYW9fFG7SdcCZFlxqg3Z
PjFyXzxL5tv4fW+/RWoW6P+FtazsU7At4+/1vijkELU2cGZdZsCTU3T74KJT1sfh
ILbi1RmyykIXfsgUEXU6kpEua0bOHXt6a8gS0au7JcKECtuhAaqGQq6xn0AUL0tr
Q5EoVXmT9UOMDaKt3qAoDioqoC5I/GNvNNO8xYGsTPH6us/mR4Alg4Z+OW18aBLC
tMzfGNBI/DEQCK0dNhWHWVmyq7gQskDQBhw2SekWdTSdX2BebXCfStG38vCN+0Fh
A/7QCgSIQ59KnP2r1OU5eL4XcBs3cVtNvcs700yCHVaRP0dABnw7SJqmTCEdWm9p
bY/sPrTCkvTSP6HRbV+A6bI4rnPl7BEAI3JuobLniyKQo9YVPpsLFLxxxTpigYrh
y2eLmtl3/xkAMSVO2f7uUnnYSwIpZDRTXB/PRr0R+37Dj3tQtJefim1oCscOjLZV
3cBN1LNbqP4a/ZW/dDQID4UyAmBgGDtJw5+GvQ0+b8KnW9O1qNrGbwL7R76QODqv
B0P9jXjJvMuMkXi+ytGu9z9xuH4KDjvIKiI8lDwp4xBQenIZDI2L8b9YXqS1MT07
m/NZmmbjk3DWrmIMfySaThRj7MUNUNNaWCr4ZGuedtt6A+4SGivAEDLbVjjP06in
pU5Akk3qdSYm0dJzSUGOAiqf3IyVjp+qvS4PW4/LWTon6VAWHNU3JoIPZpHMwHhR
oxPXgETs/hyZwgzlLyHW1VoqJW6gBJe5XIclAqO9v0NzRG1LvKfg5tu8NxcnyuDr
VXfAXkOJJp1d8O7mY6VbqLiEPvSDxqNHSpVUgOk88pbuuZUWs+ZY10ecxNMewHPd
z++C3h4k6hMub1oef8jJnwAOMTvqUpxcQ5LpocIMgQUSV7/Jpf9FRcR/BhTBeqKS
FcJdedtdl8puFcOIUA6kb4Y6rNOOm6mCGgV7V56by6ZM2k71I/XLqs4yC28F5JJZ
bwnmxrsJ/VCZYcf4S+o2BGEcGX/2v2AxX1yDrsj6+ioGFrCL7HMi1LoW3rVwKLyN
95i/g3Jy+SaJqEjOOa4/2Xwpwss82MChESb6nJ44pR8fLrF7e28D2tD4jPGKNd1/
jde3mlfdbo4KL27xSNNsY+KMDAhAOsKCWKG+U/Rfc6JSitUWCXDR7W95sHzr6gFq
j6IXZQkcJ8bzgg8NuChudU/T4TYg4pAlyoJoZ5W1s/3HiEFIkr1Dkx6L5geSZS06
/wvLur7Qb1bw2ykkivJZd5uBHsb96t6ht7hXXDoQ9abkcH0OiMmIBPbdNr9CFXuu
mJzmQMjt7i1MMbQoF/zB2J10qWIdwTI+FKZzr/zRr20CrURaVIZ4QNSO0q5yIRt+
NLqqywwSFCy5R18DCNPIV6bLO/MQGBjcXgyCVp7o0p6l+8cWUoy31cHa6KVJmlac
7vPMW3B/5YZt49a+Kzw4vUx4J6ESfiIRG+87FF8rzuk6RJ771N8+u6Pe8e31qVQe
KKVjqdrM0ncX5Gp4OOhCirz/Z0m5qz81dmlRiJqF8NeV/djsRn/MA5+f9dfylZLZ
8Ob0W8NwDt1AGgqWjVAdO0B1U++FSfFdpoCQyvoPIjz2sFhQ632uqVZPD5BOeePt
JlLU5Xue58sPc9Ie/1WLINZI43oY0C0FuAc4K+bxX51c1qx8f8kmeX41fmggMMA4
rE8uIp13JVYHkJbH5Rzn2UJODpYXTeeyxB8+7wZFm+UNzSYkfN1Xibcgx961g3rE
wjUszD+Y40sUraP+4i0psNkGJWxOk8ddO/YkXVRFkhNQGM2PvEyTn9Lj3kav6sph
AYQrFKVCe1Cj+XKBSqzhUyMXjwrwafe3HS5lhSZ7iOmVsTpMUKwtWX0QsXqRk/xi
/Lt+tGm11MmvySSrG03iCbMk3wkj09BE5cYzwMJOXE51o2sydLfTUq+93vrom+mG
k5TqqtVl6L7QdmrOBPMwFx/4icBEDNXuVkAyvfk/Yb+tRs2tHpsaorjg0qBx+/oY
72ekv54Kxp5DL9ihhfKD4SKWPRiB2+T170CdFP3nTGpkKNLXrzSrmhqTKirhj94A
HHbKP6VtBUgrS8hY/aoWGV3xXTHfV6kueaPsFFUHgbdLAe43KQIPaLT4iYGDBym0
B9lW/0qtldwv2TacL+v+QKSHAoClqXsHBEmo8HIQ+Wn2ltWeegTwjd46RVfED2dn
zieGs4IGC4QBBSKLFhDZIGrgy6jCusAIuGErtMmJGN16/5v6PBd7dPYICtC5NI86
joz8G/0/fNgAlKTV6UOWsHx4dcH190OLvRU5vK15i5pDOF1l8GevHhJ2eEa67zS8
hfaChLyGQxw84VzAPZJa1h6SfycVFNnSlXzKnUrqH/u2mWVDoYw2KaXSvllGxiGi
V4ybwF9mFASDPdAMoYWbRMrLqbC396GO66YK7b8rDq/bZcpUa7GSuSKo7miNppJ2
9kCgs+kMBlfJBd8B1a7SR2iIhADIEq9BiXpmV7g16jqxscSmPjc5+XBjP2ch/2dl
RcJzIoqHmcC//G8AA8Wm4GkUz9O+WnMneuERCyXU/+dg4sZmfB2pUg1oqWAC1Cu7
icTtwUdIz3oCBthIjDLQUm0bGD+AJ29Ak+N2sToNYWpIXIEowQ1R3yKM7RRcdMFc
cJlFwJV057hb5OfF9wBzt+QmS4aLsyIjwefsGhH2a3CTEKBLHd28WGCLxPcEc2Sx
d7NL8rIre7WGf0zAwKjwQIFAojJulcrx0/SzuAPBl3HfreHbKEkbEBVkP145dKLf
B7J1ESGBH/5JBFe1gF3Jn8bBaSE6d/GXZibJmli3jCtep3R5VMlYb6kACZ1OQZt4
9iiEyqgFuEj2NOjFeM/plHb1cgnihNXTwfdR5gzDX8PHB4vphLsq4OWhcIYGlaLP
FPJlAZ3dP913uMsRlMbzYZLiqfGBnjdM3fN4xpr0wDfTuJ2UKpHnaz1/e2rG3peJ
1g9fPf/jtvMYZeRQ2zuNNPoOjGAsEjVxOdW8428eQgxN8Vpw4kSNklCbCEKLHAXf
jvty9ERpYCCm/WaHfRGz6Bdd+s1qRYoIBjY+37cxGjTF5YXL0gcfm8C2D/dpk3a7
PgXuTdkSdxBlp6pGSd5v7NxlyOx15JzJzYOaorinpzXDhUxBEuTz/RL1Q8x6Lyne
WSbAh2K+nWdAV8Wb94uaxK3XvNHep1qpl4L+7d2qLh/wAGt/rfdOi/si++q5ijM6
GV/Qagw2TW5Lzeho6dGWV8nRAiERKzNo8zmSafnJj3wOfFydI6cBqYLzHBamP/ir
1ToZ+adh1CFViSuUj8lrkALb9h2cyULQvrYb3QcG2JNo4uRI0+n5Y4pdj+sjmSCy
iVXSPtGFzpGgy61vCjrWBru6OdFEbT3ko1kd5+5J4c4ITwSX16JVnb6R77+sPP10
ZRCQheaeJCunkmc70eyn75BHWmpHKQJkg67AvKWIgvB6OfxbPO/G0IprVOG9dGSc
im+i7cqfF3vG3bgbH/PmMOhoBfKbUCiEyDzJpkTzOqLY/xibIsmdbQ/tbgy8y+Bv
NhLZag/QBcYl8X7kucd/3NJE/nQbZ8C6CSL8SUBYmxz5yq5DXdiTMDFZTQSfGab2
5LLqKlgeAkM9ei0dg6RJnLtLvG1oXsQAeQezHYhyqwpsgBUH8UZNdke0jy0xBwSz
u4/BW/VgZZRhn8C/msdh14kaWineGOMnk7MKBy6COJ6/EpduLDH1JJ8bNbjU5Yw1
CkYVtzSnDSmW22+MUtI0tVZCn1Oqa9Yr5OO+StTmj7M0LeGY1wP1EhaIiMxTaUPZ
/8KDHk1Y6l0uE9PnDIOcbzxszhBzI7Nooar9Qj7SGr09h7eGUUqtyOXju4xjj1HO
RnzSQshZ3gSqYFwpdYTUEbxDmYOV5YQWBDyNg20RYqbdhu0FGUj2pXjuhlLIGghU
z6EkiZC2bxkEibdFT5YcHJxFEm/TRG26DPGXulb9DT7YF7u4eTY+YwFitDik+/Sb
7vDQ4SWdzWdWbC413jt70JOQBNoX/HuyHG3t5vBZP8+B0FDadKJ7VJi+BCL0ss8M
DkJhjQH5p4sA+2cDE2XlsAt7uuEvgZNH8LbMZfYnsFzKhb1NnqPrQzcvRf9iZix/
v9EMSAaEsWcq8mBs1pQkqv8B2KVgdDemUiPk/dcj7yngmYhEqa+gqIfM8mFcgCe+
oG/rzCqIBS5QOXiVS0Y7Uu4y9CAMKUPoyW5jO8vXTtEsS0QdoAM9bP07+w5jo8SH
t9u+p0fnKPVKjVIJ3cujI73P9nQRvBLkLLuCuMa96EjPI6akGqe6oH2V70GJO6rj
C5SV3T6TlaExd0xAWgJn7IXLadVCO84v7rLJMjBY812hm1XOUYkGDBkLA3lhZEE3
HaY6aXk52yPd/czjCPxkKsa265I/MtMqCR2Qe3lUVcQ+djEd0MlFLZfYi125YndQ
TmVTYGf6Efx3H1NP4ZoPSk7xyx2Iq987TWFmJxPX0AVfUQ4H8WmW7PGCtR1TTHGB
+lf68uyhZVAfTEmcqWwBFvBTjF/e/eV/8CYuTLw4k6hXwaN/7lRQhMvVJfd16tyJ
Uxt7WUwTxt5eProbS21g1GiiInOiPrzRJKB2PYV+a0kZDjli+BNE1v1KYOsp67Gf
Vs00rsAlj5udu7nmIBvQRksIwHKZv/DAzYVjioifHq4oxtcFvdfjlyzR1CCA1wiw
2lLg9eIWOzYbGiMOCLVG5UdnBXkIaC2RIA0uSazwhh+pbE6EgGm/T01pKcZXHuuz
0Onjc+9pKtdwZ+bfZF/Xwi7ykmCTErUO/EUPAMuamJFws7NShH/c6pcIcYdrLirw
nXOmEy+7VB93xgbbRE5SElA/RDngIHw15L3DJnLYp/J2s00dconq+Bd5xJGYSHWv
t/YHFYdGF4lATkEqCKUxr20q4yAAK0bcLBrGi5JwLKOg9T/7K5Z8Wf63iESUs5Wv
V/q8eMR0BfpY9o65RB/fq3KD3abQTRForDC/u46pWhTTw3470PWpVT/Wl3BirbAp
/60QATtNwgxhTzvipObfExKFqJ97/jEJfrrHjRsdfhp4EkHAEQeVZvAPnh46utnv
m1rAszdUKTOZI+1g8fG+kqTeXtEoVfmk5CZUNL8MgQdkm9IteztSMPiQhjenMnQA
5/YMviBmgIRbBSq/HpmoiAYlILxPOq+DfAP3kNyxVFpuRANZ5gS/AX9oJPjF0Baa
srPXglPdDAHcBo2+ktAtBoN4REckRwqvAzUZLlpHtWgQ/l+u8MUvEoWC6w2nmhHj
xaj2k7IbC0lNMqu5yMuXa3k0oPOCCwM5bkcuwwFaxxMajSEQ+F98Dia8i8JtJ8S/
dtAiLa42AbuFtBl8LqGgK1EHMIU7LhD6kTV69HogxiZezjmjaR2PaE3aVQp4DO7v
gJudMv7OLlardVDc0o0xMeabvt6X0m0qICPjkAQwAcxCkFKYUgC1WQAN06J/TYrJ
IryxjEk2qc2Kv+Hrtq+DuxjetDW+XmQzSKjGsh9VYZPVEqBHxEs/K1mS12wqpbyK
9y2g3dxCuNOaYInjrWJ4SrpF6aW7fxEj05mZsxmK9BEB4PA3YSXfwW05ueEunYeJ
uYEgGm/yebmZXRoMG+jNH850A9v6lHmDrPilc+TCCKUJh1wGCfd+eJRd1QUhWIhM
naoIxix2MBmiBfDwfv/OQwud2QKs++sBKVuMbEboMXNRNyx7B4PkUC7KHP0dgcmA
/167+dS5owtiMl07EJVzmvScQfK4eCfHk4+uUsNzVJjgMW2EvQaZGmgf5MiBQ3ar
OoghzmmvnsQrRb40cieptxlcuX4xJq0ffvOTJTFimiLqJe7qi+s32zRKq7ysJ5uM
ArQDq45xL3t6nvrfn4xvTpGDQGfbrgGpc++DvY6cTyA84ImAnyOCUxtaEUI9wNJE
YMFm6CdVOTsMl4od31stTDA0PA4/BD4nGfVO6wWHmWDndSA8EWPnHe0J5v58FvBl
eauvFbcwgE8XsrPEZAA1sdiKR79WAhG0nDXDH11NjQShrIVFYOzwilttzDcO00W2
izb7md+PgqJCInIE7B4TRnxtmRrtpr6x0xMZqZwPObJHINPFy+oFO7hM2jt7C+Wy
6t5O6nGJQP4eBYjurBdbpScB6fe/T6MzJrRo9SVOlRqj96bUEvW6/Oks9mFKs1Hi
XR6X/99+0GQLs73OlgK4xbGUenATDccIDRLTifNqx1EjZowKB/qp4mLorm6YErEq
6irY/ahY/USOLmgZMteyjNm/j/iKwcXEVPH5T6lvA6aGjgvVGib5UhILj/nV3sUn
Od2zRliAglCOx2Y5D8TPjGtJ7BmOlYZurGsx2gd5MfYr86TKzOxQIE9wHdcHUQiY
B42AW7cxpTxeQZ14JXqQnqTNb+Va863ShVw0KiRyTslu8KaTxRA+HPOJFzE6qnWp
0yAOyfzEpjO0wel1H3bOJ3hkXIk+g1ousyiKxA3C6tL9fkecQUyM4FLkMAEJLEnY
V5yu//SA2yA7d1X4N84gYNtqu6NGzKO2Tul3SSwPuPNNVxS++wrqy0xbplFxdNxe
EbVANXk1dDH8YsdeFdLhpFmPSTxmjCmlMfCb08EKhOSVYVMFWgcJIvUmEgNg9F3+
tVGryFkkLSqM5ckFZhkCq9r2j6cCmGZ6lQWr9MldaQhCwUrO69zoi51WgR1YTUSN
YFeW1V90MhX4k7zDGlT3pm6+WZf4NRuBa8JtKVMqdUQkhqHyyYaMnp0LsiX4Jke7
QSgot/D0yX1J6qZoz5LfU8G6Dqa6mmReHJXXaTLI5njIbOLveUEFsVNy9cBTnzg4
9Yi7sTCtgdSdAPyaAb90S77eOuEOyRcmsPN477FsS5H0YqqcSbk6AJqtuRMtrusE
ZulTz8k/ovheygJ5gltbvOH+IU8NlHqYd9+JRC2IqFjc7pPg95L318BIHB6MRtPy
yl1V7UVkd+JoVtjeecTDGzQnqtfEgpI2k16S7WRKGn1DfLAJzMlPlrBGnsd7JGju
wzmvrKCZltq7Bjdce2LPWrDGmZebXwq13d4Da3qIldQ/ZCJJDcHbyIjMjjRsopTo
D8Md0NsW9fZ6RAS4EnJSss1TE68korWnKg8SSexVwzlajNqs1VqVCf1cq2v+QW8S
ATQQyQFM4CYRJvYNX2c+rWvKLGI2Zj4cWXFXb+MXCOFxW57X1kfG6FFcdj48b0Lt
YMuZ3qb5sHa7NnVuimwS6Do+c+JTpMcqSkpPw/ChrInDabCIDcC177oBuQ6e0z10
jSWXEq9A3253bsTcSHKURuPE/pVmPCYlJLlGs+YYTrdlevA7VzY2aoRmPliHHxpy
a/DKZ0BzlSvXTmFkxUkcqmTtjnv+7SOOcLkwk/U0K1rcjHoyDoW9p4NxFRAvMIrv
HdAensH2anUdgYDTOrOAuBEaZ5JFfHjIC/wHvL+Oq6VgPGl7cF/ypc8DTWrSBDI8
1lUtg580ar2SsxpE6/MZejvimwT/eRUoXyljOov69MESgqykumneSRzj8uQ3cZIM
jsk9aVVgXKAOwHJFcSD6KI1gYLyzslobPlbz2kc2pUojwCqDfYjbpuq0BUyZyLs+
i0O23ZrFlk9wKRzwXG5UhsmsjT84EI1fmilH+MlD37hYnamKjbnaVPROKkLsyzna
JM22WRfxzvDOaRQoH87U1THWFoySWYf+gFvNgbKqQO/Jr4j3LpFw2Q9JonLQpTkd
bXR3aSbOGOMxgT4FiBrXHvi+jILEnSpwskwQRg393z2jCFAkxx5Ldj1t8D2tXuc6
RH+nia1e6M8NbPdre3Uv8dFmayUgwuP47BEYjuKb9oW57Y+X8xGKZuxRIj8L2DWn
OktCT73qrMNUWMzce8Syb0bzSR6+T+10p3ZItyoEvNQC1Q72V3Uno2H1aU91CDtO
hL4q7kBR66INBprLIByRj2LHRwF/FY9P2a1u29I9FUuqn2N1+wdO2RldI6Plu2Jd
JI3wYpq5ld8Z6wuKPkj3fo6+cNhaYJ7mBNS92mXE0rEB870G1Ovj0ETUcX5mIBP5
glAdQkPywuqRKf4LSfH6ectin4D+ruIusbrjVT+iRUydvRYdiY1c9GDzQdkyWCwB
+8gUy41Po62sgLsc91qqQH+kTeG2caODKyog9PWpKIDjvmyogfYY8zeEm19WpQ4F
7bijnNspgZmw1g6OGj4pD1qqPdyxw+vxO9ZE+PPxgB7QR2RNBM/rTgp8XzR7p/am
gwQpZA8/6RMAP9CQNHYTZrdn/tQEIRx+ZG5wrcb6iNXzaTRwCmYlN8/dFGUkWQZA
F1HinNVX0rHXUN7GfMEsg8OJy3gjg2doa1dFCVHC1xX7I8GwjwTA/qKWKsQwslyP
rR8o+b9Epxn8+SpqvfEMZhpEAP7fWd5AYrer5XB6QsEmx9egc90vl8elQAALD/Ah
6PNVJ/xHAUHvvi9Dw+Wwl0QpexFB7mF7ia8YjVeBlQgXFvZ+V6xKap7gdjDvclYf
g7CZrcgXKe0CC1cNEAmyG3/tn4cvM9Zi3KRhwrwLDZcmZ1uKVMBaotSAxnBIGout
1xhfU+SRkjWCrkRfR165E/skHe7/27rJqn+Ary9C770VB6MG2P/Uigzd3+gyfliV
EN6C9ZMt5wxzBD9/s+7dWa8e7jMhSVwhviJV6RuylotRl3nSwue3RNycfVNHHGWU
5DwoOtlSDMYp8tkQ8eirIAer9BGwrk39bfn551RoT+xH9QDpyMDyWi+rec0spnMW
W8Gryko0pe2gQCcsYztKV/5Y/S3tWdD77tzdoJtt9OpQxalBil6T2qT31M4hXN2f
XBRowlOnDabl1SI9qEJlbyYNx6aDpyFFB1vFnQExuWO63DhTa0umMPYG1yRu/7kQ
f7/DrS42YGRtGFSnnfeBhZx3GHtNCXog7yqm7UgZOllEf7PF6eqdogEztnW05D4B
SkF/B6qKOLnssz6vcPyIKUqWrYAgC4AoPnneIBRIiBjLOsgzuVwRDdZPxjUTjwlb
r1VFamc4tPMwB2/zA0T8Vcn0zjD9A86Ks1TvdTS03jy3k4HKMzGAIdcUQIlRC8MZ
XHL8Fw+dLkQVlJMOK2CzOuymkR2KFmQL+2IE9VkDkYQJSEAq8XBTKlknVFgO7zug
K2C7nUvuuBp9aH+XcDGFsStRoPWueReWU5KS+PgNkhRbbw0WqA09k9Ckwcz13ZJ3
xHKTejrTyvkw3QygSD40/CsVRikFB0TDskM5CNC9Hi1dJx99MIKdMm0kgIQnj6y0
Qn7MavH7DtEcA2ESJf17OTgpSIgae62mJTo1orXUuE7Wb3T9Q1PkqdpwLyC1MEfO
V4AEEOofd9QEqzu3vaAE2vmUEysG50eLKoPcWxYoa6tO8tNQNXBXJOjR6rZny7pP
GTnaUYlzcY422w5xdx3xlTNKhyVAcQcScvHE0YB5DmzRJbqNnEOUhsl3pdojUycL
LQ8Us6PvWquNqReEuk/k97VJYxqMPY0fG/KzhaA/ZgUfedx0Qp+xaoZK7BNcKSsr
O6GyGrasgVlxz5oRWFL44BVwgCN5hBI8Ig9WNDeG/OVYxAmFZYhOkdSCBZAHBiRk
dKXhb/E7hQ4eK56Wz812vDiTZpbQmJSu3Bb+wS4nHDVhVU4s3stVVE0fDMVJOSve
EEboy86WpYge8TBZH1BRKVDZvdaekDDGwzWNU13EsENbKntF16O0cVubcVpeL07q
5pACUp9cFD049Dv++Gxeuhm/jNWzqjov/3TbBrdH3Gt/2iU0TmByg0MM0ycq1OmT
jSa3jRc3ppfTpTkiJMZRKePBL2iDUonF1+z5ey7TzuZtv/SqI6xWa6+MMp8TnG1O
OsQAfSLqPngwrH5O4gJRrkmvZGnABbmfmOTitANJMIJ3S53gf8utt1iiuYSC7TjH
tqdnI4UIQH2MN0ILdRrYfOC4gq6dY1GoCjCVX//mHYmMcicZ666Ev5EbH9kRVrdS
9pjXoUx3aanzzaezyEm9iwFt2/2r++b/6KXP7jzzia1gk+pEqSuLIx03UIn61HDo
ZRt9aSb0Ns6PWubFjz4u9pLyj+jVBT97wWbRvwwYfZLTjwewZxdb1PyoFkDxJeI+
hjtjTYdU+DZsMrlR4LZglVWxmhYDtwhp/acLFGqkoKlzGo45ZVP9zmI72Evjj1q6
tmHFJu1c9tTWJKt+r5R3JWkxAl7AZ21aHjWxPEk2X1742jDS1LHF6mjM6xQcxssN
Z8M4LD2IPPbVKMBitFd95KdW3d6XIUjqvGwu2/liTgPGBfe/jgrWDXxaOtiQjk6S
79Uj7mTuQ/uSYJJ5Q/EsUmHi1vjO7+DthU9dVB3Ifeljh6RFb0wMH/ByHfsGHA6E
VHjavuaJsaziBYs2lBxP1iXG3Ev6nJ9s+dGaYaqzi2j8zZNUklRzYIIm0usa+f7K
wpeAw/3uq1RF8t99YJtFjMRoqnYDvWeZkqpMhFaHEnfyz34Sh4nFxH5rPC+SR88W
3nOIqiCR0H40r94HKzJW2Uuovc4nLsX3pio6ztzZC9xPGA5pREPCFo2AT2r+L8P0
cLwKETRlXyWERKOYWKSVr2I50blsucQwXloPniGHYy4f3t2gR/N0kFjlP6zTjzGd
f48DjsGG9d6bIj9oi/gCyxVBCrMzyCqaqomc5GM63rhQY1I6Vshn7VGw73+00v+6
wYmLfQyLD0smLtv6LVU5FzAtcupSFZlFKPGimKU9a5QOCKZAvTrM0ebee12JkkRw
QKpgMfO8ME+cuVAewsntk5ge6duSepI15XbIeys5RYlxBDiVmwhHikIcQnR4paH9
2aQk5kdakKDnj/e6hrvvBdqcy0I9RoiRJqDo74UDboKWyEehOuGgY1YKsX6CDGJJ
mkwm2so6oNEL069OKlqq3CnkR4+r8RhgGCyh39xOhSVYMx33PtyqpWXQYgvkBSJr
aDelfQdo1A6FC0o6AMydyYIggMsH5Bbnz0RiIJ8Jp8tLlAeY9Mvktv4t0f7G3mss
pUGtRB3Sx0nnYUMYlvHHTwlN8bc+xZOdW5EQV9XvqKDkh938ddt9tgNcWWG5z66H
ySws+sZeZF9FCakM7SzPLA2J9QlF9xLW7BN0Y7ZAFcmxX8MRzqhGrOzuvBmCHgrV
D7/zwDEnFsWm9ZvpKhJ6jRE+cIrM9jQEL0+G3hU78hPlAyuiBmUj+YXxKfxZx7lJ
+8ZQVpC93jnRImP7Hdp6ynZIAAJiqSTzvRXZQ9KgcUwqcN0ABr4AWOYP1joeNigS
lQytkDbJCQYgE7zzuf4oLtSF+7Z1biXMCbbmLGC10pnTVDf2Z5eFoPpIeI47gAXZ
P+/oFHCDhdQfWfJ2X1+qew/dtya91KgRyz7K3UjopKip0XBTpt88xzgFakI/nFeI
16oZLhz67Bi3MEmK92peNmXIJg6CF/BYBrgxMjqHBP4mbdiUueE3d87KeBfgVr6R
U9ReuyBy81kdJqSlRi1EZAePIyWzBlnOUW+GpVRBqHhv4YmF/TxxGMr/WIT2n8f6
A1mV2A2kc2M7lvuim7BLW9PxPMhKZKAVMd2ZY0cmWcZRCmwk/mu6E9gIsiU7Pa6w
MNvNgOI8IY04i3SmVI9//AMz7A0SkQV8iE0u0yF6S6znzM2UxPEo3VwiaOpIO08P
/UGIgjBF0yytiCe93tmXH3pA9QRO4OdojZ31DhUrvkfB/v6W3940RJ0uPiVVoFHY
8gUYnPEebUR6+crfFm+SBI3sVAFY40TvlC1PUC4OxNAVr+4DxFtODE98rqRTmN8C
q8coAja2sgz9ZgGghl4wQbgGMY37BAHHit8NcVYEZwY/PiziITpmsWemLujxRHgk
H1c8DenjOGwQF3qbXX5TT05p9zg5RIuXUQwdbJKkYK9JhOIRcCQjU75usVSMfLdA
ViO4UXOPGia76lWgIn8mukiAUPlGqoEXIw9XS6uiQG0ek7tRSaBevmxelnulNWfu
C2Y03BR42jJgBJACWv36ahD4bI+g8HXgHnOdcoPwjN3X3PINJPOOBgkiObz6dbnN
Ju3dFwIZY5CX2tHQeEQIl1PCgIonsNThDsARcKpaGByzA0Exd2GcWvgW5J0dDyJ5
eROBdg0gdn7UpFVJsTLPhrsognO0OdUB5VmDPyLsKqpc5AKSTmRSLHisg4yA04gR
U+xeQjaJF3UhgtTZJ5WkF2rxAgpnsHj0y/R1haTvUTGLY45rsNrJSX/oVpwBwWAX
0IrVtcDXuu2xQnRscnRDq6XTg8pnz45FRW8PfSpgyXpZkzs71VBz6z14viShdY3w
S9Ra9IG2JVS4kMncd03q8FT8RNLgtRuAIpkHj64XaxIQCpOsnAQ+yP/ZOhSg/7jG
yqTp4tLXQjPMAg7k/wGg8SMT1yYqDaDASpGiMCStMFK6qpTUNcgdv3mNRSC5GHlh
rc+wN5R4BVbXvTT/qpOOh+Hs16ySzHAZcvSR6n2TdH10SEjmf9mhwLs2ypbk/YtK
KEGjTU5h6RT94vKu63oiqvtErmUVGwnuee6zdTzQjyHGPQAIcfsB7RiEoWEgd/lc
aJo1wqCjEY8VRW6mC3XRbyy68IHHfA2gUJKUTXZRifCwm7ZiiT3RktCphzUnrHJ7
AMeooFF6IY+Wl5vJgqERtFHxpeJDU7sEH8pZrvMUZLpbY4cmhH2/sFI/9nufiZJN
UNOY045qn7UAx3q3/bxDh2u33j7IgX34OpzaaoPtCtb+iSUx0ekbA4hiacm/6BVf
aydgRQ5lwxASkTMnI7RlV3cuoHie1WyKGFEGzr7SAD7J6dtcI1nj0zA8NPA3z6FN
+OsAT7CrWaedSyS8SBL6+XuuwEs0gmwzNya6gThkcZiEIvhAdCFskse3xquNs+py
BSg2QuI4ewfJFleiq4acNvhMsxv0yzZ9R6aTllEr3xEZY9igv0CiaJ3/H3co3RHV
Z4pLc7F9tWwvwTjsjH5bHCNdiWJSE0ZMp/XYOoxBryfwmoOxmyz6mjq30zDl/cqe
2rxgGFkGhuNatuV57Gu+6XPtPMZW4os7JK2iQOkNtQ81A2dVqlPXapg/kvDtntwI
uA0x+CTP2o/lwv+LbsRMaT7unppTUyoUoSVtvmFEn/lBi+BGIYMhdsIu7PghTHPc
/yn9+V2OT/51HfT/9cGkqc7pkk3L1goqGcEXeOmb6Cg8XsQ0S4FjOv2ft9GvQZ4y
wmzNVRlw5zXiF51S3NdhZBbvRYEChPvO+A4oAYci7oKPyyDf9whQ+R03JLqvi0MF
wmggopjniBizMgfRGXhRJK4A88MC45wDXhf0P7F9bGuHSfhHgv162p+Q/0kKAeYL
xR3mqCjAuWL0YIUY/1q1+rvGZNS2w/ei1EPvyQkyskROBXPH3FWzpqs/P3hFkOc2
oy6FBaThNYuP/l0By+EyBL56IdJvnL4MolDMLz8yEkE9upNAcNbj02+9+5Mw9XlU
72Tnq5F6rmjcYWduvPxiSpxy13ntu6JmzgnzQZ3h3d2qFfyDzOEw1DphBEtMAtMs
FhoKIahCL8XF0ux6LUMmflIykSIlEe4r+CafLT6KfwI6ZGFMV+AOOA5nwQ9VJage
nUv5O8uQN/Oi19Mng7S7GW5DLHCI+UMZUqDwf9DLuoahyutGxEg/olSzPvl5P/MV
i01GpX0SnycHuFctMlimgFDp59lM/4wVx5jTstuVtNRUQuyu4V2TS6LwjWKHEVA0
mpqMTuJgsakOlLC0iwI6OGBOVEwWpPhaEJQWcCM3Qkgwv6J97Wj+ZkYOO0fMtCHj
kn1iPSdiwrrBLgcRb4CQAM/bi3JNME/zJo0cVY2P2Lbktd/ORqvwPZRNEcgSYRJo
BZfprndckPiMq7dXLznl4jIiQ73cveV9Zd1wEJxrOgGPjJ6Jsi2qarx+jjK7KJlo
wK+CHOlk6hABti9ywwLBL7uGr2vFU8F8hMPTvzj0hFqPEtr7z+gyOZKAhtMj2lZo
dQ+iq1ccESR3l45/KRPBa9wB0Pw4+4JjWpVCijL3xmIRfYQdBg0qggakMQHUFZMh
WC4dE3wcelxEayUrDlpT14jS0HrLqrXqU9/AqCV3LPu/9tSkkraUtnt3BbLwOfia
uNL/h/tyNJwH46le40bNbDC+Xi9NWPBDz9c9n7IUdefD9qzjXzlcfyd7oVctgcks
EOlSaZIl08KEFlsN8BnT3HGr9kwZi8uxMvpF+Y8KSWR+3pED94Aav9Y8nlBL7ceo
VL8gxwC2qWs7KuUcsqOWge0DNBeLxIH+Gl0/lVyIACLxo9tfnQHzF6iWcctRfMcS
9QG3YWS2AEcnoly/x48Jz38H3s+TevN8Ed4JnVlZrgk6xSVSIYCSvPZJKoSKfhIu
APliTHBaI47arbdblk+hyhCFgWOGjnW6zWLx3/640Q7ppDkNEOA8Fv81ZneTk9Tz
zOFFUph7+uByjI0D6h36ATopeP99Sw65hpHFUjQXvVkX9yF1kh5JERwt27euIDEB
QxmSPsoEQ+hWIzjBZL51FPRbgX5HFuLCbhzfmS44Rz+klmmrkMxc8OCthG1BpOkM
bNxGT0eKc+CrVIN1uYbXu5JnbKsX+vOwMUWYtli5uQ1lMUZrUr0xFkgWm0kTNCnD
8JzpqWyJL4PaaKxCKW20aYYhYL8iNlMeFrm62X8Dek5H9B+qKF8G2OCbKOzH+DLz
IC+a7E78tnyyr2G1jJL8CFfllghlI1QKKfPT8u35OcFvjqBhdiEorjM5g6UrK74P
8pgOXkdKDQU69m7UCDc57rrCzLEH9hxk1rjqx60+SZ7bkK0sPkn0iYX3REHiV177
d0ZN3xPbBwr3k8pxO/ly/PGNyJCB3YGw6dkejGccQXp6GTTq0U7hs95v3IZKCkOB
pvMg8Jb2sNdaBcZ/wxo0oXqKDBSYrJ9qAP114UhRrZufIh7nFjd/JJA48GTF7Ikh
RZe00sQBZyljsQGcTZoltJlHApVvmB/Th+qFeQ1op6tDTc1VebWNZNTIg5PHOcWQ
WVzOeppxp2A0n4V7gxSNOCwzBUzEtgCf3K8bwjmH5cNeTGKXHNcSQz0jjTAGF056
MmmVtO1P/viUkTN/i9hXp33chMgjr4PYbn6TziRTYHa1N8O/ptYvGcDiu8tBqyvh
exgDUYQnKmY5RnmUR5TidkvnC56rZfXEOp9sK0fNuJgg0hvI2zCXwKvnkMhNNdxp
g6KApsuCF9O3DOg+BPHYBG+yS2Xsj0Tr0D4vA+U78KeWx38oNCKrYIRvhsTfECZ+
MTBmNb41vBUGk5FcqpRv8McEA++4zApBjrvOK8LhGwmJymCY0WvhtImUpdUw212P
XUZhJBN5pMNOhZJOjL+o7ZCpq6pwp0mtf0iIfFrATkT9nbLFCHoamwKE+0ybjP+1
55baFpw5GvL9hRpj7K1yUqFOq6YwakuVExMtAzvyqnZg12+q/eulp/eiWSctL/+C
gP0frUl2Q6EUTt3mql8zhrL78oKjmsack7/D8ES6BXf1/ZHQTGswMYb2SvqGYVKU
qBLmtVrCPBrLi1tlEsNyXNLbGJFmEqIdOvWNQFqEGX3RlqXcL0VLe2MbmJlwz/p2
QLxR3+U0wSFKsZs2mwGx/NTJUel7ifDnut3sjIPRUUSFrIi/XdM+l2DmN+/6wi09
+GPi7pwTwl+Nsp9UwLkMSGboIQLATD2HY5ToC7DgRlqqJFhb6S09icZ11pHkUql/
EuXWGDqBKUkushBhkWwUz73U2HGdF3XgYtiqcd8O2TUpistEDLzuOYCgs3XhJmUO
mE31z6WzzXD42+bLWejg6y8IBLDhyNWM5HFnJiIU4Qv7+bTvxYGg8J5SNbK5qUy2
haHB/BnnROSPaKfKm0Ra1JN8oEgqlFdchgns3WL/d3wqoqJRwVPBMWKe8+EfFpPw
jxNlckTROO6TAbjthD75FXislIDn1LIvf8BxtXoZ1X8bJPfGS9MbEgvwKZblQjA+
ViNMkg5vF173qYnq9+UHs3lc13c+93NoUgQCoSIzRwgkNSBSJg6ARCZWYZCeKdW5
dEZ0/RPgFK69Nidf8zFZ075SSYJmRBgxbfSrCFVm38y4kholkaQQTDLVYaoWGmOw
CxvX8mTQY6PRcQb36degcG8r9GWutDwP0xrz3kfWMoSdq0pDEv38fGGMH7Mym8Xn
mY39OtelzIy8U+E1aBhou1uwsUcJgrOWM95JWONUEdrMZYPkhWRjTwz5cRhDfyNu
By12F3T/qRNJbgUwdzttb4cGr1R+TTLw3O1DG/+S1gDWsOy6R2KpmMJOkAwyegQ2
zx8y5EMenKRC86M8DlQ1i4P6aIQRNiihsGNMcTa7vYE2lg0HOWDh+wNTw9MRUwpy
S/ZSMo2wFW7Bs6gsWyUfWLHppwPinhx05hTNltG5/zpKAcwfzXGlOPm2zrCr979n
5FStlZ1vZBuhUg3RhNxDJCJkPYJhcZC1Q1lv4u59pZsdUt2wyOY+jk896nbyZgE4
WscLtq+dIPY4Rcpzx5tMx8SpXwvnR4y8X7rpmjKGtQ3o6sThnYGcg2N2HyNp4hFC
x2RS1gd6zTYTjcvncwRDFTrzlr5fWVwdNpMvCsdW7hlitFqsq2iRnrbx8zL9F960
l85TQPj0qkkT21PLLVxsaWyheRCZ+uDhseJDF2+IqXXw1d1ibdX+auxWbBKJ34+B
DPraHFLk+9dn1505VQaxJwYRJ4/tfhFnNzFrdlUvtPunOr2+2qi2Z7LUtTkF/KdT
FKgOwMlbTwdxQe+nqtt5L1+vnO0BkE+f0xeddJx919+hMWuB4w0w24p0Ta3kdwXs
lZNKXexT9cUNQez/ALL2W8hI1Na8sZwf6N8OwrN85xuNqr0ASD5X+NMqzJtSQxLF
Ooj14stxgo+rasHRwh85gmqpkEy7cuEMEPSAvme3hFlceVoGL0uqhIjxxPn0QjwG
2ZrYEnbhsgLy8Y/dvssOu9FIoXdEcqYFQ37WBX4UdrxKOOGKzqLGm46Y7sQ/eib/
Kf4vOl3e8nqME699zKYzecHRvYk6SazfcJBQZZXdIZbAW2hBRYMtWX1XqcNBBCuP
Nc2vLsBhfka6TwijJfHJSoK8CyCQRcDsd7v6PQdrDpwjYdh0vq5W/tjY2FBRtPKR
cNcsH5+/sfBphKaLFnc9ueR+oNKxqaxM9e1xdX/GaH6vdE3RntKJJLMarUc/I0Zn
Vkl44pfVbIQ4aoArW75jdMYxLnlXHB1CmHHDeSS8OHz/evxtTvF6KbBOB3QYl7tk
k9+TSNbzQFAFX0bzUwcZR/+dRrGK2ftIT/URwbIuRSjheKlasSsLimOR6S8xMV41
nog/MUCamM3rH+NuGruKtJlsWRiZQJfQZrWpmzIZqRy+yFr3QE6AtRhMUh56a0FV
yO4w2awxz4wIQNR1x4tzlyRh+tfs2+jfTvi+Y5rYsIsN0gyEXOGsSMh9DL0tcasa
Ihl30amOtTrf7Qi/EY5XFEKoX9Pfz8ZITqbaJrf+6nzm56ZILykJzbFwFsovIXYF
CJQkNZACY7RIfAOFpFx/V4xW6xGiBiRH5KnDuIwmQRPieC3ufxdn5MoKS8b5/Jn9
6W1J07eiR7CuxvmNLfJrnekBO+cEmk9IyP0z4CK4Ix3TxnrGZZ/v1QmJ/JQl/Qzm
Q6j565SQ8fzX27jvwCFxuFB3cojRWBRane9qcWEZ86gxDynFidMsGAhC/4OUIJDG
bG9RLwuuuX5uOTPPSJQDNaVDG/OztYRsVn9ZYUq4nKoXe1kwX5rkAy7looN1i8NI
ixTfuysb/Eeg3K0C4Z0BNr+6pXBYw1zSHW3BSmW4rx4oUF4O2Uq+zURuKJLCU5E2
yOu8eA4ZRh4oWpU20SIpeG8zteQqPfTO8qhakU3tvqDwVjNBREz0cTEOEUGsM5f7
9Y1uF540Q4bJjo+uODHtwnezeQdcv4f+hplR8sF8hIRyUz7UlyV8EJMnIPzo/O/h
Cko4hADL3it2KoLAzZMP7Q2g4UfLoTvdv5he5kDizogDM1WYylM16474dVWyZsEU
11eapqXqJijaC5qEilyPduAYSt8hL1kWuNF8c230EtN2v17hI2v/UYfg7CiDMQMq
ffqkFrqzGPXU1BSkJhe5u8sy9mjkA/ZnqGQH1Dqf/7SWQD6kAmVIxyuir6n6iKaW
uZDjYOAQuJCh5obEvzCKUePzIgpIWM3W9NotpZqAhbMzTLrBEng6Xk+pdcp6auWU
gzt7v9EK8LRghoJscKJg5wIAkusW+ZoLtSU5Voh7hxcVtprH5FVYcLW3VVNaBAk4
maH64LdrrUoAr0X6IgoVxuWzzXc7YStNeY8g5Gelo+mjFQ3rTWBpNf3eUHya7OxO
ubWkSSONXhFC8I/ryOo5KQltsCo7mK7duI3SYLc/dJRSij4h5KwkH/p5OBUc+Lit
8RzMjYlR+iReTJdCT8CBmRvHmxHBw8l1TN2I74Odt96sHcV+jqew2/jEc7ARDGwD
2JAp0/D/zuHze3hPvvsNEYdB00YESOhkSOYpYHSj5odb4zR3grZU/GI18RDq1MQ8
CFG7gTVTegRaPRHaACvsBC1gh0nsnMe80Jxm5FjimdOrzY4tHWnCeG7N5T73wN/P
bIyJ+ztDJ0HH6HHRcMI1sYbunmKm3sUuvLk/x+0PYP0LXPBDS6512LY3YbMFkwRF
UvncwI+JesqkwBIjxRSsfTIATw8ptPB1BJ0XWMQWPowNSNreMpyZ4qZAXvKrIrcC
qeHx4ssfCH4iIF34oXKiJY1YrCkARw6RIhJ+GEMyGLFQpwyK0EQovCymf0LN4oBa
cezQGsBN24/cWFXpxE27JJIyzO3gBbEQPGXkPOWUQZZrNaDv5veEE0SZg5Q/vM6Y
a09P6o2VtbJogxDztnnE8abaZjPRYg2RnnOrcP6JPx+4DlQFexqvCnuedU+eB2M+
6w/pcB45+eBQxqfHO6UYwhlUIPfQ2sDbk4lA4Vi2Hr/xjiFeX7X4/utScJl/sg9K
MeBKjvABneNnEBnVPz76o8kg7ep4lcLZt2WGnzpCcwaEbr21x56z7WqfwlwRKEOD
j//e9PM78Ti5fhv1u2huAG8ScDJrIl4NU1jAlst4saf+tTNeOS2f65T4AARBsOVT
zQ0FKCisZlyNCrHAMZMDcwVAC49WIK5Gdix82ydfQAuDVIcA87QtqpccSquYeE7s
HH4uZPfml8wX9UM425B/vpquaFxFIa/p3etJwdfsMhdVzW1u/ligkiVdZVOLie+G
lLciy+OPRDN7F7f+tz5oWI3m/QXRoHPvi8icReZ1jVJ0SPWy72bMUiIHyQYFeaJb
ldh5pUeoebn9pksjkh1gVZvTh9vyKthKDENEDJfhTUnQyXbTFYQHqThvtTbsm7rL
zJs0lel0Szk3qm44+VxODE8LqfNCKGY8JKxNDl0Jq+WA1RgWK2D23STdgPRUi19c
dVgxhjQsLLGirDgYt+CUxGiWVWdthgTtCGqHYXsV1h3lDRgS9IgdZRsJb3Z3IlH8
5mDZMuF8nNYi4rYdqk1yXbBnUzI+tXxEL3iSizcFYuiumsr2HpREdAxRU0EKPBMZ
Ud5vnMz4llJfZzlXQqH/QV3l3sN6JBkek1q6ynvh8r/QZnmzHvvF4GLcfUPFb4nj
4eOnqh4Ggjt2N6Hql/ndU2BKgZwuTImpQaqzJH8xoDVeN7K6d2aw5NbU2AjQRae4
TztZx4RxcqumQ3EEsh2E1FlX4gi1wyKNrtgkauyUN7fEJGSmvPiQR31qt+iX+7Ij
o+7UbCdCphG/jDoE9atwMWErqkUwMI4mEMGwdmPdxGEEXai1VvlDFhmXj6rxvTsL
q5+Y5klYUfqRkhd7wtaGar1Gxw0Jw6fIq4rxO23YdZQZrxUVt6MsLKHtt+FmFww4
ymU6Q84UBw7R5cRU9w5tiyFj5ojspPEQT05wZKYX/fnC5N8Pm6YGQA7BJWMEJo8e
1fcCc1elISyO2fGrYtax2fkoYTnF5TdEgFui0UpL4n67Yhd4EuDlXLgX4BteiANy
ZAPmtC1zQaNA8PzUTWdJxDDfj24O7BRw5H1xvNsAF/YSDrwyWUr2X3G6Hu0bbM3v
2jD11GyzqOSRVd+QtC7ROQaS+Ht5S5rLZgGgqad4JS69AdooalxBu/Zm197WPpi7
sj+NOTqtsOSgfR49u2u5i6dSguYvrNpKqlC0C7j55dOEjDfmhYTSMKLGcazyBCYw
kh10IcfurIChRTvFIBFNbGq/w7p7BiitqAAXkIyCFSz2ukGuXPYKT4Khe5ooHhg2
jHF0E9qMB/4u4T3EKoaVB6Xhw8N6p8mrI7PPtr4hOG3YXAy98/zizyeZOod4aD6r
bFYTVn99D7JfyN9DpdupfgsozKGHmr5frkKBU6c4g+5GjJSDYVLlKBwU2XwWmdxt
xRUt8PNV5ExBCgbdizOOddF62YzsfQW0Zs2i0qT5GSRDvV501bpkd44HLBAUP1ff
MwH6yGcoT0glyvzFVeXRfmqpEzJFY4EvBnutUGf1D+4ui2B3AKSZ6hMVqnB0lBrO
MvlrkO3j5wjf/zXWPs18cB6NPuUCzCplv9f4Sn1ZoPIjjZLsyvnpvqwJF09z+Yx5
aybZTX0pB881vYR/iecMdPizAwroKbl7QoWyo4c+WvKL63D6vSRDbXkyvlR5qPsD
TVMyIp/t9U2UtbxV0BnG6gIVfENZkPS04SMrcpul3XWPHdZZ+PmA3ffPqg2FGhEY
Wo8lul8AbOD0vTOQFK1DGWxdvpcXZnzcxNKPbjg+DIwo93W92iEUDCpFmGgwgpeQ
iTUbSRW04IAiP7MnxzN3aOhorNeBUASdHW3D0AjHF6H430c5Y4OLniyI1SDtz0bR
LDQuIB4O+ljFKCof9fsIDLuoEjhRLeSFrhu+275i3F7DXA6QQncGUuK1C2fBMv7o
cu/urstfchmpDDXCac7C5twT8v4dWO9IpvzKMixm6EIDPBnwOi9/aqO9h4FUjNIT
Q14NaxCCDkHY5KNS4Vivi/QP1HQEwRuB5oOgh27J9d6c5rlwhP1wdTWQKwYQaWSl
6gFMLXlMN/bqnevFrqXi/j8UzIZI4z73VpNUiwUJND/VR3eAgOYUoabjfJfX9TGz
NccuJHV2NuF1lUnujKgwO4tP2xnO7WZTenSAOzEzwhtsx4kj/7F7I6avXL6OPe+R
Zfo50mGK83VK7s/iuBAQZyPbAtlPMrR9ytAexXZb3xBuMEiz2uYtFd5j8UNe4sT2
lB80DDxrlauMOQ37j0S+vEC1iUm/zMyFSDcjQercmbSCwE8FY67UsFHw4WE/nbV3
WNAbybp9kbeVpCt67szAC/SN1rjv/l9pMfEq4eRNa055du5bxy1Ge/C00UhflklM
N4kDkVmyzwYsi4fOlVgFxoSFfSMV1AFnJ1/Cv+1XP9bjVyJ12gsaQOefMpyRY2jW
Dm4zu9TyDzzgZ2PgogPQlkLwS1gM/IIU2zWuc8qczl4jfbKOmCeRY9KyWBeryWYS
ZOQ05GVJQEOdACkEWQZeUfmEkzifvy+dJMEgWZEmWwko9X7vt1E78BK/EbU5jJN6
+/MLIU9esGnEFcZiRs0PCyK7pAVRipkpEbKAxycbDPM38Pbxu+Z7QqJOTRk2nQkb
/pmE6W+nAup/qUGUY/37jitDittte1DBxXFD+fydEaiZ2UB3udWgONHuc1pFG/XT
tncSVAydRiGUpFAPRd0iVsgNCR+ufi4E0Ob7K7DqdQl9oCv+M+lAIQjIh5/Hk939
J1iqqdu/CX/FrQxPz/7VVSi4TzAlitnuKmLrAHQf85+ce5lsO7U2H+lUMyAB8mus
G76sOO00m0aMM7BjAtcLqu3HPJOUxXwWnxZehpwYBIWYIh2Y8UTobbspBKPPefdH
uq4PTvQ0Y17FptysWOlYK4zIDtHCezlC5UPR0liU/8pXuOd/GIVfR7jJDDpEPXnq
URpjYVCRZsm+noe0BTpBRh7H5PuJ5r1XMfosPAsVC9E+4AwbC9vfenenZOtZuUWG
kPscCZT1huFJE+rQfSz8avn0xA3oGaRqnyN5g6mj9vUexMwtCRbDKfPAuEgl9dF+
1alJ7M8Q6sxdZl+maFv1X1G8pN5i34muUA7oGdJXBhWcswSWY+kmf7zWLhZT2VvF
WwMCkLPRIE9XuL+SIgzwgPgK89ZalTh5dXjyyGAms2P2Uie1tZqNrIaZ83vhUoFv
/Gal/HNoP6CqwyP42Se9+m8xrEfidcjq1pk3rz8HStfrC1LhdMgerhjAGPoWNHyO
iJw5IcTqczdg8uOy5W7yGNmlhEdWBF4ObqCrsDNJiD/b8J5AkOaLCN1v5qrSZQEm
slnSXeX2GAzuP9kg5lSTpkaWtUZgaIS8IVpz10gxIgAoh7uawBYn3yfUWWo8ZIqm
rh6bdz4KqoLFm5GdwDr6eErgX0IBFbob1p+mFHeWfzjpf+wFvgz3e+3GqQvC0Jew
77+PfnOf3tgu0a97GZdjILVY+Gz/ltsNmQoXyW48Q8L06o+ykWmGzdtSi3SS8Q7F
vUzWDCy6ytevTM2sVb6ijM2JqAtz89Ugx8aVx6/rMe5T678Ilkj7pyQN0bToSh2X
p3DGxUI/5Qj+6rc7Uc/kMqu6D4apiqRK9DIjbletmOTNm5lYaXRrvgekaY/NMb4/
cObySnmF48sqZn6f+ItwtS3mu2yvjoy5p382SUuwja+bBu6LhydKu1N0dsU8FDs2
2byBiy6nApD46NDaKwMsHepHwOc9IfqsJ5BIzqkr1UqDd1yF8/lhyTU5/ajyQPyp
okkvsp8z4rmmrf+iWz3k3UGk8WiMjBRZCygWb4MxcKx93XJvO1GJ2Adgzd3K0p7c
r17rLvjPqwBy2766N9dEjCAe32PVzI5rSX93yTVpc6xq0cme41lMPw/LXc91IDnV
8wKGJyq4/44+rku3Qo/2TkYeKOwypb/2lsGV8FAUjcpJJeVVGe4dWVNi/FT1FH0P
ek0tGoPJtEfL2Nxo7ap+AFI03DYMu8/QwrkX6stJwtmcK6+quJ8ocwrf3jgoRX1o
5B+IKDCrgzazVNS9tp41Kwwy1aOBPoG6YXJoSLRWa05StfUpqRQAHLuvtAMFVhT6
hbKZQ9NNd0slk/e+5hgkiM9UPj2WKKkE7PK6x5DoLqW3am5vmZQGSk0nmx12snBH
oXvhYkGl64N/p3rqGw1hE8WWdwM9u+5zNknk0ZP1P5qhgDN6MumCgI/KwbtnLvXF
VOd7ID4/mzof1o1iz65oIp9DgIQMDw1K8YKOdRozEsRSSmgbTU5O6Bg7gcWqUDO3
Dzh8vgDwXT5BN3DIJb+iuDXowwtkJkEcq1PpM2CbImAAg++S2/pnb3L39aju3ard
H1A4kRmGVjH0SHPJTpu+fRYVUSZLBJsKlJwO0GHKPhQ/vQkVwmftc1zV3OguvUu5
QBx4CT6HdkvDYAy1zDa8RB6FKzVs3hT5FZwFzXqyho2/uOWDeKHrc9e+78+UDK7E
iMUkqNLt2K8m7zIa0gdwG+imWP0Ptfr1uCnx1fdcik7SPOrdKU3MSDf0rtjbjD8G
jni1jn/GKbiHAHJ3QewNLaP5o/EbiyDTlJDdvcRhZB4sxR66bWTutL4EgvQ7Fpei
HIAxf/dYCiw8cku3W9VAL1F9UspTMyR2dmO+xmz811eWJQUmYhuA7D8pTrqhKa3j
OjWUoDLkZQYpDhZlzgmNYOPDv9VJllGkIud9rhM/Bf/A6pSgrkXFX8C4PDiHFNyR
gJVD2yi7HUpjE8VVGD1epm4+PKhxS5y78chx06tfpPGWvglbn3ofTViqWx9usj2z
XU3ygC9ue/Q4vhzKrw5eOFSj2vJdMQ/b6G6JRi1CUQrVFXnsZhrdvtcfYofH0HlN
TJS7f2ULP4Qi7cgEZkPhzgUC6C7foSypVXhxlL1NdMPe6uwScHEfCTFyqa6palWz
t9ZBtSE442cpFu+n6a95Gnrr8EI/ggUaco2tLZsHjSPAI71EjnsT+mGdJJME9t1L
NTlSJ+ymuCyCsKbfOMIBewfn+1d2AvM7l6cLxvZtoWhHZ2E02AyyAP4Ha1mmDsIL
p8VyVSQzHiGoWmWDLHLWxltWEAJOr0QmuR7So0GV5cp+h/YyJpG1WFIXrBXaSxiH
Q7JeN7GQ1qod+qRNYT4EdJkDesb0f95F3fEcS8R+nSH2SxQvIXAzfA1HOqFMCoA/
l1KuMPXf9djcegbyYXibf14tQcXMr4m3j+M8ucSX0sntt3w3gVaxeEUInlMJL4p0
7qP8N+OJguvklGiZutDp9QT/r9jQKjmVYEEolHlZesiCl685vmyNlTFZFHNHV7eF
nZvvX9IV2VUsxzGRy6Nr0UIRqt7XRf7G5nKydw6njj4cUIIKG1DbEKNWF69XHLay
4n5hKlhB+f/appfCJKwaw6NJeeqbyb4t7ACckhilG+eSo4HAmEEduoJ+803hQQOT
jGyFqyfC9dAf7XGRuZqMBB3ucYlt3IS/glM1VYqkD8LXYPHRWXnKw8xbFgaaG2DA
hb1ZQ2HUuK5mBklkz/yu1Y9aP3+sIf2RvVJTvBnQzK0WMVfMZpdbVYmQqGzE5Fds
b9+dRWZLK1Sd41WAcN+vhoGcWFStO7OyPnmdNcdmHxL8Iy7qlunbdqjqpFaZKFbC
Oa+XvMhkEsu9Oyf20FuNG3xBpJbAKJHci5hgvuCSM7+v0wMhiuNvHicGIi90kRxe
i5KNhQ0sO4xRVjnkp+vAzW12w61VGBhBUtYFXDZ4K6lo9wHnz76ZETktZOUDtVv4
ZMOVPlNJ0XGsR0XN1Fr1rKVlOqSg2IAjl0bjsR1k2FhmFCLw14uBz6AOi2KFbxAY
dmfjnAz/HXW6C5bjoIXWCs4KW8+tdvJF6p463ZHDeIsgrUIsXaF8/Gq/CTW7EByd
42IToCAjcbHLwnpO1upSjNYAm9dtLcb8xXYgOksUJ24Re5rAFhKOFZAQv5lrTo+h
IU9zAX9o4doMFVYDFQrM5HuCqSYF3kTmcqBfQI7FQqQrklPTjrDmo8S+Mjt42J33
aQJxSpxL3v5UtcXZOXia1Nq+Z8/ovZoDNaJP8FkA/u2wXeb+Cke+rPzTf/52q8ip
YC7gkU9p/iNOQ+50hNUPXwJrB4d5qiADkNFI08G8Y9nRFKWrSGmSzKhLoV/mOrtk
2rqraPJYvgDUXQbEVIClfh1pcFlvTj3mG3ebFs+5pkcCHgUfiU/kv7rfOykMa9EZ
4QCeCyv/Hz+ks/KXpFpe3sWcofGakxfE6xO0XQ9PBaKkVV+70MCOuG333k8g5XVK
cj5z0nj2wuMl0Qte8z2bjXB/BHKGZPxiZYKaPRH6b1hCxqzMOHygipBAjbl1VIXI
EiudgQJN3to1hV/Mcz5AVtboG8CALumM7RCo8TV3o6k0VkvzbRwbGYRXk/QQvWjd
f12hFMEkRSCQ9Bk4HsvM+aSyT6qU2vEK2bfLQwky99FqMFbNMzbqV7yiwty0B+Sy
oYJ1S2EDvVhSLlmOFvIR+XV1jOg49kA8DPlepBac50DMtGEWznPLUM6nEoD5dJMQ
AexE1p+hUDH8rAtQrbws1c2Fo3xl89ZoPeF9OKIkPSnp3qWXOvJLmRQ5Orzxtlun
ruBxwys6aEOVenbWOO30hHsR9II0IdYdcX9jxvYiHJdarrhHFt3IZNP2bjQu069d
7dp9UGrfkdc1m/P/JFU4fGy9M/iWElioHJXgsq02/ShR+8/p5DhRIyj3uSlXJAGU
4Y3AduvGpD3qolvyr3T8PHpbzM4yYQBuQb+7ETrkW3FQ6ye4fhH5wmPh0oHQNrq4
NA3Ganqm4kaKoHodqV8f+NoSxopHfR6URaxA2TwwBfXHk/T7Ib6IQwCqUwDlmRhz
lE5Grmu+LhxNtZt95HXOqTMh+Ezdl9lbGHorja7p7puqmPf0/sxSfdVDYxPj/R99
wMabDEXl4Ldd0A82Pwqoa9lBclXYB/kerxaxI4u6NzjK4smshoXaH5ZU89/h63Yx
cErKvDsc4m4ZuilpyI7BDgPf1Cm72FIY3+/ymSGgttBdbUaR9inuBlgCApDp8dKl
6xVlYd4xjvYXkDAl8SuA9UOkc6n0XkFErYRTk76JPmF2KwvfSDSGo/pREZZsXwBK
UFft6aVWTMJXTCnowrgxH+GED/6kBp/Sj7kOhL3JT2fGjjMpGnXquPvdQdSyXIdf
fzUWz5mgBD8V+TXbFbKwQOt2J4VdYR3fX+UWbvdh7eMj/WIa+/pqOpN5fv+ys1js
P13zJcLwzN1Ksftttc2sDjSQoaLlZdApF2F7vbsbjaUwV2kk9pSVbsDHphgqyrZ+
iKV5L8qKkyZqiGn1aONET42NYWza66yBY8mTXTwvKGUnafrJ6iuZGqZVIyE1bGa4
LxwmXVcof0Q1ZIHjN7TIa9a+UIh+fvVfx3aEc+bL5BJH8ck8o4rX8LKom9cWOq9n
pitOPb/2HJTAm46kEstPGHoNsc+Nztzl2wIJAmaUy5yRL7yiRswoYzi87fiOmT1n
2qoEtbkUfOUXroNnoNwWUkG3PZ8KHLcSc/xqKkbLnBlquD84AZ11gO+bGwOsEnzS
vsqlvuQ4ey/gTtoM/auOZUJlUn2z1ZxUXIErlAruNV68AqjKbE7mSmh0Ke+iFF67
tTdHfg3vukZo1ZZEtMUFVdcXROGu4BJ5KF53yZFZFyxYnU8DR0c8BwnNmUTV3ZxY
xYMnYe9UkZHcvm+jwCaOnsx+SCn+WrTlQBaA8JxMQCxj10g6pjZrmH/o/8owshaE
hY2xjjBhGn+vWYbGlEkH3l4iMKj0drRX/ViFcxDLEgLgdrDG6y72TAkZouxJqXYk
Ei7FFpuvKOygVb9s8bDGFUaAsZSAh6wQoYTn6ZzNwZv1G50jpesYsuPEuOmwolEW
SkSjDUGuEHoXFAy6LsoARqVlvx61xrHlo4/AiUM6Y+zDCmftIQq5vi68PrvmHFOo
LrjsAot4Drrh+X+cJcod1pg1glOP6g13zq5um3UzLKnIRXIFxQAt/LDZPj7/deY7
XSMDvxy8+wJLJJ+9SsU7UgC/uTJBzH2t9rxhTVx83GiEXSGyjNyvWYCnfNkFT4lx
ZQFHV98gjEo8RH+mtBPi6rzfyFZe+VB7Hj+Ael1thZc+l5n6lGppRaY7YRRpedVL
w8GGmFTruI7+BWLzRsnCYRezBLvJjRQ2RrEhvAZahcNMmYsocpN5KVrv12nNMry2
ydIQWbnO5Yuzto7Gy/8zAeB/LNwz4yc+fcPwQmCtdaHbfr2jbrWDTPA1emQBYQlv
OClzhd5C76r92sn2teZn7cQLei6v6S3rPDTktrf/PL/P1bA77BpAdHja8U5zId9K
vYcPBZ0/Oc4gisI5UoF0iNzQZCfZ9M44zPm48YNvS0mJZ2dnYL9BM93aK/M09CfF
2xBL5EvsADVzBZeH/xJM44TbxZcNRdoVS754T5ZuE/xYjA7Wi54gwzvgQS7gghVH
n5tIjRZ2aF3yWGNkWmahgGY1YH8ixFHiF/HNdcCw11pGqHh4zFAYJjv/sSGG5G6N
rT0hP8qFPqLILmBZcb+p+/KD0KLLokDB+XAbkXko8eHmeCfC9b7oo3p3sIqwzZR0
ELtXiU7kAq9UlpU6nyjmlLtt32X+G6MFKh457tFesZcQ1SmWWyEZuE0hsoo4WhD2
yGjFf9DpK2Y0wBX4wc1N0nqW9hZ3rrBBeuEhA1Qj3s+LdatczKUA0B52rPWuaWwS
Ijp66DNeuoMgnBS0Xqxrg8H4SDlWa2FjyyZEFawNNfylQnqSeMe39BzroLG3hm1u
NUjVGLsEzMp/An7mcBFdiPytkV6aQ9L7Cm6Z60Mt2dueuSmNmeCPJB/01z6+IUvO
SzneeKIYHdbRQbADvFOvP9fuY8Qdu1W2HatSZO15LyJ6+KxzN4iMkebLwEfx6kNS
xC0goOmhP3nYfZd9rBpuwulYIW2LE1Kj+nwa8gI+YmSEWnzsf7gEITjZL1Rn/CgK
HVJEjIbKmbesezG3mG0FiwVtubN5NQ//iPSnFmmGVbKnVesd/pMHXjwNO7O7ZgDM
ZtXT+zMmH3tl6NUSRz9J7fN/UtgjbgRAEe3I74tCY1rzb8yi/udMyIF8/091CnNu
Ho9r6g8KkEQsBdz7juvlC0iFhiqcCMp2WpCpYYiAzgOmhBF1EBEerX2tARrXI3De
nuopDf6486Peo2AgEbF7k2ISlqqOnfUJMXYtgqSRbB8ghxo1nWRdQbmD5yebFXuc
CIR0nj3VBwYswEbIq+j59OInXxt/bDarIecHG8MPhFl2EJjvUxGhfEjBaG/3Dz1Q
/H4gmXDTzy6drjL8lzKsXZWZZWFek6zCOJKFPGstC7VbZIDppxpdwTJ3P8JW9Yr9
eHXoRTFSprkZ3RFXbi7wfBXVCw9rb2jEW7qIhtObt/6E21UdnEEx7jMFeM+9u5LC
JRcJng6GqR8z7no55/CCw/2ymN+ZV2feTom0fvLzfrQI3bZtkwvTCHhgA2VylupK
34c1h2j2DT5TZD48JnWDNo4CFcRy9KRIIXoZAdQhrfFUMVoN4dYhZ1ES9LR2KyAF
ZMV90F/Fr0wO9kGT0pqBm95gvRxXv0HdtcWjIKJ65XMrT9ONsER6t5oDC1AC2nAh
Kw6oQRZRPvME2zBMR9Imy+k4ZoSBd/tfoZo7YLljgpTmR6hE4SrV4maMuT2XXB0Z
Vrnf2h6eE3PHp1KIMnQsRWgh+hYH21eeXBbW1/hv7dEXFSI3ZanmKH+SSSMeAoWS
q/a0WpW8bMK1dOUgtsIpp0jSALKvYw3F8O7SGBUQbRnfTV+DP8gJ9xkSnu3xOB3S
eRmFutv5yxyoqpB3dyjeQL4f759wU3nWpb4GTJWOby6DCViW7faFhA5OuZGOOd80
QBvv1PgOdO2+1jYA4X6ItVt+Fa6whDsYDLEF+8yr8YsukgKrPEjxC6nbUsjNl8Ve
NYcI+X3pkw2TXhvn+ywy4GqIC3jIEs15dhg6afvINi2BtsTJuDUowE9+8UMHz4tg
zQgh9raa53zH1dNaaogK3K6Qxa2mZaAHJWa9Bo+/fODvST/SEpkkibbj5BdQwwyP
c18KlgjmwgfOUrzc7gz1Q3po9EU/bQPg2pZMeGk1W73pzY5/nv345l7Op+Z6F0Iv
StwPI+bFVCHACZovlJ4/R6Gr0LLypeOOPGYf7tMZfNPgSuaC6Wn/VaaQ/l+qZdlU
DHlUihvErF7T9Ch6BVfbggSyVz/fPBRaTc7FlLLA2smbn9NWxkut6/9EGMv3PKLe
d9SEgMuR3PRQEkfFBTJRqliR24s7xeSe3nis8aIVwuZ98X4gXulazy0ecMqrYMQe
HHa/PP2El7fqm47H1M9f3oRCa2dMpeyAc+jULymFL+pdonxV0SmjL7xW2gpO7n8B
kb29dzUoryAdMDQkwwjITaVuLSUhUeoSJkVyrakDRu3u0c3biYQR6fu0SdDId5y5
opGh0xSHXhNfrm9TS3MjX+meLNB7sqehHK3kdNH4jog/oTFgjII6q/rFba6Vg+DD
wGH9fFQNcdBFq0B2kKgUR3zGsNZWdyd5sFOonaCB1fJgT6qYMvKbIPLe0uHZ20XW
9IRUXd3Hn2cBtgDgbbgxkd68RMAk+17t/altJ8CsznwwCM9wryLmh4B/63OK6Kzs
LXZT/eFzfJ9faNG3pg4ONKSIOHe2V5d8F/CmrCL55wrERp1roTUQLOb/Hdju+R37
AvOFRr/O432uvIL6d//uCEAiD8s3QQ5eVmHReZEdC5SnyO0xRa751TOwH2ydqcrK
gaqnW2mfHV6Enwz1LXuV778bQv61Q0qAv5uMi7ji2CC/jl0/1QpOPhA+qfO3ncJV
gd/sWqRIAAuIbbi5kN7sqjVNVcnugTL88E5inCJLgnmMjReLjC4vNvOKiE4VbOBe
gpPoPWxIQjm1/P4PJu2q04OG3BGZY7XX6X/IKfnB/e8HKXVzKIJ/134wdzD+uCwQ
quzId44rSFrIb15a9ze4fBrVGdn7TiCUF2JguwdukEM6TT1jQzDjjVswI/YOM+Qi
N74q1jdzkbPwLVvHb3RBD7EzP97bs5zdAQiE9e5es4+t/YqifykM68Qe0gSnX4on
ShqLL9+lc80KjmWmEzj/rlg8MiymWgLdGs6LcA6X5EL9cektVhb0iICDqrEaOjXH
HGEORlfUXcVFm6t4Dx93xlehL0irKHmSdiyz0VMV1bV+u7i6KfOb2tFLP1+EAMv5
4MKqlMZ2XsfAi3E5X2DhJNXqP4E5ZqFve9TYrSPQUzpcoBfl8S/bBYGcYu0sCDvf
t3sfZzfNjYRnR4vaj/rUbsYiwZe5Hw7scfKLLAqHXQ0ECUJbtcodIX9AZsZWm78b
jVxZ7y4FM5TyZJLvlxFkrDh0kjjZaHNZ7AEznnhE/2/j6EHoz+nJ0QWtON/Ebjn8
/RJDajcrgcd2tD/C03V1XLw7fnFK9u/ihisN2tdj3uhgqRorxKD7JQVVv3u4lWrB
B0WWBo+jIIKwboET0tDp8P1A1mu7KyiODX7xTmgvb6nMAcuxdg5Px2txctNo4h0Q
5EoOU/Wsf8aIPwXpjBmUmGJcOXFLLmmToOruTmViEd/nUGNe5HuA86ogZ+3W2jcA
SFKpcRpWGdHfbvVdcJ9d92v6rS0RwddPDYH9+Sd+iINCaZNW4NWNor60DFUk1o0k
UmX/hSaBucgjBlAUej/FHrGLoXURxaC/10sW8MyoofcES0Mu+ymFJReneNfOkqvH
jbuJ2CCK6p/Jv6XQuzpPzseo2IBexeYF7vTdCqTHEVGU7jopseNyLDQmIK9uUOly
9dhr/sRtpXfHaltouOMzuA6/aBCT77gF9bJ8/L1KFU5rVOnP15tv0p7nPwBrNpU2
HzuZGWA89Lpp4cqaGlYYI0pMNiZH5SxseQJB1gTHqEzktCJyEZ56shQ1mfVLC/Hu
C0Z4RPfvBtCF83B4cP6a7ctQcIVIR3j89FOTsvVmh4OG/9yF5Mthkqx62DX4GmYT
kyhkgwDte3Lw2grAyCGuYVmOkaxFiEa9+csXkmhoHSxjyAOSt323e5Edt4yzxVMn
X2SAO/LU4dFPSn6IQ2JY+gs8Pz7b097SX0ZHKiQxKYJpTaFV306gRLy1mUgXsHFf
39G3HyV+auC0WWxazfgVCGeDNEyc5Cykf9t6RNqGhlHeti0SgSMyK1aCD4aBvA5W
WoDQYaO3OE3Gf3KgV9k87uNf/HH7/5bNAHlBLK+/CbyGhmp4OKNmTvgAyTFd3+Q3
Dm6khuwm8pcWZ0sNLvSxMiPWisHn4qbC4vr4fjkL0q8rWuDEAFQJ7iBiADQjTd+D
eb//iVXmwuDSc1rk9iLP9pel1trF4I9NmMzD0BzG7DcUzngdWFnCZ6CkKo99iTAF
JBRcgYyjLuyUr2bSc1mNABFFo3DpcmQQlEyFZdYq9a4QZnG2TNHzTa9QR3DLEPzi
neOIy4TCwkNvYTs9PqIHdkveL6YHD11C3fcR2JBjIccrDNoyA2M21VXOiMHOppgp
JUzv13+ifYDWXuA/v+/tuBXZTdp10Bzqi8Z8d/aGq5hXi/DuhR6gHkZCkcn0LVyQ
VrorEL7o5Oveq9MtboLNVfeg4JSH9FQ5KE0FBDEQQG6SzSDV2Zk2QMONuf6z4MgW
vq9AVAQzXPp/xFnW0KM4d5ihxHq2+xlY/tXFNHn8kRfbT19vjJ9yjUqykcmMqV4S
1x7jwlQDb/SIAJTbYKU8OipgX0TUi86qvXDooPaeU0mte7sQ9nmc9n9PKK5iwwbm
BJCmarUmFTAUyH6dIx6aeYuZzya5hyQQ8KZ66Z12rAvOJuWiBz630XfCWVdsi3CY
LfpMiJrYmGmz0lPtX27YX0UMjuS8fdM+Bp1DYEP6xaXiD0HKGMFJQmwyVDb1iCuS
Uo0VGN+EYhKC5SoBjHfHQ8YrTG1Wt4igTVWRwYDncZaIUjAd7HIRNPmkKLD/+OKO
cCpFdDH/ss4REpIZV9evRxWsKWK9JeuOmOirg5Sqp1NF1+g05bYNVFwsFVBBhwI2
qi3Mp2W2UO5BOUE0HSmakgOAiUC+2WnX+4vrybIWcetzme4dOdfoPscwXS4igL5t
IeasX2/xjSw1XZGqkg3xk5NXATCkCR95Omd2xn89xyxpKx1E4ttm9Gc7tkTYPTDL
cUZ9hVxbIQkGf4mZ5AHwbj8c6RPOZ1Cztg6R0hMWDUcCrNGDxZQ0UIlpTzFj6UE9
ACx0OEGXBW8DBUW+pfTo6bTeYoW3NthpH36gyCZNCbk4lh4/f9biNXbAjGCawzdW
pMMu2Wnw4lyjeuN9zEfCmJdZRAzxc0Q+w8FemjDGQQnLRP/GjzV9VQf8DGeLEt2c
QFfenmibIVPLGC0QtTkBNQ5yUROZIoAtJL/B4oPzyyYipngC4pH2vNEzwo0lRwtP
mKdQEgLae7o9I1mTC7wXzijAbdEFN1gzaincL1osJzIsUJUeNaFeiyEBXzSP0MwH
jo8OMGn1pB2PstgtifgTIXJyhFlyv4ykGYyoFnJmwnM7Ysd4VJ7P4spHAIV9M9Ku
8eXVFARO9TbK5f4BafC/PzcyOEbsi104U1nmtkK2T/LRrNuIY8vWMX3sm3LQFNPe
mc/vidfONJK/qC+jJST9ePL6wmpVbwqPGToR24A9bIUQLh5zghdbRzgDJIj0k5iC
Cl7gMYmM99/OP/foIhNAhzAE4m3U7b7P2xirhz0A7U7htMuNO9EY4hqgBrlUcWeJ
tVOXS7yDg4zcJgf3D0vWegY8/znoW6rg+zJwp/jkMkQC4JQyrJqXkvakfssMceoS
1z1Rx1q55Mp9UqLRKj84IbRZjvHPiNUsJ0TdfK1U7Y4GY8ngBOOXNeyvX88Tdp+l
VwUVL1lZ9v+2/zRqLqz7NFxE0Qme0tcskRIAwEk80CCFhCVNaYoMgR8hnxvP5I9B
ByxrcmySJh1rlV3TqXkr1FFC5xj/dVaqE193CkDWpW11xtI5/zFhmyRUkXMHvRRo
6/1+9KQPcwTHE1Zw7V0AIFZb9R0wqZBsgs9z60k2AkdJaiWIijPdG8Qa4kKbPyML
dCsEfqDRVQ2NdEkvlBRzRhpU0Tul9nFyk3jBedPbMzGzkNnbLi79CeMf33JjrZ3y
03UX2wm9pzv7s86Y6h2GCmsF2Y8aeQOlf0pRUkYe780K5XE0MRmpqe5rHDDcQ8vx
HUJSCF+a35/Oo6OpYtFOhwB9DIL5mlBn2PtPMWR4se1dFXLVyWyoVVmrlNaDEleb
wSF4kFJtetGcI/JRVRRApJNWGf45EJfdoIwtFt6NZgwiR3T3/oBLHDhkPc5Mf0z0
L8UoXBpifyhDR5aR4r/GluLEsB2ueVL8cB3lf2Fj/JddUn77dK/GNLHEssQgcyaW
YS2HQbtCfIR6pIdCs6iRGNKkO+T/sT1jtBQDs/oFBTyaMOpw4yF1ViW7hAdemDjv
m+j8Z8YLa3KYS43dDIyal40jxindF1tX01Oyo2PIgFeTfg1WQtK7IJn17xbHq1Dw
J5N1JKaWjNJBHveLQ4y7GX5ExsUKcyh1dUy58mCyvEZGd8nwuXq/+WRJUaGhCnWV
HQcn/6Oj4m0S4tugTma7iXmLZ/D83w5Yuw8Q7N2TwfUzud0wMiWJGkdhsRffzoeY
n0Fjbw9OSR9LRgaZiFIMLe7XNh+2WCsRRqmPlVkSoVVuhrWJaSFcGU6YqCfsnkJb
0npQ5OjgLVANF/Rt4doDWdOAICAHHSfU/NJSX5yqGBqHql8iEFgMT+1SYcQQVdlP
nNAAsVTbuFEObxd/l4vAPESVK3v9qEN1ubhzCOyx5B2DDqHa9fe1u/M4xH7lPSTw
64ei76MJ90oNjOUCFLmmAM6+PC/QOy2cn2hH+DUIsVNdlDSxT/7Ow/nkx43F5QMd
Iw7V1n36iKS02yT8W+0fbT3nnZI8sPOD8mW5W/ZuCZGehF1P35JdIv75bGJV4OiL
JLslQnDnaR5LXhW2wBN1AUCnmZJ6//xYJ3vig/iqBTjRNFzMaUADedysJGB2BiEO
nYWvLHynu7ApjNSualR9FzIqkLmT1CMEC7tsEk0ELjSf+XZMVyTtM6ANre9FaQNq
AExpqdAUB2Q5jdpzUvuEscxuM6J4kwwV+pkmpp12k3vyguKlOsggSHcPpPofdHrT
NnAwn0QgWwOHL0JHkLn92pXTtxq2crqVwOKPztUDNVfKJqCv/JS1pPqqnIRq2H52
0ooOy/GeXDcvG2PcF9btIChoVZBtzy5jhyWbz6sRbm9ESikZbT06af/GuET6RRVn
DtqaG9l1v1SKoYAwcX0FIktOijEP63F9fPhCIBHFBS/BfRybc6pYwFuFosnR2pQe
QR+Tn5eynuDixHzIIWbd3Mko0vGnZ19BT+ybiRvIPypaHZ+/sMIuQemlW5ytc7yX
RyhAZddzGAqc7PxVIglwjPKycWaevO78Qt/yu3zuX7kYyW9vMfGCJP9ZnpQCffTD
BM6GMFiyw0dnqj5XCtCNNtiVF+6vTPZrZ2hqDI5Nb3f31zRuaStOGE9SLpWxxv1O
P2Gw1J/kUSX0uDonghT+q503i7CwkHnHHA82XgtnAJiTUoIY50LRLvciQ+7FL9MJ
AcwLtW/UYycvsr4vbQu60OLGioxnHe+vl/e4+5ncs9Wm9mIcGzMaRxoQeGfkIew3
0KeJeqqoFlB+YrXyULtD0eIk0fKsmq/fAAljzxBHB2rSEke9EgLdIAHHOdB1h2hY
s56XT5bv6ivIFZ6t/xps6qLRJ6pkyjH2pFJpaqMhFS1U7pbsGZ3NALQrh6CmnGYd
3wkp477L3/fe3MYDh42IGHzw4D8UZH+qYTO2txy5rvrPorrSD+LnvoGhgxRfCQ6P
Oo8ZPpxEGYHwZ1Xmf0wmnSrtLsv5oEjDNEz+BlcQXJKNrRZg0X0oEx6dRYRtkeHM
VHYkhMEs3TyD5cmtyv4/tUABSrQ+ytCGfAtTEr7dypPxLHhs17/7AsIShsjOuZwt
k0gcM30lOz+ut211LuASnDb6xdmx31NFrbjMrzS/wySRqD7I43NY4amcUGIhYoDw
02K62A+q1G+GJjo1zizd6wm2apYKOGu6B3KVCF56qVz7F07bG5lm9PRH1Ec+vVu3
FTGQbLNmfCbUVaWDfRWgaq+UwEtPyKXaw2CEOp6bqv9JSRvo4rUN1gLuuHhk+lN/
uIoln3OHrQkvcgz0zjjkCdvii1ZSfMrBS7uoen+o+pcHEUIepkDwxSQHW/Mr1rPY
0neDbFw8jv6yJP0JafRcCWDspZKUCizw2YXseeUVEhJJ9TTi2XEj4dEJxqI8fXOr
18er1BD4XRDyK2qgvA3t6DtstALkP0tzLFBZY0+8GPaJrrDFbp/vpOlamq8swUq4
j6cIvUVCwQkk/Fguggohp8WcZ8RVE+7s4h6JyP9/Ly+dF//mQdzufB4VDr/cEp7A
LOJlOd4waCCnyl1r/aDtkBRpN6TjpZqhdkTYxqta4KZiJvnquWbpI6Rr7UH6JOFP
Xs6KHdsVTWfr0DUb+JF3Z3ouxxu0c7rUNR8XFMkvlGnJXNhJt3Q9ajowoa6CtFlN
YeY07CyzIONLkVvSd3wNq2Oo94QYDsGT8QGHfwgtMJ6dSO/zI3MayuKa2+Rjtqya
LsBv2prt2zWRp2nbcW3r5Em3Bk5IyJUEcipqJNgUM9Xoyty+uzCkMCyM/2bwS/Vb
JqOxb+MTNZ0TZbWtkA9+b4YoP9277e1RHImGmRvwENbKg49sTSeW1sFHIeqay8Cl
RV0KMY4ylKR4ufiH/3EXOoP1CAUlArKXKtmZoik6PauIC1OHzaQBQQYdoMclvOdg
S6WA/cIV5XJGd6N31OJJWO9ixROB9O79B4SnuOoL9RtlZMB5ERuZzTvd2zxXgI7x
Ka7r3Ml7TPdafRA8t7FgJEvxl0hrWkyeiQUSc89JNmwU3Wb8D3z8mGxW9E7jpewd
zGzWfqmIb1kRpBC1Dj/IKSgVRtUr5m7Lj/PdgmJDCbUavKndb0+xp2fzrdn+hnKi
2oZ1OMGq2NsphNsR67nS3K3FeCcL9zxhFR9/mgOBj33RIDdPpeLIMXfopx8GgfbN
SBMSPMrByV5qgfBknMNmxRRi4guey25gvjo6hkrQs4J1/PFgmLa/E8YRGYq4j2Ud
f6Jij2wD5qv84ZZZJs8KX/Bzv6pUJkDbaqoSsItpXDYw2VchsUU/Uj7GRYecT9m7
gwQNvkwlqOe7ofAQTcYVStNMFqGxE1ISQ3DYV7PRAXBKh6fT15WDNefxZGWbFyUM
CcKCesRUiBV0xp8Kehdl5BR1hL8EdJgYGIHLBSOmBEdLyGoFS/Gjh4eOQnwe/a/y
CJkb+Klo91l7AlNplw2ZzR9CCxOl/yHl7HEmCgTahVnzXc6cPlYUjr4F+6fcxNmA
TRz11e1RwivvA1Gfoqfdwii/V8A/3v1KTOopv88Rp+/MJiCvL8LGM2a5QhDLvx2x
2LyrboAAPh1iS31PWNeEiiXPH1XyngNzFaAMK/Xyk8O4xl0D8NJXHYxGvjtqInA6
2zSiO9yOL97i+mTUWXj/83+4uhI34yXfoGzumlAmzIl18k046mxnq8fo/YnDStwh
S8nF9xmu7U51NSGgrV+iwkY5TmWVECDzoVsLIqUVnZUGpzCXFsvTciO8Evbrs051
TprngoT0sAZXzV9Lpp+9+cOJNhzAN709QjCIGTD2JnxAWG5OZN9n2prZJQIXmfP9
v3SEdKjutsgEIQzxE3cVlLSwwry+VN8mGwvbMgRR/QD6KenY2IJS900edWFbndj+
d/hPtrcoc727fP7YnopNT+0PepUh7vGVFP3zjeF+o60haWbP/B58f0wV/us0DsRB
4Yr9yRkBGnnXbjYnRH6cedcz2WbZru7PB2ezIUCZ0tg3vq02db04M97uIYIvmpXO
j3AksT/o/M3ZYQyo/SaEWmq11x0kQyZllYqwrAnpzmrtosuLX7AmTRP03s3NLXLC
u7belj3WLJWtGqwtzQYRlI4N8PPIYkHs3HQxc/rson7sKk/m+wPbGhG1GIt77/rv
0hN+Jxtm8sRzqdSkWGkQckHjYFFNWJv+p+u5WJ0GgIJiS6Dc6jigRYiOw3iPyiLt
QyQVqOkzZAczseT0OIsuhjrfC88pYY+K6Snubf3FA1dcnt3/synoUCNZkszjIe6C
pRePMheVC4LT88pTqkug4TSee5G8drtNRUx//LXsZO/527iMQzmmJhdYhOlONsTq
CcDySAu0hAAyjnavRCsEYXgORINTH9GTp5C4reFuEz+czGYx0uExaci6jpnPt4WO
p7/GpkSIdzLUY/5J1bMgxbO6hRC8bveMWSlNPMj00sBhNutb4yKdBXF1pfhpQGut
jqqnFUc+2rhwxWdTNcaSkQ2hOOC7YEjNyTFRa6rh3q3DPX48rVooRxsruSkq/4DL
MlxmvpGdJ/s11wQKr/s/uA2QsgiCFs0ROOvwldpJLuC+q1WIeJfR9WoZg1wmkmqq
o1KstQewE290HlU6peZGIRI1fUgtxOBU9D3GzQS84S77xL5dmKZDDDnxbqzyYtf8
7HIIUkjcJ7S29DxJ5ApKCeKTXmPlbnab1+TZyIGS1c1EXmtKISSIXkzT3ReL5bGd
o/IO4pqEpbZSmKJXfXSYs5xFkmjtEkw6DrTU3HIr6nupDn5fZm53VIQ7oAvPhAzy
V8etByqwFSDa2iAK7Nw6KQKG4lijktAZCzaTDxY3ZCG8b2BroHxHdhN5JRZdFTFA
h2pEJP22brWOgoYrjZU5d6Pcz/8bzwkvNf8wyGyfbYqWmO2iwZQvuqmed4aPeaaw
NR8IMcin1BXqJNs2Oa8tzo/+BaVuGs/+JLP2/jhxMb9BhKgSyRoStZu9vXfwgd9M
jqpjUVAPF24AEM6/gWGfxXYEYqAL9z43s4JOfETNZEviLmGs415iwkum3Z+nOvt2
lDd4L6QpXlXJYhfTgdeYeUD7eTSp2Zoaau5Aq1HdxWeB49zYs3duJZAuaNC3B6Gi
CBM7sY8rx7chNUM8wX8Gjkb14OFSww6UDqyCYGliZJ5Io/a7dKwPH3I9eN+PyStz
p7feUyDltZDFmJXYXF+DaOkivpBAMUTBz5G2CtW0QoSonP2nYlYT7pPm3RDxuP56
jx65f028PjbsdmCSWi7P3GdNw9nQiFpWBAxRC863TANvMfCRvEoD156fxQGeeWgU
wZ+qJ8IExp4MSy2TsnBTYLokTyineROdIGV4UAB7TZOLLnlqPaxZmi/MpoQ5IMpR
2EUWUAnmNvDJKMYvC8bI4utrojn6lDEZnpQ9N0WpI8NfGVbA/iuHjyx4yIDVrPEP
3cL2te58SDDrmEO2IyjyTJKMjk97ZUOqvojrl75zgEei0s1dTqUvbxchHlUDxl+W
813MzQPHRsZD91S+7YPFnANlc4XvM2Fw+1py0mTU1go2Mtw1l4A9bLur4I2Dzjf+
eCYr6oS3w4qa6/7Tzi8XXcyjDfgz/qA/QVIi0DXsKd3jEIlOaHjy8BjOEtW0MRGe
GAHx7HOToRR4t+oyFd9Va0+/f8frwLb0lbpflCAXCjt26WUApijgLbae38W2tW6h
u8sd4p8fr0YwBvipveAhI6QZwLh4fAnaSNF7SZoB0caDKUBS0Lib9gDaNUsUyPRD
9Tb8eBw33X0HrgAH/fuoBvT6eFbqJHi7RcwsX7TCU1pyaZQWpaTDoMBmA7QPL3ry
t9rHj8LpUCuHOoDzTQj6eSarMYinw08dIokYBsNqkpEs+sto/je7kRtcndXQzpM0
Uj/imVDCgRHVYnzdD02GzcM+kNTRxUkHP4DM7gJLpYzYhkS9djwxAcr1fuYYFynw
65mjy1OqS+f3Kn7CYOIeJqL5QNfK4PeebrdYVHGXcklPjJ4bXpKzjYlRdZkXgU0b
HOuWO7WRZ8Ewx8xcWYaK1LrqYij5ijC4FuhmjVcEqrN71GOhrb5KIQptUqvbpewx
f0/dY25V4YeWEkmEOUHhCleQQJ2nnDmg6vG39TyNrJ+YRn37fjdoRgS/Ig1FN1ov
8MRCzOPFgTFi25eK5b4r1/BQ+EQtraBK4iVlWE9FBQM2NfAUSKKAUbFoM8aWAQzK
QTb6DfgvtxtskFQzyNfNkbwIEj0L2w8O9e2PTQ+8T6BQFQhzy4iwySe16RSK+bzL
p0ONGojVFmMBc3SJ3ptwsn2Y0ACsJvc5tfRogjjZhbC22ChbBI1AyI0mvhxPtPB5
28yZPfhhEvXW57JRXqCakTnZsTleG/pu9RIpX3DeZMlMupbZbOUVk4uQj/YQQNP0
duIbLprn9s5/gCiBiJ4nSrsEvYJzGnQYFNavs94+G2WCsr5cd9dJHo7pgkEpXQqK
Kji3EXpa8XYwjZEnqCbyrDoh0OeNGj4IJEGAJ7MN4nbGErgYSvWLqQv2F+gr/LAV
Ud5kwYzIUwExhGla6E2HOb1o96fPWWInIggHuSr7G5fPxkgVp407o72WjweFZsIW
C+BPbXRyq3U4eMczMOWV6SHftXMlLTXFKnmQTlRUw417fxBb6bz9cuM5oCFJDI+9
6Q2wGyCdQk1R8fEUYujwr6WsRpA7arZXBv0O+lSgfHxwzW4wKb6TkG7gqaSz9iIU
QacuSSPhL5H5i/T1A1nWQWZkckdnnfF4xAIwxcufr4/2Cdj4UBZRsQRDCXoR5NVN
Yyb4ulpTU21AxRsdMtxycAkPX7Gov+nPxQM2W81k+Kx3SOVxtBb8y6I3izhIzpEY
JrPB4OD6Zjcacc7cQc/1/EWEMmb23DKrRHwWj/y5gashIAO6qnYhnDZNjTC7j7rL
0kiC6MzErgEiwR0pJbnH+wYHr8Gm7ye5RUFwv1rHx+c8/8/HrvMBW4QoWuFFPSEG
HAZTS7wHl86DRbCFTbqSE3w6y2pgLIk6w6GYaS2WKLW/P0LG3Q38A65jW1ifwTio
pGKukzoJxx/pWwCSpZ/iC0aUsotoRUU79H/6yFLHD4FxWh8LqSVMObAcJbN74nZX
t161QbqRVSAIDbncqTXbM4dwmSygt3hlTpP9bERIB9pRDdoNqAhpNjuTK+7cOYxd
1NnCcWR5RyqcALt5C3i94YIrE9UqGPFY5EOXyOBr3prNN4XXVChiXaaO46M/eNrM
BMtIFgmSuq5mT2xyrFQ3tNAWw6TQZ9/qxGF5w7aFRAjFCYJmbCECXxRmwAsOrajK
hLLTjPzy4bNFn6Ppn93/CCvj9/o//UTRhkZcfsfVf9KdixAWZyBE8EAiFtOEBbTR
s7o65MSbz2RuExlQO41RomWvvQypna8mkuZPTDxL/3gKtgYkfOax7xKmF1+FT33a
rZZCAbQpao4X80YGCBkqUlSpeIYoBLlkPgNtsz64NNQJjpcsEjRsLG4MhbllBYhD
KkvgSmL+728oR/T7O3dU2csA8XAiv0hI27FoN5VKqj6li/YaYxDgMnSyU3h0M6EB
LxjkhjAxTZmeB5xftTwVn8/+S6ct9baLIIDhR9O/f9nYO6uuFPY6t28sEFLPbYDl
nio3RY/QN/yxBO/e1qMoRkBsGxkSY734ZhVFFCteG7hobVbvugaXHEBUIvbB+29V
sa181ddOJc58rx8wRT0nqXytDcyoRQklTfqLu7uG5T8Y1wUND8kH1YPDC4PSX5HS
7not88aoaC/nsEozo8ilOlI2pZVWbZi5NgeOQQ5Pk6r0KRgrdKuVXUvGGr9JkZC+
ny4U7ZOTM8thTkIBOehbE75+/K/QAzGBnvvJSNe8HZv+MYdlo5obfm3Zn53PuuSp
7lDmbKQbg1snN4w1MM6d1zjYP3e2iiSOAVDRi7z0sFQx7qAoDcr9lZOitjzT2PnS
yWKqKZMkYLnvAs7KZlcrEKCCC+RgiogEUJG3da3JVIkwjxMAy4lmRwrt1dPv9NWI
GvYUdV/9IcLDPgqRf27uXSivZDxPg3PNR6/oGdxn+kxYjWso6XLx1C5GMhdvOzb0
aiLI7SW6AYkfJN4F1tRWgdlYncGXmq668oWn8kZcamMIC8W+3pp/wL9oEOJXjRJR
ARKWPPXEvskDIZPaKUOOF0sHXlgb3zUEUxFXvmKCUTgrYMA6k69rsaQHccH6ScPC
6ZVX4EArjyox0SuvI5Bm0+YjFOt+YYhxX4eHt4IWyUXdEEUxDLoFnZUb2+NviLCs
I9dY//zgtdLds2w8qYBr9OSPWgn6ZZi1wqGzJ7MSuZt44UIYZx9Z8359K9oL782M
FC/peBPTX9SjJ372Y4SRZkg6FNF3cADUMV865aCplrvrzhuXdDIAzS0/DAq0ruPm
NF6tVl2Nh3UJmCV03m4eCwY5BlPMTYqO524iemt1KjY21wpjgQpI2c5KueO9tlmj
6/tSRBsqFqklfnvF05rWXWPwwtORrqcuDt8d3380DtxKVpny0yPgPAr1P+uHKvTH
VwSeMTp8qjlX4bP1242lUJAlOO6gS/ln/FOPlX7tbIxQEkrFJy1RCdUF3mqDvkP9
35ewCswi9e+6Fj6aZ34cMBxq+7MbRL/KWUqrYOg9v82gSRlgUX+s0+VQVWQgqJfQ
+npcILXKC/5toaOZl1cyGlGDiiIPAayCmtxSuo1YIpOogBAVdTiTcIDKX3SR5hOk
EwKDwfZHWDlmXdbAsN8D6aoCcnkwCDbC+QwLsLUjcw3uP/TXIRf3PqFK9jNgQtdt
lWvsGd28ucha9o9lKVqwY2SbhHoVda2+JzcEDA0sQqJVJjp5v7yY7MUZpbYTIb1R
o5vBwD0bg7AA+O1bNOG2meBuO5WtA88697FVfKsrdf+flGSqmakgOO1PvoncgZfh
3fB6JJJrcp01Qk/k/IujReU8rXEZDBgWwRp9YUrWBkzHnqj91dAu9PoyqnrenNjw
khmM9ES1tlUZyJPOQAwjL84DXHVfR6T+8Wha3BRktWz977I0lez7lC8Q6htAbDzY
CAQ4qux/8PBskfZXPk7MwSbj6unuY+OiH/B5ienqWQOYYdWp6XmX4AVchm5882p5
TAibqjqJcIjqUDek1glWcm9hPyLu84TEHuB9oNhS4MZNr3sdW06yAEbkyDjBilIv
/3403AVjYcitN6a1RYXWq53koAwX2o9eHp0cMTFt4c8WI+MT6ctXnYeNQDl8OCvA
JhjVXR2avZ0o1iwZmrJ8CMQ0RXPmTxXS9e22hAw3u6iCCF0TwBBJmWkocc0odzdg
HPoB7VhNidVJuFw0mTKh8I7emMYDTg+M7Q0OhoYnjL6ASXtUOrfckLYojOu6JVes
XlQ7tuwvTJE4WvgByEDsLN8IhXOXSh2vnRIKNiZgpgyQwNt63FP+cFM8d8WsFxvB
x8hbzSyTYwWiHtx0Kdrx5nDEfXyh+/bUNAxPcYuO/y4hX8QVv3cgGLKLH/Ali+gl
JqQDglQDudHX1V02aMLyMpk6waQA0GwsSkc1agIXvgTYVQovxiFIYj5GA0jWlTfH
Zl5jeyxAnzaHjmpKt/aAxBfmRvjnvjDOIosNZ0UFDNN2Sd+fzZ5RpYuCxFRwRHyD
svZajqS+0hMj8h+r+5Qt1OoR+Ww8dK7Ib5ZR2yLobxplHK7SueWHOIGYW59DjPLr
ABEpRVBhBITdrPmicLyCJblS9OCDtRs5EEVMqfwIdYcxisHp2DWzCB7BCRa81NpB
I2OH1mS2u4MmsbUF8K3b0rSWe6OT9KzJ6k1DoWgly4DNXLe3DUL6X3un61z58vWX
iGDNXqFc+cNO91KSx8uGcEskozQZAdt/500a+lvXjIDqsdf4LY/WxE7817IrY/vP
KlVWDWyB2/NiEIkUNRizmPMN/3nsf+I2SXieQgOcXCpOpExHuT7UldJosGtTOV8s
rq6WFSC5GvLouw5zxg1jRAPbRgXzE+/ZfTc2GfAILbsujzVDgtFMiAY0Z2kPTUJ+
1UFTUCkXw6vs4AjW16To3RJFX5h0oukj/mY/8bY355RJGYqB4rf3lz9SDpP8jBEY
KH4Xtj008yvjnI7nodYRu7reYMTfBLDCjuzzIhG0Ew8qHfz5tW5nwoqqdqpSD8mj
8DzAqhE98OyIBLEfs0LvQMxD3Zl0Eq8bQvXqRudEy3VbnNrJOyCvXkPxq29iBmnY
pMMdhI9yOKJg+L/HvpSdzTpMSeUkKw/RA26tn5CAsUVIBdgA8CbtCx76QJfr9bQ9
Wve9BLaoT9J1xxshsWCUiMiBn24hEVY3tCQsEj14HHCEVuV2RwIeYhsuohH+wQ50
PwDTWC8DNRLNmGPXy2fVmI34TT9TWRG/UcPvUTaMfQ5fQruzCqnQAm3pzobGdbMS
SWDXToCx8wVUSn2DU0+1yn6KrOqu7tOlHsVI4fG9S6VNHO/2OL2R+/pGNkrdSRja
xTmG9tB/R/arZoKXKv6nMtYK32e2miSAR1vb5nh53Ub4mHovQTffpbBetX1gVQDj
sWoCEmAE+Qj/3Zqo1LdHEEPfRTrBg2hbLn9xOkmOQjxDFPKOFuXHnTuNg0gY4uJM
V32HXm1u2Utz15d4wfQIQ5uL/d/jDnRlEzK0Afno5xVZZLsFIEjDbGxE94YlROHs
WTEsfKCPTUAM75cxaEuJ3IJrcj6LJDYVKM4g+T7SFTUgQb8IQyuo+HGmsphf8pz7
2GYIqtdtT5gsnV1xRVpes0672jYYKg/sNTKjFj8beEmGjSQr7zmBvOV+Okiuy+Qw
taLLpmp78JynE79RmiTEdK5zTnLphrErZGA8cbuF1wLVFQ0UZHvjHxAPg7lgA993
IsnLv+eQgFkMgn6nsY3Jzgr/kyoP6pXZd25PVpenSBSdeC/MFeDQXLnY0cY9/791
i9eADjUDcznrg2UjBUdgLuYUh08GQsjQT6Rkpceyp/Fu2w3f2Mb+v1f8n+VfLaKB
jYosj3Ymi6vc643lQXrulPnMjpter8EqlDYd5G9QzuO4+Og0ZIDcBF+9LN7sdena
2VlCYQNvgn9z5D3BlzVL9eQUXXTjusVMHir6nkzWkjs15VRxqR3HYf7ZRqUVv+hZ
kz+Mwy13oQb/h96yRVWJqmXvxaLo/ZscioONSdcWm75drs8IDSnjSbKREHnpmbm6
O6MhRJTdXPdCoyo1HxMMkS9Nz7WHVQ3cNGnmZ0IBxnPQo8FojLfOPVs+AWreygk4
+fk6qBfgelLIFiA2sqeofFXJYhw4CF3X2i2xp8OEgOt4wWwWHUDKEL8BjrOPO1SO
c6JIu8PkUY9wHGHDvxr5/WKm+Sfzb7iqDZRf0c+4Xj9O+TKOGpRwT/ssfK7PF4H9
zhbOT9WuXJDqJCLdQ6VhuLMSK+9jmB88n4x27qTTc3xL4n/WFrXiQFLonZ2gVBBV
bUy7DN3Irczb30pWxmRG8ntmTbw96ntPNF47bnQy0ZasoZHNEc1mBOvlAPd/urva
BjowSdqI4S1z6jUF6aOHy5nNIXHwkWBtxlRLhuKI4nS7li66YNlQATSVN6MCEo3f
vGzJ1QI8VjoDqvqFCENZCBItGf23sGEU5qVSUdDg/FlIyBM5KQMdd/8Hvu7hyrlz
0tvHfSh2efVibdSZNGAHEvVYPHiohoxgj6PlSKfKbSfRU6/mHcMFqYCNdOsVfRwF
eN7mjGFbD4AlvrP91hWsP60mD72OvN1x50LP7oVnsc+jk036nK6mh0LkNjwsDFq/
X7iqOX9cJY8RRGIH9u/Y9uldX1nNaVHfhQthCCijfyxLkpTAlE2SKdKbDhlBUKbM
lCDN1sFtHoLUnWTVegkmFAA1AhkLUhp79E+STLQisF3KwD0biM38KgyGGN/LlJoC
bl5Jwt2VAQcEnGwPQNMSoAYrBvt1CyZrjXOc8eKaacgtCMJCvDPfs9Iufm/4EuGG
ng7xwYG8tmsbQ7EjP4vlZnepDX9CglNenoJC5tUXJS488uGddI06QXbHAP6z/ju3
IpJ7+xpBPcTh6XQMh7hLcyAjN58M3qi3HOes0Er0WbNMovok5yJNcHQq54ma5aP5
YXhrdy5NgYzAog/m8KtGktFpD4ZrQZHUkS5pRyBD7flzNbTik8cZjtMExxZJCVNI
nqZIxYIoq2jcyuY8aR3obD2LitN0cG2GQwvz3NvJDEkwvrcitfDyEOxNM1XAASRg
fCHKeJ63ttYtDbHgqKNBrHnUyM3MM9Kew21n9EE4AWleA4neNr6K0LTdDAsqtDy/
iLCVUcGxOGyAh2JtyYAn4XMKKK75H6aIHlI1YJ4F3K0+5eQ2m4jd2sskAfvxUwH6
V0RwDk+B6EP/5Fu94W4GzrMivMN4jMTUMWHwvZypvvORbPK8tjJ7DrD7gUoOLxZB
VzPSPPiOhcxdyQ4jgtxk2C/Y1WqtkzG8rz662syj2I/WEXPXENZw/m9O+LL6lL0k
IyACNGX76/bka6N4EGby3mrEc59VgFrQo+uQEQpMkfwIlebxFMf1M3Pak7BxC1Gb
64XJLFtT9wYlOT9JAXdJmGBQa6sKmQDFOEHDQV6sQfF7z8pNKngKdk/xN7e+e//U
23r89Frv6xJYoYXpqjPqxXuopJsXNCy9dnGaA9bLKG2cR2ycrGxdyLgoToPTC2zI
23qvTnmDoTopR3ClI3PMOYWM+xFEPI/tcyOdu1RtKp5+e/ld+kxLDBcZw/2tg54k
ZQQeDCoSV/X6DIXslXQVM7zUs8FZdm+UrzwLkH/NkEVm/rO8BEQG/msr2sHEGazk
X3AqsNcx9WH/jAzTuPzujGzJPgKM97wf4g39sSVNE/gzqQ4Vn8JMuRNXeaWb2Xkc
EjyJUXkPnQ0MaOMvP15NWjhCPGWZSDT4/KVGWpTrpvEFkZI+HZWFyCfe1wuByWod
DsMm6ZB8Nq2NBgqxOYhbe51WSrgOB46jqFZz1hApWLXpXnjLcswoq0KBaRWNKmfD
kg/JirIRdngDlrkbvgNIWIVMUN3WaWkhSKv6hsbaFecINKsRJOFKE5wQexG/0jFd
rsR0eeJ7fUSXqlgYkjgI+N/e6B9WVW2aaIGJh9alxiSzlmjxOgsXBOJ3/Mb8IoDm
Zy/Ms5g4Jndp6wCGVwyVWJy4g/lEaX8TCdOU/QQCtXf3qrmrApcLGNWYoRlh2/QR
NJPfsVNnR4nULL65yMInPIf8ecnEIiGiWVARIF/oSJm0IIW+auTHTEIHKgK9NQZ3
pT5RNcnOMCkg+radN1V8KLT3OUf9iCIxOmhO2ZFkb+4B6opSm8yJOH3PDmDOc+1A
Yw8ANkDyOCkDQeudl2HJvNR+E720+CYVEBvbWaH9Kd8LyebBPc2GMnIkwsL7CR28
GRwVK7BB9clayEkyBPGsPDxJ+hOnqGUslNt4Y+eeqpK+sVjjdDpagp2rVNvdkLwr
v/32vUidfxB2JFPQvVVl4tXJIb3u1+wwN9YyE+jcin7EycGNf7ctjsix3W7QAJGV
lJnn7jB/KVZ5WgbUQoIi1SDM71OgVm1oUX3gc0alB5+FqPhK6qLoDN+nKS8pZeYK
IzKE1TiMWhzcvYb5vNTWUINN31+u5L/rfUP7qbYmht1uqLx+Yp5AQct3vwT1a8fg
DsTItRTM0ZGIn8k1rGUwf01TC7t2kV8ana4yx6YqmBFaznQjwjZyPs/2GFPFYBtX
s2wfv8mTXVqipn/A61Ii2Hf5f02wSDMoxIAMFdC5Tgu0rHcUYw+WM076zIbHZZea
fMe/0Dd+8Dn4Y5deoa8HxyuWjmroDywj4P0zPhDf0jLl26N5YTEt0/Ptx02bP5c0
3NUwa+xZRgQjB3BB/DvDYURn9kf9uldv/lxMG3QL0dLPjnFe2gxTq0LPA5L6qcrL
LRv/iw7VS22ma8zK9EKFWwh0qPSWSk4xWAPRV9ySTe3D6ehHXMJ0a1sn5CEDAj82
VooRsgPEeB0Eogx4ocC7N3cnBjVJMYOJtyiqRMeKpZbncd7ps1lsTy2INCA/3ozb
aC7rwbADPazWpYSvwGcaUpHPgLL7GyLL3TljwwThJxoIdVAqcp338/lkLGrfgEDm
VVfz2fIBvySr8LlTyzxz+75c7R2HaxJ6AGI2hg7P1YzdP4aLb+jHaFXUEDuAzD7e
CLrU1CDMcwGchcmScfKQBgI2DkmJTzywXcTzdWi0VPFOtro6fxGkL1sBtgJH+JhB
yxz4JMNuwRDSD1YSgMXGq34pjn4bn+lnEE6afQ+UyxbBhWhynpwGo8BenVdklAQ5
mDkV7x7pOj+ooH6pBjpDIMxZKcDTyMqGGIgbiNCz/UG8LxF80wGywHIQZjuMBkGN
SG4J0c92IqP843CUHWQoJUMbfLWNF2xLnyh4b0ngr/vF9wbGBH244tqzhLD9Icn7
i+H3ynIy/Hv5QqyD40Tpx5II+R5TJkAg09H0RvqF31GaXCTqSCM4AXNNF5IqEnmX
LF/x/XK/9Z57fDx43aJXJLX1Fvjp/2WtD6OaRhFa6MhjZgZCXSvMGMA80Bx+ku2p
x6J46oXqXQhlFvQOguDlqP+QuCI/kFUKzjIdPX7gDYqTP1PtCY5ro5dU1x0/UQ2g
8IUKe33R1vv3UUZiM5HjuyxbJ3arlVpWZPZcDhyRDWXFOjy3tVv/aEIh+ytzYe0t
mlfZfB1GuQddK6AFQLmshbJ4cVpwcvj5pzacKSLrzF7eVRgcjeHlqqD/nUfopoqZ
ymMaYn4WwRQmiR35e1nHN6Q1BTIL7WFiLO5QairBleS44gmHdAjiBern2HN/DZFy
6/hJLe9c9OAKYvqW0QJttoxs6PiVGBFBGdDZ22/cxSF3WFs5WkWFTJ9/TTM/SXx1
Gl5YaQpq00nKDgiIHT4HvcCjd/pnlYbty9SNEfFGbNHuGcgECLnyZ3A+nWxdy0VM
7wf+2AAhHLRX7+Wc8iCANnGpvTmlRzM0Y89KM8HBvzRj22+AQU/Ms3egTc/G7vIR
lMxv2deggbntjf04IeKbBkGA0T591BOg0odvAP4ARdW7YycyEYObNrJjvIaAnJAE
nrePh5ieukDZ+AsUY+hklKvNnYrKjhtSPZLXNRi+9xjmK3+fcfZdXWB/WCdJyjNG
M2H7h4n5xVIKGNft6HTCf9pu9//gvnI5xFK/q75bf8Sqx5AUV7Z3xmpeWkhcLf/6
LcdPcNL18j2sXVy1carBFYgDqfZ2VvP5wsJVX/W4BlhGtATpsUyyXwa3jfePHrNF
G+CJVfO4BKuOrDL3LvkYfmmgML6GlUm9vgSk69kH7GKtr9kdM5ujWzHotBdjk493
obcaosxUH/bJC0gVjnUqrWdPiDdfw3V89sh0pwrcE7ZUEB7FAP9yxEkw5uxVfmM0
tooCfeqGFCq9Ee6DhVt/5wi5ve+DRjUV5rAO0c/AajAw4HQ+6ySx3wCzykW1qNiw
oc0qjrzHVMHocDL/n0vuMa6Cyvuz2aEf5kyHo4J2NGCIQjdAQUdYchzdL9SE0FZl
B8zVTaP0UgV+xBXj4Ctr7e9ONMCPVRXm/Ku77oW7WMUyIgOKixA7QZOwZhM1mPRi
/h+b2qzwvU1es2kpHold6gpt/Jq6VkXevtfRUb5tJBkql2nJS7z1cOlXkHdPrw8e
tcewdlUTqoLJbgUp43HI/pNQ3LfhyOG8dilX/FV8o7mop504QlCz+VR7qifwwO25
LpxHhvEDfGf0lFmbjD/Tpz+7zzMqyAn5tPewpLc9XU0+yrqjmdLVKdPvQEDLGE6W
vOzpAZ/Rrt1AJbYMS4vpjPOPbmZNC4WAv6ltgazwTqHAT+c/S4ilC6I+fNAUIj93
4Juu5/9aXQvQC4AHInvvGBUeYQILxpYzyzStdhUjdOJqUZA5em3bSL0vkG2T2n14
/F+vjbni2aXRhA0k2TOxFis+A6inpYbgxUwNYsAMOZGQ0idW3K7HeBBVuvF+hRs7
D50HKJZk1A5cPUjQEof5EPT010PbxxVBkzU72ozVJs+/BqNgSSfdUhVbuMTg3r7s
xFPxCbIw6KYeWQ2xjnVFv69Cg5hZbpLm83XBs2XrEPIJLw9cAkT4QPBDXvbQubed
Zn7FIXReE6SCN9ZexiGoySPtI4YEM+BtMpFJY6Pvoyj8Pvhmh1fX4MG7JABdutkj
zULSGGNbC6mfJaIc7WgxYbaLq+TPri1QBCzMBpsXDSutaafVZBTPeWN/kv8pQ4Hc
6JTIxM11dkZ0kFTp5jKiLY0+4VXEWPCRSSxBXhZVrLL9nbtYPNBWDEPOw95gGZ+R
KiJ8RFfrLWaDudHtKUI+vjcml7JPAWMmyKzQSSzIXUdEy5aEcaM3LWGm67Xqw+U5
+3qtLCl/jlg/sGlRLEN+oh9cD3doXJkvdHloc1BpMwrqqB/C5kHAWt2gOFXqfiuP
mxUBi4Kd2WDVIsCMnWGLDXQcgi7EMUiNLVhEq9mjLuMLcbEhEQ+++YRpzNQSwSdW
xO3O2FXpfD8Ge1Xm/mg5nx8bdSllK5t6bbm1IAciuqNHRuh92GtMGEQ+AeAnsEXs
u0Un7pr4SCw29TmsNH7rMyM7WMokMgoqv1Tbut2hkgnvw0TRhnxtvUOu5IjkOydt
T1Q+KkUYZfxyB4BzG/UCoa78BziInCVMJ662OZY5qMkLBV2MpS6UQtJEdJUB7Cgf
4uQgppyICVxL474amCUWv2uGXRboaxqD5h0ynBA5tVoIkiG8WDahpp8flQNCrjIA
21/+KCtMwGbJLZHQKu2cg2p0zQvthfNSLywxrzIeYacbZoW/Cu3DVhSorCMtUw3L
/LBU2KHvvRY4OlJ8DfJ8rOq2y+rK18iCo3ckg1QXQMGJY/uFwfHm/wGb9qL50Mra
9RRuLDDuxNUv3oCNwkWPPEedZS47Yq4LJnag3ye5+7u910nb6uHig559sXQo8Gxu
+6QtV99vp6W3Dh/jaDO8kLf/3DihB3y+NxleQI2Wa3LB+FcOFiN+cT4EALCEngTT
sw9L/VEl/oXyNUQiy79OYBSh5OVkoyU8OEy5LIQ1VT6r+MwDi1aT8ndPbp+Sgz8h
P3E9qMaoOGYiNovMGHYZdsxqMxxNcyZR6pcwZpMr6oRURSSs57AgwpCCgbD/v4YX
TFKy/iNmBhv7DN5WVitWAx5Nu0vKHjYGp/QmTRG2POgjlFLxpigxD8OHFas1Wy2b
Tg2umdQo8R4SWCMNPTvtqIr6mpZXeNTr6tiS/QEBKabpB7ox42vygCH7rEHn73v4
ivU0BRJlJMn4HfYRbaI/zC3pxAdZUtjG2iJziDOOE4qi2mPK2EMoaTtIpGM02A7i
+5YdDBqELbuDruJO+9zBiKk0fuHrbCGE1WDmwYKCT7k6lClDgBp5FDn9o5iOfT1z
fA3TTzwdS2HjUo0Bf7DbxpVHAgIihIkRdwTR/mkIf+kiV3VD94Gc5mk1/SPOKcyz
DywKuOxb0zddsEYofXEvq3cYcCFK8Ygmslmpgdecct8WKZS6HrhxAJ+jKjohXaTp
gIMXYGbEN0huBqERB5Pj+pSPRwqPHNJRYp0NC12wNr6qsPV+5/DgM3a24wz6Bn/M
XnX3BVii1PWo/jBkISRpIZNO3xGOcg/scV98J8Lw4EmKH1QuVCwwWBIEmdU4OWMK
AbfMjDIrsJg+KA6JQljTGLzFtT8pJjEBEUpHEKB+N5UCq6ARxxmoZVI/u0sS77qY
ftzohTtefJcL6FxdYtTJY6powpRfp/gwFGv2J+z1BIA9aw44Ey7VwKMqBK9U3BqJ
IfQ3vXnmmHyetGM3um5E+m82zDkI/tR2MrtbQx/lDB/e5U3wyDYmcMuibnQb0sQ2
hMTGveHiB+nwMxMSYmHgJD+wD9hxKi4wG1bIFLq3b6B8fd8F+WhoNfWY/RmWVR13
hWqDBYZ3BBCCHlXyVyUwWe37H/R/gcIjKoEFLH9tL4AGEZruh3fQqmc1hoTF7ahX
iLq2F9UTMQZ+DcVRZxRigu9qTEDu3Gp2vDn+lOjV5ySHX6vahpvk1FhDB5ja2D66
m7B/+X5KhWV77kCIwyYBP+r19YLxUDE9h0F7hRSu7aqlfWoldte/hYz+h9PRD357
HbWUff1MWrVS13LTvlIbwwyOfkLlBnI/KHrAJSMNaUnFkrykZpx+idEZC/ksigiW
X1DknOSTAUmAItZraksiWewKzdweM2naASejVv/i20iULp7mSw29jvBL3xQGpAaM
8rQ2yx5qj411OFzEEUJnzmzXc7FdJZVqLRIm5uRrFQRWe+co1k2VbskXeaFjd3t8
usDQE9MDciJKtDbDMeUDCGWXK2JbxhOrB7Qx4mf/radETdQ9KsDkmyJtEuKBfPK8
W+pgr26LkxbYpr/QRrr4RFqbIsPVoHnjyM+8ksEPe6P++ET1bdblt4VI9Ov8GBx8
hjCYsZky67pnOZe/6om55LTuZERfEUBGPdOzIOuZGeeVtUK7Fv+M1asO27jbeXQb
aZug/t2UveVF4m5kcbrkJ8bUVqG8GSUMkQ/26J/zrq0l46Q1lKh6pS8zXeTkUcKS
N88EpLdw+EqY5Ac7n1ZjgRYDEUhnyQNeIEhji0lRCY5gcVl5xfxmlX0DUHNhmc0L
nWPI7DTpXH+/Mw06NXFiPG19ubSYoCS51K9NOs3Vk98p8q1uDV0JVvn6EJT87ExW
IckgU9nDT76BZjYIuwi4ZMvrqphBkIsnLcV2QkCtofDjt31z7xUcBFKXzhopJAzE
nOhR19OSt2X5eMD/9Nr1Ghy4jQJori/CEvfpwZCdCcgHtGhp+bk4jLJtcJxtJzLA
qR1ZemLw0QH7GxG++o8l4pXFqq0O4jRziOXXiY4zil/W0PhVhKzD6VAL7REFo8dg
jkGM6msvMqYrvwwqyA2i0HMruke9qysgw5XdZWvhUYDJlp2+yePRmRhk063Fh2mC
rvmlwCxcOlbNui9IrM1ogoSduCD/ePGreI2w8REdav95rBsdK09zijj//8GP9Uea
dm6097XnlVNFT1TtI/CinQYwaFCQwaTZ12k8txowcXxZYJt95y1c0Ts5OH6WutQK
QU6rjlPYLk4iYsLI7TxnUeFyCmrmoe2CRaQxFCMoIDzlMXTjwNmxEOexCEfA02/E
ctmWN+fG7hSYZXiTjcrCAI2Y90MaW5BDLiIa+kabksTVr2wajgstRcQM/Zn2ArAx
/OK0vmoPvBLOPwzB/85IU+hlMaAmYHYgJBFvz3RRYBT4ijVinOI2jQSy7BD+XxC4
CNCo4+0D0DobHTVSAGC7OOuBPQxLzrdEEeDLMgJfzF6uadbNCGeixrMtrMFW8Hgc
IDeBICro6VBN/ByEIcCc0bglqY4rU7S6w1kOexz4yEeyHnolCVXWu8ZxG/seV3vb
/yrCGssBNmdwCDIzPP5jd9Z6c7YNGWc4Y/Ubya362yyiohpqDtMOfGXznw47jhbF
HULTUV9Z06Gya2CCKbzmIjfVn1YUNQMhMBzh6gknxQXI7h5H/K0nFRo5t7y9hfQV
mymn+mpQlyFgYMHsI+QpgLcbyqG5H6o4Zo0aHWNJ59jZWfNb/jXqEjoqRTcP6IKM
iroHbDW34qYbDmyZAAlVbG5LfadJU8Gqtz3LTY+EjTsPBaguqM4ho6H/XdnzDaN3
7zkH+FMdd60AtY+4ZPPe8VNIQ0edb5hxcRz/GvAdVhysfzcaFlANfkfrbbJ3nGp/
SmszYBxyhUfmSHAtQrbAG4C++HudA9n9WT8Ae3AFzlTNy38d6+1dHcG2F8DI9x8n
vRIb+sGX6ENu6nePDf1IiHhpGMBvrv0dlpdLxGDrXghGukwvxHItXoPjVBPyUYiD
B/+sBl7TkOdQVy3SJQlNWR/XaIQPaOAfDJOVW89GNesLoThAaaB7zi+HtIfbN4nW
WyHs6VaKHwMYErmCmkwE+qnkKnE0OcaHBnHSn7FpE83ezZw47SLIL5tMl9QEtds0
6O2XN5f5eLTundqVubQc0JCklvNbG/7z/z8XGtOndkyb8Ind+Vrs0gl/Uwq9Bal5
0mbVta/sgygN/NlhHYV1DkGtTRiBzjEUpGuqbHo6rD9heVSerP/kaILAQd8kbUE8
ypl6kaV4F9weT8hdEaldDArx/x3HLy2LGn0LvHsefWQk+Y1yCWtX4w0JJpEja8kC
AocfV7bJx1hv8f5M7bkxyZhrUYNwXR1ECSROvb6og7brzCSqdi1ZWGF/zm4eBTz2
dIsMmEa0/6gXFqmJIFJGEDWavrxMKmPNQc8MgTJyyok6Fv19+ywyKGt3MbSWJ6bw
OfpC008fMUJOirrhsuCs7993TfrMzl3cs5jZ9SrCJqAOx9CYhBkwd+GSFE8T+2gt
Qu3XUG+czW7Y5VWAmuoM6M9iunwXSOZd2R2cYb99VkAb+07aJxwzzWRPGihbObI1
iB1LGyGP13QAobv+TCr4Sz+D7nHzQ0DK09OK3o8GilQE9Z0hXjZtqmOCgAi+YyuZ
B4oPa5ulOT412vclxFkjQpCoVTpink4eKNb8Jo2NyzCxP+3R1kx76ft81AdnspnA
upPhWdQ3ocy9gFDV34L15p8H24HOARKw+qjtgfIST3J/GjNzlB7Tx8IX3C3J1uOh
SG6yyJBgtCoqJY4tia8LICwDLffgRE9EXHKjTBQ9eih62ZY0F/3oOLKOIanZQhma
LHVO1bQD85X2WGngQwA/7OnFVRhQ5AQ+7DPCMd1jKAJqWHPaLJs9MutetDtqbYks
AdunMzxSr5vtJhOqgyDJpJSRM/JHd+I2/q3hpup7y6XnJbSvNP7195WTXjkAfBKf
2fCAflGgdVih/RLHY+mrdyTNO8G4KjCjruDV+rgLjSCL/JiNrmBoR6qKH7KD2uNo
8fqFrBXXM4dQfygEKy4U+5jgKbrqXd9aL6jW2w3sweFX2OkQ4qXuWYJk61OPHaLk
wkJM/JWUFlrUgh6sq255rQcxt+6u41uFcwtD5o+0xHbJOu1LUZWx/XbTpTvmQOuH
bZMpEC+jVrzPyJ4a905wtgsLTF5X9zGtwpBrY+fA+g1RexYma/2kPaRQLKzju8qV
I77HFcNp6nNiOwt8xuoxRi1M8vXn5wdIAM+LFQx/8ziVJ1jY3RhlkaP6cFkJpvDm
737K+fyH854/ua2gq2wAS5lbj9uP0wMzvfiajDZTeNmtWZmH8OG0pdY+Bs3w2lBK
UI42sb2mV2sCEKJGiBv40p+vgnEipUcExGbfWeJuqT4zJN2o/8B3IYYjsZlxWIxX
kIOobLGN0dG3WHkXhPCNpDT8yU0hIP2mihYPGJWznMovaoRDM5EaMJQRfY1P2GAJ
LPgO/ttVMEc9N80wL8FPowyOE11xuUNPgPJ6q9NItMWIyu2AkFsGve1FXW7ymmIb
ZDcJxRHh6/Drru0nj+n7u93yZUXN/KQ0FsPPxXNOFP1ffwYu8xMguDMKJBlYg8a1
EaMdZsWxhtn5QyN6rBJykkCQVh0686PNihX5vGcwrLD8F/m2SdSX5MgEAcbbOMAK
3LYrBNnYdtZydQSkbouQIS3+H/nvqv/9bImD7XHNZBLmB+i5wrc6guWawksogCXb
xZtaNi1XcF7dSWd2mzuUckUh+nqgk1mLb/xjrUe1Nv/BJToJf23yUHGDu2BN6Pp6
8XERsFA2lPFz2Edeuf0dIz0pCX8CrJPItn3lYJVocmZ/spDsVms6Dc7sl4n1rxZq
gso/ETeZqSZadT2UzLPxDP+CobYPBFMa9WGUC61CYn1jiunUoMe7mp/5Arvfzi1j
ecPtVYDKMzAA8fEQjRmC3x8Y6zybFe0PqcLyDYVZfItRr/6vo8nG4qNrCNvRbyym
bB+S6BJGWrSPTN5RWLFe9M0DaybjY9v42MSXyrdCXVul7U2tzzdaQd17oxuHxvG4
maLyU9UNWtTrWB0DmvoEFOM/EmalkziuVN60wCmMgfYfCJn8c/x544MogtCehtoI
e/X3VXy9ibOp6TaBVozAr4STHu3zV9EIj7mopF4Nb+QFjHxTHBH/JrtiVSic+Sxk
/XvX8vDheNbvTGRXTwF37//ZPRNswqmC2b0S4tdLgE12bV/j45y2lrm6k5E7tk6a
hiWGPdIq0Y5eZ3RaA04gy1cQhi5a3e0ptJ17sKeXidNL7PHRZk/d29j9bvvbPDxu
fiYRY7jQaSUqk6Ipb1dfinN0i7AMYrIDL7mNp42NLKkIX9HdmZ4RJ/3jhOO4Rs1O
4UfmG7vt2Y/OoDu+Vf0cV/4uIDPLqR5nDfcRORP/Qv7xsPyy4ys2TQx4WhF/M1Wt
OqfUNYMr1pviipLFZ3EHIJBdIiqFL+CykRVtURcVmK/oJRIjOAe0k0nYlCKChEPD
eEbsZFm+C3AV1wRBS+vRTWdSU94Zes050TcNxct/FvMha5d0d21ewO4uoGia627l
gUA8DpzWdLoEIF+GAuurX/Mp0zXsq6VHhBDNPRlAm5I0U6F8y8AoJCvbNG7tNo5C
xuToSZ2goml7GTz7Ob9Aod8ny8APbYSjYij8Eh0+IXH0jB6Hxd22yEhtvvnnVZxW
4fstQuC4PWeJZru1soo2yafiUs05O0QUHsdZwO1sJdEhRat3ZKnswd+5Y4ucgb5q
GWahCUfo3Q5teZPGGGrT2rUh5J1N1be+j/naAJJqqZ0ON5ArDM9za2PWwWOwYnii
JWl/04Mv5jei99FJC6EJzt85WJV+4ZrY3PcYI/ZXff8ai3JSeF7Fahsa6zhXjyvh
WDg1ltV+3uHz7rZGgMZKW8z0lI2dF8gueUhNB5x044wcsfO/g8FFQpRqRGsYTHQA
y+eyn2f79tNpRPyo3Vyc60YVnL0rrx0hETs1aH0RUtM/KJZc2Q2OZ5M2JrFWMqbW
mTrycqUo4kkY0tMTlfbcYv8BtGNmziTB6/BxqXNtn/XmKYVCneq7gG1ICefs/th5
t6gs/NW9cK2g2gO/UyOH4+thDZmw71S06oXc/VmQvL5ysv4OrFzcjaCKlB3Dm8vK
o3msij+UYcSQoFnQ9JoZ50kBMbGYDDs1SthBHXL4NERI6aRo6wDKVbOk+Dxd4cPo
67uCQwp+AMcPSDB/NazY6ODCJ8Dm4rd+rLUuvEcqgcIuwVF1Vi34e1zUh8yYivR4
M/XZuJDNoU3/u41jBRuTIetG6+esAUopA6zBj840sGu63rwwFHRYOGhnriNNet/X
v/4ka1ejuiaKU5VhkzXB8FTrg8dQDhmUZ7njY5+E3yX5Lk+DjC5rR2Co2FvF/Aol
GOMeqsG4mfVfRR1Qh9VFOdjLOV+vooUE92KqbzpSQmx52+dZbiXYgGW3+xFbPnvA
IsfdLvvONOEUPptGs2OuFkeV4ia459ptoXcpnZeQXr5Gaqliuh+PC/pKlXwnDxM/
W2cZijMzmUuK5nB3mWB7wR/CS3gPMOSsUKo0NFHMbypCv35fhotlBH5f5Xqn9+nF
h091kpMeEQjQwW4nTnmxH2leLaVEu3gH9HSXaa6FHODW1xzW8BLl+Fgy6/1/OlOI
DmuzmFvI/c0Y5dMfiTtYwBvXsdLac+1l8K4B3KJYL0mgmEmEC7DFTuIoYLrNwpcE
FwiuHWiir5xqaMdzYft1ZZQnFPqGnOpCpDxwTIQHsNts2CQ1XjGLb5akR1ZJ6AAQ
miWyeFd+wO9d7UhKpIa8UGstI7gv5smAWGnqi7efCccYQ4c7B67CMQ8S3CEtIPMQ
1nDKe/tMPGjIiurYgzwvSWTXtgwy14n8VtIW7cQHwnyJ8tW4w1vrICgWJPwe016Q
8PGLBH+ZK92TECtKxmewDhMK3lzhbphEunn902+dwScWbhgJjrETQQJrvjyXwRnf
HJqIy/MiGAOoNYGCRSnZT7K9JqkUCz21TsJGNoxB4Tebla6HMFDpIzVEJVYsUxjO
3taAlXy3ps+yTkG8eiXUXClNWPRTWl2i/k18lmoy2WC6IJljBSMOzKV4vK/66h3O
gwBkNAseam5Uz67pa/78u08HoRzTBI/3IdxihPCVxELDZlNNprkfN0QkuSebfoQr
opE8Rm0/Sg7ViGRn1JXV8z84hJmBiWGleIygII0vDtDIek3sO1Iud7CdXVuRIp/Z
iHyaK5MAGuyU5BPtos4xM+9Es8qtMLMAPqqWP/ufbfGLqSC5sLpzvqZ1Yf8neO5+
nMHvfhjOlVVte3s34ZkZE5BV66gEtGDg/6LPDqK+oe7Wb7J6Ig51mpBsnYXUqQZ+
+2uFbDumlaxpgZz1rpHsPDlPSbYbq5HzZBDHxF5uelvkXpjklX8fLSvN9pJw51eR
6P64Ko3g8bbCah/VfkCHrM8IFgnJhQFZ3o5etTG2wMOTZsBhTaYYq1nlEiEjgZpp
XPS1/PfXK4JBS8l+Kk4awp5fEC0+AdMVvkXGmqmxWP/ovcTE2SiJzOHOUWU6uJ/7
Js758+tSAOpc4Bi8qP44+MMVmLgBDmawqF0m7KhAsM+FUNnDEtcPTvHVvZXX4AsV
gbr0iXSgDa1n/WUih4Z9ABj6IRy9mjkMRVLGXfIS5lo47TaXpL2/kaYW5XM4Xix3
5+k+t67rbSGziuJSm4LMsPSSyOe5yWqq6uPnnwRvh/n3l5Qwe5rMOAl83QPSRO8V
Hk5m72+mAYNhMJXNIdbeYUIYmP+7q/8WjPz/GoE5Hqh1udnxDAwGAenCqMNyG3ya
UdoIySVltJx2mrYNwCDGKd8IdN08A7QvltijW53CD5pOgqcUXe9fsv52sw4Oe+BW
oVvRky8OrRu/3ESZ4GT316r37P7sbfxIhUPkZA1OY+i0cEwao9uY0UI8GCZLHmN+
OEhDygp7KXoax3lwuwAH8U3eUEKSwpqEqmWQCq83f7HK5sm0oPHCIg0sxZtUtisq
A29RNHPVFa2PGN3GuzwNaMNPclADUvwDsrdDKNcVfzwUbC92Q97/mzD//O45cwzW
0IsAILmjBWekTorKtMW+d0N48Kpd7O9ln1mxvcZ95XFMFKw2vSaYlV7YTGY4gSj9
cJjdoQ4ulC3/MHV2OqcZSPwH/DUOxVrsRpE7KHVsEUVSaj2a4V5FIcfgEReGM0KO
EPxsJIc656zYaVlPiAJA39WHCSbDqBZ9W55nb1l+z7q0jqrld2zzmPkl+APRyJRV
jt6YBl07W8xQCBWW/xtcPI7ar6Zxpiv3yEpMDgcU4uXOeosQUO9kFkqw1k4zWg+G
OFm2fbj92/f8Sd3DAUGr4b/lsqmAz1TZJiiHmrA9gjCAlDTF77KrBOUGnKv+IOBW
zFSmRhLoo6Av8kFXgZWiaq1axsnIUg0GovMIVJYqzROrPLmME46ANEj246Q9jbZD
syZOPjKXPdN6S9/Pd6WtTDLuf8WBwpbgV9ehf8XETAuYFI6Tn6H/GhWhYAHTD8in
x3lCrOVUazwNXq7DpVkd/78pprukJrJdDUJZAs2pxxAmhAVPony6nLg8kg8Ga+N/
xjE3CHTWxOaRs9PiUH36IuYCqNxcCjT+wuzL6wZa/Nmw1deRC8b0N5/xHBtjcN08
zYF5NVzzixIn7qXQBo0TRhDSd6Wp0NPDjKWdkt/gyFKMT4+R0c3e7c4Smn9Dtvaq
jcI92XzX52zhx3me8BGEhsBoZ/kC61NPf2hxrv42P/Nldi8FzlEqLkGZDzyjHkHm
ocNJ5YaSQ8Q0acITMZmSDo60GpIV0xlnWAxM9CXQfrJvOxk8QmcoTmNHv/wbYHFC
F+ozEmK5Nq6VEf7awIElVlE7eRBtoOqf6jBxpc0BxdjyE0Zyv7qyaCBytwe7v9Gy
7hLuLDwsN7XZ0p62FGUw4zOdiMzI3uN/RKinPgoUl4lQlIwgk2eWaxVxz0AFAfXc
ugfsx3Ww4TA0p8cB8mWdiIgjH1UwY5O7CJcH62n7hHxGV+l+aD9XN4rh3rvCryLF
wbaiIzLUXgUXqy63Ydw+RDO+8xPGD8sND45X+1VpHrOKmGUz5AshX8GSvw4mBb1F
epXWCHrSca5gK3rqAogrMJ5IyYZFI6r55nO08niMhRKvVjm2Yidd/qcBaoh9Tp08
zRRxtTs8f+DQoxc0MBG46odso//LZWqqc/7RGvRM5k/fpppxPzujcXqstRJgvXY4
OFP2oagzX+h9IEB9lKB67ur3XewEcN18Uc9h6PWrfZ55/0xWQA2PuvnM9QHGcNkh
rrEK6thxCaymVYDZm1R02ogjlJf7cPFN8Jvsd1mwjEwofRXbx/qtNeP5SRBBOgma
bv3TmI5PcGkGCVoH5s9XxQadySAVqPQHp9cC/LJqFqIlsWMmQbB54lT9LcoLlkic
y54l/ACo7At6bzqxlYoQiPbJ+RivvTFxHDQ1Imo3LZ49z+DbkYnZVC7420R/wnUb
YGNFHywUjRYcukz25h+NfZYEefzrZA9vXWdAE78HJNwrgBQPv5meBPc8qMCK7qho
n9g75dQEKin8HR3v7rUyvZgyWaBBZTQCyjyNASv83u2VUcPrz60Jzey+fr2RH6KK
06eM+T/ARCLdYlPQaCw2RhRKFQ+U/880DSyfytXAGUHZKOXQKVcy0ZkFBABqRIX4
9teVxfzOh0L6xybzlnXWcxzZW+kQoXC8Rdm6SGZZkV3pR/M8oZSeJKDnlmqDFPNs
AGSOO0bXsN42u0bRvSuwvbVa2qfiSpQNZcQoYEWLDUkczPwa6d2/ij5pCbtzZ3pX
BJGa9dtpX+yhQz7ekK7zlg4B46YUIdKC2dG4SqWmtkaPtJDOnRn2pyk7Z7fbreYI
sg6OTsV2UA7xTloD/z5u855v0wRgcy5+48SfymazVdmM3e5H7fX2kfAjA/GI+3KQ
crLPOYcPRE64rxKcVdLTUdpK2W+XNUWiQd57md45wvhSCOdFOgTLsmao/+zGprBq
IHSE4eopMFJG8/F7ij5AnopbcYOoiExDIHRhIsTVwxAe/4poAPM8yxArxq4KTl+V
Hd3hccmHPWDYCLgVB+enfLaO2UJEFdRBB+G0fgPq3zQ8XUqXACQehVAYwwduCu5K
hFp55GCPdEWONgpIolX4EILw0PyiuAw5/nSc+2NHQO17UGzoJ7wrzgJ4yrirLc1Y
lkhFCRcWTM+2HLvdIFtTDl+NAjYWvug0lSX5h0uUnt3dp4YRhLSh8Ey6fwoEJf1G
cTVyprIPwpGpy2VSmMaIF4DLCI6G03tElQsO0A6PTHCwYxsGSKADCujIGVmAIX3E
t4dbC/suXJNAKGXawQi15G3Q9tEAWh/QkWOAZJ5XYtJGJeWpWe9SqDbCarVxtSEE
wNimTGoVBitihgIqlcYM8xzX5munHe5z0ksUVc5d69phbJGYP+lcyOAI4wpvWFQk
e0pw+gi4apn5tVXEYeWF9oOJD2k928uuIszejIdQGDPzh/uuYOWe31iU5sW+zjlg
c0uy654m07yk2I27aCZKI6vgNb3WdxJy4p4bi06+M9DjzgHBlop8c6MA+3fREU6Z
zQ/eaVAuJC7+PsIKtuQz1N6h/ksoHCGd2G5a1CS7OFFgJmy6Y0jbUVJo2Kx+4yrO
ATP+MReHgr0RR/1U7xUWIwwBwDScp20l/z9iopBO1ib5nRtJWOlvJz8NcwFwFqnc
3vJNExabFf8LAB+RTry+ukMkSfEKV0ALgYz6IHASKIHIsXIc4jRhDSZntVhxHpkF
WzcoJnCb/UBpZ92+MXeIvXByQhXKTQzEfTloqInE2I8bWp6NnrhoCo9rSgGXCeAd
3HL7tN1UyH7xhzj8lnYDEOENEqvwI3dWkYJqYW9eN37EiDo2xPTvQULAIyQT1Oln
IPBdsBHoKwmNuL/5NCkSkqiL5sS/o+94jJzZV14NJMMlNbghuExW6n2wvY94Crry
ixEWFh/BbfycYVvkVSRCGVw3eri/ht9eGTFC3bJlhHNVALu8Wqf1o4iKSeoU008k
s6ijOdZQoe6TFt5fgJo2u7tsYmno9bzf2yqBc0jB4uAOmhZeQ+zOJJwYmMCyWQO+
evbCj3L7FCZE91PhY5AZAFgS7iJLPiV61WQdc6DBG2mYQDf4GcDtviVrB964aOn1
JPOA8l9kOi+K4vNjIkiH8Xn45rWWM4CwcwwC2HOlqpiwScgvMEyuXymaxOhRmRaV
CrJfvRFPfzcYN4Du3YBywHrSTh6neNp9uKxbMGjgSRoUIxISiumLAxlsJx96Pqdq
jTEkBJ1vWeyoak+h+Bx4Qdo52nChutq33pwWnLOI5FRDKfwLSVm82nrVSUCl9KV0
x3MudPhWn50WBIinCsyUmbks9ZawXAKZIroue1gPog2xSC2MAjJ49eIaRly2txB5
ZlnUphwAHfndQnvCCTz+6CT8JsRFjRdSze4U/I2fjEuBlQsJZ2WI2GOhYYoKc+it
RVNaNzbrB+qEN3MvCpYy2qbr5bXLFnowKBdByhxU73yGyVJzhgKZqYdyu3dbb7WO
orZ0okLLCZ6l0ZX5A40nDTkF+YbBY8OhXoOzalQIrfNQwFNULErc+vB3l3n3U3a/
KZwrzkdqzWItcHCOBvpdbGdTaiLayA2vzQx2GISf9QuwYlmvuuw6BLuzTnQ6+nCq
F35OPWKB45dJygA4Ho/Nlz+GKty07tfEPm4D0xNF6kRgaubZJu+lAnoFpsDvvCzd
9bhQ9BRmwc7MKzz7+mb4RfIShUqk4zD7lUEtKmDPErAImvk2DFsZMYiOP1uv9aFL
G5+YMbVRwOik7dT1vJhMuT5R+f7c2Sg7OJVwqpl4wDiL1VgQwMNDoOEqMnDWKQ2f
D7hjVKLBuuzm0F0mMakabwQ2OHjvmJhd/69nPifjn+LQqytDKVTkdVl4Le9Kih7I
cT5SCy7agfPDlsd0LOSPKsWIR5gKV9putPbzqluawsGcePq99DyuGqOQPaElV50l
nH9g0Ow1bHimgAFTj/y0pOHVKJ34rf8cd+qmbhYRn8NwecbaDzI2NRa7gwkGC5ES
YEJHYA5luq0GH6slbbV69Mj43/JBqQFRSZJGva9i47Rl4mVJCrDA0vsoxDSSHGEL
w+hkBkpTihtpMAygVXx/zRLfTg350M7+Y0NlTN9rlcd+0EJPjnQzGViMvTdZpRcd
qiFhSvoK2PO6eKGf6I1tIDIonE+aiEi8kbslHAoDSht58o5hgOz+zyLlUlhJVEzB
W+nMwL5gvM6ccpNa+FOpTT8sATq4yj8HDnkoVtasOadgygq5UKI3Uwam4nuJEW1r
fI8pbbtulz96fUKeU6sG7Pd6E65iGyww9gAH4T8XqLzTAD7tkaiVJQcKhfEPw8PD
RDGputwsc409ynBOAgzd4p97YFce0cYd/uEI9hew0x6Dybm6ZeucBW76pVglnRrF
/jwXnLqPc8D+17+5tRtcQO3ZJBLMv4qmR+1wNIK0x07f/nnWE86Q6QT3PhlRyBhf
DrYE7vTRuPVW9Jvcm/uybb2HoTycG/kPomn0BvqVu4t8l+7aeUb6I4HgW+awiU4J
7KkPEzZIkU+i++sXoMXICqIcNSrFh+38t10Q/U4EZxEl/6K2rWuGAvIDnNBBsclK
IrzI9SupQgbIHHVok2maHZuHJus0o1zYnX8XJErjJ5VHMPdwd9egZcVpswW1mN5f
1ij1myqFIazFpZD9YjgR4p+Iekf2U0/6dhegBedth6zwny61nnIRQAu53/Fvs6SG
bb03+7AuuWQf2DFsQztS8bAlWlkEwx4lgB5hW5jx8U25youOhBC3ikd9adus56SY
fXxCHHl8RR9Ut1Vhs8LWvmNVV83uTMKcKLtgktQoYO1VP0qe/ortlx+ch7RfttY1
ina64pW8BdHpHB6VBrkDKpgi/envgn67mkFo5Jjf/yA4JNugaQqmyqirbqlhrPwv
L/mY63BJ6A8DrjTAsE1ta/BgIIf1+vd0/OSA75C3Z3F2ofLGlHs9Gl+uer21M/RS
817mbUw1EGuDHeSsNBr0zPxIq+5ZyG+fsuu/48HD9W6184TitqeLWnMilWLFaUSn
xeb/9YdYyZzsWm8nxB5okkb3qtytks7YsF/x4UT0i9QUYAbc9+gZKRe2DJ61YNs9
I5pOiIq86yMAmmnKeIzDOkU597xieJmC+r358UZzPRbSqZv0AhWbJ0eDtQiGE3kz
GLamLNW08NnrKYdLda6D7MiOA+zP/sDYeBmSl4IA1VrVNRT5u9wyAD4CJ2/FrdUk
EiOUI79fuWQVdBAdrqKgW9gg9IIB2I9L1A79MgS/46lAd9xblAy1oolTI6Nk4EMJ
eAZI1aSF8zcSyXHn1fTtA5CXhlSMJs3WojsPhupqV0NEInDiTU/9LhA0J1wCnma/
WRsRCVL9MXSDKTxCtlVfgtKt3gVWgjYMRsSkoHu7hUzSFbvd/Fn+yVuVKTN2VkpN
6ShOdV6M+lgS1YXdmpPJz2YrYzG1GgulymTpVfQwzMzziv8+7mPmgxyFdy4UMwnd
9ic08nRdKeL2RaysSRAhL7E0+iK3RrdiNkW25zjQwdLNaB/0w6jjFPa6roo2vlux
wmTV1NKF88KdEi4uRXHSC8XNGLPYo8vaiOWp/huYw4XTnxeYlDOEFlWOHE2bqNqC
FeS0iAFADm/iHedv7ENrcnI2A5EUqGwiKrVD57/hFcXTDKVZAjzjkqAAVrKRWZ+/
mYsqTHgpNOWaL5GaOqjPgahg9rG627aWBRAdpFzPUZs+HyDE2OMkRnjzAWu9pMt0
20Svf6xIA4p6jk+bzh2zvuQ+yAzIu8Alt9VxEv8WI2nMTCAAJ7YJflCMXz/1wbzT
buhupn92wYAFfPyf+Cov+LAiP+gD1jI2jWL3mjIQmjakWbWR1jpjCai71ykg4Vjm
kq4CSBtbVxzXi1+6D1FphafeFwqub8JZIMBVqsjKIave9fkpA+Jn75hQiG1ya2mK
3S6WPt2QsdJ0JBaA7fIQSoUJsA11DcSJoaP12Gh5sesZKIPgD6lQ3sdbJ1EiWr4u
PNpRfxVHE2LSp1ki+/kCY8rBj7HHp276fyYPYeGr0zjAAn8lf5eg9vygwxDhXXAT
ww8gdpH/rirNeOTuimFVSwD3ttTLOiSOyvTz0in7uYOUfT8fguzMbA/RJrBfI0BY
8IzI1IaVG39nT9JUAUm7Se4rReU5KTPoZtLfV/TdE20HmQHAmrifb1ExvyL/1+2b
wMQbuwu6XiHTkYIzmV+AicXHJ2k6vmsIHGrZdu5Kt/YulfRgvnhmNhWqJ9hTWB3z
zPrj1QWjUFlt+i71f+gJOFeEjrHlQTkeAIyPropTy+a0JkqWY6dxg35Jwah11zLM
Wb3a7eEATv53V2KDI84fWHldrjRHcbfYvEsdh8HqtcQ8MuhzzmkwkpCjxT4267GP
q5/MYNs7G4IeN20f7tmasX+aCD+uRB9V4O4693i449ThufmybU6GYY5E1HPWongR
xzJLF/rZl7l9sb2MHUmfAKPvUcfycvbIimk1pI41h1HYzvDQNHX2/LzopNuaGu/X
baVpeoM/xoumn96EhGFZyXAcbIN+LVbzNpDrW7C3cE1CQ4QKs3UHWeHfym9MzLFE
Ul/WEBvbquAiw+lbMg1mmQvbgkNWq8Oyzpu8XQRJLxZPinwWZ429J1ixlOxQA2So
tXX26uc2w+mFBrVG9GcbroQVzgzuPgD94S7EJDDeoGvBurMdsgyuMu7ZAOKetpZN
d+934OGkHXeOKfp9WPJAyRI52I0aNbvMS6FksqlES6hWsqq1j+dsnTFUa1OITgCX
kfbQMPG0f9/qLnhoutyzvKHy3fdid5+/88ekPU+ankMUlgI975RejF4Kf4Ku4Si4
Fqg2Jpu5QRq7MYye2IN6XHXWpz8s7DmJPRSpG7lC8T6mYzoeOWL7Dtg6ASzXHryk
J9XLbIob2UnanrufTncqlOf0azsQ8gOAWwNMS5oHyOBk9GJkcwO1VdayUYorYpPI
K0/bmWy6JRLRKSqNcw0uo4vMDIMum33DNa6YZZH6+xAV4NpITj3EhQ+5xGUu3bv1
hlEVyD43Uj/SLN6eiMMrs8BG/asSM8wbVehvJgrdqIqQKgq7IdEIGQj0ASMdoxap
WII26JQaAAF5MElrXrHU8I5jkKFfODq3t0DMgGBe6g0E1K4292m5NLekzOQN9pbA
1zMvlf0+9iyZ5UGuMABA2H5kZn8Ir900P6Czkdl0qt7KRhQEeEKvk//AZh9PX7xQ
ZBpqtiK9nk4n++DJOqIPYQTaDRj1QuAZKCulrdESyZI5hdmX3cjHDonsBhX0b6fF
FUv4q2XPNr9MIfeV+QMA2otb/dG+Z9f983BBCm6JKkJJJB3t7ZNZO01v1E7kanyl
xpBnS6K9VRSZVtOSF+t2W2JiCMnqXHb/H5wC3H8CrKNjk6siLhSPYEqdb0uZFhSe
7qK+xXg0/Z0ZJFOWnd3NE8KITgy9F3Jz6GQrg9oPd/mpixCRO1himnJ8LR32xetc
JKxopN0iJ4EpDffxtqAfJT3Wg7CvgHcLLGnUSsMVNjHyG0XUJW7yVJIrZ+d3LEih
Nc15EPxs8XqQpRRRpjHd2XjhprD9f1dimh5rhoTEXFdl6eoFEuCgqlMSwd4tbiz9
i+qC1QOQ3C33j48D6047ywEv1eKVE286SYFb6nFvnNM8P7lvCQ2w/Qo/IwAJL723
s/6PFN+WtVRkAnF0v4xmcpqgIFV6Ec6DjrTkSplnlNh/GUbThoFJFQG7ZZv+F9O6
Ag7AtbMBryXW7CEEmYKHI13HZ2XosW6CbaXKTq1syj98AcvTq4EBrybp+ajIw+Gn
u9sL/r/PY5CXuh0zsCXjS0kxjHC5shkmS2ebpINsEcLXigOGHhhESQgRvGtbpLrX
GQYtlgSiCteQ5K8K+9eT+PGjocK1IuWhpKFtk9EJ906MD7hVnzJHQB/5dbYHgBUT
18ld/yZP3M9Az6jj/vpQLoq9224Am1WUqMoLNMYok0wA0ul6tWH8dJAno3Y+SXeo
Htzwq6BztWAw0Ik1a2h1GphDMn3XANYbf6UPv7nYFHSOszf2teJCga1y5nUqgFdh
yC4QOzd8M346bafco+MLU3n8rgIIDUCXiEVBoggRHT8BjIysfw/Z3rnBBLbngFES
ELujF0SKUEz1rF9HbNwxXK7Qp5iSCNMCrLi/GOKEqwXol+ViSmcTq+uefyV7dzSv
WFp6vY7AVHPmyOFhprkOFWzLKttI7P4cz4ypun2pawbTdifLx3WJoUGvqEcfEUlR
fSNS6n6PdvSyKSW9Nf6JQ5hXkHobLIlyA7Yze7i+KvTH10olP+8mZVsIoR+Cr43f
sdZ843mih/ksYhOz2lJlXonClwmkVhmr7cz6pU21Y1N8WiINOi51ApJn0DA9SmGo
BXZc1/pnU9MLGIWizHgZbfTlTEjh+cwLcc5Sg9JPJr/Jh9ViOD3l9RqoMAOJOJ9y
zbdqWHwfCtrY4OpuL9LyS6SaZj/GMsezk/uzIiewSdeLiFx0BWPLK3iAcc4gQLoQ
K9jihXOQlXF9a1FiVkY97+zL6JvsAgr6QahujJgZj0pQXvmvdU3h5WVMztaCXEd4
TYi5VZM3lCVnDASWrI/Qxb2gsRNk/S8OrWnH/vKWl07MGNS3eXUD8zF56Z9be8H/
+FQ4C3TsrX+ER4n2GYQxgekyy4lHrj10QaqmqgZuT4B+Mfv/Dyi8avrzL/BacUrT
oD2o9i3+jTo76Ng3ByfutrhZH6u0eMANCg/HUUoLb4lJUSp3GGIOUzrpDOP1InzV
tOtEmp1XG/nSBqEFdeZjF1CN5ezD+XD5vk30oHK1GbtZc/0lL0vshySd5Rn85zD3
Qtl4cVhnLT9K2FvgrRvL23qX8aA5NDOAtVtzenT0b0gfeuDcjJG7bYNMzQkBxjPa
9UzOcChdC0zLNkYPOjgH/ienItvB832NhSR1wZ+H7RgpXIh6EC04bp1IlSvA3Gu5
SZb0YMniTRialDUq3OcBWxY0cgIhs2fivpRQSPfAuX1hAdgaPO+6Jn8oGWy1A3+E
0Xu2zyJ45oNG6BXonvjhae7GR+uFe/sJPy0QWG7hq+tAALTjJaavvsC2STP1qzfy
+qpt5ruT9nmvuBONziLOidXdngIlWABu9wRvl8BRbIkmcDIcEnUKWuee4+M8EAxm
JRtLFtpa6wa01jO1oDC386N7skJcEk7x/e+kY+e0g2XA4VDjz0FuGN1glxfLa2zD
jefHaKD3V8ppXkSQDRXzJOlhiGX0ujGD4DZ031LgE/fQCymlsOnYCJYj6+bPhar0
nKaGKXkf7ClcsycmNVQJWXn6VxxlT6ZFSGQTVNdxU8syk/PMv7C1lIZ8W/X5gvQv
3hZJ1aSvC//or9HWjJ24xG0woAM+xAh0sdFzDZHur1pLwRAZlGRJAaZPNDhfw81N
/C6kct0kIuYS+DoggIJ1kouwl2FM00J9Gq5jnxk0cQcCUtePotjY5TedfTIT/zai
NoiYnIA7esV881L44guhyOmwu6iEbH8htPrdQGJtt+z+d5WxHCiR/5e4TVgXeh24
EyeUKNyMef6FXzwF+mpUOwJpE6HHvPpzNZGIrfYN3eMjgFJmpqt6dTVMjJNR39Iy
p/uX/+ZmyG4Rgq2HndEp2Z7BFy52vLaWoeXuBWP4t4rK+GD65oFTGNAR+Ks927ls
v5WTc/HzZUM9zgBpk9CGyliRYJZtQcow7XEAIhOMiB103JgQSUbDpwm8m6+H9gNk
CtWAYsYVevl5rAg38IlSLMbP3o3bFWwsiqU+qM/I5KWwDwIk0HC85DCbRIurk8nK
V/wk72i3t+PMZo8jFK2y7oulbVPEu6Pwn8Puol+XI4b6rUNEIYxSFXhmXqL6uMQ1
dg0U5F9ltQcVWnF/n2NWEdV3EqlRJ5l00kyv3kO43jkSyBw5GZQh/pL+gVMpAZJE
71KWU/M3sga985OLgcPUZLJf3Jy4dj32xTGzlVwoc4iJNM1TPb7/6HL4OH7ie2oZ
4f+myJGvAjLKq1r2UwWtzJe9nIKHKKfa3Hz2/8JU1+1C8gHwlRBV2yID+4N3X9wU
Q2axy9iO4HiUOiqzDORfX0hlD8N47EOsHVRdaSs5MKNnuBkBWlWcOzT4yboMFZhH
pommpIeHgVIZIY+ZFbdAjjGiH0hgoIICzbOL6LHK9UEljquYYnFPieGR8SG0sgqx
1U69/ClwA3Zs/VD4yzt6sA0p407RcSOJemtCdkxQhv8Wipl/zexcIuOYE4bhWWsX
NqR0fPLElgMMz2QxfnPXfLCyvAapGpljvvbW1Y9Gw0YF3/zO9ITbdXlXjr1EzbLj
LbxqsvFPagp8R3P+NZoykDP3HTaMr7r1r97JRrxrh9vsaJfC6aCDQMobWvmWcark
kLYuY/uC/ashCjbe7lyCFy2nwFhPTai8tPnb7NPARRCnyenftZ/HSEF6t3zm4Wvf
B/iF9ViRKm1H2255Svc+4jXhR/Qku7rDKTevDNDnf+Dxh6dVvhdDWN0NYpXv0gC3
SR9mkQVDPQfbuMwnThC7IInNPtQaiYBDMUrQzpG9sa06W48R5h2AUu3OUnIEjQDu
IaoBoOPzDBMIJkMTY+kYaYv/xPVe/8cQYrmNb0tRPNDUzdsQg8I6hg1RBL5heMGY
rolQxQvITbPbP3MLTIDMBqL0jZmdZPCiZaXRSUKKeob2jkypEYCeeATs5r1QMmj+
PZGIJ7R+jEv0MPZCnK1gtNxu0J6DKfOmRhG9R2lnq5YFmzdM9P50N9IZuaM5hzE7
+GSKZtbTXHVXmYLLQyquSYISeVFcSs1MilXYWUQ3lADO6xwEjbkvWIZ590uH44VS
Q2peFY3Afi/KkhrGd7hxeGgkY1LlkavjCppEFKQhzAeNl8Y69yMMEtgc4F9OJR+n
7KK4pLkB4gYXmr64vjMgPeJ88HD9nPODTTIP4msmwhU6xhHgNzMXpYyBSNTabDvv
GDxDgpXfYciJlpGfAeb8R9MOijx+aqDw3ueAARILJ6Dr6pYS7ISmcWLY6CjR9grs
to1Sm2cn1xa5MdK7Jpa0BZ/u2w+7QbyvIuWkxq8U1jmA0FzjBrqc8SjDyXZxGDnZ
YM3feWpIMUjMXRIorT0SG4XPGlNiZ+aKrUrZaEKVCzI8x+QK1b0m1tVxZUDxG/Gv
RZOTNw5FfXv47/taveTsjhnMX2USl+Yw6k1tlssFjyNgSO/hz8eidgi8748qaADu
BOqWeTMl35IaS8DQ0TCBj04ai6uHEJykIeUCkskXUft1tJOqcloqEaxbBIBcZ+dT
LqIKcSjhHxrr0zR388rraPwEQapakkYOm0FSoHL6LEbdjkvRefQdj2UYV7BxY3CM
rp14z9xPHxH2n5Rxr+BCWANHuZO13PsvvMVlqE7rUdhyWRXTZPFNLCDRpeicdncC
82xrUqLqyl41RhJ5LRzBBv3M1xyTbIPbYNPPacz0x6g/71SuA5cnmmJ06eqO6Dlh
DLABQOgdJ0WcT3rb04wq3mtjWFpqt++Tiv6bvfRs7zNEp6FZL52II7iXgCcJib58
40X2+Rdtx1SVBXUvw2K5Jp3qaJ50kVuGbLp8+VSPHG5ZDaMpHpkIJDyTkMbWZq2j
2+rVUbfGuYi3Ias1xIhKWlTTrp/jfsqOiVgK9IMJ6xvqCI5KXBOB5YsMx7lvZryx
bhW5L5kKvmcf+jcjNuq89A49CYalmKrPRsH/Pl++t+j3TxwzUBanwsw41ZFgTXNS
8qbzz3Lf6hNOzQHsrWBdnrKjGCcfhS1mq+tRHbkSZugQ2KO12rWCvKK+FUUhBZ9z
n4zINj7G0LMdjcN4xbEtONcGEI38okudUeDcA1TdEWl/DOVMV42/fWDE7sCTjajf
tKkSX1fXghhb1WD4PfYCWTjspLVK0Jb7vFZAamKzUJHG4+D5AUX2hC2tdQRz0zVa
5NU3uoekTAiLmNOdH/jeh9FLJ+wizZAz1xiw6PzIPnpfj0jGWD0A2IhZX10Fx5Mi
WsVI/df3L4/bLyCNmSY1q8W5QtIum+FlY3g9uZHJoRsFAaIhaU0POCG8OGk08Ge6
OYN1FAWdZeJPfei5+3ivOiaQosUZYhCgw9VqNxq5lzqy7MV4194hNRihldrgPLoN
LUwFbjSsHXcSqj3p+MhWMfctgNkf3awn2eD6noO1kMoeEoPlno7mbjuTI8eTB81P
Hl0i8mXkSND2Udhy0Z+jw0v0pG0PvN3T+wZdS55g3UO0k5BbsjlK2LBYOP6q6QX3
PA8M095Ge16G7dXjreICiHclwHPIVRhbPhtaEY6qhSUr6mFYxn1EiEnEfgV3s2uN
hWV2DyKeSX12tAVirB6N6s1pDe3/g0OcWSVDB7h8vv0l+66kvPMmR+5hjuiRLy0p
Grfr3LP1ebLv29PJRucSGbpYZonjPVoVuF1By129QmLUiHhq8nnxH8ze5VMrvGjp
VBKC/OEXyhcko0qH2SkPwxXyNxP93a3H+JA1STR0Sc2wtnL6+CBPen4R0Noyuz0U
ACEqIdtlzE+B7+BxDL8qbOa8F/+Iynjz8xQWyUyHU+fWzj7kBl4R901Huk40duqn
AY+Qej4+/nKSQEzDWzNyx7PZ9KD7NNlgoU349RTiCTHUYii6BmueBCJCUWo9vjHV
uuAmCoqpeJ8ZbOLb0e0S3oPf2S1sIQ9MJzNJjq4l5cpicu4WKw/Bq3E/75wJgODg
9O3lCNJyQTZOq5UdDkBt6p3P0FVkMjitJcbUdjkcdKc2OSS1QK0HCIyHDEzZbZrE
PmrVSIOQT7btyR9Gmo0Vo/7PdVWzICI2wFCHp5i/iQykaSQkEYwoJsdLdc+zYU3d
9zxWe1/BTH9AuEiUiCpOqKrYp+8pQ5lU6CTnDUzi577Wn7UjrIM+qxFA2oIO+7Hv
vbEoJVEsvDpzDxJhH3djveGBwsvSyzRgk69sja/13v4wpCB1OmE5TWh3WWNMP7R9
LUXiOa6hQSsw7psypMKEZgEfXVcqkDVn/KqQgPC1S/bGaJ7xSWyd8d/OvHWqWRE/
HkPzg/kwuyCX8xmbisHXsVV9ZKzrN4veaexkJ9u3Bb6j6NTqnODCnyMlItufjioX
cPaM/mYOec+DZsh3SxJaX7qLeWAGz2lSxRHs+GAHafqygJbHI0AuY1Yeb3xYeVEE
9sIuxlGCFFCaGwbD26B4+o+k2kVh4qjDjpKQeTLwTv3Xn4rxyZbd8nKASE+pZc3h
NIiuvAcv52ohlMvN5z/WSKgPlzNE/1xuHx7IN0h09J6+uWBvf+ksZ/9S1Ium1Kps
CjaZMqfoOulPVi7bxTYI1/ypPK1nCcuLyDz4+XKAHON9gNwge43DGAuSYXk6XGEI
kDCug1wvvPxfNsTVgcck13e8Puw5zrYEvxSJNy9d46/eNV5v7mYN1XU7y9ioXuu3
2ZXF7UnhffHLtcwwgNKD9rL0QHdGiv/N0bYuZyym/ch2dlMVZIgpIOw4OmI80Ae0
nlZA70SGsbKAj42BJ73kqOoCkCx+bMLNwt11nWhdSibWlBUm5jcfMy7t+Xk04t5c
0TaszvLiUaaysnUrZMjs0QyYuvU5byJQ8EOq/KWDdGliXrvNHwJ9WnFgKa6nJaRN
DXcuPLvBgkKsP/V6eIB82FLegX3iYcqq738MZYw9RY6XeJr61Nbn2WC9y2Z3kBUt
aIba2J1hxXhmf8TJQjVlp3O1YyeHcVvP+D+V+L7ClEDwsU405pLAj6xcaPOVV/BG
Vi/ajg5nIfJ2VDVFaQj8vdpvGX05SqoQzaU6G/gCoBgnSpJ8WsJTMlK0jqUtUijZ
RG0XE1n4fXAqhGfe88IqB0+WF62yuPT1QMXPD9PDgzKxJXAeeOJdfOd7vwzOuayM
rlc47rbf7iASqbxNymaFTcY+E1mwUNsKvkfbB0TcAMYvfvhwAKrF27UGnSJ9G2D/
eV1D5c/zpXPNpm1PRXtoQHCndor2yhADRXNVhjw4cRSj6NXXAKAP8E5sbB1Z3eS4
lGw/vd485cXoGoTWESLJuJ3cs+yp1W3OBxJAT75klOiQ0swhA6HLWCONh16vgXyf
X5meJ9N05tG4m8cywsLgch4lKg1W6scZBpBY5jUj8fm/+/3WIucDxK+vV8g6TgAs
LEKXZbcJnpLTwFMijfGdY+K8s/JZ0N+gU6guDtOr+lJUK1ajKC+VvLmTK+6AaM2G
2tlmzJXFJiBHZM04KDvImyVKte6GlynPbouISxDNw4S/oj1pmoD8SoM45l9iUT+Q
94AC/cEr1VY3DzyzO6xzInP/PQj5DzFNidfbIjXYlKBavJToZ5z6ro3qoUXYWkYp
3FT9gqhz9eRy6ePN4pJf426Wv6jU7fNa7dAReGDPV2U33PKs3byw6CKnDQONpbcf
0m2NqCeCzYqIo4+rH5L89a/4wKoTz+0CSCS/nCvdyyMky0LOqv0qApd26o3J1Y96
HBl4UIEl2u4P1tVusj+9JRUM93Qia8UGi3Li3ZIVaUV7Z6DJiLDpWrEeFYQXgt1o
yElcP4BBoeFB6b538v97YMpWdG+hfE1yJUGND/bm7mkwVE6Y61on82sLKj5OLk/r
NR/RYfbIX1rHqJELu6viyAUPLOn2wvTIk/lI1CGkT4v3lokLWByauOO3O/tk0Ghz
I0pBHRts6NjKmXOBbwm7QOSAkBnWLhhKdQC0WApdTvX0A+m1XkgtmkkPIrMsTKuR
fTHWeuUAq4ed5rya9qKfFWaIacYAZV6ECsJc2CkAXrXKECwymU7HJTnuXu4Ec1vJ
UDzXzij62pZnqtcx0w3ve9F4ZSrRca6h5AHRonzKT7gD3ZCAJ0X3NHryVevSrJLF
t/TLOHbXGGc7L+7etF+UVyIN7iijBiWMqYSszbeNRe4Jf4McqPm0dA6zesV0YljD
jDykP3GNNR0roB9zuciAWtLR/JIAE40I1ipuVr3/2CTOFBjSTALmJx2GVsqysiYu
fRyfrJJMHigkWGQXQZH6Fe6fG3W8dZbU59+Bdv3TEaqdcKM90u6wLxPWxxRjwmxM
Hqe3vwczxli3JW+h4ppu2TOkwBor9qCl9rFA1x21/8feaubn4dnR1XrYH1yfke57
mpVO/DSOcze2T3D3e0GgD7QkOeYEzMUQOhTX7nf5HwyHdR4Nqz16LXDLtJoIOR4X
5qMv5zA0wHo8JzgE3BL0TVKkzMSbSngL5qOTizxqvQWXVz94vBsHk+5rG5GELuof
SVWYK1V85GxLXSmfdKKZa58I+oAWaqskKz8M29see1f8bW0HhHZmzstiDugkBd5T
qrjLctJYpJduUL+1pwpcsrjoOZK79mSWz8t38RX8xF8=
--pragma protect end_data_block
--pragma protect digest_block
GYq/grGRGRIYQSM03Vd5QIk9cps=
--pragma protect end_digest_block
--pragma protect end_protected
