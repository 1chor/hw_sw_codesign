-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
NROHEh7Vwi+Hsg+q9B5LP+XMihNYuNkWaIzPWo7AeOUREfp6wOxkmGw/PZNRc7Xc
K3Gl45yrCTHhJShED8eep/3+LERlJzSljzKHV9Smhm0QH650EBVWezrnAAudJuSi
NTDZDSugEikU+da3Iw5jYM1nVIkGF1xJMfxqj3Mfmfc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 54667)

`protect DATA_BLOCK
etVzDqNBM+e+SpBcoHGZ4o1D9HyKRT/y55mVCC3S8N7bW6+oFPlzwVyjjxSccI3j
cr9IR8sEpFRlkvqOapL+FK9TOTmJ8Fpg18osN/N7kSoTJchFw2pp47gjmecgPK5L
aWz8MoSRguuWj6QISKkVKk9a4Osc1flEIzMX9rMYgbx5tp/LYqZw1GHkCIlVGY/0
4mvUIgBWui65ilyDyn66EMaoMVEao9LQbLIqjFKuIBCRk5az4eD4mK79FFOa1g6+
MuRIvVTM+OQLDQseu361/dkbO40p2++JjO5f7pvAfXgqFj0SOdKM2yJDfcwE8esm
R7IIF9evT7hXU803bp7wISwMqO3Gxvxrpkjv6QoEz/uDgIxuCgsvdZQX4WbR39GJ
jzpNrN0urLbwZwt5bmcN6PzMLCUM3tJJdYknB9gxxg/ersh2/TV8cr/bs8139CeW
K64P4Q+nDL9kQjBYg1gxWrMuNiz2+Gvh2T25zvu0JRndVY/dXaDTZsmYdoDaXKGR
A+JwFTx6sw7dhQaUq/hUKB4NiK2qhXcJuGB/W83+iukZPz0AwL36R42SH4oeoi8X
2jS5X09b4RN/zcQyyHQinKxitnMFW19Qt0K4YrR1qTabHczjz2xkQJFUlMNMV7A7
VVNHkxrySHkC6JSwb07g66CyhyZrn05yWxMiecFpbJ7sCZ/8kXVJRPorCs2zS7gm
qL3jKq9fkXj0pk2oq4OeIcd/l6zo9yvvxen+abLeMlleaCs/OYqmb48EL0mNENq3
cwYv4YCqfpDuL0YcHbRVbyLKZnMG645ERPexFx+aoxawYplHquS746SrFQfW0ef6
cns94Fxy0vUFRdtJU3H+CdosfFq1hxKOQvKfXuiTyXq0PruCOAvWORz7QrHEZzDa
ialzEnWhgSxCjxFlq0jIM9ZhM5brOGuzLHTJqKvKMWnOiw1d6e9psMRsDTRWZKL8
qmAyoH8zqsfFlMxaYMP7of4xCMjhxX/LsKJGt5qiS4DbGyUZ+uuU9+e7F0k4qDwk
7Wf5L4NXbsExvu6evm2upE1lWLCm7UnGD0FjAdBTVMAndx3mXPRteMDXbsTss5MS
4ixpCIaOhJZmvUEIzLzIOBc86LCtE6KRumX1t1TTagYCSvziz3w8gAjDtbX66vjm
OKPRT77epjJVXKvkyBtv3WaVhYMDAqtla22rxfml3gxUfOXRvy+BbVxLHX+8igzF
Dog64ROFQbG2Yzha6IBtLi1HydqNWJ7woQUsjhGgYYYgRHX9NliJpZqv0Ji6vpUH
fB0ECSMI4HElULje4iDJq487l+iA+QY55zIp0IJkLMRRn7OZgnxGOoN7+dXg7qMX
y9EFxBt7TwKfl58i3U7q3FL2VaYcVUxNmGpjkDdA44e03ZRO5imhFtw4oltEkGnu
OKuE7J1YOD7Ck4LoWk14XwrWKOeRjcS3XPzDvdKZlmwEbqixLrwdkNs/E/LadLuo
y5r/bOAFdxT82ZbvXEBvVa4ENnHvNAwe00q2kIoqYR/Ga0d5WYCRNjhuMZKaOjqQ
dAogwcf9/w7yFpALQhtJjZbR4eJlssSc0YEdOgjZT+8HlZHMV5w5nJMNEUO2EfQh
UgvOgb/aj9K/NkXxvEOSRndlOELBOIegrbpwSGkkxKqC0mGD6AKQ6FhNkZb1zoLE
A+qCHmIawsla5GB9pSjA9/5cIUujOPGgI1UI3gdd4uU1ksr2NnCi/9vKun5T05NV
siUiBkG7UdyIFWwjeLhd5R4wd0//c9PlovjVLLhvljMUhNY0VweKF1Z17tgp5xVS
ssIBTwp+fzKpNNcSY2oSkJx/HL1mHO5oDPZLOdkqTmQK3kyk+iqMbPQxM2QW/FCJ
7+4ka5U+BW6bJ2annocaqhM4SpkRW5MgmVKNcdF2phqu6FB5FekMlb3KQEwLQazI
TgXMR1lxfaDynaTeEz7khukRaAww7PVDawwJo3iWCbBUGfO5aOpKZW0jUrQVBJK4
Gb/7mkOtisO26hD6+8+Qd2V9rra6SXwsAZ2+8A89fLuShGpENgVQ2Yy+PbeVV2xl
oniiCpVteiB2JQtvAPq+2A5zJ1FbG2ld8DTHfCpr/x/+mLFlBfbBkiJJp4SdBKEg
eq7ixFkE2MeaD0FHP1qwJUrbC150v+TwsllHIBbYe7HEdJ7R13q5KKgu6GoGArY9
8aieiufhuYqLSVcX0bUE1jTybu1iabR4WOJvtU2gBy79rBnJtedvMlD2wre2M1mp
TNXCRrt+EgHeRo/WslL5bNRHgeOwO4+Hwxou+C8jiEOay6/vdnSZzbX8s/ta2vx8
bUXyjiZmeZLMTHcQ1r1K1OCpxi0n3rCrsI+ge1+7bO8jPZPGezCWCK2Ago14QAks
5ISmYDS85f8ChqwXr1EDIxoscD4F2MNd8v6pvtAKFti7JOzBTSIuuwJVJFm+TsM1
Kx66uZcGpIhAZaeqESwHMTBJRyIuJS0P3hUwWxkbI4zT3e2hSbtUldx1C2t6850d
mxrrALqpNxRLo4gfIgiHtU0bYDi1kc8f9BnO5vzr8DRtrqeigeW9yRwZ+8qmceoM
hIwhcBpB4b7MrAqkeJVjEOA2fO5tl9OuhpgYrJTNXtsd28Ok6lEPkDFxeqgeiY+E
v2t/hPfvcsJ3X7lmvddAG9DTp3Yf8PmVu1BuCgqSjh+aYoi/18qDBqZ+rFSGXadj
0liUOidB3ZUt39uZN9dKXBapEWvFoQBJCY8spIZm0o0p1UV7kIZACSvys3W5egc9
8WA3d9NnIbpEf6Rc8el51JKVGTW2GNP9isc1MjyhhkjPBq/BS6dk++hanaXqcV1J
Iq/hf/Wet13VpM3ZVtA/uyI5DCz5wW3cXqK1VxEpXoMMYs76aDLG5LaV52lmNtca
6I1mgc6m2B7ohLbjwEP5QTTnakz9aFOpd+EOHQ3gegjpjmppGWmEmEUwqK5c8jXI
zXYBHazfMN925qgF22/vaINAMyIb1tOJyollT+217a68mhR9lnaqa6bDQMvfEh41
XubDo3adAhyunyMQDEZQg8dDJrXgs93KScipxYBZKBfBxPLIfeedJbZ2oCYjBn6O
oo95DnaXrfSc4eoD1c5CyCFQhmngNEmwAj/SYQW/tXK8n0fXai6pNPO9S3P9UNz2
ZPc/PuF9uN20l/w0a3VmnDhoU9qw66HlDiVEBhCXWV4yNARyc0KVVOK8Hjdfzw+b
6s+FA+Z+izDlbvkkyk5xSoY2E0cM3vbvLLGYTnmvAM0io0XjDfreNWHkc2Pd9iqy
urEdyT9n7UI/scXDs1miWdbnGRSrRNbTFcdQpXCA+AJc5hPaYNoCYDOZo7rpmqAx
sBeKPcJH0Yn+8T5iviFVD/KKAQudhkapbEDBZc6E6kBptXRXi7jKSzhesXnBtqIq
uJ5Srz0wMvDY3NXbAXemoNIArJp79KL2IdXGTuG5W4YhcWdKwR2A0kynWL1vIWIG
GcPjSbtlGBZJ/29/rwgwtUvb5T/6CKbtYW1XcdcWmuTwOZrHt7h/b+mgcvMIsan9
BSFKir2GP7tQWrp/jqtxmxoxQ97gSHd0/o8dFfDCaQLp4ngGH7v6MxgCquI4N6cc
fqmOsvDiwTNGLKlIoKy5j/CVN8FQRcXfBfEVRq+5zElgT8S7HiiMJfzyUQCosD5j
O30k02QFqWwq5Df9+7V5i2qtevk3ZcXdjMwF13RtAEWQ8x6XLnIjVRxxBYRVHRxI
C8V5VarU+rZxXqy7yWronRVfx1NcLTQ3wKqrNvJRIwObLEPZSPagR8jM+weKrUQV
0wteJmIfzsZi/urTi/w31mLH9ALxgRNOSiBcL6I6IVLSZ69R+jKf4ZrA/iPgp13l
MFOM9L3eU7F6FPGp+dUQ7janq5Vl9F7xvml2ZxQfGx6M7vLtkjyFEODN4FBZmoqN
n4m3Qw2HtGeQCC/cEp0sLp2TUApVppExXQVKK+I4E77rf+Ej/Vltjng/N/9Udh6G
3QSE2eYo/mAOJ12hb7kzodxTd9VMINgE2xreCEvW7a34vJvJe9WzOuSVMDP7L2io
2szLcdItu7ACzbWn/A7fxHOfnELC7RNWSimGDUuH224CaRqxcbru8++mzac7h9vZ
9lpgSWfi/hPS5XocCHG7EDc+eLqgPyhqNz0TeQqdHW5RLka1p/3aQGVCXVOl9Ldu
CtXerCtflP5GAmaEX21bG5ZyDhT1m4kGbZkzWZZXAEbVjlbc6kLtouLqBOHIUBd8
zegriP12Fao4S8HYB93L4qlgxLMDqINKeYPcUUvBnJANMVh5PfxwelgIww5SxqvL
xIF9c5lEleFEkGRUe2GQ+i8JMdHgMiIX0QxH64vS2/rO9+snjZfhUykWeKQD0Kvu
v4pk5WcwUBXlofZgP+wQdnpP/bcS0EbvFLRGX83W3zSGgFMBs+MdLxvce5K9kqPY
z2UGdsJEXK+5lAB7lW8t8xAKp+lOklLT9EUnIh6ad2c5MqqBnkV/oUpP7kbqxn/y
F01Jr8Ul0kZct+1r+xZgBzVjLL4WryMXJh5V26eUy0xq4/6Wv4YJ2WignemfOvbd
zQJwGL62VYyrtuCL4XjzDoOSthuOonHzd19QNsDjVnh643+5U02/d2aa+Aw8KBfQ
ZbbZ68OXrvPQsuQ4RzuYmn0Hr5zEjfqVOR54fbYRGNF3uH3txGHDGbrXiCcQHEfs
Ps+5bQ3RrAOcSfImpq92LyQbStRaUmbJjn0QF7P+jrJDaeUSMfred+CHBXBGZLkM
TQxe6q1OoI99TXZinwrAAMOkeWLh12nCGnSpM1uW/PD0sgY4mzYFAlLbrHZCNefc
bFrmiojbbdgYXnvfPMm+hBLR1UwKe8BWhAkpxQ9lnLFCpTURtdOBvO0+qvRtg6Sl
njsIlJQui3V3Gp9Rf6zZDYrm5e8JpDm2ESIqhApjv0UYa8S7vMRoGt5Ugkebc6dg
Ici7BTz3wMSLoioKpZTbyEL2wyLdvpgjIf7MujVqUo3BeTrNUuRlXCczkWC1hU9N
a0ZkVkho33ZFERppSsl1XYcfqp84ypQnSoay8bbxLcLlg3fIF1p3qlznkv05K6Xx
w7n7KbjunjkESFOvIfHDUJzdkfuuUO/rN1Q4fliN1hq4cPV8Cvvg06Y2wbjU0lIJ
A4FnD0rFHZLLuPlr8YveTkIsYEt1ITDj3aaQsVKZDkNcisCUFOo77PMQuq/WlM7n
sSmpWx2QF22/QsHGDaCLmVHA3MRN5DVbToW2imnd8rhI+emEWYB1lVmuExko9JW1
e3+HUHWQtg9RjsfUd22kIx20iN8NGbg04jnoDUiT1J/CtyJb8OVCM7vx8SG6S+Z7
Fm3EKzsX0Q+GqotQvXTFIpisL4xiejK7Dw/ZWW3DUe8JU2jqVS0+j+fR8PqaQDfV
Dm6qN+0m/whPAAYrVAdcIEHqb8NMgNcim4pio8Ra0ww/7Ym0et38C9yVHjX/+e69
cCbY1Bhe7z7BthTFwOfY05W56mvB76aVhEMa/ydNCR4LRdke+ppAF7Cxdv9SYCwx
o/8n182gpBGDTyuM10ZXaH1eOJyMmgOHWfYEcHXyjTCVaIOWmIK+tBMivM4y27Q0
vf9uisUYqkwop2G5QUa32KSzWHcLpsCFl80bMe6MddJP/E2NgeFTSmSWrzTaemVl
hycubkpg5U9/6MHKENtVmifRHQdqrYiM/+WfNTTdv3HRGmcHwz5CKhORwBPK7Jen
qN1o6vl9/Yod0tgOJeD6wQ8nD3rERsuoaXBQ7zcB6mXsFrcjDX16dtM0qTWJ+BSE
dqtJrxLUOj6L8+fjJEAdaLEbsYYEmDKs0i4+lo1jK8dGgm73FmhZsPonTK8+eCAc
cav3gaN5iMGZFUnxUckLlHZUQir6lTqbyqo+QpYRfUeWYOsolCmDmABEzaHnEVZ7
v7UdDePITpHllbJsMaR22LE/Tx7qZxOx6jDeSNuUOdGzEbBRfb21RWi0Ybf8LjCA
ci5XVx3nGnKAQXjRBUXBjvsSsBhPXzyylEQP8ubCNmWZL/0LgjpTzwc0qRR+ezYb
a4uc8V1QumlslU6X8obgt+jE8FL5dq0t7kg6mOppJ1n5xWp9Llk72UHkahOZfrcs
9I94V6UWoQC6PB7ruDN5psI8YlHVEgy1xY+lxsOuhTUrCBM/Y2ImccitKH/Olb9r
SkAMc9vLGyx0tpOcivj951umLLUUXuMeHetJ5ilVEsgxCBluevumyhmGlxoGSHio
wzGEDvo6v1+5kyPEqIn/pJHpHotGgDbN1XbSdCjKGy+BT8PGRkMftXEe5N6lpuuG
Xst4X60os2Z/BoZcILyfid9CCdAjVIhQIBe7wnrbNwDn2+ikzgZrhap7N6f3LgTw
7fkIXsNQDVt5T7zOL+hveoqVnCiaCffkIjrRKyfYHYsy3l6MaAdk/KEW70dNUycr
i5t+Ebuw21Tn6q6sNVc11A8ojzNfbo+G0S4Z4lsSOHmulajbhX4SNrARHyBGJlj2
Xq41nEz+OKblHxyNjyEFGVLai0pQmK8I27m8D1KkVSZyhcgBq825qx+0P82RomKS
WRrD66Ckoy8oJD1tEvy03ekDXWYNMkB7uXtLZMPXOqyEj2eUZyGFHX4PehATzd6p
r8g3HXeotoZmj4WrgcrqLYLewNIQ6C+9kYtnTzgh5PGVJz+kSXPmNFyKp7Oqixgr
g6HyAvQPQLfSm/YMVAlHcypk5iVhSW4eMMUJBtaT74OVPhOImE/hRAaVG60ikv4L
AdApZOmdOYYkbmcbnvKA1NybDc/vTGRI2hb9ds7GKxWUOVkwXFwZPryTJEA/mHiv
KNTiDD4jkGiNoQev0qtV2mwiu4PjHyfDltwKcKCgW4SZqiSCsOBnjph136Fq3sxN
L2Wop91CeFv8r7JA8ny9RsNxNy8m42Jr80ZgzG920TTdBjimjWxTveBgvqMy5cbz
xABNMyR8CyQrEE9QyGgKAuoWzv6AjGtfBDiQVDpj4BBd47AHLXkFcHNdV36B0f77
FvI2Ouft2bF2FnXGdD8VJnB6XY0/L/xW5R8ezWEp1SADMS09oKbtbHuyZPa16VWq
ZFyF/Fbu/KO3LHRyd+OneL38kQ6MnLoB9B5j9j+DJ/pcFNO/xBj5fuVwiuM/bWV/
+mETgv9sjrC6xWJOTriqPmg2IbFHVTm4KpiP8MJZ0DrCE6mfLW1sC6NQFb4Kd3Qz
ek4f66OKxBWU9X9q7kpTyLZpmpPCeBq+KcUhI5tk9Cv65pQRQkUaj1kwqBh3GWAw
mbG26iK4SOSiNX9C+MGrf0JRlJXHKouxrYYYteBklK/3Qbnn0zKGdDoUlIodqbjE
ge8Wf+TTL+MzodD1IEeLkkHHNeqVq7Y/cUmhccSc7xPySwp9V1MDl2jBlsdpgF0O
x4VMc2Di3Bg7GKYw7924tvbwBMT3Xocan7YucUKRIsySHJYou7JiRqIWQhVjhlQq
myathoGppN0k8V1543nyhoZQYJXXBV0257oYBvxS3Si5zRYFM9vUJg+FibLwl1xo
nYmLpsMH1qHkbK/G8sLhKgeQBQ8NbmAQlSkzk6nTzZ4dIK/iH1NpSTwEiZmIOmV/
U46VONARGa3GlVQkExdStxMOWteMzinYnOiejUTGsXqei1cCQTHNhkUpwyMyj02+
d1dEJGPV5GDwNPx86WXw9VlKHUj7ILI7vms65/CjODhiRWyWWjoAKUbu2dXiAVlG
hCAbjwpgVpWQTddRcfz3jPRx9ehD7KKO6yu6kcLhPFB0tOKAkPP/J8/g1OrRydX8
svwifhiLviD5XYZKOPGkG6y0TohxruFSU2pDMZI2zKvY2aIP+T26bUiwzU562KYU
4eqMbuxAfxJxFfcCUDymPmV9XLcnXk+/sEu1ZRiEPu7cwUKjULhS0u4IxvTISLJz
4dWCeMng7VmQYsL3BT4bvV5MBq99/rrSKNcv3mJLXmOHQjrvHGGd6Fj8yqgDJtZ2
ZcVRMSul5wirIu1F9knKkYqBF+fq9CFHMHOtuA6Gq0zgbMx2Gq1rEuqy/9lJ4dd7
tIJ6ZbuFWBhT/mwSP3PxT4GK+TH/RYKYvgNfdmfvZ5gdHdYTGuwktyPT7HKdaNlM
gx/Day8tV50jN4Y+f4WqiMB+d1eteVngHn2A8xLqkGWi+W7t2a0ckEq2ndI7M0vr
i6it52jsYQDmJqGmLYsWPK1Lz+dMm6wnwuV/Kpc0QtWoMQ2nPr9omMgfYgfIan4R
bsmN/Y4ZSVWXzQp0rKD9YLvnotnxSU6w+E3+w2d3l8nAQQXsJa72tDqtiKtzAJEX
tSVAW8Pe93cIQblujWcpSU0XtvqgcspaM1IIHXBYJOzpSBT1E2rcVzZLjQjKmFvu
gjkEq1OnZS84qtQYI56CmQ/ihye+QPcKfvM6zFT/2PrDS3GFCyzJ01oOXCJHJ3Vz
1LYiV9WsNEoyPYQ+ZYO0vr7YiS2/pmn45drRFlqTc/qy2ToNVkpO758J6+fG9gw7
eEyS/A1QVo1mEgd+tgkPbtTDFH1tuFywvjUxpZF7Tngy8VCqlRlKmlD9zOmCGLHk
+QTSaK7vzyL6rhLYQOwIWrU84RJUP/M07sVJ/GLs8wMTKSh5U6TZWT1Mk5wmG1Qj
PmOknpzqXnx8sNaJWUnOIAsyF3tw2uEl0P97QvErrjZl6d3eZtpYbAtksJlY8hzA
PbQG1XffM3tD1H6oBYCj/lYhLKoq5FKF4ZlKQyT8EkhgB6NQH2t9uu8WxPb9vvcx
wXHYj2ykl3AgI3gMEqHEkvrAzhI+LM37pJqdlMUdYS5DWaFBm0w11u+6jSF5f632
Kh/zD5mNUd9xNvqblMERBybwXzNC88KnnQfkRuAROA/zPwQulmh6PsxKrXXN8dNk
6qe11eGeXvpLyAB79bSmCla9VJj3Weeuf+kr/KOBp7G2C6FwdeDvrbQ3iHOvrDz8
VJdewzIg/p2E/iHMqZgtnPQ8UqZRM5Jqh4h1NDRLw6HzR4+dqfZVQfkp3c5HVdWC
jV2C1xQLQ5sxB7tgEpGcYmp+yXasGZDa2Mx6Calb5OQAGwo6MJYuxBm/J3q2oOGP
03dz1N7YevFzlbY2QrjgVWo7/2UckAMqxi2WQpwD6Mx4InE8t5JHz4MECQuorkOH
9Ug7OGu705Stiz+jM3glo+tgBvkUtV+8yTdb3IaOGW7gZ/wlomEcGOJRUgRGS7OF
haIWl4OmTENHOKpjk13SL7rYlQ0Pgjmlnuh3T8IHDxiVo1Fwm0P3BB91//FiJbb1
i/n8z1dlK7fqt8V4gJFo15bfl6FG5BOXxwW02Hh38YVKAVr6K+bD44NgQ+Yx81oG
WzhCvYio5+tlMKpELZblkCpQdTRtmluHX112/BqXqz/rRuG0LkuUi6NbOEpdVOaI
T99jYd44XOdaEPqU8bJ/QjmmacZ/QECDlzjfiDVmEakxoGC+TELBnt6PXowSPcF5
8f9i8V/wykH+fZDcVLfm9TklMd3Z4aTuv0FcdJ0HodE2ieQLGmFk6GyI3IJlZblA
GkMxxRjvUPAnWHcxV1Juca/NhPDMKLGafxbD9pBejoqBaW1L1nvC1vtoJt4YzyaN
ZXbTMsl20af+1ev+F+N9rKhVKqaC5fefQSv345R7mOOzcnd3hR1vtqLrejT9OMUy
OcE3OmaqfFruURqtqh0Qt0jd7og5LZZcTE5sFwm5bgft8krrM4Wfjne2ajrDdPaw
biLta5GZsro47Jzw/gxYJndKfKGsl9TPeLQviMK+r4tc6ymp5cpGD7O5Qciq7vQk
xEkzYRUj4bJW3eA8psYl7G/dSx7Xg8d/69+1W3aKRT7PCEAAa7mowmpQrZKZzg7F
xG4s+Y44E8L8se6klGv1mV89xq7xjcThQbVSL2a/rJUrCTUnxTNhLaF8NMBE9vBa
QFgpBs4o9iGWJYrpALD/pqaQr47wYb4Bo43AnRtxS4X1NJDPt17soOVM32BdrXF4
Ejtk3l0m2PWoRKLuX/toJ6+4w8KDVu35KFIz46pUdAcS+On7Wq7PGJOadI3pzoJT
S8eSHk39GR+kmLZ+ypzCXLoWlLFD1fOCQlKQQpI/GopVxLSaQXNFafvLwg0w0FxB
ywrAzhndSSD7T7oInZuAJ0DgAuuVMCCLbjsQVl3q4jVTYF/NRhqgk2PUjzF4gvsf
YYHgBYDIJZDHV9a5POIzfho0BHC9ICo/bloWBuPx8dryH+1SBj4a/hSY/AZE0IPI
29ra0DRb7+A/f/FlIgEnWM+jVX1TltuTeitCiu+CnavWsmJZ1o0rPMAHZwkUjr+t
nMEY2jbb4b7f+FdOTrpoQ0kQSTuPWMUPt95+40PeTT1/FlGUoaN+a9vna+xKvcd8
SUXxcsQIX58bkt2uz4ECjMMvq8vCmjguhnJltguMBy5+b/qCF7o6SNOacYxpEKFh
zuYzrAOP1DFPzW/IIxEKhzgHPFHK/kzIwyt7uxxe6/h4Wd2PndZ1z42DmbVcITuE
aC7bhaF2x03+ExHhm2Q4h3gLuLBjbJAL+3Sw0vrM15nxfuSK3VQkXnXPOtTRD5pI
QHF7GBpsedOowUPkS0PnhVBpXZLeiY8jr8ihlTR69KsFKOEYB26iDesBVRgq3pTM
kjmWpb3MiLd98i0qXyu1zJSGKq3QyDpgDz+MUlyxUj5t2zE0ujfu36PkOKxki/VZ
hfgJB71RDYNjlxhzkoFK/h0xrxpkHs9BO/JlVDY0l7MjUeHpJTKF61iFgwyChP6Q
P3mq+vS+/TkaBnzcWjTEaLvUPUOLpdljBqXoMKVbJu+mFkAFZiK4PjBli4H/VNWi
FK4tiAFqCJT5tgJfMujCMIGJIAkY5dDMG9GivnELbuK73XcdXK+wgAZKO/yIL+Zx
x/k2Rs6kMr1vq7iZf36Q9NakUKtnBT/eFTYr81R121jVY10LX5oDvILq25tBuTOw
VdHpjL8AU1u3rRmT7GonIW0cRjpvLaCi2TT9ispNki67DhyWlNlgD1rJKNehIF26
y0Wnd73ppsI3G3gNmyp8EP6uXxF3tdj7xuEQwajGeXRLk0cKbnQ18fzfkmTyl8dK
71uI4MaTb2mWsoIdqaX5/U0nleHU1+KpvvPnZSIfSx9HDdtM5Vk5Bl2Z5uIg7IwY
e75ZVNVFHlJGKK18CEl69Yh9Ncdt+dBTUvJvyVmeqIqISt1lkwK+hJiEbArIJnh0
cUgp3lxO65myzbd/MQP8O5bBvY6hyfrEjbn5+AsfFgrPU+7/b0Ig5ERknojagbER
gLZzcCfza+UUXSudCj2uYHWp8EeTfLnpW8hRkQUvBrlM2X/qwjvhropgpNfofmn3
BTDtueBXm/xPyGL9Nfw6BuCE9XBCVjAblH0waDeHi9M7EhW8w010pLfKr4iPr4du
I1REVsIEY/xv6icw5p/Hg1Uic3dLRcwfJffJANzTQUz8mTuIynbwUoQDrfqMtVc9
QCiiuM06Z/lyncvRUGN3xM78nWPk+iCKXSkZaimeVSnimnlksrBX7VPV4OeiEPfg
1Z4KV+m1eDAyjKe779RxrPLXyu9BQgyFAtED1+C+DxozjYjQUJhU4QrooTDRVhc3
Z2VjQfyczGgifmYXY2Cqva3CjUPcH4jIIOmgzuJtoBqmBeujI2CzANUS/Gzd9Bop
owL//OnulPdJWk4Z8+nocHYkcz6RvIA6HnqtrGLz8h/WNBrjLLI+K8gw1CEg6mVb
wsW03dbHblzTRPWpA9vXDFKL2j2f6bLqaz4T4ua7ZVWjMjJj0KNtbo6d4LqcIR1A
+hNsgsQz9epc2xut73vVHUM/2zZfXfstwJ2JP1RaIqvX3J17VGDNB9bpADpVvYee
BJLyy2ZaeIyI6jKEII5gmWdopVHaLC+BmOtYN0sQqBhdi7kte5etlzryCkE78QbX
1lqCsG9HCLxHS+Sd+OYETSflsdFDWDFqHcxoMwjcgw9CyGZfGHOlXcQCTL81ePDX
uYL/xDrJDWMje6YEAS2PKuc4vDuw8V4gaqIdDw+2htypUjjwE8dGk1l0q0Eid5mt
+hmOAjHbkQK1ZDuzXd3Z4zdzEOEe4wXQMuBHa4SD/T/Ds+OWwjRVriGrhKpvsmRZ
P66WONHNAbJkcLdnHnPC59FB9lJ9cSlu1pqxfmwZGArHnsLYOlO+HSa5NXgYTWBa
/EjM7zvCVezWT66ioAjtIRkJAAUNjeymq71rAGCf/5N5dn6DnMcUqEjE3o4SqaM7
jfmO13w7AT0tRm207Z7hqZo7F4NvA2h0+jInwLN5U5VvKl5kyzOF5XfH2Dx0zsKM
M5rqiyMkAOdS+a7GMAPKnK57NssHZXj7BnlS1z5xbkKHwXnYcZLPVi4cciVSg1Rw
yEcK7locWm2/PZiHZMkBVkevs6jQQ5mb0lshmSTiqmyYq1mg1Ehd4PccOVXqC3Nq
++/yTRGmQI1fCVAsRwdFBPlr5eWN15IeFB535kVj19x32gp97vJadmjo8fnUMNmZ
pWcTgVkNTOYX1iv32dULew4smicA3sTqX4Wn756U7BhYp8e6oEL4No3ilHomxcgD
BZ3PVpSKfCeuciEh+RfL+31DQAXeHmuKAYW8s3LCfmv6uZOb8+2fpYOhHFi4sAb5
RaR063jmZADnNLSRmKeJiky3ji01tzXScigNexVAo0UK4GowIASKFNI6EfKUWss2
t9IxWVNpdzBf76qAlRGJGsNywe+2W/EUrSiMCz5TS3u2JnvxD019U02m996mb4wc
brLhYg3Y/zojtC25yHSQ/So+uo0Vysx+wEmA/ggP4XjSvNiY7i6G5VT8VQeUoFBn
YXLxJEjDhjsJE9d5JK7tvLw3BEa2eyE2MlAS8hJ0QHBmLago8Z4OFN2VANnqyOH2
LxJDhwdsi04c87wms/aO9Uw0D+KR1C8AVYsqkcuNQSj9uGQcbWSub43LHant33RF
NGEK3cvzStg8Uqs5c1w2qbIDsT++OQPHdWtBND50e/73awKynsXehOLyORhk/3Rd
OTrg7YmJz+4Xr3KXNnzQPY8u/6YaLJoBP0aUiKVgYkbH+NrFBh5LEB9UXBtINP4D
2I1ZacYJ025Rc+lP3KYWVCuIr2aoH1IUpapnp/DAIfdOC1Pgi5VDWMuMDG9UmHX6
A7qlzW6S25YbEHsT8ssJrAWIzXvV4AF8fPcYtpVNjOY9jy1mbX1ibU/QArcrpRvg
pLPcPZhlRUf7mPjAwZJPo1aFL5eMh3qtQZaw7za1N1gcBJhPWkh7XCsXbbuYWWKJ
4heM6q4w/1tmmbwtc3jRG4mf9t450L+7O5ZQdDdP9rUAHR5rgDKadPvRBivypand
3soAUaTickNx4VguLjeQmtXcPbCQnA6LRl+BSPAw3Jwh1XE6GPWAMsQZGWourD1k
AXUIdpoTPUhCzZ2i6ajvdfQ3qz1W0DY1uTPMVGR+g9aB15YLBDk0MsGZzXsxb7gu
0yaAQvr7AuY1IkvoTiG3a5STm587jhrOvQ00CRKGbUdCjvoUgVqzal2JvOORHX6n
YulmclUD0VH7LLPtV3Th97CneCWU930Dc8G2CwBr0PGLDguBfr058Zs/R29YCHQe
yiK2WORe0puYdKtChNIp8CNJ19IJUTCklu5J2Ui12b+DM7bxlQVLnL6lFdrdKo7D
VSKjVnB+tsuftqQ9ctk6vmaJE2t90DLJpH4aRn2sA8t++ucyXlgPaiYDHuahLalX
fogsaSwhN+nykN0sPBPIoFtQQ3SZooygc1AhTXGOECyBtVIded1pjeGN8d9DTuWk
lO87meumUbPB+b3lszsZKxwCH0YVYg+39DX9KoPdG/JpHCeaZV5PWd21xorfhOTi
w18FhHx/HlaSuwMEnbgTWkoQkpa9b+F+3isoJXuo+IwGUHOgGKsCw3e647uyNlXH
fH2KpI14cLsHN1ckZUbE1pMCgZ/0QmGAcIwA/FhbaRGY4D54agJ6TjXK3jZB4YZt
4vfBOJ/D2HtRxher9H5EZ1m/Y46NpDIspI8Xr+T2A6QR7ZX0swMdcWlb2GiWLGzY
EgwhHfM0C5DwDHo2ZmhKdRNhV2NeTlCOlw/OzcxocD/Vx+jo16dE/WfwaF6V1BFt
XQMSvZeXjzlJu4tc5tGGGPXxUm9LKnPmc9pI60B50ZoOS6QZni39H0se9gwfk/OM
nMLddlgiLxxMd6Roeqazv3FP+8VVtrU1avAcjUJFgZjivmWj+hZsIZqMR2EoVJh6
5JGbnWKrMlMJlKFkv3k9dKhuIiao30UY97/P7PGEixSEkFg2+zf1iPAJoK2gwBwA
JvLZfH79cQPdejk0GVyRyj8rKXByspWWUOo/uHNvn96Ha5bQDjatVYJ1M099GL0N
Zujj28Ms3cgeWf2Gr2tsIwZt8ehRvVs8W4A+LHtC/3uKGGfVKNxfX6is5+v4m5ch
+LuySGrqwWlBVGz8Kd9ZFXXZeJvFWmvlPYm8nF/rUln76NTY566Gn/OwDXYm9Jzk
yAq4youztISeXwMfuvUC4ldX8EhlrNeZp8MxereB++RNJDTxlS+F3fkzAHJlOu+J
LV8Ug7Cafe34J3fdah5FMAhXPPNM+J0Ny86I/k83xun9jqea3IUtZldxr8uYNZdV
xjX8sEESzZQlVMuEx86Gsk8FvVXxl/t6ZSQ+kAJwRx4RhQ4uL71ZB1ZvBZ5yN4yw
iTrl1Hn7mKCxH4Jg3j57oZtsLiguomGE8X6oO5qqsSQDH+ij4Tkh7XKo8zowG5dM
gLSKhzN4zfKEo2gr7EDgRrXdW4pbZsJ6IXfn1VET7gXq2eTMQxKetuPJXcQMWdIb
ntTuGP3tDp966kYNrzL6Q/4dR2qnhGf5yPpJmRZ4QJuHt9SPbZpjyr0mZb4EYpUM
f1GZS+BW7HoXit7lZ8B8fUK7SRmqRn716G8lTb/+qU2Ag6Uhfykpk8YfI0h4WzQ9
Ev1xVZ3W2inMAWo1nlHdjSIgvbwil32v4bp6YBFJNU26LhhPtIwiytJWyWjpMrDm
xqkxZy2s6C0dmSMBTqii1fK2VmUxsH9S3pRXR+sH/e13953nIJHgKqL6kP//4ndL
0S0uFILAz3U4dDfyWbNQI4xiBNSSOC8NS4i3MFoliHsXewtwNWTDMaI0tVvLz6en
4gX6P6zVIWNWLf/4Z2b0/dnFV6k6VoKJsVT3YzTEkfUnhW8jg2vTZktGvPHc+aPk
r2HC/Gy960mEbBohlPx7KB+w/dgPEcDA7AIE1sEudph57Lv/ubtR+xM9SXNqfoCg
HC+uwxyNtw016XnIKHHozO9i2/OZ9QC3biWU1VHT2Vi3VAXfblQ/QQoiNxDA1+A9
o2SeNy9QJwKGAGdzvaY54IavrRUPVV9JKe8Fw0IzUSnEAEbg/IWCrj6xPpXAE7BK
9DT7xTrJJ/1wTSy0j8RaVbtqbkcgsT5ZTFwQKv7LaxcbEx2rv1OIkNxAIb5GHQDj
4+HlSODwpAylOO/tZ9Kp+TaCA0TucCbP8/EHBjSO94nmpnvxVmAtsg3VYwzCDi+n
251c57UfrxX2qXsdSO47GOhB1gMJ9WiigJKK9saLaJIUpN4w92VBbqzWTytSek0j
ya6Y5bu1qRgAYWAKRPQyBzUnpUaZuHT3UNf5mROO1zNl8JwZoo6VJ9REDhPLvf8g
3L8UqtYAYGUZWVQgexUctXuzSDQ034nNXXFMnE2DYwe2v5PldSIbzphocVeAPjEp
PlhJCAmH1M4UD1lwPgtBJa/rGAAutTFoKQYPyNwOv+iy5s3cpyYy6RApVzXBGZl1
0rWi8hbfDt3NadHbwh4WXVtjDX1Ggi0fUqU4CkJN8hyDA3sx/n7mjfCaTGhAK9/f
Tk9yJCdVZQ0dEpYfynLAFlgdZUEbOibTb827/rxRBn4zHyyeWilz8wmH1iBkGSP4
zFawUgUix7xXMWBouPe+fmFuQ/QcyQyHnMcC1/F/Dr6pREZ9x9DibN2RisgMhhQ1
j663R2swsi6PdXxNEc/+SLf9Mx/HtVrWXUTJHjFBLja2z4HkpvZXCwSiXgpkkB1u
ilhMgGHGAWnFSOSzy2RFTskMn1b/zSzzTNCVPlEFTJTuD5akzu79swIuAHM7UsD/
9Jyku+xMMXtlxDhlGCaNHWVe6MUF42hDvxBMhoNjly0cyFoL77B2hav0+gtY+HxN
nSiccM1F0lMqRvKcRQe383+G880SZ2k6Ywu2COOUYX+D6YJBoR9ZgcY715b7cvBF
a7qGmeMUB9nnPNEZ3agxrWkMWYwEGWwUsASqarvfwLtDGSZ/O3VkAuQlVTajqTvp
bZ7HpCufHO74bsz4ix9BiwA0Iu+qOeuMS6KezKYUk/FVDNE0O0CyYYbcsnSq4mJ0
D4qDk6Mqh0U+WNrRGQmbKUKwCjk75e0bmVklfOfmgcNAiN1YckOaIvHf63CNZ1qL
hj5skOluVhvLuzZnks6MryHUcw5/FV9Fn4ZSOR6NRx+VtMbe8Q+OyOktv0SeMNzD
OP+05Wt4u9E6F+bbPf+9hsM3cBQC9ZkL3dTe5tNDYJFFJPz+5QyQaX4CmR56/2pO
Y9Fuyd+A1Ss3wLdx8rwOHzgnrioNxBiMRQgBMyBnAnBbmVK6lR7TaVlxSdbfp8i3
uy1boX1APb5cj977LQTlxk3dAiWD8TTdUPAOCN0c0B/yC9UEY/l8FiE0DFbd88Hh
DnKNbxLP0ykKMUKoMr/K8IIgMN3yzm8SAJENC6qX1YvHaSbIQLYDb8Xjo7wEs/KT
NP5DObA1OCwKKBZEF561tLvthAGW3bIChL9HhF4Q/ZVwPI2Cus4SnxeQZrQFgfGk
+/lEmGL1N5TVCme2pZfO+BqYzB6Ia/Sbcw8gG3Us+mYtu9/k3Xop3oRWib1TnZBB
wscwW3bMgOr8VIq/E8jdcqx+pvluSJ/K1xabuVlGa4UOibslMbJKUZeXrFFNXVAe
RPDltpgjtIlcQtPCC3zmTv01tilN0R5ZmEP1ZVvRp1qO5x3TlfjH7zuUMDE0wNFB
eHkSkWkVsEEXtZaWyDlDzomhDKwUonIjVaZN0tSGVfcDtQ22557Xe3cZj0Kbp8sS
/U57ic7Mz5JX5HdPHSTanhVbN53EtzDVIc6cP/WBfstoIecy33NRZLDywvTXoaF2
Mf+cRwAxxGwKTZlm/UKEd096h7+LkbBOvsz9vCX749krx9dLMQWyYhqttu2D3Rjs
2fxIceUkCK1wq8tUMotRC70pfxT7Ryx2lLop//xJXO+WNQ9S6uiOezJLvq+npJSS
CMxhQ+0cZUIW37d/039uOBCsqsJyyQ7LkSBffIL6qotLKAeGMumddtZMoxhh+TPv
C6hrKb70n8Ec+rsP30eULoJ69eH9gXY2sX9Jk67hkHADWqfiqybdG2p7wxnErmpF
tNe5oo9qemuqqB5L6STcaUyt5SQd8NmtQs24r8UCZMUKiyroWl/P6LNorru5sXvv
qDymtxGTvGK0qiuugRCr/u3l+wRliXT7M/FU5QBHwIv8sIw8/hlG6uDU4FmHsBVJ
V8j1TMYrxShQz+jlQmG8CwaK+y7Rwd4caxPr1GxpOtY/lodwz5taoQBDB8ZcDqFp
ufj6XMh8eV+dSKyRsr0ISQLbpbqL0oOT2gU34zrq0AUTRIb9nfIIti7sIcX+JxIr
O6tyqSJux92hVOKSVcT2BWyA/2zG20CNzUtUWa25i6DQ7+mUp4yUUtOqCR9QeUiu
FpmcTOHNOsdemKnMJRG5ahv5AeAAd/UGf8jNZdTVVSrcfkxAMeQUCruzvN+IoZMj
7FO2jDNKSu/niukqZeXYt6YbFANT6XSwqa32Qg2MwXLviJMhZTCuSCcAF5fxeZPZ
zIrJElqlloJ6I0/h6oDFhH05fGtYBIsrIdBE027V40EcaSNRwTIOHvbsanD7QK6j
zJit2rJSjQRGYyEuA4DqFTBdsFyL5nypzREwV7qSmZFmYnUFcRoBhb5ii44cb2P9
WfgFLQDNefLC3k/W5MlE67Eio9QuALPJqkz1kTIxmOsBI27qRGVNjaPNuJuGhARC
A3y48wrqddKPj3fi+4JflOGFiPd9qz6742T2g9CeGdqeLYQ6jWHLVTN/mC8fLXEM
EGoWYw9XI1rGRUIuGcB02PR8ni+4p858rfd2Eds4W498gV5TMv6C/yvXQu5ELiTo
Eapj3z+dODOSgUGrVkWWkffSEkII6D+1WewvlysT1M0VPhrNdt1wOY0+valWgiUq
a/JgvmJRNRU7yJIzLnF2W3shcPMuN1aOXQg2J6y05FmKVatUCmkErRBBs0tFw9X5
dL5Msj2hOfS5aBYR1fttE5AeGs1C6TNUPjYd5mG68TLC4wMgJJWAavYuhdQJPHcv
ZCtpzagc0BLUD5rNu3vK4eXm6RYlyhC3NyQL3p7tXIj0281aFQWzIBA939yraZH9
iVoZXKTzkj5yVdXxSSJsuONufYxdGXkJkZb6gGy4FMH42tVJFdVINz5fX3xqMLjL
OzdzAKFyyuuu/si1ypR4dAvrXxAM3KZMZ2cR4gCn7C5CR20/DQXuOL9kLwmPmK7D
N+HmMXg75pmnHnITbyUPwYPzpYaNV+HaHQYRk75Ta9MfgIdZ9b5tnOe5Cv44ZEw+
/GUrRV7vjVZPh5bp1FfmXYwBjLO38TRjRmkJ4an3jr5uIEfSqG7gXEn7zaWud17b
A1ZtJg3KlhY86aZ0VFUewfyAPosGXpHKHg+eEKMbhE2X1u/pJVkL++Bo/Qof1u1G
bhGbFCq44pqy9shuStRCB39x16DCdZ3/5qi3jJH19iIqhx2Lb9exdaOWrbPc3VxO
TXoNrGIjRzS+9HY/qc74u1EagN7v0jSrP6IQhDmyYmTOwoRXi4rdGfCVBagn5jYX
vre0XQ8mWpVaaHp4UO4WxYIvH8RsAxHkDUtuTWptLrwnQF6e5uk3yMyGJPOKuWGA
e9+2uXGgML0qaf7/z9PpFviNyUwNphQKpY0msdM2R6YndoiKQr5NsQV7My6OFujg
SN13x/ovr3b3vijnJRevXYyJJXTNPQebzM2a9xFdDzDZDuh3DJGf/C1YrJz8BXTI
y2ReaMVReEQJbpzo9Yqu9KMXbe2my6fyZEnGSTZ/AzLes/p+tlwoIXTYt8qRmc27
gXTAhXCLSqMyGQleLOFMAV7aqUi2iHgqbm6ChhjVQoHkdVfVXY+nyjqaO0IFWPTH
ziuyJQ1qRJuFlg7PEQpZssfntg+A15JO5VsU7WukINjZh4RgWTXsC+iT1h0qv4/N
TlDezgudIvtLVZo9l48WvHsPwChp8wUHeaDGS3NOunm+qwynD6aWJRMSCAvkhcJd
1FCx8wK9DozXPjE9sNEJT4kjckwXxNhWSN0NAxUARzoYVzbTIfKtqFwBcrW7OUMd
tVv9xe0uM0fhhzpssIkLgLew1qSTrlUjiMdZazjAdtLYSvKtWkZKJIyZz2zZNyUa
r8BJdi9nGaQDGesI2oRJhNGb4eS10fwDDO4n63Uep2bgAceTCzeJO34REoLyyjV9
hO67Ao9g0j0MMBLs4sbe0DG2ppR1KJDm/OVgPmxPcLJjw35ehuftJVVW02dHHiZJ
mLuGLn8GeYaUwcoW6PuiNqNo4l5x6pRlwoKQ7VXV9V5g6p10FdfHJ6553HCq0y2d
4ZJbqjAIK7YfHA2eq5XIwdzjy/aTOkwXatPZr2qX8GEKi8RqrL8uyg/qbbWMcgZr
ZmeUdpPMl9JEGStzf+4+j8ImA0oeEdUi4mBaDmbHRaFWJ2LAQuJh73/+Vc8shAjF
H9wAlmYc7nARGbGDEwLjrQVwFakjbADTkJ/Y8K5XOJ2EcckekVLY2wMcyr+JfAz+
sATUSX1hH+RwnDqJwVC652eRgskk1Z1fYolIV0XXbnUVWvtdWHDQiDQEteH00Yf5
nUtQ1F7LURpO5ksv87CKj+mMsq5DyNZUngA6W1d7xVGnygz4oHtUTg7zsayR7Wl9
T2yxEIl7ornNdTRUI1o31CXoDU6DG+FVQi34T3PuelzKra3ejsH90Ka7Cy0CHtJb
9aCAiA3VjI6Q/niRjtTUfcXmrDAyCUBeZyUr/ILD8/B+5sp/riJp+DDbdHtjlwND
6nNHE0vyDPjhUPd5ROuuOr34LM+sOxBfLExaAnRpG3HGiwJOFxTUVGl481jZWmxd
ZfPWSSoo8lbPE6fW0MuHal1YHQpDIm97srlctya/WEz/h46gPvJZu+wDa0OSiQ1x
Jnn0CzaWgqFjxUF/VA7z2BhfQBogxmp9mZpxeyHAThQbvXLb+kMCfqHphU9R8XBE
kCRba0hsrJ0Jdok5NZUdETnuZFp4TBtD6hEdIjfYrAHBWapKuQDEcdgz04z7ap3f
43Bx+ACexnqJ+s9zSh68wZYroo5BrY789DuGYkGqk4ETs7qzp76MjfV6z6Y4GaaI
vjZtM8oDbKdmXCR+QEoKufavy1HMxH97gVxlhc9TBj7BZQCX+udJSmEG0btp7EaU
MUQpMPmeAKYmDyTdantz4bUqnop9OJpHI3+Zi79dA+qWQ1CpVs6ajcC7bktJ4K1t
iRsS+rro+G56etc19kMgDn50CrhZ4UeMEYzEed15wtVEJ5ZEfEq3A6vUF/uPrKlE
kXI+qqFtnXYh8T5ak5YzQM48c4TyFWZMFyCQK1hRhOCojj+7EVVoN9NN9D0U/v9X
sdr1pX+3h2EGffDmXfQJ+8hTInrARHG09HbAM2P2AZVCPxAQ6UpdBQiD6LJ/AWcq
VELe6pWrpoyrdbUfSFo4/+gf627sCA4ys9FaXFeEzGPNV+mwKHNAM++xMxdPg5zr
8tOAvCCI64QIdxzk9GTHoHwQUTG5CS1gB8t/fKu78J8rlrZWC5S6qWUceiE7gP31
/lcJPc46t9h6SUL4xij3skuOqo8swGaVTQo67hf9ngzXcp40Ii3ZsJBDQ9XSwls9
Lg/0jN0TZ3R2x34+IY2iAKahOWIFxddAJRXXOcmcAR98plQmHbL5cy0EoXxTib94
SPp6IZK02lxorXY8lUywqv70yFlaf3eIX4CVdITRwADlw8u0YUBXUHzI1VHIf1kj
xm9AEgFytptIXGadWffH+PsFi3psUTUlBYKEhvLoSFxIbrxO+WIrWa5HUhSUEnJd
dJyShID+u9biN+0pMQShAkgy5ARt2J6/DBmBMnX2NawI5rN7sqOiB8978kPXSe8T
G6zSUadkLMHNLnLB6t7pERmdbt5TyUzLauQVb7M/ag/iAzhveMxM8lmT+6vJLSdC
J5j43KMgRW3wwQLhkpCCWv+smlXVyWkH9nupcfHJZCOyEvwunYa1ee/p0/q75l3u
XSCCyRtdnh7pJPg1rPc3M7MYvDW8fyeYCo/JjUl9TR2e96BuOZNyedAe6r36I1aD
ymQQ4fFrka+zeBm7/QgDizulVCcj27hSKwdrT7g8jmot95zi6cxeJGHOjfxXvff1
03WIfd9i14FRBDspGvRtZbZki5Bpd4WWUkL4412YLoYcudeSQEqkh44w8VsaL3EC
hVWnMr2aCVQn4OLGRwpPg38TsKOuzsy/NLsuWyMfGa4GU7HNaNo7ERtwGg7c+jia
s9X2kliUjNGv50DT22L2n5cRGSQ6hFeo6x/3uHkzMXVCOrAmmgABJHzlomg2BMrg
shqJoJz4cWUExNgGXkFdaoNm8M4X2i+5J4P19VsziGKW+TGSWzi3S5bEerRnEP2h
OlFyQcKRdbiM7qcLR88M1M9Xbrn6fjIV9yWr8wAil63Fo7XHpL0Im1XBeJuhRMSJ
nqm6U3reccgQlR7BxGRj+46xwdIifr5hH6mUuyUZ3Cz6egx5oXlx/I3+PNhH7ZUs
6baypyRZ6APe9xuPtHWtfMLrPZZqRUjDN5lRkiW3uOnlpD6Sk4ZU+oMSv+ow0Y83
/NcFvzM6yQdmF3L205xAJB/c+Fos/IC30SaTWBKS+98pjZPsApg1ZL+ye/St0kwj
JqhwNC6BZFgQguuHUXY0m+g/y0+4JGDHR5Frzw2vQhcCV5UjJmSoUR45ZlG2AV+a
7eZXICSHQNU8DsKjscJ41a6uC+msaVR5mUlfAWUUk8ee0e+Ko/CXmW9NErFJcZPW
JKu/owhXAPVT2x6ZgggaDLDjjF8TdvisG2DlTsxCdARao52hObvIe+TyfXdT/17y
Lr9Sz5LLwkW4f3tot4McNzFns/Co13B4C1HHQW/N2vXMmhg5/k8aPgTpiT7UGPpk
macackEyjikPteTXDQ7f1YDDMf30Cqu/RWTK4xRJ37+F8PXqLH+/gjulT4SQGmQk
aRiP4ZLRnZJ3RjOscI5RYQ20bpPCUFQS5UXGceeEgQLA9w9cO6eBiyASyJdPyzAl
B9AL3Rfw7+qkw9UDAOTP7/IUKsAGgfSK+wMROtWV44Yq46qQ8LoNZ8z0AVhX9W+a
zNjjtD8g0woW6srSqOu7jMWMBgvtnvlnHj+hrSbZXIIPVwE06Hjg88wdpp1i6DJr
0vScT5HeQXWZJPAmNxjnNw7Evmc0M9Wlw0MBpQnXKXnHvSys3Q55O0GyEmEFzgUr
dLnBPkLHl8B6mTbJlYnv/E8A7GAVDLYGwfFfnEO7WFcC5VnpuTEFanylTT9z0hcR
D3onYhANfToAeSLS09mDM0+M/JVHXOUcxcehgNbGLb4vKQSEj8Lgtc9BUN6pa5Lk
smdyB7eilwdyxefZj/AFGWLHBarKH600GMfCtHGJ+1et819HFfU9TNpXdFuVtno7
5BoILXFnrriPn+qjEFsIVtOBg/fEiV87yAuPbYQL5zM44Y+e5dywxsw24EDh9Cf8
xl3ICuFFbHd8q6gXleL1OpOghBH11Qf7uOoF9rHrgSOVKkyVm2Or8O5sI0IyaA3J
539LIntBIq2zqap4RYA/ZCZf83sqzYyjPQlCNJr7EMapaMezHCT3LJ8BAVjEzgpY
U2jg/OHpxLUwtGfMQzUDG22Wn9TWjlavBF+4Sky3E1asAlOzhGjjXLTo3btErOJv
DmaZacIoHXP9JgZpCarKSqz2yZLK0N1cVCUgunjYkSXd65qSBdSMOBtajZg4t+B3
dhIYOJG6TzRPqOEVwv6yhHNHblXG7rDsFC3Jh/Q0LDGAx8V2oHa979dZkCbkAvQA
8zYVwyXmHBM9gWDwX3qTKgKK2Gvzev+eav2Z5V1G1UM0lNBh1Q2jZbNmqcVfoGQw
PDPG+WtQHC/pWLTWd3rIKAFb/AIfC/9xMuKRStJE355X8M3hrJoj4jCJNZOS1xBP
4UfT5sJ14qg1nvLM3ftiundHCe4X+LfukzpjJ9jnP0LTSf+RnoXFkNKgylJCOesF
PiJVeUGX1ZSBrPSVC8wZZCrwnG7TIMOOsF2bZtxzFCS7+RooWbin0VItk0B9fKou
LRMwqiWrueDq1oMSlWVuWo0UW9csMPsSwmuNh2CG1bJ94S1HdExIN0yJoSxVwR7C
GyMVxUKG7n84Chz6SalKPpcmBPC/pXctQi08ngr3fZaKgiQ3gcoskIxX40cLrw01
3R1ZEi7Y6SXQM+wz9nZqwt70wg3xUocPPPduKfGj/CGdFmS3x9GsD7m15AUu6Gvd
vO4Dnf5QpH8/mzHswXKbUVt5mzxUFtt8MO0E0tFZokR7u0mnGPZNUvXfTYze+gB3
ITWCddiMOIGN/7KCQlLKJedywb6KflrYD/ho1WDeSEMSXqOtR+OD+cz5KTJjYK3Y
Mg1a/j7oKadpog4VsYApZiepRAaQs8GSWJ7DiadeYK0RvWIMsLt/mIBW2Zc0Lb7l
bVtbUNLoV5oWno8udZ+jVVbvEALmSRL3pFGkRq9OLsmZipTDB4qxXfyw6MO93BTS
S5SsldzJBDwCTBuL0H4OWChM5+LDBLS8xYPHUOOBjXu1hc2hcmChF1ym5IwUwhAA
vHNV1oHqpfGmtKeB0CjxYa3KHUCjuOMwF24muj2+Qjp/EhK4g7mWXewMbLqOPzc1
xKvJuvZXcKO2hwTkAS8y/zrkqvDOcgVqqVoCVt5pYTJYbxE75RmBUbzJlvPk5n+g
VlmysKZ8f/G3bkd4l6goY9fDmDLZKi6PPjUljqDCR/RadQdHeAohUyEDR+ToGqqe
0umS8+Hesa6SVufhEZ1oRoMOoRMfSNoM72TgQx4gONpZrF5d2DcbNcg6ZPNSm289
Czacx8BI0SK65dC7iF4htfTd45fz757TzYTgDqtynE7z0Lq/5O1BCr6hHSIoyYXM
vM/mcLzw3zW81VH7Oh/UUUYwNKwW+eDyagjUFfqiby2G9UYzqXs09VHdtCf2fM1Q
/PXWB5kMc4wDEmv8d2BoV/ngicOdM52XCasKRcsRAG7lStTNGoi/SIiBh9IfFK8N
z/h+S8rffC3YnHTIvEX7PUAr6rFVkr0syCOXu2/ilp/mEPUQdMp7k0nhrpgn/yiW
wNuO2IqLvqOpWil5AVAEyN/J0ewfxuzosOic5wdP2RkjO8xIx/uEAqmRujpjj1YK
eKTFkKJS170uEpsSAttGFt8ZPPwUi79GYOEvDwExKgBncYlVT9eLQEn3GQT3KS0/
Y5EjvH4WneorCcX/n+2HjS6MD8ouzF+EWLMkh8GTi77RktJQxLjvn2tvboXmMdDR
hYhW8h5M5y+WWlFedn/i13Nqltb/10Gov9cGqTA8GHchWRg55Q53JGyei1RO9srX
Uc8yM4GtulDxINs/x7iO+BNKypZewJUKHjgVQMsmwa2GSKgYDINIPA5IqvZvMUdD
htk0WB0GcpjITniBeSKJ2xrHGmV2zxUdUhKveTLVG9Kuo+Xml5e0j0puWbJ8ieqY
WN5NPTVTpfkU/76ALpUKQT3VbHWK2nU6vw+hTKG+pdtYjezupNgOmgl98XvrFlj2
p0FhPx3QgOs+DqVttZoEJpvzJbV6WIkut9YXKq9XSjHEQUfCs8dtsl7+3r6nQ+SK
OafdRjyKebsIbyOA7rus0sZW46BsCUv+HcaK/tIBl84gJQ4HUMMmoLO4dJsraj5N
MczdrcsaCTEEmRuHd/zP1ZS/Nfy7fNLeM0OL6nEPLMoRR8476kWyru3akajk8bTp
YAkXkTGfbY/IWV9G9cFd7++eb5QOzuiFm/PMo3wKO9RjoLcLqIvhJTMK/RgA/DnQ
IBDVze1mIOxTVMIDzMcXsBWG0oY0jCXHYi9fqd1JlTiSke9CKQVEvNlyIjCUnSCD
nZaVAepjou+2lDpdR061ZK8ZjKhKi1d/SYA868A7f8hv+uoqtkuWIh1uI1ikRE6Q
ZgorSolDKfYHLD6LCR3O26S25cJc/ABQ0Kh2l2RgRhn619dEQSJmKpwBQmsy1+Wz
Pb3NXk9yD3DDF2Y2PsdMmgZcmTMFqu6rOU4W+0hc9CeBt6Qsa1jFyYmzyxgBcj5K
XHyT3SXFfd1sJcKpB0eKZklcqsvo57RGMr4pQ7CX3Tbg6vGe5h4pCUIP9pCT9IQl
l5QjHZzpN2rxQvxptUGr4Lxoir14RFb+D8STltJfz32/bwAKQYehWHjxXprJz3LS
wiCmLslN1/CEwzit/eYGpWangXvFTbhM3B9L/B1Xc2kuzgoNM9A7WAbg235qKQ6G
Ur4t+Etq/vN6/RGDhD/JnlJnMToZRimFHcWxiX5hYazUSIKuXlWmbm+g8PnRwhUK
xVwllWbh3k1AV2cZFlSdL2z34vojhpEiLPuOGFny6A6q8zEhDj5CIeoUSHk7CGuX
qn0rg7VT6Ps8WzsjHqMhO2sPeYP5YtI3mc8TFL3XB9fBEZKyJslfDvpfM3+PfAG8
ftAO1YkPMRyhkp9/hlqX3s7qyPoQzyvxsR8SnhZ7BAtYrypjyzUv0WMx+46XU5d2
NjJ2MBN1YfcuXB77y2jWPiTThfawYQxA+EAyPksaaEx+8Xdj1DeDy4zHtS8FeZDq
ollZj5UdlT9+ktjO/tOIhBKQKc81Tow7YJvv3VTZP8WHiTMs6xINJALhbt0YSfhZ
+e4owJ1ru03HZdaORyugy8UuxeIketut6hlBJ2j1w5bnYWI8wk6tOmdwcnBQFI1g
1koyfLsFAHkgAkJCgltKiM6oyQLxt9wy5C7bdzYsV3ua6TM0+/O5DwbDvNneBg2V
6C0fCqVWve59Ackov9Zny/oLx8VkCLkgHqLZC/J1//dnO/H1u375waQ7iQK2ZkRN
Sq4dcIog6kMKYdwqqoJvfrNXy9+ued/DGZi37tg3AFXoyTg+mcUgRcCX6ZxpqG0T
wsSQuomRsyXxYu/hm6ZAtq+FJB8n47Yq/n3g1m/7IiSdg4Xi7ReteNMH28cxaDyY
GtXfs6HPO9Nd+gGS2QmZtZs9dLZP76o4Pib+z6DBp+8CtrE5Fm9M5NF4eD+USNJ+
kaKtG8bmXcgXON4+NtDQ8EPIBExJ8cM4ezQ3p3m8K+k4JcBi1Dpk4mr3ZRt3QRVz
MI35CjvHxAoQLkn4jEQ3vu+fVvP3R6Zu7a5dO5zncPcEua96GlDZnadS8QzgR0Ie
/X5GqN1TvLrziU2uT8PGlTim/KjhTZ5Cv1p7bhoVrlGmlpI2L+BKEGR/9spu+a8V
Ezh2a+AQFOil7meveNxQH64b8jExqzy4Jg9bqKUHHRU8J9fKx1hF42HDQ6N7Q4F2
2yT/PzHUkx2zdMyOHey0skXjS8gjF8CcTrId8Z+z2JCrdL7eaiBw3nlnswBxqz4E
xGKg7NIzE5ggywTIP88qgrK0R2a8l74LQDAQOdGmkHS24AhkTk2hDjzaV8U2jqpd
ZVqKvWgCvwPB3JL+aWfqlNCBXhNP3onoyimXH5PVhz7Iy5ifxV3WduMAZor1bPns
yFlzzCxjmFY9qg6Cc5LomxerT+FPV5fTPEBLZeRtFY4RGEOUj2Es6Uh43kUA1zyX
RBbWnzCyuFV3HZ2nsNtBRFJ21izv1XBOW196A+RMXZUBtYEksg/Ch98xeA645qz/
wapjQDH4SaPCWNTBf5oMytTgwu2c7VfBXkeRJK9ZURdmgmuua3O6m3qejSCx8lFR
+wN1NKWIyaEuI1QYBZ2UPWaF9LFxX12QnW22ytqV9mHctoJuyNugJ+W1I1A5u0G8
Gu1HrCgDFHCve4BamI0qdhhb68s8+DcN7ZkVuRlBtvOWIjT1uCpHp63UWdYRJE1Y
YnoqFreUjPTjDHcOeYWTR73jcGaKXfZiNMRp6aAaXgGF/ifRtKLQ7U1Y+ud/yjcR
OTzZOB4kSGPCp8IQVIeaXh+FkZlnHIbz0Rxvvgo3Gp387LRK+u3huUd+n+VI7+kF
CC+jw8yty3dFtY9zLh/IcAUV1C4eXUryBv48bWEJaXVq4UGCCvMY1g0c3mDikTw0
pkIPHZ24gJp9f2YIjfONhBeg7dt5RK0Aasw3tFQPUbpBZKTBJWJUQEY52Gqjwv2Y
EEJKXEeTqrJICeufJNOptCHKM0RcmaRlDENFMfKv8cdJzPflm727r38/V9Z11T1X
kX2UOct/IUF3Dp+5oTLoDVBvMaK4oEoqUEptXY4qPdWmtQHGKt1YYruWDyEGVO4w
hQiCF++FEkNEz7uNiB6q+S+7YJCYMF+itZl2VZaOyQnNaUUQq3wY8CpTr0MkPacq
fyQdDLJsTOSLFP+hLXs+X4dciCZ0Om0yqw6FfkcI8xK1JNEyWGFkJvSdtJx19v7/
+vAE+KO7hZ8Hjr1weJBBuOQ3SJqbGT/EbAIOThHkn32PbGvk8JyxaFidIWOuqghZ
19m9vnfyVEpKivyRIdSwipZudtxLQxw2seoB0HhSLkWJC+7iwTey2tb5Nbd3KJBb
R3PX2lPhmoDh86osxVka1M/91WUfEXtMe4A/JPVKLtDJThSyuHEj8ghhr5pd+i2X
bVnh0l4W8/kVNJszzuwjtUlJY0yP58vgOURy1h2yaqDFwWFPaVyfecrDSLJ9Ah39
W7AL4W2P20x6Z/OUGn+RDHlOH5P3gdxxHlALpQXgShj1b6sDqOM0VitVfz4sYDZA
5Kj7aDBvKLDYKq4ERb6V6UuyLlAAMMdAks2Ogq04TEojd95cdtKcNdiscHzXvjCV
PzcDfOacRr0C5mDviTpO2/NUdCzUD/Dtp3BaCvXpy1UxhxMF4wQFaq+SXW/iQgEy
3IBk/MsaNNA1fOra0rDfnwzZLxJD+2dRPlxMhjparDVqWHOq3aTdM61sQH44fOa3
8GYDBzvMshvYFxDWZVXP3rmitpsiX95jIJSfxSofHiiZe37sCx6V8ILSGflRo8dt
LaCw8bywn54fabvxkMoTRPoqCSd2r98Achjim4yEsFGK2WsfeEqLBH1wnl4VJTSv
W1mAnrI4XITuX3pMwonqF1MdtZtLet3ixSvZn6MHcUEyC5NL0nAebaNLtRAeAnXX
1yE8zYWYthqY/lar6VUxd0mnYNXSK36yWYjuGu0pM2EpqByw1ZwPRRjAg+7AlkE6
TmTjcc5eGS8MUexHyjJQxku/WL7F6mw6f7euKZRM6co85k5T8FdsT/s0ZC/Fphzn
RZAs96msg7w6kp5u2ooVZ+qSjsO//P4+9hESjitjcebps4ac5K9TRJQH2DEZ786S
jFN2M+v4p+Rg+5N2v6n9/HXuVuFDQEDV/qQXKsl4DSqcB85TKma2AN+D7GkGWpzz
Jxa5iDH8EVn+WsMGfFT2cDCl+/cA+vR6j9kam4QDjBRPAKzuhuKyhCSlKM5wqmMc
QsnO7KtKXGaKvhgZjRyZruOBCRjroMgQv6Xro+ST8v6bEmYpELAQoSDXFjaYXKKX
fb39elVW2j+ju51r/8Ba3qjDapIp8pWO0CQVUBMJl+/Gq20NCw6ZRuKKqQtdmo5+
CWIqib4vYIBWG5ND9c5azNHludLRAtGNtwCdiQfWAGwK3/Ft9Dp1MPevxdowjy2L
Mp5ufRHw+5mV/O+7p5NDkJxaNTYmix4ClgYUos5+jh5MfmuMFP9HQm52QuKdMyYx
Hl1nJXnf+5p2/xQNF10P7ibEX4Vs9FN+MSmD+dWNaTlR8waLaMQrnhugxP4zWYQu
S5gV4V+poo42L/w24sMn81qnSpNz9VQyPxum/GQuyUxjqd9slDmiaZGjEwBevT1G
XJSYWcz0qMox2fVACJ4GOIUZ/T5r8V/9GUIsT+cdBgB2glpue1y5/zNSJ6arpg3I
mwDDoaFzfcMX5KGKCm5ha7aXGuQDwpFCPAeANgUU+LX5PGkh55jrRIJISy7h4wc1
OFhy1E+zHfHP6WfgBuOv1I3YHS5NOrqKEJlyYFC9mRFXtGibHJTzs7XJjkCKTQIa
K4OHtsc9a9H2p7oazLiwlBT9AuHW9fs5kdw1AgruwlwlsXZeGku2typW2USz5BA4
TVPY6R7kSK/5WDjHeeBbc9/Ym4ATNwqE+YQdDA+hzs4nLFpo404V41O2jbjnwos7
6Fu+MkdhjkeotZhHEwh229JLHTgqTcDqPnerZjf+GF6yPcGbYO2txYGFoqRrKT4k
vqDuLR0oeagQQEopvtsoOfBqrG3WcDk9cGcLsY6JIQ94AvdPNn0nGNH9jwIu0/ac
Tb24NSiu5ZtsLrO4Xw9oK4YuwpuqEcgmwMIW1s7z7XBohkb3O2lWrciHQmM5Qs0w
9gPcY6VZUFmXJcv4AZ7ENdLEVMAqOt0kXppFgbTODZH+jyJs9nK3w37Cqfd0IHab
yT3rwq3/3M2SOMEsTFsCHBfUlcnV7GVOlfQmE7Rh9QmEp1XSFmRls7btUZI71mLw
vgIuL+NkQMM0Y3mIFhSr6r6ZDXI0nN1jm7e+B2QnLW44VUNsEdCMi0kLJhJhCxpe
1nue9oqV01+TALWQzEqPoie6OkTMHXueQMJufBfzYLG2s5v0Vu0qft8O+A42rbxb
f+jtaMetgvmq8f5Xv8/rBTTx9nud4/DRvu+cKeXqEUuCUqNZ6Gnu6nFfg85y+snz
ZsgSUTwoBQMQ5vaz4+g6HjRc5HW20STBiZKsubTXNs+2Y1/vFKY/RnFaUvVcrLRw
IxOGcqthQ9kfU0Q9YTuVSOu6vjmzbGBIURcwPhHwr2rZd2l6U5GkYp7TyBjsBmdF
1Le79bp+Zpx6z1qW6naE1c0pUIUG5Bc+NhFsxUbsGoKF7TMTGf6uvdrnWxEqqVmX
V5yhHp3+sM6tr8Vsr5sQku1OpfxsfsHsLYA4sreugcCeqCZbgPSTeFhbZqxXcSmN
odfK/7nLq4A6Y9Yw+1bxa+B66KSal7ZluqodfFSihHqva/sVljJdgSaGUfHyY0xU
8j/w6ZhDvFhOsxeOuTU6HRhU7sbNeUh2Vw4wg/LhXw8W4PnAfliaTGYyNkkp0sWi
PGzNtEwglo0xpeZfYmS01/FRR1hUWm98maJUbupO6m4LrhgrXs9WzVOMP+SQZPcM
MwAlnzE8JYYcDdy0i746rVONqS8ev6wyd30klLwOVr06MSLwVp/T+2jQR2z2yQnM
JUq3lOyrzNRfCV6BkUfYvpvKji+JMBxnivS00UrwMEbKhM2CPmoZQQ75UkKgXFuK
WuJ2x6Ocr/7dOEi8AwzRqsfkac99P8gG9XMwYCb6AOFkzbV94/rzDZSRKkr3M6nJ
37MOXbClROpukjljZrgZqGDuU0ZmLRzBNHLThHLlCqFH7AXIKf0Qo0AoGcnHhT2y
1n2bCwK299yYq3eL7O9P1JPLJHJHJJ1UoK7ncZUXe5+/WpSVr5e+8yBNWyTwsPq/
lva+UthvTP+n58EfqpOdJfHUKgdzuClcvvbuEEY2Oz3TsfkZJ3ESKgBN70KwALSh
OyFA0dyQzIVorMiPASQ0Pn9zqd+qjG+EXsSoCa2cxgLvdapblkprHMoX3lwy1Qu9
KMepxITWaB6OXNXKvR6PejyJVUgkfXDJQ1n6tXpIE/gptdvxVU4DYOIR4er7Kf3O
87J+xOaHPW5ug2qb9DaBcZ6zksJ15et9+1SC6LquWsD3WPZVY2YvB/4QwlHUWNaO
SYne9CZI17sdW8MFNx7s2sH9aXZw+iz4UoxMWDrL+ZDKNxznu4rfrNupeV8ePF3n
cRAACCCnYy5Z+kinz9QIyH823VoTU8AHCdOx9WpMAhu7t9YvOVhnYw3eHKVFTVMn
8/+X5fOXehgvyl13Vk7JfG05/KYUT2l60ea6Hx/H1JM5XjMBPWU9Bt3Oktw31OE7
Lr1SP9+PzAzF0mRBXKsv4RoUyK4sR62/c8ZEACns3at3oKVmVCQcnJ10kJkapWrn
o3Lii7xkoeVdPk8lWySxNlK7g/ZSAAplOZtQxP54Ii0VDGbRM8hLb+DnA3P4urJs
w5tw2CG25VXSpwdHd4Qh7cKIMpQXkKIujbV2OucpKVLzbrHUqPVZtD8R8bPNfL/+
u2dhtT6VVpWEep6u2+mhst9mKIHhHfOmoeJm0iXvnxd37TeBh8xhw9cJBk8kihK+
7XCpcTFUu3kSDM4N6zBmftxT+cRH0MVd7AT//RGhAC/mi6mv5m7lwtouqO1/1HnO
AC9/n3BswqYnGNagR09b/t3cUo8EmEojaVCnz7iSkCx1eXtGqsmcRJHBbXFbPnzJ
Z7yhx2FUPNHWJap0T16xkvyDQRGgDFTK0PSdtXzgjFU0uWFcGosYJlV/Y0kSiWZA
ArXsVekcOSdQ9WkZX4ghf591ruUQ+i5nrlNzGdlov7mQN2ovWldndTph19wXpFYY
Gp9WJetVyhw38tEEYoh/8N3q9Es+6D8IDLcruufV3BeIikV05SeaUFO8ZEK/k5JY
qMiDeTQkcl56NEO1lqaSDGVcurO4SIWPJRrfCnA8lkztTjFteRrJh6W7F7lRvYad
fiYTm9dwkLmXFBaKoMmoYZgvOkefr0nYirtRubdu+n07tqIX+RNNt+xuF9eG5epq
EdzJJYepj6cIz5yfKH6yRYdCzew9MWSOuy/KV5w4aM4TTwGSOquNpRPQ6MPfL5z6
YbExTwTOwkZdU8b4RoFpnfk7NETZFgOK3WuDBj7TIBbtPR2HnpHBQccZXlXjWLZo
emE3mqjVeJ7EpqSiChaqii28/gKWCCiJjdG6EOF5ueB9bfPj8ezk5NXvII8oN7+n
u3wI/9eiomzZmoZ9l+34iriBdUwnxZypBC0qPI73KXp+bynzC4g4ogsZD6kjhdmX
XC9dlu336nyvYG/nBWG6Bfv6BshYblqaO7K2zoPwH/wxIt7iKvrBhQI2AfHUYi7F
btcsLE1g2CyXaFgpopavD2TGRDg0HaINHh1a/o9qvBAH2uwDiNUJMsoSUlO3/y6R
GNS+VQLNeiVxop1rFaCtVpZ3hLEPMBT7d5haOmLVEu9FEUjMvKfxjMAcNOvwW/lT
vf7sdcgQ4H+YHzUFLxj/RXpbwzAywWIB5KV7Crtei5j+3/KnjFvvOGfYv96Z744o
B7j3S0VUOsCV+VpQeDx6DZswKJKKO48UPEnXp/ZfwcOOZZABBJuGoqnpTH2uXAAF
jTUlk62IUZtf2VaPt5O3nUfepqSKaEG2r9JCi+aO2nG7T4aj7d5M82LCw0QDzQc/
zCzvbj7zgWImV+SMh4VZmodIoUvonvidivHRTSqG/jlODL+Li22z+osZG1W/uY/L
b/LN3u7NfIPQQmg83wWdbuxxBzHkgwW8Zv9KVVd9LHmBkjEkTAWNWsz2EOh8R5Pu
3quAcpOt0CPtY46lQegsBSjpLzJroYGgXYEf6ZNaI7St6Cn7q8c/RX65vt7I8/Z3
YCuoFkGrylxGFacaOeCTay19yMnJAqErlmzSI41TFg+BOMt2r5LIETVf4F5upvCD
41uSeopS8AHgDVbqVyfBGldQUiyipyceGIaxQVJMjIjSfPKBqTLRnONfxOoifLXS
PIS/xXk6UmS3vKmgHdbvULyOjGBlZxQlI9S8Kbs0Im8IWaz0NZvD4BQpgODpbmot
N3lPVkk1DVMLnXlwD5z0HddZ1Npy+vBnO1oMSk4f1Omdm4AEfsoAke+9bZ0QVXLn
mJStasM08SAYI+R/ZMM7tNi/PQ3DR+z8Yz4d59Ryvy6rARvKvWYwxNde6dfnMOCT
rRiYq+rTkt8YskSEOuQmlo95cJ/0oDFnVRB7GMVlyvDPghiK62l+sGKzQebzBwXs
ugAu5AUgGV+7iRMezppPiSYYaBgWk6go8Zh6a3pHxwNRNeIl5JUqqB33jBaZ9Ria
vwkEa1MuUdeItKVWvZw3iBgr6WnFuyHzso+OuhPl+6T5iw/nAbhbuaqCiJeS9mX2
oDP5whY2UhBmbJNRS9537CnFpSWeqaAABP8xdGqhbSS2avWoh0YOwBSQwjU8er4j
CNMtbxpIuJc86E6QG94UFcZCiA6f41iZ6uryUcSbMd9ymGJwhPkF3IUo1emgqqf9
LxCKAWkuWNfKWbs2FqF4N78C5qIUQ2iq7pX96aYcVJtma1EnI12FsrKyd3CkxnrD
gaQmzynNC09yqFQhjV6xyZXvDEUtjKkGhBOMQdIV041/gfqt+RAJNgq4O5xuPyp4
MgGclfzjF0VjrePuS0lZw1dTK/u3x7JmlY5dFUDw82PsOW703oGj4E735p47QDNi
qkiNsA1mSe0/n4cYKa5I9CXRvf0ZsSfbiMvqaoKkvScJoT7jkrmCH8hBKWoCFKj/
ZEDomCIIeVlyoNvD+q8aZP7GsD6cz45LXHKWl3HEEHUsbDc2T7g6pDmKdk/VIt9g
FscMjVKCopocpxjJqNHBuXOTDF19z784BxD3cTXMX//FOjryutzbVEGg6OmDuS36
BCDkIVoOntW1RAMoJ7RA567Esl/r0M0hCFHj3RD+CyYptE4TPcwKRI6Zs4Gu9wgT
QdHj6ddj2WJrttCNUpJrZGHuHq91h2IZxdIPdr35SjCvrIoVmR0gahb5hTFhNv1Z
c5FvUGMhyRK1dMNbusmhlaMDdh5mGjGLPdT11ZWR+E5N2XN4w1T0rY8dh1XlATSw
h1Amjn9eB8fMjZMbReExCkoRlrvxvxrQd/Y7ZF37Eo479pVkWoSRzK5O93eRs360
7z404fkdYieZB9nci9ab/F/PKso6mUYEgSIqLRorrNwTU9B1GYFHLpRs6xs6A4Pb
ZXCVxu4gf0wBD31aBCj3cRI48iPJguhS6q4B65VlK/O1GNON/p/ndo8pIpaINxyO
5+O+YxHVU5yySfiV73RNWqJUuP3PgpmlyOpEEOoUB3VkOpJ3Ful9XR0PTCs0CiUN
k4R0RYVVJ8ALmU+jC9O4bqxU5J32DuikkxfhKqItsw03RSINJc4HiNCr/Cj/O90v
vDtjGlp7TCatpXQbUeXaF9Nb4kAmjZviTnMb0Xiry8A3i/k4KtabrfPeSUa7JFVj
QqqXfDySZ+Nj5mmm1/0JOhDqabTnEHF1B0FMX+7E8FreJUA+4bUb5nhR7Fzn8raA
YfbxAe6yJhs+Co0s1kYu2CXgOPW3pYm2Q728KFsemn4ruebX3cLX7y1f6MT/7lOR
7alDiSJZCz9CU1IIeCtGEyTGZvv7z24nIQmhybfNb3B5ej4aCg6KKHTANN5sAYih
XzpLJxR4SzpQAAN5uw3fMEFwGmoZYfAG1mpgfmT2lTCe67E7WoqJXvturXKvfwY9
7IzfAMAK7JFzLm5jP1jK9qcX+EYqfVmNxAtd6ZGmoORFizO6bomeUmm53OlSn8E7
ZM5jrULuuys7UNas9/NpCiHMwvmgRM5ojl47BPQOtuiDVP7R8JkX1wZbwNqNIiLW
8pdU8YRHJKkcBOwr2myqT8zpiz0Jz5A7UI+OuTVr0/ig1NjT1BJ+bOCa80HbQewg
3SPPDEGTFEKMsNfAOLq+dG7rJKN+TeFcaTh8jA6s1pMQZgBn+fRccNi095fIqWPw
pIedGXZFlPH7F2J6CI86lpJxMRcb+eUnkc8JULZ/sOJOLi2UL2uS6a3pxe1je4AN
QKSNhMxhIL5Ugrx6tnZAfMDacXrHDyXF2wAp8jNkWPN+IRyoy2c9jm7kWY+E0bDR
uXjTawjBcwjun+JFjnvyrlamnv8mkySNJjQQX5goPYFOA50EePERPcqMl3eBLmOs
0T8IDPz7G2/48ukxf5weX14KU3VTg8p1NLtELgL0jS5piapdQ7QxWbZdTwOPDsFC
3z56pvWwKpGQJPa2M8KNoK2vWAXxDAtCZwhy3/ovYF+/HsnvcUCJhlBK6ibrbPLO
vA/SGOZE0xiCTMrFtpJ1HMaT4l7pLSLvhNNPX62gSYYZMqaUy/AfY9n8zqRpT6TZ
4gwt+03aEZ/N1tI+i4zbmLYryZqdQAshq0J9NI6xpc53SCcGd7W/CkNoRy0ptSZe
NWuZgkCzkjbf7eOCI9CoRvpRBCUNaj48QnCj0ffhT6XH8o6DABDdc/MY12aAlhDX
2f0EnUeruQzCOFvP3Ounk5G4o5DYgEtYsddOw+m50OXXycCO0QkvTQCLl/KKE4b+
wAcQPUARSmMdzAcCd3uTAQGHW762PUYgTQc30ObY4uHX6OgGJuXK7S4Xgw3suHJc
0/3AvQHwamv66IW1q2mHjVwalDyGV8uvxGc9MtM9TFSSL2QXVoRbcb5xwd3ZfZVF
mGXZ/NM2fY/vzOkBumzvoJ3KC2OQ6VEx8fVViFKAjFtypQcsAkxn18yNyjK9Yva+
h7tcqSsJEjaO+S0lOidm/38/TRaGw3pt9vWqPi2pw04C13zyChnj6/VZtgfmkf8j
OKcUF52cJXjDrf96viG8cwELogrujmouEAtUiFztibC3PwpnwasaBOsM99aYJH7v
GxdIQbyoUB20mhPu0hnaCaEI36Q3lNyliB0B7xyXE/sFik3y5CgqP8JAf0zrD0h1
ppDlIz8y2yl0janJTNKMuByZ1RIFrLKkA88+vKB6AyiLbo1rAKVqwIkbTOQvNQUu
rNxQfo7KNR2loWTKKd8PgxEJK1fZtmKoMLct8JNAvXNqJcMPscjs3Mf3sRLKMa1B
XC7Af3zrHq5yRHd6h8TR/iY+5wULnn6sQmO8p3FHEYCaLWYBpV0isJZRgzmKiXkd
dZs+QuIg1E8jmUuFkOFuOinb2z0c1/p4ohH2EujpJ2Xq8FI4ffM1Tx8KmdYG0Vqb
+ZoiUedNWkgzYu7NH3NSacteFiJRSFBYuA16JOECS2qoymoo1UugwtOsLbiHcg7u
kTCxVGiaYUBrCuD1gCEZp8kp6NS71utDEWWISb04AtXD2UBY4EWH/MqhSKzrttiC
10pz42DBqvI8wqlFRXSdGsqhKkEpOygJQ0WzV4+45y6/wxCWZzrppaDIn2VvVVZl
2PHdjymjiQIMt+kyObkGBcEa880GX9IXLz4ZyXNNEyoNYYfGb8esCv2BJef63iV/
M9szyioa2PaDu1Pei5fzVnLIpjBxMWtKj7ZulMp8kiH8rG3y0BRVy1FXwPNG2QvL
02JeUHtjAHGuXicij5VLhtYzxYQ0SoC9nBUKDMOB5qZwqbzzBK4uxVKPyxGR+wAH
P/f0SZvFCx++fjFWWO+i7aS1u5P4f2oWsbowXYfrfjKxQfXdx7DzyTTpIfs+L5uK
V0eYR8MA1nFl4Hb15kNaruUS3cPdOAeZpzyAuo4F3wxzfnuLfejnYLSRNid0ugkB
TwX0FmuKG5rGnbwH/Cd/AvFm6AGF0mnLaGMWFE8sAbiEPxCyeCRS9MvFMxi+GjL0
VEisU3yQEwvqP/7jSIQduPsRU/QFUtMuOwcBfZU+X4e+MqDKHMgIhEWbqmEA0Whs
WWQM1MjUkcgziAgqokEHMFN29DAaoW+EmbWpIo+ZpWDpNVZ8UbVsuzC7aZ84ovGW
olcz6Ygd173Jn0be3PHH3oej8kl7ey1S0lTcb0f4Pgpa3H1YvspSgKDDU82DVC/X
8vJ6ryVBpBRFGkU5jiIYId20VYJ5ak785ML2HaoZxWMvd1sY0TQKAYj0n+gdoRlP
qBYWdb8plPv3NDYtTBBM/zSD0bgjQzAMkvRYBprekBZRFN42WNxiRs6eKjz7gWo3
HAKBWUuumSPWHb4a8WbIzpUyc0D29vRholDVNKC/Alk0dbQLS/URdRAPSeKS7Zc3
FDH+2ylCrTMLxkcPSGmdSLWxtmQMy7vTSNJmxscomHZ3K+pb2Ea4A4exjbOmQf/M
dBFjadE3HBok5eL38/HIbYKFckkIRxIaGVOEttSBCEEf5NI5UxTHE7hXOkaDPf3K
g7avEd+znTerpH6PyDDcFOYrU90AKtaEAelG+RfpEomK6m6n3nnCc+ipbL3nRcpN
anpRETcMTOCRHAW4LR5JfRayhdq2N9c8W3o4yodQwvxdE4LplDv8NSEair+Ph/mX
4MetpNrn514t6mz8CFfJ2yh/63jdnhJLCye/B8isxAOOhuwi/tnOh2+wGmCfboJ/
k1CqvTGPiBrTbgqV2ZfMKpwZ7QiRqP3nrXvVV1ItEKW3ngWejDhW4pCnoZqIMMHa
BCXwgpsntOHC+RD2aHPEbZpkyuU2BAEM7d193hDDaOYVAQEDnNqawxqWi3DYDFDE
f5Ya9Cvd9k1MIoekNKlNhLxLSZiUtEAtjcJYc69eqEYnVtN4PIn05Kh+vTcMz90y
XymAjtWn9QTRCTcRkfvHMv59AsO9uYOSxJ89/KyEVaHTR2W/7EogPkDFa7lH3WaB
KtBXvUAQVtwSPifrbQ4L1MNM7dc2dbFqSZxc/XJEQlsqpw8urbgD0QM9OGRT1uWH
kd4PIsxkRzWDa26OuCqRJWDNvcWsS8nM0Ol0azxCK0Zz2z81UvZ6M/XGiAgOapps
styZRcD+NGXgrDe3bJt2SPm2dzA7Ovx9D3YnyKbeXkKHLLiiA0Vt0F6Bjk2HgQWC
K+0caEivDYLZh16ThM/EdV+oy+HagOLgEUCMCZkq3VudZwFQjfui8fg1w8pT3S2e
U4Ar+lG3IxvIgOcwiar1oZ+dJzyoXRHIk0Qtrjs4FDzQzhBTt/AKV4pMq+IIE+z/
zKAhhGi3bvKhKymRhnwEJ3phtxd5nQ99LNqEzsFeQ7GiqQq2P9qTiXhC/f0NbPY4
t19i2YjmiO4Io+SqJJLRL+LCZ8NP8kE9HPoCe/5x7YjJNPcG0zpu5Xii9QipNiQu
5DOU5mn4/0WsWCr82elHj2ShciOfTmdCKmFBuqwabFcnfzMO7Z50zDEiZPIdqycx
5G0AQG89kfMDK0kuV5XCPM6GqwSta+tnsCCVepEMNdtAIMxhsyhEVksvCON/cNVt
i5fd4Dppn26jOfkrkaQL5yFY3yGEISRJX+aCJCB3kBJKmgsoohvZRDUEUYjYvw+v
fHJE7CKMAchjHur2JpU16+HX0GM9Sd+Y/pPIeGPfoxBF9Di1SpAqUAjfn3Pkb39L
oQ4R+G8nr7UdvRj04SeTxrBaa9QWXK1OwmiG6gcp9nQEQnKX6GpiZn4Yo1Oct0tT
d2mv3CrEAlLeAb5akGBHuFX/og4Rfd/u6zMnRHAWDsrYhiqkMHZvYg7iZCUQSUwN
PJZadxwgJ5ZdiUIvPr5Hwejmv55XG+o6KaswAjNmbwoKHjvWnZsGPrlGyZ3yawlC
rP4s2plqGZNdW1iWs9uev/UgvPUbsiWbKh6if+pCxOseHbKXC6L49JAoV9QbNNuS
Mdm1jPW9lgROuOHHHLJqcR/lSvLClfOfW+k3XipuC5LgMczZQuQvwATU/pKN2abw
Xqe2HYeGBj6PZikY3pObxYrLv7vCjfKowYrrTo4x5LVdhrFgrXF3VOK1z1gnqGPv
oO1Cy9mZVMvGfqXEiC0mCxAfn9eZiDvIDAY31DHmAYQMJIbqxVjEC4EfKwZd7TWT
XcI0B5FYguVNK45lbmzlkhLsQp7UX275XipPJ4Zhi7dCAVo5z080dcCsrTOMsyXJ
BNZ56vXdDt8lCbZOFxYymvs0IJn5OMidTyRWYIExai2pgpzNcTUGRYjRHnVnxa0G
eTMmugfhygEcAMC3TR7YBjhC6At9Biyerk7kGOCwRvFzY2hRHldoDx3hcnJo4uAo
2umnH6VwWb4H5UQnZA+K46K1imuVWX2cy2+3l/rU16QN3EK6wkfghuJ72OsdcVbL
EFvndu6hAykCYIMiq64lIpfAge3A/TUaSqX9BGt1HHaJHZQogDbaIJLJ6hNlXASE
A+BKnn3UkNroBc/Gzr7ooYv/yQQ0x5b41yrjqr4WHahLfAT5FZpvp2DR9VvP2ixu
lQX2oriWck8LDtN8wx58PDnaZOxw1U2LMZTM0OYQ4xsSvu9tw+H4NPfQkKOCrokP
kWa6RMNNub4vhEkkzKsnjXECQfLNALg4+VcKpAkKHiJfRRz1rFUmi/0JjP+MOVOH
FVUF6X1pJ2WfZQWlyDKnHVPnmirhBBbrgKRN2LsiTR3LqOL+69C8FS2NrULVORkg
icECrrdm3y2iupISd2oJeBdklS+0e1WKAZv60aRf+acYgNlW98O5DVbakqkKBcP6
pMBTV87azna+HpcBDusG6TTa2CDthEXXkGVwe2cqUV7Eojbwesp6bRIvd57eVKzg
5h/RoSL5Ui3ZtfiN0LkznHr5lDg3O9W5ZXocZDZXl2tFKKarjpynDQISMwtYfL5L
3tEjC/x35vfdqnQUKOly7dir5YYlffFRRrCV2rYG4uB7+eK3SJmIcZyVTnMNpmjc
cfCRpUSKIGRJPs86dqsRhvSAAOaNujzxQRSxBdab0eHLJVSJVNXlMSNSSaYWsOZ4
VMZyi1GUVftNJsStyt5V4xSINbyxevcPVdRd+kJv19K7KBWip9vs9OXISyTXkHlY
Ijgchwd9oaqn1L8/aodWSNzQoSfCse8S61+i4Qt6BBvNsLpbH5wv8zG85m2W/D5i
lVDyEUmoHAm+DaomOqX85maVtUvAnWBE91BYJsD6gNKoXvuS8YYjh50Atg2QOoUB
IFxM86gjCyMMmN2vKpAO8qKGKXqynoVrjwvBBNRKAw5wAtDQ6hWNZ7lhkuNXaF4+
iZu1BtgBx10T6ELVteR5ETAAk0nqV/i7cbm9LU9dF1xnnwDR/dSa+Mix//KvlEnN
gNC4BrMyGkEfcCeAgtR1Zwy1vfdHt6rxAmEXrPz7BSckM/N5j0EUdgaDFFDnMnOT
oelZIWuBS/gvGWvOwDDi+nOPEu1pdkDZlO9d/r6WYrwfew2N0Ah/zC9kAbUaGlwI
+mUmDFy99OjVt9+gujjpmwVuL9KRoZ6m3FiAuDe3OeEvuCnBMAXfUDx6m58sdrNd
xxOAV+rzfHa98CbEYgkcm6pkoLTLak6AEUXA1vk0L7MWTTLI9ij6SA4/Ei5ioukK
7R+M5vWp21faMe+/4533Wm8jrT/4/Vm6LzfMzt8RRlWw4kZTl8cv0X/Pm+DzLdP9
nALWwpxqEqW+pFEAaGD/6gAGfxPWc6u78ZRX5hJA/vZqs3CYbphekTfKU63T+ZAc
okgC4mq74Bpz+RMtbyGv0VfUGpjxw+UGOanux/lEzLnI+EnCrQYYf1j7fTaPywPq
RlYuBhx47ZEiTLcU+l0K6pZxVuF6ICJbY9Ib1SajYg3lVwOyalPA3VBmdecssrwT
NdQGwf6ICti9bPT2BpC//gpkqJk7HLqJkUyInH7wcJXzLL8JLgPpe9a+QclwYj4Y
kg405QPweAcjs3U7AFhxe+2DcE3JQSX3WX4g9u7kne/U72T6y86IIaxDI33gNNlg
HBj+E4yI7CAFJrnk/abrph5K8j+GQaD57O+m2zvHbB9vIfybGAtmsM5ZpmzGZHZY
4rAIAob/4kkZEcyZUfz6V9WmJ+qQeyzUOlWuwVTQ3VlNQW3ewsDpraFqZBOSWzz6
C6FKucFZGfv0b9afSxIKSSdExDUN4LUr/A0+A8Y96SQ97Ake6N4PafSuASSAvNuk
ueEas1IGOzP7BftJ/4ZaayV5x94Ao2vBvzd5Zswkf9UESBOjcSNsWOT4/TnazXFa
0LoFR3iiHJg7Tx6kowd9RnSLIrhCBjqckuyPNo2gbomG5roSSIuYicrvcf+qM/Iz
ZKhuqObLBoHix0gHTySSh7w303YK7vIZmJHEA6sdsOY5vxM+yIItsO4o5ohB6M36
yzwm+KDf2wU8Md61gagAri5b3ZRtWMb2WjripdqERXkCTTAYesgJigfL9O7/tjn+
F938ZxP43S8cuiqadLFR0DuRKhTREg6wKFUxMGbTVNUEsPef/vyA7TxhLtnn0bDW
quu8ZAO278fPDtrrIOBMwpP87G+ffN5RYrP7waREK8d7vHVPVB2CoaJATyOfpct5
2o8x9APHlEkh+YFUBEVV3d500MF3lu6kjIPRBha7lr5Rg9jRLPGJCQELENztBakv
HXb9Uao+Fybismfg+IekI8SuTpGccIt6hJ4Hp/S1awerWAcxAXnMniVb5RKr/3Jc
SudtqA0cDRKt3jnpfmAk1CGcEhBNaSnb9x+lEyK8bRxStj9twBv00LYU8IsqSxgC
kK5aJ6tbm1DidWNiSgQyae91lC0p9u2h0kA/vxI+U7WGK0ymwl53v1Me6WEPfTHN
U23iMrYmQibyg1q8CU8fpipgO9iFFa2iM8l7PkmvyyrADtMTP75aG1uz2rTGAR9k
OcHnWEXnfOssFRkydKtqg0hMfn50G3J9ZgdOEGjdKjQ97s2kxjegqNSe9eED4O4z
p0mlBkGDNA7XWIuazjqv97hVMd1RXwWpGJC9mxLYYNfHxVjQvWRe7EvdXNN/sK6G
BLgTj3kWPOfN8/EM2R6CJ5/HYrbOoJKZMRVTTF+gqqM7t49tqc/xZIXlKY3WJvRN
j3AxRBjTfMrEj+yHBN6uivQ12aVQyngjthaqmhXZP2C6IUPSnt+8Q2ecPu4G1gBa
l+gzz5fNZlhskEAVbi4HUHFr1uTEYkGrVst4Pn30veq+5Ln7ndpYPynFHG1lW+on
nZO6UrKHMI8/AIlB5nG7HdHHdDCqsMWrSWTTqvUA15rwXj0MXlVHLuAfuhDI4eql
RH5AwBMtpY88juoHw6TEYfo2+rWZAT6T5xoqupHG8Hikvlskta8eaVQ0Xa9OgvSe
QHpsaWWjlTpzmDClwjDUX9KIL40X6eSv2On6ewPHQxGlmcQCblLA9JDLj7kzyMkZ
GgRFs7FPA773JKY7FlaLtTuhfLpngqcAlk5on2n4E/UW/uFaPFrNfnHZFsYnVglv
cdEwBhIrjsFaXsLrtw0b9xmmx/NFRuzEn/z/Gqiv4Q6lfz/C4hFAYgqEfFx+uCgl
+H4ipJf53Q1+JBFhatORsKIl/yCzOvM4xRH+U1OxfwMfguk756QyS2EmxrtwK5DH
ABW/whgqTJIBvLnCnlLfrNa/SbFQHp/EHcWXy0aUjFv9twlKVhpKVMfrRemIhIKU
ZEVrtsTwrDZzyt8FUYM3RruZzSn/2+aSspS2XO6Z+8qtN1DplBgdGQVN6h2TrX3z
8gME3xQGb93JbAC0Dlc+7EEZygurQbRPMA1FaKAgEO9eqyDinNgt2MfI9zkeYmmK
zgNqHV3jE8aZq1XLEHft9N9BoJSn0RZg7Cb2CazPAZ/Bn5PTBneUTRFVuBdsCWb6
fSPJWFqqZw7wKfaEWB7l4Uhxge9PKrEpZaZnpMQkwsk1NM3mxFz+zlEUwHQOjHFJ
RWipvu6GD1E5L95gCeiCpQoduNh4s46cvxcq1XZmyHcsLcnq6G5xxMAhSTb7bEOf
ClsBTZ97ph6eyeR5+vSVpiIbcMriPcRvNxfvaFM8W7M/cbB1dEJBMGWoiyr6dDRS
QwHyBQhlwmE6XVlV/TsySwOpPlwvHfVu4WKWZ9YC/VzeOxC13jEOuX+xLiol9qOH
dX4KoYduVgV6t5iiC6NbjVaQp8KATts8tUU0m3Xgo1qI4+FDG/aVszUQt7lM1UNk
24m6mnmYxHGbhgTADlYf6/f+QMg0CFzIpfnzWRo95h5n9jgWLVm0SRer/pf+H6gn
5TLB0uHV9nOKM+NfCoGD86Kuf22I7WlL5JaHHzWgXfr8I5CRnKpVDBWqZOUUwRJk
kwewIbf614dEFSEBg8eKW+l9NjTw7L/9/UJeW+JkzhJZC9SXNBh5RpTBHSjquh4P
MmyFFkCOwPA3vbwipflNdKDvN327kNulIlzg2jKvFLhlFFucHDy/t9R1dJ+i4jKC
G7xarAA0YEOgWsyB64jSkEPGItgd3kDNIC0qpyKe8vlgo9T57zL9ex+5ybimc9me
kFGE9g2d5/q24JhgyFGx3WSfQMG8r1cP2mv2qz9hGVOsX0GPQc7VmUa3xZgJwk0a
hg4UxV/X7+Yqa+9QWTubSm527VMyXN/328IZbIO0kygG7ujXOPE6EpPQ2Ux8gAJe
hzaZt40ZOH4dCODBOAdMUrUrGJ6npo+LWhIqm+0bBeXDZg7V/P9YX6MYsrrJenhS
I+5XJf3stuVbHh3PEGwOCBoxEPT3TO5jYQq/YP//EV4lf+UpLvkrocTPmZ8Jodz+
iVrJSFY0x/Vt45eFFZFwV5DPqV9I2zhTtSku5B/cvvN+oXje2ciPQOppo/5uWv+i
Gk+AAFTiHXuHfjzceQwL82ai8asS4fQitIUl5cYqcMqvGxPRVOjfBHNaQW/NE+Ev
loEwt+H5uCCpEQWoYAy6hqc2wILdMw1xj/9avD9l3luJuwqdrUo2wIKsZZj7BOqs
weJ3MoSNspTwMCq9Mc7xeWrtQlVic4g2kmckAfcD0oaPND4GjOdIYKP9EUAUjP00
r8qJaqPMQx7xqmBU3gl8sSbDjxbVJyt+4bhcamGRanw3ST7AJSANbbxBCBSvO8Uu
xczDDUPNbnn0w7WeRPkdCatoDJcDbdeJjcTtE8XKC7MJZCbPMIrXxnc53N8RlQxt
52e739lp8WtQb2VrDmoAr8OEwHOZRealiSVv9s3Nr+Fynv71JEfby26F7u45tXjK
nMNEoxF7palQL16J9KeURdH49KQnaYe6wdd9cOWRW5H/Yoia6Z69Yt79u9halU11
USHjrBoUxuaoXelGD5HwDDT1ub30cLV69eGvOy6wTeGKpeUXWUv3RQkN2YCICJ17
ha1RKFQcJQ/mhK7c6ruCgCGYuV8QO7LXKuFwGjpz8y0VKHuFjHtAWZ5fVmdwvtuC
boaBhHBGZM6FACIFUNyJCh6eOU7Ozq+gDjjCTmYUee477XhPOZVUVyDW4kVnZYU9
vYBgdMZMMoG1WcZ6mLKvPKJ+WKCk+1dQYrzPElOS53QcCOblvcO9opOKUf3b8I/B
qimDS95wcBk8C8ldDrYrZjnjjnpvsCV4YkPMj3YjktnVY9Ad/gFFyepK2mB3M8S7
lL4UNG65VI1gfiwSbi+uCNfBU8cvugpfGA6BGEP2t7Rxyn4q5qIy3y/IlogkWyjq
n7Kwirik2ZDepIP4h0fhRkKm+H4yVwQyYv6+hDeI3BEAAQBC0/VWQLNhY78nV1fP
SpdopAX9kFn0up0oXMb/vHP1FxHJ+JAC0B+ZjbHzWRU34khCmL15hXDlbHRv7jOP
YPnVYw9lk1iAjPQ1RKFO5Y7pcEbGgJp/OGANjpDmcQX+1Tm6bky3QIgTtvvKeBT7
CrBwHEStbalUWFpifAfie6kItpo37DmgRamTvPUiBMdSfsbs0/Xr1E/sOhWjg4S8
RaOx28L3DhepBB5rJGVd/py3nyRH6Dp0IQIZ5kmDLJDIlTFdPCehanlMoYD6cq/a
u9v2CONmN3Q11bk2LrqgpQRWym+xar4VgzXppP9oDW3uJMScBv0qgjHOlhqKvJxJ
NqvYvIQlZ5ZYV/7lnXzC6zWuYKoN4o0ncm/xM5JUXbg3ZqYTnCCenOdPb5mQ7tyU
h16ZgxBLS+cgKPv/ELXgSH6zCKyW/YaBiNtzg3vwGC3Fhi07PkV2feQexDG8CMxp
LXe1tM4HbD5sCXF0as4qb+3iV1JuPA/kHBfS1DHdokHl68dwerY+GLrluhYy6saL
NZEBUVQMe/SYiMZHMPX2BbEBkOS1gxtA0XpJQPCaZnweUMxHy/wCda/EuhEYsuu0
rDjZgqpEwDcYFdpEEOVhvZSHhc0Si/adddx307J7QpALOH6E05qz3i1/PTo4Lcxv
ELFIhNB+iuiEIgXMFll3v2pykTJqjvfuLN9tBiOxVRVAus0ksZk22QZSTGe6/1hy
5Tm7paMk3Yxc/VxCfs4/1N1FQ/zEbG71jsDa+WTz9RQrayBpYnbkTHOM0E3WY+Vi
8VU/6yC3MQaA/jsUhFtDY0efX8mpwQdnkrOjQ/wxqyLHZMT7Vm0XPc+5qxumITND
yvT8q+QD2dZhIILtR8cGyYcN/N7rLp2xuxcHAk3NhlE1Izva4ZcwSfmADTyCltCo
1Ey0OHyINmM7AxLTdWdYWc7sqFI6cwe6RPSwuV+Y4Q/dQn4Mx7GSaD0wgdPxTEqu
dwASnDlnqhV2XlTe0ChqLvFmFdY4Sh1403S4y0gHUd6f3z5UQMfqjNq6UfQYEqE7
Wt6/vE0IexaNBDXfPShiGJCLF3/W32P3+lVqFR2oVVd4brj/4Crq4/Wj2ll3g9wU
fTrDQxZLfV60q1L9KMj4dmWgAcUiDgihsLBYIoviAPc1Eyp3rbCOgCUScrNdTG00
O3XjnmyGpwlD6FrNW+5sr9QD0iFv6e+qEenwtDc6AfXV+ZJQgz3AIfG9ApsVQy2q
AcsoKB7EYGfRlZUlaYMRq244qgmlkHsizp6nB2fwdKbUt+drX2NQvO3VJfG2yI5k
arpbdKFgL3YtlTFnmT0P3lYg5YmHKqZF6jUT9WksB9rPFUhZWJicpiOeFIaj3WLN
9vE7wDSY+KqfyZg4ZAtU7+7rgFD//kUIZnEKJICWlmmz0fXM8pQyiTIGErPMDvPd
Fk17UiL597TJAEVPFC3fG1chG4PElRycIpikuGeYNzHvKNSTeTRu2Ve0PadgZU/+
pKBgKa+rB2fJHz988CuSqMvDPoQ0nT9DZjSBPM0DkS77Yj+O21USYYY7DBT481k/
WjbkYx/AmRKKRy9V56kzSBMSmkMLHHYFqqg4YWkJSM5HPSfm1jhM17C83qxnm79K
RjVoMDe6NfTGKP7Y6rOpENkgdEKCBmVHkLu9ff7DqyoeThhUq6dlGQBKl0AMKMiZ
ocuBy39leBVAo737QoDVfAbJhTLPh79/qISoPwgKiEgIj7kK5rwBfsg6BziofSWX
XfccDEG4h+TlCrLSuLOscxqnyr2+X9UBm1MUQn4xXgqB0URpWzWMcrpWSwYqZOkI
8lQm60p4sXdhqWPCVNLnFkGN6xkqWJ6kRhtisjz4aW8HhXSv8UeVho061Rx//eXl
1ZWAT0mTsxvroWJa25ezkgdGL8h/NQYs8H4cLaJRa7VIljfwxyf1R62nPmzY+Q2b
4CJ7PYjDX/WjjJmDmFZqMzHn/l1O0B1FCctY1xnw1RpPUwqVP0W87EKgWDMc9tII
oeVyqUUAw5MEYjGlexc6zxnxS5OIQRGqY7LfHdDhMCHOljXGuSdEo6fbwrKR/6n+
mAdarP2mKHbyKVXd8SvY6Vi24Vxi/aPNRAiXbNnOpzljTGbJsaZe669QpZ1wKMSi
Euu73jPII2w3Y8Qz+FRiDloP+5pb40hbCUVwizUuou3huCKzGhIG57i5Xil2OgQS
YcnKArCjuBWF8yI0gFzKKF7Q28IZ2cutp9Gr5KWRcIKkcNMaeaP1z/Zk99GGWIY7
mOEqbTpkYLNIoH6+FsVaRatEy51le41jCUDp3mtUeJ4gu2WtLsvW0gZmQgzn2pEQ
kDQdBloJq8y0JxUgn0cacyVR2hKh5sB6aqSYPjesVlVeFJfx5GvtjPR9RmZdR0eB
RmbIFnTVTbplcylkHVUUI6PvBsmHQ9Ijnwq6km5TAoQMnz0+4CBhiU6lQ45xLLT7
ki6IhNsjW4j/nNByeixNa/xG3LzfSAkilUpTYQtN61JMQ1kXQXsacxcRzwDxiJhG
ho+Lgf6okeEHGi9OZPt0TeKdTd2SYfjwTg3cbSHRxKf6xtcRcQUvxzyMsiw9icjn
G1SW3qcq/FajseYVPmWE4ZHHgYOV3182qrWqRVUt1CT1q+LOcAFhy0RCmEmO1vYw
+Dzplrey6+jwYnewXl1Z3/caVOADW6sc2cXn3hEKtamWr66s1pNRJnux5rH9jBTN
LVbw8qBcoUkiabG/4hMnEmgSgad9TC/DceBW+jRjgX9BJF+FTLCKdK0kdrnurjCb
T7N4P6/j8kgoQeG21kobTSfBtAfkWaQD3UpiEtMqYZXNo8hKncw/kKSy3pAduTmV
nRYICG5izP1WRsTCXiJOYxsbeOOCmesXeH5X11B7l9AYGyf0WqsEHul+JfBGkVfv
VadLSt18g4eDXodYeC9pbaD7OEoB5//a63nmZSW9fGPCRc70dAkZ8u0PP3f4q3+S
QaSc/Ed0LMP6t1YVWG320HWO+SY07056VeWf/s4TTdfinl9/4ZzI8zOgUN2MdhAg
QdXWiWwkW9I+M5NDSXyZDQWV6R/F9x84RnYdFcImYPs4/D1/EzSqr0WIUrWvvrq/
WCJAa3ew7QTP1EQ24oIbqJOIAGXFPkaz2vNf90LJR068NhJapbwUelqqkDAoGniQ
deuvjfA/KSXE0x3uGOTXs1FuVecUNHQroLFM4R28aWFIPBQpDW1mr12KhpNOvI/w
GcCyPxeMU1oEaitMaP4h+qlv9PEmfznoKaRJo3KD1hABfsyKEF58FhEF7a8qvWJx
MrAUoSC8Qn8gA/r+PbzYu8tgK/s+byD4vWXAOd5BWm1vdRTsuGgqHUXiPPK5Fy8P
YR8dkTv2wgZk+2FjlzQB/NHj/kvYBBkBfelUltIc3LTg1miXJdgai7Na6vxZzKAj
GmLY3Cv0tOQ1iTSdvKb1W+n9MgedpQGtt7tro0WMU1n0QoHdo/0QjatgqjcTVSm3
G6qLpGocakAiX4P62HQGOpGZUmG6pfIR/gZS8VaPqHc4YYb6G29zage5q5dsovXM
PCfACa1ADPJuglg9eVeGG+FfYlPUuD7o3h9wvPNJUBbAcKHnn+iOdCFmCEo2Kn7j
DG+zkS4iI8Ul7uAJ4CepJuTIGCMfOqddut+y9UwS7JDer1oaEgSVlhfPKyAGV/lH
qVV16EJ8euYlzL3rnFJLnxNk2WZcMR85jQLkJOF40ZnGdbFM21zpC2lUB/Brsad3
h7zxmVb/uxKUXZtPRTLd8IMdZXcrTbXO2zawgFrGS4t6C5zHYkAVeTIMPJK37FDL
k9S1kSZPJT4xItBrXmPtHIh6+44cOAk04bM4cPdfxOqXnXGQgf+DSHT6cNqZwWvu
L2mnD6ZIRtBKYfZkxNZEEh43gtC3+CzrZXnLMAu3pWRx6MhedbXfNn2nL5ykyBRo
a+AHr9xs5AGS64wIW9HtV6BB8/rhXB2dnwXtvJDunInkQH6+ZFos0YivPS4UgEPM
LXDkg5Kjbh2JWJFXooUn5jVo6PC12Y4/2y8Fd0rO0AtSjCUEyPz6f4qAakRGHkek
VD0gSHEZHYoz7GdcHa7Pao1XGDP9WoCqb3D8h+VM5NfOsJ/C0EbiEt5ynkFr2Vm+
TvW+B7CDArmwXzqEFjMIKmM7+hrzv8ecQol3fPch+q5Az+NRp029qC6yqXGTgBGa
59miUIptSrnD/PCB++fMkB+Qlnev+kr8sZryTlLUDFh4tQJ9E3M1eS0AaGtWVzMv
sfzCMUMXUFmEjX3FdA9WUhlco1SuGfJe0I43AI/5iiiAIxGHQLANnBFndQutCOzL
67WpbWu4biPBWamujMZu8vFdGA6/g4XCmV3+xWwjCacnC0OO6rfPK9k67g3jakPS
3aS1CLTNZ6RVoYr2ZZz8WGevvcGXZbBEjICmwY/0fn2loUDLen83l0rKfhNyCQh6
tRYWJlserE3qaTqaCugLuoQ1H0RVEbtJLV3crB64fY6nj9qDbH4qUvERlDMqWNBO
lS6tsC2V/AaG57pBQ6Xxr1pQgf2pvxXs8mEecHnyOYMJKO6SZyNKpvG2aZcCA41u
LIHAzUOE/9s4+hD/Tv8JbZgE/FLQfRnywMKXbfxnkNp2mwz91iyoU7SoldRKQgX4
EG8HXaOaIw2oYVMbPRO4z3P4OOM9agQpfJOchO66jrSfIyU0frr2NfmUx1g8rYGt
eIUpmq1x+ws546K3k2VGYnkXiBjFWljQ/fUdnMWG1Tqkdqd6kR8hbm70gTOIPYa+
3Aaptj7uI1uErajWYVMk5+weYmv6mqHvsa1PmV3ojb3fDDjPiM5Qb8sqmfHd/PiZ
Jm+umcvruoc7n95c69rchL7KG+UPGtsottPAOywY/VbzAYi8ZBAIXgazZRC9+poE
PGDt6k3qnrfQoi7+GDM9id/cUZqQLjorurycTsqO1R1E7q2w37cuSAQAd0fhbdn+
y0W2uo5OTg2oEio6dqvJeHaScQ3wciyiRijFB8nk/cQ3Y0/TSbvref8Ip8TYfq8F
J7xkHQGDdbsaoYLFtXH/ouYkR/fO31QtZxvaHscE03cPyTJw4VeEOW81U/z/Vvmn
2xCF46ctgR9Qc+JeJFyNgQ1M+fJbNXvHwAUknO19Ttkt+WjnVoBpwhlS8qEDjfV8
5FHqROIASvn80fn5HHEDROwojlB/q4d1SRlGyU243jyRzGEZ/os90LI6HPgz1OoF
chNfjV1u2VHa0Mm8gzZqmRSjgLrzVg9ZYiAWjhX6D3dl53B5r5k7kRdRaVT0eVIf
R7IUNDXVc/90fHdUOjApjBUtvz42E0fjTIZ6rSEbltkobee3oPyRZkAXkE9HYqTw
ziKLHYPqrHVnBuMV63bA6zvQrR2eTD9aduQGneeby+MGZxHBMHRswcDnQBBlQmLW
LyizBNgsQo6tuMBH7WhJfnmI1tx1b+SV8SzaQ87smbDxs6X1ABz5tIPCPD09ShRH
5mFX1yAT554+XnhotjnGskso9t27wr2xBNGKcSH56K6cZFpXHlh1c5EAJMvoZvSk
0iSQIz32DS5ngkEaSFihjl14DWk4ggOu8oHZb9l+6l4TSYBI8/ydE3INCYodDfh6
c6qdMMoOYCvICcCcbfkjhCci7HvrtBSBy2IBGblZwZe0v7D184swfGq6kaVNrF7L
ik786BLiwwKXKfcJgziPkc9krrfM0eboRFkV4o0mz5kAB16EfXSNN/xu1i3DttPu
gymQJLRYtS9zyx0lIHAHNUQrr+yvzaGLtwZtM8tgLiTuZMCwYfu02GoAD/Wblp+D
NMFsupapZdjl2RhtVC0r/Hc2GWWi9t57o15abo+xeRK3cig3HHEI73orYER5TPjq
9roLZ068v0lY9NC6swFtABP44Mz1IVcDPE1XbSGgJFAz3eRgY3FzfFitsiHY8ML9
GAl3gCaURiaGUccjTMZsuyX4uUPuldYNCs8oUHluR1CEiaCYri+S8p1wMD1WDWRh
JixmbKJQHM4FVN0aK7VfKop094YQnlPwjeW2VsotxJVd/Jzrh4aoBv4vDp8vsjJb
0QUXeYn+VAIV0yJ3/sHS4ff+NsSrWakAtJPM47RrmPWyMrnZajHQQSe+Z6QQ1HND
xLjK68mwCH9zliuC36CEtCBNHA5KvXWEtnMjB8q72Tfz2ttwpF3BQVsQCaXoC2Ym
79IGc9LuJg004/TLZD0qxSb3dupIkp2dezxCvolEr4KDAdsFyl8f8+ZULAm8zL6S
LHMZBoM+nOVBnM3PQnGVEoY7Ofrbm/3XcT5KS3DPSX0fgG85ajghytyEqJwaCf+b
BD8TelLLa8+A7rX7LV7Fh0nGpwfMcoGNzqkeOCbh2M+6y+4V+K0xD7Fhxtzq2mDJ
cvX36aZQIgEOYeKCbRqQzUcIkkL80VihRRfWFLWsxwoLaJ1DPKUZoSLwzegnyMWN
UbzozdTaQKz2x59zALV6AQ6ooxgvDo1gyYkIE7u4ImQ477moJgpBfoTAQIhokWjK
oLg8LkUUWVP1PvBsMGI25c7RFZp848iB9UvviEEUC7f9dUcqeMFp5DTACn8lmTfI
cOwcY+q48hJg/DCwt+Vurnnvo32kV9gby71ItbjzreLsvXI7uCSmLqCprrzhDA+u
h7HC/1lzbuS74oYrOQWrJu20K+2igbZJUk46VNHGlEKEb9WyKXUlMsrEk0CySEWA
uxc8mu6HUw/jbQ6f5LdPkisDtHAklOUJkWyKNTFEG3C4nPRN/Tb6Nghu/EucvXu1
jp/JHRGc7JRZvufSiQ8qneaQ0n+11FyTYuMrIUj2xtrSjUvvr9ok6T5gL8KUNLOz
q/AcK5Y9zrAMK74Jkux9cTAtrAkw0mC6o/LHq3qD9UmoT80503ECsbhZCNGp66or
LKxcshQaSGBoe9vp3dCv9ewp9hLPx15jB4d3Af7p+oy7/y6cmqEHrkPDJrLfBO1o
5Bk156jR875uuacAM1pil05/3eVjJ9dIz+iob7fyWxpy9xRAJiYq25Ezx0/YDHx1
dI3lXH5EOm3TU9cb6zPkoSuEs6yZEfGneWbUhV4/8TK4Asl3rawk1gLo8r3o4O/q
fPAkcYBCvY+OmDAjSOkaCX/MinzrGY8zftHanmuLEUMATb6lDUmMCK8pZFFlwsLf
6MIghVTg/B1+NO5gsFPS/pN9Blzwe7EIFFxFjgxmhTwT3wiPeYBrN1uOHmh0mWe5
AqxqB5FOiPWRfgdkd8vt3lHThlgj0In9KEkSzwewvQ2/lO9gr8sCjDrFnmVI8UvR
i+SDeq2NPFGyTojpu20oq64y+ftIcS/t1SADg3zBVtP4qvGXSgPIUo5jmYZBWu/m
MLlbL2QMAj0vUPVfWlDzcA6PBWjjJMTXet2bwSyqhwyp3aG0J+rNGiR9JFkOWB3B
SSUewlvPZaa8aEdexyuOOlZjLG80dhvYIsKxvRFnsZxBf1XFB0ySfqA62s7UkEmT
0mD+PzYgQpIbDTmXKRrT0DiA+sw6mBruVhZSM5K4BrWorzZjxqca5MiaX/E5t+hM
SBi67XAj4VBXQTNsQWkvBrItSuaUrHTtj9hSWWBgvC/CTSIsVHwQv0zHX49mOFMV
5r3RYzkiV4U5iQ4YY6XWSiiR/gNmVo/j0ApOdnTyLvgTUonHxMb2/YVO5/4m15l4
tgkdB/5K+xpEZ5P7KH5dpY3Ug0hNgBsyZG/qlsbCiBlnDDU0exkCbmVjYtrYZro6
biGqf0TfP0MM7QPrUbmBlv3TxueA5eI3NPDk7H4LADZ9CDhw37ktAA8bRIqSoDLj
GFABJEaZxMGytcRZ1+lK+c511wQ1BJH8zmNWJFm+6oxDsf9zA7OAaLMSKU1wnLFW
RUpUy3ZWmXRIO2EuJKFx01s6oNH3rZSABp2d0I+7AtGhSIKcybnRRU/vkXXgzHXs
9rCiA95u0zO53d531VWUiDmDxeK5rY/B3obXyPEC5HbS07aBe83O9asMgUjNtf5k
+brYq9Fn30Ua0zP0rKDR0hZubWkyWgKi5uB2xGl8toRv8eZyys3DEghDyiqiU/oG
1MxveJwkJzjf+hjdy2ZVftMjHAiugIFi7P7oMhVWq4vCk2HWICUNKAon6USXsGvP
dxwJCiQikA2OpyWGT1HLCZ5iqAVhz89PAsxZov8MoFsYrI5Qr1dSw0fsEbfGUan7
uMtI2jkde1xbBNHrqmdWuUIm6MDMMtzrVLVO1dLe4S3bXXikxq2EvFTAJrvuDTWd
IDhJm1pKXH+fyGyvF+ECcmQbG8N0kTmgTXc5IJKRVcMoeU3yup+Tcvvk6l83fCp3
+bHrPx5enrDQQ5lQ444uJClInvYKrwbIxzThOk9HNLTX5W68AIBpWq6YQ4/PTY/k
V69cXLpjqoc/5CqtclULlIjQoX6OlzNMGho0TZsbeX4HX8FgkNf5mbYXZP3uoyiE
TIpoa8yIf/OB6oR2wDmXcCj3R0DOgE69A5NCBWB0NS4r6KMdDavGOTv/xl/dXDM1
/trEoYCw+PhaA8X+ytcBwhcUeXgdGj914YR8xxqri/TibsQnI7qnwLI5pBzVH6MB
pwyStkvxsPz2tIOYI98k5uWb8ZC11F6KyQohkzbHQRR+cnw6cM67s3v32HNvq6+P
HJ9waLw/Z9uvP3oOQLOXPNG08/uTmNSPWG5kIg7Krf5kNYCBB+dWwqWYPW3rx3D7
/K65taYMzBAkDEYocGNm3BULK1qOKYFidxqtai9fg7D45Z5HeyAf4jac5vYKbgf5
pvZ5aq/cpuJiWA1KtJroYCWj7v2yJelhbZ9IwSMxSX0bE8madyMWTjWjNGP1FIt9
Xx05JtU0/2EyRFaycEXNutd7N6yhX6eqPPtaz4Jkqf59Ev9Zo+PXyZErAm0SWjiK
3cJXAMlIqdHBViZvV1OwkGzrbRetBU3QVdAptWEMDG12UXz7riQLZ3Sr/qt1jl+F
MKm6ZhhhH31t7W2Jbg1Zi79X1ZmBzTLeZ+ox1jhbArxZa40WF2srIOBb1z+RkxOi
pTPzMaJDIk84ZvTjr85pgIPkB5lePw3MSrOGa8w1p8LkSQoUQUHsSpM602U2wyaV
ey10qYUY5ZDfPzOSpGsQEvnMD+QvKeHeFgJ0stHycdCIBjq4NipeA60KAgu8/zHi
Y4VznDfsAVBpqRnHLfg6GPJ8zwL1X1es5q/UQm5SC8KoaFHDiovH99nRmjoCWtC5
DtOlDUHavLKXM+9seF6BbPpqofx1yIKXL1MntvN61MDxVCs9AMhEneUjWPnJJppO
1+UJtELDfEv3gRf3t3lHq1XXZm9RKPtXMXjdD23dPHVmsV0qrMLb5vXhGm+4/3kE
RN1s2SmuryqTXgf4M91zJZDtaK8xHPMYt86dF5/KcfjxYFySMRocMjK9vDm+2qEc
zMSFGK8Jlax7Xt1Kda3kAURI+LilgKZ1/jvj5TgqcdTzNQ8mCM+flwL7+/I0r1hI
ZgOOYeOPtM+O8r7sBZJaFWOhjVYM+v0YMMeoTStwhXsA1Llk8jfi1/c3ps3v+QhB
fZ6hhLbvwDLNZSfH4mYvUonTN2sUgMkxr2uH5kyQWu82zoGb3vY20OGaY8SfuUJ2
v1D5fzh+T5Z4dYcnMGTSwXbU7fj+GplEIUpG3P4ehbDUW+Eg3PQ/R/U9HRBeGYQt
s+hPculMPeMBhQAm+9UqIAuZmYUAOa3J7h91OimfD/9vNrUg6bxdGaHT4uuG2yV4
VlCsdJyf1DB8rGQyP0xG4zVZwr6tXFRMJVH35NmT9NDpO9TXCeavRDPE50siviNH
lB58Qy3zri9YpbHA8+iSlHnbbXX6txeFFJ7B8Grp5dE9dgT+5kE5NpX4SxWiFTou
U8i4W4+DPDx5sme4W5Ergx/xpyRnnxVcBoGx0dLAk1Qz8iNkIFpUSW4RijdmXgIs
2SR5nE1DesP/40/5lc6kklfAsOp0AfLesUyreBeKuPZe3GLAbMldtz5pN4DnOy7p
U+ooUyEyry1VnzvkSS28Nbu91yMK2BnBKCvKJHfUSK51uHPAbNReqyKtsuDqJXrW
lLGBtjkjmQ7CnH4la41Il/OFSBRR9jsxMqHWquwArrcW/DoQynZvsQQQJZGAHwIU
868GeQ+wjdKZz9f5dveRtsodF6CV13XCDRuhXyZXK7f8H+a4u5buN4w2tPiK9dtK
m+X7+bhw51JdUVGOqE7tORQ7nNj8ffgx1Q9rpYnC0G0/IDdBpQ+Q2ubv2hiGz5fD
x7N9nWIUR2Uu5HwE3LHAL/DovCsdXsn8+DGhu5d3Oaq11vDDBTk5Q+mxgMb0gUcr
J0zxQ0DoIgWoYqM3VHEEyS9xmrCNWO3DYU+JYXd3NMcb8A7EeYKxSl6jUje+AF3F
1qmHO5qD+GqvimHN/BhX8lrzTvuY/FX2Gg8bPwadal6yMaP1TrKNX3WyzptQoajC
Hhwr/by+poHfqh5DQAZCHD9Oq4TdNYeHFqbCj1uFkjWd1o+VJDY0jRpqOP3ziFB/
p6UCGEmx077Zo6uSOjoqkspfZLcsLowP5JlmmwNhev5XqjRbIaI6MrQq6/rWpHme
dSXbhMYDAsSb6BDMTcUygwzVDjJwiTeRGLziwLsZeazVShhlTiiGsNROInMPHs2K
1AAiRPJUl3whbRjJVKA9fUK5nLqIPRlhRqwB5ygjWjvAuL7+UFGYLFr605BdE//f
3X6YinHVKhlmggDIyLdhYYfDbHu+M9zEHqQkGPLnooBFT0wqzjMUHCrPt0d7To1R
KWQcvloDmwbnM6lEoXTdVagZZ3/PqF5/F7IMN8k8UQ5q1wckn1Cp2wNoKR5M/p1Y
9TE24MG/bikmyycb+v760gEP9ErX9zg62NLWr0HLFsC5HT+Fe+1ePdEWRccoH8G6
+J4CZ7HuDQOxVQ9kPpBF0Nnr+jxsPz5CPoXmDbCIC1iXLUkmYPLN3blV2thaiR4/
cRfZCPURJzQiVFQIBSfbS49wfGwZ5/8+Vsf9FJ63Uc/jujs1VMLnojXkTz+a0a0b
85On9FTNSKkPcaGVH3dN4r9O4nx7FopOT3EN0EXqJUIIuz/SEO5ZPsJgxVRd5r9H
YvzJ9VXb+MWumH8l+EtMsPYY1ud7VtoREElyqOVmK4HG0x6CE/cQrwB5/UFsqA97
f0irABL2k705JVVVx40LirIgLLyOYw4RoawYfCOWGbrkFGFWXcNTaTRU4sBQUHH2
F5W1oO3upPIfIqzvtrqgScMCxUG1JJ+vye7bc1FaUGZO8Mcjrju9VaWOKRS+kjJO
cC0c/XF+uL7Q8MtGbwyqr5frtTJjKXoqymK/kobuTouFCsJGpzATWG5DhHbNzMGP
anqzwdI1USvG7KdERn9NAdbV7w8Ve1jyeLOPR2UnGIgq6hYz4q218t2ElDWPS8Ml
7xDoDiX4E0kTCMF9s43RdHnRrjHWpb4lohh7rst5tYsYCJ8T7WyviIbyJPQ1VBjD
dpXmR0jNx6Ln+T/1LdV5SYx1uFwxKu7A3N8Bkoiydco7L1uOBPZy3HrC9pd6PdPj
+Lr7TD80GOrZtXcWr+9J81IE1dzUNebOPlm7Q4QivkcUITZZ7L+02koikNliHYjt
kioslkllXT3hlIk1sx12H7qGqziWVdyytuO0Yy2yD1jwd+m+R8XOfzGXMDZR/pPZ
TKhpBbr/CVsJMRt34146g64tGD2YQJzxvnWMFzLhEJ/TJcsdQayPT0lEMbjlAM19
KRMfyneiK/G2WvEooj6lhdDcBkWbbtM5VDQYHGIqe3W1bguyvNK7MREi5Glc1baP
4uKiKYZISYW2yd9PXgqCaLaXtJ60bhKE6V8GaUWej6yvhf6vbJnHBDs/fhgqFfcU
uOLAz1G86VzuvDqPXuIC1fchHUuwXaRMZwNNzzhuS3rY0u3VlEqlipY5Pw/38ZYx
9Ci5hkVkls7BKSgJtk6puuT1B/UFVQOSC9Ltb992q8/S1vZbiPfA09r8IDAz1kGL
crOkn6u29p6ehJsVckKG1+Nvs+BO+FUrBVsEaAr1oQbZp8zifPHiv4hDPHHbsUXD
gxiegwFYMdm4zMxXFBt3oXg4KDBTq9g9KuDLvqSAtJxW8KcudjgWzQ1PU3hKuyc9
GlejpizSGUOMzZTYltzLzic9a3w5NF88ngTAKOSutrVIi55Iq21DuEH4eKlxFYf2
D8E5mll+44oWMEkiKv/h+kEz+ZMeGz84mRJy+GuPS3FZb0zZnU60aqkrg2lZWlx0
oXTO9t8bdmYmlGYlgGmJXRmFJOgMBqjGWYwGzCi9KY2SD1RrYr7FR7CvIrx6TOd0
//lwaTuF8tLEu8kg8yAJbnQMb4akau5AoTDzXNgCZ3W4d3Ylzx7WYKWzq/ndhhty
WqGjgHOvGeBMuHLL1F3TmP0Hyxbi0rMU53d4Z7+b/yhpVrU5TNzEAugY5bF6ghFz
rWWSLKnULsUpTc15xfLz+ga/zZiY580Z5bMIPdHAgoC1KsfiR9DGUqbBMx8yZOQ+
dPlW1r4Sc5PSGUUR32nM+GPae3mpwbNYDc53ut1d7I7zNUHhP4HxkUsjNhd+D7Ko
6rhArfQ7QBVJjCY+czrAd5olPCTZj9rvDE2JmqQKxkNjKQROUiifNQ7F/oUOm4yo
kPUw7UranoXF0rRktbWxaOsPkXUxFUsk5rWZh+X3aUvl9w8SInId6MVtaVHZRii4
1RdW2VwiLsvTqmMIOBScqdaQqiFyLIP/rexIn2Pkelsq21GLAEr67LwSED46XbEr
lTS+olWQuIFAtGnPuFBG+3fpOkDk67nG06CRTz+O7Fk6tE0KkgitqjIDU9qISEBC
bfDXr4wUnlNOQxERdCq3/CLONdLNH3NZCWr+Tq547sspz3W6iNmHh1RqTQmBBeqG
u/LKIW3YoADWNpIu20lop6pDvw+lqdnoNfmIha2eDCUSINtqXkaxV4qOPED2+F0a
Q+0NfHVeUnce2knW7wk9YfmnWWebAqHmEwZsyWlUE04OE4BLL7c2OeGCkgq+RP+D
LvsYqD5Hx4ORHEtFej4cKSRRoqTfmx8+8IT5aehSvYMkYGTV83e27STBDs86PERX
bXM2lJBW7ynM65MEQYx8VkcuFpcN9zOqF8jZZqPY+n305G+f0DLXIFEEGg0EXAiI
1OjCkvekp6wMXmS4z05Bivtj9jGsj1pk4gam9xDD6vCXrqDnnX39+n7OdRS81pTy
KdQ396y2ZUDdA6UhOP7mXzj2m9AZGjC2eR+ITOmqubCFeM/0ZSGlQpiJdop4l940
8OQ7sN5RCESA4V9EJX3ft4ivNTwf0VD6teh3U8L1uVgcaWrYn9HnLa8ThCV7/LND
HttQt6uBmkrIe64BI/I3X3TS06Qrqb4odP7pxVN8EIayBzzCr0ue85uqNj4kX/9Y
y9m92jOrqpVB9gP0wxSWKm6sJlHcDkRQIyIRgcvPRLZSU04iUezL6N2BMW3iVITB
xyyTk4S50a50Cwxl9iPET7KcrecCelp816huumZEI6frVTzXWjwYbNmxkm3209kX
t6taO7/K007qb9x1n3BGxT3WqAQrbDQ7cWCc+UTtxKA2W/bQM4kGitPidsmh6Y8b
2EbtMlaKzMNC6lrw9raCHE1NM7/6oOIpiXqIRa1SqwkD4n0l4WNHGJCr6IW/W48L
v7jB5gw6uENzljUPOzgwcH4psuH3sa3JBXYCXM/RFku//wKriWgcLxiTyLgp4gtJ
azPxPiDCzvwhgLNptKVwLnkFfbVx5D7kFmh8XPt0DuMPfdfsji59HD0/0rV62IuP
zUm5feszSNcDeaO/2jpj9b9ufzhFUHrNW/zqjh/5+LsYx7MhXYuvZ0+BMOOF4Tbd
8JpYxRvSpjjLnfJ9pBPR2uy5zU4iXTn1XUXo4sqniL4/4fA+gNi+lknyrBIOeKx7
QxVjg4uK3W1VATwsG/raA69vMw5lWrhbKu8FLXfkwIthwlC9oWtZNKozL92CcewB
BGnWBOPez60PhU/5uBUctjBEl0XEsMeySnQJUEfkO/4OFBijsILo9hWLENP3Fz9b
FmJk7oQC7gfw4EYmj10yxIPfap9yzruqSvPyt2sFh1jJFOeudBC/pJ82YNiEEWKr
viXLBuqrHJE9wM3aOdknZg/TqvdfQh9mslL3XCyBuSyQnGO/UvKkpHjx2qAvznyp
icQo6pS12i69kGPAKwGJu6PhZa5wvETYpqIvabnBAiM1nIREQj+vlD0OxW/nWsIV
lheweoMnrCXKwSj3VDHB+BtJOg5ZMoQbwduqBtjt7mgh0/AUZupRJmMg0f1chBAH
MiwMRIf73PmxJw5bOzOaCTPucsJwVphJu0v/kTilOl+6LlgAQu6YbmPyaOxSNBMf
RQxremP9/b7aUt5dW610TPYr1kt0K4Vdm/849iYJM/FzArPxdheQmBfBdXHSs4my
z3+lI4NSGbNYHtDcDVHoQR4WLXG48NuYlaTUm9/cwCj+Q+XNwBZ8ngAD7mz7E7/l
3WEaFs29IOZhJMY6dooX6Dz2jm4H8cbroejTpl3sWOvc1dXMwbDprUZ5HnETO17G
MiMnuL3TDMfwrCkSOb+tiaIhuENLm62UKERxhNuEzPXtyDZ8Bf6lXe2ApS13sk2S
xb4wG+Q0WNF0xyA9iBRtK8oO00f3vmHWFte4SAO98YNqIPL+QzKSf+mzXVcagUOB
h1SamgFTIPW4Lx7REG/YIKxx4TpeA6nj0/vi7HINZdy7fSTKaRx4USJGYrNhVxgY
BGcJIYe2rZlTFIk7st6kOzatLsBSv339BlG/qDFAAtArjpQWmpmsu421yozgyJcj
PcPHUiSwhWP29EXo8ZkReElVh74wR1fTaoQzNBzKNDBOhCk1CvqRMF1rfDYGh7ML
0d5YmWLK2ahsygm9mex0KpcEoY1yr/3d4aaJXgEPHBUjEVe+2gARzf3Z5S/qRn+w
M64bCxsJCAZQ3xjTMIxO8pbXt+2MeU3km7tF2w2f1gXPj4Vx+2KOTDTJXPSpOZyy
OevdZAIULEeFXMXSAPJpKwupcRj8P4fzroluD7YphumrfSde7FiV7PrHip0/WP6q
ZAksk0XY82UdQZ/7MzDVrx6nmJr8DxUjOcVW4nkWp5u42oNGrw5qYZ13JX9uTDur
YohCj1oRTiewZYPpeek6XzWcyt40cKGLP182qLD2cvLiNo5RUcthFaHHO4d8Uitu
C8UmIjudHnDXz3nv88W6tImC/N1HnSQEEZAhhjWeJwXzrmJRtCeB5Lg0ZV7t5CCJ
228c4xYpubb7IugvTu1e8o+1G3T6aaEpJaZY+gxsqd3WxzDmd57h3feOV+WhdZP2
XudFTXEhCkrPfWtu+qN+VvKf7iETcgYLRPoYL8aXyf53dAe5PqkuGdOGwTnYyuJK
m0rAMboXTrkqYqckyV1AMolaVXsLDJlpApoVUHO9x5fKmUfUdGWzk6HS4B1MrrdH
lh4R2hgX6nTjsabBIgaveuzwOQT+49bI+gUCEQeF6SOfYWMy+oLhLOFm4++Xlyc6
mPWIGmHaAxtLhlxM3YG58FPvjkXbn8BYb/EwddnuwAG1hrlmGnYO36Y5qXvSQQbi
imlg7CF0um2KQy/2efCFVsnXEH9MNm7soInqlQZGMS+4wdbiBs3mIKAf258wgCuX
bI/+FvF4Y2HaWdaku+fUNjNOXSvNo+AFEjpBajTI/V/dlyaT33FFZlANdfnHWXgm
IIxFUbQ2TlP3PfCOw9UggiIiiAXYPSLVTtj4WXO2KG+OUVdIaa75nWTGEd1J/YZ3
1Cn7oWbTGkX4UydE3hA2dUwh+7OD9IZUAvHciiDnNauOmxub9wpcgdOshoGEBtJ6
H0Z90HFJDXomG1agBoo3i95Y5xV9lHDtg1skl/xkyAB6VuomSf7dbUAYD2UbmSHK
HQfapXXg4rAHZdFiU/jGivTEAL39vAVRoUwXC8g/fKQWey5VrPdlcyo1+N59+Olg
aAH8C3nOYekfzLJ+pB7X30b5LcWa9JNKTXyXkZZ/Jd1LtxFIaXxb3+FqeAnSQyT1
FdYwuhJpICDypT2ZU115NZC6+XBwxk38aEgBXvDp/cxF7p3rVic6vlAo2AiQGO5W
7QmkZq8ehI/QcHNgRfN7P1D+jHEZ0c6pVT1MTVQecTYJhI5C0RxvVfaKYsuwGZtP
U+HGESzGAAOXsvael0XMiOSSlXAC3RJz4/LD3KnPCJioIw4WETpZ76HP6RdacQqb
42etzGxCLHpD/e/JQsEr/kkD+hg9ywaUfo1PJCwm2o3S8VlRt1VY6rUC2hUvebQ6
UZDRcRoH6hec97uJ/fvSJ1uWCSKXCpZnbW3Jkxt12PHGRh6jYSUfLbjJJj3CiOVY
uhBLsKib4JjPy3iobchfb/h7yayZFJS8dMQvPzHrG21MX+ju+uA10fr0AB0SQ2bX
gWEHb7ZVmm7FLoCsunkK+V9jPrcrQ0RC3TtPxoLPOam0UllNNnkDyc9MNUZqHQxp
2H9Spy1Ax2Ad8kX6Sta3LC3QCbU81VNS0BmOboDU1n2vcQaBnCQzCgPYNWOZIe89
BvQegSUzbHlxepLHEouo22ZL/tVrs3ifVbQrfrMMZeuCn+gQiNbHci1V0xrhN3io
7qVSPZSknuSMdDMNTH8g66zX0P6pIOeXsCiqoNFbVMrCumEcgwdvlHyk2PTRwfvM
yZ/d64QpIALyX31QEsat6sn3zGiTHYmjrbpZ+ULB+t2D15r0WFxLSZUOOnYret8I
AHPesb4cJHlFpMzu06IENiqj6noBOsdCHb/2t+QMQ0TdxO+ojzFVPoikCdcw8cto
YjEY4F7cOSNrIWUonIA97J51PU6hmAY9pfVxmdpyzE3l9TCbLTxdFvTK2eJS6Ktj
MwuLPGRRsIzgIBBGlfWC98e167mJI/2E9IaNr87V0I348c6uHZOR9DaCl02fHLoT
iGbFrzegNH6/yC3v2enAWxGja8TQh/FodY6q21RSu6PzqoXfC538tHOOE4S5c0YH
P4vqHzYIuz+nvDjaA0Rn/NMXgZOYGR9PTQKTc1CGktcKbiJARAqD993Wgh5a5Vfl
nn7GDKMkYhiJ3wU1k2iGV//zpuI/QkWQDMDN7QuwNKjngrmlcrd9hEk0M1AHJRO5
HRCKL0rSDhZPJSK1WfTvPpJEyCJx4ECDiNaYsZV0k1wfYDEavaVyknjliCWxlX8D
6pxLavEaX1Cxytfq8zsEM0zX8hDhcKENjv4GM0myAJFgmsTYIp8aDpw4t2cdR+J2
l2dFbQDJS8sPTmBVaVqNiYPZjzRpFiYjY374CJW341JKzPRtg9c8QxY6XIV0ua6o
br1s66J+6u30oXn8tNcm9G3WSKDATqxzO2eUmStNd0gyYXhpu9ZQHdpAPvFno3Zg
kUUBi6dkwv/i2eTPXZSUQR9HlO3/0cprbIdG8BjS8kF1huvGA3BkpQ+GmW6UO1E0
b0kSTAHD+fh0J927mLnSpznsF6Puu/TM0alvNPrCgg9i2jWeE/8faT6Ue9wWF9Aq
OnamYKBEGv+e/jeYcsDe+bQOi+fzBK2Q/7N3nmi7H1pw0j2/9mz9aLVXScDIU6ol
Ku2MNMEBp3w3sL4W3OCIpClRhe8mZMZ+b1A2co6eq3swFz/YesCyQ/kteLtSDPf+
zqbG6KZgPPIaHyVTG2QmDKkCS5NXEBzU95mMfedFGHRIw+g0Pxw5nM+uFadD0gT1
g5tJP7S3wWJc+rOhwhuvmVIWIndiNpWAdpY7nCGLanWH7im3e87rkyfGCfRrTL3h
eV0/YZzPgsqQdT6QY0uaujGkKoWFYgN/D5lzWPe66q6yjd+IAWH0IVv+hmq/Pma9
Bu8Y7ZV9Qe1LQ8k1Ha8X3I0a0HTBOLf9Bzzkf4QN9fOtbuLJ1sOcNrHN9axYnJ78
xdkdNZJL0eYB7069erlX5qEx/Sse2eKiZ88qndtWa/ASvUPyyGrgvjBRtgcqKmcK
sR4Q1uO7UL5Oi20zIFQagsSTBEdYRgBqV2lzNdqN3slXECW4EefN8jYQJqiaRLR0
P67DlKhjBsOURhpHqa9mDlyOHcO+CO1PZp9P3c5ZZlpgxELW6RIHua01KfxbGXeZ
qKfuTnqQAZxjl5Xz19+jE0cX+s8blzCBm4AxoKxjYAoIo+nI1kdFdtyhNFC4lPTd
BDhoJ9rJKaeCIwjW8O2KgfaohiVuVHU8Gbk1FBSCjePpT8yzqmKTu+UIinOW7n+/
XIOh9l80bVG8i3m6MEZnx+Xp3gKbM7/fki7bBKyxPXoDpmAOOpu+VhdykR/+bZRB
GDgLLydLvxb8seA/55eIqX8O1KMbGZ1+YyI4RNVTFHfiyE/p/h4Xc/l32f3k7lWG
R9fbhAHiKFrgpGgxdxWT8uvZoPGa2ZMuxAyqy9A7hd1R06csLiPKhN4C++8hJAZY
nOyrcw7QLvQErYyfPUnqirSJNIY9fGal6oJJbAD7okW8SgsASIaWuh+k8xhXhGMn
B2yEXClRNWgYeFwnDsvcdjADtiMxTNqFbLRlzeab37CgRNiwjrTOFyyKLZwjqIZg
SGHCTtd1nS69TjCbCRgv+uo9K+3L0jDLweZqt9mkcbuiMPJiDLAzuLMHJIY81186
jbGHDg/JcdcgtSDLbDDKqZVgR/I3RR4wrEySyrJjfcGENqBiDUk0ScxEZ3lO53T9
gZqcfi+ELT9Bu5hvDBfkO6z4vHmX4rlmxEPwE+lL+Kte7nEF7YP2XdmzaYiBVbnz
MOTIpum0jDi1ZpW83x08wiAt/YAZtD3Z4C9AWQceqaIkUT+U7TqZNM/sMWKZVSpz
ii/S7dWRJrFpcgxCP0DPxCMfTJ+VSHOf6g28dtzXKsOnfyno7EZDZdwI0C+zJ5PS
9xmDKRTscXREEKeLzErXIJsiAuhf5xIVofZhJi6Rwwutwk0pZw6XKTLua8HGptSq
rMXojvpYjYV+P6BtdEKw5NmUGfZc5h96g8EiAUfkg07i/BR5KMvK42ML4bO8wU2Y
LDuOouTKAeKhIRLT+vFqtgWVHqFDus8KnsKL5ojRTTnUaYxhdVHkHMr1auZ7EkA7
9EXoBiT0knME1vGGu+waFdMXKXdUhnKkud6Si6NA9tNP4RfwDYFOWFEAmB1WWCiN
haApuNYYwGfFiJFVtM5u4GGJA11Pm3gftEOSroI8Vy2usAfgPMQQTyfmiFPcka9V
amDw3anw022DqXajde5qul1xbQhQ7gxU9srsEZkcchP8NudlqYEiB0JqNvEU5a+T
r3Xzpl694Ez10XWBieoBzkroewsvYdfiK5nAszVfA3Q+8+mfXCCv7diJPMw1yVzU
KdX1Bzf4l/QFxiYP64iN6CZDBLg1BEUkfR4V+joEu/gwTApKFvj738A/DCsZ3jJ8
eGr2Yrju8jaa9TFtYx1PAVbmciVNm8u3L6kYuhiengGEO2i+HP5Y1iV959txltOR
mI3JaWXTNOjLRPCSd5gKvzlks3UfKoJrGL2ZJIcFCuk3TCfhb7Iq/ff9wQnPF0PX
u2iDjGtan6At8Ui0opcmhSavcwL0BOFd8HQprBh7bZcSCFasu9koZXULWlgragtg
nAK4yIOBLBAudrqfgqtQyoSxMCMbLPdKL5TtWgtOH9IuIG6yBWOOqI9k/8mi/pWK
UY3x3gekSZPLz7Rykerf/QS1Edk+OeInN2DqUWL+D1ZUixLO1d0UXDm/ZOgyUz6U
ZrA41hRNr/AuoZUNpiJGZBF4CySNuSoIXLXEbUyy5lobUYd5uRstnYw22HC7fzyb
E9djMMqdhjZBh34gozEEAkNWrdfzHAeTRllpFBzDL5crI4fS3KcTltcwese0Ebeg
+60fDTk/tGCpI7VkF9KD0yMwwNuNmlHZory3A4hgQkBQKsGwao64+om9syQtQMTX
Ec96dwy/ul/DbNvY9Q168chO1sA8owL8Pf13d0GI6EJUtfnXTl3uKhMEo7uTYKub
m6KuvDHafFzzb653dRloRBMiek/jiH49ZuHBSg0CCjECHz1I2eVSRZ6enEUcRToD
1m9+PbQSMQ+4FKw1Pp4T2hb56KnStxiB95QNUQYA5QBGvRTQL4J+6WKzG/JVTPnx
KDReM1zZqWdDEdrYGwovZ+jhnviGrhVg0YCZCA78cXRN4LBDZ0r2o3+vi2x4eMuU
MMS+UBfDgWr6eOgD52AbbmwnEzf4WiAovX/LSWPwcwbE56qcwJCRVmZtBoulGq9k
BwK/9olu8t2rxyeMKG2jeGNbgKWHYpmCtsCl2Fwsk31dReQAUilCagTMeK/DFqJy
hjTl+NUZBITK2YxGMoKc9v1eLTuL+ALFAPMVVZbm+LJu2csHTzbn431YmYwkaIF3
458huHae125UJZVmhDOoDd7wtadowgBQu2vlxOSVMFm7lk40F7UA6I7rJqFEGcQs
FYRLpA4vmpTX0jQDEDy8/+crO91ztuV/GO0Lq09LbOvu+GuqLZiaD1XDrziUfPUu
jgkj4q3Lq2E9Fa/3AfY82gngsMdALzN4FKc4SmZ/yY4Ullx3yTl4q+FnauktvKzO
8iZlkbjTVKrtxDhW0+9iV74OduZ93E7bYH1PRuX9EvsboAjf619DjUM4LElDQeuo
HWcmCCQaWj3xdu+LQe/0uB4cmRFYBMk1FjRXuhHvfoBmPBbhmfulrXbS8W3tnx2j
ds4B7IAcypcyykIT9wMHyFNiSIU+pFsfP89JJP7OqlaMiE8P4CKaS0N7wjw2gtCW
uUPWW9oPBeeOhVcCBU0D4nqG7zqqJhsOJlouVwNYk/0YoUgQNPawzvP57Af6GfdN
c0JiHqKTCU+MCcQUDKLkHRo2bNWm3m687IvnFaRoMwBdyalQI3FYlxuTijxfgV60
Vq3fkuvsReJZV1C/JQOI+UgLIteRqZ2vatF2dZcU6wE1Ng06M7aKD3Bnnq8DQjpT
G+UprZ+Bh5M13OP60FEhGzLXcvGnYsElMJVsU8rfMPjYuChImeDOCE4u71gM3QNH
ZT10MpRs7Sc/xws5ZAvd9DkB5jgrrlpnDlIeTDd5lrSNftdPyFSBiJlmPxTRxqB/
CGYAlAS+8ENjCH/EtSdsyhVu0WTnC7LEdNDEEivPdWJItriLFH/FfEDrqMxij8Q7
odMN7OWVi6JPWqId/JrwnI1cSU0GoX8NhitTIQN3viBmS/UnnStcJct7vHlIz/oD
I39pGudxjVXE8XMWLfpECY1DPBTk4fvGNYSEbTIkIzr6GF6MBo2SESrRmexg1qOf
uydiwAPCshY9WajiQWmp/5Y0TCQmLFq2ZYASzsvYokmS8m/h7KHmeAGDC02twn7D
RLTHKbtN+SnNJrDQJWcknmrPmtulwQ3nlLEifA0zhqd6aaZ9ADEqQLqZ6x7L29ns
F3NN4nYFVBYJFIKRnVznaRncqFLDUSltnTiOZ2qqRH5e+7cMvl7iZSn1H6gFrEvD
Q/Sr+cNUSc3PuLZddb3578a+4Umla48+J94FVo1vhzlLNIYQYHz7BIYWl+bL2N1n
EHkew1SaafBbHREZvWHVTJvRvWaMROPL83chSVO5t5XWtUJX2guPqUv05aEIsklC
1w4N2jrwdOlrh6m0ITSymHG33/LuvgRvEo60ff/uhvmeugX17KrZQD8RyI3MkqiC
MIe5pRWiec6Qf51qZJ7SzPcCQ3UhLds0WU/p6rOXJRf5p+m6P0s5ekd8AvdZSsqy
qDzgl7wXJiVXtJC3pESSqVc4LFcOGuSasp3lu/SaO+/1Fv5gVlN3wV8jCl8R2kgK
rYNcopkevhBYCHbcnnwlT6DqafbohYWRSMyT7EE41JTJsWmrYckOh+wU4YTdNTCD
u18yOwD4YGC2/Zxfp9Gy2LEtb24TbGUuOiSCf1Lh8DG4xgn+qPaJ2L8GBDpEP0D7
9+xASWbvagyawnaH9cxscyEWLUDf2382jyORDZKHsNFEY3hrb6tgwLEdAbEYut9R
n41SoNJV7B4rj1H+KS6rfkFccHqIwPC0JAgG7cLGPmwAECHyebuFj21BvOSdXxQW
bpSc5kyThiNYX6FLeiv7At4uFQYHDbTh9d4vcfVYhrBvin5UdX3FKyWeYJdwshoK
B9KzYuTWFACL3p/v3NrRim9qNdj/Wmuu92bM/nwDykYMym6ZERa/sE8wAUnI0GvA
fH5A/sjFZilogMv3PMKcx29vSpyyp66RaFLxgRUGndgzwgtG8RPWrkVYjtQ9hH6t
tAMPWeaUsTkZxLDgClPZPizrUHk7hnbLraP4pejeCqfe3Mw+wlDG4IwOQAcqIU/m
EJU60e2H3MGa380/gKs8fLie6JQAUsmOJzDf+nT8Qv5bi6B3uhi5nuLXGPOM0OKy
UUPaob4kIQ1s5vGFFRhVZ2evLvv/XyJ22hm+aUpE8QZOikCIH76fpoREK3/N4Sbv
Ud9gKcpFxdaQpeWPbsf4e4vxnPsqtkBJPfAkTZ9FDBLp9o/5dW3tthxya/NPaGcT
eENRg7bWlknOr/vvcK9WjAiCL8mofrnb65FLa6eCiCyPGlUzKOiaPmGUQgH/djmF
/MDztIyBsg+rozXEJeiJHI13e4gCqfPrzdcd4G5xcCb0WWiaIcB3TlIsi0Z/n0Nf
1jP37YGPo5QTB3JIpYNNuq7Vz8XfGty8QZn/oleNKamdeN9kDLOQ4lQIPaT5sKd5
od+/QBSqBufnpaTarUPiSfG79uG4GVV4gVWYHOyIaIxE1wPTPQ4pR9cLaad+EZvX
bk0gG5X1zwpabOGSTI2LJr2BRMwdYdoz80mDofOawYn26PzJQ6XGAm+4y5Ws932O
ppZTDY3BeRLGaYPtjMkRxjriIVCrQtBgHuQ+JYNSHQAqXo3nEDj80Q0RD4SVj+PG
t+HaU1K7tD1GQi8KLVKmqHXIYF2xzydrIIs0uV9XiimzgHcdCaZfyKRfMRyKv/bC
iwwXHuX1bbOjVcWXmZgxz6loZOdZukY9R65k5zU6KzMAFObC3O55L1c131P0m4MB
TLC1PSdVXmdz/hMd3d5AG2PE7ebZ1dPgcu3oOAw7U+h1a0SUc7DDN3ntbgxht/U4
DnB1vZnAFKFFYCxEI7ed4mlYbU210oXuNkNOW+XHoq1DuTx6QILwbmT3JEb3aLui
BTCWJ6PoXzlHb+7fJeXzH1BuwEOZTDKISMqEKZ3WMHPICYjMmb89AaAcXxgrdcyc
eKo4roEQqlc8TDDoCNkIzOezGJ3lIL53bMAvnkObebG8KhuuoQTdMwlO5ws0/zN9
HMqOWgmaW+/K6ScXMaKoLIBquvVONdcKdyK4pV72szmsf0U0UOhpEgTEnw8UKng4
GAOx7BsB7DwgS7TDp4dZED7LnqsLfn8hl3l+y0wFTDeZ/Rew3cdD85FGhKVDMh6a
N7FSgmxxck2u4mAgyNSY5YVYIdCVyI/N8DT1B2tG0HrMw92pnvt1lG7bLua1+kXr
98M3gnDLTBGm1eYxxu8VgCEtBDMQ+8URfUD65P9uzo+FcGZuDm+RAMZqOG2CxHjA
Sg5RBnuRCsI0QIEVnLKHGtoR8IQGEUd1IGfUaBZKNKN89ykfmWLxnLCshmihL6BZ
f3gGO80ACUdlOIxMspqJphyzSdwoNkAbF7gBuSHoC6ij9oqGkEKuW7kNzvQ3H0Dl
QuKEgLS702o2gvQGWUmsvmYbt/ecrst9xAFO4LhALxTUZhztGgIiA8Mjy130A6hX
WlVtSYOLBRmk1/y5OROMA3AzVFqsMIH0yDuvRrKFiRceQLa0+HGG6OA14lY9Fw84
pygDXjlkjqOT/p14YmkGKZ4vpTa1ZnbcIaC5ZR/WmL48X8YT/1zugdRAqMLNqwIQ
Zup20twSgr5z1QnsTnM8UkJDrDRwCfmSAZXyUc2PksiGEf+lFrfwBD3gdq0B9xdi
qcxeb1CU37rDSPe5KBlsoX+VBu8jHu6ybGcLLOW5PAJ+SzTkSPkFjNGefisuy3P1
Q1SXCS86xwlQSQ2sL/LqCWwep0IR1pTXImLzRjinyOety1q8ob4ych2cAzafwZGY
JruNAxKAZTBmFbMGB9Xy9dCes+3zf6vJesGGEG6h2r5neud0tJZhiTu4/H4fupyC
GhCczjCp1NKihf8U5bHlmp11FIV5DqPjpukvX+/aNy2YuY+0WnoH6Gxa/8BoRKmg
gGw3DlSuK0w0NU+owHNL07w5yj7vS9FZ3f4n8d+lfmF/j/RcxaKJ11RQmRuRQiZ+
nXbxBnuOIYBG2EDN5MYHie66BrXtSkXoYdV6wjGS40DLYVkCjiC3QTTUtgn8v8/C
qnmiugwp9EorjGleZMo3s2+Ci79LdVUvph8+7wxuDZnEh/CmvrDkmUAsonw4PuJy
RYlMHFoxmvXpUrlzm0E95Iykw+If/F1Tuylmc98jZfVrdzlHlFP86F1dPwDUQG6b
Zu7Vr15xXtl+jidxOkVnr0DNIDW/Otmmh+HDnTw4pZXxlQHPMRjxRlLDuymeM6AO
trfbl5xsH0uCUlliZeivd2w/Aq1LBW5PdMBRk49vO1hf/Q5yo8G6grHQj79lO/XA
rEF/BeG9/+XNOACsVD+p1CMUWieH+MHwgSrhT4QxuPcIRgjr1yxXYtgxaV0JeTpd
q0WIGV7S/a96yTbg1JB08P7Cly3e0Dstlc7cRHuyQ/PezHZahCa4Xo7HmK0k6pH9
9mlpzXjb6aUqKfPTWrqXmmdHLLnOYjUW84esu/oIr4CloI8BRdaM3ILuzaRl6A8N
iSiEq0I2lE5fm5XJyBjst92Wyt29Lxv2zHxcPTWeW9oclnDgh1i1tt3TBIKTOx6N
OimWjMqg2BFT8IFPwKVwae+YHONEOj/9Bygi2VALip8MEeQg5b/L+rRMmOeo8/FR
C9ZJnKoi11lSw1krlINwThk+pjZJ0lBFlAjqjQFlS1dp0+ERZR3+51v652HI5o0Z
pQtqTd33oJUEgMtW2/7ohYiByQ7NpYxWoioxo2tA8oyQdAgQvVIn7cK0EcroXT9u
v6ycnBEjH+RqH8NiVKhCi7WDc5xTcQXmAK7cbV8enXD4DdEr1k3aRknm5Mdhafrz
d4UylHrKfCKVv/AD1Mm8P8CsYOK12ULO8zwmbgnIa7zANjJ7lEDDonwd5AJTz5F1
ytcxFeCjvktlaa6mIbcArT7dpJSaqayzJx7yXLf/n0as+Ru7Z92+/nPJAIf/4MQT
2DCuh43QJvl5IlLq9E/8mQjBODB0l28/PIfXWsZwniF8mN9vOOW+gu6udkiX2sFl
SJEozmMxdk+m1HFyBQnAH7Y1lqw9dhrEh8h6yZFNaVdhP1sHzi+jql3ZkG7cNUva
2Fq7DqnUq4OU5mmtpGC7AgoceV5kNh2dLZVYGrLJgfDrvt2DSqREXL3/LBl6+9F7
0LmO1KD1aYjexhJu05q+EbwhDmlkv+2pIokz4D/YVYyC56XlONDKnqkB/cjYZs3h
8k9n234YN90nJHF3PJMA5w9E/S4vzFKp4QTQsa028qhvIgaqteWPHxi+YssH+Wyl
Df7OPKxBNj/Gc3fDBPjDHPLk2vH3VvaDsTuwtzOSZ+IAMWnYYKpwQ4FYrcFGYDVD
WZugzVNf+u8um77Yldzwwvb+iGoa+sslt1EjmL9W5XS1jXdq7cVanXpG2IKrff5q
v79A4zHfDP/t9JmFc8qVuNhJZSBMw59HqjK16vtgqPrUuVrkqadBuJaSzqK1b9tL
mj9Y5CE+L0pUEAFfEkXmPu3z8kOXGD5b/Ews8rW5j9i/qksllJDrMgVE1q3a4geE
RYTAI+TRFxG7XuOHrOcxWCoahKBet3rDa9O37b/UQQO3iSUc44hHvGeyfzvm7qvr
FPoxbgYrbBGdGcscAHJdm4ozmtKYTjRcbTnKGFq0toCe/PlXIC5GO0KmDYL55ksa
sQn3q9TO02P7neWKgrm1f2GOiK5WwrX3usBexMEemPjVnLkbJXhyxDecXqtz9Ke0
szlWZEaFai+aw8oYnNCipybGZTj7tJnkwYw0qRyLN0dLNFpGQ/rktffjbG8gf5ck
ruaGGVxO+FOO3ratXlp8MJLpgv1obHEotA1C6tf06D/nFJfB1luNyBQSCH0HOXP8
hxszPQJuc2CnGQEvhTmV5ZF9lDV2epg2Cc2BGE7FplQtMPOCgj8NbLbpk/5HhEIx
mwfJUlG8Tkj+TP2VwjL/hwZfogDlgTBfD9ohw1kbY9RnJZLNXPPRKkj4qRovDIq4
pH8zlPq/129Qf4aRGiLXjnvukssTow1VE1+tWRDXNZd766wHBvdd8XNUpmo982zY
ORhUx/tXc6Po/+ZzdWqxytHV5uFAvhpZjcOZu7CLV+9QYJsNSfNptdPrQsHcZAqt
7j3gHQCRIX05eG9WrSLgCg4GrzQtmjqVG52M2pdIo7r7l+MLaGVwGQgnDqTe2dNQ
RgULR6RIJg7iIfIe9oS4tVqDtxocOycQbTK3cU29EoWWo/BiThndVyCUoZIzntei
g+69fURCJWZz7fx26JZJaVb9EmC2yxrej/XeodlroJvCMGsyVDpF70hoPLUGlfSR
XxBmViPr6YE3agtSp7YosbIXs027lvLfKoQiCU9DCgew6IygGPHXmU2uU9UHe9Nk
A+qY/E924eQnFNU83tGmg9c5zbg4dwEbHRUfVVV8ntenuApltGWdrYLpDZxZ8R6f
YKAMpMfh+wyjmNkb2B0jPNYakEcNTxCs8I+XF4v/u1337fw7NWu9+Uv6Y2pvmxnj
ewvWL43rlTelB8qBxy3bj2iz26KekjUL5CNRHTZszsFE4kayBcPKpo2hXptwZ3ih
AGrYP/PIZZNeXcG1b/Ce3XeWZry88XFlKLUnng156ALrKHFGUlg/1svs7hJsaZ/O
6R+1TLtRzonPYK563ISgCwOrE/mNrx1JImdI36EbFRNCzOiD7+HoHzxYjkt7Yesh
r367EX6FKFShIn4GtjZ8v+p92vAoZEPYNzjMoYfwx2TmPl1WjhCMzdc3MaJ+xQUq
HEgrnLreSNpZ1cOnyC40Z51IoIJIoVfoN4FgAFApMbTRaqJfUW3hsLBcm/IO8b6i
/onENQAmrJ/T72d1KnP94iAcXslEfcd2lNfkOv6Xh65WHZphNjeVc0xCEyhYUjYK
HWqe74nNIU6ZZKx+E5NJ4Ee7ASRLiXNzCuO/HGO6CNiFPpwVcB7w9+yge8YSRBA6
CCGz+HHBT9CTemVLCL/H+FYPMSSu91GT9afe+roj/P+xwpOozVNEZBUOr95yv6PM
M95krWgI6OoWWGUmEYfeOdX4A7h05Y5R2KN8cdJU/n+ltq19S/L8Q0Es22Cop5jO
kZlLXxT94LLY8l0I5f5DTocHYR4G3Kt8bR8c8S9S3ENXWrmvx6y8q54xAAaYlyqE
qRDgvaX+qtDi9n7Y7kZjl0HLklMouxtxBq1FX5Ba8GRRuy7olHH+4/2iP7xdy5V6
oZV8jDyt+h7dKHOKiGJ9T46329uuU9ovmLTwDi2/g7OZSQJ3UbyV0CIx5Vr+uJFu
iTkXvTjjKXD5vLWGkSvwCYHe7L/jeYMtctJGBOGmyBn7GvuI7mK1nCBNF5xBZUOv
v4ZFFKDXs2YOp9Ac0La1Mk3yCTyLrjy1oMlEChn+Rd9HHgghb4lEKsBquBaPjztJ
TXK+fV5Cqpxo8qFX1h6rlBHJtFv81zD24SmrHXZ4DIwbBb8mPLZvCVy3DfKWqv5i
jOmJOTdOmPu1a3SvvE2ZZiKlMajsV3E9Mod4zGLloY9x1L8ZW3F4Nfr4E1zGZKch
RdSMbJWQhdMBXKuiH2ZOIdwZ9JjPKnW60i+FtMStEqY0JPWSecfSDCHp88NZZOkQ
BMl5PPhhy9o5PruYgFaMoOwvyQurbzues1653HYdp1jAXUwPxn1Qnpbj4a3L96up
q1EbUuhTBzNXhEOylhVBK9zt1voa51Ex26YdlRcEUqro8zmdHwFoNt95tcMCKRnL
J/qItqC0G0uqiLza1JeYrZDRDvL6+XQUsZtIj0w9HRimQAx1N3oljAH73Lzx0x+P
MG3jJpZmivTs2TCJc9cohnG4ylaPDSWs6WHPPCp5xMAO6y2qdlHvIFuzVkb6JlUJ
RQA+NwaxgkmF4ft/7uiiO1Rj16ogGBSEUVmYawnPWAQe2TpXxkXoy2c7d3HZuW8+
ZEPDmkReOLJpDIQutVFQcuctZrejg7YOoUQpzQhd01QaPCgqcV8Z7l2G4mVI8dlX
LOTUxb0nhqfoj1j/rfv0V6sKyBdHinFksSQq+bpP2R5BuyEMqE9ahObhI01sDRFQ
tD03GCFV1d4VMfsiB3euZDRAghVSf87iOSgY6IddiWGgeWK/Td/DSwijBHUNusU1
OZ4RDXAYhM7cWSK3So6woDhQteAJ2JOEXbZ1bORc8Z3w09eL7zbD8MzF5CE2e5H/
qlMDAqKuGf9VWj7kgkBX2DUWw3zvyyPljcY7wv+GA11rqcdX071463p/gDJRorEI
3F4xvVQFTA5c/FuBtprt9acjKA5F9RQvbwOyatNPKQ5e0k89Auj9n5Uasc97tbbo
lTfI+mxu6j9atWP9d3weasBl5L7IZ3le/zF0ucb9SYyaIs7QS8YRsqxCiVSYWYm+
UeZzNp6PdUJtXElpqQI62kc+6PoPsMOFXYJhQNwp3UBIU0TsTzbAgb+Epaexhq33
aDFZtKS42NWnkOVFR3SL1hYXPnc3FwLOnU7dVNV4wUiiBAtjYXeCxjKj62KKZROK
7h+RgJXSv3t+1jVKwyFUJbH721mB7JWqaay4CuPJRaMlz7mq5NMmAy+zWoE9UfXo
Worc8uIb5HSeQVjlJB1WXAuhYQ3qL2t3iFFMIsVHkgN8XjRqtvpvj0zPCad8ALnD
OQ/ctjoUL6Pl0gTQgNpbXiwFVqMFriz2weaTIHRgVz/OMbrM2L/lHGXmYn6BKiQ4
v2fd3OvCw98WUpsCZkbO6yI42s3kr0YPmsFKq+6jdOkEcvu157qNp7HkRMb0Djso
I/lCm+MqM8oUp6NeK/WYMekOn/0z3xfVL3IKS0u5Hpe7BGgNzgZRq0vdTWOOONFA
dLW8HNIqfQpcPoHWEcZOlg==
`protect END_PROTECTED