-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ON00vraXdseGMhIU/HVDdC5daL7HT6sfnxTZXfivSOzqkMQ2w13xtbjtHnzEkfm0
PHAKZXFPHg0Q8Wx1vqlWFFA+XhVcgWqs7mqGsGbBhYCGXAVl82OBiJ10Q53dUMZe
6q5fyMAiAg5pIeBGJn8ftjEQvpwJlewjHwgPqzqmiLs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13104)
`protect data_block
i2td1cD8jogZHp5iQu8j0jkjtzA3d9D3QEiNxto4EGCe+PtiS560q8GSsRUxh0Uh
rpbMVU85jIklgocN/DJscu1WSb3AY8K6wZxX/Er12J1hZwynqL4XGupNU14j9gv9
wtyJFYQKeYoV5qGPBQq3ZtTZ/bgS7Q0S4+safsS7SCnwfC5VJ+yOC/or6nz7Kr2k
3LJWXrpBhe+qPRxPnaM3zrOZMby2qeH//bzoy+cUk0x3jipXwAXIDV3gP95PXCzg
ZPfDGnEBx2eHIuGoR3GEIvhly3MeLisYQBhd7So+LLj13xKez3/BJrVSfV1kKsxN
0AlkAE4fVvKOtvTaw6CVUWQTBF014Y2hV1Xn/7cnXK563HE2pDQ8uOyKFlqVKwnW
oLDc86JOOxl1RfO0bs9L7wtG55ybwZeity1uGUmm/OO3dZxKDorS+GJQkxWieg8E
5Z3adnDLW32xOWdXr2ot6S7G2/hWelNE7b8/dlWFiCZePpZdELjgZpovobjC+gJ6
9xLtkbOMK4X0iqV7QVOFUyzR22jG5GdKS5pvGyM0uIGRP784lJMbOFS8ODvHikte
EcNjBzJdPWEWWgXpFAo+EEtV/9WEvj0dXuJPHJvCsspz2AaK6RD+pvnEOGWFc1NF
qT3aJ6d77LNTTImjgwosmW+yvOVYjvYBRz5sag/j3QjeEUdkgeawdCS/O266qsvm
a78/b4sACwuuALQggZ9ayYvbyKHs30KyFpKAkwhlwMjsEHffDcK0O/xYP6+vpUfN
8Z6u+48a38UCUl32V1P+D5miczJBlD+5bU9O2Vd6jgNLGUn6Tgzw05NYvmb3Htgn
WC05lf0GeBK3wwXfPr61mqm2h0BoiYAnooCxFkkMb1/9XgjH0X/X2Yyv6uJRA2Ql
ZfOrIi002B7M+eTnhbOwhul2okyblZ4tQogjuaVpURqI9MRHOrpJ3YmHtxJNcQ+v
xJFtPz2VcNbirg9EK5BJA2Nwn4QC7qtvxwrtgoa+s5NNXZSjQmyF0T3ZlG2QfhIi
KREO10y/UNK5j3sYvijaBeRgFskAVXl+DDhEmir+6Y72BklzDmeoPyoKEGAn0VrC
M9Kj++bH19ngzpJysHqE1RYKKnk7itmxKzn1iQVrqH2SSIiwlSzddg8wFcMavw+u
WdVEs4wFvQPiqtIJuJIR3chLhGaXYyfAsjBS87pqPzCVe8DAOJN/gw5PhaSeAFS8
dSRPndaLVckHjHW2rcLplzCEJr17UmwS5e12m6QQKTdIUvaYaGIyDQoGoAhMaxAk
gDDwApxQwA1Hl8CUWRMV7TyPfvTV+J4jXUYvU24S01zbdOioIwiiMfNgWSPNvP9J
EUttT8JAuK+dMYF/PFPpiEENK750wQFC7LPSaHkY0vvCcc/gTjygHWBifUEEQLgP
F7gKFMTr/lGmJpNDQ+vFrhYatY/jwoylg4t669GNWBrTQwj1udHZ8E810mgNEpc/
XGuEivE/qPH+6xW3S+kNw/wLaHKgRoBX6pJWSuNBJnL6R8ohDYJVOkGsWPF08Jwd
ODD2wyk2+iKq9MVsHalsy0yQHRLIe04lVnKNBeK2r8rpaZd2qZJirKB699pRyEhM
G11x/kcR9qD5XZH+ZkcUWwf8Cz3FrMJ+W2MwDmRk6Fqex384Kk85I7Cejxy5u9sk
08XOccQfwDUVp+HWBltIKTe9JtBPInYnMKFZk9WIwscBaXvYG/VpsHd/LNdQLBrd
xhThwEqXGTjjdA8ytoyis/QUCTi/PTvq5b7LBNcpq8wIp8JiSmZhamg+AYhiJ0Ma
E/k3KETYAl0bFXRNksTWGM7svf5tWy8Q7fpkWyjpnllxsbtaMRosaekxgivh/s6b
IZ+j4ci+snMFu2D2Amq6Lg4dHgkLNJmxTKjtRngIofJbP9RQdmCblbkfCjzBCOz9
0854s2W65/01PjajG+nm7y4p9A3deYgzcNCu+iPWydrPmCeB90C4QBeSSQwzgZfh
SN4yH4+mma41btibWhMnE5yIe7qcinKf3UknLdsmnBzL/ZER5iGQ73GKCE+fllkX
+esdzROnyJzCBzjZudOR9VOE60fY6KDUJ8trL5OHLqoXjnuA4s4vG3LC3Q9GdzRf
+W0EU7wBdAcwkLJ6uSnF1SfMzX5DaffJVOHM78krkJchTEeMS30fgaXkxR/8VYHc
WoX6NFeIlIsag6ucw/MIDAU1GXtBRqJsUQSu/OqjY7bZSmNKWQmRIek7YnzhXASp
INV3MkaB25Vm6bEnbk4U/uKdeQp8A0iF/yGRFORm3pR06RQQVi7rTx/pb4fmh0af
zRsH4bxXh6MVOh1cHytEQ0Y75CxjfMwAnDSpKKz3Yi0tlZr2EMZFH0k70rYaiNTY
t5JweW+zBtDTb1Sifv4dgqSD1AI5L9MR6WWB1emlXEATqsTr7mswzHqQGnS2B93D
ltlMIpt9gg/aKoaEZIrk79gjwt7beaL1pWLU4wxz6E5+JPDlSmBYx0PpWlif9dPo
q73+r3BR/OJ4PB7UutzwfPHprOX6BSzxHH58diO8yMV3Uq13pGErRai6J4/JPUCd
Tn5yj719QhOEWK4bjxDtSHdcjn4v1hgT/lwHUqF6XYRMfVuwwwBA8v5wwirxNGAT
2C9MkK56xiquBhWZiKI8ESGwRwm+g9y2mmbWnNviZfPPey09sW+ELF9zG3WQgy/I
ARoNGkydgWa1ctmgE0PY4AHriwq/ZbrftiHHJ9xGHa30hOWb2vQ9xr6EWMYQyyjl
qZy7oX9OyEc+baLuEifRE0ekQlSQ4jfGneSxIYMB3hQZY33SEwo1+oEG2f5Lh9RC
lq46DxlQR0tOaqbgvOPq3gKUgnbXxdXgXdBJqGENFzvzrDFOybi4l0REGeWgYQar
KMI0VbQGe4tf5CZxo4vTpCagE9CkNwjZeqcEx38X+/4sPGDDB1h2gwWAIdEH2Mec
yDhH6xRQAqtK/I4YvPQlj/q8NPNE/jk71I+1DntePGiHgvSeTG4zjB1kNdbf+JEC
uf+/5J27+Q6z0Xp3uy5werM+Wvz9CXS9otijptlZ6YFUU7wkYcu1AMFn4wXcHSqA
ZWHf8Md554rQPhdbVJVI4rBymBIIThqC86RjP4OP7L5H7y4hfTbTVLCk2j0G59cS
onTwkP/lZIWS4PFhlbt3xyLIG/tqDke1i81sCdxKCSbpp/ahIiD3mZwp3CpACDzJ
J0duoxIqCHhNkehmITFfR6uRmweVHGCmrSj+PYg5+JrlJ97etEnwGJDtqj7MVMAV
yrNxBRpkMDoD/P+ucCpVVKHDCQXAAN7rI5ikBFP44QjznQFZqaOhbBjUda+Jiofh
dKN4qrm6pUWXgJLYUVa2BXgbvg4TU0DxUo01KKC1QHjXoqzBYA0B3HGds7NukMRE
tMAyDoJoLQz0Ed1zLwN2OIXMryXxaTpB2w5+18EiMbwK9kbUFKqGM/dDnUPbhsL+
MNsUwEyAV0HA0pTfeeR/qsbprn5H12CU8QBUAEMhsnVXNvu5Haev5sSnaV3zAfFu
/w1V7qdIzKfyPOzM740mkWeyn8DSej9A684USQnXkfXqcNYPqFbWrcgHLTowggoe
wPQu4V4SJdLDg4n+BP+wSShjG7+LU2MW/oC4k2AB8ITd6pk/HWJ4P1v+vVVegSp9
ugbY9HPDX3B2aA+OmqA6TJ8hnxKvUx6PIRowOdZ9RQYZfQ5rxd0Ozr77v3sRVuX/
4u1QaZlCG+6ne95kTFg+4lDcfWrdKNDmrVbqDvOsysXVLLHi77liKIzKKsN1y2Ii
n2+b8YayTOESh7rrf6BeLTP9hhTTRmXCi65bUWHRD6SWgYxDzz6tdfUw7UaddhUS
Dydwk7P52SRh9qdwsJvDX+fIuDvTomr5fqUl1pymhjfiGx3xfNbFyrY5gTYhOl28
7+KSFFE57QcOAhzyvXkLJk+gcU4FpOmQUCgANTG6/AptBkMgkq9Z9wvUBdLXBvFi
q3oMW9R08I8O+1Nn4EIgIY2NTBaH7TCwKVeX/zBoBzIQ/CkvAuDyMCRQzHHb4FHf
DlSOqsfbgq77pSZeGAij6EBrgHNBbO6S1KaAy5a1cJh2ZH22JuGrNn/ock1+lWWG
kdee66RgxtzSAlwkr6/WO72ZlKGLUqgGE56FhQs4tTOuf7cfYqlVSMoqqJMeO8mB
L7YdkNTcGp3MvYulIuFJiG79XizBn0moHa+VhftO3C1zzFOny/2XQ/1dmLrmm/ws
k5RtxvIs2vIDiIRtJtZIOGdZGGvPN/0mE06V/0J0hx85ri/WO8uF0uWk7fy2eQBy
PuUh2dlANVzjqZ5gLCRb7u0U6JHGKR6EVVwy22nqb8VJL4AXD/yR5Lx7KZGtUj3I
7NydqIkzH3qf+zgc5aRZYrke9UQ/NqNmLHTU87sxye6aKxPHk37w/RVZTMCvbdIO
LqHe1vskKeFJm/g1APkmafC9cq/liUhL/RuifSPU1dDfr6WV2mwYvcGQXCJjgApD
ylGuADPvkRxBmkPOHTttfPqj7eKHcBh03RK8fimOR9IRB+WCm/SlziQ7k14k8HZ3
A4uQzvkjB+cY1yp62U5heFtW5YcVdjSLUD1fYarTPsQSDevlJ25UFue/ev1WXcon
q4aQSAlhbwRo05IvSm56+3xolfMBeuZsR2TRJBWQ64YE/PYObV91hcuZUlBM/0rW
JQSw4ANTbpdZsbnprc0Q9CwW4WInDufzm9PsBSwRjii1KjD4k54lIDjkJlclhyHC
y785Xgj4FJLohKx6uXKiaMEraxoYWTrLsawHcOApCMVozgAbjd0Ns9WCz8B0d0Km
LOHY+qOgMjuwZjzvXZ4HmqnuQ7iNh5HtaratYSN3lnCN+Kl1WVcL241ugKcFL4/E
qRg+s4Jk9CQolcvCHU/7A0YxI8a/ywGEM87AUWBkI5h5GYFr1TcA47IW8PwJhFBq
UDBozjI1NQK9akKrO71i7nhOp0vSbDVNjhb/QbonsIo9MUyRaurHQwIyDP4dyxoT
l5pXiQEeGDwse5lqTh8iyhhuNPpsjg5TigjZvQ+i87pNOjDLkLqCAN49AFFSflVw
tapADmWoGH+MElfz+jEzKtJ40ffrKHiqHcV1R5q7qG4VoKjCosU4Ksx+QF5L0Wnz
/Ml7QXXokiqdxczD352qRkQfMIbPpqwgFWxHzeVHGbJAGQxDByQC13WjMwF/p4MC
4Yeou0YJMyVzop2POr3xT/1tl0+mvu+brutfzQkCfVUUitmdjiQLuwoNNbrCokmv
NS1VkIT3T1gt1OBrXCIClaGXtoGfiRjoo7RVJM03IsuYMEaVJfOlvNxzol0sMmJx
ludaFoLONknNLdmlUSGI7aB81PHnqcTfwUw17UnQyfYga8lGAjCQSW8Vm2sTBxgT
eBqKmTCOoiRz/LlrgOpp+V0NUVvc6Y2e3zkpGZPT/BxjUR5G1gQjV9NVmSFj/CZ7
dL6Ikh6ksGBcNoUHHrYuZ2cnKoopPeeweLh7UMnBPuPZ6u/4FT+luSgy3JMrwGLD
oIniYcCugFFmLtLoQpr36j8u21i9lqoPIZjaQCP5U6ebK6ZXggb9Bv3k3oBcFWra
An5EYGTt7rhulwnl31EOp0nlP+4h25HDEbBSb/AqlA6zupU+6QFVeU9y5zg9cZ12
tMmXraMLvCdXUG45gWnsW6ufFx9nd/kyo2PtuxJ592z7bk0ZnavPNU2BIxYtFwXY
gcy0uUffMGlfiql5lKB0wwdLi5CNOF6MJN9VXswkuZzkpU0iUfZEmAzC2H3p4QRU
0ea2LLkKr3soNS84kzT56ZQ07o/hl0RaXob0DWhgC/8qawb20DOTQkOPa/SliMJw
VL9m8giqPV7pzzErvTg7njTCgX+YbMLExSReZzt5G/Dr9PbHTvPtaxA4Ho5JaDW/
9hkYOO4GkMtFuxasZYTRpxtRIpCWC1sAnmTHTvNViTHyr6bYBR9hMVTLiQxPuH+v
loA7nUdYg75VGnrNcO3C/aNBCNpnohOo+Z8WcXJFTFGG+1RUQci7u4Ys9ftq5xEV
H2OXGWGha9pOoviNikkLwdu9tEjtKOOncZ0lQEkayMRgOcAs2LlyKbEuEy+GmnrF
eoqSuDXhfeZlLkvtl6FQzqiUffcCjfMLH4H89krYXliNAP31cdEqSPisOLXuUwXI
ms64LZn6NToXn6oNKezGbKjCXwCxtgRB4KyPUpix/J3A03ZRPX/eDEP9Hiarmaj5
El/Gpp/dm0PQRQY6CxZ81ewitRzSw6sAJyrJsduOagljV9PneF9GY8B/VVBz76YO
CUDURCSY2lRwdjtxuZu+aFbS+lK70Ir6q0WY/Cjfevw1w3SnYSymGY8fccZ35YXF
BVFDNRgKIfgpq8IhywmjzLIzyhkwrSLzmbHpFEs6c+h/uArjh2xPsrLU+U52YBZh
CYCjSVxO5mLyEm+cBa44w/AT0q1eAMD/BGW1FwEoBcZmOYlcSx8yv+X7QHv+rOxN
o7upJ/+N4GGXZwal5J3ALSYnLyo+XCWgkXp+774rcGXiooAr0KgeLJk0+tTlbezJ
9zNVPGkd8496kY7xRQ4BRbeB3+72NXMShapM6TMKFkSrSpP6E8pTuqaLiztbsVNP
Zcf1LIQ4tr7oVQpB01FN46pVRcNTKAaRfYGkGZND5HEJbCYhgII2qlI3cp2+gY8b
LVY6abcS0JXKDsTIdJHpdaMcHs7uq8jyQ85WjbRta8xHQq7KYAhbC0O+hSCMxmmX
Hj0kSAgJ1nEAPXdAxQliaGltOGA01Hdl+6M5mhAdudNgDiJ9yVqOWEdpcxUytRNv
vxcKCSujW4LY3k4o+oqFvWwSKYGj/1/X6EXypqiox6wkurOzCJaZznpfHTfdWZdq
kqbC56pHkcQSockQyArij+eES0G94OW9WQtmMtfFq1sx9oebUIjzGczolWs0kNq4
83XyaSJFyCNpSetnu64unujoiZM/1I2qy3QOl0Av4+EnWSEZlzOo3hygJq+VOfn3
NcsGiy61swXLj/vAAUQJkjbwQcmtmwOxs1iByswj9QazGiBnyNqzMsGsOZSwc0Rc
DU8oRLvve47yf6R/E/zJQtm8in2qIMJORDDB2oZaTAQrbf8elxDlMRbb4SII8VTf
v2R203kbDfEeWCM4/re+Cup7lH4YLoGOrSAMVvXZTq4O0RMqIGuFWhIISTN6PIHs
2bj8M7HWVQb/PMhGkrECBckC/ixIYKXzIBFFAInAVaJA3ML9bmwJuX8zmYUkm9Js
zPaw0ZIgc6Op94rrsHBwKILwFI7S/ee0L2inDL3jkviBK4nCSUe4T/nYGYTIfJsi
9jf6OMxvokqX6Ydg4Xce7Okzip2/dA8fTrtm6fIoGJdAtLJFw4OkcBNqLvc1AKwU
Y0THSzLDuMB5mgRjkTDvw9G4Ik5BmocvVUT4Zza4Zgt4a/QMtub6ndyDmGCZeATq
w1uyMAlkzoXd35H2mW8tMveHIQ3GVKTMNlV+k7l62f98QlL2ZEYtS7dOJ+v46TAy
La2DIVfOUCy2w0PVFhX89chiFg24prQuDf5K0hwkHTL0HDpwDh+5MFROIKombra2
7LCduZsC0cEDqKIrz1pDECRBFjlgrIuktmBz9cKX0FCBfvFEIGbLLxyy7XUlzHTk
5NiWyUWjSYyX6jPtee9jtyNbMj3o3LmZ/dYUKbdOhNS0UJfLOx5cQgF332I9OSYN
fQyn0GC7njTbHgiNFLz2kX7dkflf9Iiq7hRXifefRdnebDDOkETLzi1NsowLN2Ur
fnmBSVFpbsZD4TtT0C/I+vija8h2Cnkf77KQA5iXQAawtkbhajXM5pscI9XRDH3Z
Q2dsz+K6bzaBgJadYFaxxi4uvgrkPKNvfKZ1Bpfs2wJ2xOcAiyKTlGhyWNfp+IdJ
s/XK1/f6ar9SPUcSrnlsVFdKBrU64g521v/ejtWNCEsf4got+B/IQnpkr87SwUOL
/Ke5IS3dBCgkiszHB9htW0nfT0RQlXj1hfWKq0qeH839Zqu0KWL8YBOilg9egjFD
sKYD3UcnwusQavhyeCoJldk5pTwNTdspO0F8UTMBHRpSZKCKhfCgFXlaUfY4nG8r
XCnunhqcJ62dkbp6NnWKwS9/i6KmwfEvS827H5uzYLIHLt6wKxYCUw3E+ayHuGRR
ifZiCUk9COMdiAAg8L6V7nUqiQTJbjCmH91NllPz2B2mZIVNzaqHxIXzMhrjkKLb
azzIcC1eFvDZCUY263o+SVqCUwq36XAiRrJhxcyWg6Oy0HZPhRU5s+okO3+UGcNB
UVgi7uEsWri3r9zD0Vw3bf+GVuBE1+39WxshQLtyjZb2O0McXF2bJ93WYNXw1kny
wQsZKCaROw5Ytv+ZMWV/CNA/iv0Q51UQfFvGqNrwA8RPt2AOPqyaR3uhlbJW9oqa
4ia2ozdr0J4bHVLhXgw9Kwf60NFYIDsKGNnJdJRNIZ56Fy9Y9A/liT13kxRh//sr
aPUDeNe/s1qP0xaQLgp7mVahjj2YvRGGDL+aph+8xl7JKDV5211CLiqVZs2irXHA
zzy2rGrroKptkBfa1ggkM6BW69Us6SYin9Md7DtNefukxpmJsAngYL8XPVvIMnNz
MCWHILbMBd0mTqSU8myCVbmJZQYR3fGt1KeznmyaPGobjjE9esth+sXIW+jzAr6A
VE1bAH0kVKLAl3BhrqC2s3F/ePnqfwWG4kH84116nYX7ZOXSSYg8LAhpclnxu5Q/
kgqEsUmx0E+4BYbPds/UTVLji9P9/kRLkLzhVegZMsxcxfxYdykq1oiP3a/Yk7oD
yhtkX17cufRcvbwvxfRiPgVUax5TjC1vdfYwfkriOAsianO5fwQhqbEyS97vH/dZ
FoutbrJenyKDRJe+O15AP3hRRoS/OMYcLOnxzkgGPWIR1spumxLx3DXkCzT9Fzlv
btr2dgxlGaZe2GtqGj86NdmTHC1zuNSKovIkYjk52GJ7QKv1/tcTKa9RZc011T9+
dl80i5g37oKAOjPYxhNaM9vcXP6kJ6fBnE4g/mpvacQSjXh4VXo9WE00PhhSqy0F
JeG6oPPoJcZ4AOqA5oItle5wAzVtR/mD+GcZX936LO9W93o0my5LPV3Vzi+Cy+QQ
ztkZpwQyea766uvumMNIewnOXqRuarCXX4RCm7zAHPO+9rMg7v3NIaBPR2eIeAEa
34Et/wjIritkucI0ovRBuOKrrmILdTwgB2+LXwYbvv6f5QUXpFxZWpmGhXKZadxk
7UsJMUywTLKKHFPmoaVv+dBkHUObEqXjBAnbN9h5Nf10tdXhaabX5r756jARN0A+
DQsON8IZSQNdC2WW8d6ayofDfOqmrMkNmIdl/A3yKZ86HJTi5aSWsAZNJfShwDQF
uVr5L66IZmpOmMHDlCtMugrnJkCRkEjD2SJoJLE979s62bzBC08O+3XnsscHeEjr
f5wvXhSARNH6nIeHe2fNvRwvbMx2sXDfpNTkfpZ8mA6KxDlONBf74kWw2+RwKT8g
JPSq/jI8wecsJ1abCLSzKz11F/mVfEl3f5p9mRSgmhIOdGV7kMt+uy9h/8PHdCoH
Aj5XZpobCjdOCDcooBW1DMMbEGNB4ji1BOv0muiMwt2LMcZ7CAqTbILZkKK1l2t2
6AYn3VHOZCuJv0/qK5vUqCTSS17lcXrgnbmQum9Fornuw1CL3DS2/rm6iKyfltzO
pASBpwFoiF3V+a3Di9+4oB1/6yVZLbjn5hhz9SKqyPH1hKFXPvmYY0gY9zA+TH30
S8SoGMdo6hinDaUmErlmgdYeA2dh6Mhtb9G0tNhczmnRHcvlM2+1eUZAF2eY4I1p
abMGxu9P7/8aEIlo4gNvrKZKJ7CqUYIVzUUS/gd5p1qyv2s7RLC7RrelrV4gdATK
/Z8bILx11m7bv8oeTn8dpHb/qvyo2poJ8b1IZPI5ihpSDyAEqeIOflBW58xuKt4Q
3fFSVZUhLpErZ/aaobr8O+ZlLlqRHZt/Xz1CwJCAyOG5rUy9Xjup2Q8LBFXrM3/2
4L3JCiQCod3Ol0VI2hD3oAjD+b91abu5XZhaYEkMaGl2zB31/CA0/sQM9+OsyBoA
wPGGuT+lmPRogTnAiPix9F72wrBg8sbjo8dCx+bMt3+uh0aBh9jkSlbmkLKcRNCR
DV2qDDCGqFdt72FjQOGiQqgu+uPmbT+HdDTji/Md7oAH/7ppfYmVJrvqh7YZ6xrl
Q3X/cQ8xOggcilAGzGXBSwvz1lSDSQnbddHvLb39GSMVu80SVfAelrKxHZKIBAB2
bmevi7rMZnwx+0XEWHS3ogNekaYWA7vOBO8449RIGLHUC/+6+XxENOkxnCkGv+o+
4TtJOdL2ByX5A7/nVFChKUk3z6wlLJN9xzDf82PksT8wdWe1Op6m6ozIWHlAuLxN
Ks6ilDybSlYTQ3xMazWr7rSxxQts5iPwMtnbdei0fI/wXSCh/kWd34j8OkdGO0zG
CXTIPvKZTkTc9ivayo0LJUeXEJGewg8VhWAWZmkI5u48Wa9xNTnS+I2OK+S0b96l
LJesP1SZMt+IwnftAE/Bk+vu1K5TDnRfQyDjQ53AbuisjLcvhutxRC/QU9L3A5F3
XRFY5SUwPHZSeSXSsVWmqE4H6xS2tJ82KCW/geN0YD12ItytwYoEUjIDsOeljhEk
K9fVqtUqroe4ndgBG/u+aqc2/eU8mntqzchTJtiy1PuplEiHZ4QcfAahnpAFa3qZ
fdDPzSwug+fUwL0fT1/bME+xZyhQD25eig+COM/0CC6U0l4g5mcY/A0NSK9T4l7W
nfGjOEQt+v4ZtoNEMWWoUrX/REa8dSieKQf6o8Ve9zSLe8+NHSTjugpM7mfNNcBC
B13c19j5Za9+D4kRBEMvSMRckuqBTw6yEB1gW65HSaNkaTDiGiWsRDag2gaRdW3C
roYeW/Uic5uauew1+ggo8Wgt407RoF571S6efD6Z1FW36Cct6Ys3slPBK+QINS2M
6x/AeePH0qwshXtZmztV8v7QyVB9dEFZOaTPzAJ/FwNoblBNMIwaS5X1ggjtqulQ
JS91pmB2MA71DjJoafhewc23BCRJo1guobOgs9YCFgIX14jTzGK8rNN2i3L9RybA
23hgHsIIRcfHTDZQghx+t82KgCW4bHsGQgWVl7Evw95Hn2W3ys2vErndapMTH3on
VfWPFUcU5hRmbLd8DhauGWHKVVQaYIbeSGtKu2A2kwLf8KcxEvrwdS6uxNdi1vfY
cYLcZlq58BOLAKZHR8/eLFzEBKRQhXttyBeAfwlAsimtYgyQZWyowc3Xb7yy1I1v
H7hQw4Aw0lIxAjMVnZ6R42eNnXmAPKJYaU7Js0sMDSPNDrYMMf/KFHG5BcLRTMN6
s4AiuCzp5l7lWjXWMJg3ZmWPwEG1aJJ/LTmy7GUbqQ7A6wBMl3SHKG7BgdYKGzcZ
KCmuv/4LgcRqCgyBhy5yMGSXOFS2WE55za4ipdhRXW6sAUPRIT0Qo0k/7HemxMUT
JSWKgSGgaonyInBlKeda+KVsjIcV4mlM3bCyav45io1WUHp+Kr9vcQd8gYVyrxB/
6HSQl4Jg9ODx2PhxSGioxmLQwMRXO4DNPAz/ZBPmpUBQR4fWVjrF7EZ2uLBy9/Wh
usAI219F+bKV6Cf4Y0g0i6m9PIJfzPi+MR/ryDN4/ZK71CPt2iAc/kHeM1NFxlcj
hCLt2wBGgel9zM7n3wJZFiScgNpAupCOjphVdo4diFwO493pQmPTo4UtvUKtqZzX
hfJljA6PyhF9ArIY5zGafSpzY/a0TOq6CS4K+PfL/kUiWAN7MUitbq3KZ+6GgLnx
0mgmIZMHA9BCfiZ8WaO0FMucTTbLtEjHggsUZmRN58V3IsCc8B2UKIg8/tG84CuH
leaqB1dSHbs/52NATiZOIc4CPPpfMNpvVKP3zGKVx35yHjLNQNQeCZX0FiqvDWwL
2ecG3LPey+mdmN2xGH3L4/0Q89O1gRu2f6Q37GnSR4dP3V4DjAoUDV9XKpwytA85
7YqxcGS3av2DmU8g5w9U9NHFcEJwjMzAEf7WUkE/meZ9iZSUakzxLQMNLv15hRWC
X8bFY1itg7HAze7A/A9jvkFa2Cx3wOLpfcfTtxKLdZTusIO0iiaWEp6MeKVMcygf
Pq32n3rNF+bwtWy2Qm/z6SNVwbCGrCYNWgyDWMKgE6N61bAD91/XBOict29XoSvL
ZIZ+aqVLD0LydvjE8s1v5pyEPduiAq906TnjuxyT60gB0xB14BzyFUGo6AykcLWc
MPR+f4mz8qF94r8ruJJkrpjukuFmIaOa3/UvohXSBaDHThzh5qD53kLjqqKIAIWU
Ww86sd+VtH+d55JqpSXfCaDLDLOBjVCZ77uNUR1x1vrHeh8PLDDuBuMslc7QnkDI
nQH2/x2QI5TJ+Xduy1jG+38GO82MWCbUimMx/vGMpI9Bjnt/qPWj+UpAaWZIifuf
6cETwlCPI3j3AOeo+5TrHPH/diI3BY/dvhKlueQI2kW51Cpnc9sThnZvrB8IMuac
Im6te9cUG8tiepOVqESr55PCCAW/UvMNpWWpb7qBt7m+xhifbaskCKzZ46f6kj37
zWyQzq/vEJ+BcY7BIiMsioS2qm3uyfCURqKAWZDrB74jSa235QNrQMqD3em1EcNy
1T0cix+bWu2vmxRjoeiSJ1cdwwuc0TX6OgiU/qV5hiqhZj9KXml6jti7MTPR2Uxf
TFMlIJPrG6BYpToHKPiqoOx1XmF5KX8EEGIoVahhvIUS8fXaMz90rYYr31u/IjyI
L+cU5mhmlDetFVCbGv0CYPKW12uqWm8zg2SnCm9urbmWoRme0Ojad6FfKlEq0Tqe
8Z0h+sH+0iHimlLUqW3/L1y20WJKHVeyZajT55mkSb2mP9zjGLvskPNyhHJnqTPs
lDqVAcs2EA0VAxQwwr7maDDZYezRfTM20675YrPVvk8XBmxBd8oZ8+Xteyegl95q
3393NyDSdjsEXhCAPLt0wNrZYa4XhlTFLmzYjmpx5mFYja+Om5kGDcjScqusdGQu
0DBvQz2tFi3vFYXjNMH7YuDouij5JE4Z01rZO0/PhnLwYflpSouoYxR4ftu9HYc2
GcH6FiCcPoJu8Cl7eKYfoKwnZODl0XB/JibnpHmuronnFwiWJWUdrhIX4UcvdIly
3NNNbFlS8MJrSkUfz9WqZ/aXyXGIXWbp5p6Iyg0mhPWuLqMI/8D7f7ZPZ2Oo2tAq
nY8oqGQIJQ1/I+qJRMlYSDV91aAD3bxaSO6yHkX0X1BRhZdIxAsr6kD/ycs6s8Tg
Q1sIMtK/mKADZE72DoNINMPeid95jPtTPbZgdU2JAYDFMZu8WEyh2TZ32PBqM50/
U5TcNx6KIzEdl/1M7VKIoBkbTRHmSNBS+7ZOHXcbm7G0T7WE4bNxoi85noN4/99C
a1dCVxq6J/I8fHWjQjr+I+cvZ/N9c+D7BvyedS0jc4v8A0odmTghPFnsygUjgpT1
qzBIAMLQL9pDM0A0MFarsMCIMdZ6GzniHhqpq3QVxBc/h/b8kzdOpZ8KkTt3B38h
3Kb3Lz7cZa1roec69FM95CaId6/7FT0qLwtgV4kezXj8J6nLwLlovQUA1dH9KsHL
cKUdEtnEhzuS3m0+tMeXlxB7OKLQ4fd5zN/qc1M0uSLgYC8i0Nc3LG/DWsn0ql9P
JWM60vhwgzVZCL6WkIgWRLuJwwOBuippRiWjLuMke24Nu3a7uuAoA+ENypEuAWWb
EUXHh7kyTCTkLSKKehLu57te18KRw7RIhDvbDJEzbcWxomq7UQRjgPRktpB2aJiN
SF/CnkoRljEmjmYUIznnKo9vy9TdzjvVUJBl0kAscM4UcyXxkIMq5gE4JPmdy5d1
AhfjUzzEYEsAy9iPUmW+2aDjWOicvaDMy0NMti+TvI2Pd+pb1XQ+4vQCn9/REmDV
uDn8Pa+CqqMstxZWtLfMzwTgbdGNY26aNCi/ODrY5Opd7+p3sgZbKyoktyvp5tlg
n2SOp8nNpEvceXPX/QUw7NmmXN/giV9kCXoBBOLaLtHVYGHocweQZ9k6b2A4afp+
PS7idKeeTDIXYSuY1C5g2HFOEmHiNr6hDjGbxne3TYBCfjwq6ecjVtMAOKjqUJk1
MEuPfWp6sX05Gu+nNjaaEDQvEuAycyRkdPT3j98ofZ5SMOM7w1NsKQxytqwBs5Ye
Oom2qutghLo/yfVPBQiTwMl3NsIr+U7jn3jqdQo2sjynMUhcfc3iW/rbdzkJDS/h
NYzKeDyfe/OmMtJH2GgSHVeMdwxAkPGqkegcJZnc1LmrCJmHcLVezSpWpHDGQWSJ
aBhaGu0j7cgKq4h9itbQFTOV03251I5dDU+p1lyc9GcEtvQycl3FUyJLYQYVjBfm
YNZWgb786RN09K9mKS2ndnYRVi4X4FzjtgXmnSUvHZrUUm08g2e7tPSo4D4qDsIZ
q5LvCvtfmAWX5iimZKtf6paOSb5IwNE1m4bLMvaKFNSa+XmKaQwDLoSDovMjY7Ls
gsDLaeiUmOQjMRRwJRqAzjtRyEKF/WV2yYIlK8rx3DIr/ELnJkmoGKMvK0Y6DZDT
Nk/zTYc2qauIWofi7cQ8hKRIaBwVnlvvJQ8X+OlAciXigx3CyyLm3Ya+MrF9tiwM
A9cheWUYD/yZuKXX9OJK8wkY/Q5nOoKJ8Qj3XV3pSLGkmEov58zPX4XmYMJ9/6+d
nuDWuq9dBXttGaqfZzyaQvGfj7vGEdR3E+VQMb0ttwl3MTwSOmnsu7fTexpb0K0A
fjhimAek1lyDfFBNuCIUTsYxO7D8Jg/gy9Y83uy8Y7CrgzAaKTekS4Gt+B7zUdN6
ygINdSIkMR9Eqo7iNlWf4xnCPcsVMUqCL44GBroViX1Chzr0FP95IFyEgkaWDmwz
XhZSXVsePN63SxLW7l2gX4hCFnlvDo8sgkFpENh5EqgM+ABGFuuJkCPhswIiV3MK
esJLUq7R5Q4X/PjwiaWopXecNg6W1zboO40tLSAuTioKev1viO3bd5f0tpXZvL1u
BEN1xjD6/8ST2dgWWusphS3FZURPq9rmn97Fppkqw8ZwnnWdAQ9ya4tLyFHmLsIc
MqPEvdJODNm4FOPRTj0DRFSLJ6Mu/vYxM6XFtgEQLQwHP/f+98k/MjPb4okKp/gc
q+I1iVbNoVuOmBpV+ySSWvmrEY0LBKnKDMkLQSJajM31xEYry/QY5iQA3PkpXsVl
yVdgzaZGs/lfQ6cc3Uk0tOwBPkvuTxw17mxBQumOntHKM5WbayR0IOXXNjDj3gpp
egryjYeRUnflNLmc956B4quXS9uEiiQGq8Gye507gti+IY6yUz+qWgK74aKdoorE
cpLDo4hVzu8UZ3xm2uCX/RMhvssOk8Z/H95kWwrsoYPJ7Gx5cwYayCsqBOVFE76y
sY7M+EASG0mlW3ju7f8TLKMNw36NXJzAfKjTbmbxH4dMfRmV37IfnAPQ/2/U68L4
krViNQuU6v54DfQLu6EojS9aLWIWiL5HQoMq/LsoUy92CTguvk5PVdHM15wAMXZI
RE+i0EaU2PkoUDr8F4bP+EkGPHbZYxPjbuak6RAsoNFk7/AIxX4yxtxy9/qoSLrn
69Iyo3coGketNhr/o+LP+kYNfpJuOh1hV1gYBsf2045C5h5iU7QB8bLqZbK+M+vM
OZXqbkK2A6A9YTS8WstFbK2VlY7uWPkpF1y8dlo66CCc8GE1m1PH8OeKeEudLUS/
Bg0XJc6WObdxLsv4d2rvvynL+d2rowJb2yf2lRb+hufWrkPwEIoSRl3xACpRK8EC
0WVOTk4wHhDtkHOh6NCdJpF5HuQW3SjhhqcSUxClNt4QBBnb3yN8kPrdm3irQ93o
gV41tSbIiVWRzV3xrAEGgYUQCEh2pQsgHthTnizN9mstyOm9OJP0JcHXaiicaYIG
couwbdlTm3cn06e1JbmhE+83i6xYPhxzHe608JhskC/RlHuYS9ybfZeNBbS/7Vjd
ox8cNG/vEP8Db1SQe6blVeDINYpJ0sOsSOFD6ZbDAvbfgR8HAGMgT8cOfI6Q/aAB
atIHfApEzUq1Rg/4rQtsaUxIASpSgKvThjaGXlZTJh+wMDxbCihTn8mvGt4fSQx0
fgBanrtHaGQwWYEI5PdK9dOdt1viUAdsGRTczctiYFpWm3KfFPsQeVs/QXc5j3BF
2WYmo8J73pC/6UoMbtL8uwrEbr1IBaH+SQWVo73xmuWAWvWAh0eLH34W+15sn23A
eRi3FSJ/DYn2Mi0AEiv+fQ6tfqGoZabQpTuLsH2fP7vN+eYKKvQX1SsjzYNthXP5
26p4A1DqUA89MHx9SsP3wZJ7MYKoaLuYUeIx5isXs0PkxeKAIH0pxKoEF/aT6J3W
W1UXhYDveprS2xxmAp4+HMN7Rqj6Jlt8pNcCBsWVqA027V6n1404ZB4yreWHqAS8
YHapMfSNjnRCOEj7TXLTNKsEvtAEPwnLwMiOUGPHq0Yq4+Uo4I2pcPpTyouqipD3
8ehgAtEfjdnXFx1rvK1pT98Yvg+fvMxilx34iMOGYb5uI9qEaMVQZ+4zxEbReVR2
ZqLAp6sYt96g9wCDOCVPgRCLxpwrrU3oqhWrJ8giZTvl2rVxzM2J006JLaes7UHd
Ibpk6Z1LqYtIgvZWtMG+89lDQHebP7yBBqwV98n6lv9Q9QjdyAM1i/ywOAlrm+oy
pOhlYISUM7K8Sag9d4k3m7kc0C8O3tbFvI3+JDF7eh9w/RWhd2Tqs9fEqXY0zDzG
507keMZygXu8oIMVBH1+k3T6/oj1uHyLvbt7f49L7c//jERYZCbBqhNR6z8dHMNq
PIXhzmOlXRkKDgXXwR2BTWkdum9cveuoHvp565fWMgFnS8/KfPxDK9tZ1e8FkALA
O7oxOhu7xzeYoD0JZ1fd+XFZG2LXRg1INlJ+F2dcgRoC+xMtMx5xWFpsxUuPnzJf
dbnrzCqgYgv7C+5hAogC/y+JuFMKfwp7z3QczIpC+f2UjH4a3lZ5LxthfhmWXvke
11+SiJ0ewYjtcmGRPQd93Sd0+/evj2tASo9OY4f1Us8PBmU49EYvGJNZuF3Hfb9b
PQO6vZA2D6keNF3EWSUL7TZDKYOJPPTKZgQoLHLgimMLgSKeOw7VE22xbsQtEG6D
FLY4uc/P7WtwuzODEUY0Kevtj29hV8NiidxhJ4PTZyt+HQWXwIxjtdJkdJJw2NA/
c6L8z39p2vbxDgu+2RuqmXDtjycfoy+Ghu+44VDHzlQqDYSgvYjc0Ka3cRm5/YUL
DhqB7fX3Xx0Qaw2kwbhF3f5ZvoU8yIEg/CHqVk1xmxTFFyxml/Z/cmTwjzLBFuAl
iXrra1YIxolsh6vY16MlKsnOFipi5YmCmcMLHISmkANA3c8MJxVEME/KYajd6BY9
4eJc8Rh6GGQcTUawYfhLUY8Sc+b1S3CEJsvZTQ4jHaEuQcPvkgYC81UngypK5j+8
AQPKzBXR+BQGt9nUe0Lh6LWEUGq48xT+nFTCJCfHZ/VO+QKR/DVyih6IjwTzhlP3
`protect end_protected
