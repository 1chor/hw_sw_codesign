-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
lMMSDvUDi+d7RrKjZr52QLnVaalkq9y1knsLQWVQxBoVmJUGYPfRwIeJSI295wVa
n3eJMoNGjY4HAWUfLzigvBkH89Yyz/aLHMP9WRbv8pOFAOwuXXRWygzrcYCcUwP0
Q9zgLKw1hGKwWs0iZXbamfXlTiHaAu31oJTWENVrAw5h42GsQU3Hvw==
--pragma protect end_key_block
--pragma protect digest_block
Fa/3YPuhka5WSHHbf6hym4N6y4k=
--pragma protect end_digest_block
--pragma protect data_block
iMO6tSOkLQkIl803gp/1JIpaW0tV4T+RY6jmVtV1AVlpWGByWcw1iwyZrCwBYsZH
YlPk8N2WojBvJ9kjng3wcZrQHAufUlDdSTou/DnAK+AYfx+cxvpYyBQRsMIfSajb
zW4x2T20Qdbn7uRl/buO3m2xpnkroM2/ENzq9z5yCfV/IcMtyYWU0kzpytOoeOsE
Q6ZP5P0CUBStCzZWjuZQo5H4uTx2lqQcnK5bnDjOpqtnYhMOjbJZSxZqhYqJwOTp
hjMeje3PUJsudXGEr+1hj1EyCVikzz+1dg47zZnVY/W9h0FhNAImXnuKyYjLei6G
k5vNH23ggP3YcCaInfEZSGAbsod3q6wt7hlPXkbOYMkUBreeenh/0jLh/Od639u3
d7tH5PwSqm8EkWRIwvvCeiYXmPE/LRbeOV+YG2KNY3nahKiyEgi8ryaxZhTKAKWk
Xc2SNwBvRVhsJpKiJAt70iaRFI1rSOqdDjp+qoZGuNPRAsxEH/HhDsPSOvgRC0gj
b8Eu4ZZbiLsYLPdygkDSCuXj7KAlcYMkgQBetSzvFFPzSNW5Qndmq4kD1AP7h/gR
gD9slFl+xQKjlacv0s6E1n/uyGCT2jujnswZkkp8MDZhocBPEs+PT9wVfLFkKcjG
O/E/UmXUXwBgahQAJ/FXKyMqIjjYinSQEH28V/2TyXa6ALof1ueLgD9/OwKMEwqP
tuS4CBz1jvZ8dAXCh1HuXVuhOY527JCiyGQI3ms0LRgXlqZg24HydgjAd5/r16d/
Nldw61pHLcU3nGIR+aplz4N6BZ+IxOQke7EZ7CwA5t5j7BIjLY5Hw/87cIfjpgnV
dEsxYgvYXzp1EH4aQh2OXMMWpdnWeOTEWRqy4wArwcVJrPVuDFMhZQ3afEIrz5EQ
oYNIl62ZdVTVi5ihy0e3hfCdWKk0f2KvuMuPxTFZMk29xARq1MJrV7GwNHat5koQ
I2fh3okrn+MjMhJljSXZOZEUKvYv4BTl/Q3lZ2AcazGRSWL1uGlmqmN8uQYTTu8G
HF5vEQQDkLYIh6RpybFISbSifYLsKhCaTaq57Xq87i//eoiYaGJFO1wbSCPd5gEc
/ZGSIOYZ22I3wAoUTRzsltsQrUG/c4U6LOvTFe9+bfmwuaPQQbWlEKz0JMxhq9Bv
Zt/CTulUUtd0tfOnmIq0WokzZ4QBu4SEdIAtyEedQfUIhpoyMB7//mr05aILrAJU
cnLuTdFs7o2+hn6iB/xX2f1F3Hi48u7L/eOet94KioCcV5bsRXHX8glmhNbJSC4Y
YU1TFg2r8HWhXcOx74EyxUq5fJF7mDGOyOqVP0geBmk9vSYn+yWYhozmtHLFQ1Ya
NW+dyYHez+BZhs8ZhOP2Dz9/yLIjZu90d+i1Z9E7TAjaU2clhV5Rd3+XMdRzW7mF
iPHc2gJLDMShHJAjg5UrDuXHsrWZQ+s5cVNTMl5QKNEiSLSJWSbraq3weiHJAXnV
jtUMHZ5GP1sQ01L6X0KzGnRJVLajDNfB7JzkD1+fNNmxhN6iw3gf0BiXo/fA+DkY
H9go3oRbsFSigDbVTO0Csn5NVw1kW4y0s2Rigxqf/PrVYPCOn9buoERCRyIQY4zA
0kiOTM1UgOjFby8tNYAoQclysI8CeZVd+UsSBQAPy+Ynpht/4FONdE3Hg61xaKEL
WLIAEfABiV5FwK8qQ2f3P4I/oeVGM/zxtLI2yo12ioUfs0as70AG7Pn34wkt8lBS
4ownrfToawttvobZg6X0pzz+bZb12KwqW9KU+Wer34lEqqR2qlTQ60xCfr4tEaii
xLUytZnpTGAvLAFN3qNMHrSpCzbO5fwm8kTNRPYkqi7xvocmYsur5/PAIxd3mrqC
BvGq5c/UIHqhel4CXg3QvsLdcaWMzQs++99HLA8I05wUXzvHc/ji5l9kRbBS0ZJo
fvNucH7aFg7xL3qALXFA8Kx5wPrek1QuLFmxMi679iBMoUtLtVEc30DYBNsqL8lq
NSVEr8c74v/ReOzQxT+qWmyd0Wcv8DEwWEfyFnuk+EHdADBHHR8b/rT6PEu7t9Fa
1NwIYa91dQPub/pWVyVv3nFXkGIxzu7lKyDjcgcNy5x8rnBy8NQ9euRnFHjUwU1R
fU4KqvZZ2GPyaPy87NnRA81N5FLTZP8LUWlj2eVrG9QNJZyfqtWNzLkoAnHkEUqX
ky0u5ztD0rOj8AeBj3HqJmWZxLM3IrS/1EqCFHHrf5QEwDyWcozOIKdWwxfBqG1U
ghncsa/PtSOtp6sy5zrwG2OT5f8ryCmINsNPKMqOd9RkrOluAopgn2OxckPWVmi9
45qNfu7pKKvOy2LzdF8iXWSCI2MQ90wtdUfaz43SH4aJWrBvZuwVVOpV1+3gNJ6j
aNSCT7rI4RCWLDBIFq7/TDlup9C7RLIBZv7EFeaD+s3g1YQwgIRmVC/OzbJhFlVM
B1Pppt34dbWyazKqBcMT6uhVKEaEWdKOW4Q26kk6X1v8jyLqQ2blEd94uUT8qlZY
G9YDQsNdw9xW7s86NSxKmCFH1Nu5Ge4lqCJ3zpRfnViybsFU0FSJ2wNQgSObpqd5
H9+Tt66qzl+IuDfy8R3FWcrJiC14BQb+KEDc0NateQVtpOpK0EW9n95yx3iV9X0s
fQWR3v4N8/tUVjNIceESrubMDozZvZg8q5CAgJiDydXdXzoOPR+xdbP1fV4GsWbN
+R4kqpiRvVSZIu4NiURTSi/UR38J2OhBFF6TdHQV/5ft75jWlkW1k2C9rRBI/FJQ
cULFCA1oE+nk5p4gXDjBdBFHhcuzyYPNF3/At4jyb6hvyGbkpwgSPSVTr+5EhdIG
rapZCinAy3/Vs94lVn7+Ozq38TxAyL+2xPxdNyswwVti/noXeKIa2Gsw/aNuuxKS
9OVWVoggS+VvSy+mYVepPiKit5VlFdxobgCHFBUerTp2ut91MUJIMKUAootN9vT1
VSPRz4tg6ty1pDkKDCnSYZ/yrUVqcn5pVQQOmW7W1gxRiq3Jxu1NxQjPp2RQT68G
xEyHVarKpQHfDvmW9njJL1CX4XQY9QyGZcwBZ5x+sX4oJNOujDcTT7p2qmlg6XWu
DR3+LmUqY32x9KcZkqKkXgbInq5G+F7o9TrZ9yenzzlznZmaJzEEDVsXWeuerJhM
opzLRr/dhwfAZworqxge6Y61j8EfVMGvhav7EPhJVroegv1JbjlLZaiq2UL5+oYS
XifjH2FMZ19ODBqKGQh4oaTY7ibg0yT3j1W4wpX0sl9KhsLwxvXUjRf8hEMHjDZK
5s5Zfq3tE/gTpwPTTnSEVQmRplrve2xVoHIp2ualJqHDhiTu5f6qlenS9YSgtqd1
DkpPNRmAkuQ95AwCdvX8TxTnvv1nqsCoT7a8StnSupX7tTGkcFY30zmDXlqNKhka
qwm9zUKePf6nhtNpvoLoi+voc/yYwA6WL7Ys/A0GBraQHoy+WAccb94InEHRAgh8
UAPJLk91ZkKNi+FWDV0ugUdA41453L+tq+E428X1yxGJ9uLNqFWrsu+vSGpENPVv
yrYM/m8gWI8owrAdv4DYKKKDvrsxlrQ5ZCzHn9Pjk2vi2b3r3JDXcEB+IDxD6QbH
5jmDbDuT2nlY/EGTbmTuXjglEQ9YfmVUJGJKL3tH6Rni6JDUy/pj4vDfIf6VrtA7
5fkET2DhXPLddyDEpJePB6xzofWKz/6Ikt+h5BqkUvTrdPQIiM1XGEmb+zefy95Y
8rC8WN6JwZT0/LKPleA0ESx8CsfDSQ2DtlIo4PoJXmj/bfbufpH+tzd2sY9cilcW
uaM9+Mk7BlZnUtgsUijNxC/ZW4GWIdTW0i+C3NTiMFxUKO6Mmh9CKAWyLborjere
ILza0pYUerNPV7Xa3NN8L+XTvl/lFDH4WZmAcakISN9W3Y6xM20J6pZlypVUihaa
8PKzt+1Fun31Vn/AsnFtyOMvMWZ/8nbWYvOqUILH6V1wG8EwT4GxAhATR9LRbiv7
Fg3F+hm8MyV3pUb5oow0gmpOxy73hncR7ZRro1+mxZkq/9BpjG2qLJy2TfGiQitA
ucJNYnRWZHJElYaoJ2hW11Bp9wLkgl612lMZHDoVnkAZB9aRSFC4KKlfHQwjSKLc
+B1sy13c7qhG68r1WOdUZUfodp9k7YFyg3N/ecDStkXW8HFPRbegEL0mCY1nYa8y
x7yHyJycMVfIIJDsw6IbmreSDQo9wdAgadIwp3UZ4LYP6Kx9eXT1CCgZwc8yO7VM
3Ogq2jhyS113G2k94eWhissFAAVjnoLtbIYRSwcfj5QD7d96pUTLMRLBnOgyWHGm
ppQp9DbDLav0M3mxydFs7Ms3OCrj8c3nhngny6xWdHHKo1MW1RyTq7kCgmsWeE4K
okLx2WpfcohFrJ0LMqE1Zntg1pxKpCGmVr5Sov1cdStBkGNNNquo/WoX9ZK5nJax
zdX3IAl+kbJCM7+lu0HlhPtnGNOBajenzgJaOUHWoex0KZC7OzfiY3Xju5zXlD81
5U+7my6q/L3FZmSBoYJtxRDCTbEFVrZZdL5lSv0EfcDsH3LqT/Vso6Pf+lG4oMst
K4tMrAz9/Za3MuVjXPm9OLUW9EsrDjojKSQfUyrnBV4zE/pHKH24Ji5o7xBIHUdT
w5Di3uCZYn+yFoiRaqpn33wvdlMaCo06KsntD6ZwcZclXCdLdqjmwed7KoBs0htG
aqhRXC++HTlGOTs+yQ77ZviGZhEP7BpH1+CObgxThaW3qswqS4fn9euTmawSXjRt
wmHpdye65btlWhuJoTMe/s+pzfJ+U4mU+XiXn5YoRy2PYF8PdgL03noxjflkNuz7
ekrRMLjquIlafferHk7+N+k+OmYQP9V9Bi3DlUa01+kH7Gx/LT1WLnlN23bQmfkQ
G5MqqywpmAVfS9MpmfKCIQ0+iAph0/PGzzP8ClRcni8e2KqyPFItrLTgQlLbd3hp
iE554Yba/iFJtx7opvrACc7NE4g0uhL+Ro3NqFKBYd/PT+G1iNU1V4TgkBrfjj7w
piq/z0po66McR+47UNEacKb1J7WGhOiKDfuSfXGQC5FblFqK/uIJf4RJbIKI0/23
3c24xqbOA1Gc3Mxpro1FGCGUmctTYzvv0Gp9a0JVspi4qYKz5u0DSuv3e9j4RssS
/Jk9hXWeLrw6Ww2owku4i9OTVxcxbo/aq674LrYW5IsStwnoOP6N5ZczIpI4SioX
rW6y0pr0XiCZAUxyDdvwJZy3gToKQN7vF51sWPlbT1rBY9IGMbLPyepwN9mS9hLJ
sRl+h0NwJjCEUil9jLu1orDuBuo74/Kcwqo1K3/iqrvCNyoqLzemCYJzY9BHFHUq
0+aUWCPsp6z9JxtkHiwTIaRrOhhvdVbtR1hnO3U3bAIwCbAQfGmlUXHA/8BviUFq
ZwecFUkpwElZmcbesJsx9GGjsv0p8ZcA9jcDULcoY0GXnAWucDOeYTMbA/yXCNsV
K/Cdj1XywBVgUSaHXgdI9PVnWxDcbT0W4WHkzxqWsFZAiNyGibB6a2zRvnABQOyL
08WONzps7+tHTnPTGUiL6b+bdmwFoFpF+U69o/LXcCdSoWQXRBRyYipWkJ7aezsV
WBwS/pkaUPSf2HByWhKWHC3la+tiH3gPbq9d4N0r1Zhc3HUwviUOnWlL2ExdQ0At
KDJagkFv2uO+yXSu912VwgDKkx/MrsmfKoiziU08Iq4QAcJYBpBCjz5BvsI0CbKw
qAFDkgky0NuGxb20MmTDraquR/0n6+kQKfqgjnzNplUltgc8G7zp3ZD4BXgGAXEz
AdjuFi9hKQXKTsCBdSmn06L/IqDbTX9c4KNR/jAmVnA1uwztCfc12w2NyFtaAOx5
50+b+I5h8GVAuVNMkloslf67AC7ew20qY07uWK1fkhncdg5jeZqUG9EvSNYlXlMo
8jpKC2FOx2w9V5AkGc/N+1NwJv+WT9202hn/IafT/M3agdae5NbR0RfZMnCuIC1q
cSDQCBhUhwXf/J7KlmAcrqMpOofcLBn32/5A+G8yi/5Q092wqy2fKdfPQCHnywt3
j+/i8VparC7zswqRBMYgiz4DjQwEjyVTdaiKKFKp5U80JB159YGxsWBGbgzQ2THG
Zexw65eqh/TNUfc2UVZ69I/g3+/NWtfNlF+dhs4HlHhTeF/i3NjAMprsxKfbU6F2
VOrbRGdnmpwkwe9lQ6Nsoshp72WvZLZ3GeP7JRpYqVAMHwzgujxbRNBAS6O5+nOf
wkeqvlgeElGRUegYd+oRB2BHisx2qf71/BSoptPGW0qwvq0lwyhe5zBfHnpF5ige
LBySbkRzGdnuTIbdHYda9lRk38mg7e8ufW8pw5zZ4P/HIIOklInLcTooKhlm6/XH
Q1BmOx5Y6tL75w5GnYaF8kD5mtBvFbdTU4PrR0zM3N/wVgv3tS8Wkrt3v0sMVW+2
w7WW9zUsP3Mj4zOQYj91YZ8GXqEm5f4cXMtnV5aqNwuobY0MXNbfjNExp0GZRpxl
6Kn5FhDUsVrFkxuODQ1BlOGNmDIYn6wuY0jcT7nww373Gg5lfwUcVsRC1avefT1A
hxruON5IrE3f2HRd/soqKZocP5G+gpNzZAWRy0HSjfRKFiSDekDzXD7zrneInmC+
PKVsfLi1xB0cAXK7l8qRdeXPPpF+W5RLRaPGVpAom3F/WrHfseI1UbrawM8d9LAT
Jr9fASi4JJ8N6WyB9N8q12dq+PsSKZb0ls0x9f/DxHkcOAaGAUeZ9+LgwuHDdpIs
Vi5yaq/jDe/fhspnrS66zVfU+7s8nB8tZJ8dPDZSgDZmAux0t41DcahfZAhSsPuu
DkiS8ohxjqsAwGHNCANFsMMlLD+xQfUc3DY9wfBf5v1xoYm3No0CwJdHCutWs/7S
tsemnEH24jkzMLU5kPtJyHmRXaleU4KLM0ozjbD0Hg0HcmfXUHHzGbRa6tkMb8tR
MeYPdhrVLwcKoZP/hh+LwOX3GDomgQ1jRb9DgyaFXuGbfOQMtOFDehsFHKGmIG0X
0CcQ5jVIH+mv8GyY6ZjE/tnB9geiPsKsRz8md5QlzN/eENRCih8x22nEtvG6TOn3
r04KzBCvlQsYOny94SZJ9jUp8NE+XpPjNVVTG6dvcY386PnMXKjy/EB38Hj2//XE
zT2phcsiD3G2HYB+1NxHZssxIQ0++5c2TtQ3nY3HARXsLfS5iisY463Y32Hiy9MW
LGRfjycdcIep4tLHsTNzQMswbjk8N4z//o9+vbgQXs3Sdm+mvYi5On1AszodpBl2
OKwp1H3ytwPx6KsiM4AUq/9KajIvhAlxYedqRz82ugv7KbpXKDxNLF/GvcCtPITE
0YCicrUPm09yEh0nkBDOK7WHF8scsAjllCDzLrOAAc/tDLdIp6Ttgz95Yh0stiKd
JxcfvoyadYVDejMKi00VnHlAHJ5ICBmR3VxM6nqKtU1CFoqtPRUlcMwSXJsGMkF6
5RtgOeChBfbLPTk5shLzgMkHwODy4z8VFTUdf/+NUJVDGhQwYA8O5YNB1FU5N6Vt
qF6s4m51EHLOwygvxtqjCOJBB2JKFiOp3apgIh8ttklGXf/AvsR3DBNguLjpouB2
jS5zsEBSdUpaEbxMLhk0zE9Kyyyb8j047mficqYTDXx1LmwmO/MfLPlCzL6oJNgR
9mWHUkvQxJCRy2++lNmOrF3Trb/NSEeE1GxGNs6LVRN/k7b5XUp9qn+STEZzuiS2
4M/aAvK3dGKiriEIgQHdg6ItQTH02FrB413DoDyapdzxwA4gvG+eWLqpLMpkPcdj
Y+5fd3I8E0ck8/EzAMkeHpJ1V6qoZSMTGQLQbq1QTwbKzfviN8OVIUhB9in/4uLg
sK5BBQYFuoOjAeYmc8AfvVFNxVi3x5YFfliOTY+LOe1c4CZD8bQNXpNiGoT5yA/I
bn6cmQYvIgiaISIiAgPm4emQ/m+qxgtUmj7tv1lMN6yqnEKBCo55KVaXSYve8msj
zi6MOM6GO6C7+Y4eO7bTL9aDsf8bd5LEK+sUtSCHViw7mC0WpH7UWkYnXtpaFXfu
+HMewEk/S1BPC0rwPW7lwzeda1um6UfQnDgetr4KB5tHkC9eevkbeLY03z3sQ01V
XbKOiyhgz9+4YukaMxDXG6gn591yHcdLQdtX/kO1Dh+bKZ2mi+IOnwSpKtXLhNr3
uLvZyoeheNHB0NXjGq/V/uWiQ1DLUK2k9yYIBt0xl7Dpe8stFvuD2S4V0GQRtj4T
Jv3wc9/EPK4uVvedNn6BhsD6/vB1JoBwEnIiVO1pG8SQmwSNdZXZ4pnarsnROYoQ
ABmNRLSPUqhNMW/f3lU9dvtwCgBO+ph5aeO56r1eYDCPJFIM8SQIVs0ORFlXWWjQ
65vEb3WNdRJ5MmruKQjk8vnDksdct/B9S4NfMWGNPp9xjU9yV/8/fiWPzsKGShYD
vSGLndy1gm9qO3J3mqHc8/c6KB05M8UdbYSQ+3LwDARfI1q3TR2b1qenmQK37nqH
ENbScjRVThxmbgEJuYQ1+Y5MtK9te1XysS6ORIW/FjtO862622K+DSnzLzsLx+h4
zHz2w81VUDwjP0fvj4rf6/J2RubgKtG44KAuHIhPHdCPOHwhSVY9RbxR9602JzKx
mzJ3DQ7n6fKUz99UxXVn/2L+cPCGHNSXRmMni0ehqCwugxjLoNS+dfYOoC9Aj0RP
PVfFxhayLntpaiucuDtJqjnu93GPd+kYAPECOQEWzTjp2ETpwEvSFsaYMO1Z3P22
q2pP9pv9zmGaSVqI3sT9MA7Cd93So4KnMabQjHE4BRVwEKB5QoZOQm9uxv4Ogv21
ZfUr9ftYeS8KSM1YMW9H7D7UM8pR5Ohjt7ZrGtpJTrXXbLu04cwAMvS0DvBI8tjP
L1x6MhDAgzAAXD61rT0JIeJQqVoBpQZa2rwwc0NjfqjD1pnNQ1Xm+vp28CzTiZuz
7OJJvH0Cjs7GCFOmWi6KKk0P8ZzyN3Nv8NsiF79Rs3DQgeJ6VYdhFmTnz5TZErbb
7xSPUsnLoGMo3s30G13gmuXX6p0ylVLoz1jaOPf8FTAFl9c4oLvhkMnKOXsVlx5u
PC8e4Q2MisMas1gnvfD2aVkWFPGrERuuiSM9XzSm2q0SOvKYG1sMmYEiYM0fvoHL
stwN3TwE6aGjcuoP6Zi5CBEX7eVu0iyy5ayTsXqV1nj89laq4dNZ+Ac63DqQ2u4r
+yYZO0A/3sMp8vx4xRD3lDUu4rcVK7ibaD9LNFTWWwj2oQiuxtzVSqMU0jjAoV1F
67sKdnV+KPuF69fzfqRwDgxNH+kplSHkSyBSm/FiKI5sstTxX9QrEaQvPBnGW0U1
OHBP8IQTprABEmY+tRYgnHpciWLzk3deSowm9R3w/WN1JnWQp/mXg4TE0zRx/R/r
kYDGDmadhwwMBnbI4sM/LyUtcG0m/98quptbe2EL2fVUkPEKuxsv01uRemRiLTrn
WoKZTeaV3fEH6Mbw4KD/vHjz/jB04gydhLTi/3WJ0CnBrCef6lrBuFbOkhNgn/tY
r1FHwy4+Q+nuttJpXIdD9hFHYqz/ObsB8BaskxBaIHnifTWiC5twnPPT41aMwUl6
BY48iy4WMkH3aIGoocdJdwQJ0Oe0F3bZUeKHv9I6rfPNG1sIy3qmg0OmjLgsq5ws
NArhR7xLeNQRP21lHwG8WxyyLNVHG+UJzGQjkI/pLARN0DjGGkAAFd2JpBBtnfCT
zS0zmxnO0efrPPSRNnQI+WxhGAco9YiGHlA/OTwJtLbAkLFRh4uJxAPyDBcc7wy0
TlUeHkxkWRYPGIIgciHec+fSyxAyrmJxMBqwF6MO8jTYWM63I3HniT+b32zG736b
xzlZ9mFF2l7S+RYGymG0yh3X2/jsEN8NJpZfscPBuUgFh+cdBzW8XlQPr2Nx2WJl
i7akcc+rxlsBeBoAB8RiMDzKTlU2XyVIwqO80P869Mr4JtKHFjX/N3JVVmRw78yQ
qrL/M9X8O/KrY8LNzk62w0A4AZaXkcHnS1asOvxePEzmOij+HTWIstK4RtGbU9au
+mJ23Uj6scZ77QfJYj+cLztyOxPCER2oBVa5NLzU58fd0NxYY/YolI08qN37PrmL
Kda+qd4GaK+z7Mng0kj9RrnAquR8LufiaRGX7ug3RUH2G0x21oCDy5te14hODhvC
ZKuwQVJqOr7TrDr1aRdGApoqtkfRp4cGXTukGkwKI3xT3i8VJGFZRvEVsMHM9e54
n2Cv02VpBeNml9xqTSci+UMqQIwVqE4PiKbCvHvL5lXKylrX6D038xJQ1yjLlQxI
zIk9wP9yOKF4lzGNI9mTMxZ7+q7Cl+Kf82eZLQU1dg4GTKen6nC0JyX2/rn0AHS7
fab578QvP2DaEiDXJwBLoI+AsW6HzyihbXtzdClCdyDqn8XxT1fkeaus9Sl4kVCC
7tdb87AjF53pIunmKHt8RE5dpFTZVX+bOiurriswc1/xuvSmRPtTR1Na7lXHHZvH
cGbzJ4AvBwreYtwNUX2CVeUKjP9RPvMrVQHF0BY/vzrNjg93sWEpcK91HSZzr41J
eGzqfaUsA71mb1v6vpPDS4+6Cm+H7ACrL3np+f9D4wdiQHGbWEDyQ1sb7i+8c4aD
LuGPWoUVNo0WijZRaZLWTAOj6FGKRy6vLOeQ2p/3qMfHnmtnVQ4Bhls5F9SKyDax
E1q5H7vBYu3ygKt2NyqdAYh9e4QNvQy23nmAA6XjRBpy/c3gFTxVyfigO5jOTvGk
p0tZ5XJWafCjzCTp7rkgIvkP11oTJ2LC9ym+jr1MQ+A9EjROZxuXg/Ea/8vNWHJV
dMuVZe1ucQwu84GncYB6ezArYR82t/IWDqUkVUi/7ua5cM/qihgPDtdKoneDqon3
yWIVsgfaCh3pUABy0riWzOpt4hw2BJk+G/D7WgbywcoJi/AsJ0t4DpkITo7wXZhw
4kzLXyCUUe+dUNYcrs4gLAG7+RqPAUWTIbF0KZPetqeKcpXueLeoAzLaLSujvhFj
RzHRhxdxUwZZDaGZUrFYzgPs2UMGCUrtJeGa3fv1Th0XDNzmSsU+fkWkqirwBzHb
z5dRCCSPf0pG/lKM0Y8E0sh9Dkz9VYPlYPmbbssQA5zfxf4UqhAm7IxdkxD93I8Q
VxYwYhMRihKr7TL89Xi2yquvk/c42jkFI7vMQalyGv9z8O+hcLwH4QIXKZm/t3RC
yh9vE3ZZfv405i0OlgWxL3kgQkqbaGqaBsFrCIhEI1Av4BGnBaAOtW5UpqKOTRPQ
4OblJrD41hy3P95sqI2uYdgcr3utkqkqmfStjtrC9zoeklovGfhG3svRp98WYFq6
yF3IDYz4N3MmVnse3kbiWclGAVOn4Xqi0Dd2A0TvBWclYRsKQjj44jvsXL1pzQpV
qi5Ef4SKiRLMAPTym/n/zXDtG/N1DuwreHM85hRSCIL/3ssyRvsI3iP2GQy9EKzq
sc1cVwAr1QOc+zr0pI8oKdC/GVJoRzM5aWdNhrC3UjTnPpGmLUCejtfV0Guwbml+
uG0uFbu8zIVelINlqLBgTBrKutlAglQHJNtYHItrjvdr1/DhEaJNWZjvAbKP1HH0
HBkKQtI8WX6vkSyvo10JYJLdt3CO99y671+CDPY1TvVNpv87he8FpVX5dImD8fyh
lA6nRdl8JZH/iBnJADOi7JOzdRJFPXq//npErqGH05gSZ+QcNTXYMQh1L8sMYn5Z
1PluCZE3nn6g3oSPk16aCyJ1Bm7uuYILa926iB4bdLrFFOdNwthR+qFF6dOMfHJs
2LoV0ans7Fp28tdpv90AQPQF+xkjpux9dD5cT5hbSYc1Rf5R2ellk2dZmXgM2rCT
DsQ+1Czx5Nqh0tPUWJ8h9GwJ5lYyXbbDvdkIfWCR/44NQ7IDhnStUYsvXiX2r5LK
hYM/kJ6YYsOYYv/yD/GoJGbMzFh793M+S0dFYOHBJ4Jn27KUwTl2Z25CsHoeOVXU
w2OYb8Fy7TJJtdwnSvRT1NcD0u7BzzKn0anTgIqJMnmT++t8XEimWOaLiIg4C+qz
6tw7IU4PF+z8Re7BQT+Kx3XGhFy5+V4ixnCU3O2KNLqoV7wp8U7sQ14H0m0W5RO3
f2l66RxXHl8NrMx20mbBKb79J5El3qkRg1juaEYO1J7cOxsmDTvGNYC9ZI/o2iVn
4UKCh6w0TkFN4XG0AQ90KRcwRilwU2ZiGRuYV7yuBV9n1emmMNShzl5aA0unqy9m
nIEYD9ISkgUEIV75EAm2Ww4+K0G4H7HnTjnTM4BRaT0BNQUaowNNnFZW19v8Goo+
C28zAUqxFSr8yPIMoRMMvTJ5U2Cf+VTbuSw+bIQxcH0bNWt2Q/iAorc8a7PEolfg
H1KitXkUFe3Zjr5BYbdg/0D1/aGchai3qB9L39RVTdeZhUKqOXASJ4yRPZyv5gBM
BWJHMeqtXhhLT5N0VUTBgRxCBZGRuCHIanAPDs8bvG8fxQSjjJ5n6X3ICZ22+A3i
8kynz19sCe4kIpNZ+zfW8W/bn43aIX5azqEOMM6iK+rLh9nYMTa6h794gfNZgzgU
Glrq/L8XLQq4YnDi+ZZvxs2dLh+UC2MVPXAZuZ2IJlEJzGCWXZS5uRQXpJ4NLBeu
LXlUzFksPJ9chyGDfZJqBtFbYkv1OmfuDAbfDaRiBDn3qOyH0Q18KN9ekWiFzGmc
nDiTiIMiO3JRgpL/3xDTYqrIDEvC/W+cp96EMwZTy8mupqiViiH7j3DbPbHosgQ9
iTdSWbdKPS4nlSqmymL5qZ8V3c5fcYpciqrEJeNKmcuzCyeiAJamuZ6Ld9WSPbuf
lNs3FGaiPRcLYQWWFUyqZN8k9MRy33YiTx/4EYXsS/1WZ3kj20cJc9XPSVFWQHsF
0l1iJwDAErE3mvrsOfU2+P4+s5lvNjWTWXwHoOTJSiZTOhpQIup8ARKbvNc6h0wd
nesoZLLqPhYkjLrvx8Y78LzHze2W7B7A0F/1UB1yZAQkUcoRphX739xIEjUE96jW
FoH6HwgvsgEPIyyE60oTtM2OZFB7VmIYiQ9NAKV8+9FP4eswS0LxLBT2Ljxeb8i2
nmRFl2yQXmKbOG+5z2S+4Ak7DpYvIGJgxr3LtMdH7cievPbsO3k0SO538FFiwS5e
qJVwFYEVJdIoRjtehg0WElV1i8VvfvrM/TIe7TqksFs+WUvq/uxJUAvOkzLWhjMA
aPqf2isa7/a2I81AXlw9Asob1zNIbbVCBuuafxdIxIykKdydtZa2fN87BYGFHtWK
MGEJx+cOwGCr+iXh8Bqw4IOBe2AxV6IE0E3ezw6rC+f0+8N5rKn3aoRV3G4mRMlZ
YjPR90P7Jb33LtQkpRIC4mD9j1AMx6HfRjlGNg47veAMcMLRt7B4iThB43tu0vdJ
HudSPB34U2qZSsCs9fOR+sWUALzVF9ZxYfsouk/k00gpYaBzDC2YnD88JGk1mHiI

--pragma protect end_data_block
--pragma protect digest_block
pe5icxVXpHyCmye1H4u1zS5EgWY=
--pragma protect end_digest_block
--pragma protect end_protected
