-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SW/IfZS9XqLb0EVHzjqtba10f4CfcvH7sVZgrqXdo5OdoXexe3QrnQV1NC8cevDFc8qaCIEy9aOB
vyQOlCgaqEgN2BzQcWSyv+kAbHUiX11oxKwt8wHh0fhVEQCXzmWlOOuVK665KrBecQFgz/CfBSos
k24qgUyGGcDz2iZ9TfdEdzwA1CDqJSTFP4BHRGF3SnwHpv44WUi0Q6WfWMQ86BhOmY9KM5n+/IZb
IhTGWkBwQ/gNffEq/1UWGI8WVlLnxxLOVe/gKIze2E+gyv7VgdWszxxL2vAC9CyiS+OcAnSQ6lzf
tSPB6kp/66TB8wIBLUWFNON3kKEpJYgs15cEKA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7344)
`protect data_block
N+O6NrmVr6cD/ZrqFUpNoMC/uTlevq43UVnBnT5KT5UoDaM0CfzZ8ZJpXd0muHErhhu1JUh9Ik2h
8Be34abNSOpVt012Q/eVph/AkTuJbqnwfkycK+/VppSALhX9tmXii219LWRt7O9KQO6uvW1ntUag
Z5HLLLKd3NqkE68mXLahNLLLCLh5xr376Zn0qk2zmV/Gts7VQSpm0UasXMSK4Ns4mf2VZU0T3qn9
pvG2vex1Gj+L1htUOdSdSrCZXASsTcZxotZdT294Ja8u2CuKHJtLwPaMVYgAJb171mugI51cf7zs
4fJpOYeqKDKuMGrs1yUzR0kn7i1G20MK/Sc9GjjRN6L6VDFHUOlMPepcAWNTBxyIjKmVH0nXhpnx
SEYIu2q4i1ol3yjLKru1t3cZoNn6HVAc35eEB0UJOfl26SDcGESS59uz8962Wr9EC422pWHtFY35
aLsowEdtSvz0UbOf1XRndiS6LCJSg2egN5jo2DpkdV5SlkdqVI81N0gq83uRhJy2ea4qydFZ+IVU
nrTZX8SAra8kFuBfwIcG0TvwjbrUH579vlMbLpMLYa50MiOXA45L0EF2bhH7ao9hy5cpKxT3VHf8
fNXQoyBhTK7yL8QXvXRJAT5KY+k1udlBBZe/IAJrclP6tdK59DCJQtEvO3i0Gy3V0ukD3MdQYX6X
JZLL0A6DEjmqxNcPuLgf4fb7P8MOJDPRFJVI5E86d7RTlFFmx4iK/SH80tVjPp6EHLgiBwfRJrkw
aacZ1aFMWP+1EUJOQxSuHowsK2qnKqRl5v+3rKtICQUdTpj9+v1yMpUdJIK/1TNBFmWnzejy0Gz1
c46ima1Biiomu93u2IHtmnSa6A8z2KGQibtkkIrmjUUjGOoMfukfnF5tjPuV/sUutWYI0Qho9Itr
wKvFIz+eJb9fx8Mh91x7xdj4ZI4t4vVeLpQqRB4w5GbaKc6yek+7l9nHOmzakumpa1JC/wjuQk2p
v9YIx/bU7D6Y2OytR4g1Ss+3f+V+Cl0CfpIxmPwQFnjUcSSIO8lMjL8OfcEUtTVAGRvHszn0DV6e
ymm9Swq8UMkPKBgB96VFMsgnye+50X5hIwF84MSvKFRpRcnILTjaUhvk2nh3OFavnqSPhGEW1ibY
5VGkH4pnK6lpWg7w/Q78gk/uo1i95uhsisfXUrg5kkhH0ZvtMe5X8GD9mUVyatq2mECZdJV1gx2f
VsDzHFUeAT+2TddLxbmXRaZcG+aycFaGK2Cwj6HaZLUFRoQVABQyPQLwc1MNHBYduHwL2s4AL3wu
EnSQdZRCAEcDAI6ckUqOH/1wWesJ2B3effoj+i+42eUxHQenOB2IjZ9dkIA6iI3DSE7nan3zN5TX
skAZ3ceqmLtH1YnUf1v/FR/2FK+SG90JWZLlgskqDP5OdM/at/gT3M8ndfVHznBMZWHAyaSduasY
IEMbzjQe8FTBClbNVWuD0qZvz2VVTEvlMS5Gnksfe0YOefciurZtVrnCGB9e3EaSLfQ2edItbl7+
rXSIE2G+oD6/ABEKGxs1Wv2WHDsXlAQ5viUGbGYIrIrj/He5y9tNL2ibhJ4PIRC5NbHqeIDC0vZ5
3dtm6CJ5eJUtwG6hr6gxQ1kxJZDJpJQwM1HSahN8vy1VdKCdj8a5WeFMKmLkUFdcGPCnESo4FQtn
gjwGI+rpnWTktZeDUGyCKopTeIqTeJemXqQJbmOU6sQsaZPLbNi+CuLtNx8lWj1a2nnlmMWJl0Rk
FOEH7+wiyv6xmg+3EYLR3t8bkzUfOLQGfrp2I4K65bTlNiIzYXLzsZzbmP16/5DZWB6CkhcXzdzC
zMuNEtBZaYRhuvFIGywrDdIrw4BLTaWwf9CL+Aza96QhUrGHhrHdOuwSoMwDzUFqeYj7DpnRWuqn
F+LSqdoz2pl7Gcc2dhIiNIZn83QRAgb1JRzoObnIGVzHbXmgb6hAE6w1t7NDNINTyL7dWhBKKC94
AQQG4aIOydyCmfbNrYhdzygieOAka9UZx/VMGNozi21PaplPSRQgrGxAL+JFGbXVSRVp07Yt2cNb
k7YH+jOha4FqQ+AwxnkCI8GJvCqnBNrZ7UoPk4fNkm0HT9XdYjZOJHem2UazbO3lLz1E/gaZ737I
bJzkdA6uaZjjYAdFISOnlQlwMngh3/HgoqmLICSGQaYCLhx/IHtx92GbymMpymdQyGyxV4rJWxjJ
Ra71MEp3vahbgn4co3DdsY5lbEdKx6coAky93evie3quZq1UrU+GVP8Lhl2w5cXkh9WUBy7nxNWf
LIB3YuqSgyaRJgqM1StfBc3nLf38t113Tiw5bDD9a84GV3pCns7NRXFfY/lCBYnfVplaAYQl3PiG
FU5Wo5bGZprq2ZliNi4fol/7vJtPs0Wid2OSfX++U0Ov7IEFOcHCfwoGT2pXmpToNJhEkgeRQZYR
9WC4UJjcdjxuOe7CXqlYd840x4SiJ7WrceZIRljbytkgbNcfkcc2sN6ofq1YC6TXXkAhB1/JizBR
QrPrSnexONPGVXkGpwpiqlzrsFrOP0CV3Njunyv14r1g4eSqsiylllBJzN+tstbwwO893S896bVK
is9OdaNKudAKPuOdyHdIbWAsFdoTnoRIp/BccHPppFoGFfg/LLFqvJ8/WL8eppNQ9JS1VyAL82Y5
oRfriZcs4iWcIRb6g3Vv0emCy4y//6gAUqchtTNR84Vi+jiGCKlYXYS4sKMyf0wl/RquJeO8JDAi
qDctdqi2l4DMKWPoLQ3MpTIp8GoQUdnviRUVMRFc/BIz/jL3PhiGYthV4pZWlT8l/bSOUeBc0Aim
AHI65GllrVeio+mN8U803272KP3idtfBJIdvYaC5Ljqt74SovP+re3Xs6gtGAx1BtjzjyGzvB3BP
UDLdGt3mnnUHZKWgujztKb3hpVirCM2vr9VChfMT0n3Dc/LYQ+o3LMQ5hCrCvTYxQkpP+FySWl9x
Rc4KX8CtjU6pZsrgp76dKuPn+LloQ6RBAOsBpY3ilgWTeuJVH4zRZZFSGaQmLJaqDEV67MCnQlWr
54B4QyKVLpjqtT14X3A9936B7zJ8IwpTiRGCpHQWZMPRtC0clWumF9yck0i/pBjq8mbnjb/kEE6h
62gz2KrNcqrNmPi8rrvh3n0gbMS54dFT6FKQSzt90H97rwG9SrU4zC3nRzpDM7L1sn8oyPl4pFUI
X1UToLju3X1xuRMqhaLPC6CrckbengF+nFpCwxrcksX/bV3BfmgRkMWGN/8ZIVy484xGdBDoXDz8
mAtmOlpQIgxiEA0X0MxQhaMbBEtc/9aXQ1n5nvubDSzYa4tIkyGjWw4M42kAuaTNMyt5bGL3yZvB
Mw1pxCa8bdEkqaaUAsYvsEM7XWqtA47EMqzbUYRYG8Nf4fAGZPG+iLGsNjpex1zv+DLBCGtRwy1M
knzkepJ5DnATjhwHHqYE57Vy6bIhE6wxNpYnD/KIiWQvBfZD3318EbxrMqVgJ6sR3fUYyot/3k1a
AsCtBexNWPzArktzIy5phcRdXL1rP6sx3nifIA39cUZ+G2FL2EgbGw3PGZHWpWl4GcJzRExp4WqE
RbKd1HgntEoLl2UHYgI3DPA9k4TT8JOidrLfyJQY+y1YSJFPGbtvPRuFcx2bx6U+TEb0tDpXr/Vf
sK5T9mvbjRGgOZIAzlGTiLyp52TOO7Kkt1Fy6Mly0Dfjt7WUaBkYgzOb168SWmqmi5kWXbB204ht
Jq4siyZ9oGMybXErKrYL9I/goZF/pW3A2dsVmo8tQUsbgEcerigXJ/eozkufahv8bAhU0XVA0CPQ
ZUX+JsdcY5j2W/dQFbCyOr0XRN9XR579YZpcc5dNPBcAISRq1wBlyP/XFrnFsh83gs1LzHi66BUx
HmmVBHgXJ/4MnPK6B7WZsvlPTrMVAnLnPFAh0w4bRl423S71uNtxR6sdpkdxKUozshOy2oSHa3m0
V8A1ZFz2VbAI8veVtj6Tuu1WktbCCebyS3tnkpOZCNVvJyjkCaPsmOIbT5beRP43OBBiEiSTJ48H
ME+8jpNYBskr4EJtS6aPYpgtfGWGazyRsWXIWMLxtyVVG9ulLyWCE4YwAglmZtjjz5w9283dasQA
sda5tOeWtp1vlVByH9O92ZD4VVNGlIRK/xLFSG+R0lQftW1TLza0GV38C9N/ZN+TaMIGE9aN0PTa
BxrCJIwj2TlqFuckwNMcNH8F4BQzdWF81wikCKaJfssJSc3l6VM6pe/8L/kaEv1tIvECUjeA1Z51
Tv7qtz0isTDECK/QxRnVQs0jA49Xg/R9mE5UGxxJqY57jHzHqzQT26QCaP7gWpd84+OitOh5MVD6
+nsv9xb+rgNobkXpw+ZbapXJcopIXM4Sxn8cqRlrONbx/YnrcdA77XOjhRnZGOCjyI8flSRLYohJ
g6GVqFn68lgwyxrXbldmbTRIuT9QNGmvxZkQvmR/6fdjk7I90Uw2la2cKac7U2i+i92pkZsuRjRh
xtlAiosMHU+bdulmUZ2bMIv+NxsxYr4PEioGsxnkvPCBt95q+ZZPFS8agsbJh8AjSvSkOFqsNod2
kljs0B8fD3v11G0NeQb2Olqj3kw+phmENO80KXE5ybtr3WVUzJ0uBXFTSxMXkmmrTqDVsDhFEirH
RIBX1x7J/CEKx77NB9dJiaEjBATWERLpudqjS9UTQtmOTF0/1yRS+kNzg6bYhpJlciT5QqoZFrSw
7mYx8R+DAo5r7biiR0rXJdNXeyXqBl6GZxyUf2UVnZjyD2FSIS87zHFBuGR6etLmnLA9GXoaT2ED
n/U+ldLRUqXV3WGg4xn9v5XeITdgQT/cNSHEjK7AnPz9hVP9AcaBN6KywXx8iU2wAtnKaPFpIyfI
K3LlM/TcOVmuhc5lLgkMbaCxTBnq99qKCWX/69xSpSBfolMn9NL9cNm7K+V/m1hMR+fEoN3gWilj
gkg1zo/kg4fcjrvDpgfXzSw/KO3kpe+/fQkA0/mPz7ls3vCsjx5z4Uw1Gi96F4kUlbY5UdhYUq0y
youMM6Feh9cfXk3Ksw6hph7ekKY82AK/Rt4w5gE2kxBQGfuBTr2DCTWrMlxqZr1Avlc9cXtNGkFe
JrPTaBOh2GodJKv/1RygiDaJrgKrLe6RFv1UZLi3hBVjaWkQV4JJGIuUJU1c69RU5dCtJGBvpABc
aJIQFKO4T/ey7peyenokQT8MF9SUHq8UO8KZUYzOGfvqmgoemoWO2oBE+jqlQgOOLTqwzmkrU1TE
mu2rqkua+qCPfNPIXxGZG9FkFUuTrWdtyh+JIW2ZLvQnJZPxOMeRf6lkl3sKl5Bt6YOVqZW3pfs+
I3iR6ipLb+tqFdHBTqDPFf1RFUVc25lxSTkhs6SUuhp971EHEOLVoXvmjSpFn1O4znnuTP7fwMwA
Yb3y64CrpCMQ9AlHhir8ZuFwN9JzsNvbRWLi+a1m33d6+1L8yabyr6Z3Fi9IbNfrpKoK2DRW6B/7
5TYKjpmkFhXCLO3bwYrZhPL5A1HIQ7JXJ7Je7+y33dK8tQP79h/N4mfjg7J8PKNkP58KzUdwT2D8
MO/Lo7aTrvgQ9eSk7dpGbQOdZVCL6Zp8W0uyFsMtKpUZ7eDPsKMH+PP6m6bK6ck5Qt/HPZRnYcW9
US0Bm43KH9OpQQ69jeXCHNwGVTlSGTh3LtPYLioOW8pzSYCg9XWEpb8YpaHpoigLGf+O1mDuf5CK
n59/qLbleqvvXZ1rvoVAFris1v+4xGgLc8rXP3bxhjX49DB9tleLHXoRLCVvkdeBIbTLZ/D59YYk
INn5qfaOG6g6RCo9t7yAlxfvuMT0NH6O1Kwbsg75ESBrJJH0oIxuIuZMf8vlc+hkNxTJ2kLykXUu
TsNZnb0v3vt9z4WuXFNmpFgTOH4EO3T1+9o3MPflRSdMGzoKhlak/CyHTEoZqBK0lKEo5CNT6JJV
F9ZtIha3YRGCJW3wbF3bcn0VILXYRiPKrIz7wSvQSTKouQYcM/dBL5J1K6K4Usx7Fc02TwmBfEmu
oSSbNo2oczlDp3ViF8n8SEi1ORluxcBIzE0w4jpplCpf05k5Dpo2D0BaVjqTzv0vnwDbq74oBUSo
wwoBvmZ49DqWN1L3Jia5HXc3eZGtmZoY7ghsFpbfE1qLuCTAm6SwVlDuN1Q5CW2wxgLuFTiYqohN
Ys5OVMhgnNwCnZk++sAKloIbE67JOFJMwpIoF/tUqjeNBS1KBwdT5Ns2D3ny+sfLghz9JG44Ovrm
yOj1AIOKrWPbII1WsReXb5ZR+zdG8p0ULjAtbzZ85InYQI4LbJRmkmKJRcDhodb7G73H5X7/+SSo
r6xsyAa0/W1jim7BjcaomGspYzPpGORa2uFMlPsCvGwiu0SS0yjG8MPw3jgtorgFi0hyE2NSuoon
0ViqjbLzIKLG6Q/Kem3QWDfvNMJ6bk3LBD2zBAHffdD+AhXjAn7MnuQW3bestbMyxjpq0L3GVFYi
7aZkH8jPq1iYzTe1JvvEzYgg6OA3lpilfDB3SkJzBhvDcotcotleVhBWesrRUe/QGAMDoQqYuqHp
UeFOznxuLDBspmsPRE5fKqjSXxo0A6Lu9gFHazvKPW5GQWwPS4Lo+3JWkzCgKPwXIfFfHX3EVT6Z
9pHKw1wWjE0pZO7/BcWR6d+t7nKYzTiDSPN4y6YVbWJjRJHcgR5hNxB7uoUdXuy4ggQaFO8ctOiy
LajChCRym9wuTPXzh1i360D66noludzhJQ2arG8x2L28Vt8MGoqStUdkW/WuVHIDCCdyyTrpqq9n
O2lYrSifdktvGJeBe8eFiLByH3Hv3VBi1tukooHedAKdvhzm6z+Uykg30wZ6RcAd09+K5hcb0hCH
M+L5G1AMO1TNl3RWtyMxvewOtwAdbFbgv//pHxF5RLBIDxTg9dxXiLpo1TZlgrNJcFQO/Ha+lXTi
sFRIsPyadI7CYsQwnN961aQu3Uair4DEfYvIlnpM8fl10cqalWB/ka2zE1l41Sjmsn2bmHGcqfQX
RgOQ7LRuRNfGJmX81ufc7WzxnMrZwAXqvfg4i76p8Ane+GARXPvXH8kDAwVfHfghmXduh9SsZWqc
67CsWNk/OcqAKXZ2d/fmfmz6j0afEpokgdRh9mVaHlg3lw0TNtspzBJGqotd+Olelyakeu+PsFDH
2q1zIhBpKbDkqEDOMd0DMTtiGXhHMAKsSccX2B3eegliMEEcfddX8DX6Rik93QoF3R0+0hbL6YTH
B+FRC9qM9sm+ZOUKcb7Jjp7licH03VZqpiScWdRbrRFmqwt2/urdXlzCnrBE45TUTv/66rfhwTs/
CbjCy/fSwl6rr/dAgjOzu3c3an4N6E4bRi5osEShfoHnKTHpRJshqtjGOEoMkzxW5Xpyq+egkg9c
QPWb8xuT7RYgBdReBl+MYmLrWvQBPewkxnGtzGC+fV+HArBqphSLU40aJ6AhCHpmAf60wdPKlnwl
yJfkXcknDN2hHjIgaVMrnWR+zz1dlSH1vky79OinmfrKmhrJXpIM5d4U+Hs7PVP7bSJi43it2uNX
71zrKGEYI/TfwmLNWU47gSd+h3fD45DuIFlh/egMon2UHaGGRrmlG/HxJ0mAznrSaAu6YIPnD610
FKGHtbrGFfwz8iz9yH9bb/EjPd0X1vKZl8Nyx+btiT65gT73hDKJ/YuG4PdN1YrIgnNoQ3bhIGKy
Wdjvsg86hEODK9sfqtC3MM75oONsDVVFZNWEodF7HNJqcy7SjfctYYUiPDQ0scIdtGcpuX/pi1RL
qGOdlbmNyeyVU5ETgSEinGjCNgoN3evqIvlCYE54iHv6hkNwOSEdWsV4YWf0lrLZYtf7bYNKzcib
0S1ad7R3kpw2AR554BfW4VAK7HVhx2Ukzkr29N9oxKsHdfnmT/LMP2dhpE2awAke/9HrNQDfS31S
A/kh3e+Zf4S4dIBWHO9H3QTAYEChwV7eEdJmRPcexjUpWypS/klziTmal2iOQDlvz+Sm0xVp9C7d
TIrM2INPVaYm2quirEL8uiAyPgPDL0NW5Y2piMCfoUG3OnuYc6DaHpW6xz7UnvDyZPGNtDDpdSAn
VgFp0pi8cyEQ+7pdIkyvuM1AwYgOptwsjoF5zEoR5hXFZaAiNzICMkiOoyyrYCFiZ9Dvp2FOWANW
nW6nlJw2KmXS41sgl+sCZFI4q5Dv4RvL70xe/XtZGtByhLJKFhYXQJ2JOMdYLdracfeSDsfRGnRA
q1g6P3QcBn2VSaJJD/ff+N+rJTP0JIK9NIzLjIS1Hx7NnNKGvq2wyLSK62iY5sU8CZItSTEhPdqb
D2hw2SZC/dhDmWPkKa5kqLoXNevZNZSpQVFRTqWGM+4dqb4qqDisDC4HcC3RiNRSrYpyyba+l9ig
4AmZ9G8SEXOr9aZBZMcU5z5F0zbwcWHr0PmArpNwz/OwpUogktv9DieCzStpMHfhAuGY0DyClJXk
JAKtLW29/7lf28XyUrwXR/AnfxqQBN9nC+tXaPYCzf1ycfL/E1GdILXYR7Mg75hLjFedjlzI/5a/
rOuNsPTJ2rAFJaqLbueEi0G7/mAS93X7itCmHEK7KlBdK770rKyhI8LAGw5U3Wiv3eGNaUNvTYmP
kYErn6/AvLnJ/f4p1ARcLXG0ZDwIIOWol+X1JZlT2fZFZ7QSGVjOSJ1tzR6VnpK9ydZIvMK9DThf
YBUuCq2SKOciRoeh/eI6DsaRVUSm9tO9VfrYiZ3OHStwfRemtVENON+t+dni81YBVdr51cZiqnE/
vyeN22wTCdzat9H6Tt5jTVTQ5hu4WhyDENOdViEfgs8v6GNw3UttasFVAXRJODe1Sr7c4Gwi9H6a
QqvOo4vuxHfdOvmBfIXtz860I72PAIwPlfFYUk8c1df7p493JTMVgPx8WAyatN8XlRsVBhP4se0s
Y9oqFAtIOTUYAYvmGXLrzxv/8/5rEUY+/HParI5k2RoL2+4f/pENviLHa9Fv/WSBkT5i0wW1vAbo
IbcAnw6N690WKjopzUSYBdTT87dZiHjw3SVZrQtCqM3zkZFrTGkUNTOa0Ik+/fLUiby3SrG3YDNr
Gu1ScHIujPZ+57wh6YSmyWpOvjO6quh83MrEz7QxXS8bLw7ov/TfzNUC6DJU/iREuXHe8LdHvAGp
taUMyP3HFO0wgvlMpnGLQQ3RTDmp+TaUiCv7Yju7n0RBlV0Tv++VPoxhrlRVJukmvReDhEWevQ22
wzRytKmSOfNWLBcPFNncA/kxptBlU7Rln+h3kweffX4keJgR8frFKmkSZvSoRDYTINJ7BCu5gGlo
3iXhHJIz5hRaPVW6cv/V9RchrpxjFON87H/3zt2XlQXHzdiQmkbhzDCjKpxWulpsqYQ8UscqDGRk
8uFfJyCj+OfChXmY24WX9Y0YkdMQVDElHexrzGNhHNM7dmHRYM8/o6a9j/tun/l5F2Xj+o5NSqZ/
lNtzUjCJjhR+JT2dG+TlODDE/rmYZ4HeRbz7YZKW40QCnXJSQhkJHi1jktsYAFnImCId0TK+AWxT
pfY0DRq5/ndLY1rlOEhQrcItsVj3CCIOiabp1QT6eGeTNec5OF/Iyb2Hpv/jiaZvLV6UtAPnNRee
SK0CElohnqyR4RSzGacTBKimgI3x+08V4g39R0B2D0946Nrdz3kUChXGLe8XvtEgHoU3M4pC+/ru
1e3uNs6v9nNfuUwU3sQtHZ8kdGuce3EvC3rbny6pkkbptuSSMb3iz7BHbwX+3SA26zYUp3X43DjM
gNPFymcuYpuWBRH2Vm/+KckmZ70XiEoWeCHHG7RSBuct5r6GvCfTlDlqYG2zCNYe
`protect end_protected
