-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bVGYkdLaVCyHHWuUxjr2ovMLXVXU2bC7f0x0QXhKrOM5tyWEWKzFCe3Kiuf4CIzZjbWOexV+KxkJ
OpyS2PIFoADevenUKP40PMQe5cFFXzKqGhGLRYJteH64tWYEg1p+izJfDJGvFiprptuepKVnJ6Aq
e3aRx3EyP22/ZiwuybAZwbGVfQqU+lxw4C9Je7Wpq2tVviXFxbqYHwVhyrSYNIE/6qU865iSKdAj
htM3DVtGQWhjA8x6zo4NsPFpitCY8szMhzRFnkHo2oAA0EsUZLbBel0kUdoiINGySME76FSVNJkY
5r9lVTW5rEXJ4p9zQt/RFPCS8mazsnAJbtzA3g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6624)
`protect data_block
vE2/kWCoBggcBWEEh5Oho85ZlvO0GcFszMw14d9+5tlX85q1FH7r9wK1yz6O60MFna58kq+YZG3i
ds8VdXXo4s9y9lO8v93yKTqumGY33H25jtPCB1SVSNHDv2TquB/fG41PQLnXjytGD6jrUDiJVZIC
FO9F7jfnLFpoOvboiNxR9aNruKsfiw/y4WzE2y0TUhgR60qaLBEoYMuGrMSDpnJ+Fw1bWzgDAUd+
UoEg57Uk/INiN5LwkiXMuAE7z3cdxi6BGjIqzQFrk0UZ9wtgpPsMH2/xu/SJ+a+/SoArsD9ZsY0T
qUDen7Lq3E3v7NFyo5wERm4EBJKXPIqiZWPJe/l7Rh76cuTPOqQBWRpVYDJ3uYrHioC7WrpLbApX
3gha0EGxs9fXyPKT3+ypbSp7Oi4eeWTD8HRpLxKO9UycFcqQBqyWpHuFBwpk1QNEddtMfaYQ3hbd
YvhVcn9Q9UL4oqMq+vyMjByM84tD0c63pZM7ff7vNKdH8XevioVa/dOv0J73aX3GVVnV87L89anj
jUJwTEGxWxlQjCYxmCq5OkuOeNs9N+Q2ypWSQ9VvLC0g7R/vOKRHyi8kChguc1bdXu0Y4W0z/hh8
RgkJrz5Z3iWS/ypUeZE6XBIxraYufz0xLFn7KH/E3d3JN1U5CBfTO7RBLw/6vyQKoXe/s3OWqmOP
71nWsFUI+8sitRXIKms4878HOOsSERdgLQo+RV1uVGwf7Rz6vi/lZsm2QXzQr2lT/O+0rNKDKtB8
JqFm4fXJlahLguP2FYqucsB8KGTcLuZ+RJ6psr0QrSJyLnBRl2/Bt58Y5YhWuH9X5LaBBC7gZhWC
v+9nQLb8PvB6ybReZvPjmVTERTRPAvMS//Jo3b/gl1CNtgz/9aQ762zza2ULEHUmVUaIqFQe8TLF
mH6ZcsisnHYXKXPt92RFy/r/Iqnf2XD9eDTUAEkktpPhdpkvItWqaXFn922zlRc6hBz45rP8Sp23
gdY7Wh+N3GLu9n1TsHmEoGUVz9mgrjZzTgxeX++JfUnXJSFhjlBDee0qdvmDi+wjMoqwW2B29m9V
6P5n+R/YzX3paystO7lGKz2rDg92JzkyD/1iUwQjIc87OLm5VobwOk9YMCqv8VwgUJBuk+p+PLRD
SZVN4L7oyENRijRV/acM84TCR69OdHe9NB4KG0tZfKldjtQfOO9/hDFoCT6oGLGmzZx+Va6rNjVU
09/NiZnrvemZE6SC5JJb7wT1AOO7aRvcs4YRPDC4asw47yNYu9xiIVK43skkWfJOnicbN5E+wILL
mloYOfH+h+33HLkPhgjKDsK1SRlWi1oE+LRQ6ugbuiBhahj8EjPg5dBdi8TV3ajTWc8Up75dApFv
m/TjzGqchGdJoTxZLZ3QolJ5/i+1sxKtNSz6cT/xpdu+ioK9Mm1PBZzdMR93rD0jNFfyEazaiNjT
t3kMjeB/xk6SLFYjs9yWmJ29bkNLrakEHcihpzpP0EmYNEFYSdAzRRbQ9X2iivh9v26HcH6OCKRN
XBM8ryxdF3T32fk7clSCyigH8+Zpn/utK71c8h06LPZpQY1Ae1UJiXuKZMUJT2FWkMiNjUwChE/j
6uk6MacnEW7B6EAvPPZGL40spC3dUgwjwxmN1v5dTDKQnovnEck5VeTJyIvKhuXk0Ls2BxuLnQ0K
bXY3AtDUksv+UQOh2VNbAAn2+LWbkgWt5pPROurQfmmOgCA6M/P21udabFBiwed6l1Yt7hW5xxrd
5K0BOtgPi1lIsujsdxPNCqSuZe/By+nAm+WsWaKZbWyeOMSJxHL5rHBE8rYClR0y+QoIOiMNISAL
9NilA072wtEGEfJkU/UNuftfio1eRsvv4UcLDiXfrO/tELh99KnOIDDz+RwWQP1JrDNR0aESAhRu
B7oqbiXLxvfOb68PHXZBEgVxl18yBn1gOZgE7iKB5+rwwM1lxS7Fqfr6EcJfR+CtPc804aiXLUjs
ZjjO8NOajhQ/ipAPWg+6FWfJCOGMmpV9eRyRDWQWgQtlShkh6tBNDT+F84oAF9dmcCMRU34Sak3a
aoIf9zpswXuU/BZ66er75jwXam7MaQQCdFNgnDX5FcadDuM1OhEsKzdW3ILeNDnwEGMoMnd+Kf+X
3a0FHMnUhxH5vRlOPw/vRl8FxI9JP48l++VROkyXzsF+4QXX8hfoaRR6m5RgHP3eAZn+9V/n4rfu
LjecmStktFIhbTmDMi8iJWwMvgo4kgA/qWbMFvMuzS/ZUqRmLWVGrFoNKjfPgsMR57ft3EsDxb+i
i+DCtqRG3KcNagm16x7eTOdXwFM0QzPSBjAgxQw4CC8tF5GVaIKgRjrm2SPQKQ6CaLHtP9tl8sk5
HRZhRnnlMs3VWLBMZJJ1hfp7AtGr7jhve2+zZt+ZvHTZCWu3OUdS5NCdHSk1+oGiFJjJoLjRIdBr
U2Ps6fCXvdEM7DXygI2MRqLFzV5Ois0zkZms2egZbjBi7c9RbKWw60f+a6PsWMm8kEAEa7MVhbMh
JHur+0Hmd3qWiLHZGkDrvvhkh/ZntYMJmphx1noUQnSo7on2MazBVglANWgUe00o+8AXimsXv1+y
UXekZ312GRwJdI+tKIj1Se9qzCdLtmXOeaFl9vGp6k23UaLC76VHSK84EOvYMOb7secDjkwYNFr+
oGeEjQJmGeSBMYqGLvpAiy/W+RvtnMLPLocuEZGqq2YV2z5jJsUq3clp2XS1eZ/kP5G0d8DVyCgA
nEHE9ZRbt7M7uk9k0TB3p1BKv5bS9xikDMaCuR0AOjTkzpsjyyVDwGoFacDzzeMvOw3E2UbxyELK
qRJYrqhtVT0kV3NQyyJJnoGFF3HH+xedrDOnSGAFfxtpFrfO+EukEOLS81OGShE8P0up/QEHAJUP
WTLC9mYaJVT/4yrXI1Gnei/nwYhQQaE1M+d4Azh8uhUh0ICWEGFITBOk5I7Hx3Mhnb9qzsVpEvH9
iYbb2GyWLA7yGHBIbpFGK4diHc29V5vjuMS49QsKucAkJdrWawvvKYKoffqe8731bY0ZtfMGtK7Y
gE554yT/BFWhtWGE1KEiA5ODRATl3FdZx4woW19pNslKrN3FGoegeRcyi3PQW6+tlZBZtH7n1cNW
PWxiG7JLLiHgJeD6/ZplUuWeH7KrJZSASg4EtZ0MyegcjmuNZVhZyIh06Pd3nOD5QeL5/pPLIe6U
q76Yz1VtosS6DRPALrfvgFeltlAFU6uWYh9D+Gw1t7j1tb1fy9Hhd4kg12CJPcv5IEYJSoH46/7B
hC+3QtQvZLTVBoYq8DK0AerRTK5y01R18ufeBmG9cg/LboWoh20wtXXbMcccBrGmtBHvEA5aZ6cM
RHXYaey/mQZeb72Yfu2J5o0RRp0CJsBwCyWcHz/A5p6/ho1rgIwsUI0Z6O1fowOBEILmaGwDVtrW
xgh/I7ipg21Ruq1WL9E4ew/LPEfwI9x0ire9A7oQZYcKr5hXQGAxM+l7EoWW71AvJnTzyP22iSvy
0nFB5hapKbTN+KRtF6p4N1nRJO7hVnj0RkZh4NmL9gUCa55hQ2+Rwi6uKhXddC29ZQ4CaEbbcmBN
ZvP5Y8UlRracRplr0llg2qIIYqol0R6rLBuPGR5RgaX+lksGb+seN6aeuvAoi2Q3Jwc5bmZQtmTz
NDjWClKkBYMf0rhJ4BGJG5TWEE3xMuZeQJqBEquKonPdIfAAg65M1eiP0AxdnMcIpRrMQjA2aKZy
lgfDYWJn0pGjJ0UdAnvp4gGjVdAUtjroeZl80HMkdLI9JEAVRo4gugpCY58r43vFYQAMLlLdNVrV
K5u+qm8XBiZ7YjNGA5kio4oEhvPF8xKOd7bdEvpiEhDiygu+nZZ0+ON7VR5iqgwbC3qqqZdAPT1G
VEUo8FC9fhL8HlKVqQKfJuT2Er05EhJUB53POKnFYP2aj5UKqzK57xi6zPZgRELGy9Bcjmq+r/n+
yTi97NAUD4H+J95tDS4qBaf6nLe8wty5Mf3CxGFlXPX2g4iYh8NRoX23IP5bzxMBnlrAuw4vP/du
dYOeTWA8RJAndavzitOlCQoBsXM6g+d85LROk7uNwv9+YNI3I5WnmGeRZIdKW+/9P0Nd0lHMQkNa
TnsY2xuzXaRxVsbjgGGr5LRjcwo30rZ3GV1Rf/1VHZP0edOWBmdz041Wq/R2GnLx86Z89nX0pAMy
MUNesp+UMRnbr0Tch4l3vl2FMs3Me/nqINJPLmCioHGqIt8VIMIZnAZ/RitN7mmgmxOn/9vBHtjo
GxosHGFV6kINccjv7gbHDIS4jn6ZewikrDrmDgGcYBBu/jUOAb/p/pSYfrq3AR8MKDYmeMEz3sw6
FDhBBjn+DVpJOp69cGNeYdRZr2sWoy788tk9H0mfVcZSosbsy+hTC/OXWZ0LD28ACa8/JWx7f93K
D+FC7Ku7ERpShu6rDe9RZbptw4r+4bwIcK75GwGdompfyfJWRFoMU6UpAQy+OcWLTi9pr48N6TCW
vY1KgD1VExdL8L8PQY3KLfAVH8IZwJOrJbpxRBxvg/55ix5fa3FFc1ZkZ9qv3kmP8JxKoqUzpVht
rmAEyVy8z6a8x/BTQw+u+ho7MMIiddDHd+2RJtemaSsaw4U+eyZP5lhQs3OUnVFmZbOid51c29s5
Cem3m06uAviaOKxm/DbGV8Lf2qzT6/xCuEh8MRDQZQUNMf7MPSIYG/QEBCarBjIcKIbBd43LFgqJ
7xrBch9/QjY5O93NHBUGQD8/GgubZC315wcjiis199GAmerwRxlFVfjzeruHaEGI/7XB1oFtx/Gc
/6oEnhEgTx17Qx2IXu50bdJ7mIo29dQAFN21BI4ZZevBOLW4QNe7yrsNHAiO8Q83dwlpprP7QgKZ
cdWzkX0sYf1f2c4+kVYJ/MEWk+golSmvYaAHdCmFiMvJ/xlP0mos7mLiVkVJuI6p76HNsbV3ZeAR
PV/Ua28jbK36c8WtpinCPHVHlkH1+3y8+sHoH4ga9fVD38lWz0HDZDq5ptoAQZoIvojgO3wJYHUa
VlQS52UoF6K+GICOFrhMpcyA8bBWQUK0t/xjKTZOQVnbbYYL70joZSNsI9+ao9A3mkqi00rcEOaD
alRV6j1VzL4TA84jiDDUG1qBTWcIvoTmGbm0mi8IRBqdkE7pIbvg8Wd/2pVfPkiES++7IeaH49aP
SMevAINZ3XBYWnwzEndIJKjezaKwQf7sy0IiFft+lon3+25JawMBUjCRI34h7BE+HQ4QykYD1KQw
FIjBKR2y5bnrDXFx8NmWGop8F0PFt/bIF5SinVeV+i9DtSKHVSEHUgQovA80K1Q1ElPzLsbebp0+
OEUc/1VccrRL1hBjXPeWMlRZEtIrl7sCbpTk6extx4fuX3SAhStsLXvWYr/dtXORwL1bDhmK4+fM
7GrZrchzGMhUh62rRC026cHNeaQ7bmYsF3DhfrRoA20TrEaymA+VcunZUQfLW9wKeTVZ3msnCYFe
OLK0B4ZJe3tR0yzLicGjaMKpQqMti1bx3Jl+o+89j/Sh30ywKX3St8t2PsnN1L4AaYsvg614swV+
64B9PMojZqno6SP0lOb7R7PWwBVXRE98sxYq7wCRwOBsOzggUIisvQtuBNukGN8RBJvMz4/tqb/s
IIm8kgVDHafgDuxj5eNrrMJ/o8O1XjpnSo99QbzXtnGSX+ReJRvx1cwsBxzTcV5y5PcJh4RBCJTe
WXFy0MAYiEGNtw7oKWdCAvwcGhZ89EcRVSOpuWDG0tMcx9b/LsnohPTe7y1gemFttyjoI0aOEOF4
FzQ/+YyG73yCmuTkU9X2b9IKntO8wZZq05Xwl/KQ3+aJ3peAyvhbYPueSzs1+Dziy8VYJS0Gkcqj
3qXVnY9OjqKxclOe3Mi/Xc2eYs1PPZ4GScwkAbMDpT632e8ZjgnK3pnv06dzyVVx8U5rSwimQaFB
jfO+S2D5Cb86SunYh6phsb4tevEzbAwkC2CUGUjq7M3bF2uLX9vJKaRqZCO++7vCF5Bx2MtI81wZ
L90aTG3BF1f2WN6PnRT/t7U6a+331VX2tME6wDCM7CiBOhCR6jaYJ6R4+njBL6Wr6n/fvp2g8qpz
AOAUqgbdtV2ChyMEnwQ05lcn/XD8wosHJ7UtqI8u2uCVjltaTuy1RmX3pPdbC54Fn+LO7SPoTrbd
siSnl5kpf6a1famYPQglapmLkILW9lH67+KZo6gqHe4NhxF2fJvwhy4cociJYUTTHGgIMKOAhE+e
PcEjmqcG3a26XACUoDr0YoewGmf4yr6Ge7m2+3scb6wvMbptZNVuTzjtj0Xx9vsfg1v5b6cXGKvs
dNrn+cPiIT4+cMBDeVpa2ugargjXdMv1Q37ACJxSNPcb1afgkWzNnVIJCMP3tO3jiYZCZqnpw+Z6
BBlc0jG1WWLBdq58QVZsdfGcgCT3+l+gJxDZm3O0U12hxSc3UEnDd/W9UCHUhEKGY5hjS1sjpDYM
DNXutFqAJZVSc3PQ6lrUnIzVcyPrm4dhbXbepKsy1XPVaM+8Q84qXW6tnoNUcYjC3xdDg1XQrZTo
Guj/T+2nZHv+94kNPzNhVkyUKHw+Lh7g0d4mX0OMrYzhAlF/zN73fd4eJeEe+eQ+vDw7nJoUCMXQ
+JcHUM+/UQ2NPleeNQ3ZA48oxTM4JxrINHtNci6tiL0LDIGzCPoQUrx6ua3vzUDY69Fr3Bj2g0CD
3NHj5+Bw6uAcYr9jiwY75/PQcl3tbXdbk9gBRgtefc9xjYZEyVB9+7Hx95tly1fqfSgvZ1OpFM7t
nBceAjE2uILbh38U2OaQtY1QeEDF2595vdjPNvjLkCgIwBS+Nu4AW6GJEcsptEkfCf8xd78+io2g
sych7WxH682p3GtGuXSyP0ShQGZf5OYqNngPylzJvKa9KzMAZMVhGOnG5zXT+nSAkH3hr0Ax4awD
0oTCwvdRYvoUj+3uRAoj6HU6tu+bnCXI9Ac4T12/VfphDx+evT/QU0nl9CX0hy/vLZkArN6Qd+qE
NVHmta/EW1jKeL0qYxPGCmyfG9CSfY0GntXOx37igcrw2rdQlwutY3Hs+ebmjLd5PAWiZ3UCD8k5
o9cuSKWMCY9+sz9i2EBo+Svsw5JHcrrv06X1TEhGzFGp0H7TNBWXCtS3qczpyBrRjUz5ttdJfEHH
oVze8MmX53lWGEo1KN+ejkbtDWfCNz7nyxt6afpYIjWMMMx7/t0U7UsHpnSh1avPgPcoK3yuzRBK
ZP1/aAQJkJFeXLm02/dVa/they6Pr1B1ov1FX3Mk89PE4kLcgTNd2i49Ca1bZBdq/njZTxhOuOPe
YDQ58BP8EC1ppVjzq9w3v0vfl0iEeDt27ZqGE+iF+nKX/0cFwhnwJLdMxTf1wsBIZisMGxsW3WRY
01Ofh3TAa7FIFYFjzpAFFUNHvV1tWOmcsrrgb/zpxPqRlQcTQ/ijFYgJQZlnzYdpYjA7lAaTWsdA
UQruVRD4W9oTkNdthiAZwyYjruR8PO61EHArRkwi8RW8hu1b9FjdO0LKmxFkCVvSNBx+e/TOgarM
VUZhJGEBlZViDRFeWdrpY8BBGUim/RW8nxeIoLT0KI24MiwWH0shjNXKD4gjFwEladnHmmPCfwgW
5mc3qWeeDsKfpBb8N+xviduoKOvp0MNV3xXDoem1Ytif1onq2W3dnSEjuIRG5xx2p2HYtjgnkbu2
gTE+9unByFWjdX7rjehG6cdujX8V9ps8ACoY/rT8yKD9USeya586TKRH0elygwWjCMTfWOwltuuz
a558EBfDobsKzIT/mGo4g1aCi52tJrCSvA0+9bnlz2+vvSytcmvWltksqK9lC65do87vQnPp6OcH
3Yd8MrIT0pEjbEag0rWztE07lgAR26pC18NMw6C6Kzv9/GIZTxsebM7h1AP+JqmeUr6IR2UZlPXd
7yVj7rA+NdvBzPfWe7UrqdeuJmDwzHKD3R/Ln0aFIIVf4kAVNfk4rF13bpIZASro4+Jn2uHHu+6h
9vtRWbBd4s5u9bsY+SYsOaBW+W3himr+nLUsXkXOpHtmxrzm/Wu40GaQz7Ch2339KObcPniWh8C8
2+JtNf3NpvZQi2jCwUAbGYA0pkuTYMyXJegyKbUluHtoHx9toZbT7We+eAQG/tA0G/38j7R3AUso
yfMQi8pN8IojpMCYz+W4rgU9AS96jNdIneupJKzODn5yYe3WGRfFtCin/BeB1zvv3bZI3RpFfxEd
xCQ56EhQJSQ4IZe9incaLCJHpR0Gz9lkE8QA2HF9Zcy8CN4DdW/OAGaJWVgVuy+WWGuGBV2gHEPV
ihyzt/otwpMEH6fXpWuWil+Ll0QM23ztUL8Kv5hNTsEA4HeciWPoyX6kMV0pQtRrHZRbBMlvy5Kc
UFAInCOJzKqWV1orNQMMK7FliebQJgfmaVODCPhCOqmlDukfRE9V9lr2vs2eAApOh9zuGFuVdzCm
D/FT+4iLEO/RvMcd/fv2HE9RU6nG/lFiLAlQFIlspR4Vue4jQaioNRG8ZFlu7vQ7W+e6/GdaSWqK
1WQ7ke0N/itu60I1I3FV5gTPSMPrlfeKdzzAYnySoXGHkmjTDftTH8ocxiGCBGqwx3kLf/ihTY6l
UDejGDOZlo3/S1yxMFGBzAndQEymMl7L42+XPa8dH/JOXIDWXMEDSPcRsT98kSLqrfkFYc75U6DI
pTO9m/l1btdca+xCY93BxB2f+j066CiSsTTSVxPgnhPLGNGgvxha9tyEYHYYMVmhY9KSJRu+onEG
ppq47dxKD7Y+Azz0rHVMeeHKkFZAR5TwLM4/eIuW3lnyPA2iXGIWvvP6TOwaC8nnbgaRc0oZUm6q
LJ8GWEsjmq1oA9jj
`protect end_protected
