-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
iuGvV6amwXXy4MQxvPYEIuF5iBLXxnT9uOpqKIZ1pdLo2lZhTuu4hgpxUyB+NM3K
Sfz44OkN3E2Oro5aceYAHlls1J5HmuiDrJMzTtCe4kOi0m3waFj0GF1vuWKHSgRt
Z7jN4moW/Tbfb9hZv+uE9mmY1u7JefDBrQhaseV6mgM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7322)

`protect DATA_BLOCK
7HP/RNxDzR2Cez6K//u+Wa2c8YVGgMJ73m1f3Ch2O79VZcLCwThBUfxvtauafRp4
QTLHrwsY+CkzY+Q0dkulmY1F8rjP6J7n3Y1riLh2R9xoPUgs9KUqwAT21mBVh6pA
ZSqQTNqSqIkq3iLlZZ6lp7XY32xXwASfrsdA87nnXQzfavkIOqztSHCfkkK9Kn0W
0CufAugltIZuQOfReYZSyIUb8rTn19HlzSp1x1yV5fddh/QFmZy+6hN94OHh9qHh
16K4XrlJt8JHHZIl3XVnHt4HkpnWQfhNhjSUzPrKbhHqdLgLCPwznrx5DvHY/+7D
iz+IhhUWMA4NFtHwyy7Fg8ffvnBdS0BcVbHTzo/Hngz5n0H+Ni5URjBEpVbEpeUl
CGebEv56TY4eBjXO2JFmCHEGMIEp+Xv+eyxJwoAdZKT60ymLrYbaMww4xesBhCtR
FY/lECKXxeStv/nTGj6jL/jaoN0f+TcmaDJNSCQr8IIrYLN78xvsHQYuMlnt3LN2
Pp/n71y9ECL5QcbkL53MK7Z9nB44w3uKITL1JbyDP23MbrHRRq2L/DwSGYa7uVYR
3ZlYf+KlHxmEhHwYiimVwiMkoX+yELe6ibryUnEZm24LrxqYnApnE1yeQQYWU1OG
8LgU7KIxh6gTZZjxEBltnFRjvcBv4HlPCbUk6TjcXI8cU3nYbjiB2477WTxwKstb
Lr7EPNDD3FHc0ftrJ3twooBPcXdb/srdiw9mIKHar3RL9/52S5Oqicx8dxCIkcBM
qdNzI2ton7Ak944335qDMyTFzIsn2q6rHh/tE1XnpSKq4VfAUgIBXu1Vsswm+ygh
ZL0Whnc+K1PY3FmH3tHTaTGJKv7Yf9s4Vkd6hRHg6zm+ToIKCnEYBjImIDf0o00E
XSj8Z+GAKJUyp62CVpD2CNh5xV4Rw0t7eY8OfgEziRMUzSqjvXQMocIXZ3UWgeTl
fbf63Ps5oYE4w7pj0889b8BulsyzrNwhpd5ydl4+OrgslPdcFY2xTfuG0mRQhDVg
Avivtr91Qn6D0CTrcLYP8pmdPK5mT1TbiJ7HunvQejIiEfDxCEFyMq6lpR3bUszC
zY1tGTrexM/iIilK1ipzKdY2+RyOM5TS9in4Nz3WPL+2Gb8wkzd9HEcg3dHYHxTJ
NIjMjidQCZx0RGtxGouB8wqv3YHMgEHO/cCXGTCLcFibYXKxyHDFleyVdV3QQVs9
MMTMDM+f5tFCpI5GjR0SgZL4IRpkJmDppsCMOZIIjiRty6MHa3WxkjZN0+rN+h3s
F1ZCl+cUrJ9FR9THedyZh/h7cv0YXkgVyKGtWMH6hLmFp1L2iZNgGjl+pLOvlptR
eca9Z3bzLaoHV/ty6pmj1nlAYTfn+rRj60wuQCjCFQqIQABCedUgqyFm00Hw9j4s
G4i80m+IGcMuiDgQJl6cXbq4KKX9VRMQXMpZSQQZxrScczg5PThrrPIdrUIEAQ71
/WwfIZJ2cM3pKUMoiaaWSyXzs4ocvaaPgscrKOZHrRIhxejLenayDGrXD18oeZLy
FTLs+WerucCKI/Uhyj3Hbkf5rEqQcomMPvcPUzpIqsnT1A+QGxUQdmLjEwZD9mno
ncjVK82HA8rd5IkNue7yYWPKYVEpfWj0BILHMrBWmGU84dZWSRUXdOEBDselWkcG
v4vFqolYBYplu48Z8Au4I0cZHc+O3iD01/pbqpp4zY8bjWAc/pf02oNFc7UVXOTR
cJYe+dQrN8sA9FwntrG0DVgIVI3EZ9v3GFyLdut6j+Qs9iglQoHc6Bx7hS78hQQS
1cooWhGXPMbarzvb6T544NRX9hCT4NEGxkTWKWVKQFv6XWpwntUFXf2lOl5nNFpd
nBKonrwiSGFey06HLgGXJnMsqbDLA+RH0seOQJ2UpkWNPA5l660Y4NhKmWk5gnOm
MbRF6m07t+GYLN9+mNOwdRQuE61Fh4xPtEd0rOTvQqSNAtJK2HCuXv8WsqTIlQD4
tDmPOznUe7UhAxZzOP9cm4QuKPcRzGuxQbJfc/dyyrgtP5dLr5IyIsxrWMBTto89
hUe2RWN90Jn+mmINl/PdxaTjppcS8V0pH1jfAwJigY4Hw8uSlQV5GGi2LRNz/r89
ICaity3EADuZUMAOGSb94CN4z2ecYRgwNfir0BTIc2iNHq5/NuZih4Ks6qTNTn89
Gwvgd5KVlpkMqDqfbKBSM4HgtWUSFQePZkPJBFi3OPT7T1Y/sGlLQscNeyV7VuEt
puLNIn9yRgj8+Z3/wjkwWwf1ShvglEyLvvv+Cy2knaJ2q5rN5w35TnoUfrX8qNLX
pxRrVexrIxWXKNWqKAsIg7ScGRHIscHzAJFsJp44ASmnZP0PLSM85QWmvC+/hP/S
+tVNga3X9+R215ibXJyJ9idJaXv41N61jP3lZTUr8jzODBwVqqx9Lc7dAvXWCeIq
2DP9qHot1P4r8ZraYt8CHfhQLYKGiEInmDJBvKa1PTSxf3by5/4t2Pfh1TDDIXff
9QhpQxbn7OGWPrJL3g1wR1vWXtOHdZg2RZ6SnRltyaTFAvaGcqZgMVHqRAE6aOL9
QVtlLssBTRRjVMc5zF97YMp0PyDfLz84jZAj8gxUUhTWWSkOrJDAAIAJkICu/yAJ
k2GryXkyFQvStoCEJCWooc6eGdUlzq5E5tQCoNmRzRY6o7BvpY7PFHlqcCSh1tRE
z00xqDg3BKijjt6t3qq77LNEu0BbHnssFFsy6Rq/BgLE9PbPyYmoMAsaBPVTZKtB
9SZHWbzt7Hj5C63Ah2E6eD8WOHOlb49ivNN8DeAK6whV4vL5fBUIvbqmcwoxUWew
HOpg8kGzvmyib/8jCqfiRo43brSjafvCAl1aJC0lSb2VJXBzvd9eohGiN4x9VDW+
ExQi7S0dMTXhoF1G+SdzDHE5eQkMRlxyit5bNJtafm5Mbva4se5P5ecElO1gWPbm
JnOetD+EUzZZjrUoG8BdcDxaIay1EFparDwiW2ZMR6i3fR5Cv2lze+bzGvLN47oM
TPOH+GKtzVArkxfjaCbN84KyQCl1g+h3fDA5JKddYHgEBzn4TaICDPYKY4tJXzNg
dtxyTvyRivdyjm1cJH2O3VVXwhXVxw5Lxyo4DSFmNUAED/Vow9I9PG618SCn54KV
VhYDgCfqGAtTEXsLHcVumrmUIC+hzJI7pjonInxG/gQitt5fTmLw9A0bop3VCNv5
bZyCoArV8u/0hxlWwTyfxM2Dk6BpW7BlccTLFNaoZW540lzhBpp1h15T33kx4f+w
u6CoAo0ZP4aRoQZJz7Zyl/G2VJp//A91aB0gN1TrHgPtWbbDOWx5WTfaIm4Rznme
T0YPK+hy85RXWyqOxw1QUdh3RA9Hz+BGPpXE7bm7DaT4Dyzrwau52/TnbocIp66P
oqWU8ygv5UTUJMICF/CnebXObIrc6sIuYkseMqfYYx9LhTIKVqR4Dapo7TnKHjon
4kDugD63mi87rLWMpFhVQDZT53UbQW5sQPfq6dSbsTXRfsSlYALDom8Sh2TRG2dh
ff5+1/UMLkM3tSwVKmLYm2JCoI8q1tFYKgO53T+Nhkgk60cPrte3jwIrIsVHk02j
O/9FSICeMjh848JFGQFtlbbNtgYbGs+dcILAGnLqVKSjdsl/UXqjSZ7qLwlOXbRq
c0EMZj0heuH4/Vvq7zo0ArQRY6QuwjqBxlsfvdreOuryZ2zTl7bYA2prWNcv1dDW
0XW/AaazM8rZcQc6K4ZGSjQaXRExqPVm2OhVlYmed3C42WOLtnFIZA8cadwcxd/D
ptH0yM2bvzhmyC3VYWuCuVeAKtN4ddFDo9kIqE6oumKXhCIOgUcUsprCT+R5zCy+
TAMzmWHFcPoBLDoV3gHS0jHHNQhhB9dClg+ZoZiuIC0GSh2rFIVWYULXgV/chvFW
sSt9YX2GgIF9ox35MZ/MlO7/PoHw4yb/VPaasZvQCbRoIBOEQfjizlnMhFphZcrK
ZwyyTDIP7pjazSus6mJFc5pgrcZLtquGhHM+/BHBDXcUKwi4pRlQmMMtwqVLDIXd
K9wLszD5RZOqMAkkLpKiQ9JJR6Svarhlgmuxp35UO2qU5AI1MP0+udsNKmbkgynR
86dSouAYD8nJk3+ZZRPZvJJa4X4z/Rm+JJJL11qlgxqlAijNJBUyADQMwe1A3kxP
NtsWcs/Qr+ZwFl5oaCJU2bcM4JE2HVlKGs/QlZljQM28ehi5QunSGTIovmWg75m5
+mAciU6k+ooiGPCm2crLtsszvbpPos/W+8hyMSNvoiabMjqRTp79MBXXTDHg7xft
48vOgKWpP3ymSeJbFPx1pRo2OthzID5WJxJe6eUEfBfG5tBlk6n9yZCpEXnplXuB
9q+bOjY424zd5fjNbI9ZiMv53oBcpSj+PHzNT6b+8qEzU2sw+9e95gh1CFKGZtoS
UAOG6qHL0UED4u0m/feLkvhMN2NXdQmxsdoDOKVK29kppJt43IqwCzZ0Rx3oSEKi
jeWjZZluE2CTElW0nWlEpDFG9jNaaJ1fg9qMKCxgQHeErHfeDG46aRmkIBgPxdP0
ILRuslf2I0CKnkQANpUUEkFv/x5PZoz919rHzyMD00hRQk26C+DJixPLTWXwJgSc
74M3Q0hwmmsDoN2GJFxkNV/+BFc715RXKF7+yWxVEdLAUDrn6TOzMUzS919DH+5K
6dTNWHBW0UMwgxxtIORt1ze99OOIeujvQVPWLL+j0dbwMCZu3wUQOxg0Zjvh6AaW
et7DNa8NXa40PlKqpGFzFRB199+RSkdmDfR0eRZ4d2J29Z5y6RcKJFhhZImlb4KB
0rudvw3nm8JZZHJW0vMChduLGscn/YL5bgj/x55e7jfX44S3ceCMFncKFNyhM5lg
I19alhyz2sTYKslpWoOwoFYPluvgTQaQFMM2MoSS/FmbLBVa+3Y6wDnkez6LohvV
ffL7Op4dpaJ3N4zgKzDvQ3EpUckOfVRoVGbx5CLOc1MqsZ1iWex5APcXX37DI3ck
tFmKEiGnRMI3VGnR2/YDMbWaVzImA2gCRJVcd/qhe/zsIRdqe9Kb5MwYrg56OE/4
N9RKNlGyhHFyDmMC7aV+Yjqs7J04oszDCeVMFJC0/ZHHIojNjTnY1FbUHy24B2Fz
MEfzUyXvqvKJ1G+b4D+Iv9MMRBCy1YkOr8kiKxOJS5lT4bvj11+2BrNZZaiKkLsf
z2MYp28PhOK52NvXd5o+bdtyFwd67NQIncWoLdohJlmU8+/Ox2eeRGXRMzaws5Ck
Vd33uU2VDc/HcTfhdMb9Rda3XdWT43PXyNiqYjCdR5XNeSs3X+qESrD5ANSiahWe
tFytCbwzgBlMjXYCG23Au/ANAhh2yQ9vqqsmWM2L16r8e3thyyQEm9Dl/WXJP0dk
h68spS34gYtnwXnGccCzhP1D/ztxCXTzmvm6LAX0GWRDQZjh3bVfTO+Mp2xT69pZ
QHWAuqcasVtN2Ph1beRJAth7MpnuLL62jCeEKaPOQv+zuzBdrQSF3k7nYRi2XTDO
omN/e5vyB2zjWHSpOSoGUK2C5AlbePLlTB2PMbIRPKmsZpRFHn6aAB7WHSaZ3VJG
E8XS7vvEYSRM4JvOjX5lm7CoO5RDzOk5mXhG2HJADgiUtygDJJrNBC0UVMeEITrA
AX/WksKLt5DbDlgzOkf1Tv6c00bjpU//gDjOOPcI/3PMX/LqZl5rChD7XY9sEuXC
m/gvJL7cbLnbZJ37ZkwWPZQ6HW/lFdCQAGIU8OWK6RNi+cWhghW3vL9hYaLakpDe
d7jt2tLZgKW1YfOzezFdeSrhjkvJYdKb71y1Xu6+x3c1oqX76Q/y10oOYpn4WFqA
fLSDJOTwcgU3XQC4HdGQFWVOvdlHETlcW1NyZQ71QzEw0P6MB9JHzzrCSVcB0VfW
Lm/DkQSDmWmQsjx6URs+tUgvreVaSTH08use4qtK0X+jIxxtCWsoatCjBL0GFlbY
iB+TPV+RgJeFy1uWJBZ1cLqzajDH0wUBuRi3RHe7/3gjXPqElUVgNA12gloswmMP
i/AnbasPXW5kGUI96QrqUccLqrAHzdZHvkAhCsbC2C8uqe7Lwh8A9X1W8BYpRULr
HnuwHngrAyasZr/Hk66FE5yj5MHzydBatybXWqbWnEvb28WbDqrjinZjx8Nwc3IR
YgVeQ+Cs10wH57w0a8dtfvXY0ouaEE+c17DxVuYlKzHWXUM43aC5oJh7EMCMeMvz
4o0TE2R/sDpNv49YziUbSJ8Kx4KnEPUQxEf0YJmHNEJmYimoLKYlj+DwPEYpIzTx
a5IMrP4RL4kH0bLHYL274+EOpmvWAdzzSS1fnQ8N5iUS7oeWxcVT6r5TkOvapRvN
Scdqzc1QaiL0Ai0LmbJD/RrUvQZcrCqTxZqJp5V4kReBhG1klZRpKRu/SOMsolxm
nKfd0vj4GWmON9t2me3Ev8LeIZp+xBV1/MEdb8UDm5XVeCX9vx0pu1ZLRUEvB2AS
P67fkTwKKZznjyXXNz4ybWZoo1VmLgJk2kGD3Wv2u0YDSpgAeNNyL7Y88ByEQP8U
U34Za7EUhN7xYaeusoGviIfIWmNFA66D1ByVK/2lSClzpQcSnNe65LA5UNYtlFTj
CMJOkUgukBMr5Vnfz5cSf3wBAvhU7XY+fZ1qP1hNwH28jZ0H3gSoF93hmARIL+9b
HyY+8AR97L4W8+wKI+S6aiH+IV1jpNFUFdQEMdvCjRrmEtd7c3X0HoP5O1zK5UGa
jU2CL7eqGlH5VWqp4kmIkg5i+mcXUVBmcfBGnb8Fa2XgKWP1SEkH+nBjJRt8nU4j
rR+AoOOcw+sUH20rcPIMPa3gzUF4CpM6iDAsoOn2nboz1Ov7TQ7Lorr+c4Kx7/Cb
rv4i4ikPq/vc0ZiGWa1LLiVT6ttnZdiV/CPfF7ns+4zr42LFG8h23OUhw5fhSZCO
JL6mc7t8QHEUMtilUzE+18cO80NZIZzniWwGaW5Bb/0fE+a2HXGzcxpbV/JXNEPl
NF2w8M5VgQ2w/4lDPThPFq3Z47zKHn5DTlNmYs2mUp4Fy+HOj2BRTVvHOtdq+rgn
zn6cA1tf50bYXgkIM/axA8e3C4BmHq9fwEQ+0+x9TfLnjvO/CpI0cLKAqTKLXhxo
PuMcyNvoauj5f19t+db/HTmzhX9RkIQJ67FNLmv6quUf/beWRUe5OFwh1dRCNBF6
fFY0xh6BIgDLNIK/Knpw3oqUUUf4Y7eN3qF3dfetdHHN6MHIV5iCZEc0u0bnvyLC
BDnhMNE9kb8tVyo8OXXU+NFxJ3epAc2sQA0+13Y6o86aWTJJ05MhYyHCQAx1KEMd
aPm4E0+NxlpsvwDuzIs3i14HD9AN99Bdf51jQZmXTBRYkE/IU8gqFYubccXk7Pkb
5Kup3CWUrrimRU/g/IiS2Kqza6bjg9g9A4uK3C7ex9kC8fpSz7VmuU1oEmQDrM1l
gy/8iDyeUcuMBOoo0PObwdYbKMKiClxOFNzXUsDkSj/RgxL1sLq4VHcSk2mT0Dr6
/960GF7jVesfeQ7Y0Ej8EGDqYTMLJ5UcrOMQN1UCdMA0cu6nPDskRL5qBfhv8GqC
tsGjcNeOWQS78ZjlgBIL4eFaX3/1qT0Yx15b8yk2x/de+yRUabJj830C7AReWqnC
vwuvBCbINNf7a34JF3Q3g63ulM9ruaC+ZgpkWcFuG8e4hDc5XUm87EiTvoxYFXzz
0Pkrw0J+0admkLFslHAo1k9767U1bQCHWl16Cn+HCraRlTcMZAXH5UPOOnUuGHBF
GwTbOXOVuNnnRfzuGhB/98P2bFDfG63eWWY2Ua8wzM9oSzQKx5EmuQtD3FUcYtrV
RidKk+FMo5hn8yqrD5rBAIQIQFBnUk7suUoFRsIrNY+Yk23ePQPrdyE2GMqHeNOQ
6qh9ugVhul4imc9qRZiFr4tp+4ysGRzCtYLH2gbT5Eig1uvOKks+zZp6mJJnl9zD
FCOOwHkOBEVmbcegFIbv76owkCaFMvWVhlO5cZ1pNksP15nmV72wT/r7pmJogUY0
5Bt3Pn+JWRW1YEKDDOt8gnH8DWxwEoFF9vHnqX5FwaJ9mUBdpSTLUFwVfdvtVh+J
p/eXjek2awpxa74Qtfsg2R/ZnluEWFekOO/055TLnUHDusavb+QDKHIg8QAYwGf4
c2RouyCHRkO4fx5Wr9UVNIV2AoKAbRZJxN+Nwt8eSCOzV+HOtqNQVhtJzM7/hvP/
nZwiOLAN6+UioKTsUJafHbEWt4M3SAchP1NQMq+j6FqqF8r87bIGHb6ey7YPJYgU
wnCqDGLBZCZeS4IXxNBYRDn9QaQZOrPF9txzZiuFQHaNpneNrQV5rod/CTZ7IaTH
tl9XUNg7CyZDLi40QFFqpi0PQ8Hp1UU140NuCDi2msXHqjt9QJV/JMfdHX7VYsx7
NDvP0YIOg/RdWEJPdszPnZcJOqGDCtRmOV/VybdDgzox3OoO7fb5jK7jMRjIFd5w
FtS+CK51xh9tSW7xRGI0z+4O5RvSLmpU+AIqlBnj4UjekwVybWtu3mvsJyqlF42/
ivX/ZqIwChFLt/trykI+voDmx+rHVOFLeweLPGAmuwis11iTutJtkpCTOWtqodCJ
2NMDC9SKtC/gXeZE7E1/sOBty3JISFHNQWtDT8XNG4E32o2fsVNvjMM6cu1rI3gV
LgN66qHAdGTAXsb5if0u8z/x958TZdNM1t8jPvY/PSkgSmq0+x3F4nPs9C4EyhEk
/aUnaDSa65HNR8X8v/5xlTgESfgTKW7bgFjZw3E6AOaDCS1OvOjT5CcXNc1GJAQc
NyqH8/7dxHlwYfLC1cY1XitQ6liszW9kQ8pWOpUia/1WKvSYz+1XdNs+RFjbooxc
14GA/lO9bgYCamoJGLzQ1ib4wMIzIJR9WMuo88Z8RTAffwgtVUc8R/ZOD0VPPOB+
2/hfm4N/j3hv1Ku2CuWP44rXdTavsn3xS7H2jttY5iizCHK9RfGShCKzd+rKBhkr
T2kL1G3OUhEJAbdmjboq/2RDXQtJRGitVm2un1DkrMup7lr620xvV7e/8M7Ia1Cz
RuCzfV/ry4T9QhfQ+frWMJf05rvngWQ5ew4AVjhy6oQIB4gF7lcQ673Jx2CHt3c6
Cz0vkStwg8QTmXJTqq7CXf2NvgOSAEfb0eD10+xS8n1a2tELi/F7JC0BrMixEyK8
pHlKtouyE0Da/4HaGU/cDN66+LbBdiHtfTI7WwBjRW84NzWwALwzbp0ksNCKMrGg
DeC/JLni4PYHMW9n9qJ5SQJvXQtEGI7JjnQB7rZSno1MYLcV0DiVYUt7h44pNi++
EXefe32ZmqLhADVFQUBXNlfvrL/EwCJuEXqRQiPkk7qbP5TnyTRRTW9lE+G4P1gN
lV4+n541qRIaE48Z6ak5D7MadAfSBYR6Sd7lPr6RmR0bfx+QbhxrzvgWQvtT79tz
0QCDKT7HBub/VW0f36Ck/yjdW//FBXQqeastZWS2Cu0ntUChWJybEhxTj05fcddS
hI1kRj/7t7D6Z83HdTPUoBBKjGmzAqxzbGWf9gjooARcQbKyCdpHsL6qobW1oas1
+XmHTXs9mnifxT932T2eh/X948SJL8xqs7oceXSKjEzrmM6tzgrUfbaNeaK3i1t9
+oPtzHqF2eg9v/dQn9cMjOG3SzSDD7hJs+aUuuYvtn+AQlz6gVVn6HW+NPwbS0qH
rtvAhKePFFoZopjACDhR+6/JN858X0zjfg5wdvz6Yf/P+G/mRSr9zTdKzVojs0j4
4YyPTjbUpTppaqDwuJbwyP69cYAEwirUZujgzEeQYmzZ1D6u5ia1NYgmUdPQ6m7O
`protect END_PROTECTED