-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
U8IoZRytrZQErxrAZ2Zku+2SEn1WOptDtPi28TwG1ZZcHGAv2GtvCrQCk0CYVP8i
ZSyKl086z66Df2rCobFWhPjofRnVCxW9XxBdXzkcHNnjXFwYfrnRICZwCGTmW8hb
iu1sfr6lJb7vGGWRSucfR+JX3DCOL2tT74hFy6wKpw58+DEYa6wdBw==
--pragma protect end_key_block
--pragma protect digest_block
n6RpAijCL/OZ7U8vHbfVZ8re2e4=
--pragma protect end_digest_block
--pragma protect data_block
7tivugtwJqAJE96CJ18zXrvoF9SdnQZaadvoEAdWnUy9PLJ3z3IwFY/+PnP1jG8E
HJMcr+hXELBPLvexW4c2os091kv1NdxbrgFN5FVTtii8+wDgZrmc8Gj5BUj8Sb5y
MoyNMq/HWRiLWaBGS/WF/Fr1WWCXoM4COxgYos5d6l/vCrL8O6L590DcATjkAckB
IPqr6G1E+DE4uNNhglPFu+ND2AH6cDCmCCWQEnfYSYKQK22su/or0oLmAHp+EnXd
l9l9iyXxy1Swbqa427VROBPUb4iHwvPkDFc0arAOIFyrhPFzmS9l9FGxlnxBBshF
x2bOL2w/W/OyON3lNTlfr0lwKHNjmddzxbL+kcIYn+gB+BU0+iuAAfDe97NCWxhZ
0G2jDU+/F/mpSITn62NXB3f9ZAHptLOElXURbtOEBqKX1F9MVSklWP7U1OO/w9rH
Zhl5KtL5IzXO1+iQAINHrAXSGirLCxvA/ot/B/FScNu4TXWfaEe8/LVrw+UALM/2
Q6Z21lGf6MQ4xJ8wBmjizBbYdeLblIM5RH65SXF5mQLao5pf0SVXXwIIhAVpHJy8
G4/KXogyaEmQhTYqCkZq4ICyhQ9MGsHeQmygFsaxHboQjKmFK+gbDpK1/5P/iGIj
0SdmxNUylNV5ZmE5D7ou5b9gsuM9ZvXqpYkiwzKl4wVIvwNtD7b3XB9ft7h6dqGW
m/9uT7lwbwUAQm5hHOTXGJ/juq+GU/HU0Qxr1PFjra7xcvIfY0DY4b9pojLDEfWc
CxVMiayKC5LW+g9yZaSi/Bn/ZUb2/FAyYTrwcYytfSernM6sHOwwFAl4x1JO7+cz
JgMl+m1fnjzPfz6/D1HorShRXG2UrrE8Vdjim8qIM41tb06sNK7vCNf0gRrpv2wb
ELy3XdmTxiL0346qGZVEoGGMV5C0P3CvewCmiSB/OyuBjbNdsNROTJi9x3L70rhi
KrBpLCoPrSvlYfZe4ud8ElrzBbC3wMhJyDsKAuflIoa/Tf8hZLQivgW/F1h4OmO9
8m31DMgzDhqkYj1UArQ9FezA4jDiuJD9JHoItnmfQbxoGIOJOSn4/FEHVAVMz+bk
PWgUa7OlJbX1/q4btzYZVunFBkEN4rbofGl5BB6rAaRw3RU+2yVkjVz06gxuVNy4
mIUJBOC1VfGV9pwevNNvfYhAfOj4wDUM6Urt9C3MRwBo932ZnDU/s/Vzo7RpoNf5
L4kzg9QTmkJOmaG7WD6CmfNLKyB6U55k7gHL0qOJiK95EgaaT6pZRQXtnldSl7p1
mPG7i0YfrYS6TF4fWAVLFgcKxzGMRGiHgKcYA1nlVNPg41UrEfM0Tt6uKrezQzZ0
BuYIPNr2zzs9GJxTnUa7o8CEb1v1f74lQpgeeDZR5C1s0ZslegfwhUqRKlXTAxye
YW7b94Tf11RdcIIITrhWvhavg3tEXKQmvCXRd+MbAX5LZpPIOVDyvDehEi3padQW
bOAmm6l5xVCnPdXodyExm5Rw6IOQrLGqL9PTWbvcs4j4ypQ0RyU2R86SdHzapyHc
Zdv7JCO0PUmLmTKCy+fU1AnyJs5/jGsJjjwxZC1+2iSaVnS+a4dvbPQROsPPUJST
es2lTUoBOMhWnodx/mpqUufvVRBnPvDA9JtP+KmBBGqqkxNukIirEbOFS7OziFir
Ijk1hclyKtcEo9z0NOiEmIedTJGktjTebm2F6by50nbSwMh6axYldXD/myhrKfQt
Q3V7YboWPKaYxkMUkvDaREIUo0d0HoobLUFmCpOn2zh9E9Jjp6tg1gzyJTzJRlWA
ChDNtQ9Mq8i/56kbNlg/7P/X7bfnzXSKFzuLLOutTLPxsB3YMrQmYLtEsT+piAZK
m8Cl/WN0O4+7yRo8TaSaPh47R/dsN0t70Lqz6w2bQLnxkBMuQTlMUf+7nvaa/A4Z
Difi5YOh8lxa1M4AibeLj/KN5pGMbMiZMAKzZTsYwBSCizlVqKTlok7/SVuDMxFG
ViiKWZTvMucFip9hu5xYVeHSedYCwnBgeZRKC1+ocxNgscB114uNbTS+i//z5Zz1
NR2cXbSD68p37jUVaDVY2lihpU0fb6KwUmbsIU0yXCRmIa6cS3MBphXMurhcfjP1
n+dqKuDn9nFTh17c/yNVBi+mihxRhGCZNyGjTJjHrH/pBHPTNoZrRfClIekZwf7N
4crbyQgoMewSJjClG9Xm/MF8CXSrm3w7EYW2sYK2I4911JAiCh2cp6RYbyTjEYTa
Q0lPTEB6T6fqYyqF9oV5YbR6Cb6QDtb5jBJhM9/xOE3etXAMgveQ5A2oiyyECQdY
0sZhoWz974fJLg1hrljfQ0v/JWuNY1Np1x/RYabwK5HxT2qwiMlGeNX1io+1Yx8Y
jjfrc+rm24cO1rpqae6ryLKMA36OjP+/N3uOH193GAi5Oh84s3QJ4dM1AA1HJq8H
DM6hH4OOv1uWOib/zAWGuYSlt+sVvwNZqxe0s3iXUqEO0A5PZUsiGLAUkNSo6gi7
B+yYey0JvswGUouL+GlXXp6YwH89LdrvsAjKxqiloBudj42Elgw8vD6ox4jKMHaI
Jlkp1v3ZraIfBkB4zPjle2J7P2Gl4rzzqtWxov4majRd6JgW9wUvLBr5MAdKWC1q
9gRwr4b4eEyOH906kGhmJc7YO//gRrl+TYAv9offFwF3wwIyOngXUSlAlFTnMUfV
4CmV0BqccFMmcZ5DTYDzNml4gLPEPyGnElX0l6YQA0QB423NN8oHanVp1OKjuZNt
GoBagmPxWmzNtI23vJ60gdRwDhfcTb9tfr3X+OtMEyJPx0qU2uFUcMfTryUVgLe0
v2Zd8PNDmWwMha90+kBoNIUDP8aVVPU9t1EnXlCiG5xovl9i1EZr+3YzrU0sYRFg
MwbCsRTUp4eRn5NCkoDqxiTIlrIRl40Tdevwp7ZCTBnlWAJpWstDAG/osBvcMsaQ
prhwbOT/0m2z3oIzrx2/jkcdlw2JNeEZn/8+s8Wb/x7bGp5JgMW6slsiB70DMm55
+h5oCqbd7ENZVS65UGdaareqtgx/DB3VLKLK+gJCGTFpw1vMgCpqc7BtL8LpmEil
tDt/KKmEq0X53CnmpcWUr5MIwUohVvuLFPEp1RT4MsMl2IsJe57U5a9DN1njia85
4+M8hXvdNrnjwT9i6oKs0n+A73MI11IfPLcSdtug3/ug790gbDTvDQV7RDtnA/p4
NHEjzBXacVbAgCswzS8jSkJLPROS+QepPOrWLTIpLvapAjkn63HG/5KFz/e+ovL3
EGsxFHb0yraDr8g6DTcYPye9OKeP8Grv4dylTZz4G4YWq44DBDUbx7bq9lBLXr+R
cLDXd2uxnOsKDLt2ENMkPX7pjwaZuDoppZs9ot7Kl7ZtUNe71GDOFPT2JjBHNPxv
fateAo9/K8C5xj1MFgUxcgENaHCs6ZNVVbNeglm0M+1G6dtdhOjzCoh4k0Q+h6Ob
RIoLFAoRBnpZ05Qg0ompNAeNIZTmYvw+IOsz5ttmZc3Uk+Hzf4ZFgUWUfx9imToC
Ok+gIf3qLjTtMgeRbtMWdXpCFuCZ31LqAXCGspxdg/EuRaCINSkgQeGo9sOs8o9H
AemhRSD+QbGLomqPkxIymvvM8R9fO6Q45PrazYJq2SS3TAwLy9dY/IWQou0bdcTm
Olc65ZIUBAIDlcceZvOLwKD1wJPGY7jDqeEmpkkqvPeLKVlMuSAvFG853r5T3LFB
bAS7xbSDeIQopIUiQUQa3KVuR+sfycRTm47s4Z2fSxt4UTORvgcGUPiUkhfQqY9j
gGM1rBaHvUcPkEk8FF8Bbs4b31XxkBm5B7BrFwcH6OBxqsEXHTxAHwbsrmy2xuhb
meMDaqd8WjxF7eJaJYgVScHkJVYIM+hYLvPEo/X89moYW7vjKCD08xvxS78kVUrX
9JbVJ8fQp/J6n6P61dcTlTP0uuciM7LSum9+O7zQbEXiqHj8ojBvtgAtl2AdWYkP
5q9HTiW/H4vq0Y+q5B9aqlaXeSf/Y9owhElvnRNDoowZIm9Q2XOvi0a1VuPMDmPF
YY34a1xDLfwf5usiqPFIaD9fWoi7RyDUS3pEslK+SyYjUvlERYi0aFVAJYwc+gLR
EtceRsxL0BbE9SRT4NrxD3+0HcNbNQ7YgVSZUqpRyqcxe6tF3Rrmj6EvGrdUVKUW
l+w51lp/Y7WWCbmDkEGqfAPWGkj4lzYzq6VofMQjKS46YbEc7lihJJAXIPA4HNzN
tyQWFM1METoCfrA7sZOuyWZHAogSQRTZAsu4Z8b+mKsftTOImxFCEOyYWc1KxdA6
GhIkiz+1mtBKjbv09M16pQX4fAMq4NFV5QqMBFYYrdanzygQkspT2zbY2eqr25iR
taQ7TNmc//0pd2ZRCsqHJTMjtUXStB97ji9KuW9c4Ss+1gFL9Nv5JFUFXucgF5tc
CgpKodcbvn9GidTf5RcZWU/gcMRc31JfUZdJod/qN+EGbD3kHVJEHhwKa1mXFZhh
oBL+gJhllEbe1gSujVk5cqe2/WC1pfQJkI/InnMU6ZtlLqR21CKf2hrV/lAqre8r
gCzDpMk8bEv9GJj2fXVhZSzus/bA3MhOuI/ewnpwrpy7purXSIMKDsJ9Kmwm05Ao
EUteu9k7yfkiSbR7bzNVaCnSN+i/BDfSSC7Jxy1lTQztG/Uk+EI9Sfag5HkGqEPa
rOAqSbUCwIicnLZraocDazwKjXISbe88GkjNSfI95Dv6uI9iyiYDvSeSv/OoQAXz
RlScqv8c3VT7cIBg3OWVq+2qfH9CkWSo/Dc5oBy5mBbysje3AAAOGtqKiFVBSeRF
8B/VMPQGaTTAtJCyM9ZpS7JvKqEGo9Ezn3hUqDr42w9G1WiddEZAr3pF4FKafEgX
rQwDdUkqAac07tC1haXxL4wa6H/oX8aW5l8K2Iv0Ac2dH6QMJyAfsnsyU8oOG6Jm
7rVZp2mtfJOz6H9GnV2woqJuWeBPYyLfm7v5wVo++Ff0vPd0ouBJoJsqLrJqWi6g
ISzA6u0qdPi79xeDbq3u2nQIW4qzwm8Xo0KLj4NCqIVsc+7vEgFZ2fV9EL3PEDj6
qm1Yzsi5iLsxYKT/UqRDlsr/10lHJWirSUPVKa0RGZbIEAzXFXJaXe0R2VhmP/lL
RXq+YM1RPDVJaJbNTqC92MvbgMveUvNDJX2FzmCsPPsupULMAy/YPtljr4747U+r
ORed9kYciSZias61NtlqsAVvfHMKJQezMncKBBiYXbgjqKL589lvdjC2Wldp3OTv
CVWgVHmAa1V8DVsOTc4BsR/Loyys5oPnvEpZkkZy4tojF9fMtWC0BYXa6qV1iFD2
mOS8GP+JNnOujJ1gpoSaqTenG7t+TvaiRXJdXahn32h1nZe/bdVu4Ru/zwXRFf7K
P1OLNLaKdZaTXeqku+uis57gDyU/Mb8J78QpRtNSuF8SkJdLZFsKl45Qi8R0m7vo
3T7Mo1fn5PchZVZo0C6RiyrqUDjrpN1TsmW3U21P+K2MwSfir2AN/CnzVZ90ImXT
AsSJwL/85u/mm7ArbFJtCSV9OlJwWS42psqN8dHTDvxh8/0qgqV3phT3Ohxo+uCL
xQiaLe7T96vJUGulLVtmqsnrDI/UqulfEuRpcWJTCHJknnjOv9p8WqouQpqf+qI2
S6Z1AokzZjKUueIlx2PzE3yJ9MGQ/n8ySwY1s3+aiLjcVGkCO+5F68EMmObbIfk3
cUZ+5qJy47ntotSbF+odVXMSeFa+WygfPJygyKie3Qb44X2Yqk5BF6agzrbhIP2N
XS4yzK6dE4cUFhKvPiommysCz0EVjQRL12warwh1WJlEEj3y7FuyxO9x67ZsGtr8
y8yepPsVw+COPaJbZSFo8RbH6HoXU9szeE9p2GYf077SzzN05pFL2Pw8C2VIqr+i
lJaYIF/ojNHuX+iup9kKrLnCLylKzU4I6T5JcwbscFvtYuGF0Merf5EpDWh41KO7
t2DgYEwqwHAkb1mOikXMd6QOZ2K9J927v0F/1M2wYnUiTV9cWBCmh8RnFTvmu1/1
EpfimvD1E0d4TEIbQIH0PYymRonisPgToOzi76DRZ0NUSNegf1B59qMPRQMpUDof
SxV3GssGXeZxfEUKif2NAj7YnzOuBYht1D1Xu6b2QDqYsnHVzgRE9zQsV1im9YpB
QdxTdcjqip7CzihBL8yXDyXcPSZobOv5LN/ciuDeoKOtpHmm29LvHk5cGOwZx/6/
WgdJkc89rhS9rRHFFrGbaAwzSzHZz/ONbpKrSqWQyBIAhCBrVedw2hHRQ3cEnhv/
dtNDoWYmK0sSR0aqpVC0BqA+8akFKOxp556056G3oJ4Xa2GDo5OaJv+1WjXKwp3V
QsJLXd4bVsMQRdnAuy1XEY7VAXSVilvVugpjPzfh64GnMo7zlgQUi+hQmIVkXTiq
w5Hf7z2Vy2Er8HzI1vFqMyIz+VfkwE43UjDQQ2Nrh8/G4Pk5kP/v3xU1PyvU9ZqI
aWB2Ly64LppDOT+UonkpDpwIxbzCegY882khBsWVVNF9HesYhSA2wCs9UhzLOwXR
Mm9qpwyPJS+0pFjaln65S+/Ax67YihI/zMMnT1X48FH759oCW4/5sz+U2bAlpelw
fXE8jAGPfRwmbx4XylTHO1syxVEdnSDZcxiCX+pbDOSibT4Nr8ni02EZ/kNFQjPR
zNSSLyMtN9RNQe6vwJT7dK8IoVeG3dmcnl+DY/EsV6eREq1OI2jWm/rvoOXFHrI1
+ItOAewixupwIeibWPVbvZdR9puEGG/v8DSIcLYjc6MY9O/5viLewIuUObEwM4fj
9XqrAeHlUfRoPePXDMXL6dhm4l5DCxLoZ39x89YcOrZW/lHc3LiiHOlXtXqqHFCL
RNB7HYBn3Tga9h8RHLj+6o74H1HNTLAh77mJNOGsqSzK1cZgN/UKfuBEyS2fB2z9
fS7/NKhGSjnBUj8srk6IzYqNY6O3rsO7WXJl24rih+rTzwas5aHGv3KHTynBbn9K
/4bJrqlPawERplImtPKmP/LrEjueDZ7pRtoFSd8zGyJu4I/iHWwcgoXZqnBmdvjc
3lugHzegnaOisPSFEQQMZrDydX6BGsTAe0xR7jxZ73//SVTmXyRbZ+gxiSgMuevo
lsSy2eKi9/oeARjQO1YyEp68Ul6wFejygY3Bo0f6GUQDCIj2Ef8BoNjtWcjL+KhV
5i6Ok39vd0Be1jqDpuLSvEdHzewF1vujEBu6+DNDuO+jV3UnU8NOh3AUWbrRam1l
hV9GjHj8Sv1nHA/XoXImrJt7Tl4yvolPHjFOlRJtB/gdSVJDCLnpbtIa2a32GMX2
n34G/x72JUye+2OxAD6X/uf7d8eCTrwxnrwM8Y9CDilTIhLIC4zmTqCVRKD09ROM
R2d+GKv1Zrp5VqYqHr+LsTR8OdTT9y2PVk2308FQnd2W30a0ToWiDR50v+ZCFIIm
7lcNkS6WlyGdnHHs7sow0vkRXGsbLw1N6EBw3d9hsMmimbTKEoKNogajrG4jWWBC
YGBJg0coBz30Q6Sv44Gk4PgrBWVVx9QR8tPN98138Gbfn/pBmlrT920+m2XTc77H
YVQIrxOX1DqvLa94bjqORx2KJBW8Tu3SLqJDc8IeXeo2lwIg4OU9T+XNkb1Ki68A
8Z3/ruw3//FphLXqVtc7BA2fcbKzRbMJg+UZEt/fs4H1c34eIjyvvlAYJQ7O5mpo
n/tF0IPzouBtoadrDRy2I032kjJy2xmcAEjW36qZr6mrcn5NaUZ2qjBIQjaf8rkx
dkgbwJwBXzhLsQ9LMD6UmIt9pMb/yS2u/UL2pIkTVZDUSn4KrnjlZ3tG9BHYQfai
kUxPzWqNbQ5660VU37nbDJ4Ns4BZcjYfOPcjX381wwq2Aw826yHxfPH5Yc3+cC0T
7d7R8xVgLcggIK9HyXjaXRu2nOlwaBSoF1UIBAw7i/h7NnFgVN55Xz4ktTtWLqxp
bK5WJyw49e5bH/p4NYQyiwS/jSiyYYBtzqcFqtiGDVPgxVcoeY07i7GgVREq6b9A
0Oj8ZsaKQb3AErwG62DdZOHeKK6wXqmo4xX+M64MDWEUqqHokzz/5LYTIJZ6/KLo
aB5lYtdSOginMoQU/fhGNnVEztk6D+XAdknYtvsKMmsdOllQGnW6F1sbnXWIT10n
NQSqq2ySEwT23iMr3u9s7T0SlzirPkvNjpJclQOm5fpCJMF6d7jsY2kzugZu800c
ToCr9DqGqhRPgjHplHg5zPckmrzF/DHPqIdtyGET/9K5fsINFSyWR1/uF5Zurpli
uGiMZ3NP7HeOvPMIyxGEdNctDkSRy7edXRdq35C2YdwpVgMC0nRT/b2Sy83yzC1A
i73O+oLR0LS1VsKFG29NsYayBFrZyn+qYaoximtj5EDJr0njwDpblNWWu/9cXNRN
7//aYrlmWHbsADHgapYMZoJJvECpvCVW0MZ0NfSBjJzR2KAkipyvbwpvf/l3NOOM
NziX7brk4BWnYncyODWQaHaZvbP3rN/pSETp3RE/RH1BhXaI1G2IU/h/UpPpmg1A
qKgWUujVN+FkrBP4bfWblJCQMMszFW9sst15mgVPNHUQv06817KQ8XCa7eWz7JJX
EASXTuOlwJmHNny+ZPHjQ6MXY4mkVTNIYa5W4Rov33ydkScbqN1VUvCLxa/0f5vc
Z7mnzGTcMIBH8xDNgee+QrTyU8tRFKgfTrK0tg+hzLwfYItBOdpHHxyCV1aYMoQz
v3/UsJHbuO3todaBzImCRaEjQ+iV0t8TrvZo5G1L2NL6H56vJgCA86SL5mUCXuho
2LNs186cYLofiLenqihloHB+qwCFueXq8/l7cWeOoZL462rVWbB0dO3Q9VJ9+psj
RafcYn4BJSwmWNfAD6J2yYenMO8QYv2GdeAfTT3FuyG2XbwtpV8Kd2ADrB0QiPOV
GhkUs4lOytGVHjOe6Waqd579S4IRaLrea4WEYbHXVxAAGUW+CirYiOw1Sgz2W3T2
dOwGzsB8CUgcqSFh+tIceZgIdL6RQdizCgs0+TWpS/ojHS7gdB1wh4dPXK0Aw27j
kCp4jUYsWYE+wM16cZGSRW5CUJY5OFcq3mFmstZYnGRDQVoxHyCuWiUpaKczPaJn
+p/OfvRACdukxqZ30kPUdGmTHS+VIxAc1Y0wzlUCdpsbqQqIyZda4pkAe2gIJK3d
OUjdqwgn8pjWvTJXAOZl4txmNxjVJ5ZkEE0F2PwFu6a4pVRK1v9cY9FIXTJLNTAZ
Vb4sdBz3piAC/wZUK+an71U62RODH6pWXueyCNK7cmkZ86jc0CKiHsPZsXsZc1D+
1dELy/b0gR0Chnm0g60Ca62eQeVUD7vu6kVWabloaTGtE58OYpRPvr8ZLs6lq/SW
pQVPfm5+XnPU3dpOSHBYyMvA1RxkUvIr5GF6I3oPA7jBJzwu+PYlkYHOc5qLlwHq
53zBe5c0E0vkeqgfLQr4igbdcQlmQ5eGAuaC98BPILhO0oEUmHFwyPAIE4ySzjjN
TteqOlM2QQe/xvj9vLBeddkeoBEo3Zn9MTEh1Mjogcu0ov0iM0bn652Kq9zIu5D1
0ysTFDMeTHTuNymNHDgRf+j08BxXC2zpq6hK44l9eOL9ws7b3bNBTXy+LkhvwmU4
F6hptY9hvl+nmwN+VArjm3O0M666J6zhwNbcRpnK4lVZj9qm6At1TZBMiZBX3+Oa
Pko5xQ+OgVNYykRe7LRqQSpKKzj6O4r00EDOrVOJX9/BWKDLuVsrCol0PMq7yQ1Z
pfrwx7vBl2fHcjqs7fKJyjwhCs0hb37qtOLJvnOIasUapYUumRAKTNCLBo/nDCP7
IJVJWMQmqBnhwV7AfUxldeIZYq3WKEGrhXyBzVU6lY91QH7C54TaIDRJGXCgM6Kl
EbxLdvvr7f4AkaP4Bt08Y+Bvy5LSlQPRFTixpCXIK1M+etkG3/XO4dqpTdsLYGVJ
mAoMsTZu/0vkLkQ9q25Qvk6oqrw25eoP6X8WkARZAAobaaiIzesKTE3ln0ey1ar4
K0cVhgfXy3XUqTjF3rDuib6S6pXTX6mQMdp05rMZcyuxM22O1XqpDxadpBi0EFnS
FKAg/MEnIkJv6Q0F4u7DMMNK484AhcjHUqtVym8Sc9xHHYswGg4N2iaIdAAdeBdt
ZEIRTDT8XGC8Kv9nzQ/RF1LDxuBCophP6xdhJuYcG1LevNRsjVYzxw+QFULqJBZM
/eo69H2dOee+FwIjaX44Ue/uEjfHhkuKWIG1QnPzE1XiQYjh8JbTWQxJpQpMYVZG
I2Smk2Y1ACa3br2PcxwTy4f0sgNOMYYubv/nj3qwSSzrvCxsi4Ii7JMwpvvmc2BI
YjjDB0R9vTO+Px4ErHHxm0jU1uut+HuMjPhZtAHyIJYXrI+SJcdtm/UFdY/gRbyg
0TogR7DtJ4eLbaT9dGR7tW1l6kKusnRSk/4iJEsainy+YJCq6f5SagwBQZ+gFw+m
KC6WVJbtLswvXL52tcTJb24Qez7NYVnwyaZxEYwDRG3eC7hoV7mGLl5Busz9B98S
OXkonIIIQ3n1jgivKPckdQ2tUJ2H4sNjwivvuMM1yXeLawPQoBhR0SrYpsXN13ER
7cbcLn9DbHkaFsQu00Em10LfUORzwf3adzfBLeZhTCxDO2P/fx8LZH+PKUADvn1X
QofLHopQGR6dao48uK89ZHcCxINdauZ2SDv3p9lG5fBrMxypLkWnlE2oQfwGwoLd
qzShQeADM7lDMaUsMAVZs9RGO6bWYMHoWWbrle8iYLwT/lQ/nRscrYnE4iLcrRqs
XhoPNaiN1oznEGnQOWma7Kp5zPkgH7lNqWHmolGaMsvznx3JBCjLdaLOYb1UFhsy
9+fm6JqvjzbMJDrY8wzM+ow/l46E6q3Dy0E7szWxtCGNvJzDJq23ldIEMNXL/OJi
TmNs2f4L7i4l9G8+A53cAEpOppWohdWT3YqRihH2cqQeQIh/n6J1NEm2ubgTD2vJ
9vM98xsf+O6K/RWB9Nbd0a+2rlYpgQXml808iN6EwhIP83tvlvbM3j+g0C39xHPD
A2Z4bntWp37Mc8g3NkQAQLfUtoES2dcOjzVVuCq7Rpc6mXhRbQYoH/Bi8wsDv/AF
rXWfSLu+UKRrkLZ0lDgXW8k3MhiB1hRTZXgyJxegdK42cBdJN/ubzPd58ezfNd4m
c9e+V9MNfCM3ZS6m+nLXVDO/aknZTM1uJD4f6chwrMbuNVLooFRSCLmyV+EFruu6
QwSddbJVI6Epl2mWbpi8FkX4NzJfSpycHlGpEXMtYDe9mlECnb7M30bgZvgFMXBo
hnbvfy2Vlzw5cjJ3D+KfTNoDCp17sOHk11QNfGGb39lub0lYy4R3CiXZNhgXjkSl
tupA3lPQsGDmMPMtYhUXevKc+STFW2Q5t0LBqBRbtHqPuWa9jiZf5WtJ2S0aR+RQ
ugF8NMGopP7+f2tbxsPKyr8QdHRpm/ETCDBCVEfT8G8vSwM8bCkO5tlamcATpptb
TAaskvNVlgmniq0lyukGh7+PclaTG/NyMrcK1qyPtwupzDa6a1P1QeoY950tOBWn
J5Si4NPZSxSG049+Ex1Kvn3Bu//K6KM9GZ0k/kwlqwoIZPyoU/143Dk/5iYW5LUQ
gpy5B5mmsmWP5JURT/ILzu4bgybyY5WIix7T73mYRsUe9np6F6wuttBFPZdIIyJt
9ZjHlBep3KsRtFAYF5ZNXDCMcPAj1DgAxK9QR9UFNNyhw8r3efVudu1xX54sZ0+K
ssd6ae9bRtlXmEpcK12qy2l+qEYhBWSgbJhHmIITMOy0JR4v4cwIA/Ycrrs9OpPn
UPxM0lHlrKZd/ZSksKKWBL+2OXUwpr+wCzRdPm+OWKVBHbckjEj70Wo9rmuznbnT
fTmiVvt7uVHpCZUnFwkSEBcyCb7zlGTHGjtZtUodzvPCH4iKNKdhMSsGQiYhUtsw
BXxkmyAuwU8yaCiyoJc6ybbpCVmx/kHy9lo0o/PsGKtpswLKsDnzDwl6tARLtC2e
YeKvm71UmhfjAuKQggH5uz+IQBRBi7IcxnWVhfiAIpB5TlDpGSImLp3qwLO8Ks/o
RiVnosMTa6pprhJG+eAJMtTisLifnfHB096dHXp717e/gTL4C7atWAPkvZiW9osb
O18yEPwybbQERL9B8fvfw8KMNj3zOa7c0FDtskMa2NIxtR0x8ARGIs32WwPY56AR
EoXkLViXQ41azc6sWX6QEeb16phaPMBsvCLO4pATer8lXd7cO/NCht/XvXsK6iVe
74XFd2IHzRCcZ8VCX8RJ+2swbwbVDNBB/76WzIj3bPFx09eV86e+wpzPmhvTs8sJ
+RtkWYLzja6BdO/tCPxZrOZwjoQxgI9etTb4l0XXQ3iCUWR5oxRQ5OJlAJrntMho
wqkVF5qITlLzyWcjVtiGHpztIZwL1jNhKjLAUqzaVpKT/Nsj2MkZr3AfpGF3Uy9w
b43qhZ38Ka9vMlM3rRBsQpmog8axpgYUyrcEqhtCDd7ZzcC1JzLxHNivg9FKXiv0
OdzkQKpOKMHX7n7OicO7dMfQUSA+n+cx0t95PhVaMJxKmrCVHyJZTLFsiFusIAH7
xYXnc8M/ly2Jj4zim96NOHVGiTFycirXiACS2TtiH0T75sisafjCtbvKLzlAZOgL
bp1q3NLzvS9pISkpA1hXAU3LgiRNpmskud8gNNVItzyZBfEicY27OAaHpp5moAFb
HFpyV/E9+mM0uRvxVUwIassZGRpcjaxmVxJSSc+6+OsCVFLOtyBY643g7jfrDrrf
jPLEg+TdTp1w+InPgJsyNRvl9K3utYt4zwQeiu7KtOsa3quaWTityTmld4109mJo
DMeJ1bxd4SUD10HCnPDZo1yo1QK7bsG+BbcmTwAG+C0=
--pragma protect end_data_block
--pragma protect digest_block
WCKB5b8Dh5uvoNP9qGoClhb9ILw=
--pragma protect end_digest_block
--pragma protect end_protected
