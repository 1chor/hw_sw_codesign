-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
J1VfXjK9Oz/YxWw690wBBFtHkF4+iR936217yyHv8KW1Rq42VNsY496xKAA/p4dP
Exo/yLcsAgGRcUSwvkGI0xqY0vEZ6Iq1Q1frmktZjfxZ0L8+f1pfvZLAbNUExfro
xNbLnzmoZyP6DvUekV82lpyopn2MDziTp+pj3xgILRh652g0XCWq2Q==
--pragma protect end_key_block
--pragma protect digest_block
gS0O8a5x1pv1nmMtwl4ChH2P/+U=
--pragma protect end_digest_block
--pragma protect data_block
p/AvrsvMx+qNw65UbaHZMbdqenSjOzjelg4mKU4pj0/pztFOffKuA506QcQlvbsF
V4316i2ob9FMsg92FK/U8F3s7H92gvP7ZEj6HNjM593xiC7qJO4e55itjfe2Rlo3
VQBMc1ZicEqCO/q2f6IGtdKvZmMC+sWhJWsxovstF0nfhO2BfBxpG1iqqYDTvpJs
dkV0USOtItfyW9aox3C6SEbplhvkA3e5aKBth0XtmELRY10Z6ySm/Viw6NgjWhJd
k1mcJUgjuEuiMUrla9n2aDY44QSoHBJ6Z0AkPBp/jhK4utv16RnEOtAK8OVFfbOP
C0VhsiTo6EPO9z2vZaL0/0wUrGi7NA5Bb7j5xLzuV+8qFeeAg4qKyvQqS0bYm4fx
Qab6hi12SRgsQe8Jrv5aPqsAOw8XAvHYAKEHj8qUYbM8nk+glewin7yRjBtTLEWR
T1Yk7gk3NiruQImlrrpWLoztL6I8XIWIvRJdGKlwqK8BROC5RG3hjZDXa3Ai3b7Z
Q8SgmQ5arACrLkIpLJiCUYqbCBzlTDbfWtUgZDZ1QGDU9EqNh0NjodQbRUaYC9Vf
TsKWuDtc9oyYk18eyw1uDoQpAYYgv4ehpO0VxuU2hoxUYbpf3AjvCKgZYz1+kylc
W3oswMiE0Ouxp07og2o8UOkaf7q+waRrSVUljwwUtd/N4C091djoSwONpk4v8Y/+
SxQDvdYqt7Oz+pDbABem827jHTRrP+otXiWiDh5O80BVhK+rzBTdaPEvEyqaj69E
/fOJFOSnha6zCB+/CbfugdypGxzv0H5w7x5OYqsGcS5mWQGWJHLiLj4fz8WSczK3
nfX9KShIuj9OGWnoCe1uqUNh/0r0UWnZCsxgY0rTikdGiL8qWJYZMyg08vHU7dHF
o6obI/5f0wdmJewExbuws0jjqX9mgiy5/UT3Mi7r9OAhJPJf3XCL7pQQVxG9fsRM
HdSrROnRp9jiv8VazMEtDDVhld74k02T+Ifdho8DGwdeTuWupvYjUvPW2ICHjs3H
YvU8zR8EmuPKt8OeVtzOgyt8H8+/o3P2dcgBSWZyaToAe9IyygT/bEA8q5gME1PO
HUC9aLgsOU3hJASgsRT0ClnTA+m7egF0/gif1Dz2kEgEw4wa5nYu9+q9TgE2qC+y
OKY4nudjkEVuFwirIKxIPReJV5pR2Bi4K0N5GWyDRz0KjwBljNKj1ONFmDu4holu
9Okbasm5Jbowgu9Lncro7qX62B0A7W5t0MZWNJ3roKXUZJlCXu3dPYm99+1cazMm
SykkebgHz5VxYLIEchUpEt2MXmR/TBApOPal1fzLbbUu/RdqOKQZYnmVJ3T5aEcs
37m3ViDcuduzHQDF9PXgRiAurlHyXMwLAqUGaWtR8u6mP4WBvEydoooNe9CWphS9
uFFUraao0d+ZiZeLpC92VsTzbfR6ya7N3F+LDv4EIstiyvwpTly5pMSPFFCrEFyu
WOf3sfu/sioHunWuR367k4naUpY3rGdB2o62DrLIuA2IrmgrRM/XCEkYe+Aa8KNw
8wGy5r2yIxyrMBKQ0Olw954+txdl9I/oOxVF0wRIwca7D9hf5V/BQquoBl0jbfSv
/BUVnoNKCEV3qsDpj7vMmIMobSqNcZT9aKU+W3f21a304ooqHvChYvCr7kdAjeTT
nWfIGzZ6FZFvfqSAQIE1eQSa44ezA1woN2RWwvTiQ7Ydo+qQ+nyXgmypaavE7a5Q
z8nRBvAPqDY90oyA0PZK0bS+TyXtM4mFET6HN++aZ5P6WJg3KXw4gTu9VZxNkbKz
i93mzuU7ueKwpBj63hESlCbSGifBtsloeM2Ikb2uT4BfnBHJNv/8cB/un57Jac55
ie9yCNpxpj72kfaxn7fB4VoThIIkcofM3eCE05DO8RrsUp79heSpR/BTHzntPSCN
fc89kLSQ6OcYd8jnofBrfAymIWRTIWJTBjmBO7hUcktXygpSokChLgf9I9rxHXdS
Ek0vjC9/E/VW6/jOiGAu7obbKFagX7vw0bulEh/bRCFvCR0Clmtt/5WGiNEsusMV
y6KP3hYtDktpVwHzM2HTVocRRHrL+d3+lXfuTb2ihofb9CJfBVK8wdiFIyJL0S+R
uBlzXLao2KSYyouemObtHIJvWZhV/8JEjNTKSE9+Mvuz4i1cTEZ2s4EoT2MA0MiV
KxPEqLDrtOzuisdq7OF9wv2h+IYcm2m6EPiAsE5IkkagzS5UoJxWeDxPPWBBA89f
spH3qZwA48WE5pY1VDIvg61+vzds4vJdkPxwODZ2GBe1DkNvSBVzRbc0uVge9lfW
9fBbX/kmBbCTDq95ENbYxHnzlvw3JMr+3We48cSAREU45j3sCuxna2ok99sCUHqU
2+5R0K4J613f2Tc432NIsEAFCbKSrPuhsRDrXMn724jyLsGkMxBMLlbxtTL2ifBi
5GYdD2G1PkuBTuiKtCq9RoJytnNgvdOGtoANfnyW3/CTwDioDy66rmprgDlwKdRP
mwEBCb26hA02qiRdTmnVL/8UyURZA+RKxMPMKyxEg3i6qosevabjDO6XxIf2lkl3
82DG6mAQ6QPdly6oUSW5Gp8gkva6gCDLjo9mnYdcBOGDqnhrg90yIC0jt5Fbybfy
g+bPatI/pCCn+sKMdqYUO/vnt6Wj0jXtCA82WjDYj1glhqYeuE6VhoN01N6IuoJw
DWchhSZi+D1/F4w21yNBETtHpdnCu+ZCp3zMAou+t/NKoP8xeZR9kO/LQ3b8H4vk
lcSyKnByyeoXiQfnVlaLTx1FyA8QQPViNR7yhemZQh0oRBuvWlsiVTbVX79Rke8b
rcDkQCv6ROfhcFu8N0d6XZeuKIGODJN8fpRZfuILnIj6jYpNGQHdNja83XglHTPb
P92Z6bsGyHm4UNxZl4JC8WYjBiqZTs9+25sVfYY+NuQyKSVghcmjhNzWJT0mkFjM
5MxC23o88H7PMHjNVHLL+MedtfaKdECfNzHYv2habR7Bf7l0b1XZTpxFzgC/60CU
oDZT9ol0Z50+EhdzfmZo8rQYW4rXxn3ALicYH/i2Mns7S/2njTW62Rh3TQ+cC771
qvV9YuvheygE47y2s9TTnIcBBaQWECUHVVvLg4O+ouayGx0S05W+m6XYvj+rv2rT
O3jyLWBdNG/AcmafAsaRfcb18MS7zkW8dW+VbKw9dssHvnrGd3P1yoLo71BiPUtA
qHrutGuV0lS013aMnp8J59/OZ/ARQSk2KLXA73E2upw7Su9fE9ma4PkmlQI7A+4a
hRcf4inxVYhhQwbmCbF5WZixVikdGp+1FKRqU+31AMshZ2lT3wZ0bcMc/5dLwex0
uWHAk8WMYKMHU+CU1veUs+fjAnFa8/mR80lqiP/T7gyCnxoMDmVDnk19ku++NAds
3NxEngv99261c2ZAvU+iBAI/fCVzsSYuOxquz+yX9l1g6fSRWiYcvthEL5c1iKMs
qdnw875dOgIiHOp5P77aU44W52i2VBRwSGrKrteJ2E+qooQ3387xpOBSDy5b1VE8
Xz/n1M+gHKaO1ssg5Nc2qJd0kbnCA6+xgMHzehAhpbLQS/8O9mwDxSzj7OZG8S3l
j4ChjSUyIMw+Ik/2y8QbSvOGxFN8RyXNe7H9lAaCCwhVZ0mzusR7DkiLPc/fSaae
4jjnPR4x10m8KR9a09LoyVdzX22HD5B13Vk1skR3sHUw17bxrfuuHuvmmRHERn33
siKmzH8ecPefBsyy2Ag3HU4LjEmlXhzMOyxpfKwpKS++uutVriW44cXTid/o/BqJ
XbF1b7lY2NVajyqJUoUYtcZfQDwHi24csA8rvSC6eE/F1p0+U6/hufBnhFel1z7s
x3x2bKTl6gJSlwY7HHQUDQwH+2h2p3rh3rxvHAbj8h5MNb0bKg1u9SaTJJ+84YQ6
2vEhANG3ZuNdYgFcSLoU53PSFsxR9N+SPMXJK5451o61N9ObCIggSpQbBKI2Equv
CoN5pag3a6HuNiKKpGWNtuJWAPCU0RSONTIJZ2oapC02/IZRtgP7Cp+HQCMn6z8S
crKIac+w4IZTnR6CTT5Fq8exvuIxFd7pUZa8fyz2EoYJ/XNet23usTkKAo19Is4A
DSRXWT1xbkk2x2yAWcjxmnejFsTslM4oX1UmiH1tuDrXCHQITqtFdqrBWQIkvKnW
W0bp19p5Y8IFF7CUFNiDbyqm/Vw4kbKakjJ6q2fD0PmLfQGZDHI84IauZ4ECkvyk
vBjGSWOQzrwgeh2pxE7G7tfcohbvXMfHfzsFjxQP05wWGIom8vvO8/czk6f+t0Cu
3Wj9sDC0ZmGb/8ZXv/jIAgdeJgKk40ZGCk1SHH/zQKxpLbInCZC/Qs4C7VB8BVS0
3TD6ZmfB7ggsntD114I+ocEuBB8PPimWL5l9TRWKY1Cych7E/jipVBsQ3W6oAgPh
jY0HClYex/mL6GQ36LXGmmsaUJIOKmIFAJSOkir5u8pzynUrbjtBY335+DIGInG4
ZUDRlnFC53K5G36p7GAJftKS97/r7/1x7IQpkIus5H+mvkqf4TY5KqeoqNKBTuIo
chqngFOmD6Iri2HRCHaYHXKBmbwamRj0pc4HXg0BAw4sLAHEIegxwsAz44jzm23M
Ncoceh9CGZhMxswi6D4J70d1eUwOz3OBURnLdY3pYCfykDjf0JEAf7Vmb45s6qvR
Z0I85XuS+VE4xffAxsPCPUQkWH6sxYtEveVuzhRfC0VBW7Ba6DgyBVuOK+g2AFr4
0sQr3NYEBlNRQripVVVwIc/zTRHiNk+jTrUNBk3HGWDbTDLsauR8V14qZyVL81ny
weS/RoZOokB4oT3QwtRiMKB7oP7PsV/Ug1E6MkDlEF7tEEhu0rZT1YbR8yAwe6qL
eDc6g4k1whhGQ6BDYVxHlBwTb+JQcvFyGoNyuTjVNyWn6FUX0oRx6SeAUFH3JUFc
W2Iu2CIU5t2fAgdez/G05VXiu3RTtmWDHMou3gyj6sAZx9YeUNpsE7+lo7o6RHVS
/q/aP7CTwrlCCmcuEQFQdYAS8tUsZzHNqKaXwdvN5XgAfE79bB0YQ/7xFYYaKS5c
ULUughb1HE6bbX5GyCT+WKpiIW59BgVDXwjX+tNqKUVSgQhELp6XUEOcYJ3/bVLk
vogQ6P2CrKFBP9we5g6X09mSjN1lNTOFv/Z0bWkvjK0tQdNAYiiDztSCAn9BoNa7
P6XoZFO2Xtt3328jpL100YLwonBM+8nU76Dvb1/VBLKu+5CuEBmWpeuSRDE2bF3j
Agj8FMQ8aaQdsbsVI7XQWGv0n/0DBFzOy6H1GjiiqIu82zr1GjbeCnoWr+CoXmvn
qa+E97aBmJubCiwiTbBKeC2AjnTqDp+KGrtFIkrQdqz9erjMNSW5i4cu2JcrAKp3
KVL8ffCOEwEd5VNtKeLIsWBuu2Vg6WGkHQqJL8ydTqs/mzbTMQRWwVtI4fygoV88
2meVklwajrTPZnIXDdYset4I0CY4vsyD6Mmgp5lL73WfYT5Vdn2qotoZcrw7TtzG
CA/zRw/jYv9go2VthM731othzSRK9ZnviWdJKt0NtECBd9tDur2WqkoEAaAP1dcR
YIneRovKuxnkfTEPt8MAQBJhsc6GOTWWu/boWn9CBsIMJ4/cbXpCxrNyuhhjH4mp
X7MD8F/oLgdYzz3TRviygQwh4JS3dEuk0ZqOj3sBvjiuvth7TKjFo3zaLz83TphC
cNIg1FAgh0kvnWzM5fmVmQN4KdmclI4oNQYD02GJhwPbfCMc3twr+kzdCbEWvuM7
vNFrLrxqP9/zkHg2qzeh5VCLiWUDumci4A6ZfSnQlukNDqvDL+9Qqcfb5xWqvDfY
idJPR/XVEpyNjtr496mR+8wJzN2SdUxfaWgqqQNocI/4xxXehdcL1HjCpbkQRJWe
VK5f1+IkQMeBzIasGHJMYlMOxWZVcKM6e1hezliDeniU4FkyW3sK5jvXiVXcz92/
nxTfcfD8bHVGbaYVhjHCOH7jnoIw9nnhhKHyJlG/cviK1fxVrKwyx8vWQKj5Gou2
E2QP/AEH+xqsXkltNna/vje032+CoM2J/nZ9vAHb7LDk+Ytfvuv0H3XM/ROTDKrU
BWdlVuYAWHUZsQ/zNwZgRz0ehPMX1fs4/JQeIdaJbKWwrDskQdfzvePWj48aYwe6
w5xcfF2SCAhDTFNXsO/sFhQokRnbPoroNOxiCbp4cC1+RNzHvA6NfGwa607jPT+E
Tboz5P+3NvRQouFsh5wgUp4d2wwLBCtlp3sdy84rkmtwldCjWp/B7EQfhHjsdJg7
kBnbhqzK+Dw7kDbaAtOKU6Lcv7iPA4mCCMIxCd5plvwGWaaYzIlfaTpConmeSgd+
Q0ptFfi1eAvsU4gv7b6V8mISsGfqbF2dOGag5N3Xy5Pyf/a23NI+siCTcRnL8KuO
LUbN77ARtN1slZzsz4xk5QgZRbHdcKBFXZjDmp5EPPjXGnL39g1nGSa8C1W//qJy
D9koV9Uut+9qq2+yfOJBKzr52P8YbH7HP1KFrsUQKR86OPxKJiY8dHJP2QffEOz/
x9+FgvQQOBy6JzX7ssp6oqt/04zcYn05ZdZIUzyxVnvPuRV2pYdLSpEUaqpkiizZ
h4Yf5ligh5UGsLLFoAhg4/xtFjVXNb6TEtq3caBh1lg25nPe7D6dAl3Ordp3nmYB
GF72J32e7rBBVJ3neynFUYCgveG1k2TTbsMPiInsjQkeSwhmsnZuJBdfooFqIwV5
iE2CVRe9Srr6wfhATK+7q8RTMIOqLigU8wv4x8S+2FMxz7mKQO4vQ/kFlE+eosz0
FjLvy+1nC2P+vp3ksE/6fYd7NxJRw96un+wUqcnePrqBYhPhSX5KdaosrMl6adAi
7gSFsL9B2E9zWzDmnvswkgKvDtmC88WXfoJGMH7MUcxI7ot2Iy+r1VP8WDqaUsdF
WX6fzCEJTw/WhALbzwThys1nmXqFMBHrS4f5xNqVBLmr0/tKT4Bm+1+h9SLAyDdn
7Qi90sxCp37gFtSIE9SZk5AX3jQ0o1k4GzebInxFXc0CF15+rwIapxm5I1OJeqUS
lEZb7BNebxRVdod2kCIAtLdkJX4rWOi1WcDwNikektchLqH/k6KrNzWp26dOdgYR
UamGO6lqh473aueQOFz6kaCC9A3gzIcBYLBKXlt9KI1BEn34M6cUrHieiHA0S/SU
NNi8kDV72KEFK3RG+kUsUxHL1Gx1UcPFI03NialsuWzOrEIZJKemCpg5n7t3FvCU
QHfUXxdF/TQjTV4bxhYbbVhBBDfBnhEcfOdvg9o5wgwjxe5+T+4ulUYAfr3YwOBV
B/xfMDAuMI+VSHo/EAwALvZUEx24JdKcuCwTaI2LFhAmnIZJBXwTpzATQobG6WRc
CzV8XkrijwdX3iXlnGwYvPDJsbyniXpTDZD/N2eSq9feIJmNzitQ5TFRf8MbdYXl
ba6OIfM3efarwAMjgV0FgNGIoCRrURaRNavuq9YL0ELlH+s6sXlGpWULf+RbEBod
SqAZT1XuaSuUoC1VCmMv6cEEgmHBaBEyObz583fhSvpNSukQkhpT4tUfgsF3lcm0
6dipUvXOkAKlnAC4iXKkIX/gnIgavjtj4HL5PB+UADAz/lnQ97tKkG3/KCDgMudv
dDszA+bbgzjBPZ4msNZqGVfiKCKmXegOZDKhjERcCOz2RNifBFmE8Q+fjNz+7UZL
c/ysWg5d5Uzg72VG2xPYh5kbZG6OHxbzOr5ZgZn/YbgHX2NOK6dkken/ew2p0+nN
C/WBPOCyoWpHemxaGDyHvJJEn3GnP+HcoU3/Bz5LDeO9SHtW/k6Hw4oJrykfWpAo
ecaXvGYYMMz30xVFaL0YbAfmpt6zbAb3ZxJm5RGj/bOiFJGufeJ9Wyq5EvifUki3
pWLVGEQSYlMlk0bUltFHG6h7rCJDygLaGNYPQtaDCpiq8vu7Qu931MRnCNElwWa5
8ZK/ZrY4xCwwppjFn4T8DzhuH+tJy4hZ071B5I1fQMn3OXOQcMDqLxso/mkFkfFw
8nYbUzsMCMIivJH3BLYHQGLimxllBuOSiqlVjlTie11PRWsOTd5mmvBRn1A+Zjjn
vvXzTpJRuNnLgpJurIYkNKXo8yuL2f/gobyAknAOSXslAXhlmrUXOoNTsGqeIUEO
9iydFfWeDF7vnL19ON29q4PUhpSvUnp+kGorI2ZXEZ4DAZwFkVmj5gillmvUCmh0
KOLwvuMZk5BOGcQ7f3aFW96bUMnpf4RuTyH4peXQp2IVDf1TK+kBfHusoUcku4tM
YyrEDl2gEl09A0+Vp17a3JjwK4U+rs5P8BEORrv+pyxsacT09k5+F7LiaUKNnQPo
f7nhjFLjxa736jpHJjZXYszYEh/SxxgDkbv+GbQ53esRDdorCNimvU8vOOrHfmlv
B9Lqf356rAvt3Swd88GnW2Bk6CRSXurSQkwDBzwnT+PDm+NNmcrtRyufwPWg9tZT
g35ekWuItlMW97BBCf435BRZt5b3QtssuHdVK8Q2mykp1LTgLvhCJnCsH7CEzm3m
8kLxcoMb6z9M1PhZgRvBgI2dvJpkpo93/0PTwgIWrhEL5Z2MMpOp9zs1LjzLkSVD
CP7LtiOfg8s+R+8kdWCsQNaGPcQeokOruMvo7udcMe8MoWZMoDfoV2EC2YmuTMTJ
nhoJ/RO9nTqskEnjBjEN1wfBaNH5reTyu/KfjoLbkMfcbmWmwkdFdx5L2+FHFdYk
p9hvPn/VXk8XL9pAJLsHA196qhutn0ZDtR9CK4RZ0Ji6rsueEgi1XsEAqISmroDk
wcvYzGoM+41y/33LmfKWnlf2QxOB8Cvk4q+1q8k7WDdBYmI5W/hhf3kug+PeGwQG
Vs+kyMyTWe6eKe8ajIyjsTSCsNAHRvz6VLj+a3Sv8DdjYZluVQk7Ls1uJHsW6S+2
Kw31y8cQ3XW/momNEYJ1YHDuUFgxyuL2WkePyXDwA2DyjuGsSCNIGUlBNDVTr5az
LR38PuWZZkZvHRgnWreBRku8xmUnDFoT1YrdvLEl7uzAVjB3AWyM9LV2Ci9Y7Q/h
6lX2F8fAr9dwmjwKsPxNOt0ZsQphZZptbtVHWpuGhjsBJgJp09gF8+gBTgI+QiiT
EMawOAI6JhsmVT8qqtVnvP90tOJS7ffkBIyPhepCpGU8eC6jdeuWm4xNPzf4Yu1l
lpEXWofBW65+fVdbmcj2NPbqd8eYQ4y0PRPl14VIKflx65OOi4uFQlropJUVtu4u
gsta0vvhO3LaUkudKYkGTbpziv6cD9cNgb1/erdhXuGLX8btGXd6ovMknbfpkNxF
tNpgxYAfqIw2MIL0I4dGA/EEa1awK6mv1FMAyiTXFzlSG2OAKyXB4uGSScb+PWwU
1YeMCnaY4aLlD1D2VN13GbjOUSeaqsE9isWt1xW1erq54ap0i3EeAfC3U5js6rKv
Zj7cB/nQ2umU3zzN3l8RXfE8Him8CxLeWiR9ui8328YF3iM8dKEY21kwLkEL9IFw
ZHPPTEFSCc9XLl73Zu9sF7J+ogkZ9DV+zXYzBfo4RVOabjD7LEojsr5puBFl3plU
7xkNYsE7HuUA9LKmKYEv4srJasVNFKzvljeRMvoSKkR5UHRoegdrxntFUBSO5gca
Z0s8sHgJGPnd+Xnm/Oqv0KAbG2kAn5cimJWCYsvF8ZW4r5GeqvLcpnRF9dZ2VBeQ
dkUXenZH3BUIXJHmdsGVPr/WQxwEJy+4Y7Hc7LyzntX025hVNB42vcdOSdxL+uTY
qeMpSZBpMsTp4qFvxVLorVsXRvMq35QM2lOGMwLkyuNqyYSF53ugeyj0onwDz6Nm
9c/1eZjw2CFq19C8j3yfb7RfDWE2jsmzWGR+x2G+w1XMdU3D4SKjMjN6CeLxGLjQ
VOJqxkgbssTmPqmmbMnVktIfGvNyQ3ZUoM4TBASaBsW4HuYYnfsS0wPIlm07CB6k
22Pd0gob5Y5CgemIXseZynNEIeElHO9pfvd0cGk3Nc4YW17URW3H0Sq2dFEPWVMM
LE1wXlyV/d0IZJ3NSJ351jVvK7ncMSfZcuvhPMwxnazUTL6ZMcU3tykLkE/V27d1
pzr+qt8p6KnnS/u+AKdEEyaXMCYV1SP/YeiB3qdpRa93+rtMAa3pbarPBl9TKyXp
wn9USylDel4GmCt4HxEhcvqo5MSeWS2Y3k11AxrHvtNaze45MaFtyPzlczI4v1/8
Jh/b970yrIwqV2UrAH9cckREtAgRIJMUu+lASftYE3DIq4TlI9iSga7gH4wmiaTE
IXLFLvYRuUD3EhMigAbesrIiHAXek8dkUiBp8oiZ//oVdvR5XdzHg4Hp7eugSpSL
5xnZzGj4gN0r7tm6iKkOzXbP6lDqOjRXgYyCzN3ki8rebB3Uk0m59e4NtnYnmNX7
TO3Pm2KLEi55Ob2+I+yfLMjzq7sZy8L8RdSYAzMQUqlLVvDZ04M5iVZvWRDW3jAU
sqcflWIANEgbNvGrz7sQxLt53tTvp0W8u14Zc6FusyPHxYiHX3vY+4Fi43Yq/vd+
bVQgy7Ra5hiO1CKBI1K0DqKYVcT/ZGrsg8pJALbOU1sqPHRVZhaDvUB8N5GCVIhb
uOruXlDINAz5aBQx1WxW0mpWkRyVy43RGRdt8L6sCOpiok1jWxVjXNNegBS4Hz0K
WtSJR8gtME1V6hJy6mgxGsrQAEssn3Gtn2B2k23U0c5WSkysoVX6ZaQV42JqVfM5
aF0Ns/vkrA1a9VXvf5Hxrmu1fUnYv7rW55xO+sL3dJSGKYBCfYlDfQowu4km3+VB
K0LVK31f9oqODTSu08Q9zNDSuscO5YL7gyMayGBnlSGiQaAlU6LehVOjauvDOOmF
N9/xnLJM92cu6S8A8Slb4hgmihUVrEJZVE013ROGpHt+nCSf/1wqZXRMO4AHgpRi
mrGcCyZybiTEvRCG1KU8FIXrbKH9N6q1dFAcZakO5HuJGFPQCzVw7EVeeY7RIdgP
TLyd0QYQFc8g9QQv/PVaQSnIODC6ueRkW7i6j98/3CkvI6ItucX4ySH+t21ZCJR0
KQvPSy/rtHC/pJR1qH4ASMISo91ne0E+2k/sLv+DFkTwtUZ6Zf7AceWeymNBgfCw
ucTvUeGxRj7UrsLUMYsGHOhAQ3AP/aANOE8o78TiY39p4Xe5rNrQoGbdePlgTei+
W85pOR6JyYp7Xm9xVd7V/KYbtj0I1rgAtjUaWY1pXQRhGyITDZlDaFjcybd0Knc4
oUzAZuN1Ce26ndMe33wFtrXv8qviSQWicygs479k/yGtv46tlu8zuSc1I1M6du5X
597AUKWc1wTE91FZNBOUDcp9UrU1GSoZ//5FzPaPeQXdW5+8YBIxsE7duBnaIiHO
f//AhV373cYsCEFpCVUwoVpmItZe4pmktK+tUHsLe4MKUBlLUNIQrnQEtPotimZ5
0fDBYmRqRquG2naEYjSd+/G1k1fDo1hfbdsJde/F7fYB2fpn9+L36ugELdFSRLIT
6OSOJ0ChhZKpyPwbRX/dOzvjU6xpmKe1IQ3f8hkTuyNqyBTUn8m5MYsUT8YaxodY
EEhvCnssbuv0RMSUOoJWd0jPIa5j2VFS21h55yb4QbttPMA3keYkgKg0tc2hI+1B
StJV+iNsvE8rQmhOZFJjApwZ7z8Pdt3WxA3g42x4JoFi6V9fJUzyjk429SkZVaW2
441L42+LxMD0J6r290q8pbHyO4e8tLWjLu/QIa4e1aRYNp5MdB4vXaNg2FkxTXIE
q0Gzhan+rpTjPfgRaYWdC5w2nnX7jNB84lt8QciWMf/ACFsH51zUxKX0aHiyBmTT
MjKQtbu//LCK3sTkUSGD8cZhJwelwZa4c0ip+zFmQNk2whVAE3eHzJytjoIWTF54
3Hf/FH/OtdvnRCTg0yKB4vTH4AyLqyeDKDQg4l+lE6ZmDUJzwa4NSaS4Ih0kLc9j
0m/HUQzyZRvnn0pSVGxguga/NfD9Sw8yBioTQXamgDoE2TnqF6Ea6oYgTUCgOsSl
PqFgDV1VvkxrLsByvfRRsb4gqDut+6sMZ6oYJAUT6ywBsmNTWb1VId0NDWqgUNWw
ELcLtuF6lp02ihDM10+jo/9j2d2H0Gn81hbugmaWMM5AZM4zNUI/LHkpm7tz06/y
rlupkBaXb7c/LcGaZbt6Bu/HiV4SWkiVITNRIKoemt3snXM3GfByO8CY0EWyZPtV
CKVjIsUXzOWJ5wsxrGJz9DlW7MeluXjftYrTEgaNwzgtONb44GTXmeYAd3wbOYkz
3lOzlhuonfWIsxxkzg8+gu7DexCfjEIl10gP5COWNjaTNSQDJLCnz+AJ/HHk/+mn
DM+v8kHDw0VbwtIqsu3/sdLZuBiuv8RbsStjE2HGppTmb6TYbRsHIuwQhRATZZDd
XMgEn9Ongdyah2lZObFe84B/XcCj3/WU5HyJJ2gEsg0YkZ3qnKtoUQTC0fmfWjDs
a8SZThoZDIhjo+luTeKZPD29s8rEd2fJvZuV9pp8o78GgO2//taF7aX06H+jUs4p
6UasBMNTc3Dj5Tik6vJeyfB1fVebU4Y5yWRziwsbwhNTFG4YDHJR0+aDL1dLXA9X
42ye7gkxYS5UvyPLTb5vD521pCIshkLqjNY57Ad2rYKuIgBGT6YOayrDBa0Z7/gS
QHVEjH3LQEUPl5USDQmxwaPkLXzyZCtWvhaoJ0JnB7s5vYoMjUQswRbYzV8xcji3
JKuf94lDElbq6N8/F6uPFMwSlQJr3nkCjd0jxPa0cIKsaUasUjmH8k4O1LuRQyZK
dGk+pZGZXDWWXmCXgsmMUgnYe7hnHSZQ+6T1IY8W2kd78/2BzsPf56FAU2xWRXUm
x2ORK75poMm1RD5rLhxehctNKlL+lLR0v1iHWHKcCNWi16WSUtGUH8HjyBAqmH3G
wp4p3KetPC27YRj14kaDccJqwOPONSPdmZsV7cZkyeeg7HG0n1pnN9eHWrfykRap
DsxmyVlnIwoRv5cL6TG5jmj5wVOftjzz1ruC1JWVgzaky/UjGJNda6eOuA6UQ9r6
woSqcyxawXn0/aDfUSgQ2VBSKjfZSb/zs5dctyJrn3tgeym4uKm3IYkKYOBp39IM
lw7HDGnIsK394rEyK+7Ay4vYaQDjBTJ8h+B2yGFHLbBl1O6F3/9m07AxL+LbxIbh
UbBwB3xUdq4v5UOZ/HetWzi4oN5weF7DW76aYh5UzoDi3maUF8Zwo5qMy81cYyZH
RYG+Q/ANvrUVpk+RS0+QkbkyW5MbaEhf4pgVKC/xsSBFivOMg8ek1DwgY42Kkf39
LLMJPdVusMzm6YvmkKMTvGyVxL7zsAcguJ9+dxQZdgTYJoCmH1Pt8x84DN032dJo
Lxc5xnR2st+S+1ipFjmxJ/29mWXQLtDvQ+IL4RiPad4ZXeXdfkbSfKNAKWx2m7Eg
v6Zza50+EHKF80Ts2lggNn3ZCqfpm6c1FO7DDU8Wi7n6Gyme51hIwVNBD0h6DnJ5
cKKBzNIc0owERgdeQUTQ9y1itSHwDUyeCY6VbihpKJ53fs2siaWlKz0r3G6XCbse
MbqqoAJY+B1yC7F9UVIcl09Fz0QInlaG15jGOTVuisP56oFSkJ7hTWM5vCJ1A0nd
1grXS3ANGMRRXCFZW5Ahx8GQuXFzlWoL/tNCzJHLhDOxbC3937dycspT54HDwUld
tEI2OQitXXTZLJRX/ribKmyW+muTxKZKfa5yklxkCn2p9SiRI5j0siWvCu/3e2Gf
U+E3xOVUzHLow560DWor/rrMFO6yj2RW9CfY2k2sEhe0ks/AMdI7YGPpJCB2SPU9
jEz0MHHHz1aByOYXju+ZIhoYQrbTgByscp4gc3VQVHbV/7mvIxMviawqzG/Oeaqk
WYad5i/B/HQKnumULtAZcFB0Qx5cEx/UxDHjRJvVA1bzhw0UIyKEZnRWrJVEjEFO
WzefNymFSLrLKkZvT9ZEWsBsYRaMjmawRhOEc7ml8pJUrdWrtzZ/80Fzo9oFG5S7
GTpHuafnDMSfQSQDFAjHRZKUoSgkQPQdnM5fhUthWISSlllyD3b7IL7zJH/jVXQt
UulmL6HYTVgL0sAc4q/7KoFqycNxSja9yYIL1EVK3V3CsL1vNxpbYe4XJPL06sCs
QxjCqI9Yc3Y5G2juGnkXz9GBTfkJfenMCiWUUKtYGASGLsx2VphmpmecGG+gjtYp
dVHZuOMHmRbA9TV3JJ1kpFcF3QNhaK+LeSs3o2Jp6Q/HdWYav06Dl90ZhYkGMdpP
jJpPSfq5XDzlzPeYp08q4C3ib7jlg7UAD6xpkYqfwIfh2olo61I4dznhY69oTMNF
nBjXfmPP6pFnHeF5V9cPJKoj5wRkvmhIYXgLFIY6ln7BiCHpS3egcDkeIiHEBFGK
u2BsjLWSHwJLVKrjeHo2Ys29JDjZikWmA7H1rW8T+M5NkBo2OLF3SUfD+aDaiBBu
g/Q9QYWTneLCurxUt24TXE3dDl4kVaRY1KvjIl10ZvWeCRrHQuy8Le6Zekzx342e
svRq0gJTTWJ3NrhLVSKxy2X/k60xbtmYyGfEoW641611ZldzYkmZGzc8B+gf1bZ+
/7Jp18wKHAfLQzQ3wGgjGCpmbUkhiGlXJc4B0DI6j7FngCSSCP/TD0CW1Zj8tVkI
E5Bp8hknlLNz7GrteUDsH6u0wbr0O4p0zh2kOZO1Re03y2sMmHP7j/AZyzgOju5Y
CSloDJiQEfDDd325ow3haIeUJM2thDU7War1uTGSdg2obO/fyCzQo3/drZ3/0ZZG
LTwLvxNKZR4TkkBsBkRSvWkw8nLMKQ+wJ8HHebo7igzywXb7Hnyqjn8drrbtm7km
Ft73ZRMMXasMtiaHcaH0Lhze6HrnPioFKBx1uQmz+tPSu2sexoEq1Q/GwsKAKUoa
cWMVzkdR2WAn2ukY+JfT9iX79dPMAeCG8vB21EBTIOyEuTotcYAj8G2l+/7Fqxoh
FIZtUf+Fq2OOrTyengy4OfaXIPVzwqjDZ31CfL9hd1/MYucyeG8qi7qddUDI17+X
mUanH0sjQgfnGkU7VOVwUpwvX1MUeimQT21MFuNnb8psAH3283jD8WCiYoht1rPC
ASmMlsw+4xyH1pGbocmnDURKFUJ/8TrY4xwkGkcoJ13AcE6jD78HU1hiAIOTcYeS
kd1lWC2ahuHfsWAxOg7GOWFetIpqq8rJeclTwU945eWcQQ48FrpZ7FyxD6AhWtUn
OF+E/uBTlwoacMgEZ2lwClik67MVXN8LrWlMXNpTjsfrrHfWXK4KtyjmJLWblQ1H
3qzkQz1eJmf3luq/5kF7/jWbxPBivmH9R5MNg5rkkBblI1vVRvSEBehCXJTl4Yh/
W3OxdoIKHsI1OaA/dIdJd22ui4yHNEWopDsW7B3OXsODTi7zNq203wHEndzaWS4G
Xgno5NdFrU3BT3M3VGjZlKp1vUqNALMgtLpL6PiRWksXj/JU57eXQI6NJpc+DS/z
pBapwT/Bg4aVs+qoNuOfsGuOZG0I11NBGXoQ+iImy87IABgcVN2wXW2hm971tpSo
QZgibrFep9Zpsly4BGqbDxzt64R4D/HHF40B9cpQTW/ImgbLkVVeuH5e4cg2AsXU
DeTWi8pgtfPSh6Zrueclm8L5t83+3zWJ3f4WupgHZ+x61CwFERDS248+BpCPYC/K
KVax5jo6MYB9DXVbNYjp+fYrVKnNMJiT0WCoQMXPqGugSwhtk95ACgGiKZp0KChP
E9RR37qwwdE7XHRda6qXc8iKJqHAWusinGWjGUmcNl3cnNglUv/Kp7rajCmlc6vT
KYJW0yuugNUQOOyDVgnUUyV0KY+bwA66z3hGmXSr3fNt+j1JzainogxjeDfBm+1h
07cI/55NByEJiA44VTm0/7CQtKKDcqpJOQ5xaWXnpzJtkngpbng53LjEjKJLxpnA
EtLFOzYZAPsea/zTlaOaryVl2WBPGLEnhEOHGbdXr/jeKP7TdC0E8v5lhvJITKe5
H4Y7xBe7EMAihlsuMgtSmM02mslmxgBUk9s6sL4SZ26l+DOEOByrIcNK8ueNt6yg
YI3rxxI0bbFc4sJiNQF9mPs33HGX/aIsQ0CFgglBd0VRFY/q2eTkhBYLBUY3HP+A
HwKLlcdHsZWmloIQu1yCG6J3n1gREDoZSd9+Xf0fMMzolL8uLdkEZCdyxPXIHcgJ
dzOhJZjyKRzELguDmrcao834KhRIj1Ygzhe4KTl2MWj3G+6Giq/hRYHNeC6ojmgl
a6Srq8Qb5vzMU8wgLIPS1eCIWtBTClLAMXp+Gc3KWhxzpZz8uYQZk0rYGF2w0D2h
muCB8kOVf3V9R3pqEUA44jV0WvOeTLZLhwtY5WbchRPdjKwUnUpG9uIwGePmhSgK
o6fpd2cJ7vDHx8tz67JlcRSRsREj4I/RNWcvswny80qtVCTyPU0r9wrQv0frOra2
NcMejpRrHmqeSa+XhMGi/G/D9R7hqWJCDtbyLkR2Ai49DsmFK1n7P9p5HR924/kx
w0UJ8FNLYkI6UrNDDKYdHTlX9QKZ7vniIdgbx/6qYH6pO1/4Xk1wIZhX4k8iVFiF
Y0UTOeR8l7tjHspjyUL3sq/7pgFsotYwsyCvvCepbus7Xv4pOn9KjkFJ7aRyuQHe
7CAW2+70NUjXEliIjHT5KP+8iq15v0YLDkwfZB7pd4qe0i7kpx9XzShX+yb6pv7E
ubCwnws+17i0z0RZWRHWjlHFPr120D+2Of7J3KjGHGCokoVJeEU7klktOKVr3hrP
kDrQhBKx78ITYdymKmy4Qb8osrs4/0qjfk+98+m8Q1GInLTqMJ1ZZHJDGF3Z/35D
yCWPyB/3KdNWjT2pQvknSR6xCX45FRmGIFJNHxCeTS8ygIQfcppxF3G96JQ2/uWJ
cAKuoif1ex21nEn+u4GvoLVilwkvo73vJyeAu4NBSPeg7652SzYLEXQZdfGVZzB9
u3nbaFxf4ZGsB7WgXDGzMApNaRAL3Akttky7Yjtj19njQmamkm8epBDPeyIZ+buE
XGxVV4i5hQz0JJzbHD9GLDg6EByZhgbNcMF6x9FpN4v5Rt5GhF9DmAj8TOkxRUIv
1lWqDYxuqoE6nlQRpxM7pLOFMMamnUp6c86HXEkKlhKUO2HCIHGgdSI/c/0AnlLQ
k3fvU/wWmJ80E/n/armGfuOKAs84KXUA8Q8Tmo0NEpHCphthylk/FmXA9CGUgZvx
B+J1KjAQ7CRm/1b43FCyjatHBqnOAbAnX5Qg551+qsQ+1mduyk/2hikVR4DqdF1j
gwm3idAqmsZfqAPpvprmaKrzlx28JnaTg+N/mRabFJbIJnclG6Yy7vJd7uhccti+
JGfnQuhgW7Q/jjokPj6FxhSBBtsvxSV/c7duiX6bil/Vz0TiNhAtd4UyGb7LyHRO
B/UTVuHhmZrWWPSfpx4jNRd5l7eZWuQIj38qKPS/VwhPpI+bebqhG/BPxWNxPT7v
6dvbO1peKIRdCapv+50/qIhv4RRpBJLLPPJYjYSoRpaIEoOsjt91arJZYcMIDtTA
v3oOlRGN8Z5SYSiKU6EUv2TYzd6lpQHCqi+epSiWgWhlWvp3882vBbdWZqA856Sa
TH5CqSYRS4I+KI8x5cuQvG8djVR4TRD+pgsow5xQPioH/wIgbAz06v2zNLQNsoo0
+eyBe6OoUbDR5YXlo5HIx3G+cutDXpJKi4cUGKQUBzGYgZ6LnoZ1iJUB7UDZOhAH
pYV/p9Slx9m18bc0IJmAAO63m5K81VrOfkX+24Qpf8dPS7lz1bnKi0wxmK9U6YzQ
hpwntQEbXMIif+E0nsRYC9JSOIxZbMZMPPORx2oPM13f7ZtxnbvZXcHTU4lAH4un
1J2bxTDkNrJODwFf+MXOkpIsKS357/G4r+YyM+j8zqGef0IjMkhBQeXM1uW1uRUs
ndRYvXt+6DJdxiSb7S3C5Y/ZVkM5JZl7b1EbMrveFi2WutAY2NXDBsP9w3Ce35zP
P1jluhtgdN5GaBIrv1wBuX4i6frnKz2wEs8T8ikCt167kFle4C/psqzaQzqKwuSi
bGXUYto7D/6IzwNrdbUKxXrFjCJmh+ghrUm+3QdTfj9H3XLBC0e1NbsphtKRGQYY
lrfKd7qp1lMkMMoc+4CKLS4CVHpk5/vl7JsFgQFRcR9sHw3vqCqXWZKVxLqd53ru
C6GYqXPpEDkYHrwZD+vcOmO0GWQLjW8vLx4ymOxq34MYhJtE7A7OIdKYjE1IOTcr
xy5Yeg7uwhCH/XIhdRlZ4Q2wuxUNAT1bnV0CLiYXQ3nZZKAFE+9UhPnerKpB+rG8
hbZr/JDUjI4oScve+mHvbDhSAFUIhimPPA5nLTOYyCVQc6Tzp+0cSoNNJAvSlDLZ
dyQCn59hLKlpQxvUCdg34pOTCx3HYnBvCoRnJKQx8h5/u9y9Fjw1pCHFoHgvHiUd
nuRIsk0EeN57oPoT2/FPe1HMAFZ5/j+JmvhQaZcXIeJoiN4Fts/QItNe7oW7SRFR
0q611BIpOyZbe4nWPppsYdcmPUGEkDV+yyusfVDfyyIkSMI2qfLwn7uFTiGzPSb4
Pf4pqC9ywnzcxjmVbtZuy7RhrGrBiynDJbOAbNny4TJhxLepJcVunS1Mv9M1sUR4
jZhOXSC6TKsMNPm+6A5Nd5olxhKb+quDC9woQFnFkcLuCZM8ekafLvVZ+ZsaC6wx
c/g/S2N3lSU97bcop3wkSRD3ERuhfpaszsX1sfiV1OKyb3w2b/uAyza3A5IGX6+y
ibzfZgtv6APzgLex5y30Arza5YK5kBOd0g8EhiePpQBAudQl1/SV+8agrWdqD9mM
oHAN3kywjCCO3fHqPZisDLTG6cirLtMeHyoVt0SfidjtY6YNoOtee1GFQQr2nMMb
vk/v9+w+7OWgi0mONq5vwY2+IBXEkx0Fgb0lURboM2qsl5ez97QFM6kyRbeKeoM6
081t2W7ZzY6w2rwF4qg8cF7LUY5IMYSA7d8kgLmXZ2nmgFRgo4YFSAt4f6Ydg372
F8b+SV9OzidobWwUCdr9y0xPdRBfMJ40D/tL0pXmDHWpW14u36hyYW2emN/HdRA2
zDuSOplNrOvbbSrQQCnj17J9g1bZSqpQ3MQUskKxujx7mJ493LnQ4OccwwsmH/rA
ECbp69WX2iCOZMOaBCLQluePJGY9va6XHVJ2wKDhoy7DGSyaPgQ+Ik7zmVb/uVWQ
9OaTUxJtwti3LQvoPOnByNQn8kMzWlsZIAqhb1rjQsDa3PlXmI5TJlKWOVpmgqFr
Ls5Ix5gmuwW7/gGzXrda8vI4Et9TwNIYmmvAm8tN18HIOY/yY+AHk3TXwTOfaLX7
cyXM0TruqGBJp6BKZknabJ/MWl5UPeViJATqj+Mo93yo5o7HCRMWBALkaiBn/0oy
xX+NikPqCMsQHLAS6oIuvfux8aJFfrLYJgN9E9WyA10ltSVwyFEI7xqYWtdDl4HL
CW0IlD9kRs/G+CXfysnsKIdJTDn+k/ymmucRWp1rPeHFGHQoxsPVHFgrgJDDVmBf
/evT9hwJUooOH7eBbJr97tbL+TGAeu/GoxcENPx6qkGtb71szG3ubBcyWFP8kDkg
/p1uIMPqwuv+hGe8p1r7KMd8S31215Hwks2xvLeFm4s4VlIHO2IR7BWTL4TfCWT0
fqHzcC5Pm/yXRQpUPUgPI6Cptjy91jBpBsl6q0LdiF9V/5ssJvDQPhLCY0f5fkCo
UKqbNqfKeqUIc5hrgNoc04a86jN8OSj7ynjfV5KIc+IDMGHeNXsu7rp/OZ7l5hKv
8n7H1Q+s9qmz4jB5ilEGZc1dgduNFAZg6MoXHltsdSuOIboRFXQYb9ugJbc8VFT/
s7fAH3uJl0g2HAm+JKu4BH89rIEwqGlNjq+RT2c/Lhh0CC4Xyl+tYO7FN7+CIvyg
AQx8rX/VagMvyFAHryVAd4CrrXHjPoBDFErdzdpfHv6edNsP+oG8wGK1H3JHdjk6
eHsDBSIRgX8a2FuWB+CCpgqGtFwm2BNkPjI5SRszuPbI/oJ/oMWpWlkMBXqTbH+9
MSmBpOjnDuTGCMFXAwQx6XXyk34H8yN7od2sLh6UFdJJPrOSblUg9SfH8VQwxxEg
ikqB04lINeXBbKTmay1xp9p+oGWFcbKfDC2rsZNWl88DYjSU4I/W5iFcI7HgflA+
Pc/eKihIxVmQcGAJqJzfXFWwCTkpomEagtEkzQ2w5BPuRLT0Tusy5qRZx1gOCPTT
u/GCNthih0zuaRihoavkeRclpnDKnS/1ATleVix5LikocEi4jJIXt2mEs7fZ+X8I
vLK8CXqwSnK9GxxQdG6bcOcHVltF2ZZMt/AcmOQ5Bki0zpxDK332hKWL5rbWyk9V
VfPU3zwf0YTSSnM4CIE9nFmxAB+YbGYFR9aSDpXCZpLioMx67zwOudJLFWcVMQ4o
a8BDRIXQo/SRIRQZL1Pu84LCGJdXelmvRrCEwSscfQnG8PKtQzA5Gj0rpuCU27lN
mOH5lJr3cRDAY/rphKn/bv2xdN9B0fMeqY7NlWhKpmUcDjJ1gwJq0WYnVGONBiYY
lYsWlc9X284QctM7gfrQ73zzr8uJZUdWfmltvjNAdGCVKDOb15txbmjFRLyF+KYT
znbogh3BRCUq8asT4DB/hpspHSQcvXxqBBU4dOJqOvzoFir1o7TXYjQlxx4tSpNq
BTQGU9I33dvZ3XY/YTu6WyPzC2Esp24aatJZd0jyZSsQQddKLvcJeyS/vlHomw2p
Lvy7S5CgL00TTiz1R79B0vlobtI3GCiI6oPbKx3gdJNT19Tbcq1i224IBV7h3y2S
k6d7qqdKCJx1dD59yMhrgOJf5aI8Ynxts213zx4z59+9tzmacBi/rK0M+gLMT6Hr
fW9voCbP07L6xgM+b4ZWBk/bwPlZiotppoLmsTPrxqelDZtLnXbjboKlnYD7rLLk
2DTw1UIVQbMhcQof3ZKki8VGcEDMTPoJabeRGNI5+SstN9u4Uzr6qK3LXI028qkK
Ey+uzoiVgGQRO8Xg77IRnBlw+evIvCmujUgJN8gWPWSFfGLtM/bIoejnsaRCKgCS
vcJkHx2jDlnjVPACbA/gqcdbn3TmMsjJkoFXvMAjvo/PNxZkN281+l+h5Elt52QF
L+2xgP37XhzCR4t2QFQyLg4NnKQ2IL5Ed5mUF7UZycnR0eNdRk79oIVLQEBxnA88
ARBseM2nA83YJcAPnba2nuoe75Im8BK6qo7vB7PWUuX+Xp14BKCPWyImQiquH9oZ
hUyqdpDOya8AmMQl/hm26MYTne4rvR50+LiOWC7rNom5C8uP3t3SWiKSTfR1999V
3M6RmsySe5JiDA9sCxKpSNCRDsDHSi/p9qv7QnhKt9MfxFSqx74jc2ZwtwU+N56w
o/zuJllBnH8DJ9R5p+gxlJUtxli29Ottb8X6w2GGeWwBi4ls9RrnEWXto2irlQBd
cR9BXF/iGDFifZZ1HIPSB7fKJuC3Tm6fxrZIPKyY6BXB8BdDkibbdRTDavbvJrGP
Sxd67hbtFrq/lfvAp65Q8u/xFq2XF/COYeYqpTYhLiXZwQRYjP4hRIdYp7l74utY
Gsjcn/lR+AIJZHeJM3fU9VSZAP5py5IkrGwGXo9sSK9a89v7hCArsZQUIzhMZhcI
oQBUYSySAC0SjfEKMsp9eCu8ZDFohOHYl9zSWE73kNzMDcaUFMQ3nN6ziZMiIzyu
e6U9LAohXTVqemTxT2tcpKItcc8ACavJjCuRye36Ht4o3yGi2skIk+vAQQnQwqpI
oZyffc+M8mBTdrSXZj8XEIHk1Tk9Yhiwq1mj30IBa0ru3TDzJjsHOftRPoik3CRI
4LlliVMIoyqjHRKAXC9vtx0/fXTrgZ6jSBBYgm3DCrdRD0QaG17WtQ/lq+A6lC42
cPUoZptGbyRPLkXbKRP+NhHDCnGJR7AHfigKoAaMGPtE6tlpMiKQaYiNVv/SUFCz
Taoyb1DA42mEBNcpKi08/P5vnVXvgpI5bzbIWad2b21LtFKbGH9UvCenq4OtrlY5
3pmoGLRoZGs9dck+TrKbgKHqr4BiNPwysdVvw/NCYFUh9vxpo3uYdiE59IG1jl7+
slRopDF1faM8zhoDSKY2oTgBBopz2Dhrl12Mpy8DA5cxHbaimDYh4VOGArYvb13d
VX67OkubozTA+BWVLhKziokk25h1uveMUpjdSspy2q8Zq+/AFzd+/Ipa1WSGbxyY
I3eA4bpQSkqyEiknby2GAzoHtA9rh0Kz9os1Q4Zf6p81HRpYwx6SUYneBID8n5pV
MlBggOWAhuCKwDGDhsGZNPVrYiRXv8Y/mTrCIXL1P2D4HZRlmGnBjHCwprmv1adT
hfTt8DIJvfVDPlvyB4b9JBrRkVqf3JTw2af+NNTCUtgSW0+Og/z7nucNnk1CdPYw
mjXt1CGXOEQai2nl2Ba+u3fwVPZ2krrItFk2Ie1uGvxgczwltyPiaQ3+CP55pu+I
WT2RXoLPa1qV96AkiJ5w/jiG85nTeZOPjbfqune+vUSidgO73rOhos8hw/YgC/VE
RfGCWBN87A3jInVpMifsnnd3AIGZEOkn5eBzrZelEu+uiOHSxqmBb/j3KQX9oCNW
aIcJXq0iRw43Gx/9lT3QWIrRGNEIDarBbX1NkVBWHx6w4lMOVRIMloeapECeDPir
4FUlbBEEUYmHcxBJrvzWxohtMxxrBslFiscPkaiTHSk8T0IZDtdFOwgOa8uTgYww
Uj0OWAjXZ9IANzvp9SnFBDM5mDovRFWx0GMqptR+NLhutogbgi219r8lXCf4G2q/
OgUMHIB9KievoyawTlphjHDyeLROHLjB+lDAkaXgd+BnC2PA0uztTT3AsL10rECg
3BAIEQsDClbdyxtsqeB41WAnQYOML50Dx5MWGDU2s8rh9GwhGXNs8G/fw1+V/Y97
g644TQsOE6HvYfKahQzyqWt+yE1MbTB214vURv06gM/yC4z63MBlTO56YyhFPiCd
Ss83ChEjZGulNxpDZ30V2/q+nG3xM/nGUnP3o/dLbHNHYY5BgMWFSdhsQXLpBzIo
3tqRM/DUelnREoxxqp+tZalLX0dsoShy5JUF5g52yQqHc63NqKeJr8FnLh66MdSr
uwkja0nGSZSXScWZChsQnElaWTz/XnZkry91zA7pKFYkWqEg7EgcYQNdCv3z62j9
9KyYpmV2erKtJBSFEShMEADk5Nf8ukW1oePFIbbmR7SBN9QRt1yn4R0AYvTkjt8b
no1T2wcd2lo9hZ2NCUZbXjIXvQNTiZwrHdawlgFgQFnCrVi+gntqAY41ZdKdh2Nh
VO8Yg9pQedm7Lc4xqaFqis6s+TJ4qPtty+eRsf1fgTrnhTiBdtSqeYdw1T4FL8B1
o6zPyqYTtm+lMTfzEht5E+UGOVgR74RKyBlxDCqbJkAQTZJFotd8QQahTvDhOz0w
8Fk7oyogluBZ8CRwzkrIFZedWNdLv31gSw/lDbYHgX7jImtjfOx4R3w20G045W7J
e1uLrkl69l5y7axoeSjbMGQWFVJMJaIfU6AdkSq9OIPIC8UNG6Uh3XSu5Lx88jf5
I0Dwvlykoh0cPKKgQmQ1LAGmtlfbpB5499eF06VB2/e1dN0qMfsQQg7imw6NDjTH
yQ8FAqJxsNnMrkQ83b7NwNUG35fQoHxR/CvGQoR9H/E=
--pragma protect end_data_block
--pragma protect digest_block
jBu8SchBbJPpTyEgo1DdR4fU8L4=
--pragma protect end_digest_block
--pragma protect end_protected
