-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XNnJBKF3p657kipAHITUUtpnUSgpC3BdWi3ZOguLH02cFwk62YrYjzwbIQP93/S37wMMwyJ/lK6M
tZ9iRP26s2tn+HKV5pyN/A36jBcl2WjRGHt6nTipmSZOvQVkjUOFmYWiSXhDPd+fFwuSM7n4VcYZ
egd55oJbqnXQsfuxTkunULuP3gsnp0zMyuC5GJnX9O4OPe6R0lW9HS3+ePIXlR8TxxCT2hW8HFFn
HCVoeAOr0qCZNo9HicAb60YlNIP79xduGpKlWkEHXOR8HKjUYCZ2+PmauCEJRpOCTAwJN1NGmAFg
ippsjCb4lU3N8Kr2uM+DCZKP4i2FkW/AJuxNNg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6448)
`protect data_block
VH21xqOjqlx1YZAbb6Ifdqx0STQeyWIoHg8JiG7cU2ACOGiewJX4EG08rACZri8c/YWOwwm1J/t9
/9LpNHjkxxKOe1ipMFZzgFEpQJBoJ1b4uDnJUX5k11LJlUo0OR7MowKLJfGP5I5ZoCtltXpWZR6l
a6jWt8vF1n4scHrrshBSFIeZHeC+0ZUxme0YnTK0oDh7nVtK8q5IFhcF4n7I36WqY+lhtrGnyG0m
5eL4m8mjKhWi/0s02HLv4Aj/vctEGXfNe46KqCZCZsCvVmevJVMBLO6TpAoAue8UH8YwZLdu6+TI
I2OsgufBL8bBnNhRccApW/V5Pb8ZWdN4IAdQa8s34V0un0OctA6iOkNuvXitrABCx1cQjKzfuJ5b
4L/N/o0rGNojZyFXYh/6/awAsPLPWXN+VgmqaLZdkrVm2bYnDKh9t0R48qAhZsybKYIXXiCdYC2v
ujIor/WbjSbmxNHgrT1Wqo7VN+owPcsSGiODWzQT7iArBCp6FI9dG12owSdmbI9Q8ntCsJM9kKla
/MuNmxELgai29z9tsNRzjRyi1j27w+a3hdADlUIjaSehCmgfscJ+TYt4cxwn35FWGPErH+Vw4aJ5
cpZJJ1w/KJGnb6qZEl7hkfBhDqn1hhynxQoktYLB5qou/AJe8BLW5EGl4/Jb2XLW79JASl0dc/rc
ABKW8E3PHRYjB8S6eaXK/x3Os0sY98gOM0lNJnnjJQPBLNM+6n2SOiTugaLqSoxoTNZbYwNPgo0/
YACSGZ6jdDcq3ePtrxj7ZgOr9VYHUPn48itX6L47ts7Sv4RsrNiKAnpTLNuZ7RJPBJiSypKkle2U
nQpPaQ4dBozCEAKW/XIaUZDFcX3NqGDJ4akBsRj84Q2wQFDXzkTyCklmFf0L36hgK1mvbsufJgZ2
81UDJZaD3QSc/kdU5bderr0f73/RXzJEmgjUT39fIoEg3ethWEjJfPK8pOkr6/6aiIALEuGH3ykq
30f6YBENnWQfdzr8zkkCzYvbzh1YVX5UgaYxUX9SgO/FTs/UUoUXVTRXW2Ci5xW+LYBN2NU1xXoO
qvuCemmqUFdsyLP2iPfy8wcH/1XJ3wMGti765mm2QL0nHEAPFO2ow5USmaGXBhyIjrGdn/DSxnyg
aM4fqKtEesnOjgrCif8KXAbgBRODmrNKOPMDrXjDWDL428UwXclT46FZnqcPHZlUezXxASMJMZdo
bjza6ADlZxav7IfRsY9Ju2SiMwylkt0vquasZely0Hz2QxC5a0LmyziAjP2Sq+U2ZklnuGzb4GPZ
xKofnPXjB4gjgROO2y6jJuFSHulcit4xXq2KiWYP00loGZRyVDB2dDFYTPTTdWjOsmRN+F0R3Iu4
whOSoPqmkDxmGAgCE+DpPOrgkEwr7+MsgsvL4VqXv5a3myGZPt58fbQK7lU62hbBlUhhkGTsl1Hr
YEjy7CGm9vzGzuXtc2QtHgyC/sw+gTNMn/jEMQ0yLIKLkBsDHiyoucEdRrhSWP5Ag68OqybyqWvE
/gN3XC/B8JHLrBXEWIRcFTDMpTanqRolzK555Ycty9Wnq9Z7oVv9NKJZLrgO3UvzQDkMOLj2NgzV
q8Jc54DS4YdmVY8qVhNwp8gOgU4dm0C4Jl4y3Ay2kKeYpB7J5xceWIk6h4yo+ZBYNxUIblMhmBlA
jeC9U6VDtlvGZ4yn39bbRmHpwHlOhk0hwi5wLnr0kw8Wo39YcvLMrGSTSCpEFCi0Fc0XzrxOsbLl
J5f2mQ9teRtiCucK449H2Ryyu2IBmCMtoF7kZQbiku1ZBxPHr+oYerIOS4pM4OsCMh05cbedI81j
V61/zcqXIrEg807570dXuW0LayGhSNhGCg2gb+GHfkwe+krarIE83l/84PwzlQe8vAQo20WyzKrl
aDgc48GbK5Cr2hATQ7JNAy/LmRJ/MDi0tBOzbdX+M0gMkRlz1/sAvRyJabhE07rZczSbLgRwI/YR
3ZhJHfhebc/rFxyl/+qHTUAGhVdFlr5pFJ8tuIxLR7KjM4MToJrF5xBIl+J9YATY9qRztsfEHfbf
lxaLOGtuQMd210OilFRwAa6EZU2BG+XnWjfotQy7NI28mYpaN2RVxdyaS6nw7SwiadcbgkW3D/km
bLZL9iwHt1XvOEbWQfLtHkXtZuVHdiFOJmrDtM2i5o3hZvcINTAzGeqacuc9h494VvbxtZHJccdm
2tLrqgVB7mbh8AH2m8cfTmZ4FBRIba6Spv/14AhLekzBhMXeaBoVRwdrD3kb+2OKLYoWd6T/Y3D0
IjuH8Tx2jd+bDy1fbq3iyCWWO9SqfQjTFgIjJh580HoyT4KdjyvlTX0FBJ0zEV0u6sqBd0G3scjv
ABBFox75bpzuvqRRYN3CQ8kkL+zZ0N/JnLICPUtfhz4AJsyOagbIVgj+ljfOO98lYc5xWHNfturL
S4j2OHazwAx0htVljyrJsYXBnNgXFpptsbG9L/KrziCGDD8jnfBMbccoDih1CdQSbee0lVKXbeEW
uphrkp37ePAta6AtbSZRHhu18bU4ePBj/qhqy1sJi634JnpGc7+EBmxaICFLzHhBKoQKEeA3rNKc
bfzv1zTDBfW2kRUdyTKsHJ9IDOHNBmLXR3G59aTFEul/bMJFQWHw9BUIditWFwsIrd1PNxm1ll7O
H7CJgTkxRMEG26gqRdA62g1hlw5K5Stjt5B1EubfbRfJYJgGLdbPtPVYan/1epNKtRI05jB+uyoP
g9lugpkIqI3tuNbd76c39AbFDpUaj1FJW+TfiaMWiQVWlFQn2SouHGiok4JOMewj6TcH/x6eBjTT
2xOe4TIDdjEg5MuW6ZlxvxGEPQUtn52wkkN+MMs+XRzzcorHU5bKAhKluF+Z+1ZfIepeRWbkQ3cJ
QSzWaqYJxzTOASjuqSExogIdpnDWdPtetD3UPiR2ExEs1DitC1gky6AUMH1DVMRDJRlvd7zLfqx/
tQFmPY0lyRX9Y9PdYIBYXolhPoXjxU86GO2o/MaPnV+h7ti/Xt4FOi9XZWsMCHX2+OxBBvgYVY9x
4qlzxYDOkxHJXlzTBqP6dVEU7hd5Y9GOm2ZRN0Ks1N8pelss/26JN0zvfNI2qkVCIKf2qxpLM8bX
aXUtplogPEPqWuJSnQTKAYK57U0xbti7qPb6G5XxI5squpmh7T8RkOoLvATJ2IB9m3JSpezPeRpc
NPd0fTvkynSO5lCv/fNdDvkn1qZNEpq+8FhTz2yrvNL+W80TP+F0+KxFcRvj4XUv2dgJSGSbf4++
u5F20tgWyF2+z+5U6ECqt5k/CzItJyFFGcCnaZ5xapcd6DK2VqZRnpBtMi9pOO/KxftxkfmEfI7O
9Yl2b6QVEgIQKQOIblh4i7DAklN5LDjiNbhaZ2ilTQkLAYJNmfMUneDDxzUrra15HDdH9CRJ+WB7
Z/wOwTSENBdPD43vdor4VZ/xK2/vTgMwg8006VavGXB8lReUsPiSt5Sjl5EJUm4o2wdpDJ6nQf6H
vBS/QTpQ0oH5HcTnTNZ+O8usSC2TlJsKZERhtxSbFLWTULHfeVYnUHWB0Pk65tQkJD45psEHJUfx
4uRFLTWTwrcBPvHL+7NZDokwO6Y39YXWM74ffmoM4hXbv+K2jOU07bal5Ibqupb/lUEdJwh2KaOG
aUwwoWQN1nR35DEMN3w/KJemUWkE8fHlS3Dl+6bWjK5tn3a9jpBlHvOngJa84nixyk2avrMS9/co
DjORL2u28Ufqh04T8qKtg2pI1cHf/lLH69WDdQ0AN4HZliawUlxGYlndWUsEqeemAXdpEslpb1fW
cfYAYoBLEXEJva+N+DgJoyZqzIgRbNNNc3M7LnXGKx8wqcRqpEKOfRtBeWLaiKafXRo5g0Ha5LVI
hy/CwREp6eW7qGNIef0tGwoqzfgjTZwqlMnkn+E0l2Ap/turPzKkS+p8GxqqFlBhQZg2N1VQ5+ZR
TgGmwvc/XxzkDewHRlDFWNmHJg6AG5E6kcbMNplOLs65NsAqy3zytIRVTDfPmGsHwwZKRBw3WCWp
d9DrSe1+JmuwGPyTPXSBwubQW0G39R+Drk/xGzZQf77BbNbFY3ugkUYzk2bwf11ZibSw4704ik1T
Q7n3jnn4KzuJUxPIV1l8ByMT8/5U7BKq6lSOh5vG7g1yCOyqBnaNN4KUuVy5hk4qmASct2IByMjO
3Miqz1lneN7HtpLnFkyPUzVRWGAiyjf09G97+muHmLOMZuVz/9t4DBE3zLLPFMT8xGXomuV2crqZ
5fslyn4BIu7KsRgNwEGv0BPMaRoVXl0h/AtOuaXjcbnsuL1Ds8GR6QxkAjH/cqh6kaFP/RMGF1wM
Gdrfoq0a+Gx1y3d+d+UJoW4JkKhFafB87vslzWUFWQnX2ZwqEfQ7MEtgPLboXu8cWhttG0VC+tPA
m5d65KwwAusmR57CVhpFxVdcM2IpUbugtgowKfMcz6kP2U3Jj0DQu2RECDj5h454wsr2euJkS7sb
7dJ06Rr7DhyLXtKUwzMYD9MIdFB9UIg0Ol5xC2rGoT+/REDemRvWYtaibV5bhyGC9pt7CqQBmoQq
nwLedPT0NJ3J3LzSbhcClMp6/HSaFyDMTKZ3cLaxMqPKlKhSHVO4nKix6O/epEJGMmzYLJs18S1C
ngvArYtdeKW8841GpUcvyn9KtpnXcNLzpKNXnyIpIiwyAUIFK5BxPP/2Xh6xkkpu2pygEUJs7trh
n3eZoM/O+KU05mmoFJf63sMONexXF+EbIljFNTNTZTCnw/S3wKEvIQRDTBPYLNYSSIC90/JwdPAl
iakw3JLdSbOrHXLHyLD07gjZAEJctTqQF3b4e4yWUCtZdt08dTesC4EfryYgA9+OohYwS8k89VBf
31OpFHYtHQ+/7OPEFSuOCp2riTQF6ewCosxudieIEUBuVjSt2q50QQTXJA7q1KX4u9gke2jQIAkK
jCzUkKABEhnzjtEWHWjlumYZoIuEO/0S406Y8yB4q+2cvheKTG59ipbQp1lhh4ALvtWklt+wL0/V
MI8tFmCcZS4fPjpt+PMYz42v6eY7ufqIHiUHMti/ydMdPWiMmHMDnrWx1v5mf6r9huCxROl/c2qj
beMJW2mFQ2dzV4g9xOdl/NWHG74jDQc5W/aUdjQxEomNsV9yWdEQK45iC9ekgTFdIanRrfmLNcsX
4vJF0v7vlN0QVhOqCmgR8uYqu7wE9r8ctMzw1TqPzFrXma8C0dJy7QIxxdjI9d3EhEF0SBP8pulb
i6crmrvdDq+mUXW15jZqbxc/d3w+89Aa0eA6V9nC81VabpNgQfQybIGFYuiKU8Ugz0+TJTbfBX6M
gGXA4sEpfl3hUJpvVOyuxRaX4L6oINEgP3EkqC0uTzMx3XpSk8ihfSzw1PdCt371ya069bHB3Oli
pvqTRURXLzXn8YRZ3K6s3Jy/co2Gr+5VHS2RiRcgm8z1Z9naQVi+hs4aB2L7fCT903h/IKEsDBP2
Pa/e+ypaYx2mlMze+fjGYG98Yl28jUi9ZrTH7LoUdV20ybsziu+4ij9dbAiV/PKvK/OVrdKpUW4J
gJokWVooVxWjp4VKJb7eVbtZhodyTLK9Y671JbZerQ7sQyAV00Thpwp8QI5N7L/0EHrymG7y+5Wa
IZ1/2LzMSGW9VzOS5ly1cIuajQazAiwBuIOw9pegCsN8ih9h0fHxjYHSnvouGWtX3BkNuOwjvdhi
Cm4gcg/UtBNSyhxAIbhqXpFBiDUEtDcZa57bG9Ww1GzchVW+WE2CcFI6l/WBpCa6fsi89eIr4okZ
hOvjGyiVj7kZjP69d/C0LJ3meAcph4rGONWFnhGTVGKzaNor0LAb2frpbt0rnQHt/wyE1wFLnwRn
RmCnbTqvIqoppzdxN00TabAh+GcpYo9Bdl2J99BhI8JPG6KppLMRhmUa9WjDGSu/cREUOtjEsfak
uRK/eMsoIfsaugTG5D+8ytf+qwhXiEsAF/Oyzo4pL+mbsFr/M/7IX/cUFBfwH8SejfRRbkR3Ys3j
CrK8iXclhPgM9O+kWjP96ASAAan4sDyYVn61B6jIswUYntCbPJM+qCFsKGrK+6R/YSdOjCiyFz5V
uZdDDwQOG/rkj4/Fea5BKByp6Rp+5e2g3AXIKelnIj+08wfK7BO589lRCT4EjG/fmDHJaWsii/3t
ltV9maqvYjzkDN6/sSwYju9aE4aLozw4BpqvtnrPtlY+GilyBoc1rPSrR5967BNB4MUSF7CDvErq
ehaOCUOpqu7C36LXBixF9QQtUKr+NLfaziMR6F0+MBZpAsVqqQSvuv2Ms/zTOPAskl1NKOeBo0BM
RS6r+1ppSr15RsrHgNRNGuapACvIw6X4YRP4TcORa7fdOQjx2qJokf4tZwxQNP4SSdaZJtXZ4edl
dXv4Ye+24u9PT/yvcVXGwzhFixcYtihqEl+8bXjLHPQk2yenpkd7tLpa0LBKfbDhDVe7N/WKkJ4N
smGHFe3csQAKpqxOHpOxZopOPWElif0TeUGJlFUeDZerMW8NY5bl9H+Wmto5jAjX9XakWHYkMpFh
8Cv5G7XKvZi13dsvyp0pgjtqS+UjyCo+TTArefmOgfqKUXh+gFzp4/r9+RLONrR3GPuHSDMMf8BE
EbRtb4SEjbL4/4sFE9JzR48C5zcl+Bf62nxYEkjZLR/xpNDUGgDuDsCO8vRKvIWWXyF7F7vzUAni
OYYtl1XdYFlWJ9AnKyAzwC6jCXIBkBQkTSWrg5RAex7SuIIBcRyX5rtWlVz1aZjatl7IPG6XouUp
ij8X2w9ECuvdXVu8sEVMXb5aPgh7QZ5L16l+DmpmhsxuaAGHO0CHQ6Fz+NBBg6azJG9M2C39lsZE
DW+0ZIEhQjk0hnAZKcpVpynZgRr+GGzYuJ+IpAHaoMGD28BxDRJz/f8hnX6f+UpSXTp2BO84miXo
jPwsHSV8dFWeum22q3JPpy748gwLB3nxJA0cTHYTib5o7vth/jZlKHTvzWpYE0Y7GqiLJACVQxtM
95HCGdWEPJb44otZAUST3wQdkduIImI55E+cJ7OXVgzft+/DW+qXvgzZia//BXVu4GUh19bO7ao2
x1lPjOKBYAK5Zl19jJwtSKS5MFrvZaj07mIbbqGJoF3zfRxlo4xU21vyUwsm8Nq2eIThWFg16UHm
57kkNVngmACXmEXW+J7TEoUEP7Ts4LPAx9Mt0lDgcvpHm9SniKtsWMMs1h5EA4Ex0uZgMBVa4IFN
wrx3+azpzjEwpmTIJggI3744ByJOxar5YkLj+D1Uo8j66gKWn7q6b124vEEHG7RveE2KrYXIvUiQ
UEQEVOLA2Lj3F0do/unQshgdahr4n5Yjuc+2MpCvF9S6YawHPE44Oj0jxiwygJTM6sy+zKuFizFo
l8s9UaCM1nq4+UNrL5dPfpSwY9zvlR7U6ZAXdVfaUnbDw1Xgsvsl6ayhyhFL7mKveO/TnjdiIeRa
ZzdNzkknyXBCppH1Oc4yQfA+8yDqibxd3nsj/xfze7UAFaf6H7ztdCOFBXC0y4BV+P1Cs4z4m/zD
efMcQWKcF1zvIzwozdF9xbz+GX9QjdSoQHz3Xu0H8cjexEMWhcTRVnsgRcjrcE2ki78TFURRbc50
R/h7b/5MiE5CVIBU175xFKxWHJJC8PWN07Ck3Y4vlEZsw0q9dh/fVzwn2x/vn3Z7z+UYVwaxO/Jy
9m32+Y0fw0hz62GBQMKG7I/tMwAghTlTtq5gK31wmaYukOYDiQouChxvP919lgnK12nY5wXP7nle
o5Cq2Aw4Qeqfos1nh/FVBPl/5KFXPL0h2uTWbLpOa9mQZKDGqEYb3GujaJgHhov6RXogq2n2Pzut
KAxoABxPUe+UuMFeRJgcvmxYYngI5LlXGX8KsQ/QxLf2aC0fQgOAuV4GBogXxtMNrnPnKvggCVfs
QmqH/zhCvuYp51ujAyJfx0QJBoKfMK8BYqfsLwZWjijiCUHB8wWgI9o4hIuJp4GYAFP1hm93i8QB
RMboQsU7HnSG6p5vDwarqfAD94As7lHizq4SM8BWXQ6ETpPVOL9jjsOjNARmSHImGbox5k6V+5DT
c59p8TB9A8Ir2JkSh3b/uPavhOjY0zBOKfc/Qz2hM67doFtu7TLWteRnXQaeFaQHPgcr3/NC0udq
QPHkkVR3Sr9XeGmKfJ89GZ8pu8BmJddb+lCxHV/xtjy+StKse/7N6NN4hB7mRs5afmcakHgumGZd
AMpk8QNDAjeDp9uY9Uzm1LtHA96N+p7KFSezgnWjBGAio5oYSbu2iCd+yWeRF80/xRg6aZjTLR20
2DiHDdXiHAluE1TKnFwIThCO7P8gCFRZpT6lMn8FaDrRwKHS6A0DlPeDsgmtdsDbtBL4EXoo9cm1
4Qj58eF0dwYyIq5f65kriF7R61v2HUnW7yLwLVKseUdVQY1vrqIx7C+sdSpAbTZyiEu+Upj5vbeY
kQYnCRpH/3v/lWWyODmMYsDAYSp6/uOS3kRQvEc4ARzFG1zUe2ZD8UfOQUgzJoNr8gJ3EHCBZwCf
zClEpzSm435XXmUqBDKgKq3J0bEx1iS58RLa9F/pmU3ELVUybmUIyinQHddnaKAZEuFNgzTjx8JI
NAY2/vq4tw==
`protect end_protected
