-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ZVoitIvRCjRf1i4KS9nBN2NMlx+GlCSvQKW0GGUw2g/zNaVQvW6MSak+dV9vowxC
uHH/c5uuA49gHDNDdOhBAzgBG3YqbC9nUKv3PIabNagjSRvVd3gV9AjvdliRRjCn
8Y5AU9Dll67JfyhPWMzTx53t9XRSvCsB/F8PQYQJa4c=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 69584)
`protect data_block
WumfMA6/Kvk51iJepRxQfdf4OZ72VRBRqGradtDxgTtbj2tPhflssvU/GGzuC1Nx
vkPuUNlyonImRYO4l+Kn4AmauMfT0XiXv9+XdRwtqxKh0RsHf7QTVVfL0ZCLXrKY
zNwG0glWjD4KvP3p8lbcB4JTIV5lMxwqDJ4ZZJ/QmD6Kr7lGpRerhq+klcDJazKG
PGDTW359UmuO1GAJXMaqTycs0wJh7hGaaxv66rQA8VXRQz79KeZ7emEVG648KIJI
0c3qO4h8briEY47QGdIYvSrexda+dKgyjgcdSgp07sMAoCnOo8IuFlRq+ruGlMos
VNexibM+40BnbbNdqB3dINGOKk66UlM6rb+cSl4DMjDWum0l1rj74roA8e8XXZPL
+rCZj6OGvXOP7m9igfM889e77h/59RhJNmWZeCXygGmCBNkuvvJ9/gqVD+Ey+hqS
JB7aYyIvJtaryrmg/q1dya6bpuNDpc+ZJaSJ4io1E8gGfdco4lt/RC6zAY3B1HMz
okqZwgFO6seLOrg3/cSX6sBa/aB0fRiuKX32FQfL4RqHY7b+x4e6PxXY97UVBxaW
SS2C/LvYrjlUqcdO2FlN+oU+399v0CKtunxnV1ISDu92pBdskuL0XTzRGqJ/uieR
nfmnugnbD4rk82HtdnKOAthwpx5gjiQPpSmbx614OsQtDuh8/SqXsblpEdimmZqO
b+NwBmVYKwZh+yC0tZxAx+goytPo6adA0u1szMghgIUF5S3e8M36CkfYKRCYhHoV
N6VJ24gjPHrFh47KrkuucI3VocWsTLi3FRMScBaO9bLsqOVYe31YF+KS2q7dqkYl
DOAsKrrVUhl2OYG6b+STXS03sysSntettTxmUz3BVfQasYt/cO+jUGanvnVvCWy+
leMbBqj5yf2Hob2EMbdsbeAanpfCWWfYvEtuVRvFSG/ETLiWFQkIWSq4vUTk04qz
cdsf17Dg+nJXqOPJE1GHtYvL4AgD8LfyPxBR2c6T6ZipvS08guwFRAjKmiLgWd9l
aaP/YndHxi2dmY0lb9cHvHhmf+a4f9kGtJpr3Kgt481bxbFIOPTsAT1+LTkRTF7a
V7CY9QB7a7sE0XE7b0JY6hXQk6HLJkm4/7IaFJvYm3wcZ+xp5cHBoRvWlkyWKoM4
u152sRnhyeTf6MRk3MQTPC4vyNlt02tQXOGBSF7f/JCe1df9AoN1V2fkn/LjoTFv
RInHeCWyVWujuLCB2IbFsrdrEb2fIi6SWN5qto/jIB6b4STs6WaY57NRB0SYRVzf
hSjSxJYUY9KC2Eeg04EbNVb1ekmSgSk4A77KU77GNXRDAplYhbB2Bh4X9cqLp5TM
3YLw9MnfElQBaZ9OLdcofQyKl6VjIai2fXiIaEymEHMT7ptvoke4GqOsYfyGdGa7
VhcptA6FI4NFZDixPlYTF+btqSChw1qNQz60YkeSkmHlCACDjX7tVwsTaWQ6srsE
8S0QiVrYVIdPpDDs0Y7TlzKfuMdab/mj5feXzre96kAhwrEgQMKz/iAauB+mUmKo
dc96wP5boOyR/0ZMSVdSJRYM0vliwZ5yw7vwrnEl/oQkq9+aT/cm+vnWAJRdHtLW
ry/fRbYgr7/zMWBO6iFXP6UiCoXUBrpGMxYjNvOGjudEvxLyGHzBphRS0aoRBkVJ
3iWS3U9azfdxAsZFuChomppLwHgK45PpAa+/sNnm+Vvq+wVvf0pUzD3l5RbnOPH1
zcAtkYzIIB7FBKU9mJtQG6ngyY7+MCn7u0t3lu51fHrANMunZM8W7JtEW5mvKWT9
jAnq0AN21f3YdWsvftxGrj9zgODJeRrTmcsLGW/BmvoH5xwQwNbSawR6wdvuUJXV
T7YLgt0rEwX/mSxy6j4aH/oczqAMS4gHAhbHQlV05+Cw5LvgYf41Zph9xtvvkVlF
CpCZFMONAwVu3+wYZlNkwmy2ymlQwdRdOF/CfsgaRKrlAGAFJVcvLA22u1UwOaaz
KToYUBUA4UHbGONc2NL3xOFOSnHXQAXiDJzNTOIVAtyVNqTCJt2iOTY+0XAc6YBk
Uq9/qKNX/RyErXSE7b0lQJq1tNuJGZkXsEAyMK37pD2ESc9csdttyIXO503JSzR5
Ji5XkrGP4LlziGM9+SMlVjwgSVPZ3frrpOnTxLilk3IFb4s3r4RRagjf0+GGdBmk
iUhLuFNiN6v1yVz5pzCRfYSGENnXZq6v9Lw1ehWa88gH832HmXHlP0DDLg+KvmaS
EbWc0R1diHeQ4Z5QgOjL0qa093VBYf2kzltqDktz43ms7MMlHQlEVv382/axL0Wm
I46nhWNjSwa+EvMMrU5r9yzA/vx6WsoPi7a0uK17JQbrLrxg73I1PxVny8y+BUgI
0+2Ps0PsI4B9lnfeN4xl6Sf+ViOnx3h9JAelAO1CZOGcM3OOqVHueNIkVgrAtj8y
QWHgz8TJsNJt82BagohQAHNeH9T4R1vjpSUdo3f/gG7R8i7Uh7z8goGcevBtRAoZ
9UuZPjicBbuqqDwJ5eEMZpjLduQhOHRzw1O239K+zLILVQfVyL1/sVX0FxhsiGd7
jpzWPWgZZAx0sBJF4wnj9DckEU0bmCMB2pEW8J8Wz9sMYTCPCF6ZHueEEv82VsMC
CazpDkB6xTTCkMgh6pflHVJJBGrowjjZrlzv+yHmYBeeDfXzckT+3msyd76uEqG2
lRKuHBZp7gAWZ/7II85OAyhSVEvxn5T6/WL7Vwble1p9U2gbDd133s3fbSWD07/K
upfFAoaJzP30abs0c06PcNU1UpQapFhrl9VdJga3yrrD8oTYVkzTO+tYpCmy2cuv
5p3FAIVJJagKzydhPgvXZC0HZk+oMkI/5aoaRJ/TL1+Gh9JvUHoROExorwNRQxv4
jxq5R3A6xdSTTHHDt5dLhGy/0gaHm2PrDVx5bmrJ9iQ3rLrCSMmaxkyymkgOTYXU
Z/NCwVo7BPyjEja3ZiQKoJBy4sr9BPthzPo1q/1/4Jb/WtmHWmltnXssXO+Bl22x
XiY165wOqFDjcWrS3Ts8PNhPS5M8dHEjYazqNHNxj+kXzErJ6y0e6pmrvEWNWf1E
YdP7/VbaKXp6a29OIOvtzwM1MLaxY1823BcgvTeBi0G11YB1ZfuD1qMi3IO92Qfl
EpIA3XAkwiKagXeWTU4eEDznAzTnfMb85fHVvVRDg5z4DDfC9lut/+cvMiwJEPKO
UBiEIwyUlhy1Q5hvU+RG7XMt1d9HSFUmmMER7qUv95d5DrXDbavQ+o5jE8ZL5fqS
kU0Qgdh2M60Gh2535+uwIR1iCafbBS3D8qedg9/t6oq2N/a4zMXPqcBJlaILHSCc
qjbgg/Qml0vftBKCyYNPG+ir9a7hDzGAZPd0xqEHSz5Nf5yp4IIs5GaBmHqZw5HT
bEp7rArD4NsNGb3Qaei6pqhz2fmnWvgefhdqP+jwAB8n6B+LffJ3daLeJeT3gcZb
jaa9WORfUH597hCyVODjqzZ8AfGKH+rXmTNkRzQwkJiP+I/7gXmpF4NymaqQOcWG
l93jDXgNv9tC3M0FJCWX2RBbf/LvxEj/zAFVhexG1Mn+lxlbMigUzBAwkWHV6mEr
4kcn0O1/BewNAB5PSOic8RZ3FSb8eBwsP2trW273ZMPdKt2dg6NvLhhAT+JUzc22
LhQC9sx6M/L4hPC45wLxrbe+rsskeKqixCwShLdJltF4miW2dzVTXC/JjYGCzy0M
4E1E0KTisFd1u8YgjEgUH97o9gj/UOT9gCgYMH8Nvn46sAmF9zirKlllxWsJCWeB
KtXh6Ix5ITUP6bEMxmsW5b1Z3ubCBeSPedgflkO4Xnv59Mxz1NNFTf7TeDFCXgTN
BRJqRrOF1BA+bOtrIInfjxgcPWdrXPmSEyr4QZVnq7n//3Lves9XxpuunRsus0Fs
4poZWDxNCMVphmwWF0+ddcxGJJ/ZUTBXuITaVUScjUCn2QOilGjTj1KxKZJVxjPM
FR1PGfIkjOT02isp3prU5h5C28/LsGkt24Yxtz5wKKzdVxG00LWpIgd0vYMIedvO
5ZllGuOq/3DWww/uHVGAWByaNdA1OdvS1X3BNTH8mmQeg2HPyRj/eSdSX/k0psl2
Cs+uzvnFThVuOdWEqRFTh6TCmslzf9wiZzcG8z6/CCsSdqYqu5Ky8FAA9MrLtfwV
AepH0ULKONBJ3kdc+sd4OVypu4jR6VeCMjiB7jDZI2ocZKLe4rtzFAXf4LSaVF/D
bjA00LpD7dNZTe65Uw4CxWYhtb4zaKBwBY60B+oJxGDPAZN0Zo6GwITXvMl3Q9Ht
oCRHuTd8Wct9aXjpu8eMN3w/5o7ee/ws4j8ovYZKywgevFZp9k2wPXhdWR1lK4dp
VV3mMO4hB06IuNK4k3ubOXzsezGoljn6uQZUD+tEqmi9HSlR/KN5v/iBIL/NCTIC
D/6P1udwuMMfjiVHxqlqMF0MWdhSt1Ti21hGNo72wRlSMSFPLszz1JKGZrIU09jq
7bWLKz48uc6cR7qGZsCqzncJuA2MIv6ofn8+oFuUN8hf6UHXapMZcTAX9kB1m0RS
PUTjb6C1l1jPHwy9KeBRcczobqzdJYgKFKooCWxOt3oMZeTQVEBNHDG57P60Uily
+gTjfBGqWnO1gt/UPKqiypEhSig/9yxNkWc2gHdXSmao2VnpQUvU4VNGHy2W3jji
cXiqd1TjtCS/a0XJSYY2HahPiUadQahK4yOjZxQ/Vab+RmuIzisQUWx1KlIZosxz
8pCp+YP59vSX+KLOPJ23WrNl7UV2Jc8aXoCinTTn7+7gcswOaEXruqpK//BDqjiR
I+CcVF8oDI3/RzymHDTOokWljPyVQW1W739/3DmhppquHik2h6ZagHgZO5tSF7AH
s/3c5IHCKphg1MBGnI716nB9fMmLvCG93ra+owOI6EqDL2zfF1y8EsR8fAWmTTwA
PPZIzjs2Gy42etCAhmVueM36IOxpBsxwbj4OMPUahJVVYCpcau45cY6CULe0JKjj
4FWkjEekjLSq5FbGfiR/XRggAQ4kKWwfbM1ay3tssSq3umelonFcmQyelNqwGE67
hWWkJgcqyBrCc6FSU7yElqz/AJ8T64yeoqqgFxL6lihsliN53mpAlhq6CeM493K7
dqGgxuAsJvyVSNCMeMV9mW0pY0ml6nUZ7Fx2IwR2DR6wQPRImL+By79F3GnzwZJW
pPy1ebAjJTZWWscdOif+y5ppZa3Hs6atumN4YeBFrqJ8kMRd9XDmHNJReurA4O7e
UffQeEZtlBnNMQdLvkLI/Y1Hx1Q/tpbepYo1eNGMtoVEeFrxSLr6MYpcc6Lo3fSp
QAaLhjZ5aXh+DAfMBaPh+D1AbcptCJI7VoTJDW00V4jI6Szp6/qYwMnf0t3ZzjTV
FKjE6+TllkQtB+WSDr7uIiUMbbuMJQpu8fpYPDe5qdBdt9e9CD6gWWmE8EHIboPs
phRFqwi/Jd7YIFVJfmS8kAf50fe5S5X3Q5kLoadUWegctHG+k3YEgAvbsNwNuCTs
4tdqjoRSzSR6CLCm+O+fV9rsf75w+m8r88bgn2/ipT+AC4P62KPZL2v/QsUey3jb
4gSL8NExW5pLEa/jDabdwI0Mj+i3XfgHPh/LDOokGWZCsKvc3tQ4EZJHNMM5YbDK
bgkTnPN8UpRVWSwviyhCwMz7G8VaErkl8S8ZA5OpfcUs8cQIdVMcYz5Zh4j4Oc4U
Q3qsjcnR+xXXwDtftF9Ucodb9QsrvLvOl6RQVzVpGI/ZB5V4Q6rxzc/6W86Hu7jw
A6W254lT7EUy3La5qL6x32lq7mHfllJ4e8ShP3OpHBZ70xxavpOAYVXMX1SHsZRC
cCXmNqsa/vQrhUgrKmK+RTCkv3umh//qWQTNHgq1fI3rpnHpAipkKqUjpQyjy2Pq
JeGAl/XcuHzq90JbgLg/a0m0ZjsOplRntBzybZ8DSobFrnCvOkFn5X44mHtTEMYZ
FDrqRVW+gl6ji0wdaxl94Tif3uYAjVs5h+EfmLKNsC0RrHxwngSvRdb/rBb0/eYS
+XcFdUAwNiH4U8RoSb0ofKPk0uc9Uoblom4gZTL3uZbybcOYeGfdPOuaKVGnwJJd
wF6ctPz7lK0Sm9kLGfJDfcwTOvzAwAR1Wk1RBuiAJEqG7LMsQfa9LKYrf40Hgs7D
ut+elDKiyw+aiw4y6X6OQd2Zv6onT8k68HaCgPKbzdhcfFQxMx6Z0qTp2RjoJi3j
IOm8C566pXk/O2midesXK3PJqUAsdfoilby2+Nml6P9EE88I+ad0IuNxJ/WrUakX
031vpTFLQYGYYbqcATsyb/Q8G1l9up9tCM+oDP9AX2n9iZ/aL2uFoOyr8fUXNj9I
GeO9FLxIgSMOWx47wBlIEDUrZVhSliRvb60S6aSkIWBsWEXFStYDhSHqRZpGZu0M
JZqA0Z+4Yql8E2TFXZV8GMCVvaM2JQsB+eG5DHnnLJ6jfcZl9GgOxiknWdcyqjqK
2w51xGMKZ6P2QNG4iZYzLoRYX3/PaxETbgt5mR66D9hJ/gjFe01Di9xTjRfPHuIJ
VKYNKMGdrassZNarHHkvy9aLfEjztzbCbgSidVDH7cu76w1s7qVtavhiEb/YXzNz
Q+GCVvDLKCmtlIAyXGtxIESB9xAFvLJ67gkBjbrLn9zWIrehwEvau8rEISu6YdA/
INIXzunkeqW/SJTmUTBhfQG7rx0VKC/a5gTigXStFiBDODpPE2yhex7UGjnkPJXx
WokP+E2zhUjQ2cGOc343h+46UD8ONQVLlWQ5G4mZedrQvorxYVNLo3w7gfKLRdy5
1G7P60DhDLMmUM15F01QGtOJHIZnzIIJzr0x2h6fRRpKwlz3wYZmIS+VyGyWtQSu
F4Nxeue+FFDRX7eagKjkuv26bs27zPYIQVcnvAfgJxC9jEej6wNkFUlNyChPc2Pd
5PE2Rmm0NLlZUNeXiBgxIXpIhtMiWivN3nXV6kEBkkqQ+RkB9zf+vJqoUVftA21G
Gt53KD2nWXwF9T52ZMlK9+paa0jVvyhMjlfSoEcVteZk1GxZonbjkcNOC/4Vb6Hf
CS3z4uTa3KKZdBeSVamWd2iwLeArU2V+0gx2BC1BXrQ+wUGonstWtLajgP4iCV7g
MeM9iMeVJ7e+S5xjPnF8iGM+zTutZF552CWsbUPPC94onS9HKPscnN618x/4EC51
aK0Mxqrg6lD4/SGXaSQ6/vASHab/L/C6XoAsXdfVr1K9uygpH0C8YBvSW0ym1f2D
Nhcxlm9uNFfkNts77vWbzoIr6NGkcczqsGnvXNOfEydyqtVHPPU1xh/Rsyr2OKHe
4xkTSgjJ/WU17mlH4HknmianmU/pT7Vsf5EG8l1gR+QUc/nhNKf1//abBo26CzrG
NaQoItmHI915GChuDDu1BZel2QH7RfDk34mpI6T+DXaSNyxT5Hn9t0+jjD47aw0s
Jgi8UF49QHLR53TA5p3gewRuC3NsbPVN1jnxPZVryBBSz/ivj1lpnZI5SyiJXzQ0
E15hVj4RKkf0ZmVnV+Hn+a+/63/rIsuSpQqTEbNOZVNivErQ4DCFrmERpfqSXBj5
zsb6rRVmHn7uYa9aKin39J5WCRcO01UpWqEI9j7BCf8lDmyoitrF7LSvXQ0azLsG
WWASgg7L1HlZ4IlULJpVXBhDUh3EQKrYbANt8pbyexYA7h4s9uEuU8tK8wlr3P39
NZoQwgBOgv4d6kHhkvTJxDcx19K2DWRiSl0W6j5Cg0+FvX9dTsJVDwwHMEFSikNI
C7Iw3iAStlyjwpf9up6olj9D0ZBbgnfn3jZmiy1LB40LYDtk9NURA9BqVtj9A/Qc
Fg9qQyCmqmMZx+SrXqzoJLhxqNHHjEBPDYFMvP9cVcohUunmeROyQsqHQRHKqrWy
2GYMpUmX9IC25pxZI0D1AwTx6UK1ckpk522UF2lsbhSHntl4OXpVIHkCRKcL5M8C
ZRdbuQaDVRuY6SeTl9pwgkw8ZdXUDh8Mcw73tmQOFeTo6VT1Lx8wWICaPbXqcZFZ
RaV68bfyCWJLqVySL7WFzRnnJn0oUxdanXroR1Ze9JlOSNY5lxTq98OJcLKLYHk6
qHEpnH6RA824yUFWzmOJGh7xdtEFOA8i4qSG7oWBz1/2f/AtLqaF9nAMBDKPAzDj
e9VoODcrP7UoeoMFWR68kBXc6idvKlaLAXENHDQlVhnRhKRoTCJNGjE8Nw4zlrgK
gqd5K5WsbNiPth8o4FgIfezi1WWNcn+Pxt5d0PZ7Dn7I1ajxUBldXTjiFH5cEmi+
FfwwQxTBwmgo7aFkVLbY69WFLrR1yeTnsDxXcKHkXi4wEIX4+RtQ+cSnl+BDhhOq
Ej4jQO1864tYw87hTzZKIXc+EAKb1lmUV3s/qCjwhw1ClglA+xjn7TgsnYrtgGzC
VPAc/rxPQZvGX683f5KHFqYlGBcs+APCh/oSTx/TRDeScQAFEdAmGPVcLpAGxA0M
DXOM5EO6m1JxwpZ92oj4KEhVA1OliiLFEExuE51IG5ytGaD2XRUeIEzPK+G42YCb
xNHXCC+Qp6m7dYRybj2XHvUZaStflgVY5W3FjGAv4l1gOsxscAvlN8X0ZPPNF6DW
A36rrModfaOGdwZnhRT1LGqrwvMgW1UDv95GS01XO9bEsHzyuohXo1ZSX8GHkrru
gMZktBvb68GMqA/bE7JG4TMzBjunTZdLLph4YGUY5ZnEYdiHi2u4wMqUOLSSA5z2
uKkyqo/ug9nvtRQhrfKOLGQMqVzFEYch2/7lP5xoZzbOMjUEuZczOoIjLpMpjVev
bWgY/3NnGR2KwNcxOpwpFR9l66qCjegpqvjLy77Bcy4mRQGHRCku4d/IXTJnQgUp
B1DO4g2Kipw+xYujIeVT+moqGhR38t9Vv8Cmp/3xwClNXT35Q0EC04cWrmME9fmb
W746Idlg+SVE1Y7Q3QVoo/cLxagUJk5l33oklkRem4nuEOVQwN/FKm+V3MeoiAWi
h3+I4a7HAsRuJ6D7r8CYjcZGA38klmAn5v/8jWalY6MrIw8QRItVYcyeSNlUSy9Z
m3R7MeuyW5E0geW+VRL9DtdmoroVts6FnuYCvRiaAFT7iGNKl89mlvJKVkmQiDA1
UA8oeNzUBu+LvTPbrmG3X5UJkMfWvLCYSYU7agBiSdozAP68v9VbFxXR7vLnlvjy
e6CaD9CoBDhRUg40Y5S3N8Ms9ieKEpkcrZjiWRwkDlXj04uwV4/V6GGNCa0VDRp9
sASrBxTQ0WCp+oweM0zdIqxx1Q3MZfybCyyWKQH4rUyXmPU8j04pPj6B2SgdA4Uq
+MIGuJ71DbWL+5I/IuDaysCsVnIcjEOhL/SJXTKtAn87SOCwsPl/oCOd4qRPNK4P
f2xwCsQ5aOYFAvqh7QCakGEs/pxUm233zrDWQ4VbATHhHhDfF29As6MCS9ZD9H76
tV1O8ZUOO9l6JTEGcu4qju/hm+irT+yjzItEffS6JezRpjXuZLhIARS9pJa6mda7
G7bdWEMVhIzZ4YvYqaVAYdLOgztlZ5ZQy3rzaUdSIb3cw8jsMuDdeSRx+keHVAXk
GpqNF/zc0ADOAZTlolMtm1fGD9LU8eFcccjf3Yr9jqlgwE/24cLP+qPw9zpIEBnZ
m0Y85mteSHuj58mGkuOyqPj/I7c/SpIMGKUonizz9EpWz8w8PjgRhW5Pz7lDkE+s
8lvdi9IQQShJ1Yj3uYbZHgDEcYtrKSJGmgkyiUa/9+ja6Hqrcr/mq+TS9mJ18otH
K8ALmcYXYqkjV6U0WisCalckQ0oUuio3AwwCtadV/u0CMG8JFmhyWBI9vZ3V4PbR
CL9VSl4re84erUQ8nyuIXcdUWhWeHYNbNNzVkHzgWZViC6Qg+TCxQz2o5Do2r+pz
+tzGt0bI1Mi1t5qcKriYXnuX1N+wk94NDk1hMDrQlV+9DwibXTfoZkVN0zFokjbe
s0zLTH5FwX02dWYFExaVbGbuK5flhrDy8gsqcAtREYAD0QFAngGWT97mpva0NXTS
tG2ma3xRUkVZqXCeLH9qiXc4RcVvu8RxDV1f/HA45dlT6FnJj799PLWR1tyhWm89
glqTEdpgn4PwhKTsvRqlUaqfW5rPazT7eJTQXc9EQr+TULwNvQ4w+6522tdrv0JH
dTI81minjaPeJ2zitf+zQkIhjndnR8CiCUs91Bozr1EGsL+PaoBAddicCxlHFLC3
sqGLxYzoPpRbVhTohviOCWXQIA6SsUX9hHaj1xBFoBNRdmP0z4lfRf6ydmQGAQul
WfwhZp+4yYKDBH5HJcSQWGur7lQI3wPmkbMx2P+ykWdnsep1nvXBpvrsZo1pSnVJ
fhyJ+GWKhtEHd8y+2cXIfIDYg8ezMlHETw5+df02Y+4H7TulKsJa5fH3lM8gC0IA
N5I/97CQg1hvHZKIWPmBCXn8wTRzrEquq/4YenVVnlCQ4qF/I060IQ2CBG8LSJfQ
Unb/ZTtKsUTaSb3JI2o8L4EHLiwfBSkk1+tcG8tnz5mSgtyIBPrICTqY3yB5sOdX
H2Vy550YojYs8mu3DINFmpqox1ctM/2A3nKzJj4auqzdi+/3Sj6tRCohvCHqFLo6
dPmHOZOf+fOKOKIYJqVk1nFrOrq3PBT1ue3RUMW+IdXubU8GfUZNALsozhtuEQ3S
n1luYzECkaizjLCn1C/q9I10qOKefilpIEbjd8ZIm7w5vnJBsmCa21M7bb/rDc3C
1svOeMcB4WVQp8rua5PUrCPhTPomOZURaT/Q3Y3vPtWvkmXmzNymK20tQBnLB+tU
juvJyfdgAh+eHCf9P4w07pNWhxlAUfyezQa64K7IG92QfiJjWv9ppqmVvkTKqNeD
/RX7zCKdu40LOypLQS/1WmVPSfomUqRjbjcnMG/ewq1JJbIzXxGqllf9XVdCqNO6
eJr83uZKnUUWvR1hSMNqDi89dKLysW0E+ICxrwNiqw70Xb+X5veiHhYURmPHr/c2
5ltQVlpfWKS25Fe5tQQdsPmNBU+6KTN7dQ6nYxm8LnME6OO2sBR8/GXlvvtBGTVl
1CX2LD/9gsIeCCQ7qkV0MbsJ7dRAJI7T/q3P1lh4+k5h2t1BnDQ1LPLfCoddmzcP
2LdzIFS0T57yAFsB+Dwo+2RVSetJFv69ToWr40FaLiStEx4RL8e39wCC/CiPCMjy
xWfE93JgJIK1xU0RtH+N9FojvuL5ME6Q1lX8P0wbQeKpg3odJ4JwOJ3dC5JS2U8c
RhUJncjgCWztlLYJMgOYc4thomcZOy7sGYhmjcbBj3slJCwFlsJ7e0XVgPkKQHBj
pzVs3EVhEQb1tZdPQn25iKERWJuplTeWJy5rzKK5v8KVRwo4d8lpzn59TunkbMgY
WdX8HsVk3mhbeFiNqLEfU1/Aam5y9goPBjagFXdS9sNM6t4ejEv1RLcAXwGCTNgD
3pLXngj2xdABctQwtlTX/1G2FrXUWtFFACHiycN+woqjI2WudB/ncqte0AbteAfz
6o6PvfOs2N1FCn0cxtF81hDiiuMRjLNojiZIjWmkjzUlOpmP41aJAcyh/Jhm662k
e34fzu8tV+4YVIiOB9vITN+Njr1bX34sxYH66xhR32mUUaoaolUSordrxis8Rh/1
9Ksglp1AYxwxcdSPHUCu05xYGzi6+eZFvX8R8XRPfNbtLEtz67wRBu0vKRLatmf2
zDzzaZkjpvuXy9Gmf9jz27doQIM4aGE+FUAUFddvJzwJD4ELdgW9CHo0xjShHLcG
Tc98oiaRUdEGRVNUafgxQAL2hrHT307Omw2Tl3sPtvFsqCYMeYZKsCo8UFmDB7d9
WzmNwIG43J144BQI532m38qB6QDD26EsO0lMLzA2sH61j7u7v0lARGbiPvgisIB8
Y0zfhg0MtASNDXN0SHhjJsqdzDZgOlP4ogTnqgGFLh6vIlmScDzsgUBqKkv1nzSz
1UunoOhb7w7cLxhBE77PBukIhcvUeTuUS/Q3Cuov+lKgn50rjl5yE1iV5cRV+VET
F6oHnbp7X74v4LHWYEYimdxJlAM1Tit6JyG3B7hOEpOHnD2Riydn+HJFIQvI6N4f
qzaaoC0zmUnMe4HgWFY6tO9rKhY5mNalc+QLTm+JWfoj55eXPKO6Bc070TlfGuzo
TIqD/LBNysxzq6tlZb4BqweSSoygxPA0s+Is3HudcOFCj0TfKHN+/JWiCaOOOZmO
qEDHLPJyHrCIhrz2Vklg9bNDAvPjg8d8OeA/sBTL0fhI4uJZl1aF3DLbfqq9VeDW
KQBA0I31ye/Kwji4UlfCXlo6ahfMWBlA87NoENAJY4LZzo3ifsrj9yejt/kA4D1F
v1rtg0Ju1A4ZTMB+wOtxZzE0c3PPC0ikv+yeXqzm/zSl+h3hgKYyqLBkke3V/d5X
ir5UCXsBWmulfktBpH2IbE7/853qYfRBsWlQTVgF1kiTsIDK87dpsKAEGvodsEuW
Xp+/OIjQ4xBfad9XREhj2oGMwzsWsbV1DoQRytXisNC3WlJQZR695C9q9aBWL0Zj
F11OiWm/ObgrS3JZLWiL7vFOWxX13MVJhl4/Q3Lqo98dz8ylngE1Z7vAPK8FRly8
Q6MXKYElOUeLNdtEKjGqHOuxBG+TOvPf0fn5v7HtFQl9125UPG9AJwInB/QWG+m8
J5dW+3wizPpGvEbNvBYS+lb1FtppdGDzl8+gc9FY+r79p1bOAmJlyhQABjvq0dZi
WxRnhVKbY3QhPeg8XgEYhS26AxcIXEGjio6Nz9ipdtw0V+qxu723eW6D68pOo8KX
njIarkOydHh4DaN7wqbFkRot7EHR+d1O5R/8+taWGx4VRApdNyZ4pPA1ahzyItK1
XsQ9W/6Nsa2P6fr1VkASNAtkTG5nKqsFnC/OAVEb2S3n5G93Zj81DVnl6xgm8xlp
sBzxHnf+48Ow77V5+FT/Lv2zaFRl6nBpUWWpZCIWdvB526SFFWhoOCDtlR+e9o4n
xgXdhMYWNd0QEWvCwVnl1+RUI68RBY1eD7ab4fZCBfglDRU8i0Rml78Iy7305Huo
1R1ZoKNA/nw1p0AUwVvhsfj62MofBicaL+THoq5xXLFGQn6f7PJMY0zU2rFi/+oq
EUgQuPg5GNQGrHCUcbScZjZn+K0LL8Nd2lsz8FMPV11A1sG6NkYS3wAcQRTRCqcs
uDxZEOagnwKkLJKak3WYV3NtnXV1awWur5MHFEZHHqLaxVplqwdF0b2Ke4EmmYAr
w7DJTIdoHF7BiKxHii+UC0Je0gaxnJVkc/h/sSsaFegGugbohahiEBhSd+Zx7Ztt
pZ9c91Ppynk+RDiO7s+TMOweTWcfXclM0S69jPu6pUT6WJb9dhBaKYJYRsqzdV9t
PKIvsZkUfznp6WFpmXv/0gC/pq/EPmzy0KPydSHcBmrsaMm2sDG01i2FDu46U2y/
Npnhv7XklxeZCyS5hwqbyHZa03qAAacWyFL65Yc13tPcXIVZ6PnbmpUgd7KgeT1Q
JcyG9gfqFWgPKL21AmwUI91X0T2HSfvUrIndQIxkvXSXvy9zzBSFBL9Pt4ysa+QN
ZoRldHdKG4NTzmt6sPyYWBZ2s1s+8LD34kGzQTe0n+K9gGwLFJhAm4/CFZIi7BRs
gGzxRhkGb5T6KcVussA0b+dqk23mGCdkGboFj5GGAlb4qyf4qcn1hGY78ODPBuXP
Z0SN172eix0JmxSN9N4TZpYHXZGHreJb/iu55YpeW9LuGBxuw2LAN9DLjBiJkFDa
I9QgLP68mIf1mQxrzPkxYsQRDNgEi9q7P3hGc6X1/IPdAqV9fzVOsMHYi3PI9o+P
UOfGl7rfAMRmqmhitdNY/aGcCwVEWH32sq7bKhJNBRyk17/zKa8IbTlEXn6h1wxb
m3yZkLDBNd5fN2l+nLuzD+57yixB9AcxaOMqu0DvDjl1da3CD1t1LMqfn0uqqyTD
4958TsZMFOLEZFx98xpOG/1KfEvk2RPuybdmGyhXiTkpNbWLcBxq8CsgWt42iGEw
WFTr5umM8wTODEx7hmxwB4jiP+7zMfigAiEZkHSWluf71qKg430bgR4OQuNZbn0i
i/awvpPomFUu3CKcTzkM0IcaREfH043LDbOnemHAvh4XcgkLdZH+u3cFSJZxqtPt
gVY5q0u2HZTUB/VRkcLvIqbuvL/T6BLHNJJavPW0d0yz4EXgNH4QhmLHJR4LZyX3
ODmkes2ni2lUZbFTVk8wC7jCDmm6nwAWvPm1qhjsSDOK+FXmX/qb90/SK2OfIhlq
xat3VqRYHdz7fdOOUlrIiIg0GenvnfvQUpB6tB4ed9P/IZgPf73qu2l9mD2tYPIr
nxjc2tMgFEnr9ManCUq7XdkBrE7JKb9eSbaKI7FRKaN8Azb3P61MExYCYzf7pDQo
LMoK3ln4sbm5xI+HiZ16fUPZ6HRgGLd7zsNEOyIq6mets6LHJ/TcP6vBPDr0aFW+
3zW+38xt91mA6Qo9E7cb2HVqf8E4XWgVNkr0AuIh944M9BPkpfrPdlK/FbDES6Gn
h0yT4P3jzLxeRZ0C+6i+4T9M4AKbFs6V3QyDFqzw8+7HCisxvL9j/EuuN8NwnByn
APl5tYFdFh+ZgxpaZUg6CMzMN+GldZ18HWu3Ws41K1aOtmZKuSva45RP+Btr2bGq
gCg4wchiJjJXgW4ewO63K6T3AqWZtO1D7Vm66f9BgUBlcNqgNdUjhb9Aieth9cI5
f/fpDLzyA2w5XSSEUuSgqrbnHvWVqVBWI9EDXlEmqOLYRyfirSga6SOIieBXUZbU
DXbX5kaJ0PYp8apYjtHz3Pkf9QZonQIWe3h0QveHEXvm7jeC1Jso8fppbiAC8p1L
XRWfOWw8vkgiiYa0gJVTpVCzGBV5NeFFGOoil4Tx0daWwL03SL2HO9857q4A1ssJ
UuNPrKU83DZyg+n4M2y0eLU0qJ6iePqIFWkiqbKOPKMCprYMTv+XRA0Tlo5TejrY
zHKNGb/UjJM3whR3D1/x2H36uaGcxAYUq802Pp939nd0EKa81NRbLeOsWrM8OHbX
VbdkLgVX5CBVT/t42asiS6/UtGwcBTBnyMqDBwX0Noi9c1l6JGj3/Rzre+OqIj80
ssVVyjeoHEms5Wt4qFv4PwId9P+Xn71rIRSEkkVus0liHsoQURmhbD+Yw6Ik7GRC
MsP+meWbF8MHdZ+9C0F6Wk4Zg7/pjEONJDemj0/Kxm3GeydxyHEuNvM2FvFVMjaa
Ge6KyVFfmYXKzEn/JFfZDYWCYKzCkfMKP/hzKkkawJLHl4zwkzempnB0MyEV9upi
LjavoWDQ8A9cpoQeXfkJFGaWRNYJL6jEUfJDVLt/GPTO3mTvb4FOV+EkurhiF2jt
Bab4n2lmWCfQfQ6tmmwDOtQkXmhaErtoEPgke8YrqAn7arJ7S0N5WqJ0zN7xXy3q
LVay3Y0Y9VI0hJleTYQOXZqdHVGxr67R8a3uSq/1tqmiXGnYmPiCJZWsrUggk5vd
8FRQfXWK4kIVSsPc0kF8niW8wMPVOACFJNCraDMtutUooQpxuJo+d7H8xg+MUY9v
Udv953af0FLwj2kraggLhYG9VKCl51TFA1hss7NXsspGFHdH3rmuYaDkU0JjQMJ4
9zav7Lncgy/A2mIJz5NFZWynpu0XnSgr9tasgrK9TKyRPJEViwO6x2KkNdFpbAd5
1TgL+QnN2QWmYJVtTUcVv7BZA+G8ZuTpSTkipNQeF3371tVo3Su8sASNGxgiaSq0
UXSA0yXYBofmuaCFg1EDjwbzI0lFlGSz3QMFrp0hR+7+HkTV5Ex7S/LrjcSHq4wY
b7iYFip6Xy7qX1zM17dZFMFjaLXY9bDHub5P+Tc7TiFVRFSi0KEztrYONR9u6bo/
7nsHjNRhsKSUCZwOvlzFMrvMFqGGC7DjNLSXNmmw1IOy++sAjuSOdr024GNftevx
eRSOmmjPqWHqqz9HaWvHNz6qaYxeBSPlQJ2B58EnlTKznmMtrzU3GnyLEKLeBppr
ilsnDucqJQ2mDGBsGeeA6xGkoVygMSkVZom0xSCiBrJ35wVxA8Iq5/53ycjtGCmP
KLIKquCfPnRWaD4HiRrjGHOVI3GeD+ppcUEi74vqnvmyxFbTJRUY7aXo7QYWxaq7
xCswC7EwMP4IyVXBN3205KeKdIwrS+SloE3U2xrhdJBWU3aTHzn+jSg5UzPd4q9o
896yZ+tfTeFxx7wMKPAijFZ60ug5Agm7vLa6LIr2YR1I10fgqEaOXaX8hkCjEud0
kld3Df81euCkE0d2owLpT6skMNURpxC7QeFMqxd8hmlL0vMcErPPdiDUXBgqQIrJ
is5+RisBBLZMhNxoA6HDP7i/tueIH2PcpNPfFxthgrHEIdCpyK36MeFQxsdFevs1
RyLKAsL8hO5GRi/2FlHzmgdMAUYY4PIoeMXvQ7ZaNTX84UysHRpvrebRmjADIa1V
dYk5WJ6fn7DNle9iNFl4SYfZMB19R89SQl6ooYbMHDVSQLNLmKxYV82XK75widSF
v7td3F7TSMBSZPYyhFoWDbTSGXhW4AEBIQmvKQRxuCaYTCIjAkHlaZf+yIZy/4P9
8o9/iWjRQzIDD2zMt0j6+4Rk16x8Xs3egmLOIkMIfD6j5x5vTeb3Nvv/zjFM4+Sf
vV16ovAQfBmQ3FPASoEQ640tqGJdaniGy9COK2x4lC5YlE/FMXkaNb9RsphU3M7j
rxgutPLM3/b5MWfcKMl1jaWc0sJIlj95e7V+NMjLFSUTQt2TSQLAuZj+G4uqfyFK
/h+9H4BKR75aE9wxDpVanzZdVPqVwPG+CvGeJjYg6hyiMbnS3jFaxqzZoBr6iyBS
Unt2lhhytbwxSljRD+3jCRhgw4H9SIqv1GyGUCOkPlKGtr/aNsSRJ+Eo0aIxMEj0
1KJBfRZeuGkX2g+seMXq0DgpmaoRq21a6r8LltVSrdhl0xrI1/g10RADnxN5Y5g8
DksI/q7ubMf5ZDdQmosTO7u9zs13GM119zk4wCFfhGlWCtZujrflLl2ycFSj6GTm
MiKJ15QP4dYTFjURb/IGVUsRaKwmQ0Ha+CFprC1JjyezoCDrzTnNskzitj0Saymq
4hMynqLyFAYvjJcIy10EJyrJyNzxT4Eu4f+g7Ul8ZtZh3h4eryQAO9x2d5Q6UqOY
76VGHz/hhuiYSFe1hbC3g3+Qg4rRQ1hQyo7jj40i+DfTyLQNTkyrxRkgqtcfTOfS
sAxQ9kB7UA8ghb5uWj4FJsbcUwitrAU1ljjBT86OJG2tnteKA9GOIri4feZZAxX4
q4SlfeK6x1jozYoV7xmrGLBNN5qOOh1vkoGlbSdWpQSHdi0dcyp1AMnAD0DrKS15
VPoKyfj5cdqfcrqJq0ufjR89Ar8hCumROvr6nH0vRHPkRIlD24eMYz7MUR38PbzV
tKkrqpT7motC3zEY1kZu61T36wv4t2Q+cG0tr5rAVZD0+xsbYf3TgJzixsunnytw
vRlF4TL/RNkIFRcvc0klCRHt/hegOUxmDGj+NgdrgvUiqXT/1ZSlREzDdp2/vIJP
Q/A8mDLT9ShQbqW2/HMFZ5KjIxBADy7AB4ph+1x1yvFVGfFwPBDzREQC/QR87Wbl
s7i6Bd6mCtqszS1S02kiVQnuiH9NFvsBuGZPvBlya7nRvxeiIhNlYmcP54D8j+Cw
DXuOmkvNQhvQcuxK8DXB/Tmwhw6GWy8Iy/yBbnE7/fuPeAc9aqPpLzir30YNjgec
lG/nqyrHeXAWDZPAk/1rWZuqdcLBNqCotX472jOr5MmnKB9o62qcIoU2+5+L+btw
LiAGUlEmGCNr8coMEh+prFh51gRQ6lSnC/lq8fmy6t49MMHwNs+gH1A6cOyGeEA9
21MDNporI/KR7VeEbaTt6YAe8YmzlPYz6Ax83nBC3u7HA5+424dICkpnQWnaxoje
HkFmJch3nP9wEC/JGVUV8Eit9ADHvRy4s8LKclCm/yN7XwwO3NCzGloE0roTDl4l
m+qBVDv21MmhVH/Bvzvk64ylJoDMhtM5wWaxvmQtFvrWOYL41zeYY79nSCzYz0+q
CAmMVJxPBZUGiqsm05lkXXlzi0OS8wWfgTZGTEzjav4RSYisRf+MLhlTe96roaLL
IobAWxIMHFwlKH9BT4XXbvvsnrpAZrWvi79d+F02TKyxfwiU3sKkC3mLoTBSL0a7
trUEk73stbrH3X7QTHP4NQVwiUSogLAqd19RR8mZu94bAgZJfTBjg4LlCLb9LTDm
am9/mHFBMSTmnlpwRmf9MVzEwxZWZSwa52aSAKXn/ZYBIt8YJTLaQqShfeaXjHYV
r+uG4pUGJA4Ui/8XeD/IJSFJcpHG63Wdur6bhBbdLmwcbbb2nFc+EaLi3tTMCzJH
DyNOX7kzbzdApc766Wm6wYhiVdggYV01YapjSw10rXdsW7DoUXxoW6N58T27rU3c
DsYF2UBHjKX3CtLn1Gy83jZX7fNVNNHIq9PqtCdVU3T4qfsoZK/8gDsMB3K92iif
Lwrm5ox+i8StXhBxCIW79kzQd6MfpeugeiiF7AAu2R04LB+T7qI1xMd11W/JbWo4
zp2RoejMzUnZrjo7q6fW1nL3aFeJbI7Ij/w+ooo++Is50dk9cPaqqwXYu3GeP+pl
u9+Du6IaI7S9TOAnMrWlO+24BKeIjTdufjBrqtiKybmGbok2ZQFJpn3+69atQ76j
0VhABQuiIgvcCef42XcMKIDMX73VmxXP54uhB7gXvPRepdOGQXhyvoiXPkV+Ul/T
QrCkQS8ZPO5PsWllEP1UHtVcH5Piv2KFDSB9GN2LBI/e7D9voA/jarCFpeBFrnBG
LVYlnXBSOZOlERM64Yx63TThl+N7Np3BIH8zSncUXLSvm7AABKci0Omw6odUqlyG
vVbJOfsoRpgOZIm93DqraHR8g1O40J/AZtzWKoflZXBclWOwTdTiWwxd9aCsRRFK
WBuY4CHjfkSWMA6SWcH4Ba2PtYlxmlrzORZyuO081ImHMmwjStEA99IInt3WpV6I
XlAXfBDFUYe18a7dCwHlhIsPTojbrrUdxreAofq7QAS2BAzauQ2HMB6oGPQDYpDQ
/URSgeDrBu+wjClc4ncuYX3Vma3ldsGVImQGZ+SpHP9LQpToVI2Q01+2r8mv1yvd
RmnHkZs8AxF5HmawBHiBFHu4NLT6LHUZefQ1XOQzWgnzLZuaWaAaNNYL6J/Y485t
Z/QZHv/gvivu3d8ry9sPHm4VRUmqS1N/TFGSnc1WZsdRMlVRjFVhXAt3lH6o7HtY
gOUiDIakTGKLKVmhiL/6EHJT6DYixrBow4uvI5YG3y9wMtWm0ys1RwgdqnhNrkaU
tZhJ+ylrXX8dbuCPghSo6OOYVIgj8397Hg0S5LR3+lBejxe6TwykhrkdiwYA+f+r
AzNvXwTzCMd+B7y4L0HSkrnNLEkswZaR9GJA2ayQyPvVd3SOSho5fhScCpBUzwIV
9v/e2nM1Ipoo25EY4Se5bKAxMcBy3sD/BZzBmG81DAF2hWr1tBYA5/MR4zOQD3j9
XLNE0Qdu2r4qCImM21+3E27Wnf3n7zgeLnkXDhmk1xiqIyP4bH7J0HlehIBfSJB2
x5mDf+U0THXhThFZRRo1Cz1dC8wWoeNzGCSQX8WQs8AlY2pimz6lw4x7AUU5jpXq
v9ouX2BOBKmhBqIy8OdrxAaL0yovRnr8t7UbpflZpAvTGhZkbIGrJDg54N4v3AhX
cumxboYwRUwPVCv4Q+TMr4+Fw5hBD3BEHvI8+xZrO0dp50XR0R3cD3+gbkB65K0Y
MP8o1U2btYuV7xU3C9Zirij55WqBaZ3JJ0W5eJKc7KaOKB64vWN4AIAROrQGcjYo
lMIKkaFv7VIgh0tKHOz2IADMRdfd+hkwT/HlIAo2/d7CP4IJjM+P47DZbzZ9WZHN
Dafp42eW/nPmQPvYtgAEevDfaERF9LVP5XcWBJtV+S+/Gfjv5hMk0blHz7NwCp83
odbSbd8loEKRk34cc+FWuzeehuj1dSKxTOjpRhUqOL8Uffdh/O66hfYbf2i6Yvj3
Z1yDmsaNljlUHpbjj45ifheRUIoAyKEMQfchoB7rEUk5YnxMsI7eMIIGlUsyJ/lN
/0/siKn1Gk+QsKuDExQsNWUYAviU0v2iss/In3MfP9xsV2U7QJoP/rJa85jDwzx6
kxS6fFBQzpEFH3N9kCfw4fbhzXx/z8q3h1zrWtoGQGsyVTKgKlMLGm4yrl9vziFq
XW08NEHWOq1caSkeMFwGu11FrN3QUGdR0rfpkIi+PPhWWmsX8ZHv/7MWpB0rk7I0
EBtN8wWlVaxcDVcwzwM8WzREOEh56Yz7wuVypF75AWQHVovm9Q0T2h/wuaMnF7uu
bL/pDvKWd9FUM3h+zGefO1ZRvuaOjFDM8OMRtZLKJiSLjzqkNKawMqwPOZWBbFlk
Igs2+pYmSiyjhSve2Lhb2cWS7kk9i4iolwTHEODFWcCpzjAOhFNfPuGUpCqM8cEF
XkMJ3PT9vqgrnSgdkFwt8Tas6b7qF62eWkPPu4WZTEj7a+GkcOVcwn+SaCx9QdKK
OhrkRrtknbSjqk+v7tfXG3aZYSBd/G6gOVEY+S+9UJly0PK0F/l3F5KLN/yWP0bz
jGN6vTfSG1RoiiV3snw9SR3o/DAFRwg79UrI9q45zeUASJxCcUVuMBQXE69mD3Cl
SJtc1InGlGRIBllUUEdu/RnK9BbTWs9SWV9/Yd6FJJLxDQVdhsCyby3clht/sUFt
+Wfb0CegAc1P0p9JwPT0paQL3/f+H60W1jnKGYDe9vWRZ3sKYDHUQVfRPWnNNrrd
C/9/rTcf3bqiJddfyCCePIWmRo2CTtjyS9zZagt1rGfPzOLxiC4Mg/uc0UTYTLpP
QNo6lm+LOl6EVneILah+a3Lze8u4tSWQwcty+h0sobsEiTXVzmeoZi8vTMR4VHLh
vLqMJhFAzysF+hYWS/tyJFEGEyYw855fLObjYULH5csZf9jZgygjvl36WBv18OsL
sN+SUfHXlZglLLPfFHXusRti89KT1AoJ723dU7VU3OAcgSfxFzqeQu5mUS66Vl0k
yIk30SbMnvUxijw++fsEy++rtj/KLUTo3F+REXIGueFMhgCvfiJWOPMmtzji/4DN
pcZ79CJKLFBf57MysQY91cF06n1si8s4AtuntZAuyFC50+iZcmMaGrkxMIRy05uT
Aw1mSCsQBDTnc5VpnIQ1ozEMH4ysWMP7MZq8HgaLNRops3Z16+tmWQrF/rnSIDT0
kXCzAWuL1NLk7xEQBfJj9sog6NohM7E62TWR5i0D9lZwVVR9lQl4Q41mOR8vOlJS
QVPEIzNKr72QGPWOLpmqtiHm/xo37fymtF+ITu/tW43AKL/abnL+nbueR5rDBgVY
WmhU0PS6o0IH+CETcMdvt9yWWhkLij3b9ZHBhus4rv908WxpavOwHKVNfcreo28I
1LWMvWNWpiiFo6xEaGj6CA6duQCvsjkzb4rczH74lfj0Hgzt1mByiGIJzjyJLpu4
U3ubl3tZAwZPLDhiprO5Eb7fFuzl9XiPwlvH1tVWh5ylRgN0GQQxYpYFuQ/lt2Bn
w9hHvfpbfl61GxoOnKiDjb50g9r6R/UOeMggwVMvOCaQCOqA6gJOxRLFj2UYSh+G
6jxEne4fa+s8n8d1GfGTnd0rn+62MDuikG/PIWZBWji/9s0rwrSS8DiGCgZC7M7v
WcACufWabPlzrqDyIrbANqjSa24HwXQaK9iGQD4oz2wDSxk/8JnpwPjKgKKQRNUu
dLUFBaZnnmzg7vrBnsa4sWav37IWaDLu0upDaPk0ShuGGb+/5Ns0lmWaY13Y6f99
nv/rvsQ67hQ4Lc2ULa495tNx8ADCRNXvUZ/OZnzBH4ED9BA2rB65ifBhGLXAIowo
haJg29MNC6iTMfU6XphFsde/poW0WdMmnWojmo/dz6nz1B9fSaR8M2H5liDOEoIo
4rzwByQk5NTdVdQd8Xzm76rj2peB5OGj+LHTFn4yUZPe8/iOw7StkJ5TZdc6MdsL
QoJIIhkSuwHxptk+6dASkYq2/sD50wr1hFQrHVkrfNPA0U6i5zSOXZ8+N9h+Dbbg
o9zcPsj72oudPWtEiytm7E3m/dSSAojvhQkqMgPKPYuQ2jYJqZFfY1gTAmKJT807
NsVuLc8I50yYAd2KzLz+ZWC2gBXyC8PlOnhvW8RExwsPq/ztFKKpAN3VbqUjse7D
wOnBKgnGbXvuzxKVaQJhBrFKM8muPJ36PDiiGUtZW6N/noUe1kd0h8jFX/PcY9dP
22wj3xKzOtOYg4i3u9Y5Eg7bSFcGB64Yq5maFGsPjQJ1HQCWcEfCysDHUODPUw7Y
oI3/bdRGDsjgufS3x8ToMusfxkMFEKw7eqvf8UsAY0jHh/yn8t2IFZZ+2sZIh93V
T7h4aUrkONCx9Ct3Gsofu+Zd2mOHEWmzWhMh9jBBSDhkqut54wBEkGt3zhrQlNi/
imQsS0EKp4ytai8ljVxwdNnecSO5NkR1Tfv7NZECLReN2NxbWmdOnQzgVHkJF35c
blfM8mmNMy1kKqCvOp7oiv0y5ENC2Qkoo7TVgfSvQ8efuYqGW/CZ8vIeCtmGzIsm
bRF8sQUo0peOVnLuni7I/jtdvSwWNhA4V+AcR3mO0Xja9/LutjqcWvdNf+l/O7hz
c7VauiZfzfkZ0CvsLjX9oda3KjJLdzEWn25af48PXj2TR0famhmt9n2yDC91ClRA
a5nDKeL94B/6QeWQG5gZtCWCguAqGgLrugnLCHNBkDlr+s4KglUUEbPJQANgFCIC
aXy8IMw3yjRcttf0sdjzV9/aY+xhwmn5KmpqyDY6zvgVCfs3pltvDKaeDqn1HlHM
2G6sKkNdQkomcFlE2E8DtlutQy2FJGor0xezNx+hp+7IZcNpHYPdZYvUELUMBdOL
h82qPZamhFkTtqEBKb0UF9Sif97Yy1pFGhKO3UJqeIh8sVQoVWTYVskSPBWDddOs
SJPernTn359ETlVCrFGWOl9j2zKI/SDr2OeV+ZeKWTsG9xuEmYhsHfb4ZU4uZl8Y
ieBV/oa8zfbxWEfGvxuPiD+sfXbzumsQMEn53wnQ585jQBLGP0AtEvCuOU8LLqA5
RF2L7bR8yN4NTpiVowjD2V8xF91Xw5JwNyS0XnXDRMrhMVyknlbNvTxq1X705OvM
nFiEyMhfjdAg/BphaTJXLPxZ+qJGrM5ifrmt4BGrnYu+koUcZ4NoGhYqQYC8zk5k
M82s0aXaEhusNjyDE3CPgr1r/pKS6ZPXnK5wv3RhVTrYRowFOy9hiRwyZF+Iif0q
Cg0vdyrA2LSeCQ9hOWT9FU/uj/gSzgOzHk+WKOfxHJAvSl84PA8Fw85MEsLgX4mu
QYgOgbnEQATbj37qadeAZ6OIRCG8gGynhwI5rwCwwps4ln13ulA85wnoaJe6dHKr
qE2Be7mvZSboX/1dYshgKHkRH/1zQMhtwuqzbXtef3IV7/3yDjJUzGWm3BoJDLYH
HikS1VZYqloEyXfMwyKtoUOCWRTgN+XPJfRc6h6sM4vUR36iOeQYX6zm4xuwJWpb
JjtvQc5GLE6gfRvih0IOHlpg9R3JkC76ApnmTineb/Clt3MivIcz0MDlQk+DPvOj
oYwc6e69ZM9l4lUE/Iur9KzIn5l1WLXVM8galDS1odPgOU3agC1hNo9Ed/OK2up8
llNkbPdnjygGzzENloOtev4yLXy7/VfbKDjzxwDixFhQoMyMeFBFuA+ufxl+sM7P
7j2u2CqMA3O21bYNAX0qb5M8p8Fng+ENdrsvlxcoO69AKT3EXv5MSAtvdd2q1d92
aVdRVPClWlvGi0C/Li4s0B0DgLgUeZjL9vxL5FTZgzpem2wOM2/WK2bCbjHs9mLy
YZzJnsBSIdlwqw+aMooYabOKHHU98cSjbY8p1sE4lyUe4LlgzL24kvgXTAq984gX
t9Bld54X5/t824FMfAZRtYvwJP8jGFz0Dp75Ve83kX0W6Y+/gm20rVYjqhB50dYl
7/flLS70J3/4EiYrIq/6eePBZTqCAa+CWIk0HjxA41l3u7rKu8EIx/S//eFOddzU
B4cRRX7FccF69C8z9F0I1NUrgWlUcS9LuAzEvuYcBjO8FWGIZLMYe4BzC/EnsTMD
mM6mO7r92xyJKpzb5CNNLUOaN7mgXybr7ZpN8rt6dDY8SmJCj/SA2tgrEAEF7ADf
4XBHsxGGp7qN3UJ666mY95ixsh9afwNOFTJROO8GRh2u41p7MiyprGD4F2X4VvDY
Z7xj9adIQ3agnxuS9rCWqo9IEbPx1/aTCu+eZTUWTSain5VkXBAA7UgHLpCVx8Pn
EJ0SQx6ZtwXCtUY2tV6MLgRmFcO3uhcthAR+UGbpjmrLFckoBbT1SMQMiqH8oSqG
J7yAqXrP9Ufbs1VYp6RltFl5VeccajrXBp8LOKJxkZ3PE/re65ZCPM0lKvkCz5eK
4Xb1XzPk8azuchic6ni9MmYWwN4f+pSOf+GPCJ8lNR5zTGAfkkGoEo/6an9cq9sD
a++ZEIyMJ0+XFS5o9QXq/nozX2rQ5MHx1YRUd0JDvfVsUmRbjz3eu4TuifZDCfRz
2mBPcPk4Qg4fdnToBqfKzXd5Z+UBUJYXuXAKYLYt/5Z0xMGbSfBwZ+Rbxm4x1Quc
WHD7dTwtee7kZSUNT6byhm0N5yOMDAU9ZrXkW02DQd0cErD8q2gDFDGypdqsqMJG
xAOZwCEKxQqWMrVpRackE0WgwjSdrT4EjQ6hxoLmvEf3Am2O/1i+b3XTLU2BCCer
Tb0X52lLUW8oSoHOnaSVawxci+s0Hlh+OXZyvugCVgjwygeckNvxXSZ7qV0RsINM
dHGhwJ4ckuig3j6XCZ9VxhbVjZ/SgJ+tFEvyGPnBDzPjoywb9bLWT/2GzpNLoaFH
lyC0p5NO1uTQs64v5L0rSvvQ9diYFNVQctzEaaBONGJWFUlkFSsJpFe1iV1O6ycp
RB+NDShL2U5dJ9zveT8Q5cwjQaxlGwyQ6aKwHFSyakIkA10VSnpfgfQtGdkmEqMj
n1yZ1+ifjwZZ6CaIpec4hRHSq9ViC8lPnx63tJXqkfXxgQOEerwnFYuQbINLRMiF
+SqphqUxwfl5W5wOuvACCvTmX7WUVRcQP3xTe2wQOprsDeuQH8KUzfhE5dj885zz
3dHlFc3H2+XT80oVFtqctol3Q0DsDUSUz5oHTFvUPHeSEefLx5LMWqMsqjRgC+n7
netEwk4CHE6zlPtFp2UkIAD4jGn/ONlbZn4RH5Eq71WOK1NSLAzfywPVhlsbr+I1
tOCMDBADWHrUgsXtVkKIxY+uq0jZMwX6JZuF4YnNiFlX9j48XTS6YApBT9jedbkp
s/Nn9DC/OsLiGIPev0VfQpuFw/gEcD5UKzBkdQsDozNSZ3N/u2KpTgYkTD9yYoUG
ByxVrqppQeVvBsT797oCN+2i9fUdkBoNK2JasEkrIVpnd/XtgcqWEo+JcU6Ycg1C
wYoA6GmP9cUTRDrBuNtNnUF5yuxV4EJG13Izx+cQsIHY0g2r7jVzjZqU/xm+xhcu
hPVYq7cjuZglKX/1Nz1Apaowg2Nlm4WfSb8GMzqfzMwl3IL+2IKQ3v860nFDhXZs
Jb3epvoH0g+hO3+Qs+OTtkEBayK3bfYPNedfQCVr+9VGVbLn4F1QeceJ1fM5gtkY
M+FUiIgGd1gyQ5AUmmy8QN3bbrZtML6yxBN92VFH8B3kWgFZuFdpeq1RIgVkEhQt
j8+5Yfgq1QY+Aq4BCScm/WS3a79fldv3xR1rkC8LVnVpfCcILiZJZ0rred+uuf5Y
UaO+aRk0d35eMhFJQ/WhsoW8zF2KuhtOhuHaottfUU/I7Ew7esLGILZZflQFnlwx
81T9uqtXCna8AvCcw0o1nZ+9XClYa8L0x2e22mlkyXa7CQPrOhaajYFCpgGrNxtB
5dD8Z6VX8UBcoDyijUXEdl/7k9M8UJTg5lwPxFEp70ueN4wrLs2lPYEi/7JSaLmB
PPiVJ6K1KuncdZeF7adXkg3hoakvFdi8YVBd5QuxMtiHO0jxOQCyQlsgZlNrno1g
45mI+dCDVc1PQ5dc+P5M2hsOJ55jDDhkWDvSWBJzFjKR1VDhGJzO9Paulp/mGoo8
jtThkHgvAqtzdAE8slf3d+5WCamIfNNxcxbTL4pXEHImwUcwyqZqguwOg+Jb8N/O
45TOVnicc8CIhQ2QPTFauDyXpuJrbHHIl2+7dKgqmWyY/HfvIy26C3owrGB1ZpQb
TAxnjEmladZG60vqeLSh47oh1RgP8vTSuOuxJmowDRvS0sF+/8x7ujODEMKOYRr4
Eh8JZtZrNQ2rJ5IvgQMoFuE/UESjXcckHu0ykerVS0be5n2uK+THAX97RAL0wZ47
hOi1svcifYTMR5sczEu1b1V759HiQ/QTpRMzGx28XNLVVjuIyFnx/Eq2XuchnhLn
5phTFIm5rldeIxiQfbzsI7x2SHXulqBeth3ODtp+18++b4RRHvj8DFbgQmkPpcWq
4Wwnn82YLN66kX5TC0pXVjmzfeaHaoUob6lpoU8RYhs0A7SBnRoXONwKEGS6Dn/S
grXqCwm3k9yw92ecvEwBDvID8BY7ZkS4dVR+MwQ6Z2Ev0ih8cDlVyAUkN+77uRpF
Q1z0vXY4favxeA/an/ccG2aBTCGMqWa2d8EMJLLTXLoOFR0oKPSv5OlfpqIGjp5W
Fkbvv1VTJJ3d7iPD+eZikmvg6apKbKPg1zJWQk8i2EvZ192e/wSjeEJcHkPyNM0/
L0VRemp977BvqGXcXgk0ayqf2v9ofzmVMepVi4iJLTK1SW3nnanhgGIStm0UUm9+
Kl6pFKXQcWNR8v3Vdg+kancYyn3DJeGEEOKqsco1MiK7KWqBhLBwQUFDtN3LptvD
ehYSqWTIT5t1u6rm9vrm8R4pjdx/wBgnSnqb+n6n3VjuQX+lhxcjT5a4PtwurQIY
euzEa1IGNpMOM9fjydwwhBceoM0VvoMq0TXqJvX4kT1s8w3hY4SHSxSpAVWm+ImW
9IwfPGfLsE7rn5NGaBkBz8yEXCkXVAH4NPQZ2xVd2THXrA/FxAKTuNW4Jdo/Gd7x
BUu/Ti5kNmzWGEo3lT6nS+q1TV2LxMWAjgCMudzeehiRqIMT2B5AOY8mXXDfZ2th
rqIXNDCxIZnstcNLldG/gXB1Ql/N+cKNtCs/1n6iaXZI0GymZTmxGYLVPQxJ9FQa
srkp4lR6T1H4fOPPFcUbu7tj7lEuKig3OfwjXvRv1PIHzOeMH79cMrH7fgcFFHxb
zFZj3vAG9MHgM6CfLBDou8rR00HRMvkqErWD6nRg7ZRSxm6B57oWZg0mahJYoXT0
ftco0+enUc4PKcXYpAPoGARVq46petm0+OzwU4bDzHH/qjXPYVBuR7C89395SvxZ
vxMMWM7leYmCm95yG3NVAA5reGPeihqab8WicxsrEmLqmSrp6PpKEIDxxuHBL8C/
6vu5GcbKKn93YIEPrwCun6VYPk34jBetghWzKOJC0yWSAo52TJE04LefEs9eAgnF
bTDgUlclVnLbmcRGkWEm5EwJOqqPMIE+db0kno5O2nco8kEqa2UFeFVHCD9CQd4a
JCjDNiTlThbE6yIW4ZZ/QyvXW35CKKq/L3k19qHijfAi6zy8PBL/GqMZCC0u05FD
5b57ceW7/ovrYTXf28eZ5kehwACx8CGSwNBIvxywEWJ4p4b81JVXoRhRjfjtVCJ9
qkQubCLwdSn/iSuaDWsqqkn+oAdFcgutLlYIU4m4o8xO3SYVH8fCBlEP60EkXzX1
bd8he+dA7syqE+vMMsaxf+fVz0mtX/KArYquGTR/lJlF+ZfElPgB1B9ns9GK4gK9
E2VWqvrs8O2pksuys7ntuSq8zBHPIDFLhg3/+byjlOG3Nt4fAfVwPjvw793vvmvR
6gSPvSHk/KIivKa5kF5sOoingAOO68Mk4++ZyeZJtSrJacyJ+BkZthO5n4iccmqa
N6LZuMU1Z9uMrw25rPTbcNGy5W+a7pGI+rJyPVmy/U3NVoWlvGpqi62ABZAnLgH/
ppVpdTQcG5hjJOo+0ZYeu648OdScuhQjIONyq+A5ALbi5mpW76RSFCoLqYbQgifc
un4mi1h+Plu7vDEfDN0WtdzpvMc9f5yuiD2S+lVzXRz0OwSJ1Py34IZB1x0M3GR+
HyTHg2yn3oCeViSJ3g+ndPHHAYmHYAWBSSXnYqHsExXh0OReVvDZ853w5mnz2RVD
w/3a37zNQuGnmKmj2xlfI++CWh3PC+SOo32O2Ej2C+yog8QXNdlylYJgUw0kmoVu
Htcx+FpvgSfy+f7n42QRw5owPoqGmmgdXLIPbZUSDEpzFfQA/XDk/l5hQ2O+jQpS
tbJxkTxTaBlkuDoStWW5BDsH1WZGu7BNQ57p9WxURTTtBRfdEV1h/EfVGgLMtoiV
5rz/AGWvZtbTr+cVFVG2h9SVWDyiiJEbeRjkDHmvpx+s3UNR1hM70bWGJgEOAjDq
el5GR7SyYHLqs8cdJuXpiGCys10RAgXqRfi92H+QPEae+4dUiAVYrU0NHSFttaRU
zB/EMC9jhiFAQxKGHLgAX3W5Xie9dvUeXQcVPChAkBGvb7ek7onDr5CEIoUAbNCN
QIgDqxqygNBtH/CaOR5fjTpwOz5P/EIN0QNue5STnSH21cUiRf4sgflV1fqsEoEA
vMPmx+fEvT+X9kFv8kwdX06QIpOtgEF9B3pbgYv6Bplyods7YGezmyxAIekVTRdx
o9XUz/TGK/5wyaRZkk3MFX54WJ/+Gk1v/JAHr01FQ116xZq8nqgPF/RTb9bJ260u
JIyvgMd+KA6pQ+oTWrcrS/CQ5koeQ/hBeVAyUX19U+rpk4KIRFXd++i+q89lhZPd
bK1C9MhkKbv9rcX4Kc56iXCu+ze7Mae6ktRlDwpg60vFBLjiyh9pwtUnaHVCwQDO
SCMH4cWmx9R6a3Rnn7gSjdLbRQZpr8XhQWPZPwH9BmTvJsiMnqaDBP75iXILutG5
CWNkknH0DhR/JqwBnygqPhxJcdm9tEPZyJoTrhNQksKKRPjIlI8jtL3SIXjHucXm
BZzuIfyUx93jy+F+IFRffLjyqnavmAgWsL461ak8snXPQtxY/1v33mtYdG6GwjFf
fgruElVbWHgoed8V8SaQibQvIXxj9N9u3rIMtIKCYF77TRAdwHYL5LjGPgC7m9bb
wdwOLHNbDDqdXykt9sIhk/qv8BacCHR/jQ0us4I8ora6b5sGQon/41+nTAfaMikq
ymyBS10+rIfkqQ4ZrZe6ZRtFcYzb5Kk21cRIo+m+kCBS0j5ssPrv5UHtyngEO/Uj
AfrvkmPujXXkKAtI8CSenbA6fzNAbSHwK6siPMLCgn0TO0gV4LKssNkmniI47Qv0
m/ZxYQCGInCrss33Ki7f2Idzn2xZySuwG5w/9CQqX3dIIvLEbXFHB1bnmqkqjmlr
wrW8tH5p041pfja7+KZ/8P83ytt5UOoYuzAjwfPlGpneSDEwM4i6j5NihrsJFRRM
3aQgeHFLAqtVfPssNGZQLiqKKwpWleD8OH2zUDFlrf+puw5X/jiagA/zhJeU/zjv
wzJzoK6UsEF+wbi3Omqu1B0bql40Lr3nphWGLQsMCuJkJgP+L4PZZUayCfPW+Hpy
P/hmZAiZEk8mVdiPaDd3tl6foRMCcw7se4v1nmR9wF9NMsmdwZYMOq6q0FP8x2T9
IEatcZLqR8kaCeFbv2X33MNEmIWZ/IXwwvF8mvrzEFACXFo3U15Bpce9twPhzjVb
Vv3PVgTgEI/vDYJfcCOIgwX+YYDadYfp2IKdyHcUF3stfPR05y4Z9Ps/MlB1d+ae
SZhITTyNDQcKuixKQAMu4FizDl0PHiw0cZ9ee5UCxTvb/D0ihrWiOabGrQsWtQT3
A1FTAnLdNrUrXcAMpt8oLd8mpshKr952os3u21b7dMyZPjnVqtHjv+GXyqZ2wTkx
8TN1fOZS1Pe+HIR8s1kigu5GFvaKj3mmNLYjC5FHMPDvuCc0D2CYQzjjjENQ5kMS
ksx3b2qD7nXTpnqtLfBhvnrj8cmDiRfCUG9mMxQnJKR1uH8tGXwcjtqoNbl7j3h1
Vp99R3Sl2vxvimUuEeSBXO8FnhSnXSUtMHqGPfXWo2RaRTk8hMYmm4GGQAIQLArg
O8ED89cAuQkL82H8ABJ/yh0EH7XLExELww8harJxx9+jhB49oM9ebyFZzBwB96Tn
aOlrklRxBChx7bq0HPpQSzT3wUZWFk46AxEtpwlgAVR/9JkyYAjEagYZdYkfgeOL
yLf55gqd2+/hmTN/od+SC9My4RU0/Kei1CAkKcgH3P8bPkI/t17OpFIAZcmexOru
/pYATUJamujQYk1GgUbcQJMhUAL5gpRmOLtFh7YF+LDrzV1tkDPcpK38NIa3E/Kg
/eGwmKSBGwmeCq9SqUBcAdYFy0c9KVubyps2PfaENQfYNrM0PEh90WdoN9skmodw
yAEitgWZmzjo7uQeO4QD0LSPd3jOWq4Ipy12uB9i6UIgTwule9iC0iXJSH1zwhR8
OUjLTE4Jw7vADl9FSScacyrbR8vexx/1zvh5aa6zZt+EJowiKMioNRrdmmA9hoKx
E+yaIolFdGL2e+hpl73FtyM9j14H3u1g8fL81oAy9FA+5nxYCAFg+w1D3JZLG3B8
Rovb+0r/J3CA668ANL8sAAxPtI1EVrIRIijuCONCKBuQzbsKGdzj2+Eg6r2rWWfl
W4azViEtkVem4xUqpmghjfy8XUN7mRAnfht1Iq8YBRkUZN0QJFWmuJH522Yh5ehz
hLWG3AhAknq+ZepKlgc5GUZ95zXWjJ8YoazEefUZCqFLfK+4BiDOYIKreQ2Rzmzo
nUs2XgSwvmEKLqfk58o6RRLwnKuutIu2E4yNyXuoJ8LSpIpff+EwoIYDoHt95n6x
p3Qr2xol2aVvDGvne9sNJCuS3O4TKA7wp7frqKmql+5wEeHYu6aD1sP9mU8TPgtC
qYM42GsMLCjQjewuorfKvXB2sO67xP/jNo4of3k4U/JQ1oxBeOmW67d9SM3ruIxF
GlhObVBV9fF2/FAXoRBoSyY8yZSv2NIdaq11FLagmXrFHzgjLxJkNQmXJhyRGeSj
XbUimoQ2lhnUWSE4HMi/yZ0VQYWpu6Yd0pbuRuwSsDf3h/ps7hh7KesmfbGca9fW
ngKotDeTFEy7JDIyYtbf3tF1ER8r0ROL1PxBUbM7OUdVcG4Wk+Xzb+6zlcpBHFB9
FzMQV0lE7en77m+agTCMnOElYMY0gbz8bFdjwZBMHpBkYkmfpW8/diWEgF9ebZzG
YptSGHbY8kV6aYTYu4+u35yadMK3HF434VYUAGpRqMwvFdDBJgWsRcNpUWPHbAP1
UOEu8bbZXhGEY2zc/nxQvT/6SKs2gGpBml3rxWgL/6k59+zpUUSzvCQsc1fRFwrk
FD7mn8bU9DgiyiDSE+MwVzYP340IaaiXQWKeU34h92+RxXbSM8KkI4eoa6q4+jlE
JCf00yr7UqGOrOH4i+k66wm59mADe+zggh7RUFVeQ4RqjLNieR1yhWyMgU8ZS1yr
/j9UTz1+/Ox6C4XCSaDBPH2yUhbrjnp9EGAlM8Q8Vem1hhcYGQQCiQA7gfIo787Z
kjeQR3zrCE5PKL8ac6GU6iL1wz69ASy5NajsdCm8l06IAJABHMaLVLOY/FgLZnhF
te9HZudqsQoSP6exhsJ7KDpmM0hh7WYILI/lJbQ9yrMuhUebEnSjyXgImXzCFYzd
Tn3w9+Kl0nSdHCJCfC3QKzktzq8kys+M3ucSBWaqCq6IV5FLakabwCkVJYqiEowM
tX8mChEbVOIxJKUGPD1lKVWaa2It5mNr0gkGUWFeTk30tt8Nn/U/k2KcXmpUb/zm
bmRl/O4vuG5JgPcl9vcGUGGE6z4XeyGswUcsucMfzUMJlxdupD2oxk5MzyMJS89a
x7k+tJY+6VycQ5DFSJjPu69af2Jbn/Nf0xSUeD4ieeS8ekjcjmytncbaFTgGCcI0
E0cwe5+lQLLcYAsbA1f+IuCtNHB7rliMt6Kj33eySmiof9vcligxP8mNDLq0lssy
NR1ZL5Rqk1J+LqTQhuKZn7YxJWG4sSE3OtU3tCG0Ts6npaQVMPv+cMgB9tkY5QBp
4YsdSwtgdAZ9xxXTlzAv8UFRASLUUJeueXzllZDiKt6rea7rkafUmN9q4885JAja
zyiUAmXSf5inh/oCcJEp3v/jVC/q1AItk9HscOglNRyDefdWA7JXW7Iihp2KrB7b
+8+hZ5GGmpLxwsCRxc3ZhlYGCdJWKZRUqSBTeMnsWZJeZnvFmnGbtuZ+R6b5hjgG
evvxtB5xSkqa/5A+8oD0Ee5kCSBCjiJx8E7IqcF0wNAsAdwBYT0BiQWeoUnaDEUc
maUHTS7kGTFpEvPDAPAS7OV8NTpKAr4h+rRymUUPb09UmOVNmqTuXXpD9VQEkGF1
6FQuHE14URYB9Gxd0FpT6isvxfd1c0LTdR6sKHuNlXUXHQvdSbHMw/B1EtGIplwb
HB4/VQfpM+S0NETTPzTyEWnHSl6FdSXN9gdwYcPo3OYsg3ITdUhHmW8bsgVhEqUq
Ed6qwIDQeyuzRVj4JsrbTFg/3a2h7d0ZskcXhq8icSdlmimyShvJnadgMq21tDkH
TTQPWda5CCBjA4H+CDiAg1grxM4QiVkdhzb70mgtsFGyaUjUNNsGTNDV5OchORUo
otQVGyvk8T3AcRFwCaDbIRDYPX55nTWuq1ugfpMH7bWXqbKe56v0rRx52idvBJvI
DCQQR1sFi6hLkTJ4P4p29eV0MkUU+R7ae9owJ4IDePBAusPejwhOX8zUPFG5cD0p
6sU18e52t7669snLbdtwZFlDWMkm23+xK9JIia/PJpy6qIAI1xZnC0B41M9PpG8c
9ZD8nNpFPKn0KQLKNHFhLCgeoEqxZHQOUxfhXADNGB5H2gbIPjNiSwfeVhbnt8ZU
C111sUvLr6eOGCFlcsmYQbz/QA+Q+xrOFPLmpQBryurHJANZmCbyOB/XoV+Zaqav
9G/CDHugSsN4dqKK/aUjvF9UbClDzDbCZrvh1lxoO9iQTb8kypTSLRyeC+lsoY36
zASOHWpTR+VYBZ+dck+t6qrnnEF/F/5Bw4qWxKLEkRXytvvt6gZUBhYGrc9hToxH
GWlLJEFUVnpcgW4TzmHWFjg7usUcYP7n8IM1PX3RjqS3K/bA6VfXWb1mPbPLUh5s
pKqKw43NwUp9v/b8PCqMO3kKQPr/0d2yBnPo5zaDSn2Vuqh1qJZQshr5halUk3Bs
nRlvjhHRiEOmUfvNbzVcmrrFczgWJVjreg6f6KcbV9XbNdq8qEJOnCpSLn2FBgmJ
h+xIksbW3l8vp5NKa4mP44jjvHjcvEg/CSQ9VcQQ+/fDwAT4Px15LFOGJTNfJ11O
MECIJTubSibLgwPTg3Mp0C9pso1TifI46bjuOGeoSR5JEamhJyQrapdGl3ZOqJmG
YAbHkf65Klv+OqDlFYMlIdFE5xnmu2YBXNjN0NsH4rCpGB7YxmVsKt4TorfH+5vC
JWz9mKz6zcaQmJjN7EJ48XhZCRKGiR/6Vpahg6YNbZF4zE2YZOy5OyO1yGSjqbJz
ZmXlMyOKQqo+dsRsyFTeJC7MsaRvArBSpGUbRRhTVGiiW8V+kdibv04eWNSARANb
WIJVW713T98bjkNBrKpY3VdZo5fQ+VuX+VfHheOBZbxabwO/OpaO7ylwdyLaQw9w
aYmgNB/Z2QAfyAOOLAxVBGlzdqUw0SWHGUGTig+FEcNy4TJCugl9gNJxloYxT6yR
+tKdC5y1R0RSLWhZYkMd50JoqskXjBPRPsl8wVLWgDfuHtrwYQUGqANAaLy9ILSK
yXmjN7Wx5NhiaoUuY6M1Uur6sXRExn+so7AbRreSNfkyDuhpyMLeuoC1p5HMwCLv
usQGDxwKshJcsPHSWMQQeOuRtbw3xlvuS47nyqQqSO4qbnvT+iIKQsBsmBTPElMs
ISUdYjW8uDyXEMVL1n/rGOwOEG85aqi/pZYgnc/qQE3P1nLYvPbzczL5Cn41OgMt
b+jsIAqEZocK9bn0tD1S9Z0opAjc6Jcl1pOcCFWfEQZ5D24+GM+d5bbqNhrwu9CA
8oZjF3hc2uSHNjL3GYVpJAYXGH6pxKPYLQer0PNDNrwU/ld8XqkexeXp2k4hfYvc
KyVqIZxxElloB4xCIQZpRxGgaSYft2u3QCqUVFoIVkkmEV2gUi1C6b4sLl/y9oYh
e+utoueEsIeoqvxMA2H2WCoogr1xcf+OOxKpkRvSydABWwlp9+dubEm70N3PYnpG
ZsfPxKH4+0hMShwsIVsLhH7S0poczuOIxAMebKKMdNXSMulUhw/XCRj+gwTsZrLv
tVcYEs0kri9aPeFXgtJQLFSPAUm0m6ha9qHnlvX1NkJlcW2fByDsqB4MKKegVHWa
jRbrzMfaYgEX3HEwCloYFBDaj4sjKFgN/ESRsDx/acfssbDxYuNBIDDjAsMhwhXa
MxG2YMsRFEaitrgbxmOQzB0lKDg9jZnzWmQlu+sQ8xkHFSvL1+NcPZGG4vtpkcBQ
j8DN9Xyaim9YLxVupJihmQf4vUiOKBRQLUTvw4VRgGRy7OwbQ2AfVzbCdn8BcaKX
F49UYoWyf66neX90omQfOfRlTCr0gifBa5TbjCRYEhHY3hUI8ieBLcdiVpNxhACA
0f9emng2C36N7769JUKRCjzCjB9ZynbtJsWd+qkWjsRf8hjQd26te87Re+Ol+wX3
VX9JN56v5dKoHQV/q+s2j9N2Eq054NAi/1uHMU1x1YNxtMyjJCJhjid0CwBOPF4w
dmclPvNJElneRaLtV5CY5filfBtFhAOHYMzn5QT1ybA/OHBw/Kz4FkC3fRo5ByKG
copMsm7rIsNLB6YJQ+HrOvbWolWgtayX5LWucWyxiLaCHa5gnQHaIqpNpGKhp3Hd
AWwafP4dBjvqaMvbnm89WPyITPfkVbGnowpIKwveODxT3oj1vau2o2KCqq9cNuqG
DFpKq26PF23QX1uBm+PCYMa/FQhmOGycjfSP1Y+DEo9E9DxInNNMtqtC5Amha2Zl
7ZHHX+FcxJQ1KNxcNhk7j84eMoemFB8WHKt9OXBNR6tPAPR+zUkjOU5t7FLR64Ja
x+4tAMdgaOkjwIQTnGdKeKhFr/lcfkOfwyUEBjEv8i5BQ8zjMAzSX+K6YpustLQ2
EP1dacukqNSRXQyRF976xWqON9Yq4CyGSGYeo3TaFyoS8j4SqoA5DKniKZ+K9Tku
9iFaOEgYIIZints0nlWmtMCRkEUk12rVYMNlZtaqn50aT4mwDVq7OAelpXi5cgfB
mTT8ujgTt9XZzWzzGk+0wY9uZbR0bOppd7QUNDwc0rBthDAmnqdzqdCCKhkxh5V5
/21k8Yn7xBF0TwXxuS7w2I/FLzP5VVwa8jSTqx3jhzzXPAm0srrLmYcFapphrNph
jqjFR+xPT/VQIMlCWfYii1bmPm8E7xBIyMAjUuCdy9PZe64xoGuaDh4qdm//n/07
e2onHx6wNWo6gneE4mjUW0lpEpg2hERENY4j+ujus+32wb7Td/CHiPFOzXX3EuCA
MQD0IsVtkqxpTlr3eh7WUMJI9/MaTK7KAFwTg6bFb5D7fn4A8H97laDZtvefOgLE
OW4gygupAWLp57wtiWLZgCKv5OrBlfxnlxKZocVxD+b7469cwqx9ZlNlmiIXoJW6
MkhiNPh9BohPb6yksCvA3YVtDCkb8deD4+MFIZHlfSVA6RPVBllIhxi0pWighqlq
PXK+EGHb50V2eTSLg5r2ETSYED9pCk3twQWaQ1EcKNojw/Gq9n0Re3Gh+7EVIg3B
Zso57zEI1Oe7CGZE426KxiCo9aEI0nbs3mzJaItC+IPD2+iSQKoJ+0qX/7QVOQXI
jEq4Afe2zUd7goiE62FAygOK4OCgL/CKeupx4VS/Z5yEn90aJ8FwIOTvlL02YIeG
KZ2/SJ6JVURd11lNd71lNfsm3VyDr8dUJAqC5HZoRk/xg1iV2KKbQzW7ARtBzNJq
vyff4xZB6/4f2ksGGvfDfmGUPx75J+2Scaa5DadYhxunTCxRVosGYey053U47VGA
5fvDH4MSHKULPN7nN56rYkeHRJWqFLyba7eN2UnR2eWpoEmd5z6VSF8i/l6vTs7W
9SKiGfNPqrWlIEHprrKUNGlZpuzIMQO6eEA30VBME9q15JngFzSiJIwShwFZHleQ
HVlC9clfrRXqngQxLIiR/yUqO7cFDqFC3VOWrzCyQNGvgpE/zzOw3Czdtv2HDSpe
mEHJnzRKtYiVGr9kN5YPk01FXHn5O99vVcvm/eUYuCMSYuZaQxHBXek8KC8LmxXP
sw/P3qAgVYLsvbnS9hQcuyS2T+Vk9dPB1oCnWGY2M/7GUDYSd3AZOJhmOEv6KVMA
dpyBGZN8Ow7RYR73dfgATa09KHwWlAeOgwGspT1m0l+1q7NBKqYw8ElHXSuQ9Ys1
Y6oHLI6UIISYpiMZew6/NAPI9pgkHLHXZ2JteRiZB7JHEpULLE1V9F37krb0+mnD
mNY82ITsoMKO8++xl+A/pTGTZf0dNxgIxhEGxWlTYLXtQFiWNE8mnrzd/+uIETia
BF6Va6Ip/Sol+jQcV1RV9fWAd9u+gP1FXJ38aOrnRblnO78nxuDsaD3I/8F1OxdZ
BpmmGbJcT4C4FdyjmwyuiJFmyNiwvrtLC7aLFoEmtPxhOn/aIB1ClPKR+z/oju5j
wuZRN32KcIWIBE4z3WrOc61oBh80ZgK1YJN8AJLf+1VB5otR9LmDhGU2yasAbPvy
w2gENHb8nhAKH4rzyvOgZ8omQanQLUD+3wmwWscgqCL6OLRV73yOEERayqJz8C4n
QEFbZhQYTvei+4uLjQilXDVpCv72dPg5bC4IZLcw0pICHW8yywBvYbywyHnvpGJT
Q+OigOoP8v5glTbfRMDqOVeMnB7TNgB00g+MXCus5S5uS7BjIXU59x4ZDS/IhDLM
M2PautkN4n3tSWTcZhe/7h8ZLOnrnidA3rk33m6Mdpv/6h1rTIGu1CjzR6pTiC2J
aTbgH+fDSRgo4Dv+HJopQD7Jv7ypnkwl1p1kYavoPfK2SbWcYXRYOgfefDQYOfpp
/x78XvHIeL38+jlPTow2g7JDQbUmisfk0XSQ/kAA5JEnu9y1w7H3WsDRY1mJRkyU
MaZraa2yOaEXGrBw7O/GifStURH25m58bBZLPV2K4x/4OdzpmBpyacQp0ofoKhhW
tOGNbnUJPInLfYTS236vwVseJ82XtgN+/kCVNWxL2OjQbTU1Aft++bFXTaze8vH2
STdJakYKykd2o0mpXGOMNZTOBIoCMy3kcVT/aZf7qlPjAGtkkk9vnYP1WoKkXpvx
UeUU40tvqKv0uyRlAQQ4ydDuVNYtauG8IH1kdABB3uDh4hyt+1DU3Fk/Z1Hq4Y8/
QDC1Yn5qr4hPpouKXEDGenrY7Dk5tVXPv8WPbnnFezj0QmrjXWmWit9k2Sp30OEZ
D3GeiuVebNE5pJQK2lvachX1r+JTOpfkfTtr3N/dXurXP2uybH/wjrv6gCpzc2Xs
G/s8fwp7kxoAVxeiP5AdNcKmNnVXP02wZUsf/RZH2gkzpCNzSzzRC5/HhSwKwTrT
heB2VwzMHfQBBgVsm3eliTOo35ec0rldab26YN7JbYNpdplRQg2XGEG3d3N3KEwT
EsBeKJXJJckc2LPr30DdpqvOflV3KGRDltwEr/kEZsgOrfmn/K4TI86V8spRXRl2
eTfxKu2U/qV+wy1QzU5ffWoh/vaa821awl/FSgiU6DjuqjJTVdlmv3UHa07VO/wu
caGoweoPm7aCyndQVXJGsXvsyUsoTTxipNy8KLKdNf1EqeIiI0k8oUF4ebPlEDMm
gUNW1Bifxw1fkU40nszVvZbO6hT8QVLR7dgZEJuCNOiqfuOl1sez3PFQvCvXAlkO
2aRF7IOWfx7Y1/DAI0vZldJy8zAe3N4iV8VKEGtBFGQImG8UtaK7upQoJzFM+a6t
fL2eglR6Ds1xFcePw8PKDu6K8kFzQSDGC7D08NcCu7Kcl/kQ1jb5QeXjsx7C4m1g
ihQWd6hHQDp/7k0sDwhdfySuC92Od6RNHcGtI5f3T8Jyemzmq5UJECTZGQFrJTlY
+8feGPYvgJR+XiY8m34m4w8t10e9NjlBmAwQMZL8lUalELATBx2tEZ1ZI2Hqjix6
q6CpN3/mlccuoLi3aYCBqebdSqW63fWSYW6FrGMMzh9DEkZP+7qcPQ5vh0m9vm0W
K/A4TWOb1SDK95LM+xvGEkLVHo/BFTkozUJLy5vUmSRJrnsESgU5G0uy+pp2SHMQ
vA/bIZ4Rhn2MR2PJxrLOSxbW+qtcWjX1OHDczoHKuHWjbfYmqUhWk0ZWMGimWXLu
8qSGUUqTex51jvzdY3bppRGa/J6bG19PNubeoHDCbeWEO5bXaYEZ6Tf+7IEq7kcM
2h9ssHCB7RluALzxDvRq1KAyQqYtRl9jMsxH1byeMV+0JjNuIFiQK4T8Z1+KfR8Q
AuOkMNolzqiwUAPsE+BiA8v1lTfB1xqptFvbnNOzFB7ocHicunZQEMXl7p6VWo7u
XU9XSiInpiDWSGHr1zb3j7kE1MAKz7AvUTWcUdTKVnBbvXbD9ufxM4zvqM1Oqo85
fhHMuRwM/HpABsfaZXxcEMb+HF1SREL2m0V8Df9urf6fX/Gm547/iS8t7Ls1BBp7
t6RHW7RmMzPTNTDSgERYKH6ynexc8EnCI0e2fRkkPws5dkmnzZ3zqgxIHzfAIrKv
LTmTUQkLD9OIibdTHjLXvTFh7TAuEWULad4D/fsnp0xwqagj3wsgRSwFd+ZnpS5N
bYWIWyByDrNwhMHfrJw0SbZQ07fWtXzH2ptfLsw23A3R48ek7+2do8dySL2ISndl
5J6oD/THRAgBqdFBqSQZeBYjGjTWIgJXQrgNkjG/YGKo45pUGJT2+d5HF+Apf9Or
ZhOu807vnFHDb0gez7jpThqubzZ9EwoUlC/UdlR6xhtLrIXDE0lOFnnDq85X4kKT
xCvRbTqrvi9bZ30ODcQmbYOaanYWYwC1eewLbMgvv4ea6uWTLFrg7RxBUFU8nPKQ
V2Tbd0uzXz+EgOg2clOZbqNMkfDFP/q+Hz8mrW5e87rLXAJa9+zfaBKxQwb+jvIM
iIlfHD2dfnE42mjbowEH6SIMB/nxpu/N9nXreAqzhBE305HkPIgfdPoSUxazCGJK
CJiQlEDfqyEZZE6UvHmvwtmdDyfStn5dyO5Zg9n/LlfdfaXPWiGPyf9BDe1dV6OL
EAK6ZU/MolvW7otYt8YCE5pS176ydi8tBLt+jmMXtcAuWFnC/px/W/iYmE55WR+l
WErA9Uyoq9sLYxya4D5SFJZpvEPUTcPrbL17peawtLP3c5EV7hJnCOaQhNJnC4zI
3lBd/D0ia7v+3zwlQ91A7SEcetr62Z8ajC9h/pUiRvCIHJHydXxatuLySu455tfI
gUGQyrcd83Z5o75B9gMLXqWIFEyhHLPQL9neOwR7qwcl8ko5rUmiyNtJ3uaCDCtn
MVj6U9ENXDBBzUU2dDE9RsWAO6xW42Wn8teM4575Iufydn+dphuV2qQrZKOKyR1Q
K/FvBUDRV9u433cMwSfzQ2iBetxvSrQBA5XlC2/SjhE93O2QjfsBFl4q+T7B2mQ5
At/O8FNx7Y/n7APArq1DQbFezC1thTngFgj2p0QbLtvQs/vzaET8Bo4CZYP/5Uhh
RNATiqK6iWLaA/JrquMjuUnuVszrGw9pjBHkCfiG9kwzucZyfQBajanL3juKs8Dy
0ZaGNFf09cxMYOH2IL+8quksN/10gy9NWcRWUENf6lJyR1riZbdWFI3J00lIVqIA
mjWm3+rh6fR5a8TJGAQSFzEi4UP9G5KQe6kxeqeeBwmv9eWmWEjaOCs6JdthnTLE
1FoPenhxtovOJ2ubCQkrvG0hDLqXVODLYHVj/ZDJIKOroIH4bfW/3FdXqgBR6/62
t3J4JNN6y5WFMe7YMJPTia51D8LTOrhidRl6vCxEcki1oj+3/7FACEHz3zfD5tat
ZNZOPl3pTqizOFLOOUcFtUj4Ki6jURvZKFfmOtZ+XFOACQwkaQh205yciPJ87Iye
juWe70zD109BzJtdcubC9GWHsrFaoPMOetb1PFfLJc6mYW2s+xiUvo4k95gBQgPI
6zNp8F6SQWCTIhQktYjnyuqsUYa65tBbUS1t4sgYpOc17RUGUMbXB5GjjdiIqqfQ
+3IdpK6PmMBPQRFvgXHMbn+jNJA7QkpMpjcUsVBf7vYqEbG1IWyHSvddHwVSjFYn
76kaBvaWO835Of//j/UyeUsBHd3JfD+TcCP3PuhlxmSmGHPjgJOpkxrh9S3wwPuf
w6W6qhUbn1ImtTlMKiNtqoWRlIrK76h7Y3IzrmnQEkywXmILzFEKRjYsAgLKA7Vr
2ey/YDpnE+8HaYQzuEXIr+8n90BzmbK/zvCJ29tw82ocjvqWnWrvXXwuV+aXaESH
v1mCnUzm4mv/lHxBT/re1qQeLAact9YdPwldNkUav65KNvisa37CDrSoc2/BJtWl
Od/mEPTV5IOq5GBD2eOVpdmMc7Q4qORVcx8gBP0bAAqXs6YWmBCU/reBcAegvq82
TqkvAxVNhQiJm0uDwm/qvRvDaRsUV4JoZodpUdBHKB/1RrdKcLfBWdJadk260HAz
0wSPKR3Z6AmBvSUrU+Ivft8uLikzz4lmXQku/6NIhfnYT5XyrrHhJliiywTj5tjy
VniYpCxVeIVx3aRnwrbfcqNrj19AYWM1CB8Iw//lxEtb0FM0/D8SFIySQePtfPyu
3ZQgXWjdJCrRDgk65HMeilxdlnAY1Prp04OJBqQJdH5JIe1kPlpBcJUi7zJn+qCO
ysMBl2YlSyg1//mfJTFqMUc4cuNyiLTlf48e5Pd5x8CPol7yHWFu9PF9Vqjbc/5b
MS/fQhRQQgSZHibDQbpFnUyaJEQmEJZ7ua1QkhqO/YfHnhnCMP0pHMg+ay1XgFo0
c3/8RfxcAawIU2s7U3dmzXN79pJBaHiBCMNG2KvXpHn+FdeY9mdXTOrJzJcLmE5Q
ul6WPW/4P8oL9Ro4gLOw66YbS27JJbMHeXFalu9KZr96ZgHQAAQBKIPmFKMHEZNa
N44S2V+Edx5FjH0G+CD+tIkFTC2q0wfrUYp9MSM8IUJBZf4fSa8jK6MlSeLPXFmF
nBa8VYo07gvjoluljNyMPgcCBBX7AVqviPzZd7eyhfILfJMJUiaUdRq8Ty/fNgi2
JsMoDBY3JXWbiuxE8DyePxRgbyed/T/ohhW7EWy3EsEfQ1526ona8BA6TZwtGsJ3
wSmtIxEbIoFMscAgAqrQ8ruMDz72OLiYyr7nXMEt0MIOx6n9uhI468/BsEHCeATi
4XrW5lELmDN/UytsalsJJqBOg/xJVaf6rJliaMeK0WCaLjJ3P8i2zTMyVZn+gigc
suIj3VvulAsli4qmW4qJYPQj6qLbJGNT175h84OXuT7OrgULFB34qe4uL5vV1CUg
RyyKpu/iT0Yi9N922vdm4Yqu0h/f0K1112PjfTXpKe/iRG9E2NXhduZcuqW5B73T
XZL0gM/jrr/b7mJRTz/KR88jbGDsRMT6YhpOJfZ4OMfc0D4QbIfChSwdGbWYcXey
UAbMGXyC+oggrRizyJW6oNQSgRcb21sTcr0X2Qk4iwEYhrVwEoTW6hKGj6thxuP6
FrZtLZ6DyBQH3K1M1SkK/vXKtiBtNdQKipBGv+OPybJ9b3TsftxPBo+vifzbzAK3
QndteXuVxEb0dncFUW3GPWEBcsfRImOAg1EZ9APlPaR43lIRZxsC+u+wErgb9Goj
cZlfA6kv/jaidtEdzdQRHEzaZnuFfpBm3deBTbdrzmKEw78YRHBXmBLoctBOnjhY
msleYm3ZG3PGqcbjV9NvyjbKHE+XYeDUJlv8NpZ0eEOICi3142zOIp+C28bj4htD
POBFo+Gc/bMnSjifsnvJhkn+fLnr6tWtpfPJIjgSQnemcLx+1tzGljMECDtwQHPN
6mmAbm2N1HcS5bKYDE12HblpV1r/Eleezv6fO2V/HYCmhWL2hMVJSZs98sAqBA6a
nJSotfKVJ7Q5GrzUj+W8mpiEIMN1FOuK8oP/YScmrI74daQ/n8GCGC9nOvlO1lEg
+mjLnEr2OY0QONKHGb09xal+KCycMvA6xzLsclJjZ7dLlprehLjTsNWGFBPxI8Ia
AB+kNAkw87INjzDJGSdX6Eqx1E17GSaQnUPlH0CA6/jGU1gyV48hCkCNE3gqV6X8
aG7eZkucp5oNoEo0jGmTogvrm4tmvtb1nDcKR4JvUtddCQhkfDmzEv4TMlp8hPbl
ULthE9pPBDXKoj7eOMG+yVAiLcTpezHEou2YaYCyXcGBCAZF43tH0Z39XNL/G7C9
Ruh+WQ3q8VNgENudiA31NQ7bHvfRaQIIMdquMvIISCpn7dMFL8QsSAh64WZG+TEu
MIivJG6sR9U5/5A1r2kI5VuWvw6gG3jHjDF5Ncd/YPFkAy/EyOLYGn6rqCpF9rNY
VcD+zpWS6DpgNvoKxk2xK1LQwkcN9h+3/lzYCS4abit032tiMKyj3qXRL2knaNli
E8hNs5Oc9VwqQBkbkxUwxti95KEH0D7rbYLeskqYzqcxEG/hKod7y45hlklp7ppn
Ufz84cIkJLkfjAyH+aukSNXrMF6PE3MAhwfaOZEq8ix0O3tjSaBPQlTh0ReE8Ayt
riOKCnhAZaNW9EkGuG3S4GrkzMoRT/lFYY3cGqxDSDgRZE4F4P+zH7LDiVDVaAKv
lqv6/UxFpRy0jKBOVP0HIlXwp1DLxa+7hU+Jy11EwqkrgBCJRmnN5EbcGy5MVywi
pboyryjsJVwkNzot/yhyP5SkGRooSP/v3Szb8xK+LZHJSclbtXp1svgmsnRpt2bM
zk6OWgrb1JYdLIgZqC/SHQFHUCdjBYqf3oFg2RMUAMZ4UC/WKUoRAlYo3duYfzQB
Cv7sEaONK1RkfmvzvBCABBPa5el9u45xiDj8P02do2/U1EEBYLLRMihWwRIu1EZ2
Kxzn+Aov4qRBomF+IZAYsuOZsTbSJdPP0X0pM4cf8oW9yMPBEn6dpcZSRVGFIACN
+sqKyYTINM4lN4xYng5jHdiMObIMtQaYsAA7oxOn3g+r3GZdnVErnU+F3OCSSLLi
u7RXDA4evESOngxcrK3Y7Dsz8hV2sZueQ5jW6yKesfaWzQgv/i3srkeKphmG3oMQ
Sf0NDodn/6bsZHFZrrdFKm62oACbJmWTEFKgkyNWVBzBKHj0BqJy0NN+fz7ECEpZ
jRhbTlKgjpwgtJzrSMrSWy0cPcKvpbeTwATKOFDwNNQW0D7IO3o+aoM+YBZDm+SX
Kuxk25gWtPO0YvDW2jVUYRbzNxBfXlI8/yKuxBUUON1dVOuO1FoT93LpZcNghnV3
sQ9SPg4T4JN0zACw0tL9PhRM8IUvBIRE652JCvR1CMe3Bcr8DBAzTg8RQqXdOOmz
Qcr14+TUMvv3/QZef7zzvwPQRqqP0U5RV+0EM7FFPUZY331Q7sY87hESF52zC2aF
dbCnSYNyQpNfyKE1kLq5MnOBu75UTwHugmFeSwB4qezxJ1cAXxSuK0A0mvgp7tr0
q9+UsdRuQBJZTI+I3OJVVvyTK01Gb8JW44FSH/1WNu8DSGTyjt/9j2yhmYoKbQoJ
/iXaivwLXgOlBxbTxFCII3cDfUzfpu/VO4UUzowIdBgbKLP72tdoC2pCz+uJTOwp
QW9LI214GyqkHLE7FzJY4Jl5bdJKfsT8qz5YVyrdK0Sf8kIGthZe5ANN/7bRpR22
6vWjCkvdw4qDN6tZLNBrbwOi+uq8c/J8YrS7cpURKU1xHJYX9RfIW2FWTGqrls5p
/cbKtFvqY1gA5jcB43wWIck8hgU/ZG33ZHZHH3l4qxJqLewGK8+t+B2YOKfROahF
WdrRw1CzBbJNsKenx++uthgyYLxUaTFsFKyzxbbkIRDZ2H5mfjKp2oMBBBr2F6C2
ul/KeB5EUD8C7QO4ICU5ACrRD1FCwnmpcwqDWL0RIxyaPuN955jVvHZzkuY5o8Tw
2yDlmm6W2A40mwpU35j6ZrM7k/d+ttskRaAdtg5ThgbLSBIKwRXNq2GRBiipxSAM
ktYp0wpe/5YJp/2ElzvQLwMcpy1G6KnXLWHVYvxubUTa5M6BdvuIXRlJQjfaH284
YBAgrdwVHc14K7Ymcjz7T5m66YkYhMA8Hw7UVZaiIwXWQr8pdhx2oN0MGxMKJA8P
PyDDTi4RSSs9Taym4Db0hz8VqvGMzn6CgYlz8H5OOwJvQXN2Qt1usY474SCKTEgS
t3CJTapIjQ1Z4ZBFVU+j7CWq9J2Nqh0CnUGZCHAYoTyek9jFLQrkmYLTSwJe+YIF
oMvWn8QoYyolGE+UT04AMkDNRlBr0rEIy4qoo3lvsodl5e/jdQR1+K/MMGdrXXck
3+fJAuNrp4zk6+RZyidtpbVgufIrIXUonui3bhtQaPoGg58K50nfdRo6YxfJi/oJ
r0weFsCa5j6z4kK+hb/02HXTqGAqpJvT4GZdR0BHpcEALNodAENdSTxwVEZL1Dls
DkdejYx6pPschtzTezQYkJ6UwpX3CCCe5IfxiegAYjxrI32vlmLsxHN/3Argv1A1
hf0ykk/5fnNLv28xQS/YNQEEFRM0xPOivAg3Q7PR16ILYcUh74lUNK1WRhiBmVBT
L0guoMFXzOFIjLmdZXnyv57iZVfOOSnKwiGwUyPAy8zkucemFHa9P8mOJPLe55/k
ETix+IuKk76EXOjYrtB6pkItAZSszTDPSCspC3hnvpClO25iVRgpjk4hnEhtyVE2
1axs3P/WsrHk531TahlP3XkoYIp0l/3Bc2z1iny92O1D25UWYBQKEQegs9MPSw1x
VrI0sXlFYgUYAcwUQpmhaZwfb8mB2wY0enAra/cEukwEgg9tOtA2WpcKEhUve9W3
f9Xi+qPzLNfULBlBStO4+2/Zcaafb9UPpkIM/LN3tA2kM6/hKiWq9Vq26yf6bssO
c26PMeXzWQ95Js7NQkVB5B053Erajts2qMoLE3KzwrA0tjg6LtgJHXfLR20pZMvs
uKrKaA9ls6HDops4KdJ3a0T01lpiDH1UqQOl663iyNAaxsKObAyx3/ZavSUf9kwT
PVRlrcElOAy9wbwyHD6uEdPDePmK/RvqoOdjaiYda/rIhZR6PIaj6EEPxz2TbmPn
7T9f/67vKtXsNWsHJDmFklHzsz7gDXO8uBOOvx6m7ShefPlmCmd8Y5zvgr0ZA7br
ymj4pPPWWi7Bw6SAtwxma7EBSwlVMwF0SdY+tEePwz4W8jVC+G/1VkpR3q5fLcP3
SilPjIzgVGhoLKJfkL0DtAj11GEQi+XgnFqNTuHbOqy0PudflEsfquatGZcDaTtl
ZBs5289gRRAjEjFYbzHmUqM4fZiz9MKdJJSipgUWIMKMZEZnU5YQyEt/TkQIq0ad
5rfYZQUpQ6KNGIdCuGSdcf4I94DCim4yTM+4o7iojE0Wp0d0ZKS7/hIEoGQoONGx
CUNRj29B5gZnhw64O0w3Q5HyuacF5XvgWpKV35SQ0urgZq1X807BXehIjgpCROFT
ZEp7EdgCyeQhX5kSijiZdKjtR7lZ7ECx5C27BlVQsmt0m9LZptjGKDZ3IHrouTjF
jwHeazeFVvvaJQ9Fk5m4C3oRJBPZWFYj/v9lzuKx9ac0tqP/dcDfVZJ0VrLG/v+6
p0B4yJdcaR8qSrI1IBDQraVxv8b8hkRhoFjXP4K+91v8nLUlKokwJLaoicDdLD9o
JdYgt9V4lEZgEd9i71sNp7C6Dn4IbZ+sp+vIZNSs9/vceH7FQev9zlFewJ3F/4eq
KRo4nWQNJ1YVDksZqtE9+ZrYsSPLMveDmCjbR9z2RCMMccTk3PJBduMkThyIj8IG
iWcg90gwI0/U7lPgMhX3/WEgfpJcz7lbVWWuyhRU1Ld+lGcZTcZ7u9rRUwF8WXDX
kq6JmXck50oeAj8i7TklqoJEXgkxZc6wtgp6+FB03Ofob4K5fK5WwPWOf37uUH2S
vBj3xYB8F+PZHOP6SgZSaNte251h+5qyrYTSfkkojYhxxBun/ldX62lVmvnx/JeR
xlzzuxSCRHQjUZcCWRyJQtAZxAKEK/P+tTOJgMsqlwDDljZ7tmjKHAFyz5B+D/wL
8XdDoeYJqhbWnDpJ+RKTzhjp2UWdsoHrMcYfWmYC5T66+kxl6ZfFAVkTorienwVs
F9Il6Jly4vL/jgF8JMc0SBvb+wj/MK0Dvrvksez8R4++XzoKhqYVDe32az9x4FRf
5SErt096PkLLfrL+z/5GCivv07F0oSaMSLYTqVduWV8d2KZPjlCyeZxDEvTWO5BP
tSX8k2MsLbmjzkLElQ/M2IDHwT3z/poPCb/cuDkCMKY7hZtWZ29kYHgo5V6KgZvo
bRrTqO1FjsOXGU0rJBD9HkxxbPznKAVE3GFj1GSD4JIxnknyhHPMXP4kO7QMhM4H
H88chBe57D/vOOn/EAcy09G9rXmIx0pbz2r0G724UOO4vGoEb0N81l7TVdlOYy4T
9qXiGIKIcPEPhuIiMGrc6PtsKMQ1osvd9Xll9E5VdZf/vsHaNB3XzCdhgI4DGx0N
0JCdK7TQhm1VwhrZJX75M6wpeh5sfGq5sefQB1IEQ0/Wzi2W7imbYqDTU9SW+kpt
XjnBw7icU+BEwelQu/FhWLozuv94ROwVcjuHyt0Gi0LFXoq25JhvzjoXkbuoy8ow
Gmj3FNdDvyHKEaonaJ9BF6U6BJnv+M8JUqKUBVzQjqeEq+sDrsuSsmiYvFJyUMhv
DQG05C41P3TjQT2pvqJ/DLF/7/tUS0y6bU1uP6jEc7nFhsyfWb4plFJwmkY5taPe
QFL8vMkmeIOaWenHdu34tv53JHRW6dr5FLjErgOPVvYTN4JBKOu1bC0HNN2/gZXP
ou/pZhBWAAugv9+poRG4ml+96gTCVgzrV1x6vmgqy1nr4G3j5FslBYNRUil3hEaM
LvD8dhvLHIUCHZVRyPP3nK/cmBcOJ5yFUYzVMvBOmvartXeSqrsuhza9CRVYL/g6
/9g2X1MR7Nn5mqvQ20XhkrSyC7MeKtp8eW7LAFzlk3OLCi2aGDqGKoJ1vJYQPiR5
/hD+TwS6YxzikPuGpYFSn6Af21oyG36CFhv4XJFHS+7bD2Mv0t0R4mqStCu49S0d
sr+n3FpaxCE7lyBnCvGfFQy6AB1KkgYXWWXk7pVVBV16nOqitoKM3vY8Ll5KH8/x
WW4vG46p+enwKpkCF55UFICTswvSR/pvt39dh8cCUmicvCY95eUuZAqqBKdQQX7o
4JtLjK6QEuavqz5eap18eUulZwE2DbYvEQBct5dIhXqi2I8o2cqH+9HVymCDj/g/
5Yjf4S4ZinYBizr+m0ErghO8TIgI6TX8KxrYmKZhzBEQIdHvH8NNnj+1P+GElfOZ
3sNAe7DnZpmHPGoOmVE40p0Mng+L71WkxjHHRn1B71uzYf5ysO6P9oz/rtye2/sd
61ZhhnTEDw8pLQU2NxpRBSaDZBKr8oPX/3BuN4YZf2ajHNyFT2NRTNkhzp5oe1Yc
NQXJiawWJLOfvg7ZBv3BOp7kgwtcPbRWm5DlUtAgDiuAVMi6OevimPcXqYaTo1K/
j6LMZEATNb2gg1Wh5U0crz3Xb8IOP/E3W8MMqmcucO4apvtWFmWicxwou+m1YG2x
qITHs18TsA36iYL5b5tgGoitxBC36EUB5VQ5sLduI0FitZqlAt9iYKWO/6drJM+y
1KKUx6ZlZI+Pwfm75qvJRZlp1EsebBajheyylUpNFI52w/hbqan0CdFGFk+HrGyG
KejUtwBeGTYsCKxBc3cGwtkEvKZVGEHlPoVjgITF/Ht2IM80cwOLn3tgPp3LLVoH
A6H6XYuvMAt9+dJVi1im8wFxx/DhDRko9YdkMjUglPf6T80iai6VxiIthCYBGegq
tKwALhkr1POXeSvhWYWSAPV+pNIGkywbzKy6NkcqLSjwDKoRT3bZ2uytaKRvYgFM
hrrN5B/8TPkJkl+KjcIXD2UFClLvPmsiOcrSAAO8/CC4jbqTwQKsmRZSHT2jOiYj
8Lj8jmCbGrdl34mLK07iw/7zgVaIb8ivneHGpOW0t+6gQppddJ0RO6jeckBSruwN
es/0TYdZYnaH5MONnG5IzrWIk3pqGbbWULHATaVzGlXWtDB/DDzk1DHsWqtUJlnV
u08wSIfnCLL016DzBpv1Q/fzcmIxMrQWk9jac9bRC3tScrMwp4O5RNz8gAYeYJnG
dFbopfyUDgaPYfs3iF8wOYY+/4wb7+gka9nBWmLjpAii/cYbN4IClW8fyuIHIqpt
UNb2uCZhu5fhazh/BWNQatxlZBJdVNiARzwOKG8ryO+zj4OAgfCsvz9GKohn15Wo
79ROK6BuEKSHwPsw3JSAijI2dAMW8a1Vd6E7VTLx2/lOR+MAWG7cE04M5nNZs/0a
EuOnZz2d4dmlJjf681OwkoL2c4OmXi1v7KDvGta97dr4zU1GokZIY1YBhOR54jMo
8AcPK8OwRSonZYlpC8ULR/xP3qYHfwnPcDVg9KtbXQsO6wcaaIk6lbG4P5+VQeZr
SmiWfKcYe1bM8wDvGiqscTHejnBSJ91zihFRBi87yv3M/A6fIv6YBQSWlo/TNjMF
O2olP4rgxGriWA6MRpKpMFoa01z90JFcXaF9I9OqbuKu2b/lqSVK2qeqENJHzte1
ATQrk2QbieyVyIKQpVgADnwv0C1i6XasbSqutsQztYeMjHyvPpLYIBMCHcWG5CdI
B1Wq8SHybjEazm5nRbS4dzWsyQgRbviV6YdiEDT2Hex/ihUUs/Zk4q8kyiT4uQoF
tS1RHMSTG9kLy1eWWa4SfRs1lZgzau4DfXgMP27aeatWTO5C88hDJHW8lJdO1a2B
XSZonimipuN0pVFpJO4BUTAaSFHZX3vbFSFUAwV8z+yOKuHxAAhU/ivdaftJqSYl
LR1fltw7/gb9KQ6pljYq3Q4ne6EmTYDEE3CxICxU5SqScKidj2x2GL2HJ4yz7JOv
4Hp4z52bNimbyPngqmpHDnCvHazsCc8RUaW/N7eVfe/gws/EPnjJ0GBqXsQJ7p34
dNiu5EzX9QGwk4SbBdHqWm/e/um9a6lUV2Pb7RCBK5PEfAckRXsFcV126ytFJ0Xl
Zhh3K1xZRYqlREI6HALVWp0EjVIQk0koHqQLfPZ2ZO1XgeBMqgmznfohB2bDAlC9
8jx1R9/59Iq+mqnT5dtr1rlIg4eiiLn8oCshwy+wUZTz9uDU8WkBnS2zenI+qtMK
1Tef1P/Rs9ku2y22NTNxOuiSc2grkXCD9HZGrS8JPaIpIdErJFw1bTmLZpByu5QI
H+CqI0RAAl6t45QgdyS00EpaQMmgsB6l1qTGgrnf6y5fSHMLfhR3o28sW81AWODc
IYrWAARUxvr9EtY8SqhbS6O8SX1tgWhDoZ87+I9omItY1jU/iMXwP/CPFyQjJL+c
EFJaffLEC9IeVq2hAMRo9lQdtKa9WYBzzW7GvIJnnQTmrKMP3aR/dxEV/7E/qZqZ
9TSC6Z5Jjus0KzYU7QM38i6A0Mqd//sZD57FWB9oQEI/g0HlIJ/0EdGleUUg+/DY
qLBuega7pfYaNa0OXAf+LIMOxASe/TPrpJCskZYH5yjOr9A/l9BJGCYRLF3Y2mWV
APy2FBvbxX4Fhvw75gig7s100TXeh8x24IOPKaL9XiWpac2yTbsXLF+uiAasiruW
kKuKPaXbp2GfcuKswS2y/mvU48THBp4vRojsydj5F9JczJyaJ04qc7BsPvB9QL7B
mf0SmgfXEwDjWgCAwIoMYYcWMrxdpoFuqgis6p0NFeDiDva7ER8Fo5YjmeOMceEX
+oB9oDa/JCVvn1e1uQbUlMESJEe7KK74BGt7ezxfsuc9bcnn0Euw/1LA+hs4Bm4R
ESSznh2gNLkVF9BWTaW5DjWyxyniCaYw00YmbFdn3jI8Qi3n/nSIrJvYaxlATSVx
BKWduTK4AHX/xWLWJBykz8UhWb0VUkAxmYjeUISmhcyIPBCt0vEpdvL2LcJ3LsRi
zKr4RHWPAGKZOY8KEe8JepCCvRiES20RmVGoph/sDoX5wynlH2lQadQhT6VuF0k2
LJ1YNv+sRiyUxo3iaWGjSk0v0IbmNLgxO9cVS+S6P+Lr3yvO9N6A+OPwOzNIDE1L
ZCBcpLpZFxsIPnLnYezRKA9WIvfZXNf4WKVVXArXEHxAoWUi1L52dCQ0XeFGNth1
AqV2vkF3u6tUnGtPo9Nk3J/hvsruh5fxWSfGme0G+4+6H5keQSXO4JgEqAIKvQE+
wZ6wkMtKnouj1ioxRxOe8U04uSHYOQ3zoMEcLcsBaQuwgMHgrUzeUPwntPGjHe+G
K0AkmDRAiBfu0rLk5SNqWzFz6WzHWhIdulMBos+3SoajtLkzrTPeHeULzvVVdiAS
LOWEmA2nBWXqFlaQyMKxdGGuR2VSSRW/S+EmeoFqiV8P9iJP2ANji45FHx/Ci5Wo
6EuDKYeFFOinX2HGB5mTDVfmuVQLoyq5koTP+dEqgmcxb+4V1harsRHI1en+8WpH
rrxE1LSoRIHp7dJMideR/X8Yk0bWG6iq2WnmNsNOOZJV9FNgxK/o7qTv2KdNkM8K
jUy7IZmAgZW5jKsxjhQlXN0uuuLsHVBVOaRQjlSf1H/IpKw222JzJN4WnOyIn7aI
+BvTItnwtycAhz6smVQD5NSFZBIDFjS0AVP1HGkxqHPwMivX8kwh7gIe+tGaSEpo
Kf+pbovq2jdDBJTH1hLvW8CSM6hEEkuVB1xZt7EQsEX7GkoTfAMJJX5woo7rMM1d
GSQpb0hzKAIdfNkI7KLhl+MBUbD3PQufIAFGp8nImh5z7lmOe+b1soVtsk7vkARU
qD0+2EqSyhZ+ziRRNNcw7wvgOAe2mCAbDmc0ehV5uYC6Mu/76GlYjhrqWqd5123p
e1jKbxWLVSpRzri5vPyQwF0vinlEzYdo2cnub3CHaO9mCg9ZmbY29aP4RlVwTid/
+lIKtFD4wO7grHSOoBL5hfd0lpxYMj3azK8azIwlkmQc8StVJJT+yCWJuII3536g
0HJ29UqOTspS07lkBdpS6rxXbqSyrIKyLcKdh9U4vglXGt0V3H5kBoBY8HctVhWf
guE2IYKqmMau3sQJRE2C601DWAqeYMLp1Lvu5ptHrAYSNEmCZPWW2G9Fzo5Sp6Uc
kSEeHbx7xySFG/+TLCgiODyiHjhd9aJBVdSBGyEhQ6Zv14iW0ritUJ70micpPXwZ
ScViZMI49ZB+uyaC+694bOjfyV0+oIrG1w7oZVXF44PVuc0grfH7iy7ZgHY/tJcf
2+HXeMo6LO/GCGiRW5hoQCF0qptZsSXAwMfZtD0u8/kKinskPuBDYoTTZ4YtKEZS
vEN/in90a2lHA0fQat/tbMaY9ZSpbbuMXzZtSjt7C07epQy0DiVdRbRBdgOscTW5
y9y9Z1eT4WL5TWrPo1Um1+NxhZFDEDuofVuMGmqav+kmI5OU7KdFsaUyfi9rqlKo
yxXLH/ZbBpkcbKfbf6EprUpKR8R/W0OTCi/bPI7NTJwe3yyw+1aVmnDG41yNmSTa
M15q2i9JI3VZzho+indAyS5Eaenxt+MKSC4BjqDIDMflIcaJMmMh6oDsrrU6t5cW
ydez/MKq6dC2C1g6HgtuDQ5bqHxItbH4TIX6gpBznMFBOTC13ebgr2Kr2VHbFuSm
c7gD0Mn0VsYTC5KcjFAobb8oRMexUFjgIkIqP2ZhSz0PJ+vnD3/uExlVPIbI0EC5
8hzntp6+O9uA64+RFZ/bXfkkpNTptQYBgb9CHHGHR2g60jLj7J0ZY8JxXtM6d4Rn
84TCeG9fWS9ry6+G/36YKIeQcU6ZvKkPH83Cz4WmDKZiguhZc3AwRT8n2tcsw3FL
Ny+Z7j65WoQBYtsDU61mxrs3wXPdRtf0Plg/WyoePI0PDP2VkQ4t7FcGs3b7uZ0d
U0+L4caWLTvB9rkYfkMIt852wTlODQCXAXSliHKzz1n4/gso0kzbNU9Yql/0P7OS
9Dc6sTTy74iA8ckL5hFy4RNqZDvi0aiPe81ndy9EBwG+wVbf/byulI52PC7QC5vV
EGE4lU78TTShXayt+b41ogtQGl+CLFKiqkiE3eGhPewRYknCQmK9IODGUtXcoVY2
pUs29HO8i2QygfGXMEj2fDHEASTx1LeobUyoVSe03UnXqdue3pH3E3OvxQKvVkWG
IgIDIhid5wG/azKvId2cQY+q6GGkYi0+ATIoeepKFf6mqe7gJe066JNVrRQpHKR8
reVJ1yp3//LeNDz7909Oa8GCsGh5wXBqjzTIhNxV2T9InETiulOfT5lUqdPc+0fB
fnET1KvDK1VAeRi6p4eAmTta2fWaN5dsq0IXAs0DHeZM+B9JFLZbdblo+OpdPQnY
FmBBh9j02+gpwE6eabRLnx5zwCiISc2qrdgMSy+l/I4ZcPA+rU3RrqZgAVzd+1MR
XTwiTnPOud9C3aT5a5UhuOZX3sjw+8ZTztdg0lQZ8JqUHx0I3bGA5iNeYMstHlwM
yY8EKifwKmYgwps+QHUmm6ik2Quf+IrmX4l8Bo59xIsNgahIT2xz3Q4s3OuzDTOk
IRP0B++NHeEqM0NODr99CWsWfRLWSAQ0Vi7Pflm5ioFfs440ipD/6spcFpKO4n7u
KpVz9k4XKrHdrAQQ1xI2xp9kmhpKax4jUrp8P6SVDq1fUQUtoAa0U6i04+pkHG3w
5jOyHIaOnwqx2ydTDZHcn9DISabXOBhG0XTpl+84tNkvgdwwsuO5XfRCQ3RGT/Q6
i6LBOOqeBqLaTIN34keCkaRij0XONFkLOgtVDikSkQKmQr1ttoXHz8BRzXWs/V/Y
hWtyPkLVH0PDjMZ5IvD1Bfv+GIPLqmEggsYNOZOMvPgcJkhpz/TTauHk0G6Ga00V
Yki9tGuG+4CEdPgbuzXBIv4MBYQO6P1XpAXnGKgXAmObKrYokvaE9Y7MXnKay/jr
sIpypujQEZIwVuE83S++3ASwVuBF+3IVXuduKTEhcAmvljMFHyAjCqRZ/g7JC3lm
NTsXvuJ85e6KfIDkrcq7CETTCZ7yLjGJv4hgkX73kPSIRJWPSoiw1bgt0uaHUJSV
NXP71IGuthHCHBGhKaDsGSjv5bqVPN6t2Xq7r+Fnz37R8oWC3d9GMVgMpVGDzUaN
FJ00tmd5JtVn2j5zFk0lia3pNmXzhrulkBikbVIYqzc9mLCI1G/Na3ir5WL6dg2+
BcnYsefX6A6XifEzhfQd7fwBfLeUgmIUKOl47Aj+DRlIcSJ6t9OutRyo+LeJuBQk
wu4ficw1yNv+5lEU/k8a8pluBUQU/GkUYzYHIcIdyRRaTGT5Skf12JpJlPe5X++F
3ZaNfHJg1pVpgK+x58fgdV/XiernHPlow6IIdv7r9BhrxOWxT3buoLVY5DjuKJEd
R4m/bWjyko5FB1Albbm+g2syOQGl15hPpCLzKZMLMxJk1CR/6B0gHTPPA4G3iDC4
Q5W0//3IKFD9ZcqmGdbsd0Ns46iRPGFUdYWFeIqbfCjTb6ReaIUO2G5j7nz2KnZL
nSQZG4I7N0aDpzYEtOTaqR/j5xHCTZGKE3HDHnGehVuIO5UIsb9PCA9E+NR6oPvh
Smin15sXfXmKMjlVV0u5bXkJZxwa83qWJo3EMz3AwFOnW/OgkN10CU+LOaE4+Lv4
ZjmPSOOSQEgq3QOFMFIZN0JkpUXbJIWEOmicDysRmn9NDY9atJvrE8SzZ00/sbeK
UCyNS/sGZ+/ai4ycWMCvLJvj669gjYdLSEA5MnUqsRTMDI0ihPsBDsu0CoxJz8rE
HvgW9y+zV+HSjrnlvlx87Q7YyBSCXyEQ36HJ7fcmkeGBAAiv1nYCCNRMeK4RLD0E
dLC3eULgMyLBERlLkWaAz3nZy0DBzzN8Yk0oGFvzg2rgsVq7ewVNHp/t6xPXdX7C
4LMIdDgk+7HCm2JrBGB71DDxA9r2J085mE47GSEsn2iIa58xSGoPYI0sN2Szmkg5
jqdFfk5U5BMQrf//app7YsIJJ/ygNNYFi+wS+0J3G6MWInLp7VYoAmo0OzYNDuQ0
tLh/AWUHa/rVY6od0sWQ99P1qoNV7k7FqL+lSAlTX9CokVzyhZsnsIa7GF+NTLuP
aOrDPKVp0rATMvPnn5QJBnXdJlRZrEgUKfCzLGIHVCuuA4Ne2YsLuhp7I6LLZPnX
3ejYwB/KCC5NoBMFLCyc++jwePm+F7JRQVZrGgzUjuXZH9ZfXfwfXNaLejbvkzXE
wc9mjJOhAWIOaSGLrN/2VebuJiX0oXcYGJQogNvqSHdGOQWML2H/fJvXD2GHDZSp
fc0TZF7t/UbPcdMrTre2Fqyfh5CAOEQckRHCYCQEt1A3hJDQ5eCTBUen/f5zVpi2
thp5pugR9lWY7hblq7p/aeqNnpxO6mdKfUSTe/v+s553dLdhc/RPMoH/cTJnMett
qP3qVTb4Ib6gyi3+hq+/nGOnGWIn+TtbGZ6OJ76ckPDU7jyY1UGtuMwHVUUm7kir
JfCsG0jMx63i6tpHco/pOfV46WzCXpXAwt3e5DDwC6OsFB3c2cJBqQifa5xEF5PU
rBURuytnB0zXi/CgkJ5yRiCrdJ039gn88SwrwoHIbsnZgv7UV3wmsC1zpbpDCXII
usCzQOr4hBAwnJcO1izqYFdNtaLbiUOPQZGUIqa2K6VpyiYFlrJeeLHWsKNI9yhq
W9r+np6x//l9dWkPGvJ5gipe2cRWxw5gqCFjJcQEVyZ5Z0UembPmF1RVXS7kP7nR
AHHqdj+zvNvGpXUcIh0bX9BZFKLWxZ2LWeQ6XV/yGbtWHJ9DMAOnA5hhvH0UEfvX
UZyJIMrpl2ZaOrBPj8auKNxqsKdkQrJHWFHnTn6e2oNbuud9Paw4I7fvoly4qWHd
3AOt1d9SAG0Mox1S6LHvhNVqrcqrCgAABBPmm4GHAapEbplUfqNtXljCt6xXUs9f
kvvAv45G2pW+kQGbjhkaWts0LDP5UDvfs27nQJQOPiYljPWkAmEG5JVnPE2itX4B
4AOe0D3akrItc5ahSRafWqxh2ryUhGp0VuiIFUTaHlBy0pom9Ekri0RdrYr1QEFg
oETudAiC5o2FDcFBd44YmhKMnnc2yOewAY6oQrmGhCiNlJCVnOcmpVyZC1tG1GCw
0RkOKxhTf8XNJZbv4pqZUKxExQXUtdBEP5Occ4d9ltrtRMxWfT1n6/lgEYaK9U4F
5zs8D9gSlkhf68ui8kBctwmW0V4Go88SeUN25S7yWc8oWUE21CxCCJZ1lxfv4YbI
NqE/+1pXdMVVp5TXsGf7lhGNkFM1/PSdkVEPNoEnO+mpMO0YOBymKsGT7KDc9kAx
tEUxlHu5Wu9qabNBS5SnPQx6GIo9ju5v9UJEAW2O42rqa/Ua2IfIkk9l78DiC2Sq
fthHqG5KJpsapD1mOJ8/6H5N908qzq+XwmyActR9BzxHqLL7mCWrOLatdgWizaQ9
JKdc+G3tl/I8PeUT46YBCgfP/6dA2dtRl4aUa/5o2ejEV/bh2hnuW6gOnQMyUf5d
iJlzVRSY8frUZo7Zl2XLtW1L6KL5mlf2tCddDaCYTfPWmBa25D5jNzPB27MHEtHM
r0t5XFOHfCggrYZD1+krsrsIs3dGuFr769lTOxY1F9lIBNfxRFZZcQcoi9zNHEtL
1WIV5kvATp+CF7U+/um/IqF/EYRr5U2J6LFvgOPt8QNYya3mVBgOx2uHnGOWVILh
0oJlNCB1v2Iy87UBOFG9l+VP8/HQOdsKkHGLOq+vxIdwww3jdjqowZC2NILru2ZI
9KbkmnuSrb6INAtN4ZKv+c1YfIPgL5yWJq9ZTgtOISEG4RJRceS1e1uM0JVZu0YU
JVuCcDJ2QxmJECdyCSeB+ML16/y6dCrZRQBWIkLrzBvl/gIjyc4lokkrNxeupNYV
7yYHRbsXVBXACvH2cBYySp2XlIDEk2AUkGY740BJVkDq/8hA27EtiUrAn4YFB/m5
eESPyclu6PxKOaG1EGTEnsfWlwgcilQZGoNtrISk4qgeXkc7KCq2lWoY6KB/VpnI
YRlGxjfDL4axT5H33tmA5pQOZSDVT97SMfKYGQ93Xa3qtQYHZIiEPFAfP9Xhkl53
e8gAIRFpL4sreGFZmNQkugfJSewFenfajiBiz3U/bhJ/D34MUuqFuDGt8xuGD/hW
1OInSasbOThQsBD3mZ2B62KoAzXP14Uzl3581I4azsfXPSWos3CM3shALAg/qzut
OJf4PLoBr8Q3y1B4YCDqbY//GD5W/4qtp7Wh0RxEslABo9DutrS8JRD/NcDLEh0r
vTljpt4QhRfPsLY0D5TNWd/SW1gBo8OLZJ24wylVnoz/K6BN2SK7oxFTXlXgQIAx
c6e2tA/WALghyzQf9Z7j0bu72/oeTu/N3lj8uSGzKQsZa67h8DGWVazWo2/kOlvj
Y0t8X6OVNuBJHBSdI8fbAdN5hLEJUMS4v/3tgsmSaJ2Jda3Ysmtn/r3qAgACbD5o
KPsaYpg1ZtOp1I/B3v/+HuSpp/1JDJvnssvL5nzlmwpwwA1LiZ48ORvRs9K7TJxZ
vS3D/sDm3ZK9vwAsHMlV9UBKbpJXX/FVu+B5tSKT5KJvpCMvaNdGcZmG111Eh7Ca
dKbu8Uk+87H1+Qm4arR/5APMiIM7rs+RGZEz3XJDlJKdCGh/LrSCfheF4ohO1cAp
8Y8xK7GfH7psKQs4yrkutwKt83/Il6z+eSKQ4CA3ieTtaZpDAbmvnGvOjnvDGsTr
JiQ1pRKAQDS9FUb2sPqahBWTShwCiNjNs+UoEYNIlCh7aQvQCsqnZJtSEgBKj8V7
Ghfy1Hg4T+NTI/s4Y8bXORdtSulk4iMa5VvHC5mvReDcNZNxpLxQBeKJmzsbMh+m
aVEdaY0ZFm0/blRb3btZIX1NqkGo989TRompaAc080AmpBvu2Qp20qeKHTZ0Qeub
JRMQAGD/FPJNohMKzkZXJmUOXX08ITfGKKTf/Q8+ivqFg0uqHGwUnm6HdayvcOC4
fEdUBieE7J2Dz0428ojB5GITn5VLfqZtY1JwbVTkGP6lT0ZTbWf2o83fg2YbL9k3
WmCln1NgBr9omjBmVpcyulhLzV7J+tt3yRn4W/YIXu8mhPJWxCwuxNj5ANC0/5Z3
eAlNEBFiyDxtWFnoGApntpZ3IC9HdwWQdeQpBqZG49KAgvmujjcfgRthu3xbmj9l
XgyfSp5bVeRWk+zuOsRo+m+xKDAQduFz04r87yi+UgPky7S57Tmm3WoFRUWPwXg6
XtxAKYFrmmRNVfINk6ODnd5hqM7bgdoOmQZq9AeqhRbykgQuIcfOg0mXlv6bjL55
OkimQmEyDipPxGTUvO+vynSc3tfYk53bYnT0tNYL+vsbjsA0A9PMxGu+31m/Qf3w
QWMcn6exeXOCHJMGmQZOVHLmncYpWw2CnNm/Ony1+5x/uF3mSrsGfc27UZ49kOof
5atnwBOGyt7qtthHtxbQsFdLX4xytY9R65jobiCjzElUco1PXT/PifSNoAVLLiF2
3D24ilSuPLJEKfokY2LWFoFHdf2T1yJBQ2JCrKjz1IDeMIvo8ds8HeFmjhYInAgt
92R2tG/XJN9y2KfLdCjt6uhVHSdchDWapXL1vc9t16HIDsoI4Xy8n8RknoEpkh8s
SZPp0phszBXMdjLO2i4/bzvR+nN6jhujO0DPEH170Aw6E5zTmel1qkZaN1kr9wky
509d0jxhtay9bnIQ+kLr9pMI32A2PT2PKisLYhmJDEueC+mEUxoj5+S8obGRonTI
tP/08ZCg67ivPdkax3/K/wQ1a0w00+6piJss3fz93SdHzxWnaaEe93pO1bDaORgO
RDgx0ZBnsaB59MhJPvl3N0JXk67M0U6TeErRrj9+NtlZ3413SyXO3W+7SgLBUZ3w
wTfn+XPbkMI7z1+rkuVHSqXrHWqPdjeD9kZrypEqiiRaoAqH+ojI2x0RfdiJpa0/
tvPWfRWlBHT6nQRNdi6dvqGEv4t8kcwyNrYHGZTDDzXmJVKuCM74GYFqpcyUjzLV
uEjeMgxe63YnKXT6CfR8UFO3vdOBS2gZiHknBGhbD7L5Z5PyCkKOQTbZpJcKzRvY
d1yhdjrBofyeUYh+owDfaSe1W4M1puPtEaxcqKLWMeH9tJEuj9u1UY7OHE0nEWSH
FMbbZnUTAphBoMVgCuHtx4tZapCdiJFtFJoq9LJ3Kn/IofUv97waqWbaVd3QACF5
wjfbUryGV2RD4R9RxZNXu9UH7O6an0mnXZc6Jqdm4qaNp165+LYtU1gkyUGRVdEh
TDIdN+UUyTo68gCUjJquj4eyHNmYyD9cpJCxRWbcyVzUZ+SpKzGKYOhYSQiqWZ3t
9yT6PWNAn/2223AdDlTsUkiOVBxg7nLu3HMMmjoPNWDUlhasVEiMRzjynEe0Olsh
nSoulgN9r0UoJ9zs5YHBLtGzSSpzzE7f2h0V+ZS8YZ6MhbGVZn8vF6RriURRhNDw
AVZTV3CTTFy7BKL14lLKyhQ4mvKL0fBuC7UiMFzCvTVuQ9Cbv4BaI4tcEWIgu6ME
7mj8QagoX7UBF+SJmPCerqJJpM+btcQPHSZTe1NHzDzhwlznhb2/08LEGZwSE2nl
29DA8VELYEu1S71LOjn0AXTInxSVIzER+2Zugd0hVk21nDt9ksc+zTjPGUNotMP0
Bx8KQKX+uHeSVVEsJ+9W63vCIi//R2mMzqOwXPHwoZf2lc3sTIDcUanOD6RTq1tS
qEyz3l0CugEaPkgsa6XkXcMZhybZ10oLviCLZjbrqI87GvRVxmbWgU8mbzZ8SF3J
SSqnR4fFIRtX+Xv1WCPt14SfhfoPrRF5rlM/zFPv/cmdqZiuKNytHxo7RvFfSWXd
3z8Q1d1r3pkgl2AKGaGdbyvwxFP4VnBNPZESlIjnWeTRfuI5e39u+iRbXRPDdX5q
OdtdcEQUPRB+1sEQGRg9qy7v9lm20VsZRK/wIM5wNdXtN8LXM5+vppR323BxmBLn
Z2HOw3HOahD/aQFOfGzzt8edXOamUbW0739xK94W/j+yg9kOD8yzsRd0c4x9B0Ul
phBi1FOUVe+gxoH2Zuj6pcOMtPFJdq0Xa8tclclKN3d00lhubMlQlxep6CxtnmcL
XGQI8iGKlJPKbOGp2j2bm1NLQBq00okVj/s7FMvIm6JfihHLwTN+jd/pKFe5JxCC
bCjtaUzmOa8c+NHzzGgRkSoZxeuY0+7aF3zqdUdxp7J1h1aMdL0LbKsrbNHdXNER
FfEJtSYTu+Dh8jd1aWFu8ltZWJGpXE7DeFMUkvwV3KiCStaSDqR1Toyvh/98Rrp6
uqyVALsVju+JTdtFKO6CgHhtk9LC9/E6AP0QM5mpMnWY7PdpbTLIr3MBcHyxv/wo
NYMIawUmT+1PINBhR3Alf5t57UliqqWVeM690uAyCzEFka6Dn0N7JYNYwOucgLgc
7HxfTLZ6sizxhHzoFxpXj+ocseWvajbRbEdsk3cr/hNxCZJ9okKlCx8MRvam8vOE
7dJ2nW5uHDKteXU2zyUJoZVZk34OgaVJIT8g9DyR2StQ5iVziO2+xVMhzN3ebYw4
gIirHd+bn7d2yftxP7if99P6ZAgxSkUAzdVo75v935Ofp7lOvjOsM2wKkNpQFHlJ
iC9z66fB+UWzLO/KWpOX8gTFVc9b8A58HIw25LveqeeQ1/WWgU+d8iuPPwqUiez9
iJ0UoeR0lHcIr5e9k4skl2BIE/QHCoe14Mzdpxnv84jnRuzSa1PgvOnG6awaXm1p
OfwfkbwdJLYZOYdi2uo3f5gKH5R81ajKt+tV9XdbOOeDUcotT3XQOf61rb5wuRGt
ZnQrRysejGTrhYUCbvsYFE34cetpFCxVjK0a6NNsy12PFAaCNi7/OGPxXMFE0RBZ
VhbJW1DGT/PPqg8AWjpqSILVrKlHGGyhl0I+DcxvI+QnzJ1MJ/li9+Hgf+78X6w6
242r4laAjhybqr8n9N7xeHIBpsI3H08+bT8y9snzOAaD5W1oWSZ/TzBwdNQT05g0
4jXVzfAKUKOtb/D3H6y718dAn8Sml+d3LtJAu00/r/0RbTZady0dStqd0T/QlQXw
3b3AWlNZEWv7lPfQIQ7/+QCqx0UueOS+MKffKcm4ChFp2bB2a/xsGZ9cQzgr81Qg
ayX4soxf/EbcAgGVIBZG2fWDmVRVFmbUNMWX8h2dGhooKpA1fPMb5zerg2MiaTUD
fhZ/4sPwS6n7kRuzcyiPM8ixW3RT4d8Hdifr9rH3+eKkk+robvEIQP/TPnVcbHhl
5Ask+XNltstQi6tDigM1SLdahxu/a05YhJz21FoOCsElHTDsKPfx4NfODepNhIfT
BK7IodvTM8h6VWvKV9mDoSTVWmYJH861M5EHI79hlb7Znw8Zbo+t0K0Ji+xHfYZ4
9M0z+kHHNS7yHGKYqc+tAvgE30tIgoDTAVS9ghr+lcyjRORvxRgMgE2EKEKxD59v
4Vhzk4T23e+OsFaTmOePbL3K3kg+v3eAVkwqz/3KcljuE3tMDv83M43N0ja6kjVb
rIBTttlJomd0m5yDrrfYItyc+vLQTITBJZ68LUDNhhEr756jw9iVvvD/qoFkah7N
dwoLnN3aRahoCl0ImO6jnrZc5CCIra1yizpx9yKhgSzgDIMA5RIc3tyVxvsoHAVs
eKwJiwz1nIEq1F1IJFsQE8NFnVc1A5n3DIC7Wf0gLwE8wBVt1ETDgmTTNrIBdEdE
VGumIt9nN2SuNM0m9mWmnd0COMo4DweqAu1pu6Pi/LqpyK9q4DGIE+UOsdMnGBou
3lmz9GVNJEQ2hqVRFHMK4OQxNx0LWuGNyh4SmPAYKhlv+118wlkKe5xmFUzOsdbg
nz3PQDLm9468ydWwo9tWwA1RKqBscIEZDB4sxnYAVsJ4936MB4YWIDKH3VKLhJ62
FYWwnSwuSH5OcHkFQ6FHzaFJUPgDLpv2Nxxay1uBIm1hPHJvWmIyqX99qsN51Vdq
n6AH2dXiDi0/uNZlgbHv+2A4mZSXBZs93A4D7q9kvAqY4Szjt7IDXgw3dziH0NM4
J1UBNpO1lyuqqOVCPdB5x5pXFeYddlxBE0xJAhlQQLOlS0zGaHnc9nC5gfjOJ4gT
MfL0r2W0Qjzz1vNYDsZPw6OQkDtRD7RaBITs7UAWCkf/Ive188lA9dC0Sva0W9eU
DMxXNzOUu7LS0j7Vz8iB87Tk2zOhl6HY36dKfo8E/CAlcbJIXsQ+k64CZ3s7x+8f
q7Cy62Rbp01WeSCVzFJAg+Ib2AqjZa0Rl2ekoU/DxE9yV9pihBOizOgP16Ony3lf
w07jQRMT/waeQUZElWEswM4ANDDtTueiOY7Su/uuNZ3bQjR8487dyb+JMhVvOlui
TzbV5l2TS3TkNMeogQrFURnIZsCnbcjfYQw4s2OEWTCXwS67bvpis7A1XcinvxTB
F9adxsVwwp2rXQwWTIbYeultfgbeskRV8OZwedGJZ+rr3oltoziFsR6sYerGf7Rt
sJhW26RnJ2lwj5fo91Jkkz1kdwrb4V6TGOwOBrGgBxfrS6UmGeKhdg5G1PURjvgI
fydFe3JpjoEy392QbhcSKGr7vOgNzlt1sOimKjPQ22R9GHNJbJLbkIwKZNaSFThT
KdgcB9jALbhXE7iXSnygK1YNztVmIq4HdZtVFgX4815JR3DXOcO7bAIUqSISoIHz
V2LKoyZkCZi9cgZ3BwVa7Uc8RjqHrE1uije+V7Tl2FjgugnbycDltiJgXKnc84rq
oAxzZbJYXrtv9LGE3I//jAe8/3cmc6ntZpATrhKH8imAvu5sfU+Sup/nFGmkQgD6
XGgCRUgNouxm0PUcqD85tLd+CXSqGebPKF5Eie3JKQG3AptmmkE9PS0AEfHM88A5
mLnBbdDWt8v0aJCumTfoLUSC7l8DBogWQsdDgWkoarymkdNqy2FnHE7tEPgUcQXm
rr1NcwLH42fWkFDOqYwlxCAEKOkH/djiDgd7l6Z451mLFNEPkW5BN/vMSBu3vdCt
FBoIjfBqWlyXrWki6Ws+MA/vO4IqLBsDLTS59vOwYt88/CZhQGTPxFEJWJk7H824
7dMWhNBK/HX+Cm07nKZyHNn3xrwx78wm2jgGycDlzJnn8cnX1mAMVDC7FOfiD5NY
qOj/3bDs7jnIg9hcj2il3bCjOu4UTiUir+O7RyQRly7jXvmzEPD2wnAOg0ZzuwWC
tOrPAoEaqYtbOOX7Az3CFjzJWRxqvJy6rCpzZu/OOQ6N3S130xeA0TmgjGl2b7DZ
lqp8zch6R0riSOOBWcov4TJ9DyicYdu5OtzKFkOCZuCyd6ljgSMvWbJ0igoZ6oC8
pYzlw4rqKG1IhZRsx2DF6TCPPGWQep577VHTjup3X1CTFstrf/YXbZ0L5FbWqJFP
zvZ7ckbHmKroWgSLFpncB29fLSOtZhNyFSIKeKVn3gIKPyRlvG4DOX1+QI0aYSHW
rbiMFeZNGC7SxLsqfSNc6qUT9EkhvQ+tCKSbi4L4fXqYcWSlaX2ROpi1Bp+9Wlqa
RarmWFZSgiY+LhwPwSgEas5Terp6mTiyivVIrG7qZkeXc7WHY2fCib3QNE4ySA77
wTs7viGPByhGRzGbS+z4PWierRsTUmKvgacLban1IvnGkSgxl1yfRl8YwVOV0TP2
mSlmBza36LKmlTeOlFoqifpguuLfF+8r7uSc1OcZ4ECYM5ZOoAsi7Rot4W02lvOa
ESTHMQT1wJLS52rzWl7UIzzjT06C41S/E3lI1GMkwzvKNPX98NDw3JV+iJ8ZfIfa
KJKw8rTCs1zAqT7mZjEFMeU4HruIdyXazG6xbVhgj3Yzl1DHyxMfm3Qp51VtLiZE
2cP//UtQ6ELJnMxuGKTDMOCFMD5SmpZhTgdSr3Vc80XxXHzoCbaIpFGqvUJvDPOs
QhZ2EmbEziH13o5MXd03VfWUStJo5xOblrQh7OUjjqyvdHWq8ARR9EhWBl9c/KMX
fBRUPYR8dYc/0eJN2+rUPuKGgZyZkt5okiWe/7ETdFx9qILibW0yAmm1qaSor3pB
biugpoJzTqE/7y9RO5SZEBPVyyS2zEUvVCN+l+29po/8YlK2UCeu48L1NpvxgMJg
AbQn/7N9Rp+Ojdq8El5/zLcaK8VzFpv+k/Fkf+Ifg0h/GFXm8EfjialPf1gREsw2
uQX2Ff779kD/ZiyoRJxGJF6qmnLqnZOguIXkMIAv3kAM25zojXaTjjdac1ToTW8p
6oJ9n3vNERC/8H67UsJmse7WacFes9To3SbDtwyvqmJFMFsEFa3m8xj6LwAfFNvl
lopr+2zv1hanejWTYzx6toPxWnWTtmNQj1pAAfKTx/4JoyRGpapQvXq1PjGEvXIv
PHsi6001/ViflppgDpaK2nIqaVM/YK4I/+tkY3tar24eBK4zNwaRnA2I8WG0astT
iTEkd/mqhbo6ab11R+xk6CooqSFDFe6DHxgL7vpT/9kGPp/E7xMIVuNXsrdbro6s
JTD8RlErZiH0+ZEUFi25kb+ET7Gcs5Bq7+KBMGPB3afsEUQIjlwJpzsZBCcKKYo7
tCRloZmJrURrDpSSu4+OBhtJHM9+Y4vEokn623bHGnn5sqVVPCg+LWEyzfmm33PS
43iAyRsFZCwX69fF/Qr1wldB1tbr4d9LL15MBDwzzFiFHxagBkMSYZ5LjzTVm6CE
gbRPgiHjzplqGDsYF70t/M9QYG0YHoLe6vgT89b0TJIwT8uXbilN51gM6870ltgB
EMXoIiId5jhSORsq6CFtEg1JAC6f1Y3jD1WPszMBJjq1HvS8yEuEabnwW3BaPNKD
JHwHlS3nksbH7vfKQ7Rf0Z7dO3n+3Fincx7Biao++VyPJUhdpqUZj9grMu5drivK
stK3PA0EPd9FG6wDOXsAOu6k+214yo2vqPd9n9nMFQ4mX2npWtI7thMKnBfIzQj+
xAXO91dTh7+oONU/afdcIARUzyeVGpB79hHVxu01byWjH5oUFn0Sw35DQYmGGIuf
lDeA9IBp7nuqzsR9YKl699ctfDtOYbZHv7qE/trNgEgv5DBgvCXI4NZJag31UT+x
IrBVR3LkmZ2+brhteXPSX5Rty+UzIb+PQaW96QNxCzJYqsKmsJlb5KAwmUexRRem
h/1IN73uE6GxeSiqnjGDmmXt29P+y2vyb3jQT1k7Ll8d9q41PTbbnchDSKpFA4Rx
jjr837qc53V8YY6DsI3HozYA2Xh5A4QUsSF5UqV3ymQc2qyQtD+AnhnpUxwWAQTO
e6fqae5lP/GoUY/HVWl52LTR8oRfhkLjIWWc4nnhBgL817p9G/kfgcFIuIWfO5Vh
zesm7748NY7YR5ccim1qJ4mHWOVVrRBNKw1hEV5ukEwxWhM32gp7joy2br509G1O
mpwgI4bKUg9OPgYvu0LbSmgqY+d3pYWDvYsJwJ+8ZBNObGCuKE45oYu7weFdv7hs
gzBzbdmovm+1wGsJg3nOW9ilmvXCUNcxzgIB/iQ9tH13XFigDFkplxEM5CqPmWT9
gAbnDB0BprObK0OsOQT1wI8syO6ijqeEm680sV8F2oh+Tg2wiilIPifQyLne9Fmz
IbS7PeYzgdWIF8KEX/6/Cd+uOfmBeAwdHWip9ASoK8pdxSU8Rztdh6kwgqL40mXw
QbmnKeEe+popeY/bH6QYlF5HPJ2+seDb7CrwpmvrtL+VbeZnNurJrFmcBpa812VZ
BlT67m/imRx8RYy6O4o2BFOwjazc/7hOdCqoSNyA/h60mxZj5xZNW2/+uHKZ58xl
P/MHia/HOlcxomg5ARjrsxno8B4ixwTkBauyYYs7UTs0JLXXjBxThK7lgqttSWcR
QuSzNxARNf7l6xQMksOuWFehMZeQBBZmtimGKc0emXtSu9h5kocLmctJ7QXevZo/
1N3T6uegKhdDmApRGWL8WPYZNdCz1rwywrWLDPNuIA8B/+EEuwmd6RguwgH38dP+
dwgjmIxkSpqCty7Aws9hD9QNYgD6F0LYwPQOIWRjGeJrtApfNcwpmEjLOCq8sGAQ
TN1dk+qKgFUO+JvBUl5SGHsCOfolZfDSSCb3td/MmjmTl4ryv4S7+Fk9JAOmUOOe
wCz3ceLtulKrO+BROwLxzak2U6r99D6Q/w5Ml9P5Su25tXNfjR3b/wTf6T9C0uQn
0iqFM7LDcS8MmxcU786YMlvprNz/+/O6+fEQJRGeab3xnHcWmohh5X8jijXazbQY
Gnhf28tkITG7AunAk3irt6TiL9uC5KXVVf1VoVOxQWs1fh0Csqd6ou5qR4dJy4ll
Ago+M6bp/1QzR0Cg/lkulP3h4LEbbYKq1pZ6lF5OgbMHRvj/rRNG8b6Pta9aIL5X
gqFGq6x8aV59K27yDzc1UrLqwIuC8F/pc7m5aRMr44J9b1CTcJS/CwwpJFZiHnJ8
fnD2CqCJHC+kRTe/C/Izvu9ilr8qzfBqw4p8HGSfUGL4+Qr4JNuXP1u7dETwJkhD
8ypcxMhSP9bVRKJ+Q2ue6kvtI487m1rTXu6TyMNrY9z4Wv/F6FyZzaCCP9c6D7zy
8/vEXM2D91ltt6cakMZRvZHiGGx9U1wuvUUAtHpSYXwZR44wx9F49nkAuiqqNs8j
pqi9Ktm+Ld/vubB3nIrx8Zbd2EiDWjqdwqhGGs3cW0QVExkoAnkvGh0yTiyhm8J8
nR52mqvBLjf1M+rIyfQE3dWBp3x9ADAwqEFq/Gbsftwx3+DAnvxaqt/OKuYqkC8+
T6LWClT6XoGMQqRBXHNHEdEIWBHKYa4SxnlyUfW/F7K+oP6HM2ywjRhdW7x62+UO
0yggjSTy5B/goa+Ewv683kq5FjDZzg09nWdOET1E3ErkxEtPK2kDMnmkKIqTNpCT
KY21Vy6DMtKQyEjoftthkyY8rXRGMx1AXnTG/jzxwxQeWNYUNiOwA8XUtm3MA0Oq
9hzI15ybEABaEdC//efIJG3lq9/L0jHiDtJ7ueq4rRjfIHsm7jdP3dP+HuvzuTCF
IsIDl62Yn4X/44RpaiXejkcSj91vjy/6eEPb25jjxLXdQT3WP1u1E2kKEUGeXT90
6Fs94j2rGImpT1hMAH/9lppenvztGFwKfWWeqnV/MJGfruKi6HlBuLO9maIMByJ4
3TahRQtgBd8YNox6vSIPvkbYpv3LVqrcoUIwJFnrKhISx3I/qXV/Z+CYYwi+6btk
YY424Ff1dsP/koBx/INXKwl+7KwcylhLfNvaTwXgHrXdG3R8GHUHjBltln5LDmsN
eMoJMgxa0ruWJD28RTud5QgEfqU14QNObwR+BB/YS2L6D9qkY6jl/ngZPSMwchHA
bYaR/nt18lYqFaXM0h+Z4LNtdQtSkNkCBYh4jn8oUG2fXxeTFn5srVaZTiP+GjVR
bxtfvWDVNIECr9AAgOMOwGvxNA7DCHYMGeL3+fmXwX5PzY5NxRG/CmGUHg5qCpDA
bZIxEW5YcrpeJ0gy32pZHyU5ARBLK/OxRIbxu74iIL0+13MbYkFzrNBmS8q82EJQ
vs8hnfAOOTXavvuXpwRj565DoeZgWAD6jjellQ6qDnLHZwbOkcbcXij+bmsDEneh
Os9hT2HPau48d7s+JFwktUUKVdbiFnuzyNPnjsiFw1fZjnKhhpyIdvZ07VPng5QH
GOhsK5rE/WRXRYCKFFJUAwlLcuFGYchPcnWJBpd7SoEboHHqLW4A89KpFQ8KhIAp
TElrOM/8rwaC1HNGxjjwJFU1YkQgSnHB6REA/+3LkHTWPpafaAu7X6VshhUjzXRF
/FNrhAu0BXIfD4rbWhwpIOHe2zllXSDuabHHH/ACAZe5NIZUONBw7R0OPrMa9WHe
tDx89ZLqSlJTQ+LIPl7AI48UlPEwQqvWmSuqaoGUzUBWcMPnmmnG3m6V85kFBH85
aOMCLyKP4DbC4l4RbEoAJhdCh4MMBect7u44Xe9IasrFIknh3RhtxWzMofacFAZL
ua6F0XvjtUi4RuUJ3AvroBtF2VT31ANre1PsyW5a3r/3DN0dhyWlJakZnokKxBGM
ffgwQH54llJanDLLMbJuja2hNuZVZxxINXQpIvtVYoEvO1wmelProKJuVdGpG7Km
lVutWnoj4VX+mZJFZMy2Uj06ekrmX7mWAVWbioZuApal0YmobJZJU9uGneprdvV2
zrQnA2qXiVDKbgh+IRoDMu2axg3FhXOZcy+UY4saPYUtECBilXM/5chbqi0ME80Z
ta/bGlMZc7y6j+eaNZF99oWT56JpkmoymIDlNPlm0RvP83uDkRbyBo2UmOw3nOcX
bYtiT2bmzriLaJhgTe9zGmJjMQIKo7YmSEiZFx58bWIpMpKb1y/hrQrNo07vQU3A
ClZ9CAoT40aAbAUWotaJc+elLzHVYTakcqO01Ix+f2kkhskSTzWww2MzsRpoGnSJ
gGdxFkj479AhysbPhBX4iMmrv4/T27IZ66bllIOyS4MHmun4iNBPuvSsYzmGMPUp
w1F9ffsb/0ASsCgTna3yxVNKPqF4GeQa3tRLGLdfXefaEMaCN0JPuFGngz5ueu2E
QQo4QKBZVg6hkq+u2AdUOMUq7iqn/haXCeO2rMwl+R7RYZ3ey68RjjMk42dzyrSQ
MHheXheEnzWVMpKDy+95rZ7hbiNAH3ew8oSW77vKIBXSxu9MHh0NqnAuW1JRdNAe
9JKca77z6c7T/u22gPsORMrcPC9sgm+MAu3Sez3G1Ucc65NwEiYicASpCdmT1wsA
C9ATglwxt6iJJQBYkx8N5TvYXLJ4OXBMILcCy69WEb7MJ5rSJUoQVLb7/aiJeaeh
ry015TTl7Bdl+ta0Wx+cwciyvPrwT56St278VxQ9n6JJyFcPMKZnrKdA9Pm7tGyH
blNK3ZXH2MZCF3j1/zsVr76dMqRi8OBRnF5I9DiV/C1ivphCKHuIhqqWXby2IYax
Bc6OSzlEE3fDJO/qCKev1MIXSs+00fRdxkPts6KrYLKc285FUu5QXxN1Ex1lOV/m
mwXHCDkcsQqkBnAr2GBQabQP8+3/8ha3SaL9dF6FYB7v7Ym6FgXBlK2oLsrr3CXD
wARWpCs6WDqXlP1CWlj5T6x0dftPO/FOoDuldCig8mz4v9bh4iAbi47UfBQd/G+d
wZl4xE4T7tXXFCucPAxLExerGOSkuf8y7JOO6AE4VSJS2XBAjsYIu88h+RJyGb9C
08hIIXM9fNnBRW2+NDQTi8bo/Cetfjq5mUIXdmr87EZIF8oU4n1yV1jb+ZwPxcng
IEy8D2zwKDxzrE8s+eI9G67mCqyS5xHrOf8YJZMTeCYjMbXGrZLOa8afltQtB4kX
jklXDxXvCSAH2Alt50fmNwc8LJO06OQx5AVtgMSd7rJQvga6tVRapf/WE0eeeram
4hxkNQoa9Eha6k7dko261yV5fshkr5l5sDewTm7Z5MriBvTwJd0vODS2aeZSVmH/
KpVXPTrO9CUtfKyBU4X8vPE45MOjURj4ldxvbReXCr2bzoTBEvBLI4Gc7p4UAdsW
NFImsLrZbatMCBbVdjWeVAdDsggN1DlGwbcdVBwY3ylsuliMfWzzPQ60yS3QW5Un
SfClypV3zlEzXivHRueRRwPVu4vfCxLUBP1vDmKaYieHwwQBwi4HJNRyuAQZ3Pjq
E1zjTPTLm1VWdcg6dzSQ/yMkz4tvCgQ21ALkwWPzWmVgEf4vLc3Bz4UGR371Bvgi
9n/UorDT5YWnF1K0BTYbIeegQQMW1dmh6f4muPLWkSrS49DZPwdws35ZRXozRAFp
wy46kMhfGJEPetvN1aIp6FFsHdf7M5rhy1/5zEgvE++Nqtt27q51Vk0GD2nIGMNN
ujO9tNwM01iEXXLHN2X6UbkN/Icl1fik4Z+60U1fHnrRX3hM197YYijwdPX8r52J
5buMPtCRdMFcAXnIfHlhXiBNNDP9IzE6zwKfstaqVN9MA8M5DkzPObc7sFPchQ6R
XBxOEKD8WW3ScSnmJZ+jpF2FoICvc5djgJOj2HmK8Hm8dHCNmtJ+cTrnL2wWXty7
h8f0wjuvsnNGyVpHNZ3J4nW5PMfpUB18r+VMH2tJnTa0BOMDO4wbzDNT5gloHD+U
Uw05HKynNloF1iwWvhJEkL3fZ1MgqOz1Wc9EvwW0vUSLg/LjZu76akvvLMbFSD41
NhJ+V2nUMuxKmidfoPw6C7tTrxjGl3OYKyGL90dsXmfUJ6HFIx6wDOSI4mVWpGGT
+82v7/fl/Xyr/1PRSXKz1fRzpEvMmykQ/WZSjSLFwG64iRHYFuhgTsXgKTorZQNc
SqffoW3NikbHmddvvkOGsmx1Lnh9gxoowGnpYMJUwC8Q+JDH3Iu30U3QQeP3MoD9
nNFEsnm2u/O6X/jH06O1GkNVfXiTikzKCbpOtdyFYbtJBhJvv/hf0QmmFkZTYYay
/B7pWObhY+PVGDd2PjSl/cxzNSN3ZD+zHoppjHzkayL8fCDwwdPdsCCNXy9ZXIV8
roRh6jWQVOotv7GqNrlbmRxGCC4QxJyLCIIHZvxtRFmSZrsxR7Pzs1MpQVH1LovC
GVU8k8KR1GSvE19nQwBFGEjv692vCcjmbEgJzay6bddvMpwBuaST0VKdLUuue2CX
Mp/pu7lYa3C7uHI4Hg8Qr/CmVW4MoyEK7e5qF2xQZGRg04FxdPt9xfG7bkBdUKzq
nijrosoX/8k7wCf8LUJubAQcBXMKgBhAyTV7F9aEyvU+SrwS9x4AkgR3KKtJn0iW
Z0YAiU/c82Y8Wsu+aDEaJ6smA9nRYOw6AQK68YhkrPcxiXGx16kwq+m3p914/c1+
6NhwN6pnwGFYVnnYeRhGHoN9WGTWAycfIgl/uyBX37GmVsZBSD+BIzrSTPZgjL2m
z4MTKv3V0t6VNyepM/oqi4IBJvF2zm1wfDW6vy9M55yxV8fhQFF6bIfPmnKszMq3
l7Zyrw1Ad6G+iCtpzEvyKWq8rJF/tySt25yJawifpmlRh5fXz2i4+2gctzLMtxmK
xX8EBwSjiyrxbLdJpjU/JlAMoAa9ZTGmXl37tRfUmFZQ3VjHjCKfDazEPvNB+kIY
4ya719RP6pQYfToVJuKvexdtrub6mP7QDTCIPnsFNACp3R0C+4pZhDvD2tHYoBV7
05akOKe7lUDkhyyQnejBWnkk/gg3V5zf0AeC2TVNTt0UuI6stSfnYqhzHHkH2dTc
dTU/QuV3waLHgfsOPE+LQqwZ5kXdvjjtNKeZXTuUOkXAdZbY7JUNIUd/J0jS0L6+
w48F5OmFHK+z0BVlWIx8n/sY064BSb9D7a9xSoEw+sOSaWI197yIt9PuEmV/rjIY
UXuoOW9GXYfOYZOI6JhS1Tr4xBtUMos76lyEyu4hQRewvT7Ud6xFm7vmvsm9DmCJ
o+eNZbkmEl7TLgpt3lLVOhDXOLRGpLPfyPWOCzDIUUJUWH2jzHqWJaRMq+rpvGB/
wFNPi67W+AUr0eDUosScXbuKLrFtyAyKRRRKqRzjuSvG38sdv0ZeaPhBsoKoZMW/
LbskTUmW9yG3W4GnmLYMoyd/5SiNUkTXSqlAsBnB6equEojcOteyPmes2kk5hWm2
rMliUdYZ6UXtqyn9UwhIlycMc485TVfTjaln7DCPz3333Pp2AOGFgWX9qzZrsHX7
dDHg085yRKcOKd3HT+Eheu3xD8gDWeoadzI/FpHxU62GMLx2YBI3+chCCZICFJWj
A813a3hbleRpY1/4OASk7cTAukLwPjH28N4XFMpEZYMZYi+uCgcZpaHGP0agvEDB
5Hd1uioCuZBzaW/lEVoEexYV5QKsfanOckT5JwXr7mI/DBsBt+R79hBpzvMl4wfG
oOtQn48llMNJbyBVvpGcPAbqaMitlj9KK+9fUG7f5W08gQZWIUTwu1qSmBS7oWd7
3xDnIL1wVqgemJ5UIRpgpj5veS6IXmDgab9ztS54NFK8U0Eay5y58JKW6BLAK1bh
VZiIcRu4ztclRI3cdLvT4YRIWWKs/QL5bNGyeN9MZYEknOoD9aw6r8uo3QZ89EA+
4URefjgcE96RJkesvdgUIsx0E8mgWqXQR7EgWUSTZd34kLWpYGWgJ1Vt04jFxVVL
WeMTVYgb8dILqtEDBhE48ZPOe2aO5P6XINNYPpYPMq92CW0MslPspkzhGrD6SR/2
f88UisK89kfFMXy/Pfy8JhGYY9CxgOSr6pnW9vsrsdZUHtDm74HjaXYPhWEujuNG
JputZLJm7aDu4X6L2NZVCPh4o5wsX5p/pSGp5HgBan6/o/22wtrdNbOR6Xxln0W0
AaOxD51ZLhgN1LLgJXk/AJBs/Xg9QphJ/0rrwfprfb6tbiMkvw+ew+GXllaDa+a/
SsPSi536ASH4baC2FszSA5jifG4a6M0HutXsVqbIMuoIz6W//I3gniBLGjwoAjbk
5Furhy1Rq2MUtqczlBAJDpMFpKWAIW6qZIX7qeH0TAjuKUrrL8DagDh1hLafpGPa
S6Gb/757tRuSXGcox7YWwIJeMD3SgeTyovBbYyI1ZJJc6/FPWydLnN6sBFZQUMoJ
qbNx9zgPQQ2tfzF3L0HAQGXashFtohEf6tq/XQL+Bc7xx+JgU9cOQSLVpYH/AafR
mIIRCkQZrUDtPMN8f+ST4SnbnMotKp0WrXMCyLbsJwMemy9l/95+JW6qz31ng+A0
HNzw1QfHvSvzL6rzuyhyoXDf0WQpB6A+v6qJMhrNR1Vg5rXbV84sEozEFNh1DIpY
0C5WChblGrKjk84hkS8PJWODDaI7hhrZ4Qcv4helAvgOz3cGPfYagiSehhLJ8EpA
x+V8QxoaRL4jyKmH0Tey2nVPivNpcfRsCQsRhX08jNTwQ6R1IuR4D51+1XXi7ape
YrzuZRRbu9w6mCHknhwJ6QivD+doKKeT4HusglMqeN2iBQPTunQG9nyjBlKoMha/
aJzAdc370XhI73ytWa1+uppwFURTA0FZOdYc8JN0IGKQFW8WN5wD104GXkXH8Bio
NTmdQiFwQVu4vOB9B9CoazjoCimcazCoH34P4NY4nkod74RZS/QtSDyCcQUdWRRi
QZLIuV7QDa3neoE3+WRF/KkeBqVg6+/CqO7mwFWISqJKd9Q99kGJZ8qidv9U5kTS
Wg5paLtmMbO8KWjsLoYFFp0gxM34hmfucsaI6c+ymJ8Pd5XNh1uIpbcVBaSVngHi
e7BXFe9LrT5jJDxUWEl3j9oEtDVuz8j8H0lrdLOPYWNG/PdbWxlk4uB4XlQHiFno
7iHF00gEh9vcELRg4ULSoVBQI5/YKOjt9TbIYFOMInCL00xU/DQbxiw+0KT/XGSv
WZ5xwAcVGbgqWfqMlcea5HDhlpVLcXdccmejdMaSFR4w23rD5/uwvNxwZNDDrcC0
Q8CpBx/H/u7PboAskqacclraAJXNgU7Fr4OSviqWNwaiaSILj64rrqjw2BrCYcD0
/xEAAPKyT7j9/kAut1PwGnwtCuu6QxPiEZg4NWAUr0+L+aU0j/e0fCgpcTKlwjYN
tJx1E6kC3/ZQYOqXEyvoeQ6C/8UIGveAyNQUfbooLaSzCr3lfK1JlaNK8410G2+T
caAV8wIgc06ipBeaEDoKKD0+Jhl+ARrkhWV2K30jH1mn++YA1E3ePs48MZceCLW0
jbFoK/Z7IauymYxYOezjiVRQSbWdnBMz7Ka5jHreMgsnReVJ+nGK+j9E3NGjtQIo
kU7DdJDjg4Kwx2aS/caC9IaVfOOorAeURl+u8mpfMqZVNRuwAnB5sAgo2QrWXjio
RxcqEdcjZegP2tV5vynphxUuFrviJwuBm9NzbJoKySLqCUuw3PXMnyW9/+Bu/ZAY
LusshSlM0r8Q02nt6IlOeUbeMHZmaVa3FUwmof5n9n8erFxEWDrp2JCGDGaJRwoi
PtKfzWz6AfHScreSY1FcTvkS/LZsg+SMnifAO6rt5uteCl8uoX+DQY7rjTacx1K/
GNOG61xyu0IzHwQid1ntx3Kei2J/lUJS98FDCi1/ILxwGRGvFNwHjwFbJTFejOPk
CBZPCuIyOHHLbfBs9/hC9tqp3Ub1YvgWgmjX7ky7iMyLr05b0kM+IGdLj+lFPjN+
9EktT7jarSqp2eZtFxkDuvuymeAXg8AsYi7coCzqPxSmELEy0Yg7aIUEdpOBl7yN
Tg7bK5qRMw/awBU3MwNtBAXQAKpJVwuj/wsHYEp0elFN4ZzW7l9EQDGT4zLsLo8i
0YyAQpvMCRcRs9Fmh8aGJFhAhWOc+mmvkn2eO1EouHb5HuWvW8BT6Gcyq0Ru//SD
eKVCEVtio7b/8WjF5f48kKVNxwQtQ+YEOFGvtjbG4W7ydUrTJ28MQVlviKpq6eKH
Ep31lughDexPM8+MjDB/e37zhbshtT5sJTdOMpmHS4oht4EbcvKpalBnFg7btEoc
Gczu72vF/Q1OD5a/49GzMA/2zvoYuSDwuzxKak887OZMvBiUbmPtzvZ/ZFwGXYPw
5jFQ1NdbscKs4OLc4UhQ6LFyhUXNZ+KCLrEin7XJ/lMQSzDHlOcISdA+CglhcZDt
hgkCdvGLffiovdQ8Dtyj1eyYHB7ws2gCAGtAcTBWXLJcSs2p5uvqsIaustyuIdvh
dawPCSwRdwtUMluX5Hu/M2M+xP/7HgLPqf9yZOHa6R/eJtNMxNrTnPwNcxuYLwqi
2iYilcQo+XmZz3y7QjOtdAjaNrImsTtZQnmI5Ll54i4I+HSPwVLbD0CNLFW7hTDk
mHkAGjOB9BhboMwXoJ8P5NRITpYk2oss6X+ech3oZKRrTNE80HMSQp/ve1DjFhaY
I1toqxk/PkCkRPlVdMU922DqR0y/LkPC9GqwBMueel297fUIFCDrbo/aEyVaAu6H
9S0F2dfMm5fDcxSJR2Xw5P2xFSv9qmyjHc7IPqFYCXRNiTK37X94qWBGARCIA0yB
xWJq3H1Ohe9Sz5f2AIZLqhdlX9cLnTE/X/CX8C6wxYrtm9rH5I5obK4jVNrcBi6f
/r0AZMwZgofRHOiygxZPr/cyIjqrkFsSn3L1vi947MIrPf95YRw7/4x46v2l/YKN
pLH9jUDAres1rNOUa5xLmOBoPvAWtznUc9zXfawpVA8KvngXewVIWEBn/6HeoCvP
oaVVPvEI9Wsc/UO6Gog8vbcAly3/srYimJxw1907vqMpnI6XPHpVKVcQSei/NuJD
/luTQnlFZeasjh21W6XD61mXi7sIfHltsUw5CMT2sBCdo09l1G0PPRqxGzeteAmE
gV8TwDuYcUjiueJx6GXKnClOoh9GIYm5I/iVovAmPvltRPnIWfX9IrSwjUaU9Zry
msxVONbEGJIms2H48ynzWTXJfD+AmCfE+dvJk09L0gKWNvfFc8ytVJYe04D3v7BX
L63VS0NbI7ivKRlFDGYRyO6skwWPF7Extf0WgJ2HolB34sB4kKhTPAIwORl8zIj9
0bvLjbCkAJaCYQgXGk4d5k72k9iFa63FD/sHJ7ivShRUr6sc/1h5NDR9693sUaf1
w/1ZK0vJC8cIyYDX0QB7dv0kxzTWRw0v71oB2ggoV7rMeax2Aojsoytw1AHOG5+G
Ndet51DCU9os2vpLgPzzpEcBT5iwYNTgYKdPtMU7DupxLlOcOHQ39gs3GKMT9TxI
T7OawS6Ggcft4KZxegABiiRegy0N1+1ilIXf2WKwFIWrqgfeqxcpboW7O0u8DA9g
fQyL9W0zAVrinq8C8pL1SdDxWGdF+ojCVeyrwR9Eo7UVoCOS3jyIec2nYVHOaOKe
0vnDX3egPfsndTSfr1KRcnnYvSrD03LQt0srlz+M8PUZ0Egcf+G0hXbzkzFuGvx5
w5fX27+Nu8PLCF/uOzBaGyZlxzLp2EQQrc5bdjkxf7UwmgGKJRXaoTRHTayD1T0a
J/CO41yxYKVybUMRSAQSFEzmNoNdL2vnZ+srYMs0gggBjmG5qR6r7tFkCucWxZs7
S+k4TxJlf+b6u34O3s87BExVIjbMJv3UWkWRcpIXMbPPylfHvRMY+MQZJIXLs5tP
iL82rbTHU5z2g5UBsUtzl654y75VcDJiE7muW//f6+zvkTJp9Nlcn07zzhljSEcd
0FdfsV7DK5N6iLNK4s66agzhpdEI3SMpg3o3G1suU7ftHgchqC73IWQLIuFPnKi9
wb15rUTmQQPpwm1dwe7cDHmZVs9DiDY9RnuCPL4evaFzacTbyv3BQJBALn9gGaAY
9foQhOaxa/dUV0m0coMxR9OzSAGx5N9WH8VTt/EaskmNNy/+0jhOM7rjwb0Dc8Gp
M1ciZS4dnhAdMjemH1yMDBBzuQY6vS4Zb0fMfU6ldySCiEqN60G9vluyuelDZ9zg
sTjXt21Oeca+SrVaWVgiYliKTv8EpCr+wuL0XZij0bk0TSS/5VTwVthmGGA48BAQ
Vlt0NvirXm5K21xUE3vHoTpXRdgHNJJBSaUYqUZBr01Pa3z0a/8JVBNOq2dDPfzJ
/wpln5TWqVMiJGMsRXgzwujYM+CIv/o9wVHq4FfYZXQhK76UwguhLFnj1Hmauih9
QodXFV8FcuS4TGV4cpICNicJYnFiJEPrAr6vqlaCmFKz73LIqnm4J9wKAmPMc9kL
k3vcjzBOFIfMIh7C/4FKGTCUwaYZesGzvcr54iqZVw/MM7D7Shk5auNrkpyU92aB
lsNEDn0UU6oi5nNkzMkn+hzI2p9qh+l6frTM+q0XukF8PAenvCHN33v2PoJgYAr5
nULOCNbThjK0yHWoJ6byURGXAUSos415oC0pWiuIAuHG5j1mWd/K5SWkR0FiyiT+
yJqIx5/UrcmLLksicpkKBuca2hH6OmAf8y6aLbZyTZ3kMUOgS/ja0Z6/tLmf+Wv7
lzwSzbMXVTD9P696fss5dsPB5mmUAHUoxptn6PLy4u8GTNtUu/MgggCPu88b0dCh
fA3k0vlsojhfQZbM+98WIGZoXT9h8lcIvJWu/e1bG5VXHbV0x1f/5hQ1jm78VzqO
Wz1gj34wF6YKJ/dU5eW4EodYdIVNEo7oo/qFtvXUN/cWa8DurhQL1VlnCnyBPa4w
n2wmlRwcQDGSsZS1t0JmbfvJq6yrJYjKAjOzvLOXB5rRhnzCR9asX4NPWs14pIM9
bSaSzXfvHcAa963NZnHQtZWHRNBSJDoJm0WF2BHTfS2w+ID5UPfl1ixoS04kxYq2
5I2o7n4dTanOuZv/szrdQ7uCf/D+JVH1eC2wzAWrdSxX63VejUTkps8jsX67MWbb
0q0ji9M0qz6dYKwm4iNMa6YGxlbfkciBNDwSWZHtRwaylA3uqI1J2n8s7bSy+fgE
p6jxhOVFlAk36Cyd3X6ceH4YDp5qIehUdHXNNjy4MBONW7S+LBV3f10/x8i+owpt
dR/VrP76m2QcduLGrMR/6UXkDa6PY95+99/5dwTZ6ibLBZqYNdQWz00ZcBK7yiIs
XCT8VkiLqd+D379hNSvaq18PXveNtEcq+bK8v29/qlFdlalICtkeI/NM+iV2qmuy
tGTYMN4E5IPNbVtKVzr5md5H7jDCBbzItgwqkL7MyEzulYveNY38moTL8VIXc/gp
Eym8pxDsDsAAiBhB2q7r+aC5KSZolTLYpTvNiMZfrAcllexn/j2kGv6GzfiyfWKU
H3pftGpO4kxZx9PYZdEw1GbGWLlevdsAuFiRcEnX1WKJIWNZ/+qcx0xoyfuTwolI
NY72XFMJJL22Avdsn3nm5ihiEbugHhXrS7TSqtoAZCX7essRqaxneZB7xgV3f12A
R9bzV/q9qFE8d6EjrHC6IZSmwbWQ11DPgCltaVXOpkom37JD5DB4O9Yl7ua8pedQ
UKR9IgcTfC2dtqrGnP30iJH9o+52Iyu/mTpb09FjG42Cv77JRZLJ1QHdNlyx08fv
ImJVLB+hReKLUQtgA0ZeXE2AC67y9KTwwgUZsbrGY+nKQv1/fHKzohGG9pFZVQHc
OELyF1KGA8AJGhAS6U3ZUqfFO8rtqCGVmMmSQDoRyjpcmE93zMX03DhBteGqWdfF
wjoN/4w2R6ZgL0k9fIdreOcjA/3nDo6ABsFexS3ahRcrtuM+AdYUNn7FGDiQEp8u
MB6a0Lqc9r+DhCqyzr+abpcQVeHuY1roaoNQe4ga7zkCS7rtrGbSDsMt71UXP6XG
Xgn/heLNKif9uoTnRT6S7xZbDZzsh6xfgds3twNoj2yNwL6DHP/evyB+crT2tgab
jt8nUGJScUP0FfWAfCWza6npMCZcEUYjOAkdepFjSOwz0dN2fjIBlcRHzD5/zuP5
PhFLgLmawsK6G4ZTePMRHnC4BYWJt1vOGSFKQ/5mYBQVqmCgeXqmtw+Zu6IsMlux
5gqMcuEELAkLxMIhCZJ7QdXdIK2OVTdaGy6ZEO6QnjwK8RvCVZzt53RRTETEuuuC
GDY8BADp5OLbvoh1Spo6uBWE8jJZO4sY5gDcGthcIuOjwWeZy2WHSIoWB1loQDOq
wi8aJ4oTKsggW05Rhz1MQVj8g43bG9ZvQBFHvjKICSgrkCTOYoTFMW5VHZ8nAfxP
zz4ErRvB6Ub7NWwH9tl/sn/9x5yFOT7JKFchD68jE4ITFgf7w4ybgs/d/ZCIDxVt
Fmh8lGU7F7ldBFgaK2VghPM6vANpeddWFwUHmhUSNFq1/qeaCBGJlrepoPcGzqpC
IDhFD33qY1HTEdjKQ4zASkxNSYOvwMANVIN8SsSljjDKd7Z5NIvu/Ey511M5wmfa
8X0YNjKiHxJwO7fsy2CvD3Rpv8o8wWJg7hx70nEdfyYeqA2LCWsOaknyGajSvn17
BlhDLeh1TNTwHoWVil1356XGP/WasEXpT2aRMQSNhGrvvG/mu6ezwdWSQqKT2act
Y/4yItG/B9XOpq0g9Djv4Vk2f5o5fyWOHN6wWub9ac+/L0PFE8ua+m9wtOLRPaBo
vIdCxURO4GnMtFC7gM+GicWoSTt/tlB5BtdEGXCfUANA+fmezGzet8CcArFduYx7
TEOjmYLlrvHvLePOXd/ngMEa2n9xtrRBPgtVFl96EKY5AxohWnOCvEsKzgjGvk9Z
hcjJ/G4oIOS2R7XmiVbv5qn2SlZPRIbEGLIgim5hVaIBfOqjwlJ2ENtmCbJj3bdP
cP11BGeck3f3EqQBrfIF5MVTRQjwvS8L58l8bakVY6XT30pvfjDq13TlVoj4DGhf
5NlXbdOCNtbmdg55CcR5uGmnaxzN8N54iBqf2ZhPKd6D/u0WcAyMzbRuIc7dlHf9
MnwvUz+VF6IlS+vk3GX7jOeFm3QCc8sru374dZ2mkzgIM8F/IrXIUj/3HBE5bEws
vLWn3TojKQJlX/S7909/s8jCS/UtAC5X8B5Gp9rhkH9ms+ggI/3d0dgwEQNnQYZi
ZrSlZe+AbNNXSV5RDIZGXXWTiOnBEXevfvNJnXN7UgJQoTgqcPPnihiLDxK5HTkv
+ZdBwywMWRFUbXiSr7ZjyBMqWbDvk8JbVY38P5UMpoJ4K0s6KrwubjGr2EyGesYN
YF0nu8rvoHP9WQrhQmjSvBVqMJhDQQdui4z9ezBWc6jABsYJ9cjwSugtNBuEhEpt
PiiSfTqF4tgRqm/y7ZprsPB5YNITrgeTtLtey3LuiLV38Y54XcpNUTjEYVTllw2P
HoUBpMH5YM0HRLz3aZIU7ULkoixqsli8SIl77+TVqKwXfAQhYwk+oaL8miXwJX86
z2ma3jKSo53DPWOCSiAotTOz029vtJImthHs+XhsRSwL7T34nMQ/FQ9606BREEFv
CyNGLCB41ZWVbS79+yf0bgvHcFOJFpsJXOX1xlODQgqzxEQcw1iFhdPHehj/wOR4
GlSa5mkOQVg/cMJSCqUHrGj5MOoHSMG9XBjiucuhVsMnWSV6qus5mVXoTDpyvlLy
ruD3N5RHcUvRQW5qlhPhk+zBwm5bC4dbBZ/XPfHxKGlN6Ox3wR/Nk/9ay9mk9eeu
lIFLeLdLzC74SXFfzpb0YrTE/vXceWVgrtFcc+W02DtobCzm9ymiM47GubPUbgPb
QOcYfrLj+aLaqbTS0zWPJpwsfeO1TTfI+g1ZGLstmDaSgBhgUZhYKgIL2i6nJ3CI
TNORcMZVFUs8t36M+CVvuGWf/B56mg98Hrt5EnaTCmGysc+zwvJ9X5QQruHmxxFL
Byn3WLILZv9XLodQdkJB0vEDfisBOv2r77XfAewLUTnmBdZ62wrPRPjWBJtYZm9n
PnR4DAAbR/6kVIAyrJLYvG6O84akTTpnfMaj09djOUNFhoN3YshNAbZXzqETURfQ
TFhjkJrPQdOmVBgfCaQH8qSTiilTfIz9awG/fBKgRPAIwRHvzntHXLvRXg+H45Ap
ivfznMM7ADfFruU5HQOoKjMW9tRIvER1Gz757fT0XN2AhGPegxu1Q4c7CJGN3LN9
2KeFKOCog7BwjdHPHph7u53kkequyaTSKP5MNL52ys/gDQVb7CE7ksm0MjNo6df/
KHuplpUCihuAvAxOnuYSm77qzuaCbBPxO8ADPS0yuL0vhYytZcmN2bbEzN1WFvm5
3W2TEVTYDZErCgBRD8WX0fOPNLlTSIYh7N0a+GUF2DT5u1XWlX7jB82at5guvJR9
j4nv5niau7xjflK+DfocbBJoFGMHQP+H/YUoDE866jIWVp1DF9uUISkbCl9XFO45
eRD18/TMehe8WjrlvAoaGYW8BAh0948Q0gsOTQfVTYPKyUAQB8rcBc4xQKpotVSw
4TQgQQEncDmfy7BeYtgo04OMR6R141387NdFOWAl4yhdNaOcNNTbaHHva81uCGaO
MdIK4S7/0XVErXYmwyaYO1ubHbbkNI6HtqgFDjRdYv+G+cj/8Piq9PGLxKmIJYEY
S8MxqRc0elNDg7NaEHvXt7HlRg9suFJeQAccol1oo/H1gfpaR2oy5bi4nUSh894C
G/diXA7KsXNdZBxm+EgpSJ0PAYa0qarSMkvTrA3sluWrDb7qiTcNlpA2L8swjq6q
ua9Dx8YAlsgaQXAX6HfPN9HkLi5csGLHXXzF/rd1OzhFbrK/3g2OVc3FDa/4wxMS
Zh/50UcwVOc5ZI+kOKB7WOe0w1BMJJfpLE4OXuswc3cbZhb7WsEwTY7fiqe2RKp8
tVzPiFAoxRaVw0LyHFpU7DrteQu2afn6Z/kXHWSUqDXOb95DPf2qrdEvTaVQGhqk
beJaCrYTBSh/RY/0W4wvM1HeW9ZnGhWgxqzNI0CoecUWP+H3nK9fVFThA+ZU+3eC
vb9C24LWKNWNS9soS7Je/ngdbPzE3mpVyAazASpBs3Uulx4AYasl4LAn1rPcTWb8
E6WmvqhQL+MSnGjk5eXdKZBsVTj8Gt3axWqr9cCcQ2M/6+CkieN8cAt/1CjTLbuX
VF10FFtTIVjD1fxx5lE3tpTO5Yj/58rUfXOP2TIhskMpTDMe+Kkm9kNAtipT5Br1
pVsb2TyRdOQ5jVBjmKUExxLGXJuLTTxmEzQdXFa6vcWfHuu6njBvSAh8s+sM+Q45
/XT73ME6S7xi90LUgkD+5Q15/2QJpW+l11S8XdYrNoxGgo+YRj2sjMoAB86hRw5t
+EXLubFG/5tX2P2+l/dS+sC6/mbOtLD5lWuE/mPZLGlSHdR/iBnGH1xR6aTOXSv3
/mbeJ6mO6VVINpjk9nlIoEvnO/mhGsu3Yg9X9HL5dcdhRbs2XBq/SAaT4KT8uUUG
ryjGlCYxHZ18hkI5wztamx7qClmnopRR5LpgLEuApRQZ/otuU1k7IDDtrT9vuXgM
ttgbaEMMsT8xnehB1UAenPU+feHJE3or2i4T8xbp6Ed1r8SKErbryVJe8I8cC0e2
m4SI3Z3CEdaG+1/Rkym2gTTkN75egDUB/wc6TKWZrC4umHFRz9/R35QwnxJ7vXg6
f709UqkZ8KShZrxBA7feEySLvfZ0hBqBBqm9LDweJyX0XGPpPfmFEqlZ3YY5aQzm
VpOmIuxMEmzm+XSWK1Eq5+KUkkbPu3y93HwDCXYMqzUxdwrgFz+j1i3JBw6RJobP
sj0Ccdxs6ljGctl+qZik9JGqhK4YBRRdRUX9HSpgIwC3UpYv0rowbe7ATF8TD4dl
qDTCr/iOa4fUYMZ3zJv7kNjQ8Sa12vV0h/JFgFRDPFahMsWuN/tccekpFNSDLpkA
0B/O9Xcjh5d1EXrE9dafSZ3uGJwt7iXMoWMIjAhuPna9o6b4WtLm+idLqBfFpnxK
QcbLdrh7mMQE8bC8zN7B99IFUPPHPXrVUlJEt2YWgzYgXhZ4tPu3cvA4roVae779
vxFIwwZsOu6zEsc/JKtb3GaleAxNI1oSK5jRlZrk2jIA7G/lPX1UITdb4s3NIvBO
KQJ8DpvEQ0rGi0oTY2Q4K1iQR8YOYBzVmxU4dDFfi0BYr0ltEsJRV2ufUW7vS9fL
myU2IbYQVD/wv5FDYDwMrMPwO6njiwQu1My/GodGH5PaQ3Zh8JCHwSs60ffE68hd
xag2V8jcaee5kmkqxRJkD36tXoNypjlW1hw5n2Cs4NJHdTASibM0DZv2TWgAYcFY
selkWQRuO7iQ+CI0c/bNQpfqymbqS522jvyV+OXMXSVrFsTIl0mYFhYcBqwGuxZP
898LRAijco/oXQxOFwN2KktSGwwLYRnPTMOjS2ov/OvDp4YghvnGgaUv+6L3vDEI
BoqZJA9/lvJjqNhiF8U6n2VHdROzWY9IK/F2PVJDQiNsp1M0V8S9g6ZoMvIrqK8Q
plu90tme5WGeKiJGiQL1TqgeqH0a0Dk6470T3+h2CuJUyXeRtsLabUsfUZ9bUIpZ
zWbWUEP0DBnYlMPLRPbK8Blqkk/NXZyiL0ZEThhSAq+b1XJDvU4MMzTXti4xPTbJ
BKWsxXODBE2st4RoOmy9IwQwk48WvHy+keYYw8oQ2hl/ONTicDEYPPGSFucpEOa3
+sDx2qses79LcGf2YNVGqhplzc0u1m7DQq5+NNBpi4Ru2XuBhzsEapW87SSoLt/F
g6pBdGAqjokfqTztAv38x8xmunL2/yWegoT/k0JJPtGqle3LNkO361uY/O56Q138
joNN4R9MFKgS8d2mFlKWCrka+T5hp03PnN/vnUrwtjpEdYnx8+b++K7v3s+SfCtX
Jx1AG5HHP2ADY9iDfs/hKsTOjAouON3xkxexwdqI6U0OfqZhHtrF7C1a1D0JPzRu
l9N0GctvB+WWOAU7jxVnQ6Cfedm1DHGJB9/7kAVHYypJdB6Wfs8u/4unrot1qdbj
aPEde9MJAeZWxpoTrw9uIygg4/kOgLDFoPjrkCikK0a6QsFZ1ozAkiFZUiDEMHU/
eTt7Y4kcpDDe6AxTh2rEmyo7Agf5a1oOIgnhfNvbslSggdF/FKwP9mg+G8Gi6fJl
+r+pDKu55TR9UntEORHBDGaF1NU9xiTIOnVtiBpv9emfQf8WD691IWArEm9S9YbZ
MC0M2gR83QeveINVnnmwtpur3vXmdzP2KHG1AItLlDb8ZSezEDOpnvc/02wNIklu
mjzGeO/MugpTywWGvNtH2O2u9asn3OJClloq1GVJAbVqaqoRm56QmiPGSfxxX/GX
MIZ5NRfuFNQvAxkx4YE8b5RiUMkvvoN3288G4cmLHkxv/5PR79RK70XMNetYf6Y9
1EwZJxoAlv/rtxOta6iRCzHx2t/I/QUb0CL2fEWvtoyM9uZag33kYCe96C3uDwyt
EN52aODFq0U51EvJ9aLHdVhwwq9uWs/ALKV1R/RGMTbcKrvSI2pxdgG0Q3qs6prW
REgYlaAS1NJ4qCxXTFx9YvorZEXUAmZ+Pi99V6RXhGrlzLM5zZonshWghLG09tK6
1JhNDERlJgRHMISBWCOJlDSTn26jrGbdxroAdyr4ahYpbnxJRD76R9OPW0X4W36G
pbva4nLbXZWgRn7zSoSRgc/9iH3+y5RIfkKL5YPQsDodY8o7tFm4Z+oxni5PBAlm
6AiQ4rYsNAPS1n9T+BqbtRX4oBZ9XZimdYGC7SfS1k8I6nH36agzSsjAkipwkQGb
pxLx2F6jfKRf0NKVeBt5eycxtu/cCUVxMUI4eatnJyWeKx9cCWjTWDKgf0/1ytEc
YtN44fkuxFDCo2hjDVpQUcNgxKIHeTtas7WIBl/CLE6okMHNYSWTrqJvbaEigE45
phm6Xav2lmlcO+lPmyv98MMz8iOGWjapP+3mWOyHQ26BDaZVo0bx/dCmDLtEExSK
FYbde38KF+rtuitqZcLi9B83VIVbl7H6F9Pp/5ylXhkZzU4XBOjk+W243UNrXb+Z
lLgYls4i1spGabzRqn0f0NrHnFbsrHpaCU+7hgSssJwS4PJDAYeCv6f3d0ybhLCW
sZeXAzCIZuyIlqXB/rgz3VSb/SgDRITu0xHDoYFqfl5qG5rt4W0VyUFhOyqte55d
pHPvIQtBD7msCipjGdcijgS/KCFS3ErTIzlEOA/HQFR3zQQTzoilQYU2qraAs/id
zzi4L/9JPtfcwl+IqVRzmjd4l0X1BX+fH+Dk12N+reHntJXRmpBQWWNLkdVKvIDC
mUM0QRLMFp17ZOaa/PJVXoRw0vsHKfA7ecW7iNN3njHQaSVPWTO1gTamkeHhEfer
wZjPg0kdeBBZW6GvTZ50F8dEfaE/+1ndbMzPYY8CHjhuoOce/LrlaqjXeSOYvrIF
hZ/+AbVtJ/FUAZ6votuxAmMnh2BdYtw6qgtELOXrotqGRJWJaVr97FmaTjg2h73p
X+orksbyWnN4UTZkuTrOkcFtv/Jms6YNYHPoVtP4WViIk1ePx4YZfXVb8ny4R+x3
JZyV+Pn2a0fXI5taPyhsUeKIuWDW2oiranlhK5z4+IjCBBfFbmjlapOQmaB+O9oj
rK/V9kKmPlFJMb9flzcFVjW6NZ6rhe80e3XssvIwxQCLOP0zbEAIJitTMvbX4yYH
WxK/xq6YxXEcg2jKrYOqYbB/RAvlPiMEtS0bFMTevrMPSvs9YR23JvGN1mwVQdxt
iy10b8+CU3pgyR4FKnii1x9+EISLm3wGtBNlrWdyxJ+ImwIWJCF8JwMrRNgy4JQO
VnO53tKcgs45kf/HKWgFOXY3w25IXMB5KSkzQo3kOLlo7N2ujUtYyTvaM6sLl8eL
7RKF7dOMGQ0F0T/CKMQKtJ0GEwuV8j41B+gcPGMCqIVb1s+aCNRmainXLF62ieQ6
rGUKTaYZjhEpdfq8JVqrx4hTVW2ozqgM8zf6E02v2onu9yX3WPI4z+wpFiYj9JVf
oF+MNklHk0vRvKA3ldJCIPmztbSwEjuYhURFx82EtUxvOShjlH69U3vHZuE++2i+
IRy1w+XmZ8/Hn+7Ja59NTlHt5MuW6pNU62UFdrWcuDENzfz5bPbaDSqe3ESIiAFI
rieJWKdj2/SBKXooR04rCRACor3UxPJ3YsmKbrgSy+YSYhzn62GcEkRwPQnDOh3P
9MOf7y5/ngkdmhAXCHZ5yAAsHpZMfheZj/TLGSALUYRyaLgF4b9yCIBWmuUukVWh
S8wlvRjj2zldNsYybPNYTkmL5QaOftkborpAe7grX2BGbR5/dSIgQ7a38T72WBYX
HLVUWZXi+PMbZVq56bfV8cus9gItmKZQh+vdgk6AUa2tB7Cfay9rQ6lNnIxLTLlc
hZ+SzHA1BcRy5NtIXYcbRcN/lPK1+DeXnhcXEUzfIiG4RoEPN+7IkOiDV+iuDs8c
7xRFO186a/DF4w7rm/285YhD43Z2jNsn5d7f5Otfj6eNf1WWKq7wOnyn1dvuCYyz
tCsoz/HkTPA/RfESb5VBf9dTxuVPTHBs+p6mZ9hBxj9Afp/MteQnxtTMe4ivPOiK
M8COHJuANILUvSEoJM1PQ7vkymU66jJTTCykPC8qpAI0qt9D8UrNQHLEwPpqYZsb
Z2ocMfsgEzBdbRTNqLDc6Tu0t9M2baa89VEOgY+LD5NJGQRoDt1mj1hYJTxmwPGI
fFgCbA3LgUsJf3uah6aDtoar8bFYUSRZGDHXsZFJ2eRV4nq3YK3nLUjtINq/7/oL
XmGC+9hGR7uWAElnbZGvrQSyS/jcN/PckUxrhr96xBNUDiCOMXSbublFyA1aAwCd
CFzR+XpkmbGZVT729pKaJHwnd+ryl1h6GZlh1sxQIunkww1qBl20mWH+HYyvVSpb
zX4kacs8By4Bf/jRkdTxIlk/b7QHDF+e42WW1ehVBf0agXCq68Fb177oZt4O028n
T8v7ozZOWpPBiS1s1DNdiPH3DRfZkMYFghUENMLbO7ntPC1D2I07SYAW3+ecwH5g
N3djmn05FH+zzFSvfN+DZpRUPJe0eMPwTC5atxWnWakG5NMlVA7QWTGZGhc5UIPM
tKmWR/zKXqI322x3OSZFIapN1cmOSmJaWFrLpHs9CsJ7KJp/0JpO1YQO1LZjtKlA
N3kCFDnC1yHqVEcCk53Hk5C5n7ywQA0kyFcsRHaEFSNPgr0udnTwmTLhoFEZh8yG
UoEUyBA6SQuXr60qML8d6YeBo40HCkitA+7uIO5Ig3+dVsYmpHKV3zl1PIK1cRcx
sHZgF6ffsqekwxGq1XB4Tg6Y4utKrJ4vRbXM9k6OYK66lm9S+AcsiuSkesy8vxAM
b3WQmrh4SWDncffJTIZrOfxLMt6MzScEkS4WDYlIP9NDAzPhunzhfaXROHUqcDF/
UwiQloIcc0/NK+ZkLwHIBYSqX+j6zodycPcdZFCN6DuPrD3Q3lf+37RuxaKYboKD
RMAbzW/DK+xiSoqwy0MOmTsAq0asywdhxhLVovfl7efDTtlq1JmqQlNjED0arxqC
OSsDSKKwu11HHrK6rVwlxXkXhAF1LNZwMqBeZusxsry31jbcasEFHuGBK3RgzHK5
x0cNf0w/PDtPHDVHDmXN9O8h0lU8B2NQbbqRCwc5Deg5uvjDE47E57IAxY8bNhJH
ZQZgM3o/5JOwr00RnFp98XKFDoeDHAt6e52QAjMhrASww3kFr5RWtRKAczIl56Oj
QQbX6es+O43xmBLo8t9lIwnxbxgyJfmvieAtXd5By20vga4CSlcgAtJYg0dJLEAR
RBoIVR0D1SJk62NG4VpdfK80wT4FY/WlARVKdNHijb4QEO27KHq8/Isy5/IHvgj7
uQ/9HwtwVmpdqbqMk+LwO5+JdpwOUDv+PdXUSHuHj7kXlbuU/lvtmjmYnhIloSlZ
pDjJ+CSGBsrxuY7ykLRJHaLWHqVGQ8nat5gRLVwDwGTxvRkZ7kZp88sLcRAZ/NvO
qgnpr7Mdlbq+l4e/3zUYus87eI+lzTGHU6GZoxtLxXr6z3pNDQkKUzQF8s8ppiec
pw5ZVgUhucH+dgmf2/CXW+Rz2/uJbPmPAaTctnewvzNzze4JODV4USAWaF0KbYAG
atEg7e6AiELWGSyHoaJ0RsSGOoR5RqEnstML4f6b1OGP7lECBMaL+xRw3Vu6J3sO
iNFNAsMA74Tj9c89fhhOGvY719wGfFtrvyfvpXBVxpTwmy536KRv3XMe8w6XTp7C
C6SSd6Wih2wzYQINqd2ZOW5pNdA6XYvC8JPGMKWVphkAiazUPXsN80L+gXYEAsY5
7BqxE4H2jyaX6qIdclQwifmrnhbx1NrDJ/bc6cocMuDArfrsjAhqZkvbzCtC4mvh
jmdkjqSpt6wp2Nbfg5s9ztZ133hq8mkMfE2VaLPoWfAiUeWfAFLRI/p5bQhcAIvY
16Pp9YlYe0l4UfgbLaTlS5sDv/h4yhh5CJgrNFXRfsQu1EyMH2vfY2isje2wDT/K
/7DEVEeyE9RAlRuaY2EcE9BcgbQWQW0grRSVsqKUmxra9RLIMLDPHxC06hdGfe5d
EypmXQLO3GJwZTtlvND1oCWJVNeiO5irYfdUqxpviTEjSGcgiAsxO1de6tcjxW50
8s/N0fLqodAi7HUOK7dBF5PM85VM/tQGHWiVnYYiw5DxSi2W9KtJHI5ZDx/yG12I
Xad9OER3hWB8uHXK4ZpgnVv2nVb9XF5T+G2USNFcYOoTPJMcH+nXL2bA/JpLovbL
1S93L7AQRFN1Qe4qhe+H5jkDKQKma/+7WYtcW96rF91NoXfnprxcHLap07DDXxd4
8ILA8pWXnpkuFjrJc8uXnGygmrzGaylj6zH3o3fRD5yNiQuTJbbUvc9LgmOlp/BS
sauRtfiGm9Fa1fDXRZV0LwhSS0Biy0J8u5jt7uiLu/nMdWjDQ0enGJLgcdVXncBl
yRJIealhdPCx3LX6YKN17a5UmEy3g8+g7Xo2jLt4nIVenLM/Wt+lXPWhKWkJoNHM
0DehJoH5DpM+zIgoQlg7llRZqWGfn1kQrquQ+3TY6kojs9Gw0Kn3IYi+ImnHWH60
rF3SIlYq9f+Dm7qwNJ7vtXXN4CKZ5kdz78470nk7ynNyXQE4Ry0SKt98hWfvMREs
H1TUBKVyLo1J1ZuUfD38pc0vfgv3oP870GC58qg65+0AV4Cg8EkKrz9z8SYgHPnM
v+KFHPFwL55u84mWzFcv/VxJCbaWv+o1m4yVApX8qUcObfw1IDdsLVfO5t2kVPx8
j3vICace+v+HcAbiQHwDgS73+mnJbNpMyH5bRrZcJVXnYhxJMgQgt9fY0fgIc4Jw
uHOx91dHUD+LAI6/QdUfHAG1OJZMv83gIqeqn94ivGHe/RaxyQHa05Seir1zU3Mu
X9IOor/SwOe5cOxzOsWAf8nQnKH8rwzL1ltJQW7lS+3IdUQqCgb1Iygwfz4Qvj2o
YhXDl9vMQzr+uMADxM8NVxl+Wq3lYzyY/0EcEm3cv3cZblNEnqyCemWx/gMMf6WL
H3MjH8BQJVxNvIqpJTOIRoc/o6zqAQfsYdV24fREGi8C2MwbI9O5au/Z9GtaffXh
9yejOxsIGdSX0HU2dAgaLC/qt1IrnnK8H6mVoeIkPq/l+gwo7ulwfhNfPrWAcipB
u2uLuDdhk7xdCgMe+03Pors9nArJXjEvK7BtTqzYAqFEP9MlaYynerChGbsoUu6C
FgvVWD56o18qdmJek512hJG27jXWLEsWO1uYdK3/Q20RcGA2MAAaCSoBPSzu0uu6
a7vDzzuH1zbWiPKZUbXc+nwXxwh+E54UmcKY7lZmJdjt1Vi41PxSTKINWVr9ZTgY
y2ndtNBSDIBFIXf9Bn40vqAkmadNo3Ftfy1S9RMCEn9eFFTnWk73uH+QKeMLCzdF
df1LvIfzx1OYpWTiN6Bd8t4IIXmDdRhm8+s3SmXIGdXHHuQdGVXn8HVxKpZPOkXE
D68FvOIDtDct02P9TRXd1ZPRQ3IuAQTzIbOdhbFCdmW9rd/DabWpF44QbuwEWjfz
0Vzc7YL+/nTL0TOgjEkJ8ctUVxML1LrdugAZkgQzdbamoHKkozoyBBB9tb2/AoQZ
gEKTQFRZPdEWqRN9GHQYoPoT0WPgGVjA59vUhlsw5ACRJgExt6HazRaLYY+ARVgV
UPnbbvfrWhNBygMTnhs05Md9Di4uJgvNlaAeDdOlqqaf3EvM72GM9srfjOP2Ld4Q
smsdrc8cDbvxhKWXGEIPvq7AKIyYNN1R+s6KZxcylKxX5DhVp99/eNb5uZb395Oi
NCPLrcF0NC7GXaILT9I9tFe9p4DRJxP24pYvjMaZS0R35J5msXwP59DAKx6p8m67
2elIOanNjeUgiY4JvfmeAgXUDc19hErznH0CEqtVPpWsNb8JXi7n5G51oorlNweD
z/+nw2tdc8+KGqY9nSDc7dGbL/ac6HMBQGuQByZRZ41mSsUOobpnkKYcPdMjLsyh
mhYYbnjYVfLWLovaRgiawvKCwzq52z14KqhtMLXGFdH2amCNN+3wuk9BCGjBDzTf
BAu1225yZSFflNHxUDiXQcR0wQx3vnMwGdJ6/Y9H0+VQ8WBA1yqYWHa36XyPjZcQ
3TRUftLUBfL8ObsXYzj41get8z8dkezf9dgl9DQnTi6BnZoXZcmve1BDVs1x9UFa
rWCEKsP46SNdig08duWuelZ35C1vjXGC545pHV6EgfLLXlKOv/MGYE6oEGvzELls
rCwIgTGJuscEZUdu/GhTOSstdZ/GBvYNm2GMg0p24rnj2+y7D0VhJoqqXIrEwDm3
6i1M3NWN1NbiPeNvMPrkpstQ+uEGf8n5ThjsHcEieDoyiSmRg1BSYqcpXskx0gBH
6Z51tVCxp/sQlyfWoifZyHs3B3GWHm6vleMCqQxQAiQFPuiPDmLoaB4b9gdAAV13
Fvhnxk8XyghIg/RKH7LmaOflFzd+nyfF+6fukYNmj0pDpBlIHAYoCVkQddUvLqJD
rgbFypIB6jkCSY0vhzglyUimVm+Y08vw94WpwxErCXqwxwdlYYEiWc6x1w0BjRyj
fw9ZAKrCdJZzK/Q9Kxw5DJOK/suWo9X69qb4TffOoVQWSyxYUVsxdAYEs57L2BVz
T4FU3CKDS0qcj0kUBsYnCHZ+vopxpY21D4A2QYn2IYGqnCKOacAw3hIabVSE4taB
s9eFNCXcNA/JpQUHU5EhvqzKoFL0CxTUTL5jr58MLRLmNYmRZCCdkwRJFv2cB2au
ptTupYRvy31vH6i+PAGeWX1fL4zfQHQYIEf11Pekhg+FeP9OqSXbr54cCl0bXTKm
57+uLe0B03MpwHPcBhL7x9Rwwtn318/YtvHbA/LqroLlsGZyCt4ZIq1iqK4Ijg5d
HbIk6JWTloNl6nsZRDGRyzC0+AtUa90b67ogF43ginXjBEszQayOQ+RJjgwZKo+T
pa1nBguHmWHzep39kT7ykuaZ6JC8XoRJOU9MA5ohcApkwmdcMU2O1b6HfOqzaY/0
M+mquTdjeLXmOFh2P/mB+MsSWgcEvzNNf9+hJ3etApJaiTrV56QpMiQUiN0fxyF0
xH1nn2+PBZCS/mp/Tu/DXNywPAX2l4fGldfGFOp0JXs5tRzaPoDwHW7b31tmQtvY
EGfDfBMhACO1PqW/0/HSI9Ub59Io0cL0YVGXZ9GdfNd+Z3RAdxglyRtl9V3E493Z
QjBiB60vtonA7Oj2Wdq6c8RMlKqwVISrYKb8InbjQMQc2ET+9AOoRVdERTt+C7Hd
bU06jLk/sTxTe8AlYCqcIIIYTGepLEAhWY1qv3rj7Xc9EKqtOdw35GeRE6Xvnmup
fgBHtR2g6DoiMKzHlz+XcQdSqrZg+8XpHiPuJH4FhW2zIo7cCmJXz90MacfqtDD/
q7KZQyLH3F+a3WfbREQTzEgX47M6R+2EnRL2KSVztmSgXAL2fhNYXrdPrKF8B/Yg
mRvNS+kDCjMIGk5gRVjNgRgdbmPAHBjX5KYM+/ovafMJCkUIz6jKDrAf41oUwAYs
5t9cNiPtp6ygjd/9nrjjBA50ZtzG9aE4vLn8rrgGS6c/7/IQnlQB7z9rPaveSaD1
cRsuJKjcSTsbwymnDRsQ7vc8vjpKMTgEM1gJ4AQAVuiSYRO3Dz8psaznVJ4/eKAb
GAideShPcyjyXnkq3jXeHCz0HSQLhNNbA++xGQwyCbqoxAvlpZxDV9DvPrjY7WwY
4ksQ7/U6Fu86CEYdmYX0vYEdbIirIoZnND71s5GogqmG8PJbIZTyCTYGeJZyuD5s
wIPzpaHBzzu0L7arSKiAEt3nvk1aUMf0uUmHGrgaLytLJZylnUUUiUcrM5pRQVTA
CzqwPCcZaYM6GknvGaTZuFfO6x9YlIuQz0bIdyvSyaThBTSFU54vMf1qSNvK97eo
fl/6w1FmMarSC4HZCSYf+YiYu7ZQ1GKnVOw1IUXPlKJccrq005dkPrO+FUDySVNs
i4Bt1BotGxSxEYXeLeOWBF9d94gOwCQcxrEbsZC4fDpkWZyLp7IyMNMyvHSv8rxX
XOwtaUhlsJPrgUKwIHTF3AKGFSYEw+0VGL4GDRUcS4cBIE6v4l+L2uMxN+i0yk+r
yJeBXOb4eBQa9a0jId1x2ES+LnRPXJsm0pN+n4FfeQL1AIfPAwIOzu68k+RdDiuq
WciLGBtSntrtrlfSVEVv+8F2+obPX4vvdW5IxeFxnUd6rzZCwAWMq4YXmVQhxLyQ
e1netHecprVy8REMVQ9gf07LLrwy1faoD7QsiI9RHtwQ4g5DePCvyuOqVWQhQBrJ
djaKgSmYrr3xtlezbzg9I5owb6fod1nvCIFpQcDRD99VodVxW0xCPTiFmpPlrdm8
/ukGu52nSFwxtXHvlL8FZ22ad/6lL85uax04vnfGkwXYeuKh6rjUjd3iTqTVyvX8
JhkqzV/oUibMMVkERuIAnQitSfRir2xw4LGlR3drYpeU7GIZjtmdoQAxZ9mKHVd3
QXuYCrky+3lg35fRnHNs18vpFeGTZI2VZsKz3/ceuXrJgDlFdpLn7f5YDHuZgf71
ODt1AZ+WIdifZzqupHthox4Iby6dBi27nRX1fseVojvmlGE9vsgSiSLbNh4C2UFi
2uvqLAcfnrjOMYaZjyAh3Ye6q7wEFGEPQMek9QHjSUc9SOfzatvwWP/yeniQU2hd
P48gedJ00YedUolt94qnGaUU7SJLsVNB5Q/2cuwHWEh07+yDGNEaMa8LB+QX/kX+
Uvx10BeR7iU6BQjGmwaatIjTK9lm1wFXPN9MIXWozixvB5wmR0SWZD2jFaiGNSMn
sIOmok4SZvIlRGn+V8TfbyrPcWP5kGAfrS451brwmcCWsdRoKcmZAF9xQ1WfNtkn
yJlbCoU62EuQO8Pnny/uJ1KzBhm8LxAbQJCU7uAn4n8x4/dgsYpOIa7zPaJgMmWO
lnJfoM1WXBodbPcUr6NfPyvSujS45SQcjRgbW+ZPnRAVgTHmOm7DDLVKirbEk0Uj
p1VnF8219X9xd2YySMtVU8VY8JeIMh/GM+qXQlMaqnXNOX545MCkQa8+00xYaB2I
yFB5SEsN3w68LqSdBdoFu/55QMM06gpaqr40mO8iddbtuekWh0rRYUsIHW07gGK+
HIyKQjxrRJPWKP4HsJe3/ULYRmbd2hh2m6U5QKSxRejY8f2VUcEEF2n0X3Z/jTHC
oXeNIM89QAsboHHU81zcQZEpjgjUekl6msSClao2EauGy7TjzXE/TuSQ6lfBJxNR
sHi0YjOsJXSkGj67tlLzUfPlff921v5+fBoiWNkZpGHLmkGRLlaF3GNXSh9eWaYD
Lan+0NbWzl4SJpi3PfM8ntflOmuGsrvYPlkdhWrGEdLhM02UKZ7urMidNkov4ELi
puQ/d/lo9u1csqMskBbKfcpItXLxJPio8OWtgIhUPNkNrV/83AjbVvBdbI8vMNpD
z6IZrPNVHIpoSCargothIG3vU7mlQfhH2sDTIdhFu5Jv3DRT3PFvAd06gjVSSKuu
j3mqskAJO8retCq6SHf/LgQVn6IivIQCjZhHQBI8bSIamXyvFvK83ykp40vFuUp3
RhxY8wxXIWW018ETnLwhckixgP+jgIocN7h0N1b1nsj5dXRl4TB2C/UJwZ4elVid
HjJPM4rMOIez9XL5gdoybkKphJ2BFx+PnBji3RUwAUanvDsqcZwa+y4q734Xgjbz
MRH06yLpFLGC4fvQAU7V9C84hVVeQaiYXWMcvDXQq/lA/p0Y8tzY6YQz+I+9Q0if
KEsye/i8IeWTpJHgm2fpkMUQ6essqG3GM9XCcOk2Fx5WCVtDJkbRW60Ioh36lsPy
uEZcRDDC1ac19ehIy8apb63CJCXll1SrntIvlfo6DOBb0PdOYnWosaJS9IWzMeUi
n/L/gZrRTE8aywrufRS7tJ+QyUlqBiSmPqmf2O/CtIcZJQNUhdyA2vD2IaNaMnBb
L15fYIshEiVKFQ10B1ElnTjx5JUbA//SxvDcQYHSi6oZCTA00fRHQbSQGFQ3EXbN
iYhmmFyBtXqu9ua4P6lv7FZDif7ZdOKXRYm9UTjpU2vBPOMsc6EvCvtb+GJc81hD
OH4wVZbjCclti23CQNxWyrMOhb7oe/BdBJkMbTEgtIe3CMKH/i0xAy9OOlkfc3jv
xCv7cDXCqZsKY8iVzfl9+20zxdcKmPPiP5mlXaeH63s=
`protect end_protected
