-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Sm2/h+OcKEaqHOaj+2TZ87oL8rOUSLws2EAN+KkO0E7Ui0c9oZSWwJrpq7kjKjIa
XPbxRHyIyJtHjns9td4cDbZx7rqS4HAa+22eVx3tjl+S3KSOnSxlROl3Iv6r0lZS
cOgs1f19qmjQvgQJcu6D+twnl/DO/507vYLeMRtU0tVQDDzmjBgfVQ==
--pragma protect end_key_block
--pragma protect digest_block
YT9fd6rnWdA2qlY31ivrXhbsDQU=
--pragma protect end_digest_block
--pragma protect data_block
llTlrYA9dNzEci4EXoTrpRG1b45fRYo575xj90AGq7fHn58+d2eIPHSQG6+NyF6F
G3SRkUjpS76e77JXWAr4i4nVgwnN+MDCfcPb/nWNecd2chpj461YsEYthkdqh9fn
LWX7oXwfK/GLqpYwrPK2Hv5x+Y5StNmZbtAB5Fo3eTMN4RXKUiFECIsgnaZoTcdq
crzdNeoM8yYWRixTEPp4gDHnbXVfaswIuu7F5eL1pts+kcPvs9pc+tkUqdp4agfv
J3CLt7eGqwhY/QtHs9nGPtqcmqgo7Fsvo+1VkyagxPz+737oM2oQhwld1+pTBCoQ
jeEPN0zYzAsj8AJGpIOHp4+NsDZo/0/JuYJb77/d3sRgsIFBQcHq33ARKdWogi5a
YhBlWOtzf8myrohPxIvk75kxhuEkBWQViKrEbTjmNYKUMVnZvsyvet2uZ/J6KL6a
tkgd4X8Xb1Gh68lKi+yIa5GkmBAAHrvziV3/EkEWYNlYIbpx83Ov/VbxNCpOzn+V
hkKgiE/UocZaPVUhE80faAhvobfNaRXlDInAr2BHJr0BeErXroynLNj85CLOFw0h
aR7a821K9d3iCd0JDHDjcDTyLJMoCjuQME0VmMX08sJcFqu4DjdAGwpYAE/DC13y
kZ0gFZYGeY1nxktLJ28YCw2Qv6QpiCAaoQdyoicbiK9SSHck/StMLj5To94qTQ8n
9wZcU3A1B6WQPMMSxXWOEdFmA07QvpfXLoIgi+gcS7L20gLImaewEv2KsmUrL3q7
/P3afx3epaWcWEPqZoxdd3YqvMTMqPB7d6Yq/r2VsWEBcgDcbV0+kFjQnWdj5DK1
uxRwdR1qq4y/91jj+hObp05C/QqDS8I3KLy1+Y9OO596J9MvWUOxbm3wonwiVoWp
BbQiEbBrDXBEyXA3EQ+8rfw/sOjG61iHgnS1fWgEBgT1FbZDzhKkesVpSSoyfY87
11f6lypGhyMSXKvdY/CaQZ4PtHw9fOAjg3SMRZ3jcYM4YOjF8GNXFhONXfYLtBQk
OpcoUZZyzDeljJyQ26G1NXzHrxlR1MceOxK9jY43ws5/UKTiZNyyWa04RT2mZS/0
oPaA45xTaU2vQLReqBEyyKyKx0NoOBn+5sgiiPbx07H5GOtIP3LTmGjnWHs7Jlzs
jgcKKQj4yghh4Y1sLkOdy1PZv7aB6L+NpaHxyF/8pDfKRNjCERCugDBNnyQJFd2b
mSHr6zKt53wchvwVyaKyYXAwrfHSUFK7+uR5ALTtIbybaATZT+yjVB+VCCYtHy0+
7kJuG1vWGyl0aD4xomFIZDBXT2rGJb7D9f3t5wR60ZKKKCHgg2qDhjvwV3YjesBH
C6QjaFODgLRAJ/WHS7a7HTZ0n6OkdpUtFLyu0fq2mirK6z1dF/itg3uJ4mEw6zPL
GGllQezxi77rqjPhASQHDMmZukEXFDg1X5IFmBvnksVpUtbDNdUFdLtbwMNBSf2Z
KHgSPCF8k7ewZKUpgxa7uFXNlbtrXdAjVCS07EDn0Y3k2XE9eRVxyP6DtEdRHS8d
ACimrtmN8IZU7e+1+EEnRZ9s8D178Iw+MQUSQaGB4jEU2IVZx2XgD0Gs8UedAMEM
akwgtyo86mGBpqDH7AQtm9l/I/S/M3TVDhe2w4bWgcf5wyzyM9wgikhwwbMACpgr
V57I7mo6xudcl/jcIALkbvovy3HwZIdF2UrxgXZzq79bOTHcqO7s5kP34xhmD+6C
Z7j0zFkxRK3VoDVKfSad7QPR4jjnMoNH2UM8fVnTMyBOe7Mu6FPosArDcRgHN0D8
MQg3c7zZGOqvtHGSSBcLpCVMBDiE3jfOGMPu+0uU5wazOvEBlfF0Mq9OltEOy1Vi
3tDDyj+XPPCYrvDveqOyVpQONaag0rw51a2P8L70t0F+4NNaZ7jv+dharCmv2gtt
ItZSn9IGuAw5HHF5IF1ocogV91ZjB4vpMpdOW5JKp36cSSWZpm937L/bXgljg/Q4
qOyZbIKFUwb0JfbXgHeM8Sb+R4g8oDffltWNk6gVDE8ReEh0JUaPXDSP2/jp85Jq
r8hxxaj0vWL6OGXVmiLmLMj2FOG5cAuSW0aBXM1eTJr1l0A1Cgrxozyb8a1ltEeq
nudZzUhMWV690VIC48pYM+48XC4FOZMrHxX7vJpLLd/D7txTLvwVS1Zsx4lcvhJg
1uzrGxoJuJuH3nXb5EGXxukP9KgrlLWdgh+T99gvkPCA6/pd8VhS98V2iUv+moLj
0/3cfzrVo2+zfYnC61Sa+FCynOXr5DiV+B8uwSQ2ZEFVyPs6Fq9gRX10IZ9gT3FM
ILAXEaFpXUTjz8yxHUpRYTIr/nYXLwQ9JkBtNj1Vm+4i0vuKs9QYsscn8c9l29pu
8HHP1oA8dgmfhenvMCJfYgZmYp2PB3ebx6YQd0BGM6RtRUWvrqUENyF5ga1VcGKC
pp5+fmQr75jlZr/t+AYKq5LwIGBc6TOm/fmEG+pEx49LhJf/AFC+HTUY5dhi9oQ4
B8GJMzm8tvI5D5N9uysjn2Z84d5Fp+C4ttFN1OqSBFbfYO6P6cNLWvkL6fs9KF+6
BLScRy+/AYkTsA9+7ORB1FZwa3QcSXRueSig7fI/kRM4enlxO5EREeuLsJIK4cIj
F++4vpKpBBcHoU1PPYWYwL1TQMAFXZAzCcWNk0sFONDdSR1genL/Oj/H4ttURcCr
7dSaYDUpm1kLA0DNeLFV+tc3aLjmKhLMcsOMQvN8ZzEBMDwLcZ0tDOnewNj7IGrm
91DwlcFKBLfqpPKHZmk0AI/BlWZEsABrhDWwNP9SRizZNLUoudFvDkh8fB/sVrqg
vRmzd5FvVU8ugMbyB+JlKsTeECYqqDMxXdZ3SlsQT0Y4fuVfwLpfGFuICIeW2L+W
lhUtkRU3rKhtdIuKWY+UtfBsF75UvniCFgYCkgaG9sbo6duxi43PrEQ59x2uApww
R/WbjFWBfyQumlhhcUaN8urqveEscaAMMS6ablKbXZOiUSAxitbZk2CCMNKS1kAh
EuuELNiZivPrVLySN3vOt/gqis+4Hs+2HGwO/veRvEWRXrUPuTZmd3YWYrIxWjqG
zvrdGOPOetqLSu429XNqPqpyICARGCmm3ajIVSMpyAr4HDuTg2yjrjxBasCIYDv0
J93AzTd3H4NRCiGaAG7o0vTk8bG7w7ZvkdMqzIHkLhHkul/AW/VY1C6qj3crKAak
cmQQSWVM4X1gYK3CAmKh46SEZdhYjaHp3RiK5AX6EXbHqpTrqOlEz9qcEVrQz/+G
AjBjucklWGfMQUmQi9EwrwU5u5+xkekHYm5AmKQ8t/43Ocy8mRgVD8rD/0Z20MPK
1nApzCi2A59PE0uhZ+++oCkmnQzjdhRVumj8oBoq50Zvplbu3UZOkr62noBAenIX
wYdx13BOlZMEMQV9TrBuZTJCCcoLqfcYk3rtw08DVr8SWCgNXg/WyIgPOtondSaJ
x1TNDs8Qud+4lXuPgQvqzVOCCOaIeFjkG41l9SA3cPSxH6ElOHlVGp87JOcVc90F
18Hi4xH400/UFlFtCXwqvG+Bt9OmCZWiEGjx65c5E4bNqXlQOawyjEZdohlTIvLK
Oq+h6ElaPbKXH+UWreMChhRhGTTryIaFFrCW40dESNpSMAa+QueZJDJB2csBFeS6
2721BZKFYPwjsg5FjayeKhCwSFgXPbH0Hmg9A9r2NXT8R5qeGO3sEb1qvQoEeWM8
dSq21rS0QtpPDKUHdPVNEtDzcTYodADtKtOrBsefUlOyImrjYSUBzHRcgxOUYKjE
EVYtlKGxYLDoOtybZUSqpCWkST6R+dWK/8TIuatlShPozG3YEVKnL4bkFp9rVO5w
VCGPXEBYFwpIys96xbP1afRPTygIyc/XdGWdAIA7ukuwd8ASCPel8fzwLZYC960I
lj+fBIeeWwGHQxbUiERLUbjClowbYQm0yZOpbnSfJdvcE2P62lVlZ522Vc773fX3
LwO2SoK/mWOvlbyfhSUQ9xlb6gcmciizFITnS1KCf6DNvZJFbjmHhjZTtwNUJ8U1
HEKQR3a6OGh/p8zlYKmyD73L+/vUuiJvpw0iDIoIf5B+TgsMaiR0QjgLe/nqjcIr
AJ0RD1zS3Q5fKfw5pWNGvHZOfZ7cOKdtFHtJ0Z94hYQcLaQ9vP4+EO3glYNzzRgW
V0BOLyEXiOyw8lOYnpXlxjfB+QB7+/xPiM3PTmxGxFHVarSp0FVh9flk7z7WsUBN
UPe6KNCNOJ8/bmz9noJi/+AMbU1NknucLkC2zkn4JU3b/3x29Mht52ms8vsVRglr
ZvyPhmuBEuY4roEGyv0Gl+3kRl5wZtwz6m0l1DTDrNNL8gSa1LdWovRPI9nzjx0z
RPAU0uuzxyaJOBvnPTqP90jGjHJjKlPCOSKsc4gS0q/UIoBJTiT3SaYY4NNeQrJj
TTVRI5Siik2na+YWs4lIehWYg4mL7F9EB73yZp7Vry/hjJFGBlAwbo824v/woB6E
hvDFSC9RO1UUYN7H6rndC1urd7ZEMaY7mFg1RviYj20SwfXCYG270WG8EO4VfBoa
2p3b/LFuCHKg5wGiqz1vk7aVnaB626n/o+B47kdqSz0FGILc8K2XglTJ88Vnd1Ah
CRNAa8QEzcRzRGngZvazLmQqfzwvrH/xlqjm9QQZZI096VL1Fske8bTRmHpiSLY5
1Vy7ORcO2ypUD0IknV+HfPhJLHr3l68kU+6yzrd/JsVGVLXDUUxkDC6ULHVOHu5A
0fWDeY2gTHesIrcfO4oRy9XS4HZgvgESsEoolBgnS7rONfYr67If92XV3AGB31ss
jq8HD9WXNWvVJ8bHGMts++1PhMgRNUBiJ35pxiBuBzjRbaRP5yBf/ZEc/a803MjM
cWidLMGX0/0S0iUN46wCmcFqwkfzgRS5BCcw1+B9xVoE8bovtSlKarV5NiE/zRM/
iL6CikowMARyxM9WkEc5wE108KEAAF89Ijjx7XkazMMlb7h137vPWxTzafO8+DFd
IzhwJXdXBhBs2Rps6r8z9XM9tJeBuXmZfXcaqiswLZ9TLAQGLncsNFEquTeULjWO
hgQX4GSZvM5fKmsWgPvV23oU4oYR4ZnjLQyyg6/pLQ0nRBBLQKbBTk1T41ZcMIaE
RD1nvUF1EcuuelreTf8jNWTbxTRE5kd8Q0IVs0f3dWHQNG7lZWOdKHe2k3hPuo2M
3zGwCTXAJEzP1fG2tkeJ35UMF378HqpUBHJ/7svcpJdKw+aNqjyon/bAF22XlCcZ
BmZN5TicnVxt7LuroPNQtvcvxUSpeRlJkSNM4csv3E5dkO6YgdoXPTr3hlvFNNiw
7eVXbC7Qjx7uECvplZ98yhUS5jGFlYhOb4gFMG7gR7LmOLA8EoWy9oypwEs5IP2M
0TEaIKWfR/8ZAeAH/F3SM4QKXZMHEAyW0VONk1lHbUnJ9bdUvi75QUmjhaY2cakP
6W71AA5N98iAjhegNoIOGi7TamzOsXHT5bJ/+6K8DGvzBGTXvqJPYvcukMGNPjfU
PlAWxj90phtWtG4AJKyrNc9YjJmtELEjrp/7o4Pry0DP4yf5Zl4+uYSkQZDpGje7
eLJ2WAZ0HofY60/pEBw5YL8p9b+02VWyJvpGpI7KDaiIbGBLYE9wZMVxYKAO4LsX
ZUNixUZbbOVyA5PxLSG57KpUF54Bk0qFoKYReEfy5tSZJxHcNCvhlNHt9pX6j60L
lKkV8Ig/ucGRd+KAUu+OxkaJ3XjBxGlbY+b4wlE+89GCS9u15KD9pPTJU7IAOsUz
0ldgdhQACWBW5EVKDA9fV+3E03zFT6qH9cJrQqswI9U3fJU9H85wnb1s5f5XRDFG
BNyvwuOiIK8gWU7aSG5hbtyjTyAqk92oxx7+Oo3aoOPK05x0LKBThP/NzO2bnHtm
BOhRW02mZKT4DebteAajj/Kzk+y2jCnx3OubVVE/52mkFa/UFX8YbvrHrfTPlAi1
3l9mUEaigjRiB/PfmZgbslPIxaDOx98ZiQe6hyFcZPCmqrG6aU9fLXXsHbHRDn1w
gCq2Fa5Ao/kHzjYknNBM1MwlNfugfzA+zYugQbk1KJOhjbowZaLXXRm+I48dMnn9
xtewbzwbJKVnBx6pe6Y88mesiOXUJLt7AGc5Yl6jwjG40T7eG+n+7zU21fpNs5V4
UMWB7HkzCJ+/TjNt7rtqFo6CWNqtHXZJcoynDEMD1CmhIxMJT5+Zw0VXhcgTd1uA
OlTWJfoKWLyU0Zc9rpWr/2hMwuHFWsiJjsCLbKigT8OemOol7vyw40WEF4l6XI3/
1OPyNyVDODKOTOfu7s7PNy7uiBFJeQzMF4VRrq/iPBTno7lVnA55PRp3a5ZiI668
XRCoCbISATBrhnfVB6AC4oBi53vXdikM/Vl5r6AnmlqhQDGZw9NTcbjQBCQLFKY4
5cQ6KNsnIEa5H924ghiUvyCALHKB5Vfhy6ZYnQa8Hn2FH3Y0k+KN3S8Ng8QG4qXn
L17JrDKnLCKfFhjiAbP35BF2MN5shQoctTgnQ/bXq1jWbXqPEN1iJ8g4uzn72h8j
qYH6vs7mN5YdLsbmaWSewZGdboujmlnPquK/x/STX1ji/E+/BSOJSaU5KyAFa1p/
D4+H8ICy2YjXl1Z7hpml+ktZyHIcE1qI7ZEfFqJmHq52Ji+T/o7sHVOcba3WclQI
Ai+Jt3MSeGE4pLNAV2ASicEmviQF641p9H/ERM28LEyb5dIlngB2TvWUfMD+oCj4
3FQJwRzWuAbtm6/FNrTDTgflQtlzLBk+MeZwA8QTP0IsGUZsHoEIpPY0OUdsKgv0
Ser3l1ORYfYt7hHYLvE0LzTD8gUvQiWEya5HN1CxTzAyzv7UWk0hkhnpVn4RIm63
42E1ihoTZ1NVV78VGrfGnSOjh2++MtAo7H0RfHvJZDTk/SJs621U7rTb9bkSWtax
e7pcmufTokaKeQWL+vo+Ji54tDIyjNs6ILJ4kCTC6gDmK4q0S9GaXbe7MuCYGITt
uhg9u4d8sJN3eykYSGpLjBBzKQOhdUBpVYYjIKBVUjtTaGFvd4w6XYtgch4IfChz
Gv5h4slQqyagPU5s2+MOqIyoiAsF8Ag/yjpHcD44S1L8D4YCLsr+mkcoXUTEDsmP
QisU6Ug2oONbUYhZdP6OOMQM/Ae8L4djCXE79ZHjUAaiQx2aGACnlnMZ1d2PLG1A
iwxjDKfZGkty0jrDkEUBQsN2jEyvCrQNrcGi9Halv56KdfioYPE486dRV9eo/+gp
gvvfF1mrb667KXf8TAGcsyY/+kTyXhfrrWBO4RzaCuou+Sp1nBvzwAZJNtjK0mhz
9rGOaK3H2JCZY5FVBL8kDWlWrQSgoKCnkOFSIUw/7p+H7t99mf03ZHPVXXkaQ6nT
/1F8HjQhivFqGQBVK23pe80OzvCSMQE9O3C9h7JNSdIPVCfUWisV9kbRGKoFMimD
Z86C1+Wvibz3B0a7VjWSZVaTr71xkJZnv5T3M0r2zLKqZfXVy3qBarbnJyeP810s
7vsfQ8FBbPhOkwsNmiDTO8nQ9Dp5HhPZzjb1iHkg8tYq6kx4ynXcN9PySJfNUY7L
dhvfbQDB7g8EQsuM2LZuAEQURvYAMw/IgPuWpPS9tZBk8YGrGaKDzfr0gIEz7B8E
TPBzy65ao4dTEYimLpgoe0VM6N7dc3hllfnWcXRjSoZVv+tnKgcNKK7cx8paTw1T
usrQkAGe6fO+4LOWAhBLJ/3PyCPls1eFRUMZ1fl22IkvBjBsBeLvultL4NanXjjV
HtUEs+geP04wdIWKdYcgCoN17HT68NwXAcLFdERI0dJ2ZEKxs/894Iy0Awao+Wy1
v6w3PZ4RjaiP0rY8DLrQCx/gj90lbTCgkAkEtDGpcUSqwcHOUUstWdKk+at7wFPa
FbNG9PlotSO3j69NRtBw/LXwcJ6/VnBPAbd/LkuSqqBTcRHnP17OzrxGck+Yf57P
M/JJgeVGkN5yDlYZ7Jl44f064MfLMXsXNpwKMKPOlQwhZ99irob1DW9IOYBLFKEt
AkGnYq55HVPTEmvct0gKgn0U6vTDkzeQs7KG0YwNgv7j1ug/4kQNwDaKn0jZfUPY
T1M6YTlYugUodXbRitmKakeLX51cldu0WD2bewWmVtp4tJzSimxp/UXpxIFS4P5f
Kya3pR93zx/RL5ms9Va0oTXm+pY5AgLNSa3SqlDayPZVkVcgmVOdwyHYjz0y3j27
65tS3pfZu5hMJ3THH6TCXDNIdesnY5FPEFmy7w4swiGu9sqW4ZU6+nXjG/KwM+RE
jX9JaMlYrucFKmRqu1Op+ctWBwqj2T3LHkFIrn1Pe4/eAr1W5UaM47ZPSP+CFzad
Wu7X7m4FcWN6u4NYfl4+1wJR/s7R+RDsT12unvWGstzl6mYmlIL9xGRWkEdZOyqm
8FSvQwWqNeiqWV+xFE55l5D/ZZp4P8bswzfrATyhT1GxJFQHwd/muGUkRiQMm5hI
neYCxN5VG1MG70jyU7YFc7QMbWthIlb3lCsZ246l1stUoz6u0tSdlzbz822oVbZH
9JZ3I0cq0dUETNP6qRBsPqBdBa3O+XgPRVZP4vwt+OB03IkpRv3Zgu36+KY9zKZc
Y7UNSkAPm6DeFqFhFo86c4U25pAlAOKN8jgPrBhANLT4vnimuL8s1z86wi85FDjD
8SXx8DdLSMEYmDZi0V5O7iYpg18SArYdDCMmAd9G0tk9nHEQ+NtEA8g7yisJLTqP
qM8OE1SKRk0R/sdHcDvPtvj/F7nhpPHkKCaXFKIixJex6lSR8WE8Bwy6UHO8WC07
C3RUbpCgr71C8fQDpLDTjqrT0VSjYZQcqDgTPIMhr5BoCXGGkFI1efmF9hlbEGri
I4+xZT1tq8A1NmQVNCtgVZz5uQs7F8q1gC/TlM+y7XTBrq9pVsO+5rtin1pbCkY6
+DAjr0tsEthk8cJ5cNpHXaluYg+4VbZszMrcs+tBRBFoNlao59edDTRD8PNWqwQq
HAdbkAErY15kcR4/VA78fv0WrKGeN4WNHqKdeEAizMMxtrl1/tlq3a+TukXhdnwi
2N6nDQNbv08UAi/Xpayd7YIfrvzFb0L0/YcAcH7MFden+TAlhXwLjnSGIV+BMaut
UYi8pBctJqdIkNmYCW+EA04/lFWniIwnNvCJuDjAKwg41VRY0DoMF0ZB5lQKS+UD
YGtfFD7AcXHyCMguA8xiyYx414CuchM7q5xZ3nFQT2ma+iXR5pZS5F/1Znd3w2Wb
Aei6JdgwpYrdIlzkdMpwbrVnb7BVqiN2BevldPB7gKj2lBQqzswBo2J9PwIXhGRS
9OFzQfoSi96laXtiB4ZYJZATJkBf85/sQcm6FeWKqHyAlfZtUHGy2kjgihs+dqyX
ILhMsgxkqfAq9fejuWKJrS3OMCJd30nrNTb8enSdN/eEZJbPwJQVpAQY5sIYcUtn
FEDhcq54UMBctadBf2oVEKelUae1WrBqOEI5r+CfMgthWo/k4o/3aw3IEO+ak4lN
FUUHAb/B5yXsor9bgiDqBjH1mJUR1nNixm3cMeOOme+/ZISa2Eg5fRk++HTLFoEd
1rFOzddzk3Vj+UQtOyR+D3Bp/BV8N99TBNOjn4bPPXHeyaZOF56EAQLMzasQtB2t
l+S4O1bpgBrwyVshFXJDMKs1ePuQf8vARNu31II/sBk7vD/NuEHykwnwxoecFxSK
ylTglmG/OBNKOMsx1ETZr+FkgqTLcJmI/BM62FNS6TlVLD2Dt3Pfj8OtGqpF87AV
sWdzOuWUGbxj9yiQlkvxPTD3f/lp1kuNGZEXjhNqdhcmoWCqzipwKsFFMK26gC7q
7obYf+3VCZA2lYbyjNU7L4laxsIvfATE1nZ6uvPsEnrdK5E25OQDabIEX9ZR8j5h
6Omd7j+1boehN6/8lqwlLIauX1XshxfuQjrV73b3adEI4ZQMyPnUlWzBcBSrJ2I3
qHxJTa/2jkHq9ZP6jyognywBTGMRyWV7+5D6K18YuDoFUxRjdqIldTJTGbY8kRF9
hig334VoIMlP1T29gNSg08Ymyb2x1rGBNGVmNLSbtMgT4OsS7VRsrg/dOMEFNX2j
oVFkk1IMqJaumafe9KNXcpJNWZw9fFxRLznrdGTbqCe3dTA8Y4ZyHQkFR6fBdOaI
F+etpwXn7/UjUNJXT9rdPOyejcjvPwNjUjU9piAG0xFA3m2qFGteDf0YGL3Xgijb
QgScfOQm/ZUtDin+IYf79JU8iH2IBmuZvbCWIlw28rdnCjqNps8A5ledc8szy4d5
E8l9s8HZTBikGzc3Hj8En8efJTuM758Xcg86zXDXHvDvsCm/T65KlgBla0Abzr2z
owBYBSF1QEXD4FOqguvmQf7iKGg+BaFcqc9ebFhDP1O0UBl9j4mm+0RsnLnSp8U9
Mfe0xj+6M0rkMmVe2tK6D6HGU/QYa6V+7VzWm1NWXfyRrsAfVdLf4Yb41wUHbRVY
dfVBqmU7ZLOukDOVrnq+yxP8YVEgeZ/XE5ZSCEFb9DBG001zkUa4WQ65JImUS49w
tYNlFqpZ3WPOaeWjicSrZRFWlmtQoVDMw+km0I7khsWj4bRErQVxgUa3kd95or4F
4KGv/zuH3T3OVNZkAekQTGjOuN/9zhiZdpBMaDIqkgMzhdOL2uIAkMO0cJLwznyw
4Qj2vMu0CRsQk4xMqt9TGZkAYE3W0lTsS5gHNHpF9X6eh6bC//fbUZoyypjlWCPO
QrbOEeiZ0Eji4hDXgHSq/ZJ8wLscfpFFs2MmDd7QphuAD9QbSVGfWTf7+kwZV6Ep
u0l0Kn7+nC+bpYyq8/keAc1QGYtZpkpby/3rJQUJGnnA3pFi40kqFwqaxQLFfIml
R/5dwAnFc8CXxmGX/Ew4pq/3Iomn9jNh8j3YwawGYJMZuktSUzjoYFmhrhmHmIJ4
N01yYS0RyrTK7EOeHmBuQ8AOQFnP7updZhgWeMwz7XJSH0OMkidFNPJx9B5TafU3
HjBwYxjr6J7fSMQmDePEmQCMMfqrvXyl3I9zyadBvMDf75g4VOUzDeUaH+lp6WB4
viDWstm7y2sEOPsRrWV9AYkX9rK30EdFIpsyCAOaXY3m8B9nris1Jnkw04Ie/Hf1
l2iIuPQwx4mK8HflnjxiVa5FLO3rARKL37XwFcXeeHyVW2T9KCMGzo7ilzLnVpwg
/Z2zVS/Qje6ufV6nwsHyit+ZTMdYYvlyU/BlUv1ciTfhczpX1yv6snVjxBTVXVZl
Ffp4QYP7Rmt8Atm3vEeE82ETr0gONNnpuquJA6Er6qhGnmwokayhkqwPUTj+8IX/
dfXhgAhD+CEnyJSH1ouzfY1yY0889akfp0gXSesUWKm854SRfb05Q6uT9+MexSvm
Swlq4y2EGsN1dhQVyq/tRZcZqY+eC7tk8HNV1/ls0j9MmngE9eRlyr7V4qVagRL5
BazE7H6ewyWyx8pd5ilL0Lm/bZW/eBSmNenIMxCMGtlCClTShbQVKoG7hBDcrf2h
JgL1GraME4E8lGZdDJWuIo0rLY/XO6eeTHBg1gy3YpFUQDdGs9V7je9eFksuJzzF
ceKehc1IZxdKdrFT7ucKeFYxODGOfMeuwmENXAjCOY+AlPDZTq1tpHjViW8sHd3P
Tn6WhDvCMY9eJNE1LGCx3y9BeGY/vg3gGid9yFyYK8PSzY8xqTdZMHU9AM8lje1P
RQyB9UIfn1t7jA/eKMfg9fZzPkDT3VqueO5RUZZFr0civTJRFV/nhc1fjesuKEPl
I9VGnmLXxqcICEggWFkwHXpA8pMxXGP++LNFIq5v49fDLhXqOaIEVx3SASuCJHx+
6o+Ssx/8k3hA3aSc6ytCouRyQ05balg3rzPc2/D1UoNd5Q9/KUFS08/0TC9A4f/O
7xj9QUT9eVSZzjhUciNKsX+RF7HB0mn436eUozPWimn05HgGByf6En7fnOv2IF4L
HTsTgcNnaMxpKt6b1ZkC4upNOKalrsTXh/YYi5H3FU2mXifOcVwp6iWFijFhXiaN
fYQk7ZvbrLZHfDG+hPOoumfx77eclyPX2lLFwxlaG8SXNlB4dCl43aK7ew3RrzLd
5PlYv4rzOJhOceIMXp8Kjs5HFeknFlvYt+f4BhUYU/CP2Sw3hE9UyFmvhQmjdxgx
fF7+TJbQ8FgPi2XNQqD1Sqh5+Nf7UnziKQ4R1J3r4IvdBMA3qZHVTBKl2UikPxsk
TGSMmYVcLG7PkMxaNn0irWKf/P2hkVZzVfmNhu1wZ/HtkOo6lSklmp4umpsxZrlD
Jfamlv/f+KlFHJT8KxKCZu5J5RWedkHSsvlMoI114qLyVAizKgbu3RhhDOQcXkft
cHKHidjHcphBqYdx0GaIVOTbXEiSzGNH1l/78nlF7UCWSGADhNArWG7X1sL0uYLx
cIs1Io0n2gVfO0898qR1nrDi8NWHLP+8FqptDP+mQUpPqQRRzA/4lKb4xuF9+fdx
JKHL8Q6g88hetcJwVXhQ24ekqErq46dzDvQLOUXBcz5txLUNsCO6QtUuHE0k7KhH
XwTn7RcTGsxA6Ckea8JFadsptZyfDySglRiNqjj9C9zLS4pltpH/qLjPPXBWQ3A4
oaaSy9LZ8evgs+J54sRaDutycSHrAbKuzrjWFQMgpOOcitFMUNO1H5Ah/dBRdbjF
OFw7g5I/ahTMrvxXX0dpFVG9S8+29M64z7HScbuqJV16KeLRJ68gA9Xz/SylEBFH
wCNIuNu9EzvwXWnYMdQFGypZ2Wyq7XUc7NRAo9PpeGKf4c+3lMVvSt+YJeNryL1o
XIYTzhrLJxiD6EGpwIByfRlPZN+jd4y671UVB/j1aPAUMz35FUAuH4DmoYTpzX1z
B3Y7xZdAJd12ntrCIr4IQQd/IeosT5HRnDDrf/87fBOgJ4LnaoXZMTjaKICCbeQT
hBqoNl/JKwFbcCwBz0VPxlcwiQhOePA0mpjKg5PbgzxSYhJW6J2UTN+M/Ek2wbOW
F2DdZK7slsMKN9J+DvKrsRc/I0SKaF59F38qd9AvkTTW4215JXF5V+r9eh637hnx
ixV+cVLU+sWHSfhXTgV9BPVz6gjSPJ8Q248BOw26+CtitvGfaQ6qat/ee4tbXOp5
v8jrAzjv91DnSieapwzb07EExh0UmlWHEXXVHyTQ9puqxNi5yT9aYkOSn3hazoty
uzgrTC1b8cmcFfcaPoUqcDZ4vQICJoVyNtV88RGGPlePib50vhMmiMElAHVuxcTo
Tg0LD+mqvFaourqTVJHXy5jajnQbKexwH91GXy3niovMgjxEclqbWRPksl6QPUST
mD7cCKdtkihCVfCpo1k9tRhqzr9WEGib7WmFbfGEtKgKp7F8ATeO/EVwEUsyJExX
mppOpyGjKaKcISPwSLljCPeLl4TBKp7mdEi06QcnJkLsTvzFo0Z3+CFkrEZ6dps4
a6Z4f7qc360Wp8md53kg9pGX3cJga/8yuomdr/qpJYamabzQoN5HKVy3HlN0Pyqi
Lc6mbVaZnieDBdjLQAd0pRMTrTBX6UTC73SCRVGw22bkNjJVMEInkMR0UagDFr8U
WWnQbCdCqe+FTDUuvXBRZ/X1bL/7LuA+bBvJ7VJ6Dodig9eU6UAkTrFX5Q5sSNKT
/Jc/5OWcBoW9EA+NZhfkpo3xnHsdMJGvvpxg+KEsYz0khREfTsGo2dyN56SUtRD+
BFaB3h3W37iXSrnVrzNPdG7pJrWLE1Cir6bdEBxb/2cYJcgimJK5u0xYBrajDh0A
AG5Vi0sZfvIlKVRAh/cRZPGHTkDCpE/x3JhQ174ozrzfaNjnbV1ydPlE6XjXqW82
qwuvJyAd/dTJbsHq+5jOKkbqgrVkWjaXmROCbnDLHjeJvi/Wptcyi59R4fjZmXnu
JXLAYUO4ZOgi+v3GHBSRQW8MjPvKjgVxSp6jpEDi719krqLzm86ycxDfZmK0Kf60
gmbIFCTzziGDcC0Y913udInMLkvd8uknIycFm/fk/oKf6/K3305hmgI8pvZECbOH
zeQsaxYANIEHVAC1FM6fKN1v5O6U9l90iub1NKH2jY+pmbgAZgFWqBA7FH9bl/s1
5Q/Wkq83heBhzxPFNvhyvyoLneSGI6qJCHeoR2PMrZubV+JEb14kkCYjn2DXK6Lg
0v7ZsHZM2LM5a+arlNHqfUOxTR9m7uELxlNYi4rzGc+E1MVYkMNPzKJUPMOT4/8J
yO04F2cqdh6SbvZ2IFxF/yu/eaVA9v9MLzuakQnGrRsPX77+67eih2pVb6hZobtu
BgwVBkS/CJk3Jma7Wa+jirlktvK6fyF+KPzATLsoxYr/jtkWCNV89dvdN2fbl9rp
/IHD01fFPaqlQuJ12xQmR0swbDeWcomD35Vcp5D7z1GDjgTDIXeLN40/KTvH7ks7
EOICTTSFqJVzFOIj2acSr/lpsPE6ErOp2rUyZf+wDGqoEqTg5SVZenrYS7V5Qtii
NRjtwrbD7jdqc5O4S8zCZDL6mcIe261j5RM7jq87r+gTvtWVXX7hFjYB/SjtVpWm
kknHgH1aOVlMfDQKAK/h1PasP+1CXiJyiHVIdmuig0bInAvzyPquus1eWjpUzEjQ
kfntW+LvmrRmetDEuTY5jZD8YsX46mFMcG1R1xSpS9aGeYs05b7OrLtErPwCLvIK
6ZrZev59p9f2gkOd37/6Nhnr3+TYBsQ37FnSQ5PMIctg9vssjAhmI9RYLgEUkS9f
XLV1YRTQHTJvQDWT74pVak379d3kmCrsSGC5PoR8xPQ/N5XLvp3izwlx5HodiZlV
q8OAP8iEdGkAX1mtXRLHvGXTnMtX+tvfj4Vx1oyreD3/jYNqLc1pRFdKy1vMMTBy
W3x7hwaIuyI50/89uoS8KND2s70LJD1Nk4ZxE+UES250IEVTtnZ8ZABOxAB84ZIm
XTR7QpBSUNWexfKzoKb8JBxaPFMbvbUJSyClx4et0JiSb20rp57XgyTGuBDF1+D1
s+QNqX4OoGxxXWCUhJL1tkqKOfqoLNby3evIpOy0YreWMTdHQzth8kad4ZkEj4LV
SNOQhUYSUV1YgRTlSyplcUYsUEH/s0kr41aLXBik6Kz0cn4RtU4T0uY8E3UvdnZ4
MyQLUqX5Eu7Q4wTMU23694nxk/6/8cFb5mhx3BcKSXLw9Bqe/hPfP/nbn3pM1du2
Yqdk5DLyjuULOM43bRqq9BIGb+FhZzzb9cWDxPnr9LkZ0bU+39UOByJRtljhIqzJ
vqneQndNYlK904IQokcFHAFRlhM+8XM74lPzen2h5vFdiWQTx1mIay9tuEEGdZ8H
OZ/HM9V1qVvZw5qx2L83Jq0ij0Q+/dyD0fYqhRlXh86OYjV+O7g47Tsz+QTWbsTK
5i+cNZgWHwZRWd6KLsxX/PBegS+h42lC7WJZBFX2ccyFNpndTHwGBSXGp+mL7pM6
FNiqflOnPTw2BF2E7Z9pMrwA+byf+zmxVULFYxuy6Fm3l3/kegpAkzsQYtHmbjjx
bSHVA085XUh2dOF0jJ9NX6/OkQ9uO4wUmuob+ZMQbc+jNDJNDbMy/tq7TXzR49xe
QndPEKIFq0X9Mt9tEzmP6ECV67x0Q/SDhJwW+yEZd7ksERAY+r7VEIUFEcxMV1RQ
F5hSnoLNxO25xUCvi0yKvqEQBETfSnkro5FNgb8zhnv+18/0Lmx5xwxdmopN+Kbs
5ljdo2EZroh1lTii0oUn0zlWbPdA+qx+eB1Wrl6h+QPLKUJp0NH2iF1Xj5bUJ/sD
IregZ212QZcuVMqT0GPMdtHMyDiNDpidTOuOhks1Iv2gsXvhY/tkQBQWM9gJ5RZI
/peTLGY1GWiprMuHRn5+uZGIhUpVFHu4zArNxtwM/4xJb6Z+vV7kRtKHEByqVIJ1
CAmtyTTDUKYklMC+X1+bbi8zLjXliQNknZK6msIrrlR/xKf88bMPFp2gZCPy/Xpn
pDLDTN59R9cjQnqWBEPJzyuzO66las95he9GAndcfWvuTh0Io2UJX61U2jU1WBkc
0Fo1Cp5J//k6cVcu4jOZjQDwlvP8Xr3cJ4zc/UP+hCJYuT2l8nu7uHoXerpwoCNh
mxKByIk+8tuFtD4EoXGlYXQTasqQY8uHz+CwqBFd7PISNzci2oWU/YK8Gge1EQ5O
/cU+aoT6N3QeA+ib11zo8Lcm3opolaFSZa1Kl6LVc8448rSFJBcS9IP8u5w1UFs5
GbelS+AptknQOqrMZlxV+ZP7f0wDRMqNBDf7+BRZhH9p3dbWFtuF87WQjNhJSW2T
blGIaZ08OaDJQoP0f8FVHC/ycUxsBbxpvaNKEys4iIixCuK08UJDwOyAbhuJreJ2
jmay+KTQ0X+RUT4GDhKdr1sjprz9PxHIMgv9Qhkk97xwqiCKJH4Sr5BzWwdzFDhI
F950Igri0VCzAF/D/lhZHZVA4GBUtw6S5dtFasdFJ2QXBcMX8o1B58TUhkptv4ip
vAREQ0EN4VT8F6w167tC+OUy68Q41CcfisY6LBXFgIgpELYbHc9kQd3jQB3zXbbs
T+ZbvdMMhjfhuTAyLgH0KEwcX3camPOp4mfRdOeKi9FB8nqYgPjWijTk+BN9HJWi
Nc+LD8oxo7C+FELIO+JK438sdN4d3MBLwtUbxKTsn0kihqzIsQv0w1dJ6UP0dbae
zomdhMHaxZ9MkYrTRpXAuiiflX76OKXdwmFx4F+44dIMNbhkq8Ob8uP97L3VVca7
16Lm3cZH0aR6hs22fUlMoGrFnnDTcaEx7El6MLh9HZRdZu+n7kpxooc+f273b4Ka
fpisfYScJf2oNW2i+sYyyvYfzZrTKn9HnfQrxL5qiJvvXKgZMtNwwXFg3n6saWnl
ejMwyuUYXan27Ur/G3Jrfusgf+byXcaEcbMa7uYx7HL8o7f5ijwB2Z7bCNhB5a9g
XqueX/1qxFu87jBYPGDdw43hMz9vy8qwKR/La2RQfv1L1Cz94rdWiuta0BnkR5UB
NcmHxhWRxWCa3PCs4LmYzZ4xMEydLunIvVvUIY9mQ1SPJnEzYsYDH8WOD8uEeKJ8
GmWumSnE3PY/Ban46Rik70SDojJ4zVrt+J6XcPNuQpNuG7QMjNaocSh+RleR0YYB
Z7l4EcB90yoVubX7ukEQ0Hu/rvuCjykhbmkxA0kxG/y5EZWTbyA4et+JJ3S/RV7M
tY90twPHYzhMvADA9mOx7NclXox3vQSl8MURGnFSU6n952Dgcfk6bXJB8U+aPu7J
0WfSILbAOGp64YJDY+Hzk3J3hKgCYO9Bs+OM8YZBBCleZm9tqV4KagK74wvJRdLk
O+KaGYhVeakPxI4+bH2wunY2Jy1wkfA2Av2aUfyxXDRPqquBnrO+GnxsNH3cAI+R
VnUqx7rEd0wuPWD5hhO6XBum3PxaC/KzSzuEikwoLZRh1hoIVNAXnufhr34SqdqM
M+bjMCNAiiJDf8U1VFQY03M6O93W0ONzqgyy+l7PQEdrmyvP1UN9+36dkEmz6X9h
uNJiVNpqQphKWZZGmzNucSr1+leRTiq4HQa3mw3MqYNh2uL2BcfSAy0O9Tfesuj1
oGsMA6B+ysAqSGQETcAjfHQAYgU+0pwHSSDvbGhNGy4UijICSsG9m7RvcFW3on3o
sxNctewttQYvij2YwQkUpivRF34jz/xp7J9M/Fwq27gDHyc3I+rwE4BXoClEXI6h
zpVXqH+sfkAXDJSQGWKZNhlBHjN4hySpbeEQiOy2mZHwp0x5Rt6cemyEpVAcl+0r
3/a/8wgKvn5/eMC0hK1LLk19lO/6gowOXEC2TvTLjwNrvNVDN6FmNN0Rwqenms01
w9fEg9rCmUX5dRI1/RbspDW0yhjuo8E8e25M1z78ohGOOuVUZHHfoG6bB/oPNAg+
codK5tmTSp4MzlMXL9di04g1ZSZcR0I0kT0jIwQXQbr71rzSpudO+WWeukFuxq1m
nntpaT/E5FahMZnvTGAZqZb4i+wtUH+dW/zl2bdERliwE7NjOl1oOKrRT42HGXWv
dTPpagMlrGQxQN9u9x22FBMiYyYQaX5Gx4mKTCOPE+O08/Xpr2P2CRExWmCj5jCm
0drRHgDQNWrM7CFpt7q95Ewx5ZRIud6GdsxAwY4N4nDIwBYSqhno8TiHNkbjYR0V
kFApIfu1bqx+kaGdCC87JNNvxO3dOR6QEzZsZ+uXZCKyxDcVHpcGDXZ94r6+rQyr
aKyfLxUvpwMnj36IhNQyQAzbml9bUSM0Fdy/VPKgrUylJLponNEymHhRzoS5e4kX
9dKb73PLgbSetiKbJvmOkD/sfi1NY540OuLspXSJp4A2pw3t72tXseNcNyUR/yFR
771F0JDOAUp/5a6zztIP6ntTCdfHPybF8AN+H7O1J+HJFf/OEDnS5b4y5UuWMkae
vdjC9kWOKin3dgsNBS42WBzRc5HS6k2ePXJzbba/N9BjqD3sYiwOcXo8gYUbjMJ/
FYlZRQsvOGg3SBskCi1lM1BwIqhO+Us++NIaHFUyfG6hgs3M3DTKvF5KNBWSOwMB
lE030oG5uIfFRzB+jOoo+kxiQ9aWtpTFZId8z82QA8wAG/lxfaXmc6Y+itaPoymG
v8J/OPxkULC/X/fUpWK9/Iyt0oNRnbbpeUdSSDTxkpk7owmLnUrnKkNg5skDUYoI
SVPe1CJqwiGfT09fI5GXEi4LZ7FKdAaMegyNKXOG1PTSVlsXVFGjHFILI9wKKcAV
wNYZhFU6WYJSXcsnBij41MOmh98M9uNzicV5rzzazM+JOWELmweT5ud1WfWhnXdv
XUGUH/OLVBHj6m2nKQ/2lLl4S43rB5ECunqFXaDhNHPWvWCxNsLNvc+PYzMA+RBK
+q4mwyhvY7QUGdEdIEuAjevPAUpQ2npWFXkQStElyq46rbVz847+QLO4YJoF/2FZ
iEYRkBeVRk57Qj/i0DLZ1sbS0/HfibuARXvurnMswckjSHxjdNwGsKQmNHb+hjNP
uUfy8ASmXhcHH79lPy+eSiBGNV0tUKtE4ycsNUHfzK1lO4g7OaXauy/H9iE7mrNF
bQzrF6HkfBP4N4nPnSilXgIyjkNZuK1dX9b1JYjPa6ljM3qGlIZ08v6R4HTpoPwr
iuXK+n/KS/elknFk8A3XhQp0Amutz9PerL/L3D2cYlkKlAiTs16J9poMWn99tOXr
tpq9PvdW2e2sIif/tG1UqHEh5P9yN45pnIU9l22z8Sd5yTF2rh5Cs4W2NW4LMMFC
qd1M+Qb+GuvdHxDx+O1qQzA7GVX9aIQmH6XH5GrT5Ude/WJAR1oQ20bqOtY+ZgZg
v2FEDOp4z1TCfQE6p3XGUYiWIRGpMEd5ULzHMa1wqKiaS4CAn5V8BselFBOL3pwm
B+SSsAhuN5XMvNbRRVB9mm+2zWdmhwUuoC72/oTKH5p03TJD3bSo1Lg8wjehIaJu
fRniUetRz+6IZ2sll1qOA4YdEkQfR2GT99m8h+UaQMNdtiem+YsxXceIz+E3Qr4E
77u2Pswik6CZ/TSS2rZDUfwuCvAZdOdCDT+AyKsHcKbPbN02+bHrt9C53NlwNtuH
ADCW4CleQSk4RNCZYLtk2p0Ar3pySSWHG1PNCN2p6T9xlaHQvKuX4I52U4PAQA4X
GIbgoI7VP4xVbyr14oN+D8MuW+SMbfeXpnktF365K8aw9VENYkBjXd8l1oKzYkfs
5eT63kYXzaVf/v6HAHfCXlXo+wYNMSWmvVso50mkJJwuW3KXjUwfrBn/t2QhHNRQ
CKFLJW5a/vrfrrUU+wfvp8sAZstguR8ROFnqeKs5OynmxOyEryZSDHNJEDiTN2au
nxUcGZQ7BlHGj6Z1tLxscfZRCRFYsjz/OhNXwpILX01WJCF1sKrX9VRuSHaOXouS
MclmATimZbAti06/WvLgNn+PgqbayCyBUJPPhGV8S+sWPYpulgLMoaOGxP+AsDSh
LSHCQSXlc/UbiPxgYzHcUzp66mNWuqE5B6L4qAYSZxTR1k7DamJIA21R2mRmSx+2
22NX4wYf4hDkOu+97BPCrBa1Yn5XCMd9w0UmSSlIQCwaZEq8Ko6LyJspCH9/9/vL
nO22ZIBOmv8QAElMZWtlhWrFut9AhJOItrTqeBIxJguK4TOCIKG/DdkOQF5/RAsd
fIDvD9KC9ARYLZS0OtKfaxfNvFHZNQ9Cqs9A1SBzH97mVzQnsv0cTARu6WiUKJ9l
VfChn7CBVioGhuABRUY3IT5DYifpSpZbhCMWwedqc/39rMzK6en60ssLBFmNTa//
vvrtS7vYCmJbPApjFuXsabVjkY+FU27SMZIm3DArJ5WfyxHSiVu+hxs6wv6OSrVa
fRQmETYBJ+oqeMV+r43EMjkQ3qYYitsv67QBfsWDILp4EGXwRaByFUVBeggMD1pO
/XIDnt4h002QDLqIVkJPog/twFnzUMi/fZdJR6DI/Vh/2xD74YVHPamjL33xgMLi
uT+IPbU8StdFeFGaPwe6jdpJwCbvMqEY5ScLyLIzzxnvTV4jmZhRh0AhbRa425kB
jOQsRoNZ7zeX6xBt/p8iM5AmhHW/1BL9mKy/VrmCcDQpq9aAs4D1p3wFeINA3JFJ
kKRLMzCH1PH6C8r9Kip3NIMbfJCD3fOn9cMApOnTv8LSuGUSoZqw+j1TKf7ip19H
LBhZ0BGq2csI2IwKYt/ysZct5F4mCxul7fRn8Tr6NgXzNlheNRzBRo58BVP5oGOT
/1h3Yvw04NVvirGDBopBXTfoduViLGjl0yFm0BNo48fzFVu44ZFYuhmDlBkgSIeU
z+mcybCatm/HAoYK6YNzkyT2PiTPNjNFK9uQpv+qZzaEpCTSEAH7njk5O4xdRiQ2
9DSV4LFfCNVat/EN9iQBLZp6vLwp7r3tlUu1xMx8sqlAmppGbm5u+QdY050cQBy3
EpN5Xm2AXRA9cNUtdLQDhmwEP9ZGG2QsRJA4uHXvF33CdcKAasrO8d4I3tjAYv73
T0bWZSsKAY67OrQd5XpKb+9bMEgh2hikIvGA95QdGEdleqMzIgH5czyHvlyazjmb
ygog28qSxOwjsfgD/xnVX/yLlfZVo3vDOo879b3nEVNZbobFMYLslDu4DjGnD6In
4Vj5KM+qaYWdPMsCQLB6BTqt1az5aOO5qU8vpMe4czjydd475MV9rYaVxweauxdd
Ej4WzE0Mte6i0Ff0VSoIkDhbPijmcthVr1CIyqGiib7cMjbdMZRGpd04saGDQxOF
sFMUAZW1Q5sSzebPNP7n+7hrQYscBIN226GnZQ5KFkh+Q4o3PejKTPnTBHJDFqTU
OR6bj2NeR6QS5relOtu8u3eUqwYmry9x1ZpeZjGqhitA1lEKgTrpbc8YMIWQNK1R
TWfkyWId1m2ZNQcHxMc7WEA9xkA2A0W6NAgnOXFMp/EkekBdYOWdzJJxviqo+S4w
bx8a6K5i2Sbo+xb2bymKmoujbHMXzgiw4fIv86eLktS9t5gsDXl+cFTt64EqEsjp
B/c7qrIX376kW1llI6rSqPrzMdCzRZRfwIPCcPKrK0qDRPfpvtJQR3uGTvSFz/Fe
0yAjF8bL4iy1tqyki1PPc/MLWBQjE5A+sixj2LUplMBLkZ53Qzcu6QhrHZeU3+OW
EvVeKpRXdbicS7l+yyclU36jhv9gs9GV1tclC0maYgN5aWAa3zNbMVLReRx1sUeh
SxbvbIbYiKa31BmIGDjV5jD6SQQGudCLAy7O+93jDmYYogUqbB/PWt4gHN4Zj3QD
cLhIjz9co20Y5a768poRgBrkEAwhdBrVHCTMtb+M+01gtf3ldP1RCCDl4J9kZdEM
TFFI/NusDUXb3Vnbb2VEyz9aagx7UITpqq/zrtfZORjKW+8AUIblcKVlo1YQxM4e
D4UkQr6myRtQyG5DMbKq57ADDJiCSmK9wumGCIefY5TDsVQvMQnIljGvuK5XFk25
oL6Yhsn8XuVyzow/d/OUDbeXMbOlBvi3sTfouHDouUgrvtR6m6gE82QxHEz/yAKZ
IGW9YHIt81dVhu+djxwiDJWTRyAlSiUShuZyOJVFSyAsDqIHWWLV3QIp7o2r+BWP
krGoMtbTCGlUqUd0ZLxjM7f0drukD5KFHJKKQiBb5cErQIYgqiAvm4pbpstLBhX0
qtNHSOLDVJFdNba5xg+ecuQIYCRK+7XGRKbP6L7C2Ux3B2ex/ntxipJN5hrTrOnN
GmSebNDkY7+XOM7g6qiOxBjv17ZMglXV4teLVrxK76G1JHOdOipRbo4j4YuM1S1d
dXTk2XHeAmCxgXsjOs+pX3c6XjyXY0G3UAMbPLUj2uh+WzjCkjCM2HU2yA8j7T9B
ZgUTKG7oaDGmrVFBHCAWvfO1jabLeJAy6ey+rVjDHpdVZ8oNXyuS8DrUzeAws+k7
lWfJiDKhnY7joMc3Q/0Ek+vqYF0dsM+YyKKNK5+lTWGaCZMXQUvWvXg1NoEiJvfy
yeAwWVZMqFRT1nSdYS3gQbzvlASmNnfus+EdHfbwMt1Bek5tPf1gbuQlSvIXZjoy
S7cUr+lK1xcry+yylyi8CxhwcBM4Wz6oLQU3466LIK65KF3cXH3cgk3LQ5oFTQIC
iVQ/8g8TqoQUFzc1DMVaTrl+cgBl2xh/U6ju0jxJCpz1KV13IeFMXH8KwuS27lhE
UXACFornDH2b49EFMcNL+4oJrO23rQ7xCpLYJKcvedhjHxNDE+L/1nnoRWmp2+tH
1UaVbRToRl5eOETca9yp+EkulvKzScNW7mPMNSqLo9fLu8wgm15sh2+z+3ZqgnX0
d5tBGVq/wEysQSnzcgysbTHN0EtHESOZZGz02mjU2uMDi/oKRFygWGB3PTaXHuVP
ppZDLnFLRK2veP/uLyVs2rtsqqIM+8LmuoXSKaBtmN4gmB7ZH0Z9XTooXHx1KUWT
36+Hboql9MrFCUSF6dzKAcgWc5yM7uDxGk1qadxZz/kt+BNuLUecR0rM74s6fr9c
QwWGHEB9ezSBUt3OANOMi9pa3D0zSn9ySuqCvaIWjIV8GPaQEU/fkhZWtuDKTXLR
5naJ4748QK12fa5tRACxU9cb8eiWyg+Jr9xp2bFu2KPSyZTKwv/EjB5ocXITR9/Q
zwGBAHMUJbMtaN00ivUSVI7siL5jjTj97Vc3XWSJl5ijIxL4GtMeyIRiqB6GV6u7
KWnchp+GhIojsHyRFo+CJ9CQvwJwUc8vuvHlAeVL3OJbJ93jpv5WA6HppBwdhz5T
0N0uF4A3vc+qE5woR9hm1c0SK3jaznStImE30PCH+sYb71L/VOCawMyOSJjedKua
gWhQVnkLmn0y6IglBulczUvv6FnMzDnf19OamURX12ZHFyL6opVDA4ujiWVvnVJu
QFTGo4RU6KaHftTTc+9JXbXPCa3rZiTRqpAtq7ryEix48fmTvM9fi+E0BKyVi2Fm
/l/KulXEVnEFfHrKVPJufGAreOWj92KDsNZ6uZ2+GVilKna7QW6OGmvB9Pb6/LPG
GA55GOS92C6/zpLwSNyyEdJOSE9rxyC0RWDcxb47TEF3r88ommrqNF0GwDL9/U/R
52YpQbtOzKy6yae67zgc+ccpSnnDfyVD8vyPv5k2t3HKm1CfFuZ+l+15MEVlK3nW
4hLgVuQBppBMR81iw0r17N6QxoVvFodtDe6rWvTedSkSgg6weQesqBxCPMhFxYI1
xpajTob8z0UBq31GWz/rVqX51hrPJEfawRpEWVntQZmbJ7bkpqOUBov4vKagU0Gw
+q8mK4lR2+U02NHYgXEZ9zJPnmWQenRFeN+ZKCPfw4Qe4H/3ZtfjIMB8DiJ+9fXt
zlK1TLEZjDIppazrSlmFRLcrIZzVDdqR6/vJs5fyDR7SKqzGC94+hWOIbHKRAtMZ
Mf9o91olKIaHRVaLpUHWRvFz5wn1CxN+LPZDVjkNVKL04WeaNNTxZASqIWfb9uXH
4deVh9iv8ywIFVdvE6r4pZ7uguWvCM6q82XBVFNEPyQcjyuigAlt/pbPcAPe34a8
Ie3WYjpI55HoGLAZfnhMKwZEkDyRc1AzhBuqaPucz8QZ0PeDQG4tlb2aCMj4LLA2
VAn9eRkyh1fociekMcSAq+J369wahGDXtpgSD9GvaNI9VEqGja+xWbZAkunSly9z
Y0F8jxbR7/tbhO2GT1RBtuKx8nlFQrTUjaHESakYBE7ODPBc/dcOGIp/kmKvPnme
+3T3eFvOgzvD2ACYcIFybaignSjCUo4UdmYQZNfCgO+dzch+v7GJThXbU01hLwpy
9IkkrJx7Wh1i+5nvOh/USdbLS88urnrEQH86sYP87w78hEPa1CMy1CrqQzuZzeO+
m3Gr2pbXjUqvskFDp7QB5znDhyLFjnwnl8OYXDn+cgu4nNc8tNIY9V0uD73yNVEa
/O7w4w0vghJTM9wmVUfYCT4p6vdHmZFe7vj+M+fVf37mpsCcFoqwCTbJr8bJbpO5
J/Md5HKYM4TnC1/bOa8rOcn9iGAQl8ltflFcbug8myTuYVqvKoNiSpmH8t+Li/vu
a/B1wz7cOMZ1gPYrfk6Wt5ecENDfU8IRlxHsaFmZ4DqPSq104RHaJ9RQyvBHNfs3
nBRLJSrkjHpVWXSnkV6wv7x3+jMHwEkNFIzlOwukL+A1nz18fjes8ckWOYfYrYL8
noRpgAgjBFueMahkCHELG05ZYAZ1rvGS9gV1banwK7J5+PKS7RsDoykmxAS5kiEo
/p0/Lg1Jf6W3cRxfjNPJaMJffYXpR7hxVBCyrMiIt3N0RDKP+bktDFR396z7FeFK
q4fRqtuDmpA4Av1iDQHrVSBVFQioax5yK0bzKaapqRjmLALM4o2zFPJnOX49eKpD
lnonlQahyEZFn/9S/mj+gu9KPo/5FBLFyXtmm3ADrTWwFKKau8morO4MSu1rOkzy
Jswe0RY8ZlOVMhk9RJ2/PT1Nmtab7nwHAWeD/0mpHE3585US3TQt31VTsbNPOSEj
kJBUHfm6i03aKXzTAsMBzdQpE4uoX8xM5TO9i1HL9L8ZewZSm1SgKopgv/UNHIrl
9UupkH3S6XJ1VgpkFnFElpeYl4MjvipLgIgdjQoBKgvXb8LW7s8TdbVnvNsZ0aOs
GIiB2a6rOempnOCkH81oVhRkSspgNWNjvR4jUQ5UPf8EdYAJI0c4SwwA8AgbFT0H
mndWnDhg/BgMI0uWAl6HMwa/zHv7jD8EQ8UGSYSlDisIPPOMUTLppgztn10O2QbJ
SqukqOe7hBLCB32KHS7osGUJ4gP7HrwZcuaDKsiNsgCyu+2OkAF0I8odS/CR760D
y7E0UTnrE9oK2sIcZcT1Maql5aenD7RQixb8zEQDt+tpbpmxb2mdkRiViujNheCH
XWMBZRckgigdc8sv6IUCDIKMRljGPtdmIqhCcZ5e3n0cP/SdYlZlNffDUQj9wFGT
5mB57x0nuZTDF7Xr1PWmOlCz6ui81sgtok+wBEaTuitkEEHDKJz6Jj+qP2O5o4i4
lDowkQdhKKTDhInLW1CdwVark4FD9nmGcIc6ldsVRqxOUAMwlbIm+Rn9JmLAIHLI
REkDRAZ9b0NZK33dJq46xVv/m7U92UhtJ1yWbx+QIEmRGbM7u4klDhxzqajunf1N
iMR70BF2qamdZRpkyABAKwALLavokJpXDOFdco9Ijwc2qxxPNfw38mzA6I/Bm3ZC
6mVtShYLSQ/Xsdpj5GhtwFvV9iUAEdUCWikTxhPfBTT6pYAan6nbtPox0fPYBfox
1m8OGpz481SUG2Sq/gCFwT6AOWISDh+hWqYvnnuQas/p+fQTI2LaECeiUQIO9iR7
LkOZqIwkhCh4NaST+ZrZnE8C/2q9pG/NMxvQluut+hn3dhhdYGvrwXROmbhUiaDZ
2W2HQ9dEPs2wRp3w6EvRDX3/yahw9x6idvQ3DPSjz8zRqjN4GHZLZ7LtkkWWFzPZ
eoWxIw2VTdlrOMPYLeGz4jUWHMwxevfKrnyKOB/TeaLrPGhcySIcmuT582pQdrvA
PmN0wQ2P8xXxfLkYo17DSn3B0SrIwbcC3UG5xPXhHU0bPKWgQk1Ab/Ak6yIUPKQT
ugxmosjYecVTcRHZBl6momrT5QwK3OqSDWCr9LFzO0zanNOehacU7T3FBBBwY7eT
Y6cCSmf5P5Iug1GOeq1pyURsG2qTJGLQTxHHZSEbwhVXSp9txsuIa1YnH5pvNRkq
bDY1MCimd3KTHYqZox05G3SFtJXjknY4f8CEO++ro+AedqIahNWadYTM5ECv7sHN
Nxjq0mzb82tu2LS7Xi62HpJPftLzag/WJohaeCX537BEnPPVU14Uo/JxF5Ny7kK5
+myKhqucPucH+5ngdVcUuBTHWNtUjw07XZw036rZNCI/iK2zJPHGWcW/65TU09zJ
/JqzoSJV+82J2zXT29CCy9GPZjK1CPkq06gouRw4H7GJPE6rj7zU2iiTnLXmqUV/
ot4kkdTOuO/sn0P8N9VtG8ATtN+7CzrY75x9XkCwFEhhAfTZ2cdM96SCbN9qVM4/
3DcBjgdAc+4zzxeNLBkAm6Di1ZdboHSRgg0NJ2MYGMWxs0i9ZL9zC6Mr4sDw9eLU
BjCS6HZgiyEcExrPY45cgTwebKrdc6IWGpE9s0AfzswB8AY99wvD6a0gFtsF/egX
je9/Dl3CYsA/Bib4vH480eQaqVTjWAL9FTnfHuSAWFxCrTzqW+AgfH00iCpSIpvX
rZUjCY62iTNIZirvw9+AX7EZznNdV7c9tF676QPlqZRfbbvNsHg3rlZc0TzVQ44/
1Q4HJ/JV+q50Om/sEioNFfG0iDDY+6PEoEjtDi+3VeHTtdtaHwoYkowV7Fc3zTQy
cFhjwEmVHlJevtIN85VmIFw5yg2wRDrBjb8GnXpGLQfI8YLGfVVfRhAd9bTEMO4g
kU6MscwccFvCA3rMtcxhtViOA618Co4ZF6ApwVkHLHOY64sSupe519QWSWL7xH5V
XjXKMawvEfkcvoYzm2rfGyfq5mVYfZTaMQ3O8zsiUligN+3xb4+UfF7s4P68WZ1f
xjHf4Lw+eF5T+ao1OplJVbDc+9evrbuNYrygigSYNxpbE6tv8EsgWgJCatn97UQE
EaUfJo9c67QlInF5Nc//i0XPEnWQcYULAyFR+um00ZdeJHghlkwErcFCg/GpSmJJ
UYttIey9bsyO9lT9fxLqarubkspOZ37JMau0S8rtjw6SkRluYajkJu+sE4Sbgydc
t6icHTS8483++KJd/alJ8o5OSCcHNvyiW+R3AQa4FIfcjyXNvTRwtjVgVO/rkLvI
wzd3y16XTyrRAC8V5oHQ/qc7Yvpz2cn0w8MiBKiE7qY5Bkqt6yj8Lm1e78QarKq/
C+tjjVYk0SbrE3qvj31RZ9Dr18bqGh0B/BiuKaXCzSa11851NNA+O0ZjOCRkQNLj
rIV7pnJy9i+nVXddiaf35CX7IlMlQ1zY1vNmwp/SaGCAgpyMAjs7Tr44LHZqKiit
knFypM6es0iRf4XeuH5WNFOgvBEkKg2tWZ7Uz35VCMBf59Jpe5VCEm0hZS5VTXZI
uuMIjOQhjbtr1t0gKQBPNggn3YhLTi4VxfJR9twqly+U5ks4ztCnY+J8W8g/6E2C
Jv9mUcE/cjh/JO8Xkdn+86/McaXJexUKdn6/JIz68TFrODaPrbUc8dMXKfzC1x4z
RPcoewVbhWNlFc6hkwpMWp05ZBpuyzFObHQ+ff07Udg3V2rzHX/6CfPY73UWBv7P
dinUFtpqJ036iUkfrifbezF/i8y8NSs+53IzgGvh7kV+7VB6NbL9PSQXM18jI1GV
mo/5xoMLTwECin+yrqVUIQWJx6Uy+auftJdGxSZLp/Vso3iQGVg0+uUKnn8vwrig
VgKnHk1ywYQjI0WEZYppOl76SKZTtXrTBGS38hTwmRGKGxNTIgTcEdZVDW5xAAgg
r8mUJCwhpY6Sbt0wQ261zDsGoCdfneKH5aYm65gv9TxZO0PEIn2vWe18v1R5ApII
kuDy/T/+ymQ/M0VbiRG9WUNqAa/3zzCedJsSl0ZQTGTEb7GGCz9FWekUfcCqFMsN
LqVqfbwhW9dw9oZfO2bundJY6JxpR7nd5IOCGQw9jhdbgpmxzemHvrnqEvkOYK1d
deDnXs8PCGA17m+CLySeTPVWKJ2qqZvao3XMgqzxQP5UGvcbmLUxgfB6+mTeuPm1
FlCJkBugkgz/cWeXxe4vGo3yFlHFHg5UUCC4YLZeN5UgLAHylLxNetxBAtOAKl8L
fXHbHe1KlFNPe6g9v1Jsw6CGCpf01tUKe7bOjK3ho0hLW6p34tTRkPL7BW0vJ3J6
AVAYo+qFlAwApHsqNCXflLzWt2EYdcjAQtTdy5CeDsmDAHGea9O7VaJtHWlXR3bM
YbV9tZNLb5R7HxABxsRiTM50ZPkpTsr5sjovEpD88JJyVUEO5gDL1eCJFgGyWrx4
mOC2l6U43ePEVn4gNb488CJW2euxJSTAKqgE6P1YAnvabVSsZ053Gp23r99lwThg
1PCVy+g1HNx1vROYzpvoQjCquXm9UiIlkOei8Bgz+5aD0qw1Igw1Pyd6y8TgNfEk
nc4zOpxpa0wCnUfwut+ZHCjtSoOw9JrZkMElW6RtAFM6r7pKe6rmdWssmr6ZdRmt
c/+nyeqh3A96QXNO4phgsgdg+tDPU9kRKo3PT2YiVIEqA3udrveBZLYkstxEijXq
nxeL1c1Stpo2wUF6EZMAQzInx1FDJ5hy4YFfwNSKGJt9qY5FaIL89e+LKRy45hnP
/FxQvWBhOhio3RrScrYKaNU+2/ocOi0WRTrMvSupdoPKKw5C/JVod+5NFkuKSYEV
aVqyb19dy3sFrUv+MzazD8AJznqWZj+6Cr0fVDyGoAMEbjB0GsaV0dTbab3Tm4Z1
cWDpBj6tEqEtr9zUTTd0QekMUppaHDB3qLfUwvzLlm2rp/UFqscojuN1k0t7VREc
+LfXJKWoLzGUItSPq/y5wZIhG3n3ivBWDwiXhXcgMq2UAW4elmQTslFy7Ny25aS1
Ywv61/a3H7MxX4GM2xQGzCjTnsZfDwRSkdkoWm+6QFPT+VfvaDK7WwfF/+JP1C1+
SNSKpKdltiWKgXggSWKPUk8ptt4LJJBXszelVL6TKP2uo+3Ie5YrnRkTif5E6sAg
5WHkkbrgp0IqwcGIYfJErdlev/TbaoU3zrIXR+6FOxJ83iPKcZVq9KaNfQTsBOx8
5sRilyAATndqNJPHqTnNarfzcTO7ZPiHWzSUvNLJgXX2N2g3H9ltKRj6uhfv4O63
Lc2kUZmj7AkEonCc75fxlI0rGXLVfFEPsdLCe6HCXZ3HIPtsr9mWMMduyWBjDC7Z
JGch6FMCxQYyG/Ob/yw+fQ67ttZtz7fb45H5b8aTMbTh18nIQVZQNmat0ScLJWnY
yxhNxDFkKYIuEh7tZckvKpKsVReXdFeo8sgyJYurrQb4fIhhji98CCyx/+N9Pp2A
V8CyzPrHWjDtyVSqh/SUALlzagmJEDfJwT/xBTBa+KjeplnXxLS/zUYh4DQShjoJ
TqF3Kp7YyhEJ+LzTVyRu7Y49hTTddR3Cu94f9YwYGTKBbrtUw6mkBFwprYuKi11p
s1pl6q1JVpT0vEEc74HO4TraermMBXLJ2TZ0mIWS2NsDoJHgXw4SjX/5cx1xV0fm
t1FdfZjGc2EEkJw7r7e9r3om5afDS9I8463ydepXmRvDYQhJPNE4/kHlmnsRx308
mw25BfxgEAAH6TYiV7pzqvrN7Slp8wFtCLw9biaDeBjRuw2ISYuUTVfC1DTeZuUH
QphnnWA0nag8OCHfoabkbPC29yIubcpl76wop5okn4BS6+GEEJxRbBJnYdRXjId8
UeTq4XDgysZWRn2t/3hpupDAiNP5PDsmS4K8RGHAXgPbvfyaHmcf8mACRd3V3R6y
LyWqU9kB4srPILQByB1WlgmbQBb7lae0DwIF0Nx1J1Qr17Xcj0Z4vsH7Q5W1ymRB
66Gll7c//W9jYLciGK96piQN6qCZPMiaNXuaNd+Ben05y01LzsQ0Qn/KuaQAuuPy
t5hR538Z595Y/7ghTRvHIGg+/ypLJ79r1MeoSbl5UnFiX4bWHXRV85TkpgMGM7Ye
d8/aZNMQ9BdwgfBd48YMI44Lc9OioC5za4GzbyKzNAMxl9y9L/BO+fslXuxOqpAT
Jr3qHxF+9npZs3ZhaBYowrFB4IzvNu3YkY2zHCxJx5LJaqLqvGpdLPYxXJN3I5Oe
+T7xiVG+rYH+ypLSYHm34s14dk61MDrI+8v7Bx31UNMdPutgUPqE9jhL2pEpbVWE
UuE/UXodOotwgy4wpmMcJfPwX/rSwNWoGQT6fMcu7EEIJqaxbtpGfzi9lvJyd7bl
53p40K5gP3MxjYlYGqiaSkmkMRgh7+IUA/oTAxTmQJ32zgo1rHx8NC4sx9PgYGQ2
mME3Ygx7ux1uktCFAGXAJ5sJ1DEYRfGyGrjmle/37P5rk2/3gD9cNsniQuhjHe1x
gkOnjX8tuq33j+oq3SebyUaZMPF0kfx0DLJ/NDowW2fEPdOjFtJfIvNX12fphbQC
B0qMFwblcMEYuy1P0XKfusaDCtjjZjyCaW7x4BEks6yt++nhXjINjKPro+/malIf
MOaUhUfbpFYPIVefNUS/tnMY1NNcFgG/StRAuTSNmP9ggTXHzskSBbjHePZrKuci
EgtefWvkEfae0XK2uXOB1WvZaDCHrKWOdIfi7HHNIhXenVvlZATkEpT8MW9W3XmM
JYqQK6cVyBcqmendXs+HyH4Z/iVSLb9zBARgjtFDtafhqeoD3QHYd7aQFR26ncfS
yRz3seGcfE1jp72jJ51hvJdV6Spl3pAHwHDhByOuPs3zpmI9pfEjKRwPJAmP2zFP
KPj2H1/ftVpsf63aIfP1G0skqJCBKaKVEp+5ILiZeymqWw9zElNHbZnCxOJfGwGw
WO7MbKjIHJh1yvVZnlastgUOraTTTz5gscjUtf8ph2H+Q7R8XMa42J7oCPL8w8hg
WtwV+ztkambqmXmMshOnvJ10CDPMOi1UE6KuQnouUNI+cPsfOQAqB/MHk4OYd8zY
wSfhUDsY9rKUS6JRx88lt3enUh4kM4ORYkJ0TTxFAUYWAHMpEpq3w0fe6d8Xaotb
jY1YT1JQOerRRpZrlG2+aEjZRicTvcineTtpbCPuhA4rniu+U+9K6E5dQrT16+Hi
E3o9wm0n4B3/Uxy1V7sqS4d3YSY395A00AHEqKXlnVg54k0QGiCX0DhFF1Pp0uFF
V06sIAfQcPboC3OCmFGlPRQaZt03mzYxUB58+FmRZpo5XPp8Hsd+VKntGJsE8ppN
RSw9vyxmtF4cNBeDL8q+JpRhx/ZrQ8MCrYQHTwFkH+48Zk7RPFedP1qydlx1KThN
MKqeHd2iYDrKIXOE2HMcv6l3J1BELIbmFA9NuHJPW8xmAkOt5H1OnsuUV2vTlmXb
kAfeEdbUqjNSTXr7SlldkcBCJPSgWgQJMZPCK9RRo/4cvwLv+IMaGUe+NMDVYXoP
oR1Sv7kLh6eNGhU64GBrJ5xysnFxEw9EuJUWginFF1uWNHWSa2Bkh/gZzCFvrgoV
tjzlkWkfQ6iAJI+O/eL/l6PpWciihr14LDPxdZO2z3eWkxRJ3KhMJhRrhpsCcI2z
BrMWyS/0rIjcnS3SDQSdPeE425bF75I5J9jEBlGXSRI0zxq7NrGIv6k6+9PQfajx
VBfxdXBSjMDa8PyCcwIohmHHwiLJT/gv+Hl674a0wQOkF/WcO3Vi48WnN4DEnKLi
VteadrTGvf9R22jHhnpF3lAA3SlY4E3S9AvB357XQ+qoQJ3+aE6NaW84gWUROWvI
gVLDC5/ZJ84b6rMlWkYtniPbFbD9t+DVAHfynf/LVkQadYHOc5fZ0ICzUVMOCVXP
g8caZugVOLFf0JEpUl/9U9lxYsb2OWR59JAaWv7oanGP8pFZ9M6B0ICmhTsAcN24
nZwaGFCSuoiwE3rcjIBhq7CkylcrCoh7RzERlO2CUS2LDaaj+kaYkAL7oqCcPq2H
7Nh80aZoNe2V4WXAbTysG6crLg8ihXVnU915HTBDylW7Ho6oCHSuYykR+ecOfIkh
d6S+Ue8IdJC/HJyq32oQxtlEYrj2bTCEH0YF1i35lxdvio8SNODHzCrR1ej8plBM
9g6/c/pc0rGLOI4FyTNwf/8tkCsZr8pVMparMoeFuyFvmemJitbuvuJqzWfcLbO6
7gcIt8YJQJvYOANKlEfaAJYk/Q0sr8UdYrp1ZCczDtgg7eJcCGtJZareGSqjKAuS
b9/ucJ+thwfCs72Fr0A+EH1e3+fm7audhkRmpO5oEjwYBueLq8wfybwFFT58/UUl
GOi4TON9uYvQBF+GTHVnkfnA6A0tNJyycUMKMoSRzeA5DIfN6pwWxQCS74M0Vgwk
sqUHIeCy5SyVZ17ZoGJ9k2si6cD+XIENlD1HpEYd4cdNDPHjXFt5Z/MG0fVYfR76
G2Obia3yGpeRjXdFPy46JbD7zLVmwW12XkLtsvyN0i4SvQyKuclXX+gQB3ZGQzAs
Lzu2dFnesSf5CK9MYkR2Gs8QZPpySAys4BStHNdawLsYqJWneywYED/0zL0fYYT0
+MCIafB56z4IQiUB+OaXHzw9rBs8UjVG72XTW3DLMMhbGh31C5pnWysjWX4FecxZ
RsG8OxE+B/i+1S7IdipHGpLnjEEEgjk49bmOnlogMZHQAlNpEW//5NemRWfEpgNg
M4PMgmk6/9VIfXNuxGy4acnGb3SqBgJvTDefk6G+irJOlJY4vDRgjK0cFKk3ryYB
66H2JXZWIhuc8Lm8ED7gv/0KE3OZEsS03aw6xG9RbdGeFZBHmCVF8RuhW7izitw4
6mrTMbURxOObdx++IHoh0UPoYNa6ieKcvTuMA/bQ2CfrHWoKIR5G9RQOS87Tjqdy
isCUhQP8ifF8hsSMMbaVaYSsRv+RQxz+9FRZdMC7drkysunP8DMZ60xPtNRGQ2Zb
Wk+n82EVWRYDVxi+86upUcxOvtpwYBoeDuP9TdwddX93uI64xtRgt+4zkufIwaaB
q40FrF+YiCDNVPQvkXKIqZKJbaDl9VGUMJIi1AZOY+/GtyVliFJHqWEtVpXCsFwE
OwSp+ERdYJOTdJcZN+OOv1XD0mzSuZ4mh/KR11EGcPN+ZOrsNaLrvIk1PpO15V29
BDyLtiqy6dN5xYts5plGLpi0oJM6+GIdF2BAGyh8JDUbz2GLY0oXhl+nlTpRD9C7
jPTV1QklL0DCs5iIPbPnbkM5yNWbyTCxRBPO6hFfDFgkH+v1UxpqdYzqu0ws19Gc
ru8QdEO1Vpijv6ByYNyV/TPVuMsbvj1zy2KvWwCWx7rtIoUjKU9DCUCXD0NKW0oe
syf+109abyUay8LVqiFst55padV19K1SQxLpOib6waLUvqBqOmBYLc0x8VWjP2ip
acQdWuL2M7X2ytM4BdUTeAgr7mnBnUvHAM0qn+qMaFMp7gRzmy5E1P+lIqLd2fhu
y0utQh3tUhmMICaRrjZmL3BdnXfTH5vHJUxRd9ZlaGVGsVc1ygVvFr3uqe2LkAzU
WZX/JgXg7vz7W1ovPLDTzLAIrnw4kF+xuVn2bJvJNQ2W53UFVkcckDAA0Vwp405B
B2ij2o+dDE8VJPusQ/uC+8Km8knTmVMlqHMiHJttzwf5f0wFOIxbSmnSS/81vv22
TVwpap5yr2dUFsk18F3sm3a7Jzzm6PsLG3gLDSMkBySXa8V1EKWe6oQVl3KxWz86
ALStWsf8DRvmrN/8H505OrSvlOOlSRJUfN2NUgfoksFWHK4GiwYDtrYAJrDIKqsk
xO1zvAyp0APCGicNLH3BXFrVoElkwhIYoTiQWbAPez6kpladOU2/nhsWQXi1sR47
toskCZQEkTabCvZ6Wsb3Q8j4bXkNGzo0hFCSPj3QNaLR33vQoQgljhe/d6ID+cMr
oGjLbKjiVNBM9iMvR0EUNPMw53WeQA3Z3dTzhB1v2VD9/gdIusOR6+3euTD+q1Ee
a5tkVZv/peptDKBh52KYKjDo4Ob02qpYDlsQJCar8u8z+hlv31cEvxM1WSYZNv+b
LNms3sBpQw2bCY1y6x/DDokRNJ7GytetbYya+pz4vKK3Dp2KnRLmZft3XsvpHb1p
5JTt4y4verneWFc1h+a7YMARphSoJPLH/yIYaAxlep+sT9tTZJOEbDwiVqR/H2ud
5PuT3p2GkUkP1M4U2bAShkguY1eFEPJ8i97svmSvBqByrPiBTzQMfBmd9ASdtN26
tKtVFdlTa25/CjkUQW7UDBNnr9fmYRWlt0nwpciEHp8AAuTYM7BxmSeq2bY5wedp
yhTOiULAHLc+tvXwbmOFflx+oRrb4moYWAEa6llNvNhqmqPSgMwMGJfDMQ81MJE/
njxhWOEO/x+QJmIVqveYP+59R8ND7Mij3ZiZHc5SWYh/9A9jUvhFaLiXoMSK95ut
BUCGo3/i+A3UohehEpeRVUMmnoPSoICQ9vYbvvUWqQepZOwel5zVlFn3ew/ZKRPH
LnsoOEUZpH+qOj3/k7CrMG5+QKALcASI8Ynt4I/vS2fm7OulVSazYFD66+ASfyo0
FCNzc1rXzi8job23dZMpprc3cLgERTJ7gqlGE0xamDZ6G9eHtvVQw9bNN3Z4os7f
s6wd7f7UaHugwHK+HhfDqKFkRZUQ1g/gTwexWLrkV9wIYd1/AiZJNKcD9HK4stlP
5/OoGU2Yp1ovKQK7TOt5h4HeI3YLRt9RFdLCM8bNBKF1sW2vJXCEw99QVqRk7Hwk
KHup6MnyBtZvY+vi0OrEHbrWENtOg/W/DJZaCiHLLfB3pULOza/GyXVZerJvP/P6
Sl8+JKg3b+gpHT2Hk7T9of4mgZ0mJO2aoNZwOL1L1jZ3NCIez+XmYLZmLbh2Owst
WUB8P0HDOPctx52yCMlGr9cAKQY4GThSIZDFmKZoVv+lZAL541EOsfH4NA4VGCPS
Gx+xB20V33w9QjpLAijT8aBpQWafoLd1Pdl87iZmbCN6UdVu83xXNoH8tnuo+9eC
lE+MD92UWmi2G3nadDjWDFsl0cHOhx2+eqMrg7DpOt+BdwW4W/07QTVCJ3rsz+KW
CPA9D3ZV/qMJuKQ12HX80gbNjaHEaKhsuoMR5qaPQmb3IwyORbJsAckTszyI+Auu
41ePelCUrKdg8Jj9/YK3oo2muMLiNtN7/X3aeyRs2sxtvh5J+F7JpMsDIZOCW6Jq
z4d2pA82TI9nFeS9OqUfoBqh66EE5zwhvxapzoAO2yY7zVhwmpHVHq5B08cqBL/4
q9NGBZPY/U0mwsRqKVEOdPDSbrGlR1uJhM0ByxYHHhS7u+Pefj4TyOn6HFGnTdHR
59HIrbSUIMqlRbBbwcG+BuOHUN/MGQMKXAGmcO/+lUxt7ETRMQCPBhMeshwHXykW
n+c899RJR+d3uuclUmQXqhzbcgmuJBur4ZH1jqCYqtjOBAr6NlpPp4Qa7BE5pS4X
ywZvuU1XsTGs2xkYZVw5qPgO2j6rF12RPRMWDTHvbqmESUipKEUbGYZK2wUe/oIm
JbEUOatoy9LRUETEQL+e2V1jckfm1cbRrBYULGC8Fm9JxXJabceIvz6EXproIWfM
IOo4V56R4X1N6J9BQfnHTFUCI/KJxPKWAHWQOtvcMENj16YH6H5tFgMu4vQRfMqd
flrbaEEvarT/QGkUAQivpstyv+949/d4N1hZFAqCYqOy2mD/1Vs5ntpbl26Vli2J
2PDyk6Cv5tnpWdC3mNDfdxHcN5UyLxwKPkuPlDiyyTBPSfIfgVotCeIbb3NKLSiV
ghizuFRFkXcfuD1GF/apOHkOUM7WF0rRPeCoDlKR7/TH9JHhogvImWPb4IGIl0+/
IHtbx4+J4Ak+5Zn8lOBiGjmxRxsVmEk4X8uXQTIEeKRy+d1xottuNqAgvxPMmvye
V3dkXo6ru2FK7w3OeEJtpxyGloha32tSto6245RA+FIJkePCRUTtz/IYhWvavrjB
ASapl7sggFyWgOijMEMpZ/48j7h0naBx7BOYlfXScYrVnO8UZb2YWd4fq2J6X7tU
jsC30Pwt2az+nlCaDQDre0BBHBlDE5SDau6RWhI1C8mtapiS5s/NcIslQqPgZ6fP
qnWv/RmDm/kBoP5rwIOV8gbPmFKW7i+nKGaaSbvPFkW4dsLO8TPi+CPjgQW7M8WY
naasrEcDzEhLCd0UmY97vk9tvTnFHE5tO2TAAOAkpVx0EdRrOU83AvHu2u/6A1/5
Ylcf+1Jv72RbcrFl/G/oMhuPdD9aAeL+e68Ffnv1Hg4VE8NBw8pq7GcbXdgCAwDu
MbQQIKHiKLL7S6lGg3eZjh/ayjgPPV5Wiy7K+Kl8AX1BRScphmHPBiuNF+AFkGQG
cuYMBxeh9kFQR6rUU6DsRwLhCXHZmJOdoOXlTwf88OGcCRTtSlWTngw3i26qirQQ
PhfZJmGdsTIYGfRSZ7hrsGA5Lv6LQ38IXpkCNYP2y6FU38dJ/snmweP5A/ki5D7f
zNV05kIt3Zvn+nk4W9bTZk/4MNQH5E2cAD0WUgkZ8lYk953YZjRF/kEpuaYePB+1
IZX4J6voqhTBA6DHVyTHvx0ToWkeNyJNimjp1UF40qtY3UteZa+TJAk8l8aJYN+1
JJheSWPEaBcMLyWd8QrLvGlTIU2OivaxLLIgDHI3/V1sMnL+jWkjV2MxyhKIVZDW
fuBN9UMiGOc/OsVH6qlETUepv/gnzLTLEV4NJTp5GIKJxxPLdbTeb115xo6KzC1t
Ad0PXiBZWOmYeFFCw36uiUnDsZBId1ENeoZceoEQh8Q7LKn9bxLpqrT2utVnyZh9
HPguaHZAhqY2ivhzmal3GhyFQdXO+zfHkxpfdeHkrm6KdIZQsq2cY8WjYOAlI/oP
C33MHsRJsQOUC1wXZizrT1AHh8JusBneIdBiqRmpK2RQxeePvMzygLCxkFA2fIvi
zH5UMLqtB7iea+vbImkP2+h8A3A1Nityfi6NXP7P6mQlQcAmpbx/ktMs0y/O1NJL
SOq/BVUuZGLH6G7UiZuafY/nQng3jwO+7FrWbTlBOigW2M007lNGY5eALCqkULom
y66K5yEwkLV+cVVMZpB05XTbWuOOGRGJsH64f1KwQEg84CXU6OaqtDAnkNsM5u/7
2xRj2dSRJKmro7tsER90Z+TWnqvDAX1QyRmhwwOJUV4k/wi4USTgbnUxZqdcKA9X
FxDHHA59tNXwkGNt43NdOFCG2rPl33jy71BdUhTIouPAFIDThF+YzRASFoUs0sAE
mA2555rvWjhge0mESEi2u2mTM9EElXQqnnjhqD1T8fWXSp2loHbxAZNNcJhnfwo1
V/i3k3Nuauq3inZjkAvNYYkDqJtG3OrzHAcnuC90NfmgIOhdpdzF7rzNdMphRkzd
DDDJy/5l1zHej3QVJawJkJr4HzGEPJxL/73H6jWKUgoTE3sIIlSmjAOl9rCJz1oq
LJj7PuEtZgSNkhE4vPe7WcKqPKS2iI0EgFg2iae1X1VuqkRmvsHTPScDqPWazrs0
kt7Tyu6Mnd9yoN8m51Kck70LvFs5j7DGsBJVsi2wPA9G9wrP2As6OJvxWhKu6X8e
F6uTtjkG0PwYiArbyctRGC1w/cAzY+bXCcMImtOSZ6tF6a+R6WEBTsXtMw5eGNRz
UXUoqsFoXYwZhh83gNSLWVk/wiKrI1eWI7Jd4ckWn+NyeN55JyF6Z/beFU44kJYL
CNnCLBNEaUN9qoD2dtohVVQq2cvig25ngFn1IiQG0v7Ur+7cHlUDY7GwdBazjMnE
y0YksHoQbbIapmIrJvqGfj0vgLhE0HvvfHr5b/a2s71Bt7P96L1LiZKsqAV+Xal4
jtonDMkDiSCXX7vCJ1mVvhFn/M7NSHRnPpMaCu2kbrLrJyWqcFNMXf0aE27TBHkS
AO9L3gmQdqk5w4QTPhSf9QmdEUC0L363YHBn9zl5hVxFOAI0Mj2Zv1cckG5YZ+rS
08SKoWS6lyyzrg2L0i19/9+BnQIyoBZEdjAn0aQ+4DoIEkJzaAAYOIt6u+wjRy9P
uRYsEEzJb/RCkqSKBhUoh56Ookr2cEk/aj7HapXYbICI42xK7pepsidkt9jnZjWw
X1qwYhGjG9Z806o/Kr2g0eUOlutTaXiu/oq44OjiFxkQ9hhGnv4F8IVuHG2LGHSh
GDNQ6qVUKcghwnxC/xncUJVFod/AnboKh+5J71kkyNXOwpkLHcn4fyJv+1zlOPZd
pu2529vMNCSH4CzPX9MCscM+5dOokI6Jj6UeThWGQUJ1CntRLlffyoJ5CJOLv+Su
S7BflTd5yJEuWqnf8RysooPA32tGA3oqQPqLDtjVqRv2dfy8dUNiJq6i7UpyP7GK
ZcuOa5sQTyVOmFHfjrlQYP2giBIBQKKiL46FVGwBiB+T5yj73cFRdkJKSIDmN2vI
tc7U9w6iMmBMn8xLq0raVjUj7GolOFX0r6YllqcuROSZ1P/1H0bo+AL5PTIleq2c
gGoqo8lHKg5oXOmZaApQbPXSuAv4mFeCNrWEIazvSbT5OeKpbvSK03lE2BoiSGm2
DfUIQjCnlGwVgZ52y31MMKXen6Q6b0OtgdEm0quqbnWtVT5ogC17NEKude9E3MSd
6HD9SHL/e1DqS7tAA0Gm8HIMJAp7CHcARmWa8YpiuS3QLQxF1bUXvkmAvwpqNitX
tAJPkXE1lFKr38yTb0hPAvljfI96QhloI0bgwLEsLHstb9iht19NcTnqu5u8RKJ0
Kcv5aAhSpUmrZp5QqRP4BxWK6UbtgC4rbq6LwcZZC7PVIwFAanFpyahyLe9QIWwA
hVPvrRGhVgOYsG8ifF09thSd6q1FlQCCKs/mooTG449xXCX9eSQbs4XgGxaxnnag
jIyFitopV/U7iK97nvV76Epk58ii7oBlADSaxtNhxZ84aRs+Rv4pJ384s7J3r4CF
kvqlUaL9jO2n5vNbb7Itaf5VNpRf7TnmRZertBshsMJrwylnq7EY/C7YYaSTjMR5
gZghfNsjr2NTt0ZzDLEfdvOfmNYzmzzvC8zpIZc4OzYt8JqKlVWeziEE7FoTudYp
JdkjlPXhKPpyx28+ttMlGB9nb/6nLMfoNiG4iOn9O+1sidc4MyjR6GGZDs4uqjo9
2XPYlDy9qWtBhreoZMqgge0ZtTWfdIdP9GY7SbD1RMe+loOb/t1qloaXd8PCUeOY
GbQk4x5GEC0d8+H1JO4BhLGZulvlsAYjCcUVbhgrzV+ll42yYV1OpIDUveJW5AJ7
FfLDdU6VPntVaeuO92GDjyVYdHR0pAlfJib9NUmhTC0Fd8+T3rXK7kG2/rIc4F7j
vj5hMovu/8oGqq1GXGP3hcX1shCwLeo4aCnmtw7Tdc0CWsnfmMmZDT0G370aXyK0
mlLrhCEFCSL0U93C+RAhqhGnTF9IQCvMIPWZtDWsqJpFXIABzdKi6W0/eIpuoKLQ
aZdMZ4Fl1aA2Ym1sQjVlw/51SQRUVRBnlGw8ObjUg8d3gmajLL/rt4ioKM7zOnTF
uLSD91+GQNyjroUwtmJHjI7qhYLCfwSrXlUZSDWSbETKcIPxyqpcgNXHgn+EwzN+
OsofD1Hk1UIDtWRql4SyYYjBDew2b75KG2w+JEoZFV7X1crruBq0cGlCSbVl/c72
2lv6hMqGaT340M5L3gkbHBNT2z3ysce2Ix7jvvjkrxYDzLltx4+syyA52RWxytII
rvVI+2cZBCSQBhFbR83EZgf/9B5Vq6dZlB4lAk+/FNqlZ5dd82zC4sQBisrCo3bZ
/guK2n49gDH6jk+rXQymqzQGjOH6mGmuoH2fydov0EF/oB2rvkuPVDKwtsobS5EN
ib6RiRu9F+XP2G4IaNIofCfPkJq5BL+AQLEdw2nv2a/ILt+ew3u4+WqWjxC+Fe2f
rjSQM+ee6qo7Tcq6ZbBUmoVC3/OpLyBNJRoWw7yeNbFh+vVQmGckVF5qnBfTxliN
q0jXChTVl82KWad5CAe3Z4NFdDDyuEtNGQSS6tEN/W3Dx658s+ksLx2NepDSA3Fy
t3fZqUAi9/3Y0W+j4n/yToJSVo/VIKQD/C9kDcNNmBiItk0ZJ3xioX6E15P9H9X7
5TGyvXB1MJ8nsLoeD+2N0FMx3K5HXEMGG/rTyk3DCwoNSoKwX6XCijmfyI/4tkwV

--pragma protect end_data_block
--pragma protect digest_block
dg2njEuRVNcoEuj1K/YpdGWHx6E=
--pragma protect end_digest_block
--pragma protect end_protected
