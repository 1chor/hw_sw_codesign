-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
RpShDOB/PiZu0pssreU7qS8I91xpcRbscYA87w7l9Kt722SFkpUSd3mwecutBJ1m
bS+ud4Id6o45cv8ja9rw/zFXg71uLstd5NJUmv/9EM+u+sbVjEL9byQ5odLzUTn7
ZQV1WeuZSidmtJpfBhvMePH9KDCpK7aTJqmXbJmxBkcSRs/K2fF/Xg==
--pragma protect end_key_block
--pragma protect digest_block
Waq/AlImeFGlhZfr75l0waCf1dU=
--pragma protect end_digest_block
--pragma protect data_block
nmUd4VrfvHjBE+4spk9itOmIi9Jq7LVIaL7Wv1VhHRB0zYts6uu811w5Wu0luatX
7VxJsBy8d1J6Q6tcqayPt1UFuJFfECAybfWzE1QYHsCclj9jFv6S8JlAqwR/CbcO
CIiuxuEjJZDaFWqZi5iuZYNeO//wSFeaDAJtjfQo6vR7W4X0eBF/4ydCM23YS7ki
DltPZkbJYnAWwaja/bnrCL9N3ezRKOwRbo6Cb6XoylfX6hC74DTjKdwarO//d20r
xZb0Bmn289INcx9Q1hlqNHC6J6yT3msA1T2y9t6uHe7iWtRUlyIPKMqJAeSmu8TI
xTwzgtFvfgARV/sCBnNEyhZUnsb8VY8O/BKGRJ5+g4RiTfBkxMpH7kHt3Ye1iBOY
0v+GOhOcnIu2tL8pU8VJn/9kNQ2zMZQ3+8Fw9PhOfqjhnFV+7DDbUe7x04jt5ROO
7su+skJB1YmzmtBqZM6unjl8lOBQ1GfuQL16VmXP+Z1sYijL0zBZYI2cwJupTFul
VTAleGoKpppqHmNv/gM19Wuf75i3Uv5VgsHPNgbbeVVSLhhkLi/lTOo48AELEPal
cwn0EDpVjLoznm/SUZKO4z3885T3DVLvPuO7tP3zQiDJg7R+R3GKnzc31nom1Fi1
Kudcl1tH2vn0D6hAiUdoHbd/e2zzdj9FtDGnPcfplHMw+/a6vcAVo7yfL2DJE7PB
p/dLhoU/X0BDi/P6uLhwqNwm01fSFWCUzZfs2tzV+BTE4SULfwHj5LHjA8MXefcx
Tt890oKA24LsSCkpDDhsIcIRqzvPSDnjewC1IDuhike1OwSYuzaFgsDJZ6gN5KuX
mOc/+gNGDdzN7EFpxisekHrK86uQKOPDJQKzdiqVJpwOyFFUJEHKlVZVC1JTToQA
FrCkAqsha9GE8QP0uSdYPS+ql/Qaqm6/BM2cehcYWkIHWH92vLsGvxucBTVX2kDj
kHRkeitbA+WctBZ52RfJXAeE0yqOqmkBupUASL5PyhI+jksAhMoiEiLPj3kR7YNx
hXOaGXOMeaBxjfc5TlRQ1mqtrM5m35GcQY8tPHiZSCr78PrHMTYTl+6wRJTV2eE/
3ueFq2cpHY1CV9K9vyTcSji6+d2yx4mfPtjEjjNKgPuVXtvza5agiqZJtjoTWGUo
mYLjpjo4UX4hfReX64P+bYXL+jv6lkMc5Es6c+Lb67ucwRU0h2E4ODcZ/GRyG5ky
0CGapys7ZhLYy5n3RpwzXp8/pI3uHbSYXa+97/9Usr5pZEDGUANDBO+aTM1/QOdg
emI2xGY2pSq6+d5a2zWqS3BK9w7KSm6O0QbFFIapKixEsUpR68wK6m6ljNYtm3rx
K/UV8Ad57TWkfw4LG/4JODH2OhilqrbCq2hO+mttPiy9RRLBbSMOxq/zSRkpUCc0
vl4a9gy/zel9S4UoBFUzUPs0roNTirs7J5QIiuVVFls5vo8JRhKEI7AuEtdRrNoh
YiuNuQhkdBa3tJ8YH2n/abYZOJ7AkN+yYoejkn/CToj6LljZ8hPLpFxD8qMWaioE
un8wRyCMVsUC5V9M+mOkoBfyqzIM1RCG6Jaa9PaQse4kVCeJshM54+yIgqQREArC
cgC/Qq8ub6pmQGLE7LotITnBJCrLV8SqpeC74CSTVhS5hhLxWMtaPDBFn5SunoRi
xNZrRuFSXQ1PpDUPrAoz7dYyK46JQxKvo9nmhbkFZWbse7LZW+1ueic9eUnMJA/n
8FmCjK+bJZwO7OPn4PujzxnAZvi3wKPpjMkY9KyJqtcJqqQk2jcJ1Ja8IsllUh5/
cWuFnPoEfUJjxIbs4ko9/1sK4Isxdp6RU+NM1SnnJw2yevI6NrGloH7KuI/KqAyp
BV4YVzOmCcZpw6wiKYrLQuGGmbLyAoR+r/gIiXSygc8qkCGd5873pK5z9u0MzmUu
G/EaBV6pG69AX74BUEAoOPBfsHEx1yLs9Y5TuPyGTo/6IALXW4jM69JabNilyQ+K
5b5Z+dK4BCPO1f3XL0oYGpl9RpFWbuU72hW/tkCOmJj5PkBMHBZ5ZGXxXfhkiy84
o4W/ugtjtZga4p+cZz4nZCSfo/xCr/e0BdMO0rO9Mp1j0tZ5CugjFe32+TcZN8vx
XPgxNqvQshLBLKXn9A6nVzyfaNkCGHRs8ZJwJg2tP+04MOTc7cSU9iHQYcSk8je5
nGwyilMS/qopP2lEVwDEWw62b6B/E3ET+gscAkU+XJst+Ld8pYvG+RR/cVypz1vN
G6J9B5ikGlcBtpX4PpI49XUFZ+3WgadgAvUMJsOLZtQ0qQsdgco5/9cH9op6bNBR
8ceqHF1P0tSLWPnZgIHMEdLylTmSI8PEwdc0pwAntGWPakiHZhNLIJcPlYMbwwH0
QH1TnX1khRKmfsaRX5rektcAwxDJ3eUCTo4eUrygPzUSbEtWYJOkK4lWfICe2s2p
urQ9NCzO+SjV3LubioZKPLPAJYxVD2PRSw6NyZj+RfI9a9xFpFs+7PZe2/uM4e98
l9bq68iNGB4Tk4PC+R43c4kuBg0qLK7UwZlZq7LoNL0g993kIqG8lt0jp3y0w+u1
L/vUAwJ7S8ZI0ZAdl9tZGApqtAzDZ89KXtP25hDvjx8aV5Lmb84qlpBVCXCB3igO
hCaGJQNIcgXUde3mp7shfbYOOqAZgUvcybTPnIDqqzRQfXwn2XLidXzHUqg9OV/0
ioMO4MO6V81J7+1pHG6rcoNbYV62PcbKmaSntoXyBZMZPRVpMgyIS2tjO0Mx2wHA
OCOzLhh6U7sDpudHOFOgTvGxn09wB9W2oa4ciHN5fagk7BduYFd4VwSMDvGTIV+W
8IoT1dUhgHo8hdsGOvZ08e4lsuTH1H84/D2uTPTu9lCfgIVM+xRxPfmMow+/jjo3
Tr0xT+XVhekbERJVf9hJccO/BhrO83hEqLLWVQtYVshPW4mOcridqGtKg8fHHSGv
EIr7sOFI7nlfPOn3yoIO7Jdu6Xhwzm9Mwb4tvgu/7476kGjl/xnCxGbYluKFVKCK
IZssXGMMNigzRHtvgfw8cfirDyn9DQ1txD0Mo8PONBAVUqb6W2L9F3eE/Yvo35xi
i8z64zMlphZlwzs7iNIGyB7C5TjzutHG+YKYtOEqftszM0clmC+z+nzaJhT1zNwe
2/PJsPo+ckEcc8XIU3uu7ipjitzHdR0wGWTYS4coMsmM7ANjboqMFBq3SKHV9Er9
xIqNoMbzufAwKE4/ffdz5WvVkOD4/CjNTPRtyBzjjWPA0LQygE1R0kE3XYvxq1E5
KpCiqEY0Qmd1Jx36KKFaBgw6d1LhXJ9+yo0SvLmr3JlX1iX6E9zVEvLMsWxug2DP
zFex9qDEKzlIdQGhnA2UMCm4enAb20FyurqeVJAXH55k9rGIJc7egmTnXLc72iZk
MGpz6JH6crsm76obG0LrRDzJE/OdgxM+xmtvgvfMsYJK3tkY0EI3TtGVWd28TOc2
D0LNahol7NPbAD9lDz6X0Ov+QFVA5lBl58vSJWFtuz8JXrgjsxmp+02R+d9N5VwE
ts5LycFfLvSITav8+SQDvk/0VuyqxkGlpZBdTcG7hvGchyaLDr0heSaNz1wvtR7M
wvBtTWW4U7yM21xH9zqXiFlGhRnYJMNRqllTS5F7zzlhW6Vqe2N01nfsPpSMi2ji
qMl4W//Zxf8VuZlGeMRr+qdUIOYJs2W6OmD0wKFNxrV2wxjRxDOfHdW9okF3worB
vNJEszKsIDAKYakzV+r5rnyp618ZWw8tkHjWuh/AkNInZJlQPpiYu21eptehPtTk
1h9zoUyukuaEjLP7f/cX/RQUHhXuD73koJ60zTH9brhzFkL8Rs9f5ZNql/WwnXe3
v28YhMPr4pi+ISCUURYYXCUSSxLGR2NtBhA99/otW1w/Y/w1gEPzfqYdPQUISHJA
Mj7E+1ykmMu9Jbz9887pezJAtAoTINcKPi6BktcOaKV4C94Js3G1tS8W5sGJiKE/
tYOnbyJqiAitx+BMkr6PWmuMmUKrsd7lAM4/Dq27l60BqrzF5WytXiFffl552Gci
8CimW29+y1e50Z26o7BZN+V+xtWmNdK9IdVz5bxp+y0RPSTwtkoCIRYHseG19WGa
YerZkKfOCLGbAGaTG6Gtxtmg00tT8sZFB35YosNs/eMLKOQ2199fV9265G8C4nSU
CLmIkvfUHKY9zgteaioO1toOV09nZOeVtHWY/FhdURukPJvT3OFEaO5mpHXVhMwj
UfiUbYJkbEatfMdmAuQ3EK7pGr/HJCRzAW03T0p3TuFOf0v0fYNkC3UeGax+Olvl
D2avAgFIrqhw67aTQW9j5GvKUTSvcWlpy6pBvEE5lkkiBadZe0uqTb9PDbJTW9Z6
0r0qf7worS45/rVe+jQB0F4TEK9CaOXZ91psLTfGqTAQZnuJbCsUQrvOxF0NcwIw
BiSGNRbayRKaWs/uezi6hrLjXSEM3NMTn5jtppXJRrzQ8KQ3An20gBoQKpN/updz
3Cf145fLCC36pTF9uTneBqwIhi4uspi1FnG63/D8zK3IuFkxyBSVTdClAsIFLdqQ
kPC2Drr8eDw9fetQ1+sRAGFEABgLL1u/yJIhhN8pD9SJguq26DljZixDmGHI6Gn9
3IugnTLIiH6jWMLww1XOW5ACJQi2Wp0mwqfN+IYeLIln4jHCuZFrEQt1sM7ebufI
jhy0KYWno3QJ2NXvc1NoXEbWg6IR+GHi5kPfcst9D0lk24mP+TjL5H/Ru/Bcrr5D
bXunDPDHcQOPw9xvKtmt1IHF6/9IsZSKIMj/7u/3NskhAsp42BayHFnQHe0BHor2
HNHxaBloKriK0VwaQ4arfETM/3Rmm2jESzpjhdddZeB35evbpPE3kz4t13500Hf6
D9kQ6RKOImcLPC0c3Sx/mmW5rKPZvLOKf9100HOlokaeQV6TVnQKcV8JxU8h5Pt7
LDj8xvkdJlvu8nDSXOUxMCmXGNxLxk7ybQhkwj7HVQVbQLckcdsh6y3aGgSAmT0I
HLmTAPGQgb9VAw+Z+sTMv7T1cjz/vg0FzUoUEZdp//71T5K1SasIUw/iBQ7Nk1AW
RL3IAJnewDfxTicvvYSWh36HeLbI20c643pa/fWjpnlEgk9GGuIB6arw9S6aaUjM
6oEp9vVPNo8+2990zan5Kecu0vZKTvEWtaho8zboZtXv8o0ozl/3ONfvqGxnmr7h
dudvJUWUy4n5Bdb1n75ejB452wbU+81ljYtGVelVhWOQmaQ8zOxNTu3B4sLkxOqj
cnegh7A4odY/wKOz23VPBVHvBnABK2/00HTGMg9H65tGt004jXZaaLI8EFPNzpE+
5/OIjHPNXKfyweDTHZ3E5jbOjmGxH24Q/TbPCzdEEMMOPxU/8Rqi1MlwucViABv3
HXzLtWdH2yALFFRr8QBVl0Hpi3ZfolQFKMHUU/FJRvfnn4Dw5HOFYzKh54FIN3uO
NwkSMnEND61M+J16mQuM+T8wMDSK9mGChIdhdPIEY7L4ZlXObSYsqkWjYVh1tb1h
b389/mTzj51/0Nu//uN2coAYTQ+kkxtSHl1jGZi8zBckzXDlaceF7EIqVPRF1Fyx
ff1L3gnjvo9qN8B6kjI9dGQJWgxOJiURMg3BhCzJnYQCyOdvpeIjwZTC/I5HbcxY
lOabd5FAdKhE9kFWlfjzOHK6cxcXOYaiA4hu2KyvIWsJMtfWEDetydzEtlGxFNF2
47J/QF6wvTEeaIGGfoIAcXA7DOBamyQ6G7b1lFE3drTITBb348/k6JWyG0L6U1Nj
F6zbAZFTSVAaF2W3em32sIX1HHoPRLE/lbeHIl2i6ZclzgMvsx/1hdH4a8xTV38O
wmMGJBaiVDdUnZo3L3kBjolrLTOnz9Jacr6hA+HrJTW9Gr2ZWg76GJ0sJzEmnXek
4bPYR915t6suNWHt5ii88RwH+80Bko/cjasEnMPjY6wg3wpR6uHDJl1ohFqEBjbf
+F4M1j2jw0pJmekel6ttuv8rjAUdB1QvNQY3tKq4PXRZttsokCegtoEEM6fGKIaV
lDMgiIY7XwJQxTjRjM40AoA8J9hpg+0CJFCRG/HFGtLV5xteqYJIElIq8JIkxGTz
rHMXBvE2gEicKDWT+AoADQmWH/+k2CQ7PLMj3Sr8aLernw/hj2GL7h+DMYqYL8YM
brWEx/j358/tL8XAMeOg5PGUsxGcgW3HOvppb9B4m4K/Zv1VSBzfwUbXvmxpqbxD
/Hgyc2mNWhvPEosFXjYktOTBzkoYQcjOL4MMPOQLodDQjLlqqgKgft6NaH13FYN4
4pCTWmvBXlUCsetdZUg/LV27Ww5WLgYWFRSJgL7i8yJWn1F/6hi7aWUm0mtFSJez
RRN7PE4u3uN4kwBDeuzuDpGuhRuk8TNVgtY61rEqTWeThRk1KkyUryPC4eq3R1rZ
XRB4DdwfCJKUFUfqha9yE4YczQvy5pM2qhOIIAYPEE8/f9qWMSGv1CxiTZOMq9NU
rJZ2or3ASVcwGvfBvCRo1SISrSZ/yAdq6S0FDuG68aTC8KRx8F5/zm/v4EojRcdT
wj4KDLzuUsdlgmkA1EMbyasbfsO8dFlloQCfj50FqX+2plURLsN84XJUIffU6z3w
I7WGh1SH/602Ui5SU42otOJx+w9veMThwvhjqIY6/0FIzzOQBFvnTDh9SXKfxp94
oFyb+P/3z14wg4DBDotiTdGbxOfWKpFTFaW35rlmTv4/GquQzdADo+yS9HJ3qpqe
csUINpMFc15QFzTT4aEeToN7MmoCghxRVStp+ispzOVSFleDkC5jOD0QHabQbtO2
Fb6EXaJOc+Tmz8eoNsajzC1zaYLGLR+n+wIyQQF5DMacYAi3WgccM+BTxHZkpyeO
T8sz+iEJtRo63pi14Y1AeYaIyTgHPW9QrcT9a3OvARwrgHKbW8oCXbJL+Sj4D/Dj
Bx9nE2pWSI7Hr8LO38MI/GqWf67afDTVAvmb8OOcaONTPXwsdWIuPZVZxoQrK72H
7Z9M4ijXRfHbs4iRINoTz7hZJqd1KTLRisfgkenGCeXRHAeciX6mrdeOsVBd84et
mYv9xxGIBekg2ZYj+Qfimyso58uLNZsUYZp2U7lJ/51DRc1Drq8i1b2geEbvF1lm
QK3dFGOmM25TdnJuiuCXneM2S0F9ZRGUz06x9bz9m088kFUiSBwuhG5ryLUk8Kjm
7xjvnsdLb5OwPyFmyl0LY617SBNwDBUm9mXcofP3X2wS2wXbqvTgruAIyfyBACRq
bpKelD23lofpaLmRYIQ/k78DktwZ7EGPiCmTZVEQUhn36fxunymNUd2/eqy41Eae
LkCJS8CSrCxVahSvaX0N4cFfmYYkYRAY3b1xnfxkhHqno0Z6I45Yw1n4kP3QfsfI
lpwexyh3M5SOi6Gm6xFNf+amzFtrfaZ/jXm0jN5oykouFokN2+fBWjd5qFX2mXyI
m991p2qMg+B6ZyapAcGbjbmaA0fUb617acKBxrI9Sii/4Kb+OfTRSK4YA1unm4Cr
yZ19kB0wNok/S+cOTi+J6YPdUxsk+ZW6YeM1ZqvuVTkAeYdH6ppwbpHuDKlW8tJU
iUUCBGs+cJXA1LYwjztCaV5ZTKUAEtmmrIcncWDo4zM6zK+MBAtYaQ1xbxbJdraO
+uL/+RrSHWudo+7ohEbegPem+6exHW1c56v0/sz1ZwAECDkh/wVw5mR839nhkkDm
8kMdx44x/G/tkL0kvshAu4b1pVE8tBy7Ul8XP2uQTF3wQtxQyTrmc/AnnbTwQ49Q
gyHgtchSRfQBxW4upbqipS+nD8zEWkHLJvEV+eNxjvmw2PQciPiL1soYk0RvfTm7
Bl4Lml2Rgeqn35VEjtSy7S2BeV5aLuRC41SUWQrgofoRAlWCpaRjVWSPKhXZ/rYG
oX0JI9edQROoZD4NEELYYx6ruKVKupzGIgvcw3RSZ8xL5vNQl5oZCBnjNhlx9eKw
lJz7I9BM3Rj9SrWifaI/sbysEj2R/gFlTnroiuWCKLHZQgcQWkqvziLN2VgLX/Z0
srJTXNYUYjhw/zebQWMXlh3JzuLVcBg1vBhvgDCxD4DqpS7wXc1Gdll0wn3zvdna
K9N+iFVlASNFOvlvaacHDFzvq9DzBm1IE3CgdvUdeWRyoJQXGeuzdl6OzI+96uBv
2n29Wy1og0RCH6fiIGYKZfaEf/YXgGM5HThuwGRE9/0iJIlg9fr9suGhMHxUVQuu
EU6Uzel3Zjgw3oJQrMs4G1XBFAqfbxP0el3EEoH0/dW7J5WVcS6GFb8DZkc3KRBO
dYjDxGtkJxOjceg5HWJIy/H1MZ6cGKhg+5bq98iwoCqLujzorGgyfd6zKn26bcrD
RtMdu13X+pY5LFeiFZBx1c7APtfDpk8LIs3H7ss4WSGC/GllqSsxpM/wUQ6tCamb
Q10Hsi/GU/rFRMmH0WuuuRgB8IP3W3ZAcDjJbScja4psCvaLgMwb14SPShieFosK
dUJROdnd7pRDV36XkV20cZUWNOU35lNdw3O7kN3D/kUJI3gycHrrSPl2PbOqva/v
QR21QUECI/UDVhSgPjiB4e36vzrXcF6mK2pOV7uZdrnLwjuXfwt8tYSyDdxa3bU+
54QFaVmd7RZR79LV1c8bPITMRN8ZkmbsyawOBCMUFzh0gfuPySBmUW69dzqcxSta
YWOhwxpRv+tGv3NPq/iZ8l6qvsMfeLVnkATqA1MMHp3GheRsyAAr9yhZRDQhjV5q
yIut1bnPoYqkUXrnzChxn+Q/x9l62uDkV0AImQw/psHJ45yexW+Z62lmlB1zuSQ3
/i15A9r144ugmnFRxd6CyHJ+6TBvojj0yW23mEagZwNZVVeo4VP+48uUuwcSsB2b
EHINFRmAALO2rhpyl+jQ59mfX9p5k/6f5UWVt7d72VjYSGrbH/gVJCY7YWUs/Qdn
my4jU1LwglMPStXCchibDqYs0Ft38ZjoLd8DnP04NGu67gRHP2WgkpXGjVCK5PRK
5NMA4FR8/ZtcDG/PjCbA0m6JRZaIEui9LtEoe10xUkjYxzaV7O1JrnRoukgqA9Ag
XKyOa1zQJCkspIAUEz0RswPs4Lvd0J5bqxOiWU3dBlhUe8iNCAWo6aCaBapA5OTs
i5LaEACqNC0oKR4roRbpDjrLIJqewPKkuO1Cp2eEYdgsEZ2ZkyohmhU/iFM8mrgB
7Krmg8493guzW84JwuiS37uy/HPdYaWZnSGcNuw4EVeOsk0UtBalcFyHz1Z/b2g4
pQSu3Qvww0ZrVFd8YqTuVyFRTCywl/KDqFgVsWIehqF+Ve6O0p4Ana+gz+6uwuDu
AfsKyruifYYxj+ikZK5/ril6VDW6q1pbwKNJEYJd9kIUiUU6KUIZoHAwyMvm5cXn
3VHoIQpdSam++LV6LaMEjcOXEAVecotE6b69+4RqtSP2es7hPFyIXVdav3aMTxyv
Zw2HaK1bfZTCtCwKQA9wWOrlHqdhj76mb5AdEqbOOtsmTilpRXlzG8IJFNZzX64s
rXlMODeuN2wFesmJO9p7gVGWaqfi2VD/1jm19rVQSAFPDmDwVjBMyUaijoLw2jp2
2atXQmgKu2+pGes8mHjp5ZR0yJVOjpcqaohN9PO62f5a2n44FtMAbPR6a0iVGluO
4QvzMNM1cgO+KTcVt6a78QK9rsGBGydfTQXR2SDLXo4lPFPlmkrg2tiJRHtWd6T2
wZlLN2kUq1NPwiXRDzyeIg1/PM/9Muc+wHdex+yhhPOJhWMJQ/E+colkGKXemwZJ
sxPFEsvm5OPovun9lh8dZFvSEsnDDISoHifepC6jw5UEw3BFXCwrz/TSXmAnzMbT
LZpo9eVp3D9oR7CAMs+fDShcLKA5Njq3G4n9yC+nWo7smHfxOrgF6jq+yK5QECRj
IrG8u/CjeEl7baiMaUE+9wUcP720cfgscK/wLgTKtEhs/Qszyylt1TOkqKRWUDWD
dbFPPpmSwAG/gXHFcLdEBV030w1fxH8fNwyGYu7/E7b0Tl+0XMPPhdCMJPVJyJwu
JxnfgWwlhbY6YbakHDJBMjTT3Xwkq0l+gXLj7wFXC6+WlsaW+7KwEotLo6GXDacN
k2d5w28xbQdSLhwYR1JsfeeKY6GQF2B2GTMcIlP6InRhe1d/g2uT6Zpyn6FhY7M2
cb/RRJ44m7ovR4+n6jUT9aWHP10CxhZhDSL9Mn+gS6LjdBALWxKmxKExjE8XnUxW
lt2I1bskVs3PHMhwBKwNvYkAesYUGPTV6JW48TZp74bV9eBwufaX+921VsUq7M5g
vLieSknK7TZ6tDoCS4nZ48c7a3UQwXkhsrWqOvT58qTHhDCzmH15E5poCXglzEDJ
LjSsj9C1CCC5O4aYCIV24r7SU7nDSkqHbztLPBv15zZ6sB3lOW/p/j0e3LyFoFS0
9zzBRbVaLj0Ojcj+h8uv8Q4MID2Rwhkc/THV9DsuHK6dcIKN3qHvbJM7liQ7e6uo
WCnjLDkO0mflcISzsKfW4cJxX8aFKZiecmbiwepu0hVeHH2vlxbhHtjhv+ZoMivC
lCwxhlpi8QAkoBVUo+G6gj+HlxvMXDhLJnfi2IyhTELZQHGLYbYn8G2SauKuMQL5
Fi83iDwBdGlYY1PbIitFGZtT+E71o6X80d9bVvdIeWwQjsHiOwJ+E340jb+SFHn3
BaKEHWV97luuL42nvzB2fOQXRdwaGeLBQEHiTNBv8DqvtceL5eso1djOI15wc3q2
pfc+5APLfxlNCSmFGZWTzZecwU8q04A3a+hWDd1sT7Hs9f6+giTfTVOmxbvy+yFH
OBlyzxjXvEmaI4SMhQaHRXInJgWTmRuBfKE66nFgeDxGBQ4XIEmJDFV88hKhbtN1
vrNegFlVpQIcms7ixahoINLrWjs+VpwirHmpgbfXYnlZp2xivI1e6pWdbEqxRZzA
S/suMRpCRuGXMgjuNkW4jaqvt9cFzApONivmkEHNxkQUuoTJ0+71P90RVI1Bdq6s
hEImo6upWTf4k2Yc37cdGfJbd9vz/wyUsJINO7SCzOlIhPHyyUzjyZ5XH86l7Ey9
fstru2/V2hwIKCgNuzNf1WKwIq33iIirF9cf9x1pgGZj4Q/qh6Tf7ksMf0PohHDQ
g83YrdyRrhlVmLwABz59NIcQ4cAH/yoZrc5zkHCN9y2O6rQ208lrHnweMWRzVS6J
GHYeEmFwauk83Krg9nuGd/jhctDek7Jj7REhyw+cr/3Db9ZP21TBWJMSCfJGirit
yGk/UHN3vpCrUcCcwUrXSM0QfViVL+iZG/4+u8t6eASjxB8Q3q4K0j3uamEvkdpe
R9ZeMpxZiJ3bG4e4ZuT328R6Rp25ZjJX9Mdj41X/xNX3Dk5dnSWlB6ppVxMOe/Ye
pts49YL9oNrM0kNaYVW1w9PgoK5oRspCyMn3yO22yhT3dtydwxXIXl1vNceADhZZ
4tYlYQpQjr2lRRF+jVqcFQekGkvVWAyJqZxgAKU9Qk9hSmh7r85B49BsdPZ3krMG
extErWo7igW1EpSlIfTuQyqjWRjtKKfXXl67Cbjpmi/cACnPB+ARCyf7PDIpQQk9
uIj4RqkKWN4yfLyxMdO2ntCSGZiysOG4Pa8zquBngWaDC7L0NZmMx3UQ7v15Kwxk
ZdzYZcJZuYnp29r3k72/JFhZrqo+crvhc82wYsnybYHNEinSy7nYCcWiRDovqspW
HIKx9WLlc8hMvOvlBTU02IlWy/JQcr8l8Wbq7OtQbLgzZ+AuimTwdyyyCJaf6Zvm
o1M7IOAmlrW7CJVo14oohRincQj9bH6SR3/GcUEzTSNtqHcfeVyg0S1cm9NjifDL
08LiMMIcxEs1g8/xiB0WE+orjVYufZsB3yxbE5y85sh0QIG/wK8uSYpl3S3mMr/+
DJyfwORM8w352Hu055tLh1LOViBJsVj1XFu7mf7T3JhT+KSaFUxKkiUC5SmyVG4J
LE3HxpqcIq0jM66vhGDpkcdMde+X3vPZFTjpm+JjBD2B6nOEsQCWjOP6P4whG/mC
bWXa8qzHAboFGumhPccIg9+HeifxP09cR63MaXuP07x9hHaiL65tDgrhdiJaOFN1
WQsZbXDQ5SWlrSBx4Rtpy2VSlwkFIt5wgLpZyDe4hsjHLVdHxMXLSi+tDZEf2MeF
QFDZkhGS69aWMl+VQmtIaagX8A2swzmu7LQAs8FOZl6PGNS7hYRRHwSH+0+tTnsp
9SxAhVLmZ32Ru88rMQ7vlWCUeKpoT5zSG0pxei0MjrP1cxsUbdOIpukqYxPdHZbe
MX3ytRgfDsKAjO8Z5VoTxmf66pCgVeljtG4M048siJlUsppZreq+nRdBi5KbOZwI
M5xFaAivsVlrUB94bVO8DFRqjllBldjfEeH/nYdOiB/ufFPSZ9PR6TA9912R8szY
U3C4MQyubF8ahQTraHbKSWR8aRv21JSXER9r8Dk/bSKqwFYixJ5EcRPFjnjruA+Z
LSBDGlTaZ2wSZ/7uez5qPd0R3E++tV/XMRw7Gx6K7GcoRfRUeyYNkCTcCcwTTPCz
s5G/sV9NYBeEmxyuTLgAqI/WUMIHM6fko4hxdBaaCsJcHE+khLmxA1af4OISc+7E
00gUlwohvvVM56hrbozyXxTCUGIkhC1/o+KDzmLi/rmDN0+taEmHxSbCvZhPWLC9
xMk4PipqWyhgyMBuMdLAxnr/bfPrsqx+/QqbVtZbDJ/HG6uM196HojX5On/KA1kz
rpuBMJ+ysYN+UpTOFSnJcBGINXO0VS+UAvGlOizNiRi/47UnXCQOIfZ/e8N7J48S
teLbtraUKLGvHoRJ5mConteJ6LA7x93yCTurYel7/xNalI0gxxbAdQ3KJZA4ufML
YSqBfmdBIpwZKTAdMJJ3YU8wMCD+P9uds81IOOJRiVJ6Iht8xUPQq3tbb7UBnpno
Amxsuuz/7SEBQPdieVBty0imm2qNzJfrcRpOmr5F3sgQkEO4wXj/xvWphCgVdlOh
22GriYk2ehfGV6R6nCukvuZ0kJlNgPy+ynw83eCGBZMRzCm3+qT0HLa7MYyUWw+H
pHqEdsxQ8vrGk1VrNRSFq9ZNKDs2cEzCAz2K6IgDsCTLZnJL/Z2ZvGTgWX5Gh+1P
/yUng4cCl7fA2p6gzt9sycTr7zhim/vFHq2z64y3QPOAJwYhvYbKW4k7tRSrGzve
dTgJyRf0qhJWRdtscfEoBetWX8jPPDjAEh4Gook3aVfJ21NUkBEC5z/bvMoE6+yQ
qRJfo+mZnDIbNzDCDsH6ybSePwA/K4gutJ0q32vWCKs5DtL3UTwmxx17RtHK2jP1
lZ0i8txKJLN5NwvY8CyJmsy3F1VWsI4j9e3wIAKxTG2yo1aGC+sQ9h0cB4rAHuu9
7wp2V3GdyryGCfya1BrjgghoF0hqg4ZJlbr7kQAIrVN3nn/K+Bz15+jbGQ0PE7bt
U6q8reJv2Y9b7eJN/Ec1nK8DMVuaC74SqvMFXAw/cD+w1oILPkZqaaeE2trKSq47
BesFlLL5MfRoQt4rM1GB89uhmrFsnZE+cO8+sYI6H3oMlbzla3DLAfsSQUpxvNsa
4QfgPoHeta1Q8w1QphH8pFsZlNAcHvIVGxYB0hhs505UclKlvYjZuPZp54X0BJ1k
6R5bTj2ILKdX6b+KKdcloAJMtYGkvYEKNGp3VfSXSTxEUBok8+fGTqqgp5m5fjlj
d5dfhAjeVuczhxjNEKOObeMquqjrPpfJqmL1jjBTOTmY8XYLYqGYOymXhLH0VC8d
LLb2r/b61I81G1W4PQ0IWtj37f1Tlpq5I86SLv9coJl5oEs5GibvJzFFqEtDMhcJ
Zslqw2DQ50CK15so5uZ2rrxgKtZ2Z3YWJdsEVVSOiKDqWJh10LHVUYfhrhug8c2p
PeZRomeyKBhw6kOPoBvZZWpvocpyrjlmDQWUbEJY0l9+VK77aW0grxNW8mMMReq2
rOrQOcwK/aJEYoPWUPJNULisrxHiF4ospbE2XSDr5tip/ufZ6972qhxYfAHzbq4h
jDJMu1/zEmBsFJqzrMsAucuXUlK5VXld9j6weT43hVkQEsvv9s00pC/GrS4xzh6P
DvXgtBk5dAqWqRZpM9O9rlE2H7NNL+ewrJbc/RpPL3cDAbKVeTc+6vDjx88Y7zqc
i14v09eyvvF8hcad4LV7JDAaF9l2g1oqUOtnxa9L9WvFb28JhZHudByFTPprNm84
8T8tMp7gX2JQ5P9L43i7c/fO43j5ddp5gXCyoSOqNCmaPMhA450dSk/lZ6R6fatT
dsXGqQkEGdhFrCtDCwZbHiX9tZG44r2fLcymhCV9Zac0jFXsHetxAVkEWuatSaxD
pF8K+5qKdmy/2rQIZnWqDzLwcRDb2zPmXW9L8qsOXIo52TcQ+g+YwKADVsY6PJtI
x96hV0xHx/GTU3WtGGsy1JlB0+kBM8nrfepGw6li5DgXUs8OmxPCzPWQ8nW4tJ8A
YxkUwgTdASu8NaGNt2JTbkfuEQl+ZXEBRb26+V6DcIha4hlc/KfvEQ8aIfMMZRnk
e/mOn7tDD+2hZEMK6IheDWetUixHpGJYr0rkzUITxCt9GEK3Redam4F2GiWPGX4U
0wDUlcfjpDgTBiq18j2iTVRiyM2889xSQOlC8o2aoZQfQUYUkX+oYYFCW1qNC6H0
nzgrPZs2ib+r207hWMZaySkPhWaeLngn3QKIuass6RDStxeaxCU9GMxS42Yyvtvs
Zva35oGqifkPxTEOMQcAcJGRM6wZlWR/KXLcGd3Ei6cBBaEf5RSozAJFpN0Y5WWd
nV2H+9yTPWIVbKjR6aX3Rqvuage73xWgGKFquXLqkAKeHjsSInQFnH5VW/+Pz1kN
/bpa44NQJW6NCqaGbTNRFpWBWY7mEv7HMsEaxrgzG1cZWi8T8C4rsjOudNfjV+P7
4V89WFTenlS0veRHJi1U/scaY21VPdLh/koDAu+FwoGqG7tQtrCfhdI1M7JYGhTY
zaMTp8wTEStpo64g55iV6putX5IQkTRBkg9+xuAnzCygb8073a3thkebnbHORDrg
pola3yfuzoN5cwlp79QyceO1oFTo/GTmFTph+UK334Y80VaGydHMIuWaOEiuN9SD
pTZ5TW2diC6q+eWXmDjh4owt1hC9Z1kyYmio66C285SWSVBdfxQaxBu6OsfDzfQf
8pi6CpJfHxQr5YNkJGDe8H/2zb2bpkQ6kFkHbveVbKZRjhg/sh4U1Sq5qWMJ08tH
f7WpkIgKeof3l1H3yEQjfWV0fOICeC6N1nQncyiPPfoJy9HiDDJo/N6h8YbIUxak
uZ6GmGc/+tQu3LKCzXDB2XUANSdcikE2JRLuLy+HtqHfhA4DrMV6JW9SHrvcCTDW
laRchCLBvNyc14xIekqQt76uKmRNZTffvAUknsDOjZeAd3H6lmT0+H295+eq35AK
dY0j7x9Y1t3JhUOrH1LfptFtyYqU5Zq9jHsLsRjJ+9bUKFZW+iPq3nksh4tzNoTU
C0StIMmp97tUNY/YrM6C6T4fnN/4wixKddnG2fMgCWbNMKMd3gS3BMkDv8xIPE9l
LeLye500NQuQUYptogG6JRiC3S+NHDwvwfDpwbW7exGYQ8C9bpeXQydwtqqtHG1i
aWt7CFg75lNRM3vY45jn1MIv9tjzarYDyDrSoccE3t2fPyRF4DWn9LMZQxroNhKH
LOSGkJl3RFK+272xxdiyHxF8Swu9Igo6/NtW1WZBF01j7llnEMZbqZC+fjuwRVNg
Oldp3IOksX/zc7vY9dQNZ+wQuycJ6TNL6bgNJlwrq3b+lOHvlD2eZ0hZpt2AQ3KB
e+JC7Dr9yWJJsrrH5JQxbvn6mbGgiZzDrL2JxaJgYrORIHPZ9lUEhY3fKO83n00s
eVC9u9zZRqu9h3OGakO//lEdd+GkoC9Vo538KHaKLWzTHp6LuvRCVpPi/3TNV+Xp
sZ58cWYzRWB3nfynNxIEgfTFS1SLYD5Tef+ONGK5gFugLhGRipM1kvuScmhiyLqY
rXVWiTuA+xiT6eZmt3Tnc5YmFZVc2q1GHDc2dlEcGtc9o7cY1L/W11o9d9NeDGef
Ive8LEHNsOngqBspityvEsP0+GvWXq2qbx5YEopUhzn9Gpbys0m0hALGHYdCb+Z3
1MCLMiR2a68W95D27+eq7vR9KFiyi1qr2GUCXcnnpxEoWLFC5ZbQUAHlvVbOPXWP
7qmK6t7KB3LKWmv0z1J1/WMeOXxFUJWYoKR+4sx8HSgrnRwmrpZo90LVajs2m117
GZC+otgFowQRE7jq2cMBdNo5WPcWcGcixeJuI3cKIvasBYR+y3QBDZMPd2TVK17L
GTY+animjOOYIkZrNhwfjbaeKm4tmXBMqRTXiCa0gUHUnJDGBmmMxpSTgjoARnXk
ov0ATOQx9scSbsTBxHcsVtofrEsJGSRflbfCHJ5ZdXj6QI/C+SspBwqfqC06TMVt
VKJLmPn+anHXLNTZGRH2IwkYUx6h7SfyGUbjTyRgACai1cw79MVcAKWqeIYL2QQL
T5Zupx8D+Sl7stQRfwdeuXkkfKdqlweeeAL0+o1pmjq/3AswbqQ9MP8fZcDRoGuJ
NJcg1e5Nr3UAk0gupM4O2HjjP7ujCUX/0sg25FWvlOC3gdBNkZO/mmC+PNfMHSjm
u1qBqnoCiaM2XtOkMphnGzaAYfJw32kaYbasqhux27qiGJXeqwkOHzifq3W+iXBf
vlVvBEWFzcS4+oFAT8yQ9AG9jx+0TTQcNYDWnqIV44Ol8CQae7rnuVnxya+NJF/R
7nhANYxZduF/sYXHGjOMr/Ws+/GigXNAn5zJjzwU8E+KN1E71qGl1okT0arGvoFz
To8IoA/1ASHz+sQiZDP83VFxl5TiSJSXMmsifVpxCHFvDr94SXRpYF5z7UtDA56X
/2f3rwii3aC2J/WeIby5yEVuTk5wFrPPelZm3by/TBMWWkiExJ8tIaG72DQpLQsz
MgnfCLCImW/J1kk57wlfQXoKhzJs4eGafmK3vLUTeqteAFFOOnW5qQc4u4EiycTs
Be1FiMlSYjwIZVwmsRIc0tftOYlfR+YIi8X0vByfZK1MnY69VK648XQmkiZzl6/P
kpeSit46MMBZ9YUg6HEGljjMAmI9SpfU3VmZLhof9ajm4Xxs0dvU+NSRaqgqpStd
qbZJjMe1VRHZkIjaUK2H8Nd/iO/XDOR+ioXZdEN94JNJiRsMMLy6wsNx7vCLtmlT
yKHDTfCtA7WjJkvHSOSWXy9dMLRf71fb9PneJoBc3cwbAVVNvcDkmvmAGLYz1TdZ
3x/qYOjoouzoih/4e5hSmHYZezWJpgYT0XPVn4ofrgBhk2CwJAQTLTLDCyEeB/fD
a4DXXYVWopx5QSQTboqecuhxC/xZAEaMnYfmpsHfFEuPm/NOb5ejrroxgrNUBauF
LokYUN+GAzpp4jAczfYQSwxiiGJ5v7zF+N5Qp3P5wuj1+9mT2slWEqsDk/hF63Fj
BAyHExO3NXNC72XEzvr3yxoJTbnhybF85Hxw1wwGevWakeGwJ4wuV/PlPcUNzv+V
VNPDWBWvzrRsC3b8cei2jjPkOMfz+HPK9sjQXomgiZPiYzt1Qi+8BauofO+iFiri
mdqmDHDJmiggSBay1GmMenRV1eaPVyxjp92aYvhNItcEtq5G1rJ/lW9vyIEEB6Pv
KNNepo+3w2srac1f/+bvk6NpUuJLiy5OyR/nSkHefhCKUs9g+tYCLb7sA9FbjkxK
Jyo6EzAj6kRrZkMmjnq+GjBCDiKKA11faadmLV/ogF41s1Lpv7OuzpxKgGuQof7G
Zwq3E1IAyHYXQnQRDL4rGO+fU9Z0WjPIYCRu28x9PRwUjpwn4H6UqDdKOxZhIZZz

--pragma protect end_data_block
--pragma protect digest_block
rJ6QAhqf3Z7UBE3QNw4iXppUIl0=
--pragma protect end_digest_block
--pragma protect end_protected
