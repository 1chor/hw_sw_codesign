-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
I/0i0Dnh5XA4pk8Fyj+CKuBWP554DJLNKr7A2pdVaCbmtPbkQ7BID/xj76z0ExMc
EWX1D4DsDD1SxnlTIRFrTJ5w7avXP0GjkT5MntNpuBn1t4HRXUE3ONItEtX1XXCP
SR8Og3zkG4sfK+F+aq/FC7JC7d1FVswvISt024u/mGM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 88393)

`protect DATA_BLOCK
s25t7FFK+0Z+IVTWoipD9TJIIEb53pZCg6TKnCDY33PlPdI6pNSI09cuOJhfKuiL
YFevWhWwuYiTOCYvPyFgXFR7YYBD00/NtEADQMSy1swCekSCRJG7GH1mJyOcPFAU
PSTXpGrJgNceV2FpwRIubt5eMMd3D8TiplAZX9mB2NeaturkyIqvUfYK0vyE1F9L
1k0BUT2gDCiiJimI7KPJHV/Gcb3/+oIGzMvi4BOSpSsWNEiva1eEBin0LwE9aW91
tp06ydkV8nPbQ3y739GpbM3OWK31MYYw+qHfrBVCi+9slsVY3HLTrAbxmbFoZ+vT
vBCwK+WvlLKKzVOGNQfbvOp8W4e/+aqb2mvzmO6Vn5leH8nEGTw2/UaDXduAPSrv
enLe9CIKz+qOrFtBTcPFFuj3+u/FcMQaPuJ1oX1CHVa7sTB6T/U6MdGtoX4jxpiG
zHjaw3iIF7fGX8yNwH1nfY0XOpMAmIQPDDlo7IuekvZEHaxBswUcmXtS785V+Smc
iBsZ9T2ycfHayQ/zwv13KnbBTFVqZsXzKW+B4I2X5h6jkOhLeyz1NZMpsvR6nJX9
dVzYjqljj/zkVOQeGjz4giNMSkkIb1IOut/jjmLlw0MrjvJuyo1LxTQCMwuQUnLv
ZqlUccSw4H+by8gRiLo6E/BoK7OY7fVr1FBfVvcui1hf50cOKrVTOKejRAt1G4Y9
SwtYaLalTrqizY6Mr1IGqlxTwQFsiYHgckAso5A6SWyeER98G8IGcjyuPgqbEhSt
hGxGfx3TfuDEQh4iPAMnkYtzws0ePwW1mJvfNoucMKBz1c/FxFXLaTo4AJhwTOMI
tZLBHqQk741DHlJrgTleryQUEx3P4ivqA3MzkNyAy9O3zAOQvr8AyDQGlBnR+kvw
Ml7M4N/DCnh9ouqTywaOXcej3qnBTchdwvjMFGJQfs2WNi//5U9Q9htLvCyWnGwo
ppeUPLCnDOvyQGCZvL0zawQQS9R4wWMI2Ho8ScrB74I8xZLo7hMSPUyogVjZ74LH
jN2mo3F4twRVd/sPl2kNosvk6UzAmcATch5RXqgEwBaevDtuisWtGxoNHorz63rv
lCRdL5iepYgBy34Sf1N0SjGfLoC6NEakcY9RExUVo/3Zj/F6UqLEn5OBgVSKjJra
/nE9Hzdf6AvM94tY/f02+z94u55J07T9n3oIwakixg1nt8obf2ZdriaPKRpRR8rS
2LTGuq8LGV7lR/ii+Zr1HXwwwLyxPvWAJPtUelRbJcheX/Zsn2ozEvDU30V5xx/o
FMrzyMiujQjb7lIItfhJ4TtNGwJxK79vbnJ7Mmzpbkp2229UJO9VUesl056A6u5z
kmv1qPR06BeHhb/Nb24CcdsdazNU5eUowhi0s26pDQ6vu0HhrvZbXDigB4Pg9eXF
OOKSSFKYWm9C4AuTtPkJMoV1NWR14M/Q/OXJXY3zSDC2S5WzukLbxy3KAYjmx4Yj
gZBeu2dIyd8wule4cqSYructZjXhrRrTVxa2rcgMkrsoWX2JiilWmiTGI/m2aVdM
bKxVb9dhuMdwcW/Ce+6XnNRnkPxgxuOmF1pyZ5ei6ohs78bwvryelIPND0ETtgyV
uxC+1z9PP9sdUL46/fURysHHRw91vm3DA/ZDEhC6qSfY8JyRVObe9Bo3dLtj7wqY
CYtBA2hsCXoO5VWzZilNtSzKLuXQt/zoZatVjySo1056jsRkdysj7X35SBySxY7+
axCFYRQpSDQdz5CoNgNcPAISx8KioG9NovHfU/4E97dAIFMIu+zct3qfXCICZzhg
RSaVfqWOMJfKhO5lzJ+a/C1iL7q9QzDH+nDcBSYtVZC1MEX/9xj+6xFaC4h/OeKw
StbybS7NtdCcPPhP1sRu6johOVceH9mEQhhOE/V4DqnouEHOpevuKTE9ZtBHIapd
O0B//gTBWhFHLPw9cpPlZHC8oRW1eVLkAGmyxhKgsBms1ge6SauaqLglSpVlA9FY
9zd8oRZEA+FBqG7vYfWtKwRhug1yqnBuwspRLH01+9clcBKCz8nilaypdOanwNPr
3lkDNqVUDflFuAZ+Ren8EqiYuUo0AwbiVcR+sQORQJBJ91zjumXbFcR0zXdXQea0
6+Hugeo/56EC/UndPXdxPXb6Tz+/Ft8y5aAoIgJm41DCJj/DrYYyftXNFk9SJrF8
0TjeRzdsllhX6zgiBWGeCNvwPm9jIWCUWXJTErLzXDBmFjZ9uvOYik7mgCXotepN
aERXzX4/hILoKLF9UBC+CZrNynoW7+3H/Pc0OtUU+VffR4hUqGfnduP4Nj8+GiYR
w2oL/yjAwavPXfJj5CYyjstGBtHcqIS631T8RkooWLlYy9cp/zH9AhNBuel11Yuw
ecdBaW5DqBjE4F3j8voX9C6Im0NCDzWjmVopS9bwa+JRk4WqAF9z5p0st3TFOrU5
y/527MSM17kJLE7f9o9AiIgWa+sHmJ5yJDOEANI8818t8ulg3Ir63YjyrHKAerdD
f/HitcEdyZD7nKGWa48nPjjW/C63ZrNhWrBKWVGghUQeJ/1LL5cw1P4u1jNXhETF
LQf0zhxcHJi3/RjVeLWOl/qjyiQYu85rBKgQ00Wpi6Ex9tuZs14ZhMQYp9Md6jN/
BdemRC+6mAEy3DKUn9p2UQmXcg0wWNGxSrujXg4la6LIkMD1siypYDRyeBZDzIUe
q/r+85eei11ruKbEf2JkM2+clCJT8X+JssRawHd55wveNXdLK5wxQgszhZAFYaa3
QT8Ut5dW2mSZpF5artMDp0Mnd0XTdq8KFRgPOYNq2YttEJu/WUzVIWg+obC+SuyF
UfFiV8XTenEPP7tTa4QoOCJnRuakajgJuAsWRZyomhMq89D3z120bhoK3nAB7qAZ
3UGammv5Dgbre9bc4Gnv50hrl2mQQhqLbLK1tlHGvJ7lQOpZrkN7Tj8/rjtGAMtA
khoClgT2fn7eC9ljihKowmBL+xKGT6XL2TsmSsX1rrGu2ClN52lJbQIcA1mH9Lw0
oGTzCnIgNfQ7yk6ieBuotstQ1pp6OJVUQQGo/NZ8nFVuT0CXvK8Sf6U8nBw6ZczW
nxEs/sj6Y1aVjut1U4LhPhAifn7ZTETpnM7ZQy+5V7cTcOqHD5OOIDxbxDlNXMh+
t0MjBiQ8pp1AWlXe2HclD/7dHw8z99Mnox5hJiU9J8F3+SmFXelK2Yj6y8Ifw1zH
vME5gria4TfK3ngCqOzEOwwuj4brvRF5arnG5Rnf+u1fRX78zF2HeewLZGW1TK9a
D03l5aylFH16Y2BonyCUElsQi3dzTMqQ1y/Oot5xA76Nx8IHCf3qX3b8SK3omif6
B0g3WTKN55+ZMZnj9otSIVg9lvDU5DK575+kVPENl2ckMiRiPt+ZLJuNvyTxZP73
JIpUZOww8aeKux1XYVhPhXDYwoqoLNVrN/pnhUIt4WKTwaNaiRsXkoaRNjCa9cdY
J3wkwTWDp6RDXkSh8rMZX5eOGpDcx0A39zN8Ut+Uvp3YHFUf1Tw8Y4YPt8BmFn7v
kg4mmE8VP5qi9oDiXf48kN1eiNRajfCpq4o50gfc3d97nNdUnaluNlDDQHpZUxMd
41H5ZJf+pWTZDa0a0d4JRxYPqDXqO+eSDZ68PWTTRIYV8DhPUDE3LuWjjOflMb+9
EDvs8bkfjnMBDjUPWoKdJHlhuTCs0zQYOGuA0VrQdXqQwOby+eL0FKbfDdRpcZ23
iUlQjSZ7zqXcb7yJ3WxZ7ueoSM9rOtg44Q5Q/IMRNhKGe2QXNaDi4OEORzsKmkbO
UbuOGVQnOGKy/xUHMo6nHBQDv4ItiQZSri4obz+OIpCJAA6jwBO+g8XiT79rL0O3
XXitmCNZfpmxkOjMFpVjWjvrc6A3yTVsD+SqJCLXEfLDTC3UvDVEL8z3iW/7uEoA
W2vKvat0DR4b2/4JOsdfxmHzt3QBOu6Vj+t7owHAPzaGmcclzXqPVCBPTlaXLumo
hlR4INoLBP59JNe/adDLzjWE9tsO68ZEYigMOXZ7XZmkMyQwgDmwRMVeUZDcsg1x
bwELPKnZYGRmvAHDNZwrzh86gW95v37enRyQBDv++6phsEs5eQKtpoMh0yxjJwf8
VNnVuYpy0G7h/pT1tF5yxsReNoGd95d1mLM3+QwzzXJSmphmuT96XugaDiMX22YS
bYRvqCAYdVmx7OdbePrAnaFtqdDYBJh2j1hU7n0RmGIMz8ejmVpWYMCfMbf+sjgd
hRmJ9Izs1lCRCoHemTom4hfixcKKMQoKw+0+8mhrsMxKH9YdiumnnsVHdOtqM6jX
vQmmNVLqj5mjB26j7almuNO8w40HZLmu7ui40VFJ0I2xMiBxQVq4g3tHjyyQlPSE
Ih900u9qIfNDo8Yp2GdFNHdoSodUnulrmT95G46Mla7C7ckWCOX6UHtqDAYIW1d+
Ozx5tW7do5z7BCjbJ8slufGYFS/7vGQk0keur8N+/y8wNdECSbIK7YxuGKfelb6F
PQe1fL4JhGNq3hz1PXxgwBDGFn0j9rqhE6fY0XiQoPFQ9uEsBgzUxMNC7L/Ezl0g
Sd4VwmRlrltbkaxkmjZXijmk9SKdFcnwdz3J7GiBhKlbBij6yYPfNnCtyHFNWlzQ
JOHjbGKuKVw3DFptbDOIKEDo/qoLXhwDkPonlJjNvshOchyiYCK8HF8muJZD6eHP
SOi8ems849GREUTWaoOLjPprWKagffZmR/qRUIf0NfQBhsxUigZYZWgf7m6kNFLD
OTHiN5q9LgXC2PQpn6BKEHbzXwlyk/nTgiOcrD/nQTc9PCqVtzyQaBksb/sJ+dsq
oVPB297g6nWOmAZ1D0/95qtm+4URtJIQ5l4jwz4eJqEjA2w2zbPxxMnQhpWa2cXk
pAmWPwxGfYfkjDMWovuEbiZ1IYvLcfpDkTksb8l6MdT96pbbgvaLn4b82PdaKXTp
54SpLMLQ3Pi+k6I9Sxt8xi1kTVOlk5k/6NYk328gmk+5n2bCzP6CrFiB55mP/Ybp
3FyStjqCeIaqejy7Jhkg4xbwZaX/XqlOTyj4uyaDAsYX71+Qtzzd4DggZZWkNoy2
9yLY/lIU5c0jNMLY2kwWw+NeDiL1PSYW/zRLD4Dk9uupxeXZj6aOHGrDQ+6Q69LF
jPEYcvZHV/jfwWaTpjgZz55i+bCg0eK+CT6WeNs3ca5AfFGAEHUqQ7++vSN879Pf
6/KQ1rUJ1FK13v1845tYDIdjxebYyBWUSyCB4/vvsUJtUfTJLFE6Q3wWq3Sy/16o
RorRrYjlCDdyzkZMfc4ZrNiFUeXyKizh+w0V+3K48Bpd85eaCW4zzGfsIWMqbMR2
JKSVqUsH1w5gSL/YdmpghaSSo6qtmFUBDR1jaskvdo/Z4lggumW+A3q80/GSTDJ/
aLvx4EuBH2gQ1/lw8Ux4L44U93gj5WdCGgwfHW4IP9gqvWpaeD4Cf8WsY8xfXXMh
WEarV+9DhQ8M5K4N0SrcLHr8wLZ617mEsNv4j/77pf8eLKWC/nGCtiGyOxuhctFM
FD45J7nDmzUXJdW4HetSGVruH9/Z+50hN9odJzGS3qk1UdZ4+3g7zLbN678lYPZR
iXeJLxmBOoBmb0DgigWcEfyWKc8qUsDRwohCgaoUJtRSH7f1pzPTU3nxUz3A5LI1
awajfAQ+z9irgjj/qKC4wKeWFrK5ucMimyyTzrDDgnyRg1AMkTqoUk2gc6yjeyLk
BPWDjzKVEd6SXlrHSb5Jx1WN3u5u5H+5OScv2V1uqXTf6JNDP+sLxeZKBtWHWmyI
50zUhkkNIm+vUSqY1QNNoSa6mIAbHSeSBWNNwVZXBYj/yMdbM1roCGscZtulXTgE
hwucUpxTpDxuhAdXz2cBHtt4VS1PEzyu8FdCz/N+PjOb72W7e4MY+5R4nIyv49h/
uBaFAwOQ8i84WCM/8oZjUtyFQGWv141xWxYOaLbVqt/KJnV9ZUR1qzuUsrt9pK3A
pfvypzGUo6Gftzfo1XhQFyDaz6N5AjlgPoDvwrBX9/OoKKfgRWO78iDjqUK3wQSR
WAu8ecWKZJcZyJIplrA1PfMpd9XmCYB9Lprm8itNZhbJbf0OzlVEmcfDAfZIkSTo
GjDs8NtLpCMzk1nEzr3AD9S7pQrJFkW+QMD1rxnconNcQmkZKp+xnbCeT/+tdVV8
EGipK5RIPJ6Ry0Wi/pGtvI5s+HJETR8aqOHuWsWAVeSCnSGScOZUpDffVAJeZITb
vDkbBTP5xardKIhIZcnui0krdPtP9lkxIypFfuxaonSTrnfk/QcdH/vwt5Oq597z
OHCnvugOFlywuvyezhkD4wUZDC63P82VaauNVKKAV3FoCGI0woqBj6KPVYIjYyUo
3pYy339Wf/o6ICfKekM48egIdHDAuzWM0g+bSZH8sGQPBToaQAYL2g3KjBtf8nge
1J+lJWG67SRsko8kD9c+5NCqwNqQ4PEfAiWyfPUeaEvimHYLPTIHqfIb+C7ef0m2
cr72uNM+J2LevMsmvHQXGEurDStRfxkJxaWhC0Xuk7RQdR5FdAL6zE/KVHAgtvWv
Ha/P+bq5aJZUssVl/x5jtHFJKT3KHUkPjn5+0s+IWhXLqcCXFPQrwkN65mTk11LL
5tKoMgU8Ln82hdz+pECZTXqriD2xKXxiEcw6qfYyLxVlnqWEOCJ1w+UaYSKMxs2R
z5hxNnwbtndYSdp2nPj9y4nW6EzGjQIK8HRJ0f+bfSjDN1uk1Kjt7NPqT0YC6DHK
gFt8dvMzmRHQhGj1pZLn5Ms8aLnXFMiZW93wE3Lt8QsBPgWMBXEyMJod0Q5HBL3v
XY9L/cAPw4pjIyXzRFAEL3pz554Ql8JuA9P7+MKzT3kdJmAk+iKurMepQGsNJQcp
5igLqw5gaFITfRrYWne8IcrdqSQWVISJj5l1baI6sWhP4ryOUuBqOzaqyxRTmukg
aKN9FnoX1jxbaKMlfF52YOGYoGpQjhO0C7bAROux4M2hliXW948TXO4lfF82BfZB
/cGbg4sFMdlNNb/MaVS+dBLC3OZW9SOVzXmhEViswd+bIeQg9C02ZLXpiqihG0Ub
mwkh/vNhPe/ZyxDewKMw93Kt/ZT4k1CJ49fltvDbW7CuSbpfyPSAkt/+x4HYyUPm
d8cUJs3G4Bg+8Xz4CyCObJVkr5NH3Z6FzVpqazk5Fvb9sb6ruZj1nhpOEWOdl9kJ
VkOWBZNF/vhBwixIaKCRmdWHNfMmifH+aFS28BqjVS8FfNoa/blHU4loss7iPkuh
fUlgROA+3UOoV/RjCEzIvF0sRnCFl6eX88kp86ec21sPDV+f842utHIxCueopnKs
DlRTxfIL736MPvgZ9YHu7oiyff/Ya4BlcOhbV+jG5rga8T0VqOTdkn/6n//MH6io
mhMLmY/wmnbosLTwBCAMUKJIc3inYErPrP7cT1F+UuXmKFYFptfWbc2ZF/MDKH+x
qZzmjglEAwR3f4TP7M4/wA1Fx8lIIB87UMfc0zehFpzk6qaK+cDd/d7crGEFjZpx
joKTsVYmIOpBuUEEjbenpOwmbUYpB32Iili8Udiq+j2stMXVavSNF2jd7gXUKyAG
5MSG3RnDCNas3p2Qq/5cAIyo5ZLONHM1VTAENpo+nyiKrdYSg/CGPQW8sek0o1+B
GjQTQVBxBPdAMagU+bw8rOhOt5UEW8NS/CsgMhj8quBw7NBwv6s0C2Qcwyy+Js+y
76MAmzMt//dVNuhON4eKYdVL5oLCo5rwjfk3qeiQC9CMgrcbC+IKgknuv/5YO0g/
XuQqXH9pW9OerSjDDaQk7SFanvcRa4tDXhR5XyZNg+70H+Dfk7EbZzQF68c/Nb0X
k50kC4c3YHh8oeXwy7eWZV5mpreUs29Jp/VtvDpL/hW1BovqR4pF7y71z8ym6sCg
XzZRY+2pfEQH/9eQLZXIwxJEtXbopuoYL5GZ9PuOfyN6jtDZ1eF+TNMLDUaRBvc3
6LlpYajm/Gwn4yNrHuD/YuQO7l56MCmsl4r6cS6McAvn/1n5fW+9yq/MX1GUr3z0
MIBFXAKNRBRBSopXvhfUzl7GhQ0lpu8stv9iS7P20mZTefsOcRvSDzhcJQCcIA8x
nwFAd3P1jPjMqfaGE+ujUFzBjHr5itgwjiA93NYzAxxHNRE2EoNyaOT6N8SfPm4g
G0BYUT23c0y2L1VCkmduoetA6xS3VzcKsyxwhbqmiMjdRH9o+L6vaS6aeLWFCdYB
b3huyBmCKr1qt5g1nZsqoSnwg1vN8PqL55Dup1lbzs4U0RqZ5FbD/S2ZF8Yc1xUg
ZjNUG3P6gc401jLRkANIybdz91oZGZRGzxRBYD4x+kHAgMkrIJOFzv6hqz5b8gNf
ZN1sDKEfvs2h5tTwAIfsFgkhtRDuUkrqeDT6oUGt00YryzkbaPSlKe8ZQ+BVbQEq
RSPkj4qB6X/ZMKSvDha3TS6wq9GcQOPNrPkOPnkymamXQIZOh4P+GE/9tkR8F+4R
jdWvwiwuedYDBkZQDsxO8Tud5vlvnNfOtrKNKXwXRi++2TPHhPzBe1HBrDbCeSvy
43TPfFevkL51D/x9ReyBudqxCWYDX3Y+pawvldk8wteYialGwTKv70S64QgpcwNJ
Mrpv47sjKPWAocNI3b0lAp7fK5WQC+Dsv6iOyfeXa8oe/HB/ff3zsncZlrP6FTLO
BS5Ze9BXJa/5Xv/0EbJb0YhyZYjpFVf37qVpC0uZzxr0IhV7OUylJK0Glnno6W8k
61r34ZlM20nUJIEqRUBJyiw4u3jpz9dpyWdxtREhCQASj1VcCnfvcgdZVXFxV96e
eFcvv1opZ7YUtDoOJOAGZLw+yHFhVDJMq8dZsNjwtkhSaISTWInOSUVh/sopoxSH
avaosHC6eU8G3Zb1lx/oVZnwcdzyqJylt5kRsmdmYv2VPnOZb+hAlpULgogVr7Vw
URfEfpQfJCjKyhJYHSsM7A7Yk0kLijuU6IGL86n8YS7LSSbTkJHKn1L6lBElxE7K
cBDoa44hRdoLQQNufWTNY5JwDuM1fQpoXEF2vByJNybh/vq6f2t+C2ZwAAeZOyBv
ufxNOj9Irwg9gU4qdrCOURhR7Pyls5GdY8UuVw24SETFwitWrbkn5SGqe44Q1hck
zHp9rMWqW0UfU/ShWnF87kF2ANvNwja4GYmtcYlIqSF60to1TGgyA3ZBSCsEU9g9
2OowzRUxLgrENwfdw4gwHAIAou61KLpFN7TRGaAsRdeQlP/3DEdGy6ZBg3bGYiov
azxaBuUdOsuwsV/aKHzSXKLWAlpYEN4Mbhrtqin4fPeDwT5UvdcGfgiTKGmYwLEq
hueoqtxzG4mSBRfJvAVvJhsv94JujMdQKzuT3PAOpGCJRGSCC/gjf9funDnP5bhK
aUoPTA3PEmfipjTwvvzbVEkZCAwQGwse8P5vUZQ26v85atFASjVrmiQb6jEBi1PH
xW2xkn6odOysY6p1VfTf3+Vsfu3iHFFw1FyJwTls8xpx8nLQlogjF+jyHbtgzXKq
Ct6H8nUJb8cZiKp68hWbbZgH2BvnSf1/A8GwU82LeLOs+5jodckUBWd5hRTSbc8n
RlHAt3MmCiMH9Nw6m6BhcjvIruC1kjhG8NO80HkUOCy0vC71I1TH67a1XNy0Og2X
FspTejlhm5pFZSiZ0pIpDhRbmLXsFx9tsdHmOwjMu8qy/FzdV9/TinoYQ9PVnmSS
cODdUXdrdC38mHuPj+G3115iHQ465r+Jc3R9AVZN1FhwMggw6nZAktm7p3PNWnsz
BmA4G/ZPfy0+UT3ETg6HPBkQhyM1LQLrlloSiXjAiR2B0PDDP+Gb2ZBXOzQmRUoG
nUMy0b06fUlD5TdmMNxmsegSEwTd1W+EzaOe/nXiMsO9fxVwcnoCKs1qStR8j1Yl
CZunC8XlnRNNGAs49CkohAFhjnKEWvzUzUDA7b6XqbRvN+yrTFo7PQ39Z1BT7EaM
cIvYjZt/YGGba9g9AJ8aHvZQXDV1DxC3yaxbPiMeEd+lqL3yPn95GZFbwicTGTyJ
4Xf37u0wilPTwMCc2tUapC5W1M/gT79XPuWBQs+nEFlbLgpFW+iYwZWXFSnWFt+N
zHspVU3cDrs2WJTppWA3RO4eXImtzXw9YHGo18RulTEj+iO9odUaGuLkVJo7qOyU
kpars0HxgI0jOp76TTcO6BmSz7Uc7FImLIg0zu0zpMEM/6v5xH/WmsdFHMZ5oQ8X
f6dRKS3+cAd5gZ+47xxslMX3jPaYNgHjgqntgagSj8cAhzXDEdjWcaxH0b6+ysk5
tMEAWbIVD5lhwK9JmhHeiDICVRKYrNby/URvYyv4dEV7YSpD4vfpzGZzMLtxCnfK
TcD7H5vsEYhXdX8D4lTn+KGL9rotmczCi/RCJtosPh4VJFVS3irjU0Lm1FWK4nDf
Gszqtwu1QL2SiAFnW4O5lfINiCOMtM5+8TcJR/uF4UDYtTBPr2693A+bfUJLwMDV
vwP7jia2NSnTBmPAVbRrPrmtDv1df27qlsgTQy5itmLa0NpSALx5PNwRP2HH69ef
57kIRmUorC6ixFU5eRuhVLc/W0HXNZ//lW8Sp5O7DVDRxDfeXQc9Z4Rl4DjG7Rd8
DYuJJnYp6Ki9G5Eais/44e+hXdBB0t82ULmcTsGv/jf13JTBaOVLjtlDRiMTcAH/
iwSkPPYhFiX4KGCsoc7HhTULUUzyn/dEt/GUl4RerH3Rscwy1E/n/DNrSIB4isTc
/wNsnWh3fphEWzkXItOoQacFe0vbwNSta+dF83a2KirN7kVyxQdT83gudHN+UjlF
6F0T+1nvvH4jzyopjDg7ptZ4lPEINIu0m1tYlLqbFLxONOuWeXjm0HtybFa6d9yF
2himdwtgk9trenldpXSSik/l9Sp+ToaCpOnJrpyQrVdw5Hac5wkCPOsWso4PQ/hm
o75XXSJH2GvZGL9MTvWjhDXP02S1kIAlvz8lWWsw6Bc7oAwxLG6KnO2t5TSZy3Ak
ADDNlSam+nsW771InmVrPNOdv2lYKBDRoou65ecFGhD7ZV7rbBnkaSSnqOErAEAH
lSmhhGXZaEL5rWcemOLUyFELpKb+dQFW7Azuyzy5+yS2hNxiY19XzYJQ94hY2ApN
ro2Nbel2g5dLYDvII7clohIoC3ampWj9zH5Zd+tW6f3g5OqQAbMsnNeEuVbut+7W
Xf7RzWtDScCfmXIKPxRQr64FVqDF2+WaBV4yeFqQo3Blqn+1UEhzpntaiHwAtMvg
QsM+fnJvQZF5nU7TThVsFbBLlyIhjnEUPdQfIQ5935GJbit5kCdyoQ84hRkLPf4m
5plcsn6CPB8wJ4LukuX69Q5CLn63RBQIbaJogjbKp+G+MXLjnzwE/ThSQW5tx+2B
9EaptdkpbO1EYbXLkhXzcRy8hPjSgixNY+jlAiCFClmFqOODgq7hFgAat/YXDnqP
5GEeTKrJdGB8sSXvdy57IaIBRy+EOU5fAPIhBqwQfyNiYy4Fv3zdSS6wKSy2ny2x
vMZtyW4yBjBz7XwEbdxUqoIoBRTi1f7xqViZCXlXdIomE00HvYDgRDgUqCOwX4HL
60SPYwkcC8b4PPNP+2fobluOrXUh7B339t4g1Nvt6WQJojSfbvvRAWggA7dtu+G+
FKN3jl6hv8fry/UpOU4tZGHZBAqLVz+LwY3L3KcGCtir+rJlB06wywR45ljYienr
nnfkpktCmhRZzwlIhH+KUL1iolaHuUXguM0zXLo1N6Wzg86bBm2R5gtb/LV10qod
KVHLvcqTPCivaaefF3r4BbNoH9HuM/kOd3R3DxX0u32UMk41OsiZnPjn2hiVS8OM
U20QS+ATRdqMJHRbYgWo+iRAQ/2JNcUiJyNz0JRvnxR1ILxCenpU0TYmMnvmoZAJ
tecoAfkB3fk+GPNwH7Grw7CBU0CL2gi4cu9pgX5TuQhwExX3HEldkm//ZvpW35dl
6CQJFLuRq723rFvYnGkY34reBNQDBMOr6Q2twV7PDKcZZIybTTY9AvyLmA4qHL9s
vcqmQHYBv6Bk1HCr5tzDXVWUpL4F1etg6AieVND3xswO+0IcbgqEFXUZ1M/viG0C
z6AOyUjG3b6scrZsPp+AjtDmIJyetlr9WHMB9XjLO4MrrvespogiKgTAnJAB9zuj
SQ9kFgSdScML0e5ke+mT/T9qJwgIPSrlmuzXmtN+ks3WaRUs45jnpccHYsbU5k8M
2rz20VrZGstoeanxc9Z3u5o963fP76I904lruKHJrYknFbtXvyoJvdcZ0AB4iAGO
j+tN+SPgPt6m9n+BWyxsl5POwZ5Ib5WwuB/JPxzUozck0xbKyVxtkcSIrv5PQZ8e
G8YWLNiGZt18R29vUP7Kpf6U4JFXmhwJ2sTScJELItCBPOn+A3zaIv07M1sjDusJ
Ej1Y528Vn3TgbOm5AR3Xs57h5zEsQc+wPbfi499a5p5CVcdE2yhvH0p7/i4Q2nWl
QAMGM+tCXRskfraqKshKV2c5wS+XR8dLoQN5fgz/L+WSXKT0tR50MwpJKT0MOk6+
qhkdfe+DsPWmwwSW1k90ULvnpGJHh9y7sNVpKq3ZgUq8AW6mHnsEw4ZY46Pnm+PT
QgJA5Ko2EomqIEL/PIPGuHvl4USFdvCDl7p5to/Qx+vM6YXUJhNpPFjMJlENyIta
CmUtV8yVofGdXBmrZYRPlWS4u8pkl+6rVYjtCxDa3B9RsMlpXl8vwUqr9fUhn7cn
ECqsIR/m8klC5IjQRIJahJnbjKQZ/L4bx2yBG7p7yM5lvDe3EpDDW+JIg8BNSG4j
yYBopBuDbuSGqRUmufNE8gOqkOTDxsLmEPzyhkVVhpD5Mf76lLCPCeFq22kqmLP9
VgvniORycK2SFc8cquDR8/H7OqoONqPZA/1L5F4ZEhWAdqjLnjHq8uihI45hcPMd
nZvm2STtM0coCPbq2sVGs8ElzhGt86nRQR5lxe9sUhutBKJGfmvWrj2K4xeF8/Y3
RgdIBguprfQRvepduJW/by8zixW/bC2KzdQsFSr+HO+Usbl/VeEP0Svu/Qax/5qt
Ghs52i/KwclqCJBGWOKFaH8q6fzyOEnBhYlPIM8ynY5BDpoJkmRjct9tbpLEBAra
lVpn3pPZWMdzE7XG4B7v638s1aeKrmsRjexUpW+fVsdyGGt+hK/A98HauBK1K3xW
LxMwztWw5ONVEUwbmaxoH177PakUZeCBMpUVunYxq+QQWF9SnKzasqzTzdodljzk
G45PfLcLewj6LRq6HanxaRLteUMcQSh5adjH4uxKMtD5U4ifZZIUzyg5pzkCgehF
6kiqkjGdSzhPEkzfquf/peByD3FVnrjp2JcY3ro65sLyQjmuCsqUt+4sHLlVNH71
SjSV/BkDFCNR2Vy5jm73tL//9HUJFEwrYh6eIQM2jQP8AoJTHlDJFU02+G4lDc1e
8r9smU2EbLMharX+tzAJ7UVopS7YdZgkgHsspeOJxvJYHwmSYJ0z8M+NcfkF5SLu
RGglp18WuFAGTvNGQ3SQPE1JalrBCGgcAgslP2roT6K1sBqCa1H7KnZwPKafXfSQ
I3cToWuxg2U5ajqD7opK+SAlUppypeHjYEz0PpcLr+MAPT2g4cx8gGr+C/0T7xnR
3jBaVY8z3hM1qvSaJX8P43AJ/A/5l2if/3mRmYdjrrQsDQia4lS0ihk8zr0eVk2O
oOjscRRBlYGiFr+YIjPsT4xZXQX9JF/lsy4szHATvFAf5zeLCfHqDcNLWF+8SYyg
1gmB9Ox8SQ0HGRMr/IKdfL3nFRq91RentQnofaSMnZ6yPD89jtlS4D3gaK7vZK6B
h6Qd12UVAsxzmJ/8s5oxMkvzNdLQYrco22dVrYae6RIb6kdJlxUbZxdipS6cXEX2
vpOdaDqXp68annp+Cnw9aOPWz2xUwGGQ2rPWaKUKYWbvJSzBuy/pAz3t9cRSPMFv
jI1GXh59qzYK7kRneJOXDIQiFOE3I7xVl+739A52rjRDAqWxjnuk9appgDnwOLi0
Uxg/6WwUTbwtXRkA6GW2y1TZZe2/fxW2+P7kqZocs2k18oFzBzhRYRWxF/9AGtEu
DTwvmMkHB0x/8YYPV6DGRUceok/qqunoPwrlWH5YjTIUASKjJFBFjs4EURRsdJQ3
dR2ITG/tSkNSTTTJF8EPE71NKcK7/Wm78BHQ4LBN8+I5XQaLjbyqAarcEQ0YKlFX
G7kPV4Jyh3Kd7gdwf+7CuS7xgxeGoHr3noDXWfV9oMA9ZWXtYxZSvC+hLpG7CGOc
Luz1gMHWrYXx0O0aoiGmy4vfbGFoFfBmlj/z2wqAiVVNlX4s5PsboA6cCe6sJ95z
XhvguITTyoGIU4JpEOV42GvoGdpDn2JH/n2i+uRtygMuT4Y7WDhgtHOGgfB29o+I
5vzoDzp0Qj+LgdO8uVaDV6f574hMPhvxzw5eGTMXt+sALfXBo9eSytRgDjozjRb1
IHH9daG8nasSB1TLXpCjtYUVUAoDYBZ0NQDaT0EORxTQxR5d4NJVuwgJIoZ/KjGc
ennE0sTIxoXWyMLDBxZRBth5fEIOnoEABwVZlAJdMiCcMLS7gFxz9o6AbPUxPVoh
ECtElP7u/fQsspXGUDEZCU0R/HKHO3gaSNLxQv6UMdF+k0G9iZkbdJUN/r69TOdD
pCUJPuzHO3NHqeZ9SgIJ38Ho37yWCH5wO8zfSF7iV4CDVfCaPdqIPwVTgu7UYe3c
zb/uZRuYQkNk1XmHSl0zmau0VPKOsc8TVO/JXjoFgWOSZiw0GL3IKbHfB0kEI8/l
VdYdHEmUE8lRY/Q5uIsddluOpJlP5LhlmhkI5sFWURy/bRnLVEnsLXnoVzqqM8jd
wD5OurHCQwsuP5uTt2/u89r+wVNRdt0XJ0WBnhLGCEg7mEVsNiOgluUcMEocnZPf
Ypg5HaaBHeOHTwglUkFiGap2BFlQf2YAEC5PIPkO+TEGzHdY5ntPSYWKcIfED5BB
6eodPG6MNiWOuPQPN/flKb5uF4QIEeogTQ+q7YHHxvg+C09g16lgHbn4t8vsK3y0
DZMOhzo4x3ScqBL8O6NvIyjrrYqkuYHN03PpcSM57+wLIISaxP263163yjxh48ry
74lU+Jz5aejSwPhY7QIzSCOSlV1H1trvwnRBrH/NepozCG4ZI9cibzvLhmZnyWfM
LbI90LNxSBDtO7sbxJV6Jx/sIvkwgKImTM05Ka3E+cdh38QHZqVt8G5gGjINQ/MV
P75Op+a0h/+pQ0GZq25uOmJ+N0h3DJftnttGNLyvU3tIpHDTdEXJ7s0SG8+T8Yn0
5Zv5XZy5N5mTZ2pEyumI9ZCt0sRZPpzcQ1a4MdxllUgK938GaHTRS1Ww9PiPB1Ng
q1UDAcXDN3cPwZCix7/pxY+Tt/v21ePluhUgxAOPbC0yNrHkRPpMvvh4j2ctro1I
R06iMQhzWDajUHsQOcXzZ7ngIEpVFNTRCIJ+G++4iqlo+FAwNjKf5/gD9mGXsPI5
Aq1/1JePd3Xj9H2or3mROUp7VF/Qb/aG0NO2g6gmdJjZhpZauOT03T8e6aWpHZqy
6s/EEZvH3m7Lt2qokMjyGvIsKSJdaCflF3T9koQl/QiMA3GHmid6aofJYTPeHH3H
TjLV8zqHq5E+KIWGgX9c2x53yWHAtmKddiTCT8JWCRRFO0LaTFEow3QpRnis0zHp
YIBtr+XMKryQ1PsmDR/8wlMqzcEl3u7sWLoj1RV4ZrC7VWaAY7aWOvIllN9dgpW4
/BAsxCO7evprjEQ1c4/aGvahUggQyWIQ2EaoXHV+oHk6tIXhQWMZhgYFuqVB9Cnw
eFAuK14mc9QD75lUFuJ0d0sHGr55uF0MNa+l6JfE7S4xCHLyO3oUcRFTR6oBI2bn
MJcAle/GIxB6/m9uZPwGxXMCdvl4xF77JMQcFQoa2KqHN4yXMozBT3OJM//vSsj1
CxRSfdQDh04qMdJwgE5AnkbczvzGgecOyzsOxOW+uLrzvRAC2Y+RnONGTZrPG8d8
+YXgtLP2pYV3jU5m1EZzw3yAJIkoD8pROFo+q97XUXkGcqiAa9nt/ZwpsIMp1vNs
aG+7xP8A6QcaNa/TqIpHfb/TFZnLXCU3coQFq49ia1iMs8M6yE8HbdOvANCrg47g
efgrROJXSsda7/HR5H0s5AM4IRzqdvK5eZM9BcAf6mHArj+YnJ8KhUq/ti3yyLJe
JLLaaJ1CaPNgB9q45eWUrceedphCwIvZg5ufU2WN94EbWLXdszwWxaF/IdKSB2kN
6b4U7VFX3Bl2NRmWD6eR6YZpIcy4h5Vu4JGiOqi7l+/fUp6JNfuaXG+TPsPrxtrM
boh92Dk+tt5KT6myiVEcj4gPIPk2b6MhoyY1DCX5g2X9xReCfm4Ltzl2VDwkR1e9
hLL4zwghEM8x1CgtPB2+93pShA3Ei232m8LVJIY/u8VaiZXuh24m3gCChrR1oF+m
3lU9+TMu79f/EjH0LKfFDto1GfeWRSs+MLbE1RK/wbNhaXcmmpGqM2sKsuLLqUm9
AQiOthqLxSGCprTWv7NxkcNXnZZXsj7/GCcH2nqaVO6R3c12Fy+jnLd7jCWeNUGK
og0ndGWbECiYSd3hAuZQcA0IWeTFaxBLkLrZ/IYpFRDKjFC4v5lPs9Mil8hU/XVD
WS6CW0hKaD0HtHYEQGMksdwD/wK105P7iJGB7gzX10dCz241Sx39JwbmRjY1dwwE
ahqCVE0WOZfWj3WnBHhlKllWANpiDaxnQBNvb+SWRdsfZYALYPNDaSBLWwZNukG8
U8EbVOml3uavegHf4tvW7eUyla2xW98+A5j3tXVVgse/0m1W+u2pLl6j9RZXa0uX
3SIo012+Mgd7OsuMkNuhX+Ox2GZobUMkGTEh+A4TWdCWkm3zJ0wye9RYSBTNpO9G
alRDvfuuPEw014eZ5Fkw1V+xXfQbAusv8y2pUleFGQdSp92c3Z8WMvSYUCeL1we2
M6lEyMBTMTAe6xa3N1HeKzOXE8bXpHDQu3P7u2nOW7d2XCLamoujUEM3INkvdQjN
vHCKb2Lh2NjnH2UthwJYx588zZrvu9d3/O0D/Ud7QV5ImDpGriW7XAQUUUKL/7+9
UAtpndZyEGt0npeH/gec1tfMgAcX7zXobra83pHmFeNU93Ftqoy6zr9nNhvFIqeA
6BF3YNzNBB55/HqK7e9OO6j3CQuEpyAuo1PCUflGrwoWvh00myCuUtPDJDnyyXS1
Y3DuHvGWAv20JSE21wwKKI8sF1VDdPa+iMJ5NnBppDlaUUAOpzgj/PQT++rC5OnL
YHXuNWAnbAZSQJppElW0KXoqBVYu2qYnzTXnu6KOk5KcVbEM6Gy/p+Cvot8Pha5a
cBQpbJ5RPqb+A6XWMmuzWoSyBhWvboQ7wGakuh8ShHaGUBEWcl8tSoum1D/qkzlN
iyPpkGnqiuZD6WA97sEaMIApC7tvlfTZwQcNPjyDFkTal54Igy6Zp4YpAUR0nf2L
qzlLvAn5rAEFGUPH+hSwa9o83HGLhWcgKoVAMQcVotRJeKUublCjd3AxvAzOe3xE
NPaNTWOQ35Jll9VTNlOYxQYhwF7ZHqFz95prBd0pDyOUmr/OYI44dJu1PYdZ3Xu2
Y4PLl/g+eOWdET7YEAec54cjtKOUcHIQSF3fKBt+UfG4G9XfiCoXFknGl3+b0bQU
izsz6oDDXCHhvAPgFl2hCxT3ENh7QcbnlTH3jru1qtjf8UXn+Yj/27L7hjVEISmm
NIVF6oVnKvDrqhwDh0Whx5uLL3kw6h6Z88uqoK/if0WkKW6ZZOvLC3trfhNmR4xP
ryh2MvxWIMWCxpoG/UF8Rgp8KBeSE7bDBGoLj5oWUddqNaEH8sMZ6ujEkmxJUHMr
qod7JQScRs0XPBx66/Uul3dHpbyHupsePAIlNgBNd0dwJtbBfm/IIk1QdYPxrn1c
NRKqCZf+M5aAGhkPZ73mgK2c4qDJz4vHT+562zO64KKJfNv9hiVlunMHD11/cQSX
dWPrtRMpXP8p4ocR3GhStRwAJwe7wkr1rsAm0qEgO8bDY5q3+NQISzG8zsZ98rxB
iDwdxUkRE9xwWkHi7I/UNVe8w9kje3EkGUmBw9IM80tQcwXRHfCwWVWMpkRtOqMu
UU76WvtJXQL478SgXulCGlu3AmjhAyYxHu7JpKyrhlgM1yHTkIhLz1dusxBbLZ/X
zfxDSr74PxOzlbLimIMhpFCKaiV9jxeQqzTpUW8BvNHm8ZRFBMoRUQgz42ViUYxp
JAIzRZVAv1VxHklaOP4Hnaiu3msX56bGH747yxlab37ja1Zz7pTzyPE/XP65Tkpy
Vq6Lbp0aiJJFYpLOpQzXl2rEar8S43lKwKHKpdZbQXvDwRMwknAuy4o8Whth8k+Z
2X7BKQ8/dydI8VQcdmC+3nEc9I2aHXuOagNfCSzkxT8tz/JgeAJXWI3jdpqrzgv2
eV/1AOncnkVCq5IJR5zdrvQoQTXDLlPG0qq97ZB1Pa+pMTFeDYao8VfBymqpEh66
yytpQGmZseUvJ32irMQ7Q3+WLiixmTKR+X5RmA+RELiQ8nVCZ5Cf7XpUxhrAs+ur
z+US2fxp8sIxZ+gZfoydnA8s0k0j0RMiv8uvyETrwt/3f9Gpo2ZPPU+rW/ha0OdJ
dfrAifoJZrxnVrz+4HwW3QrXZ32QUl9SzMmq+uLYGf11QIpzI1gEaqHhNcaZMkLA
VIe/80jeRCAcGFAqOdff2XGlmMyBrHCU+RdeMcbRcDYvkjU+Pbyz5+f4V6NNPSY0
0gzIAxkqg+zfu1v/Qds11wZET7VYVdAVHpJouNA7t0Lsuvu5cOZFXw6J5X3B/FBO
dyxUleq66FvpnQTtCuERWlsvirM5m+JdFPIHLVeqGugSjKZG0ew/pJucXrk6hOID
roRlERWfq1dgm0KExX6eiuyRYICkG6KxWOYMhfI9KfJUYOdl1d70YAZccu/dJhiE
my9FywesmABGaAA+IJ79QqoDHepgyAwyL2NpTo5peWM6PbCxHTt/CFFMO+9CiPAf
rkerkopkqvtv6thF/Y1cx6pcTCPmA2n7iC73uLjXG17O4DYwN6kt2+Fw+hDsYNl9
VB8fes5I1C4MgbUxxL8enSlleunVTSAu61NdP1rkpN/UBwA2DPWJFVTEApJxui1q
zZmoEkM23r0u3TFPD1b8u1ekECxrPSm7XXuVccX+ZX+9QzYwwvwKXmCZ4sxwvpFW
iS8/zQ7q39wKX1zZVwhdQyxDjladNTVJydYdPPqtEnclBfdB9Umxn8+/jgnfwniH
5gtPgv6wFhcSusDKdLZHT7ptYaAtYXfpxxy7r6Mq5s7rra0MsgepfRiFbQACEf8n
PUbfWZAwVIZV9xdzVvzDkV/c9THw3qPwFdincH2riGNmKFOEhfnJlVKmhjrTmDaR
2ZE59EI6GOwDa3Hcy6xubZLwYULPvIrCeJ9wcH5Qcg3R+YDqbKi+z3WzrhX+9Tlk
SScDF2QayH3sexZR13Cw9Zxh18L5dHNdSFhhlzpClPRL7huCHXqHBl4JZB7OjiPX
5FPJfwJSIoE6Hv3QaUKshhUvnchOLIT8EZLHoHiYhVBwXkLLJeodbE2xCqHyn+jX
6MeVjbd2z7hTSBhQtl5Fq6EvxIoaDbsuJ0HMaH4idBV57vI3+Qdd8D34/G3hWKZL
/n0HfwygIOpUYEULJy3w5Htka1PULWtGjp1FyJt+f4WSJ0NAnq8p7Z9NhZsiojnD
KKrnOGQSZf6+Zh+UWYPb8kSDo54x4IoK46d+PPS4RIc/TJj5uK6m+J3pOHdlU4Sp
gl3jASmpjTR69yaGDwuo3hFkkhRm5d9HencUMm62lwL3d+CeXORgdsAV4oRrEfeh
U1z2+0Wl9asHSqf3g2yiUEXEFBmbTGuTHScVhusKUC6isZ72Lr0dyJRaSP6cxxTh
t4DqjK6FdYMrzxh8lQc6EKCQRewie1raku66L/VNq9av2G13r2GF3l2Qb6g+Al6R
c4R3rG/MELdxz+nx3kezCAWfXEYFlEsEcx9pwwGfHqAt5hK8hs0VzqatbLxW/mR1
BYDMMpk5/nrHt387pqIc0w17u3L7BI19f8Z4KtPi6/FtdM959R7ejZYb8wlNV2m7
XH/HDEPBh1gpR+r/m8jV3GZHPEuDu3tXKf3yQztNgCsoONR7uqOibQdhFmolu8hO
7K8ieK7EP1vrcgKjOc+GPpWZLq1K3NygtCsKhyQ9MXiFrZ+/Fc0Hhkw3TAtp1CY+
fN0xkmz0wolBDbnFPP/v+t0ZgLxhsRL9tz48vdNb9AW7UIXaY3VHlQTE4kQtGmXe
Ndfpu83ClBhYRUZ/L9JtKm7Rg3+2RSQLU7WJkkF12iX0yNxGycWLNzj2oTWbquiV
QWZHG96OcgEHNL26CcOq4TwiZ2yGYwjLCFDCEOCdCVwJ8pJlHISAHs8+LPH5Ye4B
xqvNiclggRIznQDZVapV0PFT36taZoCsGuDdqM9M4eQhc11utLDStKG24Txx4pRb
5KXTy6t573eJlCCmmUIbk8Xg7AlTqrYG9w4EQXk/T4b272h6RFIDH/n3d5Lxkl+y
3VU5hGSWUI0QsucJYmPKSGuLLeXNViFBqcvREcQpVd+QhOnB7WKo1gW15166Pc3b
kaJUwgbDLMnUj37bCTUZWBYztro0dRfsTAKT0yx+04MA/ETv7qmFn5NbHbYkoVlx
ehDQXHJ7CQyeUdlGofKT7jl9N8vId8KnCRdW/L/nKN+T+0WcBmLvd9Jb9oV0uobw
THfrolmgMDV7IkIlywt8BqVc/t7K9B3vKFVtsMEp2VqLsk0nx7CiYJHlIv6x1Lgd
cA5uvWU/dKDB6i+BxTctfcw9vUpGO2I09eeqoUUNnboroLsGECaEJ+VOOXY0viOb
6kL49SKoV0L//8VoxhrjmZLpx8tJr8e4Y68tZMV1b9iCWuzA8nqZuelCyYvjJGav
0TORRo0pXM7DuOX9lZ4eGhnOuBVL1qCpGusTHBAHILvoQwSBFacCBFQt0pcurKey
xRsUS+mHlxx0nBcCiT6bLWxd0KFFzrxdZifkSlhohmlMMzh4EyFwlsOi0k8eKGbD
tLaXOqKL6pLSkPxJI3PaNrUk5+zMATdvenjGzj5pkZeSP2BSXT/GUADTSDRwdtX/
fS1sLQqm/cyY3mux3S2Jev3VQrT7wdxZR6JGcxodf9Sk1y3AHAzCqh/LSRi4bWKv
RMc5M4wZimsnFy6KmRXNNAC4ut7bgjJb2R8go1WS99A4fch3KsvBuLf+PP/deUMo
ilzqMZgcnvNu2zMF7yR3TDWWVyuuV3EWA4BW7kQYd0hD0whMD3zKvow1n+fA7E4c
F7Hu9SNQfhjHpDjLZfjg3SezxbbDPIc9T/v6hMVfAEF7ToLzDzte4fH6VNSOc2ju
qQH6S6UBs1akw6mI+YRacKtxoJLcep4UWCPt8DoCllgqnhxSQ5FeTGey/oShmblL
BDm0HAhbsjR/93rPZZU62jUWj//2wOziUfStBHKKkbNeDnIrU4yyilMBdWYRhiaA
dbMNcuAc/HzTsRdQqsmK0Ubnt9UnPBlx++TFhMLEq3FDGFJEZfZDoTZg+YtcQh9B
qTcDR60qm2GWVN+M0qBrQHL8Wmmhtvx3UuEMuCDC7ZQXXbjybhScDQClpbcAF2bM
O5LbxkG+tjf4U5lZgUWY5RnqZ6j7JoWZk6Y6g7Ej1dZxGX2o4bRgPjf4tpMNuiZv
7t+xFGkq9v2LZElpzndpqbiynhg+wQg4j/7bgHGafnQFsqH2AEMQCG+FiSK4S2ms
T0tXPi49jFbsmTF3iIk7s/mCM9HNMzUEFCcZeCQdwZVfRy6GVhr39H2hgbXztd8y
wJg5y/hC2mYs+9g3vibNXn0KF8Ryd/OOGfbPM73aRyvXaR+8yzSxdZxrBuX0HTFd
qQ4oaCH11h9RKl9/CvYsVUGyDFhyEVpsEHhbNcGrdtJcimWdu5me3cjLWzUiAqtk
CbvM8riqRvFx4muPjf1LKWja9iCBC2LctSL3RM22JmugvrYJpdjTeMa3y26WxklB
QhTC3YHLuBCGfAnvaFoaewWd06QSi+/zom9o27j04WVdBWa1MgxVIWnsI2egb+M/
/fiexfFHtUBPNaoOhkfCu5Mbxo4WPcTcETSkUa2/nW5+9CbxSKmMvdACW6V8+P/Y
bG0+alm1QYeKyJqj6iD3BBwcYY959QSDhFJ7u0bBsXDf03+z5a0LFHJw2Bg+XQf5
C14o/f1Ck9/NHLdDGZPfJhIKiV0ummAZFaM20zVV0Gi41yDVYiAMdSq7PIIiCdX7
MzeulNFDf4LXk3DIvnY0RDwuADVpEVieZIQMHEcg2uh0TUm2UZC0ifTfrs58mWwx
2nBjPtLUk3N+ToYscwDNN5ElByk8aOaY/gA4DPb+aMd5hlrtPdqjnZ7tl72npXQP
xy4zHjODJJNb9GfsULeWBbWUs6V2G6olSJVXIDEcTME5XgWJsjOo7VXYrAtxntFj
mRvFhE+QGK6aaDaSg6Zsm88oWcUhp1uKTUXlRAdw0Pj+KNGxHmH43KVz/jURi080
/ciFxwekro89myEzC3W/yWSEYwdtjwJ85kZWPWT3zehEhfXh7c26sbSZEjlFs4eK
u1oY1XU3wSykz2E/+8m1R9yBDRxJ3y5CvI18Om80XN1ejif9dx/Cv14dbvnR9RGE
iycklgGHpAQTMPveD7Ed2+YzOpPg8DzesfjwMxxend9vVMEbecTFdT3olFrC58A0
FdfClBi/IcFDjPVLRLOQawJyRBZXg6IA4w+G88/H83qW0+wfvXS2GGqLO1uzO1EP
J8Sr09+h1rvJ5vNMsyYg7pqw4uLAdlyzTHUZN72VNRijx/Ls4kxs+RXVnmnxvgVo
S3v2W1j6PVyhNcWXTLoixGqOapAulAOdZ0lf1ZgyKTV7HLi5SJj4xP93uDdFv2B5
gmHYADK1/qEP4EV1LG1joOxPSUU7aBzbXmTuSQfXCEQ0zBO7cy1QOawHaazd8VFD
SWPPfm5EoXYAOrr44pPkFK2liworXer187KS2ZGyPPv7pwI1rdGdc1jDVH8nNfDW
/Acu7ToVMOHzUCD/nuCEPv0rg5Np3BhlsPrCvg85mLHGFEuC2kQDn37BbcMQFKxI
qTxlYt95EMna8lMTbuBG7C84uRRFxF2gmmLnQtdf8DgsKBde771d/uDNZas5LYZy
TzXT/P4APwDJvkcQqmcQW8Tu0+sivLgD70g0besr+6PIR/Lnkm8iraQA0Ak58Jfb
ALBn93rNFFJ4oJtWPXutFymL01y0rd7uqSqofsmBPEilMINOFzDkrd0TvAasc3Hb
H+29O9eei6AGWSvgS21PL8ZSCiwR4eH+TgOjmenbYBEibO0hBRsi69JIC8P0Kbx0
STpRl7f4+ojO7YGQvfkHNYIPZDEjvWT1jxL2q62hhXGejcxSHkODPMNXvp1e01gL
pTNSaWID+9xBrE80U3UrD7zXFRpqKxRRLJUp93aYYGxJXQOH7wSuvVAh3iYhONvJ
8vYETgsqT2k8qeGU3IG3eEgnThHKdoMw1U5YLrZ/NG3K++ZUYXeFyM51OA6hMUeP
OBGzkVp3MlXD5i/wxaRurRwT1x15ibbY7hgwykY1/9W/+HBWzv+bJaSn2bjHghjE
qEgozqMNyCeeI3jkwf6EjZYEw+OwywYhLKpX8kwxvxPCdDPeY0BB6OypEdD5BB4O
i2OzxJ6dDS+IH8NvISPW11Gif68PHOidARoGMfhRmzaQ6RzJeU6QZ7N+iBmlE2mM
l0WBXDykmgDYz4TanW4zhuwwIJl+fzG0MPczb5oqRCefivCQVcSdiXiw2ofFSRNP
UcxFA5cDVolvd5Qz3fHaUZdo7q08IkgEbjJUHOjSS3hF+f/PY8lMXPefRvKcEkR5
/fuTnU8/deku24BCeu5scrugduaoobMuQueVgFUE2nzfdgub1w3wXeyZLjZ6EJp4
neYAFUQYNcWBJ0anzoWP/kxq7MLu5009OfWiInd4gWnJQ2koy9b4ObcMdSaJ8soY
W5xpPjxWnw/zpvO2p1ca9Rmseb/U2CyZGqFg7Ukd9FGJ+RCaS6Fsaib3bSr96aQf
ZAl/RmAJGDmZkBsg63xienS3TV3pzR/bp5cPz8IADebeNX5O38LPjNt+C2KAifDU
ALL2JDI8e405YqleDIBJUQcyWvthY6mWW2yLScuio1vL6ZhRduV8bjGwtxmfDIIL
t+h5kKkjRBbB+inLNmUsc+5AR3rXWxIxEgv+KAdz0tJcIs+9qlTwmojgEBArZnOW
90R+OW4+G3jEet8+p+IirzTaYJ3gYaFY5VNpykQ5Xt+319EVCYI7yIKMCcj1QYGk
uttJ76/eQ5vOPa6f/uFjesYKDJ1z0sAflUg84R3DbxESdbDR/SduBP1Ahd1Dsr/P
zl++FuRJKBcoxXg+HhbamQ9Rra1k6zT8NFSUJr/a5Xa6R4aEiah9ssuBMhM+dFXG
IkLxLTUOM1RXYxdXgFEW7tTgvAtv6j4LHOTgqOyqKT3D5rxsDMoqpmUIWRRLuazb
tp5VBuHLt1i1kXl1KuN1VFAiiptc+Xt/wft4ebnb1kr2LGG0bFDvNX20/+vcPbo6
EebMw7tDQAF9aMMbtTIbxAZ8Pfqii1PAlKWizITla6D3FNOk6DDYN33DPtC9j3f6
Kuy/53HBw4R0n1u4Hg99PkE0MgOm0wAvhN6gYRelb3aT01Ooj6wxUa8VJg4AXNL8
BNMCc86DtDz0104MFeWrwKXd51DGj53AsJ66wvkuikWyRMFm2XBpdo/4TS+VmKgh
Afp4utdypOz9dWX91WwLe6UTxRuKzMSVh6bxGbYe5rPBQuImiGjxN7CE/ZeqBbU6
d3e+LRuT/iLgorOisnRbky51/C04FPxyJ318ZHqNxASxE77dBviSts05xV5gCH5i
zmDKFgEgtMtJ/3IP3AYISywzqj+153GjVsTdLRx6mnP/XvfFmkgSUGQYR7vvknpl
0JYxNv1AjoucKd/I/5HkuiU6VFZbc6+lBkfpReDjXsSuVpXWRPHQ9uwZqD0/hPbl
+FFLa7yqIb6hb5Ht8vaNi9CkSxtRu3pnVJjXvcXtU4uvEBHwVmH/tjeVYu1s1+Eo
xB9MAjwFyoyZt+eRAKVYs2cPy2fGVXcsHzaqCgfaG8yPV0kNc9mCHjSuRQ59NM5f
5AxY9LtK7CVBEaij8vofUBf6vq/b6BsW9/sIVWCy0/Fx/qVI0GWJ+dPRA3Xr00sp
qDHqIutkZbG9NfbdeocGUGdzzVwNP4B1KbGyvOLa7WJCVLy1pOLhqUTiAcdzWaf3
G/Iv2kQRZwuWEu7hJBw2Iw4vs0m5QknUYiI5i4pD3hZdPRc9E2NLhLN5+kGLUeUk
tQEsPTVM1/DwiOqaJS+oetx4XJ6A/aOoWiJB4oBABrqs8gflQb82fgZl77XV4vTf
Nd2nN2bZFbXQ8Sx7seU4tiA07ZHNKmi4Ye0a8wzXkgMLp20V0Mzi1FtzHRwtot8j
tzhIfz9WefTAppXixOT1L2lllQSE3D5Pz6CEnaHukuKlEuEzRHczeE1x3fD7xa1g
t8VwHcfXqfdsEeFMfQfOKXkFtVH9IRSp5bZubIDcaW80SIH+l8y3iy/fsJr89XRu
eFE3tc+tMiUH3kgPgmpRpXDPTk3XTnn2EicYSlo34YiuiuHcV5IMhJv2LZ9YSos9
zFF7/7gY4GiHSDHX0zeZGENiv1zvGF7YJQH4DIh1VvkJXr2ZppBDXVIRDdvH/16Z
9ujDFdsOXbOb9l/ai4HiZaarAkaY9UN9LeZsNX0pto1sDjVjWWrr+D2gvmBr6kvg
aYljc/g/4tJXg3zSb+6Uc6yltnlbUVIs9+SdJP3SCR/1+iypMB4GcusP18uL0zog
VYMfkxBbw3miHuZWPjjR6meIHARWzIl0JGp91Fal9fO3lBFo8bH++/2Odyi+jTVm
17x8LbIRD3gLukmp2D6rqYfs9krK4dGdstG+oTYHwlDBRGx+ATfrYnN2QPY/mIo2
ZvbHKecvY4rInq17/SMeWqrYFpMfATOrf9FOZDeP4BDTaQ2opWkoW3PQHczJ2Crd
4Mwd30jBf+BS8QZqB7DWzR8j1cGcnl+BG1eHiL3PtHsK9w0IqCivb9X36g1ngIvC
WmfeEm1Rf0BPFDWwR67HS99zMsB8CnbINMIlQ/6RK3KYj2JqINVcXnLptAnHd+Y3
RUQLb48usBr3+TBYbpS48RbNy2zAA2e4g7aE8VQWsJJfpmclbz7hAu0tGqw+K2es
BqYwqN06lU4itGgalXXJdMVrWsI15hnbKPKLARVg/RbRjdqpwx6OGkLXvqb2j6ju
IOYFkaCvSFOd4ibLNnziqjTLRFBfOO67cuskb3nePvuzb2mfK10/ldjjL3GTw9mV
7jl0xjUA6O8X1CATtYSGqVD6GC+6HOgrTepTo1tYZTM4xRvtHPAk1C85UnIPI+4e
Fe6A3kKxlVfW9fSmcwde/5Bh3kKgpDjEjMoPdqt9jsS+oUjV9vsZ8RTedqZ4CzQG
ZiuN95S1iF20EBeIGBL0b1DNSwLTb//g1khVmVIqtaOhWhbeLq61honCfcEdyPO8
qQpM0VR3HopI2TJQjAdKNEGVoCk45DXxUnu8GHSSN3x8tDLOMTcbx6VyxKaj1myB
nDHdyT3ZgNx5CGemXNRZZmeBdlvDDJ2lyLbb0cGh3KymJJ6ylBuxODfCS6EFAodd
nq+wTIHGOcpDh6fvjleJ++dZKanBstu2+Rk18ZsLfEGqs/wOExjBJkVDjPY9H3M2
nS+deBF8i3mjj+cZTY+j7tzLFvvzqxLxUdDO0PeM6wRrOMHu6Fy/Vqed1rUhT1nO
bDjKBEcVE5T5xaTGpH5e+4od9dWIFH3n8ggGkyP01orketRVn8tgRD1K33GdU6PV
AphtNEPjxnwrnnJe9u1MUXmichKBdPYaiwlu920iJUDxA8GEKv+bmuqcbIsKcm8M
648WhD51ZfnDYdnjy3Qdq3w7yUxW17WlSG5qMTDPaAp4rSmkyf763lmNl9aVtw5n
MWlaMyOx6Ymx/0Nf3EDDT7Z4GJswUSZqv0VmfbC9CsgVE9J/XX8k13jw1iFhL7xa
Me0OYHgK3RjrLmYisjKEJZ7qAGE4Ehh8jmTeVELo27hfq+q4Jf1WyInejxLe6BK7
DIOyW2BtFj/l+j0MgaJYRiSSmPu1DxGORE6+IJQWI4oZmCaB36JzzcB05U8gYhLS
SVEDkss1/P7tx6fXJp3wjfm1X+H/RtpsM8+mLP0QYI/reln91GjA7Swh2MxAnHoi
yXDOVEyMpTociRWjG/P7XQCXrsqVs14JliNu1WMtGN7g4mt3vd7HH/OvpWABuuPw
qxSYQPT9PVBMxb5Kus1H2YGGTV/gsDVoiWMztSuOHxh5xW4QLRfcy2u/3SbMGSF2
S/jzsx96zxHQ0bQl6PxIF4WGBALp1d8ou9Kv49Z8iA6o7YgWN3/v8NgUyUuX83dG
3kXHdjGY8bE9kJ6hWM+jQv83dH1lp2QePEaQ3Tz/PaIa9vPvds5g7pyfJGDG0Xd+
8XA4UEulvl365QnOLJojEjtZMZFgaHw+ycUYTikOaPCQqzvP2O7Lp0ZYwTV2c1In
PbvBQInHR5jRgVM9fe2iRpnuiYqZcD+8uIYDF0I2YF8kmqc2x6xaTD6uphcj6QFT
dBnCdiWL3CigOC7CaCIo83a1sc8IOW0uEopJ78IHV2b2pG+v7LS/Djeq3EZsDRh8
pUl0x/qxBM0xdg2UrEuicYCrS6PAAjc8YsjBoiqbJ+n6xLSDh+X7uSizY4IMRVX8
LuUSIi8N5Z5sihRJl0WinDvcZWVWa7LkXq84PGH64P1s2+tPHtftHHUzwrqeYdhE
9VloLFqGDT+GzlrW9NsaNzdFqO3fZJnnLknJtLEXtKfh0OA/E5dGzUxi/FhnjryN
ZdXUqnCplh+PBT+g/kKHxq9/c19JQn9OnUq3KV/0JdsTELRr0btiOnFY9xMdNUR4
0y1MuX7kK1gpxmm61ek5Mo+oNVw7Gra0y+8Wz55UkNCzAAN8gaUi6CA0Bef8z6HN
oeUhoMV2qyr10wInUOqTJv2IH11UAecRFQYwOQh2ztAQn/Whv+SeMwrEeWvJfRfQ
caz0dwRHlsH6ntq14JUMTtHajutkitos2aVVa4ST37hslap+4h2ievFLRL3Z1NPc
SRRmmYTTaZrXxr2g408cJnwhQcCap4SPAepKHn45cMgDP5inZYndRENzUyDfoR9F
3+chPb7bboQSYRQC+lYX8UfU0DJttbid30VQABpq4qvcj2bLHtJE+69IFm0L+9eC
NTnn2/9CtEQVp0OS2QRyrxMxoNlZ1r5FtHThtWM9m45MrlZukSlic6JBaeNbI/YI
FSyCizAMBxZcwEm8csLU2iVWJeMh9JUBR9/czquUVma8mA9XLjqHAV6ppUTQie2j
Y53v9pf7WaWDpbNwvd5UvhXDYRvwq+2JVacnd3OifRRN/oKoS0evt7oyhfAjnmpM
1o0+UWi9Ev66+nRjWU68OYHFuZpJMDViAuhaNXMPoxSC/jLkY+scxSah3wJYawp2
pTjJ8mnrD8+dDP5ElMLR7o9pZ1yt3u8dbJ2vd4pKoRg0sLKzAC/maRrSEM95QEpi
HYbQPSnoLosuWNNSgkOzFc9PvzF4gPevhyU0NgUMUoZ7Rp/Qdd6Aa1u8h7UxvS9X
6j3TIX6/w+IK79B7TybNMf4DFHpFzcO1tSlp3c4udmGlld7z6iE16RNU73MkV4KH
M9N6KgxdtsX0WWZYpb5svNLRVm1L23iFdbM8dfXE2LpcCi72ouYOQvoRqIiiFzhq
K8EKXs3dzr5xGqxuHyvMJgCeAsSx1d3ZfFlQVfv8NNHICkVqWRAJzP8n/fFI1sWk
HuLnTVMleum2ycvMmnPs7bJlmi1b6vqrxwVh9TgZD5azeQxq9BtShwkpyh6QuhYj
lhthEzD6cS249wH4AsElY943H6sgcFmOhcQsYjvQazmNlhnHE9ZY7jMJbkKbnfRL
9pj7JuBdHDn6bycwHNMikiXBnY3TrIET90h+6dXv40EBa1f56coUXUtc59G5O/xF
t/1sCM7QgI1iWxMwGmPcVT8JGVnEu1b3xx8LySDjo1l9feVELB1NhSb65GCLO4RC
ALIbr8gYvC76oMlh/HKBUt2HKi3/xfLD+T4s32wKVXj7h+2ASr2mt22y6C5PhB5s
uBU1N5VmEfOmlZLj0dBFPhlvrZ6JY5AYOK+3Z/POX0CoiX2nV/9bsJA2eWkiPSyK
V6Gmz1LHk9ER1UsyKOBUV9UytXqjm77b6LGXjFtNa4m7sHCbbYEeE2K1+OTiKW+K
nfkPR7sDH2ZRFnIn+oJd5DvA/JikL1bgA4Rv7G6S+YIq+okFB4IuJSyL2HMMWl5/
HKqW6tz+nBxl+mdSCIosLdnZfzNHuENZA8pS2kHNfNJAeWOY0U4ffkkeHkvtBdhX
RCNcY+vQakhalIkYaDkErkCax7/x9rgf3clu5gFDO4deHi4juuk2e2NDxrNYYWPl
1QcJ2ADST9XgQ3FxKAEY8EKMNKpQbe3FRc5E+fDy6Cvq+q7kdZBCxb+p30ozHjKY
67o0H98H6G3b78UtHp3RepLECrEgW/MbGT1h1WayAH6khLvVMSrTDRbhRblCzJ5i
pu0refn8IrIpLptlQ/pCcuytKR5MjFsuycIVuRfVwM+Y5GHd3pGZoXT2KvM772Ha
e2HBiIRgRKbU/hO7THnCjtA4r3lt1vrzmNiEvOCBRMYqMWTudtoTjMLm1P1xYxiD
F+sob2nikXTzr8jUIrfMP0+dvNww02D6iLZyL2W/DYrFLBVSF4Uq/67skcZCq0ud
L3drJJt4+kUA0iwFIM9GI/5Ujczck+xxWPd7WxOOvBdP1EaFql4Nq6+YLk/c4nSO
3qnrq/K9lQZ6LnWMFLHJ9UZFXge7xWL/gC9o6eMvk/HvwYgKSW9WqBfYTKPW5cn7
V2EFOKmgboX40X2ntuasiUiO+aWK64t9rcChuyW4uEy6K/Aby9c/S3hKwW9qhzi7
ZQAQLlufAYjAQTegKOycvKfZc61XIj2AQj+G7PyfmhcVAKJFs4sftUhOW/NwaFmz
M1+q9Mj8F8NzedHPmNXTYv7rcg7ZaE3vPjHJzFh5EDlTwDUdiNm0V0ps0q4+DAm3
TFieR0ig8OtJwu1U14JrVfe/1FcqHarPXwkTAlHIfvqor0r0pzYjxxaxMQ6Di0Ou
gkSNOxuhpOFX4Ir+6OGG27838AIFTIAEjxIXqFUez6m/u9bCyMQxvQpTPPjr9S3J
mvCn+6ADuls1JqD3+emvmw+P7Md7IuWKDe6nC2PprIFycTUB10L2Iro9OFMvgllA
6lwiRRxXxdcp5146iZYvD7Inazkn5LUpfe7OVKJjKqg/IZ/CMf/Ld55Qeu8kc5um
5cbowdmBP3dDzMwfByxZqsYqmMxWi7Zk+utMBzAxgBcCr+Y1OxOwgl4qx8a9jE8O
RXXUjG5lUsBHhK1xDTwzeZsD1gSzMmbWYVZW4eAtn5Wcl3Pc7PCjuZZ//gGTs0KC
82FKcaEvxcvOiW/vk2L1x4aKIcIYwqd9ZrXoEJH8TvN9/RZ5dBLdGAUsy/Kr9IQQ
dUBUdH2SL3Bn25JBLizDHEEoVqZlxIp94aB+U2tKdP1+Ik1mYjHmY4q8go71POLr
aas900DHBzdV1rYkTaYCcO/5U7Fep8Y03aJ+l5HdHceVziUPJp+HYdWTOlzXNZ/r
QkeIm5xT3ZQPJWkHbEDvPJRfprPfbhGzseZfXdESi/VMciL6wX71pKgc7q+pwrKG
c08NN2JuUSm9pe296nBbEjV6Nx9kjdrBsyCs27jdaUkU1BO2cU3wyLyowgCV1p+f
tkVw2mm+ZAIqE2kGse8cFTjIY1x1SX+rRWKY6EehssgYFjf+W89x29GpedXMCKyo
tXOuyvIlERRRGmNFLsiRoyGYbx7DhVy7nPRQ8iwJXeJq3psJL1bkb0DLpFZzM0tm
C6uUgGBxELx0cVO/2ZICu8VJdXhoZHVfh4AcRaQCV0tJZ4pbOYvjXmDhsKuzotGP
s59y/gDtHWVfh0mf37rguVXxtZGv/9bZDil5xW9y22tJL9HE6zInGXaz4+CAagAC
JanFOyMdVCr2Rd9DRNmb3PRJqmjhFHcskFnLPmLs6+WtKdEnOjFR/r/+iXxznvlh
3E2B2ZkOuwI2R+qXOaP3KMc3ITviyHUwOhxn5KmFHS8iQ/ZxaaxNKXlgDSFlSHjZ
HzYEDmib3X/XGJWf0vsOBzyM2C9aUwinaxJEyg3cL9R2gko7moJEVrdczM/ilE18
Ua45MM6GHKq6GD4w+n8vPFddYSLG6Aq5zbghYiOUgcC18XCGUcBeqU2e16paI++m
9wyvh3eGFPisUjddDNQ198gZvf9jMU61LzQ+VrToSYea5ppaYo7qE/Eyi+8eJwB4
xYnTq3jxjvXLwWP800PuDU8pJ3y4g4HTEkQ0OjvT28pYdmqdO2xo+0LNhNySfCPM
WYR4rhk6pPCLBihE8Sy8WFomWFMAO/hbLbCsqJShIRc9U52Gh0jBghkrf+e7MsGZ
A5dvxxVbDNVJAUG49I5rg4VOiVfpfStfq0Z322IgHcsw++wx3G3RckSQnILMY7AC
qcwYKq6sq9jxu+nHoZ/zQCT/MYRxwQayOx3UXr9HgOosNYxHLNsXzfXm3W7bZ/6A
9n/oEx2ABYm12kxRFiHltxT5T/xUMGxiP1Nncg+t5P7Ae/qTFwV7IrsUDAw5DTd8
acsdssCAqmt9wJ4M2/Dyahb+i3a+iHWo+5a+Du1Tm8qmwjSJ7kLnosFpW5JMAdXr
wDHxgpzzPJGIq00I3Dlm6Fou3nGAAFzjh7zaShQtv5anZYjkmk5lh1w44sEF+SKQ
6ePIP8osi1C2njbjR4zHrO6mQT3djP4ZTiCNEE1CeeOIPao4pcXJ2j7Q2ykPaV9+
eIy3Y6Qhfu3orsthBZBX/p69yYqNGzkItF3JKZKXHtFnVcj1d5iNLvREAvdwPzHy
uVbLK6BRX4cPVmDqKyUVSNLwZb3ScNXVVYytRunYZajz/4oSOFMXjl63MvtRQRCG
dPnzthybWdxNDAI9kISlWd1CVL6KkMGXi2+wUCzxeCqjkk7KJLvJF3TV8nW03VDf
7dGlQTMnl9LqkRMTI75wgKwlnXykrUT4ZYscHTTgaAiu+GOzfoGVMM79vnXD/s5Y
K5+0m0Op9wHWn+8T5czXDh7wNbghQf33584+XbN9lri5aFra3qN+8dR6sYab3sQt
NzRmstykl0Jr5lF6vZylxWQqLGsCAsxpNGkq6yPk2NUa0rS6v4nUVafm5EP3SKQw
hz+qTgrVQ/Vidbvm2eLl7j7ZQ3hLFNvBKyeaf6hjtqwfZml8EnAd/mG5atJYE6Me
Z/p140FHbQbGw6EPICjO7Z/wxkRsAbyXsQ3N0Dv/OAcnYGXjG9WZARm/PBHPY9ZR
F0jfU7XZ1UhiCdiCd604q0XRJCM6VrfyK/6GFmy3LGPxtc6VwTFwBzYKzwO8TAj7
I8FPgqUQ7ca+la5eXyeofNJND+e5CZOOnE7ODI/dUUNaGu3XZqYPLme1/Aw2uB/7
Snz92cwUJAaBbEBCpIieZG0Lp9281XTJaSrUYAh13rPNeyPMsXCfdbox/ApAQpFG
geplumJ49/UoyDOtp3ho8j1Guia3LJBXeM9Nz2NzOsbyCJEjtlMJJgV1LLuQTDcp
aOtfrHCMQhF22aIk9TI28ECPQFVXxw9rgKyzww+qrCxdPtTbe8BamJi3NEXS+ide
jAdPIVkzo9OB19KnFdZ4h8PYTET3FNc4438KeF0w9jl79xk+GdHAxYMZNFATlSfF
hIyeSNTKuJoegfPQBg/eE+1kS2kbPxyop+JCqi7/h4n17y9uyG+sjzVP9tdY14M9
9szV04Zx2hPB4LNaH8AffhL+yOXIFU9m+AAJtvuV44PNLB9mAZmo6flSK1v/Z8iC
pTjCjQKkTZCduHN0TuBQQzy5HZPiaIPCA9aXoDVB1yftwRUn2pFSC/1dGu1Rr0os
MFF8YiQzsxMSE5GjsioqU2PeDlnQqzC2YwyXVGCyyDO+szKG50obX7jHlbTBgv7C
F8kTnUuUpxXSmutaVnp1x0sonmrvuOIhF0aPrmn371b+BhoXP36U+KXGQVf17eKy
hHSF7+qlGI/Acr+1ZZ8Pi+SHWVmrk2Yb1Wgnbhtt4JUu4UJpNIAd2+/T+UvNiG5e
Kmc4mWSWyb/Rs2z/3MkBS5fNMuUFhoswSa67HW5D9jFk7T4lp69Z+YCKm5w+ceoi
6S2iQXlpXSTViLBuIlk6sz4mNBggHCmy+p7q3aPnawfh3ijtsR18XTwDkImPST1f
VXdC31wjiufnx46hN3uflO+i1rO1OWg/p+ab49ieof+vuqbHve5GcNvHGnVLnPhn
fBrkO59F2tZTkZK7TLV7dA+jfTvaIBWu0tqDv0EjebbO4b52L2s2nBOcbeAIta2m
vNjaiW2GTvKVyW/wlVqGl9zKplcBebEamUWvpwUcMkizlchTjL06DD4cQthMR//W
HI0KfTL288NCy/2qnuxAfg+ShU//p9vBgDJxHuuEU5DlfoUC1hn7wjPFNA742ONR
TdNxEWHD8tu7CAN2y/DgwKprKrnHvv5jOwsHvhdf4N5nlYY8T36HF5xIrSjZ5ZT1
qn7gNYaMhu+xHSRlz8GM6Ws0TSHY85HvABKE/WfPDuPnG5KhKMMqEpPrM3BImJjT
qsgknds0Y5mPdPf7I32td0rU555bMyvUs6yK9c0XcAfevJIZ6TYm57LQCBcmiiLR
SuTweQ1TH38X/S93CKFGyKEvBcLJZC1llNoOmtfoqs40BEqknjIK6HbhnXpUOlPA
gBmigPaWefsm9+0xvciTCLNpr2aZHS41dMdx48728Y4QsYqNttPa4ET/Ry+lbE54
ZcxHEfFMEyUfIiRk4cELyrj11tU9CIX1Y6gLjAw482l1U6Gnc1T7Jto3VDYeSOU+
1t8VGZdUswFhWLotehcFit4GQX6vNz4zMpnslwbgyIT4f5Fp0NXGW54rCXTvHDM7
q10+g9mztG6dHoABv7PLtQB/lnnuRMjum/YulAU2IrSRGUQovhmvLmwS+H+FyHf4
oFMcB7MbMC/0W48Sz/MYGFxfQn5MKBg8PsyyO0QfUI1SL5CW58Eo1Jh+PUN7vDta
4jJ2vuFxpW0HG1Y10fa8GTfudUzRZX+CWQUk3xnjH7ej2ck/uhYXlVuhPVb5jj/V
tlRIfyFDsQpPawZOYDgbhvKAHWjD9p6LChcsN+Uz/nANrc+orSk0OavnikG/H12Y
nRNJJfJllPdbmuQU9MU+BFsv9fUpmlXyRWWPQOmZ3q9c4yGZGuWRD87yAndLf3IY
fJ5m+KDVsRXzzJZ+sM0iQSbqYwJUb5zRajKq29eJZj744yiXgMG9zHGNzEYkiUi+
xkGJtdxZP1O9qM25vWJXNJ91bGqAa9HnbrW6XESdTq6StSArUckwyAUcACdwB9Yp
pfEEI91nAIykfosmaNKY2bgpEi/XzQhIRfNHrtBF8BGjgy298A3oyVdspCySwcw/
7DvRl/2h1oYlsTRmoiSB1LI2BzrGkky4P9e7g8L2b5h6bS4uz8SM0NqkAPxTQ0ae
ySvgB7aAN/g73LsuaXMvgJ2Enxd//sHedZ5ZyV+tIebpyViClkK03+BZTp4lLtNp
UceOUHVJnnMsbVijfT/qXCAp1XuBWzBsYl63VcctTPpd1PAYoKr7Lc3OJqwJYSYL
yXRusgLJDVh3yGHgFoR1BMKmQpzJF9mtoZNqQy4RZOGn95+1rK3x8IuQTQYQABt2
Ds+wR2wl91vxbgaKQIOPjtVj24qYKJj9D3t3dLcEU0BWt/wzqNUMud+hHXAd0KJY
RbG5zf3DLhV5dSaNxlYFVhYFXsCk/gO5l1X9oX1d9q0r+jhWFsItRawS9Tv9T2Mh
0ozjkYYaGvFTJCDf+v+NGmm+VBnzNaaikDXqUA1LPhK/6qMYjOlNucIl6L43sXMK
bELds0T1Je7s7dxyfgnAaoFws450oHqQx2vALcKxPeiNXmPLGhQ4NuV/oyIhhMoD
BEoXdZS0Htib+k7SgsRcL0ZEtb3s2t8vL7ROpo7y7P3TY8n+9ksYsn1CiLnzYsoS
SAuNUwbvG3NjXEN6TM0kUPdTuHeiL8P6/+kvMoQ1NDWsKxoTTOrSrwkM+hr4StBh
Esw3/5/8wgJMYtjK6sslDbs3uT4mKEAf8h6VaS5p3h7ttREBY5fgPUX/MhboL6Kt
5sTJ6x0eI3rxIhoTwaDSmCv8lW8B8UL9EG44aQiBT6k1ICM3gRfLQHar2pGUGcoS
F7K63dLu7Q0nG/BK5mAORy6+HCNfIgVeFZ6tR12eVR96XJGmQNHpW+aSgJ0h57hC
ij1lS/QFCTjL/ldMFfkyeHoezJmUmJTxxNV120+JU477J2q7m7MIOm2sB6ziXHmz
sb8Rc2tBkQCDQa0WF1qj8upmI3SJjI3+nJFuMgIAnjmToJfseJg5eDGahCgkhrze
IXJSTsyNrj0DpZlKeHI7dl+J9cGifOR+AR/TziP7azXTE2Ug8HOnTpvodQevSQQM
olwOmKqXfeUgHNBhWLX4cHRW5rpXm7C3O9mx7pQhL7kbdiNNn24/+EOLsPf6vAa0
E8V3bIREYvP2+cGusmxfgZ04cAnIrBqgIskL9/FR2lg9AHyKw1sBr8OQq6ukymxp
QPKpp1mDwUTXcrkkYBVxL2fkxSrmUz0kwOMhDw08fNUa88GHQJ5HPik3RQ7eeYu9
0puCqhNCSWEY/KaE0PJl4irFQYR4Je0OOOXg5cHvfcb/K6ucC8WcpYbFyzKQPI+T
tk9Gj0P918OOPKmdkBZNdHCZ/uXfsjBo2PO6U2gMyh0r5Y8vZm2JH1hDQahAXu1A
F5hwZs3p276QXHX9AfFx4+DphDt4FbS9D7H3HO1Zyy5X+J6hUqVLL9avWBsRo1Xb
7je8vIOLOdvwT7zINynmDJn084QNinfElbRFpw10gw66D2lMvyd1aJ/PwEPh2u6H
5v8y9n/pXVPboJ4F4mZiCIm41hUk+Sd4jgZPANy8pF/GbPoyeyu/R6Nyk7KHsQna
ONs5ApP/5aSS0sSsj7am4RP8spUwYmzJNYgPtJEUDXsy8CcBCr/dguqgpwl+mPVh
yGFWpGEP6s+L5eC5g2F9Du0fSFKffvw8b1bV0gRw9Y9Khz2lvTdRMpVLu4NnO5Xx
PfdkGZM8JFaHoQTVFHi7puPNC57nz5cqafWOTMCweFs69PdU6MZrVvUk0ii4RwnC
uGqwnvyOvm3dBip6psxWMcqarlpVcPI2mLZ1gJYr0JSr6RJOt4C34sc073lTMQbu
07FA0HgG5XPmViJ6v4LFXVz8m8a8eFUvJyZyjduyIRXsyjcWxlDOkZ26ijJlM/4U
ME3fOjWKhbzWSG7WRJV5uafxrsij94DTtFUhYXpm6k8iujdQlIv+FPZXyTnZx9EO
xPW0DOKcHGW5tF8PKCpx3obT4fDq8kbiyVr5c4yQrEUoV2r9LRRnUMNFm5id41le
AVK/9XPQa7jqzIzIs5DZN13A+ZSgtF3gNwQ53fOVh9cv6zwQlFSsyl9O31PovsCM
Oxx0O0GwZi2JUzN3b6k9EZzmsmOXQPILAhXPnEriB4/OTknaEJ389V9scI0sfZcv
CQ6dVVi9MgK68wbVPz/owh/CQq4IesXl0RfkHV6N6c8jFePYRS9mJFRrxkQxYV4Q
G7PBnIZ4E6bZ3dngomoRYY8l+VSEsIpve/+yrkV+VPXOyJXGwMEE3sJu9kDmoWFc
OMtT8dOZrjAlYMdi/VadXbF0jhLpmOi5tfs9MEKMjSwYZ80hH9uElveaPFDlqVGS
jUraUjK/VuJZtpDrsDnZPePasBhetmR/Lx4Hx131D3yvJC03sLRELjPpVrg2O4uK
XiXrUh/qB1Mtw7aAAl5qGIo3irGW99wz43dOpcKNTiqRNohA+oNZZM+rVH8Rp2vy
e9BNVehFd+RVSBXM29Fol7oIFuBPJxVYBkZCeYuuubwp8tHn5d1lApMMCUlj5vsG
dULooDdUq6UggdYHCPEHlskOyXZF0Y+Hzq+DXAGd0qE+yhcJh9nIMwAJ8OYk1vCe
NrJWfFDI94DiC/zjGEPK8ZW+76KpTbyxO2srd4L8Xe5eRSRbVRM4UPU9qjlTiQLF
9QkCwXr15HLB/s+VZn80irD5Rman5TJlUFOaowqm7XnlsbTkXSyW6RKnCz6EltgB
eHWEHGHOWPlA4b+Vg1fRxrYEaHx77QatSHkkPZ/J/rPYzEIuvLn5V+uxiOaQDrBp
hL4EsRa8xONmYEbnlOLOOqTaxFrdfd1szYdGgIlk/8oGbP2drNj6SvkjmdPhsAX/
H2pAvDMVhdZmEnwbJ5c54LPe37FeHtR9qSzlc3Bs0gJTeCwXzoTLb1+O5Mv5aB8D
+jCUuPeNZFX/YEGgKK2iWh0jDW7vT1DczWr8iA3d0X9TXxi7xWwt8Dxv0zp9QQOH
lOPojEYygu/FUHL8KohQDih3pu/Z883vbZsL/2Bevosfl1rv9FlA3gMXQxt+ZCVT
yulZhl+VHkwrp5MFoKq5IGAccbWYa0/eL3ksIBW6UiKMU958meUVT8OM/Jx8B9xB
QgGmUy00pIukFdfNPkO5YUOm5quGeTQwNfwLCjEjKMgkDMs1XUFOiaFlRHF/wCp8
kKP3pzUE9J/dPthirb3n57u0cm6OTTFp2f8gRInTDOaFAIEfF1nlHf+TnnNb0uRp
4dO9Bt57YtI08bN3gSgRaGOAQkBQImDe48eaVf0aLzS0saYJY60zEXS/LUKTxLu6
eU4US6GClAtxfYe1yrT1zQ9krtKtGGJa/mHnFEo7Ca71Q2yrc/xDz7e1LCoFlwQs
dXaKbk6hbDD2X/pdg0V0xtp77OrvYr8Zu+7aK8kPStzQM2iAjMZPSquz3KBa2qw/
ISOdB33Vf6iyyy220rMd02y9tkH1jqLHABxdXcmVWzNjUeNXNbjkv/NqgaM3xm9G
nti99JoiMpEUztbgFZ0JieI/IhMv37VCGA5wmrG1g7fT88PzESCwYmeM5MW2cePC
v/4nTIdbQyBv/5MDFVrn7FELY4eW9L6da0f/Gsc4XPrKA6HV6ERm8gy+fEEBimxj
r3JuOgEshkAd3C53WizUyMF031mVj9sI9fUkbVP7KTdajHlaM81t+M7tV2Xu2NHl
yh2XmMrT0SN6xkJ8WOY3iNkapUqmwufVIltO2WWDz5sO3TtDWiPaGZYj/7/x73xI
A/2i0wra82oeuKi4QzffdxS06BjJm3mbM9LnHW70TzjRsmTnDIEb2zm58SPZqsBA
MEuPSH3rU2dOFpgl2+rD91iwNppAVgbfLRWFIQ4a4MI12q9wopsekwZttdf7ekJ9
XYOQyTAtYLP8HB8+Kx05uO6tpx3gJuGKLWVDj/IeXKDd5cH4chFJwIe0ohJvr6+q
kkGt0PrBBdCdq5oo50Yb/1kymk7rDNamDtE50xLfac2ZRFuMnhXTfzL0+pp25C8J
bHqXXi4kcL20WfF5xse0ChcI7Ou0uR0budxnBOKrQUKLO3554cVZRG1iFgrWfhGg
c3tNSt3ZY6lqAEA+7K5AOs/oHDplciyvXkl18azEtHlcj73XpwOv3M2RMlwva5Ww
ZZkAZUsUejrxjcAHxHkzxw2bJBzkn0IH94UMU70z6lrjwBscLe4ixfKj1sQv4nEe
o+c6GVclCUWzr+LVf9p/A+BA+t46f0u3mwVoelky0IiDbxGdkYjn0ZO8WbOxN3y8
R+BWc+QPnly54uq+dQfpeYwt2bExNv53YR8/xJNIh2CDdhHfk2tC3A+287m4XKZN
L7ocHZdbTT7ZYzxYYMy6iWSRzScxlWKVEkviOlQy5hyznI4n2+npVfgOcg7MgVwY
jvJq4V7An30RbcmTWSf1TpwXx3a1EsdcJ/OI1UlHNvd7f2rMsxbiHX6q1wh2DLlP
fqZ9rHijAPLKl3XZ40T/luIxIyYZJmr+m9/Ph8K74cYqtdnBSo5DQ6+8dF+rV6L0
3RY2lYpt8fTFSPX+pYrGHazyPdk93wErk2ud9SSQmoaj1Ar1HqVBDfusqii0zZw4
5RBwltgvF3LG57srkOEfLPytj+dmuc56awrq/mhuwsBSzOcD2oiuU564PLXgugVw
N6pOFyGpeGcjSTXiICRwrCXT1dTkzo6yrzM5SLyTQQ6sdM9xRPJ1MfPuSHiRDxWM
lV7pYm4hm87vfi5qTPAC+HekPHk25AHS0Xc09n0YiK7o4pBmjfytEnnR5lq9dBc3
YLKW3VvBRtOrt18m/4453Rw0EnyX2sJqbdC68ZpqSD6GRFvnC18E6HsbqgGSBaiE
oUEvfs7I1oRErInEn+IVXl5TdJgvhsd7Nl1hIGjlgIyXs3mQCpADNM3uW2FiXW+l
ipIHqXhZ6st34Z2emYv5QXz2iSM4zHeL5WtmeoQe5UzuQ9Z9ed7acRgiUygzmZsb
z6ydYUY6kSXImaO8/V6045UJsbSTi5ww/EJPvU2qfQkPhaQkFCBnxlAYEbGh3F8Q
RRZ3gJO2k6PrKaGCyrpbot0N09t2jy3yPvycUNtAwKgkUzLklykH0Cn7It9RQsL/
7jpqHGMRY4Xon2zN3e4h0T9nezZFgiSQP6WROcuSl7Cx2+p6xJRvnC1weJhDZ95d
huYH6BS5A5oN2AoFB16mg47jbrhrQrTj/u7+Bs5an6+EznyNaExGa75+oKDXcW85
cR+hm5R4jYcGuWy7EIoF7T/QK7CT/55Njlp830d6cWsucCLtzTUfeEEnF8hr65tt
Dlx9sBRM+5+U6PTlAYZH5EL7XQsGOs1gWJrE08cPng+64C+AwtnK9KS1PwMcTdVz
RB7gfW2xH3ANAGx+6vAdjZykOF4Q1aeRBozUT9jJdRI3QQroz6MQq8XFJWNPAZpw
y59QKlosOcUT/TS5DLQbCMUzRWuN9b2InXHbhAjjD5cnIt+4vKcjAZzHoMtUGGrz
y+gH94vZdNNDfR4QoVNnQL8DaRrddY2pBzfIjxAQH3fT9JQdUj6qnQ3O1ZaUFo0s
OjK7yocdbjQdgEPz7blOvN6q7yjbgWD4WLXql67HTVjRRB3LwqBltydX0wxcvG4f
NESvxDolFxF9jXoQ79uZa6x9PmmrfO6PLDaqjS1bWrRuiIv3FXT8Dv0YNDtWhqSZ
GxRKXFjrWi3bjkZgfawW/Bk+EPWrLSadGJzXSSo4SGFWIFiSrQhyIPlRbzvZi2YJ
B0Z4FlYI4wpBEujIA+jsioLxXW6ixU5qwt98EIVbvQawI6x5uG3Z6jiGdOpVMoFr
uzxgnlmBTCjZrSBPN7ozcO/qWyTI0MBZaQRNEm0V4wYJdxmTFaeZQQwv9xOngaGS
5s4SqO3GOdE65AuJR2DpMySnBUwiHLx+UeFKJ8WWOQi6U13m1CC24n+tL4jxUkjG
OcqAqfJUq2FxBd00AVNj/c8UmVfW3eJjm2SQ9nue+QJQncRibyZnojLBdMqHZCLo
doRhbiafrNapQZCphp7sxcuMqN56B1TlkzhhMomHzYbLCULhOlp4eKhlE9q7Ylq7
YfPaCkvVmjyTW+DD0ZYexQKuskyGyjW2dXn52SzhjjHMlLeRufB08DwJPD3Ze4BU
YrZFHiNgj0FTLZYW677xzwCcqfpP/xDjrVaixT/zOKqltjBVtVgf7n+CngEc9pmn
qkJEiz1JK6pjugJBSilYogZ/hgji8mK2nMSnjwqCxNQ+OFD5uOV0yE47TiIFlFhr
y0da3izJTVj7Gp5Im8k7Dojdpkyrf/RXxDAZRBJBA8KsSyweLcAMM07kV0nWhkXl
hgpKtsOlNFswfVADKbbZCqTnXdDk5ybNYGNr+5aMxwXn3wXu1DRO6coWlcqNXi9x
tr3zrC5R/Kkya8yYk+ztgflzZyioiiNe1TFuQJCdiWF7BsNSlCv5nPYY+9vY6NCH
m37MunA8FuiT36UWLuAUe/uOYXMPqzr+0qKdWMvhIKD7MNWrG2sfuEbQ32Tz9yVX
x7Ru1Ns/XvkNMflt28BEt+3mevvofs4JnaNyis711dxEf5IXf/mux+g2/yUgiorb
XLpYbtnamZ2aQpdpqCVhrvU5L0bhZoYvwNDBNQgQCnVLLGrM4MmRjrpzJMB7hQE2
BPh/e/xn886jJRPkEONHAV3n02BcQ40cWs15AxyNUa0zzgEzAiatHQdKtvA3dDhF
kEl7SWmFvQ6si6oBgR7xHSfnST/s02319Bh0H1Q8wDeXRAPCzasZzLj1H2FOhbBR
KyWAno4VBPWCPHLgFWPA68ZRFWyNuw7jUezHXYpNcojKoQk//Zgjhd8VtX6xUMbI
VHxuSQyGHOTtDkT+6CQVHjMjRJ2MmqUctWwkkS6Ru2qxC0RyRDd3PrKsugcranER
QDRE+70gvA2jFs1hBJkludZt2Cel50tmyp5z/FfFTwjkmpF7osYl+W6w1YA6YMGK
bnuOq8s1UbO5ixuM4kS27OFwKDQGXXn/P06vx9kHJ57vtEJ+ngME5x7GG9gOdCLN
wgvCStnu2uOR1yPu+cP65kqbtIIYwwrgxIFN2nHWqLTQ0bPZTAEBqdhZiyqBcs92
TrMDZeRUP4Ih6I3HpcmoOA/LIuGx0S+Yt046uonkSCITYqWiKTvzrlZQf8GOjrTe
I5WDkIyuzL+zN3ue09GLiWyuBXlXxbegALtdzD2TZP3VNr8a3n3GXbXjsAdiIK61
4kmXCs78V57dkivvLIPhqgazOUfhxC6KyBKKLW2N2SN6hAj81sdRKZgMYsqthbGR
GkIgOnG5KVyyV2Qzy7Nqb5bRrgtE34PONaIYlXfCLlzkzy1qWgjTOLCdEMg79sTS
Ag85LYAaLIFGr79Ue9e+KGHAweAhEpjTPq1a+3dK/GbczhJkL75euBJGI5TrXePd
+wK3M7MJM15JxNBhDT3ZLKSFSEywQSUZezZ6LiBZSy0y4GZyaINKcK+bus7Nfceh
XpRXm5vyfDU3guDaxBDaHee/UbSwRdpxo3tPVg7/G3Xyzrf44knbInCJYWNekBZI
Yg9a+Ct68sTMkaPpGGZfVpWgzbi6OEirLoTO2VFr5JtoRrtTaDjmKit8ct/IwwsE
emckbqpBguIgRkOMDQjrAMBUqUotwRYBufzU5rfyWuceESg5fYij0rasrpGi1w8z
fYBei9DepT2Le6MJEh4uXEFy4uPz0UCpD3MYshzkI488MUyqlsoPM2hb/XxTPU2q
qNkvQT3Yyg3v9mAoTvgMXND3W/WJH6dOjfBdFrn8A0QfLtOY16UsI2QyrVk+4Upj
wG+OhmO4p1h/zIzm9FC00wCdkwjmutprZ3KXrCIQ5Gf1pASfSLceoW17skL8z6Jx
d1zhTeHjNo4MpGghs5F2WPFfdg/aX0DPnsm2Y4W4XVwi4HmpFu/tdsGFGdRjydx7
JjVg+ObrcbjZlncS3Ga86ZhFHPDwDfEF/nnXu1DGz9iE4xxLbCqmt1XNnfpvktkC
RjqKibkmwKMLu3LC5dkpAqgTV+JWM1nVfXjgfUnssq59veQLUToNuF8uexEZXz7D
hC0pk+zd0OJ6iJzZbxQNyX3t8YaRytizOIl/P4Kc1AqabVYMp1iN4nUYUMMO/Eqn
oqxM4w1X//nWkj/Wo/FHv81xizO5kgO6fKyWED4WiiWBn36q8Of8XokdY1ZqmLkG
a6VCrlX9xljYU/OH0PajnFMJdHcpMVggYvc4BuBTnJgrVz8v9hoL0EqgXLkNXjO/
Wzj33OmhMgTHTb5CHC96rXWMxEIt/yQtSEr/oCeShkn9C6bCGsjS9zvcuLvI9wxM
643ofn8J1Rt78pTCzEdnB3dhh2pX/oRBgVDgERuXrIoCp5TyDpdIDMBeZSKK0Fju
p/ujiM0qu7qVyB5uHvSwunWh5WYqoA+XUhmjtCMV/s7Bwmm0i578ZnxitiK3AGrT
tXsvdfEu4YflBI/4hOtrSDvcBd0W02YZyj2ZrQUuUT2Dl4HjXdufCiHmBq2B/lEX
KqT/beMxa8lBs7CFtkHqPvdWKxu5OMYd2MvxGwvHFWSNDW3KVBOXDXODOrUPhgMB
YVa9kUz5OWvQtveWHdmmmZ21mt76NRjmaxGIHgtUFS+0ZrrHSoqBMBCASo/pg4T5
KK4Kx+su8gUwq6vGm5OmxM9xtGGH23vL+cdw/uGzQzSr0r7LE0NpRc2axJNvUVcS
Mu5iTh0bJ89IvjGQzTVI8atFQj2QpXHt1sMblseqJBT5dLYRSMvXeQcPskT6tYJa
aJj6Dcc/pMOdlEcV/Pg0XW/By3UuoVWahEGnUKdS42wrroLbFWsJsjdrjZPBn0Ac
S480ISlADnEufRxceMB/tKQIl5GCm7zcEYqUftMlCh0U+cPquBl8oK9hcP51dTiq
fTSLb4duUc78vMmkJe7cz0Prtyiv5lKjxCVyFPvWklv+vVKc2Y1CzBBX8AomenFK
PJZdmbvQjNdnGd4xJkwj6SREQOfxO6hZXltVwfb1nVE3iEqgqeXguv7EFoWATqRZ
ZwlzNcdRiOaScFRDhcWoPXpNGzrPin8/h8zQQNzQws/hsksMMn15ZMyTLrKOfeaC
gwxnWx0rnFtk3sBJGBFy52REX/1p8WmICp7+W+uMJCdNJI4adO/8g0oH4C83tLSC
rXArVvGwdGNO6PIvX418s4eelCgppGhkBstipG2hA3UpyuIhXxvolhpHy8t6RpFZ
3w41u0bQjtigNBpsk2lgVd32eYJIF3CWp8tn5M/qir5Vcs4Ptf6v+0ITFQzvORuq
Wa3o+qPPmcwstZGCdRIPjdOXWiUTSRyPYFptQeU5zQzo5M+7vIyGTdDv5LpEOTqY
6U/DK0e4Iwckm8Oe4XZa8VDHanmfMHKyQpvtQPXq4O4hioj5jNp9vCbxKeHl/Xc3
qmm7pOonCQuGlsrPsD6J5rY5i4PSIj3JfZWEm1a5lpCTgCvkgZ36tkAAfsPTXHEA
wmZ5droeWDez8OasxNzW0dGBCPVe/5FoFxI1GywwM+Pn0yWLbiXgZKyNIKG14zTT
9xS/wh2rI3b7fAODWdeytLkkCZ62kCDtOEiG1ket4Uk8yutv7jueLC8FYZ8nP+vs
79mjodFcB7SSSj6eOybp8d5qU4+xNWRouozdWFpOs/xfPrR+7iBxrUfX54rLKCow
h8gFeytysLNVxXAuH0uPURAScQsY35YT7sn2lMZiczF1bqZr/CJ0IH86KSZAWm2P
+/M6sStEt3DfxklF1xtyPDxe0ayIOycpvNg7M1KjeVzQropOStWscqk0/7tbdkLw
GpKD8dJV9oGLoh3W15KmRqvM/1MJhT+xCI6escZzj6HAuP/yXvdn8SsLEU8Ny5QO
Y/uV+KTTfu9ztL3tMj45EebYl21sFKcJQna74l1tdIkPcLnemvF59FkEFhUdBiAS
XODx5+EDxgNTJLPGOoZpxWnFVa0kROC1JhMiYSyEjMP9IOnkVzWPWdpUdwdoJAQj
7jIBJZ35OnO/aGEcMX41FkEhUo9fuhDJSQX3zqfX8ALGNFsGhydlo9S1YHay0QUC
Q21TczcpzT23QYbHxrmiePB7aLZ99Kzl4icDCzQEW44kxYxKx9xYXBdFQQxWGFnR
uObsgIZfWYn3z2FqbIDXo4HIASEL1Sa7CkADEMN+ARzwTCdVc+wCh7hkWKFM7NAZ
0WzWJ4CWpLfbSKPF4TGyn/aisKb8N46+Yqa/YIu71cj1P26mZFQrmlKJw2ONn95y
LLK2JndBynVdHQiNknhHtPLgyvbowIGl0BvDzQcz4ZCIoLJPjK0cLyxHunFjfVa5
dX3TbLrAdPIWpRUOEtLal9uT/vAn3ZpjbVXGDxxuYPhAH/cDHWhkvTG8+DS8hGCP
5kFhgOlZSqOZZaTrhAxUmw4gXJMGmiAMQkrGQrNii43LsMQ+r+OvvtGUkli21weJ
kMgcr/r3fl19dX+X3kz6YVNnMOMoMTibib1rDgnNbZACrR9dtbOt91TqOPSZyK5j
Mc4gK52SSNlwLYRLHRjkxybjfBpvH7pHg0RSiYolOna1igkojUyIgTw4ql7VjqLV
JsuLZFCC/oh0/8VLKnKa4H3VUFCzUpB1qC1jD6DYO20802L2bZjulOJAGqCdJsD7
2OqShCLl8R8NqqR6YtAN4DEnzPuNaX9C97jpptLdLyE7OBY7iGkLHL/GEOHXi3X3
Eeh3TWcU9oxPAY14QRPC0izBI7guE4uwPQc8ZHxamL93CI7xaYd9MwaouGkRF5IN
8GFM7i7nN0JB2g1kcV5GjLSrFoNAP+yoxouMXd8+aMoKOm1CP1Ke1mF+x+4DWqR8
enOWJK9pWI3q3Ibu/7THW0qGVpbBlKvAXJ4yCiy3d70R70YQSC/YH4152MxD5rXY
Bh5Mk1JFKdhVGN0GqRBjnJUfabziu+yWeqK026eDd5kCdMwdI1rJM0c6+lwMjCRj
W9zhUHTeEWsOlOwKU1IfTpthhl6XFvparMGsYaudy24QH8WWrcEncZ4EuSozEcww
u/j5enMf63CEscxTMPp2cXaz3pDvMRlA8qdM7pBlhOo/EQRsjQR98HIcUR6PLH/k
VnB1bxU/jTKwGE6HQlIzGzjlDEqmQ4/AdcmgQGfOf3xXHfmtv04HTaXceMvLV90P
LANtlsxACq8ukpznE3LM8XhaAcpaCJaZ1LTJc1qvS3WKc0nkJqp3hM5nPiLkogvl
Q9ETQ0x91OX33Oi+8mHkbSwju1B5VYFRUqfpFPeowUuvUzMIPnE7tn5WF25YRsz0
e9p67Dlf8G4LaAQ+KQd8Dys8J71R+gdjzBHFmDr9On0q03sSCtZAVgDlTj0YzKSc
blls/SlD15SLMDkjUhTYdrSGMYMlYu+D6iDSts5gdZf6iONApxNrFewa/79/ynax
f1prl0Q48VrqkBdwY0Il+Szdt2gdhtOxdqW9gH4pnTqhtCkLiKJBv0B7+OV3KZuP
TyovoEgN9yQBl5IvBm9hhqgGdGzGtDh4VprvD3BxMZnTezypwzFFlYXsU0Afb8cu
INS2YI65W8ARFcI9Og7XTG0L7jVVV0GL1exSCwZTQAb4I9HEbtLiTz2f0+yA4GQv
SJut7goYx+looNkof6lYF9mZStLnzVSK6KPyROZJlWFpd1sHKL1GN9G3ghKFPmMo
Aprn7W3+oh0bj4x4AOX32NtRrhQShleRYeprleWzBBGoQormhziHmZIAvfBCygDT
lhAxQEStBf3UFIS+osaJk8ysTGQ3sjwpnhu126X8y/Dj3AK2NuW8f1WbRSc5H+nM
ifAU7etd0D/dzdMntJYNdwvWl6xI0aGLPnHa5OoRQ60kISNIgbIQ1Zw0VJzBeTA7
1wbGIUWeokqkHG0wZEUp2KsKe1CnmU1WvG+J8hinppAkKDHAS3702akLCxdAFtYb
fop2hMprG8ei/fZf36yb3jIWGnlclSYVTNcyqfYpeoV53ZCwcZhz9red+Te1EGJS
iBrcO4HFAvbggYLD4HZWR+PX3y1zgUentEpLbfwDn4W8acykXLmz1LZr4+VAoKo/
o5vG3085c20SkfJptysGQ5gqF5PqJKmW9R/Lh01MCrwW8WC0/8EEL9c7p0DRWujx
dKg27eWP3VfX3+YYdIoq1qS+Y8haj/WuomEowN8aYD4iHTdlTHfqbf4d1GMsUz4P
P8b4DFq/wID3XuMgg5PmTg7PCujG+AvvFASlotSJ8VP3N5CRsdf2fO8q5CDIUPJ7
1DCRJm21y/8WahpuQ2Y7LnobZJafHgf00gqyQyGzFgSjtuFtnnZFfSTCJElzWtee
KKedtmChUJuxhT9155J1MBGMbGxbJIaC+2EtMmt2dPyoAkSQIYKwH8HVVMlkTFiQ
m5bUiNqarCx69DUelQM3O+FGwjb2pb/mbHSYkWTsMj7FwNINrNLWG9e2xyIB8JLJ
pHo5FFrmNyMXqW4g8j++CA/WTNGpKnwc7j6fKWHQFv2vygWXAtytm329rSneu/UU
iHpYn8tumVWlgZZU1GtUXB/rSeB+sDs372JbaUSJlqEYnR+o5LZCkRl+HlThIIzb
0+WbCi5uAP5yJH3CQeH1pB5fErMdvIBMXfD2SqYQO9JzovW1vz7C5rFBGhpDzXGh
xicoUniNdseVDtPMfej7HftzKi0SDPEdCbo7a3Jz8UiyrpapknHwpTWwDTNnnhfD
5iTsdIzDBleLSNx0w1+z/nAImm8B8aO/HNdNolQePIqOg1vVMh4aBE/oUgQDNf8I
gkAnhrxJ4Ij07oN7jvmlIO8McJ0omnXvlHYuEyQRQaw5L5JHFTMwZtL0wgNuzuqs
4cDWqpbzLvVwSh4wnr7W4SxJ8deNGXIPNPykUDPfqO3g9+ydn+TEahvoZBwr/6uF
uhyJhoVjbM/b3y9G+W2Qb3PQCgij/k/tURw2Ltxvjq0xAHr8N1FmYsywUTG2Tsyg
nHTPRf5flvJxe2cyefta4UN54p+m0/QlxuuIkqgyXSxfJqSG6mL9UkN3WBduzued
B2hLj9V5Y3sBC7qsVGwxt7cGtM8ybut96dSG9XOdHIz3rVNQvpSR7zO5ijD02EL/
LH7e/F9D5t9e58g/IGN2cyhH4MlnCInLOXv4HIZO792rq/Cekyn+ifX/TzCLPlpx
dTzjvrNCMiBWQnMikEXvl/tQzuMlm7+6bNAzT2lx7WQPqsdahWw0FgEUzQYjl8DF
iYHjHa9FJTFkQKX9dCLV6IwBpzak9vH+D7fxnwwYKaklBJBo+8n/Lzifm3fNEuVs
KLEGUu4fQ9LLqbUjTZOGVm5OdwkT7ta68dy5mxOzybOzej/JFP7zBWvpA5FSSLx0
03xgWwiCE7/dMdbGxnElxZbDzxJ3D6OZJdivp4FiKmC6X04j+jotTeN5jPdbj1r7
e5+6gdXd14ARrH8OiuJ9+kvwKuGyLntmUoH8a/GcoOqy/TiLuT92mn1CVQxUPMj0
KTgpjryWbV1udJo37WiD/dA/lqylbaGusS3dI01470D8WcDOFBY5N6KLuEjFBl5l
xNf5I3GNiqV5c9xFg9LZxMWwbWbZoVaxsCBxtXEbxGzlK2TiRjK4aGlxPCHB6HuH
rPfu0S/aeN6qjJhdsbE2nHnmynNbhLHzUQ5NMZT3jbNV7qpCoaCcilAce1m2HUap
aNlQKYrMD8E0um9mTgAzE/SrgOY+qGMHB3I6RlnSf9vAC9Pg3rZ9vO1BEPjS2Jj+
CgoB1xboT93W8eNTNTs9qJR+9DzsT6bbMeyNzlHaPXKK/SZa/1Q36imz/OERMuEz
/5zXzSFxqdpsC8Slbk6koOxCJ4G9WpBgGPf7bDGWRALKMjJBX8xFy6A8RXI1aTH1
WVSW8WZeZZ56oEcPkELpcHa1XZfopFFjzJ3aHN3X3r6OsF9kPdtXXZhPzjOEWy+D
nmSSE+sNhuYadeHXmArpfCRrvsOX6IkU8naTrHT0Xg52m4zAwzV0pgHpSA2jaFHR
g/FMSxTZ9eHSH6Wv751akojZbw2MVTNIyzAvAE3HD73rlvsrZehtshowynmUG36E
Utq6WpPeiXH+HnpU1Ee60gwDaIQrldhxuEkQH/BHthKhnVScjLICkT3h2ITL5SxJ
FK0bEuMSq8HbepvM3bS357GjkJNq4moEHpLVVDW9tCEIe+xpjuppbLEcHNbpzP1f
RKxbUsXQeXIXSPgcGXHw+POSOMRdLlNE5R4phQqTlEfOnBNV8UXH/+lCiu9gpB4a
tfZFIuEs6i0GMJPljlKNuImBPIDVEPSJh1HAq6Eli+p6ilojJ6kXET+B6+FbCIX6
NEkjiFb4qDSk9nDSBKRSzCB04FUsK0kLuzImm1lvGHQPE5vkeAUcC7uP3LS0jmJM
uebH0MhdmUFRPo94tuqbMlCOFJVgsubM+hRl6bI0aOtgW39FT9zAdSqw+GvXlAzM
FU5om7ZKAdb/YvB6BTuLKsFHXshrqklZNkBhKFtcG3WNsI1Ns797kI7ICy1eAVmb
1E41aWoLDmsKy0FUyOv1WdlBTnhwmj66u+M8mba3FAV2DKLsvxhAJsC8v2ZzZOa4
hzeFXEbrFCUzsFFixfak/pKgmphNg6uyzyLBIJ16tKad+MP61WQefJhPcb+AROWG
X+O74o1lWdKziHD/SZ0Z/UHo2eUFxkSdK/A+WtcYGBwJ9pgUBTkAFrTh1w5WZ33y
eDzSee5L2h0U8YqM4PR8fVMZ3iN4R9q4DkLWEZmuQUJVafJrzdA1W60z9RcpUxLv
S/bnaTWwbUYdyGJGV4dn3GaxCfUEK38s8rYbWOU5KAOjWb9FndA5w12oqDj63cCl
lU9AfkxbGBRJYe/WcAgb8w5eriueXntJ4jv4oC0wpdt8R7+6JY31jhQv6n9Whl1x
ysIsDjOMuhMljWA6km52/oXlD+ba9eeqkzoslb8Wph15Be5ZKmCw4bbZJGDvXUOY
1WfEaRvUx6/ErFMByc7LxheKyP457tyYhEY+vQd8uDWlbp1PtXpUNIK8bY4J6vxS
32MVS78Z/ixTs7rsJzrCUGQu466XC/mdEw0myQTz/0BZtzU4YiL3BxmLO1xn+JgK
8xdl/c5ECEU4qEffE/jbN8qXCUJYRUqVl4q85FkxBhJw0Zf0glCrP9ZFv/lkqRwe
h/+0U3YHqYdxJfizYIHQukTgMOhDpbBF7RwYvWWMltawTOs5QG5C7qagpIbj0qdQ
bHeeFNb1gTgHl8WCGINc4XNN5TgdtDZCtOLVphAMnWD1ExpjEIIv9zP/JBXkZEoY
7fUPZxZF3DECN+ImtOfpR9xIvZti+iXD1/I33If5Pk26vnQFSkTeeUWD36FRFPiJ
odubIgVHUlBb3OmiHxr5PB9qCeDiF/VSV5wpgJBs95pAf/swSoCB4fV2GauI72T7
o4fyoYIcInLKhSP77UYScdAkgqKrqYuJkkqA2zXGKesc9WVh/co0s198IE/qilJY
gdHr63+CIfFs3zkjI6K/eEaKmvtMemmfuGEzXCUNcGOJmCKQKCewca8LyI9RKcPR
/S0Km5yKYVl7g/jr3lulVSlci4GrsOy4at3rqWGrcOuSGRYUH3E86UXw6jp6gwqB
mAhHXnRkui3sV8uT98D2gsFNDrD40lcGCSPELxNevp9FHOjIltfXJW1toC/JI4Jb
D2eT+UIkaJEa/4Dq0k02sDo0oUlForQXl5uYH7zxCxGVxs0FWfI8RmhCC2bZUbhM
k4Ed8nrLELCzZFSFZ8aiSU/Qoc4No7hVUYvGaytv91yNcAETkMZkl3oeS/oepnsA
+0AeIte5VC5LLmuZ3kkpr4i+JW/XHFd5DY1rSvDTtf8dxvtN7VKt3Nni/smCroUL
TSRmmUkzC9JVczgFZ2XH+UV6dDBvLaKV+cN8/38dpVLNNMTNJ+Sh+jsGgsmmFMqZ
bMKmAwtQQvPsyQHkMo6gSXwgSm73jx0z9mCIftGxSgnTidyOespyLws3KDSdW3IS
fOCqtn96TR3eOgkKO/yqy5Xv9BCPWhbmGEGg+xC4DTwA74V+unqVErm6Tl23WmuP
C44K+E1HlHkiGvPyGljmZVCU1l1JK9l0z4ETNCbFWrq7uSV9ObWreszTm0M2NLt6
j45m0H+TAeh+UaCJx7aEN2pATqICBuwSjidU/Vvwbt9+viiXpc9E5h92Mazce8k5
8IRAN4cDe8iJ5IpTYbpwV30S6v+INA0+sOPiDS/dRLP4076T7QjhAamPJCU6pvR9
1aIOYx6V2VjcTK7quGxR6EtLTNtCklatKWz9+Xs1+gDoHt/rm1rd7ktWcnBuahBE
HCaPSDd9wwS5Qo9IUg+ruJDpHgQARJHdtL+DuXEAvZ5z3PSiRiX7j15shoKeuAO5
8C9lFrZpcezJAxM/NJDRs0hnp3IQlqX9ohbMJpkjG5fBX0fBhcq7n6Gq/25dYK2x
qKmR7OjSkismB7/tVvkbo8vHrgMmzMlXVnNmyFIR3Jbcj0GW56XYweVILtSL4RUG
MPaeV77Y7bdV0qDGvCOzxkMSj15kGLlKy1LLRosCGadUt8SExAPh0FTeYi9FNegD
MbsTR69QJ2qjD3yOOpqQmIshNsZC/ppmTPjviOVY3bxomwKrgjLPnpfwoDnql347
mi0208keV9iy5ti1PM/2TY/3NhbpusuDerV+dRhAAjCLoDCXdXRT03ayUSqv7J4i
y4HiNg/UWUZ8pAzy1XayS6XBrpm6ikogAJAXw0H1OJPD3n7A0Cvyn5sTox7PCoLE
nrZ9jMRtU7Pu+GIbO1JYz+o9EdoXSiZhAD0lrbUdP7zwNRPeNLsVWOHbou+h70Th
KS+ajWh+xOKSeuNuWcwnSzMdq4MXypAvE1hJVeUMHpdFS7M8rrfr25lISAIhuyb9
GjVjyRebOuC3Ldnjl0VFM+4ig4aGiOsUMoAQTk2tEQo8u52F7//aFvvMDKn/k4h7
hfNJDdlxZ4WeB+gY4wlm/91093x4p2ZqnLYoFt5Xe0lvPpoccYzMd7W1O9CW9lC/
J1MAkZHDSX/t1TUo59SSxcjKwAEOfn9hxVwsa1mI2VxyBja8p4RyIn/ZSXbq0Cuo
DyhibVJ4f/Uf9Rbb+/q9DmGODNb8jGErEHU494YtwpBA5rpUeHWX5M0PuaeRFg3K
wA6622s+IdOnhFtF1Pj6hSZnmKP5A/G9+c96Y1D8BV37Cige9WbNABCD6zYNXpgz
gpIE2EgwKmsOot5GFor02OV77+1OXTH5ROBFxBEzhak+wPO+ahPm6cIs/WjOJSGD
nzyRAm2KJXz8CHmJwh2P/LsSQ8btlPPaQYTTsv5vpVP+z6n5i3GWujdKrNQOT7ne
g+7G51jNP7t9aCsk4K0RtdZ9ax3RyBW7n9KmjjsbcGi86POwbvpjKrMYm7/IS53c
80q4Tvc795LfjPUMOPy+SVvK4l8q8w3hhc3gM1niHRifKqnCkVLu+YZQPuou8uUB
4hau0OfXb6i3ugolJQE/2WGpptxyM55EK/t7ZCAzr/BBJS5t3x6ZedElcZ9dwtM/
Qui8e9wRLnLkkp8G54cgkHMgv1I22zyIhJa+e4U5Tnvzw1M9C436H3HO4DCWD0xT
kfFTLxGiiPNcZ/8yZoK1uQcNlcLdQefMUCclQ1mDRCP/TkzxddbheBzJVq66qSAr
sHZbiYJEuR7KKIrMiY3SdbmQGZ2rU1PMBRRXadhmaBeRXH5JbgSBXVVI9otuAgDq
LZ2gAT/zMIgbBc05l7kypJDdirdeYIg3svM8LcpdEVwecwXVt2Z2OutM+4fmosVV
2MhY5inDVYiwue2NBbAs/hDfYaYjR/vHxcqCxw2njz4mAB/hmtdeI/7MlNEHOId+
PLY/XsVEybb17pvaZzCPw+lZP7eWjMaWhD5A1PYPVQJ9pZ83W0PNfv8jYJuJI5hU
CwncPP3ZIhncp5UrLMFRomugiOhf691ysZECVCZJBBxZooQ7SJYSgO4HXMY+UCPK
WPkNDOivcwvbL5A9+nSAPIAhQD4Xr1Od1ZHkqTnwDvN4cKHzBK2168f7G4Dxxohn
LKYGwQDNRfKkkIxw5sfqd6oOKJSeWGwek+//jgS40x2nHFiULOaB270KSj17dhG7
ZwiIOWdrjMjaliFDOwt51kXPjp025OJTQpyyX69tcwtQp/4hAps73Eu6BiUJ+L0G
4IMczhZNcApT5/KntF2l+ar8uFWnimhlIek15uopdL1X5rGwVgSvMpkaMJphz441
eSRPiBKPrCtg8O7iERmMgmd4wFb4X9go9bT1fy3MOaZMvtWRlOqett4WuurtJ9ja
4LY1UB/N+XaGKJOwFfZ0x0z/FVK7wf/aTkgwf9ugWC7h+6jJgJpfKp4A1E3YDEPO
o3SGF604ACjproZMGkDT20L6MG7r0uYjgY3WpY1EKez6wtbXzZaHTjYegVzL6+4f
CxpWENyI0kSIdOEXWWbx6EXogR/pszkIBsEGs+kvmg6ioCXr1jYjq/QZLHa52XbC
dusYOeT6LyU0Vyp+TCr0IMCfHHYa/GkMkaSMDUDWDol42g8Rudf7bHfLgJ0BhB4u
73hPluB1w1fH6lnsoIWnkJXTp2OL3pTza7J0CgVY4Inv6RnDOZXBEpEadE7VqQEs
i7V2nvMUSHp2+iyThA9PNiYsl+Uf76EDGQucWDfpL04+3+Ddmbf0pwVYPUwxhKv0
tAuhobI8P6chWz8CrGx/2SptWPAus+yajkai3oPy2Agnw0MGb9bXl0VGw5YtvPth
vlg5AgQwJlY/UJWlrIhf2SJ/stVmI1DrmM3eOhjoUcDIS258N9mZhALoWTDPl0t1
Joh65S5ZmRiJM1MyfmIeVcplfGbIFn9DD/NyRzWOg98wOTQwimCEEME6WhhK5Aaw
UovxOk9VthjnrRja1di3xbt9o0yrSo/lbKFaJD0GUImvPXXFYvletfkhwZyh3v8B
kiv3WrWweh/8zuG+zfCFDCx7rDXaK+jUsFkf+xa69SSszOIbyKbgJ1WVdraqZXeG
74NnXwRNS/GOlq89ox0NUOac5pNZtjonH6h6OeofRXzQ+O7uCQJi3HaohpEjCXEJ
oB6dULEoEffpcWcWM9LcniJZqwFRMP7M8GKssel/Sb4iRVa4eqoLo//vgtQxAVvT
V2Rc3pzGKIs6M9GCJ+9DArtQF/Q8o46l7RMWjFXKiTf2686qTUOJa6bt6psoQeq7
rf2BKq/Lgyt4FaXDf/eEn1TeV67opPryaAmfqzJjv7YGHCbY3l4uYR9zba6SWphb
7MkF1xc8quzHq4ZmT0VIci0PhPZ2R1KuFI3yF3s8ZkPA0KZzYMpMF1yj/Cvlh/n2
zuezyulEBMPibBNoOGbXOSLaW2ltA+L9ZW0T8xIBcugIY3aSCbPiixu/RwiarvTX
/1xItI10By29jWLcykwG1pVm11w+jfHFRjVyqFbvPML4fFjIcHnQIMmmAYSUj+8s
mnYDJcRbgGdLGat2tnpKcAXKdlqjSoK+YRgxhO9qZ/+OLoD/Twr34pCh4ZRTnUxW
ftgjicXH6HgFSBZS6jej+SffLg0Pgw4PmMhN7I4bcRaAQw/3EXJhT2aoX/aYU5Bd
rssJNm/GVBkSTbjub3xN6sN3rFWDxpNXxxAy1qcnltDzhbFnPeEip8fCrrspZr2I
Kf+KcgexAIkX+oJUPfZrxt+M5jwDlqdg9fe+l4kInVApphYIckdRxjE03+454KxV
0OAJFKG6kQxqbPhRIBZmSPpQUeLacTgy+qt8US9smXez64/2F/MU555reWtwXTln
wnrU0Xg8k5iL9AfQIsvq94UfsSKN6nImtwwKRb/6WYKPgAPbNqFdHapnj3j/GRff
80ZuWpDounQWcpu/84wSppM8aXvMVDSVlWoEKkqkMlAXOUz+n2J6H44lhKb4BNaU
v/86RZ1Yd5DxEhmJ12EwINqsln+jFjT4MyhmnBjQ7ZkUKFdYCAaaHTV3bjAWmAs0
kUymlU+XFkOG03TfllJ5wmkv+6czAGIryWnlI3nVSMTO0dG0D5dbtWOZnLb5IO8S
88KgiEdVNgTurqrnIeIRwCObzSmh/5JZlQTMZxHm8/wnLJnjSLGCNIQUKHS+6p9W
2N956Du0z+uTHWcN7q7ko/RpPCPTq/h/C+rDvNhg/VOJ1+OB2U2Wg2A2XuSNMb9r
a7ybV0R9TgpRgWPllU4F4MY8ZnGF5gjoqqrbOm7RIIzOdc9qcznGlLpJVeJOwPF+
XkJdMpeuXkznvr1ZpKAQdry8wTu8N9/KJTczbkFdMUD/Gm2HikbEeMWgEG/fvqD7
yIL1oa/e3+KPoJ4Z+LucaoGtlTMUuaVMX74gTYEvlhEE3E7Y22OhfT5Yn7ZbjcfL
r0Z6IbpIN1R7+6u2fh0EMy73pydHyoJbqv+ZhcGfWRMvPNekKJ20Yi0l81RPo1ec
12SdVpplrft07LarK8+X8kdvEqRg5TohgEiWy7Ko7DsU0HMSCVe1BOS3Z0ksbij6
J6AZpWsDjrrbTNcjEJBzLalC60vEztjBTGuOuuWBxB8dbdwlMPhTWXb5nJzMn3xM
1/GynICi8PKNOulg8fbXQr1mZHf0Bvr1p6XpQntgP2wDe5vRzl1MiutUy1TVrw1g
BJor7VuBdVyyjrNuE9PbA1nWZP5cJfxI8Hp9m4bOLD8GKNhR8OJ21BKdnrihOcwU
o9LysH0RPZI2MAEdAQdzE4HePw+yl1LKtpFcTBMXExR7W8rHgWz/wrkTLqWITXI0
3bRP3zEZp4bxZvUc/D2L7W1iIxcxuGcpLXno2Ign+vy5vysRDgbxoEAll5IBYzzC
VjijgmWghXpPfrSkfq89pfmPgpRC7dZQPD12rNDLFynmSF+zYCTT7vBYHHy2pZhd
6rv9aI5YxHaeywrqFe5mJjbMnN/b6XND/RmcN4yT+NVl8IFvRpRugHBv4i3sy+5L
lrjcSYaQiU6SPxe+Iimr2iuHv1wQfUWBQXY93QgXIsn9PSXPTBt7Aen3rC9nZfy/
ZW5eTqQjk+V5GVmf6KUAF9dPQyszhAlHOcrhVFEJh6p/b3RVc6gTjV1uHwLdY/uK
2J/ButHBgeS7uutltRFJm73zHc9hmOxHCIHU/vLvwtYzFd1WDJB0dbSKlTyZhXSW
3ma3vjYnkeDSWA9nkTyTiTuDLbXbCSMnzmZiaC7E+vAkB0gl0A1lKI+ilaPHcTOY
vs1ZSRuT8nSaEUcKNIKUUwkL8fRZzhLEmB6n5IxyHJXb0/f98q2u4j4n45MYVpqi
8ev5CylyQIfC/OQKcUxbZNqx3vg67op0QUDeqPU492hz5F4ewTeteZoQHdL9aNI2
hlET0Q1AzDAGhcay4nkmZDXfa3KGV4wKhyVBHhqT9oSlD1epmiccLQKBE9vjjIm4
gpdOLhM2kSqWCqIQ4XE1nhyLCPl4FShOT3YxD86KVP1/jTF0ogEckE15ZB7GsOqG
Qrvtb80lALdclR+RQ7D/PkY9pyIDk+CJgy/vCEWGhxKWcSGlKGnttDJoynoFg5LL
QtR5tPb//CZccRdypUJDnX48P0J299QCCIUvfHQ+YX16Kvfngi9yvP+cSozhXTIf
oKzzYvnjVLTUc59TyOjm7szPL/h5/b6NCrhdppnXrzahjLl+uOa/6mmFTWwuHuH+
E6gP6DA2KIm3ZS0He/iZMHAN2chgy7n7b2viBeKBQTz6W9nn7QIbtpLOFy+bjoeG
rJ4qkncf+WoDUoZn1Us18ONKFmdj5cTWzGQjZOKCTUfYigf2tSgAImDTl/Yi55Uj
9ti0X9Bc6+qTppUPXfvJL06NjuWNmhf7WBPwIEeQq1WOL8xXoPfJ/pnhV7sI/jgi
dMw6Nl/mxdQj3Bxuhb6KUiUg6IcCZ6AajGDTofKKttgdoMkcTlGWlSXwxTRxGgUv
D84c0q9o5ZwqcO6/33PfC1OyP+GFTDs/ZqhRs51vxgnw8nNEbabtaK4fM345RMSc
+w72/5G9XPcciom3M3Eg/cwy035iJ7zEUt5NUKe1sLy+Fb3Yv/f9YOx9J6feb9Gt
5z/HEuU72AYkEzxf7ljvC8uuxwkHh4MGn9aO0Rz91JRbGQOEKxAvGCSlXScRmLED
2cHT4g700zLigenAAm+Ic3RJ4vcF+17tirCUCA38EKHsUqm5akOX9P5pCmG6k5RQ
MH92fMfY/DgoERA3QQ/u2ANVf3ECeolXOnat6qIy3VT/VHVZORFoTiqgIcj3FBt/
9UQXA9W+7olGggtjsLGjcarPATEs9XFvbXH7VbU2CWc58odCrTyuZNcMVkclLmPd
lZBwHZ7fC5Cl3i8L4idJpznngpjwPew4dVPT59d3L5isphStvaph9OYxnrLYb/7y
aRe3vc+oYtlVbRNVk+4ztfg0lbgP2SNtk6Ra+7cYAmgEZ4qLI6cdQe7keAlKC/rY
FoW8mE4jb13cc+hRIY+oyCSw6IpFb/fi4d1xPI/wbNrH3+ZcTbhxzZFQ2AWGZ2Yc
Bu8V8OOO1bc6E2atetcTxva/9lL/UkiV442gSQu3bWKZZM36roFCciwXajPlfIPU
NUyX1OJ1xIbxTpa+uw1rx/Fpl4SqZpV1w++1MQEvVJCzKwlYD1+zBplxrO2C9eCD
eOpGAfcOVvFJsmdwyz6fuZ2IyA2i1iBE4O8uwoL0GLxJuF2SqSx3L34Ii8lBeZas
y7JGyDXE/CY37qCljCwHywV0rAoDeh8C61RPeWF0RMIaaEbdkF4h6NgMi63KkJQw
6iSxAsil74Tqo08LGkncLgATaQsFHVoVlMdDAfBblEV+k+g3dZqjlgxMCzc8r9xN
/WByroyNMMVu+AkfGNB/TCfNLWSEtFDbapsjk+1GQRwGzVQbgKmMfaCcnb4loaDR
lni/5hEDJIG3nrkSNCP7jdRiOc8bYacSKffWVX2tJmL/J7Oog5xhb6MdFc60SfiG
56+Yi0t3T+zSxAtuDkPNVA+U9bWgvW/UDb+eWW6wbY66TX2lewKf/mH0z7tC/mZM
65cENwjRhBCl2H3unb2abmXLHGj1wT+8xu0lK7UV112B+FIVZvSTqiZKDCigVm2/
LKm1+X29JQutE6QIu/CFCbIfMDC7q6vUfZCbJTMl1LqE3JFJPt6NYYFUOgaSX19W
zWJnru0b5zbiJh5eFmugDn5xQDtoIl9BPlfZgig28HRS6VUAG/btSmQsSj6YzCQd
LETg4WhmJC8qs5t5EBQMejHUuKL4MsQQq8IKkdceBLm0dgFBsrpK9wZhe8aO1wE4
G8OG8ncGzLf0V9px1Jc7HWh3sZP6hL1EhA82N1vvQuvV2pKZkkpckf3udW3dtXVu
Htvwq6dg3sF+J0Nb0diy6Zk6UJxV1JOIXWNKF/s+mCuRqHgKyDrPX2qKK2jtKN1E
aG4aFKWLBlGtQaPz4Gc/Ewu1ezskFZNZtpsUVmIkSDaOzWsIa4PiLSvUozzuUQJw
NtxPEtBxtYbpCqYNHCRV4c0GhKm2rW30RRTbc/H5jEtnDeUmRTpDXXtFlJ9LIIYI
xz+WcXrk5HmoS0ftDUGHYO3n6CYoGzd0KHWi0gJg/LDO/DKbHBOvQajX9ZETlqgD
W383eKdOHZcwW8dGD+LaFHMb6uGITsvVSF0bP6gQqARrNTLCwcNI95yGbcNBA09B
Fvo2qb125xABDck5dLjObqnhLd9NmCPHLbqie2aqX4Vx6ZUM9t3QWjuR8FZ4DFk8
rA6qAshV/+zexfzzu9UTVcnn6nkg+kPZkzXXOZqorMVBuJRPwajy3NG2l/377Y14
TUhUJQyyqipudciCpRtac5ueYul0mrb7DGifxel/ROg/Kx0QgHXmvGB4JQVRUe00
gPyesOUvWAqpbOIm1jQ1ckJ8+oobES3lP+LojWaKiZ37UNLEbdpWz6WWatOdjy4Z
+DJDvN82x1if8s9BPsSQL0F0Df0D0xfFffCv45PSEzrWwDHcRX0uyu0YDeOvWXS0
JG6ZT5GRaSSIFb/CzYu2c7MNSkeFPnu+zvbgN6Ige/6I7Js3IEtK8vkoYbMXRBOy
sSzSIf01mThBSNuZbh/kf6z6eEdOQNtMXOovBzkYBb9M3UalnBu2XzNZ1+DHd6HU
RsEe+w/v5ONIlBusuh7GK8Mc7vJ91cTjEpQZjGgcLf3EpyVIREsCfZfNjsM/BGaj
J9bP0mVVpVGK23yeih8Ik2AMQ53bh1mpcvLTGdsY1suVYClIfKJLr97v2Kn65/8r
HKehB8ggHRtjTupqkYw7WEGTmCl05zA9/KsN9NixZ5UeBJpyyi+mI2jR/XS/G8j1
GKYDyjC1yHNh+P9X5lLDnpbKgq8/Vpyv0CSG+weTgZdilRexd8SSzyRBtnejIYj9
bbgVSFxxMD93SoUFTej3PM6wiGZigYGx+Mz4Q1rfzWCy4+NR/PqDcpMCPoDQuTPt
mkbZUc+WQhaEQYDVTrnYisMf1ENScEe1wRmlLIhF0fLPsB1W1VulrcFMpZbHLlzG
q5agMmbgb10aamxPHLH9dzUuQEM2muOO4ww9nOdgKMYoh/mOkyUuWryOdTyhpD9S
epm20DkiND73NkPJVesqL4W4ehYulRt55Bneu9gs9A7UaIv6SDATPGM9iyiKD0fJ
JjtqQ51IBsCqMc7tGudIzfJwKeYEZ4AI2J6Pa6Gq6ha2IGAjgZC2s62daRVEY+iT
6XuYxeUMVk+cxF+ZlJp1Q2gnBUIQkM2/v/AGtP7DnkmFLARqvsZMrNtaT7+S2MU2
89KHIyc8gWi2k+M8y0kOHlWuvsywaR3eFzPj7o286zygItPO4YEaIQX2iZsW/nfT
jbuwmafei/ZQRN7Z5Ww8v0YH9brL8/l6Ab8Bo3XX4kxb28b5FfoiSu5HQK7m4Hfs
6IfNUMOhkBxRAtrXLIjd7pjAj3JE/qQiqsmdj3Vyd98aX1EQc5vI21j77xgw0CTg
zey63pyaRYv6NIZEup4MYg1CZP7j78r+vF8y1hFSbNCihD0ttGRl88Lg4Z7cQp0+
zR2HY8RJH5qnZlfykg/ci4dz9UIRUupoTCmLA/qmDpottisHvb24nfVdI/CS68kd
pzt5MdnCnHYpUi+WFkoixU9XhZdUYAYWuxM0lokVVf9YGb6NlJYLuhbuLNKjl5ps
jxKU1uLN6VGixM2HfVZbvGYVAO78s1rckV8JBMNnuZg8v8h5Y1jRWUEfAAOFc8Lz
C6fhKb0fFeP7Mk1RcWRhLeOfoAXxJXOyTkgU69h5Wmm2d3SxC+Wt0OSHCgLNzO61
eUDzeSHqs53A4h0a+yN4aiUQQ9qvmeCi3m8GYxqSe44Qj5+eGDdPIHuzgoBGBfZO
6WJEw5NF7uiYHVg08EOFu1TeFAik9BlOOE7fE9m5PL5yphqYJAxcAEig3B+q2TIw
xH+hiuvJAgAwHqZOzhJqQOCJrycT8k/MS9IqtE7/svf2IL9EAKGhjOOTTDx+BC2H
y65SLTtzFXvpK4r7IEPl6Vvsa03l6UPG78tvCF1vzUfB/ipGezhbwkMY5WA+eS+Q
Fe8vCnFpqaW2gAMNEKgEmaxPmfvu7kcfUuT7KQxUfpY5MFTNj4EjIhy+foYlCPAQ
8boApIE4EUEyBGYLY+QjZc75G1zBIHNywmb9J9OXG20K23Uw22fz7P7S9UjFY9D/
no48X+iEjGBYde0JCFnLk9lyciqrv/s0fDvQL4m0NMtKGxMBdx9imAqVrTlD8LO0
TREgSFukeFNSPW+o91KfFYVeixDTbRa7j9oRqzSuekWG2YoA8e6shgq/zell0dOe
QcRrsHqLbCpU7Tc8FJUYYbOeqiOYIGlyU5YpOeH1NdVC61nkHRwQcW8TEc3+ebed
Qo2mqZCbL1uV+Y/5piHn6LCno9uirrrNwAAw7LuJ5VXP76WjGmXnp/IpXulNPKbQ
wzCyGq512owG0kuTb2lpE90CsJezr0wtxrQ1VL47Og/v8yVPTzaiBmdB8MWzwIds
VYjRCYOLC2zk6WDBTiz2ugVWAVW7rIGN29IEg62oX17yOyYFkYHGHfrKX6I3SZ7j
lCR/vv1r8pU9ZfCfDouB5kfxCbW7gGAKLNeASP6AFBnu3jsytkStaO4mxxIwILH2
kt0jyQ3rZgl35Ix7qGdS8PCsfcxFE62FEwbdLNuirrlsF6rxaXlp0kXz9psCAtcu
RgZAUp84ihU53pLVoGClETBdIpYYx+s1jLRKLoS8ZCLZQOx/DmQEgyvax+aLnteg
WeXenkuFT5sCilrgqqeVGi7BQmtR29pry33gnEY4a975BPWzevvr7NfO494JrSCq
IVzlJjwcbkGdHwfK/oBNHS7xcUTbDg9tm26IYlcXG7aJmnBVJbE7HJcQINgVCz22
So5ENvKKHPaEWEp+yEIK9t8uskuW4OnUs0k0rPS8vZVi9sad+nmGww7HcJoSWAoO
BQvndVANnWJHG+n4filbACF2S+jV8I1ga0nXrLZXOm5qnWCZ+hDy6eWF5fSU7Ae5
NQx39VlqCV4JWOUjj9r//vx1CW0CsWoVjtjz53rjVhIig41C1vEmUKqQRgl9Q0vK
pMhSBIZaE80Yd15/Lsgt72wXDB0hD+wfII9klKAnml8GLZYnK1nrCSH1U9SKCPTy
6nTyn2DjtTInj6Mfj5Qh5mQ32LieNYajQ5zRMDxiXpQ19uBsldlOHWd4WyezOUk/
U2Vz3szKJC68YAWP6/KjXyLEU82n0U5qR6HYarheO/FJlyrm9aCvpBIrzigeUHvZ
FK2Of8KvfwuIa1K8i8D6ekjDK15T/TMs/5MqzZQiN586GEuH1C6eYL9JIfJCcEK4
KcsvQb8jpSslSntRKO1uHkvlwaWIYHE0fM3YODs2x2ou1fmux+DwrSwElYwvgbDA
YOGtZnVl5Ekm9mDbQbCle/hEv1MOVt6g7eNloibThs1mZlVqTYNdYZvCdtU3T3tU
u5O4wppW3JJnrULz5dMuf392MhwYrGqHBCDgsEFXmZWtTE0v403+aBVy29f7+VVx
VKA4AoHwS5x9pLV2UgBF80bqXGAgpM2kBa4UA5mOPX90ZLULMoFIsqfCPnBuJ3Ht
cUvhZZdZZPdl0AHIA3So10iCSfKpndkv03nI7KH9Aua8+aXTKKuaB1Lnuq849aye
//gvt3NqOQfAB+BrvaAeV3WLjBeHU25i6/uXL/EnO0NWH3qhM4to8eRyQPFqQA6G
oUQxi0RCsyRBiiyX+56gp7ooipG+K3vD8Y3CsxpKkfhJs2bQ2MVd9WDLmnRqQcow
hMacJ3ktxLzUuzI/HMiXheUutoWoS30h1bk3F/wDvrUN1xLz52aDdMUpX298PAA0
r9l3bo9nAl1saPNP19/gNKEqAfwK7ZBDevBjrVcj+YcwjG0HXv9PBWm4klLxmiT4
S4yrwSvzq1+97Sl3ext/SPGB8zuJ1sNAWlNjY+d3V9kjPG4NyptC/rrGcx5+2Y+V
je7+9FWzM5QBkller6LZEir3u84I5C6w33Ct7a5VYHaNU6y11XELkxa1Vg0pJ81R
TumdT0WYiOhQooHdUJ3E5NothHlyrSGDcqStt55FQmx/m5CBvNUZ4iLkqH0BMLOz
D7REV+B1OIen2kyWCsV1KorL310Bh6X6pEF4tgjP+UbNuEulW7GRjl59oO/5IMUb
O+JY8V7zzBIsLINF7Bs45ltK8Y4w6VCG+qwWNYUqwT6C87QkLyzQL9kK6M+KVHzG
fDufk24nGB2oRsK4KS+ixjqRerO+BbrxU0fn2t7C3PBFspmnlzsDfndeaJCo2mey
B2lh02M7YLH17wX3NFlYZ2MGXLCdwfQgG7qfAouIGe8MtjOZse0W/965tJPuqarx
vgG5PwPdlGVIMG+r7w7vZwxt4x7/2qcJvuMlCQxoPdNSfDADEYd/9RmZ3ddGvScM
EfFt7vQ2P2pxp4RJReIB6ciR1impvOWePQmiKkk8kZHCaxitQIZfQlqmfa5kHrfr
8UFk5iKH/eUDNhT/JZ2+x4pKQWQUeOfXhR0ijfkVmfMND60oT7FXAzbEphph989J
xipBWIEaIJykMgbE9xmglTybyuIjHZ38gVXyB5CtHb9KBXYkjK9I+xCNdiV0I5Gv
yopU1GlwaoqlkvCCb7O/52riuYnbd4lIUXJQ+S3AYKb430nauBg8qyOZIGDI+o/J
3QRa5NclaKypPPP1Xwv9f/JiBQ0CzXC1jeKGqyUZ9P7SORZD2RbSIvQoHi1qukf1
F/99IeIIOwFoKhhpKF7Bi1sjM0Fpi+tpmPkoixIG761gT8SDEOQxjtI8ZcG2fLkh
FOrsKz7XoFOdayEnorfDwPkkGEsGYycC82YuxrOxr9y8NLyPHSWBqtR1tytO4UQs
JwEVvxv64v3vbz4i4YG8Q96dnd2DPpqkjzhGCZvUySIaejj9s5HODyjB44mLZHDL
6IiAErXMfC9WeiKIf1mGcPQwyGr9TA/y0w81FaxWrz08u3dy6DxIVNmddf2H9HmM
sFxXDyaXHOLCxbSg2sBUIVOEquC7/LZQdVW4ueV3A2vwqjRECF6P2igoAy4n6QHF
4qV3aPb6IZ+ZHMQFUrYVqcv1oDXJnAERJoKlLNPQorCC04hh+XhZALUpFanu2fji
wAezqTpqtC5ofIueG+12FxaYtameXRIt9sEMBSc4gygP5oAVB5HIpDSzwSF1e6t7
7IZpWujyBgnBdP2JnEGWegvaIjkIFOZtzPxXDFFb8vfufXFhpolIJQNMLQn4wGDX
d4wqBZTCGzdtHH1y3oYkdgphbsYlgbPvcZkATuyVAX+VpWH7F8VmPfKxMU6Qfib/
1f8CdcMSpReQSBm4m+YcjV1szOV6QM+2MiHJqd2p7QChJFCAyBDnIIh/5JmCA9/n
PtfdegzcaNWdMnecmXzGVa6s2OqjS5+BZknv1TmlON+Dtgj2UpdlgQjzJsul9H6o
A7dparcbhU955HyC87/bvh8vLq6YrBzVWvvk0CEjvmW3J6/Dp0AoMkGdwV/rIM5b
tIUWZFVu3gurae4stKEhYvStwC3S+r9apJaz5JXB1rS/J8lN8XxnxP/PPAv/OxJ9
I9ASbpZyPsnVnWUMtJHRZM7+obNgTS+TlHO0SS0cym9cys4ymBzYG87ntCeka8h3
KJstbFaa2ph4yjFfzpI0Q84bVTY6yV357jMBl2WJTaWek1ZGO9E71rY/hwLcLnhZ
fBdL3f/hOV6gmCWXYdB/FjtAeVuvo+G8i3BR0KE+SDssQbsMCnMcsJDPdEmwbk1k
YbWv4SjM4zaipXGnDk2HCdxWq6FOopJgj/8J3kY/A35gqKqfBfLMcndVwercSeQW
MdYfBLocCVb8pL9izanyp6NtZH//j4kFxbI6tXI7wTwvnpp18jE8emlxUKeLgH45
VfW89MdefRGv89ZJRwe0oYhSjrMLPXcMXzPtYrxjGKyKmWFeMjAdpEU2x6G2KHEK
IVWI3bBijs49XmCb76jSqPIqZdtNnGLT1DGYzty8Q9eHExLyhX28uDuxOLCB6guv
xa/EOX+BN0+aXN5Xp97PMkZ+TNA6nhiUa+s/zxkMvT8Qr2huBbE45JByTseDH32b
adr+fnDONedE7oO4akpyKxuo3K2okZmSkl+f+Y4Y50zxBCuaT5//zHYO58f0UWDc
geCKTJcUGOWvqgi12Uwr9uXWHIj5/XODFhsAAHhKUpKECRNdsYWTs/wQaqkBYUnD
o6cbiqc/pr2eE2VuMrYF71dW+0zVErCP6N6QhvXJWm/dw3tUeSrXpoy6jPhNYQgW
I38WKsE7H75ubjIpT+WIhYF6VC/4fbXkVxPrKGa2X8GcxMHgX7Nvhp48025U4FjF
Yo+HcFNYAtXQFGhiuTj8YHITyq3u4yGsgbrNqne3P2YcGSMiiYiutbVeh6q1b36a
IY1eHUgPLmfUtafqKDO3ovWez5zs3WlLo6o7Aef9BNLRiU5nAfeY708lWto4qQWe
97BX7Ts0cT7nkL0p+l+aqB96NucPJ9YiMn+bZNLX6OCZlbiphhhAszmn+ZvT7vgQ
NIiYJi+RqyAb3H4S+EYkeeCs2+uiJyoh0SbfVkGTSQXV+04f0apdMg+uwk4nDfdG
J9fNedUlMCCw+D2K5erRWv2s26Jrf8nk0h62Mvw9SmWFNKDQ4XjyJonj8A2/SMfR
9apztEsIS241w4bCElEKzt39MG1ht+5IMjEQsTX/y0JsvEZZ85SejHoDwZyyEWZd
xt/wpJakNf/3gKV8SnBjSgX/VzOAnNU021/x6YVCjeGaqQCWb79Jcd0SIPW36ops
JrLwqlNoSsl3uOy3xwO85nT4MCmG9DyVSnNE3HSujhAS5AKCisHsODfLKYnY/OyL
LoZsGfXCdLnjBpDPpjCIl79Rp7GVFzy+gKA1SDaCnokdjHzt3ZTYoMBFu0UDbdN+
LhValulkCzI54vBOYqlPJpqbq5RxaIJyaTekr32vS+SAq9DISvnD3TbiIg2AuV/Y
GSdYII7roTokR17x8PHA9P7yQAGBCBPyt53iNwYldBBcYKPKkRJZxt3yeXPrNJXe
HQpme67rSWl+/CV13NE8Dx5l4+ulS/mb/BZLJO00l9e9HU54QVgYBLdcWT8ri0+G
0MnB+N5S4ctKcRdejNYVyuz6lwTxQ3z4lW72SZ+ywt7kylRcFMeHUWmN31Y9RbD9
NGna0SCeWZEPQ44hiUWYENa+mgEKfIWuA0cvo0Kc/bxUuNfxcUgXfGjGlZjN4aSU
5Oh+eMdNIaKB06fLUAawf+4KqMh8n6P/zYYe/VVyLHzPxxoVXB54/OW5C6tfWk3K
bjqDBAdLkT4MHLBd1gJXC0C+Cco/fjIc1OBeACzkI3+aV1sdQ+5ZfT3Y4xKt0gbe
/u3erCNYK+EF4swk89vqjx/kVi3wwLKP7qnLxQmSo46HrD3ZoR1ftY7Ofz9xTSyB
yXua53xBz43l6sX5M3t7EjIxn8CAi6fI3hreO1VI+GwFMH5IDfY0xwxGmpQ7HxpN
hIfSHGDiHDcOH+kpx86ricfej2vdhSGPibsb4uZ8289fXqyiqeFASgJ3sx0dlAiO
IaVho3e3NORS6DJ8Zx3LBU1tz+Te3/YPYn2zCuvj5I47J5Qbzxc8aLEDfcwcdeuF
0oi9kjtGeHK2KxvgG8mtIhxAuKN2upQwSf40/7rdpCygg85HzgStcMJ5DBl2nE5m
Korc4ShZbNEPgtK5pWLftCbzSd47zevStxLgmkr0JYS/vFWfXeuQjYq/q6ZyiSHf
QSShVrj3SLhWVxOssS84SshTPJIeZhEty3Y6WIeAgFwAwrPFurEwBvaghJc0Fzop
9Nv5tq1I7zcPKc/4YYVBzPUdDMwDRLgKEpeEeXCfC5ABl0PfyuWkaWFRXzxRDMAI
IKCAr//jl8GqoTWvHGsUruUVQGkACNmvc5585jndVGY+nDcvH2f0x+pD3DyLmeCb
e/mABOtY0FjBmcaAAAt+bzS73ijPlTDAc7pedetItXDXNy8L44SEKrxwVP3U3zTy
jfpxCn7xShqgZQjlAi4WJlV/T5iF0ZTWiH2HbKJtSxWBu5yfJO6fCosBsZhTfpLy
Bs8Mu7EOb92jKyTXJNF0U0gbRMQodpEQ2/JiuuiEOD8/Vx0xxkdX+80ln0FDpeIo
HWfcGiBxfA97Jj4+o8bXSZEjuA4OHwtp7zjhimn+sF2GGjQ4cHM6NzpLMMtU8hcl
fOJAA6cNwgEGg9u49jzgFshD+b9cBQtA0yenLg96ph0SydyXjFqm3GfFmOg2Xcku
7XhACLhhViWVgnybSFGlsAIlc68WOdi0Ca2QoP1WouXP6uxkGgqVIQEcTKxWO0lw
C1VeYfC1Fn/jtsDr0o7Mw9Yc6/5QPJaFeUqi3bq0V+0KMOUpElZun9xqCA6ALpto
NlIx9urZjrNaDhHXSH66lcZ2/+rqAcrhcc2vuTWk5X2/UV3YlCw0+FsQuKaMptgG
zaS10636WAqlnGzquIn8W4IR/Boc6EB+rajbqgunWGlA6V9vFMEYhCFMENPsoU6y
RgxN5u7wXJV/wcN5HcYOl1Kca+mNSlPQKhl6r7IcdlL+n1uSdZckzCs79eFQGduu
MTScUj19iOZ58Qf8OJFOj7bt9DHmFAgjAb38HqES091jlzAHMw2xLSLnxDaMrUyE
6quZr3mFTMIlhMFlsxKjTBx8AWr2M3fiuSZCNDMsue6UJbQn7klR704mrzvrzXuM
QliYNWS9CVHyztljqnZ1+den8xZjaRYDMWZmndnEMxNR5A9oH7gr45dcTk2ycMWZ
8PZ7zIIDmUBPreJZoRvy8kyPUxU4xTsumFMH7CN4K6EzAmkzSDXXmvfVYnr8hXxq
OjpzGgvddS988NrCyYunajfn7beVLydvYt+w7E0mFCmzW1NwdX6uPRsgvILbFLX/
wxwfBYHo2K29yAS6RuQpKpCcl5WEI0glX6iondO0PkO5hb/GtmmOGDSbbjxQRx8S
AKyMzzFWQDBE+ohFlDUwyLS3B7LttjsAuJSauBo+GbnZczw6jIDFjRNdmyMkKMhT
lqPp2y8PH+BRY4tiNFfYQNvkutf+kMwbFZM6VYLYs7hD4zdVVrcSCoadYAWCgyOF
2zJ96hiyBwfFJcQJXgVcoYf2We9mbvm8Dd7HOBTrnrOpf7ds6kugjwj+qOMew6ZO
OAJAh6VnGCFxDxvgshSa4y8BWXF21FDVflefNo6Cgev5ecRpXG0tQA09WqZmQUQW
XDC+j04GXN3jS+rFdhkAoYF8JDFGFHNLmaTCmtCShAXEfpVqdmdRzyy5W9JG10GT
gZz4JRNqrwBOX86mYSfDzSLHfRMLVapHZLts7vA5LwjM4cXujDV6777TMZPBa2um
EXmmswKUG1CngyxpdpCMTzYCePeI8p81yvdORGauoCba9h5Tse1UOqSboJxjS560
qnw5cwcmS0VgsrIAs0GQwPvSMJrexExh9XawgfKY63xP8nJXXa0d6joeyit6nq25
cRnetvNpdcjO1xbVjZbp6x6IyIKCCZ49N3WrlRTq7PkDt5ke8VjrmQxchV9xoUPe
Me7nITbtFnbg/xg32CMABCZ6OCmYpfdcuZZll8asGrrfuy2pkZLnQtAGnw6eoYvE
rsBAdNIWoQ+1HVZrDj8ZqTeA7bb/ybClOQ5IKRhjQjen3QPmQMICaQCGSDpvj9nt
4RO9FgD0BdbTloT5/gXcMnQTVD2LQPIjwJqFtr5Nu9b9qVEVvT/5F3i3P77+vOen
mKilPANZKg2vHVqBZ1UxeOkqzinjHdDtGRUUfl/576TgVc6YwYWJ10CAUCmlROBz
vJPQx1l7z/pFz/BNav9GGo0chbUasA6Ndq0xli/Lv59DnMsTEP7HM4EHCxQIpBtF
0UraqE+Ez8MtBwk1r5X4/+9ToYD97D9I38AhZO+trhFUMMGacvGl9TSHBP0QorZO
EmxmQga+6J5ywfpNd8nbSMwRa8sCf0qRhCfGlyp4bZ93QPsvyXQNY4+AaplZzmvK
tTA7fcgkm54AV99NbnvQdUSqsx5I/S+W1UH/Q0Wnm8BjznTuGehKBM8sf1LAqAHK
QcL3worxIah8b2msaYskz+9CAEbz591gqgJRTk0A/x98zbDWlUOzD3aZoKtKmKWe
3sqgxVkhWUQDwapw4yLYQUHnvQuHQIpUWm7v0HuMRV0Z4/a+nD9NQOjCrJs5QHhm
iQvCsv/EeoMkxQpqK4NyxDWJA7lXaoas5xPqjqNO2s00Zlq9cDAeCwtkmff+i0Ag
h+qrIKlZ4hbLaU6mHhBc2IhMyW6MdU7AwBuO7xHlOzzE0iowX7TVOvXKoBo/lB86
b6PfUFxL+UysG1d+3RAEQQApdE6urt6jdz69SmGXxroa2dUYxooGLZkuYda3TJBm
faxlNA2bAa4GwPwurXM28qROC8ohWzxJfL5NOyEA7Oh/yQYrN0NVMzNliQMbP6LY
FfyN7W+J7rghYadYNESvZsM6uZ4BD+c4s00qn0y+/Id2NSgGuENtQbHrrM+BaXeN
47DlaNgLa/66mVbJlE5wkuPP5Zpnp5b7q06nVlg4yso3niLzpQM/i18fEeRRx98h
L8ixRc7aVgYat4mN6xvKdH+VHh8CI7acwSdMEy4SzyXo6vtFAtTqDiRwZShCGglM
09wcYrBezIDDmF9BGDZIKQ9hYb2zS2GY+NAr+DkoeRK+EFlWKrVrXPbk2rAmr1Dy
AvCp206wyZydsTnJAhp4JD8I/qpYlim+VGt1EwRBUFsWXqNlPHhCR4Vn9div+fYo
uNV6Ln+9k0YSe/+lGP5QorzmWSTI8mljDcgGdRIaDxsAsOZ7gj2D7iDdps6TrqFN
tb6+GyTPrGN4hUgnBbIPvqH+taF3quR/LLsRgm6l2mv0aIwAFYMHtBbvEsZJXTdI
k/D9MhdhWzgrTxQUeDxAetLWmFla+8uh8xoltHNNKZYdFZU4I81C1e3+uMkVct7V
iDT312sH73+Oq75DMbw8uDaC1UdrNjC7QaRNTJh8KNG9GrO9rzpE83E7+dcjQ2RB
0HnKbeQ4+/41qyrMoydw7Ji1WBhUG6j9I8K+0OGpYt5wwty3o3WLWM/Gi/ANxgPU
JVq8uYBVcx0wDriGi8yOarRTEZ0bYgncywBzmIbdakGN95XccSZmCDkTkiiymtJU
L4UEdx6YBvqlkEYWR73qUX4tuJDhuEE1Dcx8A6hhCCNqjU7bZ5wZ9sVqU7xLrlmB
Mj6HR+03ukwRMwtib/JIK3A+YjnQnMN7cibhLQrdUlr/u2odbVQEhsCPWZ9kKg48
g1GlGm5zACCHUUzKIEi/oxJ9Ip20zKwLfHrmjCYaSbdHVcBwirqU4a5RsdeV3fnq
inO9005UTssz1/DU49tpbtb6t8tvA3Jy6jeG5qNLOAUy4flrBwesoxw/r9x6QxLu
ZMnbQs2Xakxe1g+sxcIHMAKcODovjLI5YoU6wG/hXPxU1ZZDkS+Qpxx6TKN2jwkS
i1DZRXU+2q9qsfguev/Rg75KLhR7LkVCGYW4E6UiS8IOQNLDmC7X7xRRIxsNMiC3
bRKyeE3hPeHCQ9BllAjHbhs6lcwQag2EadZVtNOfRmnpBMK03mI4CIqSfSJrqpSt
WmA7I/fqtsgg4l36OdQE8J7CF3c8SSq5jtZ2oMI5pEFAVgTB5XoP3jqmy3JlWefP
6aNjqO5DGO8xgI2ZwUUhtDqDeMVFIdwy9riOJcoiqFwZoKhyXQEc5CtgH8gvtjOL
GM50h90jl3PPSLCd0apqH6oxUJYDjXq3NdJu6PejehuS+/LkhN7z/ZiJpYjLTuRx
0ZoHBT83zzaHXyl0cjOux0BDgaPd7Mx3ToNP6sWhvFDU1+og1554Hly/3OYW9zUK
0oe8MAtsSsQ1E9JEzAyGXZRE9bP2yXgMeUuA+LVgARtY1NgluM+h7gDR4r3+h3JO
HlIZcKOxp4BTTL3RXCV8ZM5ZlMjCnVLE15s9DP2VxBSalBoMjZ/wnzLJDTsK2y1R
UukNHT0uA/6U6wJC7TtIZhFjY37sXNhb+IDH5SbMxJT/laOu1MecyTJjwU+sM3mz
A2KIaZkJ4UeOBUf16FQF6kvlIJ1MwXW2oCqJLZDhcZpcBFnC7f/zUvUHsfmJERwl
wsTOQIbWgd48C/aQlQh0gbfty3Dp3Wssayedo+C/JegZVRhkDkn8NSRVGpHgmppH
OrmYXTkQHWYh5Xk72D5u2L0AYI2XKFoR7pINMNmZZGYki/h5jDEwFEljfTZWct+j
g60lymNYpUGQ+eFx3x/QekkGWn9IyXylV77RJDFg22CBikVKTaJPN8/i1lTfaLOr
qQjyvoJEZe9q+NPbBJzdUsNhMbtwqciZNqhxxGS5QJhRCJc9wKM5HgC9SRY/QPqi
di8YnfRRJDeX8t7KM80NCSIjPw0dGtWYOZklQ7EMKgQ9uslESeSfb0cbXqTWc8qC
IyeHOjpckx0LG0hYFSjj3CkJ6PYrKySI1gzfmr98IbvDlPuyBhPJaXtOnjlPTtJP
T6lLXINVY4HXeXLWoHQ3+HCT/BxxZyeVdkAyQ/FUDPCsH9BevEAPwox/mw9BMlQv
vTRldeERl4GGnW/jF5yqpo3B2pZva8ONFjxItFVcxJiaUqMvDavjCrDs/xdkl7MQ
buYQs8S3wYZFzxt8sX9h4aFDfJOCH/BQG2C5IgTA+gFuqu49QUQ+/QBXU6WB0VpK
QvgqcrzlgP0DrttjoAjqf/gdYRqr3BseuQvTjfQME2DLvU6FF59YUTs9HFB4nSnX
XLXGFmPB9e9TJLP9ACgfxMmqC41r77YS7tG6HXeQmLEXOsxkxc9duRL+DNbwdqUG
J0Dl67auzAMgX1sL0wrnbAIxsnrbLAfLV5qwJjyPwSP6rhneJ7knIO6WbKa63XCj
X1UsXnoosXfilzUOQ1ulqWDXWIYGLqLp0CKsWAOx/LrY2XPFhoTe4D++5+NPmO8z
Nqf1lea7h0K8dCvO5H5uK4AB749/EgnECfrqPFlbA14fUDG+98OwfjlXut/18y9E
fqtHCIow3girNxc49uGid3pS41Qil9iAXfatuGcZtTl74WJneTYfVsOt0565pKTe
4RF9H0EMOe0VMo4c3j4cgpPZehE1ZH6/zGg8Jy1K/HF24hP815gh5zuAksrg9TLY
qWXZgSE6cZF1UWkWa4em9LOE8oz1AL42kGSa8yiwEc1R6kjFy4wGFyunQBDSywuV
bxdUCuB37Bio30R9doYbJtvnrwXbjNe1C+3qD7vnepbW/dL9jKs9dTtJxNQ02WNY
R+BwbtWEl3cvgwE2yd8KazStf9Tw6z7a8A+PNZZ2uc3W5cDb3obk3bSht0PZvV/l
s4fZeEFsPEdtq8W4V9BYlqZ8qLleZa6+/mvOF33AyIyz+H+2c5DzV4adr8v8IOVD
e9kx5bmbcuD2msJaQrGZqUyeS0FhxNUoWCodM7t7Ko1fiNAX1//9WbTNkbrZtt+1
wQC9+xwT0URLLR045FkT/3oLg9ND3srkqH7rvvdBWL9cfwixH7SnVq/hU3+lREO0
43xHTDFXLHDbhcxE3S1gJOQBQON7fwoiM0LlLvcpwR6aKYaAqD6NaDmSzA7OkKFi
+e348zKTGGRN8fZ0i0zAuBdsqdyoqPH64jVWMMeVP5WGd10MddytcWsUMor4ZNsR
SG85ae6tAaYgUtfa/gnT43OSdsRS4bwTXBvBcLijFwIgOsNMp5v6UbwrU2cO3aej
rOMqgGo6FOurbP0URa8fGJyMUBQluIrPFt+Of4yetw0vro3b8Duo6+/WBUeKGB4R
HY+6L/7zRxbAmZ39O4e+qjoTHR2z4rqa9AgTmSF5E873kBfPKEECF7BgzFXtZRu4
elxfkj3rsq/Vw5+HUbVymEDaWNZ7xBhhHrapfy2Ex9NDY2icjkVYjngBya39NLSM
TaPOMRseCbSTDIDQBqKY1lZd92CU06hg3uCdTqxStwThS+I33StxN/Ycc8KmRB5k
CCSLgxt8WXxLGWk16JpwhL/7Q7m10YCnPNEYN5Le4yHjyWspGi9nnTJhg3dvHfCi
zt0yFFDUdfmTejS9eY+UrupYD75Va3vmdPr82S9bl0LaBachi7Z3I3QO2AzKzFR8
SnrE9HWFCvWQZmsdS5AIcS8nJt+bBSeE0wE5dCwG2kLi9i0vqDYFftWVObsnlSF+
TAjPMB8GTBLaQGBtWrYz4mQW9/ztgpnjoZSO5t5aRTpqQhm2OM2l1jOuZ3IV/ILD
n/upmEbDEA64QloAfB4Tix++ySt9aB5KfWVR9Z8wB8FqEUIBeVqZP+4yURAnQ4nC
LiPnERxHDmakNRoiU6jvKOrJ9/y5JtzZbe9IEhMkFz60MG91EOe6DxEc0NPkrVBa
ICqOdnBCIAZkrjfKVRa4uwrGkBCri3sVTWF3IBKzW+E1wcfzsfAhw34PgcKOZYwp
1hVogq7NxOH6pV6dXAj6Dw/l/0qZoBfqrbcUnWnn36fcI8eM7VFH1LemNSanAU3o
28GcmstsBoOoYvZp/2CRhz7PUsPqgxJ9lk2XSoi8EmoBykzr3e13biUD774Gawxi
CZB/ZPGP2d7VnWfZCU/OMNRkpbPUZxmwxCqVddE8Ph9eo9zIc7U8E/Xr2Qij4CiB
SDZExdx8j3TcO6UTsBX1Ry8dlwr+GjEB1QZQw4fBwd5DCIIc1qlk55AzBQCQKyLY
MbbXNHlKfb/tAdvoJmpZevWoBHGF/c8qU8Q7c3ts9a1MGmfGEeX85ofkEOuenGRB
mk4QMaDICtps9Rc1vNO7trrMRpFuoDi8xVx0WEC2ilGjV268HRycllgyzPXWQh/g
Kslqjvhm72/0KbqokOlOgNXeO4OCDbVgM8yRv3TE7D77m7IAf3XucCHNyEAnNDO+
FyVCzFhwQWr4uD70DFnQIowKNv3OS+aG74N1JbVP9CTuZz8sa5I4m2cDqqTvcEAF
cU0wP2mxtcWMDuAV7beQsUcOu7NjVpnLtb/aEOnsvqvDXccKUQ7owNftjPNgecKu
lnsNaEisZYcCyLFud//s5XUuApMiQoC/OcHiMPt2AMh1xWaPumY9P0v+uiJAEJ1k
re219cNTRw6aSwIaHq/pzpBivvt/8VQvuV05nbanm+EQJ0+b1SSMMYT5wGU/VhXN
BI46AkmnJNdc1Ge5zKrt/ib2+mllC8kDTKR4K5S9X1HUtU6cCvy8jo1uwPFHyJl2
5kTWZEd4gnb69FcOHfWimc4jBtnfJaARNis2JWTRAbPj5FZ6lTIaB2fV16y+RDQC
pyygYrzNboB+0bstIy3Fw1wZe4QKhcDCJ5H0XJLYvG9blOI3iPRyAJn0Czgo0vjL
rx3L7ok80HzHBoeQbIK6nX6Cs2hguA2p4uX/Kp7LjTc8dJ+0/IfhXN3cDuClEHud
AKDWUSb3x8xgdcVYAY98FIpUC8s7zIa5VuavftCC2NOuabW2CCUI2HWatYyXwZm+
2LPP+96C3ax4w8rVAdUhWm7sr9QEBJrj8vcIaAmEGj0+xeYsO6uY4VGdGH2GJe/6
9OnOD6yMQSpRgQL8phqhruTpizB47rGKQHOoYuNq8cBkag6wemkCf+6a0P0Oun7q
EPSB7DPg30aOkWi200iR6/zrfQp0SgOUzni5HzaNKPaBs3vwefKEg2GQ9FcVf05V
pXNITyScl1LLe8oUFpgMAtbl3HZm4btI8eiWK39Zg7T0a/IBHdxEk9CmUsjsg9ja
dPGSRcJRvdHET59Ypa0dUSAAM+Rrqv58wM1ZXY87vq50TWYzjxbiDLHU0b/F8bzk
skkvy0va2qFStVHJ6/gfXrNGhM/EIu32zaUvIpALnM+wUPx+7sDS/oW+BSxeGFY9
bMhZhU0A00j/LwcgY1h1aVpWSfFl/bnlKIKkPEU8TP1wqofhNc0dfW+egXu1afbp
gsX6pKjRy2oss2NmDYBdXiInT6c9dfVlNggMQKxShxxtknakBU8YX1iyOuTTK2Nn
1tvJmro13dQ2Dod969K7qbSZ9qcGdU/DWLiGwgTB+HqNcmXr7FPypNkd7aKPwXWA
6dXIvdEzyiP+1sVXlwPnI4OTMdvVUhZgkrutAOC73d6iakGjDX5OsDwgS5GrYcUh
WwrwlGBYzgvS5llBxHfZDzUHP8swLKm7U4ERCPV8z4e43+NfoW5fiVRUXM//zEoa
E+IKj4wFkgc6Z0vzROxHa0g0QUmw8rsuGiw0UyZlCKXxZupcGXkpu/bo+Igdr1JW
idmnfOamK6FBDVqpHKgI3cLkt980I4W1R2OwIFDNeRoJ1QFjb/ortXvodipLKgrg
+8zTL+1ETOleWofU9oUR3IVoUevt69/zQjoHu5+HOvrLjARgAd4pQGLZJg+KTAGl
6sJ3UCi/z0XhNmOHe1SjLriEOj/WIylSrA7YQ+UdLyCXUxkBsrRQV52nvV+Bc5da
Yf+mTfSzuTab0+WF2fsI4nofBdwYPZ2JOCaTSwAT7N46xGH6L5Mp4mGiaDU40lol
vXk5+stCk0mDwZ2HaGA/iPLOafG9JPdK3ys4FW62vw+3v6bDXR+BbXqexUGX4DPW
wFNMdZhjc3RaXzmbR4IeKQIZXXd5yUbh87zWdKc5KyBkRUHC8TlhLZ1Y9R7XqUjN
J6J4I7/NjeviC+E6G8Lhxa32Re9UASg/Ato0AnFHR17iSEoSVwQquWAaguKbXI+K
n6s0P9byZK242z1fH3XoyK3HvOrjqePMMhkQw7K832eww1LXQttoh6y1MlGFaZE6
W4HtaGcJJlIhSd6m0Zi3M4bjOneFbkg+Y3PG3H2PrB3J/eAdpH9UtPLYI9kcL/Sv
9gkw1+4eIb76ktnFNTuNTR+/MtH+u7c9YyYQCono2dyvKGU/5+puigzXpXjg+WE4
23RcGeUL7NC8bw/IMqVafuqOPb1zvqFqrOEVKMnTdzfjUp8Y6D1sljRaz/biIIef
rrSEtR+Dy1cxbcf0wpmhNxmU3XxZW1ayal22nUwHJga6krD89wgJ+US9GfIdubFr
tXipNmWPePvWrQQp3SazMTnpDKB+MuS5idCLz6h8wFDAsN//g7/n7unq/6TqhkRQ
p2Cjl9WFppMsB/m1qUPxzfpbGobe32/eaTXI8QDyb+YmF4NUqD1LQiWBjx8mwMFK
TP0pvg8mIRgGMPpx/JSBZtlpwIHftGWCroJiXNqL8pftsbXgBQqt3IbdUpvrWa6Q
q7JHO74qVMeMkxxNDaYamhbkBgE9Y0ytQcsh55xRrhTEYIe9ys2w0qhm1Z2aSsFV
74pMqDCekbAutOP6iem0Ag830bH7aZkoYwdbv71EOazoB50atD473d072ubonVl0
6suAlUjvYJEv2N9JrwEvLux4ww9NJrt8838ide0+Z0IXFqbi+c5dAG+hN29tU8oA
5R9d+I6/xkQ5RQbyt2an9waj9BAbtrh4J9mXtLoH6pUXa9ugWDijSk2PgXzkq9ki
/DT2kJZChGB8jd5p241h2xri8xJvbYCLjw7EZadDsdC2SSawgmPiJbN/gDK7QKKZ
Clp1g+jE21wzPsW4H0ZB5AwuAkSTjnMEwmIaFDXPnEpXHPqyjwH4sd/5wW9wB8Ic
D0/jg6TeLIYjVXWkN0JMIE7Oa9eq4e1IbMbOooKAeRoRtwabofoHhXS4kQN8rYQQ
qq8yF573LcZL9HMuXtBuchZiNrJi38n1XzDm0j/3l4DlxXo64yCG41b2CDym4bCi
G0TlZahdac6Jn9lmMn/oXixN1plp+kRhTppLib40dGcC2hTBpginF3HS05eTXXG1
1MU3j0Mkdplzr6SwDHx9mdyzshqJYpGAPE/WvcAhsYKaFyzWBOtbAj3x9WZdOMPv
i4jAH8FZZ3cX075+JXYKKXN5324YnoZajHt5EW9bKTjlVAvI75MTPAM37qZyTA0q
fiKXkqOADpZapFKsHqS8cKwuDPsMWimacaHXfRYHBciNiygUOQ/tJtW8Cs1WzvlA
At80edY+1t2xSktuHjhb4Lkc3GOx2V/KYPqMEIbXT2N8FJlXd3pbnL7aW7Iho0Zg
OP3SnxdH6NGaCbnl+HNh17XfsG53LQYWQXl3xJarBwG/lHr4VyvZvBplAiTFBGmp
qIlMzsa6phnmdS9p3lIHxM7utkydrhuqrilE/aSErAMFMkFkRSoDXdZuGwxGTZA6
weGABZXEbkDGGt7qJygM/Q7FUzzjT77CiQ5fdrovh4oBNzePd5ZFm1HNc/3qE7ad
MvVUXzH24+Y70+ok0br63QIGq5ILf3hR8auwc9HSJhQP99nW1Fq1B8TQRN+DX7k+
SmwhQCDV1zGD8NZ/XvkRT8t/cdZ0KvT7hvj7/ARL2UqTBHLk2thR+ILHigsEPQY6
Xml94+eAGRO/xWQGgf6rc1WYoPT2AI4TBjq08U7FOLGSOgUpXPvmuEep81Z9yU7A
hp93FWGJuN74IZuW8APfT+6oceO1xTzfqRVcLau4WdNPMnH7ZYiV/QDFkKqWodz7
vwNbXrJF+wncXStGUBtDOS4HHnIdMhXOdC/xVCDrZXLIcpjBl/x2G1KlxTfjQq27
Ob28t5Or4YjC4LvvKMW19TAnwOchw7Ehzb2A3f5O7fHBANYQ/ciYJZwSVEt4KISY
zDdTnZS3R3CB+kY1fhIiI3QZDpfiAE6mKCD3SHZeZDdzouEcJlKA0PZjW4hKmV6k
EgbIb0bI+pvEFG9/c4cfIxIgrfJeYI5CR4eEmP+xTekDN/Z52c+Nc04vEnQ3ciBV
oPGM0qedeaXvFmJCam+m7OggcpA4W4uNIHg79HoZk+xCelwBeK0e33I4se/kOeQA
9t1mEK26+bOjnTBqNLVlLapyPz+zUOOM1y2fiYp7LSi6skHStvSxUoigOOLdFDaK
q0kBxOjWf0F2foCmuX2yelNq0S9AV6z308GlYuxLV+al3mewi2tW4JE8OsYdBkoK
4BOPlpsziqdOjnvLsps9eNf8DplqPGdeaZVsOjdikyT7Nh6xS83QeWRMH83G00vU
Gz/huPFFjQi+aRRH+MCNn+LzzHFgq/kmyiLGbg5viyTV6CXOlhOr6YLOCmdWm/Kt
kB9rl8zrQVphDu0Z/l8aI+JpdWsTTQTNTujZOLy7+klx9v5GakdxNe/wYryP3VwV
9KbJg8Ipb3yLMTxXyaBUpXnZygvYEWAFB6h2fJR8GRk2f4qNUl2VawYb/VJG5s5j
29bcDtwmbgbRg18em87M5DMkCpaRfU46IP/Vszy5nx2DlizrR5xaxnGg/hVJkUEO
Rnxi+OfW0ZPkzZbmoqUkFXLuaG47rL5QubKvFBWRAkcfeqYu20NV3A4yIpIQKffB
chYxxJEsuimkLToA57nZdMQNGduZc4Uh0pjQadbbxvQtDES8Tsg23w5Z6wQcTf6F
1YCBx+iHMBiVv8COrInXVoAGoqU+2+vC72FSQv+xGcE/YrkmDuOMjVTl1BhVAlWo
w+lo1d5tui0KEDGVSCuY73luU6bwmjeKXfg/p0Yc3nr53GGhJsBE8Slnp4hM7vBT
kvUvJ5ha5QHxauBpN5x8PZTJ0djdCNpjYGdKj/6CicDA5GDAXefOYD6RzELPKKHq
+90QjuG4HQrAIvB/vEY1KvkQG9ZkJvqUsqsoNcDpyXK/e7uLh77FAPvPAF6xraJZ
yueSeCxqhfzAjl3WJ+Uy7BZinysqtOteF/ZQVRLmXrltSG6LusD9gerooff9gST8
4JG2uwSlDc+PMI8HBgO08KCJI+KR7oxjMk5REZYcBy0zbaTj9oTEhJCpTSqBmYHQ
zhLm9D416n+ZUf05cvWfc3FAW8JDG5mCwXTEx32ZdY/RGh5cPu/bp3CUjEiy2jnY
xqCSFAiOWSvrl/OtHG+niCBxvUIjDyaYUKd0AclC1ZSCXbBwsnUGBOvcSlzuKLqO
hSwhd3f1KZQYuQwZR4wC+une9bmeJYuAaz1KL3+yq9rLlRYhWJzL1EEIOY+geqRh
FusQXXK0SOhl+W01b/vdlbbS07XZTg0K7Cv75XSWCOnFwTy2IrTTJqbbzt30IZvl
JSTEdIRBHltsN0zBpArJv7/mEzo83Mx83u2r5RIUNxEMpxd16vrLVVrkWz55QF/C
qk1l1xhVGZ8nhtmuB/SY1OEXVratMM5i3IhKSv6RuSvzoFXtB1Vvu0M4xv1Xqolh
I/NHA4JMKzcXkXw+7qfDnBSNd/6Qj4L51eqDv3SUHicsTWp7h/6JFGKkD2XZrCx6
zZho0YlB8zBpw5Bkw3gJ7n78kxWics4lmt0YsbciagWJXt+vJofarNLNkIun/z85
pDYoy53kNqyvBgXNe32ZZgbeuDOilObpMAR0XkOydYeF0seK0zBL2/Xbb2UdwZUc
kzKghKxkzjS2H5krgNPTrb9JguNtJWfMT6e+r9UgoTd/q1yiLr8Y16tb/okTvRH6
5LwuaJorvEuoHe9OEltnN8QSAx+26orksHyb+s7rQ1Kngwl7D4uXYuOOoDrD9Du8
uWoohCdj5fKBAympL7ujDbuco2SOQdFMnoWwDYNO3a4shrK6Rhv3y4AGxAMr5Ft8
efFN19H5E740kH5aYaHjVjnRWO/tgkxOavBldmnETnt5dM7O7JvvJ7/YsTAbPLXW
7x1ELsTntsnRQzeg8sLnW5yHs8mqY/4op0HN99D0r4U5quhfkdQJUYPEN079H1yC
qkpPi4yHWvG4e4hbDEoVRQy4QlgkVAAGw0CVJ0J2Mu2HHvNCAedHDRr+XwWI9Gs+
qwSCv7gzILFwjUoY9m17cfY/Z4sLt4xA8RbMYqeMfosf8TVx1qFhjCBDcR5pFytS
sqft0TpySP8TS1OUzFFAcQTpOljsGfG2jIjmfUJCGnyOOSxi7PHmfib0ZYWUOXKv
ejhXUdGy2oYDb29wF29EQIgoFrRzOZQI2vs6RoXbEhVZfmjNQHtFUoVHzAEVXtrQ
DzkKW4J0cdE6dpia+MdoPuTceY6RLL1Vgw9EboupKGyH2ACCip1+JAA0B/ISwimz
Y0kyNfEr6cOKUfulM4klAUDxefakrCG5q9bQN5DlxDPOsxmf2V5Zj107JPaW/V22
dUE6/EcHJOXGEmKCyWadBF1Ocv1aGgAqqg/3ZcN/gbPrPmvu//zp7psQFYUOmE+m
CVBaKHgAQWtXwu807Ok1Pxv85vbgHXLRJTzHpa25KZpeQzMafHjOGfiTDVowkwrP
Kf+kosaM6uyqvJ6QvxD/Xbix8btPEsXwhdOU4v1mvrR1xZoPeLbOz3Uj4TC/RBLv
yWTpXzROAiAqsfLY3KRW4bDflxdJttdKNA7EB0rMMlo2/TM/ctiYAO1+8cUmZEQo
M+dplfxjxvnFbJaJIllK2ae5439s4anq2CHKeE4BZ2FdszGclkFkOZJ8xlwB1Gch
CHN/tzRS8hQ7TWxJGmHUV2eTliOlpN5HM+v+eTpTxILHOV/J9jgUdBig5kDq54m9
jVhUmQQWDwc4+cY6dcT9twS10RLgPnJHJk16LKyZARJZ9BMmzV3JX+o6DTqZV5Rz
wX9wVB5z7H//zhu5kqhui6FwvTfwyaTXS/RIUpsTpbx0XSA80sYmoryzDByULeO0
AdoXHGQdDhXp2iNV3IUMDx9rDGW12dZbUufDoZQ+9Hwm/ZrnHLd0YHRp8clrbrwc
Aw6QbqU3U1+Icu114tdz/MYDw7BsxVinISVKvFOGNPuute20NIeKFTD5XoEvVGGW
YU2rjwleGbWcuDaxrKbFtqyBKGkGptTNI3jrSOiZixoLl0IOTF/s7PHYt2pbmSu8
dq9/7U1lXYFHIIVsxUL6oXK1txFJeXlV0S8RZGpmq/+ZS43TE+ep1GqxXRrPPWEn
Cnx9bOE61g1QTC9e07Gv2sizACPapcpBzAP9pKc+PbndwpImqjfUY2USYpgOs7sW
miIJThvkZ1GplfNIG42CnJxrweVX0LIiOI7ircgvTuqNN+ei+H1oWZpa8RKZyT6U
sOjv8Qz/e5yOK8jMaLeWF/OjI5VrUMxya6ggzDo3D1IxtpAOFvIfEQ0e60JjVY7s
DkRZCMQuZboqDgKRv1exn37CW+p3y7KcBiirV73lIzgp9tWNp4p2hscCy/Gf/lBK
xV5ZNsRBgPmpEznfpouB4jDYI9taCVL7ywHEsGLQ/lw3ITIF2Lld9A913I6IQdJn
1AIj5XuWBZAzFuoANiEQGXiUymU9Lj7uReOlJUjp+lSfUH+zfYgRAJajUlbIeoVE
y1IcrN7+qnKVu/Y2sVr6DHJik/iKRtP3YPETxc3xK8afGI+r9j4mSxF/Uujl0+P/
SzqXW8OxrBDL8kV1hN2iBBYVDCuW6kIVF4gbiyxNF5S0QVnqomZ5Ia748YEQwLIH
A6ohhxXNeKB/bPAys/Ym25GzXotO4Y1PhONLkR/BZYj/J44/4cj66R6GymE5YrBA
sUNTpEkzzBMSGDHMF/UGiDEstLWFjRw7+/9AcCgCzoEbW0lBH5fVLhpnWflG0q4n
oPjrA8+ZK9ie6Qby6K+7+4sxWRiTSYjNc4TksktVEHKMzYAthB6jyIsiv0gfnLZ3
eQ6kmX4WopY+4CMmTESn9qOAcLRy9CTpLT22SWXZI9H8N9UxfLVV4XOc2tYXcoet
oGLoBb7mpjRuahy4wHIGoz0zNVM5rEn+X+KmbyHp4RBZH9rmiYB1HzX+UnX0U4PN
q2GfFMDA8KWg/tR+E4MUC498UbV/UWvgVSoxpp33DcyAle7mbMXXt8dXUhivEXZj
OFMU5KEOg2l2WpfScAYzW48kcEwI9Z98vc0vjNuD2gysRp3khq2szsrCS0D29kLX
igctVndULsbw+ePOZUG4Zam68lMAHgeGPF0c+BFcnGIGC6WqeF9ekl9GGu1+ixov
8J+O4Hz6FJXuaqauq5EDb98WLI010ii6pEWg7cENY49N62V0qO72VAXx9XUS5pkb
xxgG3yYzkcqkdBipeOh0ZZbm+xPCvnc3ipEHYIzSu9xkrwI0+VzPtVLor7FMD0lV
sqxR4lhcDxGU6OknFfFK5ef1sY4zpUf+lJ4JkNcCMwweul+r2q8roOslsfEi4sHr
0G2i56z7QLZF6ko793Vmv6RXXrdbR0nJ1Sg+EMm/0P3BUXj57dVcD6bTpYHhto19
6JcgapE3cMjBIssm3v2z8pzEZzM1Nz5WX47MFPblcLA71cAZyaz/zTNaiuQ2Jge7
0J2Qghdi9czFZK/GyY9HrVdPYzQa5kOdd5KgRD7mHGW4NFR7VzaXPEqIm2nUdkzK
vgmkdqEbtMMCiUDfHR/Q7bLJVpkaXMShBl4b25gOBUUcEw172GK+VkrQn8XXB6O9
Kjuw44yXStggcTiZO9Z9WCDkE88IuseIoeiTotV0Ai3X7jSGx/0hNZbwhgLa0XjB
bsZXhRLC0lxo85m92bkhrHzqaRLWZbGFdB1TMyHDkKePlbIshyteDtz0Gjo9CBKC
wCV2nmpTeYqxVfaUiLlem/8mFpAD/HiHDO75Pi367fuatK1L6sDKvxaOgaWr+KUz
30ectr+Ye2FY3eUopN7yK7uyHhTTnIv2Q/DgW3PPVhkzksvT+m6bTzD/3mKPrKVg
q7PzdyNrL+wLwGWwGH1Vc/+GaCOtFU2sEh0DzUVlaD85EhclpopCUwVTcuu+c8zG
Nc4AYCosufVSHeQw0YcBaMauMqOgmHj6Ivli+vAdYSbqSN8YTL3XzeeSsuVRQqkO
einPkb4oKxHRmefNIn1IaQ9A4meIkq4f8cz9XnWGaD1sP+zGFtiTtjQpftLIA+mn
u2Jj81SRPOFe903WGqDuLrMGRVSiE7/jLDpHkdkgLhToXq61WmWX/5Ad6LklzhV6
nPQ9xUeYE+1XL/zfRbRAHjj6UL3/bxfvNTFl628mJekhgjlWJGjXIp8eQtJ82ITD
lGH/9TU5jHALCWKipCwOJyprfk41lg/rcuatEhRjICHX+IofOPng6pfLzHOTb1W9
QaDt8iW9OdIRzXXj7+pN9Fsfz8LFQPRszeHFpSvyQ5alKASUPNhePgTt614pBlJF
mIMA+FhM6k0YMb3JzKYv/fO0IwSPN3oVb1leO1wBYvDwNfiTT+R0l+1TE9R/Lz4u
Hd+ExiN9utVdFEw6Ap3r/hmB+IS/2Hf/lgpQ7MLxFILl5AJFYEWuM0b42h3UxZ9e
GsNfcqPfiJKLslM3O21tQZldY8ywCe/mh5UuLQ3TzPoZ89mtCYjP2e8X4e/bwl7G
wn00ikMsmER06YaB35oms2Bd7zBsTMkIreYY4CjhTbpWMnIPlXFQGTAuiCI3kY00
nieNCyFETMP/vS8f8e48ugUTMvs4TJ+qaB7WJ33dfhVUhiEryj/hs/0UD7YutGXa
uS4mIxXzSdHJ6RdVVm+54HzbKDAj4eLmpfGfNjdClaE2Ehuz7vwFPy4T9i3uoeag
UkOiUVjyiDQG15py6D9VYp+OnsW3xairLnxU/ZI/ywDvo3vWeeMU8QDr00txf8xi
4fKC0L6YtoOxTuIbeZVNrs8Ox9to8uHo8oM0GKMc5bVTEK7lzQw6Tu59bYoLXkvR
FcZmNirpaWXXSDqG0hXKhGSmj+ttRkmgi+M37BZLAiP/U/cWcEZlxbmgw700Ydra
sx/wQvMGk1AW95ZJE1xo8MuReNi7R36wl2SKP3Nddw8OYPmW40vLs5C7aI7yxoUw
la6SjkA5B0qA1XmbJ7pLsx81XR8MMGzUmbRQYiPQBTQt24MkFCfYojfh8Umf3xDT
RJWU8WYiLb6MBwDqsN5itLLrz8Z53hWfKdpT0tbPLxEpXZ4xl4hXn++y/Tk3xAG8
OtHTW9Azj/pDYm/td4dvxyNnDTPkDMnWicSYDSFeksLzPsNreCVL477HiVqXGPvi
GeDMdKN2Raf2bC+VxaWXz0fKkKaPrKRn0T02q4s57GGvfhBBNfIXt8dJZIZno3WI
cSoK0AaNDedFutcgL9qBcsFh0UvuY7d2Zoj0pQunlGEtZFBIMLmNEo63ILdAh+kl
faqdjyxEx7NsXcxfwOfWJ91NccJFYsq4Hg5sl7Ju8XWOT2uk3XchKHZ6aUMHYU5M
Zt9fgnwYJJPzIKES1v6x1alPcwydzFeUAHdbDS9wq6pdgwFVX/fWR0SEoyjDlltu
9BPDLI9QzWvytwLGHUv74wKHCosMh4ms8RyjEGboCSJD991kfYwNJAJPeb6Z2wm0
oECUqHuFG61PjpYWoTRHkeH2i/9clpXsCq6XZx1vHrCepfHHC0i++yP9IRuD3dxu
hP1fIFjedajgxhdC6xfQC+fg6b19gXBJiSeGwLfdA5ICFRXrhXrY0B1TZMvWzHl8
C4WbFgNiLLpsLv1wBTiZKP09nqHl9NOUTm/z9zHxv8c2L1zBgGCMySODdk/tkm85
0mJIx2TjAcvfJkqC6ogrB4E67gvadpxk1dsBlDYVwoO22zjLuoGg08kjS8CQmoL+
BMvnJKOkxrOv/3ML8GlFHLWMoMdbNpNieWCergadN76IVfxOEwQho6qW/YK79ZZS
6NX2qrvOq4i/hHp0nYDsO8zOnZUnKHp2GfhCIAXgMp4xXsW1qIuQ0RMLBQEFuxBh
lf30LrF0eGf5omR5BY62aWdSrrStY0/XCvRCs7gvObliToNjlSHQKXk4EVeJoPDl
Jn6Epb2cO4FFphGB5VdkR0Q0R2K7qrWcnoMLWxmSyuMsjNQEDymwLV4S466FgUlw
+mAwCp8Kkx7NKnQ19NTfcACCF6xIo9bcrkKZNzDvMau7rmz6bjsDigia0S+ECSi7
0AvP2Pv8B0XZ2v3TA4dSWUsXo+64yyE+UkMUf62J5YzIvRIGTu/D2UD5DiJv3MdI
Y5oxKMVQth/lOF0q8VJzGgrNRws0IwxHeS8vcPY0rho4i5XYnEV5j1lEJvl0VgDw
WKx4AWKRKdExE/m0HLWXlO2xM7Dr7sQUJ9tUb8OUtp+gFuZ+qlIuDjrT8J5OJ/ZJ
rxn/V+7NMHCHWH9sbItapgkkkId9IggiX5TzThMndD8dC8ThgA/Ueh9iljQpyslq
IH+j29KIyf/5W2n4zXCAIIhe+FpQOKdXs7Wtooo0+hEnSbQ1S1fUoPkDNLKalkch
3Z+SRgVa9mVXOx9lMtXeg57d08zEsJMKUVHUhJgQQRIYVDPlZLl435etKx/Uv4DR
rHKX10VUsbLf3+AOIs7rC579PBGnBjCj+8MMaL2qQ6ThXtz10wjONhng7HwbYZGL
ixD1xjIKhTCqMR8WDDMM24EbUfMQfyMUJAbaB/py/pr2cxpvbClwAuOKgvckx8+u
KB0qx5P9BKpusJioEbNUIRKLmQ5QsGGUaq0t6PaPGckJq3BPZ2kab0kPGdp9J7gU
kbGMPWW8p5VHFv9/29jAi0EF2D5E+mfWD6Lkgv2pXzrC+R9KxZt4XbFn0MB6rOuO
NYkfmCTOb0Dc11RwLhVy2Ddh5ZZjhXUZzaQvvlCXc6FSPXND6zCv4SV9HRCPIkG8
yJd+xDa/WCfWQWJyCwnQzr26okuFhAjlbx5fOfvpoSGo74kAH5kEynF3fZHy5u1r
sZInilGRvYeOc97n0ObaRYmVROxWbpmvZMVUn4yZ5pEDg4g98yFAVbRZ2QpJc/go
KG9gMkLvzVCRb41h6qKCHVM3wSAGgCx9AIkExOqMLcnQ96LyVpXcnNspxxEO+Xmz
j3l7o2ChlIGi/UeHZ6lvlg/PVb0hKL/dwxnMcuuvxx9D1XkhPB4xgz0yPYWL3Xwe
wpBfbWdjmw8Y1ZqCYNpcnmdZxCI0OHHUKSgpcCnP2CXl0gdaebYWGtAS5gYS8Zwx
2Z+25D1lZqrhQwdBXPB5vQUWwjt7e0E2OjbBBxdI4DFHpu6FZGrApYBZkYqar402
xOcaBfv/X7/AFNTNyNzfuM3dp5DeCV4JYcF7jagVKO35nS9Df9XokHSx/uQXaQwE
USnXgfMk2I0BcZzRySDCgAUF3/p0enX5mDxwVAI5wr+kk94mjSKmJlffllQ5MXZ2
bB/mwbb7EA+Bpj/0BiJfVsFb+m/uO5wcbA8pBu8zLGrMkJalxDQVrl/WGImU3j82
dMXo+ty/v1t3SIGNMq3t5ao/+yAdeMejszNLCyNmXlIuk9g7elJoVHyTwoe2SoRT
vjI6+unlOCLHlsPGih7JoPxSIxELz/d1q1qvS06dJE+S2aus9uBrh66nfoxlNHWZ
3iPp1a66xVqFewOoPXUt3YUvjwbB6WEEtJOOH3nXkESspJkojIp08JGkKTO/bOon
HbcAmjajsFYFo7FRHm1tnSHWfmsADRBIzLREYTew94Mdh9ADCfYwnVKeHu02UPZg
6At6kF3xbAWR2/dNSGs2wWJxEu6K0nyMSQdxIOL8LFfevsxnTidEFfdNBh8qGO3Q
FqEf1VJROSSbBpBmfS1c6xfyLhgl+Ycob4/iPIXiELBO1USlwIVzVJo3vNPpn3En
bCf6p8dVfRijEwDuqazJLlbj3/N6CTIgjOOmTCtoFX8czJhbU60Y9rIBI6QbnWPZ
RFjT4VGCLO3whua65xcU86zi+s6nFFV//vEe1ahsFusOlh2XaW6ZGQerLtoKRgMq
Qk88JqyhwD5u2tcD7+P73ehR0Q/kmRpfz2gebCq439xTMbPMJ1f4MnTEY3gKwhWc
i/ekiZpNswl63zbhUhLPjLN4AkzEexC9xfe7r21Ye/44avaUWTlBBfNdsAJAWmGl
8qcOntQwZJQIIxXFdM8cnxQwtkIH3Ms0rhCzuHofJJePgkQBtrxF3v+uy/QShlRC
q389cxeSoPrj7KOpMTRYsftmtwEwgpGq91rHBuEq1GNUrF8U/nM6ctV6jp5CEg1R
/DMMvbq0BsG7ctnoO3OA1TBZjkB1Dq+wScHUlI8XaEEI4a1u4nyYZ08skfAppkc8
lvmilG5noBI5nLDjyCIrF7/uq2bYlmKjdPukKKw99ctcbNp1xor573HhKtdLfciD
Q8XFRfKgGwDR1+6Qo8TbG+t/NuWYd481P3D4OiWzk8aWfiHNQ0uHoXoI6MuPxJjT
HZX+zKPZ3ssBdK7XRG0Cam+fYHjzAHkZW2BDsiCrOPmN9rzjh2pOAuSK81RZAa97
6dzBxJSRyxR1htTsUbc0I2nPtCf/DhjwgqiNB8BoBoK2kIPFUPABFO8zgfT0zdBT
QImGsFOBZwoiD4qZlKboUf9Xgzfn4dH3EKIsBBqzxZNSsgm+ir0Raxt6bK6WbWKV
G4G4o89ICG9DLzwiDF8j5xIsmEKikIuqmOxlpnOK8vQsEYlbLhTmob9IGhNxxb2r
M0fUHv6yCfunb/M/elUEdN48la/wD2ca2UCPK6Rlzg5bye2PP+JTkCBZLlXObisE
90uhU1EiDMsKbQ8xxDLEYBylotMYb/lMXLhEXup2ZO4O8RUh7ZQYlkwpzTPVeyUK
malkYBu5JP74KYPm+LPIfYoj9Nn/Na919xUb3PWrpNMdQWaM+852eEBG1qVi5fjX
U1rwxQPlHngjMkWPGCcEEzy/yjNcOUet7d0uOn/jtTL7TDzwkmfssfd7LBFTLBXH
lPyeu24474Kh1f7AWl4Z0cEkGQ8Bk4s1B/9uG+Pd21NUpv3ngB3cKn3yvsc6U8Xl
3lDko6K3xPEnAZOwWxz7WeafG60KUBLWf612j1N0zSvpM/HR0MU/eilVwcKft5Uc
NglKak1QL6pn8FtEm2zs8mx7t2HFZEeye0r6e9+djLyXSUPgW6HmRZg5aR1zKhcN
N5JjTfaTKkSL1W5dQZtxRwYMq7n7DVnEOFkHF5kFwfwmMkTOuaZATcQn++ZPueRS
oGy3cdZ6dtrsZSwMP0L5S0n/mmgMTqlvAvM20UJRw3Z/drLBlA70yP+ppbqCOTlf
ymg/k2/wUMtmU3tFW2JDnppKK59V5nrmSiBw24aQf72ogaow0PgOziU6jyH7Z2Me
dXbDL5qxE+/uu4z4oBSyFVQD4OpHNlfM8hZbmldc6EUS51f/YLJpjNBuXIOgVMqI
uDaVi8YH1hPmludBbv21XTjxD+ADciqD5QnbpdZ+Z1QvbJnQ8eaL/gpWNH6iZ36o
eaZHgdRN9VR1RCRmPpJhGzo/p4Jq3mgFNt3/AlyzYGJaWl1+pfErU6HeLr8aSWsz
Xl7NCESpEiS5b/pYLpVBDaaskmVN1xVYTiq+3QzVFNX/4y4rz+0oETHs+qFfNEWO
rTJn/nebBizV4GlmTEd+o3rri5+DDoT5lEIos4Bf9fV+J/znMtvLwZMquJVRODeG
bcRL5U9bc1ZZENVS/K8QfujsaSFkpejQOEcY3bCMYfGH4qFAyfk3NmVER63GoFMO
Os9BA+BP7PByWLGq+F26lyhv/MrqJTJKyeAmsJ5qqJl98mrdyBF/7fa/thBUGA4h
0XlzhcIOgf9D9wnZq4oDgRZ3ZnSJdayhtFy82kdVw1sYSy/hJhJWocmW85ZB86Y3
BfP1BWjWwSZHTxxndffWELvWEiyNDBK9/x9sO2QG7Ryv1NkqwzkB6DxSmodrlU03
FTyXSAoGRCKoM75xP5N7sxjglomZzGp2vHzGLp5DBBekctjHFP4nG6cmHoGCLgX/
iO1hhrm5vJxu6993cUPoRTSSv6FPXmnA12fY9am/GFTL7hG/PQOSE+rIGwmqJncn
CAuPRIxhWynKxzSmLR6vxKznaYz0pi1A/u7aZR3x4TgBWsut9zS20sYsSzeLy+JP
oD7GHfDwiWpYYyO6/jKT3y3zmg/VJuBBD1fGiex2UAJup9EKHWrmjNjHE3yZ9Q6s
SSAZCb0nO7or6qJrH4cLCz6rbsEtt+4ehSZnuFGwuFdDOsJbaAZ9+lw2ScUaO26B
i7ugCzmBP2CNoPXbdWDEjiz/dlkq8OIGYvIeaKgIoLCdRJiCu+D5Xo0vZn4ChY95
DKr7hrHygSI7Ate5kpsplYFBTjmJagcBWxj9axNwIuzErZJA7narJ/dLKBI1YzZF
5oH1K3ILFpiu8i+e3eXUWXpOPvo5SlrZX3EGDYMTet1UcGe9+VnkNlQsRXqcjx94
Cb2r0FhO0XHxr5blFfLQoCGcV4wFl/7E7K+eE/12tcoUt0fT+GnHnbDFcIy1hJ+e
oId71wu4OH/64O6zeHzvJfQOEdNNZJoUU7glIG1HvpKRy/b1Dhvm5rX7s/B+UczM
IWq2//w4t3rktP0l4PauM4hFWa9oosJ2v+HveEMuGsUIlfdZdwTvrWRjvFLeQjO4
llQEMZHlMCCvDHAcFLUqbabOsCrONd5mjik3yN6a6KBPRplSxyk5Mxw6yP0a1Fd5
TG60uDmKSZoX/oeQAPO1aNzNB7+KgmOC/RXNlf96dxLmWI41zyS8jEjYkbiYdLIS
8DX6hfmVa7zPZU/z1YtpXKEL3KaVqwQ0tbAdVV46u5iXgr272P0F0673XSz4EsRC
Crgn7gcXRI4Da8HFVE6UkWMcG1MZLlaYljUWS87aszFynC1oL9Je1avAuBpCMysI
b+dIIDOGGcHct1rrKCPrkwKJD/n/uM1nA5Jo4VXXOwKyTwYIA39XUxEeVwAb5+9q
NimtHJ2+amBAmeVmSqV5klA4XaXJZNuggZQABpfp9nwf2eg8uxTOlYj/mnmNB9Fn
2Q7/vJk/tfkFtYhgBQJiBcucejXPbiXRu7U9GGAsmN31WorAWeyORCOHROLxpKbC
ysNo+HdIhTa9v1oLU6k0DX/MUUTBXt4hKOFds9gSt8panK9kzE7/hM0b3J9JXKi7
DzY0Tu1G1VwFAgzJApqyt4JKkk81h05F3JjopflTPqZUE5EwxcANwo5TANg7OC/q
hmPOWIDQTI7sDzKQhn2r/82uuPnFa3HHEgiazdsnPsaVf6zGnSDWUvtMxkemWhfs
hT8kqbKGQAgZItlNem3O5ML+OC/U3AsP21Ozr5ezS+/IHezipW4maIAAU3lstHQt
SU5fYcWJ2rpmXaxWGJQxgNRi2SCnADu6QqLywzA3S+JtkReusHXpqDlJiHtyhRf0
OHyLPeF4wA9EyOpbGtLua7lIW+2Z8pRj4uqnUfC4a0mMz8tpxJS55BOFFhZU902b
8yb6H8PpfwAaS5dg+C8IU/u+efyvcNFAByvdRkiEe1/ox4li+xsrbRReIEc+OVvd
zyjraBKcJ6Xdj6pnYRrpBh/WikynUFiVXoHR5sKaZP0mKAXlBs99//6zOVcWYmhQ
YGNbYmP8+IILhjD4GnJPe2MQ9gRywSxR0yLsNsE8318MvHxtUXIgloCQPOSOXb4Z
ahJzp+BFjSCbsgj9P0ZZit0a4VqgQuUCPSbfqITB2mLx4WyEhZKZdkGDkAdvVSXo
4ZCDrCGpDSNRUPJWx126Ip1pgsUwzcxrVEZFkk9iJj8LCg/ECBmfTMgUyOBxc+ii
SmI4swhQsWeffxO4ogYTqnAEWj1NAEJRbFthkD5KquYivsIAt/stbyK+hOBNTqfo
wUf9IdqxTI6oY3ty2hzJ4hhgkxbSioPkDFNAj353CK1M65pWiGJaBxvu/UmiMDgK
eorB2zRVyGq4fYciokSXHxew41jlMavFK5S3LWJAbec3P28m4YxAfxX/gN5kyBTF
QtjlOdE9yS0H3eMb1CaMntMh8M1XOVmZhPVEoiKaTj1ONPGlUZsD6ssCatkRK2UV
sLI7aXd1FMUzsLuv9CeH1s/GslxRxWDAPxGuvntyZKuArjxS0zYNIgcaNkazZkhn
0MKOPGgKSj48nZgRJxNlNMh+gux7GBjijp1s0vWt2L+AgX5BNGZLHDSmMrsAOd8N
PGGVhA2Y4vygYfB7BISSs9kapAQp0jaZo8U6bjr4G/u6Sz4nuDpFJXqY4xfTiYAm
DbJlxmcpE2Ua7f1R2iE5jM33K2Nd3kgbOk6qKJ0C8OIxRwwZT7k6C4oJGfl2Ify1
Ve1xqR0QYR7/UPuV0OCVfhsNHezea+BD8etIaywA3x4ty0DNibIISPgV4u9LZ3kf
rApY9fYJUQ3guBxnX9XxVZYjOjpMcsDvmA8tlCFhVJaAQKu54qR0bH6cS3x+87Bq
7KUuJyCQr5MZws6cPgVwUSBz+zHEzRaQjRdrdbhsVyxhlAASuW96tq9PrfHUlet3
pmsFJ0Vveu4lvg+aqzuyNHE0UdWeb4pQJpu0qogIrUwVKnkInyQNcHX85FbIiwgt
Q67XjJjAdZg2c4/18tGCBELxNEeFwfoOL8pxFLRfitklPdfYhbUDG8ecnyVyQNUx
zKGxCVd0RaCYMYhOJWkwlPPv045fCmsWidZ/CCIfbG/VRV7XToiY51E9QlaMok0z
J4vNh8QzlNcpoTMXrZtm70LjU/PHzRZK8c54mV4QbQezdc9+0I5Or2HnL7HurTmh
OWixUX14yp5wEqrOknUXmhpAaO37CDEsykVLTWW/fgi0cUpwKfxK3AZz2Vl4KHjT
yAY+0SIQ2ADQJbWoWikneOLt1lE1GoB3xDFy7ELhGm58lX97d1Y669Ihulx9QW8T
+Kxpnt9X9j4AxsPkGw7yKv01FufAu0yzO+2NVqkQmLnSBH+OkXvHsw4AAvLxPqqG
WUe7pHIotVHSwSPWKUxAA/g681rEhUplPT0JSDG6vMaUYcewEqT8RqzYdiQoB0Ub
2zKAEjq0xQli9RugWXXLmfLm/obgQqE4HiOnjHSOsSe12U6bs/7xMtQRUpSZHRKr
eGos4Cn2y3pN7d+d26NHKMXokCvENa9W8OKhmMgi2K/vDeYxUUZABs/s/PrUN9Qi
AB7ltv48MhgBko6mk3zeP5cm0Uduu+H0EQoWt8eey1w8IqR1rn9eU4qhsXuK0iiL
AOiS7IcBdBEaKsruie/rMri81HUmuG2qNHDWm2aKTJ0pT9m7x0E73X4Y+Dky2bA9
t/RNSNu0a5MDPj4nYL6JhYlddzzXhPh2HmbVJ2MCv7lC8+hHjjcyKJbNjTMSLN6C
3WIgg86RY+ZTRpYHJjUdoWWkMVRUM/L9CAm8lLnUdslOxvqMW8Wqn6SdR8QvJWk1
32znWFS8UR7OT0h9spuev20m6XFRQeZZ0QmSZ3dBM8OUaaEsOaWTn2e7kZo7BWxZ
qjmb4J8UbEdnXQxaeOae0irOyNR+5v1H9pdRKSep+9/wq9ulQzrCFwSZs2MC7Utx
7+k65oMw414mG8CZMIQGDcfg1MGGBMeeJng0qPPYM3mTz3PM4XKO1U/AwaHmi21j
FN0eMzFYHo9564acqHXlI6ZCo6Jq7egSDt7rAu0I6tdQvDXHvDXYzAPqUdKS0+Rr
W1QI2vVOAd6dKNWISrqk/kj0Z0vCJH4EbLk7o273n8htHbE5AkgYz2YUy2aNvJwC
/LKBg+S5cWv4ZKVkq+FV+6krbz1BhRp3i46Z0Cb9ymqR5rfTXBuqPOIyVLeBAm97
yLN3wh9bTBhlZ0h60W1/1dq1yJ0B4hccn77zQBeW1tvOeZUk+jYP5UEJEsDe8XgV
zFAoNVnMAwe/055wOSHBeEpDaNOoXxXVHy6p1feQh5vRz/YMwFif3nb9bWWs+Glk
KM+dA53jyHX4NQ+xxfqGLYp53vQrDMrqeiRU5BuynNdHl4gLeYK0P2ynJ24A1hTL
6bfx23Ts9Pdb6GWWKjSfxSOc/S3UGYziJQa4/S7mfqZ1AeWvmT1fvOFJKuR//YLt
Y/Oqr5+zRI8I5yPTwkwm1Q2omIMAPO8thTWx3/TB0bISmLKTiJ5QW1U8EOCF6eU4
xi0FjJnoc+TDIjNMpIz3oGrpQGSN1VzoPJXjm8ml5rnqEeZfVabf5UdxdlP2/J6I
xF4WgU08C3kAC+wg8Hr+OmFkDpTBBtT0ycOGa+24lTqAtysxyLSLpLqt0oQeRjpQ
PolbsGtaa3z4G5+26K0oCsBh/9T7hoEk7U4VhxIcmbsX0P0DPfcP75M7qk2+MUNq
YqWgDtBMQ7kyuAEYC7tGSeUjxSdJ8PgtjUWxyfIqUZvVJUAlFl0HRwpE0hJALwzj
KJ3DaVDj8jVEbeFYQhdUahz/vWtss6dSmKK81EjF3xObZt08Gn2zB0v0NkP453QM
68316U+1KwmgnPc9u+ozvE6BGDccPZ6JyXEfw4Bigxjz6mBS5ZXvYt69eJStJWSM
qZp2R3IRRnxpQAxw5oUBe4TAEADDYjJomRPCiTBdFi1TcBxE3rXVr3ozcuD1bTgZ
fGaXW2l9/u+t7I8o+L2GiUsiVUty24lzq/ZzACG33uXge6SesJxdM2VCIFJ0etBi
aFu6Sgfc3/3qYTKrfMy6YLYged5ERSr6zARCe1/y7/Ixe6dpMlf/Q3PqnVUbeWbZ
44XAwWdSc+sIXfrp3gCjOjVcH1DeM6Prt5hGqziaxdsubKTDyx8iCJV1O0UgPu2C
MJzpP4CoOgkiTANoP+Fz1ldu+84WRicXFEgyyXG5FNzfuWzWmmfSwzYffApHBjlL
+Qn8BfTe7p0BoW/j6pDiB3QUY9zz35VJZsXHDEF1BfXKarU4FqWZB6o1+1rqyMKf
ALUtsK6BdT5XuDwNMpAjFBgyryzoOYCpIu66YdrB/KFw30DqpRuMntIOWX+a3zgS
NI6y/dmP/fc7NesilMYSNClDV3L96M+sZEL12rtZWtIRSwQ1+/1P6nWB+Er+3iGO
kg+9aPjbQxlniwPVm07GogZBZTcqLpCu5q5j/uNNNet1xITGsdwo/jeDm8+xhNq9
KcEeGeBH3KnKpioOpM5cIBJrv4Iyad37dhV1WHsjzK3X9tFe34B5d+LAqNg8Q36A
lFSpIR8bMttkpc5orKXwzG67WebN2TxiV20nRA4sV7ZoPL3R4ywqN7ys+JrbeNMD
bzn425xlbb+T9SzYyq0/M6abmD4seCpvtM4gCCpWgfUCP4G+0XtpXnbflN/NhKGZ
/aw5g32R2X5Y9zgD8AzGYwqnunkFEmhWoUlubZDPrzvgrizR6MDssQoTQTlnhIbF
CwHpCKT18SeQUTFfOsW0Ldn85tUErnaUa+3Ug2JZyjRKesRe3DyCBCoD7+mb481x
Ql1dw75Of+OEtM4G7AyzugSUbi8juR5VYrGy2rEkjh2JVx1wHzpIZY0kyhGMTVCH
68j9lE0EyM7j1AeM9wHOS3cdvRvYbGOkm0x6uTvmmffjR/Bkfcfcev9zQ4RPYW1t
hPY6W6K/FF05HMKR4h2jb6Ew0WYn1hmSgMLzsRRS39/aS1f4waHwjdePyaYpXDfr
lO6F4qsGO+h2E3m6pok7Oh9sMuq5hPiYqduQb6BPHW4Dv/BpA1Tpi2U9dYTOzGG4
3nS8PT2GJ4ZPMjobeJoDAnaabdjksl6odSuHgJC8QAAHmX7IQiDp3NP2hek9MMyG
v3t+gQFrsACF1LgRXYWvDGJOOduHYlgy1zHQjlV3d2uOHYlcDjXxEIY98Rx+vVbs
z2ce52bPjfGy/A6SmH7UqjroyYZtDfI4m41emO9V3gbfpWZ2OpSIjbuv4G6nzxN/
Vj/NrTmPCOiSTYK9mQBf45Y+pGqEcXtstPBNlVedm+91kzJb7JMMXCCMFp9TQqC9
pWWWFQ8aIf+6h+lFPxInZ9998WXOklzK3QNiK8d1impcGvVdehhyKRjFjf3WL9lZ
ozKkaeJrOQiHFSr/chQGAgPSw3Qw3oPB2aOUaeiUrMXw7XcokhpKRKFHniz4AOYh
2pXi/Lkfg9XQczue4BH7kE8MiNHavsdJA2ssuwJ3DJlRzScw9dHKcYJM6dGtLJBC
RUh8/mKVnro3PD4viicTOCHIN2TlH2tTJzjRrwYFkNE7eRE6BAWF1rhm6OQKbhce
4QnPQS5BUdTa+SJTNZGY0wGtq4J7v1cy++q2I6M3MdvGR8LdhXyk1EY5tbCtOZVn
Dwf5rGlUJutUDF+FzrFRyXCsoPp6tS8tRx+4pYDusg5rnavWlDnDJsAVNGhMwtLd
NB8M1gSqWK8C00vJ6zVRZ8I1HvyOK/ryD8fly9gUyqOFpNQKFNyWaiFFNy5bcK/E
85xItgP/GIwsvnwlOumzZ0d1OcGPesPxeNhDAspCwftA3lNuKNRJ3hni23P4rzc+
krgx0Nto3z00WgbAHwYTXu8t1JCjzGoYoBd/QrhnLQ2oixuvKHSCZVGYi4AdPjd5
u5qHzOPW1gbHycEwa81JfOqk5nYi9qKmzAaQCzc0eLTLwRJ7ouRJe2ZOwsyXmP/6
n3iFrsosd3KhJqzwtIQDWBBExvw9NYaO5PrZAFrbMtXUWSYw/WFhLP25c6j2fhxo
cwb+clv0rI6/DJGn9duwMATUUhV59bAROzVwWnX1kSWAd3C9gNmghW65W03WXvkU
qCmchYmLjhwNSxgleVLTYmUvS1nq0c9rgwMvLq5CLbPCDsJ4gr0vfFBTGHm7ivyF
K/cXZKm6GFbRqgQRLr3TIfWX1Kau/pjXfZNb0pXHKvNvELL6dAuCFsZ3GR29BAVu
JhWDFOmGXOnOYtmy7c9yIf4ZspU5A9D7u/SThK0YXjm+XTa8cZHLlvR/MXum8M+A
cNzZjiwajnxzsRzgV5HxPA3Li2jN8E4MHS47yNMx5NzYD4u0TZwjkyE57Iae7jdD
b5hs7QLDB5t98BMunnY7YGZ7bSyQc0FmQ/EqD8O1mz1IgE+tkGjlo//n+qMqfaK9
POnDz7b24XPZPTeFwE+5xyVVpgrdVBEUbblgfZ5gxjK4cTrFyTUkp9cLnSguQK6a
fTJ4+mp6ZrCEnMG7GbcSeVUFFVs9JCZwIKHMhrPTfKsC9gaAa8xvHWHVJ3YQvwiq
pfSxCJERJKATDY/W8Pa3pF7ns0mThN4WvwBRNY7QYO2w4EaDnvznhPztgNWb5/Pp
m8H7wp1Rh02wTM+LCEjr9YYK3WAoQM1Sjv9PUvRimu03XsbFaEMG8f2iyza4lM/Y
m50wvgEok5LiQb+fygLbq4sp8brOn6pCN0tmBF7KApjeumSWcbC12ER3VgK7PJf0
JLdEHBf+5DB2m17i9X/JxfE9Ez3Dv6zIC+Y8I6ld7grX6zFIcdrxUxwVgsrAbifD
jSw9Pc0kXW7MFShw78Ajsp7HosPkMeftpr7uC/N/byIeYLAnjzSG/6E/10wym9DQ
BfEtLDbl+gnIw89UzMoyR8TBDRfLREmqk3xLKivdZOuqUoKI7mn+gblYWpJ9rT5b
5tnn3n+aSIyw+mHj4f3qFV7tdvbX/GK499Td1AbvWpxasguX8H/uTNgy3vzHVNG3
6BggDsRQnNzqboSBh9WuUY3kqWXTtOLIiPSapKsICDRupy6Jyw12p3xX955+0bBp
OCibnEQoq05HK/tyfQEn/qBn0+5Gc7M8OSH/uUUsDAwsRz6fh9hkv4ntLILI01dw
6pv+1Pbgxo7dN6JWiJZ5k5I8ZrPVS/7yuGOzJGWEVde6g9w44vJ7DwbOJx/jVnVv
QDwsq2+QjBU50qnpTDA8liW3m00n8f8gwrrB0u8PluY6mmHFBV1EtaFWhqwthz3q
ptfusqpRAvN3LxN4xgeUlLb2tojGmtiSijhRrCWFwv/HS8+FzGBGeFeNPhJEWj7t
tGzHLB9qSkWvBk+y4Y2q6HGaPg/9tBzoSPQWsGmDCcq07VgFFQ7tWfGfXB+/G4Ge
2B6AYwCBZFVnG+qs3KcB5bI2qED76Jm7Np7aoVh/z+I1z+gaXU7OETmzTdMZz4pT
toLsZhb35wX8bJABjcHNkN+U0HHl7OQ66eguNGWcVegTnwkUfN2AC8A8mt2T9KGs
w+NhturMPqWGynfYr0F6yJhtio4kfXwA0yBXTQIxVPOfC3BmzT6SVHp4ssBf0D8B
djOyPpj+QUm7jnpnlRnr5u6rgC1ZSx9hMlKf11bgi6y8N9Mlk6wNxjJ5+X8Tc2ts
hJKYOZxmQvHMVqumXdAv8Sxu/1uoserliuhUlQZz4b+LbdbkiKTwQaV2FiGHt041
Q2S+fhWjxXjak+fmI2fDiL31ODAjcO9xOZXClefD4CpgftWSd+gGNcY5CTsobD4X
K3Iid+jCdU4ARPTQsPQNvCCXJIDI376yXuUvAXSskbn6rZuRGA8PPvvz9CnEvbS1
dy0OPGynd2K+JkNeM+aqVPqDmAVavrLL0S0Aj6KfUR/nOyNo8SVGS1HBngaOWbVl
EF+hPgzWLYAgOuE8T65dqHZ4olhUNq4oqrTSIWyHBKqGKO+xTHUmwSogBoA0+OkT
unm84MllLFIUgGO0s1a/CHH2Lt1uSKl4k5breaX+t/8P6Z1xPVga5d3RFlei8F2d
4o84QGMjgrzLqHcEysslUj1L8S2px8vfB02Vz7dq7bOVFUvLPDzPkKnQRvae07Br
XhKCVaZRQmGHo9Ifno3i80gRzHUOiB84Clwx3k3mbjNs0vBs8BGmGxhuIyrpvNuS
eFe6qekiTPCJbY1orgqGlPWjufuu7SipZU9hjCRDMmqZfL7nwS+3SCdwFrWIANVE
QU+VqTCJPiGsF2g5bAgGCc++wxg3xqv4AvqU/dKR148uiS4QA9isC/yoCcHNqbEb
S3Wl5YcfEmmxAsvmnjJAYZ+VTxNz54XLuqWH9CY05UJn0qu6qiJrl8OwbUTvuOsU
IkNkUmtr4Ba4Qyv17vBRD35eL9IU7U6RZIzoyR3yxwgGPssU1sXyuVx/f5LCknFP
ut7Tvjluvr0bcEweUlmMpCDABKk/Kj0c9giUcAcCxx8E8NMdsDtu5skhY49vQi/z
lRJUS+xjf8NTqSV9S0DMOeitonkA201Mjs2bDgF+lHA9GG80xB3RJ846Omj1CeOE
9WQ+ZZ7DmSICWxjY7V9B9J90xL3/zsCUK/A7WtIjUmEHDiq0gZIpO/TayhW0laJF
05i4bpzIE3TckAOKtlDlHHzC27bq1x+Tfva7JkzuUdIIJ+mdKZcSdflnoOQ3H0ub
qKIykYokSNE0OA8BHnVMNA2L2APo49lRL0ouLAI/Si153WT6PME7/RQv7gd6B+ZQ
9klO1hKW2SUfbN5x3856/4Z9zDk+6AzCHQBMepbPp6kjD8kCRaPPC2a6nIgXY2S1
E5+jR05fFGaZeTBy0ExYiWCiOy8fEj8Stht2MdvuEAlst9IyVUBYv7ZhKQpGAu/i
hrilkuGhpX9lD2AO51B+qAjyRvz8TNjMMazvxswwbQp5Izl8xLEertfQVqM+ksLA
3VOZkVy10OPqX3AWXgzFuGmxPZGuGP7rFplgV8197P/axfFxsVlxZXtxR/8J9zlU
gRL/YUaEmSsc1foccYOcC09LHcw51eUQjWfEA8APcq8YFM3BJR82/f22mD06lW+l
07f8icMonPIFdysBHZ5Iv+HIZcdBdNnY9LfMHSu17hxyVvkqFat7STtotLCng2fO
ob6Ibcxy3xEBt88Z8XN5eD2ndz0VGrYzluJiZ8UFuvaJXBY/jhhs717LZsXzS4Ti
/P+2ZOAKVW6Y5DfHqpFM4gTHrGd0ut3UOFVMK8D+nOfHMMYQzgNRmm2ttuqBaetr
MlLhn04PurX2WKa+806uKeYqRw8k/Y7/cix/nwakef7VOGrB4cZdVtV6hnnHZOWf
WAd1AxmF/3K4b3FX/LhG6w8vUxoXcmghwNHyNPTkdmi4OIgJt1HYpxgVLFqS0rhm
0COD08mONHM56u78hH7DUnNeOT/8UiKvsO24CYJP3X3bWrWPFiJznfsQCY2DrJf3
SjeqIno23jrBU7yqIiBNzd1KGc74p0qLpiB4Y4sn0ShDnWwatPAyoKX0d6XZCQ9X
T7YZ1WUZ2FflS0XhBhahzZt8AVoZJHpCp/6Rp5BzHSEDg+zPRLIXjqUt1h5Pdq16
1ERj6IXroZaymjcSDq+DXJMpx6EvVj9QnY9eTMQfpmZPCownusvKhPy1wy4SstIv
d4Q0L+xD3XPVFgrT/FZdthbSD4txpWetH3VZiRmQdoPrEOgvL1wWcrDAykjzZNoY
LappTJ+LfR/y/QVBts1qsaQmGXDpqUT/H4oi5PAgDNKXiTDnOaoHUhuOvnWHZAqC
Guu/zJO0n2SzW/Fq7Jo6XVKAsS0F4VXciOtGgW5hI0wRYPOBVGPvouwDPo8ZKt2l
FF3ZJ0vcNYUuX1TXdpSwhttskDNu9IpZjkwKafrFNRKa4zaslBRqsD93lVExlXlG
by6x0B/sI5AX9LcR7qEEMZDxOoXS2QBOp8pvKgX4gNRX2fSfe0HT/7gjPVSJ8Hcb
WQkyGaNrV2U0gg3LjmcLGFpYpsenGAxrKv+FQvZRb5W37P7lraxwsG7LOfE8wRcw
f5yjrCYPa8dj5cj80m5Cyk0qHjl4EQhK/DErce4N7JfxQCZ1b1/q/OGRx9Y526W1
6N1vNcirKRwrssub2CwAFeyj1jHrjUQCBTwErz/W34JzVKCDKwQscSnbPlyYjdgM
nJ6gqZBJXc21hvp1lq29DnsESG+wEHopDIXtBPS4WoMLYvdZJmMpFMZ2vU/iOxxr
ljAqUHI4Nq9yBtiP9crIRT1967kXPlFt/yxuFNTtDlIjHi9+9/KSuPCsdbHX3ljW
VUfQGxkwAVoowVTE92T/4DSfb4fFfaxDnH64PPTTkVjwrgCXw1PZIb2YDeXbwEcO
N2mNrKZjAJXQi0eEKaQ5hQf7EUAAfUJvOX2gBS3CqmW0eRxcEK/xGhC4y4hzAwBz
Ug60FHPRWXGdELDu+vmh/F2r4vb/LvAktiHJoq8gxmLXZvrk97ktxvdxxXSRCYE7
XwaMl0r0UqLeruTCMq09Xnyy7vUwsBK0dTeCzhv51HzJE4iy2HxQGTySE8mixanb
anjsOrDIgopX3FzsratqAqEimdnIOdyKmPiuzfzBaJzqN4D3+VOQOhXC2VJCczzn
yJIdBCh4JBxBFiDcc5kgr+a9kE3AIR6hCHo9zA8bc7xEVR7AEM8aa/nMSUitMfKc
m6AyGTdnokIBs5iIXBAwlx5gdJ4An2Gk88VUu92JSFIcxeVHFfvK56FHlmfYai9i
NaKQo4XttgpinDEjtx/cINOx5J07USHInyBurVYWj1U1g1KNq67UpS/HB0I5OWEV
iKnQjKSzHMTGX6x7PXd8hS4A5LhkVKrY+gmbVbbHrpJyPjBC2akPC6gY3O13laPc
Gw0sIB306dA+Q7/bl4jiuHcD9EKwt/rreH3c8RS+eO4Ai4Vsi05bd9OIHh3tk+OS
KofeB/wRO1FvT5vINLveuutVDzzD3ivIDW3spl6iK3OILQwDR1cb3qiKxWxPw4fU
8WaQOmwBDTIakS7nHugn6Ju1vJB41WREhHfSSO/cBRmLs1rnnD9J/TcWNkK23cn1
gzmq5A2oNfydrXQsEGRI1nvRNy5lCm/Lbw1aPTer00T6w2Ldg/rwZMa3hTrePFo1
lj3GbaoLPqFZf8WqFZtd8Fgb2Tc4Vzsv9H7cZdmD89hwatR2PWDVPlMKfJA4nYI3
Lcxs9a4HtH3HbtFKXd6uq1pC9XxRu1lYt1QbftTkIagT5tdbsInpWPDgC2y6WfZJ
QqUrPd1bWEhS/5u4Mo+I4vuvwin7JkXp9QE/nSwzbnfsq+NVAGQc/1/Kmc5keT8Y
F0agtMU0ldZo+mMIDq2fly3FMjURP9Hwl0hex4lnbd2Tc93jtxUh7uueBKjeeM5e
zZ+MiTj34LqSw0taKshdGeplJwsIgTA0MsNhk0HKvN7K6R3HeMM10MZHwG3+YCvp
4DVe0GL930myRRyvm+VMZrh4E317YPxChRoNXBF7yT0Um6CK6+Oe/GOaCAADrrfu
ICXfYaN+elsCGWrzYuPS0Rhce4h3ze8wgpnDlCuSfRt6MQrtYkuQGD4c0Bn8Q+wG
mc04E6ixrkRerSrF18lCQXwPejRw5zGShKRVzZ+pvaocBHrLBrm0O3xOiymIf/F2
AAL51PBy6uDEUA0zUDnEnJwdZoNmVFiV1BN7sOKFGou9Wminf6I9GOwLOQjbqq4a
iwvTVwEyyjayF10Wv5nAzZqIcFglYrAfWzZMe5Y7w4j3MuMZaP+4Gni78SaO/Il5
m69cE7gtemgYH4QEwQWL6oDlvjIDRN8zDrFiWZVQyLNnQfl0LvuM6sTP7IT5Dr5M
sw/T6h4aEmJMJYSnVuvo9x6bit29qQjTyMh1EaqRtxla46k2Xl9I+Rdh1uizL7L7
ojIH5FIoS4m8yPrVSGqQHLUbYRQJFRpbFA6xu1w9Ik7podU3JXWM8ssPkH/ayzaD
UTt7rvSTlPyCt0fhAfqaYNINuj6lBrTZgAJFDcaxb2H/spcW1VOGFOaPZAZ2Dxlo
ezeBSHliR+Fi5sJS5APmwH3YYaiD36/bXyFjQfScmO3f5DsKqx/H2bSvuD6Un9x2
xhvYXwpfZz17nyErmkzUn1/7tm7pe5em1Gr6sKDP/jLsTW3AsBznaKhkTuZZrRUH
CFZyrmOPea/QU4nTXqx9ou/HTsFatYfetfVULXpkOZxotJKKOFNQ9M7FjQ8YDGvU
I4ChpSB+Xx+Qk6y+yOmmMjm1+FbM83SaAqlBLhT+YaGQDvdHsJ2fe1WUf6/P8Y8d
NlhR4PsZlHXWWqxYIhdh1oxjuQS2MJLI+42vP9Fmj+F/wYqODc5xXu2/JdvLNBLY
8S7cQhqZ++2PKX9k3YGx4UqoPsZ+txl/v35SaUY0XiiH7BIB1P4fai1H6q4Qndau
Q5f52iSy5WkgYoYmEXXN35rrJr1R3JDaFJ209oUvrxoLukojQR68YqxbEsYfpwgk
CQTPI330A3QzQeZ7ocYGZQWzNFEL2eALQ6MINsI/HWBOcFCbeGipo1c4Vj3/00Ha
fqclvZsysMRQVv/9RyG7Uurh9/q6+bIalizDCPqxgm47iXuAdgoEQYHUgcJl0MwR
PJoZTjjTIDh6FlyBeoYns/sykpUG7/cJ8uuta8wyClvm80FrijmYu0smiOZ9CUDb
QPLw1CUuVUlxpMKTQAU83R2CuEnJ97JD9ZaHhhVXWDOcCmFP/ec9pN4ZgV/KzCIc
lnrUDiS+TqkzElaM/7Qbr13i4wOCrtK1ZIY59i/o8qPx3ehoaIGZv71qz4w+1EVk
IGgEvpyfFGNbzL4YSFUw5An+6Z5JU3bpudImHHtPNvKofMAUs9M9B5wTgWM6FJVM
lCGjSPmG/SUFI4D9VCcn1wk7twppaI7505zdN97du6rSgd+BS5dUcyNfmTRdKGHc
FHtwhmldfp34urXBv3NoMlBpPMh8KzpGr1Y7pqVTv06+n9v3K5FBzamjgph9TsIZ
iVXpoOtn0nsJt8KIYwAUQM5Fb01fVPPDRytHMvnQoNsvSv5w+bVMCu6IMsDxlxTE
P8NfTze35jfLXj/x3J84O0Oru59uvA+m9Dh0b/OeR3L4rMmefGucCFpG9i8+CrT3
C+/CyNKq4vGOKD8vT2xMncsfvzmV5u/vHxtPtuBNJh+3H6OiKGGbQhJcZ4J9w0UJ
Thqvo3dRuigEDK8ocpdpSePoL5LFEKewf87SqX9K/V2FWcB9hiU8T6t3caUN7SHE
zPDfIpwPhp3yc7/5H67DjGocTD5Nja4Eg34tWbdA4Ufgq1neH8ALgbSQB0ez3Mcg
giPq7fXjP1ScTfVLtItMCZBycmeYl/dotLvdOXrFXmVmego7XoVGz7R+nbgRQngF
PUcBjq9j56MAXDvXZWkUatQv9lJUeiF4N7Yro2o92hl5qs7b1ikz3DsmVg3TlsXg
lCDibDnw5DPda0Vs9nqNEmO+QlEcuwe+GdoBUZjd6ue0ZHI8/dcOYV496mqohyzj
7Xl4UbPLmFgjpJ49pmF4RGdEpFur49Ylv326MK79hftpevNGxoM+Yv0IYEJYA680
pohsVsiGtqop6hvdtxyNNTnWNFLK1QcwB03MmBpnmPgY4eY/klb5Z8mfVZ891VCi
GAPq/K12G9oWFnwzT4Js9GWZB51tROAaCBBa5RjXeX3Sg7RO1hj0Q8VK+sxLDG74
y9infWG7xNTsIWoq8ewXjb4N7wSvoHfDic2lA3gGXAwBqKzcFsRKcYaHazYL6VbP
W/TNHjLOHnzy1wDktl44PBIAnkz+/Meqh3dQXpHdowxsxkZ8QJq0tljUA5gC/Ftd
ecWm3pMEaG07Qbr0+uPukqcONy0K93CscVFFCyqmCqJONvRYYswwBDag2WL4j3XW
ZmAO7QWfX2snhdntYHGD9tDgnDrVdX93yqekQ3qYntbkAm0SwaxMCn4cG2CDyGDS
IOD5U74S+/nCUfT7s1mRQLQm7aUUwIGXgjnSWUv7RtYVHCxj/MHQaUbJgzxNt/2X
zgj3MNNe1gy1JGEn7HDuJEF3c3IIVO+SIdzDI8IFQVdMsO5/zwUpRL0ZGDmp0tRf
kZnfX2K2aWE+WU7iymwXgzFMHWK0edi0AwkSjmX62TC8JLdjGIMlBj+5fkDSnWvI
ZHWUIqYeAxBTRcElo05rivmdp59VA5teyiQMCalSxPObojyve4V6GyM/LCGSJyjW
u9JRowM+DhZMjsx/XWIeAw8LgTew305BkDJBPtCVs4MpXbTyEwauWZ3NnWRXDKBv
XF1DeG35iVhWgSd2ZorW2i8fl4OWAFXjRsHGdb1hsVloCiF072c6Kvuf2lA46CYh
qJvrJwjS6pzG/FLFwg0ivUUTxWq/aMO0YesR6fEJV3BSBkWbEkMGwUxmcpdxOxLK
a9lX0XNwg5DEsqnDD4gMNvKnc6Z9e90k2jJY7xG4ugJTn21H8LorVd2jMWv2mgZU
oZ1XwhszKcxASSrVhTog1Qh9pBMjnthjWjIayR8eGYCqOmZn5NwR14JoLpHdY4pc
eu2xWnrgrPL5Zdig/zHWJWw7CVM8l5+xD9E6cRg+OC9jlV2LEQb73pR8SkYFETZ9
39UWjs6HCqNAPKztTyxYrzFQSvtu2fH/nCD32mK2PcfCJfJthc6Rf/ngYvIqGK/h
zQQbr59gBTq/zvYe3Irvg2prZdA7/culF8R4xTkvQfDtTI0SWhMEUhBKpQsROQ5P
E8nMtNYKvt0jitV0tEDc7+NV+ID/rsjKm//gRs1hiJA4OMXdnBz8KbOEIf+736zT
YL6sgIBcZsr6QoMou9su7mf2i5eP/dndgZ7qiC8Ww14W44IjJa0wo0PezWk5zhng
JD8PxVO1u41RPGQscDvC0dQlwt9EwluOyQNiCK73ClqMKgRPv33CqIrkNC1fWS/C
1SOkOjnazTUGaCB0gVqq560s8Wma5z+Bj2I/XFjZhMdX9KGi4jYIfEgHjmux7iiS
FfBTZ5HGlawD+5S2NFTZAcRdWZ8pVQk4+WTl/6v4bZSaZUfv4JQjwNUIoSllZriZ
UuiOxBrTkeTzqVZuIHeC2QU/3rPWlMyNDY6EdNg17Ad3WvVesKF1owOjHF2HXy/v
Xyex1GpUgmLXum/Nnl/66tPPS8Zwp8K9SaEZwV0J2XH6wn7yr8anbBqqTbt71ZmI
ZV8fd9JTLg8u8c0vztvAgr+eNWIaiTci0eWxQkADuhzRjeHRCbMy+CQ0/GflXQM9
XEITXMn+8tFc3h8K99LmG5wEX9YpeYYDObLG/knGeIQ2XRNpl6L8/z6avA/GQMf2
lBynoaZLfQjvY8UknYiKCBOaZN4Pk3J56Ij0P9FjKx1xJ8mSQf69LdLxV2/KtV9p
F+20eiBB8KZ2amAx1S0kNMD8todtsDgPyjl3ICXhOrZfX1i9s38Kyp+d9nE5s5Pz
2QN37bcnuhexHUdORo5XzDMBrTI07ocmutFJrzCjlq+EwMeGfL7cvnVR4hmol5/S
toje22fsgIERbtnKTGEkvu7FRTfSxcGDfovJ2cFjnW1REoJLhBO3z2IeKgN9ECjz
MFLWaOpCdTR47yRlY2TEzF4iKW8OfLZSsEzGsegQSesPYZ7H/ys+hEjF3c1wr/cc
2GcOYr3HXqdNy7bMTa1K7tKN7plbgo3yLE4x5XepiUITR17j7wL91HTMMRydamo5
XA8PpyLXurDP/neb+hi3nwxrXOjCCPUd6UBBgeH92sGczx8NlhjIjZgWFCcWdI+E
mP+MDNbm/Yg/EZVz96z8zScewINKsT1hJKcpIiFNbniEh3GrFJfogcUA66ktWwIE
d0IeMh7D3IeyK2l4STvRKyjQ/ZS80hz+dRVuQd0hv8Aqwt/Su8FzXZmPY0A3/goJ
X5PcEefiPvf9i1cGOTMRin+jPo6DT8rPffqvyfXWQkcREhIb6cINOAE/2yGu2DCP
hComE/0zpHFn9VvG13BAU8fwqZiI6DSRkOXT+3tKJcid4McjZyMgEOs/0mYcrqaH
jcVgdRUEwwpxLdwWPiV2EBbVwcW39iIQjlVHF8W6PMOtNIxPw+hBpSGB0o0hKdHE
/+Svf2ARTRHfTSgJ0t0lWYIEBqwOaXUb8rMWKS2hEts4WIVsB2Pp+jykhREST856
lIdu9biy8IS428NGiFzLNshnShw7n1ClGZt0XFuyE090f3j51eE71I0DtnS8YnOd
Kol993mUijj2Rz/MbEhyHTZ7tSBCYBYMvBQokMzP0bB66AXSCEyz5HNtIdZeWYSm
gKgJDfgO6ZQ2lMzWr1mSUMoH9dAPTcwUTmpIydcZxd5tUSbS+WiLl5SJr8s1Hdnm
8UILgnNWkydVMUNsqeJmoZPi9j9gX1N8pvICJPiMVqKvFnFCuU7DIm4Q6C8Q1IcA
YYD8RERs5PYi6RMESW1DxUgGcOtADhXNqrUVFqlP4Qgk5eOG7x5TrsM4JxcjIro6
cDC/GnxSxEJ6KAouAyxtUpR5lw6BlZO6J3RyTRKrkKS3c9AavzmUw68A53nvozjn
fQvk/1/5lAtR0pAilimHPfJARkPAZxAYBYoULgmTFGarEQVErsdTc88h+7UiX+Hn
MFCf7dbjn7gSx7KCCOfS7j536hs/KjbZ1f5rwcVPAPSKSUoSJrZ/5SJ6/qKW6R2I
hDMvhZakQemSRQhU3qI5inyry+RXHxHo8P/ZW7VTJ8l3rklALp3qqw7HZGsnTZkC
C/IXduEc4zbDo9DBufVq1deCdcyhU97jKsoYw4qehseDhQ90WL7Wx772iAgrWnnB
TFhufvTJw8694HLSGNGbhTImI7L0tuT9gh+LRisWobf1/9fKAddOqTuWY0S9yrJI
UHTmXn/qAClGlODF2fUpfqyhzAm/pSFJqWGzVSSYDgZfkTa/jRo9LCu+1guoiACD
3KfTmAigANy/NgotLKKgnZOI8GU/IpLUEPWiE/GnxJIy5Ct0bU+gfeoKeULt7g53
EakaTPc0WNPmiJEwGdLM2hTa5pOuCpkjm2cj7G+gLlQayk3ffz4nepmHUfSEf5cK
IURiFIY799MNvR3BZgyKhNY1NEhPmSMI2InPPxoti0zWVO9Ij972vb7aVKXDRbfK
w2xKxeXJLIblB9Rjd5lqJJSdkuLTbVj3fg+/dacmm4pSB4udwgnje6KM3wzD8uSw
feluqj7mzGnoMAC1IWj0yaxtTyHFIiJCSUBS0WhVDNCvmUPTSdIDmx+RjJKegyiy
TIfw+BAXY/lX8FHax2dVTsKY3wJkA8hlwu7mACs3PIRuLE4n1+19XfcaIy/wNB1I
Brrv3FgHjmK3DUG0w+7jkfm1lkmptuFl02StLKLl+BpX0tnN2wmaSBUZcNo2DwWK
i7/0ZtBNHvoEGyf2qVO41RBSEtFenxnwC9ozJdZAXaDKNSDfsfahWvg+g0W3YhBx
GzIkY0G+RZpWoPO9BgyPHal8A74GHC/K2ug7qSx/KlB/SwVBO11yxoe4xO2hBnvx
NTZokG8RbiuXeggtLnntDngVE9R0r2m6NDBj2K8XO+zvUc/amvAztbwXODsV6dYm
cWgRjGOVd3ZfKrBBntAZek1qbxNcoX2650eeKcx8pd7YL7EmiEwYc6e+447Fqzjl
u7nGnBaTIppMsMC63lPfdT0+hyY1BaWP1R2X+pP/DDL/FkVQ/jr8u7TIld/yaMJz
MJB6de2IX3FfctelZSjxb5OdN4mEH2Qh20M0FlwS8pMhfXJ3Bjlr6zUBpvjvMQ4L
pGfIIuROHflZCsClTnqEFUXsn/2vz/QDHLeJ8PCLS/qWd/4C49MgW6tJUbSt2b8z
HGyh2Bh6FNu9FVd0mAqAFOsEoMSuB1mfU/k24QGZ7nQH5g9pc9N2mGGzv/mjjCfG
qVoZcOjYT0tw3thf8TUMxce0MYq4kvV0Ov3Kkxuus5IpQorbjWn0RCshBiDMIAtB
uh8EKue/bJpZVjWNiD1kRS8sBKaJjTj0pBVHmfdeuEo5c8WeHaHmyI3pRELUdUA9
sOod11/Dlcnii6oBwpmBmyUg4OtsFEJgRv4K0/5TIO2kNJRPuK/G9mTmeusMb31q
2/tMaSL0vwfQL5UPrlJaGuk4jJPjcolz/rmtNPJ2OiNyHR6fpVftVJjOF+C5D9dC
Igg4L3QbNkyeUjKkP2WwwrHSBa3ht74WDwbINOMxf/jlVAnPi38XU886JmLx5l2h
XbehpHlXNYf7y6JAoPgrajp8xIKogeCjyjOftovKXkCLZosDNqmaJfgaaUwHax+U
Wj2+4U33EZbFfL0dGki9femFk5QfZJoYe1jjOd7vBKm+Z/pZnqRL9YtKJ6Wvuzam
le/NjGnR3hZwMGRBpY3oXMHfjqiH5F+7JJfGvzwyKFxLtcWZHVbccl3cjXhf+ueg
w3GxRISk9yFArDWSCWT8/ybiIaeXUoBvMm6qGWw1qFpUUFAWa1RCeCBygwtD0PTG
JAUvPkIDUb1ymB6I3Q2f/XfwzEHROBuX9HMEAhXIisdhav1OaY7FWkMsORzMmcBl
t5wfdQF44yRAuk9Tkxlp0sU/IVV3r68QS7IhQebI+/Z3mzMxmUaDmZVNnidZ5rj2
rhZVjhaWzi1GozVZLjM6wm+h1VRJUOHwc5/EG/6/pzlwMX66d/z5vraoGZoQB8Hz
G6RJ2CodvUOdj3CzPVyg7fiuW+8mj50MYF20N9uU33sJ6wvFlm//A5j7vgIejPdU
faCcHZJAtZzYtSXk9J3lpR8qR73y7QaGAtSHtEm7Klrg01uHXtVoprBLoU6tDLrA
F502Sxnk2RijPktew+kJKMVDorOFdKzE0xQLPSlREU/UaEFglGUoKoyu5FZNSrfg
xQXtEdXORD9i8K2ZEwV1JuAmxxLgtxeVEUhty1hBeFazQhN489W4SDThCk+1A76r
daHLv/7eHGpOzbvsSgFMkvFJhwBhzfoshJ3cCvFp/ssq/SmPkC9Z9od4DsvQw8fs
ibqSk+wQcYkqi/2AXpFFeqPw8Ssnp2fUUH+zDMU3EbL1STCrJC43apqhDF8MBeNr
1eus+zANvQVu/zcnS4Lc/MatrS6pyGgHcFXX+51atQ52pF9HeDYG/mjaP895bAo6
Uzrq7R+6izU41D9MoMfiw97A+wczKYeFFfPKpiUVIM0pqJrtSOAgGvX9R77+m0Rp
mJNx6cT5+aGl/mx5prwgL0wldDdeES30CXS2ZeOC3Mqf6btA1SX+torWncBYRXJz
4LymOYv3FpxHufUeevVN+Aw73ChkZoHeHv4PC969GROMlZ2q+Rt5ASRbVXgFn8ZU
fzBHczffq+QSTVvSDoigOaWQhvPVi0ZO5fBDD38WPB5LAl9XKzU+bCRZkrj0hHXX
kYWJp1lmrBSytw91Gtm8wmRTwCWmMlHuSfY/eTiEewtIxALdZyupegTQdeLWnVaJ
MeuYBWLCF1C9Z+8erhE1TqOKKGWsGRQ3H/mYPCzUfmMAYeETMfnoxmDCNj3G+zcq
phijGIFUzor/fPqSW2pPorS+4WnELmK+oQ7OoQ8qf4jABl4LItO9WKOYoYk+3aQQ
ixcuiI/kcOE0cJ+kjyfjRKjzmqn3ySvHEi+efS0lJXI9/fsU5z7Yp+DAnwGBiFVa
UPOsIdkrkz2BCxkVh0rXAt/CqUxKxqOp+YakSXeSW1V9nupN7qerKisLRkYCyjgL
HxNiBQRDPUAmMtRi5O+kBns/00FrnzfUFE+hnMexcgFxyK7D6t63/7Ueb7Y5USlg
39uhvxuAHwNkmD2jD04jAKmWwnTOwGiYmBVTyn//1RQlcyhI7ka6fCqPKY6/NlT2
YRHxq45VarXGXnXA3oxICYCJ1wfwjvDiBo74yp15PtgTM31RQQcjJp+QX1+2mNwP
3mUUbQHRwFXZWmp1qaEfShHGBknF94C2aMRyocuQiX1oQTjyhfEXHzsJCwHYdyc4
gGoyshcc/2gZIq/W+NToG+hywO/2psT+0fJD/NAHtD5ZoZy/rbhdl9PDJ/VL0sNR
DoWvaQLXmIoUXavDOxOHAchG6jGKEm9cYA9zbbPxtNusVE+hyyrTzRH7+fdElYn+
AyUgtKDRt/cXCHQVMM3O2RP+ybFJka+NVzVnVOsMa+9cfBJzrJgxqxX3xgaC9taT
3NwDZOZgMHbqLn2QYlytobeouMYrc0FDqiUz6KXONpQpko+t1A6/Zh63DRYusRK7
Ow2l+jJZ7d+YUSI1gNciF9qk2K9qcG+w4R/DlreMiNxnMRcH0An1hQRJoiMMSs0q
aaRMihMdheWwk4XOr5YemBVRXZ1Jw+5UOAHM4blPzsOrSjRLC2UrytGioHcAMsQy
P2jNY4Y5vaJkXKsDqmPbhb9HuQpU+KP1HyvgZL982aawxuSdLlY0OTM2gRkncsec
QcBJH2nNQTQdmRzN41SL656/Q6COo9H7hHpt5U6eVRmLR+BAflPs3udOP+jYIspW
LKhjx0ianVzu0SCmNxEQW6lKII7IP6f3shD4DQuTC5TyT9/wKYR56pRGbSKdJ5TY
mvjvXIvW/LsuUT23Mk9jKnBWZYh8UUykX2f2h6v1s3AyrzK06YF22TH19im45iwv
r/Hgzborfnx+0/ls1wrnhCY/yDyNgtzK57z71p4KMKQfPr4tLJuCL0vXonx9spM/
LPDrnE20Jv5Ag/MggZuhHwRgejNIyCGffHHYWTjTYX7g+zBB4vMJaNOL7bzrGBm3
kZMicnDucvwCL2LaXYXerAEGJ81faIoF5X0pL4UQoALIgWlAMG9AiqilNyn7jntx
5NeKX/BaLP4raSVCLZCq5Spu2ceuvbzH1jXauucXAbbGdhln9XJRL9DeDETVyKyW
2RkXVzpI+NUfAdNOrGgU6toVU+oOlfOJ/UVuc7AzJ76HqXTfORbEdxo8yQ2ZIZCZ
8wJDMLui0FLCC6iHYKnbKa5pdSgy6vwRB1qirPV5rL0QFjJSeCNO917cgLblcXqQ
jmhkEZEPidJpD1h+8e3ojiOP8gMwZ2IxjZjSsIS2F9Hz4on9ooNMLu0NLzpgCJ9l
FH+NACjlPqhVx6ncwTrHIVDxadFj2Vq5tVBnTmmn5OQ/vCDQTIbAUU4i8Kc9wLj8
VH84hPQWXY3ShLReNlkx8SbhyTjSI9Nl1hP0B2lmlQpmo980o3eEBb8vn9P0xad2
aRRCLTv7ZQluMp6WKYXQ0vLN2pTAzPFZttTir89As36ripy/Jq/YjQIp+a37Kr6F
srW+nV5iO2mS9k+2rVC/2kr3ByEuryA9hPL07rmVgSyvyH66vctCoR5O9X76Mx4Q
9bn/aox1tHfljqSKt5BTc8Ch4q8NUi8fAdxuWd50XbAncHrnljuz9/Z0cNhu5QLU
d7WkUN/fvqqpUPp/99omealXuI0udVzrfuL9hlJ5C9NtzAUGWkntCOx/+a+RRGfy
Ck9HB4eYYRa9UUrm4YvoL/JQwVTRxVsah/TewdAvvu/p7uHE4Mk+e0KtnJP8aXoY
f+4Y1bUUViSofpA7qeHp9RsZUdeY5+WePc4qTYkiNK/jMaNdIjc+HRbhRgVP/OjS
CTQciitJv6tRYURpv+ZrcwHrdBxNvCYywWN8+kVZzuMxude9mGL651eRVT9ojsa9
TOmiYmilDAh6wPSvm/RWxUQRMqexzdJUA3C4Q7VKMEDQxlrlraw1B5l+lBTLjAd2
68PJJGLq5H+E2gKRojPpvcMdxfjeiJCs7g5q+gUfbX8lM3nxBsSOz4ZKzmg9MVwd
wMBma5DfOShc7aow0NxviUPTS4LM9bIrif6zHm7LFkjGF9FzNZvEa2sNTX50wM9Y
KrRf/NVFXO2omxu9Oc0BSdU8kqgc6gUTq9O16/aRnYcW0PDFtrNyMtlquGQXP2Tk
61NUGCUjAxXMopm207B3/2apa0Cw/e65YGCTYNTeK+AxB6R6SvqPT8wkNc37f93W
ZpDvt4unpBQf2+mAIyzbqanjKLW2KfvGQtgWvriHVZkc+5bsHUdPTiglHkwbuHg+
rZHkxCDrrtIKLkbX6g1/HyMidgm1iNaKcIMAalwW6rdM0WGKz7PRNx8Mdx8CjVIl
87rGLakg0B/4Nv0ScCEMQHdqYLYxRXnaJjSk6odv0Pcy2R0FK7aZaq660Vt5s8Yo
lhIPQZOZWjhKU9k5Bu+eNewNYAUmd8j+3K4A7ucxrIrr/SfQDQ/cEyFMT9mVapFr
mWI5kIIgmBeFNaaCdHViOuPl5CH8dfVucRJV6jTl0QR4SPKUYZgi1bZYerSO5xV4
66kZIqHmtJaqvAZ39ify61V9Xfzpn7ujMBHpXRxlLG0xawzS2vzVZxdhrE/Q3QnJ
EPeIPIJKnvNnHAAtbL5ng+tu4/6oIEA1nBBineg7GZF3AO3c75dKRKWDQKoO+QLF
8/fvO/varGiToc3z6sqcvhAo/jl1eBHUn6eRKXrZ4vyTHvcHsHljboiWj4UY5DsW
TvNRusGLWN1KYFAgGI54FpdFzUYAw5tOsjlugRawslyb8dERheeEAImQ57y+zB+B
SAAlIMSjVr6PGcF5nmrELutfA+6ckB/vxsBWiXu3/9vUq8xlnHJ4zLWZkN1G+dmO
lk3NnMQpMktBNOQjEsue4OH/Iho7pwuvy5um8yoorYzahI67o2SzB3rHFXecIgw9
lnHxxc35GhWvOYCsld7LU2NqUrZCLqDFHB3/AckKKfL0qUURnkK6MMWm04rf4B9p
h7OI67I+zTwdl0H2DUNIKSR7p9wn0RK3esg8KwVlERCSKgf4TXU8+6+7L19kFZGv
jUZ3TJ+ypelMVHQ8dimbC3KpMu/QHJ6t5HS09aCvFADza367ahY8LxLPHJU1P5De
OZ+koo8lPhbjiPxqnx89p6E+o+jZZg+QFtn/x3mkrKXe20IRvwEZ1YtToDzEbGrm
aovb+OKhAkorOLsFoC/RpIvDqLCOUmtweGLwYAk+OFnP/b86L8/O8dPZE9Y3tU6s
7C29hY+i2sA8GBTQ01TSAna7gAdigaVD0dDB/4OoIRg506Fo8TGc3DOTIFdSZfUG
cDVOOJRwB9JMHU9GPFRd5oApRjrara1yMRlSbrQp+B3OJLbzNKPKeuxazYBgi0uY
oibW5m6UtuQA8R48ueeT+aLs0r3HimrrpQX1TG4PGj3np9fobvgiqo2ixfjfZxOD
L13Q6gzY7FkVz6tfv3lYVN2gqESQ3REzAgbqDU5t3x6MKVq8hXw3lDZMRq6KEJah
7xeNv1gpSKa7Z2kA3e21F2LXcOXioCnLBu6ktqSGP8VGj1lRkOhUysq5MUA3e4S1
s4epLm/z0L6TKDhQHaJCFVP/bJlXDZJ/i7tUES/xpAlTwDYfQZ6HhW+lcoH9NeGp
CSAZVu2pONkICDTTiSSnZVeJ18KSdJgY0oxYJN1Rcz6jA7o/4WKgMCYYVZ06Qf2t
iH3HKmdgQftkcN195hpHm2DPvOKbFBqs7mXu/tmLjsfyUNIuW/JJApvgtu36zSSH
kVTFIpMrlVFtsz5py1fuAv9NI7WMFLT4DreQ9LoC5k95gdWvUGBllv/QsqMLJw3s
R9WOAMo91QNgv/5FvMdC7XKar0vXceL6UYdcW+HgkZuYe95HSE9uhgZAMXx4JST8
FlAuz80R12CImoOf62m3Zslc58lUz3VrFJID6hcP16KgY1Voe0sNJ1yuNOdr5F11
6djeAYbSzJp1HQ+4TDpP7cdxsOXCCDYHrXIjkCWzQkJeOvgUB05i0xccA5+0bghf
Ro9o6F4qTsA2rl1ndS1G78rphIeT0cuy1YlC0GSOoBUzeR9n2cndxoQCwtghPqmr
dOJuTHFOCItq5QTCTS/bLHfMrP0+d9OVPC9EE7HhCtsMr9QwiFKpyQuj1Ldpz8aE
ZjkeZqfc/IKn5KxI1G+ZAAdxCfgPs0/N8f/UQcR/9DtSw/I2MAnxOycKFOEzFYS3
Issv56D8NNylhP/e4LaLJz16umo3PyzNSkFAtQYwXiD9bvqBnEANtBOy9wAgfw94
ZoYgCE44ROxagULMZZKf4EbTRTOFKhVMncwdgmavIF7ywsS7R/6G221QnFMf3M2T
2Obl5iZspCy5g15+WgwftgPv0iWY9SOcZVjNdj663Cp1hlkR3oUAZ32WKEMHOlln
9lE+U4wYDIuq+IdCcOyB0GtdW397INVHaxocG1yqWufwOsk5nBR7RblmC98EIsHw
SZgJ/AA/jqzUgWS/zUC0E4NI8sCm+PrC6YQ/csFYKm6wHCI/ZI9HnR+qNtnDk2fO
yzFKZuan4GCL8KbcecmiUhHiOm+E3iRgCPce2uANgso61VRBvUVrSDbvUnUdNfd9
VjBdW18SH+rf3B7rfOHK7Ajg6xScxBG3lkzKDrFNh5T4QMcBkOmwn6KZWW0avYj+
pHz1S9+08O31HKfdT5FCox3P8oXspwjDxufbEee4se1DZ+MOVC7UzJcOnp/XlkDQ
gefHm18Y6b2EhO4oi8y1ceG43uStQnOpUcS8MNw6eM+CmJ8srVjP+L9AUNpf42oy
OK74plMRVZosk2EPFdO5I5zIAoilnDrTdarX3g6p/jBYfqjmLmFSkjq+8KSnIRVo
l95yBF/UjdpoC4289gMCP8xGg1S65NlSdqFmflxGpejJuYhn6qkj3XL9cflsfbeR
quP0+eRUvfU/wE01vxWpRh5FCjC8WTEDf5MRcgul7RUnTNpuyGjz1hBv9kJG98CL
aM320dDuY9yGDxH0Lywct2qy7ULS7O8rESl6yQO2QstAW26hRoMp4mRKezHN7Opi
sEnLt/5jSeWYFoHTT5gHva/TQqC0sqit8fYGCIJobiT0/M5GeAK9UlkPx7ux7r2Z
kilBtBex/VceppAtCxQBtNJTNjXPlhoNaXvyDcpMqRHAehF9V/78BzryT7Ah0f9h
k5Wu27GtmaZePcbFxQRtMtduAqWtrHHIJ6tyr+ZGjmkmBUTeOc36xzErdi+krssX
B8Yf3NfOXS5GGc6WRQb+HalNvdGCEAL2BXn6YHhZwCjB7oJTzFAUBbCaQlsNxzUL
nP3wBTv4mSCq9AXPIugvVDBl2pb43f6zk6cI7Aq1ARmyjbDtcVNzj9R+AFlOC+K2
2D5NlXS7FlNktS9d6ZEJqV3hXxNbSMMGGNrYDB3R++iGRLyYifAUjRG+7vA2YBAg
JA+z+6tDxhmpwFkyHRtLu6p5a5iq5bXxR7kLVuopKKTJ1X9cEDaMv5Lhvzqdppr8
xxaDTSvHpHHUtY/KEn23aByHK0MWPXoAUQF7Hq9wXjrmZ5fL5Gp7pa4coAfofMd0
Kjc2X7WgYmBlQ6pRgFKhWflf7bAgvBybNBxf5M7lqxojCi1xPxyRgViLGcUa99Jt
4vsAPNz6QYkEPKWbq8iaOGag7jIMohocrDVPCm52ZAhPYLA+a6ZH/P24euYL7EW0
fYpTMN4wKXLp+IMllB5K62uDhvnze04b66LZkWHJT/RSBfLvlfVldkbzLI7CkKvR
R7koS/TOm1hZ2/skptMdoVuB7sKLFg/RgOFVE9hDjA/Kgw3Adih/U74EuQMR80tN
WIBlWod3H5et4zdwjB88fK6FKiOiDBFLADqpSjw1skroh7QSqCG6VnLmZrm+XnEV
GObNjxAA17ExLEYIPxU3x8p86u72Xw/uMBrgd0wYdUfCKZJ1r7GdbGA0PWYRaj6z
U1ehbwnhgCxTrEMb/BJ2/ceNOEkDjLEQ6z+CgkTXEDc97u6x1OzwdDCVLVSVb1P1
0J/t0uK+lw+Y+eWHwHhGfOT0fTo0tmZDx2jlFukhO8FCt15T7LurfSVD07txlTu5
76o/NAy8HoiiWvYliP4rQN15yeam9zYQd7c0jNMUXVD0j3S9RtjzGrAZJUDRmloX
JbTtvIZ+NHOool3DIDMUUFxNrH0LrjTDGSdQ19dJaN5sEQif/dXSwWVsmrGT165z
wOuvPcRht5LcxuLDfEIzE5lkKaVMNF9vxO+EPYdMZX4djETZ4h1Yy3/H/umGhPM6
hWQR0Y6l9BEP3ckoKs1IvAPs3PrkwiO9bqO07SwySf5QJMo1KDeQWNcikGc/mtpa
GaXas7CYZNsC84+qvZ4khQm9Jcp9ws+y7xiFTZle9KLVus3i80fWEmgVuGosbxTm
51crxQPW7vdr8blIjLjucBsSLfMm4TGUJPYyoyV5iSpso5cbJ6rjuIuG9Ik/7blM
idLwFHgIW8kbXssRPuiZ5Vo5BFhxkwSHSG/9zbX9fTHQJ5sqahRvW6TUgA5Vedg6
RJG7tHs3E5RCMwWPLjIQRWFihGwkjMA/Py5VO2Jh203CJwi+7CAwfje1aHqnUVj+
07MX7rR84um/oaj746rtIbDNFEE0uoQHDfCxhnuGNNOZbNhgKTbxKUS0+H1mun8e
cchnleyqtrtx7WhYnx+OnERLq+yM+P811ZFv3Crss5yUJWZaiw7m3tyRHVtyB3lD
wiOjpZYimUxDZQWvpFzS4R6YjrdQgWJlKpAXalmu7inJmRDiKC+m1/pZrY0XmNdx
Z8ZfE8iux1c/vzntbCoqUPJ0NhW2eQ63ob1TBTlU0qLCwTKR3oov40FflQ9aJhvY
QiagwHpbLeK8CJXN82sIv/BuNUwp5d0Z74LlaP/3itkPJsMB7a60ViEkmS9RqYSQ
TLhrUeyBCASBpKwU0Fa6pxIOwoeUelTgNNbYswdIDxT3goXBYqetAziaUXvB1cdb
kCAwcExdgNT2veqvVMI4J2/YmLTtANAr3Xq6/sO2vJtUKsaMx1qTT9kzACKTZR1V
KQ6KrBU5vlAFEUkLwnbV4272hmE7v//LCJjBvQr12AvPWSwQfQ6oiactMGh7LvOn
05Er4yfXJ/Fh4bw+mtQpGNjy0FDz+/dT9oGE6ydWgQcEhSLK9DPnkWUDZ5ewVpDH
90Y1JIYhrB5q/2a/tJFwNrLv/sw6QRGR0HyvirClnRcbLkDukvfQLD/z/I6KuJmx
pZhfZMaNKMbZqi0pFYv870mVMT9SQc+A943ERieTMLhw4PEXDH/aTOBgCIZfsZ6i
9hGo2e9ns6u8uMbt4ac/5z3HXWVohJub6e7a254J9Rog7w6tSGjxqqQaPaMnrAzj
kcuuMmaHC/zbWEsH9tQEtE5qhUew6ttbEJFlb4wkYM4qHs2Dw2qTuckvjPKHudpN
sdguzOLiAjjJ/9dn34Q7S8S/P/DKnDfQULmW0ElJS2wf0JLKbGXvq277I7ZEV6Ue
jJnE4Z6Gk1kNeP9gzK3JZrEMz08zaGSTXtqJq6H0VbqbzXND8fVYRFClKe7m7c4c
DOONN41WXwmWDGlv9eItQ3MT0jFeBlnFfCdOsiObTT7a2rDOsVxg3y1uKHslQOgK
u+QbrDXwjZz98eTaaRbccT5R+iw2Q7PJdpWxdGyRDzh2A/ZJkI5Xfq5O/xTwdz9e
M3NuO/R1BzEhxLkClSz6UgUUv+hLQJjImxbAVCAm/CyHj5zWMgJlhUemVSmed9+L
4F6OMOHMKum8+AyUhgeaDT8zth532xXzD6+FoTAeT07Waq/hmZP0qOLnWD8Nj7GH
21T6Ac0ns7S9RajTeF5XxegqZkVqvN/HnxSVm0mw5Dz100q9RZ+TZTI54o//kQI6
ramIqZ9ySVCcZnDA/Q20IdmEBUJPWAxz+9kjZqvik0na8o9lGV8r1tT33m+Rakro
NfEPHi6zS+FihXnakx7KhLsmtaceVabd8WX8TKEqVgs/zcj8PZp4RKUbvULSLJI7
gV3KtE3H+mkGIGAFD867t8wp42NFQQmiW3wRf4re0nVUvOOB+sLTnN+SAYPb/rMX
cuH+mxL5Uy7uS9mX2nRKNcVBfcSrQF9dISrGuQWolpDiGithDFTFXFVit+YcCGaV
eevnqixFPXG/OXIhGlCKdzTAG7dISkndCd7laRfdqm+xZDzXcweCAI4+f4XvpXNz
mkMyNoeOPPp2AczoD0fMFWVC1BLKlrJWEwjyKfCkrL488jOYjfTRk4QzFTjtBp4s
GTLsp9MW+0SehHjrfH4/gW19HZtUbyQZBIGRNqtGAfbA8QdCFJLy7xkA8FeFWHMi
VG4PjXkp8eIT7AhcB9fzBurhFUJ2pAvxioGlMLMhIuuPogMiSDuVqac4MdYtRLk9
uXkoFrLvCXX4fdoFFzHuFENnGG/WYa6EymWkI+UXcf49E3kpHIH/aV5LSJPNEtwD
Jhz1qTLyr9t19ghnWAastN2DTlNfL8MgMnkiw+9wVszX3E78sUrcltdmu+yRsswg
y+rggNagB2FTNlTFZOog6KHHoed/RYJDGEo2fm6/z7VTmQM3vI1PXcLyZvLXE/EY
xgGMLjp8v7mrM93l84J6NLFkvTJy4l7171B6XvSC8ctO2pD20HRnDXp4fe0cz544
rGqb2LQoXeviKYb0vifc/iQbF1r5wRJIhq9NbTCdLezIESoZPeVF6bLi5elPJk7p
OvhQVswwu2ElGhZ83WfbVtab3zK5pMaiXHCnHsKgifTm47kNR6ZiExo8a54QX6sd
Fu5x3MDtzA9Hiqva/h1BkdSamMGer77wrqtdoZEHbW+QNnn7zRez3vPymLeHzq2O
LDI8OdhnumysCUp+1kROWgXUrw2T4fsF3IlOeOcW7KNywwhmFO8rwhKAXdaxn1R/
uBvJ8uRGwuuSnCwSBKe4yb/pMZbbo0MoRxG29Twiaq+g1y8n4TN43swXD+m/OYla
I+w5bHAHyR62AIOo9zVjwFRMn5q9Ga/fHlQwYar61Cl2Kev21GrK+lCuZxxv1ArW
0WVhA+/Pi0IhlJ5qIjcSCwJGIX3yNEbRaS8ofAg1KAAwOmZeLzsOZfLcm8k6sTk8
+ymxjAfImcYbqS8tuEN7SVkOiGfS+PuUoASYij+mt0Fwr1jS3QezIsNVuZboyh7+
3QrsEtm2b0AfwtbHwmzMlJpSvPAU90CZ0uNbkiFdRy9RJmlwjUSlRn2XsgOhplwz
0+8v4dYkjVq+wWQn1i1XlVDYefQ3MlVL/NW2Xz0hB/LP7TLhBJp5+qxVUwcQqpUf
Xb4hKREac7Ylumk1W9zOTCAxYLcVkoVdK7RuVJxqcYIdbcMAReWhJaKai2bzPbJy
xmg12yPFS48oZB0VuYrOOulXrszZoywNJ1UXPbnO4FExnIMxceOjOZuc3IalJBv2
NMk42owSRhSXTsWlLzu7SKOICIxZgjTXJOL4IYPi/7/NKu0g51PNirFhgH93EMJw
DeWNf+uymO1uo3XRqK5Tt/FLtPAyZVRRbrqvZmUVXeqeEGGce9g0MP8eCmq0q1y0
j3RPK53hfl9sb5oCSkvJdU+opDHrKBhqnweLO3Mem4D2lN1DVlcLEKrznDB9uSTx
NaN+TTSFksvEzj2NK+GsaQTixp4bGilPoPd8HkyRz/O5F+cOYaq4yXlXqH7duc9T
xPrnpL8L1LZdmSYG9Z1V/6rAL1qOZ77mH2rFwaej9RBgIq3a9SmWmhFcbvTbrh/I
4VSYkMUiAo9XZrrArIJIx21L+Gy1cEdXI5tYsH4+XdXzDTHdVh4ags21ewGS9iEd
ddraI2ZX/k6JEJOqJjd+SIwYiWmbM/RPCVM6VhuAb0oG2iTSkkr2Tjk6kqb3/19i
gbTKh/qjEVNFte7poziSE0W+9PONRvSfbKZH2kpb2fIk5D6sPURTAwVJRy8ZKLfg
g6SWVA6DNz6DC0wOnBHr4HYLx0PkRHyYfmPvh9ebgiUo1g3FoKGkaAkVUe+tNoJ1
vxYQH+sgJ5I7xQK61bIOlg2efw2V4wv77oD1KodTWk2i6HHyoAUKxyYQC/I1GRfl
dutvSU6luczOYJj1J0YTsNpy49XFVci15hUqApqbkQ1jiLzqwkZQn44dWvIXWcnc
YfL4PwUubzEWyZxJJKD8vdPV8Uqb9bqPt33NMG1YUSfKl65Uyk5JUpREzROQchcD
8cHVpMT1UqRnar5z0Jvs6LmY5vJyQ06lwkaXXlFP3dJ9Boc5hG43r4EA7FS6l8D1
kumBfvGiYcxJnNuOm3NKZ/MtMkyIrqJ71qUhuTehInvg/LMeTFnby2P1MRxolu0q
BcQvUzplbNT7tytNVGTxWFk/CrI4uCaDdnP7EZ1ZDnSuJzaLf6rLaVRrECxJV/yf
PEgyPuBl3JFNyLVZWlzy8MONcKi7EWMnwyz89CXRdadV+LutgOUTH9fNG2sp5Tz4
ugfzqDSKj5t1VVPkfv9Rmi2UpuGUqZllCPRmCHQR3RxJlrKNrXilVM9jp9t6J8tP
`protect END_PROTECTED