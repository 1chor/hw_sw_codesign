-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IxSOEVKgkrCpTwH1WKve7bjALP3RRI7WpsbyK7JhWrUB3ADBmH+rAlc8m/tcrJGRK84PgAFzuAGy
NI1VGAVpTfwAd8f4bjqRyJX4B5nky+da9KJpIebcVD9KHXPPFGuIhcm7okVopuIFeW9+FPVLDk3N
T4H0pmTA7M68JAqTrKMpMuC1ncm/XxrAHcsVbYAUNCifcv8SwLhgwx1iybM18tgKGo8qNEGeeicV
yDXQ5FdtmS1rYwNRSgxIlkhv5yYb2fYuLQ42AW21wGi4MS+3zIZRMK5k6lKamhGhwHgW4LdNEfYE
WmeTnnl3q0nNPdq6cbHVXimFEtWG99wgukn3EQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13104)
`protect data_block
IW4wYfTGHMcuQl3BcysjQ31Llh2GD4kMAUaN/u03ass0b5Xwr4Yvz3A84R6tfZ5iXy4arH9XYJyu
g+yH6OIzcKnhiPDS77iah9jLGgS/nnC2w72IQxpEJ50b5TPWsxgeutUCCZYUsY+FmrK3ZnLPFqxX
cZCO9/BBEHuONPKrWYlLcN4L64zbujr3KUv9ZDNv731TsbLWkFr+oQ5fceEEVxDyae0kXxScYPTX
U/lQ065/JfN4ZP+UdOeyWGkC2CkNTmeH0U+WXi3gpH0iCdMtooW3JvcKxrg5XAVVVBDkcilblU19
Atuae3avNKXOe0fUsjf8dsv4PGEsJ5JksTD7okymOZcblDBvwGt40l7wHeO18iZ9ihsKYmpRJEmr
bye8RReqGXyNxCqvRUh3lA1anSEYD05mnE/F9rbKNwtvAGN9Y5ZoY8mUcYK9ZeAItV6nHhlUNxAT
Onj2zGVTqS9nthrC5jiJv6Lnt3YdGfvcTTL7kEaadTIE3F+Gz/sOdf2vtznrkrqiiZIUdMJc4jXj
ASggGx0DtmMJbiVd9unVwx22pHg8Shymrs5BX3Z5+GCA4nuCwKWce2sgOyT57mlWJtDCxgNZ3a1b
i051+Ci5X2Cf12cSmVWXAbqawKGh6br8KA4o2zMd1GHTdG6AhtqZfeQ1V2pahcFLN/RZ5XqBEYs8
ZQ6HsLULSu+2HOLi6cDJDblg2C4iTdshbzxbnj6Mcd89JPBn1p2ACePIif53EC0iwCyagqAvuC1T
b+w/oovxm2GpGI/oa/67cB8a/e5l/eIBrzntQT3rUSpQoowYJ/+gbqE5khpMdlzqlXJJEsHXEyB/
mfd5UvF4nw++cPh5m5IZgguLbb32flU+iEC1lNvkBzuhHadGnvI2qOhEtEHgQjYcEONB5i79f9RD
jkC29lL4WKbvgj+PXfD/2j0q776agC2nBP/UdW2QOiRhlfnwlNdvagcqBeeGzaVN+8xoIDQRcjMl
gWanf+e7GZxyMWGrKMYZ6R4KcCC9hQlB5yzFUk/2TOHtWO7va4x1MRcvOH5mtKxVvNAzSynbWN1E
fH9DDim0zFVGcwnLI4L/vzpgxcaUaEzV8fhJDoCSTR58kc2FKnaBdh5Y4xAhwCfXvlA1v/SWnmH/
AWj/nCqaIwYAQ2BJ0KRaK1mingElcu+aBqBngyLHvz9geOP724RoDS2dE0s5exLKT8zY+hQlrK4G
gWnMxhQLk5IO4qxx7CJqpfAtoak0AGm10YJiN+3nErJwdsLUNxLSGTWixi+ZfCP6bUbtLIE2QhOq
thSFRpgsDkgdj7TpDYyTxWJbEZBnNvtFoCZ1ySv6iDzCkZxW6iqcolffwgXhFX1y213aJ9quRsly
ZK21hx8ztwluYBAonwfaX63EaG2xm177Gai22zHFQKQKRfB0IEsDzGFh22KaYG39RCvV7SR2XTt3
v7ObdS2R3VTIUIzhRfspls4i7NFVTu636teuK2scsp/yPaYgL0lDesdx7a/E2nSywlELWDotnaI7
2TS49m6Xw8Nt2zYrEccIlGhVCv540AMxqVa7vaCH/dZL93c9pAjokkHu2UHlor3NWPyOf+MHrvJA
zVyTZU7DCuFgw/k6kno6ALJMVVbtPWAuuzdVhqND+8VCHRI6faeHgqGcK+m+z4OEmWQy+rzEbvol
LLhwnNRGQQ9YJPAes+MXjxNCW9MMZYwD7Z2Z3hrqEm26CL2rBdbcz368k93Gp/mxk9v51P6qnWA/
FxWGGZUcw9zTbHZjcUIBuyduUZG6xMSNshdJR5fSccxIrDDG7WqXx+XcJAc83wfzWh0ZHvcvl/BD
R7SlFjKhlybO4gxt7Hx0bQsTlAwOREIlXBAfd01Ame8bIaERb1vgAfgUKG1r6et4sNrhH12B7U22
jyVgMzecGuMw4KlcS6bFkJQTD/EwyQa+Z0V9x3VPEggFouXJdh5BsytydKPuEaHPW1m9oJmyVwYs
nTGhdhh5DnbrYchBKN+XT8+qmh8EIznt4Qyp8llf2DcmoH7Cih/Q9MEqCrhhSk0HgbcuLisTUiCx
0WbWoBY37idrArCAtSQCZY6IBAxn8HX+F1CMxHA/AfvP2phCbYkO0c41zv8dv+dY+DsKvje+GbQG
zDsSiOMHBab2/0BbPTNey/HeaAoObgIygTf0rN51SDl1SAHoUXz6uvKVZO530vhR/H2CdQwCRyOD
iCZnXUkK/NletKPwS4pu27Tr/NzDhRGtxQm6e15YOVjsHrg5iZ5QCTzLC+W2OoT6yBAiOOOE+0CM
Gq4tV/JDeWSMk0Sbb1TaAtadofkT3IaJYQEOdCSuyaMmFEWGSSMAY6nOHXQkT1V/wxCrDk96Q9dy
rHRKsNQN7O43K0cpnQkOK+vw3cz2idilFT9pdMGuFR9zeyyss5f8/BEybjpl4+T5qRqNR4f9z84D
1luK6QmWNYGpSUq/TqOGoEeTyrMEPA2ZGBV8DQvt9oYiGd7V/QEaJdZEF3a0s8QI9G+ZqW9V0dfD
izNe8te6oGTLH12RW+hlA9keIbXYDerP1BDUc3RGlk8HbsrzyGrDKhxnTE/mPrnFDMIzxdgWt/rR
K6SI+mbhaElNM8d0lAYINaeBSmHXyGfSFRSqs8qInD55Lh/H2dTsvXtj+jmlk5W1fvZH9vln4H5H
L1axlxT2llWM9G16+2GC8egyPTFGfycUKqbXuNgVsyOAj2BW35NogcL0gV2e4aqH9VSdXB63KZa/
7cnq1z7EeX3NvMTwqogRtIy8bo1kIl8XkW6uh0ShOxNHCqrPOOgUNpnvm6jWmOwqdtPf65/SQIbn
fXznZI8xt1B8x9LwMQU1goZFQMGgKi9axWFw3gRWcJ9VilaocE/RcaUbgxmZzuSj5tvJom3x5htp
y/huK7Xj6oJhrz9KhUcextMMvSywv37oU5kdRs8+lX2158fr5zrUrjkA/tmeDufIdga49w75fUV/
iLw0WwhLhfkpgSqWtMu83k3zeicClTAU73BI1Wl5PGo2oMCpNniKvzDi0mciKvElNV3rUWJ3nowz
gwH8IgJgp3PucSOlttHqzwq+Ln/3oZCWDRZHzgWOTRF5yw0l0AM4Lebwca9v8ZLpPd76C2JmIVX3
qERxLCE0fSc3wuhdXKNppPW0tneFRhbFTeKRfiasZywlSzN7hliuSKLrPEUOFSAncdMaIzm1r49+
ZZw3bd75WeM1mDjqxgMULjUgB4eqPQtocN+ods5bRXb4UehzQI4cLcmW9tDwh1CKNQ7zNCso8X3R
4cYBPl/jeA0B+FfdfqX9fbUR7SAiK+vo+y1pPsHfkqQ0cYmef+MjpP7KDZGEaXdXarbsZ3tVKPJH
QYZ1XU3pE5eMYrak+MGmBFtnsPk7TVPoVQGdKAPh2NbFl/9iCxr2Z1rU2tE+hYIPyGLkhnPwJOJe
ExunEZaM+iHahu7/FJD5bP99iT895rhto+d8OppOcpfH5a2a/LXrEdYYpv8fXBtIurP8H9Pv4qmm
B7sXE73q3Lyp0AWb27kEQOC6NDVhWx02ZKPT4R9D1G8FenJLkznHpxUEbGwTD9Gh9wuve+cWdJNr
6O2blbwVHlxZJ1nQ72qLA97NFikJ3UZXzRQkxZcpABq/WeyGUa2r66IG76a6uGlXOFkZdjlhs4BF
40p1n1+hMUpeMXDBXmXs88Jtk6gljOCfiKMApPorU2JHznXfAWRZdST1jYKCejun04HklcG6J20T
5Na6vuZPQZzuXjzX+5G1ilulBADrT2KX8IfsGLmPvrE5wVwYA7encsrP7IYvHqqXIwZv4M0P+ev1
8CiJToJoz00bgttvYG9onhMo3VGrbYRUSj7E+nBrHLfqqwukZZ94PiHQn8GJkYUkREm5wb2gmdvH
ZR2ZTmS+9nE7qmzdRPK5Z4syqqyO0Ld4sgWOOUmBNdEVnAUEDunxLV5yNR9O/WMIRUTI87UPwgs/
gi6PZ5hOKcOBpek1TJZFISphXzVUmNEOR0PjSo0QIZ7vYV4xGaWLxobIEM/1vxVuM/Q0Yu1ceTEp
osfbt4dpwUL9BEWKw71FbpgfIPdkkHqkfL57fGpGV3W9DCKthvOmIaPbK0yK7Oo5slsbHdkcxkou
PdReuMIbFOw7KNxkvsPp0G16uie2q6vEHWUw9+n4tTnhN5ZootyQHSaRkc9afZr+yJ/nJrvUeYJS
tTZXW2UGZqZlguD9aF7PRtEphk1cSWDkZ5PLNQauPVriAdplSaueT88qlfnd0gRjwMund3Nr0irO
jb89ixUAHB//bbFHbxKuWp+Qj1teC7MOEnpzziAqSBSgnsWcLi5U4dn0PWfeLR63GlLhmkMmqlNy
6QWtab4CRIpBoGRdIfJLjmKqC3fxODEwLY9Gmp3HksthLTuzYdcXGva5x7VPkdQ0TpCGAisDa78M
uSSmyy+Qbx/utnsim1R/GAYBb6yACWgcSwmJqH4IzoppZ6fhDJpQaO9DXPfx3qGb59onDy8L8EPB
6Qq3queVXaNxX6uUjD3dlv2hCmH0qneX8P7K8xAw2lIpoesOt6UO8NPaVgbwCoAX8UkU6HMLg2Yo
8xJOedoL8PS0dc/9EAQovfVTGMNJwQzPpIWM50xKchd2r+nSWgZVcZUpiNH84TnUspxkBSiQvldq
d9GqRWEETHcFxhT4V4A/vm3ZaszMVro2jiVJR7l12IZkoFTyjulhGJK1StYjZqGGOJ3rJVcIXPqg
pIOwQZ9xl6uIT9bDOL2rThufeL3d47cc5lXdtgdsOt7sAlKt1WLuh2+GhGBP/gPOPUGU4yzAGJMw
xbgfROVprEaWrZcFMNEJuIDpRNa+md52kzTW5JdgYEq4IMG2Jqdcu9v4TH0cyF2SpkUUiXx3T5FY
T3qcRc077cEuM6fpAxMfy/XAMvvcEJn71w7pBsDJwSVPN4hkbHshFzfmT2YbeR39d+u1ERmbr+rM
8R4yKvM0fHMSnaik8KA99WTwbWa1tVu4ElyddMRow8HJ8d4MPigfjiW0mfXreDSJNed9P6pQ4r8e
Xj22tOh8x8Ut9esYk/qe2xLL8Z8UtyXX/y8f9t9fXWRvn1Y2KaSjkS26sXhIeB1pP91DnLHteB0k
LChQ7tr1DIWV5CYPswmZeJ2fXvbcZ1Uc/3P3zKoNWTv+9r13MSxrtm0pjmLjbko1u3uoRjwORzNR
9cEVWvEKg+Ym1HclikMbYhZMKhJIuBkni9d1KEHXq3gfj70H+HS8Z/+8LcvZ0sw/wzEAhcrCRjzF
K9Wvlzx9GyTrHG1bjz8q5cn0pR2JHLXezp2t5PhdaEG41OpK9Ly0apIFAnnMAJz/hIcLQ3NDYCwQ
vvHsv5Dv04mWKjACUe3MiP+Z6j+twSvbsjW2egpsyEGU/egr7tpeRLdbdEUBDf6TBsXJyBgQEBdT
IaenZtWmI/1QehHF/bULIEJtTqYGVbf9dRwJg7ThVmt0LItpwUo09Fl1CeKnfk92CuDhUod7/3uH
Wz5HolAz0DQfHe03nE+0jiUVEq3DYhn/diT4+nlxoIrniWPgYJXlwjDBq9rct0uwi0RuYf9cHjvn
s5OJNNFOIYMkaC1kPgdl5m1u+eCGP575ZGeaIWHtEkyI/eEgkuCi0J+0CdSFihI/fJ0AXGHT2sC3
NGLKuX6bohlpv/uF1sLsmzemXfCsbU0KgKnwOTKraJcVAGchuUtDbeA5aZ78i+e4lEwJKKskvN6g
BmcGR+seiqYwwUbNkCHHVpD/yKn1ZTTXoX4j8PbPN+E8zhBnIJ5AlDIecvl8RnyfJeHMgaM1KM9g
eQVhiLyiFh+opm5v7gLLLHAfN81ek31z2a6KsIqkv5K1HHa32BigdOVMdOyI2XE9yA3z9jREtFoE
8DM/4046tddhqO8b2gJ1f8dHYCdGV5HEN7sjqe4uzg/ISR0QTfpb8uoDsN4bTZ2rrganiy8vgQuA
JFBoOuy2AxKQ6oNjeb/m/06HlFqcOe7q0nYrRHArQobbZF++B09EkXLGTR+iAo8IWhodTbd8qpa4
a8YYSpT5Tq+k/R/O1pewIcE7QidZgoKN8Po0WRFuy2t9LBdwwLIv+JWIPyZPq0e3D9VKrlGu3jbc
IJ0NybmX4YRYtUXYwuCcm7XrZa+JeMUB1rsgJQVlWgguhki05ZsK/R/9n61M0XOiFLwqkQRa6qhQ
qbgSfP6il3nR3b8m5s8N5dakvj+BEgaaw2FXUtPrlf44fuzVPSXOnr8eeDDTbrDdXlYRrurFigNS
8y2s+01kZ7DyCpccpQ3GlKaCShw6xBKUQjbt93J3SBN8MlPe6HCvLcclcj8k+BQ+0Tpgd1DfGnXm
cCI6oyg5V8U5sKaUHAtgDCp2J5u2Zaz3kA3BMuiE1z/5dIjRuBLkB74+hOZ90XZxFTUU6qT58QjO
cfzB+zwvKPJvmARhHmo5f5a6WYhtoKwUYEgyLDCX/fWDPDzQpl02FL/lB+YxI3X87KtyzlnEzVo5
SRFHeAqcDctZUuS0Zrb02JEmGjBvqAiYjYcA60MFX6ZEvDrpD1aaAEIIYwFV6wx7K9fnVHSHHo1O
Djd7oYUoITpnHwCBJRcu5uy4O4/N3END5+4844Otu/lRZePs2gVhOrsZkl1f9lZ0wkJUPgS7knsU
oJxWkizCiMEhksG+S/7TPNzBwd48rX7AIp3Qlznoqkl93id+2fCDAh/VYWS2EyFhdxgfEzGHLuWe
SsdcAZOPLo9nAFEno8SjdCynt3+BjCyK/d5O0WOyCcfunSrwsp+oGkuXViQ8+I2xH4tbVweAbiQ9
hTscU3b+2DUVySVK2qMRE0aWoqOxpuGcsjoR3lR5TKbrH+RuWipeKTHI3Q6H8gtRttmGwLIM4oPi
YIka/Eaz0d13NgTtjt5eFlkLCg48A//AZ2eSqDXnOeE+NQPw/lBcDYXRIRK3NchOkMY7WrlMbLoJ
M2+rTHEf4S+UyLmPK3HzPPWs3nAEy/G4CzgidIuKsjiWTkrAySY9OipVRo4+QBc5MyED0eBKptT6
IUSXlsccrR5IQINFivLEHhHxskGolSRL5pAQnJBZ3Qxyb2G73uFIh8q9QaIDbuKPhEudHFuT3kCR
cnFpv5EKxbdY6yCqajRmcqzQjNVNUygYFmYkB1lzESW3eIHvjI1XQWRmWzN67aT+2IVmu+C1cb1U
YSXmj5ay2INyg3IOWaLyon+0ReIM1b4jZILezkeI9YfMCQ4GuPa16AhjAq97mqhOnYveXVwA/N3P
apwpTZjCk3odBJaiHlu+eVx9w24iWRILrTL+duuokrEmGAXdkmLEGgyZv8GDFs6zZRDNUte6X5FB
N4tGlX9vE+9DI7LqsWO6iyy/sGBU7+8RXGJdYh41AFwhC+G7CIJ/MHUAHGkMjK673D7V+1YHTRvA
Vhgf2+Bc+H2Kur/0NCtLCNpVbCfB9mCEwmgT4aF3wlYG883OLQRzmjOTQMnFFGPCVUzrK4b1hj1y
5Aq23EXeaVmcljuNH+4MoMyduftl2dmuTu3mJF1CnSFHJBxBdTt9DDRjPjSfUJGBIftdRvmbqHdy
7uXv35Ndl93GWOFuludw6AuTFpSRvqh2M8ZV4gi6XYXcbs5e7MSbCrI24S7PwyWM+Zj4uofvxT0r
yljF/DfwsEVL8sLJ/EziMuSoziyVRs3BCkCjh745y34KBnVUFrY7Wo7yCeBNmTtGAJSBs1HHos6s
KwVZKm30Wv6l9cjJCo9pxvYmJgHO/sxXurjuGSEOusV+wRYochn+yK1FzKJ40lO4FDzKmWNRhIvY
+RhJFgkZAh3JH6wfjNSL4mq+ydNopXbUsKPfkIgcF3u4n6bBER4VXZU5WwnRaB5zj9EBvRND2Gj3
WzQ3P2pQkVfPTGyII+F9ZIkYSIpML7bGmmtNE4P+VPaPIVbRXnhzabrxr+BxlJaHB4df070qcTw0
uPBn0qc4mCloVVQIaUGksNm7X0DEolXDsShLhNMKM0rnVPZ0dhuT6CVKMG/9hkO4myMbDANPhdGG
NpWx+GtdA4pzwxJlKW9mC2SBQ08UZzeFFYsCQf/l/7dY/P3DS+XFSYiVZ8mPbP8DihxFJljyx4uC
OTJ6ROtrOtvfWFY08Kcp9/mN6MEpOXcCgWG1c8ji/Davzv2cyk7aI5JTvQQzt2+B14x7pL7ILeFV
ifVCCDRVl47B00y8TRxrTjzt66NEz1YfXufRCcdMdLuw2O/KVQbyeIRb22mVohIwrX1yv4HiIXYS
GFrtzHK3FzbbxTwkHLADn7W6dTYrlmKQpt5ZgEyeTmRF8qQAvguTs3NQp29D/Txs/jWGZnRGz1ia
JsY3sIlhkl9zd1qhgTxl55y8vIumEXzYToRD00e+aCLo9pTCSQh2PUEdkk5KGwJX2rHbHMRKh2b7
0HFzGT0VXwgDhF+6q6DxP4ArdRnLBr+8AfXvPsCXoIbrwKB2qtlk4efZtfJ5THTb2rH8C2187J5F
uCTGJWwgWWvCl2wliMkK6TGYegtHPL8KVkpOYKzs6RhIyd9Dlo8j9zGpVN3/74ggT+leykHON4yj
NlYFBuQE5lgOSMPjFR2E5GbfiN52jZC6AFpW10Om+mxE+iyD0I8+WLDT82U5BZKSr22pDWe7rU87
BOgKp1g2yHo4T8mLAHm+vyf7GK6EUiY1PimeBRV3kOSeANVu1rkoB2SY82DemQkQSd2dbGNMLsxh
fWxVZcm/BRQbNhDWu8SatYUGCScL4scEn2DZK7hON5VKT8XyxDPpPWbMwOFrjg8RSwWiMPn7+Dg7
Vhkc3pZ6qa1dGc5W/UMkrm1oMtnTHmudOv6GYphidISyYWoN5r4dJYfvrthrzVhVErzC50BgeMuD
RkIgGlzQw9rk/sgl40j1hVMDJSHFW1ahIaEAKBLkhWJlXptl9J7/ihVri7ChkzPY4jCTxsS80upM
5MeQpVz+9Rt6RNmuyP83aoagFVD2JOv3cVlj9/EjUzQltc8Wskzxm6nhx9VPekccgsfmBguDAdiI
LsFR1k8FJhkxU9BzYfq0QWwT86jS1nwqHVT1tce0IOtTtxXkOq/JSJLn66FKEUymq1RlFhD/FSQI
/MxLia5YXCiAHESYCQd05IKF5M17DUv+4OO7y8WgOmAbBRm+aUt5oNDZy8NgLYxwQLmYCWJAXFGY
0l/7LvbxU6Onh6ocOkVFkqbxbracMRZXYzB1y2B3caXG6ua3HkrkEVXgDfuqNgq8kYytQgYXo8hv
kthC8Ezg15HPiyRixFr1w8i1tWi/wWJic99SEfiFLwQxxiMG5Gm0DCMoWETOPzYKg/rsStN7s0VT
bel5AM5uylsBHs43wnSBExQN1AttaB5BZrdvOBpPS35ZUzqko8TltXbaBHpCZEaCXa/BQtu7Bcn3
FUQGj2l00uekUXoTZBhkzajbdjTNInT6EJcAJu7RxToY1kNerTtFGwLNq0CalskwWUxur2jrWTIZ
GXFhNfvYloLX1O5GCohhVikRy3rJR4aTtJaYwUe2qK92/j1fj0mJsYc0MyaHscVQMKpDMU3/Gkni
zGVfkFIvRfTKGZolJ4POq/BEx6AsJs29yiBCM1MdLfxdAcb3pizkY2XWS7Uoe9Hz53pc46SehPze
DJD9cSYrP+J3+/G+J5GRYkOvlJr/I5TGmwpgKhybWm2TE4Z+J51Eko/rpLWJBJh/a9Zfr87EUv8W
U70Uk7/M+kKZIA7X2hMykfccx6qjdkgbQrNyqlN5cBelEUhlyg9TxqJjuzwpxVoNJ7aaRWRbDRII
WYeNff7EcFdVlPimEeac8IUdXpkC1s8UEJFDrAzb2FylHfRZ/0FAJortwYNsIXYajoxCNFRkIjA8
V261s6BviyA3WYqZaUCIbGYlRuvO33YFRePjmotnwSM7NdsNXLnCLjfqowyv0Pcp7cmznd2hRRUG
facYtk3LUauKHZWRXvgPVs4tRCMFWnzVQWL1fGSaQR2vK0lhbAa9U+O9X2BZI44FdfpDN6S6wZkr
MYtbIAbh49JlTontJ6zmuXxpfzdN9vfKWkMFuHGDKEbe+WQZrCUGmUPwRV2ipqkApbAVxAmMfv0L
xOGEXvzaLV61ON3v0G/FGE24IUsoBPWLXQ59T6wKtT7QGV5ew0bmgX/5qywIXauw24yHoniMz8Kx
8N9cC2ZbYsfrBYQRMFf4suwJ6KHSXWSEEg0KqnOEeTJyXTS2TjvZjquUcZkQUFf1ogJ/0cVCo70V
lty8sXV+y2KzU3hVeh9UGBr/POXg7H+uLfj4G2N7d9pOd6Ugvzw/tjw6aMVwZ38eno78cwKhamQA
OQaNC/8SBDvOCPokopaF5A6TODLVBiNWaw+OHKJOYLuT3rZ7P51g8aJtU5aHZAr8CQIo+/kjjy79
bST3alCsr4cVp7N8sMF28iMp0b54dFXXUYdaCZQbEBuY/cZpfnhuWCH85Fur8eIiKCHFYgvG6tPj
hEXs5PSA/Py6tP8Ca77DDugOD6R10llpmEPv+XBQ3l+1zBSuXHgydxhn/tmoDNEwOgSpNnTLBc8G
JFfuXbx3XwlKrZ1na8cSAEp31u6frtNUD2FvC1C9HJBdNgiE/lHZUhYuO2+fiVsJd3m6B0VoBDQF
vmlnii4bPUP8wfIK7btHnEQvtoKx95k+whBzhVIxgo85eyYmTXZBt8f7SivPfPgb/1pb+WT6yWo+
NCav/+kg7kcHq1pEs+LJnx4Q2EKLyaJa4LklZ3sbLeyb0u09soo/aW3dxJ/hW8gKZKcopPSa1lz8
5MZnJWewPiDPaSbczTA1D+7gBpJYPT3riJmn9B3BmEsTiHS3P/zGM7VCDfWcuLpV3ZQmcpJo01vC
Lj8NP8VSksZgtNeqG70Jp5/YzDigFdLwfFMvot7SpRVDgB8ejean/mhdp+ysTZVkO1KcvtYUVpsU
TcOJI2zQRwbWDqo98JF4wO1eumXGIn0/+kimOILuUUtw2uUh1kYpxcOvZZKd6SZnYqTaP9v43iF5
qz0i1W8grl4pRrM73E32kd2EnRzM9Ap2dgETNwjZ8ijbSRkthrefWSrCfrCFBawbR1J39zjY2zyo
bDQ0vZuRS7/KcxFz9McnvCM7HB2B9bRUMNF+lq+/Dh4VUT8gf9ohFgDDWaSNRRh2yi5iNT93PZ1k
NS5u0AoPhAZD7ZdeKjyMZfwbLxVnPY+32z3Fgir189hAdPNagrQZqb7V62avyrcLfHUBU6yuG5Mb
DUoMmfUuT6M4cilMswslymsYV69VZZ27wHpgZTL9dv5TJiRZjsUC3480RO0rx7VHEBL3RK6kASq1
wOOl+YKzvx5d5Y0ALJjr1E5FrGdDcDgiPM3vSsnZXmu/WpIcGYRuqE7dfXta8dAlrhmh5dlVtGgE
fw6Oq3arqLLc5fe5qwqB4Fbj/hnW2G0/RQhY2FcQqxvL2fOzxdoOBpcDP4HsDLlj1rbWdnAnxfpc
6VJrGpCvUPMCsE9/b3GM1L6vLtDGW+4gKm1CS05qcjlK9mylKp/FPPUaVmrPXReYlHr0GRvQpG7f
kX46bXZfWmQc7+aZ28J8hOVEMvLVbz3CYXZ9CzvO6YU+sFBSQcglt+Q0uiS/xzE+PbYRuvEs/hIB
Td2ledaOsZhWpxNTi1ZlYk44qw6fm/+vglCOj29MrM+VYhW5Wy+B9HCEqgvTHv8iwh6afCXtieY3
c/d9eBHneg465rQKIla45YPfhi5iu0mOoWJBYc/hHDOi9Q07Jb3w6/q17KnV/IyXvA2JokIt0CBd
G5yt4rR+Tv8gGtyPlXP3lXcfZ/9SlwyDRRc6O6D4Iq/ZU1HtrvprgaxzEviSUl/wwlXGHqAJ9bww
g3PggrZ4My8vDTGotY2C53pElKraY3aEj7I1w8y7lU7m2piTHQOoVu8Gqu/62tOpd7AwhezpF4vL
34N7INZGhzeYoD9z0YSkaMzKgRLcVDyQ9NvX+rxpymuUnTA51z/c62HxFYMyqyABflBBn86S8Lnh
UYOmNMwQJ2dP8hf6UxQUJ51xLyALY8wjyr89g0dupx+sR9J5KUTLTZDrgU/Mh16jLPBmhXkZ9rPU
KBK7nKBHhcav6AXEVT9IdllJTIDDJLBer/EJWrEA4ZRf0z39fwsNb7SHnONjDGsP0XwRKIYaH2YY
HHxB3pKFEqGYXVcJUngIR6+j501YemK9Oao/kFpmOuzcnT26PUlk6cWJ/JMUSKZJyk+l2rrfC1Hn
WgQY+BSY2N+5S0MbfR/z+AQ/lcMHwdCih61n+DXbg4vwRDBq5NXTZWDRPVtVNtX/qSOhewjp7hT/
X/xVaSDV62oL4lRKAkFxG24chdK7tHKaanppLkJzeuATyiomZOY1+uC8AGei199l8IAkDA2ZCa2+
6njq64rtsTg02PRZhi2KXQ+dqflD4tuzHEmhE5t6geR2Wb5pk21P7ejtuCN4jg+XgpSGoKAp7GAl
kobaqlu0nxad8pFNPoGMzNMV8DH5xiTDw+SBtP8kSKeHlysNG4qlhehQfawKLbY+6qy2mEq7YL17
C1y5f9rntckiuO6OLztelYTHW5JsU3jxEb+mjaIEPMAqgWSOFj8Dj/ZFxlWZLFb/nwBkOc2gfKpP
iLnJ0t6UNx5E9iOZMK+5htVneVWLl6xKT45/e1KWtpOM06SZD4hFCc5xQW+1pweqioCWi9qZVj10
GgShbKLcXgzxdhOqC+YLOufNMGibLukiN0jB2lxCST/tcXxYsaT0Wo29aEcov+EdFXH10nyEkPOf
VfG7UJfnYbXbM6N6KWSooK5TH95m0ziuYaXUh5QdBKlLRXGls1FALS5HnDeVQbKTibzgN/Wdw5dV
mne5jOvU0fL4qfXeIyYKNKJMxEoRks0xiV62OMzPH9NtSrTxi2R3JNAgIecM+OvosCe0CwYkQfVM
nEPdJ+Mzv+Un+FyBwp+4LkWauR32oQlAwJe9oBUkDePapx/mor9+4oHl0PLx3elK/vsGt6fLCJCR
kIyxB7PXT/LzZIGubb9UdLJiD7u661g8f5PlktUEHX5uc3Lpwza1Y8rfC6bbwssHKdLtaWWWjLEH
vSxVqg8CqNsSLB0+RZZI1xoTfQSg67u/F4Ln31sMXlXR0o3k8CniIuauO8hAROQBjzGi7Sg9M3tJ
CeP85/xqRAwPGxuMkahvlfBAZZS7AaULvK6C00RYC47S2w9XJQGPAIta/jowLhixtRDyOoxuDEUg
JROdK2l84H9aAe3IZMzS5obGwOU0ZTKwMjWJjyXbqKHDky8NOFFb7k6UvGbKYobY88p3NoRM36fl
e3MX9Y+SWPxPU8WINh/GIuLabNSna6EnDNyWfWTApLcIA8vbJ9ynkf+Aq8/we7+swUiCUQHe2RDO
83PYS+2hSX0hRKX8Dps41RXVxzU+ZtPHgIRelCvySyP6xTbYfpzg9+ZQIYS8zE12NAggH5pTjscD
nGRESjPvDEq1rt12Z8OTrGn5wdvsHztZ5Ed/ZH73TbQn30bpQzeCRReV/EKQvSHonTvlEDN8+TZd
UeWjiLab5Ov59D0SiygjRaMiaILxwXzGRBWYOvaKyuJRBLsB44gCig3pEQ5t0K/p4W7gp3zX/7Cs
tYXPnmyZch7CGUTcIzH1MrKTCWtnNSLfF6szq/Rbzg0+xg0sg6JWU3gc62R6PA2BbX5dC46ug6xB
H3SQNzBpXe2mW/rPgmXEgosXERl43IIBddtYIY/eTZ2DpTlJQrBO/SNO4BTJ8dtw0KYg39G+iYXG
dpZ4R/BTG8jyCUh6LIKqXkF14U+p3qTwgyaS2YJsIeidxLmbqIPojXTn3uwQPON5OoYxq6p7UFc6
Eo3OAabxc7mxiU+W6TWrGQi9aypZRspB6GAmbNgfgjZbtR72gBPYVeY6zQvHIDmTRefBwZQZciEo
Av4H9X1lqL41PW/tif5dJOSKNdLFvi1pRGC7IzYqXY5ndId7W76zWttkMYnAc5r+dy20NGFpUSyN
DdPWFCO5PUPdJA1g0Am/g8b0EMpd4hhVo2lvyk5MM2CR9/Q12NCj6r+xdEIZOb/F5TD3Z3aKjtm2
TjfaqppNFuGPJQjPUaDw+VWnj/a2oafQsPMcoJnW/DwFV2FiiZUvQeh2ma8IlOVoB0T+rN+jXDje
WOkFU5SlXVnl3R7X4HqA1iN9LEN8yVZ68/er9E0K2E0uZZkFIVeQ5iIbB1E5FYEWP9GoRO+hUPWW
knFAMKMfVUfhPMqsy5ge/sIPpnZJYXGIk1BWDK752+rgM0goAeQjMQcXmnafoSKhX/QU0BOU8og0
7F2krdGBKMSbYXMdUoQ9YLOx3z7ILDE+g+98RiC/QWmTQ6H7JuqrSziDrA6nOvEpp5Sj0WFHT6n8
2NrgxW9c3XJql/tsbs2hAaeMANccry+TbJFkAZbICUoYCwyBfHDsFNioFAdJfIslPLX8Aq7I59oJ
9qacw6Yww+iIq2Qo+8IPGyS4NGqWUu7GHI0jN0QrdHvWhC6isUHOpHd7e8VLxu1bOecBc39lD0zU
wiMQq7WTKC1A2bdzDwMt46fem2gQQW68xEuDrrSCy3hvhr0xn5W1qLdg2Bqb1BFVerSsTZnJNxoa
929IuVpOrXQxpcvAJBIEw1bFfgf9wNR/dwOfUkOT+iUC/dLyHz4gpRAL+zeXS6vbbNDaD+255aZP
MzDbuP0jvUgVlKpizHUX3PNdPiW3I3Q6fpIMwUIOUBqM3pck5gWNlZjAQSOP3oIsFCGvuj7cEpkQ
mRztcrzDIGebuf69cXy4sGrnqeRZytdmYreFUd9d2FocKrvYBreEjSWem7OOiH33tx6ET0RMYIiV
Ojdu56vINMvnp0fBdPoSewTG2cLbULHQZFkKrN+KHabek+QgTyMYxXcw4gldlUd6vMyy2hJP+uYa
Z3/kh8Io3Y5ft0LOH+/RT9wRWkRC9Ki71OS4P8JVQLXuvzRJFgAjbMPZFb6P7kmz6w4tMrVThElj
gUWIKmDvtSvGaQfx+MClnBeTaSiQoTLndzhMN37/IkhL/s6SJK9yQmyDMVYDbZPOVql7lI3DIooa
4axqwvMkmUK4qi7MTz97xo9mD+CLb5Cqi2k7kMTFACJPHFTHbhcXh/X83XUjH14FOAj8OY15q98q
7GbAH4XKS/TsPsRJQqx9TE0NJd4iPFL5PUjXACecNBrs6psj7kHbmtchGGN0o5FFEXjtcnK6vivA
DYbYwm3Y3S0/46l7dCSoIfPtclrJ+U34H/yZt55L0/xdoBM+UJnuEPpZT9DJQggwfApDDYs2TmHe
GtQWb0j+n0iLKHrikziKNaix2l/XWamX1S0iSv3KTmbEWt87tdeifluA/pqYw1e9th73jwlDhrVX
gUWmRWXCEDefdnXPA45cJZF3kf4FtpOOZ87xCLfosue30gqet3mJTnoVh1lOxNWDE36ikqT5SQF5
m57UA/bcq5MDNYDMO3Xam4CLNkTK+PKWhKd6zWswL/QEh6e+gxY9/LRyMwsdC0YHxJtQM8fpcIi2
4xc14nKqaheZyh6vCwTz1BsE7nxZ9PK3sZ2v4RqIQx7XBSh5tZ5tLlLD8P+1A3elrYN0to5sZ1lZ
Q1sYCKz0KM2I9axCaBu2i7md5wmJcDH9YSIR/2qN97JPVr/O5klG2jDQBcYXCmRXLS8aq7qUXpsU
k5rVP/c+6HwdGoEgeaP7y/DdPVKXbfxDEi5ifRwQFsf6LoNLWmYUMivz9AXT74f9DoQ9Yrt/7608
B2lGtQIL4Q57BxSQxrN2bZXTMLEn9Qex5ZHmUm3o1A6ZR6rlvdpfYCtfmEg0/8sOFcN1590RvWR1
Xvw4Q1TTDp/stx/14oq+OPIOVPO/pJYdu3qKK5vqaxXiYBXIqytSNJLs+ul9Pa4qLRV7RAM8q2cF
Epg/OuNrNCItfakGqVVswI1b9KcJMJXjeAnKVY1Qimxdh+eIWYl3Ejd2IDzwQCdDSzKVTtIoZOtr
TsvFmQ41l9bS5qUkECmBGD+NL+2+3jT2d9NQDDD90ONDtp5Ch9jQMIw2U9re1iBSx7ELJaeMIccb
BUn8/5M/JK9SvI+0Fwu9vovJWjDKsuzhR0cL0Xd+Eu2B3F4zvqhtYLaHoIRoxor1kz/hdTr7FTJU
jszPMl76JE5gB6ZgSqFgc4TYCsKxCH0R9/FmtXePPYcyIgu3Z3kR7re+yatbye7jovx0qOvDHElb
h7cpEA8AZosGZYocGKteewAULdiWpo36ImjK0Z/bmOOUaPeSdpCBNyPXecIAl3cglkdWyPBMzsrN
huUyTSRmFtO5APV5IMyKqj+GO1HRiZYHd6/Nqspr0RYtfBJdJat9hIYKv/ypKZm7Jxup1Zy+KvfQ
7NsZTAu6EMCQfOS699S9s3l/V6JnXujTIxjdGuVMaKnKTsUhDOXW8jqtTU1GkJ/rrVRg0acV+m7K
RHkSvoDVi+yZLuvZD+tvDdKDKzVQtdsfdvHDVBQwqd+VKianWuuUzZqwBDehr/e2MvLjV9YYaW8Z
Vh7WXiamA5/OYsKzGIP7b8TLcKStW14JR40GXxpeQVEffMPHsJnVzSzn/unrU9cPUzo7PKGvsqoP
6otZz0i/zcXMMVjpkX7ShpvoclPPKQ8zu1zcNgX7xKWi+oYYiaZInL0IF4D0Hft3pUa3lys/R+Uf
s6EruMcoiTKI4M0cCeYNKEk6h4OhqzApDB5L0NITZD1AwyjAAZJxcK0Uo3Nlj15zybbDCeGvsEIk
dvNjJO4j1ANcoXaoGGxhmoy4gfNuqzX3GY0HnSCiGR3OVg0KBye41wO7+WrYGyXsYpLeaHr/0SYM
33OYBENst1pYIaAVpmGtB27LE5tOsYlBwL4CipgIjp8k/6jflOiYHG5xG9WaWNPEVDpa4biSdxZm
9mlcIjY+oxGvAtUKvGBGSlHJX/qUYo3MnYaMNIiQNk9C4nrTRkb+0W7prDNICzz0guYXY/m6yfbp
RQKiKNxaxWylzwUsmqcOk/aO4hRd/9IwHxJk6C8mE5yzkP+tijU50cqNz4C0AnWg5wz3pNJqJ3Lw
qlup/QlJh/JWC3BYsiALRLntWQE+kYrcWoTZTvaZIh76FaaAW4atlHWEEdMzR8NzHd2ubymj+Vve
uIFv3WHhJrcO1YHmZWbDjX5GrAtrvScXLKCpAvRPllY4J1sy/SQNE/9kLjt4/4Byxu96AEt9MUGW
380rI7eYNNzOWQvM3YchjLbYjZhlqLYphQV4tVXfkrbagsu5AH0LCShBuW4IdehV/COig3M01VL7
rQflDrTF3PhTR2rY0VM2Qb9QQc8OmHz8YLr5c1GZFtfdsasmKGciOJeSndZILuqMG3hT9ZIEUlwn
P7MdxVZIyl80D6snv4EJDipHCP5VrzyMSCPJvn+9ZXtlmm6idDkuifsM3rCCZAkOKFkEz63G1LUX
930FKGmHtIVGzIJ2j3IHQNidwsk8CTkTmhQw4XEJ8dIZD3fVMpF82vunwQ9el+Z1p+L6W7VN7Twk
Pm1U4TWy0q4Av7mG1j6Ni7+NYFib7S/1xiZEWupEtJa9YAVZNemJswvysG948kEhahJ7
`protect end_protected
