-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xJCivILhvFrQZ68FYF0WI9TGfnFEXvm8IE+EyOYwcYtx3ROAFKWP0MCbVQk/ONVlJNbwd+zFvwFk
8S85g5LW/ojbxGbjb1I1cXlhp3AqgxHYR7AFMhrshHXVu53az5vlhbULI9ACDJm7XLDlpQEpdDht
BjVgWNbzbk49r2o1dRQTJcGsA/rg3NHwutrWbSHd4FnNF4ceL8HMZbLEGEtXREQ/kc5z7pMwU8ou
ZSsZi2QRDRoVw9YG7nH96BrInV+RzhZNzImuf7BAr9V2zS3/TiHOUDBcj8JXEpugikbNdsZD7L2E
MN/ejfYPRTuGgTlvHt1M8F6L3b2n5sxzqsdIqA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 111968)
`protect data_block
VpWnYYe2gv3B0fykrshj8YQ8ELClrM2PY+pkLMNSUrCXqkD3j2fcUhn/oRBzisjwagYFLB4n1Hal
mLpdt8g+jg9QFWGO+B9lsYkQJA31d1vDitnUyT+eM07s25X+s02iRwarlLyWFprcvDOivorOPLOO
TnNMu2EoO1xpcvinKnlIbfFaCGEk7GrwRHAlJOalgPqZR0UaJzKZPF7NO25i+VJHGV9Odm1K9Qip
5vdK7f3AGBoobJKzdMhDV5um4Ow1Fd6ROrv9bKPtdVOL7aEvYsOVWVX7xIFSYV09eJ+H10l+dJ+e
UatOfoUhtfabVYepH3tiyelfjANeAeayMFZtB0TmG9Cmljj6qCS7mqEL0q9PjnMIuwSqswbU6QG7
TkpQ+d+ArVU8LZP06DRzWEmijTWTRRkgPOEYaseNZG1in+ZmwjqklDPTwki3JaJ2AreftL0m4Sat
oUH5c7Od93OTORvqXZQN+a4Ee8TBfpH7fqOWrBMaxL7dgo9Vs3ab3MRsamMtIAIpm7JkSuDRRZ1/
oDA0+p77pAElvtsgyoWFKq+tI4AqfbDFZ2pkQo3J6jLKXZcilwzZ0lAfU1k+POniHO3XN1TXZRgE
L6LMYM4NzZMNDtUFQeTw+epRxtFQfNheQJ2Fh33UY5UDy3NcyJqlg4CIdKmx5GFXJpYVHiakphPT
5X7DFBm7209XJKjL+xCpvMX3SNfFyS/QGwj1ucpWMRasBKhAhA8G9O5zbGruzmup6APSvYUJdY6/
OAVzpPhN8dMqSPzowwb+xaIU2HjQjK28PjXle/jWxaResmzJzZcU8hQG18SROBSNjFrvXQfQ9luD
nMxMlUmRSh1WDx9r05cjflSaYJz9MdrymYgdlbyiG++2XcCrMuo+S3ZD/DqsQeDG2/Kr20hzC6KA
wcwq+z2s3Zy1V8VYljMdtlGJmNbXttyDeNHxei6uINMo6gXx/WOhcHVi2Pwy5J5sMcLPLmE/im4y
BubJqsoyzfYxiWZk6WgKA/cq3Dz9flA89OGg1kmqVmscgm0sM5l/n+/RicZRuzwKNc3iXo5V1ZWP
mM0u5QgO8GAqWUwrG5y+rbRiWtIFhTsNwJs8sO79am4zDd/YrXmxXVDQ1tpTqZ3uXJ9WQ9QDGddK
rdvRIqvQO1TNQaMf4PTi8G3tuOen6DgubBYozucy2BuyTMWhEOrtmh/y1ezSk41U6miQrw9thq77
xxSs4UUPh0gS+v56EQKhVsMbHiEOyT+K/r/m7oR9YQtf038y3aa9X4NChm8gaIMWNEx79gXMQGGC
jsOEWIMtO0BrgTlYKB0ih0BtK293cGjbsM7N3cbJRBr8tYBAM2kqXd7VDADtujC07rKrD+hEce2a
iZYmXCGQSAmtbLEuMedgwsPHtYwTLwpwdun+z59jBvmwAiThy5uzJibx1MvJrstBQztCKVgM+Ry0
wBgiUfBH2jL+GwsSSz1ir6DlRto0KvHtk3eOUQaEd2E4gnz5/470iC6U85d/iOxOxt1mLql7XQQa
LY7dJOAGi96V+vCqfVFkrazKk5PYJC4vDuVyMZVLO8QBUc5JMhEVLg40OXkT37pYo4DPW2C94Eu/
mrXWX+ZZpyS3uIEKVEIDjTt3Pgm5pbtNaXMDaz+afOQ0k5xsEb2cYLRbUQNFYvIGDTBSeEjV6PU5
LXBSXVTMSZXLlvJu40Rx9f8E9J67mM71lnaRPdJGvVHx7GBq1vL1Irkk7nbysfTEqItBK09saN0z
3q3NONjkiW6h+K6b4czVswX31W/jqoo3UiJmTyOdsHoD6iDyjkH6vwTpgIJ/ZmRQmvDCE/2ELBTn
s5SrY5dG4Jy8qWNLnT39okZO89RmSDv5+wexndrknhDkXgz1GTIiPKuyaAkAXoddCgtejVd1gfBR
3xeNTa5x9x5F2HfzMG+PLADauFaVZqf8dauRVHkU262yigyCTyDRjcbKoURJfTk1OrdAoL7Z0QgM
8vj+xPJ/kRWSM5ni/fcrFBVItfB2TH76wTgEFFgr8n9s4rCcypnZVoTdpp+uElRCm8sTDzmUZjTi
qgk+wNkTY3qm7X/MbChlvzKS6lYIfWiQVVyPWWBjFzkjQh+UmDZ44Hpl4UwtQa1678iT91XVQAlc
D/Kmaj5NReXtJbOudphb2jak9hhZNltlMPP+ERXJoYHRPeQA1fJOj3sJI9L7WsNTjKWzzMQTsnmy
A972PVKZKB4uzDBVg4QKlEIlatY2HQfB3g4zbZMIaVa23kEObkGuNXHwsWuaZbp21nJQbUE5ZIHj
go/5svAKtbN4MVO9GDTV/ynRu2b2o3oRP0EeYPWLt3Cga6DToIXokml1O795sc69A/QtlZiIpWB6
lb95UxjPNjaZZifqk7YvisJuPFoO9F+g8QRhc0qyB4FSObTFDmj5RWNUR34AgB3e5cdfC+1VmMMd
opVgkZcGkNO5WEFeN0MiSu9SDO9uj7C2DqW2WqwJ9EspbbFhB82+yiVxXCGenm2ZZlulIXdoE1L8
3Qz2KjAORmS4KH3FoGzTVZpdxsfyr9GXE7PTO2xxg0UFBP5MI4MMOt0vZ3TyT1hGZQZtRIA2ijeD
8vqCmJ0LlGUGXYKrRqSM/COc5CPDeyLyJsidQQ3w9cf4POsKpHJ6TK0722K4i0ieTVdJy4jvKl0o
ZEa1Ti+z2KyxQUaqIl7OvsEOTWK/5yJ44XXRw8PYX7KG1M9rtBeacNQwxv46UKcWYtbw0QlGyOR0
3D0kR4K4rX6iWMW3wxBLPJFtdvfp2nLRF2qmWyD6EpLvNwTzvndX7KDniYbP1uAPxA/IbBLrVH1o
q1qLShTlb5yi40jHoB5cXIVTB/PEM2p+rj6TiUeyyGIwt4HjHu2mBZsQEwBSZrOPuyO4cFrQWszZ
m/ju3oGwG2mB8/tZ7pV2KWIJ4rnEDt8E1GArwl4XRPO0SPmRG3/KFZL+tVB2FFJD4ddEoVw/FxyJ
MzPKzmsO1tnqbH5xIca6pLL1EEkHiPpSCCnw4ipk+S1zw0wIZ4dcQmIUxv81RvZ619HL1XKSUJwc
Oz1HB07YyIoxiF3eRANWpB/WNGs4q4O3RvkwhPPzjUfO8aVM2TgUKoCiPhFvQWZ3GDh4oFKj1ROz
dVbtAYE6jqMoh9YZuXbOWUmUTi6htFSPMzskwp0DAfSyEh8OiBPMt+EfxkINNocRX7Nxv25BsSQu
Kgmd54BXwFla0M68D6pt2tKtgIzSAoO8jBrlhsKvcZ2EfoyTObL7sU8zFTZ6X9UJg42cVe+/TPBa
EmNfGgX+maBUFs4yP4SAONyptdzOPHJN193SDK2PhJelGGabzeBL2QPSUJIeL2iKqBRZtp6ALjYW
atw7UvYbyus4YbDM/dbxre1FCUJw+sv/nYuD4S5SLDRs5UPHdodwWAF1xEIl7w+lBsohV1JIzp4V
ngzOghPi2kv9s5QBeBF/c040A5/U3xiSEOgndP/mw5+8AtaTYKSWzGL9lIhI4MUKUj7T+3zfIWtJ
QjzQFhKUjrGM8E/rsYyZ6sGpfDuDpOsjYCNX1qitcymBveZqqG6qukUIwcVdsxO+t6PqO8mD6d2x
wFwnOPkJaH9rvZ8L6fmj2PmA0m/LTPSOs02tt2I0qBcBf3BcTXUsUazb5kBXbk9gXMhq3AZ7rVg1
KtTkFmKceX2Vo9chsTup+tM8vbU9jb8Y3rFfgSkZB5DKZY3gvOkvWMwrtsnadkFxkwsqagFVPjC5
iWSgamZJEic0bn/4d3vyLI38Gu6kUpjlVpGIM770ozUeRvJt7peWoQXAmu47Fcvb627b7F17l4Xr
UvHUPyLgWYOGWXG2sK8UhvUbVPJiVYYuBfxalXrcfVdcglAmkmogvafVZzK4V7QuhgH7xcg2KObs
/2bmOCzc8g/XZrU8lFtxYX0DrnI2lEThQlnX4L1QfbxVtDsiJA6KNE7TR4/TNfVPD9EHt/alXkNz
6/aEOo7vjJOdOzU6vjTwR1OXD0p7kZgNOa+xaNKMfKGkj8fS88elTQpib1ItgD/39GXaG0DxCh4O
9E9HPm5DPdXMa9+N2WJIjhZ28rAgJqedR5bYWzQxg/S5rC8rXfeaG+NIX3hNqmu9FQzItPZ2CvD8
k421WOTUmV85kgnPmnEKyalVxjm2gwBRIFkNXBCK6Y1qJpMoavK09m4JdTmKqJw3D7wO0atm1SVH
N195nmF2RrmdfWfShbF/rSO7Qh9FmYWcYMmYW8tcbFA5IAQ0smzW47XVriCc4fHPod4WvnGB7Zli
Pxh3aqj2J+PjK+J6C0K4Bvt2cG1c7hlQZcEU1ExgoSLnbYdeUI7BI/4teL9w5S+07JnNdyJkRN9O
CSXGnXG8UxQ9/hYS/so4eEBPffvgls4kp2cg1Y7xJ1Yk9IRrIuZK2J5WD/fhzPsqcgyVd4gi5DpI
xnzyw/KJvspxjEek8pX0sa5jK85kHG9QwCYZMuGrdGWtObhjL8kBkT/ZApUUetXrRZ8wPu46V7zI
dbXHMeusRTMvmZty9aLoJyLZ2OCMt/dbWncLBcrYb/Ja7wl4t7ZVb3fK9EZa6+/KlRTnEYx7Ze9e
k9SSo4IGXqmY+Sis03Q4HfB0vTKsW3mQj6Rn1kr4RkzZauEw6xPFC8lvdYu30DNZ0wxM1M36eyFA
sWlufnb3adhxhZN4x9BnGVOivhc5GYMeQlK8nd6gOUTbi6t1+QSktK9CYrI8HrsEX/hq5z8u1Jgz
KTro87zSIR+ygp39pUe/+iZjSOSxpHpTap5wbisgbOVylkWdgav0EOLOjD5XizEYHoOoYHFL8p6/
2ud+UarMR2mOIOxVCS3OY6st9HQL7ucbOt2z8Y0fX+CqGSQXfRQ552fJ8fHKlHRricvXUvZo9BvE
pwUpC32i2F1oNe2mLrGTyGZzMrUDcflpcNT3QqZ8E1oDYzAOCBdtaD5izg1g587SmSELA8rzWd8H
tDiL2mC+95qLIxRNE2pvPessggvSZZ3xLLpQKRFJQvNLdALFwSuVbVGsOsRST8RhdcEtvmPwb5/T
/G8B9DimO2EqIiO+24eZlUCbBon+5JCL1wiNd+hfi2UbUGqsAvAc24BIT4g6/kkuDBvObJvc0GOX
WhB5F6L94RR/XwgizF5z20wVSEOSbbQaMiI82gc9Jg4cgFrQIEDW8rb5En2f+kE8OcufmN1BEu1n
oVG8A7yudvhER2vcPUrzx6gwm+5qThPgNCZR9TpT0HGFLQlGZxQRhduVvnyLB87xLKJWfsGgrVbv
GyMeZs3OGAE8msPEXidlwHro64USSPgkG058iWrHgKdBd8MCvEaQhjYFG+Gily7/IaRjx2AgLtAm
HDJ1bjS5Gx+YSM54pDlzVRQWZIkVIzipC/R1NbC2ng/nDfbPXFgHRLx4MxFU540Cpr8WV5XIfnNL
9rRYMKTbdH9VQM6lR9LU+ly+cKrhWdAyQdK3gWlL3HbvpKdAVumCQb2V68XRo23E3XTt3Q49xCZn
71EytfIKULtoCSa1JJV4TwPaoz7yeXHvaICv+9xvpp8RGHsSQjQR7cltABLjZDThqPs6AvBf0MHD
gszg1Rzgv/KfrfWwGpeMGn/0m4FHZhgzN23SCNmNTcwL19JMt99hsaUZQw+BNAQebnOBwFn8XtQD
bB2DJmnwmB4G/K4+bniHcvy6BLzXuGSx9cj9Z7A4Rb18OZU/P8t5xN+ita3rSaBaHgo8oFmFHrMS
Si5JXeCc+FilMOI1NaHAHsqkcJsHyMGUWaX/l5HhOChJY+9LhNk+DxY4nrBF/RztjdT8ewCdXOzi
KFBU/jYzdwgiartayox62/Ll0aeVOWD0cad6vcbYaJL3bfJtM3/OSJiGNDnP/cRrNcUcsl6c/Rj0
voAIsmrgsKKzE7HN0TlMg+Sun18rh+rG3r4lAR5xzkvUIofxsryDQ+ZxbbxkMjA+Yj2PNY5djzGn
p6gWhS/m56yq2zNFCzl2/mbZOXY14wxN1iEGfXtanAF7S82D5QSDrDXqhLBJHnKMkZCzreulWCGk
z5FxPzhQ4rqmMNp4pYggSZtqImT8L3zgopPztzEnW2ovSxs+EXln+s5yuWN94FdnQXC4csD8M22P
au0Kf9IOIp0os5vDa5GrYRBZO/+Fze7illahqxdMZT9ZmsYhwAoXL+U6VLD+n/+N4onvtD3iTfqC
mnXXr5kXYnB8CfJ4AGIndZb79Zu60MGtngdGjQ6B1dWaF/1JH94/33u/m4V+ls4pAKiYKpe1C7ou
fPKBW9pwb2r8BfVCUaF8KpM+pIbl5tgK2SQuZwSiQajmeLdUTF0f5NssQs8upTDLc0Btk1BKxyRh
mDCqaLCRqYva+ofGNmd/Bx35hgImBxIUtroQNIIMvBPJMf8sYcYprevv+Fewj5oqU4DLy6/20lHn
0EOmpBHCnvDY1zGJai4HupoahySJNPwYyht4/P4TdDvZsJ+tX3uiCgB836s1IdwC1rw72U1FXKdR
B70p9poToujpwpo+KQzMKdbGYfqBSp5muNVv3YBZiIH9hbtAZ08Phn52QC4VakjFO74VBvZVo8B6
SGRLGfwPvFITrVbh5kw33hw16RJ5o/qKDvitarAZImP8Vlix+1c6aFMYb8s0n3wkJzac5RVLo6A2
xggyPEIaLWIZn1TsdpRPjSGFYGIXNUjN2sWen9a8BFoFsjU30PJwaHU7lnBSRdCpWaJ5tZQQHqlW
T0xu6UQAqXWxMsz2d3lnpfD0pDMPqOXHo1l6myMIEXyDwOkRzSOrYBgzrJTB/SOHLaypFRIYCcUa
q0TwL+Y46iGuGorwGaNLK/U7/HkuuPAGgYrNBQkMh+ngfRH/3pk3HVbU7H3MqEKzUePSDIQcYWdW
fC5wEx5aXTJYntHMoUeBFaBUOOqU9yWKmyuQuZXcIue32N4+PaSvXyH9SK5DQE0XsiQdveGq/vH+
7J+zeZ6El5sbp4DnDZlJ4qbDmewJ4qk4tJQhFU8Z7Tlg1jbDWlLXA0LBzK31TF0AUDqeud6xjpSI
dXW1atovP7/Dr4Qi0GDB5kmBolIKZPECv+fbAo+CKUmeB7MtZqL2KvrOK1hMTvk1+4Qbbk9Aq2Eb
ldBENtwNelyQLLo9wcUNzWwkjf8Lse6YaXjhKcIslYosejoh0WotEFNWi+G46aPx3IKCROJ/PsDX
U41uYFppmt6dVnkE1Ng3DCnThVEOor+QAqkK2YYiJ9XexfG9ZCwLpUlSLpsjG/lEYwjtjfYjf0HV
cwfcSZD5zoQXzHr+trP95q7Y4CH1zX7THCL1E7vSy4M2hB8rES0iBtlW4UCMwOORuXI5wu6iGrZY
P2t3WNHzh00zJXrPguCNiaP67OtagdVQEap3sUh5P7rXEXdwEQkQhzWjOyXN2vbKpnRLY8NFjSMS
UmrCFw3nGFyGUA4gm0XuCKYgQ/L8mN0cwWAC3h6tswL8xhhaBcEiQ+XGgJZ4TMmp4l9hC7LimlUS
EPrE9g+LsuOjoTf9j8J//Tjtm8U6eCqiEr8KbPeJYE5WnHNExH5FbXxQ/lV8YT4edNK0/lz03UMB
WYpqh4AQLFp2qw09qDSniawVO/69SuEICGGEEPcgqoJ8krGFMhdaNwg83H+83MZiN/hOo7yvB43S
qGWbDaLyeh6ym44Inc+QvHYAHD+W3S/89y2yPrHoYg1GAliCu4WzpRI2nwr6PPGl7ZNnv5WSNJR+
Yr8ZadrOzTF1I30sRbV648cmcunatAK8pA3sqOWb7BzMfkOvlw1fKFRqC7yV+mIpWr/rn5cQuYl5
f7N6Lxf9vtz0aOdNhQl9w7DD4tbcTY1frhhAzgP/6xW4fJe4T8XuKN8eOI9OkR2MiIbIgFtYvZxb
X1qRySr8RggFYT7vIkXqulHi5nW3h9RwzwgB8RbqAhpTSH+jId/v4mZt8Ep0E5UAJUslvsIXCLcY
AXZ2rczIXOIu06NcSjpJJRpW/SbeVBJ3fY2zNlH7wLX9aXfOdKVbnJbTkR9p7w8nSuegVkkvB0NR
g22lxiakUHGmGTLZASjbe4awf+ItLcdjrl4BzWE8N/cQ56ZRSAYuxloJqeAXAR+soHO4e/2XE33+
BJ56OGN6urRryic7x6VoDxmlN1kItz0U0yR9jFpMd1OXTpvoakAlTksHxPrrBpwrRnJPknEEJeMv
LjV9tMEMzPug+U/WXM0LPx/NTNiftvyjYl7utbQ4CGkw+jQJJ3MqNFUsc+kHvthxS+J4GQiXJ8u2
O76Yv0SVgyhquIA62keQPe0YHdwCxwtE/rNVjIMJruK7C3lEnAK7dnMbL+jb5cxiK9e2qjXg+bYU
wW4FGi2lNZkMKNVjbE5rjTCW7obA5y1tkW8vKg9qraxAQaiXAzJjW5j0q+dO7aBLWFjP15TKzHoS
5qnweTAPvc2KJGiwj2AANNbVWcYEjnIsGIjGrAXPAIjAzMVx584xiGt/I7LsCbyjlh70WoS4uH4U
3Bquns8izeBRzwZZHEiHMIdBKZpdvQE6ZkudMMK8tl3K2NQ6Jmm8Nt7sMM45190a8S5z7dsTY7f2
pFsIwGsxFGC4Arj8v8BtXaALjya6uN62xnH8HDYZoxWIzJagr/vVTuuRrr01O5cUiR1iP3wwWRaQ
TvHZjkER8Rz+nq3YynbZoD2BSCj6lekWaDL3nfegeAPlYjUOiSMamILPBZAgIw5dDGsRB+s8utfL
G+FL+XDIvxcDnzE582uP50TLWkt7q1eDtx57dn7+93qRJYS76alWizXRWYxvcbnMegTHPvu2mQCq
mp8IhPMjhxAxowip1FTKWGoAOCOV2xGlaB5CtjjQFccb45n2XwDQWiJrFR20e+5lzWzEYZ0VA5id
rV9DbIfUyyFlBwJjmxAmcHk6IP/LwlS4SkaytvFK+hJKcM8d25L0/UKn+cLNh+M8dX5TGfD/f5pi
pO5XfqWTTbZVAi6kPlDgo+6lH6uw2bR7HSM1oY/saYrBr+Z6KjodQhEXAllo1WdH3HgT39YBVkGt
l2d2g6xjSjWFIgRdCttF9D/RgIUUBBm+h6Flb/8BvEAxqdSkW6ETwqub1kCbVBuzypt4II4tOp37
MWTLrIlfqa0PNFSuSar2Wa3GSOjrodZSuZRoedn5YBGikf89wBOxvR1niEyHYwBev4jsJjDYjUGN
rgBDYPh/TVyGDSCKonzMHxxisYEPOiH5VeWYB72TZ61GWoHv0gTvwZzhCiPHMieQ80ZGT8yrzh8e
R0dzwDB40evetd2Gwz2NzuEyXA2AJK37voWPud2AfdZwHeDSCykoyjZqd+tpla5MxdrTWiSC+QZr
Oxjrs0EbkF7SlRu47jqbHmda6XHZT+NXus9MnaTzx6SnueohYAO6fOU3xZ4wv14I+CBCcSkB2Hev
DahgS6/6lyueTHRXmbvk/ROnjKWKwQkOnyOfy1JuiN9fqz7ZtmeAaAKEjfTjhMEIw4ng1PmwqtkI
86Gu7ApN8oDJSPGBSvdt/pFZSGthhaX6ppN+o7fHm7ccs8PVlxewiMIDsKjODVenlPZEuIRmbllV
bRqt17AeZEdRdGieTWIkHGdiO86sypAj3s/71P9g0kpMUAubVoull9JLO9JPdAV2poN10wQJoHJM
GQChEIhiMEtmIEabE3PsiP+fZ9TyYkqyMWrTcOsbq2hIK5/yahsMkna/416MwdsuSdW1ADYSZhx9
uqk1rNGnDn9JRcF/KUX01Z9mfPAc1Vy/FEVkfv49Wh9furXeCaeMlyCBOEGTneIK4JnsZP6MBTlo
5e73MP6L3teqXtS6hGdgzJBdODJyr7b0G0m37dA5O+6po1gsxahjgiF5WzbweuSyKm61GL72nSBG
bi3cNHAThqb+IQNW176/t32da6qDCcy9Q5LfMkSOZdvtbIlVTdHga89XuO1fbu9Cgw4rbNGp1JYZ
G4irWWLB8Y8a5IAi8zbrWpviUy83mSvG8hKyIwXxm1Vq8VE+wx8m1ZI6H/I15kFVAw+7UFEcSrXo
XxgDsPV7xK2uERb3YSWVdLDHfnCnG4dT8h5L9wurj7j3b2tIbNrxhw6/DyYalNBnF6EcRitiRu4X
mcg8mLzG7RkK13LsJehQOizVkb2D2BiW0vWS49LkEwFNZuxprvk5Yz0jBVzKzTpssyYzudH6WsU8
WP7HLe2dL2lM9E9TB+cFnNIWUxyY51fllSXY6Vi2X6+3HDZi/z42Q45GGpKmjC7CLeDtXSq1d1sO
Qe4CtljScZK7qRJf62blcvHf+/UFoZoW4Y0pxJdUhwGpD7fQOABg629xQQFwPlm59HCs/ORqP50B
+0o6i5jN7E79Loiospj3suClKPqXdgyw3msJeHNFIph+/s/RT5IppOwcf5BTqSeZp6qsisafPsEe
LR/b3pGaZePAwx2ITAj/2D6HMnHa9P00oTylSWuknGHWKlDdxzMdUhAa59q8Opk9J3t7L3yaVX6p
yL18c7JA9pSrY7yS4lTMmyfjleM6wJNIMh38sQCr8vD9JewrFq4NYaQtA2A1JnS/SW8rvb/MKzmK
eXhDN1odWKBfXcf3NqUjogmAMy+4QpXEi3ZE57cvKa+b+qlmtMZ7xjkjFaxDBJCnqq8ZabApv19N
XhGG2c0kbE7cutHXe6td1dHU8BeDZxVvQetPKyM4Ih9aFqs3SFgO4UaLa67ybi5ucGx9/oIvcdv4
MmJuOopYQIypbgSMH0FqJHQrfTBUQ9LMpHkp9VT03FFD/HPI/AvwMOnlYQXEvb/mO/Va1/eWuLl1
0CLbNhBa25dIFlcuIMIz3VIlyc1m4rnsr67yr4NBY9mZd6qeWQPvKlKXRSCaxlwj+W4VGF45u1Ak
40FnKRahY+f5AEy0ruV/83few5PYwcqF4Yb3ayTPX7/QmIVhHPTevvFekyhE4NDUINI2/I/mh8IK
r7wccsP/YFd0YLQNjCUti1odBkbbAyNrCFODfI/5IzOI+VUx9V/izzixfce3kBAnZUTWlpqCzMh2
t6WVzBkZSUIqRY+MwWliYFAIZK7YP3gaqWAXKGyUF3neUXcA5WeiW0MQFq22XWiRvWswkmoQj1kj
r0ShmCtUvJ3YYiV7P35QmEyyK8fQMkKwPm9NwKraN9bSxWa3xuVv32L4XMjAUEjtBMEgNv7Xq5t2
7bKoehncNy0llbqhgSp8EqH/BN4Q4lpHonmbX8VeXcEzdThUsX3HF3yIenT6fGznPKnW77yrDBdq
7yPNtR7DlOD//rkROZMT/dCCXStq2xXreFvOQYTPenEY6GpQIo3zCSO/DJ9CO3ixqf9oxhO9T28d
b/acIowBEcKkgLoqp4sszVK5uQkcqjjm0lmHPwDSKJGIyP6aDhAMfiDmSKjsLqeE5KN+UxvhIZ43
vexAy5hh/Wny84O2aM0Ewi3CKgc6zGgZYyph2h80b7Svcs2Y5r5pKP0IOWigWISYcDG9QFZtL0js
X8nW9YCctF2J33WRPdy8AFYFo/Jra1zvS0s5tVnDtdWJNx3M+ur0Dk1DERowuJGHvEZREEwIUwzK
ffWRdNVKbnVpheoM0BlyM9FtA8oqTyqED88cdBBKosWzdIXitQrOdFg3h855nGZ72VQOuByP3IGM
PKjgjLXbh2OSk8bjQ1I3TDRBTx5a4CbKDgCt0J5NF/3YHL2LpxyFMMYzm9a8ZlGJCYwYOBze1OSi
HtyPI7sHxPdN7qxlZz/SPCOImrsMuddtRLSNIr7N9it/53DFrRdprO2GZDcL4T0SSTkL0o6Xxw4x
vOKWAFqSxquBDByvQ5etmR1yryXrUe0+XyhudaGfJjgWyq4HtcB7aR2wf+ULLjj/CHtssoHcmCAq
UyIJ2bLKr+B5Qiohv8XjUuMhpW/jJ0HuyLT25qiPa+3JVkMujCRMaDi8enjiaXEvzxWDSvNNdfSZ
l9dm0zdkudoZPatAZBXThJ99tfx6ym8NygdSk/2mbUBYrMCgriemimyQ/OTFlKvzxkD5ecJv7H0f
XsKQmHfrSwQwsYrR2iPxr7OXfB/aMLs7YQAKKasxJvdrpBa89UthYMaVxzfv8HAXj6kwXoveH9pO
GL+6lFZm9b9adzVwkBilJPYWPKDnz7P7JC4KOhjsLvXo8Sis3k1+rc2eGopw3RRsvLVmhekdSwXV
ThKEmHDN2VKxqu2JQInDQ2bUY68m1d+nfjCfmm7hI2/od/qXU9ctDfGzI+vHdxP8KSmquUvRxyNA
GtNAWd0P6EzyyOpy8xs6GWu+qUY/UELxcwYyR8YOykO2hsKrBRMblscrKFkucVyQzWNnUZ4f8wo/
jhbXkDHPMrXyuWyXDBjHNCJaePFECJIUmUGOk0/Tbs0g9fHNuboEZyF/mVNmkXuwOqT4UDzUliZ2
J4E73DWIMBSfsAa5vMmuWzLj31LW8WIgDy0+Hu4+1EptF8hI8oH1Zw2Z4VkxPN9Vr1VumuVC8o5k
YUx3u7ZntcOUmW6PrN5G84wU28toLrvIpzO7SFo/YJ59vtnFQU6Z+LanK/TnvOru/12G6pz9cMg3
pQWlzj5RRX7VPq+tIW1m+KgBBLuJvd02d9/0fRALcpudBgSsS1fyZiY+wQ5PQ0N+ikaP+dH1WAGe
DRWHs4n7zzOwGq70Dg0CsZ9hNw8e1bms/RioGER0cYDtCEAJjmuRHUOditWaPXhGXH6kwFlG8JYp
k32LcyY69TjzGPvCLJC725qe6VC6D3t1/EYZ6iaykIZlnN2LtUIFzBs0NBMzQzntEa99vsqeY+SE
adKksS/wXnBqkVQ8zW9A5qFZKxN8RcZsNoHewbykkXOCVyDimSvuIc7fTfsaAEAeFmuB8P2lvKEH
UwvGvX2GJmjFiN5Hg5Swll40VRl/L0nKrL5OpUtvtRnYMJPd31vMXiX7fuU5e1gzkmOWarxmD0C5
xNoJo3OxVLF7Ju4s/tXvEBIgp0D3nyQBKpYiccJyyqqDrw2WZq/10otX0OHE00v/qzK1woNWScV2
bJAxICNY66TzTktXjsoMVZZAEVO4PjrTcb8XbZcp6t+hCr9Dg62hyCwanKBngoopCMs0OxNu6q/B
cdND6os/wd/sTYUlURMEax1LVKDHUzXUtXYIRkKFIEjy0XFlOIrCF8tqnOjhnJew6WhpOXQY9kSP
moog8joiXDN6OW/jFoMS2WGravhPTucnoNxNTTfxFOlX+zPnCmSPr3k0jkgoa/WAxDbD4cWX+2EW
sod2bBNvXXbtosC1ZHKkeONtdiK8EZPCTiUxn50ddjXAIJN+wiqZGIGlzIcl/RwrcVgulidmI3n0
W9JPwHx4WUWBaljhQXAkm/iFvAqyh0ErGLUj7tjqDzq5rpJ1tiu3BHJM3OvdJ3YK0wkuSYmCDrUW
nsWoJ50+w+GQ7553QalQski77TJlPmZ2tGkxukm8CXdFTSauO188tqyIIAkCkEd6X3w+6+hVhXPp
pF0iNgpBiXFQioHFIAfZeSg0+6uHK7QrrpqL5VwX5KWVdrIuKvc3bcwSkVnSnidUELaxnOsA/gil
LVuG5PRgyEqgVL36pehY8POG8BWgTqGwQLbMW+MEdYEu0FXjodHxuRdIJqlxxsjfdgPOfQ/zIUSz
wdpnjtReTuuvDE/uQwru/nVfe0BTA/U/3RWdzlYeIL/M42FNIt7eZUatObj5EEscPRMgF0xoOU8E
NzA2OwsjSQYhSEBKocZTX+wp2fhcO8R3gje7iFKbGTnVgeQuOjH6D9VGCBHe/HAgaa7435BCB7Hi
BYjFJF6k4FfzconEj4m+/zHUn43muiGa7efY2YlgoZsHM3JTJuHR8VA641qjdWYmMT7B7kBdZL5M
axP5ybzy2JM9Q3iZXeHDikhcySuXjrv8tY5PYWYMtA1NWjaXZ+nJttUoslV4751NqhsSSB3y9wOV
qOGEu1rEQYTPf62YmKTRMacxD1QI0QofQDHCO+rwIMQJlwzV7g7nNWBZJUts7vbe2PwxII8VuzO3
8T3GUtxQ726oMcPqkATB84C8jdxaVZuxKBo6limSBLfOPv/iBYMLk/jWOO4n1zJitKz3n8LWq9NA
7F96G7HD6uM+Vm8vXMkNUWi0JBopZZ2OfWMDVbQ8Hne47teJBKxg7iAbmiGxHGfluQnyl2lvyHpK
pQ0K6Ece7sFcgdadYUKWORteINUyPkOHo/qRYSpRU8+qvlrW73iikvQTvgizoy4IFYoQuF6T65kc
YcLMzBNj+f5Lbsg4BJMgGnunPhvtQstYIRvLNJMsESS9w2u+W9frKPiJX1Jso1WSAkoS2eZLGQQh
1YBMpb+/v3yIKNzUKj7iUeyAaYFv3UzbbJqrVo2VwoTTxombMqu54QTEFpgLRYw0siRRr5siE8Ms
Mp42uAGMTJS/nmM2cE+TplUUX0IAUcBNxfJByQ0jc8Sutzn83DDkPB6fQjvEf4JsPyXhaqRFjIWa
nW6IVpnlUWOXk8uAO395bu1G0J+FFSjf8EtRqy51Zzo4XqCgt4URJ1bE1i2+h4T22zmPjAeg4qrB
rFE4SdULJdjx9R3TycgDTdAn6ChC50lNaPKnfhrDvFGY+g1SaHcjHAWHY/LwffC9wZSYc4veTmuk
M84RRNgCgkjz7P1ZvDx7IttDkN8sOQ+F5RTicbI+z8K8oMIgWIHFaeYkREZVr75UwjVGWKvS5RSf
jXbdjgDIntkHUV4lOYrQSlr0rnns/vJzwYdTBPXV7Kz/to7fnepArvK+nR5dpG8bBEazoYknHtGo
bsb+rjuEoHGeEoH9novu2U0WTYP0b14HmsQ2ZoXwhiqWwW/oF5dOHBIvJ8H1UjnSttc4IU7nrc1H
r30f3F5NyakLqpQiCjbS0eNXFmPjsktbNHEWpao29iMf6RlPbRo8vZIj4S+DEL3mtqYsN11p4w22
T57j2G0nAUy1yHjfE0UuJkTr1WHQdrRQMBRK4+E3TH1rBV/JlnTjKXMQEQhWnyXWABWuF9iXdidE
J4A/RBRvXITBKsUbrNT2SudZ2tvuBh0qddTyYC58LGjgufR0UZ0wg+gSHSddSRgOKvIH0IFc0TtF
gqXfrgtFx5O2/5TYUBdwhB42+hkV/5M8SIrJBb/kOXxrhHkCU5SZC2m+cyAejExZyojlPXnlNKxT
VJGmXCdYOrHP1f1k+DvZ5XZW27LVD7Wb1AYH+hXzmmaT9YmGARUj2rx+EzRL6JQPVXKgxJGiIwnd
RNzEtfyMQLme9/1/sYorg017D7Kbt3IPeVwwkoNSTfGT1snjep9gSLdJOCDYWcSwmPCcwdcMg9wx
GQ1rAaYbqenRSrEGDclevgayC260xIXV4Fs6tSIgAaFk1ukabQDZnoLkyp9Fjf1CEy/1TiPVWuQv
wcN5jIaOOfhrLlCGqkP+v/O2E7tBe3Y19LQOtb4feinnS5Qer0SQs7m1qsob0HkJcNT8oYhwuzYM
X3xGHhjXmLPj1W93VZdGqDaGESjKSr5dzNijYHeZH8QrNjHz5hZW+QZHD2OiVHFdxz2qMWknhoii
RsQn2cU29Ut/dGqaBvYZ9xab8jfBMUv+TBoPi7A7/mAls1e+Y/2rOyrQ8sfxCXiqCpj8cgQxe8A6
++48leScdKcXWKM55lAno41tHkRjePQtkVRRJ0ps9KtJCRdAxbZ93UitXt+dHM0PtX8bfQoUfiYs
UaBjBZfw5RdcWC+znLqZBCjD4MY7JwBYXTszwwGlSvBJB6FyAqIZYJsJNg9xAqvFDBAZURA0espL
1fZoH49pZM+bEjjofqQSrnFOJvce2Jsetr4m14mOL1cfg91UWdajo8WkxIBiSawB/ADZsKd/rE8c
U8aM1V1LxxoKPhkt2OH5mpOGELG8oPe3/mp3dYPzqbT3JGs4zA4jTEV7lnZBmC15u6MHpOfSKQme
AKSyazOAhFS76fqsvxGiGVGSRGiv5mqsi4l1UX/3kp815sN1yMYOw3WbgYR/bseRhWeMJuipohX1
2AGRbTmF6Fkbq/aeLbvqOARQrYmXHrdf+6YhRErtvXKkwVdpigu2FFgRk0UqH7k/rx1xz1hDOzNS
4rkiRjR+Exg5zNJLfoyg/8qkmDeb0rOn/zI1t/xnTxr1qTzglY5ZE2lx+J77yVb7TQaQ8eXRBQjd
VFwiazH7jcDRxV//BDh/z0TQ17wnU4LoKLmsZ0vGsKxA8PsYw3UHs+ye32G/HlF99UYFVdL2pdm3
HzKH9nfJlXLl38O7IATO7tOQeur5QoFrIwlQI9c1nrlkDo5T0j8pv4bZBFXjzTATKGGsTsUxsLqK
lIgJ6YMsvetTHWykkPhmrLP1oMJd17RgcJhd7tOE4zVo4vDZ72ZYFLVsb/Bkaala0yhdj5SgYMhP
qlt3i8CMv/sCghAesNuyE0OvwruRJOnf6x4b46ZfyhnRZnx84r+Xoi+camDh0U0ZUDXregMGn+uD
ATGX4/1V3RJX4LVpiXiWya4X26HggcLQkD6j16vyxjIw878+waWs8VJSd91PVxFPJTWo7NdZ7TO/
eaWHcnatYGCtMNOMrnzqlSKx83R3cNqbspk4gWdq55O+z0U2r3ogJI995gJJfL7SdrjYc3NswSTG
5DuALP6iKrGYQp7kR2Nvtt+AxT3zh9m2w2CGwyUrLYRNPPe9SJDxuTqw0ZlhG+C2KCcSShRrGt9U
6x5TzQKOBEmZ96hd2ILnyNha2XXgOyoOCGCsti9z/qDnm4EZKbolVy080+TXjtSeszxf8FOEAB5w
TMBMvvidjFOIQ8XYrSoW6sZp0CfwRPY20rU7kjRtW6KO5PB7Vsgn/dyJwvRr0Omxhrg8IhmtvkcL
6jOMfXv+bZQrG933x9VBlR7H6ohGgfb0tHPS9NMHzbTjlUCUn6O81sRs7zbK9X+9K+oJOPCMI3V2
IwjTy/q5b+mLzwKtXzSgHNlWwLL/KCS1oNLDXBB+XsSO3DtJYM3PNqMWIn7EnCSyiUvlXvz7haqf
TRYgCV8t7bvdF8XiSfIm+CEoQ9ji6MLpv4laDq+CDGwsfX3i1NmGwck+zWEb3DziCxc4PkQDNePh
K/6h5CttHTa8QdjjO2TRJ9syIVJMTBzvWRcIftV8zjfDcNDxw/zlqBIXo/cumXzj8bEF5JJMxkGc
Vl9XsCSRMV4xQN/MpB4OE07/SlrNtGms4ddLl1VezJcLoI0oZ291ROzGeiGYMEdJWqEZFNetsJmt
9PRpEH1HyjiCQvjPhQOzWa1pamHFUE4mFihjD6N/bBxNQmZWmool+8vI/BW0NqERwh+rBA7EdPv3
SXVp1VWyY2sHdHYt5gSg8Ie9IE/Oj/etWXBtpIIFrnI9ljur9/wq+ScRA1Y0fHZc2yPhWKCfMCy/
Ww/8RW0i12+rRJiG+NXOdM3ebYBww7MR8+7+zHfu34Gax1jQyPcyoxU0Ia00XDvHc7+ZduJsNwr8
QaOBZpZFOjsnCfrgevNJC8V8/miVrpvoK2y6r4UMf4WGC91/Ma61lqQ+b9+GEKcUWvWzzK7THbdJ
fCys+0imHCOXqbz/OPr8GKgp9AQQ2vzOWU43Flua7LvVcQ56Xo3dGURV3rx/5nf7B7vVajJaQYZO
GUq3AEwWKEr9VrlGxND0sQDaupD0pBOMtVdWCRVtso0743qSdj8VEIrGzWNe3dTT2xmOstX9R/ln
KMnEB9hZdVvP91haktXqzcKR39MlcVk0N9iscRP7peo49cReRCOwUyhBzkzNyw8UhibHGZOPWNqn
mji+bXPV4nqx2f+CNPkrUhDpFzRAPOgt8g4XS/SvuAcOAN99bydWGFWOQSfXsiQ5qMMOwwkn6F30
vfxXQkpB90BCHaDq/f9GvMYPM0tB4MXKuv9t2JYBd7NQhXC3h1KU97E/6365m+Yf2a2t+NOnZ/Sc
PdvZvDYZbck7N8fipgLqBOBXuihF5ryYZWFrJpD4jnKIPA+iNRJpKzD1sZxpXMgc0923BH+2SP1w
ATT6tS+8OzPPQbTtmNR0kJ2Jlovmo1ov1AkKSfD7lc5thQM4CSrabO/0wO2grVyEBGcA9bOUjetz
U3ucq0E7Zfi8sSgOjPKFjGBlPO1LAAz/JYSgq0In/p0luA5DDRAI1eCSt95TJB4Doag2aIv1L6K5
eVPyPsGDbQU852tsoWcnDLI98RQk8uGvLbMWTTHDHfphguB/I9nupKPQblyHA/vfzwOrigY3xT5W
y2/KrYKDRIz3GKIr3rHMLZFhiUdzk0M3p0kScnLCU7Lo/dOSQ0CvD4PmUqsj0EFbB7bHk8HXzDpl
MqltIuZu8j6mFKe3AjzgHZ7h6Hi1xoyHZkbCPU5SVW0EkJad2Lg3iqYBxwhR6frW/Nzmu9Q1Xf+d
MKt+4ZO7qJWmujFPkSg4rdKOTkvFJEb5Mxt+p/o9FX9KX5qVkilYgKxaSKOUrDLp5Oi9DdgOua6i
IPi2RxVomfLfgL0FZpC4rD8dQP4H4gahG07Xu59Byo/Z8SbudltD1VCLGzVTG+ZKNmKV/eeExthb
AJWGs9rJidUah0BqTCeaG6fUAPun+GYuBqFdwokLCJ6mqxTpJ8CDa4r3/MdMU+PnmIS5+J050nC1
a4YVLZjepq8GmNBF2zEXW7SOlLmMhW6TKhZNMUVu/AwoGMXt7EL+wTNLu68mCcGwagAyY5zJG1j3
TWE8SBZCSNpNfahxMlF5aPq+hXgQde2cX5OJj6GDEO8R55uJ8baav+GNg/DIsH6bi+MRKkJLFRgk
SSVoM+HAsawsPv2PuoqbmdwrxxSKuo5ZYiYC9eVy7l1abZF0Ke+La4m6G4rD+FonkmjOOAaSl2ka
9B+UxP3ZuJPB8Oo/+w6xNGPrwu+3wS9oZbLkCsw8Hr6y9y6SH5d/j8n/42LL1767tSqGYJYxBAUq
q2R2zgZUvbtKWT2CQlBABqcmTQtQLxfeFaopbkgZNQ6zlLKck8XU0h/qaQJK7HtoKdLpT+P6Ax0/
nzCT3VqUG8erHaI5KdwBCxf5CVMdI9uzt9fO3juwOvJEKhrC1ob5aAuKGjBbjQhaSQX/yPwxEWWz
po/M0EVjj2gX7kPpqNeRO7KrtD8f7v2JKlmlrNHKLXtcLr5DA+spusCNqjDl3dHFyt70KMBgVTy7
fByfqECzuckaVq5voBGhS35lO6bcyEUT6RiVmyxixQR2P4W0ZR2rpjvPj8Wopmkuwh3nJiz0f63q
CTe15YuP9mXvfAM/w58gxasSzara3lvWeYDmBBykJr3S03tahf4LextlmEG4KrwdiGHLduJGE9fp
Bd4PeBq7jRmXNLtGylIn6f204idlQY2YrupHBWVd6lXVUkNR5+odnNcRX1HRkjJW1Hy1217Zamkh
bo5gEKEo093TU5dQdcCGQBtVc9iY++/kd2aLby4vx7oTFu2viGN9KrmcX0uzNJbLCClu1ZvZ9hK/
TCoZN0F9Byd5JoNgksuIfVSfhOi1LCl/mUPB3izGitq9HVqz0mjhAzZizg7osgEye4+NXlMv8t7+
B4JP9rfSzM+b5XcIKAZJLTg4z7IIQfSnIvai4nQXqpfezxhgX772PvNn24DeFDoh177we+b1rV/R
rmaQzLX3InLnAy90DUkX4/dlq0K8K2JMkpnQxrcxiApqK03Vay1o27jFZf3zuhnfS7+ckwUR86O6
e2aVTCL/brqqXo9RKFYjKO9gHpkZJZkk/zEr/nvwE1EiyQgaGWPPkK9jl3PnxUV0bDnV0DRwi7PP
mqBaUR04VYvwO6TyE2DI11HY8C1aCBR1w3VkTF0Ks8dOPhSJo7yLcT5LUBCiGsFZPVpk0r2qIc4T
upuUTUpHVKHxmM9mNRHKeCUKLOHfWFKE4VFp93WHJANt0MfkTn+cOsRMdKjAJprfQypGUUGYJ+ut
nzTVHsOkuX9WxH2tpltoZ9wSQSQXts71o7EZ7KNJUbYtB+4xSHcBvkECJnw8QaBZc8442RgjYGy7
/aEP5QIxXdeQDbTHb7uuV2Bp5G+2NkCXXQRkYFBLFWj3FrNcXm6hiNablm9Fc597yd+ypTXGhP77
SonymuJAflJQkWZ9QKAhknj5QE/2t2TfIVrbb8U9H7LFL1JY6YOHT/ztLPtIroGcGf+eXcQNd+jk
69+RraUKBr5lrl39D6TnqtqR7Pe+zYaeXf/266aOZxPVYgLWf2pset7nYophGxkza5O+8XLERrmR
8Ya1q1xzFuxt9E2ogQ5YRDuurCqCi//MHi8PWtKc90ViVzCNjRCJyv+4PEYzNDRvKZP0I6Stq5Tz
3E14l3bVenVYiypLgnAKtL5ZTWTbtQsp9NcLcohwl57hpQ9aAA88Luaew5dV1lMZGa48u8npJYqX
h+6hsGnBsuGwAawRvtP3L9Ya4vasDCd2Z3Z+I+2hanbmM/gGJ8GPQwlK230dAGjkKZDYodC1n77y
942vzfCETt/DA/KQb5Tn2E27WhMGNeJJg3ZNntcWb6iuBDm476s3g066XPd3ai4aAHeBHoRm8M0E
k6uWb2QNiBiiva6ZjUnOZSOrJxxeyR87gmYuI+nnK3nAdKvaorQAICLMx698CYiIF1CpIIKzVbfu
gstmH/GAdg5mOxy+s15989S7UUtnKvmiXiHWUA7Kp6c8dsKjevFW0pJ2tO58FX0gyz87RUIHKqWU
Dm8OW7pNDdUGLsshyi8ynNKclq79hOVDIzOu/GPsXAjDc6X7W/1wwpkWxv47tBnSNZN99LyqR21R
F+o4J3iNK5srbCQ1gT/BF02453JtuiqHagLHRZpm5prLDySR1esnaOTGprpF6qOwzLcxYjHdmvQK
a/4Cmoxbf1AAGll+TmlcZqn8XjL55IUuUt2vt3g/mSix+n/scyNyYmUOXniaY6mZYTLny9ZBfvWG
sZ3rPaTxKpMcU10635ub6SfR+RPzf3WkYOLIYZHjTyQ2aw634jYlkpdHf1aattbTVaRIkrbp1KRF
jnKrmE9H1hSiIp9TugXBOhuRvY5jvsVYaW3hsvDeDTGpeouPYtMrHQ5D8dN0BYQbeCUjm8JFg6hZ
BNVYfDBBhfy7ZB4J4JSIZfpDvq4xroCprqGJK1P8M7m6XYdo8/wPCXygMTv3mcooCOdpmIldycUl
Vw4CRlVLP7DrE2uT0P+cRMlpBeq+ku/KAGGF6Jawwc5xdKjBuJxiu2DH/NqHMBCFNh4SDN+UCfYx
AAoDihs5RctY5kD6oxcye6VRlaFZUxF1D9yR6+BFTtRZ+IzmWshtbXn+rd75spD3iXlrWO7DK1JK
RPM0hh+kDANdih3J3U2ZQo7iOa1h6ZZTyrXU/t1J74bmIdinGDqvFzysuDMthAebl8CLM2jumG5k
w/NWnkWdDkCGlDVdhBLVe+m6Su0uz8N8cwZfHx2y4DAjH55qs34EYKcuky0ZgaYtpK5iGLEBa5lF
ofMg80HmlOrWgw8BW0erBIsTawPEjP9q5GutE6tXWNZbZbN3gLQPHB8Gwwany4763HTAX0ZTNXMZ
NTYXPBJq0FrnI+hQoZXn0Ir8/SomID2XK6j2TRol9yFGSQvRpuI0wsWLb20uLJqixQZkwG+HTt81
RC7MYYt3GzUR96KHfCLDmE8NoAdjtT2pYG+1IqHnTa8glhfvA1KjGfguwOgeqiTYNd+DhVZx7dgg
zAyoXVijYshg+1D/hfDeYwKbk4lFRFAcsSzZiN/yo9z6udnHUU67ZSkiOWQ4/J9hMh3Im9ckF3B+
/7b8NftyVI1m1bBl9u+NtHBhfRPCV1Ksrf5+UuIzeH5wgWDjpsLwDcDcLwxrl3vBADqg8zKHgXBq
gTSZH2Fr7v1n5Y86Geb6L72/SYz2eIpfUXdrPrlNeFhYk99CSel6PV6jlCEqWlduudKglyEQfL4t
Hm0uEkPR8r4PSm+aiJNO4F5/Wiqj3tuGE/y4LrJkd/WDgG8hnft7S+27gPXXTHir4Y7cqhxtQ5vZ
Q3vK/695zoB0kHJdMKAzsLT8pDtoy2wZXtq5+FND0hMwJKmqs9UsEGwhvQgL+isNPwQv41ac422H
0Ar/cfX8bz9R8Oa/kczz2VxzrMouNmfafKY+Y+LM25aCD4iqNu/WSh30HoWsGwM0EKHjJpFMFow9
oru7g/3Z3ulBCvZ4UJh8p5D6bbkbQvz7MZomeniXuz54T4RLa19Moj0ovERPR5eZYNOE/ld8Rzpr
mhkxsK6QQnO9FxRStUPnNC6z+WzJXKEJAQuOqNoitEWzmMtmomQ4jlLJUdrv/76BB04srohfM9oy
oSSWmRGlm6c27FE7BeWNpKmbcjcuHcs5rGnbvzG80v4eECKoObxBPDVee49sBxzIlPeWVhAe/dA0
oFjB0QH7q2pSol4sBgaRPMK+Limy1Z/VMYwFD4WN0BblOX6GVT/TobUJplPyi0Jua+8ntjSOMmfy
tj3TdsRIg9YXZGTwapv9laD3kcdFhLPOPWGeYEpOETkEgHh7Cpp+CYKxWjUd/qNkgEC7h4/6vC32
47AclqVz+nP69qA+n87lO9bWHZwtCk9HOgryzoaS04aTixd4iCsUvgtsO9YLM60HPDCd8FLsXGJX
O3B8Uf7873GQZ8HqKWYVYxK4sfeBmO37n4DtJMXYfv5RMO18Bw/YkuIEqgvdL/EZmuh1pD/mffKn
YTHD+NaTN4HgpVQDIwSNIm+7rz6skzKf6EhBeN6WFRH7LQNuAX1E8BdnboyeULk4DcT5/aXty9cN
oBF+8fTpJA/pgnsU5QCv6UPYJYkPISNe9WrvZDjFhGWxj4k0qU3TKJkmSx7oFgCfziWWSig9YOjH
qqF/R8/MVnUSXdQIlVtyYEPqparS+Exw+7PL1Z2l5uFSqmU9o/n3qS+z/bWyGNFu2wLH2LJTN+Rr
9YuK3tDyhxtKXOhEZ8tcNvzdIQEmSRKv8c2SNbaArBmyn8nYL6uPciJkphF8+ybEnFRo5hE5l42T
zTejGCmXWfWo82xeMRcARe3RKxIT4oyLWQ0VZimN2S02BaGy6a8cYPvP3aDiZ/xl7cIaFJQwTBtp
9mBf4NXIgrhhLHuvbuYQK55QP8qiTsL1WTABnJ0PlxbaT2oI88AOrH+p3m2SiZnXExnzf697Y2lH
Gw2SWr8YGa//ItkE4mXk6nPTa73ZOxcqCOSUM2SR7H5TMgoCEXYyNzWJD/isrNgfcZ2JhqPXgNHY
ClITUiSMcDOrvx7D5wOsLJCfpCO1YxgTmvBf78pWDZeyCW38ZMSXh7fg/obNTyx3DpXlt6ViMuId
KjaTDj2yDmHvwR6bbHJfOXnhNJhJOC4h2KP6B0ub30+Y0mlIvzYdYD7HC3/u2b1P8FkWiBddSZuu
HbicDqJRBd0kaMNumjiCBq1WY3N6JVJWb3la7Y/PHGjw+N1+FpfnCxH/vljw8/r5O4EtUO1IL+Da
1Wr7N2ua1VCXNgN/lLAQz5ognTlwxHuPT4PKViqj1pMgTyDKS72JyFGHuS+Y6v8NfaG54uGyVBZy
oE/WWMN7UlawaxmZwBIdPwqDcJ01l8L1nHp7XKsP8Ia/magtupiaoiQv2p7AqOTlgnOe2BmGwHRj
qWYYxDHmv6lRlVeSiL9V9txEN+xWyqngAxbK5z+P7pItOcTCcxe14jr5c3EcdmIaxi+OnhX80mjp
qvnU2krx51ZTMhFQIi0mhHiUkqcvbJDghKQAO6Sf2B/dXvNzjyVMIqM5UdnxL+TeDoBmvk0qDr7H
J1LmqCWnX7+9yV8hHfGPtE6NANR5wWJNNiq7eHma2jMGeuYPpm8HXIMDjDOJ0nXxSZEn/obVDunF
ehOgMXji3ZiW31ZbMZjVXAv+snJeH0QAr2YnrXLy1+eoKn8L2CCOwJlfFsFh8E6pa08+Gqw2t6IN
i1wyx7JOgT15Nux0oU7AYq2kMT/ElCXOl14Ka4v73cpuN+rECFPnE2X/7Nq8Fg4/uXkCqf67ZgQy
tiAGqOmuAYUIVICw/SdsZP2gmq/Q3Z2nSg1HhnMjsRy5c1Gi4eOOl5BzXaasagzsoZ4sxveb9g1a
KVEoSQpoKp5Kgz16Wbdz9VNTXfhSh9JK8kx0YHK8V2MqESa+kG5/9P5LZjb1lCQLBwWso+za1oum
FrhYcTq2ud3JaGTeHQO2B6m3ZxCl469Stbv/+eA8A+eeA+s9nCeOBk4VEsAOROuBRKDXxZ9STgHc
gBGKLUzgiNZxbrWAauZObOdRcJjXHWa7UyGI3qPerMEX+ZJ+ePSgotbMAoTw5yiIUXoY7kwj//1M
4xVcMfnsuTHOgMggH4Z8b9j3xbkzm/iGgETSG9wpu7rHxJ+Jo1bl0KOQh8HGdqVmT7jy2q7vfGFC
R7EyWC8hAEIeXmH7ez/atJjGCf9dsbL2pon/kG+LNj+pjUa560aseB6fri5E0uKbZK8se6WsZbur
3lE8H9rJHKsA/9RXDL+A0gk2ZJTeSv57nORxP89ST87vinjCe7k9g5Q5dPbMN3BWY1RRnhm5X1ie
LW9HPYxX7ZetCUV9S6SRwwB4m2nIb0Wll/6g2wO8fg/8Ktk08oUmiemoODqvp610JAeEf3+TTwaO
RuHVp6ILLmOnCu1XpM/MBKXZnN0ZNBR2Qm6tU2l9xqaoUkyKjYS7t04w0mKkngSuQJXxgP0Krh/5
BnS5mZ1J+Bsa5VnZu1FAjHEFJRAtAxbpWkIOqw5pMEaUptVp+xlQr2nLm71Ybr42sXAmJ5FA4Jcf
S9r9oywkPH1yA1cx9OLccps3YlkYvjVbhwX5nyREIvtxuf1cLUrLk8ZSJsv/ZAsAp3015cEYblnC
3TjOI36PU3EnTWsQ8iLBoV/xNJSnIjP7o/7w3//Jt0HavXSvMl4trR0MIRoo4S3fFLW438kADh7Z
Ho/KvJuM54PI15fGJ08AGTCcezqAIH8qlYcDFdfuNX9oAACuMNBbi2L8IMd3JD7XJg+D8QJrFoct
5BAJCtJ4jdCJaPqO+hFTdvQ6OzRcjyHQVisnPZsHvZrB3Fp/rgpH7q8uK2YFLA8zNjZHaYcvLYYk
KjZ4+JKBOes1RjPCBruDL2E2QC3Wh9pB7ZmiP9OVGQw2MYQ+awGsA9iVvEJ0cCkmDl7MywK/fI6m
MfPkJLKm9INWCYpcMKn88+FUNo0sovkBJy0ifCoiB2mwtFjirDN8gh5v0p2W2o4U/oi5UpxnXRB4
WejjxOLFa4pTjsLgvLKEukS3vjx/BF1hnLvIJB4Q7+f5Kox6R2FKqv4UzcLAOqPSS2peuikRv7MW
rfJ3mOnwNMOtw3EtN6363XyyFq/EbxazogqFqPFHzyVaGbpiZgyK6KP6xrnjDGjEMdYs28ub+MCe
NrXY2VcA8dvE2doiTcxGfPReCZFq+vgOT6phjKKlRDJvmEF3Ttk10GIzZGu1l4SxHbCvHF8SAOmP
3KyqdEcVqWLtGxiSbTJfcBvySmwtuT9UxUY8K0TdtVPL4wo2n3U6hmaFPjoggndTawF6fxxa+Fuv
jUxRn5K7wdBpoGC76IvSxPCcD5x8FhzgnoN2lg/Nbq3k+XISJgalbYqgCuJKCtgYg8Rd9xb+yPni
8nuYXDNfu17mYtuI2h0zP0tQtZ6xMKH1IwYmerUA3u734neb6LiVrwpDnXonT8klM/AyHUwcHkF0
xGCzN75Vn84BgJHhrfuv83hqediM+gdfJS227py9S7k5wZkZSvrtKUTQqVMlj+6g9RelbhkK1geZ
jhjPNpX0t10Hez9RtF/8Wgl52072deWLRGvimLfCDygvkd8SaW12/0Li/oC2/fUkF7vfD5JP7cF+
Us+52NwONLPqBxPeBCmBOjepGLAIUIKtMW1ovL8pzUc6NujNpPTFMzo/w7DF5nLI3zztzU5bQFS8
zYLpyBI+/RyzbYoJ/6K5GasHfuEMx6ToOGfyOovvM5Ub8zuzBp+q5cxLMIs58xKJAJaojXnpFOu3
RcEw0Zptp5bKmtoDfQPupt0ofqP0Pram4R2HFSj6GdNByCfRiEktgbTmbPv/vk1tLf3TTFhC78Lh
y8ljiCkz5YrK0b2JZqM6pFoikw3rjBZKmSF2UiWDMUyvf+QSV2nard+eFMkpoDOQZrV92NC84vGa
j5LT6U+YtlhlY0oV2s0u3d0CP8FfA4l7d3a2HB0sWvlbOxioq7y3DtRF0/kIhNaxTXeFE/3UDaSf
CpBERiBmOIqkVuHvTetf8wDsoSl27r6FDBq35F+F3kdjGMrU2V88A22YcME8KtBWxlknNPLeZ5kS
8XMcp0a9/euvs42gXAIPbAPYFmG8BtwDagsFWEKHLLI28oNRAQRPRBBkYWBZWhhVKEJOe1rJXEuv
qNXCzhFvN2QePNc6rBIfLOkSw3HaQpoLmW+6FGcCUC857glBaACfWDSeGyQfS70+UXZS3GN8xW4T
pOjq+sVUq3a5AA+GuSfEJebybBq0maFLeHnhw1IhYXKm4zVX2ye7rj11xiPq0Z+HcXroJcC9qVY3
VEd6XNPx1A5yPTnVy21Vp4e8t6A9ZiQknvp+rp7XvRYrEKXZlYTH12aVifTGkjXSGQug40kCvg86
dK8Ooxa4k6HXH2uxq0Av9oK2loPB4f0adXXHKaKGfhXJrR1lUKwCjfyYRFa90J2+JEhSQak3PE2t
trrRV+YdotRIoV3SxWO7WC9bqVNAGBp04dxiBGgeyBh3PtKTPnHCSqTsevBq5TTTuVGWhgz7t2u7
25gdRZbFPbOde3GDV1JJDgdFyewCbJabnJEOKQJS5Z5PhF5O4H+tfL2ORePpKRpooTv6AVFrvhmq
YEE8CUUers99KiPvu0U3/dgLrzk/BpmeRGdjfTl5nBPfJEml5UJhF14jCyuOnuuEo+xMeS1YmW4o
8p0sCJJC+KD4EDi24Yx7FpqgWGL3AEWpjSJycaZq7frLPFzI3AL8Cq6JV4LFfVyue34IhErr/vEp
7PXxLMGXqXqpZ79fP7/AaLKCjxziXo1XLdrCmL8siT5TiSA80P1h9hyFtAmQUDF3uZvrDwRFmEVv
T2KUFY9dK94ANgPAKbMX6brVrVAU26y7+ODWSB6hHqkRlXQfpc7rhcWklJAj+TKJeN1hLX/FiEpz
AXLumP1uhothC3uMX7LasjUEbWlC1l7WSDJaTZ02E/i+vHPBwv7ug0cFvr5+i6DZVyFThzodelq8
DlZ6MDvPaVibUqicH8UN7EHId8Qg2FNLHnw1k/2XHUloQZ5aM5NASA2y2KjxhkZCNyCPZiUDTnw4
7zazBvCZMmGCX658lKNlhKXhbb64nvBj1I0SSa2ILNEJadr7mJ7gg/M3jGqPN2GwA+HQZw4nnDfR
9R7b7TqOwqBSRWwT+eh/WGlrFXrq7lUwU3FtrYNX1CJvEZbUx0QG4Ul7fEQ+pxA4dLMzsj/+JASV
/vN2eohjjCOGNUA6Ig+P7hWHv1iwJQOCxSx0w0ab8qn+MBkWJ4lFRep4BjDilgngQBNU01yufeTy
NFa+J7duE/IjqHOGvMQzFN9LK0t2VePkKoSYRbNnwbd3koqqMXwEIABP7aYOoNfQgsfCYIPPiv9Y
907vpAO21r474v6sERD4Xjfw3Pmz+FNLA1ptNKjl948nzyJdrIJPbFoYpnhoJu8YYBAmU0RwPReX
dkpfhmYPCE0EzEfBYwn4ibLLdTGM/WN8/GKOFhduXMNSB00ElNbZcg9lIkaDY9VLjN2raO1J1K/t
DcOJcoKlNZjEbDR8H1GMn5Rjv7giIzMSFpZUgxXZGWVbkUJUB0utTJqoOUq/GBc8jvtsxMqeywKK
0+WdbUzj8iYm442/6rQAQhaRc5O0N+mAgvPf4rhpxwKwJqT0mFkglsa53aLNnzjaZ7oGOzivfGJa
A7ARO7BBtBLwQZMJIyJw7HmOBjrTnO9GpIkwupt8iRyzsQfdOLW5NOGJqmT6wboHonprdQgU8vQB
AweoI/ouG2VPks5tVXwebFF45tUJ2x3Zm5aVJpVhbTIzXazO+uX9HwAzYY7Z8najqPGEW/zn+QdG
wCEHy6L/u+MIPt8mT1KrSA+ze0S6c9LLIXuyMzUXNAy30Ipz1fn+Nl9nQVs+tHTIZdfz8mPittkl
VNwNlzR8TgREym7DjIcw4CCZGMT8hrVN+QkXuqez7m0WFHDONSnoUQXS2eHnD5aGMHrOdrT0bTw8
UqDj9/8IE9yr5Gp8jjCcVtJS6W29IczigbKYZ8IVkl1vcLtdfRgg7+8/T5ViZWsaT+z5jWiCKtxI
JoVXFnLqKY7pX7OIqkQi9FjJXXKMCKLhhktdKLEa/oPmLN262I58ExL65yngMFlxYZnYCJ0LxpD3
rP5bWfnIOhPx5gm0VxdQ1inB7690Ej+q7EDn95bIwtLv/wZxbSrZi7q3lHajH53OvPXMLoo5tNh0
Xn5I434hL7Ds8rwKSI9StJtLbuzttUqg8N+DpFNV1MiaCjnXjq+m073x3NZYG9xwat17bW3Yx2E6
mt2C4HKTzdTFEuWbMlFEbZ5UakpFepd6gTpyg5T+JRUttfjPMuz7Elvz4iPDzFVEEkkkcFNkPyVU
cMYIuTCAwNvJLwLIF2ofK0nvL7x9tgnrjklNdyclcjz0QgjVxMo4feo8CIF9B48XChykwxe8CVdd
mdm117pytSedksb9NiiewylOzxYr0rc5YO1VrF/7iWzy2M6yCaLQopze4d+AeGZjFmytMewbRqPL
QoxQm8dvfoW5cFAt2KoDC0KbarklC7B3JwIiSiRjH0w3Ok15hZHbh2NUu8JmocBuTjJKybMyzZvm
ZB79inQP8DrYABl2Al5IrO1d8ccYiUGYXTF5R9q83GD8EH8JVhKAgcCH+aCXuwNmlDgr3sBhn0Rd
3VqO3HI19GwQHXmFIVrV4sPmMShWU+kqMgzwx/BeX0V7gHtqlAkQSlRS4jNThxiQCx4bCXVKS/ej
CtknNOvD8vrQFPyGF32CL/Kw7cJh21B0G5pbUyzx0pJtliaD59A1aBzV9ud1RmBUY7pBdxVNLpZ3
+DbhWfm0qr1wXLmxTI9iHWYQR70eFOyoE0gUMKAeuRXbCpGSLXNtJHYG1ZzuouZrq7BrOADrILJG
1Q448wtIS7mNqoC/wLTZbSHOFHJWlJSuD+7X5UPL4t/3qExNZ8XkuFUa9Bi7/9VWx48iH+AE6uDH
s7atzFMmOR/LBEMK7qx5UbU/cUEbZEA16v4z0ZfyN1dNO9qErCdHAOlIrjvFTPpCPzwgefwxP+XR
zo+hPWNamZ/GpJB5Yb4PEfiDWxtf30WtVueTEGWBT2bQit2YhYyl4Rpc3WuYzC56byV04iZkncIe
wkOFAcXX1d1xgFV0JY99LhgM56GD30n6oEjP9g9nUlPDBRd5wzxVcIlzqf8D1UO5n1x8s8pBuo3U
VhNEd1H66byoHR6M2/4YYgWfUnCrpvKnkN/qnbcyBLMTI0Lj6zA+KK0aH8ezcybpK0eHXTnptp7G
il+xjtW6oIstCiniNwW5GwwLaFhV+jniquXM2hXamTeF52pzzmnV0PftUQmBJ6Jg1vGUCBWeMJA6
yeorncyKlsIqCB13a2LtINiWL//MNkM5RVzEpoc5nia2WtEfjbhe03HHVgadPPmhOkcDggA2UHo5
/4AJRSHEBIuwVtJ0jaZjVn5jBANSlArmUxnaE4Pl8uBb1PEnB7zq+NKDmgfbVNyMzUUTgAzmGPU6
PboFHUD9f7WrA163uAnbeJ+0Hfssc68TOg+gZ4W0X9dH67OZ1Zg4ANgTsfXOiQcdJqLdoCpHRN31
AoZFQHjqRdwIfBakMt/UMNQYO0sNedzp7psCT5fKKnSXwlwtG+Zw92NeC4TSLEpts/QtEDBgLVXy
7vhg42XA6pzPhH8oB/MY+am80/3eTNiVed8uRiAjgljgmq3E2Dr9uA3zEMvFa79NudfhMDakebB3
SOpu3dOBzDwrN7yKfHBNiOB1MFlxr56F9Bqd6W/XPSOhE5swMy9rfBv1RQ2O3ks5AOQv7sXB3zv1
GQN+tgXu8Cyzm8kKwtDoWf50xAf3XH4AN9H7hynpoqIBYFmvkRcAJJQmZTdofJn0vVlonIbxOnxp
HiQhioJt4QT6AVwg9Q0+6f4nO4NpwNh/lV7ULYoRE+zRwXs4ByKdb8g1a8JWK9zhKmrCUCY3lKDy
HvwCo0yYcz7Gc0bm3Y3hEGWn5NfCW6frkZW5byNupJBZEWaVr3juMAOJbVjM44AoR+mh5TV4YTUd
iot/5l4DJk3tSYgyNoHmxMWIkXqKXUrqtyAFqw75k54s98TnguKIWlzEG7mNpcuJIhluqbirwZRg
4EIBvoBUA+nJ0wqBrMkmppQkpDjqYKJfuSwyzOphVFjcchMyOo+R6E4/1aeb/A6xCYunxRi8cwMl
ZnJXf6Z0ewlmvNvlEgZVM8Cdu/StxFOQEqi20CO856JQjlDmooFCsvXtonmj8gtNEqVvP33/pd0j
8OW1hmMDdzD+UBCEOY/T0spEB9cmFOE07Bd10uIlam1EpMSzhTlzxC4W5lR1ljkHw8/0a4D2zTlG
/VcDnUdqWYBaaLqDfsq54EKLyiA50mu0HA5pjcFALHCpaVgleuhi9+VskNiENvJAyYLmSCkKmI0A
qgf9rsO3oOHAhqGxl6SmOc4r5rTwgCjK7DsEpaqGbtzgExt9NWIQ/mdSjNW/5q31ZmU/p/wfB9/E
EXHjZz+By536il+/s27tyjAVtFcmmFPdv1TvvQNLhs6lpIIgq16S6aO1+Mz0Su7sLO25gNoEF0LA
rKvVE/52+dnVjK7B88utFJGEQZZyV62qcysP+qsh8dpkXwBWj0GHAsntICI61x1oRsYTIFEq+MUG
qQqlWf7eBEnXqkYvpP/Pjd7iNl6ibV3aXDnXh5qAl46+GtHrg3U/O+wo1ZCB/6D21sc8RCizV28w
7pqH856JMr+wY5zftYmCniU5TS+leM5lKgKaf8RQKFvGFNvfBcOBZ3ZHGLlwXAnjSFTJTYbxrMt6
vXKLjVGUlI1JjzihJYd0Kr8VnB5NfMEq+PAtmrFmPQiRJTfvFJsmzYnrmwwblY9pBrZc6PNb7YXO
YGrdtlR1Pv1ZtNwUXh4k5V/TCqhvjmrS2ULqVEUAfqtqhqZHNH0ocKGPieJbBOQe4jUemGnHT6Na
VCO/UlUeFF4LywRsac0ytxnmSDytk1JV0JiIHw0nSjuRsL+4LUbTht/oDMotX/e9qquEA5M99QAZ
wJrKD8GWP0HfAIRgalIp4e0Hll5TbNriNpwTo6HBixaJ6VpOwzryIxJ7iJv575HiYx78VMRmgn9T
0Zax15Wsn9Qrzfyf51I6VEESqYQlXdrP1FVEoIY5ceOTk03dsPN0ydcId22xzIePFYQQXlERY4Nn
WxIFXPovsB9K4RHA0L418UaZSsVlK07J94tulC1ubMDM9TQn2K0hWOLLvUdtPeGNxFW/7nKDJyja
S250Iij+3SOlKJN8lFdrSr8UnvD4gI95TovLv0zn1/Y4zZQsvkRtOn3ZRGhC/TPhVMGRHhF1E6Fj
1b8Y6wX22Da992NhyE987JzGdLAsIb0t5ZPgdC4gfPSaXBxoNJSxbGS60K0YxH/iHU04iYbDIUia
7c2F8JGCPH1MgnoBQORZ1oBrrTLy4u1YRu1b44guXmVxzvPOKbc/ltHFxFZgw8uXrhCkCqjcua25
aqgkAihFI7gLS+7HbsSqUrKyc/MOIs+x550BIgRJ8lItoiVVa7jpKXPnpzwl4H/ooDtFSlXp3QFP
nd/4hz0fKMbiL/9oyaLSvDpfelgWPJs1kOEswxDbQAyvBbhLOE1Yt/rcSItwau0wYDrfXv6g5AMd
IBougw5i9JUwOAni9SIyJVy62ahWgI0LnJGICUI19csPwE/CWo4IL+mj3rbwLgIcAXUu4cqBTHMH
WIhbLwP9v6bpRoTOK5wxAD7zj48krnpUoJunOCQDZopM67t3ORdcGq+qu7qMOJMQTur7otWL5Rlt
o2pfrjCv4xbNJymPySprnAplaJKp934W+nw2djf1a4zrGn/bkwMWHR2XSou83jJRbwCIK/xjj7aZ
zXQ6ISNJwicC4b/caONarLOmibutciilA4dJGqoy7ST6HiANCqUf26IqC2TVRfgaTW/TQFwG2ajM
my6EXJ3p/VlSI9jO/Zsdrips3O2JxwtJzk+rzgxC2PHjzskCDsPgVXnuIadoKwFyfwtj2HjpHSAM
nNCzmygOIkJ6HyElaM5ZBrYOvYM0UBF79d/N3fYCLTNhLHG/0xbFOTGOZa3nsuQcHVr6Z0U/nf12
DIpleXbYxau8Tseq4A3tdWT6cjzdTDo3UZkD4DD9BC/YZsm7A3io/0zTPwi9qLPSMXtQHeYxA8gX
zPPHyoGgFHyvnDhyEJwJ0t3/oVndPYczoso6fFzq0LqkKaq9LwJdLKgfw2fdptJvdHs4sEpghMzH
b5GnOMf4AYs91Bzl29vw1pzwYyDqgGcmwoh2fkx+Jbo33JKkakeojzUUAPQ6blIcbwy0fKSTynKJ
DVjXxy7EBagkz9fzbTSU8pWXW2R6KO4zGbFIFs0p9n4IIKw5yEnO98TxBwvu20HGVMWCjA4HUHbj
qvRn7IjgulsAYKD4OhjfQHQrIClvYpfRFQMMlx5alRuGrP8hGdTDl0p5gQyycSqTkkt6+iVyvC1I
2/zdnRCAe63DgvL+gwCCMYOZKQ2jIsWrkuBScvqJT4OESR6lD+n9TWnJFP1ljruan6+xkitxTHYz
XqMeJgBQD/Qay1SXqw6+xDGUATtG0jtVCnpyTdNZHhfWcNUHWjDYGgyIpvfDU4ZFT7rGWDfzUfzX
Ol0g/2arUze+/FCsiSdxUChNaFrj8zuHK9smh6m8X6mhTTSIW+ddJ2dqAPh3lFkDHA8aIX/jyEeV
6jTJg30TI7pP+i3Tv9gdwXBstmViOZTQ0c8LZuxyLMQgQUBw+kOwRkQ/ohqvIVS/Go5RaA4AWUHo
dXYzM0YWk/kM0MtJ3ud/K0XnCvyOVJt5wSahfuNf1n3770zYrCY0mmzu8OdX04EsSzzGFG4ReSrI
3IAb82NYGoIJm/DOFAE8S0I5B9bG2VGi8V1MvAmfq4FUc2T2KsqjGO5fiAyv+4yewHAr6mNzNjnQ
x9PES0LAOT84MPwBp+A5mP5sh+tmHu3Qe+4Dj24bR2s7/G3r+WrRTA2wO8mSa+Nq7ldP2KC+AOQ9
WB3OrsphtwQrg5o6ZlF7sE1q95MRybAXaIGUwA5ywdr4ouLSdij/3U/EnhJlcxfovklMy1xDB5qp
OVULdY4ECEhZvH2nfXCTC+NcC+1cFDZNAx5Nn1F67u7AHJ4O6knydr0xN2/u5A0uwROkpCEpf/nG
JkbbZlvofYRe1+aL4Pvcy3cqCDgDiJOol5/SPguzsMpaoCnaqaqGRaCS+m7fqfuSAJGvLvL/sqbY
LMavo9R1gVnllS2MnaEh2h/IVQw6llylzH3gS1VyEI9WlhZ6EPMqG98DE0hBj2tzuTMByUrYVLsB
CYSS7HPTqdoydyNForZr2iEoADhM0W9dHGHY0BYC8zqWvgXMHu6/PdoXkrhy0pYpO/4aXkiibA/w
q3igBoulLb06QY+Mc6VOQCyE47hxMwmMXD2kZzCiCzTDQxLBffMOcfyehvExIO80XIB0YuT8rje/
afti4LwsZ9L9slwHwma99JZeQ7zIFoIzM3bJTYF/7o9KeCrake2O3CRG8qxQdn94930kULTAqxot
oG80j5IHTxUJRVdcfWCJZwsoF24bCMdQ+QuU95oNZJC27qPiW6+Aw2I+fXb+z9fUZY7L42lzPJJw
hPYNOfbn8ti6GXAYwFlghNEci+4Ex/WpnOe6eDhLpPtyaQsswU4ZDQPLXz0hkSqUtuukEU9228WP
HhOrgT+fWbe8Z+cxNofFUhv7y+h+xj0Qwcx7kAzDtftfsiQhBWjPNu784hxFuXVnms+iCiN+c/nU
iITNPfhRYnXrBLBTq7uh32XVJcUHqqSTt8r39qD2MtdlR/+uwhfQG9nafcMGLmmBgPiRwNXkPliT
9Dg48SgEH+tkh0+7CktmlkAXWtl1uZ2AHrXWLGMJYcOtRKAZ+BWe0I5xXjla1Uv8Qb3GUuCatrBR
BoOL62bmYkoxaS7i44X9zeTYFgKRzE9izis/RzpEECofWkoR/CoO1FQB644i6S1kLcX9Nd5a9s3c
pKiottNze35PQLMw9jQo24FdEc10sT4sYqCDMTjTyThRRbLIT0aZRFoV+oLDa2FsG+WglMmpZ/1l
lSKn4NalN2M0GYZeYOUA4ukHtkSyYzd8t/y46JYkal5pi5vzG1uzNfokzLKlFxQuVYk3vTEaYlQR
XvTJKcx1C9BmtkfdCSuaI4xGFYvQsT+xidy+4uMyPAX/ss8qJuwrYiV0aOz631DyllpHroDWCwsY
CwjmJXY+ZN1IzOlh687f38qFt83OMopnWETbCiqzdFBSFbmP9Wt8UOQmAjevHDFATD4zzgFryy+n
VqY6F3c/luhfbssPjJ6Q8fasVGknkWqlsN+TRZ4dciB0pGXvKW/x5q3kYF9v73Sr4LYoDYFAZ3Hn
0SmFNggAGbhdeBTd4889Pxs6A8FAB8p8dI0FUt7vyhNOdjqU/ILSA7pHic76MOGraztDOTqHzCT8
fYv/4ChY7Oho3gcyWtQj3lf66NT0xgoPm1gwVnzT+WcJ3RzZEurPOn27xWYufiiISfJN2zPeVk42
oYaktcbWwLTJXb4ZUjYRHa66oGk8kRhYZfEpD4ouayIYB74zkyNMJGGfG6Py9qh92FqWJ8DAdBXH
CheQjujpWt/1AxlguiTgHyZcshXGUKtVBnG/rFf1lIReaOlALNqpbTMAssvOuoohgG3WnCK44ch0
2kyYKUnfmp4wSSlEbI2QXIppsNA2DXBCDlg1tLobtuXTYPj6lzx4gKx229Ah8qcmeHlBgn+0ZF7A
sNnJNb464S65ysAFlILe8JfdhhoALpW1xo778EKZ0t+GTEoKtt1cKfJEk5mcQgE6ynjBnhXJt1UK
uZZGIazQwOJCPt9lgb45TUmM6N2zmMUf01mxUoOObU2U+SMAdqvBYOYxV/gJm9Uol7m5nrRUMmnq
SRnAzIfwgVGLsaSzO1iNWSLjAKkYMiibTAu3iBh0gFIBjFDIbPrEs7Kkk9H05bNqi876vQ4oTmWJ
bLy8LH3qFb4l25OvXwsnHTBmbpluuGxBTuw54FDFWYnfKJ/psGspMOYvvZLioKfMWtd6y6mlKj+/
4VX2DIipuCrMdtUiGJIVr48otB/4zJwtKYO0EQUCW7o6kEMtUcT3KnqxPEu3qOmFX9tIDNCaTY/9
FRer906eQ7TKHeD6x5y6JYwp22DUmbd0gX9+zHfmX9FcylJtAlx6n9zniPmVya3TddcaF73//u46
BpCAY5F8rU2A1+qE1pxSxVcWb5Ww2MEBzFpv0VRRLpwxxYOLUVTGQC5jTV6smE9dlgcoYkixAnAS
/1bilSf8eoh4RD9KLfrxx1LCW51MdS52SvVlOIho0IZ44uytBKkvFeG0RtBsxe1U3Pbvlp+yTlTc
Kn1qLmgFiQ4v7DhB3qsl6q2C7ppEi7sXJm+dHFdFjFXdYSTYOtPLO+8K16xmzLHCRrBZjzMhBErc
V0uVcMrjQHuPtl4mDKKvzTqXGnU7Ii5JeEg7+8VEW3jmj2Rpn5xnJuqikLdRbJzhGnMQB8yfwwoc
Myf2uwd7jUyI0yQ8OOR47dXDycr6vWTtYrUMEsRvs1uNb8yaS3ITIOJKVypu4MmQu9GSKvz2v3/Y
2s4xNQaEByqN7XAw7SL6hHl7GfVm+ah+IZb0ciC6PUG8huHlAFF/B/99qFDSmPS5I/ITFZWTC0xP
+gG3jypyYrpNxlhM/kd9udtIe594YhCHUcnxx5oCtEQ7fWL40HECYo5oUo98ZwVz+SSB83/29imb
VCnwRPa6m97kcQRWHNk3D6mzvu1drlo0bq5DklGlTPO+wQafwWykmvWNwEs+TatP7RZwRwV/ATTT
2Nla40oOK29hn6AEWF5RqzfNqyHsNoL4eXplpGVgod60Zsgt1acforfIha8TyfuL+UGkGw1HScqp
qHDhc1lEQLAE7UFxdRnR4+hVLdKhZ8TNhglupYBO8fdGR9F6j38YXji7bTqclmtHhPU2mM3D/iK/
F8w4gyHYb57OUm60tuCkv/Dgf4EmszPx+89GdraxPhMXExlTzXCRd5gp4fw2uEHxPH6yVRCnQlXq
Qd1Nho/6LqKA7bxjNbxFmOWxTpaXjXIkyqzEAnIyDq4fwofBQUE/JzPpzJ+ADdUE5nzYY48fHOVs
mJHr4i0ZxnuLJcDdGeI0fRtquOn40Vn56/jAmzi138JVZfX7VenL2XTyk9jrTeDp3i4u7BcwCl+H
5DKPL+yK/FvzUyaLcf4wFggcCkn3hIM+IBO8D7ZTGrdhfq7C/asyDIVSYmlT1k2NmhlbR6gLZDBA
BFf7rO1lqVXI0f/1wqy0JhulfVsDC8qQsTPWRKccyLE9e1/5QFIs3p/ralV0E+grCjV9sjS1iBzp
2oy9J0VPMQWhwBZu8ZW+ZSQwxagPOqKR2RSOrNFgOLezMjNGI3XcPoxKJI9L9mDPxmAcIC2yV26U
trpiEuYdpi/+HqbOCnewmkEi3+JctRKqF0QH9+aiKPqiajSAeJttO64Gmc4al0VcgUk8RnQWWH0j
1FZ4Ca4aOdBXp9xdT4GmiHqHJeWgB+0u1+JxIhwF5FrUzNzRhZqBPLPzfrHSt0Vs3idkquysnRqQ
5I7yUZycgRXI3tP5nULDtt3vatKdvfsz3MH767FtGkSd7PclxgSYcFSGYXWBvCPsFdFch8MTwIJV
h9jA/Kimcwe1/YDmBaY5DEvuu+Bc7XnDmxMw9LLb8MmmRkOkO+hJoJEUAhcRk1V6+g5c8UGL5Hmb
62f7v/dubkcf5QkE3BVvvId54hMf6b5t+eY/H42gASRTQod58SmBwpZXyakTnqXw0IMp3gp7uio1
bm98vfB7PA2oX6eNNu5GrC12QDXHfyctJRwr9vCuyW/JnLYSvTEz0lRkUw1ny1BzpMhHinIbUpbL
HkYtLFtKLG5K5Tw3oCDc1mnanUBNwoxGgbrY/6PGVcJgeGLnfOtoBJXMrm8hQbtVuG4whQLaFWlx
DiNW1ccjT1Tb8vV5Fb73NuwMUnwOc1Dqo27zh6AkLAh/X+45JkGaYNHOvy2HamOe5D1+r+cwiElQ
B7SB+hUE4QD3sWiE5DMx0ulDItWC5zmBDSbho5D9pBZXSZ7c/47bwR36xiv4G19TnR6EoZ1KssDw
F2Tk2Nb6JICZY0/zuS/mJ4tC7sSzvP3M++7HvGvnV/TSOZAhIRVe39UXdeIaeI8dxMymdarOZS/J
rczlT8pGwEpLA8E42KBowUt6XKXx4dmc73dYvTKzBOOrues/kMGqX9YaFCDtm0J9EBIvtNqAlHrU
zQUGk5d+fKoAXXO/opTQnovFoQdfceUpIKUuE+Z4CYLRDcFjppKIZaA/JSwYAhejRkjm3nv1OzYa
RtETAXSbYuoPVsQfl+j99q5QTuzCSgVt9sJwIPGpW4LrdBe6GrwIfUQMTZNK4r3OpG2ZcxHpluCc
2PNL4MnRaW7wPv6TnIAbDKUSnLZWUeBsS3HH2ZuI9vh+yGfZAiveDgbZR0Qo7JqrADnABJ9xI6Ve
6tjNYUiijc3NuyOIhiBo4bhx2GEzliCX7heL3egRO6WgwRto9BTV4pzCDV18F0O3mZo+sBoAEBCo
dmbpjUnEGSA5+slzKmJwYIkIl3O/d7CYDPWK9DuPdNp1dqakbSJsEHLC6WH0lHbr1+Zfy6y+AxiI
JtTjZRAtj9dP3UF6/gBuDplIqBjhQPoKfPGOYGjpTrjsaX7bdki0KdMJKaRAl0z1r67fwS8VBdyV
+Yw5/i0H1yhXnqlIXllyLAWWLYBGR1rxg+49QA+Klm4Fh+nJqBi3It6JDIDqqNUgTRXkycjn5FRY
jXKKmgnDvh6i0q4vCRiRHy5cozuo4tTS7JzVpfIO5SK1Hjkusy8+ntgzGcHCb9VfEluy+BN/xkSE
uLAoAhYhTlUb3LeHY/WswD8jAg3gIc463vVL1Gwr+wiPzSzON6go9eyk7sa2nZgX4zKMZ1LfzNsY
0yUBHM4C++6W3lo7u3uR90kEgXXLqQGRST3WmN0jmnMXrCGhWJZp39CcapffA8pG2F8/jshZO6uV
WnLV7BylAOLBSjtrRI3QSKwgoDEXqv6G5MeHhEIxkgeom4Poyj6WfjuY1jDVHQuFeneCCAigOJs/
9XjqWTuwB9f72vXDF7HFg4mLP974/YkIQxwBVUXD2DYLMn+WrDr7/ZaxXRocBOy1H2NWZHVT+lrF
sYWp3LLkefvSU5obWiSYd8rQBdYVn2v9DUL1SpGVd63cL7gG2dC30Vo/yVmOOktgui2Q0RL1I9CX
qk2vgCsLvs+N3ILESW9t9WwdB6L4ArBhxlk/Xo4NgBYyYqE8DoXoIvG7EUGGxM4rtA6rY0z6tR+l
Wk5IGVEMMPywhDPrIuu4iBRd//tWrvstv4AQz3nOoWON1Z5VtHKfL0LkDcWvkZms1Lwat5FgmSyT
eb9h3zXszZ3J+VGNafnO4ATr5jN0JkScFngknNRBQl9min5hVnNxjRgh676pih2vrfVdvsN51NEg
V+XFMjXpCioPJOcOYUlhT7vSYwtH/ae0Pf7EVfWwUen8mhVjk3gcuGVu7tifhIhpggBiTidUxi4F
ThpI9uj01vdlbZ+mfRw4076OhPXKjyDQHoFhcTJIiqkjEUiK16c+AOb2k/bwHG7fZtzKsZqFiSPs
lnoHE4v2Dbzc5y0kVfLs6p+doPA5uJ83IW7QSBzUaG0Oj82UAAUEdzbGyu1M+7RJK9leMekOt4+K
OemVHq9CZhGGlrIv4y2XRq7GwgrDTBWEkJYXcZOpuVG0i++UD7/FCEwK3Y5UnrJbJ6NtHjT1H6k3
y9fWz8pg7Pqylgh1wKXEFGdqAa0OHiXLwiqYHiR1FlU3NhLo8edpWl9ggea6lWQ/046A1SIwfoIw
lRA6XJxLRQENCyJMjrE0/wy3BBvFuv45nR8VwwEhP/gElOuCz65r3Iz0SwIN86BEdswPBSXApbmJ
YU4KISWjS8H8mHzhrza3J7nT+uwHLFPpkoRE1H2GvIAGVb96Bn6Nb8/9kgTbv3FEgNQL3/Odf0Qk
qeg+NwNu/8gomDadorMG2Cr6WHZCgZ+P9/Gjjj4NG1xjlTmWVtXKWte7Fb8u16VmxXh6uJoAYj+b
5POGuDyWJYTTyxrp1NhhL4fJfC9Vf0M3SY9WTI9HTkAEs8M7jrpZ497Te1JpMHlBMxQv4cWmJwnh
eXauyfoWKrBK+zr3sCXuOXSfMqvvHE4cqp0thu/AEQOmkB5EwpBKhSWheoOs48UcZilqcAH+oTHD
rEILgb48NrUyzpsp0v0lAXN+Q1Xg15opdnCfC/jDBdvuu8A6aSa+OLTurZmubR+v1E02tTXmQjAq
q7y06un+Xl5NSv2O8vDmOjd+DraCYkoiZNnfiz3iKTfdkvOl/tvY/63/I0f0qmrdichwYj5oCEej
cWR4vQsSZXAnDHj/N8/j2JKBDqNtOk7l0VcKaiz2YWFfR5QI9aDuFZt7XBBVJAYed1HSkNCKjm4K
2/PFMPvE1nxUKqNtwzNxNIcpUUK390pm3DYtNWb1VdxIvYQ0dhbOLpWjd+NGZEx9F7uti7yXT+9z
DyZ/zMtpMMADEmVDiZaISaZT7Iek7CVUChCGGWzhJ3e9EjD8xOrrfNXuNVVdI72tqqCOesIqdi4d
NDrSrTx7e+vXbWvm1fTr675Zc/8mofmpEIC+o1xFToEVwPaRFvYRVsvyxO2N7kgN1uwHk2CLXLD+
162IVeyo0nQot53jrjLBfAnSTNk/KscBls1/j9qm4OcdapjoME7BgJDz0QwYj2+3337DYQbJQegv
27Q7xMq3qAjlPiMSwRzobj93PLiKU6hU08DroJd9LeakGmxIKa1SsM22UAoJSnvD1lDMxRzjcHhb
Sh3tt0iQ9nR5rOJj4UoS3RbGFIcZGcMMgChCYeu78EAY8gWvW38HESLmNT9InfUxUR5Z1uNDCxCI
u0lNZYZHOCJNcpUUR3GfwFNymu11lqneAyCYSW6SvIMFDlZOadU8FM6MGK6uu9+t9SJC0Csip/0u
97OlsO2W94zfI2NJ9nU6GYwQHFYKSBO/bHFsX53OqdWbBJpB6F6+3zBi1a0ROfezf9Z+gZHsGAar
I6u3y8Sh+W+yE7qfRFy9aT7hrMF1+Shr8OdC/2dltjlE7OOAs1UQq+82CkGV3MWhvjfhCZYPwAF/
oAxExE2kH8AZlc+ersmkReJZh+R+0wDfMhMWYCH2Sv1s7tIQ6ZndiksvtGVSywoxCoQnV4PqotYt
hQIAQLEMnu7dJwA1s3vH2/ECbiQoBhzc4KR9HDwf0bGsdstGmXlFWe8cxK579S/etiDIrmk8yX6X
EhuTXlCJlGE/NF2suskh4ptt0/J1KLDjQuFHMlT9yvk0czPhdg4oF04UJA0KN286fFWQtucPosIn
g/WHjf/EJWvpJVCbQT05vdJCjPDbvtyqsnB96GO0HIEoTkHyKpB1t16qLuLGdTVIu/kUJGLTePa1
G9panKXaBxglf7q7MXZJ9dfZTeCuo8yYVWxrmXfw68rPS4jpbkY3xAOstrXiiPBmuCP6wTCi2ayF
CmQaTmfuGtQVELqjEkwbCex/hqnVMvhUPW+u/UQv+p2i+7/Fx9Aj4rzasBGrqYQiS5wi8D6D7Y2+
rZCDhN57S6cN3+eCJ2msi2T4Ev6FiUhU8ioap9i4/8M9EaIAQWRmS46j1L2EOgRW4UBkdqJpsL8o
Cl9xCpmNmPeBhSIzho2gQQCj4TUEFgOTaIeaWqwDstqAgwPgqnkvqoQi8DEvR+SvwL/ID7+k+4hy
7BpYZy3m+N+rI0Svvn+m16a42eF633BZuhceLR0ijSzIfZ42B0sAqrmIEBYTLlapgH/95smCJYPm
01A2p0JtgPcVBkGORXTamjsxfwqulvQ5bl5h8L5YyYM9CesbS31qefpSS0XXYEQdJzGdL6QQpWuN
/6XEcAxGAxID7toG65YUGrnqSCcLX8SVYIhPRIMmU+Xa4O5ihSu7xxnsQ5G/a27SS2tciNYBpKPK
Y8wwEp+bPyg9Jq1L2+AgxlZw38ztDa4V4RFh5RPLttLXJh094DTIEroCn9OfXKmKWv8aDA1H8Zw3
zJk8r2WgZ7kzGi4LQJmTypnuMvpgwSXcKORRUCTETk2sA08MGOj2azm6TUtQ2MOvLZ+SPg/HsQ9d
u+3M2tizU5ClZjenLOMIHv9N+KTbiwgx61XM3A5gyQCluJTZ3l3/oDhe7iPeN3R1WnZugvs3u6JF
RPTVOMZcjoDj/iAABOGoZsToN/wr+CqXrpsCy20WYlQUGFEQnjCjck5slN9kzTyGJQfEBm7G0nPf
rE6MiZ4pQ5F0hDMimQNS6ay3EysceRHARgR2ZyBgY+iKzfIvx5U6/cv3+PvnpgUXhoY3SVoQw8FI
BEc4kcbMD8pdA7wChfasJodS+zl33bab0mJOIkUB3NgOPKgoGJEGYR6j36ErqsjPNf2hdJ+F5DX2
6MBl4Uns0Rm34frFq6YzMBjt2PmGTW+JKiN09J0TXTJ8SFlwz6fiEpbzGpIzwlgjMCdqsooEuPpg
/Ayam8WRTOM2WWlipo9RCcboSPcBQn/FDCyDwL6z1iRSwwypd9ehPV4Zlj2dbTWeMowLJUsGR+B0
0m+P+mhIAhhXNbobQ3xvRt8tblvGL3E7ToREuM6gUn6bhPL9Wq7hjqLhEvszXBptq4jgIf/p7BGT
WRbgiXXp/8QxJgiCITnqROi/0H+Rain/2+g5oIkz4xNLNYpmLXJUzB3eGeYGMcS2XDPM3v6zKa8R
AXLVG8PRUYgEnfvtpXcsua7ypsZjPzumxn8ZBxUEboGxGNplYm3OtCkIHIOjkoY7FIrd417ltZFs
40WWSrL1sCz4pMdmaq4kyepEGvpvYajji9rVvK8HH6rMgKYV2ohItok4dayDTHIEgXQJ0tU6GAXS
9EG2CP/5o4+FXP3DL9mPb/hya5+WaY7J2YKUKwP56sHW3XBEICgmAYcB+RPsP9OgzEENhy86PWdz
GkOJ17fF2sXYHCbqG0EgHsVX+Orw9qctKl/jbfAMAti6SwZEzyov2RfqxFdUQ6J5dnhnttnOK6Nt
9aDDhcdS5lmIAN2yII0RxHhPJ7wqc/LDw/8eap/G+qSGqxZ03Br9VUzKjLX+rFn4536ElfFR2IsT
pEXny9/u65P9Ck+fPzqvs+1w9/n/FiN2X/fqzv94CB7Sn3olxv8bIwQNrDf+6Idz6tWtPSSYKpW5
CteIYeqkyARLQdj9tc1B9wKinDny6UmQBN07KRRgJB8xgjg2vKHHAJse88RVMQhPeoB0I79DPlf+
3EwbtxQnuVzfbtlxkoJIftai+ALMhYiU2NuElaGCSg5bzWlrONzZkMWKFUZa11QLQbT4TM14xnNI
bG5gSHJ7BxOPnjdvaPQjsX6YCoS2wGM7+ngpiQZ1l0sVjHWEQQ5N0xmss76g1SVgxEq5XCsj3WgQ
PwbzroLkx/AWo4zuAGHBqnB9y2AQ+deUHKVJjarU7E5BMP+1AoKlYghHdMaGbMOVHME8MWQyGqh1
F1steFMO/kA0YL0Fvf0jpN1vkFwpUp2rgZliBHL4HZR2Y7RsRdWI4MFU1tpFka+y6kB1PKITB6T1
Nl1kZ1HvzRE55M+VAkqSuUjSXVOfE+rVKeZfSze7H7NhNY16Q8g6dHazwMiO6umPr3PFJR/bLEQd
pk/15LJSlqHR4bFN47CVEXV6VhfXGIB5x9BEJXhSBUKidUpFNu2Nhf19pb9G8f00sDnMkpUZrduO
eoKorR+oUoMxHgI9hyYELatHpS6huHYDEhhIJM7ojHPTTnZzT3dJ61y1DhEnILYCzwsVp7LxeJda
1R7idt7e9xVSeE41PJkr4a396z333F+ZqjcJ99dZJMy79quuQvtI6srEJd+JmkoxoavjDmOcS13t
kXAzhjGzomUkLGS1eoiA65DvGIM699F7X/b5KFBzu+DKtkml7oHFFG0oWViyxSgAWLeincuOOO1/
lKECvfzDHHWGSnFHrYuDncMbBx0Sof52Bgq6dV+Jja+NHAViW6a+EZKGoxiKyP8jqwaZTa9guoNZ
sjtHdff52TZHPEeymMa5zPkQZh+XOSJFeD8OUUFyhHbXE9fdBvOzFIlhIZczZE0ytOlZRqKjhBEw
wl7in4Pgs2u0SSrznPAh71phkYR8DWepEpFxzzgAARLuBa2sAt+Evm06sbfVwlYAiI96fhbzAjO0
d/OEJApj13InOXo9iOiFGOk0a/yKcNA311+UftPUtoU0zoNNTom9gEuZsPS4EwUq7G52MvUP8lh1
LJ+8XY+r6ix5ZaIFZHETnI6m25L0VBk9gr874Z4OzPj2Uq5oV7F9zEql4chKtAfnInkGlKlOWsaA
C7jRK+cAKQzgcFaqZx85GRlQzrzu62u+M5A6Bc8cCzQ1CFUSgxVlDT3XXvRGvPjngcYDct7vgL6Q
Rou/zX49KSRycH9gaOVqC8TiKl7ne0UenLO79lxJkm/yiiibl4j42k6fsBHbU1EcgiPcsTPltxaq
CdzSV3eT8O6cagHOnbygu5HBwmVESgVzP7pa6Ep97o3TeCa+GQ0evVh1825sBil7XXMLEgu5+0iI
PVZHYOxCzaJxc0pct3bZ0fv02gVALmjpvKzgFTmJeV5PlH0eQS1lPYHEzwr6hZ/fhde362lvZA2o
9FiZlTKjOAZesvPvBJEQYMP0Vg33yJZw1+loTMUKo4Do4XRST74tHr07PsM0QXqZnKDTm5V24OzE
F6Zofp3I+DoD3jWj2iNh+OzQu6pSssjUv35YkTb63iBQoshILB3qfer49iJSVxIvJacQUxwaMNbm
1YgRF2YE98eYEmNxOaPGQIgiR5S8FNEBP74G0tdLl5oftP67RPPRHoOA4UungY75npoFZ1BuIIQT
i+NVkQcM9q2H67NA0eOBitwCXpQPvbW+nLEY+l2ZubvN8O7GKkTEc1eJHBHN5sF3Ju1ugtdOu8w7
20LhfOD9Fx/aNvaBTZsL2rIufTz2yAcol1cmRlbXpGKRritHYX60Kr/qd7do1X9C24yi5dh4xSV5
4L9SromYIMaYL3CASzq8dBJmI4Xps+BLkFMMAkLcq0XBgGBsf2Nm0oWeQFuJmLl/L+STdyhXPASQ
wQ8JAUrhWBuw5gz3d00JiFCxFBAdQYo88ezxihpX9/OpY9yHcHlNHwK0KLzor5GVobXiQB8XXq2s
RzHPDOAYCasV2g7TUKImPksZsotIZj97syZjrEh5KmZepNnx3PatVQOFOhtbfwwj5oHasvbEt3u6
Q9iv5zEkVuEDHnjbZ3BYMdzdTHJW2TZ+cYjMWcp+Ai2/LaBeu7UsFXmMdcsj4VxxgsgmdBMdkfZF
VxotsR8z8vEMjS85XshpcoU11dJcT7jTP5JYuMTwOs8rIcX/xrNvo/Ww8zcaukgJ9BNtM/e2mPUV
nhu+jjwmLtYEuR4EDAlXL1zkbPH8hvCTPMW1gTngCd0EWTmWZN/VZhHU/oeuzCxF992CslHjIBIe
oA288XlqGaYuC+P8J8pWj72PxE3WNzBEB2eTqcULundHfqWKIlIXLdpb1eixi0mMcbGo1o8Wg1EV
5XVZ3Sitym/kCOCZwgHxB3Nef+V+Ls6ZVfGtxio4Fp3FnQ+tAJsMCaptLTo4/qx9essgOena9tIt
9ecKdoIbYMI4GvdV5LSFwRJEu58p1sTdsqURYVqwQjxPfvKGNNRXt3SzDojKgErb+0dTLf3YuA1a
nqrfG4YxnGm+p+Yy3rvhBkgdvQl8P03+uRMzUGSt5EwNqVeAc5gawyS0DobRUWG7paC7vRT3GNMJ
Vvjlxr4q9BUKpjzNDOeX8krehKhG5SLt/ZJGua6Yu3yZj7CYrh2uJKeI0oHDYsxRK6RYoFOen7Hv
2ioHPwyaZ8HyZpBgAr2E//pEKIvFxl3OItMNSdarHIiw1A1B0TA61b9ZcgAbZxNs6Ur6OVwjoeX+
uA+elkasqQJ1qRAkpGgfJbtEhfzfJt630DTSYcPCgMHACOvsOmuuNC2Jwz3wbSi/v1oBDi+hGThU
MmoUj/6+NSI5erqFhAUiZz0btRkmEJWt7zVYxcxYrDA0CzIW3sgGuDXK3INtoZFiYZNG1+al83P8
gMS/D0c22Tb8rrE8F8h2QdFKYXYdAAkmN93yOLaMfgPj+YM5F2ilAgmrzPsgXNv+D+ducw2LFdKd
a0CrwsCloknoVTWbk8AOrDmvS2K2znUisvu7jKagZyjEiLg95PbaZW9x1qFGKl9q/cu1fx18mzn7
L5fynS9Ioz6QH9AemFxjBR7d95/dSvt0vkG4Z3ikFJsQfw98+88LizHAaUjXhQRSOw+HUBAlPP6L
wErzJXBTgCkM6TW5fF8jluoG48EXCtNMj+AHFyvGWpENfj4tZupIIhZ2rJ3dx896iF31sIyDmvKK
hP1ARha8dh8TMQlVd0bItlhcSVsorh2HZj6z791kKqh2gVV4dCRrO+HD1G90bMQ1bPs7kLzfp+f1
+tmTmOXs6foKDTGsJW/EoPQ6wYXGSkYgJvcP6xRB0XutrJDU+QHYQUtYTQJa0L1YuWWU0+EyQj5K
nTv0jUmeONdLAitthCNCMEbhiTmsgwH7VM8sQmzT1NQdzB/t2KN+kwOHCrnyJQJhBm9R4e+vnOGw
lM6ZmYFYVAOzwZ3M06QyXMkVdL/k8nmBaAzADjK0hMWuGLT8bbOnMJvoDYP3eB68c9IpZlnGfbbX
UH4pvLQZj1AdXvsyhQZDHkq8Pzo3EAvg34n2D4NXI9/eMozh0u0l72NunlLgHbWQuIYRxNVrPZdZ
kLOjIQGi9BPShsEuJWjcNrnV536o7bAzGMFmtv4fnfeQOtBdION0J+InUMg6+fRAaV3bBgkc4kE0
xyaVURZg6bnmQI7nNvFMcPIvgZrxANyA0NdjG3NCaVF8mT+GlFW4J8aU1pBPf4mXXzGSB13bxWoa
gNLUMCoZZjZNbA7ysvXD+ZSDRPIQxoH7sPyg8QY93cyvGiKnbAV/vVpSDxzIP3/DaJlnQCnhHxP+
TIotTywX7jx2faeO5PN8bK1J8Jr6Z+/e/p2PNovBz8i/TLfjDmB43e8YsZOi5isOvAQeS97vk6vk
/4IlHiIGWy032hgtL/idhbD26uS2gEIWYP7QmCIWaP+NSusmoeGcu5gW2QaCqbXkYdaipEi+dMlb
E4ezwZBEW1xeVZUWLcLiWoTRR8ZK7OUP+pcTyeDKTYrYKC7Qpz38sH5B7Oq9cd6824Kgk9vJVn26
N8qWHQ3REKIpRmCk2tM7UOG9oaUAsL0YPqwtY127W1QOvwolsHHi+2ycQTVMmslPZyhQauK0znmm
DKdQWo3F8Xwy5oGlCxnYnkGFBgM04OraRx1rMQgzC5zy6Ml9ZBCl2v93qYBZvULLASTErtnSznbn
tY1u6pQ+wcdUNleepBoUTkMpLj3b6NlqvCzK5e1Q5agJSMQ+7HzO5ZztbNDIRl2gtMM7WMfwCxDS
q2hx2TYmIMp3qONiFwQnD5VuCoZThxJlV/JgtBdNwdqSnY+aQDwve7I8ZsQJPV6/ZXGgM/hV1MLF
1COGYjZRRVWEjPxU37q2gmJw3UJGmGPEgXNrCGLuicSczy8I66dUlnBQU6i86xhcZtWvR2p3FQxk
EY22rhLnm6w+xXar1Twoglf2IxaZVYYiREim5e/WllkPjCHWtzfueUM3rYRNTfb8BkNzuXkFBZhJ
e3g8Vj31G0AwxC6weyCTKIapJEKYwP7jPvHOampQ8eFAlP9VVQD21sJuzO3SGIo3WaB5nxJGOzXG
+vgnllc1yK1CwLXNtpd1fAICf2FR2ylKOqqcDS0jRjuJKYMZukkmDoy2JTONz9vjl8xgUGdIx4NO
KPa8N06xglB1NSIAZ4AF3AwHeD7FTIBD4XGBMKkadU2AV/iyTFLosQJfRa86uWHcfMHi6CM1tMxD
w4/OABkanKSckAcxHkkijau6fdCZpwpcO6XKYg4XCOzD3dGFUn+rl+fFmBh4XVB+2gaoFk480/ln
xQy5uKdxGAS+9BODtPGZMxBvOIZiJZQO0Qs/+QoIlNomlnyVzeCjrJMvYTE/SQZLe5M9LcTlzFI1
yfMJZYry9N6X64Ini4TXV0T7t9mqLO352hZb5t3mTGwb+CEbhXS2u72CUnrzHSEtsTuSP5A7YaJQ
UiX8RrDTEFwhJ0lzJ15qL9j/gJDhUn4n2YYCUmCnKdImv/gmU9wxGnoJAQcbGtQcs+HPlv3pDIVU
v+S68ayjaH7Q0LBU/5YLgkTiREQL/JjMKceOdKsJt3xSf3Wp8/+2M4Z9yQccICv2tC+clBCSlLW8
apHg5zDHN4wHtcVeCo0Cp/KJuO5giShzuKnqr4NdVOX2d1XxkCRjqit47FnYPjVuTNhxHa/5uiDY
l+A9O8ocNXvwlG2bwvD78dC6BqIqH5a0kX+SNEDyGrIkqNVTzx5PesIRueMqN10w1rBesxwqc0u2
z7LHZLiZdhM7YCydBuNhPrLj3DXiWoyZCyrBkZ17O32gRISPBdCw594YffiaZeyaRdscT8ZVJFiH
04cB5XTva7hSLYWSMIPmgZ4cy0DUImPa5fDQSIsjiLB4fewHPiiw5asySFSrv2NuZYar/Z3CYmuK
SlsKyGnep1bOPF+1+PBD8fp732StrPQQIlHm8rp0j0nropADS5c1LdAY4fRdfAwrc/fh7HjGakdd
gHCSi1Z3OUwz38p3mLHoTIShiZLzrFVMDhEQDCwZBuOOQNYlLBbxtKF1BgMhE4S4MA5/uXKUVPck
V532QJOIgkR4V8R2qHDn+X0lQfMHjt1xBStdIPAy14T3N4V/KYtgysfjuPKRlJbuhFOkZkgiMuQ+
ktrhPDeBIRT3Fo3OqNqc5eoyM7Ol7MdiV32SLt1PC2hFTAEbbU2eFpVQcl3EfrMu9rXw1SjUTdm3
+J4EFVBQU+O1+kByNGtbAuOakU+6UfQOSfDiIPrpurGuoqNlRxeCbhDcIZS3/eKtdGCJzHAZICtp
twfNgerW9cg3LIlMy0f0VHtr9rd0tQ6ujrkAXgKBEEXLplM4hM2AAv7pneMZAYlTGt0ffDFB9Bc9
4RZEtNw3QSEdDEpWiMOBp/JRpLySw+M701ULGLIEMYIl3u+r3+GCCfrIK+zifUcJVr6TQAel2UJB
l7VOiWwcTsmG6PXRi9R0nDufBgqoDq2C69Zwr+cszmsNPtKWfnXo3/Oc7LHZZmNjWDrtO8l8f2PO
wkf8m14A4duxDXFqsf4RwABjHOZPqUIyj3tutM356reTGZRVSzHrLqaWW7hLz77wnxny6Jp5fz4y
XOc/Ew6WnYHcFvWGpyd0rQKClVTSuc7ykt1wc8ah2S0e7SPBvfgHINEPCfa8FR5XvdrMkJA0Eebw
qpgnd1EiuO4gDhDq+TuEKdrv4f7fG2Taga4eTnx9A+AalT0haWFRFq42RURSpMmYZjnVAhotx6nl
NsqWR2QkFgBnGrRkxdatdCwdfQSGwCmwOMq6cQh+F8R247RmdcoLKMWxAJoanldPkS0A/+BUQSF2
4eXnE3jG/dHnPAtrU5+42fs8ek6TqMxmjQG1J4CJrdurCVvsDWNRuHOrVKbmabGzKGI5H2HJ0dSY
hFr2W+DbMOfYagyIcKpCuOFGpWAdWGypwhQmyrhG0yCb8OTySZQr3wXAi6d90l7ncoUHwrUPmzhM
ilhAZT1DwUEfwUihbOvnJkgkNlfawS1rVaij2eC/oJosES8CJy5+JoBcIG0W0ZLWIAw6h3+Z/4GA
SEOY6zdUFWSu8QSurMnhs2cG6adr7CQkj7hZzLaM15VOmyr7MPqKsjeamTTZR2sMUMHRWgvABiq6
YpkMwoBUu7rgiPcmboevfa8I1n6V1Yk/3+ZKHDZzHm3cciNFKYrxSIeNs9vQ9gPAtA0bomp0K9rH
yu3dNgYv6gIgyCdJOilJ/pzdpbZ4zeOZEiQp7K9i1GOxaLfjQgHgF0V8rQMWO2JzM/dUt+mFxznX
42MgNfZDWZT/DH+O/1lkyEBHYm4lDwM+Whe2rJmYSzXAhiHHqGmS01uB1jlzm33ZC6s3q62SIhru
ZFDMfrM4Q9rQD37tSsgMdf5CDhdFJfcpkwzJQGprAGALYxjBoZSs2m+2V75oSp2kKEKDBTXj8fjt
wJpZaCZx3I7bxyKHKB8skcLVpjv8o4pAxcx3helh7iA2CDY5L9dzyKLtrqwzEFqPuB0avNtOYWn1
HgnWTmqLmQrFco1egtgayXL8564l/6aguf+C9x23s4s5ebAaFA4dTfHSczWMsvbjAZSuByvnPleA
S1UMJWjl5aZ+e+yvjs584PnIoBPmxQMMER613ze7RRAe8B7R//Zqpt6ugoAldKCI3wOtPEzpkUyY
8i3aGuHPRDSKc/3tg2id7eQJjB/PFLD5SGcP0Uq+7J8SMKa/Q9k98hFD2Dk9J33v2vLy4mLonZ/l
6LQ4A4PezXP8JmjgEzJoPYvIcY+WdPlYYHWRC02ljl3TGsnImEWgXgLLKtERR5axUB99/SIQV4ni
Yh7I0I6/oRfz4Q4mLbyEtkf1/Bx+BsJF16FTsyy/1f5V9ff3yJ99ZnQzXoOanlqYp5FLiZ5ge6aC
+6tYW6xZS9ivStUfML+vEgLRgtRtpjv88uSOEjSbYh3GTclB0GkhG9RB+iKfTJGgghYqw+I8L1Wc
j4PiaBNbm0DtmT9ED4astHvffyavxeX83EZLduO6W/D0LDrWBMCbkHr7o+fl0eanbmEoI7uCrXXT
dei0Ahi41eJ1ooWvouRFtd9I/XycoT2IjvhGYr0lHZbAREQUeuKybNAF///8m3LmIOwPK6wvLCom
20yrhgYj2oEpGHQGMF7bgyh+LqZmiQXOZDXpfb/gQqijlGXWX0i9yduGetftG+0qNAQ5kOBXdijD
Q8GacXNFpGyIevBfUDw+9H8Yf111VkAW1FzwsO6RRvH4tWjIB1ZqPZ4PJDWPN6WkTNAfc3dtGWpG
UcX7oSZUaqebAiCXf3qg7ouu4KQ0/XqcvlB1JCWpE4MeruTTedCts3HXeIbmluXXEhWuAaf2FZvZ
pvtbz00+GsATfT7WQX1GtV+Z6s+280HvAGhbapR4OpuL6PNDfS2OFAbNZ6q0ScVx7SJMbmeHdShp
vPNdLZOYxIkCLDbkNoRk9dOaZ3eiCq2uCDJ8af0U0ffkFAW61JgA8i55dorcyICmuL7qE6iJzWF2
qI3XQ7K7rzam9T0unhHGSYBxcZRVVwP7olULVm9vyj27Zgvgzh6RRtGeTzmdtFaIgUsm2iLcjgo6
BgpRDJLs9n/tT+v0neyK98nbR9Vz6J8Osha+ohaS7bE967d0PtyvKXK2Zc91Q/4FwaKplAEqf++S
dA8XoAUx/g/btodnKawbBZFUP/6GVpLs53ovsoCSwfMjNP+lpud7fopZbb4N8sr7G0bi24MO6OTX
FyvKip1zMetM3cYrIuee6/n5d6etgDlS6k+pJp8bf/x0AJcZxUwxAzetyjIegMqBB5DWocnt2yTz
Dsgz/1ya8iC3DwEMliPhaIpeI9LJl/orqwKIGufF/dD/FOk9gGAZ98eXwnMqPKzwxRX7tGpeXmAe
5O4Ej2XI5yBm5X+l6SIToqvDTpRHtJ6ccg6tPxjsmt5MMX70F5GIdzNWdw7+jE3d7AFGAl+JsUth
1XTHWiMmaTvJiGfhTItkvu5bvm0KbcZKxH99jQ7wm1VpPatYd7V/B+G0HzePx3CHJe9qlZkhzsiD
GQJOJR/9s0WdZHPiw1Y7xNmOWT9RjsJCBSrwO/zwIDB5F9nLIMR/Nga47Ej42g2bfx+g4q/B6ETt
S9NJa3FFVKUKv2BaieP1CL4PphRvo4GhrLoGTi0PTZk1NUhYMFkKI/t80un7Tf8DkdI0l3iPFODz
hX6jtpe4YxKGkZdzlb4yP4DxHmGx6KP4cPgoQOF8BOdWkrZQb2eu00GArEdstFXYDvCfPGBi3r+F
u4jAONemPsIXYfFzj7TgLnEQjuL4c7nb/AyhqZn8Bl1waMrzRe5beHhW8Zxg7T5GDn4DWRaCvm13
99zVwuPOOwm3blTHEAIUEmdfHwp26ZoRC+z11ZvbzoBcSp5epRfBpJqCWkSUKu92Y27ZsdjZkibz
596qJotRA5TiNcFpu7nNx/s6L5+K92XyXq8WqkrbC5L2zQHPYEHiMLQ9laIvstuGiz1rvYtV5rl9
mg8uW11XmzA77iM1iBwk5jMl8Bh/VSrWz5/wbwea9Y0rPzE4Y2l0flEUQ3zajBnDQVqizCIx/p4O
NcW5/GDSiZGa7xdQp0TnfT30Z66b6nm8tRTLxWuSHGzR947qxiYSdK1uHaSaQBo1uzGZaN9l0mE3
1SKpPuxp72/8vo8trIq1QGUbmR4Ga71I2IEuGKNPxRKUKXtsz8p1v4jrRPDkGB5vBlgZ57P8zZOS
bn5N2a214XC4e1sR79fovsxdlfuL4sWbgNo4GKW9CVlRdD+UEVqsbMW1GuJxznlDyi9hpyTI3wWp
yZb6O43YJ2lQn0LgL4EBn3U3Zcwc61s4eC763QYITvmP11z3zHJQ/pY3IypC8ppwKjvJgVCT4Ng6
pCJJs7O9Xqisos+AiinV90c6QMwJZZB6pur2Z4meimrm0hJ1s22X/CuBfoglvR+bT/S3q8LxVuw1
fUkroPfh0Rx7eVbHQ2BMLa30oP/O6KsOYWWCDIPLUJfIJwjuj4hvRvf+uSrI+JNdRA2HtEnHEBwl
75N9qVQPRWr4RPrVVRRUc1wrVAZDWbBzgxR7cEWo49AFzTnAIlH/mCXox6vTF/owVq/2KC/IxiKG
+eA74Oi4H4U3D8yRM0XJLbNSKoRnJgsuCDDoh30PzsV89dQp5xv/mTjbO8dzKuM8l+u/ibV7YCOP
ZfDFIO/nQZmmDiel+UD6gAZF4izLcSczeleLzlUixMC3wzzBo7io2ikn2nFRZeOQc/bJ8UkdM1ty
4NMWhSws9O6aDunpp0MSF1aL+OuKn/sTzKbjbFuaAZnbPjarke0aoYBmfOqOGPbIk+n4VgPnD9aC
Gn/qt1RsEopp9ZczPyHYJeyEiC0NVH2aR8gNoCisEhX1u9Xjr+JB3gF5nFGN31CzxLZx73P+SARk
ofLL9lublHp6f5OCZMEJDKMtNEiNNDEhtPHO2mfWR/V+FQZR6YjQKcVJ/Qa9uKF/o6j/ABgBSVKZ
dC6E/S1N+eDXLwWFijfObKiSuWI7kF/FRdju+wU4hw/nz2RetkV514iCHh27q3cb3bMjluo1G5rj
s28LIkOJhpOo7sLtZGAxmWgz6+g/JhTv6YR+O4AINerjIJ1nFxpe4m5GuRgrgbg6DqEIQ1lytM4L
pHS79zo8f3iFnumZPuV71sS9Sl75kQ6Rzh8c5xNNXVStVJH3Md4BDuJtOJ8Np4eExBjbxsI2iwoM
BQS26VYUnvou+bhTZhezQlMJxKFgK6d+Qfg5keCg3MC1C+C4FkLwrm2Cicf+51oqhJ5bZJl1TVEW
I5LPepie6Q8HdyXVdxW7g4rA0OkTxlk11hZTbK7HCmfXzBuvpr+iuI0q+gQWXnsq+teTXrm1Or8U
vXYj9GzhKJSiJ5UhwI8ekgh0jSZLrSBXxz4a5+nZR/QYxUQph712dkqp/U3CVCZn8crpmvc2i+kT
vQGTAQ91pmVT2RKZ4xOcacquzamX59Z+0SUiHHfs67ffJOw2pCLVsrl9jWTQb6bm93EMrS9AA3wV
LhSXsF/x6KUDgZYDFxi7UwR6sUuI98dhIUvntlavtyC3Ipj8derB/hlxMEwTV/o4/Jpr9lJitJ+J
xTKUxAJPwJYYVyDuGWYkniEbB7VJLsDrhhKiB3jfSckDzUffuOdRShuLz/WQTzzc6TFKBZMZoh6m
qXq1zm+PzFyBh8VF0/pKPHeslCRZZg3Wwu8eZlO4y8ifF+AKZE44D9S8/lZRUMsdQLJsYS643OVy
l05Nybhxx+QO7iVr8DgmvrRb9nIEZ5cGyyBGZiIYxSH/KsUjG3BfJ2z+VDQmT9i+oj5Cyi57dTVV
Btw4Np8YITF1SFdEXrNRlkZLDI4amvST66RfFXFrQRottqr/18Ofc/UzkRlMkkp4REfDyssiBT6Y
SRXxCjU8bkWKrKP5QPIuM9Nt0FbdQE1wV7LUYyiY/DnDIQojQf8GHd9f4gkUkoPssI1D1ryC8dnj
JbOTQUVkBsvHHdR0KOMCIFaj0N64X+55RSW5PUmD24GJD1doCySBp/HFUgXtQ+TSx1TjpUpSjSUX
vpXxl66i6BviYGvD9QAk8XiiJtrEO+sxP11p/PtAVhEvGL6PXBVf1m1dnJvhvpz6BihX6u4iz7cC
R+NOoaV6StECNoLuETiAfWoqgy1VeKvzqg0id4A1gNC326bWue5Lz1eW98qa/jtQmvzjjbCcyeiL
ARuJQjgtTk5UAUXEWDNyzfI/2GngV+nCLX2QpeqAK8jHvOP0VTMuMqnuM5Lxe/Pfs4a729KGCASo
FnJNExsHMfO30N9B8YxD+og6hjmfQEEhlWBo5/3PZ//YZKDqV3S9pPnhWFTOPiIBHnsMgyoF5o2Y
LR0vtxjTSgDETF94Jh74kLGhfZl+08nyT1+pnHeRxLiJBhBviCpkntLs+Gti3jMODhgAQrHRVlTt
zVujBx8NvTVfHvLVo4By4U3jwAcKJN3PJJM1qDr3l8FhERNAieZ+rjF/m2x0zg+xDh3bhO9cAbFi
BLSxJgiQtRyaHt7wDcEzYnvh5CXYpVgtU7/Z/3O+gFHauU0qL0JWw6PZCdF53CEgnPl16oXYdqm9
XIbCAXBDxXGVu7wvh05l2kXZWHoc81C3o+t6qFGsD/Ix0eSH4qLbj7wTzTR2ikMvmngSUs3rZNyb
vhX67DvRVtUIvahxK3c6jRQcUlpac+STVXvcHtD3WN4a6G1GdUkTtBlA+GnsHVE6rtxKB9gidbly
5WsUSElxReqrTOq0LmWwreo3WoiDWUERUByguLANtZI+MG4YNODrmno8SFljNo6oM6q6W8CEK4AV
a9cgmsvkYwxPylzjgftmxDSvlhSxKYu9IFt6Jd/gX0jVm2Uaa5w15CMs4nbx3fv8MoxN7oqliYV+
jwKBwBMFFGaNYL/wDOxCicj8NXB8jkpZoPtiO5a6InOIXp8xlmRDUa3HWGmCwREQnUYqWbLiv+Qq
I0u5xKV7Om1CJ68WZozl2uCF2GemHuRir+JYpaHaz5iXJEBVK6dqrDJIkAfuCGGSBYcYnWnqOdYq
69/3JIJfZnhWIdAxTGmPUnBYKxOFF43JEBaf7y9MIjgQH35PRDVNVmLH0pa1ljD8oYRCLzLN4swJ
cZpIzEdoS8rH2U3NQwamS9b+ACxOUGLNjHH8C8wOU2ZWHOUtMGlhSzvaZriy59/aovPGW2xzL30r
3/tK74ZHuG36Q9TsnZMwFh++Ziv7fnOjNMEc4KFP0B+TijHFWXHvoyBB00ek+xCkWmSZU2Ae/q0d
AE2V9+ebHdzl4DLhShv61y65DXxIQnLfKtO7q1Z12TR79HsrpcZi5p79jev/c/BekPfWqO3tEJBm
gtW76DFwJIB4Sj+dRF00A3cgsWVfxnirNbm+BgX2YbkLRCCWvwzooP/TUNYUQVF6regXsNiC4as9
K7gDkq2WQNcknY0HMA1t1k/qEa49BDJzMMXFi62kSyNvdwofOO8HW/Pci9jNJz3cxJzBXjgeqdpJ
NeAo4aH+ottzSfTCePl4NrtIlf1VfJdSG1MisvMougTyqc1mJHS7rBQJ/pZKD5TdVFwwRrgJhdC4
DG6A0uor4IFkxbcBz+QaRAtZRbWh8V5eS6z03nk9G03D694D556FZNZffnEY7NvhVyWfzrsJDJGb
bgPaqdcOSQlZweHYSBnQiIQm3VufLVBRDLGE6AByMxI6W++CugL4WBaRWb9kG0QyEqtLk5If2+aV
78rT2WSeL2kRfCxyYnHG/UN5N8B/X7eY17Et6t+BDZmbr80nm7fBavORvVRMAYeoYU+CQy4ls57g
GqYU5kVYZODRFq8/vfi/e5hFsQpyzRTNsURpoXJiRDn/FxtwPLS7gDDJRQT8NAwdk8Bzu0b1mvkt
oENInJes0D8y+9yuUIumczyWMSWdLuj6/4x9c2EPw8mSiQt5Y/iWEp8yQKeXPx7u+FYV1Old1zpz
zEPwvLnjpr4ZfrKcwLB+VRFCqbpqbf3+Y18REqv7Mf+aWBs9ucK7WnFGR0qqESqr+Pk/SPPqW5Ia
TQLZwgVnPyoJn97G3ULv65bE7POmyPhd4+Ud2rULB1oSag/3/Bsq7mCYmg6lHUbDEvk1lko/YZZn
z/Mfjnd8GchecNEDY7J2ciFPuC1zRBIWY1/Q/ZgFzMK8PqHdiSRW+YMA6cot2Vc9eo4PM1+fZZNk
3DjLLUwQXIY1iXCCm7JxIiI48PAJdk6JZqhwVsfdFaX+FEfGnm2lS9FA3qMt6qsSFecbKMV36HgY
vhlVgCDYTpmd3RnqaHbunLiV8JabRWgryLiOAYf9+uiid5DFvuUA2Kd6PPmyHhB5iBvm7pXRqxUH
bb55MF/uDAzLZeSSeKqUy8e5mjmvCdNR2zlxhUEXat0cZVXbJngDOLFeJdt893Tr8icEy/6X/ROo
moTR0CmHa/2h2K5gfj3kAPHBYPtlkETbEXdE3T9nsTXm6ZK6t7ASE/a+ue8Lt63W2j9cNh5PEIrG
POVLZilghyXNTBkThKDcEJbsUp8q/5ag3+a87U2oDSHvmXxgMYbWYG4j3uM4lGSIxAP/bAEPDpjk
oOBCyffN/D5kh6MciXS+m7vbrFUeUp0lWGPNLazpqJMRmhw5Q0wa/6GCgUpAnW26KfYJjSnUxulN
KnbqJHNNMD8trGzwHUSABI90mt6hUpn5hC2gSqphtKyT8svI2WwBz2KIHrzzCrIAu/T4w6v9EALn
YnpEzcvTbLWZtYs6UubHab/Zy8GLpZIlEaazn21slKF/YBU8aig/lz+tD4SETTCCUfSwPKzOR4Lx
AWd36vt1RvoeernpCueh0Wn6FFbPVyqptifFYr96unEh9H3elritXEHp/YNkCGetC/M6K8/YAWkd
nidjgAmfFYhDeM7QjesiL+IPkB+LAcQ/EOVGmVgyrIqffBxMmoHxcTgDRw+nDfTDOMWFA7o+MSqD
RmxES8hSMLh0slnpRMGCRMYGf9QynyGSYwZYzPaERduaG15azz3VTqsW65inLW9MBu2zIW2+wKmS
plUEHUTicz3Sk8EaECra64CP3pJuxCPyrYqq2acYIAOKCk30ZiyZnB1kjH1IXEt8kTZK9BLFufIs
ggJMHHj4slZ+HjfXrVNvMyxioBF+cs8DhGILMG4OAKOIm+aWyx1KzNG0UJnh4bWpYH2TMjeQBAN8
PgyllU2b53Tc42fIdTz8BGx95pq4dNbKXAh8BX2+GrDvZ3atigVrAP9pC/G2vBZrVtrG17bibYGn
Yra18ofwObwpwQcCF/FtM7h0CKvYZJPwutrQhp1OtIvhVwUtQm1N7R07e0UWqpDBqW5JbTnQY83G
nlwmy7uXwcbGL8GWGMernSrySOmCgM9/M2EI+l2+8CvqOy4Ke4JveFeeRze1uZBveUGR7iYgzOzb
elDxzF7c6VYTHh8tCtkLt1qe2ggFIo8FgrgwpFjneAqCZPsjtCYwi4W1hRwoZCUBl+s13pEz+r8w
wFIdiiWeQoS4v/Wjobfuuvk5xEILunyIOvYmXkQlPQat4PswKlTP9+Gw2XyGUjoVzjtiG02XHChT
wrvqyTkHDEUxHpI3lCQO2SmwckSK1aieHehkFvMHXp7YCzzo0bk5zMV/M/nOBVmdzWDJRT/xlyBF
G6WBnEghHwfumZiR8HMEggOiCtRdgAw4LM9BUOgI/QWkr7UUUEQk0MBkxGz2ZN0ULZQdx2k0P9ok
iPoAsBGtoZrSHyjEf/ME8ch4IrQGkXQd4RPqJxEw21Xvjb2X9k/8Aeec98fmADULFfjtMrNN8q0c
OOoBv/O1m+zxysV5Qxh97ddH9dSPo1AdlUyCjW/ARAHEqXuysdYgf1yJjNv84Jy3c8XnvJqeGjyq
nfp41MhdjH9vpQQZKVxAxCbnDLX4XT7TF6MPsAKyO7WtexCRNzInhrT3No6h1ra3gG62/yoPIfF1
0zy0rR7WGXSTSXd7cTjgNcuto0S9/bKVULIPgt8kIQAVZ/gQQMr+wrJeGyBx4E3YjlndKwgyWyno
Bb3tOJhbNC5w5whX0SVuEGrolAzYnfgqgchWqO7WEO9llOHnI+c/mx2aBnnhwScIZLd4igRM+dUQ
zOBGYOYwlDYiU13ro5A+j3926QMJZM5WtyOrux+sdPJ8opmXBTXRbjIkaNO2F54OeuMtA2TJEmL1
lekDWFLlmzVkRazgC36grOXwc3jSfAccvc7IsYoUVMZDWe+FEaxdWYPVEpHNTpfvhbW9nBd6tfO/
d6dSVA4rGWGIu6Z46knjZix2Zln/qIeDMOv3yd9UnrX2w95SoP0LaAD4NT58MpjbQezwe1vd/kWp
Z1iBx7pc/kPRO2KFOC+6ImZ2QT5JvB9ViMobDqKkauHpvVL64UmPFUYWDA1IgnP4YlqORwVoSN4i
wn4X4PmSON2bTdYiqcEcbu0m2I6tBxqsItV8xLJ4UAxs6tmbbJ4b52k3MOuxEZFcr4K36L5r70Uc
BBF8CoA9AwT3qHkfKagV9MDeY8ulsmiwjj7M9mNy8OL3zU91gGhrjFTZwGlxrQbtPmAgUsQC6S5m
gU4qcdxtF1DMfbR6g3dSRRWqH/5ylDpWUAaqffHQzCKvNg88yVJBTwJZAbpa+w6QLYRS0xagBExq
mjziGTOauzM13hu/DZh7gXw0VtaJVOBwcVZ+N00Zp+J24OOolb6yAPNez+4FR1YQ4tWpDhSKo/yL
NHNUPa5ijvO8Z/lSYopnw6WBuyJJ6/yH2jjKzRhunZXS0ynqkt5qri6xaH2wyXs3l18fTZwXPSP8
cxDV8sOEUqDjbBouUO+KV+bPWhNwcIk2XTSES8+F8SuFFD7uw03teZMuxRfDVDSKG6jxXdhaVQ0w
wfLJOiDfXeqcrOUy/IRa4tWYeYWCgxjcaI0ilod9TMxo0QwhYEGuI2lA+ixZeNT+h0TOVYi6yEc8
I1rD/nc+hbMcvkM3LQ2k7vJuR5mmjf5CYRD9tFjoUeoAqpH/xffiWAhIzcu/YL+YOm8tkmgosL+I
U7q/L0zsk/Hox7E8TScisQYZbZ1cRTxzCXQzzMi9oUcR7xLOPTHScrnWMkL3xuhpVKNFArcDbet8
2J1jaRjssQCqMKfMa+40fKwG/d84y+ayKfkE/KcihXv0a/mDrKJP/yK/ytViLixtcdIVStTjhQGb
Hxlg4HMCzuqP/ZLDE3I5GFC/VsnEnoXD6MnQoUTcPyrOsBqzBnPAX9necUZh3LF9CufOZeC9HKxt
5XtNoDt1RlLi/qgUclpd6w3oorBXeokil7sDiv1SHaFJjrVfLDEZNYeGUkSqslddZQEKWuqboV/4
QWzkAOFR2pTWgq2WOFRx2fosZwmh+2xfhvez1k3o2bXAr7U/fhJ1xtdjRSOJYiZ5Ux5a04jU+B9l
3Z7tJfTmg2O9xqxafVAnj3wnvnf6X/B135jGF+Uo61yNpH5CUatKw/P3nsEM2YzVQa4DuiFBe2Ca
Qe21bTabjKjf1RZFUfgXmalju/eQnaXMGGiavoW3AcXE4knyHZhzSK1/1vzY5FdhocYMlVAmKnqm
YFBUIHwHhYFYsCVY7DaI2+vO4hKc4yCx3Kp43d3m/2VEz0g7SlbAsREY+pmb8jotW1b+DmfabyAY
xeiFavSrYghBUhGZXPV9w4fQLYmDpndxpxoxvRS5l5Wrcxr1j1gtnMaJ8grWZ+ggC66jn3Js+bSg
NYBKKa9wSbQ2r3LR7CZpm9++w5pzbinaXeDuBm5V8xi4DjnRlsY3Q2f+C5qBzQLg5Hai439rDzFA
zD39E6Ir3+Ec8T1dr6T7ycjcD1q4RyASqHOUfUKGAm+jnZi5l/5jRvbDniIwj+pK3f0N/M8LxJd7
SC8LC4Ypcmu/lnRZ1Kf57EJh5gEygWLaKS+qjXa6udiT//Ef9JFW5Xgt4HPZyKU5UNBH79pMrBXn
vOzCUxMBgDLU7EXHUWCmxX5ZHQ4QNFUSjat+Rx5tA1wxVyMVGIOR72rXZswut1wzXe88wOvm8pFi
Tn+FQUjSs7FlRVwzjc++juSXD/hJ6Jvt7rTWk6Q3poa49Qc3YCWSKCJ7TMiaqmQnLypexiBOdV7Y
h0ekdh3jcXOExTaxr60jvrfgEuEbBGJEkX4uD5/Dr0Cvxb6P+lWLZhqkOwrPyIdkJOq/VyhAJnBP
C+Yh1JT5ndoDmULz2QUNbM5OKiln3HBE+yTRQ84GsrBbun6WMFcHVQH/VPNleBZeFtWS/h9eutjz
+5tofLaa5Wj7KT2JaBIQM6WABplo7GV83Ks1NAKawnLaxhw096ELFtd+KAy2jfJrBNweMaUSFU70
saJ3ahb4uOQarLt8YYu8qb3nIbJGsXwuyu+0/4FZXTQfV9lFUTsB4C2ks4iC/vP9YJjdj7OFVkIO
QKjebHgp7jOHHL1GvMZV/Y62mXiosKhNSmZToCm7VNYiWmfmulKXNjTpuBdPcPTGcmIzWJ6HY20p
zmwVpMkA2jUc8z99Pc4wXdF9QvOpoW9H9dXf1o1ofIfEaK7hfbwbT02ZBkLtDnK6o+W07KRUPP+1
fSb/t6wMdkeRXonwkRzOfnetC0VZyxMWA+GyTJPVbu2oCUYf7an43ACeyzusal1hTGuVhBmW+02K
wDb315mc0fEP5DycsH7YY5wh7LoDP2U8FkAu066nS9+9gsXHXC8msfN+cmB0gmsFkuNxtvIAAaPv
sthWBlx9EkLnsJdpTINwUvkYFN1cpisOZksDmKAfcBI3M734zVr3Be+/g6/QO5kUNS4GpQsSU7mw
oFZ56nrfkxNvRFhVaIS5IxOmFlkzKmrTb7gI8b3JD6sHnfgCgIT6/V5ZGN7ZQkniWDUbdj6hQrDg
AXxlc3dCmX3TzapwGqt4YVwk4on47HfGmq13cOL6va6yFPBvFYf7Qmj2rRdx5ricz9OvZf7GJ6N2
G1U1adW2q0kPC2hrWHZdFqcS3kB+y5j+iyIMeh9OQ4ip7fAMvxs845R9SoVdOei93E0HTmGEjg78
6MUGlFIeZ+t9lDwYYNfMSTP0A8n9/O82FmBqwRDZ6uvd9rcujXlngCrshNsQ3XrB+XQQFp02FVHB
WoYs8L5ERdkT6w0Ehh5/V833eWumNuHWmeSQ5sXhxiXnv5PCfXPPM+hFDcCLEDEbjfPABnNNOl9X
hVkDSexwtjJDzvaQhCkOwKNbtTSZ2B8aEYp4OKiulF+ONFRTdIFh+y2vRGAZDPm4A2jico1rxD+R
1MNeAJ8PFHINg6L9YwudvKsNGPdlA3BGvMvl7kt636OfRNaA2F3QknK151/8zqQhJWi7FD8Jff7P
iJmQw4GdX84WRRRX9hOjmHYnCjZtw/eBwh+egvMjU1QqztDf6IsdirDKG8F6bl5g3y3s1aNnVoot
mY4qJ6UXagWK78HY4LTjQpDM8aJ5AMy59KulkGYorwLr9PZ/nDz0vnBzrm6xdsArp1uoH2cZLCOp
rusQeP61plEMjxXCmt6OTKbRx0gLTDTWmLmWeH/CMbomu9OEEZp9Kb22iJTYzpy7riNm4Hlm+X7M
oqlszo5i7duIUasqPfq0s0xYkA0Rv7Jn2D5MD6XFXCbdi2+NuunRUep/iZmb97wuft3zhDrTyo6X
pyk74sWDbiWxy+/DEYphA+WfoSq2suv1czdS6xaGgTBiHw2898FK91xqd7zLCXBDkFDJPWcoJryK
JoZNaLxRKQFFtEcw536Yb702RpGl/7342EUlj/Oi73xrLzG1EtGQ1o9eOkhK2z0IyYBdT/o6Go+6
yWp3cYxbV0NQTFKEhvA8nqlAy4dvWq8Wpxd0CUhluBmrse0hV+Q2WdKFw4BiHgjlHG/8EHG0+EGI
LYRxnD8CybMkr+QTsdF8fqJmoQu/M6+8j5esFB5FsqS4hFOvBZP1fhcwenyqDLPRl22L5bAn6BvB
8mQ1xn6D2CGZhIxxUDf3gD4Q6E/OU42EGnHBMcIRCuZb2VUSU3b6WznG2pCWpyo+7NaUcRWRuKDz
YOnVULlqooRsdtHHXB4PR2ykVu8SWukz6ZBLUbafCpBwtfgpaL/Xr0PgwsFsLH7ChBrbl9k4nsZq
npV5NYPR9+iZSkI/ZaLoHNt0s+0ivOUiPOjsmtfdxxn653T8fz/y3CFUd9gnhSuqoJxyc4FhXUAH
1AGCAACqg4zKM1KX8A4e7/LAXGFaxngB8+A8e8zWVeXvSac0rHO5aGeRs2TW7EaZFLZgi9MdAvK3
svUET5ed/5BODFrkGIz1DJl0XbFkrOGafnmTFlB7tiDonu7fWMiodY+5o8PJBcCTivpt0+a6ZfH8
1q0av5qie0A+h9YWWjtxJ7l4rGdGp5/MvOIWOU7eA8wIs/fHUjUKxnso1ZQWNeZtM6A5Xis4MrNp
XXBYN9B3VDEyEmyN6toH9HYYg8UhknB6c2lRZhSu7yP0HG+38ubchVed3/UPF08ycrmLJEJCu6zs
y7PhnbiIhqYYI1mzb1SLwrdoxxDaxICwlzjlWjtlKNNRwspOr1cQBpY/ehJwmsCZg9E/LYT6HM7y
TSpLye/QB5mp/fKf5PkD8kVgsaziJA902vFuoQxCqRPWeEt31RUFhE8v2EnJIUoXfJ6VHeoprgIA
VrHLDldx2t7clbyl/suxbZBCYddtRPKhUMhgFqVAT8G9vNqsSzpC+0iy7lzr7UyywM7vLG2GTPUa
uHFge9cEISQtViMn7QjbHuHtl4QpK1y+h3s87AayG/pFcGYWDQaYSufs2ufXrlDrj0LdwWTTwYeN
3G6MQ2/zkt2WrRuo7QBmW86e0PsRzXXuXfCYUPyfraVcsFpJga8zrEMVsPnTksvDJndV2Dc2UxcD
QyLu/VQ8ThXNgouiWuM1BQejnrMVvOHYhKJRslSrE1qb8ABb+LG8/7rShHj34XaOIxkWXe5PfnjU
9AFncmvgDaUgP8C/qf1u+a21KkaUd+q9dz2N1/Sb+R4Eyr+56ITU4RSzHUF9nUFCBMCjvFUQU4re
60dFofGwxYdaqAdEJGln1wOpnEG5rdcqvx4UZCu1P70tGrrlnTaz8GZr09+SrtKCTlRLo/jNyEAg
drk8w9Imz1+vGGlcZCK+iwueXzPbyZdXe1+9i68pkODyEnUzUt8vUOr9DgtNVHTyYjvQkBC1551X
MjVf43Ctoio43JBsY04Pl3nNp2O7RYC+EaSj+84pLwNdIJeNU3HdJ4T9ZXkDsYeuV3DkF5IOJshJ
8gwqLzQ+71Pc7kD/ThXphY2eZsBIeokNAZPAJ9R0DXVWPC+BEJF5ZaBm0JI6Ms2MlYs5A81m8TcV
dzgNGas/p7/DM322kpwXmvWcYrW89b5p7sjU9WUD4Rvzf04iUg5fDa8l2qGI7egLZGr9h7fLE/V2
pwu/e9a1wEAT/syGEV7RRFg73s2jXxFMnbm371yMt0Dcb8lYFFiueqx7fe52IXbkbyP4bKcOjiPh
s7SkeZiiJuk/8/Lyrc5EiBAVriIObSImevFfcuL2tXvfnDYiUBsR6cVUnfi2ASwmXycMs9yLNBb7
mQeRC49hKtbmjxWp/wupKFcgjWPsYQfr6fd/bm4Tp25fdh/VHyT1AuQPl1ng+pYmHN3ZACtnnxwq
qPTGT6iH9pBLDWoH96fmsFg59wWznnc82ylPeW7vXg3CBwyYy3u9M0bdB1edb2MQTJ6AjPLtHwux
iLQovpDaoecgg9P4nyvrGwJ8C2TMfeseuzLf6vExB5TGnVPP7dYypD16f/+irsrcGPeXp6KyniXq
eKJgVDQxJ3xtdIwL4vWASJOkjow0tKni58rs6PwMDd1rY12SSjA91UbmuN9ZpkX0Dg7L6Z15jy93
8zA6EpEHnUsIGY+MMMGXoLE674AYX4D8VUg1VSK7QuUZCpPy+bTa7epZBdqYtFD7ZHdtSLCFYgBs
Chjk6dq4plNzS1sy73cGzShUqRBajwFRsH17PHiufEsvv3c/mHYbCjUYa+PaE91u//vpbDZizedp
nj2/usD8Qeu/Sqc4EtpPiOubOQhdLsDxtQu7Zjy/QdRf1kBLn7gfux0el4OYO0CD/jq5nw2uqMbW
2uHvx+YTDMSa0R0yEoP6IP0e6Og8VQ2yGTa0wWP9xp5qsx5fkSN+izek3X+WW1qWC/p0rbAnwKzM
IH80HBPoynzKBoGbU8sVu12YVEqu4aLFcxbMz5jUlzZimRdBcsWUsh7z1jS69ZYiov1PbUZGQNob
SMpM5DFiqncr2epZCedNJ/nA6Bop7/0W8EzgivxNDRBa2yGKHJpmO6IuX+oc3c+r0rdhEN57vGGc
K5a0S7+iolt2WBQiApZncrxyhjK4DpLiUALbFU5Y5WTh9A10MddN8LcE4Bul3Df0YF/nhU0TJ65I
cgZc/R4u+qou9kPCQg+pON+av/hqPPfJQLrTo8Fd9AbV1kpFDXMZOdJHoYEpmWwCzekh1G1X3HWO
d37d7tHxuy/I+b39YntpvfgEjZ9oNKhosREum8qQ+zpCcjDa+1kGZEEwLxegvuW1To3RvckhTrkd
eW2eCi56c92Lg53H61MUjNDRRpohY+G6EMPn0sQVKxHVbBfMcccrAvQ+8IUZqei+HelQ4EDx39nr
4V6n+5NTHVcV28p+KkmeJRZrnvH0AWnEOdTwgnYR5H4yFu3xxVT9cN8loG7aJm5IYXUNb1X9sf9p
Wtxm8NsqvHDT7uywuNu+/2ocnKKwuAtrn9vhfA39pp/i68Abeq5KWh525Cn2hKQYZl/j23+VjNNl
fk81c2xDQm/mxjXysHaL0SYRzHV+yTvS4Xp6DGFto+xlvdfgzVQxcIivAKEkIclZ23qET9reKUaw
iJkj7T6jNxrMBGELj0L8gLbpwFG3Hh71jklAq+9H7NdwBa/R+LbIpwFO2MVVWKoL+PB5JZGIPuvB
Y9lVosmtgSNR40GYUa6bded3S+QIAlcH3RG0BGYxM0w1cw9RE0Ucvajw13kfX8cY369NWuQfDhVN
J+Wum6H8LO6G1D9Z8n+kpMAG03plCJadAq8IBEwvknr93I6mxLIixtUWAGa9uM/L26UsGfCD6okC
Xg2JLE/i7QRBoG4zNBeNSgvPbQZkgKNIHDaDp35VOOyzbhy37To5yDkTvyxEZsAvoZnWbUcN7IuQ
JhR62ZihAd3pnDirxrkRe2EpiXM0ciVB9V89sV4rb3o1GXwDLQ3oBwypjDTFRIbkz9IC+qovRxkr
BRaO/9gkKRReANBo1RVjh3zccyFQwxyidBwVlyRJOWJnfkh8lEhPGp2JTBghnzN2idNQYRp2nKae
44H3RZRNsgOQ9tzVq6VwOn5y4HK1dlRyH2a7quHqYZveLnRb7eeZ7C7HxqvKaYnL4czzYMU+vFjv
7GFf1SvH0iifuU+7NlNnTsvMhTLeAv7h+mEGnPma5H5J6RmjLmV1LRVhMYvXP1jwe3AW+fwlDTGN
dbRkJ4BA2unQzC+O/4JZrvXMupi6Klt2Hk/z6hukOLXNj0F6bEwPK2WXDAKntfTgS+Sd4P7CkJ92
PbQOwNlfOUB3Gv99kF7FiQxlz3TqFyGae2WhnJaVYsG8tDd3kC4CmVG/5YyUPdP+WIMSEkOvimPc
X2700yVdHStALcPT9PSqi7caMKQN0MIQuBzhpaepiUpQTpGm1q7W3aVkLrdmJpZAKAuB72Djs4+0
+TtUhtxIVubiO0hJNcY1AmmMgRN73GSYsbXEIiuL2TZgO71SUdwjV2GaB4jya8BJgs1/Sbw+hoQ0
4MYmquXBIh8AHgZczMJhFhkj7j7ZfWl2E8sBdKe13DTQYjhGmc4VB9ohNkeRaJoSaqeuclgixs2y
EenLswMqKQRM8CIj64rOHI0AMbHTdd+dipanyZe147EMzUSOEQLajMxMYYuJsaJKBkpCuFaf2nIl
Tspbn0D2NApwiXAPSnG+zqPtZZVyCyU5xcXzZ7o9StD0mpzF1hYoq2x4uw+hIqrTDd4ig7M1vCnA
phJAnnA+GvqtONqKh5iF2IUqt1mml6hxQ/YnlZp+SP3kBaN7uJKL9cVcK/jrTiGlxNi6kLOokGKE
eqoDcMKrRt/ySClW2WRkBC8bkmzzm7PrDHZI+zJsV6HxNotlD0QdRTtZLdcSFV9YPFWo2B6xwSQ/
sgV0HbFEgOXSR2doXrp/593ocbvSWuhvJUMP8MT12Z1NfJW0DATDyQ1Q6zKLFztGDWLSJpvalHOJ
93zrb4EknKJn1dPwf+DHKTL1PrIbT3E4RAOIMvJ5zk3+UZ0M0tILKpIFhCSayhDwPL/ByUWO16hv
GWjEJblpKoZwnKLvWFcXPjmc0ZP+NvLakilsfL73nzjS2Droq1T2cefymxDXcced5M7bltUwymxa
4Pn3RMmYau12/SqLJXFPZUMxmqysqu1q2tkgNCkMOW0UQKfQbHifHCRlha93NDdn3p2B9V8aYJL3
ktnFxlzXraoMQ1vBf39FU1nKhzxGK5LSzra6R9fa4ebOUAxm7Qnc6zK+LwgD3vUS2gimrQNblzVI
4ZD19HUI1pMi/NJiC+0agZK4a0rDSpzRGJzPctTEtTEzxGlej09B929JCLgxfLOHlofEfhGvcVuz
V3ocPHWJrgQpeoeN05rw7tSsWWTYMuPNpVK4hhKmPsxN4rM5SWkjpWHpM2V+8C52GnnxC0svJ6Y8
K5mZPDqs2dGdFygzWZuol+f0W68I/7JNtH8pOeFH7qlrB4OviGSnTqO/sekur+pJBXUgNEO005+o
2cNlHGa38DRFtUyIXe7cwpJsMnTT/rM+iIz/qi54LsG9cB2JEpg39yt0oBZRrG4nUJGZVESG1vjZ
RQwqEcQFvptoYh4g/yeq65hnjhSSwRFnklDOkOdDCPYniCaHBF4OZiVk1MYpb98tIDvS2TkE1JC/
7iOFqG3UYfwSE4lDphobBffXreLvvGwSp/2hewT2d7idp36ckkPZ9npBybSRInOEOWYGTvwnZ0OP
5yfnax+XVoECL7qw71HTK37YDsbGNxVRJtCKsIDcyww29B1vx9to1T6WG2wm0X9leMM5r43SM+fb
C8hv6mMDGOPeAcvAitoxr9UnL2Q+AR7SSG0J3RzVOTWVRuXZKtEFSeuo93RQ4K+M2uhOwKhzSKg2
WdYCjla539rnNtcGgPw++eGKHB83jFowkacTORW2tvPiJbgF7RSQrN2XXwAHZCGxl2o0rNJvuCRE
FLY+8Pao+VhmCASMCCnn9tYOhKiFoW5TMWoE0oJhsmQHanD5h2xwVBTkdUXjneM1bzkxSUnoMFnA
86yQBEKJK3E8NUbV3MVyNlnbZXI0kgNvafoFKCj5nxYEzg1XbiFqzkkU3qh1E3EoLNXNwASx4B/X
PynMtOSMWxq1cxZrKYrAZkCYQhItZPqJfxTRiiV793Urcn4Tao5vy8l9M1QTAHFJWGrNqe0YieEW
YoNzQJdBCA8b3pgN62qm3OTwdOL0BTWaGJ0nBksdUQgXQCtPfn0QZ3rGBdTERjakjPHQEXxbgdgV
v+9aOGrWP+wNz4tpBFd3xVSQ2f891VOjWcz9cYQf9oOyBU3RKsJlVHytc/4StDxHSc3pLzGEFNBV
ha9noAHoWsrXyEiMIfzfLq9WimS4mhHkhg2tEV8ZyHIHeyuEyg7tdEPnx1lwiFCo4oZSQiFpOgcH
TvRS/qIZLIFUGaCiS1oGXZw6lL7mWne8jrTSVuwdsO1XCkURoTtmaAMHDkT1/A1VS3SURelOT+W0
iJZ/HBn+NaJ/mhuxpTN+gGHIY+PrBml73F2fRKx0qli21QUwQO5ik1VEg2JaITkbe9SjIC8LPVWW
YrtgFimIPw3F8wvLxdVaqCBhb/SdGIGzNXuNoEx7rLQytmf682jqLuguIWHemppGCmj1FSoY8ORu
Z3Mfo0lhcMzf3y2ErpmNGADjMUM8Y9vPike3G67vgdjRlU9ND0igeJtNFUzfo9guCP3FGmXs6pYd
UsN1aZTQX4yJ8ySNEl4nVvz5dgkvTI9v4JrYqlQUJBTS3Y3POVcow9QCE9RKp/x53cVHAi/r3JRx
bcfa8loKZnQHXpgV7w3TPSHP0H8d9QAJBMBBfFcZ1nH/t7yZYBH9rpiH3NTO3jVw0LLpzTv3GXIn
dhGQLPJPwTskSEFj+WT1jY8WJ7LI5rYgsj6aY1PoFk6DUBQPj7liAYsR0oUeT6XGGuT5h77heei8
uhpWr1loqAAXlUq1LFV8EP3U2h6JVUwSXqkENrt448GSGAV/mj836J46QD+k7eE3s1C5K3l2djZw
RgMymI7AfOfAVQHF9r4melZwAyevTQs8x8jaYuPJphhTMhsDUBXtYmerdYMVqmbjjhJPo195T47z
HxvrvRAJtU6gnAFUNgGsHUC4NRF4jcETg+MWsUaZLLOhIpD5VXhj5Ny4Ry2dGo6lAEqc2kG7bVVf
eB2cN8hyB+6lBkb3F8s5CP0yiKyCbh8EOyH3o+wx5Aq0bJmIuNrEXlQ6N4b1qQ4yjxnYrx8QJhZw
HD6tak47hu2WidWd/KrYkIUbKBmvu5ba7wM9+Ry1Uz/GcTUqd3zKSPlQMe2oSW2WJ5KP2d69NzmY
aP4BIjZwrJ9yfnjGzqmnVHTgWSu727dlvGPt0IYCEcSXwe+L203Ze6LJawxTBvTaM1lVNjnhq5cu
/tTmhNxCpahp7injAaswa3TQ9OrSAEFR9pLkJ7cqWL+9nrqPkIqPON4wdakzsKgqiGgf/YVIhs3f
o9ijiwuFcvqmu+ixUcSTEd2rbceqWLXioCCdOD5YY7A+WSjzPWiHYbJ36yTq1yoUSOdziYd6bdtd
6znVVhg58M1ydsDS8O/4cnC2cVVVMeiMrDHXoF0CW1njuWYgG78G4vTRHpMWP+3+wz8wccXZGVh1
hFA5XZ+nQNMt8vSZH0cUdHalr/2Noik0ggwv6UwSoDSVM5UgQjnQF8QsXuODT7s+tUVkCEmqghZb
i7eYgpHGgeJod0a2T8cypDgwlFm3a1XUVmDxSdYXdzzQjV1zSJnOdZUvRrO+ReuwRxjwouinDEPq
Ng9gJlUsKQqlPjvZIl4ZhXKYCvVg7REiEoJAdZq/BEUMAGN8zv5C1xLJ7FAKXlWZvccQw6cjG0EX
KzjddSwO2316oVRPjIX8rEebtdCKMznHOfMz12D2wO7PhPwPva2yXHsaqqvSPA+1mLt7z1X3BNad
DM2QjZAVXb3ft7RIh0E9xZwancbadGLLIC3lxBWZNOWNeZEIqIA4G3LbgdKyMFpOf2j7bkn7M8oG
H7j9Z+9w5bIrzDa86sy+3W1x/N4s0C87AGIOXtwPPtfV+56DMrQclH40dsP+1qNmH9sE8RHO5nP9
10Ew/LfHBsPrSEnE1J9m4R6MKN8YJuL/rlJ3vqJ3Bq3XJHpY4AcNoJzYmJ9UXeNhH8PR/XrDZ+VM
Bx80gQhK/Q0g7w6zbRNuWT85Hj5nVADz0fHvT5fXZzcU8aazDILv6VSLrFz490BMKVIHEEjYuzCC
hlkT0dmEct/qqE8HABM5GeexgXvW4494nM+pLqcysOQFCmg62layw2Xl17bpk2WBabd7TLSbaqKK
IhFl3CazMEdPu1xHmVFbFEbAsuBr0jne+PIFRNQuPrDbMuhxZolB9EAQ+OTdyyBWMtoIQ+sCHW1D
eQO0OQwuUNc3GzLXOoRiwhjlXcwEgvLfNoFZ4MnjIZlHeX630iDSf4uWnMey/DbZKo4MMvpW8m79
1Q/9ugUDKDusA6EsGXVtH7glGNGBN91JiaBoy3Oiwca0s/FdbXGmLjqTVYUQux3189WJ+rPVemnu
flZC/lYLrMRf5UX7ZcEdIC6KmHEfMjOx5oUBxPfYIkTzfcWUnyXOg3ZYOggp1//W7zrMCJgnvGvr
YoXGoy43g3i4msGYfBkvbtkpjPpqEC+QYUGUweOXnVIPZI6rPkFVHXUKC3ulSbr0tKKnAx9XwePk
1W8i+jbIqfv2MMoSZntORoVqgnAZE3BJ9SCkXreMY3f0vI5bZB4pxXhksWOsEi9gAOHKzVFCnuqH
cr7thobwM71e0Nk1sd/tCNt5lDaeAKKMm84nsVDpYbZhWFQxxDOMPXrZjVmO1pTLS46JW0IF5xqa
ictBoO0Xj6Kum+20OgCWaMtd+sRkzZirQFnIhY4MPBlx3NGGZTuPZR+OTQr1UbycTANEWjFH0DVT
MkR/1yUK1GAqHgRMgtKGyB80PjkzMRxVUs089YGoPSlG8hEp7xpfBX1U5Cv2rLLc/fKCS2IbUJCf
nDt+x5l1p9A8/iusLyppuDRxPfCc9LVk+b2JHSu4vmlp1AZ1hC4rZWQq5++UDMSwV1UWpGJGybZ7
pzRqjYSog/LHrqTnFNF87dzr3radWinhmzzrBpbj1Lp0c5fqFjRrIxbDl5oB2uNMCv6rXa01uxcQ
hl0ncaq3PmtMAaPEG65mCGEjEDZWB+U5XXYsgfNNWlC/EDS2byhIfgjse4DqcVxb5RRckTP/XUu5
cuT2ZTg5UtXhK6GOoZdWQxcJAzMj/51pdGgcIsI3DJpJa1geF5JjX8S1nkvSJp40UFTYkBn7U437
IOamcAEvH9ypEOsA07JpuIh9Da1r21VS2UGH/PJikJnyy4ixL0+c7rxpfOM99JDreCQuLdDhdU/G
gRmrTLN/MUSA0SZ+utYgjKkg0wdHiRj0abiM8lEfe5VFC18IC14zjcXIoFGCEHUiFTJW7TuvQ4rx
kUnC6BCTkntpuHdJXRP7P65KzAu3OQ8WyKt4alEWmSDgJnhMnYqyShH2zq+H67e03iMXEmUAsLRm
d1YuhX0cjbAiCYR774ML50Z1MHorSgYTCC4nCecFRcnvL1VggIH7lPXOol/eNlhviihGa7jdBq7b
xOwgJyISX7dzpjhTU1oe0Zr1eapqE1Nx18+r2XzsOpMI3NYK85FqwABRbYCMP8FFoykZcqlDOl1B
1lOWqLpbOXM8X/3zxMaAD4DwBvmb8fQYiJC17K3rR5jPGz5wr7+nvJL7AZIP2vkMUmNyZ553misO
Y3kB6xbrC2PzKCoT+tCjPbDoxYwbus+krJ7P5VI/9asmF5wab4zJv3JvNGo3omq2zFoQ4WhjpweE
lSe3FaLFdQkuI3w7qtzpj0G2EcfHODPeEFPh1Txmqit6+3K/mIXO8vjqWmAImmv9hGb8AWZSlx/s
V09yVZysUM5hOqBq0hYjowzgizDD2E391plSta+ua5hfZ81wdJEcNGwopw/Z++AUKNSesXDwrize
f0ydACFbHVwoRfE9643sskCtX3bUp4vohEFJqrsHLkqV3M4Q7KZUxTDMsD1FFFNlcsYPXfGT0rIW
1y+HJAVwuTTIDMnrOo9jA+FmZzRHfTI/HoCVMeDXsyd4AjAwSdsA7ggRwjV+oWYzAd5wgLdEWKTI
gG41MNRsTF0XbmZJ9znkCmdwqty4nOw5UmqKow0ohQYq9Y8klH6DDEyAEUDmEcd7dOgmJ70BKfRg
jvUiWEZjM2KaN4FHSAZK1sv0+zRGbXkwmXKm9eIHYSYa0FPPMUJ8rcaJFFu525WmJ8Cd7IKapp6j
CzQWmrlVtEyur2Ucmkd8aJ8pHCDIgW2/cQK1fMejxucznjZmoQ+vb88F6K0F9UD2kC0jkKCe4idy
I37cL3lSLR2RBG3RQ27ZY2kjU4PYvHcX6hMdRlD1W1lsgNtko+DSA57HKCk23zATdwgfNj15vYM8
g6bqBtGAAyTSY17J2lkZRReOabT978C4HEygrAt3OBbMA5i1k00QCsTQwo/h6l6XVwlkeoW+3Ube
XJ5IUl/6sskdkijy+MBzpcLpY95TMTmJJisJiRjUTpt2Ob6cgrqmtR6qfxRf8x83I9hWX9/6hwY4
i+GTsblTbLFgK5aNM2QH4M0MiNSxTcOaPZ/Yyp2i7LeU+xUqTg28gJlN9JVlO1f+fNEvZIsopklW
e6etBB8Uc0JKGMQWTSUanjYiwX+Zu3KEgVrgqvIC0FW26jZuh2yqy01Fxk7obxUXsIsQoP7ITfQ2
g1JlZq5oLusdsr8iDXqLkdgRo4M7lkkyQv9aFClxokJ9dytmxSUauyEVARKIyzl+RA4CAx+v4at9
lqQucxLQX94sr8pFhgUhfvR0wtwkvB/VBDgi+8vXtQj7Bep+7rBU14A2xWhrqWBviEGGRMkZSKgK
DUefZXumAsEUlHC3qfSKcZbB95qZC6gb8YMaOFPzRtyTOnolN0FodxbG+AVnRlHsoowEc1k9lWmf
9NVPACNs5MuHz/7aZDwvO5Fch+kvk8rggHhxyfyx1KHg/QgYgZJSbY/Vm2Yb+QBr2IxKW4YzDmJd
sFMs0F5jKNjKXk+vqSWr5VUPcBvaY1G6GPplsR857XfzYQdlij26Yjys0Bq1taSTOl6b4GvdCeIt
rdosUkFCqVmcZhyc5IS6qwduyhIEkP3js7kbKpCmEhYvBWuzQg9JbqKor1VjwcLgMyd0h8wxoi1Z
NeGFBiup8Q+qZyFgENg4oBqrB3KWq1B8lO3z04EC7BWU2H8SHQMp7fPVjrrE00MfBH7FhVq32T2P
w8FdPWgXZupBAVXKQ8TPYAR2O4MYulePqTttku2WGPo/ugK62GHbS8gstmqLL+uJBfCpK6Isygn6
3seZcCjPKLnW/EUB6wbdX4lmptw7o/XvT+nP7w7lZylVUMqjYtGswApy9xHUnTGayRLZgVN9089U
IQ9bnfJ1+loAPDDqluHlqPZrOWTnwySkElQCkVE4BMhwdqfin7whieTQJ2pPV/OP3jRF2n/vmGJb
sHczTlfrRq+zKXy4gLpwdYjH9Gw+yK0rIIW13LM+Xq+ojNfdrNLIeER8MKlMWKVbVATs7h9LXJmO
gKIHJ6bD5kmngLqQXtrRtx15EarozNafZYbH+qpPRfdR9rPW2XQK25DcAtNWYOyrzTCeiNWq04jg
BEWqb3UR7SMySW/qP5rJmQabANFB8SewuCgN/mb0+oKBaQ6/dFnm9ZLNDp5aRcBoxIxIthaZeaHR
la2Ed/7yOSn8bj4rLrF/wk0zCgHIQkeeFp1nKcK5+Guh5MONFQVlGrkGNI41+9dWfwysiytf5U5k
hl+3KL8p4apODCAeNfUf6hzKiQ1ocRL7d4V38t6+PEFDRUbh1ytcjEuu8zVTFxQQY5Qmr68CBxcD
uFEQ0PuGweUP9NBrTP3vGKca14ExXsw3fU95Q4UKSpH9DJWcUa1XhAV7eT896yYCMTRI6RhgJQkF
Th5YOT3diYLUBE/Evj057XJ5Fgs5UILrKa6qzMCbW40x7A5TGXmsbZeY0KgJEepjG0tnLGwJ2UtV
uKhwyG1QW9tXQoATsu7fgRRKYswv6gOPFcFIGKo/3sHNj7fW6oBlDsHEw+Vf7gDUuM8j5jPbjYkc
VQZI7F2713LZvXfXDuG0m0vmfbJ29ZqBFX0qsa9YVCW5jxv+ZzxhWK4tjbFKULT0m8sy2doB2Jn6
kzJCv+CQZH6gXNcLJM2utAnf1+oX3Zfa0pZI+TIqKnhp7BpCFdrUdHssqqNKJzoi/QQBLtOGytX8
a8Mv0mUhvJZ5EXWd1V99+7IYGrK1n+hTYkUa6SJwkzcexUX6AtYolxfJ7OdpaCIIhJnLl1HFrQQ9
nYpHfM5+b/3h09PqBPlGIzTa/+0UEsWVHjjXkB/chKp0wCmj1PgdQysg7y7PKs84hqfGIsp3Ohxb
0rpBZTeeqEZEvuMZx0nALtHvufPQhvQbbtQWgCxGETMNexYZu/FQyaMwLAtvTj2oCyhhgFT/I2J0
X0+8/U1Vq8XQwEJIAxJ/gxZKmZiJ5aLH3Rpu2GCqKz+n1wHu5dwNPyZrggouwzoQKO7w9bUNGhJg
SNy9ndWs/wuC0Z97GGVXfXCazseLRF54y1HplbfcF3RWlctVTzixkiurlsS9XyfibOmnILxWcngt
RMyd1i1j2so5yKJaDcq9WPQGJaPImYTdSHHbg6NvhVjRUYzip6nhdfd/dAcjp3eq1DwM9pevcK+H
5tCdXMqXJ6bk6tcYNa40mFKgR2Sxj0StHHsm7x/pFfbXHccgPu8uWyfGzU5gw0uMSdZCbRmUVfAr
HKO1NNgEMRg8OFDwaWHnB+0Ffck7lkSBk5OIgFlcFJicpioGxVcibazDWalsWICMmMmQ9hbpWwWT
lgLW1HH8blrkl1nrGDF5EBQ3YgAwuhlIlK/4Zx2eZHkV+MuFskuW7hStZibmfPnlH9I0VFrDHnHp
ZT69eNRcfs0GfMghkLyeRoCPIN+vN/2NFVwkPbHxN+U0TkQn0mCiI20poepEBIhkI2Myg0HioZbF
07JM4dUdrnepfQhpM9iQSN4XV3xs+QL7wuBNTEDy5zE0YQkRO2goOG/ElbhHMICP+7iSPhYVCpaP
gRP3e0y0NbGrH4xNCjCBEqRIW5RHrn23mVlAiOkpbkzsf4EEIto69dd7SxtEnOwVb1/l+dvbOFlv
irwUKYazQc6n3LmB5GQUA49rxRvHwANFvTtgpnRr1Uu8cwox7eld8SwPd2UzizF/vX6/goiydeXH
J4vgcraggr7PDIRbgf+Np+jAeInogAhtVn7m0SiFF9/XK4M+0I4SOIm6f+8apDSp17CjdHwAZGWa
NroUX5+F4dBWI2wlqc17QVzFZIQ90dOrlP+UFE0lLYVZAUq6B46pFI4Ur4ItH76FeiIdmocFKDPE
5PFA5HJY/bkSB/j8kc6XM5ZkIc+aAcvVYz2RnAXMQ45d17MbYn/HUN624gV9GfIaPpXUi3uv0k6h
GMYuo456hLg206F+gAG7tUVlb6Nr66EJYoiSDmPBP30MdR5oklC9K3OS6Rog0LzhJ7u5jQOODyT1
oFUzqTCU8/4LzQvxIasre42bYaTnFan7ad6QiyPgBr9dBuBfcpJEhw2eYykFWqd+L8RVdrPVTvOC
KaX0K/BW91F8OFDqrzLin8fFyjhNBK26F7UFPh00YXbwSjdzVt7wrZQt7/lggc0DIYAPt5wnVDQ0
EGJmkHj7BxsZymUI+l0u1Qu1OLicwmjrHgPlc++zzwFuI6W6pJoCOJ58KwTRYS4Qn6od3VTWH74z
R68WIi5oximSRzOrp0HlCNGUBRonla0FfMKQRD+uILxzJ37RuxhxsA+0KdbOffGQiZzUm4htcV6x
tSWOrj0vFGq+n1RS52AFZ7hLpN7YXEyphQbaAFK1YNqVFHRlldPxaHAIOJSG/DSaNTW/q9QRxo6Q
xIb29l6TAH6M+LgB1KAYCNvT0DOf5LTgCXMcsmGm/uCUCN9SoHULzxBXEpCwBN3cs/kq7nm/nzX4
Fs2Umus75+pm40Z9o68Sa0ffKvPTtGHwjBiZRRJDifXT5VXIEn5/y71YozH3gBWO8CVf5SQWoDZS
uxzNCa7OAfqHbkcID9cXx5F9Zil1mLlOpYYEGCubcSdyJGIZb7RZGBGPNFwuJiXhJB1Q/JHcQsrE
F2l9/4X40HRcEjAiphWTD2dTxX63JE6qJiwSXUu455nLFR7oE0SuHNv3dM4vEmxZWKD7VSsmn3D0
5+/T/c2NX9QJb1cPmGeLFLUGob9BqVAhFdz1eEbJLoR6ZQm7iGuyIK//YTV9NJxbj3QXWy3VArwT
/hcYomBCv83DdgaKPOqkYfP9XmvozDpPl0ZECIWFAqTfQ+QXPbX6rPLlUotaossA12hhyYB+q+ax
sQteAUYcJYSzhcXUAie9w7nZzH7FqvHxvVkNRAsBvVQEJ/vgonMGeuIB+JuY2IgahKjRP+YRTOw1
mNQSCNol9RW7+jhboz9BjVJJNo++gcsIG8knWifEjdSCJCrK6zha3pcnPjMd4PVoWr0iESx+hU0R
0K/LNg3aXNt/HXvUmGTzb0Pu3yhpbBLmiCZzftngamWrOdV14eUVDyjMbWJRjdRhFs6RGRT7PBOB
oJQFweuL/NPz7FTroTi/aT2iRUH/TrxXG6GZ8/kT86YQRHBl9R0TCx0Sdy/2vRtwiDmpjIn2xR2N
dCqrl4FCbyOR38ke0fJ6+sDepQW1ev1b6dt9i4vGRxSfVbE4bIZNGAHS0eRTbE7BkijKeW2T1Tcu
/v+9D/3iqh1nGRU7yplOHP+crNcXU1YxYzneg8xukVYvusq220/4TCeAou9pPjrhWITwu3icW6sA
q60HBa35zsZYFIHNn0crsC/EcwhpHbxRed40a4VisY34AhnLqyYwtu3mD19ow9C1jZ0D8Cu1zCek
XU5ejfT4m9wIRBb6LljlJZguMoeI41vm51kQZleoGWAvXdWYx9WsN5K+aV2wPyrEISkZGT14LmSd
ClIu0EeqQwzx2CYlsPC7p/p6SJQnzyyUoYVnIxTaJm0z/0KdP4OcvZuCv9oOIlHsnDN1Ec5PRb9C
cIzF0Fejh0Jct3a1iV2vy7XXd/cOq2nySz8NThUiSu/mKWctdGpiqkiHOpxutkVgLJxT8JYI7EHC
282iseUwz4zpyFfgL6dbRwNkZ6xcNrkmHyRlwCYWDXhSuIWIpBJUp+tWPsM1MeFrCJEys15mlIKk
PgOPO6sLyawNttwfglS6pz+48xGcwPTcegyNutVuBjE9ZfX4G82MWzH4mqZWK9zwQ/zjMJ7+Rypa
lpIyXcUwgQdhknD1iASXubyJiIV0NsRC2oTWeVTQcsy6MujSU8XdgKZ+UsgamKDkDRAHfgBhst2W
Hi60hLAqJu5TByM0WD8IQChwF3C3xAufFo99huO3MOmqOlEwGEcyMJLxnu23rUtnnavDLjgHFzGc
L2LSFCrVKs6KufbgKJAgBsr5X6ZiYIwOh3DigmNAJEx/iGlyfvGFG5QunPFBCXd4NYnwHzh3wQWA
noThDS24wYEfQ6wqdfiNmJe95mAjsyWHo87NKBhBkWMoK8ysjQhU9tVjAJRP5Wo+xiHiRS8hyPN9
Ib9Qpcac8QCxFXzohceq3biwexyBwBZxjg/b54+jTmPFb7m0bjJvi4OXj+CefjTKfCjj/qXjn+ot
2wSX/8aey1kwC6yDF93xe82cp7P99Carn+nsXo194tS16MErgyoaLI+3Cb8/7S6m02WJvxx4r3gG
YnQBdLTmyQQhgKqF+MbAXapDSgScbMSEtxQfND+5Wi30vHCxGtcAVJKdAniDkAd19r5mIkKDnCB3
siv6EeWh4kByCsUd53EOG1yKbJNXzv/fd4clv46YbQUkjiw9xZMM8jZ0V45+uG30JcYytXxOgX43
WkSuhMa3So1tibTExsMJj2JSsyF4etzP9Vq5mkZfPSV1cODVXQ0pvPSf4vyXuiRb2qrbJa1pCukY
7pssBf3M8c5i/Xg0wGtwYfMw2QtHsR3V06TilqkWGklu/nEFc9nbm8fY9ZTIMI/gV2Jcsfvn/ZWI
KgBV7kSQdjXw4XGf5CTpvrtYHLT9TY1VLleS4HC1c3rJ9SBA6ulnOz2XGA8CQFxpmutZaoI9HgFp
xMPj6/9g4UrU/lowZksXnGMSg/nfEgAb6Dy0YqJfqOyGMn1y5nrvIJ3iwLfU1f5KTXALVOGRyc/X
qzRzWcrecp8Ld3eNExSDSRC5xgaxM/OC7ST2mY2jzEvi6CIsRoxSrlGVPcDoI8QpCITiolkvDGcC
7xLoVILh+1O7zondxMb7lkfz+FGk7Sz4pqLTtNbZOAHf9biYkyx9X1rxwUG5S2qyfPKfFmzjr9bB
u4bLaguiuOId1mijZeUK34G0KCghlNT+CPdMAryRnQ8+jL5VMARlcR7qKIFE4YnZbFKZgmlnp/+P
TZzsdyDVQrkFDdwoq8VrwBtEz7BBZr3NUMZPNEkjvROs+fhPG2tyJCxy+QrgnDF1O2Is6YZjt+YZ
vmkkRxVXfWjPkObrrUG4Ean7YcPi5O8kXvTZyU33LPdDVgisVqUx55RqlFeo0NcPEYYustmu1tPz
UdGireEZxLtVugm/TymN0HcD8rCSAPlvqkITa2eOUsaE9BNyXHyAMpSzHFXWJcR8zcZVv+W1rtt1
fdtYvVKBxXWTXQ9zNQ5pyxE+adpsESBi8mODAxX55f40+y6hCzsNhocOAqQ51YJqmWrxe0Y7g7Gn
ZxrgFmBvp42pDQSFrbqB5moteVFIrxQIdU3vDhHD4nc8hsSGqTcPnVzm4FKft4kut6zjMZt8tqNI
P+ehygVg/ZK4OBeHHMco8/zMI/WAKD2qJvuyRriG+AVyRdG/G4ANiKP5h5gIsqXE+eeUWy10ySgA
RXOKoTO5T8Dzepd6uexOwmzZWpo5fihsDvm8yTpTtPfmyXE2yzhrlN9kKdJ/Pdn0fx/2uJFTI57u
t+t9Tyw8tEwoABSq0WieKMhsL4amTN3O+PtNVT3NUy1/ffUqzvsNqspmjeynZ1trLz80Bu5o95ma
T+iDBUAbrFN/wJ9kvPPRo6aWL6MNavZNVdKr/c4r6NXcOPWTH2YtVWJZ7QmSXCjPx9kS5WP6SdJJ
8bhKOPwvJwEOnz/X+XvCBIGVCrOR/lw4NAFRHvJBMjLIcfUCWaoo9BKSzJS91/yOvp39Z+Sh3oVN
BIHvcncKpUyoc7+eoKZao5k2i+S7ssGbyImRu8KMFsQBzCgfh0zZDYqWOJW317JO5vrQnEB0rZIr
1/bLk6tJXQjaHYCCs4bcC80UuhMX4L+S3XIzTIu2OPHMUHhyENi0T7I7/9hi5WYVNzq8/QkF5z0q
bxpD4DvQGx2cAJbfR4ENcnC1L3uj4MWchETZXcr6XFoXH4cP0UvTUtBaGtdu+P2kWMTOklFxrw+x
wiYahU/Hz2hrbMOxVkmV7nPG+TGBgkFHtsR0xsW8LtLZpyfk0LnSccDCR9arMQ4HhssyOaAY7u14
+AM6EHL9CH9LOyOJIZDp9RltKqGfjl3SjIpEZaNLkYconpXYkgB5YoSLNzmlqoetOMWcdz+V2iDf
oi4Xtkn/zBQTbWHQTlKSPjZAPcYZoNzmyn1PvzNAt4XsXrLbBdfx9ZhwaDtIorhEX+Ibsors8f/E
mdHM4W8T3cdGs6tAGjxKvG3bAMWbxmv7G7tQgT+bFkHeBFcnpLt6tZi8Eg/Dr4Fgi20y0If1eC6j
yA43Gy6yct6l7/s2MKO9XUqIxP18Hjw1znfZ2yjDhMQcX65h/cM9YbPF76s8nSZweDhfNaXyWbpd
y+Xp2meJyvXvlfnYYNK2u1J9wBjEtWlCNEl5heSgVgPBItD6i4BSLXCZwoqq8I53Qa45NRkqibEe
loETCDc2zOmJhhBxRLvFjJiRDXzO6tPp9JEvJzNDOtwSO8y46akQ2WxlNjmIepoYsiF55NGFDw/M
bqBjS1L3jT7QSs9+71PhPMGb7cvshr5KEpxZANCbYZPkS8jnysUwfBuZpskTtAiqYuG3u+Rv3rw9
ePelL4dEhuH5polgJCX7t+YQFARUdVwDtNbQ8u1mRLVWmfZRQZQx/0lVurvRM3xk6wCjyVcmwLWB
sZZXp7os46qpwzOzBSuGHvHQWUaSzXoW/zx5zEu6z8aEQ17qhaMJnwLQXtxCCACi0bVjBtYhvDOu
CCDVFBvLJ85RhILF/OBn9RjXS7Ocf/KctmEcOmuL6zbg6QMX+KAZZV5jHVX/gAWpq5rf8NsiqJY3
YclM/Knf5FbQxd23wLRFyKz3YXFC38keCFeclqI4bRIQJpM01gHxtMc2E0gSov9gpT1O5ZNROHF3
ySxsLxWROZMUKs47fQp+lc2lgWYbPc1F+Yf958I01bYk4IEX71zGqvPbiANr35FhFqRmF5/chxO8
6jWXbgywIk93n6USvkc0dFMMLRz7XbQC6jr+5Q6NJH6KI1j21nb87dfnA3kgJaAZzsp3Ul7p9ZB1
ZXXHCJUZh/Pw06hQZ1x2qemtfiLVhGWEsdzKqdbVHpuliSRowHFllH3vcwjz75DTe3bqWAf9FPHp
ZePWRjXdjT2oUiZNkj8ZxOfpVvm/RFsNtRPFlhU32XggFZpeOUUlPn5FVp51O5OCKp8oeDcYLYyD
40MLW4RixniaKAc1v/333GiG6+cC7M7YtxBK/yMKc0OCIdZbYSxWk5OoNaxAncMVFbqQPQqhYXok
LkQOHs0/iI+/BJqpqJ3WU1gvv6nSuRj3BXFWt345LY5snzvUdHOdQE6SkqHY3O77q77tErtgWpbY
v8FrAAgqAMRlqXoxWzvCOZFG1rC6TIlclLQL47CNAm8USskMXIkL2UjUF/dq0A+M98p9h6q5y+eN
39eJ5HjbjdFZkgzLrNf27UGz9ARyM+PWT+BfUBU5Y9WGB03rUGuZiJ+mrJaGRtVSaWNq90GyFccT
r9rBdBX6dyFO7Tp9n7RtYXzT1nXtHlaWVKGf+t+eZVRj6gZMmSRcIA04tc6v4Q5e68XhKQLE4aKV
MfSmfxEY5g74PBfY293tqdbiylPcLPs+Z0vkL3Rqa66K/GUXDY1os4TviXDUjfRP37T+WNRGfxJW
FRG4tbFDK9HI21UlFrCW9zgzTPC5Z6tnTXYSKi+M4JYlZMmVgCIhf2rwe9PWgXPO3/N82riVvARL
jFPJ8eaGetoNHGqxfvNXlHNuvSlC4ypBQDBKca03DCCNc3UXTUIsEPunfKxPmS5u2ONabT6kerfg
BLSrF1Rt3m1EJXTetvH9/rzCpfudj9iyMsfwO2D6GujDAn2P93gldVboxZ3ryDI9I0VHHxEXIQTU
N7a/M+zRkgDxRFlxjqxlq5RN8/2tFZquP8a6Jsz1Mvr/obLS5TncD4KPfE1HTRJAocTnQIPvAYr5
0bdWPFLqaWVOTNzb0iLsUGnWhzMYbv6leHp/6Q43hBBP0pQKoPGlfTvL9dmXFcK+VjC7EHinw/W/
AnaiaIZakQ+zBuLDnEIfc92si1Mwe9+v8aUvtcKKs4+9+2Xi98gY616DE03qDYhxijkKqTQJt/vi
dzG8o9HidOsDZuQ/C0jkteY9M6uUo/PqoMQ77aH/i305XJV2e/+gXUkFRwgOBud0iYx1UruG2vPG
lQD5GcvEXH1BELjjklMHt6+fLvL/B/yoRcA+nU98/TdL8SsJqu4TsYoSf111eoqH7yR0r8sKFNrn
dYMepMxlz3NNZ6lZggFRhdi+VAPLsSFPmpULaS6Q0pxNAk4x+qOBIaZSXXHM8HVAXIjX5TzO1tEp
pYHuQajcKyjVtGttvl8GzDXCMjbAkEuYrJSNl1ccHYx+Di38df/8V9KWV+uQcTWWHt8Vak8qKWi0
QQQbkoUx346MhVMpyVdYpx5D1CN6s7T46YBHQS0WkkX1BgyEFBoL3G3+SuzRaxyv2XT83RT/Cbwl
aURs5Io9dfhe8eUtC6z6w/XKG6ngkN7s9i4tx5KlX3sETnN9GNvJS7WLlhHrxETidwEAkIwtvzI0
GY8ur4mp8R4y6y5MHzKiWMe+AvejtMrZzUG4upzkDo/9gNTAgM/yk9lG6w8fBmEJ46+WOIMOPexK
Rb/c/Li7B8vkcywVi0j/7CYDO2ZSe38YPGGLHiHzAdmpyTmODoSnHGEL7YQLo12adr0XjSKF87A6
OoGEzWynWnH7h4+DQt7DMb7nTZW2xOrCARMUUdZdtpzg+0x5W/1/nKtDPHHDfKD8Nw5nTKtVC56c
c9KIPWz8ZApegFgJuX4dLJkYx/Ds42H1YbmwEDih5hdWjpc8EXeOPS/GszMBFrG8d/lXXdOOd5C5
ORISDPssyhJ6YLYtSSrHZSp7TSYkp1Ahi+eOXxnfs9RJpE69qhct7NYc9KKm2h9b/P8Iw/K5Pz/i
ait7DfNBIWJ6gvzMpVpxYTDhPxIu5suCqYEeEKVNPyilG3cQJ04qLut4RhowbR4mzeVzyxmDNMWc
Dhe/OKq7OkB0WVZeNA0iuh1qtVKQ94+l9tsaNy+o23btFkGZRewbxe8f5ZRjka93eVRovFeTwlBi
GvCsUQNnsJHOGhclTp2Fm/Mh5sxzQM+HyczRX/n6JL902jNnllEIJBOrVc4v9PtXF+hTIfLZr9WZ
Oswu8koqV/Aejf9Me8w+FVxuwlO60oh1sWrcaY2H3SvrV8MmdSxolMkG0+UeP2vquvdOVaRpDrUB
hrGHPl8VIwuCMw0BsW7u6i1KnFlB5mwnk/V/YykDbPpIycEJ4OD+PLUKo29TdEggB8HzcyM5OBXX
PzOYqFPkDK9FUx82HmIgo23T7zZ5VPvST1Zt38B+R0MpNEwMoVJyiVg5SC8JHvPEHoV5FZK/uZOy
DYAKgKFAH8NoHMQoXmXK+ekdrWpSd/p22wZoGAXYiAMUCq/bijkv5c1dnmu0tqXPQuAcJ19PvPqu
JMwda2WNMLd+iul8qpnq1wlpW8AZO50B/oGEzrfUGLEAeq2SlED+KOlmT6PEvI8bAaOIiQVslf74
mktDYPyOGCu11lAN/jcd6tuDVs2yjn7vUuj7kW0G+JLSUy3I19TpqZk+FWAYjIT4MYRM39mZ3Uq/
e1sB0vijPz+Qw7KddS62FzpdfVoqxiOND1EMLpUzcJr4+a/heBm4GLWLfh2V6TEwN812vL9RlJJI
5g2b8cwCHwZQCtKlO8pr6metDe6RAc2Dg5KjhhvMCMllySGdyzq/tbwM2tYuF2H47pXrDetxZeHz
n9Wt0pIijRyI/M+J+GaCeiKOD5kdiY6aONCd4BuaF/OTk9p1sDN5C95vXkMEwGEB99cc+Ra4RhWW
B3f/taRYUBcUi86CGT/vQ5q9duGTnm1YAHXWO5aA6zVQDoymuv5E59xvMGzQTvwiXbX+i1byDILL
PraL2rAgQN+MI3IbC4iSGW4xsqZ5pAeiF1i2m+mKSsq2LCmSyAFx4MmWWw65V5m1mHLNCTm6bIyM
jFguJOZ00hUpN1TGDyawYD44YdqG74KKjIcUpLeb9YD8TTg3VMHtmZy3A3aW3JatgS3bT0LB3TN6
r2OOvaee/DKjQmDRV4U+qt27j9MZfQA2U9zfKo6b3DQg+hn4cZ/UM/JIyR4PzFg1LzBVCV9fKUlP
8CCAndrRlWlqMYBRzM7nWXml18iM/YjuGL79mDv5XJP7WmX2CSLAzox3ON6atBcSTPFdjiriRF/e
KfsXtEQom58h+ERJf/eZbjXY9Da+sOHhhvukjn8V/MAwDZjEUv0qFfIMbJxwfWZ9Mlhr17nrvMsT
CSQnTC3WUXv9wY0nQCuI0+WOAxed+cM9I6g7+pCkjzhcRGIE77opT5S/Bd8EVo8oYIxFdO25gP/0
NfmL6jzAaot6jqDc1yRgYkgc94/NR3jhjLpyCYctXdKpy0GT5C+TZ5Z+qmmuNMLIJI9RAYskGwBw
2fpq4aKrOt4REYSFrKUn+TRIFo8G+/b4iv1FTxiOwV37h5BOuGO755NQNgWf8UA9Trtg6l/fu+Ww
zbbcTiLPPToLVOXxPn2fziuql83fWaTe7gis54GWqsdgk27ys2WFWHHCcDpJpaKbDzudya+VQd6y
SwuwbK9sbKtacLq2isdkD/OE3viQxNLVXIj8EuKUSVQUeolwv7ZvE49+Zin70l/RDDecgEjp3P/Z
FBc9N+7TeOr+GP+MbQumS1fN5wW7edZxomHQ1kRKoQM5+S3Es0ttTtIXreLPTgCjvla6jBr29BDb
VosEjhqlW54i53jeEKXV1ImucsF+Aup4jKfW4lcSoV/23OG25mKgDkRiuIV6KAFyQdfXg1g/b2aO
tTkEJSr++CgmefnXPyDL3PDmcnTT8KAevx+5cp6Gyizre8wDaxpz23OlsQWxChS5NIyXORFqzrpc
/UaPLqoNlKsyh78u4qD3kI1Wmnwnv14byXGAA4bJZTOV9mkIRzqwdDfuK+gS9XAxHbZikWKTBE2A
aBVG+FTlRoigWn05N2F/tl99xHaGbSWHBBGb92EmFlah8NmpPN34o+StPwLjzUTGfdYqqV+H29NO
W4iHd3xieoIN9G5z37IyZ0k0jnvSokbHRm3ZTZHDzMATythBp7xjbH3wG46MJ7Ohg5I04/Pk9vp8
IgGwtisncrVx/NI/0ySQ+80tE/CyFqlZEFxLHvd1L+D/VU0dE38WqLzrxk1sM94MP6bskVXxJbcm
Ko0PKpF2NzKq+wP5d685bUhyJjdlm63tO1NqNM42y6x54dBTZd2Y2wprMHlK9vqFMMEVOwUg4T4x
EfPJHG3ebwnzGe039xGMrVa4DKSvO27nubjRQbwSLahtYXxx0QnISZpXnxtpqtP6fHJLfoV3pwcT
/RTRulCWuSWF9c+SlJ+gdiQGSO2Ceo2S/qvNXBsMNpIfxMWqPDnyMhz2RrMD8KTivpClYjGmTsFo
aZLD/cMNiDT1lSpdFyCEjFakvGg9o5bDpVYFTVsrE9SwbT0XpzJAWZzm6hAqwY92BxIRqSanJE1p
xf+0mv7mJujM3vU9fd3hf7BjBMB843NwJ2T9VJ4ITN1LWYrq2S5S5RLd6pAUj3vDS512RoJ3GDQY
v/YO31iH75LOjaFpbEBZsdNjGOxJqmxmCnJgUizo4a7oku7UmfXMmsDE/gUzpDKen5u0r9Jjyja5
VKU9GsvDaTwhFg8w+oqrwKPn8/VJ9HIU9JU+4EBxZRNtG9yn/tPcdxSHxo91ytg/tOaiNiZ22/rN
mBv5exo+q6hzegYvioCnxUZJHhH6172Sir2wx6gU3zmRa7dx9jNRUSPP+5yj8CouK4hMbtuHu3DO
X1mCcHKyV6ShdDQcIvxjLLpX1huU4wMVxe3Enrw6Bmnvjr9Fcxd3DG72cspWx3VoyFiJqvlS17JV
lFvgJRohjaX6q/AtqagI6rqvQu4DDnGefc2hNdl5tD4OR00J+rqoFeyfJsNv/3nMO2d7mGOLnwjU
UcHdwnkKIzq4pwNLxQVJngab03ue7OPZFRdQXwbYMWXIiKb81ZwJ+SQmfXT4jK6BsCv6wQkulsbY
6lWDs66g09f/HzQ+YvBwFx6lVGMDWPZFIigpltpiosi6T0mpo0dSEN8XGHQvbEQ2c5DACTjm46j0
vMqnYXcfOgI09XcotAGdTDEUDRrlr0IFvMCYolaFb/PIl+Vzq1HB1MNDG8FsQeeUoa8C6KbqL/at
7o+LUJmhsUyzO9WANj0LU2XRXVvsUkhqcruJspbqAw9oBtXBKzMop3Qw07w8DTwPo27wsFXU2KKL
UqNgizMd8GsBHdc06w49pE5wkhBRieil7DKVA9xyYVDf38tqkBCcEIRT5MK3+sJT9cZ1EoCcXHuM
CwWy7mfuB7zA4/lhxsYOHylO5UIVOzo/Ov1PsPj5CHaUhrQUMPtj3Tba1BdcA3M81aKeCIhopi/0
aXxV8rVo5GMLGnBHz3sjtTYCNB5mHY9kxs3EZ2DBJAr5ybpZj7JZMoVtHIPl1PVR/LO+pTbKuuq9
Idw93gFoAIwruUfTloiGhQCaLXTC21hqsQulzG1SvdYkGp5szi9SItTwwokz9ViWCKqXE4P2YMtd
dKGy4qe+Ou7KqaWVEpFOywpmEkE/wvaUq9XgQO47IW1Y6Km4PjjJ4HygUrarROlDeUYaCA5i8DCW
DKMjdNmPQiAXHSZ/x6CY88rtxZu2lz8F9vtCRlcKB3DuIGdTFdCaKLh8zuIJKKMLq9pJQC8IeMGZ
FeTjzqbYBxCCNKm8VEB67CH/xp+6ebW2vRXH6/ocxKhWJtubEGMyqlg5RSpO5x6D0kDK4I2HxREo
3NUO7XtC01cBgc837VB9i8gwuSqCrrDNK2M1CQ/T9xCne2y+ZW9ru07NXlZHV/nch7MuSepbemWK
RWA3RO7ppQKRgHJgXwtPcGA/sb02ZE6y7iflhzvDMI+Po+rf8wOgSFG9BZqmdlIv6tPbR8rhH1Q+
NguFyoJKUVML4+dmQ8hy7LmRTT1WATkIoA5mnIAuXAhoYlYrGp3dUq0xPs+a8nfsiYlHCsxLSgYe
IsM+xOR9fc8OjuebbjtJA4GDqXr07e4g5th88g3CfRL+AJKJxvFdEuXjY2l1Sp8mrP/+ctFbY6YM
sH4K7M0CWPP29kf4fnBCoKj9LRw01GxvUa7wfClMgsIWQlz9eiIVgXBGprBCT1t7qxQ1IQjuoWQJ
FtcB0cY5FNqioMbuKDjiUpJLwtk9FK4MlJdra6xbrpi21opBcvmzAstRergjtNHB8sULYpodF03A
8LO/FxMRINBNmhshVMlGTRLxU/AijJDv+gneUotky1br/RAVWQNp7KhFaWjKAdNX5vieQ0+KAxSo
x/7eka2VT2pQBUdoEiEwxvr1bKBBydakXZg2hFJbvXA/Af6rnojJU35QMpzhkEqxo2FFt9tvy0yR
7J9JxcxmqeN3MJtHcW3S24kXsuOT/TiRW/RZT0ruSW43BIqkzz3BoMAxp3quZtoNkI0M8AgolQAY
5nHIThGmYiJ/v/qWEr9Vv735SV4HuwP0ZTjTwONexWFm7VqilttrLs/NVKqrTBvewJhn9IcxYvO5
D/Efm3TgYWcA+f7JRp+MJVY6iTzQblGHMN0BIpRw2rOFU56T+SCEnp6OWob00l7Rue/FM1J9lid4
rqj6Aes5fvAPDcjV0eztySVc9gl8Iu/A8bED7C4KmV8+ZH8QEr728QULDcclwYOAjpd5CWUQCzQe
CbsaG9S3Jn7dupwG/cIP/l92z6RcRDaaNDQQ2/pvW/zMOYk0Vy/ZkVBIFcafqEWie0KIWfTCtlBv
D6Cd3mJw5raaVCjRr2LF8e/7Y2upeUfYBxGj05iYKiMZhXBoOGT5NSB8jxPgR/PAO6zu0cK7sQuD
sEpUiOXon14/hjOTzhLLBuT3nWOacuj3nRBrJR5rYXvywSZE9Vsj6g0TpgCITfRtHIePfPvX1X6v
MxCKsk+Yt2LZSgCg1lSZA1zO149iwPq16vRQzdG7K7sItmcevOk0PE/nLa8/EDqAbgUPcj1yvxb3
03kaW+Iimo1soUNtSow7EcsbjY0qdyx53/Lmrrn/DC6vWVz3faAOdO/3I7f3ahGBu5w5UUHTLSS+
FDuRrQltayLFMjoxxziRhs+33WV1aZAdw33PdTerO8b+W52js5DWmI2LEDZzW9/noUr/tPbk53xN
/Zno0h43oXXFKgVueFSqFPz2axOZRUPX3lH7G0FCeKq7/5XF9sUILpixoAjKUTW+KoV/Z/Py0ltu
ldLL7T7Oxf2hVf46Gb3gJnbVVHKSK8MgDBvnkGe4LjUBAnCvCZjnZfyp1G8GlV6fRMlVYOU9eTWF
tgeJ128jm2rhvsm99RzZohdnlxceRJv+4nnTR3W/Xst7WzATQZk71PU8tLeMZZs5Esb8LRuTFXJW
wMd246s5u8fh9LN8X/p5cqfzzjZ/LLXw44sj5SmcRIKOnKQlp8W4qdnyYGINs52oAA/sFnUFCtop
M0KP8JR346zs2O8ZNJ/oDVTVNBZpbZQdJNJLvnGwQorYyNtHMEUyGoE31iIoELku4UzUnGr1YjB2
mWsRpc+JWZ2/tePILGjxMihCfNlzABPgE3Eg8QhQMHy82GuB8dxOnhozm6oleFbqUa/pcZRbS5Em
T/NEoWBeyfa07yCRhGMLBfNBhgxO3+tVw6j3WelMIXQAFOulHyVqcRcXr3QsdsF6lrWl9/Bs9oaN
1SVM/2tiX8E/St/0O4G52ITr7euJRkSDTFNaOfemrwVm+/qtiUVf7NAl8+Oo8g5KsbmATkeuxOEc
TUzKLpTL83Sa87cxLSpF9n2OqwTD5b5ZcH2r4wRnr5OhgZJfTAfMsocxupdPGggoxR5v9doRYngT
Gc0dpVO91YGpCHTHW0ChAtIa1iYQYp9ggn8qQo/UJyZSnIQGGDaVHISnEHpwhkc4REJ/aM0RT/iA
vgC7v2R1MdA8PvUXCyMcuGMnBgkA2jjfVJCCxD7B+mJ6ZiAjtAuGJQUq7+Oa58NriSfy2kkr6S/m
gVHOAcbxvvQ2lHSIXJ8xuQOYVMFgbF27vNzybuWlg4kIkK1GKGoFO/JQnXKx1eT1jw9em8+9PHMQ
sBRo+paQwhXvUiNv+UUmiIwIAi93T0Lfltcy3ecPSL63H53GLrM2OQ7STRllH3WEIiCC1xCjY9Yj
kaZoOtR5DgfYZ/eaXY4zGh2uyPuQHndiWyPkPf19Ws4UW0P9BBnzQPMtFwAw0dt9HM212hx645BZ
ZnEMDzi3qNW8SqlCCesfSw0+RhljuNOKZ6eI9n30ohe6y0KK6aN1w2w0rQ82yDMhmq6C1LzEQ2fq
RDuJYm2iZ+4/+/Rk4GjbM9Spv1A6Uy7ooSMg7I9dMvanGhYnF9USMpQVWy1CDB004YXJ5Vt57kqA
h2ETgtQlwFnoTUfSht7nb3Sp2eLG4RLHqgklqyXxl6AekEziwaGPATEqjzxOpchBc99wOT4GS+4q
SqgGDU2ixDrAeysMNXAyVCpvB2UMZ+xfQ4cjI6rCWWJgXoURbyY3d6oXLT/jWzgZcP6vvTYO1nN1
lA66P9Q8IqjyrxT4B8Cja5hCav/kdX3V7SaoK7wgQ2DvEJd9ydA4XpDupWHBzu7L1pGgLdDsitJ9
8g2a+0hXupIkoC4vRz+YJ2wyIzveKUdDrtPyJFBLxZy3kskcvVeFIDisFtKV8+K/KxB/z8qLZnP4
eQEHQjuTBM2RV0yvMrq+5+ieSdTJHnC0oFYrYnUA0iLRu1hQKd541leToDo0TmZrHaGCkDFjjshH
u+lNc39M8kIROPbJoFjE8Q/i+JzNJGx+Ax5G8tISC7CUnQqiSq+pwNSbsTXFiZ5lQXPy+YPubgj/
m+E2JgWcnMnZvBKcMf1csnohT+IRxnuneAwjQ6DGvJyKupjWOT/oFl6bHRyYSoiPH/c9JqnZoHqx
0zPuv3XuLI5/tU1SyaLO680XmAotj9OBK9pxCpHrXqN3tLmbp0uBCwYVGmzoxUyk20W9rGlc9PXI
4w0Ku6NpSNTwagT4RKfIP6U7eTduAYGW91L+ysH1n6qb1ZU8acgY4pVyNzocNT6NhI7eyEmJyQo1
n9QDCCxj6JvmyY1P8TkMsm4fVDekFlJ3qXMt0Ozq4o3jfND8qciaC3p9bSonBtac9n3xy+J+6le1
y6mHvLcE50NxtG+I92zeuP8KlCt28Gftks8lSe3ENPlHjhduKp3F1tCDVcJ0hyV5ayIBaBkZBenn
B83434YPkNyqoFnQ3KHiDrRirlFguP4ncqmXh/Oe/IwNnqRX7bPf+zaEOFoB6N8pX71zvuSZha14
+X5nSczi3fDl+ga9HBIKDkQhTSAWyzv6afHguA+ptcWe88HpIISqesRDUTgntToRQcXRlpyk7NZK
l7kQkxbK1kATyH5Aj3jIj+cfT/sZdGgrPDUmRP34URNJmXYdEqXxtEUExG6gQJuy8Zjg/KgxNvx+
TA65yDzBHSuu2glFT0j4Ub28yHPee10vVD3WFefqrehNR2WQqIDTR2CJ5W5K+EYYwBhryKmBWE8f
MvOBkhOzWFhK0Kn1cDvUHNOjxKZogzhF6lIpMHt5WkPqzKrJL1wnKdTBLWWD+Ek3s7blI2pOlwgI
wCVeP+WhCasAgIYm6TVsfem4ygKQ4Xa3JsF2bHD7NQtLYNz690mugsbBONrOs0ZnMpgJX33G5qUO
ndLxNpZqY4w6uMR4p3kgt7646e0YvhKb05HLTLNKazLASvuSpO8s/Q9iIi4I98nJ+L0N2XuNSUKq
p8YiEMGfzUkpAS20dpwhh/CHxgqLU0DKhToAjTnJHXZyMWU0/uzD/idp4km8/m3YuEGo4kUXkxlV
HKUbZmNpfVsF/eaJi5gf+51qrbRm3DAHKVM2SZn4mxyHK0uSRE/vLa+NexRhXfIWVrX2qMpsAXOM
47VnI8Xgqq93mAKI7VVsZEgTBhREGeWTNZZ/PdghM/F6kZxHPp8Dv1QbNM2Zk31rhAi+b2/YScQk
TBWT8xm/Bb8+IdNrrdjvqGM21FajREwaOOkzXJV9lsg6cZTle1nAZLlFOIFbmHcHtx8XG1K4qAFx
oaSPnNR0nZfhjRxNbsEl0R6RnFuYKertk141lZ53/mz897SUKwkITT+viu9WoK5rcUJAakd0hqp/
E47YZog7meIU+XD+kktDtGOHxERNSq4n/OjfjPbeYyJ7HSDKPeXgXnGC5nLRJeUByrMAa+oT5+R9
D6kDNSU+ztXet8lN1GTnbtks42DfMUna5ZUZ3cfS6jWnVbiDfTdR99sd5QOIzFZMH9UP4D8IG0L9
kfjOEzgjXwcxeMPxObfUgym6nFMkVyGAHaJSNL1NGkWi0mbBUZI2QVNCUeW9kZQFjwilgNXM+pL+
+VsydmZO5R0lu/jHRqnx4YIIiO2MhSmHW6pg4EFsBY3nN4ori2EfUOV4YFbi/zzPYu5BLQJKHj54
9GEMTVBw3tGGgnIar+O5LXokt+wVEF6VDlPzDOMYfnM/dgvxe0L3Pt4LX6F22zm7MGuUthJU7J8V
xqAbaetNFk4L3Gdr3FRPovaqO3R0ao6UUhHl3bWxbb06f38YmKqwHWiREz+fkxjff+vXflE66G8U
AE54bfKVIQrZF5VDDH69OVs/EWxJP8RXuWnXrJlJ9EdScq8v538kknL1me/B8Wr8Ln0BuodU2Fx8
l0RGqxnOBjWGHkIbDYk5hpVXtGgGHDJqXtR4kO6HtKGDfmD1RkGm6aDpRuXrnO235Zn3TegrWFGW
Q3FjnVogcv1Uj4LrQ4WMCrEJfL6J8l5GO6qtn0S7mmcBZi+t3Eg6asbO8xLYZmArvnExS80zPjoE
3+RB4ZoAEmFkV+LvtT5TpZvjLhnMCuwre0p1hhcFEQ0OxlWvfFrAbOUSYFNxDnWFxDTzjMAL71YB
C3uTnUlIuV1GMXLGjPf9vyl+PxWLMdPnTot+EAAGkUc08PzWhDtXYGmM77OzYtHKAdAi0Ib42PX2
xEZY7RVd2Fy1oivikz7s2SaLSMmtWfRu7slXB2SoqZ9ELm++1WE2InfXkAxdxEjJ75ZqO8kT8t92
9uytrfKWl8krhU0tiy1porCEkXbVyYyZuyUROIzjxfYhVrbjG4jeANzjpoSQWzlCljtfeG/vnoHi
BUw2abVwnYPc+t7pcPzpnziaZcYRJ6kq1QakC/+HG1h8pGd0bP2GbjHp7imdrHWU3mgmF/nQ77QD
yAxoOt+GrmyiJIy2ZiW5BQ2/gZ9y4Pj8ANoIcyJFW7l13Gzn2BgZNkpOfzVJOwblvdbVirb2rS9N
OV1bA9KnpemhP3ski2Tl0gD1OQhJH/XUOLIAzkOY6D2NwiDf5Hc9ZkvELkOxHLQyRq+JrPI+HC2L
dmtYyq4x4XWkaY3XB2XDeqQbtZAYztUFVG17fuZU8XaCGFvdLLa5O8azrigLAQfvaA3uYqHGgmoQ
jopkHtexSXHC2oyHqyo7gvk/sriBerPvs1mh4V/f9LrBXS+P/K9qiVxPIUy/siMumOWKSoslf7WN
GMfsn6gnMzkRqHgi0Ydsx/6th9wpArRTXIxjRoJ6LWNYdm0QP0TH/97EpRbcnS+NePjvJQstLTPU
jrXUfZ6dgte20whV6/KzTkFbdq4go6cO8H+aK9hyluAa15trl4Bz1mo9jxYbN81MjG+ki+xfjH+3
vclFhsnIn7K868KHfnxMTAysp/34sNiKKXM9rxDesIjZgLr4fSFZdTO/93KBvtWvHE4ahdW+ZlOI
tUNRAqb2GrWN1ZB7mB3irdsd0ECgxVBG4js0supm146JtzmFFH989ktmU8hBeoIhUHspoQ/qb7MC
OmblnxP11EyCa0OxIMuUr0Lj0E88XesS6tYybQKMFJEriq2LhvfCpmiH8SUZA+myY+9gW/H602mK
rmjQIWP84OgJAS5SFkiOcw/8s81DOu34Ze1tehuNBcHuO2gIL2gPuluHGNK/zqXfz+m7z6g83INh
U8wcRib0ufH9S/pvQKQLaETIjRXYRAEs5r1uUm7CUwTytb0tCf0K3eqJ7RJaM3Jh5ZGagqvImGD9
ecpq1gDF3xM80r8p2S4t/HMO7Te8xyeFiilvvfthZ+6ILim3FW0lySIT9hDykCcqwY66jcfZ5R+y
1DXAGR8Ix3MEaqdhzuDkpF0D8q6y1DKjBnSMS6yAZlHLPhuDLYQyvqqSqpPy2DTnMYjPRsLKCuKX
vxGvIRQsfwH06MR8280IUaE0lg4JsnE9+sPnAwmuOd3kC1+Tf36WTY909Ha68oHEwD3vADsAdu+u
m45TOgnwIno574n4n+GUKfO7QJ4HhAruRnEkLQuN8R/G/eR16p4R6LYxjRhYAtzVYb0pKqny8ZTU
qzrdA8MKV3KMrRzWohzOFMr65fdlfCNlepY4DyE645St9890BN5M6CbQ3QtN+GlrDZjF9eWLrQU/
eAM9QQZb0kjQgVZPZISaPEKWb/MHOK4l67AsQp1kJHpV+EZz4nvfNfhcYiEkhIO18A0pq5GfzYdw
in1wNQdnTygLqoR+EaP4sp/6ZGGt8+aoFCdpa2RK4H4nD3JGrBWmDbz6xstKpKzj3caTS0takTkW
n2+5XtaFV5LmaSjpyTXQ8LH+Xk8IOpMN1Z9rxbPmk53Ci6vqNLU6+xiKQa+/S4hmcvtT/XIWH5UU
PWx+W0U0G+NJVnl0OOPx1A3WhaFI3+U31E5LgHA+DcfqncihVHDcgE+vP+DtdYwaBPM4jMGGu2aO
SbD+Xn9UIV68wBE2DtGyYuP4M4Ju1wz/RSCdTEcvJ3+P48ePgmr0x2NY4TkDvNfugBxzkYTniky2
55Drk6SJWCBhkQmXi/5lj5lVBDsztf510RC6Nerr36QWF8EtG7O3ghZekk6UjOaOu6cJEsA3O1dA
UW/Fba5VBXgfN4ArmPoV0dGi3Yoc3LqAj5ofxXaSkMKyTziLr/7/k0Kg6OQNzt9qNcll12vjUG7a
Q4Ibt9q1Sh3henFzGIP8GGdQz8lGt9qVor5oE6z1mePFgkYKgwogmb1bGKdT/HptXhPFn9da4n2H
Sj/p7qkXR0DLAjwIhmR4G1g0wgn9M2vhLhyjg7wtoPo3SvsrwRVsknFZXUqHbiCqNlp2zIGMEKwz
DrbMjXpf5vT0o9yHVgFrEQM2x/MfESYIpaVWVze4gHnX38oWzxSGVAd197e+Qi47EOIdlMBYzEng
SKPYfLMLrjHxU5+gByc1n5YYQv/lUa3HZeloCYv+JqI+HFex9CGtIl6AsoL3V8mpStpAHoSJVbdj
7NWoh48K95TVexoV6zCjplZQ2RpuampWJY+/mDqb+DPMEm8z26QxvrUbUJgqtIux6OeHEKcqiMTa
b/UL01Ds5rnd6+iyGZcnHocPHy0xZTJtjkqh0nQ8e+CIq5MYyGo8SAKgDo4+/+2QJxkOyvC8xV9Z
My1omynV4xaRCISzFAvoA46xbPQSOzzB+2q9NPO8x6Mz0OkhC+ccvPrQq+zSyXd9Q5DWK4lAlZ6I
GqfXniqQ/kdm5AOAEhUFIL5zlSM0z/59iPlWdNKzFKVV92Ye+Ldo3RsW/yGHZaitchFpG9irvj3+
Tfj5YkGniY/FNczmrsYafisJouxs5J25eRcibSaEwImZ/gX0Kgfhfhfj+MUL93vle+NM3diNhfCK
HKYfy2Ix4Askc/g+G8fdkd+/C4e3AY63fV0kiQycrF4G8uD+8P1mYLN9upqIqzVi+VHygHZhlQ5B
FnEeE0n3fLLfD7L11ArViJGkAmvne+EU7PJAmnUCXae5p+cwViebZISTIpyZhCb+eXL2c1vt6C/z
dDpN4f7Yfd9l3m4PZB97EboTtZoaC/aERKdOhjEy3kWXL0F7cArnfZZD6WJYXt1Nv3G7YlNj8vnn
M2iaWsVVmlw9lZZzqRXScd/7H8C6ynoGXivamnc9e5Wn3COCsg5kUmRRSWda19Hbbn5JMeFurTyA
7I0rJnBUf/2BAINBEqgeaUQuRLQQlM7SS8q8Gdvtb8XATCygihkt9HHRW2W/7Q14rP4GLGyOtJ+V
WaPoyWtPC8MTqKajNk/FBHG6KRkJF2jLElJ/KhZoxWhS8g4ep7L2Uv77eWQRjSq7Rl5MQEDYIsqP
IIt1SDRpQxpodRSkvZuYZM993/a/6ewRIEjonlJJVYqmp2tjXuZeOsr7/mLVIXSeyau5xxi4TcAD
/lQ6+Z9RyEKvKkF+PbeW6aFiH5S/30pq3OLfZQ+kx2MWfTuM5LrMd2n1WmzFSp7SMwYfQw1YjqPI
EtwIB70Lm3EsOZw+d1skGpoYCz/xMKGUoj1xuV+9+nFm8nV9G5f1MBmEDc4QRha25urTnC+ya0tU
61guledOn3Uj6UhwHBDCEUdk4QedMzZZRoe1pW9PcgeD1v/44FhGvMjrVwYKk8HuoNwLHcaBNNAu
wQQawweQfx9aSvBYyF14JuCeWsbrdii6/z09x/Wpd7X488AlSkaqYRfmi6+PVy2Z8BTxkphu7VDm
qUxWeMAcKlrKJwKnO0jwWq1rfqfLgaMdGOS6x+w3/ohIIW6OgH9MY3wlI3CDp9m10ukstJpFqYft
ROexiImj4wlvUrbO7R1MgjttkHwwuKdhIO2Sy/eeVT9La2VrrOtihyCARyxVApDv9Ksz0cMWxfd/
udL/d1RXU6BtMyN5DFSWDFLVft/OOu5FUGce2AwZ7bsbuCX/lKEjTR4yUBEtcTna6daFAxD5x4RH
oX5H5kPE3z1a4RfhY8kmdRbJwzySeTxxPvILZk/X3nx8OXkdBS+iB21s1+G9h4VA9OyLQ/cXJHbZ
1gb87VJaz25PLtNL67oXwbVgTSFNQ5Ia5bxG6p4WpBO0IMXShrPFE9Ts1NnoUAbPj8MCLhi4PsNU
Tofn63NN0IkmXDl+SXMuegQMsiA2e3AuJSwxT941p6/pGGLemlexddbwoklZVGoNwnBYLZupLZs+
7154wUESS4221dpGwdka8JG0c/4pbKwQWsB5rBxv8y3xGMNIcwiI4e5Sb4lYp1PTTvjlBNzgCNAZ
bwWYLfmYUM1CVGnY0Or0o5Nm/BvXg16MYpxThNeoNXbpX54/cc2EFGoDJ+aPw5DwfoOm1sdvvlEE
s8tG5MArHUTTIiFgSkHFdlIxZYAimTJ2ZDSDmTkhYM41z06tMkuRNe7zEG4p20FI1lsxFGB5mErz
rGegGKMrMsanDeK3WVjaB5K88YWXF6DblDSxNVKAh5VJRxnj/UP1OJmMW1DlCrdzF1xuzdBkAlFL
evAIOZXDOrJAiBm+Ir95t/AdyNocS3SEtkk9CULoPRl+IJPZpQQWxRsY4IXmPtlRKt8Pbprm8Tdj
j9JLfXxNCmOxtqUlnpTJJkenJkfOUSoxCNllLks4WcHpq61vZgNFve/hy6N3mMCsaxo9msRCWPWV
HpjXbJ0O+0AYg+P/djMw41KnZ1PgdKu5CGbSS0ezrSxyoMxDdZ8UI7RxmR4ISsY8wHFA0C86LT5G
J6FtCjARjxYfdzf1cYl8OfuqdxDei9BkERFhINRce41LuTekAGTPXDfucImv5zc3r5mjiLRAFAIY
SIAZoEOjnXjq/M9jWNJG+6/VYbIOY+/QGDLgV22gzzPoelGFuakpQfjTbqwZxOd3uJzUbGw2EUC/
JstWkeTmdPwvr3FFw3YNHmVU+WNsom2Mkk4ylvcPPLDMq8O0jzI4px+li6Fo4A57JV7bK3en8gSR
WoKzg6UmwAoBVQ6GgIhbGqeaaDsHJD82NHnsX8CVY74tmbJmlh3kTHkg4kaT/CVCur5o5363sLYX
gjxj0Lu87g7dqshBD1p4ohM7kecQ08yVmR8HsF37LpJ71Mvp9598AIR2AnUoSbsTwSS70fem00WK
qFjJMLAV3cU2fIZuiv8zIxQLUhPSZ/bs7JuMNu/KLpoB9snJAsI8bABZaLwelMGjy2kQFteOElMM
r4FDG+T8OFh972n9ptZQBEDWDN099drAfDLqBD/waKcRJpiKJqmJVkSTw453mg0/5iBnsAnwjyqS
aDbkGPx/QJOszYi8NVqW34LipD204bim+3wnkeOnjBYlr9DXCkzMhwTHgN29uEvjQx8Pkb4rSUsq
H68XUM/azo5K49GXZcSY+95fo2V/aaK/AWjXIKytvAxlNtRv81rgYj+Xq+RXTHZ4So2BbDXo/V5Q
ZYPPJyTLn4w4R81ZMrITirXGJbNj12zZaHxzc0AAAKPyQzofNyz3HHtDWwtFt9zjT3lgTF8XRkY0
y+6ZoD+TyyTtF3Uh9vrmfMaV7l1YMT+FAwQFtuZ1laO+sVF0HP7C6Tfz1FSQqQwlG9zb0wgO0nRX
sKYvYrYhJKFxXOyfTX7TvhlF7bIk9+s4qnUD9hODMbYY1Opwty0OvG0nHZv9IxpdQIMXP5pNNOZB
yQ6grsqaC0lyYJQvyKfa91tdENTxkUeWOrBQPdFDv8FqSbg7t9Jxf3rivKKKnygyO5S93PJJW1N0
Qd+5aaUqMjkbNxNePUuprFcYgdR8WKxCWta3UnLIBXnzAAU0WLYgiwXJVqJstJvWk4PypK2Gl4SH
wEYcl6A42yl3lZEW9o2TEkX9hHyygKsQQpoanU5dKOAThds/qAuQRBBGKOPgKKsxlcrLSYGMAYtC
bSi6dcOjaqOnIDbauvx2dmKZ5UNjjNoz9UyK7JKjlVizH+wY51yiTfgd/GKplntnlk6DyVPyXerG
66ziuu2pFcisdSH3qENP48EAUrd2pOK1/s3Yd9Qr2WkpZVdghbRWw5xfqqoTU/RhLXYC1ql6e6iY
6wJUaHw/zXA8ZVd3TLvANHut/LxAJpx78D3Y/RaMSbZOs7kHsTxPfRyoLfcd5UVWoNSRcaFspHO1
Bd4GkiKAgHCunPT9dFn0o82cEDGezNd4cV4sa0psjfYbRBaQDnF+kljdeqpDfvPyBokFUqAQBsiK
Gxh2y3K8ikOEBht+hn7RmA4keQvKoN63Qjkmj/ftnrHhSSUHirySN7EgMfqVOB5GqvIBWLFAG+LL
zqipWc8Z2eCux6XBs4Oh9UbW3FexGYJizaU0tGbmEQlUDY2PDW3eABqBfnpH8evNn6y9bCl2rI89
phblLCdkLvEEaf3fUvXW1kzMiZoYlotSDgpNKCZbJ8DPaybxomCi561mUlYiVQvltdwYnXdgs5an
UkrLXBmrWM+qZjNlYrVDTJh+U0sVfIYG7vlO0WEtuRu/DGwNBmPDZjQT4MpC+U/m71iw+ZsuJODB
GqIhA2caCtTKB8awaC9P4E2VEuFHzZTx661v7AZzn0HV7AuYRp5uzcgZzMFOy91eFqgrF5+jgKIZ
g2e4KQxudAWWZVJPSBH4XYO0j39VY55MehUa1hpnCPHn74d/6VQNTZrTxhGQgARvleGGZg3a53q6
DEyH0SD3ub3oLyZ00iJJX9I+QXa0/q0pPzwF1R61xG3pIm0tU9hNTcoj6Q0M/zsyLe3ZkgQlElxW
ZSD03g3rxeSsdZ8OhVhiw+ZHozm1ZfBkIrgkwnduDwhkNexBb6lUR2zASpJf9ouN49BkyRlBCHVg
CKObEsuDkKgdawcdBIZEH63H8rUwyi4cmyKWGQKpm0TYRtIoNprQzsUf9FlMJfXmw2aRCorfoHBm
23MTfHFzO82TPcxIcP6nXKrpQb83gfWANeytxb695tSfKVkfjyV1ed9YI82b3NZKnpg5+kkTJHJm
LM351xeLdJxn+YgB9N1bfs7S5WDbS9+gzDK2TzTmqCOgQuQw5sd2OTLRx/Wl9h60qZ311963U0W3
lkqNVOljmVJ9QwxMlapQijUC7wOx0XHJIZeLnHa87oaKWlNjtMivOyXMu8hnLfHRg4OGXJ6bGu/F
zKuz6cQxAHiOsVgYlwxPhTDNNhqxEfi1VzHArffUI44xrUN5BgIqFvYM1T4tbzpOPyxaya6SM9X7
Hsjr9RR8EQw8mpDF6u2c55tiJTwg+o5pIEB8G8VUfi0yY+D/OoBVbj9GHnsquE9dl5TQj/Q09Gmr
mSSsBTONMErmyknq9f0kfN6Lo+bMpz7hoxaojyTKUG55pemwawcYCRKXJc9lp3B5ys5+Oe7sIeIh
2KLexVP6wySabrEo220BRbqRgP8CblR+wrTud/WBao+aiLUgoGDcG8zjcM1/JivUMwsZWeTFiEYs
aQTD1/LsquX5cTrBWelMewRGHDzAoVSz2PC4Qy0a1G2B9h/faqX0yvdB1A9zWPtxwgqacZq5+0vb
1b11AZVTFcMeGWBhht3h3YIV0E+bHdzytucqDJ2wsvaZ8sUNBvy/3nmF2e6Q0eDyIPxbYZEnDEkh
TG297RbGQctwSyzzVE/4XUVTm38TG+iepTgpJjk6+4DsLRTI7aRLc5pEgsjK2FSRssV7/NCJYyyb
7JGAuQLZyqBMgFju7/yU7Riz9rO3O5oFovcZwBKpSoRTliHVv0g0zPK+rgy7rUmyJ2Em4LAUhVxj
oYWpzIt/ERIis5kXjhjdUhCM/O5hNoX/ucC9ZMbU3whgKdMYofFHTy8Om3F3nk5zkk581TiACUns
tr4K+JTks4tpwO9esz34RO2kT/zN9evMW4ibdB6XFqmnbbHB5vpYFXtb3I+nBxB/JTgBfTed4Z7g
CXQ1vJh1WGQ/Vylt0L0aDsd+vwBS64/ARO9A6xHioWrVBIBA2tuINlNnf5RqYNs2Fsye+0BqBu0E
ds5Vx0nEpDLOj4Pifje3xBHqS5Xu+6Uco1PAYky0NpWp7SJqxCL+xj3dbev0WkCZUBbeQs5wJYAX
Ud+Oc92kc0ugv74zbQDG/vFY1UNWNUuxvP1uoaVIz2jUMu2OY3ylRqJKPQICD6KVyKLFMFtRPJQz
uF+U2UdGECStbBtDZYJpB5wK1/e5SUGPw55giCIOzP37y8HIvkGyjfTkYv9zuQCiH4xt0A+983CD
xz3GsSlk/uAYx2OwelO3E72Fnv0j/s8uIhc2QNzPNKt2E9uKZl0/MZorWMj2MlsHSwKr7gG8k+oj
J847iIPoQ28cJ9djfzF5uNK1dQO/hCWxeznA1gbG6B8ijnqbXx/pwN2vF60ztYxuvTmuGDOFl4c+
1kNbUgnFjLqITCYcHx5SZX1Ji8xdsIgIeqhAjlTP+WhNNwQFEJClU5GhEMYwlBjjK1LacR1DoWNd
cZYv2FWiUNYIo5EugBuCIfek4SHnMit8lwA6uREuu4AkiLQy667i9WRvkm0dv8r0ERG2KoA6zrQH
vJpcfTL8LMOf2SrBV3qx0WTH/iXUBAKmvNPlpx8LOtmyLLdVZz+mnSr0JAWo8R2vbcMUs+MRtp+5
22rtVRboEJG9cPKMgNdHQqoYJx/o6f3rRMkaWFrceZdsflmUC/NZLB42LXeq6cEk+OdPHsBj7QKT
0SWfRAEdtAgGTZCUrbXhnAkY6HQif04ZGA7CHEs6r1KyHun/+pAKCmPzijDPmfyn0DHaCB3Q/zNr
SXXxt2YnYrWOtslZGujx0JWc0JQh2plHtJ0+K7FJPEPFgPmb4voa5LoT8fq+m4dL8EukjJA9tu2E
0SbVIPz/uP7sWj/fxxeYmFQOsUjDBV9Sj5rKhSdJL1d1JtTv75n/KtmwWAk/DiuM2LixCxS4PojV
X56P6qly3ao4c/z8XhA742YmU0U4QEe55V4ZLAC7ITRWv3+2JSm9eGF0hH50LRMOByf4G0Z0fS3v
TzHv49x2KV6Nez6dIgZx/wZDLtZTLtVIgGs6W00iB8O6UwyqeITekEQ/zloP9vVqDTN9lBdcusdH
mihaT1zrf6ReyFZKzqcRdQ3S/X1bYU5SbmTExKvGIIURQ8OY5ahyDU2rRbkCbdo/kiHljqEjWfH9
4/nTUimZTjuUEsE6oHoUHAt3YgnqNgDJYF6JRfYuvjNdgY54wKAL/BwrteDy9ahrhKfEsa7CDETK
rV5/Eb8g62zRwS5342F4HI0nzvt5gv1hF0dvlfpm12C8pqnMRIVJ8GbMi5Z222PeMcZVIxiiPOZ0
peCHfQnc/DRWBHEjtaORrVD7q3TvrjZ+PLdbkP+IuNQf1xVgg3W0IozN15xjRJ0W70TGi5jShhYs
00iVchre7m0HG5D0uk1d5cjwEIHAB0uXp2RKhe3fwqvO0F2PKmzLwtnT4TSJycTPo3JBHKChZA+P
4tMp7MUHBw8TIcoLH0n1iFIkh5qtxU4/QyN9Q9gGF35Uyy6jfiKWnQGUjmvGMTAWgDTy84rdR/WI
MpBDqcd6awbAh1GUKlbFZtaXs/d2iX0YaQ5ShNTOxSwkKT0GrB3D9JtVea/oyZFvo20nfEI3plUW
osC7A/x3vli9paUlNeR91nNy9G7QPkfMGET2LPDa2azcxWMe1ZcoUnbecunAUJLKSHUQEjqghLji
ySiCKu52cB+BXr9wi7rw9YC/ItXERuZgbhhmnhbKV7jFKQcEQQxmyFqJSPiN4+AJj1xyulnGtiz4
HsbYGJ1eSl86UjOsQop1uijaiOGE5g57m+8K8oxEYoh0LDO9lYal0IoOkAGcx1HyJ4u2rLI3wupb
haXS1vRrOx1GURXlpUIn9bUziMlfaxRQCDCK1qjZI4bZ5W2wN8Fefp1Mp+i4K2ZnYjgQntskXYWM
nvlR+y7V5Y1BZSDnvNvx5QjL6y7CpUUUSCz0urstWNgsOn9SnaxgOK9cAealq5u3XsN5ogHwTJ+P
kpLHJ3CTqq3zKVEudtlKWvpsBmduZi8JtHZLHHAtP75WlgkxTs9FNcZ4lwss9kAxFHBCAvBomUYS
zKy6XkH8z8hpXfHV6V3mm1HQey+LS3l2lvzIV/pasj8+XXHLZ8UDMomELM1cFw9UOpcpxakwR8Se
N6vlzVilVjLrLAZjlU8Du2INSoIi7tQs8J6yexc99futhlioseBIBw0B2G+CDV9wJpNG090mVFxW
pU8jSnAO37fv5Ag7VQ5Np0Thf/KSLpcrs2UO8ovAjHOBd8nExklubbk75El3G+xXeb48YJSFu3mM
odCZJTcC61gkzw30KjyCzbinO2CWuoNx9rWR8jSQgGoJFvgkQ+FpPXoeQa9TX2xaV+EAS34aJ16Z
wgEIkRKPk4lFYf7AHSGzLpKdT4ThqoSdNfGDqZ9vfikIi/49ThiGrVx650ImK/swuSBltSbhvtNQ
5CFWJxNOEnWinnQouG7N1MqkUWkzvR5MfBoMHDzplelcrx2iZ8hxxJaNtDMbEPUPEMcG62d/5c8g
8uy3pO8SoszsImalkEqWh1+8QthxRBT3YELh32PF64LCqHHd/12dJ2o0rD/FVfXoml43/Ml4RJWV
Ha77gmJ9Jw3zEVR8ZLyJ9bVgvxmaFE84wkY6HMzarl571J1y1gwfI9J2Fio/QUP8He+bWTX4pdnp
3j8X1I0nBX4zTCyuUpbm+jwXZY9B3ALg10U6O/8RlDcYqAb3JxQdYqPaaMUfCf35TSkuVhaGwl9W
fcvw96HxxrrF+M2AcJ+NynkovSn/WF+1j/gVjyLobR2mN7zYBrX1ZELIHJpEWCd/zi7nESUTncsD
WC71ke0mtMpCH9/1hjNYuz5tMsdnhKMnKXxWK20hguedinLFBmDEfNFctlGUrjPqb8XjcHvLrUuh
zHwJm8x0415Z0bJw5jmrzfBmCJxSxCMhRXgQ4LGzancSLaKZNcrLR/MnomZ6rsnp4bYdkjVCS5of
YgLBR37AQEsEmejVj733xGWBcL7I8rcP/DkVLnydnXku6C7qwYSb/+JJXWBL49zuQ28+nLarieKv
50fcBVfXgLwv2hqIBPRVfUaFCn16uWea0YMUeqGkdHCJACtIt4tgsK49RMCHAVgeZg4O5Cn4zrVa
Ot9u2XFeGGIfzJkLJ1Nwi2r+hLsB8QPD8ryb0a/ITsvsFn9oCjuZhhrrxBXyOMhfwZqKLfIH5Wtm
kW/KO42ItG/zlc4VvkbZsokACNe5dw0nR8mUj94FFAXgz9YFz6mG+wHX22kY4ZTHGkRd7NqIs52k
5fG2ZaiK6nJct3Onv6CqorOsKjrgV5QtbbBNwuENq7+1PRy9eERw28N7/zh2u8N6Duap1GkA7Bkt
w+ITg5h3/TFYF05c9uoga35c4510ak3bHJhGxK298UQT0J/BcB1cLSUhpHBqTcoT8iohOmjdRs9V
iTqoLS3NhBkw4eLBY48fUnKsQFpj89ZePJAcpkqRNtB4bq+WbeN+SmX797o+AScQho7/nDPyqBXr
eE1zDDTXTMpu5H8RW8Z40fOw9d+Q7txhgJyPEScIpasP/QJTYKL3pMlfRQDeiT1l5IPvCnMO9Ukt
pHhR1o6IwNJKOIpNI1aiHjMzf1Ey7Ps7awk457BfE21BQT3VTLl/IODDIj73A2KfpYqxtvneJAF1
YOGYAzQsGs6mBO3J43V+VzSHic9BEeyf+bP5S7gJdNogeHQXo8apDaHE/V9JUULwBbPqjengPsLe
7nsGN44kheiqed4jWqM0jQ/iKb+LjMrIkw0sKy4VgNUQmSbB/4JquRl8qiO7eTszuHr4w41hZxG/
TjwXk2manIiwqbaiq5ysIChUuSAR5VsF5EW7kSpURHoKukyT5kpjI+Dh1AhCwsAYJY9Zu5/h1cVU
QyFkS/gl5DA8t5tP67Esr9rXv/BBCv2BQYs8t2m5GQxdQPIQMpchHOKzploXPZkbopReGRQQPluH
ERAjY2+syLqMUR6UUP5kYsQsfW6t0wNEnzVbLV2kRVFyIOh08nXw+pTgUFmQM3FdY8Qm0tMMKGrc
xNFIy3vnDuTzB7pO8qL8ctH8X4EijGISjpvpLQExdl/x3oNYTBMtzvsynm9jblovrMqXJ1PvPgnd
XAYPuSu8Ddqssiz1CWJAAeNXZEdWjBoGMx9kBqc4QeZamYSdmLxWhHku6s67EhAuFnCCladpZWCH
8LJ3oOEb/tkOGG7OUBkuAdwBiK5bAaJyZKpe5WFVTA1ocbF4qT6KQvFv1y7PSUxBIrM7lFaGmmoR
u1nreKqyc79ptMsclqbHwQbESPSdDyUgfAm7qy4MFv+GlhMT5yaA2BVeQc7fCZBXDJ+qzgh1+nOP
bsEkE3djygqlz0GOvc8aQAn55NGss7JwcF2/wkHtzetfjf6l2Iy0DQdtCmFxT5rNIe/sTXDHbuZI
uhbva+n9mZ8j/bZSqHRzppVA1KoiEJ1WtVfvjslxENE08ayt4y3JEJtG+JRdIEhmMJG54ZeFe9aM
KQB0CD0BJycHsghdjuRTaY9F+oXDNcKEj8jjr4qZ0QPEKnmm81ZekNc5+Xi9VUJm07wO9KU3nClk
8N0cMTnoNsIyXPonLeJRw12wSARBPLxwFInxizXKKyP4dm2jRo+ZBU7ZPNTa0KsQN0zYT29dFXQi
9lxkt6D+6dtfVTraD5UQTLKAEz8Chixe29VJdvGhE+EApjKUeFhkfURsXseY5wW/IGpRVW3HHwrj
xmkgoU8lE7EecP8hNsIuPE9RAc5jEmGypExILRdhK6wrks3w5mkoMlK+8lkwWYMAM2Z8Dtcirnwg
T3ypeB/SQcErMk2KVoWYDgEszqRta7FXBFf7onlb3XXSa7BVfmgoZqiJqPgdUwIcJ4vdbmQQThLi
8v6y99p2wROztjNVgqmwCp+bg1EbHEOGkr7UiO7a0UV3dZlwO+eHEA8JBKb9IJ7IiqcjdA2kFq5W
0Em9Ttv2r2A8OM414se+YhFzsf1p/KHxf5hgTVj19eIBywED6Q01LuK8aPD31MG5LGZyPRvmhTRn
4Z3HUAgkCiofMZKAnyOwd5Cku/8vIZlVY3bkE+pmxQEyQRatl6UrrWbOajl5bTwOy80bRqjLL2OD
+VFkNXTl5Id51YZ856+Ts4XSmOMsuY0tsolLbsRRPBWg10P7ujwxFKFy1PAs9MYBXYeyGqe50jLD
LBcIcbDvGQv1lTw4lKQTC2kVHJPhPi0fK28Ndbc3DmzhKPQlDNDRL3EeIXj7e1MjT7NfZIz26nZ8
8vjax1iezR/AVSuTSlRi6uHtHQXRMT4bGX7k+oGD6YM2OhuiHjHB4Gt/SyMNoXKW3cmxR1bDorhW
colpAaw5jVjzbGzQIgy3mb1cDQ7ips5h1nyQySPJoaIHYT/VYU8oEHUErsxjRzqA0x1HYfyYCgyq
NMAYwoUf97lDdroVCYDG+QHSFU7XyPCWADMeYyStfzFORMsLxw76kAtnGjjJXHX42rU5Ab9v9B/z
RIxB+lgwyvYcL63JAQGckpF5KqW8QteG7jD2iTD9yDeFol3NgZCpbv316houaX8Exea6n/o9UTQ0
u7nL1KQtKuTZjQ4M0G9I9F3NeWQXIfddOn4ORrTDy+Q7YAqqRTZyucv99onZuBF1Kum/UJmgQauK
d85zbnAZCTjipjCLMfn5f9OXMpHTVVLUyBpyl3BvPckeC+XOuBP7lYioGjfOP9hvxXtyK99Fg4JF
fxKDMD5pG+rFb8vKkQSFKOktvtQbVzP2OLr/J0Q6KDIyx1R+dTpqRZMiXzYWGz1ZNafvK2Xs8THQ
+N91ukA4knxeMVMSL5ZwUaRLP18oWD5MDtqy4E/x52yZQ6vgil722HuYlHEh2Ho9mXdNxNVxYnsl
StHVoQWkjuBe/EFHHp4gr/wxMKsKbQE2eVR+gzCb3ZzIsxFcKSmiIdOuiDT55qYUhDN+8Th+rBqp
0jYyCLt0whroZmb8pFAj7gp7omZ5dnASjhM5quTD3ykNFkaAeo2kWRF1Q+drBVk6lSoW9nTh7u+k
NXMLXqO89qfdTXaPYC1L7rM8qd98UnD4diZzNToU/J0oRVu0PzwJIKZ+d+wJa320D87wrIWiYmYp
cEngdG+LAo+U6jlMgYfm6Vj6qmBr2wqK3RpVTfl2h4T65rVPpK2+RYqXM1Nnq6E1wBzNp4wpU5A0
Xyks+XAjN6FqgQE318GoL8cAzMizvxoCKjqwRBB0dRfHWd1wely83VFZjr+ZO71U3UM42zZ08Smg
hQp1a8G/KYP1mldmh4x1mgOPLwW9puQ8MUttb5+IHoEIcb47ysfAN0G1rFv8pVT7ZVM8iwDNY9XL
PBvAMQ26ncwrJhOTW3+lEqgUxMifUx1Tg8nxS9FBcQ6ddcCCIToQOFEaXAnJDP3qeqrNm8sHFAfL
KiQOTiwBaXHnYnJWj5akW2TEscgtuDYpB/zm5AsEl1kfHpjDWDOWz+3fuWs4UtG+tuIqtBBDM9Wp
JERW7vAGm6IZdWWfAQmToy5jQNYMayagR3oUBU9WOT62MM1JzM3+CEeGriv3dyVIhDM9KICSavJH
SvaPMlqhO8OamN1P/cGyjnyuTYamjTB9gi9QACluAnCi3Lt9PfzhGC5OPO2W8KxjXongqR2VRzi+
dWlMAenRq8JAicD39YBQax9Mj1kS117Q7rNJLDgyhDXYIoQ06/nG0UU3wN/Vv8D+cwgJjO6TOP1q
DzhdFeGbz0h0hfPR82DqzGcRyRKXQ6YxqeZnRQlKPEPfaFJU0ncyFQoedzpKNE7nNmtFDagNUxpb
/5+63X67qTPsCwWgn4iF3NVvAHCoBSJhVQqZKDiCVnch8pkn13cwp4AnYkWxUXzzX4gl2dq8zl99
kbC4MlW/i4CyjeDcatEDuy8Gn19RDcGDrzK3ttHYwxoZqRAcCL4xwlk0/ljyERbbzJAvVoaWCQM0
6pRDgpUa/DuMkfIsiNw2vONTIBzpgiOv+SykVbzGRwCF0kLU4NyR/sKWPdkNrfkSfdPQ4SqmAJ1Q
qdBNhvMUwMXFFc/zFo9I4Ca11yt58Srjaaw7FE+0FEsX9nF2P38k9+d/0utkqoqaxfCbpvw+W7CD
xTZdLNM+ZHUo/cFDL+eH5NjEBohFbrkL8m8gF4BGif/NIbug3W/hW1qhizKN6IsC2TPmYj3SjwZ1
npOoIZBhoLiSmEaXyW48nZsBH5RLf1PM9zhSPY84dn8r8OPd/vlJp5uhi7OL9ucR5w9oP4APS2Mq
Rw6X2mbm6O6g1ZLo67wNUoF7UmgxYMbCYxzxmnDw8JK62v2ROuWXZdriYiLW8eM1/yycH6Zm4cYx
e0U7zmK69R541++Adc8NBl2Xr30S8qH4gv4EWYQsS9cOaDiJSED+JFpfLEJVXAG077DeNBU3Mqip
RsBW5Ry7e35dhj656xQLkz1iYjUHRmD7xwOmBjlBJUwAKnWRPwFb48kRB9TFpA+nAutGWccwd7BI
gDXwEHn5llaqqJcB06xIgOPHtJqHNBDAxXFqHVb5olJACdnwcTNIQAAiAHhXeQlUjZTyFpnuyYO6
gZi/Oa9lw946CYKNu+UunVb5ruIzIO9Cyoht4SIs8g+fIyRwNLGgFTz52+Mf90P8j4rjhC8vdh9L
thPS5Yz9BOrHUxvt4fRVac4wA6vIAsGRHpVUX9Bch+oS61BnGbW+MiPk66q/Xpn2Vz+9SbfqHEoF
aDIcAjyNM/cM+y5xjvSmdSl3/pHUl/986fEkTTEJlHHuex9EVNQFNv8qr0TgHmOxdm8My4Ww9l9h
SsPmj0imUuAyiF6/pC6n2ubHwGA2nMN5aW2PaJtH/kxji89sawmczfnJ+QGYVUrsAqDevwGb8YwK
XD2z9KFovG0d3HrbFARP3UP8XWTubhP8AT3bl2X0BdkyaAl3ZKP6YoNblI/oEPelPMrFr/M8znbJ
hdJE/CoQ1u5r93+DZcvOBZjhXdLfnGgrURW5sGGrABSHuweliO8XfBF5SyMYvyTzvbe5n4N5MqR5
u4yY5i3qse4WgkqW/MGZD8WcYrhP1ZflsMQxg+YlXK72iBIHyt7YrdkX4bL1AMKGWG4e/hQnhqiB
tOy32Bz+n+dOZsc6M/xLGEC3QqtyLBFZwCVdCk7cLmW04AgnUGILNPVtJZ7ie9S+DOcxItbOrHQV
WWx39GmJOuu3uDS7zC9zMFtwmwkQBDUm58eAta6m9Pg/ScVumlBdJ05iXyq2SuJ4kY5ukzzRrZx2
DlsO37lQQXNSDQ4ajhRK7QDuQ6Bfk//I7wBCMTnL1jzW2yOBjm7TSeLj5NWx8q9JwmAdqd2Sjafu
2FRZkc2wrCrV5nWtD1Ov3rSMOXHgsBhH4PHMHs4+wS7kV+cT8QKmkzArPiFjff0eUVPp2ucP83al
ZkvSIxHHPenC4CLfgUo944nbVUttMpvJLYqZD9ucr/SZ5GGGEPxViWa2KxZyl0lGpVcXm7nUoWGn
kCKqI1gxqG11f8ULuDJL5LEsYiAUcB5BYg8je4TKhnrqDa7bAMnU9Lyu5wGXniEeetaVEZh/Hw8q
ckuF9H/6NpOC+l9GBPIlCJPcLqoE5hLd9ffaePps41o+BbmcoJbc9rJ4RcOr0Jfw87VAcRgBOvIW
yNjMcZSUxG/XuwCyAXl4r3YTF6Bet7E27+HqU3XYnhThQnRq0SKE3bgZT37Bb/oMvRyHPQIvr8JZ
MZiM1TpCipTQUwe5iwRGXlQY+uVf4LUfVs715AxJ2L9Ygi90IoZoxOY+Y5lbwOQtQshXGJ99cwDH
lOnIlpCp4gKqkQZaRBWlZUNVjypIq92GAp5eV+R5I1uOL+IAzIa/94vOvrcOgBvGAMb28rHtZMP5
DXCqaIL6vuANIXOoEBa4xpmWBW3Dust2AMNBNWA3LMyuxl4IqsMRBodQWYGh2jyQwma7zCds2nMC
AEAJO4OleKwOJShqXdz2gNWrc5FqXEMbLw4P7I8obj/+BDquVGXD7PyEZVMf0M7YJOHLsHe06xgx
YHdz/lx/+P13OkLDzFBsfsaH2tSNXaDgpxlB0lo5b0WMh+HK+ekEr85ATZtyfVu44+WQe3z/t0Da
MIedHD6h9ztawgA6cyIyukf9PplJYz5Qt00x5V5zXeEsrSV608gluvu+AbHeNpsFeTtR8REMlBqX
RmrxhcC3+AU7NoN3IUPpzKpuHPdMoGmxw9pD4Odn3RpEEnlC0xUGXy+GbMyI72+EyY6ed7niTk9h
kitHBu/hRc9up/a1MOx8+0PvgSUuligoAjr30GBRi80XgelDfgjYSSDVbH2JZooKlsKFOK1ojw4o
o0+geR9xu+Juq/tK0sZaY84ZeE7GHVLfmYLaQAFYJxBYIiEX3y9jIoZmGjVyBVgkAM1DCXLQ5JT6
CRdRpsWXtlXnkuVHLc80SY7gcKEHL2FffKcgm5Ag5fso3OiCIdMbuMWzK7F2IoWbjH8ta3g9cEFM
CYRFfLOo4lXxJpMobSuH8qaapTIFPg9tFXbdcqkhnHTburoBPwSf4JlmXG1p2Ev/Nkwc3LuIFVm8
zHXdXN27Z2DqsjY54LibJMxEctuo8WKSWPXC/PEXoVR2ssmdNUyIs77z/MqRp2J2u8e70ysc/YlM
GBdFIk7nsVpRDYqmYcX0r/H1NuaiOkYEzhhsmZICZ/ITWdiUCJDPtEYW0y/AGUjOGfqynl2vCyrb
Ui9B6Y1YHHf0850aolWOgBkg1FCu6A4er606xEj6Xn0ayELgHzM0syJELlNy2NG9qPopU+YNvwVF
ponmLZgai5Ci5kmpU96ESy/NHXJasuuKPTFBrMwZG6zv8rS1HWlrR56iU5/A9+bZ1MfHDobdFUvX
MeZsvHDQ6Z7+NXkOpe1I9ttpg3IDl4naYoM3D0AKoAubhskPN1/iuEyxBFUrtwbQMUesib6BJ0er
WGGEjiu37DY5QIcHCzSHEdfihpaMgSYxKtmOR5r44m4hqChemYV9UlEurx2ZC78sIawzWe+Gfqb4
/3HXrGXNQRcqsMXD8szmLKx6AtrqTCz4oFoS/pPF497WmtzYadWL8ehHPCN+xGNa937OZ2ZEysQd
7n+0oTe25tGq1LAw6sOHeMzZ26GPKIgSsDb4iHYODbLXAAh7JFNMB1t0BpmpKTlnHJbzvfpn/tR5
JTwMsPkxWyhwH5l25gNBBFMsG6sZfBlGivYQj2k7UycemR7AjiFhVeXk3c49AA9LUpfyQa07OaYm
0yozCCcyKamHqwrvPoRYVZn4FD8ownpp00GW+mjKKdHNs5E0OdvgeEsq8jJD6vMco/nuVZAGcmBQ
IeZD9MXZhMlGmRFdS2NcE7AVTg0BH0hN44EGH2dG48uhGP+CHClM8m+NPEH6EtaCHASw7v3oXCl7
795oECLhekLx3ckQzpP8gqpGhrws5jD9LJvXjyb07C7sU1p1AZaDfbxzer2EZPj7X+7PxWn8QsbB
9I3jQJiyj3w1khFehymtqnuYrSYdf7lTPZFEXrnwr4ZetMlkYXgv1njnQOloGvZHyWKwfVIWjHCd
pqqW5+FCdFiTbyTJN//8YKE7eXXeVmvs7EoodSHwVGQvS/9Ds+rIH2HR5bJNjSgmcW1Xt8Y6tWhb
jb/AvLAmCLoG09fZmhJBc4T/yoZ4j+PK5+7ZjYiOpZ7P+VGCshLjisi9TBlfNeQo3CSzisfIN37n
qhYgIk4ZdneKZ/ilYuYoLn09VuVyCMhXc9Bh/wwarHpLOU5fMNvpCxWNNI0m/uFt5pFiF83kL4bW
MOHGrtoiS0VqbCpGqLTop+LVf6wmULopqMbAPeCNiQmdBWubG6GjhZZAXP9/vZf1cTYgKyhgb2fR
rpPII6/qgePIXqg3U3X6dLTQHyONLd6XiuMPcPzYuQB03DvmrfyizdJnCNoSCHB226VZQ/uoHoQd
3AM9yrJ2QXU62PJOH0WqQkLs2A7Il898bre4PpdF8s8/ERHbkmTdMUuCEA5y8rg6g7msqqhs87Pq
RXjL6jtWrCZ50H1T1HpQd0Y0Vd9BATe5qf8bwmNDQMExmLz3ioukZT0zZx61cVHSS40KIKH81p8Y
G9ZNgddyQMoXWQQLyTXqmGpqjeVeXCkDtkFrCEMUSIxnrlUcuPz2k7Aux48+iUYZWBBUXo8g11Yl
rHe2Uhfx5tGiLXA0q0sQRALt/gXSTLOsE9IA0yxugnJbR6tdgt/PymRoOn+diOEDMbGktO4RLWHV
JujCpI4zfDxcSyZGDufUC7SLkRUByNMl56vJZqCGF7E9qzv7GccJstROYfM0Sx1TZwbndeU0Tdkc
P1RKIHLII42aRNOCxh9ClImIBIKR112cHxxe4HFc3gO9+noSEfb+Wg7ftB91UMAntbHtVOaU9jTK
5j90d1VxAIeZ3MFpSM/xwzwpaqInB3odkcjRCSozFVvxyJkqqU7Ma3qdUWfa9GukC0ZlENrl7jvW
vSbEoECDUyX4qHUTQUSeV2FW7O+lVnCOEvZ9XpQeOCSogCDTtYJmlCLdZBmu5J61A1qYMDGSBSWF
X+sMfeJ+AtIUkkkPUP4SiRLQzvA3D+90zTH5uAKHxL12clu5mcqNkMXvGyEuF3q8zgFkTv4yCiMM
gSkDC883l3FDFMF74E6k/1NszneTiWyL6vx16OPKKlM3Ii5yDR5SLwpRlB+qpZA3I4AmBTyarnpO
+UB1r/5ZqDMQlnXBMAgL25BE3DjOaryDlnAX59oklM0xGeMVpHVpvgmol/q9BGt4xIu5wJ8prNrO
R41fbUt7y5MJKzCFZ5HKHX3c/fafyXiAifb9SHkar5ZSBMeOhR2frDS4VsCXuAGveVmZaWyZGRSf
hehXGcnQ6B+5Pr2r99DU9acE+ORo3jp0R6UQpUCGeWOmqKHsvNPKiXZpl7BgV5e7AWLjBdSPB1VT
hfMnyp9AaU/KPekMiteLIdVDqWL0mHRnUM7wWQDR+I5F8UkVM4Kxxj4jwVZeygz58VoTyBycioDg
3Dr3PssgLHsHYazi9xL+viAoHa4sCnA8H4HN6L2y3BDVRc1tN72nqM/CFD5k/ONsZEEQ5u87VChg
wXl09X3e990a4q6FisJAEIu3p24Lh+VLohT8I4hDMM578auqzv4vYxxWmdtbAqfmAoXlmBIgGB2i
RIsEhHh2ft6L0DtjpGtRjord4F8L056fTMesJ6TfolinYAgpFsRgf016Z5+gL8EsbhAD0HjVBGu0
LZSLfKPe0nTy4j6GNHG17VDeWzUgLx5t5YVqwBeJlFJvHP0QZ6doS4n8QGPuUt0E7r3QsXYBqyCu
sekexW5MTBrLtX8k6fOMY86gLe3Tv83SWv1C+76RG9GlVSIXMfgMJRNqDplglFywfhb28Asvmv8q
DxWM6OTPztV/1h6DiCSpLZgr7M8t3N6Ko0q9ZpjqqXKp7q0K2Nj2Ae9SzPKBtrs2ZnX0WRzunTGe
FBHwh4biHf11U+rxoGIBTAxZDI1CQolf17s/lf39g8VFuVikKf0msnyHzWWPrOf9U4soYtVGeJ6U
nKwCauAh0fDDPMTMf04b+DpKbq1feUawSUrPMzu7ndBbE2eifV98++AvNoNUXYYma5p9GvX889+Q
8jZ5YTAMhYJ+lP+uV99OG2C55I0lnkuYObBQKFmbkWLE5OUmUEkEtMWTJy/rCh/cZv9ixVmJCtap
hvl+qbwQ4E75LYX8ft8jyy98qUbM5iePz93T+kDW8TdEXkHljbdfctrgPsGzfwQUFgsVwjvlqKFO
5IsEFqicsJmMPTNYo1Tw5VhpJ7cWTvJRS/6ai+cn81jyv97xqwNXvUq0Yc/QP4zq+i10rrwr/V9J
i1RLHiA7PnX2Lv1elGcoJHpTK4jRZ2G9rq1d9QD67sXu+JMk4ayJCFAonGDvShI4y4OQlXRgjX+m
2xl7QYZe9sdraB7P09lJ+oYnD1Ld5kP22RNq6ecaRSIRpsId2KH1FunrSeKp1iH8QYN0k0Yyym1h
bSx/1tIGuNkq6uweHW9DptUh9ZuZjgKWnE/BMyn0zcTUo3F0U5wt20QDsO5Pu8TzZZJr4noloK+V
5U7iM7rip8/fvUmz40Pq6WrLoh0rf5HplfVlIeDuVIWlnnl6jG2uSCRy/G1xp24ZbmhUQKt2DcWn
uNpkwoRcf2RVLlwDKxLmYPtB+m4OXK2718FSatcczq8ZN5eJ+mmNuMQhqN0Fe/iXqGyJmkjMgmq7
TZTcuP6fGVonUruD0Xl9SaCw6vtnKdkhVJ7SsOat4EnCmIb46Sz+/AqstVhgz0MB5Af7Fzk8kFNA
fMwpd2I9+f6sc/N78gnemCfpJt4RBhAxkBQjdaqENytW0LSbOJsjJOaWf3y0lD24l1KeIBXzfORq
2IuiQ4gSn+bdn47gHW0dHw6BXaJ+ee2JJxy2HprP58KGYrPvcPLv91PK9mW9IhCYE5GvADQ+6GQx
m7PdpO7SBcCSVm0SFJ1kCA5GfQLikAMljWzVUs683mbrRs0OlchAybiQ7WhQogKdBeYOk69/nqwL
sUtqRAz9o/hTAdao83JoyYNuyNxeA12q0y6TAgnFmsi9HNxnrHQX6hvU+jF0Vf86BuP4EGa41iti
vBNkyZ87D0NasBGzh+oti/AQCrTK/X0ckl6S/P+7BhTjNRaS0av3O8metht1jYji3EI6gnreVkL5
p+fgushpFhvsdAcAk89e9w8UDF1xC/XQX8ikTvca2Vjy2Z/7KT9cY8BI9Pt65U2WVRiA0if6tWwC
jqtHFlhPkGyNmNrroMp97flJBUJpTKoL2PWLvKGt6Gxu2/cT8iCc55zu77qE8PC8vxHj5pozKuxq
JtjxLDbBw5SobHBWct5zs3a/KY2H1X50WOy1qIP6rqDrI9St+u42Xk6cXo4wLGpiMQqtPoRxfAYz
FI03UumU84U9A5VCM3jRyAjj+IoYbWoTyXnHh/fs+msGPoRaGcqqHlW6V/4Wxc+JxpHUPtDzmAW4
/5ruhElO92Ehp9XlgdKW6jvszTe66iLC2dHsFokfJsi0rF8rEyf97wvtz/NsMD+lXHGlcxq72pm2
MJno2KrnaqbFbxfOLxaAynpZle1PA+25XYvhxUcXEbqpXMOIdpqmKCcMr4JsrgNu/LPT981a3rUE
G1/ix/1fBfIdZg8AZXvv9gRLgdO0ISfBlgaOPKb4pRNTWY/9OJrrpAnmHmelQAwqoa9KwlPNvFc8
azqCrwyR1qX3ARzmdzN3WpC+ueSYLezbmH6eZWf6KcRFjzmHDnSA0t5nNNe8Mi+zOb4ZkXWrbR2A
MIqAOHsMk7c/ODqy92lcdGSbX7B+suvI2yVsA0Rf66FcFAi189v0Caeg75272fzDyA4i6kM2RtD5
Yry22qxq4fbTac6ZiolCA7v7jlASNWGC9d6CE0LkCLIrBxdyxH8XWudGMufUwgCk+YBc19Ewa/nr
v5+tHzDut2ED0ksE3Pcxcx1FSVNhqdGuoNjpAoCdcvl1lq5Ru6ctje/h1SAhN+lqbEr1gNkyGEL/
c3bDsb59hcrOs9nnUn1faCgAIVOQNzd2BAxQTOaTxhWFQjU3Wq3nlwrKYvcVq6RLJIa8bXqriu01
yu3JGI++muwXnILc3Yiv0r94jsF9HGGPOQnw/sjqp2eJkShfB4y+j24LlYx1rkBdKXmukcxG2dQR
e1zu/DNp+SAgCTC0fM2RsnjfwqItrq7sX9egigqqtUP0nDH2GuE7mEq1l7sJ83+HUWOiIOVf6iYI
Evbl7VRuZLWTmwTtf87gssuLilw4GisXDsGpYeZVMvpSIuxC4k67tN9BpJ7KsYIB2677fN2zn6R5
+5O9//9InYPru1/sIyM4VDxBuXL6GoyBJsQYyvQDO4TLiYFZCt1J948mmPD3xWPAYHfgb13nX1kq
bXCboWwezD79hINMDXAaa5kvutJJJiHWcxFJvSV2Kz4XY+aH3ludUSmzQH6JLcM+CuH8Xsmcg87D
2Ykm83C2x0Kzou0GEbHAlYNE8ZueLvnMeHEJFgcTdXjljZEXJrSTJvckUqJVW8MKg20mstzKvY/K
FP3eB5CzPs6d2z3Nc5NVw/1log68c99FHoEgAVYC9uN9DttndpC8K+/A1wSBRgPhhkHh0ihF1fv2
xKLGGf7iiA95Nx5JWg82qN1SOf4W5uRh/HbnJVmluxrahGWHRqh/mHMAhYVRMD+7O8GgKPmlJPRt
ozgGWOzF4nrjzW7QkPL7lTIMvapLTtOLprjxI1YTtEFV0ZQ/F/hiGFYj7LklikEF49bOpv+7ce2Z
4496J6nNQsdRMQuPYM0evKvG69dFy8zJz1tCkQzcJfw0wwmJYCxGSPad6Or6CP8IHyJbySCMlVlE
E73XpBRNlHGYU1f9O0slwXjG/xz8neCZwUuI1GYcG/cXh5VKubEmfiQIbKsGMKFzfto38Sr4Qdb+
Iwof/4tIW6wLZh8BN7d6ZLaXORHVV5VSRfRNzjE6ifpHIShE1ExAgpCbCxSMwTehfgYFvat/ndp6
x6gikeZlzOk5h6wkxS2l8/kj5cQBCgasHiEO5hO509B/qgBbRE+A2FRCtP9c3KjGTF5WIwqmhSg5
x15pmtKhquSm+kxE3RVyj3kjKpZpzSy/2r2QyKdGcbLt5XLx+Q5me3NNl1M4hT0rwclKNYYdhsyT
9NOGOQHtIUhhzYFUjps42TLsoVQXppQIW80Zd9+tIJ6SrSmtx8xVIyNNlk6meycpzGdDQQ0xnaMe
b6aWJXE6BcYbArzi+AYdUHVFkTQpUBHJO1XZB+U2+padMV/dhsaiLmCvLkvSx5eVZC836HBGVUcM
ACKpkwf4+9vQcqjWRACAqSGCTWx0yIofXNiLmjG6ZIqcTzJrzgti8Fv88a/Gvd/iUu9pSrlWpCtb
+0Rvrsz+A7nHt5Mztz9iNFNtNm4U2DXBZh+qdw7JcPSdlnkhuwv2Kd6y0VgXZtw4G5NZC6jTpblU
jGaAsnDZj0oKKBYmjY6BB/LiVJMN2j6nCyCeGTjZksshdciWX7xnMtPSnzsmbTS5WZ7xjPBmk1j4
XufRkjRYLj4FReExSKTL8SY4eBOeWHsHvDwC0ROu7dMDinnWLKyS7bFPt0Ft+Xx1db9OXfJILAJ9
Yn+CHj777Ljp6YE/wClZ/XqMjj/mVq+3JLfrlXr11YEKMXKOcLRkH99ceT71v1gwgbLkOYfBjL4E
wRvUTh8bPZQF2nXDTaCjkrfIex81iQ5LDGkmBIHbd92I17WbKKR71ytATxOHib+m1OETlQJO3ROO
8knkX8QDtw/mXKXnwQ40Ikong0/RW/0Pj3n9I4Oqx5R6FACbKtI3jYL4qeB2NnSdlfsJtfLyB1sr
/35D+ZXi2fJD3dPSPwuGQ0Fp2JWJDNdCq/Hida71vJ1inWt3RAA/LpJrPGNhUzoC4X8Cp77t/it/
Nl54xkQREgBxZq9s2t8BEqsorBRcHpvjb9q2Xt7s/O3f5aQ3shRMCho2Ax0pqhdo1IgpKZwAL8Gd
UQP9TV9VdkPN50UmOWLnveasN6W/OeFrgxmcJlMQpFwuqUJ+FOUXxkvNhMez0hrn/n8j6Ikqqe5P
1jg3x0PTynzZbbK6uVMk5CJ89pE8AcqGT3ZpIqXDfy/WGojfusvwTw8k+xlhggrDiqDl1SlNRyZE
ehnxTRa2yXlQSY9fyBj/rRNutZcvvFBponYiTODo8dNpmIPQTgM8E/4I16iJjWfq522JERjTf5+8
kiQ0x7tvDjVpWQnCgIJ7BjyhVGxSoVEgNKQVBgkk9RQ3n2X7GdGK8CVGCv6nQoLcvI8tgjyLZU5E
k5ddjkx2yNRZUD6hl9wgJ/xGfwxJtftMc1hMPFFiSkmb3p5TXfdYX1S5D/2/8msbHDCZ0ZAE8zK9
3NTCXTkiW15WuaKVciG3YUPxH4dJiXFsdufgJHgkihoRsoTjCsQFrIocDDLN3CCkUXVhzpRbsbKF
1EiOIE8CTYCf8cU/RSuqPQtyILMRnkDrTI/vmuoSbdr0A5of/XsG+Fwa2KWZHfgnkn/Mg3ko7Qiy
KnlSYyKqTvDKq0zBy9QxEOGFH4xuwaWtI91ED3gxbzlGQ5ospKwRD0Iq1sY47JQhNWUerlPEnDAM
5u9Tnb2VHmOz9pMAdLJsZ2tZh5e5k4PwC/AUdST1eJ/b2CvjWnvR3WmWVZl5/Snq/xYIxvi++qDM
35kbs29jTVTeQxPi+KdzeGDRhItI5OiHThfijntT8aeytafvQNNYgbbmIPhvoPSGVPCmhUkbL6UE
5scakSDUReNZYyVK9CwnwHIRSLF0gVK/T8nQPj2d77E72zV2jMQq0AaLqVgH2Yyak4MGyuuJ3fUz
WQ0/3GvpAv2ktys8K4eP8DBJH1MNQTHZXPWerb1Vtd0rnpJIiVeHJiDoG60Y1PQMkW/K0GsKu4Ao
Ih07LfMpVWMR9z5Uxtgbzb6i1NvNhhArVY5tY8RbeY0FOQfgORfcJH+u7TFhy4fiA2d8WI5iJJh6
mtn+tswNM6eHKRhUAK+bELsW3PQpuPSBp5f3MDwthsu72AsjzlyO+jlgQ46N0Z0Xygm1PZOcMmrJ
BwfHf+RKf/HX7htxA5/rJ9j0BoSgNMenIB06HmiwFNsXn1rAPukowLOIpt3MsqeD4qvwDytRg0qe
0JchVt9EPfibrQhv7S609JgypSR0AfQ5KDJqqH01A+cDLiodS0w/bMg8WYFxwc60Yu0DOz7dvh5y
pAwONKbtIh9DvCe69bKXAnT8J8BDhnuXkf42zNs8wPCkVmAKCXVHnJuBaR/GeAgiNkOPNN2AL/z+
GtCE+5Xp01JmuIePDbJU2ClO/Lz7kgSBs3nZZw7jYsF1gUI6efAyFsTjgSe3sfwvDibB3WOrg6Aq
aEpztWv7USHXP5MRH2VD6QYqeuqYFJOfX1QXNxAopO+2aB3uvp1G6JzeeEd+6aBGcNp00LxOUTCO
egVJg5jKjNOVi0uxwp4/b9v4mYawawzLlV1R7RZlcZvRv9ufvpKQhlYyE84AbSMj2WYUpchTIAQo
I38krWiJ4B6ua+J4aB/GyxfZaJZKNz2BQBHiNz9zW50kK+E2epXm3blmp9OVlV8esdpHNOc+F+wD
DrFrlHkiY8O2g/yCm1JWkpKDmIRnW2vqWAt48MLXWIsUHZrPDEJTFYBFiKsQuXkdiVICvVT9IWOc
JDfvTjKCqQGsIaUpmQ+plDA9TO6nXhMT6Smq2F3CuxS0KVQBPYyo49/6FqJEI+l3/prCYcMVT+q2
fhWI07XCwjepeq2FDOBqdMCK97TcX+Q5YcdD08q91vUgRldqreS6m6ZfuNapk6un4EJtHwvZDO6y
kdqNhpk5mkZLpWBlKUA33FjJU2K0sGcwJIeUmzvut7dyrDKEXYF5fUWTpx8u0G04uSOUPhHeG8kk
ucqDCTaaD/8IQ+wV6TXpQFlSzG1mr7XRx7DStmR14ZIGJHKJtp6GN+9XTf4EG/EHUSvZdw8056aY
ql+9uBlr81DEetUCju/3RFyzJB8KFE09VLCAvxDwUOHRZxesQNtez3X/Zt/WEaadyCPetr0e66Vx
gnPUmn/osepCpjE54yruoyaATfFGD/OzQqxZytP4AIblJcSXhcybMCvk2rxemsOJfqoOOdEWFJLQ
EUQoHiiE7AAconMdcokyhVzUBPHMpi9Q0hJ30flgf0ghPHwajhuMn7f7GSrqLC62iHoqHbWw++8w
2WO1EWa9TsOzfdWjz97k40cJnhYgfRU7KbGdgixQIZ1NbBlmX/yE7itzyIma+mTGfNiWaME9wncY
zBZtiPFfVlbbPLSTObJJwfXq4Z44cQ3oHsQDkGGhhZiGZbeZBbpurOgpk34BA+50JeLT+PSusFIO
2ga5rlup72vO3SC4vbffOcdPo91L+EUu73kABaVn2ohByDuPkmEhQvcFpkr8lUxXIgyt/lsT89vj
BasSIeIFIkcoxcM4McrdOqytGPewm4Eghfny9ynD4kHt2dt9kKzMFdur6BBJOZpPUEJ1vVr5uNlJ
8ZofSgk7OUN9h0iAJJMxDOxX1XHX42N0m6aOncMFyN0/dgTzrIAmtjMNHmCQv2r5flR77UNDd5TI
5YWsvffJA/NVCawmla24vK6SIQdwxYSMDlpzXLF7Fpn7XKA1qo/GzczWAuT5lMEeHKm7sqmbXW80
BPLrXuWtTROX3g5V0Ijo8xjfOiiB5xoWLClfVJTgajC4WYwZGzXQ4vLs2x3UO2XmOG8hb3SfUyA5
V+pPLgN/5hUIrvP4qs9L8lIAp26f3yznE+oZyVUalBDaTOjJPvRAu22f3BE3sKGyfAtpeLfcusWx
adaYl3gwqpHFGMKJEM6PNvtvcJtEKTaEjpEbgXDBM7bAkjKcclQBS0A7TIA8pFbYw35a3ROs4SNq
jeeNCMrgelQ2GoduGvHprb7kGdn4ZroY76L3R47drY7i5dme8CPLCbIJ/9yw1mGBiQ6D1kWQYnCG
cIsD/X7IqQ1pKMgGEZXMhDacT4fFiP39ls4jnt7cNOsMnTd4JxamllfyKLeHjsu2zviHa6H7t1JI
5NuWnOfVNUF4BXc06uNAidAs48x3leUUFc82veiOHXGeostO2jmVOJwv68UEfrDUps1P++Wc/Wju
kdIGAtRNB11HZwh04yf/P41kUVnKvYQIhskZdihsyul/4uNy6hEg1J4fmpwQE2IDLbz6dYMlkw8K
PgCfX8uNDdaLdgGnD6Goi+cD9W3pa7rEuozs0rVV+zHdDQveBL9osJiGD+7ctKkBLVaiLeHyJ+Jp
HkL9RLdxc3WIBnjohzF1J0lGahTP8RQsnvygAAqwfO9P9OYvwU7/yu5iOMbjfcmMaYFAq01yfHCA
l8zQ6JmzH4sXyB6WYRJJOmsoo3fdGFslztmjCbUwGJn1baZkJUuBQ8d5MT7AxflmdZ/5QzCLz8sa
cTSQTQYv9ZOPr8k4Oz/LV1nKeBoT97e/v5ILMkzf+JZo3KSlfAyKXJxENvLaOO/RcnoVK3qdJVjL
MMuFDhKO/X/z2znI6Cs94JhYy4gM1rIKQjZ41d6T+zCqz66JUzbLtNQssZllLwCmzbDnZTQZpN+f
UaR1tylXUoo7f+N3nDXGhGLAOR0gcQ40r5GafOtRoIuQ6j8MrNcqZQUayKuw+FIO4OQQ/1qDX4I3
xV9aMgQs4+HNzEX+SVMc79DyLuK30j/lpb2fQFzIMSgo4vAJJsewjNvTVXm8eOy+TFMaViVbMHnW
TO1A867m9XKTZr2vgMGaC28ue77QqwKt9bBQ9QVB4Gab94HmNQoZCF+O/UtzkxW2xzXD7++o6z7s
VsCVThITWFnCO3p3Pg6TkS/7mEbWH5NSJf7+9m5fRx/bvdenm2s0D1zilajpACjGXudI1zzwodSD
yLlSkJQxTQ6CePBXK0NcZDUhzRrEVcV/216bbX5D3pgeTRXulCpvIptyWS2PB0mKJMRRhZDiqlcM
ZTmBxxd/Ss8mW6yoqyVOKvpeI7PSc2uKuBYO6jZ5jgB7ezWSD9NUJgKpcHuoIG3FsMkpqjDcW0ZP
tpggJ/uAC3NFx5IuQKH66ZOc0jd0kO06BU1UUmBSg9I3re5226bBHUxq+9zewh08sDpvFur4Vviy
9hX8n8VIIZhLcAk2x4QtJbnAxkFHL8oqIigBzfVLbGHdrd/UTxcMjpP5pMaN/4XnNWENegAxSkli
T6pC9T6q+nk8Ihho4hbsEwYX5Rp4AX31Kyuc4Nb7mw4D5Gpj7RjNZcV9jFPXOG4G/I4G+3OL3liN
wJjOckGz8IMAUiySaV8CrLvEBAkVwiZ9ENhKp/dX5OvOpdcb5Mq6H4XhpcfUupGOsNtz5DIDrt79
S6oTMZs866JAic4wqBy39U05zoOFNGUmP0uPRMiGuDM7Pk74zjben1oCmlfE/nrUqaqxvp5LPfw2
KNKO8SdSStSvW1LXHFgaBEEHNYuzQot/nm938dQmT7ge7JAjBI/DL5PK8OXfgP2wrCHioD8jf791
dnHIekGsSVzUvgTW70nPBNFtZjo3ho1+H+pPyAzqNDNfhGBEeqrZVONgIT2u5D+efQtp/JxNAJxh
HbIlc4fIluehWECLDdNHm9nafP5gvLQ2U1l9vyrFrHbrDvLIYGZxXt3ZXLWkNl4aDjO/6/VNQKP3
j1/X2biKno3HmUyHvt2Q68e+foZ5MAhPwd57rIAafW82p9v46vuq9Pg3aN570t4t/l724HQbk3dI
oV+cRkSb2tGxHvGbuURXIU4d+LnQI709fumVzUX+ppVQrjDVf5HWuKIvDpZ3m/UQO2EPIyTbYPaY
64RBSDzvto8Git1Th/nqNyyC7sR7el+qZbEUf8PZyzR8uuXuzQe/ZdvRX3zPDGH1iyuucc3qACEf
x7rDE20vvCDBw1zSexOK3F4Gv/WW2RSX8jlm0kbj+1u4s6Qp2yTx+8hVD2FGVXtmeVYjcvdhLTBm
vEEOD3cQKeNqa/MhDPbzRVcIlnhnp56umn0c9k3Gdc/4+BFYkIpQ25vmAx1jsqVCpRJUge36WckI
PO3YYPv/fkLwdEhxK7R68jTiCu+9BdeK+teJQJaQhDeey42MGCMzE6vOSE9ch5vK1J7mp/UsrZ46
diAffDlOzZac+ap4tKLpBDrsYham1Ul46HjbUcVfTFPXHbOG19xjuHVYepDjivSdiVjcGItMY3kQ
/b25laqWxsAyvenpH0mkOv/pEt1tJatVKa9xd4XNlHNJ/PxKCi/Ao7wQ0mH1FxgL+fHDDc88KLA4
A+SJMTzSXBeHRhGSurJGnTDOQrJRzpT+kW3V14NP/AkK+LUlEUvFkTpFiIgDkiMIHYqBBcxrXNgY
IGzZpkKbKGOF2v9JdaXTCQYTQUcXTQF9KvxXgMq0hEyutntmJavhOuY/Cu92tspC+kmogm5hKho9
0OcRYxLMKSil67Ngpq1sf3K9vQkFxbjG4v77E94PXboH4W5xVytYzPuNFDUEnV+L9Ko+JkZ1Ek8A
qAnnaqBZmdevEvFZnCNrggnRSqYUX65Gc3cORP9GR29cvtCB02eWgGqfeIIPy3HIqSr1EXzrCXDS
WrgViho9VMYYistOz/HfnayjctyGjwzhkkS8mJP1qWtsR2rfDAPI82Ka27fiYJr4zItN0wQmrn7t
yLU+VgCldT+K7OigoilIn/KvCVrlnG0JN73bYCsNG6mvHPB9mCq4TMuGc+0oVXTwK/SdyZ+A20Jn
MxKsG7V3Q01cKEjgK8I0781w0DuxFtiqAYJ8r+CwkOhSWaJxMr6qLURYgyPN4qBRIgKRny1WHpYv
hVksOPmbvEQBZwnEMdUnyA/RylD+6RhOCL4AzAoZR/kofyrN03J7d4xM+UfsPfqzuaJK8fg257Nf
YLOA/Ytz+Isck3L4UN6gzEM/JgecuinC2+nBKb6+FhK2QyaF061wqf3tFx8opqPmqkbjTBepSWMe
f2tZYHUGMy8xxpWsVrEVOrExZmf3OSgZ7YO+ZvWg6mpqO2rfbZgNyKjP8b9V5o7cS1j0OAETIAXa
WzPfdFOSb/sGYCs1BEdyvoumLlCe+gQ5rAbWFe1UtjYPm9Dba7JrPp6lJkbMGGkokJUI2gJ4UWSu
AHK7lTMyLsVGnTdjo6mHH8PBj4pl3A8h88ZELB2q4HPInWWqb6HjN3yW+gbbJdo1OJFb4KbN8rhd
hL9IxWZEz0yy2yFdGXKcQLTU7TwyyfVe8nx48a0dTPuGfWzfeESc0jUE+m0UNqZX6XsbWNI0huAJ
E2qMq11BVmuUUk5E0cywxT5f26+yW/Djyl41L+WW0LX4NiunbgEdkwwNpujQfy9AVQhT9qbWX1/9
DTDUUy0qKJ5nyKEqtF6HjjEVA9S692drAxLDcncyPlaqKoi24K4lDUs1+eR3NgjGJnzF7g0m9Er7
IJQLRnKjx1nB5TrHhHeuhUHTTzDcudmbuhKq0pu5781FrmlFblPzX1eqAJWrL1GKnfEbzTl2OZZk
1rt4JvLVVtw+DbztvPOou84Hsrg+oBqvEZoy66aS5WXFwuGXUtyBZCkYOIwTLLDla5UhK0l9SdNM
vLCxLwJu1LLvacDX/RJnrvYaioT7yFYavH+HJvDmcjrMHVX1nPzeTkuTaeCNUbXkXfmHboRFbp2x
EcfA/HtpNYs2QRdkFRloPaLVZCm1bC6w/42JbcahNQSkIIqrkv2f1c6Kk18dVmx7mCW8S2WVlA5/
eeqePLb49UH0yR7ilu6UG+A4bP7gk/PHslgJsE6bG7ou2/TtNbr1o9h013cvCC2jqfVEIm1jlQbd
vwXTBTYJ7f1bw7pFg7+9mAYDgZOmyZ4KqAL14VSrhniRlXzb9tXrogzcNmmpE6BSdh0ReKGZsB71
HcU5RFR7P5jPzust8EwBXgz78j8HUVweX2NNO1gpBw6K0bEvgIQMbrAQsiBapFKqShfdGKnGM5yd
UQuxGQOmIgOsmrTMATczxyCkOY6JUsaYf6snoPqHSv8xlijMsr+Uo0lv0HzUTcxxmAIIZqT1rrX2
+I+AX4y3cDRdyR0Utp/SRQUGD/B32C7RKeoSNX1ApVye2VmRJVeqBZPYhGno4oPTt2971vfDQ3Dj
bfr3TkN+UwjU8Siht5rwMBHj8o0VL4ttzO+0FG5jHtaArKtAR58bFoHQjFBn0Ie32NUdEKZGJTgj
d2m6BsFmIoyC7Jbf9duIRAUqLvCPCjNd1mkvhfAYawKr8Gk0UuiKEPpqLIyg1YdokF0v/tZHUr6r
iZZJnFOfopoI3xpzS17bolK0IyMpnDTpuqIHAC+FkECu0s/e49ZY7SDQTRDqzGcFmeFh6kFYNDR0
4J1fGvGc6WfbvrDlLzxF2VLL2kR+McWdrusAvBVjTM8HYiHLRBknEa0XS2OBJIpQDG2M38bST9vT
/hY2Q6il0yBVoF0HpLBqcjQxxh8CjfWoxWVvXhYcbRMd4m+nYVaJu6e5hORw2UnAqhuQEzbOaNO5
8Ra/ahBadXgVf1gZr595PyX3FZ/9fqMQOuOmvyBK+G5aSLMi9jg1HIoZ+g/unFTfLuPcmIU9yY6p
gkEpdhRKd1DhJgQt+YlWELRo2g3nNddo8VCGmXRBxvLoSHSphsvPbwqUrS1TZpKWmBTdSJMKerVL
pjV8FX6F8PFSrOR+nSlRGo04/u/ygrlfZ1urb7KuROSK4M0EYhqv6N5i55SWOzaraXBKJynWCeHy
42cgt1Oxra386rB5lGE3mpFHttd+CP9FwAgSr21/I5qqWnImh706HQmp+XYk+/kSwykpJ2VUF0PG
gdd/fz7O6BZfoPcyBSTXs4yx+dGZPiWG2/I6pdsJqkZnyP3MWdUL+lzmN5mV4hSZ1ali0XjmYna7
6G3pqD0paIR25lyUJFcFocon7ppScYMxke/LZa1jxVpBru5F2C8CF4+kJ3TOu0+HXlUdpzwg8KHc
7K4Pb8ceRiRYyRVR2S6wj5Nd0NA22S/oW4/eR6JyhLmLTYbL8rBKNnormttQ7d7w9mZA5SkgftD7
3WDwTlsQKFKWuAxNYkpYAthdL6HjmpjfUagbcU486aEJlZoLWYTyoanPuYCZ3T5s+Mjdcg2ae9Ut
Vtf0PauDjeo30kcrmxB6oCEIbfnLVBFaDMijMGnoypCekHFO5ZoN3lR4QANTJZEE1sRQm38P23LK
GAqAAclztqFvpnYlHg9RCbEL/MLiyOaYHMB37qOVP5drKW2JnZPFn1uhsxkz+VKo+Zf8Tvh3Y28B
pB2BKGQt58NmN94ihpAlCdkRxqCxS/tUsaMgkcoO1+Ch0/uASBiI39Q4zO46CcenunSuSecf03OE
jOHCTbb+0o5X6JsY5qdkbqK1yYSkVpJP9qgMiJ425K/cwbmzYHVvo+N0y8WQRyKQyIcmVCeIYOO0
2PaUV2hKPyiI6WTdJi3SQQcNQbyck/AoufJ7a9t/pb1Kxr/Z/7zEFD7xiyxOjcMBkaKDjZxp7sgH
/kXkiNneV7gg7M6xZ/npSA1TsS3zdaCWaBT8abJZlssrTimja4zXY6tyL6DIw6ChdFOBuqEtWg4L
GA6p+aCEO4F8PtzwGCsn+KzgUgQQsX28+/OJS75Lb/J3+G7afB8HYLtlfpUh+pR+iUy/Ek+lM8V6
3MQ4GI+MLAMFPXI/9Zc/FYZ1XxyAK9GdpzvzOcrSgRSG/62iXHJEM6sw5uV2JD7lAmgfmEGw6jpA
dg2s7ip3ZW0sZHiAOlfhhmy5nvrIoIFB377UM02TbWhIuV5NvhNgG2TzlrWAM5P9Grg+5+WaVWIQ
ZI59KF93FdhI5S/fOHIKKJEblyHRpUy/tsqVNuvfefghLCOy6rHc5+i+Zfk8hoX21Fa387YR8HBD
uV8KO4iz05+D31U0d832ngmvvx61EoakIXuPP6rNGw0EG8NQVrNyMo2GF1YTQtLXVCfQe4wsAU5n
PLQ3NVpZ26PmFKdqWQu5z0gFNWtK6Qcc+xyuITPfSdN4R1FW3dFXnXvjhuDoMfY+44eJTKbDAEJz
QeKysxqXazjEQ5pn/dlTaXC4kOts1PI7D/7+SaaPteMzGTqBPlBZTzKWAUvBhEFeVuWdx7sV22mY
Ifk6YQwgvYdKjt/8X/AQQ111D61Zg9NjRBRp6VMDjif5KPPuefGJp26/hk7nzVJgQBS+J/ITDjni
THEdse0RV3f2DYMJ4oodK6G0G0QxDAnp6rRTDylVWi9HHsVzq4+BY92fWW2i/xB0Lcr+vDCt9qxX
rRXNRj1ot8AnwSYnJSPagCo3gK06LsVSm7dvRILLze0uJZzmIM8w9MHCibLFiKw2lERepTbVzl2V
rjDK2nx570VGg3CVGEP+WlHvv2pKxqmaoWbIHcT5KXuqZr2YDQXZw05yrd5Bf5zwCHafze29CzH2
K3h4i1x+Uq2iP5cyx+S0rPQuob4Dev9p6lZlRTsf0hECnzHN1JS5pgHl3JaS6uP5DzoyRmql/Ziw
Mz48vcpVc8FUyFvvhN4qk0KNntGdp9rCXlnDd3jkmfPQBQsMwAHpG1/N4192b+bWuUYWHrkiRNp3
RttHmJ23d0zvqevNokO8Bn01yNU5e5mUl9amd6g2vCd19gpncEpl5l3nCH4NT4wBE+JYEBUalTsk
Rb5fVbcutiCk/fCHMr8erOgcH4N+KlHlgYN3JItNaaFBzJofVxS+l/wJq/2n+P5wuHL9CFjLgOfz
d7wWFv/NdMltTEPZLiJFjo4XX2G5mNQXCCbbYcOyew2sPpuaiHuYCkRS7OZTgo73tVcyJht/tFjx
H+FGHdWv+1jA1UuMZOL+Zdn/iNknt5hAFWUmN33mB2zJIhPcjUQQ2oFKquU8ULLrCf5kfedKR8qL
FQ8D+jNdCeEupUCSIWiSsmwUmS2YEoXymhlkh1IcELehL7qPI2zXc4wG177FpHkliY4GbnARllHF
zTCQ+WmfGrcTgUoZqYF6BkrJNKb43QqmmMUrnDsC7/QdTlmooAtuyWNa99Hpphur96yybQZGGk/Y
dv77CP1bA4wDzsSXPX829CNNZ0idkXZuYEc2U53/2qw3FM7RjMTIHS7Bhh9OuX8FQaCQ7gBB5N4+
SfQrlvg55M4zj/VU84sZmA3QDgDjzEbdhHy6DT7eTfajffIFoEm2BH7H1TF0+XcXFGjx+q9X+bq8
N43fdYE6GzBS1s1Lx8XCf22EXM15xrS+ig/fx2hHDnMcQctrwaWaf3cGDcMofiVj6EN2xcV7eeMf
BKeHfiFvW+cwaTCVoKGXfqW14oUo/LhVQpZALgq8wsZuVPKBgRpVZITMktqDptkCQ7VeChZO8+Qe
7LtZiAWd8S2vy0UfaP6KWMXrtrlE6g+Adck82cwP9JuUxZreuzsRFpA5dEhhEuQWBac/9PQ9NrlF
Snk+wEZ+HHlVnOL21bRc3PTXMH8gB+59wdq3DsDVm0xL196SK+uo54Eh1t4zKMo82dWFvpR+twRD
+93bgDDV0y/hE7WRUxfpQ1mviu4tTyjGpG3+f3XswSV/43p4H3hN0EG/bLcNK4SxeZCU0jeMAfCv
hwpWAZxfXs7Ba1cue383wZra2GGi5vG1ztZwUv83ZtuulPjJpWT91xUjGuZOP2CSOULqFBNZDwv6
QMqn58vxXn6K5KUctcSYEIp4SoDUGZgL1UFaRrgW7QGHp/cmk1zinaYxQL7smaG8l/533nKlYZco
gpSOAlR+9H1fGNHyIgANL11nYKkSvfecaJecQA4pLnxNZtSkIrsWFyQYl93XFpvbEoNIE/WV1561
/s1Ob9Di65CGn4ickFR28rMUzpyYVrrM/aPo5KtVRWmXdlR8O5PDMQTX9SWZIhze2/S1wsdDHmT2
7+C+8LmdrjGQVe50EAdk0DMvm5de7njgzo8Xq2/dMCJVzPVjcBi6IfjAYSzC2cs0RJ9i/WJgFT5c
Swv7H4xP1CrlNErmW5oSo9m3RSidcihx4yEErEaDLTmyhZt81FIHuvlGLP61QVqMZrJ+eF8jH+3N
YUghD+dRK0/Qdlk9G9VHAf2pmGtza8OkV+JnefMf5EDjdEQwfTGxdTEWCOwlpz5swgYIHey63dvL
vJg3W5Lf+q0zn2YSPNl6wlR0Hzfc11j2xm1CIagLnIzk2O81KVr8H7fC27glqc9UYFdRl6Ay4190
u2uLgH5YTcAdKHCkHgigSZnM5ayRTD5/NVEtOb8G8pDwVCIdWmVb6Dj23tOuS2pJpJdNSXJnxhbr
+hbN9qjxHNO4rPf+rp+Lan3YELXsxJt2DC5dHWA9grsdSeqE0/4LPVNrmwn9awPwRxSwuTY0RNA3
mGXrgLqt+OV45m7/kV+93ZhgRVJ4Oa2mm+Mxdyu8n+1DWeLbn1uEcnhqJ9ZazjQhoiqtYmUoQHhT
PKqgq4pdMjp6M+3tuvoBBJlra4jQSEIXFQn9vxYuC4wsKuKdIS9/154fIiQ0VLtVxfTbrJd56mXf
abMoMoW1x+h7k4+YY0tL9Yu8qa6j7zYExGmnCFhFegnV7qtEJZhmJzaDPSQ8qSB7GVsl9K926ah2
jtlSA4sw/57EPqdOj0XAl3Ky6mFIIi3VKM2Jk/inpZKwZzggpjO09lKNuUrMADLTAa+YEbYpKSaj
udTrhiAd1pAHMA+Rrg65aoGTFH3Au1tlk3vngUU/uPx5dqK+4Hzl6iyQXlBqGRMNFzmJNjwrNhVO
8QGpWtkRecQnV27r1AgYd708uoqugUmaCfmtYetcoKcHbBBLSfgdNcnm9ubKbVra7n+99/+tm4OQ
0Z3CCj7cX800Eji71WpxMsMn6yD4m0Gb0LEm72/6NIltoPt7/OJz0T0XRiLSCo03ASHTdiLepihI
Iuh1NZQdJI3WkbUjXlq0YahRivMwlW4jUllpIJ4y9keOEyOaaLyFaskH0+iMLyWRat9KxTPzAY9c
kXLtPPIUWALl6Th1kCflKQ4VYxTFp+akbXWR/pxXPq5F8QLGYImrGOI/rao7jXnVREdmqexpUrUf
2bF68zRuGdbtOPr0O67CSLiG+mGgHNuHSxajMN4Zp3wRcNIVWScZ0dTxFfeQxUXV5lfQxRdizIw8
VdYoP54AXxTK65hBZ2M/EZtASE6AzM8VfGs83AI/9R4pfivmaR0eOlbax90oG7JDTh9rr6G6Jxoz
dOGHIOVXoKk/LdEzugOmg7LfAgR4SJOfLNk0geSiug9FLp6mY9JaFAtncesjo1fpO0KPlNp5bASm
CC3XZxKo2Mm4t2tlzxfd1QOzQAVmzcvDA+qGzR/2Gq/E9nscUcawUVrILVsy5XVsQFipIdMcV/e0
+lO8Nlgwhdpj7F+KK2+BFAaSv69pns0AWF2PNn7Oyv2CR1X+Q5zqmlD0O+mwBYxO16cJ/j6Ql9Ui
cnpQwNBDJQEM14VJO/NGdrpenNXBMNcuSWrbFnTGsnRnZGHhXSBx5cBtpfLO982fqtsK6SsliCen
1ZgwNNbc7PRXYq/Ulu0lvbAxtRGqAHheBIMTI00UOMxj79mGBVGfVTfYxEFsjMZYjJFusqaKgTTz
c1hETX1+U97iUk7INRIGRiqqKf4OVxxXtYevWuf9diCbc0DmrBzfQRjS7gac2HEmNfn/3G06kkby
wYn4xoBJZejRrmLnF1tQ8o+ZHW8fpykQHGowUc6tv5FN/iEUDRBywgEGOIIlrf4N5iHcwkZbFfSg
3/AXQN8VAgxyWTMXA/Jfp/1L1CzE2kESL7k1mwTytUZ4IzGbF/4vMYyzNMnClD17h4Jk/ydrLCrl
kWoSSERBrzReNO47Dzrljt7f2iawNBalKmH/8pBYsOEdAEQ8nm+CgQjQ+4zPlZHW6e9zRulGS2uA
4sdEsrmeYJOFSVuWNv0VJDQJXLw6SpI40twrA0GmuiPzyZRbS7uYNW4LVbyjc4xvPd+bBK1K9rvI
NS2gqgek9q/Uunw0vDaJiEtleVwdbWlferDIfhNpZD4hOUXe7nNFxFymCGZG14HNHLvICqdBsnwp
S9flz0Tzej4oZJFNoSV6fhARSKOlHT12rJRrpNNHhgjkuqPD9Bc3b8EU5jDY4ULL8gYAEMj7stj9
fxb1/F520lIObyXsrkV5bswuO4uksqH1RG1l19BkYPPty0Vu/BtX8D/UEMUd+H18FDbofxVIz4VE
/ykWdNJNLjJ1uoRKWEMPKRgbQOnsEwpU6mn+f7vVk56DMpiFaYt3kz5/Om0wWEr3utzpuTBvptLy
viBlTUCPVGFuM0AYmSLlNDLaW/hwfiNcnCLYDn3gWRPTLPJOAKYaAQI7+yF5i0lHRPHpWKXny6VC
5RfQ5nACIcoVXIdJOPdkt4kkaut372IegYq3Zvx/r4n1kNfEMpgLoAtRxLQ14mIegdSHflRmV2Hr
D1tq9j3qvVoew2HmV3oakLacioPFdLu66o9EzGQlQ3eiqKTCDxfZeI4c3/4EOYakfm2fok7A+uTS
VoqQku6VRbAZK3VjCi27AIsiPUlMMGJuRxQPEQU+XuNWOjWfdUJUvKG0XnhfW7u9nv+mhQ+2Z3IH
HnyS/e4N63TXXf52iTLAP2+tyxM9U8OHZwZqNIyLwo1sWWQlUyki74aoZi22A94ieNAO9kP1AtXt
+zWqvmGFxmN8ZxFpppVf+Ve8R6S8ugAkib3pqW4SD2mTz/e3Y7jwCOicl0M5EH51SBOPrQUVBdf+
kcfPals1hFN/tZMr62erigr9mTbwIbg0Umufmp1h+c1mvvA0WLr3mcHNHJm+XEn1Br/TVbFheFzH
Lz32skLLCNgR0iLw8cTZ77ZfCsLGA/LPMjREm7l0uFQj9GMPZ0DSLxZgYW5lJIzbyDvSKeNmFKmt
MjH7mSCCldMuamRLX/FmGatj9Ymaeld9t5hsQGJR+JefY50oSj/hRn9JmjMMCIj4OnnoyTWqWC+i
i2AljHrx1T/zO6y2JheuyQJraTkECntuTk1D/0QD+CU/3oAzOz33OeGhuJ7mQ99NBjvjN654Lv4/
dp9LUIwWe1RAVjLNVuahVXJvx28+iwYu7iYiWp5pamqwCKDM00KvwBq3mHyaHLORajMBADuU1DNv
5VmWCDznsUirozLJkEuFQscbkdCpF343WMdda+1rjkgPK7RDoWWXt7OHOKPMdRpx1Oz7XsBVF6HQ
EEjAVBG10hIoMJS/q2HaKPhfVv7cZrdbT2xiS4cZUC5NBoHNcxWKSus+numtrrtZ1j3NsdFQhQqp
Jg/I1EB8vXnUgRFF+7CFiY5W0C2blh4juqGMKkhITBptA4trjGLqccNNmHTgdyvoO6rQdoB+ypxt
LoajBykDbnsRG1MbOGjEuFHEGLg+ZLnlMp93ZM5uVgNTJyJ4N9xN3GKa8jNinFSqRHH/jGDwrPBH
8iyxs94NKgJmkUrNsQmYVNtQRAULDnh095FRTdTeO3lNAY9m76YfFI4XC+UhEZR3mJd0TIG3Yemn
t3cEv4HrV7WkHqz4/emK1jM734R40rHbsr6obUDINmWGc39eJyrScqyd9CK+tJKgG63tdDCQ1jx+
2v24Zfsa1kT4xmtlqoLwzC1mQMONW0r1v7BErJnihXQZ0baZfnNSO5k7/7rgRe6ZvRYz6lVvMkXz
vm5jyKbdcpV7KufQZ+/tWKsoxidySoUguWa56+Pztqz8Qdwo6tH1ZZZO90vkPwyQl9bO0ogoCTXr
9UaBKRIHVh5LA3VFoMrOKtLo1iIKiPJA3ta5rm3s+0bTRGQkPKsQdpuNnPgIiJ52AGKFrDfSahgZ
CadIK4Ylx+7GXfpWpK0YFZ6AZOCcNhy4XFm0+5M5GC8bb30td2E2pnak+rQAO+AyM4yCWtTLViO4
U07FuQcUrvZ05PCrFEliwJsDIypWMF0oYNkm6tCyvJQIX/c9NKdmsor0qpXXrZgbWOw+0mFrUsvM
Pf13qf9MmC/CBUI/33aQ3XeDaCB7GP2+qoZIVIytpEUYJoMM+na24vZD/hWOoAzzIh/giQQAupkF
/iw+hjpsnAyw7gekD3/E9CBHD/ZDCuZgWEa0DI3dzG+eTICjc5WdJ5yFXEQ2gDwkeJb1Rrv/ErRz
jAlMeCrK0O68R0l+51+QjlElQuVIv7IFKFuRWfOyyKqz22WZLY78rDtuG4t3IRYEFyshue5lrTPd
6EC8K1TAnnTRiSqlIu1Tb0lJPeWpAk1ac4EiVP4mN/w7aIS2CmS/sjRYzAr6ERGLe1tN87Qd322K
uehQ+yMrdZpWr2/aip4e56fix5U3XCNhXYTJ2CoaCeVsHx2XXFR80wZAGDytqFMIw4OYeVxVhFHE
btLfyJpHumwZ78qpYFXPyrxgIN/hS8tvtFV8sqec81R1a0BwkiZdynV2uqp3phRXttmzrl0Pe1wF
YRn4S8O4pJ96oibNHkmhFIG7tOV+Q3xDb1zVROEDDGQ1NFC4G/7HNSb4g61rbvpW2lg1AKm+EORX
mXk4yXaj3O90Fhppqt7JLWDDlLq38zR12f5Pp43DfWe3UJ2Lw5WUD0O2GYG8XaP0+UO5QJ7DxUzY
wZWnQgDb7HkvGR6em/i2p0yto6uy9EuWDX5z6a3zelMNjgeuU6590jFcs/RvXjhj1SNaQkRfyV55
eVEA9+QLaZnBIr1caJ6SxJn+P1YasDWKf+CTBBhNDWDQ2j2/8tXxcv2mwAerTt/x0eGG7/9QSyN9
OZP2wvyRQsz9EH6xA3BPQdT11wTz2j0GkFvswqaijX1d3psjrp2GN/s5sPDSWkVjbftgMjpJTJTa
UE06dTuJsecWI/w7uhTVeUpdYQeO9iiX6KZMDoOIE8ukBK26U0s/CkUXjJW6K62KCgcicRB/4ESe
xmG/WJeQhmlbXjcao/8y3PsvThpbC0anFDrsueB+hN/FySAmjjbXDHSOkP8BS937qOi0y8+MYuSy
1CMzo2cOTeeINNRth+qawvI9xpOkfp6Usa7JJaNVQrR5MKoRPqs8rDIzGu3JpheonAzlqMPWuJAI
xP1THMvS/CaA6cOgw128qNDrsRgd9xR1EbdtPr8a5qXwjIFArSkFVoI80QqDvrk0OnIV0r1RMFv0
bh3ksROiO+7P3N1icyIMSAyUa1F0fQee4/sHsATzENFwwdLYFQ1TJ5Ux8+OW51XDdisQhkV+hEIX
8wbnHePPryZM/uSdAHo51/DI54lzAJfKqb96Du1azBYhNVccnzgfZJ60qDAiQUAgg7qqL4PKmOyj
oq/pbchNXh5QdOv4bDiAhswlbIGMyiooQurf22SGfv7PEGpL7DOhjsJvAx/iTqsFJ7mqDKEzK7Mp
AQtAKJ1yJg6/+T+9S6fw2abXr0fEO7yVZMBOmgc+8ZpN+R22AGVSN1566XgKs2T55cFSYBeDgGQJ
xUYMtsNYqThzKi83JJdTolIx6MKFvNfVp4ETYFOp33LXb/OAFXGubaC7Vc1LZ7HbrJ04VjuhlhHp
KG14ooStrevQgiLxh5bbJwfqivWwnWDQbHiQbKyDenxK1MLyL5OZR1c1um0MpKWCqE36S9930qae
EVyv8bWknaF5OkacCumn62SVBRDBnIAOlULxMpRPrrdW4nBO7Qlm8DyGVWoDm6DuLj2TL8enMHQF
lH+CElnMa9veJ8/OJy7/kLLQQJ+8+v1gw/1vwMdFs47uxl+imAht/o9Ons2dU2ZoJVKim+9MOMgn
DPi6bdEvXGokzeLHH2hrh5HN7UnWW3MfnzkW70XuyY4W/zMPD7GCWg2DpXYeP3Sl35rV1gXeg466
9DcQAAPGIsZHDNrlFqVJ8KmTxZtFIIFTAyapJcrLpsZ3neTdyIOFuVctQfu6PwujrkLr/LQiiuK5
xkQtk4vuGN/dySFxg0otrRjON4DWkMftcnoSDigrxtBOBHLQdhS8RZW6suVmB7GZNfYsFtazXNio
RouXfSGMGnztZe9QQBgfmmStIZDGMk+kiEhqgR/GqPYt87pkx4h51EdteDtdcpxBydCUNNeW6TTf
2p4FMds/Wxh8Q2bSpjWMOPwVxRmDB7u5cTHQmjUlDsSEMc8SxMjNrKIacLa7PCAzOJbGod+cnpRN
eWu0fUPf7horkqUPlwuhzByATgSD1ChvATxIz7N03CKnemC2ehQV8Nc9RdsxGmy5OzDKWAhnT5a5
pzT5SlCj3uXIFBYFa9qLdlJmlVYNALikhLNxx1VSmFP1NXeyI5zBDJf459MEH/phI/i9KI1Ob5ER
bh2M4cXZVLBJvXZpSayzBcarilfEfmlWRwzJYHHbDLRqBIY9FKtREvyDyG50cr3YQB3M3+1DF9Cf
V7VmmYbLhZlRq2KWilWG26doeFfyTS0vpuyf1uHsCHnpzOTVfu/h5KkeVyhnV0Sl9FqfQggtkevd
R+EU7TNwtyCF2S7fcWvWdU8n5oSoqHPX8kskpjHlBdtJJzAqVmSLdTjj09nrHK7mVN4KkBjWJazx
FWW7pIcQFUo9nzJIONs2kNnabrHivdDwkTTXzGLTALExy/j3tOvURkBTIfcsJqAH709H1UcECARV
Pd7aA0EUTTnZKjfxr6gPpYyK5wP4AGdYDhRzVFsmnXq+xZnXfDxhuYbSiuS7hM3bOTEQ9NugciH4
qnWiG35L4Tp2lqg9zYlEMZ/Y5uTX0S4tnI6PfgaGvCg4LfN0bYiKoX5CN3x4FYLuW813qmdqudh2
AU/2tmLS8TFzB5P165475kGZoInz7kmSJlGOK2Jtt+sD3xuI3kUKsMmOR/yHHzcwj6J6O0rV8twk
JxoJpzFl9iWW9k7UeGgQ26aR2HCane0RBb8XjdiAvlbvOJVoTtYykw6zpBwqXa1NkW4nTP+gNkNf
L6LNoVULdSmewasDlWqr3Q6OCsnyLGQv1OP2utQeuyvZuGAdlJKUwTuRwpfIeUtTQbqg+bO0p3K1
SDT4VFirNa04GJt7h3smQ1W8afuoj8jd0JP39v/LSBdqzz/6S0lYADnp8IQpBG9FNJl0cp57sWO0
CXyXoHkzuPBdeBCH/ggGygtwNAd4IKs4EEVtM+6h1f6ECr/vcX4hMj82Nj7WaHFickFIA8ldy5EX
uCpY7OPeaBTbh1NIo/UBWm9KcgyNQLD2tFo9WqFX5mgHEEL41c3r1MObxg8yNGeqQmqBqNuwNXXr
Zo7QvEGMIqekOphh1ogbUgBws3/6WzCttWXJtE1qq7ATU02OZhdTCYDiQGa6agiD+79OXvsWC7jn
Xuf3OD2IHjr2WA6iL8MUEdR7rEHGy8/qUG+wLUJbMwhgEiNLagjb/UQq9adn0KoIgHuNekdb2EeX
HrDgFNAQvzZZhoMMkTahE5M6yNmz/KXofVkh7oaMNgUldEozy7y1Qwa9OXWbUHY3u8LPJ4DQeYkA
zjTEsbUCMRErT3O/4TbabCoONDJ7YDabK+fPNhy9jmoomgttcnHL3vNg4RxehJNJjNfbmoFgnand
ZHNVdtJ9peMuF8olXlDKyyHRL4LNCjikUWRVFgkZWri5+t50m+ydaLOqJoudDnqwwpY7OLbdSxn9
9Jh3wY5rNFn/ZgJ0Ln3oHmdpKQgu02Xe+93Y29lJU63S5r9NdPz5ozVvQARF+Xw2GTXcUxsAjzTF
KohMMxYxnzA/CMoT/6KLd73zoF2mkD7+oql6y9lHzjUXRNkiboaJhlCsDfJOeDLeEc2fYmG1Eq2X
l28d2uvMnycZwYl78vIuJqxZ2AVfd10mPe16t5kQi7xNyX54yflx3SA7CFVXyf+aULPoiV/OZbzq
9YBNU0bKqMvBiuyqnATLtzMRaMwr7Dw0SeIwjkrddfc8rSii/POwkQEfaZGT2E29tR3uQj3Ltjvg
c4tUglfkcZDvjpJLmxdy/RVsXDmDY0gZ27Jbzdm8Sx2FkRCN3IuILEneWcYMRTvN4z3TRPSFB/LG
5XqtBmInS5TOkWFQcwxPI7gYgXftcd2XJcsT+kWvF1nEWMrkSeggVw+T2Ohg+Tl+H2fxS09LtX7g
aWJt1CcqZmUjj9vnaix0tEjgWRJObF2U3a24WekfdoySUFxMECp5awPfkL9NDFLn3yjaqcYdti+P
qQPW142NqUrVcd0ms9wPUmjs1g1XM2kG1ukcgSjv0SlFyMbMvx5ksBJ+4eJwF1NJwa8p5tj76UeB
jxL9YsBNSYD9JJ2H/D+MeC5fM/irl0Kvaii907+Udo96+UU2X9umIv1n/BzkqWA0x0d9AXUxxIDh
MkzGM6SE3AhxpbSZzIMgTeDZUfmqozbtFZUmZfA41gO6nocn+KdfVah7fPX53NAWs2mqj22Hl41V
HH3iRynWRJnYkDlVDDx5cjT6tCIHe41QGQeF65bLCOt2jKC4qm4lLTYXks4+gcn3WlAnHOOlfOh9
Bff3MGzxVC4G3q2fJkmhQp8EvPDV9DMgFbP0VfWu+zMIjNOF1eKXSw+jVjbTakzERXO4akbxg8dW
9ZC5l5j7wuzWK4tSlr3ENA1uJD1t+KLMjifL6L2wW3zwgPRQXi6yTipkRBoMXddfqVDJKtUFEbg6
SUwrqSzC3enKYMTlGUaHQEmdvTURF4JLOm3IHZjHEjJBNKUqSWTk2uvuJHthtzXM0hlFMbEEkRbX
MEUgyDpoDqYfVWf8gYmPO6EZUO9o33a/H5MePrylWlt8yrpN1uSxQ79wAF0m1rYF5vkEsOHIl03n
4gTRMg04ZhaKNFGj0fgS+eavC0jE5qrPokCs+zHCVYVEhxXXzRhCHzvcJ1Xa5zl6JTxyBfdPGNW6
h0R6pPTzF7I5XdSaZB7uJujWxuMOzJPGJKMMkwuow4b49cjTgEDE2Trf5oIjQJTetnjmuAhE24eA
0tqn02y3ykGYo8JmU+GlU8mQF8xB5yqsHt95xsgJGfolgUsfqd5/rrn84WCEGZ9W28UyHZsdbTOl
YXf0Qg4NjDutyJSK3JOUhHcv2s6YMZr5TUm9fNGYkPLuUfh6dKUWn2PdGjNsIDdXt9OAggB/ejv5
VdiNbPX6MPUIvD4yHPN5SxwU6G1HV3mVUyox/G7xYYBw1Hrb+k3elZNINhZRtyWIOxQ8nXoVtkWJ
qjjWW6YG9FbDwygK/gW26w+q8su44Fg3J11pDdN7NPU2moAwdMhJ4Gy6RpxRhzYNksdc9pfHFJoV
vIXt11gGuO+/HOSn0fZe07xm1ib6l2tDrAHbpVj/zc0lQVCreTqxBSOEW6emqR1LiOb0gnri4WWU
5azBM4xNtM5q72S0PWPFnMc7SilbHcSvkXU3D8MrGBCKm64tHiXbWeg6wsEK8QWeF7D9YI5zsmE+
FJBCfN8ENL8THb+Tp+WmSwfDWcfrOhj/MOjStDP4VmAmPTl6/UeZDtLMWyS2cijcfvWDsVgGUtwM
LQ0xT8oUjzEZ/4Ueohg9JfyVNqqow19u/51V9i/X0aX0gUlycrIw5W1T04kx2LXZFxXu6hfZ/RlY
2yt/wLa8QwjjwoQh1McS7BxP4Sxpm3Q6wPWUiYpGuqo78IANdWJchPMkkD1Uv25bQPpYWk8Bn4e5
o4he8rPyzqnDm3/T90TizXdM0dSXyfIMNYbLOEbw3bpIr6g/xbVJw9ZZfUSHlMi2pLYdj6GSY0B4
6R4euFddTkXFal19JGLe6hLNmtPD2NIRi4yNp5DecIvEuB6p+MwjX3mSIntT47NbBLqyzxB9iWux
PUC3YvnPVwEH9AXXHEiSzW8PTc3+4cxT8cOIGkbW+iuxxDyVoC3ys9rFBH8HqbC6LDkD1jTOeThe
Gdzf502uV9ywXJ+ub3CNjThqqtromdvc8iROdCicBxYvf0cZQ4HW/2w6Hl0CAUQ7zVP15bi9P15U
QTyLskHVIcdMYCynrpl2MfmHe+vD9P+pLctHiM77hrWa2TGEEEBVoj81f23KUDKMTHbLQKBRT9jw
qxVbxLTXW0/rNtH00pPtNzayPQlPuQryQ/SI9ANPjr9BQ2byQYyTar4GxzdW+l5mxPodhAg0VZmF
YdcJf6Fvp7+ZxfIS5n2DgZp4aEB621/39VBTAjQUwKmpnWTwKy7EhvtIcOpV+yU2RI8MGKz38xcE
V0kl5iLRpJ+yOSQrZecLM5vQxexWK/6VKjGtR3+XXOY5yc05wqPmXGh80eflvAdEipeAEVq+bSuI
Ww6AEPC7t75SjLw5WYJY6RDbYVYuDLDKd8dTdNv7LOJVCCBhnOFRc0b7ObZWEitQhM9JAttunFGV
7OWbQHqktAuO7cTLADO/tYjVqoVzRbjOaGTiMD8ZILTNlLRMN93APFCHEEm8j5Q463OgRWr506z9
d5TFucg1l8RGXuGCOcEY/YNUx4Hsw/UbG4VfRxr88JQuuQPQxRTYj8leRLIdAYa3wOrIpJZxkHoK
g2SxCQTzMJhJHbsp9L7PXaUHp0IqWBa2xr3xojTNseZev8ntBB3KH1wkCh8nWzhbg3+YrO3amq9C
B7PgxiNH05Er7rJzlujkGtQ96oNAxcNen8ACApgayg8lCOR1ivaCDeSWmsHjlU/RcHUUXFhq2aTj
2KSgGd4mATJ69ZGIUVwHkBicJeBJ5sXUOZNajqwK3SaJpYHksxt7JkFomUkPI6lGqQqHWbMDNSqi
aLwUu3QVWtySxfSw53Fp/uO5+tcVwfM1zHyc3sszRPPVqjTA1gYH2eIvBPPazwtf19khcXgOGHC8
OmFwgt5QN0SdVYW9O3CUWsYQg/Cencepy8HDH33z9OpeH3DR4ZqTiL4RpeSQ7bsl2rVR4PZm1Q3T
oA44mQicSH87o+BDVUQmXgkWbDwCmBvvDiB76i8mGGchtpx+Ub05ICDto4iA/Dwol6JrzWYFCsUa
KGIIBBYgFQibGlOqsU1v09omjHesG84Nt8eJ7ouB3H59Y5qxFl+TfGzlBvpZMdZT2Qk+keRYLDDY
wXkcA2ysKUCIcUmU7WReBAf7JhTf53efR2xJELJoGz+NDy57fpmOSZd5OVzq3wXUbnxv8gQ6maBM
qYrGxY1QremqaeKWl6HqX0re548gyYdRqQefiea87Dqy+Jd/LJEW126j+5u3DoqVLst8yb8qQR9n
L156xcn8GhyzdFpzWMuwu4MT6cAZjedeTA51naE64ZuSYdHMSezAUlFLvI1eMe9qcO1lnGL0y4lt
lx58iGLRhVMnVEuQvMN7rRTpFnMCcuK46jZgNoXDTIzzEX1i96HLhIhE9Gw5M4+G0DMmPTOVQaFw
qKcAS8qKSmDlFudZIAGYZdlE/1hxTI3fCcBiA3vN19yp9yqxPeda1+AfHS7+U5NPs139b7CtWjTL
WP7ctbCBMud1xTMRqzs5ItZSv5FtNobVX6gQajYlVZQcFH42bXKv4UFOq7TKK5xMy60LXOPD4ZOI
rinuemJ05BEhLWWbpbrKCUqUK3WCUdLCiCpgCg9P5YdR0vY3Dj83hg38sVOKtVFfbjAaVO7UV2rA
v2lJ5CyzW4ZbJ8B4ZNCsynjUNh7nLgJ6EkVdZe6Pya5CpthKKmgaVUy8gtgdhC198FB9biS1UPMP
nKkhqTa6uRCrYCsoF1gQAHbVwTHURvrZTr423DwlvaXY+xg0AfYtRztThfZtk4lU05/LeFnFNRgA
Efde8okACfDzVLMfdlvm2WCulfS6D5Qhpy9D44tcXZn8cPuXx0DOeAX8IU1wBDgEo/hUYak4oPOQ
tHatmg7w5thcIWWorMveMr3Hw38Lj26xq81VS+VbN5GCOqzJcPFx3LHzlvIYyxfmD1RgyHIRJ1GT
jAiSYh/6lrar1yMqcY9t5SyREAY3EcsSRlncCoDJQi88mR5kPn2NErSGr6DQl6x0MBE9TZfv3eaj
Bb7i1S5JFP/ygj44mBJHBI6mE5opa9Qaj44kr8BxBOSopRvLrx9ht4t3hABaE8pT07Hxh2kuWpSd
0OxbgoBE8O8JdcAZW9hZJ90w9F5kqPD9voE87ws6vGZDBYmC8tQ25U5h1S9WynokVmz9rtFpgbyp
zBDWJbO3RcEi6Mm1DU4p33PiNSzKErCbKziygYKr0q8KWTgtkDtEIO63QRx4uC6SmK6zMfs/c4OQ
W2SbSlK+6Ean/f6yDBLGzggERhUGsKFi79+EEW3xptB1BKM5wLeTcFbIsFKyB6ufLQrJibt5zyWS
NsEuBsO/sfZiA48pK32Ti0mFNHUOL1Ik1AuXYvrWECwZLsLAeTCxcAbyauxyLdLqrRwPt3k4b+q5
dh+BX50gyl6Aw5jRUZ2D+ByvW6yINj9a4GA7AUsUiAz2aKtita0Ss5z3yMSLUXSWXfmAcHpXJSLT
4hQCuyUrovd9eGNFR/JWDUCxBeoWUYTJoTMyh2Dk9e4pAfmDyD6Vs44Y2UhU3ZwhBWYN4RxB1ZvN
xe7eLL/xSt1FtjgAE3rpQBUjyznTtIIiv9L6NhXtdYbL6JavfU6uAgQftmBkXa87MTlRp0oMZul+
Fyp87xNyDvTjEyvgvyPUD5XVzCN/9v+aQlxMWBe/2xQUWoJ+W21eN2COOoI92p3n5zH73IzvGmh4
EmT7RXm2yibNCkEtzQgevNXcLRFWZhAmjYD/xzUv/DTjp4RCF/BJCEb9IX9ZcDs0HIme9rL2VjEZ
H0pHQOnquTaMQrCsZ3baSRblUT+RDUf/bwGxmBqgFnBREwZr8aRzOOl4YawNHGuObAy4TdrbAOrN
+H0bh4ghz7rtSfvPPZabo5CHBTn2lSXnQ+nfW6pNYN57ZUzJj6is6bi7nhyLCa9nEdaZ8CzZgegM
MNLlrGZp9lrjDFUptariGoPgOz53amCkHKKEu3VMN8GYvCSzjFH++QsHxqkAHSxtwTAs+wlE7ZgW
CvgU6iHXxxlftSJ/jsf1upk5qqNASorqV7cg6TVH2cGgmg04Pj7f4SHpORU2SVjhpRRJt2Au9P4W
+OfwYJjBQX8JW5r4Whzybn6v4eQ/MBhIhcTzW2khQVHJ6wxi0EpvTmTFtRjj5GXV35TBKkSy0Cfr
46nLtHK4mHsVYs/R+AAWijOmVflKuGaatWQ8bWinDrYIbniV5+eObwBCkd1LmPINCcv6FuVryi7U
5J9LwJsXPji56pWTgqFzHGChAX2ClThzFzQWxZps+KWpztmie0JSdQsgvlqA+aInsz9SoG93KUfk
LRuaCBRmBLd3s2LJf+B56MIzFs42kzMbIdOX2Bk0f/Yb2dbB6IKZhr0SRjSVKk2+v42ceRgroJ+D
A2vm/2L1APrsCgc/N2E3xtN6IpEHRnv3QPCZj+tRmr+POXVDcbQGtueFQwtuMhLe5EYGCVBCsZfQ
VPgyzrB+/Xl4tTJGZNp5AhKYe6r2l/GAt/nSpd49wx/X7vP+5eXLc95x4wQhHlt6zbEVm1Eohqw4
WPIHvTO86Tr7LAhuaEnRMySSexcgiI2LjP/dF2OuuNFxobsrcxkUrxBT2yK72pVN62GGrUAKvEKe
899T78D22QVoXsFkiIhrXyzH4XU4r/YZ07ExF040/Bh7M5yOARmUSlKns17hxmCQJ0GwrsKzcKvw
MfKq+HJGLhT4hFvJq8gi/0KnNGOb39Gmy7yrFlqyhWushHGxF2Tj7l7UYXmkP+NtDq0BdDtEtjMO
ZYOTVCyRpQV7x2X735W3ongrkfELJUuqjd+MUi5oWgCtjf72tdffCNm4hC4aRNBbotC8rsZ/O6ZC
pKTZYELNrCG6/E0Zo4VZO6+EgJsSM8OIYm/7pPM7G7nv5MChMrsg4DoGNnE3CTZgNIseL1V0Voi5
SrNNnYGMmfsVarDo4pouDdW5gpwahMn0ve3spC7onGeK6Y8a/RJdCXfogPWFEVGSXOr7Ek6TRevC
X0fArCuNa++IrBtTiz1diE/ndIAWXTpYwLAMs9viaqbQ2NT4h3//L7/ioLAAgdDUMUv0kp/eo7gB
KSjgVKnVOmGA67UsulWlxzvXY65IdhsqqyMv1vHvFfoh2Q95MQCVBeONXnyBQOfznrBjAWQWEf8f
wKwwPOod2txz4N1RKbh6kr2GmuurIayVPxJe4NJAC3LscjbtM90mhBy06kzeW7bdUOOq6FY3X110
8lAhc3QrkP0nAYnHNZY1N8UmoD21tIRVWWCUGaG5QBEcKbw5YdnkGNZxBFYqF1bOtMZx5oWb6/U3
qqVI2WVG9aQHRIQ014DrkjgbpBpG9PUPpWeBtTg0D2JKrjOE54y8k+zV97mKsqxtUrrGSMWRkwge
8kE4eAvWLGEbV6b+EesnVC8HASk4dHavGjuHw8sQxgCLkjjtrK4NaIlKv4dgU2d7qLMtRnxCjsTy
mStGk/7WHnUxw18lmrwNq2WQAENj4CZ3qeH5NwLWnFPLIFwdMAm3MUzPF6h6jVC2PWlRzneBsgga
Gpo70nmNyjpo8Xy4WK19T86SdmjV29MTiU9DLB12zoZWlLYeQOMnvBPYVIKsDE+y3lEYEoR1ap1a
26z69MscUPxu6cODEIMolYFBo1htiJL2Bi+wfRNy+MgQB5WyE1UnxikALVLsZP5JeKdXPtHnqr+a
kCLC/uOl1pN0Zpkj9MWAY3Ctmk29/layi2fipYAptnrjv4Q5TsRep0Zh9CBdNk2/D9/RCToT6CGz
WtOxexoLwHn7BkrK+PeeKKlH2+ZSUrNo7uwC0kDa1bTieS0ZQccMSP52T4MpCsuWufzPxSVZKUlA
bnnZYJ8DIAJqHiKZpxbIa3MVgHmnZtdTvAAs5p13ARchNjG/5OJOLB85JmC+TaSs46llVoXBZ/lC
0ZPX/+pE/cQ/wsSE1zPbkYmOdFLucF1cs4fSdALIoXKKzyapPUJYb4VTTa5/zh0MFC4mPqeHFekq
X22Xt2h5HbLfPxfltaaGta7iZ/JZXfQAIWP7QRefFtXSyyHEnRqhZmjW6oPBn/6nVZuFP8QZR/0U
jWi9wHWa9f6mqx2ceR+RSBSTqowvylOY8uE4Z+x6l21CAmAAdLiKea5gEjKLlFcOjwbXXMn1Bfa7
QHzHzmlDWAyXzdlCSo7kRzwa7BbR+vjZifPCPNrLq6DCUyqMX1+SeiduIoyqzm4rU8brEAMXk6eL
AAzCAobAYhvtSu3OW7s1neu9KNQxJ/lxT7/z0FPwjJWSJYVIPlf6P38q6jd8T9k59VE9bTbU/4im
/IxCEy7RXthv2IeHu2bYcO+3lpclkuRntiUcngvo64vJ09uwTmGzKWgr1BbI4KxQMv52VEijEDpG
+unLSS6jIsM5s7Y0NkxB5ujeEMI4nMCV4OxR3e+lMz402dor5KO6edtjV0ysSYB2V7YPp11bBzPA
ctjoB1WkbMlxddZBhGy4oFcw0xkKHj10XtZ2VDdPTYPPcZ/ic3d4fOQ4gh83jxukN7bGM/6Wf85W
EjokXfcNBefeb0AjB0v1Vo23AB7zx5b7N9N/psAxe5kYk5U4lkxks2x4ZEv9l7psP53GypOytIsq
Vr6nV2GpfV6mjRLWNwPJKIRrsI2SHdYPX4N4q+/KJKEm2bRnGZI/EkQXVLP7iU0MmbEr3SsF7cZQ
oJaWoSJ2CmLDCoVhZnOg5hS0h9qPMC355V5ODTweJix4NpSzU5RyaQFxpg5Aw3xLULzELbf684Kp
eV7aoO9nDL+LkRXVx25vw0fCrK9T3ZmiNKOhybG0mFuGFEyOkjf1ptXx51C0wfCfUgZiyaDlJWkQ
HJoZ6j0WMhjInsHDVoYqy+vGlD32qUnx2kRfrD2Cnkf7xIG8m4TIxBsgjRVe/OszF/i53fzudi1Z
ov/wPRQWnGJiWy8+4s3JwtO/5CPEirKb69C1BMKAi7GIL/E8OHi8dc4JdW6iAugLEJpGU71u/LFy
JVfDTWGcgPUt8eiTsiNbcza8HRe+yscoD7KRKCSm6c/6G5HoAaglh5G8fcNYkhtB6ymyLRMawd9P
pVvkMIxn6l0BrrHiUZa8E827bU8mpwy5VJcsZJ96hruxZyLpoU1o/Bfz9pS4VrAuFeEMjfrto5FS
zzzlHpXbvfTB84MOnLo3qjhFq4OkzU2JxWg1rcdH7zPO58H48qCl1hoKfFmborJgyv9uHQrrSAYr
olcWgin+isYkjMHezxqYnmAYX+x0FQuEQkxMcRgTcdien8hhYM+BSQC+9j0GwBIeVCwvzV5R1s62
FC2S9R9SDvUQjmzU4/puQ/9Vj/FbJELYD/qF8YEIsOAPx/AH4vFf5+AoP8IfngV3/FvSuMsjjSQ6
sXoJ202M+/mgR5qMISy7f2Zp6xeocxocl54PiS4xpWJJVZniAkNnJHCOwl0Woaht05EzopJCaPoc
ht+B2gSWE3dvRgbriz9LF5kAmJr04CfuMFE6wZi8O8LbGRj2kxKh6BTtiw6mmp4ndByGlxBGHeRq
z3nFacJC1hV/dsCJ7HjtOgkEn1pxX2UL+j3mcP1ChdtIzl1lvXCSADwV3w/V0zIDO4YotlHWnAfA
n/c7VLQDyVTVFiPK/obgYMYoExtiYwdrI4T5JOsOpoY94E9ghjMusG6w04ICr/46rIO+qtFKXVWB
/0TDA7V3xUZElzEvnAhRDWhoMba0qw4yB4xdbS6njToZ37YAMqxSjjkDzRActjw7qZvCMNnXdDvf
8V2UxLqqLzTRjXDrse9ngGE80AIACELSwCt8lANlaVud6HYiuEgJIZ3mldJGhghNoZN/6I4MWafZ
bP6uuVMjVoqSgaxbs6Ytlg7hYUCrJ+vJaOadv2SKMG1TT34kwUTTmwBMvHZlt2GBOCzujlrr0Teg
aXUJZSG39EEcWhzOlmZ9RJgudejpwNgt7s8hYvgr3URooxh+Oh06OtwXDLTw6BpEL5wmpFxnVdRT
1W+EOX/IVT89m2VU6Dg0hYdfCDQJ7N5lCP/Q/RMvszFlm0qJ3YsHK7jeV5qpj1Dk7GjxaUqgSG96
oeL6LKXFFp/P8oqd6T4IbAqVfBWBBRt4J8+v0pPnewIKqkM0nSrRSFPa/PPT7J3PiaxRVHduQQA/
y6Y4HBGUYv6mn3ORd1tM57azE76wNuSQ65ej5z7VfBMKzOMWinqiBcPIDUw4hCUPfgDe4te9t48f
s1HblJH8sOBXF/Xx1ukDzKf3Sw0WBt3iYxeB38Bzju4Y1r8XMq5/z6Z6X4IoTy6rX6NqHqnev+yP
q2wEMrMmmojK9foYwdhMwRnlxSWBEdBje2lYD0eDJd+lNSiVPg3pee7wtneRjaNefzkEeHVY4ISN
HTcIDjycM/DFUko8Nf5gOqWC/MrHQmPoCJ6Kq2tVTMk+9DEFv11VXDW+7ryH2qWovblNX2o6y60H
PIcV3i6gDmsU3ciEaW/8hPW5KqNFlXEnVA6RTwBX+TIBPVGPiMLwa9zvK1GqbcI0Sr0trtmBsqK7
KpwqQqW/xUQyoyjHD1pqaQl6vyxPEBSOfMGXeJsZWsKUvwjiiV5WY72KC/lXfzLP4lODvfk7IAmq
tUeDn7EUMDyfrWaR8uUZUTCMCCyLviyj6cYdiWYIUeKixZth2bi1javCAKySW3gGmXA/IcoYePXG
zclivftjcG8DJ5C1yrSWJOiQ11u0djw8RwczhAXGjhWLMaPFqF+rSjiy8Lc6Je+XBN2b0Isz2NEU
XJEEPQ7OKMrD+nDF/wi7iIk2td0XJ4tVSE15S4HdwMxVLQwyQMrOJt/0DIP1k79xiYUpQRI328P3
IeJUdrvHZXTkytRXZ+b1gETOP2M9X5OmgosRGjMSrOVnkd8yNsCQQy/p/SDIWMLwKXkYbPrFimZy
/EyDdqDXYP8xOqWloQ8sgB2UTZdalB4kcnE9o6CjyYIUt0S/uSrlbGsNOFnVhlg5XSNqTDo/j8zF
GqW7BApJv3qyOWLUTl/6oG7dbUMrBP9EQ4kIxeAzePfxKm2+DQGmFAep8oM8NOeaWD1epYR6sqFS
7ENBMsjNFG68AfBohmX0MAILDCO61juplBmXdI4XkrUX8DzddyaL3UBdQkMokqBiB5eNlooWcw/Q
wytXq+Z4QzRuiyVniv1sM1sn5QQouzJM3ofsghpTh89BMvKtbzlxwZ6UOY0OQ6PFYD7wTUpxd7dK
gldnTgaUrEtpKj1dpoiolJJBnxz6OB/oIPRT/ECtIsZhX4KzYvHtbeFxPmwjVgtca8y4wvnqNcff
WzBAYgX9Z6IElqoun9LADEvurJd4T9l8LRFqBFOppguFiyHlCAMQMLsdmHSCUPwC7QGXJzcZYif4
alTcWPrnkDVS04zVSrUy+l015JgZ76Nb2ElK2VmLJcrWrnCyoQPOCqQew+etrlv078Yrfz2nRssT
UE9VGEDLDL56TXDnRvr1RMTH9yx1JxxBcNsfLqxuI7cK7YyVGKTcNU6rppuWilKCQ15MVy7O98lm
dgKN64bLJ8cu+AwnOEUglDAOR87TtTg6PmWP5ZBgZvmm1PN9DNQ/RKEaC7RliQSEJBt0Jnmo4vO0
zZtuXpKF8XsKHQvhvDKflL3OVjd78+a2vr58Op3/GG2bX9Ia3HTqlXmXLSLS1XurvV0YjLr1sy6W
g0QTtz6OFSfE5qlkJkP/lEUKWw3xOUeuCQGnZNrvkmx2lSOZRKbDLfYKW/S6ffxqOEgiRZApW3ON
+eYhgYNy9qmuvHHYGyYFHHJOH/tF3l2vweXSJrulkNedJItRsay1MYM6BQG2ezC+zYvBDBl1HPCH
UVm+qKDmP9tzOcdkzRqF12e1chJauORVyC0i9HQjp+FYiRgoBLDR7Hlxg7oaqwa2l9vC7mYvLF+N
Qpop60oGxbHC07FKBLUnvB+asShWdsVK0X6SRdObrBVHx7gys+IWHcFnW3ivxzW/naxRjdYiW1SC
MtNe+dzsh2RuZTVdjMxdu71FMb358q0dulK5y1ltwqeimOfmD/6IKAtpgGaENrUZPvhow1rz8+3q
ht82py6xdVtS+76RNmYc3CmBm+RE77rB9/cIWXco97/fluLVYyC7F3ctKMkxB7CL790Gyv0oPyVN
EdfHEE8uVItzQPRdPeVGD8QQa0POmn6HGuW9zzNKjtn14rsQtRP3LugqO6E+xM/3RzlJYxJUdVum
nWhkAES6aUDSSThWFZyaY7/qMEpXKdIaKJVjXDHmeHV722x+0pObEs6gHJAqKwsJ9p8+YOlaboEV
MtLXNpEQcmpW7glbxtrl6a1ZFl/EH525CehmvKqvV/BAw4Z5S5MY00kxJo1D0NlOy1J++yg0LNWM
hypFEdDzxOfJbYLUBbINsS3thq7R+QYEGJR9Z8nlwsIeW/mMARrJv6TbvD/5DM4S0dOFherFzRn/
utMkRC1arZcxIk6zPZMK7XxllZQzlxw7X/IdqxoHUwa3Dqi8OXsla7h0RbUrUGYlR/JkRN9JIWxZ
wd8AHrY+XAhMtJf9CTtOkAa55MIXNHgQRAlZS/Pj5PBVsn1EszLLLBdc8Cq5dZGvkhmn7FZTSoyg
SDKqGvlbIRouknZUXypIlgkeAOtM850kUbRQ2qhDy3vRZZ9LgmVbuDFYO1Mz9BDGCQAubi6xV2Hw
OrwbBeaXwS1BbF1d6XGNKAgzpC1Gt92DggneqNn7DxUsuHVbBuD+quG4y+GTdqeoxl7N8ty49d1H
iCK4WFMwgFtttNnzAggmLo0CjL9ktA1F8/90GR6KPuhHEG1ia8nlZoUFuxa9vwJeZms9zr5W3LbZ
WFQotl0G16S0ukA9LPgtnWDyu7JxmMmDi8fCkANCwrtzFNHPY+29BelHvFl/20Km3iL/2eH2sqAS
7btC241WHSYK3yUGYJoWEJcPbegNlLQ+f0Ryd1XsOfGzVA8FrkcJUm6yZE16TLrkNmtWoW6VbICe
89iPvpFHk2U0bXAfDFIbD+zpbQUCxaBe/iW5O7u/4YC9mk1Q5xfXdQcwiDFuR78TSYhWSAwIkiWH
1B1jVs3Xz5XuUrKghDLeqXEGqLDQfW4SwqlSlpGuUQ8+NUuNjKCCevFmAWBOHbBAogpZlVnNrsTe
8XHSS3uBKF0LVbXLi4DGDYCCQsLBizLU7ckdGeiinuzLOFFrwt7lndcaCoGkD47Aula+kGwnSzYH
QpONNXZplxzqjN3YbFaYJfmzMdUc75ILV8sGqZfLmpf1DJ9RaCghqZeBcQSXAqhauKxvOHnDFTZ6
pA619s5znGVp/aco54+r1imLFiYSwSe/XZev9PV3EjadNIwci2xXb1Eb8RZ81UkWhuf4s21S63Az
S0xccLH6xKnegNjMfZ/xfzq6G2RX4/Xw7y5QlZlB6lv3aoxL+GcSDwP13GGq6F8I9qMEZb9ciOvq
y6vWCbqYj/eerVVfGFJj5pa/KqgLpzDLq8u3s0bOhL7xpJK2aZLBWmXndaqsHk6NNGU86ZYdnn6N
w9EzYn1kYgLjrITfPRzFX5Ds5YykJ+WRKgobDuB9uPLddZpD1wnSSF2Is2fFXWXt5mOGd3IDDjWP
VQUwteZQH0Gq+ce3SMdCATWGx+6VuGomFFN54FcWGaiTf7cbVV6/qpL3O41AuIvCHmWXGJ9HxJAJ
OM6AaIotJV1LHupvWG8pUAXwKlc2+Egg4xM09KHHaZcbdjYuCfHpo2eXsZVcdQgLrfoRHZIF28IZ
CllIJYOGcfZkg6X1NkFU2VaHzWra0PeXSzn3IGhqWNY0AfLY2sAqFuerCsX/n1ul/MSXYirnsJoC
mIVz6mLQTsSQtGShmmV+ZPFVFKx/Ltr+s+BEfobxvypZC1rCV/s1cg2vdZ6JhLzs3ywiMVf9BeE9
xSD6eL9S6Sn/vZYxEjy/7DPsT7hucGZKVu8TR7MMH1cmvcbB9HXPYn7hr9sivMwUcE9TwTo3mROH
FVR2dNvn4sXBcDZEoohPOnTZ8d1NDIPyeWBiBD8WG/X59Qp5NLbPxIYpQ/G9ly2cEFJgFsphqX33
mpYZGOFM58O2KxFKmIPmcSPlQXm67nlxXWxwiV5428RqE2P4VS7JZuEPrJbgXKuSAriBujDVAw7q
4TNTAEv6j1+p8JNYgIoIJwKjLPHqknSbmNYcsLEVxMMKq1wgGmxzIhNKcPDoOISSce/7AfAtcq7g
PayyCbQ+G5hXFICebTBoEu2WwWffydEaD9u/ENcdwA6oUQ03I3fn4zcDUExjSvNZTxZCUTLIs3Yw
8CBtBbdSnLohGAg6KPiZ0Yp1qqYlcDr4IXceoWgcb6C1ePuV+idnioDmHMvsMsJzXwa+XTiJaDhx
Mu8xbtS7zWBDWQLoz9ivKLvtP3LbMJMiJ5Y++SqCzhvTumsU/0NlYIgmUueV4lnWsK18c0RWOIA3
Y9g0JnPt0i8Xc6l8xQKNq738m4PQAobt0VgpHQoHMf+yYT7pJb+pZdx8Di+YN6v2vH8W9SU2B/vW
Djm9u/0IwVvzQD2y78BHD83eJ9qgyi0EB1Ls4y/mGlV9XatA/V7SO5FNuupEg+tfEdkZylhzvT31
FqWn9BbaLmNDw2gLTKHgdGx5IuyTeJe62QjwXAV7ooCuWJQ0DaRs34bcNVO1SC+mxIo9GoJBU+Jd
5CxYQzktPchXNps8DJWvcJQcP6f4A8chgIqlXw6R5Xavx+5muZk1tiupdzULIW19SoA04qrr4huF
QbEOoa7ALrXpCO1yehwkK7Ifkl6dpVw+818ZBcRCDswRhTqJ8cFW9BHsvibmEOBkZmbFRQDLEezc
nUPieyMPZONRzkMDoSy7+ZQGnJqHXVRuo5xoM6NMO2aL7R2J1cgibf6cTATXZmuciaWoISdb1wNJ
daLO5oS2Vwsj45RhHUskjvNf0QZC20NDO+2Eii+S/VNGJ+xFiEsh+bnkxLAzIRhG+9SmNj3WE5c9
Et5WkfeW3PFGX++XreeMMr9/B7ZqmRbHOjyida9n50VAA93ZL5Alf1nf4p7lTxWHWAK6/BejeC+P
zFJuaU3xUPw2WEcg2/9xszW6Jeg5DCvu0BnHTO5mSMksb40Cuf02+ilzZrHeq+Ruv+aCJlvyldsN
17Od1XHTmMszNo1hQuJDbrdFMh65QGXxmoEBoK/J2EjBdowA4uPBg3jqQzS8/ag4+d8LaUkXJ0Wr
2FVgQjb+KR9Javftc6EB2c1hvk10QacVUBBQoFpPctTwtnKA2jVJ7rF7v28x46xOiP90TqoShuPh
zaE7uoUXMMH1T2oGul1TJA0GDhgncr+S7XudmmAga98U31M4NYPQWmnVNw9UiVAkUW3hjhQqBxyv
Z0oTTzHMXBBIuNEvUNTQMG2MtEMiY28rUQLA4C3qwhEVArqeEi+FyD6IWX5/9Ph/+S0nKHM9nVPw
dFk3Fp2qmO2x73CL4gkr0KpOY9DYRbWw8niPsZ4/dKqujcfvo4qkxo5K6QnW49naE6iUYu/75Ju2
syWUkTXmNc8X2zdfZ5ABTD22t3N/ZPbEvzJDtbMg15d0qC4M2Q8qelW1S4NkbF4Wq29+X1c4du8a
vEXwV9lOTku8P6mzIAjRtG2iSxvkawpoi03QPkki4SgMFWmHUupRDfJd1vDlt3Am8o1ChTano7z2
RTKkz71psxJgkIs9aanqSko43XR7bbif4zNG36nfdF8lqG8iuezhBbdXqwducpsPBTWHEzvhY/lb
m233yCLcTidOngl6BTAsj5s4wne1z2a+Mvhwl1SSNPxMi6LAN1qpbXEijfBGnTxXLzK04jitYhjG
UElUdUmXky/gZtrkEA4cjlAmC+5MHjVKzzR1NxG8AaqT8yNFyixjqSdx0gT40Od1flpc8oozZXvA
6Pofj4tWYeuw5xkLIMAivrL9fIZU1Bp5IY7C6HyEsDqQI3UX2IlNqTqi4rDx35bD1S0KkAucD/ko
Py6N5gPXVvKQc/tfiLVVnpOZfHgh6d1TJeUBJy2M0NAJklJnTVpf/BgyqyF07qnIvKdZkTmsx63S
Rf0djdF41gwXrxqHG7QoI5Pt8v4+S/2z/MR1d762i1slWX74y0dHKdbFGFOxbj/gXfNo1TgIdJHn
s0VulaAnYDVxrd88AORtauyPhxBzuAwZ1ruX9XDmFs82tuckLxuGy/oX/UYhXDIFkSgG3kgGYYcn
Axazkn1WgCgdwSh0Jm9ZztFehxr7iEMydrDAhTweOnz0xjkVdX+Fztg9SlcbtG8QcuEGk0Pf8axd
61Z9UAvKvi75f0qH4ekzjlGKVZkOIafp5pBOke0kl4PDYTXVNVKOqv1Rh9qnAp2ZoVtoDRDqW0eT
yM0526PKYznxmMgupZ/B+CbaEZVJ4mDEJsYVCrt+S8szYhj0uIX6m6v55ujjRf1DN9sv7EUnzqaa
0STwIJNA1yG8bwRTEQjorUF6F3XwE6iEQB9sCEmKrc2FKgstKoSFOJS/tAIBgrSZNCLjSTisJ/YS
5uKmylGtccw4erpQ0jEl/DZRI7h0S28OWBjGp8ROpKMs+5/jPSq+RhpyAvmrVlcNO4fWgf1iUd31
tLT8pnt3t7S1FrPwTtWNfE2Myt+3a0rTvvE92LGP4I5tbCYfAyJ5LyofVWAGYtmXVCSSeILe4NPJ
oFSwS7OfApSR5anUkcza2levtnoEzqzpX2+151aYfoYMgnB5Rud30m+UUxfg9SPkmvsAhDh4nVeN
hTXZx/8abjb+4CI26EeQ9WG/YD7Mr4dJ6QIaOXRR5MK/d43DFM6exkfQ8bhay2wTjLkyCwwAQGI6
x7bU8Zn2J4RFAsFly3YnSdQ+PZ86rMCCzfy9uOQHMTa7Qo/rRm49JfIjIi3bhTw612Wm9F9MlUYx
4pj9EcOdcYzlb6nmP1wCk6Y2UfZS+t21qFeRzoAa6eRTGRclTD/M9k6sVoAXb81Fv8ZYJPJicsxd
SZAQUHFwAQixKjkUQuNlJjA0zz1iIiO477cBB3LaRQTB17iz240lRiMf2TvtDPHnS8On2Qbid4fc
KpKgj08x6S6ET1ER3NCDgXTg0gzwJJ71eFZ6KTtUpFsIWvVyVuwg3AfY5WzoJl24jr2u4mvyH7Cw
a+xrDUcMIIOD5amOgipHWnR2nUxhz3vaJmJCGMBGJkOVtHxASlxbaSuAUPmdKN8sNju2/oDwQKMi
crf0KQMNRMVGOYfkO7Jbnfp/fsWXvJZDeBZ2utIABuMZMikV32g2DKp92G22jdMQFogZnrutWnEv
xudtpOG7S1vUC8afGIswvpeg5OnZkOAzyejMaKLFIn0FxN5dZwjLCEyncuv60HDtxvR5R45QXng3
ezMjP8+MWx5ipXwGyRhh3HwG0uUnxgnGsqUriT/Se+aC2uetfsQq/R5UkNkzp/sJ/O+n/zR3aYxR
lbfRRo9KCqY2Ox5sLFEk1ucPOtUbKQoFKMmtt4ileixtCl0uSZRPZwOZbUDp34PJeMIJA3e2dfif
hKteFcxkAWCP7FL5jLODdoytaelfAqrTHFPySnC9qrjxWn+BjqgdIM1JdYRhQQaKStBN6whf7baz
vV9+yVLmh5J1t0lki3QpiIJmWKC3zR9croS1RZBetfwDPMfzsv0PvGQ4Ckt/os1DnDGqJU6MbgYR
f8VrYVRwTbi1SRAPDPQsjzBRO9ksofQvRBlGN+qRqYIC36Wx12JDt+bQgGpSQSBtRQzegusPciD5
16AoW+sGb+wb0Lft3kiOrRynTQPdRvx9WRPs0YnytwoJcxrZRko1zscuASuy/64U9N7JhPhbXw4d
AiwiDtVYto839ZU/mUvu4g5IhcIfF6QpnFmPrNERArTXDjVBZnfGwEq7b713Zix8tWkMpOJCM1rV
6FPMMJ7NDzaL2bHd/yMkNfvjMXI=
`protect end_protected
