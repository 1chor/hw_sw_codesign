-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
hsdtPZSi5qZrYl95UAkgThpNg+zq9PF7GY8qHdMBtYZl0VySueaQ8FBj81JU+F/S
4t1eaUW5li9SoqZUzvyx/vc8d0Sc8+j5Y7bAI1DkOsr6mipKOFj8Vsa3w4sOuaJj
Z5p/soneiDsainljxXIuI7qy03TkgUlIanaThGl5PyY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 36496)

`protect DATA_BLOCK
l6AmKeBtsxjbu0+nlMQ/XYwk3TzvLyLOt8BfYA3G3R5ZsNCwTfpi7xjOcJXniffD
PWTznQSAhnU71LIv3bVTPj1wF/fe3BhNFnu2BTXXQkkXVRoAHtJxn8AJU09lgoRG
7SYpyrGtk/pMW+ajWcG5h7e9Eb/uS0j/jU1HjRRR78O7C1VyJaTMJs4PrkH2pWj2
HFN01h6pZOjbylll+vciqhbHEH49DmYah4OxvC8KCpFHyyavBnzAmAUOVhrkN1XH
mYsGtYGqf/mX5M5uIZXnhMbsSFSxhwq/w1iEEb+6DKyYqo1l2Dnl36JWw3NgGpIX
PZi2apuYNvD+RMH9kD+XZMPqVJOB2RexqIE17mUBgYI5VpgGS6AUoFK+d+1AZhmj
gQi2QURKOf6gnmdF3mimUsL4q01fc4TDXdPOzH03g1i8B6bKzBYWI9DMlhsqocO+
PEq3wr1dyhbCtYpvGbuUJ4yNa6UQcGV9s6IINMKewD00jLgdYKhf0/qVkwHpSdzX
i+kPisEva5lvG5OfRCWPPZuzUGIYM8bb0eyNOQH9UM9Gt2pd31YQCuK9+CjMBKhR
dyAvGM4tyCCQBY188ncIXg0qeQg1N47X2h1gO9fS4HsXQCyMv2EBALyjPF19nGku
nV5iccgCQzESsIIWg7fLLkwEYBvskWUHkkoTqWuPMatqAy7DVDJ5mY862PwXvJla
tpumDjrIVC69qq8Tu6Rph1qnxBfQeQSH4LFDScUO2fv391rGKT886xb1jkQqfmru
ku1Y2xYiJqHiIzRIMhPcg+Qv2CKSr1YizjwrzmMB4JpJH9PFY4aOv4TDODbTpjyk
bx2fq0TD0gYRy4tv4o0ZgFoyqEZVpHOFvQr2u0QX0nHTpDQFpKeLrTFPe7kjF8Zv
3kzBCD3vFa9t/jLVsNhv4utE11YpWEre5sscAm8aVSxiVVp2GluJgyppWeFNKl1s
q80CvswBXtW6Yf8OdTHdla8s7xs5CX+neyhHxTsgAd9zL4QOdjdiX9vHy85Ivul6
OjPCzECOMUsdpNnJ2E4gnWgxHGwXHTQjix+AUiLXGIyVGoaDU6oMRcR7C3DWzhUq
IYfY5JFcCRPfZ4syGlsr0yScPyGpCKsuR0Mn/qQv2CnSoTJdErzRlh7jy2THJkQh
xpPXolKxOwNE9YYYKWXu0gaSY1gqo3+YuyFI5nAzchRgEVXg/T8N5NzR084YtQFF
iEOAv8gac30yLgJabciVD2I09fJGTmmx4rjv1Sg4MonxhOcLtgyX+UdYeO4cU4E9
7UFgySphmnCQcWK2wKshNL+gNZHi99GO/yXr5YqJL9YuctWpQ9sFfl0g5pEZja6k
SsmmHULU+qfP+jAkxxNVG40QdbNExTc5bObXH6p5/Se/qJggfyBQ9/fWOPCmQlPW
6cEQDHjXbgRuhEoKX4/VYrMjiSn9JuSOlAB2pZqplzXvTmcDybfhVlFccl6vc6Of
r4VKVXLgz9K3jk2zL+/tquNQlpTM1T3MbM3xRPoONY0+NKQTn3g5BBq1u8oHsCIL
dVB97aTsUMZCP9PAFAJCFTktSFZ4EMYAvfopA9VPec1mnQMLzRMMiXasAfPZ9LE0
BVdZf5NJXz+0MIBI9W6h4xD0D58xr5FfxV9RtLGVDsiUzAFXo+uFAV10gzXeblTR
ZgWF/ZoVExdWJOeH9gw+RWl8KgL/A8klewfpQ/Gr5VeJRqhl/HtWBD/EfX121t+w
Z6EZ6qgMms0tcXEXF50QecTNMGXEiVl7J5C+VCw6TWtV6GIWASsPdGDfGePNYRyK
c0cGB1P6t6K98TF1KaXY3WWl99xTx29bFG1P31EfvQlW5mGK5CEwal845r6uUjDh
XJkfAB63YyRasPHRVU7GKD/tMn2tdUc6nr02V9kzlIB013c3wqp/FSThqDYIKdAu
DpdnwCGeWC+17ELo2kk/tszcq5Y9lhTb18Wr9kXuofjcYfS2zUGq4P+o26DP/0nq
PgmA/mpgMmfZwKA6UbVuwcVeHphqbbNOznzYTnxvqK8a6kJtCmv7EXvCZiCVMhFB
hDaSG8atQ1JxXDdRrfTtXWYkh2m7AdDMbB8Sd3XKSztzHfMTBsfu/mlwKTo7lvlM
UUGOi+Y2trsbCfjZAu09BQkPBO9Pp0x0CA0rkQ+UsyYy6/GKyNwddZPJfwE6CpOS
t0/QHDdKYwbzR5h0KVrsrmO398TGX39aAtqrqGSWanqOpzQmiVy0X5yLLJCdrGPV
rSJHvDVXV27w693r8DN/wtP8qPneAj4EF/fG8cA0kqX2+sGEfJq0jPCIjoAoJ/Rw
O9zAjR6RhnR5ae+mMnFcuIr2ap5qOYWezzsUIxcUsOKFzJSiBzBJ0aMsYnD6kqPb
lDO/QRIIFW/MjM6G6+1rAojCVkToS6h+edG+5kfQf7+Yg6pz0BcvWE4TzEGD+SRG
6z8iRiyfFOQpRclkrKxzqX/sZTNz+s5eti+/+GjUcDJaRHtohnAw2BKxTWZSfbo5
dsxIseoBxnjZMzReIb0StDvFxVQSP3+pjTBGE1yUbLmH+BwalO3jPGIcqeJKGLnN
f5GsKbtvNj2tEOlXP+GZIj9MIp8HwjG0sBzqvMkzyy1bPZjphcSfs3gLDZ7DVJtB
MCcvFo4FBQ6MzyxXtEgEojjtAcU8rO9uYSVdgrUgAl8J7fCs3SR09svEZ3xdHWDA
XNNzjCC2Hlk7JrjKwIaLMOvf2xD+x3TZVVxugjlangamkVSp5q3Tpy+vY18lsqB1
pvTRBKinxv1+I4QdH9VBbHPLXSRLnnAHI+hA+ZamloyxbQWJxk64yl+JyoNOE1h5
ytJC/hoShgHH4IfOYNt7zH8XJDa6hlLT4MD6Bz1aVYNbsP02SH37fX2jF07fIG0Z
2SAWI2+JUg+NovjOirbRdtTcoXZYP5pu5qBcmKKkrlxsnUB/2s3Q/BQegKoaJSrV
YlPP7uKEH2YxUwwW27zgk8ynGPZBJCD7ZWUD0tle6EO1m1HoTf+Bu3WnLFTA8fyO
EezQsMHLfiG3+UzrlDmXbUhFKNSV2LE04poHSyCENRU3DYg4VWiGhWA1N/rYefPP
9BhUd4+KILP5SFRM8WrCdpOYivZycKy79/o5cEpZKJ0sV1Lu/ABABExNCK5r7PCq
CiCzE4g8RuG3Dt/QINQOH7ujS0wwon4v9dlUpGQoJt7bvXTHi+w2H2gfgzG87imV
tUGPWsAVt9oKDKweFHthZr3cPMy0njCE/CQ5LuEUl6UVfKVLyfvuWoNT89b9MVB8
Yz70XRHwvKM0hmWifuW4maLVjeA9VeELozHUvkbfmVGm+/vIZPyY4B1YXNNnLWMd
RU3fpZbeZ4Tk2o1my0DxXmL/kEFRjEqRzKUeeXZTKAD5qD+wH89V5eaZ7danDWqK
fv5W4+K6zwj/LT98rU4iLJxamw/+8u9bjttjA7x/Z8SNSZeQyXe77oMv2hvhchZp
uZSzGw5FauYfbTxr6Lfe9sTp6sk41M/p2WdHaoo1M717swozKvYmxe1qdOowE2Ak
HZCfEWBh4gJQFq5r1piqOQOykHoHW+JHBlqP1XMaFoegCUBrOHC8AJOQfVyfjTFU
JO3+8jX5BMiVfw/3zWq8Hp5/wtymNixS9eZFbLa25F/ShtR7k7pf9oCiCT6pD6kG
aOZqCz79kwPlu/+mdQh5OD1Spt2myUhsVSI6KjZZu1PxV+zXRN0esjJNDJHS9XlX
a5yvjwZxNK5mevuOm0U3hgmBa6wMCP2TVrfYO5QqCQ94Yc+7mcThXsAssAGb+2DP
nX+se7l+qTtfTV3uhFYjxYyp2Kt0yIX1wx7VYdUU81VvxGGh2gJSLX580Tgl6wFP
Va5/fdQUCOUfLRiX25dsAI3C3PlwZQBEaKRV2leBDxfRUOuZFdJ5geMdeUZd46bJ
5AFs6EVDVbjjLQg13G5Lx/GJOVTmBlcjkHatCCuASXtJf7jblGvlhklbps2QebML
Su/MmboPm9EaP2z+5V/fFsCf5eDd/SPONevHzrgMa6M8IxWKrXkjGZ4jBzmmklOc
V4+3nd4DOjp63jwvZo34FVH+bD6z1wv/NPcHhmgOMfJ+ASHJ0fqvyT8EpnuLCMAG
cF/qkuCix0syQ7lY18vOxdJDdcAFZERudh4GKLEnvs4jaH47ptjK/QqZkkIUYGzq
d3l1QDZn5OgL3c3YaBq6rKyeEXKJpvSAFjfqIGVq3R3chveVGNW5wR67AcHIP3Z4
tTWznzeYP6SVGI6jZwhqLS07akv3D0DHdxZuSOQmlBqL4EWTQ+jeDSbx7DjbNZPO
esFvAcDuiAJh+3i+UC77cnzrh/GCBGhiohhWemZgW1Yt6H7BlimrubGKMwV/SLhj
NRseJDwFHR2MZevLpZGME4/vYuKe+/oiPCtQX1WWoE/gleNKW+uBSCMNbKfgVB3/
c54pbC9YoYUwqo+Hhw7TtnR8cJHWv+lzBujdK+gQ6DLcG8B6cjg0bWUj4vYl7S52
MjW04v3T+eX4hfT0YvHCB5kUOhh7rZagx9zXMfeJh0Z5yQA/wLDVh3gXCHgxd/Pv
7v+HT1ni5y0AMOTrZKWyqJxXICcAYDZ1lMPxGMwkb+OWP4ojv/N7W21I4jUJnO12
+ZGmzXrGcxC6Vd6zlr8iZ3insklD8TYgRDFnIhzN3V2/jD7tVXEYl+W3yv4Uppyi
4Ya4d9E/tTcERzIXSk2D5FCjWIWg2vzYQmEM579Q8yDNiQuwmvBviDyufxC4uSDd
6l4c/vJGswz+e128wwVNC+ztN1i9xAcZ50XQ689KO+YdarnqzKEBcjuSyD0Kxlbf
BvLOchLCCSAdJ+favRgFe3lZLHL6DqMcVLh6ZmFy1D5Ha1nHEUQH8jQ8+Ex4o7hr
o5nZbnx3ExFHOk9tcV+zpRw8dHG43Z1W0O+OUZm6Zhh6fq+iamHWH82RPWPS+mD0
piEEPb2pNGbqNh8qFXk/w5VbMsIGxsPMjd/joet7hlXTkmiM3dkyVHT+r8G9GvrT
VigdnZQsU2n7XFAV2V52QzwmqN/OIjUPueUy5gTXGnL0qGd5PFbzMDE+TsTBU4tt
xs97K52bILwbCiv4uy5nq4w2qQDHMECRWRAH98w+FAta2cu+uOaQKTRNtOTLrBTt
EGwM/VOWkrl7Drr1+nHjG5wXYTFH2ynoUUqDO3O6U8DuuJD19nhPPFGFqy+4QWat
+NDQ0d2CeY7uBR6wmiGTL1qsqmTbvuZVIn4v1uX2HanlJLZuGSwsrI8jMrHoI/eH
TKyVrABvwddgGuHMWhEvDSepbi3TvqvoYtVihZEjfSe8GfmEEldhy9DZ1VHIe6k5
J2DePgBgHBgNqJMO2sgkbPa5sMo9L5KjD6TOq8Qzn8mu5/hDCRYm6c+DZWvzvJvr
VJp85C0VLpl/qPDnNnQJi/gtIfYOC03r2oKxzpXkZHgIBeyqPGU8jAdE2/ZrJZ0u
8HRdD+VOXMRHrTcjjerKaASkJQ1jGiLVgrTPZ96gXud5RvmGUQvtS67/HECwejUR
N4xtRA0Nlf/qUMjD/XMLPlMTrbEvq0XJOGrjLE96Ve8smPjfNd73CdfPejiz1E29
ucIZv/qr0qdQv97b8/TmAlh1AkD9IJ8bQUOH/i0164SQPqWDozgjvRhBj6Vkc+fQ
llJ2jKYQTFXOQypoUrMEllYRc/310Rg+yECQOqCxhBsoPakTGu5H6IfXz/uJzse+
ACGmPVDhv8AVWPYeefENsoev8u6xVbtLgWr7B9kL4sq9JfqfpvBbuzB+XKwPTx/G
yocbjHPa+pQs9dt4+FVXptFr7GEu89H2zb2+7HdNIffn1X/DNVvvnQSxX3AkNuX8
iktOYNEYplm4mcOsqjRPIEiUOK85YIeaAukCNZfOHyRPG7P2fQH9kjFQWbNFZZ01
JHdIcC0cbEER5m9kHKqKyslSEvBKZOpjoovxMi4+jfKN5qMmizhDZg4WbUp4Zi2e
kiqJiKeLX9qFtCHwpgo/uh5ayn9GmLlSuXpaTOjfpZSoDWcXotaPy+OIM3qS4Lig
rSfbcDXaawLP06XVb6C+2KeUQuoC+wuoKh+BRxChJiDLbaZMGcy6Tw88/DdITR3V
B1ngaY+u2eRInrHYysR2s+PjZqW2i0kTp2vYa5/nxWvyNMSCgXctCf0/WgKLUhLT
1CP6eNi1NKJzO2v3Kzwo2CPKKGOqle+pJ2wteQr1/u999vzkOtZlVXfom/4GM9Oz
4vegJiYdTpDlQQqJOVE7hcknUZQlXUDQHnOJMcGNSw+/MvfYKBWDBCWp4h3W3Ik6
7CDoaeAvJYkmJaXgsPFcrHc9417cTmAjFBGd1NGl6xwWg3LkrdbAybh5beGhvax4
JFGlrOjZ5wpsDhlKUoyWEFTy2ezXIMDRmqwe0ts5K3IL/dNAdidiT+1itCDLPouc
hSlQYgmUREWTVd9xVp2gEskrh3xl8xCWXbo7JyvpKGNzSWo50mbLBZitvWDDucqC
Cw3LPSFtWQsYFbxuUB9E5+wfqcY1OTIPzDUQRoIM4rlIy+Imu/XCTkCMqApsLQHY
IBlL/QxL3RWrz4jG/OVjjr1xHRjRm9z+58iZ4QwIoCrw+uS6IOhFDJNzjmjlOfvK
KVkqB3EWil9ohMgq6QcPkrfAwmsJHuKR6SmGjc0BKTDWqxZ6p9+fFWqY4qwPXkfs
E2n6oT731wRC+5jeCzw2cORGyeCBLR6AHvNPCXkWl7YMsyx0qZDifnqkw++zFDEu
MSWRcU1avQqg2bfmqGuKwVAxHWdaHPScf+OuYdLzYl8PivEO5NnU1ofE+2qpFdHB
OzGP78urvne9pO1iSrWRavOtHcymGMh6Dy1nApAT9v/3N/V+rRwH3KsWW5Zq8mgd
0CNQrmNBZ0AKVJKt5/OtfH45w1z1oOCq2vqEKd+Czbvcz9dIzSBDntki+5HCn8Mc
Aqv8vuLFun+HWxNMr/6QHwrr4u39XVTN+e32dUiiT4njz5qfrHk1SrUOdF6/MFVH
ClJ4v98jaQny1VMAP5tifBgBdkPvCRSaWeUeb4wjcoG5WvvV+s97FUfGKhxEjZZS
z32wBv7+qX9kMAbqHUNbYnsbJSoD9oIbWLyTLbEjgssvzFtUht4+V5hLeDLsROes
R0cyWD0mge2scjfKF0nxlPtjsfKmrTiXsb+QueumNjFRjyLHHK94/kWIdIyCmPUE
QSF7oGvgyk6RKEMvqWKjeQp9MHmZu8VUsfemXotFRxKJjTQUA9gM0PGD6/TwYZza
BjxvM+mGNnK6YEh8pNb8oEhuIOjcKE7p2FrXQlGaWwVKBdxvCH8TYH2f2JbPeEwI
C8evreeUfMOknkAeOU23Rx2Ps8eu7e7//zzsFPxI7TVMwgLws0i4xswB+ABko5b4
zmZgsRrf/F3sY+8WNUR5KosUqEiSeU0DhLg2PiQfhfwxC1QwcJd5AzwNDQcTHKAY
t47hkoVWHIvr/BbH7lpoxteUaw7j9bN0I5ZKX5Ene3WW61IE/0r1BwxJnHu9XzOO
XYx3NE3KLIPXyi7ofJ5kVPDyM3X40EqaWXSZjZO2XbIVSGEA0tC/sEHvGvTW8afB
aMvTg4Y8y/Pkj/AquplHPp98kLyTmfo17nneNNDUEfuk/ePMLD1iNkU49+UtAYO4
5AWkNQS06djsozrMSitxwI+IWPI17MZf4gMTyEZR3RAGyr7Yx11JedzGD04UKG4I
cVlD1VfuLOtd205JAQZKomTLlSOT2Usv0nj9yh64IVQR7L4wYLZY+edinDLxLn5P
0iDzVOYQu1TdDsdmITEUDLW3MfGXf9dLBkcIBRAkvVwHJAIs6ioT8gi3zPq5L1VL
CyynxNkq4Cl/9nDuoCO6LRX3ulfqMVvq8Fr6GK1ySXSIu+1ybsN4iTOYpOmmEHs/
b2YVIMRhdfuQci2tjogW8VLL6pV6UnU8YM+g2FRiq2qXNJfB5IG3Zd/2g/rnfS8j
1n/6I/YD73jiQBP2GYvCx7bANfqm7wTEBuAEU8PvGvJ3ujzJgHjCJz/TEPFP/SLO
wh5QnuuQvrP2Z5tEAvrkh8+7LBoojqBQ8A2HLJtWtOei3/kntPM1lvzuQx2v9Ulc
qh+1D96pjtRB8QyIjBIv29/G6KfBNy2vaL2KS+WtKEEUmSO5p9weRcdo/tUXmvvL
6dIDjLxbqGRrKxmuwby4CLY70avI41Thp6JuWERhynjrcIV8PQtzbi52CJDq3+60
MEPmNt3pGDsaHdsGGS0ue7dF5IIew/Fyj1q1BF3HXJUM0VIAgQKAFVl67YDHaYCB
Een+pnzn1VS/FS69of7eL1YjJ4FhhOML1oxww9SGUC0kUg1kfcU3w4unqAAk+GB9
Zpu6Gmk/qutDu2+Nv8Yjk5SMQh8NyFdc4gZ6/WCxPHfVPnHLc/RxPwZacU/goMuj
AgCvVvTzCr7YRsM58wPx+xK1TpzNscDJmdBkzxGeYzKFgHLdAGy7/EonaPKrqRYr
NmjmIFZZJurSYPt30ZMyepABJaiQALUb3kiI3OyfZ9mDwWOv1CRfS/LIVmhNOVJy
HfcCCGRKXcOdI0GLk3LxUy3YQ4LGAm+kpTST3qVbkVAypBRe12aNVn7lmUFzk4Ps
i9inn6nFVqY5UnnCE+iYC6S16OOYnVtKvfQ26Bk01FcDOSRXpuNacuFzAxCwHVes
qqP48BI0sG4uzU5/BFcTiIQl92/Jb8V+kkKP7yyZazm1tmHAQQA4uNv1/KTOJwus
lALe45EDhwgF23YgU90g5GrKUhUJ0uuO2oB9GJZmWkECtvReo+F5JTEUf6UgsZh2
833pPgMHS3CT3cUY/3/5Vv7kSeKGQh3AarTdm5okXm57sKqFa9hN7/WGp+agY5vR
WNwFVm4cjWqiUglN9puhyEtvHuTk1kw4MJRZVzeXebEWIb0nK0EUcEh4jA/9UFNS
t+V9oTGwetcWef8EMZgHB3CZGPegz0clN5OXJ+OLqCLtcH7mFkOnf3n//zNRnQjq
s9zf0BUE9CRdc1reAA3cOA7YxmJkjpjEPMsJHpuWSK9kWkyAlaa3GIK9oDUS9d/v
M1kttn5TrGgGlNWj+3PhtgVyWITEavv8Qmz/CYDmsG09WkCodWNC4SEN45w4w6Mh
mSFaOAs8QI5p+vAbDqRpN26N6BQsSOaWKoWWD+ivNJ9mtBI/TUCOPp/TjRBDDrG2
4l1X+DquuTlMcyoJQQj616tY7yiImpgK28NhdK52RAbUWR/8tD/5r2vJ35OFKWZA
8HlGcqYNOkEpGmhk4JCCueVflGUG+PhY0Qmd90+6QxT2WROk/kqh2Q8m5btU0fyk
o5zhQZ5YEqXFZbZ2xy0daDffLEzRzqMfqzmQodYt5NXIBSkMmzcqKQxHfnyx8pD7
l3sG7F7LnWd/7DJKVaRphKsDGVPXQXHAmu5iTV+LwglAu9aS6mNM4ko3t5tbsjzS
XCTkln9ZR88ZeJFsRG3UgisfYE1PAK5AYvEC3KxS37SeC/CeEly6nDEtJHMaGXI8
Ap9/A8waVzu71YyEN4CC1KLgh9bSbtkq/kHfLhxwU50lgLqDnOCh+MSDCF3GjGMr
YSiiSO8346upBMXN6sgkXrNEFNZEQVs79tgamRS5aNinhgUJkQtKCGLtLHVazeFC
ynDGzG/tmyKSwYRqusAOxozB4YigjHWNA4n4DL9qYV/ELUXX3TIlHDSvpyQO4+M/
2IHzfUb2Y1WXV22lOozcY+UdpJyZwlW8R+P4dSz5FQLEY7RhyS6snWHu40jUh/pG
3w+vWpQYyVDgGImARbrx8ENM9TVBsUMA+cX8ke7+x1aA49QiPAQZKmFUmVhAiay9
ng3Pprgtsb8xT/5XYcsce+dRMuQiPd2diJLT2V9qu7Pjv5NEl8p/bnM2dJ/zPMkv
77YH084W6HYaR2heH5B+HYWN090FJYBCw5hKHYljqGPN7nG+kIrtkep3+nJfE6je
H+La0JGDpzSsX7DhPoP6j4MDQvCyaKGz0148eqSKEJUeai8Mhpqs4ur1wIcYHBLi
+sVp79UXLuinyZtIyVXP7NIX1vMuRLKtrmTzyBMwJFZKaKjrz/vuZswvEgTcUHuH
8c/2qRs7P9y2j//H1ejPnsEDWYRwfCd6ZY3Ft+qqa//9IY87LWIO+7CBShiBx/Fg
NhFSdmOfHhjCrpBuY9lCW7y3KqBLH6ycLMX3Ii0+1jXzhz2ZVZtKNc1ASOjLGpnx
VgOyC08L6xfNuw2Ta1iIanuJgmt263DdZKvkotNSDwMJecadC6RnEp7eb7QGvGKW
J0sanMQWYLkXmiLYBjJF/HPiMw/PvC615w6BrK7YI1glMLV+pOGeymo2sjz9R8E4
Zp4Ggfbu1FXIeJEzDXGLca882fildYnYSkQRKE+vvwVjfZt53SnIQfMoecidB4Lg
TuPpCWC6/UA4Nh5ZtfYAlHvTZXPrJ8/ghngm3KldrN3xgRFp6iRE20P10JAumBie
4y+nxPNhVznnmpODox1Szt3SODRe/drdjWD/nYKnA/yBZJtmh72SZvRrm2L7LpT3
7yrE/FN2Nr2LaKD6n8fZBo6gD+2hY7cTHtIWTXemKNSkExnRs51GNd3xI/QIsREC
Zj6a8OFSuUa5W2VCcf4HH68wLEH5Kq5QYmqTidDtsjifbgC9pauE8iwj4zDtUruI
3np5RDDFdbfZ8dBnzP7t7oHgH8dquX3v0ENt6vGO08DsrDPNkgYP2seWhUnTDgGJ
N/5keRkZZpnt7+eUH9LSRBkk6Rq8g1f9Pz+D6GNyl93dO66qCJMbI4IFfE5tYx7V
Ho0J4NjBWTzBceQBWSEaqpKaGpL3CTSklo+cYykaUPL3BA/oF1DOx2Q/btL8r5k0
PCrui9+JWqvu92DCJzMPNcuoGFfd66vfAaj4ltdsF515SJ3zIJJi6oQrMPWUr34t
KLm/WZULUanMMI/uwvqP+QI6okYenjL440R1sj8AQeRdEiP4w8+Qkl46ZCc+Fq9+
gzasfLbVjVigQlDSqbG5rgGJP9E7n78Pc1Cz20vKWHMwV50Z1oQT+DWOGvNBnUnd
sJ9X92osDpsRRVK77yw0wQE/jUyOlXEw7KTyu/pnQ6qOvamqVRYUSsOelSokYQgL
x5ug357m3XwULLw0it40YmaQCVTJMbYnxq3/JMEorlKMPmoFP6w4VbBRw4HnqAKh
BrUbWkPxe2WMUTQNQ+gSbpnwdfxvgMeql9fb0kmbSMZApoBWas/7rwn8oGLwJkpy
bAB2mAICz8OlHLwM52nfKqQpYbWBhSVqUJw93BAOExXzW7j6As7gN4rk/47ef/IV
3Az0zclJryE5UBsICpHqjLWTSRShPDLqrLtHiZzA1Yii3Mkq71dzbUYSd2wsciC9
J4TBTr3/6BWQ8C6/C2Rfb8ZfP6W1Vq4svZuhdlemO+J4QnK3OqfU038Rb4HkQlUZ
9vi9rV4t/OX5BWWK2mOsZ5m8dW4f+psYq3yCrV2MjJe7RC9grFosAc2JbVk818xs
O+qXWl7WoIyJELZX2/lRErMwTcvsprc7Ihg1UWQ6K2Qm9YHN9JpWkfqk67CXNFcT
vJ5VdnCoPfx5jys4+yvvv782pzId4NuM/2cd9Evx994DazQyp87dDmuBPa1rzcDR
XP8t4CDbJZqpJQtlqXGK9EKxsrtEGXidcOtqcVS99ezIqN29b+JmUG9n+fpDiDob
x9DuOJRT/wcQ6dkKRxdLQ0fmGnGszlUYek/uSPE2dXk+N9Aw9YcPJDbUWZknj75/
vEDG5Undm1wFSQpeW8dn1grG1w73aV0GHZs7R5Z+6HMgxQwySolljpFrjaT8DyRK
MVZHpbFyC5HppYQzS1Zp3sXk7H0xNnd/cvP8u1GKMu0gf3rsNZtMtQGl4caYiZqy
AV86DG5PrAOLs004o3F/azlPLywrbdMx9R5EJMPUVZ77kgnBoh3s2iisFrFI4lGd
EbGTY542MvfT0kuPH6im22dCPRofOQm3MG2jFkcs0Kn6kH31JxwrL1x4i7TZFFiB
vqZaiLncoCbZRfJZLe/sCy8pZRHCP/Jd+dnfT0vBKlpG9w04h7i/tbCrV3YIMhZS
EwO+8JF33HGxytgPqTjM7kScxoBo3PdHbiMQmltrbCUQe4mehXzvbQMTy1tLAg3I
wrcIxFgLQ9EsLBYpoHWQCGxg0vEp618CIDv3BPiBkDyynoBjTw3IqBpQbumFh7ua
gLWiA7U92wNrjU+kuWwAYOKJLCkqO0LCwI3bDe2E1jTWG455MWyCKMqQdd0X9qkM
LiKKnxyrLAfV7dBZie0kQaswjNpOy8KO9P8etjf6ePbsY/S/MaOZXZnat2ZzgBUt
xPULXR91HTJzEBhEWnYhEK/aFJXA+5qpnZZ+k+0YHQOV4/641e/8BSYQMeIep8cA
jGVirLxBq6RxM6frjQpFjC3OPDX9rOc4sXyW6gfFclbCZs83NOISKj/JFg1WDP2S
p6itXzedtPYLEFLCMF/ThWuBjUwnodhVv+sqW/BA/OXVTcshdEKZY3nT7V+nAmJd
f4cEwIDDbxNMp+akFsoMQzzkJHUzf3HaG74RxBxxrDmjs1cw1BcPPiA0R43U51rk
k9NoMY8a5Fh2WrDYCgqyKDFnKz92MBQoAUQ6NXgnvg1vMsL5/xCXfrAJab6IDW4z
rU0j8JKDQj34NddxQgxgmErE2vdnDjaRD0PB4TbRX4jHPHGt/X0aw0qbeyj0S6JD
NKIRu/H5HkuVw1JVkuccnw+SiAsLjMVekjU4ihoBFYRFaByYiEa1wP403moFoyl2
/tjE8qM/bSxSWAo0BMd0mrERNDysEiTqYF9k2j0bhX/Sx4asNbH1M9uynnCMojsw
fWQlgIMe0uKq4HFkOX0bwSQfTgxkeDkozGbNOAGNsjvxJy2Qt16/OfnHGmXmSsYZ
QgnISCyl+PclE6pE4lZQiS4Headha8LJz3qPMOXIHeUQmFPkiUQ6883o423y8rdW
FMB4HiH6ZTn6L0gX1Upgn/mBg01RIooOU5VJrSDuKTvdc8BwRMSc5M4g0njt/UbS
tjrDNra4bBwb9HlQGxNi1+ADhnYhS7YGKb24d07MrY1lvcWIgArZ6NgjXMchRmD+
EgV5phpXEN3rXOHkQptbo8uEGuulbUQo6s/Qszi11IN2BOq1L0JN7Vbz/15soW+m
XWJRX/BWc+IOuTqxtPPBm3E5RTpICNz3JaLvRkDjKkicbpXYjgyEbvckKqQ2gjCg
GeUJ/UR8tjxdBz/6D53KwplT7q17RPl6H9F5FKSDxUE9kX7qWDuJP225nKMJStih
HvmXCE3CKqqGK4XGJaJE2MjLzXJRHzzyIQ0SFV7Wi3rvBXMVE9qZMv+8TcqNUOfz
SNZc25A80yCVXYc9q2sgzG3NPqme5XVl/ym9DY7PxRF7RxTNmGOrHyIDM+ICNs5W
jN65CZOLvowhRBuAYbFsFw0hoT7BUbYDg04QC4J2CSgkTTlYRYeAtdccUcbBXzaY
Yj6pBMYUoMUbEbfUWKgV7M6UNN729KXnts+Hds+FAcm8zYZr6y7Y1u40fBWUsWIx
+j/MoYWeMysSQXppVoSXoVEE5GmDsXz56Uot2C1/DpZoQHvORKIO1zCzr+TtZMpK
tmUXDfYwA2isrUZ+9e4XESRiaio7wUsgT/15EDGPtTOiVfcehvTQc/BcXOtywkTo
uHIkvxJHccGRgiOzTcZ4RycTKS+etpEytJoHvjNSLTrU6YBAUwKLMUo9zfvGxHny
8NVJbp8zXAZnOtV/T+5Q6pd/cdZycjYsKB4eFz7ybTYfv0qZ12QsuXi2VpNaToGe
qa7ynEMbVZLR4Bmkgx2IQPpmBtykPFEMj2zLI1di4HUPtJog+Jw2psqYAsxf4YXl
pMaAwaZWDbwkXRIiWfV7Mrgzk8GNJ9e7b0dC16i9kPKLIWDbqKcascYPDVScoz1f
42rF78sTl5qoOy53Tm2EiVNOVIZIbfZw4LP6hTq/MwlzH1e/AvqCZOiRHPNDMnIr
vi5Wmz9YF7xVP2OUDK7kdLg87kCtxXwXdrRHqKhoMmIM+w7P9xz1Il0FxYFGHDM1
o6KU7YausE3kx3phw1HEiTOI8RMOk3ShDqNNBlP2lim+uiR6cu/eNWoURW+F5gJi
UluoO2jCO2ZLnfeJ3WpySkAYUgnD05sMDGR1l6hEIyaxkPUQZo6yD8hs8jJ+xUKY
KBdjTpWf6q4aIEGPLS0HJTlCDI3dLIXSOAYS8aprc1R17gasczddFtPqj+xIhKL+
kJdvMD/YTOh8ATeJGUHCTDX7syXZBdfzA5vDn49nmOLFX1ErnNhtIo16Nqa6Lq4R
HgoChD7D7/KGs/W94a/OZTeNy8EAW+Dd3QO1yiXQjEWyYpmKYm+mOKuHE78kZPu+
UV5mYHi+qrT8sldJYPDVnKytKd1Yi/k2h86wlym3f/VjhB+R/S4XWf+FuZV8Kmau
vhIDyxf67BFS1ctH8EvfVitG/5vChg0ArNUl/TLkPt3g5PKil2uPGzyh4QPvQdCa
HXDpw0fI6WUSL2q41IL2ap8Wvgq1MWee29cjr2QXr1IctEd91aqzh7qEwULnGThz
hmmO8Z6kn0TsTWwXPLq7AGdnYB7YCxBqte2OGH5qWcKMESGcobtNrUBxs4IPG0vr
6YcYxKpzt1twRoeoC1bUQMqw4Z0m3wwYgtoSTAAqxQYDJ1iAISYPNJZg6JLf903u
svG0evdX58MUvgx1gAQQmHDx5tnar3KcHuDIi4RBbYXiuYsCS8t94ZEER6AxQRa3
AU1g7QoAVQA1FYqLcSDzr5y43oajrOGwKdFI5hZZ1/wpQutE979Gn7pf/SbESb13
x7P+yw5ismuMVq5Ergy/PwdaHtuxMuVyuhRvJqhrCynZ/n73OMLUvlVh0f0ZrWso
gV5nmQVuQC+JXpb0uskZpgGkIRfJHqRUutoq7YZUKxVxzOr5VLD9TmjAHj9X9Hwt
MHupDwY8KwsrAFvgkabiTHazPLqQogux1cFLsCxErIHIaxBLU+1wEN2gzx3iE8qN
gS64kTZX4SFMi15hGQH/EbjwxKZhVThmtqjYeXdO60sUQfiikoe+vlyfpvBtksaV
w4qgUK4hNylIjULHIi1kQc3keIIPZxYFc6/Hr4CJv++TAzEJEiRi8sO6/HMIZu1d
8itGeTbpGCbgd4AWx8dwYQhU6M9PyAeJEgvWQyOs/6nrFv3wj/5Z49av81JxUqJ4
LGr6JzGzHF/ydtLmkz2JjFqVEaw6PfIfdkNJvwLk6NfJVqiP5+K1UyEyl7mapCPo
d/PogFLdfFB0TIGy+JBonC+ybwE/TWQ1juITM5l/ES0j87122hby+ZAGghZO6CIW
7XlaiFtEFoDYSAgb/dQzXip5h6UMuOFnLsX5Ztf1Dcj+xq4DI0uB7P5s+jpV7Uz/
iOq6qX+ReFo2WEGFO2D2KWEjQ2/s/MOeKnOKzaItiIaEScQTvklIQwig8/ZzSy1n
z89aCtRbSGCrRwqwuz+hulyiDv5vquljeQHgn9D3lFcg3aPooGJ1+U4pmTPa7DqO
KCOkvBPm3rZt6hbP4ksKzFkTtMboBN8KewCxngGOZky+TBBOosXYHCdfhIjixdol
HMn9R0R4ZcCHKy2/3U/Rc1cap4qskdD1UGTgmbzQcFox2Pk/LBYzN0hj2BEYOsih
vb3tz25sftK8A0dnGRBXt8lJLDuvFxb3lgUs/gWX/7aWcL6citLEL/CpAbwMeOTE
43mCC+TrIWtDm16BCYU9zYNLetp7+NyuTDxnRASbRPfrHKm34XNfcp4Boi1e0TWi
3drG8IFJYqEQBZDkco/vVcnJxS59PUt2imyRsQHTmIPqqEt4Jd7Z8HPEhpr59c8n
ULvqJfq7FR5WtsjSvoWQfVjhnWmotlqZRebKEHr7yuKb7gCXt9i0csd+uMbqhpEp
AWetKqGF9Zn4fFM6VZxJ39cEpuQjuYAPfR/hhDRs0sRXnm/M733X8IprbAEc7UCC
O+2DAdrVJYKMwGEWRHilUpfxCpqmWVvvdhD+a3Nfpdy8ieXc6ReICCbmkk9ezk01
Sx/r2d6d1wNixG9y0lba4wC94rd/HLf3Ub5DazFGDcoK/eFBmk06CTnNd6JDqstU
QosJ2aEvil3F4HoqnE0JTymxPEYb+b9Uj4oh//rhfZW6PL24ETEecxEKCLCeZpYE
TpzIw/cUAhD2ylEJkoQaX2YlHsMcOm25PS2fyfobILIEIGYXwKIxkew28HN8xOhL
bcflhCW20PIDPtTzSa3AkEVLDQya/xpWsHqjYH/3RjgX0r6wEFjScpeZj+IJF8do
cuYF1wWyd20CjIsk4xwNZeUGhIXmX7K3vlxA43SdUI1twrArxKDKT+kZcCPm/087
OISTTWUbBsYUzken6DGW+jnsdEmuG5FDjxZI+UJFeAabXiPDgS2FJ+BhRfbHnSGf
b1BSPoRVnxKGl+F6n6lXObdE0abm/jtzWxnwR+6uB2IDHxOxzYX2tQ09q0WkbiQv
rmYGq6muG2i2LahMRuIRjgsBQJeMFojiGu7Pd8wrjklxHXIE11ZY+lyL4xe38enm
unKj7UUo0kgx0lsSFZio1MEVt1gB6tZ0SBCxuoq+nfaB99jUNz9n9SmJ4laxG4Xb
Mg7h9cj6Uuyf67lpcbpPHcDylGzs5okpLcp/+YONXg7WOVJT0zkeaUZcSDDnAZ7p
vEuKC/7tS4gUfmYv5eCOz5qIRX5KHWAqadotha/6SdaZFQdaa4/6LmGuZ6wyFkZz
f/HPvGb9ZPFP6F9ix9jqGYTGDjwrD/DiGnIpeWtkA/uMruNc0f7+KHK20fUt/NHv
rHOTzpheKXff4BmZWorg3PX/J1439pMJDREHqSwcK6bXzcnDH0K8SDH6CjiUslfx
ek6QC7EGl4lwHisfHF1BMTvaWptAn1TD1q0MdHOOIf71X7MTz/qvERJDxvRjBZli
w1qFsu/Zv1kxV7I3U0i0F/HYQefcUyhNh6rDSZHu864yfmEMdke0h1dubBEf7bRH
BN2/60pQSF8NaSOaytTkS/t652k+CQBnAwJaMfLwkY7CJEepuE2HIZeeu0w5T5BX
HHeFO9QaoMIbfQxZ3lBYbIW05JVfZPkRHKHOi/n1A3/aIt/eXPW9PBDy1sEQyG4P
3B346mWetC2DncTnWAVnJfyttJv5xZU22zrBNk/GzmE4J+x9gMN/CNQWGjNVxNSC
tOd+npUEoC8K2gjFikd6B1G6MbDlcdkG70VHna5OJ579L7jY49CGsLzMTD6gq0Of
9vgc1tdfPBZ0aTBpL//xjVVMn7Lq77puZXCse4Md3tM/F4gNCe/o99gnbMfLiO/t
0DOCVfbBQD+t6AEhnkxH5sKS7J89PuQBEvD+xj8lHTwkLao0iByn4yGezlVk4t0P
5ejkFn19kidcFp3E9jgw6O0jC7jOhQ4Ff85PCFdgQAS5sC37BDFNkdwN64kcUdh0
QoWDbV+RjU/SnZD3UaPgmzGGQnnNXqtPfk3K7e5NFWRA1Vw9ZWj2+4YPlnGz0pZP
G+GonX8pv2IYovtg3f/rVQtTYMerQY/vEQopoWcxmEr/jYtgqo4GiKYnUt4jt3v7
cPARF1AKJlnjlpCPulu0B+Tr+neSqfjkdFNIWtBcQdhKo5Nx54M4VU7Mh7hnbE56
b2eIt9TBtrLi4bmINKFkN1dkB9PW0Nl1BdD1ozcCn6GHcDGedEOkAAoQ0YjsJXqD
yJ/TKiOQ/c1btMGq6noJHSkPX/RD+DrH66Gjvlg8498MezVy+/P5kCcxegQkuqLE
EYqQbftd7KTmH1UMmCka2IgerEBRUOj2fhkPJ/X1nS1yNnocXKe8m/YC0srSGFUa
iL1CH0ry/23UfdRqOH8Sk1tIWlnMQEfd6CI4EaliKSep1R7t23RhR9eKM7TjNEXL
70bpZYsa5IXxJlkrYsgvB8TiSJnIiCyoQuDvLpW2YFCQTFHYoVSgPgqy12oYx+WN
EV41DACFn/ze8fWvcC6Wt9QMvO23+IbTTVBEkEII3d5AD1frIpBqsdXm2NemdPO6
VH5X5W8hq0EtcnbC0CN/IraoqhGh9nGayOcIhSP07LsrU5kg4y7WLofsZRBE18ZX
9lDy4SWzpwTAUDSJgNM3nRMVFEVja4KwS4skIjlAX4GeIRBCkWFNEG16hl0fCveo
MgGwTJTtncf1WI3M7AypjNRcBayezSMQ/Mp7HJqttGmJLiS11No9XtHBu3yg2jnG
a2CB+dAukmk/J9kmgsGdA4ma7k7TRxOo3xoirmCupWE0hK/LXdHsBQ9x+vTPM/Tc
o+P9lnDv0dihm3PGu+P09n5bhh59g1SUwj+hsvu1fPaF4VclHu1rruOEulkiR8l9
dNMtkJrV0bH4UcGtXeeoNwJoMqt2G2oRbO4qM/d8p7NL90dZRlrkfk3CQV5lEGgS
PPksu7rHhrliIHuozyYK20hAppVkJ0IOOaXnO79ofmFd1BYmBIZkcXx1Rkx8MhBG
mR+tjx/TcTq+bj8uLINKMbnBLPm+HF3kC0hs0RWLoom/TMofG9IMsl3Ji/4t3jgf
sm/EBlnVR4IW+GyhNymgu45nOZC2neJmpZohPTaOrq2FoWTx+0adHmdHamLeN+oy
qCLhNpV9JVMbjGzzMCl5P0Vlh7MOe0BZyW5tAGZJK1tcog9I9ozclrygTBKaz9ed
pxi3ZwCAFvyLOfqNHbML/Tnj9md4UD/dCpN8okqNgtOJo2gsbfRf2aNpUnoQdEYU
e5rIWWWp/OJz2anWNmanmqib3uZcHQvnC26BW68UwCC9rJRPXmM+Mp5MVVWMYgtY
LQdDJqPmS2/ElVri6NgqKeWPd8f7xgN61qSwNhav/XP8Kaioat33LfK8fykxAAg7
Xe333YH/K2opAW+tozqbtS210ezQwN2KqYYntRkpAGnBs6n7/7k+Njm2MsCSv+bC
B7DZaV79tcqM2lyrjc9LDQZBKGrbxQjoAgFwgzECRL7m1TKZzeo493nslg1ml++s
2n1XobLCjHEvF6ECBxauq0C025Lj2CAEU557/3f6ei4HsAi+P+VpJ+HfrLK1I/uU
fP5eQ5yOv73TjjjjP7mBLxmGEsH/2nKDiR4ktDGhKExH4p3UqcDDXaNSJrnZ4lci
6Bhau54qmB130nFhWokbNVm05oqQKHuLOJPTT501lGux/PGXNHin7uAid1uwR0OJ
YkE5s1mTF3lRTCM55jeo11d/qvqlpLA2jwOBlfHu+44JRN1N74739uhVvP5Xn2jV
2PENmO3u1WB/ccWJFRJlkqsvM/B2e9gV791m70dCUIWLmhkkFtlTuqty0qNxwbOW
e753ktwrV08qpXFtUM1n59Hv69EeWfCmW1xg+hLZkY/bZC4As/HIxRct2Fy8yrn+
w8H7nfujQMYHHkcoyzCC/oBsHCdz8YcHKJfX6oNlHaAZtzU6+B22DqnG+jHPxpwa
QjKWuCLx4XWCIZprbBDUYeWFf0QFuTGqqTGwentN9K5C7acbDu2BveBu9TR6NQBr
otJpEHsrJkhEwRxKkYIschk26ysp2tDD+3pqCGnt21mhEb0R9UQK2PNvMyPXEX7z
HlNy8TsQ/qqzOYDFTOklkVRo7YgqdOVpTsvoScZNk68ixTrgr2Osc9AossAGnUMj
3+34s6O6mKjaUeEgomtL91QIWuu7ifMwiYQ6g53WeMe5TuLVakoho/cVz27ANEkb
tVMBw45DWD8Iki/rKVdgQYlS81uIVMqqKhhCoQe7QNe2nCBiuLT+0SiX59cgNM68
1h297oOL3CJOkTJCKVCD88qjCi8NDAoT7VVdnM+S4N0L8AR1grYJzCDmXeTOfP/d
ntD7LYCHVKlu6/vap9ciVchJdQev3GEafW1pUApnaGv5G2fsnS5Y+TzF7tCcr9b7
5463dNPQVH6xS/X4ijp8mieBp5CQHe5yjTyTt3YnfIXaYxgsnwFLRkom/jp0UzhD
wbCL0sn3x6qhMntYeNcr30/RKTJ0dtoTiecKvQEvw9+jYZE4TWLHu/CHWfil55xS
wJSkOyR/UMm5ceZ46MznQQ3b7nsuYbwpE/gKzfFUtWDikZ7kLhjs5ZAiro3lyrdp
IIKLnHnq5o/SK2WBYrHF02zrcpWb7IZZsEKy5N1Mp/v0iPbna6b8FZcdWE+xSmQX
RNs7J+9an8G82zldtllRS59TcTx2saE2E1U6VXq+k5fi8mDiVBba9yWOY7Pg7daU
40aGzbq7w/lD8zat0Xvlkd8l9sU2ucnEMNEGbDEWhc/cjy+ayX27JJtvZyB4sK8x
wr5iZ9pX4qwwi5AvCXewi1LYRNthEpX8P0iLCk/BGxxFHNFwE1HThR85jyFY7fbm
8ocgKH7pi1z0mtKhppDRZXAYXRi9QnbfKQ9CGHgjr/k2w8fP05B5mMFhJHzId6Bv
5MuwgbaTpw7GQ3ab8zpOB434dt4Eownk0qY0+kzhvNubEY86+i34Tb3mIWUwi/np
O+JV8mmwjno0Dx3z+P6V9iR6tAp4kZYbPrqJcs2M4q5XvFLGBxrpniWUnErrHO+c
tpHUnY7P9DwwBgfkUK1C/MJ7xtp1M9PttuZpNS8/GmqNeo9Tui+zIuVxYVWgNBPb
zuR3u6hUh8YiQQ/0g5ohsR0RmRg+hRovDEFPX2B7Nln9sz34t3FCb3vWti8QlBv8
w4fXzgPVZ7BCCby0ozqLiqnZeR2nacvz1jJYHbFJKYYMonto732EUb7Am+1Lka6X
bjg104/osD6aWHm0wXvp8y6KVXwE65Wmd+jfy4vYDsxfO2Se42z1qbpvQDgrfOvb
t9zb0niE0dBAUZgGuMNMLGIYXCli5mm3p+8EK2iojiq0W8VfvhsJda7FLbcjE8T0
imEEmusJmjWkyen5+YDTJvQ73N1HisGDMma+GmXVWU1Q65pJvZEnwIng7cdBgd8Y
w+05iw5UqpUALAsS9qvSyD2wSfe8q1OApeXa5kaP0gRSccFTvHokgWUKtmp5mabr
+A53qY+UTYOa1Xe0OrntobLKs0KP8XtkIRDPB41fKxY43eKXq4VSAtr6lr6k0bnc
U00ez4GU3b5mpwK+1JD6KIv/xDCD4pkJGqFNfcjxWAnScGow+6x+E/NaeJ6ZZz1z
zgTqO+ye4Dka+CjuDNrNGasLpjfTBrLYnsQAJd9HpCMzqZ34FY2/g6UTyu3YYkKn
F7AxHExPHJ6o4ir2y8+mH4bcsF9eTIK50WkNmCVq5fYOV/lRrbaRgdpm0uA1k89x
lgoBPPBEueyC569uvm5pUb7dQUDjuU/o9UpFzaTyuNoTzEnR2OhetPcI//j+a0E3
C663ml1H6Ke+DO1Kc2rGuEI/EJBif/PKeI2lRZZ/BfhnFDl5tA+rMRi52GrraQhk
R8Zspz2ZHTZAnNaStPDTyI6lVNLRVsCKCAQXewlRBqbU0rRTH88ync275WT40WTf
trjxRcFm6hYYakGFprZHRZ7n3AO5ngdfYaqtG6XZvz28UR46/rOvrOgcywJKNV5Q
ol6dSDYzd29pMQF0R88e1njJhHhqVEkEo4/s4I069a9pFZczmv6K6abq9qMqDKtW
no977WvuKEqShsxPrwKkifyRyNx0jV3RAK8gJFGAf5A/ULkS6ZliONNp6H36a/h0
b16be0qYIQnpIFZn3azxqYiPROhHCgJkVDU/0nlSeYENijiw5b/+tXBnc7NyUUEZ
PRae/5NDMEfB7sf6rZ4cLUr0TrFeAT2Gz5H6LqiiQEExLNOjIY0L526A9EbgNCbU
txmAHwlCjqPHFLISbl3CvBBE4nddCR0uv4mXd79/VVbhXkbVKzwGpjBFO2H8NEtp
1zhK2V+3gep849afM93R1oODG9ud8yMGHpKl1RzB6/H3bXxxCFxJ5HmExyYhIpH0
gEwpFGAg1NEtBReDj+FBXX1i8wjL7LIu8QQKKu3zfJGslrWdgiFlpxukTlwPTpIk
2dnFj2YtrmYGbGYgdUBnE+a8dF/4ipYKyjWWRhxrHmMI3FdjklNRPXkMRleiygE2
FWfq466nycaj79io6R1D1adE/wmWadekOQkSPZ4hmGxWGC5v07lpXzh5A4pZS6F0
T9vEjLSpYTf3hNZZxZr4pDCRpASvoCNC8S7Zvks2v25wqol9G2HD73JJT1ilgmCg
Yq1TuA+t+9Fli/LxM/915OLlA3ieYG1GKY99h6u7Xm5rVV7Sr4riHmidrLvbLm44
2UTxPK4U5Z7+fxQXB8eOPDwWzdCmcK9xFhX0VLUXnZeMdDE7EwQqlCTGzhGPBoxx
xvPWKn5+gl6qK/fs8AzfoQDzjdTO4aBvY+b+9Nw0XLtWQGlthn6MyXzw2g6a5qSI
RZMjoHdNKphPobhM+CUPxjLBs214yzBINvzsklT/vM6GSzrgkzJ/oOC7Cg6OK7si
BElV1uwsc9IDQXhheg9PVB+AsFfQiBSA8P6GUKLHPmZjWSvfmfLcC6XvVSR6k8sB
yINY+6kPnkOQ0L9BpGZXFVy7VGlFSfcfh7Sbb2voN382I15Nnu8esBHjn+74zoA3
WYO5UDocSembnIyVEXVAxjkahrPwi+nUfDaEFX7cE3z6yy/tDVMMqVXwPFjU4sq3
E4PJV/JkPS3oLNOsF6CL0fn9S1BXH543hEXI1Se0jwYzDNpd4537tcKkqAXxJWOu
vKB6gmec03Ycr5SoqhkrtY8rCWAyDfGFBjwYTpw4nXsec1eIOJDgxqZRgZu31AFd
VvXlDwwN0pktfIfriPF+ExgbvKKCa+BOIYDY3Rd7WY6DlQAoDwOL2mlp2m0AOPcK
0g5KN1QDp+5OOpxzPQcAlyLH0cX949Mjgt+JqO1kEwCEpU6OrbMgkuuy0LJWvd/9
uZGC6tWm/4iThBWBfxGgWtVxFFeCjz9D5Sqj9L5yLqItqOa4kqDEV5aCjacfHZxf
mchUbW/kwlO4EpLJ1oX4k9ifX0MzXNgWi5djqhH/XeFHj+rv7VW072Xk8ionommh
UuS5MmA9ZSaPiC7qbxtRfOLBSG7EAIt0M8j80E6OPtIC45bioE4QXR/mW1EZ4dJq
dE3UZ3xTrUHnq7N7chC8PGgJmfktHrD18sf+FbYmaSGCfGENv4niIu+eu4LdIIs4
QTIVH6ayj2A2K8+uBI9Eab9YgkmihTX6RATFP6mpcXtJhjbk0142tl4VJBS84tj2
iWLs1bVm9Y8g2kHMfQOY1gTq+uSm0iE/elQRw6jaltRZOibkCRKVS8Sqbi2YHsCa
0URDY3F/eMRgKrcfoCe4abQ9P4arI0QnPcX8/tptXd81KUp29tuWZdPtfFyPNcml
jXMTODAKSreJ3lHVB2iraPYpqTRJx2QsqB3yKI5eN4hOmbM9ulwhZeUkUloVS4W+
N8Bq3bja+BsC6/5vG7XAFQgGMGex71eJ5rLR+cXRvE749xbh+MecXQXwNus2rIIz
X+bbfkCBnAzzy1xgZqwgw5Ofx0tQflsFCaZVnulk1wCGmj2U+pz7uXqVCLCPjE+N
SDCfos1dSlUL/aMFWCWS3WlRQeEPGrlS+fMWoklD6Yq7lMNlMISvAhdvA2iAK21l
00SKlsBPqorn5WsO1HAl4IiWmh3ci/ql8fMMsw1UnjAkrRYfjt9aJVFjG/7sua46
tnTtrjwBr9x7b1HjKw1dmT0PpXToRX266s8jTRzlDzP8z5BV31ISUGwqVzPsoaGg
yG5EZz8MjaQWV2FT54u06/vpcEnub+9961YNQ2OepdGWL5wAEqyVhdFXumHhg635
/+tv4wFRcDn/DYFXci69hCdcGg/vrNzYcuiYKep1TVHp6ynDvvbmigoDRJA4xeSn
zj2Se9Y5vsD0ctbrziyPstpANlS2Rq6icyhHD75PZ/KI3cOucI78e6FTQ+6TsCNi
cQPaOGa1OUhZ4ka1ImW2QzhTsnlFhqeamLYLawNTLwQ4yeo63huwY4fsmj7bbFnV
jWbZ2qi84n2i9qN+fu9bCUmeL8t3PLXflKxJf8cHSPpiRHgBKk6Qtj+CfmRwom9V
1YBnlAumQUFdmFLwl6+4sxQP/ed+4UC0taAfLT+Lx39+qW1w02Ev/GGubSH4LMGY
imiHG6aQY+cf5iL/nmpIrMsZ9jHROKmXS71YU10FSgAuwq0PnB+Xog4cVNmscIYo
sRHZX54DFWqtq7ujp3/vQQdUTtA9/9iXHkcfgqYEM93FOym3b7ZRrcI1OMBEL3r0
RLxvmeWv1cg5/k5rePweTseABpTJ9JAiGQ/sU26+o8DKoVxC7r+NwwSLOKEf6RNy
I0+PQrnIrWsqp4t293+v7kYJD5MuJ72b0u6akvRKB5K+rFIf4Uo/6+NaynhMF25J
yutuxbSnjxYCF+HPxhMTsulY3oqxBgSjIva2q/nKvRY+V4IUiPn7zkLju7QqvAZd
CWSZs3Y85WZFQTUhbhq/Gn7ke6KHG3ItOnIl1ncB+IQ8+hQccKlA/nVWjjmYvk+e
4ZK+gzCRdwPoBoxic61f6RGRhBj2yz3jIAOwAueOPmVXHfAvLveddLVPqkcx+9jk
fPGDRypq49omAxQOlpVWNtCr5+WuLWn2MKGS9oKy+vGfNTMUBh/DW3Ywp+GigKsx
JrwH3p1kDtC9y4cGbA+JoBT5G8cbWcoRwbrOUR8VSTRvazFu7IIsbPgWVDzF618g
rbeTHi/9RfJ60pguqZXi1HrC+v6cXwfEwYpdhnVylZMlCehiGnC5f1WCJzesIRP1
cGGd/sguSFVp6NyaUDiiXzGiPBhV3vBz6F6aYXARnSGzNiXUaMMCgFVtYXTtBSlj
XBW295UmoJwjVDszbpA6BVnx3HHEQlBU8jqUNX6newbu/DLQLBrl1UAF61b5DR36
DbfZF0tiyB5ZvdkdX2dGuNBtKtYNY1g1uJuRXeorLhFZlmxdcxsQCsGxc8v8VUBZ
Y16PxlEvwMAbWJ+ExF8u3HCjYbfhoJFRv9wc9UKU1iwQy5Ig2Fb/xsrVsS1WzKsR
YNuBB64cO5NscEJxH59FE7/wa/Y4iSx7S8BdH37+vURqlLsJhj8KKG757Te1tD39
rAzDxsjaaDNN9ZlsojOHSVwXlV/stolbtpNBnY69MwUE1rgBAhgxdfE2lVMbNVu6
K/2jm5zLOzcCzi/AVNWG27I8iSOa1kJBGAS83x/4dcYXuAHJNQ0b7Sp5x3b1c+P0
6B/hoL3qHVyMrzjhXN1Gu8pCGpxnYoRpVbt9Au2fpa00QgRN6VILkT0O8w7n2qFJ
DNnhw6+OFHc/fkRdUDWZW2NXyP4n9Fx3suev7Z69zuhhOGLiBpGazd/LvhPpapqQ
oX9f4YccWjfzs7mBJm5aKqwArB0Wuh3HJ7upE2OUSH/Um8lJd9A3MTED6rdfw1it
BAUs3XgVQfpgcO1gkjv/QbsKTaFGRJd5fU77VYl60g9FOk9IEJsv69iei83y0XuT
srtK83pXyur4Fiee208fepF2XOZOkAi7YrgFsvcCZSzr2LIvXJntW2Iiba/1yGXI
EhmsNiBUyLLDqwpFuQYx32IkRVFXTFMrTWmqX8n2LdP2zAE951iddGGw7d03jvv/
xazXDyBcYEDfp6UBH4FEvcNBMp/6pdGy5K6HX5N3DZfkfmdrZYs4kba9bh44A3f3
FU1Y0Wca94fACEy1LetYLNmc8Z2jU3/fEGNWVhE4kEwpwtzMFbbBoAZWj2kEeU4K
iU37f9OV0LMacfM+i89FUafVUlih3Jhyx4X4LsOQ6RPdmOv00vP+9BnDzVJfMZMG
efEItJnc2+K0QqZWVS60Mq0r18o2ny1NnWVI3mWNlL1DCrNlpOE6Xk8GxWQkuikM
f7rlSAklNbXeApK3eMgpJFHXpqrCXLlNrqjFmRB4UFE6yDtHsokCR5BtAdPKj6b6
GXDclHehUrriissQDbvPXpxfE2lnRRJRwcc+lEoZ66Eyxr/jNMW5EKdQCbHCND7V
s1e7zcTQypz479KFUsnIXvPslFYXbdo9mmfSiQv/xLv7lO9qvsEB6ef+yY/yMWQJ
cq37GHOzrP2YYBVejtuXjxOh/JGTTSSPNxthJFw6he4Bpa5E2w744coTkshkclSX
qp47KjgJ/XAQuwhDGHuPjUYkuR+ohFjEkRxtEI0pJFsrnbqaMbjappjxcTw4h+yt
YqGDfvX+2WGOy1tOy/3IrhIfDF1ltHQ5TyVVHzfXWbq4iwbb8tMyzrePeIKgWNiA
n1YpWTeV4abbb3evnXvshz9o221eAgnrg5kb2dUnEKO9RJfgqs/fDZaDIMJHM9Ey
JJP2P+hYKodq4nrqM+9QkhqPc0bE8WyFImj/w/dgf2dXsfGbaqmBB1kt+/KHP5Zn
nYdLyWhTPn0Cd9m+sinGw+VH1FCyLIoHfQDVPIUIRV22nn3P7jRONIINLdmJvH6i
fOMKZU98p/96a2UUMPG6GrPVBwqEGMrzHgYTr+dITO0KQl8tkYQ/uP3pO4slfXMu
JCe8P5eMipB72H9+u0ppVgLHapIbcF6/TsFgMXzoqT1jumOpXH0cH5I/X0aLyCdR
wKCs/o8Gryidc5RJWhhmreGF/u9qjUDZlB0XOsUehrwWXS7LjDx/8otyBNKVEfio
aCm5n5B6/kSfa8j1DlyDcrqQ0kBlhkcJep/Iu6r3Ut2JkbA5semmoBrbajerOaJK
WzZDzc5NQ0i9QEowH25NhXydRA3tLi/GblRsWtxb6wWkzG97I2QWDOqJsuzfroAP
XPL5Lzzki7Jn8O1gZeojGxLXmG42kShH+zB46WIsY1fZjdtbaWdb4vc+2jvsAabw
KXawG+Lrf4Vj4Pj+oJS06zAEEjXsfeK3UqEenUElBd7CM4dbscm+Iizq+Z0buH/Y
J/hOG/j2Csh2ntRPhhL6r7PsBlUSOS+E6CP1CsfzDYX9nBy2lkkcmftWkv7lbOaG
1wtCotTM+rNdJfGy9WS977PFidDS/neDqFMT3IdevhnRieX0BDPoORWiTF9KChS7
Do06Cl3pqP15P8R5z/U1ztowKr1xbkoJom/j+xd2T5msyY4mr0m28IDlSRo/ASW9
2ajqPJs3EJHJ6qkjZ8SRiZkt5Fl7LJGpfYY4TRk68yZKCxTDcqYhVEiR2Z/83Bpy
4qv3m04TBfd+y34VTEceFirOUvO4XYSIfShVbYQisQgKS2iSB/mdgyBXm+2ZMszk
s7w5zZlBtsWqHDSAd5ePb2/CVYvbX+1oZCy9Y2HGCcHll0gOtxUBcG32U0N0N7BX
LPaG9pbqQq570olt1mojROkesXnYfopgAs8OENZW4aXlAWtMVdGzOP8T6yg5p53+
UEF49ySylRcSi2n61K5521w52W2cC33kGcgnLCSCveGtlTBvP9IGd0XACRgTTsm7
gzDprHEeohcejikPgd6xzghATHOTxsDuKtDEi2Pqjyh3c+BdR4Xjq69lGFE+l+bi
oZm++HJF2ou0ZiPFagRdIM6p0qrljxGunhYk1xW7OG1EOVl7cNz2WjVvpmM4TOqO
5pXWTNbpfKWMmShUwHxB+mPL//3zJjodGOXDH8DnEV+gaSVSbaDC4w4K/MmYLXUs
xDu101P3Mmg8FvYU8BIS2b7xa439tHRLZK/KiLdkchMCmmF3Cc6p8VUT9hJRH7Pe
/FMhWcGePU2juf8WndGAgWg4Ksiyl6eSqqzeAnLHYN7ej1BLFc8OBnyeEtg3p738
XqRWc49axG2Gasr3N+RSIGVKySROlhDpbRopW6HdeuNJfJLO36a6QJYjfEEki4CA
JAyN6CaNuoOBnWeq0VDmFAriKve7PB1MGxyX0yTuR1On5MVYBdyu7rL3XXNTsW56
b5EYE2nmLAAoghSp21GBMFQjDqZLJ3K+r4noDGPlK7TzlUehsXsxh6Ql/memfuf7
XgJwY6QM03PHHfTOFzAG4y2tRI9WllfZ9s1WBGF37QWTs7aaaGGoqmWIz+L60DkE
Gh9vbUzmEObr/ejzZV0Ch13+AzuvKIQ16BFkwRTI7Jo8c9P8N5bpwNPIQeBfk07v
OhzYjEpZwoD///rEVQhQcLuGI9BSIluBxtrlAWa3w8X4sPDSXyy8Z9NEXMkfgq1I
equ4gPnox0wGNrfhlW1n6RK0RMKWf/STTEx0d6X6FtQ8aut2p6vUWUm7U/yCTdmL
Ypi5qLf4pvZcsdBErYts1UkG43/JAv4ej4+mj5Mf10J8ZtjhRr6mJoxXqS8p+P1P
KAbRisO634my01KVwzZ1I7w3Q0ixX9pMBSc2m/4X+Ulez8nhO05XEesLDeGKyFh5
wwrta/Jy4HzIHKnNfgLCQYIj1/YZ8It7bZMEVC4GpbX0Ivm/u6a4itJGWAavm5x4
tThzSIfoYv8rUBvJFbpJfHv3qq1uxmpuqPKsu+hvuSuBqa/SHGMUVVWCgH6iQxuq
5Wsz+OaVG0JJZR8oLf9GZS/6bqHc4zsLIddiBfyaHte20MMBlM86ehjy44UCt/Kp
NW2xA/ETH8ynivvAkKgOIHdW3HxO89C8LMjRVsOzKfOL1yNvdOyVhuJZlCOp0grs
iPaHNElzghC945Ozl55RsvYp+Rn0v+ek9t7uPkMar6Mlp0/HHwpFxGhhmJJQxz5e
71QBaIbNdd/J1bvxorzRtuMag+26+QQnx4s0a+Qgukjz9mdaYAIUvTCPPc6TStXp
pmGxhR3vB6zii/wwN4CGwGL1nwl581Z/E8GYF2UfFfJU3biUqZPPwGaENYNNJAra
Yvc0fM8JOdiMCcAht+LVcN3PXEShjPKTtEEM2KSZFyFgRWiIFUmTu2vIitlb7vQO
FNpoBH+pGZOaRNzGGvy+2CvgYP0RaROnj4xbhdFKbF74bCDmA25OcDV87bytj4VD
yUSlqaQCd6zRaeWXmVxWhRDotGa6Bs2aK1X9WZaLvW+uYY1ZzEfGmCo8+tOewIfC
3wYNOgscIk/X9l17duF1q5v/i2d681PJpW86gnFYoM+3GYChkbMD9/XfhOJ0+Gpp
JDJwVGxL5c2OljCQPtC5JrE1d0X0uxOq87ALzbALn5OdMXNruTHKtY8HDA8EQuPJ
vyQByayKBPeI2soaRYD4TdNzXSbF1KaYzrsUR3LPFswJTxbxTEeP/YBWhswX64Xc
UZIRc8ptmFny9E28tHnmVP2y9UD4ws9/0dLKHz0mM+TTu6QlYxkjbGxm5+GDtmzs
sBA3e5emZs9ERrvctXsQFxEILNAW6BI2eynWYpUJx95gNMDBYnCoqKj9e7IqyQb6
snrr4Z2lk+F+9nJg5+WlKQCuMeHVg0z6XBG/sxwPhxqWEH53rYVpmGge4pT7ZwLv
HkdpIYF2qpm9siBc+CG2BzCfdzm6vtuyB5LRpPsA4lfqOCvhfjUzNq43Wu9xAeYL
QDKQiWNoNXUJ+5O1B0ICPKuHyMq9MIfV2TfcCLbQbtpPZp6rjvjRg8jFtZxfq/L8
TlN+Xvt4UVKMspqDM1wHc6zEFg2peStGYF9VsoWG7pqyfMkf5FsRgA76oO/VylMB
QAJetyejDQa99n7n2NncM98yZEXsJaElbhBPH5vcsc6/1qxIKbJMiYuWWpGD99Qa
iPOi4/wA8T+43Jw3Gy0NX4c948pSulo7wLqBH0dWpIAcgJ7OV60sXxxtirPyx8uA
iMMzbv8wWYCHG7u1Oa4VyPJiBZjPyjw9WD4msxGbPJ+wQBxOyccx0maGFz6R1Krc
oqYqCk8lV9mgjIlLz0Xgb0tF8ejNaMNtXwck58FuaJVX20SCCpJuPGJJATm0q2MS
yGE4QzHhTUKDPjy+t1387gMqAhPWh6WyzBMBbkZntqPq2S5fhW/yMjhIQYSh+1qU
Tkm8t9sMq4JLrMfvN3N+QZ9XlZa8r/79lH5PddDCvKO3Gx8GN3x4nJkp81GRAfqP
b4CI3r3qiMMpJElgepPiDc4Tjkkk3aFjsKHwkCFylmIpDwBDRr70sH+GUnQz4cPX
B9tJoKr4Jo1jPTi2GGD5HYXUe4Nkpv2VloRVpkv43tBMQFi0O6MuI/id5vqLH+Rx
urXM/oeaOxy+o5tGaSImwVMylHbQaTpTCQ/YRyWsb2MwOyNUGRMLv6HBXHmmOaAg
FSd2hq3dQN+0LMRm4xlqYqMehhIDZI0Ae5GvVD1HKk7xomq+htM/UgFwbgAE/GdK
JZksLHpDod2HxBrQ0z8IdHUhCeeb0OJPYiZtBSkWu42ailulJAfyfj2yapLwDowg
cF7Dbwidwf9d4wmcc+he3k3HQ6sVY2zmjP8crHsSZwMejHEWWnDn+xnJzwveJpkk
2N+IK5X/sdWJ19GxvK3/Noghs9TyTMxpALxRT8s8aGLBwnsQ+uhyhpLz9Gm/wL26
xRpRsePOME2l61gU3dyXoe31SYMRutF2FMGoiXelOJYCfg+5OrX0Ja5qagIgdEfl
9j8OKMqBGflGCkhzZPW8MfruI4MDkvHsApOFc9Iwcl+ttpBI4917r9xVUPLvyzpV
U3uWTpu9fdisStxKEWEb4HWxQcMX7r1MnMCIdbsXvm6zAcMqPg7gUyLtKP1mrsZB
twLPDwD7FSNjZ9Do52lblHEA3KttcAUG1b0UbKhhku7+T0VKHFXH3S57mAFGBGaw
xdgdfVsN4c+oFAB2ub4GT/gO4HV06XBaCgpIuKAQ9dfjrK2R+z4JTplZoesoZNjt
IaPeBk9yTN6cs7fBoZllS44WE5J5m1h+mVYnLgsrP9zjKKutMPNohZ63xuleUiO7
knzKJKmC/DQfnyj6o8RwUtvYlgALfFe/Gky9qbnLj2BDb8x3l5sXWlzjI58JPivU
5FyUfocwmEwq/OfisgdOTU+O0gDl1770R+H9dxC5hOQaawBhFbe/UnsgGgbcK8UV
U2C46hyqHvsbw0+paySENAc3MSIPPvK8s3LXw7RgRDaNj4J1apEYVXIdmwpUNDW2
NuS0fwDvlPU236UEew/MgF6Zmu1x0B4p57HV+SkQrog8lyyPCciWY4/WRd7ZTtxR
XyLSuS3k7tXgHMq5FevjJsjmynBAoSrp0tcW5rsotFNaedbPyj6Swyc3yKnztrHD
nMe8xui3VbOvM/LQqCQ+xARvMQGt6H4+NVcDqHxxwDku7dVWfP1G9Txw4kdfWnDD
jzwKWdG58e/+Tn+Py8EXx5a+4EJiZNwBCjJ7/PsVUormtZpugAPVE+plpm4Wkl21
Xu6QcsA1lkdBkwgPb/Z09WeMyikS5Cu9LADHjCfTM5Yy1tCsruDOz8FWak+lR4wS
tEqGnHm0MG/mHQNMQUq2BJbiUrsnPGAvodvy8WOC+26H0PVdLOPJuAH2q+cn8TAu
meeWCgXvQAJQkuz64U9gZH0fpj6uTYw6Ox4f1+mV+R7c7QCchbYJZgPo93tNJw7x
casAzT5/jUHgk3Y9A8Nv8/1ohE88fNx8HuVyXSXdoCCaHl69CgCoM6wVOYoUf0+t
dZE5xe2itEx/Q4/LvBJVMI0YnhSNSmoMOzRGj51c1rghlpnRYJ+f6BkVxK0WyFQD
uBKm2EdVy91NRww2h7m7vUWmkqeFBaARe88kUx9ZCqajY5cVbkAPZa2PqPybzXdA
7Y+sUzDkYcJC/tEvNrhwrVSSORkWLscDcumJCPRtqougvwR4BYt4n4uqnk18Jriv
PFuRaZZoZUJ69Y+twEZT9+SKmjKpsTm7Kp2KgCx6e5bmEEFVdl0tWXYqZfLrLdoz
lpsY5NQykprpP7md/SvEgZJr4oUwOuXfWcJw3WtSMhPUfx9UzUAKhzy6mVmFaWTv
1qPYiE24V9RO14wJULSO4H1NyGcE7uYIwIX8lNTc8m1xbOX1b370VL9MRswU6Ojx
WQ5Ci4oO7rZVbdJ2EsGEiWEy26SCU7EMltqrH1KiO7+o1dCtr9GZyHvmdkx4Sw3z
8wHj5EioI5w2akNuGSmDoHlVetKZCHev6wKyZcCLNGyjGeFvNlzS91Yn4sZGnvlp
zInbZxQGzpKB6UiRpf9jPpFN/avZjT7rKBJ4fPMMUf4IwKWwrhuDYo3qrQpbbHcw
RVaN5v6iwrga8EE8T4PAMBNSECwe3noafKLIY8bgZHYXIIhrVHOadiGsrcHp+Gw5
rWcychipq1aweTTQYHeyBxvDV9erZJLyy5qfXCmBy2wkHDSr8m4RWeO1faPcJ3ZO
udfNGEAYy8WF8fe0ZntJm5+sMtv73lycS+Sd7wzmOeHdLcyQIM6CRVOMXZGrWlz8
kixwO7HdZiXURUzVNZe03udwm1wqk2hW5WhZz8aTUPaLXFfQZeDu1fM0KDV506ge
uquy1EAGDokAmA7VTIieB7t60hfJOHeVd6cPYW53C0xDBaEYIQG7Pf1NnhzVS8Gj
TunZitZs72ioHH0meOqLrzfYpjh5rezb1su9mxqP9vxPKhc8U7ebLe+FPre5e8XW
uoIK4jfNGO24skqaFtx2P5YtkjeBrTW8QDq4Ui3zEh9Ni1eU2elWFk5OAfzKFnsP
RwfsgRk5nB/QmlxIXE9Rms4LqQsE893AV8gOcCJkrzRlx1G2TSqH/O0Q3VwH20u/
hWFnxwML9oLJQZWeY1j8l0Unwrc5/760QqZKb/6QUO1e7I+cr3v2S2d2FafpQnQp
cPkt9sBrrM/Kgssfv/tdwgu1DoTqaQc+3kQyHEKHBKQLdXJmz3e44yg5b2KhNi0T
Ujjd1jA+cEZB/dMmhZf1vHIa91Y0CeP5ylwK+pzUN0aYWJQrMhvPBXGvni0ocvlZ
vlaZ4mDo/AEgySizDa58F5zKBc85/C22N48LSp2oL1arClb0yHTSP6QGmyAtuNd/
QXBkC8+CtXD3zngl9d2rbXcMOLos8rQ9iR35X3U+6QTDJMpslkxq+nD11r1dRr4H
TUjiuzIqN4NVh5M2wRQVPbypegkeaLbpLGzD3vVvSn5SSISTLeSuNe5JxS9kqGX9
xhPKplksYKxBsDUG8Je3pSYDu1/lORbQ3UNiL/KBY5f75q/kTWG/RVbUo4sjdEkA
TiLBj3W4UWub27KOz/5xxN5pvPP3UfmnnjOU3ayu2hxdTjNv9chxppFcwAEi5k3F
cRYCPfyyVWs6YVTZ8lNWV/E1VDwjXZcRNcYoRWQu731iRgSvJFGaTHA0SHQjxDPf
pUigsQqoRCLwyBfadVuaFFkgeP93WPoMEZ0s49t7nnrsgBWmXJcmJW8tgXsHJT+U
b6AaN7ClnnqwF0NS6iF3XDo7E0ZACTWGMC56f4sh45WpeyX3l67WPJnj5fUMEppN
uiuoA9kuspUZs1EDRm1ml4MVWPJW2LSDCAXbHW35AuzXlh4LnJ7h5/b1F5fm4N2s
97Kg7lS94Ac6PQfDJd9UrvSiDM06y6j8aaF0JnT0vR1FXgO94tnQK4TLejYpC/bh
7I+27uEznQ9naMWKmS9Ju67463tWfKzZMBgowlPVaE4uj8KpvFRS0EbeXJJClug0
Kakekesm3bSNoU38XMWbJfdu2DBIzizslNYWmg+nzZBDnODErJ/gvXKGuwVldmtQ
8wLillhMC0JAnu2HyYPtBVZ4Zhk5kX3gDSi2x+sa7NqdGHb6lUF66JuKKg8YCR3b
lZ7uFnJmhqfwg5uTBaZ8XW5riOt5vW6yKajYPEh3FRpPqcZ6Pqo3sPSbVtywm+9R
kByX07aGWPD/LupKgluWzv9SyBIdix3TxeQtpLekf/DdIDEB4EwAh943K6OaNRKE
beWAuMdJDexViImFwNrom95OEug4pCkdXrhUhqVDw6YeY92uIvoJwfnLL+n8mlye
2q/Y29hKwVDdAVkWBhawCLe55KBw1XKvG8W3vpiRA1sWX62YvZiqfjBlZ9Skm1My
Bss7Xnmvr0XIP9j7U/VwxWWtzhsjXUgj7kYtnW5MOQjudex7gg/c5m1ARTxe2U31
TtinF71mdWUkzP8GwFn7n5Uh+PEXNfmrGz+4iuQ8VvWjYiX4XLT9BdxKYNts00Xf
lhpwV0U3x8S8a1gx7Ot9rda71bOmTljKLNetAZsqActIi6+IX2Cj/X7WWVvaBa0o
buWmdLe7Vhk49N4yTwQZcd/45Twvrm4P+Tvpy28j5BauDKJCTT6ioWRtAmWj7zxq
9+ffllhd9UldLW+L6ErSo+DZ6d7GSJALX3jdYYpxPO/utxhtOGZgs1kvPsGNhLZk
qlVA9XM/lVGID9bjIM9arN8/B6zmnZtkl87ScHodw/y2IIAJQO7Xm737CZJVFsYR
z+RXdhEXFXYxjazt/HhUApkHf2biWAy1DyDQy3rzS7Gtp4m9x3tXEzDdxUywkZfb
79CQRDC0mIUFxVOPbToD1jNAzq/Lert3opyrx37QxpAPjoU0+VcMw+qfuveykjQb
Q+qK0uTfURyQA44uJGF0Buoin9Fo4rhGlMM3Qc2ShDv2ERqb3QJfXxQIs+CPMxW+
ZxxbmmzOH2qmY6PhnR+ovYkoqWvPLdn2ooSi7ZUr28NvOVTH0qaUHkuNpGu8j69V
7h0hvy0KnCUntaunbP+W6q0POKBdit4kMVWdFdxpE9vSvquQXlfWbExesawZqhKL
J3M7dRsoUrHT4vwqULLig1SV/ornXpnapoQB4O2WQPXBDnlGto/nUGGyvj4tjEPJ
RaZjRZcaBMPrZKFwZBlHPgiJCsGvoefjjpumuEJjZzNK439TOOUzlm5afuALAkpX
UHD70/WzV779SnNrAzEyXTykNkaI/y3Xd4dAr+Oe7dJKacQQj6M+Util7pTbadgR
5vgRRuNCWSU3USuIHOMqvLKtEmzYTb2Hk/4JO5mSdf2rEgNbb/uybU+eLft9LKH+
5bI6rNPFkJHWsYATGYENYLM3DVf1moFD/yk857FF7+OCM7jMFgVKdm0MJsFqETLP
iKzplRWaiUpP59CHOBYtqmdq1ROWU9D8wPz2BF7KCxRo9eY3kFqKxT5TWfx3hgCe
mJkfONEUFFcDzSAo7+UeCEXBXNquwiMCOegmNdODSuLkW4mY9l03+Qk03pUCkVgZ
UAP1lfqY/Meuh9nk4I/LZ4Q5BBxodAo5DGHkSMOctZcwDZd111ReS2IhLFeCBFzy
jeymOITXYAAZCmtqZOkpKnX2x3K1V0ECJeJgWkoW0gww1GH/laYvEYdwi8O9he7O
m/v/z1TyEpQWuF0RCdIXworyWIHevvy0LWNxBVlF0/pGTCWwA3cXDtqOsBV2BSTJ
jxC97c8Va5u/Lbe9bGBH0S8G7uisQmjzHY9zpTOsIQsGjn68u7INZIsulY8jGCSg
ONxRzOJ94y9I62Ws9oy2rnfMINkh1EVPLOoa8HhOImqc0fvCR32d/oPetZdVdXNE
Ooqi3k5PnYdMtLxrc+bGxpweW4E1MtwLx0vdh9W1Yy01dsX/tEYZYhF1x701j5T0
TwWcaXYpX+ADPMNfE1lDdFYxKpY8D+E/zDdR9PPufb0hljREom8ouXA86xlGBh6k
s2zijHwBEHNVq4P0Ifvq6QjbMdiwP29MHxfeisPEn8bJ1MmPtuavfNpfxBfv2553
GnrdM4ncJWMayGzmbVbmzivcITau21uPVlhDjSUAKWsQHxnD9rECQUrXyIQKiHJZ
NcPqqqkfV9Ml0D8y6YCmROhbUh0WB6M52c7Dibja1OYUSAHTGSF82fzIumU2RW8q
Ivx+7W3N+I4k5wh5ilDw1P5VKatTUxS7R9MFtzOrPq5JNl3dIdvAWzPguC7jliYZ
QvQsTy1Pp+CLFI0lpOFe9m4XWCyhy9eBWJp94P3Wqfb5uae5/6zmYMTaR8OA4my3
nmtwqhQc2dpknV3bajsin8snshbnED/pRM+MUmOl0F2eoYYVzJo1oFApJYBRcAw9
7otxQg0sH/LDgus893mSLspzEKXVTuqhQJ5JcK1ESDiPq8xLSrrg3EbbmylwwaiM
XWD+Qkf9FiZLattlOrATqyWW73SmN2yXw6RGtIGWBbz7gGysJmupf3OKQfp3mpvw
FbL/KsR+ZW4JfHSGkF01UdRP9Gm09SCOFJbf9t2hf+ifw2pMUQKwvYFg13DY1ue0
aJzFjxoRMRg7jNdXYdzW7LX4FtJBiZpmDKWNwlMR2lIaeEWIoRll4/G440MJZYYc
Qxmq90FL7cmg+jfuVwhiSXNm0Cd5i/GjJ6wcx3fpcvFJClGGv6y4JqOxkeTh46ie
BEB4bKQtWg3M6YyCJlCP/jCRrcz1WHEx5oXBAowPTzgbpystJxG2KAyw//COtQhn
B7dmpAeTUOZE60zuqwwFShVNDSrKoh70pjlLRHRIyQC/cBJyHLIK9vy3UiRCiJQf
VEwZxA8H0j750WkVpsjL973O1Y9Nr5/Qojog0wjxvn9vFkEjQydxkYzReWZNeV8m
qskBdDvDltULAFMSAGPr9fn+NHhzmhQZUc16hq7LkY7igH3xfNWHX9sZ1Z9MYiFm
XphaRD4riCEIOYeAblceLYVYHZ3nz0sC9wj9ZHF8vjO4RA6nwaNjtDpkGJCO8ZDL
Byr3VZS6Rn4eWkQUrr5/AMiuQgMM67jwyzkqAbM75nMmOjHuEnn/sWqak4Z1u/Kf
IQ17dPDns16kXrbr0sSyJXQiQjUZPT+la+iqMB0DTHsXe7pGGRdXcttufgWW7fAt
NXvgusi4MSGu1AGFOcxsx6nNuDdWOcWX5CsnzCYwsFAIq684CKJEccRd4otVAJi2
sC8YgvgliPoAXJk8DIKae0NFX/ZKFaLU0Ozx+KMzyUMeeKI3vBtzm0RyFv6GTgmC
NcOf+Zzs38/LR/Gz8wnfwCMVTpZnYugstMSqz9kUGB9tt+frscmrdSfBRWpaWd0q
7Jcbqlz5+TleRh6JhLnjfisfULQmY5EE1ybOTtwFbDQLaLh8237DlEvHFdnOHIa0
uXuKWcAWotgI8Rf+cR14rCXnhui3nKYrv3mb7C5L1dfMBmbZhtclZPewONvBYQEf
azYw2MxXiN6p61r9BPCvtztpDI6xqlZ6JJzyWxNln3Jb6z82oJs1ioFtFTEt1UsW
s5nccDpJU8fKf71yYITHr9bz0rAwTUGof8ogdl3CpC16QptmL1c2x7WMnc5egseK
8f0wDaGsDvzfutRk445ByRWRI3Xc7JstVY99whxqXZRKo22WorIQSJri3GrbdeO6
rBKyhmjm2Hfj+8tcSvu8yyGTHyo6xiqFilRyMgGuXScn6vUml6kS6Mw6ySGk/Fbi
zYX6dyU360qJNPJn8yFYF0wFiz//+nxSg5GQuEW+9itZK0BCvuPZxWo5ufJ4rF9h
D7UmleIdAB9QXX/977nAcl2JGbmrLjPc6Fj1HTGDo27nsNMMecpc9cXadCJ8T/Uf
uPlohEQmUtxRZ/6DQuGX9xWqOsdh+XqTgGkF8xns15vI0bGD+i/oPcJgl5Em553j
gcEuZ5pNNEqNM1rUYeHvAntHSTsLjnzyU3ZoANpglL5pUIgckKnu9KXX/+IXNvz3
ejkXUee9RMEglCIYGx+mtRPw6bqpYfPJy4hVF7z5muW6qsJ9KtUfnrKuhx8iuZME
A451Wd69vRpEQHoiU8dHyQqmz885v2vHfjeEUWPUXo0rf9iSgGkkqBhQTquAGSAH
xCCpd/NjpQX/+g7h/6106qfliWz7OIwpNdQxyyDES6qY4xxtkwkV9fHb0xecexir
lFLtGi4arGH22sqBY56rQiy5kpNXodvx3hmefEK9cm7yZ/0ubjzpSrOt16S41Kx8
nXZiczXMui/etgGhFSUBJFyHk0RUsOzAGNOzaMIhAi9ZiiY/VI6cxno2FyIHXTny
gzgT2jq5a8q/36K0zC+xjUH2msIRcp0Ur0HU3Tvg8FLBptT9TAmNGSFgajzne2MW
u+4fXqGcWYNH6gihUxAPtb9M9L+VsY9S402nPhRAwS1knn/qZs4ikudgHwENCGNs
uKgaYGxQI4NozPKqdzgkVeGqmC1OJSTrQFY4R5Hs9CEAAgHtdn5ZHVzp0DGJrJZu
g65wJAa0UzulmXVvuuqtwJKKWdHCW+V0Xxpbp12EXGniBaGh1DTiUWDsjvyNeYS9
JRCMr7MGsfYWzq/akC2pglnwwgecqYUIDWIWO7xQBwekRL6XByfdV4BU7ndPur5+
43qQK0CLfAo/IoECpUBqF6cTMm2WRnxz/6lnWwms0SoOskqF6d/sS8PDCWsc2ynj
bAFP7NZz1fnC4Utg0U2GSjToFAO4snW2gaiFfrn6uNFAdm3JznhWFoaZil6nE6Sm
J8Gqz4MEaebusL/x6xvRE6c5wsW5WKcSLcpyOOTuVFwiyzHmyoY+1TVg0XplCMgl
7f6TSMfw9UhCmZGtuU9V8CfQGCfPGestoLosA7p3gzKNpYCyZh29bG81CO9YZd9o
Uo4JjoKypL/tcYATHDciFsXm0Bmo+hfrBIljmEMeWvtEIQVycq01MbuP0WEsMp2t
FmfjzuzFXbBwx7ji6H6QKe+fCCVzgcBjSVqFks1vIYVvsMOYsfMa6AxQj8J8rLII
e1r95o31jrHtsTcm15WINtZjw2QniQq5xtSOwM9m4oKWj9zOF+NmQ4fDwOviX96n
eLhTiKHaWVfkBezQbO2a+XcVvMkLP5+zmbetRvdiEIvhscTtyCmgQWt901TuK8Zr
kytLE8SJYvitwgGFYpDqGBrk4MxyWt1El8HIfPVgmtpkIdmTXVYVGNSCCIzrZqoz
k2EdC/SbE5r5rHSByt8tOd/pX+rAYN3h9/qttyCFaNXO7XuMzmLn6alIgpocEe0C
6jnZPOK2pH0074Sm0V3O2Z/7f2bKsxg49uZF2NThIxZvuHp4Er9xqe/yxrm5ceEH
07OEGshuO6H+HvCUQHoT0lNbzz9evGzqu5Jf8MaBlYQzWHVfr4sBLrRsFxMXM7FC
aQsFmt/9YHVZCqhn8DZDeqPtffwy2k6XTnCyFqwSmyutd7OE/DceuyHZ/Ml92GjH
+xjM4YvmdubTHY8Ok31LH8xL20k7Xgob30ItjLrFTOrSuOsyMuNm4lgIOJGDgghZ
pORRlewcYvbrVVNrspCQdT+Fbgk//lVydmxY0d8MqkDwYjTOokpdqATJLwkZbzq3
2c/6Ql5/qWH7DKSoKhludPph1HRWPSbo7SVxDm2Mt0G9bAFy9Pq67VcosqGonSUp
gNoJ4Jwon4otHyoZG82arNHB8GvxXDnwroEq54zukMXXSU8M0QvPl9zYQUopOdjV
If47GZZ1f+JruNEHPTz2OS5ghLSu498eNORpxkjqeiubSFkZahU6NQZzgSIaBb3L
ir0zh7Kn2s8R48xIP3JCFF4yP4XaRIOPPtwCh5SXY6U5sjK5w4ULAI1J4zcAG2uv
8m9Pj3Yf0y9tG746ifXiIsE8MblxZBeDsWtRsUgVdZnNjlgul0z1ItpF4+LerFhU
k0Nb+27pIsdwxXL6M4Lea/mn37zD/rFrmt78KifJapRpaao8tQG7KX4YEBIHu0pF
EuIspsRfjmzl6GiME9AOzENX/qhYznZ/VXQSNqZOp02hAbAblkj6FCxZgWYnVi65
Lyd6YoMX4z5ctUx5topMoxgYuFVIMaDdFfAeeJKD1xtstJ0EpOovPSIlLMRrAF/t
FHNPUUIkZRssvJrpcabbYWvnhF9IAlyCw8OQRNLcyk1lsacFryhogW5ZJgdPYZ7j
A+wO5hOEfOYU1J9vDQ9H83CuWtW4Vz2o4qhm6ip4bb3PAZU0Yy5mYQhV+9qvarlU
ta00xbb5VluHn5bziOUFAjc2fGbOJ/GL/ur+EiVoQOD569SjdP7kTNsBM2hsAJZf
Nq7q7NxyhxQMyvJDHvfPiDyYgEi8JuX3Nanoj2bW5d+ftI3j1XLU9wJ3XfvIMr3X
nLxLhJz+sXRRqZc7+XjHm2+uztuI35MN1r98cGnNnO1p+TDAtuSPSvS9Ch4X5Lq+
0i+iqt1DE+hMgG5TThPRnjfwlMZEDdwOFh+O7Xr4yU7V5jzOYlsEte3FYgKBUYbR
vQf+ttb1IqSc0hTvmvXrj02Ulgchmv2id2t2cuR/ZaFh1BkQ6dUIbFj8y/k9JFX8
4Nm43YvMWkSsMm3FFxbmImTaZ0dxz0d21id5hZqW1PrYtQd5GRgAsP5hTPuDXbTW
aGAbGtErUmaL6BCP7hWQe0l16/p5MWSkl7v4G0RCas811DtKR7KTtIM+3kncBweD
B9ks3IL00vVhwredH1W/aYxO9F+30zqIekhC7nDozWxFkFcFX7qnllT3EAKDoZV3
Bj8toMZmgwDQo1RKDYoW/U2XPUt8cUrEG3P+f+84yzQqL67VfBPiBzp+3HvxRfRg
3ny24QOmIUkSxUPyziYU/cWLv+x89n8/zZwWjRDFduYb9gT4pqLqOhQp+iJhv8XT
OeoIV5XbH4cG0Phm1RfdTMM/4zdRDvs06lDfA3el4Wq/IHcpxebznWIOMiOzF93v
U+BBPbflARc2ih7E13KDOGsmvcNepVvqQmH2vMTJWfsYfWQRAveMn+muHZtwSaRP
q+8pl77SmGVFHf1ymTtF0Aor0RjPE4x4bPHSLI/XRka/LR+zYQehiXxHLb0g9peb
jbiwKKnIww1EwY0W3U69Dk5Cy2L+Y9TFsGpOyQYG5aGlVE5yprU7fYu6n28aIHrB
Fp9BQZLPixK9gF4X8xCCqHRGzOAJlf6LXMaH422n+fXvc/htgNXBQvwKt0VsDFr4
X3JLULao9MaO5cRKALG+kdxivBFX/KlseeiQGio3XyzSoHFW38Awsll94Dk7xS/O
Y7n3x888Tx/kCJZrXnLt0pP3ddcC+nAonyYwFsBXmMp2F3SBAfY2fJZrVsuOi+Ss
5JZxt0Xp3YoatLZTCOiXaPu2WZAXMiB/xBdTNiOKn4u2WIOA6gaSCbxVEE9zXSP+
t38zge1b8Vdj89T3xjYSgK9l0K34QSLOsKBzHdEe2xwb1Tw6oJkHTcSoEKMGormn
UOBAvBbNmz4xJQXrybmYrVlp2pnIAsHaDWaAO5XWnuVDB26xx7LcoHoPnfcEMfqo
CvyW3VTX9HjrzhYuVus/eGRlUZ7OqF74I6TFQMMhloZqRpRH1l5ytgMjjlcoAVbb
kl1KCi6/R5YgE243g6gNgbAZ+UXQHtrJUahTpMNGUMd56Td/bIrl8V5nASr7iVrU
C+5BkA0OcvlHgyYZdm/RdQacWNDyMcmQn6GbQjc4Z1pxHvkHe6WqMQvar58u5wWv
4yCOyH32sY2GRe+P5hVILq850IlY2OVZjajf3Nbqg1kw0Za61hGtPEBSLwWAU80N
rHhvz05z7dUis1Q4yRgIvf3bJbM/G/kAFiZWir+IA8K9pXn9R2bxaVxBAVPcxi8O
wwe/R/BEIQAqJlsue34H7vPJ4eLQY/ZRpOgtx1ljGqq1i1vDyzEEzH4y7BdvOO5+
nRnkqKeLW0iL51AviUkvTzALM/WU8wCHIHi1qgDFv+CCKyJWeEF/vhAXrbv2F1nw
FuI3EgwKLZUmvVZ5/oOX5qH9KD1VOkokNzC2b8wf9RnAmIX2x9xCN6Vuv2HABSzq
bZTyPbogjk72nea9m0CAvByucL6a/f/W4riRZqwK/bokXFbBP5EybTlKtQMZhKU+
PGzT9a4P3xxaI5aVJDFCp5G6H/UWXJpAMw7y07LliIx63yuTTPzJm8UQMaZkjeuN
Ano9YZTPnm33FmLeYROBaHQ+8nkBqylPkjHtT47/pmnjVjhLhSkjzhKrPr3DWIeh
sMFJr5C4kzzPqWKyPn4dP+da1hKmBuJ8kgXgxgKJ6e61ke9fr2FXUaHzKhx9Th0Z
S+buFnUXwmKcKDjRYnTLdJ98i9VBKF+aP2puOo9jXLlgbbKQNkFFmNprwlW9dclu
RJUHo+5bG7YI24xGkXYIIAtRLFbqYb/kYS/RyEoE0FJL1TrwElmSQr2eMlLxqv6w
CzEqBlGeYdJvwc3oJdj2ZQvFAVkWsaJlnQJxEMFw72TQMyPsiXYYfWMt2JODg2EC
iChxE+4ATjLjTBlXT4F9HM2j/TI+NI09vYpO2ZVz0X1W3Xf+pZ9E6BeCZhr03KtS
Q15r5H1JRJHJq6oUV6ExPtzsYfu7GSCHKqmsQZmSPP9aY0sdkBAAnw84xHteCzT+
TyNKYlzfbVI517sua2EOFXMMEpptMFt1MeQ58sTEUY0L/3qJGRZ62UMJ8MeM9W+i
LfY7xjEKllTZh+ebkPFUYiix3yvZXRJWZLqjy76AmLj1YFSeS53m+iVPOM1tYAP3
6RltPFgAXw2BkHZWQzehS44EIs9QkFZxjSaoKywb1AVFuuY+YWkzxhRgvGQ/YN6t
CXOYQP4hX8pyk2wbf6dwp/f5mruww0mO8Ea8BNjO+KCKtfbHizvo5L6dRgrIMQiM
WNpJSy1+Rk/GXqbZxmA1zU6xhoqP7KcNsQRmXdgdexrVXLllMZTDa+DtFXiUnWoJ
kZAihJjcTmnr8b8c5p6MKdcDCAP2WlNTVV8nVlyJVC0y6wd9y6ppBe48Jkz2PKZM
Ya1TmxWbHGkjBk+UVlVWDd7fCrtTYRnaBrnWFY0dytjroIdTlr+M680XWH0l/9+q
o9GS/WapFRrivjglSEufAku9cuazLFgfR8Qls/1FoeOOunA0k0RCj6TiLpf+55DI
uiiSMm/ljE1bCNrim32diSAt6ED5iD3XzhayaqfBWlye0OFAEKnyjvIsMryW6Kri
XBCaVacHN86bpBXKaf+S+2aUnFR68plAj2Puil7hPcafjtPGcAVKbbjSRI27oop+
/GoY5vNt/cx+RJwT1HNwsyS8UMCUuhmNnDBqrvtBXXyPHqCbD5XUsvgtQsLpFfoj
CSJbW0tHFD4AO6QqKHzH5OAngsqv6F/SdkMz9SUm/jwjE0NefubwIBYbrelTNRFf
92UdHrMfjcOKNOv6iIpUQkB8z3PUECNjEY6MmhjVxF130g+pX15yNHfZu59L6POm
X0zatTNhs7NWDlrqN0h+Ry8rxI2FDgvu2Eg45B4mDlnccrJOGjqoKPD/iuo+bwCg
2/If6H5/sX0/EYXfRKA6QPgvvTDx5WUlHMAvRbLCL3tp+yHTgF4aKmuJIJPfsVwJ
j8jMF3LZmGjO/e+sX3P4T8qOvR4xcnhK54u5iso0FnOADAfzA0Ax9TAsL3nSoN3I
fCzQZxaDxBduxpvpJDpczdINwIwip20wTJ5A70oVsXIIQ1VZuuRvdeqY+svioDNc
rPz8F1kCV2Dx4Vvwq3F9fZ275S3lUx5w8ubkij37NPSWqPreU0elG4VAJth0BIFq
NCqYGGgejA1TMSZ+07+hWefz8z0xWsSDR7G1lXRpLB6682AKSqiCYU6/FzOLUVzP
ilWk7VkKticTDTFhRaQFdiMmAz907yrPr+bGO/bvEFsLbk/qluqXmJlBfGXt761d
BFWmoIvD0CDvasNdSMxyBu7e1GLLrjWu/CDe1f9vn/Lxdg7R1QQDEw4IhgJojshm
2vy+6XvduxsrnJtm3Mn0BPeJ/Px6QudNbdjP0VpWv7DoXDn0TA2mTJ1zfna5zImf
pcCyb5eG9CdTNURkxH4aiCaafGwwRZ6fpAczlZWNSWQPKDmxxDQhkFQKw/0W2MXp
1Ve84XtSGKv/xkzhkzr4JwrhU7PZG73q2e+zOxVYXk9J522SV/IyahRY0H38/me6
zRVarg5G0ch4etOaRGdsTYyhp9R4UhN+cFS4+WMqAXGqfDVrOXZSsqcD+j2H7uAv
1DDGY8soIycdgpdHq6eUv+jp4ygRtnxffkAaEOgTuNQNMdiDb93W2HaFjz9AztIs
RkcM2w55d3yjKwndmVmtFED9kUIEQUCN/Ch+lVMQDKRMAOwrYv2oXZz+1jkZdVIT
LiIFyVtLqIIfj71VXywHMjKws+kE/4CWrJ5NddrLFQmyJjsTIj0/mWfX6gwLnW2v
3KRM/TXm1GtDFZ4wtq3dT0vvqNQA2MBGp3EwW5gsatElyAF60Y4uZDAm3qklZPdN
379gWbcwOwul3lerFJD7bjtxcnl8FjLrgtQJ1dNaX2GDzrnBZ76dv3O6lwblO8ZG
TiynSkE/N2Ub56vefh8gTKPgz5D1E899Aip/PWJI1qoQCXspOC5s/KI2eV0+BlO1
QiC3QKdaKtKLRpvkClmqMvlnzO8s+0IS9JNZdjT+zoql0ornnWA1Mo2+/1gaAYCZ
jcB9WX1GzkrNljQYhCEi5mrkBgJhN60pX9LXwLfZA6Zkguvik42DriQh04er9nI/
1WxBzjJ4ZrX3Gp2qEkToXep8QPBsUmgGLBqwdk0anbHQ44bZ0XIYfBF5dbxC45To
X04K5GrZ3cM3E8X4VQZgBa5b1s9TagiqJaWJB0JtstvAnVC6KpCDkIOr4twWWRbY
z+yB/fOuSf/rYOJ9WBFgzGCTp9pskzjnKPpp+qytndkXoV0cZsxlHZAAjIWEDNmW
m3w0TLltcGAHKZS/NNGKG7zbeQlSJepxEQkPqR0RGs6/0ARiUxI1apbbU59F5Y0F
TnYS3SDKWU89YFsmHm0jJZUmG9Ew7m07UNAk4vaXoLpgn4WtvOqeCsSIG+ymc8xD
JNvkZeJmGwkrMlUDVMqJOjhRMv2+OlETW8b86G4FTWFD7q2ukdcmAlqjcbdnAubr
nJV5uDc13Mk+n4kAciVL7l1Wz/Ev/VohFxMwGayaegbrhct1IqQPKy3NkG/2HZoT
dGX5gmg9VGG7O7cbpNG/gAYkUwyS+NzNHXW+TMM9zDUfsxv7PNYlkEYmzcvxS3aw
hf133QMlPelcvYl+HUKWVEl40AGvO6t6HfoEZHCeNccOkzfTa1YtCdahdGMEnMFl
mJacA1tbkU5cDxnCxTbVgKBOjrG0xQnvJFMEtR/OX4HObSlAQ/3KCNPfiIKI6Bn6
kvlkcITvZRMmuaKyivol3lL44RhjOtcJwMxlEBxeP7zQqE5+LNUoXLPFDBJvYx53
WFHWCdWMR+IbbDZxDYCJ+WbsKDlL3dzhlMLlPvm2KPBZ2X3+mnn6AZ+hmFxJS0N7
Arszm5j02NpT3lylR9niHOTJ2qCFZMG/L6O9nqLZzrznkC6NEISI/UpSi9OnnXjF
w7GtUEA1MlI8TW1J76ku8fidLbeKozUldoooDEs2AH4oaRSCkWu9iTS9JdhgNPMX
i924uqRfYGA+1qKuhW+ufpIUBcWrMGsF3eF69R+cMFUB1DVcJZZrip9eZVf2Vu10
pfWmdHeiKySkM8hJzY6WTwM8B7isBjglz7xhgaPMwPgBaaV2m/u7rMozTrSXCmZi
xWt1SQ9vC5ERbBGkjdrQMnjMC3HxlKFIjXjbYWpB3N3uqnUqHMs5nxiCw02lLXcf
ElUq2MxS5/0BDUVb+dKm2Qk+E1XhXO47RIXbQtfKhoikjooS5emMp737XNv2ORK1
GTG0YKjfw6a+KEgUYznKV0IyhNe7mGCbsiXxHIb3kHB+BJr75EmE9GMSZiDGr9CT
TIj7cdV7b5RjOFcYvzX2uGzhOfEDLjQZMFIDXkxzZkkoEvSrfVXb6CL065fEuLSo
6xLMbfkllXYLajdQslIF5IpOho+bV6vY0eOVRw/rdGHXSkq2j8I68La63R/uQklv
trFXJHdA/sgIOPAezIj/Y0s6w5tHh69seAEpwc1qcbSivelNKecYwImi4bKo262q
l3PBDMJX3vvei3aLZ5pu8WQf8+b7ZFcl8cll8U2QBM6ySKo3HUb0EK1WXsFregRp
m5pLNVrsFjYMPGQwRcUxm9od5w0ioEqoAwrQ7Mg2dSsh53QtOAtU03/h0RLneXCh
picPCZFwOwrMT9S1oR+z94PHaYAKxEkvWf/mxXKGRvwm1muku7Qkjosw49XCwKmI
eWVU3wC2ODNba0EzhgWM+xpRQaWcLIEJK1RhIA56UOjo3NlVRoT+aFSqb+0skOUB
89KyQKesaKGsGdkXPhASCmA6dcQ7tyXyqX2eyvVMWcpcydTmVlZJPGcvB44VnauQ
4mmXYZJo9zMwmZlk6F6HoKD6GveOdpzi33lJ/Vc+7PFT6VO4fA6/oOUJWnJYjQoY
J6WUrsAwZVAccIgXbYgc4Kd2V2bWFsNumF1JKYgK7PHaMXpRAdfYh2Mr53eafeVR
GjC+a+lx4GuAzdK69v6FhXwIBAHeko/as9iADlRK+rHla/1ASiEuIWTqtUoiJicm
7EfrpwNB0SNnPiiLEeR/vBdJMCpSiV/X4qXKExmOZwo+T5B3a/A8nwiWyKzKY+S2
ggSZa2acg4nGDZByuWCVFr1cUKGk5EYSNDixP598hOTo409o/TcNfHM+d9x2VnTN
muvvXVDisLvcSQDMo3EGGrQmLBl99EjY2LLxiUmcDY7R2/Bu4rmTI2pWjIW1bfyG
FaVUg3xwuybMEGjT54d67zXBIMr3HSUVwJK3iqhQ7LjwMaL6so1cosTklMDRsCeA
J+Td2yT/QUOk7ODxqYVVGKB/3fXD5n2OZkM6kHxd6w5VRhIQ+lu0CZlDvCgBk7lC
8Mq7X82B27FZnNw65gSXMhX1ySeWAqxhzDHM2Ns2XbOXGzEjegZyls3za/dytTYh
SxB9ilREhaSY0Uhqt1yfco02G40ldQWHZPtknWJMXpotxBTdYoPGwNVXSM1rj5Sh
jDU4HTubI4I/EbiQE3puXRu+USVFGFj97K061Z0RSoNQCCCZ7axZmWv2YNk/5nFF
Gr2eyKGP3WOlbDcfbdNuJdgGyWjOvctO+uvANJkgUCDKSrda0hMZw3Jspjd/SvWr
Ax01joAJvtrBuv+3NXeDP3UbidWEOnzvVgmk44xc0XEUlLd/qC8oqmpVbrcrAE/0
NR6VT7FGak7Povp1zM39hy5GblfthG1Uq8RGjeWP0KG/2OGypaK6Ey+G4u1VKrZM
E8uVJMTDdAyXqfvLc0UT5/TqePSSnsXiDRr++/wV7Sm529P2xk/09ZAGu7YuIpff
jWuI//TEndmN7M2eqGtasXtsmuo5CuBkT5fUOmZtn++m/UnFHiElTY67YY2nJ7q+
eihB2XFie8cjhFGuV+dw0GI+uv4lcH/CZ4OllvwzFn+dr64xyH5IKbNCL6MVOStB
qsaIaKZBz+84W88ldIPsbpr5HJ2SFRKk8m9/1NE1Y9ZsynR0caZZkar4geTSpMX2
+luss1Cm2J4S/V5Y7FcSaP45Y4WmXLGTlmTMM1VzU0kMpdrFpkbA7akfGlB+pXRy
DthXAXSQmVGKvI+0kGiTzyIYaIO6ifvCPKtNBTQEEKJTtiWxP+oVbEeBLKdJyP79
o6ZIoJuIl0gVAaREX+jojr6xMbJwlr03cZpM4mEKN9S2UAn/FMnOc4xnUsOE3oBl
T0lExLrQaeK9suVAKaNpigT8WCachrF5puYZNQbKLjIIxiUPg4bBcWmeys+P5hIO
EoOpet5kBvePkLi4hXk36+se9xlgjf3T1jZVF8znAlnXmTpo2Tzm6/MgVn0zAz9M
xYyx4W2UlAOrqPFbIpWnFaYDLRZE4Uu6FGME/NXWTAffcvWVkwjul5cqDzVipjVo
IusjHZ+jg4XW4kEwPMmrVLEss9RepeYT91s0rHT2AhMAFO6GLZcucjqf7Yd9Zreh
6EccCr+1ZkV3IcWv5AK/uvy0zvW5CAwiBlg8+w2A2g21VrdPfQtVJsdaThBoY+be
HpzQEb8lJc1PDLJ7X5JqYrXBt6dESPOGBXPU8LhR/Emnh6OjDEzfdCSoH7A5kyCi
/nkSpahf5cOXXvh6CLoNGY1MZZ7X5WCoi9zK395zPSDsyLNiB+c9RWoowTeY5HUg
6MUjF3/w+8Za00MT/9S2PKsp6AWNN2Mg4HyaGrp/w/sky7xXLkY33ZWMEbtcZV49
3ejcoMs4jJH1PKJCth2y4/ZjsyZbPvR9tRr3J6rn0UkdvXPQrGuLEx2C45RYDBrM
PAaXDnkrjd3oR34dB46V15cuFY46SL3DtB+fPqZkXDaLpnqBsosd92PCMK7Ue+TZ
+V0RLzh5nGZxf4LfwzsjmzYPtXOyyYxHN7tjVezscpgGKRbntOSgRJTR7O5GF//6
t75dju2oxzT5jqdThl9YcH8ODBfWeevj1JRDVFH/NpY3tbY3011Pidp9k4EWeUmX
s0tfy1P8YQqgPQjNoAQjwEED7Rz2QD83J/W76UAXZeKBl4mZeXSTIjQFkN+rZ06r
mkSbliKO5a3FReupTnTTB+/BxWDCPgFcBMpd5sglgA6kDualHMKTW8xPL9nTJftW
+Kxuzt+tTvUCnyFxlHZaj5kHZEeP/DGuL3MrFWNkHCruzC5Tjrj8jNPmkm6m5LWa
nvO4oum/X9NQQghiBcl4y4kMS8SxvJwuqk2C11B011dKZK7lgVBVldRo78E6lwAb
2YQIJoimGpJUG2x2OIgrQJsM1Q+xLg7XQVoCcWA9O/rIr9MShgJwKymraBHajukc
pkghjaikk+6FjJ/c2DfQA0Q9GztqCTXZFBJa04I+NQSqmbXI1i513Dn45oIk65iY
TT0S9n/lr3O0J7nfac5Ii5VJnOIgUa0fA1ozai4GbQjI4oQ9Kicao8238DTHJg27
AQb4HXSZHLckX2e5P1CyTHBn9z72XobUJzJCcU4n7GCp7rq6cko9HyR7teCdMIZo
2GrSHDtargvjYUUja/Cqock5E29CosIrCuNkkhljtdEMdXdJNh/fMEb7lxuZlj08
Kbn7o7mhlrNfsH5SJ7a7XJyDJBTATwUEREbfeCFv6jG6+EmJ6iYFv+Vm7eUupEQm
QsFtLN4J/ZBpltJ/EnC9Vyi3ubDhIATVWkrnJML18FNbT3lOarb889/tsekuAse3
B4ppwOg78nOZtsVSy408FMp3PhY4c+qwjhk+tLjtWodjfbJK1yRei1hQQHZL4lh1
0SXYpeiIDAI+Q9TYp7SFyyNNtUGXpgjWiERxPh01GGgUcOTEAEteGadKl2bSc/Ov
9cLNCQT8AurB/FwzjNzV2p7zh9ONMMaeePEzr7yHNl4PLJiR38jWRU3rcWDFQS3E
`protect END_PROTECTED