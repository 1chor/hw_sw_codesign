-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
NWGGvKqgMI4iwm2MrZgXcsW62+f6yAuBnKFhu6uwlbM2Zpcb9147qdoYPjqgauXR
WKUWEnk+TBi3vgkZQMevJovB8t66mKJyYkr7a7pQNpt0lR6i6/AAWGh68hxLPRbL
LLLhvZBB9xiMSGe1qezDm9PezmhlqioaGxXIGkIMKRs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12544)
`protect data_block
2U9K9t95qncvV/8Hf4A8yyXslXeiHu3T9jpkKUuIepCQ8GuSYgFq36l8LzlUpYUI
tp6ls0XFxR/WxXJqXiutWcgC67URx6KJgVsubW91MX3vXkPNZa4bT6cI5KZfyJbX
Jlj3s3pnA/bx1u6lH+pBNAAyDWFOLES2v9RHj4EkWfPRnihH5haeUVATKWgTC9g8
2SlssLAQBYG4Or4NCfBZOE07qq3PZ6Qmbk5ZzfYpn+mqEkLdUIVKYXRK0wDW1GqI
Q3+5ZXMX4CyP+NgVdqi2+UnsHxiiCmOcxBhwtwylOAb/Jj0OFdPNySuFzsOZkbmc
XN961UJngA1hSKVHktz9WTHf7yu/I2RoaWC+IwoxFsfzP2DhnaRkK5G7zseizynu
ZwPzIb84crCHByXcy+1oktucMbrSoFiVNyAZGLsL2JdWz+k/Bg7L2v+qjv2qGB8K
lwQH+QBEkOG/pN9UGU/WKxsmvY2RdyBoXjmIS5+BRvCU2DLtq0Bxy2K750NaKFw/
yTXP8Nl0XMJrOVi6ic59xL6q2Z/egKasJiB6VBjeKGdqfAxhusFoKZ3lLmfoRPJD
VTY3q2NpiOtn0lMOglHa/VTolTONV+zHJeV7Cp+I2ff7/NPj/MBaW6yEfNIx9Z1U
XWyw56TFL4Kw3t/HGjxJxMdwcpgHtjkR45SR3TwiRCWfok3DzMSrru/BVnQ+q8kH
9Ph1mpNKSlZaKO6GQVVARqCsAv8MjmTvOFTHPFca5hxg7VtBJyoUiovMDumt9Ch6
9ILuqQC71U8PKo4TEhgbpEqyRzNP+f7m6SfZGC/Hwtte28+E3yc3ElvvMCZttM4R
8GpdMJBgeicsNHKgXqdYQPH/iq2auR9LtIff9HSCVHQKNvPm4shnkmbIxlb4L6o7
rSc6OaqrSkRUv9Y/SJbLas+705gBk+9Ik/vb/Ngz+X1/p5CbNlICuaGX1sLE4Mpi
eM11GT0pBTEb8CkGxlBgoGMd7Nt0UV5d16XmcRNJHsONk/2JBpm3WD4cKoU1DOkl
nR/PO0WmQgHtloV6u7KHkg/N/pFZFErIWxKMQskGM5+EvpvcMEAbWatSZ+kw6Yz7
MQLJHe3H8RaJY7O49n08MEgbCHlPzmOjoqHHIiKYwdqQA4zlY16vcd/AHwZVLXgO
WPrw431xy9Jto44mrxgSlZAP835dkRmAfoYBgV5ePiYafDDcbuTKLo3zopDLkpIm
g4nug46CANJLEw84Y4RtQVnp/ZP5pTyxhbtualj6gkmeECSzOWo4tYnBE0na+uQX
PWtoorcpBjYYVKp45OFcFR7H97m7x7Tj0DfbwC9rdBsUHpcxCXXzqXetUEenfGIU
bIeaDX+tFfzR663wQb1Y1uikgvIC/IbrsjiMffQ+87q/n94lr8SBQj4SJTaGPfT2
N46mLFol7li6T1aph6jMfATs1i4OMmCNGsy/DVObxc71Z1TWLfHyS4dSfCt/lNmq
Za2Q8U4p4lJbGtM2fPDWC9QBbgUkcYKbZdxTTqSjuNylFV2yIEKGJkeQOb/DSoCe
DvRAbXsEKeq7FwcFcLTYPAIm4qazOsamMR25E3mUc3GOdPi5LrB9ADXrUYn978g2
GuGsXSM+Zfu9cafeMbWQgKhjsK6Q8zcPPmYdCo0ifz/7QM1Pc9LGbLUvMVP/mp2v
NU+6251VnxJgx8knjyBkA4bhLEdMx+7SuvowU+pa0aTz5H89WHSURK6a5geL2Gsg
Ju7yiktiwuXpz02NMwRYg4Jmfs71KwjYKpUBJc7RKkkbuPHSgG4+tkKnPb/+EL0m
HSKutIugdZZ7pS++USbWFqRjbQRxXm6AMG8ELRp4tAWuMVqG6xvcQkz11xX754Ap
FVFz+OCUqoK5AbOx+pwc2+Nt8Zc5rml7BQ/cpUx6OJUqeI6iCPYU3CxsAvppKvWK
ky6LCm6eXXYnrovQ082QGas7GH/RZ4aTSCGQsuwQ09VzV7OqUxJJRoEIumPz4iYo
z7WckHXCU4aPGf1XmcGKf4DMg9yED26HSEvbGAPFmerHbjJHcokLlCkXB4+Ldsal
alxTiCefxTJoVTkflWRxciYs8+F3iI0pkrA49m3xe07RZczfmipN/QosQFnpItg8
H8cEZUpNZRHJ5W8tDfMFL9wHU0Y0KgqzDFe0LV9YyDMrlnssNbNi87Iyfi3tV4zF
rdqCP+pWRlQsk+pKzVaYoJvSi3vdckKpRFNgWDykMhK4H9Mlj8zK6DaU2+qrPjTP
af0g/WNQcYa4RD+98W0VlW7wGUSAAR7nkWYCMkxgED1ECPzIxzNDvZ1HGwLhYXih
+x6kA3dpkwRKutv7Mh+QBYG5oSjpC/szO4oDvA7gv7yFX537vx/rxQjBZHXKIvmf
mOiJ6TXXYYO4IjduJ+VdZAjpTBK2wwtwLesP7U+WjsiI1VDYwNPw63EFVD5Jk6zu
mhlsEk1Fu0P9VEOJ2iuQ63wj77P0ppvKc5Y1OFPkZsEp2k25fEnsVe3Iu+XZ1pXh
k0i1SIJMjgmQ/0i5qE8DNGwmoc52OOJvvS2l2H0nTTOzRZuWv1er1vR6dVn15IiP
1/n6V5Hy23UU1gbsWR2XmrBeErvRTLSbcyHDsC+02WCIDgZ2bKmuM+qT144fU14x
Zye6CaGod3PzeES+4dfKM/Ys3AC935l3gEPrgvvYT+OFBE5TlH0GIu/Tw/AtS30j
OE2fBZHmSy4kNz0/l9p2psHV3d9Fo2wEljxzfo7/PwTzjnq+k7MsSN/SP9EFXJb6
+Wwsk+5QlOKY/K03GGkB9jkANrAh1xF+gXxnDKTg/R7g9VwT9c8EwzimpWduZZCP
poHK4HuNDxy/Mu/qi7IOBNOEThmeu7M+abakRDjsNLT+1iyuhN5g50pxhrxRzFNw
JKeD4jOssGQVh7HKcs9UN2apPQOnbqWqxiqw0kUn8Ug0g0MaWQ2L3WIMdvTk4hi2
n187VqjMsF5LsKVce6vVkcZ9OjxSJXb9DON7VdlhZBXMtkv0mTVedS1fX5Berx+b
XW+9RJB6LUBntJDXXfnaXWK0pnJM0tqa2XXzabNiu5zT80DXgU/OM8NA/xQhpwBo
TFgevemN4GLJVTtj2PhV7B+i1cmQxy8CSSIZZIngcCuXvCs+ESPwgy5+E9ahq+0v
SfvyLx330TP45XcqfxK074Iqxm9AGnjBUqwdQTDM+n6kDALqYLN28BmQL/uQf5Fw
YEfcWLToGlgXYXZ5pJN+smRCL++mBPbmR1QVmi/w5fhSNUzISSnEMYE+8Mt4QPK/
8v7mZh8CzAG/1IK1SIjCBI4OSiAaKajEYH/TP0xnpzr/XI9AnX/KddfMn2X1g0YW
vazYeakrfZ5ZvYGCi42JYMugAeScz/vBfRNCYCTRrv7dcH1UlzQZj7Rz/tBaJGQQ
3GH5OI2ltEtWuDa9EYBycVZRs/QTqKSLa5fZ6XK8ngHDaeu5j6EXp15aCzSugioM
+daP9htJUV2h6kFxGDCHj6E/R9QckV8xi3xK5xMC9k15uXigvmEuyPTJ8ogFGfLJ
AKA+85Y/aexKtadNxvtWNwZyD/x6P6US7ny/QgvpXm/n7ZaHYXQ6xAa9y3oufYKW
LByuu4o09UUg1MpfviAJLE4oeo8g3WOZuZD/+4ZnUyv7ueCUr295JHJC+/NGIHlT
DBzdofn9M7/HQd2upn1zfOazKidRVtXp2rGQSVyEX4zg9V+6u99/zLvW0J0cjg7F
C8qanOnyEt0MznE4zjm2lmqEMDqx72CTSaNAWnWsYLZO4qoanTPHmW+MJagaHxG0
J3DXCNhoVjO/XAYk9YMrB680yOl2fL1BgMxC30QoBi7hTKVUoorjnQtJjhFBHxQz
ZUtMmHWI1q5Zv/S+4ZNFTZiKjd77GQJGdcC4IZGl35pujtwL13igbYCaJoAen/r7
HMju2jhn5VZGYkFUtH16dUILfXEsjMFXo19PEFfM65s3lw6+eet2riz7c4gbJ05i
UVChEqAJvE1oXHdEQ06BeOnzQ659UcdLef7Qfn2ZKuXKmRb8lHLiY5wKxy5+4JJX
mLn43dYkNBG2pvuzrzrpKVmY8weLwWXyWTQJDIUEFAzyMz3bsDT49BZxYnMU8kuR
je/z7D5+gtz7eK04yv3PWLTHhuOOScGqyauwq+LWwMGf4HtAUk1cHHXUtGncMtX9
sXjpCNDa1JbEvRxn6lZt9e/Wx+zbSW47nsHIlWRev0N8k2Y2JUcmgTJLIvXObdnC
cS9VpkIm/09g6k86slj4Te1Hou37wfAhg+feVz/FH9/1dBqv5iKRnGnjCIne8Zs5
d0ch7Wmp4spJO/n8ayfFZ1sUXNSCwhLsnd76aJFGM2QHATEOjHz/XndIdJFz1MAr
Mpn0so8B2uSEOTwCb70xV5rv3shcNxbAmF1R9MFJgqyrglltjv6MwtGRVdrgnXIt
FQlyf85jZUKm6LHJCHrj7ek/O7c6iergIddZhKwmjhZvQYvCFdHV4gRiKKyAhpCR
+iI6LilfDaVmFwJ39NLCIGwuAZ37myiEIPOfX4+aA5nf9t0XL3+7VuSa6k/eeTfj
Pluw3z5Lr0ymF9v7kuc0EoxwEJAmVFY/g1rHiBKEDxEh3seYQ0znixONDkaV1KVc
ZkKk6oFmlYZkrVlEac2mCpax+k4wED4G3HBoX7Rit6k0PVEair7PtFeM50dW1HYB
pgkUE0KTmVae65Gb531ifdYfD6+tsPwIApuLZV2SrdGv4sf4tPua8Sf4dd5E/z/r
/jK5ASgqJ5eBS9HRBANGsRJofa3yNriK3Aigby8GYGaO27plj8wSrgdllibGsW52
7g+q1r8/iCgbWxn3toIJKcujyxArCkMPHx7/rUxgWXklI5x2wTAKFmcG8pbOKNgg
aSmPj9ICz6UQ1NennbCeS6MWEHILcXPFrGo3yvmXS9qpNroGEfiLgAFGXI/UpNab
eTsfNyqyR+0og0gj0fCDGFEGus0CCncN+0Mye94TbtFqmIMV+a/XlkwnDVOv5hYV
YJszijSZk5wxsVkIZatVLDgJZXAZQPZxusth9ziKiGod3KC4DUfE0XBN9rxw8OPI
sg0RFJXk7EpwCizXKwABzHCGEXY7mui/FxTZvEffzphSe5cNWm2qXp/fgw7W+4g4
T3VXSTFzfJwjp/aKJZW0zh9YTKjyhluc6plqt68hpz2ACExONZ2FrVs8aNUPg0Tl
sflKrocBEMUs9byGL0dd6cDE/WcmygekP6Vd8l9L0N/G37S/PRr5ReBKGJkbv/Gg
dGMoYrHNvfGDpiWKli4EF4S7q5+Nt2/hMhMWPwhkmCcW8xvEtCQ6JZO9W1B6NKbH
t36p/3UOG58VUn2zEdpNjki2XPYic1Z6+5QYfkgiqZHo9uC0yCWfgGJF0BYLXFKM
dUwot/sbAmSFiic9j15GlGl00rZoMMEUBshex2vbRcsuIX0u6oR3hUBGbhMQZXDm
SRbftdseTz2LeaxFP0Hf4vA49A5e8kVK0R3hPMhtf3LDi5YZEPNsJh5+ifM4Uj+d
HNFg1zVIkFkBHxHsHVKtlvlQ2D95c79d1eL8ReiOFs3AfnMP2hdquQ9xZRKSLqBp
bv22LSyOOZUja5DwkW5U3WaqtSpf8Lna+fI96ovDdCrycwhx2ONaEdJKxrBY3HMI
GcL7FRfhYjqud2/O4AI/H7w196CZtblrCOqyvo8+a9sp/+nRjHxmcPiFMjhsGbHp
nuv6q+IcdT+ks/4GsAbW5uH4sZl41Sj0XVgPeWmkvZUMEu73PlcGO7fKTZwyBl1b
w2X0wfLn/Fq7l5en5a9vIfB/ipZLYu2diqUQzkKGl4o+hyxCUH7u0dw4NbaCp6Bx
UqoU9fsOEypOaUGQmkH5C78m7ey4rV8yEVDAh1IgOPqb8TzkoEA68LnSTK3Zb2hM
r9KQ24jXfKr9o8/VVxhbe1NZFPyx5RG+kP9xMN7uIrWrc9DAB9AO7PaYyAil42j/
aVEQwKMtJI1Vso8KdvlN8LLUdZtdRtYnMzzj6dsHj+0jdEjc7qxuIPjd2sFEl21h
vw+v3Xc2eQwc+V/DU8SS7YSFnSQQEwev7rgTCAE0TgGw8qQ3Vpy9+QowoC8E3GG6
DO5g3R9VE8SS/T/wvlH5hpnNf1vqtYRagihSoSsq94nVMLhZtm3W+6YuUB+uUgPw
D2EMxeETzzDRfnLjWEuzXiY2VB1BPvzaeLbJV88mWNL/H/cdGbUmHO44f3YTuHs2
CzYCQ9ZTwruNLY4hCBoBEQrGyk40fmWqs0lg7YVakjinpBwWeSdc7WEogRrpIq/p
IVhJl2AkwXRmSmM7QOHm19zpnFiMZOjv/wAN/52cebT3kC7vjHys0b6N/Lc1RO0S
8Hc5pp+fxlVfAwqYsBpKx1zCUaS3DI64T9l1bvodJ1Jaw5K7NjD4MiYxl3sUit+M
NUYrN8w2sr3d3lsM+wOEbJUTb8+GZGlyP417mLmfr4Inai8PEr+DmFX+8tvvcdVL
Bb+EypVdEY4dbNtblfBofVfiIqAEa+YbIQ3B0grATCiUCQtHhQmU0IdYTwSK5uVM
96jeaYcvulKqBtRJOVXGts0TzJfHAz1O77ff8yCFSch1ro5HA743osnHAku0clvz
x5L2s90KB7BrInD7riadqizSVql3EeQ+ojaCvTQ1MFnZFgtFgAWyHryOI27/sjL9
RMU4KR//f+rHGyJujJpeQSTcKhxv2SwG0M4z6W+ilxHRRpSo4Ki5yGxKM/2eisfR
i15XzoDc3ObmUddpMSxPWj246aQTnsYEEiKLUJNwytJZIWSOnntXASk1oLDqXi2U
PiJ6lqAqaHXtZWFZwASIN396Vp80umUhk2NhIeClwV4xttsE7caxAP7jS5r0vGNy
QDPEZQ7KMCCekBcZp0GokQUo0npecwCQ/O5Kcz6EUd4Ob0wrD9fUenrN2aLi38nL
WrpWZ07WqphfAMIan2WPxbpnP9K4NrGYpAFt5ODGg7iIhdULQiuXbLst5su/TbOa
FVP5B4uJ1E9mbQfFzqQC2gOaaLhPOhImJatRXckQN0FFUUkfdkLZXbKtlshSFuNM
K80iQQN1H+Y05rYa7XcLXt3anxEO6UrUcB79U4bwuCDKyKbBGYXRo1xXhD9qTQCk
pXogDBIZKxmzNDgEJRA7BtDb+o7dSh88LmBE+8paVOq2Kpayh7odp/plK2byOZbL
C9qQcPDHtxkL4fH8Yx4fq9r8W3c/wgMGkwiMNbwqK9vkaMNzVv7CPlPART8iJjoC
TFXFdb8hkYvxhpYNd5kNdHxCnb/fqa2XmUML0JJRX9HUmcduzTR4vlNb5lgecyeV
FQZaVMRDpyvvLxILruX8shT3abpMNST62umakmE/64beRct71ClyKcMaRzQnSWXB
zg/7PWs2MIRCi7M/endJuIrdsGq9tR3Qfc/G446pV4V6hDq3HJzN8w/LTHGGX9e8
+cW0vziOiKKUJNN5H/GMT/iOOZM+BMECxlTbYqiEijbVLoT81eEg7JcK5o4Sv+Dt
79mJKTJsLfNZdTLidWZ//WsMkyk3R5zciOZZpUA0dbbXZXo139Kdu/EOUCJfFtgl
2JUa7b0+N8lU3dN3qDG6rqQqGH95uy8qaEzxQeIUg+OOm86CmOKeie0LOjhzusRt
0TZit3YqtAxZVtk9uwPEMUHAVGfiFaue5/xfpGm7F3mv2SIJPa7XIoYbk7XSaYUT
/8gX6kul9BQ5cuvxLupXtjysURne49vGEiAECea6cZhwVAwJ6Xo1hCqMVZeDGhE9
zxQRyAYN0V9aIqWWlQeZNH2RpF6XfP4TB9xKYzB3QDmdGv1akaH3Uk3uZTAfqdVs
MynPek+miv/5p39Y+MV6qML/e1OXbTkBukkrFEw8e1nWQwePJ9+xcHAeTmkgtmIo
ktnYdJrEAmI1rmP/Rc1GALXaWCSDH2Tc7JuSl+hxlSs1EJpanGyYUKz3cJLsv4T8
OP3PFdrKboqjf1JB/QCT/ABTQ6NXOx1DdKk1pyi9YZ+UPO/eBbA5T07g9X3KdDK0
zS8M++JINT30CzVDCJikuiBBnYe2QhJTQpv1wdSYPt3NK4Q8DE+CNWf8v2xtmq9M
g/5eJdbHn+ND1IqyaILJD4uLKdl3yQFGDAdP864OeQkponDZL5fCKhHEqdxxFtmZ
Gco0XKRr8s3W0y61dx3+p9tDqWapo6gXT4lE6abzs/V2qmZDfiNtOGPAT01L6jUW
LEmOHNs+9EbfEjJTaUuBxzTv6lNCvat5jmYfQChhwotksD3OWO+fXs095ML1Se1E
1rYCH1pMn8VYq9W6qeigGwYOfRKC77wVXQkIHJLfC/oD775NRMy94CxuDLdhrA7J
Ge6Xm3eOsPfO9Fy1xY3SwYRgjoCE8VYcYz6qt5kj07Tpmjw5402DzBbJWe1eAkux
8aZw3u6FsOmpMc8C9dnKQkE0tUUn3OB+4LPxkdYNqtQeHL0immiPgcDLJgENC/fw
VFd/27XbPwbvfXV8cUVxgbT+iw933WqwZxkt1dvwn9cuFDRimVhAF/Pu8AoUrjxN
LtU/I+AsNkqnecp5M//DqLTEReQc5f9u7DPz69pzmaffRZKilTw+dNc1YGv8r/aJ
Pm0GEEE+6k6oFfUBNdhlXf7QekVV4oEAtu7Gj2BDvDjv94cxAa+MAlKydHfmq1QM
pAEsMSel/EaxtTPIUl9HHOdOjoySG0J/KoISloqKq3ixfMID8AnYDGF8yBg8rbQS
Gr7Uf0bwzWF/DGUxvqZiwZJfj1Frh2d+kr+x61RIVy4/ZKhMMBzhDDrUD5ixA3Hg
ODbuyR/MHuE/h4TxpXSbnjYXhZ1xMntUvK51sHcDLg9TSpMfsHOGjwZPtyvkOSBD
RR9k17wAmC3OFi007hUeikqZ5Rx+bQjT9LCMoK0nKMK+bSg1uvCcFI4tr3J8IyIt
59ijUmXNl/hzbfqxklX9JH0k8+gJEbeCi2zuL5pdltxP0aHyYhpdcPuZ/5XxUerV
Jxz+xtN1ySV7grZUPApmijXcbZ1mNZunAxY9+7BrkqscpAtHiepaYbrp9VzdzOtd
wdWDusMYDdIcy95/jPr/dqyAf+fTa6PnYS7NPFBK9VWa5gp1EN4QW65ixnbDr15z
u8g/Tl7bAsA5MlpbKCM792nxGG0fTzoxv9SEmn/iGzbJheTTzAUO70JaFTJVLV0W
G0DeQWpHU67v/fcLtJCx+dPdTn0a/6aBNdktfucfQIyDa3Kx9OqSkIprcD6E3WnX
OTSbZZB/S0JkXwxRsRMnK65x5gZ02DWvvlfjQeAHN1eU8MQ1v9oa/eG/yQWzrx/R
TPxfmpUPZe/0kK2QSb3KOJAILvhqe1oiQKahdIQsUPTvQjthl1yyFEXRAHSest1v
QI8VY/t3lp0Cra2KvAthC1SmOgq4SSmJ/WxNxjrtbuZE5R3G4igFYHWNDugk2zNL
3ZDU8cQTKp7tktV2Z+Y4LnsbEgci9zMfhpy8QT42yrH0mcTDGpHgdMt8dlwy/M4X
W0ABXEEsWwUhfXb40ET0FbReCjH/8jWI/oe5psT5ujyH/MgXmbjcOOLIHSdRjx4+
dfFoTl0ODrwMBf1eymLiuPYG3+CTj7w2snwBC/CvFYpNi7r7X44ZyQ//i5sflJOs
q2slgFN7FMOg/9q3jDx8vc1vflk2gCS89pEKJTrBFca6rtHflHRI78PS2VBdbPrE
ZQ6+NK5hI3++2phN2XCv+6DuvgMTOVcxhTvc2LQgJPyiDPCqhvYCe3StEFtercVJ
ejkHYkjrEgsjfLOlt8CntR0IBRIPo76r9VWkMcqQPykWQhTK3DNoLvu8yAQpe1zU
tYuSvs9DjXamGFGlQWTGbFXg9Cj2FQn3O9wX/jq+bKjfNNjLcbnMZWiejfJd3Jek
TUvaXCzZcrsUre6npKIXprAhQU3ag6KL5RfXaHW+AVSqwTwGqGJuD14RRrI7FITv
hRKpbEIKUQbznkf7Krls5hqQvpoooYSPzOBb/z27/lr92Gqz3WUVj9UdLeX9gyNy
7FG9px7U92am/GK7aXxVuaKnoluFh508a+0HbcrOJHq/BqCf/IZCZpUPlarqQgJ7
7Zjv4duURj94/tZ0CFb6eDR/5DbEhpoXApH0ILov7wo0wZgT5SX36k1nk9Pjmyfl
30jk/m2NYQUZYyl7FK/p53U2DFhjUQI0+lURldJTQHLmjJwgsmCeqYjn5LF8fWSi
2MsPEG0pR99kDFbJuHmxL+tV7bjt7M3PRQnrJzQffPxEnbohTM5F2l3yamwyUOb4
9HT84s0nPk+pYvJcaGdDQHhqMoF+9hd1UhnQWF7XO0jAcmCcbVxU/d6814VVgIta
W+zTpcw6JyVTfuMpVLl5ZW83F1cXwVJJ0lsXtDpPP134F3GT3Dt8Yz0O8cGUmODD
6qIOiJi6gqB0llLOwaKN2p6aILspyNMoC8GJ1d+ams0W9UJgEqp78x8sHib9uCuh
6RU0FQpOaWSSsizuq20iRrg8XTrqEdoOw7x5/cyXuirHHwhJX0hl7vYa2fVrZU5j
X3jVzpl47Y3+19N8Dt/BSUYJxY8YJo16xepfTqW+55B1ENt1SE5tIR7JdVxMXkIN
cLB1CnWptBj5PqY6/jqmFUMudXEYhCLsfg/zxrOC/zwtEj1wn+gvUiP8C9a9tX66
syaPIi2EpiV8e0Cyqt4jyBQCumV8AXmRBnzP2Y9jheDu6YvOnNCV9yUOPxewrFd9
41sIunPMAx75EW0+3zCC79XyX1pylfn8iR3NpoGdLbVeQ0B4CIwkQQ1dFA46wxaY
hku/6goL3wmUKah5FGzBjyzH1d2vKwEjuu3lZwNe06KlMdnYnfBMAGI71tZwd77E
cQvRf0DEvB15pmqlHz7eC4P0goye7E6mQMkCRT4HWNFoCGZBoMIWbrkhlxG22V9Z
OnYtbzEHYjwhF0I8CYHknsOZcwPOHzYzkT1kxGqXl1RAgDDP0QAVrutVB9+xzp8N
3khe4LlG6rvuvWSWuys2xEeQaBJ5xz/tU8Qfj5Cmqvl71UrOL4xwH7Uz3ob/3TiJ
FxeQJEyFeYnRV2Smmww3CqDjGxthK67NSagilhiIuRIFh7Mdv77uDw5xc9M3EuSi
5MDTBZrOqj8nrlRJvumtbR6koWElQJPWceCypPB5NMfsvgBPKU093oZqaw2K1maR
B756rCbDl9GKE66f0x73+HnaYHkFjvsAUg9XJrNFXqtZBapFGWEpXrZFJle6jTDB
k+5Q1ZfBpdX640JuxRqqsQnmK6OyuPzhRCf5J/hBAYLapIpwdnD2lePU3ddapqZz
PN2gKMbtc0OQPH0omAUbnVcqW5zKTFvbwSqg7qbeE7xdMAGea2tNbCmU/H5h+ufr
pkcy8fnwZh9FPFtq1sQGDly+6COZqFL8LECNc2VaWEGc5s9D6fMxDSBByI5pbrKp
hr0DHl8GogC083SSrRaUJownOrnz0MwxnKfINGY6RzuCorgx7kg7bND8+nB87+Gk
jNouys9a8eBxSAGCPMpjsfpqgmQuCfPDKO7gpoxfrHGQaZc/ABwwVPkVJ/NdKnoj
BwqAH3sJHljjwx5UCjwPpeBldr9WXFgYw9fLV6JBCybBXkmDy1rS75ofmMj6ksfS
e45jFz+kWoQAYZiDc6jHcQENUamZt5FyQGLSPa5pRTOylKMFFgyztxgztJO87HmG
m015GnEW5ITVOU5nw6yQLEudR25X3QS9CNqxZ/fE3KDHTO0Yn+kOkt7hAwnBlQPm
G79VsYSzJSKuwODvMAyBTKuLvQb6xu7EvDJf2afJubdMPyey3pTxHdQ29aiTo/Y7
9OPhIOU1z4tVFzmr+/z5qPbtiX4cajEnPZMVFRO6whUz/tT6hN2H8Gn9rFf+OhKJ
C+A0lo982IIx0Fk5/pAmsnjPhmaHZCb5kl795lI/3upLqdOQxXb+GjAcWD/hxVbz
Rl6lLoHLc4/Pc5dQYmOMUMiTSgdM9idC1Urq7U7BSUPd8D9UERd1gu96pSmKt9zE
xa80H6EE908Usz0BF1lsY+cHL1Q/Nm7mevtTPPrBeY+FTGAw82JkOH+AlRL083uU
4ZD9BaVdD4kPEGNosGiN6HoaOUnvT6KE7yBb0P6yMm0qHi80N41z3vILrQrS8OOZ
ymN+0IBfGBaacGdKDu6ifFscvIbPSDbhtI1BeiERxxj4YJ3IJEkHUwG8L30z+d5a
5rzv4QslT4xldGggFXRysdtTcI1COetGyKI8k+e11Iwk4QuZYyUTn+kGXH0O7b4f
/MEPs91rpyey4NlaVFVa32kJvVhgIVVGtwH8mQkgX2mPfJrKYapTZqzG5lpM/Q9l
0Lfc3i5qfISO4eS7oTeZCsfoXPbd84AaKnF77VUXq/IFVXNKcYlsEzBDMJbYQqa8
1RvKcDZ3EvQsxGfS9aPrVsy/N/DqIgI0peFXAPhpAraR+ETjCIQ7H/r7X+7WsdW6
0P4xoZx2CvEXlWXGvbmTH3HsZw8ToEseNM9CtqJW8/fJYjzrx+9BLLSkwZAJlltK
1sFAI8DaTkZPE7jPjK4IO+gMnuWSOr13tqh440cOvYm5389/fMIN6wO10BkZvKeY
JQOmky8kpGIT0nKlRClZg3U6gFuYJx7r4+jmp6dALHXi0N4MtzxGVTXRvhcX7Qfn
g+AhjGeBjqlUu/b+/osfvMMFftwXZPokCLS4lZWK80tYRF2YBVbrsQV2eOJlWx0Y
JmFFbpMsayUN4UghoAAe0eNdsvWMIeSXOgTB7hMXdEHiGQxTbFCtNgt/JlY+t/+b
TZ3B19/DCltX5qPPilQBAq69jpc1QlgeVwChdqV3t8VndtfIZQXRdTEvFeD6ADaS
N+BN+nfZd9J7nKjMamLFQ+SQll7FcH3Wl9ph0416mfBEv2KYsO8dN9cI1nFfdRAA
KEQIfUWM2M0oYKJy7PVHNWlmptOaAkai3Z3ddVNJerWIaKhh6/DxUf8qk6JIwDxp
HimSzpxE9VSJ8YXR2SwH78fThLFvJKp7ntIpu2N7t0DzuOkb6Lr+MAL2/K/ZIEVf
x3Aeww60C1mayKUWiZbD0nnVhjGqJgcEi+8ZUPno/RwAJVi6LxgWWEibe8HnKsqn
AdydjwCnv+doOmbdo85NGehFbtm3MQsQwb/Vt6okoCAtfvINf5N+Jb1XngqM7Spr
q2Bf/D21YFLS4RlL/hxv+gYa3SrqwOS0HV7b88n2BpK3+SscgWTuz2QM1RWwvOaQ
80P+3eWqGajlj5SQPewHAy7SXaTslAtwGgUaZHNGXl2GR6h/ebTzHri0v4K/5lFR
Eq6YTDjsENxQhmwUwBuFAkiwhNIbaIAdgAPgEzkavrXLCB4LStJ7NwvZSgfKiKFy
5zQk8kuLdQ1Tc7wy8LsdlvG0bx6QhaZx56PyAd6EdRruJETsnaYB/LwE+Du2WDxk
+kwTIVl3wADHdRNGzwBH4YGh7A1vFHSqCkkSY5Lz+VezD/5FAZReV4Hj+yUoR2XB
jxhQkjJfqVl/QooYFCA8gg+KALCYopZSjtG1ccaKlAlfubC8t/pUEYJdHJ0lrkr6
sXr7daFc9FuE3f1/nhagyQ1q+cGluW5MWB4PuDIZmXcz340D/wQmfwoslyuJPIwB
bu4tknN3M2nRFhCUKlj/ZUVsmf6ZRspDjmbu78QYFfauPcbaLhV7adxPCqQu9N6c
NdlUUmEezxV4V1tf1TzEZ/hIIbpUCRFPx/KU3GJw3rsSQ3rKTjrWdCJwciZzenj1
slwvFdmqdaH4nPIuYEY+ksp7jtIF3pH/fXx4Vf7aitHerH6EQkifpRV4VP3TmdPd
NJf6LNmfhe4q0Cd+sjF9elCqQK6migVEvs3uGMP4iEWUeegSbyjumB+H2Go9zCmR
uBTTXPkX56xm8Y3V134o7iwYhQzVCy6H2Mi0kl2kRNOZbuVNy5fNNtXSP0AZ3f9S
itBgAQ5wjoz1P9tO4j3nkeJqs3uixgoii9xRMOjWn9YpGwZKIq9AeWxwcf6RcbBj
93bqjOf4wvOA43FScFg/B2RLVsHSc75762AbKpfDY2Ce+qlHUpGbFpEbYwrha3YR
zjt7rUvsf1SUi00gl/qI57jFwNhmXUO4sBd3Z2VlPCbUCxiZ1jq1GL36oD9R9CdJ
ildaZj9nF4aP6eWkdE6AdbXPTlCn/ijI7WgAX9Cs83wSKb6K1ux4G60z9AYoZUJP
4BAoEsmXVy8UOm0gsXOGOdMRgsIBvwD5sfwUvcHkA+JP0iA/lgPzjCLb7ZeL779R
T9wVFSuQ1sDlOdPbW+XPtq7mtk0Yf/dd1Qcg3mWxVNPBFBuq0gTuN9IWw17nrAjF
5NkXXVjmtZb6vkJ46bGsMZYjYBXzZUnG8hWrB6gQjzySGKqruhkts1nEsr5ZvOQf
Dkc7MD1EK/QngfEQbut2lY3kflRlI1DyU/YISzknIoYBnQ6MV08K8QW/0nbFjPEK
PM4aSv2rCRBghnOd04LoXVh8fDer65IwuwiaZpjhKfNWIXcPXBhAF/WO8KH3Oxsy
eFnajsUX4ayHh5C90N2wEbNvouxL9dx8U9IGRnhSjqbX91vI/zoTnPCmDrhiP1EM
bj2MO0CML2FDSIrlbDjim5DgKG4NL60d8INboFt0yYyLkoFGSmhWyuKYlELDOCsa
vVS5DxJoPwSF853olYvUWxohSHs2CRyBYDE5rXbXNMEAYG79FHQPJ3yVwbtr+KNt
AoPWKIU/+/6sYIcebXfTkSSx9qek0qP50ohYGqqCrROdSQBwOIEDS5ZLlGCZVlqI
eJ2rfD64prpB+ivW+/Mm0esf7JlzYfrcBNlQ6FkckPxMNy3Kim3HQ7oM8hJ/YQ6S
OKw4iTwis0F3OvdhhFwvUdRgev7cZDTdc3odexiBpM+iO9SGIMk4yUTPWtdTEjr2
RxAJMRpsVyPCUFhOjaL9iYz9y6Kz/JrHxmlS3viKZyaCR/NJpvy7rvd6mRLKEh+p
V3C4i1qJbi983j5QLu+89UkxiUc3SYMPVbZ55BpKQIEG2eHVI8PciMEGLQBeIEOf
c2dGCYR2ZQX9bswzNQQWY7gtJ7egikxtzR8dggJlUmJ+DivC+Yxl0ADu/mSP0zHi
7nIPdvlV7D+VLvzWbAMEwFg5O4R2bdBw0v7tNjwvvaF1lNVWfjgWcd76Y+o0OTNv
8Pui7fi7mSzl7vlWAlfSodiKO+aJlzV0gSKEUf3Sk0/ztitpVjorXnFkGq0Iwu9o
VlRc9fDPNKvXX4xa7STHVEGsgT0XvtoPHeVkvOMCAYRWNJnhFq6nzUCM26tBeWFT
47rmnbmKKNW5VRlOaFnWAr0X62X6vRSqbr65CLxH1FcHg0qG56X2uwP+Q8e5v5kU
Uqw5zsQI17uoTQv5+UlFO5WiTLTZ26/ISJKXMyn+dzUDMzh3HaT4/vxQsL8QjewZ
4164mP5t0teON3XiQffaLw3GmvQaqERkPaLqvg+eBOKDURAlR2JUx2/0G4LOmpNL
+tMF4B/JFTYxUvpB6yzreMW+q1niWACxUwmGn6rVY2yNzpovGWOVjkzsJU+9OCm9
L6EcsVpPsFWW1mbu7zIvLN6qzKqn5fX/WsSBAq3RPEtqomjuGSDcv1aYgAaF3pJV
W9xZO6WXc6jbf/jnkt+AhZR38Yn1sZfvboqqxEt4Df4RGv9lvAHpEl57CpFI3+nZ
WI98Gqo6XZifJOHXbfKQB6wktum1D/L5ocjjvXGGUXEHX+CPzckQKX6wPiXndiUd
qmcMu7YcTTM6Fk0dQntqgXSxAPUOzKjCT67TGD/L/hiQpTznNejDCFZCTyR9H5gh
tWzWRCTBKNc1aYDF/ym6jbG102Yd6NfULd8ieCIquG80Lji28/XrDPC8pso/7aNy
tMFcQgcT1UBRUt2hnRXRlrVXL+cHfkBBBKugY6XMpeD9g04y6f3hBCPfANG7arSn
99VCmjcVKXK1tqHA6Ti3+RYKZ+PjHgALfpgNYj/caIQabkjjahtvfoYYyH2zd92y
sJrrGo6iFrdOItTCkxHeaUr/waHsa3AepUthbFWibi28OH2wuOsHtjk2ECyb4nwV
MKxn5A6GcbpEDL3lSaTO3WStO+LbS+CSU0faY9Vzt/OXkil8k3IpWBPL04uN0fsP
8A3gMyMYYEXAZY70oQOM/88zYOWNJripZrv2jZTyrKWWjpN+q5qP7Yr6+NDDpNgb
KpdadsSTXYlBfy0aD/eZvyp9OYotFYSuaI3gzzBeigJtzT0/Yttg9pQY6GBJDmtc
BmAjBP8IRcw10/9zRx053bwwvCUf/jx926kdkij7cr7RQEr4zYammyZBk3LQIQB6
JYiFnz9Zoic1IAU5Aub1nhBfKBwgeDyFOCiQMFeokHzHXK9PM/5qGIwOMZ0B7TZ0
7PYamKrEYe/1DVOj98eExnP44ic3nQmL8X2pWBVlJvWbCviUc4/eVL88pNyPsBKJ
fTwbfEV66wPxfWUt8UZdE9U39y9tS7bCZVtJInfHErtKIXE+MU93Q/yt0aepcNfd
fxebMQGYrwvrhH2P3XYSb3ZmQYnN+uB+0sB/ojSZe0jRJ4Si0/cpNtE5VtbgBLhO
bK/tMjVDKaki+Bs7TVSfoW3e72OPy3b884qOftetIew2uyvTh1cyp4xoUtvUkqN9
rMvIZKseSHNtZz42HyHF9Wxf99SCchPz7RrO1OmZU2qVcSDSpGJnJUW0m6sQTzb+
T9Abh+2ffYF+OcdoZLTeJ0tEZO7JDVrv8AD6XIuKIOMlN2Xuz3eeqeOficZF0TBe
T/Dwxl6rqrBNLJ8NlxhC3w==
`protect end_protected
