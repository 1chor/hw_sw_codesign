-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
mRnyPfZUF2+jaBGTMnNIv7CMNLvKhGRRvrfKHIFS2HFVh6e2Ubh/PgBJ2aOl7uqb
ZiJW2B3IWhVUqyndJ6hw4+6tqu24aEne0Baj83GduMA1ntHGg/FnmAlFazcCG5tH
gcQiVK+F7AncpP8hy46buA3lisg6uvQ8p1aeQlY5c/Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10336)
`protect data_block
2AohZ2Lwn2ixkN419/jzy5F0j3fiiLzErVew1sH+LDb4T41zbPWVQT4TemB762jz
d0voH3jKzMPGM9LOenOxzTKfMJXHyj2ZSiYHr40OqLPA5C0TTBF9rq1xKoCDBHeY
fopmxSd5QFK8vNBW9mzI12KRZrihanJNs3aGDTE2Bgp62RM4ZBlb1iFBGKnOmCwY
T4CT8kmhe4wJ+Yog2T0n+AzNbv3tzis0FZBv8MdjQdaH7E7l/vTE7H8sBLL2Dcmh
E9UtWqciJs9r0THJclldFymwwvb9nsnzA5yqAlKt48uAs3lWmuRYjYxYgvXAozpq
50wQMUfA7U4oH8cELZz0geLbXCe8ntJsCY5ULIH0cJEYJ7WhA/m5TBOi1jI8ofe+
n+beYUBucEcR/U6EIqPMmLE9aGxp00/OrqD+kEup7sxCoLx8Y7HIw6IudrgAg80s
KVmHSs89Unc0hhQnDDMo8Z2fPGeIo4LVDc97mxNSQ67T2xfqfj4TuMiHvaQaskRm
QhEOJWm8IewgDXkubpmwjy8URh7MStOYJgqvmB+BgXTgCwM+mgUg205Gb01WOS5H
UHpp+SE2mqpearZ/c2I7vWu+VepzZD6fqosXQMVUDPzQbiR5iZltX0uiISGJrw7x
i658BMy1WYC6mxTPVn19C4M/e/ZGhhDnmYJl6sSpiNrVSYlLJHdwwPgI7OVy+Wce
LYGNF7A6WWISzUTqERLS+EZFBmmT0wqfvKLtYkV9iuJ5KwH90gL/1euqGjsRB3Qe
eDhZCnAMs5ugsl0+lQ4Iq5Ykr3Kv6MJXELBGE2RJGKEGBxMgbEnoaPar1IHdurUK
Ik7tcIpKd0v5bWQOVMcToGlWsX0dgnhfBU4+HQbFGJziIH3/UStrW/YN3b8xkX4z
647rmAi/8D723kk9SYNTJKzVvxVoJXcF0xgbbavXtexdR2ZDIH51BkP1XOk8BvV8
JaIBPVID0A+fxgVqLul8OqQMYkBBqTDjMbxB5ThPInhEj1Ewip5t6AES/u68YOGd
y8GGlS5JD4sB7jY9mPC0RH9jMtqq2em8pbRYId1B7N/CtXTUeGLpJRdnMOwuNCpb
yYLg/xye1AtJv40xCN3suOiIuz5I/TQanmgAEtXsQ0Qt97QX5xz7ZfxjDKTmHo+9
Va/p5xVq6JOATWLgJUcnIWaYFWiu047y2Dsl4jV7bTzoppGaQG+UAx4RhyoUytrr
Acs4K7sm1yb4hL234fgK4G6hr9KD1toQUYYiO0I8Ku5vOJcAoNrrOdkgDlZbmbYv
Y4OMPFkpBrh264AIbeOy0mImdXzF7UCRbUJYCR88Tx5vbaH9C8C3LV7zYmkbdtFn
C/UpMVKcpyw+8hBqSdahiHpvCuJxTP38rRUA2m78b6T9chTqiqvuHq1pqkCw4vU4
t9+0acfHNiZYINiDa1GP1xZXgUYqs296hNcYb7uUOmsaBWHNlKebziP3O1nAGxMP
/HQE8/Mn+c46KSUPu+yfmFwA6hwbTGiJlrSkD+j521P9rNzH46viy/9omr2I9QFt
p/IbxrcFy72vukZ/kDGrYn7boMV0YPbT101sA2slmU39oS93QhmFwCRz9Yp8lo3w
H6pPsNu7yU0DBfY0tXET2G7KVLQFozDL7nMJZ+GhmwquH0s+8lgXSICe31i4mZcn
VZoGSSz7Rvj8BBUspIETbiUtJBC7vMFX9t5X2f0a6Xhagg7nc2fGKyTWBaJKsJTg
75FO5Cpr1bZBM+iNONJgME3YgaqOC+wZEiOa/v3EgOfMDflWzgvwHzeGSlVkQMZ7
rqfiDxVgyffVrgmNr4a3Txujwp4NrqRt3/zBmnY9MaMd2Sx5n6kp2ZiZHr8qMjlH
8RKmFFTpmZXI+k033XpNRWqcdmlllYoDsc/Ucly27OzBb0glYm9oQpaYovgUB7N9
MMUCc1dfSwtryOqGhHlHjTAsQIOVpJc6tACcgaPnc1TR5K42HUdOE6RSvtvOnKd6
Vk+g4CglGnYx178BFrYlWCCuvq4lGZW18xGxu/jodaUSOlTDqvd9YSYxipSpgTM6
sD4sun3sA8mCFKqL3fuQSktJvnKZm7WPctvP2Db59hjc0Mv7BtxJREA+AAStu4l0
bb8xaSz0mMrmswzrmMvEj3ioJ0FxY9W3TR4gBNBsNNi1j9sfihfeLvxtabqXeVqu
OpGEQ9uYEQEugEQXy4LuKGTdZlLE4Pyje52yBBacq2gzEo06tPR2nif1za82decz
vSXHnDTFHsXyX7GhyT0tCkbocT32jpbQBo/uWBp9otxz7XZ4saFGj3QVTiE+htdT
UX2/ovtq1mgLyXfW9VCdbAmyb58AZaxYsXxEIjrc1mW5XvIHmXIMGS1YXEHF3hb4
vCycKNmiBPRTq+jukUT9WFn8fi18a3kNTGbZF1qBRXkKmqX+BcGWahuE7Aq6E6lR
bjdRTZ4H4Waxg5++zYXa+L60H9Z76nkJBA64SraOhJ/BNCIq4SDHuumgZZ31zLhR
hHYAt9t98M5GpELCZjw722F8W96etVtzA/qwft1Wik806po0pP+7ey5t/uDwo78N
nT7vqMNgEc873ZxwIxmlxXB4JxRq2DrmzWZG4V3r7NmTKRs7TGSXyXrHhouvA3cg
NSdvOLb7xLbx/PZR5cr5QBSi8hffPqaJGmrzpgbI0orl2kuXDl2fjbU2VNnkuAiw
IpRmQcq7JMG4QDc13O+wmC6LdRWdHwScoLPYC7UcSUOU5wxMKSDEhT+pfkEL3T1e
NXDibC/8VtOJvXsVwmoKXv9EqEUTE45gsc6eRjbvWvBp536BCyimcKsGDfO+jlYU
p7/yQp5gxsHkm2fzeX4c0y6phgtpuQ3BHBjBXzWhV8HS8OVXncLJMvCqclrWY7Ge
RMk+BCSk1BgmFTNOwBm1+X3POF7rkkX84/DIJJSJYBK1oi4j2bhlA80gxYFmwtsm
qs/ARuFnbQSJGOgBSvyebqksmvPRLpFjB8aVE79n/YePL9d9FKD0jCAqs5GURkyP
x9pIAAREjesOiDVQo8rQrKvtxoEqZZQSOFM0GLlup+YU4gB/IyuiNcQVmtogubO+
IannU1U53ucMq/F4KXgO2SVzKjRXttFAFEktnLgwLFfLX68rEgHGYLSe1WJbk5ec
fH8eLbh6hl+jWBQvVLUZtbIBt/wV/grqybIB9Vr5Xo805bPOZGTdZmz97b1MPLiI
phAnACcaRHtas5UeJI1KgRshmLoUY5oqSn+VvnWfslWEk6JUs8VlHL9yVFQcFxr7
aXfo9bzGqkYxw7fhqkfDN0Q2MhCCx+IEj7vYqHJlcrvB7WETF66JZunR+UauKImY
1BIHX0c234ADhqmrvGIz7C03lO1ZTFpRDe9jSXkTR176rqEjjbSQ7onWLAkfsWM5
jwBbyu3o1NjzFQ8qGkY65GaUH5J/2MpQllbJ2qOlQfzNiK9MKdyv1udm/1uV1cO1
FW2gtndiyZR/8fA36henzc4NGuIfbDnSnqA1Txv8eilRH0UxI1RP7HHbtGpHLS0k
pRK8kIQdOUKSuBfcN8pzaLZ9qVhJ1fE+sXl6Wdv2PkiAEQBtcjvH7EJdpPdGcc1y
5jhdOT9fY1+c5UMMEw+segzev3nIGutiKs1MQWK1cLb/WhNkSY+l3hcrTctciU4G
awJt6A8XJLymetByCccaVm8rAwLugnkiUhh7UJ6ivUZX8ttAEqfv8QqEVtby5N1j
lZ3QbPshOZW6Tu2ebzXVRs8jAVCNMe3SyKynn9L2viVwKSNbyiNtpLKEixyCI0FE
j5EZsWF0tDVc8t77u51MJrVrDCesjSKKG4xZC4yaEV2Qzk1MDO1LB6NXqI7W4kn9
JcUH7TrmuvKcCg3tZdlv/7h10NBS45A6RzoKt0VkpRakdXJZBWeIPVKMgfINVaZu
UssrKr6/R65O8VJXzhHpEW0wUAVrZ9uaTm0G1U0lxMGhMsaXk31yJYJCGmd1CmfC
UyKazKubpKjhD3Qh5oFfOwbOgAtZLjNk+4vg+wyAEk7V4DF6Pjbs30XXCSyA10AN
sy3o51dBVDHTgVvH8ISPQIDPA5T7jNWRkqIX5brngkhPHKsFN87zfrcx5dTf06Ur
SdzgcZCXuX+qGzRSSfYVdk0pz/HU6Ps30AMH1k3Hs7xqjjOg6IiEUxMWMmE38NJ6
WxCsSoUnFOptDXbyPOcv1js+H0EIY7aVOiajbdGfo7BZowHN8OHKHBad+NsheqOf
tG4J5ypYxI98VEnbRezOpTMqijzZFakhVAaHJWX/EUwalEQU3JkiZmFbVDJUYAyL
Lquxzhnork3jcRxtDmKFsFbRUbDqdUr6aK0I/8y1Su9B2MbB5eqixaZIiglvCW8a
V4k8HwcLk6ZphtUzWbQjiluNfF8qpQynP4B3txlw79adhZIqEXU02jzWW7784V19
kp42Omt1kyKaXquY3cCBjFFAEMYVWbUai6LNYaw1r9z6fx7YTmcgtZvUGlp3UY29
wKba5RcFZMxSQdrF1tfositLBqHSIlLPEAOxJc7W2CV7gpDDMdxmRdwdJcDH/ZYR
K+5X1oxyXNTkFGd4VzEjlvoXafO964VW2VOoZ9VHKoqNRhMMlWJQrDI5zYAmF3xt
683AVFMvdKrNii9M7Zp7hyCMoyAH0+CcvNAOWYCODcVBt2BPlL5vRjTOqq5hLK1c
/wRVFkBpADYoeC4Zc/bHnUttROnaak52gpnTRo59KqjYBKkLsORbpUY8IkP72KeE
QKuq9E8Y6atXVuYiSSzny63p9AZTmNri973Jx3WhtnHCf/ulEuPVIV9/3p4KFXaI
0BuLM9RduUuB0ZYJdc8MWYPD/qarz0iHyL20oP17l/3KfV+mTAc4WgLaf91N6CLu
FM5t3B/BDbC7+3hEcrEfpdjCPOrEeELv0uA73Mae2BCQyzpDXP0b0K0De3F48uHo
a8wyQDURnFlrKvJqTgsHCZLa68OXPLcI9vsd1oAesi1pidV7BebjpHu/Xe2cl//k
GhH7q0nZPywJY5q66r3A72Z/c/pr8SGkHmiXy2AZ8H/fiBd8Tw1YMUo77fEkUTy3
q2IdfTQj3TH5wV8EIbANDEybIPtp9Uw55kcXa0t+ElUpiR3i0gHmxjsLi80Zx3md
PfRIfd17Vgq9M+5O1pcJ3U13TCZVwMAmz/IylN/FeeoRCLwO07cUx2G3bzOSkg7Y
jPYK+X9Y7dTevdlgD4wN/l1NKA/E5WQ0sYoXGH17MfMWuiJrFp48GfZ7DfZnz4Nt
0g+CoPe5X2X3bl6Egin8Wo9vUu2cQ1pAbJpZG3Ob80da2gkVJpHrJGSET6e9sDlL
r+r8NcLMOxbVcG0m72pDMBopq9J4I8R+Rr+csmTQmQ9DnJTtuJ8XDOKfImFRZsgL
byBFJYDN6msRnvcHykW1eGbxEvZ2Bo7UnGV1b+s4FYX0hDYA6hHpLak2yIS2AXkp
qtD2aEuvvRS9Mpt07e0WXiL72ajfje/KkJxSoOIaB/NcIFcbXRHJtdDOoAAFoTVM
Z0RtnVOfGLowrjWA3NxukIf8szKzhP63dQDgQFFmDV/7NHsbNj/9w+KPVXW3998i
fGS4v1jEx9ppUYIEBcoe0LdPxvMnXLr+M+dtGSpVr3l4dH4G2JTmXe8WDS2+BSeB
33MQmi70AmuslznyRuF+AlSQyBZ+va5+22OEqR0filHc0hQ9b0rI/B1OjiqpQn6o
+C8wHRcADDOHqQTzsAnz7cEPHiN9UqiaVpK8Uj7ZVyd5wEMJAPUOO35wDhvu+nm3
L8XU/v7cb3V162alkMadNw+fKeXTnzErOgjGK7INBuwgEeRm8SXynyzkH3PaAz15
a0ooUjj/D44ONYvDvDIWwJUCji7Jrw3/iVUp3dzhfvKg4F7zqBIpFY61WkLSdfsR
skBsyiDPrOCKMps4bnoNKAqOJR+SuhYqqdXdmEz9LyjUOytbHjGv+mt74JIgd+rl
QF8vsmH+7BVX8spE6iAa5AS6R5XqpdS5PgmkyyomYrckiAf6foah7Ib2+TX6TTz6
OQLxRY+nfU7ihKz6+JHylMitljaXSJjg89QsBV0YeB4xrLi5BJJpCaG+oBYwNMlC
4s3t5TFuxiShbkeM/4G2uonZ46qwBZPBpYRBut1RbUa85iOlKHFBHc6m2TVqzQ+2
KWBw23h8H7R7BchBpzrb2yzM+pxzwBUqOJU4I2s8ibLR/g1WQx2XmEUwgKvgt5gS
+FHXidVwUVxVg4ojf2UkAVDb556OulD12mzoZkQFp/vjCACme217VuzPhQ/YDq+T
Aj4fx/ytb2bqXqnc0g1ZHxWcK2kbhadHXEY1mimd4F+t55EUelF9xuroe8e+kgAd
1TbKKuh9DbmB7lWhgF9GgGHIDGDbAEyivsuxtSvT7lJdRRaW2GdKuxh2Ondrz2Ip
j0UuDtdtPn1qrhgoPlcFUAusf9UIibOy1RyqXdWBJLzLpa9UogCuLyzDdfMd/fyK
5sUiCBfvw4YW0TjU3xUWCqEQziPIDWkbqrIHh+p/AsQA2ERGdCTELD4bIfVfESIC
czLa81XAz6sjQxt+xJVgKYdswHwwasnTO3iiAtcIzUIQMcg46IHul90tyXa7cMsB
NA2IX6RtkXoIkERAlf5T54zlLlHnNqdgs64KC4V7WQgHuam8fhlSyPCwZLXOSOK0
+x0VZU6OGEych0+O4ZSmI9+/PaKmcBcm4osVZ1vsz4WT7HGwsRBOMqd003RGj7Nm
Uc0xjUdCB3NK2CwT5BcCn1R7qEy/G5L+hVxkS/x5a0VRkoIWT0QDmdJuWJW/Wb04
Gy0UPe1g19EpZG07/KNFE6hH6PqRR4sV614M3dGnIz59sFlUt1mJPF3tQaEEbQO0
8/f5mNQ/gsHfPqT9Ks/ORicz1Uc9RSs0Chxt0EqLnh7CFKXcKJCQH+VtlxvRpLPr
vmvZ7ZOsSh4HQ9LkgARB0oINPvP0bUQS9u3lKcoG7tKdaait9ztNEdZUY5yDCe0G
BAVA4lpDski64W8MAVYjnb0LlUziqeXYK1wd/ggwbivg87VEL20sEPwFz73KwUI0
9y9R1JX8ULYoBZ5C87K0RharRW42tJ9Q7L44f8wSktv7SvkMEum0kcUKD38VI2hd
VexvoatDnaYvRbJCnC7/7Y0JVODSCa2puIl2DF4CvLFRHZIPVfVaqCnqfKWEdxv2
Se41KW8qMRGy06VtvRgZ00efH5I38MMLnDP5p6ab1brB6UqJU0jFV5Sjz6bv7Dts
zpD1zddb4aFTiyYRoawE7yUAtEhjC4gkho0sP6Vmi1b7JXPqvuhq4x1tsiXb20J0
g8siDSm3K9bizusQuXc5bvxZd918r6ne+58QauTh1GvTKKMB+Szh+F5y5emSAnvJ
I8CipS8FE6r2PBoCAfMUfPHu+LEtBnISdu0AcYsRFbSEmfujnkY7a7G1QqLQa07Z
Py6TvbMG8uPbAKe9A3JqktE03RxRGL8+vBDJXJkgucHG4qN+QQNLbqwk7cRw+QrJ
8nIxYfv7r8bZlzX0Co1WcRXo9zeT3VTjaKP5wKp4IRyjtToEp+/FFU7cVBX2uHGf
9W2VMjgyOtgREcoAruxFkmQSogMEO7+sikhjEsJpnjacnAIsFEVFspoh6RZNz87h
0YO3SOhGrnx0mWK5msH1qqne6iezJB/6eu4kpYAxnA8lbDRt/w7ww6EKr+tY+lJf
Z/tLUaVaXfJeIAF6xCtssv/xMV4F9hNGTjgDKq1DuWzVx5iwhCnSd5FeIesLhAqb
e3nyyi9QNp4D9nl4l5yMgGPXVAESokzLNIXyvoW8L5F/2Y+7zfNMdJe/j6Plrvg1
zg0pFRxQhVJnCpHq9Oa5pN53beU+EWFvAdvGI5spLfwavLYXTjGOtN7FfJm+xaJ1
X8ALBLQQSnG9OjUUf/UPNHrVITRiSG6Md47HaPn/8ZSBztODEh/5nMAtexuPJOB5
OOaS90JapQENapFf/6ItmUlCMhvhNKWbewKtVyMdjYRkosr67HTQ4HCx2RRVzAdp
fd7FAsaRckXXZ9vkqRumTxKSYxloGPgEnW4Qp+j+Uo2zNbhP3hX11L/PpdT/++je
mGeCh33ubb7K2T2BiDW3HjYbBiGmG9f8Rm9BmqwgQIgaN2+2hIc5X2qwK5yUqN1l
wguWGdwfkJbZGOmtCjjgc1SdYVO1EEaSN8MnQ32NpjIThfzyYAB5OrhUBlbj/r+d
NV6XVkwMb6LCAkgVJneoBlQJfqKmBM4sQHqhOhd1TZN/SRPKHW9xTPzWo1DoNv6P
B00yOxK4bBYoQ2MpsxRWVYT6oU0XtHNQxc+AtiIthbcZrt20fqvA8dCCCRqBHM36
XgZnCR5OQkR298MTDZYvnpmIaLSe7A2Bq9Zr2PCsVIZWqpPBEVpNmJDnc/vRmuCU
fulJtAIpmaI/e8Oj7Mexxx007F//Kp4Zm4Zj0oTazMODJIq0MA2fHuqNg0uq4Ox9
InuAVVDW6UHH+08JaUddmxT3ZG/upry0RC8H09ZgkRjrJNhEzRxzNT85U1vn0H21
CoSX9bJXpX7370p17BjcA7F1o3VbsuhyYrKGFr+/iwX3AKZa/kp1W/4bAAY7yxVn
hks8x8oT0xfjsJopmrWv0RyyTGbP2Uyn5jCDwJZwGTdW+6VB+WLCZUbtytVGucdv
cRMrJqDKetO2VGMEKrpalY27F2Gpq59GkkRXZvjiNZnmrFgfK723Ge0szZ/7WXZp
axkJrOfczIXC1GUvpmjjBdAuT/dvqVh12pbdEMw5Qp/Qh3zCXnZVJ+eoOC8Oy9tj
DOCbOUCERZUsDJtRPwhhEoh9Oc6pkiMSl5MFvJHd6VgW1CTW5nO8Whdfz1Qk/7Ip
Uag/UNECLQlq2Aq0bT5WRyxI7P5YNA8Q/+tY2DJIDgVzInOlVMVqn+hupXYQnG0v
YXm8BnYyTVqsHnY+ykJRSFjwCH8+ljkN8oHn+ckL9IvMQ6pUg/lK7D1ZdsMAR/62
YTW4+46b3yZvs7Z7nO6NnbOd7epGCFykkU1bvfroTgevSHQ9OwffMg5arB9MgdR+
BFLRhvBn2k2vQpY0amerbBt/bSsSzcqkrbk1V/X8Wv9rSHsC08ENq/HdyHo2kVHD
ibGoNNwhJeXnhX+HuuU4tc8gBIm0VNDKd5cF3dbbIfPVZgECWEhWZZZ8w8a2mVfG
dsfoSCWVCZap3meK3T36lxc6oLlaaDV4SMRueDp4Ox1W/bz2/hn+tFqFMspI6q9m
/ygjLNLVlDU4V4zjuoPgE9wmTQKjHsuD9Y142glL/qiRbPhCRcnb8ifIiGxN14Cy
+IS2UJ1U+/bytis6yG526nC22QG3EpuQjjCPjEJnzM/w7MObAjUnf9zgU10jx8TW
mnP8KF1TXLBFTDin//eD7kny6wdr75HvQRZ8CZBV47OwD6bzKxaMQpFDUyaUbbof
Ec07/SMxaFIQhSZ8ZjufyBu5axdbtxycxLQPCYjRW42E1ZUj87Rpt1uk6tnpdzkA
Pux7Py2cyDCTTjKcZGGQgDwPJFG2FktPPjGPwI2qwEBRcNpeptwpCb5+pdbEfO12
IcZUs6zjs7xXXUuggQdU07rbe66xMf7lr8lS8bumzXx1JKWRlZG0Chq1fBlElsGh
kEOPvzDURcpZ8LR2RipqG+Ipe89GMGd+j8x+RpdXoD7TICpJwWdali+Qua5j4osk
TKB1RAfNDdvv7pH0tXDsBMxDRGkWdy2uOykt/VNrWUExkmg9Iq25UoYa9ax9IETC
vd0Q3LLmH6j4N2zM5mGI6eJPt/neV+uSGZTtT4p4fvgZaRxz7ugbuNsdh7gr3Iv5
HQosElUHuumvve5FjRtL/vvwnDhH6l8AHnhKkTHzvG3L+vgSIaX1xZDXXGdgmI4Y
2y/egbBGTGodkyYrkTSW+A999Ls2VCfyl12CZicSMR2xfWmh7592fpD6wLigvOmS
V7L25JUMSmT3v3lJR/iQQZ1YZUydEUBwmfDzrGNGkFgLq8CygxGvzijAoOBnRp5G
X61GajMQAFXctQ28jBVYRsoYVmvnXJIIf6N7T8Jcc/CvXqxSTI+TONy5jIs/FanL
Y+yzFzno+hEgo/u4WHj25gTJ6Rxg/CPy97t2Krlgy60kbN5mow+kLnzp1+2ahKc2
fkrGMgio2tVKa1xLjEyGO9LZQ03b5JTDhT55nziFu7TjiBl4AwN84JAEEaBs+3/+
Dhsl1vatFWuxAhDpiPL8v4DcakBgNSuXxkHORxYTp27cIoikOlNEusvW3bwDMPR6
8xPd/LKgamaxBdf5I0gL67dg2N2ZbTLsu5juaLbQmCofhG+2U2ElJZyjKQYSBw6Y
cYGm7jbYpMIzeeNasVivbpGfGRcGXhoBStsEbuStDlkk+5+3WtQpbVno97IBc2r0
rc3xZ1BZYsLWtXp2jeWLLTBtYBgJaVaNljVnpC4Bl4N3Ix7TPfoAIFIhM4HnR0XI
DM7reRv+bhtC8wjovLfNLgD7MfLo5MPaW+4P0EqijSSgC6IYmSpLdNWf3/U30NWo
YYZ283gpy4I9vj7yHq+A0NQME4NvGsGCK5O0ZL7gI1KtCBGrMCLlBi4IIeSejNJY
aWyQJNBwIgmBOY/xoz27K6buGLBIblRNU7yZcG2NZlSGHuHlTev/Ak8pyg/P4QCe
NwhDDZZHOztnaIcLOsobMPAKi5lred2oconfOZrYhELTt3R0m1p0fZjLEy17gvBg
U0uEEIdOH1w6g4nw36pGnLgodgs9nPCrdGOQV9qqBHmzR8NAedagIv0uu7zlVqCu
UIQiyPTwCykeCV1o9u/dO7t5CPJIOETX20SpVF/0nhAxp8RGfvPKkCp9vsRroDAy
WQaEPugs1eewNspV6fXqrIea+5VdeIuqporYcETE2toa8vEKwaEZRblfB1WRR5os
YfPkb2GAzrJB09NN7rhELY6WIJuT8DTksdjH0iZ8Dhjx8SaZyZAqU5Qzz7y7m75y
0Pj2tYTHkz4SF/nzbxEmqOAJpXDaBaOlCdzjia8VeSFjoAPtN1d5ZCXaP4kYErkA
j5uqm/IEnThbmHzSrOOYRHsEf9yqCUAq3O+x26Ge4uILGBIxKzKNBVG1psUbfoOC
gz86kY4o+eOtQX6VJ1G6Nr5Zf26Fyf/olWKrWl2twyqn88ElqmZdmDYlvi7CL4+6
e5KwWhEOGgAM4hQ4zViUtHiuY63w6ukuYCApVQMG+tyaDiWWtMmPT8yBUzDWTSpJ
uER6ph6bu/mo0ttbcsGK9fBmgYqQrTN0K/MddOAu4iepso0yy04iWI6RpEk8ILoP
fZz86Pjubeie5tYmjAGV3EJGaslE6jlAtfor+WPSocnNBZX1/hljoEEZAfGxvAyB
FIHFWiHeBwMdVOTSXFuhHwP6Q7kqfQz3D647gPfFqPlBm9iD792yb636tFhsqHmL
qErBzyI1Z3WgHDmeEqJCBBLnDI3tThosKNNssHj4jSY15ErzWOeUOjxi62YKyE8q
p1NdCaoEOjMkD9tTqQj+7MJcT/JkovBpe8JwaIQsLdh7A/0+LrzOuMTelkxK+J9p
3oW4yzL+fGCW3BYl0u8HpsMpgDlPLTUQaQkvjZgAnsNp34sN2RZlCfhvpqOFhvFg
POen1LN4KNtebotu9b60P87ojQ1kGe9eK2cM59wN0ZcstlqlWdqaf3UNme8O5SPa
uQnPM2j83+TyC7tfcD7Nsk00h1dhtGJkzVHwDrO16UoU12nWUoRuiMYLjQ6AslH2
b7/hWU5vYIBuFxpHJsQYUhuJU+hKCUssSR/UO8RjP6m+BwyEjHmzCtkfpVZ8rbjo
wFFH3uMBkPVy0CV1nwQL/uuNMfXz1AV64PAonOIQpQ0AB7Ui0oiSJb4uk/kQApCb
WXyTVOOjVytJWhMGjMSUyRi/9FBJUIAIDGMtcmAVS8Op0ft6Z6a9cjpMJb0GcOt4
yrNNu6xPay1N2JYE7vy1u2h86WIbYFlh3M5tMnIe5OjuPS6nRQEKrAn0dZKNAY0K
j8PZdFM7ufNF4bUOeBcG0H0GH6XpTq82k1YBmuuvngf1J40HDcAN1TGgpDz8hAKs
gubdz+wiD12LcZRwn9PiOmLzL4fXqDsIYE5y47op3lYR3f1w/HZxe7YSLRYG2WKv
5YK1K5KFqHKfTzcCb82GCw+YXjtliDidNDaa2l3kzwyWrvwRkOpdx9uxyB6es9sc
UF1oVMRGlh4+6tMwlYDSYz/SM9GKKaYEWiIHvi6QbPthscP6KTZ85TcA8GyTN6Mb
BwUfeZ9DhkgLb02pM9RgHdhekBaCeQjS3xpsDLpeNbQxfwiMFrAuqV+k6e2XoftP
bwGMP1vrV+ANBYi304m3Dm0ikUuF9zQVOwA4+2y8yB+7LYDRZqT917Ga46BJDglA
H9idAFavavCbEqhrhcBtU4V1laEivCx8673uQ4VLYsPIXRBv8lp2qfFOxHoGrCBB
QHww23MTMYpiRX6UJQfS/aLvc1jeJnkAkRxJANt9hcb50Ru6MCM4X6Ez2gQ24JDH
rmxg25dMAujylwYDHB4+GyXuW9GsUVNp4M1IKG7DjBgAmYhwEk9aslRUnIQji2VB
ZIWsnKpTpIFaIdqgKhd3xO9sEqNNGk9NWJZQZN1kv5s3a72vTQEwwSKXYTmhp9dz
y3sYFaQJUrS3ACdxlT5l700umXvAmje8kyYwKi9w3vNJz/M9Mg73eNbNYv1zoqv6
QhftcWOj+H5gIL71O9k+z/uhlwFk2Q8qcbqn9KU/WlUbvAHCfSD12AIz97snwPBw
UdzZ/VsP1rnBBTcYY1V6B2S0B6B1xY/9nHd6JfoWVOyzo6jD2hQ4d+39Ib+Rju5w
MNYAQJVxNlgo/T12Yu9ipks97U0scp3B+Nzl3NEzlN/JdldLZO12bfoUeucXzHbQ
oB4k94zudP21TwumwSCnwlue+f8DSjYnlk9LYB8RUSHNe8z203jKGdV/bzfo+MPm
R3HofQ5UVpWo7N2LA9w72LMfaF7zC58UdCiRXHfm3wLGyIuM4idqccMGQiQjpt9U
OQF7qixK56c5M1KGQwnqTea47YEoLP9CRF6+wkDsuxFe/uJO+3ul+M/aemQgppU7
F3zbfaM1lQ+lsMSAq10ZgKOfD2CB3m7Iyhyh1dTZAIGdlNBj+mNeHEpMA0EygKH1
wKzf44t2khwKEYFAT1DEmK/3dfUowUNWp2b9hA+9KLwGjcbhaZhbOfuPuMzG5XvL
CiYczaYycwaU4JqMUzHTz6ISKes5xkaxaH+uqPdPvm+lTzbpRPyoBRoVY5MNYr6q
T3jcK5FfdUrGD968mY32FuBudbig66X9ssdgDY9vWl0XfG7ngdhxdQq6c0wom/TL
CVqU1z4UT0OJ9UkAkdz8udhc+jyF+98f4zpJ1EPyFhF5dao4ebxqdgVajc7ReY4P
28mP8mAZ091Dst8EQv4+ZFmGQUsTkYq8SXfrkTj/NOU5waQlWQvZ1aK2lZEZAFRn
MrHwQu0/b41RqI06rIx53yGD3fEJp2Z1ANcxBJlqnRx7v4pcRPn1xnxMIPvFUSxb
GCuZZ3UVXtbY+xzfwhBa849I5mpv51rHt+w+svUGbXCuzhqNZI81TRtgX8n2lmcE
ArK9oBzyitwa6FNLTHYoxWcH03XBVcQlkTXzUzUC8U/PqrC88PB5xC3MRCAWhxI4
c0/o0yurco63KNnmxVv3XuVbaaQuefvHTSRh8Owa83Jayc774wWUTDTNJi1bCIk0
qn4LUc+CXblYZxGXdK/ae+Q7/PuwJG3nq4yeF1zUboSs7QTZiQ+4RovuXtksWa3Z
VhO9Ucy1eY5l6W01JuyHAQ==
`protect end_protected
