-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1oEO9r+as8hk2dM2yrGe2ZsY3v3cBatdrqZ5HqT38ktumn3QFiI2lOLByWzs8xAg
foJV7Sl6Ncojb7AcGYQBJCsd+JmSVrAoiyGeAtbvWcuWRWFFKFLGmMReCkEmkGa+
jzi1yigdk1xXDV0w1b46hiNCm+VMIQcnFGjfV3m42tk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 84752)
`protect data_block
NN8yRUu2wpuJgQf0r2CcspS2N+YQjwbElOt6VgXdIiFGbl/XEQbwzwQdI87CHzhV
NoIYvMNcpAe+L6++1mHK2OXCahYvx5joYQM2IesVPfkCkoyHJzFVUQP2KlmGpzCn
OzJ1BmN7S5t5uOhiqkKVYrS7+XNsv56zRCffVBbsmHZXMynvQd/MrY0FTdF0FfBu
kzUFZhQXOfMpv9vgg9V+QaIHlICL+r9/TkmakJUt1b/i567cmT5sZ4rc6EX73/W2
BMHXJ1sYc8I/5ulvGMXbRZyRhr/OzJDxTWPgHU3HRosMgGnHTHakV3dasOw9Y9fD
euwkPrqN9FScwIIVcAX3kkds4JrGx8rIXEodPFVYrselWGL9u8Huhhz94BPM7is1
zE3VZoFYI4TMCaH/ByxCDsPYGEDPMem3CfNeTw3VAAoSwK3KWPbXak7pxWUagPfq
Sf1+TDhOg3ROwSC7W4+/Llm0guyq4zhpWlT4EEaIlrD5ZbpXddWet0Ii/g+sBA/d
1Bd7WinxdMCBhIb2w0iasQWi/O421t7ENWtj1JQqt544n6Qe7SYOrbgj2EVL0G15
9r8nuBdq80qhyK1/H4o5m0koxEpO+5e+C0cAgIfakH5rOyO/AYcHdgn+hJ8xY9Ah
2EXA19JVeXDq2kV3dsSvp7sAdz6yxyAlXfyXcfbP7lfcydsUuDPCvxt8uk0OiiU3
lrpiqitkWHB4mpk0ejFWlkG0o9QGJN+rtitVJlLnAvmKNA5DQW1GAZU4gXs1bZgL
cLryydGzEdKRLG7Du5fzH9NXwztJ9ud7dKZDOBPAthScxRhkoKenNJjnDj2wdXE7
GyeXzPJbs2Odx8EDmyAjgDijbfTuTIw7D54MpXjtSlx4r+Uy9xA6Oas1LLOxwWQB
Xe87JduOyNHqtKLXKDtEaHdHSGFdNsfslD26fSodOn0StgzBEdrPfhMOn2bJUmqe
zRvwu++dWjHGGY81/PW1m0q+qZLMDoZIr5lcDwNwld1IsoBDJ42q1iAxl62TWhXk
02ElOJspryXvAwyazKzThtrcqqjngpoKAi6SLqGZutqANL2DXWr6j+f6m4rLuESL
Em4lSEbto6NuvJxsCZd0oLj5adzL3vJE2bR7NzLSYB3Ar+hwxwNt1D8YvoadJiHE
6wfoCRlabQRwJzBICT2Jp0iYNq1P8mVQTeoP1EFXtqzJj9uCyC+UbD1ZVyBi5C2Z
6Me29zWhoKsr+cPpQCJt3nC67DqVPx2JTwoDVeWz9X4igmxv9kPpRbpWNpc98wW+
2mw5YcO0Ej0c1YjtSTAdJ50eXeIy9rKn6wyppQbRxWVq5sW8VEwLISXmeBzqzCzy
zO/ne5ntkkIT57df7I8vRodr7oB5ty9ypNC8n3GN+5GuPRIkWIKVT5BlRqbYO4W6
Bhtxs534Aqxnm99dS6+UFGyPsUkvcH8pu/nSjiY7uEuCN0ybWYLu1KC6HQ6zpXpr
h7SE4ubX7rGrBfBvK5pEnlR9naSX/HeqMD1BrWx3MG0G0rtHy+a1sENLA37BI5ri
9KbB/q4mQqXSaEns/zMKNRFInXLQIakijLmfKLYQL3nVPybIfIRhB/EsuwZ3Zp1r
jBrpTD3qTi4+aSGfhjUmm9ld+nfVAQq6tJ5LQEbrJx8RDd8mo4g+DbUvrvkmHe1u
W9PUJKEp6GYXYTBSBnSyBJa5KgJ0aFIErHNlyLBodkH/N02T3N3cnmv9OfFHJGLH
7PLPWv/4Lxpaoehcq7ZbbTVJB08IRpWe6Y5K4wj2Yyo2vF21YPbm93H67niSe4NH
1fWoqX1PjMKPbg1ynLz2PXkAUR/z0PAArRwHlvovwFfs1EGh8ATRu0Awz5/bvjtA
C+UD7F12P69fiyoi0RDKzcEk/XyzL68ZDi/ndbM3m2/ZZ2JOGtqJBd3vTbjFcc8o
hozhNzSWqaqRcXwiRFl+o7kSK6ZJVXzfBZX3D30mQrpZsbrUX+wvRbNmyZyR5lPM
CmEzHAbDZC4C/4zNdCGoAlOrmJU6jVqbhG7eVv2wPbD8meiK3UyzA0otIR9dDlkS
Z/TzNRdNn2kzHP+aDqwQ1OiUtJR0pN2Hs4qXVq9K5PsZQ/S+97mYguqrWChBOpaD
UbGQzBK8M6+tEGfr8ZsQOg+UcG7CPbzvVSkw6VtZgWfM/gVP/daFa0l6nM5xs0ev
BlN+q5TaFzbXOIWolqIgkV+drwC9R8J3hDCG+6yvQToGgi4qyZqXqkHNh6R+wiRx
4VsotKYOeZQc9HEYHCYuX360MkQAAY/NueeFxR1dTgqoyTDxbO/fvj/z3xxzgr+8
NQqchviIBFLHkfwCexrEAM4TnxRhRzbqe8PhaXwCi+mNK8K0Jsa8tnMVAwoEeat3
YKQvwFopR+yFXcW9qB1weW3kzsmgj8qRJH/snhfMYvUoIm9/avfYfY6n6f3hrPKn
mLrw3iSpFHz7giA2sMSjLKwWNstnSvJaxuBwswhxegf50JfC3xTeH2abHQ/5GF7/
zAM3aG4I0Q0LMF3d2K8as9LK+v3UvqtDVcFvy98bWz4gHexqI0XLzK2awfu29cEQ
MKCdZEz/RlsXmqQmPwrPR7N/4YmrOcqsJxQr8YoyRlxyCTSbBddyI5bF5Dn/KP31
dX+eRz1MNEIi4GMrQ+Xkd90kQIG0YwlfXvJkzjHOP0mB6FNX+Ko9hitXxFGMQ+hE
7iEVMFm4qaSb/EoImxiKqpn8xVgXIjapu2igCUl8ndOzrBKv4N8tJBCTV88uUHoQ
m/aRnrDddwnKZcnopNuMHUaMYJjTAMiApYtIYU3/pVloQMBUmOX5POGCYFP8NI7o
NPRjFZQ+qXmCfurrtA4AJZ+zCZGpM1+z5IAVKB4Mueh5kSCKCGO8KUPzO2KZr6Bf
sGFH2P71LcmsY37OGndAxdNldpIb/lV8JhiVojbDPdrbbDzrIli0TC0yc0AeSioG
vyGX8P1PVaJFtsMgk7f9RMOPmrzIk+j/NQfIz8OGtuYA2HyDDLoRBRxJmjEuCns0
hoN/ryJMrQVze+EuNLhp5F2/pzs0BPPIGiXDVLzw4XnOfVMA9K1Q0G4lcl/w4cZ2
hoc4szDxaFRSuTj3iiTk7wA8WVMymEmcClV9Z9I+Fa3CqZP1Cv7Ms/7fyO3s4+wX
AWaGqlfyNve4J7alKRiQfhUrpGHJa1mlGSqjKgyWON+xE2F229pcj0RDmxAd62Eu
y/sEauYM+EU9ZhDjek4RzqZfqQANYzok+ITFQyv2k0ltn4ydZ4xTnsATcX6BgIww
DA93nW6Nm31YVGaQLlmz6NR8vfWWCwKg12/ktKacMP+4SWzusQ7q3v9OXT0RedBm
iGCOiEytFwrTpb3IECuu2esG0akbPTtw/eqbUEonjpxmY4/lAvwUS7eK3IlEntjj
mN6+I28MlWBs3WQ6q99VYGEpQ5bi9wEH9hiUWYfeu5WD38Vi55bDKlbSXAQasr62
Tos/PO7YtAPrzR0EWGwLjGLV7T507c4qzsTvRhFKG5Ar2BlLOOBRbaVxHjcTp7bg
0/KZ5lMAcJZr37XrnVK7oDwWJLyRDqFQl18FYD4iT7EbL/N9a12/zLaJDUFfkeEz
dG7ME9v2/JZv8sRM4qzQWVSfHMTE0FKobCJr20K76NWjEP37RGa/pT+9lhmpU/WQ
Bll5Yy2y6DQ90n3+UdMD7OZbgsmlh90+lE81Ng1k/qZf5p6uiYzGFzbGbQT3WCpX
BhilP5GS3rccowWBguESAW2sU2cD4PaV/fFcVpznGUo2rnxhb21La4lhTD0pUfSJ
GCwgO8+WvsI8Jswkk0Re6LApx1JcT04mRYHuSXLSQ2hyjGRz5JO06gjjm7R0J7oF
5ByK55ZWkEE1w04PFjCJj1XrNsXIhItwW2E3VoPp7nnG768fBYFMSz81phWKXLXo
QdJRCggrHNaNgHQrWcL2ZSSJ8PAvmCcQvLiTr6o1FKgVlZ5/WawPS+7jUJZ+ZYBs
xce1Tvh5rDUr6fKNQvbwx2Fn97M3InMU7HGAxv13jrgzil3LCWei+m39MaoIg7lj
bStdD+Jy57erpT+8QZU1WKhWG3jJF1RwOl3XzD91+5Hipc4UBvFAWUr7eZ62lH0D
zuAujKzwzGnz0EIJp391derEAsoZhGaAUn2+Fx4X6Jo7wgSlmfIRBLar4ObmTV/l
3kWg5Qpau1TPywDWHQwAtMzGwwbkCelsvOHAJIn4u/kgh+R0T7Hk6IkXztygmKZ3
kPldiXojTkWyeG7Ex3BMYu/+5lmxTimuupXnd7bIp99v9mmUenTtMkiCwFYGA6/y
Vx0Eh3Mx5euh3fKDkqcgrd73sO9nZjcSTrFy5B6FE+HPZPlrGS2zfZMIz+r3/CYJ
hCJL1D5P4r1Grxas8CkQ4t4iy3UAI7GRtX5BfynpFgWDJquhjxNBIQmorB+0CasM
6SqPJoEWO8nQn4/+NnuzSdqfd3iizH6nUa36H0lDKY9MMp5CeC3J74wjWs+78xkY
me1UmM6vQSiqpBWz2Ut9VaF1rwEgMgAxzB3ihOh9Wh2WTFJwh51OqrikGWFkP+UV
vABC83N0OKOPDq6perPgoXQDFdEO5j+UHkLLCUQTOxncgu67oslq+IuUJ43OHYC2
TQs7HiWNUh5fmknV7ZNq0HTP4cpzNQRLksxWc9992aR5gWVFuxloW4lfHjftENRR
M84kw0YTP6j1b+XubZws7QMeb+/jip1x73GuSs0ulOLRyDMksutnDSQhWLPeioo/
ztJmhzOrR6yPc0APTr/YyjocNbtmUzurW+3fVnG7dU5A3OhWtuo48IL33fED9Bf9
ch86EQJE1XObFI8Np8OrkAkuX+u0mo6Yg6Xoric1sAdxnNEEYsbezGPaS64SchQC
0lYblDcVMoNo3GVIe1qg0U+l0lqriQ7lIOzNOve2USjVlhyTGUZ+PKgLhfDCsF35
xXXOydI6BTH/7tFip3U2/LFfITnTRuh18ZCjpeiY0tYp9ySCksEN1n/0UUn4I/aI
U902Da+tiBwsi6ADA9GizOvkpwxIdLpwb3UxE+CJY1e22BcrbhRPg1g1opoGpJjn
cBHLHIl6cPw6pdj5sTLlCeCGNxfkGflVfQcpo8eXZCAwx5np/E7Vx3qebt6/PIbR
0uBXSO5NRTEKSsS5UZp6YGOaZZ99wx0b95YyjkOhn+QTZRMFQHYSGVZgWngDniLe
46cbvPIgeKlRnO3G7f7ov0VXjTjvhevYDK+WzbZBwwXTL0rOs47qNN3BPbAd9MyB
UmCtpO79TGRt0tYcWN3Ai0E7ozfY5El9VeFlkaCQ/n5VpcOglEsO1kz3wzXd6MP+
Vy/FTesMotfUVBtaQC3Wm6w9qXwxIgPjqaQCI65nPI4SMzOpDUtgSgygngQyjc0c
g7WxRmwC8u1iIHZj7OL/BLCdjmKcqLT1rR20j6t4OpaosRwCdicqDtOFU5meQ00u
p/HrPiZ9WIZUf9bm5NRL3LNAs8WkgULYAHp6Ggmh2h1yZ9yWq4xAeBOZySnj7ti+
2+LTT3V+kJslrTc0IvzaAjjuxRhY5KfuOUXoMyJJzEc9L9M+HXJceJkChN6MwSKI
xR5HyjhYkmUWxguDYKQD3PeodrpJuHgBCSjd3NP+Ln+K6R/HKqk0aeCRy2/ub7L7
sFf5/A3nkyk6VgqLlKMRkBItL/NQzfNJey0kWay/IB/MU2a+0V4md2SEQwxxA1lS
pQlcYgssGtzxpJDjgKsA8O/hTqGj7zEO0uNYbSnTA7+HsMotKfKHYHuB9yhRplhg
2S5OpIrsWaABXGHjORNzzl3BjX1Hd6WzV0LT6hjipcA985zXfdYr8BmDIN7+usl6
4/Y59bWH879fbxHCZAxYSCVBPKKWNPZhhU6YWG6UUKkVGXDvZ5/NYihLaA0cW3Bz
CRtkHrjNe5ID3Sm95vRLGJH7MXOGGFZi45+2N97mHGa1GfGMMMUCHfqBOk9AOkWx
2YlofDj1BnspRVQSm68QgnfMYOSB2HZHTvWQ7HQka1BclRdVcEzUvRPVvB1eid0A
RVzIPWihRcQUoxtkCXGbZ4THf9PRmprgw51i5sk6wdWVgq8u9DAX9BxEdSo1/sLY
ThVyuuTuXS72B9sFWhzLuFwlC7RP4djdBtPnrkmPGdtxLSr44Biol4H76Rkl4rl1
77a6AJyP+4aE6MDZlXefBK83LzHCMbP5b4J5H6aKvtCMICuz+MBnw5ajBAhqHdw0
JAwvyof++C8cm6AO2k+sD8n3OzvualWYbW987pqJlvMOtpDLoVG3XgSfQp3cDO37
5Bw8a4o5RCtM4DvzkXnDIk4f1N1i4lFZtdvrd3e9+D2NCwwiVcDA5eFSyv6I88BM
ty/Dq/CoC1Nz73c5xp9Lkj470ZUq9gYmxL8m3yP2nqIs3WO6d7GDPkTUwthvRT4O
k3iFHqOIgpeze60zkEdu1HQ5vOX8ANanU8QyKjnjbjq2QgHFwifdU7+C996OUKDu
JGu4P5Cr3166mS5QqS7hID9krTNz+62Su+x3JW0+RqA06MJZOonEWJxC5rHgHpJV
0aNHoOpMv0HsQ0n3TbvENJOCx65dZFO4N9hTyDX2E8FlMT9v+9CUiv9vzdiuRkPL
SI4B4RcUxg0obG3/RbcqWPsWW0kWc44mPxAi+6Rd6ZIGNuIsvIqi19SwWRvNRJuo
AEGxPqkIwjKQ1OB9wpdGWlHunHJ69LWfe9Hbyk6Vs/rszHu6xXRnxy43RJ1IlL8w
6m83xTAognFIX0ZVjoERsQCa4Mx4gehzVwjkDqLmYvBbdLmf5+WSuXRA4r7RZ6Bw
bcimsvxWj8cHQXD5n5cUjvsBmA+X6EYutYO9OAy582k5FIcN3mNMw0wCW/uWXzR2
idcilJkckEdcrynPi/+Ddx0FYeMkPEvqBajARobjf1OFeT8qhn/c+HWm5E6z8INN
7naFV8nJb31QP7pY1C4b6YglPLCZBJJgNrhibm9eL7LVjctqmvw450xwcJV9J+5N
xQLx7FfHNG5BQcSjU2XpY8L5TJdIvyBGMR2WK48vuwe3+Y1sfoKBWYk6cr2XQspw
EIr8wuONPMQt5n7OSwrP/pXV+9k8pvsu20CYB9W2kBMb5ZEmU/tCj2UIWWpTnrq8
oemAjYNsGPodUFMM71oQYJMaki+PgmcF1FxUunJCNrVCgOlFkKYxcRPr/9hKgGU+
iZ0Cgjqty+9XuB0+gBiVFEMHVjlPafJW9wkrHfV8wc81qhgMsf9C+gX8HL4TZogr
UFIanJqONqteyM9/ljMwgzRzzyP6TBM7752AFSSYlTd5P60TsfdMb7xhkTKMeu0I
MqBIZOKYm1Ih9/2T5ZC3MkAXP7HVp54yPcT5JX1hjpo1piNJKKiJRlbLoOCGHHGt
cxzGR3hrR7PkEg+X4yj+i2KleFPK1/YIvm4CIQKRC/ihi9KQtzrgZIHG27E2YB3w
G+Ex95lMZHGee8eo4GuosAhq3cE8wqr28cLlhDWqhJ13EZ5M6tzNcwx1ZvDSXddl
Yi5IHw1V/J1R2JHQfXaheprmwwwKHXU5GXRoBtEYWKeXKp32F6bmf+2G09Xnfz+4
GjmYESDoYgj14PUay2M9MHw9QvcQz5hhG5j/7xnoSs8y3/21mZE5ydc7z8v9qc9u
XDtSNGFfMTaLwENPAg+DBTcR6cfLfKB6rzoU1esAdn+PzChsW0D/Bx5WlfUar1DD
gjMvko0NJcDcr0DKjLK5qOaowixCqX+jBmo+zWs9H4OrKPxvC1FE5gl700xllrRq
4Q6BsmC0R6qE+dwqNLuke9E0iwp2M/rXrEByFyStXc4iEg//BCWP+z9Uw9CeGE/B
91JDBQgltIyIPyeI+z+nCm4BARqxNMi5eru9sA0oQtPg5MIWadMun79huG3i5NhJ
QN5ySuZBB9b4YjR9cr0riM1hpVhC4XyBAzm92KQL4n7k2/0vC7QpS+YCXl9NDfMh
QsVSi/QKKzLRophaAjUYxeHpZTmbL1vNfKvtk4LCx5nfhcEEpXIksXspyt/04lM2
2V5zxymMKvylFddtXIeLDGGkEAtsccAsPOEFhOVWK7n947SPCeXCUvAE1YztOtMK
jCYiDq9wt2XlQiqDqWtS1u2kpZOSTrMnv9Zau7qQOfkipYcEZFPjAkaLebclRU2d
0tGu5I3hJWVzKVUSZOF+kvPWRQO7yAMbhBt6Kvan3fxJLJcEJ6CoW9Jm5JxU8hnr
F5XJkDcLm8mYXnSSY1nA7EuIw9JK8JvAf8WUpUFR6DE66PJqftEteiOhZrmDIZta
/L9xjncy9SlkWvPHW2UGJ2DLBU2XpQPPj4whW83qqgtTcvKAemZLpxlWMOEg61GV
5wjr9BD2JJMgYrozd5qLyYP00NfOrZbcuprBImOBJj3Hpr/TgS/Jgsj1ShpoxMXN
vvZDAVBvYejzP66SkygyXhLI3L9XJws1SjR7vHbCDkym65mIWH3FSwkaPtoEWOFP
x7x+nVpRu6Rjdk+pmLc49IMMaALGvVeyXLCDSOPA2DDx5uDYSN3o262VqPfxCJxV
yXmx6niO0BqaBPwIlriCpT1jtoWH6G20GSedKU/v7QDZmCrwCOYskem+eU1y3/lR
33rN1HdvICMrj+nrmty076I6/eMnPdY33mr8+t+h870NNXMghKm5KLRXbenbkKcC
cBKxX/RooK68F4yZRwK7EZynZtdFzzVOKWOuvVq/tjYkRm8NUB6wlveQTSlGNyuR
jUrjR/Wgm5MQesUdFcFM9iFr2EdS+C6TNfTqv0bDomUqPMZHdoA/D9j/CdvW04Zd
beERZzcyazpuxhoL5D5/+3dAXztZALrZ8Y8zxphLCUk8WRoMGYXgwCx5swbErD9J
JaKZY+gAL+BpQ5AuB822RG+WAv4c0RlP76UnnCK6KeR+ss93KxSY7mUjOy47k+i6
UkMH6Yqeilxtdj3l+nkxGf3iLLwI/FnfciFq2Epm0/KnHj36PW5e0AyhB7Z6pEHX
9oY0x2PH+YA/BdLzzn1oZBu1/Q7Z3q9W6lGaiKII7f1JeiGMfLDLjdgFb/Jg+Ccy
VTgy7JRd6e7R+laq8wjXqmL1yvthESRf4c+CjRC1N37CEiDneso4mYolk41chmap
NqpfJBkn3qAreiEMpNAOEQ/pNFECHBK0zLtoqQTxkDqtuS+RN2f587PFOFOh6fLS
GTbzR0SwN+xjBjVBRfusOF1Rt10BCR7i4Bsv6QjOtd0/Lu4rAwV+9Dkk0FQVN1DM
30jeTpcP4+ao/mBpod2YBqfYEuT29FZbcoUp/L4bd+QyK5g5FBWV2QO/pTz74t2g
Qec2rH69bANIV+Bo09Vf4XLDA3M6Q2k0DHcMYvsTRcP+PjkoSx8S1N5WBNV4bOwt
OZYJvCfaCGAzksk1ggenL0pBouHqzyq/X3ODQtOBr6Jv2vyfEeZe8L2bn2BsjuIv
W+UbLSKmj4aBZlU6ofvsNhCG+4BcVHhWBTtP3O5uSVpImmzOB/7iGAFQh/ngvMG/
ai8gdEBZoKDXuRJXQRstrolaxuF0Hy+r3K+yGebvSlYeQZCmIo0ZZhb1bOjeId/J
PI77cELbirH6rD5soDrgXIjctwetFhy77HyqOgGEMqJN2MW9TFAqaOLv5p44nvns
m9ubUfqbphbpuv7ndo1IEe73shRMe4GODLPEgKgkKpNo6Zav1N4r1z/NaU/t6NZS
EqLGWO5HEBMcclnioPAfI6miBJf2rGh0M1D0kCxbTC90TA7G6lhE2sQ612cSsoWb
RW/XTaGehMSnDxHuSBWU388ZyFigsF0AB0b6b+HY+EI6uZf11TGDq8AP5tG0lW5c
GgFa2bz6KsnAViuvFIS8EtesScesIaArHpYTpJatjMq71N7+wU7CPJmNOscCUmxP
Z+pu1RXUVELDPRwi50BJH7ck425aVGvMy4L/4zomPtHxXL89h7YToAwczb21CI+1
HFERvFKdTmqlCYmpdEvZVupyU/WYLyMEoIk/Msgn43FnqEtcUggA+jcmcnyBQ8Cj
Dlah7sojQNWkK0SSrRD6vUqYMBVexS5Z1Xzr2mZ9mwau0wp7QWzo1zxED/Vem04i
0Zlk1wcZAe7Zkjm72fQ1OHc1uGAr9g7WO5zMVTq4uraVpZfV9f1vowyFIzQL90Lq
NdnbidHfsMVQNlsGnJTIBMg8u4dbz9wkDYXMbrQtz673/QY09t6b+59iAFR6JoWf
Yi3AdOmYX0IfAZqwKW6ROufz1qVe1OXquTLQjFg8+V5M3bP25b9pG4MD0Dlrmxnj
kwJiRBBvoPhJsS818rdLYKuCbfNYBEYDsRDQEjw2saa4qMjTK4ia4BIOiRVzm3zS
X8aqOpuxGbDx0WOBOVLJtc9l4JJ00nEfVcMaj5y1VVchy+AVVgb6hgALE7wBcZ1I
AwE8Z6WCaq04sYolm5XSyO5Y8Px3erPtTcCJv7wAjQAj2MSpEZZPepNR44f+6Jgc
2rzIcYYj15SbLSsyImPmK9BpMi40P2e3EXFkxw79L2O80vGPZamCTvnkZ4TlusD7
LMTs5nMWxrKz3qY4dXNi6HIIItrpKk76Gd3xRc1K2CL8jrD7pJFQSzZv+X2y8c31
H5G8S9uyz1JL0BPytvAg6hWdjj98R3EhX5qQJkzfDk8XMqUBsmIvmjmib+IVFcsQ
LS8BqTToSZMXN91/NAf/XhudUNntMv887BR844FWbe2wQzqZZ9Y/w/5GBXJIm+kX
Ohp8FHaZfeu0/M+9EvByoO75JVF6sc6ygIUlb+nZUhWxd2oMvCSbi7pp0/Ru/4cg
wep36FVzgsXlLNO1MD8BoBFHaJVNiMOKLKRdr9joO+X+JmuljJRFxN1UhxukCf8g
Hi1F7HcAAWxcOLwoEAQAKmg68lhSYCgfD/M1fKcDb7rZ9lznIZIn0g5jUvx2r9U4
d4x5wlOGRXMwCbIWmyASXh3j0VJbvOohWpLyZfFi4Wohz8rN7CkdRvT1FiCoRzyV
In+01Udl8NobGfBD1n+Acc2OKEt4dZadKtlRufoC8zD6c6SvNq4oZBkwXSZ6TLbc
BcuDP39ADfiGyqSqMlGbiAMBhJGnPQgN+r/NlsnNy8D9hrtYx8rp++7DBetPnz+A
7TKRW5dyGPHpW8Fyno1lUsNr5At4JsM77clqPFSMw0bewr8M45gKjz+4bzeSjUr7
6pIBKvSTUt4fvNKWd7OYm3uzT4f1YBL+s5T8eqTitaUxLx9TeWBqvhOA0Al5aURo
Ii9n6Xaj/TcqOf+LoT7CSVt6ghu/JUwr1nfI3zsUWDH1DSf8aSMaibo1Dsezj6EK
ujnzVsYi46DQLH+i8iCF14Wm85ekMa8CueDK55OEyvcboRTJ8hcbIeQMwUjxf2DE
ay7O//ArKZt8KUcrnHUrsB09oItDj4wImb7zzqo7XNvX0SR8mcOLGcUi4FAOygVZ
9+l3n7E5CjVFgX9EdH8tHuVTsPOJ0m4w4pXIL4XSBJApechB/tl0WplQ3toEZCQ/
xZDny/QUB7kQ+S41W/69Rc5zpAscNkL+Nqzc+EYUVmbrq1XEX5cWJkGzLDPlS0aQ
pm+ZeBtwW4bo77/5gd1AUnCl6fydK4SQZAqu34KvitAMiBJFoLViwDyKrf0TMXOX
Ful4T598tVwO1agk6nFY5qPh9wlNF+v8dXFjf8BmuGuII/oEyzClXRE6Xd4IfQXL
rERIkC15LzOFil/MEPGffmG84m6Eox2vXbQPY6JTKjGO4ssWhgyZbiujKJLqRjdR
mVwOqaQXPoROqggKI3zhLJJRP9FRH6FDeR8dIgXvcD6GprIrY8kFxR3NRZ075Ef+
gQUPx9kcFhlXOkDvRXhzEMqsRAQ8/mf8iZRP9YwMBVUmgPO3t1AUkIac6VoZXwEt
sb0BtlHEI02kjuXk/ADMjES4wXaND2owszS9b/KMQMw1VCuGd+6O/2mIlk4Fr/qs
8IZpAv3w/xP8IVuhQsXWdo7YgFfkiRvucmZZtpcdnpEUGU0tS+3I2DORaypGs/Mu
oFZfrJL8kuMG4y+BLfb3elDNJBxfng/LX2S0+Ud4L9HW5GuOyNRTBYulubUxxziD
2sH2Qt7HrKH4ea13ew2sPIlIU5TiU7oVFJZt0yi4jKq/65zkgYysX++5PsjbNdXf
Nr07yf4hy0yCUhWUuOnkD0HT8i3QLH2CAHZw+snVj0LqptAsexCAGbVpGIcRzGAF
bKIbc3+qtm2JLEm/hwSHG5LK79Z6O/MiKpbelpBtjsAem3PSrBkLjEYj51HOgJkV
56In88LQo301m1sRj6YVITT/jh0AXXKRl6Qa5sIdQnUsNffX0x9VlWiSTW7OG/Qc
8Y+gER1O73beTzdLhVJaO0knx2a8SNwwal69CNaQNo09sN3p/GZsFu+Z5jUfYMyO
OwaTpUybwI6VUJ7T5u/zb8y+hiIckGwUulIodv8jRIpcNDw4ArhH3S09n8KVrjLG
YeJEMO+jVOhPOveItYl6lCoUCT4+fbBzBk4ZeC6qBo7bFEW7iYvmMrVwh9MlLkDM
yXSL40Kuoa2LK34T8kD2INz1MTBsKdvtenKDeCxBbXjrc066HFd+8F76fARPhjbf
8W8Y28eBL5ywNKqK+lW9FiQfsEuI7LJAFhegvLc5gYh+bljxnwoz8GIwagXVXiVn
KjjkWxsMIBykNZDzF67m5h9gstPNGadA2+nAnAOvE/CxEOAx5N0b/I20h7dwtPwv
LQniDtwBCBX8m4ZwcWtjWooC8Bf3kFQGjD9eCgrKMbPyYWHLsHcdVwQjwG/ClNXI
IDlppWTtna2WNe1HsD/k7RZOhnfYCt0SVxzZfk6EKjnqjyuavy5XY6IN/je7VApU
UY4anW2sBUXqblxmqAmE4YaW43ZVyg+1Va3xAkZ2hmUz7Gwd2xl1YLeDngoCtuYl
C3DTwjs6yDn3I1d/hkMKLlGke0kMhXkAYvaZuQ0Ihuccxry8j5m2p3Xgupoh5Gr7
MgKonT2xlsQCNDbYfd7cTziGB7j6iMJTECsyFdH7lelE5bIEJp0CIeZ7vIxgW4bn
R4PmovhKvZUHhmA0wPj5TaBco4UlraWyXLyGXwQqUt1d00gSNCxXmqcMw/osMwqn
zP31i0Q3luTyZJdTkmS6GyemSaJHDUabSXQM+3MbRdvBpu9fzKfwfylOFNjwKAMQ
PkNEvEdMeIQb5Lsr2JfnV9Jm5Ng51hyIKPb2Tizn1gT2DieqyqLdF/Hk5jToGNjN
F+AnhE2dU7uruhn8QWbP9RhCoufegtYX0C7+W+qXmAMomTs3nWeqw9w3pUzgSbVZ
KjqU5S3t081LPOvRsrvRP/k05fAwb5DHpspGVmlDr6hE8cTMiYQebeF8okm12ad6
KWcg5QUYBo1UiqRXJnO8DkrJ/E1cnqHsVAwgG9N3o/nuNiFkWHwjS0+8DUPtQiQ2
3Vj9yGzU12T5yCn2x8YnZKvvquo7eZ0+Otpjgh/0AzsL8rPPuPEX+W1kEI7fZnYf
0JxlYZL/62VcMFPWRhQlmJM4HjK7zQLT/LZsMMSvMVO0C/X2EctCd/4lkQmTLwRC
GK21LcqSTyul1B/o7zNdIqiUtQMFg3fLvoX+Xi8XjfxzbSnxW+oFn8zGxk7lryW3
r6EdCslVxEBln6454joU5Y1a2w4JoYThAHzD3E9lY3Y37rRVWqr1GQ9f3zkYdDZ2
uQX+aEW0czo3+9jVf3fblbGntx4lkMEm5Dw5o8CyArA6V7TThNC3pFU2MXgkqlHf
MWkyVbO1GKSJL8dBpNPfPMeSZ7f7/b5icPZ9I2Bb7wqrgPvDHC+XYn3SLDpybc0s
POy9m1RAfKsuGIeLR+kCtiafE/eJRv+ptrV7BDaUIj6fMDKT0FZDKnoqvlpnKT2W
Kz3FqxdxrUuiVqevm6otEfkGjpPOwkc1gIouleNbBVmjL5s6yT35z1SHj8+gohLI
ViNCq36Ar94sldtFlPR/WiODCdzlALO6u0IWSu73NJ+V9VhADvP/CplRG6E//wAK
fQf6p4ok88qcnFHlQgg4YumSXHTgZShFBtJ2MeKIKwa5hfxfAyrMo6EMvw/ptX+y
ekTJdlAEHKPfaMx/X9Yzdjo59hfEh046PGMgpRmMKwV9ip5Ho4F58xvXb3ShmWiF
4RJlMLj9igyizgmFwi9GGb/XA/x21IueYpdkoCCopawsauCtKejhE3YZwvDWK3Gw
xKT46kD+zEKdbXgliCPQzuRaIUfvBgoihGURz5kO4Apm/uH7kH7Fcw+ONUV2xES6
GfPTHpJUYKiaMGX++UAEAbHnD9DUAeRf1xwATDLEQk2KzDOYR8HZz2I5b8YYq4lI
4PfCh9nRgauxDI5odxPthtw3Qkrrs3ScXaDSCflJv+9zTaN3sIlcmGE7d0l9fNDe
n7eVvbv7IJTG/FFa/yUWORDfQd7q0NhmzTj9eQphjml2nEvm2E+bTqzVcUFkFtkh
ubPvSbwTAP1/xEgt5s1bgJ30f3E4fstv0VxDdXpyLOCkiNIcEeS005UvmG40Zapq
+r1i6OfHKPdjkQTAHVfSvM2/o9z5zvDktkllNCHy38IRG8dAmbYIY/EIYgMERBXA
Elb9hhhohoNuzIrPmAJhSdf/9XntACKO6CkLnEIlWuqxJIj/4SP2OrPxYfEbAlhw
6G+OboM0++C1PJgt7a9QhSRz586SmWRyrpzke/f36APjK2/3v+Q9xiAqZDy4M9Ll
n7NFWoK74cTUf4GaHgK6R9aCOYiOXdLxKD50hmf5dc+ZD/jL7VMq7kVaKgeKBdp7
pE2KsLhACrlhZDBkimgwMILR9PreVn7dWfzFOLSkGBkfm7riks3Nj4loiwC48ETt
xyxGd1P90RxKNrs/LdmpM/GxXUU4WUwqVcTnrDX7LdIyVGbQrolgoAvITsvs18mB
PGhDKBQqw1sp9YUx1ajKW3cIRuYWNT4/JgvdwyycKIvYINZL+7ZCF6ZuWmcjQraJ
GTrgWuhAVKOx85dVVmfsHFQ4LSf8JvpUIcTfYH2kToWBpYab1PFC6Ylsw/8MrXTs
S6Rv+qjwL8uh6JV2YjBmjYBpKCxc5G8zOlGWj6fZroO+eGqhmFSdguPfpegxeCdR
jTA3XghOhNCLowMRcZlpNlimx/0yxNLIGgVh6S3rROa0RYfb9Qm8EKdb7uZNK9c6
dN9PMNO2djyK/3sBpBHbp0obr+1K4rWffuu/ok4pqu68op/TOJ0g46m8T0QwFKPu
ClHvO2JHllpnhMwSi80xsvy0M93JFg3l526j6Zdu7k1djfcPCQH6BilHt6fZFSqA
q9QBAWsHBS2z5BBQULuuo2+1PHGslRr2TjGu6NaE4kyH13MRH7IwPYrOkLoeeVO8
sWTVw8CO3UFDOdS4QuQVh/emhKvQVI3L19CMRQHecMaLTOgJMGdeXxmnS2SHVZt0
+IkkZdi+A0KTFogAUNeW7mIKegPJEVzcb1yvLnzpLqZ4gw51+oZI+vIyKaK11Xk8
LMC/xNNJW0k0XbiJNWZK1oMnbbxLf2ImNO69xME14JtL1n+0ZL7IaNUCFamLylOF
3j5GsHEy/lXAlGOo+07HUv99KmPoVLO8NOCDJk4UfmyR1VAt62LQMB6tcUwexPkQ
4U3flj227neQp6Cu1uabs9HPB5BeRAFLyyrKV84ZEPwRz0PWpx5+FSKnrYq/Gm6K
CdXLaM4heHam8RBhqbQdcYF9SDs++AT+7PaI9jflLUqiy6EEIsdLCyfOp4KD1LXc
wQzAfvnS5aPA24/QN3yxDzKPDnEmrMgjtHO0lw9vf4O7Mc8/PPa6xORVhZRATDei
O9qOv2NrY251mljsJfW90/3yo924TSIrIPsYH5fj8zfYPKq3C0XnC44XfezO/A//
sRcz/wkhLQRE7T5xHXccRZTCd1yFMJMSM1P+FP9LsUyZzNGTVMUVJ/wcSMwrpf9r
7iKPglaCkuod3K9JGBbbSeAQEFn+kX89ecm54HsKHK6ffMwJ42+bBT6feEeFj6Rb
iLZRGKgy9zM3NbLVWSMqw4NqRXpZ8b8xfYtziDgaFVU/ab6i7AbgxSsW8e4tMjXR
qfKBqHJWT2CjVzsrBmTAAvEjRFYhcDXH5Zu2cqNblDGiTL17RNF/6y4riu7oNCeK
p2jKfkR0QT8R6iKDMZwiSHWRfoZh6SYMaOuNLLpXv53/At2rLhioE6Bd94BFHvBe
46AmbbuXc4ztmqFUEec8ebeJyiSjLe9luOtJLQXsrEf1fwL9CaiD6lhn87JAv6I2
zs1JBcjrrMsqFP1HVXM2VEBngtUxGd+ll9lCyQY5Woy1+CEQ4SnDk/uVRo+yCulZ
DBqB6RugDDoCdqAdRPewA6aucTztOALKk9PqRqBTM/eJ0AdkdGze59J9jReTkKXc
ywL76CmGaZvXGAhU+FB+P3V2yd3g/Nx4KEHyeEDkCX6l5ABy4oPttcSLglRDYUsj
VbKwlEK8YXEx9iE0mXydLw4xYL0Yn3x6WuSJtTyBZZ3PU5iONitiXEs8ew8e4KMh
Y3/q7QSBChYxFCPipEbr9j5P6dkHxmiYlHyKJlGOG35Y/zu8d1HAHtRnfHUXfG5A
77ire+hmHIwtrcnmFI57Us46wgYZIkuBuL6J3u44aOwY8zgtl6h1Kd+dapMUtX4P
0QtQOpwEsVr2Ltxs5f1nV52/7ms4HAsxWmjaYtqqI4YXLUrd7/sBADCZH+5v8ezF
OhpCZT6L89OcLr9ZEB3kbohKOuXLa0dTehgfWQnp3F3/1Fdc/Yvp2L+dmv6GNpLZ
Z921Br0VmCM4djrUXOM4kyJCHRE/acqdQQejmqn4Bch0zLaGmbDVUZQxPo+S1RqK
6uJno9eRfUGg3U/jxzRFj2KKK9M2awjVbA7EKSdTnruwvyP6LYV5SOHRMPnPVjuq
mplgusPW9ydDi2ZDi2eWCMwgtXZaS4gx1w128clDuImIUPJ3tD9dghB+02e/TRYo
g+iu+7ad1tMibmSWiwAzvQ6uVPNA5tw2DSxMOMi7VZ8A6cciE7DJQTUrmAb35xIE
9mGQ3mJFLKNuQ6fNiKx3bZKsojywBatWDhz+lto0e688hF6IYSkyO5CDUVmPitYq
hGXfhVVoPkH/4IX7w0bSbklrRgo0BfgO9KFZmkrGsG3iy7B3B5pH9zgV+xKRBeII
tF9rKkw+2YuNWbzj8MUyliJ+IAk+kUmWk3U4G6fAFxP4R4kyekDub/fKvSKHqZau
kVwxsTIujavQ/j+7GAgMUEjr5/vtWnorECB8xfIz/LfNhG2C3avLzHmtJgXqiUP0
rkcJvQ004KgXfITjVuoayo/Y90z2lWZN6VMqDcKWcrppZ9zEPfAwuh9VJr5FEskT
IyaK/XPsKPoXGKbKHFeuwNLAIq9as+cDRPt37Yh++2SZb/u1xk41ls3bBZVAoDNp
62LCiZVyQ+4fcBKjusXNydMMutjSGCQVpq4vYs6JJdWazb9OxCKPIyxXcZQ+pOhA
8pzwy5YpilCpbbKQkFqKkE+i7P+qq9PE462ZLUs8Prfz+fB3HEeFIwmAOpZotEAv
CdSzjI5yvYEzbbLr1MzXU6dfdSR7Qnb+BDJj3ruFdLN3ulJ0/dXZfH6vrIj5y0J6
TH2MOyRF6s8QaLmM0us6nFd5lxTVW0umEAnhXTIlL3FnYd6+w5z18ulF5eYJGBoP
A+I0KceeAvfkgdeNWXgNGqAZvH1JMxV+7pVkCIeb6NUKlsrLhAIANdyOFbi+PN65
1wqqlr3NO8JxSC0NMNboNnl3BR0tm7A6mMFbBtTVfK0W9BmLdlrl3YifXUEAqyHN
YYsvGQaqSbp8bMchRQNoSoA7unwf2sCIFUtUFt0nHzQ8vAra9nzAfI8bM1jyTf8f
wObfEwCGA1vKy2H0UP0KVNDbqMzyIOyd8CwSuDze/16JZDyR13rWPNUbsfVyMHdI
PS1jOHdUEGbNDYPP7VASV1Y3UswapFep+gP3s50RmlgHp0wAsU9PiGKSgtz3pxP9
aIddzRBfZqEonz0dQIXRbiFGBnEQHKPFmOzbaEYTapMi79Now1OR4GPsurPVRTfU
0qF0cHYxpWswHrYCGQTAArUpL7cH+Vf91l2e0jy3MB+f0r5RSr+3yWlWU4IzXL53
CNm10PAa5TrxczaABegecRMsZTcMlFfKiKs5z6ZzQ2clORzUPv0PT8Wlfvh21X7N
3TaIYpjacunzKR1cAnoSmVUaD9Q9ZenIkLRxJYgb1AuEolqOzsg8/WMr5hKJ/fNH
bc9L/dvV2bWtX9ZUTJtq93B0IY1bCpW/pnJM4mXMuaqWdhUQuqDKAiCugR8I/Yvt
v+K3GRO/BVD9olI6oR39PgNuELaXi6gEh5JIaSaY9pAz1SEiJGYqO8ILIx7RBlIb
ZOF7CzfBW495kE5TQfxtFIHZP8esoGlkpqQPUfMoWqcAnMcUpZGIa1phaxE7vSmb
OvKTqSzFXfp0rGBX07X2eNiZ6yX7nfeNSaxha3zRGtv7zTxzMH9PhILoFYZtUUdU
2nOCI/pu7L/dWo/v1aN+yDbwkmEWItv/fgxCOU7c9Se8L7xYSY/pMS30T2xSDhvF
qvz4OKlPbSCFi+3QQuOye0c2h8b8xBq4z71j1lrGu+URevjwiYtAn35XxKLHfkq+
Vl5qwbDYDgRSlY5bjc2N2ItHim3UhQoztbEO7y35cLmv3ztLoP4V+mFPZFf6AVXw
FYyy1YNE0fdqz4t4ZgMh8RFyuyP9EKQv+SjlRH/CEmDn2kwOE27LP1MhEustwV7d
R0zfyqBAWJ0vge7DlM6lSXrxsoRE3GVHj4CFIlMo87Z4HcHWYGxDrRvFtJfrXZM3
JvvXmfYgAgHi0XeH+RCrr9UUeykfL2QQN15ta5nN7VV9x+vzogZVUwScsZcd5x34
j0fyY4xCOoTvzK70jNLNYK0YMh4sSM9hPjLvhWc3it6rFt/MmaSPoWWv9MOnJXRF
u2If6evO3YUxARcE+dPy5B2Bb+0pG5aogF/lgCk9Z2TA/8wlTumh3S3rkJmWwm7X
aGw6EcS3TS2HNpn/5LINtNLe3JSStZKeFEtix6G50nxS6JOpeCq9Sv8wv602Wp46
L/zlskZ72cZLzavjyO3CXWK58nhwmlCSmHc7CfwOhvPPKHOtEObluRF8Xb9/oLQn
zGvrZdQ4vCTrN+IyaAhWUnuxrfTq6XX6oFKIsUH/DtHiPthcTBpSEtK40Wf//B9R
pb8jCwkjy3IRGfrW20cfK49mnZZy1Oytshv76BXhxGJn95p+ekGBTK78EP7hAQw8
ciDND0lkr/VNU1PNDGFYGosIsIWfAqL3dkUipZSAZC6Z1OAxbuWfuSVoecIDCc/N
pCnskPBwvz2fK6eIS8BXxbJS9hUXQSh31YqYJS2mfrCo+HbX6ZIAz2dF2DaHC9IZ
Qpz1HjaVQffcATmx6URN+HtPVpJkoBrdmxIlXTie28bI61lM7fYslEA4lbmXsfD+
Mr3S0BpU5BimpqNJWRY1vtvBMwqk3xQCz1VOrBPfjIDoi70cKxSgorqRKg3rVbiW
SdgfeMPERb6Y3iwWyBBqd4viqeTVOHEw054hjmFUmThkMeU+CSPPqHwVx7CjNSfj
bESSkgiTge0j2nBETO22sjzrZs2Gy6k4wW80kgUOHzRfZCPiKwfhT3w54fh8wrYP
Yi98TF9tTjIFBAjAnDtRgGnv2cOcxQDGvUEaj+6lCxcrTfjS8h1lhnDAstHno3Fb
M+FqK08J0bbO0CZ/s775lQLUHWfW6E9FkHaNkR3N8G5kNVMIemC3DRXzILkO7q97
tOysluUu1TtDJ4zG3ssMVNGx9fN2feFuHcbNlKVfck3bXehVLvOeGfD9LG97k7mb
8rhdd8dnVzsQWLP4odjA2yUHvRNWqAbgpMr5UCUw22XbziaOXGFjUIXaVooBbpz0
YyXa5Ldl4yZ8zB4UEGNduwsxjwZeSnCyGb5CS9NTJoC8B0HigpbQ51q5AjXfaaeT
lOLuCeMLbjnU+0fWh2T7FgmMHJW36Jhbg3tf4GJvgHglUUdni+yxDxgSs7UENPvk
VQfN/JfGlDsrFWUtXYvPH/41npjM1aKq8UVuB+agFgeCZMaDkynZvnTrd3Yf+EBM
c/l1BedmWtYXVxxBGxpgWux8AHTHf+jLXT+g2eoPnRjaHUwjWtMiHgu3r7Rl+9ss
O4QfO1kC5E8fk4eS0qMwJBMzNeQJwueRMLwQc1GebcJGhZQR1/NQFrd1E6zQ9+PO
UpjWq/FcbflKhodoYsIVlnyIolTS5KBW8z/io+eaZptkOlwWHG+YkHTQZKEXqsmG
8LxgV/TahzibShyB9xuj8byp/FMAEN9iwz8J4teVDECME6Eu4yuPBL+sKOj6T5AH
e30MQUEwJR9E+Rb/D3nkrnRLC9aNsN6hmcZlxsGqOQwO9kXf7pwTZmeAJY6WZ0RV
Sb8XCk5J0Rqbc5VnmMhtYGFxXgx1WY1G3dEJj9Q2mgfF+GiLnS6TNgaEIbBctUcI
aibS/DMzJzoniQSWUKXcGCJJLKGt3s24zDObMUrzVAcZD6RHbnU27Shi+btjCY+h
5AG4E0T/ieJCfZXwew3tueokupKMZ4IZebINsxugqDWTEC1KsGmW8bL6iyb8Csdb
/ICSTwuebuUSexmLSrby4soFnwlDTvQYsiFPhAAuRwt/aKo+neEHVQr9UY94+Yhl
BVJD6oD77+Zq8R9NV5OugWtfrE/QUkn41cZNAgligTY3Qu1ZOc6uQhV5cZWYMJ4h
rfSOOjY7YVapBaUsaTIUm1MlAfieuj143pQUWLiVUg9oc9D69Bsn9UJiWimPxAeK
pjBTSVf8v+od909rhs0iCPm2dre8TOU66P7Ah5E0RdNmBun+/1U8riodwzEB0qfs
MfBps2YTnUvCkp5JwlzJAKS/EEnYdqpzdwVrHmGNWKEwpkinhaD+Wn9IDTYkJCWq
mb3nZ/P6oE9/faQqMtmVZ1AhqrhMQXPW3UUUZPk6lRPP1Rtkq8hr8Iq5HqhIvbKs
e4ZiIB+uk/M0UFTkgoqqVoswyxkiKwjPbBC7ixH/vPVHjsRaa0WslLs67CnBllfw
/a9/2jakhFLu2yc7WggQXuWJrLhIB0oGfAPbF8r7Eh2KLvfvbo+RgEAHU/hXhiWf
J39vOaWhdSfbMLSArbGjluCwBVw3DBzxwIpOLSG6Dzir77OVegEFYzOJ4skQruik
Ifzc5ueA6BhAoMANPsJNq1YE7yPVMFwD1bth4Cuie3o5jo5kwtywCmNEl12s22FF
B40UbDUnBU6G3sF0aTB4knaCzOoXzFQgPohLH+vGYeJ6Y3h7aT4SW57AdBjwRUxS
WK5nZztZFDcPvM5/2z/uh/JsjJzxsQZW6tbNbmH8m5bNt/CKevNpuGLvgaGNzFC6
ejXM2wBhI7kd2DSsiMNvPI4AqRTV7JxrdmmWySRy2wGha5u8KsVXNFPhC0l49mzl
9Zw1TMzzMTC8kLn18Ruehxg19QOpPyp+VBzPe9gh7XOYUkMjBWmE1I1k+BRiBDuv
Bm2oJpmHzzzubJIfcoB9zHtq4t6ysmT3XKOMf4x4GT6nGtFezEFUaJL6V3FnXqIX
AOhPg8zuIYSSN7m5sHccSUvBlX6MoLur1yKmTEqY2rFF5bS6h5RBgkHzwhDUK8EF
rKYxQufDcgXLV1xF6bsagrjkw7XXvNf8rkoSeCouWskIzIZfeex8b/dBA4iRs3ZV
wnIriQunC91K6phsH0Jj8XvH2GvTOPzOUE3VUJLuf/Zf0SwYOqIJoBiOhaFXeQeY
R72qVvpgM3CUBTBRMOb9zuxsWr2BChTs+/zinf/0XIuyXnYxxp4RlEOMIr+ccVCu
bmO3iYqrruKZQYA27UCwM8Ly8RfUGws7vXugHf8+hvyAvg6MYj8rzIEuKA34KCxY
5wy3uod9YSJ1uYzUjygfT3GT761XWGlW5fW73Oim2tvuh8zChOfmuZ/hVjqhgPgr
nV29tbMQ01lDkuKgRu2GLeVHsJgu2NPwy5V10Gz3OdNTLTlprCg/oto2OlaPSrsb
ecG4nD+C5BdZIQw4UXXTg0zj4+80g7DBzx64SKfOZU/+AoQb5SdsWMjr9M4nRjyU
gTBnSU6q8+ejIg7btIe8NQzri7VIcgekHNgTn8YaUJhGDcHe/QgfmiVEt3LwZeyq
GXNYpPyEJ+rsFo1ArOWY4dC1TftfYxeXpm7YQpwwRXDXGE6Od2O51EWmi4thd6eX
HGeY6ZWMIu4e0IfX/w/Q4cn8J0pcjl9nd038/4gCVq3W3KN+j519NaSN9viRLuq+
ul7Dsga6aUbGENsMCV33U0ITN8J0IyzjbLAw7krTAjyqZ9ilntq7Q+voGLzc+Y/+
SJ0S3C2dpF3m2otxmyEeJRLK3dTA12I76zN/08RtbW9tzo2RT6i529NlhSRxteQ5
zN5EE+kp2cmWSpqZ/XtZAyPuO6+zKHhTlIDl2JXeA1CexdU4VJAntsmaaWmQ9XDR
iA2eZn94ZXFeRlTxqVULUsfYzu5s5CIusSoNHFefykiryXkNG7fTLbgHwYmbDtj0
DSVpqwVjX6j0vTr9xzHEG6PRzPhr19tlbZ6B5jZPZZBklFl3xy7OL0DqNEtlyyXN
JNaeUHTdo0KqJ9ws36CAMw/WMlLHRpYpB7v5pVe7LF5m1mhGxxDk60xxIlYAc1/a
QgQlp9CIViaRODwE38l1etVbA5rbv0k2oe+P2bzsucQPPZcl3ujclnS6mI8rebem
5mTbm1RH5ISGgg0FLSgGm/VH1Jj36io8wuTLGT2RtJbuKIBiU7GleiaOlL3geB9B
ogJF9dXiv0gTS6i5gqyDHB2yVvuX3xt247NppW0HXUnqkbpd+uIdWNeoiS48kEEz
CHOKStKwix9Cb/pRX66HkWZXnWl5acmI8kXxiWe8evicGoz0ivOi9uWCTszm077w
LcmAtLztA+cp3rXJHUopSyTNwzt7inJ6jT3O0glJ7Gww2m2T1aTxdWvQdl9VGh1c
ZX5W7qwuPIsFC9w/kjwKOuwUnbOJYZXsIHe3kPvnTw+qacKW3LGVFzQiOFuMzUDV
0HvklKzxgZoSAEHo7MXlHtWGfYd5TqunnwRQ7t0CBpsRW+JHibEeQC5A1/AN+3vQ
dLvf/Thc5YQZAi43Fs8+5tNYSsR9+BbNBDaq/M3RcktE7dcCKMAlSHIN+jb9pfvr
UGFsL2bcN9HBHxvFNyHufeFSEnTSXnaGlWZIetQNWPUGxWdIa1/xwfGIOw6xN4EC
2gjOxvmrueVtM2N93MCRgHBs5hKxYl/ORh2ZBGxcdIDnInCcQVhxoyv0+IqwPXye
pWNcbZRJWX0oMsIDXWD/6FcK9rvb2L7aexoG1bcyNvsHSDPk5BmJbqUNm4Qb8ZoD
438Lmj69Hm/NZceM43Db1SUZDq1xxJLXN0g9jpxRc1olBBihTFK9/7yeTN01u/je
umyVWZv5Vm0aKoGcqlvDv7UZ5J9ZH8vOKLEMOOwZ32/QCv8Z5QXigOvSynsqwCYE
HvNO5RCMW3HIni/7/EDeZpHURMe2yOM6vxR7QA49W7oeHnpNekmkNFVMfn2pDrUf
IOgiOGVpvVMn1iVyISsBTrf6YGWIvHD6iIOGgEYfy134yx3nEHWQUa6IsRGNoe8B
I4d7Eg/QwwRFiBlS8rqWwXYrQx2hkFUaMArm5QoHUQ3xuLs4RnQqeKQJrb+zBQnk
j14+nK1sj3YiULP9DEewC6wQCYigIcseYlifb2q58yxIPwwH/mwr5KBxYCXHyW01
SjMoaDl4tXCv6qiBQtNusKIXsJKNzefelvOPXCUa/19R17pGbSYAWxkKFtTXmfUp
XvTGmXlTwhRvUrT7jzUImFLByZYKF8NxXj8qT7VQbGzUJq/kuWKQ6WI2QElhC32p
uWo7vaLwro1yKRl/qV9qUYeyo56/IZsaWbzp26nxLhdxw9F+loP+0gUxJMh/FF77
pGWscep8biYrYnpMFUZb7xnbENV5FoRmzWHNOeCihmdYlBOGMeC4R30NeeZC8yio
grHnRg44SjHlFmRycOCq/Ww5Y6st0uYE2xKpCOb8yhQU8+LOeSorpmZDIs6YeABq
A4e0zalN9WDRAPxyRQbHY+4sx8WajopOQWJHfPhwueN4MhYuTLa1Vt09tr/ng4bT
DN4tRZYNrbKz2GL+Ogc4iz1laEAXdys8ym6Vu3qejbdRvrZ/gNIcellhQWQb1i8h
maRE6xyC/gIZ2Tw1ilcPLMZhAt9AAHKc4uEWMiN8Nvcu0BCNKIGWYCE3lh7XWkFz
dAm22zPOkdQlS28EI0PwZW0nLAwY0uMIOXM6RK2+J5WWQ9FVsK58qLUcMp/YH9UQ
bC1HvZsd3uQgGT5qJ53LHe24HyVrpigORy12p3cYTSEDXJvuBo+tf4YL+B2b0nwX
iniDY3/gYZY4d9AnscpvMaW3xzjfhGPnifFUcsiK3cQ9+XO6ITK/KsTx2AeZOe3O
CnqRzTm0hCZqfgf0AzwOx56zmx3FKQC2V6zXbMc+mCAIE4bzlp2QyvrykXR7vN5i
uPYNdR4ACW8orOQGA9eSOwjU+vGF7t5i8PNiiTfF7vX3B9ydu91PjaOiFwKpOXwf
UEWFUy3QmVgv1o/OyTSQ/d6gFV4H4R/sJyv5xm5xG7Ekj/X/m5wTL+z0LvUobQ3L
hqGkPxyVl2Rn88itOXRSC9JeZ8t4fiUGfhUhK35FN1ZoyE078jPsz3oesHwOs2/J
hVJA+7Dqe0vWwXqN/eJGS+mogqgW9QCepl+CV7I5PoyiVXLwOyOLsZ0mwNxgmwDH
UW4dHjjh+M7EGvdor3/N/f3cJxqoXlo2bASgYZ/CRSFLTs75IS9dbIZK0nef07pq
lHneppWow3+kp2GB13Lw4RlSnchdVs652eQ7hYS6QaAQVQYDB0fBfCf3ySQ6xAYb
8aD+ouaV+wajgw+Gjj5jBPRxYyaQ1k5bJUKGYpJ2ppGXI5EfQ/bwjJmT7JCRqeP7
PeV5jnV0bs3lFwUEPoctdRDUZ0lgKVKTgQwbhDxgxTShrZ7MgO9PvxHUQU5GuFjJ
0sIaTU2iNkjMNwXHSrkMuTnn9sk2RrLxPbIQT5lNSDu2Quua7EQL0fJa7VrwwNoa
ulVhjQLlx7VEk2lLjx+nCnICpzTnyzlVmwKruWjlWoUaakAwjEgjkneOwH3l485E
N/+/UskEjCIdAOoRCaUQYjeGO3408ZAlBhcMNU4yHUdCHDaPas1LRieGqWlEVbca
02EGK/D8JFCNVr7S7svUmUXqXiUG9qv+R2NQ3xniiSK5I5scg+A1NMUKNLSmK2EX
z2BFC7vEUbyiPHQkUT8X/6sir60nwcDxV7lK2fC66zPSG75qB4/B60qT8vi8Lyi5
OaP1HEh62gyV1sFOd0QqQJ4Siu945MLa8o+xALVJeeqW9THNBORWoSGL09OIIxKY
pUaOPBm3eG0DBSK+XZa0bjk07cLQL82G6CftPNMckydSluhvlBMuOgqBXHfHmGNN
b1HcoM41/gMY72fS+EY4tAS7gFJxNy46vlLpU7wUDUnsJs6p5BkmL1H+EQOBp0Dq
07e6x1ucYdmtGBY/twT5OtzLVPYl24k6AfR6ZaekcIAAV0xpsF/Q+roM0KZD45Ys
QarHpUECxa7q0jYPISAN6bsx60ojHc4Th9gPl5YnAbzP4CNMslOQ4nnlawXnYRXS
Tq4hy16Yi/Frv2bgu4D09Z3e4T0SL3ue/5ms46T3ESw4MBcR9dyGiCqVZASIKkYp
UoT1+bI/ylWCi1tJ77Phb8ORuOiTKyq/50mrRxedhT+EtHpoJWy91GA6G1Beldds
q5ZyAw5okkXQN3uDQunF4SRybXFw8LXzVx/Yu0HBFeK3krRS2Ln2b41wG279pROU
SdmwAZnXrF48YioHKBrwViLit2/BhnnqoseA1tseFbmxmd+nNwNc6//uJDpTT4D2
rxj0MqIdMPaXbB4tdpe18f/k7dUOFXz+PbsFMcU0PLlIM93h2HqpeDUSnOdc/evq
W4kSgQYa7z6uVyv1zuswEpDIpndLy7SyhHTE9z0a6TS+BoUBLC099UAWCDzBIfyu
sr0YhBr5b/TbKx1cDH/RuoRw1foEPysjnrAOJz77ETyCK8e47YbS+DbPFePRKDhV
nF0L8EuXj14jNuxmFtvF/BEDPsAdva0l9xB2YftBE5xulUSJpF2Zrov8/Io4msGA
WlP//eTDqFr1iylcfgnOmo7OtZwKzsTbtOMYy0+e9930rqa4Kwr1upXynTRgnBhK
+DlswGRK1KEri5eFnLNvggGDmPCPJQGK9O4xNlPxVX6uY/zbEeRLxQdUcDQivqqZ
a2YdXvgsPdHLEtRuk4al1zBEP3KfkZkzQzHoUhbNMHJrSxxSfugDlckrwCilPjN1
PLXxqEPB8rUr+tGsu14iu4se65wzBr6QkhSzPLMxP6lsLJKet676OzX1bKwaWO5w
jNrRkP2t0w+8dZVUZLJWpto/0Ss/muxi/hF+EXAX4/+QAYs3Ioa2cGL/WNDmdl5+
MnWguyN3v3gwKRSLtmiRd++98na9LvLz6kV++JiJ7FEUIcc9r1Vyw6Hvd/qvsEyW
nyUbeRG8qeOWK4ER6Z9SGRepETYfyhCK8J9i6M8KyhylIWqrawMjmrs1w6uT3xGS
QpFRebMON9NZBEl68kFb87s1kfdUhOteq2hqbCa6G/FNtWkwEtookOm+6oks5fgi
B6Magrua+TLIgBtP4pE2gJwtnQ0g0MdepcVub55d7pEjBXxvKKWDS0kT/Y13tQq8
zckPYZtaKLyU+5PEF9KEbz5DcCRAw5bqyMB2EkyRs6ifQdQo+qGO7/hgLMV+KHzc
/Pk4yhFhCNxdF6J5s6eALRuNWnBS1ofg/87++pCRVYCPFmrlzkA386jIXi1mwi23
inA7HM105yEobn/O9YEFYLITM9HFlAcoyV2VJ1rLowPYrARurLOMcwJyHhIhAN10
qRGD/KY47gazR0GPWzZ5oTb4asDKigBmmNXKG4j9ejsW7F34iMxiEmkeAK0gRlgJ
asG9lAmP7PjYn56zTi0HXNHXf8VxBS/uSXlGiC36KRb+O+TsXLOIbWJkPFBgcG+Q
fWXzQkz/QwEd6WMGfJG29Y7XQECp0iDimr4tup/PEbaTvXlzJfnNviR3TTJMuBnR
RTCXOsaj9Fc86XIdTDKnD0O0aSm0yHO+siVDSBVGaO3z2yjueJFGuHJ1KfbxgUFw
VwwbF3j5fYuUCtkQkN6U2my+VkLvMrTDStJvjWszI3NfbnujfAweGb7ep04dngQ9
4uRk9QOogR4EDAlqG9eUQt2FKnGdnXNMsdYRQGVLQ+tnqnP+FHh8d+Lf++MQtcyn
1yAlBCLm3R296JvO7R3wmRzvCfHi5sIJf0p4damc9PIJWzV/HbpNErzD2xiWzIjf
6SX/HntljMXTTj7P43NkJqH8LJsiiuywmHdLW8lesbCib1mxCojimwJapXmXdFgP
UxoBu1t0GsWOYAW0mNwQMBnAoVAUVnXJ6nydY4Uau4ipQK2PQ8TMrfgoNiFMkYmU
XkEManj4HOYeEZfpazx8KT3h6lYTrKgB3e7VnwXLFgpxWREJ5NHcbB8UNxGu66MF
/3UFeLFVLK92AQqpcgxZHTmtiK8uAbiq90Guzd7W2lGCYbftF3vcVU+bmF2L9FP1
rNf2stMbiGHQRecpBuTV2jbIRSU99/AQGD+MTJIKse0CHppuIVHYNtQQ2QIPZxJf
9ERUdQHIIuOM4Mj2omV7lmVqAEmMETVEd1EMZNR9SLUPBqLe0e3mZUhcDNnxlPki
MLgRYk1OcsshBeQuMUBBJo16lG7Kbbn+5YtAUA7JJLwDe0yad4w8ixS50xbLxTqf
9gEEZDCgg5LYdMdD4UKgJy80OflaOXoKRLER8Hc4vzWAsPgR6Pwr2DLX3VMYMba3
0csWTVFzvbd7VENjTRTqPtP7elzsYCq92LOhO/A2Oszdck+X/7DIUSsZqdjEWTsL
Cs1K4QZKY4zDWZEsKvB/l1pdV338G1erliNq5e2poIQCQyMvSszDvqPGe0xXlrhB
wOUCBVEZoSkpk60cs1I1ulMcg2ir1or83Obfvi71Hyind4my1puLiQId/y39/qqM
+coz234YTnDQxNC+Ta0zZEE2c8ZT8fLaXoDOXZLz7bizTH2SL0NnV3JmSJv4UBNb
2HDhmUnTNAy4aAMonVyxQjMKPlzRpgTuiUqWP64NK2JFqEX3wdNe0bdr0vtymIOz
FjHF6p1NQ9TFV0l+g9+7G0KURVDizWD8AAODblhD3rP3WI/0iiebQqSv83jN/dUR
W4EihnKp1Sj/0Ats8XE7hSqAOMlEhfak1BcbAV8b7tnxFGbvKD1oWLjpSaOMXOXn
jprHXWM/h86pRqaNrGE2jrITWtVy4XGhCUCL23hLq71w5SvVrKa5nWMykPs/HkQF
85FKLt3uIqf9OTzZ/Kdn/A6c7SQmG+y/MK6wquaPCV/rY5T4fHwJ1SFCPv53AZRc
bmr9xAAsbgdKEpc5y7Q/4ECp8jGmlbnGE1OVJyZREdS2JYh6a5z0FhOTXr18xnR7
+uIgUtlQqvOgZgFFUGW4N4KV12r7bxpUseko4bLVmbGvHOiyM92XH/i/wIz+naxy
UCuSxIoJLDhat5PjXUY1jRdIDLh5nn55bTZoqBGq33Lp/bz2GF9r0+J0TLlgmxt8
HxNqzAqm905TxRb6uNzQ0Yi5spuhXKO7uex1sc+60TDSJYaj/LFu3PQe4f5sQXAy
4O0LIpOBbH8hMBMiDBqN2qa/lgPTFHwfZSkOlqX43epy46LreMiShNfp3ssfuDnU
gHNc62S0JneRXLAWA7rOAQFsjwL88tWlLfDkoXx23tqWp3o5hQM2rZ2EnhBUm6J9
lXIDsvd1cNeFgal+Ds+QmPOn8qbqCoXpFdnBwNVpSxxqAUN8W3RTZopbWjZAxand
0sc0MCew5JYPVKCGsx/bAFW0Cfn5nS/mBdBkO9ilqgfyGpoPHgvWL5uS0WArTP4A
fO8Px8n6+a0+Tl2FoVu4E83egbeY/5x0+wLX8o4p/7fY/WN3UEe7mFfwvEYVx7Ua
L0vF107BqUtRX1QiZcwnDa8o6F8/gDxRUgDQACZVffNp8IFY5krKazAsbxTG91uK
v8arYMNvTtmYBESKVzlRCPIaqL+TiTUR3+sXBIsrlg6c0JizZyQeYYyLNnj7HIik
RomxIlRguBYqjlUYVlr3lxKsSWl7ZUR/MSr+C1Z0Jwvr5CnNRUEGzxsgmeaHuf9J
Q2ng1pu8dtipxeoaQ+w6w6e7hyTpLyurJ04ZWXUfBKLfilhJja9CyUkNz12ugKPU
A7/ekzV9f7+s+MYkPdlhqPH+FMKvwqie5Fsu0uiUtHmAcyROryCF12XceijM9G46
OsnqRJ9cdIkIEa44ueORcqfCVNKZjNoy/48Ntyow6vEaqyVX1p8IpZ1WjveYtaxM
GtqD8jdfC2y65nXvs+RWfY2B8eWjsX8ty74B4BQfqEy2udaOVydsmMc4LpIk6NYm
e30g+ddNtN4c0ewiKHpYRd5YGcF3TNVP+AoC4ilrbpPQ+vFZ3L7C4QaQhO5NWS+O
R6y79vm3M8kUuPieNRI2SzPNzadh6I/RE5A6FepB8VXvEr0OrjJkNdN1RsR7QP/4
f4avfDkAvb0QvIhANcTSUvXXBQM7UM8IH/24cP+H2jPkUBTk8rKTc18k3YAlzcAu
jHrRNYgfqrLhKAyCipvI13T9zB5ARheqGW+Z7WPlmsVxI73LdlvnB/Mkp2yAW8XE
ud7ZuDgnyjp2ZFVWGBAeebgaWmxs14ztjktOw5/q3d4z6Gz3kCXnaE5EtZ+zIute
GiqY7C0PE5LhXG3pSxrVjoEF8X/mIoe6eINF63QJvAv59whz3wPccvcus8YFRgOv
95aFzQDul6agyRZnxAVQIx8x54ET3aXyjksYL+uE4tdZd8VyVsSbVwBABHGG5HTM
YyC/VUiXJoGQTC+v4aKQapASMzMVhiZCyPOC3Lin0BML2+HRs1UoL6afTe5J3PLm
AlE46kgHZC2v8k+VGNITibjYVY2JRBqRtfqoJplEo0z8WQsLhg4Pl+WwYOA1oqIt
GIiZhYHrTmAqmMwnPO/dsEYQjnayTMmcpN11h+Dqz9FG/6PVCVwa7EkIdN3BfGNM
XOAfQyQmKAgoigg5bDnlbOte4jOxdqQqSsgy10Ji6vc5EzUmGNs6RVxkZ75DXD1p
X20kvTuj3o7RpF8UkPMFRckqnOiXPcBWf7+XZODJLR3vF7MfIdYr3BvuzRMtkq1o
7tf/LbWiVyA53MgkZ3nXKpJvkkPMt8nn9tEBkG0R6JtlPCmx05bLAV0I6wLzdADf
CUz4Y6AjydOSbwIrHhXCyFI7t7UB01R1/JYt33xNVIgRFO7/0YFE97tATZ0IGe1m
0wlEZSxvYmGaIdpQ2h13KnfcfsFI+MT06Q0m04BJhYZpBcEEtMF1RQ4OEuK9u91Q
wPZkuzE2Au7CS9vuQ6+XhKdyA9T9IM42BSgjedN5pUR6d8NkUc33kuNhzq6HUjyd
9BxJ9fmYMz9GP45QQdyNHWs3cLhNcMVv1F78RX5bTAKOQWNPJSb7BQQcy1zIciGC
HHzuOiv7pPGjWgkcjN2M7jkTeK2Lm7JgqkP3HJK9OBTtPX6n9RUMeBtijqVe+2Ix
jVot8rU/ksQazi+bvF4C6l6aii81ZL55cDs6egXaFPIdqm/ulOTKQje47QTP+nfi
iga21bZXdmK8pZ4o9LHnleNqe4AMEtTZri8kp64j/L+qDYEvQBqFOITQf4S0AS0L
ajdSGQpItJPd7mg0n6A9okvR19QKQ7c9OCO06Ldg9mPgp7X26cRl1BBRtKEmOrcC
8JHhmmCG6Pg7CVfZzIXM3pfdgo/oXO0U/s3MCh+qLDnj5TtlAK4e6/T/bK5KVPTp
IzePV8Xl5mkAa2/QD2DTngtpsE5aWFhjJSRiPQSyoRR9Qj9lr0Kn7NeB2WcWevHk
QbHXDBvsF3s3raHMZjzctrk/OShSCF7ZhQpsjV/WV/+JfRP5xDGkHZ/tYhvjDX8c
Z0d8+B9EwuHMSvXl7qyGSEPnCQ+Glm7ei/xmOrk706I7CDufthIPhlh6IZlzvLy6
DU4uksAUyTgCFpA6WHvdkrO3DkLMENkbLbWMWRwxUBoxC1odATmxmRvXZzJxSKbm
QUG5SyaOk9sccIq7FbG8xhEVwjfD//cWbPGBxJNd2vSdq+KKyQSjAjEqppJMxs2I
2ELBbQZmuazrIr3d7W8s4L9kQbgdAjHqBR6HdWXtx7EMvxr+/MAq3hlZGARgVHMf
ZqaBcJfRgBO1b3SZBAkIsCjDwA+ToKwhDMb1I4Uvk1KLpdfqrBtd1ILC8baUBnik
0ILpIYE9h56Q1L5GDNxt5sAiQx/qGZ9e0jlfDX4PBaz+R5lVUz9Ncf6kf1fpf0bP
SC5VBVtJAYksxZPCqiVSGLl94Pvf0Vw5iX6QmRjszFW65UEdEjkc7CHWuVFvfSfF
vGld+a+2s9ZH2axg3B6iVhoBJmwUUlhotUFoDVHUU9O3DFqOAl0S5WGzxJnH44sy
0i+qPrWgj65Rt/nG1vgiSjs88yCGu1B7ilmv+jLAlQAP7XrQ2nHaskBSXsxb7xJN
MY037uFbFg4o6NQ1LlDODCCkMBV7/HeV2Tq4NrbXkU3beKAiM5AhqOb46gjIFbV3
qHjYm+D05WtAqR47kwiN/YJHQLVLoZ8Lzks9vC0Wt9WVoxI8wDBXezu6DsYYwqyz
oi+xwC0RUQdg4owWQMKd6wB/xCxey1qsxcvi4KpGMQcg32nf0g6vEZH3nAc31wOr
CnmG9Ihqrp1iy97TO9NyHzlMvJhmDJPNam1qpDpcNuK5lABpl38DsPOsNaZ8z/Pn
ZPXcqLFzRF2shEs/A5Tguq4FEMwRY+Lv41Rj5PMs4Qzw1Q+OuOpvW7rRrJGRfvYL
7RMZjdeCeAmbwcggAyExSFE7cRn7Tt+0E0hRA7awS3tGDchh3hsiXEH/oyObYqFe
JoQRB9WKb9hw/eYZQMimqVpfuO1P9CQ335V66OmrKB3MyhqRk0y0XDQiJlgZb0Ft
Vda6ibaX+fWv9+HB009BRPDA04sWwA2ADCGRFKTGM5D8OLHdbPCWGN00I3u13yyF
+/OVPukavq3kVv6B01TWLCkh8HsC8ZQk7LgXLD4LcPrJKSb+6eNyWk724w0V0Nfa
KXAlLxedgE4FxX+CwnOH+gWWn+ZVr3zN8Z64ObQnJSEmqdeP7TOM7Eu1aEylpFY5
wmDQp3CTPlOnYSWfn4q0G7IT+6DmbEyDVolmHPUtknkswF9RMqHXlULgJJ2+YNar
7xvmFi076BvGeRQMIkEZI/HwUcgQ0UoKv9dX34zalYb1WD2c9ijxB30J0irAe4/H
wMBr1nh4fzNg1PkMezj/DdKdwUE9d/zGz2Pqi6sOvFrDYLrw+mzoGmJfW/oJSV8j
bnDZhYqJURQQPdUbPv10v7U23gC6mBLf5UbA2OA6wIowmRCxQhmgFn2DuFRPOEwT
i9Y9K6MHAF3S9ygLYtPdD+GjzhX/rABjSBa2503HvelWNf7w1E9C+D/fQSw9YzmS
SpPBSY4dgaeJSESbVdyjaQa/ZocfYm3HmiM7vFT+lFK0GlC0cuTFyUOviiczpy/g
+89S9y9Uk3/2QbxY7yp2ZL2cuMsWISI7wKeRFczvHdp2TPiEN0R38I3jzW0gwTDe
BCYKA97yoMp3Xvl35OTTmgzJOSjkTbj8NIyTpilCQCVxZsXcrRPJveOLpSMvgG2h
dw8dfjO1d0bTteTc7VYb9d8QuwtOjB9cmwVPkY0an/y434w6umFx4nRpnY7l0hSM
g1/i+SNnRD1CixcIwDS5hiul5jeTHJu67jqhKwMiSmfNdE/wPdv3VmmqfheYtQ6i
dRDJUxogIVKj/e6sSbRAycme8Erf0xcpzSaY+XqS/HChjX0iiHMBbYveGWBsWh4s
054o+55tM4sZNy2CUU5vZ2spR0uATQIPscRvP3UQVAuIBk3WSzSCZvLeJete7dXm
FlpApaT64E0DGpJFG7mVBDLcODooQbq3gFYSPl0QUl3uJV0bQIPddgKPSRPsUU0n
icmaXMO/nRE2pZ2qj0T+HBXRcCCgR175xMbo6/oKA4JOzgZvN99p+iLZwFmWsmeH
I7zTmxjnzw2/T/hYjBkKHzquyzWLlE5bgVJ1ZQm64byFEP5WqAKEwpVQpCTws0xl
KW5ucegkrDBydlrIlX+JgEACJVw1ZF+x4hJvfvkVsx9lLBok0CAQeQvE9Ui4FUAS
ljahq2SkZtLYsGbWJYTPT9qnXAitZSBrxR8VJtsfaTtL3bec3R3jBMsHSbh0XmjW
wtSkiMw3RywHgQw0ltqdLQpYUxQ35qz3tTeF6Q4otbQbUupaQo6YSKQuPsFhy/Qv
CfVDgZyDHfre/7kvtj0fQbcyVl5kHgiQqJ9jj+W1bbzylJsoJc/p+C1CBK5LdEF+
Ea2DaQI3gcPhJLnYLfrpJiiZQQ4KOE5PrEB+ryzyWlUQh+LmgPPpMjrNvcqwXT4h
/JdoDDTP16I5RfgyuNts+GyYG90WAynyXxQ7tLg/ENY6XcCo0zuNzIE5Jvyfm+0X
imUh3Mi3CRip2ndwGXfAo+X6sVKNmna5HXEIvX9ByXIvv0iy9ghHRykwUL5k/8Ia
8xh5PnWp0Av11GV6tt9zqeFyMIvPi69GbmT/DdqKUUMpCteAxCZxnqWPq6EFY5Vj
lpri6DnweitFqSxqlKdu6lnpHydEkRZy9cf6RPJ8c2xVJ3nl7utnipKmecBMRs9A
l7d/M+XTwg9LfbDgKmPUvdMMJWTxiOlcbJdgzFF58St5uxq+iovewIg24A5YBTvO
koItD4ZmhYhvsYxUbgwMZEPQBjNeRE+KeCJtvmcOUZ63blf/hO49fQKcReTHEJlZ
UgZdD3c3VQO03fR30RVB9c1+wtBUnRw5AAnj1XqCbEoAjPtKq4m7F8KVeCWGoqGC
FFrFGA2tvcvT5tVLI/tJdQqxJLVkLAFybA1SNiR/S09e6Ag4Xi6mGASqawSUdphP
9BoXr51D4DhBpjGcb88cvNAl73lxI048YnD4IQ4TGlhGTzJlAF9cK0O1Wgqm5Cv3
Ne5eDXgJ2M/QpqMXz+dkXLcF2XIUVFcLEnT5+X0alkOi0vzatVl7syH5ruC73fVS
FuVru7wySqNGThuM736pF1VCYtqU5iWAY+3iJFOt7tbmxNotDgX7ilrCi1T9V5oT
KgQLuUtcA9qjylwFa8II7GxeiXnH5GqHZW430Rxp1CrgovKpK1dKYn/GHbqLESjL
VdMH/Ls/cQMsITucIq5RNP9CjTe2ZA+teu6jBwr3VoXw5yr6w7dunyox6EaKYhH9
Sri2c3MgBGO9Q4bUe/9LuOW8LPnDWgowRcLRO2eBJuePq3WcF3YfqwzAXbtgxeLg
UrsNOTOknGp/n/x6l12TvzrrqNR1HVRJnatmxTGNcEtT74VDX6F0pr2H7Mk6Bi3h
rjVXVx1tK0cYHHLhWMaiHpEcGTeJwrLmXec/Wdu8HVrC9ViLaM5ojo7PMHYdveNj
E6wZ2q+mbqcUNgZl/ejLJHJx1JfSQhCGJZWVk/+bnoXM2QXVkQLHW5eFwfWcopH2
CDJ2jb5p4B6H55Q6ia9M3wnYqjwVYk0Q97bMmTkluNvbVwp6koEq7qrzoZEW3QOT
0Z7bfHeAwqBBZhFOpGHgo36vpv1XObYJ3pI/mulMK/Jz80i4rMtuQYNIw2Tt7yv5
FT1JVuTRoqhZHfVAhgXv+RrC8sSklk/aRNgwa7u+bvzT6qfQ44TuWe/ez7UoSe8r
dc7YozQwy0wrzCksRec/9eiaFqD396ns+OmZPBZcCmDGpMTKpNu7ZWifj2EXbclG
dGBlBo4h1OHQyXFfNnQjr13DQiEF51xurc4dItPAWyudF2ehhwQTaxZZVay4BslO
9m1LcC7JrxuLa4YWzpSoqJZ1wP11MyN6Dng6SFRxRbsnElzyRQk4B5/F8XTZR5k0
lJKCGG4uYWcmfyFNTtCaFbhICFO6lys2Xn7nvx3ew11yA2d034VTZPQr+3Tr2UJb
2/Yo3pNzABZ/WEkhXuJpzXOfSTcn9n3RYhwHbmnKI1sBWWBosg2HeVm9Wye54JGp
DVHnx4GlSgk14mMHF33xOqaCqpFNKIb07glsBKWKg0KoCvh342t3nLGrEthcPy6e
+7f5JPy26mBHoGhtcms3yK0PpxhRCXiNy1dgNNFO5Qqbb4zMyQVXdex23I5Zb5nZ
2cppNaT6Wu7RpOSGw1mlpwqKgYq64IBEvvEzpl+qBjMeppQFr4R4xee7dNZ2LYuG
Q/3TiIxdDmcmgrfV3c+PNtXDSVVdn7b3H8lvuZ4xlh9Z+8kDjoXjWbvBylMPjHLK
x07xLGRAIyCztXgy4XNqlSqUl0sSFau4vkEcFT9lhu+BnzKJh0uuFuE6zR3xEhrp
INB1eHEjLT4jsyRCIKHNUNG9gFJWtzVUEaED+ASX7kvfdRBhlehVnGDq4XgSy7Vh
dG6O6AzOq2fGXNw7LCdtZ2kphTKfG4efhI7o3rWzPkvQEWEWrhmmwMZ0/k+lXCzh
ST8HCvM/Te+moJZyRKVUe8eCQ9X4fFT8Q+xn+T4CwKFqGweXstFZVDxaeK7r3LAA
gl/quJdQZfRP55aMcqgPWNWRJCAAjnfAQ1+jIqj3SvGI8AF6sX8zhBhN97AohIL1
epzU87gRYf5oElox/JCtiFcooEuLZfkekkm6jE0Zod56KDdsxsnuri9qcfr0DR+z
jHQCDIjqucG0WznqZKK7lOfjvdhrdf3YIpRzGaDvhxGZAXuQbyRY5n0Z1bLWlDhJ
Hw3HUzF6sTeE210zrR3K2sK9AHtyRamRCIa4fCnFn8extoCHuI/6uCHRJIPCAm/E
OxOs9vzkNwiv6V5YjoEKkKs+qjUqbRy3Cd3YcOfmmeNPSprEB3ThiApbdV8uu18l
fxt+PGv0pGes+NY5vAwQh+Hyx0On/GpNjFlWZ3mcEW30AAM2lODzHdKoBX+57p1H
/h47KBOD4vLTvaTQ67LgMsMX2u+5LRvQ6YvvObjkwbG/Zwyu7TPCgW/HIBl5Y1yc
z3lFldDQwxSxGHLANHeooZV1qFXabq2lrgLOXKgWsqC+yosrio9UXJLCEMpMJG5V
VbjBZyK+EFAaIz4a7FSkuI3HkdZ1tl+4YiG+Q6qdW/+ra0l8CzXNqIC78aDHxz+A
7v7zYNzqNYBXp6LHBpOT0gom84ngNSA7JQmNbp1LpojPV4qma+V9e22QzsiuGUyg
tF/jbSBgT1uXsh2Wu54PVDqNcBa95kdAgvmK86D4BjppfNhZpDg7o9WRCgVakZUa
FoD6g2mQSdZ1/+X9zSnBjahURovJnqaA4o8ogKGRSljeye0VoYxzOgwZ0JKGHO0q
F8f+plYaABqIkiPSxPQlAkMv8vJHte0RUrPDZGlqX0HHqQANmUwTtxLs9wsMrMUi
ChVtDfHJv6mhV8Xup4BgHT+E2cWRxvv7xAX/08eznMb6VWEGvH9LEkxdygivH7YH
2F/G9cP7nlcElvc2IeQ+AhOtYZvyiaqlbcVbLTcbgPwAlwTgb+6b1IMOGf/Aa9da
QaJg8ah/piJi+qabdL0O0zt55+LqzhufmOteVOI+szUKWQB+h0AV/WE6eZ+9y26Z
W62o85VK2sw35K1FM5bbEkGM93gA0njZhZOSFlGR0h3ovy3QXnDU1Vl2r+WB7vVk
ZKsb/cn02TJYL40lMN5ybjxO5GYLRWenhwHID6CzN0Y56ghx4nsgCM9PdLXh78lx
O+h3Ev5U/8L+gn9HidmwLcZWY04IiMTkFOzAQVi8btjNP9qaKZ481tZfWrpJ2Ebc
W4x9mE+sQO0p4QlD6RKuGYiVj0W1D4ljpD5YACTdCEUje6Waja7P/hjm/G6SWuZ4
Xc3rmglmmC3SKSw2txHJRkhBSGNYrT1SHCKgfubN53oVIhVBSB5xQU9Pvv8omFTb
9RLxr0kTkK6sUybF3uLGsp7Y2fkmxEE1ScsergDlt4nH+MJeFRWW7W0MFvQ+bHWk
m8uM3F+aKAu42dMETmnhMe80h10+mNx3k6u4WxiFSPJxYBUde5ahoyyHGcFMhepl
YfmwYEJ36mdgZvR5l8UJrK1awi/Lack0HymOni4PZkjWuxcgNyzI9+2g3cZi/4d/
blsrhEfBH2IZruNieV8jKYD9MoBo8W2yNUHypxJHtWyVWJtcidSLjmNvaJvP/+4t
Q//vY0UbB/T7Ky4vH82lCds+Qwy0Z50oIFBB/5wiaivPlX9iupM2XAHsmeh1jFtH
O0y0WW7TJAOx3N9nwJU+BFrYnw/v1XOlDjDfomEn0XDNWmMm5tjbRgHU02jRX+jo
eiQYQPVff1jgraZkS4ChsvtuzX9T28PcmnQgdazDKNK1CAH4JF2GGK9DfwbRwWX1
fVfzXlKuZAqBpVj+UmInDZrElOIdzK5qIt++S05ga82vClEDrXKrJMhjgvAcEbIe
SsVxmEreCM890bcivjT+JDytSziapfRiNb1HGUaQ/snxtel6TyBiDQggV1e4bltE
jFY2SgFIu3+kvU2ewNIy/g16BVtMpJWybBGywgyfQb7FahBWRiyhrnUhwLojeV4W
GcSbJKjccHqJ4rRe5oLIFbEwZTiee11C9BlmlCupIAps0k91Copx1bssmT1Yr/Me
DTNkdNY7xydNPnV9TmR42aXn59fNKQiJW9K9rdPk2KD8n/hod8GowN4Te0HHPoe8
0JgTv8IXz0VQlsGH5GzBzOaoNTbkKSNDrrlZNXf2CH2xSzCY3lJlIWbDrepxWlv0
0/vTHnp+ZIta87mFHa+iSeTDQGN6RMfOQSgNeDMjgltlOiGZ4teuBLAXkfN8Xmd6
SA9onh6bYFZ+XLfX00BZDmlo1QGl6Jf+aFQ/iUAjHJN3xOyJHsy79FL/75ei5LUk
PYWO2ffNq2HrGg8Q2scOvn/PdKrqNSkjtx4crQ6kUfNhAVw9y/VGo9QphhZt4a+x
GEi3kI7Ah/4G2F6L7ndxTIdPkJIh9CqLT2KpSQrBoZYks1z1jmR3cJD541nFHi8R
HJC5ijPMlm1p2v/Z8ckLvY2OTdfRZbNDUMtNXdqLI52JOwYL4vIkco/Qh5BRKXij
eh7jvKfFHhT57aKhpJDhVuW/VvMdAQqsWnO2bl1dm7dqSm/hUw5qclzblQ5d69pn
KZKzlz25iGjx2gC79yoBQqO2OEhYOk3GV2A6Vliu80CrvEnHBqyEto50rrlsNQGz
kLL5l+fJblhxsiiraFoHKTx2nCJNTvUutZESI6inWZhpkOYb09bfqcVYqlpBVog4
Z3cQ8Ezj0yFb7wwDFWxEE5BGNkdQZgn7Ysq5cMNhIylKSDc57eLwvZCaKb3fZFJW
bUcE8f3MDWKC2D+1dkJAUi15HEYfeq7/Eswl9knRu9uAzqseavrl/St2ynmKnVEi
qLYxbkjI+lGnRGOg5tmN7VPeOSnROrfdq7BP0/mtqTwyn14iZrb3eKuKQ4HGaMdX
uLn9jFSuH212uIr4/GcYiUBcziChvR3ms+LwfA+6YFyLDzqQ9Ep/XS/VlBs+vhtT
aFXndQdRtMRP91/ruHiJoY70Xs4Xmm/XKcOBML1RanktHByUTLQyl45Aoxf3nYmQ
XRphYHEmLPohF//6RDAiYS5MuMSvVKf95BDvN4P04oT2bcZteYCAZtZEPW5Oh0TH
n7D4+nzWpuwt4goaypu4VJs4a6C69o2zz0bKAcrlv7HsSItbcqYzO8I85O1l4WoR
m1Hd4Mux4y6LzJ+9+v88HbPdajeyRPe9aPBu6x8lMRazNgps+AUz+M+MUZWrM0zO
RuEqWDSCptO9R6f97rqXvlvQwBjK+gqsAJsMvnBo9BjAdj93NDy2py/cRrbBkWMu
GUpoA8meylsQOdibKQ1qfWmTHYQ7YhNyxToU0nASnESEAnlMh2llSKHg3waMqC8v
By0IRek0eowHkUSMQn4Gkzy0BdFWI3QuvOQPwer+Xi6L46tdl0uPWU+prh0BBObk
hVZVExY59f4Ic23kpgUSa577RwpiR/dPhGzZN9VIQnYdZPy3c1zRXpux5hRIV0CB
gEseJ82Kh6n7WjLk1Kb+bkWNTJtQonkCoQZNErGFA3WVWjyPd63i+R9N6SKLfQyP
Kjn7teuPUhwX0/xY6pj5y/xhI00W7XQZnFQPri2cvq+qevA/Glt/Cs+o4vEF3FTM
JQCUGf/eXWdB2pU4BoNdIEPJuYTbHgdTv3sMTlL2P1XFYbdEOMXN5t1ba980t0rn
zKxW6RhsFt1blF5LiNafPQNSg+PhdHb2lIBrHZTXbxrQIZ1RTny6cN7z2ckzKd3U
ZwdpwK3FjfmdnyMsKktvBJr9rXlv8IUUOsPtdQ4cpfAGsJbZyiqXBDpZoxNQLkTO
iSGpM9ST9bs92Yb/CKqnK5DX0ymywUIyERh9NwwhjiNu8XtldYfn8fBcuxr9+uIU
qmoL8KMiae5H5wrsZ3scpDw/Mq+sBbOOuNLKnUZrw7f7PMPwulR737Auuea8vX+3
dFpxE/H3QHW3WBxREmqr8HZM/66t3S5SPIBh93VEflkcVM51Vql20W7nAbTco//W
eI9gXiRl9S34US6tkzc/UhyUJXrK15zoW2rF/Aq0XrlmociFGvktWEQFklTmp/vO
775WFjYnZL3UoQ3nhL6S46AoQPl6zcSkTonNd+BfBIFf/sve5eSbVt8sW9k4CVQX
8KpHiGVCniepEsFZIJwaBv2IpdqjeLfARuG7KTBm1/cRJF1C6GTaJN3V+K6x6oiQ
tzZJHMenO6X/UFFg3wE6PLhIqtNUi/EycRdVBu2mDWR0/r/K6Mq3mkN21UOPeOSj
JA3u2m/HIPHFU18aAeDuL6nnpJBOX9WiywdREVSJKRnb/U5Gc8KDnDTW2QGPe4p5
81lRy9fV33jC54rUsJF3ux+fX3J41JlzBjXaky5HdfHIRlBzDPTSrs+tqfb4RK7t
FKFli7WgTcWTw0DvwV197Cn6R7du8My+KgWEMyIMYrFyWibRQ+BWHVtYrXKuF0ow
09aM4MHWXFxa+1yHyOcS/HZiE+T4rDJ+oS3PBQxlZch06Wgc9VNk/fSPfYBWl+k1
kURZwYFHQnRJKyJU6AfvQdvXbXzHe/U0WUEpS8uOz5zvq7dSUWFeiPDyfao1E1D0
w6X2NNp1VQcYYKLui9qPOG6ErRc4yNYE8o3d3880E88Vy5uLKYU3hFFHnKj2PPEx
BWWyS6N98rO199u36Hv8epZhNCya94ru9ifF5xwurAKX/W4QeG+TJbIrD5kUZKeS
Msp9nsCWSCL0KBcsyWD3UZIzi7HpUVkQ/P8xA9P6KWJ4WcJZWprKTSuxQ3dJFb4A
Fr3afo8QAa3pTH/j5QlNnjdxVVYwScMRJzQmNYbVoeZZFi23IiUF/JfBt6qu1MzN
N+vk6kRh9YzxpX5czqI//+Tp75b9Oz3kP5F5wmpAhCdyFj4icdLaF4fZpiiJ8mI3
YIi4JECBVbsZ34QHiezDzVBFLL1DCq3G4Ob732+HfetlW43enN7VQvMngDPw8B93
ptEPMSvm3jGAy/pEoMqzzCoZRLG6rphjj+tB7o2kCxGu5ikyKZKFO6QTMuSTTcdy
SH243FP6UgiTSKDQWH0pezDFtv/j6GYfhEyAqFbDms0vCwneuKdjnj5BZhkjudfg
6A4VimHyCbLR2r5828nGCY/wAK7o/5/zlIXmsCo4l1qZVv/HybkPXLozMtLqYhkb
3HfguMEuUwTOSwS23IUBPAxoVeAztXTxPFqsPPLmPiNYvy8arl7G/LwCXzoKB/WN
ACXE5Nwc4R5ZHaC2dWAsQzWS4Pd0y3yjlB8+DhQuOaU55fsUYRFuglYXbOJGlCOi
MjyLXFB7drgfbHMN7GbFDkeMiDsfsf/R8fB+zYF1EfuPzEjlqVJ8KeMAwScgo/rE
+HOob/yWlWGynLARlcB/O/s4fTWAwpIa3XjqjmJVb0VUhMS97Vwt74R6ByFreili
csl90JnWab1zWSuRvtY1P9PVPxGPZ3+c5Sb1kGV64RZm+rTUtwe0hH/hS1Kvdrhe
0oEn1tFre2n3DjuOlbazsvIADs7c22lRkycOUckIlUW7CfghgmJmYSYesvRz61Xz
sdQnYXjHH8XM4hlTwMPQ5gYhXrxabGRaktWkpSwQC7Otr5yhnFo8FRFjCoxvHusm
QVO7nI0PR6r0TjYjH+dk4HnFQYkcg6sk2NwLvDsLZCDt8eRvvkmlmSvDnC9qb8Kp
E2FWwcmuu9/s2J2Ui/c3a00/EqKw2554K9Uph9JrAy8zWB0lQh4zMM/7RHV/DR2J
p8NX8A5IfhwkGsdTRJ7kaXUY8DbuXBwXzkOvhcEFtluH/nVZFUkjsJXTevKH5hNf
ERUu5yzpH+Lz/9LICo+c8mF8tYQlqaJn/FXrNIVK05OgSt74FQ6qG3nVLelAil+7
efGGQfsX3uG8Tzvouj0TidxmbtBUNedjccdk+rZMYXMXZjYaAzK+Mxme0qWtCwiV
6bfVrLRyNx37LHv/AxgY6Hx1Xf45W46W9RP6dkFz6E3I/jM4F6k5f7Gfhhy7So+X
Nn51J/8QzGYhEjAiLkMt9ZjttBk707pWtSradE7NaZr9YsYmeANkuDbprgX3H1Mm
/ZvvBhebGjZbF//gkV4FAKIGYFVX4HrMm7snkCoci2QH8zyuJeDUFHKf0BXseq+Q
4baAhBHuTBTVvzt2PzkXQavweKoJ+C8Ng38Uf5C4cpQM40UKPlgmJXDUtWlH95K6
bqYEgUWRMN7B5MGaaXucGSk4r/moPWJBzQu+51bEpCoKVZlNRAFjv87WcMTEyLjO
1+4JDP5pccL4kwaVW6Hf4dDsYw9c2P3etyW11/V1lnyKh1qmHRlR1jYIaoS22Uk0
zwHwryBB58FaB1oIaslklQMbI4coOqE/X7DGTpmW+rSf16E5DZHyMmVIePS/P+5/
iM6xkhAlqgNesKodI5YedGFNYC1hspqGGcvOuK45Rt8gqgatW88fzgZOVn+oa977
50Z2FCUxXX59I9jvnu+wU1i2Tm5kc03/CwCJnlCtdczvFMsmNJXNhLscZxd+T9Sc
qLyFuFQtgFUFCSiPj/VhzoT3giRlyPzi+yPrLC2On3HbBp4MKjoODtgObcMrKNDn
BUMUSKeb6/zqxOkJZpyVGb50C2UwsOJBGGcod6L8v0nqOdHklyGj3LQG43+pNWKL
sMGw+yEvXt13IqXykrNKOscOREYtS9rlDNFO+woBDiDH7HvMhDxjvsxrRv66K/pQ
s73gvFUSjyZ/qUtigGGn9B+upkwnF4vbdfM1beXrny08uV6vX/4OCGKHEw2Eq38M
LS192P8wCtOXH0BQg9E3nYvWBf+E39b1dZtye13zXyTHKLEipsITN6cH+LawOu6B
PkicKN7z6TCghrlM5Nze4vbZ9jsEfTiokN3p3Wspc67Uiv6pvEupyrH3aa91IDeO
st+AggLNZKiEvjfWNCesH4X0Z87h1G6tiTLxtawAW3JGBLmA5g+1zVhWLmn9xQxc
ZSt0hwMudx9wQZqVxav/DTv4ZCyoPOIg8/CD4oyxZ7cLu6BFsgKn6R5B+bevAOlx
QxTkM2gB5SbJGNcqrAkgaNjT7d/PK4v6BwAI6KaEm2ce80O6CJEgOoO2X9L+fFRj
sdO6+VUAwyuwNc3/IE8DF6h+eCSpFuO26uFctC8lWIOcmg54mqrV+vV0m/Vys7sY
zJ8iDd+qvH1snoDcd7K0BH2WzpqtVPru4qtj0yJeV0uU9NDE6MrGlImHox4Xfy95
d8dS0chE1m8aFreDqpHPTlKVoqyrNPb56ChP5dMDwe8BVvwxi8q3FFeZckOt5nVK
KzYRDI61vwF0Dh/L0P+M5xhBnsEZvhv0OI6EGMcH67pDIFImPPJvfVPDNqpY6SkO
VPPBlEIim5Q/2bYzJ9/GlB+fl2gCGVZerxR581bg6155xirR9CYEOHNLPF07Lkv8
sGOSCuGwmzEmRQAwygsUVW82OG9MBCJzRPJ4BOhEY9r6FyMTl6rOYmg4iUZ/H1vh
3dY8EwrvgTXKY4Ud8K/Kjol5mJB98U6uG0DicpSp/jXAt77pid7wef8ph4HGZv9R
zTMLh1nf+1iAokQuoMuniVc17bVr6Ces+iDbjfKUytYw1hCYDxAaE5l7waqGneNi
kiHXcNYJWbNLpYFKFgOMQ6MTypZlfzSSuUxXFGrPG9l80D9DMkbwC/hUxA6GeM2S
e9c52YeUx2WhkgaGsjo/DSRvGwqdLUNBgPB4RJJWUb+aLLzkeqiQpQLoCy6/+bFB
+VBLUxPtAPqAG8nmWU5OJ/hLWBpyUdy+iki70l7dWhd2DNteg8D+g7UbQ7BSDiJH
Ntu9DFGGZHNBrBWkRR9O2CiYNG17iLnEKyYIYZbo7xeu7hKP97FjxPsCoS83g+OA
KLIuUhw2FZmyIumHbMczf6uN5NHAfik4edmB02HMRevW4J5DZncySoILViyAASG5
/mHxK8hdI+81shATTnWrfL7Kyf3hlu7ZrByJwaumoPc28e9Y3d4WfUmwBxmhX3aq
EAXYcKXToL3yf5+xMiZ1fH+tl4+I4hIHgQdNDqJC7d/t0w5im0Q38u1MZuJ4Ul5I
AzjwTNHB4ek4md2VD3wMGQSIuiB1xgtNlev+6Wq3vHEnR3rixbZjiZyoxrWlJRSX
D9HkbsKS/Ez+dXCjVioQfLtpXxH6UZuZZT8dtEMMTGyiWdlRA3SC7UE17cFT0Emj
0GCMKDZ1POsrB9+fM4nuIoQejUdLwfSnOQZ5cpE3vC7tfhyFgE8QzLQYnsh/CqzD
Z/SjApkIz0DCKZzjH6POO1OrZOVPwRrNw4y97ddZKezoLyNd/OVIDQCU420H9MZJ
vxN8dVj5jMRJRjfUCshwH8t5tqM+1fYCAb0j34v85D1GrVzD7TcryefbOSEsUYzc
5Rn2H3VYS6fFVNOkfJRZSfVtEruije/OcCgQNjrb5Mror93mxTog7pOYoPlhTOmg
Wy99r3OVAgMytBXdD1EWmch0YKIVbQAhZqrL+7wn4Kw3z0k9DVyzPW4rsM0I2kU/
srK7AmhwWVECvCSM1HKafYs4t2+ecO4o8dLlPWMu2Ok0VjIHTYk0cB7AdgVGlu/R
lQ+xKZ2DBM6DDVcHEZxlzYcVEyL0QGA2b5Ihvv8rkq3GOk+uHpQal0GdCI9P9XZq
BuuM3XtiAT+p0RyrlqkJZkhW8dJfBEk5K/YLrOBFXm/6lV5k/okgj4zclgZdtwz3
OdmBRBMVIiBvWp7Qz1wgca3iVPyHJKF0GM47aVWRRSwT6Ch5IAgiLRw952qxj2hd
N8/XoDr3FsxQEespWbQQ9JcvG9Iie37aeREZ3AyMYdH9huEzfnPJN+e7L3X9kS23
WIilknupvlPBRiNU/vWkNhrWFov7+tACDqSRHKd0Op8byjVN1sXi9egMYX1hdrdh
xWgsx2aj1aRA0OwcLUx1K1OVhwhkYJ95uwtvOL+6KLFJOQmq076+hZ0tDdgAT0/w
yoJEyGh1x1keJAGR5qCEjnkvOS2TDy4BhtoMUYJIwWNyfKWMM7czigf3OO7T5jo2
7Y0dOBYZAtAMAiUbBGLwC+zK0nrW1+NbGY8kUnVUdOFy/A9REEFnCWZUEWvkfomt
CBuvy7kX3saoAh2J3e98q+otXbh20lS8LVIGSYPpWzS4xICvnVGDf3LdnwYE2h1j
gGqTbbZvOMTVsZ5KGsf2Y2hR9LZN6U8WoaTUu7PcEDGaQrRUZPFVgb0iBShkEy3+
F11oFJ2GGK3wFvI26rDf+83bi02t1+k9BmW+Be1yOsO7HVWZzpRGCd1yV1KfxjBK
0LuSx6fTK3hMvxBmILaGlJd8+4jJw6W6duEoWO5UBfiYK8x6+uaezyfYverpDzjS
Y3f+vncFJMFnxngkQXYiGDo25VNqPjYFjayPBBXhBUHnTd9mfPNOUK5bzgexNlh8
VzvC8t2s4vg2CV8+NJR0fcru0Hz9MARCd/9hcyWVTWpu69iWPn3it5oLRgmQ1Pv9
DQ/UUuYJaCLjBxvG/7F/V/bftvv/nA94JPw//EAREO1OzFfjHLunqPxX5jtrqn6n
5fOMBOBkJ0mPq/leJjW3U64QfKTvYT2+8VL4mzEQRvV6kemEKzhN3haR8kddrjfu
Iivy9Jv9r8UiNQ1eMUFZFD/IiRqnAhiDIMIDEvb3Sqc+VSupHmDtT2VB8SG+csYg
sQjuAhmZwHxTp5OTRQ1t674u7+NDazS0xTp7JbT/lb7EXmnCPjlEON9nMabKQUPa
hap7ggoOha5J/JPDeep/wBes/xnMXecnGyVk3bJYnK4Ra6xtcZzyzyEFV6xILhky
5tFfRGl8umqN/p4eLiT21PyrunPAkamCQJOGnnqHz91I9OjQRMo6+USLyp7k2RTb
1nNglq6vaHTlvXSDxon2ETdFbRQ9WyIPRTQG4aQQBWSh0brgxBk5rzrSF2axmTKM
rY9iFZ2/yV1cvTJx4ZFQS6YjnNPf9y5ioXAZmkeKTSOb1RFatueKxrVwhAZ4PZ5J
JRmEwxsY1weYlJWXcdRznQAPVGDIOb1Hav7BnsxLY9v6XxtAk2CRfsrBSIrI6yHi
8PXSWbMkq8UT3H1Z0Bm3fMC4XYfahZLlXyxK+iGyxZ/4b4Y3AOdZreIC5BLSti05
pxWXL7kdmtsVW91webcg7xKTU0MM7CcWMgs1k2ajPZoZm38MXdHsa1BKFE+2yRr0
Fkq02w7YGNv79cSzMmHs0UyN05GSjTl02Yh1OrKrujLm+aULeeu8Lkscbwq1ApsK
u+p7DSye/FHh/wjCl93V5OJjY6XnXJgMcVQ4wA9z4TYj3lT0p6HKRT2T+YrAz2Ds
zbn6QUwhlT7RLcJZ7y5ZD240+yngQGcuKi+g7htzgWMbM1lTbfhYKNurBjFHAsFB
gJwAg+2CUa9CQnIin583rIldfyPiJS6BitVklDcAri7CPCds/evdPyCA0ZneSAAC
KRbVGegcxETYYLSxWRiUMlz+LtfltfuXWi80pKin7dEq1lO8HAxffCAhnPPhmGW4
pYEEOgXohPKU47w+JbsPR9H3C7fnFB9Y8hrLfpXqX3e6G8uw92pZE3Kp9kP+xevD
uZqZFEQEEJ4+H4yHNXijElZzJtKx9XnruGCZQ6MRjAcd2hnHWadWKqjQxsj80NoI
Rpj2WcGjPHLOHLNjwrCt0GlS5E3VNIOEkYhBfoujr1vMXH3VQggH27KmpHu4bf5o
rAOWXdY76BwFFkrSVaVeNJ7l19T8Ok9/beYGDnfkY/A177wVj+SpQ9Ix8cNQQkmz
bO+dbZ9t9mLPIu+qlaF52WuWiuGufo7pvsliLd60usGhNqmPj2u6snqreHIuPIpD
rc3AuOkUKt0auV5kzvaAGHTMh5B+S/xUVRn9wlDl/gfJSglKkbdIrBELc8uKjejx
KX3Q+EvUfRVtAbVjMy0Ptxa/zDO9OW1jRA3Xs8NIoq9wj5IAhZQd6mZkHcoAZd21
UVZH6FjTbkbf9vu67uQRVHqcVESWrSBSHVV3NybTz4R//qG6CRdjgQogzVU4FXbs
tw5kYp3mOuKx8EEsKi/LscSaPOBZLY3CSHtz+T8Ik8hBgZCSerxtCTKwDArwIQ+0
VPrIKdnLBpB1Bqit/CLBNVasecwO+6KVBIHjM1R/liS29PqvOpHCzibtlislCJ8F
rwJ77Iq71Jjx1Crbxyf49HxBxhCS44YsOPib4+MOjdpYEALs9NT9QfKVvE2YHZTQ
YpuSDvWOx6Hbyyn7ORiNwqzxXecJWIpOVs7SDKRDawvEQ/5Xt4hCqLBkIK0KXw3H
/tdOzi1uzmFJYcnn1GkFTJ1sBQF/fGPNnMr7pT39gICUZks9joFH0aVmoYoxPP0P
bQAA21m/T1BDvenKiXlBlMPhAymHl4ocYV0G804AbFvBAoxUUoXc3wH/pQaDq71F
u+wtj1WzClE7RXlI8TfQFOGEQGgSWeGJF/t7RxEzBf3RAnHiretg1/oeMFnCQM8a
f4WBV6MTYA1CeuKXgvzwFcxs8mfJAU4scJeHvaI0qTFTAzIl4700aFUwCc8BhOEc
4KcNR5iwxOVm9c4wMtLcy3eza8YKCT3FAa1U1i2gN2t8W7YPNIFqwDb/QKw/+8Rm
FPUIJkNFBUqpRcTziHl8b0/GeXT0dOYAbmvIyZ9yBjOnll9aIAKpivwdhaIquAQV
DQkANicncwSNuAa9FCZCxvesASPDb5wmNlvmklWrNpt0li/Ntg3Qr2JaEEqSXC13
q6CbmCRwuJbFGDYzho7Bjs1hJXOWmfkhOxjSEuRHnX303GtEte2/bjS4cJKrsudh
xJxDvs14C+NDc8d0/NHJVFNq9/yHTcuLdh+34oUXaxhZPP5pt5WxTGvd+9/IjPUr
ENj9aVWy/pAJwZ8yEUHdrWs3u52GpPjTTi6oqv/lJtkCxNFz+XlEpTo9zdk6ZZjI
yUymg3E1iG2z6/Eu3yUZaQkDjLFevIbb+u1nZYOfxidBWF+QRP7T5uTFYmZkOGlR
mYq90aT7s5UCUgf3rtg9epApK2XtEfWTIdl5uVxDl5jnkqtI4vT5iDZg1OXnKBVk
66lDsO8SY7jTviEBv3ZRGhDDTbkmT5uwteyCBkjJ3x81yUdizEVETDzpMRsjc8y+
tRtfkNzaJgYMW/rsMIvjb2xGB2whmReErFmgD9AB/qrGkWA9L9NIgYf4HtSiGtyJ
LucTn0uSl/KWJE1AeXAGmLW19s6zQGc1H/aFMJhQFwaO6nIrsvLenXs2v1tcxQZX
GaT7WrxMkKDnwZGXifywe4V+Abdn0JGxQTWgqU7gdutb3apQnxsZG9ufLfAwslMr
NT+jTZ3mEyR2CNB+sJ+5V0Bd96tOfgf7BmSM09+k4qM26tccj+02YobvK5f1IR8d
+usBrNLiKvoiLoQQjcS/fsIyJc5iGS/yCEgMDkzvF8r7t7bQFcwW4QNRQlIYWg7k
2ml6ztf6Tg8pFvSJfUMwKeSDwL/l7F4wHe/Dniy2TbR9Mham1jP/3X6pq7zgH0cn
8xfZ3w18khrrCirP9NsqiVzGrmRkgOXL5dihzM78vnwkOwXyY22Z/sObu1zttkR4
lc/gFPjuZe8L12hUBZnTouRJBVDDzqTx4QSbMmn2dvXHa0C9yq8FLn2y7zyBIGIv
paRxaM52Z0+rZbORqEh4oVBxv7NPXuDpOIMuZ9+K/p8SXslqFNKzNrOiFtm6WWQ+
B3T3Jow3SWTGGeG6Z7DZMUCojJ4WB5H01ua3VX5w+xbfOD7zDdzDg7rdjNmGNk6U
glUmHHqvuWnCyANI3gUnBo83IW3OnGgWcuE625d17m54k3ssjZTQrqPTP2v5i+7a
bQAYZeWUsrSeyUwSgyzuCxBBZ7RYB3C0Pb43GPagXD7H1JiMYrwcDbUC7Ydc++Yn
sUVDYgL/gMj4J6NOhD5Oq1ozyCRz4LAZ0xXCiHzOoOT3T0bVU7hKEu5MNG+XGitp
ZeyNomkxeJqoU0dhiTldRran9IW8A0Fl5Dz7y+BKbVohdDINVVmhy9T6/B4J7ZtB
xPXHwyREiCu3JpwGcX++ASvN2xhCGU2liBdPB4B8cLRWq365EDybmltdhFtF3wHJ
r+45lEBO+Bkjv8/fGVAuICT++GqQKBBKgILsJP8xvV7ARxqoZG+xdpdoXNJN6aWb
y//Ez39g7ZKEv4RaBjL3pGAZi+85f4G1ZvKLqhEb1cS4VyI4L8s/O4iKzcC1KoZ5
uOiR9KG737fpLk6o1E9jOfshoqQL2xvj1mJRDzxt8LJfEv5vfUCIa51OYrtJWeSB
YXh9MWoXVCpH7TIfyuXx1+iH2ak0pAiIL06UaDpXChEWJwwY0nJ9ivV8O/6aEQCz
G0/01UoXwHFekopRhCnOCvwpn9gzzASWfxU95a+8Svo4J0WoMUDlifYrxCm5mdcf
qJX163UM0CSij5+WGc1FTD/SvfNO3QhBg0jMMsYalKjB7VERruv7/8XGpsNY8awV
dzThRr308/ss/p65e/OuYytRkA4KMwqvNJjMo8LsZqgiTAmtvdaBQRAEqYI4bJZ5
gP9AiviAG/sOCqYca1bZ5Jf4o9bxMuI3ky+8E+48+TASS0JOfFScvD1aOWjQUNu+
6cCOVjUMNN763F1vZfymiO8TPjcupr2kf/xyqayBd4jkAwecrhAsnuTjA52rcwfN
2mfJ4C9979fGQRkitECb0SGRaHviHSz/DlAKdnbH1e1qvbMsmjJP1UoYRSd8WqdW
EdWvYvf6+PFvbqe+EIonfLSa7JmEAucOxTfZ6Q54JnPDtZ4npBu0lunVMSXB5kID
6mKx3z86BMLcRhQ6ke+hQKDm5GZu6QwkU19lh1EGDyyjU5znkUgWs4mqYnzlbC7N
EU2jJNzVMWtBI8AgDjuCAoO0m90MnAEcir7r0/rpr6AhfSL69CkGUqDCVnVQ6iT+
5MZLMGRIbSKSgFmIFK8cIjV8NME0VOwZzf1bkEp1z4CLfTzbnju+LBB7JIKwXL3B
e0QQbNFPs1bTFsCLDQQ1WMOcLxD9GbiJS2pTUtClOM0/Oa9FIjLaJFD+/0LVqNnz
o71XB8HygEWLLY4roPX8GAWBuI55LTbg51ZRF8EcV7ilrNnmX2ldDqQkQSsHQ6l4
08owCl6xyIi6AtR49hvk7FvnLeGjzEovFcdVz/HMF27+nIIaXlGgY0R582uAPmj+
5hnpAY5MGAs8cTzMuEik06+S/9T7lNIU8T1ZKImpGipU6Wcwc7ahaLUOuEwFpB++
xOhohQ3O4CdUVzWEUu7NGWzfWcZmXJeXa2L5u8IdZCyM15oFmMcdvqdFTlwcpIfA
npHEHr1EzBnleAoCZe1VHcBnq3uD270rqDnssJM1bPDLYizMBhHQ4C9FoWK2jKP/
3X7g0H3ImSv56plNJsWSsNGuZvS9jj2NBxx0JlBLjewfxyD2jsuVFiT0Y2aV5Xks
e4wpRVMCvOW47IwlcMr0yivsS5KOHyMjeZHg+Re6b3xeVZx4XfuUSazz98NsGEdo
F1ipOBaLpMsaij25Up3X9P0BLHW53czdz2tqOwIjK9LWwr4wSXrb4+J1yufEu05n
sYVBkZzo5Azv5Cjdaq6U7xc47f7iszaVYkDwXxR0zM/PnMYzQI+CHHv6Jr9pmkXK
QEeK2uXjDaWGJP5wPvI70j16Ruq/S+pf2CSyz/TkeZnCkRDfarwIMRKnLPwT5aDT
H2f539Ekd2LtdQGaSWYodTYQXEa5m+HgIdB3vzVmmrpMtFysy0HmaRQo1WNHLIqA
gL1x+QGzgMuYcb1F2I1V79FrnHjzOU5op8Q04Sd1GgkJLIvlLDNVo8Og1fvBGFnY
XNcMKP2zB7p/nuP5/N6e86IV+y2KeVn4nxu1B8HLLa+18debZWAWsGtCHRz0Kwyt
M0D7Zq7KpKTUw2wVEMwyahdFmwdMV4PFUQ21U6A+cDIajJXHPDoZK+p3vNi+f1sd
4GSuX3SywSkH4M2hwVKj0jWtoeLpvuRI1fgXQoVsQaYvVEwTVzi2mAoff4t5QFIf
hgHFkl9/zraISFl+PseRjzQxv9jOVXikIC+ecTzr+NaiTeE9DZgH4ztGoebvH6j+
pPXyIfC5i14kD9YSvNjFJ91AAFcqSK6Y72n5UnJqpd4DNvr16uaHoOxCPN8C3RnU
JDmLOchxeJkTkmOMA+tFNeQnCYuvkWzGfkzIu4T/kVfO6V5fpQKQO3CE/IpSw1RY
X4gYNfcpB34/yancOdnDugfPHMAj7YadFxtNK6Md1kMn9yDvXmKE07XgECDZHW+q
Uo4i9elX0TRdkjGWtcddb+5CuSofZlb6ZLzdElDu3PUwyn3y5Rh/2gsd8EfZdTaR
3qolqzTOgWiZtRte8rUdRibHsVS3CGIirPzeibu4kYKq/Bu95fv8lJeIzCIsPdJx
Ks7ycTOqEgMB5lchLZ2av4AJIqN0Kr2UNd2FCBi/tF48wDqAPuXPhX75dK7JjdY2
D72raXJZ+RhZbEUWeJTMGtESRrGRt5hr8Z1T1/6sPx0TEz9pz5tlTUvweY2yeA3/
s0rcydsW7q8Fu7zdKuL/WZNdLufA3G3B0mFKDLNkIZD57LLA7+EKsZH+p4TtczO6
v/2lywoMv5cggTXbnoqBFAVz6Bh8URHbhWN/01s+E3pIBhGWPcEiW2t5zYcOqbK7
+03ehe8CpQOckjztjtA5DL9EBzLx6n5zyvCkGE4efVM5q2ShUQqsT5SmDFu4TnGO
st1AUvNjKILahMVrbfx6PhwkA2dOph3LUOJYAzgkigwCX+Wayv5fh0RP86ryR0Xt
kVEE900vyE8Qy0LjaWoz8c2wEtajwIIaezWMY5d0Q+Dvt87i5uarsRwAlCpuPP/A
yKotgcTiiTjLuqgAM+Hgeszs/PLuIzvfbW8g1/bnuNXk0SFQtmZfK9aDO1gV1BgY
2R28i0xFEvPIaG6iakEnnliCPjNfXz4mpLAeX9Uz6MDFuntOmpY0/Kjp0lgRMhc5
HElD+YZlHTtSnn1f2cInNoi+WaWwXptNjl+LdyHKqY4TMeuA2nqT1aTolrJ2fd3A
v5LYwwCbcq6aiYXdJnSofY5pT5xTxqDuJ7kXUHbPSJkCWkQr0nn1ukqcapnuvf4H
mQxupNF4b3VSSl4+RynqthBy2+ZQBP1uV+XXp4PnLADNMkiSTrKS8povIk0Bj3sn
L6Ce7Toywa9C2WhiPd8SlZ0Kwx50qq6lsmQ1bAMO5th5VbXhCr1M8ZPm3BIyMBHM
Yht9ykNrirNykKdCD4EKe7ivzijIU/jQo2dBRVG1JtKyA6ytkpSZglXRYgvrVxlS
x6lBm0lGnnyYZbQQX8+SfDmpCZMkgGVeWsfQyO71eLoEcKDtYb6jrNQ+yvLySU3H
xF7dIgAM2keZehBMVSKoRzBtIAyXPki94jUldb5RbsyAqlEUT0TJLwUPJ/+4Yyen
7tqHpy2nJHspm+L9YcHUtR2j06A5s8WnYzBwn0/CWnnwNnaAM7U9jYYAQeuN/v7g
sv9rzwV2yrVhLUanZ/F9+Ol9sgqn/D0GuLx2MBeSW5KkLEwLRgo4f1h7O1iDjEfH
2qOieOA925p4eFi9G42ln0HZHPQke39FH0+93ZBXH/ldvTrqzhxr1x9cXdZmpkX7
2wtlGuLwwr/MwWgV1KkL6uNkwboShFlqgl9lnQO6sRp0Hz9VSDY5k6nlktjnbMD1
wuQRgnQu5X4hjHibUkfvIJNgVw8w3nSNTypHrZVpan+IfTk6Ivpthr1zNGD8H2F9
Z6FUyTFsHGaqcKl5GR1av9iJQVA1IAZrkE5l2NMTCgFpZQUU1qsWLOGkXv2hIF9k
EloLFOT73fAFnMfwxa47/rCAvN+EDqZaEM5eHAo2iff/vklBhcE55WqD76C4ZLnX
T/6uW2yvtPzSvVvW4q0IrFRj3cqDAteuUyVckwA0AA5tXgCMpkLBg4rDghH0ZoOF
cbmQwYoXoerh3rNkijMEPaKdOtcCBZ1uksS2ypRGCzpdD3CSU6zkZzhMPfcHPwru
3Jk9qV0biieVHNt1sWT/VekY/Xh4HOk178J4nInsltHet5aEOXLON6WpUpeRAAXv
MEdmG3F/9rn5AYSnsrWUVJjlT/7qnQvOCJXwMQ0LDQDMB9I3FjdSc2qM7JJO/HYB
d3AyDTwS8HJ+UzgwZ0eEqiq9rW7d7rLbhtHjlrBZldKCry+ELt30b2ClBSoaGAcU
b2K9d8efAWHKtS6U46zhYIiiI1ExquJEne+jPUjjTCk8MR/Ex/2LKc+O2DwBFmkv
s6b+zzff4Dzc015Z5k6xjaJr9h/P071u6Kl05CZDEPWUotzKuWRTLPf8txf+5FrP
z5D4Rx14Yk8bSQo39L+xqiEiRFhlOKYH/8xicdsdjif0uvWDaZCYXlVk0Rfh9BdY
Z9IZI+S6zhjomOoFVMR0IWAc/rT4hGSGA68Uis2t9OdQuP2v0/Ww0VzB/Qs4Ij3u
v8TsaxbHIL10GjKe8QhKt2Dw4ZWh34ghqrHBCURCOuB5g1qrzz+auRh+RFQf400R
MBoTdW3n6iTRJSPfeNd4g2yJdZF3dqjdAHv3WEOpCbcwUU2HIvn8TGkepBHq7Q1p
DmMH6HUVzGIhymPJs9xkOXj5L9+xO4YrQpOe9cwswt+evZ9TnDE24QYt43YP3q9n
JueOKe1YK0Qmkib1yBvFJfj/a3SdUdCgl1r7LPpPbzUE27Hhk0oMe/o8Z3hjLlk7
lW+1KDUAXvNKRQjGGt9oxrTQvv4QyyyM35lcLsWN6rcB5OeOZmCUV86zofLl78Pu
QtQNp9Wkx/0eyMkP21yYi2eBEwKD9zpSiPXrmMG6nJM5Cr2SCdg/xMFeyHQuSb+e
ysp+rAnINMuVJalIc5GrI9S6fYBOKaYAE9BliVUMusWakN7tQL5ts87o9zSmGwHw
F2j41tnA66v/VopRL8HcgIrx2hmVRtzFxlbP+nD6WXQ+j8QeGE64VuOkWIdlRXgw
nWGHbw3Xs5QWFQxCyE19rIHESv/Lp1Yolp7r4PtGPaGOi9XRgCfHArv0sLwiK+pU
Z1LSX0UejuRwp8BsWsWNzMBuBLWYYkzwR9X8rzkndlPIuijEVgDWvQi36U6GTgbM
7swJuaFhwbz3LCy4t1sfzHi/qRfrYS06WKYBGEENBSdgTJNqqb6Ml/tMwrd4hwSd
sjFIEv2ezcx/Lx7hv2/UguIIjnWCo59sRkNXPG1MNB12slRQD/HNplg1TjgjJ9Cu
BFqBA/mAKYU8fMDbLEmi6cHmGIcvd01MlNHH7XjMYy0vKoPWglroWXOw4lujk5X5
RPPrJNhDWuI4QxVjWdQeEgBWpIv8dusox6YqgcwmXXnopxImpaQW3+qCVdNMmrR+
a1pVhPDSSWrqTnh/HYjnLHAjI+7bM0bXg04cFMgtVHeqgAnTPXiS8SITIOrpdr48
rXGbffiAdGpPBz3/XtDt3WLckuLNblnmjYTyeUbEO1PvN9d+EKXrjTSj9QD+6ctZ
8I1pXtLdpZLmjcEh7KTt9gIkBluwX1asfzG0HDrCstuebOtuEC5rXvfvFOiy37n+
DqHx9Mmoe8V94Ei0g9n13Xwj6+rlaVMxiJzwegcspQ7WjU5bvaa2T/AxUGt3n7/9
L6NVUxtlxyDFWUFqMd2wU1PLbR0U1DuNJWrNcwJqQQe16Jyxyd+2gEmIa5jebBjL
YyZV2a7hOsbLIFhbCVWX5t+0Y/0IkSw4BCVE9/oR1CGZ2uDJd1Gopgi37mDyIPcg
jCSKShIlaWxK0vGNzGg2YBstEujIH4pahYqe2wHR9oRJLHIOojWTDRHESCK7+S2c
IAq8B5rQC8Ei02T5JTIWNBlwBbIybf5G7DUjCcJzaV9N6IWTZV+sdqfK4PLnJup8
Ch4HXygUvjBLh7aL8pHkFyrI07OANZICkvVvtiB6z6IyhnwGaA6DTiFWawggEyC9
bmH+HOTOAIvltDBxcqcRdH5x/aoPWeC5pxNJgbXWbiRUN7lhE+fUhkf/G4bfvh1s
btv7NaiOhyShgg3wgl+xfuvKigNva4ZKfPJFE2N4SRbxOLxR3wDL7DF13KtMnSN7
uRqgkTN1em90cueoNFeK7cYxvGePC3u471WSI6je0kkb4B4Zc2ecoNjeRQvAGCgn
IwCwcvcS0IVwtN2HII1gtQ1S7dnjZvyoVxDqQrmgZYCjRBpIGe8iKZBYuyB60J7n
G3NE4Fc06porKqRRhZYh+zzqboySK3XYzPBlEUureyM8ZtN/7MQCM3Qu85vsO8mk
WSEGCN2v4W0mAzsubvy7z1GmsyyQVjzaFO7qyrsk3ZWXo0FQsPyra2IueoZRB80Q
XOc26YkMVA6WxkU4DVEoPqyjHmg/UnEw/+712zJ6L02o9byFIg2zSamun8xHrl4I
pYC4NUkBx69mO3t9QFLn/390j+iK9TiOG7A4RDO6Kjc7dIMdEXkvBWzhFXE5uddj
2iBZEaJXGkFxI0CAVrUmdW8wh2w3uZtrAm80XcXve+RUgIDZPF+dc3I4Ws5JSq/j
YCKoWbASEaLZUVKrk39vz8CpZIoO3RhXN2zJamNg6my41oiO41wqYCJOo06z9tcB
/4RgYCNWYPb3J1LgGQDrdXVTQ5fMWfnVy2lSNnpvEZgO3V3NOKvx6Q6+Rpc2eLfy
kkw0e8PJ43Tl6FCtRa9oDJYqnWNDQ0zup0vrvkmQ3PbxbO0Kl7JNsBHLVrXlh8vO
QoiYM64dlU3D8PxKv3nsGqjif9KuyaMFIvuqSRJSdoozorDeMX+N4SoSdq51MdCC
31M3nnLAgmYgacWBXhpsd+Bg4ZzA+VybjKiCh/D5LQDgA6NuvKE4DR6n/RDBAmR+
gmTgmP967Ys7DWkCHSeEDrwEQYjQ69RkSQRqaf6gr/iW6pt+YXD9o6kIy2bKBtpT
95CgktvSwpJibFo9eU9jn9kaCwS9WbsMnck6Vi3LwWb56NvLe0wsKpsRC5oYxqfu
JvZYXvv9qBQjyHlZ22bh72sHKkT9XcoUONzZfmuMyB7cjFlQvmr9daIPGGVOnafx
Ym7vmO9O8PS3zWwFW67n8qCokM6RdeejUYXtA9p34OFOnyAc3q6ChKQGnyxSuVqR
ncgpBti2murbZxJE8soLQZCmLzrz0vlocxSlkWPPlcREWBBC17lWAKFtHvcrG5Yd
URGilTr3Xyq6Rv2G8mLxgB5A4gx2sdYihDCVCorCLLRJZ1zGM3izB+Yleizvcu7X
+NEv+nQkISvg3c7TnbRDOGSs6sBlpt7CZAn11ugbsXxvm+DLgp7OYc92oUM7crFe
Xi+Zqru/P57MQg+s+AXcjZPLOvB0DOYxtuuhtkpE2fEzZyU8OK7Al6dT0GIg8iyu
K67fl6i4pasOCd+Zz/fkRo4+w+NLn5NVUVwiY6d9Lhpb25wyCl/07dYfiBsX4KFO
CkeHeQSdIcA6h/NQvFtPrWJD9rclKqHY5Q7o5rzVlaxfXJztKyJUHrLdkOlvRO+A
CjKRvRYaVzSy8KtBx+0Nk5SAcvpJRpc4HaO/njqxHAizcaOas8tD7AZvoVBBwFoR
TzhFT0fFq7VSQvIOCCZtTKqdflnzyKZyahfkNIEXzoezu8P8QS0tbhEfGBkJ3Ouo
qU0nLHM9v46lvWoWJISMvS8PoDfws17F0DwquqDb5PpLor78T0r0TDqdOf2/27Be
WzEz+ZWat5RPd4knmj+EpOhjkyz9L/9edPQw6cKU7JQf1Z1sT57uMG7/wAbABqFI
OvIqHmalppa+ouVQ5bsVvewofcqhVE0faqdH0O9QgEkyrAXnEYNIjBrEAfLyO10A
1jJB35r23Pi0My1KuCrR9MhACy9lr73dI6zQ63XPl681EZoPoZRjyMaPG6TjSNFK
ATptnSwMNnENx4Kv7b2nCcMZcqHORWBqF4faQGdIvmoQ9O311oRGlt53DJ9d6mgS
s/o2hDVJQQcP5E5ZsShQqEFS9Q/fDzMx4BcYdn/r70LSwE/tu3ZtscegAgpTCN3J
RKc1obTDpPUVwnvU+8mDdMf3kyh68WzN9DhpmQBz7Ul6HOQsRd/iDzptTDvifHOw
1RsbKcwqcJBsDaFFE+cVn9DYtVpxaGtoG6OxM/U3DGMlH0MN3m0ZYfQtXbmxj+m3
O/dKO869K0TvN01s55zGKWteouw+//UR4h4xPgSz1p0Z01iHi79agmgVfDU0J5ZL
nlxOc95b/cc0CGZapD3RQl16Ula3QZRseNcTg3bNFS2IZ466pBKTI6PPoAXOBr5R
O/ZUByyFxR8Lf6oBbVUdFgOpst8ppASUuXzXEWlghASJc60XDTkSfwRtCnk3mLJe
8XHQ+Rek9EQPQ47fe4I52nc9uwwICvjrNQAyc7nTIvN3Mmby4zmn1PxmlUdu5ay0
/K2Qt8i1U4NSmP/DRfvKAD+PKNSMARlvbxBCBi7rQbXNuDGFUWIdwL69mSl7bHqG
cl+qUP45aqUHmL/EBzljvVNQE9RVoDjwtbrIhMpAC4MTxMMQtUmm8QKNJEA1rney
9EJoJW7PSuJ0FwTpopkt34l6Ta4M+9PQH3jEcz9vZc703x7K/cYRAWo4TUj9hBvu
sBAGDG5KwUobCUQUNeS7YqxMH/6AIjz4mgS10306KzGCLynAYr0Gq3YvWHZ+PFar
+705DEHreI9RTLeElor1NR+LnXZuE8DJXcDSq9al2K9ZvEwQHjNVFdpfxQCdbxrc
RXnRHnaCrIsTERi6+NYGUDa21SiACVzCVLJ2laEfGP/lqZ0tS/PWU5SIlptEUZA7
eM9BEwEo6yS+3SaSxckUSJ/7hrD/nZGjZ/BcO8+xJ8rCF9LpY9aJxONEnilttvnY
Zq1Njb42qmAido/RGF8VjOYp4j0jqIZ2uG2rGdweHBfmfbaC77eRejMvDkENHmvF
4YNZpS5QzNqfv4zmDAAZVZICLTzpqMFB0narW3QqKxkeZCcSkd/0xczZ+z7uaCZH
di/qRPAHqkbdpqRNLOUk+1d/JJG1GSWsCarqY2ecI07Jw0oN1VLFzY+2tI6Q1ix5
h5V8W5cuXTksGEOIgR40wMnOVaixtdvT0FAsre38f2tB/z7SY4ma5MGixbvBP0EA
vbmU5Z8vW6YcnNgoh5rSOuwDaC+Nxbssc7qvLQndf5nM1aim043DbFT53dkuNruz
p8KJ7XS7XelT9fEnAau73oldD+YSsvv4OJ97tsXIfIme4zZlnG/7ubbWAcm270By
iMg6fjLA2Mw2ZOKb/IRo+YNfIa9HkEIyqZSEiRREFNv02lBoKNtq3R4kNfhpBjBV
osmAnFYc2QeCKoJ7UH5iAo6j2FGYP7CbyMXYJ7clXsA2oJvAO6lLF+t8nkPp+8iS
Q0VgHU94iaiWakumGpc7VADZFFjKl/sTBVSBOkxplfW25FLhxEfOgkLX3LQg3pAn
TN9k3OaspMfllkMIPToXZlRqGTa0s8XI5XSaITOV//6L8EFM146S6XlC5IGMlEtO
m9OtY63PMa4hliVzyFS5CKthLETFiaupPeQ0xeITNIeeG7uZ6f3/JgIWe92u3Jk/
AFbXRf4gH03TSFRN2TAgo0k2pM2GvErFp0WfUdV0GlKDl6yECCW5AVpRPxCIWmTT
aUXIf3hBPkJDhgWkR9xzwi3Wj5wjrk2Y6R7uT7BhTgoc/YoFGrjR+GqNF2a2ccpG
Huwsjmjgsy6IX9MhEQd68RwGSQB0cXg9jkkcv9baXxDdmhqMlSJeJ3WWBS803pJP
At1so/jnoGq73B9zmDhKquwk0uidi1ZvMBBxZtH1+/lsqeEBsPNsLYse7RuH2+fm
0hWEx1rwf7GrV5XL6IiVe02bIUu3uubnclrkejkJecVOtkojhvFS84khUmJzs6J4
vCXPMyNlDKiBW9eNR0eXSlwWz7Odu9eirOJRRIMdrW5VAZ5UjlYhpSvG3XIGnwr2
FhiDoMcEtC3CaLCrlzq1kGbVbtg5MZu6V4JQ7KHjtk+/YWZ50js7VdF46Ccqz4zb
j6I4bJK/86cRRHB+3Cuee4895H6LH7Mhr/yD4j9M+IVTbNz/Qk2lpi7csBtiHovm
BxSp7T8AtdHsVkUxqcQRMcIVqZEcN9XQejxVZvjO5BcUfJB2ta3xhWirrN1klHx7
qNWIjxzJ+tQpFrfHGUtuJI6gEfgdm0PU6w7srx7rS11IJIDlOsBA8htzdqCyxI9A
XTrFAhhIAY85pOdIWeHAPx/hGarrLy3xe107d3QVXY5BCflzYtQPE49s+rY+Bfgv
0bU0fvdvAqzVj2cUhCLsWk2ZiSYh+3K8tIPRVkjH9S9ntqBS2MWf2JFEMbWJWe7i
MGbsZoJoAzuACvoWrjrNyPfFABNinn84tHmZJoqRTg5/s91Lk8DguR2i4XdSWrRh
+SQd+15DLFD3uYsB5eUPK8Z4ZCAalyfm1Yzpuo36LFedeQS9RT7dSyjMbGY7xRsy
k7gZjcjbAgZ0VEblOUEHTc//Mb5LCAD9ltB2ksRHHvVTtNADQHNcyArRQ2jJz4+0
1zp6ZnKmN1dJ/wTPZTBS1A+OJsjOQox6czpNLS79UJCvM2MaHftd1swZhtGuU5A/
bnnBljnY1WlO58kLhXVrn3P7UhPssjozwnTNRToCYmOCczrzANH7YeM4YmLOCXsL
EBTrNRyeZsKTUG9p9hkdY1Tan9xihTGCzAQlwMooU3N7kSFEj8B6sLsmAc6rzUHh
LJvSklmKcxWWusEn6EjcoRx/ZPx524nYYygqw8ayweatOERQpEiqUbEzxeQJ2Yac
x1zWicfVoVexc/j3NMRUD40L+DjtYicDjvKVhRkXZ5x1V/k3vU0u66LqKO8bcxmj
S43E5hq/Kt9+nUB0sZAfSDe9mD9OrxbcBGG8ZUzwPbea6aY19L7I2Yoye+E5bYsx
m2t8TvCAH+MLn0gGrocS3KU1Pv0nsBIHxRDtdWkrwk7NEiVIn0vneC85wEaPZODg
V2dap7ubf3dAGy8H1QrdUWUpOSLrKuib4G8bAFSZvLz96W27oNRgeYPN7h40ZJIc
OXjbWWcmT8xMiMawCQjcFUIhrhaI6Tu0hKGG/W71SUVmhJoJn5tr6YTEkz4H0dTw
wHCAa6FeInXI851CSydo3YcAZUlW3MyqxNTP3Mbf/0hhwKKjzobbgkybJBXFbM5k
lPNwvGFpCebhfFMOc51GKmbpCkx1xgzU40k0Rw6SqY0somWZSWEVr4PnMCsYkeKt
Kc0VREL2iOR5uMtX9cL5uA1u6fyH1ns0nsU4jy7jAGeyKd78+wtaCSfxJ3gBq21F
pE1vEkf4zvKcm48tvUD1L5cdxbtE9s2/UVPA+i/pJ4j1vY5htwV7kSKKmx0kudOu
Wtz0sLAtzVOYQnWHguVBnPIWTXeZrNsaHLZXCi07ZjRtb30spk7oy9qNRqg882Oi
tw3WntrqDUjxAPcq0kf4RW7g686df/N/e9u8l0r6lTuE+m+oxvlkRYqXN/T67kbQ
yzcS68XDdEjGBcCVojPIpj32Z3VCTfgjd0v8gFmG0HM3XuZxvOWr22lUCYV9lVj7
EGvp6gcw7QtOmqcNBRdhrp1kFxtvtC08+RZRV0002TdzHgAjM+tdxGNC7ceZO3yT
jZ77A3kv7cI70s55Y9kE+78GuHY8PAV30EDpKj6GTy9u04qwf8zsTjE0L8nCf3JE
Yabv1tLognJm7OqSD9lYzBWzd2LqI20iWS7qrX7D9cVM1lX5+0V3w5e6d9bCBbaB
OOpweTW+2I3tje3LL62bNyxI+uzsnE65CW5X7O4sZlu8VpIBBgz/MZen/q44qZay
v3NMNJzRk5eX8tQw3Lo4RgPa2RGWshtybuPJY9zT6e8FVY3tkYDxJwVNfRxc7sL9
ESgUPhWc3LlPzOeyVrqWm9VflJrjFGdYQ4Jm8X7xdxqyDv1O1uXnS1ZaSVsS6gf3
AwtJdw00+c+CwaO6lbJjD99plfxvywek58gZR/14cDmI58pBqnJ4DmP21LHXS1ib
GRAY8b7+fSc+iQ1EY8gNuK6+QHH5UlsO0Sl0LypvOMyAGd1WGy5X9dOTLQsJywSb
viO9hpOM9L2CA9smjK4ByByUeh5EGVxduNiWoEyY2RU+0b6aos7tajkXJBgyl/jd
HDxTPikPrepnKbQe2jd0jOZQRbX76zVW0zFyyhIAFIVo8cqRRgPW6ZUccYupzeVT
VGVjcJfBHSWsgm11PE3NQqBzcHqJwmykNvd2J7l83iL49pCQ4gd2l8ekRA5k1AoP
eyp+REoJqPidSlwXrBMKA3R252hllbY7Cv6OanqrpBPZpcl+WcWHw2NV5kSAqZbY
rabtR5155Y6N7Nh+Rj22NIUlq5qBYSgaPG7u49RC73U64laHYUgLorKJ8NlJIHJs
B1ZA+KXy8HkLpDCUIF/8z5ceLehB7+hVZ/3VnVzdMOlry1hBq28dEduR/TSbKks+
2ICmJgRLwDhxopHyB500Xi9BOfM6cxSUXr7sTbZUQwoMlWYpQP4+53VnMMQhmg2m
aWifG3UwtF9RyYXHYwb71rWW0eWrg2XEq5BNNgOGMoUKzZytpbiVK3jTmJEFIup5
BpL1rcZpXEseowDNetp+YE4cglgq6XKhGtrJOtbeiaC2kTEWxVMthJuW/l93rK/C
bdOhgCJHnAM/yDp4YuH0XG1U8VpwnwbDGSojW5CWJGJbsZ6omTBiRrVlHRxLXR6E
LA02OyL2QAXM2qGDlEdIMCDMfHo41fAtswOfmHaRYsHezy22/6f5LmEkumIw0o8g
ckscRBhem5Fm+60Ku6aKVPesjVqSeEQe6xAm+9V6CiHUjM0ugOWmZryufg4Jlu2I
3U1ltnDdMq4m0xVCRHjFOX8SHpQ9jyQYFn8BfYX7BQJ6iFM4ohItKRbjGfc0LvmU
+n3fc+6GY8VOtSMH9sjCmKnWZ3571xbeOOndR4MpyZBHP3smr0rRL7KFEQtBM42U
woiSm8ikf33X+PNj8v1j9ifkyLAcQD0k8YnY7cFExeufmUhfMn7YJQbmoOvgIx60
VQnjkFwGnZJ9U7IkS8WHVUe9iQw5JSbS9I82gdLe+ROYzNt7tkhxCX9lrt0L0Qk9
CWN0h8g1eF+NUs8o39AhD9gI0tFOZt1d62zhlzjTgVM/Yqs3VzO6V85PqxFu8FMt
glDACpWyt7OKHiJ+Zq9gH824YPTnb2qbysk7N/YvHRylTJzP690gQaCkvFJgvz9O
FGO7drIkEF88QYjK4B2Cr8qfiS+RqmklKbaAZHpACxE1RU3phUNxTDSTybN0dr4Y
2t3cUhODaTtGOMuDvnKivBmvpCYCX9OaD6JgNzIRzhYGkm61d+MIO6D0Su8HvFcP
85wEhr/e7OQ8I8/8jzQPATPTaiza7/M8Hi2BIo7Z2jP/33kJ3k0Uv3H9qrweg34O
GuQ1VlM4RESx7xzU1x5A4ByOQ0hfD4opO3xUnQbA+V4ihLEBw9sbSAt5tTDOsSmK
MFlRnDOuEVkQI8SbW0sasDGG+HuA9ac3kMOmJ39qTzwYu8OkX6xUo3vlVCETnUIL
fNsnLRYpwC2bYsOLwZZTwugChVCW/jm8RBCZiIlVOA5tyjhYXaKNtpq4ewRh+V8U
HndYIjnfp9ryhuVlUDQOok5v28TDpdXq46IfHf6zwgEe2GWoiSkYJ9Sg0gbwtkqu
ZoqhSqzClcQ0aW3NyyN9yly4n1Bp/DaxW69gYQmP4T9KZ/0iHpzUb+79vE3dbqTu
AHKKqHY0bybRxYNXbemguiYX+9cOAwg5CZ8cR3xW8oxkSJ6WLcSn28TfLzbBorR/
7mDfDk1oQPzBrjxk+4dpIj5NUFt5BYK9f9LZGMJlURmMPmdpJ/pQKphVlPYhQumT
HNSUUYXEtSapNmj7C8hVOgj6YXNpnkrhy5gZR7w3b3ktlJQ32Rx+1/Yzaao6WcZ1
WXIyHEqYYYPIYxa69/vOH4LjVtbk8Qoqa7xsya0HZZXlXXKUQ1Ox6ptJkBvmhSj5
1PtIAvIaV64Rc3FvQdr+YMxHiPw/sxAVj9gCywbVYaXNDBZdssxVNkwCobQ9+v2X
pSg6eFPHu0jDdz5zZL6JXQrYrF+GsK4f4jUO962G59erleexEd541idtEFQFCafn
dOEno9hkkXcPtWDkDdN4a8rLi+MU/0JIP1mn/8omwRD+tHsErJdwlo11OLwmUrfD
icFCVk+T0aY0JIHBvIPczU+eY3tfJOS+voWV/ad9lR4AXoiSEfdEGqbbFzBzTzLl
ZjgOmi/5IwrsdDfC5R6pbJuVWDDg29HJFaEGSklsAbFr2A94kgNWG6Ei06AOkVCX
OvlePAILVvv2sZ0XGJcp62EzFmjRiiSGve4boqNHtV/mRIJ5iu/Pe/ZoN5A46tfA
Uh2S0lrTRxdgippO5XpV2ibCPoxHd9ZIyFg3rzh5m2H92e0SKLYciJUXlpuxXymF
+sxCi0ggyJJ4l48T26oEeL1Fkp5hj/Xn/0NtmhhJjaUic38+FJOWwVp1+SGGO+h2
jtMdI92eEnYazJ/rmXqp0CFBAryQGyEhwzdo7kmW/1YbOWBQE+sDGSAwlV/10/AF
mB4AlN0PgpPBLCd+2BnpFdaLBBBJrXc/kjwRYeQySEt2lE6nNOSBO2CUAm7g3+ei
F7YJhFwaU5k0STc3vf5sN8RhpZ8P3nRh9Mjn6yPTGbVVblvCxfHE6gPPZS2ITNb+
KvKuAh+0vLwadaKDNrOjib6CqyrSJVXnntKDzsUZxSuQReAgYc2i7qejb4RVObgG
4gkZlRa+/OVlKWv+rD+EVwtR4LlFAY6la49vlvyhKNCUlMUTQZZ7hkFi7YcivRbj
in3V4/dFrmT3ZxK42fdePzePOWtXk9UdcQ/3wrGjD0INCW6Q2h10c3lcBE40rZbo
s2lXehMQW/YvlgAJyZw+QlNri5ngVPVopXm1iqOK6/QyqPrTAtmu1cPrUUFqMEon
QI2OKLpKQrjpUP2nIEIduonU5MuGaW51U6ZX12Dfy7oQ1D/Da6RdwT4eCasIJ3V1
rpSnPu4FrwtLd8+WTv/lF3FTg2EwWrkT94yMuAvBiwyQwp5CCGPSTQB8Ks4UcRus
uzuyVT7UzDrTatIEDfiWrSByKqj5bjEV1E8F1uDwpaUebtblSC6ro0q8xa+RjMUY
78mmAHC7/YxVcw4f5406K74hWh45lUlyhtuPJaSscX3pysGZ+lRUXXa/QY49xqXe
QRja5/C6dQUFfX1fUc0olHVJFjm8zBfo9irzT4C2Ib8ZRxhExl8i2pfoERrsp5Ap
+vJxsrEwemRoM62VivReV35lXczStJBk+JZhS+MvElziq6re0ffKdO4XrcW3FevQ
KPYuYVuiOvEK14nnd0K7rAVO7cBHAPdJduaN+9fUWKNiZBldfdgkw/iqSpZSPF5K
NK7lhbXi1LgUqjLUdswkOcvEsBBd/oHxNI2jm1+2vK4dTUmkY9LuPd0aogHzj97Z
tjU+1C3Zfs2P6oEk/bsrU+wyjq+2eML3Htp+vDEG38U8UZHOhTpRVhDfSXKcF2Fw
BSeDVyPA6iM7dXPYa+pmzywGOKd4FeX9pMc3zHfOAa6xKfQTUUxz6VXl5UY6RTSW
Y1Cg6M/HFhIc+FUF5RecKQRxdnTAE09VyjPD1cfkmaRt762EaRZt6U5utkCgfaBJ
r9sp5z4Z3e4Hk+TIUzW03lRZIxhXASBc0p4eTGkMsiE3U5wM37CgvQcfPN7QtbYm
EaLrcHbDBaMpgMBkKnipc/A9FT+xUXEKBEgBhEOAQkkBc/SmOVDQxX02QNDmMsOm
tdsOvat3ereijm8b+ciAZVzvJH4ysehqnqFYKJOwPEPMgpudkpktWHWPOnGoCC71
LA0MhSbdPLUnzwJ54z08sMNQRkMMCwUTvz+tUfP4po58Bp90e5Mg4AkuR3LfOB4F
dUI7DZRJohJH94OcMigY2JqfLHqqygJoQmNm9FsL1AIlLy7jbne96GfmtP9PRT0X
Eh59sw18/poqh2Eq3AMp3oodK2LVRkswV6J6f5KFm/chNTo4PohRqN0mGxejZQct
XF0dXZHhq+2d1Gmiq7CXhX0WuQJFjnzIw19qi+7SbWxJmlCYwH7AGnvFtNjBSTrq
AFCzqQOkaLqAzBRcmLUhQMaqSY68nUJKvIw1M4Uatm+N09CQgdrTineilNbwnfHs
l9NzO/LQE4eN9hxJ5QM51Zf77McNby56DHK5V2RWgFuNnyX4K6IXUF0Rw5hTYIcN
XNLet4Wh6bew+4C/nd324lwb0awpKXhd08vMtRciVv6v8jvcyLn6i9sOtJaiUooc
gOeUkpXa911qOFq/kdlcmfc/xMhI6gszP7XTAnOMswAOYfz4TwRmrfLw7gQRBg4M
34+0OzjWN6IgDYjW/kUTx2Y/kHIbA4Hu3xcjPYz/YAGjRR7tFFNmlJixMvzuykNX
DkEtYSF8xDvRXR/xuptSrkDsDd2X9+2GjwdEr3doAbE1GciNIP4NBsaOBJj9E34x
MTlBCcJSVew8o/0UDbgKFwaYWMj47Cpn8ZkV4SLhYTIQtBCLooaPyf3QD4F6sEJU
IQqOpQsGUmErx5GIn2pREe5oB760slHLBJDPRQHLu3iQLxyvT6Xe0Btjg5nBe5HV
bouShsdCewixMjI2DRAsCJ9QzPy7zozjglhd0JjEYn8IH/IermZc+QpYP3TXbwS3
f1VB0L+afuuCXHampXBSGiUgITst3JsIKkYA5qq6PFVPfT4cpGbnAO3YCdTwYuWp
aJrPDOZwnRkermtLGgFBsrf7+Xp4fpxThYJifmQz2PEYADw/IhUTEr4ADpsv70fO
BJrSIU9rrawr5Shs1HXUmu7rzGr7E4NOGWEIRrgSaEuKqwFZvUk76lyysPop5B17
MPl4yGC40nlxR1HnS/2q8Rewiogy8t3G4YveR7jx8w6kbWA1zpcj63ZagzDb9PRU
4IQ+g+mYkQj7X56Y7wRW6EY4U20CGmw/E1FAiYglfjC3uwBrYUi9uzkteO03C/av
Hu1aKWK4LsRHgJxVy1PXC7WmvquuvU/TRW1cB2pEAZ02OqPGrY014//jYy+2fv4M
07oW87mbuCy7Hh78QU7QZ13dDixk+xQLJm1Mk7nP+RDQFH/wXg2xDRb6cqdVBJ5o
Zv6Cs9ixGB+CBMX5g+lhIqtKj+lqYrsvMbOp8bDvAAEtYdzL3jX3FKUI6nehycPH
Et30DQM10kI4BXVGao64B5VR478yx5gTwBcKvSCCjYjRAEY+mwk3F+zrA+HPXZ23
D32aOaIOTTy31Dyl60TjPQJjyIYowmekM78xPSzvV+GkK9ieQvgyPXGsx9iyraPm
Gllc9kgF9n7WBibpEXzSBxr1fj14WAmWQNt60FYhrqQP6kOY8Hl5JNLdLhclRj9W
G4YtsLeOMNuXALjPUGgORDR38NwgUdV3NAkq9I132+g6y2LTiRdyctJ1dSYNTi+J
QOmAMGM6oxzcgIien8ChBT+f/qjjW1ArSswu6unqY2+2a9mx2GH+6Fr1JdCAMESh
kneQh6ivmTqIF3Iu9lV7tzGPpYXj2dH+vMnbV22AEphzSC/jqVjnWBC7HSP8zPnU
YAvVt6eKgjXPo3q8HmD69uPQbExZyuIRUmnXR9RtjCj7hxZcAtLA6DO519u8z9GR
4Qic2ZjWLFi96CcaTiJXdvufJJKMg37MO/nPH0QHUTsVHNH28sbhjly/FpJcruMn
g0s+fmPozCuwbm2NANfD7joTEo81Hz4UXz0+oPhWjLHdj97ZwGf1PsYaCFu7/nNM
qYehuGnmjQZLx5bj/NmLYW+wsYDwV3V4lju38wxt4qL4GxA3JE5+lO7KZPwshz+E
peNlzD/EEV2xp3f/9wwcfAnfxOfAtJE0vRC7FNQvae6mZntEluaLhPzKiBKb/GvT
NO/ktT03xcIm3wAVWbBM4MwNlYt/2q2j9kN89XEEEPAw8k3uU8FdqZ8SlIZp36s0
1vSdnMtRkA98LG39w/C2dAD51RZHrD67pzYJJrrC1T/Uu0i9WLxwuEVqhkGgpxCV
Yccmg/7bIcGGhXhXWMUXGWPb39hzgNVpcedpi71AFDThXS3HksrWNF/tklha2deb
CIdkYkQ/l61U4Eoxt4TrmPf07WWy4xXlGNEARyQgpgLkE5L5b4yWluVcx76EXIV8
qOAi8s9Vm3zy9PuKN0suGU+zFHWCrVL5C+0GJmUWLJXmhVXqlvxkJSMH4w2bIclH
ZE3Lxu2xHu3iOn1WzgGYaQeQwxmLbfYCjFMYvIjVjZnCON+0QGpZHPgGyQgSZ8ZN
BB9N2FqLadlzHZI7E+ll9T5W5x7bTpV3ntBroOMYFC2/iKilfsK3/GecuucEvk/P
rHIgyA0UZgazhKFwbgkyuJRnBbJE+opMT42w3xYTYvoN33OXrOS1/3fTl3IYFROo
XcB8OH4S00USgwe6oWex2+ygn7XlHMyk2Vnw+kL/irfSZ38OrUy8LtT1cZ4gdAvQ
y49y1UpYkUyEIJeIytIB142Kvxl7j+tg7UbHtorKLCTGz8Kji/PKd7FNykpbNuG/
TqBgng66TtsydZAaSozICcLkEEJViYsFNn6JiLASB0r47Fcp6o9xuIWTp9Da+DNU
ZATAjQ281DLeJaU3McZq2KmGTvZMmTE4WzKftkbZ/Z5gN3wxu8zOtCVJ6hwq/jgG
v1QsZrSjbexhMjVI67YC21I3TC2HvbeHci2ndkywg+i4rsircgj7uYJJfSAzwSuA
l+5LdppX8AWNaDZuLCNi4qKrI7wMiTEflEJhfXi2r+B3ztUA3pJmqF9ZGz55luiw
7T7xdiXDF/NiY8LhUeHux3pG06aheJPz0fMZx/6cg9D1ATuTQMq6wXqIrG34VAHN
04iKUF62EefqgYNfsEyi1e93IAOD4D8fTQHLE5j2rl32QIysDfCsawotec08SkQq
tPETIdCC089aPDikr7loPGqG34hxTI/eFjCytxkuXTTEebak68D3uy4TH0DVBrye
bTjqkg5GEXHTONCgMrOY9X/N4y4fq0YZp6R5QOjXrW9ddrGddXT6gsWB6SDYIPNo
1+JfM9mY74cXhXyCPWd3Pq5Q+R4zB5xP6kqXtwYfcwAoMsiqZlo+JxvDe0NArwwX
faaEk/FcoMaUl3KSO7t7nuQTmhaLK675JIhGV5pxos+QBK1Rg9udTy5SzdFwHvu5
d4SV9pDVyjKMLOvbGz54ONZHoDzSRsMt/uKq2I81m1Z63IfDoN3W70PQR4v1ihVO
yVFlTSN5n/67eSCIb05npqvaDGJW//TFppTolNbUWNFmza0UaQRPDBaIx86IzvdI
bwZFDVga3Ex1mlnP3f5BLLDpe9g7Ldz+PyqeuOLBl9KsMFY00CifFv8sbASYECIt
mcV0c1xvg/xTE5A/sXSUE9Hu5zzebdPRsz/SpRIck9UkoU16EDbWSg8Qwp9GOFC8
KBjTG8mDdPOQzMVOfZglIxBCurnJmSyOvVLrpRk9hOK9pwpDhzojA9ken6G+H6Tz
sYBGYej7HIUdR431KSQde2xZfDNCdL4n2lLqah5VX16Re0A46PHj20887uIlF7uF
rYRFPyOYGPuIK3xoPJfNhuQBRBaTLrK7dKkZKs+vz5+mI4iyl3G0uMIMcSz/3SgZ
1BuyF6qbIQMTCvavmu15bWD8EhWQ4dLJDKeiIRM+u6BYzD6iTQrwjV98SsJLsuYK
M7KBxPRsw5Yye+1CI2vr2PWcCbKBR/vGU+QVlFOlQTEfst0VD9axhV5f5xsumnog
22f2LXOe+m6wE2EpO1OgPj1fbuRXIolgIV2cXi1om99m42E9ls7GwKyKBgpX4OAz
qiOU83oKZF6azMyOQzUmIbPCH2ebx0JS0n0LhxRu7VLJQD/vmiN/pZh+d3JQS/cK
N0H/nY3T8WVWdTUCBLCA2Jlzd/M/cWscxj4fvFf7lcY5oBjkMNm7GBl3q/Ho44fp
XdsD6qQJYZJZWtQ8y6zs03ruwy0wtqKvwSXU0wmp/MzdJCRTaHmZ4flsfa73ZNAg
JorcOu4N0hh4l6AnTyDiobNhmD2vwOYmB2InzuUEJKSFnKaP9dH0MRCnUMAKuTtB
9v9QB+iI0B80m4K9BZ5f9+2r7L4ZmEYav0AcrhNsLk46yejnqZaMC6OrzFeWfmZo
fm4wQQRQD9NLp2Ry4xhfY/FSYpKSV6J6SBqGXRD+GaJMrThP80o5Rj3sFGTdvYnz
Aefz7xcfw7ud85ehqrhlveuT+AQ/Nmxht9llkG/MLAzrUvE7BRQy2yUU3M8rmS44
Cz5x/Dd9McT6Hvt2SCxoKu4/hMfiTXLTJmP3FVaN5VKaECi2QtPssv3tDcQ4syRe
v0CY9MvoDKurs5S8ZIa8IjSY7gNjvI6uP/tyI2x5ZZrKXDVRC2g8VfiAUJByp9bg
yiaQzk3uYi531fdBiJLgyPgv4rQrzlZD52EWrdQ9aLZdzcw4c/TPT3x5eTv0NN91
rUnWzsQmCthwuoLWQ9xLwDu+Ne81DM3V3RHKk91wEf2U3U5MupLGFcDq3gXJoB07
RdlE74LdQeGDottfidArOrLLWgrPesiVEFoVcyWVzxLGrDih+kQS8eEwUtOUoH8f
fNvfyWt1DJZOhhNUaO6ExmbEqkQ7DttX8EJJaYNXXtl+l3Tqp6waQHSsBU5wHIXC
BUsjAF+TjSybEaH1s0WCuh/H0l7WJroLnDaT9VxeqggiBIUK4yEIaa89e56YIWpD
V2C6qjhz+7RRyoIky7GospAsU+tdawTmCevOLa11XevYvSG9TRIJZlf1vclDOr2g
HyBz2/7sJpE4YujYPnI8fQvmmzIsrctN4FRPAwvuaAepIkjyzh8pnlNGDaTIZ9KP
9qtPGwwBBnjTLonRD/iy04yj92v+hDyYYW9PfvdGuqWJsAK9+SLe5UaotaFcZnvy
8xz2u7xSPchx3N+gwTRMg8ij2TWo6sWqEOaeZsI1M8wSMyl3Myz41lTEnwqfoq23
pz/ZY532d17DLI5nRhg6sOk2f5a3nL7VsM6JT/2s0/sno/7KZjp0dA/PVhiZt5BP
AW7aX7Jy2Xkvba1+k29jh3U4jZLgypGrT0KXoo6dsKGMzLOZsHjpULhO3AJ6oPKE
H8OBQ7aVlEyjSXUbQwMcYBelODXtyv2N0UvcLnjqvXmnC5EwIgAIn5c8g5ofr6n1
5PgGODVZZZKM9vpDtmit1UkkVQfuea7CgtriZEpqVEdy5oayC70viNabyTudDGqE
LB2wGJ1EtjvoVUR71kHZVHQPIkKYw2xizmKSMszUBFH5/9qgVDqzNGWthh+f+vhr
uDlKWo8+GAXTvOitAyTBWg2n+s8dHHCiuoJiF4qdbpgzq+qAQO8si50YYzbRD4G/
BEIu19zdpfW3zoxfrGbqAc2v1VrSrVolvUPlbMR2J3EQqQBXqWjE9qEGOHFNCngv
5rywzP9pVgpQBnK7Mp3ZfdBdTL4tWD8oQ6h+xlUTmsa/p9hoG9oZGCvROeViO5/i
hLEriaMmek9OMj94N9u2vx5s8mpCTUNqcNxeFLGPLrwMzJwr1f3BXcXahSJx73wq
Z7v/kY9W96uvcIT+Ot4Z1a2CcwxWy+vgRb10HTHsAk22wiXmKRoy8iKzN6QufW2Y
EmseJmt3FM9XeWC1+qKiUqLD3zxJQPvsoDQdt2ur+y7ORvrEWuvzFybPNhCHlp3s
XZ6pI0HnDWFw7zKxT8JY7KhD/kn9boCfNphAumqmf5mREWcsNIT7lwCkkqmsGyDz
lcwNZGSoR677hLacSeDIN8EAI0PSh4z/77Fo6og96cP16Iw/MMiig5h1Qd+18LFV
gFarub5saAs9Q6rfDFuqYFifwTTwbtCwRKAoztwGVxroBm55aXXFTPZoCD9NKjm/
7lf/v7h/xHd6RHO6XNeamAF0hTxifflQPhdYO0RE7d4UlrdV9z8d4uFGRL+38OMg
vrT2AMPy+9958krylmNuA2hUDH7NZey2iCczMGKXRTInwLTnuve1aTlkcNs3tYQB
YGL6yG903Om4t/U7nis1nRUjoLYF9bKHDBvc+0prdxp0aQfcVw9apIl3Tyd95R2K
0IlgcLPR3OrPTG4pKsVLtnsxX1+vKX6DQYmzUpwcpYWS3HPqn1JvxJIi5ofABfVj
dzFhStvvMCJE7Lf+RHLIcwz6Oxlug7YqyIGyzd9uN2tK7g6YkQTYbk5pyZYQyZrI
+mDR2obU2W7AnMKkee4rQ/BHuis5WmC6Qzjco48DJ/btZnKfuAWb21IxfKzG2RB5
sCS+voU3IzHyHYFdaacyQUOppfi9DZoe3wJ70VZTZ3ZPbkXLbtHCeC3cK9o1Xqdl
ijJAjGO4sF9PttKYRG7AcVQdTWiL+y6TiPaszdVm9CWFx5qYF5j1Ed0q4XzzWeeH
N3E43BctgLXkOovPNktMX9T6Zym0VZ3R6dLbMtIBSchanhBnUDMCv8/fi1jrOHaC
72jCKhomORf5r1q15v3jGRGmTXkwJCb3bGauNpXv46kERxERhKsJDDQyoQi4DNdb
6J2AZ6UtMeS5SQLy3gNhrmHOUtgXy+zO4DcyJDEJfD5ttswBWpDL4FGRPULfNWaf
eahS1JSSJmk8mMKBF8e5GBlfB6Fruyn1ilA727G5FaSGrPgMymarrftTTY65ihc+
uK2jvAJOTogjMpPVlvHbcS2qWbqbITiO3KJEBp45l4CEzF3QcVvL5QDlbp//T/qD
oD4FyF2J9CuKRuEy6nVeqyHVsCDxUA3m01jVHk81RKK6gkgXlYPktw4YGJLpRZKI
kVErCS/tYJTLhIH+mXEScDi6nT885EDYa2VO3YQnZEwS8w5BxHLZP6IRkTrWudEG
mhugdXWgfmGr2eAEvivDRV4ij1VfYAOkY7f5fa7ZkBPjzVrnjQEQ+WOzaew0/cpc
IetFCVo+BDpT5ph3ClkxwIKjGljR3Ya00k0fZ+cbdYBQ9kyGGBMW1QTv0okjP32G
WDIKZx6U0yGYTI0wB+biTtsJ6OjKY6ZbjP5rtbPuZb1bPTxZHGQ+vU/EM0NiObDz
ZCnkXVBTMOZ0JoZRLZxOsIQ5rmGyoTUnXpOLHboYG+XbQzzGqz0CSqTpddpnrh4F
81k2a6C1EE/uSHhEytrpBEuFBDiWa2JEC3RJLNjaTozi6KivOOBxS13p7fQUTHe9
wqM19TXer0PYCeaFJyDnC7O6UUTqJROWrWMPpzGFJI08VK8DdCZw4vODkQJU0qQW
RmPiVNplB9DQsyTbwWY7+Gk+qVzKmPgPKfz4iQ7hL7Q+9HR3tK9INH9QxrE1H5fs
LkpGKNEt7vRa+OM+P1GidiMUCy7WCWSIEXo3it+FLjOHrAU4ftR3s15hxFuOM20l
DMnO5zIYqdbWRM7grnlIjxurr4X1esoxi/e+ioIAj8UWz6ScD9jt+N6lOYIfDBKv
VLD6cANw7kJZGBnjxjMIs86IsvQOqPq3LrGWSYhAMcbQZQyhST8gI58G6q3e9sdM
Nivkaao1BkoGI0RFQ6azNCar0F2+3s99AIeyRrkTbqqdAv2lamhzXIf8cI6Tg2+U
y2/CAifttgQGuOmiur3M3/GLQ0CFyWhS6X8BFN29LffIq2bMUBktc8KSpZ0mlRPU
gd2Z1zffq67xX6mGe5zTbKOJcuwwNLhBEaA4lG0j8eyXCUmAmrijKx2a9RB9beQG
KB+GHnkrpMSjkkldoQujg7ZRNTlCtu0H7poX0ZEELy74SD8i4KhY47XjpMPoQl9k
6YjRUEwR9e6y+eXk4FDa99SeCAKczvCz22ZK3+KF/8m3YnsnDNylIFI4n5Fp+IFW
3nJJl4yrTPkLsSwJjvlMZLRukV46Aw5W+9M/iT6Gt+9ajytkFEEwo0qmjlXiqmjC
a3JbVdQKy+OFrslvtIdJ1BZ1Th6qMUZu97o1DVxnouszz4n49hbSr8miqc6s132y
33o5meZwGT4kvratAun0D/eSQXY058xa3QPoxYe+3dilJJ9PLhmm/F6kJxZdHqga
uS52oAY0KaTxL6D2GkFcFiaRHGzjOgSKZfqopUlJ/+FBJ+76mdS1GHVLulElIlz2
S9Po13J5f2U8k89BTy20Fh0smRVbjzcO4n7MrZnqp0IYvz9b5rsnXvwIBwJR8Rzf
9432wel3zomTED9Otg7DXoCpaACcWbMkfRxSR1Wc9Kl3+iIK4CkYGkSe1sTqvhbf
br0yW2W9F07QsXhKaRmhB1BnOn3vKxCxxTg4H+eFppi22OLnZbeq4tS2I2fr07XD
aKO86/kTlYdPcMliAIe4pCXO7m/HRNJXcoviovHFGO95v/ZYWxVz7CbPWDrtg67g
t3CBPH+2LqkJYRkDQdpI1TY14Es0Yp/SU843JQS15nFhHSyQONtUGD6gvOtL6734
E5PIGbPxuLKY2oDKiLbp2brqDGdyQqUAmv5+0HFuwwaBeG6wNsfzouvmG0LOAx1j
l9UFGyj79z5pxpfZ+CchJ5cj0LdKdWR2evWqrEM0cSQ1KyK2Qb7W9EhREeFwWZKp
yp6/6InA7tjdCgQo4NhsIFWaAxQWNyRsjVRjxHRozKYcN2hVpUPcFRKb/D0TjmgC
n14f2g8kKzj+JOkBKyZS3iqd0fobP24uugx0fKR47NwbgLbCxZ2OEqxzOsuYriu3
Huqa0v6NJ35Tlt6QD45WVkAhXSEfbB2ETet6lAdmZL0Bloe68wTZT8VOAqti8wzO
pznqag+uuLnK5JXASPZjZJgX87Ei+UAASnTWWn5/AlPvJmjLco9dUMt9A+UNQIdK
exbTANK0BAd3IEyGmofJcxtqUpSiLrKcPYsZtz8XNmAs+AQ1dSo7Xg7WpWJFm76i
L6LUH/4miKm8zJCkdvsgf/8oKzT3hR83jPVK5dBJmEHg2aPkSl2WzpajRu16pREl
I246Fkwoo4SKo5EBE9KNl5kClElvLoN6KimT9TNBcl+KPnCaGnX6U1EOk8h2NmbD
11HJiYupCvPkYh/Gyo1Qk5F4hIrKr7krmrc/Vg0fSWrAW0bzezxyHxc/9kfDHmLC
iOdKGzoiQRMbhBJ1dJvnMgth2vTwibyUcQnfku0ckhdSKDaAytR47vvjTUJGzu33
uYWwICWi6iDpxVfskHTt3x0A66BN2+WLGZiabdBro7xtO54qlT4NgEnXeFCMO/lQ
TfVTHMv1t87qQXxXn1n7F6UOHpPqdW2y9fo54zBf2dlvqB+pMi4tRFiMj66HD6ws
HTq9Tmj1PRxBEVEsx6JQiLGu7Py7BoIri1MjjRvFQOrBj1fmdgMCmkpiYEHarHO+
UEYwinVRp6h1t/iwsKBXd5fnc/ajJ48vBOKIVIjczE8IgET6QAlnvY4CuuDUSTea
BcUA79pHKYzfyth+5calvJQyPYo3e1f9GBUTD5Wm6YvmRLsirGeqeVRtjeziLqQ0
FKMrUtu6HHCMf3NkFAWzebM0Go1H2y/7wbk3TpFfSoBvGfLDOF7qyWw5I8WSbf3D
r4g208RM3ncKD08q6oawAKFubr0S2GSqBH2onsvdXo3p9sBAwBCEfgMSAowXZTwL
HDE6MbnOf6/3L795Evyl6t3Z5nN6WPPRtApuk4EjiOOCMNiJZqV5Zvgjsbh7DqX2
7BCMD3w2mQZ5UqX1XefU31gjhBDhZmI1akIqOeNCNO1dCjgq7FpCP2xXHBgRKXaT
HanIiEDEjr2NHy7SHz/0geNEq6hP4EnR79gmX63u50Om4L90DqYZG6cSm7W67Y4K
YTDVXRtoL1lfKbtGq+XTlFfWu4pVTKUrKD0MksOFw+IJUPKJ66mIRq6gwU0FWtub
lcD1wVeCadhb3TOG5hMLVchlVnhe+h8p1RklmXRBg7LbqrBNc8rB8f0/lWEn18+4
VbeXveAcM9PuAwl2gwosfaBLhBXUnIQQ2kEkXgNpE7kYdfkbVQ3g/YpTu/9SKFFM
9ndHDYYQ50/CjHjYWjHags0aCMo3nxfHi2SunInlQvRv4w2nIk+mplU75gcFP3DB
QOut26Gv1cR+X78eOLT9i+qmof0t3kRF5j5wkqBOKGoUExcwSqd7tswTiYWq+pd+
sQ4do/ea8zjm4PP+b3++Hv1qoLTxzslEbpjfjRYwmrLfDvAIpWaO1OBuCTKjTyjE
m7kKiYotjn3K2tkSgcOaLK/Gd8n2Org58G9qkKknTZ7ocpJvwb8AlpcsUscSkOWx
sSJtimcCQSP4a6nEm2wLfv+U1HMjPPx2REFpUhlF6nMnQmfb2YWDNFHzzHY52ufa
MFoWkU0EkM4Dsl0awgdgAAuSQAhChryH181GVrqq5L2xhyqRBPiyYdlvkl0jouZc
cgnSoy8I5se+0oEJxAfb9YlfPCXoFljmVIUBdw8P0QkB8i1xAJRyb8eqqdThSYh0
jbitzDoNwP043R/hZ6h5hFD8gHXsf1uWG5hPzu7L9/pl5E/jXHxanUQpLok36atj
wZpQl7C4NiGYbIqPqzBNz7EEB1cg4Q9GVJ44HX6Amb9Z5EeWeITsGQscjFIY524a
xUI8GkJcRt+g/EjmxiUPO/3vJHFwnmIKvtLsrTHyRoaTMFMyDeYz+RN9BmAHrBpI
RdcVvMEgysqZXZ6lT90nbxu+v3zWKmQ+45f1zVfj/dN4hf+q1Dv796039Zn5qTeu
R/7g6uf3p5ao32IYN3x5vHzkc+38jU0Icpzs9tV9jEULfvDIZ57ZMXtBCIsZ9NDZ
0mtZJtOoUmubp1dm/i0ZEzvG7JKfHqsuT1nMzgkBfWhaVs7JJg5B3DoQaPnMagCc
7xWuNE9BV6e+hkKeSjqw67NXubfxDlrFpl49GdE7QtS8Ycwl7eKnRQ27VPFEqOPJ
LZZiKao3lpTXZ0ux3kd4EftxY2hbdAl1s9QxxJyAgriryfPPEVEP81vniBQVzdGF
dKJWoCCEcK09lHPxFD6O/kBuxBsYgSpaQoMqhTUnIxoMT9V0CceCTN4WA8YjNgMw
INPucmXutVW8T+ne1ooKil8/GpbqwkbJ4Ab8Y+I68cv25bROnXkCM4uzgrSUSECy
hxF30EmI34YNjdjK2M8c83EOmHHz62I1rsmEUaCnMITiEpcXqHOR0kIxi3wZ0Jfk
5PYL/GPdeKIUuDZk7UnmSmdPHajbC/cp7k4mvHpOiXY82RParPkUlxwgN0P6RxHX
u3l3DJgx6vUoWApoQxPOm/r1ps1Uiekqyf4Li+tATxGKsv9NGs9KXyshB82Pp2MJ
rW1D9Zb4E1D/Qm9PzgMgNTpW4qctH2K12/T4yKUMmAKOT6VvSak1+2yGgGoyQwdc
ZQzw6PIR7z+RAHsyg2uNYkoglBoz0lfbWrhobsjRM1lcp0OK5swEjqmt5pmH3kBo
5/75DbHC19VWh7G3a8ede8dQ+FjtLjA4sJRQHKzdykj13CcU/s+Js20APmhejf17
haPcWhJBPmnxT1gvzGkNVYqih36StIwHAlZXf0fLE1QKqhE0EL8MlPxthkCPPXs2
1hA7esj59RNFCR/AOSeLYlHvuG9wZLTHOMYoQMqynX7xCLZqTnqg6cK0bvG416P1
DmG3PbvTTA67cWkWheDmA6rr8a90MCWZLCAz4zWC9HOuEhN4XMIYYXBWXY0atmIy
cUT4o4PlCVJP7MwzVd8JpYRiCD6gjOpsgP8k4ScBTHuyTv0ku5pecig/pD0bQBAQ
CmZcAdjAkkKnPNYNoXXaQIkLqO5Y8nrnTT3twKtrhDtQLTzDW7/51DXHLzvNnAxO
VvtDmKzJk1PFyl/7pCC7Il5lQAFHPuGdSVD1iJW98xNh1/2Y0Hs6M+KEWrBOQhmx
vEb45vlRegcU++AJ0wYVC1v8JxCdWRz9NDUi8g3tStpYZdDT6Bzz+cUItxPtuFoi
gr4HBxeqVxq0yN5ZH5nYW919Ev721Xywae3COvIP94rOIUGhwvQ1wl4s++w6JwFG
GHzTOECmS2WOvhka0XcxRdVU0TthT7YRzJ26W2pcHvY0j3dIGRyGGj+h/1CVOHE9
z/51CJOzQc1AoTkj/ALwfgO8l4pbe4W1r4wDd3r7l+jyWvJigC/l9h586VQCP9fc
B6nWAUzOwLTYIPCp1oz2tGFwfJkhL5R9hmAgNMYI8yxXomzMmUpU0+7cFcCqaU0d
fTZpIL9DeO4FYPzajaSfDmcOl9HSxeSZKx5rCW61j8d2qiwpdp7yj7PPreBytUWN
ZJV6oQyQskBFSly0GzSHzqMYjIERpDaGIJN5Ump9Bi38UJIjyrLN7Z8H8KYzXLtT
Dm+QpyckQ7DCLcpGBMQuAZBYi1jN/8IE00zbSC5SKsqOqq0FqgfvrYVNbMZCmoJR
xnC2f5YaMrEeNYMMdLktbOdqMGQj2DH4m7W7PDUFLYsZoQckSfRA3MDcpW2USFOK
EWre3gh4PYcNtlx0EOatanAUiV05m/Cg3Z9sXhWNVx7tJ0nqDpyQPoLCG+y/i9yO
Fkluh+dbRY8b5glpQLSF64Sl9QDO4Yviesv6hWC7+nZrJi8OMH9/83fimD6Nu89X
xGpNsDi0qiB4yx4q4Wyk7j12YMlCZTVJoRODwkITgOUslxNHY1Su3GunVg5vCWBp
gvtsEbkhcn41C/8N8xtJXbtBuVkbLEEzEvXCzsRnHvWO2SqN8KKihYS1IoY8f6Rq
0DLZ8/IpxbSWyH093hJJvA+TILoTpUAmugtb9VeHYufT/4tDm/i9FisA9vxlZwzI
5jBV9eDC1u0r8tsU2pgqQXa/dvIuDlZqHA0F9HpFDtEF8O8ouS1Sa5AnImXA0LZd
H0TsWHgm7nt12HjNqApfunw898cEhEGLdCESrrRahohpdvQgPMkaOedgZz3tXcAn
lZ4kbizjJHG1k2u4LYG/gp4oQiDczJrdKKmwdZ6nE8OUcd8IZGyOrT/QhNgnsSNj
Pluh43GXx6FKikl9IXt6GaKdf2QoEsnVRqQB4FnBZyyE+/pS0ZhgOASORLH01sIV
/FOI8TbLF729NwPXBSV/+Me23iIs4xSfr4FiaOJkVjVCwyriVDVEA9/SQZJjaiKr
gjfEdNXk4xE8DGHZBKipsIkZhrwRRJPjkSRV890V3e7ergF7lnlewviJixTsK51/
wlFLKPk7mJdLurNKo9js3ijaZgtmm6F+5vsLH7bg7ar3bSpV9wsHmpTPfVQhwSZm
D76XSADyy3mCRunSNMWwbDjA/JpnHojj3mQ1hwyScZBebxUPrbSXSwzwCofgvqEl
tXX3DNECAwr+dOPaAlXtFfHOsw3oBZKWrnAib5I7n2+m7WNCkK+DsqM93Rs1IOpP
Z9FpyYU2eIe8jHLoUSAOTnew35m7Pi9uGwlj5SbKP6Y64DIJ4uNwz4uk+HS4juT6
JknVTKvsC/W1cM0s3uuSgrEHpAxN6ar1+rtkGnkYA86yUXA6Gu/+KwwbX+Cby/f0
xfqlVnJjwdNSiROQ3Q3Fm3vQqi3Najq5o7bs3LG5uTT3hk4xeWRg4rjkv9nZW0FG
1+cc2DQVMvAousoW+5DkQo7zXBLUBTyqO9h7cmy4pRb4+ljDFRX7KNcDopPEdr0H
m2lYuVzg61SdgFzqpStEmtM5zL5gaEWbXQZKJ/16PeKOUIgTLW3bLUbB/Q/fgg3Q
YjHY3cXsdmTCSgzxXvr9rV1pUlGC3PPV3h9pbLzaTMqlcKiX+faPgvbgX6V6a0iG
7HbsrVRL1xXKWxwXJz58BcLlaUJ+oBT50ez1c8f9UEJTPdT2tZXAuARo4UKaUHdw
l2LvmB87iEdJWZ/I+Zafnd4XHShxmODmc37QiS2uOS+HVtOf1Vc5fG5P2E9OHRIJ
ykukL5af5oJQ7zLChCq2x1w5UdDUoiAiIa7uuZiHRADKUWbPkkjilKbN5U8GO+3b
BSlDLEa3puy7q0U+yHm1KT4u07SPv3BsNX+rU3sYMKKwn13mzUfiNIvMe2vo4aFb
WGqk7BWh75Hd2lz7JPTPRX6YQqFAcPGWVB+wb95y2HAr8xf9zw6L3q0Gw6D6k04J
bVECGS1EdSWQp/YySkQZ7FP015Te/JRzSG0/FOF+IN0gerrmogVRlXr+J0RuJaRe
3fhJrE3A6lbLpIiur1qxabOQH16dYpW4wzcW/3LUT++67Cui2Y5nIaXB9291kAKR
iNfvTHNPL7to4i6uHLJe/o1o9daRV4104UcLmUAU6E5Ob1/5n6whV2Ojoi3jO3gE
rebMTtYVFxitYq4GuOSHs1rhE4ToncvoXFo5Pf+9fwSLmPJ14MxVhs9Rl5TpgRiH
igCr1BRQUMvSy9vLvpB0HyUXTAjwVz2PAvLITpZr9lqZddUiMX7sKLawyCAmrvNJ
wB90YS0UICNxEe74v4vEIoyfDxCTvrVQNcAPyr1c868DZBU3ajCvDXy2Z3cSE6c2
39SlgcLK2gSaLG1LejqqSVcCah1+FKpX6Vzn0mdM8SuFIf/F9hFOev+Pmu9mk5bO
RQmaIBJ4RncCYimoy/O50EuDVZA3a02jclUgyScoRSW8bxb+Blu3tcDiM79RpT+o
OKjwAlfeoMvgC8qqZMEuh+b1uD/EO4/3LQLzOghSwo00z853/4zbJCAalqlp9Ag9
v4bqXP41muKoevNNSF5XyMBkE1uz3b+Axsay7hdRnMmrc9bNrvJcEt/KSxwu6PLF
vjbZf3OvEbK1rKTs3AhMAeFKxAnV59iOh21g6642Hba5pIlRt8vgd1Arz2f3YbCz
uYPkMrKqGEHnkdBiUUGQYncGV5Zx8onZY2iK3aZLZhRn9OAiRdkZ4wbVZimMacjW
cJPZW9Xf94Km7BOifKbVlIC5q08qVFAenBdi32SRhAF0rknHp2Ygf48q8mh/uaAc
ediqIJ4xAO0UQyNGMEf+IZrD/ZVtVHA3DweVAMUe14b1U16/m076IMsTJFq75fLR
2ej8rxoFKCrJ5XwImgNdqlfWDgWgRIfCDtmFFlCbI09tPJ6S3IOBMJogzKCdCWeO
y5Q0H7dieqrQiA22hDdOLiOBD7waWzvOFkBPK2p1PB3qZinfEtlD3sNql96eFD9z
D6UIaRrgRQOkkqLZ11hoBv8A1Bhz7e/VP22KbHvlpaqEubtMiz/DV7wG614t0H09
dmiWkRp1Zf+vtv+KcPd+HQHovsc0HnZdUrVRiSXDZKTmHx2/OBoWk3ybZQ7i97AP
xiFwSmQdjiWrFNE/YiOsETuSiNRyZa6vxN8CeBygJBlf+3WTXu6ke0VxdQcd5qzS
RNI0qez3UrzJpMdgn6b2az7iXzJ7H/UaC5xsUSKhRJRRTCZOe19aVRBg0M7s/lVP
DCHKqOoILZb5SWrrt0cUz64jz8jNjYgizk7YCyBH6DNBXNhodkD9saMRBp+FawhT
YTz1hT9lUpu3Ado+5yOrBWYcgzFM8t40jA17Bj3hoUAKa5GHqHmwWmy8HBfa/icP
6V0HGiXZcRcGGueDeJB1RVbQ67ogZD6k88R3AgMuiwJmg2OeGlJoRarpOnOAD0A2
bHBNeChJbEYbMf3ai57u1y9ANA0Wcig4bUXHr91B1PiKBub0I1fOUcDu7fc1+XAJ
IVVQ32w9pfoBGV5tf7fFRp6vEoiJn1R8pfcy2wpPR236JxbAMA2D16smL11WJDzy
Upa6NLLnLh4ChY8Uu2OPBmBgO/hGsWGaZfVNDT8G7LxG/MUggsoJoDXOIfnq/XpM
uBgeBDfDDqc3dWEBDjjMffuD+TiPec8Tqj+/zg236TGWysi/LNrZ1z6zZFxE/65U
grpiIWo0H/O3UjNpsY7uCEcIgsUMa9CGcJakIhIVOsY4EHCI/OSoShfOWHK/cKpr
Lid25M1N3GFaHUHwp+s5B/UZPXP46Ca+CZ2jb5X1Sd3nxK3KlyG72cqOJd/aUodr
DueZCrmO9NyVj2myZs4JFNsYXEPNTuQvWm20suwjlZlq/KqfJ1aQBrKStKGe0/Sy
86/GKzhZJXsCTlZnf3C+2NaNl3GkiFyfi0aw/vJGHWJFQU6KgmwF6KOJCSBpsNyU
7KfQoRsPKL/pXYeAo7mIt3t7fewOWSrEbhZQOiUaA4NkZcYw+R8BckTWN0kP/4XV
zRCzrL/X5qEuM71pRMdQLwoFWzo+lGU8JX/cuvevDXKtkhQdNItXrhzWeRX4V8bI
3RBS/Q21VCvvpD7m67K7mhdTR43npmJXVCiEE0zaZq2np25s6aqbA79Dd1ovBMkU
hnnTfQ3mFHsObKjH4jR0+cUgpcBCg7r33/cTE26bQmQH0Ecbhwg0l7HaFQKMGaSU
JEvGTvf0//2fUMVO4p/SxyWukNcUVyBsLW+tB8NJm1Y2pVpgYCJjelYBpe4d/QhL
tGAHy9ArqV757HXODspJiwuScq7XY1qNFoW5QHj7B9LUUggMqd4plVMLuI6sDnjc
HStwfT3Rq+Rt5OVxKlsWIQV7THYN83HnguyuyNq2g1ZLg5Wleq5GQgG0CmbEBuui
4HbIU6KrrEPpx4IzfTQs4p2vg1dZlfT10LhsSZFUt71GG8P9q1ucnfAY+fgKoKsI
xCOlsab4+7h1qmmLtlCWbr5EgNwfSPzKX3QD5ErlBIAT1qQf0r1R5wSsI6T0fP50
urfqpftLR3iatgjmkuUlbRqqmcNWWvysNRFy3zfsKHFTfEHaw/vGuc4XIj0lpHEJ
zgCpHkjiAHILK4MdgCjzrm43a6FEUBVdSljKgcKdGXYgesMMuMehSQlVSkimcdue
hmZsFrckoJE+kxLsgDv7OY3EBHa0gVdOANHSSqRo9chg2ILjODS42xVKMrkxrnPE
Iu9BUWXb4y7IdPqCwQVv5vq5oYN562N51A3UawqRwtojm3pZgvaFPa7hj+DW+1Ha
UfjuVE+jo2DyeM/Pvs6pX1fu2IB86LS9W8mXwkgnhXLuGVEGSov9pf7R97eazlVj
q4mn9Vn7d7P9BxBoLTtYJqCdv4U2O1ELsrPPQgngoJGrUv9JqUDxp80cE21Ch3Oc
j5mrubH0zWadtIZq8otjZImy3wvkKJNCWE+0x/v54PJL/vG/DqtyH/eR6DJEHtNV
bwNyWWlB9vTWZuj23xkB1ZP0AbvG8vONYyOa+VDMpLFxamwRTkvFgAAitEY+p3NR
9KBHQ9/t58MGruNbF1Xv+KFMy94xiXS1ZzEd49LpUNCF/z+PyDrZO8DzfM6a3yn9
Qf/6XgToIJ+lOSy6/PgdoI2wpUJ1u5Ic4E9YYeQM5YTD25kpGcwRt/dWCySK8Dqy
DMUZsIMFreYbokfBGQNI/YdM2RhrzQwrh5FzgV69zxvsPXLYWWnFHKB0WxsnDQV0
xzaKEEc56/fRfz+DtuyUp++q9iGrxLH++ObcF2Tx3GHYX36DymEdNHOArm3ia/J5
9+2lg9k9xmBl1LB01Ki5mQRRh+W8O+dA5oYWM8l+R97ewXVxyjQ9KHun4OGIa1ok
8ScUsjP3sfHL+rFkenG3YOvg1oauZZY26Q2nDAGf4GJVnbT0396sTsNNcbwPP0hz
wz4T90Ff++O960oUVF0xM19d7Wp+yvyDhcmFGDjSneY93GftqH4a5/ymrYRIMRqV
xTtR8ms9NYOcn2xCTh+D/+4WZnt+9Nxeq+wQMJoHcagqPcz5aT5UZ7N5Bxq4s+Xg
fLRUJbaF5y5sNGmCNGDIffIHgcCVhtGhay8+8AIf7p7C6n1kgdce2cUYBYXuILqI
TwBHrZ+9jDN9i4kvNZZaasra7jBQSkd8483rgbcYYeIh535pPj2BnxXcLleEdIEz
NpOsX0vV1IpFTr2xTubnWUJLAJFI7gGsUY0QUJdV3Li3J4CGnHki0o6K2tHzYFeB
bQompKZr7v8bNDpMLJV3t7S9CoYEYbP8sTv7xCsl6kY76VXf3xf3Tu9MqZ5Lyxyc
TLHYf05cTKXIV5QHTU7MfeNBsNvlmlx+JmqsRE0A3kHMLiaF3YeMiROueU/4bwB3
4guLOz4LtTlj3WtArn0xVP56I7MvDBcMYLpYMkajDJLBN29LKawxts/aMy5dIT0X
IG90ERRPBwIbFnYR+C9ggNW54yKDF6y0+fDYvcwRNwgKK22Buq8Z6vLynn3+yXlV
Rbja3J4GJjQNoMcqU7fdouVHVaE/qHfCoP4sybCNUeB1CM4q5IG5uH+IZcF856L0
vI8Ii1FgGB5JeyH6gaWR2Jntq0cSKUVGeqMqPLMWe9iCxenEEFxi9lN+vo1NQmYj
jifYVhUPqZCy3Ve8LAJjBUh8+oZiaxTVOj+tZCAsA+OXmZF1k2r/5fCr5PQKXq9q
lIkg7+V5EBATPzdOdf0m3Kt2VNByMYvR6+LBV1UPfiddYhU3TP3I52mIvmTEmTiy
OFlO3n6ed70rNZ1CQTdYOi/lPUQLabCVpUTmfODbbd9ZV83Ao3n9er8pLdq2cL/m
uIffPeRfudDdt2QYh5y+59pzvPrI+nxYeMuC6pcKNESteml6iI93smR8vBrvqhmp
rOphJDEoXNVL+INWGvx/+DD2JoZQ8zH1yhLpKB4E3IRhoAU4V3zhjL2zCX/tHeLv
5Ebf0S9Ub+uZT9rbDT6fWvn+wEj7d4OSRqRV6U5ssilr73FAxso+PLOwx+Lsnvk5
OwfZFZX8AN6MCSynnZ8Z3QjlsoGyjTV8JfiE6SMsxLfgET+fDjBwKUOzt6b3Z8G7
riX9eSN6holSZOKgqNSGtw0skFP8aDQK7rXYQoENqwR24DlIKlnB250XKcXS1v4b
ETy/e+FdP/73v3mhKGH1U0u3cxDYwEyTFOp/vUQtJhaCe5BTv6vRYhx5upfOAx43
gmrZA/697CSd8EcKeP5Fw5kF+EwND8F1uAHBycsB4lmMdMl5uZx7M3xgq6lo9P0B
fwUXrtkn/boC7dTZ2tYTBg0x0uhXMy/ACHpDa/6k9VB+E1t6bAy5zqCeE/uwqOpK
d0WrnBrnov1mAojT4zi/5qHOR4vcHbgs3eWGA3w7yicLwBNNpwbn4kUverDPD4cg
Zu5j3LlJdk+nXjaR2v/qA2VOG5WMleC5yr19WwuBr3U+2rVQkpiiWyKVqZwAM31u
4XN4nCIgsHw02bAJnNR51kGiMvKDYULKnwJHeMO3626c//shYAB3omwHJRrGLqGl
dPuUbAWNN49ZGQe/dtoHdl9zhYw9N9o+mf7L7OYWoprbKSF2xDepYvw4oHkrqAg3
z9d0xTCYvmSHwXdwphPG6QmwUYKcsh8rrhlBUzGqLMwib4MRz61LebPmUGlp+xGy
xZqVHaMCV17SkBNHy44xKIlAebDjBoCVvpJH+mn3mrAq0GJqTwHfuG8Du64tG4hA
ffSVTYGcePM7nRAoPPW8lqvfVEAT/0KS26pmnsFwTa7UjycNeNzF9BMFfu4gpr6O
3WZDre04AtP3kiH3unUfRKGy9T+9VZaGWcXh3t/00T3sbQLXoJLxoUyYYv5ZU92r
iaEADwSTIxuP90WqIEV3A6nnv7HuMWPGrihFufj+WUGwyrrFyI2w2LiXi+r5ga6f
hHiMhPt7CeOYx82q2rEXiQBj3FPvIK6K3erL560m2YB3X2EGRE4W4alRtz5a3kke
2aCOrqNkgqAH6ShPwPunVK8ycDcRIPaNiOB9vXEsWT+WeAQbWGj5w2fRhgSlpM1I
QIEvbmyE2iF7Ik4p3P1rJLNfEAGzDBha1g3zzU4vUWsGDPVSaVjpxH/gobDcIyVf
RvHuMdiIiuAFQ0lBk8zmk8ZsLzkr/+28qPLg3zz49E6qJi/gfoQEj7QoftjlV8A0
R+HBLGqtJcqD0kt0IKx12vG/Cxqyja8FcW2kzKSErgSiVSH61enhFyft3CM0VCoe
Xnr7vimGjRsQNr5F1tXWz65QUQYIVF6BgsXTG9wle0lTL5K+t4iPuGXl6iJRkAlx
ePvaF5A9jprLXWaNz0VD/2AqHY19wG86y7MQzAC6kMOxdsXV3QNtRj/bPHypNNq4
lPvlLQiB4Tz0p+msBRn3qayKpHLTJDYNFikVZ/xBuj8KKCtf2DhNk08mVmJchizt
6WHTnKNiW1AB5dvwVBSPeHVonViC4r7wuL8A9ILh7U18AAG2FEwNcDW24oEhrM2N
LaQLXpF2MOR/okqoh4F416cO/f52VfJxBXYKAeftGglsbJsvNmXs4XC7JE9EdAF/
ZTlkqlEo9jaNchtS0JJmH0X8XkggQFx+LvHYgpXi4p2ZqxO3mHGdhXOoz4b4bXoT
cB9xionP0+E3g7VhQei7hYLYe6Yn5len2rdjSqu4QfAH5ILGv39sJCt27QYBqGNC
OBPq58E2vd0an2wh3TtP1idOd3dDQ0d0Va7WOXyEAzDFTkxxi5mvqod5g1oGFPbZ
KEduNV4v1zougxpUifVx/i7SrYUHj5a8e9s/lIsA1oqzsV/QxVlBBi0z3FZrCuxO
2REP1/GnfCZzxb9/RaBURj4Uni6ewD9biMB1ai9jIdwXA8vbJbjfPfwNKSeFZldZ
JmC5yhjjVkNAuqtccSSRnxYf/lvzqWsRvJxYYbQvHjE5rqEKTAl66+vzfX3ar018
l2Frb75gOMhbOqzyfO5I8uxas1zeY/EGxDaJV48v5dsOXs7URda6RUra1VMDNDiC
VPc4Irt0sgxOcxNPW8npb6tPE8rXwxBfqHetJBiNmjhub/3I5eMdCNdzwMW4QrBW
U3AoQOiR7m6o52KwYOKHllNx2TaBpcwRpiO3SSSGiZGtb0TcnAJC8ZLBizsMCudW
51WeWZa8OgPSnsn6J90Y1FyfDV7CpRZV+H0xdxUDMLS743f8tOXJdealbaV6Qz6V
6viTLyyjIT2WzvhwZecEspZvIzq+hXt/waCK58zIXfxBNqMFp4A7CMpECrT8L7qD
BI4HNQGDlo0nDNWeds3JGx0szxntv2zFpOPItQESrpo+4z4meBO7DEDnmhjyWuNw
u91xU+LnXHYZMlRu6Rgr4bpNjN7WNX8EhGXAtBrCvMyQ8CaR/EMH0TBf8ry1VwLx
Z5/V4VxY2NUcf3oWi8Ekw1HgksKbBMDtBjosReTGTjLFP9YMcXabwdgfsTip1kqX
4XynBaX6LxDjMaBJPONFtSXcr+MiBJbqlv6uVB27IdsAUOm6emXq3v9J5U3XLJCR
rwBHq351d2wXJ6+tOO/Kyn4wF3rP7esc3vNdO2hmPT6lwSg9iOT3khdG6HtU7xO2
ie8MNn56Kc/VaYP6nrp/r2791WeoLoBM4S4X1E+h+s0UIWVwOaVK0ElayLR+gt7+
IFBXgvWWPvawtc5QoS5/KA2Y9Tp6GsaRN0jNJZiyWBMm0A/rFsIErjexov8x1r3P
Nv/c0U/7o+YNToylEAqEAeY7TxVqOAqLgrzAXyNgZD0x90RMQxKp1q00JK2jJ0hT
FAxxfHxJzrWu5gDupn0Lg/Ev3rgC2r7uEcLYhNnOTfxNQZjg/Rgt6SG8FeEbTcwi
TI4ZtmiMATwnkya1nTRd01dGr1Q/03aye/p2FkxiKzgoTCSRnqSmKvEwOPNaTCMD
R+/gI3Qo28YjN9wDcIS7IKAywB/aMK+HMJrgvOelkNGpyfYuuLqV1+HA8ULkQU23
66CYoigdKQx7/+ebROtJ+wFTugYGPbOlD3ucKcQUDBW3UzNTxIkHrzvTd5Xty5wh
4L1vUps2L0BFnewVVYE+ZWqHDcIk7EAeJm4VY9q3qTkLMsEGJoV1v7fk4fv8z20l
higcJ/fQMJmCshNz+ttnFzHVN0ErIcYv1MIXjnrNJEXEwL/pYg7PhhJYYw8LXact
5iirESLLhNRGQJgg+l/WaiXY7RW31eW1gUSqCIyJK/XZgYy1lGwvKvJXImKkmoL9
rz7RRn7TAkVh6+874GJUspxnsW7xAdc6xejyKU85/I7sf3gn0f9QEhzZBxiZFtKs
9fLiBYHUgk/2m0qtoMkHb+tLXqlM4w+MYjCMeEolqIirwkznJpK+pDyTWdOGg9nj
2M0l9e4rV4uHGUkmTpp9YLcLgd5vj3Kf4FWKJBCYYFkCPxz09ETskGhNRHhQ//YD
PIQwbLLzcpBw+A3PsTTpkIjpU7bEy2aXFSUasC1VFA7KkoOcH2ct/fsvkAbEtSSN
ppqgGE10feq0hcU/JzJVObgsnqpN46cIE/gVhKukzZQj9oetCqgiIwag0DJofU5F
akSKPghdqHZk6ziruQRwOZX0n5TAFNvHU2NsRf571DTQvsiTM8pKhTw6jPnx9fIG
XFAHM1fyAE92JaUlRhLUuc+FKO1Or7uwRmqXOk14zlLSwNQ8C27IsYaJbmxORDR2
5WihzilwCJzA+12DwW8gQ1bgOEC8QJAzxxoPiqZXhWx9ArPXHmT4jNrW+b3Zy84Q
M6bOfsVIWM+3TB2C1Emwfj8Fm2phJEqlmp1dgH2Bib+qs7qol7Hs9S8lEDCf00T5
ikMQhFb85DyDd0nmtwwmWUoqq5WEfqD00Kgo/XLvjF1c0rC9xMQ731Pxr/GZAzO+
uoptfu2eNTEfVmK07D7prv7aTGhNsG6w2Z/iJLi8fMRbB7Yz3DWk+Yf0GX4z4Tit
mbBmcTu4bw234xVVhxkjWBmvER45teDjhn1l8ZX3sITiXMoFqNbWwdUFUBeoTRnR
y5Fiu3jooJ0fAoqj8sPFQikIjDhc8d36BUDncltBbfHXkn+Aby1SUMn9IHeymdfk
3O5faxYzW/MC+Q2G8ER5T9j1LCKNnmDGI5BhuzKVg7ymNxJYKT53hyOJfcyOOSzZ
ZlL+uToD9YPBHlKYcA0FalMYcORGfh/05U1RIuRXBbxze0euptJ0L1rkxkO2Y20K
/ke+JwPUlFzL08bwORcNjTF735OKZerEUmKY1qLkCj8FwISp50/IBKxm6WryUPID
C2Jc3ebGkmzvWcvx+9E8dtA7pY/4IWomFw5Djrq87GXweKuJBgLkxZbZ3QGYhc8h
fHa4+b06DumoUMGd5Cryi3Ylb0BpGC2kACXbehI52jom1AAZVE4BF9HgBvBFjvah
SXe+MM/IWsuNIgoXLkzK2FUjvpA2jRZrf5APQSw35cWFSYu7Hfh2Pb+zG1iGNo0j
FzpZB4CB6czjQ6L50JO4o9yReFnYEF+4eBLG2nDxp13Hw1QfleVkCBliyj4oNA3w
/k+XXUDo3tZLXSlg5dmwcW2r9Tl4vWBpz2SZf2P2tyxlof1pweLW3DTrPO07YBDA
E3QguDjg4wh5SGlJpyhpnOJS8sfpWxTaBpM9+epuoTGhBepynPt+0jQxdmMqXrXO
LVMb4oA/JpSKoD6kPpLoyBz45ZwJ6GtqgEBTdNCTT2gZ5oxMsnIuM8vQpovPIdgE
6aUgwAZ0EoUCNcZ+6B3t7urPVsy/tuO2yjsflDE9GZXAd5gqCrsyLIucrSDnUy5W
cnf0Ue9BVEH2cWQ8h8XFL1Yt0aHDoGYjOjmmbIeZn2nj8YcO0p+MVVBzFL7Qvyg0
jjkXwHRSoJEGfRNmLJiyFnFMNDyuLhk0MiaVdWMDjMAsYZjMFpobI2MwmJY6TFzh
iPnn32os8ynYZGazF27VdaCFXgqBB20ECiKOY8y9Gf8kP3j70UXFQRYK59BLG46D
KJAg/FrDKdgeUhlmtiSfULfelC3sYsB5j7iyPQ850OZ2/IsC6VZ6KFBNwp/Z7jGs
yqsaqWR0opB+An6uul0Tko2cleL1cXo12FBLRedT8TrfUv3pPHg40PYCl8XEG+uN
hFzyyKvarhsINLP6fHyoOFjpx1hqAuWcdD3UKN1JBDguy5+ZcIO1fQXhpnGRcve0
56R2kyb0e1BrQ7mtqaYl73RJDVfJsKFhOOB64cxaH/YJ3lbjSYuJBIi76owORyCH
0QG71NI+Jm3/2P+XGP9iZa9qt6CX41S/Mvu/GKzRaKqg99p+C9HhN+y5BYi/36GS
QxOEytF4sQj+ejLQ0y1RL3vyazmmedwNGCwdR5bH3I0HFBNxe+TIyUoL7kWRRVh8
R5DrZSP4ju7WHetOXNmPi1v5sSKIg1son4389QDsaY/VxtXtKYaeKqEX7hk3NWMp
ldd3/w9lYrxle+8AtxGb89NKsfyn6OIHpYJKk/YKwPB30j7TPa80yO8ijFvPra40
05GyEFU/6J82z6eQ5As4JV5a3eti1Qk6us6BXwx7jt5skxMt+/hhKYB5eOwE0N6t
4Q9ruQZgeX+uuCrpEMtwMkW0aoDcjjy+kzdU4TjeVYIUlKvdryemWUaagLqr7VqB
GLvT/XlTMXyCSJTLW3pxpCxXQEwE0aa4wvVXYSmKjs98Dz9wGBVHD3SeAYP7VeNN
P5w90+JlNE6td2+1GuCZTaOtsI8Ct8gcJ5KBrrYI3dyFO1h0CqOoWPnwfDeIX8lJ
SZdvLD9OJUoAqhu4RR1KAyZc8yYNACIK/85ZuiV5Ym3/W66WtbzfNw1s0rFg1HEX
OzdEl7ZMxygCrbAF6mEPQ+yGiwl6ndYyONs07OkedqgA11vhIyr4r13VUw9QxRjw
x8qTxuTu3LOI3Y/oQhRMJgdfcPRmrG+BlUDQQ6LoM3brKft6LgwpGX9FMlrc4B/A
QDNS0YVaLO+d+s2fSSMWmtM5itMYBFKhRRa7cPwhkedPxJts7SwhcnqUq39NTtoH
uy47ZHJJY6Kz8DNR8tcOR2h9t+ZbXVXhEQCw/e1jH3KMgwKmafp0dF6fScNe3fYE
C+9+sgjnVOTYv/yfbsw3Q19WYPiiiG0y0XDKY+S1cgG91fGbF5SfwFNhD6y33cfi
lMKoX9ejzobiyWfZdqnNANFKr0SgNXGpBX7GHVNXL38bWodUL4+bN5fJ5sP67Dh2
2Th3ZXSChSl+HoV/wMWeEwe8aOyAn7nC29EqnMFb+JhV2GDO13h0HUGR6sERFlge
n/wbJF64JIouB6vm8oa8AXFEa0K0Z4D5d9JXpQz1ZtYBQz+/w974emhfqUR9s3W7
lRmBpoDeFPXDT3MuNarcGXNjmKPzy2wvgz7yzQoAIwkfNNOnuOdVdkWmbTJOA96q
e7oqKfx3/op/tq20+X4ORmyFq2DAac2n3cK5lkzjB5n2ThyFB2LQ8PB5D3DkT0fV
p9vuvRMd74tni8czaKGDygRzmnKPWpWtEz0wGVzkuRJvOQMe7XqXQqAjJWJm/59C
BJaGH8I6yh5iIMCozst5lIErVwjE4xpiq5chfzpbmArElfYiuNXLqltDYXx89lBR
LSJ6aB08u6zSuUeosTO+565mo+rfVAEYGqVrtVru0X/K7NXjZynG8vKMANupSkvj
Q2+9FPnMk6trIDO2xKMLqV4GPcDAol51+ZXWqQR13zvHnDgJCQ68hFOswwbVOfvX
LTJF+Evmc3gEZgjWw63jBeyEb+57Bj5jyC46bS1ol6JBabk2xTS2D7+YYiNIMX2f
ve8DWquaPrjhLkl32K3dbgojd+TJr+abGkp17r6UHPr4eP2LtvNymvKwIIKyeo1P
INYt5po1prrbSiZOUZN0gi2HQTBba/ui3/nEFzgYAYxNkybKtKGrDcCFPlaK7F5M
OUkUS+5PWHWu5gUtyz3HungmKGP+D+Nx1ihE3hjcsBncLIagIocs6z+bje8wqJkJ
Vl6XduARdPlm+7en633m/Pfwl1LIk1z5ZKXDMWf0aP9fX9swfqSroWIOqGQHkHvJ
QIxKgDqXuvrA+H6fxEuHFwZd/hm8/btPaquPU3yK4xG4xD0Al+tSiMqemXgCqvqb
zIqgy96odTJmpVT9bAnBYJ/mcEmQXCNN+CV1/6+4quHrgGrKRsIdluPx0VDp6m/e
sO9VxyiJOWQcweeFFdeAT1D6awRscO+YW3YTnqizrSS75UyK25QYPiFLVF9OTF37
4+gF83bq7ltEjCEpvM6BpoSU1SjzGri45kh0c++yuNnh/Co3x+M1q1NkCKy0Z7J2
a3efKqdhelmWqeHhF7kIdQ9lDAmrMZhZLwagqkIZ3hVSF7CSxRvCPpD3V26/qEcp
BOse5ZEwKOjSM3CgWOOEj8XSo7SOhXUW8YkB2YcV81i91HTR3h8GBvjfgpVFay08
h91ndlv7p42IKYMdxMdcCJA4P6Hn2iF9z7W1gOi6iYA6xACQM0G7j0aywfdQa4cm
VNQ3ht4nbZPDHnhhhdrqtltLiCh0FOAoiPDpSlagFXqMV8ryy8z6zy3BSkRj0wru
Au90ZPyUwqgX04Q9q4st3hP5BfhZodUGoAHVHSqjbnk9sX7PYfzUCst5FaDWwDby
Q1ecEVumX9azh9mLT51XhBansZ184lbRjCcfyrGPggUcMvjEGdtx1bc8uxjaFMR/
B9RwJVsApcfQRZST4LKfN+akX+CYauOhawWipQ036Rw9hf2vXWife9PZEvl0OJg/
qXLWpfDqWFXHF/xxlSKDdDqtg3f3D90KqgPhm0cOWMtJJp7gKRppckN6SAjA0T01
AnYB4U5+gKpabuDGrzW0BYvWLQY6mc3k9t3K7YMRY/bK533oyArXjFEvxXanIIsb
3gk9e4oKoY7UDp9QxX3Wyo6fYcUPMQIfkSuQdd/t7t+i2rumfDOTvIMJDmQCUz0I
6TBay4e59KspbNvEmCknraUt1eLSNskxGqiNrIEbxZ/FXizWg6JytX8X1G3T5Q9g
tNIulrZ9YUj/bqjlr5USSoJf0F4NytWDHwgvrRNzw3c16ulPdBAUQELdA7ppxxQM
Vmw3svfpNBUQ7oPbpIh1KSTY+coz1TlzB035mnU4UaarJVL/35wgNNjcJNKOH4mE
iXwwWS0fj3zzvgwwrRUBclNVM966GMTOQ1ywMgZGsmOaLtwZRwHYH+DkVvdM/SsO
t11CkGKXHC9HkFMhOfePSAeHfUmN8Adn4OMu1OmmwByvwnEyZxC/GOdBY0mCRuuv
J3ec/QW9YCZ5L1cPrixSYuMyBXkD2zdCCKSwW7QO8qDMPOeQ1N9+jYLSB9sPPcuq
+kfGUH+oMDl46D/ovB3hIzhoCdOYIGoBp2IFF7ae/bE3UQcFbxNAeZZ0IGWjdUD6
WXm+qoFegUbc/onWNetv8LhQtqRK1c3NS47ROjrqiUtaK4YoZwfYixdWO62/1JD4
OYmjW9eDWAmtYO2MNpOy6h7Rgv5oWvHTH+6OZ763zzTryj0JfE86xJ4dznEo5FB5
0ETQvnLFPYoNtVJmkPhnm6mmklQQSBD5I80ZGi6msRjwHowL4eYv001JH3Mp6Y4k
tY4oQOy1TB41pTD0fTTeE/7BbghDFZ747wo7fAQDW2eqhJ3VXQDY3Z/DQfDSURbH
VF7oWO1/EvlKB+0RjaWukpZh0TBWbP00f1xVydPQrO5CxIn+mZkfvmqcxViRACBd
aL+nRmM2tlSAC4xphjtyuFB8/jEIUZxF5Rm5Bm+gSfqldZiKRIpBeSE2gElI8PEr
vmUOlC0wpYTBLU0oMMEOkBPXHsizvXxeVxNao5sYuM8HJ6Z4+ONgjiLAS698J57b
Mr2WqJZzmrXGWO5sibRzyviaUZoXzQvkgyexS7gvG/JWYJ1bu2uoqoWLY3oN5d9G
7L9OBh3Dvy6pPoDER4C2/43wILWPqpo3n3YfjsodB4FADp8LRlhUJ8x5OK4BfnuD
K69+TSbAxLzATwB+euSvC2u2PHZFg+G026BCnkICvsIqzw28gdjHOMis6JIr8qLI
DRKefs9ayRHjN9Hc2VEUmcYf7Vccve2XgQf6+NyMS/MH5KoO6/VltjLMelcMj1A3
/M+1ttW/DCEyKmmxZJLMRSqEf+7Q1x/hPwete/LAFohZHGjbHFPNb0DtF7wbhcU3
/b6mdlLACg56ELrbL6Ea0cudCrXP/33hJw7j+PKZiS1Pu02g7lAoi1l+Yh2SlZ4z
YBCcrQjwjCQSHpY7/2eljjZbKiiQLHxVQkq+z09KFtzORSiy6pjFmpfDfSgVoo5Z
0PNh1kiqVG51vlffhufp69KJC/+ueUVdRK7uijWPrqwRqL/DYS4CyXfflY2rSWuU
AekD7/kGwkDpYCY5B618YixJ0ufjpBNxNg4V33SJOD+3lhbgYl838xlFBw+KpVak
7tT5fHiBo2WjZ3kTG2KmXVhYKu5Rl5pi+l5ErW9Q+fsKnRQCOchDeWu3EQKKpSJo
Y4As74sc6UHoYcfhCuznBsxrTACrvyiwogakqi6sHTFlOHiPW4CSWY+ySQk7QIvP
B787eF6nfoq9kn64LcLlKgixWvmgJQfvlttlDfSpGX3g3s1A9KKq6TcKS4MgStgN
uBWMVDeW+2iY5hDOQpxPYBPfvsaWXXUlOYVrN6uLN5AAJXW172wAyFLcZSu58UO8
GkE4XsPu28lP/8K42IOIF0rLGhzR4JOaFEGfXluizrH04R1KkPfouU8dRPUuzjzd
N5aXx3hLZaeLnSYJkzGRN701vEVn2WwhoYARNxpmkOI3sVsGvTsn9ZK2eIUJ2swC
e9qD6rAjh32LCaAv2ZGEfU25MZHQ6MFLTPTuHF9bnFX7p9WueJtZmAx7l/4gNq6e
OovkKAFlPHWzc/7bC5h1K4jMC/WCd3vxhJ1lODowbKOvaTs6quQ573M/fQNENuvN
Zuv8f8Jk9Y04mIG1g8EIkF12VD9JVsBjfzRBbY1RH9jM2lrveS60P4p6VFIoqyoV
VkNiqghwFdgdBqo9k1gv7mcsyX4fktR/s1z9AhYSQIKSGjweYrrJdGysV7vlHvtd
aCuYqFKybjV8UypKbo2qtTC5VLyhngcI7yAqCa6sj0qObPVoc81fHUgEh2uk0cfl
lHHWVDJ1zvJ3UmjTbvqsncjK+GT6q3dj4Jf6k7dH0c90ZO0zK0OLvHp08oDMtYF+
nQryL7Y69oivAdIRP95vBdWwK0SBe9qf1xpCL62IcEgFcKhLmPIPxi7o78N/07HX
kmGJ3Id7JvBKT5MC9KSRJAJhL7kuGDT12CiY/R7ROSos3Bb+2deruT0EqTIlaBYb
ClxIurBB7NNY3ux4KQucwRPs4epGH2EwEPeF9kE0CX+C4SnaadOPOGSpCRocQfd+
d5dWGJTxQjH+rtfy7jajL1acEjSd1XaGp/uUdT7o1gFA28UGmHnUU3vtffepSq92
8cu1xdu+PKu3L4xjyx2Mt7eHL/It2oha5wDVb+lOiB30v+kbRo3qfrl8kYAp5TPz
717KY+S8UqtF2a541VjlDGlCPb4QhKcbKxCOcRsqhRyWvFWeY2LaSiL130B8hfC7
8NFPPQ4ucytfDBuPgSxVSC2qfV6Z4dyOAexA1WazopQmJTKomPaKBav9KJO3t2Zw
Gr9+JaAHUM2oYyu6nexcQx14E6Y8v1DLK2jAleXZeP5kBSM7feGvf0TkZuqHMqEA
ubMXLYcZUWsvKQFoU2jUzttvup6yEoesET4tLBhO5pSXmOkaSQAvRxisyZ5NOIW8
CMFGtwBh211jvXLlVEWCEm7a8LtIiPPqUOiDTZhvgnq6p+1yxo/haToRsDL8Alc1
D5NHJFFQT14C0N2oHKK2shVVB3/bYAOXDZXXstMSTWrgeem+IW7qmUSFuekvK4zs
gYWZcC8D/ex0bUJi54NkSUbi2NeGBvCDREdtg2zgzM+O2RRQAsRMQXTrf+Jhof4N
E9E386jtY2efd1nEDiZ20feKIB6gZNGFqAnq9ZdkJRNMsR94n8DjOStkSk6uOxs5
67+jRjx+qURe7QVCI84mFkr6U0oHMTDOX0uhNtMWIIaRsdUDNe5S1/0KwWSVJQSj
/ohFM8+qDuI6FgNIQnHt0VlyQLT1OVWHJ0Ehofw7ZMcWK9B+jedsJXXlrEdM6Rv0
aS0MuFFb2Rjvmzv4UpbxVaIcp1WIQmM1PGkewjMScEcMuLd+eCeBJtvqx39SQAMv
SgqlOcrCUiJVpl9hyeBLQHFSIY/dYFNFxG1hfJkJ9ZX+CLXFu3Gvpdk+22NC1RQJ
UFLQTOQFiCEXpmsuTHk1XmozgV+rAm0miq2GZFy2AG0uYr/vHCsUT1SGoZmu/8ga
skxJIGkpzJKkjc89HcJjewvi3UKrWFfFPHhdKSIC/Xv6vQpgY/XPcCkX36qFHoz/
SKvcHmB76lkR2aYnelfakGupFq38CqUgskTmi24fyUK611z2Do3hQ/F/GiRd28nr
l4clMV+zx1P/TUZi6DvH8ana45P/GvjxzREc/iy+TIpjzOTX/VdWuTPo6cPGcrfO
yvdSS9JcUyJzxYEDvUYN8BM8AKV27+rhLS9fLrmGPutzYWfVZyK7+R1LH4grjZqN
tt0vvU+kMOrW2O4X+1s0qi+7bnMnD8UkZKGoih3vIcZRkxQ0N0VHMvw2gY/+A8bi
ViFoBZH8aI9gSgyOtftjR1x548UvX6c73YNssYwnc3tFWggx8eW1Vz5t7UAoAcmv
VcV+eIqg6QKXxuZGT14rE7pcYM+m7dl1xsxCvXd6NSXF2QxAcxNucqMGVp4DT2Lc
f4TFAOHT5ZrRzBnzstPte5ggpwGBKvslir3DJL4U5HZ4yjmQJixxZZm+nAsFf5LP
x6zdpq2J/4X3GFPJ1rtHw9eLyiH1tZ3edwz4slwYLOuMcmeu7oEd/XPXIDLDB2lW
utQQWTyLhr/90gTdq+otTGuqizafLwODegRBY2AvYl4QXu3bDHtghSMVdUnUqo3f
W9/pdY8YIrTN0s3u6mrQqCJS9tcbpqYYNWU3NCx9ZmDIWsF77aSakboYE/zhpcWV
YPQcemrIcFCK3fBM3EslkQ9CUr3uuWQIRYzqQh0m2nw2eS7pJebwOZLaboNhNIfW
xhDmCzs46Q3Sy8xCoOcEV66/NIg9R5gM4xGSUdFl5qtX0lHWH1/BmLW4bDVxTJ2L
55zY4z2WzY5dVvOddxbeSHofyjKWyhlo+JnLivfMR+QdMcdoOIsnoA37tpxLA3Ph
gvHSQ4HmPhrNCM2Jgf/xfoUOf0QB3f2l69E92qpqV/6T9cVZyL5bBNie30zLPXkh
WQCpUadwu6vqD+vobq/a83Jw1OWEN+BWGZtJCm2/iJuShQbqfAkYaP3ieV52wiDu
tr0U+hc4ySNsZ1UxzsRYab9D273F6mVyYx3y0MLZA8h88ZohjJBEOQDe0uc3UfrP
hbD92cpdsfxoGj1atAhI8WObPEYbk4bFpSBHpqklmV6u8dU3BPOkv7HbyDzF0zBD
NxXaccsael1dkugrovPOHz+Jvr15rn7lxKmwZfid2rNFU6OTf5k5Hn92Vn8LRfrt
y3XKJEIZvbs0u/ciCsjkkKshdZjTqhifXlkGvZmUqiY+Dh9hzckOfVxykpaUnua7
o9dOPUaKCejcqKb68JRdGDXzzjrg0C2eAaReuQbsYDmg0Vj3scepzbMNTR1cvEpy
L/I/nTPNFKf1neL5c3XMzVNEnDQsDpq1yHa/UIgKhTBudud+yzC6ay4rcMhAejPj
DUraGy4LDtPjzfWPaY+OCzq3FmQi9S2SYELYomRh/lLBRj+y70bj/W6xUT0P6uCT
OK3SQWaa+1zz+y8O3/QZuuB1LmwAcTn3p393v8Oh+yFI3Z/oACxa6excf3QinYLK
JqdtFcNiseYBd6DbMGaSXh7tCcUypHBkvEEvkXxcmrVgRzjQc1xoeLhVlKx3kzjc
y/4JPIVin9kipjvpfF+4LhR18Fo6UFThuK4BmbZ/gfSFNhDSGHPiGz2A395hYBef
TQfPpHyW0X5TH+ukk8Z/Hu8WX5KnACII3iP63J2nV9UJMQjJPnuXiMJ+QRlza5QU
RVVY40rYMgyBJaNC60ZH1HyrlGrsAj/tD3Kpo28cJirEGRtio1Jf3qh78TSIU7kn
yLy/bnBEUP6A5mObx6mdcPV2lNdZIVpmiEsA/lkyXSoKE6DEPoZtJXpfCilJLv3W
01lqSI1YqAS5axtMDS/34fW0Pv+plwEbnm+ViCjgR3rd/CjQoI0HlK3ZVfyxTU84
KHtl+OvbipeFfkgnCrtkL6xdTjt5dxZDF6a36wzfJwa2vlGNpem6eLyhz5z92dUE
Gqb8izNdntdrPF3q3itqxUk/OwimRMuTkdBZyk/eTTHRTnSpmCA5bsV7DuF4tJq2
14dhfSbGwSBxPWwnqmh9+e16jYWl+I5L98b4l65z3UVzGyMGHjjjruqSsO/p+vUb
Xv3dTFd3UdU4v1+l+mwf8B3zEfw6yKg/L8jFBGb+9jRtkFRDdbt6PoXQnvbfPCid
HarJGpa1/6hh8UARvYCgCLFRK36Q/XPWZ4mFLw4HZdoW7XCwjv8NqpxKgSnP0GK9
3i6EOOSPdApfCtWmK57jveUyL/t06FFTWiomfnKKRGU8SmE2AEFHC+ahG000vUJL
cwObZYe9sIX/bZGyOz0jlHUHvTSgHIJ7kRujY+tmCTM7VsI4+ksCQIeoisB4UvB7
u58dWfnEmRVZENwESEsS5QGp429cGlcJkbYJVbedho5+t9+9+X+JFvxHIqM5RTJG
QeT6nzGw7HQJtRypt3T2JacsqHQwffn/jscbd0fQfKdf+FiijZTq9liKWQWZdIEM
Ui7l25Ts2gF/s6Evyylrgiaq1GQDabHlVD3XzXr/BXAXHXXv9xo6gWmspmDalkWv
Iu6A2fDLs+iuwTT7lX2aQ/S9jjicz3YIy6XILIxWiQ6ikZzyY5gEZ1h+ZpESYxAE
qcKfr/n90jQtImemFcISESM+Jv77GBaHG+zPX1+sxr5S3r8UmRyspG0GyMK0vWa1
ZB2iIxDhsu9Vc49sgCTre6g50aBIrEcuDmpLdI0Myozeye2DmDy1xIm3uWpNZzej
jh1gPF91VCa+2JZdicwMcG/bP2/cNsPaFtYue+6Iw47vU3DPQWrDb+dwJO+eXMd3
ljbLoGPNx6LXFaaOnBjDDM3hFLqdaBOOtp8XOry316EK0RnO8CfRDQtSV4dbTz3j
JhgTWh68BS2KyhvyOZI9S0yuoJLDejZnPM1LYnCbJRWXPt78+NV40p5wD8+01cDY
1zvtbdGyhX2qEqMbwYFDm34Au87XPz8BM/dYGqhmf5xTGgjKZi8gOui/eW6is96m
+++snzIvhWHrEb28gc/Hum1aLAhi2WTam4AIp0SAlX+Foj/pp1kvHOQ5ENk4VfVO
fJArTRpcU8dtmoIRClYmsNuV9ymqhpZ3xgncuEwTzunUP819HQR0uJE6HnBpJsPo
vQtZCWRsTcvQAnDJy3hIrqboPdBmCpvY9MchD4LHpGIWV2oaCi7qwAcusYLKVIew
7FoMtArC3qNH8A3fSGutHCXiXcMyy5vwgxqsqvFAa5EcKxiIAXbwmt6mfpqKoV83
ZXRRGfddB1O8fj257H3LH48tExc6ctnDEet6VDrMoETor3915fKVlhUZju76GPyz
r65kYq68olHYDqGzHfscF3nKUZkWCJ1+vkqjqgcu+J8yxg8QZPrEiwDvvW31GQxE
qOsE/iEVaJYt9WY4ottztrqOKJEuDaagWXsh0Sc1FezR0P1bpFPkpbn6mSpvyc9/
Lht4X/R7H6tFRlFR5EZBQGAiRoUurc6eMrpLSVvxNzlGQcaVATvbtVeKvZAHt3le
NHlAM6qnz3hajr0h4i7mfuICSECbsXcTLpNAZStXtr9PvtjzRKLeSx9YHQZSqnf1
hrtefVFkCGh3twx9dd1+s2wm2TCF99GIm3YthhpaWf3jUgfmNpFhFTgpCWl6Aiom
dxfVo8yPpqL+Mr2rlhd2M4HoRGpY3uQydvqWQx1v16Ww6GU7L6xQy/fVYOGh/cQ9
LAWbhxXm8x2o7//omIeGWKignXhDSrML8bSJPIc9YL+AfRd+5jrFSEFars4t9vWC
CifKmEfhkqcewaf+saF3fh6SQtF84M4VvXvXpki2PhPTq+vT27pitPl1B9XqjQ1b
v1wlMKCtAyWbORKljntTPr5msWg6qbhhflkXVfV+TlzPOwRCC+q6gpbDUH4BCmZQ
cQkUo5GRHr1CNqFe7H/6DBsZrWtyQjkc0Xqa/zZnC0Z2tTahjm9RQmqwZWJoay7a
0HKVEz/UtGqCWyD/TgFkHWOkbXNWQuoEANxFUbwyx/2uPHW0Y2gZwY9FFVL0FbFe
LDF6XcqrZcLXYBCMrLxPBjXwPQsrbKUoDcFOkZag7XzBnw3AQ5IcxGQG2SkQQn2o
YJuANOXub8yrUpxmphSr3No9Qo5bhTDWAhKdndhYhPeCBsyKQ5iIkQenUPeEb/ff
PGVP7FciQajv/l0jKR80za0scJZt9bNL8rNhR4VozXmXJvz8Eo/GpxyRiiEdqfsv
TugKYcaQFRKG6vPv9ig5IO1eHbx58MG9CWbMuc+BwWP/7pQa8VCXDXOpswZJqKhZ
/PaUAXGHy5SiCN7YMKsR5cFJzgUM7oLSDtBqVvd2dUiT8UpPYDOFQsu9WEjYqFOR
hQ3F0YFHt2hKf0lH7wg/GeHrK2ndD803l/KaO14HBXvbIWAiJ3OuumW5RVtU7ZoR
ORRoBGT6MPHyQcmM2h/3o2wfOLb8lyq7mXZa3WEUJxQEG99Gc2lrboq3AuxYWRX1
N90lZ11E0bV42VY6idISu+gOk78QPBFa4Q6kverpc/rh94XkGMhxe89c3+8rCT/9
UJJp9Qe7gxoscMI10J1eTqUj3mQQvfwC7NBF4nHc9Cx3+lftcaZ6CSmv/S2nO+wm
HXbmF8KZmpRlpSmkanrf4JoRR15bhKO00XbZpBaBH6PvREJshWNj6HcjccnMjC/z
YUoCVvVjUrueBOYSWp24z6MDE+u7eigp2uvXdecBMhLbRjNSS6s57N8Pf19sWN4h
piVz0/luXhGVVXovp6uAgFyHwIsJ0b+l/8IHwmlVwZX2408pMUD0h7UTTRx2FqiG
2wAju8DVDZbTU2szbcCq+l6/XFz4SOwk+Inx7FmKAY6ATsoE0DI17r4AT7txDhy4
kPf7r2fnErV8QN+fyUkxL317FSWiSPbzniK59yAo7b6o9kfy+iqnQT4SCNTj9st8
rkgNzZ3k7jwqVs6DBOZqmaQA1vVZm6x6C/HxiwcBrEKPgEpjS9RF6oMXrrrKWvXy
hG2AQfxdQJ3J2STbn6ChaH/wtaauVZ9O6y+tDBkvYaJOZtLsDiQPCxHBIhrHimaG
Fe4w3t2sQDljY8rUtvNU4Jz48ZlWjP8EfDwJkNyuTbkRtrptCIHdTYvlD2C9FCZ/
Ffgg4ZW+GnQARBt40XKcjvGZetcXPsKcZgYr8hscM/ZwIyB9Q012QGT0TUUr7vBn
Rj1+fLAUmS/lMksVh2tSidAD+31xeS0/B3UCuoLeIrnPDwmIha7bMwqqnF+Oj9cY
UyVLhisPfrBTsCu3fCxHgNScTfXT9BQWTQF9S1dmMk1Pjn8b+z2ytylwBAsgQXw9
EXTS9hO+s2GKltd8qddBGYYrer8fgTFM+rnhTFxj54ZpBy7BgCP1gNgWn7ywBQBy
H6syb1jhgll2TduTQ8A8YEtYSZp9WGxmChgkq+s57ZD3lN+hA+QhdSDFsXqpIeOs
H+hFZ69excyDGoAo9alIxw1bydoA+ujm+ByFWKsllfNLZQSQWkvenQQkqxGOFD9I
T1U+7sFMiXCRZIljteLt0h02dUzZN8gO4FismLhAHHMWIwLY/rhE8GoSeWpmN6GC
Jh9XUkGWv2lEBpVwAIrtA/+opCNf9xaeIX+9Bea66tdY96aOoIA+qjf+zxXel0+e
K5/EQlcG48wbigb47BlK9ZO8hlDATioFi+9lR3ajfvzSJXBY5ZFaxdQ9QCAwLD8E
LsWVgNibS2I+UA+VeIfxE85OIjSzLYnQGSFEsLohNneewgublrKRr8xgudLBC71D
l50CUPzklHlx25KfFUK2s2A+Xkr3ZlW/anXPPailUMuW9WlHBfyRtkxtlO6UoGH2
AL73vh2hsaU70H+nkgqGdAHnyhUuvM6nJOIGVXCKbPV8kaZd8znjFQkHCXFGOtop
pO0wT5Vor++SYtdYdzUO+/+4ZsPl8LvvI6K+WjVLMwL0JA+BC/RW7iTCcDLjahg6
PjTeom5H5dntjAosdHdRGJ33Ki5a0ZxHWR2HzZ+UbMXPFsmwSqwKuc9pVR/qVvPz
8IvYoRb+fpEq9EyEUs9y3nm8AHnZZGRsqiFJMijZ7xVwIqTmfpII8I2OonLffZpi
E/I9tIghRZvo4n5Y3bN23yaQq/bSHRyiyAMohEPz9lrsnU6vMhon4dxWjbpiUhat
/NLEpDlpIhpKOWOvDZ+7LPVySC9G05bkpjLBs+NP0xSx+0wk58sSK2Xk4CQrZtct
ZWjBOi2HpqlbQhQb1I4XpU1SSF2GvJVNgsdEri5FsJJgMYbL5UIaoypWAItbYKFZ
n01zc8t4Prh3CJgqOSBPNj4HUpCCIoaEYCnj6xbSck0fY15gFB/enAhuO9gDAylp
CYQaIOXbzLN7YL5TdyhOVlapfMN70q/lDhstjBXwnbnkvNhECnJnp3WQMkvHQCqn
OXPb5LtwxVEB54vN4LwGll5MseRPTxhPGArujuA38LGcY/Sk4msyJNeYFBkru2At
d/HEmaeoHDEMeMkD5Za/63DgOKxT0iZoUNrRSNeevA6szjcSEhl+GQ6k72mZOAPd
U6g76F057jN7FoOdwufHIddjTgpvNlL6nli6FukOEUt/hm/0PLtzYD4dHUZqG2UJ
7GsbfwM28/L0J883hRSoIa7L7lOyCs8Kr4wrOOli2bU0ZgFV76RVg07uZxDrfp6f
mLy/igjBd79huOnhvZOEiShEpKvLdMBwJOfoQ9hCrxoHklD0OnRYg8NVdUGXCqJ/
dl/mwNCB2aiwNoUZACmwTDr2AQn4RSt7zaJrwiXH3a/6jl7ZXBGg2qhwmDIxylw1
/xpqWEcsz9T+SkeGakK9MMe3NOOY4eIlFEWugfahRLGDSJ1lzVjPzWen5Z9jkFaX
Wx/e8ZrvQouLu93tMsx2Le9KWG3LED1dVlzz1r7mHSEXSrAfGMguKNjyvhNxQov4
qcxQ51RBQnBUJGX+7fZJDR9xt7zNR0V4KU/toYsxDn9L1IrcawgQjzk9+i961tU7
odg66rwJ7HAByKKEK7uXS8DFk6Q/Y6qpYBlaUuTX89Ejysx9ReDlTJU6a6l5MELf
VO83GAB3HBzPuIFT6mB8pQd/VnVRMlwUR1dX6pb14ynjiCOZTn4BXuiHGSzv/Iez
qHQOfLAXSXNZu4vEDGXhuPnM6d/JbqgWq+WkcO/8zzESSggBb9g+DWJRTYrbSs5E
DiiwX8MCCxLrIJMjXKlJZ9NWTkd2y+JpteTTqVpbJLuAhE/lv6LzNRUp0DEXgi3Q
ZyhM1LQerCJn0uHIzBDmzyzDAbh4XgbrhDWAKI368+lCFXoevXJayT+mPLYVdhvr
QZE+SWX65vCAN9TqHrcZKMEb3blq38VubSavGCW4cFPFngx6OWmA6s9e5ySE2BnB
qBUnaH2L71YECuYK12oe+2ADbXRcR0s95YZXrSKraFYmS18OGC9nKaFpOg76c0pl
Bxj7L5AC8pW0Kl9p6ywfwms4L29YBmKRXV2S6xKvR2AiO9OY/Xm6CPQdJ50W9Iy1
1/xgyro+SOzVaSkL2ow9SvVFwp2nh1gosSpF5R2PEfRTYhcx8cspp0QSbW5OR0Lq
2P5WeTgcf2kPAMJGad1BZxq/wK7G0zMqSFYTJJyalwA3zllcCHYF2NtpUEIGm7jF
gtbi2AyzK0P9+BQI6arVSoMTxuuzp5YiIwJmEfGRjKX1BJWQfSMtgsWYeV4ZbcL0
TvyDVrhLc0aXX9YYne5EjikJTzBj/LDRS0wo2Ih3bmK9GM4j5sGCgIU7iTQFJcJ7
USP0wzO2ky6R79XMBtgAB5qM7tYd5n5CF3oIpvYlO5PiTvykTmhg054GeUH1ciLo
AJPbma7lBr6E0CXgRTLD5gMfbC0Sxy8Eof58Dj/rsLRdJayz/y8hd5u2t6WQQHji
M56S1Wue2Y0I96PqXjKvNstIYwv+S3G+vgStUscl8BsB3IxzybNwQYKGIsgit9vv
LI2L+3LJP/IqpRJ1WqlV914Dl71zAhQjDT7t0JrRpy/r3E5kTPzUDDanrUJjufaH
4XKsKPA8/SJVVC8i1xhZngkTOpwAhf/U2MRo/dbUa/t5f5wfuzArnw2i2ZWzRH9g
9s/Bi648tUXNJv5WwA8DLVM/zW67UsOYXQ5Zla3TyDrdxzO/HOzwu6Ckhwyupfs3
ezLmOacGikBQ1z75wLeEiShagZMCjFnQuPwF9SUVQ0bcKKgbqWonr1oZ0DGzBnII
Au1swhk3FUD1xP7gsELYtLMLYNO/Q9nL3ulEpZ4mQFWxxoczvHLsROxrbRqVbNwJ
AwhF8WuQKuZlGXjtlnPUufNTNl6UmdlXioTYXXsNpXcoWSByewlDd3g3rU6hHRI4
dI1qSKvT3fppf8E+eUBvC5xyZgQ6N2FC3xFNyBAjMNzkephjEsqYsBr0YUeqCcA0
Yb9NMl7kUlUcvKpA9n03bvJlTnfN5Jgo9tC+VwFPduWKcHAfLp7hqPNyhSA8GCaC
EgtZ9ZcpQAYxfCz3dnD4V3AhVCwOeZrf/bCUCUssTbhA6EFe8hS2y25ayk6uRfKA
lEi/HKhIvbmsjg3nLjc2OdYOKnT6dyUkwDoXe+1v4ZJFICPT42d+zZ7vtUIBlOEQ
SxRPkX1EbmVmfmrxJtP5hcn6F+ifrEYgJXXHAeRExhqh3+JLXV6gOmv9cpwUVC2z
8IQMpatbWN1Ptv0Kba7hAsM9ruNXHNOC25+EWvxy3nt5bTT/drFGJVmQAHHhOE0b
gFrpnylQhzCki0ygm0onL9l/Pr3lqf+bp8ywIsXCkWd1n4AKzTBgl2sbg7rqK75+
CHUYNqEY4Dfhnc2LxdEQ5M96vmtPGoMyY9VbzNmfBC7kgv+17eZujP3RFMP5SMvp
HfiHP5ZM+4HEGdBgWhl42SLJn/hogTB6d4RBimUnyzU4E8M++arZ9RN8CKM+QYVQ
PpJ6GW6VJyZLl1/1hPapFfxY+aDI+7yERG8l3zN6yzWb999xBzDK8xm/WI7DpaQB
gQ/h6MZfncQod9MjHRlXslp7oKIUMS5TMC+wf5fPCVfMixE4UpUnn5JfEigWg5ds
7wjsuQWW91zEj4rIvP6FoFtmR/rhBhudmmQUnzeMT+QxG4ldoxUs6cqTar8VNUqw
A1hMytfBoWYIr57UPJlwLvhLB1MBW5vVN3jwv3jYqtpWafATtHQgv7Az0zUTl5rn
dpdjKD22K117PhAXQGZRe6xQdG69D7Y1BqAJ+is9DyCrkn3bT9WEwiUm3+9Y4AKC
NzQ4o1sFaWpzEzls5WvuBeO2VShZXoMG5fOf4SuSjoGbizkNm+SP98ImYSNipR5S
iBwrw7AI15RRm86XEbfP6qaxYxiQtNCBDCsmcJYHuB1DNQNEGmahWBguLOKnh41A
ugDLuQ/OPhxLMn6oc4hiPfeNKx6tTVEYr7LeB7Qjzf24olOOTF+axMHrHf+999Fo
fAabTEEyxeRmpHs0sTK+0UgC+x8haT66srpryeBev/eNPXQo+tBBt00XBdEpqB+A
pcg85hvT2W8rP/Ve0h0lMBflj7R9ME7MuwZqSnPaak72N8oPFSCxr+NAFrDl12Qm
6cNFTnEb0JVpYVQZBE+4i3rq9F3NwP7G23/ItV1+mykusE1vTkfZ9InqtY1I/2JK
+BaydOsn+jJdz4kXFWz9kCkussPJY94YurOHm9x37FAMOLog5e2DnEyJK//lw0gP
Py6YS2UM0zYshhvxtiu5vACMSaYV+MQ/c/xv7+6+4ieu/NiKVoKjc1IGVvCjpmI1
mFwg6cJ+I+V5Z4w6Nek5H8mKRGdCGJv6BH6UhwrvWHQ6nt0kA/FosVF8KbFXYVrc
a6gG9ZWOmRi9Dsz9sOUdIuycxsk62x4VBeazTaKdzpMcY/SE9a5jNASgUebcphqd
EggRe+4ZKwel/ktdhhJzevfmhK9gnoSXHXFEaJRUO3gWlHmXhkwwNOakyhTOYg5r
PZPG5swLjB/CH9wnwGcOI7e7TOo2AJudkxYADkoYKGT0WqjNKXRIyUjbdzj6QzqB
L/THmGP9HL+nBmtQVjWXWCeCou4lhLb4bQocMluNQ/R1r9SQhZKcsfCM3i+8KYBo
lKIKDA+0Xo7aqSMo0WQQqSs0OE4qY/8Das9fOgcy8xI7jiYO2hEIBJSJUvj9cyEt
8DPxmQEv7fBJhY8LFltHXGB4lxG2bBcxFjtGHKIGYWmB5u8AgxhwHJss2lYtNPkv
+i2C++3sNDJ9EaE6gt4HyyPvTA24N+ITjYNr3ARHoYFMb3ROcJ5620plqX61Z1Wo
9zu2SK3mnFEE2StHCBkRDw5bIG3E/RugXV8woUNPnZNxfmVwAtT/5apEynn/60fK
vriQz3y8As3CDHKuA7abZDKWht1jhdY2P6jLzbaE7JFvfZ2S1YozSW4vC4Cz7R//
Gdrn1LauS5+noVWX2YOI50c09wKs1XaQOtA7T+PkTIa1Dmi21oVxEazmJ3/2EGw1
57DSTeB12V6ekMNKuAt81iE6x1jM0EAHsHT7E011GuO81pJipeh/700WgWSINKqr
DlmV3NZXDfJVxcFaeJjR+hGcPj/z0eay4gBaTknuTtBzFtZEVXwLmFF6am/wy3YS
zBMGb/O1FhF2CibzA53GClFQc4OaGxyzrJq7c8tLbJvuEPMoHc7AdBMs+txAafYx
o+y0AR0Jiqp8F+EdkwRyXRi7d5x4BRWEQkAYmPch7PnIYC/iNE769cmg3XEZYxBM
sJIPS8iy6A+8T/Cd3NO6h3uUDz27yn+mw49/L0/ZWzUw+dR1gy3ijBI/txTRJVYD
xkgOP3rFjIry41xHdUw6EUCNBjhWGFvfcrL5m2XM9g5saaifuOW3X0tCIfkpoPeK
s5wwTZgkNiFJ8RMpyxAosUuj8ssQL8xsz3J0z0gJfB8UW6FsOlRu2p8C4ORtV236
dsdGlUDh5Di0gKc8m9JYC5Cj3/2RU68dEqmxIsj+6LkxYjD3X3DUGQmiojsyik9u
0mLlrbv4zAuhv4ZFqUtYfTsXSyjAUsQFbUnnr1ye6Vc14h8p2pPME/+ygIsmlY0O
82EAeBRGJEwaxeyavzsCUyFP+ZHAjS9zEkhV72RIliShG+OoBRjEDW3KfxrKlojD
v6DAJ2UpuWteasMupbaxlScQQuZ13J0SIHBs7PNcl7qpKFptAkEA15CDVzgT9nQI
VRhiRWqO8K7umMjNSmhvkD9uD81otXkp7ZCnMaUOr/Ppld+d/VyF/PncEnVjsEDE
G0rnoGoJjMJ1tdKcWn1uo8lPmMcGWXDv2bWCSGEcGfralRm6UrEYCdxmjoXusBy8
C1A9NvkrkPhaJMwdy7MykvIfku9QWqlGP+M40qaIQFj3tCfOJehXwg90ERscmh2y
UX5z8ru+9fQoJ2v6WHGn13hlYGPGoTmfuIkLlH1CMD/W4OvFO2fNVRbbgTUypExG
u+pcJjSjCU7yyyJ0sqsB46Lzq5XsDZKlPKy8uH9jjmBLrsr8b9Z7sc/mucnMpyov
mhbAtj8JiEeRHg27ZchaY7Mhx1Kg+7rJPSfB1rkGexbeo/1qJsI+i4Yh3vaR8kmy
phZ0gJu9AgrZwNaFRy7XuEpY/PJew6sZlHGmpIAFXgtkQval8pjYTb/FRQJ34ANf
PH1ytUd4/fslfMns6YJQIT6KZu3PLXaOt0eUd9ELn2H1lDQRmMga5rFPviZ6JTN9
tOWj7T2dIUJStc9GErePFv3JIJnI8kWl9ffekwPv80myDx0ApLfNCjrcg04lfsta
KVgnWoMY6xk0pQSdr7G6pJgA6TWDMt3IqbCOqrstdyguCzYGsf5VYQq+sPyRFPPc
kh/A4dvcn6+0qRTeg5KNw5yMrgYmzV1bxNqYaTLIVTtwYbcvZP9xLJ1t1fh57DJC
AoL2RLrVjbJWgkzCF7h+72tJu/MpKlIPwdUXh0ngzGmR3X/QFY8eX8ZHic5si6Km
sjeP1cOf7RN2XDbx/u3vRofA3BkJOLSaei7ZVaMSbiLUQ47LO2PQIlj4Fn1z2kjp
8NdDAmlH8cGgRVE/RCSxWAMU+qzPLQbGYcaBtmeYoUpds/mX+2Ze5ibnJbc/pQl0
ZTMyGFQ6BAixpNO7FrWQfiyt3Oy/wm0V/PcNC9PttUAG/DVJoE6nTe81xOBD3ep2
cSgpEh124o15nZ/aydtN2HqgC8Mxss+Il7a9sWfFNGkS0RxZNDruPeeZA9EEqqHn
jhmqH/hoNOaIQtVf4AIWXPz7cPGmam/sX/qA8FOsEM6ken1sHKQhpm4NkUFwk79L
xPmUOxoa8mmYRo9nU8nKlv0X8/phCXRh9o2LhfqqG0N5Y1KcP9b8jbSD4BtNZMiR
4Hcueu5SdAYFohpd1RTJNA7/uOHJ/tEXuSAjg8efM5FTNQaqwN5sBpNu96jBWnee
aw7YOnPrpCf5VwoBrQqOy+q7SPBZ5dSTPaS4M+GU4WP6layKmtAhMbDjV+Rk/QvI
q2wj1aol7kBMDu5QHyfa3IzO5272drf2Ducx3RHXCQya9Y6HF9j//EI/lAaHqp2e
7OyXeVtsZpHchgBD0ra3MPeWaO3yB2Kbgxgeh2W3jzcovP8QfOtyfqAfvxnjN2Ca
egX4YE20xB0EgPx+jdFVCTQbSFV0uIGHcgnoxVLsfCiBIYOJNan4DvKrxn4CEp2P
8MWK4zLwbAxW8Iw2tJ2LQPFrPMyrIZlwwvDiwuOAvapmOmfDuDwo85NLAKx2AKYk
V+WdUzJDvTHcF8wrXImwmoI+b2NChVOcDLdcOueRT6laY9kaA1aazc8WV7fraR+Q
fDjQUy9QVzF75y4HldIOfIJWufV1SZIVnNLc/KzeGTgzNVWd8gPqDHuADAhNPjOv
/5wscKV6LkwKExYF1En5JaGeAuto6VzRsNbDK8FufLYmyWFlp9ph5hUMrP47bZyj
LGKMjBrUx7teCUERqAB4JjLomZOCb+9C08F4QxLYS2US6mYfpxApKYZ/kbEovjF8
rPSXRIyzXlyC7H6lzHvhqwwI0Gr1JRTmxzn8wWmmHePMdbmclwtCC0CoMfYRz4/k
EjsBSNwfWEcjNkOH7gBd7/IJqEjT7316cVnY0AQmC8LoeMu0FCPcQcjaDNJJHS+v
PlDBm7Q84SRnBsWl9xGAgSc0ZWSTSMb2RYGbixQcj0sveqffWvy0I7S1od0+AerB
Vd/QxZX+tPSCntxiW+aFGc9ZcYwTIY+5+Zp5fuOi/8U2iLPP30hA0IuWYRd+qyAl
vVBKZlMA2nB4ipCQYFcG65P4pR7AAdjVFo3lpXo6PVkRuFaQu+EjHanoPz9O3I81
5wYgRcfHyUDBe6m4e4Yg6wCVsA0ZaudcJoLla5P3cD3OqThl5FU2DfYLGHMBgOj6
3ql961vDZD8Az+Q/NhPfeI0cjSsMe1mBw/uBUW/Rlwsw59oEB/XCnr2jXqe6hhjb
YoG7QMrQnDpbhvaVMq6JXPkJX0+8rPH7lVsbkyYLUqBIYRLZgCItjDU3DGUjRwBa
US2t6bgBq1K11duXyynjnYJnrFo5e6u6FV9sfAkoYsNgHDmcPofpO1QMddkWf22K
ie6atKLyW8wKO+w82gsYHe7E5GQe/ubbSi7OlAJO++dz+l+zek9bpumKJ/fCIqWL
4fTHGWFW7Jpde0RXE/92rF10ZI8N6OKZPJzX6xHn8YrcddHpDhQqvH5U35LYK78q
zrqc8730QEsbimXuymnHJ4jLwOUwYT2F+n3LzRJ8hvP9mQMiP3PZm/20jFzCzwb9
pzt1rLIMRTqXlnf6aY5W+jsEYhQojcWPUPP23S/WT66juzeFr5NGDRtc4YJpTK09
aVK758Y62EYj9hZRZCmON/WO5uE3dWr/OYPoxeoLRFlJRIdgjpFbSVNDShEmm/Gw
Zu2bWiMKieHu8lsNnO0RLytK9vOGTxvfzozC4YK6LQKyL27X9AtkZeWNBo/hOgEG
hmEvLl4UkyZlpqnSR/ab+PMH6FHNW43cBBUQtuI+YFhEc+qnW3uhC5AC+TI+LLDR
K/7aeKB/CyJCRLl2vPNiej8mydyYRXj+Y+t1iA9ENWmAtA6PP0U/O3BBCPVbPErB
/jvhtccH7Nza6dh44BKTXqRiQahsJfUHP/1FrIhYp27PnQJkn4jcJBw0aonNlpv8
Q02w149cdNmrj144mbM+fcwsSPZcMzAmSDuoYqQqlah+czp1OKhu5t9gZhyQ3nSO
SqvaMcM+WLZkAvLA8E98yR6GZqeikkW24B5fVYsvmbDGY3u1Y547PHckYwNZyoMB
oWoHWQUkyRNPpepUmpG6q39Z4egl4EaFWXf11rltSlKC9ZdIEa9vipPh/ESOQkC0
2yB2JuJ3bwRauuMtaqfOfRoZL5HI2BR+ItdBGyyG/xrDRa5Q1M3YXpPA3gMDB/iV
ciYF/x6dbN4BE7J1dsdZK4EeCC9pzYzHQGmgWOEyudbp8yQc4YiiGPeXpKmJldET
CRIXECkbydk8Z8CmzXniKwUl7JB+89Le0Qx8Dox0qnsc0C7BcOgH7fAaEe0HrhWE
28EONVfti44P+O4hagxr0FuNPCCn2UJvmUavSDEUKfCTlMx5DPzSiHiN3Me6dzaA
rl6zTopT9/v3LYUbzhCqpQqARxQalMRuxgDPXbogUNiyIpIo5YFMeTQkQZnPj19f
SRYVx0jC+pg9TiHE+UJAyfEGh/dc+xqzrZqasDg42hqMV0yqbLek3HNX6kQS347F
EUyen6GVj+NEqp6mq+gH8w1Ip9cOf6uRf1E2XlJDlhsmbPZk9kx4SZ7HgTxAq8lU
2dRRHRAh6a7AN2o8R0QS7jBCmO5CWuYNad5r796UBu9QW364PaCJQP6/3XT51T9v
EGNrke9EXCbp0ZsZss2jzVks1azVbK8SKwm76gcYBJnD8DzlqPkGjluKa7WxkKVU
5MnLn99qFCk3ryNcOKoaxD9ywBRQQ12fSI32xCnmrX/nb2i/JmkkBC+tj6sWv6mL
MeKDt6gcplK0dH0w9Ao/bcOr7mY+XHWgZDr09VF7TajRUB8Nj0UKJTEk7vL+CW0k
gLv1P2tzOrXJAupdpWWhqeTFEswA1LCSrWXQm9dSr9QcZTNwTOE7b0+DdAGmewQD
/aMcv7hLV9Aq0xI9PyHhQxDH+gTCHdFIjmB2X7X3SIMSgm9ERCP4fBDIQ65acgoS
rNgjsI2x68i1IwhrWITJMBhsyQQA08OnK1NfalpH6SX47LOm+tBkisDxGjLL6yiR
rtDoymMINIlWUJqxbT/BsR7driZJIowYEtZ8Sp56zqLilGQ1VrA3J0j9RiHq3B60
t03Wnyj/90fmyv7l2Ricl8YCoSsPVES1p/8UJFk8SmVodbagXurFbLPDGTD7nNol
vziViK4KMqO8QTmJmgskbSnLRCy+HPH7eHrZiamqss/u94ODUQVwHlRcRyxA6tLi
/ap295fRowKQuQqEjJGHq+ksUCzdxmw1PBjI+VwMcJbzgrjws/pZq/pMjMgE+pUT
Zae1aPbHhgkKSPw4QQVzjgJqYckS/2WZH7V1rDDFjRG5FoxkBOOdbad96zPIH8Cw
WmH2+23nVjyKCgVjxuDcuGFAdDohyz5zV1WH8iuGZtYJz72LCPyqg8BdFuQYPiuF
X3x1c9NNsj2w8v5PYuzKmcBYAVtDxaZcWSMpjwzwkGqYY7qTP+Z/FxrzK8qvCEw4
tiKPG+RHUhdivJsiOsy1eOHmNhoshr6g4enZWPyPmocz5tt9lW8dymCt0/yPiBCH
V6WmpqV87thwGCybKXTkB5Fk6sKsBjGiEo++BxCvyxJNkeEQ/mB0z7Jvs5b7pzOQ
GmM7rQTmCSQWEJYFeYJ247GQktlkVHf+MhNmQLTy/bGymJGx0dKDFvRVlN0A6Dr4
AX2/hjnCaI5T1//TCAElpmUNYCqLjMurug1kHYm5K52yggt6TNrez1xC9Uy1Qgd5
JRx0TtOxg66LA6iPKEsklFErytC/8mvwGiOpWxHsN4sEvtLUvVC+WUy3OiviRBR2
FFLL8ulr6yuAUPAXOeXzRNKfPM5uKexDdECLQirGuG65uEGHfKgbT5iYmH30L91u
oaQ/0Puv6CFuuYDVQ1Scm0/4szeS0USwZ6T5Juh3AvfY0u8jnbVz+r40vJLqfyFd
FfulEEReyO6FoIHwh1qFNfJvR+2+RINDrJwpJkrn0FN6IrC+17MfyOTxpxGtTAgg
/tsIGY8S/RZ1nZDVtfi5D7IiQcDkohVBUHcmpFv8o9gqTBQmU1bQWhJPQvGAbc7/
WNETGbTf1rAzMT+td1/s8l8Ewevb4LUEP7n8XXjr3tTVwMBhydn+f6Wnz7sqk4y4
UkDA3PQ3TK77eaXRuRpC2eLhZEYe3xl5AwOdGNcLbj2w99NL7EnVOHGFFaqQZYmE
RdXe4FWJYc1Pz5xiBJA73eCDeWstoLd96SyY34R5/i9jwoIetvyimOrHptAa3Hk7
SxDvP/wRoG4JLAPQkEmduKi6VnYxEJ+4N0jemAntUx5JVYcA1jOPZ8uiDVCSdWs9
7VqhTqL4CTnNRMBZ7GhkkazdBuTxzwwjSEpBP5DfObfWfjnG5orH2yN73MaShnDE
XaH9E3n1kHl4uHvOQMdpxjQq7KQhZnOCchRJNAyTHB6O+L8u2zjflTAiFmBmqIeE
gzVoFnlTSt1upWyfaWLM5L/8u4uggetx+RCsvmijwqn/hyuiuCg/7+40uqjz+8mS
CMkJx/BkVUjlZrlOby7KcCjIm3qfZMIQYfQXRaqM3Qp+Wx/OJPO/DhKklkUVogg9
ybiUB1MIbUfGCGPZKEynAAnhFss/eZ8uuCTfBbTy8irVzBzX11R9AGP3C72xZ1O1
F7MZvhx6nsTNr084SsGMgdrhGFQKgNt91f5B4TD6VSrUupIG1xhDG2f4RiVPZ4VT
CCI0Cn2XQlP/LqUkjfLRcaE2Etfa7Wto9Bi/HgaPCc+aa3LjE+lNJPQMM/rfQWbN
KfnPVISruD2k/rzWF2yUgC9+4jDXQ+pu2WedOP7B2GaJUC3xCw+fTesYTr7y2EN0
Reh4b+1+3NZip9D2gXQOuKL7UooJUfOUEoioQ6a4VtS6YW8Uk1sn1OJznyOC5MpU
q8hjHkS3Z5mgbvXnkias4d1zzZOuqtZXghWbY8lIBshabDYRwvFfB8TkmrjhmOSO
nUxjnKp1OiPNKxC4zdGNsmK15Y9e6t3r1CayUAVAtTFiQnWA6xkTjWkuXLZeRJIx
ev88/pksRQjk8f3jvo2ZqSRwy8bPgZ44Gs+miqlkjyc66dtZbAjy8mpjcUxIZpMx
Qnd8F2Q81fr551HjnNOrkSFVE9O6ilGeEIuTmxy96D7uJMUvcrt8C4zQy7ZAUx58
U3SsJ6YWAOC4DJQhI4vpy9zSD0jAvcgYrwVpkfYrypTfEBlmQrXoE/rhpXHMzM/m
4L5Md1mlJxjjkEPv5PcziIHbdBQ51r7PNRm11g4A2+syxLIx6wPqXHDt6xSD+Wv1
wldUjzPbmvgkkRU4NjF60tR+mnQ6aED+QJFiNmNlEnbBHq5+7wVj6S66s1IzMax/
LoZYa3LxCoW88kwTtV3bCXZmoc9Gw+lwcGAvYSteGewF1Y6gK5T+LlRXZrnnpqSV
RbJ/LsZtjZHpw+Miji1bHk9GOQ53JjJJ6XRqsEQanmSr64K+ydoAr322iw+1mA3K
sH0WWOqL1N/ZokKK+t/AuOvPg8IIExsgaUyB48rqKh8z4rBFtRseCoee6gpRJevG
q3+6wmkhaZK3JsqrRUCLxKyiOOJPZ86nnebOKZ1p10ywR8RCx146B+scg6QsuKW9
JxsDPmSjQBH/EHzFtK0cQsGk0efG5keF0TmMONCK7hKyEQ84JoFcoLQeRzZihQ1u
S6/Cb43g9ybDzC++jefM6hPRWthZWavSa8wpaNCNIFBqqYWAmvNoScVdqD9p94w4
bjDB3oyDNdZZHKEoAznUvIhsQnCNa686f43BaxaqHov0IUJq2QoDR2JyIZvDBEwl
8vg6I4G+pUTjimsEQT5zLjp7sZBPtocKcrG8g66ZDZmBdzYasxP4Cr1tnhnsmaA3
8fdwmE3D6P+r6qlkoVPHm7LWMMqc+kHSFQLL06guGFLb0nauSgMbFmQd4TVDZluo
ZZduxaNMQQ4g2zjgAtw04NYy7La1u60yA0lzntRtt44XTOpORCglDfo9vnjjfcoh
4B/ht+m6RUtjK44jCK4yJZ569J5Syuv0MqAlFw+N4HfWI563hIIo9A9IADOffqkC
hovBjSAG655+wV7tBeb0taJc2msNjCePG8KMn8A3OKWhkm5XvZd2YaZZHMob6xKq
H7zDD9+Nz4n1+3DLKWun8zZT5e7emptsweAbepkHbz3P0C7WNPjP2bleMPD3sLzc
L5wiflm3Ht1YOR/79C0w1rwNqz8RrMy9f7llo/LGP9ePE1je5WyiTBA1CPzxRX5o
zRa//Ui2wuHPW6X0r4SeijUm1VWCW43CcuaDsL1CYtY5bIwc6lYbLVQtAD5sHO9V
FIWgokxvyhLolVivp3IJbWEYgcMVSwIxLxEqSK9B0KmRSSkygvxGl+18efaga0dE
qtwSbUHe78GsqrWru0boGFFn6sIWULGNMSTMT6fYJmSa1VuIckLmIJlCQ5X9MtuK
AuSgeZTlx/J/7HX3Vc2URCxR78Z0pWUb6hmZACH5kaR+wxZO6YI7YA2CYG3PKI7S
7uj0cThWJ5kmfpmZuVVBc2QRH+rG/dbF1pjHKavU+X1oLbGF7kInje7/9Bv3yMNE
8+jxfZQaYQ+PVyOjrH4k1p16kNwYXKd2atT+5cM+RpH2JmL4IkihgPylhlILA6Ix
wDY7YlpAltNC6dpKa1zBNbZdGfNo5MgC+q0pSmZnE17eVucRmxavDl/jdhU9EI6o
IT9ZYr66qM2u2/9CXKWwu8kqm0cLh1eA2fyCjD05ps0=
`protect end_protected
