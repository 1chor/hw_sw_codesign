-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KyUCtUFTksNlZqL7R0AXyT7GSo5xujKNECHM99M34a9jfirM+z5u1Xvbi7aXJAawnerZ5WIRqbW/
GkSe1JWXx5CXR7xr3PzCMBYFRFQ9eEA9eJ9Nm9McKuHRWbaT4rj7ZvSF6VI+354LdPvCdokuSJWi
g9+70DPjBQ3Uhi7kPecghL52B38eiUomH+AD5OTzQkbXpOdqAmZLLEOO9n/9IdkiN4BMcUpgrHlN
8wvJyxp+2/1qVSbb1Wu94sde2Hsnwwnp98a5L3i9lLZLhKMWBHKn3nBmGuob/Tbt6yjxiTSvjFff
gLHJPTPswoMDgNuyTNEjZwo/gPerSEP2G/nV5g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24384)
`protect data_block
29RwTRM78or93g34suqRmtbq8zPgB/sm0jAlUKX0iug7e4OnSR9Euw7e2LQrraVF4AJmdX4UJUc/
tRABnGxTH8+SdZF26p3U6SvX3FoS1ddhAYr5VOGG/QSgZhaT/9FmdHn4MPaU0IfH6+93F/mpVemU
LIy0TgrGCyKJPZ2kBWZElj791HKp03u/sl9OBfuUJVIxODoHDCRG/hDVsD+uev5B2nrb93G8xUna
9B0+bVCtPuCosDQOBQTNv4Qm0/xfYP9ycQ2ejmT4gNRn5AtxsCQ1ARM+/Td3pTcIKluypXp72tO+
FzD+xkNynbFWv/uaq/Qa1WboYRD2K+jKSAvmrHBnKHXBOL7sVTzaeajGdQ1BhwWv6ejq2U4W9VJs
fOohL5nfp0kSomV8uAzXKtRN2vlosscV5nt3xDBY58RNJV1/kHuHhmUff/9PJuXGBCFXJiuZepST
05Md3IWAjbtJOI4UYWYfoOgLEayIuO20tGXDMNZE/sM/PKaAVAC5JWeQtMohDk6d8G9kv5dBCR3J
4RQ59JMfad8PDfsJfdj6QG2CgpNxbGSnAcOo3DhbkPVjuFV9k366+ejXfp4CSyz0l3QSAW/ljyeJ
p1vkb8Xqb2jbE09Nen5to8mgoKuZVtEgZjYODfo3lGyxqFmpy9hbtgjfJ2NoulSp/Y/5BoZ/dvg2
bJ/iuaBriO3lQIiyO2FfGX477eUOdLLuFKUC5d8wbu5iLw1tYht1A+sf+PBl3Tfs2bceQVIGLBFR
Hjo+gGEBrO3QpsELAU0eVGLqh1ADL6Zbryt+KoJTmiZ5meWNqopsngEZhkwdhH+w8AqS56MqkzOh
xfbr2Nw+/qe18s/WWrgmKEsg2+gnfgJCDZvMMOf1N982gy6fFvygdx0mBVlGfknP6YPlQGheu+tx
NFLzTjKkCsmnOqYdPOAABQcDSf6/49PGPkO5PkqF2tddk435zz5VjFv3XhWDbiBAXWRYQps6oAwz
ItTS5BnHPhWzHXCpYSDni+SDVeduBM9baqlhzMIrw6RzPRoU5MMcHQesV+1ddYyRoYRnUY79brA9
eD8KsHyMqCmy5MdGu40FlTuSqM6WuToP5TFj11lrMEi9MH0MB6DtN9Rk+PcoTy/Ft61u5EvXr1xB
V4xNthszzJ0hAuSqp27u1IIolhxZiJozVuRJtGTujrwy2zRKgZqTg9WvXTP7y8tCq1Lp3qNqLbzT
KypAogQKbh5E4mEz504emvvBSMKy2ZFT17uzwRCJoewjmHSctj6ub+1r42KYdARBAqz2Yn4lW9fg
jLtdRluxMbCYO/Jn5s72LDCt8FhcM84varL0IJBGp/JQ/odVcQyY0/ZAshO33mUC1q0uE6YPBNt0
HJkWce4ZvxSi6CUen9MhTpNiFq0a22RF+N7VtwXU2Y7hRo9M1mTX5ybBlGKoqxw+i53PVvSZrY8A
LDmxRInxxxqHKXf9Zd4H2gLHnhSms5j2arMNkwRJw51VcRODdBbvb6pGDagNkWN7plJLgXGPaRz6
T0Nj/1ZDVyk4bId+6lflu8CZeUTD/FCDN8l96HhwIPe8ObOKMk46x7sd1fF1s8iLlNPmKZ3BpgI7
nJd1c6/wvW9huf+i+LtwYoQdjkyLlaCNOr8zinIRQshd7eA4hxd1XlLPXWP5Pv0lg4CLXjQkmB40
i6oO5F3li9BaSe1P/V42DKWWEk4tuGCSkbW5kJUA3rywO8YIRG8SM0nUaS20gq+Okj+SJpUrYU5/
j1CUTkk6lADPw3UIp3EIuMDp9q3WyPE5Tr24uC0zpanuhzlUr+WX5brJMDjkld2X/nKil+XOBSYH
RVejF7DZ424m7lGhLJ6iONBnXFqKYGy2v3yBUyFl58s7LQNx9DAagwsE1zA6fjZZDl4f+Oa+cC6X
ZZdbcoOAJOQsk7pxMFPh+qvivyv0qZGHcJP4tdkS+uId4MPvOFSdhfudF9B21C4aYbE5O6lVAFMB
HS8zwZedkuDhFlNbNw1xTm7DEpZ/7TdrEVueosGZvgpfG55lIpX0LNPgr3ghmy1WaWkWnwfovZ1J
tYRkh0x/JGCHaGH5GJcViwzQYfJvsOLS7ZPUzz5thsKPcizKA66rSnwBh0uZ+RenTB6dd5zbPGPR
dy3Z4TDGrGxJ6i6qyB/+K8b5hsiKPyO8LTmMM4wR+tmJIBX99KNSkpzpWUtf8Qt9L12UgQyUUo3r
uzLyR4MrGNJLE3gV2433g+EUDEKgInhQmwkZ8Jt2jAEkXKcUSUItalWsHKcroUQSdlbP/Av9j5sh
izBmhIb/YyS49GMYjLoHRpNSoowTu3g93q30xCeH99IDpzBNDeulLPE0ijRRycPMN44TqlC657IX
Gx87wtCw35waC4kWfrEtcEN4gf4RNGjf+1W05TgaaUdIYuMQIVERR1zp2om6/jKCKigZne5SYZub
8Anbfo6rw4Ari2kPDk/0DtLnjoaT0Lk5lCLprlpVefmDjO8MgP7nGYZgSinFNuDlIAEzMoEW3xSg
EvyA2/oa1TWilbHhU/ApH7dLFP5MFZl2IYEeLO4zYVCOc43J1GKMvRnuqZSEaNJeJ6xdR7izp7T+
rh6Fm3za6G6OXoY2SE63F+fJ0nTThy3UdwnsYOBxcT7hopj6NT5ifEzsOa0dACYjVXmbYa28t/dp
GrhIcm8Wthqn201eYXL7lnp2W5UEQZ2wC3sukGfXrJWaITWadzL7eM9MJef2uVWthQ3B46S6iNeg
9qUYTHE7gZueWPCtlcjai1yEOz6YF/DT/XAdGVcqqnF+Ef7zIC3RgOrC2ABq/VZ4Cr3tNYTu4Fh+
hK5ZUiIcKZZ7SBQIaOg/JQ1lwhvHaBF/xpEtFjeF8USclEHCdQTuO1657srqAjHvP6xgbXEfE5Kk
8lQNaLRa+b5DAlVRK9Jwj/4Xh6LBRm7h+sGDklgKnIwspbVZi+4txYlqYCEUtUOVeweQcaiQ8pzf
p01Bd01YaLQdmQfXbmfBkDSRIM+5y++zQyvoCK8+dyeysjDkfJg6PY19icI/NOWV1/isk0v69IMR
LDPxL6tsFd7VRhfgH7uqcLhd5PWAhsX242j/M0As5YqainB2t279ZJrIJBSsefMWFgqOq/y9QzyY
klErWb0LolyNH0p/wBJJvWkGLS6Fj/hGZSfmDSE7rG7ZF/D3GfkhescMeENQFvc7y4AsMegAu8wd
s3gSpxzcv3Y2loAuKmqA2lcWLU42P9aB2XeYtR0SZOLBf4nPx6cCm6kXEPLV9EM3Ih7KNpnAt5Y5
TwqwSirRPn/d2ITd6pcIZl0GG0YIYGjqd+/QP5EQxPI7QFKdZtaOCkaEweV7QOBJDzy93vKa+Knz
jayUJ2034RZuCQT40FXg8aNuTJCpFsHOVsTnU4C3L9akNy5v9aFzQ2PfEOqrMEIVj82lSR2DY4T+
bn6uhxrfbu6KQYeIytwP+i17DzBGeUHMst7QCXebzMowcFtdeGXf+a48IuTjNEgDbTpG1O2uJfMj
Hc9o5t6/npLaIoqKzbZofubY9ZVm3pSELfuEwiabWQTjQpg2NzoNTVkEu7b2B5o8yYIVLbc1U0jk
8xW97PIJ56Z7nDUczCaIhlLasdNXOVXI7U9I+CniikfJ5YJBKx/k5khyfGn9he9fRndUqN5dZe1K
a2+ME9IZBMxva6gDmZbvSGJvEKLMxGVr8F/GSSdA2l+tuofYp/fYDB7pTPzGIhNNw7/5Yj7jXzZD
dz+PxoDm7eZlerA6fNCyWq/MRhSFC5NUin1LZXHiM/49ciDGv83sxLpyo8Vzo8SLolnQVsKdqC5A
xvndyvV65pWjtxUrxE9VDhGXY9/q0SWdoTmc4TROBw0I+jPeMxRywpTtRLQ/h2/HCqlGO1uPmVFL
fmnzqz8UAFQa8SPVlyLbiTAwVzgxg2TcWDJ5bmyUhx9sjVvSuyvs6eDbbscJvXNVI9kwkpL7iVCE
18/H0+4cNWWCke8qc1f/KSIllw3BtN/WB6nHmS1/4ZIr9xsza+JOq4SQvYGP7hsh6hPApykSZqzY
ISVAPbMZKylXyO0kDruHgfra2rVvVckQaW6I+lb4GF/f0id/SL8YFfdBVu8OfBdfRGFHjGhVdguk
qjERRKTlagPAAYWf//zDdJjXDwmZhdrMe7Q6mjIh/BwJco1/Qu7swRlfL9vlLm78pEWfiJJJbgFw
IZJy11gN48bwn34Dk1VQCVNhfou4OA5Zd91Un9EyeIFZrCjEYpx/+z/EQhpVfsSG9QaErhTIA+HJ
4KMnvBWMY4mnTykCilGaKLXUWGkJRlMqfJ7A8R1CIT6T07bl/US/SUAi+Y4ov5EfAVNgcIpSBfOR
4arK5sVR2ho1Mp0cJXSjzJxPP2IQD8J3OMco7bNEjm5eZO3sbPlu1RUVSOcveRzhmuCASfMEACWW
siv8bLgtKnI7SV5YaM4v8KDwE8ix8jl43xROL0U5m6Qe2B7BwU69i7D28pSiMmbcvBJSpzr3uINi
4XNCuputHuNq9phBEsqJKP7sYXvuHQBSdADRlrszUEG8YKugs5I00hSmxaDifAqc43pKIKK6NRCa
807bOiZClVmVWL4N5K0UVM87/Y0x6FuK8rHNd06cCi9qv0Rff4jgaw9QVSLSX1CTUAHLNhiXRt9c
6syv18ntteWeYQX3SLJ1UOSWf5AkdKo9MfwLeOxvTHyqLnY087V/k5+OyPz0ittIq0CkwWQpWOa4
hnAsH1pqoq3jABEGLTY747wjlFrDeDjrwvKAgvwkUHyPsdNQRC8OHDZx6GX5vlMzhnw3dUQ5NwaK
BzGfDqnCSc/Nx4McijxdUaAeMz9ksplTRAZ7kvUS9K4BbHV8g2V5IFlT+p035mSaD7oyV85z2TaY
pV1g3bNf0+M9GeLOVbOTxku5+/zvrtj+vzy2Z/aq8UOWGbqXvyup6ccShcCGZl2oScCJR3O30IqX
512+FCgDbUlwDd+8dAFKql7N7HQeCK/nSyzZbv1wyD/Au7hOtoc1XhlBhnEIRfZuQAlWMZPY2MWG
R5Kh2wgaR+Og9Vz0vaVo1SsdLAp73TrqtpKJ958nHeQYL9YqUY9S07DgJ4PuYGhoRTSlVj7sfLJr
kalT2OVJ4XoXheLmv/213oo8GcIeTo9o489w+ZZ7rMqWAi1kEpoG/cZPxOVmreUz3BHqXuonS0U8
yklbv3ukmG+7PTycGmLOmaMGZjcnPcxCqUILK/4DQf+ZlLN9hEhVojG4oWedaWEcdxs4EqgSHay1
AuOJm3GIMTiklQ9THg8LECa8WghQuyZc2FW4b0LxLsz/sKDknrPZyWRNIRky77aJzQl2koGcHgDP
LVNwWGFqZyAkpCwiVPUEXMhwTCTKP87ISwOU0Qq3EauZDZ0gOitlJ0RteFkrB4lM0tRp0yls8jss
TDDauEns9R8OWF2tkFF/mtdjGxdW2KKnD3/FgfulAmMRhU0HINN8XrbHhH43RMfnaGzHtAc5OLVa
Ged/6G9EdRurpwS/rHZVRjpyHW0URbZ/8jSWmZ8R/n5eh1bI9U9o2tM/Cvj6PWWFV+q3vF6gGQ5i
iT0wRyK/RyrNjA9xtGkbZZu3IGfsAFZcSsXRK7CDsihc0mTtSuYzke+WPUtqm7X28eDQqWH7Oid7
LTlHgCh9cYrtCozEtZynQszNQuVyr+Tn7XJQ5imSEChd6bzFzwHMOvwzuerM26Ek8R+K56OrCoDs
cAqHVszFciohGYboy0nRu3jq+Ldt6lqpYBmxMIlLuLH/B6pLZatVJ9gre26vD3Jrb0aKGNUo1UB9
h4msOZBTC31+IfZMaBeRDrT2Y90QbHKZkjlw7PETaXMhxFX/f5wLVNeIvMuDu67CJWBjvrZL55rc
86L8IxKG7LalEDOU78cJrA2LeZJYXISZK8lhqijCsUzpMOriS/nRD9vFFWIA6SPkgESmXxtvTpSp
7MVDpuFR1cyIhAGwW9z7ABL3VGWIXuEMqOw1Vn6flLjJLbJ+ytdv9zHU7TQpz66V0LZPGexcEmLy
EOHNukW8lNWQNS2hSRXi8SDKfHTP8ZXdWBEgc/IThzDTREZWP8KQqrNKxWGUy/+zrzfAcFtcIiPB
+7MIB29ur/H4DQ0ZCt/XfMB58ijJdDmPRQtvDZ0mkH1zLrFET/Vlzigo7UBgVckSjNiHrRaV436A
UeCD2eGuH6QvIlzkEGtdZR0Eo/VkWQPIKvKOLzVWibjQs5Z3B0dA0M7J9Ue7QPqGK5cDu/hGz82e
tfonOqiRxexq5NcUJNpxK4fzyq0dZQExNSsQFGAe0ZRsfAC84E2rKFwn8n2HYrX+Wfv4IZMb4LGr
+zaGJ4S+SjARUyJpPVsdCP1DOy3wWYIRHw1c+wuXjh184mX5V1wzW+6Ex+xdZGUxBrsfD/D8fvot
kwEq86CwT2NKavujaTsP2aFxw759t3MG411lJOR+aNYgHKig+OAIzDsRq13pofB+OY5d20AA+jmy
HrW422hVh6xYFOGI2aCr2UrRiP0bzaR4py7T2HcnIjiRZRmeIi7dSm8xRKBS72yu1wskCA1bV9bm
//FzU6oXS42PrS1ThfLC/KrEQHAfGZORt8AK+Ztg2RAub47mSxkK0HI2wzOCA85+J1ojpU3za0ml
lpN1OVqJ00YgCr+Q5RERyDSli+qMsb0kPuAtw+nXp7sh8BBVPdl0wNxBx8Ra6FPdHN9OZWFeZXyr
LQtOeVCw/M2GHTA5jK/4sQ9Upw2bNxFEAaLfSxj1zcWWTfmWrwOusO0F/Gph6qceMxWCu+Elib81
0MbrwCqWhzFYze60h5LcHF4zQ2Yp3hdm8S0RWSUXRB1mV+ofujznYOgTZI7Burjj18WTjr5L+uvn
FrsXxW48935BaKDGQCaRzDfSWdeWWQSNK80HcP85awUWb/1jvh/Lj4yh25abs0LTf4M2z5IrVCBD
8A8fs5Sn6hg6UmYr2heI1NRobbuWgfb0c7wyXg8fp4WN8djklZTi4CFb0x/+x/7J9QfjPHR1n9EV
yN0/U/YC6HkaziM04w2nM69griwm9viagVLpW00LfKsGJy2hLzgVPaE1WvBY/0WxPs49inUocBpW
6Kk29ckjm8X8oWti52AbAtg895CrA9stMmk40vs/idDXbOI/LjevUApYwQAjEb7DWBAR6eGVcGpQ
gBDE6HY3Hc+RsirmOoC/U9QMvIudrWYGcL1g/ZSZ0seQSG4HwZVemVhCuVtnirU9Tu5EMLcmJVXm
uK85X8u6eZX2UmQP1hcCUyn/xd4INqMEVECIBu7T+wM8LhBs914Ucmc1RxtXlaaEfZo/mbVrfeM9
l/0W/c8oXtot/R7SmJmTVSGedsBGzWsDsbfqRylYtPptfMhm5E/Bq8gg19UAvcA4D6jNXsHXD8YH
T15RQ5R44s7swc/L4I7qVVEWqzwc2Clo8xjwQgN3khFVB726zmJNYWXYbMZXRM1QwKGM7wq5yBUn
vy6AW6eEJHj+/AGTQ4+yvIEnsHPOK9w3kUmhPnt2YDljG6R4+42jhTU3LAwPtx8MK0GTPAxRNH3x
psjCWc+eMbKSO+4448XC2GoSwBx69LzQSENgCatjxcsFNsVnKjCaWyRqYnLAP/0pgvqe7hAKoNb3
mExVtJNkKi4ylE/lfJnbNsNDdLTyNwmTNilgjgKOTcVZkQdEc6dPMnm7egS4Uplav46hV5egPe/M
c8p01v0a27MrMzW9BhXAst4ZPZlzmU2Sd89B9wIxpZbiy8O+V2D2+dbxwzDNsmZf+9ock3XPXxwk
0dTRbr/I1i21VNsDBjKRNcs1Zk/wD/LF2Pt0S+NhYE+Go7vpofU0n/ECSVdfyGnVWIo5svPZbRMY
T9vHicJDafczux1DU5Or0bylB5JL2bPeuARzAyCfm9OGOhsWHesTURF+RJvSILk5hY5spKeBJ9AB
4bXSCoRxFuLjq08mSjewTX9nguo0hSprf+C21t/buaZd3XWcH5nJUIWh7/A0v7FIEWW5INUB9/Ad
voXEI1ah7/1Mr9jGWe15yZQcG0Ii13VleWifXk118avyGq461HamFo3j/Pa/wEwe2zadj1mtln09
uK4hnc+jATXaPrVrEmMbKS+4Xk4tsXB50MPomrg1j6qsK6M3NyvmIs4QKEMKA+fTs4N63HQqe4tM
G0k8bWxfq0AE1F4C7Poe39UKTv37dyLsNSFTr2hne19y/Wm08naCTLOtp8mTAvoi5tVZJaBHXJ2P
TxjdjQc0HX2i27Ds6nDrXmcwzGO/47YxJ9KcMZx3Z8/nKHegi3Ge1igIlaa1fGuxOeWOK5UvWUs2
W9vN3Qeisrf9JIS6ISWq798P7vkuruTCJBItO/6ro8XHBQ8afZI1Ua2TCvf2jCojLAH0nTDANRnV
IhElfMESqBDxhgC9Cp9c7rmyFHIPL/7GF+K+BeyOeYaxlqKClvzuUsW6MaRlNy/qgd/fFuKVavuK
JDer4OFuBLv2zbjPN9etgYI/FLi8tXnarHYlFlkw9c77ybHMxFLF323sFzrIgoMFhlJGPhlR/CdG
PQkdPGpXdTECPhMS4og8I0ZAz519ADSOJDuGCg/c9K1tGIqqwZEuS+F+e6GdOOt5M1TdS7+Jfv1y
IrGn0OTYtFtVaPxLARX70SQuTh4UniU7mKEtiH5kRikPUIzPnTJbRfES7lKxd2M/Fg0LZKs6/RLt
sMZDB6iya3Qv3DQmtC3tjJENMlCK4+dTnW+jLqaTBAXpCUPVcUGDqTDV7zzNbNHnfUW6uLsrBRGT
w+mQ7+57YEduiUQpf8AzniT5obnIwuihQLDi9l7CzLd2Dz3I5CLGaRjI6ECwvUgTGBGh0xhgUFUl
GP4Qa8n8yJFHJbwH3AtuXISUs6ncMznSSjmngTJGuiCNfm7chacYS6sglsWphvhId8sB3eYyQYoS
4sKsi0trNjUzav7UIk68e86h2Gf2h/RfT4TIlIxu4FanekvVJaj76xNAUoR6SI3B26NFTXC5v1Ea
wnrbYn3iTsYKJmHjA+FJ3h/Xhbu8EaH8/PyhuKD7rrHhzs45kZ5RjylGWQXg5Jj+cqVgBe0pBXSM
FG7TvV1VxHi+3vpl1l3CFT68X4BU9CdPrYNoqH0nSwWiEq6aYAHxDyTVqg7JXfqTFs4o4/CNUpgI
vMHo3QQP2Jh7q6AB83dxOMbkkIi1kfhzOVrB+JOOCFwxt9REtzRlSFXO6MKVd3Ohar8RADE9lv5u
blKxfh+qMBwboL+z4vYHKdbkE/wsL/wzpk8hHs/LvsgB43vevzDk+yCM9Vi4YOx8oTTXRrIWAAX/
LZqZuRRKXjAbEwFL/h5Z5FliMjYLzf91jElP51Y6zhDP7us02MKbgpFzlr96nK40c4u17ks3QgD9
kdxTcGgozO1NdwGYIdPFru9rCVT6LY86TjPxrEkbud/9eB3ZvNeA9pOvFEUQx5m0ft55qfubGfqd
D0V3RrnLbL3AlABm6zV5+bSM8UImOw6aJxqd+1TsLbkCKLVNU1FztsLwRLxjXxWlyhMsAU0L51OV
fLGltbR0JJfWjYh+Q6WveHnvvB8Nh3ED6wVbHXXLk4G3sfkn6khfSM4m8ioan8+weNI6Ltdnv7OF
agumYZl7zbajxLJYvNcv/Q8bbP67yVnfMUGHvSGMjsOh0K8/RWaCqvZb7CLJcJHkTUo/EgAxDWM1
EolzHXPte1SYUezA3KHkMTe9r8Cg26wJLrM5zKho14OqgjzBb1KKFhBKx5UJNrbbgkssJoJ/Xv3e
DDFG/DeTYuVqLC/DZverroMxaIg3Pj6dmKBw1BTMBiuMIl+6lMUoYfatzLzN6x9mn/P+4O5+k94c
CphXk406prBOlpPwVEqOotRqY98z9WpAvC+s73aHVMsEmh9P2EytXhN01XrQCp7K1ZhUIKVkuLBr
6zOKJ37gRnrJyzeCjYt0LZqHHJToagzXrUOz1q6ioXZfEre8Xgp8eKRmjQ5Wt87pmhCk2N2sAQEw
aAAvoNMwswixTLA33n8jTctEfTd/z2dAoCWDdhQJbDiiKjFKP1wkkRO1HP76M5/hVMyjEChCl95f
VCw7elhWZyERQDdXBqn6re5dVItPJG4QYodYTLJCFUuBj9sgbyWW0Pdz9pcTz0BW5ZTLUTixKdFM
tutheGYD9NTyDdFqcdEl6lCOEzB8MQ5NycWbKIKtkWc+hCz6PCHDiJfBViEbKrsuVdfAZVEksxex
RRq3oPrxkafAZrF5oXJl9KMHy6+47ooAqAz9TVMUrx4nFzsesn3L72312gPDdqffP3KP2xMda3OQ
eb+uChr6qO3pDvGcpxhVMpVaYYOi79hOe/sA/T3nYIrb7hSLz2wjAbD6UsxIzd5XSI89H+GmTcKg
1iNE4Ge30tYuXlOPCFuWI1x4JAxDoUIsvbEVInMxYBkgE+KrWsGKt0mkwNisUCedDEJKEcO4zGNR
H+Va0zgj7xjCKmIg9eNcq+ogWSAAnR3fNC9D6uY08vEGJq+FmTHKJ1bzj7HJbU7/VovZ2RKRzR1M
GCDT2e7kqZ5R23uz2dAUJBWrvT4D4+oUeqKqhre5au5HZh7Ofiyfifnxw480jk/hc+deZhLWFaiH
f3t3QLFgTPfrhsGnxKjWqoLOaGEO/rmNpA3jytVNQBJsDG0VPbNAreKey8gdCn0bFbR5d9DVdB6r
3d8gIJicO9o1bDW4pD7wyGypJTHWy5wTKnhi8NWvmSL1X3GvtnYWhzMvJ0UKoBdsN7ifkH2ExGN+
HOX9lbXu1JpWVeiqQnXoPKStwQZUnWa76HzlIHNV8/FR+0UaXDIie4pHvmtWyfqHTzLT7prJ+z/x
i+AUijjbYZEscl89Bi+FCHE5u3GYhXvqvFW6GcKGCaAdI+jW0gYY703utbtj0I27jBM+lxQg+1tm
EuPVTU4jbV1rmbfM8ViUn7Vlq56AJ4yShNR3Oq8lUcL2NR8/x1jE2FJJ27Krzp8pWrQjG6mmHjpj
EGTrJjApCrvxDE5Y9Sz3gRHE5sa5GZ83PfNXAbfPp+vsrdedsDz2z7p7CT52nmk8QEt/qfeniizi
dW0ltKOde2pFus6R50uCDDpGR2oba33UlzhGMNNv6NrUQHFhrFeigsheXf2NwlNVaYXcm8xgT+lN
eA9YR1WBjTtziYpmVvpo45iNDhS9eIVUKUuWasRmIuDVe554F54k+o8M19HWRd2zmhtwnpBJ56Wp
q1Q1zZoelmqcLxfYavH3Nj71aZkWCAFElpVXW1PV4dhJoAVtM/QigJSqrp0fWNI9B0AQxl2UgLmf
cAcxRS2xxnVBZn50YtAvxuJGBOfAobyU0I+3wQrVn2VVQN6aXsCQlQoFozJ8MPbtLgFvVO8Fdb72
ddzC+kS6gkdK2U/Pt2nuQ0L1z/rEhl03iXrw6Cuvlp8QyIt82nTbj4aNfT2oS3y1ipm9wtBtttAm
lq4JVOycw9MrqFkj1aP7+fisMDyhx+KPfuxtnFKcLL004K0Mg3NJ1S6CoyOVkFFQXCYwopuhqY47
HDCLZgft5ECwit6+4UBR+O6bcNomzps8CjtQzJH37m4dP5asg1s9ixXnmtX2B6rONlpQWds/8+HU
yUAbmsPkhN4mW5rYceALs6Xb29HpQSC2AGhOm+1o0z7i/UgTH01q0peQDJV2ymRENKidV3r2xIEB
vot6j1J1ApzB/F2gtfBM37ayQIFXicMqE1DsaFeV0FbNc4H0S5pGplQ0/mKp881uOFAXCBEpfdiM
kjMEOE21Zx1g4eRWJusr7fJPZwPBFxwR1hPz6fmRbY0Ox0ZNSs+/scN/sRkKSCks2UDLzFxkSw+Y
921KkXzfQgtCBCT+89RoTt7wXxOdXon4N2IhC+X3ysYPI1zSwdc4WPOOO3hY5bwJOTtYNlyti/zj
R4g/dppcExRlyMjszE/kJyFmtC00o0xxEoEKedGkxcH5Ds8qlxbLNHUHwsLle44XkX/oAM3O/uKS
qPYly/V1Q1jMQnBZPk/06kmhAQbHA2Zdo+I0p3XL9CRF6ojn0u41nXuUpcL2TwOUeUhTHOgTftd5
saDqIViBGyfs/m2Ck4YT41Mkg/i/6KYZTZjq1vc0wHWBzbaJFtBI7jR5H9PviqhiI7SxCAN3rJZJ
XMVV0vA3ej56URnzJr1KqRThm+iSHC2mbRisKZ4Aes72rc6yU4DkhXAfTd8UDqNPLqtFTmltiLk5
6FgnFMVXc1pRW1hu0ePheaLBTtRuSjCZa5eG8W4iE/5XtbKTUIRGNEvp3mNIr+nnSwn68ljHgf8m
spt6RnjtRIGbJtKiOtNe9kz9tkk5p1LjyhqVKfJAhrzS0C9ScHAe4MBiGMsw59s89ncOeQlW82zs
r48hYfXS0hfcx2+MghvbzsD8Q4Q+l6INqJ5KG6G9RM+Qg8m7k694zU9rdqkyRVSgBZKl5aCby5cB
6TzxFhIoojkSqaZIZE412F+rPgG5Huoqw0aXoInsbX2qjwl7+9TjPkZUQBKhDtAvcLEv1NxFR2Ui
oePhtaSURpOPWkUtATJg68MZgIckBGmxg2kEwPZO9D/p1VAsbGazjdFTvOjZ9K69M+FvziWcR1Ic
R08h89uwcOocbnQimdUHfKIsybLxf5v4SEVVXnjncL5TDk1RLk1AGQ1lI9rQqnaumEPMH1vXTRmO
9wveoucBCD9zR2ZKn2TmF426ZM7kU97V1DFBZMZ/yUpWZbrrTJC7h8A69lTb+WaKttaLQHu5ejB1
GCwGLKZzxPAA/Ku4UhGNKluZKUWh7DU+/UIal428IsZLaJZJtdQfEemZX/AfTFa5GWa+zEbQNXFK
1h4e4OFCWscen2WFKA4+nsAEx8B5CAGMruxdghJm9DjYYwibzZOQfucOjcmgrVQ1VHChaJebclVd
SzPEt4nBjPA6qcHdMPvTaSTXCfYZx6qioB6n8LSL4ogIhu6z1QGCygBwbgGwCSQg+g++Rceq+aU6
e6cNYaTt4+ROC4gb7n/wF/o17L1Fge2WbhX9nsPl/oOiQdeXxrM9jEMIH6V1USD2d3cYtBm4H0Ji
lGkHtew/oYwQAwHH3s3hu+1k7YMWZhPsvmj6UiRMfPXyGRZJq51S2/sbyi52nXE0DIcx2iBFEPlL
3rDQF/OnjLcrdsB/nmo3wYkqB3HTNQr8BsRIJv2kDq2JQsFdj8rMPNT/025e3MrEJTU+thOQnLGz
mhZG6gamdOfO9lgfpRDsKN5y2QgyoABFGNoDhCy3lTBDslcXUfG0YUvmmbqbTL06QnQEoV6fWdg0
tHvqskawr29X570QJqq90eCwng3/Y/v0dZf+SEmJ5ulTh1T5VN4vr09IhEjPNW5++v7YZwjDgIKO
K/bcSEqmAZuH72XnDzQOQrycaKHh/y4jW/4KKF3hp4Sp5WsylVHV9TYPiVB98c3yrv8Nb2gXZXu+
e+9xP/adVsqDceeo4DAOVDMxHnfJTlWJKJ5+zbew4/wdpCzqoAYwbzDstyoLbGqjdoRmNw2ZQ6t2
d9Vfxb34HWVMQ26xvvzng45E1iIH2Wr9a4jLk4Kg2lUF15EzSPnFCw3An2S4yUSf7S6CPr3yppmQ
ss3UCxzm7xoKp30b4/ruHzR8GB92fuoRZRlg6/PKJyErqvX97sxbDCGMBB+Qj+fE7opi9XPoJ8lz
0CDdbtsmDEro/jONy32ilDzAU6LK1opjxzqq2Reyr4d9VolYxg7GnqXCBpCRs7BTnw62aQy0NdTD
HlzeeswrfDPlcGeYQpwUfszoogOxA3RluftM74r4y9u1bvHcx08BZwQRusMIO1NK9PDmFMaAW3q7
IFSvxtklr4G88ufVuRuGq9vlIyVVgwlk9qyg0/InJ4atYnVuECXmux+jtjBvYrWF30RfDUlwLYiF
OjeNxSqKIChJqLsLtNS7pHAqmHymKKxKQ9sDdufvCbXS4p/LrHtzYmFSvOp63FrT09Xnhh6KXbvi
L/XQMdkqhScFiQkqV/hHhPVhXT6SCPMbr2bBCeTqVcdpB/CoASI3hhPO/rwASuOAOEeKXXwpfsfT
1tYJJVTFE09dGCijaf89nGTxR2sk+EQOpMqD0ujCdqyOkJJE2hepOhg7h47Mk72OQY0s+w2ReZzW
MYdEhYdaDgcNVD/jwcng/WnMuA0u1FZmt6Is/WeIEMzC3Dpm68+/zq8bbvsMc3h+n5ajKncG83Ji
4hP/tyoyk97yfx6zZahkV8pwKkMPt/HA8FlDL6rnemu23jYuP8fTfJwuRPt19GW7OMBB+EBAlFtu
XcH65BCD25yo75DkU09s5KzG1feqJC8P8iydiYfV4rIP72ut75w/1IE/42SWRECqdnurfEV6i6Vq
kxvjDgLqvTREpE1td3HOWPgDzV2ioJGhDlblN3p4MkuALWmY4nkmuEK3rntGk9eQ4sa0C5jwCX1g
LIMyzNNm4wz4eRhJiArIrjTVVkH3rlZj7wqx8pJ91EWGlHKYkgioxXvINlX2RYwMKxVevreJ+ktD
lUajBZKxEQ2NUv7grrW3GOhbpch+P7D+22/YSbGUtmoiKtEG0rbuwSq1PIp2uXdt088DugpTFHwJ
lUu8SUFH4jEs13IrY1uL/AuT04/SZNLhAPR/Fg6pPrQBi3rmM8WkjTq2x/u2NsGhEisPQCKEO9c9
FiRMPkamRKDnNKo6Jsk4CfpNCSFdUfPDgXGoiHjV/ylMfOeO8/mAXxCA8DIgYaJRyyvAua55BVPD
prwaekVn6pBNUkjzqCTfmZakw7IacX8fl+7XerhdliVtV1yId/5dsRvGuKqOLcWLzZEFai9A00OA
Gu7ccAHDlpwqFHvZgApEiYPBF2RBUf9hInmP5UgWLlbbToOiJFuCZbFbOGStDb0s8huX1TYNyyhO
drGSOvuDBBYgUY03oFLbCY3Dlvo0jU/oLHFTJzHUkp4jW6f42EYGEwK7HcAmnIVvzFjn0FYCxhps
Ig+Hlx7ansBgzIbPRoTRPsHhsJWcNq7kHZ5aZv58T5svdvTEqi5yGliYc1oZDecSpsNX9uWNztpL
TOkO/zK6a9uz0GQizgGVzx1E8IqAwDqe3XQPI/D+g93qeJHLEEwxCc9aSqkOWLZp6XslfsqAt5i8
Q0VyMQXY0Mvq6UGy9yh0F7b55Z54HN9p2sPyWi289H1sr3zBOOJ0uy81KALixqZ29Iodm6iTpBYT
vhSXp5cFzLWh/rqAaOGjbZM0QgV+rUe6GfaxCAsQg3AU/vQsefBwv9fj0qW7nhGaP2XwlwVq5vgX
TSpWWWA3m9bjH+RasaSN2tSvl63bd29Bp0G8heEjdcbNaWIjc3ksztkO+qODxBAOAOeC79+TxIuV
uXpXysZOjEWh51kHhc7KRfjuCXm0dUhthG5Q8Ljp0mo2lz6ZONc+toHmLLC/QerduO3a5HbWOt+n
W4izbfWatIzBiH0d77Ko82+KxW1dTvaOwD0INrRdxrBItK1QFPIdZRsX7mI2GmObzPQFwN2/ZkZG
UIWLUPXJdA4+/9WSlXMOMC4KQ7HbLJn5nr46KfC0ciIJBb1F812qdqVaaMzwAoqGhQhLsqxgUTAh
7GseOzGE6Zzu1dpgNqMvTGoS/rMjTUbJsFHidgEZ3pUMwJOWdK7hHXaHBfBjypRA7BUMsnscpBwA
JqPb88Dywvx57xO/8zTy44YHUNR6gFWhdAyWSq42um/9q956+u/k3AH1afvUISo0Ke4V/T46dV2V
d5T1SsSJtJoHZ6jVACHevaSH/mjNVhBMA4H5l2CmAy0Fjd+3Cbim0crh3m+pHZ3iwT4A3FSizBKK
5zesW5lZTlbWUBzvtj/OCOOsytSg4tYsCTpHvjH8mDCHykwNz0/vyGL/3X4Qqmbf46JfbKpGRjdT
JKgYlCZEK4GQwHDpz9m9DNkbylKt+9nWkmRMZn6VxGu7huv43qAGj45o5ZPw3FROaDK9pHC9AhnY
9svD/Di2zDaeIP1CziEc3Y89RT2wc/gUy7oZxkGIfHQQAF3rnGsCw6gIcdHNttlZ5eyby+rM3RHd
y+BeFZJZkwFhup1uIk2M1VEjbZUA18Z96cKj7RJElSYqvX8sCn5khV4pJiKvSLg6bt1aOiQyUQqv
Nb8klqQfS4HPusjRat240w/ksOz7y6S/VyFhAyrDFT6tyyHu+jNAmoGD2vZbqeIAgt3lIQaARnNn
Iqwdd39MyTthbjbdLCxYYGxFOtCFLXKK+XjIV+5N0g+NXXuHuT70dYA/K/u+K71fLVosr6Gdr7NR
a8o1aqvLSv6nHD5gzCqbceZmJarcMDXkCjgu7+++v7PFNRozzONSm1GQ/QjuwHHWQcs994VGbV3M
d6G8CbYfJg6ugvS5MQvefvc9gW1dXWkvUMz+XXE3lrZ8I0hr/Yl/VtwIXpf2AdgJpif8lSiGxc4t
PGwhle4fSMAwW+lE3UmdRbQNv+QttGTUQ3eAgLiqU8PAJH1s5jkrkJVByK3ZDcRsOtqHrN67DQXt
WMyJbvbpk8YOThHCYLKAqtxO13tsbmqquGKcZxH/jFSrdpmaRFsBP/+fzjDTKFTZKK3uK/K9lZY1
Yh+nYGtV2rwbKl1JZLn3kiihMTHJZu2JvE4WypHjfaNFqXvOTPChGDaC78seA1sE22SamL0xNKNk
tqkAS4EJ1LEtxctCyp3RSN14luVhTLAOYx4h1D6kTUHOhOxlwPJ+IcKPl2uXuTmMqJ5SYH5XQNuy
sf6aNdBxzlL+p/XtuH3SU1NBJvEaNorwkSYcyLhjfdBv23auA6eJfNqQJ5I1uplOt5rXOlU2YmD2
4FF+InC8jhhBEBXRnjtOq2PiM9JFheB4C/a5pgpTr4Do2Hv5Ab1o3uCmrSK27LmYQmy91Dpx19Xm
KUGNU/+T7+WOMU/j/Am8qA/5fSzXdJNkjYpAVafRyLK+IyS4R2CSOtTDZM0JqGVzaZjVBT7szjyw
IqwOe7uiD6PSzOkxpe268aa8pnZ61QzBRQ0ASKRC3mweL49on4S8BUv7M4UFFA1YMQ+70bXq7OX8
3ZogoX7M97XcaSmV485xDhyHC3nKPi81PqvGBETBZCgLDCZKFTXpogbeNOI8fegdgd34gdb6bKFN
i6GWeG9sAQVRp7VqTI8Wqj+AEnLKDdbE4CBlNeOJuRUeaKq2zzlD6QsrD3iRZj5jzJokFreL1TtH
i6GOPMcSR7dyVNKB+QQKnYEW9nqYyLnRLZXT3vbm10XvHJfLeB5ppqBGytofXZCeYwOe0dUlqnYQ
EwGIcOoLiDa8lNiBQaMx0WxVXL21hPtTAadVAYxXPpz3dAk9SaOF/6OR2NMrZmXwBZC45WSqztUl
yCQETIiG+F/SomM6ib8GQixVxmLvbGSTrxgJSOh31IqCMKhx+DLQ3tEYFOHsnNLmuS6zKszq2KEb
OrwdgxWAWCesg0wkZQfo2g/QiRGP3SlF/GMAjd10oKfCAay5318+l5Jyb5z2T2wOGJAer2i0NqTT
g9YUGkWm5AsPg5V6TIY85FbaGQ204ptEONXML1ezOmg2yLIrlgMocDmH4zaGurBBZvlTedbFKO2r
6qVnCm+HLSS3E0UiwuX8x7NMOPQgYuWqGNgUU98xbhCPFUBoSAQTQcLlV+NaJAINcLFCM6uBBPzw
CJ8po6+dCp5CnRNScG/0ryI9IvPvAQhhtZOoMlST9xtGs9DYyyYIOHK8/Jb05TVXj1rPSctHwOnd
pcOG2wzcWHhfmVzQaUwNImKpq2PxKKtUbPL04uEZjCmyNuhqmHMdKdDz7hxkhG1bixN6WoRzDtyn
ZAWmfDvMNJVf2xD5EunoXeu2SRJqnTAlHzdtRSkESf4k+jutGZbsJ5wm21QgUfrZv8wxlh0t3gpX
ykDDcEuL/83fMkomADwWqEDw0ivBc4Z3DVeq39g4A8iueBJuObHugPhROtJK5N5STWMr86mCr1Ou
8FP1/WsB70sgv5mLG1L3ymjuO2E8o3YdhYMouvJJ03H2tpnWPtbH8xQAlOvqdxOnchhcPjWp3aL7
o2L9Xcmw1BknjSB1m0NJK8I40vjFzjpcJp/HurrrtVkYA/9QkwLvmEGhpEDhoPp4QabSslMOVYJZ
rkzQAIPLnmL/8qPLpDA64G9/gnurtae6vBzgB71fxS9ymURY4BrDKfByUZUBUCauW+4wMfhvQMsk
uJKBUhn4eVbaZ8Fq6ffeMLADC4O4NYRMM/ciDNrYFS2c61zg4QKoJePGEBOkbHs/zMggJqxFS7Fk
CLRbRB5115ZHASlwy6YRD2eNIESALoLlQNncch/iXpVf+n+9F7tDKKShiJyskV/nz2JyXhu84rjG
OteqSH+Ly/vIYzzNSB778rYbgWt3dyRALHR0t+jJG9KfuN3XoS1R8drA3XIZi9uj4WJaHSYQlJ3k
7A/DXjh519VpuIEmB7yZTPUDzgnptzoTUtTXPQOfygHe9BgVUbuMuoZZcQpC0k1MepjKucpi+lzU
1QSAEvR+AX9jylJeCzER694+LhxvfEKRYyN18KNsuyLfjw9fYcDvyPxcp8O4HYH+zS8oKd1P4l3j
U4PuGW8LKBVAYhnu+5+WGfLmHNoWcB4iZh3oU901iUQYNzyGHhxbNiWoyQ9E+oOcRVUBU5GITcsT
jZHykc/DFec2Sap7w/jw0h+JLDNQpAX35bKq6OJKDGzcjQCRLZCWfb7zPl7veF9PYiMg4w9I3Q9y
Hu7seWp90XetWXtt3MxI7I8OqLvuafR5LQp/s6xUAlSRcMUb5I7tIoRG+0HU8ilVuXz7MCb69gXK
V2vOqet6RtOcdTqZUHQelp2nWMBWdT8XZ8ssXXRYSIoG7yq9N3648WpuzdqwJW/t++SFscD+CXQ3
hLm8I5G1XwPuamXsESgErW1+olUxZ6gICDLI1oVuxoodDNN/icMVnXC/EmgMxMpJhLQO4FWzyPU9
HrTjUG2EQsvzq1F/um8yNT6jSOZ2mHc48K/6ivgq6UnPXFVKrbyAvySki1GXFo5ShN+tUn/xoW/q
8aXT0OkhMDWK4CAP2/sHSXh62FrJTOA05cHO4W2nkttnYC+0IwaJMWEL3xm48w5oKHs/CwcmrCHP
OFimGFjJO25QpdfUxM/pldbD8WwJO3y/KE6wz4UQ8SdHV0bzePjR+ETa0FTnxVieRdge77qYIsXh
xoM50GzC3ApERWFM10o7jxndJYzERb/BT6q43qasDodqlDmDFi/xXXwxNWipAHMgCXoDYAfCMK1S
3baIJrWe060VsnSVGBy4Y+yHw4qEpMC1/+rpF1Mr1WLNTGBirIyn6kF9y/AT343TXPdITXUpwtay
sKqjv4r/FvWjFJxFIF2iu8j8OttEo/a3ER6obTtyo3MLqFIMuaIPYG32NahB9P/wliIP+RgdmxAQ
44IEXjO3HqBGDlXlrveaMl64OdmIJNLWh7iEYGS4Y4VCdvy8NA+gWN4aLF+9BnD+ADbztWFoPGwk
IN1qBW4m7VWX81w3w+lI8ndMJDu5Ec20a546Q7ogm6OIjAHvTW4RsYDTSmSb+nuPfTMnJQ3sk68b
GtgxRih1PPaaYtVcIsxYXDJIS27vkT94htHMYI3+27TFwpRmr4FrDIZWEtZlR/YzkYMdbISzOOE4
ktSGqRPw06jGJMkyfzEZbEne4+WiOKwTctUPkMBxpt1jRyrECbHcms6t/YMKl1jB1JnA9eAYDax7
DgtONN6M39znsRpWn9lFEO2+8x3rBelEbZcvUJMcKE4hDUb/na2hAsFcr8R5k3SkSbm5J3WhK0Zc
Al6RoPntB3IIhzKb4FBTLs5D4qk1DKJcC29PvQPkGjVj0VXUNtC8QcRkewY8RBzYDXR3PXtqkLkW
W1QVxM8Q0S6G8ssHXEfJxL9vYrRFJ7LK/4Hd9vjdMNYN0a8tkAByjlbJ3LBq6HUQzagkywDNQ4oa
GjkpUatb2Y+agBUG6YchupGgtXNPBHXmqoFXHccGTmX6lV2OYnXY5A6pkBXjUwajixCGMHoR/HEB
smONkKqBs7o0oWXuk+U2Q36OTdf0KPKTFi5idAdsD46pWzJx9jDaqg+QaLkTbjpDRYt0SsTGE5Dk
t/B4iKEUrbVdnA5QuBzP9VPmNfW2yOnilJqCoJxIlhi5oXtN4Y4OTWonRVGuq6DWl0F8hjfqCPUg
FmJ7FPCs/VyvSO3LClvfAjl1ZvhRj4esU7vZTaUnbKc4LKpWSWbpVRZaePk4O5XLM1UR0F50KkzF
rjC7n+vzAt3bRubiTkmwoAmky+CjOMMWTvJDjCZ5ZkrA8bTO5kdUyqn+uAfKAo+oiMkEUwWAqUcT
/l/ivYodHS4z8kz03LWx1AHiz7RG4YUtQOPtuliWlwohrNZ7CAndhyJgpOc8S/P+W67TQLb/4N9D
IvHGXAwNHWsuh8t3T8+jrqlGtD2BljwdnIeDZKcA1KT5aWFwtR4WJR1GT07EPghn/L8nVMNT2U+x
RA4qXqI3AEg/IUXCCLUgpZ/Yx+E3+NSzi3F7RxW2DVMGjJoBiMqPzxd/nMdEPuG7/W9X9EvJlMtf
3qcoEQzLLmCLRds14PVo+UDfWbsWRpa53jtzIekEEHXnIRv+Ucw5AA4d4MQdXLjrjeSS+5Vil8Bz
voYkzW6lSPoqVvwiOJux7V+ko1oFmcynGlur+DjeV8FnRu7jMnZN4QTi0JE6tY2FWLrUTIyLwLZk
jWf62ImSoINMSj5Bs42KDLvws9SbZx38ED9sL5x2DvCjXec3LaNpxlva6/tdpTrItjdJc+obrhiS
1juoaQHl4D3r5J3oJgD3QbtguoeZBAN3ghyY8NlptNDzrQtPoHZkTLsJ9iESzRqbWRtMSfVbBCnA
TSrzJ871fXUW8xQNKdBAltcXWA62raSm0RTc2Af9h6f65RVKNfnvqTRXHSsirAMGrtzKhfJpSInb
aDouDwQ+Accz7FeR0r9Be2JPdbK+qwg7I4wSRpJx/YiJ6K2+vt15RE0dMTcmINahRKnhwsCYqhix
3i4siQ/bIpQl5flE710ASA3YM09h/wordNkhORoT1qbgNlhBZbEH8xH73hSP7Hzyqtk0foJAkPRk
84OPherPIgolm1HXQ3ni4gy1ocqIaLY2xOdxy4NGl47wPT4UBoyuh9uRMpP33AYJa+tUz/A+89zu
hrwnbT1YGNX8h352djJUNON3CH014gFWaMZcRBecjX5JAQzec/+hn4aME5mm7dQuE4UFgx5725A2
HhsGzem4JQGcaxB2pWzIfrZFEtEY/5qa2j9Vsl+kajZAsU8BHoTel4QLBLbsLNYqDN7CHqK5HHxK
vzOawa5F7dswLDSh4LHMDa66DnQ0Qg28p8RlmhFRV/deZQwg9UeGWHA7aC37nPMq1DuIjDNCytL0
PftqhY/PA5GrC062ZfqDZAt20Rp966c4u9TScnVIFnY169houVeTXSobmQfelHE3sdLjvPEwX4N5
T/IQaAipIrur0bGAcyCBrlSuzhw0S5XmblhsuZ52KQwaSNeHed/yRZ1DugxDEZRg1O9NdUvJeAf/
OsInsXFfmo03YCZY9/wXPivI3HnWk+Ae45cLhu5k1C6QP2gFAMgKEerRRmXvdniTlXE56pQ5mOy9
Od7j/xJw1eEuh9ZdCH4wC65a1rY5F8j6Z3RET0WPIGuqdmygL5Eqr2Qei3m0ujj7E5g16b24AO+X
4b1FIKvQub6OToGKX/MYk2qudUNjXCbYAoTGPbKD0cFMsR3sLzC4++93JMJhkxLs04zXSPGbgUBF
B+i3Gfzz9GvF1ekQR8Q8ZmLik1Hq7tUDEoiDV8b8m58tHEPn9VlZF1Am1J4fKa5a9WYeMwBWr9M3
+fMECNrJt+5v4aNvFpjR2RaYwql1ZR1nOAoePQNX9Gz7RqlQCiz8zImD4BHsjsIpwkT8btRUIdil
c7tY8jCZ1dnqa+0bU+IWMBT9Us1ZIz8C/UDebjV4hVz+kbuGCvb7PWqsDgzG9NRSdjz1iqHtyiS1
SaAO790j2wlYK8uhY8FDsCSKYTFbrp4gXaPsTbhsWQVMrFTN+shBAntHSaRPiKai/QoEh4mGNf6c
p/PfTN5nnrDAESU700deTpWsLhv/fD+88HhFG3/EUM+vZNImGBACvaqYSwD5EOZDjyag/sTarCyC
9LV3nvjVkvlWxF9GeFyHsDAmfkLgo6VzVOOtU4O5nsZ7wss2gcNwie8KwdiFHe5QIodAxEl9Seck
efZ/wyjOa19DCpgxx1WGUzil8A+7z5D0UcXg2b/sLeXmP70CPU5xv2WNnom9ySf+3jIueHBix6Fn
CCpiNlqX6FFYsbXPzfRZH37O+5U8/2zjBwblRPWqktXFdzfoUoA8HJh+727pEqRNJCmvaKmJKiGp
qANmkSTqzTFiq7GAXrz6NkIWrCnYG74Sd8YBfkunzC5ppbbjwuHpKO5tdS9wQzpqYF8BWx4iYuFq
MXWeammiCn3v6rGHXPk/0DoDc8WG8vyp73DExIs9uipjgLbYKCFrm4A2hmjeSqkwAzYsbhNnBoBv
O2txL8WmB+Cg9p7ege+lqILmbVPuA6zn3/oF8O6ZKfO8W9T/dxkEhbeaHjDgEuChih/5MsS4UVkq
IbtLI+UsfIjrl0haLBtS18WsmzG+E40qTkP9qUNAS81nQykOTVL4MUrdyOOCjnPIV5ZgmaBgEdCf
C7kMuVPeig3/jRuuSqjJqiQR6zlIWvgQTwWxTfk+3s/Gb760p8hGKRd9FBQ94YV5smbPpzy8qNZA
BglDelLN57Vf3D0cifvMJXF/sbQU4SkOfeCqQiRsML/vwTjYOeu1tpo8BWBadTfAGQ/KDsDgvkgf
I1ck3wzIkW8+TaQouUlItcrt2Wr1YoW7bVvLvHP0uNF+s2Vyk0iN/KNE5/iSt5zXDXGR3YmqRXms
nFscCey7vwo89EhujNNsSXv90biDsYSJu48C9Dul1OTjIh0k5a6HYXeSmgfNLbFQfld2nQSWcQLQ
dp9xmXHVoPlok6EHuamCsz9M0mhimyViIOEB/7/oP6SW0hFCKu/xJAMb6fW+X/s8usxbjHY1DCF+
mEP9VP3A1x26SEnKfEft7+gjsHMiuUORhUrcBYrSM+9UJ3oi/0fYDyeu5VmCh55dtrGIdzd79+41
OY+zHdhFASwFi1oIwNWjSlqG0GWeUcomixxwWSBWpQ4AFPUhzmjhcgaJL4qSwnMNK/SXlBe18hee
XGOF/u+MCDtkaHF6PfI7vSZP3xdLUlyVi8q8yhy50PG4+rIkNDOFqtHGxCNoDqWZO0j30YWkFKqo
f1zA4LHaatxfvpLSbDsJbM75v8bdiPMOosMSBOlo7iv1XqOAJrCsxde0eQVXnibnGi7o+6wiFceC
zjYKL3CDuqZphBMbxz3GQif81YVFzwT/4n3ipeFo8sr3HxVXgGsYsiw5LmrWzwrdMUL0FzKgnBYK
EAq1tp8f0LQnGicCOWOtGUHfzjw+REYw4Yg7QgeQB2soUId+BOclCpv8QPTk2hrIAZOZjyvd2Ttj
ydY3TrvCrg2VDA2ebXkW0n9cVx+U67ta2NX+C/miiBT+SCJhCf0RsnLeC6Fb2OFGLzrLQ26543e2
Ntm1WLFPufVAUbRC82+5Bzvhuv5/iV4cMM9hR7LRwPtC5VgSbNds69gjoSiol9wVY+aANJkJHHnk
vFJAxNTONmO1v1FkYVMnh/e/HTgFx5Lvwt7qOZYBBGx4e/mqwvB8KxfOJ2FfOCCCiEECYqwpscTr
JnD3CGD+8RTecopGL2MvQvhm1w+RBCALhZAw1nvb/BlBgDQXUGqZDpxqiofNkyqoXiFgeqOQBHJ9
bmvbtIpDNMm49jQlKIRoLsd6cfnfGGKZZ5TzAuTpDkY0UaVDxaYWRN1tiy5EH/8g5yH2QN2tWd0G
Ofgyetpel8+mHzeVu6Vu0aiDaUJVBQvamSGrCN/Kgd6kSqt2TYPe/A6Zznk/bD5vMqq8mM1j+/iq
dDLT8dURYyXLomBsaNaHpoLEmFWBhloK5VKOWZOnRynrJyvvNCw34eF4nZnZzGCBlge+lmc8p0Po
JQtS4vr3bdkKov+Dp3+O254XkCLSpTTYM0zIrgjZ2gG3yb4Zr/5DNbBsuQpS2Pxkg9Zk94np5qzg
CU4hnLehrusg2O4YWW2JEQI+jVMMI9BUQW8D/IbaWNfpk8zZ8l0teiHt4u9/8pK8XhvGgvzPVqkR
hm7EUTqHNfhKkrV/hpzhs1T716NwwDLn3bZ1cdaL2qyEjov5VhxzfkOFAuaTS+IRfgEP7wVHKjA+
4IiBAdazky1l46SVwT4Tcyib49sxBhKlP72I05fXOEQEwal01JODmp2JYgAydheQwS8wWB9LlOeL
PbQ/9nzvzOxD4SrP66A400srpAZGC4AH/sCC/Hu/LVstzCLwD4gMriPT+bC9aQmUzQeNcrvNLhhi
Vk5Ky5N6FTq+SPj8QyFZHnpQPLfTgyf9uVcmrlh4z1LqK2reEfVWTIe4LjoizIH0ODTZtG+MHGwM
r+pmb8SIYI8AfJq7iI1gMIq/lgLvv9T+QY2kiME1l8xzq3YH3+86CdWDTcpNYCHllq/yzQVVks1r
aKpS8f1OZpO3uUfDFzFLqa/8HkVU4dD6qZYgYIs0iV9hYpkjKkMhlZw5So5Bm5JlPXR9K2UA1mji
NJD+LcWU2k3r4AbgTyWxJW9Un9HDWxHMQZgMCfyWGf0Tpdz3YUpDLpLo4wGsUDSDxcbC0sXDVFrk
FPwN0f4rJzGE5ejkIpa+k+cFHeSfN8xOQBIyRLpV7O9F6NNZmilcJaKuXD/Y97nMDgVZU6WzXDZu
RtrIvzDLJXOmi/zM83EVAeb8dlkNBdfbB7GR9IxqTwq+OhObw1qEJw5A5YDAlz//bdm8QGXrfHk3
iStJeKypyN0riWodJmBRVxrGM+8KTmdTc1j3Ni8Av7wHlMwso6mV54a2v3g7Wj8mTVETZsH9bBeG
KNxkkA/c1IgAipTUJ716E8OdKBuZgtOxMZprCHeImlYMA4Ldc0lpUmIaeOnBLWNWWy1VPf2WW/K/
pnemq6+sanpXQfKDu9usPwISYRKqjWwo8B6fT3VIO4xZ5GDn7n+JqF41GOrrfGmv1H5WSbzeyYjd
vf5NDM2kIX+HZzRocUtaTMFVWZ9AXO5DmpNo6uLUGTATBUoiDAxzOxecaJB16gThgNkUIHDuqBPV
kc1jABI2Au9/hNuuSADMgG0qz/WpOydxxIka5/AiEYL9E8wUY6gXevQx1GLvURDph5QvoC4crdny
1DwS0NCtg+5o6aVkQi85UuQsOLDH7Axy+6Sxsd2vcfMxZQlDZ4RRjqqzFDTJe+y/6DIY9GcxN0oC
FJ8Mvnt9Yp1PsrmpkljXsmuhLoeIv7EHeEWQhPouyueSpEcFOj3QSqTzy7xIyqg7HnebNhSVdN01
JX9jTd9FxYx5/DpHmapi9aAiaRMs8Mg9Gkqe5CZ0c+OEjAsiUxFVKuy1s4dkwaRkTkOFicNaUb3u
hQ7xn6YNngmusFzAZe3nMzOOCjatfrzLkDIOasBqF1mtXxcPVXefo3vhakFoQT38jLb5jbt3b8Px
FNAxcCvhq+Ep7rFvMoUz10faMbeiIilOha/BGqq2bqIUKlI2mX2mI3pjVtKPL2nI6hq2IVDlS0NT
HZNtGj98KIq+9DtXCL3yF6xktXvKrxX7qOYZlEhckae0ebPnNz0QEjv6F01cOTVzfJz85yqQNpMw
+/aaDQSyhK29v/LBn4C3PwDKP1ORQqJKDm+0Euergrw0rdND8BUw4XNy6ESkYUqI1OwuWFrNn73O
6EC2Nx0ubY3Lr+liTPq5g9sNN9PLEoXXCnPcvrgHdPWJmEzzwDptLl3YJdvteN9Sis1E797i5ZMY
SqrZdPrsCs9uqYE40BiKO3K0I2rkpYELrdseP5BVsKqwAcB+Ced67//F0F/XLyyoJxY5ASHO4e5N
cA7FZnIy6G1BIj2+WRL871rryv5C6klN2hqMZSsPpU3kvPoF3iLGlzXK4tshvs57kKyQQMG5J1NS
0pKouf1tAMiGisi/7jaCtPgG8t8mr6iNzOPNR2T3zbiR2i7aeJWF0tRz+id7tQTwLhdWVLgwOUjI
M8FarSoL4lwSB1mOd8J4sep7o9dRnBSEscI8NV4osDa/elrt8PwGkKuwDMKa7U4D9MkFQ0bF+IwZ
Jus/Ipgcutd/dI2c7x4FD4bSq/kKi6rlttonVea5nnkRDO/dFQMGdUUFXcCxVi29Gym9Nd35LJbZ
IHzNeM+/0kq7wO+u0rANlugZKw2Yru72Mafg55et+DpmAQR39JQkaq62waxbsULABWEkwm/kTz9O
Lj40ho5xcr8V+pMdiGwMlCowBqZWrjpW2+Bz62yCbZCCZg9pPojzJ+aufpE4wbGU3Fwli94WBo1s
ao/RY4s7OWkTWZ54p8aUAA5W1CVaczlxDA/EsXHmSlNQJYL26f9LSav4xQj9fwWKHuKjK+hIfKA7
A05YrpFzlQHIvhAf3XLqUNw+BFRxR5Q/ZT8pZ/FgWLSOEu/lq70EOO0Oa6iLTDNXpg72kU2wKDS+
PPaR2b7kddNe3ZBzkY1LGG5P0F+vccdBxmZ/njq1HkchvAZ0Z3rfw1oZmB8uOqTxxTSpVH+UoRuN
Yd4Lyjsr1w7KqCJriIWbNgmt5uuB6uBsBZ0pjsCU6Oq4TOmLKMeqLw77S8jq+5jbQBfW0ZvV35XD
R9uSqLGTjU7O380OUhUd5uPxSAL9ykzqOx46z+xvZ6ryVuHbLZb+hXWQN0YdigSNNXpaiD7yAk6Z
cG+aSIIFrn6Jv+KWAr1JV1mTdEb2ol/cKkgZfkCtgiQn47hNqXL6aV1qBfNZDADj+Zh3nEbw8say
xZ0QF9rTq2MPCmTHp320njx7gFl6HaiaW8c+jQExbARhjNpkn/MiP5JJnbPCYoK69HcQT+/LC0Dn
L9HUizon4nAAL1t7w+OMW0YyDj4x0FRHIWL0Vm+AYimBwhYwPoiQKvURFF5j8wDwuAIWRvCLTEoX
eHWR3A7KLYftL2AjCyqQW88Eu2BrOAW2Bfnzicutvnk7ovPsAzvFqgL7xTAuln8UQpwxtvw+4Tg1
UIEJI3+eiVlBtUF7+NVvc/C54JSKaQai/cjsqyLHIJTso6X48hacjwToTzoLupsomBZO7i8Ppo+2
GtKI/zuV2GwLZK4ebHXb+zLCTKEwryidfXyqipIClcqUZ/L8YFfmEpxPtM9pWGMp6NiQ1P7RtU++
3e+Ik3lK+e1Pn3krbKu11eXwzRH0ZcJApLgCIv1W7+RYF7z/L3koPV4+mtvm32DT2JhDA5pSf4MD
EUNnGn8j/unH/wp7omW8TlSm43qm+UtTYm2jZPhuUzYg1GF+0E2DhdD9y+9PHKR7J45LhyKXPqq9
HC2D1z4XQCj65uYPYGOr30iKpyzifNQFSpkpKVReWRD9CyHXHdSBfQtK4iBoBBcdNjnDfT9qAOFE
FGRiun8oAG4kuzPMTXet+uSaMJnN6isrWBWWyeQxm0AVZaChdTCP9ApWzjn+HWWTDqWjL5k5SXHe
BDodgdr1YHDCnInZNmbHY+X6KgL0OKJ5Pb/2HF5lz8UEePLlaLzgqcWB7yIXIlbFFaKsTUm6CX43
EINkV6tSPeIbSSVcfZgRPBhjEsa0M90X9tw1S2OZ7xsSixFXqaeJiYwskxWZy/GGV6k1vDnucvI4
+rsTNsgVKSo57TB1EnqHKoWnrrl6zvO1PO3xKBzzFqxC8mbLMBJ4ZaIMNcenbJznXRo4dxcNXxiI
cTBYe+nzIIDJ+m+VV4vM9K5yjQMe6tSWNRBTJSOUP8Spbo2r4DadLyko0HwDRCcmqKMrzqA17GNv
Ua3MTderZO4gezQNy7t5xgKctE2OzON42lOR+siU+cL9VnEM6trG0EC9nr8UVUWeStyphkYuPiAt
XIh819D0iIuuzTyWjeZiMNl/qunYE2XpvgLG5PVLvlNZCCILYu99+GxXbLjs08c7+8agee/9kfWg
EpcoRrPHHOCCb1SQ+1IJbfFief2sYUScTMro9c/HxRWeqXzdzOxxfGEFrnfaGcgEqCsu8KeiM61N
mJnyI0cJEp4MiV9llhRoYeEJRq/A+6ESHdbs9B9HnhwPGhJ7A3pD3asYYiZOIdDht76mgk0QbbOV
7w8xywjhZky8VUOg4SBLgPk1aTw/BMsaZ/IRTesLnl06YYkZBvfFI67dWFdIVzAK7Smb9CKvOg8S
oyGjkPDgh6s6tnBJ9j7gwNZI0vCgsfzKdQHywPZkXBc+H7CbyZUI4GTGI3gb0aoe3rx+/+SKAOJ2
LpXTuIQe9w8/kk7VSDUJOP2zvdHdoansKGQBjBjuef8WZIERq3ThR546BGo3tLSvEFSVYG6oSnlQ
udk1n0VdCvGuVMg0N1kdOC/8JiHkrORGvvLSff201yqoP9RhvdxlqgQE8IcQfZzUSRabizGvw+AK
t0AIQ7bh9MJT4eFYnhV1zdBGFiXBcIy7WBtZXJFp/F2NWQdf3CgAaTf17Qd+sQ+DPaIbP2iU7uE/
MPJj2QB2EJw9pA/QzLhv36RM0ieaZ9/THlaI6zQixO+s20AqJqI7clDWHZT7uGTX4M7lqbCmBm+u
+z12EUoRqA+HQ7SVw32PLoWete98a5OigrASmEH2j6ZDNdSox17AJD5w/l6t+1iczvLIxLpHv2S6
Uo6lktuivIB/wpHwCxGr8auRyT5pXSkfE6ZDYLXCibIkaMrWjGQffEL/iOa9X7iIVMW3KZ9BfE3J
jb43nGj7GJ48a0CxQlqRP687w7+tqNCpXsD1VaJae2sVE5JW39frl0bsdBjkkZGOO7ubuBjF14Cl
UFC1eX671zDF0rM6ckQitQ0h9fst9xTACLlFrobztKhDI7q3AVbnw5ikqa6T4KMGf9eOoA1OunwP
SgvQclK/JnTICnoqPLYvPKluriMBD3dphrdER867kk2DByrpvvOlpSDdC0b3HlrC2K0h3lqUVpZx
qY1Q9VrZJAefilQuu/lEllEzNKMxXz2eh5ctM//VfAEImBO9FPBT8GUITm9jQoSWoJVRGvgeVn3N
gx4xzdEoWXM2BksS5Tm4CHmh9k+2pIcc0NrQnulv/MAUfXeSiWPz+7yyrViuKQMvRN4ozavOUDC7
nDgHIU/vFEFYYD61IIy0YBw5zGqxYOUwSAesR6P2ApM9Z7K9aFvnJJrni1NNGNcrNRw3YsSjAwt6
gb1m01yAOPc25YaNCYv1U72mnJoJLUD7JGndNYsAMnvqlMP6S6phpgfat5LmB2Tk4j+e7Q/vS8EI
KDOeEjIJIFG96iUiqIxTv3L8Eo6NoIRwJjG5CsQ3NxVDor+VO84LH7lt72vRDrNgCXPnF4Ymdrcp
42Gh7s5/RW+7at9R+hxJa1qhaUPQvY0DAxqe5HhEVgdQ63Eb3T97ZyNTgwAltOXBNOj4HYX4nbwQ
uGoyIGIxKh2gI550i0CPz/tF2iRdVN6+zWjSQ/nK+5xhuiJO8QZP/uDJ6QrW96vTNfR83SjazqAs
QgT87l8pugVzBhhTbmdz1CP0ykHHtCg6a/nvjEJiWqvZuPPaOzW8ETaCyEpZmcS7tPsMdSa8IJhy
/aXdwwTb8Xtcd1l0z4FLCXbOcHP2Ll9sUWaiYaXqjjOXIvCIVyT506PCKw9W/t+kQZcESHDjMHPD
JVFue5uWziGyeEWROIYKKLSaLPJGYutlKtgkJOjws5CSNV+5WLYGOhDlEFPWrD92uNlez+TZWszd
cuIVI3XGpb3xJD2lUzlBtjm6xH5xenGKZ+wrKR/iPPA1UBdY5WRtJdNnxSnu2/iYu5sWXVNeExYU
CQuDYlOkZeoNUwYcHoEfGdpGAmYeyxUvot2XtO7Z81vZXOpS1ifBxq09LwP84byvdzDowy91GUFy
pG1NiOuvrPSzGWET2HtL8BoRrfH/BZSqiDdjwJsoGmaaNhcACtbQLuqMS6NzyaZ2oTgKZtesMT76
llTzSSd1KotcGYnQx3Thr9Bu2yxfMG/3wJuTLnhD7Tt5fpJPpD5o/PjOXGDDO35/12taB/7tNgKj
kwXVuP1G3jDeCCCH45BcpORWJ+iyrS8A/My3oyABT25idQByGrzhR+B8K6yQ/vTmkbXswbliBGgo
U7W4wr5K0K3bpmnPzp+KgPEB1+/9JbYjY4J0h2WXkLLu164eMfY8it73BbnYVVmJwZFgvg6LqdLR
fbuPvU7lKlxsiXBmJAnoYmasip79vjbO3bXguWpWaReVuTGIlfQO/puZqk8zBR2JZg9uYNKoSLjz
ZerhqPURTk+Q6ZAvIR4kmtN5Ed1KsH/9so+NkIF1QpZ18TwfsLXqXSA5pc+iI65P1JhOgunew3V7
7h/2tb8so5lECBvB8eedjJ46qHBds3QKzGM8YgkKR+WEJPFAFAvdr5ZzN7ZEAy0fJj3S/NinOqmw
30mMo/0wx+SrpR5NW/yQAieVMecek3JmxWolZ35wCTbp6DlYnyV9gWOu/LpwoeYli6IVNEbYotU1
0Kwg+nq0FcJYTJkSILUAwB1BrRfJaX6wt4uCh8X/2F8CxHvcMUTcXh5mEn2HcarUg75TjDUhyGci
RR7opRYIcsmWNJbc5740SVHDmIUqhqUmbIHJOUbH6qcVzjCdwSUVaB44X8qXmzfVIRCbVye7lWPD
Y/vgIQCGH1MVGh6eDguJyV1fr7YkkRTmyy1oWdFKE++UuBp4wgoxO96BvVsWqzum7LFOo0zM52sG
Ma60y3SSNwTsLrPrHyciiEXsPN67pxFHmtWz05o4QgQ9/dQ1AKA7HJmN2ABAXmNyhKQHlcrX8FHD
oDcuDhLYqp2Ca/zNzBBnruS6qDOeE8FWgNbvPGRv+sG4D0tNyShcOszGXpKaIkB6Q9JK9Xt/x5oa
R38846Kc67pIUVhOB6rzf0YKJc9gJRg3yZJJF2u4jbV9RTOrAfN1uMU0ifA2R4DdlZHpPTmnIppy
6gjgrgz5fgou6sJeV+itSBksKCwzHcC0B/U2mcuxGtr7/fobcZlhFMsBqviB593/K/XZkzefgaQy
8r+wSowyJCq92+LgdTT3QfTZZUkG4D/aXOXtzvWBxjQmHiWnXeN6hnxnFR63+eQ8PnQpXfZ2d6GC
UzDrQY9qdq3ub72ckcsUaKvvtw3d4SY/uv8L4r7yuNbzyt7mf6LCZJvi0jOoG7N27jkZO15R6kl2
eIb1+tc5bz1ZAsUfC9pBJTr2rPofYoFvvNytJJHl/ZVdCJr6NcieIByfkWBbA0jWT+ZBO/htV26O
qEJbctVYnBlGYksL8D8i58E99O3R6TouEzMchBc/PhgnZtBoHWxbsgh/kyeBhi0eryY955OiOm9T
dSs4sxlpYn0gWKPUn6WBXp1P/hKwVwaOGiT+rhmUcSNBtiTHYret0FQ5OoEP7rfh3eDMWW39Pto7
7nLnVVYqr2Ozau2PdScg7TxE2HxiZijTVqwO2ET785fWqa/Yt8tuIdTF7Evoox4edWO6envpWDGH
LZphODchyA03Nfh3k475JqG8X7ELszjFHcai81evxUXcotwidyakrcv8FAWwC+wHlHr84We/wjZX
CeyDu8I2DXwrrZtAxx4UZ0migpAg4gBF0dWQb696+Dn7A35qOb+VYe55VaIMnPyd+uV2wJeqAMCm
3ifIbWyLywfiVT3B/fYkLLeWIT8BhgQF/Pb/25I/PGaWA0RaM6khlPSAEqwcg3jZtDyo9suR0uac
r2Xv4ugkC8HinYl+z2wydcYH7HuUiAjaq2oNrwqUTlOF7UoqHiMKOMdFCv8QymDDe02jx9/de5gn
aAMB2JHk1NYyb7pp3TvDdetAS0WvopQWvPyhrzwJioGTniP2gXozGDhZTouQWWGarjMOjgnVdpyK
6rAY2rK19T5aULrfFgJCJCougca6EvrPAOtEgwgwZF9ReuRiqijt3FJJtjUsjteaegwnT86xsXRz
Y6ZcrAjXtW7eYiCYg3ct3Vxq4YIrSqX7PS5zjt0kyynNdswexbu3zuNLtLv3/2IcizLf7tJzb3oo
G08gxwqYVxLZK8H84CRwGY+P1A/y0wazp1ksRJZHwuP/WpbP1+j8rDe367iKiFTz0h+iipdFJ+vj
yfrJlXpt7jhAtiwNkPc5wEkZvE3PzwT1kSVca3YOd9yjQzJxOOt6kdMok/bBElOV8SS8ygn5Ap4O
CbZEk/Iz/bpaxenahnaVqPnVwE6tz1IQE+2grLB033YKvdGcK1uyVSkfkTqS02RpwOkH2ahJy5rS
/NrjRTUu657SQwy9CxFnquIH9mu7e/zAJmlbed2hWCBoxZ5Jm7/N1RYMFQr8x6xE0dJDzMqbyE8Q
TJQBj9EtSERP4sDgkBWs5Iv27jmhOceu2KR4Dk864ESsM5z0StHl5mPIUYoTLTpM51N3dKy4gt+g
6iQQNUsuqF7hN2EVSz7lS/HUx3vJhaVcrqiENBhuFvB6A2VUNF0yX9LbPfP4RrBu5IZP0G5cKhmg
x7+yE3nTzG7n8IUQfiZUmySFriXQqOhfVDLDyAqWhDKbjQjIE1qH6N0MTpomlgrXvAw3Cs6tvtcG
/UqBBh+oy508WNe8tG0iSpkS1AU3VGNJnm1wW/xqjRHA1f6tQEJrPBewCuc/
`protect end_protected
