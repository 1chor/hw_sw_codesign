-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ha2JkmZwXrcIuoDsn7zyWXOCPI4ytcU1Nzrz40hpkcxtTBNUkOEBgQ7ikuGqH86t
3jtrBNDQ2FHIQhXpgtrtd5YZVn1OdzgMzuo1TrR5d0pRvqitgkanMsHDLXuDlOkb
vzBFG4Tp8CXmGmvns+7wfHk9+DteLOiJtzuov+dd0L66tqvIPWqlsA==
--pragma protect end_key_block
--pragma protect digest_block
n4Z7VRvIRcosnSVTbp1QwH/SHkI=
--pragma protect end_digest_block
--pragma protect data_block
HDpuyKaMh9L9DgggV0SjOhNTa9jsFbjBpW/6wo/OoBLauB1h7pcmNG7PP3GTzrLj
xy98y5niVrj6OGAa4/RXvJt/k0tEiCWPyrLfpsiDkDgKjja1JOi2YZ0YXLJh+YlT
U8c1ROflWTYFJNgpvilzd5ry++1S2o7MsxGquQh/o5+qJW3Pg0fCCd9mPEnZW1sJ
8Wfd+uZb2XfzwDlU3lC1cMiyt4lHwQJL7euLMUAZPeLnueNnQT9TGVhCBLhu6MKl
ixDbHGr+muQWL1pKznY7SIWDhZXmJIRdHP0k6Jb2eNIQvIFvGBr6/jXdSQgqqLeF
NGRIsBrUgf8H0dgiapP+6eNW76sMJPtML2dqvOn3tSUCTn5MSKQEFwAd68BFbX2p
h+vVDVc2HgUL28/G0VI3JcaVhjhuf+vLyq71ivpUi+kxsvQplaXWjxIW+KkWc7er
nNd7FWBdV0nWHjfiXdD0EMDQCEfRlw9BqZ5pzUPwUtSMtmFDI9sNLmHlhhX22uEM
Hz5cdZfMeTpjunQ5/BmYNGCIL7ReOOxGzJA0UvKzBYWFQDU1WBfyzVI+o6eUAyfS
dmgz4j9meuIeYdn9iHjvngo8/qZf9XZz0qpLyvzvCd/73lN5n82FkU29ZdMpy2Gm
JxGbt1p3QfSfVGYCJa5iMJw97fNfwD/KPtuWYZxos3u/GKGW2Nwg51SCi/pMl18P
ppJZy5riE+M3O8D6ISLv8uULpi9813L0d+V+JbdymtYIlSgM5kYRzIVS8PF/TwoO
6c5tTk3rOza0PSPdtFjeXdPn2PmqpKOIIfxDdETI2HCv9UEWmhts1B7pzLoSspm1
dnnyvudVHfPY8BO9foy8XA1TjWJepIBxQApPE4dCmYSWUhbGrC4zeo6HOqYm6FWc
3oxzc6OB90F5OTOR9I/4dROUg7omu+TDBHwYRbaL8gabL8VH1jJOyWzjAhZi0Hl0
MP2o73UlGg2QBHNCHJYf3FuF5OUjjFbXAWxKMSN7w4Rwq2VNvfxPHwQPA4Nt/wSa
ixEF02it3vLv5+3cJGz9p7Yb+3DR3pvD5NlKQx1LpBvPPtSPMz8bOaXTFcxBgadu
A6DnslelG52eRRSR4LngHP64cnhKo/1sjKMEj+nqFuveYQsT37I+aDrADNpS6Js3
9WGAy6T6KO4/ihTYzeiPVYJJVodOqWBYQDe3jetggKQ+tx6rdw/CNO92cPJEeFz+
4nvKfKPhaP+kikOeMoioK9gjJcLcHNO1OxcC6flkLFXCgv7ErfcpzaOH2AxxBojI
YH5hMEdSh/8Isu3gwe8mcydSMQ9D32kH9MSCz2N2l4gEb/Z8ZCTuMWt02H82WwZo
9t9BdWZqjS3DYbb798lmf/bkbYbcHldjP6XzF2oQ9tGhtTkKAm0DmCP/qe59lyPv
ebZI4gukXDpHp3Wt+ffjphhMVF5D1NDhwH/YsmIkUo/PqEvRxnhCj8jymXR+NRih
MItpfUl8M6QHkgewxSC6zWqm8IAsSHsV1Z06eynDz9RH03A/uwBoYvdUIhGr6uFP
mzp87VhEMx8bVvvQT/BiKpgifhmuo7ZC+7ZW7dHirjN586zYCy8OXYFYAZg8YMrY
VK+5f/Spi3dBXnnposgrPj3nH/HVnMPhVHnCi07ZOr2DWuuKOMqTPU8E1MfRVYQb
QTuU8WWesZqOA5ShhIl29gwCixXbbQZW/KpKNVUTw/Jyy5Vqb+UF+jZcWBcDj6m8
UgcRs44kyQJGtHt6rrMWyl4933qe/NcGGT6HPLe+WsFnnUQCufmtxPCzbRHUp+Ri
0mGi6vaBnZGe/ETa7N0dfiHQdgGujuFSQTWOQfDFjHlhy7E6W51JvjLroUly/RUh
WsDABcuS5RCnL8Q/U9RZ8uGw4yW5pexefBanOIo/GtAj+f6LucXgpsryfk5aSL7x
yHsMGenZabIvMcj1fCbRyuS/zYZVbGztkiyDzZCRBOQBERkEWLtT8TEzLdsMT+eC
Z1nCJnPBTXEXUbyxKtQz1SGoT2hatGY3IqyEUpwVnoyrHw+m5kgULQHPDW1RbZSC
vFyZPYrSkGZtk7wULSQ7YUh7hLkmhYcvVFoCOCOS7r3nEgJKveVqyS8TpZw2O3Jv
T/DXE2sjL3kQucDizcDqtwdzpq3pduJDGkflj974JuP5mRduaaB+gjR00BDQ5OSg
xA5i0vPklaCpbRYUuutT50Wg13cX97KEmzOCjMwExfNQQpdFGa9HdZIXnCX/1u0r
QmKJJ5sxL/oQrEeRtrQj2XitsO8KUXnfQowdcgwXRozW+9DSdCcD6Q0VzKhL1RXb
Ll12nMS1KNgOgVBkhgHOdo8cDPkFMxZJVy3uDY7eawxqUdYb8kFBmydho/NooySr
y6BIk7LDFVb2iUpNabU7RFDpc1EhtMFS7rb1mCHjQjV3yAZZXdJK5u9uHZ+TR69g
0M/N0CUu/4GNQwy2dhv9/a9zXYtncTIk8gADh//PRry4Tlth9UnWtu70MdGt1BSM
SHs6v+IA9dHEdHdI61X7EDLSbFqp5RqjziUSrccxdBN2y0SL32m8cme4y9Y7c4Bx
p9tIXPFkCsQn1q7iRT3uOSLRwVSG6hpeBMzImgbG/fOShErSZlV9CkHGcZNvn4M5
uYUBIMSND35yVait7sLrnzNPJ0piq8JIvb67oOp11h6TV3HI/UDdkwoddA57QHWo
MPr0XBB71SpLJZEX8/0Pdxr4amWzzABm/D/Wrhuuzh6dG6zj0wr+GZgqFP1r8d4Q
09KUl1iKjsAB9HJqpGMGaUse9KmFMMJnZvtFdpm/xS8AJFAO5ZNkzZ4bGbwrhpDO
IZlJdoFqApKQ2Z444AJj2RUnRusNLcsKb9hfxLHdOONLFxCYqmj0AJ5V9IO/JhcO
Qa8heEx2zRTudYsYAvCA3OypsEw/eGIOknFZsNgrrSzGmK48qJg32aZpg2YrItJm
Cc7SeO6jB6OwomnGNme2rJKrPYgKd4gj13qmW/IMMlF/4W+5PCR+Cn5Li1MNQEGj
0cxqfI7EcngDf3dZOkyoRTk4HJUjgHSwuYbXDzDH91W2IBmFC0aZK4XhlYIqqoD+
nAbf6EIUwDWn+YquS/sfjM6nVgbS0NrEtpVT/DOy/6VbXjNXFWA5t2KquGMeVnmp
ZBjoNT54MrgekYg4GN/d+3TN0vinVTOmtwZtev4M0iNz7KQIIv6Sxc7H14JcDLMk
imXqEeFOj/4f0e7tkI0kgd9Y5o49rutnVkR/FyTNBHCpBA/4EWV7Dx+yQNXhu0rU
ePa2uzVTiTQPYnxwh+z212gx0WKV7B2f6q8rn5PmmITZPnwOx6vXqYR0H2NbBblp
2AGwoGJZu6H8i4A+yPQS6ceqO7ZprGt9arHhk/uQGPwENVzQ7g2ZHnu5o14ifDxp
l064IPbbgIQTdnCP+wzXdllY/R1ytnyBa6zlPDyQRhqU7Y7z49FL8U2UwibawQ+f
zzyA4e8BcShnfVDLLZDoDhbPEakbAx/sRLlUIqgO7dbkYTM1HF1hqWA/31MVbRLC
MYQhxqLoiMEn3qdjI81lBQvHDj2FledfK3qW4Dthr713Ws5aVaLxuoKPENfi5Y/R
/oxy8ivesHAho9qFlgzFZt/F7k3Bb2HDntIayMCQAfIDUBfKRr2DlaVghMDc5Db/
btxTBlRew0t8Vm1DYwV3hXip+nr4bXD/DR+o+eYOLcgHpo69ez2tTcI7PlY1ZOBB
FtbikmK1tlTuHod+R0uJY+UNoCyeP92VDV0zaV53sxtGa9w1mLNbn5rHVAPHB+tp
J5SXjordmc8V78O5eGBiCX6GoePdrtqxyLii+u8sdql/ABpFk8Vn4gN6mpPARvvu
dKkOqO0kuim8YhNXIpDHJBWuNS3xyJPd1pwpxKv7DkJ2sQ4kNJ6dVLULcPqJbQ6e
KyZUGJS9yYA1fyta7nBvv+PjQcvvdujmJ1FIcnWB3owzCGznKuekMag0xar3AMKJ
UHdAAUlNPdc/FUgC97QAfHNLOZ7cYAU9MiqyJW5F7+KXI7e9x20YDLS/B645moU2
FcOkJ4mb/TV1wtTFaOX63YyJ+3RCQ6Q60lKs9YyihuMPd/rxgUZ3noAnyLsxC/+z
Ytt8dMRvhk0B8QlC1M+ZxCzSxtdSQLQRGZ52OkL+XTIT3EnvidAOvdDzyksWj0Bm
aeiZ7wqZNBeHAnrsQom+GpHOviRth3tQsKbqd572GeaqrY8Bi4EddfOwuD5CPM5J
BD78gcBnG/VZlEuZdHg0I8UWOrs5WigrGDENkxCv25NawpXsrDByJlUn/wM2tMpl
Mvpknq4NtCI5/OtQmKblJ+SSutyGH77qndjfWSQEF040aAhKZHYykN3NSWsIP78B
3gMdDvv0GoR8YaTJizeU5AXBx0NRTLxWaopocFvII7XNDllgL617UJiFK9of3iZv
7xlKdb9XKjHun5C4PIKXaWA8Z8A+FgPH00G5tzSj7jokWL9RzGuZW6hs4KBVBqKW
1AHyn1ow9vhRL35LJLgB7W5oN87Prj2VZtWipfOnWVWFWz8yFL5R6H/lJ+IG8S0q
YpieIFvkJJbWrVMWeybb7dAIWsm+T//fejqZCTTlinvXxA04lWE83JYHUepIHgiu
Hg48zZ/KLEusDwfOWJOcwl7jOtll43KxRzZEkREBfY9t2WF23L+5q/tTIvE01KyK
ys+rUdBpdnIcw//ykq1Ba6aTbsirUseLHJFPyd68+8s2KRV9ixxYHx03IJUCauOA
axKq4J8GhRjcgXuaGfYq+jUQQyXc08SVMqxqb+7mcMLYPvnofp5LOzGjWW1+/UTE
e2E/IHj+mvW3CnJALkNDNPJQcgUImLR9Bsw2+FPzLGuobgO4g7vTePLi/mRqWDFE
8HpCrKdtpkxcVQJZ4frz5waQewYocx0jBpauxVgrjyaLV2ewNv6oL0O7JnSgmLa5
zrZ14ZrS5+P/8PtCHQjlr9LKmkIyAPfRHS0lEEpiqQWr47dJZkERG6n96NdQQgl6
4qv3Tc4u5JdxpGmtYAEzQlDKz+//vpwq3WABXAidQG52pcufheqcCOgs+9zPV16p
yaBKNzHCz9l9ltwiDvGTNf8uhaT47GFW+QHzHKx9TATlu7O4994dcUVhmaYLFxRP
GeJ/1Ty6FRdzyQc4wimrVYXzDQPaA95BVlCiGO38G4FIi4vymomFw2bFa22bUkb4
zv47iO36OvSAF9fRyc9GIGUFw6ER7scxAPy2EFDlk0vQgH1STzWBJj916ysq0tz1
v4i9tyQbv4FL45g4EdnpZcx8Btl4Xa/7ZMf58+wKtwonACLEhz63UoKeTkxdUMVa
pp6bQwKdE/79DxUFDqNbN4/JJ16/tYBKSD1fgk5PcP283fQxCuJaYaUEh6kZiO5f
4s8lC/aG+duzelCuRruIHN9xlywU/IAFuL3KW8dxK0HZZP5HVTvK51PFwer7WoPr
ub1hR5wgJgnKaUIaQnpa6nbxJh2rDac7U4CndkPRLz1Xuw0booZhZHUO55f0XMeL
+kroTMF1R5dVnQuaIZXklKDvur2ENCBeAc5bqVDSZ44EedxLQa1c8Nb2t7ABec5j
3QZwRfLoeGs01O7GbBve33hM+pYbqFD6Qi/l+TmN2RCoJruhSZ5wMtOZltudZYEa
aSqqx8Jv718LTj0TaCalu6Ql0Q4uLyrI+MaDLTmxsLhM7Fgp8WsY2R8UR1twPUX8
BUZZvgmid+LEfSHyY2US4pcxr8wSVrYoPtg+/PjFZgFABxPOzECew5I2YBizv2CB
sHFq6oVQlJvBkbDQO5Xr8QE8tKc9xZUvihBTV29zs984gQ2ST61YP3brfujXNJ+6
VLSb3t++0q+B4KZLNYE+EQACF8sooZGvEEliIHp9eTj80MQ2jrmm0KYCmUABkeyb
ttRBrZO7EXf5bOlun459sAkYlQ3zDaLPiA18qS+Q0pjdlTuDKA1vi5evvmlcDU3S
i35oxMqgDSXzdpLN+bVlVb4aaoERdYq5nZ//YjDr+K7lqrHYUP1BLw2PDAjemc6x
zUs7+kAED6pQIlvbsA80yIay8vny598yEMkBbx058r3rNPsBzonBHtDykNj4zblF
J13vnbZupESGlBio+dHGbaTpQHfNKLVK61ArhqG7jJawLzD45lIS4uDO1wi2sL4B
5OkLHOG+5R91coEfyy+orXf3xcfI+iBI76L82h7kJrgtUPjBeemSTNrksxqwWvu8
6cEzm9PixLEJrFvdDhq3b0t16mnx3G1+oFbCFUeNEOb0FAekQrR1wcz4HcFGF3B6
/ccoYA0G1RMKvPNNCQtUPQw4DL5NUAbdUPakl5smNkTA2fKN1OfUln+bL8v0Uy69
I8l5TPCkDmAV4T7N+ue5So1ld+ChYc5UlRT4kgk2VfMWxhWETOuIYSoJL4SP8jXU
j4E7BF7XJlHUaCvQsB0dJsFxn+rW1gMBe5hlT2MA/JMm82Rz5c4VjcjC8USK5eI3
I+g8csw7Tzy1KABWBgNagVpRs1Vg7B570TgbmYpqGxxwtzRIZGPTqemuakfkk69q
e5oSG55L7Zpo2pADExPEOzbMs8Si0VaU4PAmcnq6JZ8ir3y1jrvGuY4fnt63ycdD
ziMpqMEWJemS1ZlV4l3VmDOwo9ff8Jr9wwae1TqoFyzNRZ/9iii1C2a7UoZsJfMl
yZIwkuftMtDPOIDkn+CV43kh4xQXJ3Jb79nKWnduzL6nbaaEhEy9P0UvGjhnAKcH
U6oL4isrOU1gIlN6WA5w4H3P8dz9/TwWc0eb5INj5T5oK3MDwquNosLvKtSBEOo5
LdnzCCG4O32Mxc2y6LCzKHTSu5kgT0lK5C96AOghIPR7GygnFVexkGJl3pT0Vl/u
jlQrx57koGBkVziQqPvST9HNUthGHOpqHffeMIBoI3KrSzZqmy+BwA74DhSVwNHo
n6tpi7HpLulI1yUeytFw1yYRsgeLD9ygB1B/dPH96c7qvSgkM46tgEcKiVc0vATG
YXFXwJIm22bYgdbv9FPvNJG+ebYtvZUfQQKnrUX2MHj56IGe9kwrNQIe1E8XAaEi
tU4Ymd4BOmAGcAyF70YMpuN5o4U3gd5hXi9SjY0O2SeRZWuwQKp4nGpX14l7FpqP
VjAKl68ZArCSmAbLKNP3JUM4LR9lx0b2JOk7UJSTR3VjneKvHE+T96pcR6Dwfsg2
Ujer+9CyD25GUWDCCAKDc6aqk6cXV8cCh52FqDChyfcXVs40/EYtNw+H3Ae7Px/F
H78qjcN683wEMAHZFFsEnC1BChspjc5SjLyM2Gods7mUxvvrlALwSfa2sw/qjuSh
JeVcecdKx63I6F/h6evbQskJVJZMm+rIB2tRygvpsGR/5CUp8W1NO83Hl0GCJD/U
MnuOMhvend2B62Y6TA8xEXsnrRPuGhU21s2PAnAZ/eC6/CNT/VGZETO9FX9PGs8p
WMfhxB9jr0MAzSu2QSC+yK78CnoBDmNdrda4CK38FbKFE26tFoMQqyWdQFh5sNvF
LT/SJjERX0UD1wGAR72foBX2V1N9xJvOHMq/ZCkZiati700J27MRMsguN+bqmddM
phN/PZtDMOrV72jYpop0ZzQlCqRNfrz38q74GtiLgoB/+xZBOpyVymliFrBQ+uYg
OYgYdJmp4BLUKwx2SI1kgMl3jUxoaXogBqbZCvkOPieQ/i6h+w86xjGN6VmIv7XM
rKPpDgHhfLHfe5pqBaf3jAEXzTBCzhwucocTtCvgSyZ/aT3tCfigR9EyC9olmz6Z
pCrbS+DGkT/6gsBRHoMqa5N0W7Bam4zYWjlXNy6jCOxXQhLAqCKCX9n/20S/jzPR
yyX5hzuAsi5mpaTnaI0/SnaqRK17+FsxSQj7n5B1lt7kv0kJKbzv5GCJ7YiNs/i6
xw2m7cbzXw0JDg2PO4A18pdOMghdOO+hlI4aND8H44b2iKEfcd4GNGTwz6PZNOBM
6ppCtP8cWu3pPaOew4uzBS35SkUU1EotS57vrkmqVMDI+eR0Hvfx1Plj/xP2LUXr
kbH2wILZJWishYFXm/k1k4oWTkeKtZDvfChfmBKGndshzpGE/k/ra7S0D+U0eCQr
jNV3HfITuAXM/mV4jQjZ8LIz0RTDeyTG01UtHynzp6AcS4n/Kya0MNrhijKIyUz9
7bwlfzhctX+357OdRBiVEpR3khbk7iAYtYp1tKq5MNOIDdPj4tH/Y4QKFb1YeT3f
h3uM6AqzP6UXXh/rvn8gsrArDNzmnp8n4muKAwIImQ1lWLGSTeNCSEx9UldBFvUi
Bc0/8u8bpOCBQrrp1FaioI3zzZIRlybyZMyXLN8qdnNXNgjaKw1+rwZv2tCY7j8O
1Vd3IoHLCDDFkPGMKJTVai48QVyrIm51HGYrJcbcNimUiWkOvO2sHVAWMvWZqiY6
vrCzRn3fVTNxJvf6ddrLhj5UkaJBEHxaZ0Uwpw9h9BcMU8YBo5gttK1r/dkA7/qh
Wx/0TQ03sy8L5aKK9kLdttqfbaGEB337AugZS7vruvOxgIVimDsG0OvJzbGXv3xP
FsuoDsEHf4Hx10kxgEX5CUkrel9CMoEakMVdRKH0CXQVZQSE6fd3WZFsDZ/PnrsS
4uL7HEdaVBWj2tvwfQdBAPHl7kg5LTjz6JsCIDD088A0h/7KkSNhwagXFALhVyyC
nNSFv1xLk/DYxv4j9VDUp/eTrsGNhXAFqwinnSEk5BktHcMeUEt76hpuEc+lFJCE
qc9Bl8GO/OLj5Pwt2vTFbfLZFAIn7yEk3XiHJbkTFaMQlijKUoyXdkc6luupOVRV
K2GfQdg9ZseLemTxxurmg3eocmFmTCW+fp+S+U51Bc8yaswqw+J8O81Cjzk4N4se
WKVMDO0YOdFetkytnCJOlsDdSX2lFPuzqwRyPAMmgGkD5gxAn2krwVN9ARW8WEJf
mFwiYmxcC4vGiwhDO+wgCsVFygLRarULdi68hkIUqkgHGoTLxJ4eOWa2J3R7E8JT
TNW+Wz3kcm73PnSAftwEJQXdm4AhQrisYPxGx1IdqRXQsmHbjDoMUJrG96jsGdio
jswGap0t8D3TlP6KluGN7gDBHsprnF6ZIDIxAAODAGCnA2P/M59kYNxTI1CtGndD
nfy2btWE3N+rauqUVsZk9/hf+KoVnR8bM5qIbIbMkdpP24iqOecs+4KKOJvAlN8D
xm2Yk98Oae2GnKkwQX9XKGAW97m/T7HycBwosqGJxn6aQUmWGu9bC1b7Qjs1+rYe
UGbNXZHTdiP6HMIzYGCq6DRdxgVbs02AxcGj5MC6hJwgOAWURgKtoObCrlHTMUwL
i7ZTHMKMTFrjaS0tBQ4vS6wKuUZS2U94UKCUsDuWDyx/ZhvY894bcHTf+AsEmpNG
wED6f+MNa0iMwOVq65M0w5LdAlNWq0hfBLmoIv3g3weOzWvcshJQVw1/Tloy3lnQ
AE2EpBooS0q88oT9i1u9e8weQDevdXz4K+Nry+kwTt2mmbHzyNtEsl8rMbIQIBnV
M6Wl1l9iqFMxBQ+PFNcjpAvI1q6vySresSCq8D8cbV8OyPQfJM23PSo/aYnr3azE
xVlU5q3hk6+nN1Kf4GNGk2MsBAoBLBQZ56DGRZXEiX6Qf/+FYEfs2/G0/U8tzUMw
gTra0A/9kRPRdP0IOHdNdZvCFAy/NQNARx9z3id6hlAOVWjKeQ7Q33hJaKyH0/la
Pd5ZlivpDsD5VQv/VE1j5wDL9ncN7Fdaqt+FOhnsxgaO4PG7jV2YfgNX77/d1g4u
xnUfH4LDjzH+2/1JF6f/2Rexqh8Q0N3p+j++Vo/YjQKuxiIe9UgcGNLSlhMqiSux
KF8NpmEM0wxTQ95ZSLjO+rr+RVYuGKyJHdAv5LvZjb6Pd92jUOrJYu8FoPkfT+zW
0ws/tATgwEnma/ryTJWZJjaJV17PLRIrRgGDDREW6bcCru7CqbXq6B4abAz1YPdN
7u1TCcqk7VTnrtVX59F3ty1c5/4XSEnvD5QPLkbXlPaFRMMoTETynsMZc/2l+Qp/
eLaaOZ8TvysYQa5jlGlOoLk7Gt4ZvU5TPBunvRDNMWFE0HUqn5F7fakBZQLo7dNA
X0YsxA+EPP4iuawroq0utCuiFcGjUvr8YzBMnIT6qc5WjqeS1U03/3KC0BYP5qLf
6Iru8c94gBUZnmdMUg0LBGQ3g1VXK8DHPbOKyME4qxGbQzH9QmUla3YG3V6mjhyg
+jaolAk2DuDhnE/57zyUfekgTykrO44evUfbQwWmtvumZG+jvcDhcM5o3SAit/WP
Nd8IyR6si6Af8UqqH7c8qFSVd+AO5bznSw0GMt1P2Lqw67QHHItvKodad+3P5fQE
sJme2pJbgH1LwYytsMh53DpkoOTvxITLQHN+YUWqRxM5UQDgGa81iCbv3waK14nF
9OVcoX13HWL+3QhUe4Q4K7nEji4Pl29e43/VZaqf/qX26E6zME5mN7h6NFbavwXY
a6qJV2PnwV1jA2uEGioIIvudl7De1jIf+wK7xze7RIBiIpQSYmMlOpsBiJFRp74G
aslW3X04i1jGSfXDdMcWIf+9GTakKKrN/41kMIV3me3TMatztadxa9lBfmV9NHtY
gKs33nH49zjrzdwMHShnuvKnb8abLVabKunGaLMb487Kw2h0BpMRX68xkAdeXapl
E8oz3rH1fKjaptZ2IEeIYmiNnfPUEAk9zf00p2F9H0RL7QQqNnCFMVYmT+lSyXQq
a7EH5jGdmokuxSAeEs0EMSuKpqigJ1Tjv0cwZs2YBSx/Ztg4GdpjN3M1marZHF89
axldk6Ul3ZoLj0BF+SkuSfWrUeDmOu1XGGTd+53vje81uxOFy0wNwvgho/d3yr4l
dOs3G8yjjiFvRIyJyLAKk8LO/SRWlw2LNiD9beeQRwYHT+w/GErBsZ1diEY/IzaN
CQgSmY6YN/6ZBZcUK5C/A7et9uIbsk74IdycY5YX+S3y0KDpS44Wo3dMBWxZ2v5g
49nUCp0fv/QaxM9n74bids5jLJunn4KaUafxjAKRWzBF5RwBIxCPwQMj/W2hKR0M
hBnTibvCVov99FzPPgsi6B9015NBy5xddAVHaiVEakMARWb5W3oA/K47R6RQwiyp
S1fCewMSl8wlmi8TTJmvm8Lwmii6ysI7l+JhqdNu4V9H7h50f1Bj2pr9wmGyYW0n
VatlZkHex7+XgirN51gtEyCAJbG4QoCvszRvx8hlJdcdt4gRh4KpxsdX9dUqY3S7
dCGnyTPcMp7Nx5iEW5e8XA4T5v0RKHimln+EZuDELUjdAq93cKBjRcpo6XWvsmvq
K05kX/bch4fwlfU+ysEUmNk/GDyQ5Qode5w+79o/le/3UOa0+vWYBipdZQe9rEp8
ZaDfYRBdQR4JoyOOk52WdaS2mCTsa/Byp0atpMlhYCDYsrlVYhS501Cfuk4cWCSo
JbaculjObN7kVLOWGy9U3vsBJEv0/uHqPG+3QjsxOMSSuvmnSn+NpmhIDbWBKjpq
Fl9pOy4OpMOZ57zhjTdxAVnMshHKbbJllpuUuJOnRzYPXWaFSltT4iY6Gt/4zWDp
fcAnyc0zKnAJuyqRf9FCzyBgj0kiTxu+IlSZ9E9DcAVsaT4jaWxBC7NrBpp0R+h8
3suDjucltlRN1ogDuKF6SBN0ZQnSWvTFxubVtxlp0QPDhbMarv/eX+SjlEWmprqs
RPBUxYRaB3c15FAIlN/53NfKCAU8tKJhXtGh6bFoYrEeFeVwc4Gu13J6TqzdloBj
43Ydy8tlmk+nsAdPDnj2JP/ip6fSm6QYbCxP09lRv8syTcuRrOWC+iJYv0Ts9sQd
TiMVO6P2dEpR7W2/yuyTA6NdGK4NrIZNiA6jHZkMpBBhaLPm3OaT3OfEfdZqDzlJ
tVMjeZVcKmAE5sAx4ncxqZsRc65d461Z6jvUJmHy0/oH+3LK2aID4YhB6V6Q3+Uf
o5mbJpSu5p09jSlDn04Sj7wQ6fyCgJ9jLZkuRPQRqgev9RkjOJYzRt18st99ZXwc
OZx+ch+smVZFMgvv2f4ODrqGq1+uz56AqiuFnZc62p2xcY1tQPc3v5Tw0GGxIH4i
lxne166IpH4czbbtCcwtfMuZLGVaWyySIDvd6JrpGWDRFoHLKPlCwRMYyzgFxXlk
Hnth4+39M2MMjZNnJGgvZeYZ2upKjFZnyx3azjKqmF7PUombqIbdi9AydAqeGipZ
0I3hlBr2JGjLVLnec1o5GPGPOOrlUjrBJv+2Agx4jAkHLlXZ5hSd1XdIEFHuOFEn
yw6zV/I4GqfZ4ynnbyg+E4/2vJAzTbYSVQaCbg2AdNGmTvYt0EmTtZW5eJFOuUZH
kx2W0wTLsqlW9Q8aVwZA8nsiJSiYjSV6F+pnMC7fAvwl43e7foivZhynz4TiONyr
lCdw5KIlK0admnaS6QS4hB84Q7U98/yna2YjVrj+zkfcOZwShZ3ochCjHsA3QboU
SFOA6+u6pdk94qsHeDiTm+j72pg3HyaSwKzrYWqPXp1aB8E5cYN7Mcf3eNvaGLkI
uraXe6HJLPsyRJXpGjro9VekTpEjD1HB059YrhONlH54CdOGAdoNMT5YxvE4ub8F
QExFWXwOK/026xkf/mTfJAn+5XTOZnJG/xR5TM0WDjDrc4ZV7AR2FVL+g8Bbl+S6
QRl4baADBpjuyFRTNLNKTXwPsSXeqQfXyD5S1zyihbFs7xlFCDCzIgPIYmPbz/Wg
076sFQeApLgYd4UzT/SfSPjjUXOxqhHgoJi5mX5QvR+mapEG2DrAgf4+FDmuWrvf
ticx09cTr1vzgml2QScITGHeSLOtzPZckehIvS8jlidiWaIA6gdWL9zQdbkDvihD
1zbQODJgkOalHX9vPRo1g4YgJ+xaGl/vw6P4WIv6+Ydsmwy4rN1+JzwuD5XX5pYN
Rd6pC/t9Gbl6yB8wizuB3mtL4mhfMy4Uak4MobsicGlIvDTSBj1Mm0aDbSq2DOER
qKEBTtTwY3PdKhC70zTKYzTd8v2K8T5TrdNAMDfFckO9jmbWPjCKrv53paD0Wk6J
rFbLgBkYfiSjjbpcrUAVy1gI56QmXmhqvV5LhJVHA4vVk9F+OVBConEzKHZMMOjJ
RjXfuB3Jj3h67acIyDjjYEsCCy4yfCDchp2nefDSQT3pUQ0slIxeYuVkCKA5kvP/
/9em7rbwlmslcH36G5s5qivCCJWhcynBG0TJUD4qzV+9gjd55h+r3yOhvzN3s2ta
MbPiUNryWvXla8fXnPxHwI6/GdfH8til/d72a/45Hp2g2zCg9VBUhBhaiAIBKIa7
w2ejTJmqVOm26qgbuEqPSs1WKvgroPf/JTmKqo1xScmFCI4AjSpFj6/dZyE6XAMQ
UUeAv1LgEppDqaQP4RVEZhF7pSfsIFyxfdYmfvf+Zdfjd44kQ37oY2QglHjlYCy7
NXn9ttP+czjjJ7ml1jHJKw+xNzno3Gs85uL9keJKZSnBq3w1ymn0fM/jtzZB17sE
M/8BsPy5qY9wa1/6STf5fQ+iKte7xbv2rqZwYu78weDgYzk1ezJM0wMxhZ1T4KCK
MQQEhMjS5Mpf4BCLyQ7Ha5dSLu5iRp8Ne83HXU1dkEcZqhYsxAhh5FwBOW2RBs4Z
2Sg03xiWbivCgqw7bVtmj40ft+SqdWVK67Pl0uyzcsgLI8G+3sY/G0JGzlfql79+
QjNAyCcRDYtf3YuH2pRwfXHlIT5jbra16Bx3Sgi35LqWtsSzVeeMfavpexO/X3Wd
ELman09t+hl/l2oehRpvL2+DsSZ3Tsy9+fMwTfmle5uliB7PrYELv97s5K9bFLLm
zJbF2oLkEYKRdEzuwvY3wmyhG57NQ1lB91cXjTLEmdpJac0alqSoAkY03HSZBZG4
fDYdgzI9J9GbBoyREBCFScIO/BTVJzgIdcy6e0CipzzJ8J+jAv59gH7Ud/QOamHO
EHzAE0mgswVyDW9gjOmjWWObyJ9K6SXXTpbYAR6dHuL8rxBSWdXD9VptAJcWoOW9
kljdBTaSReNUthitovlksAckvXT8vH/mR/J0bVJYQ3+2nWq8AKC9rQoxa62bLFnJ
dxd3zgnsUla1ut5qJaiss0JqXZ7aPqNeHza1s96qxUBYwWfVGY/NuWWmiyzxHZ6b
YFolxys/idVr7DszbQ191KFhpmftkjk5BZ3BCaMnp6VG/8VHQxT0q1QiS9Ay5Grv
VMa4wTJdRmSiU3ksTP9MEYLORyj/vc/0/Wsxbql8uFiN60XA5CmscvkdF+xI3qq4
NWLGzrgr/T4fdKZ9dYhqk87wRlaSakk2glfKUasNnIGdO1jqh4WRQqcZBnPxEkhW
LOja8VfWIMDwvHcusIwIcgkJ62VvcIJMCu2CcwXGcmOS5ShBRifB/N62pzIX9keO
+x3T6X5bd3L2PhbQfRPJRAQbHQOn3XJWtrjcecAO1dxAVVgI9HQHpA3M0Evdv0qX
AbGZNS3KuBNgQ1Vj98Uxc/ia2k0roT8WidyWE9HzGL6+pguhxv1AvCFj+xL3wATe
nVj6KQ8vh580gtaHWAqey4BvJikCy9weP2adwxELV9rZf+4czWYyY5z6OErjIiDl
d6kwdreziQUlibxgF0F78YANUZ3qUImHD8H6uTSx1DV5kTGaJa3I1AIFR2r0EXQl
imrSeYY0HDKUUg2pd6E6CVXDLFUu0qF3cV0LsnfFju4xb/88hMNSe/TalncSx5sz
FmX7qM6asjHC59D/DYGIx1p69y1dL7JQ2P88thE/8E087R86Qt2mD9RkWZjKa4W9
XZRzK4q10Xo2A3v/oKbH5gTI7eCnhr9TxbtOAmYBihZqvnHPMlYiWJfm0bedNuer
9/+Uyxv61IbpwMzswEWSUqKf15xD2DP4YY1Z7j9X3iobSzNmULVH0norIv1/bui8
QtpJavnnzC5ljaUTZZMmY4adt/Cz2344AjzI2+dVPch9PAjsM/BnUVY7HllhfBg9
Rw0yxqoxCiKKhUQo+nSvQEgtvBZFWaJSJ+jgkz0vJyikINMTptWx1b8U0cJe2ynO
oy3b3bJnMQ8h/en5czkL+cBDgSSX4lHhRAPt6xaAPCRKV75viXLX785TVk14luYp
eVccp23fKLlwes7GlKvditf37hMEgj26nsPTolsR9VluPAYs3QxD3MhThxnBHWrz
1TiM+aLMgCIC2Qi9Xoil0LqgcEPeaKKhzibt/Dc/500qdqJI1zAa6eVV/I6zT43N
Uqf3lt+xwgXuUeoOUt9Jebad2cR48BskomOwFpiowAFgosbQmZEoLRybM8MyC/EI
j8NNrQFg8F5YfRszj6YcJ47fEqzqIvJhMp//OSEVnoEw+2cyqIAeP9mSLtYIGoo0
Gx/OhPLF8V36KTNuPSTwzxiBZwRjflRnQYEsLGOwYTIBJA4A2UnTcQvfqNvGTYtp
vOCNOqwJbCBSh0NApYqeGcyeEpnwFRIq0ZsLGLMIlLuDWIU+gtywRZ+gbnjBQ47L
EvE1v3B62VwSD7p72o7sxhzItSqCIkrxJsp8n8aQUL0s5clN/PbFQMAEdpUkb2/k
D9J70xZmWIq1DKxHFvSEccP9SfeSGl/ziDeiFlv0PN4gREzsFj1K3ZJCX04CUNOx
Ih+sKWuizbMOQX/w3YhWvGXbStAL8wCZaXsEGDafRajs8dBfDz4Kg2t1i/2izsrv
8hd1Gqt2IydV5+eG1xBKr894CdJt6IrmKKpQp5tckmTcMRwu7MKXSA/xh3gBVxE2
WdFxIHVPrbAIa61dxoC0AvYp9pTYE4W0fjAezoxlJUexTj6mY2xT76SaNMvTH2VH
XWP6U0UYbmIzTWZHdzGnxdUPaq7NddWi2GAQWu9IWHMUUzynCUDcdjhjWHhl+hhp
sdHRDOa8NiIrXNr7xieFzYu2Rz1m8ZKLPjRsgCezYrdty3BDgsawfpyaG+C18l8u
SBERKP99dMkUT+tK4jBFSm00gmtd4TWyfcdra431IJegq6NVLYN6i/9rcZZWH4ku
xrzS1DyOsyNkz8ZMnSJjkUzqIhBl6zAILaCl2nO7/jjfYdJNCB507cAjfeaGBjOg
FuXUs9sCJtNcn2Z62FJ+NH4p1LAMZSI5Gixq7kIUAdecviTzdIksXZUl9nOg7mFS
r6Ji7Hm3Wzk441MbYEEWPX71oVZZJAmXnEDh5Lxh+mMU+5fHX6KN3fE2ZpI2hA43
hQgZ2TwQrGl3kSXETRoMKZijZz6m1WYlymRGZS9y+YuXQG7N4bXsOZC8gJHIg6nb
mH7K1Zt+XlvnSlFnUjOm9L0Gdg3QecUwBipniKmreNlkYNuJlIyIPv54+BSCUVi+
24h8ewGzMuuWzRDfB87eGLhpgSgaDr6oWJqlKxlntd+rVD55RGZiWAoHWe54OG9p
K7mjQqsBvLV6nNKBUNy3GJA8luSfQ7pxTMsBTtyuiw1LewoXbAHQhl64LP9XdMtk
4on4OYiiKIiX2dbB7tAstUNVy1Wl6z23fQOeeHc58EYNtW5py0qbDSm8939M0lJ5
0QaXgBZJ4OR16bqMYagdg0GGPZNi39PghKjqEEbfOrp5j8v3KtmoVgS/OFbka25p
MlgsrZXWGl0ePDDZylAxh2gxQsDH2ZVkih7o5aNSodronF0wauVwQx6LpE2p9Vg5
8ldwpIWujREUqW7o/Mlfu18TRYvaPxr4qJ24nif/3yEqeRjYqxyFjUIPYKpMZ2CY
BUZdCQjWlB4YX+OoToUMSORgdIM5BOUBh2+qiFZheWxdABdYqE19e1d4RPa/kba+
K2GGEuZcyqpsy6tEzcZ46g0TIJyoH645prB8MYARhH9sB7lJlWfsaIyDRYnZtWkP
pkuZrEkL1HfVXy7InQI3+9QV46jFuyawCRkEiuJrVQEKy5KfykJwm5U39ZiVqoJQ
iyVtp74R11UkbO2ZCmJq3X9uNT7XGZQdCsTpUd5sEf9EyT6hebdjG2aCFWRY3kej
N7/Y1PoOE4K3EgbrmH5z/27pM9uq0m2gfNStsPkQJFAhzV79diYwsaECJxDU5ySG
J0zE9ZH+cEWlC8Nmwi/Qm1T4zKfhf2wgYIr6xpZp73SmRFxh8xuWWU37EGoS4LOG
uWQUi8yWub+Rr9u7YjAjMCYow1s3KeAbOHHSAzDRnLHEL/dBsKuh//yswSG+EY4k
DrdRO3PCBCNZ6d1rqmtSrOAqu6xqZPft1y51zJFTDFhZoWQuRR83BimjXMquZ3pa
nIcSXO4WOopIPjLzSpzgGKgRdPLXMNq0tXoHU4Q5VioYYFiUjoycqUriN/T6swHu
ngPi/X3vX33Cc5PTq41eMiJcxwN1NYQ5ZWTlxY9S9Qkq2N+vZRTlEK/9F2GmvF51
+Oqg9Zit9mW50BgM6EgUqY5lB7sRTn6t/JknmHlDfvEWwqChTFxeyLZgqJeJ7rV1
YUwVJqmxf+CQCiuZYYTfjb8Dnm1v3JUnl2slc3sS+cDwWWflCzBuE/mZnCUxay6H
MwNORoHw2/s3OjlyCYMaXFXqUneIpemSHIsx1Vaki7epxBhyZv+Ckwrgf44/Hu59
/iSKQejkY9lMiGfK5Qu1T8zCLRkix7PJ1q9XGH7W7fdwSvxjn8Gs114Wtxue/8+C
7qyIZ2G4PorRB2Na10GzifTWAPz/QdnMQpOgUGxCRVgiaxbHUmkekC3iPNeaWFzH
hLZkPPuVQUWIIUXnw1WOLGw4mEfM/RIDbkXgZaWE/xSfgvO8b/TEm5wdJnrragSJ
xLI8DdEeMac3SnQvADIQT2G8fIBV+yj2fXvv8UcXvp9Ynln/xQNgfjXmgDVC0j1F
tHO32e9o7d+ceHgQyrnXzcPmn1x8krJKKDHYvjmnhKSKVsvDS+FENY87op0pPRz6
MuyU0+PTt+sGD7hnU+0CCAlREbxTukcbmQOVtouwGmX7oiL5kHsKuVbM4Cy55vk/
4zHBx6VEyYyr2P4E6RjA1HNQPa/krXyxJ9F38wLx35A+mlRZ0wdx+DAw99kQrXn0
cmDeAAaUdxlWYR2MjHjrlA7QJc3q5LR125ZVgNXTIkO6/1uTbFKmQ+kF1dPO7DIE
4cMJxpqgEOPzZIqEyMNsFFGXdZCMNMNdRnoZ5uN4B+vGen5mvC+zbJgGg/sHW7cI
CYx5w1rV8muyYjQ1LdAZhGk8Fhd1sb7r+1kE2kEmFcPMBDQBZtYnRFHi+rhWiwoq
606zrvL+6AbIK5CyqaPfIDAVTND2tIyWJORFDVoM/F87fdTkSgx0tX88ZLQqRFRm
fPT5+Bv0pPJpPWU5mPlhLKet2ETm1EArPnrnpnDJ2nHJBleXu13DHlrQF7BifWqE
lgLssY5NSAzbhS3nn4EDWcTpZejliV0NeuoaTCxEJltUrN5LNEsb1/e+VbwYNEGI
HpVo7+DZJPYPBk9Mz7sejgVDjpBRflbbtmug+BNID3P2au9p/rKzayw0XB76p30B
JMb+/mhnF8Gj0tUPvuShDFe6pv3vgD3B/O90Ul4vwSPXciFf4ZyKpy3eeYnj4cQK
Pfvub0u+nZ1gHQmILIh83s1oTTqTrIYhC818aj+c0Pfqir8jhc2Ru6/UTtJEAkFF
Fd25cl1/1Gxv8ECimcWy8NK0su2SwY0O429bczuSldcJHHdA4wmlHRX2iA9TeJMO
gNrJu/CbuWc0Izs4kNTV1PCP3Z8mxouWn08jpi5G8TxKa+hBNOjitBfpH+R8aQLO
09JMTvKp6JBUcC1pRGlHuKf/O4fgwHqUz+FAlkM3dfVYFCq6jx2rCFwT0yUr/BQk
Qe6uAMHlQGX4VbJ85YDUj1xgFV9kCjn2HLXn4oRznqhbAGTECK/UdDMg5ZvH7G7v
Of+q3GNezO3X4XC3TM7W3WxLxMyeOe4sHg+FZN/phRFH6gdGOjgorWeNc/xCilVE
4r3S/a3DoHCroIOBM4VaQpMzsmsMVowGpzkZYQ79VuPlhzooGbiDjilqeUWFq8fR
nKkhZZdAG2vG1OFxVFeE6xQFQE2MDnHH0I7weB7Cmv5Ik0jQ37MXi/WBTQsryMq2
ZAFG+Pg4AHwlygL7cgxpYkSDOKHTIRg2JGU+zfvsPXgjaq5Gd0CrigT2SozYkcSt
VZ+xKq8PslKT1daeBfMVswkDmg+5LDlXQ2JUxagPkdQ+RlZulHJleQLDTFqvtFDB
h2YO8MfywTxTCOpus8YcjsFRyqtE7J2+TzONG+XMEtbu9to6xW43Gps8CBFaYTQv
cU6wkQWLLycQm2eNidWH2AB6lxCZSIJMD9laabiNfg6UpAg0HlzXuB19sQwa7laW
COfE0xTHGKYeFvVGjzHHRarTel2w3OyPgEtMCUqFs4NlZOJVDVVdlh/vjv/zuxi1
iinaS0IzoZkNDlzInWfLVS1QMn3x8cdvOYE1K+4HrekNv+fMlJCB1Uefpm4VUMWx
0dDwlCAyTVnf4QNKb04iRs1RZ8PzsyJ9hZ0wfQ4Z3Z8eBy0gWejCEx0QUZyFOuat
6INq/+u39YrSRmVyO/9X6Pt9RpmlGcUT3T3NLO0ubcWYOEy26XtPMe0XvfLKPZTe
BKdiNwBbKx/25q1CHxt7YFsXYUjr+mpdji9O5cDo11/KSU30oQiSJis9bYMBxvdV
fm81l15l2oyAMcXPZhW25QJSgLdQHA2UL40BPtsqL3azqihWKhnkvuaioih79amb
O7Oge00f+x2jH/OIR8D1i0ZsRwPcs3dxprcv31SKqN/4cVY/v1Aw+QKKDBMQx2QZ
4B48CPvcQnB0UJcdDSu0hQcqsEXAP3ewL2TVDH5z/dbXelGvNcA2dlX4VDk38azg
dVsvrd+vJt40ojxhai941eEekZo+MWzxsShMusRMJDi0GGhfcY3LzbR68lZyVrBz
QgZOth5PjraoXctOixPmQjr9ZtrfZoPQWRQy+f/EmMEhGyTIuWwG1rZuYDFy5bL7
TovbxrTWC1I62MZHWA11Yqc1lenrTGBejmhQhnPQN0RN8hr0OGyzyi47cJOKeOME
tcO+pXoYOM977l9cYVxkv3RIMv36/QkVqqMdyjurkfe6hnM29sixRsb2BARxd3y0
zeRE3ratBMH16bJfKS/K1avg57dQRJK0s5WPNw7Y5Vpm3A/fdggt4Lw4LZS4Naho
prpwufN7fj+G8S5aE06AqsPphHBDQGK34oVU31GgO/KGqsMPH9ES6FJWsjTgfYUY
nsx5uj/KC25TLMH2mDij0+nxbON8m21IluUqlS2ey+YUZccmOMdYfTV8ZDK0mdE+
nLiCSebCJr2xI+cFuhmnV7VG/fFPA3Vva2sfi/zSqaruEaTUIMLAPquRZzQb3h63
nv9/DeaSBmP1OXAnLn2+grct6pmaMHGa7ZgqbEjieO47t4onA8hqiAKcrvQ3UvCW
qgLKVbrm+H6mQazZFotYo6HMZ79HA4C3/fDp49ZwOT6G/wD0QCPOrjAOC77l+VL+
jO5fpFF2JwlwGFFQ7V5wvYZKfJ0FZojSdnCNSlJkWjOBCTPp8tfuuU2cjXZ6BgrO
6stebXpqkEf+iyGFzsm/V14EkHxUXTU7vzsjB+Tv3knOiW3BKfpfn4bOV1ONESSu
mw4YLBSLGdFhJMZQ8FaMu0VsyfLMTiv/HatYo+pgfXfpvpIuMw6quN1QBszvWZL5
tmAgGPoUlL+7RoQRQ6s9Tszgsm1XYpX1gbJa3MPVU3QJjrD5BmlRLoS/yX8Js+In
EG93G9Wxd4JoQWm6IpDSeYznu0r2Wr2xuv9w6AKad+UWSorF6pqoi3QidOIG8UPt
1o4OqH/QKVpKJ9zaXQXQuixHC752cwAU9x63BmUfMET2RQA1otMRbQDWyXJupiZk
AfK5LhHdHUxsnpMb2Tz+lM00+nav6Kcor1BasuAsSYxFJ6A7w8razy9pnBKAnir5
VGe42q3gDC+TewY4VnpgVKhm6Vp38CFdZaCZAbu9ura/AmcA9cOC/7JfLvUaOxkP
VnW9F2Hmm9NmzFjGzIYzy4A5WsmdF5rTqxhPbXYLtb+w6Nm6psZ8SV5b18oQZ0Nz
5Lg5rUw4wAcO3zGU1L6jgP8kAiH5p6SrY32AyeI5G7Sja2pxeGchLmICLQwd8seG
HE+Zilf1dXNEoYxGPou+yX8zRCsebMmbrh3FlBQEVSFMmPfmH8BxveO/mFEp2d2T
F3emNK8d6xfSedB+wxT7FNlpxj0jlLNXHgaYJmJanooB9PkpjTzqfLSc6uxWgGlD
6vUoEFkycIum9PKFjkmz/NsmkiVy+WZrJe0Cw4kyqpry3Zh9hcJJDnS/2krb8yBt
EP06a5nHFPArRPkjGR3ZudvoVg/4OKDVt4KM3ApTrh53/LOXJNtI6jIngzimhqiK
mLZZ/v6gHjxvpnbUsBjsPf+lOl2epKYl3U5r/lsHaHi6dgER1kmosIW7EEfSzE3s
nLLJ0nE1xv7Wx40J3s2I9u9kI5MW/c0uIofm8BQIB5E2q/2o1o97PNJXzYAlqrOX
zn68IATDtArmDm4SZcDF8LbtVoTOAyrH8HYEUaL9wMS+4KAse1+048rWi8DbaL1D
7mhGpcHQXmO6b5ODH9B5SvhlbNEmhqw6lHRJg1ts3u5DFVsVOCP40JguWzT4EjlI
AU2N+GxAS3doKwoJIDxTCRt0seIjek1Tl3nmA6Ub+UN3HhfrNcVum07FNTWnT4Oj
rNEOY7qVp/O9Z7+wNF3PC2Kogr405S7DJ0tFPxQZSY7XWs7PkTe1Mi8NhJB3FLRS
ue4yDIn+apdyqYn5hp1omH2okSyi8knNMW0eIeoXmatleb2bs5RokZtWcP5p7KBR
TJ+L57ndXBxY//W/Sbif5a2Lfl+hc5kKdyfG8zH7yGBQL5PTzVKtksEFcbicyii3
B+4PhApXT6CZ120PmRvubFIYbpKLCxZsutoJEd4WMstjmiPVjZsY1RH9v5e4J0rG
RXa9MUDsHO1/2rj5n3P26rECbebc/XMuGzp+s9hUIWAFMZbPioZbDvzu3BjGM9IT
8xc96qsN5S9kPrBeImGb8kpxFy9wbS5/RHZl/z2eROoAIDSMwLKVLSVVRiUeQ+to
ebuq7aciO2k40DL/07gqm7UW6q+/R7ZVmJ5La/34fPRQ+kkTLn6pTkCKFQSMkkjI
XMIVIRcSmpDYBhyRjV6MqVDrGrO9D4eQpFnRAz07rS10R5xsmPsy2qsyz9Kusmro
kg+GBC445K+YHUxZH9eF+CQNPtijc4wPWxZXSZLJa35/8ddwG0BSngAcI78WxyOg
TrBgVe4rXWnPiCxg59JnmhvT1DhzxIlmF5knR05zBY478Ckq83QbcSdRI0TtFN1a
yQ4zikcsMGH9kBMbOKXK1isJked+Al8m4sUoEsuJkA7i+9PbWx3m7IfKAxE+uX0r
lMCbMtPADf1MKJEaZvtuCCrZWtrcrb8XkPF11svhtpkWHu35QjxDwWTJfeq840xb
+eVhdU7hk3VT43QpwbLQfxxxLTNI9oFmR21acmj9CkEDMMXQwE7BI8tD+IA612fz
IITyBhVD1On4f1ulQS68NGt83dyBSTvdFYTWVVVwtOCmR6qgn3ZxYQev+Na246Ni
uYjLvy5ewZKPKfng4obGN3pGzCFxPqxAyrAHnBSfEDa9LFgJ1mPLnJOE0aCNQmhP
1d5iZhuotTcR77n3wNS+GUIwp+eMnr4u93FSAFvLp6ztMrNfkLjLIBW243o+jH1e
FmtddbUXu60XFJEJkB8zuyiNBNcKR/sIV6drVWNEG6A/FqS8056jZYWZoGFhkzjR
C6J91vDx/BltXLpiRQwaX4wO3fXJKQX9+qfzmS+IraZUT1r9JHWfvqsiouSGtGkw
o+n0hF3XSvon1xzE0q2yZHIvLX+lqTMoR1JX0oxPw2a1zQN1YJYXNHe4GryNqnYo
H3kl56/gxNxzGHz0pPhpYWA+q3w/56m/JM2XTGVELj/y+pbyyhD6qktPnqo4z6Ev
Ae6ZKSaQgnhQBdxUWWJhQyBSIy9l29vh9YFfCsEr9POCY1NHahiT1X/KGd+BbAa5
/zwbZsMVlRgmiIAip+7oOw7Ht/yu4qoWUl6DLce8tdYfEGopJhChmduGcS5+dhoq
+K++idAwQx0uxXsE6yH3qC+fyCL1ajX+fsdpS21dVP1EXguBRPkevsRA9x1+IZ1r
BpgJ+nS5vHk2DFY6zQc47VPsc4C3VNAQFaS6GklKu72keXkJhlfkS/NWoNRKQk2F
LI+wHuCjyL4sZlw9JHssupUk2knj5C+Ue6D6ZiyzcDtaiPO4hRNDvQb6G0+Y8PtO
/gRkLAqsGckUzTfOLePLcFmj1LScYo8vPv8QjoryS3ele7KG4x7lcf4sWDikgg5w
/ksumyVppwrM/OZA0cu+E/qCfLbvJTtznYiNAMzgQ6cDpOBONkvG6M0jZk8wSQn5
+MzOODwenaCY0yEeUnXOsAb0M8V+ANYHxvcSQBYRZBpG//FF9xOrVlezi72iBhRp
QmE6l1QwFDrtNUJ8zm4azXPs3hp5Zro8/fgFSr1faL+gDk6mlE88Gqee7vUEOjP9
8qkbVu2QXiPlti7cDUlCVwo4IFHOrKoNBNfbJeucbxCZDZGAWDYflSXrzqW3aj3+
i8K2GSavu6U1UySNtuuAHzzeERF+q6xZWOSqzIoSmRp8PCzgsI4Arkxtf3btX9dA
yPt7gMOJO8eeyZsnT0tIhp4AccxXr31PV960hwHL4QlikY2vt9plwmuH8qqhzUoZ
unsTOga6wawubdZ9KBgYUzrssvaAqG+4W60tLChjELgJ4JMWEA0OV1rFcggW4rP/
2arIPVSyfKSJ4GQ4Kzr3whAfTxo7gI1hHl9uWNREBtpqPZhYax4MS6F39NUcv4Ls
kR7B+oJLhIjLgt995MUg3HbVWehEPeL99t9OsMGwxM+LJmnQxnAPLdfNQWpECWPb
GV7quUvYjIebmbQ48+1poboS7Q6k27MrU+ffEVN/rf8n+O3rc7mBnTrBoVG1Yh0W
yhWwPLqR+dn6Z+rHB3fs3vI3aTd9i0yRdb5Y/EbOE5W4Wx4COEAxaQZ4BqltS787
9/g5bkkM2nWoOBbypOCshVmwa7OVIvle3ov5h3Bp01U80YA6S+BEUIvCVAOioLZK
XKBtkx9VW0vwxAHGxhg+AroGP3j2sXcyRebUKZ06aBBXeQw8yg+dW05/JkAmVukC
6tDHsmtdtILQ3W2WPnUdlI5Ph7c6ytLH9CBOb7w11fC+tj2idBXp55wCADYk0tgV
AAtQbvWxpzQjTt1Hr2QOmnIq3N2aOGLAk07PA3IMVssPyrYBxvumL8Pl1L/nIjkF
b/IT10B8ckKVX2vFYbOZfNCbWmDiwiKOzDoZj+tIeYdfxzFXWZ0HP+tUFGNANGl3
RxSZ8LrHC9JA1sCw81czTnK890tZeMD8Ryzo3OkdthH9czs6mrbCsQRXR3h9sgbI
8jg7ZKiF3Ufcd30pHtC8o9Q0PM/8daUXK80tVNhrAMAUNPKcCyCXexpfcPBq1QMz
2DQuEaAwixqPaketOcJ7ORo4UBqfXHi69/ZaNKaUhzrnGAAwwQqEZwqJbJZtZcif
91fF7mxwHTVlBwJa/iU2kWJ1omIwFhgf/S2S8Nzhk4NajfGVd9Xz/7UJwszk4frH
qpvLI5gNAnMo4/Ob/DSXOyGOXJBAr+o6Lo+nLvUTHUQvDzzyejk1yRsRzVKsoBJK
THgWp9yBrn2nK6eRThQ1oV9xCfuPZbfz2Z7v5liD2tKYun3kYeKN+QR6vPwphoBz
wkai6/AmA3xuqBIKnIry+Pd1MgP11t5JIjM67oXPD/aKUR5wRuRvq4Le3ukVvvPM
WGYXYf/F6E5236EUro/Ps4x8WXw9+22FbxVbDHQisP2xaZ7On1Khu9kwk8vsP2B7
sYOioX8tC83Mlh4PmPQ24MLeCvhrIDNwrSZroCY1vxGjGjJF2fMyNsP38LrQSjfn
Y+SBfVNd0qyxHeTxls5MI08gXppU+GPWpRLxE7fswQaHqYj5n6iaAo5t4l1Wbsrx
3LPb/SD7Es0bgBKVDJZQNL1ajBMfTQMEOlF/hC1US7Fsn0CYSU7mKSsQ0n1+KVoP
D8w7/1AIKfWNi8ZCRojUutLa3qAmNSw5n2J+hGzsUTVf4NP5Af7aT1hGvlGKfD/M
9V19OF++S7kwEXisxgkV2dWm8UfRvhhm14TSrxVozXvYR+YNhOFVxuDjWQHyZsGW
PiMMaaC+rzAINlWhXDpY/4EaThMonFEU1LFO+VQKGWjx5VOqPMN1Dr1YWwEony1O
s+u8iHu6w869NtbN+a/yoI7xCOpU+E2mxAcoEDtdD+KIA8Klg1cfzjX5rM1rrTA8
0TcG7z2ftZj2mTU2bOanJgMT8xqcwWrrfmj9JUYiaWXr6S8h+/USBtF0pZWxy7WB
+dgxf+IVDgvCzQH8gKchCbbGACLrgDQsuGjjexBkpvETlcfCLIAXAsVt+F5eAiup
Lb9zbn2Vf5Q9rKFp0Y3M6Z1XZZPPq1PiOwG8OhZfxMm/3Go4xxE3DDT4goAC2c+7
qDXpXaXlyO3DM5VvCpxYD3+KuXh/qqU+Cf4rlBOSr58Dw+5jX5bMSvfb6qNdg0Yx
pI+rBPz3/MK46c7R/jaXpBBmDjW83mHQkbRFrwKUzm+d8tlgn1S0bvabTDlXmqs7
EcFhPiggt87HTrmogzDDIaqowYWivsFSLKPYl52tvNFNxkw4rHnYrKhJ+IwmBu3o
a6ynHteQqmhIqykqR3rlNun/DHmkaI0EZYKjLztYJaF9H5jjPo3eIIZ7cT4QbV82
CWu1p1Yr/Y0AIl6UcQ7cGvd7NqMLyEkBZ/oXXf6k/Q5CfrDbj4/A7CaqWvE7cRAJ
UGZYaVBA3PBWBMNFSE2m0k0K6l/4SLfGE/9aJfrvU8syulg4CdE49G1PgHBNmsnv
HyaI5di7UCl5dfNAtLnOFPOXEOJqpoLWkIw87D49oyZWijBxZQC2CTkGeDbtj46A
2Sk2IomHaRzHqlwoUNBDI4iZSrKky/1QnaE5WPxcRVN5V7Zawq81xSU24VnqOyYM
WkbH1VrqcIUcEtRftXWSncKMqOftKO0eMYX03dvpi6EZXb+YExO1qU11xocZ1QjD
tx3HesB6rKe3lN74pkW2FgHnqYQR1QV1MCINb6E9MhFqLUPwEbzPOufQP+n20G/r
sZ6fM7Pr3xJ/YmOtKtVPGtNxwPhY+yc9T0xVDIfEvu0tLnKVH1QJZY83FFFH4wNR
/cA0lH0Opt5hHA+ZJ3kPvKPgfZ/bITUHb9P/4+TtSdirWJAp203g2covnFBS0I5E
pY3arHU1aIaWGXTRa/pwNgEiXBd2wOpQyw2s2IcucNLQZfCbZARhgFeLcUDBACbn
ZvQKFayO3DEP/odX3GVWJbes/rtAftelMfQkZmapwDlG6VmMZee5PQULhrlt7lHB
cH7UVpILcuSwaSTP+JiLrbksl4/yrki35YszqR+rg+Q3pSKxL8w7TwWqs+a16YdT
u0smoBAAfpzgidMD32ixVvbvCnY7WhZaKx9Fm9fOXAd7Cz46KKKgAZZovsCSUB5i
2pabNaP5yjb/d0515YVjiEKgFGQaLu8VQ+IIalfU6p5hJFQ9ewnMQBoc9iNOAc7I
1KHJK3semMeLqGHs/R92B6nAwAQkZIC/nCAIcaw5NADnPl1ydGJ/3rSrMX91vMWK
IyqoKoXJj3rXmlDYMcS/h5SwlGptUkox7epWQKn6yQpSoWNBdgOa0AE3lx/vQZCu
LgTg5Kbpg0JM1SAhIxDtbKr30ve6RsXNJCkl+70gOoDJxSegwzaYA3puT2AbwtKm
zoz/T9uca2RIKlRlTeo9oNJiJnJQop91x6on77J6jJ+yp/ZWDNbJniDSpKPjvKK8
5tpJU1pws9WRgugFgLo4JpibmwLkzGQQ08FP308l3d7c52OdKTTBIP9JTydECU5X
f56y2BNUKAcAlWYSkb/tv7fO8hdBp5v19mjBx3th7v9wAw8yENof+G/nVu2IgIw1
LJEwQAfyrjVB540lG9HbiAhfxXXsTbIwraRvHLxhtshp6Aq4SAwiHPIstm+1QtUm
ocmK/fbcZ/DvJzFmjo8+x+CMVzoWI9OkuStEITldGnZmg1peE2nClCnsttiSGfDj
KnYhX3jfp8tY+eXc6iBC+4OafptXTnEXrQ6AJUDYQcL2NIIoXKuje7N32JTpbqEx
7Af4iHHhrgmfHI8PAtsmgMyXdp8GCkQNoaRB+RQbcsSZCenGA6uDfDKVrK05qhu/
VUNoZjBxg+MEBbD6Nsw0tLk1PXXEWIpsR922UpBwFRwElfUNF/Olt2BbrsYm0TGE
3Xk1FxcToCKeaSMxNehW+ZL1MdpieZtBIfwWZNchph3SLcmWl8wMjBXvg5XNC09Q
nCfSE2tanwOazGuzwDdx0Hp5Uvc3dfnBth1imXDhRucYo3esPpn16kJBVm6PW1kv
KA18obanfXI14Qt2qedOxqQv/1HR+WZgquwnw51vQVOImhmS4Q0LNDt3Gcn4r5rA
wmNit6AYTca6Zs8fXDXoiD1fJWIknOXhEsXUKq2uMxpf3nxuGQr1oRbT+TYJ16nH
tZYURdcJmRckLPZrtpz2DPccOtcSFayOaCABXoDpmRc63NGV5h+Hm2LdpQY6pDXa
xO9D/TxlxCNgfCPznivXV+WtsgyUgxLt05W5pXomqFm9j7yA2J4dNJM+6dmr/I7j
MN6LNqKvX3a6rIqkgNV0szyPoOgfNbX3Dhi5DRadcqqgbIS2mqIas6I7031mA2kF
NQAqjNAGx+biG9J98rJOu5z8H9XfSPN7/YAD8A4os3ickXJsMlrnHjS8Zm0A50eF
acEXcdEa6ZhSPKrKCmB3NFYC28G3Y3EWDqnKKGzYtNKDfkZqClaJgnKQ03uJ32GL
V5XQQ0YB5j++OjM0IuunAvlEJulvYZ1SRBpprMwlKUTCe+b+tEd6qVR0QuJ1rvPW
A2TFW/urneSWii77sgn24oxhfwmq1qfr0KyPEBzCQB+0gCfJ0R9Lcf0H2UystJWn
+BmyvgrLnZyAnnoWPJE1mxaUmD6QYqDtWEE6X6T1C9nOpdEdzOzLawGDzY4UUu0A
FhwJzvW43dU0ul+Y2uYOYQ44gMc41Z6HQ9ZSoGqybQizFXUDlUi+8mw6lFyrHNPz
VnL6eVpNDwtDMRZ+nksxQVB6Bw9OqrUJQ0xgeOWtgKxSLk0jC7ZSNGbwudlSlo+N
HuqKfahwC+CctpbqV6gv76C81/j11N1t4BjccuclmCFDlrOnlaxYDnzm8xG27G3w
UBOp5fM/iZzT8QaFR2CjIGOQ8P2KM7cNKu5yQzQASDzhtSeVqTgslRTrfb0B8YNq
PDsfjdiwJh68uDTk6MjUtqw9V4Wo7JJ7q6/lMzWn3dDpMm/aUvhDE3dcaL3ci1eA
9GKkLUj/2nncJODp+AcJoR/RwR/tk8WGSrxAVl0aW69IV/2snid3VIsY5vaN4VGN
VFmgN4t1yUcTwcELal5YA1md8wr89cpjJvedBYQzZz2TriJZSgSEkIimWr+DzezM
1+SkXHMDq/s9xBCEGgtpaXwJHwrg2imgZn0efA7r+R00DR/soLhukJybvmNc0OcY
6HqMMzZHXhFuI/8+bbDBdQS4MOEUHGc7A3CZwNf3n8+bbQtdVB1MPE3xb6elaUP5
jGMlS3R9nn2Yc7QGkGFiTxe0kAWtHJ4fUfsG3Y/A9qN03n2yftmkUtCJ/OzBsqXf
r1275d6C9XguDUVXYznG4eBu19izjcbchuGFtLhKfbIAks9xWdR8KbwRYwjN3va/
VlrF3Xq/IIGuehDlRmBQMuTtzRjKgXZZv4CyqxvSpKuMKAJelAiyfvTy2I9dspK0
i8RQbC7BNJkYk3bUNku1krSC57PBDiNWKq5/hqNdPkmt1fRjCNZwDV6rZY/imzYU
BJCBwI6fq7wZOq64yWCpofEY18eQY0gghu18pkJU2SO78MpOmCzNqKJSaZeUBipW
4pHxEZGGsFwCjfrIOtgfpNDrj9YyctQ0dwnUekAbPHvnqkCwLf7Cm8YPU7uFPfAk
64bSpv7mX3VpVwwOrTSTHq9sk2W9xjG++Ybl85XCi+vFxXczgWb7yQmSaxoWNZm0
J869ATJoSZvbR16L7UvsWAVPGRLCfZ2On9bpeB0DevlCO8aXHc3k2+AvZ6rPUi+i
YsSJ9Kd/HcbfIcy4R45+yrg74ofdg8KFzCR6omFcGT3ATO4BvDJsJ/RvqpzoR7jj
4BQMiua7IAgzc9TQZMdzR2Px3/I7A8De9lUX62EUnt6viNe1KDVil272IeJkLhG4
LO/UoMTk2geB7j65o+xjacw41GQOVZc/fRrdvh6wiXrsV0yYBzN7sxX1xg7JFATt
jvEIZSjw6g/t9FaYhBKsv1woM5Tvs0r7cC6Qr/ZemgtS6lfyf+mAlF/pe6QrhIgR
s8cmJJjRd2RXSNnkq7+Q2ODyYjFoxPKNAyxIkeRWOFSTn16Mio13M58A7NTW/PNS
o52xFt5+sqh2Mm8qPb+gAwl4BRwYY1M7Jkt/dd29NQ1jRZvR/4JLniar9Qgz1aOX
6qgcuJDSq36Pvm70rX/ugCcjrBUU+S7XQT4jYckB4mfDZeD65S0SlCCWKHhF4bPA
V1cptdeT/XTf2Ov7UbCbKA55G/38wmrzBGDR9PvDp1VNSaKbMG9ZHKtAvTWVcItb
Jc3KT3CtcrGXO8Yj7BkJX39b+zQOK4L52S8LD1I+oIahNaCr6k0R/TerUlR9Pa/H
v0dG2g0DM6xvceYFOkpHCYJV8/PQyAnxd3JK2Ps696dJ0t+CPAp7uzHzFsRHOKEh
PEQ1rfYqsfIDn8Aupcy+DragVNoysGS7iXqxs7kxwvhqAO2WZdw5fWH2evte4NJS
H3Mf3FPv50KL/g3tNp1YX8BEjBrCYQcEg96OJ2jXKbp0efB9mkIoRrQlnwgkj2+H
Lp7fF7zs3kZgOYsaXfx/yhMej88kMbqCswsQWvv/mtQ14GiYjtKLvkltXd0DF7TY
X/qvfa3SrIctEVS5N4NTDLYOAvdYDK6gsBKZcLKwSuFY3NB1/a5xSCvCdA7ye5VA
D8DQHLDWIC2Uztf0ZS8rXwBopI3nko8DqjgO0a5CxWgUkWqUIuwE8jbr+CQqCC3K
LIrrUMc5p97rfEjJX9Qsvz9+vwz1SAS7K0vkXOJatXfUq+eY8477KCz0CISf2V1l
PW6WOMvPo4i8qIypvgujy544DI84WKEM/5+8iWSIPy4GujL7jf+WFuMZmVe0tZPG
iQjU+H0S6xp9uRqAHsHUnO+rJV/sPXRXhTwFYvhSLV3Xa+C/KoEo43eBvX+a314c
OrW8PJSf0WVWiJJYv2DX72TLmbghCrTxV2z8W0R2gcEox9R6n9KYj2jAczshvZCn
Gcx4wH3jltNhdjEBY9Ecc7pio8Gt8pUHAFGnAGTzlTxu/UYLuvznmqUCY5J+gNsJ
5mVZDVrtMQYkdBoerr/Y7hZ01dJQYzYdepEW29UFDdETUgVDJMKdMg8TKSZRivak
q1ym/KifdBtgMajPbRU02h6xrF7X9FoNaaMfdwRQhWyUoVOT88pdqKQwmr9i+j4H
DQy6jKjroiUvwBde1+8RGs94iPt8zpls2ysMK41XmHS7JGhs34RZjbWUIoeTHXhC
b8MiFba3YYzvAfPpgWsot3IdvlzbW2jA9UiAiSx7Ztv4trP5oHewdnbD1S+tUfFd
jEM4gZQwmdXl0BQIVl+gqS+hGqd3sZ65uDex74Glw8UkEybwIJPF3hR3czzlVFpG
4Iluhs/M/mRS+MYn9wVPeu27vTudjCBOOPB4FnshTlP61NPu6mtoPW3KLfjpzaXE
P95QEwGjtMK60u8d2EbmWegdPPye5Drhz8ZJj4say/fV88ClNlEA6LVBTHUr85SK
kFiLN0/9JkgDBJ30PjbgI38nmMt+3bdjBApNsdvGxnnqk/cN9tsv97moa7SWQtT4
v++Kf/i5+TjGgFCJemuj4KAvRkxt8moO6HkYyuXR+2hXVYFHqbyLuMFl3mJU42AT
DQ6kGJ7yjHUP1IsMNlSMh4JWTvNM/nmvTXfT3zX4PzgdtNcDi9pNcF61zZ1/t6ZS
LRDh0pmSBk4rABmhQClK12GqxWU73U8CdQobq8FA17SCcgZjPEAZtFZDqHm6oPAh
sVHbS0sz+NuWcTz6WuJltcGi5qnTaXTG/g+LrGdAVZ5QDrzg9XCNrEGceOanHAiF
lUjfHVW89jo5viOvRmVFwd4YpMSL0YTBx+Yh1sm6k9wFmtXwXXlqcAJ8lkbzG1Q7
dd7CcZ+maCYabVI/1l6p8IEm3hOKdVT8gdtqhWGy0osyfn4xdTDjAFxb05ZXKHIU
K8obzCIaj0Od2USGAF/AgwR4IgZZiWvQDXz27STfCim+sUYhMnc61iYbEjPmbPEG
o8zAJEhag+Bep8kGbkcvYRdEUjGtglFjz44ZK68FxpshjEhfgVXncnzrPgVjJoub
b5YvmNJgQQoossUD7xTNIPFk1QzKwZC1yMyKV/SMz9Tp2jcM/O3smRURroLxMbDf
ezbSsaqC+1DYM7RKIzlPwcst+BF+ILeAUC8SxGSdQjXivr7vyFAHdYQZ+uv18g8q
47ZS4oYKT7bjYTaCxFHNkfyiuHO0BY8QSJnGVpQeoJqMSDFQx0P4cuJsF6TCNci9
4J8M6/scyvUGw3kVltWPI9Y1CbbZCXHkTcBkMXDIaskYsYhtb6bWKJDBjlwxFP89
WoxYFrwfm9YLtM5VHnxmd5ZQIFcj5aUuXTabrAfE6OD8Fpde98VFue6hHO/DxfAD
3LzYF/uQoDvuKNy76WSKpBhI+sSXCW809yIkLIOTKbqCLEWki3VhfRV8Kl35C84E
554/9bvgfIwK52551p2leJF/T51P3bh8SXXTSVi/AZZTrI6VDOUq0/yNf0KemQVn
OjcrCphM86KWpmGzdleQsEVXDUKnZ1wio4W80emTv7Y71l9tc6lAOhP9emwM6peI
kN8IOaoatAYi8JGRqa1etJiT63NxQu6fYXpT/eIMPcypbjDLJYqrDGHXvI3xMKsN
LMR/lEMBao4QUPlX6KRZ+uDmxMyFkVJmBpTbI9a56/SQOgWIwQGnFCBQ3/zuukD5
nZSuCSF5KarcGRVyQsuXpkX8ah1BW7l1q8LBLSGLW3twqZhzxW/t1NGfbXBoriJv
/+Rtlv4nzirx5xEZFTaNIAkoftX7lNYdaaWvAPNXlTLl8f8GM0wCaui3c5tFoUS8
sfQLTOkyF11rwg9OT/Hw8LnFin2vWF1glwN24AcYsSomMUu9Q2HLkPojpw4kY0Oe
nKVPDAewHZPl9TWjLVSqwzo9JmyX0TLS6eFYauu1bacgv4tS59pk0SRQFg2RxFzj
nJgOZ948lgd5K9AkAF67ZE5g2pAJ6nAQVVcs06Gv2B5JdOMWKc7j0TehG+SBP3br
NU3q157lPYWALrwKGso7GX4AKxSsCXCSQSdo7+X54NSZZx0cEHDex4YMayjEAj5V
ULIzGKZQ+rvyjhSdNkgupP+yXqDsHewNqyf0eaRGO01etpYFWfEyKLTjlY+2KiSw
/DluSrIrSnAqEVPUbuLqkE4Pyn0IILZoV4Z238tia11qXAbRz7yrAZWirtjUBbnS
FZOEssVgzzfTG08u+7BaenFbMf1bjcxPX/z8bqSuY53OzSgnQ+u688/eGKOhuKO0
cGRzoHDN0Jv//IuuwabGu2Ps6DCe2BAl/gs2ZXHLdTig7P7ToiHZnjueJQtWlKbq
WEE/MepE2q/BwHdC66NvI43mKRAuX1UfvXMx0dcOlwXcXxDwA70kQ8ZXt6pUirWY
ULHFEWAj9cGlkUCcCEvL0XmVyTmApCCaZEv71NcpMrtGxu3sTXwEsstL0kODuz8R
w6taurEPA+xHbPBK1WNuR5v8en97INl4HTLYd8WpAFCYOk4/FLG+mRHntZrjijF2
UpZpUPMsKl736pdbQ8DKxAUdmTvVaSOhpnP//m3uVMVRM0uoEIM4pQVpivkmpNsp
tDU8xL5ol0UcLAhSY5VAUoflNTHIYffw7/tC5sh0m9dR3/XYYuPnNVNuj3+Mk/We
+NQJAhjuQqE+sxN+oFy6woid/Z8rIFF4tdxCQvfGkqRLsvBMP1yKya73d0TQmWyH
lBCxrguaKbdjCH43S1A/94vq3ozIFGNAXNl6Apr+1mj691ngnfuVkic/uRgE/KoX
RIOqMJCUMzx1AUAmRqmj/jbL6ZnTEwg9i7BdoV/nA9vP+eFDcWO3eKuf0Pggww9c
EqNgFrvSU7zITIMVaG9o7kIUx1M87I6Oj1itTZ2Jc6rb13D2VP6ZKSHQxLNWkRb7
S1gnZ1IZlKDYjnGW1g2EvbUBB67/1pVb3dT0xMmD6bgieaJXLYWka0/1wcRCTThv
1O5ZD9TgHUbJBXtwnwWi6ki/fnNFibJAwtIc9yKp3Gcb2k9m3VDrazuV//haFx4Q
t69iFV6lbbmJvvHCB/GKCQQODS5s9YTJkVxsbXq92cXfpQLAYdVyRfxKNco01Xa1
f7Hiz5t1MiXjvFdjeZuvbuny3Mh5pCq/0K+GFFNc4Hh/HpOPDsVY74LaNsHITD/H
hb21n54Qx0hXCqbwiIGmT3I7lXVAEEM6TQrZVsW54Iz6XAhOECkdzOUIFoUHaAYf
idGNAsE9GvwmVwSXjsVokA9d47v7N0KRjtAKTJyqyZKh4nSbbjpjXF+QHeXe1K4N
3fRa4+uOdTqzXFz6RfJnbzH4ywWLxtkK0hOaJuu1eh9IokyU7Mo8O6+EU9wj5XjF
RR2hKFooZnyd4DOsA0ZLCicUdUVU1cVixIfYgomTA2QtrXjvEouBjUQJC0ekVHy1
g/1a57MTrVtSQZckAvsbZvW8aQHPYSWulQh/cwt+h7RrYPZRJ4X2zheFHCAi/uFK
RM7Hz5I7H2V7O+QNoy9xg5o3HtpAr6HeGusTAIfFMBuLmcR53ovWFZYDYiksvAMm
P/tF8S2cDwfK5/10pIcYrItw2iJsMst9Of29c/7u+cTixuacxp38PjdDZwFelFXM
sYD97dh57dKm5L5bXcVzVS+ClaMBud1d2EZo6WKfzzdhp56Lzkz+AkfiFEmgIXEz
ACAtliq/ntjhuGmaR5NvOVDVMLJX5UM9wJJrRVqRmXgBhoq+JY797xpdX3Nl8qdW
kHhQiln0q19ZH65qSGX4vx0F6Eg8UpdPuj3A1m9hlsDDgbD8IX4H/6RewmR2rGo8
Rp8Wb2cvRAqHdnunOlGfYGRzdfngaCzb7/iBXNADmqiF8yft/20JJg3z/qEM/B4j
1A82NBiJTOUqLZM6Je48kStYnRHkSeQMt0xUzA2zXKuQLf5GCLhfQ24CJBpfuw2V
AvHIl3sCJcJKo4DPhf52Iy9BqCSY29qeezRGT5pO0jbZ2HYrpDx0hw8EQHjkLTH7
lxgJVK9HdovMgrO3YRqmUtzq3mRHNDDdMpU8CIPKyYoJJG9vlp8in8unVimo3uEd
uPiBz93N60Gc51iiT9LmpmHdlr0RgGbd6DBB6T/EfB9/UKDOJOYu0PrjBYG56ryr
aCYb9XJy0ZmrwJfwXhEWZolMtkLpXMGod8o3AellqrDTuBXQPXZbxPFcu+neDHp3
6dpy58guoB2kkylRUcNY8i78UTdoF6WP/KenEsnQdthuLfO/e4x8hpOz1tAcLql1
X2q+UNsHxl5rKHuKlD0+CQw/MiDyFZW6zTY0VdSev1KFe2SP99RTU/1ptrgnrB4Z
zKx2Na2rkoSS13N9maTpkemazdabgr1VW3yzM6q0e6/1SSHMbWCKU3vslmFT1OLL
ZjX2g2x84xd756oVjbdBTZb839uhfVmjMr/MhSPXozj5TUylsj8skm2LrfBaAPoM
TQs/S+XQzTkCKRfzFfHbteLC8VJ5xJ68AgYZvy+PbwtYH4Mav0/W7swe51YsvP9Y
49KQ3O4GFN67ryi6L9j7KZDrIh0jP6F4OHoROQCmWAQUP9q//X6HziuQx+PmaoTk
hKkd59/m+UOboVmlWhWP2yAqgl/MKjdWqJOA+IGVObZblukG0TLJ0LXUPKrReXKj
Lxg5XgycWnsSAIda5DX6QMKAWWKZ8u7QzHCZDVqTBNMYwcYKA4viwGB/ki8VhWN8
eMBJP3sLPJbgkM/UcZfqldFFUA4Ty+pIuK50Wy0f+NiQG8zuzQ11h/Somm9Jw2nt
USSc3o+SWjauXsTluCZ7OEHV4xOD7q3eATGlpxIPj2K2sfi/5CsiNSoeHB5OQAal
fgEHGe6rjMENvhkKFTOBrOa1cCtMKTPhD7zgMmA76H0YQUj5cELZK26H3u4XPxoL
YXafoP3UIpljQL5M80mo4fWjsEFSZs495Z0GrO3sEKzEaN7LlE3bblxAgisZ2JzN
Q2IsUqd/OQi+YBg+qyCt73DtN6vjXioKL2jgvvdKJP2mlkijMWvbmvq3UtCCJDR3
ypuQT0zgRH6D/h2LCjvhdaCsKQu62WFnJ0X0KhTy3W5fBZpxz/1GJRonrwcHCUPv
WXBv29nNQmeri3Dq64XX8XI4pdUBLD/PRajXa5/oINgG2vEtpGhkvgPgxX/8YaWY
fFdlWi939YXn7mcP5H8n+63uYct6Ir99z5gBfYyUbFI7uKemm8hV3QiVkM89sIDs
Pj5qNk1bG3r4Re5dyQf7hGAbKakcbD/wSyP+wVx2gr9DYGQoprAeI5MAlkr7TtsE
usrVFtCOtIEFqFZrpAJCgIc/rMETrW+CrnTlsDYcqGooUVFnmv7FsbzqP0T6X7L5
Ai8QLi0H+8PEP/qvndCJ1iuTxcEyMAyDMbFUpr8e5+o0mI6yVO4lWq2Rg8P+C25x
TR94fVJ3aVlG7VhzUkMkmDHjDlztYD/YyaXZiVRV//l7+3RWJZp02tKOOgLpUV1g
gmMZjDXVQWZh5P4ECGoleJpEam1ZO32TnY4/Ex7gj5rmZ5z/psThrpt/+7krxuqb
A5z4f5T00GMl1f21YXxUNl01zNYwntlxPBKwp9s0E9HRdb4RXYAXPc2fwy/DJma1
CVSgKtZbHHz/cA7I6r+6qjPp4parq+7yDI5g/jhYGpKqPBx+5Ji0s4AO0xbxYVvo
m2VD1P6bagF/GlMoRjEYDlBxBbMvDzq/yHIlalzhUCUxtyjGXuYdt0HHOcJyik5J
I93AfbVpYI9DROwku09rGUeyfv/VNj39txSb4V2zgPXOAbAgV26Rb4QJLNOweNcO
/ymZOvzJcOkAx5GGiTWOflMsnqnSZ0297WMib1m6vTtcc8zjxTV369uO3xDy3jEd
oECt2/xEsPMSKxPtsCo4jalLaPq2yLA0hxe35roeNVZ3gliiWDEPVH4YTxWCNJHM
m+A5+meNGAJamQPAIG0azfLyVW/WHm8e52R4RVk+sM6DqB45t/3rqWQ80MEbZvTq
L+9a7zL0ysEvv2tqh/kqibzVmYOnzfbLcr0uuYvxK1Me7QncLEGq1WcirBmWd6oI
QiuBYgKk8VmxqMlbxf/LuRBRP39Y3hf7gztkrUUhmdn6yDMLxpC2VZKkFMotkZTd
4gX4m6hbbbUGl4BOzYAy7s/4BZt4kxgQJlUdNb/yn9By3clDUJj97AeSQvT0+tpo
GOvNFyOYmNYzgVjZxFRlgtEH+R/O6gw1Guh/5JaB5jn26ggzjrGLxs8Mf6r0aTsj
BN5OScal6M4BYnumfe4SDR2HYeuNlbpdh93R+4JpRDi+fiTHMf4QSkAL8FRhWuOn
CiZqZkisKJqM/p7xu84jbxTVMkpdPn5BPXWZ4ntn0GsL8sv/LVffIpEL3lItEl3J
HvlhSikg6jdJ57jDZ3o/WGAQwSYwuvm2LfI/jQgT59Coqn96LxY4uUsffR9utA1n
+mFl6k8x/scTELImQTV1Eb1CT/mui5hGaCPfbiwJBejVccMfQJtjHBuIus6lmwkG
DHo0JnBIjV68u2YpY/+hSzsPBM0GKK+bIVxaEfAdz8xpZJSDDGz4je/2+tnp4+a1
5xYyvnDFZLV+bTzzNxi85pZuUUmdQi+DBV6NrQnufjUtASAUKTZ47+3BqMecxxZy
YNccweRPa5j3ZNbvCbG5bOY57WEZmOYBIaMC2c/pEcAU1RT55GEcrYzMccXRyb4/
GnNitc5rW8Z2vJViGDgr9IQTVqA9Riw+BI3tn+7zkleR8ZBge7mKrNxf/iaxJ8K6
qEbS2x2lpnucGsjIA3P8KkTqT5xvqrQ0+jTsaMEC/M8BCkVyk1gNCH9YFH1TSulR
NYmObh71s0bB2kj9fbnIlABU4IJmvomJ/6MYv8wcumXlGwBwEYuAljVu2btBBkXX
0xq1ZxshaDHoLg4kkaaiPPuJkaIhbTuBFC+IxyoKrJ9ezZP1U+tTr0uR8axMuzmQ
uEhUZZXUHzDwDDff3RuXgXWmfDHvzlEAYcIoIddHue37FgqFsTnRJXgrjf85Np+n
hzB7N/7x5R3bmIg9mICNn2nIdRbHYD/K7TgIzwJ1btCUKnIw3BvTt3t89TrOpxFy
XS8gyF4gAnZz56l/r1/5VMWFnQdq8AUKNoApUUbuZSE8+y5/Nuy+rxFd1e3dimNB
z5MqdbLey29SpOsVVONN2//3vdMM1dNDKZR8GA4zex44BtU6Wq5ac1IyIrbORe04
rjCcrjBRhRli39BUWsEIF7CnWi2HvVaEV+TE4qO4tpK4FNmxoxjq2YyR/SU6nEP6
POFxYnaIcgmoZCbs/JENZBqmwk0igJESvEJgrzhBkwgln+zei6H4kEsxU1Xu0jHv
GaLtKW/WcQKet6zqNrWpvQbBGuskSLKyzbsBngvcVHyM2UCaM3WW0UEqxu4UxJfZ
whLPHEtqVta/QB8HMwjJso+moFgrmygFx2KIJRWGiFRgOzCLEItDd3xrRjfOI4hM
+vvvrpa43SWqMNkrKb1p/y4it+bcTLou27iv/HaAkBFGtcLmPVrMtMUvaOZHPrCO
7oAEhx+2kjUG4PmJfVpP311D3glBtjoK8PMIkv6tbKZ/PJVjQIdeM1riaJhmUAnW
LxDq7vm915yC0cWdaiRRFAwwhnYw3rIk276CrqPpFIYCpb1Ge/gRi2cfGjFUNERQ
obYQgaR/BE5vxSuodu8DQdAFiZjqMA6uZ+a7/6N7sHFlDBfGpp+4XgOrkFAsys/S
s3iKjfF/hyoOnaAfhn84+pF3lF9SpnXPhw7d/7wytFxDN2k+UPm7tgYNegMOVlKG
K9S9+9u3btfd1CfvXlrdeEd2WKDn6ZV4o6Gu3zLFhoBhqK69w4RHt1lXRU/D3ZyX
ya9k41/9u3g4GpAAqcfuhVex7U9/K9d1O7UYs7ZyUv/9Olvl8wMYHwaI7Mge94vI
nvMTZrdgFkl9rP2pgEV/6MwwvF5rFJzOggRPsqy0sdlbSrWO8bpMWcuEeEKvq/1J
23+FGs8Jad0KvQ+RwB7zzRwQAdPZTGHIU7J8lZF51Hjj14CUQhkPDfbD2kNxMY7P
ZqcJn32iPR75DOI++4IXftzF2CjtDkkGdNFi6ZoX23E1HwETh+kzKye6Z3isXX33
Vp9uxdFXef+nF/KgYwgphe9rkhUq67JiUbV4lrl58LcvmaqkSqFpdT6XJWQpCe2I
YzVfPP4wfpD9fR1dXJFZKCvCZdjjfYNd5RSRB9/s6Ue7MCJaTbBFsGYBGrTOzir2
80Tq2gcYchLjp8hVlwdyYmQ7+FFf4f0I2jkAa33julWKGyOz+jjwdlYopoEDZXdT
p7VN5oBCe3OYMR6gbTb/Hbl52HiHNjrneHh2X0U3tlm3YeW26mW/wY0QKuNqrBGl
ARuwCaeExM+fGN5+nV32s1ba63jnCwnPTPuA3hZZ+hhDfAmQ7itAmUqJzx16567X
dBvD7E43XP74CQzME5mmLe+mhMGh/WhPHRFRlPHeZwXMsHowZtKTP27gYI5GXwaF
7zjot1is/CwDY8e4XXddeH5R3uvVzOti/WcVWc/P5fUroN4Z241IcQWpJfvvCpk1
cQAV5tadeHfM2AW5ifEExbtCVh+ilmdIEFky1vhwuGqoVYtgdppKm/EuHZNNuaXp
a/f7dRGKAHF16imMKYYhyUvqrVJTXZWlcMmAX2/IJRltOZ4lp8V0pNeF+Q3bmd7A
deQ1KFujtuJ7sG7ysFfllTB304F+bEDYCldB4qAvHvI0/fA6y2IX+bL/hv1w+luP
5sEftmS+gVvUKnYCEFdXS6H4AcLyEcYGtGdE+LSmd5Yz3Aj5a0swzw+5kKwGLFy6
lpijeG6tdi1hiubDScqYsI0gAltZ1Nxe9hOs7A46c9JZNiMP8VpfXbSAYcZMTRtd
9uLsN8afRKFEHCDiGx/nGhHXOBnevwbbyjVvzCzyDnxZ1LQv8pJEL1m2bzz23vh1
IBf2rsaKgDE2lIXzAUQpkY5ZOFIOQnwQzZxk9hnV31Zzhf1K05vEuDvq+DM8N8VP
45bR1VB+2JSbm7dF1XZhzPtbbnzoB/lbH2JLj8BPndLXHYAtCp+qbQMyRUkYoZgc
gKWPDfh4T7OHUsYSMk5LmYt+A9zn8UQ/Yb+ZtEgXwFItJ+Dl6KiU6Gmo2/bDQFSN
gcPwQUvW3VX0FHGmfRrioOrvi3DV1tlKJHqj2EV6XlOqgA+X5PQ+J/LuYQLeObHe
4VH2anMQsCEc18rfYj2HHVn/qlU0HD/WY8KEXTOMr17yrD+BzVu46wzKKFG+aWYQ
cvFboXPiXoDCu36SkuQ7ihTGXsv9I2fkaD8PauBbposLj/xHwvmb57UPi91IyvNP
r1U8ahaTAtkvaACFSPRLPsavBZQsLkP2SEn5nrUdYEAcT/DXQJ3pKlg+f9RtmA9j
JRtmIT/I9QRHQzjR961ri/xCaYwwYmDEiDQWjFkaT/WfihDQkZuugm1Uefn9GVwU
FFpPK1hMwU/kXii1t8KcuRZvtisbLO3H5aw44HNlXJS45NX3R+JrC11i8HFRZ1UM
kJPfc/qSgoCaDMk7oAnA4CrMmasu61UEPViV1/IVzj7eVRQ7wdSJUzRvYhk1gU2q
4f4AcukZUmCMHZuy53Yvs/CW7ifLWAL0my+tqWMsPicH279WTjSsII8L7HdsPVzV
728tlR9jJIhO/p3MBOYHtjTKPZ7iJX8Mlat2Uq+ANGi6xxT55Ln1bEgIF6Hl87Ke
3th2/PFx5wknkPqNWk3wNlJKsrgMD/18RCf3I04P+Lu99LZO5GRxn8CFZNVuuZgf
6vfkAS9a7j+5TlSddAeiy7mDQagQgHtfOQ94/78iP9BWMOiHbv4jofyCeZeKMpIs
HUMjqm9zo1oyq44a06i+uXNm5aPujkE2jJUX/0+9MZrByDg1+2mpHdyIQrhZcnBf
EAkoT8vN+jC2oRMJ9WEnGDJbD7WP12RjAQKBUOWvzHir8R1JMFSkQbaF7AIncv0H
SsiILYEJBDbSLMtyfNIGmWhZ0GqnN9S/xE/XLC2pBtZjGN2WvsC/nQqXMutqg//W
P08w/zsOY6JOMHx1HLVSDxFNbQXH0dvhIRJ5nxZGNbKPCikG/W85vgUMi/FsY3Zx
oYxWm6zLojBXTKl6IgXYYEEoS76Kj3WTvHzEdJ3wfZr2zb8th3r0g36DwFAbqOOV
r7H3XZtF2mlsu4BHmjSgA+P/M87Gqh7XgzvXMEMayPnc3F4ojD2xCwNs4oORc2mN
Nq1tlg0gNdDzOvGmAK7E8R9yIYkVWUXG0jSc9cUem/VBovU0FsbsWwhPyAWZaQkQ
5y0QWSZs8ZkyxAvs7Hz7ZWGoEEndahimRk9e3Y24cJbC+ROZM03LR0N2Rx9MfRqv
Osil+N5HOLjq17JMpSZ4lAWsR8fdOAZd4xAQPfvjV9AjQ+sHTFjNn328JserUYqP
WXVlaYI89HmmMClC9q+KupqW8590DzdjZtT+NiaVAjpt/4HKszscPfnE6xHSMtxT
OnEyOGS0l2IBAdjaIdEDHco13XwWj26ninlJfHiJNOBUGiLX1oRYwhTLtj21B7MG
pP2DUTP49FIM8xOOK1UphFv6XIRShSz8K4I4khdQkhTERsWUyo50nptSXtpKU5k9
ctLCMCn1xB1QGBcvOYosFy2wcWcpVJ1SWlrdT80Rb9Nhr90pU1ounwkueTsdJ+9a
mWCCcYMnMyCclgjBmtkThl8dbnHTMGbkVT+hza5NTt9ShTkCn4iVfHxL1CKRmy3B
N9pqU97NJ3rIK2Is7ZwuH4nofszzcEdKJUcqCG3uQOzV9CVAwkIhJ0rlvF1TyH3G
SCQDlE8bhIv5bMb5yjzhc7BjgrcQgGL36PwNtaLSBfs4PKxawMEUg8gj4FYfimE7
hLzRGceYtbrjV7jLoT24XX0rP9ihf1snamz3EJxlxVIS6gfgYCCb/BCsgA9B9yQa
xCr1Wq9z561UtxoQIDwPFvecol149HVNaeT+LS+4irM2qIMZUokn5r0Z9IMjiEKX
ft3sjrcPgfrWk9S0More7mwd7HMgRGCfDXrmjZeKWenAdPCp1QsJbjayRKubmGpZ
1lRRoVruHKlb4ZhdXm2wlWvmJ7lEgReJ6g410cUouAOMfsLoNGXOOOvIh27jnViX
xRthp+jR6+x9tHEz0rfLSuRA5CM7Vx3A/pCHcEg4qfv/q/hoq7OBXaByRxBIpDNt
rEu+OTMCpG+fx4nqnXTjLd/dPkPMhnr780husQt7a5zoUawgbbM1vAuNWCxGzPmP
LgSIE3ERzg4FA079OR9rUTn2AQNYJOOGAjJV/c8RdXG4ZMzx2d2lX8YcHUCLOe2b
Cl52RhQzU8lmPq/AaL27hxiC0k5U7MKV+z1ghegsqByT/zp81HxeObvNzw3rzubN
4N2bZYf/ik+jBgGn4wcK+uUm7lJMJ0ToQZ1tF1o6kmwN3js/LbQ3a+h6AmAdFAQx
p2cQXZuzL4pkCL6NzP2CDTL3/PhZaMRnjwEuSfzVLqwfd8yDflmqmOILpzchkAB5
GdeQ5TCDe8PnlW0fyQSWM/Bz5fwePfZWsC7zATUyvE2FythIFnFeT0DyxHYZbt/R
K8Q9670FQ4LEMNZ0s+xGHKQYpRljVsXwCMX5nFeszIEBV649v9LtdRRaBYLozu60
TXkuRsbFMDk7nH4AwHOYHD6J9vmuAGU5SCpWrT+a7eMVQ0wWhCDQgU8/FjDCNC/L
1lgXH0oDwRYbok66UiFlj9WFCwknegNyjCK/62WvDlCpNzXYGtfYwvNp1f3us4s6
JOf4E6qiYasBcJ7GN3RRnd1B5dOSNCgwJPNI59E59EsGyvWJbBoYX/jdN+jXsrZK
lnXHzUr+65JGxhELLrL+mIEpggzB1WaG4a98m/tZ4u7905YWug6XaUYHoSiXFAVb
DOuO0FLsv2ObY9opNkP1TalKrT7PfObvKdIkFjvBGDP0a3Fj3fw8yEOWwF/6ffgj
cByKHu8NpzwMEScnTXqDz7ERF/8eJzgd6ustyfb2cCpHwDNKFEIWjxL3W146zD4h
xUpckH4ZKIjQU4lsZZVHgzfoBlpgiKpJGw4t4oX2+HQJ9S8Hb4Sy2yJKXUotlVhQ
4yZqhqjwj3ojyddXzTqFQGbIAlRQNi1KKDITeifXoDWHeIIWjWUWvfWKZMJtNt++
C1XoyYHDALih1pvlXFGa+7p2KHak+uKl8VKKhhooiCFb1A9OfCnxvnujsAUe5IV6
oOz8YdD51CF+mcdgFFzAX3zkx+a5SVYkfpbOWFok9mYwArI3aOJ/Q2/x6z1J0qds
0fMlzZTbdMskdpYYjpNqqjTtImQCEyYDNLCQMk1xf6NNLFaND9Zk7cyBy3xouL/O
NlBAsQyD6uril+yAha/D2M1i8qqdXcVvPh5c2lTQ929UJxVwY5ATlgAwOXieNBVT
H+I9qPKILJnUe1n1urrFdjkJQIASrwWSjyHYc7DCj4t4pvhpb4hNOBCvfYNnKA7k
QbFl3lrPZmHen2ElFRr0IyNxHuNnQU8azUpohGDOA8gK9bKUKiqbkFXtwWuhUi2B
AriaSdjLbd+iY8j0lI90eoPTDhH+a1hCSRlTTdWp0ibDrGFe5mO0kJzi7xqskFEn
3MbLT4R09KqKaeSCntw46+IiaWw0ae+TasMUAhKT1rkuLZfpx4q3TNnhm07lAsXe
li20AbpBQy5n5E3KsqPiS7HHGVsZ46HQB9S7B0IKnhtEsy4WMFzMCzRahCQTmKN0
PIN3f21fVidwXemRkWL9ydJTy5KN7VysZ5H728ovmRirkWNJjifK8KAl5dkc04Xi
wIv+u0YNu0WgN2xRhMSwNjWkVLOIxZ88bq1PidqhBHigts8inkyxpGCbnd0foWdV
eWF1TgibdAgpk+vWB4Q0QlzLT/mJkp2OZC+xj0bm9HLZDJpD9G1AYFuUa+MF+jqJ
4lGOWXmgPsJzQbXVe25idh3Z7NRBVKfLCjxFQmccRtd3uzsaMkpPmOy3ZV9ioR1V
rkVy1wPpJoTxW8ZMTnzIsrpbFKPurowU9Jo4XqFgNYBMXWC5Ruvflmdh/wGPqUgf
Ucin9x4imeCW8gwENfGgv0zROwJBewfkd4YIkSvP4OQ5ohJpYscbi+6ZNcZY/457
abwdWpBKa2LLxcUQReOdq+MBCx1FFhriMJXgZWxvlkg42RWVW/yBwEHLSex/AT3S
Ku+KCEE9PS1L6t2tyrEJVjoelEv/iRDwux2+ufOFBgYPOvGjfiqOSd1wiQTZOBZ9
VQe1lOlZD/2WUpH6exR/ltImUnkFaC6phwQz7mTPKNAufBaYSEQO22sv0qaUPiR0
F4jO5QavxT9dC4BbshU08VfJgiIoMLKxWYp0f5haWQRe66G5Tu0W1EkmOFEA3//j
0oMbjn4l1/3S78YGoFOwz1wMVmCKMOZD2h/VU/IEckjlVwY2pjSNu6HNsyPtHdub
QBxKdY8gpZfUq0sxiFmoxqiZVAkZF9GCaPoMtF+oPnjaZrVmPvwtIXsqvBdG43/Z
1aAvvbQgP6Q5+JQWGJgj0rmEDSVDuVyIekZInyWFYia+kxJHDBDs5FE2kDPhvX2x
mHxdQ4AIz5REsSLg9Tyc8VsEWQ8pjqJKInVa98dsCFWSJ4F1NVZn0WQuaa+o0M/A
uLAkSzMGThLyZJsO2TO/P0K6RUyydA2Vk0kjKsQE3RS6RoumOd6kBhLSXG1tFrcD
iKRiCm8td6mnfBgPLpEUAnYkAVe+EvuTB7/eMZSXhRphDCCif1/av1UfF1ZF/8sx
Y9qggXLRGGkfyc+wnxcUQCFZcSXKpKlXkjws7o1DLbAfMqG2RoTIgxj+KCwbRZiU
mAjLmp41bMZa6l/J+Ok/p4GCS7ha5f9nzhF/lu27QcKQWGFkjTCsvOdLuEhWPs8n
TXzluxyt9lS3CMTuQEGWSAqu9L7irxlwlBE97uN9LAP7pPZj4oGQN/A5uMjVERIA
KVBionxKVZvMbdzR1wz6vHRREHOVuY94bo+j72rU1whUydj0UZz5wcE1MEYBB5gJ
dStlQ5XbC6RE0j1mkMi5m3PnDZDsrP5djuPn2PVPRJaxsGAPRNCWIfZx2ygXCt60
N15KNjcwkGwcXXCirseTP9/AZhO1NH4JkKuFCsqjGZeNhGphTdcszMEOPgzWGenz
/0Q/n55fsPjiu9loxeuYKexgcuNrC1+QI29/bI5uWdf1xLERlIiLH+DoVssKQFBQ
GfHa3idk24XFgLKY8fGzU961Ng2wP0ycP7OQZWmcaKWg6he8Drs2objMQir/T4B1
YVDOhfkBm0+P0XD5yweD7WJ8M02hbBoJ04mKijFm5whAFV9fO0bdgeZyCnrHZTi3
NDaBxvUelBXwpb2VDvbSQCGaiATsRlpdK05zXCbbdbbwQEuTWlgxC7EByw1YOX4z
JFFdK7V325si+4MTIXNFMIWZyvsmaTo2DG/mEg0ya44Nt4EJUMdOvLoV9cYm3i8B
xHRcjQ7q+HRAkc67HbED/Lu00z7k0Dx8cktCrQLIFp9bIsqiTeDrsBxlG+kAMhjN
ItSTe8B0fR+4uYDlmJ/tS86lxREcEtUPrW7Bz3iPLa4cgqf5u4O3BS+rfcib56N3
a67t9B/UV9bn0ylIPP+Df3pGNzA59h7UH1r1DuaZzgT7UD3Jc3WX5tyxNZF8eMeH
3sm1w2178YKYluxtV3PcpK6yD276oqgnB7Bu8TTvocgCQ0vfA6u81e/jFyqN+Il2
zScF+et8fLqcGdakI6kP2A2E1buv6n6G7fo6+Npxj5UnKCK+Xgf7yaE3u2lLPP6T
lRvL7sIPFrytHJq/IgG+c3YgxzPDCa1fi0qig95vB2OT/mGyvJUS8WVbnvf1/iAL
TlH166iNOj5On8xhki9AFwO2Mzz/2sGXCrtdxVwmCVXwOVSn2LrTioIpKsUKSGuj
ic5NfuGmY2uqWTQIQl2YRJZGg8dVsi3Fupquq5cVTMnojcL6CwlsLZrMeT1Nu/IX
WEUh1eoLlN2Gu7yMJv0nJ5WpwHCdEIsIMee/ZdtXU63AXz5k4Trvt5u2B9uraW6H
dHvcNunB0IoAj4GAVmi1SOuC/zOuyAuGQU6SaqRtrelvBC7GOBXiGITWvgDizbiA
AiZtue4uJqScgZLOKT1+xuq6BHER/1JnA/WP5amaoBZszsi1iccNgS4KID08Fs/t
KEfMDzdv9g0CauHIdv/lppmq1OsliOXdsJ2rbtlUBOAFLGoklQfqqAQiJ4ZvaDWl
tuCfwuzKKOS8V8d99eKPK+NJFK/3o25BON4BffyokXne5G+uNvLX8XwjGcTAgemg
+2QKAutxJ2GtQMu530Uh9fAP6uGdVJ+9sI6WsZL8u7NjXq+1sJxp9MPEhCZ6qnPx
FF4QrlufxzMEL/LfMB+WnBDoiJlkIbAg96BLqPcs3B/K8jWVN51uYoTohfbiE9GX
S/aamt6gGhzMl8x6o5hmjy/UZtLh7upr3t6FXxYPjdYmTEjPsF34Lqh50Ak8JMHy
6NL5oa0NsJ7GaGO9z0QyQbwrWbnJ6CPLZMZ2LIfZJ1dA3mbOmEkpAjEMCWKUpGIc
jPdiCsYJfb5wahTPZ7UlOIktZ5M8RvDLmL987laMg7GD7td5leYwod7r0dWYxI4J
KNZ8hF1IQOnzXF8DhZOZnq3l9dNmVM4kqRsGK+OYw9lqx9ERJEV1vlZmf/IhbaEZ
JuCSyXpuvx72NRkTH6KCNXhu+AosBI5gVXHnZtV9sksrEqUttjR8aw9l4OtCL1Pi
VNzvCUrXBwOcQc2qQiXt76AVvKxKQd8oRqS1BJA/ugUFcmpVTjSUAINyXfleRqQl
/uQkRrMrhslpCMCdHGFPS2SA31XSlRkK/VnwV3VqYcz7oVH0YlfQE3p4RHDNQyQf
3t4ZyrrENqDeiYJXWS7vBTGl0GY91wIsJ0LVClbgv4A=
--pragma protect end_data_block
--pragma protect digest_block
MfXYcb3KIUlxyuFZ0/0OBfbfotg=
--pragma protect end_digest_block
--pragma protect end_protected
