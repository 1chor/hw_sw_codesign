-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eJoaOund9kovsC2/1o/y62s/2VLrC3Hwt+XtHTe9a0s5iy/H+fEoBieSB3ueoCXaBwrxgOIFhGg8
qxrFVYienPao8QiL0afMQ52UqcKr+BNLLewZrvWnbb0jgNPq3w8d4k8GuN3i+ai+7ts/DRJKWABW
a9HhN2Q8EK13HkKfnhEscAyH1A4DyfOZ9IA5BeZEZT0bluW4nvi/a5l4mR0jb9iTG9JXVo/Ukwzp
xFE7vuhrq8A2Q26CZN+aGsoTjFBgO0xafT/EclJD5QVKXe5QD0S/Pn/4c10c3o4pA2f0Yywm8mXu
hiLutOAKHR/C8cRhzqwVQLWM00aCeS+5BBWjag==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17472)
`protect data_block
DBmzkaG6AAIBzFrSBpQ2CE6z/ldBuMKhu0x/Ue++9oZaKIv+UzZwGAG71fIV56x0WBJkbB0MgWnj
G/iorzZmhNAw0wY9cgO6qcotqhrGCVZCh51weV4eiIpd2d6hh300kVcgkVTkr6OupLPUApl/R6xM
cCU5YrHwj1vp/6T+zlEYnZ2C0Es4ynnENCu+7isVXLkxSdfdXdPGCMn6qCIBew35oCnSO0h4nQdj
7McTJ4xqtCvI+TL8S8cSueKUzZm0O+0E+C0Jh2JS5U30V0IBwpC3QV9ac8XyNe3geoDk6NksQuDl
WBJ9s8aA5cnhmb1VfTVD64BO37aJDQj0fyVZO7KdSPDW9qxy232mTnAlZxOtdENBuKF5ZkrH1HSV
h1vXwQyzhXnysYqoA9jmev7sU2sB1dy2rhy6ohOFv9JdXOAK5d19T+r/DstuChE/nJar2ITeIg5e
NnkkNmnS+q4/yWyVKLWNnOra7t/UL9k/B3Sf3jWcdY0xW5jridf+Yh7c9xtA0dTgvy3McQb43ERE
l+4JWGCIkXPHsxEjCDQIrN2+jez5KN0U5cpz6w+kTCY11j/tL9HoN1wgHPZFn5pbKAUPfgbnt2gV
QV0SxVVt2mOSUis9fivJ7nLBbfTH8BSy4dKIb7vT566OD7y6sIALwtLzvn3WeETyETCo8AxMZ+aB
PnXrWuzaPrL37xrwZoE2ObmsQ+TlNAjBzRP7Eb6EoOpl333yCFPtcpOowCM9io23+USDuJxxwS8w
Kjq3zusMmkCE3ZOoYv4l5mpdzOibesv7T7J2W4JlduSKMDpqmMvx/hPsXb/7zRt8ioieoDVHrvSu
Fzd12NtKgQ+f+pwhE5FyvgTVUtxMv4lHGYFXSU0FxfJBj7FeD3vKG+tLUB9or7ZOUUZ4DtGaFOry
2PQyUMygpaBYpxFCMSjha9ZnFFeBYocbTZd9v2hWhDrdLBUuNSayyoeHWWeR7ImB6eRerGlBvNpo
fje9pePt8iZw6tAJItahf2vjpJFzyQwMCljS7Adpm97RPECqAm5j9+Zji4r1pdxAPbM8MNs13JgE
4GduukBO23DmmX6BtnQdkGoAFkLkT+R9coKh50zxJWagohLGCbYvwlnAgWeWiHBWwrcRYUSxTQHK
5B3DKTUPprefgGMPrqjK+pXP7Zu/X6iS7yK1Qu74YyViJAmig2KeB8llk2xUW3Iwj+5vFDrRwhS4
0a8ch+Anex3dNQ0+jtrxHzYrLe6rkDMUlBTVXhCdGA7OTONfYRb9D0+9HrToBTr8he68ckuXuy27
Ye3ae1t6D5HIuJy8Sb7Bmk4689PmyBMRuAACn/JwHGDvUvcrzXoiqitqQO9DgjqhV58gUOtTnj9D
H439Hnhqk6EGRy0SYvueYhDCh99pAFjlGi+t02Icgg+nU7AJKnMESs7Ai1gM8BWv0GhMDgxoMThO
Y/IYH0qxJZc72inymFGX/qdxVfniHoymfirhqMduykiP3qPJJUwwuJO3qJTcctvh2EwuEZhD/Dyw
jVpTTz/Wtkk/d2+lOIAfrrnIMIXVu/YpNB+9ErcQXi65WNmwS+mFfp1GGIC/+e+aojhciM8KB14B
XXfWFnyFw949CdSkkhGJC73DB7BwIgWD5cpaTIzWoEYJOytBhVfzHzlPky3jRHZKymhx06rpiZv8
LfyBFjm+7+4pKW09xgOsjeSIXWO779Ng9aJO7k/dY3bIy0e8sE/JHK6cq9ZT0Vq8vnbMczACSqNR
4r6KHPTZH7Qe9322pWzgHJEnKcRmhcLmcon1UtbB/Jg1LqjBf7DLIAxYQAwVSeWmMZozDs2jhXGw
2+Bm6XfRfmlGXJpmqQ3ktUilLkVdAFQo0MYDAmTVUQN8y/gYiQqMmH7dtsVohQDAAQujWVF+QpbI
tQ11X6AJmWdOHQWL3mn53WEUo2PsdPchaFD9Chg8g31i4r2TtuA9Mx3E3mUtkQRftIaaH7fKVDkJ
5PKiQykG1RjmsCj2CZADSdJahiBE02b1xg5oiLrTBnfxzfLWbuXOSRMLzAMM+OsphCQApDfvdOPG
ncQfdC6AIcWhZCf2Ij0/CnLrjJ5H1HfdlOMVnQPpOEnVRzQwrLUqV1N6lZxLYNrUVmVkOUdEi5wJ
qkKyxLKTG0G1cLyqjAkerMA0L9DHjHOMTgQSdWszfX8cBK/7LfyjlTTpgArqdrS7Brb2gXxPEGtb
ZMa8yBveuKzX0go64TWsmOMsFw2J185s3zx8OaXmnN8FHvs+Hr9SZZGrCq3EG0eKxhWQAjHUP0Vs
r/nt/hOqhX/mTbHH8XtFju+NlT5DiB8mpYkfcPCFEvrOQSWNJnykOlnZUtMTfb4zoNZTFxa4qKJv
0v8QLdBlJfBwfHg9ROshUiwMBh+IRHeJTU3om/helUDWboPQSTKhReQ2h4O20aRTfSiKbqfdIUq/
GBBVJbm8MiUC2DAHK/FG6/VIqPcdRIxaDAJFe9ix95Og/sMEXrEPh9dJCWGRt0kBaQviFtdMWXl3
EoyTFA7OGXzPzsyJ8euz6hka11bWM+hHG72n/IVjquNbptK9+21Z+akj2zyEZv4l9jamTBfnB3qn
m9prUgSfx26kqk7GRiUZUiwzCF7I4MBK4F91x59xUtvTmQPjiBI88H+FtFVHRvhRN1q0ceojqLd8
QsHluuaCKfBJXD0Ir/06nfwqSvEC0CMYjxaBB+onltr79ux+1s7FEYU8pStC0eTi/+kqb+XcGxVo
uO2Sy2Kd3Q7cR0U8p9uEDEN1OU+jR9+VCeNAMSvXC11JZn3aEADIP4MxVroDKWToX53uHNwZsDwQ
LRv7DWv9ydbJkuZK4MmunyYCHLTG0VkoVsLsYe10+wLDcq9cIJhKrX45IdWUpsoKOzKeVBUP2N/h
Tpm8cLNngdulADi/jkiccoc/hFdwqFIJ4FYkHVCkuiqHHnV2THaon/WBuLMH20D/kJu/7KGSpuRr
5RFWj4Ic1aPqLs4QjFJOG8B0S7G6Y0Pawtaxw9L27s19/jfYYvsUmcZu6oMrcjfNc90+xRfPTPnC
nVzPC6525CBCmWJ43r+qyS9IqET2krgkwNHJlSzN9uXkTU+TSR7UozR8CphCDJg6+3zDDTXaLA+0
KNUFU4fj44aXYkX8rUq+thSK+0mJs2nPYdtsS7gFUM0yRDB/cYZLEWEemfACylT/HCj0EvOoiCSW
G5AGa2CG8yzoZI2pKNFeC5FLRv3uaM/Q8YbfnNJFe+Bnjs7lwCjxM7mezS6tIw0Wv2w8SCBBT1q3
cN8KopquuiWIvUSMxPentW2J4oUPBU6+wRY7fGon4xVidbOef26V6i4+cJHlqPqj/7Q4BMNlaua6
epu+m9DRrSwdIld6UYD7SgJBXopzo9fO6ROXpzT837fyz4Gh6iZ5VArhFCPDzDAIu+k61ga8dLR8
JrBHzp39Tx3fixY+P9H+Rd/oVjQjykFWJGRRbXDl0YN4upl2t+8q9hbVSEVrN0spYFHGXnm2cJ3X
I4AQDszmyEVgWKGP+G++VAFnx8Mx6Cy6ZDBawWeIQeYY6rQ2RYfU+Ue04gHHepSXbKxtPFlKYvQz
yiKwt+JTsJgAvalDdmRu3hsnd0rjOdzbFlwyBoonOO8wpXvA6tTBaILvoL5xmBfkhDqDQN70mEUS
yf3xIL++y09///KUiiRAgDRY2m5aO0M2Y3b6kr6XCnhbrqNuYI+z/5AcAKeX/p7zbUSzhwivuMAI
HpEpdFrLEG0xd2b8zI2I69OUjL70zWBcldJejQNpZTWpjmF/UrhpQd+4m63euW3Ij/TLvjLkFNjZ
UM8Y2tuaMstPiMkw0uQ288R/T5TCw35e3/dnpFKEkVbf/5CUp4deWKxhFbTNClrVqlZ3HeYngVdk
XSMy4X3yj1fT207huTlEBTVoo7cDox3riHgRb9oNPcPGit4DZfF/rmMHblH8+if5IMhGtC8XeUCo
LiKFByHtP3o3MLOeqYgUSSNBiGGpKKznu1RKlRu/rq4rttjtKbVIiJwyekXfI4lo/w3JRh47pMQy
ZpF0VccvW3b11RtR387hW0Va/I9gAvyKYeCPwzJeCdqNmpXHPRYxiXYTNz586+ZSwiWmojzohN79
MrqWvNKHtkEFpSCK5ZyOrXLNvhqNFi4JDpFKOzGfGZa1+3dp4RcVpxo5XtSDJF9gqCBIWWjhyWrh
b3rpumKJ5Cyd0nk9e+y71JW/2/cqFG7EEGLdBYXhpXvroJeLMS9WFYJHpwCN2l5vJzwf3aQ67pgG
mMBsKrZhi8ll28irH5C3HyKyQDImZR6hVeZXbLb6apj2AD9/0j7knv5/4CYxDPC/9O1yozobciit
Ma1yqQlX9L3tIqA+Sbnu+BQ7oNAkHSSs7PrO7Iv8Tmz4+AaLskEsAPCxkXAhBtTiTlnGWhdW9Y9Y
336qrupJpt5r0yB0FfH3HP9SmLNAPdrhO3ci1nL5Qebk6z+xtOWFsIJdQdGTlNBREWcUEvmMTRlr
pN7KYyu3gjqHov9iUsCzWhrWuyL4TVLLtETXcI6edcOv9tbKIfP+4uXboE1EUdgV3yQUwmg4SfzZ
21SkiPMcAgx6/Cm6fRwes/7Fkk4/YhcbsqkaUnTsgaL2OAKTer5OCi/XZ2k3959Z3PgCVwvtsGSY
u6JBHzibw8qmsLYEhBUi+kWbeUc5gcllCUmGmSLsnIbI38NZ+zDVTRfIrsoUy6gRGESWU8yRYuXK
ezX1rirMCpPf13ftn0kkkE0Ry5mJ4xkposOo6LUn4n++T2mHRgRpryOuSRuwYykDa7/p1KVO4AK2
2cQjixs3j0t5US1fXm3Hsg2b2LcvdKmfHoBDR/wsoKYo5ABoq5E24mP4GD7P9qTViljBpUMQeroG
jZo5L5HWdaY1gp8rXWRSlcgy82rinZPhggYrDc7sNMnAhGdGtYHjjXO5ElM929m3nGX8XJHYnlgs
yGOUp14LuvdQ5akvoetHFJ0UN3+jzGTik7avfCCL4RLEAXxYSSy/7LLisxHgcoHNSTYvDEIeX2UH
iUjtftBa/dc9vr8UITjImZs3svY58oF8elnU2zgbPmZlcstI8ErZ6xtBVZzafh3aGZT0t9Ax3bJd
30viRQcIJQFtWj3qKvwXRw10y35Jeo79K3ZcCVn/PbruyvzPdcW9jK1pe2/O+Kc5K7l9Czp83wy1
YIAsxtQoILOUlKJpFKZz00DJOwNoWbgFcpJQlA+d66pIP7Q1E7AM08+6ZtNeVlW9HbakJIeiwvrW
lhGXxRBuWRHuHEnSWASLH/6LOSubCys4BndFte/Jjed9JoCMP6NODIBV991aiU//AhWSYXAPnmW4
MWLMWxV4Wr/MTUtIbFLSeRJh4NShVxLTwEBhXx4+mvjMiz/fDOszzC83UXDHewpx0rntpJ89eMxu
HiEPwKmEhIxhU8XHhLo34h7M7lz2Z6+6YVS6eBwcqka1QLLGYYSi8ojNv+XhFeMxvrlM7FHbSgTh
JmOkRN4areRRGk7hAud0+EsNyWsj0pYYKTXTb5Axl9jMnL+acMTEf9EX6or5/N6N7xYRmoHgNHfu
wXmU81Tc9cbHinI/R90fluMIK/dqfHNNnFZ31pG/5IfUHSNc1e8gsOFJNJJWcQ1d11cYc/J8aF+X
OrHO6DtUQqvZ1ZVCkSKfs3E1zjQeLZQYz0oFMwy0dKEFuuDk8i5WbLpxCJtS0hvyrCqoEXHYPss1
4eQmuADHm4YkBt7SbIJvD54bEvkrwK5AKPKpAL9ZpoPiTDAQWBkFraweHoBznKJLPhSvo6Itj4R1
ko+bf369/XU3Oq1/GmYfcYKhyS3T0Hj3eUtFopPzwXAwoC9lkXPIYeJnYLO0/paQYXK8cJqL3okp
duBGRfD9ol52tnj9UWus2944Y384KVj9vQkBcvLT4MEWfuTGNuP4DTbEwBb3/YSTa8E/jE2sA7o0
zRqT7h2H8vOg/2vKAu7QzBxP84l1RQq1iEzC6AJ2vujetj0lR3k/mc005Dynw3B5w4jriSZjus2s
IJGYNxzMgbeT/YCr+fm3QhlJ5RfZKBS8Ic3oefKDzRYLdDUsP60+im5MgvhdB+ODpvLQZRqRTGgv
HeOeRBufUcBTjr4e8mUi6Cnt0JMMgidIa8zJJe1HXYtyo9xER01GpUhJ1fxR7L+vgKRrtmehZ1v0
bfbiacrTx21zj/iExQe2PmtqIAk+CbHi5zTE0aFzjS2KowuCJxYcM9hNDt7dDJtG/L/Ju1zx/kH7
UJ6xX3NkzR0SbTxm9NLTTmzTcqZIpy2kuPu8ebdWewVJQ4RwkDou7LUkr71tcRC5VlE2x+PIceo9
aQHs2JN4oTSbgNv4jxwtrISzjHwUN9yR03q4z3Z0Qj/3GfsRB9PSb7gcvzH/IoA083aweRxA7nv2
mbHPiGlLqu7j95U2rk694kHUr8w0btyyC0Tw4vOFTqwl2D45Otr4LrKuoVFxHvLZD6RlW+lkI7w9
A3ciVm8T3doc5lzjnTgcLD3xZiF2igXetm5+BLFqDQKcw/7CE1PsXbNyODBNK3yLnSVbkcRB2LtQ
uSReNkDnMyoQMSQhhVs4gt340VRdCO3ckgGMlcUCcDb9B0guqvhZyAp5mgugs2EHwAP1XenBZwJg
tq/58yAW1wLVo10mrNNlnt4xn/ziJKoukU2NnpSY8n/rhHV3C4dqVXYFb66yW4qw28VEzUU5h7vz
RG1euiEUMUR9Uk2+Ik624illLiVcnlbMkxQpeFC9pjbGtxgiRMcfeaoK5YisVizkyZPJsd0xbgLr
ieU5gWXm5t6b5uzrnFYqfHs3C5Xt1dFqnACkSkDvC4SY9MaS/zCOhAp7r7R74jWkYX6HmvpfagXQ
FTS0FN6EgpF4XlBiwlJPxyEZ4k7g/9O1SlAkyBPYGMiJsdfKDlt5E/7rYfIK6yvEvZbu8XUTRo7i
V/zsl6xNUA6bVtrjNaM84CswHCoks9x+hjIIK984vXxlXlw24vNUcBJUJkPSU0jcsvY1wm/8eagI
zTGjdLcI7IGkOZaaLz8Dj2nLEINP8dcnoThPctQ4VSGYnSq5kbJJi2yUqujay97hnGQB/fceEp0z
fUCY4lthYpsyci5sQMehPxa5LogRvYymgfDZP9YbmBmo16YdbiGEy/6sJzBt211G4f0fofGyKpFH
IP8eYKp5u72QaFqSUmJqRNYyUeZkwmASiOSKcIGUtAUeWRYBpKqwIbKBIppRhXFNW0dxLaZW/OpX
5b2xT0XB9LT7wY4Bi1fQdm+l8NB/HzASFk0+H94E5nEQ9ngxbZp5kytuDulTVAc8180FpDA/Xxfv
utenQWDRsIRpyIZnc+sIuj7Z+1aOrO3U4pKiTFlPW9mq71FJ0xVuQKOYZ9b7qQjkINKJ0dH2GPmE
Ihlg8J9sAClfPdW44alLb/7f/xbxbvtUJGctPMM+LDaarDQKug5xPV4cqccJ9w0hR664yqiDb83y
KythCoEkZU4X3mzZsVqHkNjoOSh+da/ShtRwDhxy2Fx8WqpkZc5kgztNlkwCfnIoca9C73SflNLA
cozM4r9TADP7f3iGwRH2jndbcllk8QHg/Regq983v5vDGjRMLXrOyFV58u4PPQr056ym3ug91vLT
U8KxEjTYx/Mn4u8Oro/jYUGKGlX9G8vS5Up4eNVb4RTXI01Wzt2KDszGzQdlJMTuKfZEPvTPpbS3
/pDNC+QpXjH28oMA4hwnKxAW/yllK+9rNPdlrh23MDe2dd1kYlHy7wtHIYx45b/lPGQalB0Qx6kP
xyRmg/0dBHeiLO0b2OLCVg2JUc8QhD8PG/g9tE8Wb1FnysjB1BZ0WIyDiR09pIMaqhGvArXPuTRD
W5vx3Oe2rDrirClvQiXKwR5Mzc3AVgOPiYvaNDxxrQamPG+x2FTi8xc4iDwOjy50K9Y3HefjG3hq
rPOei2GANQEQESiFrET0XA81yM4KAS3Grw6yzPEecrJvdXYUZkSNBqedScWrUb6M5mWqccYZ/ql7
ZUL/MkiM9mjze44tm6L3Y8M2JNkDt5on6bmjkQNa6AoXiq9QYogtaivYDGv5MdUILs7FwvCWSmwZ
4SKHtg56YBb/ZvVifDHXBna+NFRGRakKqppeM6/iOhhxwiTqPXfaMHuctJOAleWyoas/phRYjcs1
P+UA8kT/uwrzVzOfgsBsOZa7+shREObCp2R4kdWGGHokQwlSuSlIQHK0pjH7GbL10ezXj3zfYurS
QNFxBxrxfGOy0C8moVO2WPnC2RqjjqxTxdmJIUkOJ/Ym19DyYhZNNlKkosdjrixDFv2wH0NMNsHu
yW44Ho2yC2CgSJffOLL/rjq24d4SQ78s+WlT517Tp4ZVZ/a5fK4pvtg/psCw5DZYM/KTTRHxOjlW
Ie8HDboqU4DhJ3IgcnIB6P/fvnYkdavQcY7mbnTPf/3qiG/ARaOyMjS6pmgrlzefxfxQW4pHKpNB
RDHXQwu6FS4jyxtRhSNF4z85MYctNOdzXRQwHK9k9wbWjysKpogJZYA+rJAliMUxf21FLp9D7dO9
vHjAvOIAXSKYYgoJ/sA5ba0hsEFWS8yAZIRPqwk+Acf5OzF1FJ7CmMVY4oRv1a8P/D/aeMulmZZ+
psRvYRGBBxCgX7PT1DqtJR4c0JzgVvggoWPNiS5n6AGb2eAZijgDpQjT9OuLejUzp8yhZSmK1q+Y
hDSo2AVMY70PyGpJ9RvV6caNHX1/FrO3/7ozsQjmwGGnsKMHVyIFLy8khPb3xJAPW1zTZk0XiXJY
iLgVtJYQJ982srSWRFhwCKrNRn71vMwtnEz+RZXiUbCmFaBmEQ0wVWZEXxtpcx+mlm+ZzF4EI4eW
S9SXdpFmbNM/kkLKJVHo4iE6Wbmio/x8YhvrImTKnxWVVfqMv/IDNUIexo9DYOlQJzS2mBs3JFE4
ORWY3Q8zS4rOhN7CA9QKC/ShfvViIQE33JMa2BnTS+ILJoibLCL+5WZ1iBCZkebPpNqrgbEVFQeR
fo/ZRHXAJnQ4k02J7CT8E9t8o3LXGEULXKuJLZr17oW6mcF7i/ArgZ2gv6BE03LBFwGXrQc9koJg
AVac1pVuZH5M1m3JEnmgsfXJqOWwR3QpOPodhrhJspwKMuSBaGnF4cONBjOdPTU9dOATT/KXwEAF
WP4NaAeOZ6OUB1jPCYkg44TYCpXRbpylwx3yeZ63TGrAA6r/F6eeqfrpGcYZIWHiuXgl3tCB85v4
3V5uZSQBlM6PPhzeblV1JUwqDid7nLGMfGGuvm+oDL/eEQ0lCAdmFcatO3DEMhwJUN4tLjbj0Xg6
v5lBOMwFPpfxwdJ/J7i+QgKdRioyktGPyRCA7i6ljRGdgutT67CQM/asfM4ix7d86dW//sNp26Gs
kkPgRsiIG7moOBqoMz4WaW6uxvcFZj1nC1CD3uchVvczE+FetOlDeywOi1gum/2eo3MftleT9Lty
8rIjhuqPL7R9G4AOESZCM1qW2l755ifoiK+xAEAVsYp7VenPgzu1cNZ0eJdzcZN7kiOGQCBcunT1
hCnZV2Oha0zLUh60CProMFMDe4KVXPx6xpP1PsOfO0/scvwFWPzeBRNBeQvG242LlB+rVsHVij+R
f0uN2qQdMIWtx1wPc11aXsFkkDho6DTWsltolGC20QdZGRKo1PjmQH47Xk+q4h6lKcR2zABOHTnE
lO/lpKpehCbaI53stc6ywVpVd3Ay4/gOVBS7JLZIa/fCc+jaMOdm4+d0Da8RhKs/VScHcycJAKWF
8bKgtTmDl2IszD0ZJE7NZtycWRO6FwKPEWY9TfPftNWMDuWbSXXxuQVP5eAfWjRJhZ01SM2KRIvH
r7xU60Wdp9ugOFz4mNKsN56UvQGTyFQVvrwROUafezizT2qftvvQGlUGPJ48r36+3+o/wM7X6fZO
m/Sh6vCCblmZ3ZLEwhEu/Xvl2OJepeQ0qLJCAKm039cK8F5r7s0pBfhJA9mtXZEOxFN7DLOgcyOJ
I0priyG9NEeQrmrgMCV6kDwlZduUapuR5SuJb+ManZ5Cvm3EDPJiBM2UpW3Ugmc9OFP6Kb9EdnxM
znWlNMeKdIHyoKe1z5KHtjQZ1FbnZHPRibk7r0OBrfxxyW8xxqpMru7edNQys5QBSDF1LsiBWMWT
LJ5jSSuaalRcWKyCo+vTWNCp7hN3fjJ53Fok9s4takghcD97VkEpdHKBgC/tlmuYHDYf7Y7zuVph
v7Ckk9ckSzOGYfyn0+QIcJv+wbtuM/RcMD6rCQEouytmd5GVjMdGv7arWIbatU5M5FuPi6DePEuU
TXMYQCgufjy33jLTfDufgFYyQpy54012acWGg8rUj7mlGVxohW9t7fYg3U06h3iKGSbpXUZlkPcZ
AlZXNQG7It19obXn4zw9JM8qfMC76+ElMNaiWboNzFV/V5GuxKYVfw/bahm8389k1JNhjOwoZ+Lj
UHk28l7KZqZCyz/mcd3wBnYvNzSfSIIjTzq28kyWptA4T7xfL0vgwC3s45/bm3lS1uQ5+14JE6vy
UP7pXA86YZktAz5NIRYr5e8g7Xzd+PrCSRV+ldneaKX+z2xXAM5HqVWgSKD6VKGpZdmTgcCrGOd4
9oKgTH0zNNiU/Jal4OUpfqHumMt5TIQrfCL3NvR7sbrd7Aer74Wmt8A6IQX1QR49fk5vfKRDtLYX
mR6obr0LzAfL4MVh1FJ8PwSuJ5gGctpi1/ev8Jw7ymd/ocrjvqk7BbXj6cZQs9RmUwefbxVegyOt
Re++iSpcYUOz0TyKNVx1TNIBpU/zlRI+BG/YZbaLfXRrfG7iLhCsaz75YbBVMOrrK4JVs6LZVlu8
xWdeTf/jfXTI5pUBtPz9k+zLQdelc1bt8Gq3RLx8QWaDwHRMrv1iY+GkA/wMdchjST2eMv6ffAQ/
XIh5+k0N+je7+fZa1Saf6baCL++QjNpfHxkgLR5amr0xO8VLU96nAsPH7zE2YqgIcXxsjXoaBo38
hlUXOfJoaD2RqzfOnjHs/HGsyZBaIaeiwKiJFWstAK054AYXV6kYvyVT0gClj6xX2fPNpHfzI5s6
4RI7QvWmnGR+ABd5/Kg5T3AXG/0+Fyk0rZm+8VHZaDtWNXIOLSo7XAbMj5owtWSDv7ulC/DOrmOE
4ErRj1l4rW0i7uMxPIfWpVhUDJe5yWYBRN2asR1lr7kMOvXVvO+PpC8HuBF7E1VTE7JfkQuyo853
WIZzCRbaUfvFAeOeeSXQHhCYauPMMemreNwRdxK+l7mohkJGj6s/oZL/s1YHBAyBym58fllON5YK
iHsF9SBMtZXJflhoKLW1P31EVcmWNPU8GCCysLjMy4QCr4Dz8dbTsEztGv5SNTKmZPfrPFbk8KGC
MBhEsjG6EZBGsoWmk2BUYIE0j/nK4RyxUEgMabvt1SKXlOt6K6WNQ8e4Tx77ejG6Hgn5OAlC/Woa
qwDWnkigAAmJ6Up9dbt9NhWz0/mjc+PoF/LvMNSMN7EcZdXT5YwbdNg84TOD5lX4nwu4uUf5rBQb
GsrDfgC/Ae0bTzuBE699DFDJzp94huGirCRk2S4rjOxJ8Ti5mHruv9gzZ0TJHWIS0ZQF/wqAOdXj
u15f/kFX849GX62IIpemh259Pu8HTE7VcV6ESt3i3wrBH3kVgmiOvlpZBcwaNHgHwnndUGxBBP/S
XA+aHbUemVvMl786Mq3yPbTPusNamy/bWvEqBrEf7r+SE6y+wa8QfYIg4vmGo9tlj+ed20VA9qX2
ZFkWgkcREC93USU4VpJoZe3EFAPyaQ581ckt/2EZaeHJply/sHmGSJbdX8EbwDLq1RaqpzMD45ny
VAOCoRS5fNUnn4ZqmMCkmyrFzy98f0Z/SQvs6YvlRxHDxr+mNhpAhsuyifuzzdtCFtgD1zYeVy4x
9XLjeFA7tH3Pxknr2M9EJdLSlkzdmYxFSEEmp5BBXPwnveQgfGJj9ixYs5yFTqOJxdqk/mJWJtkP
6UA2aJKqaTpcHxVxRV/+s4gBXafiXuvWpOvD4g2/0/G7ZRfPj1jcROavPMsVDSO1IOPnbZkzuJlF
BTFXn4toIkkdHWeobuV5EWx45pggRhXW8m6WMI+rYDeFmDsWS1t3+LifGnvB5IZWnG0ok/wl0pJC
u/6VROIdJhPpSbJg0mHNK0PZQMoOHxR+sN5M91TLaHVnVaCrxD92nnFA3CYD+u/iAmunWKR2aofH
TW8uAKmyLN6NeJ0Gb1kM0+pL/Xffvvd13TWJdstMY9LqYMzXqm+YEQ9r6tFIm0sqtohsXuoKJoh3
cyJRO3P4N02mKUwmwZfvxwjjNEQ+klcNmMeFzgcHZOJXL5AU8RBhdVEWb+lVywmIgRwvWhObNmv7
IKm1DiTMwlKovd53FNV1bkWoUu8vu4G9XWJdPlFZrCGkUtkafK8ttr0+YmqbI21dEoqfzMU94J4E
m94c877PZQdAAlYc6EG5NC8dqLNaNhZKK6uWs8FMTa4+DvNuhAKLs3yaMzIOGP5mXKdeHvT0VUZZ
Y7hGefHd3Ro1mF45TgR1NPCqEUGs/kPi795XP8PBDYX59aDL7Qmw8n6pX6fFA1cvhqm2UKX3mYzD
SBiW0Ee6wvrYruX9Zmw9XbSAvCISPlm6oLGk/9l6mlwK/xDeYU9RquSoTbAR73lVWp1f+/1lyMru
iAyh7fL8pIhpByCwdO0Rv5KVr5jfiAZdva/P8MrIE3gieswTLDVg1lgnuSTO5OUwhmrSg3mgXdKd
DeAi4Ciu3w7OK1qjRzlC4L4sX4rpDuU9NGayf6nyI5J3WjvOaPKGi2nS1hKYQnuLDkHQwlbEld3Q
aqoR/X9A1cWG/kdUwShf94PMNo/fHBaUsjlh/YxQIjaRP1jM1uxLDPoYKv9JrA5REuHz2TD7QJHJ
sUZoKhFnBSF6nuSajhSLhmqwEPem+CmhO0dmITQLFmiyLKPqugxJyHEjBZqGPfRPdULIJSTczh2Z
xkNoawQRR2wPazT/z3qWWEWIeY2vbsoyAo3fcqy7k0xcsLg0L9bqSiDV+UaqIB1XwAonhOvN1lSY
oT8mD4GAM0ql9hH5efaSVkoMCh18rU6qi1gUquj9wAxR3v1bmXXmO3+6fOBVAPUKY1kiGwPMbNcN
XO/PMDwRVMDPLBIV+58o0gucWpeEOJH9Aa60w75eMtittTmLfQaHGrAlttFaaefJg4eqj0BIILl6
d7Ql5LafEGnW6kFN9zaIkc0n82N3aRG4hToLipLVIVs//dzv0jkGpKya8gmH3O6hB8jj5fRsJQkY
S5/VhuRh9AtoXhC4OPhu1yPvPAB7T+qkcMAmWNxVlvMWmuRfac27QqABos2+BDjaMr1zJWvpkzol
CYVXPZkt0sxvAbJILbhLOdve0HKBtMBEWuOxXifuQOzqlHZWAfN8o5hfoh1Us/ZFgjPi8cxA7Frp
EEmNsz0tQfpqx7/1ccu+9DSZR4zX2a9zw70ttjUYuH1DHvCiC8e9qA6Eg4TesGe2Ilh1tx+OzrTi
V1j4j1FZOgPTVuBBVPRk5Q5ED3Uo8C6UlcRdAPkpIOMGospOAwTlLBOI99TOsb5pxLeXdp4pFmZx
gN6fPuReepkBL5wORM2pqaaqb1mHDii4LRWBeXfK4nuDmnb7PDreQSBQk7gbgScOgLr5hsVSKtLj
TcRXxJxZyg0swHd8XoxgtlDJ0ml1+FWDMhk0UGWQrvWwe37tQvMT9S6P+OkGWeiBANu4QqyTUpZ8
VmBBUqD5bdy6GxR0aceYJ/Zvg5rlJkrC0l7e2xD3z3VYeg0WKlJ4FO/pXXOk8bW1IWd20kn2br7j
KehSTM3RMAUnGKlrqfAhq+7T8H0eOgdTWYhoSi4jT57wm7vgxu9jYosDS9U3/TTOGPgrsGh3R5KG
y8wYNdVObWeIF8kRCcGyrcW7CBDe+cJHcvtuQTcoGll+GhXgf5MMPpxQim+vTTVldItgvVXGX5XD
VO05fxidiNIEpuROGKZKxNOGw4SySYdpK+HwAKF8xz35yndvRTRyLdGs62zd6AqaBorT+GNIQUhd
I48Gur0A19OFxhCtG+UAxUslH2IRcJ4zpe9XGy1NAGay1DOsvtd4Qo8yszT1hVQ2sjrZKjfROK/J
++a2vkLYbv+Z7RxKLe/BHDOe3Mk03HsePPON9vGOgjRuo7cn9/YGO3sQuwGk1oHBYOxIupLmqX7Z
ZyTKW/kqmlxQ4bz3qR/cnNKwcG6KpGC+4M2zjVfVft5QJtkFK4uZQ8hC7h4DPLcPJ3uRUtfSMknI
NKYWkql/4+7UOepTuH6Q66BGz+u55gcYjzD+65wIcGYMibNdRvXZuKVS2AP1Jx3ZBWzr0CRctAFi
rpj0+DJHuKmE7TZQsAPfCca9WC+zZ75W6TL955pLrIfVYt/ZIAVnyZS1ceKKKLgZsOysDzvslO6R
NcbDBh/PsLe5BV++HTSoaLn7u7dhkXrU9dB+VeEo791XwqT/2sMUvTqmPjtdFgKXA7WbBy5iMz3r
isGTNfJJPDnmb+NA8MUKNh9n1F85KT140+jtZrdYuLfc+W1Ya8q9F64vAo1yFa128jNQERWBOGqR
T8zQteaKBEgO0QI35b1bT6ww9aEfcG3XNmlQknlFa4OUj9sMYDJIJn8a4KZv0JmwKc22AAz0rvlj
ltx3+dPLnNy4TkgPXVRkG1QwZGY6/ae14CvXi3lUs5/kcicxhjNuQfW36aQynrLiwMXQeyrCEkyt
wKGkekD/THIxiVxgG+quiuBlU3OBVmk1+/p4boo9s4zI13dohll7IFiA6coW4NvDkE/swYQk/+ZJ
gIoWvGjgN4/TULxhXgOGxqvcsI6iL+REFvCUytJ1IruZ+St3FXUvnmr5GiYjH4l0/AdralkFiuAq
4Ua9/8yU0ftLxLizd5asb1n/leqlPTZp04dLXzh4d8cFF5/i4Ju6z0HMLAzhpGGKvab0Q49KScQS
MUktIOeVGAkfHjwEnyQVGBTY3bgZfdkET9SI62eQiQFbsVbjw7WRletmYDufhe7KF41ulJMhX2/c
YGlIg5dokSncbOWZaji5V+0JF8ZFs5y8y8e89hyWSqERQ0vvI3Y4pgkbHgf2THr/xcSID3Amhcax
/eaNphIERlA9Sj1gMJL49WHDH0TLbCY1CS/gZqs/cBDPVri6OcBg5yLe6n1RJB1equiBtb9gbIzs
blfwma+a00Z9WoLTsl8KOzKel+fJerg9D9LCl1/5ZLHM6MX2cbnyB7jVfMS1qEqBEE7YtVmdnUz/
gZfDpCJHNTPmvoBxO7TxUpv81mW5V64H79B6zE5M1WNu90lrQOkDVRty+6b5B/psXhU4x1Gk+bHD
oVk9jbc/9GnuDgU4zzsaredKJzXdrM3M6zFB7QDpyF8jd9vBjfFQY/8+qLa/oo9+BVzc/H5chpvH
b0kv6zvQEnvDnpSa++kEtvepCVa6ePgXhImzfu4Og0BbTnMg9ZuP1VOqYhyiES0CcLwIs+ZwSlR+
hV7YmSjLavmjgQczaUq6rGs4zPCKtfHj/zvzvjbWrru467ENi1w7QGXmmUPk9ufirnr/KRiLLQxM
7NKpw+pt9U66fv7rl/3TU55M/RF1WYS7O6/aKOZFUDX2rJuWKGIOyopm3YMukC5B21TL5ModOI7F
PCgxixKwQ34n1HSMdUroLeIaQE/4kwhZKrlhYWIGLPWy2JL0BjNQOoWwRsshwqr0t4EHhND37/au
DE2Bz40TAMaX8kpVaK0jn+6onxeAKvllnfbPGjlb833JfxfV3rv6CO2HmGt9r1F69fHAJ/R2o2xp
SGi2qeXEgIhqm4oPlh9W29SWAcqaeBrGGeL+9IHgiCx6KjfQvhlYXILkapOH+0shtVxMZDSpagY/
EiuhYsE+kySZX3bLLvGD4V+xmweDhmv+ov/z6pSjlpQpJKx1MghQGZgKkYotBwIs97eR6iPqDbZX
rDqdTQwYKlVRSZR8EUtG3IR81j2W7AyksDB5kwAPVrpZWafEhIBWiCbix1NgBlCKCNCa3RnlDPEH
wsD5+zaorMe0x2w/DIbHnKqFaSfjwEvrQGyG5+wdN6NTGPFeeO5gPtfonK13ZrWwtXb273yjBzdq
asmkMA5jp3fBWchsIBXx/JfZIvCwaqWgO2yQjmf5hqtDB3ZJw/ymiZtuXGaTJq3XOnUL4edXvX3F
hn6Jm8WP4VyD5Z1kYwpBw801Ewu4gPGN/aHMJtwJNLugOdTgWLXbgzjtVy4pfYhDD4hyOo4BonWr
qruYyAwGWsKP4dObr50vauq9FsUqr49mMCu2Mk1csLJSj3n97apdHbr+TWzpuvOT+GCOtNJBeZeV
1yWyqCi+LHGI034OnJ6MJuscekBsrVKVOyDZ89oVT7Fe2zxrW+8e/gN6mVch4dAMMvtvd1FE5U0k
rx27Oui2giIXzZK/c6JXxIrF6v0RcwwmvDvBy02LZdti+e18r0aa40R1pY/cDTEFcQF0vi6zI61L
WcIdM4O+V+8Ip2rf6h7Vms7xhNtwxnxEfBQA61tz2bHS8wTDK0vPiFB9KrPix3ne4/4/k8earZxz
c1pIViEPD7u8UDW0Tm4Q0Dwkj+it9oaOyXGmvyRHMMg/r1vR4aRnepOKMt6cv0uYMeRqAPoWhOBN
jh1IEpoDFuD4dQ59gEy8BFCqr5ItKYdOtqjdU45RLQbGIRygYtCgbuytFX7wNUkHW7t7ihzoZYcW
ZJlppdYY48vLY92y88VWWyz+CDZlnrqlDvIj833exgi91nwFx8HZ3N8esn5RjEwjVepBqgrTPlUx
q82wgb7EgQw9PqdUwvr9jVX8Tgf9QfBI3VcMMywXXilBblZRizbqYNV6L/21VO7hjbbWLSZTRkeo
KF9sEpP6vvEYaF1/QdWN4MGPpuMHHFBsitEFOfXrPIvytE1cdGpnBkqfUN4q/gV6tz04BChcD8kE
AJTNSALb3WDUjjTDOsNrxV5OVCsp9ItE2waInoivar0BuoDVxMOlE0tOpAb6DFCNviL4EV+kduOP
Uh//AGZDYFLViecXBpnRzPLLX48rQDJed2bzcTLlcUNbpaNRTPcaoHY8pppyisEFuH1eZPiR2X1B
BCvV2E575UBpVFTQJUok73BnNxESrgZV0usCEnFyH/CLOrKCuJGk066I4q1ylUmM77LFSPGpQ1bD
CPm64RnMsTzm2q9FEU7mHU9k/lcEaRkBujsXAcM+oXu7UxlE+KgNdNVn1sUV79IGh+HDj4Mk2RAf
SEDuegnupx8ZBxmz9VyL18NcK7HNOLQTu34ZqcOb/d0snAmzih78ngujXN5FHvMrG3OM4zSgEZpk
SIisRpttrMaHOkpZjJMqC0i/ZCVBflGLv982GByBxYB8AIOjixac5qkRC9ZJK4pgF5VxTn/8R46E
tnN7KfqJK0fIdGZzf6oqU1jgtZRg07KeDyXHX9kKsL/dxsHItZuMDb1W2YGHNwN00XY+eQQugo9N
re0dffNOXTRX19bhfnG1UU9BQzb+9+uh3y7lq9xBqnP54yXDDDUccc4nNLkPg4b9FUaQ+hcBXBZM
oYmyq2w8GfjVsfI8ovp35N0XojDTGg6w2otEX18U1oXX39mlIVu865GEx7hbeC6mh4YRtkKRfAJV
RHjgqCoNmHaC1rGXIRQ1GiJQHLwatkAFi0tPNZ/4oEeMgYUvgzvFMJGzIF8dQbYDZ5IBX+F881tW
MAhclp4iAGGapcwEycBthRkjbn46n0Fvo+hfyleh7/hWPEU6MEulpuoJdmdxBIfNwdlb3ytsTPUI
DyXI+sf9eWiKrd5vAc+/9w6X+QUySeNwdx0IOLHOfbHrisqUYHuFsAC68VDP3Pa4lol5QnPxzJ+a
FRZTgM/bh2byZ3tu6kRGbmNddXdd75u66f34N+ud7aNI0wyy0B/e8RWa4xHV7mIap3GWAYitbh3v
+zws5zdkzDFbB2ZkNoDelsmvvIvTaDGt0TZi1h+K9R3ppRq9QasbM+cw/UC5nsP10WKCWRlRQUlH
lz7eHKjV4ipaJegKYeFqeYbHjMOHhfauQ4CaTOd1cfhd91c8wKWx+VD3F8rnq5RsM58O2XpZNz0u
2TYI1W0lUFQvdHl8pRmbMm8r3qIF9AtBzKKSFnyiKah4t/rVrE9EVzPBW0S8xml3g2vezuOwM9Dv
oWAotSjjm7d/zIUm0f1Dq782JCOUXA+KAAuGQndUUYWCYOspJ8G+LVbXJuQ0RfC2lvWGo4EZreMv
GwVhipXrI0JvB7Hn5Sy9xV8jwpW+x22hCrBHNKAoewOgWgoJ4uyqTOsEgH9JFa05FSzx3rEAVSUU
+hYBlIz1008o0lZ1v6vP9Pk/0knuASKqqefjfpeEdK4tbG0uQAImqceMZHmaI9OMrWE22kzNS4Gw
9pyErKVD7VfQxq/x7sy93WP2dWqC9w4f5SwCEgp70nF9dYt0zxKpFbxSAdHen5d7bdnvgdi1wv1d
JWLjUfMU4I9vlPzm8aADOEyw8Jwd0z4Uf5C6YyltHffAJthyoPdqltZuIC3js6QxSQHPJRIPhZiF
MsgdeWfxnw++ygz6sE/ru+vcla7F0tO+m+Jt204Pfo6bOIIJvHAKdfwfJUMpTa4P48VN7V/dWC3j
3fQUZqI9gy0zN3XlvxC0HBPaLGVqwZL0OSDqoI0hzL+0V91Bc15kSDzYTO7tuzIJfmHya/lEllu7
6tNNFgbH0CT6WglL/6LR7o5EbhOtCljIv1MKYSpEdgy2IE+NGx37/ewCaVo7GxgKI4RFtd4Ewylr
kT0P605F5MUo1D25iMvI+Uw5AvMEGyDMDBp7+EuLmfHhLngLLkXGbY//iL+1p41rFrqMVMX97Y38
thiqBaJU/rFIDS7oVUusF/MBiM0jdnq0re0gXhlXXGVtBlH0bKGa8Yc8M8eGbrMLeFgd+RMq7hyb
bzGFr/B9hXhdikyBaEZcUnCAIX9HxqmeKW+h6fB+UY8Uhv/8BDPhTzQ/GzYjehWlydJcxXbSUMIZ
6LF/8t5/n6o7rVbRRR+8/q3Sy1jH9ZI+1aeXgd2e17aRc54QtaHRPFLxRVJZ2jGj6R2wJ20YEuBu
szlPNPnyvDEnTJaFVwoj6JpdGNW+d4+Jhvdk944iOaM4MMbd2AaxOt181xlDpeT3vZFbwTfjJlfM
hPo9mh1PiIN/mKJcB+rqYjZbUzScn3qQXpUquq7MWD+cilp+q+XRzFdkjjiSo5TNKdfcvlyATYEt
pSNuIad9KnJ/cQV0OIeSerpmS/PzvbaUtBVrPiuEdSlt9o59rdiPKfcta3V+npk3ao0nnIoIw4f7
TgI2lDmPpfe1IjGeI3M8Ga06rmFSM3qstKSIa0SMBfV6KwNTDciRe7Gokl3lUqrYmEdnMuaJUybQ
nMDDO2MJnt8CgXEureQMhJFaZsXgW/YksE7YWTaltS3N5gZHS2Mq840X17+apWDCuPqTw8tmondM
FJKANebmYLwapfPSmCdCcSp66OUX7vIcgugMDlFEJRUY0taGxUXde53+j7nL8shkxQWvuKgauNyD
2EYzo9ZnzpedyhICyIOIXa8NuY4ISWJd7TCG+s9fT+TCpN+jgACAANItIVljRV/skc73JcvVVyCf
YJSuxsEnn5YkNp3ZSvNviT6M3sBp8KxfmeEZwn7aBY+36AFLpAHFaoOv+l9sQCPrk5XH12ZrT9qV
EIkVF3cSwL0kh3Y/MWmg9C6ebbjfR9PkY99FtaGDRhG03SAbF6QC05T8xmzKlkbbadbcynwaDOHH
PRpVdwA6rvfxJ2ODTYAfPqaxhG/Cixhq8BjJt9aBDkXtqP37OFskGkijD6afZLvBrJboVt/twuuE
RDuZiPf2THxpRvui/vX03SE+jv+GTjEs8m7/E/TbowqWbb+8AMYBlDgnC+5RcR0kUYGXAiFjBNRj
Ca8hWRqb9iuQtQhwPL9jy21CbwSEmFHgNyegTOea62VbByaxgIEI1so5XyywEGt5pIQ5roYWV6Kq
urloHcZPB3Gq4UTMHXt/QYqDeqrT/ig0WuW0ZU3cDNJW9qaZEerJmYvqhoJ/hEq2Knt7lSC509K5
9z7NVTCHof5UU+pJ8oKTIUNgzoGzmChC+qOtT2To5rPhc6ZtSz0lJ9FR8WbNCRnzXzEDmTYpjeie
Kmy/rBnqilSxcNICzIJ0uA0jwB+54O/mgxTaqBfWZiEc4ggUk3zyfVH59QMUrf4tqTakglZsyaVm
qi3edv87W+nBFCBkn0W0NEHCRB2JrWBBTX9oGjUbo5GGRj/XbYlBcLuPLj/XISDicjbLjyfS7kx7
mfKbtvfJJVrtJmqw5H+Bed+TPbGJROBUqOgcPt9biElW39+igq04PdDu+Vzj2gbW32RXXKwHiyAd
rn/iRR+P2tlmGB8mneFqMDeOGqQ3zReeY35jTWjJxJWeUmnZONggI6ajCJbPuVVucQ7LdIWOgLwn
k9TaZeP9FoaIMHXWfMJDRkoMaYnW5sD3TPaEbLFgrUY4Z1B3HtldWXOEyr8hhbn8L7fLSHiDTEHO
wNcuJhYaa5SASjvKZSxbCSHPMd1EG95MPoa6bj5k/M3c5YcwmgFy6ToTfGWrtc+3c792CD+99A2L
n0xOhxZQveiwCxM7/JN6CLJ83cLMQuOeGeTwwCSCKATAfieJyJxpzPbN9x/+Ux8csyfZPJVyBplK
CKL9Im4cYMBuF9uR1tF1T27yhQMSEudNrKWtYwe1LvlEUnVAq93zQfym27rdFo4yAEM8YlQHHx9L
nmuF5ziO5lS237pkRYxs2VVwVJfSIyLTTVIdi4ivJkvPwTHY6F06PxhK65NeHEXLK1SEXIyy8d7K
9iDITXmtf8nk5dDk/kEulmZQfEte2jh2lrpTPQpGXK1NYd7uMw023M0s0c5fArAiec4BoQf/ezwy
sA0XJCvpNGieHfBzt/HZ7gSaeX6mWgWFak1+MXhy6DzjPZADHIT4kqhJpbJUQaynJsJcy5+Dml1G
pK9DqfSAa1qvaV21ZTKAD5/hDncF3p099jbVBeYoUXP29Pr3/D8H0CqR/+DAIlUk0n54pHz4tkzQ
mSV6ipG6S71WqJgXQBQob+uT/8W9Rys035Yro8R2yngLxnMAK+kECEuc7oZaTB9qasmBK+6qw9pM
IE5ujcMfwdKKIDzSnLUDnQVHvl8ENjCl8b5MB35raUPoxjyFFZ8Wwi2smrgOBx18NsTOuyzs5adK
WspUIhHFQr4dxrGp1WPpnMDejo2CeIHSjzcYahu1WMpAXELJ5I7y6QRIph7MktCbWvO9Rr+/+S4k
UbcvjgjaUHe28RIROq6htMU8tahmCLQ5EhVJTkiRPj+b2IHv70iPYf3HA7xj2V0kSIGcOTALH3W4
rXAx+S83zHTXD9al2iq75ljYoeXjQrlQFWc4YRhsYhtfo7p2OPElBkzp4/Fgbc4N6VZg9SErTq0k
4osyALcE/Dn/McPpOZVGtGvi+vEysdrvaWYDxZv7B6UpYIxSgRu9343l30OmYGL/zxgD1pw8b35t
fMz2GRB9SzvlUoF3WeH8nEcMKrqfzCe838bHHdnNeWDLpvWoBGUhZpnxyLBUhmwa2bmuMgO0GP18
MWZy7byOJK1o4IKKue3iHUeB8SF8GsqQhdWspgCQPD/P0ZwOasUsHqrhVMgt8xHF0FEI3omAB0KP
w0INr3ZS57l9DsW8Az3FxipN6f37u3hxicRCxyMnXzA8/wim8PoNmU3yl98QrzEihDR+W8LbrzYg
95ezCfbxWhiHPI+dfCSr6CVtkPk7qEu5RoAjIr5NsKwkABk1rrbSi0lqlTYHXOwMARha9W8mHrVC
Zt5/+lErne86+shSZaCuJ2W+aZsmhpESKu0/3VgsY13g7tcDdYOcprAU6R7H/hA0Gwt4FFhICkS2
PGe7keeiDo0x+c3w5haOEQTVhc1xUrJ4BDijXSHJnGv4Bb6zW6UOHd3wR5UUs1CArMBFnK3u5cRb
ZvCmvvgbv6zbAZtemxGy+cc0akrW3vfP4Xs7IjRs5HxYjzj41bMPVWKSpJu13v65Pi2Fa5bg5q7U
P9siNCIbunkRACZCGMVd+kDhS+WBWO5+gRgkpcq2BQQMuRUk4ufWlcMLyhZxzslCm2+kE0JT+CQ4
ozP4YegtbmJr7O2oFSU8voyH96NpPKHGXW6cxDa+oabwgezkGkXGD77YHpmRsUumjf9p4gFDT6lp
u2W8vSrCIbL4MVYgLBghY8eBWj7qKPjj9ay9XcdtGStGa1HgjWKw9ASIBLuB0W9b7KeWUX3JjtF8
/hiow+sB8AkMAeWTlxnmXYDStjiypjadDmLtKzq9bPRPv49+Le10vq9s8KO/hS0pSYxY5+QoonNY
ckyfDndnvwmqDEhii0fCPJhgYMIqXuu1vOg3HgPWDhB8cOKFjCB50h3bMVMuZf1X75+D9tVTsmQv
xi83MQgO9tg9VpxPgfOnoY7pMgaauYCBbr6VWYvzcmTw13sWtFZjQha/q4HvR4PfgfyOypchaezj
MyC/yAnXC9QVuqddwzffkRv5+NZLGR4GetYzpscyFUJmilE2YdYQTiOTiMlIVWGeX0PiIJK7EF41
NNmOH97oNJX2nG76d5amHmNfy3BcMqZqGBy+WMB8VeH/icQ1j3tj5Fa6X8ptVIM2kr0Ix3hXFVzr
dt1Pucw2ttb53BmoIIVzbZdG2An8J/dIOz9QQKatyQCpeTmM3KNNOw+Pzd+yRR9f+3ogFRAEmmgH
+/vFGo3qpTsQzSm6RQTwJDexbUZs9LIJKUp2J+yPeJ/f10uyA9sav/DszRiMe24HlxR7nUlXp2vz
jgSF8fDH1uZeXPmmer9nV03kLK+1sBSeN44SFtQDrgy8PdPNyigWSY/tYrP5pSzZ6OJT1DNZ8hlo
2qC6Yb288TIXWO/CXfy9rSPJs5V0/1PFfoeQ+Uidn9CMjW7RiZUREAuxJltuw9HtlOSiLmDsN6SB
8BnSXYW/yfECfOkDODpNA8EDqpR8FKdobXJtZKcyovlfH1G07lpRGSOUN7MvMOKHeRvigPmMLySl
s1amKRtXLToru0KfhhEVoGSr7U4a2N89IoUednilku3liaOa0oss2gJuAUNsavFfUGFrjBLo8+FF
2vw2TkUUN6hHePIonZcHkDK/8Tg/0ZZakCHk8qbbEn6fxMfjcZOekQwImw/Tul5vblD0cCvpixNb
rO67hnDVV/i1eA+1ulH8zgxVw7IBgliFy6DR6LUfwoFBaUG8iKYtDXs5VM3AUjq2wZJpE2eE18Po
x8QmK33l6PPUHn62ZfgW1o+qlFuLS3up1YgyEfvUfdyybLdCSOhD5pyrnGBCDmBazS9WtWOKZgY/
EjToqTReHB3erVxAcd2CjcB0qENko/AG35UidNa8
`protect end_protected
