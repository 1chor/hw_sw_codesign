-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CbChLfUpTp8nifw2StN1URJ+oYn1OQfpNRpaNqacv/ikBlbh514ptB58Erf7MI/A
UvXYWlCNMCC2cci6vtnnTgUOWqqUvdmdbPXMI/KSLj2l+RmFz7SiOY3Rmk2nY8Et
LFIb7SnKI1cfcAiEvviPvYPanTIOVw+9ML+lnGDspuw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 69565)

`protect DATA_BLOCK
3CtaJRDXYqDYrFWsIBMr1ItSHl9zxQgDX/+bVREygS4iZavkI1LHt9wdCgz+w6QC
CkfENajHYAMsBWcl8WtjLembe2O/QATdaKbty/AT8mGfxSCDvtrz/QmlwjtKdFhb
P/cq6vG2IE715/01ZmVlJlgnXeUzsl6bKS72CJoF5803sJlgBC+2b+fEf4bJQI/s
idVPwuOLxacbx2xAlrF1aOrWEmdOcTQFCCs2CVGLQSySGal/9eJpm0tWvda1pOJG
GkrXPP4pNP8XRKGW/sb8Zl4vIeswck51DWmetGhe8wWpNxq62FA8oLOk7jUhktEm
GFvxOpgSjCbHJvR2rtunj6FkLG/s1CzLbaLqasAKAkObB7h1OWeO1s4Cj9tmZBBX
H3hFzF4lAhquFyXLTNj5LXAQotPgGW80MkYVFFF/jXRonLet+iLfwYN0Li1dRQgo
d6/501S4JJDsqeUJzhKDe1v1gM1BZfs6oHlDm2OihAVqCPE5Z8LDz/7PwEGO7Tin
EPzNDiu+9JZ83/ROAaVm0QxtlTgmAqqr6l+36sL+u7F7+9ICvY8gZ+Q+XgdHzubP
k6m+HWgOy0p5mpFk3zoFTr4SipTDO0un94cF6QaOpcAwCysmgmp71Z2F+Q4FhUT/
K0Inrh+biHJFw1PDGJdO54hEsMt/hYSX7yErBwPMFQ74W5MK4rV0Dw2rq4g/hfkq
Ab2foE5qNIMo+zIGN8nksx8NW0NEKOBo2D1NHPrT2QMGNfphvXnzIF0ARBOJmDRY
UCsvp+x63UCC3aII7QiOOMKD35DvQd80KIj2IhK8+P+4DzqUz3b/rXPdSilzubT7
cbExkZ1lgF1AmSenJxOVclI9UVHKkiZhq9eAUwcI77ez+MmAm/svniFGDbSDNNtg
CW59voXAwXXxRMdPgU3O0Y65Wkny/YIxO/Bo4yesf409sEOjPLFtsk4qsRZOG9k1
+tVZhYKN2uhpRKjY83tXkH79adcyzrBoWQzDbPpHjQDfa89u9oVEL4WqEWV6v1+O
iOZYPdlVnNuUmpmt7MqlCahdQvbxHCwg3Exyfb783xuttKRmtIvszLdXUKj6KoyJ
FXaAS2P/zRUOna98KnDa+6jse5NaEx4/fOEMQUp66NTyQCLa1AawoZXNRPsJslQz
BJ166UgILxfmaWuYQmR9tpi8p09NJGVGKZmCkiN5xSousqshcILMR5a7x8VrciGQ
A2LJgh0X/6IR+I9kKu7BpdSgHeMWONsUn4YoTjkSA/rYKjvSbwq1quWos8vHv09f
JlWQJ1UJw8E3t0G4KKmbC26eWhhOf7bn20aJ6T8c//LIknE2O50HxOKfg67janWj
KGU7+jMYgyhJORsLvjE3S9c1/YEXRGgOS1IpfEdew4Y+tf8QClU+G28UvVhkTdET
LHAabohVLivjFrMwa0H+8aDmg7h+aGW9IQBAIXa6nNuoxTtTWsF9HKQgtuR3D+oO
x7Xxy+Tnxjz6S9pJ9t/TskMXe1bXrrc9XjvFn/SYEyIX37F51Y0UgUE3suG4/3Iq
jF3fj+K5jo8pMnl76owUEwMG2jn+yoO8K0+9YovvXHPq0qoJbUf8G3AGkbMSh4+5
5P6WWdkFkzeDN/6TWjue6W2UVfZ7gPJh7ysZuGx5PNXwWamj8gWnpuS7cUS2vPqK
xkrAW2gf1WqiKKpdYNZ6smflhUBvTvUW1XNVsQVEec2Z0m8WqMuAMrbAgBpFje45
GF6ZjtWNfLyyZHtTmAxKhrw/R2h/5P0vK3blcHi3ivuG4YFe8y7ZzsFWOUXSpiDQ
zfXYPl9kmsJ1BP49H/H0NwN3BmtzaPE4t20JH8VLZ4iwgHdQYdTWeqXVJsKBfcX/
j1SP37cW6sggsZ1xCCAAFOFtgVcBuSFZjUozcbt0ZWxxbVmPV2kC1B7BTT64TSLC
w984/rhZpwU+pQBTytaVsLuS7vpeH7zKze/C20YviXXGGSCA5pOxXcu2Mrh0byOc
9ha39YD7FNzUc/GbZEx1jzNmxJUyyAbs3K2JFr/WaxSmKRMMeFzTrAJeMqFkCQjU
FFEg04SjCCDaAb6IfQDtlhTxwe9Wbqex+UgNBXvmjwiQ/FfPRrorG4Umgrsz6+F5
6GRYMrXhwu3ehPWFHGMCih24LQ4MCaUYCC98NNlMTotWSdINCI90oYP4CYnJ10oH
qm8zO/Z4AEsBc9jhYT2DpXYqMFOLSigPqwIP4kMnCB5RnvIWSth1FON9BLLu0Wti
vkgeLWWXQY820d5rrKtIqF9dBQ7YHfdacsIhisOmV8aK8nl0xoXReVGrBrJ7g9jU
Iv40oNtE6Efwo3fxxjo8QXZR/M8Xggddd3ugrH6V4IyhxT1h26EPuckMvUIaJuCt
1SIKDAn6wL/OFOeiC2A03dPG1XSTMG4KGJskzwyQXhWcB9v213Okkq8RtAogbIOw
32cDClq34E94xAzoQM0wd7baut6w+jM6ds6/m5ocsz6BY5EJXNJYTodLWGkk5rTE
n9+sJUyl+vFvRBpoaQhXvFX3pSJN8DSBuDuLnV7aVmoSL2fTihrpvYmePpSvboAz
Wr6s6DEjzYADQBIJh8cbs+GywcK+0mibkQaqOFJwUoJt/K6PeEm50m2oVJhCLPmx
evlplthvajSbFmSI5VGFbdFbhh0WH7RxyjCjNvE5Bx9LHIE+VzjQnQji0VL9eL9E
k30jj8JaNmqfzRMHpUge6mt80nLNb4/OvkCK7cZPhgsA0IUF82iZhPO9Iy1oCKYx
qYk67AffQXbpzvJXhOps9FggXd7o2tVV1pYXjO22uz7599KoU8b7LQJ/rx1pcJrx
zdIOg98eURVb9/Mw28eNXu35UqIDdBVyZTtgzyAfNqAC+qWpSqry/Z24CPhywLwT
BlxSUCkVq5+WeEzg/S19NNVGq6ql0KyVJuG2WJhZVWW9Tby+t9jnByHbY6gw9Sfh
cskW2i9hjjTD25kXwSz5WQJNJG2TXkGYmYS5nW5+WZldIjXmYFhCzrlhnsrVJPkb
dgfpTg9YPDyB9lKHmKPWRwKjIvAJigwzwRjz3UAgjMqqDR+jYNoTNnS+Uz6AIil2
R3Wz3/znYe9I9OMIALO9uGNlO16z0fr2xYA5zQhIM57bxMiToKedoEWkZpR6HbV6
cmx4AekJt07i4QsjvO4vVwsQ32/UTCgE+8EjxNIqzzCRTTMuEfkJnfDhRd05qeWj
w+lCfeOJ7MCH+7uf3hL9QAjLA+S125QSb+dDbI7T6DCyX8wQuRF2defODvAWI0pt
N5WONHwyucCB8Hnu1NX1v8UfQ/z8Z1Wif2XN9wYXrFyR5OJa+T097WyyDbKsnf99
ceg+jsWSAKQdLBxC7SKuW8F7I0Y6z5umZhaILjbgwU/5l9G3SgFuzeIHMC94owJl
8r8gpG3GYmc0H/Yqv6Q5iNNE7L3KXb45NGZJ2tdWT02wkc+AZwLMlJfcWj0pffMf
MZKHbunNRU+Ca9evz3ZN+mGWo8E2bd1m/a++y0JuGrgV2XX9Sl15LH3OobMqNlLB
MxvL/AE2Q6qgDwm3h9vAhR/qhO8xnDn9UI6d/rzfma6oKO4aAAmIAjWR+av5zi6a
ndAMgvEcFHKR8hIYenV/chwNBSNjp9YVP4fiIJRxpkc5hqcbMUJ99MVpv9oaUXzD
bXvuwN1ixefHETQbe3NoFXg9ie/V+7uOXFZ2hykDMYtjZNG8kRD4mfX3iECo7Ph+
zuC0IDj2oR/+csecRhjbyShohD1Y5vKJsKXPoC7ruOQ+v4B96APjaXnPzj1mlGz/
vHngvWTlqb0EYiETCPnpDzpVOxlH8CtGvHDZ3+UNDpyOhWChBPCSeBY/xuPR9sC3
5vH+w7qVk4b5J7/YfsXgXkrGwCdCY0JDesVs6hDSM6ss4U4FxGufbdnuK3zFIn0f
ukrRhoUB3mS8+nX2HxQuGEUkxkIZl6tuIvn7z5F6gr7/ouumIPZqFplqJcUAfMG0
mGA/Ya2LS+20cVAIwixziA6hQ8+JTJqbxzydiACko5S2BT3nmDB0LnNaJaOvcLOt
zx1CB1qcXLWcMQ17ANUPF2GOL1OSG0F5Jf31uw7Fz5d9Ynlm/1vjZkzzcGShHnTq
raWhGyodAZtRG/SQllavshVPNUvTHbPNYcztqXogeVCbzYH0ZGbASy3WlXuEqNbd
TfaesNVrjxTcEpFw3kNkOWeAOAlaUfZMoUqsJgGuyN5UVQs05g2P+SfR8+KOK4SP
r3mgH3stDYBN5gW9uOdEWGrOKhM3NBqQM2KTcqxfWRdTOmn/csUfZUth/HCmhJfO
quZcMOza/7CCDl/lG5XPsDvb6I/ThTnSMgLdxh1qTvweczIg/jUXhxdjS+uL8Mqk
NLIsy/I+Xup45NlyeSKL41jl8nzYAqCv34JxaQCYdaSEDqasfNvxWH7IS0ZnQRj8
FKl0w5HwMCyN21MDgo9T3jQy74z4KwaKJOJm+PfM+m5N3VWdS3ohSPuIfjVui+cz
J2VmYz4nJXYJcZLcS8PdDq9uuXXMVVWVZjPjEGE1Znt4/FlBToTTbcDx/Or4JZdt
sY6WDxX0THFgQjxceq6Y8v1yVq05GOd7+5UpCgXJJ26wBziZ8Mk0DeC0JNefXBVo
bQphRPoWKe9mhknOdG4vpU6+ZnDXy0lRueqB7pykN6KjSh06up2Yf4lZdp7X+sMy
S3BRfxQ134ortG/6Z51L2rXK+3aJRFtjhgS4dcjigkH//W6+PsmYP6hDLxiuUUWP
qdlmDWlNs50ooi3M0Zeed+O3tgrHyxPOrtkNAz6iBQNif1jwiOAHrsZQPDP3F12i
T1wc0GCUDJt6NYE22YM/4v16YYjEl5r7hHGfy6bjfay2IEibkSDOVYrsuled2Lp5
SfjvBwf6HfCEWWVxT45ryvuS8nTQBRLMCFlUBzzRDIIqIMq/KWvgiiCyY5VqB29/
iumFVsubkA0nFlPrcIxKfM0Qv9j4g9LEULHOzlEG7dxFVCSUpPj5DyPl/US0Mr86
bwAqVDb5VUx+QsPmY6EJ3Dvc89I69IkSNg8qVFDhY+o3phmdy71esm2Y06hxiMd8
EQA71+w2y8yC3PynbiWhbVHM8Sjjous5bzYYgLCJ6NZP93sVO1Q8yvcuYmlhKcky
jGAyRA0O63mo+GrUYitaHTQ7SDGY+jIPK0IaPK6M+d4fNSSHoJQn3WxdFJXYPGrx
VWspNo5fDudD5m3nYgBxcJaGo4lxTmlBXlprCT9E1Ip4HdnS1CM9XbpAXm7/53id
XTPum4BJjKTpDyBKoE/63Hk5BrDXIltTmUYH69QPztUzm+5XAnJfSf9g75afnk/g
SkO2soIo47OFANfWlBrVtADMsaD63cl4rEP/L8pTON35qqFuX6QBKP7JzWjRtw/S
sgRAQzyuayHFZQv+qWFWzIueOKVP+WocFXQGCwYzk4v52nOLLZUbj+omAqLaVtZq
8Ne54BkRAs/pAKsfTmAMXdiHyf6u9dx7WOmd4Jt4ovsn0zhjOmbH3UP/5gX/4Aw4
U0/k1TzxI0m+wnVCxfMJd2Nt6mvVZ3Xsi0M5XVe+OhJUCd/9TOXapryUOxADtR0Y
DBeSp4ZhO4FIAunVK6lFQxeUw53u13W0roY71AcdEwcfAEoVjk4V8S0iBC67cRAJ
Txc+EgIsJovydBeAwRIYYellQPSCPYYXPS1MPY0SMzTk5xNtEPwb27J7zCGLSN5S
2oqP7jPU2f4tEe5Z2+JGRo8SK8XULoNgwQFre6YvG566DYEU1qzOM39BqJZdhg/1
HwJYmMz53yhL0jJwAAcH/QPcXcrcGbvAzbWqddcnChqOgZZ6f2XSsQEncUTeb46H
GxgKVINHysWoNWloxO3QHaDf71ZxxNBnrqRSxLnub2B3nr+tFEd4o2K2+8HL3scS
yxv7YgeUq8adnrxps3X5Ceq87HVmump4t2y6U/k9HUTbwy+KKNHsaB0LAeTAMdVk
aE1H7GM54EMZ5ONL/r1NUoqwvs4lbd0fc9Ur24x206SEMFtaS7jl0G0RkCo1GJ23
8J/bx9naWBeA+HJ50ktQuQecdwBfUlzkfyFx8Sic0Q2fnSLIj+/DAfEhOGVTdtXL
sDafTApU9rok0yhiexwujyDejP4xsDpk+h1rNnskH5avv95148YL+nfqLtNjqEna
FOt7rBP01cxot4pd2rsTS5kvJzjT1yS+6z2Yno9NBWt9Pks01mLYS5uc71zRKHbU
K8g9VhCZ02f9hqTO+nkMxyLmx7NcCRPW1vRFAiYH3BlB2u8s3msa7PdWO6u7hy/J
XJJtXID0FDtqM+tPZHc2ZyHUA8/86aJmBeqIHRgu7qPmAaNlDzxCYw1QWno1wVUj
wrEwyBXtabz2idMP1WKhTPa3hkvKJcEe0Jm3Iu7WJFkv/b4dgIWyeTBPBZjQEVZG
F6WI20rp4IfIfz9IYRTT0Z527bRJ8IDoOVzq8HngbUhqdUCKvFriMbm3S7h1puLM
MXrqb65G1z1aUct3BBaDwJtDExRXGQOtXfN9PHrAlX3bD2wuEWOBwYFgNl/EY7ah
AbS5n6o2nXmLvDV6B0yiAMkYROEa2S4fMNdcLAizIc154i6XLb3cb84+T7mazuV8
AOBtsEJnSu+lebXdsP1E5iLdEtQCAe/DOS7U0ouY8wbAg6vRGmnwN9buS2jvEQRk
bd1dKNlh/SwBbm/Gk/DOdCpSjEQ4QBeYhNEkJLlv/2hyi6uhmF3eXAAurkgrR24f
Qg3puPNsOKhwRiAjLGOrOtk1IMyXe1S67b/W7yKGUCsxTTgCSHpBMp+0cpk1fq9k
2zJMBfJWrh8/0MuoQLXSkgPvIfJp0B3hWSjA10OdFltQjya2WzAzYBYuvcaGaew1
VRMECIsw2lka9gRSLO3usljEm839vW1hX2tnd7/B05L6TFwS+QnjUv53hzu0+iqG
oUitt44OVDPeNuZ2MSHn44U/qXJMS0fyNsnwy9+X+Am+fCeEo4tu9LOCgfKrmWMo
UHySqRRaOSr0IhETP7V4itbRwcwbGVJM+SOGuIFwwDsNRVCg853TvDRIlFh/ETik
Ex0kf30ElYNzibaQoZmHmysY87gWsmfEX+5ZFnm5kJ308AH2Zj/T7kEEpgsz6gG7
b5SkLponRDXZHlA17qjjxKKxw6Tw0AkwF5a/zl0AJWTU+XvrDbX0EPr4rGGkNu2c
6YqF82Renk4LjuGm0TpfNyLnGgHqrjrb/86M+sGRAk1qi95K7sv9Z6u5kW1N3n09
a68kxwdjnvdJXCLgKRNUSv9FqmSWp3zaT9gt90Si2iJrCe1FCogqFNe05AoPFbj8
Xm+fdXP5j1RfhiK71wHyXZiAkZm9BOc1tauYFwjG5sQjJX55+I6zrvMZbiUVUcYI
Oz6Mf6eOmg9MAlrrgSN3XD5X5G0em1gQu0dWag6FDd5lgBjpQ5Q4Koe0b9z1RVTR
3meN4qPrGlVHNzt91ch7N+2d7O4wMgb/+4AbQzZ++0AV+ROA/iV77D6wS8DpMqdy
mZcysuH5G7IKRq+EKoCGUdwgT/Mrbcn02cUfPreLRu8YJU+Z1nnBUAZUj600nd9N
emxnx9/RGCYGLmag+Lln0LRXvmAW0oFgNRSfvZSORa71mXeAOxguJQlDl1Kqpnkc
cb0zOfqoo3QqPchVQYMpzfqHM1/4ypHRCcBT7FXiIJyMcxncUR4jlZv6asO1k1Jg
BiLRN2yu1Gnp8/5HFEqB8EMj3TeiZHsm/RxHzdzFYpQ2TeQrGNx2jwsfFMGEtI1b
V0dSiztoQ3VGQ0oSKjh5yJhHQZbmGeAISEgeDv2VdDqKXGB4FoXWIg59c0ap9lDG
KsaAraPFhUxHnUPOOUPJo4jUgA2KoWXlALLesSYgACYYh68qYS8nXpQOv33kNx0Q
iay4oSOghO7kkRAjFuD6RtXeh0u2Nw2XGWOgxpcG3s2VxkgR6A9z2z06D1Dv7CcQ
7Np+73dQ2KV1Sg1sYTdFQkFJQyYanTEPe++OSXFoT4Z9cbZ/9LY0Z01BpGUe/JwP
Y8Wiff/xE3uLaZNbbsNq5qUQsWu7IiCPpmCrL2DaojAMjHJ4lnuvNsGMHB6OekB3
CcN28EFI1XumuuQd0U/0QrlCFlKQHKfYn4jHJprNvVFiIvZiDXYTAryDW10y163K
ufzgOFgp37PARLrOvoD0Uj6HlqlS6FNNvbJMWlXZ717acezOAx8NcUmzjVKKocj0
DdzVh0ZaP/vjKzW2UA/FRirEgJnBi+eHO6Mu2Vvcdnl4EbVvQx45nl7z0gEw6IU0
dYvGqtbC5xkRfdCIb7SU74398M+1QXpkmYDvZdV+UKjV4OuLzyBzV7Z6eHvlbu8M
b4AuG+XqJmZ8teOP/FaXbrC/yBrEsbhTDqR2ZcSngyMmnfZz6Z8vAyAoGfPuEH9Z
nEW7x8y+e+tD6Ekl65uG5VyhJct15l4ddNrWXHLQHYGDSDP5T6cZxZhGv41fOpXq
pn4ba38rOV2AMIXIHs6yzY0RQ0+A3zhlMikXXqUpTz9KvtM2tJkLPlWAfg7Wgfsi
wqZDu69wXKdaDgrZnRjW0UXqN/VE+M13DY2jHO3I8s3b39J6n4sC7pgpBpzmtYtk
KVk8DjZqSCny3ueeKfu9WcyPJJQcD/dOKEHg/i9iNDzKwgOz9AcWMQt3LD8cgfeC
m10Kr424elq90haZgV49ZnyV5LnSm+IEyrdcI2klt/md5BdlSz2TNQB1lu5s3sF/
X9pFxtTSErd3tCuHdxIIW3Y5kc8FujB0DpHrAXey/bgL3IhBPg1RHm3wv41IJt91
KfDCkC01PbZkkRC35wBOJvcnQwGhrKNoRr51ypIlg+11NZlCz0voDPkynEocUseO
5d7UKfVwfFdHBtt/xCguj2/7x89nZ9IG2tP1s8LHdcRW30hhMP3h0Nl5kRR1W7TG
ZK0ECpzp4qYz56mb9JK1Mv6JbEj8lUPigOoycmcMZaCOdyndj/1T9a2beh2sor/D
NjeGbTWAsb385x8IFKskCpEboXQ3UnlYNrhOhK30X4n8rgnR7bCt+nlEqcM5xdk1
FN+K3e0tSfiKAfxEvnG4MQRvx9yb5arC0gyPkxDxclCO+XzUEdeuxNK8fNsS/nrE
TlPvG5ZXX7buiAww5+F+GewiT0j67+A1JzFg44B9WgdDBuWcilRS0tedK/fCrJ0d
pGh6My9OCZlJRYV3bJJskxiDRe1F+inMtlPuDs6PcuUqzcHXWzrFYq+Crun42LYO
H+KQvLBdEKkfeVzOqCThdV6vHuhRy3hDzyBnnP8IBNW+dkcYFbgNKNvGREuXouPr
4omxPgdpwY62s4Llgi9QeMZj967M8LY/1D66KVMeV/jwIl0ZI5s7Pfi6bvW/WZpL
WShsxvdVMCM4VY/vmhsRO1CSXT21U2F9BCKEsTdhSCTTTEqoKdlrzwDH7l1K0FKs
JT0I4fQjZCuq+p+jwgyi5HHyMp4LTfZRWXDZ0ljLn0YeR1C0vntkeI6n8Mrv3Tgi
zDdRNi5PL3TzoMOI7d0OSMJZ7D5zY9WLFu02n1OXpY6+u6F8W7wDSCDiT1VelrKF
nO15J1K6mibQmX0PHD+E4o/Zz1tY7e2q7fGFbD1xHIcX00o5H83JK5FtTLgfO4cm
9wET9/YmjAP5H+jJW4cg2NIa8mjKE2/giH2c5EgUn7QY0COi2w7UYXbnGAaehE5B
CttgrtGo2qHiKblDkcjO6yjez50khQNuHMv/vrJ0CAiGK1wn2zEJKZPdYVBkEALt
Rdxsymy81eCFee4NY+aK55fAmU4MSyFBstCweqESrAY2hhJE9xgq5lNQ/JcaB80Q
GE+WOnlucHpqJJNAxClZOa38UWcJR3EttrtPI9efWwhxAatso9Y0C89bbfjdHGQ1
K2cjs5qqKB7NCn9Yz9Zl9cU3KOcdHsNsjPv1LBV45inuDHvq8+ucSKeZ9ePkjZcI
5kMF5p3HK04901UZYW+FrDAz1ge/EyriHM1YkF7Nn6kvPWN3LSUtEVB42f9YpSKk
wnStkc3ffQMPtXnAFK/aNUv91NW4ojEqoz+L1k82cHiRWdS4sUxkN96xZjQnXOnh
RTyyr0iiOLUewjsUrP2nQ8oeWC4++mJ81bp2oShWsthuqXIeX36NWsBdirssmNJD
jflNoajfyWGco338H83RAPQC2bont2atIZEtFMmjClNX0HmHhjSLMZID8nTflMWc
w1iqRxtZ3gPcaJwbw5tcedlDfzMMidXbZytaLY2Mg5IhOzJ6cB9WEMih4LWGNPE0
C7tZ8RvmyGFhBu/oeikkcjHAEJq9jj/8wOvWd2uDTRUFct/z+9CiDuOVvKO2YMvy
/0i3a0lLfbTkGg+SBtp2RUHXKGocRkIB9tJ3OOrvgLRt38TI/f9ydofLBIrCq24m
n1fmzAxQujkppV2wfSgb7p4GaqIEX3YC9yBdCO+HIq637FvlE6BapmjirPnGSLnF
RST507aL0SECCUeQPspmIpjj938U6Rkt5M31VShJ7h2iqtA5zfeGbm3l8OAC6Wil
2faHDK57EuwvNaABnXsjw9D0+CcVzN0A7S82rhbFXbbJDP06eXAlqtAcH6S4K+BN
0Nm/2e65hKT7FaRbffrWhTBR84mBbDMRV1H4WYGCTpFTIUO3P59PliMVbl0is8Ud
3bRwD6dhevTCBfjPkaBUxeEoKCAXj2PW8ouQzFzqPCWe60omla2b4NCZpom9SHyM
t/89sxsi3mLZpdJ/yfKGb4MGeVAxo2/hALCXdOjIB2/Tkf/QXebuLr9kqHSGVAqs
jLyi8JTVI6KQVXweezQjsQEiGY6ZYbFzxSnGrZsnv+masXXjHt1zE3AamCBavdIl
Zc7PSGGuMnywBr2ZQ7Wv46KTwrS7Y9fG7csGjyJCoaWRuBrjZL90ZNo7OzHOfRX3
aZy9V2i/sf12uhOsnRsyPVCzBZpW7XwVEqrHXjVWdhYHGe+g0P7de9ETpNqM7f4g
VOYMZpamzaChlvOOhqI1LPbv6YksxR2weWHlxSbgghevoojZ2PBjnoBh4XAHRxR2
8vtFK49G/hPXReV8YXkU1PSZUlrqkfLP+rHCEMpx7m5rdvVOOw0g84xdEG/8UoTE
rRbhPvw+Y0gsHy4+OiwrAn/BNMbX2ky3HwY3GirHHOubtjpQ1TeSqwoS1MD1/nd3
HGOrSLjfcdy9iwYOfszlZCuD6XYjPBzqSVVW33LYEmke0WTb+DMBjWKP/Rv8K4b+
ACB76ttYKWXCFHmRQzhnqfxV8C1W2/RMCSianaCG+M2+RXgUx6RJ1p9gY9vkYpt3
JCj9O9hwzkT1DDztif8Xz1rgVU0P6zsouin9ZpCq8mguErlQZU8tmfAc0WFLpKvC
qN2S60R0h2u+nKQUCTdjpodqk1UgVEysjZJET13cgqqamJLAxKtk9NBEZga4VET7
WwPPc4cPzUhvicEc/gRyBsBeQLUjHBOCWWQYR55AFblu67BHziVmuVf/09BM9VUQ
rgDx8Ygg3C/E44EdURvWvQ+StVTQtZxR42fQbGPeteQF9F+qU93/Xh2nn3D3Wkuz
NCFJviPB76Y4WppwODv9vC+2J8wZGIZnQB+IPJMKOXaWrDnFGEtqAgy/TLb+0n8s
X7MpIz71EfnTs2ODKN5dcrXTTEKUnp29KUu6mAkuqY9QDeL2g1xC/3U6UHHBFNYe
FzS66uXyIp53ftWLgX29fGZF0DuNnSqrcfaC+iL5etS84zpgzEe3p2uEIqLh7IlM
O+8mqW484VSdkf/fpBEq4qdL2lxvDPHsPKI6/MGL1yZNelGOKK4UXTvDV3g7PfMv
uxdnvoIhK0iK2oaoAzYS7EhxctlWQXLBO82QtD2RtkxItYJvyOQUjyRfe/2FOMGC
R/C/i1HCHQHwdmIYbbezM3MNbNUpx9Ks0U3WZF8ewMJBcVulGoPQWgqQbP+gxt2G
CNIB4RgjIeN8i1gXV3Zb+ji1tt/baLNCWWN6K9RSCw3IQ8ht3kvZP5ggZ04DAG2y
EX1eNd9mWtQasdlTCIHOyAkKFSVVjh9pntVSvWH5p+InlfASrPwiYPy/wfNam5Gg
xEe6YkONV2XFXCS2R5gQ/HSR9W0bTRhYXc9D3KUrqImRe1XlQjS8c3tBlSKhU5JF
9PBRCsnQKx88Rjs+fKyQZpVPjNfjrL8Lk5twf7WthoMZtlTQI3Z5AvkjWuAgZpC/
w+L8OhyijIUAmL5P4e4k2jEW1oTq5sIq0yx9w2UzyRxeOLbwxTWON+7AY1ZhEsDp
ffMBeMtdKVUFlZCjmJ09gci6fJKw+HvoDBnGcytiQ5gJyiln8HSxcNKwabtDr4My
F9K90IAV0HxTWTKtrKPTICYLj8+UeqDbWhiCUVhxpDr13uRogKXkt3SpLpv3tdwY
LGh6ewunb7Sh+Q4Tf9PYadqB8lUdf1pfBEmv4azQ4WvOniQJT8X50y/eUVv6NAg+
pBdkwv4LTgjiX9TRlmV/QYPI9xxeLdWEDvDRizu+irDVo576nSkXPXggumy7qoLk
txffqXDRSczmiItNPL9rrqe+ioAuOJV5oAswd7kuntZenrKI3ykPWdaegAceB1qy
2/BjME1dTmgTvlTaS5KrEW4Azm8KaRc53u+6jrfq1MIlHyOo6Sp8WbgJwAKXcS5C
9F2CnEVLoUWfoQWXUH71yCbcLXWhEsm4InfLQ+m60qFHjnUfY4nZ2O+zKRf7++gx
3iFLG6FI9d0lIVSN8X041qTZxjx1Dk4qgQglagldLr3bqqvNoOsW3RVraAsHofIP
MHrKtMQJovceFFAauI5fgf7WEkeQj9bqpwIyIyGHE3yAv62Dp4Fwfx/fzlxiEw6F
9VCdL70PZ7MfFIrMlaxj0fTR767eiMD5hB8N025uU8eSP5XjVbbGRvBLBFPvrTdr
4T7cADggVj7Rg+MsY3+7J1erixvVvoqIarnuQgIf5YN1BntHLy5Ja4/Hf5cHs/fY
5RvyS4QrquTNC7h5rG7yKpHHiqmHar2lRRx0S8C3iJTXH7lFYpbvZgGPvTxVF7bd
SqVmLVfcTjwlh5le/iDo/VMfLer2yxb35Slc5SS2hUxsfMh1BpOghnzmzltb1tJv
sm6ijWxbepYYRYqOXKhWWxUDHoqAp9OgBhlF5f03cxx8fq53a5GJII44yktMAz7s
vuSfLbLC5uoRFw3eEzeT0J+mpaEs+H7bN2VpH8mXqxC1VZkJixqsr6inlptfv8rn
nmuwdMjZcoa9993LJC79CXBV++KJ9ZmUIXPmhVBQVKSHfXv2w+jMtFMG5ZtQqI7g
Dgn7FoxuCBZFWVDDJoRNBO+0tpSQf1GaQiPui/NNq9556RnOs0hrCt77M4xQ1u6f
XTE3h0+9A2AjQ9wjHVwbbKtsmJihh4EunUj+TPNhOixbqM3qGKHq5bROofZW7bl7
MLP31hwEEkoGLhisOfKUpfR0By4bMatCmyL9nsH+CpXDfl6D14TnHwEby498YOtI
XjWhyDeeEO0EWYMV5wT9zzqdhX37j4A0ANIrhlIXG8fBr4KAsTjcr/5FlDg0ZfA+
fAA7O0UdoXLU7wYTYiRGYiYneGnnlSfzoaRs4hSB0IfG03QlZb8RMzIFhQwaebfb
Irso8pe4vVsptKYCYazMGSDe3fzgVWRSiR8BjZgSPhwuLQu9uF5Lj48Sk12UqUuZ
tPnIhvWq2oHMCA/1GqrmYMv5WR2kRf8dMv0l+PPcNBE9zcL5a/6v5NzuuZTJAUca
NWh1dapwCcHedVmwG5C5FvV1JQMyMWMt9XTIfSvCKRoNAPwxJIOX/G/D55KtLERH
H6iXXAeg0MKu0W7UO1kYP8JkvgNyE1mj8MrF9saGykyU2+sr09kIapcxw0p03yYw
xm03evvkNbfMGwQRd9k3M24NhwzCxJkb5L15XOyCcH4BGIOFFnAvK9lWo4zXP6k3
uPHvP9UUTY2OPRFFPCgjctyBoklm90BMQOy5cc+7YpN1UTK/sjUGY0rQZFCSLEG+
QgkccYlF0dEKC4L1yw2I1KJ7skOlmj/xz6IxFTvWefseMF/iliqyHuVO1sZsXLPu
TLJAJtKx2EJScdg5XSwuIcQW71YO/prQeS9xv/ez8vuhJXf4yWeYX/h+Yr7dfdxl
cKRwCrtJc2Bc0UBM+VT1vU05XoLs9l6RSDXjJSJgjb3l+iT5G4kX+ytZhBTct6s1
eWuT/XtC2KBThW1CG3vNATp5pTp1/dm89+dKp50gLX1VK/squEAC6kANfpSfpWpH
1lliw+RrkEzHR8S5EWSL4zAf4q3eX/KYR1seBG91URa42OEAZkrpx1A7gk3atP2p
3EEy2fzCCY/7gUnMHmR2JPwg/vyvs+FUFzocy99XHWAKnu7Q+3XdkqKVtoAk5PBH
dD5063Tk/XwPBie6TIVdsqRHwPtlHwlq9jk1z0BuzFHdTJ6cn6pJlYFVi95KumEc
+GG5lT5Ms0KQAEZ0hoysrqmUpZLDPExWSjVKU4JCFKJ+U+xceNnUX2SfLK2gPkd9
xtvkF7rr/xKhTYcRnO4OkpefVKBNd/uXkWW3HFSesRr8LQ7QkOsSHn9z2MyPry80
e/BlkBYB6C4VaIUuXpzPji7PP8XcCPbxHXDTZdt0sZScEFWnpEBPQ+alnkrR1yNY
RnAlWV1G/GVitGBKI0JMreSeFqN0G0ZiGGF7sMFGejqRp76Rx+boWhwix3Za9eiM
OYJKnnW+I87TMUnWTuaf83AJ/TABP4QBcDfhb+4PJxmEOA7HRtByZsrwBNxvm83Y
sD+L18fmNC7hu8WB1eiL9s5L+vbbDKXbZhYAuaK8p9a8beDCb77wI4KFfG0VQSTV
k5JFNqH2g1Ado1tOlD7orbyNBUYQsHIxZfF/yLu7S65oPqgOX1LTLv8+9NEpN0+w
Lkqit9jsGv0BFii6pxaL0xLghDkaIV6ngk9q6pnMT8VhDrZQuW3yo8DjrYxr8ARK
fAp8Q78Xr/qxsRQrKXUnVYFzZmOxcuoL6N4PYCM1faSFzJcCczCUUjm2kSdygNXf
w2YbiHz7bFjqs1NWnih7aBNHZ1g7b2A0uz7eYRgf8rpnbBwMqv9pASjGg+klEXWt
IFByFm3X6YxB25FlbDbBduJ1KmXxkr2aE0QNzFSFOLOYtZmlB5Ag3rScDaK4nfVJ
EAxqVv9QYx9MBrbRrQwk6XMUu/7fgNYDfuZfUFrjK9K3HxE0GFAOpGN1nxEnJeJU
XGMd2MHfr4AuqCO8ZOhjqEbNg/9hAuZi3p3in7nu50c919e3skInPUIt2C619vR4
IcgmRUZMzJ/eql2NKdLubtvUuYv5ANlIXAEKB1l51G4ZK3gQx7jFqT+WMbb59rEr
KpXhxTX9Yc7897EsoqNbfW7j8XgJG2bwUqLhNrVIATp3+Z4xacAeX5O+8V9u5KH4
r2pzUnvgpLnxAlzgHkeR41oZ6peSureum/wLL8NTDK6ssFRHF9kCUC5QGyyduA5+
D/XNMx81mht/Y1T48X7UtX8Nx4ANvrPvt2hne/PrLNeZ1kKACUNUxOyjK4+6CHQw
kqPDLE6pughrj++GNLvfmI8CbrlapLFKc2J2rWM/bKPmRQWabpQ9VWCWHyj47MDi
qqvGj/oZ9kFAQm4XtHRn8updD7FkZstnypwry/C40aSts6BwMlc31HrDEwuSu46v
5WSpC4/WbesNr7Of2O9MkCDccuBpL0H6TUS6cZ2OK1ZseZGLAc5l14lOb1gTu1qM
ypZUaKLAkrBGNbTFmep80QqNqUpdcrBSUXnD45hAzEr2OzKvw54PX/iV4toBZHcF
FzMCsvpC9kIb3qhKRr3fARgJpN5yYTjBpfXD3gg7u/0vAU9JHEE7TSMDjQeu4Okz
Q411NqQfmmlU3Qmv2IUX1XmCQmJEYVCPVqck/VwRESKe7OB1RfhTHfFeul2moVQM
bBdBGOw5IZYPPj9tzf+GwK7ILTdWM+no/x1/+kXKKCOOStCOzkJ+bJnj8x1/aOwD
pVlO4Y41LMj5kaFOCqFuRa57mdYendBFGZgstT1SnDghQlhBG3O+f9mxeJ9tBHHi
KjTTxdVCT9YcQwKZCquPVinhk7FrrO732OEU1BPGIRkDfyHw1atlPY6V/vV6b3L4
qLgnQEhNmZNVLpGoIE6qCncLMl6JXh53al/9LErxmx28q0IA2Mpfp65KDD9hK0+O
00bdAHQfXZCGmJrnUyalV44aU0650X1f4Hul1SrGTLBSoGw/NrV8RvPH12ONVMX/
g+QFbUkNtD2M8oRetcwmSCV3ezA9zuQg0VGb2RdswYnPMKGkK8f0WNbFGf/8H2Lc
UT86mPiSv6Qldwes88lP8H/12YBGf3PcBFMZLbHsEqmVBEiqA3zBMoay5Vwvk1HV
99uUbQB5bXWUm7I4eEi1x4JcKi4FgmUKbQZGifUP178ihVZaSn4E09OqOH+4PUFT
ZMJONQMiOGHzbg1/C+TyLxelpS1k+TeqiMLlhTRLRx0c0sQEBUaioTeXmLi6S4wk
51ucEC+YHUbslkLUtpFkQSu70NcaA4TapBC4MXmZ+7jCvJG3P8iohXApPR3GlWlM
Qt9CayJFNxKYq4ZGG/jk6LkuaFgJwi/TJL9lVnwbE6oK04IMreuXhl2pzBcoYM03
NrXHhFroWfZCEITpoU+IWKoZtGiHBqW9vm/63/kOj4wVol6hQkAdP2Pm6J468hPF
5H9dXK64lE+I/NTTrKnhbmFitUfGR7Z4Riji4WcyFusx9CqNyo74TaWMW6I9h140
zn5XuA+DK95DvMXWM3IcmdhW7g9ThfELe2+MZRUwlar5Qfi3xd2iVUvml9uN1NnU
wEdc5cywpdaMaCsMdW2z+ekevlmmGhDqG0x47dFpJ4TlC150HYEHiZkREVaKyvlD
dZxslBcG/ew8cON/6DHohpJgIm4PVELGs8hinMNTGrwIX8DLpodBe81ZUcLOMe7K
yFTeRicUxW9+ab/PQhJC/SZR2eI6KsnqWuNjOjrh/mhX2ULo3aBU5v+PTZSf9tSa
OGSV9uyLlNiag2HJTq8CTfRZVQJEmrSflJU67N+yhgvVmCccT4MTp8vVAAhzOpOr
Ph0binHYvEzdkYYUVxLrhwa3vTcHhFO7AJ69+lQ2a0t3CIybjY/nX2t8dEu4tovO
2DzbWNY+l9N+2t+hkxcLNUGyeA5HaayyO7r6THnpk8vwYO5BzMhUoGRPwR1xHHYo
pc6MPuyI0o9EuOLc0nW8fZCrTmgTFNZQiU22LN2iqlbbHUob2wpP32/znDQJ1k7e
fu8f6G2yHKGuc+wKMRxmhpo+gawU5xpj4xvR39krIhvPzahHF/YjZ1bW+UzvKIEX
om9vFvAC1V0AKXSzX0jTqx1CGJx3Cdo2ILJp46N71bDNI3fISJXj7XoBXQ5aPtip
kQsF3kGG9FtQv6wT+M58ecU6mMsN7pb1p5WJgX2l6l4oC9SHjZtmAp5ISdkbxcdS
2bn5vir6QUIhyJ5yQdSbbvlk7ZZ1v3ODVNf2x68Z7KRaXcWmScKH0YBXgLkb78JC
qkz6e8vA8muVXar2M/HWzY5kKfuv5CokYDTmLkAnRjM8wiVSzZmnagOfAXRnZ7Hk
Zdl6mAe1+TttDhmofcsXqtqNAw7pkfoA44KTaQD4fLsgrzScuPYJPFTwZZpInBfN
sNJvhEXr/nF6S+uwIZ+Kh5Dy9D3xny1ee89sigi9dTRET9D5opzIJUlVFnFCxau6
s3iNunh6iDNu8GcTODizDjcxkayoxVmJ/XDP4/KOl1O3dERP9L7G69fLmlbEptWA
lUG8QlH6kloWyw9DQe3CLTvkW3+KeSv6VRKl/JxgDqx2CCC9n0uNIRiR3SGJSif4
Im12+9w0F/6w7ln1YrJFmnrZib7Pq4KFPvaslkzYZ0MHaPes1uCEv0zyij6enWkq
eI6F+byJakvedxFn3Z+4s19M74V77dp7uF9XR4t/ryDFIWFTqYofp4ZtBIAWNGlF
5OoxPn4R2jnq02mMbKqn+zlNJsdRj/36pCSq9/kZGnWCJ2ckAh19mjFd0WLnv4KQ
EpfxipBzYkOrlhO+jJzzoRtJ9R0FHVKcHYk/bcpQisyXwgJo9jUohes6+RJbhNgu
m21xJ7VcVzNqDF7DohaF+QRpFcTdGW6dFJZ7RktJ5shLWNwLWkG85n7w4FCiZCXr
Us1ti9XWJQkG2uqZ2evBs1LQ+D4oMkM3q9vVJEwhLXjcIMo0kb+eh8MhiJ/W8Ql4
wkUcJFWNungVcccsvFz8BJ+7kFCS25QciS03qDJMA7OOS/mGSWlylOIa4g4WUTRl
Q8KekbEbFVYZRHdIE5K0xgU4EPqEPycOjF6JjPPs8PR0g2/Kw2rVv99J82PwP/sy
BX4hIOhni4iLSKLOldbgSXyd9LcNIxMGM5DUgrHfR54Xa+czWCmeCqJEdn3EPDbA
4F8q40uKeP8/R7elMywChfJOnZSnFuBRDp5txl7Cdjy4SdqU5Gho6/d1OQTXqUgc
Qahz6Z9p4whDD/ea9t6ObpKk+Ic5/5r2W9sxdH8x5ZxKfGjVjbK8xzqnRr17OyM3
dPjp+TbLTyY2QcdrphQSbtBC9EYTB16iCEWOs97VxgqVq9IUbnNjXJtPyCWSxWDx
4oUV+v7NV7J4gzyXS02mbK+Ip69UZeOSb4R3rWD8ncEzy6Vdxhauy3YngGztbHy4
302JZafTrNs8bVk2ueFp53fawcSelwqayHKXDrr+u/a34cxtvwyxMYY8yNZliJ4z
FMcmMY5i3gOfzTxduwcsIIQ1F/lCYF1Gd/G4viWX95f8/qw8lkF0vK0KUNmlT09o
QoqpPcYvHQdeTwB6PgDoeNwaxMKpXt3DB7jZbj7urri9nfbo7QGu4nismEO9dHYY
QDiXqWiWWe36AgcvVNGOnoOofhy1FBnXro5V+f89OotRF36E3J3/7cSnDx6DcOM7
93OlYEFPmNLYC0mzel4ba/l2UbsM+ZYqQt/MHIMmCrXBx3kB2GlQeM+6G1jVSZIO
/Fy4HkIFfT95ppKBLZr1AaYLXN59vL5IBKAD2mldHlnb53FZBEb2NlkH7H5g/Lch
jP1bykK36cDj91zxsExbaqL4M4CcW6P+sABJJF22wxuQIh7eEuaYMFLCQEImlYUv
ckuw5szik33djXL1OsTc+dYGB2oDMWtfiTznT90dJlnObrSb6JSo2LkTybIrGur3
wW4pgHFjY9qX3PHnC1uXGrTL7lXBtrS0DEwiVhv3ul8tKa4FUDMPYJVhHqc0Wt+l
d5vH7k65vzr+fgEzfEoXGERsRc42FNb7jBOyB+iyFm2S81stEOJtKjjrmgiQ58/F
KbTtGEFfC81+1nCc1sG6RO5W5VlWKyas30iry8S3v2Ir+QPennU/UeGtJirgyH+r
D5YqDfrfJzH3LNu2Nqc9OaKds04KldTH/j52l5JjnO+SExorfTiIHkpdDeIH9AHf
8i+fTLEvXIRpKtZ5QXdnYm1/nrji/c2g4avSqpzJMkywKD08PPGzXFTkZVmndTl2
VWfaf2HlZ4rTV//CrUONPsBjMDier/AX+oU+WBZHnbbM6newjFv2T8Vayt1ui2V8
ixKCMqoPdt0nGVr+PsSVD8UHstEQOP8bL+RtamdfkqFSIF7aTnxJWbWGU/6dM4eS
a8ILF9/JPamjwfE6HbofTZzlT5PWSiXIOUW/VCvicgCFlorcSxMzT3MXO7Sy4IGm
5bVx7wiOdnBbA+mre2Y+IvbgWABRKLS8jYT9nHHywF+pyHzH9JW1v2bRv7nrGLcS
ffVSfbK/iHoOg9nqAFzP1iDscKjjJLUMGHRvjy5mN/mDaYyITLnAw51XD+ymLRmL
O9MNOmfj+sZ2st+f5mk37TF5TQaLoG9QYFD+5WmmtwC813ets21bYgdPAzOldydc
KEX296MauN61szR48SDD1JIJcuNA7heZp9D1C+5vItUSPonaQY4RsDHDIRui1fm1
EIcFuLxXBhWzkCrJZwcwv98owl815r6iiKDqQetQHxEbW61GsAvUsxHN4xlIjKi1
HWdylV76rwkYve55v5JeE1DY39jjoyckmG8NFl9L+0/DL6APqPDIxeVjbDpZZwmr
DTVwQtgEL+Katk7nzr5Di36db5gH7mtqFOCbKxrtb7NMTv6Fxbn2h8XMkNiHu0bR
6XqP40T3RE239aw7Aqu/alV74Jce/NK85xUdnMvaz0JhCf/JAdOXxkuVLsJKv4pU
lYLjeCkkH4kzUplDeS5f4wOdnny3yNyaPLYE1Qf5T1eVK1X3ux5ezczw3l+iwq1C
jtaqAdbzoov9QxsJQn/tDKuvl8XNuCZeObGgia8ffqrVjEvdOKkEfb6uNiR0esVN
6w8WDkPTKtOAX8sF5PiGvUE6dKX3kvgAmL5LM2Qh+WOumM+kpuwSO93bGigsASQN
B/4kuQ8UBEXPAQNSqF0uTkzVI9HTk4/i4hnm4vQJpHnSuGb8EwpFE5aPX22HdGNZ
cotEPdt9KJB47jyrNq6UkQufeTBKv+imbCG5GZnfq/dg+odHUZyzBvHkeLdWuL7D
Ugm4Ot86seIIxA3UQG+Zn6O7MC5HL5PtsLieOtxzOPK7d3qJX1DbkUqsNnppnWio
2r1OO3O2MwrTMmlFaCTbQvqIQ0SafMNBExA2Kg13xV23vAy994jDgVWEQuYkwRgW
BKnJbrxRxsn23ufU6ymc8c0ytHG6vhI894SCNMnBt60fdLYep9uxruWelELoUscd
y5RhM0ya/++eTY/rCD6dik+8B/h2tdBQgvzgWJ24aI9OTr3lohhasC1MKd2UyYhf
9SZOw9qra3ic694G9AtKOPykhoeVDRITrZYjcY/XcHyBFvw2QjUoW+EeIuB2E/LU
3RWcvaQAqJw5uT6DEjozw/C6ukcjAA0R363/3lP2tTOvuj9d7rT1cSq0+HbcOr3n
ShCxoCPyNFe1Gqw3aDMIe4zX7etSfvhFN+mivPVwa8qTQO3e1NaRR5HeX1LZ+M4B
k4aHgmWyO4yXxuByPMz5+DYqU9APzFTr8/ef3wugO1vU5HudE9Xo749C2Euov7eo
AVtrprzKoytJ/FlahTh8JRIeAcqvDgMy0SA4IVzu6IxJVO7r/sdtn7wkz2y6fOhl
89hjNbUZReIM7+3y8ajUs2Aka27wGTqx3cyaIkCtmR1DRk8CBc9fhdsxhQ7k0Edn
XxVFMiMvPxP4pIbe3zmhmvHGgcTvbs862zw6wz04rqZMYTLQR6ie3gDyAJMd5OJ5
SJQh5bX5xQ9dUDek7uOeuC7SnAFhLPiwlobbNyhNI6XZgyWU9TjhMWayeTyMZWtz
o68K6zkYnzYqg/qiC5nl+pnF1PeMVjpV+fb97NGuyFz873j9ll4W++EUumrX5+jz
fNnldlANsWnZ/lLu5mKcqKqRDH4jm9QD9AjCDhZMuhBf/Rck/mzXsXU4/eJhknOg
9jg2naYQb66krfzFncTMzWu2biYedQA6UIfEUJW6Ga+JKTHNll6YXODYJ413vcF8
5xowCWUn4Z1hbezQKYGSVs5/Enex+Ub87iRjVRIghtlQqLLNK8+kDper/WGilgzq
6Hpwcpo1kpsO5XIxZh+wLJ87sbCoky4/8Fdjr3EJWZOHQOiFv3xv3CfAt/oRUxHW
QQDXGAGYdg30vD0ri5RMXQcO+sGdswWsiBatP9fBL2kZwvkkz9pyQxiU2bNXrn38
cxkDb/S98BvH4w6H8cm7OF4xULq7hEJYrLq+QIt8M2b7xJk4nr8mpigZGTFATAtA
IOCmksqYviwXtn+HoP5bccpfly4z3bM9sG6PI6ZgwfihE5Egefmp+U9juF/UGzU5
cLiYvCxortliMgGvhuuX5iO9SkA4prJ5G07mRSCyS3CkIkGWYkXBG7gbSwI7RcHs
ZW5QxzJayU04FoHL+6aWogNUFHle6235rFnjSoSMlIF41EeYsqrJtfxOGuN783B1
7iQcaRVj18V0dvnwWHkXFpTzNrWoU85LvFQx2uYpVeahgUn0GWC0c3oy9977vr3N
2KqB08Ogr09TaNjFu3UTNcIvmoz2Mgxx/7g/lx3v4ui/dOskVn3CQsoQbAG4qmGz
om5G8xWJXc/J1LVRugdm1ohdKlh46r8sEGzVTEsEJj581LGnh9tZJzsywghhfVqW
0N7+OMXw5ejwCMePvUpjCFcpcjr5NDdlWI4FpPPOvrpSIhNeSBaPfjignrIJNDAZ
q7dllZjccZuLu+IxoYx41GMy0YFRCWJNzhUh1OuxZrrsDZZJDZxJ0XwUjN3Aat32
lU/CKxkuyj6qslyFFV6jKhfh6gehYJMj5e8mm3095aIbbzvHOSQvRPPcQaqXzpqT
2Et92fEvqb2NQklXPoA0CivUAXzPcPkyYevBV39/m1pP2pSjPP6K6x+4cggW//9P
QlCz6f2RdUX0whWTDRdAUOw6nCxs7JuL23D6VqH0ZVD7IDCU3qCOZGJP5jyAkd4i
2Td2VamvLQm6djoEB1Xdk4INObGu56tUaRq08nvq1BF1vQa97q1GyY53a6YpYdIt
0tw9ai9KJY1wrOt7Kf5C6XRz4y8EYWFa6Jx5Hs1zZW+0Fh3H4sTFDZCrsaJW2aRG
biS23Ap3Z6kssfM998VAn5x3OO1zlDVUTOFJEsUIGpz6MjtC33dlWVzLoEYATOm7
ZYfsaw6bHahicVa7E+VBrGfZNuuxhDVDMYkKeqgXw6nEF+hHwqRo8LvYYtMT9zd+
W1DSHmjqH4zaJsDBKxIEALyXXteN4LjuiomLYreofgN5rhsswVLsgfNS3DNA8lG3
zmnCDUOUIrwkmKsfI8Y0j7jVdt0uwcyrLrFRVfEHDbxX8b5TI/ILyX7sonxK4Jl0
VkQBHjzdPrpB1CMieYGK1UFzDya2QroAtdVff7ZpSw323Qte0neMb8V6wRmTxmyr
2GZq5zbmcu8pvrLVgD63rdwLO6Xp77wigGh5nNnJSA/rRo/CDs6zvavf4BupE2aR
rdpUZ5hBHRez371PLbGYp4KBPPw2c7aiFFv+kGSrQUg9YZU0LGNhlhsXGtk23JTH
Ir5/yIXwvhcrLTmAYrh8g+N4bBWMYHCsCoGwIcAuw1VuOaeU5kpYDuFfHFTfId3o
qPz7zrHOCI5uPwZeSpiYTRkbstcw/GdcMsRi8r5ylfSJBoO/sHit+oxRNeo/adBR
iQNRTDWnMf6qzZ7yHGlZGvuHIDbwVdBQ4vo2DG7XOfXzRlYPu/eYZXIRcjsSrdFn
5pdbX1U5OPYZqzjbp+ar4CR29QjRK14YhsMd7+7JnfBGOov48J6pdaL9wbRUz12C
b7fiDn8X2eHu8v92QNeVwC8W5DI1qhbUDSCcmB5DX8n4OxeZjBxHc4B/oo48ug0+
Gh9+X4Gb6ZrFAE12H1Oa5pC65EqVu/ONqN+U7Jawn9rncKP7B31g0SmNVYBZMaxn
wjXno50v3CM5Ccnkv+C6Tl+KI+JYMvlwWtQazrpvWIa90MUNUGUMFBgh+QAptf+q
cpKY3kRwbXemFYpPq+/UKBVVe3KmM/MGJAwnvLDojQQGZkTaIg7Kv3mdgJy+ZjC1
KOL8ICmAlGd6Ov6nfWvr7V4cuuz4HAcgH9xE3iELmoKRMquuXPw5rD8SoCCVHEC4
r2QB6RcjLsh1HlFJy8LU0+qy69r376n0dCk/9wnlpJYycT2A+4FQuM5l2w6Sm8Fu
SISnrQ4KSKYX6cI3teOxMpF1/Au4iQNXqu2b1ikRfF/NDxxF+jqcIAcy7YibDSYe
jlV4S7U/aaBy6XjgXhG04xc6CzZmlPxysO+Ac6TIggnUMfD1M36KluTNVRazvAp2
ySchZTEIJEdkdweYq+wcbsiFH5pFVVO1y76bxRqBBchMr50RsoqXflwXrR/Ig4X7
9AT2V0mOC108FgdlRqkBfPnOet1ekcwIxEAdGO+A1tumm/SxiCBVSElOpuqDEFkP
AdxRXWqNnvUQr8WXWNYPLsc+G6s5h+iqVKBGZ8wlQKYWiF4Dap+jtrQ9FD40OFz+
PrsJnpASLoYTEtue6IoZzQMTGJgY7oEbqZikN4LD+xZxwmzaNT95aYTlYxgf9I/0
XqNBMyVhUEU0JANyZcyTHWQsf1yzm+wE8sTXXHOyYIL24sGv95/ZBlteLu9lCpow
28zdsgsBYzselp0f52rajb5ru01B2vh6qqQH3N2s0XrQwtdF6IVc3mGR9XT5ZiXD
+nOq0uqXmZJjRKL9QsA6aPDVFis35/f/e1FjQ8eQhxA85B+o3qhNJXZjGkJ9ZgoJ
elUKlIlwApf1JIoI/bUOX8vS4HfODTayjr3Jpk6SWEpyyICon+fXmPFSyMXwQOPg
7jTbCy/GOpMSHSjhSGrCm4KcCa5+dHVd+S7lQmCDysKcKp2ULXzx6k/Ov7VyOwLa
NBRHQTzA0apqLLN8Z+O83lHyxclh8kX5G3ud+qyTUvuFpd7tmOMRSjmJv6lIUbOx
3vNrG/cG69YQ3Jrppb3eL4+gLwxObi6R4SafJjwKBPdAChOFHbig2K14QPHDWeym
UIUba9VNS1t6gvI17tW6BjhLn09ZCYwLrY0thJNfgyGFapclnZP2iIKQjZtkeCi4
GBU1vOrx/u1RHCPVTIUQEuRKOMDZWz9F7LJ+FhUZU61VUREd8g9n8nnSmmBUmjkO
hecG0viEEJRZ3rcYQ1L/TYHTT4clxVDyQP/kSl3F6HUXBY2lH7e23IYkytyvkK9b
OtP055OEtRNDaTLvptd5I65wR/mVr/3KLC61C46uxwEb01VClAgSls3+SVCsbSPC
KSIvuAX3h+XHtN/+MIGsdYajh3az3i3g91OKrIRDtOGFm6vbcuNQqJ0mF6pZdKsr
B3iIdQ/PlsS8GpBNkFdCRUslCnFh2hIZvtuz1AU2lr5Q8ewJOLQt/wGSZ5v1t/kd
5aDKMMySgxotOeBHo7L/GCdBDbxNig3pBCHf6DfTjIWZ6YJiNtr74N4sZWO3aQvb
rqIqvsoT7JFFxv+eALq6lMH1zeVJZtgDc4A+ybM5pFWiW7ld17Ilt7k736ct1V1v
meupIZuCB6xoHXjniSYhXuxyjM0aKBESCxaq/RLha5CDk+d6MMBipyrx6F73J2HQ
SZgef+b0gCSY/rA6ACmeprAdjAq/MOqdp82EJcpDualwMKYa0APtPHHm0YT7RaEf
BcGDNz9DYjpmJOuge9PXQ/Sg7xHPrz7zrExf0buhtC29ztzRpvouz9fXLDzAPAz8
p56KXAPz2oN4wYW2txvmGCYg4yURdeC6EKauDNKEdqmy+6GKaxl3Duaz/IU8qSL2
KFEMohWADdgzGlci5/MhrhmJuBOsPP3+bT8dMf6swxg0S8eux/MFTqfCJFxxaiFk
lJWrVw+85HMkBuPF3WKTbbEVh3ittDS1+2K3uZ+CL9O1bxxfYzaQ8SjkThtTRDhR
cpXLpmtNOnJPtDRm5cpxnazzTXiveAvRmZvO8J2UbN16wndvEWbtDq15OSW4kHQp
9lblFdZwp2QCLj9JgYX968DFd2pFS79JcE/NUyRyN+4lt+5OUAWmWSvucaeRs1cg
LThbnkV5YGupn1ykjobB2SQX0ehyKXmAZKD91EG0KC0GMiFWHoGXVAzJ+Lko0MDv
NnKlvLfcLkwChw1Bm6PCk6pTJ7NChAs82yCXWxC7MYEuDtCRofA8IUDDMqGXSdff
2ba8iLrKrS7UbpCJPWMrSQ3ABtg1qjBsUogjYvooFS/i0aNkQbFeM3VOHcOTomLO
9rJpYVm2k7rmmOw6eOgAF4iQZKQfg0D/DFINwgDyHREYN30FZVrApQ5t2xsVZMaR
Mq/ntyLhfjrJAo7396R8b2QAbS+x9nptMpnYWI9MIttbo4Ek9eg7zOHODTaQFyTi
jIc9m2C+iYLk5DupY5jygs9noqJEKAXkH7HFZ1w0e+I9LbuJhfpg4HlyEeE1o0O8
CLm0cgHidoYMtbK5Yy+nw5lNBVPDxJidST/o8oyyQVl7TdolBS3MAS0vtdsVFbKk
J0QOUQ4xloL2lXS0UwH2x9kdjjuxfUwBEP795h0uCELu1wV3PvItKUzwnJmvVAA7
zsAxy+Ean/iF911U2Tp7CUSuvD5REgc48+KcNiKm8lZsHr3lHA6v+9Ro8o2yDJFM
6i992Nysn9jXWlvV1ed7dl7/vgGkAiJMcmZ93EbUPpejR1haaiWRavEP+a51MoKX
qledmPW36v4J2umRZhP4p8t1VN0ckwOUH/TcVzR+9EGQwRf2BTTlWFZNxJLKsNZf
Tpj0N8E28dq/lkzDwIxeW7M2KCkKL0rD1wlpuDQ3qlpNpVLRzxdnAMWCmq4Z9EvY
5etqTvRGIbRihSLp8pejk59rApqfJAkUqiY9vGkqI76eSUUXyTBoZih9QUhJhRXr
OmJR/Nm3qMdqsyPxlXJxy9Fj8Fwyi6wPT6QhZEnufKUV3n2K9d5GBWFHdJdp1FLe
k2khWfJbe4r97tR8V9C4PHy+fpOxAHZbiBoVXUCyH/EL9WKBGQ46LwtQRrcl9/eZ
TD154ceWwXDuzjt//vR8RE9pofHqug37xNhLksPc0bTFGNd1bMFPz8GqUti2xist
DM0OXM4xU4+rrm4UMdy5/5TmHtTSmbX4hbjW2mlgkR0VZukXwJB9+8kvyOuEIyXE
oX0A65Q13KV9GyaXSZnuYJ8qGwT2vWSoOec2spNCIoNsyq4TYgps29Sg19QrerAJ
Zam38owZfX/f/B4HYx8rFhLqXp0U6wrjdc/UKqsMPUD2TrRnQPExpbXhJ1KL8A1S
wnH9pVHCBzFO/iNaypIO7FbiAJB/GZkdqccU2+hhV/YmEd3chh8HTzeRw5Oxguem
qpaCrk0PRX7mR69ZBRjSOOmH3AEduEbCIOEI/IjgeEjCxOazzPwvx8LTyEYRtptL
HqwyPHWceYOLPethxv450Oc5foy9Zd+A+IhZhEuOek6fENDvU+dsKC2suyOpHQh/
E3K9Ng3uwcDbHCMG+satpcopnsmAYp8kyotyfnhzuG3EnUTGnjGC/HNNQZnAq9xT
tKEicK68C2czx+JvtIjAAdjIz8PTYdKBVj7qT7l0WTXMiEvqlzCvq+Fi3RCYmjsa
o3EgST1WfGy9xoECY8Txwq8bdmYu3f3qoa7auz6/+GZ9e45mkaEHIF24gWwqwrqT
rClMnKc0YUAzf5HNemqu3VtW1qKy8vQmkMS4bIp9EcDX3bsAoiYgsLQi66VyMzTz
9B3cIVX33047oXsXd6bXDOniYSoavahuDl3Otq3oNj6CyXTX7GVsNJIXC6sessvY
gAOMQMA54xmv118hHe7VjHeu2zbb7ZeYbnVc0MRivIH4c/iqKVkEg7HD0B3uNExy
VFyhh/4hGXp7+DuyfNy26YEo2/rr7Ms7oPRGZkp7H3GWSwkoAJ2bJ0VfFrKiYdqC
CcyYw/1UyoU9h8amhl3I8p9i9YbD8FaOBwLxUHPmIuQ85RAowiYS1qJXl72nuEKA
vN8c/rM4vBtfI9Vtg2aWKteCaqIOPOzo3FXhpiCbl0N4kAGsYpYOqy6EY2WAtUor
Zxj5PUFMJVCgMCnKuUnuM5L8hG5+3X4yOHii/VgTOa2hZa6AZFod+ozwU3xa+PAe
TSFDFGRH7xbS8RwrapuxgZwb5+Kme7lJPND/ctYbZUBL3DRJT6T8JQxjHdZWVAwI
Q5dhgd64vweRSB7EgYg/6dCrRXfLas7aSxXVFAlUNjuaX2w0vHqP+MTIMjPjvJH1
dxxb6Vt/9dmcYvwje2+JHaO/1J40hLCNHhtIXHuQO+7APLaWqcRwTvWfHJ5O1tE+
IXbzNtkduYi1AlxU/axYMC2evD9BwIl1CTWYi9anuAMZKX2gzOrtb2wGOfCC3oQl
DmKPN1G8FbYVEew12PFpBMiXiozeTDMGTWMUo05TgJcZljmh3oBmCvN7b8speqSd
s8GY7ICPcKXogvEO9pvJCEbHvprcWAdkTu8X9JHFfGZoCa/DADmJAZUdLFvGYkWE
DO5pgLgcsvnw1yPBe94qogVJ4lbWICKuap3B859AbcFRKFETYJELxNVos43VoWQq
feHIgOGre8ikTxT3uSmgloSwNUESC7pNVYZbLPVS7o3cYH1k1XUCMfRCGo5p8LeA
IyefK/so5XOBugYdfSWq/u1jix7mmb3yGqFxfA6R3zHtyrSDaYp1+V6Qa94mgxFB
Gu2zYuluO99CwNHELA+SuJffZT8cZsBfDXP0i37Bs0QVhATnzDkdmSJ6wZgMe4ON
FO1TftgEMXJ/U3d0Fz6SyCimnEVTxeLtwMOdSbQ0iqYFsNEqb8paUjRi4llb9Xrg
GfTTcrNj+cN3cenrV7Egou2tkKSz5Wz5EG9nNAjH0XN6DA/JZNQDVfgaG8Zehhxx
cBBjMiouHAid1hiJqOtUQGGjdK7pfQtj3Ss9wacyyVRyVVQ+/mAFi4cIihzy2ZGV
lUytqYM2XS5NwB2pq6hpvoFKP7s1s+kVFCbyD17O3yaQFUn3jAsgO6EdVc28Ebtp
IHnGEaswbgGafNrXzuOwoyYqu+I5dTc9GAjvOV+29E4VH0eh4RKjTOmvVeo+vk7Z
Lw4V3gMWMInYChrj0UwQihTNMLfYOSZTPnvViMQoFfDEhTotiDZ+HN1kP5PJK1H8
m8Sr631HbNBRnzsNF9f9oiKPf8edhzXzGAqDLeBxMtFa+CHZVDKfrJmeMavdfgw8
N2DCT86cZAVJuauM4YysyNmLAc59CnpL/Vg6UK0lCipK3w1fZ1IEdliyR6Bs1D2X
3gJoQ19RMCPtia9Qtg7r7Huw1S6WGKDgVFOXAaJkZteXGh2fyBbZSZzLICv8c6ZE
Q3i2sDEJVvP2yOzEhADAoJimpK7ritar0V8Z4pC3Y9u/RgdRaq0Ja/P2QB4oEv32
fJCbbr5Da35RTBGAGHPA3t1qyPERC/4OuQ61ik1fDv5RUsPhziHzJaxIAfDOvW8Y
21oRzRtOlvmD5ri9PhhoDL1nyZGqOPhpQztEa1Pn8G2+sPVDagagDuBRh3CABur4
qFTD1OFGCQ4L3uWkM8MslVVGn1cHA9J5IyXIh8UuNpvNFfx4pAc7QIOH2fUjlEPB
JkCVweVy+/T5mDF6YjhzVl8WgKmHsi7UoCgK+NmPBWNlxSMAtWCg8M1SHHDo2sFf
JYr16IV1nguroLuJskipZvfxLvQAzkRhiCvrAT+gkgVpE87FWfHlqQO2+HmzDxQq
dgOdqwkfbJCGMZem9jk2wc/z/0WUACDr+INnP1HbpZYhLvCQW23VCbUaUCiphRsd
rVzcs/XQompn5S9EA5lIWsqHU19PxtSdPmX6UNQ9mVCUoZzQFjqhtREakcRyDofg
wMJuaCUPCm3zPXVCNaDfiRzvWOjEfT9c2jgjSiweg6ymmzU2xzee+xd9tKQc6wZP
u08AD+C+TW2nklLlskI6bgE1YPRw2v46439fJYL+jRYf5wlaGOCJ3DlKEMxhmN8/
cBCqjFn/eWCzaFnsfTI2dxtK877SpSH3/EVh9VHjMfUoqcyKrH9K3ogxVUytIcTV
EI1no3+mEYNsHC9yFN/rXH5byOAYVQuNmxlTE2hGeKZmqQLY4kmG/zQ6IE3UyDaC
pKv4m2PPynYqDyHNTUJrluUfFo0AEeKByhf9aHBa8c4if/27rE8SaqRHXqVSF0CW
cxyTplTr31C0Wxwc4teFuxVSd33OhlTcGFKIeGKFNNrV0272YZiNs66kMied5BNd
23Vnpyx7i+qDMxgyso7lIJI0C12BAOwVRj2B44btbjJuNXk2Y+/CrcpE77FjQJ1v
NOWXlVIApJdJSHTZV+T670UF/7+2ybwrvhGeln27GprpP2xEAaJ7p7IvSQ7Obxm6
oTrEfr99dmXBCrSULGYuWNZqRRqyQI1bhInmo79P/6YLrdrcwBZZYuTioolofZL0
moH6QmH0o6RnXiE7ZgBetQmw3VR+CQTBob9C5pBfE7BsTe/a3CEO85V730104nsk
FkvB5DpxZIUTMTxT3Ccjk2QGJLNtHkqVpErmyrIq26nbARgjOOUE/Q+3UA42kq4g
KovMSaMlZij5X/VVzFsvjnDC1iNhw3jGoOSiu9/t8sQFgQVCKAmOtZD2+N/oDTWT
B8aLfJcEOXGpLORePlpqUt+3C2EfykcZE/6eBHaikgaMDdn5yo04YvgXv2dO3R07
2uQ5sOgbWPk+M87UejdJ2RI7076Ds3i3YFe8Fb9vCvCD1yY0QFQK0yJv6ifQ+2H8
nLRLqHMqHcW8jb3hwcY3N+4vImCZiAOlIgfL+9o1pI1okLrPfd8pi8/XV+MT4t6C
56ADkMb0IBaz6JCgrcUDgpDYdXHpsuOlWONN40y1t9tcUXLMpi5buFQHz6BL1Coc
IoAxriXYw00leI9TuwDo3NfFVj6oZ12P1ssaiVIzBhU8Vav8cPa3qs8rZrTyRMmn
7xf3KTYDWyqHMtEkPGGlfV/FoIgvIqx3cMd/TR4hvuV1VeG8qGsBsICDUiJT/pLd
D8C7QczE7hyBIMTwFoEtlq2HQPFgcVM1sIp2d0OpIE58RAlCfyV1G65JyCM4jDWH
eS5EGqDx0uPh6y4DGo6zXIUCsDd2MRlGeqW5F2DpA66M5yzprJ6/a7LsjgSx1MkM
AvjjAczkSF9Nn3Kb5y+Xv6/HA7go0//178qK2y2KNRFNPV9KAACNki6Xh8EepXwY
JcsYXljaZYyzD/Qf+D6+cPKDAZuGKs2rBB4yZ74dnK6JZTiGqpsPpNvE/2+AOwbX
shLmzXWvRFe5MjnRlE1uiJrz7ta41UsOiZiYGCf28BQiuHXAnml5qskNaFJDcq7A
kXDITrAkFyCosPSHWHShBPRILf1HHZDtYBFBkjFB83wTimYztGqb73gIpWKZLJo5
zfLU4K5H++H+56fsw4KjQhlYbfHRNOcUL6/D4PgmYSioKsRaB5lt36B/x+j3YoGF
UVfHKfh61B0wrGa8F/x2EAYK9EadzbtfLKsJy+fL+wKqPpC6WmWeMq1mujoQ31JM
OAtiSbNib+59/GHbUpQOpVZ744wSDHc6abomCc1irqer65UT4W4zQMYJttFGl0J1
c9jG7EqQvxkrQt5kGrvPCR0EJrGRgs3W7kfmi6jsuBF0CqVs9wvqOgvRqCmdEi0y
5Feo+h/2cB/6A11Cry9f2mMOB2q4OZnjUVk6DLa14jCGiPQ1mh8VeC1tkFIp5ajd
SPBzqtfJZ05sURlKZA8XCTrKNpCVwzmpfeLr+JynyUEti2A4S8YcSnsK/Lb+uSkT
v7M79OXL6gjV/NTnXzyXGcvr3xlLy4/s4uTOOGPzb++JulmDSUe5yhSI/bODCDkC
07XFquB6tn87cK20EsULMIZycVfPRCQyT7OivcTsrLnEOJcqPXio2QsfQYoSro6S
EsjXkMdQXcBKr8ieMOekvdQP0Df4jGNWpolp5lDWaW5SjTAdzZYtLnRaM9oz5yeo
Du0Ya6vjG6AFvaR9jfOt9l7p4Y8M9Epb7GhOCoHh0vlsYCnhbAzBHGyI3pNLqLzw
qYOXQoC1KS1jN7HeCbB2GDAJ4ayDqhGs9GKtHxxpfzg/9zGfmWx7fo8HFFtA5KT1
ni1nlYzDP05SZ3VgV1zg4ZOq2Sz+MwNiRfsQmYTM7Sm///UR8tvh+GkAjTK1siH/
xiNptHVCOLtakM+0e6R9Jza5CNcoqoJaJvIu0PoP6wmz/jS34XIxcVr/N/nEa7tQ
MjbsqUg4q0nMqffioKs5pflO3XYng8xLGleGqTqhz8mFJ3iTOTudC/YYlpDhhje1
Yh6DVUJY3OdzMQgcpdub/PTpixQymMMsA8UcXVXfptOx0K4nnZmNLWwz7IxRxZcG
4+8iEZFKWJRU1fIxdMuEE4iYocnbADwiCtrnwpesKvQJJukam/pS7uCGfNFbgPJB
hW5wzFyzZ778dCU9Gsw14prMV2pt1iy6P1Z9URG94s1lh/CF9VHlLIkmQlX+t3Xr
eRnZS+Zyk4ruoYJ20ARpDf85NGtYOv2hCWeR6siRMqV/1VpWuHq4c1Vqwp6tvFZH
Mh75Tndnu1v2s0DZEezIIMHmRdzGaqy2QHTTOSvN35Khd7qHsq+pKu2zCgvw2vpD
4iUiS0vMJF/cZ0ZBdUGyDc65TGNwY4j4KFbv/SKHJTX6UzowkYsPQAUnwqI+akCP
C6rhs1LwfNLC1zdZ2qaMT0ZxRjWDrcf1BXP7hCI2wMw/uBsbUYxxeHXyq9vM/zI1
ebwgFe2eYZcl7hS/V17GYjcORwxgO28m4d1QmS/Gy960beqaR5U0H8bCm0O6XU5R
MT7SKRLnqA0mQVxT4HL+dINWHsATnenv9HJodDpZ+PPclgMJyjc8oZt27oWGwVo8
FgYDFbpXqMvGZwCTm4yVfTklTt1ApiAOXiZPKfg4fJsC5ouXFkyXm+odyVcfkBDI
R2fFNfx5DdYZCwmuBkilhrZyg2uqDHw9//nSVLlAEpMiywJ3vwqTHLdPGlGyAchz
3Y6bZXJZh8hebRQj2pSZMXDhOuNN8M7UqCqyQMgWEy0TZE6CLHUmT0LmiTnZCq01
rV4HN8cS9tBCE0o9kCTzN/2bW7ZsXO5JBialNQ4P0a++sgtDPkgYjQ2KvXuXf5FW
M3Z9px/DvrjuiFNpEwc6oHIjF866LDzcCh3uBWcSuKJKDFxtwSIT+uqrOn06cOB9
jISf3oU/edbDROFPlTd5sIhixnpi5EBH0wfUTQ4uKcEIO7Gmgu1i7uzppDiDfxVS
KfTNlqrD1FFeD9VdnHLaEYPFlERGbl0/X2PGOqQpxgRqYNEJTZOB4yw1lHiGGpY7
uDgwB7mGAhnZCV9BU/2svS70RKy8oez/8H05d0g3ykdxzFx/0H9oNSmsCHbnMqDA
DsSqU41Xr6fXQKTvaM4P8CTBT7XoYT0Be3FDYL0fbXTDj3J5SQVkO7cKpDScvNls
gtTZ1WHgr0cPMBEyn1BoTlnJ24Pk2Cg5EXg1tFsPa2mjrZWadITnzp/ywQMjbU3T
MQBkhmRxfyCX4Xqc7mY+8MIQFCi5YrF4ReUTqOD/3WXk3X3dp+mdh2UuZCPNid6S
BVS2RQurOk/D+zhf4I2Nn9Cw3bptOF4RK1vsHAAYPyCmxvAFPqwz3ufteU3/WAFh
2eqrGi3rafaBGxVJRdYcwqrBZQSO6k5K3HZwahpj6qWas9Ib8IdQN+dHqbbHKuDc
M9jKcOOpWaHn/0pBVPC1RjyTax/6ajZylgC2RUHJrLdFDj/+4fqNiOZhOeIamxpJ
FsHNswkR0Ex43dUuKE4c9kqnA1lj8XvrdcmHZdPSvWTSkl0UsHLOZOwObKqD821m
ee+qo2m+CgmOpZnaMs4ikHD+uJZa7KSPzP/pXGLCheNqfw0IkIm6lwvxCMajJoBQ
4jCZpgxV5OYIxaNlgB3sMul1G3110Gv/QH/Oh1UU+YeM2mM0JOMdrC63TWmUHLrK
JkBsMGGMMfNh/agsbH/JDcNYGni0/xg+A0/H7HgrKyDFGOla6TWwaKsrm5WHAgYk
/FOzdl3UefAzTkNH7riUAd5+00KVGGnULjjH+8DSUWrSK87Pn81P8sd06e7nP06f
JGFsaB2WkWyxzETrOz3JvXhEmMWSPYCW3XR/3cluiTkpdeQ03XnEdhQxlr9SFGZy
PxcN8Rg1XFLTTZc51/grEUWIkf7al83RGOfNJii2vrioX9NZuYYp0ohK+zG9eJ9b
Ugmg67+A+8uPFkueJW88pSYXyHBNlVN0Gjj/xFcM3ky9mHoDq2B9Pd+Q5sMT4ypK
loTKxUyEqGMymd5viUTF//By86xAmnp97VBYLdlJCxwcO6mfuMe3CHARfOJve9xQ
tpXl/EyT7jKUMFUOnPxlQqHAhUT3pyfyiXHh4l1vwwIdyjwWQ5k9KKECjcuGfqIS
viEX4VucFRp1VA0eaEjb97cfBALRuZC5MPg/Jyq36uzSNIa9gi/IyuMlkM1Stf6T
YD19o9bR6z4l/p36SRBkKnxbZ+Z8HqBUA0BHthovwTh3BV/bn2FPwQ1LslSwDPmN
beS4l2jFI4dbXOUnN9QstnJ3TrUL3EbCb5XkF2phDTnq+j4YTWf+DQ8PL9SJALzT
thpf6iYn8zAyTbjvp1Fdy21NlocRlLTVXA9tFEco/9EV6cYDPhd8chKrcGZbH5q4
UMgeJIFNpmW5++suicjYFhppUWexeRep/e7MSOLP5p02C0Dc1jCdsOCiZ41O/uUY
c8Q7w4WSDZ3dm4ZgY5eYPMaJN0DRmuoRqTYwo8Jw6CbDVYjP48IwEmnIFoLbaUJG
Sraa/PBAqpRhaCIXVWnYUQQt7Ulrzi1soMbnasVL5DHIRnaWVf2uGWEUYjSYOCpi
H7yabO3j28MTmoBJ6iwVIuUg4ZkJ7HCp1EJQm4VYBoFKMPE2sbmTFsv+dh94DyIT
5hM8Pp99cqKD+zNF3DPkHw1RwaFfrJhorSRQzfPDw6/3qM2XKruID38BmMWn5Oky
A4oN78plO6LRZW0sEO8dTNC2KXGcYGY4UdXWxMILyBBmxbuOsgwvBbHOC++nhBkt
V8X1vJOYyfzMYK2Soi0xKs+qEjxt6yciVTubF1281CBmRMdrDbSB8qYFsCt6+wB7
WXY4Btnfkh4TuSZa7lDPONoJYPC+xn4y0hD5/21jxTawPvvfzhHW+k7i0jjO6z3S
0SJDi391YAocudNrbFnlOCUOHpL0UZKn1ZgdyVidiZNfv69Dm6gnGTw3o37jxX9L
ODyeqwFEN/EsqJEYM/QxjgV/U4KYv73xK53Itb9J1HNfb0UikUUpv+c9gCVP11dp
yHSDoW7aujlBOTvhB731mbpZKWctwxETpk87h9B/QjktZcr8LuV9H56+m9DoENE1
ws9eYYdaJCqt42SyRgd8cuZcFuijYqCiolN4jlR1Se0ZZCWC4zsk4vVq9IvKxFlC
TXVfC8WQzaFYYSdbnIwVJUhER9EIlexEigE2F0T3ukMJ3k5Ev8FIp3IlKUHjBrbU
SfLUE9ZdkV0W9Wd+Y6/+eIZgZgQBRZXdr4GDSHJVmUN6sBUwwJve3Cse1WwJt9o+
7as+JdhkkRLa6UPFsc5XdlKB9EkzssglpmI4QWJue2qgQs3ToJwctBy7qeomMonv
E9sirL+ORNOVUaFBLXMVusBP7wLPAcJIDqtTXf0zhkeA6IiPCF3XYOzzxV+NiaEC
MaZvUHqF0p6yzx4BjQyHad/e0mWMiHxoa2Nq98/kWVb6BAxmryZ5kH+ZerMwYW3r
yKVF+C9gVurOMD/0boXivnm3O9iGdfjV65BEEgGGStqk0ijbUR0A2hf1nWlDdRia
O8f16vGaMSx0HhGnozJTdeKOz0heMqLLFWTojtz9GsRFKzBxQ9pgcuBdRQP14A8i
mKqcnWdczZZlFPX6LC4i4FxOefrF5+wQw3cxb292X6himjYuDgZ0lQ0DIe5hcZEg
Dyj0s0OqSt88xwFNJYuADaahQZCgrLLMTZicAG6IwZl2euckExn9rVyFxjXc3pCU
JVe0eoKWqmLhIkk8peRr50uBBZC1hyhJYNeZWVCWi0Yhqu7rLl99EoMTLJQnFqv6
3HJVlPnR0WzR6u75VL7AJYaciDBWMcOBg5DZfPn48MvcMqPaHp8Tm8WBjN4bcTju
F4qlnDtDBHdElTnEMVARtx8egZa3HQCe1/NLil/GvEWvZL7rpG9iNdCkyP/77zrs
MoAXlicshsCxSCFIU1vBouKnUaiAWjFfr9SuvA3pOSzEgJdECXE0O4+d/4KSzet/
GcZh453HGWHszxT089n1WHtIb+JQyGnMoviDxb70apHVJOOmbGIPgddXTUMjkXJO
cKGlGwcqeJOh93vGVr7hChZpC3eHGdNdFwDtocg8WfHoS7/nkvwtsuCTgOu0iTho
YlGgEBmkLP2IlI7qZ7VKNfpU3D5Hsb8MO7VeDWBSdtUfqS3+JLHVJhFrxbuR/enZ
AC1ebLQ8ONoaovVfnzOe6vlySvOudC6Je8bhVjxsgMCaDKobDn+lHPG8VVywpurg
x5p2zHvoZxnX+howCppLdI15y4EXsQBVFFsdR7bZd/eWUOcuKjt2W5n/YXFhohSj
vUY71/TEhGHM8PErk9XgcLAO2Xpj5h6L5BM2G8K58YoOjtT/cOcTabl0tFAfvCKE
6Ml2BcyFfAC+BPHYvOha/QY0mUyF6HTt4L9bbXGL651Q2Y+0+G2IvKQ4XPfuj7X9
5IcPPa1XvW1+FohMjY83kGVmccZOnfRIjYfO03ZpXEh82gJ+acSQZb8kfWlxYoNO
kw3ksk7kGnEnRVh6t14nDlFw99o607YuBj/jSjcyYbo44qblbHR4w0uUcGYJuhYh
ENB6rZYam9+RaGH5zCtFPPfhvHrX/dxEmghpH8+8g82uOm6oJIZXpsBRSukkwJCd
cTl6+xw2Tioats655pG+USgXll8RQwcnqy2zwdBykuQqCKaBpbEG5ElIsD7MHCzZ
6wBcUA8GaXP2A5LW6d0rYv2KOLgextcTF+xd0nmWitxt/0kXxbNOHwBPxIwkYRZ9
kyBXsB0CX/zWPNiZlU+TfrArjGCK9MuvVJH+aZFgMvjwTKeHdI+erYCDNM6tp6rm
6RvjTfbZ+m+5uVx4cCsNUZ6mkezlGWv56gBbOSASRkelvDe6wyBcAaLn06ykUFI9
SSJIzhmkO6+e6QjUPODw5mC6EsluJd+aZmN/10V8d7XuYCmA2anHRXHhBYs0YJwb
Xb5GNSGf3YIMV2eBVKVAYWOJ4huO0BTsqNFw51mXKl8+2PAB3zHTpRe/sC3g64HQ
pIlSPG/2u99bPTVO4QeOC9cPsMYytD5neaAL41f6FqEw168fmY41OzYl6PM0/oxq
DW/yc0yjtnAZ3uDfUkxP10NNzFzIFpL6210fDz/Dn+7At5VWQ7a26SwAHSYUWYWg
QXX14YIalUxoaQyGO0IKa76uRT75woUR3RO1lM5SHUE7OXYvKI3JhZrzNwqw5E4H
n6Atrzajkwc0SVoTRxU2k8oesegxGiv1k14aFPFqaDHHJ6nOQh8fi/rgp/RmbnhW
nZV+fyLcsf72aP+/Jw0X9UKYTni5GN31PkFFJMvRW1do06co9+POHLXAxN1TYfFa
homui3C7bLnzS8/67x8iXra5eLnksGAT8ljxg0qxMLebYnvZAiD+B+eM4nCdtizi
aqKtW7N2M2ctVZJZ05YYVaOCrLH4scrDgfyFxI6nErOl/G+ubLnZbGlD8ooL75PQ
wBhg1xKf35/XHgGbhxjsDXePYIJ9Woe5k+/YGfSX/SntvNwiZW1jOCk3wNbY8aNM
t4ARt+T91bX5KLb5rqIpgKkj6qoYaDm888as0+XlZeI3D9+PcIPrDSCz9EWtWqhE
BBypZ6zF5kF3mZys8afgCORNK4T7gFoTVLke120HrpPcVeV8d1T5lL6xL5YHoQRe
woyY1mv+UlYkGNtr8ZA0fECwhHlGl8RMqrHsIuNmzIM544VL4TdFKc4yJ1p/yIiU
UedL5HBht/Quf42W8Cgzdn0ry2s5sZE+yQDLkjVvMIoteCyTRYspO+ERjSEkIypA
p78rBN/pBeSN/2zXcyqBMiVZNgxhy4PIP6i+8fmqfdqhItxTtPqLenrf9a7Nc83/
kiOHokzgb9988FarO8tMno7OiGWC2LeSk+8YZZIDLqqYbNiIUWk4Z/iCyf18FwWy
5Cx/bYRKyKCybQMQO1qk3UQy/Yiu3pfMx4dWk7KdsLVNCEkNJdT3Cc4wyfYSBNfO
bdoK0if3iS54f0qNwhq2M/patYUjRJPAwzrnGY7IuD9M9ovTxg9qIeqKvTaxssdF
MJa1WxVQBE74o6Cy7VvwPO6cJF76DwAU07FXKiyBn2sOtyGi1H4Cm/hocDY15fTs
F9s9focUtFmTbnhKCcasdJ2MzKs7ygkuRHoSOp1erGdZbr2eK6c0lQndPiEZzlBv
dVVQr5SHvQcEBTKByG+n2ts+SUG/CROLgLndodkwI4ljzNO0kXcwXUzLN/Lx61RG
HiaT6B2CCqgqOJSo3YblA4ugpRjYVyPOhwQMAYLo2P3TDTSLNoCmQwUSTTIkL8di
OI9IyIOUogSGjIig+SRzytr4PVQyQbmjz3pTMEI+H+6wZfamU4vwGyftboHlvkgS
QbvH9CgsU9+7paSvgetQ20FTT79YpmAnP4gFgY1xoDMgoRpMaSEbdf6Q3V5EtDwz
Fg5aUlSU14aOpyHxnEFpEO1lJgA3PViGGCOcebaBC9K81ho4tnZSFPPs9ztWdwBK
tvD7w77RiOSHcOgsp8y68IomIFi1vhImr7AOIlHGTwEvjrVK/EL+qAmQS+9vHqyz
vAQ/s/cY2cAgzTX8SNSYVp1XneixgKhmYbtsgLqvVySVP1DQvPj1gvZAZqjuCRPR
QJB/UFkQT7AQs3Sa+iG8SF4sV9P/Hx8MJFj4lVLuPvCQlQrX0HirNGuNULCAtxta
5fOPxts8TtI3cqHSZLM+2UahcKt0xHM+CBJvqMJ94YctRwmNCNpsYDC6rY7k8Zyp
WIkhiFaxoM9SJybWdye1DmcnOOpKF1xVMjObR0PBXGRuPzRYLeH1mkQInKz+jfbx
uYRF6Dy1z/sLzYC1L+/k4koyI/ioZN3BgvSp3Ls2X08bfixVUlMIKblmxqGIUW3S
P42Ew2ijr27TyT8wPWxRs2uXFk8xXlfSuEGJhGBCQZAxHlp9blAt5TAzClyRaEWb
l9ZzR/SA2Ry+Csk1lfMKqrHm4aYGTQa72wc79550VqCiqNX+fi0Od7jUTF0Z2IV0
KOKD3NlQ4rVNE9IryE9Ho084gSWDiWldgfeMlXE4DtToc5utvu5gfKOfLIBhXoi9
UP5xiz2zYnzWK9lsFQCFQr7RrJcUv2GwH2pIwSoYXasKvOD1ERV00FguNaAZuRlg
4uK65yuhlG/u8s4zLK2srcdcBbFYVc7R17c5LexCI1hSewge7rJKDRVqBq+5TsUf
1JwiHftutozT6hRaT41bYRGQohb/ma/W1UVGSMYWngdW/54XOWMCpQoW3FSzYOFc
7yDiNPePYu31TRqWTRFIJo2u0uKEffWEpDS2UCFUQMBU6ErtwSTaV7AKucBmZWBk
yqih1qSYyPlOap1tdr3uTUwMZLA1FVbrmRKcKxYNY/Yk4NMmYhpqu913PspEk34b
ld42TzyGpp5Q4kMlaEU3mqqfmlTQpmiDP/olOuuylCxwb5gK5YHMGI1k5dmWcUZe
RU7DVRrjaDf4QXgA7PViibWXPdHNwOV3/Rv7J62lF7C9HdSBd4gdD/SP6sqjPLL8
V4Cmwxc/D3+BqDo7UU7az7AWMkbOUFdB3nFBnWpPCJubMR/6qL0V4NDEQzYLbXWZ
ctUeX2LQfHO0sCTHlA7YYvPvoUumNBMUxPfoi5CNIy2hPkhkjAllBmwN5aGptP4P
6hcnsbhh53phb1ZCmd0rRDnTej02+8AHd1HlldnTWkCH649l6TLlvnGFKziMESdU
RTBUZz9QQfXekms1XC0xSSLKC1a1871yT6B88wxZ9FEfeSr5YfUDAUWQEeupDhM8
41xjQQqRuzTfulfWpgi8ga0gxR0di0ylfUbGA7CerXtaeb3o96R1Ran3LH+CqDtR
+QgrjtcHEFKPRIxk/x3HWTy/pv2XVJ136dEMSFJaY2XZDeLD7tWdBfJx6RYxDxSG
nGZRuQFoygC3LQDcx0hfc9NbnV3QIpn03VNh4LN55LK4xUsecli5RgXKzBpiQP19
BfLgWi3Gxsem/r0ItLO/eZfsQHUmZ27fXRVzvNFwtRQBRhJq1XTqc0E/Eu/n273V
zsxWDtQa4u+m/4gz967eBMKFgmTQm8kA903ix6TJEhiZgWZZFRyPCK1xbq1Ebldg
U0T5AY6MqhMSZQeoW+DuRvnGZzXn3S72PIXYdJu9MTi0Aliv0CA9j5N4cJ35SBMw
Y8PBQRvOUI/aEIASoxTwTphz1hV42WnXgmEqfaZ3uszX6NoP5AF5IUeyC7FaCzHy
ii59J0Y/Mo+iBLTgMuvFgtYcBYv+iYfiXek5cVjRUzup5khL89DCMxRJ5GnTBuT7
cB8tHPreA487Zv3QkZ+TtSUBG1NesivIQcLPYZ+XhFKG9Mzarsv/lP+s+0aIfZ9E
rhsjdLWDuhnExkjkOkg9iaYmxwe45lVs4bZiuODwnSxeb4losHJ8/l45yqicJaRw
+tqSZGFuUH9bhX7nvoFEJWVuOeb2fE/h5tpbQCdNimXn/KOxPQblh/mK2mA9+c9x
euvaWPc+CWU0h4SpbunM2DVFEX/QTrsqoTwAuGT3Dbttn1BDnRVzZzRkyJNwUZWT
6e/uw7FPmHagJjhVcYEx+7Q6Ei5ErHECfHnTfkG68cWKHyDOBwaxaZ55ZboMzjxG
Z3aRMIUB1pEM0H6YoeTUbAfqjm3waSNWy4IB81a6ei/h/iFdNf9gb0HnoAXTdOWe
W+OeiBDBvkMEo6CpT8ojwqUCn1jH/C1bIV84V43EZgYlJRl95LCM1uMEQwbTcrhK
7vW81y2EfUlyAb/Xj4TU3qV5qaf6qKY/KRlY0l3YXFW4iRjlFTw623S3dsEo44L/
lKJEmEtKxn/IJeOeA+37tMo9hrwc6rBVQ3QlwrFtFw3JqdRi5tr08eTgwuaPKZBD
A7dGGsHJlKM8XP+eMmDggMOmxTnWKNHJf1QymskmdiiG7zWzZrWvrGZzOthBvbgU
1RzNUwy88NAMs+CiN9sHa/DDU5KmTP7s4g4rgUpL+oCvdpG17hhgWY4si/Pum/Ss
3iS8VOtKpjOFWGMhFrQ7yoniEeb2ZZyG6fbULouOG2UbBsm9/dciK7wfS4jxFDqE
bRHve+yhdE+N25IPKcln6sKFYKWtl//dqxNXkScvV1279ru3UO6jDJcXWitbWBCS
LytQ6tDU/zCDIvgNAJud5scUB8LSNhw6fi+IrJTlWekMhSqx9EWVVXZSOj+wCERw
EWbjGDewDgpnUtIlOqZg+C1ydfbXUJ7pvGZZsJAIDtQbbtR4Cspp6gmD6qTpN+1r
NEW4yWfXsqzrVbRR/GvRSCt0lo08KkZxxb7l1gRwbvEowzWpUfqlRvCAyQXpyR6B
Q/HGJ2BR8t6at5y2V9ic/wxXoXLrHfqbF6zROHfZIK7bsodID7+fR4326ZlkAn7q
2wrLj1DAUSvd1ZDJMx4f/B0GJz751P3gSocWNrjLPjts1JvKvYG/vCM6L2Sww8pn
jUlkJKaFedZhZcG80EtMiMWVq91BAbL27IMyW4Dg8EYSsGqoLFiStX0p800vEfvI
BuniHeIDuEcNhFZEkKz5k+7wjErU6DS60zmlvIJhKJ20CCYVswuOYpKtMhRvv/nU
CBX+vWwWtR9iog8k/VBc4w88jFzYDTgB2RaFHW3OcOvMYMAr4jkBGpWsWoqum6DB
w3kPAotRK4RiYy/CBFOSXQBBrjlic/GKuMCxoN1ARlq7080DErj2LXre+YlXWGlV
cNzSa5zkZAqUqJCJAaQGX4+Bla91+SsTB+mmOLqKZAlBp0Ok5LkKZILUOe+c0pYq
kLWIlapmbPFHOQfNDf1p3a+nxKAYc0SGXRKgh7dXrJe8eoo0CDM8BWgXcZOYq8Kv
XiJLw8LQQvWHmyzPpsSxKP6apIxt1bwQnHfrkW4piLz/ruzTbnr4vo5q8qdMcOwr
NLRCk8dczKx3qFJ8nY/8y6TBrY1GYkNKv44yuLKJWiRrkub8XCDKl85ZQDCEMUaZ
XuOwQsS4maTrgmxIuPBodPdV088tUoBfw6fxjX4xa/n6tMz/0DU2ukFG8EkhMLd+
aH7roUYG7punlA7gonrnAcTP3epK+pZN4hGsxNmJ5YGlIp6SpcM+vhr/akHgihmN
DWu7DEyTwg9mYVhmsm9/iNRk68dduc5jPjz4P3NxjohXcZ39rRQhHeZkOjCifbH3
CLLVmhHQoRFg49Ybyh57uaxWVmzl1FB6pX4WAScWtkfMcS3dwltxW/3Vss22pWBk
dDVLf4hZ7+No8CLaYit9lTmeeDNH+uJu5Xm7zy4gP2UopWgE6F2ZfwWs+ZyxUJn4
ciH5lCnExJwTcFB0h+XGz4iuchtHMXuJnjQG+z6zjMXBNhUjWvBA11y60BSQ6JlS
2qOJun+siexqnqYgqEE1wvXArBnpmvTQJycWLraYsYbXnVFoPXSzfXBV5XW1+z2n
/KFTrrY+bDzBJQfuXFfC7s2ShOsz8A3+xNYc0Q9NJflNB1YvF8Kl7GJALjfy4Iyo
FMHDfkhbnK56/5mReCV03Ovm3y2p+lRGYjZYYVvB6LNI5M3Knze2SmojUKtsQoxV
VQWkCVqevdCkto/BzmGRpWPDzzOsxHh9zogksP5T6ePvwve68Z+cPpJ+++apD9kM
JRzeq1WcQSibi43muZvKKa+BUtbVlyqfQxeobspPQJwO8ixRs5R36ibp/6BHqTMg
4Vuoc+jovc4bxKZCMTOAeq0L8JWYnKz0FKcldXnh83vPzzeU5HgOx0j8Q7vpcyFk
bjYrKKR33PxBfVl663XkmtCV0RaIb0YgSF028Jv5W9kK9Xq8/G8Lpk9bilZP7EoE
1CGWwoIoOK/M0/+YJLVQEd/r0qc57/h7zkh65YKYyoHmyJNV2YJreNjtDe/ueDs2
ElXj8Zrv6mszvuYYwbPVierAWV78WfYveLCPcRP+WggcT4AVewn7BSGttjJu3sxj
uNwkvPMK50JJHHmuWTAKsj5Lnvnguv2jjjCqecWehFwM4Po45RvDHl014ivKZS80
H/zBWjNmZzDDzZV5GVJ9G6bbVJk4ABGMunYvzu0WwMrqYaWKvhfbGrjVOCH8LutQ
h94LErqnxWSP/GQ5aRTpkQZ6pqYiiTsxhHRUWOb4UYfrcs5XkLZEcIhaX948Uc5p
Lm+gx69Ua7F1hHrH0+TJzOoi4f32vl/SzTsMa+Sig4lPmiIEnnE9MtDySXOTFBrI
QzI0IZCM7d8Og1wwe5G6SsUPqIIpUxuasc2xeyoASD2nMjMPUei0q1I1vmGF+AKW
oze63jLyqZ7VUf/MVgaAxI/+bWADWzVJ1C6L1w+Ys2rWKhRTlK3/dHAJBI4fepN/
NxJ5SRF9PWfxtLw81GkqKaIUuxXOBk0ckZXCp2r5Xs7lK4sIquM8IYr673KYWp52
5JkcG6g61/1Fsm2s/UQmf0r0+kki/QbqczibpwTLtKPzsFWBhgcKLGqRry/IkloI
JAkkNJ9y/uoytytOVUmH9WDl549Vwz/sP500R7IYp+zHYrwRGXKBzp+XmCleJ0ln
d0VpS7uyQu2VhQXABxeKrT63czVBaB9lLsVhAXKvxXI1SmnSahiZvYR0/cB9HA3j
XH8K3y2HwF54kzhAcKypzOrGu/KNQST50EivBFqXvQl32AKymjTqnJvKEo14RuXo
L5zYB9qEmocA2AmwIfPy++OyYuGpgKTBmcYrZMvWR7jriu2Sq+mb+Mj1IAeRoBVq
aMHC4WJluB2HveoX5SKD65+O6oxwYTwqwsAndusKo8rwDUIssQEahZSpjNUVdYiW
RaNw536Lm5qb71w7vTmkKoHqiJC3STgXznFZhv2IOa3C9ccPjC0XaXo/X3rdHR2k
7C8AI6nI0jPfShkwzZ3H5goZNESVuIrrMJiXTFWj9jCR/iCwX1tjMNwWJPhuvmz4
NNk6DTiMW6EsOFmMoSAniixhHU00z38UW3gkhmtqQMIVfHtK65Z9fer/vzAY8fah
kf6Xh6C94ba2DopoqEtsYXd+XcrZDxoYv+dC6DOo3/HALVzyd0RcCvLO4XDtjR9s
kxQwl1jVxAkiBvZXxUNGg3JHjfnh18vxAkBita7ng2Bit5p5N111Ul4OpZ5Ie7oJ
/iGCfpjpShXvGLfdnbBNNk4V5SBKaIBfQuF5zxyS++s0jhdDUUHz9zDnlZ2UxT/I
Yu9njt6WvM+r9+8NE+AkrtkGWdH10Vb0QSwI6hWSftxUi8V6zbIbHIrfoL8JRt1I
GGNwEzJG/QsPKnRAEtTfCgll/vMGWXfWdN1JI3Ck/bjMoQTtOvMmNQyw51a4im99
Fqdra7xMpzUkbEuiY5IxJ6SZGLmffzimcik0AEl4oKsBM0nvirt626IVsG/KJee6
m7Q5uB/hBVA+Ho6qe0ziZ8CPQqCFAiRZSiUXWZogrD87iQmerpHE86ND09HfK8yy
LMYi5k6BANHPgKhLxQ1pgS+08WXiaxrkFJKlqnKjFn+BrR0SKK5t7eOmVTJY1fji
4Hq3kEiil0auDS9tj5m8beraMI+c5ooJ3pE8saA7JTdFidjK54q1Jr6VslY6KTon
d1202EM6bYZroFnKVEy8SfEPQc+Fq+84BCbNwmoMkxfri3QqIg1rBtyA9DSYvvca
b12JnDGVyfLV2ORFlEcmwi++GfJY/M6ckRW6EsnZmXi1E7Is+8TohymV+12qeYiA
tk1L6pAa4ymCkxVDJebKHblhfqlexPqp3+obcV48iGE306O48MfwUOOT7MUGZqui
q43wKj9BF6nnYdSNSBxnPqtaATz8IwdfXWalRojl1evoxSdHdTZtrMBPR2K84D3V
s1Z0q+F0IltSqBKjtleV6+FsTHP2LHEBoNgoRDib/iMWZ1xmbfZGBxgnIw2CPyVH
O3ZqoQWbgExJdXZtGouWR8WKA+naq7mp9v/+7AJhtdAElql+BHxBiR+JvSG2ydyj
0NxTCN787OY4yf2lUobX34jzn5OxT/kdyPnb+n23KL88rrm23IYATH+LpjIhGcU7
FlcH4fZD4e9A/W+O5/yaM1vyVPDKztyGZOnzGVyPmVpjTdAFh3URw74gImK55p7l
LR3TIa+dACWxNbpTyGa6EFEnd8kD/vRoPC+XSRBb/MH4UhraKwLnTFnM+Q8Cb0jv
L68eHDTm0mfPEn5A33v1QpVMBmtilNqSLVBAMwwUd3hp4ND/RML3QBH8MMmsTqFc
8YnSxiFa51MSewhM8YSlry2PgBSW9mkuOd/5xN8hTEmjCCLzz0rhqS0pB9msJxc/
b4aMftYVWuoM3DZmoZ2aBQ/7yzuamzhHUCR4eCQT2BYMGkrF2UxQ9GDLdwuBLnkl
cDfTv8SrDlx91SPWtx1aHoWD8D1g3m1oIOpu8nFHfu/1nhNKbl58IRbjez/Bt4e/
6vS/6n077u2ttubUDHABDA59lhLCkhoFu223qhLL1Yk3WX4wA9kWg709ggxv8qQt
5AfuFXR68yrdNPYHbFDOyVQOmAiwYTCFEH/65l0nPhkJBtJpj7IhhrJxMQEj0Pf7
dYHQFEtOTajkGnJJkG95k4HNlNsqAHDAfUrO4iUd2oxyo2AjewWFzSQGBYQjFVNy
+jiyzeVkstn1kqtVNRJ5nF5G+rKMWBy9AUU6cfjDXIXYC/Hm6jHmgGweXkkTCUJ1
Djb9M35iDYzr49AKul2TVAQAWrmbbsH+swQaaMIlkXegSXICEHZygFrQYZ5SWsL3
MBBy6J/2j8LXRlPTVEtcbwB0RgtceVr4RdFlMo7b7kCZBWW60pzMnDEWV697rxOM
c+iGCbGE90Tg8jKM7q70ZF8Mxc8n2xtaL8WOEf212UmIFQHZE9XHM5OpNsG1wIAV
OXuo3qhvGzGmi9aGL85zCZNYkSLQR61wcxoHgxHo72Zxox1n+ZXKNXgDr/QAHCo+
Pio/+6Bk3I6/Ry7wpNsIQ+hYBwxnczc/2lkMnKSDY9NUAI7nCDYMiGjlEoEBr0hg
JI8csQXjdHK01pnu+64oeYDEqbeAtiLd3reiPPkzAOIsOJ/7fNcqucxGhFk1BC+8
2RJLjlQxRqXR5A0So7u4XE6Td9sO+FVpd+omrewlfQZcBIxDx9BAI3tYtzNKGY9X
SYgCOkOPaD5vMYWowFimwlPjApQ8R1x1FeNMcLkp9miAvfrKxWdGqeRrU1KXIpT0
Y7GaWGjQ+rpmqQvTelbOeweyxmv6SBFtCRYZ/NB2r+Po2g9USVgEoKQI10ai0WQj
HpdEVfk2Wa/Gzwkpb8fNRFGEBgae/CoB2sFlQCd2bsaUhjWt2TnOomF4N0WtTt3a
GGf6GySXjVOcVxLRaIvLI5u61SI2rGg3gP09MZ+LITzzD85/G2/Gm9497X9QXMwg
7KJs17t3nRw5iviAA2Hvpxl808JEr31Dm6SU9MY2bR/5R4/TRBEnh1FKh9qMHSYV
Sm2+w2LmKvwCQr4pwh7vh/rke12oV3cEU4YvAXNsuSRBO4sJoURf/LuebYDp+fUM
R6kXMaENpnuitc9dXiJqKvnL228sX87WJNQcD8Q1oiH9CLPBabSm6qA5j4LXBFE3
tr0rb2ObLxBEokZb1YLt8RS6g3fzJo+ojGMvnRvU9lWZ2EnVC15ssP6qzTDbACje
xmQvzXVuvLvPlLE15hWKix3Qu2V/UtXSo65KMVyQta9k+rMmn/AkuLnpN3tuK6ci
Zj4GnZaGyfGPMWB44UBgIfXYrqRbGlbyRDLRr/QcwMQe5Kk5ZCOgCjFpee7KJXA4
OZWCdeMy9Dv4lwIea9PACC8eKWmVSpu8kcBkTOjm4/jyYG2mIo5uq1mbpxrElgoP
sXlPVveaesyyp0CZknN+xbwSNHpUB4GkYwhL7ljG5xzcoCvEC8A34hlJ5i7kW6rI
B9MRQEEgzr7EYZXR+aqCnarFsqHuJUH7VrRjCP/JkNlcXSNLhAkXLLyTKtqJa/tW
atjafTgUaRH7fXORNDaJ25dvcjCkVjKlyYsSmzOluXyjh6G9nGIx4iGGmt4wUCCu
lbMnqarugg+l1xrrKSVsmIA5U0HkWkAxNvltr+jJNjaRrpkMzN83zUEilVNgJiGF
JtoAdWC+aHHB8CmOpxbDRXGTSdOmw30hdtiFacFLU8sP4X96HxY8xS/R/ByrYmlo
jpvEiarY9Cd6z0WnPxSfz0akE3t5Kqt/9r5RE1NZnKJzG0tVS423QklMgMUQjY0r
HoGuTus0sxPR8I79hQiWHQNbgUwp6D6ZeRYr0bLy1saAYwK5TZ9F2L3p5yu0Xez3
2N3mJgTsTzvsffihYAzXXAdCYZkGbqUoorOkeCzyvb57n8o6Wui1CFFO9oSTVvf0
II3AbDSvVecQfgG1m2vDnHR9ZRsUpoNm7RStA0EwZP/qlUUyVBNDSPUfck9/hU7T
UW4Uv9EmZ8y+PztRcjhj2fYhxiPytCESEnOxXNkCvctJdZmxdB2KVWOz4WgT1v2v
R60ez+jTe+uSISNTNCLT0cfVhK74CWUiq8PQ8xk8YVQmGdb7shtFu2xkuqDZ5TfU
Vh5nVbSI5jqdtwppoQpa/hx0ac81UkqcXULbXZSBKRNaeF31qntEM9GLTlm/uND3
Vp2wjAHB5E4GpyQbfUhvOpW86slJeLCHtR4nk6OAMEJAxk/dtgnFleGx7hNk/u5p
zUbDhQIeMxJq4Iez++Z7+I881pOsfRpU6MvRJQpyda2yDEdX0BNriUFnD3jH40Ox
xAD3mPD7bBwx+YCpaReCG7MXQ9HxWE0pjekTHOBif2aWzSHlr2iNiTvn1Q07edfP
bzoX2cwUb2wmgE5yw3nUeqiHzsNXbgNu6VHGhLoqYIgfcRM6UvbhUFAE1DGt9oGy
AdbKiZxRHKIvU0BaIoSiKVc4eZ9KIgeWSoOinzS5E6oeswTaeO5uEpHIJvUopUNy
qE+zV14ylGPGUfq47CScMcZQQtYuE/QWMcwyc2TLgkiRqUe72+Rd61gktcL+EwZ+
vwUdo4jLJKArvAGJUFUCw7GtP5XWs7l0ai/dNBXyKaEsqvlZ4sQpkCLzZ/Q3JcHs
ej5sV2Bef4z80eVqNiHIMy7xuN0cCxyKrUOEyEiVZYBtpU73ShhKm9YdCR9FymBD
HtiYJoVy66+fM16aI2ALTblemF8rmw6lTrEny237E+ot4SJu8xijTaQ+aj3z8uYa
1UBdg9jJP9Oks+zuo82S+b50CPWXis2tsG0ygwNMPg4itu7cBxH+klOshmi2FseV
WRF98AFebWGYp8EGIR5RB4ualIBCHbKd915oMsp1vXPVXDCbUJEIuAW4hNjZt8mx
/drrER5Ojez4FlbV4SVD6HCrOxLIP4sfoJzt+epcKyPhJbjI0a+IBmE8y+rYftbU
ztwXrd6Du8IVTDcKwDDv0v+hk2qRjI7IiArZl0WuXVv6X5q1NH/+T0XxcY1QFCsk
4c2laZWtVko2PzsRHa/tLPtIgLm5QpLhDIR1EwB5X3UAtSFIfTTfSAJ8mZefojSz
oJngsZBHTV82s9tkpwIGlDpkl6yLVgFq9EmePE/lv+IFFfFbhgwOj6zgiloii4rX
wZ5bvAvhkxwtgqzOeV++Rhr2XWsVsVjIEkbUbXKKmCpnOyS/i7iXItfeMtrszOgB
C1vQLcBBDTf6XkNTXrvDNukal8x6m1fWQ88rpcgM71i96kFa7OUzsfIezHWPvj5r
KsyLJx8J7OKkOul5yJURjY2aGNKfRdQzQBAK7+rGgED322spcFCG/qh3j0xS/YYF
Q6ygWWUbwkQRZCSwEtFq5fEnGYk+AYHuT64/BmbzaLDs0AAeYZNGvxYDBvMKK0Lg
Wbtm0xerVaTi3F0CEca7R0H5kOYhuAjyDYA4x75XXhES8UYxGkYTc5v4925tAb6U
3zF+cpesWTXz09Tb1aAgXHhAltiOpVHGfSC8XfvajT5CICgoyiYAPJNjP1CJy3v4
Dz3IScl+Xg5PtkX5nmUynERM++9f2pBIzD5RTCI47GU1+ZRcxu8W3bMmnaq0yDtO
rLayT4GOP1tP1t9uYG1hDfZOazU3A4CFLB0IHGlH6D0z888qsijjyojqbs1U4E6g
ul/n7F7DNFOse/Wz2RBuoagW98noOgGs8zUUigDb429bqRa0v6IxytOlrWtAJjeI
FZfkmbJLoM2fcCNOI9UhAb74gyVT3CVGmJxMnjriHt5no3J2a5ChxhImlUfLqNiH
+F+KGgUgQ+o0f3jCHVl2sYF6sqEVi9SUlWt4FvtgDwBZ641jbHjf/z4CmhjXYTr+
2fOwYxsNg+cTRWb0KV9LlD67KQk70jedSiJlgDnS1ayGSb93uI6ZW1fR8bbGZ7Ko
8jYbbbSVOn4kRPURDL3cE2TS0jeUw6fkn4HzztJB38zjgT9HZ8C4kQudvhoiHniJ
H4bPJjjWAxSQOV2/3Npd5Iv9wPvluJQxT7ivRtzB0AorNfOsnab+J4AHIlVzw89O
6no2yVdwyiul0VbzXDBntTDQfsz+1n2tH4abkGPMEMh0UzpmsIz0mslR2k9RhBlN
vYdWrwMv0XweIWyZRs3SH8Bk4iOXD/LYhvDgQ0yqXLP+D0X4TPD+a6FKg257Nd7b
fl049IORQyOOoV5TZJIUTVEEEzDIYO+xrFhQe2xZWYqqhTIksEVEAHsQC0r5cqA7
WUBaO6nk8usSOhKi3k9zbPl1omY2p3HmX+t6t6YWwvneAQtFE4+bvdJziA5yoruP
BuPe94ZU3rviCwn0VTc9QnQNFze9llXuazh9rr+E5n8CRZ3NiPJ5b8jC0+AbK2ug
tIdjvrbBLZtPJ8gfFV0v3kFf3l1Q7jgZ2UbWuMebscMhL4yiPcgkMrT7I9lQew43
1/k8N0fT1fsa22Fd7k3xVmTXx/LL3IZUcsx3/pNdFizpEJ8dbhl1AM56wjseImur
j448MQAA2/i3WPiG7DsELtF4zZ3vi3E4l+S04ahRBTZF4UfjpMibw4zkv3kRn4sy
z4C+mr+jUAiwlTfnwwHfobI0NMH5SAI0A1G6Ba9z1H61scGab+5N+qevooIVjii8
4veJhMybs18AMGAzQ2WXWLWjLnPtpc717ZhbENRhTR+KBLafk+wnV7GdkI3CLjoJ
F4T1Jhu70N/QwBq5vc+rXCq6NtecljXyopNbxWFXZJjiunebcNVSWEDZdmEMkMZq
0huHaows5U72eP1n2HxKD9ReHXLwi7mrH9Xd7VDoXzK5DBeYguSL4jO/aUe2XWfX
loJb5nsUqZ6I3kxRDIFC0HSwRRE9X7KT2on+7AhDNR6qd7DsVXU1Pr2Xp4tYGpaP
Aoo1f633sTXzrHPlVTLtWZasp/qXHFH42guNcGBs2dRqJX65AyE7XyNnBYcOtu8b
y1VMAZdWByyNlY/lSPyrQ27svIKYbkHuc3lwvcIwVkn5hjj8pV8PWZqlvuq8T6tG
yF9qIhlik1FKLOsyha9OH3jhXIlmlCg9RSr0FWM3aZqnKK2lUyVqUjAhhKWxOPoJ
X30NrD7OwOCCz4I4KR0b2xOjxJkDUypKHAIAwm+HWeZsfTLyj6/L6rDZBf6R9uWJ
q0z1zaHtqWAW9P5nw/DRWhEOFaLG42VKInq2X5i40tafreWd1C5KJXLPmFvBOkPf
sY07Y7vOL+ZsPTETXxsJ+OTaWpWlYj3+35hpvBiMUZzp09F7WrNPR29qO7KHgMoj
XE8Me+wtN9qjkeIx/lmVgtwAopD5QTzVWvcfZTpfHRBTaFAKDs1SfolA1shlti78
5WzP+AqqSSxJ//AY9Z1qXCqrKA9A5nXeC1xxUgUTQM1vbOQQxmJPcbF91HvORPU+
0sw3OdrSCPQHfK8ovr4h6HO1y6gtt/BF5pzPskMFkBrk9KsBEwrBTQoqnVAyVh/6
5FiTdOYcmHOa/tYNSrhqiLloAzuJuwKReXligFt/WlIB8Gui6ib3qNw91YvTGURX
Bt7l+bnOwHFP7rQAKsBuupCU+lO8Iqvkpo2aL1SB3b6fa0AbKN/LZgUWLmX119Yz
cEkjEPHe4DQ9S0FJydNokZZBBQmZm06smXckkAA7iAcp5X8G2KvwndzQEPJh1dBE
TedscSFtVGmxxzulGLKCpTLgReOjQuIfK8sc5VY5127YID/3xJzj25Bf7krdbfP0
s4SZQT9TILl1ndfWxOpSwWOx+16JxND369kwkT9dpDL03XF2LSUOIE3yRHvapqLC
NaxEsaXcqGtdDetmyEOFyt1w6UV104aoHYJmXlH604kE3ioYQPguKhv/+cAgGq/O
Ofv7dMT44dEu1GXWKSkWWqymqg/moFaNUGZdEikRD+TiGIY1w5bEEGaMLLCSLc7S
e6x+FG1kgAJvNP6+DvHRX5NppB2mRo+SG8fhHC0BNzD1FzNbwWOiNKoh/zRu4kCe
SBv0Ug822B1/xllVhZ2O4lt+ukfYXF8u7e8dLYukkAQL0s/yEKSNJ2jY9Aty0d2R
FLuyLyMrjJDLD8yFyLEEvd2mvktT3yPgSq5uo9ojHqffe9AQ2Np8ucwPe1GX3vuB
wBTRH5ZDEAp/YVefc3il4mu7xQj4qgxzAP1WGyGG1RpLa5QjMRdhnB/Z5S/2GIqI
TPd1rAEZkVPEAGeQVscJW49LmPUkMSpYbV4cLP682zZNUXzDe8hcLDn0x0UeRwTP
ZI3c8ZU43lZIW1WBCrYP7CDLtBCu7x+vd32UPX/HOBb1yU5GJEwIO2nWtbf0+ZrN
j2tKIz32m87ZD3w3nF8uzc8c4MVHMc0YHoZh6p885VYF3Xe3X9SIhMny5rLQHrYN
+lReyuIG2Z/BZV/8tdPGGrNO1MwINTfBoa4Q/hRMhdpvJ0pScST/XJuk0g8pPIgp
iPG6iQQJdBPtyz5r4eVorreTBm3rjAMoQUZtPjJIE7U+Uv4F1PvBuUUmY5CKuazi
Ty+yXby5ihXmBM3hKjw+GCAFFFwe8P9MtUAOegXifkCFf2oe7s7ac7TQlslnmQxs
dqXwXfBR+8d6Th9ILyyWP3CjKUs+f/pIKzfkKWGTiIzzZD6zMqEFY+v3M1NeJsAf
8sCM+7vGKVD54gTzbYZ3vv6XfKnNRtvyKECxh1WeR3NZ1cFuYOnHz12UVfZfZQPz
t489ossTsf3phGSt0O5U0Maet7MRgGXXwdK86Iz+BDNX9Pc+drwZPfAMahk28y0x
Y4Rux7GxhlwQp2UzvNXL/+oFF1p075GX+zQ6UqXDlSZ/Bj1CCoDynQOJxAhh12f8
LpZv/W8+p8n5JuT56IpXXtOfkNWt3o0/lfaQEwJ57Uc8f9prQqmZeI6XsHE70XXJ
C87/GA1RLkJ76Hph0kpWOFAZNT5IdSgCMjQTrUz6e/9mZbqZATJt91lZxk50S+3z
N1BKjNd6tqMwXxIR8Nm0u/oMBQ9MM2AFzlK1Dd4ry0dHWwa4vOF3DvU903tklos4
0Bqj0VJTI7H9maRDx+mtmfVMaLGrVBJ3hX2g5HSEdi1inekhyI60S6hCyHff+ReY
0gX4kG/EITYtktiWz32qkMMejvyIAa6zcUSle1RpAU6MOgyDuRcKbpkKj8tX6gP4
jCQTLvc62PFyQt3GE0eodPHRJXcQF4SR7DCpBsxxSoZUSUXIWb/S9JBaNCGiwzqn
D30gLM8piy9QTZbZo6eZcckm3hP4bCI+50IaZl46cVNWDNSXZQzvhhw6qXP81mZS
o96ojLEWtW0VHAMDs1h1mRIsSmuoOoDEdXUWEmF5q4kp2ovCJ6WHH9uTsnxMh9Du
vPxeLUark1z1qtf3UfRsceuXpEZbS4scTQnQGQHOTrKA9vGORy54VEX0tYUtd54/
WCYs7lKx5ZEgk0xVRnvHJ08rAPK4ZMcuy96Jp1Y/L3Qi3+F9Dg0xiBzm/vQQGnHp
95mBz4JZkcGbE5yBhAQzL6sw8x10GhLeqijlBEe3+63YIMOKoyBqdvzqt7EOcTn6
K/zZemqMSODmX7I3JwYkp+7NQcmMIDuWTNc3/T+bxy36JH0qB3PTSP3jL7D4cc03
xPO9pJsk6mncBxXjDJbhc99tIWN9e8zlTw0ISl1uDn+z5cFiSzwMw2LJ++GHd5yb
7Icv/9qSwvr473nHkFJSCUdZ9IGLU8FZ9tAGMdpjiJIIydSVBYSpnpLVtZUrvJVf
owXBp99cu5KRn8QFwgRuG0Nt1RD7kuD3bjZ8Rkty/d+OXL6KZxaSejbQUrC1xjm+
4fDIAlDu9KdPBKKLTKAOd/JQqfv8Wpk1xsxZ+gP5sxYGMa+uoHmmNZnBFms6bZTI
8GzlD8UrJFCXVCADS/JqkE/wadFk2iYdir9ZU0dl75T0FDcAHZAqnO4NW6rL2KmE
84yTIUgOMPBDNETBJ9xBJC5ee39dJdTkcH2BIeF+QbSX6nGCArjCvt//AA3T1427
P3ais7Di3Js86RENByQlsCI4EY6rkV2GtJZYVsmC6Pigu6pIDFwNfmoUYxxJjF6a
TVmL+sw6oQLKHlsrQqQ3QuoO9j7pWQWjvzzJai5B9aBdXUMoauId6naTFnX5Imcq
s8S32OnVYDR4wwTu3xjo8uxDXwehzxjCVdf4RyDs9lYfrzj2sYpcyWExOf3nhLcD
RC26vOLgGzclpL5VLFP4tBg072n0aPJUlfE83/2dKdN05SKyJ1r+XpQe+A1fs8rq
E3XQcqaWEDfdt6dmQgfjIcla+kHF4u9fGy/U8PqCQiX448/8VD/8dBeFABZymP71
B+zeWH0INu4GcUuXyQWt18KzIhjJ2iaqBbH9FKMvmt5P4LVPdYIeG4EKoOT/D4gZ
aq7LHEeBGBykGPFU3/jI52OYNGB9XQDoN091yVfS2q2Cpftd3Sf4bakvUMUOyPLd
0+keRwkaU0NSsrxH1UT0Tixe+cx78rgPEgXK5hjb44bT+VLc83i26igIl2SzasjC
22XCq55v9icPYHwIoRrFRMYTR7Nee7vj/LKkqLSfoRl+5hu2H0jEP39fZcalmGVg
3aUUqK0kSS6Jj4M1xAh2xwH5IaBpdpYJUDd28dwk9JSRMfZlNAlZcppFHYdbThk0
xqq8xbpYZ8TjUIP2jRUuEmqoPzjoXyE5iSup1adtnEp9IoIyXkJYYnG24xIQt2io
gB5aUp0TmJr56fRvhUGfHPRMgBOA1L06vBOQQ4dYat+MIAb8LS1avqDL+2mDr6ql
uKRhFdPhwps6yLy25O/iwFtNCcJZ+7A3/bX/Q1scgUGSU6fxkuvXJhm/jS9alhDT
+S/2XqoD3KF1MAd0pmKvPYT3ibbWxu7+TbhPH5ovVbhE+CtIknq1J6Dx/nkAlbAw
WsHPotyasglA6OmGUoX/2yD4QJyGFeXYBVV08kxPPc8mtGca7EtBnu6tPYp78NhV
4onN72pxpoAvn7VgJ2HeVCJ/W0kr3foeqKv3x4s2tTzyskBBgxvy5RkrFRWb/HAd
hBvPYJuy4bPM6k8hScXDNNnysgB5qq325vGzOL+aTuwtHTaRNxavhpNRAE3ZLDDk
UfMUeKpwUgvAr28cUMkddid8dDY1XvhLz5nBbbC1Bli53tL/r9dccHXnpRMi6rEf
KFDpAD1/b8O1k+iVD5skWd/pMMVdM8WNBrxd1A0UaYlU9ePEcfyqKjdLwRx2HPSN
ty8aFVhCyuG/dlBgPuk23QVxnYa+WJ/QLv7aYf7Iru5xjmHVBElA8qRBZuvxjbRa
8cPoEneT7mfbaLVovbIP5ws1mQjn+bUXYS5zqb8/Inp8pCECOmN7CtjMX4TOD1Et
bjag2ynoki/HUcm2DbKRpAqm0fYULrqKEmg57AuR9+yivp/OP6duOSkskWZdP3a1
Qp/cRCGd8AGW0+kpN28fJuR0rZAZ1CCJdG5liwn8WydEahmc9cFcVkP+hL/V+7Aw
PqOJAJ5sbpTI06eRFwHF9KpKz/yRDkmcsVGDTYMBLntOoajv9MSfrCaSKGyzpX6A
7t0ZxktW/kEoOFwnupVv70Z+QNAf5V6oqCv+/CVBA40GLqHWnjthYlKOolVyJa3K
p16JV43xFaC2KwjxeQuVk8HW2tLAflKzIDZ2ZHo+S80jT6cVt2fglPJYLf/zBCgw
3dW7FrVE3p3ClOXh68nwKx0T0U6qpVk68jMczEI9r/ucfhya8MPPUiJN6dZS20+O
0B/krI8QeJxXvN7Fa7gYa2rinu3am8zueCWT3pgW2VdGwCR7d6lrcyLiSj7ZPbu8
B1XT6CVAFCXurBERwRSfTVLXEinliX2hU7Aq1btm77dXpLD4v5ZSMsMaMeAHkT2x
QWkQOHKzS5+pGtVPSzcZfANi61L6M3AwW9qyT+Bgjo4DitAa4XRIVnOsOZrRTtK4
DFT/9NsEJ2ATOO2RAxjFIIzfhEnQ0QpMEFSXFn6LMEEq3o+msaEiyXh6lfeXtxZN
pdUFkgmspA+Cs8YlJoGimtkbhmN7SepsHtsy8aTcqTD0jBydaAunNW0x9kNYdt7J
GhoHIa/DJ7NT2TmdLVd0EnCv+scEH4vR4B8Gs+zBmftmcOnpN4ygnYystrEQdQq1
LBYrR6KsqmgTNtn/ACLjuKZuvgHAD25E7/GjgO9kbXJPpTj4TlOJC5OIgjYkHJGX
iKcWnH25/oIexRA6W8zpWEkM+IXoD9DRhmsDrTPTuAVSyU4UrOar+dMQVrRm/pFG
zLIq7tvauUUWYKptIQjqgSmqJE8sD5VO/hSf2bq/qJmigBfYh5C/dUNPzcBnI5In
la6lBoTUQFxp+lszOgmwiT5JH5DiCaZnFYQ9Gbee2EW4mcxjwjco6L7/L37rxhFE
t4DQBIMQpDlPNK6Jtp4F6mjhdd/kxTDv/6Ds/z1L5x5wlpX1yGkKYHZxMVRJuMMl
ujX0mnsIA0trttR1MZjdOwjiqhzQARG6oDs/oHHy7u2ER1TLfhAzU6PNEZgevPqz
29xThg0ChZ8f+d4CNMeJQQbxQWY3s5hCQwOuqir/l8QjDT44KDzwd1i0zNB5+eHn
t5tpRVfTGvKmJNfj5jjTFDsEambZCSaIokl5UVwzfW+wbz86mYVoNbudcSwNCpES
+gpmWWshRpVuk8tHpcyXYF7fYMxD/7akqzeoIBavmIzrifBFSkWiyWt/D9qUrL7p
oGhA/w/bQxQdC8VOcpMF5T5rFXT9200SwEVpa6yGoM1rdFIgNjm/b1xkreWZvbtv
JZdP+C7LYNguyPTHvSr+jgGkbpZh4/zPsT5vU5pWhBefHrW2Ul6h47BrfFTYhhIZ
FRuwyk41wCPmZeQnvXjVzulxG7mtznqG2noax13h9SglebJbkRypI7wxU+h2Pwm/
yLTU+16huFgtMw8Uy4oFthcZ9d+5Vm/yGy84OmK8eCiO0rhxvgpG3xC+gk/k4maZ
b0vehy4XHNXaWiavCp+xStiKAso4ZrbUJhHwXZpbraSv+or0B5FZLJgL1vdcIPyJ
z8J/UDREYTNO1rF7NK30tzIUGO0BXbMeesJdFk0EPIDWjz0CEpqnhKSo/qTShSlA
1YWfwe2t34lO6QU5l1XRFr2NbsGcLrQVL/eP1JbNlcRGe98ZyQAiWpwQx2PPgZv2
0QplYvfaJUYYvWW30shwFbSh7XAqTJ5dnz19HKJXbksWU8v5eo6O5f/p36LRsK0E
paRfqj0mDSHhnJKnVuCF5tq7ugt5+2LD8JGI5Gg11SE3gQqcwOQyETECGvUk3Te5
fC/HKG83jUYufzp5+BHQJdBHZJ0k57Y3yaSfgpeFOAaFFZRUhH98GRPxc2GL7bmF
TEP71aY5sWBcx1723pzxiNXAW4Be3ZNu70nBwxCnYYhIFGutfhG700e38QiZm5Kf
Mr07YH1r107mxdyWr1HTaj4rDPgQQ0i5uJqXjTD/AcamP0re9NSh6D+LLjJiG945
TSUmKpM58DBRIu+TOhZ1mV9B6Hytk4/8InTO2OaNX92KZqFqgIzfLjGRLL/cyvma
jDm56qj9atL9QG2ORw610a2yBX7Cs7EdY/583vkFun4t1SYJ9MTdWWf7BHW2qPwE
zUPO//IsN0AFsLokg7zuy5rMFKFQaOWlrBy09MsIqBwQB289GZDBbh9T3r/xajlg
QCKE77asyPU4DuF7H4zf491FHEQUxJW2UM84zdiY1g9L9vN0edZEqnoOZJs6870c
dX2ahtBBbSfw6coTgWx8BD2KBUUCJD+ZqOgnSCSSLVtR0npXkUtAeqW38wxGYKSd
SbGz1ymeNVlavxiooJ7AzMPmhrQIpOZYAeK/NuognBXcn+58m2Y9lpIFwzLZp5wT
+g6sk87GaU90KQL+wc2WcigavmXrC96IR6LjUIw5GJdovOFWXV+BWTag0FlUrurH
9uPIEwWc4q4xL+EkR6EqNI5EelwtfJRMGzhGsVTB81MnhjndzDoufWWFqddyjQ2L
TNAATQyiKiIcGndxnxXmokrYSEOqJTi9pwzqZaIVEJ9+1loj8ZBbfudCnBxYnPPy
IrX/aMBWpUpcYuAQ4xI04tBllc0byacGV/wiwPi3k6UCJNmY+ARZk858/1wxiUA/
USk9WttjsrSnyBqmRE14kDGnhphs7tXVbRPtOCs9RNv9esg7BmpGIWvngIjGN2E9
DBRYDu8vF0NPZGFWYCbp+8BGZUe8Hx5wthN+vHvpSJDZND4lF5psLHQX0QlnQ2yW
82f0UK34sBlOa43LBNVl4cn/JDpdumZZYBCM5CijGuDyQOHhWp+tNoo6yW11Hjb1
b5wUGZXS21mdmv+J2Xvb4+ydU78O/s6Ygdrka0T0edyF04OT5yr1YqN0T37QTLy4
mygCUIdKF5298CkyJcr85BltEy/yEX7dLefk5XL7e1Zzz+o6OrKwy9vHLTXTbi8l
kNzRbgXKMhb6olB6ib7IYNFEzYgo5MMllnZ0BYKzltlV3s9U/odMHzziUAzwrNba
hHyLqGKGiF8Y3tX7ikLWcbdkIGgnTV7af7HRcCx+jY2BgRcB9Uoq//vHgXei+pAs
bqd8vLXp+rXEiVo9D1EhV0we95bAg7OCIHBgWvdbfByVptXvSxMRfgggm/7Ll8N8
XAuY30Ufo0gzLvXUwxQOeRnvW0V+BgtAQ+wJkLGs5Iyqzt74pXuu0yvnDjBylUGl
fi0AWTW7BxolYe81Wzp5t2RuGOcwVsuQZoSbqUCONLKYWRLd4Rw7CaGsMxSU1vF7
/Pg49TV52ZEMGCUJR32pLbgTp3eMtfioYo298GHlnrP5LyKTV6MfqLITQjwOoPDx
XEPCUH9d4d7Jl8sBklgRYBW+MrlH1LWhiMNAMIW+8eGcVkwRs8mjcTdQv67rFg8R
ewOizn6cCr7DTf0BHL6VzjTEKBaVbdq8jQZWkh9gASRIWD7sxQarEqhI4a8/Du3t
q+Kr04tcjfNGusJwQklVmi89yy8qrJEAaTAo5hXOXfNbQXltnF8K6ZzQKne0uMJd
dfH1pvJUd13qds5W/DhQUQxVNdUhMcKmHsX6zMvFGpsllZqkfq78hhcvI+zIKfwK
j55E0vJtRbKtj7SpOkd9JM6W3OIOV4eCqZkcxQBViKYPoeBReycfG03BUW+oYaXD
PrZA8sDdL9hROqZQdJiSo4prPHgJj5mmKyX+g9ScBDCHVkvVAr0qLuVWgGmaGvRm
521y2x6KG0+Ak+PSU4p+O3WQfHQFj7tijE3PVBU052GATn58ZHIrqSYHsipZo1Up
rkbeDE60EH1dq7lApTnBoBdUciNmBTmBDZrDyPV++a7ETIxxp1hnhPwfSZCeE7hP
oPWDJldJEQc33DHEVkhywD0UnpeKGUeu80DlloWaf1tw4FS1LZFZsRlSI9jTCK3U
tUxj5w2Xvww+3c4mb/eg3axKFhZroLA8GLC9nngDqWuJQA1X6ImBDpzgN0bOosx8
VgVlV8M7iBV/4djgkh5uY75bc3YUw1Gwf6ZkwDjx0EdYIXnv7IEfLS3hp3mBUf2N
f+EokT067XdjqcFFwyksgIigGIGGug6aDlhvoEOJ/5svjwk4b5B+vWQzx/r62iF8
78AVNe+gVZJdFDpTwe8IhvjvzDH1hNAcdrb957e3Is+A7DEd63akwsXlY3Ctzien
wGSJxVcPNsjD3p+0uCw9UwgLvRtCbBfYZKd0lrb73zCDSKyJ/SBkGOVhk7kFtwRP
uDdt22SNgJjK8A2dh08fu1Iuq7CoRZ99ljNIl/4++irdoBmscYSpph2kV9DYopPI
hAmeEnvZfrGcohTY7mHG0OavtqMJDBxwm0UdkjeU6kHZzBNOvIC7gie1SBhrGtKJ
UIiK7DDAjSI5XB5dugYm8qld0V4t7R8GwJNZHXqKOdGzcVoc4m/svL2Y3EiOoXzX
gvJ/2ien7WXAew9iijL9EqMWe0FgIOYATB5Vn2/zEoyjFS646Q4m0lrsMoa7V75f
jxtd6KLntCMrA3g0Tx825/8g6MCCdH3NbrwaPCcVwQAlI/knYR5r74YmyeewaJfg
z2yEvvcbM6PvPDAtJGCk2RpEDEtgcEeGt0QLBP0QsKeIqprU+Obqygb5qAVS6/r3
lLj15UgjHIaONp2y+e2y0USw5oPZT9TMm1SnDApS7RXrIkgg+dRJAg/eLArHoJIo
tiOgfLXpIpV5/cEovfB6xQMQL7g3qFeg2qTioKWAcYgSvFDjgGMzElF5QmgfM7JY
+FcsP22Zz3Csx60HiX8yfDrgIPhyvzgiBID4lkGs6HUWJ10z3BkpP4bb1WgMo/eA
flV3fedVZxNVhX8zNwTEbUvXs/brG+mOMM5eHM5CzoY5QCaouOlFWxgg4sOuAaR1
l8+Z4fnXMD+QRDH8sxhaGR5BiO1r6avKJQP7r8uH7QXkPy90JVgXrHxBaY3pHPpV
yqNpiebiEX0he4CTfyebja1o6hgzTtxsDW8d3DVGd8h07fMRuAbyZEyw7VU3jpYX
lbHLyw/9V30tluJnjRFeUBTr/a2QM5jqB8kShGLAf1PCyhjl/zMk0WOZUm4Am/cF
D8TgMumS+6aOGTLq/mTQR9jl/DWzUDfC2zT9hbLtYRGhHa2QFSan4bNMdjyLi8GK
5/eJPeU5Zqt29cv4/Iv54PXZxxCsidMs0fUwZoGzCMxBiQCH7l9suG1j1sbdV6+6
PcJLiQW6p77h3s2wiUjZ1+IE6jF3Cbmu91tsT2hr1CMppE0APwBcTI0Jb74vbN6o
J4eQXbpw/IAuGLA1L86fdru3xi2CBq36NC+oxfG/ImQvl7wteAvjuOHBJJVOvoLA
cFdvdftBrRdkn+CV1XR6Lz5LunthJCzMBzTqT7Cd5iEPr0yMHQx6qvcGUOH1ZbUd
XbH08nRASF2ECilnXDekdxIam4k3gPG5lxBiCU+DfXAewPFycxz06Obnw9n9xKQB
aLRjUwz8pm0adqotQY8wb3P4vOjEl7EXMIC6PETPL//F14wLSBY/qgtfOeRcKyrS
KPtiaAPhTQO5yppZ0MWKmB92DoHcNZ55Ab2PTFhiHVViN3h07xKvm/PdxM+Wh7IJ
4NN5xVLtR94PWPsWh/4kLm3MTkNMhEnTegZH8ac5Gikv3URWB3CK59urmhhM5wRC
8HbZ0JeKOHtAz1M+M/dRpZVCnygKN7R7yjCgzXnFFzJ9405jK4f6H9vrNFMeAD6l
DGZ6Xjektc1fYeqolcY2Iktm4xI5ZAYvfuyTEN4vFD45ApUcEy90hI+AOUXtCaUb
Q6cGQZNcuR5if36gQQw2+Lw+YUXdwTQprAxzMVf16pTgbCtlXcpfnAnf4iycJDW2
F/LDPRJkRyC3DEZZT0ky1J+LcOQBdI6qE71b1OTKJC4e71FUmDQou1Wvr5/daXfJ
EzCiN3N1hwbDj3OVXeOavxd3SLEJVapfeFg+2c160uMS6qViPu/3lPg4EJSUagvn
wlI66XKrUnA4rFOTjLDf/Z/OJKXsUBzMncSW6ymy42bdEOPsnR3mVXj0Q24pmTF3
p6TsP5lO0RnWcTny6Cv3CFG6zxWiCOmGl45RhsOdxxdJsUu0MfKfwa5D74KYMYL0
SYDG1X8o/Er5N0TNtcVVRJQlibZ0xCWzzJIRmBfQmurlKQ0TsHiNs4NhvI7tK7HV
CdLQ61cUVcniM8RGcrQ66lRc50w1q7RpPkx5UgzjMWwRW0KvKoixMH1F+Qk8N/ZV
WX3REXiInmX3xYH3gHxYO1p/UM9Cj67sznzRBWE+At4TQaUntsR3yL7EGnQfEp75
+Zif6VciT2uA0oMCJH8wt4gmv2EGb1oua0aYtP5pp3nUOkpD7Izcgjb7mhU/yrwQ
hM1DZfe8K6dje4zmR0tyjLiUuY9j0ZLjZzQVph1HcIU6R3TKlOhfOY/V4ol9+q9D
2WJN8Lf91QrF+MNTZoD8ULR32uke+DAXCa6ARK+jhd1EQwXNWr7bx1ykqEJCSW4y
n9pFMdzJntCi2DVi73dfMOWdqHf8mSEyeVxif7/sOwVBwced8C/F1o8StRMwpkP/
c1CS9+iJvrH1BsEFINAdq/l8nY7DRG7SBNGz+3kolOYShzh2SRWp2qnADz9IwJhN
rdM5dWe7QV/6RrKM1bMdEtDvzh5jXWnQgCISqcNUi3BaVkoMTJQzQxBXONKkUlYD
Z2MhdYqwzAdvj/n+CvUZ+pKVBjcbhWYd076PAKG81EwBzyGKxuhOv7d9t/X558IV
Bt5J3uz2M2G4Iw2x/YyaujU4kUSt++ogDoQfDxUUtiZZ/z8QF73V18/OGo62Xmnz
ejzIHKw5D1QExTeyrljEXsGSiJ3sbjMEE9eF3nMlkPG/2QcDxnrZrhdb7wt0bL0S
dhWdQZkBPhbUp2qeOS9e6LuSyc6IP8eEIsTbORzjRf0QqfEEtW4e5YqMrTiaek1K
B5p6wwmaJiIjwltKb9ZWGYI8hanx7eT8VZ01w5BNGJcjxjUiPq2BqZWxcFzUGQaT
tmMq0sQIHOsMzjPt06t88t99bow/7h1OllZIo7zGYXPJptEFiroTLnIS4CvoCzCp
2Wrd6rCsDbSvOGCmVPQ8sHgnswbKPYf8VZxSJ3Mm0NNq10wFRnT6kHrF2DiK/M71
8TL6pS986AvL1hYKyFCGIrC6Udi6zA78D7BmRCqu3ELRqqAjddRfrHozphw61qeB
0eGPavT6jNFkX5iTaO2M0OS8B+y3FgN6B09gI4HixuSKHgu9OzfnA4QVml/cZgmj
EQmHuBJQzFK/APJpxmi7t6fd7pSyNh9DL6c9QnKLuETd5V7eDvJK53RQ7cKxOCz3
zfmCU4iYo2My3OGeGfuklSXyOkU3oiwvoFGSh/nW9D+l3P4UD4fp/Sl4xPLcf8/Z
KHwLqIgLaL9MIMwVUe6IDtkNepqc+HmTfrJOvmpf6IGvtcngdQOdisZ9ILLC20z5
qRiI2wLguPKOoFGY9wPV+L7IsFnFI+luMNffHQPadXUW2H5GjZzd8RglDSpH93KL
d9DBJlCsPkonKrkA5MqejRl4qaOeVcr8uYx2hc1LBZ7viwf/jjNgJ79xABdH5JUV
j9XNlYBJxzStB8ubwMcteziCNuXz9uCfeWPI9Oh9Qzvpx3Wgd7aSJNR0rbLqgo8o
bZqv7J+I1aJkiJW4UJvE9DvdnL4drqkGRl9Z5bFLi2qs/iteKsGuH/z+83vqQZJ2
KFJkXAhZlhmS2nVr1/RBim3/SUu195bt0L9jxxJe9kxqzeYHbSDxrRzvCMjv/dL4
ObrtTNPCn07Bm4y3IOQS5pRA4YDKOUbYpmkq9bt8fciNL6YPYc0SYzjX4YFrDog5
j4lXe8y7xl6241IsXQIpk3qFT8OZiScfpT0XBX2WRBiiv/qv5UehYsn+DCgu10lL
UjvjNe3VT7afwdRwOpB/Pu8gs2tjWQIjDm9l/vYK8/ycj1QCksNm7FL6gTNoJXHF
nd3+IRXLtV2vmJVNmwlKDPMp198pVJ1o1jLVCnJHDKlUJfwJdNg6ZaF+6tp/7X1w
dtxGqmnVfk+smuQNl36hNOOJUk8FMMUP3xoq/i53vZTnESlUi2bnleqUHi4eoCP0
lClaE23SpFVz0EVFdlsdT4AIgOqJRmDm6fhw4SVvrNneLOED12u+/BhjUst+mpXY
G6m6qfe0fyfXlgoEu7WIltvb7AXxJLL4wI3J/xmBDwfAJN/V+3gKrUpSp4pL2NdV
VKZjNaCKh2aAw8mdi9/RMBTERyiRCD+lTBy6oYfRMDD/9K6OpTzqK+9Uzo1vg0Gt
8AGy+1Wfx9EJq7CzeWtiAasfc0772W3G60lD84Vwt9cwfXXjSJejQDBPVxIUsI25
HCo9kjLT1fohnBj83bvf6byngyhkqT+rpuYExwjxw1Z78fB8HNML2QjJMYsILesj
aA7xVuSosIBj3PqcnEAzXAVJbqQJDuTHhDARp+SuKI1Xi0+9d6M+O2fcrndM6ngI
rnIEvUUis3Qu2Gw9X9FR5SlOwWM+dJ7ufCPM1mrr+DYUnGbALp7CGTnLDtR0NMan
GVMSU4/MBrr9LNoxSb35cuIeQkvKqn4jKPcOgvA8q4X0ATp4bpmV78X1oQy1TF82
TcBDISA2Inuh8TokUU2mVOyZ05oT4ZqmiS9PfOcAtO3kZAXge2GI8JyOgLu4hpQx
7MqrM9jIhdhcbg7AY1reNYm646s1B+OaVeWpNfff57hhFUMwbv/etHIgyPueAzIQ
96VBpMOqK+2glehGf7kKA5Tj2Se7j+yCGH/wlz7fU0nu5/vPDAHqn7eRHp7vcvje
fAgiCcJRAG/wd3JnoUsfDF90M/Jr1FIziorbvyFaZZuhC3u9xEKXMQKU4fzmv7s3
7Aw0syONtdY0IHzUddYt1LLDBndKfZ7FHwq/L5RAdbo08a978nQvSSJL3UHBvvQL
DcyypvgkqjPoFt29pR1NWq5lGJ+NlPrT6o8vdeN80opoFycaSusd+LcpKPTrCzej
xf/rY7QWu2KhGHF2tNHXKv8hGTzKUPBHkJhcly/Yh+qjyqviffbm2mOxs+1K69rE
dkxyso6HccABmAbXfdXJ4z/r8ZH+JWvz49assgqqnQrYdfX56iKI0javJOmusF9a
5eXrl6k5O+3hRCCQo+6W8AKhc6fv3TmUTLQ8TM1m3zbwxyIlbDAoMm8ZWg0KNs0M
KaENCkS8wFF7gCc1MVnmx3uGqavF99Dkhsx/zrrCeJbyTYMpNXkENf6wQEyFjRy2
eN7iM6y0K2LIPlOu9KLD3vms70PTpTE7jyHYDEu3TmrEECr5tYvzQCUTgvNyZJMN
te3MpAnJmd1e0VZqZ6tdcgRORtKr66fAKjWaWGT8WwKvEdiNBHTgPr7/FgaW56S9
pAbHDstJw5NsCorApnSBwFCjEwHdDxVLRgGxwv8xRNTGKhxLaO9DBRxbu6BEFmoK
jPHsItRvcHGS1qBLzlXoio8jXUUBPj/guCLBhjTNbXdk84HtMaY/tKKs92eG+A1S
K1Hpf6MC+8LrCLhGMkqWtP5MR4VVdCGc1VG2BvqNzdh31V33noS03jPsXGG9Tnzo
NCEdlr7YmIHd40z6CfxVhqUJEq3+jdrtP+tR0hpJYin4ApEWq56Cy106c0wionCS
oew333s8O/DcdevLc3E5Mg0XodghSLK95tCPlg8p+tneB/uSbEcDA5cCa9nLfnsx
/OavI1nJ+fVRW8iN7nHnbwt/KiQaCF9/4sYfJX5Tm7moUcjLjps3TutmPv48Vu+g
k+u6G7tmSVsyFufylkP2z+sM/4pG1h6uKr+NFTlgC2LXAZ0q4lhAvX+X/OSa/DYS
yAcGCT7bAlev8b2rcfW/qMzqCRwTnmFdFAGsofoB8s6GKHKdrOHOAdT+NPuJRF1O
KPBsrjvmit+nhZEqtzjk4nvquDqGx8KGxsRfXDoghk5CRmjBrJLKx0hSPj3+q+f4
lgfIu4J4Cs1XL2pCsV8Y+GG270yVPNC/S9xaUvRG8LYjX/39Oz6cRLG/LbPaFFU7
njIHhuZUghNcOOR6cgYk+E5E1ymWo7eVZOwM8pnV+rbtN9ze1lfgYL/8tHqQha0o
bDFQqwvLGDsh1BCdwMTTuKNZmCCanlL6Gwi9WffJDx9gJ7lCqXTmzJyO/RWMKJZR
JxOCRVdnGXnuDfwN87mjw2XJFS176WffPnZUB+G56aVRIuYLrIKNKMcad28jFWjP
Xb09edTtaB7OKqy1eJY/PnCkmzd/VV/a913cBrspia+H+aixL0ElUVwQ9EbENgYR
Fnv1fErfAa1tUEP6D6L9CS/4f0zXN6uhKHiYk0+ckU21v7iAUELZdo9LpuVP6YLa
TtrB+1w6DdE7cPDwzx7e7rgF7vptO1/4DZ5Md5kJMuYNMKObdKCDdwKQivuhAv60
b3VmQMAf1vdTiKbEi+WLn2owb6xJJBBBCp9B5hwJpako/Pkc+/rrf5bEBztCox8V
WBEBQmQ+9/WRwdZSooyPiZh2JsWrROEJtKXQCWVKFkQC5c1tKEqpgYdvg3/jZTmj
Y3SM4Y0KNR+SVCV6poxYP/zfsQmhIwwA5DIFBiLLS1KWxgNWOCo1Ij60eNzKiAm7
MYz708m1mZY1FW118x9z+3Qa8ESZQKzKpMc/xJ9P1hGe3AhlPCbliy22NeKqCutf
cGMLhTD5mMUcZq5jTVv73tElqKnj9dETiLLJyj/TkjoGo6CzdhpOxc7QJFF+1Ymd
b8vKT66+ZYSTeHoH0G/w4me4HeRtXYugrJVQ7mfRjUsoqRBSALmv4VKSh2xKjjGL
DLysMqFA8zPBZcGbgwuodJgeGdU0uEWSlbbsEP+b43ufgQtNFT3yDkCLCrOzp0q6
ZANIcZT8VQ8+BUKNhGOjBi3077WSSzXyVldwyRpj/HwB8do+a0wtGqla9H0kjAIl
MDKmgWLnPDa4HJ2mJU59m0P2e9HvTG8SYoXmNhG3qjALbLWWpi682Pb3CLSf99cm
IWs8jiN9cLTmsvZksbM4AIWbnsqPOmyulvw6ea4cxyjcDKdnjReg5oix1XCE6UtM
OEBtUGo6y5Ik9XCrhlSc5WWv8lDGklfk92sNwd+H7np2N9fHjJo2mU5UiSbqu7NG
lpscIrIXuYPpMG0g0t6A4pfnXe3cGJOTILxDiTwi4FcjTXtj71ufHR2NWR3tySxJ
hkN513eJD4IgW7/9sTnnv3Kv0MHs23gQ3gi068AfKcHp+sgUaW5doAO2f0sm16LG
OkED4WeODdMJw55/0HqqZWP6rTZ3B8ntllwk5HWFC8dZWHhE7Uki18PglamYX2p2
BPniw2hBffSte9gwcGavRBMnXeZ9NaOIS1VFlMLAjNOBTq5KmDLyubjFWSdELPJc
Z6gRJ1CZfFntyhjWRXUnlqgv3UqIQ9t1zoC4nua1br+hAkSFEnASuRD+m80/wYsZ
JD7SkuxGQCRQXO30R2zBQNmQVXT2oc0F+8ztXnimJwFemHPCB1jlFayZRukQ+/7e
jOz1t+shSVay5tHfhQG71mh7l+wuIwLvi6453N52mpmrbqsQ9ANh50nxuPeuwAXJ
TUs6dNYaIG+1Pc7INtRcHgv3YcVWstTdsDS/lYFk/+u/UwOnPavBG/zv6P0bJ0XS
XN2pptTDltTqVIQ2PInlJqL/Qzdz8I06nIkWZ2eNhkXcCsr57D8wxwoNWyKOQNEt
RSU9To0IBSvENc6FWLCnYLvqjIQV99tgyWDdNmT3BtUZUbswf14Pri7JREV3S33X
qNut42hsRQ2/8AbzXJ8bmkT6hmjhP8/BnArat2NDlSMmaevbXQO+JPXuqy8jDUcx
LSQ5wbZEy5W8/bQelml4PmYAB7pHPNc/kuUJWI/quymQEJ1kd51KV5z0A6sFOaUc
zPoAF92aeyDuzQ64fK0jJs+ZPCur3rrC56tvFUsqXP3ZxwHrAWj2lieLcnJZV5Yd
kOQd/kkduB9prXBdHT0BvjW/XY7/Ohgrz5WwfYZlwf546LdLDn3nEcC4bq+i7so/
nCIaG4A4mA/qlFQ4VzFN3hkcfLmZtJXPBP5wnlcBtpvWrBL0CDctOs7OjZMhpjhZ
Xh+Lc87Oqtp/dgvV1GmEcEfp2H6ocFx7d53p0ytJuJDeGYypzCVhj4+hlvNiSsON
a8ycHh/c4BdDzzHw0Twp7KFkFyZqypEK7aXsssaopezGNZs5ZFJPLmxa5T4pFX7W
O2cs49Zr63IKxbQkrrCvwJtSGD/TdA6ka3FP4AvRE0huk4sJzYRdtHYkVsy3ZBGW
9TJDya0kG0N0WTcGZtXvztAdrETNz1G0FHwPwasr8aSQjlcdVDQvzYCoqxfviPZr
hHpFwf4nLoVOE9USQx0PRKKCfi8UwPFklOuYZHCUDkmX9ND+sDVrUndR7W0YTybX
Kyunlf23T5BbtAhdWZoQYT1NbKKn1IrdPQQHw0U9Fvv+JhBZaxz6FWpem5jvaQzU
xFqp3qIxYAKla88N3AOVHaFVR+XSaGs/NZ82p/OUswc5R4h7zXxZTwIyXbiPN15/
0AE+PMLc3S8CKCDmzuswqqX/8vwWczC2ZWQDrLyGtsf9qki+iYV0R/Fro89gMzUY
dGAXoXmFUgB3txjcdJcHu9+kzSy1SW93HSt88s4ID7xoJAv+GWS9aOReBl71rCak
nNYNT+DK8n7t1Viz8pJmXgqYaXGIQ9KPaBPI4ddze3tQBMUd8EuGbZzaRskKdrUS
FUJpaxNZjtar78k/XKlihMmL32j2/yNL7uVkwJWUcUijHCTfyxfzIlFodG1tG5Ck
MkCu9Y0CRcHnc084hlIeHxWgMtJ8aI4kmsZMsiMcg5VO84Lo4CHiDJLHjxD9oU1V
Wtd7j2MT2cZ/WvvoLyTB/HCJe3tchBkbDXNRdPO71LKfG2jzqEk0Cpynh7oMyHeN
/N2RiJfTMJmxjt2ZCl70B6C8+S0bf2QJHG/Qz/ojJr+6WMzPEJRwlA4lxka2FNLM
kKzgD+rzpUD65jBrVB57LRatT22CJlKJohV3/NiHOcFIdIoMhk6k4y3+ZMMqaLG8
EZRAKP7QpOLa79gmQpTgU5e7LZgKic7xW75lHe7XEwB0AGxLC0NneGqEU+ggWK11
yEKwEM5yy30JtHNmlFPRPcGyqKcgg15jLOvUDYEptIg+/B9z9pXkJYNwB8rmmSo4
7VHxoCaa8mfbpzLyqABcWH25LCzm60sd8yjHXYaK138T1XA8K0rdDuxHHPLTe01b
sCCpyq+b45vkckELTfUr7VAwweret0jLJsxXvzS6QCcjGJ3MPfF2UMIjMWX3PGhX
AhJ8JBZqj1kfHLeRVsfqAP6ULiEHf6+6kANg968429LtoqELKVWKoJWXzgdjigWA
fU16TBjPAEpExBy2IrfkLNYv94dbF5dTWFDEksM9Qxu9759n2PNX2vXjFPHvh3EK
iQE7uZsKheWKZ06jbz+pIH7xXcNNlVUndnDJ3TkSuhcdMZUVrPtLlrSz8OpVOcZT
LaFWi8PbljekMAfZLhxxgWBad9XP8xzCJmkWJNg7fbE+JPu78a4ByaQs5C9k7y9z
5bxILSLl/5UPqDpgitZRFMFVe8uLsRMqulDso5N8/Wwcn8iAnyjCtVHSCGqra0sb
Zxh9xtNqr1NGGPrmTUEmhvT8q39papwFq+PRhg4hgbRca5NUohbhP+tmajJMQYUT
FfzOk51zC4kNUbb6HmVWgE3QqEkmkfh+SKe4d+0/bPMojaLvlq3/xQEolzC1+eAO
XMok6ZPAJrH0vekDivozXwB2TIGl5RIetIAEj3LBeKHf0zxLQuxg0SRpN2lPd4AZ
/4X+7RSdd2WM2exhfiRbQN78rmtSqY+16wgl0XrkWT35Iz5gyBo3YTNLOXE1ShOV
dMWVQFPk53dkSv7dLWrbDf3mISvx7GerjelWIr94n/V0x3TgX5/ECZiIoN407l59
jaSzmz5j6PnzW1rONVzyCWKiBDI4mud0oxLNWYG6RApPpDsq3ncUrgaN93tkdyc7
4ohOt/Rf8Pyx4xPU3npfxW6FW+aQ9i5ccB2fh/acYrMeADSIdKu5u53ngQdFVZ8V
KYJK8/oj9BjWWg+DMpI1MFXDnCdAnO/Bl0rQEBbER6hZmvgNaU1F3Givsi2y1QGQ
uKGH+pVWeMF+y3Os0msiLaHsLYWIndK3R8a1y67t3fIyb5BT1+ItJ7TQIRMTm6y7
qDIQ2LuU9NhHwSZbQyadLpd4Ng29fJwzXiQ7+plBbYVfNFqV67uyKLApeN4JTpJt
D0+NJ+4tm3YdGqVsXWZq8TQoFBLcj0hH2ObgTLc0kp3Y/2Q4nEPsppD2uUpR4xbF
/gy9NDO9BT7V8gY7O1tVW8vI97vKkKwMBWnUaItfyAFt+5u5sMDf/axLLxjjJE6Q
4/W7faEqLau5I/l3GXSWbvJ6QWyVNRflfCi3afs4fqEkz2RWIrAMGUthgAc66OcH
tGd5WcFXhQuRyTzzslPcvGUbob6eQIcoZmJbX8kL670sh332zUsTCLWw+Oaj5ZPM
/exZlGnRH0mTCiKxb0tU4VvsC7caS1ShhWlzr8E1WXpmpef4r3LiyrqLz99Z16zx
nlUx++4JOcFIhsLs9LXrfKmnoenEi/vOnhdVIpXIlteaUHh+lkUtiaLzn0a/IDNs
eJr8pnYqzwp0QZnFKTtum/kGsHl/qR2MtQ7+z2fhjkvNYT7h6862nN8DdqPZUTNJ
k9TIygmVsUV53qTtdIzLysUK9wUr89kNSFf/sOgFggYVAB0hr6DpQT5T1UY3Rts1
+IanKIZWy8JqkATbOmWFp5L8XmoZV+2RSA+Ww/CGgk1FzswLIKKbw3JaX5EaJ+E4
VSTU1Rf1uQtawVA2sgdCEcUTnFwjG26M4nN5rJXb8DML0RdDLr/Czns5hYuZ1JNI
91DtHY37ME5DYByuo/Q/cqlJ6mF1Onlvm3fxAwdawhF0eVeF3e7z3aXrBjuYFdjK
171KVFRWG0sks1nFbdlWSokZfoD86HyExBLfHKMIZuclWG3bP/Nl2snZTZSEWqCa
S1vfJ1t4NQbosr731YQmR1U1mkbq2Sf1uotQDkGd0NThM9/kDRcybJLZvXKHXJAj
6covw0fUj0szFArYKAisNea1M+EUqb3GCTWFUuDyv6Jgmq72zKtf3MP4TurgG8rm
H0j0tYObWhjnkTadyjTpLi4mVhmq++uBVUjt/fnGFeiRi4SAiqOqo2BrKFsU8L4M
yTrlQttY9uLP95DeHzAww0af10DGLGyU9aTCrJr/+47d74b+RhM6YFPGnzStt/Dg
9o2u6GvIQ4cAX5l3CizA/FyYfr4r7sGfV59d5BfUIUD0RZcG31Tr+pNC5nIIe9Rc
b85jfpwXKHXqH715sk2QUDrKqMcVSiB/66SxNGn31cqZ+fUHElM3/Olk6dRzIiTK
EwuLVyeRxwr1cu0US00AdnkVhnFIgFAg62Y2+PORonsPp+QdnalFunmhXJfu9aUd
QYq6XepeWeWT0zPS8fhau3OjBnd1IM40dFkZwOAA1gWjv+I8cyOFczDopdiQYcAG
BFKXNB1ZanGJ6G4jZIYOWdXNhsYuK8ESDADwMUUqF21qRmWVjQjFZyYTLoeCH8i8
nSezbZtIo7dyS6FdifvtEyqykTGtBDHobJ2FVF5ZzpQ0lQtkvotFK2+qtJwjdwBS
xeHxS1go2AFC6N6SfZyGtpW9At6jb0EXtu2kyfqur9+5m9dsg4j0t5CbHNmZqdbn
uDY0urYaTyvs1HuBXStoUCmAgD4Lkd2GWTpEZxuKswJx5AXx/bkIWNIL0Y90QrZi
35ichYw7P6zIoIBeqFkAErqazuwA74G1tnYrHJwHtfuBT3UQnn2qdekQHbvi1ACE
STuAbvCnJJ/6FT79z/Vl1NzF7advVxwkYQLQrPb/3Au69PTnnR5Y7UuxyB/fbBCm
NBBb0o1wv+QylqkU2Uq2P8UxnbC0Cv1tvQFXAV4uf2vD3065Z4SnXPjzQPYQWpTj
TZbS1owV6eexeOHLJgEc3QxIKBYZTzyzywKeYdmxq9ex8slOEX+YpJ2J4zgutqUZ
msAg5Jo190LKceK9naOBl0h+3ie4A+USbul+ztmH2Y+3U/SMbPhcYowGIsvCxYGT
KZzcYORgaatuCxX9TSAYEHT8Q/9yEBufGgJNebnDRPplHljB+GEVAlIbIdpqsqxL
c6iPwqgm22GGjqPM3Mbj+1+CgQ4Nxbh0PuDEeFF68oRVs1fLt1ZtLz500zkZCev5
srN2hsQaxeDKK/Tnpxj72ly4Zhr0kVXVJgMjs+atdtug3z+2F4pI/cQLm8LuAp+d
5koE0M5866cxac3WTRpB/ZspPBV4OB9ThhDpS3Rb2HN1YO4aHSZ0qzjYMcRPR1Ga
6wqn8hZnOm2Qku5x/UipQFTiYcPz3jFPy39tv5QtJJxTduU/QTFnr8LkY1ABfu7y
LW2g0css5tDgPm5cc9PwwV5SeC/+DXQwKBOTfDCAncu2nu7/u+pobl70WNNbvYnk
Kmz5/1q0TTY+BC63IGoPWavphdzr7tBed61sd7gKU6cMKnb2jSI9trQmCgsuEqRT
/Az5ajhTeNDT0AIR5iXG1oPGIb+uIiKk13MltiYwHzdSz4ZtP4c8dT5GufDZgbNX
/y6cWDgUCIYhBEh6VgPtsptHG8w9RxT6C0GOf8SlozKah9dFv3K/6AhgI9PGQYeH
VUjuAM0YnocEmSvNijjj4HW3SNlhIVZifDmfsBB0JlZ9Ngcq3XRpkov1LG2B+iC2
En1zPUTS02VpuTFzcm3GJK04fpELSd8y/aEDkuqDjL5aT7YPOHQCX2E1ehBLvSqP
WZNf5mLnwQyBMQt4Dkex+p2iigc7vJ/LVY327KqiaGmSRcrz8k9ZeooHiUf9YQeQ
DgHbDPj9359fa3Owt2KvYhV6Vs4c18Ju13JMiW7pEKEUE09m08SjaM9B8Y7/ybfN
hU+Y5aEExuSmSKTBl9MIshyBLrkS5v8smvySTqmPJ2TLtcbklLnR6E0OwXdB+wOD
1y/zU2ghEsrHS4VBwZfzbxVnRUNvTfa2nDtEe0TKWcZm5+PnBxXGT+lFjCIIJREm
LAj6cEyzR6mB4z+sIuCil1ShfZiqjrrYd/30RISgchL97cWLBT7KxTBe2XYjYNAU
U8kv//fIT3NRB6Ce1uEN+jPGWpJFvovhM69xQlzmsSXL9+MLstPafgTWY1sZ+IgH
mtN/+0b2yYXAWLCH2n1gZTqvWTHjUJM40ulSOQ9KI4Wmvuzovn3JT6kD+yy/OcTo
ayuR3wFN4HpTmaIMcL/HCkxrvNnkTfXmtT0DIGuJ0sBEHTlVSrO0uR4UwZVKHxOJ
fD9b86u312ZwIfD8Oyz2zAfDAW0lSJD7pXcmdmXCUD482+AoUjNmfadnoEBZcoWj
QBt/65zIzdVM0paMFPMNjYU7xPjvwigf1x08nul29LNce8E2wFldf7XGgk14QwTZ
73xlNEfOxAmQJzY84MaVfYx+nvz8NKnYwVzMKlgeOUXc+ax1rcB0Vsi3mNHXYSOW
9IS5830wrqj6nC2VNjNiw1yROfwUYCuGLk3y1Mfo9sNcD9BGLSuH7SveV3awSwDW
LgLupqD7M75+BM/U0YZfHfpJl+jzD8e2e5gRMpx9qDL+Uh95qC0oSSF5xYCSvjvj
A4E0ky0iNmFFVVe/agCkEmpF2p1ZMWNe0zQmCaQaV6e/JsMQlQAiH6cYVMD+1Biv
NcBLnET9s6nMBvtLvz29oC2fr08bMauAW7c26l0a6L2FDXb4n2+QRQBogIyWPhem
GiyWI+PvW2Vu/aHqiilZeXw1O2ixcTT8yEGk6WPo3wEE1QUHZDO4bHNd/VuGChv6
jqlanMrj6x1oVE7inmC1xPL0yJSRSrTD+9Qz+5+K2y64+nTo5JUCk32s0XJc1tAy
IqidbkkrdR5eyVevhXMahV0EiLVoBtVkaerHyZOQNr5FWTDKvQFxYdCBCMzwXM+P
jEIvHqi0XbT+/ltxauzLMEWVrwLJehO697g+KW5IrKOHOIT1MdSU4yxGGEUX3a3P
sDQ8DrRs8PWAl+BkGnMUVuLykQAgZkdnibuBjFSIj3jR/Z3HBfSwasNlSg4D3Apx
GZawqUkYtktDHgEiro05l8auZPwXuk5kg+yA2pfgbilyf5ik3Nl2DjHHyFIdakQV
JL9CzhkMQIGAUMehht2KZpR2w1ViC8Os6V6+rBzkNGylE7g4aus735V6Md9b16HT
vWOUPrRsVFI586nW8IyURcv5Iv3lydxN6FtKPIAY3DbwBL+o8TX2fisLbgE1TDrt
UgXDYUmKRxsELWPNeHQjYMf4MsB2HVJQCwS+3+RBQ3U3zpsqGkWqOIjVxftbq9Gk
E38GwDXrpWKOq8uZd7cIvbqwARMy9TOAgutxZ3XDznzMGNJdHW9RsOB7JUjIVMv8
eDIF+69pSRG9/7CLbLQEQfMf/wJWux/oHdaHkjKTTmT75XF68bOsemEPs17S2Jgj
p6uQWc1QHBStKaTnqH9W5iWZuK0MeXCuEDMyvb/IUYGs3UxSbzy80KxRL6RM+Y/2
FVfSNQCq1BOdMvfULSvJyYlGtjdqyJc3YhTsY3gDWFijZ1ijIErzQZjwHft8UP+/
D6HZIx6ZNsRw0g1Via7wu1/610RlcVh8cVRy7ywV1RDm45z3Drsi+qZ/xx5BQIDW
K7zNrPxUe09Z60YwV569kt8/1SVv98vzDnuR5Cr0ADmN0sTln6pr1yGcdDPXWQiI
TrZmBpwFzJ/jGKHxvFSqFsYEw7k6vJnWSwV8HwehbzIXWCMcFRxA2Ahs31cE0x62
R8M9KhJCxG+evoyu0hsZIM4G0q3S22hfcVsY9E6Wl4fBoOTSW/sVHBlT+wyB2Mdk
VtPPKaHK8M3ZSkd7zw0ta5k9ffvQTmYiIL2fXQZgFOq1UHHL48xPnTOwNan7gDO8
OqoJnk8Tjq785bK9vpDOLw/BfLigRpb1xOeEuaXfI42NyAdoLpToc8+joqhfTy/x
b4zuFZUR0IpIa0T1KvyCkm1qs9HX6hDBt4ZIlnyY6ue4V1bVI9OveehpGddk10M6
TwrRkdXvcsTG2IBr8YmPm+WOqtZX7T6OKcABiiFwwUmV8qjHtEM8V6mcwM9FTdOz
k63KGKtWT2PnDupYZupQnghabNEs7YyFMDr+D81ka132mot4TLR/Uf3IecNnALq3
vM1VrCsdf+VwXqZkGpkepilDjRbWVHQEULaczAMZbylkj2HZpIGpY27duGAe3sAR
QlzR/mif5SM0YrWfMuqRU/YeoLvt/gaMQ6q706lRNqI7GL9N/vA0KTWU9/WJ3ryz
uqXb2iBfwKy4QMJb0g5BSH5cwMqujnUTv6bq7T/QenLou27L1VULfKFjuToW0Moy
rqPdliYKW38R1ddAL4epmo+c/L1PfmmETxWv1VBSEEejqYp5/pYNiyGgiw2b7m8o
NlZBJsVzHEIayFIoJKCQqzTcmvnh2/QZ7DixzkrV8lYpPQhZKgl3PX0Gf3HsXH/u
JK2ytIFBFcOJhLpSBB4DDlYFiJf7DHkHQrwTuiyWtLN1Gbnx8WN/oQjCH5m9ppgg
3e3SMVipvfaJifTe0fhqYj4lBU/PYWtvU42Gi4rgMCzO/Yvh5nobbB08UQS0wsjg
MNiSi8B3s1mvkDubN0WCYk2327+A7KKHpJBcRRKcwinsTPYaHyTpxTg3HkgbfNdt
FIsAE2OAVel+vSIiipjDUAeVZK9WKOgNO16C0RYbRdgWoLrIykybUBibPwQfrtAN
Rns3Xi3MVXNl3K1T0FtE7+ZnimBHBtu2imT1GcaguSL/EkPPrrb+RraCWX0bRWoi
b2NkXsNfxAHKm+G1KaUtR+xFLXzf2nBi5WGBWgFZlHkuTTMfPkM06WbY01iXZXhr
Qx1Kr9qy+A+p2LYuvH6WEsRLSuPPPZy4Gv7iW77em//8e+XTfxl+075MrTsY3jhW
NWyFUq9XdtNvX3/T7jIshBk6YJ55u8ec2u13AGz+1bA7AN9++xW6sGbiy2xgFhYL
44zOTFwpP9XuPt+VENLO5ld6M9vR1PRmbaf6Nn61rBVKUM7rufdlUYswZ4W+CEC6
oYEhknuCdLqIyeqwxOOXFWJ/LBVIqNXV0+xBOh2vIPWikRvfy2J9g6eQLTDpDyEE
EcQsop/e2XzMreJc0ujgPAgod/5wct5RM+npmNBLtusfba3ayELTRhVPHYnrueUx
b4NVRZcDY3FIsZTIy6a0Zrj33jBB15tu25v77x7/wuDb9yEbNB9sVx7zmhQTWHwk
rTMR+/LMZ5pXGwglL+tPVAHVR/GDwm5bSqNreErD6uy45o6iFvlrMYptj8Dw+vcN
3BrEyPR5Kv8SwAeHbSokkgM11rZQpa5lNU0Mna157yeey0sv2AOd7Wq2d1SP+RHO
cb2vRvnzumjvRW2dvB60zJO82n693CKnxWqO3OfEBvUkmEqgUVvzXoJSsUul4GBw
WOYlftENeiFZ6rMdkwBzZzCCphgpiOhicQ5y/G71L2fc9Kgspr4IrepPllgyfDv3
5WThrwyutrGfHdcFp2DXcNHZKrzbtvZXWsOEPw+gGAbv9A4sw3j26xVVECLFVxQ6
XN9riz3S/sAq8/N4tdOQ5U24K0QI60hJsCIu/JjwLWLcbVEPf2EeJZtCKMEPtSkQ
4P2GPR9a01W4PxaSTVJBQboq0CRJY2WxtWMt+kcoFJcvoVnuzt8rtiughnvOA+sG
6KV6VG0dRTL4nQo0rrQPTCu/mZJQC02LpHUKBtpmUjehuwA0a20gA8ttRkRMaUse
GsSNbkjAbj+nijzp2mXxTxX+u24XmtmmPDhevPfKCRdcvaFD6yit0R3ai+OsiSVx
ivbB7Lje1VzRd7BhHXR+aNCd7rVfLqvr/77+HoH93TPGUeE0WjgVrfsr12L9fMLj
0PXlGDBZy+LNaMo9Fev3iUvFSRXzudPxhkhF6eJGtITmHa5EMlKT7XDlj7scHDvM
6kwdtjWGEpk/C2JOaD3MiTW/veH3d1TQdZxQJjNkh3TOIT6IVM5k7LXcp9bdRIA/
SOtFZXYj1QVhG0zNyfHyryhe72SV8drZfw/5d2K8e7c9ngFPmidrs6ajK5LeCImQ
M3HkgLSdwKXmwg0FXTUR5TYw9pjX9+AJrM7RWti5372Zl32eVLPnutV2TLyX+5T/
UkbJ+vttZu9e42Nb8WGGRDA39nwZZ2XXbBG3Wqn8b5m5LGZuTvXWXOSm0paE2SCH
httlFKZ147SF1KmRWbL7mAehEIo5wrCx/QBxUrLGS/JSrmQ/UUZdyavejvggaMPW
6utha7Zo998Z9/5qoD0q2PFurP6URbR8yGEVnAIudClVUx8TPdgdY1RPqfx9hF74
zQU+QWui+bPT/TO9nAkK+RcxGRMAftNwzeYX94CsrPVezkaVEIaCjF/lJWinldu8
7BlNLHMF31Z/gnnh0TLnOzvQeo8y/Zw+EcXWadFgJnAKJJQfnGbW9LtrD5vxX7Ka
7eiLp86Nkq1S0FeJBz0y3An0MuN6e6nzX6uMfqBbTPbIEg5nLgq1916yGahNtZAQ
Hw3uJAShLcxdYjSCR+ozQYRRzjQOp+OxdpWqNQLDRIUcymHZSFzVZFqnkDBrZM/s
tVoSDSs1r5WwkwEOYxcl23PtvCE+OR3t05qNihagwBN4V6ywkom54pNBvxCf0Jix
E9dURYR7H/gIgz76sXDnMwNrA5V1dxyIshA63No8rSo5zTANrZzg3dysJsF37gqu
GDkJ8RMSoeby1hzJX9GgkabSVrb42zQf5gek4D+/zqVsIEy7Ik3MnlL8+0HcWdi3
d4aXrfQeIdPg/o8lyb/V083IZQ/QY++1J+XNF/O0OFWuKzbJ5Y69pfy7zXXWxYAo
/DxMPQMOqWCHsmZq8VR2lg7EuRcbiUQte6ESaXm9YLrYkDGucYA5UcwEs8rox66v
CXdkKzM1YBYV3ZMAfNuLIHNIxCJPWGdgFfhNt2Mg9H8NEWFOC4dnhsvGDS9q4g+Z
xQer8uc/L+xfSIoE4sImdl7w4kqFf6sJCs/KrONS5LMKfsuW1cwscxPtwjobMZQ9
yJ4K3rz69WBztmrGxHOxqjOXovKlul/Uqm+VO7mdLnghBHyaDpT567K1mPmth/Dh
DrcU/hdiYBxL2XIGRg6XoKsNmmb4hb7QiBiw0EVHKiva+JiqTa8XZdk+BW+mLNIZ
WsOmMS06T7q+izJU8I6m8Y9CgZQwos9f5AvW/K/Khd7qNxvaLQqhd0otxUmTRrSU
b/kkxFjNxuX86siZtoXwmmvstBaSgfrMrcF7G40uDET8onAG/mdT8DH1cbYqxwm3
C4a7VCZrlgNoE4LHK5mpj4VfYGFlZkMKvTRD2NR7v2c2iuuHsOHyUFMCJQnD9JjY
mfZB+UNhQtay7QD83A1nuMi55P2qIaJUQ2krDBf+/unAcsqGgxg4bXsBt+lQkjWt
H300Vv14lhCIPf6IrEnEukWiHwJJPH0b05aA1MEfJjzzUWoOMc2amPUjXHkm16/i
CF5Bwkam2ZtPw6kjgXThG6mkq0A3lqXkZ4nJ3bKKX/KF6msHgADtc10zU0hjXu7X
9DTTE3/fgLqcRJxK5Dw9WodFOQs9cbgHOY1qOp6D07Ll916ZuC/sPdW+ZzaYkVpZ
3eVDohZp4MNsdq42ARpa7n8BnCA58hUsYX7SBfLYNvXreFvsyKRj3K/6ytBTNkh8
mUIXSPu/4UzD9Y0Wq0WMcI0bJ9NeXu41enbEpKR6E8vC41+AaQMXpN47OBv2w8n6
+Przrg58pRIMLAcQ3Bv7cb0BKOke1QymlTKyCwqj+QRXZeMkHYeK3nNTTS+6qkQM
euhN/DzmDciVEe3F/J5jfzAg+eDJsqRrJkXb41drABLrg3iUHaVILWOBwu5oJ/8y
b1Gmb8D8zcDVPRXE1cLTWV32L3ux9hIADirOOABKY/D4puQV8MEWCl0DyF7JQ3sR
4hVr7r+SNzDPwZPfe6pHULzB4A7UPkjqu7kRYhC7CasqRbsvTcXS4iMQMh4ucNl3
MC19H0yhUTzAk/Qjj4iciqeq3VZdG9i9ibYw4EMoxL/rOEX5/JoV1jj8dNXp1DN9
fL+ezwNqXf5eW+O1FNyGmAlpkc/+Mhgz7DVp/UjG2s1KF3LroCpnaIusQXcoH8Q9
c1TJ3kM4TNw3UDvLtGQBGhkLP5G29tpwb08mjA0Fb7tAQ2fJiHOifCLL60SdkmNa
+OOmyvCIXVVGqYOnaX1HXPeJ10Q/dOo/gia2WVRGY1acqjugEwvDS/ndOpRarrUM
v3700V5wXi2HHDf76HaHz1z28UgufJ1ZusGvY0EiSNrwp1lXw1KFKI1wwYn8mAXB
+QR6kUA1Xdw0xNvyjaDxtZY2TrmTLlaBgCDBbPNm0Sbou3/UP1Cz5fxNSP2oRgyc
Miwij8867taEfelrXYQVwiA6LY4LdGW+GmntRozz5tskAt0qO0/Xv13OZoWQOxIK
nWivBePe93OuO06tAAbllZ6hIAF3W3kQoL/lffaD1yCdWM0Se9Zswf00E9oRqluw
l71Z5fTrQ3UiPbMw1koozYLelmr6M+b5AUj+j6f8pHFgvlAkIFVaJNK2mJ/eMlnk
X1zbooW8N6BuD2LkS7SrNvDKH2PCFVPe6/OwuCsYc+9n5LMrHDAdzrFAZPkmBKP6
WGxuiRdqXEdRmPmOAkjCB3ZRpqkxmKWBfyHUijIqyjoTxIF91kESSuEZxdMYYQxS
Kl/UIk1JSoBMQLeNa6IqS88V7HYzblN/vdcsIZgBD5EgMuWA1aYFEY2nmwja5/QM
muoWjYIUz8qECL37Id3iGewLTQ905U6hkBgA/P5MSk3C9BUIB+9+/lMxD+fWQaTi
9PSVzcw4DT67M08gOVfMHoDngkXUNvs8A7Qrr7Hxt0ZZAznNZivKMQco8LUYKYh3
n26S+b9qh89bVAAjGe5h15+H/JnxF2kJG4//uwwY1/WLktUeRyB96BxcY47VWy/P
bRBOEUJtk+PuSZ3sS5wxrsk1af5boeC57RfZxKjnAcXCbMp4mCZo6eqQh7GGDFLw
5NxUBEY12dfW5D3+097+DfCeYiJpXtF4Rg+V/qP6QAGnpC0+9PkJ3IJoAIzfe1oT
yLny9JQsllk/cYMAIFMV+mrkTUsjaX8McLEbkkW6M/5xqhC/LPQI5x7Wg7hKOiXe
BfP4+mK5QWpNFkR1U2jsJDgdRnH2Hw6/KH9hLl3OGIeT5y/KabsBfVWbxoc58S/e
ccYxo9pcTcAeiLiuqWP8Sc3qwe4b6jJy6LHxSyKia5Nel7VK1AwMsi9jMY8fykLC
8FYmLnq654rUvUY7fYif46UWZ4ORgazlvRXp6L8f2+kbOm20utlMxKJajrprQIZ3
6qaRTM8BTlseShp/tH8wUIakZ90QGJnB9vlkFn6N12gskRNdgzUSjMHDaisMMM2L
lAxUE0KSa3t8Jc9KkYsmdFJ6jp9sHLVwbix1jWI1iMFcm7tJaFL4LD5xfiuFDlW7
RY6CTzPTaiQVhQaCEliCGkc/gvbMrH0UVRfqYgSHw7v1lGwiFHh4ImpqIUGt3/Lj
6gvagQeeJriEyKYOL7F086Wdf3ibYSEEgQuCSBr6THWMYCV49+ZOxfSivzoPjKTS
e1ZNlulm/6CN/K4Czg1ejrTmYSw2MocnXL9V+DTpLvnx55WajpIIgWkqobKx3Eqw
XbxjeYmX4X0QDF7gkrYpYp5rMZ0Lvr3L1TdSR6m5XB2nrl691pYGtJgFkpxl+Y2y
OwMWZeYgb3yCa6r1d6n4jzXh0B9WjxJSklebJwrag0h2cfZjFrW4mzmhH9b6f1l+
rg2jKOI26BI7mUcYWSjgSTSRf/w3UOUnYI+Fe2lkvVldN15QkgbFhB75a9BQslbE
fEwzrdEvYbXVeDg8yOBNJ5FQLmtFAgX6tRml+kOjhmdoZRhM0QBk80a3+Kq49RSl
yWr1/giDRH+qTATpw20NQ+slNjiGB9YUNferL+9xJbOz4zSm3H72lteCrE3Im4Bc
EHJLa5BTnOA8+XuLQbm1euQRv5vRFyCztrAqagupWkYZ2KQBqq1tyniWV7WXM2OA
D6x8EXIry7V4px8gg0ZEsfhWXgrs3faVNT2KSNHH6mBIhX1b39q5XYxDsyAkdBuu
wuvHmQPuK+xOIOXyLmmfd7mG/kKs7f1EYzRObPJm3tBFycJIpEHa93aoRz4N8EcA
L93ZfkXi31L2qSrQte9brIdGPxlYEY/ieR3te14yteTdDpcChyF8GmvQHGK0AFmS
rMS7WA3ulKphD+8XlL08DDrOc/oAjXxtx4cwK9muQ9MFPCChny352HZrq56AWmAX
qzagV4C5mhxa9Ri5PUZJu8jXWQvwwLz9tmqW/FBalHm2axyYPsLH/TBjAZRTd+HY
DHdXs4P8IoLdYtl8xfgcDYaBZSseEYXTLLPgsZGetjSIHWj4595fFx3UPEUcV6/b
lKEll70gHMqE8WWLW8IR03uVSX1S2VrOU+tWVmdBpFixHPOIz/jGfhfwrhY+SPrZ
9p2r2xFQZIXvlNGVT7VpsZPK/RbtQK1DnzoktPhKNBnVY+AObv7dx+7cCPooW9jg
fjHrjwG094hWxHlY4vT+9cbJZECmanFQCJlR7o+FgH7zJLglLLVmy9CAiRGJNepG
fKsiV/gPlk/z1lAtas87o5lhaS7Ejd6iS9zcLS7RiSeNcvOLGQdQCDIfsPxRCUjf
Ea1ePbZt05pc/pgA3AzKymcPhPdyFgHTN1gJzmla38tV/JAUV6bgt1f9WRhJ5+FJ
PHjFU0GXBoAn7HBjGHkqKsQcvmrL4DviCLz65WMTEaF5dZyoT2ovNmtuJJuWfBnM
A4EO5FKf3yg0l1MP4ExPIoWM27VjsOPh0oRs4S0mWzpRUORL+Zrq1OXSmOaGy86M
J46EZbFnYpPRogasES9VBLc1QZIxBePfW6NWo6hXKpePEbbofkhhdPpG/o917+MB
u9ZESL9S0a5f/mRUYAanapjzRUk1dAwI0Whn0w88YSfm8oYzXMzMxd2+mNU840kR
gQ4C2AE51DjuUp6oDp6VMkUmFoKitJqCrVQzQ2H1+kA6RJydscqIOWYpvfwTgUe+
oG2oULs9+UzCLtqzAroVStljmPZdb+tn0Fnde+ubets6JwbCj+JsfbubL9uu6KVU
RI1iYO1gJruJp0zEaOkS40aprpoa+axt9elEiksoWxVG3vj1qmtruB9XEL5mllCF
PD5iNcdA8wihVVAekveyx4UxGSAaTdomTl4OA+mQ1z2iS2Fxx3LZ7lBL1L4J7fXe
4YQvu3UUlRcV6nqCSY9W/xbHuTjp1J1tjtJuzJ8KRdLJtk+0/JuVKbBepPZkHJ5W
sDqHJnIfKWYNKf2Dn1qpOBI++LylEr11ONgqPjE34/sAaaH+xjUgPDkEZ1q6l6KI
cNpbcoGOgZbaPH9V502DfrMlolm5e70kGSCSlPon3XdWb3U58RotWVC707vrvf6t
iwFbGfl+FEJu2c327jw0ADd9lVsnLHV9iGoZxLsrzJHWQRx6eVjowJy5cbEg8FX7
99mp0ANpouL/Pm8aLzQo4GsrQjPY43JmbQk3iONsosgOCClt1tAOhZ+Ha7rur3ok
st+Gj/y+tFsQc9vkWESYOh5n2XgvwZwsBpE8SZkUVFZzK7yVG7a20UQKGcLEuneu
guJTlaaz8JrwWaNVEgBcM8sU3UE56bP1CTGhggMn97RCbFOE8AQFzWs49sQHLxT5
FAOrmGD/606brl1tF3UQclhbHSo2Ixu90irl5ZtDNzFhPIu9hh/fp0P97x3R16Dw
ZYEiNHrfb26du0En1hmY5Yq9Xgtw5jTaLpG21i9Y7IQW0LpBfclkKTnlwho/oyrK
wfv8VAzgr8v27wjhkhsvrK4kiqYclC1Ve5zRLXoGwmBIt2QcXouYhvhZtYjRmX4l
V+i0B1RZJxFAKNRSvbxut+/Crkih9v+Wfq/knphhuXPk3uhbO337zQVpViZfEexI
5UJoRoVBulndolOEBNjNMpkoOWjacHtiQ1QYlm+NmmETw3E6+WJIjLFsUvnUohdw
I22B3iQuTALBnve7f/K4hgSoHIhIFmblZgSJc+9tgOwzAdqVlk04EA/hMQssvlQj
Tu/riqNDp0iGZ77jBopKxcwQ8OqAN7OXuEfxrqzeZrr5PXmLHGlL8g2f8LFCmo30
wgc+KulHBHVkJBOL1IQxQxTfym4uCBR/aPnNoEJ2ZSsRmAz3O7OwsWYOfmOI8N8P
vCIztc83C+1OpMfNKnveNPuXeQlxYvuzQJxGhSs9T0jRITtnPW4mYwK5U0UPCWbZ
/70aGqSlaGiTIr5Z94IWDt3PEr+sl9HpIeLz+KUnLbw3pa0+vyV4cz6nyzQx8h48
pW8K5q593U4PWVUiNT+di6zBzyR8XM6vX+/vuP4TrLcOcuUVYnEMUn7RJiDJUea1
9NjvFNLIfLs3b3NwJ7R8Am6vnYzJ4b+o/sU72qwyHkgpTg35r48E7F8xLk/SxJ8S
rcTmBy1R6S6TY3LQWu8acYBx0alq3cyyyNmeV0vrTUAmKnXojsWLICGwM6WFPdSK
K1OBMbzCeTUdyslGEDtj0PC//CS+yw1zXgApENZN6cojOpudkNUqyFxuXBDHcjp1
0txLd2dWEyZn9HhkrWL4LALanxA56HHzWgItdp6czROkDjgAtLryNkVznZaMqNQ6
UBxIZNWgZ8GBWzREZ9XY4/MEedEnyL58e+jIPpXvFmuzc7HIyZ9nAgtLJLF2jAte
NMlj1q0vNTxFKh9b++xAKQuX3Kuxuh0W3SmaSRO+P/VGpLCsQaiab9/zXaXrLGWN
AyhL9ckdRVoFvdRRrlzmg62UrYy460ObaJt9E1XKqgyVWwqh6JiwlLCL+thxui2F
SBT7BFRNYUy7MeJGIwm2GIy9uYp9RNsTgLvOy7JUxuaHUeDygunW6ZRz6WMlgAkW
U7j4d2aWWXJ6YZmxWoITdCH1eXV6VEuvf7vG/7fYnzBb+a+ggLmKWLcW75FvsX6L
8SREdfWN2kiCORgn7qoe8wEoGircZ1M5hiwq+ihsRaJEFahX9o9fl+SuNlZPOiT8
hnyctmm6/699sZR6BApErFFPe9PRIJVos+CxvU2whBiJYnEIBgjAS443T0biDzaP
iugNmnxfnh4z092BCo0eGjyMQASYxO7gt4T88IAW73wa7eJ8Il5tpPz3mKJNntKk
bNQkV/JB9/CEDVwXOoABSId8LBGawyvBegpFPIkV11zlDM3YggD/nhhcYIbq4+6F
pRDwif3Z4FFN+eC0NJD1oPen7d6kb6uTKQQ2sFb7ODFXI04egD+07zniCKoZ7N8Z
TctALSB+NLB2fITV1Rh7lMImLCxLdEm70b6A+wBVJ6XRDWbMjQZutxblT/5Fi1wV
A+fn99PfkvIeTfnikytW1nZVKcMLmXPBoXB9UWALVN63nJiDIDaHHbLSjh/P6ZW1
ZxJShLn6s84urdOrSZJX3jrIFTHGZpz1jEgjp6V92/BsGoXcfAScxVCgqpkCiAZ5
5an0USbFrKZVMy9lc4hTCfcqnB/mQiUwUkH7O1gTA52nz7Sgf8CdQCebsre05exI
KiJlD/+V0RUrLJ/AjflE+6+A/LE1vTYbeOzXGfCuMZq7XeE3yiC7aS75xdlanSJI
/DoA3yj5Us5Hs2pn2jYF7DLOPRpG2/hnOL0Vt2hp5cnZzlMpmsxu/CmeQheVKN1f
35AZPkwuWMJ6WhcNJF3VOKeXM7lRKQjmXrfU6enhf/SgzPV8WP23a1xjWRUWKp/G
u4CG05p5v3cbA07nCf0kUJhqKr72B6NIjVKa/SxltzU/RzE4piev3lkN64mv06/E
sTjfRKa8k/vWQw/djcmz9pSbEI/zU4LAydLw2ihrxA3ebOGmG7Idz+dV1vCvKwnN
LO7XJJnHEMi1PM+1qblnSvMJzAJlc7A2XIA/IfG4McNOLFOV7A1OGPcoVT2z7iWf
pj8fZYODWisn/NEBdV0dGHJG4OlMPDd5GuW9GfuvplpkzO3lqgJXdNh5I90KNM3F
LMryBzWf9EaXJBiGB8zc2srf45uJCj5Z8wurnM9g7qI5gxM1MYGAzNb2gVIu/nqB
33kEfqygusZvqWdfHk/JTE7ca+qGjS4+vjiobD/I/5saML8DXa/x8Xjvpm0a3IJb
LHdb7ZQ4JCnN/IBNB4Hklo6i4O71uK/fvykjyn6TK8XT/CEH6ft01UO4wM2VZGku
1U23KaxJeYO0zyxVB1/RgJbojzZpaPkV7KEs1+7jv1HJf64NhxD9H9QIwtkhYDyP
D8aURWeQm0FfQ1Z2gTR3uvfz65A9f7b7jDqbkADop3S1A7XykZqNhBc7P6FsmeCr
3FJTUGtmqRorN/6DzCUfOhUkcORxYVtAX0EtMhqZLEn7crbAl+7+9F7M7aAE+W/P
y4c7RlAaSm3zyqLgTIXwPj2t8DU1Tlhya2Cjw9lsWzfbqxbO2Y7+pJ8OItF1Vsvj
kMYT3mYKVtDM9PvOrMTfZY/vxKJEnfCS7hfZsLsh/D1/jdYOFm7uaWwG8UOMvm/n
pRDCUdntB6b0UiwyhdQwd4SPN/JCiQWkQNN1gLwXR1cvFfN/ulq8V0DUDGoqdTo7
hwZpsj7sDxhlSXWQMAS6whUD2GuE2Ex+T9f7co98Sg+m2cOuSCqjYDleQ6Y/9bBw
IfKCowaoVRi46hfNNup5tCHNChJNDHj0kuV7b4j7XUDTb3t4qpB3B9YhaCfdPfO3
f+w3A1zXAnsKQjudF3BLb1WbbsZlp9XyhJrDBMdppHw2nU8B7K0twkdNnWchmX+f
Lb45U5zpoGCu6MJdFaig+OrMb5zdQpHhXT1JRnF2LTqzFCPiD11mrEMryzpiIsfo
HWr6CYAOLBeRvsj8DTnscz9I1cheqSAz4mTb4EIwbUybz9Mxq70OUtkE7qPb+9I9
ccBb1zwFFMfdQgWS7sz3pBzDV20CN68oykAigNzAP1491QKJasLbYqXrv8ptih07
E2AO5JFCoHs4+zzeGl0N18Sr543VEcRc/sHLSiKQP+juUsKWsCxIfkHpISai5LV+
fUa/rh5FnWcrYODglDWu6j/rfrWDqgZgYp+lDhtZRD1zoC63e+i+23ER67H4CKAO
NNBVYEd9trqch2e4YVS1E6CFtGcLarlXCNLjwrpTEAPn4n+TfV7CXaJ1mp9+yh4+
J1iSUNEzOQryuiqcKy9YtWDWtVeP6M+tMJ95ZRclbG9Fvzw5KjclJwSe3SsgI7gs
+AIR5i/+nufXGnkF87rDptqOiS03L0XspWZ4pzN0EUZJ0+dU/agGo9AEp0pDpwSx
34AkkYz4o25wETD3SdZqzGLwVU/l0duw1t/U3rHmh22SmvR2k8ERvjsY4n/Y9gtg
3+bzXPGJsLktVAJw0SGVKlUkRIz25bLlsCveN80XquHFmHTvOPwk0EdtFcfuJ/ei
Z2PhyQ40a4/e2d59e6poXd8PNLx2SKpFl6gWs/soSv7PAGWnZOGMHNb037KWIsiw
646DNG9+Tqs9XuCoVudUwLDlyNCmkhGDnUtkM9hoPpqgqc6nikj7JSZU61TLoXMT
mfZ0yswhiKwzSVIRt4gZqJXdhAhOEBB7O6UMPhW5FLVWIHxXdeldiIzFFhFvf/A1
mTy0yy/kc89gJhT0bKbTwTkrsXFSsQSYy9I2CZ6vrCs4mctRn1/SY2q5j3saxCL9
T4q1qGa2/uls3GFZPeoMgrAjUoO1hOJZ7nY9vEWY9I1aLCIs3lNiMe0Cvd7qERyM
ih57nde0ZqaBJWH4vcYsSglViiYPggFBR8FKBVoNT60Vy1amaOWvfxEwfLFzWzmX
hlP2A6kSpzSpSrwX0zKLQi0q0MUwAdyh0bFTh85XozP2u1nAbDP4rXz4+jgO9ybS
JnLIU3C/RpTx59CQqmwzuMo2Q1qW49xtrbncvBqhBQsbTUz9u0ol5WzEG7KjDyvk
Dgn8tqyBpJJkailKzT+M6PtOLuIFD0IDlWOSAYF9w4Bp/jmyOgHWfxK3RbhCIZfO
aV+guSo04zfdnVyqGLUDa62/vpCgI3+CFfCcnbzh/vzfZXvUObJq6UB67wu3TdFY
IexI8bB9InnkmIwUtB5TIhXdQrRL5fLfrP9lkLBVfZ4oJr/LOGGreXHsGnp/42VD
RRBul40wV7N1MHzCnyXAzlIqLwzJN+/G8Glbnf1q/Dt4yxwTqHFw3JPCzQYNd42D
U/n4DttzB5qvxOr7ANG7l4RVXEtm0EVI/Fpnsj/yeDNiJfcxeArYbffKwnRZx4Uu
EU5ZftO4Ms2BjC/HW/Ra8uqij8pAuEkvXGrHs8amLsFls2EiwKPWgmdx6bFKN+ms
ujz9/vBdjW9PRe+Pe7QgkAPsZrdiDzMo2dvmNyvqS6nt2Vijtmz0Zs+TMrRjKtxl
CzZmytEze//eklaDGYq8LIYiB10QO8zuCohYY/j4j1o9oxRKuDKhN+INdR4Tqhf8
iG4QZbElkiXKBUDY/OkYTAnTXaebM+CPlTOqWA09h9I80GcC0zzwtik+kpEuZlR5
PxOsZUXa4g7iyRCrJR2IRuzVYlBMxfZ/ckPMPn7DPzRn0OwbJGRClgVUFUfz9DXn
RVcaNC7D4NuaEwE4vBNQEApSc8ayOzgyEnJfa6gOQBIym5fL1jg0S7Ivp/aZhjf+
3dPNmw1riyTw5C1mRy3FPJeVcPfnPN0Y6eF1jVUxNVrGkP3jDWAyZpT/SyjL0Wgq
uANwJxdfdOoT6tq8yA7sCYGUpSY3dAmgiJnB5CggIWhMP2CaHqPusP8icHLr3NOb
u09wADBLMHTskZi9aDlywlCeg7h8Uve24KLy0DZgd8xjU8ZrF3AOOmRG/FZwn4Nx
tXpFF8vy6n2QcaU11SKRdVMBw/m26aESg2hmPyzdEQMLUw3M1QZohVFxKWMbPo5z
BM3qzULtMg+aYuBu8HSl/eKKi9iDKS6am60w2ZIadZKeo8pFrCVq4N0QJyjpPwln
5vfdaJQQwncdxjxpG/wMEBQ2kShTlJDvFW/ZL8tcNZXj66A4FWcvZeunaPIwqrn1
+nfz9zqhf/4JsDCKE79Os8vUWJgMPgEC3j6U/pz1hUOSe8Kt8jKuX6mXJvl2Yy08
8RL7XGOVvZdxnJYHHpZy83ZpU7m94hktzL9Pkw41qS4K1NxIDndXZ2/vZWy19Ygl
cwSKZXoeruMAbyD5VuE2nBb+1Va0GAV6wkpYPKsIlAh3gM6x2OwwlZs8I3lFaV4d
pAlvZBuKdY/Epd7bqgqttEMU//7wLt+ftghAy8HRBMPhh8DjGRpu4vP4z7mRroIl
uyYRCKVfwwx6POSyN0Hp8H6zS2+iE1iRkYsQCHUQzYDz5xFQ4QsgOXl5jNtDeBfH
VxxJmxWk93XNwYsD361r2AiMICzghrb81SqUC3Yt13fYFr4uixcyrQTT/vM1FQMt
pGrx8EYCix20FjUva+Qvd2STk/4UMFMkYYRUYiRG58nhx1xbPVpLhOw5HqK7H4YT
FwnfRTfN4WrxbJslUXsZo5DyyiXc+QF7UwpTlTagyLV62EGleO2BpmL9Ixky2wN+
N5cur2xNYaFKIim8GUo30uWvYQ9HMlGPRZxPAxlBD27Q+/l9vhuHvLYInCYQaODo
P/IDEb8M2qz1GNorLl+s9c47avLQMZrBy4mxO56Y/IBOqHHk5LB8a+j09FS/BTJC
ANHzqThV3UqUFWja7S+q66ZXkIxKYKQ9LH9x20OsirMC/FcdALjpj+CgQM/wfTsj
p8p5EuOleU2tCwlTAWGL02PPNHr2V9J8C7fqRM47uQSFyDY5hE78SXAnHRU9w+aV
Lg2MXis+mqHGEn79ft4wDsHKL/j/BLtdhwYPct3rpv4dDlY0LPcBpJ8blAx52iKS
ThTpR/bEDAa6Sc68+tbpzZ6t1HVH1BWljyFghd4P36TeRpDSB5xaH1roPAU4x7L2
OUNRfqzQXKkdOJgRbyq635Yp1XGLGXnW9qiFj6PbHeBiE87Sn9tMk7Wi+8lH2nQE
g7AnEVSVUh6by9O/2pbU9kQQFIAJdePCRDh9IIErVoPrahZxt7xd+8P+6ziXzfy0
NwrM4MbCctRsneRfj1iwwafF/lw0BWr1cbLJZm6zokPudezAVmuC25YbOapvj98X
NEX/Ii97qVYBSbbKN5gbhotWElDerH9v7VGLwlKcC/wEMYXJge0gzfE+RT6IKu52
Sxau/qX0wmv8jhrwP6lWYZBFCSnHY7yJBs1ayZGeN1yho+vggDQynAZDFiXsYtHh
U0quujpObw/c2uxhA8kfsCfzrdAnH/tLUmfgRTJQV0uaumWJNMeBuFsJS8AmhrLO
go6He8JaqIcA5xSCoy1Eb2/ZHZBnvbglhqAhzRJXxJlVSMXvpYyuSe0vg2UzefA+
jTGaYZ9RUvsw4ZxrnLDhFyDv9CDGJgljY+80kjPdlf2AJrv9Zpeg3ewALLZi9dOp
LRFbWTPofqEMHE8mjZdneO6tq0+HEsblcstGvrSBinc9Hyq1pYqRHNYqrhGbNGjJ
uskQYiHLNm9RhwuE9yfoiSsppCj/jOGhCQa5GrbbUHIdQI9sv4KocSkAZsBo7Inu
h9dYPHhsiNX7MNfkkbs81XTcASbGtu7G4GgcsydJhbN2z+1grFHbyc32YIeI0wlT
mQm+KQg6LTazLxp1cp7r7qX1Le+5Y78A3YSHkl2/O1ATHCJ/9+JHHNzZHXZ5bEIm
8/LwL9DC4mEeySE3xNxaaZVM7tqYO1qZmIenubKUwzvW449VnGdikbFz/+h4UaEH
0jDhYcc3rCHegSBUN5Hx0S0IU21nt7hXRK78nF8FCVDSIw9evx25hzzjYXLOFTfu
O/Ha5yN2kLJRTlMjafnCKdCRvTEqd/+g1lq1BRTy4P/G3bjQhZUMI5EagBms4vzh
k5BQM3Sbc9gnls3HQksC4guDiR9it0/eaqEvXRudaHm/k5vNCe01uAjDlCbJhHLH
UweweA4uWF1SpmzZ/JvxbFV/YnHy2SHSpjzdYV0OZOBOo4bNGCqG+PHWdcK6TZ0G
JOdBG8om2qxfpr1FHE8qZTZKI1qMRZVQWQ3YS+LvTf9rnRTVQpmG872Me3b2LXG7
Vo5c8cHbKNv9oDW8K5HHxrxUc6+BxjTIPj7LjtK1NnnBxg3ju0KZiJuRzdhUDdbH
Pr1d10Lw+i3ddGZ1TmPVa9MzjOG/pfVA1KTzqThGYmU01msqpLWcPEqmJXbTByd8
o0hjqP1Pd5jQ8LtVYf5vUFbO87Fyoe2+9RiZA0AnHIMr8WM7AMNUlyRlwFLWFAZs
kw8zSfyLNTaz/y6f5mRwqB+Cy+NafPWDwq5xwxkRSnO6CVEHarEqi3Ex4oAQ1wGX
4y0R6/6OSVNs7SnEMvHDe514HFJ0yfswi5xOoftaNZTqiOpHXYHsd0j2hnCOgugE
nj4ElNVoqDaLyZRXqmwPDYLxxWh2dm4lx8BU7mhIHRMjQ3bFuWzT7QSsCc78q2aJ
LEzvYm6P+vTjEquE3BdhZtu6HiMTn6mk1OlT7+rKEI8tG54fciCDIj30kvK8novg
rTUHVNQ9HhP1SL9SlGhQ9F5dK3pV0vZy4RKCTJwu4kuzLTHr+RKJAOrDr/MSkon8
MS92K7XrXFy8ciHVj+Q4pw03TrZPUyTh3tRR6AebjQb9mmgwPkwgyHnAzG6R1/Zc
LnlTvpC3yYlBAhN2Eqr+/cBWT+i/9Y2fLlurgXSRUW7rsnNIrtbdtYCvR0f8LdeH
OB9UeJp3hHRIGeblhghM+Gy9CWOlHWn971OVlVExIjK0CR3QVdDTsdCARK8hx1Aq
bphF+PGlt1JrExa489qG7POgIob60YuzNuODLVDFBkhNNa8TkUCOL4daWPti1K0F
/HPh+SctaPrnO8SKpvnXqZf3kP7lWAwDs546DNAPjRg9wav7K7MzCECbZz9MZEY4
5J6Vno8okJ2u1XAlg/pGt505v8bbXlI4vSxyNXfy1qvhm5fjFTV0wAuXGTzy/pOw
t4wAvfNqhT3Nkk9GvQwkB/GMZ8Im9ytGwUTUT1RWkz6+6/LBI/hngeOGMZb3kT0p
niKFuA23P7b4oCg0sWgzGt8N4UF1idHOLReoBYCiOShyDa0Th9fo8t6f35a97gHC
V5jBpo+sarzUH50x4U+XyUg3uHaNxNGmGXjj1ZAj0VrwDNkgcGAS+Cn/LA8AR7JT
nHA2RyZVMWxefyyyot2GT8AulHJxKBdu32ZJwyMym2Hm/D0QolxIREqCaaO/oOyN
zHPcaAIAFvF/uKLiNTSmsiZudqtJCtrIimZgimCFfkVTq9JD3NLx5rSj3p6gkM6H
rkbIFRrGeOMQ2fn3aU6vpFUoEGjfBKmkmdngp3M8Hvoxi1S1e6hhf+HcjeMvyj8N
PnS1IzcvxuCJQ+RWFqdLYCai2j9+K2blKEsFoxGZmCTLOwzhRevPrEyPBesHRHi1
CtcYv1X3mDKAQ+veolvWcsX7ije+H6lDQ1et96arEUXAlmdAqN0eJfJ8+/Ii3YOT
OEcdY1uoGTL/U26Ade5dJ4fTUXy4Jetn/I281XKp0VhOlBEkg67SCqTU6pC1PtGn
nqyThw1e30HOiAcU0mfMGZiY1NPb6n5v0Af61zcTrTRgJXU5IqcYRo2rxDbdvL3Y
y90gHW2yiBYmaVaCHkqn0mINb4lpZNdX6Q1KKggeY96P4Z1ES6+ffRtukCsCMKCD
dSC5wgNY8Udrbz3tBkfX4N9n70xlxBD5fMQpH7WTOh+ExyPts92vQtn1q2KO4coz
KxpD5gEpw+SPayK7VsL1A5uinqPjig+kezZzATyJc5836lgGsa3eJavlfyKKjMct
tgBM2oINBs8H2oU0sgs6FyjLU0I6CMPIT39Gf4YmaswHIN/woMSCe1knspd/dBal
ce/2ItBIMECQLqsgquSDb6J+MBrLq8G607rIrbvF++NvDCn9c3R93Z5Uo59YRoMj
kdDx7pIuY6oeGnZD9Xp+fzxiJUdLPi8XF/VbW22jrtMFHfwa4kJXmiWJj/vad1+3
IQllN1Ud8eySZqILp5dNYDhPPi8acev92bDcxzRQb/qiCguzHHudgJXq65yno2p5
GiKSbVzXANzPIjL5GNuGZNEeckmLMcaJahpBhf851WuWaPQD83KzsL7SIGzk+SNg
q/s7rzW+YCxhHlNqxDnobcuG1ioMgouZITaMPE3IS7rvKUd6SqEjNe+VxcEfIPuo
Mgp55kQ1oKxVTVaKqQxEBjP5/e0wrrRoebVOra2bfbC2sXex8gXb1bwb/fH2MF0/
MLPRzwT8DDdb3fBUVHF0cPsIS3IpuWXbwlFRAEb25tEV3iIzsfGb9qb6LcZyxJan
ARCtO5oRdkKqP/qtm2bVvBGAlXyz/A0Iwg2fXdudOgzIZ9J+C7TadGXPM/gXbhC5
J1uoPjjb8rJPtfr1ZrXrKg+BOvJ3eoWP72tL/cBbfJJqpeDnONeia0uaNRJQWTqK
7JBmOX/DU7qUAh2IJbBkbf+eI8VME6PmvrGbH5oCa8aX2SCB8g9Gt4vyLs9mG+nu
CNaYkEV+zlst2ZoUPfFSxwRkUfOvrRvFPoYaM2cBqjGNdNqxjHb/rIQCHpUMJKkr
lzVSdHTpkQq8aV5PuxBJhcZmHEPPsA0FGl9p86qkL8ZALsX3dWoPs4FCqTMNSTig
XQGZDAknPVpAHGlJ8JeMIhxr2qFd7vqCVxy/ofx7lEc1MQahRBVjjgvv5WVlFyhX
3LpYiCJjbbdES8i2GjIZ/6anh0kmvXsqMKQxdJITWGuvwHfkPICfjO2IRdGZlaoO
C+PpTn6P/5lwCODQe1h88PJ+T9y7ty7ndIWbvKZKtb4cUN4zdqugjelXFU5Wkv0j
nyct7MbKG8zmVmb69m07IKnbTvqETk6vBWa34ILQnhudPjaI6y0e9vbJbmVYDc48
pZNws+B59YvCfukYLiJHgBYMtpPPosutf+5OY1wK4fjX4ujYuLMMLBU+VrPc2bUw
a/MmBbW6DmAinjzPde41P4r1BRaz4tLpQhzgyZpz9Zj0QtgyqS4uZzOcvZj/dR/6
CtZfRYIsE6nWRlIptSL48k7t37ixgoOLzNvdYl1I2hr5/asTvOZ+tr2Ojeh3wDkz
kgIAVIya9p6EK3bwjWSTcjLEhVtVXiSY1poAOyHBlbRTcxagGbyX+uxGSUm+SJov
V/BPg3dQOzf873UHVNmwW214DyDHm5hW3kZvpx5dAMtuv7LTQ8Kh7w+TwuOsMMTM
77EZw8calFo4a2xeopNcyVEapJuU1aZAqcGOIZYkkSJVnLCYSP7K5rWhLJi/rZAY
Nb7AvpTkChfXG7cshiMPv6UfqQNG26zLVUs8rE0FLpZEoPoVsJlAkGfB1n71C0bz
SDZp7D67BcCU18Oc51FVRypj4SVhTAyN4/WJe25ruR78FpCM75JR0Py0Rkr0cdTC
q8iktyGVbfBQsVGTc1uDz0gHjT+AAULCvO4XXsnVWVs6s9w3bQKiUZiH6aYCAP/n
HsFdFTbcZE5XOP2ulo/oFhHwZXll7hmycvBBODluOFp+crOXpqRUIGLtLk+cSChR
LdJowgYTnHKi8+5EWAiuoqdDUP45natodgToiLhUhqGSjpQZZJi7BFRzc028WlC7
VER5RkWJJCmhcQ7qC6DkENVGAJJ0r9IUKujJokwYv4u9FWbHffy5WkSqsQhwMZg2
fUpjuhFMim9TVO9FIC9wXqUPv7sZNPCkTA24hqZBkQD9EGY5lAQIYAHHJC1/+S1r
qVhEeOYaq4ETW8e/sNchr2/KShyXvM3jPolWVUBfRJkuT/r9wnANFJqr6TsjKiGy
NbmjGTLO0u2EpL14hKQh09VV62PnX7hcyNzOBdpDSKs/RKNuo/zpidGyvP+nPglV
VofG7NJmxmfFf6CJ+tnKH5RmGOIpyicyVARj333el/tzecfQWfP2smg7GssApGKN
xl0XOM4yMvO6LqUbYPw1yOOosGXi3i1J+Oa6KnHHfrqA/uAt91Opo4AfQZIGKPcL
awis8uq0dMOaQ77NzDQ8UvcsXhVpUt21Blq7VAZt+vgxmKbFQuOCK6nNmwO/Ek+Z
8xC9cwf7QhX/Xoei1D5w5xWrPEw+vknPx695L52Oqoup9HAm6XxkAbqzFENVJshS
gn+nvAekt5sJeQLfF01U/xk29XFXEJ51SRMAgHW1Cmwe4GvfLib43ddVJAPVRBRE
gF9UFkJTNjCghclVePkIsYjYxjh2bEBR7RTVLQjsKCC/6x9kPOpizKpF42A8dCvB
quZdwZAgs86shNvqvrFuhvqGQCn/0TFc7JA6UIyVCUAk0avMIS1HQ1eAVeORT6DE
EMMrJShf7MHaNFdfMwSjULKCb0n6fZzMDOnRPYQXVAuYwrAP7NH6MWJ9YYraAfwv
KTzrAVEh0yE/ZR84FDDXMli/MX3PDIb5kCEgILluxp8=
`protect END_PROTECTED