-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
uiy/mcgVPJ0gtHQFj0mVC+lft7ZZi0Ye7BTFMgH3o7uQ3sPCqdwrEN/nHvN79Hao
vLIXurX5jkHaDuh5fXpcj1mP4X1bNSegnVVY5rshXGqJRf3fp+d7QaeklEFG0/5O
iPzp6ua7YtDlZHoFrFMYkF5AtcxbdOWsbbM/CGlcWn4hOSLpiZkI2w==
--pragma protect end_key_block
--pragma protect digest_block
frTWYtkfZ52mlUuoqHXx1fAgJPQ=
--pragma protect end_digest_block
--pragma protect data_block
sH5PmwgNK9PMVR78pq5DrbafjQvY+g5AvNwjVU3P7jn6sH0c0qTOaJePgvOi/uCV
uIrcyKn0foIvrbgu2P4WLLIRsqtz5m4iTP4pQOBOD76c4ryz96M0aIX4qB4e01zh
epuRwGTJ8dRu2AKZgAoauLAfSJ1P2RGqWPdGt4MpZ3aRD+DPNfPXUi7IorMfEJny
Bks+YLpqG9h5OosEpdmu+/mBf0De7s9osp0M/0ic1ct/m7SMRlt4UvVWMBOD0BPY
oZ+5HLAqaSVco+T2YQYO9Bcw+Uqd5gy9slkOLyKlvPPAHXlVWAzmo8/qKMRgsMAD
NmbO1qZjFKmutqLLf9ry1ZHRWZBqDpaxzi2HqqaDy2X8wMvDIPuZ0jsoqMzsQjG4
k7/iYHvu9TIjFmBumCdZ49r6fNRT+u2tqBTMv87jxB0rBOnQ8BVR8opDN9PTC705
0TTWHhLkyyToay+5uMVQeMSyVab6/3Hr61dyOjHDiIADhhCV48E82nTjCz89ZKtE
XeRo7oR4UnpbSDlYdHMZJM2tNgb9epAS7jYVHYNZX5gGNUEs+xmcD/aF45Zgr7W3
8E/wRE30SgttyHEh7gTdyC9NO2bLplbJTgWNmbKFzNJuBKWlW+KgHJAjfi2I+fXQ
erA2pjxyJeBjyts9AscgCj7veKHEytuSAr3AKB3YQJmdbzfJtQFiNAAXWXet3fC0
4n+0rK/RoXQiBtNs8dZi1Eba2rBjznMHaiW1cD6WR3w2pb2RZ5fUJJ+pPLMLewtv
WEFVDGHIubaF9Xzw1aONRMtE5gpUtwpz07PU7EQXHQX1x0E0uU44YcBIb4bZPxAl
ddHU0Bg/yvuB4Jwu/srAmASS7/5i8L1a4VGSzLbcyoTs2VbEtMUk5PajWcyIoniY
EHbD+l3V4zksM3E2bUIYyDqGwFbQ9R5bYvvneuN7WfjVsG3aGZRr/KkUtAHwDqX9
9RunViMieiZtgtT9YCMP/LKVpYqDPshI6/BUFwqLeeJXrhfnJ4jnnkxwCLtwXO5m
uH32swlmasUsIZgJBre91wlWQISj6jfgUqCUpwyWIEmNtdRVirnh0ghA+E1YkH16
fFJmq5JrPN4HSVShrJxa3Xb6/E0LbZVVMfpg+s2/HUGmC3xoSJfwYZXdZ14NcJkK
aygAVka5+MSlF2l8p3gyq7FEerrIRpQrtbwcHifOD+Pfb26REvs2tOfyWX8snTPL
m8jDvLyGrdNCWhkU1l9if3tX1GBMgqazMKUyogplnE6d/Srx3Hi6qBAIcWRM+yX+
qHQjKeKrpXbY0H8FzvJKd6DOCjTh6hMa5bKsFiV17Ehuf9RBOo0E0ZtXfxssNwXe
cE3qgo6Z2vBkkK78dtVrs17T31qABhIErNIoPdE3eDsWK7gSEw8OXRXR4otETIPQ
IcuOjFuE2uIyCDJh+/m8lEcqg83b7HzSswjIWb9weOur5F1FrkOREI9duJMi/Adx
l8+avNkVkh4bfkhDNzSmhZioq5N65yiqYRmm0QzjzLRbuOAYkqNgxGagTMmJ1/9/
OjySuAY1kfjRK7FErssLKrmXj88qoVu+SvJBsREOauHlUsCG2AfW7P2qW34x7EAv
OF221ULyemqfmw42A50CT/O6kAFXC3CDHdSEgNddhXANJNdFJPucslCEILmgJb07
2LaOoMe/7jHTr0H5u7Eq7TjrYLXZPTS5Bjl2rFE1sGn4uWX3hQvi0LIzHl5WzJp7
eofiuwjbpg/xhQWSv0j5TDwwkP4lfFQYJG23eESSH8NMWigmxB6nW0sJnU6Xvtk7
UI0yayfLjoRnuK7Iwkxw6RlwTLCg41atmhsPgG1WJ6XOE1LO21ADEaMmra3RbVaS
fkqjpkLtquCHsKTW/Tk5MHyKeCAI8Na/q90LcxmcNNSws3kHFFRIHS1v0sW4/JJi
g6MeHvjXneaW+Lkj0IJ0hzohryZOa0dJhSTtepTyuHOX+QshEjcCU+OOiIkMxg2+
4wpV2FQonLdIUJFbngZQBDk/aK1A715T6MlS0HSh392oBVeGYKhVjGQdlzDn2Dbr
GMcbIQFSu76hjKvigcpCFS3AYs31z4LltQPL516li2Mh6nHkzP/02uTkzt5GaBe6
iCOnuOTx7oBoCdDFse69ayRG3/glsvzdR+DtbuUmhdnEQ7DDsKCSK0mlmRj8vmKN
actgxV+/6S5zKMKs3ynEzRuTU0UKC6zWBKtbiCSwKTQYG6YkpIr0VHjVnsiOkYDb
nA5nuC4Ql73wF2pAeHcr7y7f+Eq7TtiqpPo0Tm64zu3TVPfEhtRJZzAObWnoivl2
PVBaBN1BVLDbafvzNwxCgoTeZp6lO6WAjanCtgorkeN9/hRqadRfHYPYAKcCmojZ
sCsK8/TdbX9gJ0KAD9yqXLKDQWBgbc0mrA3e+w/z8GFEJp4RnurMf+2CBu4CFx4c
L3YOFbGH66+SE1ptNy3NpR45WVC5a2HUmfn8XAFwUQD4pr82zrE0pQtG12ZJ0OWm
PCltKO2Rr2M3wABzq5nCM9f9pweJDj2K26s7X5W6qJC4qLyHXc2jfG3LDpXds7iv
Tss+Iri143sDGfG0E+yQklZG3gWZm+flEy7JbLJWkWsiswr7F9M+8ybI4jKyLEvy
ebVupiaHEHloqwMTH1cjvPUvfW+DCedi3Ek2xh9KxdMWbeFiKCGNZcF5LSdA8I0+
vKn5LUs6MUfozp/N3TENcjT/mA+2Lwlhl+WL8W650S/JNURK40kdzScpJZqGLoME
w0H7JSB2Pl7ue2/kI/7XuObvmWFCUz4gC8ZegBuGMxibP+JQn43zAVb4L2b5QLKS
bTbOkxI4cqUTPT9KoBHuZ4aFzIbFQ2KwMtnXPUOyDz7JGP9fffWC9t5NfQiZ283u
zvGLXoMOvY5Aem9nie/VewiyLyHcDVDcTqihYiteEthHK3RjwQlR6m6AUX35nwNr
gW6EFsOyJUO4Px7GohH615naPq0u4fDKpC0afkOchNzAjf968zw3GFO6Y4hPN5PF
i4d9hGm08KFFEO/JHSsCbX1gsUIlVf4CefJ4XcfQG0DeIfm39q3hJOZYr12gsSes
OzoHM5lUhjpaZCJ7iHDzjPDt22j4N3V2Dalhm0Sh5eAv6Hk4ALk9KTzn6bscqFmV
ekJGOiVVHoux1wUyYuZwZxt2rt5DeHC0IhBWLmAqxvkSMmOqcLjivMTr2mYI4N5K
Ivw/DlE5yZCuj601tjcUH9kozlw0pV3r/dq0jr84gd1efviDUpt8MEsYvHV+yvD2
BmhXGq7JMeGV8SPUbUpylBProwLsupIOgp6CvJK3xvZ0teHJDRX233JfPXIcG6I0
QvruYOhS4tixBaheAMoao4Vn3CXz/0h7ljJ1LVUGlhnsSoLGcEgtbv6vfwogt6/8
pDGUFry/bm/yWe4/bxabv5TNipohomzQZcyK3mUbiBIlu9uQNGBOxmwdYwupDBzf
Xxo0tR/mJKTwZIbjpw2EukO9BdGyrZmZGpF111RNJ5+oZwwiB1TBceTQ8qzhJzVD
tfyWA9ojJb52ytUHW88rw/oG+Nmxa1fQ+1+qUV58zZvqCK38Nnx8lolY2Rp62aYD
Ewxr5TDltyANcgUrcihpdv3cRWeK6dE/J+6DMF2AqhXsjElw14Bd3hhwfdDyR0gN
K0faq7L8D4B7uj37O59bA4Cl14vPyf32WDVBIWb+E/o9KFojSGL/7wnuxboDeM5G
fiJPYZyEiX7tQ9JnI8UnjqL+fMqAj9yygbEZjoi0ysN3T40DBslcZiuIFNcT5STj
Bty1ekBL8I3nlo5h9B3JaLN1NvtBbzdjGenBKRDNR/W6khhEm+abczUviRq/BeCU
IznXs4HasxCHqoG7RN/EDgskSEtBwFRyS1yu8a5mQEXgCxbYtANvU7F3L6tjDScu
65GI/4Qa6S10OIPsKnF7HdRuebls9SGOpGdII7xpLMU8/Sruymuokkn3ghb5UQqc
SOC5EfDUHf9Rpey0+a0gBCzCksRqpfIDDomrqCLRbFRBXhFfbzcst8JIO969P1sw
ugpl+whLKkel+FS2Ej9fwvuvCvLKrB6mXhOALXz98lT8nhgPeqp/vO6vUOnqRTSl
OXmW1vAhr+CLNcLbzL/GhPiQjjDxJUYfgTVkVpkBSIrFDFJFGnJrvXk0pEvgOroq
48WSrKC5CCHn4GmSfYR837WVhkzWaT9hK1QjJRy0k0ogJ24JZT4BpDIbfYd5oiAO
5iSck3jE4nvgZ0idrdjtbhp4yGGmY+m5XZwI9sL/n9vaR7ne93NR0ZVf044KiJcF
wF+WIn+0bAxWtBpD4Vu76SFC4sH4qbGElcBnYc7I6rCAhpIQvNsxojktkKcMge/Y
qdbWpnts3yrDBQ5iVTa8y7xs7rLmEcqxrYNjorZ7PUiiWMQPyTqapW5ipEneMzw0
ZMBkkAAt6L9+dD26tOmQoWV0jFgDGbJaveDnyhikBgMKdlnGwsIPX450F+isC32d
TABNB+T/SM5bVB0rglCSCEAGfWtA9najq65JI4odqJAUPzBTvysySrdr2vuY49hi
suWx7AfkTlIYTsq0cIkWyA+sKvhcL0SBwVHP3wpFhdGGapnScu+O5+67Sm/4waJ5
Mz/7Va4nllootVT/e0y5TQWBpiKUxSecZCds3y6HcTO3xReh3nNlj24cYBB0svkL
UowQdRJTElHuOY/Gi6THWu7T0bGj4rHlMcEOBb9h8afLoRbQzn7+26/j50+feWq7
uMtaJKjFiWQSFAzvzheRe6OVAw6pn54Kl6QJcnMVfkPIHGm4TiwkHPJcogG/e9jV
CNVP6EcoXAaJfnmmuSl+SuRVRxWCUJzddJRiiRzb6y+oI2ibRJAsz0mivNAxYZdb
uSHQ5Vx6sjMDq8TagXG/L0ysAtqKYI1woSe/GGQ3LYI+VZS+677tzzvp9QUZ/5Rc
yuA+c/0Abx/L65PukuInjVKuV3xYX7UDYJygyLXXUz93vNdZOYL85D9OepmubLNS
w18CD+pPVGbpkXDueweNJXglAdeb08WYPz85GlsnWcAqjFSN8M8L8lwYOYmybXxp
m8feEtetDZtWd4b5MpLkj9TGkYeInRFJo5N+pzaZ3Po=
--pragma protect end_data_block
--pragma protect digest_block
Whjm4njCGBeikfS4ke9Ppx0nHxw=
--pragma protect end_digest_block
--pragma protect end_protected
