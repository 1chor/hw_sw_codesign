-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
PljbCNLwQ32g7q8tvA5oHCN8Yn9gjQoujqQe71YbFdmQ9mnufGuZhT0MPTxdPooz
neOE5qpskXhcLtTT9e0halDO4iIqJCKFw4T5VqCKUM1Dwk8kj/8Qv8TOOs42A1CM
7bkd6o/p/zT+mBSgyB4Yz439mrI7q9xa2SX5bgqD8rQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 34470)

`protect DATA_BLOCK
F+XRu5LlO5o2ebOPs1Z46ShM75CA6/6zUedv5zetl8eMOsNw9cRMDvfbrLHIS+TK
4CmNBXLpu/jtxrMXWLr2fdAWDEg9rbArUgVcCh8nDJbx/GuLYfGn4weN1lKtDRV/
VcbdhJm8RB+gfEBJsncevvT5tKn31YHoI4qhlf8IlhU7JBnr4ivo0buHa08iL8qD
u0z69kDyEoHCBWdJgG6Oy6UNTnQhTdPd5tcJVADB+8y3OUcV7nGbTYDN8X58bIUI
5XkI9Rjx/tdGeUMZl4I45ut5UJVd7DplLcDWJDWI5BHq6a+FHmKobJhhU73Movap
bI8P0kQMt+hO8tOEgKo7lHGfTgROm5Zq9t8+pIbUp3DemrnGpQzPWzswMQpSv1Mq
QBd8smCFzDmBU/3570dZDe+M8v3fpw3/uZ2zLdT/932/S3helnuBUUDXH029AilU
vCWN+ZmFdmfwRIR5iiMBCGu8LDnH59V67+LK3t00kJSvZ0Pvq3G1m/kLFfQLAtwR
ZrSmcBai3nRRHy1OSGQNYSFg4xlzkhmg70loAswHb4/dFYqxyY6jZ+deVtYAWTaH
XaNPF3wYa3QxeYm7VLqven123RlLxQO3qNrBi8k+G85UkJ1mXXFTGIHXPB5ird/D
b/rx79vkZ0BVRj5lRQVXoJORPlY397xpZATQK49T6IB6wdgOTSbdiLNBP8ZAfohJ
FAqKvXsfy7SAglYLCaZenijybppycQX2QKMuit+QUO/XFskK2+txH7s/y4cLsGrC
KpqKCZnW2vpxmMN89Jma/SaGaLjpjL840wzoG4mQt0SEl7FQpk65+qyOaH3+JBf3
rojwSDJUKiQZOa6kFijdvqo+lQgrlvPh71ULLnV6/e4dwXkNoqbyujFPf++rwT45
LIIGqIg/qLAp+67d1Y9Y0Qrt1jJsu3oAdeWjCfOC5UkuIOsHZXTXox/PMhPXIFOJ
pMp5cOrxmkUOzHDXzqW9RpNUH0iPfdAMTngcb9qpRBWbvJrAauJ+WRvwJrAAsMQj
5ONqY7OoZYKnixyVUtuENOIB4UCmASRoszWK3DZrWDhlIM83nNhQg0+IE6K0mniW
Ia1EIA8H3qi/d1vl2XkA+3eTxxs8eGr9twKDPOqEm9Vma7D7iDXoIpCkmwiiLvWh
LPnk1LvGt4yjphF3FZKrE5AT0VpfmliOIHzZ5WAeYziKgFo8mNwyHdqJcSHDIK3l
NWfkXJ1BXakf9rzlXucdbiy635oPJft4oGrzybwT/NdSbYjRv2vEhmXDdeZjMNC1
fhv2V3VRMDfyNbr6xTnq5G+v8adq7U0jUPzZylEYe5SCzhAcBPq17dRq3p8r1pjG
8g4barhv4F9sxAXhdoOfHgs4NFVEhZhNneNq/zgs4HYcRvIK5ChNvnh3HvQRmRpK
sewFYhKvL8m4zA4SCVGJzRt9U1N+Jv81Wngp1HtvNFdQg2+Mij8+mpTatiN59Jha
b+344TOTw2ejn9kxtNZ+5YrjmthAZjeVf+C52cqEnjypqanSB1BHFPWgM+oX9dPM
kgQZ0yAn3I3qNRwRkoByWwGQUJNnb2nIjMc3+ahB/jd7XyAV8DlssDiIv7kpgRiu
Do7Yl3aHoL1yUl8cJirqIStgwcBcwagYB8ySOhoSFqj0dh5rZWDFmdhccySsVRp3
XQWlhZ76LFAqXtos36WatTiFtA2jn+H3dz1q0LRNkcIMQqj4W78tES+jImMU/knN
m77j2zLAi51Ix70IZcHyPYOUwkcYi+rWkard7Z0+WLqNRdGdeCY/pACqlCBFSZ1Y
LH5NXLYVuZwDAmVxs1GtgrZyftDMwndSGXnGuccXD6LubsFZPPbnvM7UK5r8S49h
PCOLGeHy6frbrMg+It/L9lJYQsBlV0ycFG1VEYSQtDhflUPPogbXN2l/KihCCRXg
4mCR7wvsT18RHOmg+/rF+a26XZFDKmz9f2zcGR5VwsBVy5P/D4fVeSHa/+c84fk9
KvHGV7TEbeLWlR0OO+Ihp3wsJ4m5mDZxDna/VQEjBHsXKEiyQVJMiEYuHg7UDazA
9e1v1cPwPDccio/stbNBxruKlFc+KEjcwq04w6qvGC6mVq38WNMNz8pdzp0FvbXQ
ZzKW9khPomBhK63W3OuzF+Wk6pVNBnEik1c5vKaovLsmVYu+dBdcIGgRn2QMJg89
KZD98tbPv+pUMlRasPbcPqUDQj8pydyHE5agHopwUp/KQKS8DxBHNaTzmLL6iAtR
W9kPRIn8u/qT0cXrSvV4Os89n5ruN1i2SsM7UMCXonGnU7ugvXWSNgE9mYVYW1Fo
TF1m1EeCYLHkBYuCytIw3XTHSUenK6pIn6kWWjlgWVGFqhpNowAuxzT1dfrw4xJG
zuTYBFIRaBi2R7eThWDB17xHkyYt4XvUZ8QYoda3tk1FwABClhU0Yze60LPmN4xo
t13MxGjBHMaSnyVadObxLcgHFR6kQF9L7LRvQLLx2yjsp3Fgmfr0Sd36N5N1y5qm
mhtrb7ZVlD9fl54eGxHyAo8nuS14Vyw46teNHpG/fHV29WG8svyaZ9pans4n38Ma
Fbwhie97b0y51JQXgCke26FrcKNurwdDT8yiWXO3nI4iDoxzlZXFWajsUCtEGtKz
NJsMg2boF02a5d6Lle+21VS8MGeHaGngE+7zT8RTXih/qxWeYP1nyzAop8suS02n
ZImgl/I2eKX5LRWJ+xXs4UYp50gU7jniJjrU1IoWXCvi8H1And+oryRj/UfTQNmQ
6CZ+kVGETcBUs5G7oBfRrNufZnL0w0USJI+3Q6QAY3d2WEqjlX36SCnWXXw5DkMv
zydp1AQyUPzhn7UbRQag+t/ivjoCQFLHlGJFpmqdmttDBcz0W+iQAN7zjhezslEd
qRnYr9T7ITGY8lEEwXcUmCSXB+92Q8rjWUTPe8rEriW/41LaXkBS761ffltPPXr9
dYhpASWe6PqEwvr7thHqaeOKbGnDtywEaBZrXIceZJ319I3SUHX6Ds7aS0GSozNq
1/C3KqnY2PG02m2h6OT1CV6ZOMwyJdfN2klsYzQdu0AgzJvk4SacGPkCJ/RmZXCx
4VG1smtN9AtRKoAxpnj3KhL3jrPsc1KYVIR6wZ4YCl8elpSBkKmcC3alcbzaQaBq
KQCWwVqa+EGW7JGZVMrrCvrgtTazZmBFy/Wde1QJzsjRij9CZ+B2u2AlBCBDsSzf
q9kfvh9d8QTlUHUQl72F0F2iFFNLm/MLqtlf47jXP3I+viQAcugOx4M5vaUX6rgI
SQwmCxK9Am6iuMDRf3YMSUA23kiYSsfC6p83Zvt+ISOOPDgsUPFbWpQ2rFekiXiw
GWeIwt+HHm7yQ2cKcF5pVyqfGD/5E4EQ6Cq6GLGDtqBYjVnIVJRILxZOCVwYNnwB
MmLzS+ZdT7fxGDL+7xt5qQ1aUv/wza7wTte+9Il2GNu87B/EG6oW/9ikbP1rE7jT
E/Uu+W5gKTjOouqEir/FKUOk0BJQAe5GCprKtK8sHzNcFUZ9KkIsfSSyfEnlUZDM
L8wcAteH6hS9XLWLKVKaoJpA7gQgSQprTCg5uRYvOtVo5TAj1ccqj4btK++vo1EM
9KhcQYcgf6oRtqYF6IkRiskoQkWgW0N8sXyBn33MPSblfySF0PK9s6hVWySqnD2y
17gXXkepdI9R+W3NTB2BCeIAvt9kQ+Q7Be3855OP8pc0wRMGuSvwTX4/rRB6ndZY
YJpng30/YXzKc4tCKgTQtmXg/eZMsRCxg/PXSbo7RhBVz3UE+Rt4FFj3i051mRdH
dUlvWwHrBWIXBY7J6jUyHjTSLixXMeRZ1wYNDTxN1jfWCuaaPx/ffTUveFJ8Z+ur
vFbXimnfD0weKlwbq9NvZsOcwIH6eYFuz2SpkfQl+XZV7m4nU/zovIoQiud2yD6w
oZcDN42GqEbZ2FUZf44jhrAyX1rJeBNLEAwyLUoEUpIpduhpBJDbaWyEP0AETLof
Sw4DmnVpFAG95flqwM/RB5Bmz61AoPcen9R1tlTDP0xjeWoNSsK+yIMyzEwr9ye1
1jU7xetKJs7So2A1yqQgx9ia/g9HC5CwX1tN2A/acv4FriSOWM3KiH8LJBLIWYo/
Bq67i7tM7Zzqg1NFIsFNqWCZlK+SuKbwExKcoYsTIi4mSMiQTJQyKF+qE4+0vvLO
+x68S0Awj1AC/Ks79PCVzPMJPUz5ZjMo1VZLk3S7F5+Rg20BDAY/5bOzO81uWt8w
LjhTsUZmN1ZlF0ghYI1qTWkxLC5Oag30l8E1afkNlVYZKanQdYJHQEidpqtC+UbX
miIQyax5bEo79jf9A2xsOaj2AIdavv0wtZio7/1dvtD/0L4e/h48LwiMJW/szfDO
P6/DX0LNSUTSYmKYNqpeo2xhfDP/nNseNHoq4Dtkb9wxUkstz2sU20OgXgmIumoT
GLajasy2q2+yZmNe+7oN1vLOvpglKARkl3Tr9S5WRKVdBEQTZSuwdQNl45Ygs9pQ
I1tR0I90L8/svH+1PgMgFVCltzvNWLXvFleLGaSjYYHMvWrP2BpHyu1Gbis2nCwT
ByUU/eFiP79Q9UiRad2MIvkD17qekeL1PSk9zCpmnGPu6qItXEqor3zKwgOrf5or
PHQFmibElbQ99oxotBNU6KpgofwhQuzeDvwRRFAFxAXtzIyYTg/clQzEZqMrFcAk
OpAF2LOEqijWO9mE81l7UidPWnW595ueZEV1jwyCFBN2X5oJ41rcGYheBaN/rhxZ
GI0zuuqQ/B7RNuVoul770eAeBtiHcVJqiWJeejj5kpfzU9UJL06ftKzG/vaAS9vw
+I2WJb2elw4674TdkLQ53MUFwYbdz/4ZyVQSPNsPZQMQ4mUxkIhXDvg/zOwzg5O+
KTOOeRGWnkH7+vtuWBlTfH8RLwN4D6WeHHc0CXM/3j4gqEiRKpzzsV5pi/qQe5g9
ChtvQTCAS4hBpcbanMjeTYGY5XJfrt2jw9q0wwow+u0q3hAYyPR0EuiVKnLAAy9W
t+wzYHTWD5EhJrLqVMo/a9LFSLF776H2vCYKRsidjo2nsojA/qgrdt33xGhyjw+0
4KqkjT2Ld5TFjUL21AldEi6YB+YS73hG96AjLsrC0fSIG0xh6s+ULldcOthl2X6A
MoYkuFp8kgdT626ziBUGWo2JrojXCgBlf3htB1RiMZO+/Oy6GF8wPZrWQxIr51go
gIDKJwFGAbxyGB1j1jtRfYSz5ie29GA7XHciD+u50LGPhegBQw1SaHleJCjwnUoo
6C+zONuO2V3L2VLfwePKJnml3m1LjghNP2eiLGh9DpBegOhI2gwPK35tyeF3ZwOo
lmm18rQZNBTUQCz1GLycFtjltunrA1u59AILjbsACMy0QQ3nVwNFNAchH/6WgTbj
G++aiE7HOJslpBSGvUjJZUg3wNUuz/qa3L5QBFB99l4mJOrfG1AQhoHZiGh2IHZh
7T4zkIaVnKTksTgcQKbyKMtcx8Ibs2rVF6eRTp5dS9YVum0IjdNwdQ33IBqEM0nC
W6ij0Tt3nZWhx8Hmsu+G469eIopiQCw5d49vt0I3NBxerWWxA4NFSYceyLmfv/9c
Atj3we6+u2F6u4/RJ+7a4SFhw4nOyrkhrIk70h7Id59oB2eEdWHZ9bTT0Eg9EtW4
8jnyyq7UncDCDd4As76PcbOQ3q2bP0yTuSJ76PS/lc3wJYjELeaV/ACl79kvC95e
AF76YEZUTwMHEF6fLCGVfZn4E+u7oVCy1dsqG+TBoLcQcVimPSqRUgcG41K+PmIb
9bT91wAYSdgv0dI8ECA1CR9Io4uu1JgpYtQ6oZI7wtAXOXJGtz7KYBnZlWyTn8iS
jIEV9fTarRgLBWYB5h1kCQUGV+MH8eOefMixE+D2RS5AbRdYWdhq5/2xlKwNoRvS
sIQaYgRDjt9IIiupeTbIzsky7aDO9hMODVzDUBg2goZ0saOEVVE7g9khLcQwnvhT
C74JbrfqkVtiWXuqDQC0htDAoVYsLVWf7HoXOEBCu1TXzuWY2rHbufyHp+/KryQL
DVRqS1/abWqKUmPXhdcjUSgsSC5ZdQX6INRsgMql7vtB2LF+6rBFb2Va2fnkQkMu
l7P4NDdsI1VyB3vdkhZ1TwgQYMPh0SavMH+DMTzQEdeCIInLkNe3wPXbWaz8aRaF
SVAoTbvDjpuYBnEtj27Yd/lUtcAG1Gt5bQKWyC2iWZjDwgP24gL1kTJJjB2ChClp
aqFSDJCyi9R0Fzz+cJKWczl4D++xtynxxBzwSxyCK6qpzAch4OTgDpiKgQySLaEb
je2a/4E4m7hO63F53JsZhvtzSpw05Gpep3XBsPKZrB5A21nrxle6dBbL+Yp9Pjhd
tzvEWMUL0N/l1shhQjGae65/y7p++sH0NMvzjw+0xBqwKSRAP34ZYSCgsEwGgOBo
VBrzhTfPdF1i7T7JJq+Dx1fT/6I4g/EfmIk7XCM/to/nC6tCnPuDTdfON+n17Qi3
ODwhjfa41b+MwB9Q69ZeVGV9z/oCC/9DHJ9GO2GrT2aAJyThAq1Y8EObkTZ+pPby
eN9UqXwPf/YnnTaoU3QolOqlJLeLdZnMSMRyGgDjYsk7v6PG4zipMIevYprxphO6
9hswVaBqdKNv+AFR8pBdJxwMfKl/d9Tvbv6ErcTs3frlS6FX0yrDi1KYC1595w3r
OxqH3y+2Es3QhegsesQ/wsj7JAMNLb8ejOhVcCGD1nbgp/kXdY4g8IX7bWzvwV6+
hFGAIQAEHzVSG+lXwk7VOjAE/rImDNRQ9ENbSKvfE13ti9sr0N6TsI/YpOAy+ut4
9YjFHowuqGPD10E8Wz3VN65GYuCqZOCtIkENoiUEi+8Ikxt2Cq064Ht8V/KwY4NS
8Q9SAAE4hV/8tWPDeoqGr2ZTmaq3vfLAJ5Y4qBsyAvesZZgW9j69TxGOnOo5gTu3
7MHYVyf/Nr2eUDPr+nDez/19VBGmls7qQFhqvc2t/i9pFqXMZxKe2fu0OSeZSQ0t
DUg384H4h/Wnlt38AsvZYiSJ++so82PXGS9rIBZjFn1LkiU1uuKOs//9F3NRk5Sl
SSQRoVFQGNGcSMj8rUXQ4riQHI9YNq0Zr67zl5sDzTssJIkeODiaNVEhNkBuINZi
iruL7cTpQxli7i5uRxiN1n2t+vqkcGI5gKoZhT/b1L0bm6Ma5ssUUK0+MM88+uuJ
nTOeUV7LTwJFhldy/jXsmviewph7/EHyxwaqFa05XrxPK7qMc60I3g6Hr6K74WWy
yECpn53lI5KoBhBb4etLZ2qM4hUKdMmxbJX7DItqdk25RM/AskzKFgi0nDYZcPSp
YxzPDjDVurKhapivQINt5eXFRyNG6v310ox9RcFmz4xjCnX7GR2gW+GdNZ0S3ei4
t2bdHPtMfyS5Qgkx85SVrmTXf2FZw4iWCjtJhjZTDbEzcmUisOvs1sZ7EIvYOdD8
IqPUuQ5dZKVJaPx1cJc5cdykCoii9fBWaHdn9RUbEQRAPozoVWWgeLw1TbZrHOFu
uVenxnA/RAPvkmXloQRawKNsCw7hENlIBRN87TuH3YrdgsIB23aMupr01gT3FMiU
ka3t3dAzNyNjpbhzcydDjmN0ZOWGoJKjYXvAHu12imeRRhy4LBx/sXwuWYLUWT78
DtkWrUOfEhHqAbmQote5lU1QhodZjtrlBJeSekSOR5gbyAjwThm8kFg4Axvckdqm
1fzrMZgEmTMFchxzR6Io9TYCrVfdUwggIyTfFC+mbQYxfDvzYfrPRLW1/98bewkr
ID5MIwVt/TR5wvlOwdz7N+hSgEdR9EJKfmGKut7RlESItamwjjoE+XhwcymiCaVF
LFk7MfLZx5bKSxPCX6dK2Q8NfKvolCqbl1s/n3q9RHgQHCFUkds6S7mb/8jzQs6q
P5QZIQzyQ0Fo3AeGKnQ4eMxNjuAUiQ4sudeQqFULxY9RvEiH1uE1L+SLzUaV3C7e
c1JoxQpmXRW4vlmil+5rcHTClbKATC+nApg3fnZcqogc2xQBNLR7gutQUNdgWvnN
mzGjjkWrCgDd+F0vsmZ0aOWaZaAb1bLag27L6zF6/AOhbd8SybewC3ZWXyrxZtda
edn/Pca6i7cQ16lc4ddJYMDBq0WJUUWdcMnf8UuDofIHeyfA6u1xWKJnDgZOuzqG
cRa11Ztz9Nh/UOHHoMGNWcS49QVr9xisfgpsfscTTyWjTf3NX3l8C1VrJAzff8tQ
PTQ5Qyywi2NwKxmr9O69J4xjP7qWHHGM3IDQF3ikFmrJd/Lra9VIOKHLsNzmXa2Q
3kSjn5ogC3FdC+GFX+/X4yqDnJslJ00avBkmVuv6w0CPE0Jh0G9ELeD0jH7DUMFU
DWqMxwQDbFxOyoInkuQ75PCmmi6STTKSF+WLejsVBXc5VBl19lvRqQ6i8DN/0Ogw
SoC+Z6BcwFmsESbXRFLU6WEGwxgV5bPUW+quKJEMP6qgONcXQ7/t5jPCzdzy+Hl+
782BnseGBhKDMYl1rSkUi3WMxB6eHsBoec/DWOHfidNsgN9AXSIYg3FlB2ysnh5r
luz1nU7N+Xs/M5zwhdA7rsNu9MlSGXkdT5sUS8BPSoxAvYdlHawXqrvuCqyJnQ/A
eVfh2mxowRH92bi3nOXQ5YNEU/rXO618c471mxBYqd6Q6DcPjONB8biSSJmwFeKG
raIzdEE1+BSVNqDnPz2EPSsTRM5REjBwJhbb3z0EJgBHt28qkstJyN/tdDk+iwWx
88RVVEXq3kt9dWsBw4TIl0D6ePCN0ADhX+o9+/o8cMmfBaJ37R5ylsAyqPNvS0yv
Fx4W+JhMEwHsWivF2ab0QSn/ma6nrj/7nFAAeg8guEf1yrx8+A0TpDnT3KEv6GpV
hROIUxIEM4JpxcZ17NDpwip+q/gy9CQ/S105STykLmYMGkXdZLCZEieS5zIsRh0z
wf5KJi+hXRv114oz5qgp94Vqq0vjOE01Z0gYT9LYjbR2TtG2PxiNdTH7+4Vj0PmZ
LE+d55YVejPQPDoGj35xq+SsJEg3vH4zBPL5qAaPnwl6Cwacv2JPOPSursPlg7SS
lBQCT1ZrECU5suMh6eJZGX09JifsbE9o2UpxXFlWj3ZMRWZ9Q0NV/Fu93taObtQx
kucPXGMPtkLuvaJEGncx7YkvatvK7EmJZtTT2C60ByiA8Il40pRKo4aGN7KvytYA
rZPAZ6t6lf6QiuDy0lr1B4Sp/reiaaWj+JyCT9EuOxRDHAwC6H6KmBXLLSE6f5cZ
+QGHFmb7x2hhNFbYLhatOrpDBbGE5b6LDqdGasDbKsXfUPWzz8sW+6oP7Qsw3aXt
0EPLT12wRoXYIBSzCvyvjT6wuNywaDG+tylNRBlHTcDaPDkLW3iBEw7UL3ySIg0x
Otc5BoY5mmGN7XjaDEyBmM+UM6A3Lc35aCBsKecgLEADNQzNrywnTMSUcqBO4WdO
mHo048qYSAKtldZK60cMqPYw1kFKPdQrgPtkv/w/naDAUiFmvGwIHgEYhAYrEQMx
H0TgiwOQrMBu/ZrwB0PDi7iWbPZMxM3Ozc1cpNFKLIPSyPzAzgrjZmLTpsxdY2vn
RZ4oiIhajPlbhKmjppw3s25TAEnE2Q+eSZqre+e9+dMhttcT43y4MqExmKoB9P6R
/+JbRtaJAxM1cyGRPWyVAqBPXbGOeNU9jCqzHnaxqi4ikI0z7cEgI9GcdS6fsb5s
db2y4+7p7w7tOqICJ+vPlbLD8TayQk6fT/6s5qrXZAlnqI0CRr3RI/dX42dxiMdz
URNP9UeQvWNnh7yRsohYHRwT8T8P6/x0+tKppBu7srdac/1r/oGjpsQxluNxBLqJ
NODy2s90R/VG8uDYWhT6tKjS6uw3dyQdxfBXvxdwtJjLvOeexV5I06UMssaiq4sn
Y/Gi9JlZ/2fwhc6OgBwhWd+lrRhCft8dibsQ6LeMHl4QLhiedBomxaMOK3RXt/CP
/MvRnlLbFTGBSkpgd91KQBqCB2YiNkHXnqfVhEpJkH4VWoxKlXEr6TeLihYVmAyf
TbaQwuMpTyKuby3CbuA2kM8c7vb/asPPZv7n4qfEupmDeliL+DSJ/c48Vs0zudaz
sNd3Ii+ix3RiqTOQD56ie5bpIQr095eZQaoEdbSmEAHMSGxX1qTBpjznyD5UWWS2
aYAtc6BuZJ2Uzjr1gGXCPvvRLa8dmHYp8d1NpQQgOw6TDHgkX9SWW7VdVRRjsvmq
nIYOTaGIEnk1BloQ4n1fFoaaeetHFiUw4Uzs8np3Tq/5Pw8inDeSGqzPz4uCmGkr
lZCnKnBgM+AMY3BxZbwOyoKQN//xxJFk8+h7waQtafjb4aIx2+nWlPKmFrnqP0nV
hbpBahsDpn8UzMx3LX+CklsIsHb9+6jT6NUTabuLUKhJDrargv8XkZfQqfm1I/9c
pA8TeYVXytONwA0akPl3t2K6xN3mecaNM5piIwrZkg3WjybCkbI5XVGJreVXb/ri
upDj7TAdKg7nkWg0DOXf/jxZSDr4oHsAN1jBUYgHU9JR6hMbtMcrjtBbFQILT2x+
sGBq92cpmbeY8L/56U4bF07E2Yg3hxTOwBPU2z/EzcG55UiPNob1tP9tHThAhY8h
IaMhaiiTeYDmDzRpmo6xNIALmEZryNNovyPmbu3Q7Fr6rK7MLWN9YIhceJScI3g2
TaoJJETE4rr3x2rsOc97lWR1VscfvklU0KDiQlg/2tikFSBtR6MtK1mrsyHDvySJ
WzIolayCap1ye7Hg5KpAinUiOtoDyNqNkaiMYestAwJ5wr77sfmiO8t1pBYcl2KE
wwiyo/0jH/UTCtA1JBvao7CgiQJtU95tJfkLyNCK7uTDYSqBIVV5GkOwmrUJQHbG
ehaLUURExhke2jsrBVKnOYKSG/cO+z3ywDX1660vR//BcfJtEDxzNOZ3jNc4ZSy1
fL6aSMrJWajRPpTFnS6vdOsV67JLjNi9q0Z8X8Z1EqhjacKJydq5TIzfdT2oIbxb
sOUwjfOizOX961ePqCtes7s+IHSuJSmS1pcIOH7vLmBCL5F40/ggDgU81UYN0wzN
U4zMEBZUA8bsG5Sl1gs7cb8/QkZEB+fQ7nGLAA6tHIqVmgnfci8od+mQ/FbKOYYV
5oCyQhCUWGrU8fKLq2ywgsogglobpYHZVxHfy3KZueNflgWxluxxSAwII1+OTAen
7Sh2X1o6m6h7Bl/RlFXhSghaQvHWGRZJmalGgeNLdqn1LLqxP/TtOnA5A0NmnXzY
wglYdvRv1RmgsovwK63uTK1tavIQCfoDSjoHCx/cz4CSVylQ8JUgaaIyt6lOP+Y8
82THxzaQb+83hTVcLVSRqaKTG9bGD5aFzMEdf/N4Tt50nQ9c+IK4s9kcyv6MUvOG
vTnTCg8EOAduDCzuuaPbCv99Nx49SbWzi3MO80FMAz0cdxgm5QLnc25w4BNWjuIX
HrnECE7Wh7dxtK+rg9NJB3WY26tpyE/shwS9n7QHZqmTEgKrFqqz2bO9WVfSIDew
gRCp1I9hkRQFcl6hOV1vzfvwhAFD8GoTmpRVAdY8uu64FW65kSFuia5/28sdL6bv
QEMurW0M2ilqjHyiJa06/f7hhZi5gQ+yZPCDY6k4kUn8pBdpfPqXZzmI7lH35mnR
oRpR1oQl2OqZWr8NaOOcubwLw6Mz59PofmbiUAlpL8PdUzITa7E0dNILyEss7fMl
SSDIMW4oZ3lyrvAFPyJH8Jj4OQUWCHIaj5mZ9Xep3u3G82OxQn650+Ue1G4kj59c
1mcvHmX+HEHimd7yJqFnlT+Goz4uOpoLRA8h+/njQ3w/DXCmhoqRyt4tcizPR+ze
v9Zrdttt1ZTCMDtR2+MDD8kXXWrUr1kjWHxGsHzQwtwTLg0yW1CkXq1W5NuYXP2K
VutbtPLXKala8pCg6Sy6F6C6RtEhAC9DPKCCYHUETKk0PKsUD6QNNdAA/6pYWxcG
kVO9ijN4crToN7fRr3hITqoG0Ii93ff6NoTG0pAt8GBL8OrtoGVIMSrzJ0RbxeNH
6/5SyZ4jEsZ6qUjmPLuHQdD3YPTl4QWTO/Pq661o3A+SDXJ8yH4c6iwYiFzJ3+e5
4Oe8ISp0HpvfzTBDrrY3nOuKb8+u8XD7SESi0nsG0zMeJRPZKeBgywZbOT4MSw+O
6OUeRzn4YXfnDX4z9fniaewqgPzsOAwZ6TzF9wm5ZZIKjZZRgePKhpyS+60375Cl
OwGf4NM8K12NC86pFOQLQLES8qdjiFev6QWx6OMwazS8XoDGgMpAoaypE1B3m0lI
loWfLowc4Bodz+AccDejE9S7UvPNVQ0S4eHq9SK2cqBAzdM08HReJp+fdB4zbyg2
M/JJA/czWAPoaRTVQSEeGXrO9FBkrfnNBJFiMK8ujYdojABn2YlKHnG4OlB2z8Ht
2yPdLCQXGFGSnA9lGHsSu5elVZgAyA3Pv5miMBW8x3HFKLJZBh2sznLj1l53qloW
4ADkG9dNp6OLSo+dvaeI/SMPU2XVycEmO8WF4TA9vNNPilbA9LgLRGeita9SH+lD
0/thYUtSCP4XQ3VRbJHmZVLdHMcxV4O/eEqDXCDmgPMOioAiNvsQ4lNquJxF8nL5
4lEI/zrWmdS7M37yjnHzQeweY++mrOMnrjKbYWyIqaqaCDgieho4zKgHNAwNCybC
04nwDTxKZR8OQbPYyK2/jjaDNBsQaJAritsUh22YjiGf47BvhHLBmgA/9myue4jF
hNRtUtvOvvUUm5b2mxJDzqGxKy/H8nvZJYEsQyCKpdDaH6thCXeZsaehXP+gajcV
6l/xgp5iKWdPXZXPOUKc/P6H9jSmYZdPKE5DkHEdShRSCz9BbYYHSbMOq5xXgPfg
bDxRITGXipvh7NOtr0R9gxE0k6HNje6bTwtjvJmit7MepksToZ4KezdfvQkU+tee
9d+zkmvEPlsGozy34KohIQ1DrEDClE5rCsSv/ihH38H2Z1u5GGJgmgRjPvpKxKPQ
MKe3m9ViuMIvgsiZs0pUp0FDwwO3YZ7XvTVYBRRxZ7e3MVt4gcTCZ5KoDD4ctrZk
ICE3M0Ozyc+iF7aA4HsDXnavfpGfT9hdJANjOrZGR6exGQo+ZbsWV75aoE7kURTP
tRGSS/shcupBijRmPfjLqbgeo1g8oL79YSsHKmWC92ynJPfu7KcFBh+NsxKvHmSf
/OnS3cfJw41Y4iy1KKsfasvrdz0AQYr1rG2cjMO1M9H7RRiclLG+LsXjtDyUIc9P
7bL3s9eb01OvyzvfN76/ghH42Bfua4Z/Zf2d1hyfy+MDCrCkV/VdnXcIkoaSJp0+
B8SAOKD8L6wlpHtK+6B8gq8lq2dK2v8xYpdedkAIxPZ+3ZlTg/CzA6vTnr1sOhZw
nyjzSkUUj4TBhHxsVC8S8yS2KlKlT1IcSi8ObcyIAXeWV2NZ8jPEe7vI3jAy7VeP
fd54Jos/txJtd15U4bwV11afmWHLqXMUq/gJ6lpRH0mRTx2Ie4NSrQWlzBsvq8OG
sMyGSV/9NiiZ6H7aYLQeW0aoowpjvA2F1RtF/WZqrhblT4kSYvdWOoCMIXWK6feo
jPyIeFSp55h+2TfM4CTnuT2nSqYnsQsRm2A3UNBo7v16BlzVOgWILP+DoE5K0iAP
0NbuVY5zXLaQRZHPzgonXiy/mTQ0GN2p0a5vwbXaior7eNQFIO53Uq7fPLrzBvy5
L2sVN/nMdsxkn2netnul6+UexfZGzjMhzjLCHa2N6Q0YLLR2nmmMrB2X432OejKO
wcQVfGM4Sya3xIL/LFzhuzkCvoGi2p5VQWJH3YSjjw7+Q+clrLuvZn9XAwmoj+9h
/kNqs/QfVi9skBzsPPLHAuxdb8+CsRGx93qLFvSEWDPNaSDVy4pre2m0NE6HuQMt
vFkIssoY9o+w/G0A46SB9mtmT0KKQndvgBYSZgIHSktXYCj4rsMqCrWJHQEyPeKc
/ysdDgO/NRwyKnRkIZDg4czZ0pCHM7XbuUvSNZC7JYS9h5mh5k9x8C/LiLrslOz9
8tOmf7VZpSfI7nWWeSlcyIIvfmrtdgcAOJVvu9hM8lieS8B2teDIY624WegG9b0y
fS1Y5cE5O/mFWBzCDtqC7p87zUlH0AF94Z9floz2NWjLw5agCClezXczHTDMwgCb
LsEm/bUNBC/SS6EPRBIebaSPJI/y/xYgGDMyH0wd5xBW6wrFdklFW2vnGSof2djK
uG/+tDeDS4v5gOJrYUsfFe4kAwqNOnxWvRh+U6Q14B0rpJP5NhXhQYuZ6GPtGgVn
IDQjifOTKnIhBSND3TyqkjdG1kXujCCcf2uZsd7/zOykKnpMjwiIgsu/u8pwHL/U
6K0pWNP3Q58lDBwCwufkpEB2IWe5lcf5x0bemWm5d4Y6ZeR4/6t8NrSy0DtjhLTy
BJwuzbrmeN20Hp/yrbhqDmvNGB5UhN6DPU4dkTN+lMf2iomuRzwccaNYqTDAkJRR
KcYpZzo+CBOTluQuaBc0try9SqZsf7CbaI+76EeDfKZrN48yvQs4XXQvSgWV4uiR
rUQps3zyuCQ2eplPpKuniUx1EsaOnxkpELE9CLLGEfXrhXiAc+yPVxMJI8ZYDIZ6
9Bv6jvQN3KISM6HEEbcQYQdcgQ2teT74yrr4zWj3RDuk7ScUcBpiVPOyZajjUuxQ
lOSQb5BUNEuZf2knvMkll2RPK5frQKDtrw5uNi1i/oGWJTbAIMS6a+uRi9ocwCg1
wL4xnQ+CH3Li/lSmApWMb7ROFoC2ylJ16guRZYy6JvnLfQVFWDGYPInbIWpPdJ1D
qGogUbKbXFpDPxJEmxtWKBbMiYiBtWr94HDhxxyY1orpYqySXoOCmIZ0ZHQY7Jel
c6UgDRrCIk6UPO452I2FpgmZZ2tLdnnLYuXnqwopWpfMucYzUD0q8uoNdcL0foT8
zZeuBZvax/oOHPcQ64z5fc+bF5lcsoMqOgW1IzUtvmtDQzmSQTsMlw7qTQR58HVg
jAfX6D8AdxKHcEeSp4sT2Fx3NPb3FuHT57jRSfzrNvwNr1aCHP+0v9SRz3865lTJ
fDFjtRIv7NqyLwCjqLD7KzEGe8rTjr8k8IUlGwnrjfuVG4ur6gAXXaKgcZEWQoEt
pVIi/yCqxNIMjkvNImaVouYBBTNrMYAJ9ZI+2Jtearo7r015MWuKbNAxNPvQyB60
/Q1CG7NsdmXgWSefgZay9hQofitguhGsnEuN8+K/8FIhy1vBUp1jjLJDGC24TxBG
srtwDWVDF0J+bfrURvbihBoTz+N9DB67/1A34ASjSI9fsUgaidt5mwuf9YtB0rOg
jTOhXiy6zkzH2gm6e3vyUxXOZ9qvLurlRlOrhG2jqEZOlah/69OT2KaU1hB0cwH+
hkcAokt2oup43igVctidpPnmNPo2YOJjTmqXslCobIOOunTn17SN6qotty44F046
MQkLdPzurVc6hL7IA1HzG6l7Ey0jij/rn0JHNmqNVD+O+TgDK5QTTDWSTbQV13g4
qzgxGbnpgEC0LJ9Gql8wOhfuXhlv12YIU22p8esUtNF4UThxZY9/pRITSgqJGsdB
aEOn1DffgKqG0o5EShSAa6yjdQ/54qIpEuOSERDgKrepsrKEW81ieFNj/r2GTRka
Uep/iYh2B+vevxjJp9pvYTUkE/iLz3rsAs9YH4AIhSWzuT4NG3+1nj8S0lQyJ2V5
RvIwykoh4X6PjocWf2JdxuZsyzOtDyngB/WIz1oo8GeYE8YdkWtXLlOTSFvBS6Co
nNKsqxJTdSORAZ2KoBb8EEtx+GbUDxZkXB8Zv2uuG5V8AefQoq92kmoRK4+LG3Z9
7WBSx7grjIt5G/rxputinkdYjrRjnFu54b638f2NBCbofIH32kI5qDVV9HUs0KW6
D1BKhNWTnODFAC14FZG2ZacljhXhkDHwmxoeAYw8zR5ZylrsR0UHBiKp4zBcEowB
nT6FP+iaH7at07fUkyYOmiy9EtMDiC7RbDK4eu4SykWAbpgAxXk2LQXigWyYfka3
S6l+R+7gM3Ilnh8KSEbM/X+f5c7CxmD4wQBzQXmE8PDbgFP5yNFYrhRcuhlJKRuH
1fu3/Y8PlRiuHxZY0NZ4pgcyxWFqcbxGOnh49/Eq3Q5ekM/pqcZaecIbWPIIsrjT
R3gOx3+fO/t1g0+Jj2wgwfUqv/d9KtQT6havzY/xRow/4ovADZqqsQyuVKfQRcYI
KjCKvPWD7kXe29jFll6I7BkLXc9WAtUqpvdDL+j4EDj1kPW8BMiorSboLlicqGiB
Aj1aFJQ6xNHBrzro2RiW7EM5gU0APXqIzwYbx+dkkVsuh6PWlKEAgk3zpkSzb1Us
PzX2PiENDTHE+yvmYrdumMuYlNFQD2YQaCbWDkVxvRKBP4BomD57Xs5N3GL7rP16
sHEA25f7pb1xo88imcjCp4F1uZ0GQ1S+W/pT2awId+j4YcgsIf1I9svjQWtvVLjX
eszTtPJVX3of0dGGEk/xcHJWCu0ZkmbyczNvTcq3zc9Xl9Jigz/atHBtiJo0peS9
+wmF/5+9SjqnSNqWo7Bvxhw8JjrICjjtgZdVX2kmva44QFG+dUeBbvhoxk3myemC
j+nMWmzM7zBXNxJ9XivYDuTjfhWYWeqghw41q/3l9HLXx9pwMw9uuYyDTjqk1nck
9VB7UFrmlmBbwX5vLV7hTHjIMeEt7LKsOicQBh2nru+OElQvoEqX8/3MMfMaOP9/
E3r7EnWZrClf9bnjxQC936F0CjXaBLmTTrsJCQLXSkSfRmY3jUfTPwKLSmvOB52T
dpxcXLClC1d69XMYsOsWgjkKz2V6mo3dCVAXJwbdoYBQsuBkwwPJGQ89LjjvBEQ8
/+TfE1cy1wPhR3rsmo7tzwhtHWzr9/KUiGWJAoKLiA6K1sV6AZsMmqTSSDKGJSYs
FAkHeUpnAn7AKzwxolPagxgcNyQJnK2rAkJci49y8iIuQ5+gx8E6UWpzBkNV1I7y
dVC89FViZWZL7tgh4EIDtbNJcIZ+MAlgNOFb+USIncf80TgQyRMfQALxqgd513Ab
Yxy3icLmVvI6QAX2LyQFczqGpOF/N5Qak2kt66xAt0MUsh3T4Vrwfdsmk2lN6dwy
gGW8zIsJDuYCGEPOV2FKYHMSFchT2XdgrdTzxZV7gbklioz1PMJSDrzs+Y5rq3i6
4mZ/lIyFS3q/1lqAz1Q4NdA65eg8PZuFs6Ih+v501ez9qtwwZXOJGscRtmqSON+N
bn6PRePP14K0aSAc1wQofT9NqYAKKa1ixBlGx268tRJmB8EfjmsRvg10rdYhKIB2
3oRI0Kx64zrOx7k9BMf1KYduecrW83ObXDk9ivayWRgp2a14j7/O37mLIF9Cd1d3
KCU0DJzRZZsgfdbSszwdd2n2V8LuQOCIpj6PwOW/FoZ7fMuFOd+ig7bv0A4Iw4KJ
4Cqjx2gqMcvkbktagQRXjRvNcdDdC6O1F8cJVc1kHRpA6nhI3vTg25YicG76f1LH
DkJ7qaIGJanq6niL0afncAGg3ZqpZWtt8sZME50Z7P13JAZ46kRZoI1SvxvbjU1i
6RzMKvTuuPovwbYmOJcNMFlughLExtv+UwtjvYnUTzBwOfPdaP3srX95Utj97oAe
xKktSjf1dxncmoDTzu1CEJIU032Gaekiqm8hX8mwozhM8Jpf8kRUAfNqgnQotumP
1WWxpZWUxWur/oI3b7C5sbtm7kNWw267rdxapdz55B++zZxfMVvkR9cW5F6px93C
D+amUfdXgnGYk84erXiOplVCzN5+mgOB4HZDVVQDSB83yl6T756+KbFlncnVyIRT
Q3eue4i18TfRYm1yHU/PKoNuIFi35e+sf9zBg4y5QWzap+HbdOJcA8pBR7/8JRTV
J58TkkFO7kC8POmm1VrNvjMnDUT6BfddBgKaPx7jR0I/oXkbrGpE6isZ1cPpFg8r
jK+dHTh8M04fujOcge7bCRASS5B5m+W8daSc8NFGkw33qoRKeHQnqZmG1w0GfvUl
XuRx8XzQ4h5GD4a/3B8aUfhSnTkhCdTIGxwdcwzTXhLe7x3wvdLBYZ77tXnD1bEk
vgiYswCWw5fLHP9tbIeKTizRwBKVYWdddlQWoLPTBEZ1Nz3BzjhYjBut9Sv1XwBc
n4dLn8vXn7bK/yKm9mvrsU9qswpYcqZmg/PqS/mkOUPLj6z6l8LDXNiYrt8OV+Qt
jDW4zYdmSiE5EZou8dQh1TVwFO/jWbk9CZEj0zogrJcykq+hSEzrpycbNeu2ZspQ
pz+qJf6rIiA85NzkISs9p2SE++/ksr5GT+C/j9XxN9B5no0TSqeFx1NMuxlKfMVM
n+GQZUmvlztbVN4mFj8QM3+HxzKH/hHJDJP0QCaxaDi/BTfKeU9YDo5VQkVXff/9
GHq6MPInkF8LRtB4P7COrUb6xQq/sFh2Mc/FKugoz103GFsbLriB6ykYWD49IUfk
RuHquDkzX6GCUdjMgteaBrJiWFKwOWgfUrp8L4P9ZohNtqgY7OpK9tXyPMDzEyYQ
kHGPtU7Sm++9A5cIYtJQo1+U6GKLlPxNLJMrDENqCJwbuJ8P3jI6DUEjFjBcsiLJ
S6VwAoDvFpKDsCNa0AH7iXwWuwxXDE9aR3+/qnGMFD4GFNo2JEiTRZneVTJhzhwB
Zg0A2upMyk/XSNVUo8ZjD16FHexMvi0aCoEGVT1o3hDjjHLo/0WrQM2q+kqyJsYO
y1mA4cUVCxXBNaNH9eF7ntVpGW/OC8u1owpTD4+VKxC6MpS5v36sHHaQMZ2puUEZ
el0w9ojOCGNNUDqsK9TXfGGa6vL/IRkueiXICosvELjF7hkvESLcr31hV9sTsiy4
DAEk6RZM1mKhV+dBFRIEdsTmsBBL/qJQK0HnFS5Or2zD59TQix7QxzMB1eKJZsSg
cPOHvOkpsCfgWqqxFUKi5Oa0tGLH9yDF1o8s4cJycAyzzVU4mN6pcJe05YENKS12
IZr/7Awu03OD6r0P3h+q59WxrfSz4YSErkqmB4m0hyejM1N/kjGUaEyqlx5WU58V
cPJQIAKOdVjeLJYDWXgI+qzvs3kqzFuzchWuF7tq/WIKDVoX5gLlR7kz466heKQ5
MJpRbBEFwzj2C0Lo3f70pemh1pGK6XzHE1hliCpeV9tfYfPGO0qPkIv6YLWUN55o
17mSie40jsMq8KraJZRty/bOCzLMUo2U1r8gCxVCen+1BndQxi+uimFFvs/VOgnG
HY4+CCKoPux/6YmeS//E2BGHRDlaToZR149R6dkCdiT/Gh8A8hQnlA7yME3MzEOY
33583iQUYY+AuSq3ftzxIawdUuq8OnXm4nFe5m75nKdN3ReYzPLH5J6MuVpQdiY4
hjudtUpB80xFK7N7DusYjfQUj2ZoxUQNu6CSl8QjVcNsbWfjTRK/34y7Ozxg1d5B
qMYuGjMDzjkNw88mPAa3sdEFyqzPMPmDCictMvgjZbM6obo5WBav1kvx3N1lHE4h
8P2liITuqezAti1BzVT3aaXzXfxfEONUAlUiAd24Z0fvSfPlwrj/JEzwrRsxMgja
dlQ/N9bn/dbADIxWdkWa3YakIvfc3rMONPTPFWExeHdFxrP2U8Cmszz0WabuvVno
fFQIg6xQoqtNVnEtJ+PSv3wDaeGmLCh6KX0EUucFViS2E2+8sMLljgYhmMyX/rZu
nsFva6Gln315XLxzweGxfNN/ninEoNefR3+lolvvry1KWzTyMGY7lv9/nqGAp17E
KurpzY6OqqS4q5WYnQSJLWQutu6ePlj4nE2er3hLlsd/K+oUBY0BW9saxCCyQKdm
wfi3We7JjWYEF5h/jdIRz5wScGAnC2f5p3Scl3MrxkKiqTtXKKkZWKiGSS6c6HlE
0YAqpS4KUiNgC0whaOWUFr+aiEtkXOquYUMJVgbhmeuKw1e5oC5X+PVppLItmsZe
m6P2lnHbccWyM/UKbU2Vu2w2tJTgizPTK6cnZwXQXn+bmcba9bOkcEsI85ziHvz/
yVuUdkMQoUNH+AXuoYQAollTrYf3d//R+uuw0k8eRM44iibqCGWVNvuHyZ7Xc0zo
4Ft5kIrnfWeXRaIhbMJMAmSuoLeRvjdSpRlh9sMDKXFqzSK0iajxGS02nqURSXqn
51WwR9vXNHCUWyMcJ+ssZ7B6d5RtGeVkSw4Rl6bxSv2dwOgZNaQ16jo1GkQ6IZY1
z08b++TsEUV9v0MOgjQC/WJkL2uzm/iUVmYi8CBsVQT6a7Atb0V5Hrgn7142/hTR
eh8aZtq6JceVPKLaM4v6ogz4xTFqCE3VnHxr/QTvmWP3QAJlszWVE2/b913oRO3q
S8BUdDofYAX61lXJRj6VA6/oy3ANfQPo99wfnhahEt4JBByxHJK2Jv3iW/GARnyV
H+n8ZRCH+dy2NR0gLe7RNDNGUH0sFTfIUuPDuEYYBy795srRFSLJGDz4OZUuzE4l
A+sTUnKrjg5mw9KN0nyGbEFy6X8x3N02zJ/SGd3/14NWgA95bU0koLQax/R8mLKE
bhgg3Oxq0LHotKTa/EQncGttW1A8Tcl6bPdP4Jcnb8bqERZw0JWadr4oNCWu8eiS
R17MLQYnzaba2qtsizSXDoPk+u/fA41zlz4fX8N+tyXPoSnNtg4664BmX5svpurL
a9ANWPNcqTS0RpF3he2q+FvXZHex8F2014bOuhTcncyTbn8vGjhEjU5iaJAOtlVB
d+hktB707TONsrgViQjv/wn75Wgjm/4Wrv4+X0ErrPBme/XIG2NonuRcLFw4LcFs
MHPO3exUXZpxQOyACT7mYMyZzMRsLTVjkj3gkC4Dg0lIpso+QCISvC2gUHMEbX2i
09RW3LhFm4YdKSDJuVi/cbfGljOBBYQpjXPcoc6FPRr4Q1JY1JWtQ6RoU9SQ+ajO
A0faAWtBsCYCMBR+xstRiT+PEcGbbC7t7Yb/4EAfpMo1jSiitqxuxynHXpgAasMO
zfLBiKbLoCKrleYaznTzsh9SgEcPLMkznP5YzIGxIN6lxqPtkobf9bGSZ1uTI8Aw
OulXHlpJ6gnhLFA4wLI/+u/6PO7Zy8Og0IFSFzeSWg9+xz37uCr2LRuizo5f/ByU
O6i05os+lu+dq7KDpSxcV5CStAhUn9m6WUyRIsNk9buZukKozaLAHF0Y5n9RcrR3
aF0YyJujhOyPrG4vQDhJXdiYDGktB+cXieJO4mjaaqRnAEjQXw9OPaccKaOAaIO/
sg520udEoXreX6dmeypiV8KttYxu2F0Wqa1CEaCic8f2S8cG1gnKbOSyCkBZR04d
jIrDmBSaKuIC2oEkv893KXNnBx5LBBaW5g5c7Hp7Y3faMvoF1M2iDl40KM0uKJ8o
XfO9uKvKtDOsSXiIcm9bNJFB7f7tmlLT5tPxdX8QMJiXKWzb58oKDUYyZ8n8pVog
ic8jcfFjbo/U5RtlFYAbV3X3lyFf/t4GuPEDeEEdnTQmCqi9yFu4WUq3LSvaJWKO
9/zVCgqEdnyBxr5L0dXwI8uKpvBSxbGIYMagBw754aB4P7ryx1+dwdw/o1bXphZH
VsGbJy3ksPGFsbpfiMkg9l76Rw98MZd9DmcW14bdlj1Zl3WVSfC2H9tTOTuhSe1C
6Mvuv2LeuM0zUye+3ZLCc4nsXsB5GSqFEGkZbdoMBegvDV8dg9z02W/BU+ZjTw6a
/BrHtAwZKpktco5l/cJHVApQe71z8s7qXJgXfNrIpkjD9NDIJo0+xwcTvVET0LF4
gOI2AiYWveFUOqD2L3Zef/vTJWzhwZ5ooBiMOwEzzD6BApokwqRh6uaSfQr/gOuZ
4AQnD/haltYSzqZazn/jdB2mU365YjojojeGk4BbZMCHJBbH/SsP7lq95gXcPfIV
028A9DpuVAJkyM1du68tAaBgURjDDwZvxAxU8x+wWYAAUGuOGkYO3cuD4siFMSrZ
KFo5B0X5vGKqlbF6HNN5ZNUW8baiOAP1VfXC87O4snItls7/sxq8GKuSIw/IrrF0
gBqFQTTtLnkjJro6tTkDO8XXtPRJScElq7stZJJ9NgDhpTSOLP3A7/2bd7P3ZtKs
YiI0f75MSMwvbTVVpZLiul00RlY/jwPPTO9sqW5KOhcF6ljw0ir+kjzuXEiJ0y35
MMkrxh4lH/ybTdmkDkwrJDF/E301flZhPzeq4K+zHhjLpqkrbkDZZEwWHy3PggzF
Qxkn3YmXejeWK8sKURK2WIwGxgDJ/nLTUT+NCRenOoMxFAuGUVAQwv39CmfKym2K
fcu9g4KDASy9ZD28IBMUvxjPOZWa1YHrmMpWvRjBLeqVTwYn0U+wIIeAxsDztxoa
M3L/NqAzPkdJrohbiu5BTdkDs2O633WobuFBGBwyebKfgQ+7Qo4LLwSTY9hK0yYJ
rSfAGgWZfLXy+8/0Yi8LXqxoFuDSRGWpmduALdToitX9HT9l0kgfvvsFlGGLUlzd
9coMgTZhGOEYHn3wGt5mbTiKgCWMtV3a1QKJ9ayqvhCKg5IDHNZkgVksuMYedRbc
AedPF7aCWUXepnmrb3I7CajXi0d76BOBCuoUHllnttR44r/hrHbbU0+ux+THqu1A
s95t0GCAxfvXXOaCoj2mdZikOlcG7wBcl8muzbkMzPd5z67H/wyC6pxbeLacWZRV
C0TkovVSxVHNo69xlTLswkp+X/poMGqDQBefkOMwcUVTXLTTw8aqZnlerxx8pSYw
nUB0WBWsSWSJsPm11qFxxU/+junPS8av6/3gg6sbbkeQTZ80yXGrDlisUu6SvPKa
mt5zgjLK0vfYs9H0RYBZ0IUx+g6D4sTS2B4Gf0mujL47llgWmG4jq+tZ0vS9zoDW
i7yblDkEH8nkhGFGh1K4DmSe2NolfwHJHNZq85C3EaQQSI6p9NzoQYilyftGxEQ4
iuOcDoFMw5x2DL/WGRjgrTIiGDlqr3A0hK1vTV/X8mMDO22r4IdXWgXyz8F76WtE
wfHVU25Jykl8ECBsnIjoROPN4cIiQ39dPp0ukISj2RW6n5rt6ROMNkRiuWTENWTO
KLJy2bPzn1gs1SBjZuk7hbc7KVL/65Lp4UlMRBmyw7tp48LkjzzQ3r36WrCAUWFI
9wWO4bRBdFMh8Tz0aonhJ8uM1S+Atx408TekowruFjGFBG8/kGeAXhf2HLNSN+1F
Yalnkn/76SqDPyHddAexgIe/yc1h76dBya2F3plox7caxrXRi4vTbfmspt4p0cH4
Mo4exJpXv7he8RAgtm4kjEaDNLz9lkADV63R1lPvgjnyWc/nrRClYJrVQJjJ2Uxv
jgaPbAWe2UKTjk7c1NrKRwGTWfdqY+Nfyr/TZC40rGL0GLolWFB6S29TgVvtzH73
fNBdLeVtaQR1uiCUI4uAg8CMI38AjC8EXHjroe1C6F2Azb7AS5rQdLUiFOt+DDz9
n79RxD5qd8hKqNfRx9lf1thmgH9Ur0ACtj1AQ0uyKo7TVt5JPnsINw1Zb7XgCZkw
NNV45JxUoI1VmJaXH9qlYBUGgroaPSd22OWQ2GYfNM82uFvGFliox+NlYmCUEU3s
tfaiLZx+zU1ZksxClcw4LWoKBzKgBhe9LHKBQkWNQizZpIMjhSY1+HhgakPmUuat
c8Xly9EVLLKYpCkHDw9x5B5TNodcb6HgOgnMezO5NhIjOZ9OemppT2TCPkVQvvPC
vJgowmqvcyVWbewCoCNxzYWxPH9aT6SCOYGQFa1zRoDH5tGu2kgm8nwY4d21iH31
2fhE+j+tGaFhMvtvjNZ5FpD77PRgjM0mwHgg7NVoPeTVQ8VWRcK1gUeE2kKCTqaq
p0QTgEQhzZHfzXAhpec0EgNsnHzUrig5qedU812SW0XQDTh3OK0eDHvvlhDUpwmd
62Mowetfz2EzfyJ4o1okSgjfflWWLt9EEc3EtQlYTAZ9BCJtNJo1kufzqDXttNFx
QxSzZ79o0CY+e084X0ak7BZ4V/MJAJpw10QUG7ytcDX77P53w7OYdsGx3cT0AtB7
uqw/eg9/WcnMQOtdj3meClh4QFomhl3NgIOLwzHGBWsbL0jXodatKS0C+lxeX3iL
5wZ8LVLgT6DY2EPI7q9kUscIaG0JmIbgwNtlocDZdF/mf44TyxvM8Do+csUtKt3r
K6MaI0RUFneRKtemQOA5/y5QEDjWx10OiRidJbWN7HN8UwUJh7/sKVNx8sl0A/qo
UR653TBkDNH+P338g099qESEWG6kLqg9Er5vCWBKTd/aW3D2+zUVEqrh6/3Z83Ye
B3t/GD1mBFOYn04j6M4HjtdwYIJHNKlHBzT3QTqHP7KjQ1vExtsZ7ljYU0CbbrAJ
jAkecbePPMz7XG8mR0AyFywu+oP18RewqUTBUR5yQ8gNK1QYW6qPCCoL9zHVdFsC
/QFS6Wbbm/vPigomokwWv2KTYJUOjd2D3C/yZ4C9OCilTH5TIXkPLT4CjhqiHEmF
TWEa75IPWkaSWYQdoSFbMFTKvnIstZRM+fueZn5cx6qxwShN5Tgn7GbP4J4s+nq2
cCCU8isc/75NDbpFEJDmK6g+GjVzqb9YzqreGJPghzzS1Wb0FUXEpv6zbNBibCje
F0cKuupunsXUEC8xPoRRxD49sQdS+2tik9WdVQAPnxvR30JDjnjah6KP0wSRS8S1
puyEjFag75jKbuqFtmoMhjTIfhL+NgpZf3yi4TFQ4IgQI8ugfU04/aGQbpcRNv5V
/ETdn1a0AMSj0jC7fKLih8wzCES5XxjlwFPCQYHnKMdlsDwKzr0wpLdE/V/pEKIe
A0e8OZnzagKUmZis3oMdZvVhKvbVQXS35X4Gi01i+WShZ7xwCqHnXNMgGgVCL/67
HzvZe7A7a67uqOWEcZvYsK0gbbAkw/LZjLkyLQWSAHyCDo510vuZxHosDbQ5vpTM
5WvFAqpGPzEGzITuIYPdQ+RrMTX53zsEHQD2URFg6ElUqrBHw66vo2kMWOtfV/Ia
q073pLpXqz0URkWPqtFG9+/nEnJ891pxt/PjeUKX5CLHLyX5WU1Ezd3rlXX4t9eY
rFGH/wNUK0Nx8xMFzaz0aYyIp+q/s42p6A6uSXxb7oID2wC30L0eTxutKrMNzyDX
9yRRJjSikWqEcETc3Ht4bq4iBvP6cTP4P24gvG4go2wjXV1sxWmlBHpIMQLBmOO9
l5hbgk0ugXx7vZOthso1LhUsZbyXgj8Sg0+srWP03+6QwB+i553fgTryk5ph+UTh
j2B3zx2bkMXLsZEZCXECo9E0+GpblMx6WCrJzSZtuLCZnQlPyLykev84ABAGNYSn
8UgJCnv9kSlDIKD8h9zVo1WQU/jG32Y/bBRX15fg5Ue26bFqUZFlTIf/0HZ8K0FY
UwKZJsIU/dY6JQyzKLvQTpQCzKry+uWv51wD2MDG8FovQHv4Y1q+mZWvSwUxYYpi
gndw22YFB/iPFn+VDJDBPKyuivec2fD0OL8SfFRaJVEPmaJZzC/CiuSOTpsBg/Vs
pcPb17W0M5Pr0rE9ptOHgr2fWCia9GUK0hBxaWcNNxFw7B7Vmym+FrBcHlf1kCE5
wWShHozlZGs4c+YGZ8RrLRcOX5suH3NY81pSgwcOG37mhjWmtEzFTcdnoVdY0orC
z21UT4EjgH/viFZaKeg3BgilTTJGs4z6T4QSf6mqvTF6JUthT2STmw9ljeOtsLtO
3VQpaL+EtxaN8T6XHgnsTVVjCtXmqYtaHb2lqOxkscdnsbECjeN6X4cmL2h1C1dY
XCoYtOHoKdQZlpTtvREDMG/sM/fm5J+ag0XmS1JJYgw6Y/olWEiHNiR8i5s4AOmE
FAkmJWDiEZNu4SnDqnAcJaMbBZfA+Lkdr2JpB25csYQ9CaT6Lxo4I4D3Ryvu08gP
1cYvojMf+Lb4vnPvTeItF82yWbUyIM6y/Lbg+mCV+YFspJx/f+BDuCDN78ICedZb
iWIS/vHuea2oH8j0NDEF5Enz0/Zh9ZGLTEv8j9qTkXAGlnWf/i1S+dhX+sgO7TmO
m/ZE77xiID/OhOcxwzz00UMZWj8Pt8Ej69R97KopI/ZahGuGlLG0Jh0LKVvS4l35
iTahOG05yPj7dObABIdPEry6W6CBXROtS3daaSWEZe7KlQHD891TEkKrgZ7LdTmg
YLoj2rj+c02HNTxEJ/0IMeGOUGLOCzCNGYV4PUFHVESJ+e/VVtjiEZaH9v3lLYWK
9LFYfRtvmksc/XYyrq2mK9VsIxPgA7bIyUCTOESt11mcePIJ6dfmb9aCVqSj95fz
rqNlKHXB5WBrWOA1EpnC4jtV1YHB3Zn4WKpKtT+96v3eraETfDISWCP0a83nZTey
uEI0NFuQqmci0a/MowBLW/9BNMRV6S0VhqUMcEoK50Nvm0LfClEJhetPnW15+tkp
oetMs6y+1P2/NXX2WAF8dUOJKeHcx0g9Pd6bkfKCm3QKze7eRxOGl2/RNo3A0E74
VTR9iT1T7RmEMoY76R8keOxo/1yY+VaW4pcNz2XgSq426MaxPTP2z9c9YYiaTsR4
FLpObryYMy32rdSLd2iwgQU7Z9DCot7hQrJCedP/LtGak3HSxtSkVSo2KA+LI/Bc
LYDjexRclSwdwJ+b7fu494aoBaxM1wl3iKXNt053KqJnwmKQgF0KGMTHt05wpXf4
fP0uSKc7tKA4VuZ2SS2bXCMU9PDSBxUta+NYWRto0YQ8cr5ba0rXgKqNnavWjJCe
99UyWuAifScibqYRAmQynB8BYPEcTxBGQZTgQ1cvaclgYlM+VbT1cpZqoJw31ZpN
BfsXjAmJEMWWwXUgna5AEgSd6CVdLEvMXM70dG8r5GQvKP7MqfESI2mwGWHBI2Jd
mD6IeKwg8H8IzIrIMSxAPxfWLNW/jaNkr3iP5DMnxu4/xPBrlhSv1wzQDlRCgkbz
bOhMAysJiOIPriVEbA+vFywYkjUPFVMjtlWOv17VtXR1WylHdMWCRVxjTTkgk9iN
JQSUM7ZSXiuEPiDCmEBRp5CLveKF7fk/mL/MnzOWcll2KBS3qJxqycNpMiSw5uYl
6S3Qlu4742huDkvFGo5eLgjya5t1uOM7v5pA92BIawne+FDIWeM2JEUIuxfcOzFA
QPowF8cHEB+NKgnjbYlDIqOdLK7HESr+eJvRKVzhfNu8PrH276Ofl5eC23Ur5BLJ
yqNUZWeQv00MhU5XuoR3QZydhyXOU6PZiWTpZ3SKqSKQcmeC7tdTJgn/aH9xyss1
VLlZ5eo0hgB702lxIUGN9UTk0db9VyXFX2WVNxIuEmXa/tfi8PWy5D7+f9EkVXKf
3v0NlzSPGO2zm5nBlDHlxScZdZZ3vHroineh1C5jGZUto5W1OFbQUg5n7/YtQmcM
plcWUhhk9D2loRgZ+vbQ7rD/jqPXh2F231OmjmStEtrfFGI6JHyv6QBwNxcZjfQa
+W9pR8ClzWPBQwt8CQYrt/LUi7mt1SWZm9d/d9fSoBsX1ltQlmaoNlSAVVDUc0Kk
Hb0iHwv1GG94ZTYIiXu9G60nivDZ2vkjc6yuJp4ZCzDCWc3B5s7PcIix+X3bNAB6
jzUlfi3ykT2Htl7Zzj3qcKJF95xVh415d8762SQHbbhp0h7CzTrkXDWt99GM9HAk
eK/q8B9l5Qvo+UNOY7A1huDnoT0tk28CJt3Nee/a7EKhYu9sNDEVN1LcVRmjLDt5
9qTiXSBp0qN8HyAulEntbp5KijCMv0PJx5ucgUwj/Xndamo4sjWstjuQQ5574Yu2
FeAyx665A3yfDyNX6dtvl+TpGE2Nx69r1wuaZWP5x+Rwvryhf9jENWHKrdx04hp0
fGvNa0XK82viOPoYBcqNAubv7VDSuJ7Hkb1nGL5KbVeqr3FF2tyJQdzYdxdKkTJo
B3+Aoo4bP8clUIXHXg7Nw0dh2oNVzWnqH+AKosjZoxed9UxeCiTTx2e+oLhyNo/V
cs2Y334DUN/xCkQe1SZK0z1Ocaazu9tHafigelOHY5AYfafRSwPcmqB6BglZmmis
mL5w5bZH/mT99fWsM/XwFDmNZK6BqbeeRJ+9uF4B+RwqgU2hTV3WAA0kmjpUYlnE
q2eiiphxFFBrMa5yKqTce0yrJt01cAeI6pqda5X8PVtOsHFJ2eqewhYWV000SeLD
+p+5OcGO55WMjtnljb7I/G5hUk+sA/RYiR8BqO8kg5uLZuft7Maub49Kdd6yz7af
wN6wC/WKFn4U/pDy1gYf5uExd9fPlOAVzcJHaJfuAcQhQOtWmiuv71avVgl8CINd
mymC3Y04Zh2jrnabwv71bPnd+dDpRasj2f1WX0Q6GyZxxKuggvNvoDAES3Fu8Ncv
gp1DaQDOTTfJFuotMHsIeHgVbxYAjpJ486KgV5kKJ/Bl7XF4snsmBsJvpFeXO7EG
o+GJlcS9rtxoOQZBZ+7zUkJsmfbGiBqaKsiy3kU3Q57SY8BOkNpYAXq71xqd5J5A
Sx/59tqXGUwYXSkuWW8SnUnZFhnBR8A06JOuj29wKMddWqrObZ0/vsss/3+ssCZ5
wBR5ps1iOZNikAQ+sH7nauZrg8z8IjmvKeKhvvxMxYsBvuPT5wv4sjZTTfkFyHt9
114kSBs0qFJ0BDoHDU/S146BJeK4SBraLevGG0Oj2rU8wgKvnxKh03CawSLK69xk
9mKnKCzs+M/3U8J+SaUzVjH+f14tFhmAY8J+0ubwhvp2Lby6GPzlqt3epWDQzR+e
iVMiUlHOSXXpQLVHLl/AGYP6pVdrEKNbZOU0xJY36jKK+8YvPPkgS7rxDZRYjszO
z+R5ekG72oYDwKMGAf8opwro59z99VaCGr5T86QIdUWQrgalbXOhBcmA1ivXdkBh
+0uFMuQpxQp64WSXwwLhUy7E3eNd3qcJAqTSxTqiZd6mbXZzW4CYZA9792f/6gQU
GrO8Kow2xnVcEKd1qB5dPcWHvxoLday9HtLDiLez6If+u4Vcen+pvjftkkfjyLiR
9Bw10HFKMldjLqTMqhLhvyjdLYThPQmQMlkaciZzUSyZg1iorAwia5TQPYArQ6IH
pXu427sD1+9jzamOUqUV0YwrZhP1nYtg1Qnu5tA1aPGwWStLAZ0jOa1UqWT0Sye6
hd9IuGSOTb/JVb6kaIwa3K/A8FHwuwVXEPWaRGcCzybS30lVg/w7nKL7fRXMf1Zs
yU4yIEjcpOeyUdG7Cai7iJ+pW/ryVLYdU1nUfMJSmKeAkVFT8KWfrddaG1SUSfyu
9dLyHWi5V69qn3L2l8ELUWdnQdfifpza0UnUdYAD+D4EA6GfQyAQtJwFoCV1uAlJ
8ypksxSNbxTAdLYHcrgqm4zAXQ8r7PVQE4+CIchj8x9p41kf4P7ixBThwsxacZQJ
qDTaMZLYKhnTE5K8A9gpa+iUn7cBcZ4PZlIggMDdrlfCmE6GrCQtaC6XOcU7AwwF
fLeLR5b6zoNDch9iG8apNIiqSbwk2Zm5AkIibXyA4HAa5z+sAerV5SWcoZEsctEb
dTjUASteCpEJzFvWXW9jO/EWaLbtmElq0eQlX+OSMWyHoX0tnmOP5Sbb3OLTbJri
hFucMO+qVVwzbyMftTuGrWhb/R8g5dBsqusv8S9fW+q4VhCxWomvzo/4D39KeOWi
L+GKEOtk49AT3k7W2e5bXeoZYgHZAPVoTwLdBQYb2WlJGLm/xdQ1AHuUbZNIKCfB
bvSsFgLGdYsJ7/KNnVKcFHHkl/ybYmyIbDsfAB6qTeJKPwJWvKh8dduirwbny4QZ
8Kzd8XiMz/KPrwqN1a6DHUI1fPxlyAe9ExFo84G8Z79gMf0T2GSJrYnhe2Qibi/5
FxdvUpYmkIkAOkBtlpeZezfR+N+DuHWq9T6/qgq9e3VD1C7Y2niun8DKowDEAYr1
qicixutc+viClL/ojVG0WmP/reJYWH15ZiJPKkxBKU8cvcmKoW4ZyWvTqTPsHGJJ
HLm58syFcc/S/JHPxYiEmpzqPneaidLCuRGtd8jbk8F/FbJkTHXkp4VMJzmDqGhL
jbQ04vjesYbZWzVhrMSHrUdZmpRMiUmfV0n4vYGdHxIBvjxSf4KWKhcmSRdu3ah5
tyJ0+oXH47wFn+iSTSAA+JwhxkRDrVk4HDepEuTm09UqvM7dHFoQLLmk4FrH+keF
6PMCrWQBv3Z+RTmcHDnVKNN+jKiC5sosquOXs1hPLjEfwzsMkoS9k4sbDHQuqz1r
s1iLLdngaKC+aiBbZNXalivPd/R4fIZL86Z1Pt6GZaWZNYosDEzjv+r6H2rAgd/i
uUDOAcw5zLY1SxRIUUWNIMU9nHm/bb7b26EAtbFyK0Fve7mNhivNKTsbeS7KjSRd
CQDJw3v5N2ipaSq1JN3QrcPGJ5/fuM48GBGL83bxvIedw7nCdUEjENpW82ayoMrZ
nfoZ0BIa/1zj6QMk4uUDTq8pikfH5QPQ0q8kE0/kf2PuhiqaFrtqKlbYnuaA9Ob8
18Uw7vzeXKcHeHGgz2JRtEfsEhMIWpTqNbP+CVQJTVU6ZwrB528zM/H+O4XHT/AV
hmgwTo5+d+rL13els1/CS1zAMbqfTtxJQT+fONkOkTMbBWEq32ja8A+x3SjbkoI0
KoG66cz+YiM38vZzNWOhu2xGfIozOOy16nmrDwVbvj66syc+s0MwKbUN0kWJQbqp
xVatSHpg+L1zRoWYSV9zg4nZ8YufBEApvN20CQk17Rt+z+YPjGnaPRZBMuNfyCjQ
4euu3hdiqFt1RDimT55DwRYhQjuBg8Fq/8zU8V+K7jRA+Wx79PpR6naJOsbXW0Vo
xOll5tBkoxebb+MTwQmqoZdsGWIDpMZDJs3p9EL5j6uLO74yxPaGyl6XKdKnXjLl
PTjyLIY94lGfnfQ1oL25RE2ONDl9Su061fiuUJuOzRATE5OJvfUDrythC9AekwS9
JZjkjpzfFdhBzIv6KlBzb6H+Wv5ZxDcHJ8/28rg9K/ATujWTagS+8MiQ0/3it2qO
EHBi1K1KDSpUh5a75FgYenMxfIQL7cOOUEeRCY03faKKOfZQkMofNUrcRDSA4F9D
Kb5GKHFHLZoMhDRpqZWRXl4AaCH+lqGR+3+xJNrgh6Gwebom6l1+EGP9nqovALed
Jl2P4VRU3jK9ws+RYFUjD0BxuyREUhDuq6ndUTLngOpTo5E1Uk8atwdT1rhNj/BD
9As98s39m2IlOzqPjy2wWVgi2VgJrhvLe4BB4iVqG4NZTB78bim8N8ASwi0k9TcR
HqHIXS81ozDcXuNjzeyhEQD+5/pT5SilK4P5uKZU5kmXYKTYSnL3CvOfq6FyjrF4
wOUDVvhLPn015Dxz9ktuYUlUGyCbIkFqfyvVWK7E3hTg7nqOw0+GmJzx3EUbFwR4
1UBNTPT9vh+yb8USQ0U7LoMJL+aawi4kjC58kW9soZ+ZiIPe+1KTSDMBPUrhFLRp
dhfs5ZpQu5PRKbgE1pk33Mlwc0s5tf/3AY/TMAnVCyPON4rKG3fVfyNzyyoap1bV
w8jmw6//qwH0cJGWYkig+YhaVsEomh5ck6o9Px+W2WRPStYhoQETrkdaUdb67CSd
jkL15AXOBE1okCfCpQ4ATx8Zr/gp9alMgOX3p6mOi2o0weB/8Yu6HAWAVTKxEN+a
QIbWjhRyxI8zhKXI82BQFIGLNyw6U+d8ib7zwqJV4CuCKfLNQvovThL/TV0+8lK4
481Z5Bx02F6+0Q2pLdMafGEARrxNgrmKBONvrTmydFiyBndA475w9gBHPSw2UOAc
qG0gBgUATVF8gLQUBQFS1IJDWMHPic6aU6SntXOHyp/TvXMqx2d0tfDnlVMmqaHF
fCr6Wc6KkBZFA9dYdZmvxu9BugH7/2B0INnyrcs3LUZlpsuT6f9G2cZuecloZyHo
HFKbkEZaYhzTjjh40HpKFsRlowmVBDv6q2h6AL3zuO6OkGtHbVyLS+LaRsLTQZfk
ZhWpm+/kndaIfSGdCJDZ0SksjhfscP8aJ+8bcNlR44Xxk35tqWRqnWv2bY9AX6NO
bOYKKkEO0Sn8bLbi2hCmlQzarbI3IhJOhOfJXHkOedKP7Cznkv1+virWCPs6pwFH
1UCv2yWyA54DtThNMvOGzISUFMfwhuke0om2hJjOFVwghDf7YZZKj2OpFgp5ZeY2
a2FHn8h1inexqIq8syYYG+dV7BiwUlScY2C/mqL38GUiap0+veApcdYJAzFawTCj
HJVwr2wh2DRgdTaZNvsgfRe/etaHSlFgUNGIGp+m/6PPOQB3JJgA9woKELKIqSjj
9ph64gRZ32IIp0y2jbSLHaGWumG/zqPZ9sQFSSmS1eU59/94BQ+aeLPY3BDE2P7T
5lqt/EP6kwCQZa6tkYX5gje/2qbC1D0t8Yl5g2qyO59gHo2yyir6fY7k1M2bNQtw
rLekN8MKWxnq46M9dHYFYvh9RB9AkXWq5X55MohzlA0ICIQHibER902AaWG3PjGm
3SfMwav1ONs6pK5hVA9+QNqX7Vvlul/x5QwsJ79jYMEdTwLMSd3rtnfDYn9NFlnj
rs3FLUD0Y7Slphs2YSuJnZ3pJYhWwuMJwybqMLn7krtm2XYktbd/ZmCpccZ3c2Av
ZaZXj6/e8BopIyFX8vux6ikPCSrQp3aCFGJTYXwK3VS4zie70O3xZyoL/jKwYo3v
PF+xcii7nrL83tCQD+eGJMnN1PH8kSnKSWuZ+5otWGppOX4cC5x6eBgNWX6oD2es
XcM2gPyzRr78tXCzuWCyAttGJpXZt3BewvIc2X5ixyx/aFeT4gukly0xS/me0t5n
sSiWYrITXITGeZoAiHSdnR1Iu5kPiNHNZ9FFKuqX2bhEngrzhy41XGLFGmEZ9TLg
k7TzAtb5t8xki2uYAUtYsrVrzpMcb3c6WtHiDzVfzaZmWo3PEPOQzhmrQPiWh1M7
xgj6svbisHTfZzYeCpuTa5DfhuLHKPNViXblW/oAnsKyMDXXQcwsuiWrToxvlAcn
/dp/B7N2OsizbdcPy7uEMdFkcTEOJ6PyUcyn+vHein7OPQ8/TJgDU1ynScpUF17W
muBDSW7vGokwRC2C1peu/0NYRdgU0xqA9kolJUHPrpFCpTvpgj7SCvcfSZcFS2ti
IoGTgI/UU0ZpKstX4yeA5oDJa4sfzyBzlBZIKbXHjj7QhoOq1E+xXvZILkU79wIl
bcmx4XwzZzLoLJu+Y2/hLpQ3H960Qr6tUeW63Rl7V2SsZEDONfVGfCsGI0lLHtiX
cZpj93ASxqN/zQ1hy6cjrq2I6CfXjWFCk4zU5/o+LtSsXJ7m+q1A6kYwE2QgdsAv
hsxCNaOc5TbRr7uecQSljY/04m9w2yunD0tzMlODCnZUc1rvmrMvhxE7ovwpLgFG
dWGh3AJRhh2CdjPCdyWAbDz/H/gneDnf5OBQvmTiLl7P5pMNU+xQ8kt9bieCCvid
ZBF1s+81HvXrxFQuvIPpJZeqsjFHJeF6mVH91GeHUnvRZZvPgQRHAEWL+24nclE0
ufkxmC+xDaJY76Bhm4UDAk3bttcp01NOxNhjZs4csOUzKkmDH3g3wHYSscsXc1eZ
KizLfdDFl6Pn6w/PVhaWckdFKwnciYQJRhn93HA5T7yOW+BZkqjvUHVffzSKgDFu
oJUSIOmyyWaE1sRd3FH2wTJBERj58+ULOXtu/PmXMhnTx4iEIKvDaz1T2NBe1rXP
HhF4r3WJTsoMdn0dh0Ma/dbP4FV6ENavzZ/sLjGq3bNHlqcmrZCTNakpZnWTMo/a
GPltuDNICbofOD0ihgEHrUqx2KfMlzyESh0h/4DDi2vq0Fs7ltMs3cS4z04t6mrl
a9qFXxwiAra3+8CeVDIBqTfUyU1PcK8D/B2Nfyv0t23ZOdJVOAoCPwmLP429X3Tb
hA1SpthKLc5ZU6afnbdxDq0otasotniSCT33t+STFn6W4FaLMeSSVfW0ZEa66MQw
byTdeQaIZ0GvzEYn0rD0sp3wBEl6rX+kr7U/pcTmJV2EdiJ+KdX65vHjU9ZZTk34
yOfSmth/olVP0ArCKsM/jnpdXGqzvdNA14bALBoRJ8M8v2sExMfpZOPtMS9nMDoF
vT0Er0kLh9/aH1+lKzdP+AUw+aKXbMUTsD4nZi8wLusiD74XNwG5G+sTyTUqcphR
EfDqnQ/c0uKfRRG9Vzdy8ccfNAZoculIPpF5P6QmDIxADxv7TtsWSixq+2xxW7wO
xutXYJDPIr7Q9dRI4W+BjGeqOFvIyPu3q8yUpgGGAHzF729VOiNk+oX2NXkuMNGX
7h4ZwdVAeL8zrfs7VlzdYUpN8e3pmxbvFRdwhGwvFw0dJ3UJ2NZgojxuaQksiuWN
oB+uSBeIfVuAEUQy6olyCEosMHbj69A3Iged2AVL4KbTOcJMyrxplqlxMNq5Ah3K
ISyDr9U2NA3wf/p2ldKj0DAy+tbL8eepTo0JEz/+VUJNA5WxJwkYvCubjrPvR5jz
/wtHdMRXjhImos6g0F/vU2ejJVgT+eRrISIduH55/qtFT9nxp/mtrbMIZ2eO9xKq
cJ0aDk+aMBuhKGuxHM9O3L+a0O0gaOXbeMSo0u/H57BF1uYO2dCRNWFyOz/PFkPW
spuiOiEUbJTnl502xWwr1thL+zfNDUQ5o0ls5/fUm9oAWs1A11qeL/Aksif9Mpx6
a1yRcvywwiZbFIeBEzx+bQmP9v4iPQ8ehMqlX9g3iX07t0WYgf+hMei9IlscIjQN
puP8tBrWeq95hGOIWZQR9R2QhBCEqEcY7LWesa7ZtVdplUeA5lToMStmiX6jDEcI
VzyyiYZbtn8YaDg6i8u5JTlerZ+1u5WpZUppyN8hCrKYclShY0oK/vPk+TOvqGDg
DW4mvqRguGl1sSBtJcxKAAkm0hNIH5ltgjk4UUllOw1NgSJIGzYo4T62ozE8X6xl
Bx6iKAOb6uKDirM6k7BKsVEusqTDowM2qh2TY7KM4rgHwIr9E6UlO+kowzXQS/HG
DDPUtPeabOr9nmWcGx1uvAzIOHuYCVdYyVGB9OTmVnDKd7pKwmqHZzEuc4zMlGNs
w4SJQdv8H81Mly3L2oj2aJM9VPIa/8mthLRS2IlXh5p4FRsY5oegfoKcqWc498n9
aX4dBoNdKVmM7Ig49OSDcRJDH8ai9ULSN4ki9jgppykvXbqxhlao4NtLyiKJ9/Cj
1ipOSDZzqqjZzMKCyB9R0NHlg9mAGKW9d/NQU2ZLqw5R4O8YBnrqgnM0TbvTMZIF
5uvquWY6ZnFPXL6PWkTUa20U2azWaZThix9W5v4hUoMzabmJ2pUnm89+BaqNlQZa
fbbfnZllIhrlkEsHFSH8SuqGP6gSaSywz1fX9y3jYz0Ll2bn72apwFUNL7gcOgXS
BxhALUCMg5ttwMxg2N4ChSJWmoReDOpnlqmAmrt4Ans29LemczXoclYHnYfc0hdF
VOGO0FfofB4y8b5+RjZrsA3Zk6n9L6btT+jodPufEkc+UUHhlrDCkWM/J8dGEuVX
gwKqLTsmJDfSS6LRKQp4O/H6PsU4TV27m02Fb+d0EwSOREcBW6XajsrgyS2wBhg9
7pUJhF4+INMYgOfuN1VGNoAKLPKjqySecALmAUMhjjloSacFRdt20IaQrKL7EKeJ
/mlnYoUOgagiMyh5+kWyPQQS2C1jo+0uQFJjA6VvlC8HGZba0ZFqUZBfEIKHQld6
s/YLW1nVXtSb6hLmKP7G+AFykhcaTuZoDypVWZmXlOgixGFS3F8GwRGg1B8fNRz8
h2etfqoxPMm3bavoRCwk7eR3WuNsUyIHbL9CEevTRfmKvmQkwF75CFX6jQEHzsEa
HEzsEft302qMdJHIdFQrPuwSh+xn1QMOyWwFP0SigpQlJnQw0M2gpSnnlosyUI0+
ec8SPtIxLNmSZ0cMQmLWuBP/EaZu2rLaOTpj5qDk7ILiFMRetCDIqccq5+/3XF8E
8FHtYB3/nqaBoZbqNKYVvRjS6wsmLl+wIWNZKjbsT7BG0T46VgYaLnjBJhSP5Lv2
o5qJeXu/cmO79kQkopA527dFauQlAOds8Y6h5y/Kgn/uTU6Nx0uh3y8XNL1GvmDS
0p0kiO+BRweWZHtjCj1hngV2nnYexvtyfa7g+AjCnMMEG1G3MHVpPGvawdz3oCcC
0ywnPeRkDSqt2BjwcGhhsbPYr8XeygXz6UzfNXv9xf3mDWjC2qYMaD+MPNwitQZA
vZmE2DV7Jh9pigcCPaH91TunVzE8rHWH7a2UNsQOmBsrlz6xuN+X+RZ2M5pNoGKu
rkbCJfwYKBDhKPTFhuXFk+VdO3g85DNdKFmETpFa3y/u8fjhKy6Bh8O8ZJcip8tV
BbuPgjQHLknRqoUEl6jHeRgurrSnMCrH+hN7LN/PO+qPBySjLdHJln/kv6HuLqyq
FJyGYYjBjmZN1MD7hlvJkB0eVRQXLNN/vsBUdoC4eOsM0Uuz4YJwtRJJ0f21HIeB
nN8I/OdteePToYnKCrBxINhJYc5dsLoVmXk33VJhXHV6PIYn0FwvceWW8g6Rj6rI
ADS1Rf3P/gLKOUM9NzxRA6iZtcXmRzggcUlPf8XYxVVosIA83mZ3yFSg1jNGHuCc
u+vLDwbRdsGA8kBQjywB6oX8fW0eJfwUggpnaJmLqJeCKgiLXvdJyDduwY4izdQk
fcYNxppub+p54svp3Ctc5obLzutdD/oWmD7LN7jGQX3R2PeynztkoK8mW6LlGXGv
S/3E2JCz0cYBYqc99XplZm79cFjkkLwSzP9qLF4KmHoLjp9zUVbDvInyZcuuJv5J
x6ELCysEU7BHsoXaTIcRFZJP04ND86TUsKKNcFh/6mnWqkEiAQ1VMEbSB4cm/aLj
TCsG3TiA0npCMN95nC9u4+4eAdKWGKtwxsb2d3SI5wmHlnqN74oUmmGU95BlK+TO
I0rCyzGMmXTxgw7skvdBzAHVEz+wrrG/DhMqrUmXrb1xBVSSjEVixJ9zsxdWVEkz
Q0gU8qOd3Rm6EywrVgylvGh4bXlRpPOarGEsW3tyYi2xNvbu8GyNO94AwMelJgSb
rU4FS/JRa0c+6RDl/hHZxOZ8p3UdxdRq0LWbjtERUhfDN75tCKaMtD2zDI6Xo/IB
RkRhXXyfxPEl7NSRpffYA+8YtIMQh67CSKB6mTd3+Eu6mz28L5ahQHbUgZT5ZuBN
bPQK5YMISNjfQ7P5XedOZZtA/Bwd7+617v8UyoiGS3eTT40QegeSqKx/mG1Kle5P
1c3NHK0qatnOBTI+GJDsnVzwhqwRU2a7CcCd2T84HJ2+KRhxoXN7PDNAgGD+/fLJ
JTHnL8aNfwY0XrkHkMlxVkDhnAmJuseDT+CUCmIP/frF5JXK6VdI3HSc59wD68QU
ON/YEafOIB0kC5NY0P3sQgqv7HHZq+8FAA1oRWDpyCbVCmugZQXuweKQ8OjjxLt7
uvyvh5o/kj5YuuMnQdGctDELFWj8Cs0Htfy4mNdv5hE2oqA9V9x2PpQak3NJLSRo
DnbH+XKPOWD17XCavNCWE0UdBG5wsYC73XemMVW5pB6ikLThg8C+BTAKA87J9U2Q
mX1WY1eTd6pN2YRbFSqNZu63SeGFZxfObFFmsCC6QaFHXZanv3d9YyagaaRttks9
IdQeggk6UxFYcKs6iAfBKIEf7Ju/Jw5IoOC56c6xRsurMFoc21xnlTH6WWevspfr
Wx82ZAOLK4ShH1+L9NOyJ2nEotH0lOKY57FqG6cqMx/QiPylsb/Ekx5cM8u79g5C
e9MKsaXUoSgEIkBgm6fgjLhshGT+ASU/jec2dv/k9zoPTe7GkwNgw4LW5MFj2dST
hUSUhj7uGJVreHPqrTkyDV7xrhKHpKT9SIJ3o812vMyGIBPoWcPTAXBasxsPnGEK
aueq7fSgnJRYFFFkA4wzBUNnHv2pGn2lCxlRajyA3OYj+ELfEIM3jtnhx32YlP34
yYWkE4pF2u2gmLAc1ueIkhIdlzMcUW7k7t1QljMre8v44kWxylRCZDl2uf5+bzxO
k3YxZePRtch+MGNq2RVz7JyxO/3oKStwlf0daRxUgtx268unoSB9vq5ALh8j4J9l
8D6xcUfLGeZBnfClVJfP/C1rz6QSQZjJk6hoe41h6i2Kf62aHKtPVDQ7DAUvK0Ns
sIRNDDyIdtcZuubZCNLJoH3dT2H6gVqnHr113vSgJRHSYERTAhvLH6F6tUIkEPW5
X3NqimF82/X0eJwofSZPVFA46Ilol3iE+GZjZ72+7nSC57qlLFQA9MA/FbejpqFq
gzQg6iG2gKnKg2JzU5f+tcmEtiG6e3DPKpBnUgFTsjL0e1z0+Xoa4NFzlzgdbeLo
zNv181Au8rL2wNeZf8FH8e+vhlye6I6jrX6VVvizF5pC8zRUaKfyl1JSNubqKfYK
vwd95hUNmRKsX22mprqFpB+kep905tCKR8Ftwnn+XAx7lSOLEpcPEgLB8eShEQ0h
EXFnmtrHi4I+OmmnDh3To3ctutCMFkNXocNZsB4TcTTaoAcU1QZjPh9mqlDISTcP
FSrceMe+NUss6Qi4y63zYDQyyBoAFlFEAPNp4SI5W2JiFIYXpq2QudhtIp2mjwH3
mDEtCXdjyk6n5c39c4vCPX+R5lrhPUwgj10SzbvLnAl47nbGh2xp+nHI2umZnpeH
oSjt+1nYJ8e7Lsfx+WQ4tUFCe5idt8JolZs9IVWoWSAaHgt0/ikGxtr5NfShOUH4
iT1AWL/sv9Y0aT7g/FToh0KBrUwCjSYNwaqe0/2L/um1Z26UqaYKSaQVXQKabbnB
WgbuaFnDKdUjXAIAk38wMSlLYnH10UvnLYyxvvhpsNs/zO0XGGWKH0A7CqrOtB1M
yK0T8+Sc0Bs54Ojj5LiD2OqYcYC5InVGbOWCmp8WWm0fhDYu1PgxbbnVNzOr0s4b
ShxCfzOTojDC5Dl2cymTZNMGwOSTX5b3eHmYRLR4Qk9VasA2swFEHwjT5eW5QYH3
5Ut0LSOwHw6KZs4cxTahdqTMR1pfAnFbw/D53qUcX9Te06pEKKsxz0pMjZKoa1I7
O4mfa5isiw8097CxA5u2GPXs+I9CRJe0W7JjTY5ovbKe3ZkyngD4vLrsd3lNtOcm
pXeFJneHNRrkT3HZ9pDhlip3V0Ds1LvsXK4PFbJ3SQ8K3M34lN8Z0Raa4EBrSJmA
m1+8L7YvzS6pYRs/M/fRb7RhESH5dI5a5oWtaV34VTuEABxVTDmpWGzd1royit//
ad7wjgSrgyP9jvCe3Glnmv+fgMSuYT3vaAOvr6t4hnfZV50IY1DTvfF+1/5fg9bJ
oB16psk5IfZSRpS9NnosexnFHdV41vBOWCsKz8hQVGpLnWaBmG6DOaYJi2XlT5YU
0lsJVmZI7F90B1x/7G+jvQFWDlbLsfb5yRWR5da5v+hA/3Xl/LJGWOGixk5EwLWH
mJNKegK+LlhdAvJgqsAdA1gG6VTjuTLYJzfQSrPXkVtC4ff97Urp5KyZpYgMr3ty
+BnUzIkU8nCqC5G7GAIyxQwAi1jDaYHAZ3k/UDI6v6FOs3tOssPcYSYuumFmQwRH
9knM+b7ZEUaR9uVtiJOcg0KmxqFXRPMWD7pwDhh+vXOYAmlB+rXEaJw7PC+Jbjol
19mqdEVbWam3RKyk3TdGgedJqGqSAWHACFS5pdsHu5be2ETDbxf07Njb9mnM3Jt+
hwUAnsu8sEWJ/p5f06s69fZB9YWUXb0KmsSqZwwDOM7OZww3W1BwgmFjmOHzRxbB
ywzV5FapUROPrKWGaI8L1+grllp4Ev9Ge9g8nfmOiND+7NCFV55icKuwj5Rl/BWy
rERAJ6hJCmY10HF29/WELAtH8UBLS9fQwkn4QGZFRUCJHMEjDH3DfOpzhzgJQEk5
JqGOgLhYQi++Hlt6/PZ3hwFDKTGQ+alCuUw69bSxO5TiSk0uqxSbybNLzazrfxCi
mkznAwo+AufeYfyIY4gG6LbG0/2Y6ysxLM1GkfQcCnjqJs0CjeV/7ZU4mlv4Igdz
qQnQtY9QG1XA9z+3NvuMknAr8zcM0LCYBGENl01fvcywP+06JTziD17x/blEjbOL
AevqmGgEgqLdPLGxVOS9CvodEJIGTj064ro8vpu5evc59DFnAKFJDEGXdmaWFZkO
QZ1M2cr0uX/O9vqAK0QkRe3Hqmw96mVytAm1HB0NTgNp9GU+7I2YFdYzUvc9nolj
ZpslYIFQDXkqlzCjMj9+cZZUx4cKN4C51a2+VzkuwUeDJNF/Qqv9tfByjQUN67ZZ
8KS4CMGurLikC36/mqAka9TeBgiP3O/0v4KXh6ywTbLKU+oF0ZP2Llb8fwc3zrhG
++7DdnKufdjGbAxm7HHw1k5NxZfjwy+t1LuK7QOMut0QnonfzNWZY+ZT1lzunEGI
1eunr82J2leVMZ5lJWC9sm3rJx2blneULbuRXZROuDFnf7l5hRFTbCad4MDrhwQr
wfnD9uw5s7Hx9oJJ1UbAfJkWDOJo9OFHklotopCXwStiDsZlq85bqUxbTVYT2Qb6
yQViZ4c5SFBS3+3G7a1pbppUxN4F5SFTQFY3+WsqxZ3iD6RI6qMSNxjBkGQjeGeh
PPZtU9uwisD4OOuj1IKXsX4KKkC+qrNqyYrJRhKhTanI5fpuFbbf2ed9rYwQ+KY7
gjjhuhFnjnK9lCOPQV8KAW65VgbpMYcMiXRbHwBrd3ICvH6jHhdJGiVCigx43VHB
sGMD/9HesR9S/bpYx/amZ427HWys8D4BmezvRH4IW3DL+tOKj5HyLirhjPAiUyyI
WcPWNiGbMhxQo1L+VxRKIt6LE/l9lHULjcOH5Hzkou8S8oQUFwPwnHApm5/C/aI+
FNVynnREX3+liR53o69gpSk6d1mKoP8V2Q1F67YHWsD0IN8EZGzi0F7867JScSsI
y7iKrVIPOQdC0H8nqcO6r7SDEPx22yGSeuDnNR6775gRAN5zW0MgnVHJIMH1+j47
0g6K4kk7VzFAH64JvdEwYuRyIlhnoh7I6TnEYsIIx/98VNBxZ99jm01iKDBzCnDb
xFIxkfcENy76i3/rvmtW9Px+zziGcHLL10m1Dms4vJnACJCVK6FCPGawMMWd2auL
x2e8tE6AsLg/mnMX4pnmHveos2HSRjj2sSVlv6ueudnnKvpv0bQbzU+eHxMEPnh1
9lZpUJgiB7mMFcTUgpiFz77o107sa0gFXM7THy4VTOuYNSrb/iqNedcwjW4bLh0C
xfzriUSwKvOJ6IBV2gprlJP/WkAAF40GMwSsTyDRZKAwuINbp62s5J/4zHpV3gZm
OyeLKjhF16qb20WaqvTeebpJ+6pJ/tNxM9bAflaj/50k7cGrd+cNuuiTTj1j69Dw
FPp2hjYusCnTAc9+Zols8FaWMz8l3w7oL4RSt4CFbIEGdwHEZqVBE/IphU6nO1tX
mFmAp+YdLDIh42/kvGMnMcLPbjpKjW0j8HWVep1mitPvh7UsafBiovTiui0wpBP7
nAiW+e2n+Ish3sMKw5CFKpT/W6g+WXOPr81k5tlqG1SAfODOCi6KADRS9ThYsm6D
K8Ev2QSdieQ3S5BZEQRsUATFhZnXOhMuKqWtEEkGvJqwx2EOCWLqel0YiF2PDUKm
JgkBO4cZc+eIcAWVoSUxMnhVrSmpELOeeW2+qrRgIlw2AfQIQ3flPyJ+eRs+8pb1
t+VPjOKcgf8JS9TYsUiR14Q2VT217TQP5xiziN23eQssGW46mZWtSGjyXq0qyrPL
bbPZ1YkN+JQRSGM5kYnlceMHa84Gw0TPyZYdn7VY05QlQ88P9KDlRhMLIWazs34q
xEGYXKrVBPFsDaF3mnqO/SxJwjoIPv2KveWlznSfaiU4u2OCSk+FRs02oRawYSpc
E1/W68NGucjB/2nnigWGzcQHcvFkWBfFfgwPGcIuSzIeKoafSKMpACu++hyW78Bp
geyOd/kzfzJfpm/FOT7se+TIZoAtbOf7j3AWm9VSiSLRj9aIrvSFAxBJ3D3n3ugq
u9skL/unCyj33H1yS8snb0BsAXCNfPC/ua5HvyCteeJasKqE1Ri2UM1T8xrJNj03
Mu3yRcu1jxRhPaW4uIUiGj+RJFWb1KV5p70p1HRiaSt6vVdtbixI6cEF7152q6fw
llucjjQJPOhUkc0OPOdWd0m9l9JmNmhvVRGXj2uoybH/DiObkDjAJug1xkOp1V8z
fUbE+leD3qAhb/rQe1l4nJLRpSc2sWuuyYYpD9e5m+aiSbqBHhuAAqAvwEuiJQ92
odLbfsAx6xumWRRVRqL03h3FAvgJfnYiH+t/l3f8j8hyTndAdJFmyCAXc3kcIJoq
XBK/ZpAXUCuWjmlxEkL8FbegytJmkDWU52toLhuUwjdMTQ3TErTETPu54F/xRtnJ
s31vvGrC0seOOkunDZYBVK6sSg9CjB2NV5AN47MCFdpfYbClQnY5xiKkH5P04DBh
2KPSbzedBm1ZTj98EXd/WYZH3V8rNBo+wrITAv6ElIcezgvPpwwHS5lHc5kxQFup
7VLOiMrx2bfd4OX0XqsY8ILo8LFVR45iTXI/lCia8/VU5gaOKl2M0jjP5CbkF2bJ
4RaorpCkOBp36A2ORMp78vSiG9Mk0S7leylrIoRPhQNX1m5cpXHCcKeWdo/6Arp6
H50z0iiezK+TZ4hgLBK1ghWOaFiLKKDx5aMuf+9GXkVyk/lOeytQZVJ+xww6AM60
he5U285rdGFWt09En+RWoIxPQex94W1JKGGbC5Npqzs+bs4uMqXJ7FNzfJup2eSJ
+U19SOhvYQdXNEnGSaWRCPqSejx39qRKx2qQLfjRktiKq6Wb6RLgh0RhPypCAGhA
uYrxJGQxdd55WdgYkBTFM8XrYW6i7D/dz3Zh9r5S0OIn0V3I2JHPDFZRh/S6D6/1
RJ6yGAYTmmhfkA0DG3pNXoJq6TubZYrISAl1YCIGxp5pIMTak78JTxqR6Y1KJmiD
k/q4zkLR+hhPai4f8lfxlQpRMrKD8GtWe4yHJAmvsGQMWIC7ssd8a5fk+V4YRHBU
FDWiwHuvkYsem83YkWyOUW23jCiIF8vyNKOgWztCi3+cR0EdIYfm5jPjqDsENhX+
08iKEKRX3w+yvbmO3jAcnvO6y7D/TXMuF7EhXRgSdBldoguZVb3DpOZ5wAum6X8G
CaxWif5KAN/8lPeRUM9FmlEte+lpQ2qYx1i0qtm0JKQeTLkMjf6mPewMKODJ2/i/
ye4qXawvE/tgjFeMBbV6DgDFAuCJYzuEwSUaRq1jVQpM3lQkOo262i/bmJHtRGSl
mGjAw8Yx0m8J4i/OLbVCpNz6rnH0K1Le16QQqdx8TF7Ig5d6Vq1paqmpOzsv3DmG
+4q5ZRnCYgFmNGDPwkSYjaxQVY8u+feICnpbk4fxoyAKiktUm9AimDc0e+Q5O4qV
56vMa+uv6WEf91iUFWSHwe/LrdYFs85FZr5ba6YBxDqmqileob8oytXgrUVs0AhS
dw3BqOKH8wo9YYv6GDet/lGncTMlhegP9GBBhGXd6CO65144oGRM8nmaHCKURV+K
BmhKuBMM4m0mDhoS2hzK9PyjNI9iZqCEc8Cby5Er9gZtdltQ0OnK29hLNoWrQxb9
/cS5gA6qyz2G0R0JIl/+vW3FQO3N7WMLl00n+mapGCY2XcqVLX44ezNG6vA/aDcp
FFNhyyhjil5TsVqU2jEm3y1UMo4Kj8HXVOdu+oFgZ9w/ImTGDkVLtklSJA+iZkTO
/TvrtM7TfxFtFMQCeTWTHcRvIv2N/INxaxSn12DTSnVgkcxQruYCd0lXCkkpNKj5
5M6G//VbgghlFXrrl1864xsuhX22gGP+XBAh4bV8IsTOTvyzAJxOuiZVj17m63lg
avXm3kFZkEcweFQkrpMm/pEOdFM0Khc0qkKOIBwT+ihlserbeZPB6s55VGJFh2HO
Btz0BTzeR976kGuFYhzhZaYnY5Ty0H+ujAm2fPqtQnBxmaQhP9aev9M7dc5AI9hk
ZRN4zouX/M8xkFT5Fu3BLYW4oZ7bPOfRP+YfiqBSchBTG9lFIUpaLpuNQaZMkV0L
vLYvyOGS3yos4VAQN23+S4aUT1yq0SXSYRCAr+fKQfBfdXGY2r72umVKvDATdeJ/
tZTAnW7QBNDVxNNzYpUZoOLDT0xKGLUJU/TINZxN30ppF9aam9bLP530Ny8ve8My
bZgJoGa5Q5VQ7oWiDireYW66x2JNpn/HMWjM2CWEjJFju7dNDZlFBWeA7QdscyXi
CM+3Nb3kPurJO8/ID2uaSFECluBSP2MtxZY9Fn6Md+xD8GtPl4P11NiY+yR18mCK
HrNCva88K4Pl9Ddk5Jhw2Hps4GnrSwwLJUtEPZbqMGLrSM7fjoPc0HoQTrVBg4Ki
oYt+ZTpVBtSzOmv9PVSeOGD32US9dx/2CTOXlRdKZ8ia10z3807Qp3UZzR9iLhNV
O9KuB6/+ScbF4bY5iVe1Y6XUGHUcuqnqx+os0mCvBt0BhUsmxkoMRRYPz3V3tXFI
crOpi96ME4Sl9VmtaRLMfOlKPXHxh1yKmKXMka5rRMJ6y+clILzdxxWbA4btFT/2
hpp8cj+aC9OVh/FwP4k4u/atNb//Sq2dB/EcVBs5TTSJCZwQkQhDjId1HEJKPV+R
zqt9ZCyRmeBVK769GTxfa5u4dDJgxqiKluWXGa3Dx1gqUwHafHwsbxyz4gzqpgHx
1bGCu6CWb709vfZGQvrw08LmAiGs6NiXiBKgN6/f5KL+T0DjXt1sOQtiu04q0k5E
aRDAMKQ4eLcTKED45DPjRbH7w2Ty/UlR3u+ty5+SGExmNXq/4Fd915CoKVtu2io4
DaZB9PBYWux1df6AU9TzJh9fpDkdfgimwll3oEiUlbh5wwJUmsE6c8tV/uk63+vC
e/S/A7Od4W3XzHOrVMoZXGcWTqhVAxobKlu4ghg6Oz2+r4sjYoR4yq6WJ2d7Edde
AR0JARGTojG8StVydLDSROo7/FUOWNWN54dX4kW9yR/l9UF+cu+4ID0VWlcMTCox
4hXsh6eIL+q1VCPgMSwEILezwp+rMXOUl7wMfZW5jRtt4tqsSJc92Sg7C4sDaeua
Sb+Gduf3/2hZGmDPNrcJvi9dTwizOx+jsZDnuSMTo9ZutUJ8rbtIgNoFg9cqJE3T
Lwk6G/nhgJiqXjAemDjArKPa5sWR0bXajRSrB+UJ5O4GnnVJYiwiPx2+Zz7WDR3t
SZRanrzB+WoGAurc+wZA57bc4FoZJfIVDx7DCDCSJNvs4qag5tG5eS/y2Fap+z5v
fuVFW50lxxxre4XMauHniXVjMFRqNQiTm6Z93Wbe/zNrflTwwk9xwVMR+anTZ5dU
elds+tn+tGEZIOiidVZDTp+dcTagrHcpv+iKvDDaaYQ2DipNnxhxwdEfU20IhEsZ
4oq0tpHpl7lWJcERTOeNH1fPpmfcofFXguitJUzGRGEwKXxdEGgiz6bORTvPEMc9
nVN0LQoW4/DNZa5hEZVDn60HF7q2Kf9rPlUJDWP0iNFuEncTn0n1lJmdiWdGchvv
eLJn6TrCBKs/5d9Vz3ocB+Bk8cuCf1QXuSw7H1Ir8OcWcM1S7xT1rADYmUoUZ9LI
0n5xIC34Ac5RYtjfngJ9PuAdjhBpkRV98lrSYkLRdlvkftykcaSI0Jc561EXy9L0
x6T/r1qqfTYRo1yKaxeXIysj0Bio6TFP0HVPsucLIDjSRqkCtmQoZot5L8oRRSaO
nojoF/l0JgMEBNp7b1lI+QgSoOgOd6jABRoZvEWQwYHDr1XwONwleBq6RVAgaZkb
EZcrGIT58xfeItDbK308ctJjW9Ac5RA8gFlpWagWojiwz0qFCUjVlkpOZfme79Ve
9eWZA/4pMrXcoebW1XbXorZ9gQeQuOjmnioMFmkFWgljp0paRAOBe9tNDROcrfpf
fdXjaU6j2aN9XcBtCASASG36tFS/bAsxCrP7b5njTFKBrHMQRrCENI0uhzSoN37E
jmrGa64U2EvNC2fEHSpavKZNqtYhzJ02d5iOvOZhbpUDrHIxBu58is2IKlsC6CtC
zBy5jlQ/UltLTGumpgYfCigPl/O+3Owv0guHgyuDVbv1Drbn7RTO+V+pcYwTGRTd
nK7/yz+Kpu3cEPe81fbinoxjKMdQRP2j8ag6B65Vty7hK5ZUyuO9/6HxmJBtSgsk
hbQRGgF7RbkXg8Q1upquMd3xDSSGfEw3gkHIcYukgYM8y/Nv9WKZiveMmSre4Vr8
EU4SydOqOR7myWrCqgQt0LgA2RusJPRPyFyfwrJuUvQ=
`protect END_PROTECTED