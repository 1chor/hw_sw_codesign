-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
zy+PvcSZ8o70Fvg4SrhTHBAxXho5GWaKvLA1IX/ryA1cF7jA/q7l/6bD7h5uLlVT
bV1y3BSTygVJoOH1DkNuo4TocvVeHHERYsOZ4liksm/05koK7tHkmIIxj8Lbp0Og
+1HkJFeuQyJCHC81c2EdCGpCdsn+zWGJDMIQtFMxzCM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 36528)
`protect data_block
WzMXNDZkzMQwQ1xtPjqfGwUjX097lADF7IRolY7Sj+o+mjqcTBLGOkM56/zXI2dv
Q0L6EO+2lk+53Tlk2ELEYZdsE9gOmhHPXkq02gTpNocy0maA8W3rv+BUIWGtdfrZ
vt8MD5+njqHZtXMtT/4bugqFOaPruP5692uHoe4U+fmc9q8Enk4H3cDblaQ3WqdK
WUm7agwFD5dnWGcysvUXgnFp9tMmguz7niDJIB1Uo/wmRgxb1UcFnuPrxmO/cBXv
Hzofrr1gkCWwB6FpVztCaqJfzWXdZ0yB+TrgJnhBGpzpQup+LtXmUY4v9fAgPWxB
xefo7rSxk1nwSQj0QvOBmm/hlAk6/CNHkL8Woy/2tIZHohfFy51l3QHfiyaYsWEw
DquTEJzZPHPNLM4DrNwWCab6pApCNrd+sxMHhxkAv/ozVEs+AJEHBwlv5WgImt6i
smjoDD7srsbYsB1/2cs8aLGSKFVQoGzNEVtSz0GV717UAOlxBr+6Ipij5Exwo2vO
BbFdujdRZLYFiLsC4ZiFWC+bGpgFxgMDAZwEvQmeh3eIUljQFPscScmbwhgV4IeU
18AGK/pQorEH5YQuCEUhe4Tp//r7VuwpkwRZrNuC1N0Wq1H2lV8q6a8oO2Uld2Al
g8zJE6jLm6mz9ByyYvjqbPscdQJjFBZaKSCZxOi+LV/4BNXQKeDuZJKxYNKFa1IE
eTeI5UPCmX9R+cP5CW+x8Lx7RDMbD2dM30uREIr1DI0aS461UoppGEiUBorYRXOq
m0NLSy0Td6cjL811rnYAo9pdC5e0DO3k16LjeDqcmptRDS4zepHPL1sLQQ5GjHz4
kCEi0mZ0SDQTYn36mvB9hVKhDCl3KKrKD85YrDc0+Tc8rUBca3AHOG5HB2zdppYm
JJMG/3Il5zkylUJ/5ywjydNAq9bfPxxn9So9N9U1zYk9rV6DwtNawloGB32/gTfc
0Bg79QdFE0Jm17+7r5W/IypRnPDfjFj/bc8BYa2kKgvm42D8PbAtUhgabrM8iJA3
N9IsIg5xZVrnCkqFMvrYy4iph6VbC7UWjAxJsHQ2cG1uRF/yetV+2CzSeN+6uOr7
xdI8xip7EIHe0ZZRGTfVRu4ysYY9t/HWHJmS3JkSrTrF+Vdb/f+Y45/vkZa0Vwp/
Ck3h2QxjkQ0dD/cSbSd6B6ZgE0q66elPeUgOai8uZZXzxEul4b3MFBsJx0A2oUjZ
/hIPFhK/I8DWQ0ZMD0oOi+85VCe2ILJnVYWuZvUf2Z9H09qo4nLxK9h1OTmya+H+
FvAeXCMlEraFEtGylPeDGQ153CjCQVrPyf0ZWxMFqxCQxynGl58/2ppHPDSfalbz
aMPgmc5OxmogmcwJ8iaHUJWJl9mqeU1IEbF9zs3fBjUpB3J0vlOMmV+rQwqOD59G
U8GvEuiaxaGcvGV8qPUTX3WkV/0P2oaxZFC9GP+YYTbD4gDqG00LyQ9Ji84pcj2A
WxDMg6iiBbg9qHvLzvj640QlTMmY1s5cGAuuiFML4FBzIuG9tvmcLb6QrzC3tLc4
FqSB2Od31ElmM7nAdjvlPKlS4qGT1j8cCehulaVZ3E4VMuDM/4XuI87wYqa/kVmJ
nMaS2rh4QDnPJzHrLxz19sq8BhbmCbTO7Jdugl/qCViwoha/amNomCUHpM9RILBz
A4lXCRBumK/98QVXU5lKXxr06KV6FT13OUjl26rhehBAlzr2mrKntcToci8ihO5f
dPSJnZZftOdzTJ6ecjrJjQBVO9RYix3upA10T7HQmkSq18FzVK5VSwaBOc4WAbs9
3bqD+4p3Xlq/byG3se8jlwhRgR+fu3YEEpadu++AniZK866bGyHhLSbjUaHdKeOG
P47ESO6R7xMeUxM1rUz1qdIErg37terONbHfXsEAe7H8CsMvaPRpvkqyzAwFFKhE
lUThIxKfUDSJGDOeYTiQ1pNZTt0F4iefHKaHSTY12icIVBV0EaMHQ3WvmBu7skA1
SEgqaHkEWlSQPulUspIPDyhQfg3zH21qUOSDrLCub0Lg7wq/HMG6JhKl8eTuIoZG
V/2q1nYudibgqmtMYWvH3Q27cLBGtass2h8m9PaHdzC1vqnizEHfTLRF4TjbjjhQ
dHIluANmG1/YN8zuQWvkw1+Hlr5wpXpqS2jGH3Rio7ZceBaWSw1YUE7WX4AvJWMR
tWIJVRQj9TuZfezrvR3FgR0G3lQzv7c5wMiKulSyJxaHOHwqGncuGZzB17qvSfAd
JpySm3noCeEZUh5Ns568Qr9GE0O46WsMHFxbcVRedAUOrMEveunrdf5rGQ7UmX+R
jsaYz4Y6Z/gUvIr514BkE81SFW+zurWnfkrbSCFRLJHO+Ll+xH9WxGGr3j19kqn5
9qzYdElWlZFovPp7+Uvgt+GR98EKMsKDakAHtnwN5qHOzdvSkEXGlhc1v3fNhjx3
UEMk2fvO1AHFyXNFG7nVS7N7aKVaxwgvnIPTF1kVMxGWIfDnBEIxm7osAqFRRV+b
GLpMHCBkqIDE4NkVQQBHhB1gn5cpEjRSkexgBsMuMu717ay1WuvppQPSlBnUbKBR
3L5NCy20rsub3GH2sxdEuTJIB4EbS4AeBArZ5lzhp9vNsPm55CtuGTzJ7awRVBGg
Y96ehcraW4207wMDiTPQDR8c1KfQhEJY59VK8pwI0WejS143Q4KoZn7GV6bVNq7t
HbkYznKzmCXNt/PiglX67Ts5uM5V5ox3pd9Kqy/bVMGIxv9MokktMrk6tyHneg3G
smI2BTpRRRbtr/I/RwQ1rsznU+W40kTEh1gF3elPm6aAfzrfHl5GXejmt9KWsGdq
KsRawIGuO7k3yTvQeqwb89iiFC/Nk5l58mWqdyMeFR359msFavbSB2PADu8zdoqe
qbDgOFQLkrwoXxukN28VNKcXdtU4okEWDWlLYZjb/48IahW1kS+SF7RftVIFeXnC
FH63laZ2EzB9Co0GL6ofO/zN5oMu4UsU+34uKooX3dKbH/uuGugcszILPgB4FNkD
2wA6T+6ngQjml8IcJwyEF7SL4KMpHHY3a2oZJ+bv7Gi4Ppdow+0HMzOPCyt/w3se
RojZjIaZh6jHfgrJoWzUtTlwTKePQQBCGXiSFEEsTXpfWeqajo+UCaAfQRrQefpJ
5qmtfsI39GC2DoMQaI+sOZWTicf9fEOxHGb3UQtVvvu2rLtisaPojt5MFBEXMk3y
xOhryAYoBo1n4YkkOtBD2P0xyl6EqjDmXfn+DleHR4w00beGCT2gA9pMSSmXKV+K
TYXEothVzLzPTrTXjCfLvgK1s9Du5Ptp03FSSU8iv7rWj6gV2EFbngYlVq8zmRUD
3mGBCOIjjpxSekumNfv4OhdMJedeinXrTLtRKBx34cpypGh2xZLa2WPBOk89Ry6W
Xw4XqkF+nJK0jn3i2YIFhyFwc3mVSjWniR+34JF5v/njrcP+nUUdP+uYGn+RHaMJ
8GdgIXaOtCqrk0oqVTAAZ69UDiPXVSsDKX4u9js12B/DyRDILl322mGphbdPPa0i
XfzlGE78ka/CI161bLcLsvA2zbf1NF/+S/psY1U4cKmsFYoYSNjeBuOyB2vc39iX
/+vaQUs8Q3Esh14gspFSf5iFUcfNLObg2aaZjxG3HXX2bTDWjcvrCA1MPHqQLaHa
cTjeZhrf7LonMr5P9+YDYIt+J+gIFwSjFAayhgSC/+bonNMHyRhybCIl0JpfTbeK
dwRb/u7eNPVB8ZsoUEid5cAA++jMQdTxodtt5SV0MVcqvBYK1zd/hrokmfdL7M7A
3Tb50C+GqvYRBTQLHQjSl3Z9d5qhC+niEzU82k5BMExnQvrGcju1x+PK3C6JkoaK
AZrOfjUateuzAo/bpQiJFr743NXqzTe9OpyW7nwpI6u9Gb9GUbUvC+zrEGR7QO/O
jO2mMyzIFaw4B/tw+OxI3fI2OWQ1L6AyLVlHqK8AuTM4XaaQcHNykIYiMgMEOcu8
n2ECTyP14f7In7DoeEdZY00uos72onpUwig6lJsP89/dkvx8W3aVOvRa0vYNxMsl
9wdDtuFsckr0s+IGuT0cJzREyx+cmywY1S6ytFscdCn4cgOCcTvBcnF1/9AUIp0A
r4OgWwlKCLfLLlbsJH4BTcFKu0YbbIjDZTYG/NnvyWCI+dsWoPr1/3aLvmGKie+8
FqAhpOa1HfHpH5mDJADTHsvPt0Ie1hbhBAaCflQsw8eFEkaU05pPTnxVzFJxA0zW
z2+6cRzm1wsvjwU6r02m4cdBAAos6WZ3pagjjIUDuodEmWZPTZM8LwyJ6EOVqzmd
6sBXiTGUhTUXBq4YjixESl1LuGS5BQ/N/fdRvXggKuKWdLUjhNUwytcbCzyt46ul
isUMTYgIZCTNEa5ysnlwXTzLyIbH/qF0j5Y0PJMe+93myq1YJi20G9/omQA96Mo8
TPlYZePKvLJSbl2U7j/XlnDUtVFHYmQZF0TauSO9kGOtTjnLAlDhMD0T3LSx3Lsq
g/uJ6pw04tOYbZFQUhUkjjWUMzeQjF2VNZa8x+zeNVzXuh4xGU4HISuH9L0iM3/t
3TgruzDBV76guU7VJcy6h/9wQBe1s8+p+npkKgue7VHIsFj6m+5wKR2HTzlSoWth
5pSpWvlbN0YTD5I/AAPI5QBqTFiSZ5jWYAfMKd8U89uoQWjd1P4BNC8Mnl/F6ZxF
V61M/TS2SPq3e0u9TFW7mTkMgtoXo7W2z5i26DxVspf5vI31q/KQXjC5DhlFPJWH
739TjLrP64UCwMCOsi+ALF3e2dT3DpM/AZaVbCyyLYOebiKVtVQYypJk6WP0y3Fo
6Ettt7OY/gWl1vjvQWMaRMyBaK+wusE6ii2Fpz3xg2Es2b5t9fZDtsFy7vtOIHDa
Qq5shOacPV4fgj+BfHA4nvY/nKWDL3XgmCH0/tDg8jZBQLHucwdfo0VKj/c2nDxO
e9WGYlx3Wd4MKfWehQYYbJdMhkF3zl/0RtZG4ewwSV2DVc75jpO3+T+nY950Y9pd
3KL1Etg2YCktcjWr3CB9OVIvv0pADECs/9iG8ONRHa5PjzcU+CGsONRyPEzm5F02
omlEzLrfM3z3B5J/1MqarT74tTCUx6XclrV2+dlRU7X3iQB8feWm9Njte1c/HE9w
iZV2UAYVwF+r2ymM/ySZtrNZ0nKek0Erj2y246d36KnozSF90tl9VlpaFyEp96nc
aah+o/g7eY5RQgOzZkhmB6DBTebOT6mGyW4HdoR2tUJrEKQbLogkO/+648EPYNuV
WFT/zCS6fDGshK0FNWEOa7tW3C4dwCD2R73kLZgMZhgFTzFE+dgBIPSvl6+R8DVe
TIRfGhMiaKCoUa34GBpfyYWSudYQSaOUgeaf45h58MiZtMZN3c0tRQFpqD2lDQ+M
+nIF3vetuE3qlvn1625x3WcOAMob2M4CrG1VEwqXBAmHoue9kDzvdEX0KMyqgJJX
Cfqy8YfqD8shSQ9DgbYKWXJFB+BYh504/Ql5ChrRXXTKxWe0i61yA7r/t4SAa+oq
R8U3qRRq/iNS2Mjh0rTCbPxpanknMCq8kqQiRWFSa5E1o8AikFteFA1ZE1KspZxP
FGF1Mgi1nQFBfgDup7YOz40qAFcU59gcDgn/tU52zJaKJpuKTQiCDdMT2GS6Ctze
qisqlpCAdqCcb/IoTn4fpMjbEb0RrF/8zA59ulmy4K+D/rCEHOJz4RHIRkeTrfao
JneTuN+4pzEhik6cDUIGfCVsAlOg1HLhuodfQfLsDNL301/yDPuP6CvDqq0NFFAN
bHhNiBApRUmuuk0pPdzIp0ziYNW+cGO4xRRAxxAw88PO9rV8qqnK4OuC3G5nTpUB
48a8UVALOMk8OtnFI/+6YYqK57ikVdm3Jznwml+sNdt2hWtTC4Zr3Em73WTDvI7w
+1CNiX3XWm9eRPPq0Wlb7LHt7hBjk2DOHgVxyigZPU4l10XwlQnFykklBWYV/jF9
n6j3LhVHOoIjzuySE9ARgJfauXnDk//8X1y50ruwxHzUt6BDu+QSaAu3SA//x6aB
vxPeJ0rjNHQBvvv1eKPWCrJOWj39Is5et6zzy1yHREg+cEIPw1BZ/Y0AHl5Kz9uS
4UR5CRwVA8FxtRmzsQYpER3FF9EKonCVGLNkTpRzdI/4hTJxR1p40U6eSR7ViyMa
Hs4lxF3gludS9DPShodOJY6vc1GrgxaTrt6O4Fm2BQUg7Q0dnP3RcYCoSVKpXgZq
6RKit/nZCt+ITXNg+1Ha9L3Q+6k7ZJz6Td+Jqv6+yQ3JBGnawph5A6iBQsCYXPpH
wtDX2a/27uChymz1SgXbJLQ1uij6Vf6c/GQhSbVQ2aQRAoOzt7tbJkNK7fzlflnJ
pxIi9NM6PNwxHkjxQpwK+u+2tkHM6b50KkgJfQ1m4xZPqafYpC98taROThqyDbLc
rYbqlFN2jf1JHng7ku59Q/GC3vaUTeXhz6e2MNAH4cCLGOBArkkMkEGEOaJDGMvN
UiyvTd09v7HkBTG+mqdcH75r+iWObXB6pC9PzMI+t9widAyhp0Q3L11p0I2l8l8t
B1Xs9EgjDvl7j7Ue/axV2CKEFMpWlS2lQXCWe9lV9KryXZw/PZ5KUMhqQH/6tF4t
K/oR87o2w3rsqxrqRwn+dgTsmkcW1B0LVRzHRve1kbqbI2SQeGDhYhuAUhLAiVn5
34Kcrit33IDthNReH9tKl6nlQ6uwkkz34FW4/HC/4kOWNkOgLlXzDJUJmHy/my1m
BlRoI/dLLtEv1Y0yM0CkuZYxIRq0hvFYi7bRa0DNFgcjVZh8xr+aVJWXpb/mBP9Z
TiCksn0I/Ao2LjekRrTRVpzdn0nzem6I7S21ge9y2fuGT+u2tJcAsOneBV8HMNA0
k+Zz8DiRaz2ym1KMOGocnftDJbCCbCKKhYTuU6olXlxFnUj0Y0pbc3gLtIdMsopK
Q6J572fm5iZ878zLamrswV+KH9iwZrJFXzI4IC14RlU5pX+JjFm6ElyL6kI+Q6aR
0SRrDs7bHYkacpLAyW9RsUTv735fa0b8iQAU+dsEN6uhM5vaX4nenb80BXsJhyBw
PI+nNZetZsL3nXJqYG4TWYNFAO538Oo0oZCKrf5wT5v4pKL+zNkm5vzHRIVNyMKr
WcHOV1uJKdQBX8TCFLXHDAojfLRvyuOjZYQbJWM3p427AEktwizT6GPw7jJQUy6/
2X8NfmjJrip+iSKVNSKLr9/h1JLfPPbyAgm1hiFVvaSecQNhyHCZZdT/PQhUSqiF
ra2mA8KzZYvr1sl29I28hr95QJ3x1vty9LmoeutrtqXcmFr1Aa9qkG0y3DYYkE4T
3/tC+Fa2mmSTV0DzQIZnDDJYekNcXUTJO+C22p8fFpzoJ9cU/i8PUxv0y8H77uEK
72xkl53d6OKmRnbiEyUqKUvYI9oPceeXyywR/ND3VhzC7O7o7idUcjHofT+SwxEe
PaQMbOsxKtRONpem4wAoVQdymxsbnlLxm2m9TLWuh3Zvy1Dw/JvQpXGOe/DX8iMT
g/jXfwOgp/G/FVsSE9bIANp3CzEtJHruiJ9ZpbE6MZHmdXLNAscY3NnVoTRb/Xcd
xMZ6x0RSQpBxQOKzx5YiS6U8H/T+YUUkYX3tvrakZiZpvKqMPqQsMq9bZc2N2q1p
YyO0hNHo1zPAtYE5cVhs9F31mppukQWVDsFWk0FGlmfrsI1GtrTZ1nGU6sgajckn
uC83ue4hAcoes+mUib7pymXflgr23EkbF1QDKR4Ih5d8rvfLAtyczMp1uX5k7vyT
TvQAB+fWxkAwFJXFY26vecegUVDh+Rwak217siDZzA92bPEpwxMAh7sB1aWTleGr
dUvZq+kBT9s+Rt7lyRFZAkjR7tssn+SmpL6vMzenJK7FRIwtVtA33kn1nXDfXNPp
XeIMq7Q3fPbDE8e8daC+Yx+GQF1wxf4xig8BrwU/SMRZLc7XblWCXlZx0tMzyoID
u4O4TZKD2gpvxhN7fJSMR49pfxEKZ1hevpNGRqeaQUju366njM8zgeImqNCtWeOg
0t8cXOLLvZHAt5t6TYf03ceCUAMQGqddyQmlmSHub7OWCjFZRrbqkQe45BalajYS
0pf1EZkxj14SkulPrTP3U1ih5taWWuH6BtJTCh0Hp1OoFslcfeNEG6geWPL6q2H2
m+vsLOIyCE/w9Yyrga50poMKJoC5Q+LZ1AZz/0oScvw8/ZvqSyco4Rpde5CTM4v5
2/wNKJuomm3xZR128DrAwgEQgaZjcaioot/KVR2MhDK5LSq+YvktIV6G79h3g+NU
fi4Ro3g9cjPSya2Nd9ZcBtUjHONuPXXd4YqhC/xWgw7Ph9P0EIXoT/Tr3gP0m3Zm
ytlXiHeCxgXj5Dz04MtWYmzUFY6xzB/pe0/Eh4MejYXQHv2k98NJerWFWZkQMCQr
HOtowHkCNcL4t4aYU1YrUZXJQJ3DW/TfzTcfNKmmV0SLWQp6ERp2qiafj9MVnQev
tD8AfuViloCOOT9tVvSdHB/egdpFxu6bks8iEhlWon0tOMNA5dq2U5oKXe3AG1IK
R+vh/xvpp6YM+DSgcta1hajU+aBr98a/aeiCGTIFYArv089LLRvLfrSqRjh55AZf
E/SdHrBf0YDQaIePYCCW78Y9c+U6noehLAeYowbvl8O43i1nkrl/8Ei5azRSGbsn
Ey6ReuELuqT92P2jqPXxT6NHeZwNKlfGb0MSohn3zNVcWIiLk2tndQ5VTuTUlY9D
kZE2HCdkg6vn3xGFbTpBYX5jZVEMhum/q3KfZhzy4l9dyG6impbDPMIkIt+iqeFd
6sTLP7b8Vqu7XHBSU5xZ+LmkHTgPHmgqaG2HmF9kiiTBLO8PSxxhYkBNw0oO2kBY
HYnf0SH//jP4zzhWLsltL84My20uVhq+Px0TCF3B0GJN7SEgHU7+XtB9iQ91x8k2
ifSTEUjoNG8QY6TkZMH/j92IJawZR3wjyHBWOR03GzfoAsqYgNjOCTolUyOWsfqW
DdUDpuorYLsHlg3UL8K8O56EecFTigcr0xQ9r4UGPUXNaS0iwpVyt3qPJuAf8tfZ
8gR22FjDYpxUBD6zg/UOT1uxhsF6Kq4Uslo6pTJNprSODTDj1AbTO9nXYH79XFya
pN4X7V1nAwaZFTZs9jYaXYjzX/Hz0T5FuplzMKzzwrTuwCGnjPdfyqg5f6G3CtF6
3xk6v+wN7ASapzwvOIbYmZlTVgdB5kmUp8lWwSUM08tvi+1XXhiDQuUmJhCkOCXd
j9vO5BNJnrZYOV+nd9skZzuv/O1EVZifdJRAztnjWejft41iJPlAtm188ocm04hC
QMpVEznFqTTAAjvldr06ucM0RRm9wCFEmdJBx8PO351Xx/z1gtQ36yoNBxhArPB6
bDeSfZ26cBShIT5jdAPypgAmqvgRndKCBLn6rd4lhTq22PN9BqglkpEv87TULy0k
Jq1+ZRLkfnDhwjqKopVimg5vD/Wf3+uRONnN1oHlZgEKST9NYJlB8kfpZaBQFwpm
y43s/b8iSWaZ0Auvpw7okAKMG1Ojcn/8Lf0OLA/tfsLIGC/vFzbSYJLmwrD/Kgxf
EyNUDSOVqgjojfDm66Zz38xgSZKdTf3vV5nbfx+KkDzc3+P7dpNIiTFncReG3Q/y
y8x7ZMGpFliecVkYOuAIMAMtuNOSJ2GMzWWhoQoA3Gbn6sXxzPMCuT/XvMFmYdCF
eSOhVjWxcxiASFeeFWAZe7l5SMCByeeebZK/gniNmUoWE2OBNhZv5lFExYT1M3K6
eIFOCRzkx830Bo7EWet1tA8MR51Y8KimCX4vHXO9fHrIvF624iOJ692ccWRxBbWL
a0MhWRJw381f1RlKC1cAmfqGsmU45N7bynVW6hmtXFTnoTLMjVdqGGpfz+q3TO27
dM79EcoPx97sAYPv8iaSAzSIN794lmsMYgnmjK6FMEgyJo7sT3uyZxCnRWq3B0VK
9DIBcS2g2c+ZdVvvIJ6ad6//ykdoE0E4o8vLrJ3JP6cg934m+/NqA+5S1bXP7hbH
SZFB1JgHMNlktEQkcaKe0pFvktpsB18Ap3m4Nv4ogXhjAcgXbLq+h4axh62zyRRo
EIvRPmaSKfXdfceb4OoxEKqEtQDCk0cGfEhLuRaFrvSDaMNyKa/IRR6ir7TDgU42
2qijd8qblaRVhJiU6dVEwr2Y44BqA01VWJGtscr1n7Hkf3jc7as3b5zi7J2fPtua
Xe5WpCaoJlFnBFHrtiQc2E7gzPBSaWEUg401R++1C+cYSUY2PaWTBD0yMNv0vXoS
WnkAhIU0PpyQ/gXFo24WIdbP3BY3S77NF9328Sup+OX8wm6S55ruxWu2ydkyA1E7
1xbQTKaja74bPOYQ3ALdKZ/erAGeFBD6W6+8ZcXPX4ELvfTry4Er41Fs6ZWPQZR2
xJWGMY3Yp1DsFZNZpq66ioNwdEMO4Fk7uJgOlQSm4kBMZVHPp1uJwM0ia1sFPSHI
k7RpGdMO8RKgcms9y9dIT3LL+KDHQpz3dTEtI98Tobt/dvj4ZpDNeoP6woCfepPs
DABPa4DJRsng6AMXOHwDjPQNPZ/erGz4NvhpsEKj8P7I8gYaxBVx+DRW7tRtmFoM
qGy01hpObgA0CJM+qUqege9NuYnqE477nDW0mtplfrOkFhs8YkW9No42epou6+HT
QSM6RIASXcDWHf9DHI9GIZavg6VZN0fqaSwhwoU3G6F3gdsckR0l4ucbbxMOQRUY
iOpTNqDYEk51jkwnUNe+oRkz5FAW394COt9yAD7Nq0A8ifGuQr0TeKOOR2mMlBJh
W5TyxMqyAseisyHVkAr73QL1Lsivk1x0fnOcuBTKwejhFQMTBY33xWiQdwE6xdM9
eb8Crey/R0rYj7K7eS6VKb7b2F6Dnnf90K+Q+DybUHo8+hvBKdRIziihtFGV3fZW
7h3avBGBXIWYDEQNPGvOvPcUbYxpiVzxb5DDzhAamhfuWhu07soDVboi8en8ebsh
lLZxx0zXjvkIATI6fNPyQTD/gO+BM5uoibuJTToynxZIcSa9jMwV9DYzqr+e15Sn
0a0oOWw2/Y+gXofhMw+Seg7CV4TXh76WbFiZhLH+iXU/+2UhUXfOgL+dbnacSpO3
Zz0RoPAizxqqNngI9ktNksCVi9Y5cX8pwoZ8AatEuGN99LSVpZeJbLDmiN+VJcA/
tSYJtOGyiCj84SGxQNXVoJAYQpCPn6iyMvAe+RZK2iPFkkpSvMb9pOsvxxrQZr3a
h3fmU69Nntj/qS3C+3lFjpPKuua9M5pBZ6KsrTg4OqSjHm7UOX52IAd8YgVdYbgA
cUt66q4LbQvh0wbCVwjyRItFa2SZyHVYZyVYs5bVflv+EmIshUIEU1squ+zMqz5K
3isG7ZjSdSqJIi5EnAfMF2Xh+VuLgvHS6oyjM9OeYdlrxJHuTQoya48eFvhTjE93
SjkFupXRfKpbTGTtqGw4XbgT6Tw5rIRaaAHQFvwWG7i3s8ZsKmEh5uQ+nDAPF7Ed
mtEkJFmJIllbAtC9A4ioJ052w15pZX6JEKWzW9sJmqiqXVFqjdmdB7+qhsBxZdcC
QopEQuOmIyare7ye7iIr+LzyNn4BO5gfV91L6ab4DrouAFeFlTcGjljEizwFWCiS
3cU2KZS4nz3YJdGtoZsqd63HtOm4fP47kiieKjEYTvkC73aN51sDejP65BP8ck0J
yq8ufQG7YbrmRcAPM4Asx5ZkAZSf5ju2akJ+NEAOwyEf1ojbhvwXabZQ34vJjcSj
4xnj/03+fP10m6nuUF19CYPekhD0k//yh+YVQtR2KQj+ZWGY1+9YBp8A+aBSRbC1
2jh71eGaa9gvCqGkA2ugB8VQ4eMtS+LtbfRGhFzec2CY2r9JzWwsBCSMZBx0+Sb5
rmlw30ZwrnrZvZsP65QWFrV+UXZhObWZA/VASrtx7DCIxImd53/Kr8gQT+EMrOs0
Kj3srYb6DJ2Mtt0PbGkfnzVu6YuZUXGi4zIh/S5X7MJY5fnHbfg5xsxkiH6zBzba
6ACO6b/l1Dl3SKF5v5s9OLHnjblqWZJKkwBgC3Oe3Euy3cv2DBoa+OZATptMVLNY
bONPZYt0wvRAy1Hdrb0YYQzzEvSfDXA+HYmqMS8VDqqhBv6CbW89pCoM3fgj/PJw
Bm/Gb6naZgTqQiTQatxcgMq25DbA8hXow+9I+Jm56nknrt9bmeF2DIhIoX98Asva
CF/h9L98mZ19uHuq95DzxdZHOsY+Hcc0M4cSvnY+hY1jG6GLVhJi/K5Hn1SrbK+a
bK4TLJzdtyRgHdRwjeIXFDXOanRGOtnpjCTAdF/3vM8a+DloSeYwf61ndLb3mIdw
xpX/9vbcaM5X4cWvdz9i6sEgClVxlea1Ec/C4JGj4hhKh/My0f7371gb03TkHH3h
mY3RAapxKVojUldWd5gZ0/w7l4QSmw7m/qjMqE7GS1xchrUOK403H/GpQsv/IbkS
01Fkq1cRvzimJ5prNUQ4IkqTCyok3q3xH2WUO47eJ6iIsupfEH4CjB7V6SVIHPNI
Q/K5HKUx/5XAPD15mIAZIIPUqWMcVLCBtA/tlsqmBMndxGMeTxgwmF5XWgKy4qVS
4ycmgVtiUSlxYYYAl9z635bFVE9vqIvK0kKUeBNvnr7sBrXa6s+FipPMOcqAIfwI
gzP/B1oS/LjYsJ0IGdTcXou39R1AMonxmDHGXOo6tUw2iUktc6eJLsUHsBES8Lxn
PX2K0wfwWZ9happNPlEV0SAOQ38DcHGVy8d1d2kLFOcY5QuvUDjD1TqrKx10HL2X
MDJr08NmwjdxEs5CaZFpn7REX4pco7+f70c7QQS8e/B10ACzzs/yZ/xeQ7z3fh/G
rilNR/L6jiF9HZiuejRsM+xuvXunUPU3YsUkECIBd/eVg+GNN/RvGhSOhHzasIYE
wx5xQhb2vyf6E06Ox519P2AbrGMJyta34gYQrWwdgfPf59g/wZ+NZE7W9BfgcXTr
MVZXvLcYVd5dHRLloKKRRwyWW32+EtcyRl7FEW3+3wloxrMWGuBF/IVFYfbBFxua
HG8tpr0JcKnNh8MGIYERiEOA+3NPNDLZtAcqSve3Pi3Q4DqfJBi7RZit0aOev8hc
dWxmP3xCB+nwou+y/Z5ncVWRSkWSg2kJhqbTwIthBAy3N602X1kiPK7N2NDnjv/Y
zN//gUEZqydV5PRiV3ip9pQTIploz6sjuFrg1j4xnuQKqxAlz1cqKcrFINDZ7thX
EZdw8EB9AcU/U3xeDOQa7Uflhzvyt0gl/mQoQv1tm5ftyfLxZvep2KVAlfdSVCFg
tn2MwGpaMHlO2JUR+Lz1o9s6s3hgUh1WMAnW6T97dmAqVZoRBlKgJOZsPtP2p68f
oo6QmloTRR95LzJimiRKE3doVU6brWQVC54gWP0bq9Zy6qBH7ZQP7ZIlfd1Xtnyz
GZBp+ZH/j9LB5VUeoQn++/y1N3cNJCduauUp+2cUfJekcYEoaL4gcKNKNoF/+0hO
f8t3VqGi7vzVY4FfAjbtR7zyInj63VvijSDV4IFh2+a4sYLWh8eZeb809P/UU5si
a+8JHVQOKDf//zEncmDcos1s/1r2MO8UXCZEggJs0YLf23b4KGn0OJrvYqbKT9d+
YKG9+dFH7aD53olUFo9567hhSOcwzVJjMQTblhvm63VfDr4CfR8IAVx0197ptdWN
eUe5wqPYsn/7W4sNAjQUfSTG8fVj5w0cZUjkJFsuHR8ve61D03UmvILQcKKyz88f
lprGwuNAl8O5IdeY99ySYprNK/I/KGI1wFaZK6F8QoBRglA0UfayQ/cruhotEu6F
uNMxJqAYhCJk17Yxfw5rT8kFP7ccQh4XOogedqFDw5mFhT8tRDpjQqrNoi08I8ai
5mLzvpnmD8Yt3q3yWQdZ+I76gMJzyEbumPl6MzpRUEhJaPJzbnWbR+aV+2qHdvjU
Coln84g7zJv10EkDbuRQNx7DVvKBkXePR+rtUyn/OsHohx6FVbjiio3pllGsJz+U
ZMTqiA+uYXm09uWeSkQ+A57TOe+e/ccL4EgQY5sadycyctX6pJSG8I8X/fNO30g2
A3/mnsBSeVY0oZk2yApdt2Q+CoxwEebSTlxa1GQB1DXM5zf16amW4x9kzBgBTiH0
nP3lB509B1qLIa2nn2uaiCqnshLbf9J6UMynX23xpfGFtSkhkbMPmn/VUPhIiM1j
vtH79d48+T0KErtKn1gNXUwJby0hC8iWY8wSSfhyrkvHsV9Ytu4ws01VZhxiP9lp
Z+MderOa0RuULu5jAj2fq8pxOMJimmDUUefelvT8ZIx0ykzz1mickMxULHTpRvkn
3aDZKa2HJrl335wdU/qYhZ7wWBzzRfirDNnpbSWUaoYChV22yFFEg6WATmDzCP+N
q9k2kN6cAEdBBy9+Y8mhNzct0DT6jq0U3dA+LVTs+0U1mXDkWpoW6RFh7mjoUhR1
OXV+YoFvEfvj0NPJdbRpbe3FL9umFI8UN/M1Ff5MHzXAIcd0B/YpZ/U4yoj6Vba2
Hm73GJqFXxFeyipVdx3epy3rThpKiO4OXmXNarUSgblGNbNxRkAe3gfLKDoGTTfx
Ke64+jn9D8PGaHtJ5JgkJGCOSLx22KZN/zj6sPf0jEQFNAxzsHLWPDLcnzpgcKg4
0gjMPG6KQm4capwovOGhcT/5VVg7Xr4tBMLwSrh9Xoi4gk7zwBE5o5bVYbXN6g/j
hjblhEhqCWg4jBhhLqMSgK/qMJUeJ4Ia0BxmL4OXtaUb4dQL3RQhpPHwkofRFFha
VBgKV0l/rqya7kZxXWAASHMoYnTn4u2x8MU1LmhS3jGR4M64DYWiY3Q8bNaoBNIs
ZbJyHcvU38y78cxPoNDbZgs4Fi/96bqg0fcLL5kjbxyt5CWZFg7ya6WrkEyXWdqN
epicZw0WB+0hay3XoU2tIvsBFQHTP82jF7xfEsXlkHzsTxHdRFCA06Woqf5/DWiA
317jUZtHEdch6jZgL7eVRNQAbhEmUMW+tA311VdkcHT9fHD9ucBaEO52ZeHJ82V7
XnNXn/2stzp7zce9pjWQ58mX+DCdm4AKO/tiXu63P20K+6rrlDPtHpUP2+Ukx4Fj
40XyWAex2dNFd88/VWp0XaL50XCwbgSveXd9NYVfxTbqRIzMKzUgw3AmanKXuJP5
Fsxc/aUZDnAkHmngh6XzcoannAL3Kj6saAgVBFDu+ig96CFuviJ/qmSfj/HMO8QY
rYHfIysWfsdI1LGp70QAsvrS8tudSLXvfsdml252mvln1ZRXsXCnE/tr/TMc8w6h
hK9H1qHBYHlk4zxoUfjuJeIt+E1eO6JU//TrkZEwE+A2Q4A3iEW5xVPqB0i4EtaZ
ymeCCfWPuI7/Vo7lyYu2XY3eA82K04csLn3FNQPzFUwswzkNqMSG3jF+svVrfM6W
cXUYrC3ry3G3rz8aX/Y/Ag8MybC9RZMAKCyvnEd1o/G3/Da2wi+1HIMBoTwnhy3O
HXbvsRVr7PaHfFFBES6VIyP+uHeWAwG7LwcHq6mzLHLdzT4ANGy5/eNpMkQ7XpDw
p93slTIEvt0CD55aTMFGHzPH75/9AGN98Iyq+rkjYEx0ZuPetKhrjQqj5dvAxAKD
0jwyweh5Q21/rYlN/tZwF+ezqFDDu+DKRk3S7P/LHQK8p+TgofHAF6nI0py4MsVz
NcdCmOjIUh55N/ALJzgBhvNxxyG6t36vLebU56pWSWR2twnNzOY6XsRldBtGyHi2
HB6zUAA5RpTNPHwUO+ODOS6VBFfUxZS5DhrFrZzcGo4k5B9IjNcxyKEKQxlWI8cY
RDMedZSZR4rOSE4koCJ/zygyr/RjbwQinkoWoZneUVEywq1Nqz6bPD3iOIQ6qVa8
l5bSAw0hRQI+GtQXOb8RON1+rLR0PwhOOqRIgY5vFmGL0t4V6M/6CrJu8CWCkYP/
PRj4tGg9gMBNo+Ryl6ekNpD+pCUul8XbzxALXWRG7PCvW+joU+GxWocW2lNwk+a/
PqVZPlW7qclcenPoAtreIXwDWsuwTqc6K4eRor+8lRiNrAW9wKDbVw8otrb2i1rl
1aliJ0EsJIKglIPwwZ2PFH4bK2l2iuFIQTwEVxQImqWKWIkQMcVhmIxnvgbrZ2Vg
Uyqw1NGrd1sZLBTR8WKYIpH/92zY2TnzOFRyoCHXiUtxMy57nBR+Iq3iZz/Om6fB
taga81sE7+5DLdNPCxtw76na26nBSfPTszgVg1wuxSL+E2vn+Vj554Fx8w0OSgg9
zb+rFKVbCywKy8G85rLjuxWB+dE8oM2tscLeWh0rQSvJWRqOd9X2byUvC2aDUPYY
Sc1E1tHK2vsAQIacSxpWEV1CF6WrAOmHiz+/lYmBKLr2XISA9e1eVzMDUl/4TQfm
eFay9qH1UgG2dCDqtSeNBKGvmJPtpMJ6GZcupcvP9xsL/s+XmEh6QqzKQilvb+Zd
JEDPgFsnspiRHntBnfVotPwxXJkZcHY66SZTj0BaSwL3YJkuPGsc4BEgPz98/Pzy
BZcq8mte+fjzERaclo9vfH/KnTOJoq88rdAr3b0qm7URRdWmBcx866cHRDqNxNML
AXp1ZK04KPoKaeFhAa6vI5HLohMIGpxfZmm7tUDk2TNKRTiGmkoS8PkL9NQOeQZN
eziuIAenkgM2aY6oKLPaUwQPvqgC3K63XPwCj0MqfLa79TUqm7zsV1Qiklw0J/7E
s1OdQ5sdQBFOGybS8+XDwmiXSA9caQZFIf0+oTU2k1pDDTISANu/7X66CD7EywHj
JLPaRcgzCz+drwsgBpq5Cj7anVYVPSiQbjG9AjP3dbMEKUgfgPI3fONZcLixxGgt
edGM+8A1230BzdrFpCXc2HN2Ht7nvCnzLY8ujr9p1d8V6bJ9hR7QcbaBlI8q3wR+
YWRayvdlD2V0t2gk/2fIjdhL/SJwcikpIsjxEZNg1V+NC9aqYbo+oQqVJEkVnbnN
MvnnLA/iJ1okkQExoIB0vWYmugkP7RLJS+0kB342/4HCFFT6c3M0D+ylUsPgYd6v
roRpxQ8tXTYOhRFxQ1igsIaaAGS9e+3pt+elkU/SIXMT3HiQOPjfr7ObEgUl9+AP
fhVBpPCU2V2z4Jd5QCMXdUlNM68JdgsOL/rgv8/CgJT+3SU7MKA4iveeLB5AaDna
QkUe7RuIIfz/a5rBr3mqRWK2O1QILAlqgF7g0AA5a0sphY6tVXM5QM9UOphQ2/4B
TGsuI2AoojFYELDwepRlD8oVuW4zHaFeRvzaexefXBZhCA81A/LGeBaECEh9n8tc
+dBPbevRBh1mbVLetYwtCaR0cCuTdiB8sxUZdBRSTxD6NOba6OjG8NxeTP33rYDV
+eyyyPPaJGgE9ZoloyEzcm1e0mKNjOecjGmzHbogXsKYSFbRPVEZwU6gbbRsc09T
6k2UKTRniwiT6oKSAg6QxoghV+tkv1lyWykMQ6EkNJKK3NbLqO1oqB9TV/e0Dtp7
hDK0tG83alffhu/J4WjG9C0/8546mAUUzutkoCN1u/k8R4Ywu5mCr3/y1+NHy6kq
zDoGAXwWUU3PCsfB7jLHohVGTUpGzo9ojUlyHg9vbJla5AQIAPjMAKRGfYWINqd7
KZjuskBiRbndnI4WAasXqV5Ggvs/nBrqydOapncIpazzDZ5Bo1CoptpV9gX4rPOi
XGo5XudINdENbCa5OB3KcHGiwdRmBJaIDNn9yxvljt/KzAGQ6eHdxAcJUGrrT9mt
MumgIv5A8gNEApS0/uSgiwg2W/I9tS1yu2agmHnQoga4VE+UliRiS5K3oUKik9W6
bAk7QerhAq8vORO+h24zGQrGyE0b6+CXcMdheOHxZBYaTJdACXWRG9My8ft2R919
0cj1U6EjNm9tvq6mTOWyFYOBwNzNAvrxVHqsOHhyVm92x3vDNOk1zlccP5QBIrCS
GBgNqki/kqBse9JyFYot2OnKeLSaZUSVMtNdbk3+R1iPnXY3CqWJB7dbCVEpK2jp
ddKxq3sn40+yx2luXrl3RygvOejtCr5mhj0Eirf/Pnbzpc2HMw3RSlDqLfNKv1sO
pO6SX82AlhH0lX0Xj6lImnLnPxgHRBiplu7M1bijfJ5zB7Ln3oUi3RpfJolYm3ao
aRXw/AzuUHZY8tzX7sEaWjHYgDgvMnR2V/3mOFZJM9gASYm5i95MhUNH5YDlvGeC
RI02QLRppMJMdulzmJgNkFY1bvJKBHBNMQKqEyMZpVyS2gQ0OHHgFkMnHq4JLLOq
wHW3gA53WZRDHBrz0VIkoXEsd4TMurBWYpILEOybPJTYhXQdUtjWqE0XBxCTUOs8
XwRmZYoZql6vCvJ+RJbd40ZX659U+eFZsTm1urFgQQdaaUU0ABMf+LncnGemBqL5
SJfCt2xDwYsKHU2BNAC7n4sIs/SaEHQN6GM2KUYQPp6z9xerQq+KhPScUY7pXUDN
fG4sw9y/gEXKv6kxfZajPVvRDuk6IazRSlXqmQouH+u8VqcVuRh54zKC0HJ/Hkep
l94XJSI94z9jVkaXJ3Lop16O/MvHzItqGjEE/6COOPGahopGH9EdQQzoHazNn9X0
fzFJx+PBMrezobXWL29bXoinxpIAI98gL1vEGPoQb/Z2vD+C58Hia2qEvHrrQoEy
pW4jnMeAf0r6vKmKnlbbKdfIIY8XbMq3iF18UA3zl4StmwcQasB6ygHKhLyW+WiK
DsVUuTRCVgTUmkSE1TH0/HU/Dsq3zBJSRB+ejfWKuA6kBsz93VSqQVCSbb5xIUwU
KC1+/V1BvQA2raWb74h/ep9Qn7j9n252O7QVBaEUlXpJhHnsfhFkElHcbcj5VV1N
NqomFqYm9qqbgtAZJcibMelorBvRuAc5pzNl4Tx5ov+ARp0eQr6DYqLV2SEDSQmO
Y7IFyOU6assQqCpwfKAsO1alz48wq4gsBX7HZr7PellepCVEB7EKac1hngiaHKR/
/Ge1lLSDoKlm544KmU9CQoqLNncTEjyTrfmDF/U0xG5qMjZyxgu8A+h11xBlLQqW
29fKXKsJ1kOAggRa1z3OOSl4rNk3DenZi3m4Lj1NPDnzyLwhFLqBkGst52fRH8ej
BS/8CO9usBnubeqCfVqJBSqdx8/6AnxGAE7VTSJbdkC+vELGx9awq1prYKP8DvsP
UHGSk68F/k/padaC5LO1ePEpi0asGgxO6lBE8Ms7O3o0EyoJ4AX+RQs/DnzDydBn
GGb0aux8ipY/BDe+oemdEj/JGmxlZfDSSOWqGgT7XYbfgyWhB/SRS7+/RsykKikO
abEApX/E+SVdSzau+LRPDdZxGbz9p2CozmXDaZOboEaPZPoKhZaJquDC3+GUN8iC
z1krFbd823XnYvL/QYfkG5GvnNrem+B+7Vl9dWfNzzQQ/QBw7ejctiMx/SAm8OdB
4MbQpjoU3OYj182KLSEqEZe2SFgdec6dMMyogoxPmYHpUWRQTsDHh8xpOcphoE59
HhyZAPYh9U0VgSQtiyXzK4bd33vfycChPebeJuRFDGcNk3StbS3crN1HHs4nlxm6
pgrXp/fnDpY1obBKf1KYyeMDASo4TWaa9ZEMZenhyc+IxsRdHmXrluyh2OQvd/+r
U2DPmyJQ4D0x91f4ZZaYE6iGeYc1fpSKKJvUKwGuSBG4nQEn/kpW56J/y+/W9prm
vu+gdsnZEYO9+qCC0gZNjc/j+eijzzTg0ith5Rd/tVjQE+iRxZzUTkX3dA4gNlzN
SQhWCKDhS6nL42hRJcUov7sJuodlj5eaUYrs6LtxYfVQbNEbZcPdxYPk0KD6D+Xd
UCl1XVcH9qjxAqI0+cgcftcCWiAaxvdxRPq2QXwPtlYZfLBZ1QziD1dzno2nQ+Dd
Um8u/jvCJ34X6TFRW1GvbluU+/F9JOwIqwG2fc7AZPGNsvAwcLwhp/RV1FcpfvyW
+FctVpH9JfgpCTUbtRmdYccCBsgYEKNYG9LISuk5tQHF4FTNXnsUZpGOgR3Yi8PT
t9dIS1B3S4CFRDEFF7uxcynvU7k6Kc4p0v8Vc2RVlMflngsrkPzOigcR4MLO+e5Q
TB0aZHTRN4V276bbgRYTdmfVxWesHSsLShECOrriN3Vuh+GEZQpgTDZBuuUxphXf
BxuT6658gy3VuSphD2iUoxrBb8D1HZYQEFvQz/CZRDWPkIJtoPMo85sUv0eE9V5D
feCk+2S9PSvXF6/S3FcbVGi0s5sIn9uaI1Q0r3AQSkIbZwjY/VYoEmj2m+h0oILn
bSWS1JftWKil5yjZToN1hdIRKhL4O5lpvMeg5ohpvM2VCbQ+UW5EmTzMWsv8Shpq
xq3YtIF0Zhql0aJDZuCehHJc7uHSx03sQQfdn2tOBrL6S/XFJ7nlpS1eNI0+IkTB
Gbd2VCHEg4bIGfh3cZnLXZHCh8feyPh7Wa+kygWtoA8acmUiyC2zO838jxRTTXe8
XIY+dVO0bNfznbX5x3yMQ+rgqcZr4yIV438yxz9WpTuntn82hhsg3YWPOM0p70j8
NPTZPFdP1K81FhvWxumGIP6IZjBjNJ4i1VUvifAYiwUL4D1pT51nPMDWY0vJF6TO
r0JcVXveThGXg4wpnDAKP8KKtLa71KWP/9l9DdgH4pZJzxB4fWsLd2mZ71zHWydi
4gGYlnhxCMG0jJ810e3KQDaLH9wUragET5qAJWoISCbsh9DCmMaD/Z1nfZnKhWMP
LI9C2cfb72zUL7w2mNDbwuSkDbUezaPK5AZ0hz8SmFDhls0QVBxlxrjCKAlDfOsG
TecSUpylqUCb3DEg7IwHKTV/rRzaUsdd38EtmfNDOJ/xjU9MYw6rSJpSQsHa8GpK
Te6zgsdvVnzoHLJylDI0vsZ165lb99zSXkkXZSsZNoWy8VAed3XU/W8d71sVGOnI
m34xY7WDSWVVGZjwexyE0z9O+zNNJ5SUs6Wt7zVBAVJs+8WcvOBlZ12uzqdWmofT
/mAXn7guEQeXldwSQh3P475MNKhOZY3F6KGBE9ncIK0EA8jYwN2hjUlkJ0J5smNg
0UnPt2oyqP52C9sYiys2t2zEoySATA3MswyGY/QXqP86Th+yPeQPJ7bUMYnEKgCX
7nVih7crJLC2eS/zHASTG/T9HIQ3diCXkmeJn9/z/q77B434ddBFwB6XRQ2Zj+dR
k8NdITUkwxFSW06vUfg0XKPK119Akthc2qdKyXYVCxIcp2c9H6HF2MqWVA0SdBNI
7R4iwjGoKjP6jGRHN1If007xQSeErPM6hUaP6pHjCUlSTOWgdR0YPFeMOae56TL1
I6izlGa0d2HFH3PdZH+OdFDrcSIOgKfeLKg72Rmw6wDTWfoujMF0NFjAF1An1dUW
Jrr4MMQQGQqWOkzv7S/PEwXGOWqh0nznVWqPF0QsykNxplOy/CQ/uNQn561XIFMT
KKzYjWcaKTON7YklWJ4hrLWhhBChEojl5XvnkPRg7zVo1oDYpm3Jy3N6EcPOkkCF
mN5RumfP0wPT7v0uhKpFSeuj18DWNFjTnMSnCh3RFkkCgi7pBhjJ1UDn3jZow5Ld
ZqMZ3Vr9H/nNyuoIsCxtPbUnjOcxrSM0GiUi62Co/2fi6n7uzXAjHd+4jtXJzSTq
p2a0DTmFRzrzJLGMm5V58eBFakd99k1EmcORY+2lX51bCdno1bINCWDsoMH5QK+G
4dw5waupmxKAYkFe/Sif/6tUoz4HE7/Y6+22PwWZ/iQS70dS0632Bf8Tx8obsoxA
MP5JEJMFf2Jm/Hs9Fc+r7LK1ceR9tmipX3K7KDT/t2pe04n0BK8JUwKCVbvpsCxs
ROTUFf0NYx8i0r9UX7ejwOCrMokZXrja8wjoN8OVtU7kCXv52VT29wetQQ0AxW1z
yNyY0yew5tNWKW7B64lX1qlBrrsHHTfPJ/2E210pGPE66a7KfFrYk+X1d2vPqwQ6
d6PVFy/c+ki0ZqkrlFk2ZaGVkwOypKbSXFaKBDN3jHB8cr30UGkI0DspmSVZiQmA
OH/BQw9DMzYlbpwJ16q3Ym7bewjInxzzejlTmndfNCQYq1LkP/v141DfFDDRplCm
l+X8NlZJl8cqhESiUDjjvg8UOS1dOP6A9Ud7BaWIz8qXP6xA53ClkYKM/mbChgte
ZQVH8RapS0Ph1QqlxRMA01Uw9l/6d6D78G3hgSWKBePEcsMuxtqwUQfozkmuOTst
2sIN7pQYjhdT00p9evi4xfSSINjnOPpBiy1M3qFS3utSz/8uCTayMS9WEWbtT1Fb
gMXeOpZIlCH5/ZRJhRWUCiHMbz1fO9L4spy56yaLxsHI7aSeJhMNCHPN9uZCrf5B
c4v5W+GsLr7C5UIZZkTY/0aKl6KuINhXfovghi82dPPqIc8kG7vY8zIrgXFyKCAt
7C2Hp860FB0e0zJ6hek+gB4T/t2zwxCKW7PHiuQ94x9niPXS0aJTqp+5qrmTSbVE
npEy+h8ZhhL3xFBYn9eTa/KImiyskxhHiSlhflJeT6gBrN3A0gKVLf8TwzM/r31G
uzzyfZhoux54erdh9MGpmBHdBf1hR0Vma8wVPccZtzpdwpEvqzc/UjKfT4E7bj20
XHsddXaGsERGRR/JoRQONpeMxU5x8hLtqRIL2ot6Ho5t1NWeeya1DztBYWPyK2Dt
bgqAAY5vJk/6/CtnRrsiZM8SW3O4w27c8E8Izw6R6sCMWilYpnY/zZjHOPhzdaNQ
jMG6JrwFNZtrLS0AC2ssl32P+ujVkNW8DlKdeHGiWhFRt5zgKutSbF4yejHFies8
6ohp4+bZuwDwXz0sECfYMXoQyedbJzKYULeWHb2wb3I3Iu5xp5Kb0yMFHzRt5rJ5
x3mHf3Bm77dVu6hNJFnyTYhiBhy6ylZaWvhFZhcSz/vOBps5k65ZAQc93QEPPR8D
7VCJ9PXavLsYMiWUn6UdNi9skaJSFE44uPnEqFnQxzXyBCkTG7LXex2Gu1Ah+Osc
gNoIASYYRiDRjndp8roWPXZq5ARPYxFE9YyRTNrlQD1bHWzoESbsn9r34NsyYSpR
9P5RO9qQdE9AO4kWNizkzTjCXQ4n3u1JKWEIbGqWpT706wEPIoJaowXzc67M1IPd
YxIO1AULISri0hx+/Q4cCK9gnIVu40dJnB+WM+epwFJhfaS0HBAA4TSesvIyntLs
l9lYpxF1/PEE+qQzgf0yYE2jvO9odBJQuNPnni4cUdzeCwX8CmgV8s2UAE7+VP+F
yqTBZ/5z6K6bPpTI4r4HSFGSk026eULpXSOETFgD0JA8SrPINWgNqFnDk05nC3jW
yeTwpLoDje4V1H2nYGCvzmCKUlzINsHrR9wwWTcl/bxdr9zAvm4mkcaagXy0kPKG
lW/HGClvhxIkcxqlslZrIHzgPN4JSNVS/CMvMPfIXm6Q6IDLSY0ARD5DVJ7Xi7XD
/wwPxNvvg4/8xpijuSufSij4tyQeUGlC+UA+bErcazexQphzmqpkxu6OOtitCdW3
y5AUUngqlK+Ux/RM7am2BqTBadR3rWwiLsGMDUP+hsxv/ZX61MJx7mjJDSVP6FPZ
hPdb61ufccw+ch5FI/x8OEGYajnaJ+UnEot74MuqC5NUTuZUZsAPRH/UHYoYFpNH
v5DxFgPtb6sLtXvTxuFXrar4iVzA2i+8BEXba2S4Iy4uKif5lsg5t0gam5gSapRO
0UVuDeuFLUWSgfqpANnhNJOqP8VNJglsy2gU5brWIGKJRwQu9laiv3xaDzTGvziy
jOFizENd7Fvlf+V60dVZk4mWqOXJY2d2B65KWnTGyJaFOCPgQB7f0lGZETwFmI7R
G25/wE0ZlFTQlgM46tlkNWFWJM2WjI+tiOmnRlpBOjARbLKKUIXcdxYgs/OHdAWF
wWqj9Ujx/hKK5we0/xjshMrPH99PM6fyUqKEKuDlbWT/S7VZem/T0bsQjRCeX4bM
/WiIl5LYUWQMxCnj7c80lpkw6p0yRqLKU0Z4lRWW2rXADgSoxTM1GGfXesiwhL/M
AgY5t7XgfRAZcI8khPCSJMEKqSGxJpW3C/9/hj0i342zJKkIzVoY55zxAYnclzzU
cFXNM1b03s2Hakt4jVkjvLIziMKBYCIaSM+QNZyCku2+rbtg1vTic5v7HdSv9bN0
b06p1xO90VrJrhSNVGM4GwdvUPAMmy6R6GQ5JXlstHqqnvVKEB/GqYeCM+5jlHi9
cXbLugMdhACJh8LedUXo54OMUWKBdGVxdaNSMr2hMvDZ9bzQj2kt0KR6d8nJMpxz
hpaarA4tT2P9bvGNZEtXrfeWsXIwKzYXUT/Sc3XaHyJQh+80W7kClrMTCqAeNb1A
YlOJBoUxMHFqJNGjtBswcRe3oKXijF3N+OjuQD9UH/2brJqDHjLxzVCjOZvSSZqY
JRu252Z5hO0zEUM2zvpU3/Dk8ZG8xjO+MelWGllXw9JeTq0fc3dKD5+9Dyoe3fTP
XcHA1G+LESdF+zI7bwSNmUQiw/ljLM1Bu9DMF2HpcpFQvPTYMlDZn5WhlDemi/Yc
slfEmvnl/LAh6VSXGGRAlRDKT104yKQCZ/oqm83GSGr+mmTfaqFL6xkhRSyx2rlw
zzXAVTPDRxdaH73U1eHwDSGDUgD5Sb7C3nC8Di2WFJcT1//8oB/KHEky5px/1ecu
B980/+9trzMsmH51MnXlHe8UiI4gFq3KhVhyC5U8rQO0Ggj+8iO/zBkwFzqleWCy
hwWY/gIOeTmVeUyRUnlZdZh5GyiUwJHX26BTwpdmTBVZ+wzkqN+z1ikcU82Ide6t
dhyliGIGZqIwixVObUDm2NoQaAaHrowUfZzZIBzg0MCnIsaiZRPtwyPrgR0lWM94
DG7JsTg04voyuO/hjUnoy4g4miiGTErXvmbi0Y85FTfebO+t1YPLLF0fOqaNfAce
qfozKLdxOw/4a2Vk11VliIrc9AzHRnYhDlb+GKGG5tD8PxsGjob2uzuQa3ta8sPz
olL/G7HDj+pko8Fwv47REG47GmdUy/2fQ+YbLVxcSt53c0g3U92u6mI9v+bNBif4
WN0sJ5TMhQH3kRjR3Ksn+JCi4Q1wHiUA8hWhY55Aa6GXK9UUF0D5MhA5dAvfptA1
u3P2Q8GRgzRzxg7dRdxw6TWaovVepZuVvSpT/DGMDeovJT5uPOKRSt18z6+gFQ41
joa/m6DVqFbgsJ102uQnxmRl8QJEn8RPunMetgEKRBNtfK+9rLHg0xMQi5LVPjLS
cPNsQNKEzh9VSEfSN00qW0pJ8c2PAgqJCNZ7QYP8T783jMaZxfq024dHyxPXp2/Q
hJFFPlc2oMYNE3gay3fe4ekhKcFwOmx3n++oFWNLulG1Bkl1robzmt9Y6lj7v6Wy
G9s80LIcbUOS+kGiLiFmhrOV/lPkeZLt5uHtRnuX562YWtX+MkB7geP/M2vku+02
lTdxuy5lrBO7ESxpqJaiCBPytMEfWzOG+KEHfKswS/rdVkMtpUSJYaKlb3JZB+qZ
I8/XIROvp8gwA74dDvkaZ03jYpscdN0SnON7xCHLgPrjHQyQq9lusAljPAvoMNPF
FvFTZQnFcbjV5NPvk45SyPr+gImRCOCICeRgiCfdWd2pcGEjZJ6O7VpnnMciMTmh
o5Acx0yMZCtzBKMy5KIVgmOFVxovDzjjUufV14ZuFBXK4433KbD5x5zpPjWiQ0Oh
awsSevmqajKPI67xiXhsIuADzX2Bq6Txd1MTl755DUTfiVwmZTfQ5J0H6h4+AY3V
U9OqRJli71kYOQFv9NDHygxcxf1IH/oXI8M6EOkAQ+bzUblbVBnjmswe20xEmFI1
3Rlb31VqosnA7NoULrkIwW9riX1Io59C/ZVuT6UocfZ6aC14dVj3CDKIzR90WRkJ
NuVAc7uepWlQSy+yalPVRG/Uksi2+0CoJbY2yN2R1n+B3vkIC6MoOs/M5ovEBhH9
7ZhwlSiZgztKhLy0US8PAuVXRyAtSu/ltJEWarPLkbSbjxhMHVTjbKNAQT8rMLwA
Lo7s09wajw97SOW8BfH4om2BrSQC7qXkdbN9ozit6ldJ2Z0q4ph0D5R94aHSbfJ6
7XlwLefenWGLxnNrpm4Jz1qv6ESlWer5Zc8N1QR8AGqjUMJVDeIFbItIXcEmUj4o
JSBAn49Q59LJtyGRvT2QHqQw4lxFnu4FaxwpHN2aKp41iyM4AhcD4/sJt61KsLuc
sIg+bbM9gPUIlwHvhVjbuocvlawrem85E0o2+EP6a8jzq9U7Br1vZVbSC3NFzsk/
urJv+YDbzKkpvgXF9zvPhJ6Rg9WufKwDrDUx4t4GaJ//+U1clAqV1PgzDXwFjqXa
cVT2Vy+UIvfINWhzeAfK1ni9HkNNT+R0TZW9Q09YhWgMb19CiDN/smbdFlExUpI/
mTfqWwg7MOHEvAp4JQrd4Fs0aRv7CbJWy6c/HOcjVGXWpxvhgk5JbpomAHYED55V
0RaLs24ci4VHhkQO1YUWGzAVkPSh9n7cKa8gGc+zXD74xOCmJRc8w0zhCKhTjjlZ
+VrWk4Cl4GISArAcejdkD7MNGUve0rbu4jek3qyDzsr3NgQPR9GEjvjXQxnxLaAp
O627UEC/MTzpexCe3ju8XthBL6tATxaolghdnECzC6stHl7sEMaCR8Ldt5GKI6qC
1/fCooILmCrsGAbNKnGc0yAYPtlRmIXkxBLhdOQxxajiMXuRR4QbO2SMp4if8lI7
7kbETQdKrRx3oYDZCNm6ULk+CNgiUWjV2tMsadXSN0phFFVlckXXRXikGdLNWsg2
E4KEDdTF+QQwXv8R68jLPEXT52c0wPw1jjIa4Z+HudVwH+5d7KOimXuVPxcZLf74
JigINo00Qft+XUV5GnDbN61ods/pvExDgNGuUYTv6rGhRsXOWM+m+FdX34bBFVgU
Eezhth1/S3VrmdDB8w9UyZ+TWR6T/cJyzrg45CqE5CHkpXZx3rMWMKE5c6PdsuO7
fYISAKHn0n8+b1D0ROG35z08A/NGuVwMNLWbbfKUKumNgdbQu0o+mHA1clt3D4/O
VDLk+Ci8nvxgvPQQIxDBLli8RjoMlOZTeonq5claiD+wurciCy0okBEQQlE1Q6LB
pIuBdXpHj4zZqL4lyShKwrQAmvRG+olM9/ALyXx++RAr8mqTN/WB/uDk0jugrN8c
y+6kPHHlF/1hnjzJ/TghL5S1OTlWA77pF2Pntnxp8CXWT54mMu6pervpTr4qFpQa
9aab3lLP1u8SFA16bSKu53QMqt3NkG6DW/KD5pF69NVuOBt4TMvlFyIGI4pnvhWE
x5rxOGELOCgWq/ceCHuT0Ud80kFaReGjPeGL+eaPaJ3HJZrb2UUtNleGf692w6FT
zk5QsR3xf85YEuEt7iG76tgS95QwMQHmEbMdDLPpbJFfu0rj7i7e9P5ZLqWNdDHa
dRASixD9VRtZjMzxin0XyDCqL3trFkjd4kI2SpmhOZjxxfdLvHrMsI8o/WapMZGi
UdtZE0tJ51x288l0wxLdoiDTjNAWI9eFC7eVDvnO31H3+2ocu+WK88Xi3iONyJtu
C8ztM0pEtQHNADbHftGdB8spWA6c081oIt08cDalA+JwL1aFHioMM3VHyUdGeMHZ
GSbFlSEqG+X7UZCSu99Fx86GNY/0Z/Azl3un514jdyypqKrssOEdczAhNQxgwXl3
lnCaBX33Vr2r8siYDwUBobmTQnPUFx5YAr9VJCFTjzdePdgVlRZ0whjk5lCSPhW/
szTs1EU2mAeKRQfzvWTkN8a3YBDNAWv+8l74CJzS7uQzDp9WlctVQ5p/xM3ybK2B
FfEbnv3WYu3yHnv2XY9hRXSvM9sOgvGW7NcLBtRGjffRp4vlvVPBbJECOCByvv8+
ETrFZM9Mb3sqVFdHeX0HnIXizlitiaRKfLbUdHLDRFoOZYcpwPLuuMnMOY4H2Swl
Aya4c3qzvOEd9PDqyifEY7BVMy+HLUyE5Uk5/NdlpASnIub9xr45i5iBqxX28dvA
xdWSYlNLmLYo5KlrLWm2v8N2yHGR3wuFXWx0EQ/PZ9hF6yB37h8N3VFkdthJ0PcN
DE2i4BrjBmWsyjX7gYaJ/mK5rEfOKk0NYjxGzqu2CqMQm0/ujTE8a/DTsZoCq4C/
ASo9n9v1xcnYzWusM/GpsKc4jPOLF4WaWzbprsuBzTKnOV0AtFiL2dj3LPhQ3Uu/
7xB4Xtu0GbDoBxI0vGMqKPyVC/U1jBpm8RXztfBJDHodN5oaA5ExnhltR9HHcq7m
AXYoCCgqlfGDfoLgFM2c+TRDMzyL2ds8pGHIGzCAqHbpQVb9C+RGkiGIrUnAWsLy
q7Pbyz9HRZSFPX4X0k35WCRYSBoVgMmDYGZ/Y11m6Itr47b7DuV72iMtJjTHxCmp
ixDzN/dW8iS2KJE2qyUOPYHLOyvWwL4QlFbew3NIfTh0DwU0pbA6aQeziJbRjTa1
y0KFf6gvxDmoQIjbbgz9y1qOHj+gFN1AoR5EPNL4GdigiNtnGeq6T5hc9SBhE+F3
XfzT4LSrVUF8oX4rznJoIdVb+0pRtPpcrAwZNq1eYWHHEvtfOt+e8EfUQyRv/plw
AdOoqdC3HkYvtdmJ5lof2OpGmwyNWMQmXu6wCvBBYvfZnnQXFu5fSPUVDRZHCJIA
nuG8KYOHMqhtJOAQAiKcl11omAOQGE6VlVr1A0QQHHjapv4gjMp/IIKuahHZim85
KCEUXPs71zSZdsdr1JzaN1F8e1MFZIFqXMTIagqv1t/MMvWlTHwzDzGPZai2si+j
QZE+9He+TVOAfF6/fn6cU84lZLbAxv77GU4qkDWZx/nV4VGrcHQ0kvSYdgPs0Qvo
zBdWyzAhq70ckINeh4mEPzOD0cabRaLAa/avCawfknLjjwJpb2wuxtjwEaF3DwAn
a9fJqOZrSjg/qAJn3tYGanWZHtKHDBqf0CFB7Ou2N1PiHLHU0A0wb+T0WXvbJXU3
82qjqGS0LxgUg/tnPu53cG4bmYaDFe9ItM6Vmwo3N5ApEOdiz1ydn8h+0y6ayyfH
8H9txsT9vSZ5VizwALObYqorROEL00bn5iP+AiDB0DFlGXMWbAoDinOkBn3U6hqh
p+ukMrokS82+GoEOhnr8ABQl8SQvPGTbXvVuXOyLCwogJvuOTFmZZ5du8QIdPb1T
sstTVWh8k5yuOtvGRIyzxttg4ZR2lFd//f6hEMZm2nbnZG+CrINGtFi9iX/5wN1R
bsXPZHTWT+dIYIOZWV1jGNW0wOksLB58+py2r7o9pZ3qfd1osSTmhyu3kbDj7Uk6
o0yMco9Ds4vSURjQJFgVy4qRyKua/pFBWOjnu0pKcmD35dOsiMQ/02X0J8x0VrX1
FxPRQjXj9K+Y+SUBbWCrt+WxrCAKW5wJuFOcKFFzpOzhpARqpdPkE0kL6VDeYgPq
t7yX88LDiyuGTudsUpByaNSQu5iRVhbM3D114+7ySg/uERY51rn4hq+47ueNxoIB
4KIUTStp2KFmIfMOiRtU56/VE1CpdQk4bfk0Z8wk+a2ALiUT76dUcDIWd/t4VRms
kBkurgMheZ3FdWlBGRNinN25ja9Gs0gDcBpcIjeqUlydarp4mSPoWHNGH80RV+I9
0cUWeXZz1+sE1jKSeV7uZ8W9Y9lymqIcvuSbxCNkKlVkCrGH2N8SrFUl5nMks0qi
bz1+L4qphYDoj8K9wDsaFA11Sv/KADaoJUby3gZkgrknB+fHPWlwZ/mTEXQmagBh
TcofRDNORg4/TlaxfWOVsPX2m7avf8u4iazzx267n7BY1ZxiPZVszlDnchT0fX0b
SD5WSdFrPv7obAhpjjoWD/S5hJiCOkqOOn35s4vsMsWHZIK8C4wTe/cWb87ML/2K
B3GPxQ6tZnPSRrz4vXi3ZAgbwTZHzRwxvp2k9jpVklJ8Uxy1l9ahs+IC4RwAcAMu
4UShWvYxomFXpcCpXHJLLVe63+2VtXOkJuKk5YPOevzjSv6GiIrGof/V7HkYxvxE
tyu/5fWO+gZbMIX2dUc5eITBzk1+GBEZX/9ceK7eAFUcGVayyRcUmAQmRg1yqdvZ
ysfbdTyNMZlNXEOTVsInHGzzAtEpGkXmqMeiwXiEpip+qv3/NvX06nUa9ha0WOg2
kL3atdZUQ91aWG8uz3NNTOvyNAiqAw3vhfB3JXcjhIR5dYElTM7vFhbsgrwsFm3/
QXgpQ51KOnbKiohZY3KDQxiO2vCWoDwC6p3k/lsio16c6EH11Y3xpZmmmA4pFGW0
rXxAuJ9m3LTMoJpLusXSfuD6I/qJ91z0XE3KHuTT9CxVh9uUBP8EhYvWFbxR6X+T
2hYtxQBckTdDOtJ/JFXc1cgrQNSutGGaqSOJqsSCnYiHcmQbOv44rSr97lsZkwAw
roHQc4mqDVeFmMP286/zzhwI9+0jx5QE/9natqPU21vdl3/QHr78vGJq2I2dr4MD
E6FllnNyQR7F9kV1yhFltx5qgHoQVVSt1IBsqb3mzZMMOBeRmaK7RghujdbXlNkI
BOo3hR7GDje/79PNkjUdxWe/TY8GLE0ljd8nRxiWvQYPo/LFC/CL0yV7uKJKgYlO
4TO8XYkSJ5j5ejDTw/1TyUhmUFLvgYFjj9D3CCSsRcGrfYWf2SCrA4o4cw+Hd8rD
vnmZLuHopGJIdAqR48Bu97uOLAMIEpEEJOBZDp2yQDzrzoOcws15v/15JdDSpsm4
qn74EGfXSlvdWT6bPxWhg2+bJgh1vWfWkI7wZn4imR/2xY/AnuXo+z6l/Iwl1Lla
6tcNsKJrusTsiswujTzepyG2MvsRCnP8vTm/yDyrzkjkb/9QfYeJRRmojURQ1L5D
9HoFHvyWFXrHcw5wbYcyr4HECjy/oBamiREnbvUCP41Krf6y80OiVGUVXUfte0Qk
eUco0VHVUojCDGHUlisUvyeZbu7n8boF81mSjSmNb/LgKS89wjWTE1mwxamuoMq8
5B4NpzMwBrjdR8OsTHcrLgacdd9KDtH+o5I6z/WRy/ZBoMSmSR4AHzvut5E0zH66
29m0GQd89KcJS9eVzIe14h0cTxhAi02L6AyS1Is6mPVw0kwPQBpLwcKwyn033zJy
AmCQZLisDfH2KHx8Eo8JkN/+WHbfTL3JLXUE2c/K97uprQXhBWBE3bQY4Jht6529
o2rpP5dKDvuDMLKazhBbyUjNHDgsYS8qj+L9WZWZkpqBTVXJmU3bL/Rd+WuXiPZD
ZVYw0OkyFZDiXf8yg091Dvu3IsOhRZWaCF1OFj7HkzSGWupbaGozgL9uh4/Qq1pt
SPHBOpYkR6S9CbL8jATaJ8tzFnaovwhhxjaXD2zGefbcnFS9YpFfmqP18/AjGcPx
aiVse3s8AUuIm6QxwzbGyeR/fG1+WpZ0tt5bq3kzfZC/O+8tU0yvU30iHcK3MpUG
GW7+Ld7dJAkahM+P41vWvO+AfEA1S0GvDHeBkqryL19BZPFupwzG1olfne7MEIT3
udIuC0uKPmJSwEH6rlvIaNPSYknaiY4GbEPhNTxvPNKIZgC/RWtm0rgBz2dAISNB
8CJcc/TWjh1kT+0EejqbQMPUzO8qYMLSA0ycFnpA7BKDrEyT68AzkrV+QWSV/rAt
oHxzQiNEggycUnyG00JkULcYjdbl698d4a2QjWN9XD7a9v5+/G6q7wGlgPSY+2lj
JXW/Xh2+DAA1XYZ1A8+HdlJyixdVmNnYauGsYRkZ4KkUbWY6ySp3Fa/1Rj30BrOq
irkXHANMbjAfbjd/tnc7/4oJmHcn0/0FfGoidcuqDtfCU4jeHWRdcQHiCNsgYXw4
Rl5fnK08IXPDDeTevtlbJ+ZnADKolG/rJmjpyyK1LvlFFTUNIynEYa3zjTuF5vLJ
Bl0cdBU4C8bFe+RCQTUrOvLOx2sPQi2ReeGIu99Diaptd8vvtRbZi5BlOoai9O6X
JKHE2GhDtgGs0pAGdNFDZAtfLI4/88wfLlmko8DWNOyKGPD6oiAkIHpOKHeZX5ho
ePf10eevBTJkK2y1e7fZZlQNb3bQrC+eOLB9/bsVtA9uMvkWHbFQbSuhwYtG/y4Z
oJUFGa3Yt/C3/yxvGWDcQo/Ym/aPG036twezOvRfQ1Nv1rPldmAcfDglJ8/BctM7
jceoLlk8SQ3dcZYhevnWhGpe7bLe9TRpAR8cX+AJcIThUuJLk24mckHQXlzLKzWT
caijss3v20GuttGYQr2303sKtcRmywTOhXDMKMJ1kDGLEbiCI3hQnBD+cjsYG5/m
MeUzcJcSUFddbxAwCn07V22H6CzywtZgXTfsYV19cYX0TFkLKhtNTkiHvUudLODt
Wp5PI6ISUAWtgPoVxLLyxqzFkIr9PnNj8A5wlh5L1gyrObNqCUnahBoV+xX0vAoO
tGQeoy3kXT2YBfPRIFCSa53WjSYjIXhoj+3U7wZ+pWho6xnzkpvgFYM/jwuEykx1
V3X921RP+ZXnnGAHq9WFW+DdHVQGn3aaUVCMPSnUhhdx0kN+CmUVNm+7Tr4Lnkd1
BrRJF1qXop1LsJjngQHt8Okaj6e0ruEq4hjFYUiBx7yMBV9HVjp2pWbaoShEKsZt
RG+H25SkSH2a+Hz455Ie98LhWvf3G6FsrfjNhKaBQaKBE6fHq4O9j/wxKo0CMk0S
CHunkSQJENIzbPcLh53ez7asc47g4GpkVq6dpcLAQO55DZzOv6n2sFpMyy1zaNqD
fscunSUrB+K3AL/CUbjafDsyI06Qlq5riBVG7RNiFGk1MZGRS9mn07pgPL18ZVtV
9J9vHba8OHAQziDo5nEwUdHJDKrEYqS8LMDY1LrNllDLbio6y/kPNzVOoR6PBH6l
YvGnVO8kVRZjutycp6Yu4TP0Tf2CPt5nIbpBROkqcC4HL05FhQxDv3uzIxeI8tGQ
tEu/uJF1PxBU4VtH+kBXFY5VwryPmw1NKcLScFrAyBVh2pef5xjk6Jgk94aljT5/
k4JPk5CJVJgvUnA5PrAaUzZNTT8QjhQg2MJhHh6QY7xhixInZAkRz0NOwV9PoViQ
X/RUWpZjZxj/tF0gr9zM2pUcBji8r1+S6mlJobCCV7nn4jJwDa4z+tW0JJ9tdR0l
YF7WoFqUDVQ2+bAnTk7s5Nyy1msYc2+xkK7yN4hZwEpmKSH3XXRmTxwURzRwnqsz
4MAD55d3adMOrM2vIBrvMQaqIMt4hsHMelT5o5slcNy2AUM673QEEFR8GQ7QK3qJ
X/KnaBCCh4ODEXRR7t4CFpOBnZ+QiNu4e+mRmaVpkqkKNPH4X3CY3C+vfhzM6HEo
eqD7wW0aHdgStE3AulanofrG/mIpDL3Nt1gTYwTda7OiiUj0ScXqlEeUedbGvCDm
+zLkx8dLEjUYlDgEQSQTMejvf7h4u7b0Ra0SqmqCUzdQ42tc1E70nGkNztzwiBko
76rK0+FTwJd9rZfIMZigDEKrOpN4lK0H6X29OBVKbv68aw4WkiDHsA9xc7nkPw6M
evvbwS3FH7rsFhS1DYXJiEmb3nfI1qF03bdYo48Xnbdqgms5JBRkUdASxvDbybxC
OQplrPJYZFevEfSY7J92Umfep86JTB6bcpTy/QOdCMJBEVUN3Jm7xEdG+LCTDqiP
pWKB8sXkScsx3X7Mdq0B9iZoEFtCSyOfpTmeDXt9E29o/MhY3UfpUfJXHzSySICL
kSG0KDrIW1wb8wsZXZ0olO01hhDNpZXcNaqbwL17G9AGL0a5ix4HmZ+k4wYxdNw/
w8B8bltEUP7C6gIayzgIZpWIQAe3AP3IH658N08ZBAkKBFvgBx53V4LHQPLqdoBG
ZOo9nvX4T1abML2v3LPtD9kihB+mXfj357fugeqRqhHsb1qFNQruU5E+7s7HY8gu
7AEFZAcEMr3MoCyNqd+43QBQVpFpbZenQ7XQtqBlp5HHhGF4Zfb3JNP/APEBtJc4
WuaMUlm5XuIzdE00ZVG0s3cMHVdmdu9CmWy8p5FszdWk+d0J8wfkhXIz6sCr7Rx6
1oLjiMWAfDZOP+AOWRp51upWBXJcncvnvQEw61HHmwrWIgx973PyevVyNGUPLltM
YNDCGnGQTG9RRgTejC0/LoseNdW5YtjzfsEntxJANDtrgjQI2t4OXue2+Zz5xWKK
CMImwGFLrWOAomx5f0daYwPredvP6LhuZ7w+zQBHHw1r7i/FKwhojbKfPY6ce++g
UAwuuf3UsikopErcDKTZOyQzgd4pAf3KI7oVUShnDvrpSKesgSMssDQdEBObBf8H
nj/oJfPjOwtq43Nj2GjTkTsxLyUfhhucWhKMuYIbAm5Owr8sMqHnlcZrcMP0SLQo
O3TvZ7yj6BVazfspQRmzrpFHln2vuDE0zS1D5SCrg5H9SSTtgAzo4dDBWL7XZhjw
xDiwOWNlqv5iXNxX7UwaeNfGD3a1VSftC0lr7aHDKBQ3dp94JryQspPeH3Rh92Oh
XyALkB/el4JMPtr5FCw9c/77/Z/hMQHYbe1gPFF6juttkdmJbP5frocLckU2NcKR
/uor1jM+dYm4SD049rytF2Low/AxJkfYMumLWBGe/9l89nHAz47xnzuG9KCaaE2+
Ho/I0b/DDYCP+yi4TCnFuGvtMdYjDF83fFtRIqQ583Y54SLOEVna00Hp7CWKCtJl
IaJFL9co45IfEva+KFq0EIwRWYWON0yy+Sfuo0tezOEkq9eHIm4e56N6jJIp4O2K
h6dNmf6bsekQKnciVTXfb/6r79s5iq2KIDJKnlmz1B0WJIP6JYN70fbNkUhlR9RK
n9Q+sltz5Cjpf1HGd4Ap3NylOwsuZbiMyvdGURhky7MhorzL74F0T31LY4H/rbXg
5NvCW/QJE9I1ICFjmD1KS157x+sYQUJJCEjlz41J21j5A01xi9vS0WDdYsajLn0M
k0h2CEooV66P/bzQTFYJi1xI5X+WZuFaHp7YF7e/4nMKwDayipNbCfO7icOk6Ne0
yAec+9dUReuao+QZvB77cVpv4MwFDujlOzdfWyfYYMADLCNi2CA+446uGBMStl2W
0ojEjlrnk8tmdYJhk1q0DHwW9B5+iK7xGZiCPkywISLRTy3gtUsxYXt3ywGGhyqH
6MjjFZaGzZj4NpesvuxPkGqzumnShl+4rw20pQsvM3hRn3GW8biHUhcz63/RXgk6
evkzBIjEGprlfxO9lhtCqfcT7zvC83BQiKd94u5pFGNBb3KN3tMRliolPC3msMPj
/Rx3cGAxqBLHIldkEuHbuBhvNAh9wvzCUI15vtxKD7io6EV2kpy/gzl7rSiiNvcW
Rf5kZRHwCe2phlQZrukAxP3f/YmuDsVqB5LPPhwMcYrf+kvC58/yqD3hrPCn+koy
xIbBFKjInbscUygJGau6u/CLdw9IAULCg/sDhQbBlN+a10AS8qGsZiaq9sujQlY/
cv2gaVuQ7h+UOfTcr9H2pNhXoQ9kAwL6MwiZmHKL3YpgvyRIAwNla7P2t6HEuJ+J
IU4YaYrHoDU9gvmYxbzNr2BazEWptzQ+6olMBiMvlaf3uG+aGLspMVtpRMWGxUtS
kc0NsxUBIaI0m9TsMPtzCQT6Ugut1rNxU7LUaGLKceyc/o7cgX9nPEUcwXsQi6YI
qjjRhp3xMZAb2kQkAayIAIS2bEocLxN8Axa/diZFqizwKhijNFf/d13ySwe9Yj5P
o9JsGYwoUT3GY4rUA4+8MkZAOIqwmOEPKjjXOfu8IpTRwf5fkfjZor3x6MBJWDBD
kd9zE93a9fqS9mi3hPybGp2tlvAtADGYKCvjbKkMcJUiwFT+TiePPYXtBpNsG8iY
+XMFkANm7MCs10IeyAX9ZbaezbAf3X9zbLObwP04/m8LI4Nf7L6h2pJrHvJKbfs8
MOzyGipwmdjWgSUibsF788/yIIK7y6hPrseXD1q3wKCps6e1kI5MSQ3nA/9Fd9YZ
VYRPnykMeFhLTzamBfFrsHXdCo9d4hkRClhJk4Ur3nH7zi4hVcfazpeW8PJZyVDH
BmFFTukzXNiEkS8PJDS8g4u1gwj/Pj2E0B+wSr6Wo3GSD1Bs6ymr5ERyexNZ3JES
/ZZIYeMkXiMwTnvnISd0USAgHBXfJJ9oeKceQ12TUcRhSqCiER4CWHzh2QeHw6VP
xs/1mo/ae3nLQC2GliCyCdqLQMfHxRMy7/c55C1nG3g3FMJP0jAuJgl00WjIUzFE
+Ibl9IrWnMhfPrFt5A62sQZyorK+KNAEPo4YS2quZ6M//NuIQaDo6jRV/W4FCcug
ROgp0DrvaKx3zBnedYPcy4pN1updLiAQd4nJ4Vsre0+xJ2wMnmIKLfa7mUdmN+fi
1p/ppsSz+1q6ox8hgliVbFR5GWgXjYxo2snRy7J87CXmB8KZpjMsFo3yxxiEG7Qp
b235wPdkBwF2hODhxBqZ5u6hsiedbr+oOlneOm8HHwdK6MwXaBPNtagE7qfizxRp
ORDaOYOyy7k6CZPAa+GD7vy7Xpcq2W1WxnqlH4FCiU2sZdufkQ8ZjXJpw8bJRWFB
7DJwqzAYaTGDtdlngBF3Tn5tbeZDNR7+iuaL4jT0ip22mNogiZH93h5vtOOp9TYL
6wmShSwOMrb9iET4FptvpSlC+MizC/tKgMKZeg/iCK30GnNmoAYUkZl2JkJ+rB7s
eIn2pAwade49ASOf4XA0HPjQTwoVsMn4RA8qls8hpRnm7+ix6oyeHjEh9q/caYZJ
OIReEU/xF48rN6/ZkrDf4hstU+jbA/KxsXpxrPNiBKay13x7W2sgbIc4QTRnCntj
miuZp0K/giVpQQTm+pd6K/rajbuIkPmenKtNMxKHo63Pbp10RqKHHGLr/Y9NvRdg
jQ3GhbYSHZ82bkV7KWin1a/pa5ISKi/4KSXUz6kypJod7hbTXyi+qJKZvJopzYEG
cj8ZM26qqwi+JExJBQkK/OmoLQ80AcIJtAFPj81JXczkET/8dcWJAp9uo8hB2ZLt
AxEuU+aKc847ZOqDhk8hhW/HMC1FBTE1TOtXVztTEbfW2sNdo/I5Hvbi2Lw2CGZe
KZKn5pz2MBy1QD20uDBgJtjY6ZlRnIniW8E3C2gxuPj+RJ9vK0fxOqdSWFZ8GkbN
adME9JlKNz3amIicqxIbLNauTszwVlroVUAxAiytKFciVPvNtH2xMOCl0NmA6iVX
6xLh5ErgJ2M0QpulHT0kSx1CZjFS/Wxvz4BW/dqZoQio0YklMFtz8ZsOSEssURAP
/dPsh8OQe7+5kE6Z7jJ33tKWAGMClBV45q5j16kYqLdthO40fgWAr2WI8CgruPAZ
uF9d3d7LaW+v8EPxMowZ/2yzabvmS0Pf5oxVZNsSVoj5TPtfbCyhHZAaIfg8p1Mb
HE2HQWm9t9mhwyk0b74MuIatEGq85r8K42Wc0+CPy5dq7OTpk8FwK7NjjJKGimL4
vJjiryyZr2rFx7gt9h3+RzCHGnhjt0wPxH848Ye5ScTPJUATeuIZ/9tt6H2FrXZ8
XDuz67wAtQbNC43Sd32AEDfrUGXxdBwPfvlE4VDih2jlh/3VEIfJTnZ3caoUMnIF
b0O/oMbPzfzmq+aVWFYfqgAO/2UD73trMpQWbfPaAugVW/PaHhOH5vhu3pDsoeT+
ezXimYPMh5UUb2ycgU2ABpV2WjL37h42n+vYg9y1jYRZAenezi9ikUF0gVkl8w8w
0yNohq2ig66IV0NZB8k7aSg+cNGbkV0d2O/eqF6J4eEVVEUylvwACdhqQsagpoGE
cGRCLlF9vSYDGStL95bsfhoH8zhNlEbIiFIx3eTMHjvsKdjCHg8VyC9mdKTKUWSO
pwfrunXOMRBtmKTaMhtzC4kj5wukDqnImAesUUuZsLqgKOmQOdbIf03cnlEmHIVn
mEieZY2dYaGMPwhQZf7iA3Oc6SGPHA8vv2+IA5KBUsEHdnC2wMtCxyipmnEQGXD9
aFv+Rtaxj/hdW3mOgsR8hBNOZLNjHh89USeWhYL0U0o6itu9o3wl/Rghz+TbxM9+
J/gSJhJKZfPlm8xnmr0GUfew78wegDcQ16Uw1bUeGozlRMHS9auJMboDkeJMf8b+
5RYmM4GZIJPJdn+JO2REDgX6H4di3RtKG5fQgA9R4HBDwrZvOkbDmpHRh6ZN0bYQ
SmxJvHrUW22JzYfitTrh3IecQQmMJtOz7fU1GN5hG64oIks/weHg73nLBv/aiEVZ
u0HG+7XA8qPnkXsA0wPJ+O+nK3NiY4N1zWNeJySMeHo2UVGx+YuJ9gAKwSImGZ2I
BG2mH7n9MqENHPd1Y1Uet9f/irpZSbqk31p8uCtHz2Mmqj0nU6VLEROSN+eps0jX
haQG0OsCmqEEzkZVTwa6oA4OGUS8C6SBHFDSzyBnUDYSRxKYP9sE9OUHG+AxJiJE
iAbLqNU88Z0rygyZ4Tp3FbHuT8cAogsICEGjXFGizidRRACiHjrgNb6+I6k7HK44
9RcKWxQsD+bftzzdN3EbTJvtgNQ2d3igm0O5e/12gPaTAfUKO+p7ZnDQmOQvQnL0
StVg2Ur+E60WEER6VTYkcUPyZ0K58/B1j4DTtoBlCVYsLvWcPorPjdE7VOBxMT/C
5PzaRupyXztXE+dFZEkuMbNWoR9I3b6gzeQx3FiGIh3RxR5H74pZZnGSGm/SoZFP
GgAA3FOp15A3EYMkRI7Go8ZxRXsSFp1viWq4BTZ65mwaP+ExqqYqq36Whs2lGNUX
8gxGNuuo3WxxRxTvKYOH24cvYQ+M+hHOymvQlHEHbeA/pRbQ8RmFGO8KUjTdVuiy
Qgn5x2FQChTFDFi+togOZWDHWIQSjGcdIgU30gcdOm6sAlqxVM+/9qzcCyXR45nC
gnZB/Yo1em1XX6241kwaHZjqG03vRzgEByvHdS8byy227m2fonA5SWko5OSLXvsj
OUw9oU4ENCb0qidnDhwBb7g/PCmYMGHByxMBaIFnSSHF7VM9epsXcSOBI6PPKdB1
iSJRwU0SM6AD9j3BPHjmbth97YuoiaEW6QgwuBtAJeCLy+Fpx2ZFaLPElE4YAf05
Y9AmGZ+mGj1DhjpDQ58xPH2ExGPJHCZVBMfvV/rd1AC9yOkPUQ5lXVKaxZ39LFLZ
S5VznB/JKw/pwGHn5U3sEf/M5XdF8RH9Z2TGWv7OPkv7aK8u3nO+gshOcujV7eEG
d5wXZWmF71gzSP6mNO65kcpzQKaRX5dqu/6P/apcixNxo8R2p3LVKlZGxfBu7QjF
nQs6PNq4IqId54fSw64R+YxvLHvp+2lvQCn/M0PiwRYDUjR9Fb5OPcjhUaltFnE+
wIJ6+Uf4h3TJJmVR6VUI7ZLZSfp2IqC9NbsMw4Y9GE8S9BXvsovXdBODDD3+qLf1
d5oMLmSPrr2SxDmVid13Qe26k+4nWQU//u+uZHOYhAGMAFe8DEGG6KSKk91r/3T0
DyFrcfTtyUgoYepg/rtVFaptHEA6Yx8Ytt4VqFNtypZ0ht9IdAi3TaDxe9CDzfY9
o5eA4t3K4fQxOGttMQJkLQTXyJr/fr7hroN/gsz4OXeKzew/vprqKHzaeE31egn8
jZj57yXoSAtfiENxKJ1HG5i3VdEgwlV/z9mQxNN8LODd723trB5junOY30sPITqI
WNqr9rSe3K9xuBkcMY3sXbptGiXkEAJACCqlRwuoMrm0VC6K2yBUTgfGW35eAW9W
Xguk19Bzxl2Q74kOzJmwvvDF1zbosGDjC5H5eTQZOqBjyPCXHZn+2gd4bcpz+5Ih
0hadjvO+sInvbwVP36YMD4xzOg/WDrgFaf8oaijVLulNGnEaKbcySakOpDhFBfRk
0IZOcxtDfWdResF35zvXbWVGzWZT1jCAstCpMG42K93eDjcWFqaY84IBuMGpz6pw
PXiCM80wcuHSgA3Gw/5CGD1fy5pTn2YvEyq+Frp+MyHMeA309v60tEXwsWOPlDRo
eay8oZs8vKhC/8KKVwdF/EVq9E0fJrXOrCZRJB36yIq8gMymzbn3ktEzdX+XzlA3
a9+kGSfUxmveuvBiBntPJhLlmlC/SqYxaeK4IvB/z0QeYbtyYDrSqD28+2y69F98
Ygf/XMglUfM5YB0uVtAU3wJYIiXFZc10d+gcUfplWsHkND9te0kox30ILW2UNx6g
hGa8QlfVi2GBfa7em0ehycju6bCxE80UQ/2YiqDDB6sbShAZl5pTqrKI7ZEuoe/J
5/G52x10xZ5i8cN3EY0adf9LZq66zqBWjNU4s/f0eeRk0OmmYNqHk19sVu+90pyd
idvXo98FxTdUwidPtfxGk4Ghjw8VBf4jquTgJmICIuHgBw3Lzt5cvsbiXe0l6hoU
IKdFTgU64hDSwCQHj4C9UxNDbqUX78UI+AbD4+RUjUjQ2ku0EjMU+dfJ2WjWyRXK
omScSaol5MqZuFYx7DLBdXuwm/964P8KAFcN/xYNu6QvyHrX1Jvfs7wdbnJgd+P6
OPsW6VvuuPJk23gPhSEiXf5Jb6oj2lK/T/nunbbLqXnBL3fnPiJ0whpRUPiMnt2R
rK+exZ9ojh3yzxW35yOAN/qeLqjMQ8fzxu79RQIgJnuaKlAn9oNAfupN/QEAyHtn
idDtot6mif8OK2+2PNc52sq2LKooQ4ZQUBBd9+uOYivKlBdvIoYm80yuZGOmEOIR
cp6W9x5PLVW4ejCWKrNZbnEGdGpwiEMGUd/Wpnj/RcuV6cMA07mOqFsbG42KusbI
K94QxH+60GvlIh3TaRbBND0zAfad0vmrkzRpWGldofKMFeaJCM9RP28rSQEJtBZv
yyRyk2937M22Qa6jfDEK15WmEpGDtLYjmvFaMNFaQHnTmhZcf4Fd/GAOOdikdpYc
yVKzLuHYogLKzz+1ivRqA4gkaY45kTk8NiYPEbjmmPdXidyi0q3hkQSlqlbaUFDm
EV5sfmIrHWze008HX4lkgzjUJwoCMFWl2aJWvuKV0aTZbou0i4c3nmx3jTjhMKT9
a7AhL/yqbr7lELo5Va/GlqjKySE0e6ddTmgFwqx37JeWNpwozRlc/TUjJd2br63D
iL+7oo1xQdkdVFHAan2KJ5BhZHyy8ZXjglPhtxKptkAeeiQnQdnXruKqk8z8vbsz
/6M7csvfJ2pgJKfxWdln1xV96xSoiJgtsznbqH1JkiDVl/z1UGR7gt9lAvTTFv8Q
MF4/4Blrsixce/OfSmQ7eUFb3wzZrZSVz/XO1pj4qrekVZAooE8swsBmQ79xIgFZ
sgwe7L1VPhNrMlxmsodERPRupRb7c68XXr1R3RK9v1Lxv+N3yTTGaud4yok8nURl
ZsnU+hkmZLHcTNuGsdCv4Xw4RrALkzsaJ4ppL8k7ue/X+xIB3bAS77JNQrrDBOnS
STGpNExlZKK13PxpDjAkYdTbSGAYKWhFez+bOcVo4Bj6aZmX0CnGKL0+nAEwrBH9
JCOrYURliyfk3sWclYG7LSb9gVCDhEuwKi1TbUmWvF8chPNH03o5M7wAYf2bUojn
u1QPNCRQoeMafWgKf3qTPKfmRdv1837E5DgG6BeN01fdZXl4QbgbhxV6OjngOSRJ
NDrniaoHvJV32tLDdXia9kZRA8ZgAoS+nVsCGeqve6FQIDufez3qOAyykQgLDfWB
t7kEDWOl/AncS0R7G5RcavhVthrxyVU5OrrtZ0H6YCgbqv+SL3PowhCYGYIIlDp4
KZj7VnaCm4o2sT7qqiFYvizJJ6eoTSat5OIhvy/eeWhUngmgSmF8SyBbH+22Z5ts
Zo77lOY6wGP5bqITPKjUK4WSmhDFrIzXDP12b/MPKv0UTd3PiWwn1zvCgM4V6Q0P
ZvFHOSxDl6EG71M7ar3fF0e6FIhGuix2DPcin6yZPohYWF9kPTJuvKf/gLZM/Q9G
K16ngSdMkzZmNQ6H+KeMqUHSxHKhU9IYiv/kujiMQYcWOYCD8m1pd32BmRDVovpu
oZD7ZURPS65QVU1LEP8bwho8YmOpTreNC7gGJPyiumW6Wev8eAFKqMURy1YwG1QE
Vdrq0yxV8U5xGs75PeRS9/9y8zWtW8u/4tr5qEhJIpOxea4x6VxmK8C9Q+cD9UVW
zrtXgHPN8yF+JB1S6aPnEJqqyq5u7X3r31EAf+3Ex7Z3UaYlAJzpS1yDAwqJYQdj
fmuopnWpd01b3aJbc/1dSwJgT8imW/QWddgipqW2kzP/0Htffa0Fr7f/4WlJPhnX
Gd5BCubAuPiIb0oJmFjKJIQmH3T1XICgLn61+meonpU7s2kjRQ1wSraMfzGexjq2
TRKh1CZ1Fd9Q1M3dGOffNdFExaDG9gZQElH+DEjirZHzDb6Jg8fFsmB6+yiTUmmc
HsyPRCWIYK29Q7qRudrG6mqOXYpCGKrSC9zwbV3VrSOgmYl7M4sLAaLtn+WdAGFO
9KjQlCd91GvIdX9gQfvEBlB9lHq7QIKSKeduj0c+8wILDHhawGUVI4IsW6zkOUml
MZ/SOumjYDTKp+8V3VGTkmOMvNQhFBsSFjOpPPD16sE0OL++3vyafEHkVRf9yWMH
dGsnWTfoE/l5DF3hTXY2NL0MVy70FnCfn4feHyfO0BgKQiVKXWRK/ZyNJidEI5rm
dul2CXTEbATdHIxwMFMxdaC/OFfnaJgyLSKr/WpmrVa/iKTKv1yqGAYA2TAHFFzz
yqehYYIjyWcKS/T+Ya3DTZ21vmifhGaj/n2pikADinwoQquLYrz09ZCtMkxWonAR
5LGg3TnDyWN2xHu+v9lq0+NxTqMdbS+nispjmLRjBz1xSxJaD08RDRJz83m4jeWN
maNaVA6BPleGhnfbCrOCvCcwmfefyqTz9z43/eags1qF0VINn3tD8SSoV6+lpt07
pF+ce+8/YI/J1gfTdj7B0XEQEgMfEcIovlFWFR1wh65BUdGswEqmm/dgzo+DgNHa
5b/aj/A/mEaqURjePgH7PjG0LQHsHlq9GprOiDj0XCSe3gOevBn3vxyyeBERnYOV
tO9+c8RoHNfnOSU0Go1PTs2/nSWVlD6Qm9wyj9otn6siyvVfOgQxuCYlzVkY2/uB
MgovG+kwpue4HugNpn7wR+2oVn7rOtrhRznHS1Dxf5g6wtHuiqHiPdGmJ0jaCe/r
Omj4dObAdSptueZI3d/TmnBKoG3+/3Qz2aB54aoLCHQk+T5Itekcrl6vNtb/cUxu
eFolzVu6rlD6K1P4gLCgpUaBY8/Liy8XeajC8gAzJgxCMiZC1IIQYotfAFdJyduF
meBRaOG2QVy9Xk4P0GO1MbKDl2UhQxzhv5rR6bEqk1vPpls1dja4BJ9HW1Vy+sCa
xXdzT+rBjXbHcS80g9pb6ll7cNJsQlXqkzbrIpGCgXV7tRD+VTecWde1GAkIRu06
fcGZZTdAiE4aak1YNNfDPT7RiW1oONErFwyCe03/BhKQv/iT3Pan/VRSQVS5qvoK
Skqbw4HLedtP18epojU5HYJtoCQqRiJoCa3+iUw87kI2tYwwrcgNjjWxnaCDa4eX
h82P1QQ7RYNAgZSBMEFINkSO7PwqnHlaoDNzJ9bPRR3BKCa4DmxYU+e0XYXl0dQ1
yMTMJ7aV6oxUBHeDeix61wEZByUaZHVNomW1EZ1ONiQGnh69RoJuDRwpUfhWv97i
cB2Mykny3h7xDo3oEZOywPyX2LbFNziYZlGvkC/lyk2tdzm43+mYN3z02pjNDpPa
1gm0bCK1mnyoREw4xbUl5K/Y2o4nAyZ97zEbr40+0voP0btb60oKi8vPETAW+Ybs
OwRBScTnJiJGUB1Ax1Y/9jP36mNsuFhuLMznYPNpnKyQuQwiDb/jfoDVjm4+ORIC
IWi4hxQfi81gpjRnqcI4l4LdGXzGciblXCHSMpFtcG42/izBMSRhhyv5NYj/OGTD
hrG9Q7M1NqM4lZgxKBKyOWvyHQ1crhha+p8mVxpVI354yPPIx64Cq/LQWIocFw5J
Q3hzXgz2fkpV93jkz3R6o4vXcUIHTSr4qoL/xhhLoqMeHZOrpFCIsbIYcJXX0QzO
DDcPKiXTagCEdPnKi87TNqrZa8pQYj778xn+A1lowaDaN6zh4kXMkYswuo+bXwkN
bihWnpuR8McP0D90YGpu2+zCQOOrKxQBSs1YIoUEpATVdTESrwJHLUfGVev33b8U
lJ7otiePMTJgfG0uSwfkuc66vATXLN8RnaV6kA3qYrA7y2fS1IFAZI+XSKoUKmAd
SziCgyg6cok/k6nDexSPutBhgOgyr7Yd/UJGmJTglIoZpDlHeHQxq3noHhS596Ts
8bYMVIUgkCFEwH4M25zyeT83mnn4Cl/48LlHuex3KagJw6A2TW70U3r6vS0SbFN2
O9UmSHhbRtqL27gqENCqiMxTMEPt/Kdz+zK3JeK+WpOrG2EMw2z8dSTo8IlcJ9QU
rEHt/UJOc000xBqx1gP2Lz0Th3Mpy6y9stHahhVUK4bALF7tih+qvqRiPrTMZKac
s5593EJc3zqRBmmmZNUMYs3ObiXb9mMg8zJKQBLOjk/Hr9aBTBexFdw5F5fwvTxd
ACATv81Ql88xg6oEF1QyeIBr6z4KoTUhwplv843watLHEOuvUMR0lUCy5kyMc8Jn
qtpNtXH1B3vzfX2BFhpUrh07OwHButq99N+1oDhe8pM9QzKiTP/LOXWkMzHmvgKB
/qCZmgRbN3+iPw9VwgLo0dq1aF5eCxTGfXezQNBBfaXPJwoG3kYU2h6GmppGiGUJ
fBqXnyaNwH5+Z1ezBKCFjJZtFc4zJN9FRbkifRaR1PfEXT1V3oujr8SxpQbRtmtS
6tKKsMAcLSJWYjKLIxItzMwP6k0suIMQ4bfWUJ28ZW3wMLUjbPU/HBuUZWYscYXm
scvmgFqYpUV4DuvtKWEr+UMTE9AdZ7ZZkukyo2PS+S18smjp40cq6W9KQ37mvw54
PQuopjBvznE/MrP4us02DvU0FE3VM8QpPispBlw3xC3GV0FPLfy+leDHcz0fpS0R
MXZPHA7KM8FT1PRGsl2n6VXHhrJauRlcWXRHl6x5i2TIKzO0BO5ga5U0+0zcM8Ir
oy5m9+XoiIPei5wtHnbP1UPUk6GsDCxmapPWO4SbwmnRG+V7jZMBew08A5U4LFy5
1MQnaH8LJ78Nbwl5JGCGhH3lAmE5SjXf03rIapRVsFWWfCSe4JGUGL0VBYB8pMNu
0n96PtzILteOnHKB2iq/8wP37nufk3Tte6TifZSO7EutubZe0AGXe0xCp+GB3sd+
jUjxkfycL7cUg/Brh4jsRMepcjgXMTXJT34kURDAs//zR9B1YD0iGQ231GUN/MS1
R7rCv+D4GS5/k3a0UqxiLuTlSWnnN8ApVpC3vAOoZBvDJCBl5Jpz4RDVXDGijI6d
Z0VbXE+HyNj/hICFyt1aJ59QDrDbjYKkd17UDCFdVNhVO19EaR9GkE9shWQIENuK
W8hZLK1xFY/0EH7OlWh5Oh97pOybtZ+KIXfms2VPTOKBuvFoM2jrJ4eTNNnYoLuY
torUROQqJpDwB/roPVSfSV+zeAQwOHs5my2n01Q7xro8Zuhv2syJZ40yqzWDiE9v
evcEPNSTQLkUnidPvH8CAkedNXaYZNoqnnQsdXa8PbYlUERTTncxgTuWYvgFtw7O
RfkoqHaG/9aKlAPevA9w6w4o4AdxPEEy2BjntCNepBcHvFBBMachZlocnsFdBb+K
EEGcD6J2+IJKvkMhq5716rSw7owisxz4wxs1R3nM6ikRrr3HxUqvkwOOSvAotfdq
4Os1O7HOo0Gu3l67KKqvFo81wPWlssS1kyRgEGzX9bHNgjcvjgC0x1x1DB9Y15yR
gjtAbGZ5KI+OygB8jmNYNpy0oC38ridmkkCe28t7RgInr3DLNDE5JnlAZ/AdAiVZ
pPjPqT44G0OZ1d9/qsfrm9PKIIiXIrtNxzJgrRjtP0I8h/LCCkPVNlHcX590UzFw
ipIUvN8xXsU8hxeLOGGyX+t6NVo8NjgVpgSQB534fwaBmkUgdoenRzwaKJtCfrQY
3EsJ7qioGMyS+0SBYd9prl0XsIN4jGyBmdBeXaclFrRp4hhyQJhOLCRkzSa2D5F2
hLWiVS6lcNBqhjiKDGDv4MYxFtiW0seLCFq3WRb6Q2f/cJC7BdYnmW71mpAc84Yb
wHyJXZRn5Luw1UU/QM71JI27ZI/pobjGn22mrXIGntI2lv633ll3BcOGDaKGeffX
dubhv310a3MvPVVvOUBcHnhBvpztPk0/mc2eGSSwHyBa1H13a39OIaBuHsGl6MkU
gEU6W897hz1G/m5Ww0MXPgGoPxQmPrgvteBa8CxTMclQ4MJsCYqfl3FD0StAv6ku
0PIlU/GihhsYi+HGx/NFQ10/jgyMj3vUqoaCNNfhCeJ6uHyJX3vOaI/T7q3joeOH
D2IDKkGaTqloScyOfu2EiE1KjN7Rd9RZFjt1WskXKZgnUdvapmubJhvx2sTPFwlR
e16NWG5+l0T0bRo/7Uz0NPdXQSGpZrc2d9zqkjSTo87JZALX+OuISF7eTPKJJM2Y
3FUUEsFXkss8Pzi+Cse0GBerOCZWFi7yTu2XlV0D5JjRKEu72u6bu2CRqLNDXHiY
6aCKLm8dVQiVjhOW9SbX3oMEvWrRIRzQhm4pKkAV96br517IXd2LC256tYvkXFwo
F1ItSLLtiYPRt9mQllE3qOPeoUCwfrG3BOjFuDlC+3bVnFma+FpNZDeKTUTHRztV
178E33CIY0VvTNX/Z/KHfab+ev9VCrvXSl8/OtYHRycVfO5rgx+bYKOi1gBfTRxm
A+/PJ9oVZHB4Hj8qG2Va9XP735eQX1S+mv166P1pM/BQdF2u3jpz6uTySVR/Fdy/
XzUtwhynMOdK0bhQc0afPyj5BSYVQmuxFNAJkVEC8yzfKsbFkNTWJYFuBuipMwwW
zcBUJGHvPWnq9hWoDnBTQIBqKiakc1j2qeuXEos9Tk8c6xiY2WDx6rMd3BWJgLWM
VhhOHRCzPu0s7OESzbAtZLbI5DzCTEYiln00s+vHl6h7jjg5HZaGuMvOMPrJ0Ixh
R5QHVedyoonjPcASa03jh20rh2Ya8Y9WwGwB05gIHVaaBdwiVo9yJwBtqiHLPNO3
YmbBDWIXk8YaLopif1lf3Zx28nwuo7swh4ymtqF3qKed88D5NKwJyTUUikRkq+LU
+9qruPAaeuc1xHk5ken4Yf6jM6jVT9YotkzCp29EUi3D8DeO8mcJLZphlxekDm7P
Ez+Esvt+mpfsQ2xLhFNKrghA1VFksacIEC6VD1Kf9miTrbYDFBtqWgtB+Nvki4w/
BPT2qL3ziCpcXL8KkorvOQJhNqw9uXR9Yikqt6zqkRfJ11g7TytfoSka+D+M8Wl/
CV5jqoE2opNXS+uZeg29miQV+jYDNseIjj/8GHNkm0B1Vp01ZSSZACBKTeSi3dZs
a7D+CW+8FddAcaFf/pb3hZny09dtchWfpTJgOCgEbgDujfJxnrec1dXzMBAOg48Z
vc9hp/TSbUmOyJ8wrmAGqnCAudugjwKF94hulGOAEB8YxGIh/RWd7ojmLh8Ai2Q0
Bc8XDP0KPphA/MQjU32jOeErqi+7TDwaEQOwmCDbWaYQgVbeeQoaziht1DKD4HLr
G3l+sV1QxsdXd6oNYt682au25hlBhOtGWprw8FC79+2yXAlVdrFcx7cPPiYCGod9
4ddIO1qbPuJ3CjqUAWuTdfAhd70xv17BJ7ML5G9Lv4cIKRaYt9FiAivMkOLK0b+A
HTNKmCqUNp7HQi2o02mNV9dLb2eLd5kUU/zZ6OUkheq2mDOHyPvfCd7phP4N/BD5
j+gpxQ5v+Aq3gBM/COQBe1hbwx7L9rWsAMe544T85/cu5NFUQUJd7VONH2EdrQTg
EEsBVPKNaY9HYkV9F41DklLXfNxwoxwgJJZg9VS//qgE35WH71QCqmig0/MlPH3q
QZuuuhE2OXOCHVeDAPsvXsFl6u2U7YV3R4GRGT9yqso5D52EP35DrzKWP3f2vbEE
RkBp4SqcwN8+02YoP4SrCpO+a4jiReRzG9VUOTFwPcWZylLaUGAkuAqeJEeNTt60
miUVmQI1PihT0WfYP+hUti0ChWiEI6/vrP4RlTvKdNb+XtfsEQ1nvS7mbVuCA3d8
BF1iNCmevT49ayyULXg8smjMk4sXy9dTfvlsd0m1XjAdUkTvQ+KG3CVChehWh+qE
+DGd+yVaa7K1VkHFgYAZB390LrOpSgNgE2CgSbAs7qtAGfUp9C7zSgfy6mvKNUdQ
C37eGerp+/efHoMQMoVl3grVeklYtQQCLHfyTUa7xJAE8vxP8hgR8Zh1/FIzcFtb
m1m0aegLrIWkW382YsoIyUYpF42uN80NElsRx0LjZSoa/qa/UuGMkJpIYT7qQ4Pm
l8mT6vrQjM9a3aUDKWnGU6SsCZ6QmqmiuLxeedhJTNzYUS/EUistEHqHOAezGYLf
MlzihcqIWvJJf+AM9QFj5hOpK3zIMGT/W1KYoeez16IebTUEXHjVPCNqMARyCbnh
1xehVvn4kuvvk9ADpZvJX4SRJtxrf3fsDUw4YH6F1RSsoJS6trB+B6GKd8kQwpny
9Q5wSXcN99syEETtuEWWRtDg89YELftJrE+Hezvx31YU0YJO4xj567wcjENgY8vc
Cvduqv5OIBbhkczSs9uP1xq6Cquq04KxUppSCJ6xJAoGrtFac1DvrOJIUwdUrU2G
+FDLnJRTTqFQ2pGuQhw2Sa5sfvWrUFgxuVpuyrm0Jq5fJPPtzI0O8o/mbeewsFJn
h7AtDQh0nSCD2h968OEEfo2Uc7MZzTPCQtpy93qwZWg43s8c2LjXQkqSVwbK7Um9
ujEKCZVck322DVBYMEa9Cndmt8pz9P65qphg8vRBasYKI/LjxWpO9218BQQjVaTo
xrHnsvRVu2vt8hRJYVCmRdDOGxAcGG88Y/3bzSDTiK1WS8WpHeuiJ0JGlLYP9NqQ
SLrgoHk5knIt2mgbKJB7Jrq9b0iy5fFFAWFUYNw5NzbKkr/DcGnPvojfT0jEX7Mo
`protect end_protected
