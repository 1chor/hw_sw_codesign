-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ZsWhWGk6JSAMIJIss15zVtYr12e3LSK2/JFHZFvU0c0lI7GZ07tqDzfTG1iWU/Zg
pMIftMbatiKVWuxASIqDoQenifshUkw5bQbw/SfHXRzBGrnP3fGPz9E5pb8o1AtX
rZeXhFnJMxXgGAXXTNz8fv7aHxOxh+tA1yCGeQTFlEo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 54688)
`protect data_block
s2iYKX01Q12oyiJu2+T44o8kR1eMmvWLOe42uqMsfJ0ENB9mOKRT7Igs13WdCoML
yOKu8Z/B1ykSBuQxGbUCVqmitrI/x///MOlZsFTZrg9pKgr/etdIMvMzKQyoclMU
0IirwKuHorBGP9xOXki7umEfZF1wLswRagDTeJTjhlAVEju336YS4Y213W88S/uL
q4FzlogKqKivppnYJHrPMo51b43DQa3EhlR1oKhQRKPxbzwn75WTuD2pt5yyL2gN
5JyzOWlJZYXhyRADOwbvu9j57DpTW9phSwklmVfuFJy7vxlb8GY4GzS4dzoiG9tP
ZwthsqQuqIAzXqSD7acw8NIT5fWeeq608Ibwz+MSj6smP4AFVfUjMuGpKwIEyeyO
2wRwZDKibH8YRiNJTYoXeV3wmUNZjvs/Ecu5wsEY62Fpw0l1PFe+9N3PX/OwrMKl
Kot1AlMuAvb3JO4DIdd4unhkGv8mDMX5NjrLVvjh/iKyuu56e7IOpqdHD2tDJDNo
uDv3/Ju8mY0HOa+3jVs3eH9DaBL0sQ/0ecizr0RAjjdXevs0/8ooWCQxYyrbE0mR
VCVAXP+1OZtNjseT1Z7Iy7ilvOY/HALNn8QukLY7Ghc+UjUGG0GpVYBFc5yBnJW/
/5BHqWelfxsR7UNAQuVzXyQfTQl5WX7qe+GgY+TVv736bqw7jSeI6Vs/s0cDzw8F
s2l9hPbLySVaRpPeeDvsLvdJ79YYBS3/FxvHBnvcrqlY+acm0dNa5uSOG+pGsTQK
POdvjcvEgu7w60ucqOk/B0TTmB9PlsAufuAUPA/Sx+rTqRJm5Dewj329iNvRehjs
1aOJ97NI655XCk5Wt3xsFHUM8eeybltYkTTKT5Kpp87wajZdZJQHyOmbx5Q0Pzjx
RVQoYWqIsParLIqmdangGv7kuKL3w1lZhDeVG4ND/tEVyoKAyaTM+BqeW27Jp1Rr
lyREJ5dQQx0OwrervpNMReHty4Ii1m4RF3pEET71bVk6nnRzeAZZ0kaxjCKsh4XY
xEmChN++IisvCPraV+JbeyShDEAHYT3Fcc/HT5TODmq8pBbhkwX6J6O5YSvcUVyz
ocv718wjcd8yPUD58NGFUsYPujbmFjqxNC6nUAaDNgO4xlu03zEgLdGIaxwOznNB
kITJ6QYk8qM36cHSVm9UZb1YOk60fn0peHIQkJXF/GzXKvEOvkVIsiEmItYxrIXS
UEkmoZEZ8n+PEseFczt7gMNEKXV+IT9oGAgFmiv5rD7tYkqnRAgTnD5goQAGm1nE
vecqYV2haBTRNUTGfPyRGla9cKP9adF5SZMfdu/+xwEIMgAiJvkpAl+eAX7fUXY5
b3sP+CsJYSM/BKOZS4QGdGWckq0EHq6sqrJgHit9w/puVShhet74mxW/C7CuoaNl
8lgCm1vGgNgVPiGUfvCIbVM4NMHAawNNV4Qfu/JN6efw7e63gSmhiSh3AmyDAvT+
CrEW+dyltFI2Ir7tQO6bnhEb71zdjvE4eLkvQYGOdW8ZgpJhvzVcBQk3lJXfnRhx
ChSUvdMg2N1DIGMW2l20LpvvZqt8JwhSxndXFw5EY6t4RXO7DVYLdVV2sEzJmGXa
jc4AaGEzi7QXeS55F5XQw+wI7BzQa8+yRpgDF0Djmgsfw/e1KQUDciBdavJ/U7NI
RdbjvlcQEnC2WvhND0OzfTngpOQUAkqf5lahSRF4jATLMR+a0TL5bMCt/R9PwFMH
k7hiGgaRpRAXqExchbS6l6f8oKdG9O2NDrDAsRUM62bBZDXEPoMoP4bwGiYi/gt/
iHXrlYEif/qjfs4lDdIKtGP5UEXSFOsgAHgOv963fQlgiAF77+U4ZRz4FvwS90IO
oAUO+T85e3IjljumHETkdSaUHW49/kPrk6iZHgY7WdLCw6wKnNvJ/IekQJpTxH97
i0JMivGPVgGrxs69N+NU9LPbmWtOX7xk9nOosnnmKK0EBwNuBkJRHT61zf+OEJEU
IqcTxOyBauCf1OYY7oj1zXBBHDczxsDGuGw7h32YNZuTcjIwbYIesiDx923Rsmi/
R+vzGruQ9nw2X3OaYJ8FR3EEvmbdCh2bPupxOErq0DZy9QYHJPsGmz/8USVq4sJD
HqU4Vhq1wDQLsN+PoboWAHbw+1YUmKrV5kcswDMwx+54yNQE20L89BAYdmHCasNr
vHRYEMpQ/v/vVDeVczNfnPHoBHJxY40I401yoh5SB4j/LBhWqiCA5ygNfO+ojZjO
oaY+JDyY3K1R8uQ41OFotORSOankAqODQI5uQw3giDD+i6B+qZnISJR8ARprPa/K
fypbHPYQupwkUb/c8CclOdHxpKv+NwAsU12ey6n+fSYoLQLe8w3CNFXbM17Czg77
TZQjGejOa4MeOE2QxUhoxH8sbzn4AOKTDMQdxzMFiKRX026Nmv0r+ACkzpaFewf3
uBFmrt+IK/NHo4UXF5dcA0AtPVVAAA2pBAlepsvwq+gmSMCe57rJe+skF6CbxGUk
6KMLQq4IZelRyC/sl3aR1PvexF0bLZENZNmgY0caThXWJph8KRZaNVvr7kuPf4YV
RY/cfhw/oOX3muxe+Jq2zlxI87mZLOd74PzX8ZLX+WN94V86aV85awggY+LoITSB
ZzQBpAr0fUkwIIJ8Ma+avMQbZY9stTjH35rb4o40OkYBSehG+c0r140BqeUR5L4i
h6+oq6cddB+sZ4/hrzC7GLJDFcFPnD4b1+Y3N9oGupEx0dcAL3/nSHx5pWzBlZyA
cnhM8/7f8ImBJqKRNTn4NRvybCFzYO3dLqxp9+bQWP4yZI+0LBVsVMt+Yv55Tfbx
cRpX7teBbsN/+PJnGuU376zYFoEoXxAnhg6rxFDMFM/c94x3VeeCfBaASpTQBVgs
xFkd5/eyUT03eH3r+XtpHl3DVCYGIp/7jEvE+A9OqE007LKFnz7jllqKUs07GCCi
nB4yCyQw+zhGc8epsTbqkUl4JQRFU35U3mJOFdpjpWQP+K0OJcdPvoB8d9TuEWir
/FSa/66a1p9wDpSu2USTWkKPN6HmEFAUo1+lTTmw5AVySxWDaKmJU7NqaJWIw50Z
yhiaYn84L9iClNCXvDLOdUpV7Zy4qGcJjYiin1sr+4Ki/ALD2WGO6p4haLfXAagO
qEfaX4DR8xsCBgVeo2JOvsXeFcprn9ObtlHyHdVyifcmp4Wbz3/aH/K/vqUhyv20
13aQA1D0PFG561o/bZJvTMGdkvgGi3M9Y4mgbDPfX0HJVcHVHFNLKF4TOY/cnzE2
LJq87y/UUc/iqeIqe4AMGvRsW4H+Pc7R77xvT4nc7iggr2xLErT8g6KUTFN3ubGg
PRz5tp5ZXhBV+9Fu1Vsg2qTfQeSdRUM3SSJT79bF5gtLx63GeFouCh6EGDB9QKX8
UfKN5NiUX6dWEC2g0r+EGXTCOo7PgeSCftAeiyfN+hvXSBr+P7wkNLekmqdWjw9u
21gmdmWO8aDu4kcYMJcCVawnjhhtkfEJRU6BgfjFqkelqI0SbRNW7CP96qOresLf
nI1Cxmtd1IWvkOvkUqyUf6ruus3c8oDh/u1s6MwVln/SV8l57kPYmPoSaE9gNw54
q9sQVSLByldwovYnx5upYvVrsGdpYC1mRNyXYg8f3Ie+YrlRFu7c1sc1B+W9EDcM
e7YovO5teaWnllEWilcYTvZqGLnMm/bI3VCHGtzSGbXXsbG8iOWi+yPkmeQS1Jlw
x32eLlnKDYSEJ8cCWBoKaXXQ7bWtinYDhYEAvz+voHsRrr9i/Erz6uE55OXjOofh
Whm8haeY5a1tLSCyEq3wAGiD0C/hCkJCgjgrIepiKaiPQPcXLBfGsEuYOn0rrsBm
ShQEgurG/ntORagMOQ0UrZD0cDfM8LFiYiq4YXphTG+BLAT89gI3lkGfC2wPByEk
rOGfEse0uttkBgXxUSCQAvdw/oToKrn8XtaX67FPaCqHP8k3kB91MOlwR0sqxxgO
4dg2MPs2+H3+niUErgdrclIJ6ax6IlXehwAP7hdC+C0QXz2yvkHmDqgtQyTWaTjV
T+0Sz5OxfvCa33wGoYYStDHAkE9s3YQUrDCtMf1+6HN/bfyettw11jLz7Z/6zuGa
sAgB3FZ6w5E3VYmjj8ofxTNNhm7Ex84MfPzcDo0KoMggbQ8nLY7DFpSDsgV359/1
Kj91RqgdBRhpYcpn70Tcu+RXyOjvVAznYlTAAQEuUrHIQDsCJFWf9rI5RQG7r9th
cHewyLA3dq8G21k2a57VRqoEIwvZFPma+6I5a0dTc1ozKuY+M8zBR+ppneXYD2MK
uDIMMz4HL2FJuyFDfPCcgVgjPK3jftJbns2NiPMLdN0by4YV1K6Ti8BUQQ+mxhT3
/w37I9XrT+9Uxs0F9UfHYxoyVZBhmHKoqmvA5x/cfuhQ2fKuTloLv8Y/AWMmyX5t
R9qn3iypyD+w1AdvYH65/CH/sXey0jTfQ4j6+uS9bB/5LLsX+Yu7lmxLKW1UDQGZ
L2V4FiQGSOPWK2UbHuD0v16xsM92yJ02ARJSfLZBNNv7nZL1VEhM+IjgQ/+SJRq+
GBY7GIjeeaPKJ42sVkY/pXxFVMczDIR1N5dn78kXJrHtsIyaQYLfMQkxo+UjUa7i
7RJHoRoG1ClrJ+/Wowx+dy105WC24c1+wGttIMUekdWO/JJHXx+yazQdl+iYzewl
kHe2zDL3aIQojWTp6KsiKYpMTh/TSOmMLVA++M2GhO9DSj3VwlL+SDCGskvqeoAx
sWn5SMv7ZJE89MvZunlHsvUSAwJMYe0gDDTZ2Rcqfa9h+evdPsjMdCVmhVp569tM
ZrHpTk3vhN9JY54Ltx42F3jxNvYZKkUIHCuPnOIVS5HLOmRr7K1xrilJL8dNm2ow
hgyH1iBxt3C2JcJifquUokUUfz65Sum2VtpjppXAu3uuBJUw4vdRXSdd/yOHis2r
xOrwyEeosp6ApGF4aNjQKv/ZT4yoE19RkW01bFW2lKDe9L3mmRb9RtMkSDxyQYBE
h6jiRu2+0E3zzmm+aNifzO1AWVmUGAjQH5kpwcLo3TeNWMRb6zz3oERMRBMNU6iK
TTPx4WBesUdeJ/lis+oS8vkBMhxoulTypDRxRHdt50+yyuk0skhR8hX4+SRcju2B
we8DNc0FLgXNkS6cHTWf9NIBKDMN303WAl4gvvQkro1UqUeQRSONCxiEKPaA28T1
aea3raNN4PRzdFO2L42kHsaqJOSeUuvsUkWQ7usB4Sgbw7Yot64j3MEb1Ft8+/tH
9VLseqVTkdeCTk0nAdcg/5u5v1WNH++YkWCGJ3fximQoJuSe+AGewB/WT/pH/1M6
kV/ZeUKdbwnMg9z0tZGECEip7iSuP5d7MNaYLhC1n0LhWKvBv3PJHD1vhIw7NBgB
M8z3WIuNEdAJnxllDyuuwhkD1dpEOSWEaHRJJ4mJYpRZ2+VW7Uk7hqx3fN9jAzru
tvNZXiMT823ZKweClSaW15CCmvrkDLJVsEuArfYKhDpKSJYD17ev6om4id3bSmhN
DzaJnmLHUToaFbRcw7PQmHRNHazR1mN0wEmm05qkNZZ1328bivmEuJNPBvZ4e5ws
Tf/BygLUPeuI+CviWb6AFhiDt1OravYIwIFFlQOG+TSsf5OYySKChClIjQyn1FQG
SBIOqp0SgRQSzS5x9ayKLr7QzFhOXJAprLTdw880Cfpsl53ScjZ3tGoLGjAtgpFX
exMBrB+KDOMLEHJQEzUyLDnJgG+f8GCMpaVNCK/o7whmBm5PHOlBEMLLmfThHjP9
tr+FbMzB0ROdWW4S/a4+Znaq856Gf7VaV4imc8taHZNoqx8hqlM/IGGd+bHrbN3y
CRV91ezVdw4lugCmn4peqYtiiH5eGcLHKDB2423+ZStQ4ijxYHm59KrGS5+817hK
3DyfyMfrWzFzu3IevEok9KolNoHUxJCvYDVGvNbUJosUzACoNXJhEH3fLcO+b2/c
Quqs2coYflZV2BsroX2IJNUH0WGqLfiXB0MYreNpqJi000h1sWKDY+nQqkRJvKSa
b+fq+cpRc630m+imtb2cR0GodZh1vv/1TZQOturVSwIVjx4TDEcrcfx2NFpwOoN/
SFXG3OByOuX838CbfgxGB9ALs+KidpF/21jXFiSsSEEAzk1+MfrxPQfq0dvVA+2n
I/zYUOsNZWtfAU3yLdlC17w1XEipoq9mTjB/F54ynq6SI2aS1JOwTwpdjMxTWBsD
NSqxe24NwBYakazgSjjF8Fd+QHr9kPggvfUc0oEu9OLryRsjNSrr43YoFAypbFJJ
JtWCspDUut2Zj/OGBV/TegFImwJg2vinEY8cIqyI/FVVWvpYyM2KvFOgAKbwrbxF
ZQFZS/WhQicspaH+aCAe/i9bsC/qI1TO3e3mY+DflRTcSMVSTgW+EOHfwsjgofeQ
VCiz0HAVjdAj5p9LPUHupYrIm6sAQAqQBdscHf9UjZYsTPVIRiX4sCpDMZoU89hw
0RVbYGZvIvosVatF31HUN6OKomF7C8REIO3mT8CixJvloeEDP0borWQvvZei5mEn
eKcTP18FS9OMM2UH5VgUKrjT8P1KDgJGPP85uqbUB3ZMT3Gh543QdZTC/c2KXSpG
1SANFDSPkLBN5Zsu9TW/eqHFTO8KFNO9JI1zwTvaLapkffTPFrjwtlQPNNZgNj9d
xBaRUeGKz32Fui7pBVrQvdMzeBQG0akpgSni6c5kAdGfUMS8m3OziRnSYeegOhvV
uqfkyvbK8xQ//ddHk9o4DsaSMDgf/irfR00ud3kwa0ykslLrQnQMfIvOioUk/PNX
H15NVISvkkRIS9bZIwhLHJlBGb11k0Up2nEP0AQpWEIYmvwX4XCF36rBGbOfktbv
Qmk1TIMuZblUnalUd3k7NxyjJcjH+hgb4J6rsHkOyFljBioCKNWU1ubHxdS9/I87
nYisYB8NIU3224Loji6Olak5euUaUskE+wtOWzCAtpYrmOxFYSWvxInKif0z/1V4
iPSwxiTAcov3di/SXMkJ2SubUCg8LwjJMyprImrDsKrES3baT8dfeN2hpb6tDI7y
eaigg+vjJcAyd7CfEUHG0fDthO4VAa8axWG8td4YrEwA6yP+1hMePg9rIHyef3bO
+WC5SsiSy/GnAvdDaLK47rVN3FQG2DZ71im6dtUstrKJQNjLhTm4plci4ZIPst26
39lYSqwcYotT8FdxCQ2JnUMUGeB/Be3Oxz5GXyFqYM7TcULkPstYAc+yUAtWW4hK
MAqKy+RKH/bgK3FSWd9H2ba8rMZSo0gzR0AB74zGvxlJEi/Fr4sbdxGNZF6CjWmY
dvOovYUXbBG/GPlTskKyTyBOlCja2Pmp4lSvPMUHgRMoKf82zKIfR4znnnE27wm6
V+K9t8cKci2CCYrb/Sahh1w8Gf98xGmyiP1BSsB+iG75RoiNPbRzjC1nnGVb6KRz
HpJ3NkQ+ORw4EqJGLr7gtR7+xJFtllBedj7EAX52YigUh9uxAOL8Vm4VTTU2VAAe
6Ulzse/WbVtPW2pf+CLctCNnytkUho6NeLm3NyjgHAFUtw5KLCtL9ATN59ljn3SJ
5y+PKdMv/tgIwbQFI7q+U+LI2lMFZuHGxcNCyyv2zIm5v2M/y/Qc5Nk9cHG7Qzv2
yEdfCB5PWGT8sNwog3xAUGTHwi3svSyx8yPIAUTHmPSI2fPAaMbMWfiV06rxoGKR
2VvA2ile01EC25PhzlHem9ujWwwnvcB7BctlzU/2qe1dbWE/YK787uyTKVoXku4d
JXRV+3Cf+aiHgsRXkaIRKUz4r8cHhNqyOhVod4W5oazHkIOQkjhEb5U4l3OXH6EA
1QIBIXxUgrNuf6Fl96lDXffOMlP0otwqxUTE2TaQHHm1q94GymVmfZTpfgRS56di
/stGNGSp3qv8y+gNimcGYkFdnJ8HKTOTjUXCRHbKdlk5YUUcbuoleDwyKOW7xXc4
Ql8yrgx+kRraLslH2nrJD1WDLxTkWJitOr6KuZg5rr8phPMQU9jMBdBoB+HDz0m2
pAP5OVxQ42EhJY4OMysE+rwgxGHPOILwC841xZzLCU9TWrlRHJJt2RectARs97/U
XcDZR3jlO7wF3B0b2g9t3WSEJ1QkPxc3CxzzP/vgyVGeXVgR2wvwoOOm01RVn5Jw
8wugredJ4zl47mdTAqiHHaBGK3ImhZ8NP4g8ISLacTB3W5yav/0nowwb4znyvJ+c
u0u3LmAheZWCwR3dFoEoLbascEmV4Vi3XhJTAdb9qhiqIVp1FLaF8yQOm2TicMHx
tHCwpdaELFKI81rJZBxY4KMno4ScxXOl83KkEXm0Hzc0BbND0Ji0zF3BMhRrpLsM
c5sOxCEIFLTRIMfWVFXxnT4Zgn8F4GSaKyRw1Avn02dlhNFRqInvSiy+19CeyDpB
LXO5mSGinFUzP45aY2o0JhkomD9Xd7jsoztISv+iSbaajwFeqHbPfMAQ8oBiPqGB
G52M7yuQBJjvgTHHf/73JXH+quvjEzk+ry+dqm8KC3JvO1aqZsXRiNC5q+PjYoyb
YW8a2CrE9008+nbs2dScIg0WzhB55saXBortoorgS5GBPukN2QgFrehz0jupZ3da
HptuIPW7n+6FYNbcNE6G6fUxgTj4mDLBSLvj4KbuxCh20sZV6kRdrpwtuuTyyDuK
SsCu6BZuHjyHvczlDt7dJrBdqVnybS3gxyzwTX+f2L7lU89uqXY4OWpgadxFObyI
BlPbzUZOq6wJmwdeerzIZuVvlbUoIa9z1NUP6TROZVA+NRCP+qDd7dvCRxBNMfl+
HyOfCZgYSyurE31iibUUn99b1D1O8rbDYdPCo/AywHDjf/migIWN/5l21ECeg6wu
NIaUD2h1xukV5rfW8tYiFC931AvX31HDaf1rdV3BePSVzd1FKmnpjrDJyJqDbMUZ
MGBzSfFPK20MavcINBRkFYDHzlqoWkjMVF88kEM2I8/FG6WuiNwE/bUFwSsdYFbv
morFUThpCZEX7+BpfZ9xO7LUILVqOzQgqJPxgKRgjriPgifqORrfOzfjjsGJxcPe
QDq5SJevu5Rc6aXpch58LYUClF/GP71dRL9fpcF6tcwvb8cP3aTlN4yoRVlaku5K
9qcjkGboGINN1QFoZCP9NUPVYYmquQbsRezOJIT5kBF74F6KZoNo4q43iMGkiscm
BM3xRgJbRcP9iryeqn7fyISxBVCdsO1snzp+QPf3RPhTbYv3BqiSeYPGAbSQi02x
FeLd1f1xKQGXek3/Jy3DVcAaAV9E/RvK1GU5hbcMMUIp5ChsGQc8SEYpWQklexdK
lT8vbNL5R3zPMQ33quP/VYKdRGYDVu8S9LdGx23XekJhJWW6DCfKe7/4X10/ZDCX
dZLiJsDOxmk1BWW6nDfBVETC3V7m7bF+QApPGQEDjaVrj19RrmVcAEF+O/RgSqa8
EztniQtoWc8m2NiwaxWUb1AzaNZyLxtbXvJwwRk8NuW89HKEEvtxj9lpGD10T0Gk
JYfyo7c0J8Rsctoso8pg9QPDhhCzuDp47OqU2L5Id4UEbN/nOMfvDx8YZcGHDiV+
/A+1Ob9XxkhnPceIJZsddMUbMZOMOb3d+loYZskhDBwJBP88sFeEs9lJlZgpaYCS
F9FqpL3PBmFLrOR9ctx0jTo1bWaQLt0DpqtHEnzHhZNlr4kShRzChVArjp5HVHaN
e+1HdKKIniExB/MTbPyJUlJBn0LxY15pF2i54yFfBsUDqKiPjdOwFDrIUrzJnPNe
14X/36p6iTO4OUK7kteuP8weMjpyNEMA/K5gEcte1FpiGKm0K0ETrqA2IOT0nSfm
04HYBAhKhD3cGuFzsh6+JSCpGzzDcthGClTv1f8CBo7FzNTQqspe7ADlZJg0CgNh
h6YOjXSMe7fbDeyF1heC3vVBVn9bbSLSmycWSJ56L3r1nDA5Odx6F0kfCSVPi/SB
UjJDor0jU3Jr0grIR34wSAGTGZTxAWOa92SoIoISjPovbqb3M7poUdNhWdO/3RPg
9120pyoP0VVBgfx7H3dIJ5tkIaMe4GNWahQ6B3pnKvF8j5sO+OW6AJQsQd6J7RO9
HEJh1X7LpGlYNLEcDj0+LffL74pZaQ9jS+u0SMtnt4LmdwYwN4PVEg+R7tpmQyJ8
am8KjIAzsCpEvBKPsl30jAn5Hmf9iHeS6pJ7VGjxPqQv7JfeEYzZH4l+CzDSuaWE
qF0eee7Tz10UzJOYn1BkicvvKpSb/Aqhe+pyZg9dxPaJZecTi7UvZee/WPxMrahZ
IdR4QFCtgg0xpcdxa9Azjg3QyTrfyQQ2SqYUvqmfygLkTtOs4njINh/hd8x9UXv7
ai9suWFJ792tmwyhP1GJ5qwAtnkQ0gv6Cvd9YfNaks+lf5fSnr2YmombGwjfX3ik
aks86Sx7CsMS0Wa3XdZvng6aihy0Sl73NllMyBOSEJUpoN/q33jEVnb2BkVeLm7g
oA8fEHVm3aFsWnQwcVRitELdcQLAuAC5KuKOB1nAiWsqjRgzG4mceROVjdYPRUCV
o65LDBdViOzW0Z+ec42dREImS60fbq7u2UJVfO+1zyLvH1hremaqnoVrnlnfCl6i
rVQ36IuZ31n5wTU2+4SqJUPCYKNUSEF30DaiJZ8U2Cm2VPY5uXxuR9mAq3OenDMW
EBqaY4DEgYyGujZjvGVCoOBs7eSY3R0RXuiGM2YWXpZhPyeklEEIA7CowSl0Mj2S
Mq6Uhmd2ZBtxAvmYT/CsP0EAh6Ntfzo1rWDfLjC6zfHGRX49xOsfXDJd1RyjleB1
Oh6jHV5HFvZQS//7/iJYlxY2q/8CaKqyIagfeZQ1cF49UQJMYPBc0Xw9wavqneVO
6Ug8c9KSiopHM+4VU4zhss5DgxPRfiyKcVDuBjdUf7lwv2ciNBW4tY9KgtDHTHr7
ftrdR7ix/K+Tb1HwdEoBlrdPPMq/fTSG3V+rBdWgJSpI9kaZv8rZYEgttwMuyipM
yOCJMaIlK9IPw+8nBOln63ToewQ6NgW0F5KKPiRcuMDXnrpH9Q7p4HoHLrX3NMR/
0f9finx7+sDoOYZwGLFhSmow+uiWIJNFTZtD0hrV87B8fNnmmhUn99tv20smWr9b
9QURypXyXQ459hksA9vDaerLY+9empMGEof1FRm3QinGbC6AK0QZVrAKCc6xdq+S
1flJtrQgWHh9OCNKlBnEqP+EvMBDzAsImIDCd2YZ77jhVgfCzOmh1HAhqJe1l/xe
rhVjgdKUqu6068d9GjYogPXVLOLHQF2y2g4tYbQRdPe2peAIIsC5BNnRLIMjNo9B
oJLNUdNPYLm/JxnFVZhlnzqDJ+MCdD1XAtwC2/i9ZqkR3OzuRBVs+KEWh9fNX80G
qh7HMa0oGbWW7PNkxOKxEnOA+LSq85QFRGTqXc7VBHiOeL5pmnoQ5XjHp+LJ9493
N2QTIbPJwIxQJc5YQTJqels8AhZuCabetfJfEUKCXowOnYYFJ6M9IcWbpoJAUmpd
ze7H7WDj+6OVkyumdQeUTiStAYthHWzcWaQxbXkrl8TyQaFR9lp1++hv5X3hWiIL
dCTrn5S+JD8nBEvyUJDV6kGawbw3h+9V8FMPJl+kwmUxXj/DSk73iFD9dAsKNoQA
pk7ee+q9geTXIXYGmS//3eOnXKuwc8NfZvqOHZy38XWiNH3nJfd/P2jSxJ1my1zv
wb07zDmp/aPKv3d2dnnoXw8hXb6pODYMf2pfO425eQSe7jffc58OGal4CY4Gpezs
UprlAEaEL42Pj8odvNA/XEHQ7FF3D9MxGETAerIhH04G47MQPOKQkx/OL5hnzsGX
AwUSj2z1tGWHEDTORK2FXcZb6p6C09RjraaT2fQxcto9oFf22ivyd7qVUg6kB914
h1K82SwCHaC5/XSG1zuoQdvjkj/59bbKMTq/k4LawN4O7Az+tEk+L8oHYuUEL2HK
VhIpxozrO5i8KrFBstfwjENSNBziTtEhSPXi8AuayJnsXnfGmQKulInp/wve0vjW
O8E1tU7Uqh5W5QKS0CpV2oNUq3mY0KswklxOonBCUWYNNugaeNLNosZlV6Y2IldE
W2EPmxdJj7d8ZNSIHdNeIPubiolTMvMcn2bJBv+dsgOYMk/rndAZnqiHsqg4RVHI
wpS8h9FLaAIuY/cloKAsxwcmg7xLJAezr6vcwmZ87e+DC3YMYiy4fQz/KPotGQMU
amRluEQajyxODTPXo5GoD/oOgxTGfKiYngj/8pJwRqihXH29Fbuys2GkeHk3SGUZ
1g7gFEpRnlu3Ag0zeu1ZYF65xjmOHah3VEX7cljFDfqOqX3/g8ICOjRlx88xrOW7
VSAxxvLmfPfaPqeKqD/+0XCIZHyImg1Gqs83ty8oSTJPtoDLYPeZyGxcNumYz8KH
faDvCJGhx7ddQ0wWlXKvjAaTpr8uMOVfOf9ZZW6HFGT44DUauMWKchzEQ99efs+m
d4B/0iAojut3E4CZ/CgB1JdidZwBNXN/y058+UAImasd4zD7jyE0zG5b0R6km8nM
fhyqsfxdxD8UpSvNaB9J0f13UCD0xiV470AlzirTTqjMWe5KQzIwhH8kpSUEiaE8
HS6q3n7Xb58yD/nLVuqv18jYp1AuLofWhCk2zwgd3JRjK2SE0enqnzEO71zmcht5
BFUN34Ij/RK6gsltVIOGhWOER31jt0LgXXCAdVan9nHUTfcB6zM8ELCQ2HlGdHze
1SCETcVMhvkfGiJrj8wJIfXigPt1r9sydTCnBgBvW7B7tFBnoGGHbhz2PseCr/by
u9ZkE1/D+yc9JsO0P4/IAwYTpw4JqorG9yCQHTSkRnV41DX4Ia3GM3d3wRvtrA0p
udjRMsdT28PBlNuPLUlPrOTBXMQVJSqiL2duHGL2uIt6Pp9dyOLD24BOyW14Ztkm
eDA9st48ydyvM/MAVbAL6fsI6q1UC2gTdTbI8Fs5y4CM7WIMoEK0sPbeNGru7mdD
eWXbCC/jZ9B9/VMJ2p/lRAuZC3f79GbE5bAeU3Y62+jMZCXG7CuoxUMEo5YPXlYq
XOs4JGjxkkoBMCc+1E3mYtjpYN13T7TVeK6BaV89r+LDGk9FR4105HZadGPjXnfs
j5f0/DVkQeH9i8A8T8ECdKJxGoAHLGrVcve3fvjyiMlDrk01+UHrJY1tphDlcZP9
ibfmGCXHHjWb2Q+7d5sfXZEOVdqBSjFKHiTI+vHA+IUB1ehu5CTGgIV4D3WFKjuI
yE8Rz5bTP3EOMHZu4ke0/A2VWgWQ5w5yofXvgdTAp9ubKERSlJWIk5ZBwGPIvl52
9Jdzhx5ErSz+4p3cksiMdWlseM5qwgfxhRqLU8w24fktlZ+UV9D7PpLb/1gtaeZ2
iSuddF+qffycDKjazYuosB1St5XVr9JUJDG1lVROY0/T88trE5cQ2mT1+39XJpmz
akhAygqDE5MNLmKUnHSGIo4DMWXepXiXB0wKDDs3g57I5Ns/q3Tgn76XccmCDFr8
2DBguA8PYMbwp/JosMwWlAq2BSPbPa+9r0W0gy4Ln23Q0/eEkiIotpWbe9LWaN2W
/3fZC8/G4HA9IMHyrV7Tuuya6fhK78qXjf4LxQuIG/hfuu9yWKAofdIROsoTYbfz
aKVliSJuwn2kWdRnMFhKvciWMxEPrsmTZyvi2M19yDLvRsbq4TjWCc7KiapxOZcQ
9Zbk2dpUvCepHIWcHAtow6bb/Nlp9UvfpV0I4XK0vnA2G9myKgGlTPcOos4C07SN
k7QzmtfwLzsIo6ljARJTmj8nxf05P0u+8JdDTuYgOP+V3PJcMpyXHglfYJmrJxWP
bCkEAsT31TAtYw065x8wgbtdwAC4NZNyUso1B+nX+tSGWeHIBq3pSYPLxx4K4+00
c66n3Un3Ezas/NPV8fqeoJ0H1Az16ZOJNgrCmy9H6Ii+A87ZIU18+hNZMgxkWta5
eJ4D1H2S8+JUYddYMDVDfCDj+OhOc+uGaJG7K7oZv7PGIF8ZAb7orPvnqtlR6uzU
sXBTk0n8+ae8racshac3Lms/tNz6nRPQKTGoySYVF4wbS55MtCYY+UyBcw+7TA4v
RPRxCtuoswYwHUyPblERfx1oaZ7O0huvdqXsQ+89MIaQScVUUqaFYukfH6XZouw+
R5dRd4OVsZEZ0ItmzUmH46hZ+/Sm596eJ94macV9K7vEs6tmtvQr3VkNcb8QbLIc
+6uA7crIVrrzf1ain7P8h0mVd1UeK22/Vl73A7959rjuc2pvzQ1Pi4XylsVxgECi
nqiLAcpznTg3gUvsKGIFUlVGIdXeo/ngCSMmAeXPM8iMLBECUO3Qzkp/df3bKaLv
3eAV/lJdBbwVeS+rYBOArk12TY81y8SwmbzJ8iF07S63fqRpImObiH1fitqB89Vn
snZxUgdBrSl5zRhFgjEKUJOURbqved0wzVq1XuBHoNVutoE/v/wF5xLW6J6nNd5t
d4u7NRnnvUT0iwVhr3QLwk4fLa5XVgJZGsfmd9Zp7TPdjhhokEM+l2ZmTP4bwfsJ
FZgWhvl1bkFV/qU2enIbNA2cm7zGIQLL04RfHdPX3ErF72ozDODYldTdXecLcCIE
mgmLN+4jNhEMR0ly4sEV1WxRuDiFtYof2PEVPWIqKGRKOxBC0rbIBJxhX7DQ5Rgq
t1tyZw+Q1Bv0A3QfbOwfmawwYFpdY5uaj+LNlXwKlP1p4aHrEK8De686RIuTijXv
jw3X4A+PhMn7jWtXcDPMAHTKMJqIQdSb4Q+ydCtAfzvei6l5PuYEU4ERuQkTKIfm
WOPmNYWbrU5HUnvvAelHzGJMjA33YBmfOcu3Pcvth17Xvax28GKiC/kOh1KjR+fy
unUkxamXiQKv/4gOdsOSt3HHF3cxWCsPekNS6AZ/0fnOF42dw/QFZGvdcSdL56h7
sg6jw/XXr2Jl3yN2aQ5HjhLQGtmre8r5nCPtXU4+j3SNcroCay8gpEjWs5cwCJjj
jbwT5uMc1QUDiI3rHfR9KfsQQH1DKAR3ANeScN/8xjayqLKkbqGhA3/DGwE6xn9H
bj64evlD+dwc/7xqa5XXZHLA/teL9BUtKCopTv8mvYg2much/XMcCXKbxFxMmKU3
mJXED+0+oQhs8XTPA1HRprynV5ySRXT9C95glN9oE8tZ2/cAOfdQ6MYunPt6Rq64
5BjVdR4JQEbfMOLbHM+L3A1f4HiT6poWnpqu53WpuKHS8rvzgwbGVQ8O2mvklvHa
WLpzusKejdMFtCShoHE7/cxV+CReb2VNgCLyXWV4cAHbHewRUUNX4LVLzQqvMeTL
vr52HJL5GHChlZw9THlwlWgFDBRkC3M2nya8KX7p1zouwoc3zFw3d6WAsZIZD8Y0
7c/x0nSvMXhu24sq+EgI3z+2YzJc1VEVtLJHLu2a+2WLXB1qCs4cVx+TVz8+MhqK
+dTcpfNT+LLBX6k9ois9DZZFyrV2cbNA/W94/jW2/8AxYCt7ZXKnsxjIez+XUKIK
xGEOxhxFeiYl/gsQ8ObcwrdvruoOTKYFJRixUqRGQUTgdZV8WZjuPKeUJkX/kRfJ
BbTow+klbBb0IAg8j5JLIUysT2G4duK7jBpH1XdR4Znq3p3uZhv9S0C6vkqrmCfr
0I0/wbhYlbP9XtySPMDXPiqVLUHHYH4GIsvgtsgTdX6C0+C1jKyZq1mTLUL/Gn0a
1FymxIU4i4Yb7xN6jG7PqcNPg/7ahQPCK1x67ojVsrn5XxjSDZZ9AoEEyvkWOkFc
3/hczx2tcyF490rSS5z85cfxj7V0XaPi8KvahPOGj8kwQyqejY2Nk68KwWIJJ/PW
4WxAqpbILYmgG/1ZsCsun+NlZZnONc4J8tdcGkyy72ko38O9htVfvgYUuV0Vm3K9
pL4X/Wso7oq6gfGWKV8d6k5kXxuoR64cOMVZxdG3PM401EuBBE5ucW6qV2xn/iF1
LyZ/4ozPcNZNoR8+/HnwFIhxQBw/4xrca8dZjhF703Wfmt9ScGfKe+GR6mI++W/K
8Y5DYHuPV07XAv7RZUDLPt3jYd74oKyYM3KtOlmVWNmF7PPPpKksU11wH2st0mAI
TO97oiCVwrY+rb31KAN45nNBBQtbb25dJLRrTPFCsrj3JyzJgyYh+PkbJQ1qJyJt
k8x7TJARSqvp89D1Zct22MUDjos5DD8yGArQJhFhkM/GOi+5xcSAAjtpA7GcyyKT
HxxQsqAWWfQLfw4/P4iD6XIHJxACO6BnXe2nzrD9AQNCbqlH1DcxQ/Csc4OgIjJq
FwjSV6ZUvO0s1eIVmxchw9rLbL5LhFCy//kdN2pFIq3IguQLYsVEqs4ZxnysxpZy
e+iFwh+c+bkeVE5LZjlLBAIRWwUbzw0F0AjOi6AcXbpLPlshYJfqjyLyzhD1dnZq
5Wl/5OIGqUqbz75/Z61BwD3nzdptH2UipvRjHqYc/A4qgJwZbrwY5y8y+dfJyyE6
4ychRGALCuqz3irT+Gu48U4FZzxuh32cIp/nqfRSX7YJ+nqDS0KJAZ1HeGTnJ5oO
qxxETAm/twICMnnTRYvZ+fy4BciSf4u/LNu5J0XpOTcC1kfFLrPXuj6ypvy8JBZ1
QToBVH/koEIAJYApMavQ+ZJta3bttqpAaDM+Bu+fQupi2Z28ZhDC4nHmDPqnfNUi
UFeDAseYbnBLH7fu8Cu8Y6I1EQCQAKLNO/Zvb/dsuUxgU5cvkACW9+bGebPHEpM4
8dkNElLrlXGVBbPOEoux6sV+mT/SQ4jsvR/F2b+q0FqJgtSrWvM3aGUzQBNiKV16
dXgP/KfG2x/79g2kPNSGxDKOv3lnnkwdSfcRgBVUBOwpJApXF+MkzulqNp3YJ4dc
vPr1gifpXqu5Mq3AWd8vi7Tf0I/6J9H3ppj0uKZx7BlO7fhxrw5764ecWLSEUZNg
riThRprLDbySpHf3gJNVV9trhgdjkf6vF+P6T1O8kVQAQxBw/v/j0/Uml51uo1Cj
+rVbNiQkJgNgtZff+7mi6d20qv+U5wROEVKp7axy6PCidk8PvPDxzL4diwhxTfKB
pAK4miHrIuuJwzo0TBhBhIFWHYM/pvIs6pnaq/OP1Sn/s/9cA1gY1MsOe1cAAqa/
NY2KLM0uGFheit5pdS0JRC68nm8btLdmETTTh/kpLYCXpYGZpHLyVKYhvFDwINVf
q1w8G5Y1+zpCt7wWuR0Nz6f/ikXM9cxNbm19Vh6zprA+SAEQP4Jt2JTojJJVE6TT
/HydE9zSbLiKMxbNfL40hCi1fnnEokuD+eg5gVCd8+havNOUEk1pTT8FgYdCzNVI
K4e35PT9jdUQmbIqxTrugAvhdSLGxLEwXy3YAUdpDGm6Km7XN/KOSo5NRRw/agEP
A0ll0Ll77nrqvAgV9gU+MvrcJogkG9XYqwqA727tusY7BrrU4/6uJMau5T9DZifx
FZ9h4K78sy156wwzuwVK5pPggKlQ5PpguVjeyNKWzWWZEGhlESKdHZI47DiiI3TM
vHY7Cw+btIv/FaYlEFCojykaMWh468OgXQOPDb8paJ3I4B7gkI7bDro/gJE6Q8c9
iYWW3DAotAYhRFxKEUVL+B4XGd587FofR6TbQ06qUUc5mT0gV4h9X/aWKwi/acAM
+T1sICdLm6lyNFzzYRLPncNBtaCn/NRzq2m9+dUwz3E0n9s3B5VVGrAqZxbDoodu
d8XtfueEHwpu1ulacdGfCcZEZTUZ/mJiQRXDkN6e/hRx6XYENgXID/tCAuKdzKyH
kCmvGfXltounCIdGhcsCHEixwQhK+39SOFNpq5n1pzyZ/UKp6FyDA9FCHbe1ES+P
lN+u455m+1Dw5wdCDd5UmXFQgzmOfIjwNDY8kJHxVTPWUMADz/ijxPcDEfic4NBp
AGgYb4fO9ec+CDRzaQ1+u4Qi16lt/kZ4n/dPw2W5J68Rgo7AiVL1kI02wI+uxHIn
C9yRy8isJ2808E1frWdNyd/ubvvq1y1HW6Qb4xqbAkZhax7XBfrq4QVyjc7uzge/
JPKwm7IyEYwghacHfcv7PgMAL1V1kkAS3pgzm/63Y8qLOd8NLvvxBT+dre0dxOhs
ss16Auu5DW/egQdfzcDCbFM0W0Eui0SZ+DWoOEfxIv9rwwyxPHoZ9LGi+vkfsKAg
5FK0n07yJfHcPEyZV34mn8wG/H81N7YgG3+O9e+GhiJ3u5WfJXPoxdVvx992iOeM
MLkgQ1ROZDusoEY3PBtlRLxvchJ80t/3Hdkp+QW8UFRctIO7RZ8Lq8g/I4Tf4n8T
9pHYjBthnBfwcf+vn7ZdTOntcbkF064E6hiktf7FluPA1dClLHnR1OmA8XM+4RYQ
cTTXc6hy0D8o6bxU7ry4usIpoxZyKy1w6qIcgDyuAngTOcALza5xET3wTlXMTLSR
d1ATkpHEqfovSTTAbMT61ztHipkqz98CeWtzKVPXzTFSMFjNrvMRujzjdgfR14sf
RTV8u/+w4ppEpQNFI7CnxEA3cEcJGZBBS9J0SPW3jz4pA7sqHW89ZKIdTozlaQY6
/odZFxoFWnZWoXqfz58fPPTAa5aVsBF6T53OQr6oeOds6IRG7C95UAxJ1iRGIw6B
AFRWxghc2B/TC47mKO47/6OYXdGE0IFrD6hY95d9hMyCjy7rvHLT3YCszwiV28DI
t6H9sHQIKe9p8+rdymCtHuCz+pfUgYcE+KylvF/wD4hGycVa/CeMJJVVqI62j0n9
nO8L2p+IikHqrJNXbIJOupqUIApHLdDtNhqsRa1du5QN9WSzCI7vCPHxj2G9V3/h
ZJ/j/OK4S8VDk36nGBwu1wdC3tUW4GlmgAFWhthNTqw+1smjrtcWwSamvHwEETEM
hkI9H5V1eSGOKnX8cMyUnwko6Drm4YRiNTO1i+FaoGii8dsy1OSJe/eXYgMcTqh/
bNAs7FAcsSupmbGJTDknhYSWslxq+ibHfrmBrtormnvRGjEWH/2Y0UpN2kfs+ZZc
dgDGFmx2RDqDHoXJwwfKKqxvfJGU038LeJSFR+tgvYqznswZRhQ+YyaI9atET37H
r3RtRIIIwpBes1qEE0tPntHihS3Ov9nvlx80bGO3v9mBNXiWMabFZ3oGldfkKlIz
AhrQBbs49AVP8Dtbf3qCO1+vPpriKSWL48CQm1lMw90cnAE6wZpaqwQXu4uasBnP
wQrgeOCocH3mP4hBsIpo+0jSbsnI7WneyFanP7Bv0PKESKSkOmToL7SzDBDCwhH3
pE2sPurJgqiABINnz/F3YQdZIfIsyUG3mIcaePNbsOrb1loBoAs9TsBxnrPfdyRF
LbHX/+N+vGRTxLMQdzI0c2onzvutJ1QHMHDIohkTqr8bDrvqGdHRd6FzmdF0u1za
QOLRP7aSTwytXaPBq4BcY7cO+Ja2rp5d4fyMCM3F8LoWln3D3pW95y4Z/sucrviT
TgCvLMYA9VGx0ag+NGzxAwGn20QrqDumXBcenoduUlDEaTe0uIZ1T0JDO2bBHcDW
k6Pef8mpPfMTFQT9yEVEFZ4EMTQeORb/zu/9qGmerB+62rbdbSu24hkr/dEyiWEx
bio+2hHMME9zQ+cZ5L0wZRxJpGPggkJI0FzwdpeGF5vr5li3AUYMIGmnGOk5gNYv
LhWaB7TOzLxeHKenm+A0Okmn5wnl0TLHeWW5/ivrVvy6Wd7tio/aAgnms0PjMb7r
kpyfHlerDzDo3u3TmPEpo9GUBLTNrbRbUy73MYQ7upQ7iUYHnr0TgE217DLhliOz
26egomQvqj18dYJ9QV6D5uB6D777zvGXFcOoxmN/u849NK013IdaYOdePMkU8q7a
hpVAPntMWEPS2JQEQq0vQzVsou4j85WGQpa7TMZpPqkPpO6RIklV1DmOH1Ec5CUe
A5oUwgZ2DZi5sgIm0VaTigUoeBQkNzspJ7zSDIt/hjWdRUpBfjmbRnmPnJH5zMqO
E5X+XOVcAiq9zB9Y/Pw9bIv+bkx/CJHqMJLTV+RvQBFHQuEkonhDVHDZV2m9G6ba
CwPO9tpZKawOpBm1U1k07gXZwLNkP7iyJMHONlYEOHaJzmWAkmMk3r1nLWiguMbf
I9goAspml8SNKYLd1i6TspZ+urAH6/GwcNMgf2pHXDyECdwYm0FAaUmgwxBewn4w
35SZ4IfHLYeiH2D9O8qO1PsWYDdRLlGjDgbUzZiAshVxpGatUvjeWmj5xNw7ej5u
n7Xej4cXN8A1z3mbZAB9b9lFarc23cM9E6OMdAvoc0GzF936klip+iEP+3hkHWNq
DS42PZazvwvqzhbme96q0uEZt0khxmR++XLh2KG5raZlAAopTqX6qUePqMZdnd9B
LC7ch+PxbB2hpu4BvkjE2Kzu89Gjk2Nd4yBGb2lc2hD/5grUUYSv2DXh7PXZ0WL4
Rw3B4LIODoJ3gt8ObNPxzmRLWGP04aXG1e9qJF1Cwu114KIPxfdeq10bMNg0FXPD
0VSWRIstPnZhj0KtOqAZCOtRyKMCUsL6x4aY1I7olqmFGFd1gPF4uNkIURJVgiBZ
OHombdMyMuqymcCctCAmxLYiB92JJ3VMhgL6vVSZT2+sorkblDSY0nAJ0D1/NEbK
JPW1RMmXsQt48IGBxUs2w+7+pXd3weYNqAGnb5JIWwdCKr4tTTr9o3tzP4HjarhC
fuRvzx3g7G5uQjOVYrz5qJ7pA9fbeEsILO+ixSUNaPLSV0QmS+CifN/HuOqJW2pb
C8YNrwiWVyQabpDvViILM0ivRF8tz4nQU2nKA2LqwHm7D/4XA/kR2BpLsyGvPvJF
lkdpfdTnbYKjQ+/YsRYunidX22K0QsO1sHPd3Zu5Zk1G4taRAlxk6uScJQIH4yW+
ZrYCCOIFWLLvVHTQM1INssAth6K9jY/ApbcOaKz8y7LuOc5kJVYy9Dwv0Bh6R/1F
uVJlwS2/pCToJMwPXs0eni9LasTJQFkwDIY/0S+x8QyZxQ9NUfL4Adf+34Mbz25f
W+PmEEh4OzEd1x/m6e8xZu0VsbuML4QIEIz0XhvgaOtmT1Xn1LFbH5Tlzb+hpnVL
u2ArIwAMjSIylQeFukfRNOzEvPhgt9Miej1efrMJcrKwrrZ5n90GQN2sIfj2gSpq
c8gJqb9+RMiH5N6AB8nbrr9uNcehJ3mLg17Xif5y7SUHf24G3DrddTgmRTSpMqpT
d/JvFcT9tCyMw8efvq9VvziH5k8PB8upEr9s3lGfYBbjjRZGmAVxnDzfRz2faI/O
INlfchmsaA0XZbkWSGq0n+pYbypPT3IUhGtDd7Y/Sl6fcPU3BPnyV/X44Eddmo5A
qX5HnuZLvFbBormzhnsXLpCfkrWtGiNnNeUfXhj6v3CTVXKfMgmJTCoBniezB+pD
EX3Yt5tIAFINhUBusma8CJ9u30BhB5h7fRyxaeOAN0lxgR0pId5AtLiVvCGFIA4K
MQ89FdXTcnTqUHzwFEbrS3Z0sUxeQtP730FF/Ff93vH7O+YEcAEKv7BtsgWRXy9b
K9/UKQYwY58eJ3oer3o2kGt6sfzxvxtOjittOgvrI7WWJJ6MbHyckB+5MIKV64jZ
2PrR85Qs1r46YO2uX9v1DJh4gMaJCsBZ+RdF7HPQy5+4kg15m5+XBzytALEhDo9u
ha+DmgmBvRwkfsFTds/FyCp1YOYo9EZY+61EcOtFfZfeU9zjUut2ETcq4avI8e80
vsVMaYwYGjRdGLjQuqolWAaVgxdJikAJNOdoZwsQdJfjaA2xm9z7vRXI3CzWOPi+
H92vYYAjU0jDGk7SDm/a22ocRdnTcZuxjJCYm9DkDfpimtwcT/2VLmGzPXe/nCBV
rSgezKfoIR8ujtR0XF4GivMEU+4BhpI2Cqq67zBxTJze8/NoY+2aCTSzcr6rvXY2
WASHBksH/Z7QEisX0HqBxO4KrWQN2PJGwjYPn3EkWr3oPFQBfk+1lUPSbkD9z5O1
qTFGDXHebYB/7oNx6oK3aLra5ckZUvR9JkZrwHuoO7LgthvvHKNCz+m7ftPup7wx
QoIXK6N5qcxbMEiUA1vIFBzFv4A6pvx67uzSbG40LpNOkjIjHXYuLd7EXaxUuYCi
HROv6EiAdXOKeUJ6S7U20oSRhNyo9zexdivSpzYExy+rKwTMGkvKK7Hjsg9jNW6N
ckPYTUpJEM8CLavl+FtMoYL1GTU86NHwXKhVpUDt5MKofYjSU8aI/IKjF0rr1PWH
Jw22rUNL8t56kRRXuSzO5ySxUdc+W0hONw6zJQOAJyGjXNSg05ziQVbya/KkmNT/
8uzaZnfmjyZlDGfwCaJeKJ54gTX2pE0EdKSrkVSYUzWmzjEooo/UVB9MsDQBjoj1
mMqLsdiWJsB4Zk2ufvdKfEr7Ncmf5nsXtGFsQPAnCR0x/p2wOlmsm115lCVh6e3Z
xQ+p68pRQt8Q22Id6lccLSvfv0AElR4t28utkQqsmQk/sfBWAJnv68K9CxYLh5hX
t5KCit2UBUpcf+/f5NIgeswlLxh2K2w3OJ0GPcX/c9hFH5klNB0nCuDEX37Nvn9C
kO2nv9vVDt2hf/GFPfOZo2tJFE4CaeEKjEkYsyeRg6Z41aQ000o+xRzFova7NDGY
qtFLVXQ1ms57oGwz/KRCnRh9ezVGfQiKBe4gFTgV3uqustp16E5HT78UczRSShMa
elRbQz6FCXhiuhIqXIzVeIPB6T1Ey7cQaRx5xQsQAIKBqGF47ML/4uaDRtAqszan
mcvsyistjsdJcWtFeysPu9+aYMyzQc2D67nyGu8cJwdZTVx38qC4945MZqJEz+Jt
64jg4qiP+UqyJMd0UiyhvEcYtbqT/OqpzPXU7RC+/o25wKURRwaTlHUPvuHV3afE
EhpwPRBCYx60RvQ62SumtGDDzqJUJkfD4mEp1DPSpol34ZGDViRoYkQhLL9WUdbe
iXg6e9RKm+VBgV5O22Pezg/XftT9UpBNx/0PfwaTi0UxILtFGHlIzcpnVEQ3M4BT
tbhbSw0blAgtu0w6Qv0P7z+zXZ2FIui1R56ygWKVAcIz89nwcSRX5j85gl203qtP
qcbCVN1BqfBVyK3RydProih/JJCqe88ZCP7vyNERTZwHw7vNvqmsJ7Wsnt7E+qhl
HLg0/6bq6Te52TDUmNqHzFKooC57x55rR3bQE7MXjL/PpqwjM33luTgkLm6t7QWR
7Oihpv0t/e4hSG4eJ9zFpTpHml/yQ0vnY4ttwsbSkZR9Z1cd+n2FYmXvH78WWoww
fYG5fTHbGyztzRm3Y8pb94lPckxMtsEsR8wNMX4hdVYzLmRsSYxMYxV6lMCgO5k4
X8EMDom2e2gEsMucxbiOP+efMKACz/NYSdRP0G7Kn/B96iX7FSgQ56P99dWmWcXD
wX9Wl1x5hkBrLNS49kmo5WpULt3p4uV7W1R2ZFe0uqbcTeNuEiofC86VXpVNR2iq
bbzjIn7XZkSH1S0+IR7CsJqPfU2OBP1eEvwqeYXdQdp+IRf/TL7HvcpVrwE4tyTV
xX6DgZLSXp5cgSGR4ODLrKGfqrkWBU8x5Zm1zky+rDULQsrNj5IEm3wh+OWws/lF
7p8FBol01o7Xyx1ljYUaA4kClG1r9w32PdAkdaWCgBvebJS65NR1VBMYYrUzdasB
DJlyNck1w3Ztw7/7nMARTVeDBV47zd6gTagCipBrwaO3XywLRpTafdrQRGsQDJHm
1iNri5PYEiL2i3jeulHbHT5nrhojVhaLVtOj6362ZBTD2ezIrv7jxP7WpBAk9xBG
FH1Ptr7lw2XST1eayI8ErdzGMkh4EvpkVfD3eYHjttQGUbwrBE0MQau9ITTWXzvW
AegKiZMJ1ewQdqIHz4muPm8Bcc2hHHtekVt99kQ0SMTEfPMFom+DGmz9MI8XQYEC
EcoMJasu6BTFGAqtbrT8gfpSh7TZsoblZoygdeqLOlJpdZWEGeerOFdy+5Xkj2FE
sSRQuT/9U+j/FqqAPaqUM+d4bxrE55+1aN9eJo5FIWEyx3TRxicHoN1q2qNCSkuc
0AcBTOmmYNhX499U6N+uCXoPhS7V8Sydqd+UBYC2enLlz5/XjI1Oe2FICaUrXDxi
5NiphDf6ExaJvTIKeX6PMT21F6DOJxYCek/1FgeFnvIIt3sgoASurv8U8wHq0B6i
41iKzlQEOnRZul+XIdaI+WuQqlv9hTMBrm0v0fcem5t5/gfs3yy6mMDLxH893wnw
CD2cdJRJw/MnoFs9sdfIjNnDL1CGUzuankRYqNQrXn6eWdLKcCL6EArRzFwuYSLI
lCGpUAQL9Mdwc+K+4I6p/6lcJMwMHxbI7rfvT7WcxxL33zN2+i1JZ271vRwAXroR
VY+ljPlP9d4Cwt1uygDFn0gS9DPdUw0uaSzpFnU7zm7F6ZDP7BPAy2mLMN+jSeNV
WYhR/ZUHu6J045+/lhjTQAuxVD9aJRkiJpOiPSfRycTWBNmp0NL9C4ATpwvlAvde
YMPThxHzdLzgg3uYa15BfgH292S/rLkXAFYz0olWPEXc+KW+eszcqxuTN/sYxAYU
gI2H0d4EYo7t1WUAR29YnWewSb4TGQm3vHZCDDvUCQkAbgTxMrADXqhFAYwYjlHo
cp6Thw3rZAHZ0eqqXdW3Vj8T9w1eVi7POpWUEm/+PpJjqd6w7u+N7FhUQVR69kj+
mkvNSIdU8g2ikhDKsV1irUeBPX5rptcgIHFOKky3kDFuWh5heSRbaEe/3BV3PEUX
UnXdxxFnTeUW10lMJXLL1+7uIRXqmioLCBJb2UQtmQDSgNPHSoYm6bm8mRYVeE6/
hue6cCGEINLKYuC6lc/wwTJmcvUlEhSIpmxp0Ag0vEvNEKpX9BtPwru6mPLjwbrZ
Rj8oZ0lDVhzadm4N5e5v0W4fgHtSCP0wVIXIC73wwh6nHKE2vXUan/hG8s8hfxxe
qmnsPaJEiosLgNLln0Sijl8s6tqdC909hgoxmf+j0WehEPdXVzgDfcF1SpNBLGYc
szUduwVnKo95MqICkohrTg6tyfboc7ykE+EbymODugYZt/ubV0PFEz3oWYsLzVmb
PzExnDMRVXcBUfLBBJY41gGA3kdlejGQyQZtGTtYIq64kItvIvNsmQKU+HKLzn61
HCEMRxLe1gcU4KKXJiVzg5Z1+QG4PZgS8HEqoWqKP57mo5MxAkTFHK01m8EjVC3B
9hl5rVc6BsmihjPP42v1Fjz3sA1yHBIU5j+QcfKB0ro3rHPJrvHOKxFV6IY8ybjR
nWXd3rPLeNbJK3dGb4JNqYa6yLTcl8tHEu8p7B2wPVonMASs7aKsKBChx6Tq3lAo
j8wb8jWDvy3+tC08zjrhnVCUtiYwFHbAgCQjnhmKCEM+GzLyv40jufMq5nbGmrcO
pDvSl3hpzbNE5rAJ6VysAlBpzlKNpt9CIxjWWP2Q4t8++yAkZ9m3kjetbFCWqhzD
SFXnItodg2ZgzDLMEYFq8ORQsA0Hkq8ZLfXn0nIIDcGZvz2/niqaQxBrKk4vcAgW
RGpAUdW+32bG6Cd769bI3tXej0QuJ/n7GtVT/L2/FmLk1c+rKiOhJIzlnUgxEFTV
bsCB/ay8uY1J+VEsroP1BfnRYqSyjvK7AbDSm1vbCzMfdOrx6GGi7cid5v81aCYh
Q69gEiwMZ69OLuR/4VHPPuvtqX+jZsQsVAx4TtY20AuB42IgpEgm9Yb1fvlgQitP
I1t+hJKfrtUGGniHuUNcavmaoQDrv/8VqRnnWKn/2A4ePBAgnXhFtN7Lc3KW1G4O
PS8Ru33G/c+Ea6DBdWiIGgA9FToQMkDmYUlrz4cGYg9CEy9L+xr7As6+tH2Drcx/
ouOhz4EOytsq09yYCw7zWMN+clplq4MwkGX/ADfBWl0GU63D3OT9U4FyljbKFqkp
utNmwRQlVnDiSdGYibjgABhSirKRUeYdolWJW2Q9lzNASQP9vAjvYZcTBdeF9D+0
9wvG5T6VFvPlVjVBNVwaXbpGBAeix972Qj3AqwcJV6rPnerFQDjmJu+HbJ0vNYUw
p5RADrRrtFEe0rXZTWf9r0mwB2WUxBWT4Fgp/nvZ6XkiRt9PiQt2QQ3F/Xv+zEW+
SqSpebdJaR8ZRKBGCyIDCM86saI37YeSTJDfvInleQDDqtwqGRWG+TAJEcmSGJeu
rf6g8KbHoWUQfyFbTrxHzWQuEz6uGiuEzgCBhtpmfT/+YvyhL7HX6UpxWYgegRhg
TBsoVomWhWJjzxvqN09hRteuVTQuzVEPPt9AJaFHpYwAn7TP3ZAwQ38y2j7FRhIX
4u0IajSPt7cxRuhm1mXzR5cCXvQ41jZKw+njFTmPNUdjScYX7j0fPqeEDjFnvJdt
C/i+oLW+7CFe5C1fKbBa3xmpyflphJ+LEzIuRqsF9khCzqQcXND1tqFxYKG/ifcC
oKNThF4k7fGuzu+B18yngZVaLy5Zx4AOVs/usQnz/FjRvi7c9YTn/P2zvTQBbs9F
KCB7VvsZvyLoXkBwAUhFXnkQuYMsiDfkKWmWP2HzBNbjI5xppffJpFESOy+D6sL9
meUKCdISW+2NjGuDJjcAmMfLVt1QpocJRunYBgtOVZzyjhHvgY9bFGT8eAa2bPRQ
2snQd118SkVuekVCHXQt5Qo4siWpnUqMZJ1D7iGa7bSY7mZQLQi8UPk2IqvnWCGm
tKyYcS0M1sXnvJcB6oR4btcsSOYIpDAqk1qE47oVRBiKZLfFYWznLUcybc/O6WvB
5mQGq+cDkFVf5PCxoqIrKQvWBNKbvi34fUYiEhZpTR0+S/Mj+OGvd3X8FR1t9l0n
1Rt815h5JDdu8JGXXqvIL5Fcl3UzFGTrvcG3spmO2gc875UrCNCnoewXe/MyQAEu
MeOts7hppBKR8w5y7afiV6J8HuH9G2CcgDXZ5Xs9yDgkiW/VL11CqtoB04mN7PG0
nTD8YB4MFlbnbdKUzNtmGzdCWldPqNCeL1OWclSF4Kq51uvH044WoAhtfJlJKAQo
SntHk6h83DUjWPwe7L5FfLAaJRKITLT24PSz9xWHTj1hQPHkmOJIjPP6E3/7d+qC
ibIwAdnMWyOYW0cJMAznSi/8eBX3ig7iuyEuCiBsh/8/Q9/vLkg9pfonW7LOsSJQ
A0Pf+lONBodbQiI0a1UVl/aBxNha7Z1fVenpt3meViFBC4ytq5ddA8SNdSiIzwVM
bDpdUKowupCu+mS3DZi7vU6i53B+/0r59xEEK3NGHWUHAnHoK+xmiOBmWl+/bHms
cIqC/NhBJSuKNJGrkeefBx/CtWkmvd2LB0addpuo6CE3y0zROvGlB1wltxA8mu8m
dDsgwVJeEwcFgYPiZ9LcBEub74muR70nGU00zEVB/JWfwlwLGlLhNKDaEiawilhW
deVXhbMMQT2RyWzg2eNzIWXLWRT7sb43mse8kJ1J0tbAZ0LtYMx+2agCsjtvjiYw
F5DwWrsUfJQ5Ve1q+XxKol7eLSJJ2WT5E9c/0oVJ1Ji3jWVuR2YAqgm2XA75GAoG
/MSHux9anpS4wtqDLceVAiCiH2tilqs9iinKEiS8wkOsq1NTEO/c4ugMbzjgTt6n
iMCgOBOCpeXGv4C2x9CYt9jMPqB6dmph8Um2mutPHOQlaoV35axweXrvSUNd+fIP
mZ/Q/bGAG/Mb/0ifW6DErIjAMtagyrXtMwRQaSbuaKx9DV11/3yjNO+QABBLmNEi
A6M4ihnlQAbvLb8yUe82Q8kg6y0dUzk7WN/PU2ALkscfbOFPapXjApV1xPH4pydk
3+GllSu9+Ov6k9t22TixuJSUaQimwSXfLb3wfdUwzc4t5vrec8t6lqdYqTxT2eWB
uy4GSetyltvphxKSmHSYGSkAGONSMY01FNH453ID4Y64ENqOGrV/7UHY4R4ChPgP
4MxvK7zv2aH+YDGYYLrPBuD21PmlyFvVvmkSNGb1a4jdlKxlSDF1y61GGZ05g+SK
KRwR7E6aqNgeCgqgUmHn+6L1dG6VXe+UO73MW4t66yPPyzYyUC2psjO4Dzns0wrq
HUy47lDZjf34KrNJ+vzbxjlZfVYI2MH36ZlYrj3eIIkbmxULaarGE01YNv3Fm7Nn
HoUg+i+vfB7EoD7iBe2Bd1jy2LaicJELoK8jerBAsr5Cf7L6V3Jpew+r23l8G8Ru
zDqSuIi+Sr40ybb3+LIHwLWOlJ0DLj/rbD579jZlOU62NTP9CQnfycJtAKRcYAKy
VhQT4zhWFNtJIfeM3k0PBsc+44r9wkJCaLsRGmXr0AoqNb5+a1Be/sO6puU78f4i
tMlOJd/sg5RBbd4nYBfiykedHD39gtFtK0TRzG6shPmbwrHhvvmTPZrFhIyo1712
YSwfj5XXrlXwhH7YfwDfInt9xnS+IaYdLl0hVrMnYB8HIktzfEVjuKh/P8lafsVz
FLtru+z27+1QYk6MJE0l+l7BNQ6z6UIlVyRnzNWolqTj9zKJf99aF20HxcYK1nJX
j57ODVCUm3w2APMHtZZJGPEUtMXob5Q2rnaeQHmDgoRrs7A9z7bQKUqGX1z9rdFx
CJZwhJcl6e03GrGjp7EkWLUHdKd5jhqlJbFpYQ+evMLM5TYImB61nYGPVYw6Y4Ue
ZV+JFWeR9cEj4QoJo8t2nrFH8kZuwO3tRSa/YKrS9E4UtIN3t3uNheLxpgTewejJ
v87MulGtX7dxTnpm+0lVsxhymL0tq0eswXQJsQbfw4g6CJ1Jt4g8kkWjWWql8v+a
oQg24mmik4DBGecj6JYtSi0Pb2n+LlmnikTbNRjRKfkvFdWqf4xivgmGAAk6ZZly
INfkPhJBU8X/G45VettRqxfyb7OodhBhg/sXRL9iSnen7owSvOqM4XdWH022rTrj
JG4R99xoZWNmE6pWZa79xR8f4+GbrjOVKzyz43vRupt6r7X94puek9qDpkrXoNrR
p9mbaIVvpXGi9/ia2QF+/mvI27AHq+h7w/lqLelISw8QnFqXlo+j+BVm5pvhQeZW
kpmriIudIF2BOKukrM60fsoKoFijGLc7P/p8GoSz9BlFflXU5W2qBEa/vxS4Cdlx
LdQ7weeu4WNk9CRrEXkNSBiOs38PRvG/nQn9eTPnvto1XTOg+SwirFXOGxWOJmhP
jh9wTIYrRMxpPlHllmmVMXW75X0o8bkUKKRZ35ppSGZt27G3O9viP7YCYDNLrKu5
mYPlN/ETYZE2j30MAD/9PYJm1wumA7mOH4lmytOCUoHrlTGVkeiYjOjWUQW24lEx
0b8b42tioxbgaHXtA/saG7ag6H0SgxrSin3W5ZA/FGwLxtJow2HcjRNwqevSPSkj
qJ4qtNlu6qktQA3b4Y9KlsnWtNHpfP2px9H8N2uwp0QK7hntKuvAeGVnuNX1JrSJ
wHPGKdKHNGsZPn0YeajTr6Y3bO6VEu1YHoBFXaQ6M/BX+vdio89PCo+tfTKOj4Fr
sitEtdTLhGJ3XDm3r5EWUOgmwciEdWWakgHXAONfARD85l+1HmqKcm8CntTO11CG
surF+JbhbhUWTPrcpPX2Cwu6osmlUB8d57Ad5mW1rDESCTRcxHvGJl0JkUyyPr5t
uvWnf0jhPN6bH6lsx9l4kgdAafDY30gFN1bOwCJNfntoIY6vveEWwM9ICviCqGZP
5z2/7a4SOgjCbqEWlKeH+Of6CGYdLyVnH5wo5wMBva6DsFGLPzUQTBj71igZwrNn
I7JsBnECLIoJsdoQ91OnIHXfbdXUDDoDWfDfm8J+cIzk/ahXN4EYOjH9cQxUkKty
7dHpr05Vu9expaGDSU6GGba64YTlxlYRjrUt+zGEhT85d41FDYxuGQklHmdQ4Dxj
6pD49XMEgus/TUMiI4LO2cshYXEo7IqvExvjYnENmU5Cxfv0UVti7mGbmTJF+cKN
aWLen1tX+vfLZa9pN0mCzdW1wv1dUN6/KAL5NpZr4Ubegw4MiVXflBj58iGERoYO
Z6ASN3gCRzJpeQrvr2dHBdN09KKZJftkonsMNJy4DorSxMLV8xXh6eZmWyZrnAkl
Aw19U/Jp1Dbiql050Kd5dI6+v+qQNR/7eMLe3PtddxZkglpRDrehyG7JaY0ueLAs
RnRkEXIg0KD0TZObAt64cuLBQGrw2FJzR66PZI+6iR8462nr7OVyMTwNv1ECIoYa
mKDvZ57PNhNIk+NGe6vvoFd2E53oU0HRmxh/hQS1SqmDtnxRkBehFnGZabZOsb/a
ApFX5FHOZ4AVIHaOKdnbfybgmF0LDncTEhJWc9eYTsNF7PTOqEaN82Ggs/3A28F6
O1nhWRShPdMO4ijQJ38MgeUNQ4h7o4JQ+IwgOLYDHdLnXssFaCMFpqpFangSfrn+
yonqv8uKwqZmfVax2vEjvCR3pzWT/yydkkRwqFWj3IQhPvMpPtUQwW2EJVqprU1N
FtZdd0vS4of8Z6kM48CPL7cnnrnO1m990gbWmtwTyUOUhWcCSKeu75/fPjYL49cd
Tfgh3FCBDGxjYKQ3dBrUKLYlyITg7d8uQu6beD25w3Lqaq2x2uL61+g3p2nkpuBg
LGKkJFktYiie0u9zcWTabSyHVbR+BpAcE92M6JTbvU7OQXzgJd6Qe5CJiq2Ogj3v
fSDPPTQxW0q4vU2l1pIyqfjEIGIr98Acw2SC2XIlxxFUM8hQCnDIED35drh91Oms
ERmBPWjdX9SyiwC4gpFTxk13S2M7Fd+ByMgHGbANeyNwOd12z4Bq0DGihziZdA53
FytxV8hYl8cnyVXqXZY/JedXuoM//e7T/Ug2PMmxQ1LDx1tz4110DRkB2X+Or+Tg
HSLzOAdxqEI7qovfQrT4fem0FYymwQtGnX438gfGkRmdDq5Q022yIpl+3/kwgK2b
oSxRp3++0BjqNJUMNqekXfghA7GtBFNd+nv2QS7dzaV1+MioFPemTKUuX5h/7kKX
4wjjazJh/7GlCbgUXVxdPAJVnpjdM5IYrNzdEPqk4v3osvdjiEgveMRYxSPYsto3
tVLqbfhLQeYr3HuwvPOyrcgzi7OKQjHtum40P68lZstd/iASp/z8KfvihJzIwbQG
thhFuwIgnSCWxxn8O+3ORsGQ1xzmVuvvmtexxKw6W9BT3CFQdnSOL7SiDAOxeK2Y
3rjmkqFZqBVJXlpcqXi7RrlfIoSFFtqjjWcD6EeJaA/mO+kwdJteljvhN8e4zXHh
x1X3c9QhqbpUkNs+fK3dfWHgXd9M20qw0Hc0jiyCmSx+YtQKTNphCCPXgw7DkNtt
J2UTl8RZt5wjxTuLLaCef23TXNhCeXGUP3GvyRuBp2ADAJh9ggycMiHXyKxq63zq
tpsrNPfQEdqyeQV6HcUza/eFmk2UQzjHh38RcKFkYtCPlCLBWFLGDL8ThYszT2T0
fjg/N3X1dm0KeNgXzk7stlrAqGvHVE7rp7Nb+LPUEYA8m8Dkwz/kaLR0ApgnqP/o
k40SESSfSxfVv5GtCRhw1pBI1w43gDJjfR3SINz6iM+kP8wiYIVDw0XBqiCbof+1
nQya4VSp3hW1epC4gMWsRqhTBWgSNP4StSBMZCQKeR+ZXmBXpJPogsJXZhaLQxLf
w7CwtIQEo+rQNgZNwxiq9EjJ88QU0OXJPcOMRRj1SDZ4kN7ou6KvkbiDNrEvkgzQ
V/BBbwO4tBcbJ2DffaN0RtV2b6p+5nTa2WO6Mwx6+I9QkneFniOpynosWKX3AhJI
qF0lDulK/WkhYVlwWRepcARpCpCvu8lWWCbdNbPQVJqsbuPTrkbd2D2eQoerBin6
hdBBZWA/1VKSXf2mKJS/T01ETatQBWAQA/7UXWzPcj2VVwoH0p7R1qczgifjWuDM
tzUBuwGF0kcY+flfMtbdWkpFgcjrh/tG3O8cIJSqnDDsacDg6m312Oa3kMFG3Dea
r/NR5XdkD1EaB4DEVEMCe6UCTZAzIVNPIUJ7ZO9tdPDIpdKLDqzLxIVZiBSyZyBx
mAtGcHJRrL1PBDOOKD0ih6AGMpzfSqLmu8L6wr5f9dt8j81e8LTeaVCxpaslYAuC
qdOjUC6JVwPv6rd3EPslX6V/IGhDswXkOC0edqgBzizx8ZU5tOhKPzasl4tR7Pd4
4WjndiIjwdQl3kgPlqv8zlXyqMMcHcRSdMVr5Ilj1CN1lv4pC8PSZH+3v03Q9ljS
8qGUcwLsuvARrnHGGodDJ+UrQnkatekkthwAJxPz2rmA+1XTlRLNTfiQW1aUkzpH
GZ+r2uhExr6I7wnUJOZ7n7OOnEdE1ukljTSy1IA9Ld2xC5ReCwWX3duFwiuYOhsZ
qvhAFAmS1q6fAokAn9AY2PK9QxeXt5azdgD3Hu5mZw1r3TAv7jdMQBDzrIsx9C19
LaJB5pPzDlF5HctOgRvF0psMkG12XPzriwj835qASmoYckPTgkDR46CRp86oWit6
xDB7FfAlEGQdk+mb/t2ruUCAvEBdNtTbDYICD5l6n+Uf+eBJLkiY574Uq+fkmXiy
WWh1WjJHGjDqCch2MqAw2TkBIphMGL/AV5tKIIPxJMMIdCYrlx9NndhP9oXaD9KY
4cnZMqLTc+FGuXxzZEz66Gmon0qK7QEmLTL8DqkOj+qV7enBKuGrEHtoOaJvo5cw
NzKP43HQMmRYiSlgGtKxT65Pn2Ex2OWiX2BB4zPo1g6zwH7nkzrm20IqYULygFgD
NmrHDOcch6m6HSEEtGgGDDaHAhOwfIxyEnEYYDNvmFYA9TW8nbrnP7TCPzyxUgKx
cguuBLryHao/VR10pg3cqAuj0FEvGsmMVCt+OPhlpdgOEc+Hnpx3g70hYkynQxWJ
0EGGBdiE7N9tQ3FS/IuABeTkLyyb0v5+dNgr1htz8/ZUNmHIawGjns4Ebp2AGPne
Q9jEOxvZxMbgkGlclP/orcihy0kLD3hygm5y5miymEZ4vxXvT4xpb6aVUmDkPri3
2GnByk8Ncm3rOHwo2AggcwMqVbSzMhpuLDmwHktXk5Jkks5/dsjVKaYj4cwmnTqT
5v7XVYJ238FOXb8lLlilHvk05UU+ExGxopBvirnNHnaju1bfnohxozD8TBug5It/
ujxFfnYaNd996PegVgmB6wT4W7F17o3s9uY6taf/Va5x/WNKWp+9R7SNxQ+4yebF
2SU21tZtzh0Qm8+N7UMjhHvtn4HDcUFYmdR3v1p869WzLldMJikY7+LvBUf7zzyo
XEMfnTqNQOVOkyfplYXbK+cUsYhuGYGsQvhpwvHTbSXHDYDE6TOvCISZRGi7pyH5
xEl2s9AoQ0E28YQD6TCIojMTIEc2qDpjTeZkQev7WxkFbmCQ6X9ALqeioeMnCtwS
lXKQKu/2XAffl46WwJfag/zXXVf52eHA2dAjbxKQDQLR4uyck3Smx/HbzEt2SK0u
yiUzirVoY7SmCEkEDGai/D1udTnB6O7189qICM4lKG1pMKSFId8MR+6Zos9b/OUA
XdQYCWqCeCMDzdPtblCh++hpdDA2OWh6KKOeqzo9VMC976YgTLyqPwnPDLYCZDzu
WKzh9thfWnoeCoIFBTH44IAhextOFI8bfTRja7MT8cl8JU4IrPGHaUOeSzQI0H62
XhsnS9d03LzPtXlSQ/c8WMh5mKiVeNQTt+CsGTeEi53F9zoP9JtF/o4fjCr4sDHG
tD1W/Z+nSRcK0Fhn26olAOHZgZoM5+i63pEogahPrb75yUwV2/YCxUwPyvsXV3Yy
L1SvISZCGYtE2PNYd3qN+zvd4RUzsyTvLqvQzLBmHSpZybPGBTOcxxfHlntTXBR9
1StNuMyzdqgjGeL1Vq5trKee/w6CwDl0rn7BZMOQ8DG/SdVeEW9OzF2HR8yS0oKd
cQYPY6lEJ87kltJEwZZ6P09vgsV9KyMTLHq4WLlE/UyGMxSaAbIfH888h2+/fJwV
Cl5KeVN3h6JyVwDCAP8frX/bGKGz4NbZ7WCEVZA15fcg+U4uzReeg0FG/VBYBWry
tGAIzB4R+A369G3bQejBpof3VdVVxFT0fGaa6g3Bj3yMKRprG6mIkUWNJsmfWL0c
g/9g1W8ikcVIazYoh6KDOlQbkaRjNKFWSv/t8CEaWnb28L87jHuICbvEZ2JmQ7NE
2bEMdFuhbrgn2XNHKKMdAM9DUJ8VzRRuRjTpiB7qByoLxrQccuEkRYgfZQNlW5gX
JeM9tY5k/P0WErh8TWbRBf7tnNGcoMiDaqI6IMQfWSAgiYds5lFatrlVw3cPdZpX
fFGOyuOV8GRTDSZOV4lcnSXPnd9WPztNi5JS/pqWXBybJXzacindoqmdl+rg2dpt
JdWmcM3duTLGcIIIQG1AUO4iTE26lgNT1KyfNfwIVtxxQwJrdfWdVhR3JfhQ3Mbi
jYEUv0Le/uDXHb9vFIOCyg/BfXhTe3TsFmuWlpJIU30n5nkGI0b5mh32Q19QH3iI
u3msV0sWCaQz+aydwxPr/4yssMYQl+TyLYvy+U+eg4zmiKMs8F1oM7q5sQV4ICmf
m63PmRK8vTS7DhoRml7KClC/iBfLso+MTRLEVf8GS8c86VXKLOSEXyOcxACX2ewh
ux1jRN+3fvQlatjl2nGEZ1EZCNz/yMYmtrO53zq7pUUB4mhYsbcPVT7kaouFiPbP
bXU4ipxHI54IprfpSymmi0RxhIMJa1EBqrDNd1pvT8bxLapJ1MD6Dst+wP46hUrM
+Fy0mzE/1xU30jfXycgdd5g3OETBm08mHCEXEfHd7xWL6MBjY44xE94IILlpz5z6
qvElk/AXhI1W3CV6iQ4W6ATr9TyqppzMOpuJmFM8n9Xo4n0kzLPHSxB4N9jLWM+J
SRwoBzoZU6Iqn6tN8euX0HK5ezNRjK6D1b4DrtcF4KbYZpHdYR7868W4fq5o5G3m
yW2MTTih0TU9sK2x1aYwUWUuznxoTmQmd39qY7qw7wAMVtOS8ekXHALD0M3AMyVY
izALi6vjJSitygRQ259fwFn7WZ5v7lDRlYATgGJN6sCKklvf57UHibd/wXBl3gmh
7nSSZ6kGXEN38HmE+ey4L1l9g3PZkY7O/sY7Z4x0/UvoWpFN6HAbHzQJAsxrrOV1
d1m/OUl21LTnQ2GnTQy12DXd9TlD4Eys2ro6R1Y511DEZzPVUJVLS3LWSJQNCVjX
++r4JF7r+PnP8HtJa4Y1J3YJ2wrco/z+Z9XBM90DAZsR7tKmvgnUHYek55M+Tzwn
wSzb/QhLIipX04j+XlzKNbeNVFSBxBMlNe4lyE/bEXP+Q8FmyJjbehGtBcIT2bYb
1WzUngfKoz4iHjqT+uSeIE9c1gRSK7gDKQZvh4q1w6pQJNyYIdCttw9dJFGV3sbN
nT8HZakKh3+nLt2Az7KVVi79gHDbygCJbRLsf4GNmVwsR3c1Hu6aKEx/V8y+6zbt
BgnZgzXCADwNFD31bqPwtDtbRQYZxpKWxWdYWkp+LyxnzfalKCU0J6j7MyJ+FanQ
c53soDdDGqgpqleEHPbmxW/GA2az1DkzSoYMefYtHR7MR5SyTdDwPANyQVtCtPQe
xtBL7QkpRLFUUp16RA73TQx/miHCSV0Zip/tpqfjYopdx4KScEwh25Prqs/GHvyr
fUyBYJTCstEBccEaC0jr87pnH09GXY+zuxGroitNC0rBCUHV3NhrH2vCwFQwx2SG
OeW1ojMsb3jQ57oh94EOsfLskDqFr4rbIi5UbHpDa2w7cd/Jfc+5Es7Koj5APMHt
0rZeKcQtAebcH4QZlSdkh51ycO0NoGnf8hBxkuoZ/i4QkPUcADzKa0d7CG4X2lpv
BMZK1L5cSmnr57wotiiOpHqrJqOe0U239JtFuMSBAYpT5gfGw3VvvkVEdlTgDV+u
tb0ZVgPpI4XhoK6wTX/rlicGOVJOL49Qe0WrP1TS8aJKnXiBaAqNoQLdqg+18WIX
2TcG7TW7TG17IAQHx6jZXhtr+VeJBNpS5fL9hhk2C2Q0S26N5AvuMML27pHnvOEh
n/BD2VeJF/rkA1do9ObTCg2kgtc/JpMX3/ZsS8DeZahhhIinUiKkgzLvCT503xuk
95uarZNBjNXsWUnKo/YMp4oAazRcaSuruGv5U84D+i4N1W6Y/ZVvLuKo9LF62tI5
OHmYzJNjot/m9FPorRICCgFmGS7f/Y00BT2isOD5EZ3jkweOWwpVKR7oue90QinJ
JiHK9X2IlCBVwYCPrRdIZXQSxJvh4v27koFcul2QR3b5dREyUWlykJeg29OCQIsD
nJZ+3tA8xxlezlflZzQOnvxlsFQRz8CAjxFpwA2ST7MfXNQtf8EaHpsrHw46uGqX
wS1ulZGcxMzYZ9RYMLyjb4K5ROxwUQ9OqQHZi975UPf0j9VqF4SfhKZyNc9TSyhJ
FP6yflpd+18/enCVNfnIHPMv3OJt5Pib804swX8ULv2IHaavQ44oD1qs8su+3JBi
KWI5gadHsFRmLxQYKVeYaXbpBpHS4f2ympUZ+j3mR25Z0Obidd6aMiCCxTLY7gWU
VodnQ1ZIK66XERnOb0J+v+MYDk/5svjvfnwdZNYJAM6s3ei0kfYw6BI2tGUaClBG
2ob54iIB62RyiCbthWN5tnr45P9Gcco9ZhHbx8r8uAoSPngiN4bisLc3vo/WXCKh
dH7b9rXe/SI3uxVs5iFuqeAAUJPq841ByVfy/o6OLPkOSUI6nuQ3cLRkxkoOO/S3
Qoctr8J7n79aK+OVvIuAB4e9wwJqraT4ivCLSFdjNgN3AjWfRedStuhIalfA3O3Q
FULjr+dFcW+iJvLJmEgynr3pJjdOHRuSzs2f4HlsOSZ+SjCma+bZopBfI7TpFksf
bX63Z6huY9yr/SzfKOov82kHZRGb2ACRRq8YS662LOAbGq6opv4uIuRccbF2uVw+
+Nt3c5n9pL2jutI9sMfztJvZ+d+lEFYfZRq6MK6syaZfWEdjn8TgQ59IZMlxY7lo
B4bIQB9SkcaPmjN5RHmOSOdFCZMYBygy+3DEhpgBRp9GQQYW+xGbegIKN4floPtW
ixMMzmQOhFqM2ipe4Vm4k3DiJX4jtGXC9Wlra3L84BQ+3KGK2mJyJOauUZJSNxgX
2+h9OU52oTUQuYPaURO/C12SP4Wag93F7SgElNkQ7gGcHCMVsLYIlaSwDe/GMqvU
gHXpz4Aa33T3aL8vB1Y++ZO6N5UHeX9KW/u1nDEaoCCrcaXobKylTaY/yilkqFDN
OEqML4Kt96nclrr9ZssqvgYJYWvrpwSBQFt5ZyYI8ogcJcaWTyOzd03bCcxGKJGn
O4xtdrmvo555vHAk4NRuDAcQOnsNmqtmzHvU44fmWfZqopjhWgzcxyf17lBZSzI8
LsEsEkrsGy5cVjPKO7opa2Js2x4J8sIOYb0ircYA9oKbnm3f8oOSC3jc/sA7lcag
UNp7VLFDiNGaQh93CsXLKamdIKosyi75HWimxk0SmVdrDvIV5Zpi0wDzsKINPAF7
K+icPwfllvl8DYm6e6YtcqWnU/b1NQUInl2KOXjkfAUeHqUvH4UcWHlKJEdY3W5t
8zmNugpKD4XO1eAYLx75rftTjeltCEmn9U11cxrFadH1PrhwwsnYz9gTnefwXNU0
T3F7ogzkneS5onQiGQSpm/vI5C2P/GXh2hni2cPVlJonkhUidu4/MxprKizoDlpi
07BsDm8RWs429fJQz4Q2dBNIgCR3+21U9PkmoM7vMCf7dZ+HDXo7evWlDf5P9UOu
6k5aWsx0zWh2bJesWtJ3uG6YLlvL+NtN+QxrpVsow39kvzu2BKjolX3u1idPNMYP
dsQuLzHU1mJaxNRZkUKmXwFoto2ipjOIw2JBmIURC2Pfrd3tLi+VrZMmgBsEPg3J
X7V/lFVg7jidXxhxSVjYtuTiXMSZWJmI1LXGo9v2S/90F0NqAhGdBIA6CbQ2aqIL
kFhkUF27WeN6beKo7LDdrrkAkp5d96R9kahHCbIlGFLXuvH5gMK7rx9vLXZ0hMRJ
9hS26J1ztu+RYySfpM5GowvJaWl4YactwDAE/9O/Shi+weOFuw6sGzo5ZMN7gek/
Yzm4+Ta121kVTMR1UblgnU+sHVbia/aRDzKvNmcic3Bk4r7dUL6lgz2ltf5HTZbZ
IbcmDFzfpx7VxIMlM7/iJRiGewTAxQmUUnNWqJofSIw7yoRqWmDOebN7QTAAmqi1
6ZRGh9L6LRb/zaLa7XZuR3n0Vwiu+y0fmSGn6ta8zAL3rMOPEtIOCHZWjkbFhrQU
FVdcltMfaswQ5luDvmJtVKS4SCmVT004RU1HNoVvf6PhNruxAgR9egIlaN5T/yZy
q9OfCOOc6DCda+JAHNb1LvrhVMS9F0pi8wkO/TTUrQ26KlaVS2W629gFb8fKe85v
CHOb21Y1VUT05DFlwCQqKy9qWWd9bnlQBTcbvkL7OtcauabrZsJEH7M7WSXnJFaL
OT6mNCA9wzkm2CBe42ae/BLRJIfw1mQIhu43FTId1ayxNJbJXKa2dGQ2UvD+zcaE
J5xoXycmQLKtDlvosj0Upu//gJ0WeN8wKwFHCurOTBFJxY8g/XyrZUhO3jiObYYL
8L52FKd00g+bl/i8TaDpbWXz9vngxc8MoM9m6DBnjzzYr4kliVRvD7cWpeM0VHBl
aay4hy2VoH+hGVc5LqrBtFNI/i8wyUsBrDBIHvhGPDoL90io5S7mc9XwYqKtElPP
vSNqKNGqFUPV7se+SinGdRc5pRywZQsSudzV9ABl10KNCv6XSBNRu221tCXu2TQ1
p72tGQeDJYR43jWbQMaaE5LrOY1GCFOa+HK+1NYr69u7kHiQzjYBnKPvB8OYUb7y
UZht+GK4kf5SaaS6ZApkvJyPAMe/yBz/0TG+kLrizs6xWZqGbGQxIOZM18HyLpdW
WP35y8OxU9Vo7L4oD+xBDIh65jkQu784IB/oJRlRR0ptiVBR9Kzi9KWMUcxtSjMm
zpObkRYBNB7t8iMiOdx/0XhnxRqabU7MWl2COWKFhr0XU9KNNQU45rVkrWR7AICD
TwDakuBSRkVqV/xhjWNpwP7GkLDqJzVDD5YF+hOBhxOHCH2O0IB7EZGw73VfbR0A
sL9WYAubiXDA6G/tKkcvNu1TNy098hHNv0VJdjWDBy9l3LtXXel+6xdKbO+r/ILI
3JtTCLgKqHxiSNEuW/eHeh4AQAO4zUDkkVhjTL12Ps/mwyE4Gu7yzHK20Ecl2w2j
EbaHvWwr1WiN1AfxkjznNKh1/XWeAvExxLzjIgpX0N4AdY7wWeSUhLSypwvDmFrn
U3TvX8BApnhIGZ2zju+gxK9OF8omY/h0UVSpASYa7DYXkXDL+Vdgi4U4y2H7zfS2
ym1StWKh2HC6YZqoQtI/h+gFD+skxE2qjZUhuh52waglhkt8Qsx6TGfs/QLJAgps
+QQOp8vK0Y44zU3aNSL2Jge70qzGhaKv4PHFI2QNrM21rPNrL3aNt0+72HxOJplY
dKd9H8M9qLGfNMGs8HD6GJariM9LpIRz0XTlz09Fgg0eLbwuBl5zy5ms5CzSDmCj
i/Y7vcoeO6QTMOm6VaNlfW/+8IKBkAWAuYHrA6ZTd4/27JAgi3JQmZxQa0hbMfXW
8QolaESF6/Sjs/L+sKZXZcOOOnS4o1LnUJYGilt0aPxVcxggg8U22m7taJm5RkwW
xySLEuyoQv1EFgo12tanAeX4a4bGy2+YrJKLH4GbbJMsLFZ3u3vjKaxfSGiefoh1
vVWzA7Dqat/vSsvONM9ko0MEogQJQlzXu0VJjhPwVh2D7+Ofbqn4Jpye7ACUgSTq
mogN+NuwuTCDwXhxm3DmqMxQI0ZwLOP81cspl6MRWJIrJc735D6+iNfgTPwbe12g
Ymcvw5BlYc8ot62hD2GzQTkolEvtCKSt7MIujyRnmvV2a/+51phrI5YGVfPEUx8t
a+gwuEruj4P/GC5ARgXpUv67vmqtthyOTTv/0leDdwqagTah2hvOWetiOZBymV5y
cY4yJfNQO9G6vz8w2oMRHCU2ADOrE8zyXq1Sqfl1ikOGiVf1AMaWLRIGfwsgYIQ9
xYRlK4wqXnOffbww+FdTVB+z3tKXih+YtAeTfbteWISrNYPoERVvMIZ5oClAm7AS
Xlv4PrdZ6cRI73PxFh5RoKDF+GwzW7bsWJonFf6I0q7E90XgTHofZwZW+ZTma4A4
nvCJaqYXbkHLQ1wUQ8PisNWo8pWozw2G+Hdovrs1TmLn9PCM/QwG5teLXki+y1y0
0sO3ZJYgsVId3rAVG0iKYEOppckikVUVoRNch64caye42IzyPaT3+bbwqa/jW9YD
CCqnvfsXbKynZYW8do67FgXFFFow5i72HifIok2TScCzTdeKxfT4v6y2pl1QaDlP
xhcbg2DaLfBoIhRtL1E5Ew+Sua3PfN+kyIKB/tSgNzOzor7hyY35nptiwKdizeDf
YSzNG7NFN+93DjUVvzQHINuVo5cYDaE9S7zB1oZI4sehRyLf+MpsD9LsCHZ5rw+l
pnHqV3Cjes6jIrIyyG1ZyRPujiMtyXohMb3u8gL0UvEMR/X07TJ0tYWWOPMKKljH
q14ao6Gq0JhYqpiaxr868TuqRCgzJCAIxpoocaWnIPLtpshfYlLTpk7GXQc9X1aB
fgMMxELEwqbL+Qg9VYHDBqOQei2ZGdmL5bV3jPsPTpMsXKF+3yV+vfFhGEUI1Xr+
Z2eDJnnxB7myz+5D7EBqY4hC746+R81almvvsa2RF11FZ4CDV/RaJDtI+hf+YG7h
QIvrHhrkdizTipw715aq6zhBF6OjXsSRqSvz8m60osGAZajFGEMyIkcQs2e60mbl
ffQSRxOYZLe5ObFOEgg35C/MRZvlSEUnmgftOl7e00Le341ppcJuQ9hsbgDr2JaP
OgofL8OMvZiBQhtHQnh8vpwt+h5Yk3UH2C3wXaCEZ/CG7N5+6P3nvg3tKn3KjuQE
sev9h/kIaKneISOmy26yIrfOZpLg+TbcS4XugKSeXg+RVqtQsislJ8BlKAhXS4lF
L4qhkO53X1ycPy80fcddsbU25cVvVT12+5TvPqsH5FzgIPH6RlitiKaTQk3NrfS3
wJN+xo6UtSwxK4Jbti64AsnVxcuMDT9pHAWXFF9kWjkAya1RdliHB7CFhvQHiA4N
KdOTOtIxVKnbx/qXZ5NDgYEzsDdTnmcC06W07W9GNBjyP/v2z0vx9o74NLzVNGzK
1RM2vPLiyceQql8ABJ636et/CTuH18HNQzf7ZBcaQ5LBpNah5n9ebexiD8m6dD85
bhL7IojkFBI6Uc5cWeoTVahBMh1oorlGQpZa6gJvCe0E3CK2HKQK2fCPsZOEjLgy
fbZwA1MTGaBXLZ+AIZplEksDL43jbvBdhEkb22uaH6X9QG/R/BtB4MPtd5NT9+Fh
wSj0Mc/OOstOKds8mlBRAJrPCg8ghT8wapKJ9FJ2EL0BY4ZYnxzvhUk/ff7Nbwvs
YRxiKUfV2Ci/+33va0rf8ggarB55/7lqMcVLmoDwFBSWdRcPfPJdvqyrQifRxGRH
ZyZPVROxXBJWSRwvq5P3T3y7djMPi4w+0mzn9DDFTLB6qBCP6AR76E/P18NkGXNQ
Ih2FE6HNmpoJEUbKnCpe9wHdvRM9rWEbxs9saU5vxg05Vle4Fy1cwZPg52h/XyJW
tDgesADKXWHaXwla58AzeoXNElAJn5iO2mf0QaUjHMpYs9UJaOOwqQ+3OmIwDUN5
6En/1fI/h25Xxgd8RZKjLFAxS1j8fh7G3fBzY18jHiK2aAmXHSqpsER8f/y5MRbe
DX1BQUG+P3c0QO5zsKqxOBLGBlXlLVAIQBumbvLGVOgM16eUeLWxUYQ5tKmmvYrp
6d/lhQMCmneMqSuu8/qDKIpBBftL88c/Eqy+zHegrJGVp8sd03mAEZDENzxVJ2Go
Qvq8AfxflAcLZ+3PDVSfDMCcezp7PMlkC3K0mHgLFKU/aDutYeyS/BTDujhjeO3a
66HR4PO63Ujars6djg+AUuMyHXZSBxGtmkOHcy2i//GRP5lJfp2aIcfqmM2+EUt5
Y9PM9KQttVcWL2fS2E/miBVaGkyUP0Jcuv1hW6p1l+zjtq/cq0m0DcZ4/cUh3/zm
5iPRtfwiphCKHWBApxLCu2KHPry0k7641Jh0bEKDfZZK9dFLTcFXe4860CRj/qxq
VYmb2vYAYAm7xcPGDbWyQtdINXP4z3hYiypTKjC/kggw+2gCkgWxrAJU2vk43cCI
+IZnH+phfS02QTSo5vER4xmzaMUg6kFcPTK0Cvi/pg2uvGmR1CoUSZB4W/zn8ba4
eJqG3+cacVAU9gmPI2jTeY6jr5cGvpazmjlj8E8pPOK49l0tOA/G/pTz+YXOPXuq
4uS/NhuZVL17I0sl0HtBZiq8cZmIxbGQaBX8TDuLhipidoV7yz0t/xFSmDirxai7
gTxTUX9khP8s+PWiSLkZNjKhGTr2GH/EM4+Af1o6ngf1buHXQI8HbmJ09/jyhqJ2
8k5X87tLOifjt2BEtN67rARNl3ZuWoX2329s/+JTjjNq19/n+CTEMh+Zt4xrfr5E
k3BHVHbxkyr7M9Eaog0HeoZsaaJ8FJAcgom03mgPg3vgcO8j4GxDCcwHZm5eyck6
rJW0cBSdQJXYRKgNVqlkjgJUN7ivND5tKfyQoIZkCbbDCyblMQ5pPS+g0XCC0Tdt
q9VLIHKLCigrE1WXxguGel889yPUu/YflihX5Oyeg5ByIaIKTOK87XGKtBa7RBrr
Rl2pn9IvODpvLKrJx5k/SLN0j962IPGYFH82IpiOADSf2RE2Y1LKEIS0KAFLZ4ND
N7xVR4XaKdGGSA8ARfRQGPg1FA61PnZUIRV7YZ3svbqAlIRNleEyCA4DTWVHuReW
DI4aIYvxra0oCkR17WqVXjIb7p4gi5xmnz28opcE5KZykKXZNQapW9jtQA1wR/4c
KHRYFow3c0gaS+ZmY1kJluspwRXnLUZu1vc7HJFHFucRf3KVvvOE/KXSQq4S3MfK
PZ7yTWUcitP6ff7R/AUSv5wzwlxdm4tu8qPF8V0R6g5eRnESnYe5a8fmzOwxf10p
+XimdCNylsmvdZh8/ZuHRIAcVo+8+kBPSkC3vEiHr0lO72yFoR9Tt+oKhBfuScYo
Gkj59hb4ObYB+L+Bm+JYqwPRBgnkLIFPyclC4jHE/5MNjmSnrTWVm6bj9QLH4xUi
z9E8yZ7dUUq5ke2ow0HICGmi7RKcazH4RfnqmnLXBD3KwC2Yof4tthpUamgnoYXt
ZIqTTFcZ8wxrbFpKtTOcnn1wWzbiuNqz9uBZETIWlt+ftDgfaGEzOc5Bf6MFoplk
kdaEV+G9bYEQ+fe5/ApGgzpRlBmKMzcu33Ztmj8+pA3GSOlpJeS4P5KygiDapCBk
kfwHn4uLLmNVOiQTWuk/3LdfdkZFHWGpj/PFKAp3bp6gfxPDksZHHGSOh3635Bbj
FFqFTu1E5+wrQdI1ymFRsM+A5xTarM2NC9lWdVfryFxTe6JjM+17uwBEoIbeWreq
vfs/xqfGkjWySe17aoNz3PCdDZStrlCqnUs37tyKqe9eh/gN/X1HVZ2eeBWfJF+x
8jCgaRplSnjzoIlNZKJwXRUXXSviMCY7i09SRlwj4IGOP0p1kM28vrdWNA62iXTK
m3UJN+ef//hebBQtlmYBe2vZjKWm9Tng45cmlijAnOs5OKf7n9Roe2kpprU0NCJr
0HIuTxvGZsqeFMni/ovHaTyn+R5k54VGnwVxjNgqPHORfLGXofZURdrv8pnm7ikI
X+PJou5Qg04lXjOkwO18e5woXJ/3U8YmVP2NiN5dFP2TfRbju2rPlLe0/U2x/O7n
72LWRKGFDaYv+ayrzKgbSb1Zo8ZccKQUpoxW6VIhh123So8iU7sVBdCn88P+Or6R
QGxixxd2uJFqpqHtnPwlpxeXq9ZHCdet/IHVeBCTODHvMD/sNR2YdxPde5A2A9HK
jAW9IhYVpsucI8pfRSXAOBIA42CyTEql8x1ovuJTuS73J6fekmCzDTx3fycMUCh5
Jrcv4y4PGGEaPQgCSqq7r6r3MbVNVCxbodXMuWZSAjgasmaCeGQQ/UYRlzqhp1R+
QUxYosM184Qu0ZimxIdLYRDbrC5Y6xzC8lvCrf9rThJRYQNDVfC9BaI3KQciV6cY
AfRBxWRiBlyyCM73oBBvDF2SCXnSKcA22ad2BF8cs3/R04WWB93u0qRu6qpdPHzz
EuouftOTtha+z9ASWL3rTZdnmeCiQKKLasiIBfzumtIcSXeAcKsXwDjk6rw9z7Rz
5Q0HBU+UKDJDeRN00UEaC6sEAE1ZGx/SAt6W/i2nSggjv3cpYUZBS31j3uIMmr36
+bPtsQzVp5GaGjBd3dH7J/KSGK/uswUAFXhTPET6gwFwlhDhLBerzOpni4QdL6CU
ZWzS9AD4wpiHMor3EWymdS59usIxanuGeKLtoG2iX8A097+fbxpCSzfTdOdRKXys
cTQyC0U8jkeyDAPfJrAncvVmh2irtIYs7d8Rr5ocsXRMuRtKOqEonUjLGw0gInPG
ZiLnzjP+9YIcyueFSPVkM9Ju2IyTepE1dVajQAjk7T0XqKOoOSvcKyfvgy5ZkR7K
C+vXRWbIs2SxAO0nHpWdIAjipFIfId8VHZmdMid4cAKpevhoWJkO2lR6wBydacfp
pwNLltEy2LjEZCvq5AQ4L7hBbcXTKA8GSknsCxo0T12QF65La7xhsOYwaOXN/57y
hRPW2dnuGANZUhoaxHmSbQ4FKlNOduYnz2Hf3pDtUVpleJchWsBmrUh+oSBQZumI
Q7yAtOuqJpgHiEoqG4cEgefndoFF+W+oFQgyPtdRJtxiLDhZ/cH6EzDUkMgV0szF
MPiFFMSOCcxMiYiJbQRkFWoF6ptetds1SUcFnBhv9BFNNzHLAs5lah/UHiXx6mqJ
GQplahzqxIZCEpGGMukGZ+2GAJJiYpVzm+V/0kvYi6wt8izS7PzpVhz+hP1l8Vz7
JqzwAGqCYP78hFGzCAq8sGY/WveuP6d2wpoh3rPaMBJ/5B9PeQx8k7MwNd3QFyRa
zN17lOlVjFqW6Za2djDng00R1ZzheR/U7tB9iHinDALj7anvU/4EwPW49btXHhkE
EMfrd3RcvuAR3vkrhPOUjfL8+sMRbXmwAi1NQNrX9OyvHwPsnIlY+hzdygs/3NKe
v3TrFvA4VOvjmV25l1iohlH9d+cCvA7hVkk99x3kr330C2HYSymvpUCBz7GN+oca
9PYV4vdGm8S8SxpWKuMcw18ejptCcu8a/lGWRce5nOJkd8qdzxNlnoZU3IUXUb05
qbBqY/mDy+j569pBUvOnnU4qdzvEzcc67lP/V3swG06iPjXsWD/s3RNqIulE64KY
bPny3uvlLGmu+zx/T3ISX9ox1O4GhzCov+yw7fK8UCvX/fOf5IqhXmNdZYzIhQ6i
8TxCd753Hx3KcJ3iqw6SXsSEVcU37ZR38d3RaB/cd6E9pWBjp7zPEthVSceX3kSo
V+K1oRK3hKRcLruazdm26P86dyRPRsiwXtNHY4xr9emOFO+5IAUxAw4cqC6/eEes
aveZ+HKiHHpOxVtpgEPEgUH5BBIMq7vhbnSctiQVG/pz11hYjypeu4eYb6id4p5f
9TG8p+LyMWudcszHdlhtonOqWhv9nfxfpYSUVmxxIrXl8cgLWjvpIMH4KRClHVkR
h+suPVArhK/686vLwkcDebUy5luAASE88UJNg3DZrtxdPy43iQJCZTRyCsmNqs80
TbU4bHfwjd5hYMV88kKsnjj4+CZ2eUj3nmbOhLSVMuxBALmZQ5AsBpmklNg06r8k
MI+TyDU9wLqId5L8P8RznzNGjht7ZG+Lggh7fccu4XCKTHxpJ+DWOQWn8RjHZ8EL
o1lLOjREbDopjkgwSUalyz7pft9b/K6TzxpQrfk6BmyArqH/NWa3gL73bLolVMZ6
mOKhgbbBt4QIGAB/kjH24MVWV4VBu0EDFCwsgfaTfrBL3IyyA6A23omjmZZGI+b3
9zlaLfipINaUNryJ+YQhIBaSt2J+rWp33765DVpL0OcL3raydrxXOP5ZwT2t5LE0
v5AgYyhp2VYWtsbPKaC+J36mO8kPfEY9I8s+GcfwYLbXAgmD/PDmEAf2O6H+N4Q8
/nhPTT3IP6VS9KXPx53KGkIVGxdbpSN6JBiOZ3QYVJ1yChG0ELCFZqNHX0jy2Vu5
17ZJCJDGN70sR0Xi/X0wXRf2/LtKew88oFYFrhd0jVFvp9pIlVP/cS9wowf9DWy+
a382S7CzX/LqzL8UeHI2lXxypGMO/OrJle0MBneZYGY6o7OA92JDCvLzq2i1rb5y
UXOO04Vv7Ev0W78vh85qx+Jd8E+ub5JodoP07RMftQQFSDJIhTdYLKl3g7w2JZQo
SWgHvFiF7d5aMQwnwe5RnJrhsDABChXAXvvq7t6viZFcOO8jj1vYMqggkp2UVbNg
tOAOgPof0vJpf15p8jIFl7TY3Zq3/NEhlOyix3UMBZcjm0l3VGT/I0pLTgMawop9
8y0uJv+rw33Wsx9bffJuFFDXWSYjHksPGFQ8wfxXiBps2tYskqsPLP2uXG6KMCE6
vs+zfHlDbEBQw4UZCGDq1WIzGf68jZXzbTqapZb4y5kB2Y+6MNp9ZEWFcIZbq7PW
IeeaoS4OkAEtjZbHvU6HTQ303NolLPNsHJW3pPMWzBFU+RSbGfKvzvaIMMNPTNlj
if7EFNbrRFwfjCX1pNAh3RIsmg5MP18lLNBLl06f00fLeRYSSNhzjAsEnL6r5pqb
1NlKGE/h6Of9gjZHU37mqJR0dLwIWhn9O4v22qKCeByvT0MRU7PEL84e2HFFNHRm
P7KLdziONR0mFfIm49D7/Vb1e794ICGE+O241vaXhiuCDvXpYXSj5i9dcLFi2tkl
W1nrAcypFo2/k7Kv8fktWErWMbYUOxoRRDpD70KumaGtPnMNu6+C4KdmlCauJ/vm
t8E9OC+joxzjpQZTOMvJMwNb5Vcc+DfvOwZHF/CVNN8nDfFmi7Xe70n8Ak915vdP
BjkrcAcfLrBTa4UwXRA8sPBRZc01trsQNxG+1OoPfZuxNSyI8hQ7JXQsVkBAscKd
uTjqtVdvL96bqbXt7HcTab8gbZX+tRb/8c+2axdnMlqb+gv2HjFCNHUjCbpT7tFq
93jG7igHP0/UZSnNyj0UL/59EJDZU/8aCLzDCIyr2jaoyRv0w2vMIimqPLQvA3jq
3+zH+gBnMsKXe/QtyDeCvBWHmTIZ70+VAcyNUAnpZAb6yEDiFsAWVofhU+vbifKT
PjWleXvu1L2DmcPfL49wcJvA3+MLgiqB9qAvbEjf3Oa4czviyw0jClDi59WGGwj4
/JKyt1I+MytpOxQbXKYu9wYh2S54Ppuf7fkW4dJyMX5OURhEJci0nsUEvhq+r1Mj
LA4zckug1WuIMYC7/N1B8JkIFy5DYwW+oxpvwkg/eOGVs5MY59sCTsMlBw1rDPf/
lSmK7q4fzXGVhaV4aQN0qnnWGeqERMbeJ1xPwyNMtvo6et9fJp1q9xDKn4IzC+Gs
Gn/roubXV0OkaO9oBhWSqhsT5P6G0JYFfuCulxtGkFeN5yl/8vag4IrvAOnsxLxg
JLc7nQCz+d9+wohJuJhoubhP7vb6BatDN5X1YlZhjdKOFfXOSPWRSs6/q9mmqIAS
88IGLzL2m6EmeucF0Mv3/wZp2VJF3AtzTKb2JD42hXcUW5+pdQONRQ33zQylwTX9
ci/ysYd40MLow0fZgqvtHrFd1hSdp0s3b3xdIqcRBHtPFHZdVBTb4sBp6PG78hEY
oVqayqfFHT8p9pv1eRiR64EoDo7Zgnr+/IL+jUtKYKJS4O2wzlrSMiyDfAqssVZL
fa56VxkuHERKi8BWGiivu/a+CXx7XbmWOXQzQsxx/7aF/zjRBSggTfBRv5YJEL45
XEqC9EN1IoV2xb38ypwy8esUB0+aHtzuSJRKZ9I25oQSmpNujREVsoUY2lVhCuT7
8WR6c3BOLKSDX9Nu/NSr2yOWK/5hZ3sk9AgaeDAZmnK/TztAn6LGx7/L5yAs6z/h
qjLXqSYkR4BDmnx1vbebjqV7W17JVkhEXfwJDHsOjrffs3Wn+dAJn4IZ9AXe/noY
bzow0sWD3w/3jobhYSe76uIqamSWQiP02VXxSUH3VFIxO8MfC/PCYbKM7aaL0tYC
5C+HQyk3jsLa9juKJrO+a2UJW4FvbmnSFqyxCsG1kt7CrbmbYneJAkqOnHMNTh+Z
+Y0elnBr04kGK/6J2QB66SVpMPXUT9Pva6U7470w11wWkoejCjAbEYCLZDdKsEgz
1V0LH2JxhXFJf12/p5wZMTs6+MK6CbaHJ6IUJm1DIK22/9/cZuZyPnJvhM2UNKbS
aRwMrqplyDK/klq4c6iO4Cr7FPe/32JWVTefo0Dr2iv0i7FPQQ2loLAJBiJJoTos
AJ1plOdXYG6ajDmmjKY6aU+WPt/GHUdJJvQ8utpbxYxeqn7qVZ9/Ih7RlzrVOJFd
XAbDcuvSTAM2vdV9B1sj2h0HY91EkOf3ZeKpNlj/pR+sF2YXV2R0ETOFQoOCODeG
NpRKpmvrF80zA4cK4MCXTPXsoYn8MOU8P53UMtfQH09iiFhZuC9GvcNabLHvc1+n
qF+cvO8PJ347gOpcAmzmSVMFsDx8lWos02TqWbvVFwJwkI4q5uglJEF4a6meIt+E
j6fIDCiKTmTnCwwexsF/eczEu92vRu/xOnua0YdLBi2TpUCgqqNHkIAdMIi8fSLh
oQh1jMW9jHyDQHe3LcubwnpLMugqzAVnBpcWmcpzW7RivQJG0YnGFHDOr6Yz3EF7
KD3QqQEmpku7wPDilFhvq74Q1qYDps3av8yFAUecjc9+5PsS5bMYDT9Y4lCoFhYD
tt+lu7JMise4IwQ6vR5/Ypv1UyAnd3+pwFgJg5Yj0cvoirzBsBAmojGRQm2h2YMa
JAHnK8h/+jQIqqUzR3ESNsfhOKIJEw5q9//dsLlrgHdIK8vEkQSkncMttoJuk+49
NBfFQFOu3Je2NTU7ggcVF+OQS3jPpQ7xBF58uIkXGFEq4W6ObY4kXtWU2DnfSPC6
ul+5RsoWgCnP3ixmSyIFn4m7WaX53TQIC174wFtc0kyBneLgQo0yGrt7RTUQdiL/
nmOuVtzyXY2iq8fiWRo2HIfrNKZmHJMQfNaiXek++CcNOnqyys0YjOzYOJ7phTd2
+xjBTFM8C4mKBXsCTnq1yewc31FWzNKDHs56BObAGu+xHHWTQ/HQW6yAyfdO9tkF
I/M6BxOjMa2fRN8SRfLfzeaiR8NBPvJBVXYLjoswfPYd86D5bQt0siY3PUSih9qL
jIDVYiqt7bHr5hefE3Q6gwNgeBJpJSphg1Fscgm8sdubFbgT4Eg7jWQIWm0ihOiE
l5wo41+stqGuNCynO+dcRF/GT3+jvGnwhhaNz3H+vZvG7IZFS/dP3fGYMvotq3s0
pkJD8kfF4hcZ3qaPmvZ0FJfRT5EJNeLNYcUop4T3v5LtxE2nhCAzadHOm22EY2or
sR7i1D5Fd+ksliQfNpzJRyIjbMBwUelRrUYm2hQGl64PAOAN0d78d8tDxg1mYV5V
Zds79I2ohuOzoW8jrkSUGaBzMFpCCXUcjCrL53iym1kaYpZQRPf4qg5/OtdreCXA
cJ7Qwy/QVUPULLzlkDInXrtfZlG/Mf1NdJ9RKXerb99RVEzji6NHnc0FTO9YyT+b
TsY4NYyvu9bqL1e7MIBEoR/FnMg/ggDj/UOb8erjSmkD1csQG/dMQ/E1SP3VtzwZ
zlKYGbOI/D4N5C+4VtBHr2+5ebTxWUxTkWWfhnngaqmABDqloOn9pe7INF10WAZw
m+zTTlZR6Uqj8VnLefr6uMcf9FwIAxoE9ihYJCZRQvvltMr3oaD8NsQvj6puOEJA
iCD0h0EqNeDiLKqf40rRR32dApl47DTYB+YIwL1AOXmrxo/Nf+8kSBylC0wYazmy
j8BiZQkkrsxl4bvWC2S7gQq/hNU8BobsXabZwOzeOsuAB3AYoRJLADMCKfhYPm8K
IXVLyXEBaoXgHAnQnqk1kNvt9fQcP0DrC0x4NxPO5lqlxUCUykIZPKqmDSSa9lrT
8RsrmpHwnXD2zM7ZEzNHYdtzk23Nk2OAB14VEICtWJ9GRt/UD2eDq7yIMGglxNus
5xc23DgVY4MECbpIAVW5DOFPfPIsbNMMrnCOVVflcin8Xny8Zy/Vs9OATVtpbJoA
xZi/QFfZo2/XUfrQFhxSfTI1IYMwPhH4LN3SsrQ5N9xTGPYw7hWDVKSPyPcKbv8h
0vqZFC7egCQHTQRHPGNkaXwq9ZnM2dj5IaXhzIuL3YXFSARB6vCdocNXwo2V5AKH
608P7LpN/sHun28WFAOaDPFdR5ziPtXzGtNNIQ7UghLc5Lhw0r2lXJMFXFOAv/S8
hTJwX8Hoq18ezFiQ5zm5MtwrPE7x4PEBJHcVvUxp5chtDbWAsjQ+duUi7Q6Vq9Ee
02konJd1De4tTyD5heKSEsjS9fdvz262ZaXcdXgHYFe+c8WCAns/Qlms2/ZkzgNZ
/iYZ9G6rEX7vByj6WuHp4adv1sLnFYJh2/wmvfnoZU2p1by0VfethIubfyda0IEc
c4LCG749kTfmBu726U161PZeKIV1h0ArPdVPmaFBeC1krut+jRUcxYx9zwgbj6or
RQ02URXCnYvEnIWFXQmTMq9Dai+7N5Ds5oi3ptdq5Uq8cr9eGLp2RRdiv/3T9ciG
s4IokHjFK4Q2+ix7nF4C/PRCXG4Ce+fqE0j3vOBms4F5syTOy7VlzwrrUHHGpXfo
mDlmKqJ3k4BensHChGZrdwQW/wHsikIwei8gRSE+rCNMPyTKRikgsoIjT7q47O7x
dSiuTmiKmpimYZXWOMCK5y0pZpw4lbjL9W/5RQeMPu1oEapR6zE31p7Rgrf5c0bd
7PXK8VTqXwM84eW+0jScR2tHqZROBVA65mvM5mue+PPKxxoSxpbqtF67DLT+wCaX
gB19kH03dlrCjK9q2P7qIlgGukqj6ca4p7gHms0PrerNPHdbk30JJeBx6/z/Iik1
ulTiz+u88s//uoVBa5luH01Ja4vO3Xw1OHr0To1O69VN8NleY3z3T/WaSCBXyxaC
8WoDyId2GkfXVirUwY36Dokwm+xBHgfxWRxbPkAdSeZvOFqjESgKG6veZDwThECG
mBXrt7Z8J4pHIDMrH6eo0jLhuI45ZDDMHtIXMSIpzK4CJ4x+E28rZWDZxlHN8iwb
doaSW4kM3KIg/SZloxtDbVD9Mjvq+I3KU1G+MxokQsOCXOoTz4rHTqSPGFCdNYMG
NB6EDEqtHxFPArqq5VKKlE4KB0nevXnLzvzbfiAuo2ZveOYkTDxRj7nwwMxlbouF
6NatvCh+t+R7+2uk7mntKGZgbkJWpzruZHGJlvXqanHI1XkIVJpBtdGQPrhvva06
9talAElaepzdLm89s+EhU0KacIPHoTkWxeX8RUzubn8N78wad4uLhewJmstsJXp2
A64O3OlVSWdtHBbVa846QvC5BghUoKWdf1bsO6DV6piernmM+1PpvYgYIUnWoL03
IZYkN67WaE/X4pmYoQrsqTEI8qfgnpbFDSd9+VyA3Ab4QLyKXAO/38uHxQuWPOJK
DVlduC/p+LlT4qZh8oEJLIwvMxelScl+W1yzma83p2wPXzNcfZSLax0L4Y2ntzK8
gHNhypcPelQ2qom5FXkVOrE50MQaaTNfseM0SNR5jlnevq4y43Ghh6ClS+d5C/FL
Bp9M5A0QvXmF6379RtD9NtYzT1kefUcg2azeQQlYGKwZ2ue4mYCG/Sug/4PjVtht
Ccs/JtyTvXevWmtlccYSiqqxi36+3qU27bdt9p0qpZbn6QxgzlVVjEmkDHxHShI/
Rn4R4O2tlphnw4MPRRCWqfIjZIOQUApDc0tfJKTKNLgCnZkkf8coUhD6sqI/2G/Z
KyJvHPSDdqgcyNbYoB0rAMorst9Ry1OW0G76G2/uSpFy59rNgZid7kDcFYzPVL06
4v7QUy5BELtnZHnORd/xMUm9oKFWlxisQk1I/Hiq/EI4t0Q7Cg3jnk3sm8dHH2k9
3SA+flnxUhmxLANLYFeeKm1IOoeQNWP/En4T5ye/Vmwv8rXaKst+GuYoxOqNi39T
mYay345AUPoySfmnbzL9e8QOCrAOw+Sy9i7UEXelM238eEJ/LvXDMy178fkP9Qa9
dgRSA7b6xfxsqCt66w5RO4kTKu9kBbquuYN+b3zBjM/cM8IRi2r02f8L4VtE02ch
kY0lrLXgzY95WK0He7QQElBCxY+cfURolgGmWJifoQSjbA2yMam2ACwoTFs7+JQS
jHbfzRZI0QDbdujYgYs23TbkVVVsOG4+MkRB6jd1NQm/M3he6PZnBGUSVwR/ogte
J6GhckFcZm7a/RL04TcoheDpXsHxgmwH+tVnqbD0PcoNtt3vLiEcC/CC4EKz0ljI
Iiw2eZ6kAxuYD2rZ5q3YSQT4CCdGjeIJ7BXvVXAWfw2JwCJCLGtHCLMHkb4Y1gg4
wnPWYbAlJ0JkrJhIUgVMNRRE206A1ju+geCZqL52CTZpvj3Y0QV3s5ckrDvC2DX2
h2mn7BWkhROy+2VuSAW1iZBzTSss+uy40vIwgjmeYoQwdYMmJUP3mpuZk+/y3L1p
gKe81KNvt0E05zCc5qp3QBBKMWLawYTBvfQWTp4u/zk68Z8Y42gsszIjsUmY9nAn
jQ20gChYLwpQy2RuOvEIobWc8ffCCOwIkbOZx/2ekAUN3T72cMHy615u5WFlLHmr
vZ8/oVqZIU6i1QdVlr8z/8ASzBffQLmEweg4oPL9rUVNAj5IeQKBuwd5xdSsuU5F
HQBChBMqZ7hqLYjB1zKj2lUfv7Tw4kCuU6ztv+4A8LdVwtmAZtvkYOzF5EmKXPDQ
95J76fyzOJs96bzw6ldvkKXDVftdMuILZxad1PbaHDT5t9u2JgbFOxwdDttcgfBD
/NhdvnU7fJdeOUaf0qPu3ME69IWywJn9qpgJMY6LmUgjn8rymJ5a40HY77W7j2YL
D9PKz80tv2GbZzUPb+pnAoRE3vuM0zWSCHzZs/t7UNqXGGdbRAe2MsdP+UAXJxyB
W6dcbTtR/UZwPNvpM/X2eObk2rfwCNX22eBUO7ouRJVDdkN5OO1LKr1+sRR15mto
9FBqgPCH47BP+w0JZKn30Ep6KeJf761eJD4Fhav/dOxWpZ6OWFNVYXDIcYdch/xU
55XM/oyMheGvlBSgH8LNz5K7cIxBO0bsN6EPj4/FDTbttMI6CvRAeyk3f7q8VWrq
zm5R1yQhv68m4ETmCnWFQeM/MyPBiJh/gbO0x9Xe8DjV5fnGSEwXbyIupRVuPPcB
r6bQWBvfq+8E8E4gcEFURXzgNoGoSmRMYjtH1hpmaWrgHlVpDsGRZw0UUIO68o0Z
e2P0kPxlIpymIukcNQBMonVzf+fGBpBpmOfjfX6r610xbKjLp3N6fBJ9mWIvkYwd
yG4NuZNEcKh1E3RPDr+blWH6W7IG15XrNMWw2R/aIdJnzoiZesyhRMRD/hlDQURU
W1OTNOzPviiZ/lXjEu+gDbUNRgkuhBZG2guWaV/OBMmiLoE9N2+2SwZLH9NIJg2D
qeZkK49JZdInIE49BqSMcD242Z0FHcmfpoUaHW9E1ndow0r1sfYUKlltNYDiucbZ
A8NZbQ/iwliavhDZzDkK5xOEUQPfIyy/DCfUfW9tQnX+wEec81+PkTdRdh3P4h0K
rUwKsd20gCDsj6sQ2xCrddVTtdeJ1Ru1bmuTYprmHWqgrefe5diHyAbmK/DPyCeq
9ee14NbWXIPjZaeCtnrWwJ8ez1pp528qD5vJ/OoFByKaCUEKGcMxwfQcCKdMDzzz
b+xs2fUP9l2S7UeMPSlHY50j51gNOz3+dd1Gnxq05xdLSwZdx4yix8TRnQ8tryEE
3l4cb47GQrWvoIIxFInpQ6NFYu8tz9RFV5tuE21x5RpYJM5MwmNQPKd2Mm6w8kzq
Qr0BBFaVtL8kuFz8rQC/LHFRjvMsNYt0SVJbUMopw5KpOiCpmyYtBLJy7vIjy9YA
b1bcQtWkNpTDA2w/oQ3ftQZGEbe0jlDa+GkqzxcI5qi3bcojRgH7UwO2PumNRd/p
ynjuKP/CerhcgTdZ9seSt2pqYxzb680fIHwAXfPWpLWLb3/RsMvty/HqC+y3Rp8Q
bWq+FSl9Ud/vuyr1Pb28DPq4+q3ZHfWAlrXhvC71pDLClXgStIFY2B7G1IRdSeNe
SkgOpaUD1HCLVayFTe9Q41oCGEj8Gq69o9qLID0vyiG77iWm17l/kFt5MmeGFYTf
/GzZ8T3ZK5iGZ7wH3Vchc9d1FvFafV8V6JI1Ga1XvVaq28wPmgViahm+rReCZsPW
WMs6XeDB2w6i36DiJCZqIGqh+Mvljw5c4l1SOzaii29Un0JFUFkz+mlqQMeuFOaX
DcsHSypEt0Mu/nh0PWw4HYJe+YE4vbUYjlWxNF4VAl0EqDcYpSkbJnj5W7/PX4Ry
RlkysPRd8PxhtUXWud03UayCihkumBfNv6fqDjBXzrKtBlKTKu3HLXzPdTBtgdq9
+m+UJNIga6Y5gokb0qMpgoeEuIMYjFA3oRFNPVTjaiEiCQisAomOgBm+cxZO2kEi
EN6soLVJ6vdeJujwoR1M550M+vsNGCa/J8wyYz8Hv3CApBPIGpyrNxPKk6zBklk7
SbSqkRGUFs1V5ycG+HBELmh8ZpNEMyaPLSNzm4iiTKgL7P9YEwMJbPRIrHlpS2oz
0pwV416sCV9+J7+s/VDw6qOh5mJeuerP7bt1JP7iHFPwaQRmvN7IZdP02rvzLv7z
pvE//1anOgHXbKbK81WZQzPW0p2DhDywq4vwJ+gir4HzvilfaZG9WIJ3BvosiB+a
EhpJbysWVuUaxS4Z2H1dBIG+F0ulbQR69U/gz0zDC76yJz9ThQHjqI38GWNSnrA3
0buzH75oK1f/MAKjQfAuZRYGTqLyAjeo+aToexMQiTElKuZEivya4WIsQ0/eChsp
YXOlDKpcHfdGOxE1V6oby3xhi+B5pqAoqG9S5L6KZsZSkzQd8iJN0cqraF406cqh
NzruV3YzY8N3AQhW+v5w3Z/dUACLTX3aENl7f1998Uk9BrxIwNigj40hx+x021Zz
rDJT++IUKyQlTpKoP3/xWMGTeWV8zMaQj7ag7W7rjFDe38m82EH8prlw/w/11smI
Se2KH80i27cQTBR21JaBpop1LLYkmWxvjKcv4He+UKuSbRzdH2Ga6k7S8Nzks1Xs
ci9IRs59KPZgWEEZMT5Qk2/F24nVqSr7E2K01bB5QFX99Uc6OdV8m/wCtIxv0/fF
znOl3TESp+HUJAqoWIbtDeAe6VId9A5yea9zuDz2mAFWpXo5IpRTI0gse18xfNE4
4w2+3ynpYxCnbsEJFjknkxJlsYM/OaDfDBdzt9mZ/UbPN9JnfHUIeZQHqoSMx/ZY
zC8JBtAE/cf+ukUM911q/bjBJE/tc+9d0T+2JD1Bwq0wP/2dzOGHzJuaW7jFiLpH
JjuM+SXDP7QOGuy3IAcwmLJSMMg+sCe8Kmbmwh26uEDLJd3eLKWva7ecu7wFaYZR
FOlahmJC9whtJ6cvCKqDwVcl53/9o0WB5/REuPj79Cg/0NkrQY+psBhkc5lM53za
FZO0HOj4wMKYHbqz/cYSG92uQz9kbO8gy+tudrxNKx0FrTijzzYM4dLnPkxpFBCH
nw+dT51a3Gytde7/GNiYSOlj7U/DlQNb0gzQ66qFtu1rtl9gN+ey+WYBCfQBz3Px
iHOtEYr3igwwK3oThPagdleW2x7HB2fQLdEOQk7+jHOyqrS08HIAlJdN2jlxVHOQ
rIwvKtD7xcwS09DvGc+pQ9epQQ23yUq/TmnLDJGdQeIl4BmAzgy/cHTocKexU9To
byi87/rlB9r3TheSQVfm0YeLdanM2wLcEVSqNzUjJsHRfjPx1UnF4Qo6JKziXx8m
z4XxsAaHGNS55I+wC07eR+9+BdqVrGKz4yr0hZG9FeG/ihj/9I/T1pFo/x/KDrYd
iHZ3iFBb4K/TVdcsTcBQzTGF5lg9Pp122NP2pwV0b6TFTSxUcLKqOr7byVMkHfl6
0lvH9nHr1YZeDPrXKjujEDjHx462uAaeJxo2CAE2rp1QJUNvFIDPqHXHutumk/Sy
KSqW1Zc+Lge+qDUk100td1K1NwEvmWy1EEQw/jwZCJG1RKbDQ77JxV8n8REKajw+
ODMwS1M51K0V/XVSSZGXVHnVdGfFDvmyL7wMAkwoyo/e9yguFm9OlSXoy8s+w7iT
wYdfELBlI2LPBsFJT3/8FrPzqYn5yZcvu0Kq3IBub6ebgrxcpedlnLa5DooFSPHo
2pTkHaOfQDhChIElE885mUnmHbfWGq/xmtXuEPAzmICNJHSd7GZ1cj7WaVURocz8
hFdLGAsARhUGYoMtHrHAgMW8Hex/3MDaGue3J8wzbsLcQTeOpL4fX8LWnC/9ccDr
FaJqvG+ljw0+d3JVh9lQj0/kIjkCuQLJjqDhhN894dSVVjFNAv05EHiBDXW1jprn
Rwin6JQ4vkby2L2scUMl0qsXdBmkzueRnW3y5nVz5dhMUWShPn3EbteMwvvHDxab
Noyxur84f5mOUuxLaK6QfW4TpEFVSn3yFVc39YFK+dNTWXvUx/LfzcFKRI+S7wA/
yG+DfvdLLps03A71bbNlC/PBuCs2X3bAkqX4a7I/2GN7AZ07bGTVhnVlETaEi/gF
5LcBo3Z7knswV/03jmEanWN68CdT9Iu7/wgnokOGDh/O2YzCpD88nYaXa9vgGllj
lnAL1Q0NksVvabHC1v+i/9VOHXbA9mhGon0h2qb4bPy3pR2J5pclmMYjNHjEJG0H
gSsSsEyvIS7dbbXnMjY9cqGPkS6A3c7+wijIIPLhtW58orIJ/M4s9m3eb+YQ/9Y4
fpCFdOTIStlvIQwJ9eIjBrn1gWCh9GSd4SOqH9G/JYLXexjuy7TQZtM2aJhLN/wG
nXShY2/OgQZ3w/zJBwU53uON1Zq1QZ5IKuiPjRItikup1FF9OIvgRqnlLx7KoiE9
WV7n0GIYZoPY8P4UCmAedUphrWhWxaxZ/IsN/cCfx93HWVRJEE+Z0k3qPsPlCUP3
X3aDvbHhH0E+kreW0PNsANq4ncRX1D2krc4Kh25KMn3227UP0dfXwge7dpkLPlPB
FYBpUuUL9i35Y8yBbk/kzzyYlR3GfhaMxBcIQlQTXoSuUaEvG5tQw7uV1E1IRhPx
Tkq+vUcqJod0LKSQJneG9oETnqmQ4r5V9qfwwsRV7qy+dlPWUX3eKNvSzHpFk47L
JB8BSgPI2leVPnHc8oThu+0ZF8uurbibFflXUXLH+QXukgag7sedTRzzt1WIDXpc
jpg5BMqbeknekm7t9xhZdhX/l8yM4IE1bvywZIYmrLF6dSANaCBCPkO7DA3OUK/v
7wMCTiS7Gh55qyy0ZQ5MiWpR8Xgx6rt1p4f8J2DF6F1sO7x/7xeL1ETKXB5Z1o7V
w8C336q7+QhcW68oJrQsai36z1wDUxBkNKOE4wteCkVDAMf9bOv6Vthm8gkC3Iax
W11rsI9FZXSEyf1NaMERUmcgGoPk6D+F51ZLACe1F7F8q+Xpzalx6DZ057OfB+3a
4YZLU0KMpAmcmndbRTrWd/lcJrNfcqTKR02G8RKjjiPcFwg2JuC7+XBuXx0O+ogT
nWJM4uHk4PRb/RzcFfL2oXKjpnV5FD3xalzCAxN4y314kptpk/FUO3FVkNyFZYni
FxfFKtNkPIvOMSyHuRzm2UKNgv7B9J69/TuTabkkSA7a6Awzm7IRCXTBeS1GZaT4
HhJkwli3Mnq+SgEw7Da+dCCwHg0GnY0c7SXb1vzsi3POrWKTRQbawMe2L4S3SPVb
w/lQHP259rGY0ckzrQYQXGou1iUjKGs9rV8CjlPOlw8PDJBXzemDG/rk/UZngoYp
cRD1wkwgEPuXBAf/N6Phh6HN1EHNPbVX/XMS+dD7CXxnZXu/jTehjTqsBVeRvzM7
t1Q303MgHuy4gMQO8TbpYhVaMU8++ExMAhtsAW6BF8eo4q2ocRuHJ0A+tA84Cib6
ge0TiM5wqBbGWOluVZ3SWLm9DxJ45kIPRCg6JUERIzuQcw52dorZR+xEqe3ycPgJ
yfPVLynrTVQmsLH8D6Z5E02foCNlVYkz+lrqHddfjD4LJ3A2XbeA+GdNoOqcw2Ed
EH9MErjGSpX5daQtCtKVSpgjPSdZob2r+Gn352M5pvk71akTcWHXvdvKHenuNh+9
ms2LrNIJNSfywkieH3ywZzueGNhHIBeVWTZqCOaKRvae58AclY7dmZlKvbUHrKmJ
68JXooYX3clHmpnH4KqWgxvvsctBCoTUlJXmHUi6Imm5etQfrdOv46TerFuKQ78+
06Df1OCxPQb273tGRoJYFetQgb7n+SPKWlyc0qJTVBnZcvJ9uKoEM3l3nczul+/G
Nj3mNSq3DRK6L5OSNCCKgV3JT2gha1UDrdWA4IPzuqIwiziR7kvAV5836yNRjLxF
PRmU+/QAZfRdC7se2ngm4zGOR4cHphoEwCc+dbUg46DzeijyYK7nyGlpo15N7AOr
2z2rx/sxMteYW5kNKVYG2qNX81aVJZ2pPhkFWR8+cqactGIAgH7JjJQxiCA8vXeg
AhYOZqXrHcNfTJT+na5aBfG8LJjPfBqDCYMUDYYQmyIslKbF2qmDctLTmF1ECuAB
CJ1wwPNnhKbYfH/CqS2cyS5M9PiTKEzVQ9+pgM0yXef1jLpTKXCfSsia2cUo27mN
6TzhC2rMlzGCWsZAIjbZrmOkH0N81N7kvz7pxAF6cgEuOZNfHC4TFWw3Q/JLBux2
it8zB1OQMiDwE8eCu/NoaAsQ99dwg1H8oYbEV/QgncmmfEtYqV8T9qP73fLnz6IE
2YMkEpW38YFPZTzUvW29VrYFRQQlOVZnQ4Fz/WTZVsHhp2Hrp8L7GCwT5pKXZD5z
jieOG9PP5ugp+ZlSCmB2nNsf/ZuP1J/ZpgmyWeD3VoS9mYWztZaZL5iae2Spze1e
sQB172pOCbLaUGh9VpRbH53guSPfnUTWur9g2pm4ZXjAN9nqWMhR5PP/AyMCauxr
RNcMvWfR5+Y2TtWrBefCb/yyxX0F7Q4gcn2hfxm7QgsujoFgvjrkTJNz2dTQYFci
gaEmDgZn0dmdRkZuTVHWe0+fJwNA8aodkfl47VYIiIAEMIx7NFAr41hoPKKwohKj
1UbnWZavXawp8fDglJwThCRBUalMEmkbM6UFLdxPiRqRzWzsL6FHI7wlDMVDSP7N
BH9AKjUS8lcFrrAD7SW2vlBXn3+MYkpfChFzH89zpzFSf7w9wDF2zjKDudb+0Itu
sYTzEd/3tzzKiQvJtVQnpGPNtVGz9ZffNp/Nr5g6Yc5cG/SQviAdzXTd6oAaxfLJ
NunoYADDp6DXeqTbdd5zQOnnds201q04nxTbViqHTO6pgGN2ZvVOPFhfmA3getSY
BkVGJN1bNNTH/QIFMvbnhmCqZ+cyzFujsNOjM/1eAo/D4jSPrgxNtlLnlIOBoNVH
2PZFoMTXMg99UnlSjPfLA0I1WPPj0/vq+Ch7IRt289Ko6K7PG8L1uA/vHPeU2Ilp
5NzWMU3Ap2bc1R+3xoC70ibItNJHs6O4Bi7TazfK48MxjG816wq9X6WxZP0VcHhn
uFbr3t0ZqxlYm6nv+/ipxCM7ApNvE0h950G8V5xHvHU/FOsBPovmZyqKVtWtAsAw
m4ohyTji/lH7uen6z+bNkGymKITu011ruGsxWtDjyU/h37IXgrpV21zzK8+r4Rdn
edxLImNAWLrBwLFiqqYIEIPRMm0NB3c72eezBG5tRM1yCIJ3nBsriuWZPxqgsOrp
JQYpQLPm11U3kHZgp0B3HNjXUKsvwo4ZGGNfABhYjIojK4h/m8gRKwg7DVvY1LwX
XG1x5XJvVXcTo/Pe7rZKXhIfb+1XxDoNgnIATNGf7kJ1vbFVkhyMZD7hCIw6Alq5
hnX8VOO+9RmtdPK5OG9gfUMSIBdf6U2dNjgXuqmonBZm0xc4ta17xrZoYcEBghtQ
B4kxxkaVlBuRAPBGbtxifm98d+EME5NceXbLiUnvmo/59SOkO97LajJbX+XrMMT9
F1QICSS2mXaP5bCSp/6H68P1kF9jTVjxlqL+6PwQ5KpPoy8Eo7+bTxwNtRkhjOSK
626bbbJvuxsSiMQj8bUTP4wlSTZ0GCOne+Do+B9dtpjNWDy/h3G03Ev81p53FMGT
83pe6weB+FFvi1jSaKQLcRQa6sXNbptIx5LH72z8AyT+Vrv5t4FYKsUwsri0XkJX
sjKobQQvxHw7PmFfRi+nuTHH2ohXEh86wOph0P/l/hg5uaVkaThOaHvOdele6f2N
5m+5wTOFNaXOvMUGif+yDsIE+/x5jefKnNZgMz2Xo7+7z+M7UUul624uYuPaRMui
I3b+qeSumvmU4jVJEhxSBbaSbZPjvZQdwEmgc+U+luOubNuHxLIZ9SoU8LUQxpfY
Y4ld0EGNEkqPUHNiLoRuDQXjAMaA+Wi1MQpGOjuKeLNT8ptgBmUpqFS37oDmGGAQ
jWq/1uCO3pVsHzpdB4XDt9Gea1F9ug8/Lk7zOZbG80etTzEFKfxdIinKPKhVnCLw
7eTLad74PqdZRRE4IoY84540aDZgJoA4ORXnBS2AC4ENR62qqs9lb+SU+qPejZ2t
jf54wmReLa1dT94Gcv/e0PyBmgt1gysv9ApuHEe1QeVRXS0fXDw9Mt7RctAKeph4
1B5QhlXQrj2kjg5PqNuatDDMnatBjjJ2Pi5m07KmMoq1/YhZuU9V7b0Qbz7d0A9L
7OtkAKwTQyzcvT/3QRvpMWYNtfD9ta3oGbSqDSLGKeqm0FM9ZzHyV16lKC4tnQSE
2+iISTHk2nQXJ3kDyOB7/26uUC6Uc5nHFK/+NT7Hs35ABOTdCPr8cWVD4MTb77Jw
MEKFmlg4I742SsF4FMtaUJFIIBJ65FSW2gJHdCpNiwoWRT6w26/8/pR2+Ucj43fO
MBFm6vkPTM9HlUjVeWeWP8AEeyf0EeQaeKBru8uBd1/c0/621Ucqw4CR/HDBgfG8
7JASrSksYriuNYZvZq22yh1IZwoOsKeNUUvnW8pr4j7DwSzC58a6jknLjpw0/h/3
uHcs8rbe1vpGYopBfGw2txLPVJwhHnKLmWqZf0sN1tUXFffOf/F0cejb8AlaeG6U
JgM+6Q+UpLjr6z0gaHw29ChUwRh74MBxs7Gzl4lHHOk15fP3jtOA9w/JH/5V7HSo
/jodrPNsmQ1fNSOuxQo38+0K/xTZJGgbDSSI5DdZsIxKAYCesvDWsGA+jN3OMoUj
PbuMs4iVQjmpvmMu1XM42ggOO0LwsD1ek30geSVteYco0E2OMlTZnmtWPI/yEOIJ
Tjd5YE9Xfdh0BEE7SEU6NB14uLQafqCoqgUnKB6qYrjaRqz5S90u2Yt1hnclGN18
JouL/rGn9a919JIPKr/wduo8SDG5UarSXcMrp9Fkj9RNkS9U/D6KVyBZGmqHJShJ
orEbDQRoMdEu0T6tih04WoDo6L7aMOU2Ei317Op9BpDocFHcMQ0piCRZagmiRAD9
QgDhAGpOqzTMxBxwjDVWgc/D7Ypd1fvPqJ68LM0w5GoY5GzPJJ4wA1YoZL8A5foA
JYiFexalB1tBUfcM6Kpiee2UgKpy2ThYzh0rkuntx8jBQk6+Q2YDrRUe6IS9DFGk
kGhhfVUelSBfp5//05bxf4k6Xad2kUNdR32pxGOXAAt90328rSwK4U6cUcWJo7yK
1ySKPYMm4IHdLoZ4W8e6mN+6EpnU1ySs1EvNmJ1G9O7MQMSiugaGyGot9r8A2d28
FbeuTf3vHJF02QnNXxz+YWAciAHcjMk7o1vYA+JVYFazQkC7luY7mURgb+fIVpb+
4awGoJIYdqDLhZQhtyw+/ZyLxag1ONWZTDa/REPH0KIR1gLwE42xjQuASAoNNGX0
RXe4dtqmj95bQ/TPXKwQ1SUxulh+ynPxsE9fRVNkDcF2/gyoCH/vZenefLlN+xTW
0qlwi7Z7tMsVabsLwlQ3ElnO3HNuvcfzOCUfBy+zJZ5BDsaVgfVy5M2ZC022gEw7
jeSJ2D7tMtFvjsybC4qlMsSAOmZo5CCGVKqWW4mdxwUxss8nKGREdLAa+bK6SJps
nyTIWyuHiW+1Koi+2xsZjviMsE+Sp95yI0W8uIzoZwqfs4/dsM6E1aviPMeunuuY
Jo2shLbw8jilZHV17eXVk7cn/POvlzGtJyuErw6GMk0JSx7C+6NvlfKQOS7Cstfi
Y40CXADAncYRmSRDe2FE3uJSuQYtvjPtrEYrKzR3ZrrOssGSse3f8VyGpcV0bDzz
IYX42GsnU7XJXf7zxbN1dNFUCjOGaY+xRNnlJ3kkIfeNUmDDTw8L0Jmq7a29mTMb
6+pki3VJ3SgpPyyW8Oj6nxhf3DXrxEg76UT8Z4A7lQUcm5lJmxqMs00+qcKKo6XI
ARWIT//+yY9AxJq7FVw72P8i1jnoUySA7BxEITMajzIOXyvrM6dd5NFMCXEx4YFh
sfI92mJAOrQEXcfxu36Dpe6ySW/jziXG2KWV1FxJuivFQbX++sQHV0RAew+IhImM
vnbbMa0u56EK/XHv7X90ECpPh03JYJnHeLg5Zjf128EOPx9KZ1MrDvRoXD5hrziX
vAN7TyjZqyuzwEvtykXglcvpQU9TDpcG+nkLqK43VJoJTtUywY04Hp2m2lgwCSkU
jycUEevtumNsiHb/XMKVtXnToYwxhB1Tlc0/YTAQ6dAJnPBIUkSqND2rV14Z4HWU
aLIlMJTAfI8b/iAxjez28vI3Hbu0ErLzGBqr8k7750e48HvixmrfcKnR5VdIGVp4
KQxf038UF5dA+GijFBCJ+Na4R5tdw3TAUOWqh6td9hjoghAHRCFyVFpyU3eW93eY
tHkgdb9V31CYzXCglJ0CUKOXDJbNXs+AwDGc/lc42Du+MFXqHMje4N2VJPO3NwVF
Q1B6mCEJQ2RSqJ1jUlsi2vCW7ehwLe4BhUynL4LHAtTMk0/uFX2dD20WuTKYEmgg
4qJtsU3KGw7TD8uVOOkUf3wdQn3N8ljxSYasnD0YnFt6NB5JusW8a1A8tB+umdOe
nOfXLnQ7jxd5lJlaje3FLBeWENjfPqSSzywSDd7/nHwk7f4xVD8+70jpWpD6hqYs
NWLX39UkRIrFbK/8oV1nkm1ENPEMsrLzHAfmMod4YlC2/pkHwKF76KRA/lfCoSxp
+qcLSm8Yow/+YKobzNUifxHB0NdL9C9EJCfvyHN5yw2pGrs4lNY5OvTdRWe4PxSD
bF0PXHMwmrqSBQjVtLTo4LAPm+FcUTp4UtzCAscLeGYL1p9EY7F4aIhaFcaqL/pp
F/dE0QRCfmr/miw+aEWcDdxR89wiHoPfiMUWbIWRSWx8aWa+dUHtVIDzf38X75qi
CRSBMRTF7PfsrCmV7hqqQu7hYIPMsL2mSB6iUhy30jQrfEubhH/d20WYQ9IPGnEK
zs2r0P8SyLWigHVl2CG7JQ7bB47tmTlXecRcQ732bxT7xLcojiJq0OTD5ywE06IZ
lSXJqjd3YSACgA42zUNy5/Q9mhx3ZmEVDPaajzH4KEUQJQqS4xdp+dQaT6evX8/K
lLJBC1HmUCh6K7o3ivDITqZEbsZNmpRfmNFF+FLHKJ1CwT6cb/20PIvcoK1MMynY
nkAXVxtd+Y5DUsgxlOUm18mjul5y+eIu4aKlcdSqRLAFWcPLW0+hf9rrTz8nwknz
IokTOkw9WnK5InE+mNT5j8/oPdtIbfvOU94MT9bZax/JRsotf9JRcPR/3g1C6FUW
9HGpy04DrwaoUNbnTIC7N1JR396dFfy0IvvJ2O6ns+od8WtPvdJGfcJecQmuWg0M
00e6U7H7JMgzD2rIdksF3eCvJygPjfhRnC+D3kNKPTBXWVK2Rua7mNb8LawaGe1l
Iy1mILQQTXo/9uy5l4/7QFxGP2Qf/7/aKOpV0EuzEVzDYz4cY/ooIMnozbwTgC16
qxuZG+XJry+wJ4OY/IV3WHrehs0/6BEfjC0GvA0kX9YAldgR1BHvbkfqhJAo7yrx
kIifhmR9TR500wwy7YSOpz9D7yfKZYCbYY+ecWjylZHn0zUT9N0luGTUKlLvK+h1
1GH8eYNRE8sHqO04uxEBmAXOMufw74g/OEVzBIjT/8LbngoeP/7cbiRa8JWNe08t
dd9w4y1uq+XocqKfbGLkdZ8i9BEENxa7T5MMI9DNpT7MJyLZcScfRK0RZ8pAP1nr
aSIxokJ1WN0LeGlkvhIfe/wMqDK4+xASAI+abfHR/meBPYFsgdCoYU+/Zmh1Ox8E
1vtlN+ni1bWolkkq8w88WU5lK5nKneEgPmUFZiW5KkKd7PEgx0jCrACOoYoOvkjM
Eego4zxxhEpZjNwfiLMOWueApjcclb2D/JPBVkftcVMHGOAGNOnTmkOlw8HLOjOz
Vx091PrY3KzSIZDtT74d9ozcGBuB0VHEHH0YTQ1JGIkVx8FfEktvh/OPAb+ENERy
TCBM+GQ+Sd9RtpcPW6FhgkVP8+KZhFTy/dD+T6IUMtzEHCmdreM0PWFYtfBlFJeo
Q8BLd4+c2lYDwgzngkLyXOw2eI8F1HSzVbkYW9TpGkr2TRqoqGelCtaFwJLJtyf1
5pgqjH15/E6SgXg5BHgukuDL/pY6xfbot/1wVGbpPuB+Ev5NVUIaC3Ayr6pgl7c/
DLo12qvnWMywN7t9AqjBIkneGe97c+7golQCZieHGiltATppeDwp7QoWJvU07Fcw
+HUxq//zkU5BCBia1Iiu/GhenhRhpPohiTIGXyqcby1i6U8/KPwZtfb8l0AIAUpU
J5h2OJDxH75QbskeVrubq1qk2i9Nh4wW4aH+Lor2YkCM2q5Uf6aLabVXU6sv5HOA
FU7AzjpD1+EMJxEqSre7ptlhtszY2LwEwtfXVXnwodgLyuSbFEmZ6cvDmMH/vlno
LHqeZtkX12UNPvR2jte+9mVOvkw7hX98LsMxJxM2lLzN/ujFFnHBWiyGPwAnZ4Gc
9a0pUnnpqYd/JXjSYncxmiIBnm1QLjDiXkv5DiYI1wtGdk9Arf5sQ39ZQlJKaHVL
HKOkDRohgpwSfQgRcxL/Jp1kT2dYF5qf4BG0N4wc6m6jN3NB8YR1VMVBt2RLiTH5
6HFyJMjMD2Yrsf6ruNnGMp6rIAHSHK3BVZjKPjbfFvvKuHCGwRPJnlmLakIFDXX/
ZTvLa3sbWXuTWcxe4E/LrMKOexIGqFsALsZ7mqUlN0uxh5Im0/Zjcrq0O7HUsd0L
aPP1UkWjMxaIf32N8UTG9xQEWA44c7p2RbsISGlGo7g3aL5hn0b/cm+Hd6nZGD+x
cHzQnFgNcNrbR4iCP0M4a6WxDba3eEdwey3Ani1fR4Y7n06oOOhZm4TmOVoKmbC/
EonqU3mJZpyToZvIW2sMIfJ12zekoLdn2BdMGU9Ze21cKQRxZrg3gBrTudyOI17L
6XVC+kzfVNAK2T4hPxEbq2Wrxd3Icqe1Hyj1QLpngDJdWFwLtfMOaeGkGVBLm/Df
a8yyLTp4hI8aV2Gk856s56cEgdADuuOBGaGfkep1Q0tTkhPTgKVSyy4QbWYxED2a
PYdFFH7QDSamME/A1CDXlY+BTIYuYDxwybvANDTNnlADs8EYkiEdGPAww9xUJeau
qOG3OTBH9TiF86+oYfs5OxQC9/hQAhP/EgKy14AfArgBtiwFXzyG+0M+Ki3EOb3G
WCC4UqtQ4PeutVhVE+cW7JSOWfDh1QZC3ERWhv9EKGbnUkIxEgX6Synt0sxOeKxh
vm7EKcBmsXygxX/7kbwlF2xmraSjjAfW4MY6UW14iRJyOw7/6irKG/At4ce8TJtj
DwpMpTkHc1w+vy4iBa7nibFWBjQf4A3X4/vP8teSZbT3Hzzug6bbjtXDpEVZoKcs
irgKv5ome27qb8M655S88wa+VOov7beViNLBSWCyT5h6KjgqmmDXoAvd8jjcTE0s
t5g0TSmvHqpYse6poQjfrYU6Bw8Xv3w+MJ+/IQpOcGOFPfeGANGoZqQOuhjVrhP/
HV9Gl5xMnSkr+/rZN4JGW+Az/4hz1LasBPe1jCNdde+qPJkfXSpF/794DWjmZ8x9
G0IYviLjZQLuUd4EK515WUFCsULCBRjroE0h2+4qkrrspWMb1d/LP06WO+5xOXIK
sn3kJFQKKsrVVMkdxo6WttS4E/tF+K8E3Fl4d9EkVncgDNrSpR8FgMy6q4LcuuM+
kezVfEuYu7sqevBNugRSwA/2llWs21ar61gUWErwu/RNbYHeT7dHblkZUfLtVSPN
zFFUbSjft+o+Ijp4hjGmZUNZcwvEPdg4I3WrDqVmjha0oIO15jN7hOr8yLC4sCeW
UKez1RJLJ5iUA8/Pjheo375kT8idcvCBNGpcaGBzzDrUej2u5jrJf9eVbnjZIyA8
83hWbghyhyUJc2ciu+uoS3wGFbFZZddNtYDA2oCH1HlRxMH+nbde0uKwKqbnigZT
4gQYDkQ8boqTE/54oAV88BoLaU3xmJ3d2zmeEvBeBblZ2pU4C0fMAXu11N+68WuV
4GaRyxr6FlpCVydzVEvTD479PpPFNeGUSmee4skFWYa3FVTRJsH07vRyk5ke9By4
kRWSYC8CrCpNikkxBI/6UnGghGCxUW85aVy2SkimH8GqwKnKPVNXBhL602sRqKBW
QQrZXYja/FKB137XMi8jpXbpgLBAAQPZVycwktUgTYCcFedZ6UDK2UsZy50ZWUi+
smBYpmFC9YSKpqe9USyyPEzmuuwT4L1P1Io03HbHowvQUWZj2xGnMQPhwLBKGM4Y
kPVfWptgDmOLY7Jg8nY7XGE273STeV1wYys0RvqCe1ofatzGsKq33FoSqiuzS0M0
fSPi6uHmNQJTf0DgjjeOi655oRAy/JAuRrNeMN0hUTYWO4Hnz7hqkG9gz87Ls1Op
Xwr1FSRe9Fl0oV3AT+AiY+x08ok5zzu+L2L4kSGnSH5V131/542OEmcW5yxdIpRO
sePQCbF9xdh+s7MstCIzC4s1890dX/tvAIJnROR6yRq14on8iFWio96Juvwbm0PG
0UImkT/VG0m8W5F+FJjH/g0FaE+OLcWvXMgZ8EdnVEEDi8p7wNhAfteOYc76coJT
r7EbNlMcmc/OMPOwXsFU2/2PcMy/QLZolRXqXqFTm/PxnJzRv0fJ79Dc0Zhdy0sZ
67FeDxOUmfW74Q3iyRS0f+hzN+cnYxLIFwwDqgaeo+ukuyt6giNp/kaJ3d1TBLrh
Vi+cpIFMXB5T/ndrIOxyP5oqIstedAyXk9UUhZ7Tjm9MrC+HLvrFfvcgPs7p9+7x
YiZp3o6jfIuAa60OqkHVixcRX1KFfQ8+GrGETYffcuAOK8Hm8VX714TtMc+jfxkI
eVmXWWtyZvbQKVHqnlq6e7HQt7rRmA4mmnCt1a0egrbRjxDc/u144JZAfUzY51Vr
bgGqnDg3IBxi5PATRH+i8n6HpruB2oYgQwNvtFiZYHcBlKdF3QCvGnIFPztyW9n7
UjDrJ3k5fltLEZd1hQfwS4gFxaSwobzXJGaxdP1S9nxGuoSdcEKZz8ZZg1Cz+QJg
TUfP6rYK4OwggYnGEpEihxwCNdJ6OvOhAQxf+I6jJ2K8WvlFSVfRgwoFP1Ecm5+p
6GoeWVUsHEQJ2It61yn7OStOvFbAN8ef0N9zhsLGKPAMtIqwAy/w3sxBBib3+9Wo
g5JVfAa2o4rwZ0ry/hjW6rlQZ9RsPfNclFjblVcBJkAmzqFL/C47jQCkX5yK2/Jd
Ft6+qKr/RM5/XHXJrNYpSAvhnmX43qrYvmnbHGUWP3rJPnPjJH7+BidDY9cudufH
JOxV9iOrruBkiO8X19wPc00gGzWfr8WFAO0eXP1lKbX3cC1FdLJ9X63VoxhrsOyt
INiwP4jGpLm2MCRMTpz2B+Y8eQLt3fBZEM2siEuT6JXB8/HLIRhEg5+ZtHOM7TNd
VGB4LxcCNxBuVNvfD5vMjL2YgpJserYL2Z8BWS1rGnVi6wmTjrxefuOG/rzKnfwK
LaKtpE9ok/f+LnoJt9z+qBNDHHKyfCHM7GQ0BCj3eYnQt0BGJYMkDp7zrHiErSPs
mgienOeIL/JJiRtSGFSrBRqPdLjrN6FMWZxtxtZezkk7ay4oGB0Qw5+XlOCrrTkn
E8m0lg7P98eZsgtN0mwgzppilMZbHbWmOq9RFnn/p0UyUWdVFlj0qgwJyCavZgcn
ywZM7+R2UojicnehQnG2cQT+GO/OMdUm5vUWGMgwuzZfnwDa2BcW+TuyJ9QoH0eG
QdeV3PWWQ2muSUf0uPP5zuCTNuvrOSULegna6LY4PbZbCnbmD/axfQ/W6wS32cVO
DI+Jg+AbtKKRDBVpJhWct8yFqaY7brwsKcThE2PmFUAM0rZU12Ev8Hi4CeEUfkWV
2BEDqyUDEv5H9W+2d5Y9wILQcT2o79qQY7TXs+Uz+rLGbXod975dB1nuEUlN59oI
nknzjn0HTmQ9ueRIOXkKGr9r8OZnsE3JvLW5gIqtD/iddeHAcCsBqL3CgGiuOU1M
m3/2VmGboDJisPmJ0YYByAJSLoQny/oMGP54/5m1q1H9Q+gahg8P9IqhaJwIdZhc
R0YsRjZcZ+Ya4NDEVqP/t4pfnGa0VtfhAOL8e8ggjNJj+HaqdwU+14yxgHlSMoPa
DJhk7Z5ufDQjknSCMvROBkIwy+AZ5cj4FlI3sulmYJHhJkxLz3nF+sopu9SDWsGv
jdQWdthwvsuPrFVLcNuJLtEaOZ60TJmCbhNp7U/gGBEL/byef8bjsIlNUrO0M0Rj
GHYKve9cdTXg2hCtoG+13sii8oFGOD0PF9568pfWAK/zGEqkmMwT7gz4BUkm4a0m
7GDyUXYVhU4JyIlFcXiuopfyP9pjkIaCKQLI/wmhTUFuXga3wtcAVi5edFVTGW5s
v0cVi42C8uBbX+hC6jSa2K+AMl2MPv8qqADaORzkH6R7Tg1x1/VmnLPYtNRlt+xg
cFSZe4+l6AWOvPwsKyFDV+4E0z29ROW13S/76l6ByaMcEJq4zIfAYXCnrPXkx6EP
8xcGElnVqx/QUlb55qnR8l/7wv1jhxd8DRURKsOhBVyLsnOLQgRadVJ16rGZQ+pN
ZQjxtgTBrJNZ8yJiyyHThXwhB854SM7Xdtafr9qryf/5y9C1Y8TmdhxEHTzjbPr9
tit0+B0dGledqI51qDmh5Fv5Raa0yfkZvQRb8jIsnqZpWvkWC4PgVPlA5PhKDbmz
H3Gqk107CcjilfudvDoVlsKIgH0UTvJR+sUBR3eFBsnY0D1wYmPSwkeASeUsLa5r
kewFAm4BDcxbxs4A30Rg+wOZWM9H352NCTr4SwP5lDkxHhy0EP4IkI3pSBMuMjZM
gan/Zxf+1ZIh9j03f3+74bLIUmOSXDHwU0bQD99ODbjXZJMBth3eX/+PWT1lqgUD
jYnqmMUlf7hPnEqS4xTF6qLMdf64nYx78hT3efxOGbHXGi+Ld71pbDMuMa17IrhH
/SwStd4SJU6jWlXA8J4L07hNF7GMZKzAIDfy5dhTlt7iCDzMPzq5YaIfX4Jw+nZF
YhQdODhYWp0J/ihaXRFWIxI9nFjz42gnLe8xCOvPDKw4LbzdfUwjuW7tZEazIS+l
KRY6Qo4nYgt0CKwXe4jJAhAd5JHp1FSYKvWMXmCT78lyWdyyQgmUykVGO8+TylrA
MKwgswfV0FNPT/JMIxly2EKFRffAaPpXUvb20XEJ8JW8gd86U5mJewP2/XA+39G1
HHCiNon2NVQfBUosfab6mPr8C/w8ZuGHS4Caj9QoN/gYeDsdKPN53eay0NerkKYt
LLDyH6O1xtNm+mCnTrqohI3Pl8L292lFs7Aueg3S7Qjj7Rix5O2nN8WH59hZHjsg
6Viqp6IFxMnOCXOWBNGSqRcD2tH0p60GpQQaFHQ6ls/R/K5fCx0O46Xie8PNp7ZD
1qfeC6M44zn/ZhVBtWg3whRNKNu4QcbQ2uE1OVFYQgqRWntoKY3KRvzCf0SlQTz2
mL659FsSnmeRHUwvLoMUtaj439ODtMxBqYbKJPJ7377V2dK25/f3dyxtVac7LRTE
IHUAL/fXn0mvKY102sJHbiNGfus6xZkDblkt6wZ77Lbw+bEiFGf1lP3K7EFh2bQw
de1GputW8TD9SocLgMLhuRYAP52DkMTIgJnPpHA7HNf+jGPUJo1lW3TFCxsUzHyP
fhuxsusmtgE/HXPuSNkPp+gg9pE/rfmsv8ikvEyUV+EqyljWElF1Ep6zeW75p5Mb
K6Xg7+RGLZrJZ26Oow+ezIxlakClSnhspHQbz9fp3FIE+b89Vl0Wa/dm2VuguPTd
ktpthn9orAuFLmsEMqbcFrhmG/AxJj0/BfezHgke89ILrEuYw4+0IVJDFUtR48UM
BPaw2Z+V1zFOExXfGUayk/IuPuIGdTuXXcwJvxyvV/l3tNFZMW4oOk15tSqmVd0O
psb8zAmb7vCvWQ/VrepEyupyYxUcgk6N+z7y+2xO0fpwk+0FfyppUNYmWYB/OZJZ
Dl5pv3ywOlzod6LbVwUWkww/WiRRkUPuFdZWHQDSMoTFKiP8XTcHjGNoiE4pziL9
Fubb0nUcAvQsz3Oo2pYCQN2ibEc9LaLS0w1e6oMtwTqwTkcSCkqce2uz+gfgfKna
VfOECWKyt2XWsWXcP4tpQgfNXBBU/UNxDYtpD/MuB5rtwO2MUPijY1LpM7WZ1QVJ
ytfnur+Yf24W/VoLR7nDSPtllxXONXNOa3oJtS9BrUakJqagzRLc4PkK4CIdsPGb
YfA5FmXouztZkC+Pr3ycZyBEkGvfjR2GHKG04859bseuglFgpqUXjPKGDNcN1hj3
Wh4PJl0K6cvoQc/NGZGSdjy51pf6aOYzP8joZjgGX/BhMOnuitBTQS6OIVUtImkK
ctLoSjfniIaUTycPya4ZBrt82i+AkM7acHu1mk9i3UUL3eLyFzYRdiB5r5d5tQBY
C2gku68nJZzpO+MYxhGXaG5chX8SLShDZSCclm/OHrlwv2LYRTnGwdjhB0muE0EB
SPxAgM/uDpIImqLoNYrkJKqLV2Xy64vgMeDN6ADD0j8dXRxikzcnw5UoADUDKP/o
oWWbYiLeFgak0uHLOcbrRPxNsBvV49PXaTv49efPUd9tpntW46CwEjhdLzmn3yjx
WBVxHelcjIA/YOdHkEe85/4C5xVcNK5v7rIFVR/24g5byChIoBqNs63y5oDil9lG
pW467nV6HzPoMuA9QprUfSYq/tcyVMz+D3A1LJQ7Hi83cAdW20JybtHA0ToMhbv2
dWmMbJXxq1+BBHj8O3ywqjAReMuf/1Ftz2Neqb3MD0Gl0vlxntW+QDRrqfKMDzCP
R7uUB6LfM6dwD6FPjbIq7rJ80Jsd5s7yIasAsQ0Ih6oYoQmgnOIxDcp0s+XKi56c
ccD9d28n2UeOEBAZ6ixBz9dp/vX51fgvwHektBx0qHY/e9LYCBWZmfwnT011e3eO
gC2WuMFSmkB6U3M1GoNgkonjJRP4ilZlIFebJB4komJZdApXISgIKuTlyjAkmDE4
LaXWVDA5/sUgmLCpMObib/Fq42rPNGXO7KtjWPlGTNKQntNx4V4x+pQkkk9ZZMxK
Zfp8TYJmrba/XocKI6/iDU9NN8Dpnk9IdSYCX5JmXv1yNULT4Ik62jCVzZsZ6gpB
6J03uIIK3HlA0xbmPiUw7SkLjJfssZu7TQW1o0svdrMIAvH9tY+0cdde/1XtonXS
LLsgQKRX/R/YKg/NufQog3+B/0nnv0B2Z2QM6xF9A8xP7Cqn6qIVGhWgkYNZ2Hij
gELuulU9NwAJ/bGXS4K25xvdnFyp1gRtxnUYEcNLie//kaHG96h/YS96dtWeHOGR
UGGhJix0RR1nOR/mUawKgReD7SlQTMQ2l1aJ/Mj2HZH9VzPYdtSKU7JfTcKOk6+5
eizpBUoW30NbWwlVld1i6baDLnzhMqpfkjDFGkVx6K+/DT1MuFX7pyYipX33JO71
uxaM29O8b23TCWGsvT2JK2NJm3mZyRmJPnlJwT8a4mYulxUynRb3+yWfyxZXgR9c
ZNOs/T7/YUfVmKRqnbfdYridAL1PFaFgB+ux+wOl2RgBsn3ir1soZ5kMIVK/4QRz
VQlO/7KT4GD7k6uG60I+OY3GFVRng6N28DCpj4sq0U8QVF5pLTpxne490U5T2ncA
MY5HU4ES3t2E1HuWNIpIVOxfOZiekfSjawyizl6d+WaLQ7Zb8rvW92TjHkpBXp5n
dicefpeNgi4a6QnI9V8f+3ZKDzSS+tSG2zJBY49dWWkdDJ/wkShy4DP8zY8d9Pp1
XhA0Q+GfekiiujpuKr99eOYy72YGaXQUBKOIwB4qbsF5CA/rFiyxmExdHRb2CW2Q
3NZETIamLWqMnjr1+7jWZjgfuxSJOkDzIUutjPfOQ9wbTuJd2mL865GdHYJLV2D1
LDFwa3QxpwMoCM4iirhKhNvhQ0z8n3RPx8/qzqsqkNhhGnqa9Gu/Nsk2NUjWmdC4
xEVtLHEGCEgvPR/Y8eM1bhwWbo6K3url35Drb+T0KM/0ONtOXrPxbASdjy2elDtK
PMyilUsB8ASMaJJrc37ag2OcEeDElDD4jqARbv68nT34CdyGgemET16wM7bemnDx
3loBEFdZnQ+ynX4lI7/gzw5fTInbHN4bdt402tDmioBMc6J1yXII1udKdko43BuV
QjV0ZrMftFMgNAYONUNwy1obnXLVxo1kF2s4XNWwoYIybrOJ1v6ErHfwC1/eg1+s
xAhSkMxdWnMRPuM2+W0zzykFt/qErZ4g1XPhCaCTxyZkCgM1fHVhAq/AS5/znHGM
/kK8lOJrhSZc1L1y6kiKbcSAgH3ARydRKI7to+i8N5qa2JGJDAhNKh+wvh0OIZwh
+w69bS//mqVEaIYTcsmdrm2zFl3HFvuXVGkrH3M6WfRnVPS1B7GMUhZ0xcOWfNeB
rRthGqJq4BmTy+NjeIO6vmFdTms3QMxKFrC2eetJh40ylyj6AirPhdgh8ChfZGmt
hqnNjKNRfGuwaLbizvkzxmSaW0VGOEwsVyjltrVBGxTHGUEVqsj1lj4bHDsZ9T3Z
+o5GN0duCTu97/H1Yg6nCo4eKHoqibeQSmd1UzJKaX2Z7qPG8+3Nt5P7UNKfsLOT
gjkJsXUe+KfepJf4xUEYaA==
`protect end_protected
