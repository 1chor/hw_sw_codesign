-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tp2eHzniOFK/ZM61u9nqtV1pUr04YHTs3boc9gPnHfqvBR25Lm4FcIyX29sliEjQ
fPQQ3CNFECn62CO8ABKagAkCNhslCtC8YUlJrbtF4wTxIJLfSNMQTvCeq6gSwyz7
IrtoKws6sg4YCG+L2SkxVC9EZ8SacrhbbgUv2zBmKXg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 11632)
`protect data_block
tMkn8Y0YwdUYfueu5xWrD1YsPh3HpPrUFNnRbLgiAwvWL7j5r30Xrk0wfBG5kdEe
FKVxZSxO6Qbc5hXijM08a62EzGBgJ9WRBW3Sx2fzEJHlg1SbJ9OqkeItZm+QZrpf
Yi4MvH9+kXHTDXPbIyr8dH7m95P2PoGJy54psT5iG44luCcaZcR+ZYceEZEvCTAr
XKrf9hqyfkp6yP25088iXhzZTFKbcbsdARy5WHmxf37rXLuSr4hBO/bSqFkWcwqO
b36s8gdyGyxiVc8wvWcIRdOAFFkHqeHfeMKOTiblm1zIaQISCKXbx5Og+tWX786u
Qt32EVOqDSo7wG56nJ2DuxxykVw47Wf+VPZr/dS7AZvr7ksGc3/H+1Mc61dNCxgj
E6VslEvoO38pWndOQjdN1ITkt6NPRqviW8rcXECyGtqq/IyB3BN5OUXMDAbUFEzl
poZ5AJ8Z5Xe1YoOb8EnLS0/y2lpErqaUVa2++LSMLDxeRivUx2WaqJ3/Q3uwmojh
NuT/TRjtn26dR19AUPtaSB8hgHRsVb/R7pW5hWyoHGe6fgJOVXR51xW3c1hvImNB
5+SI2g+wIQqtcXV9Pr/XvBygmfmGiIdpLtJ/sK9+eZC3lJ/9l0Qfo+aIebqlETRn
/KnKFttyxOz+iPRXCbeGvD/5n3zUZ/5J5zdNA5USen/tH/uZSUTnNdA/QR3LRqRW
5fljp/FXDzV4jqPGEbiNDkuBCWLvDo+qSbxw89/ZRwT/VPkoXnb+PdwkG2RoEQLH
XNLV0maIOTeoQA2XwK+6ASCn3jvdIIabMPTV88+pMZFw9mMNtt0uO1IXcrCa5ega
zjMRl4XUxJ11yZG1xN0kGX4m+2FipkJ9NLPaixRyK7pdHnDiNvHyhytp3YNUPhaL
XRD5+iNsczJPVNdZDNoJUMRqFML647I8A0Ujx8mKI0IlLJFnEMVwaaNBZhNH76Dg
KIRAUUwqC8dMJX1n32sX2OZhe0T7bz3bmh+TtIU5RJL/C4sUSWMhsmkoykwhFrfj
1Zcl2S0JOgWXP5ln8lPMQ3HsxKDAF/Bd+VxcXSqTtLGThE0nVdA8irjegV/SmL3y
1B3eC6xDvO8zyj5/xKW/t9zKG5RYUsyDs8KBLO5ryU+D0BlcO0C3FdYN9pO9CWui
dfcKt3MZeNHivlnCZOQ28QfnS/Sio0KW3TAlWYLBjocQSwgkCy+whmYP5KP+YA9S
C0vERrnsfAA+ztTsU/2vvI7iCp8fRCyeozgR5k/rwSHxvVej8vyO9aofdDm+EiJL
nf4h1mHf8uy0sXRcOF9KUzLC6nX87f8/3Ee+V56mTBcPfXR19QQbfZWNFNSP1oF+
chGKyfu5URjCJVOBGIr3yl9Li95ByoeTsteU+NkYyWNpo0onBBotI42fJppk2cFp
FV7D53HJ7Rh9kyjguHPPfNnXfO/W0eNPGjcpepx1m3rxkGHLkgygW4KLQghPZvwn
C1h4zqNX5Ws8GWo8UgUhH6XScs9uvmAkX9siwnVE3e5Hz7ftIeBr+tH6DV1a12tk
ivP8P5CQ8BTlNjL4zB9B2JqQStV0QvV05JIpdWzguzJTEO/42fqIMmbmzKzH6DXM
jMnid0kvjapmidS3nawRF/g5uzt6BiCyVUIaoTQO7Zqtarajo214eGw9ecHYyDzx
88ajL5stpiasl89chW2zquf6TL8yEYnYI7h18twAkhF26ua5EOWZ6E65H5GcxTka
BOafblnsqz8HSHuLdLN8nGB40tvY0TGUj9BoRcQk36cNP02LiYbGKidOqXsXpGp8
jfq3UTNWn8RZb7oeVCev1sqkR8JgzUTlLnPV4H6Z9HvCNqHmKZmh3K2Shp8ty08/
mwlff8Db60ePEvWqE2Sdv36+VNYah1ut+cnyA8HgG6l6BxjGXSU8SM1zWLm+a4Nt
aCFPNYGkIPIJWs0OyCIvv5Go2MjPVyuM9I9c2bdJIyy0A4MwBNA/b4PopdW8WeJj
znpdbOPCmVYzDqh3kkbBwCRTn50eiQ8uL/T+aXSicWmiQ7OTVM8ydT/CyWCEOoYS
hl4Njlgsv4ILJspLMpKCwtkG8O1P7C3bEA+uimJ5OIqgbBLTPJ4lzgZSSgrPOQy7
t3uHl4xCbHJTKYrUDtqTe8NZSN8S6PZhPyRfwH/QFxGBJPC23EmMKUpw3QX3nGDj
inWbETK/5GDsOd0fxizP+WF0w5wx8wl+nzoAt7nLPd4fOrxJ9GpyJuZDGiQf/M+b
yS8LvECdzH0Uhyf1wbMZKvYtB2jipT3LAmCGqzlRT5Qm1js6yKOaWRHcpT82nxJO
eOoIqMc2aNElNyvUHdDAdslgHTmG40aSilDtryzI4s7xMbFTeKuVNX4MoTOjuDuh
WuHYMU0LaXXWwju3N2XaXPhUXZM3ID7K1Xd1PGyHmhw6KnkcwMSDGVoPl9bv92oX
T5NKEOoMLYMF7p91QDTIBN6UJwooQ1LBalSLNcjlAEAolnsMbRE3kEljOb7PJhtz
YfHGyzwzaOr9lGnPEdL/7IALmoP93U0E/hC7EFzKf+lafn+BNonxO0Ao1Cy+nkWK
D4klODu9RUCsj9K3HzhvpVGRA7DRgX0sr29Fugjz5witxwDhSBgeaA/bvWQAWdf+
b3uA6neiwSXof8MlhTmFkytforBT5mZvBvOG7RM2OJaT1zTJ1V9gQ+HPg/PZ1H1g
FS3glffMOjvIl2SDzSCQS/RtGROAlV2KLS2wtG5IDID+i36YV7XSvvexafpphKm8
a1HdD70y32WIWtfB9Z3i2d2DpTB7VWJo/0HcjOCM6QxWbKznjJsh83IC2SnbT4VT
kyA7N+T9lA9RZhShsiRRFOvtFLA1UtmL3JunqiT+lL+Vm4LhQhM6Sho4cM2USgI3
NSGAYZ1DbweP+2wYPt+23M4T36RSsTA8hWVPg0diAKHEHETHugsTL7/BHSllKgqD
G8cLVGsX6X3Qoa8x1m5ga9yOdqM8aWhhI6Hhje0T7VBqVxQQKAyeB6Wc/aEWYI9J
XkVgrYgwffojYjPAc1I1AUn4B9rJxqoYs7CCBQzIDx5Mw3RQneV9f/Kzbcg7EHjy
5iy9to8mnimFwPnmBOED167ZdEYPyK/pf7y42fwjmCkPCwgFtFgrV8SKn9taGGGH
mIIKOTaAS+2ds5jO/vWkiAuhS5gYeJaPyR1v2FLPlfSVjpehVl2XMnTdVHOLOmZ3
ksIEpX80yHL2JwM14dvC9P4qyDB47wytZGxFSFlz9oAjZo+GYVMfWo8ONmx3EYqM
R7cJcjskQn4UPfKsS3XzbOjYksyF5WsmKF4H9IYNkRufG/diAqBQvE/dbL7wneVf
dc6IFeh2vPr8hEdXamg2yDg7Vnq5c0MN338hiprstmCQYhQpv6tM6o1xh4bS5VPB
Ma1k9EyBxVx5e2TP7aTCXvL5CvxNbWE+p3PaRJYPuF+h89DT97Npqr0IyBxmYqck
8xey+ibKRmyUCcLdyRI9cJK5mTrsygOs4mZt/5yh0SC2bEisOWqQzC8+ELf2kIwu
5SKMpMBwBXd4f0GZHHrM8kX/K+KCn4XNraL9/IGAz9ye/Fyh2kRIfYSg9PzlwRcT
fnjaf29Zxkvp8+C6cWWAa+9FQy9L3qMr0zMQ87yKzHnTbLd09mZCvHTb4HOTK3hp
WQYyce/H6xhkHfypUSnSVbRY1GpABO3CEDKErP3IH5Ieyo0k/UfiI7eCVsXrPYZ4
2lJRXfLuShUQNlwuobswZJGnICBjQETvK6mxmVY20G79SBguBxIKqt5D+AJ9KVkL
qUKQwfP9/rTgFz/zTvo6m+qNzHR9r+LQISPGbMwbHSosRVwEpDxjiuddJHl73t2M
deilX1Be7i7JoFnkFJHXS22YQzFmB+dWBVQDjRhwCIVa/nmwskB0BQnAwUoq9Ee3
a20oyQ87RJyc1Q74EWNYFBU1H6jci+6hwmveWJbg79Rdqgf7p4KZvmBOvzWcpyqn
9Vc7984QVYdOps5r5qPBvrTRXpfJFAB/wBVF8tBd0qLUOdLQK6xhHTpQanuTZmxv
b4+8YZX6eSXZH8ok9edMoigJhs/tlJzzOZDQgaZN3XjfXd4wRdZsubORxu8E8oLc
M2Vd0/N02NLXNviEgp+Fj0BunZG3AfJl8cyYViJdC/9RimYR75heWnbkMw2cG1FP
ABI1yIuhawfzKvYVrnK6OredlKIWxkRHJrdqunsjLWRJ1/wmalXOrHxm4wVBTVZz
F/01r3PSMIJHuLRJ0Mh5evZ+ed1DtrjxB8huNZXekbUG/5OHCXVMJYgqF39dIldV
YxBSb+7p4AsPjKwR4YGNV11fljIUE+sYDdaMRMdKXubKKzhtGnAwjhQ27JP8jCLD
uzfckPTOptoyWzYJ0kZyPyi90zP4uSsdnqseBBF7CbfqVw0aqfqCr/TWYBJpV+/P
z4pJvs5BS4GrIKySaWomH2uptSFzMzGlKXbFGI3ltC0WrkPMsDo2q89v9UGpTPt3
LzgRnPeIbm2CxDbprf7NtSIRnGAiRxDItQltz/TFPmUTNbOr1vPuWRKTK9XlVy32
I74cri8ULAZd/9/vLCdkv+sXinsjWK5KhBGSnv65kqGMQi32rnO4+tgNFiEGv7Tp
s/Ck1mako3kMTi7hKf1X/Y/s5vetE4CkdBueQZlWnL+sWjMn+MsiW9MJIpsP2VIu
s2oCYPbsz5mWwfUmBJttRmtfIluBC1xWYRZQzTFFtNmYupYpexA7/IfBINkyI7Hk
SldTkNFP45eoaflsGnVE1Q5i4dQwPG9tbUJLODwxuDCpO90rgP7JZifxEsIjvNkJ
R2z0cYQj5uZ/Do+R5HYsQNdqLQLLxaqTaylu34G444mfJBHp9pvd2CNVLSJtsrMW
xGRqT78dXO5pieqF9UGmPW+8IqHb/APBsBcI/9oCgGnWgqXFCXxAGoytO9Ial+wP
0aNwQr3/+6RHvDQHmu+O+yxZFO59tROmrJ+Ikr5GejAyD9HMhXrcYfnwMdV4T1RH
pXT5io23qrbs2JWdFl3whRTohvJHS7Wq8tPQ3yLxmSFcAttec2wx4aPYct9OVIWe
bm5rGhABBAL1maTr4immYQv8/dxcXMbKGWSZgx7iiRykimUen5vYYidx7gn04Qvc
r/W3YlNvarbvQASQKz9IgrY94fD7jJDgnbPfDCd9lkIvwsY1da4fHXZ8f9LQYPGT
qsruHunQbdknToKwF8/6ICCR77N5fWHp3Tqe4CNPBtXVLJ6MnO+8XVLkEFZXJKy0
9PKU/7neeyFtbhk3vFCCJxdmnZiuXvwVFfCvO1atNeYTMiz/hDbLNj1p+T8zAjRZ
YLA+tmyd6VpDA5qTc24STVevw0JKGRB7i8nBO6Ycx6mCxZQjY1fMGVxysGKZda3d
7SJo/f8cy3iLBtzDo47hARd4sXnwO7JJroKx+JF6OA/qWklPClxchdgmaIasqTKK
sftob2CQ8UxNyom+Mukf+hM1KbXZXo0QlXIR+B0EQ5PAEryKKF+1PtDOLImC133+
GsyOA2J12r+ddbXoU+AKx1gCCaMh5KVl86Y5hPr5o0rtxvt2p2ik1nN7nLO+2EmW
F5NsUm5GdF5C60fgf8mtZ+aMDMquEpu3/92+NPrwGj36crhTpNCE3wxHyAxRye48
sp1f3A84sxckcfwNvUkVvDzsJpKQv6l6glkWrXTDad+gOzR1MQMRHJjxdkcv2nG/
g0abBjNzUJSQe2NVWoR9/6/vDWjnfP1a2Lk7/QVzWZAlmzChk8ptHjBmUNudGxFZ
++ij1yerioKrBsM/HvQJSwfCYyT9wT2PqPqEs7rDxdmrjCG0iwNgcnOe8rPsFQPC
K8hZ/YmH0fxbTYULBcU02W6ZkVgQ24jgW1AlCg2xyWSsZ9aXsUb44mKIH8yGgg9g
D2M3rjQlGXxrsf4jOC7qzUtBDLUY81hQtvDOLGd84FyrBgOEFGpvJ13XOoo13xLy
WMGmR+M35VkQHF3ZQn5foXnOSTaJX7nzX52YaZYny2PQ14uI8wp0v4miwGbWni2y
MU4v0i3qVlmpX4Mk8lMtU4BRSvTerZFh2bmc8MWIW7/NOAnjHFlJBYrv/+hiZdx6
1dyVIeK3ZOmL47MTQryWkHRwE0Bl3j+DekrjRtV/yFILW4A9HScrpND6NZVQSryX
R5c5uvQZpX5sq2YFojnG+xdfwp5oMHxvM0WerkBr+dyKv3zWkmN9D/feTSS13gRu
uWR9nwGGoEloUuNHPckZQiK+HYZtjZTDY0WCde2+4faxkhQJ9n9ER1KjMTNwrNxx
BVo70GQhixdhma+9QQEWyMnLVUQ3xnLZox1JrozQuT6IUOXJbgNEabxiQzs9KJY/
/Sp0gqqdFUqWq6Kjwjvo6PJ8ceW9oxnEUFcnaEjeDA4WjWsRreUfN+vFtvUVUb+b
I6R6nkVO74SK+sqhoOtJkAYOVpAz65NOjtSYVGRRAYgZ5Rd5/dYMiMIFBbqhnAu5
QD4crPqTTc7kDva5kcd+ODqN71w9iHQ/dJxuFB/Wm61zv4QjOfWIE4R2+vJ3IdXR
ZF4aAtBxMiXGvrg0O2RBNLkz068r8yPxN7wTW1L8uGcr+NMB82QMmy2AOn4dniYV
d7xMLLjlhpn/toR81tp5kTffrTpKDKu98AP5G7pkBEtdyjeOq6nDOIaa30sj9nL6
fhJV5ly8EVNKKXmqOfecyHsPf5V0JR+ETgAcffr136WayXqq2jxft/6vO6qF/b+7
9h0rd2sG8iTpDrocqajZW4mh0Ej9DSp8/elFP4he+7dYYasq64KTPl7i51C3xBaX
kLRnk87c9xuxNzDIdZGdKzUmVlZ8aBap4kGQVU4lVs47aN+QG8UtrNQZcrUvg0Nk
szVqvENaFwIcCjpOkUq5SKUGr/KRCXslnTtzwhN4zPmNpsDcS7wlXUF12Eu2VEVV
e3zfLN2MfOsgi5jUkP1DgzAlvtZ0ZnA80lThjyyF9b/aYkVfS+MyfGxQ/F6KAHuZ
GgHqFHGPIsY6g2+MDrCcbpz13aOMRwNFNqWVlQlGC11roT5Cd8EBsH3RE3REI2jU
nBSk2p+Q78qOsLKlXYPij6jxfa1V1nTdREJBV+lwgq4vTW8kIakvoVS+PmQwviQi
0bXqO6RONA39Ytb2hNcjD+v4FCJguEq63Mn22akBKtAGWkf2muBZWwgH8F4MVohu
fX4EvyAFj2poZJwET2f9gjjpt3TQ8lt8TiXMkdbeGgnBsi9ziMF4H++rDj0BMD83
LALgyFQKySnQI7s4gRbj1ebF3RDAxqeAjo1bTW5YBpp9Mwj01sW+y5fClNp3kEBW
RZ/UE1ne0hhKZc3vYdjr5SOxUhbX4vU3jdJk+VMj4nMmLnScPEbegFcFtXH3M56U
rfjORV0c+BmXrcXOfNxswDhz2rGi7lO3jJtGFeCFYZj/F+qgUB/e4D/wnAly4TSG
mohyiYXd20Y+TQGOO1gShVEXZ73cSIJZv69XgR22RXT8A52Ar3gfoSDFL2QHEMBv
qitW7gFcGzRsexjMN28pLMEPmouxprU2tmJYD6fybbkjf3cetFGVggLnTIY/335E
qbk0D0anQx7e/zci3q/Dz19Tdgn4sm8iZEcqhE32znCQGRnQ+sXFyed21P7HSuuK
f2nLDt0YLtzLhTqx1lO5sO9mgD0IGDbCUZtYLEApcxCtWH6pKpJvmodX0swO8fJE
kj3G/uTqa9ucn4UJAgqzOAJSNHwetdm1XacVmYBl3cUJMESvzfNPAUPM2+dyLS7J
LL9h3DyDzkrWCNORJGp6jqAbtEpKevEBm5zUzUWs1ec28GgTHRWG+LObTncpta23
Q012Lrn8cTgmYs0P+lXH2C1dFUjiZ0j/6o51Q85gmk6xRPO2L3EaGkNENknwZ/PT
x87b5qctFjRyDBe4Oma6b5yq8mRO5+sG/A92d2xVZ/9iI/9OkLis6wD2g5SkOAJB
mJ2l3V/0oltFlOZZpel9CWbxM7CvtX+PxvVmnqALKUet+Nm2lv57SaDlTY7teW8e
S2QlB9kOcUHxf/ecQz4jbGGWZdaj5TW/g9FtfEtW+xV7aAaPtyHmizI7crOr72LP
pDTNUI5VEgHPNSptLqSQWagMivesG/DsTVMh8ou4vEqHLyZm17HHZckcQg5eGMnQ
vOHLY7KkZM3zJApqNWUj5//3Km9ZYBy+O1hP7WlPNcZ+iRGmQsCNcICasvAtK2Jz
6nIRr+8dF6Ziygi2I2aqCkDea/Ruw8EzJESgkNkfZKIMUDdTuf0wWlA6bqEybRL9
rHMUbjJQSpPUcxbs1UuB/0UScDF/63YL87GJcAqeqSVrvVzHaXA6GsatSjlhUHOL
YofKJuaPAkitiFpqr/DezdEGuephiF+9Lf4UZRZpoWg/g0Zlt8v/DuC/KnaRh6lc
dptT2ov/qEx3t3HiKNZhK3PYvwcJQ9igACZ2DOtLaCYlCXxtMGspYmB9BRsA4HYH
uJb9S0XW0e3np5u+P7g4jjqO5JRN7RLcSHyoQfOQ5BiN9AIgI5vQtB6wtFfJvX9Q
fG2mJBB067QQdmIoc8iHlmi6iXmIPATb/U44wlxRPf2gQMaSJ1kGuCm61AnLSl8z
ljFULBlCrppJJlduPr8CuLODjAVk1cT7PlbNQlL/Xv/hZ3XZX4860VZHpIqXaUBk
Y3a7VdC1q3h9yAn0+rwQ0+A+GfVGidkLgxmR2RQBUjQVTZWJHBazlPwY3jl2qyki
wzlv9RbJaW6QpB7RTzLYyJ0Htgcuhq8Wu1h5anKNQSFggpqrxqpV/8XGMbDMoOt7
hTni1NDbwxlvSUdgr8zpbvhgipgMEj7a+EmUxM0841ECZYXZ2RIFbTHtmfYL/q07
nFQsrh6LshiYpsIgRKTlCcBFh4rw3Ex+llZpJSSZ0yEspO8pBsffKTHqWHafMfY5
m1aK+pUS7lW1wULv2X5/Aw5dXc8CYM0BYuqE6BeM5wCYSPmrOtZyyjPNLiY9R9Yv
OyTOtzbevWB8yPAZCiavxgnouw3VDHkqtbzFsrW+F4Gxpv3gpY4GUUhIfau95xU8
ROZBgyUfLQpFWCl2hdT9KBCSP/RACy1E1AAcajg5gKAKiMeWNd6iMVZ28Q3TlfFa
k1Ux1S9fdKmMraXAE18eF/T8StKC/RpSRxiqG+t2DFrrmBTZre49yG/90J/H+5qz
cMqzXaXWeQb++VpOzlvkRAbGiN4/Rw8/Ebc94t+9SbFT+xNop42x9qVsg5qZxMNK
SetKOFsN6xUTVmqTBpKl6YmN/imTQoyZCEGg+CeGZENekw1wwWKx1hO0y1IOy6Fi
Sd9+5me8u28/iNS6eD0tto17bnShXAnDKK9Kk8We3dZX0WyRuh9E3VuMY8dtWKyE
oCBhARYWrG1a3sJAnS671BtiksTEPla05EDBSQ0jbasYST/Ok1qEM7zxG/GSEi4q
Pnh+480PpuJ7GNY8w+ct+bIQjV5lO1D7YMtd8R+eQMvFBZehQopAG63xTAqExiJa
hbqYQaB6IUp4BnPvQQeS1bjpJBmTOHv/faf3nFepqaG6jBjOJc3CIHygE3fVOkit
sby+k098DISKpjWnnNCjJbq526QNNOYtYb/vYpQacZ94Tyc75PRyMIl4soDi2IpN
3XWZcaIH019AL9h+DK2rqeKouSb3AZtCDPGPZ5Zj/FvkHz64KP2gdAFvib0LwXAW
FhTo9NNT80Wl09tgt5cheJYe8hiN0TGEgnq3Nji0v6Bj+X/BFFeNaOGlfpSwhmJ3
uu3GtR3OR6JPl1l0yK2Kw0+R7lZkZD3W2bo5HGPx41IL3FseOtnsRSolBU4XdXdL
B/FINMIfE75gSa/wWhm67QVdoLFXlg7Tcvp0rLR288MxT/QhgpPs/L6+jwKTB1zv
nmKybwDLBoOhUun3IUdxfYc+wTRLfTXvX0tkx9BlU7ikLMiOMPiDgwKvPHj7tYXo
/lyLH80iPZhSaULn1LZEuAmp1/XY2WdXFdvT2Q+SIkw3vYRkLkNwl00+LQYt5AtU
niAopF4lGaJ60f/CQHhK+wWl8bDy4w7BMTzzgq/EyUr94GYTnAw21tsxrFnYmUMN
8Fn6k5XzMIyow3r5eiEEini2ZmwkIBa2qub7X6sSEtBO/o6PjtRZpM9dRM00Jyr1
aTFeePpQ7kBrm10c3HstG2Kphoa13ivUlMhBsad8q4nRwSyysBJ1q5HjCzakKoFt
Zw7o380zPfFHSrO4bfUISepzQ1i7OMSeMZviKvHtgSwfld//rhWIKo1D4n86N/AW
jktgWwJEdeSQBCxt3P1beVM/TKuhXYyMZs7Te1UpSHjMr9pHGXsTvGl47Cbx4xb1
FvU5LIndLd3ZUPBuhHdTyjzUnM885LlS4S2gqYy1wa/GhIn+HSuo/X7/df+1j2ZF
l8PrgiiSeUpWBDQZu54Ww/7yXxqpBdyB9XcCrVvoDgz2tc7ZZKpLTDezRcKJ6N9Z
MdtAR/j3sQ1RMzh9h7Ucw7/RAesQs2btKIWMUOZJlOGneDD5ItjJn2aPDPbpwvSk
uSNIPG9AgrwWcTKYUdnxqsCCOy7aIv0NHLuXD2wiyv/taCO6FdqP/PlwwtEYfIem
laVZylHXDXd8YLqdAUc8+rAWI+luI+ha64jvzEQCcKWf/qumbWlHURAgGs7vpROB
8Bn5TyfzXxKMoGVhNb6MGk6ORcVE4LFUnPZy+Z7FcIGjagpKFvi4luKvLCAOJq3o
vr/dNHV4uF1VKYsefSbSt0mYpZ65YJ0YalKn8ybH69ue/T+grBovknLtpP8efKjx
rHGNo4tBlIdddxfz0DMc2kJCHIYHCE5D/ocJxN8bbamUst5UJwW5K7FeTjDsp7MJ
HIqcZHIctCP3F6buiL8lWPjNVWyqdlKLLgFa1mh+lC5nCD7up/qovyncgV/UIJtp
90u0MDI9j7J+QJeoGevMw40JfN+/SefyyfQbROArSWxgWpLYMUxC0LAuSoWf/KoN
xEvaM8fGTnipNrye2IP9uX0DY5LSaP+GHj7hUBQn/4vJLNUzwx7RV5ZMZ0UgnjXo
PTxo93fVzEfSMirHtfbN7XMLxlWLbYSN57WZ0AZ9bTLELf1ea3C2MuYQWCGvxeI7
FPF2bbuYAy5HEcqkJVHHXFisHDX8dwzdM1S2rF8VZVYaNcls5vP1hb9Ovb1GgDu/
yVCEfvXrbVRzmfO8eE2U6ehbrt2OTYy3ee1yn7QUK+auIbBq/jJwNnZvBMM7jFwf
pMNsOEJb4emQoZmfY0b7gUNc5yLZ77IAnIW+amDay3B754FXz+HzB8WprIpWc/aH
26JNijAJBaNM+UTiaAH+dCgjRs/yXRNKo/ErNUy7YeL0fCd1elHyb68jyQtdXuSr
WZyaxkz6RQ1mFbcEr/30zqbate/6DO+H9a+q3YyLfOO6F5vMRJYUG0qu9KMfPYQe
cV7+bxouZ/s5vAd9FQgu6Bztm3AoT/vkhUOYDsEgBTruIgYqfMuYTtLfDRgwCTih
KXM7Ujf0+T4sJUdcwJIxp2vZ9sFKcN3yS+NvLqGMDiSZ9b/wJJNQS3IRqiKyDESq
Qde3H1PMzkd0IRzqZ7f/ev5DLTedXADAb5KXCAxb7Gf+yvXNQ6M0HqAX4BQa0TJ7
GiE6jyTlxvSo32t+fSFqMkM5HiSA/PH5qEYujX51vnCxR/ggwFlaeTKVvB+m4Mkq
akyuMXJF4crR+Zp4k1ibjOoeq/W032AE5peM9MqYYLd3DexVKOkqVQe1dEiKPXYJ
a6p0aALrKghaZBbcUF1e60AyUG3GimJVAe+ZSQGWUInZc5E4o3M9DlUA9C68FRV4
92YMKGUG6p3L7F/Ubl9wN1oL2RqqPQvSazF5/zHRQHaRMUEG+k53R/O/Yvn/fHVo
qrbduq6aQFBuAXLjIUiOr/Ts8w5gJLpUUyPYPfuUR8ATvx1aoXufuZO04UQ2SiWh
mP+1cF2MjpL1cwWGUtcwP6TBoZyzOknq/6p+7q2bW493k9XeBnNoI+zCoeL50DF/
KSc+V+ZqVM3/mzEstLiIUV+1V5M9Aa34dIkRCuszQSKaa6iRmbxJtsko+XX77KoP
jf1NuRXOaJ6qyX5dRqsQg0lVRAJpqSytv1N9GO/U/EZcJQJCHqOP9hmw2tcJUJaN
ILzQEuxikU9jerTXjmJ0Xpsr0uN6o6VGgBVkO/tCT6IPlfnzdznM/YEedXyevXY7
QxMvISfQtJ8ol5tB22LPHaT3AbLyBn4hlozxYUdwDn4oP8PyMvRXAFitjyTiDDVW
+gVsK5VauLTwd5RfnQLoiysSMoy9UU5EXJEHo+ty+Vl4IRa1Bt9hTjbad/Vrq7fP
5RBUh/EDjfSsNFwese5ywWaKqKRaeKN28ZxUL0TJx7595emDJ+396fFcQwo4MlYp
V8j7h/8L9Pw0VkQqst3c9UJzKOgpqP9lsa1s/fUQYqNyT3kw/SlFMXLaaWx7xSZb
BNZpXfLr3bfqQ/hKaOgrSLE/t84kCHcHur4ap1NYAgekEU4oy9mlz3Ev86719qmz
vu6a8UKFyV1gN6hn20P9jLZPuWtTJPjziuhuLgZXQejl4TylrDC8TF4ckV1viM9M
usFpJvnmfm723zGmSbN9u0uzAcMA5Ag4AlMjDvIvcCXNj2Lb1I/sbg8h2Bquzaf7
ndj3gE8bsH4sfAMfPqOcV1tKtIUf4abEbNrON8o+RfFcJ1ulbM44etpaIzpKcu0G
q92W+7LBb6Ri9e3BITB+UPW6lKtNMz77wxrcPqQCS0WMA/xInuYIlEbGHi7X7NOl
6jedWThEk0aRtSNQPbYZoAEsJRIdQG89uDXnqlJR8PkN91gf59140TaQAQxKHaYd
9ilMytkae3Lxf5P0P7tS8ubdFkTZgkYJGX/rbvCbneFlY7M/atPGl/etDjffWErU
Wv29yCxs59HkTz5ArMYAMbryou7uePoSPuHhnVsy2aF4qwEVlcfNR0Z7rf+b+yi5
SF5eBcYy14bWPePzKFe/auF3xZMVX4Jwjq8KsWKA8r/F+esNz9DCD47aj1WLWLpU
468Ail5+2eoi6+P1O9wiRINUDbL4/t0IL0brtCFkkyJmrgC3aVw5WqBRXKmMdtac
bA0N1yEucnSb1qZHTy1uKB71Gkegc/H6Au31TZ3Jg/qTZu8VrjMUg3wF9F7njfup
kLssR5S2QLwvX5iXG56+kYiBGBiHamB9lI2m13QoBXMyxWNaCcZe/0bhAskYH8wI
G/k67HFZxT9nIF7qZ2KPDpYt64WvmYvno98u/8YqcBC4OY18XnjZyW0tRGam6PNi
J1f2ZW8MsvMXe8CQ5+eotqMkYPnJoktMI3D9zLEaCAKKPmSrV+2uYDg8Fps5u1R0
dwuOUCSeBfAYjmfYzPhoy7RaYTWqLTgU4aP+lJxRh6HlaFXNaJd3XN8ydBgPk1mM
9cG/ubK0dbIr+Dsc1E0sVsoikkQlNRxc3xf523YsbG9FKHleDgYdff+XzUUPMpjE
9xFCbbzG+GYQrHqNFDNgtzr8lPcPj+udsleN3wt8PCR+MuMqZRCnexOclV0NiKZy
5SZJYUlfMtQI6cyncOu90/lzP33Lfbn4R2No7Jg6eDg+wK1pijkJzdxmr69ARrb4
yH1FqqrbJ18tWc1fa7b4NbrCAQLkeF9v8Rn4BuMKpx9dYHgEQNx3rfCVBVt8rgbK
z0uiEcv0lngBmPTksC2KcPZuSy1U2MPkMzUILQlYNWTiH0zQ8JZqBY289RanVA3n
WidH+IgxmQ1ehs2/2wXvLVx2MO96uBWgAGIjY7G5g4SD4r7XynUhTX2xvUwxXchG
0to/TrOHLttKlzo9L/pjm/mDNkt+nkjfFVFE3xfLM0ZtiG5v+l6XDLwHnFueWm9G
/xPMs+uBZK5HRFJDZglObVhNwuwIJVsAq7sI8SVEMqrGS/SW+g5+UKb9da2hiD6K
SS2cYCGJARLThCmgHMZ0CWv/u9MxyhkoHOt8ORc9NVZpujIJH1LjTqyek5W4RI25
hUF/P/zboiwtVMTZJ+sXZDabr4MmKndFgg1NMqAxt53ko6Z2n6Ue5Izf7bHyB6CR
GDgMU+Bz9E2AJ79qfPg5FddKX7497jhO/pNJW2KwkYrF4uP44pOtkVD7VJXubOup
X8XLjC+TfQe99LyDXiTtIko7mvmHtwXa9belKos6JM+/XA8r3XVPH1V/ndbRoa55
G9Zn8+PLBMNj2Cqpvi0DxS7WhKT3wTbuUQr8ecMZCI3HJFYqG09pXTL3vKZw8Yxp
hlIY64MWbfRas7EQdLdCeWtaOn6naqc3v8jxpIlsLtXVClVBDg3+RYCMbaUJQHoV
G7FonR91+t8/YjMheok/NW+nFBAyQHH/PDxrBEJPl+BdSlqzqVHQ1aUfe4MRUFSa
x2QBRQItPAUZvAnpazNYe82Gtt1qAhK+eMNmqHSr/btn5gAXw44yKpaF25PH+/Yk
Q8X1J9Ci7HgTxGgh7hmN+6ZyTp+sa3dHTUXx0RqEepPcVxzENcN43BZ3vFyCN+2j
6oJ1w/0VNDU3bSjSSMifTy17S4nB+f8I9TlCbLJ9YRciALw0/03m0W+UgDnnnOyv
P6u5Qfc1WqSn/VlKhW1YU2sTWK81SrE+gkpW062+fPLgoj0AukegPiMFmTVhG44r
ih9MqyiD99i8bn50WfmHJdCLygACSkV3XC/bJ1TEvMSYqfugu4FbWWfdCqa2nCnN
feH3DmqRuTUyW+wt4QApka1gW2KQqyA0+nVosip7ZlTeMLGvhHiJE8ejQvZoZuij
3dY8zzpO0vW0+0XzREmV8zqgcUQ+3yzeLK03b9BQwm0NDzmzbHROIIMSVsxKH6aL
8s24n6sSb1iqkQXaubWGaRhSgzpfM6qGQh6VUpqk5TC6hAcGsHJlt3lcCMLH2o6u
fEMPu38FG8rN4sDybs7DrKz/h2vRsWkaVPhugcsc+LDUsg0C4ro0juSpObSSLEJg
4MvUYRtUKYHOJVvQwAD8/uOWYzCEMheW4aULbz+XSdJ8tKqx3lnhVqa/eZozm2lV
ItducaI+5YW835gYUiMZ2YKZVXq+8nUudDR26pDlcf6S95YH87HUaIQ02eK+Nme6
5HB2Lm0ChxFEypkwmHLb85/Sh0J6MJqbI6eOXr1VbOfy83XMH0WeGZRNh0quUngp
qhLr3Cy5E0qaiR1L2dJeLzhi+pkuBUBrEidz1aOVklwmr5N3l+2fupSFSBr2choq
yw+UfRmcSZ35L0oQC7B2v/ViIMgC/yDMgTQv8JaaBF742UliJTjaIdcyGc1IPNQZ
EctXgZLzTu2kSBeodIAdj8SRCVk4bFpdpf4W8dp3p8FgW6+2yDVArKGqEqQXFSPQ
d5xiOawtUNutBBps0nWBEt2VCLDJN5mwekqJOFg00pHWXaLAA9/7ezAF/mUzS0fq
sXqJZG0kl/1d2nzSifU10NWC3H9xYw7ULrHb2iRbUHJzx99werNeql7tZKWkniWp
euw12An535PbJV3Df6RTDl4oIILhIlHI1nhc+T6DFCf8mNsvlCQiYzxJoFK4JyeF
ASkR16gOGQGzODrEpm6AmA==
`protect end_protected
