-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
V/DdSQQFumZ+kNaEOmHqDx1fCiV2dv1KlNPSLb7wHYm6FaJFoQmdvADDDowMpU9r
bEVwgyXNT6oKsR5RY9/oBkdOWX3jxLqbuhNl2Dydw3JqeDaFMKe5MwdXI3Jhhg8a
9oBRCxnoREv6JupiOFSp6+JOuBfcidLg4al7HN2ECkU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9217)

`protect DATA_BLOCK
9uFTd9ujokuo1hh6aD0EXRmYEM215st4Z1mWWAKu0WKdrMmU2cskwVXazce3QF1C
Q5T+Hoi3m4D3CRJSRm2jqj3ODpl5ky0p0aweGgF3QBAECtWsNsIvxpLlr1x8dVGI
p0fDoGdik5WfYQf9cbaPvcoI0wBdLesLMbGcEVh5CZVwKbaxc6ZnZkOi8wfbaD6V
ftKRosUEiA0BhcWPMlmreboJoXL1qh/N6sXP3l5r651ekgWwuxLlRkVIMWOUqP2C
Tq8jIPqBy1r8R2uFwbXEZpUu6/4CfTeNZqkq/RsYuawbPEbBAbbZRC4++7s9GDb3
tsKeh/HOwDUPzJ5SBjxmKc/j+FN4dQiz3v1yM7POXymI2+KKQttWC0acyOUNP2cw
F7SEb8HqEpAhLL+17wten+zURDB9U0iRWEO78nnUBUSknkpXLcB740wTJTN8K80O
IUzmAWkBTuMuNKWdc/UoPBqP6sXtsVju9KpqdLipzwaCH7KhVYkpS2wzpYKQbkSY
IIhuW+8es1lsrqKO1x2O6GfYzRzG1RgpUhHjXtuw5tMi7+Wcr3RRJYDnTEL+0BqM
sSwsR5WypTN7UzWZNVy0OKuCDhE8HeXhEtHRA0Lsyj1KmF/v4I+YlrRjpD9n2W4f
4p9vZ2vNLtw/fodXt4WKZfF1nd01xsNfLUxz1OD9pB9OUHMDcTDhu8i5VuKoTGGl
WAAv1RwqPCh4GtF/fbAsco8nGNiTJAGjTT1T8ahX5ZhkL3x4b/ZGjp5qqMhD4L+a
X6DpMPeyPwfn8IsJu8arVmPRDegHEl5S2PwswVX6XH+tUywcAx011Mmkbdq3qvTl
eLGHsdJ+83zi2ebZ4robzhipgJv3dU4fmJ33p0SZtiZck/890dD3e5WsO8SBZT6s
D8CW/CrTfa69MX198xUTTyvFAHGZ9vRyVFzCt2DhpEusMAhzwOvbNH1CR4PFFzBD
2jZTw/FLRLhYZX528XqcHYOvNhkqBkJloqYxh2ZJg6JEV2n7JpvCxgTz71bzVRZx
yKC90dbSIhLKt+KqgnrKHsDglJtxASL1hVi+htlnEzqK05SEFekQAFfzEUZ+DVWJ
AIBYIAC84hIi2ukvMnOqPdI/MPP5VIVgULAaJWCtbJ3NlD6EB9E8UR30WKh1sMuW
SWMC3PDD9Z8DSPSrrBTA1MKP/c/JT/dqpZK61Ix8cNBvtJnoFYIFAx6ST6dkRwpL
p/reHz5je+GgQXDQWGVat3G6vBz9aDFrqGQE2FbFxiS3HiN4HECQFK876AVTfH2F
mC0MPc1VpAZqLHDcH2jXvWaAwYq0bt/CIrUQLTkShx0FfDeAWTvELAH5dTcOWBv2
dUjD/xR1kpUPfZIYmuqSrb0B46vJyScvxcwr6JQwmsTogRHJcVBRepwDvtdcHZsr
WF/SXMZ1Ukm1vmnWB5HNIk2YEX3pQneEoQTnaQeuzW7CDi1nCqS9cyJAZSo3u7u9
Go7C0zr7CN8qfoHjTxy1DRBGW1UeNUgQCjXEmirWMOcVR9Xbx3Ply1M1fR9dTV2Z
LdG85d9BAal4hpR5WHzd/yAwVVExs8bKpPGPTHUKf6wk023FFtaF3RLOahppzYJs
u0gFv1aMHwe31Ew/68YCiNddGZYrKO03yvnwyVg25BrNENbBrsuE7/gWpyZZZ796
oju7sIztEQrCO31KgSzZg8YkDW5raE36wRmjH1avVZKo1aRQ2YDdWc5wTCsMebCs
08U7r4ytgdVpJ8o00CibiTjXw6BcM+Fx3OIsCZYseatfbcgW+o2q6/YELime13Gk
oAYzyrdfBHn3RqDqRocOzH6ANAOcOFx9VeGhdjDPf5Z1ANdeaSYia2ResahZvLHX
9rNjroHe/erEfNA30VSkCh44uxFww2kT6VGzMhKi2oKAkS2uyiv00jJacp4k6ZWE
bQHk33+TcP3B0vbv57jmf44J17XnE0EccFlZ/BG1F92yMXCvtqbQvHi1oJAstGFo
d7P4PA3G6tf1UQsJEQKiJxvpjnAip4qle4Gci0U0ZhO2L2ACraUq4/hmXcUx2bAv
kBkxjIvVdbyam6QKgQ0pn2umC0XTd0IqdQ3Fr4FynR8VP+XCCbRwhtiQ4DLtk+H3
EmUugG8q44VEAZ0WMMzcnb2F9XxlS8rPBau0x+HliVniFimL3qgsWbne+E1wVv1I
DQ4bM6qv8VKmtPHGIC+fzb0+Z5VEjNlqSFqhiRLm7AM/a063h9NV2kn3swIyfMdm
ZKrL51rAFMPG6VEYfZp0dZauhjF9u4GWYC4ZDMN2JlW1Klx9/gQ+HP46WlRZ1WyM
duY7/WDlUyBsieqa+LL3Pj6jBCASn9CAW+WP8Sr9qVCmS2ArdwJ7aOMT5C9+2ZOJ
uOBoFVQD1kp7RO0UOnEGWKSvKxkqEnGlF//SJk0Awm8alJK/BiMBBZCcfgr/N8w0
IR5K0qXlFBUZBiE8oKe7iZFKTaqSIVrK2dSNMPsJq2cr0p3c8gsqjHqbJrMqvJ3b
Rg1gzdKeXRt+wOj1ox69NAh8F5lm2q9mCsiRnqusc1dR3VCbX8aUkcM6PsZPyN1p
7+FKJRRg3IZAHqwDOET6kaNiMDWDVkkUSJGLSN9Y2FIuq2z5/ojiqdzLBmUFGTl4
YEMkdaaHGxcZ7hTyWROjAzswKnZh8qFBQs7a/TYr+G4DgKzr575xSjiEifSMtWdQ
sxyATotGjGrWxYBtTIzx2u+WkeyPsyOq8DVHxWWT3yaG2qqb1LIDxNkJjV7jMANG
J0lPqY6RkDgVa1MTV5TQf95WwcuMc5yKGbPrQkmUAdlRN/EP/Z2d8mGKp/uzIQUg
3EyrOSc1HRW/SK5F0Pe9iXQIUfy3YtEE7Zow3PP+/Ty7v2r2MC6Rp4FVlw9f7tRZ
RFhZ2Cw+eHfaJEwnd/OgeMc7Pf1uY+KPIcNqKHKEoazx6BmT2lIdiKcbu7BAXGZw
pDlRuL7KZKqWBRWCapI1AvE1bwLfrq+rHyzNXESyGwgdd6JcnLlVW/Y1Fet8M/ZN
h4AsSjiT3GddxGsoW8IQnuJOdnHornLrgEu3AeenqGuj1QuKQORtwcrOnUjmegqG
lSxNst5obYMki7Yk0oNrZBWpu3FJknPnxNhjvOGNnQ/PQTCuLRYfSvkINEs18u6q
3byVw9T39VaOz6AMLcUhAIkFA0ighYJVIraUY6B37gbBJEujHq7a9V3p4g1mKImG
jtV/0MlDbxhBcYv0Y365ar0ErDp2+3xk+NXydzu2+D7WjWtotLwuZbi5cxH2cIyB
Dlw/3J9ZZKalXzzT+oAYarjQIcf+A3GAY8l8Ww+8ebRnYvho4zxm1RX3xzkF/P1p
F0cWDg0gj6CGr4lgMtQsVxpyKc3bxEyROc93VSbh7xICK5NLtyyk/uW7rRzxLyG/
6tjqUYOG4Fy4aW9N/gdXKjqH0MdzTDkxbOVkblpGSCbkdrqUIk9g3B63ZKZbfVn5
qOm/phhH+PHpgDKMFZvLa2xKfDQWKKWEFk0OwtY9xw+zGouLEuz3ynsgV8GnAxyp
FJaXWQuaOoJwFcD/fD5oEoBOu2nQQ+LKnOPqhIvt3uctlXNFC4nX+wiv/CxdayM5
bO0dofCpmsT7eEnh42Xu4DlQZ95ymg44nw9LTVjfuhGuX4WcwAQHuBfqg5QWmdvg
Rp8DM/skl6jZrgMS/SiI9VQcRQm79K+TkRePd9XofZZt3JcSzEHCVuxhrWvT1Yhv
KddBZQ0ViChsqyyLJozCS4dhIeimyaPomzq3qBOTfVg8Aaa+g947H76oiUeb3t5b
J1RoMR9SHdnQiGUGAOWr0Zbee1kDM6SA6AYglaP65b7FKgU4y/vtw5BKLy6foPCY
BoclLlSDNjdvloGbhqnsanSV3Z0VpJpjS0QvcqHd7i1+bnua+2NRcQKWih+sI6wo
ujDKjbW1LCfQjLoeRo96/QCt1d0hJCuLWu/lQQx8zrplQQsAUExds1Nv71KSJ43k
k5KkUND0iZnq2/Ijo48nKQXjJ9FbYSCgINb4I+mwbwymr0bPk+2DAxu+MlKR+N6K
pxy0nx4v555hgwpJ0SJRDJLh2i1e3qyGpiv7KRySxKgUhh6MiSTjshQeH0q1wukA
vbE1kW81Mqyqh9LZ3DiGnWWL1UEPnkJ/YIhnsUMjx2VpXpNOl5DcB6pG97tIxfUH
nVTc2/wI7bhKp9u/Giiv3p4MakG/LOhDI9G5xulM0PqmKIcEdV47nGw07Vef2YZH
O5pUGbycyDjhII5hBGrW3DcWY8BFAAgqdXkAAGcqY4BaGwHrR+UhI/GRoB3rXMLM
9v7w+ImAe4s5zcaoJSYLPFg9YRoGXs1+wVuOjTdtpA1qmzQ8aJby3bcOuYKaD64n
kCZ0+Fj+fI1jhQtJEOlQmfP4EDI5UL4J+urGgTt+ev7eGPsCLwPx41wrvYETmtnZ
D1MqudQf/GbHwPqlRhComn+TooqME1dvQ7VZmR42ZmjaAR8oOAE6B1uARKIQYHhK
s39isIcOdWZ/Chddq1qCUhIGhNiBIm1oENA5IXBsIKqrFDBArz+iYSBI7KHvK3hq
AOCOlhXp3KZfPPKZuG3/taoYJTI0QEe9/dU14YMHfg+NEIxAETJ0PxXoE4FQ45To
X0ZHBLX0i9EpKjTgD4p7ypVo19B0EwS47qciNUm+cATgV6+kFRWfdtbXOz1gO2nT
MbPiXB2w3dwiXoZmKNGLiFbFOxUG+jQ11cxMWIyO0Hq0QQ4wg6+OtI3T8EpE7J0q
Lk4qeh+/lspHFj2tbnymE7zRp0N7Zi8ihXwuYRFj7cYZexBicBzmQmJSPLLkbCBa
U64hpGZgaTfUtwIIJjTuMXoNLVwUKWMtCaidJ8i0KT/9XQdLi2NBLVsNlVVfaEFM
qvj8m2lZjbR+b5i1ximFXSmmGIxC/7YhjgxT7G2ISsWuUGriBKbbP/RJCqDC8pFB
aOWe2K6mrgS/xFy6akX4k6oXxq8Ep1s5xuDHw/L8rG5SEL0vYjS+sKaswSMHxSCR
vNASecUmDwdr40YTQTfRu436EnNJK3LQLtXimAbkBJU8Nm4nQ0WEdKkE12glnImr
DU6OAe017KH94jdvBXv+5PJkrBgGFuqTTWff9ZBRhklCXqb402DHzRWGoxNLqEMQ
PzHjaSolmS0Msd0mxIc2eeDsbcg1fFpepCQCdChDjqXVHlE9A2rFpdfAKR8EtoxQ
88X8ffCWTmysPJAMt9P1AxULFPS8GCyIvId7NVS9vgKjXZ5qnxT7v27zmfnGhV3x
iovevTBi3pHeVHixhCZS4g/ThBrTCo8XhVT27mN4p9o405ehDnqRfSGeZZ7RjMhQ
hHzwViAxHy8pklqwef+hSLICJ/Es4pFjqr5tjs4j8o2oKT5/MI0jzeZrbrtDUlzC
j8PTMuy9BrROCrQB0ag+PNXLkyT6jRMA2eOzchSLVqQPWZ261h3kOcB2lKE/9DYP
AnEU2HHtYrJw8C2+xs94ZJCPYSx+PxMTQyQaSNIsxKPHNeFfTOK2ogi65YNk8aB0
VIRQ9CncTxPO3yTIZwWjR8gLDsH8g/HtejrBWpkT1E72FsDlH3qIKCxaBaS7F+MM
ZB5YwXH/YDiOPgobQHrSf8VrjmWywUp3cOQM6kxNEAUn/RY/GqAY0uy/4qrJaI8B
k1STs0ubUg3oc4+7gjl1AMC5Hs5g/Txc/M0wTyJ3lZvkyuAz4o04E9PPx+990kFD
5msUKN88Rg0hs6x1uDIlIrXfNOYdSrjwQKxBH2rJpbdttt7lhuLSqK+E+8Eu9shf
7W+Jk/eV7uDfy3WuTEE9HwzwKeq4r5LYWXOZQwufUBmzr0wHmQM1sop1qcB4YsCQ
KiXj1TJx0ljTuz3QaCFTV+sBmavbOY0Yx8xsyDiorDlFRCPm79Cqi/fp9/7qfaL6
Y3xzZ/TlvkTkOgMPCM8F1WoIjgn1Yr3kmqaS0eRdOXvoZKxwdy/KKYO3HlDmY9aG
5QHX9x5af4qLeZil6UNdrZe93dxDRkZpgtQYzbg//w/e5eVBfsP7pd6J4e8PTIKu
1DMU4dzJhhX5zJPAXm4RWItrZ4HUkl4XVRRvO9lJWrRVwbhFMTrkN8ydEmf23gLX
h7qhTqs3V9bgw+WUaiQV/b26ey06uH6875PLO6RHxQ3FJzZAcErRPUUho7Jw5giB
FRMSiEm76oQnZBZJas2Wbbn4GsX/u+UG1iKrw+R8LeUw0ne7t7GGr9+iUPUFz8P1
dBEHZnfAPgTacTbCvpVqIcQk7D2IylXnItQfcRJ6yFRL7MMUgHLxW1nRuN/bv19d
JK7OCB1mgxY4fVXbA7wJwc/+GvpEwUvtoGWD+K7EiKBhU0Fzw3GUxs3Wl8c1xruo
wYh5gOfhmxnPNrmFBI/JD7PHGOE1cEx0smbHsRwPQ9xvuti8JRMqAKlo41zflvoA
qDHKpomAfuMVE0d6YTrt4EiAY/1TPtRL2uOVM6pd7GMNPJxUqw5c0fj56aeGT11L
Hzbh9Vj9bk8EXlBVXSbr/RqjkDfmPIRwhN4CJok7nj7uBEgXzrkm/dwsCwGuOsdm
Y0fnEoIrIxvA5fF4Hb/Bsnj9EqS6JHuGO79o6aU4/wo/mUuk3WGxrUsaYMpyKyeu
lp8bPuUQZmMwc9yYs4yNx9Hu1LND41Pggm4xyo8m8RPnPVH2PAeqymJSGR69Ii1O
OKnW5TT5BmH9ohmjoM0cXMPgdG/ub9T57jvzQuq9lpA8wbgogBHaz3yMGxo4RkuR
y9z67AzuDOhoYeyzeJIIj7nT2j1jzozN4HQELlII3pN5ZamuTdUSsLRPNNLaqbYw
qPssaArH84b0kFML0UbvvKtLG5EKnuLjfw5bBczIyho9l4pLq2F2fTQvasEMwGsc
SWduhQZH0Ylp1/49myDZBzVODh+JADYHzqSCzeemS6t29+zL8iZagoBpMgvTo0Ar
V8Xs7UnNmIrEc4gutE08CZZI1uqf3PBl+PqEXMUiQOJOS8o++RytANAN6jmPuLFJ
/v7fd6CiP+W1hLJ3mZ86pw9KfUlNiOge3f2IjgECesnY4locWrZIG02XaoL1DpSt
XhVXuAaAzbTiyVZOdrART1ble6KjlNXiw8OAQb1P6x6Iyn6YveFZksBHay6m8WJ7
/ipycfKYoemLvYbeXFNe5n/GqrxfzLqRM4pthYUe4XEXvGk0ZIYIfT6Kn8wqXOXD
LeJPSOLgPJLsiOpIlxThlTEjOcifnpo+2x0gNKXtaEoTUDXHQeUAl8hbZlmCQD/Z
k5q3x60ERVteZ0uA1hIK3+oHOb/QK/1Za2ewBqhooxv5Q597sOUhN1W3Siy9NZwC
eOkuUwOZ9ZaBI6Jy655OiQf1nCsRHNLOsXrKyK6nBQlfnwW/taS3pquRTvR4wn33
v2ara4sDLNFeCcUSeDjpXRmQLk2d6u7AewGNCWyvckmHSZLc65pp09p5qMpe5jIo
SQbu+GAfN+P///8DtZ3ZeabsWobvUg5G3S3eW9UPPQ60/QTmU9AgID3EXb0xXBHO
KYseyJLzkxtRLTRzdn3/LWETroQM/rwojN6xJooSHRxB9fgiOps3SrD6PmylqBTv
0SdMSFKZdAKuIbp7VTUTG4ybnG5Nac6P7WSkJVtc0YEZBNbYmnVgbCSOYraKpA3K
tPgMpN7PhGH1Vw6rzBRN/IRkTqiywP+6YaCnOmm7YqfzmZkL543fkvb/nQ9dHGNu
nI7p3x3HCNUZ+Qtmh1GtVK8hUJ4ntoYVegDS85YZWtH/KQjUpKC+U/SiQYlg11iv
y84uM2+KYvETLNf3ZaB/PmPI8+OFrI3lLxh1OElwtWyHXIq/2euer29p0nx7vuAc
a8duDXMy7hY2b2GYky0EDtTnIAT9ti9pPRz/WmHW788Ovmqu4kU8OBPb4Ym/Enwg
QZi8hcQ+yk36sraroToQh7WvVxKXpFmBWSyZkDjGZ7iSgU2gN2neGSy6OjGvyS0O
puEuUjbda7UBoDA1ZjzjLMkmjOWbHdafOsc5Dyt15zBCYahhvnNxQGZHY/p2CEEU
xSo9AIKa2a6oCMd8O6+E2jkXuEMxHKIYzQFZuPmeneZQhvduO1HIvcPw9vpUDD0l
eSOr8qSudGJwfZ4tIso92ndmQHniBMAYO+RfkaE+YIZaPlUmhpDMoYLXdGAhE392
BxF6AxBs18KWkLYpA0gxUzZ1sN7l5LxuxfzRvKDOTyfat4+KvXGzzihu15SEBqzu
4XVftc4ctT6MS41tdyyf9aBAYAkr27nYN5rFMb0hvtcIIrFuCcQADYlPvWO90K/7
Df5ha0N+nIRl66N54F42T1MEnoiT1DbvBcGpwQkrgtIQaP+2wioj9/wZctA0xBBg
eNFZbpXwmDdXywC+4LYcmhh0GA+X5pxQ3K4eVOGrmGsG6BBdmHGEwHVGfvpWkocO
9166N+c1JtzLU3aojGDaEC86OvWMBrBVtpstq7mfOUmJfmVpbqDbQOlmlbyWahxI
MCghTuHL59clRBJt7PAjBXbFQQq4QqYTdO5rdK3JzqjIhd6fvYicNBZFojYij5rA
y11r+ZVRNYeQqzhrlf1qs/FfrXb9LxLVegOOFtWBXvdgPkYP9EstTQLp49IoKgiH
s/gEmeHQgv+dORlH1XcB38xs7Jf8YtwKvnR5b+BfIyn4Q5qQLJtzTbuCt5hmjBub
FJz78qkkRISqenKzYZvyCMPUZu+41TtYvjJMUVbz4Si3J8Df4FXJ9LsK1rmtrhuI
BsyGhUjsfK37BiEiTu6/MfE8tnBsk14hDV14DSDQ5naIMfIoGBYePVWUKdS8UgAL
TzN4i+WkzpfuW7UCRM9R9o+MA5atb63zNDn1R2q5lGDq+BmyeVvcMSIlBkE1fFcJ
63gQ6L4jrijsucbUUm0Itse1VzxTDdC+70iDQtOuXCUOki34QEX4UbMZoQUp+u1e
mChzYwDoiq5DuHYEF7TRIhPFxuKg/Z8flAffwL+c91kDjhh50CXC79uFWSGJ81Fn
Oi/wbLLPd32EIohum7Khz/D6ARjJCfjZiAim8jiUgZUOsisbVYrbWQXqv1TRlvZ6
qypTyvGldvQqrEUH34Kh0UmsVh5OxaMnLkUhw1uIH7cdjpOlSyNhVjasHlIzdqDH
ZKo5q4wH3olTGe3oiA0sG0dTMLnkeiNMLVviYFu5HVDozvlRyJbkI3YWwEya7gmI
odv8NbhF0m4Jq98Lqzh0qn0MIhxGUfiD8Xm2Rn8FRpFTmD+DztmrFZNWqeCyNX70
zo43crqK/pONFTTsG1D/w9ny/znDX6PhpQ8/j99pDEMOC2VSJwq2FQQ9zQipSeHG
Xsfyo/2TyqXzrQbhbNm2MrZrONqS1sOpY9eE1511i5KQvsywEeb5EF1KveHDV73P
AufJgfl46hGDs+hWgeFVa6d6bba00DysvMg8+cbIg/6AcaUR5Qvb6tnJGxsSDJut
XSANMQmFqKlB/ZOFlg2Y0A/GbMipRxXELMCO3cAIeCzHGVhmCo5Ejr+ZZrD2bV2R
M0jIchq4B/1T4YfYhk0M9LwCARF22BguqjBWREy+iScsV4Dsp51k/kZOBRBHEyv8
/CXXOY811FB42Hs2k5VZAVPl0tqSiPB1Map6aCXw3ZtCE1/kfsxdihSFOovGDQ/I
aDV1rSibPw6ig2bFF4txziCKMWzas4ZvABqAo1YZ0vqGiSNuEBJUUmQdPd2NRmr0
q2E+Re7hKx2aNrHpD5YvvxCrBcfhEbThdYEKhxG1TFWnb/7dc8CbPS9VB/3DjPc/
GF/AG7TmlwyhL9jQ/nC1iS9FD7S4B4f+RL1fpGMajsO2jY7Hzapf3AeiGT3x0KNN
4zcI4H4SAW+vaWrMhVrY55I9zQExfDvUgZmbntYorsNV3lRLr+aKJ5BqXJzMhGoj
9ZA5//O9JEaf6m0/ldk3dhVDi/8fID5CGc869jkZ0Lgs7i+HxMwLnz3iarg7NPUj
LHyILYdecm8IpUBncrKNG7Db+IrOldwnF5kS3+lKRDGTbR2QbaSQ/SFHoPdvBwE1
6jmbUnCdpw8pbOH+i6SPjsayNDK66zV99lh3DsVEy187zswaFom0fJH6CJBj7t7R
VyBw88l8bOsIP6zjYiAUNqDfL2yW38TffS12nwa9MFZJR9bDuEr2UVqpjKpp1Mrf
+okZp4TfIDTeQD8RkFiFLJ/Cja2gsgCtTaAnLqusMR8yqxNII4Z43bMT7jlMqL58
tPsHRm2xFcNCI/P50qSqvmo4aqXDAVjj3RS9FJQcnLCjwwO0v8k37M1BmKLGT5a2
SsATIoyiyYlraO/K70RpK4U/dzCKcYn49aDPac0W3JIjpdrjRAQx3dzKCMTWBA9L
wByMTVrFqiTfDEinjWt+g+/CNNHYUD4/ixiDjsZRsgmtQ7kXlVGjp04rBo0qfVZV
YdI5or1h64w/qZ5U9Z818OPKWOYClnz0dDQJdtKqPwS5Yyef6T9/dvT1uRb07hCg
3y+MpQTNKRpzQUdaMyX0LnD1zDsKWbO0VfkaRp4mKpy+KtT1jGPxyPxzRmuHrO7+
y87IV5/MVHS4j7PeFZa+ohhhuB+zcmLACPtHFd0ZS2f5sGuOzMJwFO2HhKiXXxc0
+znoJwrLbZ0zyiMqHMcTvgqFi5mg2Sq7M05YoTVUOjuM6x9G4S5qZaYd2RYB2iz6
hZp3cZTFL9Y9hPsRG4UaTEeHqES0E6aiGq0UayBugqDsQ999121+qLQg4ERkjp7j
ocTsKSKzoJVEvQXWEdMSB7uaDtOFj4nFhF3O+vEMcULphCyhOsmegxiBZ1FFZaUf
0AYkX68SBSi+9DjBPKelE1d7hn+pz61PIXUFzOkBEQ+k8IOJkPva1wnpwHLirn82
4e8sY+ULTORA+nofbVUTqszbZbkxSUJyyA609RCxIupgkmZfY75nu5wJ9S2XRdt7
/gCzf5qv+JPcx55DHo+Sg8TatOMTWDuF9prh5GNUg7wiEsbho48MzJr53vLsMBBN
kG8qEnewkYKKJ8Utq3jGe6cRM/OX+sOowaxg6fi1xHWIQ1ZrzkZbRX/dJ1kdE+HZ
WJznu6LWmed4SOC0TlRgP4bLWubP+xNM0hDKIVRbOu4neZzrNOn/DOLSZxByWcM1
Tp8niCx+4UfPDggjGZRUkcEvDrry8qjz0Z4BiD0Nn6LkKBo0LbyevMzauFCj0huJ
0XgNMkVIjHzZd4hFchnJek8OJbGjWr+ND1wbIO1zkRGa1RJizvcyyA/Vl4wFdHxk
I9k4Kg7ZTsmtFb4mgYj/Kqh46OeJQFRoEgAnOnQjKRwQ/OgBrARB/cnO5CcbRiEM
mV/zGYi1uZOI4IZ4iiZXpxyaT5d8PQm5lsaa+f7TYocpD47tO9xk3ObthWSOJ6Gs
IXZQk+2eHLnGA9v4pLQ5b5bbEV4P+SEbqTYwSD/PZrR5/PTxcBMQ5/ntOrRrmf44
6V/3S2jrHObAxfePuhm/wzul+P8PLoGeJweD1YaQan2KBoA/Z7xpTygmAbrqsI8U
esBWitypwhA8cHjK6V9VHAoS6gppwO6oECL/WeWl6/7rfSJIwrYMKGGHLZyZFepq
Lqf+mbIOY0UDyvOU2lLQhUvxzB1HZdeDmSZYUcH4nBWrANziKjdHc9PRO3mGQkO1
Y5Z3XUdfefjZ3dGofMwUcgwzIzN/IuckKl8IY11vm8LLH9iOznKtYf9/KZR6oYDg
Oz9ccMrvIBCPRCD6cn62Ol4i6fPQD1IIQBDjhWRrAOlTtjtVGNW+dcNWNAwWD6WT
j/Ynov+BGjTTQe/fragtBd78oHiHtdGan8rBrqgdeoy8PJADjfjF96THh8MQYSfK
yBW4VRHpJg7L5xsWOV76isPZTQIfJXUii7tpP3W0NmAOR8SQtDkxdJGYjRcsfGkG
xr19uG6TAYVXt4imxxHBbEcxtniLJWM5xTGn8OA2tpPlHhVgvrsHfO67CLbOZBNm
VU9G8qKjgJJlyDjNuZrCqEkSFEE4aDrDoMIcfMhCembktXp3+47yfoZ7yTPLhjl5
7AmD9cKa9JOtkozLi1GnVPYXZcvmest69XnWP6ClYsizPFtI1wtm2fqz7iraRD2M
m0SYsInJ7whfOntc4Mnkr6aVt2DB5njCXmRBlTVolyn9QKLvYvxKp8x5Np276ZLD
RpMiJw+V1YKZ0FBqYreDIa3gdh4+HnQcr/pZGcnNo4m4hnaw3ZMpp6GgjpGA6q+k
eea2+5Yrc75xtBS/hsxP64zH6SggpRoC16WtEUH20+4c3kdQJgxqSaPQigsXBvG6
/syZ8WDTx/BJO7wsAMZDaxaVE8g96u1gHwT6eA8fYvmxzLHcnjTiMMQ+saSyemJC
axcUrvJDQWlLBsa6DNleJ3/zz8DGfs4/po6BBmO6nFo=
`protect END_PROTECTED