-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0Lh6/8ozWg2Qlw6DQvlzvCJUoY6erg29Fv1kC6cx2Qp1W8MPrEg+ftms3aGwudskPmvIDXBQf57i
pAQZzmGFsbs/cjnqd/DFvYjCDQFL/gWgcWdHOVd8WtQpDQRCGJIdEcMG5wxLA3fuMEMpvvmhDsH3
JuAZVKj1tLIlkkLFBqmIFDCcfUMK8Vc62663xqXIkAwBCSqJbrICG9KD53ffYjK9Q0ThHU65e44r
RHA9kkjKPiEPrqhOyJp7SZ+3I1++ziUj4MlqC+gk21CrlS3N+ePsyM20DnE6G8Ut7s9aPeXat8bx
ob9x7a6AF7fkVwWY2KXbiM3d1jc9wm2Ne9kdSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 36528)
`protect data_block
TfXnQ8+DDl3n5oSKBlgcegpe4/7dNzSH8YLVfKkqyvE1iR1xqq/SHTT1lWQX7EDDpmKv09vvTIbe
6vfQ1KC84a4wbvpobZedEdKSGzRDq4KPh4Vn9JLFdDRD1geJVYFSI8jm8enLx210B7uV5upzWXG7
W7jne5k8uZe1RzuBbEfreZ5PUw6d04aJQxp0odw+7Me4iPB2aq0R3B/9usxrFJ7Jrxh7MMGKuMLO
gWjXboPIMRLevYL/PlBCCbaFMDBymKVL0IHFH/Um4e5CJ9MS6PwfaqnSUyb02yt6HDaVHT9L5cW1
eQojHsfpPl2tHaaGlvt2Y7582GqZBWXK54KFnqxHJh4PmV+Uo2cyOTZHJCwCgwMZ52GyqOYhuMpy
y914+boqUgFOC6umllsIseaxcAMMFwOkuyDbrI4WL4FAKObxABZp7JqScMxNkk8Pvcl7zJJwopL/
FRuNst30nT7mBye+dszWdSWjycKZr941It8bzK17Cc7CFaJpVRi1N6qOGfgoY/mCQ7IukKhLqjED
bOFOs07zpojtF/5RJibdoGzVGTb/ThR1yZ93b54P+dZt1e2rc9gz1RUZN4tH9wdlRMBb9VlDwTfO
Awtvbe3i+e+hfKp3C/h0cAq+HAeFhKKv2ysSVcHExsROpARr25StAhhmabkEKrFDAyij35yIHPPO
7inrumZ0x6PhwuPtYj25S0F2G5Gz1u+ioHorlpJT1np6z/OGwWPe2tuOpxMf3k1JaHkNJ75G8879
OQtDLJBo56bXpJZk28Ty1Dpr8ycEbswZkoJ2fjjCk7t548oRHfupCTjKFzJDwZs9Rz8wlHdw1+0w
FQd7ucw75m590MH18YfzrYYD4/E8GTKT3znJzPUfauCF2EX5Tv6dz4TQQuuhU0ecMY/f5IVZNTrG
uoAR8Bbcjf0mchE0YPJnCNMUivd9rI5xkiqkj6E77OPH1+FMVqouDPhfU8bZyrlGc3NTA1tlJHKw
1E+nDT4/HHeOO344XaC79DLC6bzj9Te7hXHBxgp+2QrK2P47LMjucZQo9bOZN0cxscyc5HlImH71
DzX5wVm0tzmXQq7dGb1XlE/twFTPtcKRfct3q9cHzIF9A2M+un7pbdXN31hvyACeZbylwyBdYfMm
P0rI1qAuGhytTqUcHzsahyT3H82h7noCnVXGZ8p0ilbuGPOlm4kILOdyDK68B0lI5Rrv2PR9bPKE
6holyCvlWbC97UP12sjY/mbD5bzoljJ3ggVkM3nSouuxHJJyMblNloouGAobkMH5+BvqnvzFcxDT
8cFjV1p5EHN6ouYxq9G/yU0l3taWksYXVkKLvu3PY7BD7O0qMy2Ic64vh9RWxERqhYsAdxoMPtZ5
1+3wu3o7it6+WZwLDdlJtTspryHXGTrBmvg6MM+qCZrXv7VPqEGd78mcjaBPN7sGjBKY8+Wm6fJj
6QOdyqJ72p5eucfaHVQeqJ5cMMBuQaJ5c66ZKPF4EkQ9omEp7MwLEOls05zlFoYTxQlQKL1/pPw1
G3ChtGO6u6Q9VOQSsekdls+sGHwFgawam7hvH0kHV3eFyGSotOW1BIjZq7/57hF/Wzk044AT9wCj
BNKelnbeJsowBJfIEFqSk+0FoWoo6Upo6mBuyVB69fLMNJKprfqp9TEAuplFe/osG9+oJJ4lsbU1
/c56kNMVM6R3M7WdrwLtBCb2pTP+iO7YTOV5L86MC5rtUWflQoTeSVU/sx3iNqQjHSGD1vp8maVc
gaO/hIRV1HGX/RRVLLPOgybjKZJNcPqLAKDRycUSxW3tkrZXXqxFnXdfGs+zdEYM756xS5pvSXPz
UK0iSYP1fK3cn22LXX3AxmSBMkUgbpbHk8ynRrWYfiBNB1do/c023p0kCOWas4h7GyFZzrboQHGn
iLXYp4qwnEdp1SnmnDufA4L3StEjNDb7/ZE7nRmCrey/QKgD0vSroLiVR7wpm7b7hTjMNhZt0bP7
88NhUMfRhKbmmhgzvl9J237A3Ng9aVokygSbjgxR8mq9kYDfjURlNb9gEjUZjnIywrOrqJ/RAEBH
WZIULf59b67/0mTa+oF5J0A5ZlQOzJQn8sMMWrwRZp269z1Rumt561INIwGz2uD1nYiOOM7sMZRU
tljJQPy02WVsJU6cnxVjBo/hIwRjS6YDiFIrYCfkNd4t3aVcWSdyWgtwyWqSGyWnHvfx5WMC4X7q
cQ+exZ5mZIKfD1qh+qO5Bxf+0Z6nPkDLDTy2pp42AJ7vaRohagQXlCEWNKgi+yRShlaOz5ScWUs4
zIV6mWFEVY70U3S2G2PXrnV5oAZqTJ1rIq4WR7JJZOb9qMT7ssvv0Nx+O6q1ITI4GeJXxl8T72U9
Pvi65Va8MNAaGsvU61lEOvysKreFyf0NNV9l2Q1/pjnkg1KZVuwyxjaJqdNHL2rtYFZw6H3nTq/J
Dz1ZozfHNhCEBXB0zELjg/B5YDUQfvBN3GhTHE2wXiBkeUUshcLk7pdI93kbY4SdPA963QVefD04
oSTlrcFpvcCus+ysA/c8WTGB1KwNNo3cdcHDsxajVGvtZhkOHkg5wTVpf1AztuaNDuG3R5ZQY8xb
prJcCE3ET2NDAq9uHTL+H6mJQtbuPoGEJL+1LCldtExLF3fr+LrmwIo1b5uwRsu+/I53Hdc58za1
okG0Dk9ZOROEEsIZwgcsPLEm2zsffYcVbpo5mIWmefE2FS4VYvFvpfk+BWBX80naTZIRcn0HGipD
Zte6YhyZq8qNIzPdqO5iTh2ivhuW/DdKSfzaZajnRb9KPTrqUofRX3CmrnjHJvSoHK0FXIMh6FoR
IoI29m/Ac5C4FQVKBQMsjiq6PWvaUMAXVEsgHJH8zqnfF8s32B56qq+npRwbcfq8E2z14RssFxdj
ebHagf2IxfSRFNviLQmVeVlOHPVC3KCydupI3G6b3xJeky7wk0QxZl7QEPCfHzFE1fmSaJ2Ob4p0
SGD2pR8JVZzHEw5toLruRuSAgu9MM2L3XIHyTht5zynZa4DbWMZ6x2GgY5r1wzmXcMBnkqqJvTqE
tu1MkCOc5SSF5AXGd046jK5Ns7+YRXZdINYTo/e+pvehCs9Bdl8tH75Ki3mAJcHozet9M+jJmG6n
pnMvcog+V9SzhqjOobvXLkWp7X8gK/zbkgsJSLEYKO7F3d9vsO6AQDy4P0X/FdAIaYMvwkrN4JQp
VDGzZp+RrPelGDTl384Iuws12FhoUqoeC9ngShKkS6s6s+Z55XxfaV80/7DqmqZUkzWor27Qw+y7
B/syrpGdI6eRJOLXqhzEGqKsgHXj/lha4fwZQdXMSt8T9kcLDH+rOyxetLgzNKyDWi/NjAjkcXg8
/8mXs0Wf5wBn5YpotkeCBQW3KDJ1/NFuWVDHoqcWwuggUDO+OjZxkEfbuZg6WML+ArFMKxdqEIyq
WYjGqhFU2HCo+rPieouxP0N1RfMKqn7qiOl1kmqHbQXaUPt0bUBm/p5pCL6Sy6TqqVxK+6Xuu+Nb
78jE+WQIdnA7UbajDB512mWgXoHBeg6NnrvnLpBiwea9vLEi8HU3QpXHYaGr3crr5b72rBtqCSqf
THVTwZ4e7CdgGg6SumvKXR+ix9+ydcYNrPrNP1lDE659s2qzVZqW4raFaUqmCSyyc1zBYDFYEy04
Ad/1ti7LetxOV0fOmOShH5le6WsLYxuUyvPHxLC4qS3BCsBteqj1fbOkJjo+8ImDaVc8JuAU2+X0
+JmqvzWhDqkL2tz2VTypHR08sjAzDBRzfuj7HY6vXveAzN4FQ9TP/bga1H8QMrHkBoRx5qk3dQEq
5kpwYa4VSbVXH0bm4R8es6jpEKm09AQ5Dq7oylAv6tMRKcSrv3VQgTeGEWyPKzMI/GNo6ipf/XPb
9aoMqbfWn81903DTgowwyt457xVWD9puwzvZkCRtb3Dg53aF8ke7T2VXGYFESTNQY2aOO29KCs1Y
vAzEI9uDYSVgQPJcSUdCui/a5tCc+dD4pySyJQ6TX5nfY+8h6RF7/syyfu91CL94iQfyhvVZGam3
nmoKq1b60rNoN3E02B0ClaVxoweYBEA9fn+ItN0Vva/v8g9p0u83sRXNmiJ73ncHGvIzbDiSbvl7
O0+IcsOBS1hiswSvC4r/didVHfi8XmKwnwrQiSW0gDcQ2JzKQjWdyWgF8f3SE9aaAwFKl/UVtelf
wma+rWywMa74LMVUQgW0X4EI/ttlceUUuYwP7C4omJ7sX/vkw8ewE9eW2dMDC+tapdXhhl4nVagV
PJRWtZbq4RBtBnnSezzMkiiRTnj6tqaY5hJ9HX/q8257rnZDLcwg9GBt5yzfpz7yoUC99xDfehZt
fztEZgfT5cWHIW0G3xL9mJB1jtbC0rilfyV3c99/Oi8069tvgNgk86+GiTJh/lOslpNB4a4EJvQM
rKhQ20bpaioNZigb7z+y/JoayGf0eeWhYtDcU1lTsXpY30cX51PmbRkLzP0UZhWbVpU2SQzED6Wi
sx+xViHEhxoqtI47rmYRoCBIXBW33zq1Fs9OrRWhglXwRjsSk8XijprLeWAVPc4sPw5hh43Rf804
SLatPwV9QlEUNuBFrSmUQQlP0tGZA0Qm5fCY3IHE5KpzCZZEFb4QCKed/vFo9zA8EhPDMp7CpcxG
J8o/lb6CWlLR22ffCl3mEyGaYqagJSKf+QLdq/wyndYZA16OJ5dOtK/nAXdD2EqHzTpII/59wkpn
nG/gUAs5Gi548iDLR5RJBbWUAxPLwPrG7qPjtvdbhFVwxbY9fsmbOuMthaFKdPkLBzWDpY+ToROZ
aWpotyGEn2I8X5ZipjsqIwdkse7sk4aa214bcpDIdMIoOniW1nltSRx70HihJ17CqCFYCXhw7bDK
vgbssQ8sCoZ1xV1exA7WZAOU8aYKWaH6HOwozOnSLlU3jxSpwBQoXQXVHHNVjm2imvTt+YAoKGef
+MOQnE6S00QR+2hzhTM28amRoAj/17sUqkxSCvKZpUFkHAYi69zOw6jy9cdhWw9f4IaZirWYcGDP
jskI8xZpqMkZeK7v/2sdgp3p3Jor8VQ2uZI4fN6IzCnUFAA7GSeetJrzh5bp08Sfi+oTMN2KVb2e
zVnoqxYPOJ+w7iuukGY821l+vHjGtxqAkgqziKcgij5XKDvMJcwzNbFN6OJk3s/Zbr3jI0MRk0In
zyw3vEnE1ZbKfD2GgW9BP8E4uRdZrNxgGALq/JRoOcmcmeqUzlnCtuGxJN660CRkpOtE4sAk89L8
X8pmn0ExgUqY/eLyAFjsRIFnN41N4mnFLhzqpvfcNejJinjOmRkgMwh7GWQl0DGa4FrrMGCWqLoO
9kV0vJFXSK7qm1qMU3V9i1uzhh3qpVpfBfL5yaJj1bKZ65ckB1hB+rLe/OYYRxkQ6FVgau8qdD5g
hpQwj+d82Lr5CmX77/zbV+jHf2xNImDS3g3lBlUlaQSPo74aobLfu0jUF//19gzT9hAFbgD28dAN
HJOWee4VVLIuiCpLwDpoSPeWK85siOgWGCMaP1yQ0bF/snpZvA+hmYeFQZidVI95ikBPHOS/42pq
m/SriYAbQRItZE0qrcsq2T1+yX6MhTGsfxfNZdSKtmyz2Gyj750zTPbJfOUGv2m31WASvJRuWoWv
/nrQ4zjHnmWI6fRYRrEo+tQVHWyySFKvJVxYuvc1S1dwlftyL3wY5aW5CWf7vtwje3ZG5atv/J7y
5Hbp5t2r0E28w4XTMYA7Q3eID9thCZMKR0z6UAAGp54Zejlz9I1G8g7J33wCqAT44lt6y/WkiGNU
O3ywrihj9CCifMtpWeaP43DAluVsHxUBbCZZMHHCqVOAe3noqBYpHJk0yMogij2O8nCggNVOmxmc
0wN8qMeC/DHh26SqV+qUbkIoMqucwG1F4C1EJnv3qU1Has+/slvwH3+SA9rIFv6Y4xhAolKojQLZ
5YoI354jyPc8Iuuwb5T6LFLpTZcLq7onOZ/7P/36RstCYrP5bsln0R2QtlBztfX+PN2HD2sWAXdt
C/kE93NnptxLCX4ZllggGaJtM0jlPS8GEjwqv8spgrOds5Y20T8qwX0zO0IyBy/DKA9BhVCNGaq7
Hz+o3RQt3smAywtq6ZErF69loiyMTWkGeGPltuKLWRLwqwQM6XfQmkFR+3uFdJcDogPN5ZSgMEeG
icvGySOz8Jftidz6cn1fNMe6kz7aalE9JluSACYfGymcxgqJXz7Or9BpSvFw+ogbhVlEYnYHp0Ce
4RJl7BtMr/l+W6sVN4hH4hZ51oSj7WqwOPPtJ5RQe7baFID6pIU4OBl6hqhOn98WLcAOvlVSP0Cg
cA9jblKSzPrVNf7Z4JBcBWGVHN80ETu0Ltb10cxrdOrquiivVK6oy4+GGjwe0uMz0wTHvesG6i44
3GSRsQQvCv+ymFilQITuD1Xb09TwoyMeqOdc9BWjX1N4YcacXZESKTXV2QpYiKZoPwBTqhtzwJOg
NUSnIeISmxANiqaqfAHCb6cD0z+d7WqaYmcVFAtQ9/Zjg4GLyc9yLzJxu2fMgyPRzVsjgO39J0Kj
q15ULw3E0Oq8ZD1am7R7B+xEhx5UZuIvTg0UpFrYJwBjODxWCMxlvTLL/olrPlnprA58T47jHlIm
hBQOOGkvpEMrO6Qz31ixEPRBXLFPdpBqQ1auqxcCn2kQPY4MWZEprkdbs3eBzKhRNdVqu3q1U9NI
HReqb2/Yoy2QLfcbws8Sz12e0CqwYzBfXw5OBbXHnVceiAhizgrINZHIdDvMt50OExhyQw/8+usM
/33/9V/4YCd8UMCDLyl/WWE+aKs66PyxbHY+jBKSICBIUebf5gunzm8QUtmWsZDIJcwjYAOViSjc
4sD5JJd7/5mIqLPs/hPJLuMKk384nVpKEaVGcgQ6cEZ5/bb/UmVekHNW1UEtEf4cRkwp8cNl32gW
ri1vT3KLSqwMwmhUWMnpGLJvVYwwuseuJvX4ygimZiNOK2NJOkYFtOOI2Bx1gKxXXH63N7pXtkTY
yh9cM7vv51XGMtvCDYinl4uk3ezwzljL9VSdhi6Ytm9ea//QKFqQav4FhSzhQ0pdJrajv5r4WxQb
N+XCe2H7s2TBUqrkwfdfnrv/lTYc2xEhPeBbhz898ILtkz1LASzYuO6wx4MQ9Dw8iJLjTkpXudvY
E1Y0nDSbQa7UlInQySPncKohxx+JfvlotnQ+3nEWdnnTadsLk5yO2bi3fO2/F8leVbZWFGLu/2ae
Tun0/bHuwePyY1w9DGtj6//oYDSYWTM3vBVyu9RA6pcpaArEhLyzO8MJIVPYkqA/PjYeuT6QDW45
JEG81tbHQ3jua1HKs1yllioofBMEdRCMuBegz5fmHDfQRYon1nJGaiDM/AfOduCtr1iiOITbfZ8t
v6DHPpVWS+uFjHantaG+Sxm3pYPEpDt8d22GhCNYoYFlyYsEPjdh9AfY+LjFSnJnOP2EiAIVTc5M
h5riFKm4/2cRLcs2ykly4eDfv5wYmaN5l4R3f4INz8GHGRG4lAXub99eQJS8ymfWuqd0oOhvuBTB
AwQonj3HI1JdUqvRZI4+WlHQTaH6AgsadWgqbBas5j+9E9CGnEEPzKQ+n5WAvflM68haSzUNxZEI
m1SvCdkX+awbjiLeGjlWnY9lTU8yjOMCBp3CJ5oiKhIJOekqcE3DHF80K6jeD4OP1SGg3rYl6xzT
wEsq0YsB+obEc5c99GcykhTM/Zwjr8PudSLr64l6YuE4doD91Ux4uXkIM6C6RHiXCWAPE8uFHeue
N5kwDghz3zWp0bvS7NNOu8vVv4yQnniUgkvZEyZ3Oqj1Agby/KE3Vspc+alk3+eFDyqhKI3e9dLL
87UMoX0ok926LBb+BOIjP1w1oRWKTZAZExdVW8wtSGTyRDf8h/44VSnRIdYxcILN8+7JLlfGK+qx
XoRCZf6mAMjQEGY/EYsSnIuaUTaSyP9ZbCSHKDP1EIz8Fh0eGqswn4DpigY0XZSxdFGdr6oIcUGF
SlF8adMgWfL0LGdunU12ntH/a+k4hSF+hwqKsLYj+e72Xdso0yLBiTpUKzc7VPJ+AU22gj3uptym
1/py87leb6NkUseIvtcGCWTbw96RcpBSVJvvAAfox6AJy5b8xkgoEPu8qM3CYI/88fzslSu5C2KS
hAOdIGVuXrwBe+TK+G9eSalGGVHu2LQAdZ2TfgCBXvmu5sJzboAd3H1/2UkH8GGD4KdfCwk1c4ot
gVr1nIr9ozwP4xIm03ElgW01/rEMB3/jLxIfSiGwY6XZ5d7Sjdu1XbNhoeUdZ8aFl47NQBiwmY9M
O00aVyB4PZDufj+0PXFZBZGRZBpO919qYKbMNjjlJNvITf2ig03XPdw+/YRIVic2qI50WaZ89ePC
fYq/cfFqFfSEsn5ZUrmgRBTQNP98JpwGeCQ9r7ovDG/10SKd9gi8ElO1OgRrf6OWEKM1jSWO+fdc
u5U/5PS//AppuEIcmzyncE+W1A+SeQE+IRmGukzSvzpAbmSVjMBIa7QiWGL2aLAYu/pHoywMHDxP
c5vUhOkKOoez/ZpydY26wXzPN6/oQQsRt+jRyiEt47artJhYSzTiOeNvSEcdJ3kS9c9SKqpu6j6O
/lvY25ET0qXSs/2skjAamrov5UPilBxCD+0vUwWp9d8F4LpdrBplQFnd8WOtqhafpeXdEHjqfJX+
kksGtpdB/9N34WR35OV/bwC4UdrEV4bE8QPKQSd1kQmW93M26ZoY8awzJb9fJeO7AEju7kF63NZF
00YSQt9pwnLhRBN5dQzm/nxOcEurUiX4PpSseFTO5+48LGpZEdFDW+4t3OygAdSKHfo1EYQOslW6
nOwxeml4yIk2dMRMStSA8NetCBKbF/yWsZLK72egNDmZp+d1h7FqbytMSydQxKSqxqHFB9IeKlNp
vuYYdOi2NMat++xjn0uxUPPG0WbCCaI7tYWoHXWLUVXSDsNlCNFT9uR1CAj2FGBMER3rZVz3ylsA
+E1jlUl7Xvivk6PdO7OGVNDPwENW9qmvoGaDQUuAzgjIZXIiDgejX0MtdnY/FwwkcMDBm+S/zPIo
WRtMGicsg5zjr/4Pq4tty2ft+9ViSmmHfDrhJLU9cwj0Hm/O10F++W3UC72lEbA9Ael2JPjOfXMn
2vk3scEskDdbdmUM9GA/dRfs5qbBS5RCQ2C934Yphuf5082UM/rIqHUztqyjAge/cjP/ceYiI27I
bVNTLm5eF6BPTUEQFG9k4vUSIsUAs2gX5q7DScxAdAcU7bHY5jjibzEhwwj/oOV7UfuMiO+Jt9pX
g0MqeuNZYDr5eDmRlLiNf+/GjXr3gcz5TMKYdIxXpPcw/LMTkbdebDK+Vqv5J+J7g1gGEztLbCm+
yk1R4wuWFDcwBXA+iPYiRD75VcR/Ndb+lT1hcPWxHFy2bUXp64u44bsLe6hgDKdZaOdZGxTesKkz
DwteP6/8dt0gFCqNl6Ss09X9ZomHRFcTVt2XlSPopydHvUCvfmbIpoDJ6GrEsKNtZTHhAKzFUEYq
BjXQFTSPHkwyTQ4PekpAImCD2kRAPhkaodngkJtR/uME8CrACAFrgws09xDIj8R2ZDAiyilrVtrB
R7KILzqSsYZBbWFNuHqmJEwmEfJDZhAq90/KsUD2l8/AjP3P/p+a9cYr1zNoM1OdqBfJXbamw5kW
0kPbnolXtLkibGM9fRCIaiSMZCGJdey/f2fgYa8R6xFu+Dh32nFlnBI8rFo+JFRjifZPjhCpPZPB
kRvi9MiGYFXhezZx14DPX9TfPYTdUOpWmzMqlk7QhS3NXeFv6ApKzaflROJfyrssZQRpFB26M0yk
lfJy8E90tgP+LU1iIUbd9luHquUAlCm1FD4PdN38w7cutvUYaRhquNsArR+7ezxmXXfJdtd0GZJY
Vzo7sIlvIPNvkr4jh1c4v+kS4XgQSbpZ7ON0GoHwi4U5QSek3kHDuSE4en45ukx1gLbPZO/hXhR1
OkpIu+9duzPuHQquMQUx1NjmQU6yYXwOPKJRE/lh/x1HDvgbLZ3ngNLdU3tkWr5fC+IlY1v/L1To
Ci4Gq3MK3OFjYpq51odw7Nzh4Vlvelz/GgM422GnpnAKYvT4/BmbvwI/wD5CR3/EMkvzthSJUrmd
ZlN3spqucVeiNmIwuv6MombQR6T+HgEuou9ng6cdN2aTbn9OCLkN0+9I5j8mskbBXQbmHxyrXbCF
6FW6fTQHlIrgwiDPWdGsGniEvw5KjqIBuS3z2WwHtEKWl/SHktU0+7Z4ZJ1gHUzzmJBfqf59Z2dJ
niGKByjRfe1om0Fl51TvOh1JbBEdUbOLWn0+YYgxDzxZysvmWUzsrWC6W1H3azAJ0qjhfz+wDC7D
Mwa6HGmSnJQutrWr3KmBHFQhrMCtLFssZ/gzWXt9MplnsCJAN6C2qVvAmORdnveBbuRAKCY8JZTq
47q0C/oYhg81UL4mgK0jQAD4wh1mCLN2DbVxwHDsCPTBJZQ5BYWPxV34kXM9rD36nAFF6RIODkFz
3jEvFY40aZOieMSD9pco0euXZBzvT3jBPihlsswea4FBgwROychrPXHF3NrxSetAA1XkY4ZT7rPy
xJr5Y+yTyJ0srKkBEJ5AvzjozkAJNqp0Qj7/xTLMmwkiEi6BbMx15gYNOPmdie8NG79t61V4yWUk
7o3D3PCXotLQKOerYCMREFKhp55XhmtleqdU6B4b+4o2iG79a88qpge8kAlaPij1nCYnuVyDkpJa
ij24GzlvSFBPObhnRtaiSI7egxc33+d9vGqQgOlpr0LzYKhYAR9vg/0w7Zm0VIqzKF6NcxBNtT6V
tdP0VhjR7BKY2mjuRq//Im5zNmoWbcBrJhFw5c16FG/Mlef9v5x+m0nSl8kmAonT/x4c8Iei4TEs
DF23e4W5Tkgc8/CmwQVMiAOto1BY5mtqDC6kfivWuLIO72e1xyV0Bm+RB9VbcpC6HHniXh1dtnNg
BRJgepGtm58jN2f1WR9jHOGJsYFyT64JzrlRknu8x4zwfRfac4aPDdnTlg+9stfT2sMyAYXc3R0u
ifXTiRQW5zLlAxLC5sVxvgPno6bKqcA7TZDj1F1WwrGJgq5ehSlMJsR9fl5qYT6CcxB8bQ/GPAX/
oIFioj+swVoMePEYvRDQmIFSb4lYbQ3Muvd4nS37sVLAR/Y94IcN94aC5luzkZZes6aGxlZR8+bm
FqUMFC+nBy78Ix+AfS9qu5PhdMhjFFmRLflYNLL+k36H7GvMPratUUhy1XSKJ0AAepK6KotVwF9O
Rj8Gc9A8XQTDj3YDliCr+SdlKXmBdBfKf/tl6A25EcWJKEFUtPJqdRwnDe0khchPIabHDNd/xQc/
7A4HRoulQI2QLzhFZpD1sRnszN7fXVc9M2J49m/Dl40/9auMiIlOU8Xg2B62nS8Vp38GKVmA5pCa
fzoEkxkJAE5R5gSgZSwqFpealWwsZLSRLGffmnmI0JcSpT37IU0FxNByTLnNloIOtqEh9lH+zhNw
jpKR05iISCJDjNY3HffmGZBKHx4yAohk2c9ywyg84Pq2tvguETnUZycKMOpZeNNGXa0QSofHYTOX
OOtPNhjC4IKAi07Np23SjuDlHoVCWQqcsLK/VkqLj9wRiGr8eK7Np7ngd7y1eDY9ghbYjbs5BcEw
6mmo6L8YqAc/6EIiumqX2OQjnE3FDGSKkh2t76yotMzXq6pYYOr5ZLZUp1xtDnD/IrP/AJP9O+lc
cH4jXdm9ScZSk8lgjG8yMRrIirlaylabwYEXAblqWfiWfL14WTCt/XSJihdNuxSM+tDMcvA9VwPv
9HSM2yKrUeQGeEpnys7kkWEYhS1iDsF5zQ4jxtjx8UgAObhg3FJ/QKTwq5V7/QdCAtsUSwFc7H7S
yiG/B+FqryjB5JTqRvuoxNQ1GNUWTGHtukpXTR16OpzIIwcIPrE7x/054MtjWynrnKy5RJvH2Qmk
wej93fGFw0dOLIBXRVqmF9F1roPK/yJ25LJFp2z41AoPNGVxpZExcXj94H0mrlI684dz/rxIyZke
j33HNtXCddSB2i/2W9roPh6iLMMXTFvkUsTLj8tRSB5J+KxO/4qUX+MBKdQFt6IFQSP8/JYwLGxw
6k5cpceKeGrLjllGtNB+7OZFkOcTm/AqjP0VtPKnakibg2a4bev7Yn5051snFa55UXW4ShlNJxtg
ufZLcu26xueC1QoGkS9Xf/IaX4t2BCHtxzcXN/B3lQaMI9gMJ2hSJsNkA3gTYDEaFyMD2AGOoV2T
3Yq3JMrGHLfjnP+wYz7kDQnyaBb1qjkmyycGZcspA6cpxJElXmwe4xWQuB8cQIX0Xys6mKkm4Zja
E1iZ1vYd1CeUbaK5gbGBrd/gOE6vVgEhb9iVxu7tfpV7/QVf6NNCnPI2M2doEwBv9ZBlnHGBMO+5
849v513zrM9hb9WFKPCTXYDto5kRSzFb4iKw6SPYoaRnTTEpjEA7c7DBnEzRBxnhwpLzoboLWY4Y
N9wIiUpM1JKkU23+r0/1OX/3XZ/fviZczqdf9osHqgoxaWsTlKFSXv2bzb0eE5u0+ewnUFuW9i5l
o6zTiwsWF9uACCUbjDTGs0OG/ZJVCTGqG2Bqq0BwJ9J5rl4mK4PftMu6HYSS1YXOIiqiSlSi9hkq
HaDFg0g07SV6Vpz9aaECN7YDTIh0GIQNQ3gyrVLvQAsYrm/umrmCyITMupi4RCLglwwzqFY+HWVn
Zc5aggbfnrwywgnvKoVBYwgmVGNBGFzidKyVIGf77VITRLQ4k99OwxoOfjo6YDgkvpULgj4XeA4Z
Gr8Y0DzG4XTNk/l+9zjq6Hf38oZOmYVGzdhEhQxSqeWqVJkuHQ8HUyEXao3CqXgKKNOwSU5Kf8sz
6Gnf/Nf7VElNELIc1Z1/NQ0Z0fi4kwQtA2d9BP7EmMH7dM7+osZZiI8cg6tCP1aJEwxkSPZysKSt
Dqog0Xlt/Om8PzLyPerpMu60RIVdW/wEb1SX+MIxUjmHA4xLdW6YaFVcjG/DUYrnD6UioLAJkcGr
rByer0uGbJCiLi/wVUotAsSjIsnbhBV4IhySWBio/7I9O/p/wiGfzCv61BQ6CtK/uGHzRkRkddMN
Wq7wtvhVJ7Oa95SZLQcQZ6jaXVyXdcHkPk/xM53xNbkdOg7WRai3Iyl5hL20I0eECRGy6LVhKdRb
KzrWTEXLm8XKPxdI8QUxU9iK/tNjYHk6GIyrOWBNOD8enYveZQNEIONnmxk4kAwkAs02e56kBR6T
QTBqACEKqogTiINBUvIGv79zWS6h+kDHSvUUsPX0mIf1EDDfnkU1+wfy7ZXVv5rCcdQYKnYem6LB
aYJuNaswp4AmaguqZw89P7XF1wZpFsJR/J8DA//4XDG0pUT4X7/isxdXLyPNNa1ug+rLjHtGAJ9L
EbL8DF8/u6rOnOoQM03WCAjAxRX/Sfa+YMeKh+fsr1svU436MaLiA3yGVuiNJDiV+LNTwIjxGDxu
DW30r2V3hwakfk4BiuTtGITOHtOkV/ebyTJxg21Fb5ofKVDOq0/iXEK9ToxivgB++vha0pjcBIta
txA+pJDR02CrrqrgWaoLDum5LlQAAacxB0XyitSa+/fnGGMoKDzxjsRGAHLCJeR19ZmET86DifjH
71dIDCRc5CGmFZLIPhhI41GCYyaK5IwGBsVL97C3RRKhpkIzmJ91sX2VBmL+UQLPENNourHpxkGu
3oVtBq18Upz6vDCq3A0mzCwuYUyto4BdExeAxzBxfyAbmqqgQVHtztIytosAPW4PJKGTh3qHH2LC
zZXaHKAXZ2g90IEyAL9e5+6RlcZhgKtMMUjaGr1AJOkG7gBEX6t5Nfd7nQtaeyHXJLEhHEMeDlWX
nDEih+OpCQYsu/WXkpPTQw5HGSpxdc8seO1RycXAOLD4aE/iUgxutBjsc+kDpXn1DD1GqQUakuh5
Qc4RiDakO+CO9BKN2gRN1hqgHMAgrqbQrunu43E4Mi+fhrE+dBr//qh57LDO1Dj2nHcCGxJYbBdV
y+8j1L2B3peL8+SUM1NWWfJ9zKBGy44K1AJ1rimuMvatOkgyI/M4MivxKDHMb/fsJ30p3+GKivBk
3/7MLJZae5O5b0TZPYbKUdtCAh4krwj1D7mYuiLcgPi2sxnOVzdhtLjI6P2QkuqrEfAVQhFkYauP
2chIoFhg3J07JNeehkfu/Xzm5oT3RuiN5+7PgYVZgACxi1H2cQ9jgFnN0Ejrenyg7rZQNw4Ryo4T
+hJHYpHWMdopf4a3NP9pWRrzsxE40cAGHXBEkNk2SnNlJmmAO7+nbIhlbtJIlQ4kWQMCeGq0jG1/
XRB3wKFaa2hKUnz+LsCFZ1KwOJZ+mjTn2CTWhe6dHr3nhr2mezH2xKjTTtyVnoKcwNmvwJe6pmxN
/cN9GJrE+R2R8HWPlrZejKDjcXZiTpkvN/P+GZnR06+YHNp5bb9p85aHB1aMcVE8j9ECUnmA4L/L
qqD1wqZmjswnDdVI32+kUygG6qE2AMgmhx09rpBNv5w+cKJrg+tZTCctC1vRgUBknol73aqxv5r+
g926GfGLWT3OdYYzRqbFv7qdhFRivVStLsXkXRs96WaxnZ3+9BHd0hRBI+C6ZgD6VsldMmxEyW1D
FTvDgWYv73VL+hnQI06qrTSTPKdE6FtDY+gO2zbTOOiaTZU+zGtPDKzxDogDmEvdG11vtl41bFRu
4YArGts5XHMXnjhIXeGe6oJYkf71xuqvh9Ie/3KSCfUyyokbt3QIXcrBnm3ZRCKTuSL6d8q+v3iw
xTZ1srYYXKspiRhgOgRqQMbwZOZEdIWWVs6vdOnXRnY/pV53LoLpC39BDBaTy4NMsGPkHBtiVgVo
IbcpLAeXanUHH0KobD56yf47v23Mot5Gn0A8UExvUKLV2h9GqDiHCvBuIX3DKYPNyiWrCZ1fDU7G
B5ma0Et+mXsfXKxYY1qYU0VQqJeXiI65wAd9uil2lHW/ot3jQiACsDskp7W8ioMBEJrZEYrHpYdy
ZAdSmMSuKc8pcxx0VcmBxckNFgZREGsTjXQ51IVSHpLHjwkKv2O2Zv1nus2amsiooSs6ZgyXufoh
OSO10oTBm9YuGjI9g/78umA+wHOrbMHZx5z4vzm73HEB/G3FTnj7PNPMfOpktVQnHVMKU8YcS+fS
mfOK7HdWSWi9BJ6XHE9mbAli9hjExG45Z1TPbFirRUgkxzTFinVSr+xXWI4NmCPvUSVCF1+rQDZP
5Gs4kQZMX3lq8UMPXFzfhNlUswvGkKgfHpO3IXxF6stNibEWyVkz5xlXjNWEWmp7vY4GfwWgyCEu
SyZXE81tJv0PqLdp6zV4EBpn6uT8jiFGU61cTx0kI1h/8vqAngsgAslqMCCiACYEiTnDyLx+fkOc
IwIyiX8A5pG75daSKgg66OHGHBBeilyTBKy+ywh/nrko9NPbK4q4ha2ruFRm83YFYebvSaN/miky
tM9InnLtid9EQYjrq4er9XIYuFAeQ8C63VFLmE5TMnSAFkjM8HJT2dcS8c0ZjhbgToVvAfYYpCUL
aL6GHtw0cIY3sO0l8mltOwOniOda3u4q9Dutvzo0NGY9nPOGzEzErhBzCiT27NqUr8khc+QmiWiU
6Em7ceeL0Si25eB9X74X6e/QUM/HQYnVRs3jfHYq12AxrwgEp9lYkjFyfI0FeUC0tH84hPu8Hz1H
H6In5uXua1O2XAXFYskY9UByT4Jf62+G9UWlaiy2e8wKKerT8EYf2XmdiyUjTH9/inEMyY/j4kBJ
be/ud1Y1Cz+XUqtDiTRiQQfxKMM5hPNJcyBy6RMZRUrt43NbX04jyoojenj4eENGspAKfNXkZ0MB
+MucvDGTa/6nJuCPWDjrdmdIJL3ZztPIoOhS71XdvVwLxmbenROwWL4gpsXMkrROUeng5wl0VXSc
VmUdd8Upt4F19aSogKEJXUDSmhGxGNcHRoKZPF9nFhMn8HWhGsMxQGwsmg1jLC5owH4QRfO42RUx
hF6Ckl9GLi/kTHjQqaeT7VkYX1vVkmco7teg9CxnXxCvOxFPrpBsIhNPcG1o54wx2qfoAkd9TYZG
NFebFTwWkSa+zp1lJNPzNF/1cBP3mUyeGxDD5AX3dAFXL2nfh1NO06LrkB+ZGexba3zPKK8RCtcA
dcZZ+DBE+oixtwxnlq8FzYYvro3u7dDvPiKy+rOaytN7m3gVRCbTBcafBvH+fC3JOTaJLf+vYjsm
EwSvQiDjA5xfsRrlCT9sOIbDLR17W6P/skpBz25IF/sSgqg0HPdTdeicp82mUcd9sDr/NEGyer+x
er4lWuC2z3aRLmWNswqy5lD7wuvPc37UpK1A8AudKLBxbA6Cn2u9714Ry8FMp1p244VT9DVZokqZ
tVKZGEUevM3yFrjsUmHacZIIm/5QMzVGvnJeFrFXUPJRH0XXlGzHBrm7GKshXfWTiLpIcGN6qPuq
/I6HXDmc3t8OwCOtf42Urja4bW3h87PbJssnUdUqGbJeEU7mExEFG9sMzuZ4vEV3ruZgeSlNKzeT
cIFSkkK7QxF5tkqd7SBVLg0I12banHhB773HhVwO1xGKDSXdWGrEpZJPDszi0ch2GbE5ZCiBTuJH
aq8poUguiLbt/hr78D8qq0tdboiYt4J7HYyBBjzDzdKUKHO7hZrVd+Vmifqdu5a/2KHIRC6gich+
m5zqe+0OGo6YmAvjU/Yv6BE2UP7maVdZzR3jKBpICzpiXzZvt+pc3LjdIFcGcamyVsknGyX4rPDw
LBNxecy8ZqCf575ygxV+Y37gcwXNbs+WZOfw20SyvM1I0OOaBE0A5/2hxPAK9xm4c4QYDqZOt5zq
hvQREAd6tTSRbUhSaRF0dtKu8+sMU4DVsmn9E02SZd5aDgqcrZmmBbXHkPeVEKS6lL2wry0OQpSx
oSGO4hueGAREuOXG7dc3bQnLSc4sT/31BzpZ/UsrKbSUTyjfcmF5DyKtJbZHDTxZsOmGjkmsQim9
f2I5zRA94OxR75z35I6pGr5+l6ClPpXUIXWKj5wqJdqunA3nl2ECbrrQsXseQson6/IzdgFUp5+z
zTFb5u0q3tJqYe0glqbn071CvlL6SEis6Hzp1YTk7+DAlu/xIG6gJRv6swAtdkEwkWPX2gjeoxyU
fRvI/fmrLhj3gdCKS0Sl5KZuWdbAHUNt2eK6NB9YfzUSkKU2/NKjZowVC5vB/huzqRh3ZGpREtC1
oUXhYgEh3mnE15qsY1Ys8hM8TCbLXc4L38KQ57MNLQskHgPXpkPL7FGuQrFgpiA9WFLAJczrPy9G
HfRKtYY6V6RmjH9LADodYKLF73XLo1A9TnIVpyrXVR7JQWnJ5MnrogZWjJv5qdShEoGUZ97yPMkh
/tX44n7Gccz81hvjDj2r2xzjMGwqXiZqUoi95uza89pfvmnkrOFjJLxrF/QcKSV5W+vJL2CgE5/t
LS+PxAIsqhATUfh32Vd/m21fOP80OFqah7IYOhAr0ZWt7uvrzVwhDE4tOL+5D8JQmK3pgfXEFACr
gVZriOi15N1yyzR94MI0EeY4wdeMzMmTyWpzAJBIVkLW6WtJILKig6yN85mjP65LiWqSp80MQBAq
howGhPLveSaZlFjWnFHVc/jYdXP+51HK83UCFKoFFq2S0Fjr71mvdKyxdK3aQXE6lOX0nsjVNtiy
w3J/oXkIHX3rzizXiYLMlRPtnD5BCoC0VoBpkAuJTTuc6+xLAfPVlz91MAeSCMVTvMERAQtaxDbB
NtGaMkV5/WhmvdyTj60cTTXDB7tXotHZXpHEiKNLJQEjqRYsOw0szhtcz9B3m28nBNStOM6j68HE
Jiy5MuZLxjJq2iFcuYZ7dHmKw9oLHPiRepZ2zHPedljzCOWw1VqWjFT7N9KlXzCs3ZBMft/TrFsP
jXHhn6uyguxoeFTsA1XWybMAN1YDGG5K3mdvi/3k9FBxY/TRIsS+rrFrkdzM1p/eTrG2hqynjMwZ
cU6j40xx2lH4VWKWCzUh5YdL7qiDxzO5czQ93MrKtdZDWAfHhuqw30xUZ14K52PIYDbljFYT7T56
aUhLbBnr8peqTK3+Ltw/FpweCyXy2llkimdj0xQ8sqobn/ijZQ3jXWY8a7Oo9bNb3fJH52fqqu9c
dVWeyIyRcF882FqAjb+Vxs6I7iKgoEZZvMGFjPh50Wn3NfBHikkavq/dMjW9eaaRJ+H/z9NZT2VY
BcUxntmKR8syIj4UnXovg/58b6d1qoHGYTgWFmHv9uEdYBMiu/DkwU6KqmkjSsRW17QvRmg1iFHW
cWBHnYIVw5tnzQ4b6YIWjkly2e1bXq1txsjYrky5B9GvzCTWc1MmV/iPIEtf0BwpFZ0ECGCtcsdW
EeRek5izx5PXbgh4DvYVkX0U3z8VGbNm9rWAr1JNNq8PDj7FpW6z33zGvp8qwgxoNbLsc1PFIcIK
K/m1KjzZ7O4tFybVrQGuL1pB/BjjxYTH/qaABmMZS7bWhNLgUSn/Fb7VHxg9I+kObuNHOwB0Cc84
GgWlndHJ5BlrEwCMae5X7zoTD4wWLE7anUfCz32jCZqxwc1o/ckWMDno/hfpyjxdooYaY+UCo89k
UonJD+M5H7P7w7GwvdqpfrtvqnM+7We91+IZWeZGZ4ff99BBAQAfkZyJVDWXgypYcNwJClUVv1D9
uEY3T0jTCRfI/Esf0loTqWgaqkRmQG+IMp8bESaS8PduKbPQBqvm+vGC5gfZNR1acBoyrsVf/hRu
BjjHaUxqexjsH4Y11+//7cgLA7nh2j9+T9DlBIOMCDCPl+TderRuPp7s0h8f9EozwZFfZeFjltG3
0zzJRYo0U8Z4rk5L8y13JBhrwzUaxP+ne+2H/c587FC/H5SCJfNQg7nQC3+Re1VFMG6BVpD/9drU
Q2ZfNVvy0Xd6grwFg7DqVivFBYiBNkuNcKxonA2BXzhFoJhVFn24G1zdgTzNSsYMcv25iewLPibw
MUXMzD3E03PgmmRZVIVrsyaavRVl+SknIhDB3wLXV2VRXiJiMfhl8JSLSGO0/+YIAeZD3UPI+DJz
/fahtMgZSRFA17ZuVhzo9JjV6kfDP5OFFo84obmFUpMQ0ZhrOlykDK0XyMFJ2wjqMzmxRLJ/NL1b
ytuzYI0HOnR10vooJ2FtoVHRxXdDbJcNjpAODa9CCbriVTNmZbpoMCeZmAs5XdLbsRcHnfg7drol
9lyMnV+xAfFOaHLLtkTaL2mhDmjHSKWnogicizDHNj6vf2/A/TSv4w7nnd2OqqMThK3GNxaTAchv
7MCywYRJyQWZgk/L/379GCmBJRUqnzGlfGQKvjiKUEY6rSG+pOb6al0DWXwAKhhhgvBYSNtI5WXA
HxNdT6cOqYJai5+ZQwNXzE32Tx2vNEkGGDtsTpoY9V43SPSw/ishiReza4FuAsdq98GJu2+nOlYa
kfcCyhByIsx5tb8ggZybs84bTT40qCkWiCW6AWu1Cuc3FA7BJJ2Z1IYWTh86tH4r2kD192vA5NGs
4ti8tYM9dgtV+qa6HMDYl0Y7jntko6Vb3XBHCDkCzViQws7Mld2xRY9pPqHjLVfpWTNvff9vErcl
BCtdWpdzyTqMnBniWmN8agbmZGLYBqwgHYEnDf8fb0vgRC4YFuH69iUlITDA5bh6ctbjotOXbkdw
Cot1HUgN+Be4LLaYrUnK9KJ5OUJJAcYQchrnceH9RZusGozZIHhCQRvRbjzIQnn3gYs2Yhe9kYgh
1ktXMjZfy+jC7tG/W4A2S8//aN1iZRrcddksIGwj5nQLsPvJe7HPx2IRUvC37UFvwYnLxYsXnbhp
2JHirPBO3nuGYzwUs73q+hr4/ZCrdWPwFqZmOlJNBRd0j/hSYaT7gwbNaGlAGf1Xcm8Rewskcrqe
2xvYuW41nPuQR+CUuzXuz2qGZWieGu1FDem6iIrD/euOT5igyeTkXqoD8AF1T+9z/9ekkkxdBg+W
9Pd7Gr9GFEwG9Kv7jM76N59BMBReRpkswEhN6YPnQu05SClNKph/RcqtUB5nvWbDEcEvta6bVmma
NqfAk+kizJLoR236sRsOMJ6dfpK6ALRy/TBbzAkTL132Y1UPW43HFfC6VSlx7OHXDPNzHYrm3wmt
0EqegF+2FiE1FxZ558XBsI7bizbihfvj2qVpE0VIqC5oBzxt0dtt0y3sjNkuRRyab2lKHhi9OL46
Zm2n+amKKaYo+SgEQdOKMjhljAF1owfj9xjY0AbYJHvA36USM2TUhxOv5sqTQdfbhyxnKbF2FbCa
R/rQLOc1C2mJ4YQYFuiA9bT2zzMhTOQMsncTPTOfYHeF5eMsh5hW7tVPrWY8AkXV8qoxh/XvLN54
f8QJeBWkvjmbaTYyUn6C0xLLwdiJITO4NA2JeziYvt8KarcI7G4A7mw+sTArLL+htRUi8jjaDxyn
URecRaxBho+BixFhYKqUKNf8J/TuE3t3WNKklNQ8HSchWt834HcDwbQAXsNVB3gx3WKE1che5PVO
bo648R12Xf+QLYwokmUJMVF6GA/RkP9NihrTj900K5nvgXz1T3PiQtDDzYcKDQI7GUhsDJX4fEi9
R8v0W/TrO/QiPuX1lH8DASb5I4Ol6jIPTWo4fBOEuecCPJnqOQBoStmgf/20sbhCQyXPog5lieKT
+rFQ/7I2yzDmAHM2GcsTZqoYDehn472WYs8Ao3NjgnGOak6o8pGhHMLoMCVLOqeHyJGryRyILZA4
j9HeYFgVd/qWLob4KpzFl1j3LItJT/rdBSBLqyO6UryeJsqgPxQubFUtCO1rDcsKXd6M4lWc6kuM
Mul+wZ6Wb0k0gusBmXtepbvA2tQRJYLWLkxJN9DUDdIi9IlQ4p9oyCrdZX9DPCobmwjBW56RnHI7
3LMpMNsz3bALXvlE0WMigHuLSZmPxdkjAyBdboeI9tjORZ4/DwB9qBI2d+kjIFExpg3+6cfEZ6Fz
z9A4TznZ90lCUu73FdCGP8zz9spYJKLcdkHGo3TsJmONAN8EHijsmcnWTcSltUbtsLrhGseVZ/Sb
pjohzaVsdxKCdiG3N3JimyT/jVJWcUdPvjcBBgIko93b0fBK03Z9/uIrvANmu8v29QdI1pqoYFRl
h+ElnHLvXom0Y4R5khSv/rU2JzTlu2/4KC3IHDCIqR7n8jQddoNzLYDw4oxKCOqDMTMprugdV7z0
gS4yjSryiysRCw5gb9pRCxxD1b2XeToeIcRbmqMKwiNr2b7OX59Zn/ZwPfC39SkD7GI/0wsBzibP
vquyVkiDU8anhliRUC+OBnjkO1zE/Keg6tjSCpdz4yXVxeoGGbRKOaa7mp//s76Gmltdh1Y80RyT
EWqIl+FbNp0+iiUq34y1Wov7HZn/Z9beUAuEdnel+tswZwk6Sq5F/jTz26SNPB9sJhPxTGxLaorP
S+oHIQaS1XCbObCuHNNwy+2z7WGDBpEPSgKvQWWP7LA8Vc6xdAWmvs6T81f9Mko4U2sJhrZKQKvF
SWZ3K0ob2BMdz6KIo9/Wc9GqcTjSOVVFSnfn9a1MvcILDL1JohyrZ/bzirZIDdPp/ZRzAvrY631j
YstqUoqt9FcRdwPC3k6HrHJ5E38xSXuC3e6JaxHsA+dKCDXU8uMP5heiFGGghnENJoAcFe4cjzqF
WVx1aM2hxdCwHWJViqVt/F97iu6sxKHfKTLML1YbwZ/7cG0L70+Gf+LoiymdERi8ohMPNPEutsRc
FK+xWjlWOhmD57kDjTVdzleeIL0uQpHGiO9yjXZCh2px6NtFOQ76s4oz3yA5MavmLqvvR1+N7iSx
kIaU6ZUEqEo6HyN4CKZ6x7UNdXIDmHxZPpbIUTrqSmUpPEsTeYWX1Cq/KpL5pK1go6/bqO2mp1Gs
dDW20fRrIZQZxaKzd/XDrQnabH/BP+Th1W5y7ubwMeW2/6akXQ+DgnIgaqzvanjsPn6JIJDNovWe
sohy8/KBANXTPHCXJLJnAUrrtynl101Koot4HuAYiG5z30CDiI7vpmWbeLWQ5YLoH+6cgpYyxSIl
07vt2DBaOYv8FiKaG9qcO0DLEbFQN/qtQcYzgJhg30+FdkFllhwAp+wZ8o26JrTq+ZwRUrQDa0sl
MdC9NYcsBEwbZOwfdeEp+uZpM6I2zcn56arhm+pYtRZ9C5PqnO7KSqXkiFZtEMIs3noeZjnTlSyJ
/1lJg+5DMHyfDlv0e96HkaUG8NLxJ4D3Kj+r6IDcj+LDDTYzx+2feeru+67d9mxfUt5kHjgXKOht
C0kb3WQro5134AmIHJt5Q9XOtsxcdaNayxoba23WDM54nx1LqxxcyaAZ6chIyoEuy8DgMjDTEKA6
PBi+mi6oPwaLSkdFusLQH3Pa1wOatP74eNOyfyxmDJb+6OtssLNdF0Kas+xWktEW9u5PIGJU/Gq7
rVc426kw2qsIbyii1WUQovpouIV/jsazFvMItpGbdDtnkuTWZicmZXm0wixoSOGpR180OP1Zu+ES
CokcZNicbyfEPMIuLTtinvJH3SNjJVH7Ckc1IaHoH2wp7mc3CzX56lQYTtFaBi5qw7Di63bpB27g
TRVYMlUY2aO9ElzGvNLP6sFzomZPqI4my82TIG4WjqqZ+lUteWfm5aUGrm0dNmPyLszAoAmjGdA+
B2PvBwCQ1D5mVyMKfIDaAKLuWjnDLMy/gHWFTFvNE8Y6H8jPsmYqzb7fVeu+XmrgRUTaxQ0mHN/C
v3QX477CM2WjOcAy+zU9lzgjX2cdnBmaLW7N10a0ZP7NWCjQYmrX6fxEDbgJuQ8C41joGzamE4w1
Zxb4AboyScnDYfA8CPywcVuBl9C+uBvuwN6OHW+4fmrap+stzdsaJ47mIDE4wdfQxBGZY6Qs8Xqr
WeA4IK8jdk2/sz1RNRY75TkLeuSvtl7x6M4ecWd34dVgz4368IrDIZUAgD5rHl4pyL8N6gavhJUP
Y/uvq/ZRMXCOMfHZ5va+eb5nYRg+Bf4WwpxOL+WF9cyPIXLw4nD1aHb5H4cGsWpor1FYsGRV0BRW
aYNSUpx+ezmmVBSGBTVtTe9N7G+q/F1qUrYnf/+x2vsV06rMojA8oS7NmteXnrtA+dW3OKTMDVhF
VIR1tjpxC1m+m4KbNEim+pwwjjW1zC9080s2nt9MIW2t9Y8NqrUiNIso9dEFnZp1fhbXzfZHTq5U
Oaa9gSVhmLvw1UJdOhnlCQYKfXEVdjkQlVz8qar+Y6UoTZfE2xerdqEXnp/jybWHMGTemgfRwxVC
yycNXCU9S8G1sgFUQxmv3J31BnpaI/NrQ6c5FG3tCSIZAZbjk9V+zIr7ZbSuzPbPLokHPrZDPWJ4
D8PZOJZpQa9aZrc0qsGV1D2GKPNfBXJrFpN+klhBjVskrAeg+I9PS6T5N4afgyPAVmF5gXMk3Xem
srR86jydMzmDQH3W51B9bQNWxw8N4Tk178t8O+OhdROCXt4BTS/OuA9TBZuLESDc1E5Bt8hHdFH1
n1BwyZ929NOu9cFitfTgibBf+GCMnAaJx0tC6BeNh80UM9aQS9lBI25I9p3fUCx2jyWCpKMi5mq6
m0ouScQm7Q4+jcu6pso9ndFYtTELrcqc85foHLQqMENvYvZUcCdRfSWhEcgC0V6gLaejQ4tvlqIV
z1UXF7iiv7LkpbtlYnddgpZtsmNaEEaGYvkhqcbGb4jL5XA1qXM6BQZpfSAM7slR8oF4/fVFGsZm
TmRGPXDEQull1GXRk4JPJY0BTpN3lbQw5Xm8lnfqF/gmPPxjYAaUllTqcv2tWTLSfxmZh112sdJ8
dvH+yORaSAUwSm7nm+F/hbVe6x4/aOYiUoKUKpmNIgMexCV2+7Zv8ZNW3z/Yk7fQIa1VEwec416Z
73EBBkzv2jEW6W1GDTjrCjtDDXHBXIA0BUnxziFf7q9k97of4TaFE1lVkA91YfIUx9d769o5piBU
jzNcByc9Yv2FwTqTDCI72MduT7MGBqWUQbJBObuUATDFfozog4NbybI17YCeTW4LMioZXozPZTyQ
1iPTa0opWUctPD3vVI8NwO8Om8zje/Rc9WzAL+DbXufe4XMAK59aXkCshrr0ytVOYxvwPPyeVC97
yPFsUhI1db65E5SUzxkqRHAx7Qx1y9jaNRt1J5i3BXx7CCW9HF9SJ3q69HPo+DZWau3d6raxiL0o
pl52c3OcOda3HLR4Jw3z6+VbQ07XOL47znY82lJpLEG/rWW8qHl01efJs9vkjr4kgb0QceSBTVC3
6SUKMHVx0trHNmdv+YEmsJTrJ7tAMBjtJBN9SBmrtLitBWwiBjtDTHUHtT3gqDQX0Hpb5756Sjr8
DiQ6CRdadSccUjNOTRYa1DognzHwNwLA+OHNpcfb1GblzpFxA0haIeRd/1CD0dWmTBrHKXqUmGhm
Q0BRtaIGSbxV5Ol52rt+1oSVvx9JGfXlJSeBvhUnry11fMMNNGLNV1YBwgeZht4wlDAQXMwoQVAQ
sjWDaU8gcf+YGH+rH1577zltu3m525bVy6JWVc7vveOth6em3+FeYqLXdASLNBIxQeIS09Naer+N
ZnKUVjf6imRQplTw+4E404IjQIzhDJr+nQFS090jISjMbPrzvjUwxHLCQTmstMpkiJhhh0EDtTHR
L1g3vRB0ZuU4vnqcbr353sdyju536KRwrKI1H7CGeASzmRQremx1BZRhSA8SHzScKxC1ILqIHap5
ee4DNZW6JHd5Na+d69cRaf/JXOZv3ymhCMjxkS+kNh2Ldl5yjp5nQMpH2kOS/aFToLKqtRvoC2fk
PEFKW05qfUZ+G4aQW4IUT+ZdvRyjc86uhSXK6qgSimQ49A8hFMFlcO5v7NNSWxnfncft2IYxCDhK
L5JKCDat5Fwa8Q3QqVSHkGw/AZ+xNCO41vkpf8+FG6tsJgayLlTnEYWY8HS/Rn8Bp1Gpciz5zPoi
6pbB9QP1Zvpq4S09tSEGOyS3C4eZw4EI405xuQSZp03z/ctlYWNuWMWXe9U3X2MDc+yaQgEtMG4k
SU43Zed8GyF4wDjCX/RvBIrvWrVbDK4kIy27uGw/gm+SO5qvm3abqAcU69XnwTs8/hJaTg8Kd98X
mhKt4RymokRjkThGg2Qr36HiP1elhQfEKTrSSA8HDU9ESv/VGLtFj+0A+welR3uhILYhpM5eFb7A
eVEJomWTYZBAwDI7ygoJoMriQ3PFKKZU7gJNGharvRUtlYNhreIz9kfkJ0WI33Ty3j9O9W4Bbq2m
5jVHUdpSG8FeMp4F5hGKnZYT4bZVQHIbwMQR3VEcaBBKxVySTNsHilf6cmLjMJkQ2J85wSemdVVc
XtWFJ527ry5wDSTGMWbE8x0KKwkYeUhiYAQxpuCikUuRPcrAcWgD2UOpMLAWbE0HHXyADBsxFdtk
T3iPdhY29G87gzDmRFJA9OCAHUaRec5QaSyODpIDgmt4T099o+mEAo521hO61LoIEhMuKIh5o5Qx
zaVlS2wjfp9cqL6kjSyn+rlA4QcGP+Dd1a2+uA8U/NpOD1EiPG8LK5wNPDHxz72XSOakTqcpwiv9
yumrxdwimdJ1zOfXW7tS+EoMEJ3uXJv7GexR6WlEruHSefWAtFmpTe7V2GtBmo1IipwowTQJhOgB
PRsUGS0TQwB2SA42MfNHf2CoLIwfEIqlwi6k7P8CRqjRRyBJF2CTkIeKNSHsqxSDw1FI5+FGPCLz
nIaEiP0UF+RZi8dB40P1IFMAXB1270rhTeFM4ts7OUAIy8GeWJnnSS83OFMknQPT3nnHCBRCj6+a
QvEWjzTCsAspjzr+/PfdNHOkolqlutC2f+CjB284Y4ojG4J/gbE0T4e9WAxh0gW2GzY2R5WW1Baa
NIpZkBteiOrVzKV6um+hFVV3F/2uKhEq5VISxuus5wNI9kExMtla65zXJ01TyKbNnkIPetrbcMCM
73U263L2PV+8MEMRUy8ciZkJU9HhdbykMY3OcLpczWYlAhB7CnoGo3GIun/Nh2HyBi4njMV3Yn7P
MuCOnJGoaz/oSEMSqcb+Z6DpcoUpeOTJiPYgLDc9pgs4+/wvwOcEQW71FbVhqrMUsP1DwaQC/hc+
ayDyb2WRxj/+tRNNTTFTYB1A4G677T8zhCP9HP2XS/1qtcOMm3+MjXULvpfcLofie5aV9rEJQmQa
9D0cVxXC+Rc/pNNLQ2+1rAdIQYCrDBKKg1dhHRJ8UYNoY1KkrVbWr2cWv0FmqW0IS6idEKsnnoqi
j1ULhgRaivUs2f4eK74tOxhQqEtg8TZAE5sGrDdcrZFAHTRQqwWM/RfwG+03QRv9Qmn9HPy+fU7q
clzo71s5bIlQ7lCz79fqUrqUhfCMuk85APDnROEXNWC1zQ4fNRWCNaUFvDXVgWehiQ0Ox4c99Gsw
f1zj68R9G/PHZpljImdUnyh3cQFu2KmDRbe7Mf5R4naTQveyhfDYrIuwAQk3R84lKNEL4/nf8VOf
x9RYR+KPqEn4fdeXmc92So1TxS7Avb6b9yOpo8YeiHEkXOpT3Km1qBZfQW9q9Jw9l2mgRklTu7Z1
RTiqSEQHb4CoGJHqEHDIkFecck7fmEJROxAzFuXYbpGYpiKMT6o9vYYOswrE9IUJmNjsNnsBtuFC
xMZqVnJ7p+UZ4d4B0ZMfuC/2lmpld+H3JZb3fvaBjj0qtnvgljjyWg8W06KDiOIHnpBe3Hpk+Dmn
7oWM1Yc8DXa0foaDzLEUDTOKYMG5MRDZ6v5MtXq1FovVTN4o3ITPzwC4NMHtkYSEE5x1VQdYBYZI
wX3aDLxoU6PhvsiXG03PdGwrKqzUkh2R7L6oiOsQsa3kNys1d5qtUb3BKGxmJlrzIjZ7GIkovS0d
FIHvEp4wSiu+wytzjfO03iJPEmwY4DKhtUOOdGMQzPQYtn9xcmSKFxdief872XL+ZsIU+DgGPOCK
R9PHGbwf0N7sII3/GZ1sgaIYuMXRkTYKpM9l0KiNw8V33pR0usuXx6i4yQWXjp6FEdt/oW3Qi/R8
mzDoe4AcoptOGoGhnlhgTa1SB2dEI/xKC4a3U4jJdD3Y3xdnD62xRDT+gca3jNkBcGqFT3jAkwSP
k+h8pAFriU3NYPAO3zt9poDXas+s92TNn0My8L8kdCCkSiT0uXMPQM1mvWtB1mwx+O+3Lgp/j2cu
j5N48rI2E/NCSL2j6Nw1WV4FYZM7qVE+R1KYROgA+woj1XZhRPjn7acxY5VGgXK/huElO0/yWF8k
QkQmNqVjFJc844NHevxVlLKSK8yoOkHGRrdwuJmao4GCwNvVPs8OzdKsDOPNdy4SSND629Pp1QZ/
pzn+6iu3DyDifN0KZZZqzeq8LVrc1YKJRQwMo0vo1Nx8/hk7d9bvovjZyuwgyqHs05fq8nq5kuXB
gJn2fcTVeloCj+hAqhhRlOtCqC+r8oMrP8xeGmqh5L0r9VmSMprk6Sffn0ymPXk5vRjQOb7e9tmX
a6Lp5tgKuVRO1hxdGEZETw9uKtrmMVjOkk1LBT6YlLT6pB0iVdU+rmOi67MHO4NkZYOGVxIaAv23
oVB2bs3l67gnBAbWZwzr9JMKymcbnjvLunjnGQ96EFgpaBPvtAhruRZ/l3JdKDAUZnXEjpHk30At
dBiIlpjkStDdsV3+UJthFSOfl4cvwKeDvwfFS5WgEeu4EUjx1wB2ad6WAUb6Ebdrd9OOovOqMxBY
HXJqbeOlmtZmmAoV9MjZAFMqWjd4GGTO3kZlLP22SAtroMCh/cYOPOK9uvomy9XQDYxvX394bned
KEteBbtWwoEtrl/OC24r8qYma/Koqqf4ZJHdNjf204RRPhT3B6mMYLqjybhKHkuJkOQ2X02CSSPC
w+rJEkeTXE0s8z17O7kF9jUIydE0mLgNbAqBvdwHmQUQ+cyJVnc9FUFI8874LQcVsbCb3QiatqcY
vwO4TP8nfz1+Wemz+QpBJldepIf//E2JMIdkXpR8AsMQ1rdeZaduujdXunSFYqQp15SuBwriUoGZ
TqDRlQjWOlt1b+4b7VDYXMOLa81NqvfoTYl8/y06MgmOQpoia3Rdn/lxnZ+QTEYrL2WjvdCCQXtj
MY7uCWh08CjcnaAXvRExPGBkYQ1q+1sn4MVoBums3TEMHAB8DxdJhjVlWEnPS5COotNn87KTdKgg
AyesKF56VnAatsUYPgDwd38U6l+yOz2B91eWTIZRaVlaYnubl+NspA97HcO0Ioa/j8RjUj/fIx/W
F2HfX5J4hNSg3HRwruG60hi9nNITEN93ft5SzWe9lDI+b+OaYWRnS45CuD310ZB/5jOEk0k/6B8T
NlKEEQmOzAYuIQFIrboW9pB6HdGtDYrRU5hqxICfhBooyWlVxyElnNtTjF8uK0Xtp7x9EKRPPJEY
N1hGGYN6krHVRj7z0GQoousnmOpsc8q0Pk9oWjJvK4YdKKBsiP3dkmIFR+vpdWCfVGvfr0srBRqV
mVX0B4nGhBJV7mCDj68XcrnIXpI0kvnmBKEpAZlflKmgDkAbJsfN12hzgRjW8JOxq3JbauM0Vh1+
Y6ol1IXyYhGtwHWsD9FP68CxiW1mdUR8R4iNQFv9Q7z4rGQZjzzuQ0VS2Ug2L6AMBlSmFgOXvg+q
O8FmW+vI9k10sVHrWytX0ppJKUrZL9l4pAHRMK2Z8Wuw0d5iFyABxSpz/IetrPjThBm5Lf+SEp9L
AXinl8fyZeJrszTnUPBwssoVMPoWr+8brUqXieMegqFEwfIjg1ZhNyFusq4xM9NK0wsFGN+a4z9f
eztcW8KAuF7BOjg817MncTVZ1wRaZAd1+zrJUpR5hDnxLUQAyz0nsfI0tGcTDYYm25tBydB3mYDL
AkG6CuM2WwWnRyaMGuPt2xFn7LUqQgH6idYMzmEjuC0egTVJnLg7LsAmch06XqXuTIn2vKEjhSdJ
AWUkXf4AD1sNA/zJUAtkFcIwJJiCNJmLltTdYHcO/9EODD+yXtZwYyC13qawonAJmf3stt5hCZlo
CmzMiTKfiSZlxnh41p8d3XvpUoLj/VmIoB0is1V7N7TvTYDHx3ORntDhlzcd0ohvX+nKoFGWIwN2
3rkrzin+nDrAJeaTUriQog5lBp2Sp+fA+qHBpoVk7VFEb7I8/CemNplSy5329nNtsh3cUAywXN8U
ksTGVQjuUqn6sUzwWQLMYI8xwRdFl0uEZ+OB2HgTVhYOG4PTTAmfrtcpdXQhKE6Fgeqzo4ehFcXd
GDJwK2gP54QNFSgpml7fAXGy51pGA7YPobgj7msHEIhzibXuyxTOwC9ccepfrg0nNkae8+gxFK8D
L7U/IyOYr1/JEhzLTqDx38DCBFRz/PzkfSUPd5qOWGk4SHTauCjoeSr7BDrBsxAihZ7CjNPHTMi5
LleCwDo03dHMf6t+qzpCcgtHE3lD8BIe8VrFlEi5zQdusvi5Ppbbnvg8hGrCJjzQwHLrpUW0cnRl
91zaYpAIAFLvrmt7S3XCpRgfPFoHrb/1vgHDd9CZ/Hr2r+vnnRlT6qduS39E+hQQN4p1FzC6riy3
DGZzasjx6Vd7PgH6UptiJfSDQ1ca6GQVA+0gsdKwZGw71wjA1L703YazDn0AmAk2k7vW8ueXPxKR
xiDGTpvlLSsyMJUMjorNYnjjp1Q1G3rQYDYEzEMse7lEz1SBH72ExmpmJ9YswTdlOx2/dOUFQzqr
9D/WbuocnJJFhAUiW4wYZWtM1qCt/MgFKBzHYTIyeujdz/qY4QzHQGsQzh7prn672fA7argzTzvC
QJu9403xDk3Ce8zURvq7rAeRo+wqdz43BD6FWNT9xBf4pGXW6RnI9NbJt/pmFrqJSgMr9aIh2f6t
lK6nFiILpnVH+0nSnFENUqzhMwdfeNtgD1pZ6aYgZ9ZJRPtEM12rRt6Lqe6gl2i5no7/blwHMmq2
UjhhgiKNK2VGuDTM4Qpc6XkQYvXaaf4BYQ/JLa1pALpDtcX+yMpUV6Yj6mqcoCJOz08bODWgr4sI
FEShuEOLULdQ4PiA85j+e4YKkWvnLxc3NKlyWBZbs4tst3UPKpiU3LRoFUNXM/jhBZxS9terr25e
d42+pkdflA0GfaZifvZ7BRvxGwKjPwFFMs7Nn4pgNROqOZLpSDn/68VWv3920/d9dk4LxJicYX72
EzLCETgX52WXeMGd9vDU7HuYiqweOJrIQko1BC+ktW8wugfKqXECIeMr8nVBtpz2lKLYFLXOp2nU
22+FdKQTqj1SGnTDwXGuIRQ3z3fCKWbo9ezLh6XwyCssOJctVjhKDhP4xLL7e9+SsnxhIiB0ICu7
WDlUU8sC3lglEtNHOwLT8+NOgfIBsPuvzPmvy/c+z8OCNatEiC80xVrtcwewJR4J3HVeGNZH0xfy
jBh/TIEQzOtPzKOrm69YOEoOmzDHGIaflXzVyLmfC8YrwzSWI6aZXR57PbB4fP2ydWM1P74ZCjrg
U/ipyiMjLMyTAdTkotzItW+argCo/vCOGi+khpHO3c1KChjH0efWWal23ZBSeUdYMsgBXWxGIO+g
nnJDl1FFbRqb9qNS5y4KbRK8CA+Q+aM88EJykSPzmBHyad2JyCFrqU7JRpfnzfowe2+CeORSNsCU
r+O2m8OmmdIY1BROibCx7blVNI7mwSn/X07PyRUY67nN+0hA/UN3TPPHghXiupFsVS8vUSnR2Cp+
Knh1hXbs1kmP0H+iz3OAidNq66yXGAHo/AkIdfDN35KXy6B0yRhUmgd/DmyzzeA1ev2IfKnhgGgE
KUrQxxLa0hvBhF6gKWfsmVqo02Dq+IG8gEvtkhvVCw1hDSV0a+wBFgO2bgFFv9Qs09jAwlNT9ySc
nlUjlhIjqipn0iw/UNhvBXx+MksFqleDxeJ68Gx7AZYlhnnILL4U1cIDC0/y781etN63rw7Unzko
BCWghV0f/IcET3+mC8PtW/L6zkI6ZdHZBV+GoBpXo20maT85ZLaYYQgraND7VOuxBBRQNswU4zal
M+Yrtf6CrCL41nPAn5cK/el/Nup9evsknPhhJWE+n8Ga1my0dc7mZRwxgMGsUfiLijjv+B2c+ASd
4ru/mPpb0gFnxX5zY8hKkgzjCdVde233tKd4KnQn+YRAzKFPODIvrCyTG+/ihEKihhPO5UUVqH/m
ZtbuOvZagVAGVjS/+/pS59NymD9Z92eNydEmYKm6P70AOtlQrqbTlOjlYTXOAFKjv9JeC+brEQ5n
VOEr8aFf9T++eIZDTaV5RnPFwuspCEC1D8v6nhjYTsGEObKYguKVFcu99MtzKpnBs942DPgzwHcR
iWqYaU9z+F1xQr26VDP2l2DJ3UlmH6/SDhajxE+CXXvjeliM1tRfPuGPtgQ5FK7OczGfJgpuN1um
Bvn6STIT5Sn1CSOUozGAMytKK19C1BwO1ByTde9LTWOR+og33TwEK65JjLk5MlJ/UYbOVgoTrJhh
5IHB0goE0AHtNCGGs6CbZ+Zc6Xj/9XKGLfUnsf6jSuYNjK8PL4IRjG3ooZElwki6Y+Sao25MoB8r
yMUdZl50iFXdQm1MCkBlc9gFHEZPjW8I8MfQbqbwx5vVhtFWGZMY6/fIb7vx+chlfwX1OQ29i+GP
QkpAjlgeWZS1T+HmXVzm0MJ5ZhdZl41Q6hzzXlQKiwnUhs3+MCaE7+FUAzAyWKhUccTIhipHnF1B
JLr25MYDbWoABtLa/y7TDcs48mVScKQpEFS7aTiGCanEleRH/OmMfWXHG+Y7sVI9ep0eLu786UsC
PLfrcNLyBj+Q/yMKQkwx6BV9DAsd3gFUpVzKbqUY6GZJWutgyOKmh9Kz6m5MJPRUNQxwjxY1iKe5
BySbpHRumlCh0Vm5wG4FSiPauP4V9nC6s5sVG/6iRbadzzhQpZxGUjTjuNtsJzQbQnpktoPjz4v/
M9gDy3mNzyOgtBoADBNhApE4/Ej82XAmHOm/qF90afE87FDcI7Z3VmFyvg1QXjgKj0FxCe+LemJr
9Az+8dN7rrITFazvFTRZ4HBeFrBZg5cWNX94I7mEL2S5g7Ao15ZdY9dUyrP6lKdawG3UX4wDBT7d
W8zCuEeVW9xdiLqub6MBrC5XkOUDWhKjJb6+t99HCqDZXxxZSQkc0C3WDgX9zOd3lRoyyJDz59dV
UxFyf1/iwOuM/8mAnk5wxQLxDRNdm85iCFte01q5tjlHsS9XSWzFr0uGMfZkk6LMmpJWFhsdWsEu
FhJB0ZD/zm3fRUA18k82f+HPwdsWtyHU3g6JET49wCxkRjStLk7U2Z8Ht4uo/a9LeZezxkiycKMc
fH5+Hp6g1P/ujJs9M/GN2yAgVMiKqO6+pQ1SS5lzbgHiTWCTvfMYMQ7MuEgfhoOL42nntXbwmm7C
dRpKwj3mWzzUFMwRSm+ijanOAJR0AN3iVuq8YG7UbD0C3jYEL4oKrzPW5zTWOoswR343sY7QPYD9
sjzOTfjTZLJFhha50Ijg8CWk0xPamAHoo/P9GJfmN8Up1nMqCaIP/DarWpKT/Qug5/kzBdhuE58C
Z7M4nInTSTC/wnKMqw8PupX13PzRNffGjnGTA0pS7AAK+H3EcGE+292SbY8HgDJD4vtjBgQ6IvZX
TUMPqFcV8uXXYUP1y3w/GF95RGSQO33TWLjQRGDudekmGC1V2axKQW9+ePaC9xDd0X+grw6OzWc+
nsdPRQyY2XYVo2jbDto+h9SiMhzggx3+gKBEvj8CTR54ORSfyuZMTVcoVfJ13iZo88f1bSIkTYn4
pYUW8n+yoc1jHBeKxKdaREAPTXcCQ7jfzVH9lD3rTzxpwh5OCBnSugvt6ISEqS0ULegBVhlrUUDr
j2990zvK8MQtTseteDyaKUNeKqWzGke0+ETbmANlOGpgPkOXfefEM29vJ1gkdbV7Sb3B5uvkn3eb
xd4Qli9lui/tLNBqo+6KkHqD4J29MGfvRhHpkNrVw62+SY2wE0oPfynOwyoR4GgoZCk5w+/i4rsZ
L65BoVCKH4D1PxnqkuK6t+LzEIKw920nxLjJy2gngRm2PhyzAz+KsX0Phq9EdCBMMM8fH+Lt6Gez
JZlGS0AQClS/ztb2PeeKPechBUQbRj3O7RaVVLtJaZXhrB/Xk4i3/np7gOcG36R347nsfqP+UDn4
67f3J5VLEhjC1FcSJ+mWrI3rfEFvN2WuXA5NNKcZdyWBFjr/msvZh3m2hxJTHwnyKFxTC57h4Pne
KaeKw6gQFEmUMiju+xD4ZSmlyJiFpdhRApPGKPKkfIr5DtcnCKfQTj6i/hGXl9RQPTmkFibk5pLJ
QERbM6tekDaroy/y5130vNdC0UEba0J0bdjNJRxdR8/O7yNYhEq8Ciroueui6HdcJ44NkhRjP8O6
gv3zr8tcW1ucL5Oj/b+PHxRsnEL3m/bevNk+38/gP7FmHkOhce/iIW3TJRiNPOsjZmldhDfQPpR1
cDjLQuGbfBjTMOZk851jleAW5/c45F7/R/TMBkhUrFdnYWr1nABEBA4bEM8YSa8c+FgP9ACid/X9
iNTK5y5OJCkXpXN2EvWGzlq/Mm4UjA8EeZkbQn6zJ5imdEK2RHfKDTD0MEbMiEpN3benBU5mUhJW
KkYWkvW3L8KbUcoEGwpnGKMq1XoUth/xTSuijKWBuCbob3jytnc6g/VQpN9YZFbrFV6cZfaN529V
NBv6D181whlNIurgFuSB9kYda29D+fOvxkiYuAtRhI3PQcQZX+naGZwuU+VPlEI9oare1AeWyomh
DGXdV+lSrmgVm3ayjjda1V2k/l5G/9fxKyWStooFqNVn7XyDpsjU8UvZG+wUnjJVfl3x9G2F3RhG
EFylkWvMCwvYEe7MG5gfyZxAFnAx0dT4Sj2FUIKRSZhRCo6OnNVPqnOBnKS0xTtVckyqQtXQ//Dv
BcTLwv/jDciiGsF/YZCwBzPQsFYDogyDjgsFGE8kjWpQok3j0xT6DMS0Q8WTDKUD8lyXuD3d/c+7
A3Umgh0j4O0Lrwcl/CClIXrYc+u8a0m9SpVCI0p3AM8slElnxE85YH61DIpK+/j5KDEld/XfyjeA
N23ge6M9T/Us1xyCEsf+bamjz4FZJzlWIwx59xfGMAWETtG5iT3eSEO5ICxktqE2El34oo6bSgYS
QJXlO8/gdH8Ve4imNgaVPxn2pJ/eqvRvvRiAiC6uoPOr4cQ9lh+QPPfda/6EyyfgzTad75LkVUCn
40ttUTvfu/PFFf7btzfsG05Kyie6/4noy2AxdRiO4l93+b9CHwerTBAguw0ZWpuL+lJ6515OfTm5
87/ZQWX2YbopQnVUTVCU7GEOwV8vnvoGChxywh+c1Ix95c6k3TjEIw2fnAL1B4cZbxO2fIOOfBh6
DmTYcQy+Zme4nrbrKgFhejxL2oeSHHlX2yS2boqtVd4ZhcHIHC254Kso6j7dtSNAzzeJib+RZphG
UUVT51yXRlreSA8wuPrKDVgqU7tfTp0LQVGOgHGodfeLM6q7sZfRVeQuvA5glPA7EXWMvOOmKMCu
TAacmsmLgh4Gmuz+o6hrA+CXk7DUyixNmMAY5UHjmPYELh4VlT+tDqo6FmR7L72fGDA5hNfQPT+x
uBK/tLTaK+u7Phey4zB3i9mfig8RjmFh5CQO5jgCWOrb9KDCSqhbEP8/LxMZbGUawZY4imGaytPf
bDJKhLjHKX/RmPmqNGeGWtesQ7R6rwWmqEeXiGcNoxYQpR/GdcY7EYK/phu4aLYIl9HoDyKnlf1+
mzgveDitjnI8uJnUtEWqc7y+BvBWFjsL2waBdnssAJThqR9xR68HFHxqIbY1whl9mj23TMAILAb2
i6w7Xx2birTb0iQGYSRFnBBdUGimj3BA8LxBbZdezFTN5sVhiR5f0W3Nzck6zDkfJFLO5wheTGDP
yXc2JpNvdXq1ehPZtVtj0ik4hcPDKnQ66qAmDetfvrcUBe37WI6Mq/mmn0D3lJHXGrubs8TlCjcn
MTB4SZyqQoGgG0T/Vw5DiO5C9YjSMZs4imvdRUTNaX5N9NjsgVen4THiNDu8Zl4f2UIZ1E5enWBD
Rs3igRZxrjZpKc+T+2L1bjVO4SGUB+QzKa6EBspzUCqj1Y2lsj1+kQ03OwVZlU7DvqqcnyLB5ScS
0YCXJlx1vizlLFrLPAbQYsCG6b8Yym/KzYj6w59wH9MDWfqi3UQ5TK1nVjJiR3+lfKDIGMh/6bge
wyvWWuOUjsiM06jM3U6h6lImMzwC0XviZsNjqt7nXcJKSvRNHcTE3Bd5eg39Wx+QySKnRYTb+5In
TFfYCCH8rtfuglXetPXd2sXyYdq7gViz6IkusrW1zNJT0HfRLQdBVGyvmwHAMq7GMpCkvLNo4I1i
9tJ/TdcpZdlWmVPTN5iEf0mZ8v45qOAkNpAU3BQfqWEWm+EYz/Fl4Gyy98fvZekgPEU2AjLuYTMp
HjnlAu0z1noKMNmOeyBPkFiCGmCCMrwB0aijo7sci9L4uzLwjSjuMsPmZUXkZVsXCbW0O+w7dgUf
47GlP3k/l4q/wdJy1KO85hVkEPaDMpigcQXJdrPo1HZ6Ya2Vk3OzVqmtxHP40o3Ozdssg0Bo32rs
1lKlcMm6Oiru6WenMi8kFqzHldEmuGkrEpGbk2FvV3qu0J5U7niGzZvI64eRCracCYw7C67oqsWO
dmmDZogc0iMTjlEgFieMlvBhXE4//LUtHaG/f6uel7xMNDg+PPaa3DB3QOKMDLcBP4/kpcun670A
ilgbJH69tJYSriRxetrkvBeYtpqw+5YcMm0heKed6zi2XVxp0W8G1VD/O0I/DNnzFRirRE8XAQwt
ex+WKn2zV0p9rDmVGAdudPBFKQzgerw/PJdnAsj+s1Bu9potLtc9rLz3OHtvEyr6l2QcOLb+FC8X
7EvZtNWTKzHBvvNuMcwenUnQIbTFo/mLkxOPojdIKTRBhW8JG6uzjmfDoL0vUh2RLfBhS4H2D4u4
4tjkvBHmRbwGMiYvz2tOslEooDZq+Yhdqy70gPdxzp4AYVbCBfltHaSibqzrID+xQ2lsjLH7RA6t
4rc5ZoUkCvwvLyn2Uk/WuXK4NhbXeOKs+7EcV4SE7QCB4FI1tsAAbGvZMS7DbUqxUJtLr/ss7i80
IGvy89h1kX4aC5W9iVrF0a6lntjsLt3oxwc5rHrA4WXXxQsubSxayeUkYZNCYWFk7AnP12MB0qj0
2xsVWtTbfUQZZ7O+nuLsoFWmGxdPCvV+an2SQQvNXtGnLqVmJ1Uy6qqhNB5pVwrfJcRriX7FMPH3
EZ2cjDwNsFykyMFtcW1YLgTiGPkyXrBYfhSB0cronnVErQvb9c6tV0YK5tyLSeeJ+gnboZAqVRbW
2FI8XmeCkFoMLRKlEg2srib/HnipRioJ+nSmCMEuNzu86JEaq06dW4qJW7n+yLdGCu9/ObBdOruh
NDSKYheyfVPgSLYhbbTDP7+iI//OFvhYPj7rbdR9PicBZhCAxxshlG0P6iltAdf+w9VJafJxnytz
FG3rfmZRoBUefJYTDpXd3+SslYyIPmzxW3k4rW7nZl5g9AQ4AcJfNl18yMntMkwXr7eM7ERkUFBw
Y+VTSGCqhyaA8BIM0VX/WewkDTv51xJMxTtmVTetBs9aqRfk54R+KPdn3MNygw5jyFon474KSiNE
endCtT7rc5NlyiAmBiwse1XWfC6e2vOo4nowKIK6/vn+q+sPu6Z/yGn4+j6xayR1YIZJbFfaKFs3
FTUUsedjmXyqgr1BDdQzlHr2MeXJ9LTCMi/aDlybCfm3M9H9BQjrAB41O9ZHB6wQ5BFrH/bh+MH3
lqQHr9oNSBXWpnVoFeT6BsrVmElee/ZFEhpy9rhFhpUpvvoW+NLcSsqc1DiPOHWyo1ASddd+DBo5
iGc6JOdAdFZIiTTGc65jkdlsZPzeoELTdA/W8ORSChfcZqtb/t+oNFj9op2e+dY1j8j4fs1+lnPl
QYR0IvIvNJY0pgJZe41akBSmtQEvO2sLDc3Jm5Y1VslMJ1yviHNJQZs+pSOVObdpFXIJPUwE1b6M
iEVU4O36Kt449t9hZ14rNZDcEvXdDMMKNth85FUpM1iqzLi1CGml9R09Ba+rD+olDL67GTjRXcyJ
ug0elRbyuTkwweFhgbLADz3hViI0MDTarhWvz72FhRXRUa8IU4kERhug2BA93K8XuUkN5jgLJzsz
cUvxbsh55T26QGoNJl6DRjYw0tRi6MOCASPuytjyKnbQNPW9P3bf3uGX5On302RIkCMR5FkEKAgK
KhKdlnVm+C4KTI1RmXZlTm9yrWIP6Gio10avagu6KFhnvoCSJe8yoket60W/qnGR79EF0M4n84RW
OesAmnDdkb4BhG2ht5aHoc2cm0l73+PFz8tMuqqXNMtcM+PAEzGtiXFfrRqRAVs46e2bL7yDRzG1
v2SOHI+xIXCM2ZglrqgDCpwo8WWdKA7vGZPVcV2gBArmxApTlcqzUuQzAiPlKYaHWG0hYus5KX3T
2lkwWV/pIvJ5b0J2+hy6JadM55y4ifxSmX6p6rxkagaqY8PVvgVunMhrHVpr6mfibu1EA9/h4iYZ
mDDaxwbL+LnD/upWjjkGYTXMWafQYAMP0IBHX8nIozpHXhvbwSK6W5HhUe/cO0OuHvJfrfpxi8yI
+3J6AlR1jCLWv8N1iO5ryvZzO/S7bsLAWFdJsnJrBo8NZx9TULCMP+8xKEKWtghqTraB6RgbYvwF
d0YjihDO5j1Ur38dklQN97zf95FQkeCj9Tgap66uFkHS6nkJnm9Odnwdh2Z12gdCsgLRItvhworj
8OAYjD4+bs6VBIt3CnqiJKYHHwfeuMOxr0RD0vOMbt+0v13NAxl4C7c9AqG0J6rIeoisiKJOY9XW
HVfkUXLCyPo+PX36pQbcc5lgrhqNSaqeOD+qRvB1nhxxLK+zhJgG0sbmSZ6jlmtKMiURfyseX9DY
LErkLiz3je17snn1MbeaDm6kdvb0LDB/uc11ABSDA1eUmSxFu17gpQaBHWVOfgwv2TMMVdfODskn
AWYYRyRkMVL7WCogFlx90nrUkWb0qmZleEj59iBjIiHlS+QWV1wTTmRIRo/pAkmU7pG94egxO258
d/4Z8+vbm2p9ED2bwyZyHKgbtDsNvc0e6+jYkP5zJmxRUQ04ig0cTN1QA+aDnFLnFk0b8ysn6qUk
tPmvO1DAZoAJ/IJ+bSai9YYeiMTL0w1E0y4CbnTWH/2BlZ/GOfoznYtyM+D9MNantFfSUTqLjQ0C
F8lpSDn3ykQ6hZP0t2XACTS09Eb+EL3AR7LPMfsBRL7lCBYIDfgTFPfyh9mVbViCCLYRH/aQysy2
zQsL9aXKD3TsMIEvcjTIM0pGcx26iMpSm6xMCscOos8JtlucbziMwWQhx6qKLrZiabhnneCvGQpv
Z3iiO2rLeeeSsKQZuyA3WjkDzaINP1I62Hj4ewQHghPNgQL/nk4WdYhPNF4mrZS+as1wTuOlMQ4W
NCB9r+xH3HDnAbJzJmkW7z2yRNYpmOFiYAWzIED8bfaGHuomAfGH3eGIhh22WA3T5oFV5+GVJZuE
Zl2GPWtoPhwhyexTT7nDASi2a54vQtyrDoYaIgBIQWWgpWGz46pRjAFNfAbYC6suBQuQFN3mE1VI
Y/BSlaPdmpnL/l0KXBKwjooaCQGi/RzUwQS5LAGApEgBrTBQ93V3u+Z3BCa0ll381OAPWQ+8Q9IV
EJyN8HUhIeIXhU3yiR3jQZPUDbERXO5WCHEFwQiiaasnua1dk20UehFTonDHftGPiH5XgkFHSeHK
11AaYr77bEy3f5A3/svFpI3l2yQKyj6YiItPeSxcOfqFad/WokRGeEUPupP4+52jeWSHd6DaclhV
ydEzNAWWmuf+Ct/Iwu7Zr/VaHge+ionwybywZnPUhEOOHPYxakTo3Ks4VLS3O41j5bbvOBZ5iH0a
rW5T67Hl+OA1wU1i7nldMf8C9Q3Tbphx+H3DV1AUpuSvXz+RxOOkj8vk4AudYMRLfOQS4Svd7y17
0s3r/74a04QhMfdD7tkJ4xOsDEEwrFKjs3jfuNjR/zWVQU7P1/499/vIACzSumqyz8+dToiN1e1Z
ZhDFAZ297+30cdIEuBcUQ7Ahk4oGYs6zLrkxUPyAWZ/uCfMYS2Ux2njIgQygqQU5dBinswhly35H
z0qrEtR1f1q20Jl5QnmG1Qi78im2oq000V4zY3t1+6BBmEsyyvEzAfGLtGBQje+Yx4VfDpg20sKk
+qlkDaJljgezcAChp2lMpf0asFrmnLWb8Umxbhu2NEVnEdPS9kbZYc3AUzSmX2GnsbEmXNld3zq4
LlFmriTpq8XKwqcVIa5CJY2/qAfVZ9LgpkIrEXSveEWaRQcaI/PnF63AHrDo9MnU/zakYnGds4yo
d/5nntL5RIpjEPVzhsw54pg4Ppe8kizWS0ko3dPW1I7/6fOKA4GzPufx4fE9jJirELHopxSXVb4Z
DzfNnSn46s5uwmO4pqSNSgKtDwsvbFcLtXFGdMMyBJVtC4jEuzQyUX2H8+xPGhoJKKpK7wXQqMJn
IwaoCogocO9UZaPrI4xSBJDc7R2PHk6RQFGXqCNI+fxColnyP4foq1h9eUQwDxz6ys7RyXB3Boeq
+xmUEFMQFbTkMLhkAeMtW0hW3KvlA4vRF5KsK0t9kNDZRvW5OEgSxuR75z7qqx0xlII4dv5C9fM9
MTK73W3bk1x0p6J3pnLT6kppgDN71VfapevCBHJKwn2k3MLdWhELXxg/K/YZ5UQRPlNe14VI4E42
PkISxC5BBqL8zwdZhrhFTnoEPI7vyuHY0iXXdqDVuNGFC/A89nY7xy17nbC9huvvY+wt8wuwa61J
1b7akO2hCc0wl+bgyqYqhQyFkoVlMOeM6ypeD50FIMzERRcV2PfA7p1tKnNMAwKXos+SqOhRfddk
rqsgPTJzePdr2KiyLt6xDbfpFFTcllkymskhIT9HTwaMA0duUArnA2YLmaSIzXNGxMwRd1D3+VTY
5axjW333qkydM8HYKmBsZsCxX9KnOjwVivxCxQdwNHYKlqehkMjjKyuf5Y5rXyC7CE0++37weuX7
Vz2fD7hxW737pjA1gpC7OvN6b8nEs3vk4+KkyUazBGx6NqR2RugNzTOfIKKAtPZiO1/XMQ1I0VYS
H+A0U1kfLuEQ5u7qpRJkWlKruVW5gs5XBlGQOmHx8UhbvFKlC58M8xfTDD3sbR6o+reuR8T8RjzV
XXScaXnLs+VAFr8MXmDsWmb/E4AkjRn+0qef7Ysihz+IJrLTGW0NRlMKI3MPp/jCKvwQeEje/oxl
ibaXVr+96zkG+GNFw96ndR2TOl1MNCUxPVhu6LX//c+pfE4er7h/4hnc43QX3D3kOtzfvLrsCdNZ
3rHfl1nqa9YIbxUt9jlNV6sDAM6oODHyuidY/N6oT2wrdiUMY7Geb7Ce3KQIHVmFF+Mr+R80L6+P
kWvMXXG+Z3jCgLh1JnacWzsvJWebE7dMr0JdFfIQkGM3hWYxLc4hPcGIRNGxha+UbWkQNMw+4eMp
Qqgjn4FNuiMP2p9VPiIAHqGpIVUnpCVyFJ9MGzT4rFei6wxgaGxShc7aKdVQvVnMtZgHao24LbjT
7jTgKJGdivIVzt71cU9kqEvjxDCiUmT5gMeh0D9O/n30Lvbl7PEZG3UxvL4N0lOm82L/8T7KVOdc
OXVlis+L9DRTDueaipBJJqnt1JhnTqKluh0zJsNBGXHWEp2M95xL3Z7RqRrz8JSBdByh2LfFRYrF
0dmkKt/irzjUpCNazl5T9UUWuTruVhU2gN1SqusPHIeN6Gl/cN2cZMuzSrjsNkKGJYZYZAuktLhC
TfgT9ql1DXwO50RlPKpQVo9cUq7PaIYsXU9TAbdcOdVMHa4N2TLPDAx2O4+7EKRdeB1V4vq8RXwg
EaB8k6se47svt7wRSz8rMIT+9eG2pALmEdRZ4Nuiu2g12DpbxxX3k9h7zzwJg/cbH05gQu/KBfNS
ARCKcIPYfGtFvKDnpECIqma4GP0IkAwC9P9STmXRqvxxdnISBQoTUe35EodjCUaZCwbiMpN9q+70
UXtyQYm0nq66M4l8RzeR7ZWt2Ntrq3QoR0WuSMmi05Emwgbo4NbWhjncVWos4hS8Q+u4i4+Hqs6A
r5sjaG9lO+DIMV5Knd+VL5P+vLnEXk2Elrwg2kDI0nNyV8yYw9BgglP2YSDgtbF2l7q+h3VNkb+B
h+ZHUAmhnbkKL2ZcwpbM76LRmzGfTBWeY3R+x2Z9eRQs/y0URSwpxkSJWDv0BbkyjU9+oML4dy6I
OhCXDp/43JA7dqIu7aG5UyZR+NexgH9Cc2IpugtP7Bb+Vl4cnq/QxoJ3QlGlIoMED+S5JUKd2n6K
BBcVzEbPD5FuTJCzB65xb+XwSAYcJm6I4wtAFnp5EWReWjAyisykRMVEIP9Ukw/tsYutQEe2pnpX
DCMYuBv47smx8YPcqeiJO2N+69zKnh+LmBxSgaNt+12mH57ePw7PehUTj6DiwNDr8KbXnmbU8IuB
vcDVJfPqHoLVQqlxsD3jE6qvHsRAXuXabsS9MTF+u3RK1PT18tli1BJuIzafgWM1GPMrZZjYPOXX
vfmNWDTd5YuHwQFckOFvVHb2Phj+8Vh05p1FpiPbr2GtlwWzPftG+FqkE4c2Ep2GDRv234m0yWvd
vMydbClZzbTsvj+ptTVkMa7TGJGeK78k3FwaPUWtQSjNHBAbYHEKkK/dt0QQcJjBwq+8BP9H6pMm
EarsdaXDp0fCEbd+V2lfLyppGVX8qmsJIXmEs1PVBZhqkSAtQ3GLBdjPmZivHz8t7U5s5mOmZHDd
FmWe9kjNsGJE+3O6BEnt9g8hKNd5rFcwBe18PbflzIY79u0HfuYgf64KMO1yquM5ha+ge6ww53lB
UhrqAbwVdznXe9kRTPB1+QYazN46iSUxHJNBgY0XG4lTDEjoZc1i5YEcBsvX1FjiiDN88KvUqqmb
Fh5qd5Vm5b2hidrPE965hEtnWJmv0o+ZHLNd5rlxYRgVkxF603RxBN3Meh8LyEb0VUWSSQlyPKlF
XBWHLdjWbeP/zntVhcah7M8VVhKpw7Us80K0O0YWg3e/MJqigsIaQjTIyVYj8c6GJk9jme/Izbfk
pwL6w1Iw0P90vUkxnZCTpjFosrkxVmwhQLxYq/Ow6e//sm7Z6VV8DFEuSnNOHV03OHk4exS0PQcG
GRc2xlRL3/rSWMic1hRVulvs4X05WXyfYEIHKEW149cJRFCv6f0Z45X0IazPjuTvkUTCnt3fgkPd
R66EqKRA5uf4iqbOG/ce0J5DBzvrpDRaYHsi03JtnUT+0BnU9T3kPFkIvbh6c+R6pg/jcWv0o9R/
rWT12ukpsmklfOhc2G4UiHpx3E9wriIT5ir22q9fo06kIuvYM4C2xXOeQo7RykvxRk7XS1iJEkHL
55fBNxKrkyn0OEt4ft8rLjq0HEV04E3UVv49B7xrWuMFREer9xr10ggeosl8F5/tTWM+lg6TwVWe
WJdm9HKg8qOHi5rd7/bb3oQyDqvTIpzg6fzm8GsXcFyVenO2qh6cJ6i5v1485ujw0tX++odKHJxP
413CUV/yYB2z9qLh44u+GvKoZy5ed9s9wmqXWJQvwvU15hMUWIOaQ0WQhGfaWkNlB9Add5j/pD2J
dvvW/Sr7l4QFfi2xITonp/1FoZ8CcT4S/6O3aU0KLoK2k2ptQZRU6w02VP8VxVpRIMuv61e/oyEg
d2GK5AnTOhQIKLJD8U2sPfZSxg8RZ2Tir+ihk00uXzNAu3j+4phbzHr+QRBd+nQL7gCbqvwu4eL/
lOVAO4Eor8enR+F6w23LYujzagEUERciC++f70a4EBz7xKqPL03aT2cl7q+QRVGK9q/uPiwg/0xU
D0Vp8JoVM+hpLfT+vAq0mKn7DVXW5V/dZBdIggMfCHHG/VJpMgADzrAOBSX8oYumO+a79dMVs9Fy
apYfiPg/MAmCoLjXr0TLwIxsXyJNyt4vwg2niNQvbZSSRjdUjDgi1i+ltDAXbrAqPEwZCcH2xMHY
5XSjVZe4H71JuyPpTpgfnSnVLgP2yxOJdkRHcj0USpk0j4InYtBaJ9z861OxZ5UfOkLzhQApbRsJ
q2Ur3OCZxbt3g99yH5+Q0bFaWKKlu8dkdR3aT7ysw+lk4Lne3cEuY8T3mq4cRKOXHwwObrDRkUts
q5r/e8wKgU/ELmR2tVFrPiPjsuUDT4HdaO3KvmuXg62Cj1U2A3zbbczlAgDvRgrYhhFuTeJz8iS1
MW9K40IpJXDLxA0QUfxL1B7VIrot1yrRyaPwqTzzIDS/4WZ+QDFMhmxFfIhFiFPH8mQel35J9Poo
G+I78kLNDCeEz1EuuJCAwbPJ2tp5niSIzhk83aTSq+F9uj7YsfenRvfEeMzzPaNCEst2iSGPPfak
Lvwo0YJPId451ICySlAvt+EdbYqH2Sp/R6I/IrzEPR2/8La7N5L0n69449kk/hJKKexf3MQ3Cjfk
ZdTLk1iHn5J3KaVdsU2IJ5CV0Qnmtp1wZD7KaXb+E8SwXsm0k++W/JpiNzemwLe1q4YRq863UFPl
s2RkhgxEnEX0zSSS5HnQgMGPcelUI2O1oTyoIl2XhMS/F9yd4Aee8J/U/HSs2IpOw9v9ZHDwDNwk
GwfAS/Q8dYxJUlp6rWLRySNb5cuhvnWK7lzboCAJP3fBaKCrYlKoVTuVeMV9avrm//th6fAJ0oYk
zeNBgYpZxH79hg1HrwELXCMxWL6KmfJo11bdvwLW7NO+zb9AC9x/LrBIzmlhnObnod6n9ot4KVqQ
TmDE8XWPE6SVsFBxS858IoMf6hx4zEt7YUemIJEhFC4m0ntQeFq34CeGWQVlQ6DsqEsemkvTjLV7
quWZIMlTCR6wr+GnauMkAIjqt7n0690DQ5yxRGUv5+Wn+ykWex1NQ5bdEPOAPEEtr0MSTp/3asmw
HYrdvmALVKyUaLEqD/DJnxev+sO9rE68PxTchuL1drJEMpY0PKjvE5ODjIuIxBF/sjNf5hPZpGwn
++EBBsTGEMZSFIzhkPh/EkQKmaGhywDl+Yb5Tv7Isjpyxg0fsBd5STUoyqoQPr1sm5OSq03oXrpj
1nvkxb412nfvsYgfeLe0TXfFNwz6RoqOmdabiM7XZd6as28tOk5duVcv/iOsaB6oIc9JrWT4FifG
xQAZ35Ba9WH1NCHsH0BV1Gr5oahq/OmsrIYEBiU3cKWhecbx04Zxr64bGjMTMFMGfsH56M6jA7z7
HJm8Su0NDqs1DkgR3Y4PNRkPmzo6Z1V/qBRm6imQDrOnpOggHwienSg4mu5OrFMHnDWuFd8YujWy
Tamc9I5LwG2TYPdN6BtD+/ZUMfVKdYDn5MLtJbihbGGRiGJBjEw/A0K9cLQjO73Rac++NgG5BWe+
rPXTF4roi8ml2EZpzCjXesJtK1x4Zg08jTtxONcFk8wRztkfa6zjNzeOMcsURweEdMkvJduZR9s3
E4N/sv1e/+wLPoMiBGRSDAxggHjCv7G4ud3FG4un7X3ID9s/AufR20sFl54sK8ux/HS6bw7hAqtt
gbZRxl8/ZGzVCvZjLBOBimek7WZh9ikVcRa4Kn6ncaVIV1CQaQvUTsjeDkqXHdKMpyNV/f7R8yTN
bijYKEHJTBP6YmmnIFYFqJwQyWM2XNmNWp6TvLCPP9cgNVAk0H2K43ezljImd+eYnAXpHgNhZzoy
h5r7LH7d7OatlnraKgekF/S9SMuATzsbxI6zu7tj+ZUhw5rPVMcHyvUMkZod7c/8dYinTWtL1+KB
7KPWap9nwR0QlX5ws12+QgpGmnMQUur0Zm7kNWpXHho5jlqpEwkWTScxc+eF/MElLHyTQ3zlwYbj
OLmirENA/pnOK2a9VMv2yE185F65JngN4IXTZRVaUSujlGzA30o978uAJWqnyevfSRzD3ROUQNiS
h9odZAdCxXZt0i+mUNZB778T81SBc0OALQIrLGJsiiF+waY6fCA3p5LgvjTRW+Eei7jxN07z+k3O
TKhu14aJ5o3c6Cqd/or/u/ccXKrvlG+F0kIufjvOl9UhTgPKAgCwl5IpIr+Tbs/OoPI0zwsVKkiJ
s3IyBsL8UmqxpbPrx0o7mjfeX5iTyD8JC+r5iUPhBQkytIRaoDzAIuFDsGJdBp6RpiVXVKcAmg4Q
KhtKP1hrKHfHFs10JHmQzNauRym9KptSu33i+MRuLP3hw0djybwnespus2wLf2YYWiSPg6B3Kh6t
LswfJQoUhA5YyFlD3vVjjEKoQsi2dvE9tO+09v3jLkHHDKBi4OnSzgtSOzzDDcsu/wbVU427W/Wq
m+Hiyvqn59zRU3zUphF92TnzdkRgdCdifQrxeqNUNEJ5NMwXqnk1IPSvEQs91O3Qok2dqVYskJuM
sbH3tShiR9oCe1r508T6mVPY5laizHSIhQNCYtwH823gV9Mxa29lC6L50Lg71f2WtH153OR9RTse
U2BbPFA4qW0YZKazvKy9JDpLIq1s/gfo0+fnWa1tTacz02tJYDUbJs4KLYRBc+9jGtdY8sD3v+Nk
dndDCPE5PzWI3s5Fvs5bCKzbHSalHfodKk3JZx4bv2gEgBYQkGp6BaT2jbvn93KnbgSZwYPyjlSI
JnONz4Ohsnd0JqDoUCkT5aWH6HGcxyYzLca/PpiRGgNzZigPu9wbe7tumPa4XxVJSzXBzcTLkmNz
+pO2BRbbpscYrci73NFtnmShrvy+AC7n3Ts6gUKIWzahercr02w8yK8+3ls+X9K+Khl4hGGFHW64
FVHu7sfuujKVC0wCQOMGXAU2hh9qilUQF2539e51ETOlyPWhPcex4K7xdq5zJnT+6RRTQWian+42
58st1LZ3RCVB/8O8/OZWYH9EXxXwt9c/C6DI8KuoKV/e+qH1ukeeQb+4RTul9HeuGI08XKDY4m0A
qOJ104+3ZamhjvO7w1wy4ZAXK+a81xxg20q1GZTDVtXVXnozfMeSd35rJ4i+/wi69HmjuoofTFWI
sHN6iRV85kCSYvLuZqgVXGF0pEnemVySTppXiCU2+M0QWc5IRIJ3zaNjDlAbxosg22+3ephxhZ7d
FjXmoP1Y2lOYj4j87sudXTJRCO0kKSfzclbJR+ftP6KNRPWt+WexYamMHjjbn0pHjshQEqE/MfGj
sGT9xs1NPxdlz1SqOilMnm9RHBUksIUG5OCWQKc/akl1d8oBSfsrECBEywnsBTcPuKhXc7LUckpp
UBTpMy7B/LgRjnbX72A8A9I0MySKvjO4tAf0J++51JolsNvco6G8aa2YEZGBkJ1HfKm8Vo5ivPE9
eKf8MhGtFOGDOeGAioNc+SnnoC5Nl9P5/KhSZEBNxzTctxpFuu7dLvv2PRhLC4Wy+nNI37IEBTNh
ZR2czL1pJNHpmUwcDw1jvLqQZDI+9N63QCqsV4FO0+GB8DUSfg0y4D2yGyQ42ZDZH8oeC9wTSBT/
geVJjU0atvhjf3SvbaKmU1YhxzGuWFG/A6Uq8yc6NXVThWYynmselZ979ifckEpitJvenLr/P/ak
XHz9f6IqeByJemmUnnjnRG5RpfEAabDhK8OdHb1OBMHFSIhhKyFCHX672OEZCYE8lkwraV2qR/lG
VoqLbB6mV2+4oF+PsdBrzEY+s4QvJsyyso8avlRpfufEU1PK8EIw+m1RZyv1Hgi1EJWbecvQEijr
UvoP2NpS3uwOk7uqZag72NYwSDMB8rkGME8Ifyu+1hpO2KEAFKO9w3woGuqDJ45wjQYb3HOpmojA
6F3ubCW253Nu4y4CsxIyzGdN3k5r3HCDoQsPpmK+JzjLDKFRfAsF273d6HYbKClSbOI0fZQgRG8p
Vi2noyXnGl1nboWq/xM0dvLgndgYDed1dkZE2TYUW3HFi26TJlJy6gnlROWGOJrD02UERydbqP5m
zjBwBGPHYxANNXN6HkAEtSpFinEY2pNzSdmk4DfgO/v8q6cMv2qBK/MoKJurEko+8IovYNbCkZ/2
XEQgulIL76wig0Y9IwbfSdlM/Mb2q0So3VF2YFv+25rA7h+mMJLurSICjKQpkBMMw3fCvDC+VWiC
R7bh3NNvglNTyei1jsKfRjUwfrhBgEXAp2OVh51P5g2fHvLAEljoG2V0FpEXOTnKyMGTEs3Wmrf0
wiLAWf+YiR+KhrY1e/9rp52GHUq9M1tAMuNpKdq6lEg4BHmzdD1c2Mzpy4y711aUIH5FjwPCcwIR
gLk2eKdc0QRwaIqXzalHN3zopdHBo6BmC4gNv+Fd53+Co+H9X4Y11f46ScUW0K2qvvzIGO1oAYZf
00dhEuLZdf6r6XgHIDhTVf8z+ePRrUzv2oHnW0xwctoAmrGJct47xIXW8VKgHvxjzpEnn0tdMVzt
EP+coYDTSkc3ZyavAFTxJHZC3qHeTMjRhIOnvk/iYAO13MawQ3ZUm5G+9Qvly4eRsHTSqAfsoEQe
5C3vsv/uTmdDs24md4kUeuyv3qwIYy/YVybQ53cBVYvHQ39dY+7qocudOGjRkU2u10Gcv74S9Otz
jVi3HLMpUUvJJFP0+MviwAPQrpgRrrTBz1TivGDqTUNv4PUof/0Gh0qeEBBfTFr7fUtEDiW/Schm
igCp2LQcy5u3TRyJqwFwdaJPdYhVruyBmiW3XOYTZIzC6f9Fd7OVbJTz0es0/B57s7yXc/2BufDC
BuIfLaSFrzEjOiEkBTN+pAlb2IJYKWemfeZ3VJz7ZNW0ylkQ3SCjuwS0qlogKJ0zD+JgR0j+SHkP
2CWEQOieOyn7lXA8iprNwMqyQFMpdj0BfJO04f4Ld/AM/viqqjxsI0+sOxnFezxV09qhQJx2V8a8
jR1BKOHgtDbWcseJ1jBqb+DzOIGR8an6hlJn45DwqsHsD6RwrNZMkIcP4nB3LINxnXOJLXC5D+dN
wB4nh0wXVAKK85k3oIF4KI+TVRjLvQV6azsieWiq5lwSEJzH7WBJoiG7a7c8oays+PHuh8Fl9w/S
QsB3DkPj74K3wEddART3aKEKTYZzgNA7kVsZ2hY2rsjgRT7tuZ3ea810AKbCnn8hL6X1hpvHrwxo
oV6Uicq+kR6ey3sL9ioNOGw06riA0wMBhxuVbmojJgDt+E3iW8ziBfoLrUsBWgLW+8w9yy1acfIR
ePLATniPWYTng8c0av8Uze4oZPmH+AnAYnpEUsPVx9sZ8ZvTiSJxKISZplDjBZmETvwCZ/BNJOEy
mTXeFIgwla5hF1jspwBZ6wyScY5cl4ec8fqhsrIZbSdZS8Jo0QLJs6EGDTcfTf3LV/7mYiSvzqov
ndP/jIwQC4N4qx5Pn2yvslTq2BTPK1PmUD8lUxpI07939qf6HjIa2Ka72qLcaVb3q+CmdQqcEAlF
koJSktWho4/ohNMbccVUldCrWx2p9CYO+4uVfdIg/FH4Lfhl6Cg38mg3rt36reIqzzWoPRN1aTn4
zgt5Bdco6VSLTEuw3bWdFBhhmEgkRCFCK1+HCweWVyk32HnfC0Sfg+M/a8ptfPGDgsV1ZYY3+zar
beOoNNVUXfR4jwl/5fMEB5f+6OI/k1WTDf3dlpJW71mwKevcxpZWV8tXtTi2dTk/TfY6iHzSslFn
svQ0ToIld4SY1NFe+BEw9eyOCgAjq/iDYHDclxOGLUQ/OA+w62terX82wnQ3nwm/T1etN7L+PFeP
k3GUixlE4juwH+V/b5Lw0R72IAXBp5T7EUDMH01HBuzvt4iSxAMILNJBdzsQ60MC0q3Pe0UJnN55
FQmshvOKhxScQzV79lV2lS4OERB11t8/hDRqXBSooZQmdwuHAWMniL1BLUgh9wHWnXi2zc4tsQXa
hzoyuNJg0HlRe8byWm4lU5Zzj5Npt2b0OXWe7p+BSrjVfl6WUCzgLRM2RT6xnoj9
`protect end_protected
