-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
L2hgnC205CVm80LMWKz1dHFxY3C18YYIYtjoGM+Lm/zaWywi/+yxDtWI/vEsb4y0
Y3K88pA2Ipqj/I9Gnau8lBxAJpPD7lYpUQa8KVvF4HBsuTDFYbk2T9sReOsEQGn4
24Fu00GWE92JHE8kCU6KJmklv5SxR9zw82tkfSMGfbw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 20227)

`protect DATA_BLOCK
kIabHJgOj3PfyOcdnKXFQvUf1eQo6MrkabSgAbgZZPHgSqQKxeKGTOrZzdxmYaOw
DKJPxy+yIb8reQ5ZSwVgTot2C39Q25b3vMof5fikxl6bWq6cucxYaP00kYLFNBJb
+hTvrXDcZtFgIVtWW5SjnssC4gBciy1K3C/yaaCJzXjyH/QZc0AKTO72QKxCUSrt
Ab/NH9tPYXqVLgy+jPxLs37TyoHV/HdP98TjstMA4+d63Ou3hQzfMUj7Euv/2G3x
LlxkbmRcLEw+7CYMagcqB1eWXlXm01M5BFKO0rSxQYqiKsORelapDBYwzSKAcOjl
xLc/8oGzRDCIPOMCufyNXGzub34iXHW5FUanFLYPlAp735hRbzWgUWljjJUuwBJ9
+Nk5svQCdRvTHqby8MAdQ0kk1NyIaFS0Jr0Ejt1cclVlIsEfX81BrNVBtJciEf5Q
Kv/Lk1MpINCc5qSg1atwzH0gTs331SQSK57l/H/uMLjR5W1EQjJusmD5XlfMYGOF
JTxgyQcXvGhsVj5UiiDjNZIHj+P4nEs/gq5CX3+JDPQMgHVxxCVMKV9NjZkSPeKP
KGknj+wTeriDqvhli1x6FuuG6NyyFDi/9ipC9CNc2tQgfPTZrWPniHsavY9gRMLf
wjgILKCHZLn3GYg/iUNCGHLFQHhUa0vp0TzyMP1rqQ5yD+tvS90Pc0pHgP3SwJTz
eX5HkVHT4pGhs6EXceLtybSTWWU/5jS6u+26GIwUWUfCe0/QfLO5FniXu1V1/JfX
sG7N5g0dKoxluKmVAlvk9WZdp/doNchEsQ639muZktu2HSFLQ6GBqc5Cn675KsFs
X5t7UfYZPogrVrb4NO67id66jygK2eRAho2kZL3qs6Sil2nkPC4ern0asUSQoSfm
urgSubBgt04z/wMbSaZWps6blM/UKnrl0mSnlpOibHjCT6qvdW22+gSSP4544iZ3
BzUCqVK7y/Y5uNm8PCM/YBUgdbn2rxx/BAk6q/FgUHUBCVqDX1cCzNDz9DobyQL0
XkrhWr+V1lWSCi3iTf/3/unRreGqjazDF682ck2J7KRBRc+7XX7iYqp7vMQWz9Rv
nz6JT6K2WWHtlK/b+7IvNp4Pqm7RLIxOyWvRcDBUypJOIhmpYFXGyiH/a9wQHGSy
iKPN8B7A8DaAsyCRD8TIFRMeiaYH0ACKw7sMY/RnPpDHqE1cmsrP55ipR4n0xoIE
R+iGMwcnTlir346oRvYfLmNzBby2ISz3KAMMJrspbIMMkYYcDr4L9m4/boiAgT49
qLh3xXFxXKnbKSKEs1bnJ6sp8B0nLYncMowgUnqqxUiBjZQoKGmFajHM6kgF8uEX
aXEcqx/QIxFlLHT7MmxRjeFBsA0O42YMZyabJs7iVZ8y0d3GevyAdWenIhMuyBix
2SoHyUhFd62c1y1Cjmub1iCtlCl3az1LOgsPpu0ERy2Wm89pYa91p6RfYQhUd4Y2
NeXu+4XPWCw58K1DG0vD6FH7kYdS+Koyv9SycbzDKJTqdzmwE8/U1P6rUbIzmeZ0
hu6KyhG7NbtOgqvEwqw4+iGAe/kn6W+0NOZmwzI1DTp7T7ZyEqqW8690pfY65eeq
o5IIxjSwfHNvkkK4XYeuVOiJ/dltkeePlGX4o760ceBzGnPa6/+5rKQJs5viomrz
uKZjovBeUz/P/UQH0AE5YQeN+RH97ddEJDpA6mUHkPJJXVECG6v36IgQRxrqZsX4
w6aXIvcweQnggoMsgj9CLpFtWSa12k5KsYXtoYs/bNG960XGZQX9VRhZfRvIUTLV
FCjVAQKMG70l82bksB9ozNZjTItiHoX5fBde7I2OkqIpyjaRD42lZ0vOleZOHnQv
esxzrwXgJr0dfi1b2hsoteafCA6EBCzB/Cb5SdP8MxBz3CbP/xsXWoy0NmBUyoj/
ErRhFjTJntN9F+XulweGo774m0FGtTDaOz1Qb98HgqgE+KfOcUjj25wWyjyseTHQ
iCT0BY4ib6faItGih1nhXVx9tf+3fUzk5KRpnl2jE/XOsPpD45WBtekwD66pvvoI
8IgMe46OmBmTlF4ibQ5YnIXI594pm2oRs3ktrEIP95y3zmPVYjyaQl2YSl6Tf1Z3
W/ldNQdGZlrkYLWl4ZtLDu2vbGDPf5SEQ8hrBAB7CchgMOvGrk6Q1KoxKzzbd7si
lw4y6UXJIUCmX3IQrnoV4p+D5OsMiw+1lrh9PDD6cGVM9SpPn76QXQLkc2pJZl+O
y50553XdYgoRoHL9jD7sjAIZwN/ySDTgTSc2HQDC1qGv0ySJAArVOrzeFSEGYiIM
Umdqe4YCOHU/rV4DtVYqhJNXEFur3XYLRm/a91//DvInhLDaMToz6dGRt5SGZu11
Fqofwh15iwCRo+Zx7vjPVp9nuDs4GxnsqVrclRxPiw5C3qUQmRgtHuRhtUQ8SXdk
g7vk198lSsg6Uu557+nDdDA30tsu04eRvGBQgdei4vtbjOsVyMXJwrsllLr6y9ry
YMbXipVyIj09PvZIEVsc0wwRximGBxbrUzWeCAmAYoR7+Pt0ILOLvWmieDpplBHh
5Io7bsI/cYgRLiETYggMxvLO0YbL5c/Z9hxCiVRN3iW8xPZAmLL/D4HdKZC98HpK
Sl7OW6/e2oDBEXWJ8u/YTBmxS0Ikj/4535BOnck8KRP5de7bU/7UEhLi6F0R7v1C
7l7malxiJY1oUInZs31RE0m2Tuw+d271/FFUs4a0XYwDGmmV6Og+1P/rXdyEMglk
aHyOw3r+fDZW06WVboQ+srwFOxUwdGjDbQC3iPtHC9PmiVpxF22srz8UfglHfdaB
HGdk40LY5zBZU9xnKlYo1xVUKUYjSbqW41FdAmAq/qd0TFBmHdKZdKLnoCYcuD05
JO+RhDLARW/wI9glgar1fH1E6ZQY2Wakz2T+BZ7LJumzhhJZoxAqQFk69tm7aLuG
NOUUvR0/Dn83+Yw91eBJfCg2sn3YhTcWGBQ5XlpwGftVdI4yukz541gs5KjqLAnH
PEq65xWye+9GAZCb5fL9aFfZDZk3E/XoqBx2u/NZ8gO3Mk5exhDjuH8lbvf5DwrY
tFl+bxDp3nbcRcuA/ceoxNOz+Wj6WOYRHL4Y6H5ju02Mjs7ogki1sUYm5wY0Xwpp
tFDVvYspH4yHqsLSQDuBBja76DFsaWU/cN8KJKu1de0b2kgOyO4YBcJJgklTmJd9
PAa6IZ17+f/OhZKgbW1m2u6t0DqqLp+YnGjpHIvwCfDIoo06ywK3X+DqEbFmNvXQ
8pOQ1TXU255GqWmUDP+GlQMGb3TKeWng2NiB4VTYZCcE0rl4BAyiL/MFi8b7LZU+
zDsiZ2MIFr/xF9k21+DBanSZlBhvw1PhrpFsolcJBZVT9RPHuPPGgyjDPPSGKCyZ
LsFJnApr0uJDTj9Mqte5ZKqL8dgwL9pED0aBaKwB1K3tToOOqdVweMjJIUWDXWgA
IHyAC3L1bP+nvCs7QGkECSQY8MeDxnKJH4I6xaFNAHFBkUTOjWG151RD5aLy7w8J
QqA2XuY3NG+QiAOUmZQ9fTtL0MSVpkgXOuJjGSB29bkdQoMcp2gAzUFS3E2V5zv5
36m7lNLxgWSgzNKrXBcsyGSNgLshOX9JTVy8VG68vTV2FLv0IjkwyQmdan06sZvU
OBbO6zma5++qO6qrp48TJN0ZWBuF+xWyT5JlH2b4k2a8z3lG5VolkYo7d2+C1OO+
rv2Nps8dbzu18/SnGYusxYtZ9i+2OzItUQAvMmuzC27rdgK/N/iyqPWa6iLGm8zI
h/k9vHaMHnBWJTJiVwQ1YMXpsOpu1fGN2MclFSSwftyEUw+bwecJwIwvofsU6Frj
iyKFGDM3XM6P56Po83WwHUBUC6ynDzsvvFAoUhC9WvBppH9KqAA4ZS+1HZ+O/shn
gfSzFSEHVlGr+EEgwK3FzFDiejH9tCPncoYmw6/oLHRyUD2tjzmXasM9VJRRJU7Z
OoUWu84o79tjX0f+ebTSxmrHSM6b2W5F+T2+9QCM3zwy1+W8y4f1EA3I26KaaNvx
6JNgDflwvIXGhLa2sAN4vR5VwGTDUVJm74n861RLMIHisTkf5m2TI8ighr5aUozv
g/Oks+Qnp0wJM06VDH5qW4M/hBkA9y7Hd88IEw0F548dRNngSoV2y6dkqxvM1KpW
bjybhfGj0W1oV03OE2Duu8WI2PF0q3KqQedD4BGgPZTcVOvxSy+iL73YxelkNz6d
HpsNpyDU+e0ySsO6w6/QOj83J/+eAr3t02V1E9cYBKH5tHEdv+47x2OVLsuZWptV
Y6SNe2Zs1JJHMRSlIkZwBC5WwcLt3azI/e7EvoE3iSAYrRQ+Ku0bIUd3zEPx/Gmr
CTl8W16MNavbapn2lfuwuOr7rk11OeAhe20Akmvgqv/GMJ7F82MXzYdt0rByGjmk
8X11A48i9wESbXCq98xVCk1ea70q+vZ378tJwFvCTrxxysNGTSHAzJzw3kzmJXKy
y1xUDUVbSbqcEnjrE6QWCMeAyoDnwv8cOM6piKazwr1ZNVv+THXJLBpMAZRvIdWm
vSX2+ja5O69QtPQBlUxImT4HQ6eSjpR8Og8SL1xyw40viMJm8c8jNWvkzEU5hRlD
gt8oqSKUrwPACrj6ge2/MvJ5SVx6I7YwvYRbFKU1yOezooOhVa3EWzQwBfrwJAjg
LTVhXBjcLiA1ggYmAjSv3Nc5qRf7E5X5wyGfDr/Ou19UpEF59EP3dzxfYs4ZdW5r
yGG/05+iN9E1xBsGZQ/vSnp/Kwv3Nbt7QzIxNvH077ohUjsxuUl/3ZvcMDZpR8T1
ZKKb7y5ETvdaZzLwwH5rMLTtqOFWMye1K8fHjO8PImZlT7YG23Y8IJDypEOiG187
xs9vlwSUImKcrRAbeVas4zCChu6wvpAm2ht7o/Tlv7tKPevuTzFS9bTaM7Ny21jm
FUsKiXuyTM29PhnSEg4JNQdllgaUtrbIYpvkXsOF8JLaD6IXJH3GROeGXFYmvpSb
gAt4FwwgqNN9yIDWnZGWNjzRMa3ouiPlD7LNW5wHYau8yQUxWOxbthhU4Y+yydqM
S5sF/ufMuulZWVbUWyN+R/n74dr7bJpBLS+lvceWft2q1pZL1yNtWqGMfFb6vonC
c+FGjLuyI4/Zax/t5gdtf0S7RqGbVpuLiwVcEP5lc066/NvQHC1/ev1LYPQ8EIcO
45N4g8Ot+LuMMe26/RnxqBczdc31tT5NdrXu96d565tHb44LC0lHHTAA6h6LoNpq
AhxmKHuA8kf3VlDBBvzRd0aSEJ1Mr76RVk3TSVcErJS/4tdHdWAgMyrasgBhp13R
tODNd5QWp3u6GpPHD1QLZPOYiEyqqlMd2Ug2Y4fg85OzQH+Aq5Z+78RKYvlE+UMv
LiZavzYIagwp4INagUoUHRTaAY1P4F7WyxAjy9wzWSFlUpb8rZqHkIseBbVOVU5T
QPiQ7wteb311wOlfQDysMEcJt7/DJOo7MQIr6JDAeLdbh2mCjeiO+DUm8wPmgdrV
8J5kA4GcuV6DtO9oGJnM0BJd7jr4SC1p3AXLD6fiBe1DTwh3Xxr2pb2pbW+kAUn+
AzX1NkDj0YKEDpK8DMCh//SzTyiCqPoVlqW6nUQaVJaq28BwYw1jAiy5aJgDj2LB
EQtDWRvc1B4la0tiHmwuUcggKeeYrYmQONRejnIeAv9IthHNVecrUsu/yMlAX7nN
6FhWpPuQiosxpl+hQ9cmfFLq2M8kTVwm3MmBUrXKHTtDwutQKsQXbXsAo3T+FrBZ
fJ/mJt7xNU0HMjSJJVDxw90a4/mGDCk0/Cplop+IEP0CgKyF3U+LismOAeTmnsLY
MBTx6EAY+ySx7OJnkCO6FckK676PffFARjDMp9fv8cvZqVd0kXzG9/aiX5OTRbb2
8xC11kYF/eO0k4IeYFCLi0KCx7hMm1wOUKcqBqMMcPWPoiYJuWA9ZqcQ3ZTjNQ2q
YKcB+CBizgD2N5V/mR/NSvlYXVFxSuxPMv+BA0lH3mJ6/8vXN/y6fTk79hGFwnhV
sALZU+LK/47m9/B7XCuajdnGQ0YOCxEjAYaOHO4OhMerwbXu8fiiykhFYkpro00S
nu1h/d4Cpo0wJH5q+Dj4sk6jTFU1GenooyBdH8GRtJV9vzNFfbJYsSmtyvIeL+VJ
0LdIt60aQdl/Qh6TerOI+9Lmep929FL1sRTGyWIhZsSC+eYqHrp4gbrBY5ayn5Fm
l+u3SdutwWq+oq+T+F3KNDhLGvZqFheBnvGoDdY03AZo1k+RO9nRip26AR2PXITF
Vdse90AslMooSV7we6MRG3k2933Ecr/NS0vOx/FtBUuMuQdMzyIj3ohE8P8oqJXA
UrUa47SwVG4S2MdJK7Ls1Ro9n++jg83T0ddNT9cw2cPAdXX9my04hv46hxNpYZwT
d1lLWcridl6J9usFmSQnYNl2m+g50UevLxN+w7eUtrkywlU8wHNMFCBfSj9Z8q1M
0uKhW/sm/SsZfsqYxUh0PeZwW518/DxDZczIeY4EkAR0ldAUf3MP/76XzS3hRqYb
3wrJrdu+N36KGOk2c1SvJkVGqsAmGjreil7DDlUSjH92krqdr8QTSFZ9aHjbY0mi
3fACVSVL5lXIdTPOxPAtwHGXczKkSLBmenZI9aiQXdn18Jj2Ywvfl6fhP29L2+fy
ban5MRr02ET7vUndiGaBzxuT7bZ2yuoBgt4S92LOF72hJqpQkQBW72EsJEShW+Qg
jWd56TmKlF79ijzaZsUK4Di4Sdfy14hVgTA7VuhiwVLSpKqzBd+gUTJHk41W4TZ+
IJfr8Ywd9h+T8p1WGDe42oiObgiHzT0qDcG1RX5rZXVWR5KWLRaOMCYUHWEKpsnT
xGltqagXjQsOgpLvkHRhdUSG48gUPV+FJA/hj82QaCeK5QSUiwu8ux4ekCCHMFC3
GbxrzTVZJp5yb9ShFkNyHSnvPRhAGsG/d7+g6/P4dMMsguHZOMF21fzLR0b5kjq4
Qo7gKjThAvT+j8IzAqHMaCP/R2N7+fB0UUIFW5P/HuW31pMhI4rxtxWvEmjdOAdk
LZ7kw9aN0GBkwfmbk8hUL39iSqjezIMCn19GeQka4D+krIYxnvKSnoGK2OFQmo/t
9ovT2kj4rSwNNmiBgNgXMCqr/R0/d8jDGJKxMOGzdWiPRiiVZc3O54URt3NYwLTG
cv9yaLcEUj+Ro0EjzOMh5rzOXCzJxsC3fHP4vor19pSFNKE+uC42NNwszXUiQRBS
lHh5NVfguSq6R6TTmVxcsWAsxQzMXM+gImypE0Dni8nALH1PBiTbFdnMsyx2kEcW
Ucd6fA3Fj+hofcqOoTfYGbV7zCy65Z51QGtiLSyTskekyJe0SS/TOgNvbmxGlS20
8Vf0XCBadhDHyNo6K/oXkiUnC/1t3hrhHgJt0fLlOTm7VSjtXxJG67TgIBxm2f27
xXXzbAwMQdfy3ONLpvpg2CWJo6w0HwVJOZAY0P7ExkGHvPt99dWc8qm6jQGaTk6L
cvtE7yhimLtxtr1cJjRqux+QBk8t5jav29vG/6Cdj1fWlsDJ7xsXnfMDyGpAunev
50JaEAC6L9PIoEMngB0jI7RJ3IjjyejYEK1hpe1hgYs3xCZtl/GeOp3G41M5SNPz
I1ASj3CfNdBZrIGwKcPTXvyzuj4XxqECzpKWuskxx1fFVKqQo8wa2nW30jBQMFya
ik1KFtcedoMcpLJY/N+9ofdpZrQZBME/lC8qf/svDEfvtn+6iFH9v2wyVlK+zsCH
HSg5/FCQzq1r7BieLbC9UQm5K1CjzZkfSoPxt92KUxMUEUksbX6J1eiRvCUZ9I/z
X7qfmmzaoi5B9i9g7VRqdGA+3YO9GS9A3wtvxabH6fDLh4izK3ED8ay/ObSvi7Aa
NgHhwyZSlA/q8iu5+nP4N9d/7REkN9iR3Ab/er3vG9+hOzWhWLEQrzyAQnWznwqL
HIPq0ef0fRX1FyCPQeVCdfeIeyLQFVkhqYsUG8NClcoMvSfuicO0tDMCctl+/24c
Mh5PyYwWci6e8FsyoBTDNUg17DgqXBpd922sqNJ78ftDIXKd32crHITpyhSOO2uw
2pYjz+TbdQ9GPiOYIcw+wMvpOlkB7EFAmzm0EKskOS9eS1iSIoCOl5rDeOFmABmx
vrWb8aOzS1g5EmLR1SRWZ+uCG8OZB/ZPWsQJxcJcWNPzTfmfrL/t+7we8HwKPztX
tX2REY+SVZ+BGfteKGCFr9woNCzMgcc3WrsUxs1zOkFW+h0eK+LRG9VAntG8ryKA
5J5Wx8AB8uA0YkoMczuA4k9uDWurMpM9q1Lk83xIByUGDCle7w6WeHhYYoc9xJtV
1qvA0NgxUwAJAH8YEW5j1ZBq6E1tB0pNvbRx0HNQfNqg3FZ4zGyBMArymRmeYjM3
SkKP64SztA1zg2PYWiBlNtlJNDUBFrKdQfHpXtveHesDF+iBm/1IWJIwFKiLpfV6
RcNsJAWynHKPXWWqJXpElSIwChwgV16scpG3AVkizLELimtuKffN1iTE57wsG0ri
sXuTkIJzK6FYFQ7CJCFhoO+aJOoD34MPaHbv+uLCa6TsVwGWkkI4ibeYBzCYUrS7
GQ80yEqvbdW0N+kxTBa+geSiuep2eKIH5okAIAv9UHaTh+Wfdk7y2CmJEaSKkkV0
9kPUJgj1ySOFJrii/i0gvevprzWBNHLxPNfpxJkzFnfef8+7ut+YcYk9yL4k0NXb
jA2OkV9+cMPY/oikd7u8a5qzHKi58gL/FWB5HCXe94SveGx6gmVnE0AqDgmt5uaF
Aqu1kgmxN4U4lYB4eloch9rTlgYi35W85/+2J4QghlLwQVKLh6BdGfGf+JXqikxN
tWhAt/fvTYifMm1+cUpZZRNsWcvlbt7DwHXjwUd41Zrq7hFhKVjUt8dPEuVb3Ybl
g9qQb4gbwiuNsLgTYbHrbLGXutGi927gOZyg1VKKncmpU7X4KVprpTzF2oOWUpfX
8wnHI/54+nxq7EcJrpBG9RZobiiZs7CH1a83qh9zGb7e4k477RfnpG7r1rxN36sM
m4Wq5RAUs7Sig++J1syT71wNkeWL4QBRDN6/tfSZ6geLls9kxBPBNomQe+gFWdjq
cQfe5s8EaIA7XQal3FqnKo/ObmNz3hafjhN+apZysRMoNvLF2WLsBJGt4MCPg+ae
IaeFl0o9fFuBkJHXcluuRpfSTSY1vKlzdbNmXrUhL+BWwNqeZSysI2fb8smtMTKb
26FcfihPzyjI2OWENkkomH38tSY3hig+lTEovnflHSsJdhHgJtZs10Hnc0mEFWnu
W2zv7KBN7VfNhWc3Hh9OyW1L7O8K4gFy4jnyYPYpVYqX8TRogn6JuWFO0NiPdG2D
dIGFJ5a2C3W+y1jy5lQYH8wqFu556nRXe9QzNKvCEkeIHLkO97GamYohgEEMruBd
E1rw+NP5TV7q+gOEFOr+WUDNqH0RDPNWB8XWrBu7arbLHeesQZnsw3VDW5qMLugG
XqgojD3A/Y1Q1ABwejE26Yh0uH1/X9Kns0lJVcVAfohmowrq1HbOA5OTnjFqcpPZ
VAnHNnlZddSSV4yQR/i/qBDaNqJv1pFee5UAgxcNPEyBavh4BnoI6gmb4gxB7Yoq
0miSzjkUplidlqwdiIEU7Ow3Vt48DxHZ3Argk9zDRtc7Ran1Uk8bhlJGRSNeY4m2
ASW/U9l546uj13eMj+6HXq8TRaKmtqf60WhBMylYcK72uTanEQYF4RL3Vsr6/DDN
G1eCsDJBOu9JnO6k5Mt3Abt+041QvE2nXJW8618Eav4rNoYgyVId1u0uCxrAwX8F
POytef+29M9x+bXnX6B3djTaDRPvLMVz2+M6FeobwFfQaUM25V8Y0WCaMkwdf+SA
Kp7crL22dHX5AoBrcxeR2vNXPG38xFaAdT8gL8XvWI4znxXMgMKLWSX3wKqShUCm
C0P0TRSiqOBI1zY7vqd09ZRDhbdGkOdwAJtwNLthsEmw6ZbC6cB9eyLjT989bXsE
Q/Lpx9L+lbrjZsK1u48kZ6grAUTSzWJaxI19pExf0Lc7kWxZZHUT4YtJQdHlml0p
Y587PQ94zJkni7ucgkgmnk8QkYU10gsxTdOJLt544aNJrHdfdX1kLzL4U7qdUD2G
/V7qQqD0QIkYHn5zxOs2mDlu5RSNBGkm4C7Wa39854BfQK8rQzQHCd9PkiEKVsMg
5mhE0gJVk6hxon2kzZXXktf/z1FNzSJyKApxxgbxQEHbLHLsfVw0WX/4pjlyz2ZQ
wD0gVCsIXWI7tATsS3fqbvDW/qyFKGmRuqinKQGC+QSukMvhpW7l4CZ59883IiwN
mOty1Vd8vdiOLL4iC+JahqxVlRcLbOxolSbKoNsGiC3gaejieA6NZMVO5Jbumv+a
O/r3rHl/iCDLZIQ5bJn/m7GMIlzVdGQw5IqBMyYse0pScAS0vTJGrb8CNKIVCm1G
0RlzWG4SrLdbVLg1yYRivT2KgmLfOWTmuHX1z1yazMsTnfeRQN2dYeG5g1tgCNek
SsWKrZtxbctepWYYZF+bgWJLAooQ585OlsjnUZtU1O/3qeDfEMWmX4QYIwccTyU/
CZMnJ+WQPaJgqP0EufVWdXk9Re2t+e1qCa4y86yAmV94Y8+IorMUjCtkKIcCyKLv
zVnrjIrLm26lTFj9/cPhbrYbdXNycV4M0ShbNZXLgMlG0rAKerETIyMhgdfbDi8P
pc5FWz5M/G4DZTU/BfMtnfW8O3hD1cjBETuR6PR1wVjw1UpJf4mcSlA9c8qf7BOJ
EyaG90MU5+1ylciWUjjPNiv7BDBkZQM1QHWmd8iGLfHy82lqkti+/cn0MkY/u6Z4
mq9Klpk3rv0vDSolVy2IY2y+S0FLlwgReTsURFlVTR9mOPog/v0tbuigcSgbF4oG
7jDysI4pzaL9vfjLDyEdqZobvkCwKrc0lm105s9xcffnpUECDPcFsaWPrZwA4+ND
BO4fJPZ6Ie3XRVRLwpH/EflCUBpSqTg4q35pRVfPQpana+nKoZhyrXoLFurqQFoD
6mN2ZqK1zAoUr2HUToj22RJaEDEYwPH1Fg5IVV7SeK0ePhyzzw/0AywsDwZQY1Kh
y/VZmgHyO9iNoeaol8aAkdCmJmag4z6KjmSeyw2mkU76/hBGP863Oc6sA5wK41F7
yLbKuiEf93Dd/e1/yGyHGjKE4e8Igl+OFOrMhPBIgJIrz+Xxo7BIxZDp5+gY8WoC
qJ78Fuo8YQRiupj/WZRQ08ZFv7mS9yTD6j+bKxgSAfUxziJkB2/E0hgelbhZ0e4b
1zrpiU/4Tj+0IoUrH+/tOTVq/QThB6gyVKIltaKv5napMz5V9inpnB8YXed+ildc
pcAdjBbsbuW2gVWuUcTivDFtSegfEHuW13O9EoRVtL5dC7aa7y5OopzwlyBTQuR+
KAT5Q9i0zJR1jOsEXpIBHyrnIEsDi3jN7pB6SiSZH6Qke8ioVAGULXwySI490f72
yVxPSH6uN+hF3ngbW7uWDutWp0fgvolEOA2w3BzWccyhN0KXiWOfvQIxgVixlxIM
dmUuSrx2dIRc77ex3vacxs6tgt9aNYAFNk9+gIzuIWgYpYBBW4EanDGrg/WPT6lN
6hGPgY+5qalm0plX6cVfsZoZok0no0By3IcF334SiobT/DNmOMzSZ3qr/mMl/SVr
OARmaLvi0ZUeWkstB3kgaJtwKKpZcrzZjAPt5M+4WconpUqoyTK6te6xyaCTSAsA
NSG2J7CrqWm7UXSQOkQVbs7UQ4JMXqfwj37/976WxrfA+WEFnf9aHUZylFdA6N1m
1IkAE3uHFhgizraea6GfrFalnwCthFm0TuQpvpVaPsw94vyjilNmy5/gYoDaDMmT
UxQBZVSIFBuJg7H1Ui41dWpEu5x+tx4YyqoB6FL+wWKcZZuk7pwelwRZWcY86O8N
yg5zqtsiDMBhx3ZKomBnYVjJrHn3z61xx87tdDYR8btudoNCgU83ACF24Ge5OUmD
HDiv/B36GZsBYDFE0qabz+r4c6/r8b1pUOfuSJs2QCOKcXkNUdJSkCYZ5As/aVPd
YQ0citx+ZGGKFuMiVVveclmm82VUU2+BIwNjcM6tRkUtc0DIjMVQIncJ29EM6YPw
HWDm9wi3t4fjFqzq1UV4h9JWnuh6AtJ4gpcjqNoHjle7+Mgcig3trz38tXhQ/BTU
4y+39VHN9V/Wb6vuc58uyyLS2ThS0R0znt8Nl68ALLa8JvrN/wN5Ro1w3Icv3yl6
fWAacxMZYM3E9y+zZnoB3+GByI5CnWtMXTZaslftx2AVV5FI3ctXp8njJygo0mKx
IPmXon7WS9edGZKvNrNdFRYg8nntgNNNfWerceCvqlvDchUUpO6yMgNlQP/1DT1/
6Rr/s+C2lr88+RihXbdOKSUOh8YkRqh1Iil0E7nMBz+b/i/P2LThY7FGBC7P7cOK
U60XN9KJ306m6bzYDpcQeqa+Z7b9IH/8DfBT1mCZ83dGM0qoEwtbHFwrB9tX5TO6
/nLS3zxWfLS/vsoATRJY5rOwDxFTgGFcQIFSCDu/XjlrZTUegBs6yzvyBLPbXToL
/QCCvWHZameePe7/QiLxx2lqp/wNubYCkMrh3Mhsh5ZwPcLbCQAwCTYMeo/cc8FW
s1Crkmoz0k9FpAhJZPwAXGgChnwq1mIOzGsPVskbucGT8KBiy3pVY6KGvIs8VNnQ
oFJRRJUtVlF/8FCY/HCziGoj7NWIF+m95PkGS8U5tX5gGWTAJesrfLjMU19K0bGB
QCRIkoA62pDeDZSjTTGaNGJ2bhh++F38RaEEytC0N68V6RVDkDORzUEN2vK9UlqI
Cg/A1VigFWdRAUtz8mCa6GcFQUljI72UhGDSgGvB3f29EwDGPFfesli7OPnaAn5Z
4vBe80sGFtNutnVFJzEnNVmPKy71F+j7/2Bw+rPZqsBX4YyeYLboAWNRo5tqAoPl
rxXVN0K6jr88sR+K0+j3avC8aH878alkzTXTfCNyBFAi7oXxZZgZo3d2bIEP3pr/
XcavNFdj6excoWstipAvQhnxF99v5qRElN7QGLtP0/in2wu5EA76urLki8JntoVX
X+ey7ge3C4sk+qS94AkplarF6lpvRwk8MLxZXioYM+yeErDUUyL/CrXuU5ykCbiM
fGSd1eKmRW9s7KYGl5CsTCGaVWaW7nkCdgtaUSulPy4JtYSNZtC+0BrM8KhKgh4T
SpghLHuC+adTQ7kTDbdRgg7WjOIkDAhsHxuirMOtjMreCZz0s0dHejeVuoA29IlP
l8sAHqp7BEpC3Cj8D6RT3RzQDKHcK4NY9X4Sc80Us5UwQ6FfYsItVhQskTmeg5yU
VG6+sa5bkg2M/K/GmBix5BCCaQI/jig7Ioelo8DPPcxo3mr1nOGy2YfSqxsaP1WD
hd5iCILaO7LkyCBC3LR+ophkpoqDvqsHpmnzErCmnpywL8JPwaPX2NGJjrIiKlSV
GAH/xouYL9SwDwS8ww5o8DnbT+FlTgtqYwsq0Dt4TXHLZaCBkwMr6bEDidkD8Avv
mPBMOeVHTXo7sMZehToKI+gT4GVGkVxX27WuhVfpczAMglyw2cX1WPWnUTqCGs+4
D5T+TX8t2BbT573EI0bgP6Cei5N4g2FdSmBCi0Mg+bNq3jZ2vLf/WIWr3Lgs6UCJ
ei9K6HjVUlsG97XMbJx6Q9xGnHLlpwdRai07cLqPBhF72AfunzivE1hBePAMWihu
TRLkVSR/gEgn2wMyO/QwZqXrKZ+a1PqCOTfElugR6pO9rzIuft8O6ufIXUTB1YVe
xTA17LeMgZdYvpHESt6M0dc0Xq78C5O6etUBgkM0+3uN4GluVW1F+v99btFU2AYY
pZQuZyKg06cmtHG7egG4ULBsKv3NxOh7zW79Vt3sDaFQ7Jcx6/DrrOUJDgZg3x46
+rcgW6RopVF5US0Ia3Z1UQnNmKTS0ZajDyMQCEODU/MLM6IC6w/FHHkmN0xZY/Um
lX9vYjy4+bEg1oRcimzzJnQCv/o99ShHDpVy7vwmj3gnQf0K55mvEobZpQyEMOBZ
yWGfz3TxAFA8AW6AjnRVhwXEJbAGCJsxwUWNV/yympEWSN8j2KhHvkavWpDjae9E
rhVukAMEtpy7ll27m3dAURMc+8Pi/hOWzhj6DG7YnKoX0xYsRsPJOna+VB1Z2paU
bQltnCx+vPMHQIjqh7ZqKBIIlY49d719x00jC4rmWt2T3ffj5UZV/jRlecc6l8ku
/4lde5Joq6ybLuyjIE1erocojGfY+Yl4gPH70wF6CUCZoVoGduU0RAT9b204lKKM
G7QTYIIN/2kJx9EqSS26TEzmDcAb455y673Z9YFtga2BAPTBBN28gzPrSK+sTj3b
GnHJCOF7aE0m75rhCAtzAjsJ+NISwU7gzSEvqzn7hTOa2u/vJJnkRSQe+yhzUfmj
1mYNFXbevmKkkxui1IceZgUcn91NNNjdqBeDmBsXuSJ0V3TqhGqqk8qzKzyR4JRm
KVUJrXzptrQ95Mh6xIqLHOfZ9t7wzAvBdAlZFH/+WPyesl5g7XQEdhC8xmzbYE9T
HR6UOXVOnqOsl/JhI0pnDX91hxBOdpwxaUXu6le9nPk9z8i+RHQofMNmIGA8TAJk
IEOdPe/zYoQ6V+WR0pajr/Hs2bfFhGoQS7F0d1xtn1+ESGKk/fpPah++o26T5HEN
5SXoqUklSoyIIfcHWIgPcfMX8wfOxBQEH9Ghls1ebvaWIg5KjTCpSpoEvlW35BBg
dqyA+Za4nKFw329w51uoh9gDvH+IbJf7dztPTWpKet4cZ/7F7P4VX9lCbsGCNDFt
dsixW5fGzJz6rW5FXa2TjninCw6jdKfxYBsFU43GCUDCwCg2qlmEORr97wb505Z5
UWpfmPJ8nd9xk4+F8rG3M/A8ZKEjfrA6yIM8sHq+1UqmfG98Ln/e3In83AIRWyMJ
/KQ3bjw/czkhJCZxqcFT+5ZRZADeto8tOVpqQFxH3+6QAQFF2Vo6Vx/eaQCgUP+J
Obv9V6WlQP2KmlUk9s8cdqxglPSdQSavVBBXSnTun1qQq8wFcT35ArIRjJkFGaFI
oknvMhWGDaAMHwby9Cf1ttuN4JoWCcLQZZet9H8QdDmSx2cxPO+Nq3aS8FaGCNBP
svX6OHuofiHdyc1+qWHsi5c8Hm7SFIULcVTAMyv2g74arx7QzrPzjXRMyINEIZBX
Ho2tVeRsWrdmfCQCg5fDOLENtuRkSbhdDtVXPawWS7a2ds4gi4hiXz8BOkPCABD5
SBF3omML2Q5d8deF1AziWN5XWXcizoXFLhIhHM+ore//VAajVMXZyNWJgN57S7jd
8nFDjuezTVU9DEIywNt0XQxYQsDB2f0Z4QQA7gB9wHbK6Y2G2kY9EcP0Ys9eljmv
VrEK+PS0lM5yS+w4bykD5VsszaUynex1RAS/bEa/37rlnaD4MhsgaKnNo0/nDfaR
6WTcoHh8LMGpz5SyBIvixnr8NPbJ3H78rWc9AWWmlxK1WeszZE0Y8QMn8ID40QyF
eo0znxzZVHv+tPAJwfuLfErV78SrOcKFKR0jNxCP3BfFgywUnEglDw/BvzWqOczL
HD9O0Ub4cq45D22aWJ8uSVqOlCUItiICn7uAFAYiLFB9T4bqHaOazM3+Be7nNoXp
Y+6khx50GYSn4H3HhKcZncSVbicyhpukbNM45QtHVQACIaNiUKMrP7ZCAXw4JeMF
8Savi0yF/6gYOo9OGTuiAvHTS+HT1LrfAfKCSzwkixU/T5YoIYankBUePjVYijOr
+WWeJ988JsjOfISzKpXHuI3GfkbojAneNjYXXsM8nSER2Dg2Tm0WVKGYLhUY2JzW
gg4Z1o3yaEKQ04RbEyk/BdDajQFqhV2mUnQgCBy7EjDDuXBYDBGIsLS8RDIPuywy
YAH8CTMWJbVn0U/W3x/uiM+zss/Fr5RVv01D1SS+ESPQVIGXT6v8hieqCXkt7A/t
bwHSP5KBxfaoylLuwZSqm81vj6sWxI8DDcyk6TIYg+aMBsDlKp30UuEkAGk8z7sk
af1y+MBIjKMDF1OqDq54b2bsIyifzGfnO6VUM40rPAa7kcsS9layxXkAs82ggz/V
d//h2gog3Ly0/EYXoHD9Zb7ldICFrG4UG5Ea/AjPm+Lt7/a0V7+Lnf+Pmv6mMcgK
dzPmSc8pAydobawIF3b9nOhR1i3iA5XC4QSW62p/9lMxxaDXvbuQ0kluOBunK1e0
hhIALnaekKwdo9P9KR3NG+TnKDM0ZIJJIO0AgS2IEc7qAOAkhJzMl5FTU2AW9i+n
x+vU7WtzBmgnlRjuVZVUTE7EO4HltOsiphUYJGv+mjxC7ALLl1dkYy1Vh+bx2PFp
0rbVJtryIDGBUWTb4KZ4fAjSy1G9CZOi+QY2MThLryVsP2JPCCoZ/g5LyjU2hXJx
k0cpDF1KrzrH1olfyP7hhoMaZWyE4HBGenbmIp9TsDHt/KIfwzmU6dkB1BRsItoG
NDt4tsEQZ7VWkdZheFF0yPVHNNqsLMwvkgan9qh5N/BoahvkotSWvB59uKNAyW89
5KhWnCtaRbARjanC7OHs7k2OYCx2e1DGkqs8y0SNsanZf8FQxzDEu4Y2FvkG1zwF
8+0TMGmXbCS7C4TVS/Ma8i6KxND+o6j9w3INU9JyyGtTR1dfTznoT4bM3PDG6Uuh
3BDFZwdqMYjVCXPeqgnB+sR4KydEyoR/kspHcwM5RFdMLtCEFMXMjfNmg5mo9oQX
viCtJC3Ml+WuwPEVv9vxiQQNRmUXCoLLrivYGj8Vk6MquwUU+D3u0YZyVN2MaKqv
3wvOTp9Wsa2CrHZLTcWbflJy+CxYY5snmXfCc2atjP/mzwZUKxTeuUe4LGRXjb86
6WbFTRyi7uwzM3D+lsFDEOHBuCt7vLs7NFtRdg8dMCujtRaKzUTuhCAOiZZ99x6A
4oZvRjsYNuHTI3RXSF1FX2ytl8T8vlOFkQDv0HzjqMA5EFm6oj1nNZULv9OYtB8h
fB1a7MUcTLCeqvN3ZzAtO+CWSnroEwGOGYM4Jj9PWkd07mL0yunRBeCsh+xTHKFi
mUDc/7U5Yhh0vCzFWvyseLc5C5qGFSGRWu87O8dHd6okZA7a8WlN7brqt9Ipb95U
N3YOTKlg7qmdVhYJODvEUziZW8RQETJJ5J5MazAsXeGWPZoqJ/7BdXjIfqshLj7W
mnvVKcCKw+teleOFMuQ5Ta36dJoyz0I7d/BbN/nEDVajtU+d3dRsbsJoovYOyADG
n72yK82LoKCRj8sL3c2voq0NyEyykqbr5ZisuJNydgITsX48wMzGZoALpzGzbgjW
5qOClLKBsJ7Wcwmb6N+pnj1XeUto4lZmu6zDLRi4tInEz7KnOu1g8KADBEXKjW8Q
eguPYgQOCt6Ui0j/EbOxSJOMZBmS2rEvTUakk+CejbxeiRpAYmiFokfsuBPwdeD4
kDJxAhnbECLDTx1OX4z1qCM1c+ZrgpXTaR5lj8jefonqayQtpojmtERgc3VL+ukf
hr7CJHIe6NeGxAdgJCKzRNCsLb935fciPXTXSNPpYKJY76xeSvMXj697yCOABGmQ
uXYX13e6dWXIapZCMDcg5bK6iOPNwyZT+VEkngxt7fhhp8J5b0JS1kcZr6DJJobg
zD9WIuzy+X3ggPYxI0LhL4ZtzoN2l2qSIneuHZF9e/phd+EH9OtaCDsLBPYHzji+
NgdaF/Hjkyn6n/EE28Om6xuS5iOtnLs1EcnR30GvG0RELKTqzkq8KTmVFjzFJwwe
KjvmFuuuq/0lFsxdgUep+QZ+qVjCicqIzMJdzj/tWNbWMv4vU0unXpT991PP1SRS
ThcjxB73vnUH5xsym8P1ulsuvGs1EenYUzVRjvbwBGmZfnIYixUQS03Vk8jm+yof
SknC123YKgWe126FRp7wBQwksR6RS2tIMGFVC2a8kIjWfQq9DBZ04x428bnB5Lu/
/+TTXiottdpeu1wmwfYX1tcQYwup2wfsV2uElSysvW+CsTWjEvlV7MhPQ9qWgjNO
b0iy8DxIU7vAldLkA1sa4iTAugiG3OV2w6juCSFPizltpNZueBrWYSvhcYYZxT/4
lrTLpEM+ttwPkF7wCtoBprpnyy+/OhuAZl80XN4BZQ+hGsxG8FijM+hIdS6txo/D
1v++zgjyYCszvVWJx67Zwx6Am0AXN75PrYnUNMNgyLDfIKXc6YM4be16slfSxybi
LjnNB6NGI3EUkhJVYGoJWnuEyyWGWFRFrnCktLq/qR1P4HjkxAiTobML0zOksA1n
0mEZ4nOJcPmpInhQWDWLdHLhCfrDwM9ud+DWF0LFC3mJtyLuAwq4J0U7kV5NIfLD
H+aiZ6vK0Ld58/X16eLCRt3ZQNuQKpO/3d7Sub8U/BzL17F2LCplcwWEJ2jVAYz1
YmGwocfTaVZk22A9SwuxbAyuk8NqFmSmK4kVyRW6HaJ+CDXtUEdCgCPaoyX0fDYg
V9hP1R3v7Q6NWelyi9rTG2TkwhvC84pOR2h8RRbXOzuac9AKVIJ9SdUsyxvSOhEP
P/PsjvX1Kzi6XdOWLQze8mcKUAGms7waIwMCwR9lcZxt6+Yov0SpYjNJVkp4Myus
uBbQwDkWDkaA6loWXJVZ7EdfBYz7GlZLt1QS5jhFv5Lj/bKiRKEEZNi5ffSjD4lG
MIsECWpv+JYNnvB5iv1poK8kojhFSl1tWwTKToLWRB+q816Fi53Z+cIDVD9r0PhM
V6yoMd75WxYGFyY4TKcUdCFKQuuarL3ZCQ8qb5uxsBUcO2ab7ciQlrKUAXcH6fNQ
YToqW/683reROH4r2hWTGkZQHmeMIWD3CPNSAydHm/YnRKTuHobfykJZNoImEOkY
XNfgN04NRhNUi31l9Ryy8sh894M3aSoovqh3kNSXsHtkQ4grE5rSQf9dRv8AsqQ4
ewpKhGRbhYGtIvfPa4N6ITMkZevldi10jmEv0oDaEXX58g2ShstOlDaAVEDMtBLl
TKdnjUXvA6x8PPCStgooeO6nKfYd29Ng1AMZ8jyfR+tNyHmTeDDBUONSRYouqbmm
HpG/h+4wOKVTBRlPagFHkOu9zmQUTE21d/mVV5GqXLBioSSUZX6D3ZHx2NntSB+k
A+u2he11yrrJpKreBySwxkXHfpu4I7P1Z/9KQd6PiNasTn3CeABHl6/waxHr4jDM
oQrmciNBSpHLdNA/r5yDfUlTXwEbNMKIb+PwMRcy5nULg40FSGQt9R+XuoS5WHtZ
fVzaSMeKADQlXghVSgY8lCz9CaEyT+qB/9mc+m7emGqq+uJH/ue7feYBKNbf5kAH
Hon8EhR7yQ8uQ1au9khzgIMD9kLwXmzUnam7j/2mwq++mWQrwGPOgs+G7yFSwzOO
/OJ2MMg/oAHXl4RbBZMHBcZTAbFduADPKn5RgoQgLJLcsQ/HX3RcpGF6Ug6FHhwl
57jovB5iGG4/8x2iHCvbq8ZglCAknlQe8b3fHgxYslO9GP1P7doRzfpCj/jgv/I8
d4rnvZ4g/pNcryCZ9LOq5qmS4Bv3Sg7DQLW43Sd6kpZd+7zc22cdBmGHUkyGTJpr
wYMJscuWe8IkgwWteIS96UE0+mzUHAfBJK8L7XdmOJXJguQhxVQ6HL/xZl3OT0wB
pIJd66uGkCK796lAyrlRAH4+7Qzv6kjI6VJKcmBVuTPFoodz48B0qFUnLcvCuQzm
igRTeLP2dzlqHWgcMKYdFvgxJ+IdqlvmYnmQngWZf1BuxODjCN4Cb5FMI3kEe0y7
lHl0XNWWixTux2yGmbv7xH2ZhR+BnSmd2KfXdj91A7kZTz0kAkm4BC6AGid7Q2bq
ZEWOyZZnPKd8+RWQfp/GLDDkopvaMNDFXY43rq1adVhEz8bqUvG5Snh+vJgYpTxD
NUCxiZv+6sc6S/Kmc0ZhgzEHeuF5LuA9ePeGPB9+pVzGG9w+unB89jTz8En3kijd
vbpouTmrSkyDAh97WSxQz6G+aOhCk/H5emqH2Z/Xj1l/YDvypN3sTjN+28VaOzXx
9B6+bB7T06ZcAdCHu3y/TrQDZtTuagOj25Q5IVYDPy3i2TwoqTiu1dENnMOtRRdS
9kjNOk2ebeYXHMjoxXR6CMb8byZyP2dsqSwBDeqViBX5felRLV3P/VyXVE5mGu9K
1CT5/G9r8a4kP+azC2bpY7IYY9j7E/cgws3KkJ2NhKVPRsdRG9wqoRlcrpe5TbrZ
LZEpaMib8/5n9LFiL/70rW9fDARsfeWlSkfLEdrix2QbJnyssYmeBWKy5bjwS3DC
qD6bBXByuY+wyGayVNSvCCUPeYkJGd4NTBVj0uCp75CiSauiUTZNfweagKwTSH7+
fku0rXCzKbzzZ41aBV0ZuKqGhzHluS+L4EcvGx1joIuyhLbhqK8sVjeNgSlLliGM
kjLcMHAIlfG8grhLsK6FpD9j78G/ASemx7sW52jMkVyxhiL/EtuuuIoe8oaEeEVg
+yb7Clxk5xl7cMZ8uklirbd+C9Z3d0BSuR9CzczyKddzPI/f13CKjZQAMcraVWzA
2dlj95K+C0//PHaAzTD6JnpT+9+OnqHpRrkuTHl4RepKYiPzP7ViyaXfXESn/uPH
mFaKhnCg+fxmyE9rTvJt0DYxcE+znxQA0BseGmUx/KC6oBhvNDF32vK4QoryCbvy
jTw2efoL7/U8RhTsJqCaBvyZV9hZx/vPezl2nLNqiueY8DLUfJKtOL6erW+DHVmS
l+BbOeXFuApqCJb3HNr446R3yPvJa4ceJWfzuhUmGXLT43vskKi/0f4x4vUagxFe
p88F3NHKY5Aqm9m99wGNR6dEFPYYZhkXcYwrotMCH8zw+oMS+E9BzdQBnnG1uWD6
iXpoLbhMc23K52Hm8++x2sgltSP4IpQvLZ1Vl5fkYOuL+EIx/acFseLkSVEb2HGO
0D5IGCmwnyV6+YE4k5OQtjapoqa+kT2xBNc5Oowg1HPdpCFVBTs143YaHKOP6dCg
AjuFVIRQl8+KUAKh/IzCvOO8Wc/KJMzHabLOU1TCWRvRsma0nL/HSM/5iBrPajuR
k5h4EgEGLkdVr5Cw0P+k1ix7F3DsiOf9ZSwX8HljpiHpsSrly2p8i0Vu7QnJxn57
KirG2a5gc+TMsjsxJRp7koZf6zVvdUHslPHTo/g22/wmHXbNAx6mo7f8V8/BSP/b
P5ZhTRLLrTOkGMqXw5C1o/JIGh641ogy5Jn4140m2SbAOsfPGsX5N1OPCxXK1Zq5
u5V7wqOEm0e2QzSrfbvv0fW4u3LFn827JQKYNS0zraYuV39ZKUeMp9BWS0XdNHOM
uc7ipMf5SURjhMRhQSUVdoYWhxnqqx0qJRxtj4Ym0FzfkLlf3mtIvbsFqdOBEZQA
UOUdFej0JpN4kSwL/4E6qxggnv15IOepk1S2eCowGsuVDeiu20fatY6tIeoRIGrB
DR6wG+D16uj2nSUrdmrYoO+eMZ0yfXwnx6AjE3b6gsfbLqBYPUrBSNRzYVTOvaT9
DHXj/saLExk/jBFyngrMUNwwhXtZOj6fEKYJLac+e13XXuj55fBixa3LzXC6DLoN
IydTfESwCNT7i9t3WEYGIJuz6cL2+L2Bu4N5wi9uaP4ld5GNnqYTjt3U/9l5zlXJ
tQ7GP5MQ5jtn/SFu9PNftVyZnyclNTdVYWwBr5Qgmft6bcbMLyfNh5Il4zmCQKzS
+Kn7GJdCTKxvOsowtlD9PiIzkdxuPCQ7bQwBzvx/nMC3X6g04h61IefhS/ALlyi2
B7G/GVEPbodPgGjj6HkGsoUpTeCPhjuyc9+g7FiwH6w7gt8Sue+XQmGJZuXhqPXa
ts2FSXTJC08xzV6nvHRrPC9epfqy7q2noYyIp2kGpDQgS1S4myzY+GhtRU8cvz+G
Coj8lgEAk/wPg8HHVjkwbdrL3SnnK874OD7FfiY5HPzwqsCMqq5RJcTaN249zvY2
/ZQ/vNAEKvUxYDYWhuFvk0VpGfjkgIk6T5DJx5hssRdyFM4Rcxh1KJtv4YZiffY2
GmHVQl5sl3IGNcnKtMRu21Oz6MjW4uhIHfuTlEScc7/DyslyYSDsGgPONBzjVMq3
Do17kNqnkATT4W/FoJr96vdyh82yh+VKeGWgIedE/v+wBVo6cov9gBeYCvgH58Fp
k/G/NYE9iZ1YUKFw1oQ+L3HWVeeqb0KCECaNcgFOCtU1qLgXzOX0upyT5+PvX1rT
80xENYnPp7RqRjkmMassQfRzlJRsRhcVTmSgBVbFtKa2qcHUPds/ZX+XSFPacoPU
Pb4sxPq0LUIwIq6tQAObzhHhI90Xvvons/dXz8+9CPJGEKh0hoxX6TZ9A4jvWnL8
eSxwlzmX/bF5AkF84ZNO+lP/i94bwXsxEBedE4143vaJyNrX3iM26wRvTT5tnBDA
JaR9+Ya5L44YvwRXkvnWphHBUaOuKhQqeujq+Ou073aoR9XAHEYs3R58ABVz7nov
GjJt4ia7DjH1fB6mSORyA8ikrdDoFR6LgaN9PmsvxjU3k0UdMntqxmqCYRa1C2wg
+nwnUc7H/T3kuotkewjvcZKDzvqyGkUl0qUdVA1flNLFfvR4OhGGHM+TWL6A1NyR
XlC8NR+zOuDk8412/QGWrjKcNtx0U2Y82cCE1WDhXIWB/R4z9Eu1tqUs4iN8/nUf
O4Hn24LR38BDmnAkmsW6RDpNeoD+CDQABYHG/Bpz04VuP6CUUX7KXY/Tadt+8S4j
gxstHzEDtt9dwKHfD7u9oKzikoGhnRI0hBbDeGNtLraV8PwAY519Vcu94bu9inPN
wmjdu2k53n6GFQZ+ZKN0fTSH9XRn7TYhlhATP7e/l/eN8OL86/ceEKJkN2na/VeK
Ynirosoh521uibcWS4mLZfVvXsC3vPQdLofF/UcYFFomdZuhx0WgmDof20dRsNq6
zy2gU25cweZQJdGWDSGErlENkNVFBestXVcAzkV35R7SCUcr1ccKOnmNByJzzixc
sFrmhZ7C2+Wq1S49JoxRItu9LH7XsH6d/WE5r53DFIKIZvWHt1Bnu6pqZ6veHV1z
elb8OJRVxunNcsk32RkUqJKS2rWE3xzgQwgJ/DtXlDcqq0IBWn1JzNEDBZK+5GMD
OI6mLMKwbOJNGCxbLSvIgarCSiRaFkTaXgOGZLLBPrfh7FgbIpUVaHA1WIWosSFQ
ycSiAJtRetDeHuUpuFwVlBNKBHBWaY55JhltY/UJCY+YDVK6gztq0UdADDWBx4HE
Kbp7W5U2fwKNYa5KuUDt89GQvuPZciVw1DCOPqGOt612mERJfksnBBhVegHUE4sr
P2ZoXjyrGsC7OMHWNhWGqrikXi2NxPl5fl6rWtfzcAGyR8OYWPm82PYqQzO853oi
9prJwtuLxCplNoc+sxyPFUp1yn/f6UZ+l2onc+JGMrOSM3vQ14IhAgi5BYBXLCh+
9eDc3kjoE05j8Cy8VlQRksM6vyfPm2JeZaYFEhQ1/tR4eMZHk2yqJmc8LKT8jNtm
4nX8h6xqiadHXk3rSG0gqj4P1+3PsQR30qEttoe5K/u4tJnQ6UTbozLo3/rjXNtR
m7OgctjZvpc8uP6ALy95RpZmYoMaAlt4RAZrb5y9LILV4WaTUWPmQZIYrl2f5c3e
AV7lpKyMI7GHhjzgF2luL/m92vf/JHOcXYrwP9DRp7spinAC06hO086uEM8TRe+L
CQl4lCbI92V8T69KUeWb0B0eJ579QzcjSPBcyrQPVZ7rNYW86ORluLMzXeNfUzhO
6dWNym2wWE91NXUGHwyudFp/pNFrxA+fNtz7YBa1hgb86ZpTDXJxFOuF2zK3px4v
jGqutHahsLzGjbU3CH0GjnTBSr3zK2jM0jLYAoeO2LBQdTcWDZf6pCi0E279IOM1
mFGrC0fZ8R6i86JOgqYN9WAJSKQXAFFox3Qqf92FHOwlUuRI/8+zHA9FpYz86wNc
9EwM7iuoTQ1U4Pdbdhxle+MTCBZaw4QOMa7VVJhBcLRKuwRk4OERZ1rwuYdzFTYD
lY2k84gE5AvaVs1rXXMbehJd+JY1KcDvDNMyPLAK9LfUVPE8I9aL282WIa4d+Q5Y
0wvcc+vFN08VC0Th4bRXe+j/JjzdV+K2+f4/OWB9UkV6x/zDmu7m3wEjukedlK7i
d76g87Uv8uWggaGPL0A6toT2KwnmL/vcke671Qcm1bFNqU8bO5zIBrTIXXJZA2ji
OJnhlyLv28Bzrdus0Ah6uvlc1+/hIsAlahbTQk902H91SsaycMQWELNJOgf4h2z/
CnBya9wAbiFwI8h2Iqiuql03SKs74VKM8gvmVnmp5DcOtWf/hHYBN1wkn/7Rsa4Y
mCruNmyMljXVpkbHRgJVlcgmNLyuvcU5r0QU5i+nMo3PUdru1kd/JJgdy2BhKPgk
y2LQY9eHuMziyukq70Y6gJGVM1Wu2P5IjIJd1c3hNMRRsSXsylwlkI+b4aqffXUc
RTU4oNPxhnj8f4bujziQidyjzv0mtHbwxkxANdyYvFPRh47aIHn6Q5ed/d3FHNJ0
DGJSoR7S2t344/6moHKTByNQTV7U5oOBSgVYTKaaLE7JULN5MLOE709IcNt1p3KN
MvX7ySv9+XoW0FY/L6O0nzcUhbrhoOSZWAoHzHXkehMisrp2x5qJIDr5f38ns1vw
Dh31aC3O+BUnxuonMiJHP0Rl963k43i57Gytzc7M0qLKFvjJogsctU3IaK6XT6V4
lfBTCNBJJXnvYa4YXRcGV9pLbWAZGwvNvAPZqMgvsfQacFIBKHXwPRErqH/Gq0Ek
aMqFgd926gaKXB0Yteksqojf2LPSoI/WABdX4QmBzDy4lF60M6yXkn35y3oAywzM
tUvXgv98LI5HNqcHjdLoUUCoRJwsK1Ca2pQasC1BTFKDuHTQw66XV7pbwR3YgwwK
zcSm+WNYP8pQgbCLNnSGicj1UulMC+kihSjROJvoX2BW3HM9Tq2UBtUhZcTsN90H
iaRYCMMU6gm/lEcgGBfIo+NJxrT4KApcznDLsPxamBlllE09h2obQ3kNwcK1jW+Q
o3bz7bEyfZipmHyAn7kBZYUujWH4phyrH38Gij0dHfN3ngGm3czbEopf4zMzTXCg
EtrOxslEpxRfAvC8W2u+qexNMymlMWQudWFHuWBDE1STEhLl+6APGwFMPxoy6tLN
G8ObOuEWxBKBeTIGXk3u5fhodumKm4kZCm/gDgh6/oV4mw9NNn9ugzn79jLFc07E
320R6aK/OSltGLYQJdalxeG9w9JzOwZPkMuI1KgWFPeTUqzWhHLrd2cfmOpwC8ia
QaR3ZVo+KyUOSZDx2vEw7+Rstz4Gtlqm1oaCc9ZH4lVSU4JvxxiZyGRqhOThsesc
G+4One5M3/9ml1uAJxQYzc0i90opYBKu1LATsSJmauZP5bysNYjqKB/IiOI7vIjG
jVEaz68lxavpEx38UAY5FivdEtriA7y6z4r4UHN0YgjzcMHyLmPwXo68YO238DzF
2A1T4pIlQL7KjtfeYgfwW672im+rKr5wvciohQsRmkh8N/ADyjS9QLO8pllqb4wD
2xF3FZUEWVBq/fO7Fs311Mv2A9i9Bd+PU6eSq0P8BscoIWX9ndsuR7LpuG6ArRuP
LylFSsCeVsPNBpIwj3ix8kLPhQV1Fsc9aY7AbLkbeCzUsibX6nPn5BaabLOSotXe
F+HUFqAzVrMD2k8m3QPNsxwWEPWWu36e3H5OVJwD8lJAYxF5l+/Eo4PUbxxaBPY6
7J5rpD+XxFnY0Z08v/14XHG/k3xv/kGwEhVrbS66SWLBC2Qx49HHHMdNUNB+VOjc
4JNiiCsNlCQMhyjqqRx08q6oCh/QP89oQBOHiIUop+6kT/D/IUnLCaDL7AXMAbJI
0pWvlAL5gibTaPqJ0qx7wB3P02YO5hjU3LynLNf8WpcRHdw/cAJgwoDdgC1/S/V6
TEB665gUNFbYfvqqZsiKddecy5YGtmCv/rnXmB7bDcRuHROTmzHPvuf5idsc2X/w
l0ApGrxr+qrDiRt/UpUYimRkpwBL1cev6GrRTsHHNPatRElccq2SwlYjAQJz+9GC
3k0PXMLC5gDD0CdIKSDKg2EBb2m4lXIrw26aVF2Qh84V+prFKKj88dzGU7YuD4Nw
cX56UFXfnkG+tz/Vq9E8DWGWMR6WH7QIp1YUZ6OVQ3O//4mo4gsBCh1OoH5lwKTt
VLd3Dpm1py6OOuQ1aw4NP2oJ1/41habyuYup+gMve8am6phsHBycSKpwjFmHJNcw
IqHjzAvcyspoA6a14kLXxJGaRf6k1u1b02ZfQlWWOERN+3jC6CKpX8wXjl5b534d
zdWaLNnXlKoUpRfVChw217fjm6OqJzhGJaS7xlEAEIAjdAmRgBH3glVmCzPcLJSm
oNlPr2HqL+fNaspEkof/tuQfGWJkmyCuQJLGPMEC16/ic9+HzzkmJb33Ax/Br3Zs
WwoIjI5uOeZlSpm47aYwDp94Nl64HI/A4eqRbJ4Z1MVLoDyhhB5p1riW0I2DKKvg
Xsb/W839DZ26Vbeg/kOuJ8w37T7ECQOtQ7HOiEToGzg/1Ua8DoyhAugKYStDNO1k
AP2YzC56HJcO/xWTZVB3+njtZkr1LYvPkcIC/HgZSe6ymlx9MmA529bq0REP6KNb
0GR+7yZbgZC8J1oYO+3ounCTH2JolsAAqOMLv5hSDO+Qa430iiotAwaEisfdcy+B
Sf/nDRfYLtvJR9Yylxcu5y6P7ZYMc8oiujEnq8yE4uQSkY0l6mZit8OQtBIkfVY1
m7eRf149tmT2u6fkBMYE2ZpICOZzsVrUf9AmAEIMoFKcyAcX9JCY2SQqAmdq1cIZ
tam9YH4Fxz5quQIXkO8Zc6HG4f2obkZME4T8/+iHX4vhmcd82YAELdpltqxFSm3U
89ciU5jWq/6j2SHkrNXDTwFp2VZUNozVlXVct8/alnIQqz/6wUnANWVKP4mrJTEp
d2gjKRR2GRkgi4F0wJ5xcHR2BRCtsa8KcnBlluwRB2IVwwzLFxlEoY61uQL5kkKU
xBrHsk0DQZeLBMIgYHCnITUaBkWl5glDsDQBHXZFf1uQ1AHCJzl9eHHDQyy3r9EL
`protect END_PROTECTED