-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Lbrx8ixLjneGy7/WW+1ysfFzTrKC0GvD9hEbb3G1Do/shStSyyXt4+wE2zzZ+4KH1sXUOdS+dV/t
qbvxXnxsVEnksdeHUgT7fnx3Lw26RLERF5gVVrxTbmbBs4mVQW005yifNYCaG+GEvPvQ1QElDIxz
TV2zN43LoLAt9TWLzruEF6aH2K2RZR2Q9BcbN9UsEGZqRaRk7WN0wMdeauCwIamv5mDRhsoaiLVf
ZsTfrSsdbO9edFISH5258MQooL0/8mqlPBStvhjKbhhJCPnJBEtmPkoxrVU/lx7D/WDQy/YUsA4k
5xfxzg20qt8c9Rw/6KjflUQYKovX8oAtoOzIkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8688)
`protect data_block
g31idPzBUfePhqTmPxYrcYx8hz9MwsjH5IMGwnpIoH3fQI0GiyXfcFKxpI5x+jCg1tfZGg98qDIn
AUpuOEmZhYlZ7MHF6/3cHMXjF9ooX4PQmLU2uTDiU+icqybYyyXksGusYamphbLIyAXw0xrj+7oV
OX3Wh8Dv4/dVI2xLee0A58Iq5dnHojNPMyqxxhPCdbfn7NknO5LhAXY+SvYJbxaG7Oyr6cJecmZB
gbHfgWVss2ARZyZF2XcK8+stXKaQ3qMKQ6ZO4U8toTbmmEtQVGOISCrGVI/oSnViy2EqD04+4Juv
TUjM1suqh/OEBjkDc6ZcE4AU6pS0H8BypFpdej1cFlZATIPDyZ2vyMUA07Mqf40m6b/KwCkJ9o2L
54L3E8NSOlpDsJpWC4ZrFVED2+zxHNviZ3BJLgRYyUL2fjfD08w2bBRlljVPkZ0/G7m69IN9zMkq
JkU2twU51FxN4dAmxLVUL0G0VyTpy+8qvBmNiNn2Zivut0Nghi2ec/Pur7nz2H3/1xxHIsXO8Vil
3z2SuAhM83/7rr6yKSOHZBmzYmie8/SRjMpnCR5xo9IeMo2Yr64lPLBKu4R4lMPkFGz1U4MAARin
dvmVVmm2+gFlxBIcgcIgmrfSoAT9BqtSX41+jWCK+JsdsJ2iHYf4IClEBxBLSURYE/paoI8rbJa3
KK/+MX/xGuy0IXPm7i36DYSZcmu9WRSXq1yl58l0ilrxrc4of1gYywADZH2Or/+JFp+MOjnv5pSd
g+pCmTFVCmaw2G2Hkz3CcZviHRffMllaxUOM2WgUBIobZruoG6kUhxEoLsVh6Y6aPy51JFLjzZUV
s3Fg09RY39RMsB1cb+EQGPslKABnGSIxBX2eR66iFiftiGclYSvxYp9k9JfI3w4bm9e3kNSvqVCq
6stBXgeFAoIfsWOqKLdBWoNCn5wl1V+Mxp/CI6y6Cq6zjE35HjuXNH2aj/Yrt5Ac3/PYfswhSXX0
fx7cV4Z6fU25h5YvbcY4uMScLZRYnreGAVVEgTWvtIlOrAUqlIGtcH/h85YLyRmhj6k6xiqPDWUe
8RsFUDjh8njbj7ztpfx07KFO+iv26nQ6QF0w/sZJXMPHsasoXozRr0nlaOPvLRXJIOD+XYvG8jCJ
qylBZH0M5zqMnNCDQcD/rFUBW8QQ7qPbCJueYRj70k+qGGxvkVekDJzN9rQ1z9rT2L1ZQpFFRK4Q
wOEmaCRQIm4XqYhVmy1cwMlS2Se7KlvENqaBc4QP0JPv10H6JTG/SPEHbf9Tae7t4gjGgn3V+IVF
cMcdKRozAw894elLq5w88jpkIWOqsUE3lQOgL18KSRG5mTHn8vlp043EpH8gA66VUsmtAKXpjGK1
KXpcPiczZunvkNfrcJS8kEa1oRcBVosjqAGFXbQQy5CAGYCXnDZowymECVzAxucCpyBo6OVcX1sq
hL6j1bQ6vUZk6qitmLIRaDJkpY6wmShlKIm3Z7/le5pwW++jCNKm5ZFS2IJKpd0F/VDdkqiwCQ9S
UJ1oum2IAKdEYRw37xn81H4H9NXjN/XlcGo/lddU1Vx2OJvYr71Ca40sOWSAmOwbrZe74XujZOS6
DiWwIOobxiQKGM3OBZ5yYBNOzh+Y2/WmKdUm7EupiWvEqyjeCVnv51rmXTeTnRlDc4zaEOIwVV/b
1Lnl5eaMi2VpsXVufDPDt308QgAkaztk40gJc4EfAoFisVocmHDDIetO2zunhGb3U+QUp+1/PXxy
M+d4gCR4fSq0HqQcduQpQQEdflSvdJeEw/mtFtk59tWrXFioyzX7uknJgn+WVf2uMMbFukr2gHb9
Ul3gy+HnievXY10L14IEFKGLcoppQlDafYXY9JVvUijvPGG4wOwb1lAVvwxXjrUlZpO5Dxf+DSEc
Hgh4iyZ5wivNgMYgqXEZcwh54h0ZGq39qaG6ysnY92cP+VYxnNARGHuGCJXr3dORwJ4b7Vn8Dogo
A52LjRNxmZ2y6Fa8JPQCAyfCzom3QZ9ZgdfLidn+7gOzHORb2EQ+yqvEy+h5LFoDeXfJd/Z3aqk+
sxJtsV+C6oMYwQbVyprkutcl8aKeP5XnCbJNpbLt/zvdLJOMlYa99LcsVIHASuVZMhQBqsOQQTNW
JrqROXEJh8o1gQGv8iRFPV9z9Y/JV3UmbaTw3LoP7tFp68ob3YjtFIzZLjdB+29V34weZ5WM0jjQ
8xZ4KvklLhNzwGpqPuc+MEEgFjOSm11L2GxYAq+sHx+MYlwcdAWdiz1PnQZqbrLj6RyjQLVDVf74
9YD32+UX4MztqDcn/8YkqA1mTp8F5RbG43nPRxoHRRDq2VbvDE+QMnzDiLp9D71YB8aI1dGk/8Xw
ynfux9BeNAbNWkvyUYzceAgWjNNIbyMORWJdeIi66An79u/uepjhJReI6lQdg85SZ8PAQqVmK5Yf
z1iidAeKTBvuW/Z+/6MWAUYm2W4Tw3+TJCZMVs9hwcrBmnD0+YZ7Xbozxl7WyaePEkTxCHfhSwSz
EeHgNSHx552E7p/IK4Di/rrG5hmd9Sr6TfQgS+3dtBXGE55VaRvTlN93b7SOOGukLHr5r3bcmrBc
VKtkL6jnn9dJ3pXOoHE5lIh+J+h8nvByZcPh/8wmASGjv0/BOpX9oZc/JXvCzVU93UQYJkMkTsXY
YEBjZ8eem2W43+AkDDlN4UTNmiHBwTu6NtEVyHVmmA9r5x1sksDGkAzc/WaPDcaYYb6t7aqqws1d
LcrghqKbNWUYHGfMruthpiJQIjW4+8erQZje152/mZeAaEqgKC8w3Rt9KdxfdnnD1xLbr8g6Fpaf
glXkJDkY3YETFE45N9T7mfkgWojuIH5bHmk0WKX9MkGvhlpl2xjwOxZvBE91vInzJ8evja9jgmxr
iaCQLwNpKYyjNxbPJMC+BULGyCJMc6XeQr8XRJVzpV9JiWAi4TVkSPtkm7AnxRULIDc0l/nz1mnM
JNnWkmB58qjP2KN37kHkMzIt3l82B/zn+7E46YP0Qt4hiOpC3ShNFbi6qJ5zdJki2KwEPV+ccaxL
7EjeijAsy5vdQ6AK50SeZkMh1TsRg/47KuDNC4ZRVecQiemal0JMKxKX/thpyUtZ+lian28NA2zT
7ME5L34TU0xH3hguc4bzpzDFlIu8cG8MmKPBsqXMJDEjDmW5TyJFmnAErzH73BT70pDhFhYGGPGn
Kq18UNnthw6rcDq6AhqqqN5EZ02CDOYp3+ccBbUlyFUKUxA185q7aHAISBKrDW7itueDImK0z1uH
UYPjAs2xClvHAB8RPrP9MhMtVrfC9e0CvBMfM5YoY81K7ddKFvDXroUDfb6MTwA9WwkVyNlavqtl
cT/S1JswNwgHqkXvPMm3ltCuXixVxlBVD0dBAIz+i7f42jCKh+7PtSpjMM6J8KlRliUlZDQN3NNq
9YxYVRsdSikhhN4psjbeEcfzHv8y9Wlykl3EAddAIMKm58TWQI0LjDWlO+K5fM89AF7pWS6pA0Km
JFQmRvznvHnDLBiufGeKkAQZaOb7RNDvS1eWv7oAoPNpVvRmwPWjGgO2W9k7OwGYpvso3CbMjfL/
gBADvpVwSyiPye5OUzk4pWl6v+fBHwhn0Hhx6LXdFHszuNY2+lh2IlWDuf+J5pW1wulhluaPtqqQ
eJctuTjScBAmyk6duckQ90rdqdUIlRYwJRKZk0v/KgV/AMYq1oBpVhVf3SO6zpWfRMzfWr0x80c/
apqbx2d7AMWYxyAsqXfHWfGoEs6LVt0jgi3bvw4lTYoUb8+09SGBvUSYjoYyjUsIKHmtC5+MKMoP
JjIZBk255H/AqK+gLeXGWGhgEUV75bnF7Zy6qDQqA2rLldixWlds5Msev7tBdJzZR53Eii+XnBF5
e72TWJ2RNb/Hyi5RunqjaIYkzCDr8kBnTohAdM1eqH4aSLxF0NQOJRXR7IeCCW8wfEyP18+ff84P
7wb9vR8H2L1LjrOlSgUU9PBsAmWdwNs4bFFAmUDlol0os39/XYfMXqGtjMam0gTwtw6B70QK6+Iv
3DwmXfeoXlzQzMIx4npzz6XXifZR9COrhSIuQpFxzLDEVL1ccOpH0dsbsfcTVA0eBGAl6H13hsgm
OueDqHOCeDlk08xbo4Tu7Mvalqkx/kceyf6nnLgD6fgQQ+NYX8Jeh1RRxQHYnvO3nEdzk02ffTMJ
JkdDJsbZwywDrqqev+V+98E8h5bPnwztC1fzV2Uzz8NmZkTAYj+AZfWP2lL+6Ce3RgfZJ/9CWpgo
BtvZq5J1VvxPeuHic67uml6+Rbx+BeX7+pNfZaznamwuA4ACFGUTLkub3BeQ6lcRENhj7x40SS5G
WPgDSopHL1EGzm+eXS1sRqhopvf2LVuQeElxyQgr5bMtfpgqCp5MkMXO6LbCu/KstFpl7+sq0Snx
WzGfDNNSRUiDNbpOSL2D8H7MvdU+M8Nmmv4vT5NSqTLrUp+Ekj+cDS91L4O2oIzf9a4wIf4Fd6e6
Ij+/dXPNuvCBbCMn1fRipZRem25c7M8XKoTgfYV9xtmImnyVLzvGexosETSnIR9MdwxGTL4CwMc5
XID6M44XKdYOiWektfYOzCnz+OuncSMVTGc3ceKR81fKhzoWa3ANE/aqDRcgA4sP10e+F75fojhz
weuByQc25Y2W52KnY0TPQ4SllA3UOTs/FLFrAD/q7mjmpyOO0nirXAyqEjI/4JyE3ztdlSeguz76
1flnQCGTIy1xowp8lPbHbXYs5mKMrOITxGarRlDZ/EVeaPZFp9fngUbs4WkUGr406Wb5DNHPTFx2
sNc/qK0JwVcGOcSYEpP8r6scjZKOxxndL4wm7aogu1PUTUmulwmveX414vHxtvTqjGtHlfEkdlPw
1M7+kOauLN3dYVVOHiL+agcZDwc+V/IkV/pBedgMlW7CNIEv6CWsMpqqe/67rVggjcOYA+6mQw/I
YHLmcVMlD5cZns9ATNYxVSvRWstUv/x/VnA2xmhQwFb+vvVJ9bzRa89jpiSTKf12PZoz+zdqDTV2
T5F0SMGDkTowX8sKHb17srOUaIggm3w0f7I/gYmPGJjOPjGD1RvzYeymnshWLu9XWetpNtGTcBPN
HK9bbhhTyo+dVrbjefrOD1/fq2u8fcUpzifHg8G9++lw+UUm5cXLtGYJdvbiM/jfzv6xn2D+eafM
xTqnq0rzjtpbDNOaSlt0ywuXzSw/UeXkPKsTho+pM8ReeFaOg5PX7RvFjhmH5JVVVy1b8KmDlH11
tMh5s4osInSUEFMUBuSTGXwRwUqy6/4nF9BlVs4gDvWvbHMk0V7/Qbf0iy2P3sWbgkSZjL3a+y6f
5KPTKZcylYB9kI/02aRfxH6rUjU8cmZky7Sx/NFekaoWAYX4hBVcefDxjArLcmau/lYPpljZKDeA
oA02VY3v1MNcBPq3gU6MRsZBrPflol6eZycYSlLDjO0ykyphsa9QvEW5kDzs9AheeZSldFS6MkOg
bDhisHNzAq76U05NkpCXziPXpfig6HKUvcK1jwt7VLVhPVrwmb4Y8sDvGhXE4C9NqArSUmgUtY/S
qw+kVPyJRRcIEtTIFVV1cVh4rLCSWiRUlvjQoYZ3KhPhlhhJlqrmnxcw8NO4+iDhBQ/6mCi+Do+4
9AnlV89wHxS4bJKLrzYH/3uzMog5bD5bBz4nwM7JTKO2kipSf1V6mpd5to4pCIJzdG/WSvq8j9LV
JVTlWN055UQ95pgKUnH5MFkMbkLNdyUtI8lj9KLnfz1FlWDjbmrrshwiLypFdzrFyH0AvdKUCKrJ
CCT+OjxRImp86knpIaeSqLO/bhVLH+dz0j0gAjUlrChuijcGKRKC8NQoX3eu/rgifGDJPGB1qmka
70AU4tJ8XFIBVIRoZedPyE/xW8R8YQ4aJOR+XZLCRGWpoPOhakNAUM/Vl6XeaaWolw4PK8Hskzkf
5GHlevkt2ZNNwIZQJp6DsRMI/5YacIfbfxDTAlFmYdjnl78uBbrD6/L4AjN+/jzZD5Gji9NrQUEX
Ebssw0dERD1dhIjH7JzF61HkX3uhhINiLAIiTwDCDBta0snbrxCBmvUblhQKUe2zimj1lggxEeIf
ZAnAPLDCGj4Ti34DZBjG8mi31SlWzjC4M3urTOAfL0oPY5HTq28dhZe/mYTIfbG0DWNRf1bJJpno
NJsKxNoMeNEpxtOYOlPjO6lKfo8F+B7uCWYMScmUwrdvEDbVqGKoMbUZMas8VYIyvuDGnS5zcRrz
a1XaVSdrnz+Ou+8wBsVlTmCKOEYcjXVvt+gBYusOACH5gDKU9tg6xDdHd10Od2CQ54Je/hvTwJ4x
+c9PBRALgSGCgmDucPgVTBDBV5/RbWsF40Y4QVXPSzQmGX2k1Ux1HyHrp9/gzsJIVW+Gegva5n1t
6TTpGDeDAiDiAXHPCDLQRdmmG413zD9P7Lq5XTTxjjid7xeO8pT6QHI2TBZSKb33UiAtQegaWb47
45AHluWOoXkJgY/3ZwPiSiqcogiqj53tFI8SzRjKi/+3pUCcbds4yzL+AOfFCrsmQKk4hBR7QgSd
WHSrcMYutNVAShm6RA1udMulDtMaCp++DpunQB9JQ7t3sqp7h5GZ581Lydh3T3VAOpkLtWdmax5E
X2Pf4iUW3/Oyca6cOCgIeUNW1oDhkwAaH07te3fp1IU811R3kpY2dts072hG70VUkcPBfGmEKuYH
56ntn67+naUkrZaqvZR6Az+9ybuU17c6tmYt2Pbd1wO3ciNNA6gLSJbp76oYHzzwect8FzjpKKE9
klzJ2r49a4KhQwN+kXUoXsO8+lr7jx/UDnb8Foys8TFHmJwNJai1lA9dT86p9ztlyAQlChlT8y8+
2PPDA7YGETDzk9lEVeYiZiBLW8obYpmvDbGpLFqljp6ZPy4w3YkUR90wgf+gNiUTwVs00vDWXRY1
GQZWBSoGuqHZWOS46X4yw9STR1ccGAmAXH3yZKs6W1lNqAnsoJtvAr2FCpo7OCbzBkAt1o9SE1vM
uTiid3qIBNYDrfnVX7Cy6i7krxQBmWflet5n+a8imhsOn48ei8hGfnHIFGT7k0huif58/qdKaaDU
8W83ZYEqoql/gbq9qOcwAevoHwRbe7LXt6ZaYzpD3BqH5VOplPcvhqTe0MXVXZcs1ENX5zc7oaI8
qObEGALj2uc/vu/19A6iYhEJrnmKmkKAO9mc2QeHXlbQdDxjuVFYzZ8WBXmpRpK8YRCG/H8fQ7Xu
kTxxd1XU3visD79VXyc2+YRM6z6hQk7WWmaN4aDWQqkKWrWVG0r5Y4wWmHkO+wjQCAfhq5kclurW
pP/O0VYaKuLWcyIg4WAj9r77Ytm4wRNFBJxYwkKxwR5aGLoceYN6xo/dpdQ3VWJTDwf1M6QvYhR+
3OlOKhRrtcs5ZKocl435jJjUGef6q+EvbH1RJpBVIemNiXUEbGICvw0ppQ4Vq13lFqKC8wUCz1cm
D43trxMSJKn9lKgzCZGfvGSYg33g1sLjvVde119xD14XweBroHj0P9o6GdTBUGVsCB8+2UT7WdUL
9idP/vhdXSVOwPYhsttuSWnDCrLVEjJzvhP/PKf8Sq0/2g8cMRIC/ue/z/oJJ6N5w7zeURypgbFU
YAo33dxCcgmQ710azNASYvI5j04uLSFE92mTp5IgW8Y52NZNgd49NtNEeccnYQpGHOTo6ddW39LM
YLwuSISJZYnAFC2rb2q06SwK2u2sBIP55FjRMbUxkNZu9whwdY1Ya2dChJv1nIpwBHibq8TohbbZ
txo/wwbkZBl8xraLPljG6yQgcQKrj1uWalGoPTc/seVqJB9MYrX4cOVzMOMemlWuqyaiYgcTWuw+
WREP75/09sPH7O63MvATwKCVUuJP6a7HvgK6nCuRkmnAt0ESG2Y2Zz0TD0XCtJ7e3cu0kgpSDsJ1
4hzpjPqEMAPJhenWSEAkkVm//SY1aAhgoHKehArRys25taRsKED9ygzhHxkpwNqeHXvTKqbm9dVz
Ce1vRFlrEk0Doivbpl+cmCHjqXAtOak8wU1tM2C7+FB6P1ZlKy0FDKzwbB7Ol/fLEgH48SA7KhCe
/RLsPUGAna9WlZCnu9XSVNDctN5PoRL4frwxp+SU9MTvbO6lwq9uoSPYYqG9ek742SXJbd54L16o
jjTlrJsStoAYEC20pucfEf/HyGraZZ9ydM7rWMnP8VxnljfsyYDuV1uqxEbdf6hNFs2rvwF24rNT
aNM1XJEWlBe7CR/+BFdExk30hDiZP0cos3UHOq5+svIIr0r3i1LJefrYF79M4IVv31eyndBJ3oN4
TAYzTPSTsymM9ghRw/hVmZ/sNrLSiDwKq0b4EVBfgemL9LyDcMyPggJqUugJmc7kYysf4JZMFUWW
axK+j0+SC6unfhx6T20++e2P5P8HL0mVJkn5rLDtfUeRswXAnDmyv2EYM27dklPPTRZuegH9jpU5
lhK1hWpVgYKinoPTHVNE1O1zUGM+Yk3AiqoXG8+f+1to1tsspylKkS+t7+xof2ovR0FhN8LoNupl
+xCBmyHch+XE+uQEG+EA0mKmFw66hPky3qaCU+YQYU/v6rC4YG4MXg83NNIiDAeTlzCaopLXkuO4
BXXiNnn3nSj2ZbArX1QVYOt/TX7hu+XTIMnqJin2pDMf20nOHJQTveXNNkO3ClkqWxg19UpF+Bf+
xwJzMIAvFZPXur3HIvLbhKT0PYxt9yx8jFbb9ikxI9ZgbpopuIrOu422stNPFHRDsbVB03LE24j2
TbEqsmGjMeRqKGGWtVRmMuDNj8xZDpwcWieYFV9DiNm83HfJcZpCLPN12OT21VNHft879eKovHHn
5m3WHh6AorCRTWJcH5+HiJj8PudewTbQzPMYvUhZRDa5O7gIbaCBf6sD4Qadte1TIZgna+qeMpa7
s3pZB0UdlXaTxPtlla+sOlYC86bQzyh3jxY6yMqwURiy1IEQGBgHwdqkzRTApjz16SbMgaN7rCwB
ySSvlNguu0He0/PTxriEGV3Q4m0aVfpeBKXvPo9Q6YzUJTsFhEA92bCXNKht5JN0ZoyvOL7XFjt8
9ESwGaqx/+9h5P3shUyFudcBq01xxZ9UwJQGSUzkXxwVJ01PONDgzkBy+/EU6JxZM/K/aQVlbAQt
OfJJPlkQ9bUB8uuewH1NvoFCF+W0LQFufJ7y0bmutAjRLEZizmQG+nrxUKGli2YmU7A9n4yY83Mt
kEIDqq4ZjmK3c3x4gCHcSg5M7wg+6MRMyfQuVOWE343ygcsvJZAD+HS/F3c/+c5ccWaNpFr1fWKx
kL9Cj+epUpweq4dO5gp6QbRQ6nqcjvIqa24D/muTZE1PC7S7nCIft+a+TV/Wy7kHLurkm696xMBu
w4FVBozf8Ov+9XdUkjJOEU0RigxNrhPDCQ8yTZAP5EyBAPoRLCezrNyvUeAf93ObTQZWrRIKPJCH
3ArViyg/RIEusQdSSzPRf5/Es3Wl43xtEDQgjrhfJ126gZLe7hBPUYyiHjl7QWVvERuQqrhu62e2
RrSI2zNSdsHnNLHXNGhX6KBodOu8T4f7M4FfmmF8z54lmzKdcyDuu8GsPSieT1eAO1nt0ayweuJx
cs+4yPNZaQJlOPulgH5j2wdjoHqwUu9Alv1aNdVYyqOQLFhd+OzMDo7SceNecbfm0P8VJR2Z3uSm
HmLN2uNnOe0PeVAGO5wwi1DMVtOi19xvpAz4uqAE24G8NKprIdhh0bJUgCOV/15P13fWQLfs2Qt8
IM2LN+muDq3MBp9tEVH8nZ3lzhkMnWaQWOJHf5+RxEilvJXukSWgXAn45/nI6GRnBvQIfSHdS0j/
XMxcB92STeBK0IKx3T62pMnUCnKpoBQRhtjRfeFmk4n4b2iLzOAzu7/mlhf0r8AlZ/kdNPCqHtfi
TSh55zgCHw5H0zHIQzrBRq7ipGCpYintqISKa6t9QfpfQsN9R1a6Ue3cYaznjwqegbDOzAYpObDw
K0qlW52a3HfgM2jaQkOAfHH9MAwLLzyv3dQ7XK6gj8kHFsLNfzYXYFTG1PnDBWeJNjmpX0hBOUM/
bydKvcvwIiLFBhT4teSSTxFaYj6dgrS3RdZANxSCcamCj3EfC6NKgcekdw+kX9I8CcsAwWjutd+b
cUg+l1muX/MkDNg3jnnE4FdVn4w3+ByfxSvPXGY6TUnUkHxwMvR4rTrr+MJIfP9eXTnF9U/E9tmc
T7HRs2Lb0DmQuBB7Pzah302BKHZLM6BQbehWoC9ZUpzLMyVqyi1ITa6rzVGTlNDBCKQC8dTTg519
kamhU8q9hiU2X9cAlrSmPUuSKPLr9LWk7GatAoleOtRReuyb9nSAnL5gqFhu0Aijo+8CptUIQQAv
UIDhBFsKw0XbSsBDWlfvhKBCDxwo7XGQYXT8EXrJrwvYt/Lqa0JD1yNx0V9fn9ETGj6Cm39SjLW7
X0fV86w8IRTyWdeIeAFIk1gJCbaDZ8bToHZ1QHc/nnSGuj1SKJltdZiPrRzI4qJ/X/X9ErGrCT+q
dSLr8WhykH7h7WJSimDX+HRb23wQJSq0nh77mRpOtIhRNYeUbqWMoC8AvVjY5/nyK2ulhj5fxgaa
JOzxxZu/OV2U5tbk/i6yYTU8iK47jPuhkmCr8q7FbHH+2vzPKSaQ3rLUGrpfCaQPQK3l/uKjhmP1
1IkjczgI/cCZ+GR1oJFwtrw68LZo3jl2r6JMYv9FtBWiAB+u1ntOyv4FphayXLlCXvYKucPF9K4X
Qs3qKAHETOLDXyKCOu/OrJOp2icdnNYwxywXw9iuBgIoqLBlhnfbUr267wxs72Tzem0jBQMgA0Mx
j2vnvQkAR421IYW3y8kk6HF9AKnBFK4Y0P0EelPCKUVsN0tlNFAXRsfykIy0HNdHRd6jjR66zWE8
aaMgxeMMC11u82Z0Q0Xb94eiZwcMT1A5k2PBAt2ykj/M+wXIR+1OY7oxT6vY7EEFnPFW7v8j3/Je
3jl4+qEyMIk2yIp6LUbSBgEYSgT9TEWG48rTf0NiEwRKYdrGxghwyfovGx9lTwAwuR9Drm18X71s
MMhnqCZo4YdgjdIko1YclX0g1E757dwVjQ7+cAavX2OsaXGTngJlQI4ooupLO4fnpkOMGRYagMTk
27nmzYyc1imc3Zy/B7+X30Kb14JN6leBGSXMlEbk8bfCy9UxQLDcuLESjIucNCDMTUq7fJJ0lGg5
JCMwC3i616ALLPCM48vojMgPsLvHd9PZHgTNV+BY/Q8KvYisagvCANn58+bYQvgZKs1Ru9qnHF6V
vZ2Nca9zu3v8+ew6z3QsyW3FSEQqqCnoT9r0k+2gqDkzwwB1At1SJmcFGtgFvzkzssEsHuVW3ybO
DMqYTRKj2aBHfWpbv3UFuOFxOTv0qKKJQVz+dvdri+9UOUcVipX2Ghy2LiztZSTUpu6JvUTaSU8J
p1o2ujhOOjuv7Mijh+TWH6NwtQu1iHf6Sa9xU8oUpw8P+Sq5it1lb6j1Qyqcl/PojkptnxQmZgrJ
45b8Z7EsJMyUrYwszs4fzKpNsHWtJCFarpvdPPE1Fbf5oMpV/fqtiGQ5iw0tJPc9F/BgpIJWog8V
B2mZ0GN8n7VLPWt4UGn16/PGYVp2GFDK
`protect end_protected
