-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e0VhUnuSLetxb6/KRGBGlIuRubljaoqxKkSuMUsXiqtqyLDLqmemukZmaQZQpXCPqUkiHdlfZaaW
5SOz5+gekPW7VAtrrf3iOE3n3LQ6FN/vP1lVeRmuFs/I7IG7yUdu+9VKcHzNAJRteNx6SIaArJGR
mSS2Zi0BPwWXT0dLMX9shWvPX5W+VA2dUHuguAL7r1G9l9kCu1AfIiSwifUFiKkVcVQSCbf+WpXY
c08xI8Ywpzk+sHJoPOri2hoIgstZ3QJYK7l87yalySkHUMTajsmimyFsuT8h2XlvSZKZODuC4V10
Ov6p96b5aNgKQX9m8lpoOPNAChb5fOv1fsvXPw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 54688)
`protect data_block
PBkCIcrdXUWm2+lQbwz3PUHhGQjAw9rEB63C5htK6wV2i7JgMTyyD82gAVRrU4GluhTPPeFS4uJ7
x0j+12Z3gWHnHcqSFxnI90AAHW1Bs04lViE84c4tOcS2Y48FB3jITAlsY38hM2TqS/vNoz6g6zC/
J2Xaf+SbhpQ7YON0dZ1h7rEVr8sdrtIuqYaskGmvYBMFmuFzMdlm63eruMs5tv2/BANVJ//7Q3lm
Spp3DtXeB/WUoX0OJPrO+MEsWllX6gDYTnz/bfUovKqNR/R541FT4TW34KTbItY1QkCnJmD9dEo6
ss3g/AZ6ecOmG2ej4vYQ3PJdOmfl1qfPRExEXXDJTqYIE51V3k9EWrHFShMsjuAcDghew00eWJtf
r990yMrkMJDLE0cCaWzVXdwWVMWTg8Sz2UyZWG0JrqA/1p7RAzgic3o9BKzFvaf8cDHYHEsVLV44
IXpxBVyaiSlfZ+JVYAiBm7FhtiKKRLfG5gAAtKIV/7RGCnI4WaSIWRAA92Lr/SlBJsyrvlZd74Xt
9D0nuTw1IFVodEGNJt7cYCtdr9kRktl2sy3ZQbtZzHFOPtwBOcHlBMVHUtc2O++vjkKPT0ye9FHn
2CJcglFtaDm0qGqT7axxwAZxDxWYzzktVxeclX9Ee0Qql+prFAGXR8lh6/7jpLrtysYVjkNqNEVL
u04NNxvy8pVRxbIw6ATUqHzHvjU53ZDSpxukPr4sZyPdtvYx+PSmGL040ciGiV5M4NIBmDX0IGsZ
J04733p6IjkLx7BcV2h62Hk3dLE1fGZ/J8QiHxcdei5JjiW7W+pfq6auw19L5ZOh4j/cX8+sbtJv
fLgCFYZVM3aSLSZ+Xy5s6mv2kKhI9iOi8Aap27dUi/YfoiyMflNXlNHZ2QKu9esSY3h/bwNJ0Rq7
oEugDGHPLmlJurUcRZVCXCpXZABi8pRZoCveuowvTWv9/clQBgUvKw8ty6hFAiwCzx7z42MqXxGW
Oj07yTwEAkAyYB/35nDcY41bjw+s6+/Sz2cGkP0fSgrIb088dUATVqUMcbLHrhUNi7nLpVJH/7EB
CNT8CPIH4aN81f9QgS0apgS8/fsbwEkdKpTCw6CBFXaeqmLSofxFaQF7+udqByX/RbBmq6q7jtx4
a8JFrSpM1s/KNa2egtCU5tuPu/bi4jZctBZvO04eRXbmVts41GlCdwsPrrkncZJl8ZvMl916Z14O
wi59R8dttJjIvyG4Sf09j2JZzAT3nwZUe0zXcGLy1eqnzOvbiqTbIPZxdK3DaFcCBvvLK6kLWqr9
MojOahcBnqz5rk3c2DVkCKY7TvzodngdtugS4nfffzL3eCGAGqFb12yoJqdgA05HQtzdDrXz5Dve
cRTIus1MoZzphlmgxHOQA/YCSPi0F2MWN+NAAmyKjb46OGyh+as1CTuEEzo6LFGNHfNPk2xz4Sj2
cQTGm2wpCbzkuoWDJJOrYtFDxf9HFW+549ZOh/sDNkLdAFyl3KMEll5tP755eLnFxM8/yBUOvh2S
kz6keOruO+nd1Wa/HP7QoaO9blFXLH/4n4Q2MOuCrSMlgvxXvUVKPITKzeW16jiU+JuYLkJTS9au
J4hRksKFcrJ9r5CyVAjQjlzEAxlQw+HDTT8eLnQjSgzefNWJe1RMTewrHYc3x9c+JiRaZM1phMK5
2iyy7+YG5oAya/nrDT1lNiRIQKDutW3dd4HBdvNIgNpkctZEaojwf652R087T8QTrP2dFguF8Yi9
GOiDdtwB58uLX1woGuJEXVAhAHTlJF8rncN1EojJMeUPf81/zGb+mDOyF5B+4ivDKhJBh2bkzciv
gEAGUItVAoAb7R5ETZSeASkvc486iBIHXGhDPb7uP7jtDCCeRyBajiQHYySXyrE1Buk/n41a8uwg
Qapz4E6pS5lhSLTcChlh8Vdp8X726I3+xn7L7pSG5/0EF7u3v8mVa0fwlEeqtamY5LdLKWD+XWhr
VRZyowSYBone/uvKzTRfZ7W3lfcGGyJhrT0Z6nUc2xO6OIG30zOa4Cx8ia3J0b+OuYXnJI4WFC/m
FTbgqFPzSRW/ZATeVDfBlb3JgAVrTpoQeojQkZfg0Eo2keVQLBh40Yy7V0LdT0eI2gk3VZXOaQ6U
0C5voddtUwe2IthBx/Sdu19s/mdw/sWImjktRSWssYxgH7K+FPLVZZWo5EXA8ap8DO4bx/Whhj/h
/x7rGVs6XO4nqlR+G1m+2M1Em7sSusfPdwc5xtNRDafg3YKfXzLprKmGz8Qn9TPpruuXH47K6Im1
bLDxpgI5am1GmBTkpaihw2xVJSaUqGCNO0xEO98zeIX2EY7csZRo9Xb32f+N5iu1/p585STbq5zn
V9U+2EJLBQJQ5Q3YQ90KbWistcqIQtcJv0YS2PhXN2uU986QXzM5akLpcJUdpBD9EUWczQWuCFNA
jqKgDMSQzU2f6V8LOcFCOsItQdT8as+qiXAXcY9hiSmTEGYmz4oWB3jr/TeAgDerGN6c3+lSNgdp
+sZ9QvibT3IUfk/JDyJj4LLg4K21C9PGf1bJrR1Kdp3c8i0pqngRqrAQJZ/YlNa8K94l3liK5gl1
He/oyFXchYkD8vxhgjZi7u1jhjxQAvmunjrIN9fIDpMBpmpb/NGamnak/pA751AKO4aqSuigFT+d
k6BuANNyJMjymhHRAFgNhvmrWJH0pl0oSNrT1ZpScddXlCQccnLBmjpUhR/b4JGMQvq7X9JO8PiS
vJz3d1Ncz7d2Z7janGxbhE6r2w0a8bryr+cGW6Ju6cPUsiIdMUukbZbRa6raqNPc+GY007obvz7l
QmnnHNkFT2J8QfrJG+x7+AaXg+TGDS4q4svZpnbJa1hlOSTsQ6YdNMFOpUvLA/9KdhQR+qGVVhXy
D9IUn4QWAjkd0iziqivOTpq1LD7eLr0OicL6CQMYw5j7+GUIwVhzE5r3D8aKhKZGdniIfkBMevsJ
DgrZvW8KR3syAhjnjLOWh/85LtJ04jIGMWdQHqaSe8+t6mfBMG9+X+A84uMMWKuKefnnvJ/XTnFT
Hn0ug9TOwbuvPE0lpu50OsCnWo83jZ4ve/R3X5sZKvn1k3GTQD00EAc/lHZevgERn/XNXq1VO0b6
vPP9oGkaGSUxN7NUyyJ/BpdMFi891EPm3XUk3WZzPU8rI5WzFCsP71Pfo1QKKwobPIJt+2M9JQ/O
hSgksfeY9s6j9SsbUSbqKjlYXUtzhGigzN3VmIhKR56AnAkbgOv6eghztQ4Ez/Za2A+xKR30LuTJ
isBPv2MCYJOPm41LA8AquKquuJ1f8uHQLqdM7qv+2IBzPQoUUpvAcugVGjQ4p0I1pAuudVgYjfnU
4iYn3t5ebjp9FNa1NYHnYwc2dqc6sYBv6m9DncKtLfwCj0dd86k/5H3qEnTNUrW/wZFCt5kAWOit
iIW6Hw3oX/M2HHCxp0AtrE194Rswadc3mHw6BNe1nxbui572G6Pe+3f1k157JhO39kQQ6qsctytP
jIl67jYkl42gGlqN0mqCelnE0M+GNex/MHAdBezDrpHJvrSSden7jofjCDldrd1yHN1qf3PkQhp9
xfeC0pkuiVTHh4W1l8/l0GYgD1Wl+zffIYfYEk9iXH6Rvi7tkwNIyZ8fJek2gVtRzcrpgre0bsur
HdYlwBke8zwEXM7cQHZvLtqvXkHxcRcSG6RuJ2TKekMudYSc1bEbZlEsEcdceafykTS56dbE1oLL
gdcmR4wkibKYwmaiEd+EpMXGDCLqKS0o5ZSAGMNrHhZI83gOSqHO2bgJKD+5VBtakPrWp8pHqQcr
kNTRWhj4VnQ/nOBibG1qkG4MKR3j0KMGLK/17DproiKoJQ1zhtACDwbO6Zr9WgGmprbFrwNtO9Kq
0PzWb1j9zJUwv3bGIr9TZGgNKZxXaK+eV2dZx5rVDCGFQXT7u2oraWgnKk8m/yohUcfUNFzOB4Kj
leKvzPmyXuY0O1fgrnRawoJlGVcqCuTM6QC/XR3jKgkfCt7DnSjvdl7dZbsmKH5fyCtJRVqQ7JHV
WbD1RBC8296dmGgHHYQgxSbHTh1JXJjKkVMXVxPFtVw8pcLFhQY8X4yisJX6pZ6c1iicOBa5ZJXC
eV8NSh2mr8QEUTSpfQAmOpr+bctzyySNEm955rjQX2w23cSQJBDOD0YOek6Jw1WH9n8esvcad920
nlSSxRzIJKRcTFRyeI2GIvAmQzMtn3fcY9Vdm9vAKsrbJlztqK3/3ew6jhoAc5POy2i0NwbpEY8h
hpRM2IadFrvdAqrlX82o2ULgMmUyWG71fgYZ/Y+ESNLrkSBUoGOvUlC81w1u1/e+ay44HXga4/Oj
xLpuz4w8OXznZq2YeFZOnZHzPM9IdstoI524hj6sLEl1oaoYRO8za1g/VWjXJRxo8yINRciTGUzQ
fgLZEh9f0+S+xbCOGLCeVUO0efMb/KXwvqJuOfmhJrTe8sVP2vTzjM9NQIhw1SPNBagM6W7M6vmx
TEBKRk5UKI56tqyHQo6FuAQULRDVMM0XWmQHcDwv8DSQJSTW9c3hRk7uhZoMrItYqtQTaeycN1t3
LLuBwESOHKGlIaHbanKAU8jpe+uzvqJ2p7EgczBSyzt0UFvp4n35QdQfFAEuxbwAdw5w9KUE4jng
3ZwZ8W+ffdPhHHiEeHaDZvtN2NtHM0xyACoiqmFGT1uh6UZdQ2SjE7kQrjClYD9ucMuas3lS9nwa
FutdjQHPX5nxdDaWaEOg4RiLUCLZABQTtrpOZuZY4+d9DhxCuz1mxalK51quhbNLZLvdXZjeKrgI
w+XTT4YxUOphEi4eXzWZRqMJJXFQ6zzytnMGNHaUnv+QLRito505jEM1XzQK3vajfv3fTKfk+B8Z
Fhd6JKO+dOiaBbfBUEhsTPnf25xeQFYL/QN1T8KKgEouU08yY+cJ9rsI0rjReKWKJjMcj85rkYzT
1cb4+7tgGpVnja9qIsKOf+GMToPAQ1hrKWTnVtmfYRGHAib/YHoZZ6HJqShvbjS0tYPo+Q+E8ppL
l+lxkQotp/IF7aEfb0Tiq6PJr6/cl4Q9tJz3qFXnTOSblUxE/C1DTuDX8eDTFIRh6AtCSgp5liSz
niSufK9XjzKPoCV6yGyvCpvNur2HU+M8N7mOpuO+QcDck2mRs/NOt0rKlIxk2X1kdIqsnWmn3Fu8
GMvhUyF9gGG1Csewxl79qXj4RnT22OSKl6KdYLXWxpnxwTkRcTGbx9xLWouVCwz+k6CZc+7pPZGW
NBIwK4sQvF/TZdksJXDiQXKWql5DVqcy82HJnlzvxc9g8Zm/BLberM+TqNJvQr3KtERjk00OmMVi
FSZY4A3jAj2vXp7Gt64hU1x1ne+gld0yXHhPIL1+FBC1EcURp2qUsChmW73/AXW6ekyBl8Eqlw71
2K9j94TyNkNBP6pfeRDz3lzWH8m4UO1MeZByDSjvI04ilL7s+A09mMyhFAjAws2O85zpDXinTdpj
QnAAqdzAc5LRm8fcguDuYYOH88l/aRlrJQEmFqjFwjKyuHjj4XB/YDpkwTTfTFuPCnl2pxS31yw5
/NNdZa5dNFjN7np00R2W/xNRG09/Rx98bmhwrPEtBR5Umq0fkP3DLch0dVBqst0YyAmxT8uFjJpg
3tjaZC+lrLOeVKmoNXNTpEIuzITHRqdIbib45v/GiY17HshqJzb0P/beFCh8ep1vXCWF/ESvWvzc
RtAKj9Rwp3DxWURnQrJ/mX11ppOTPiMWvXlgGFFmU67MiQfJoy7kBaM0HAG47dgib5DFzfRM5WtS
kQFHBG2lkpPObnRQkBQB7ge9VVX5jNTwsmgc1MBMfGGfl5/2cCyCv7Z7V+r10eSteD89/i0cYyXb
sKunNAxO/VZhGexrglsqY/xZ5PrSUNoxzlXo6gZbYxH9a/T6b6gbBkic2a7KbtT/ECn1P4barpAu
GK4e0MZPxI/Vf59gMtxTH3Cqc0pWHm5Cpp0Ele0xURy3uCncezf4H3ExCJXHVshlcm26nok+b/p+
tYnFElYJ2gyzw6LYz6omsybB4VDrcSY1jGpU2Td7lpF6+mE3Dy/I6GQ6VuqZ0XziGazxy7PgAMwP
T8qi3NonYFI/ayL/fMQPv6PCLcbSVRT1rFuO6fb24rUVsbFeols2Uz718Q4LUQNSgcPYA5Sp3YOR
o7rOAzJWsKzQGL5T83pmTZnKcidK7kJDt6g1mF64iA78FQO2uTonGSFjiQ51kLLAe9wTEWBGnT9j
/G8S5CdaOlB1Zol3oP9tAkprszkchsl9vtcVCto8HNU0dBKml3rl1MZHij0+XVxB7bhTHQYbfINs
PLHxRWY9F+7bitcs/cPNjrZkD6UHRkTFjuCKHFTEjWWEzJ5q0v2Tkj84tcCOor2gDnihbi42VDd3
BBYsJsXLMAAk2Y1K7ZNlGeXS7V4fVasBulVDcAl00Es8Ip8Ig7XTGS3IeU0SSYQl/U2j2fX2v2h9
RkpEo17BK5ETUAXJOCkhpC9oAgTKShmCqxANU/eS1qUmpvGYDxAnzH530yo702mqa9oDigpu8MVd
OEE3fMGOcxfTb5Jdxc4PPecZVY3+zLIbrNM3Rtn4O6gxxIjV1G+3xRYozp00XII0wkHmLSknxUae
oSgdxrAt2msJL10J0kKz0hduYgcp9Ydk8QvbsJUa/Fnr38uVeCp8JQ7D6NWh3B0mR89ddOqqGl6J
5iqRdo0RdtBZOysm7B3qUgxXqYzMl53R3T624FDpgcFUbRcnFRZH+H/MjvpzGMRfdJmOnRR3pdWR
KR/HP2JbtN7s2exCJwW/ds5TI/fkQ0G5TGSlN2R9g/cfebeDiSMIbvrnPAJtuChEbfUxJLtTkgk8
0PIwYFl8sxPl53Fi2hpPkcXG4JkP9MgAAERTxQn4eSN+o9OmdiKFTHSYjVpAyteQiuCiHqFFPw07
mYLHJjXNew2wIJypDqUAh36nYLhEPoifzuJoYKwiDZda+pD2We5nGIFUKLEN1wpc2zy/xf74guKC
c/8OJnnotT2yC5seXY8y+SFqBWlYwrvFxXKJ4Bmnk/U4culBs/6NGF7njvCN7U5NLGMC6Ey3PPvk
8yYX4ci/rQC+fVKK+JQSQ1XP2iqwvPYdB9Gs24Je5sUNDmKF/Lqzwh2GGPOYgxUbFFF6d0b3nzXz
ky9mq1GD9wg7lSlk+dXAz2qhJSHAYd49yDu7E3a8kHLx+ZscExbClAhz2iRRWmGM/PjWOzjKvxZN
WqyQ+4ZiSHE6S9UqzAZs6sVZozKQRgg3hCIi3lAvG/afS8mOj0IKZEcOKtTgevzY5NJGDcMiy1ME
EY9VzOvWf/PMQI7yXSHw9vGo6iyi4QcVWXRjC3eKXFa4Km0ikL88mEkCEXfRYRzHpG2ky2InWZzv
cCQGEh60MQCzzejOJNZ11Y+AdNNdE0sBzu61Nu4Sxltd0Fz4zNJw7P4iCRrjZJuI52lHAsdg/oaF
scUdQuphYTQuibSIwc8X3DVSIm5NaLIXDgFt3B7Es/NGuDf5bAhD935Ug+bVIZjlfwC6Qp+UXM4t
e9R+advH1RrZkEkgKtdq5pDDBWD1CkGjOkUvBG49iehW3QuP8jXG328+LUtekS58UXpZcpPPVdIJ
5pU/8MqHTmhIQsHBuZ8bdGeSIg5DcevbX5byj3acacCJDVvdi4H7dsNbK9UogwmDfoO/vP9Y12Hy
/5RNK5OZrjhL7XO8Cxdw9kyyfBRg0pVJGnW/Pul+117FpL4wIv+xwUE0Ll4DfytGM+qdz4LDyavP
2lJCj+HpuDQlCc67VBr7l35pjmo2oXHdYjZK4pJsg/ZoyVuC1lBlpO7M684ZZDmDWshg/+He8BWv
JffVkULxim38YUc3SWhe6YL0sxYLWPQXYDdaIU0ZcemoHrP6NkKHufFf02FDwa/PL3hOIe10ruNY
cP7fRmrko/gTBXT3DGbRxb6Reza1zxlNwBtbj0hXya9iTtt3dkQK8CeCUBoCB8cpnIOEuYQHK+my
n4k2lb2vmFsGbxqHM2hNlvy0tjGE3lkaRIDU7mF6avVuxGyfWATQ+19jkMewpNi7b23BFlVDwBAG
i72J23t2a9JH+7t+H79r0TB1goVSsdsCuxUOhdMstIRamOfqLgvOGtYmdCAXnkUAN+PWsShfwXg/
n1HEtSUp4i9Ctpquf0Ajh9hkPKEsKwxF41Lg2FG3x9M9zd5u+uHoVTBYZaOAmwKnpSw5tLaFyiwO
VzVoCS+udDht04ueP4wtqkKA/pE6jwgI909RyTboZ5+zQuQGQSbQDdB+3K9escnTEceJOZgcllkZ
FfqQB5JjBrdLr2UNaKuPD99WynUwtZZSlHvqz0fWf5qC9w25ug9Bxv9v1Nh5oKtGrUkJ8wlEE2AI
iRuZGmgyRQ1s9yn4d11cLa9JEhKnjj33YOFZZgtlCfHVPS/TZEbC1caGLcO+h7N+Lhky6mOEnDnl
ZG6+B3LHJqnkKjfi3EocqUaPkSd1uCZ5Ydr2JzkBBofHA6WJFHMZ9zh17+BHGQz+oTtJ8yiPtBKT
9XHVQlABy5CRS0C0Makb41HT5FGB7lfsmgA+XfzfUxqgEDldrFNCyvJ7b1FJVrPOmG5DuWLVcsG6
AV54GIENL+GqBXRIPEx0AEsZ/BxrQ8xeQMHi/C8o8K/0sLwIsEytZhkAV22c9PnHZngCs4whwH4M
7gI01AJ9iNmSpouxdrk2hN9EU4CkHs0ADGfdFY9PAg6znrtXoGLSQLOB5Ig3ipdXkg7e+nslWXNY
E2xmqxayiiqClt6EEfewYF17+iBI7Xn9nItHOhTbpv/Obij2ZqZSbXEL9/JEmyW766Y2LNv/DFAh
c43XEJt7wz7XHGM42aeXaLzfdRJS76gMyzwEd9cWqqiKHfc7jdOGbaeeGE9F+IH3TAobaXHTRBUq
8wUOKnryPpCfuAu8PZX6yiM68XfHrPstvQx+o1cvBpPLZlPA2geTz2VI7JcnsUvYhVy/Q4Z03cla
Stf/IMkKvKfeJWXLu/+sgsJcqFUHyDkw6HJO/fGcf9J8eg5/Im0CjU7uafdKG8WD9UFk/HG5ARZp
xaFuTrB1V5jHhEzuXmX6x/fSLs+hqzQQLNxXx2hy7Zvwj3BhOMwHVT0B8YzxQ3KbcUAT0J+xophA
96Zm8TkiSUenSNUFtbDsfydlHeaX7aHs3mB0GIwTYZzhQc2b2NYROt7+zAAflMP92sQBPbwSkCLg
lcE1Qa3IRMXoAkRWyThBbRnM9wz68fb40Cg3SzJ2Sp1F8l1XLKLBgYok2hMxw7t5wMHkluB9Ztx6
RRI6P3QLiwcp/eqZDH6sMmYUF7BHnj5JB64/6O/4bqCKYcb62bAggNIfedm9wvyr9ER1lbWfjNBk
QMb2YEwT4RCLLymKfqjFWS7hnCytB5MU82q8mmP2natv9lWTvly+oEhY+HRvR6J2bi1CT1S0Sh5C
iEhsvuNq/4yxXMSBru/UT6IS5b316o4Y/NfwZOHTY5PzY4yDQTXkTJiFqsIlxYomiWMD2ua3zZDS
fQWW2JCSSpIv6HrlhOK860FKeUvPBs+uq9GQEc6a5w8n4h6irhsYZ8slO+xF7xqZIsKUe8CoOSPS
Y4GAuZ7q3sSt8I1XISCE5gZfrtXIuVeHEHbzodLrKKMAiq/dWcwH5+ohwWmaMOKUJypApV52qVuR
Ou8TbLnTHfxeA8L7zt/uVqORTt0vk+7CectoCFFfcTPlC4vWvK7H+RoTQDKC5oGrRvl+cP3AbjNj
n4yx/oG+TvaGfmbJixOBkEBFwzEpm2rGo1i/WJXH/xEod9bpdnAETYRQKZIK10BweqE5yv6ppSF1
r9qA7xNXEynnQXjkBmu5v9TDdymnX3eS4aOlAcFWNE5yJImDDe0+ZFLqlgTEPeSkUVpgukaHc0K6
qpF/bElpUmx8KHveKETGJCbgiySRjMoUQibQF+dhGCSRTABcqRcRNs2/gRBcIi8QRccW/CUz0OdN
VvUcKjmtqsZ5O13iI1hjFfTs/qMvvtCLl8FJG8mkijjwsI7fZgxpT1xpnHVX+7/6mj9GIq/KH91X
6xyOwJE+DqKLPAobjNMXXlDDtmsMD7Ub4SP0OxG9lpNIDJzoikCcbzdA73iRklua/80ca6lAAfGx
GGarxv7gyLiJwU4URNkcdobNqi5zJw9X/Q33ZuyhQcZCLwR+/zjsqsp7UE0YzWnZhaq4v2GMhyx1
+SsU/hWGcz7hwGyas9+vZYrcVm2eu3FhI1v+4B4NBe4NTdptUiEsJIXFZBJLV6fUc3Zjpzsq3xTt
wqeyfE+G04E38ViPPN1x+quaHpfzy3M4dUZ1ko5erU+xis77VnOpjvdcTzKB2zSQxaMXDPA5pAVh
ihxpFBCYP6mVaXhmlZe2yhLLtAb2+qiCL7dN+ojGtc3/gm0H17dhsCoY94Ip4bAun3JCQQOSVNsZ
BZMIqyVS3OPyr9Kqm0Ch+N8JMwmUukGo5JDjknfCxB9oVnMRikNKBsUg4RN6zwmZ2d+8bDlbP5Os
rGV3iMyDnLPFpdkq5bdPIuhTPaCjSFqYFmK/gMn86suYC2VYq3yOMSEM4dycKhTkkPvDRxtu4pqZ
3o0NLs4D3XODgO4sG9eBgDFBb3F1n8AtJB2GSIKeD4twlGDht1tW/xa2KSrM26klqr83e0d4UtLu
g4QZfS+9k/GrGR/ou1jay83fYFDDRQR80DjC9YQr6LwzOmGknCYthhiUzjhgRq/NJmodGO+2FnA5
b3dX9ug0HXc+ejWUq9U+hmkVxPuA8aqdaAicUwS8U7Zw74GOsb1pIaEhTo6ieW98iG64sKb424S3
ku2eQg1QLtfnATzjD6Okpd+1cNH17Qdph2U2Ej5Klkm1FQOX5TZP9ctTPY8jmtAXx3PXwaZTU0wR
BV6XUyKlqZpQLYsd4Fjqf/LKKJoO3ro3v8ff77s3F1XUQb6Zx8zgubHIKpc9raTukfs1xwUrbJ1S
HtfsxW29/6Hh2tglhtp99R9iNwZPlN786/wPdyeOV20qiweDnFIGghxb/9NTjReibtkoriRR42nM
VE1CSH/5qC8DiropIBZx8WNZtN/zgg8wMiohjbvwBb1Xq11mvm6xRU7KiqKzG2akLbm9q28oPJka
d+nQ3Pip67vEp9bMQ7zdR/2Y0YKieBkSsEP8mUmd8MWUW/N23Z0lg4vIqrCSThYMtwf24kDslzkq
hNVklkoZlvbZ4bKkqhCxRty4rlLxAsnZz4VrEc6eBoWVywcibyAJrSxU553sXrDgMfV81pI3NidJ
BA5d/GLuPGZR1p/AA9QpgiX0p2uA4A0WGB081yhFQrS/7a8VdPvIMWaqAFge5bPuzFpAgv/woat6
cCn+6zVwwhH7wdcxbasdw8KxcLfZSpAtjhJ42euqwV4CslaRi7RlySim6W7ALBOpSt41FT9oo+9l
xzhNuG4IAuLDv7p1XVwZFT3APRfn36AyDtJbPr+YyzAv+BzG9ONG6gCthaMcZua/Yy2VTdlcSAzo
N5RKwVqJ2UpAHM7xbZPHZEJjrrMfscLArHpeaXqDBd8V/ZHo2GXnMXZxQ9gNmZc0gD6+qCGBuCLl
0/6Ce3y8mZHXTPBPpbzIcx89bkCHbaPSRrrLqO8pIXb9WsscnQFISuLP8Ae1b7LrGGEPVSyy9BtA
WSNCv7s4gKfx+l97EFKLKgTGeCw1lJP9MZDIakbxdkMNPyS2jDclJVSCLUEZ/9+yrBsFdZ7DUMPE
4BsXyV3PAAi4v6DuIuDoJcelaUiPQpnEdYSoeSvdNvMBPJkXdk88Yc3S+b971yhUN3t0jotzvPs2
DPbreIrilhBmxG7yRpOszFVr0EREmGSI4+I4YfpieJtpNAfylrSLkSpkr4fLdfOiCSvd+OpB1NHF
mWacdLTVeLTAvREbDQrvZZw5gFTjaoTbASoz5k59sqS3Ss1JPj1Jd6sbp9JZ0szkS2uzS4uuP8cR
n1ETdZJRZAHdT5EddasJVafLVGrMgaB8GSqPqPBjMzh07UBCGTIxUWy1Gv1l/I1YFV+mXsr/24no
WjD5efz33UXMzV1xSiKOVP63oX4R5svplP6BV2oCDXnH8i0Qw/8gUNoJWFz3F1n+ujzk3yfnKMM3
5+wYFz4+z2PexiiMTSmdP/ZiqM14CGsT/bPT9NItoq++pXBX+vbu9A6U3Z4IL5PLFnvSAxJ1J/IT
rbF7RqKiJ5yxCN8GpQ7+qeyTWnH0NLXzwjGUFYlF9Sq3H2XpgTihvCyf6UNDrsrUHgRZGYhw4s2r
Ra2TmLxJaed3W9TFcFP6YFo9IFoKL+vigvbqPp+q31Um1GawNT+z/zi4Cu4rL8wRnGAdwgVi8hdJ
wzQz85Qm3sScDr7cR/2l+sjl9EDFw0iYaE4CulPV3qDStfKQ9c6YbbgEE/0PU00Ex2yxjym6EGrZ
oadO/oF5Va4+2PTN+yXi69tFc0jUyW2zKIUlOjeI6EK7oBzb6VQoQLe9Yk3OexJVbiu0a5geDGf4
hGmHabDzKWXkdwAlA+U0XgRo8Fm8c8awUgMjHxDDdHPkNlztw3aR2eRtyXFuSV2Qnf5ZlJZm7/JG
x94Qq+/KabteeeFSgN73+aEzs7qz6ZmTf6bcSzreEDOxtL2wspTar/58awseLqG1wG+xXBE9k42e
1SKUXy5MIhg7OerH57YA5HCcZYw+T4/LOARvYA0eSmY/hFN4gtC9c0xdIEhMhAw0tTUFw7aqtAg3
ZSHRTrSIlfkycUGbIPg0Zg6mZPH3VF9Q4ZgMq094Hb2ZlN97grZx2IqGYZLrRyrM4jgHmvR1Y7+6
BBbMVDEqydL9OJKGpbO3qm17IDmBRPX46k43hCGN6rpK/8IRzbb3xo+o1ateUvsaVpCx+ENG0VwQ
x/8kS1UUuY4javBrC/0Acgd6q1cl9AjPvnohA7Ofm2Nw7DbIegUlpkXQ3sHo2m+cV9GwLPRBaswS
LcvjHdRfBGlAmMzTy7WIYFL8/2LrI5T/MmNk6L2Ims3j9XDRQbmsnqLc+5hAYpDtt1519HvVhp2P
84DfkV9mk2aJkV+DDUy3yV1wfEC6v6R6F8jGj9l0IQZt2j9E4JgVawxTYIDFWBZRMZv/5sroChq0
v1B6NB/XYpS5TubYyw4HeNuVMhcnSI0qu6u7EkvnPMeJdyzojAzJFs7OlpLPh+WAXsPn9Sg8v2+h
WaXm6/YNx1yusBzNM2cdSMwejshQ29oVZccO7kBdcQ9Dwt+4GT5e4xomF+cbRTR1tFu6biwQ3nXB
kzdCbkjLpWx3GgG6hPf1NB4UoT8XldKhZEB7kbg0d2l3O1hlDIDqQTYkKQudDQgEACHv8ft6zDvN
LPD8najDWT/j94F98IacRvSnadwYNtc9WrchVZ0ICiUY6tiSh2yrEMH+Cy5Opqv1j+7PxgH8CrCL
dpJzMtOrrXnvbfl2nAFe+CxXJn9JV4K6Epjf+uzv0ncTC3797jizWUWXr9Cn2p7jptR8Q6qQaJ7R
Aeslc1FR+zVlTVdRJYIEXh5ExkfgmBqqSmxAj+MyBIcaFe2FJYgaevkWb9pOYxN+DnEXEiUMMK57
pS+adIkfHxgoZ6X/95SAs2uVksXmL4S7hWrILZvL5u57a49U42AQFo7hiJRG0YwgV8Eg3/2XrNOc
KJxzSNsftbJgW/emxdl4zaxluv+out4vQ1l6hyKSFvxD4HmcRTGfLFXU/fawtM74hiOF1fj8279j
3aMQR1nJs3JxBTEmQ45tKI1ky+ffhHGjEoMD5t6M64tCkmsOf8JEL6QIUIft4jBYZTGukQLCq8bO
Ei0a+BN2f1ys3xcyzKUSZiAEqklUY5RsgRxhqRuih/ortxVMn2wYIw4UKQNgZmPLiUft8q5E2zlu
S5HXTv7JloUXC5q5Wy5vchpS2p5qpCn2g71wa8A66hlpbCtRb147mrjnO3kpC89HI5z0HxFSO8Me
koA1TlRPUuxBzAwuJPRfh+mFb8uX7Qg6A6eM/mYVDZTORkcami5nvEw4seFukSAP08LQKnmrXgeS
tiT15XccYAPSF06BTVESl7O/ahSlQy09pQFvLDlKGFtFHntGYa4vsNOMcxTn6IKMCCaNF2YgKSdp
qa8l4F4JYNLV6a21BYpxE3FN5vdpSu2YPxFQeYue3MZzRpIISVf49qBoxu1JH+eHUugO1kbxSW3y
himYLSetv6HF5I7hhyP2KP9C1EeuZ1avWdAM/ZU9o/jdhphxIDvLEhY5+idpINp2eZeX7xietJOH
+ZzL5AMqQIiNIozkYmrCgCDBw/BxoxI0LGbXFGP5gFALgWxxOkZHkEa3ImMHi6P4ZMxOpiRTfylo
dvkFwa9Jq8rRjsbdDZbo7bayJIVuGUbU5WhufxbpJVZyUh0n9LwtpgG02DVT3NqLJrN7l8FAnvhK
iK7nPwXVASjo9GCJ7LxHdoJenD8sU8EWoxWzuiwrHQySXS3pYy8DW05GAUBD2mhfTXVLHezjkor0
nbNXUbeAGaW6/D6fhfDmmUo5yOJXFvm8s9QPShAgpImwKbYHK/S2XAEXjRwHvnsqSSJPip8atl6E
uK3ZkxE1mV7uylTI8C9flJoWuh2/+OhYA/pKuLIr801XvIhWLSQGz4oQXdlnj1llC85ivcBF5+vl
SWaAOe3UF18806eU8EdbhtrCrN3QS1EbimsX9OV7Cu5bXRJJV3TBTLEGK9qq2dTKe2Hd/mgICz+2
hqUnX+pjxrbEOpn5BmWKFWGA+ljkNikaykb/7T0jf4A/1Z+uBnuLQuRKC7SffhGHOQibk2H4fcK7
bLO8G/FcIcbmvpEGcoJ5EVPV38JVz2/WW23cJVOt9+9Ke1RfKZjBUBj7MlfFuxrXj0d7z5WHQA+P
H5MW9ZcRDEbawjrHympSpyVFpmHKQmq3nH31wltmtQ2P9KVaiO0finK32GSoYvm3H/skWPX/lfTg
5QXY2iqSWLStvmSly0oNs+SXmNxprtNMtspH4uMgO4G69TfH5jCSlmuOLNrAykdRYXX25JzvyRz+
z5BCouIFyjd3rpBwsrI9LkJAWjebXErCiQ9mQm1zw3YOGItDFXyASdnWB060nTrQw2KDz+ZfvVMe
bBWUUEwCVe3btudo5EP6zX3e66EKPRLIC9mouyg2HLNxCnFhxWxSEjzziIr+1HMoyKhVXu0D08Pb
5vGiOdTXDzJ25GQBBm/Cm+KDTSHkDjFm66OSJIJlymJPaGRv4gNQ8MxOoaveZ3b1idaH6u48yuHV
WuUKBVqzj/3WNYgQRbpVV/dfZHNDk2sqErc/1HF225pthxxCAVYlLHXSE7f545kQWkXYvg/umVG6
pB52aw5dGbu3pryiHGz2Rox+m5NNmlSUbYxnZNA6ilcZu3oWCo4RJi/5bPvwjwB4Y0CF8dM5aH06
psP3azwmQDgDt0rLuNP6WbyupPf1H9HvOC1MKV4mrGF+fIlnmZmAp2kuJKekP5CY84/cQ9eAllIE
joOay47pLEgPmedZkZ/VhCcQamajeh6vMrtWZolEzz+DmpKMkOTU9V9x8cQICldE3HeQM1yiR+kp
/nqTjvw42Bd+HQZxFFGl1TqGY6X8wxz55/UqXeJZmQbrOP62ZQTVrQ0v7tRDeThVCIjnvHhfu2hy
DqeafwyaeZiC/S1ZAZVoZNTJdDEtC9yltAuwE6kNBFJD9Q7b8nPUfp56DjUBJ/efVq7RXkjI3ea+
6EYTAgISnHl/tue7EaJ/ptpD2uB9k7p1UWmraNXwKJ7ElpocpI5Glyui8osFeNlOYdWU8+DTKHTa
l+jy5mKFNmgCstm9OykrUNDWt4dP4SOZYoLqdjhZKFIuzyjPbjMJ+wKCiaoIJ9r5XITamY40woM2
F8MJle2nEOBcKtl42r4ad/BllFenWwrTtAmT/5QLCsX9MuYNKSD4VXM8xsF+WEA/QCVHIk+a/4g9
ZP15rG/goLTSbrDZZ/VHlDLun4LIAx7sbC0gJuApc7faPYqzXd/vK1uU547n1C3pMHct2EzDj272
B7IgoJS4bs4zlF5HRa2LheATrFUjHxJV4Lb6nj6HTSw/YZ7+poN8OXSWGC19lll5XRqXFgxgAvAT
2rtHzvjihPWONbuJD3+L2cG5NcsOC1gQ0EoFlxrsbvsjiGUSpIDDG4dfqQy9TIK0F6kKoAWqs2m/
CtqAqycBahitG36gtMMta1cd69miKoyJPZ2jTarEaHAOcdmQdmzZe3in1BHNziUPFYfIWbLoAvbM
6sgyHFF7KU9msCTajnUtwwM2gOguhh9sC/iYwT7Xen6osrKADGF+ukhzlBKrVeI+GYGbn00inYjm
cIScICb80fUR0QcKI86VaqjyeAHlWed6Ovv6VQXUYWs3wL2ONXPDzFox0DKpOwmtfJkYxtYLMBBe
WDR2o8XjJaDCc5VW7aMfK6/1H3Wf49egcS+9EESbmm3szq+oAzHGpyJiVju0YsQKUtnyoWCFUmEX
QYqpyc51pAMa5mQ7jp9LkhmTXimWJNDIsn73zCqIQrjrpTeLlN961bbF8Hoq3kh2bRvFINGkChtE
5x2QMhmXdp1Imu7x2m3nl1yX68oIdZyEZemV5UTMIiCB6puBVnaPMSW4xFZtqOjYp+pakPJ8NIDK
CLsAScUBz+Xu1XWq6GapILg0ijWTmfzdcB+NFxHSbEvXeIXMcjNxCHToVVOO65e1ssKZ4lRHMt73
Ow/1pPYQE5nsu7SDpDUXvKCTlDY/1T/E1hj/u/kywbf7sL+bfyd4i0Qgc1lRWmZaZsmgcw2WRfOD
7U4djjlMfOAlaS6c8M0DzeK5NoTNftFaFfA/avU/Z59AX2rQlYTGpNXwcXT9+xzYFPfftlNKaXNZ
jXmTswfqQbVA+erKf82PfxgbjDnjdyQABkVot6DZRLo4wOz6r7dXO7ipJgwyfWwDzb0impOxZ40m
REOzgjlk6YZ8AW2eo8HeSIlOVND/zsIH+YurNOfg9sg6gslGV5n52x/MH2GoQdtW55T2IV5HOR7i
HHAS7Fh2JJdklnU32WLKVtj7UkpO4AwwPQPu434xlWCYS6v5ud7Bx99oCwJK8f/itm64wcZtFu3c
ReJjMPot0jMu6Vj02khkr7y2gOs4ANVI48MeIKoEqm/ESCh4UyR9PsykE3P+DEtd442R7kYJiB4w
lVoQ6KomEZ0wYUPotyiaVWg4ZoFgFvBPIxE6nzipLPnkZdk3GEhkmgmFIW5ZYCBCs9twQsBkzdPo
QMq/cAFjNIRx9CTmn/2rFJ8VKLZZtxfoW4vEVH4WVnwQXAS6EgnsjRArwlNoto320AxuHxPd48Fa
od4E8Z524f7bmB7p8NtNOFC80CarZULKg6uCl31FwwgdwlLjxNlkTEcytD6z7CjbFlekXRInKhqc
WqLKkX99EdkKQkQfRvnmiczuKsoDpDcNFUQ1gilX7lqD/+dJTr1bQi9ybIYSiwkbhsRKJ0S4v+sf
pEQ5U5xvg+RCXJSEvO0nLAyfisukmK3tdGR71W1msF0APnEcVccnv3F1nz7gG9dL5EYEKQ8xtZ1K
terJhJbixydRCGcXEszWyFa5AQwfNwPTVLsbzkNrNO1OfNXTdsqlP3X9vdlIc0onC/MKiOZ9QN3D
0tsTdf+WyhbtFk0vI7L2WQi1S3YFj5PZamqrz/g37C/UlTnwG+HJ4YsfZB+3WpoInvippPMejrxt
hQo6lHtp69wSlZcj3phzE7J2zSp6BwdG5jR7+aLP++xaSXzkzeNheTUP+rnGWJe694q3vMTdu180
5aBL7Trls2uNHfYo2K3C1Y/aA4xFnjsXsQdcs1Qw+SELwtnRvSJf3OOFoK37i4Xy4HZSzFADvcwg
9KbRxQGJeJJ9kYcn1karKdeSp3+6rOP2KB+PtfVYnuk6+sJY183K/TzCQ94/57pXCC7ZecrvhyIg
DAXTM0fyBiR54smNkHT2p1S//VUB1ZuaJH4o8LGlTlTR0s1lOaif2vLau9bdBEjQPUiXaUzDT1r4
dj4Zhp8o33x0ZoUPL8CR3HfAoAOV5TvDX1WHTYq99hYmx6csitBFnDCcHicDHRMEITVaAtt6mTQN
ZrpTcC7bDH+EjjeNWjDZWWV3IC/OkVJd9v6sXiZ9Ot2BSmjEU40oq0Q9pJouWdQm1aVcDvze/R4s
dN3KzSIkE45TAZyotqKR7Kp6F1zyuwIGvw0JwAqqSpyM8PfQfwwY7YZlNVHVPnnoJYCHyxyB20/+
xwvJueg8JIGYKvqlWDLFFOtFz/CQ+G3ILeS4zYq/v4nBhCUJiv1D1YkVyj8GtVtICUv24DTn3G9w
c5QSM2V4ltVw/xEimJM1Yp2cW4NwcOti5NEv2Sr0U6lXhJXNg2/tR3GJJsyg7FJ+We8fgx2ntkvw
5o8wqRmLryQC25gB/evjtBsoZo0+4jyw3twGp7bM9Tr1D9dmU/W6/JbJuVQ5rdHktKKuEM7qL016
uhlpiUE2mUNdRE//tiFLjsxPvAHRTVOpE3GF8peyrrH7KMuh6oU56JnXbnRFl45eopCNaIKNz0dS
IGkWK4/4iMrTut9P0KEui2Ou0625Y1Kh2pSViyC1LRNBpx2xRUyrgKdKar5omKocrO6/uBYcelO/
AHqBElkmaJ/kQbZ7Se+QMRu7b9FgsXTgOtBQBUePz1YF5P/WAYEVj+KF6VO+yq80fz3aIpvf6THq
6pJa3j/GnKECcs5ZogJceLjesgwzvdnoAQa05LvvuxFUvdiBa90wAAl3DkNVmtKTIWAXbAnZFVg8
3QMZHO0vpZgjQYWuq6PGTZMU2MZSalEnUSA4eiVgfoJHb+sdu5zjd43hazV9JTOlFONMxOu8Jb5V
qhD3sslPVa2qDztC5/tRZnCd/S4+d5X9Yzh/SC/oTzx3Vfwx/Inuc+Xfw0GNA9ab+GgUReSfPrig
OZ3YhvRUDD/6Ek61geAlVmUapehLx8HT3majbtr0XQq5btzZ+AWM/HERpRdkuYUbKgAu4rIjQjzG
wOH9I3vpYUj6kHKRH5zRn2qqu8A8BfAsjZ5ccVHAj/c5Jh6EqbdGLYtrGlgwgcDoV2A8KcUPViQo
LInU4Cm3tWhzskOXq1uWZRenEYWN+j1j1ckaEMCqPS7biHJGOpZF/kKIlFoj7NDrLUOQex45LLyR
mc/cwR2nVLDZIAwHYaVYV9t/DN1XUiWF4GZiuogW7CoOndYaZ5A2h80PiLMg5kDw6uMUS4huz6x+
Oy0QM266fraZRH705So8qztj6p/RXHWPVQRc/HPmMUlF9Ckn+LaEdwcrYwxLS1rVOTCaT9ifxckr
ycGRUqk75cFQxVzdH9L2EOihpjNJ6KyL0DSXED3B8KoqfZsQpukC0qvjLkHLyrl0C0o7eQbNIDjT
CSBLWl43vRYyvbW6x3N+ib1lukgy+EoCRN6rG9wDoU+XLbbsaA0D05Eds/6PW+L5mLoGv/aztNsZ
FXG7lbwIdustN2QYnroIxZqcNtMhWbTDLwSfkL2llp6ghtn/J11YRo2J+1Cb/uK5JrWoltfBHACN
hsrXbmwYMMYbMNNwccDiMwtZ89/XMCo6ORCmEsQAejTtyeK6Yrc9XKlk/Q0zz3Lb98x8u3R0tLzm
4Vxw4RW0PtoLqqJmUinxJYwRK4WJSmpmksJHB4AXCFbzrx7djPv10GFfDc5rRvonMyK7RWPTzJT4
ZdDrmaw9zMVWVRqHNJ79Ts5vvoAoDT2xmmPROfVfgjbEe/dUZGwPG1NjrA6gjBc8XKP1EhlaoFpQ
oc95R/N3kBG0mbdIVcYDHaJ0NBWnYoviA04cYKTwGBLTz4Y/PptBa4vyYTJjz8/aplTeAGAHcC4+
eIPJ3MCpVLTwR271eK2lDlGgPLbw4rOqIh9y/5e7/izwPdA3Vc8OtSmR793rWhgoYV0bZo+y8qB5
XklYgDS5ozQRYhy71PCKtxH3DAORtN+k/8ilKImt+B1GxLPqsQj+xirH5N+U8n0WVpdGmcW+px81
YyRHqD13auBb9paX5LryCyaocJrAk8X5mdfKqHf0qSlmBesg74J3haWUyMHMJPzk690v2NLWQY3e
I4CmgCHZ22K6RaYCFXNBMyStzUb4YT2JjGYHppDHscIZ/wnNE6PLqmfPIReHejsyE78jVIyGht6z
aDwEoqcpzx1tqlAT8qHvjuW0JXeCiH6LoKSae3+avDiux86laJEvqnh5KmePRvvKlFpLUucxVf44
E3vPOztsLmQG8OTZEAt2Hqqr8AI7Jt7GkIkZHa/4ib79KgyTuJqy7rdNb8rwvxHDTfdDdjWVfpDl
mvEIRCteivtL+5qRtOXP9zLK2f3xAtBkeYatZblaDvGB7sWpCYTHp36P2nf3ndj1aJ4cqUe5w1Ku
Q2yKohm4ul2oeMEWmlpanZXRJjGk138IlAuBphFc/fRW+a+2piOcvjJOKq3FmdmEutwIUEA5wGrf
zhdZlrQA3ZfMz1ExVxunWSykTb29qywV8mv58BWDabpOCNFRdek3mxpPUyD45wrctXYN8IchCheH
XxwmqIgeH3DA20pP4luM5DJ70vWYFOzZupPn3geApJkHLsRExWTY2cfuJS0ce5mYUZSvlE8jD0Ho
gnQ3NpKO1sJOxcwWnc7dPkPUNyirgmypanGqWlY/3+ltyK+tMXA3dmvdsUgUcCCoe6tW7WYdYMMH
QaLpCy6LhVfIApSXRIVBqeMbUjATil8OTHMNI5dryeSrqMaNG8nqAoT+7AzbCxsHOauNKDSR0nAS
PwuA4EF7TKyEu78dDPta2Fy4xtLgqYZS+JShdudQTtxouPnGgeNpSK4wtBmAg8Bh3aBYj8k/V7T5
RCCfx6u6CLXjklKpfU5u7w0VquUo1YVj0/zqnbg3JvPlDV7kFsbUGVkyxrUn/GZ3+p0/4wVELbbY
ynTa8MjyrK60Q65WGqfGHAkGZXvCAby0f1fCzWG9ivDt5JMn4r9u6nnqSlrcEVAHxAkiBpl49ooM
jVFREHVU2SUzDF6ekHSOeFDIyBnGBSCrpXG7OsaOOq6jE0mtU8WncEpv/2wxCEPRFkQGfU/+EUUr
YHw0qV2uMQU91LV3MHiDjpUZhEiKYDESj2+YDhgHstGFZ7Fj0z8PIjTHSmDantW9X+A/ECPnjFMQ
VaO5PnFgRhRKIzhuHtWWcj0pLSRvfdNWemaG4LG7yx3xS9Wq2bv7zgrkxivo0e3wEMQ7mzio79nc
MAqut5amG7Sd4PRxwPK/VNl2SnDIfUi6Joi5kNMGNoDIWeO23aUu5OcnZJsc2XRFQrv0Q5EF1qEU
oosVhzWUEYaJJVGwNF2M+jYsd+Zvv26fXSWWXNZP2WQPvFGPx0XJW9KpFkJf7uwN6otloHUXf31E
kKKgUEq+0hudc3I9q4/bE1a6Y+CiFJxSM8KdGYvVOotGhgMzPARfSDwB3icwJmK95M0NgVcLOXxj
c/0QXnRJZ2rfKUx4nqAbj5zVERKd88BOe1Qo5GinXJkfyqz4hEivuf8L8Yj1LdKjkiDkU0ciiR73
uc0WfKYXxp7i9jGLmu314B4uoEx29bTNORRqwFYM3fawfz8KA43dcotTVLRzkq3/X33y4Mmm+wsz
EQDeRucmL6Z8b+YtRkoLoq8GLBbSoOZFtDepsKz6xLNIVwP2iAROjbeLFcsuAjN7btRAlR0E/j7H
p0mUYs5bXt92aXB9EiQLYUDip3yLpHROAgokSnS4c4grVVApEpFoHV92+X2AwStZZzBeuZhJQ6NW
gHn4lDXLOGfZmivUzlvpSpTsXERuZ9LnhEhN++jTRPawZGIqrXD5VhNEnZRbvXJ2ADWIfMoBNdCF
huLAFYwdE88JRo+CaXGaiFcTvpfZtcHNd4z2rZULf853+AsIbZdB8pKmWJ1aSie9JOQlXpIMc4iS
B9xi6Bt/W1P1l82+7FH30dnJgtGbGnggsr7J8Z8rnobhKTb6yMytDjAJ5IVGpQ+/h2JWcrlOzBkr
+VHkQ72M89P97VzVKcd1Imti3H2N3nqlxTuBraNb7HiYGuDfdg+Q+w4n6JoRWmTPqovbNKz3QHki
xyTG4lRyuiVA1On6d4O044b6t1kplZAHSXseZnQAy1iB+q6p2pTebwJ9r6QMCXntaDv0rShKhQWx
z8rKa2xNwikaFV0U4xoFA6fl3bIVcsQJhuVKF4tNMjn9Bv8nrhUdrhcXzH/FbxHBfbaxbTL6LtqI
83sHPInfiHdArOPcEvUqHALynyNTG+yimN4X2TWP238nvfGFO15280nrkODGY5wAiaYuxeTInx6e
JX4Nt5REHju3iekmEbNBfmZbelreD+CezRIfpDxu8NBxWdIgPmf3YnpQCcQ3XuTuWodFPYsmLeFB
BDxfoHAzUBvk0VbpY9D3zoU97sZw90riH89XQj6GTdetgpKJFCG4KpBpgG0dGMgDPdMQuaYhDhp4
LFuFwTwC8Q1dJq3tW5BPVfcvs+v4fPfIhOn0ARCzGm7TgHa2YMcfZXw3tNOYfFIlwXw57AieCJb1
9jKGUV8GP3M4gsob5XlaNMDIvrdEbB6AYSdKzlbSDrmjFpixGx/lLJZKwYuqF5f3Bhh4e0PKCm7v
yZkAflIvFlegEtxXdpz5kct3VEHrMlyn149yc+N+Ycqa+xOSuB9Tj6WBZJqWURfNxDAZeatkSktp
hh/QLljjytwk7oLQfWCenXZ8e0kwI2bXrQS61OvQtl3HV63/yqmi6DDpmDGaVeTXN8uXAtRmtwDk
gB61GcDOu7tCt/10Ccts5vglyv9HDpbof3mg4zWMHYBvYm6nw2Pm/RXF13Dvuwab9RP08MtmLZ5Z
zDyx5m6tYGdrQZhIevyvyOKIl3ABT6HZzLwdbt2NJQfg1xsx7HgTvgtAmh4fmorjzxTLLhK44hVV
4oaWodV5o6J4u5NSmN33gsAj3hYDRne04CeEHAUlkY3CW24cP+gJqBZ8beJiOsvIUkk7UUX45LBf
j43IzOtpNs3vA2ZEcyKhVYqVbamdqPvgc9N+KjH0UR02Uh7gaHQeC420r3vBbbfwLMUkVMRdWNJW
rJiPiehP/D0FmdCLFUjrnZRCU0gwnGc7eQNqCSA99do0LH48TH1Em+jP3rwh9KZGp2DO/ZgEZ2DH
1dcj9JLsEJhryyzKxrbkndRvmu8jfNdc7dFrozNmvumWy/La4+Rx3irHwJn1eblIFdMVRWKBYyZj
qi7iRU+98jk2ae2C8tKu0D30es3L/2BDq+56GRFtUetG0COIf7iXYaYQNnio+HDHuPtO2LrIubRw
Nxd3Xrb1edpqzH2UgbJZ03MBKCuUKiiVYoaQVeh7AP/v5Dpd21lwWS5n+jVHhFKAwcA9Br5SB72n
GcMdhI8TfSL7EyRWwWj5Bcx43V9k3QPlw6+jNtB79RkVnJIlfnlDo0VF8icoB2F3ME5bXpTm0QTk
b9F8kp1NA8f5E0NUKGmO8qHeUgY50O1SsAiRGDrUIxYG4wbUitGtJqmAVI+iNMmBS3bUvRaCXrdx
aY59s68PU0fPEnqYu2a0r14a2U9nFdSmo6Es5Uxk9eOZcp4ke0Dtf6ndB2PLI7UQoaKO269+lrhN
4LKB/VvThc/KqNdtugC5VF2aHd9wSnOZvk3IAmtgW6QTo2N6bKoFcfq/LdukPAmw8p4js3H1C5Je
P30oIMMwiqLaBJqTbiAt1XU0LXa48YZo1Ii2mqaroFbF9PHxvTiXrNCnLyZCA4+9uyJQmwAMPaQ9
wYOaj9QxhHexYjByyAymWRLA1LYAFf7dDg4eWIoDq9FIqxNOeL8wTWStSU8ZGt2wC6hJzLg27TZh
IW6xPyYej37xE0/efMMghasSJ6oh8Evo9UyYkc9NftT7zy5LtnxpBfLI9EVzkQohSR/jHmRU457R
GUpXHJJX3uyxUP9Agnl+Krsw3vDC194FO3HEY89BgLIkMDyhySlULp/CzDVr4E+v9BUOn92rlks2
CmKIvdxMNpe1TEydSIaI8oZzhwGMDsagOAYu4X1cQ1t5VVFekGeLLmoko/cjUoIjOZunaNVXPzNl
Rx63PplnTa0CwIS6/9umYaxknd1eXrWDSkQYWnLcPrCyzFXh7gVa6YysyuiqqcSSSotmbCiY2LZ6
jdiRlVHlh8vDfxnc+ut4EXowJWsbaDW4++tLe16/qEiNya+Iq/Up/HMtBlkUTLzMJ7ehpVSiDj6u
WZxnNg0PgJG5kVSrsQ+BUzyHepYEP6gCsnC2y/Tq+TnjoPX5Vkxasom6JWO9C/Sy1dgxl4ddOs6m
H2fQyjxBpg/NfFs7elyf4MB5tB+y6GzhQsbaHfEu6nVKOxmBXy+mYJzt+dIPXV+k3QTMt2kl5czv
QPRslyrvNHgZxcZK8vQN0S2/aBPwc4nm++0SwcQZ3uGgeR5jP2lCrt07ALlhrzkgQdFs5SY+LNu5
HC09aOlJUVmnMIOKEEBteVitwBxNTPvCdLEIXa97Q42ET83zXXHsJzrfNFgQ6rk3zdRWCZI2Y4TK
16o/KyWIQSoghPy8Bv0LdICnLY6V3zR0D1GZq73L2SV5oH6K+xQ/CVRxOdv5DOmmSQyQGJpQ18sN
VljVWSFSeX2d3VPiz6tkFh/0zkKJBtaj30Xxa882jJ/ygpgtuZjmCJTi0SW3gV1ojdmxMou0nxgK
ea4ZFTnuxydeP2ZK6P3qotFDBCCw3DmB80zV25DA80D6JvWOPLSfPZ0CnlVVm1gQaeXIgniRQokI
x7Pd3AENyEFwrQaYCJjRmcXUmVDPkbKJbq0zsb6JSLBr7yjefNPZOReNquI5n/M5JHzzUq5gMEYd
/+31cRkeo0NS03UsnqYc79ft1y5nDWhzcEfaIegt+vtc5OzTTO0P4iiQAfEZxNnlUVoPYQDf3ft9
DkI99h8akPBfg4E7Vj8mHYTi8dpY1rD2j3pqbQbKUYQkEaMdtdawAOl9D211jVjMu+rKSXL6THau
grpeYt3cRB6kG3aDLfrcmqkWrk1DE4AuEO+E0BmEASmzUJ96mNlYgGgm14zTSlOJGYNQ7kmzWkxO
TKxaqojhOXFpSve5z1QUSzUMuIjjkUatF8OyQQJn1OGtd1/OfyN/5tcqynxGVFw0B9WpuggAuDjg
Wmtprg8rM+BgPn3bmg9ZUhlHmm9D/efUshv3KDlbHALtn3P3ofrNCnHzTQF+K9pWpZ3nqt6BLBP2
hU/EmNYS6/GofeA2lh1Mzuvw+E7VlQRq960UE9u3hogOuuEHmNrv2ENyTPwJzO/VVH8uYguMgjzN
QxU1JeKLtnsJCMeFdWeZvzR8niMg/0ODOx81jfB7kAogupGNbDxe50cb1J7o24MzhYJYE1zgZcdF
s3OQkiLr3QHxRU3pLKRae0P68SavXUkMCPqXHK9x7zNAGQOtFbVNNxlIDosUG3Dnulr97QSQontH
QZBvVE0hYhommwHNWn/ppkP0uA0Nt4XGzdlMuV8jFw0sEFnIMmHwILsYbPjZFwcgp1VfGAkDcUh/
GWcFTabnTnB6RTSKuCpf6CpFkWenO6YFNsl4a0cWn1NeEZ4yx2v/DPhrLvkPxfwmS8hQN8bCRBLi
egrUvmnxhsELgpitbYkfexSHN2UA3kppmgMJcwpEgzzuzyiZorzKnohIPZKEdq2oEFrWoPYkIezP
Rd3XGCxiSjhTDOH/+m+S1uf2YZur/smSW5eQ8CnvBB0gEtk1YWwMMWtQ72k5F08j2QIATSTefKNP
u8GhvtxbhGMml1TQ9hJLHgxGZ6trmVms2smzdFBA3Ilmag4cJ1bFNwbT+3yxp4yfVNfJUiOMGcNQ
0GRcvnGaNYYcDh68IuGuwc5lbTvOfyPWMs3Ta5oTTkGc8H+yN8YOllEihuVbRRsfddWfkKILNSZK
l7wuWB3MkdWOg9/avJRQIFuEvct0Pn2PfaCBQXQXxZY9bZjrDr3VJfN2o0wI6CEMiYbqO+HU8SHs
ThURorUisUwXF43PtfPptaHnQ3bHsbq91ljqtyVnxdol0o0KFT4Hrhg4nqlyR57/Yn3yOQfxBGfu
MHNVtSi57OczMfGXjqfTw0IpvycYDt93R5ME1KJyGu4c7O+SlVkNFp0Trzt0nL6hp9h7J4m4GIBI
le60nSO7kdu81D0JyzVI0fTRm+1CA79SpluJagBeGP2oL0egtLHnAV7sGitV+z8IgILPQVOepAtb
s83gnVwOM5ZgIEzaXe4q6DS66P2sq+UtbczT46XQNiqmbUvfOFtaQEZzt6Nh1MUBmM6MO++Mtz5K
/UEZ5RCg3dYexFRhNeB4nOyLDEo6XarcQ+f7WVeOwhC+qz9atmD8C+CnD4FjWHqbMTluiVhEVxo0
1wa0ik6IqU0IMB0L43ZZ89cMFTjIxCtPNKU76uQJVJV7MZCrlrJ276/RJ4rGogoDOTq957GE/X2b
/YQS7ypB6hpc24sAbX281MW/y8yL9/t33YHp6Y6AYA5PeiL7avHtW4YiHU0a+EABSwz20xg7s5UP
3dila3gV4DyLMar65mr4EyG1ECaFPYPVsY4pqv42Jgv78YDmtYYjjsowvRR+1EccnhKl3wdRbdqg
kejefUlyHLqSYuS5l4ovsNhLoeSAKicJu7cHLKOG8z+4ZtY8Or9TCaLvu4O2bIGO78Liii1gt5WI
iW5/unxzy56sF7Cg3PINYZkec7AB/gLnmSCcpXDTfgcCW8R1CY0boaukF6Jpgssq23IxXP2UZ7b4
7KbYb5pvybcH+hWR7Xvgp76FOEDeRGB3OZehUAXBevUrtnQKyAOKdqKlCLp37p64X5TmHwjsY9u7
9FP9ooCBLlwoqpnJyh5y7Z2EbITwJ5K4L6Vu4qlPffGMhQ+AN4ufJT1AfbCMoY597DhWWQ+BRGSH
QTbCYem1V2ul9ReYJAN2iETir3mjqEh4aKJN8BHF1rKEu1bJemC6FPmwU0juFlnLFcUrStS7u436
kmTA8WYoR9GjWwsNq5OX9JoYuqM0/PM8kiQ2YWIx6HmbVQ6QBjoLJHYbjdu40CM6mR6OVGx9hWd8
lBbzImvTpmcbWKAaRcxrB0Ko2mCtGJ/Hinq1FZLktSRtTdLx/5aYr/gikfON6CgxnfKuRBZe32u3
Eez6u7Z1laZkAO/zqfWz3FpjIHBZAWZKYxU4nUBhtOU4abJM9V7Ut6pDIhCPH7EsfciDvKBaqQbM
vsaoLKX4Kubb1530/R0qaGZASrMRIih9S4w3oDW4vpT2S/Aq68NsyWOk8HRCaETiyElmklhZQktF
3k+qzzfxzOwlntAUvo0GWLNO9XUhxEqF7DxFjyvgiTyJ1it88NvMaOyslU9Tj3dB/UfcPe9tSweN
ZQ/LQxMILLkLzhB5sV3PjWmGwX82oU27o3FuGBa2O7W/jUMO612UT+jvg9iGg53GJONMsRDbW16B
YpjttyzlnrVV9YM8EXQLgbwns6e18P9A02SPbr42+XyLq6ezXPqnpiqOaiY7FwbPYqsFMsz9B8Kk
39OjseCxX0vwKnhazWlIN60KgtFj4kbyV6mNHHnrrW6K8x4aBEdHXOhlWa0CYzk1hL41p6z2uZf6
5Zxmv+KLCEBpvx28LJ+u7O52CIOruiK6IcrwVFkpXeVUz7W4MB44D9hX8r5DjLifEOqxWFkaCE7f
eNjq+m2Zlnwo5USwVrcEQY/VBtqAwNDSov+5Zwr7V5X/4qA4PlHIL5VVIXtLIKR2XApQF3wQtaRN
YdQ8hGC9GBSAcB62bjqpAXytXD9lMG2cB1bCEzsu7rLa1hCTB3/B1kIxytoaewPajsIj3HSisSha
F0VyHu2ZePN+Qdzm/dlLSzLIZ9DGgAQSGJrnez4rDBG1JY5yeTAkSaOsGgYZD66v5WcJxruHsaoI
8T/G/iISfr+uxtupMe/W4kwuXH5S+PHhqu9cIWnVoRG/xqSfkTKiVCHIkhPflKQL0mGgQtliEVtw
7AgdFx8GmL3BiZCFHkfxZ0Qufr338Wa+BsZNa/EURcsO3uWPvkYS9H01zSX24M+G49PhqimrrXQe
vMKS/dgQGY8BJlefHjPLVTuihk0J6FLxriNClzbzhIxvZENRvlrjWSPoajzlJLZmGPub9pRNde2H
XOjf178YdR+qCQNCF73SBTOLLF51ObcC7NTFHnY83FxpoD4IpN3e3llI7L+Gd9QoBsnN943Dn2V0
v+7Dthz+/c7pmaNNQVCbyhNhzo1HGrrCyIaNv72HeEW8AQLTLJZDwrPNAXp5pkocCQtDNteaMgVo
J4SMMU3bVo5sP7eyldXqjEbgacDjXqQ46Xtdc/z2fASt0DeWZyEiYV/uayMpX2iw266DE1uAcH2I
atisW/u5Cke05T4VMRvid9Od2e70uyA8D1DNZuZyODkrB37b9SNxlggfns6YnYMLjUWWGP5R8nqk
gWC1q7fFqeOHdbay8UxNgGdrGKqGLHGKu/oaTlvaADAju6xSsAgB8Lfv9dErr8EWLQyrCT8KA8u7
BXrWlySrSAgNTeHL5Lre/f4RRIMywMQFUFh5OvJ9kjdQRM52UpW/p7nu5/DQtlTTemfF7+MZrxhT
3FOFp+Lcj4FwP6QMEeMcqc7WtpoOeNwNVjtt+FsojpQ9H87zwtXhZ0ulLotWOC4IRSFbsFWeh1mI
g2HFasGQxFhLan5wnKOMcP6bbA2Wd/Ow7dB2zdQDuecV/fAwaIq5EBJLoer9UNh2d5Tdz4eN8BAM
/HmH6DC8KPNY0vg+8lyEqQ4DhpcZohfo3DFIgcWvMmMD1ToSd1z6AHJoqkZVaa7YKPjAqf4iE4zT
LbT9IEfyhBVKV6XRfXiFbT+EAK0xz4gNmD7IFbekqgHVh3NwSFHXmPoVznTfYP9yv1RH4hsyD7XF
CT0RAQo7DSZGbo45f8e7s6vZ0oSii+7EHB9Pxf8iH7kJfx/y+4s8laXGbqqIU7YhFUhXOYTvpzfl
qL6MTV/sHE59SBIr0HK5PPRl+4JabnXir5oWMexOma6Ty89CNgi9e0A/hLRYtmvj5Ax83iU3l+nb
EoSS6L+Dyw6XVyRjffdGjpkhLs/4rs8ROfWYIuoxmZRPrSo+L/GrTzXIe5a75uwSiIV5BryCyywF
TS6vHn3izUJiiMCOOni4tsg2uQwqFxUMyISt5R9tPnCtZxKIZ2c3JeBRyj7Rvw/ZUOdCsUWQGFin
vmr0NXQ6DwzHITrdSj50/0yYO3mmDXH25WRnr2dkoTimQRRbNLxCplAdB4N3Au5gdItWPzbHukqj
R1PhoJ4iXPEuGFaYGunOZHIl9ns5fFyaC7ZaaRq6PhrQ1PkxLAACz7tvzxV6lZ47NOCEnPWAgZpk
C2iek+2rSV3gX6VmCErfsfgD4TQltQIyEHsdHuTb24hR0ZYd7cL4oJ7wBGNBCEQzue/wNEwXkzpF
Pq0Vo6pSnaiI5bkk+GjzBWxcpoOWIz/iooONot2rMO6nLBkZ43yJm/qQDgIlyqhhTxKmSwmOnLx9
70NL2sZ1mrBXUjpAiJgaABKPXyB1Ju5GqkIEh6JKnNwbVWw5Gk1+0DJaSzZA7b/AhpqthAUrAEnE
Rgu8VZWbQKJRdjQbKvexi/4ck1yrnZ/W7+JwY/KNg67FzwjkQPyYYP7qr1gIdnh/gpHNi7+Nvb8+
LBnNTXWpnHjOO5rCOzbUYMobW30dwswUXamCrRBNiSCNTmpx+/cD168Oko4OX0pWyok9rninEP/r
vtbCMWvhqDU55XL0xHKfn/SnfNeOrRki+DwcZzEMy66QZ+B79wlYkEl2BaQ1g7gS9FMX6G/uEPX9
QdAginBmKaL/605kY51eTBHPJVOorRvI3nPU/lS0SRKth4x1l9I/FCWcgvPwBkLcyK64yVYi+9rY
e0Ze8TBx6iVTOFnszaNuyegrB+fWpcdcmlljikJQ5yCfRZExTSwphZH4gz9KYTR8UrODeyarKjFG
cQUzneQI5In+poys83lP98/iVjXJtNyhdrHV7vjZPU0UTcsh/dIIUgUucwNpS4gZpQHXAD2zuiT6
SeIr0DwN7CwlSTFXMACm6Dut/KLexAbZoOcH+lgNNd5I71Mab6IMW43o4QzxIjvOBJb+kYQO2fcu
A/twERi1okS/6kitHdX8LbtliImhtGkY5FweR7xCX6+Kpeo4NvCsgmHLdmNhByYLzPYyXHYNwuDp
ABRzzeXuXANedF8UFz0eaZ5ip0MyKJGiuQ+82VC8jjlLWRnXf/+rCsH5uCduZZ5GE8GRpqU6zUyv
rm8sQcMDzu9A8/tR9nEBxLD373FHM5fsYeO1hXd2gJtUGHR3TlPSolmuQQAP5T8afx6Y67S6qBFV
tW3sRQXReSEzJsEnEk7Ys43NAQFwgmWsBLbKbh/HuiO4E/F2l7Qn1nVioNiESY/XcrArlCXuAMj+
0Y3YjBA+kKISvnI9lqGFTJXEyJ3RxK5/BaLQXPQH9mL3oaaMIh6aPEpUy7ffUVZG2f2Au+pXinYW
+EXgbwD6jxSeeSfhVXU+ovxaPsEeika1KNO15kFPqILvFd0wKCm3p6CcLSMBhlhHkO6e98H5xntW
UVMnyYjOQLCBNILPyEORAko9YlcFlGHNQuTKORnfBpMvwYrL4wILFnKiQtglXN0XqziOe21NZJsK
JLK4Bj5Vxz2Buq7xxqfud+GQonbxJ9YMHHuFtsMLvBWiuApEZDkEQGLcQ5LIJofgU40uIISdGm9D
BfQ/zTg650GuGDRwuUqVVRk7HWBtYu5TGr3SKymgEgly3JPnhY+GuBoUgyASSlQ4AEvLIxk9RPdr
bXyi8JQN6/ZKkO3usCysQfMnyY/XHzwHGiVG7IYP5cL3Haeq8sN/66TEACj8vphdz3U3P6T/jx7y
BV3mchWlbNlHq05mQgtnl8QJlQGY9DHLWfxL22qDeqVqxkyAjBQkthDmyzDaFtF+qFYiiBfCU89y
LnE7/Sh52ekV9rrUp0HI35SJgInM4eE857rNZWivO/3id7nhG7ji343KPxZqRHdC3h+OgE40MVB0
1gZmOnWJrDNyu5TudiPYLEARW2XXa5PQP/Xa+P/JU3X+6479H3o6GeW577BAkVxOtiY/VbPgjxcF
JEWy2h3tU5fvKVYXtJifirgORdq3y7fY4zAdlvbx7NoRxPqTqlhv6J2hmdPW16h2fHazdD0fpacs
nZmEXWoD5vISXcvTRjhCsvD3GufCFZSH3owONmZIVTtPztPOvSS5EyAac4upmhV3MMIImfyYawDf
JzpzQJzJAVUrLPTCo+Zf2uPMGZ8sULwLfjSR6m87BPDrmT1OlXd0Q2GOydzC9giRsOHB4eNEwpgn
gH1y6OF4abDfkJ9bUT7HlTBOl81S8UjKdFtQs2CIzo7sy5+Pbebe3l+Pjp/GGkxkq7WtPgAgsJoZ
u9egRYiId3isvFLwzLcHKDTGPKrUjkAWvtEGVq1q6lTfDqGqjix7iwMfT2e39JdRgjlUGPXI0s0V
Wb2nDYllzAxpWwueG0oUrlNzm0+71IP65Vd7zp0OdaiNEo/02Uj/18uixQUA8+C+VMG2QJmCKgsJ
+HIvRJktzH1/mevBWwq28q3h4Nz7gtvp/dkcGGxhjkoMib79qcP62LqjE2izCvwn0FdjI6GJMiJH
lnlI/HlDbD3WhdfbFneJt7nQ+O5jIOuXKGVrB44wxKSyFsTxveaH/VVTToTJOZH71gGNbNMbT3Ub
akIZhlMPaKdXF3jIIpqv0dN8oLxmQ4pEWsDQGi+UHMciIdikHAeC+ZHjWEgw8UG6XwH5J8gA6ZNA
3ebGU3LaGlTQLvOMpf6aNE8x+GO++WPhQRxj1a+KAC/9viCGSFNEJJiA9sy+FfnxKzPYbvOLhXVz
gEgygwcIVWuHwFX4id2wJONgwC1R3YmhzOt7ZVtOaKiF93THIwSEuNqjhbYXMaFc8uFtIiwtbX7s
karZvkK0dQxBvyO0vmGXCTUCNEoHRQJO1jJrs81hHf8ThxR0ln/YEn/gDsy/y6+fWNhl9zIAVVlt
yyu2G5IehzT+VMQ8TYuDC9CkVs6J2me/yxDttrR4Vjwif0xYY2QlO7k+CzHERjyv5y4KJZqtGXdi
RVLylogz0Of1cLNZyqw4tiXz1UN3AqpBhMPC/jnl/t/q38xjZNiObV2flK9EGn/lKCl3UaegC/Sm
daGfk1zfF4Gnlq1njjhpuIaaqafsEUzrEZsaOg1IuUoPPHEskGglhyNapdlEyytur/QgfzpJYpeX
b7CaiQY4PiXxrj4de3CKDt9JFCbgI+s6VTIpqjEE343P9yxOIZGsV9h6LYEWlpOcOuebD2kUo6eQ
9CLOSs38t1EDd0bSToy4cuBWHJh2nQbPwmZa2dLuerdhKZw4tfLqEG7tA5xRMgZDi/scDFCsFfbK
jdKYzl9lPuCIYGMNLXKFiqRN0xH7fm8Mr74JOREGxHkPm/3iwWWJ+85msz97AxRgNIDjL0826Lm/
61jUKz6ATCnz8AF+2dgI0b/SVv37zRxTGMgp7Pzws0m24YrvP1LlAqkIzEk19GluiFcQ8GTYOLcn
Lf0D64nZLDJAdwsVeaDto2FMH9JcqQPMocbOgeElPW1BtAf1kahdTpL0ofJs+rl6JnPqhE0yRCRh
wsi2dp2czKRrqLsdr4wF78H0VwignQn6b3myT0HJExVHt+4UxoaSCqBfiQIv8solMZTBbjmWBDR7
Is9ZJbzhtKxvegxXvt6sT/0RD/VClJu+dBOGjrzREymdKW5TJYrkbAAYr4ZZTk5GSbQO67oGRKkJ
gjT0HOhO+hEeFpxEgVT+oM7hIOkWBSF77AovHNlwC1kWDQMU4Q7nGiIdZDe4enlUK3WG6P3Gh18Z
S54LxhaigTYHowdY4wUNH/RZ1Tro02/DzGHCnANnVjTpKpHRKVpz0eanG6QE5L7JNkkurpW7VmRo
CClIHhxP0GwwKuEgJ8fItpV+/hcfzZ7Vlg7BXYuT4DLH//mwucUPdJRWmtS64qrHZ0xQrdTN2M6A
C8KxwAfLANpa84Yzej7Jk+A1bxcqUhBsYN2F6IavON8xgV2AWiZnTxzGnAgtwFZfPD13la8FvYx1
Tcz3WmyEVCul16Z9rMJ6y82HoTiUfAs93QBK1D0csImXKfSTK5V4U24glBfSMlF76prZp2MBOYb4
nXXWU0mdIyqd5TWXWol39VwekrAcjcyfhrN+eN3pTAIA91tNAYl82EEfmCPpvZIUh+SzDy+B+MZq
FbY65duVeehPi2ysDg0HHROJvFXNrzPETMVIAbJQsvP8PitSIv5F5xo88jSX356OrSCkN/HrUpL3
miKqNa2scIIvZlxays7SjnrSE0H/BKdOVFbNgcznuzxHwMC8am/zIDvIEIiiNuUkRFFKs5CWKu1Y
mjUTNCPCr3dONosJKfICV3tbOQbG5l9MdHoaWJGw7bkRiFmOD4DVepM5AmqJcE4wkGJNqbg7EjC5
VUXQ30KiGDLC/vp/tj9aFWQa8rdCBA9N2i7sAI32u+GK+7YOWZTkCpNBSAGW5CVlIyHLOE8V4low
8rc56lRcpF8R3OOMAZ8GHuQ65QQhuNg0py04dsiPAqTemF2jQtN5BTrB+4vPzHBYien4GWHxqVqk
59HrazxMHNdMDt9+RBqR8pPfNS0Ny+zsxMP74TPCxTesDZ/VwIKPE7XJL0svMWKG4A3gLBQymWbd
FfYx8LAOAAvUYCaqF4QrdtEp6c0dKNXz8Ds66nfUqsOQRzGV4sZcDudpB4YP23v2PJRVSbL1SoxG
eUgz6COr/dPkVSA/jBREp+mwfykcA0nZ+iZAgKWC6bqS0qlfNK4zN/e/xKHzxUvFbTJ0SLQTBtgP
cVgFeZV9yop+lgZ1GXl2PA9jjozoKEfEiGZzJJ6NjxnSqxI18OAyXegHjeLpiqb4xFGctVItFpQZ
6ttwZM/9Wq25coxMBjK29R0p5Xqc1M+l6CCMjdyO8+aCPfDEuKUC9V5UaKs6KMKH8RQ4JwCTf6WS
Z9A8fgx/+WWC/ShQymsjyR1d8sx48jP+iVFXtqdiQaC2b2XKflnllUeB9/dVTBPZb6JN+3jOYahO
cuwWAWGmqDK05U7YddvJofKG4amwT8sxITIHRPTn6oAG8zhHOi44okTORRquuNbwbtddPNtxhMth
CjX9kCqgB3vHziQcL4UMO2nVUQJGlFyvIeiFGE2BZbQgCtet4ibfoSwVbLZdX14QYA4llJqCpRzT
Aoqhz8iJFGeQl3ZxPfobQuQVUWLWb2sC48Y5c9N2Iox2bgA/Agw5jOgjgYlFjw3VtBtpBzaecweK
FS94lk6i3XT7EufcZlY2xcQqXLFtPVfa6yDide4n+6ejr6QQp3LGvZzk/gBeeqVgptyKld/n8AVH
r48+9Qiz4/GDgOnC0jplBskfeO+FH4knrt2KJYlGeGMQtsiXDNYYhSXnVMSAHJUxbJNu9htPLMoc
yTtXMJNzt/sd3CBrcWrMPo1mljz2jHtXQI4l2Pf2VSftRJM0siFCtZu5T+nAJExkDTn/XKLHv64m
yeAyH4bIVX7a9STagDGBeBALfv/6KRcWOwkxW/1enpRZOXnDiA6FRPWbGIGSha5eIMQd3orkuvkv
Ri0/069U5MSaSPbPFuAo6hKa2dF6p7yN03b74I5a61Q1yjRGUKb+GHWXXC9d+lF5O6SMQOKLWDXV
XI1bgpD9c2UtZ4+XMW11pCZiU8GAvkPH6C0o1RO2MuF+xMJN+R2s41lm2QKvbldtmc5EDNNDW8zS
6MfIbHVLX8nL5Jtul8d18y9rbZZkfGX0TtJZCXuycsCMwAdk2q+sbv2d/rsl36w+ywG076apirxl
giCY7I5NlcE705NJkelF+P7qhHRwgF0pncUOJAQhq8YusX6Cpl4fVwGJAGKwoE+VoLnVXAMweNqG
GxiBZkpa4KBJ8mcl8G/CmDBUwG8Srg6nco4iuBRTQCDY8lQiaYQGATA1NUhF2RFUsNY3YZDZAaWp
n2LfN4oC4KYpC3OzC3Oi+6fstJj6nWaJjG8KIkZYTuWWKsP6307F8I+jgtKqSWVhd/1zIgpeCoan
joBHAciUgbfkPIayGUpDyBWXe55xaCmgXcnXkjVFsm21V2PdkZfOZnjcANOK+JudMjRYxCO+EljL
ZJbrkRcRzMFHFEcyRcqf4QThm7XVSAxI231zAgyEcG9Ve01wBhnnCFShJbcpU4RiNEv0Lms7u6oO
gA/M2nG438RDeoZyhev/hW7xrLMSTyHMdft2BNZ8VNsZUSrhVHVG9/9xiZo0tDVuHZyAZBYgQagK
JY0mc7J8jDuSkVMD/S1GqVGBhtNkvR8TiPE5UTzvKi7QulGXRYoe1d6DIhFN8bzU4NCjNiIeozy8
gjVVWVHiC8mklVUVx57jNG//IuOKhoYneJUYlD2Ng/XYGosFunVThI0phE7u9AE9F5sCpptGMhQK
QPPnOxsd+U0sc1PztsOr6wYOjEqoeCXkREBjZiQPTVNS8EAteBZlQqg77i0pX9g17ZR6uN/xCvDB
K4ougYg3oIhhYF3wAKi/vVGyseVTfQdmH+7bDTvySjBcw/Emt3KQMTt/nEYKfMTfhjHS/aOSSwAa
BookbB3yvnXFGiCEL3LXKAf6R8nUtse1e+mQi5DABi+ZdFCxi/AAywgleU1Ec/sis4q4dk7oMQPW
D1ouLJUTwA8pjKyjEETBVO8whXmV3ou5jeMCGTVlNf26VY0dgXkjQfCfC/kWB05E/EKPIsX/NnO0
JKCXV7O45zUia0MiAKDLDPbfqN/WNac2g7exGTn2sU9ryrCRJzMeRsiTPZ7EgGRtg1NrTZDCk+fR
MoLpO3egHebf3frcaxX9eLAKIr/TJvZyy418V4wBocOouurlvVXDIlMKQdBvunRKLW0IP7UQX203
6p4onmYVUN+HzGnUeW0V1Cr7+iv2quFxCwg6A9JABHMBN9fnabtAQE2tGMdztMf4sFQdQ7AuVhqf
jfBN01MpDVF5SICSz/+CCvWRgDY2qeimLOdmv/n5wofy6UhKyj2ta4mVWquDp+0Qaght3Gvptbl4
rjvNtknUuyKzej9hamORMR/JA8lvmIizdWOOSd+nqRTrOlFFUF48GLP+B2o/d6YW1gQaMyxM2bRo
fsG32WTvuEht0PqBBVA2v7lX3CfkVENavtBa8HfLtMBYqWMXlHkllM/6Kv3v0jWzWIMroehZyHZ4
eJunAqGV+PwNDDJrxoHPIkyqshzZsgFPsTZ1Ah5T/53U48sn3eIZeE0IW8QSrxfJ1ASkHw3qqUI6
4P/651qjLFhSTHFvEvGRKfsH7xawoza0Tersmo/fu+244mbS2FCHiKFBowUaj6cWKQDQ+h8Fwq7Q
pDxE2o/XXATch6Qv9S4CME6F/x2OffeRMQlEE+CKHGjp8S3fclHpejKkKnNIfGWnF+RT3QSjqiv5
MU9TEPPLAJiADyOD5QpMXM87QLw/hjxyhW4tvDn/jyaAaIiju7sgvqf7VmeTaop431vrv/3WpnGk
/0kY0oACtuKWbkW/3ggYN45vXz3l0qJDMzwQCn2O1vejnF9WxJrxzDF6e4W+PaYvKp4VQ+U+QQ0N
goimoIuxUtX76eybNuNvh7sDirjRjD9VZt6qrNmDOaR9V0Czxg4JjyldK3FO/kirsLLc6HrAyL++
DEXdQvE1MttGsnnokt1z0MN08ffDN8beaWK8wCbty2jn+y5MNurYm3BMOa9YptuL16BKcyEYP7Od
AE+tc0TqmtxQoWV8TlsF/VLyaiyr6neKTxnKTL0Ewt18Vs3fU3pBS8LDeJm+OVPikIDJoe1VFqev
eUc6sifco48X/7+6knnvM9I9vdwPw7UPnntVRp5FBW4n8PNR3WCi9a0YAC6/xgeKtoh1qPVi5l+m
F7UxeUj9MsOXZ0PDuF47gn/niimtjrngLeE93OKBK3mfH5k1lsy/MSajEQEq0OT7x+QfL1QzTvlq
PM1E8573slKjVlzAkK8S+iweQwHqjQK/DWtya6V3r24mHTekVSIIcAJpmB18SRW364sMAl9sMlZ/
MBr/KZWOx3/5lRREDEsiRF6Leg6MtATyp3kIgl3wbb4kE0VEu+25pz5meCi7isgpNxqgjKP0phcr
OQrjY295ah01AoCJHXpJjgP3CnDsy2j9AT0A2hZysY31Zp5TPIyDw1RZuKIKtaBFn7gIwCcP2Lgs
yo/gfaSu27shBc4136THrczHfaSScGby2b4aRfVO8tvVetBsDGFWEsc6qJeyk6lN4EFV9PZK5+sv
0yX5g+cd4XvjpJPtQi79ApMHEK6SRpbU+QawCReO0BBaw2iu/7jQOzTHs80YHU2m27WmVlD0PnDi
omojDCTBuNnEzNpMmAWnwCH/Lio22Z5ek2MuIrJMvJGNoStLT+YQdV8oEE9kgIg/sVgqUKpZHvZQ
UyQRxZcsOizfxO6XbSu/ZJgKFdnqYjeAJPDUPGIyB04/7gtQpWbbA8fB8znCCBBILfYfr9vmzLtT
mGSEFqYM2Y0T3jWsNA+Vfc2G1Ksz5ZlNHdbY65LPqxzSrcP7Rp7pcXJs4FORj7Pz8pDD4Wm3nuqT
qOfPzh64gRJufD0Gx0lZPWWCSKmFFt5NTn/gL3xkTPYlJIe60GbmXtZVpho5VkjgZ9rRrGJKm/gC
s3VorganHHnM0OxKmGCYids8lDwxuvmRFhL9PcHkJMHGiL+NMRtwm8y+0MHSe+THYvESpIQtwlkv
JgAijyk5gZS7TsgyEFCkBBLfBEB3ROVO/RHyuDSGK4N6xMCohlHBhdIp98a4LqRgL7dwaguwTLA6
KiWGx0/31OmNb0I8O1PSxFbBMuIX1vyeb1D9Uf88Nx1oD6oUi0WvrErCMzWxpYwHxbEmsOp8oXQD
qZjq2smpyKdNPcHYdj90erv6q0eU40l3Yzz4dM7DlyeDpb6rybuNoeZWF7EYSjFb8BW2LXO3UrnB
UL+2zRXq1R9LWZ3FzST31oNg32KwqRDjX63f7uo+iJeTzn3rmPOCSkv5Oyz+ad6ANbE3AS2ut9v7
io+3oKlVolByvVFct+XjbnP+OcvMI5ovGnLoJW1TbcSnllX4nxYriGK7DGOvxSDDj8vOgArak3p/
XRDhj66Kyesc6W5f+8nlHAigTfgwaqcGsY3TpuL9OPRQePVTq66nrQU5YJXTEmTRnwlpfJzmc7bu
CT0TvkVPUiTbJzDcp/Cc7pzFa97WzUCL7h7mGYgB8J6rD4S0mupacbEh5IH//Eh9phe1/luaoLH7
7S7O6JOo9zk043XK3aM6QvTbr8lEXnyo3SqY7A6X7A0lT5z1Tm+JRqnzzLpqLf8T0huY48sz62TK
sEILAKabaWsX2o+Ynmx9BiaXVhh9VJXr5p6bHrmrdHrs5a5ve9X9H0XriD2Iv/7cA5xkX158yyp+
pqqy4uBzTAQL5sttNMAJ2YThAPHiruR3YsHyEJkv0I1DF1VD0p9n+AY59t+ZUHuIY1B+sYKBiV+f
kUVt/Uf3px4UYKsTEhnUt4TxU6oazVE1jonPER9kxr/9TUFHuVBajq6jtDImj+U9DwfstnPxNxZy
F4XSKnS7+GejYyCIEO+B7kh6nHkS8j4m6s1EojQ3+M9A8F+ARWIqhjPKq/HQmEPlcoowZ3MqRDbb
XvUkqu/BE90v6ZTWgcxUQG2mBmL6iQ1hyBwifpgfqKoi6lWMPtxgJ++fLLXKxqrzF/J6vqxsLutt
Tdjh0OBbmfpVB9wE60KD4hwuqJJGd5W1gBM7iMqjfZbDTP2YySD6BnGdof7Iz0SY+rSxiKDzrq67
vDJ4WlfSCi8gV6d5UbNyBVwCgw2XfD0q0RkzeGIPG2A7ep30x48IvVL5oPd2UfrOt2BNouG+lj94
qIQAGsDDBjr6+UTxGg5jYFZ6aH8/MYYAgCroshWQaCRrQ7Ur8PYboxntEs/fYtuFBtIoceWb5eY1
X8PUh4JLyrC12MchySGibyFIJNRXSOIwlTWFfN0Wy5cdQOw9B0fwK637MkboXIieIZz1DE8AbmOT
kwFeFKAbiTHUzJ4lTK7gqa6B8J3NhjquI8LLXcOwsIOyx/6DA5UqLPDSK+QC5dj1uzBYyFdsO5dC
HqYEM9TIJsHe8hcgoZYxa4QX6uZ6nkJHF4dnSKTfjVL9oDX8nrC4fTegLJWTjoPRkE7/3Hv94qEq
qloxdXl5+2W0Wg8TYhuvFI3vsdMusxV8ezQw3ajdRMaO6BLP5K286RlBdUu7KKGW1FKs+SHW+fdt
c36WBX7xen7igbNyPrbl5xVGSlYykReKRJ5lMXxQpSkkrwYv/lhcAAMb0JiyEMYHVgZY8BIyWqVb
vMLquUSBxqU1wu7CTMlXwcTiSJ8L73Kodx648uJshh4PSCCSc6lB7Z4NTXaEiGrB8IMXr+SjwKai
+Q1pBjO65y1Lm1tP2PXudH+Wmpm9xOv3qAWQzti7B5R2h5A+LGzGPGtQDHFOjhin47FlZsDmjC9a
vvDNKUUBuxuWgiYF4zzCVIy7WT8UaUYNdnirb9wEW1kp+vmS7rbsoUUDRvhfk3OzkTI+kpVGJLql
LJyzuJlwCxFpzuzuqkNeSk1+tSni6kdJFmjnxrEZiaQM4LiMAc4E5zMCTSaQlGScapbPmHLxuJTR
TxEyoPVgIkAeS2rqksjlSVGkfVvk2jEYr1XA60Ayf9s1ArdVhmcm4J+f1z/sl9IYOJcrbbPsftjq
GnJWBM/y+a0ppfcUt7OE+Q5CeHZ/SoUcmlgtRU36EmXGNvPbVtzCdsIaZS+CqSWDhcav+5lRQpgZ
BaF/8y2urjc5N9qyonTZIbHJ2/CJc/QFEwN+KZFACUS3xbwmWIHXdoCCbYJZO099GCvnB52FEVeS
NWtyOMfvDg8Fz839A29IKLs0TCwaKXb+DICPE13zk6FL4g/REyaWlgXMrNfL3aShvZmTChan5Xfq
lHULdCmYAEoN2jEzHb/jSYfKWnUa30VKh2Ss2/BEyWH5alh+c7zUf8DEFsHUajkoyyvlMsqQ3O7c
KMv1gvE9B37qe+Hu+rrMJxcxQXe3k4QzMOt5uiIT8E1IwqmKJR4Y0iZCfm1Gl92qwBxNoLC3Rr6Y
RFwzgsXzRsPrhLfeaQgUvn4hCADlpu8Z9arFjpcCbKHY8Ky+Ymxe2PkoGXpnggZKgCW+mIKAs25m
urL1SSmVEIHxXbIDxzquvJ7re60TyomlK+gvzJBQ3bu8/62hHieiKQCzHCuHMgSeHCtEBHMioFUA
o07OpAWxStToro1ll7IUvF+zVrEH7nwtioOXpwYL1Tqvab00SkXhz0HNWwBUjITeHEIoK62uKXCx
fMkthU8Bs9if2IWzJzy9rqX8145UpSNzxMNrAQRfI+ClKIMeB1YomP1FjDRZSPSrBgudtSaOinzo
GycQDWAWZBKYZOV113pcrTZ8fXbxUhu9u9/N7oOCpYH9TIZAQ1slWA6PUQp/TECV8NCQdtWNNV22
0uLk+wTx+CGobpZU3yojsHpeEAPvmIlPp+uuo3UW7h7zRqzk1R9+2i9FYaRwV6k3R3gHA10UF8t/
Y49l03yqrksrk0Aum+qVQDJOIgS18Q1unxJChe/sKSj93848ct+1el9QhqXuqxinfBr74OZMQYOs
IsmiyLHhrFVm3fz0yfKn+9e5jJzmfyZuXhTVwrqVdpLpWteeZbNikgavdylF2gHTwCAjhpa9JN5Q
pCjWApRmiPlFDzd+4qQ/VGg2qc6kgHMlX2qzHXXKRjtc0eePNU0ciAuHsRfV7+mS4uTd+firjAdd
HEeHw76jq098cjwCc9mYNwGmaBNZRpPVkDOb4cHyesVCIgQqCS/UDIswFEEKif6TnTQQhMnbUiR4
auZ31wJHGLs9tUmjs4Wp3q83eSp0TAxV+RaIt+gFZsVTgANUxBhhdhKsI8bav6WOF2cgnATEsHt6
ctBrsVYy8hvI2FZeMlesrf2kAMGDiBwxNKbPCGzM7z2LzCEvyFnsyNPBxEXuXkCdsU/cl5AZFbYu
jld8w5By9um813vKpNEL0yqGggViPhZAp4LdaHHNm+igqtT2fPB6zj2V3FP6/O1HIY/8fLy0SS5D
+eT7hPLrkd0nlWIcfF+6IIao3HjtmMcLs2OpEtjST5rNd5jDC6jnjdhm5RRSouzvabFHyMvvfkz4
Opk0JtLfKqgo6awkGYewZ6/BYi07Xkdc9G1zVsB32a4N6uGAQX5XKJfichxaRCOm6TnR4ant8uIs
oX3HK+oGpzRoZOQAE1tp0viksx2QCHy04Lyzh5MO3UoXVYjingxwMnyfpCP1eJhV1PL/5JUQBeqE
Lu2GKriQohe9ytpqz1OnXzy30ZA+vQahMFOHexPmsNZftPnofjloahHtNiQh/RsyfJp7fFxa18Zo
m8ZSlglgZpmAhs49GW/3Efqb9ENklau9+s2tvU6D0mW8Q9TnWiHagFA+6nnvWsaNSa1DjdT49zYY
kiRyR1HZ97poejfGfZuAhl6UgOhdCf37ns3LEIAw7H2QZKP5r2j0R0uPfbeob4TL1sb1tszI2UKX
nGphJXKceCjEGXM80VoEY37zHahv4b6aQxJNGqj19JCyMVFqBUxhSF1Lxgno5cl/5T6RvyIcfcqO
1nk2vJPcgW+71fK1xwzCo/D+GfGNZuTBZRDE8qak95D1v3x8GALIiFeIBNbOEIxqsHWvUHjL+vUy
dR/7/n0s36W4CN2qUiqcWDyhcMuj+bE5SZb3sllQCMQmy3osphQSYuYPFsYa0/XDgmhJwsLerJz2
T91RWW/v059XzuitVU0FH8YV2+s9VI4kc4p57cVSgvzr5uBZvUoLfPPbAvtkcSUhKbPtKmZg+1up
RDZy5a+zHaeA2pb3Z8cw6Q73JehgDcbuEL3rDhDpdiC+K2QVA8HRUMV+M46UWuR0tPbC/nr7JDaH
v4O38WyDDKB1FV7wWkrxd7BoJxiDrDAKiSg3gZmSeYDd1RaS2PHvT2VRDqjhKUFY8pWA5+Hm78zz
/3f00OOZdBETkex9E8YgCAHp4VuWHmtOxzVt/OI6XMVK7FunL2/mLJUUqOk+qVicM8qLDgl4uMjY
4V1YOrLjF2JUWc61GJf5ED3y2SFKroTto1K6cvwhAMzRZsU6aJ/R+Ejw/9tLRzElIixRNxCE2Y1k
XzhXmem0gOzgDBOjas1Om102AptmnlTWh0XrdsYpvHGi5sfNEaDo4FKYhYUwW2SPOa1FWF/pqZgn
Uc4mxEQbtdJV4XpJvFN4pZmO+vhm50MnwpZYGjc2axb6k9ujYT2QsZg/gqzuk2Kh4NLiswtAt1fT
4N/8xNxKFPT97P0L55qv5BA277/7p/VUxot4WmEUOKWD1hUqorMCnS0ihPTvP0qC9DRyjENJ/E+c
WTCp/yh83TzXRFkVFZU/NzFD0OQ4v57sfIG/+wLmaewg42jgTNlOJZ2q2J/gn9Yy+UUKqMd/R9j+
fVtFxKWrrCuWLL3A9rBDJyPp5ZN3tfBb6KC0/cYuZnTauBJIEr54PIFajSmv13JUxQ6FZSHbIwpz
rlgQfTxbPYRD3i1PYFGtu5N5NsZycTUHLMSKfJse3D87R7E8xOud0obFQbzFxyvwCixZQfFv5awq
zMym1lK8X1hYmwyHQmuZJAsVYC1IODPWuQn5xgK94RNSs73IW9hLYuEIMx/6Q4wSBDoj/l11IRba
LI26NSEY1Cl7RMfMwcAAFWRcc4tCb4yVdNFqbikH0Dc1sjaP7wiNVjIPNjtAnOW0N+WP2OFir+L9
s23VtDYyhrn6//uAILUkc3snqpud+6aSTY3KWXW0EtHzpUAKa/kohJETPtKaUITSxfFRJOB4xxMl
2NJojmvON2zvsFQcD4Q59HZLXSkYDDZHSkT0Zhc+QZ0XcWWHiBVn0uqMIGFQFEu7q1YbAqy4XX/h
loKk32vwPIlYEcFu8E4K/Eoa8G75+LL8eCnu61CwTGoV+4IG79ZH6G8c9gWXI1Z4lQJgw3OgqyYd
lPz/5nisZmhIesuBX71x926YXkbMU9ZdlZznQHjxrKO0z0/M8mTSikQqglOPq/mdU7tk8Ho1hM6Q
xbqMY6dQ0nse1sOAXBvMooUP5AH54+krpEOM2dKJOoMdv+ZSO6KXKKCXMrs15NBB+VYSPuhIiP42
XhX6OD3zGae3DcBCs/eZ9U0EoHY02rjsqd1acAfHTuZ2sYgb3TUlR1bV3W5RL75qGc1kabNxL4+n
y4Tq85PeKQvZLEXuIKY0gO41w4fQVr8fvVm7MiIvQYVPMFPQWqPcNn8KiiSOXut1RkqDCMImc5E7
M7ItNllCZgG+MTNABZ4+qZ9E+C3t0izeodxynnPqgXWSYvFg686XqrNDVFc/O4UBTpspwL3iD0mk
SFkTh7Ggun0LeQkPO6p0TuKKigqVX8UVRYKxEDiBDR4vncSGrXmOrBfwHzxXbsVG//NI30kQA5a8
oqvT7cH6yNndxEnLtKGbRKJXz90zmoqKUqNeQSud53JmgufLbJIL/H4A3PTQIcW4cUPTZvnyghzU
8gATXMa53+x+Z/Oc0TMk0GZedlGSlftLOqnGPURRgojoJizCy2JVH5OoYRq8od3kb+RaLRICt1SH
YZVgeM4Yvz5Ti7+VATMBnVvoi9YA2htloOoc8fshyqCDRucudO3p85P9Fd7ZwS+cIQMzeIf0sBmk
A2d7HkA/qUjDhbpzcsT/QFl9E1Eqd1cwa3EHPiCfB7VcxfgLYO/rAg8tI9M9cIpu90YOXIiHq9RW
XDrhVDpjBJra9Pjv8+k+ZW4DW4G3A+ZDQDikTPIZDfjKcOrtb9xQZLwuk/hn+1urjWkHKl4du5kU
sIMd+svFpAAHWIRTzNOYUt/gB809VCFEoQNA1Ql0POrwrZWuq2o/C2H9X33hr6vhLhD5JuB981at
MHVq36wtZ922GPGDus8xo69SRYUFBA+EGNTgqmrSrzRBF1AkAkQVWxo20H2+26kKnnAk4LmDilNd
lpaD43Fo03NqyZjEVQNkmKt40ZkP4yL8XMKaaETBKdCvtFuzDove7DwPqUQb/4CIDOv1/Juxy7ZY
CmF9wjH0jgMEU/FisKMUc4McFyCo+KBfyBailcpNlnQ+ysgYI0o883X357X6iGCNLRB6apC0TzR4
hJ+hxcYURg463vr+8y6nZZzfUuGcTJMwnrCZ/7SdWGUQW6ykpHpDcwlAp0A9UMyhe74kRvoe06ry
/+T0OXpIYThqiPfBZxBdF3lE2dbbsx0BVjBhCVWlM4dEd5ldIBIAOFFl0A+R/hRVmSlc8sx750h/
LnlYiPWg5TxrQcZMHQDEJb56xzHclFRqFH7v8MJNjb1XgUq4CODFgcFtE12r+kt4aeRgHqcqf5oT
ax3B/zLqOxg7VjZyURcoglvu9RzTUsVRCy+ITM6vPix9uaR+4HMx/hVUZm45qh6c5tSoORgNcM7D
fYCXn5Rdd5Li/vqOC3HDXfH4t4RdKnec3bidQq/SPLARjudy6QGi9GNPgs+e3bR1iMTGz9ZwfDXh
NW3MX+GbPiizyYQIfWGAP+8CvkdEfm4wgE1yVxe19XDiqoHeaco5RvxiPwDe1qOV6vhTYIZTI22s
rTFllmMnAHltZGqHrFbLrEPfLo9Kzvq5x1NNELR0pn5NYZQdqLTcHzfNjctjWGqQmGUlIztRlsk4
SR7i3GGZ10GVUiPpt6M3J6g5C/ELRm0PAbYjV8pTylt/xhppjyzaQ4yfrQnqSUbbjK+L/aR+/h90
L56mvYnumFtKaV9YWWJ5v3uW3APMC/gthXWoLVGede7TWT6gfB2Kk8I8hahdnP+e4t8wf1MgPITC
KG2NR6hHIpC+cG7eeXiyoIqxLuC5HFDDK9bUBYRYV2sddC6Saf0D2HaiVUnsxP4OMbNFRLSptBz4
myTQu4lzmimVkZGCcdnYSvLT5HdW/ii4q0L1mHDliPYeQFPkCwjc4/P8jJSidTPEiZI1mKoKIQn+
VcVKCKIIC+jvPabySHOXMwj2/kzn5EU1o4YdFENFoAwxtAdzvw2QaKv8NXJDnN27XRXLfREMwF1m
e1ICbIDGfacpPw8097ADdhfQp2ntvseiEhc4eVxjUgn1xFje7AojI3ZZGZXIwEDYluyGeKwaIafZ
Uiog0mNosdmFwCrgJX180sNV/RleFWweY4t7eertAZ9HA3YL7zQ9Zj4apBcEarLipEuvZCfFuk28
qb6GDm8qAXeYAjQVlXj7gG7uI28WQzAYrdw+1kai3bdAL3Xe+713dR46xTG2tWDefT8Xouaq3fg+
Q6vJjnGrxrfqu6oGFE9FlnwGLzCCcrfIs9wz03JKpX4se1nFz5HmeKRun/d5mmPFe5loUCJHcH7c
pUrV6dZ48jqN+MFQAgyCKQE6rC2ZQuxr42McoqbBvN7PG6eIP7vPmz2dJk8lMomVgNJFRb9lKLsh
GXFmhxyz8ukOsFL6yHiJ0piTvxfzwporRDKaNToObd8JymlPKSRO/G8LyfJJfcjXbwZcI4rlHQpA
iMsg6W329aChsWDs4Utt/IgZwAIagyUk2mxpvoxVlg3c7JgoxLcYXujvdILXUheIMwBLYPu6S8kQ
MupWDo+Fii2pLp8A8MGuTbi/8tteoHomm0jHGNWf6nw/Azw2XaAeLIdI9mftJlLuo7kEzG0c3Gis
GpCxbuxT8//wiN1xHCcKu5AdIc2ZlPH8YTkjFjnEekGodUV+PuF0Jtvv1ey5QpFKPNavQ9EtTaTe
MiK8iR6qR+NwJGNFItIdlj+Idyp1H98hVia9jjBIOSn+nfCf+rhIjMQMpQiP/jYrfG6h5qfPWIkq
uYkhAI0zsb8ZIDE3hentuujvFgvY0zWY+8YLy3OirVCkZmJabq94ttmEFbLgXcZWooT3Unke1qxt
rJG+gio+PeHklZck8EebDxVJUN5vuDSYFjBV3R5UOVzUV7MbHeQMTgM4UJZor7ooJ/5/G0wO7x4p
34WszmqlMdrlWJ6LyoGz3iinnK0/B6UvwDsyrU7S9D3tl+K5BX2TYrqnOyJ5fanDvy+PxoZhUyY1
Ftb4yHhGtNIW4WfMlJP1Sr+q++tZI8zMOxgZry3jsFvrt9DOapmK1D4PJ3bWyRZQJlGmZeU3a80z
5eGzDqq2a30+y137URG0LWrpxaJsc6f0D8YkvBS4d3Qvnq+7ZoEfJ0A1ZmvcdwYsBYfBQIZm5ZwQ
kPD+mpPhw3PxcPij7qqi4qErfIWruXQTTEOh1ZSmzaZso1Ftl5uxI4pvE5JSzY7hn+oEQ0pkobCQ
r8CiSKKqlwU1rwO0aNUHBqryei9kmbgJBU94nkuGToR4xEDSYzfxowK7ec63hBZnyeHz4EaEESRp
wFtAnV555s2R/uC/KXseSm90gwaoQdg+NvW5FZDj9UorjKnsEOmR6xQrXeNxS141sq+TuTzBLiVb
kCvdd5oU9KAPle3MggX/s6lFgmke9cF9Jtbi0ZtZqzG7484wK6bdARq+WQrTxdrNo6hqPo/b5VVL
fBOYdOHbPZxQj3Z4o6C+Rgk7cbhWrt03V9RS4BNKj/O5DVDaIJ8Hknx8CDekpl0QcyycWubSOzBF
/GgxHr7ZQ7M4SKAr/aq+zfo9dgiVva8ZA2Z+EaBEUGiet8CFJlfj2+Wy45WhNuhYGT6+82K0kTmC
FzuZjpoIdDYfIS1g+ixbGeDIUE9DORMa/E03oivEZkfOnDZIL0taJj/2mCJQ5q4QOdEO6DAPgXf6
FkxqJrw98E2XwK2s7vhIZZpzzVn4nGVMgQDwEtfgQ42whLcwoD/blxtfF5EK0LvOvfvHjWLJrDxp
BVrlGdfeE8Ab2+FYdYCBKD17htXXkPIEAm28QB0F5fjN0zEZhtsa0Dc9ZgLMSWGjmVU6l0yxwUpD
xoJpQeXyYbeUxQkmCh61UkrkgFNKRLGIpmv+zamu1Kvnjb6vlCJaanNciH/pK7Ym+4BYxg9DmOjJ
luj0/huxoOaDTyAMRx6PQf14PbmOue8o24w/ytWydaqqzpIkUHdXFaZhj9rCR0qvYXMMxlww/GqC
BOm0Eab6Q1zRYvMPif/BCz7R3jjViVtG/Tb2JUbVWnzpc/Vl4aNZXPQcs6Nby6+zmDa59SbiSU15
uTbwdVb66/v/8efpkJpgiNhhpXaZuOmtK7axSMJL3SwHdowLdXDgu1LDHfm0/Zf03YtdXSXhxS2t
XIAjrgiiGh3SNC09KcgENkoWqIpPiMDDGjycWxEguAugYx8qKgIy6yzzgoYGiKp7tvgGmiW//Oe+
BwgiuejC7N7R+ahyFRWMd3nbB8fyIirxKDaVt6zKbek30TSPDEVOtZU+RsrnzopxWuUZrlrzaLmx
8BuvZCz9+Y2O+keVWh1Hqr1gvWzjM9E10cstvPn+ccBrmS+35ATkaxeDqJXgUhNdZUBl9/QGFfSh
Z1qIaW6EDGh+KPfKnoneKhALQgnAdwwwFOYQP36CTy4Na+4EU7r4X0hF0cmIp6gNcIjvqtoF7vOe
4Waf6znv0VRzFvbAG7YaonnRpjol47EDsFkuaGl6z+QF9JoptMm28O42waa5fjTmvH1qGcvBQY/U
ULKTv99tVWNs6GB1LU3Y3M9PU7GyJlqWuCoCI+eGq18/6e2lMj5GyzdtQfNBh3xGs6hp1YWe7ZRp
JR41Pc2pBCM3kYAEDjpxNGxRF6oDmnBjFHLCNrnTbLidH4kMPM6s2zOk5COBmnJobw1QeBv9uheV
PoAqZG3tpj40AQK8zXV0nQaoaid2+lezjYTpuSiC2UYQSWE93KxdQEx80Lth/42v0a82bP7unvtq
ASc0Sjjtsjn/0iLNgAstn+tfUITGkgGyw0j3/urBHcHVIgYoa+ghMuANbZ1vt0kzA9W/L8fF2zak
YuR3QFsgrstEDBMDcfu3OJz6qjqhcgPg+bRoHHb5miD85hSuYxluB5lt8K1q2oKSQWpt8tWBOBcY
7khDTRvyO6XzgFFwgbaYGxC6/441E6PhEK8ChA0YGlVdrE51tJvzOD+VAEiO4RcUK3+LK4OrovGV
N5B+TKNk54JA5iQzNZjXEK7Y80xPxQq/Xhh7J5Y8FkopfsMDisK1XCyYaR4Vg9+6qh5toxqVVg8r
xmpa1RGoJA2N27B2AWhTtfXjrE/GzM4L6BKU0tQCnbOknpezlfkQaZL0fCBZjfWR8zEAu0dpMsqR
aHenkDDwHBRlYQardGQTA7rCYd4YuHge8BwpeGrrr9OHn/l3T/Sh5RTF8wu2E1N/IKeeunHAld/y
T1hz1Ho+xI6MOm/m8tHOQYL4i0JtEfcOyINCPb1yb5zcwuTZ1G65FgVV4SFZzfvE0SAXDuHepttf
+FAUOOI2eIYi9bkp0xOa95aVxlQOMbdALJDVqJovHko4Z3qmwV5ox8AJtEUpUwcVnBV7bAyNbwi7
ZGXcEm79+wN7CCVh2Kbsh0up6KGJncRmxH0bLcC0AVDFTqvmyuxNF5XMXlE5+8am/jXf1PE/T9Wu
2rgjiKPzd6OXjMnLePpfKPvdG/WodvT3Wnzh7JVPRfIzoMeSi3lMoG3TRCjT6sXgoHP+DQ19HroV
iuGaU0LS7io8ljfd0awIKd/2rAFIxyvz/cbfH0dStLLS/vg7E334kXvlKhcynBZx/jDabLSBUeY3
od7EY6dUlugCyi29bWcz5N10ecrYAvHm/wXZf7xCEpVkDt15aHGKBCaWHj8BIfBAwCX31qzP6dJ3
Teiqft61U7zd9WuG+ND7VYn3AmycuBXcUQGf4O39gQuvDPKmQ6o41Z+bhg+ULbO3jj5ohDqXz8mo
EXAPXPh4qEEN5dO2WaWL5J8VRIshOo+ofHbtzCCTwEA7PiF23kSmnimG3uDWyzknPdpMJq/TtgJ+
K1NfcvS+CfPDYdRxpJHPLWHW0hYk3vn/1sRNbiTCap2vN4/p1URRVBlzeWAXpuXQtxCRUNuGjeyd
tluI9ehWVyBGlJUPHHY4HzF3WScptfWHAkONB7ILqymCbYkMYYTS+uhzCJaflL2lUROMk+6M3I90
mtAUG2Sh8bYE59DJawwCmhY45FLi3qNWIa65a4eNt35lE0rozOdNt28hBWghgiMLQmqoffWyNcPZ
w9ztlOtKp9IqCBWQVVVgR9V/qOgA5cxtRAG8slliqXRQDKORrQNfeN4Ex8OJnEuo7mtLiC6CZCfq
v3/HfE0MFZ+KDn9fbNBXJPkLyxW3dHOWTH6aXdH8WaEAHL84YIT4xhKHV6inTALbRnHmlibZZczG
UzTqESYpjkj4jX0P4PkFtrXpeCzhdZcen4Vowydh0Q8UVdFqLgoqYDWHkFAqzC9PdjFTmRkRPYKc
3zopUr74Je1CzuFv9+8qopfkEps/ppFuRWGznS1ak2JVeqRo8TGH6jBghH4MrOjVg59WIhv2eeCi
eHZxl9kB+hn6HydvkXD6y8hP7aJwsUzF0TncrFSXVVPxAuMwyzRcrh2nT58dVVqJr7BIMc6drTHs
TTesAQrdSOT+CWl12+BggEMVbmqzVqNNOydiLXO5K+I9X8iRRaLCeisTZNa4osQMkw12GOtNIJAi
XwErQuEuMaflXfWnLA2LspivZD/aSdr7TQHqS/11N0k45GhxodgrMf5EpKV6XUEQjlMsIQ7MY9py
ATUCj6D9GhM2eEKo/20A9Fk4pG2j3lfmPr0BjGvu9rW1IiQrwuxb39zfFAAhPbFpG/z9RXsfLiLm
TYMRcA3Ci0rbUxqPxoTEpItHYbfQ8dl6lQ+y3gpdEbJtGxzZn6i/Bl3BRgGqEdV2dgsQY42c/X3p
gLpDQ3kWK69FnaNNpNiw5fpPXCMQMltm2DHNO+Rbf+qoqvx+QPqLtxI4RSieQ8G3TvrHqt3UWskX
BepQD8m1oibGV6welXS6wlPTEOHxSG5ru7avq5Xc6lJeAE/gdncxFeadbWGAsorWoFnjY7xz91cB
cEjSqQUc7G4eevKbW9LOWREk5xzhc1aSAh1ucnc0NqToLv4OVi8MzXq3VDyjpVdmQy6oScOQDl0v
gkr4wNmnaQtcb4dkdhktQLMvG08rZ8Ooh2w+4+HLoDAuxJt0rmdI5np4ptC6N7ipHBRehUmeqZn/
aI62L5IkDp0256JEijugBhU1W86c/WhxWiOipM+mfqa6hsAT5gM1408MtuNPIKzOlwPsK0Fkm5Zu
9dIsDNTuqUkxJ8p4yh/Kgxj/YOlt2Kar0NkaiJpWQ8ecw6vz1Tn8uhWH/u2b/k6ZkdCYo7Bg/gnA
uLRbCJOcGojp0JtEG3Yc8Kk0b1yiPDllBLx5RhfJUGljdbjfFXGbUCTQPSJ+OPKehvIHlgILp4NK
Xr2KqUCTAjZRRHtk4qUNlNyFWLVNMdxpHTfIkWEsZqKHmPyM6lKxkJ7ljFnlG1p0dUT8EDB5rLzB
gZ2vRpTXUbWkK634zECa6SzjWSNHvn9MEPifSxvB6XtnmsemCIJ+JdfpHcTBwmh9+14osLuJuB9U
0iosBcETM9D0qpLnYmRu4Xz87gf+G3MNRlQ4R4STmlU8OHSjg4U1tRbWqMtGZW8qkWrsGVb8LQPc
0GxirYCaG9lT9iod9ZzHMZt/Zpg6WzQ7L0/Wr4jOtPZEaMTnDIKqa0Oq5fZWCnGQpOeOoJoPPA21
LWxvjT1hMzhKjpkRJO5HSwePnERUT0PNxuzqq9fLfWTvP836gL3E9TM2v4MDloOj7KwFl8OkXDvB
OnUP7kDs+/TX8KZY1uykdEkFOYWeemwX17ChXCVNBHrOzctY86GPRUQq8N+Us+6V+N0LMnINyN7C
+mijEed6r9R7YKDX+ZDvXpMcWGETM2RdIIN7PNVXU+9MJbxpcY/aktmLbt0VJwjnh2fS0HwPMc1E
NPCAxfLLNySLf/o19zXvDRHSfpsQiGx5i81bwMoBw+SYHpfu6ZMGdpW1tjpJmQ6SsXc9wE1A7pcG
6CVbTiUzGEjfsmQiQsqZ7taeQiYElVnkrJhSFd7f3sy6/3pkTjJirvGhqSxolcXeZghFJ8yQIfCJ
T0SVpjcBWK1XUKUlagw0PVbVVMcUt2HDhxCqjXbUeHnq6N6z5M8+ZbYYKQ3Dhsl2ENEUq2RI4N47
bOavJVgMPQpqeW4wCieb6p/zeWw+PAW7tKbo6Nf2BOIph6Vgs4iN9JqPtviul9lIMn7c2dwOKfgZ
ikXSxYwfcrZpSTNLZf1h9Jxrj/PK+CI7ppXdGTg80eJigKjhdgA0BAGBZa7c28SdiXDOjQd0EjcB
osn8Ou99JhfSBFtxAlzK97WC1lrTbWcMjybUwQMQcI/M7Z3dNjMMT5I+bM+q3u1kEOT9957ixBVp
YVOZ2LOKx6Y+cp03WOSD+mba32oYl0c4FoWe9617A0kKVkpIYSuZ6g4gtgtil0fZ3CxAlQsgPqvb
e6AmF3GsYrHacNw60B7nu6N9jyNSN1B4IqqhG/mLsvER14/zKyq1bp1NPGeZUpx0MdiNUJ3lCVVW
BD/Xd7HYvqDJvAN+34eWb6Oa+kEsf8NBskJ4Rk3VaiQrEOGfXOKJ06cdsLTfqCMdaleyHl91w4nw
SZFjKIaWzd/lftvifWs6IirjD8fdzkZlxyOUP7W7G8eCFYo5ubt6Pb56sZzk062xgtb/WXShlEdu
a3n3jsT0NElmzJbN2Muxny9XTLDozoWbQyrD6jh/WCFzXKAe5V+c+VlpR9NKgo/jY+rngIhxeGya
UnMe7GpPb9CNyJvLvEPbyfvWVgSPZ400m/QVdjzVsSajXv0+jbXW7t7y+m48e7+WktQkEGh2oG4c
N1iW4T3MVk8rp9afrI4IizEIId4zNVaoJfPI/2smwwc3y5TsUFhkNagNZB18y3QzdV1a2I6njr3g
Nw/pw2vggupma2IWSJQKSzVxS8dPTaovFu20gbZ7AjgOaD+YsYy4HqS/NyX5Z+5N7k5WJhf/RPjg
YUwj7/j9MWiHj6MKfLCAYc6stxB1V6/Y6TVk4yxjV7WGU5tISZZ4KG4rqqTfSj1iFs11PFQ/j8TI
zM1Rg0AkYQrpOV2Hs97iJhHd0qzzeQUboArTytfSxwsghDziNQSlSzUD/kUtlb0PzsVtgY555gy9
m9UeV5oRf+hYn/ZIBIhXiiiX8Z/BZdkTMa/1bNkLjPt4p/0/Un7XGK2I/Es08srnBcrISSbbuzN/
XFW8wjpqhFlJmhh4IwsghWV7ePpGjbsNrlnUWLePnDii6eMLcgo8KajVR5zU8W2oyhn3uyDDXjfT
FeBQ31ibm/3f5j2J+6JF8lPydjtOJ06a/zSdRBe+rd4C6U6kPWZQlI5D+sdXnaK0eS8vjBoDXSo8
5fzz3jKW0yL4O9PlDwb8IJ7dKLszLZGuGCeiH66qbrxN0U0GOMJ4aMC8NpKz7k7urD7k4wwiEVaJ
KX2Ttbv3RraV6eBsrLQYxFRabBTMpBcyghK5sF/J6iLArgHYVbB0gOZ6MUogM7EDb49kl6aa5GQo
ISjBTKbLO8kV6sWCzUKAfYvCmKx30MS3NOKmqN1qnpud7T4CGpzxXfzFPfCQ7Pc5FKwDLhUFuEMi
Daq1/kNT9NtvIAMWRAtoaSWtLRb4/45fwQ/a84Cmfc1aBol2sYmqpM6EV487YSeA2ghQAMwC6S6g
YVdd/w3s/9hTDBYRpVoOcQElkRfJ4Fnvre31N8V2WCKYC//yoPViVFCl+jgrSE/z3VRFn7nRyRCs
whS/qnYFZx1lDwUfWe/Zb9TBjgCQmnJH70MhlXIvSqGkZbZ+Xr4xobOEmzxQkyiSGgCXz46m2MQq
qhJNI1gEkUo00oo503a39CxZ8SlcNGJSYAoM5vYTLB0z25KpCPAaMraz1qtH32FPQD3G+cjrJ9RH
d9gLq8UyA/q2OJqsXdBCHCEIPX+XgjBQkv2hvZiHciu6WCdPoLOAW1axFA48mMliDkYgg+BcbQAj
OkKosrPlh73rk5gK/2ag7FgBJIjGZ6nMnuyLDsGyadJ2RbPA3Fhr0Nu5ZSmRynQ4bMNMd4h7GqB6
bE14T2p/RNv3JGecwMtRz+I92KwwSUXCKMAzse7bNTtYCZ/W3umQYuWTVJV4La/YIpWdmG2xntqH
lBtNWngapnQDzbHOicVcyc4v1mfhwcuzkbJVl3NOdLj6jDnPZYarM8f1YXqea/I+C6PpJdyhvhcH
vr1+4+IkGnnPJaNnHKKY/YLhKb5nLSbgDIV/g57o0JJ+hVokvfTJM1F5jmc/tzt46+TFdVXm1XOP
ZyHkfFBlTqNEwLqQS/Wmn2nP3xPThD96kXwSWpPmiwV/nsMp2Xcj9uFH+ZquvdXhz6Kw/A7gObEv
tTy8QXXk2owi1uoTcinVZ9lnzvhuhQ34UC7DrgPYSEObLmm5BIWKuVH9Pg5EfDqZ+uxARoyIfHHz
mIzAeL5mEO7Apm6Bh9N5OTwlBVO7M7OtvsfSH92zoGt9OqqQ7E5S1WKqlHAdz9SgHAO05fCcOYLJ
WrR1zA7gi6nd5XGLDQgTB6DHPsSpN1K9plEOgLlhu61QBMhYpMRehs/isEa/RTXhY7sI/fNb+B3f
Bsd4FBAaLU0hG6sz1aLhXhi2QLdp08NCaCeiHnzLxhBVkO3PAT1xfkCf4rQHX1kwMK4btmmx8Pab
eRK1aov6yDqcbXt35A0cjouz5709pKGAlmJAzFkrHnAKRhy4CGY9HDzgIFiSnK4HcLWVtqx1/dgl
uxiEMsQPVN5Rm16ZCJf6QaBYlh+7yPtehWPDj3EVjtmjmvP/e39LuCmkcuq3RwDmqZSmhX+xGUnJ
kx3ZGwQVI3VxbL7TQsQsyvhqd/CXxol3snz8pWBxgRTh0elpxQCArmL2OQXCHBq2W+7HXs0s/ML3
6AiJf8qZtcSvp/X0QeBP5KQ8PYnMnSvqacQZNx3RvSLCKX/Z4BDovH5cUi108htYQa8qEL/+PwQZ
PI1ZqzsUp8xVwiD91u/wmm+rWZPpzkdiYLcXzWjuN6RGXW4kb3/R+erQRyWPyheTEM0KHQ72M2vh
XK0cLxg8hu2Hzhva0y4xE2aTKIV0kcfdrlYsTt4u7WMW5s7vTh+NVyFBBFCl0I69uZBHc1IrgfVJ
/FLaAsbJsSyzboyXZvjm7GE3YltieIZdyAa8JkRKUMPPcqVy1eiwC19XO+jDNNysJ9mzRnJy/kM7
4LiVCrQ9hm3OFG+c9HLgaqBofRWDz2FnaikyMVcMByEYCDaQDBwrXmt0wLDN43dsiQ3STuAIJJ5B
+aP1Jbre8uN5XuExWyDQxu+w1zeDBucLtwZaH9EyCvF5VV8qkQVDy1HnSx4e5aenZddcqG2rjxta
TjKC5cpdG5pzjh8jo74vj23Ascer1K+02iMT442WeAmLYDNTXbpENcMlDuqFhdxUindrwreFz+h7
TrHahqUVtslXEIeNQsr/JtbVQI8C77HlwokLQs08wpT2znHgEQ7stMPrugcjFIdmnfQ2sXQ4ns9/
TqNsbUWFxNBE/J2m8g/EVXwnSE0F2x+sw0dAZdRfq/6Vda5wFQyHBh6rcueXdb4eEYvGFlGufgVb
1zxev8zDUPm7g7DZzElbityIOCnCVzBSJhtC0c4vuNa9rxwIPO/WFIsLLfAYWLzbJLuHJqGXG9Lc
ETsHC3HJzI789DoQyr227XVt8eL7LxG6b9c1ZrAk6rbijJedI/nacXUP1IJJziEyE63qSnZB4Y9Z
lxCPcqhWnkIM48GfZzh8/1rj23Rl52YBKJC2anFghKbu+OHkyYvxf6BBP0CT6L803Z2gKgrekxM9
Pd0+WtRxUPfj3jZMgMiL/JMgnU34sPoyn0EIrxFb1TgsY6quBZPRikVSAeqDsaFOXbZ/Cyn77u79
cC3tdV6PuJ+pmVb8PPNRMaBlmktvqyUfJ89YM5Yv8XB+x8TqqK3c9mVCByAzdY7fvGgYfkgFPhjO
FFn6ZJBC3DX2YSGSUAWWXOL8Q06jHeke8nwMVjz8OcdPjtWJNoY9WtmFK7zMOgdw6B+d2ykNNbG3
pbZgl+9v0MMANsPntovqBngIwcSSw6830Li5/AvKfc8HUUBDJeQt/yldmmRr9fTrI6oeSENwIPun
gdSLnFHrwyopDG/kfnOvnQvm/CfK6FIT5HHlKZemcMICDgPzWGDN7yPE0C+GP4e4TAl/oxdZGlLD
/SRn7pxCBFA6hg9tJWLUu3JM5BmxqaSzRXoaaK6SDb68Hbzn0LFyW5zQ7fjfQIg2MDanXaXiK/R0
Voll5GKqDk+x+C+YhFeFWDefB1K+SE7NGavI0tF3Spt0PJTBTLre1bq4gGCnVzDZT95A9m8GaKXH
cydeGGWhH77vo8yJ4p0r3WpsmgVSYD2Jiaip5LzN+K+ZqqLpaMhB/wcKJJgHbyMpQbWKh1NKqbWx
DqVi+YwpdgI1QQJClntAqSK8C7mUWoyV5P/lvTIYkmGc0GUsso0rwHVbNe+tkMiw+eOhuio2bDsV
KJzxGCxG0Yf08+OmoZnamTULVVml+WpztHBjD55GkJwh9NKuyvUULfKiSblHzC+1M+MXZhalF7F3
TRtaGKfrNIbTfBe+dQMwhQ6UMGysT0iakqKAF90LPp0OgSdcTyo5KZX6H9U7z9SeYgdRrB20DCbm
D+ETyPHX9nQnrPDkR+LoWdUt6H5H/JXEN/INIhnpQg70IJPdRMEgLA9Mj0FUaCYhgYv9ZLl7tiTj
12U8vIpiPHLoIRVgMsafpf80rHl8GEHDLazgm0EHYCrJT1hfZ+V4535/qR6IE65RAxOksAHMPJ6Y
jtgszJcRmvQgefM2DbNtJUd8Mck5C0A/5Ev0DkAVNiwjGq8XyApj1f+IKPNpVaPMTWp4KLIwnjBl
io7eonndCt5JBp30kdp8bkuuuKR0TQ/MH4RrA0pmTF+X/l/5jNp+5L+dns5b7bAUg+EEYRQDY0aU
b4pAXHYSDN1X/rrWRYTYk/dPEb2tTH5flOXi9zHuFVpn8OlZ0Hb5q0tIVU6ECv2nEpgvtJZwX83s
6MRTG2xG2aJU/R5SaX1DP59z4SpmvBv5IhhC58LngUHWUoDNcgrlbBrnAMUQP35ea7mbg1tiStL5
Aahf9qLi4W06xsUj8gglVRtWZuhHQJ/ahSa70JOMNCrNzpg7RcMhbsKZ0ak3umwbwyxNV3/0D0e8
aqTg7/9RdYMadxiYqQvt4f/n1ASWaVk7yD/9OsBtBe5c/3HmEeOMxaUwFW1sFIu1k6uV+PJAzC7n
qMz+THXu8VV4rTTZZtTS7SzchjqBlDeCB0yWZ+bM1kPDBrdSGa06ww7bd/ctftdiKoB+5cEBD571
s5HNkKefwzC26eCLGsRtBbXb10sDWuIzgnisTRaoQShw+8VgJJCV7GVuYGft5v0TahlAFR1w3F5m
EAdUJqdJtLEE0ZWP2TlMSrSNbdeh0TS+CCuBjvljJzNAGMdurSTeUcZFk4vxNpv8G/nqKhNnzXiE
D9Homru1M5WM8SEDe+o/OaUtO1BNf5aUeQx0UKDMXiDpomP6Gc+C5JrslxLWm5iSclJE2XN7VQUt
0jMCi5ux9HT5Gb6yu3S6/5be1lmaC1tJIBmN13gww4eK+b6VjvkKQ+1DjCpRuALnjOJVx6c++QX0
NSthH4ZGO37889vUxpHhCTVLLdp0dy8sKMkAW1CzcKsQU3UY+Ann+L4qMiByBKzdKdqKk+U6JKh1
HLIgaMg1jrUpYTUn/L5/FnZAYvdeRTS11f91NHu54zwkxvSa4qu/96eUng7dlD5mWqtBtz8rqSX6
MAuu3YTeJOy/NGJjxOECxsPuUwakbZKXBNb5WHRGByCtZNUrvnlXbButLLFaH5yN82vO0eYPnx08
Vl2e+Djj5zwrl/Ep6CDueD7PK/e2FLXea6y7BcH8/8E/20r3hf1WK7bpUFW5fk/Sck2LXS/hSfEk
jnqXISYoykKcP9Exj9hlT4vuSVNVP313ZDqHravPGu3fEyxOSp6H/M3kIFQHDXFFdrmGOS2gj0e3
hFo8bCcXBiscXMhm2hU4/IquvRHdqUAg9Bx5fW0ai2CAp7Vrx6EcLunQQYgyeSP6GDrhBPW00v/9
MINZEQeUwZXKa2YI8nkZCV6I7bPU3eU7icYt1wUWLCriTvemC0qBVEY7Z7E+7Fh/4Ob2G8Vx2t3X
KpBFZYn9K6+oBiATY6kMriMZSPH+aJdNg2oWwW8rZwC1NghqRJQgo0b8yseWEhBbyIAJgCGSBQ0t
uTpRuNF5ZRw0nYFg4u5P2g0Ol3HEfYICLUXnMpBEBPXhp/i1E52l+8sq9fy+eHI5FYjmIwQAJ9Q+
0GsJKSpX3IlqaITKB78iAdATQnOhj5CxocDow5zU8xkVa96Um8eL1HlfwOL4EqipRPZFplkr5ZjY
YeFuym7eIbDIuyPzVfcTx0jSYY24576TKAsfgpLiORc63MUsmEQOZPba9DWpYR5N2OZ7aSx9RxaV
XvGXxOJkoJ6HKryxutorFuiOIglv7BgjwNstRvrEIuoy20UzpuzPzrkL9J7Gn+GCc2RLIgub76MJ
8meU4Llv3Xx+c/K0rdtoIZFTHoEfcJTlsrrG0l48NEMnqUnpZxSMierGrooWVOCfvXEsgEA5/PYk
4zwARI8kqWsG3a1uB+6XOOmzBIhYCkY5tPYYny1gFmdB3OT0ecB5h9cvF5/2wfnnx6obbwR9Qbp7
I8dhsrGKo4dwx4w2dirk6MWPKXeD+lNjsuKuGQ26zlA8/cJnoVTreTztF+rOxdssYl2ZkSm6COMX
DL1JDYvv99c+k5YrP6nJoNlu0u2lJ+X72ilMxBku0n3PzQ1ZYVSt4w+jIlIGtIQu4x3Pq0pcy3c6
3kp8uyETZNMEtD8C1bJx8aBJx6763+YceKCgzA4+QjlkCpCqRwO4XrEzMHy0xYA3+fAtWbt0QbEj
L50iW1YLadzuYrGcWWGE+JcHnp0TOJMGI9tjw2zDKnZk7tnWEQZwCwsFFr8zwKZEIuCLRMEX94cX
8fDvZiD0k+0/WghjoQTgFAfnrlNfXas5VCdiyeaXZZnp1/5X2vDblCbPqJsPasqWkCfOHgjFIDEN
6UMq7QImd5i79OHqNX0xo0LMrTt3AxZ26q1Hfu4cYDV0Gwhux1lEZsUxqPcKL21XZNit8YyH5K1H
7ex93JtYEfX5+G9MuS3HLm7QBRdpOuxbTzd9/MvKlOrqnETt1/XUVOGZkw6/rjV73Kk9LHA+S6nd
E8lywgH3rPlzE4Adk6NSokKShC/Csr4zisVbn1cmp6c2EEByYc79jZjV9spVOMKBpPv98dQIl3XU
HhqcHQGQloMmAONAc4WJ2/DhVUPesCI5bO4axvXm5q1E5fglQaYmXkPDllD3U+ENxDfTrYmPjynK
/+dFWlfmvwsVf8rl/b12PciVyVl8izCNzBpJ+58Whp0lRAmDDsUPpMu3S8iJV33dXR9YkWF7823I
6OIgRm1YAmeF4apP4vX7rGqXhKC7sb+/RMaUPoFLTJb5RHi5cVgTytp7+jsy0VyOXiDos2eOdouc
mlUpQMFiDr8R9qN3W0R5V48rIO6PD1fKULsLYy6R6TbUY0Ke3T6kB68BN8KfLuS62R6U0VBXmUSd
uMxpevYF3euVWAZlzYufhbf0Az21Ys2SqYkCKuE/5rzXLsU0gS7mPD3UhgGm6FbYlRT286OI/qR2
mAb0rFNLDghW1zD7LJDlCnjkLWL79d/DQSVV5KuZPHbM1VNs/2YrXByH6wAtKbKu3HcAe8ExF8oi
VAR2KTiF5Rqq1pS4R+JImkleRsLq252q1tjMWj0UJdUeuATAFcYkKPGZqvICEw2lre/MygaTKxNh
dEct7SuY9tqORAKoRGlURhB6wl8HWuMxxgHK/XwMhXTjbz9wP3C0x7EAgKQbhZ3qn3joL9mUHnol
ywOAbGjbL+PmJQ7NGILkVTiy4WNdPnHezNkBxNZV8yDTV6RpVTdoGFi974FDoPaG4h+jMKyQ0i2X
cercxXEP0azlCxeNcdieyKvV1W+48nRzhjyFaf4DJgnrBzieIcXcP6EOuVvvCJSU7dLIYGjftkC5
bY/FAvmb/6cyHahuNvRXKcbjgRAAjU/nqj1ecXBoHSLO9Qnc8QxmPkSZOyM6CttAuJo6L7EY7N8T
LWWiqBfa9dAItKPGFps8mwdujCo1yqcnu9w8/A84XhI54YaiRg4TVuIl8O67+hcOmuiren6/juyT
MYNpy4e1JqQoCDEP48On0HR1HkVM1JAAqx+8a3UOGWlyDfaMGGbspsbGLA8PBs7RcgZJwjlwxKrI
DVeS8sXvoYK5KswtgJQc/Llpg2P78B4L+9rlJVLf0NRXC+6rji2dREgFGsFUxVzNrdrOeU+V7uTW
pKYgOlFY/lnoztsCgQHfAzyMKJh5SvJueRI2jdbzgqJn5n4oaYGB1FL+4E/4LwJQUermfiXGTa/O
l8BwyB0a/l+eb0tZUySx0miloyu5UVFG1lSiy45Ok7t54L6YlUZchzazAANpXc3qQlha/bI8JWHr
hjuCDYVMGn9C67mE9w6Vv+kueEQY+ClBXa0axiQJkaeAEaosuTAw0uzArKxFGlZYYzuZq59eIj+t
pP/6ljy5xSmrGScfW2WLq1Ih44OiowsIlfrJRP4i+bvql9NObHdiN0JKfriwfKiVSIqLwtsCmDrg
Klh/uqTRIMOvBYximh4ztGs6eteX5GOI+KIeAhTtDIbTd4mgFzDVtRxCUX1/huGNBWVE0EDTxy/4
59oUCUwh/DqFk+zQh99qcrJLsF5jNuyttLiCD5BYVxGLHY2vRUKljVvhaiERy0vGyavTerRmPWpZ
EcuxUP09T4xB/GBei/OKBXhJVkZl8PCbsT2Ig5c+f74c67as4oaVNepn1RLxImCt6eSMGpUCd6Yv
wNPJTHXvPF1yAkxe3RRC7peHeiRpHpPK4Vlwi+I4MRayC2X3cc+/YQ6frlNqyot9BHTqJBaDOxIY
283shPuqAIK1jaA8MW9Brh+q3FyOKkGoEmu3t45o227wq//9CN6jUOxAI8459X0wkh670JvmnJsR
fTH6Vl99XsBgXOyn8vkRyGSfxtige8URe6o/uuVDBQle0wN+VUO0oM1C8PLAJI0eGEXoZxE13+GG
INw+4mdyb7HUA5S1usHuu6Y3vmHK2hWv0w2sNHCKR/AMe9PkIcBOsD6dxpGGw7+7w3Nbc//mDI0X
qh/ZWLtrwyd43D6FzKRqD5rRtvGUN6zwCbmZa4X1vCN9VwwB83ytOSte70a/j2b8aHIkz2lWNN5n
4D/UNHet71C9xRDoVk8de7tEcMgTw2ffQ52frNpMS2YfHy9d/qDfuhYBVQlnubJy+u/yU1SRfftv
GFMsqkKVaPJMz7M0h0C0w+9A7eOfa1e3pkilCNd8frzXKep8vriRpjVitwP+KSbm+nRqyjn2gTaP
w5D0OsJ23s9OOu1DAeERz5zt7sOXX+Y/GAJTHoWaaAzfwCp88a8f5CDFdxDK3JUsRp88/N5eZBUC
2PNU9yiMH8RHT2SY+19kQm+PkVZU5hFP9S2ZfzXMzYMlwhefF0bjDvF9tsBDnkG6K3fhbgvD3q4b
I4ejpEnrMsuz+qCwPhJ1DUI9ba5nrP22Lo+tnox03wUlHnAXlZuJOJZOIwyzb93y7aRI4a3K7H4d
e/BTMzv3Qkv9eZgDJ++6etSpt6jwaFzCT8KGTjoU/o4NQiPhWZ+nTxn2OsENlVC3PFr0PjryG6VO
uClo9+dW/JA7EH4W3KRKsfR22efuKEgk1r+9YOPh0xoYFs6QrlQBteSdIOoK8aJkuO2Eh1LEbne/
4XBS13YkP7F9d77PX0wsU2XlbXtm1yeNQTvHh/DnbhyslLUGF1Nc2fmvfdewWCTyO8rYCLog7jex
VT27xkYyM2agh42Wt7DeiIGnpijFnlyYeLG0veY3C7r0uqCqc/O2acMbjqm4NyAb6up2Mk9Q3ITg
PS/fci9TiWYkUUVxbFD/4IA1ehKeimug9lol1yDpYh00BpSKr+xF1oqsaE0hb6IHhFRQH4QTFPaK
Pko2TftMAcEljRFPGJ/4m08GDZwP8WSZd+Gy6MlekT2UUSGtojTYWIJKUad494sW5KesSeEaYseq
+k7M3dlWHoCDfyBFU/qrj6OiaqL7ojBm81gIx6X7E87JeGj246FOdss15COtJJAWgVVbdrOJJ+zR
LPduwWZ0ou3FVSP3P34MP51svcsqcN/TfCUsQx93jNh4KD03YTRXNf/zijxCj/sVu0dYyghOP6ri
S9+kRCYuvRL0nKGjRTnoZSwnp/efmTzS9rNgjXBAuRnysOpGtQuBPPlIU3ONXyjFKyfWvNwL1u7b
WRr64ikHawVSyrcxd9eYYWetay35lMX86wZKDk1dAs/+G8VCKMVxHKKkGyvbpcKhBqATTizdLXjB
C+INpvXvLAu8KALD3XtSsf4yP48gqOqadYcyFHivjvB47Mz2I9VGeH1PXlegoO/9jsIXZ+H/PKLd
ZqFCDFRqzexguxw3yu8MuEgaPS0TM9g6YBwXrK5o/wQh2KjXkxPGGZhF3Cc5Oj85d9hAxtA2rAjA
8ixKitW89TSAfYzEvnh9akIRCJ/VkE2dCkX5IePAGQ+EhgoULNbfo2mwFmZx89/UX2/k+sy51/mD
C75AU2SzBFbITyOlQCfJMkoTaPHoJw9F3vAcDEYMeuL1u0DpEbBVxrrUFCpuPHGARkMwqA9oxAkW
yaVeAGE4ljVaN6l7TW7paXC2MMY0526zK0+gP56lJ5fUWRcX+p5X3ep2iLUHnXx5OZKsnUk38CRs
/HsExMvy5xo5Gesr9JvW7oI1zAo3oI563PnTmJPNAt530XcpLkEm3Y8t3nPuccPZ197mGM93D93G
gDNFOhMVODfRIeLsM4Sps/0Y3D/NgUUok1vf0kR26W5YtCM+TePoIea3SmGAhk3HO3rKDqNP+QXs
wLyvCKrWU5dlwYvCuEwu71omijHg7XVxI4VpROcxgcEvP6eYpiIhYRPpsUMdSnFdoNZ/+lQHvvpT
fL67vpOGToW2V/8TeEjNLe5H1LoGWwf61lhfSoN8K6xvji9IpKTZHcIA5lesD+AOW/EMrTM6SIlv
lrhTB6SoipNvnqVR6G4fp5A/Sn8qnVLcUo9cSTrEmi1kiFDNJ/tiXOq24XVAQdZlP/Nf+cCaq00N
PuJtxVu8zfJ2qLN7dDAz/Li56PuO3taa0ORiXGygKu0of1W7oac/L5czWqpZgkg4/zvaamDyOY2x
ogsIkIAycfhy3qEUldshpatKEhdEkxODWEprj089y/GZzgKBmHBdqqZDIFDf+6MQGYxv2fs873Ua
oLO0mHRdbuvLZPPB+dtBynXqeb+KpeZoTpcYXNTZdjE4pCQnlt6+9IejkLOAKmyO7rayLeaKVG2h
Yd+N5Ri2eG0X8Zh8N4UYDOrMgOXYQNLEgcZ0N1RDsEqBbOIZQsxQK3GLEXSWbRBi5qT8qx193TR7
i6Y9LMva672mJEn2UEVkh9VyCZgjTfPVpp4/lp5jhs8inweinCi1nnt4FS6c+4bg5ZelK34VQJBN
QwoLN4cke7iN/2vTCJ2nxGiCwHF2TXI4c1p4L93LYXmU2n8gMuD9mRcKRmzWnIJaBffnO9Lc4Szc
YW4dTEMTViw3Bt74SOwm3CMdZDC8nkeKjTKWSwqh5/2L3FxkRzEZOMYimrKSsaUnUs7+nkRmGZNs
NbDZZMfb8CBm4OUWCOedCELA0xrkgsYOYWGWPN8QpdNLXEsEReUEiq5+SfksZTlIXLyMQV8Eg9u/
fLtQX76hhZvQCurEhbnOhWoeNwagzrtDs9HBMxJ7MUExoGJxVmNvM2h0VIDQgFPSJmJikjvjDti/
MBJ467RWHW6mJfxlMYPHTddxm8k3uCPhJsCRSgdjoQWZQlJ4dEKUYqVbmLP7NPl2SavDeg/j37db
9WfXEstEs6bq8vbSZKCeOCTxR65scWTafMshuiT8SCiTIhSSEgETT+gpYEgnzqkadDM7U2pihICX
LLfcs9QbdMJdEgEWZXAyTuEs+BHWJ19V4g9ZCvYz4Xe+f3OH96IE7arPhhnPUH0QxsPggAp2C5ha
OpIVQTnh/m/hRTOIdghxe/oVev1HlSoDu7aYuTaqazqnug3pQcBT0rrK5Bg6+bitt/pZ20gsTAHG
CbNrm/VZr1K8PFg5kLpmj5ioF9DURn+nvf1Ct1shpDfhLuwQo/nikHmfzKM02CkFnltWqDDm5u9N
UBvBQSsYIfhIOGB7Mik70rEMLtzEWFxZDGUWi58PmOpMgp/68abGXwMPWkCaGE/2eHnWoVwN3DJx
oKxK8HAsolPAZ3oGuWuIHQ3gmmReTf5KTtUQsp2mA8VKmBsH7j8nfL/wmdiXTH06RDJK6JmF1zZI
QT/I18W9lQHdIo6Ua5wa3rUgSf2jCguIaAHmwc6HRK/ndAr3tGslWCWa1poobyix2hHYK5wQwPH7
0+QoLIDv1hKPyWTdsDVAhV+s1rXpFbpc4ZCOBWvz1P/zuvFhvlZdbC8d1vkDtFoTL7hvzEBarvDi
vIs8tt/Rt2eBrvnTGGS3oENKydMTtoGoavQaC1Ef/7z66XncG4b9N5fLYUSlGsbawVOcEhlySZzG
CT8W/anhdtmMiVljPuMyv5pOewIoxVm9TRvnGjwYk/GKQWxe+DhzTz6x7cQHeGPSyXHMcO2PvQ8B
uVpiU9mrN5iBUFdkAGpJSXbTw+EcO33Ab74RvOA7dLY6FPnl6Tg8p2az9LBvR3vjcamVH3zzQoMv
V3oVPMdj+UpbK2Pkpp6Fizj3UVfXFPesYRduuxuh+xhOpgRDmVBuUM/R9pImjEXkk74y6jFktM4e
Xx2VHZvp+yDxF06H4vIy029at6miS721V7nFOZbVCUlF1q/Wufo71RBILuKkzzObVrrvqJ+Xp9UR
UhjqO1S9ee+BycX/ecsclhe8G09OjzOo2hfisWSAk05IdYLyH8qWv2y+vHYjLrp3DIIG6G6SRlKL
5bVCGTs5fofqkn/Eq6vSD2/LgcTjGOrZo6TfDm0m/M12pWnWCccLf8tKJ0GGF14Xwc0JJVwOtBOA
+kCuypVYId68GO/ahPVEVuKZIVuznH3VaCysAnvABf/NWDpHXnSxHbeebbwPVhd+lVOmsPlwrYeV
J/I1O5A6cbs10Bc1WuGKLaoUyved+LAxsyBSN6Ud3ZQcHuPYeffwsY0jzt1xfqyWyxy1y9bqMnxu
eEFjNGvQnWnbZ+3w5Yt82u0NKYSfjZMtMzcEnp/Gu3cmY3BJvXolXzQ5o4Opf1W8IvpJIk/MRLvm
FLZkhxlnMX9crKge3XkmhYqkmCpHOdehISB/d6DNH4FbMCFk3GgvbTKLlSIZ1IN2P646NHGJDtGM
lA0SpjK2x4qVhvBkyyB7E3a3jiRf4lxBRn1m++jdNszA9mmb4xonWw04f1ykqNeF4HHYSDIGt7tx
HM5HjJiydPo4hEswwwDVX3vVZFKtxMsplbuCZafLMSHIQYrWHkLzZEHiSx9iYfhKvKtbW316bSNh
4H5GYBqMoDohGVSF6xv86kfeMyo7GlavyWRLZEziC7czAAr/GKKhSZgWfk1kLm1uluZmDoCqug/C
fZJ1uqcu3ShXOFDhoyiWYwuE3rTVcW39/NE14k3qwWaMVzWtrnySvFSkgBnsW9MxQ+1YZcz2JLZb
b4ws2KRrc9G9I28pz791BOx7ec6n2e0hUhXi3DcKu08uMxw0fZg0KnUUFP3RYkJoqyVL4rflE15q
/021HFZIKAtdF8be6oqHNdj/JaHRDz/gml+w/Qjg+zPxrn3Lv+7nXmGeohTXZ9L9b0S8/TTMKZXk
xDdtKRnqMYIVg+9Z/m+3w/dODxicio1iLXkcAA2AROv0HLvv+SNxaxlly60oIHDp30wtvxCFSrwe
AEcSf4r1OQlBhJdcr+CRaF2GIONV7BMG70ka1CwnzKeuU1f2A1xhppOBWnYFATaStkNlKlOxZuql
Ppzs2s+auk1IQs8CoevxfwNgFyHCMLJ0nDrp1HNo5ymK+rPH13UXUVG/BtKt1nYaL3t6hACH/ZFG
MTwpZq7T8O2rKlZQeePd14kvt+wRrYc/Qx0z4UHQZi3YD3PFgwKxEabp8bI/30qX8mE3LEzCYvZI
Rf67wMom50xc9uWI/qHLTVCgufTR5KZzfR4V73CGU5tYXxF6wnfbqVR4ente28VfYywbPv9u6I+t
xntLRnOny64siSWSlyQ6bTsVMRoLNnpQuqlo2jcK+D+foqBjyOAncOIar6ndPWOBaf5RSACsR+Ms
O54y/sOwGu1kmZtyBTLgMWMg4OrtmEh538TR4lJkKUL7T6wGaUJEV0EYWDVWpglc6guH+g2rFsHF
9y8VJmV5u0z7K6ZauaS6XG5bOxQkqPmx2fntY46tF8NwAH8mvrNuHxCEt7RAUHXpACM8Xmm+G45N
pDGPb5uN7nW0buFl3qGICeweRX/B6ypz+se3p9P1Er7tVufuYqVoF8EihqKzQkaJFI4rhcTaN9rq
JY7UOrG2GmsV5S0i0srVz7ulBiufSdmC15h1KxhiCqzkRC3a0ngg4YTzJkJ5qovaEJ83XTL9ZgLR
DIqcGQnx9LUva3Rk5Kz5SqHBdhgfjdhme1609PU8Yqr8R/jOKrlYLFr/82imbmvrAO1nOZj5YaHK
/96S7qms0HqG11JuhDU16P+ccwch1vm5EvB3rqjsFM9SUQW4KPQEwd8jWd8ollkmpYf3Wx/THWcE
i8lw0BC5LUHKFiaDPwUnrmZPNEIDHMPK6SAusphCQMvw+/KiAvWgYxm0K9p05iKKjZ+cl2gGyniz
A8mgSyh3tQSEpwoiKtjAOqgtC3R/xQXuB3y9+EirsBvkE4kEDRtw4vVeqA+tp5NtIlp003N+Z/ug
QkdLMsIWjHvxo/i3nxGrYjxwDssFZeqfR7LRCusWXye8MMkRcJbCTWNQmtvdllqzyxlHX8RMbmRw
PdY0IgOPsw9MFLIM3sf230ZdFcv6Wn9yUNFWcxsV/TSUNgMk/5ljirPNi0tIB8bvoTQ0t3g0Gf55
az1sQm3VQDjwdxWNmbEuXN1bi0KE6PypK9NmD8KAavQmNmv8q21dIN/zc2tnrI3xqTnxIj0oAmNj
9KmYEIMoqKdLE4Mxjv8y8kIQh1yuZ0kcGu3Mw2a/UdhZ4i/NfLzBZWg+bC3UdjCPVo2PruP7ns/m
vNi5etQ2JUPlq+AwF5TDvAwin2D+MSP9fac5I14ddQum5B1aKLX10qwu2c4a/8za+ZFJEOSrOjBa
OIQmAtUNYt5dGm1oOi2GoBJjrDG232dGH5c7E9nA8Ut27Ov9m5zrzOis3ZfEwp2uwtzWSKWpnyEk
uS5wgiY8dOymIIFR5mVeW2b+NVK4FPE5oqko8/c0Fq8wrI0aF4n60XuxXIH2b2+wFGK0e6V8+jZW
qDwDhek9Wwh5hb2eORV+osO8ii5dX9yBuWIpUZrpsyWX6+8MBgBig5WgPXPXE3TTRUO1iBxVx4Pj
/JlUhK4PgUl3RrkUwkli9gEumQicV5w/akhRJq2OJ48Pny6Dc10OW1GNDIjqwe+cnG99srH8kH1R
h+HVysG9Fv7LfCpPMkhbraeXOG59T8TJWtk6BtCnoYyNWUKva1rtN18KJyAQ/KEBoHxDG+nO1gyp
L2oxtQYNX6wa24HDZR5k6W6qfjtixb4fISWNrSznZb8muuzWBMjFBUgp/pjBqKAiiXRpWjCPywej
gT4KqP8+27VYcipj2L5UY8c9K5XP2ePfK524SDssh7IzIgQq9TZIhF3jrrf4xvG0H9dmT3T70v8t
ppDlksCyU6UKnxSnX4dmsyHIymxREpiEQiKCy7C1kqWL0MrgJeezl89WoNdXHCfqwZO5GGA6D+Ic
bQ8fU6Y/6jpOu6hUktntNfDE9XJsEDZwjUYiSAM3rYPc2fhkxCjwec1XraSMjSM0LFM5x/SvWWKy
Sl7/+AleTDSEZ4IJQJ+xbADBlA8Nmj4MiaLTZ/JHu7ZlqVCSud4/maFlINjh4YscKmXCM2Alfpgl
sFYqbNOuPIeO7bd3kE2FhDZxJOpk1nWGxP3oaaU6WFNIAqIm9TLc/XDrRPhbyzMvhmh3xoZz+pq4
FwIQqRRnS37jTBXRNvoYmFr7Hw2DSQKOYP2I8J+VPBcK14kuoXDPq+iICyCsZutjby8i8NYOPo97
U3+bxEQo3mxXbxHO2BTcQT4c6Z+1NybTR1UkJK9/mbjiRdLsgLXoDvJVJWNbUHHDMnsgXqUEZrYx
tIjU0Gow0T2FMr1ayIXKFT7zB8gOp8AU9emY8tsIq5GJ67PpgRT2qd8YCONMY8d1b+7gmx7G6u9c
3TTDh1GohY6FblIKBg+4nTgbgAdR5AzWK8h9Vaq0ctASqo+cCDFD+n6tGsdOkdh2YfWB4pzalX2h
+0MWpm9EtsgILxN0FzD98oMWTwL6BHLqcaN53tbQNiquh4au1d/xnsNIa03akwiZNOLF5yTWMKgk
j4K6rTZMaVZwBME4+L7sZiE7hBJg+kM6IRZkbuyatKiR7EUrVv7ep6vu/vIfkwwsT+1pzJGwH31d
FHb3aZ6E29lxitXzX+Gbe5hpn6mBx9joutrRHCfMHZhAe6e9ZSpCu1QRw8YwPK9mzMBs23sVce/0
V6qTzbs5oHSKdZhMIGhf91s70iSjVImQmf977LiV2HKhDx+jjEIu2XlFgxX9kz2bbWJq/mPvLaeR
AulE6liBjUWthj9llpFf3kb6XFrQdBIc2mFuDZvfjR1SyoMgiT0ywy2+ULs54t8VdO6XVvMHeZc5
qRjMsKAcxwazLcUkTfWqPiYtt5G5huAUlrQR29G2KTxVo0NLeKkD11BPZbibl52oaIi5bbALkYs8
S1S2acGnDjD4GFS7Yzz8AicJIDpDInCapuy479JK5yTm2MLfcLbu03+2XatXkvG0D399yhr8Je29
qZSqhtrnJOt8yDbn8+eRUJcz4wh09IlrcUeUr/7sJxC9GyPz+FAx5EKCghWLoLXUoygXJoTTuTH9
/3IPkMdIj5gpiao3CVSa5m7CrOUPN4xBIQ46vgQCTFIwufEdf6u9jWWh7udxISAOOYIuULPLwlTA
4bAirXcAOl61fYAx+i+pubryYQ7JTOtjiJFZFAyiGUOP7jh33nY5hiyo50+MNN1Q+/A7JLPz5uVv
PMjZ4undbd6dip9n8cexY3SRDEBjuABmHnfju1cchNdrCidI0bIz3ZNNXHwVhMdaZYIUfDirodO7
880KtYOOwFp+AjMMtub469bbtywJRYerkSv7y17+iViWdYrL9fJXtMt7EPwbZWiRctWNcQ9DuAhZ
T++b1po7NpOQKF1H/av8POLS1LwOvzOcmKAf2zT1c1hikmu4JyUyqCQeFVocfH0kRjSEOgvxuOS6
yTLPGO4T+Z1bxHB8/5MvR0FlJvh6DuVgyRl+xTARKOa6nbgip9FZkQR+8f+SBqSgPeLXjOJd64H1
SxoqBfm7MNbetekih6fTCH1eYbC32YhEjjIDPFv7VbH8uHWEhm9Fuz/IOkWxPmZyjHgZloOYpJLP
0FNqzEDMh8lowPhcqopT/5HpNV8VYik3vr2u/Uno3raryOPMdaeTfljYWsZ6RPsoMRH9AlW/U84M
s08RqBZgHSrCqKz+QJNIlaKLZuTa62AxBR32QsEmXmbGkYkbFaiEH8LimHs+zNkjjmZdzRdhDKLQ
k9ZkGnfESTbKebPMw8EjWV0xJyHjYNV1+eO+yLL/vbiWJ5Q8sr2hS/WRIL3v6/bdbwgusns1O6M0
PkxajAAzYz2nuiYfI/M0i3E9pQ+TNEYDxIoOl8cr/e5ar1zBt2xaJrzCmTHbkASb5E8onKcBkzWs
d5nqkdU+DcKh0YkW3zW9XYFjbsIxFBrjI/nGiZ3BMcnwbQ3aFqvqqRrkrM3SDAqNvAFAcvKa8HxX
UPIFQH+P8ObM7Vn3ThszD3ZWCmNrxS7R/ugyPqhDY0rceiqFSEJKCM7qaU+99R8ouf/EFIICiEtG
BOko+8PUtQTOf14gbyIt+Yf186Ai3KJfgwiDOdw1iPl48iaUIqXUwOO1kRygFUVelB86iY9suEf7
TtS0SDtmQ7ID/qo+KqC6dbjGInf8cLk0EySwVwwslHtuRegJKjvQia7T02DYwk2OpuEjKiJ5t4pz
Yb6yGOdKZ4fqLGJspkkVYs2e9QuSzCfI8g4X5YEU5SozKb7CvMvda2N0fP4QbI8QzUpNAtQQQdpj
qfWKCWoU9dRyskotQpZLt8oCe/sDYtBSBTTPdG4sC+9Updz8cnI7vnuGKSBypIQOAq+j7De3gyfd
DOZSblvhQQIRzmk4WVA9qJE5fU6QCFq5aM6bQiIbaQaE9u5LUye8ZZ0pP0naAYOz658o4DoNZG89
iTNwb4xcbJWcec5au4t/Vh6n4m0GK+mfEUeF6tBTAOlMQH8RpF2DJyOAABUP8qDAbBNtPcMguUTH
eSxOCd7pwzB2HofHIuHnERVJkerqbPG4KBf1SvNU4/T/UUk2l+PW4G2YmwjTtEyIFkGBrfw9XmAs
SPtxd+gxXhI7dQQyrwKzzxjn1Qry3gjF4nVfig5nCCUL0qXJnQ7O8hVScN8WxEcD9ePGLqLE05JX
DvSpNSScG9QSxOlRu8JcbACcjUQd708MpOwK46gHCXrnWKbVLPnU5dfsqpY2IeGEt8FPbxKwM4rI
1RfaD1vvirZzZ3mgZfrMarPX/pt7VufGfx8Wov40WfEsXqdjeP4InKT6jAvDrxyC5gUhmvnkwC8f
28yDlLt14AJdmWRTodeVwfSIQ/gCrM3Jrx25MRGje8osq3wdsZfPsPjQWL1UsGvX4J3Gxarx6egt
Dl4OewpbclURX9Xw9QpZmFdsL1/w9+o8/o599XehRhTzpH6HgtkKW7i6bno739oscyE6uueFBeMu
tG3rx9SWrHChVAIyoIGM/Zkh6wjx5DXmaz5nYAppMmGfKxpt58TA2baQph1kaayDfKi9RISZgN6E
PJDRIRv91Ai9kS9B3P6iZc3/jSSKWuXbEaQ7HE9qvTFxRXBVuuLbNfSaq7xS7Sxcnm/2VAGMBYOP
JprKaj/YwPQ1PQSoKhVu0BbYPkWy4kBwpriqvJ2LB2qI6/iz1gqfp1wU99M1mu6XHyellwbH5KHz
l7+2PhnI9PF4kzWlySKh8zOEilYLtofmqtyl+OQmVARHdRtkbKR4TPVdZUVLlw9jkBISVcjjhPXZ
YbdyPSUudvQscM74Aa9Z44peieaXZMlRLjXznRM4MZMgPFKZZ99VDZC1HJQilP6XeH5CxF2jwSYB
7R1b77M/FVQoVeFpEXVIWFH1UErCWVPVAUgbcKcAUWk2U4EX4M6F3NWngDwkYk+SurzzcCXvnPSX
D7jWkzmAA64Ot018IepFjpsV0bJXVfKmP7tusZJz6+0BW9GquiIb8H93Gcj4M4rvYe+YwKGC5t2H
eJw+Xxu9V/xCrOvDAWudOYYqZfMaYwWhZldgC2yPbbn/qo2vzqDDpTqJ1++bl5ehqHFslO7ATieC
cVvXw8y36HPwAXuiM0RWJIVUq0fSwjAPuLrbOhL5WsM/ODvqKJRZrrDE+4X6bUfPVqKFW7YvR0iq
hpvdRZN36/ThDjsbMb2oFqvb3WFvWuCCYjYH8k8y+TzwoxlHCw45VttKug67PCkht5JL9GX45qIi
/7gk1l3gcYiqU9jUnhHGa3Vk6/olQNrd0eYa+9a0PzZ0QrORXJ/af4tVRZCFMs0mF8bIlzDNHd28
LmcMPDHop92XuD2xDNOvHeL5S5ccSREEkr3r31qwWJOm3Cl8EzRGGbam4oOLz1CuYYTf6lmylDLO
CE6lMfk2Se+OTkF0tq8LZEVUBEQw0IJPPCfz61c/3x4uqbA5OIBWRa/HQpXU/w0sjiKyTB+g92o/
+jjQrgMr7MqsFd97JU6aUVnbFJx5uOYo6weUlJLTh1sfAC/3fWHQz7zzg5hh2+vhPm0xv11M//AF
YE4skdSulGamnyIbcIfRNrT2g7z04GZgQR3AFM1rrH6xLUohijAShS6TZXpP4JXBr3nziqDSKVgz
1uJu/2mjR4Zdx4+USZXFTQxPQ+4Mwej2GqvH5Bdja08Ze43N3A/CCLvj3Qd6XFM8nVF1psfJYU8H
ASwADO9frF7SKVMtDbCbuMuh2JBnPzxRUj1vTSi6HGwWszC6DqmXPjui0kjAXqyrMZv/d3EN3VmD
tWtv4LIU1cnhYtdDLcjUPDGy4CKCDCzRq+TDbgKCkLmkYn1k93yOg1I1zVosl/Cuyn6IowHldRYd
UHgx14G5SgcCNbmMc9R3cSbGLfn0ChPINbn5axqd+T4Op3j8u5AXC9bG6e482KdvBE6Vn841e6Se
blSd9HjLlrud+t4IIZl0OkmlW4w6OG4lGh54E0UuzGW/82UwRmVMWNEJ/jyn7VVUXXmHuMCLEj31
gPI0eNB/qgTAZ5njzd9LnDwmlIT4c6tIUFKW5dm/u6yfD7iJPCodQDEzfxjgB7MQXti8/EwV6AoD
h8FBnVTGH1RhnQBR9Q3HGbNwFBUr+KT60loe1pZHsV4p6HyCN9tHlIzas2dOb4BSMLpJ6rXL+3du
ZVXgyd3bWoYvqCtBJSF5sASalrPe9T16LH4RsTJUsjyEVwQvwiR2Xql3geMkjMRAsOSDu3Pz9hPP
lp+8qU+FqwuqvcOZVI6MGXOAOoNbyePaHdqbUmK63zaXwRjawDi/IPSXuopSwC/u7wWscJJ01KA4
tdaqCkMqnCruYF91+EjZIVj5js54+JlrJhbqfda8pOaEAn1TGGTOPV06wkIC7N8hvt9baXKt+k5V
EjJdNsdJs81WsRQGicEJM5G2NTUW2/odLO+bskN9rbEEHwrPfolnu89shSBewhgbml3QdsDrnH8i
HraHk/It7R7xazFA1s2AzK38wSR025e5JpQ0WgpB+5ODY5om+EiYA7TjraqenBUeia+bSwjMloPl
7hpuHrfEh72A9gpmEgl7kB3p+zQ8KwX/L2Y+HXzn5wOznj3Of5qf8UQnsLr9dPrSexlGmzcHEYiW
Qcq2PMyqtRMbdCtbVN6Dy5UaM4TeZRNHViA7b32Q0nri15OUlbC+HOYFpM61ls8H/zXi0aH6VI1K
jtNf3A7ZIRM3J/XLuwwulNQzGBG9SZiin5jJgJwbW1BCt4LozWehmkbnWamy52v7TLqtuPDreB4L
2/3DNyjyvrpCwFX65EPYoERUl7aJkhi3TlOW/Wxd8vsDe6d498NNE1S6JqGFbFGK/ADlc8Je9evR
tIQL2k8o8dVoR+W7N6T6fKDNAdM2eTS1w1VLRJ5UWerNufYPR0RKBslXDQPGK+H2ZKPkEbnMQnEu
GE6fJXoJhyXZ8fcMFtdJBeWclJL5r/OHc4fjzxktGyKO+UcYhlu5mUlLxjLH9JGavkjOhgAAVj+V
+gxAC/CUpR8+u1yK43/8vEJjUpuSyA9fDOadI+mqRQ46alVlPtEhpSnCMBQYKEKSh55NGmSpWR8i
7rdBTjlsQUYOey9uveacyrQ4O1eN2ey+UluNukDK/UzjedhEFDH/9ez/PcZj8Loxjoh4A511ZqMn
rvVWOxCC8stnTLqdPlDzrL1UXKQ+APnPyeazpOV837Qi4wDu0H6MORaYEAwYpj1dJH7R7Qekttyx
9lnV+EVfRkojNcV549W5F9MVgabmA2Alc8wo6oMK0rF1tBl1KSZshTogmu5qqupnG+k50mlX1c72
5AVGMQbXz0m59m9+aBv2XCgEJDL12e3wng7lj7uHtiX+MXHxB55GTXW7DedL8upN2Lpvs7hcqG2t
oA9zJmspDASEGWk7zvR2rSpTkHzbFMpc6I2O2yZbiL7WdqxjFGzNoIDN2jtbcO0MYPYOEVazhZsb
lT1HVZOP+bY5Fc4ipntmVLVrnc9kUDbxxFWNqxv+p3I5ENuiLC5vpLu7OCBGPUetpJkYEFJQ2aeg
76kriYMOPSb5b7PqardnNwwP56hzFQOuGfmSSftcr9+ue5tbgWreQZkavF2URo8EZpKnPEDFe6DT
tUjfC+l0k/jGCQ5BczvitYs7EbmKnz/tnpW5X+BGJcA3UJL8hoa8aUpRtTHGaHi0FcSGzC1pwoPl
CX/WWZUbWVDdWrCha2rhFru6X3T2RqOmnQsFs4SNhsIajo5LcogWZ7JYSVmVQLDYKceL1NBmxrZt
GhUnz2Mf1QO0tx43fCEGztS80tIz4AUd+g==
`protect end_protected
