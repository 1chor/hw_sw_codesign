-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
1YlSqP0CBquQl+CTwwEZxfGuP8ua+JJlv0pVXRTyiD6VfJlqpsOyExVsH/jn+bbj
UBgBL1c7lSQ8KfEA6T7WYj08ni+4BvgxjHpt7OTfoDk43nF3KXP9wzGNBI5IXXpB
AmRQWdIFxVT7RQm9nDXIA/X1CLNT0jyUQryQC0xIgSV5kMc4sk/kaQ==
--pragma protect end_key_block
--pragma protect digest_block
98F9K0CMrx3Qn8sEMSrsYHlbrxU=
--pragma protect end_digest_block
--pragma protect data_block
6sJbP6qGdxYg+nmkT28POO9v28+lX/HM9lz/l1a8zHHGnvmarsNvpZWeBRAIOkjk
mwdbV4a1ODBw/ePFEnXYsA1L8b5tIp6er93hPttxZbAvJLkcRT2SKZ2/QFsDc6JI
xFOQS4UgCtOmHYrRhrYf/hKUys7Nz8lm5bTZh3grR6043dQjaje4515ezuKZUh/7
wsPsLA9D818pGlppYE4qCWgZLGcr6PLj7JWPT0H505toLJQml9w8qOfD3zljq3i3
fE2F6jVHqmhNmkP/HP7AQlrEChkuxfmW1RCg9dUqft1owAfZNgbOuk9/cojEbWR8
oaVFmetYBmCgI7zF2uz8SN30CpTvGW563/ox3Kzwiz0PP2R1jiNERbxPk2B1Ltr1
mwTFgZ7/7IMEJsvGtM3+224toaLVMfGupLg6pvVNTGZ1iw3WtFfp5ULbq/Kndr8r
xsSh362hHvXrlrDJ3VY2HCozEk1VaCS0GFbSxOHMSg8uaA1WeIXTKLKELhOntVin
FzmwDFTZBMxknB+opLGbdylTOptaaKUvQRzF5UGkqr1174w484kNqGmdzGNNZLnc
4VHBOFXkQ5xYlGzkue4w7y6tE9KoncA0cS4Jf4s1/hN7VLLCcZTOX9wYtHQw5NcI
oj2jIKCRfjMAS3OSoQ2+vQMw+uEAMP2hAH69qffJrp8HZvxfasl/X/1H2XplsX6b
BieCUo4l8wN4ByEpKVJjX8ZG7+yyTR0JplG9m5iL9yfmQHIpZ/DYPsJPHWnd45ii
MxkHz6+YNWpUxtQHHcZ9fj2PQ1aAPsvUSXQEwnDB6nBJQzpBG7Njv+DNq3Wy1zzU
h1ylwU19G81SV6Gc+2M70eTz6I4NeOyHhVEcpZJGdHJmFD/rkGTUtHnPlsItgn6a
+J8Zwe87jCcikTmIh+XE4EuoHhDog5eUulqFXkeVsFtmCXoV8voXRNYTwE/GGkC+
3Nz1lc2/zCaJVLSXJpnCMFqKtrnkkWeBJiVVUoEmxLLZapkgapQoRJygOAqA5IaK
C1sglbiQtx0IaT9V1id7NI7WYiVCQfxxasGpGWEE4dNys13GgRMb16rCXIvpx2WH
Ud7q+VF/andwrLIjwfwakfgiG7SfNIFalOW1eB96mohH0kKk0cwRHwmQReJEwB++
2PnQGO5blvfRraZ8gqBt39vfYwsCs0NjLlUH5ekW3sALGJ83YqCUZ7Zd0jCbi3M2
ubF6w9POH4koUhkWqzzd/Aee/Zi3AIa7lZDMqO2FZsAcJ3qbDPoss1qdDviO7fFe
2/BmknlE/fgAAX1hJ1pOY9hU9wz4NF/QNFrbcquSnvVkLcWC1YYM1Ht9YVTDt0f+
QkeI4mH1bR5nHSV4QxuCmLeqTlt6VAuEiWNq3CsDXbU3q6cwHTrY4jFQ+3KUctiy
LS7ldtgSFgwknRfp5MMByVvCxWykCXTzLbyn6hENYDZvkiQy6D9urkznt7zFrwof
Y+wz2hEj5ejtTk2YFVfCUEZJ+CynesE1j9+5iXe0gfbYgvjqaytDDaN9sSaIBYgC
I8S48eFdssFSA46N48OVDCsf3HES+XA7d8QdEASIvMg3z6CnZHrymSXOIizM85br
YhuQD8Al3N+QBsf989BaJGshBgVy5w3aILuRNgVqUyFksPZURobbp+aGtzEztlPZ
R2spKptY1+vlT2VEKzfY6pkPnMmsMFewogncVfDS/fP9YaQSsWzhsUh3Gr2HrMQv
CJO9Dx63GgVe240nHOdPkIQVjA5RRcKga1H/mwdrVi8aCjtBLLLO7C3rl3NZo/9p
JfW+raUohwQ6VHapGWUUYmd2sKP5QSm5JyYZuhW6C+RnI31aTz7MthFl53dzXOtC
Jc4XeWTCua2YjzQg++0C9E1ds6TG9T39EJwOSaK/jjsxRhyXSR69ZhZaDiXKnlrH
+XX1myuUJYDFnuO+HHzwEmB5mLJED0TvBs7dMpZBDiFztrpWAnjI86TnGITZIoeS
OkELcgpW6551V2Kf13FQYl/hXw89sDW2A0vySS6h4SnkVxd38pkoJ/XsPsaI/ojX
zG6xEo6TOgwQ2LPwz7A+V9DAPaqu4fNPTKYyLYk+/wqdEQGsdEGniz4MH5p7QFqd
f05n/XdLY/8cgPL2V97566pO6Vt9UGvtjFK7/St0awkVEoezgaWAmlnj6a9YOU+U
ZbXl0Gu/AJ3J+w7+HR2grRnTNot0REkWWaS0YwYlDt7QwxYvjHbSM+AxfMU2Wym2
BJnXkpG8gOwBkaPlyQF1PVZz5bhAb9GJDHQ8jrpmhc0ISm1Fobms0Iiz0fazN4KD
V89Uq84HPyHM8JY7cK56P+GzZE7qBSrrWvkTbyn6cX1OOhNTTEUyNlbPpF8juUfR
1/mbGU84Q+q9eZnNb5abKxYKE7j+lZwWIPe/gETBAYeIe3l9iqfeoRNc5SkXtutp
N07YxMmGCtrdHGyunV5yhlJfR0quaog2oiefbwxqEsp0J5+xJfxwqLaCMZ+a9PX9
nitLajKA7f+RqBUP8fmehi3vDIZhcDsSVk/zdkN539MBu6mVRxemZwtMNI951dhs
6woLBRxTJnASPrGTV+eX6EK3LI8wI/rkLWLW61nQG3d8Ly9Cy/kSjQqe7kqsuvwo
34LVZHkqecQ8yu9Z9++T0O+EIGgMNH46Wj7b6rSbCZ2bjLxnzx6wdBDcBqGy0t9P
LSTd9KFPvQju6qu59XqGbgm3Eo03u+XvOVzg69Sf0r3pKSSpV8S5ozexW6+EU5+5
xlNgzi/NHwAJIFZsJHKrr/m2yPhAYQwfsIotb9Tbkn8D0xrLJUwfB2+wAaQquPY1
2cI+M3eO7O7vK7HbtoLB+Pq/rImf0JZePCIJeG/Zo8PacQt+PevQ6bHiqiLSb0fo
NniYQjd1a5EVLAWM6TMiM4MI7EZhHQbB5roPfnVhKUhupN66QyATRO50xN2f+e19
fYBu+v758CuylcYMaZz66u0ngcT3oVuOyES8Jz6cCtEXfBZ0A/HQElvr3M7TKZpa
kzKxC935MBwRopW7/vjry5ohDJnuxs/8QMWBiKlT6oNAVq2IeEUIQcCGyvoE5Nhc
XTi4EDpRXAfO8jM1GlhE9guxljr8H7YorTNz8IPWWbQI8brmc88recebVMS2IjkK
MHFeq9ajc2DfqTGVxKcw+v10t/zkgX9OCyj1xjWSLuUj//g/X2DAd8xEf+hWdhWQ
TVf+6JGAAr3zYIBuhFwL+Ha7bvsD5a08U+k7sv9lEzSJED9annO8wZU2Gj/UhZ6F
0WH+Zs3WBatItnAJ+8FskA6lQzr7rdr/yJQI6jW/nmw3MHuZjIOcf8xNwRnkF487
JhGayCKZ1G7gByOfQc5V5UCO8lGC2Ne4gj+R/SvVTO+BFbxxhssjqCi368vbBn2P
01mHPGnl5v8LMez5NNWJSkv2s/4HONxGj16PIM8sMf2L3UJmZTl+EJ42eGyQ9CjO
s7QhC0LfoIQwMdA0vvxpAoCr+F/DlXYxUYB3IdVzY+FokQD1d0oqWiIGCcJfCCAu
DinS32n193PntHAepdSqDh4wsIehJ7qZ8YeW/MNQ6NlnLMgFwaMKELNRWrl1AgRJ
uq3NNNjSPnYfsmRy0S5GqcUbNRF1Tf3VEwuRsltOsiOjPlpko6I+HJuv+MR4maLb
4rGMv8OLEtrpcLPLa+B+3p73TUKSS7KsgeOFCl4D1HH7ua4xIU6cUmlZrr0itLlv
FZkK8SvNU7hpBS1mM4oW8WtjoEhbK4GADJRU50ucYZwg+f4PtlsONlPt/cUZJf/Y
3zRe4vGcUfVHtZV0toQydorE+4dBaDO+ejug5nv6u24t2bZ9JyHg7gsept+xALFT
B/ZVLvislt9FdInsm+FE9Sd8oSpUilNd8az4q9ffbC2BU+RpDcudKQTIVBaDUjwN
8OQ3UVsa3RqMDB97iEi5kIZRpz/TEMqQBwJ0kuqlvJL0WnQijTBLQsCMGnkOOw4o
8ygK1YwGz/Lzk3CSj2rv8823bPK3xsrrGrkSOw7Sz58M1BIdpYV/nK6v8K9aJgTD
8926PwCmSvcgtqS8cR1+++GmAOFqNUBecu7KCMpAvrzs9Mz+dSIuIU/NDn2fxx9A
tSW6a5p0tZYp9F/teHiImZ+vgm4wkn0y6idbmQNEL5S4giJRx4gmrMwzER4Z1dxZ
jEDDbxKRvAIF0O86C07lmV9DMZKotpJdbc613maY+/vCLpjjZ+JNlAQk7yBAwxE+
4Fg4hywGLj4z+HQSab4Svn0QNuEl3hYOrJJ1vnrlzZzbYI3zJzFJhUV3/44LbEUd
BMwperN1DqUJqhkljoB60kjV9f9aAu3ISr+lm+KeN4xPDowAk78BGpMRyurTGkRI
hV9h1U34Xz/K1lrSd9souP8iX87o7+ZJ1+LiyRH/DG+KvPhjTpOFNG81jx77ruUM
u9h3Urkdr5pDA3jMPM7mMSQ59Eq+stpf20mWpIfp3MwskNbKjiG3owm6bxw2c9SU
yzLmQ5h/0Bo4rtieXzOvdC+SaopOryQN9y3VItOGNoR+L3iLiyQeR4c1l6kIc4zm
uljYrkSvuvNwYWEKCVBwcuaVRSJLea8LI8acTJ+y3zCSRk+j50Nv8K4f9SWQc7rw
BnkIW3KAhvoEPb6OA6pMY6JauYhNDqbottAYxjcuTI14r0BSWyDhRT77SAK4LyzR
skDRIcK/ZK2jlqo6ZDKaajmXeVxe1aK+QYElYO4sWboXFlsjio9dJNJKUfl9Emv/
gdy1U6av3FTEVg5NHZIf0pc2R5HhL7ghO2MD93ZiD7hjlLg7FlDikATZ7CyZHydl
CtxYWjW6Km1KT5Js+dQjVNwcxnCodHS7rSvdlEuzBLHGhUwa75fypfm8yxP1joWV
w0OVbLoTF5wt/AuOv1xGbqQ+NedlRAHyN++wv6WwAxy7Ta+opu/Hie0epg16DM2Y
PpQ4uspFyGKrGPgXW1IisTIzOnoM2N5Qs2yscozmHKjnAlv5oTSjecpXkM4U2OoE
y6WitlTiUOoJxUfQJFXyTm/8ZcA61yh6Vfx5JXeXLds8nav7u3llB/gjTUPHLaKI
ow8b9Dz9ThaSQaUqXXpEBeLau0FKrLQTohY8QpjVtGXknjLocqpWfOqSS5MKwxwH
zEOzHpblzxL7sczQUtuzDT5h7BJkexxvmERUuSLXUmNESiInAY6qim8NMcRhGsmU
ytW0Gz3VNLRhRNhk7P3KLrJhm8muQJo0QHuxuxKumUVVlAJoTsHZEj7U7QQesOtU
Kc5sK7+eRul6Qnw4S04DJPJXFLoqHBWtFe0IkTTqkWxAkszjJD2fzEOkr4s4LTVq
nHAxXxFTpgce3j8uIb5bwfQCWbqie5WinpyD0dyL0M5q97p2Pn758MbsHt/AUNjW
d79EF7BLWv8IwNq8RGFWHodugIX4nsnD/qcbr3E+ZtmZM1nurRFq/nfvLwU4X80j
1P37/bVPmSpnKZ1aCjqcwS4yN4L0+xyz8pMBnsWgeZYDdIUdABjSj93qAbsICNmR
n43easDOcvh+iHhBqJ1aUw7BaZjqigc0BeGSjoScF15ktaY0SPpNQXGr7EtigBC2
alFUUQC31JdVZSwHbkvQYFRtvCFqdeCOMmqz72LSFF01VUCPKgYSErW3Dv4sc96w
yS2qWrB9r3PI9wPX3W+nqniB+jvg5MPSspVnKTWX+CqoZShq/qngGxOzhrRK4PTV
cUKELr2bubghlS8YLLJkVQTXl7PpXybINrYeUYZ8I7RPmeeLUGdi6ipLMVUHftAd
WrDAFwiN9pzOrxOHZLHjbsNmz/RyIGcA8LfAHjEfoxeUsPhaguwk919XWZSm17OV
9vU/aOuzd6pvyaEJ8RpaQHqZzbV4knxSYmnTxzMPOEi/ucu3gJreLasUAB6f0dKP
Or15XR7B1NvePO8vE3SFzh6X8pbbxNqhiXpapoLXgKS/zXl7lm3ZKsB4O04L3QXW
XpZd5AdEk2/cp0uYqLfHxyVZD/HU05T2NmqN7ux15mihXkv2puZK2cUIBtfrEtqu
vvXijfxvVA5LW76oHwDy3RyjgimgM2w+jZ575RGtNbCJU7jTe0VGBp3VEcE5iEOC
E70hKkm/1wWFaAI8wul/vHMxC/TpuSU1VWB9HxKJnf77QXdEvryctdpbrGQqg9K9
VGJtHLYkq7Ezs2nuyQkSP7GvAT2zSnitKBs7d5+PuBQDDpGvrmJlLkopQfo3OxWh
a54O/fkbXIsPTWDB5362hbKlWjslpCixR69f/odU8jhFULJKJUj3CFRUt1tt8jKd
vnv29SJdo2j4GlMX6Hh2jdypCFxlH2ekMMTrHWeh94YsTVecno+4ebu8oH3ST9c+
ty/EjggupaUUy13FdEr7lzM6Rb/Gc/sxAYIWmk1ArUhRdmeMSKmDu4wb8/WBAuBq
5h0Ssj6up4AdHrBMWJ8SDrwCVZHZUqdEUuCOTFAY8l582WQVUDdGyr6pjH1QryBl
bzy71Ai38KfT4a6f3un5UkKBXoQVtCfYYV2WZkCCjonR3ncsr6mzcOPTJLndQtzn
1L6QEOF97Eyx5bMjgW/bUNvJIhkIzZWC7Y0jMi62mcaw7iXi9Z4HKMiGmg4oe3z0
p+2KXmHcxeORexOuAxsIngZV0zchIyJ2AocGEJ6aUH91V9FoJh9XDxeXw3vikhAx
hZWKtEWE+CI1eBmiuBNT4S9Np2IGmUgQSImeVXF5sMPWTPGdZ1vmHYRuL6JHZPe8
n4m8Hdk/9+hLcn4qojxUsv0P7Zss7wlJ93mheRWtuyqPQXT3gEFG4G6PEkQ/p7E/
izip0KKN32kmqvFB3IsnkiCTqrfc+iKhT0lGSg9lhyHX8dk6Q9nPrlX4HDOvx9V5
lGl+E3N2V+SsKsxEy3v4zzy66t6WSM8vn23/OVRrVPuYmoDR37GAvuULUnAaQT2b
TLiX8mpvoCStZPFakgsHFods1OGGEjzxQTd380hnz1rdwl8UdH90TYolyf4NWw7K
McOoTHwm7UpKXWNZS7QBKhYT6Uzn+p3vm5vrN5A8elUkxbY6AyPvXj+3t8jA12py
KyhEDWJ56QKEviimyFb41JwvBWt4fPrC7O8pWV39JZQwrM80DTlcNNf/XhycjNLZ
CM4LJpLfJkzEv6D5bDCMB7pvqoMFD1uCrNS8Vubyt4PUg4QeBapngfj0YhlWMK0r
V6iMCTR6K+lA2l6eRaSkT5FWZmWdQri1nSep6CwFWgfSYSGVP4OXpw4/Dff/srnT
4b/IfyP1I7ImbuMMMiQIOxbRn5LzBcN1aqNQ1tJbw9x5TOyvZ0obrz4TJb2ElBCN
ZyLfoCN/XQEJjFEGEhH7HheCwXbLnL+srD/th46dVEtE4eyFLVzQYMx+HNes3XSw
7CYSS9pn9hsHUlXBMVded3wNrJXOB8KjaoQzXshUPqm1H29s60Q2BeVtGM3dEy6W
gWHQWOdkvl9Tqgz2fbh8wZzi08JGvJo2a1VQNquHWNgB8UFI2zJb3owaBLW5t+4I
FPF0CppF45pQrAc+T9aBHgccXfbjRZkFoJhZF8jiwYQtOSWniLfk4V5OswpgobkU
uCegdgnWwhR5NZFjxtuQVQow+RSe3xgagT8RdQiB4DZnKx9aScp9D/e7ubYZfXOH
8swZ4sHrh3KFV0SMK2bqOta2zw4yHjhFVpKTuIJdR+bkWS3xnN8oN8ooCCQMtq/M
GkNSOxTIK+MA34he4De+qYqjf972CR6MPfvD7QY6UZvODpRMitc2cZTV0kHuDbCy
MkHVUyz6oyOamkzniOPtZjhuwx3gTSrzHoSYnC1mT73W5Zgh+a+vigu0hbhQLAm+
Ng2A5PKAOd0bwNasxg9Q2qHyPic5NBeflaiFDcKg0SOil7UL9Zvwy99hiXWhTQ7F
zAAU0lXu6cRH0K/QoYx6NwP8Cq5Ky7X34EpUkC/0eLuJBp/0ycoDLjaiNWFkfleZ
QmeVsWb3A3a7AHWTdCxRluB3ZbdmjJsnHFzG6DXScimcCeScabRt5Z7SuBlKHZL6
FViE5Uj+MaMvxE/kSqvN6TrKj88JaqcpP+nPnyNHfoQazBreMoL86I/yvZdip19p
Y7zQGe8pXuNtFtLKaiiGWXicwOqL3TPT2ZSTZn0DLM9vrZj2fPyULXG0dS45SjFg
RyQaiLYhCVKjgoIHh7gT1IcuQ/kp8Mxa7VdCA46au0Y55vi0zBRoAJY4oWirhWzY
23p+FH0AhosSoBY/CHwkBT0jp13r+J9JOUzJ5/6C9EZuOe4OzOaw37WnouhZ9ZBf
5iO2U2iV1KY3C4HcQ4RmeGz4jSiW1n6ZzrruvBfjzvKEcqOX+Lig0LnNKuYY8leO
fiHGa2DOFpZhH2m52ic8g3DXLWDMsyYt9kAEbPyQhXiVTMpkvUpJmWKhsHmu+UmH
3YArJnzjXnWzPsB1s+W/mlfrrhEJgrwhrsWi7Kjz+6N9R71sH/ar1DnPxvX+2zUc
TbyUloXHMddpykIixVbqPmPapsRTjwqrgXUT6nUPRW0+nSaH1Yb+ZJsFxucClmC2
s8pBFFrTwrGy81lmUav00YMDgFSR+R8a2crhSMC64Y3eP2yPRy/GZDsd4pE4PfZs
jJ9T2BUfjn6y1CDbEXDrofoiXYN1jakj3atAk7y5Fumh4nCytwbKDUVG6K81sgnQ
v/5p8hROVmqw0S5iI5K5t9vrm5tStszc3ADP5tFKXFQVpWt7kEhumSmDkOUL1xC0
tcvRN1pKfiDMV2LTNGjCJ3KKRUQ3jcIm04FS7YJjTlGNVJYS43u4MJP1W+DGpmVh
AKcWKWtv3Xv16mjDZyYoiiJqfCsXhMU2pVo7ii0Q0J6CwCXrnItX2V/KVvI6MPbY
1gUb8FQJr1k9UqrtBiPwl4Lz8NSVx22EEy9heVNVKZBEG1MvN5fif7+CWdDvGN4G
h2uScqHF5uo/Qql2k9iB865hI9FcD1pdOwcHLwgUWjHkybQx+y2qcA38JsE4EQV7
ZrkM+77Bzq2ZKZ4fT4W5tb7FCzAw3/JN6RfxdDovFOHQu2+bjI3r2jO8Rq54llgW
NiUoJbvtjc11FifDYjsl0tZkv9KPixaw07hErm39OSbPlS30KBkq41ca7IDczhxe
WYw5+avspJd7fJVBvUcYou3YDhJKUwv/xs/tTeSQyO9xYhJ06dn+bLnWIrMG+KSG
BwWpxJzLUKHBCRQnn/RAY5064nJ3W5BN2DQtiNs1RVJ25YMzPK0ocetOF0fWA+su
M6mnZ6Nox0Pcf3vMse1400lfYczBgFGivJjhmXQ6EYWcpzPixptLLFIGhRJKAtTG
NVVId19keb49Yms9MR/0Z9/o+HFFBPe1srbGL5XDEoiPfHFZyV/hCxGfMGlVABoX
fPDq6sSu7S/sPVtsg5uwawDmCMxeJEQcKhSSDgJkYzN2ek7sbLZMxUWXdDrK0kIv
qOWzp3gUtMLUikf2195ciO4UfBF7A+NavIgS5Ph40Q+HdaD8p/0bpRAqhlWgHE9D
1RqvZXdgV2sX8guzZLrKy0LqZL2U5DtNNXXY8YB1+3B1aFaZW/T0kyWzs225vuMU
XN+5e2zJG5UXb+ZZAkBsnHIcAUQePuECW+Ar25hhjnC0WE44ill7Afv4c8dQD/v6
LBpKCXpAblIHSwHZYqSwO+VEadytsAeEdenOp2XTMQbhLNTImoKbFDHQg74fDWeD
luG3tyaSdBGCPvWfFzelIFekRYaL1Rr19AYivXfARGZvRdOCVP31ZH1pH/xsJAmk
qtIUJaax4HfXi4ImjX3fLkJKSOJzJcAgljE7JGzl5N0JI+9qdvl4ZRqnm4ROgtr0
m9zEF0KnSlQiO5WTE7BCJVMchQrjmbimLgAbb9P+eDu1fPlWyXWp19OHm7BLLyfl
tF+9SNwPjg6F+VS+oUtDbmdN3UKyE7GBfdXCSOrC07nGQqffjSJhlTQXrxolTUA/
dpskH4x03W9JwlymBKSFYPNYt5omUIHAfNqazj8KLP8atVjYL8v5N9/rC0MYtRPs
daqHkGBqLFkvgDD1mhB+BDm5Xr7mtJADj08iRpsdnfwGbau2OctUqaWT+Jw4eK5U
x5nKP3aOkqV5JIPRsuyPJfcdEJadyKgxq3wsU60TkQBSIAtbw3BV7dJcs2Y2MEqB
39eLfWpOngbxeD/7Z75ztjU2YcHFlsf1DxapIWfSwbMBUHSM/Qu3YTHQMDE3okyB
KwYimztTh/4hlFErHfrk6F4FJ1SsTwjg7mG54lBjP4y4jbzcF79rBHBdQW47ZaHW
bkhWym9ZLcfw4IoLU8hEjM/QldVVEm1spjkXvrfF+AX2Y00T0Rx/zawLJLea75uJ
eXSlqvTnRobm4JsV1YAo4g5ILYuO+Tu30LFmwX3UR5S3KfddLJmKRppkwiS9kt6m
VuGOcVvoTmRfilVxRKAETmbZdU0dCyso8nQDftiRJtCp7n/NWLf0DaaTl4BVhY76
r502t/Ijk4JKL4nSscsRU5wNT+QE6Z8IgN/PuB3yJzEuaeKRHw7gPd2F6XXCR9D4
NCBf5gbTBY90/zhjzPgMdNlesD9agbD6NDTMt5Z73/uDs2BqYjYJMrIX9ECSDYnd
DzZFq5NBTeadlaaVmF7TSXyPQe0Z3SRnErG7fwyy4SOPP+dBxm5ieATAJKSRJyEu
hpRys0xR8mWNgnqIWZRv1KojQnWlqxqLIHpHtKJbQODz4U+LT2dJ1mMgCwXToScT
ozzlbsAKRZ48Tr6V+ZJLf11iasyE7umCL+Vj9q7+k6MzXJFFFpxDtbhMVGqvCSnw
Eb7KHqVX4G1qqjfu7vK7OjDGxGugers4WPFDrAdLQYu0p9slp2PlfX+ubAfKZvbn
bEEhQYvr/hobW5pXh1+XpeZ/Z2C3bHcod5npXhch5PaXKpgB+fHfaDcD3nj4x/yg
Y6BCkk1HGjGV9fzuFZxeHEOWk8RPT3mbtzde5wgvwrYMyTGU/JrMGHeGE1+iM+kD
aULFPsH8N0s0dJeVr9/zYQCYvWRwcrhSxMtrRk/VTcwzwkrPnay1tSdnd3kF8aFk
+VVGivhLSMG3jmAxnFJ3mpfZ9Jk9DAa8xPJlSoQBYextbFfs46MF/ygBNwUgzAJx
AVcTD5QVZf+mHLty7ZZMLeNBVBGZBhuyAMxJig9jHypUiZw+fA1G1Lg1muhWLowm
Cn8+OnhltcSakI8iZ1VbxtDWIEN/oJqtSmNCxNrOWb+2FDaopXJp+ImAi51hwzwA
1qkwNFjNmEP0ZVVEWQW87vPZOqDRv8n0159I0UgAJo0/edW/MeT2lX4UVaIIGHWR
GZuWLEDDyNK3AWZ+f+cEuTFfLsagOAuQZsYjIfB8X8Hb8j0Cij1/XP5971E6GIVS
WIOTixVmqis3ECNRKGevoZvsRwSzB3RPfWhUGOeNrRlJ40vQ9SBQ8MMciEOriiEg
J6KHMDxlGt6scKcPXoGMpaSgee0evrdl/6hLLu3QBkJpOHs3+mhYo5i6r5HaRrG/
R68+ypbPZnhgnf4Ra83kZ5m9xWL8mF0V236YQ6EMX2bqk7dgsKE4A3Kd/hI8OZgL
hXum4mw+vNtkdxCkPO/dRrvHZUYj8hUSiXGpWr47fxbh6TJYuE6cgSOkgeJbIArS
eOkgyMrrkx0TS2/NkzZ1leFN2+O4DDTQdor272ZqSDcTHMgx0fxfGZPtIO0ZTJom
bTbDjL4kNrYYGK2oVK8o1LYiVvytXC/5u6Z9VDRqufBu3/qR2UFaDAKzzp5bHnqz
xcFLTb9XQ9NYPIa2YhsggrVv9VVHX1PW4oTs2z5LkhQNAmX3FkZiAEKGsP+REwA3
WT196TSMTBxdXN2J2ina+wWufQbC+NEJD2hf5tIVdH/krZ6KtJbw3uMY4QST5sDW
zi2aNe9oQ0vCoy+PRAKGMOd8aKpLVgXySM4tl3ahfZeg9bsn/vbslMOlALOS6M1P
gT4FizWVVLjUXGxCpYvPGFwUrd9zt9Ty6uTxVKJTo1Byh3ZZ7AMHpGjvIx/MzAvh
R3vtDgSjrEBC4LCeLn2p8RkVHPkljAEbdXVHB5fc48upBdJRIA7unCSlx15wQiYu
x4uqfkhb2KxL+plbiY2jNFywC6kccb3RDPH2jjSy+s43QUFekly1YGR9GvBMYAgA
PgH9h8PqzhEjemFU70SjqPvDI6FAt0e+JKYEfUfqvKbLBogPrCLJBkLG/e9+FY/3
7v7Ex0GWkxCDGiRnTTyAG1nE574t/RS6W3qYxZwHDGjBac9/3t+vExHzQedjNNQX
zZPi7MUgtp+RLuaXdI73tPn4CE5t9KlN5bIJCAllg/OqL4dZCyK/zVpC3NzEZzK2
MiMJXvTEs1vDWnJae9tz3l19gnOf3FXlb20ewmgo3CUs0907yUwHYP5JRL69aXN7
PckcPJRRQcqX1R1TQNSR9ydxNt+7aSbQy73SShoa1YKkgJDbf3JDL6cqptoI/+GO
3gxDfOoQ/mtFPC98z114vSlzKX04FoYrmmKXQGEZwDsPRfganwBFskMkSh2EaEQB
bnxcYRrwzAw90sQPpJGegwiWheE/kjhlVln3e0ozp3JNdQxS3XtLqV60Be4apDG5
tDbUxvtpo8a5q5d8kFCBB8yeQOYLZ4yTPsJSE3u0/Fjm58BkSPlGWuqYKtaXyTEp
gFTWsMG95zQhkqtwM5Ja2hxlCg0dEJar60BBGebZHEuIAImUSNmpWsFqp9mwpaxO
nPnR4hzZ1T4eX24enYNR9s5lHeEVwkCucbXTWStdrRvsecX42MCPUe80dA99Bwud
BZfrD1NBJcS0BWOrJiKuu90V38ZAq8ikgm7y6rswwicr90KEb2KHNxm9P9tKCVdL
HqUjrE0XBQdXb5VfCA9IdOH90nzb6jeBa80IVCIQjgC4zaiILsF8/vVFx10pxuum
ouhtQ/0bnvPfEhcqC9AMAO2YAmACNdcpEbi36bZj+8wdfM97YFgVcS7wSkXPwGvD
BH4J/ZXCITokJoHYP+MYdCPr7rrsCH8GCAEnonDd8xyo00IXJJCOI8jC9zF3AlxT
+Sdvpcx0GDl1/59V4Aqif/w0vHwrOcUrmh/O37ERSNtiXc1SExpop1zEFw8T1U2D
kgSMd5AgKSnC6Z2r+4zg0c8xp1do98+u2YRDXkFD/vsFmb+40cmjSvFKNatFMPfH
cP9VO6lhYUdDkD5UGRnEYxCNTtQce5X27QLhPRb8XqfEDFsJkZtCzrmLfeBji4ow
2OvOe1MUL5rnBDA81rIoQ3RN8T3wmPSEIYD04HdaUy9/Sz67u98onkmUx6fIhMvh
a9D7fvIb+vwAOjXD7AS7uhegHPGuXpzZAF1Hlrml8yCxlOTZMChwwyLBCUoIVD67
4MwcqBRzSJ0Gz8DB+cKnt9MDSLVbA2xdcxJXDjOid/xCFNfDgcNP7c6B5TFRbXaS
I23b+DavwPNmNSw5RNHn9fJgolpljVZ0VM3fD+5w58M3OF8O0u6MbxqEmaaiJ5gp
hVYdnWvueRHuLRuQ6ud4J1ujuAIqOLIwL0GrUIVzUJ/fYyWO9W5uAG+kLawIr2Zt
VPJH6aTx8ULt2ZBfLCQTFOKBEmvSU6yFi+NNDrGcdjkMfgfG9J+tF7ew1ZTV4KQd
Or1Z2PmBBjlOXTNZU8B1YPtSa731kZqxPS/1qV81Qz0xr++1K/jBwOP0R0IBlOjq
l2SJBsujt2/IY3kwt4jmrsGAuz+l1BFiXBlxAFbBunmOnd1MzxVuwlshUP7tWZaL
21YfJ6Edwn4rmxi+CcG/XR34Oca7GsbNd0Qoy7ETRVpESg58DMkTwe9owT8PTDPc
UyZrgj0Nrtbd/g5GO9E446h2edLeXekg0SoSIkH35ajXDZAPcorP9YBs9VWJQtf8
oRLiWv6zQEuI5Kkeu5gHRk2IvNA3B6l7pwTXl5By+4d0AhEPzCQiC6wrexu8C4bA
gJiHFSetMhuucSCvBSwCXbm6unad8tUg/V1lv03LeMbc2ACa70h29Cdw7lUGID8x
VuFvyXDoHt6yhrIMP42gRPtrn3jknIr7ANqbvExle0BXCB3xrbV1+8FkyG3EROq5
p/6NaEybHegAxnPRDIZ50IRCcwjqlExlk1eddAHcCQ7g1JwoUq3IoZvvlnlkLsZT
8Wv/M8Fg54YtyTCVILsQlnCTcbwSaWEna5s6pjWLMAHQ7nPzYWQ2lsjLjUIcSay1
6lKsWPb6BmyIwzxnC+L6/dP3QeBkSbnV/KonuK0JsdAPKGXh4+Ks6FiJC4RJyBFm
0BrXYfwnqq7ypkELQTZe7iR1rJmZu336aSQr6Jd7SOgcoCquK/Qzn3DWWf7qZ7UI
kC1ZgSVnID/MzTvylEVbaKK4NKIgSVl9PjOV7TwvNA4pYci1up+hQvyIYgTKWeyg
P+Kt3UYwDn43nOELQZ5InRLJhP3oof+Yp8ELMIffA6aMcko3U7u6onhL+8QtUEP3
cejVv2uNXJgrQOn5cyXxzND6cU4Pl1/8Z6KRvDgkBLGJR3IdpbOYFdfwXNhLuXKX
KOo/euNaZq//hvdEwuF3OU/8tPG5Qw4U46wv+zsoDeDQRZx6+WGfkBR8vONSTNrV
mn+xIgvkt/TrsHOpIkbp1ppIpEnPVTHvTEg4wN/Ufyf659rxoVleDtat7e9vnKRE
tBLqHHCN0Iusq5UJflUADJ2fmnUjo40E45ii1PZt2NkxZAV5iQmtDhbTy29Bnr9f
m1Qz/essUWBg2ZCYwh/lZvtiORFEfygcYdPR+rK0N3g7fa3FnXvx5NT2itVqglS5
Zi/jRoHOQh5Zpb5Umd+ykDmi3rXt/hNuXCa/Bn/w7A6aB2rSzozPj6h0NQCAhClI
ZvMy129TlQwtCuqa6jIRaZBluXRgKN9Iun+ZOUJhQcw4Y64MC/GxTjqGgvZvFPe9
vhWEGJTCuEUnRvCf5bEhKclzz+kggvfWk7dlUVMEIZRLzdwzbQplytyYew5bse7p
H/DG1UbW9ESWU2F079lUuZarroBAY6+MtHy4NwGxsHmQNU0lKrAoMID2yLOQBnpt
C4c3lz8M4c7b9oXBDw9+UZHMZEuRPfCyrbJtZ0Rzl+QUhasho+asBsVvJjaGgHIU
OMBWAU7tlE+HhP8Y69e43UPWHPIaFpI6fvlOWLUPP47+VSfSa+q55uxS/u3aOOJC
IZ+rUq6kCpEwR1jms2+fdXKIgcSGX2c0sEmlF0yNg06hzhzpFYSljXhBji+2p8FU
r4GjWl0LXyfEJK69kPhThesUOV9M2bFukEKjUS/xxM5v3dB6WVXtVedRao/XzLPI
wy5wZJrI5FMhjyDo5aEBPtW48HsWzkuQELa03urNguhwF3o1N6Nn0Y/grbkMv2mQ
TUP17fQ56ZzSlpH1y0wztr/kK7WWd+vVio2wd852Vqd1s3ei4zBepRtgxpJdhXf6
cEquuKlaCdYKa2JUW+7WNLIYxY0lg7eibTBLNd9UGerg5w0G6HqgGUK1AE7t3aKa
dF0zK9qgK1vGuv5Uo2FtqyBHuX2j1Vu/zWIcOnnxuUSuwKLfh42d+OUAebDyelH2
TO7nntoP3gJbrzh7z5WNt9jVGCIqKFF3WZ16KUIjFL65XCyGgUhXByVXpZA6sIku
U02ZxvhrLzzbw5sMKtsf6O9Ku1mA+1PeDBa5IFmdW+UmrNrCyE2K3a7I/Ft9o9CW
sdEnzo6oxKf6CzSlY0SlpjZFVhTe3UpufTotl9JyupU7eSIrhcf8A2VwdRNm4us2
9aGjMQZey210TrZgwwbQBYwj7vz/lQtY9FxyiLA1eNrcArCeGb4ScMEb+F7W8S9N
rqWS1T2i/fUsorES4WWxl5osdAX9X9/uk5BsfMFk2EEgNDxsa9Mn26uwhpcG9iyN
5QAyQFkClwW+KuEgiZ9Qj3awBGpf/u95NzcU+hP8IBoXcSI49eNbylWeDLS0i3s8
kwLqGTDzgL6Hd9z9HPg/7Ma1k3ER2ViWpuvQFX+bKcTkIcrJvxoOAKCy9M7e+v3F
rqhpuOnsV3GdWndOOEitULVL9aJokLG3X0RRO+0U0cNu9LJ4Zv2QiKpIAhOij29I
clxupeU3YOTPhWOysSMnhykYeQSWCO8QKOrthkmUCoJVrNI0x19oA5k45CwFBmmg
ipjuz3po0YnaY5r72b4uV5d8C1m3BfB05H+ruUR5fKk+hcovvinxs3y34pCOjf68
3Vbbvd/6DPCWdyKeCbqFfrsPvM3s8A+12/czlVwgioDFkGNpZk6k/gB2x+vqo0fS
mT3djiF9XpSGSQ5pQPETwQpRSRg7xknsF8lad8QXoM9pkzCsa3ToZSt0euzC51gM
6HtNZ3vq5RxIn9FOMMFQmZ4B4rEIyoAOwS4NXDNWf1rQQmNO8ImszRQXAuuKG+z6
8dmLc64I3Er5HhRNU8WFYD9PPSIZTDqrttWN/owaVKQitm0zoHY174rhx875N81j
r7kQNE+K4Ilrsln4Xzf+YL6TfLX0gqNMA6U+icymmJwJ2rm7d+f+NXxqiPriQqaf
8UeuCAcnkq5rUo6UOs3AnojF+RBwrt+aAxG7Bsoy0+iQpEQAsTKnHiiai9RkKUQ1
KoJmKHfj3UVZ1JdCB+yODthvIvNHGeHeV1R/HxZMmXop5tu3qS84/BGu2ntchvVt
RiAZif3zNJm/HzXhbPzQos9UrL8ZM6TJe5dlfpXnQBMhTmHbXH+4BKjikc98fPuG
3JPLa71/O7iJg+EKQlTluy9zAt2MVSpfJWUB38hsymgtgfOBnm3O6L2Bg4O9xFgD
JVQ64D3SgoO8CzFUpCEHrJLtIw2sRL+qwNKT+36wMeyD8ZD1UYvYGjzfwkYa4OUB
2HrjKlyCYHdFQp2/GbyB7MvgIv9kpUYaauYA0CNQoI2uZ1xamlfCFFr2ua6QqFlX
5JW4fxVGCy5i3ksHk0SPWtBc3oWLNwQCQNIe+Jozwd6jJJf4DQzZFdwpj0FZ6Thh
Q89Nu3H8f2J0wwyOUEelR/QojlvFhcntqvytp4VSzDEjV+nryA66PA9O25+uvrEF
GZkftBL+OLiJccM2Jtz3q/TTJ3Wdabf88rsNBxTKPDb1XOmV/5bsxp5S9Cc1sdaf
9ISjuHQS2c4S/c+hqb0I7ltdlc0s3dmUEMKSID3S3j0CnQ95MTGdbhu1jthUMZY4
s15vBjgItjwkrHvWrRIdZYL6xkgOrU8848KV6IDcyC9uSOsfWcit05PksXZGYFUQ
MP27NxVS04Xmfy8tcIrJ7OEE4qe61yBXM5bPl9hixJ61tlIiJJUi+wAkZ1GI8H/H
gbGqCVr3eyUxqF66qN3yq93XCqNK3f0Rzzm/jlmr3/T6fM/TwclajaesvfiHnXud
SujTCE6dvhxAHa41Y2wKhRsxFsjP1XYfeRty4IVIcJz/xhRBt/lQa1+us5Bs9/b8
N5D4VEqCDDqPKh3ZwJovuzCWnGsSjoOooKckN6IensMya0nylsSnyiJ5PsMMw4fx
uIy9z79L/SSbVBrkrG8hI5JiohmEWV77WOruFmdRq64TFcHmW+bYcrZx+/PArukL
sukOOBHAV9P3ernr/Lvb6ES/W1IssfFwAIKc8JsKR5glDmDLq/oZa4ckH+5Bwr86
xjlKGulYtgjs8UnVpcOrjGN/wMjh9OvxcXDwadp4gil67cgUDwoJHSm11LV3GLG9
yotF9wk84luYeVgQhChEWIJ9PfSIG1g9q7SOdQGZm1/IUj9d71CuC/B1b/tTKt6G
mOr3H7VFQ0ZUNjR3RkOAyYdtoVVHb8BFoJA3hm4o2vIRLJtfbGJgCkgFNJPWK3de
IIZR6oDw3BgRhNtHyLs0ZcoV+UAyhun/52VBoOM4YUk8wN7sVOS5rLmI3e2PEaMk
m3jdgXp0gl434cUXF25COhdxSFvbUmmFAQzQ5euDk/UssJFsp8zlRF2MEnysyXUz
AxOiun3IJBftsOzPJvoRYz/75OFH20bEXbQ3Z7muzFQhA5p51yj/8Dz0Dr2MNC2R
+MGXnYLZMifZio3woTPbHEjnGXFXmDhMGgig8nEavFi58gQvC8DLvRLhIMb9gg7h
Fu2dJVgHYvNhRHKhuoJi8nCHtb8aP8P0xZlBAmIfzChYwjY/uPbc7paP/ZUmJJkK
P5sMi75kkn90pC8sOdBQxSchGD3Dbs+eREVJqqQY+ZFAJUMZf3xcnF17KdPRz67d
s9Bj7NjNvn9ROcohFcX1x9kbWvkYGtf4CFLkaCuE0xHmSwDN0XPelyYPL5M171Av
mtJ23VClWHtm5U5sKfrayvhpA2668BfCVh5SNAvmtYc4wxQiv9Twk80Ck/FNyfYk
I8q76i5VpNgWtSLk3VkXkraU+7Ku2PeYxn/+QE+qlIGMbCx8wRpnclJfR0QUzA1u
ww7SPj6wZE0VPXI4SMd6rZN/kwQTS0xJgMGqVypUhtP7hTdPd6U5ihcL/fYiG5K9
I+dAXGG0etpPMrcjuQ+t5v1SD1hKiSfEiRV0UebKHTSurWTR+b0TSZn5Kef3z0PW
rSMMhocrwtDwV6ZNep7B0Wq7v6tIWekPzb9GnRvQkTp2zIOemPJ+zELSQBprHMST
Q8D/vUvy81sMCjKOMEtU2vyUiUEyyNsydMAfKs33b6e6gGM8S/l+F8AQw+wlfrMD
dkc2bGoJVdgJ2uo5ufNw0rYtny3kQL3E+S/bHhtANtOaeYcEX/gs109BVksEbgPJ
a0VHXPPF/g6u/bAs5Pe+r4MIR0b/tkOO76jjbHEIFPz5NRWab6R2Q3dze4698Yp0
F8Z3cZERAVSkMZrRB1fu4f3CmVKy162R5xnkogef29+JcTw79JLE+GXhVOuJEGE6
ZzLHmeGGn9e3Bi0hrOeYFIJhK4GUZjjYiE2g8SFxJ/UnIHizaO1vUO7//Fy/3Unb
Vp4weCW7lWYVcJaram+xv/XGL7gQ/+MnG5YbO206up7FHgWc/BBrm3ifhty9LkGs
HR++AWlIoZr/eVyJaNVaixui45NEcGrsvX1bIlzX4mowiOo5/lQZf4hhVGaQorau
1AWZZ4VSA/MS63hqN0LWXkSs9HPAx/dcv1TPWz4iIgAw2c75cD4rCb2vgTqR/J0A
9aTZw5pzRhkzJ/pX8DISMM/i0mEpmbDclql5FSEuDgp0Wr81C6eNHCegUME1jIYH
V9qWPHDdUCZdiV9eIGFwVHrnlOcgwKxkQEdNatcZwmMNLxU8yHA2ep5cvlqBfNea
/E/fE84MchiUE9SExuyWdBb4xeWUy622ecVFJGrO+8OcCpWfPgOPzbDTNQpfvmGq
ahBObVyfzQFtxofZNTGVdgc13NHOO/SQCyq9aZHF+eHSe+A+2A4adMbjj0bgNcPK
ZT+d2YIKYLnx2n08IG7axv7Cg6s8m4VeltW/TpfJJiyk1XlJCdvaHPEXcRptCdVW
/DpbzOFdL+eorJXYchr2WBSRKyeGiH3h+bazNEREkEKvRnhpb3GXTSyUKJaFRRHe
2bNB8EJEUbaqm6rWFdQx/l53pAle4bJ8EzQiF3+sJp7MoAq31pB70Egu89FUaiWW
2hBtlVqS8Bqv7F0n3pCJDHRXBzs4oof5WoBIaImtRaWBUiWf3avMWDlQDzpDWKpb
gtgnPg2kUEj0UA3r4ZAuSXIHxqu2opc4hlWDE4lTq9OUPyqbBpzBd5oHh2cX08As
mP6Zc16LSMQH6l8GBFxQy3kx53J/NpWNmlFkVoZCHqltNFtCwlMaKq/bupsdMCbt
qjV/EraDrWzOoVDgoFgNwybZ8kzIFDvMzS4ViiU7pUly929kEjP9+MUeOjwbCDMl
/3Gjt2UQ58h7BdukaYgSXKf92whL3Fgs5jWFm4oO+HEPQzweZPDGHr4I0mEcEJjL
Wjw1VjaAywdzUM+vCAg6akPCHa68x9BlvVOHkc3ZsdWbQvLYKe3mxRfiGBopcgd5
MaFLFSAGak1u4JBAWFSExD3RmxETuAUhT8kDXsCmIto2ZP8hyGXqUNv3c1RkhPnk
jYS9ckUlXGEnkqdnVWOGtyj8i4ww/AV8nUoBj0yVAF+eOzfUh7cdRcROPkXwwPcZ
3BqQvKviuj2bMCkNHtoZzC3HhvaPy1xXIO/90lKEnC1opo9GioIV7/fTYTevYyAG
1M873VcIiqhw3LkRNDTeYrWTcjeSSjo7f9x1s4HFp/BUcHmsXsQFz90p442zwQ3O
sxUOphh7+RaBRwE/jtPVe+uP+RJJjD5Nf6zzezyshG4XVOTK5aE2nNfWdvJoOk0U
BNFIniAfnOhDLz2vLkTExe21o6d2qHmJwUVcyADms269XH6zy5dL8Y0GDmFdUgI1
NrLgYLXmbaU0bAAyL0tblV2x29yC8VjIbSafizxnNJnO5hpqzMO0EAayvXSKrLE6
wN9b0MI9rw0FBnbL6FT308i+M7b5PH09XmmQjRk1+jGl8XyRQbruHmRvW9Dcufc0
TZ2CW7h7Z4p+3w6RJZhnC8mUrBaxGmefkwLxn+N3F/SBMEuXShEzKmxibHyhBWYS
pElzuo74kxkmfx5Ky84Z/Q52FHLv5JXIEgXgDO4eiUGteyDG/CQ4I29d1jrIkMTs
qayMILRuduo7jrb/GokGT/v6rSVLdVHNc7WBDHuIxvzaynqGuyU1yq9HEwt+MNsu
9byr6n9L74ZZaYQtzK8zc7AXSnU/yt9imsamU6KEZ4rG6qQLO+1yivDFzAwbdd4+
dnUkXQMp/jyOQqrOjimk6M/qQRa3Sivano3nC/Bxg2gcBrUxqhx4h/Pxd5YS2HMs
YW8oHVogz3mvjRrkFoRUxPleNpnALVfGGHhOJs+KOib7W71TKrVTkTRVgeaX8sQU
T/krPrf4GVZSj5Mdx44E7z0jYGqJlfindwX1znWI+jCCile+CyQeFKEida75tQ7X
3B+kKhbW6V3PvKuaTfp8XGL4iATaLEoL1vnAKYiuaTNOX2unZ1MZ/L4PSYDAlof+
6oRTXLQ/8oQX5RE6hNembMD4SUeHjj+8bQ1k8MQTS+dqPT+n4VqOlG2EiTyswmRW
ykyFZd6LsdevJZdwGZZZiwgG0pvCgHnw+gbrV94R/ORlbjSmx69Lf4sBG1TeX3Oy
rkVuemH93oijMxexyTiVucttCz+d/tSOlAexbkJS4yOJvesw/A7iTKRBrhBxckNc
jZBnbtyeP1udnsug/lYeMdf318GP/QJkyGZ6//fFGqoOK8J989IiU5N1wWk9L8Jr
+luh+jTwua3GIoWRSPTOcBT5kn2RMM/C8aLxaQj9dKzLbSuOpvzH/H/FStIRxwuP
ZK7jjXiu+rlp1QapBMy1Y7Pf9bi/2/AX1MIjre84sa+hcxNJk8XYVDvLa0hIZkFw
0/LgNortRBf1lIqPUvaghcCLlNfJj7gdVJ26aBgtr588ZPwvzUF+a466tb3Fs20D
ndmtukOtq2ObztY8IVuC2vjC5j71rdQ73fv6uHsmKNIC17ENEJ1peDYmKzyd+zr2
SPyJtVOBx74o++QFFGUG3auCeFGjjja29ynQe3yaECuThTBgxtJEO8u/pwgH/dcD
IvFvgolaq2l8QuncgeQhk9mZ6T83phVMYgAravIXftK5+fZU3xttGmgCc9jAu9+I
xw/I4eIkBoOikceiueZJ8JI3hHfHA0YQzSNREc1twf4FHWT6OEBWkf38kVUG8XEi
BzFfyJvCXC68qhEBpkN1VJFBVF1K17LO1FqgB2Cjts+EiAqDKpe4VhOA+AznuqgE
wcOkVyGMvdZajeQla8LgJY+T2CwqqG6PLTmKI/6wQ3ykrJMyljAToUgfN8Lg+15s
aFesd/1KzlRKLnEEQ090WR8IKVl3WrnPPiTsB0dpXv3XKf5+OcH3DN04qL1J/Pk4
1isdxr410jrJ9vdwnfQJJT3OFqCUwL49gNBcd0cc+JZrgUMfjDcsbM+7G7Jup562
deH76UbE1irM0z3oUPOUfVMdqm+t7BPcqylHChWOaGfIUv+E8xtNkbGCTFH5G3cx
yhPZdUStY9JjpxnzqC9pEavu3pWuAqm7pGLTRIhUzrA6cBD9Vjayua3pzgabpSqc
wTaN6NO/PiKqasZQnxkqHDgLPvt6ZOpZ04zWB4F86JL/oel94gMGJ2xy/nh581ZR
xTb62giIQzFajCHRMpPNvEAs6hgVuK6oM+D9yUmOtbfzdgXCJyQzuhGK5RV2u71M
zCBobue+5psSO27r+VqdeX1PVZHZJH23oQ8LGD93jdokYM+JxSbhSjb/yDPxg11b
6hcOcNH309CSVv5x7pI2yCD12lUgPWCwz/qErQXDtbCIMD+y4IvkwCUmV8c219Hy
FyKnnB601l8BCFnpHVFWSk+r4Zb2mN3TPQ/3B4OHJZpuKoI1zyn8oUbt3jZrnlfl
3Y9PlTkZaaj5dr3bGHhomES1xrvPXwacoEosrbzChloBofBvfK5pffAnhPnfGuzB
sGsdMNltSqJxTfaW4bxeDKaw6Jh80UaEu9wWozRElxjw0OxNg++zdruH5C5aifV2
WfwwE2Bnmb7VAXZZvdb5cLNeEc1hUlO1Y+EN18NIGEabmRAsgca+F6BeyH80CI8t
SwGzpjiZzOdUB8YcbaJ6Qks4iOIMcZvkdeEdAMBvsgM2yI69SConinXdDc+gt9sF
DV1NK7e1XRAsHACLD4lo2oQzKRO98WOeDNtBUmmN3iWoEuacd+FWkykFyLT16prc
sk8F90FJWir1YtqJinpbOdCLmkr7IvBdyl+6V0YT5Adk+na3ba0aeNQOGi3rk3HI
KMIbBf6/K/h5jgZw/Wk3Mmw/zmuYLTJTic098rWB9khp0R6bNQWrHUy6Te4AVKnq
uV5GeasrYvIUiUeaMpPR75peXvn0x9yoJbByxhKVoaBnPTWov1Rs/ISORDOp8U1p
7HEQpRFvxtf/1BW0WftqEzJR8MBqVcMECqaiNCh9wzFP54e0VKpztJCTFpZwpwSZ
pHHBujcdcYoS1kfpejUB7Y2e1DLMFEHo8lvuejo62b8p4z5PmJO7ohdaZhCDRFA2
VFFDTAAz/55HhznSTX88zmhvuPyaYZf//shaxsp+KQeIbRt3Nro2DAsdQvjKLrk3
lcDoAYD8WP6PlvsF7DbxURZ5IbndxRvk4xyju6+icRNU+5vSl+MC9sega9O8nxgJ
Zkh7VKsHvUB9mJCdA+0EODUcngOOhvp9+m8Qxtg35KsjwwEzBAL+zcTrvl1q8ynw
115i8LIBHKhgF7oTqEtAgf/DhEsthO1IXKFGor3Gp7sI7SGbDZbyRHYjut78mdtn
AWf3h7WLnTlNMuoSe7xevNMpI6bj3Z8aQZKBvBlHnFGdSLRhBd4CfQP38muOXzke
iUSBY4s5A3BkeaGTO84x02coGjbwZU35qwhGsVZuoIeyFnqYovQMqc87WUWHoCxJ
GL9t67II+WIvls93/Nh/wLQOufBsgRsw5LEqCQblGOgLFPVzuy4eFn64z3/7Os7l
1QVe/SnotdzLCR6CnjcVRdrxhxoMl1tHXe8BDV91R2yugf2IEU9W6ByqWyFL34RT
05q4XcD3zU/6VnKw8dJbZ+LEh+MxDY6ISLZTz8b+G5phRiHfPKNYTWvHq97xBFLf
SDj+qT9JSOeI5Xmyl5idVFIqypiIuRKb1CJ2ik46pWo5BlKK1RaajPbsgAG2rdCY
qGUfIdEcE79Pp2njeNEYM7GBcHPMgRPzsvTvDtjCLuITq4GPvBp8AX7ArsHJHxN/
6MzkgJm030u/r4ec0bPvF1swjflFVpHodscPU8oJiviDRvC9bLnzzX7L/J6sAAj+
wv87F/mmDOBc1exOz64YUMWDaUWJVN3NusKvtJuOTwPfc4sNoEEI2HHp7p2WMtrV
4mwakJu0ULCPmhmZuPL4IcA5ZpUkHOSQIvZ5232tqpMnJjzSMD3IAHrbp/o7NoyY
X8tDsECScbIVE4NrppfZFNNWTPqJWYv9Don58QHVE9cVLQ7y6VOWivOZjVSQxU+h
Luf+MSUGCb1oiEc6x7rj7WQyvu4onJecpy2BcmUO3wjm/WL2rh0g59WAmJ5V0aUN
Ssd18jnZMOU73I4/FTJSd+jqT0TLHzQnAiZaOdBdgdFaeB0pEn14vZJqO+lp6UvX
iVtU+WV57956/i9gTDDVbXXTlxcpddA6NPdrHF5eu7nXpjYUi8vbI/5QMOym7ggG
rUUWOL/PjLaZYiLuu/6Wu3JyU4N9LZ/z7os/dbDA6M/q+sGKbJ+5++IwHuRiQD6r
EJHsLT7Thg29iVnrSF6acXPXLhFmlafuAvxEd4eQnQYMGDPm0F2+N3XWqNH8SUqJ
r6RAQsKyBqeU73Zpw7Gc29JzDoXZB605Z6omwruiVMFhEo8I38+Yyh7wVavoBfrZ
KHWxgcRnKRJriNe1OaeWpNJhAXzLzS73to24K2r5Hb7rQU0w9R1pk9HVyIjlNs2j
19RBMbwqpmh8BfXgE0p41Q7pCyPimBeam7B+OVZbSgwFwPjZK+vhfkIhavqWvLYd
vfZazdCjB/bLUgxsamlVrAYHHmK9eOsJPiGQmiGfgLPcCLwhPbOZdonv6OTaEhsl
ZZ8xfCQkJXCYk0TxcpNkkah0ABANesk110u/vdDx1Cgc+HqtlA0tYx5eIeyGVUfI
iVYNxjBALmF8DyEz+p9TWihW8MyZAQVZnqt3NOMkoEnaLE3uqnrFqlPjwEupUlIU
xAOq66pQB0FXPE36A5C0jnt11mVCW1yPlXSY3TZuG5cDysCGhGEovmOwpQf7I8rE
k08A3rCELn1zxEWTJu3n/jPGNmxvsCkgSYJG7KdbyanzMieJI++Js5VIhULLJebp
X58ZbPtwqm2SMniuwQzbeVn1WTPNbr+JWL4VElQx6palrx3Y0CeKfYh76BZ0eEUH
iv29wfv2LwtHUBGRK1buh9da1ybepahKDS/X46f9Ue1XgmNsiKmqS3moyU7ws9aX
n0/vrUOkP+3mjOK591AqQpNgWQSI8oCWu4uWJPYIMenhk9v+SVvAOdg0ZT6UAtgI
ukQBx6kQd8Jeg0kZj0Ry/nB8Fp2z15RYi+AaZmxAUub+3QGJx5PBUFyNvm9IymCh
FkzZ7fpRlFNuF9qU+dk3RAzGtxCeIJ+9IkOsL9emhRTWsG1Vw4BrLBUyb5RF644w
DqgvcMZCkiIMfWORmnHnPyNUBEBj/B2wIScLGcHi1Uvkrtcstc8kEdgjSEc33ULD
3hX4YbUebxS0X62LC5Fl9kosD8looCdMjThYbF8Zu0b8tJ9OBI+tMe68aFHLUhGL
qbEebqjg99rcR0Mhpi/p5z0PA7kk1NZUorDM0SNGcOoTFIXAin1MLV3aV+LfVgNg
sSF9AociwshVD0IcKKHdW3V+bbj1EZWTib/qdKc3twEcMg7qDdOraRAI4gMa7Fgo
svSGc5Cp8JdA7oNeztTtlvlSV2JKg2Zd2BoB/xhBGPh6IG1MeNj5E9CKoZ4EtjPu
Guvo3e5ajgyqWeAH9Jphx8vcPJ1CoV4iHxiE0HHpwQXhgvbteEmN7eW+Cmexd45X
PGQ7hZVgcTbJYkUl57jRAUrpAyPdUxL359kyKfMkQAGiPG+JsOHM1kuPufbym1sU
6JWstimnoTUV3tx5dqaUbehu1PST7TBPYX6dnlf13ZDFuciCs2dSIp98npU3Q5xp
DCbCroB/TaikFAO9SpiR/6S34we8ZjBhv0J0jKCk5WYCEh8v2rLh+xfH34ZusHU6
jFu8RWzOO7SGCU6XFjCBsOsvhdSvgH5EvYcQWd4gf/YygrRjKUGkFkFkUZiS89pP
AjJmvwCDWPQWUppHu3otccpXybXdiKeQsL+4Eoq0Br6JjurAX9b1hA3yYWcft54u
oQ8Ar0gydjEPdK5KfcV4wq43o7gfhx96GM8JclLPRy408q+aqFPRwFTqJxikdBad
UZTVscH8y4+zxpExGwGhcHgmPj7qHENp7UH7rt8sqxdT5uzzqxdw4EIy6l4EF5xV
EY2u+9pZNNieEoKEXQunxCX83tOAziZACMAnSZwr4Mtht2UcCaUhQZVqJj5BKgMh
IZuXiOmO4fpf1nZaL//UwPvnEWNFhvCSWjtAnJBktbSGIBlMZ0sxUUKsCm6SzMmM
+gkaCGoMKGszoN6Tqx3iQMAHlhRodLdws9DrlNPQSVs0Aup4o1J9rTp5wz6z7Ddl
ei6iY5o/lOg4HXJ3jnxtLaHPjufcRfhJ84Rck52LDAETwOvA4TJFeuSb0tWeqo+b
ApqvmQTwimRLLNg1uRqo29dDgH/uRMN+2WIROacRJvNyZHqQSiQGZ8zRdex+pbHV
HeySTiC42t2RPK69koxU3b5DQkJtChAz5SyJxlguSEVwheDUoL4t8sRKCOmnSKTp
woST7UK308pUGdWwcNHGN/prGpmiHfqoZl1tUWMyDWqXKtboEXsz3MU49nmU9eJ8
RM0Aov3QvCYMkAwSnHAGir/KMQ0zYHkrJ3ZZsH9uqF4D/uIbxCSV78Ms3sN4eK/U
wArz4Cv6+EFb77DiCNkTQprRLka5vTnmlsw+G+8i595LIJ36pPq3KnUCLFhOQnpz
5X2cVkNaa8M4iBiMk1HzTr1vrGhmzIRCO4Ck1qyN5WL2BYFU2Unq0GO9+u6JyFlT
NC+HebKtrmexPkRG275SIVgPDiAF2w5nQD9w3BDPo44AhCpdNN9jJ9icLDcWJHGX
ADBh2DLrjBA/doU1Bq5QhTZlvoeq4oaml+M6H00mH06eNae0dIt3tgKAMTglojcQ
CIKzDkNqmg/Wbep8DcjjeoOGr03GqJfjvKoajtqJOtLgWb85zPuWnODXvWe1lCT9
THV6WZx2L3dB/FIt7uesJkcqGCKeUuzbSprtzqnIBn5/jqqoBR42f8sE16JfW4R7
p3kNp5YbBrFc6A3h9HuwxJ7M/qJPMMox0EDo3AsUJafsHd8YBuMfl+oPH3ZMgDC0
bkmTllinVOHahS/VobQRmNVQmakysPiwAZByMjrKyYnoXFNg7pQFfIX4BGrKmZou
DBZio0YFi4gZE09+wCECZW78fR2EWSkkp1fyTryFwvDTcDbcU00Oac1UMLat4Yw1
hnLh93IUcxN5h6Yh6r6ZCgxVP4qgwyz9HlP//bJFrErks7lm3YHtQZFKiXhXG8jE
n7nfvBc/wGxc13VepbQvw8CvFcFKIJyAwrSC1W2KLLhY0f8vdWM4u1Fe9PX/n7AO
Bveeaxlznq6SpHs9UoE3ax8VUsEFmJfLixzym3KKpSNX7d7EZ8tnau0LPQmMXPwb
fiO+NyNJlIFoRdh8e6bHinH655x3n/30QkaHmKMgewT8u3MVYnnndv5hNWz/p6yS
0WHHvkrAXz5CmkdkICTTGGKZNdXemWU/BTLsT8LuF0nn1h+S09GbngWm+RAYM/01
9aOXPN+wJWC9BmjyPyBD3cxC6xwtpQZImfhI/qo8l6X8Do7RiepnBIIqbXM/T5Bg
ClijMomoB9xo7zwT1okJGxidNUsP7tKt4mvM2pWJKORlcN4V1UvqvMIaorhaO3La
f7Z+BrNiRnRnBMnk9HvRzc8iPb2loJqsIBEAmCkSgm4oXsAzatQMNcicPBxdmPOZ
2hpbzh1HHL/aNMm8kAZBtPYUASYXtTQ7y3PJv7ZIX98IqJsaF+0dZ4t7eCJytKbr
vz05aQpyo3hb1MDbiLx56jZwNyYSoNrNfC2Y2iotOnpRXb9DZkZYITebF3vy4fB5
/g+IOeYPhAD9JJ6XBlDXDaIvmJ8NycTmiy9Y56I9PeutxEFMtqufNtnf9EatPyQG
8ShOEVuedQjZeMM/RKziSVbyZQp+wmPFrZMytE5UJzmeZWhK2/xkYwkr09ok0vdq
5Yoe0pzYvNhuPPus5v6w7Wk3A1Ud5xvhhkqMVGyOeuWqn4mqUaz8EXDlizaUy6nZ
VppeOeoYHLuL12dwKqntfKhhNCXd6UX78dUV2sZUp6kZDrszc0YZMzTpgAiVlMXE
TTZV07vukkf7/k9qGz5GevTbcZhO4PxMjkYTh1o/s3uVtAp7uWcvWCy5h3Go5u+s
1sbt06dLRj4dyf1kcWHQ/tj4rr/Cz4aPuLzAYFseWaSl8WMK7wesjJcjMkNB4ljl
l0ceNSLTsdinmmuv7VdnhE9mREgrVm2Xq/9Ukd6fdP3KGyViCrt+TYrs1QHyG6m0
iu30+wJBo6I0VZLMh4AxwKeWPUZRhwbMKkjilLGKS/R0732Q1fP0CwUCwqDZHpH6
OOKxJGmXfBFf3+8lyqpR0VkQqt8zVeRWtE4vJpbjBQZjra4v2YCx2WjOHx9t8j+Q
MBUyADzZpeSI/gomOL7pdQHU3ouDgM8w+Uk5TSP++tALeYOC51qnhbmhNEMAHVre
10lDnrmoDO8cI+eGpfclyj4LFEsTJQujzB/9mmDu+J0s9YZSiQaqtCr8mL/TgpDS
XtLPUGdtz+H1ckfoXfNyhOKK2IQ/o9Bje+a/xVPyuMpDBedBtdSqzzLoaJ29Tfxe
nawJwKm3j44sMjPd3FS16GxCl1N9v5aBy0B7uILr2L0IrSZOhA1ZxjKCPyTWj3/W
EBrdnGlirr6Jyp74eMXPKwpYXO0OVQlO23oEc9dct0RbmcoVznsUB83HfYnQ/DB7
yU4WN8vvNBkinYsJht4p4iw7qHuoZjJK5eGkbceRfRW9urZmNNsIwUnKv7UavbxZ
WjIquZLtjTMkVihhyMtB0M9loz45VsLWutjJNhpOxrUjXYfNZcDJjcsKWYtraack
cAIlsKTei2iOTvqwuFFrHHSU6GGOlKCjyh2DlYO9a7mk5iWPlfwnLOEz1S53F4qE
sdkDhy3R7H20tlipoiRrztF/DPerhhdmKW/5mYT0OT+5hKjH1pCUtcPXVeKIIOT+
22tCjrxBFsKHMm9Bq6iuIR87sfft5wJZsZ2bNxqh7y8TWKPiLEQbIHKK6I/g5IOx
LnANIUvEwhHMTV/UQdWH0WIBdWF6JJ1hpAPtytGxVj0UszajSzDL2oMSlIkbEqzM
5lYvMv7rD1KkOsXU8ZbYGwL9FMn3OoN0fnm8R/FUB+CB0TrGI5kssbrwTgg3VC43
YsWG8lHrxKPwAJ46dOJwSJ0v8tKYZr0rh06DoyHWWsvg1gxITLAZlZspFwVX2aKY
ejnEV/yxdXVecUUZtepre9jjC2JsUX7Xr1IOHdTkfQgFNRvi/xcmEKWKT488RdCf
9lyk5BruY2iuZTHYnDMeAL3YajU/VjZf0RcTGBU/GeUCN+GXebv3JY2zygVleQvW
SFLCZt6grW4yavRt1VW9WYpfw6wv8Ya5oKIC+S5Rn6hLH5SuRRVT3lqvAbNrxAXR
PKdYtA8BGfQ7yyyFU7nY5pLNoHH5AJ3my8AUVDQYvGsB0lunQWhWDypFeHbRuEOH
zbHU8UWya5aMdOggK/avRE5TIolOLApC0RLY3+iSLygyUns1FgSiXRIwq16E7AmY
5BxPeo9USPxDAB5rF79zz7YqhiYVOA4HGiY1DFO8m1kh3oDrRcGeOJn5iH5ovKhw
0Q+NO7ScQS356IcJEWzUzbEaJafVy8E8u4D7T3fiFdKV+sU4U4mFbvqur1qjIIOV
jiau2TuPzn0NiCfLi6Tp7ih6pKgF7FurOZEzfu/ElyChszXgFyOcx088Lnpqt2rk
xs/WAvPJk0w3clBkIEJhh8apEQisHHu4t5ZCb0VtKCob5k67wdCVXtBktCR4MKP3
8EUl6nbtAKvD3JEwS6DORnIN/7/Ouo0k4TbBq7HbQhjPnkU8cOgdp4SRp1Yu+Hc/
jhDWLZS9TXNs13ylHAFWIwshrJEvOoBDyzf5WAwiSgia2CXU7x4aKvCCD7nr9Ngb
l1WNhI95n1GCz8WfTgEsKqWynOlaSci8/6K+Ug3PuW9lB6Kj4DKdQidKRPAuYmAV
C2Kmfd9J+1BZP5t5UP9RAW6Y791Cer+xIru80m2b2tT4zFg4ZIeTggDVWJNh7BgK
es5tZSfSMmzIwwGZQLzgSPhdESUqlG0dSA8a5RpyrurMCLPnV3u43bXL8MEBitql
U7IckoWLjvnaHy+BSEKepgFTnfRK2MiGFjTeWOyI2qg5W3hEhjTFNTiUaqeJa+ci
jZqlHK/1N/dxHnvD9oKFD+6GkoM7VbDylgjp81Gr3MWr5OVN5wzIa3qC5Xwi3Agk
4G1hMhZ6ovPDxNaNqWwDpVmML8tgBGGam5fQGmrT/TtDt0uWzpFXpaCCkUgY5ZXo
3OS/3/8BKXW9CT0I78eOvjGSDmb36CqR05ZG8IRvLztHu8ANSzQpOxYjdmc03MRJ
oSpsO/iVZnd0Cd1JsqQvqZBjuXLRHWVEpNJqTdobY3p7Sv2znrDaBKPL4KFlnrkq
Yu2AHrcSnm8njplwfnHphgAa6CGBWnwVNuOvhxwQMIZjlfQZ8kXJmUFGjgn4CBsL
vlOQi5qJqtbS+t7g2jh81FMjGi90WkoBtJ8w8Ei0Rzn0sVPZ94ohdv5fBeQDAhW9
ABvUfLdvRMs7VzTJseSWa3v5Xm6RVKrHhHtFemdhVc4vBPpY3xjbD2cwDUzxddwn
pQTZW6Ytgi54j7+BnF/5H+GIZI/xfmD1WeOhx7lAL3/gMhBAvmsg2BPJEo5g3Xk1
gqpXS4TfjSWIyFSRMuFeUEkUqJB8n2EMFli7IW9aq+DlXeyJsSektq44sm07imvO
IAcIZiMWl4XMuFi45qiHYhEdH7F4xSzFuDiRjYRlCYUzp/SgmGltAqqtu3/Jzxf+
n2MnVJZy98vXjMlHVOwVek8tFpDFJNVICSvP4lId6hIIQHc1Waf3L378qxIxHVDu
jKOs6Z6ich6+FbkkZ/ih4kpOFhWnTppgrobUBbu8wIHl6ehw7aD92Pm9Kxavxh+G
T2TjNwcD5DNriG0qFXXBRnvt7kwfR9lwQCzCpySMnlkYXVg71rqhmITSqDW3ZYrl
gcFgA0dKX4zUgT1fIZtjOS/ed9X7uQ1CCYNhRZp3tamZC7v6dIJtBNdMRcNlret0
Wu4Ob4cr8g/WGLJOncaLkFv6f2i94uagIx/qXBYj1/2/kS3SpO3blNU92uvRbC1q
nJi4Q6sAtpYOudOQrjnZSMu8LAW3/sx4dx2MwN1EeqKAG8JkYt8XfXbIPCxGYGFh
V+dPhC+zXc/KA4CqmIt//F7uavA0ClxtWRbbyc+ew0Iyivho0Cd/2TgtCouueb8n
3xejYCIELnT380XOHXarV63dm7ioKf+TDjHJTdF7sz+4oe2c3+SalVL6Zgn2lIsE
XDtLXPJwChH15+m8LxKLKaJYGJyQ4Gv8H3hI39vmEVWGHcxyMTA/SLARary6GAHA
qh3cSdmGKubHAZYMAnxEKl7wBwFHWFrBbyh9Rwd2NBCEeR16VwsDwNvwlTrPpirw
NBrCw3k7wlehndjQCyGVds0MD98vdbopxQr7xAHkQGKnvBJK4s7mVOdAOJOwlgiG
3oOuc2tPgvm0fqAZPQZ7D4TIU8BiODEOM4Z+aBjh/F2zjdJ3DhuYf+NUBX/2st7Y
yQCtLjnDSQJEJzdxBmjByzFz1o72bzPcO3j6oQwE0+S4k90BRMqEyOkPBCGRg6TD
99hpe7myoxsx/eTXYysxKlOZC6uz9cRs1aJUT9QKUWsufrEsaWaVGtdgDYMNL6cg
SS2uI1OqRaRhWuKkcTX2ToyFEr1a+3+NGKosFLqHLrSEEPpNPd/6XobdDiREd5I0
gdBU0w2CJg6fZnTCY08bFbrqLvjHihmUFCpDUwj1nd3TDvYFCGqt+vsV4NcODvf8
t9eCPIRXn10dMp8IgdvhPeprS0nJIQDgvdu/tn3jja0ZrZ5nBGEjmHWh7SI0Hsf4
82m3zQJsOkeuR9NzmVxKIyHMiV2oDkSAXVlfxdKrqsu+752LYHf3LhAjd+dbFUke
ORIrKOCRlZakhz7NFQviWWEW9Z+waQnJ9EPnxCeDOg/SEOJACR5S2U2pJZL+sWvI
d5b4nyY/RIWKLQbsCzjaF1TmEy77U9er4fzbBKOEeQhAel0EQy9Qbsl6Hx8/laAT
akH/Q4eU+AHJ7Fx8fQYV0uOIprUymiQ/MOwxH/DXD4l6X/qd0j7MIH+Tg2L2qdEg
RQPH/Y0DVesOrvicU7katdFMqdXVzr5td6NS+Egqu5v8bc2v8dCNzI80MKD7yjr1
JwvG6lQtgXIrwjkxuOznojabIl2rpSfl/pGjfzskCUHV2hPOnm8bpCoBRprs/Rbw
nky/CMx4Di1/XB3qDkrg8earKcVJ2iSR3cbLywqNRnq1uep3iu+IO7uj/kvr0teZ
xonVBI3iurq5Rj5kJRR+xLR+f/raqcEws34OeSPiSVdckXJehpC8NYU2D66xAu04
q2qLjWdSDyresP5etCjyNYOIfJQWl/USnHxrhDaQoHnBW8tlNyCs58an0sV+EvOk
f+o6WlxQY4cC2+uSDmTr0Zh4L44sBbnr5/ZovfKs53Ll7SVHOq/+0d+1mj0c+hA9
w1aAMy9UEt2chwIIIJAvK0cjEM0u4i5zaghtPPW+EeBgToIODij7xfOpxoLsBAJw
XCUGoQO+fpzvOFneaBDUimZ9nRxmecO+3vZTeGe2HEG+FegGBrt+X9DdYdKU0ROc
uZxy6EYb6a/1dsMl1IPsYma9XAPtGhDt8YK6q3V15RQxuFfIN+rN/N4Dzo1qZeen
zHFECoft1XVLVHcweJq0fW0nNrL8BSRn48fNydSIWL6ZE0dYqdomPbN4IAr8vP1q
UoM2deAfYPLtd9X7F9kkwPuHmIp4IDPU3PiBeNfmz28v5GM68S+rxVG2+lPsBmA0
eiAZPQsymlKKQBAs0I3+mOAGouU0fCUAO2WMs1boNsh2ntCosan9+m7REzmK7zCX
xMdjT18+Ms3RfzS4QAsMCANxul7K8AjLyMKAP5UziR+mco4GMOqFwpEHFJmTPbxa
OElG2PpGjNY8jxswuz4jJewWENL3kKWDYeCf4lTY5Lksmhv++qXx/THAG0p8Xqke
BbA8HKt+me2u5B0sl4GQ8AcZK5jLFwY/9vw1ibszyNrmslCSjJcljw7amFHeDTgT
0d+bY+8OBs8dTEjsqDc2vueXnHgG4h9DFgNpT7zrkUk4h6HYdiUlbYu6ni7NlTNh
ZEM5xYuZPriQtAbgkVa6Mu4t43IOQ3gx9YthYD9CozA7eJabMsu1tYaXLLOn7GrE
xwicU0tF7u4woYiYjZZ1fQhAwY8If/P2UDWOvJ0QAHhfgNpR7byBXEamdC2x/s7o
D58TcrxXuQvTmG0dG51Y5FHqpQR5rylFnMscIpIyR6hewjdrLvjMuoyLxXqXC5+M
yPwv/D+8w+9n1he9yu1a084NEk85AHSjlOoMny4GRlOFd01iErd0zxLmuGoBgbmt
xHOTZLDnCpSyDcoeWqEduUwB5YgYKAesGr6idYcEVSchwf60ndz/lOsXT7lnQHHt
0NQOSc+/A5tDC+JfEdi3t7uJMbXIqD7cFrtkPyngvxGwZt7URyCabYw1uXChWrom
z9CBEfrI8W69UfpoDrTPfF7CDOuHgG4mzfOisnxDxXCSQyd7u1f9MabO9pPShwGv
S/QqRdhNfj5yXwiN7SfJJ17WoVCCt8PulUqfKiO7TnfLqcIPbv6vhRVmGC6W25Pv
EipoIt0lhyY9hHuNBvvKKtGHwdk2dSev66TJgfc4AOuWYKBuG/DCRcDcI0DcNtWJ
5MsFwrko4Ug1xRed3BvPFq/c0HTTAJhms7O5iOqwuGIRZi5kFqrMoh3Kk5K3uNF1
En76QyjDSdVfACHy+V9PSmyxaoyUeOl3DfiLyl2mWGu+VjkX5gI4f2NHgYDKabRr
GkXUqEbdpsOli8g010mmGyhgpDzjG/UlHisd1YDkAL6Fe8Ybj568kkRWJcefg8cu
QRlK1zJS/FBCeD9ZybYSSWwqt5wqjZwB1p9i9cS4xd5dEQpnh6oMIC9Ne3LMoPW/
KWMTFDmhmyOMamwyCt71FSqob9TLH/VpgGQnnPiU49ns7zCW2YoT19L2vSbCIvDu
2wzjUhvGTppYpwmWgeVjCszaLgvopwX5uIpd8tRiqKe3JTMHv+hryOkGuCObVYSv
jyb4DEcAaWfYcdB200f7/PJoe7SWaOPri66C3/rSyMNQicCnbIwaoTRxx4nP+0Vz
ejAnUdYuG4zo8wphKkCN5sDuLjIk/yOlutR49+mNixROeoax6XkjKO+YqMQz1M+i
/YnG5FX3kIQk/P2J9u1v3JvU/wQ2tOOwv+PHX6BGFFV0imOqGUYNxhzeUst1V48O
uUIcWraIFF7/P3cHhB75lmUVb63U+CnEJqes3kAA9imKGvIspIaKa1uEkmcVTgzI
8LlHfo+nTgTyRTs6Fjd/9VDIlBCbOOZApEFspPVgOoV7YkIIRZgimD0XEEFsQS6Y
4s8G1WzIIuUAbn6cVZhjHqClv+knIcfu/HaY3xzqbPUjzhIDKTGb+KRWP0KWx5hQ
UWA35UkoRKBNdbFbpw/mfRXnp3Vdzh2tOK5K4UXeeOaD7mj/O16Tic3wBFejP7mm
FfueX+HoHgVc1chvZc8RRVosHMFdoJW+0LZSJwBppsN3bnnDtf0+UKH0OLR6md7d
31SGrsH0rHkLZfa0Ya188N0Kx7jbIxiPohcd3Xqm6nyvNA9hcBBGaF5CvZ0GCeA1
rjl0rh200GrpvhEeheN6NrqrkirJHn1krmPs+DE7sQZbZXcmUZY9VymqEyMsORQC
aCvSMuRDfy0OxDTKdLPbQySqxGABcqRM8PQ7yCodHbEXtD9daWxXvSFGdEHnk2Bw
74vFolo/SFFCXFBiXm6B43fJ7Ek3dTkx700Ajn89UDSemWHMFP3oEBKYPDcLepI3
BzxgJj0DYiS/JgI+t40iQhbE+xzrbLgbH9wIqO96SJD9wCuQ5Y6GC/sNsPUcSR4p
9nW+StA9EZQosjTXOxrLylJoizScvdm0u9X2/HZP+d5+mTpBvFtaR6W3n0u5HkI5
VXnWVJoJ2E8Sq6pvqtOCeAe4+Dr8gZwqIGi7B8+AueooLIwECKx6CS6BHJi5d3RW
+SwtHG2wohLz8oFys8ZmR16nf2hdAC8HOWlKx1gX8SCBAgahQT+A8pizDX8UfSZE
KXwsraGJ8hLZtX1MGxbWOwNUwwB9atnYOrwNGDBj4n33q27miXypIcAbD9OQcMFj
rbEiJbWsEZemuFRUMwJtcAIYDOwHT4RIxb5WVvL0XqhT1DnmfQPV83rQeodcp6dz
ArTFC1vYnnIGDDGKp/QkPCUKve6hzsVH5qi44MjvZoaYrE8/9EGKocuN1m8/aQu4
0UPdjOfYIG3sDqH+Msjp31735frh3mYkFgfV//tkdmbHcVR2Hw3hw9L8x4BPLEXJ
qdeTHILQdBEVNQPg8WjiI38jRgXD2Wy9fDye2K2LgEiEFYqInWKDFt56oZWqbiIj
DGNuynBeD/2uSQL6SuDTd5355XK8/MZQTzfCrTYW7riRjwmv9D/KhrH8PmdGOj4j
wvUoI+6Pr8xa8oTnH0TDQiHU4SjoB5Igt8BEOQZZqJvTEnhiTc0cSth65p+z9T44
6/0lYj92YQnFxTxMewYNEAUctXl53oxcsXXZ6vZSYuRoIbpHVabGxXzQPVmFj28n
cnSWBgw6F4hN9GC0AzOyi/uKQJQpzmyfmoW/mCifLG2XVSFo/CPnZtRlEm4Xks/r
B9NGVGfYMlqIi9yut0KXHR/hQ5EM7/c3TkzUwsI0Uy1LU9u6dHkZvQunOe7TPfSa
3FnSEtzS4Vt/gHgBBm3xuiojDvqvd7uVPoOgEiSv/QLp6NOfDoOBzEm2OOTNOgdl
tpiFDVmYyH4EIdJf7euw7KRHn3chK+myBt/BuV5L3rY654kBidfDBaqm0ZC4eA47
mZEDkqJdmm/K/hx5Z33g8yP9JMCMSAKJT54DCBCpAbVagK2ycEXIPZkCsHwxhR+M
a7Auwht30PUa6ej+vLizalc5kXvcjGx5zlB6oCEywWSXm+Q+VcyVtSNqQ5Na9Omk
4H80zbQznWqmQhvpGJVyit7cXbjAvtEXY4Q8c6scgMHD/bPnmD6ocbY3kpUVfyK+
s+HdCwVNwDp57zkHrACKEOeKYzstHtITeJE7EMllVC1/rCBeH0apxYsyk4pe9FBQ
RjRfVWPsBVBplvo+IxlGw7dpT46/86XSsUkee5je63PrzrlgMWMIVSEX6ygWwcvn
tO/2YYHEwXpxCTymgYmYVxbGBwfY93TI7d7sf2KmKR4zNTHSmIcBaI9mZik4G1C3
Skz2R0Owozf5+fAh0P7ypWOSZZ6ObVFVlcYU4338USvyxYx5lUlNMyk3C+8N92Oa
GLNMFr5nsmj2+E5A/wT23Qn75rmqEDsTru51plk2oyP2Lz/KmbiFsQEEMofRrguj
jcdkoWp1t3qZ6EgfbbeTIrvydLxFZYw0MPPXM26wZOfEBYc1RsN00dC+HGjwrO7N
4bDYOzEPCoXLIpN+tnxRA0x7LsShmU5jRLC3UCHdZMLshrVihyKMMcb85ltqOku2
Zdjpvn0gtSXOsbtyWeoJM4uHhtWps6rQAhXNrp9cw6WhSOrb2ZWmGJHXagooMLPR
pXUQ1YWK4B8sex5eAZ9QtlHQkhZuurn9ve/NiYKOaDs9ruwQyReiTLEi96HZyku6
RTvTCSY2cDs9wj/xjOyH6LZ0OhEs2gmbwhzVWeNnK0N29YYON2t4JpeccdZfgvLx
GC5CeWOEOEAQfi4P30zOJVxYEOvtZQz0ZwYDp7ssNKlO1T97pPwKsaQ4W9a8Gap3
+FJoWhOvywvsjzQHOhVsHFKp79Ry7N56DHfLBxeNFA+vLsyCtp0t54pcE8zQKBFW
B9q+wYSSkdc6JraSl2zvFbI8hasjjFcSGTZ3sg4xaSFwOopbGjYixffw3DOYTOj2
kPEm8SH4JKUfHh8nNBTcEq9rB/skAK7nzSdEogyxM+SHERMMTgePiOrItDBSFT7U
J63hY15k2p64dT30yRaryVgblJTqo+d5IPSWUI/BqekZGrRslMBx4YN6WmuI2NET
YM2Wvcgumu60xFP00FPDq9UwylcrUB8JXF8nE0sibcV/ckd1KR3X1F/B+4FLLTu1
y5lVXaRLJPFn4ZGTPowtE9B1GL6BLAUDvyw+qTrSqkJoxuxkYLbyOJETA3IjvuZ4
Le4Cls0F4/YZfz9DfRl/iD9+H0xSgwTC4vpRz268eh1G81XqhnQ5ShqdT/bsylVy
p5DfjVFiR8XpD5OYS38JPKI3+waJdYi7ImMovsn6Qp3Vy5hh+mULz7QwpCXBlFfO
haSVUy8NNu1bRYOCLbxqZYEvrUPInM5BEc9gRjrYUW2dVwCDnHsn6Mo4vwstMCXz
vElllgtsLbu2ewgaZ/JrnH+Rr7+8x2C7Bx6dxhDs6TIJ26IApZKBYwptnsUrx01u
75+knVxk76hlEuW5xqTCyo4MkzuIcuK/VUHt6I2N20an6ymrAXfR/c/y5D5km6XZ
RU91BeOV4MvoUoWH8NgSq+clt/wSv1XDlWG6busHivd8wQ66wTykb0moH1AucbSx
mapnZTWRPgAAMkxTJmhNJlYu9I89JS9lBk3HWFwHnlyUtYGUZOmDZyZGwKRK3OAe
1ZZ/vhY5rPujXGkDuvW9h3TKUMbjruFM8g9kLk03vhzRxVmuFKpSLXD1nyvoB9Vk
7vAXrrC8qeabNb+adEcLcgym6D6AMg5ZoMkBO98phW9B6FUJkFqJM4RuGkTBkIXP
UUN0EqKiBMuJQNaoEFzfullM7Tu/uU71twbKXPTXJZMwVxUsufhBIgYxxvKUArOO
d2+fD1/N5xhJx90+5kf/h87RVq2+XD2OqQXalT7XDSsaco1XgISzwI9ZIZEPGhQJ
EaHq1lVgr+5gOeifDvDekjxt7vpz7qV+NPV8/S9351JXBHgM4aiy4F4/zDCYsM1t
R1rd1NDWYOrqhZeERKcdgiHvTQ6OMvi/JeyqFwbaoTq6+oonpT89y34gAgIR1l5P
UaVSVZWt4a7eopFiSHhhAHkXHLcukmJNMXmwZIoQrSQUcXNJt0oNPz6mCd5A5+UT
ydsNEKyuMtY1/rsMwiXc8FgduzB5HrTu5/iK1/wn/JfFLA/LfQ7t8aWEUkQ34esl
APbyBD5dueu+GxuViRrjZ3jOp91mLxsBxGbFcAkZBazGtcRu8Op7egdCSJjjwYlH
2fX3tK3PxmkfbX/o+pBQjymaVAi1tc03oitpvErKa4YdkUYXBI8b/z+2ZavHQa88
OHE5pkpdE+RYP4LBo7J0WWTfztvR3f0gWMRi6/PTPjhGuhl9ruScTP+scVtSygnG
3l+Avb9oymq3PV+eD7HEvnSYgsSSF+vR9gM1+rXbNUFZu5oYRjZZPUbaHMoC57W4
Xr6O5uqJP0KeXYAscwd88Z3kAo/S1MSG8439zDgYn4cyrChgPrkikNVMtMxYwaHG
G7ACi1YItvqThtf9A5PhoGpRzpMEVHeNvpuQ5ynVBpxgX5cigTPexn47gOyO8qQN
B6brxCQpxRcBR/vfX37vOewatIVK0o11f9a/VmT5Wwps1TJmZm/Tx3MK8614TYpc
YI4ho8gkgmXDd+DcalzCWdh9LiqxP8Ul6EM0bPemP11MFc4t+JB424cH3SRwf5Lw
qzk7A6nrNvOor1D0tkOH9uCgDAAL0vdtVTjgjwr2WvvV/ccy6irfiooIK6+QzJ6R
xbPodP6qdbeWtO6h7mTj4v+pTuPZrNbjUS87f9C2j1UUYu07J/4VHN1o5h43V1it
a3K5opXWSQlgSwV2AjeIaK4Kj4hJG+Hh0cFlZQBP9vy4/kVswU6oK/iPTpUBAtfQ
aSp8/fb2QQfOetVI1uQRO3aAUT7247BNMOgQvy1psw2NZYepH/fZ9GXDUmuHgOHo
F8vYFApmBnTPbbom/s2oMoi2SLPPxEPf3VTNrOkIO1rr6lDZYxhhCzZhWU5iw7O0
42VB/oqe3ld+YMQZO2dZgsWF35jkYWtTBgqFTy23u2s9ylUyT3+z32aLYNHM3sCB
MC8HfUK8iOzftdqfnNnaT0vW6BxjUJzasCcqoisbkbn5WtArnj6n1zsBrrdzs+gz
wLKdDG65bkmCjTuQEFzgav4UDlgH8nvCPjBQoI3YkBHt0BQ7jWCzybizWvcNhXni
ifacpydUMnhHljjNmoUGzSNllykRsoPdn9VASErgwB+BrpxPrrUWKvYYkw1O2+ua
DKHgqdOIci31Kioxb1d9Am1h+Zn+L1urEkYyv4kiuydeUA2e9b2l+8ddouEdb6kX
M27CkoYUppDgAdau1K4qw5nfICF91ZQrt2bDRVqKsKASAaMkUt5OYlydv6hd4xac
lX1A5fhbpP2WiwjttNbbVazMbpEt3OT+tNeH/cTgqSCdAxS/layR9ngKRxqW+CJJ
oUC1g8/q0+BwjlPQlZ0eamKcQ9Di+uVJhKfWjPHhdSkhax/uhT3+/jCNI/B5MOYF
kjv182vPXQl36ojR1J2Q9TXcwenV/qqeOSpUR3p1jrElHIydZwiDWbz40SoUG1/Q
mHflk7YPD5LICee0oOfivivYAOOybExXz/AkybrEHG4OL8czKQx4zzNtwmgg3M7O
4nD7e+QnE9SiCP3cfQK1UvQ2lf8HwyQj7ng0/p0cvRmpYJfGOf9y5Bl4wC7GWRAq
beC0ItlzsQJMmC37pPh81AjjwmWiIrDgRTvpqMFvKzJIM5gOe42ypIkxzwHx/7sE
vYVhZl/o0r8R3WTYDcKb3EpOROn2hql29EpqilWmHxe8wGJ0VU8aCzyo8k73G2Np
u47HI50jyyF89n2QL96bxliMSxXFzDzhtNnyvdeSW3egVbn7iGK8a749MeENVOY5
mczmZxIDPN8GOLU49KGNeGgYVzxlf5RwhRjqyn3yhgaMuazn9DGP6XDV3E9K8ru7
5FRE/4vsrVJiba9H+XFEzvO5rjDG57MWUaHM5nopEqdk2Tv9a69Qomf31+WmbkWQ
06K1l0f8w5Emz/clAnxTim1QblJlO+/cL2vAWBc390bcguM34OddDvGfb0U8UbDk
ToCDN3DTEIg+oPOj1PXSdrhAtWd/oHmk7DGgbB2X5IR5LVDG4dwADH40QXEYUnmR
gGYzIXctuVvO+0TkwAyv0pc6/w1ipsYTgXE1Y58exN6vGtudLDIrDV2go2tct3I5
GLuRls0DFrUXtZ8HfVazKMQRVLF4sjQ3OvatQcfw7zCgAJ4XpG/RrUC0g9me2UrC
kpZ5VR0Ze8QwhKFpilDl7St6a4D7xhnhqlOT19neeLsRcmR8Y5rDjhD7qQxq8fXQ
rGpDCenHZEST3ACFECfVTg60xnTFXjodunxMsqIyk6eiUyrsqFrUkdqK76qLcAi3
kSMO5rMsENZNPseAMRjsU3BpdkvqWjtEeGn/Dn6neF7gk67rMrOvQaPn2s8bnjB2
2Ybp3KekesQ2JPslTU+ZBnB/zOEwyNfD1ta6kbWeVn2xfl2AZhvQDU3QeNU1tMIs
x2GPHIF9T23uR3nYcIpjkr5qR1txUdRNv+wlK92S/XJsYnjDQEwdNcJYjhwBhPgC
Yyy1sscd4e9a1jZhg+ebMdoWyc7yeBUF7vseFizBDYvGWk6FNDa2HEV+KgRltxEm
YjX0hSy1ZtoS/FcNSABmCsUVooF8qdTZSlc2rq8K41RtOq+puBnLWPWjqWTE+ZAE
JAsqaWNx3iWfrjTqWGNvQsJ5oSSlLEx0UoAFye4d7wgDaHPnvlXcgomw5ZxuzzU9
gWTUWECEXJn4mglfRSaM3HSdJo/ol5bCZ1SaTv+AzebFknMSNiCA/9nTB/9XSAY8
wBvupa+FYVB/LZcCaon/H68wftEqqSDyHrH25b3C7tTvF2lKWDLpHgIYN+aqow0k
KbwcAS7/cnAejYttpNEtx682e480nZXfVLcOWUipDxerIh8gn0fc5eFUfYtyFUO/
ku0960551Kb8RuH4p0xeoLlNpIH3leIO96pyv5TRQw2SoOljvBx8g9Kz/lP3GGk1
cbUkbz5ee9xayz2gjTSBIb1z6IKZmUaEk6/KxgBjFb1UC+pYK28FBSo77839VN7T
sJSyp19mrSbpNeyHqsBCKjb0x/2AHu0XCW5jkP3R0ygt8VuAckhPCTbbsRHxnGtN
zHwqttkMjUb4Bbcg39I7kXVtaeB+aIYwDscBkVP1dnbrcYLUnlnxN8AWJrgGr/9M
J0dUFx9CUxDkexx6zcjExQSg0Daq0BxiS+tT9Nzia+uuQp3i7nLOAabprlBrHjk5
0kA7PhspN2VLlizRf179CVk4WXpe/Bw1l1unW8sIBiB02/lWFEPNhjutG2RUgZFX
8wuNHR7rwAiexa0NkADW3c44klAp+AbciL2u94ZmTGp0/qmeJHUeT5kc0n+wC3I1
n9FfnXkmcO6g+EE+BlYpuGIxQ+ZBZ2lytsJbU5piTTOFCJymZRVB2bfwRoNVwYxD
fWmoFjbwzJ791H3vVQlOMH468oF7i9sT+vv26+im+M21FlN5VXYp7GIHwLkEFpMn
HZj5dtlrErejvZ9Vms23XvMiiFsLWnZEbofpYbEslk7MOPy/J9wsEaTo/Je+1Iim
bN9s6tQbaxp0RAqV/C6tfxMufAy6mBVW9lNiOAlq4NkPMAgyXpte3DtSeT5oQIYz
mmGRZdvkKi8uuYHmVSAjUg+BkbFHKHIC6DeGVFoO2wYdwXcwz6WuxHb0qZjvJqr+
W3uZtu1Uftykpkyqwuvgk7AozxL0OyoImxSslw35n077177zDAiuwe6HsKxSOfM8
iRMO/AWKwY8TLnx0Eo5JbVT67ZTjZ1HepsF1eQEEPINg/vCIQq0o/9fWl1slVH4H
Ulhvw+2VhJZDBi0Pxtah/4rZsELkLgeq+wd1kYb4MeGHd3UmpsWv9docppKcfsAH
VJXKijMegFlaO53hyqmtzfCw6jmmJyLhW8VfnUz/+/flxS92JQ09izyQ7n5Ty9wW
UNA2ureyizuMFBAsmqZzc0WzG8I73xRKZzyI0pBEFLJvS1UsmjWcoXH5ULOJsiPc
vpj5J688U8ea+9CmHHEhuY/cZqCUhwJWPS/PIiy3TiBC0dJ/z4buSERZTZOVzYzx
BNiuaNNN4Iaae2y08vVVV3GxoRrV9aR45YuoIwbivoIxCbt/nJuPTR4IX9r4negH
a9YxVokmpWHCI+f+iYPCCJ2a4On18+ISeFFSYL6IC8C6Hhp8tUNsP4tcuIk6wXVA
+LWhUoAD1h+ZVVCc90vbbVWzcYwE82cLHgo/XbcmzM6k1qWGhtWfoxFc/lcatfvs
BySDc0oD6NU37tkqOC6tg0M53ixSx/MXjna/YcfWE9/hE8FOLDzFq74IcHO9Wbxa
yBYp9e/8vXgHx6tf+cDPHjaOJzPKqIShqFYorWfMwCgm3J/vwi+KDTfeM0nEd/j6
yDXTKGS5ZBCGJvxf7cbZXtyqhzOaDvvgXlaQDVZ2gfrH8CCSlJkyhcKtX7rqYXhP
eBMezEnNJWnJ9VRZiPJ+YIasESqFaWh/07vzaZ8qkV3mTL+jGi+qYjHmjpKjswws
zgWdE6tF5D0notAxf/Toho9fJ7wUZYb+lbtd5c6AcwuuYXPIzvCN41GxyIL2IaXu
Ab6WrtjOghmDJ00CqpUQ2kcjizW/hDEMPdUlqFyAvSe3nbcm1F5ts+ARUKLFjWII
tS7J+mr6Uo57aVjLUd9kQCSrIDycedM4+nPVHPAtyKvb2PpjRFa5ievZc4lJBYZI
l54sREB4JTU57J2PwqiRIuJV633dh7vAoxwvEhQHCCJVJrWQygXPvznTCp4ZQNFg
TRraXACX2koO+fgaZgyt9xEidcPJ1KF0HvtPB4PoUsr855hG72c8anl9NKbPfQAm
eXETzQ9xTum8bhHJFblW6QcvC94gsWXhHQ2yCCfQ+hMP+EhAmHYqrq7npUjHij6a
RrIGDjc5nD1eWfwZJ1Y+YbKoE4PEYG+TbyNJNgVSJKfn5gPLUZuLxB4VtL/hBhi9
NiN7xQiLlBfRncQ0ERvLjTLc+qlzr089Xd8yPOw0+9uXYb4qG1y2LOGq01nvrGxv
4y/gjdGTGEYLarduWzrVK3TejDEDrqTqdF56mnbejUkorQ7QVenj/11pggA1QQ+F
yJ8ulHkkWElwagz9dXSLB2Uy0wDBPI1LcmDGKgE1AkXQvVa0vystLlmhPF9yrZBR
GrzblxS9FL1Nky/q4JJ8MZ2RyJtTRqWsFvGPvNGMZ+IGyS1cycabm7Evh5G6z2/N
9AzVt8tCUQa/HwcD3Ooj9ZHWXFixu9OBUy7CY3/NLbfEeUdqgnkeO0NawQQf2gcA
9FSdb3mk/LXTbaXjCtOKCottPyOQv4p254UqnUanwNwLP3gt4DB8MLzcpUnt7wJ+
wzrz6WAN6S0uWdemYoTkIFeCLkRHzwvvbDxXnuoiRaAqjVnoI399yONPMYR9qOox
m1pSfeqLNVF4kOGLCJmTjei90vHcV9sk4aVlFX/Nrr3EVxv0IrT/3bDWG+TcGEP4
xpk09919/sX1H2gV9634BdCfPyinPzGp9QnWmLT7C4lPWPQ//a0Slq7qNUPXi6+C
HKKttghCmi0S4agevLemvCpIQmm0iTcafmGGtmBcnCMsAZ5g4x7OoT699TN+mJ6X
XtTdG+S8Rz9Y7h9pe8caTQZWbDOkUeDRp1Hc3fw7LMT8cpl/ntk4RkGYpSJwWykb
ajuJDqYJNVYN8edLvszYgP8H5vVwreiPkimt0SPtdwvG3AN/4H8FPiWOKHJwHxS9
qvFMOp+UAbFP0//oXqj2bntldBzslcp4sIQBZOLmc4/g3MtZ80oDB+La1lHrVf6a
44Y0NQd41H+2nUGmH0GYGiJKGsz7IsaWY9Q8mLq5xQ5ygFcMYUJyiaNcLqE8+sgm
IADutF5DDgK+3xQzQLboUVhnui1CngmfrIPCSfeL3UfPuZpqtC2rBo5np7g4yty4
N8w+itXNhlqio8DquGrXSgCm7GVEs2gM1vr20YpE/eyqKWz8tbwOo8YDW7j1T3kS
IDHbA4PMF4YAiNtixqTYG8Z6cha5m4jx+q1v4UEUebyDTHe8/UXQZ7dx2SY2twOx
pGpUB1pnKzJFNmpTco9FuagFtj1zrcjr2tv7Ygxard4WTjqeKH45ug1nCGFayhbN
NmwxUKrJ7MpEeFYYGmPxW/DbfvHE424qbGaWbjh4ZcGEVPug0iAtPI0HZtA3jXJt
fFsIXQOCKjEdDR8Mn5dLSwZhbxCwzsKEL46Yj/9KGSCRYDr1l4TYHZ42dnH4I3Ww
Cjv8xbe08N24HipVebWuQPRHXk7wzUlizVYOuHw2PVMPrsSD6au5424OwR80F5L7
IKJbK1TLbMe7rwTWu3t0fQWBOU8O85VO1M0wkbAgTfChv2dXiy3tfEwLTAoXsSfl
NogIYjvPIV+DQ37P0uLTcJ1vgilh4OhuMzN9bHWtZwi55UnjejNQutIMSt3C7wYH
Do1ZPskxUTT7NhTuu9vjidmfggh9rO5H49ZGUGLd2jc5D0GSvT+DdjXAssbEzHPe
YVKXkEp4so2H+pH7HvbctBt3WWPtq/qR0DfBNWdzh22b4l60y5r8pwb+XmzQ6M29
Ktteh2r+ZOkLk3Mvhd4UCIUyTg9H5m+uiHZeQlpolxYFP/aH777OaalQPxlkBkck
kjcAPUNR1sdLgW4vvECggDnonKWMaKI1TTabrrMNrFpbXRlRQc86CjydAuX5C0O1
L7T7F2mxZsXY5Sd6eTFQF8XxvYTobJufC2LVyYMzYuKTaF6/lqxzX6zB41J+pGJh
TCIdbpj4I42h/wfHdD5AuF/XcU+ZzzvRUefdF0HOD9ZL3DD9gS5oFBsi4389bBOu
kc5U/bJgGe3q/ZCIu1TGOe5DsEgHZzyW/jNfLm1QkXbZ4tHFpuHC/dyh6eRRHjXY
id4p0N2mlgKYPMC/Bu2jJMNiurGwyvmtZdjUHWaUDFpc1PS+RFneDYQx1oaLDW3Y
coK+eBbiPq47DQ5TryF03SNxBjlbWwja0Mt9DKY3o9BnBaMRbZwyfgk49TcD5ery
kL5Pt9h/iTGsujyaQRSJHs1wg/hxv4B52mH32Fcipld/ibHvdXGdfXPLzpV2iR1b
IvDscHlpnMqEdrmJ66HFa2Hj4WOCKkCpLVVWKVCiYBoV9BYadWV55YzkaH0s0Nux
msqYx9zR3v477kBVShMv8T7m/hmv5YYhfBOHdwNiHhXTSxWlok7SdM2KVeOeZQ/0
Ik9ds7YHDj9RVNqFEpFo1NsfpfVeka/727nZt5d54jadulhC1gwYGNXgqokITftC
++aos9KhfLDb3n4Ze8KrbxLczz4pqQs85FaxpK5x87byX/hFVD+yPPtPeYxSopwj
RbxtqQ8TePxz8Xyb+5aTficQHAIWM+XRdc3VfpGNHRaLibnU3rVAvnnzktbBCdjV
63qkdPpCOiQbAYIB+sLiPN4mg8qgeCey/8GIWxl7BwlsyONq+PUuEd2DVCVEVgZT
VN4kdIK7stynV6Ma34Lr2eQrMLM/KSCQOCD2Wcf63OMzFqFORla2a92XDPg7sq+a
Mq/7TLOUYo25IaWFfS2BGw0xpx+l81pUFWgsEjzlTfbrcHEmCY8KlN3fWmdYgH5v
M5WikrZ8uYtrQlsoJdMe3ZbJUg0Vn0Tnd/JrXnvGWLHomVutqBY6LZRjlo9DIAvR
JanhTy+laubmFyK7MhTwH/9j+oy+2pZtvfrLLAIELw0XlSi5ZStFUhoOUeGNvRz+
dGrQEFVIzMTR6GwUjTJWJ4SONfp5zW4DOXia+yvmE8TmGYNI0bn8zegCyZjRxu+4
udz0UBFvv2XyttR+m17DILeGCJBwzrCavZGmNhACmiiR8o3OaVpEQvz7BVEY8ehZ
seIz7WePzOam3LcuhOY8J5hDjl6k2xWYjJo06GcIVV/2irzyYwJsrFTRGF4+tMdh
8iCPVepV2s5g0SefK/WIkZBqPiSZr8CkikI/m06RbG8lWay6skshXunWaXYRCBqV
DcEyB+EBG7Vw+RgkLRKoHaDK/oPsim67B2HOlVLtw4Y0adoKNzXtwhNEjcrsC6Hz
aqa+HzaYRsSLpF3wf6rMcap3kyIv2Bbh1BP6WDxqkdH5FsGrnBTjOAOW+sA61LOp
olVdhNs6lHvoTOQZogLNsyNdGmICgR8Jb1LrqYBM0qaxXh8mTceDxy5yRTZ/7Wau
jUUaTkXjqzUL6Ecmoh6vTZH7zR3tyQfr0puaodsZkgjUf2gMKs8h+MZaMro7u4ST
4+/BbJYtr7AtXwe64vlIoZUJbImR2JITdI91MUFZ6rjB8jiBCikHyKxisO7enwrJ
YKp9r5i5tT3c2Zr2EDh+ZRF5MuORLSBBV04n0QIg3fs3v8+Uml1H838ZLjO6qLl0
6ng/eqJ9O7/VXR5Wicv1DSqqHZqlTfw7CizvLEkn3aRbhA8OhRKCXtuU/BV2NrrL
fEl7yau7w+pudhdIAjWRpLcUsFHZdYvm5Ig7aGSAsfAvkDKTbckPOgFm3LKUlG6L
IvHO4H/SZS9c9G6ReaTzDQWuJFKC+vSuvN/ZfL1g4nIZiMFO0CQ6pvSj8L65UFjZ
4jTzuvUNF8ahrSJB9KQ36VaA8NzQJFxZD/PXscKm9qGHGqipRTkkH1PNVpkqheue
gVOuwXp4cfGswQqajq+z5SQIop24sMm5KrBiHYMYPgxgQdCf9I61LBG7pIFG2YPR
vvNsSLKUxyM3XhTyXUl9sIp1aNAfK5AWjJMxlt0Pg3qompGv2gfXgkiT2HHs7IE4
CUDslRoFM+IUE4njLax731MV40hUdThHjKM367oGlCJbUFonMQBIWjM0uRoGdsuo
eUSdaOix8JUJYla84uQA30YQrVQ79QpaST5QOv4uMJO2xNmI8uwaVwHpg2l8O5Eq
CnYxZaVlnKUY/9U0J21OyLlyn3+gDGhO1Ifh+G2Sj1Fv6GFZCPunLsfQ3H29ZvH0
IglnQJSNGid4L5X4dNHhs0ZbGTcbvJSBrbPFH3cpElyKBHrdN3aeoGWN4M+rTxrw
zxT1zbh7eaI2VWtBmWvHjg7l349x9nor8G3JCOEPsEAV3IftBNygbJ4TC/U5nb6i
hQJlWnfcKvWn9181ncqjT/h6J7toRI24NM3+tlpDXRKPlQ4KuJMyX0JZcGFb97YD
cnzuHPnK9/+lFbl17TM11weqojFuLq5fObZw9VQ1X6QMd4olGK3ovCK3DkBd31Hb
YHTGTpvND0nMFU5Wst7kyC8V8a9872AuPwoZLJVNfVKyuFJXgfNePXe1/ST3NMPF
P1dDe59PeCNoE1iOffnWcvnJG2QrPHGZWMlOgJ0j6OstkArLFyBgwDUFXzyXU6S6
EqL4EQW0Ngd0j0VbLp77/CDWy7kPGZM2F5MAoolW1dZk+az9oL2QkWxMsi/VFfcS
QeXN3aGnuNlDU/BJx4+kOwvTqalxdZBchywh/cr7R/usyF9Uq8EmqAf4isuUHWwD
Ns3ui2vkq+uR+cI01zmTX7O/jVEdjy+Ag+R1WCwf0+ED0tjAb9PWGh7iXsIEYzkt
5tBuux0AmITI1akbjdDAIduYK6PujrOsTToAsnTHdAL4s9rciTGrRrSGvYrB0cH7
sTprzG2vK77Lz64E2NLIKHzXvz1FIIETi2Cbz3PQqe9/+wyo8WNpGvs5CDWb48cD
92Xqhl4vr/OWCvfVe8pqAb1sB9h5eV24a2JmKrtsYTqlQY5l7I/LkiOwWWMXlkhM
ADW3XOXdUr6ftyprR8+57HmlklIA+lzbHgfDR3Du5LVIoS5hCuax2OMeIENwKvxU
uIfaO2iRNu71hPatnMFmTIYC5y++d7UnDwYEEccnuWR9UrofpSFi2nD9NSuRhZ1X
oVciNWEWcknzBxW27RzZUUiG9fKSyikGjWv81y2ayps8+OmX9sB2facFoDUuK6yO
n3JD36iSk1FpdE85qyfJ8PPZor4CT1k8dD8cvIGvO1xMy0uwSsLStJ2F3ZbTtzLH
xTx+VMoK6+xJITvFvaVoOU0/XvL3m0zkvu7ElpxoZAnBW3VBH3Gxwf7aMIa9rdsr
oXP/Zs8zcYgbPQoBzyhh5X8Nxo43KNJGs3mgeW14Vkn5a+dd9R8fZxcORce3pmVB
lT857SzoLrjvAE+RoRKDHSikvuH4ju5tpVu6CsO8MpRq5MAub1FbYlEQ8TP7LfH/
qOuF+61OMLzGS1TU0Btew6ld71XaSJqJDXHBXNx6A+PUBApzTIiMrKjNnNCwFeim
6pzulzNFU6MDBYIeFyeK+3HmlLz1+dy5Jt5SPVEo1Dg8ANu52dWWCQOowYdp0lSp
SI79OPcYOM5FXFwnkm9wN7VSEPPjmAw18M1XQ1lywMdqXWoLbOv/6FUmG0vKYfDX
j6dGRn0bd1+lYeKoJivfatIzKwEzhaQZ7sswOGBLKYMXjE9IZqRpfJUczBWklB08
8WZj23P9CWB4GKxKh5QR6cIunp5OVjXksWjFk01YpxM2SS7H+4GiPBLg3NZRTHeW
y2Sf+ds9h+wqAZzYk9T6BtB0jTaV++yg4tv10OEWIhO3BZCR8jRWm4cS9gQdC9nK
ZPy06k4VlR85ZOSJN9DNoHj8kHpwQwA3Ibaxd0FmiDRlZnC9ot/STmeza/ggkspr
J+BXz71E2k19+PoB5w0wuWMW1uyqdjzIffklo6nQWOnVJisVU/fv79shnoybkeGg
Eor0bJqPl6kIv+6Oz8bZYCnCuhzSNj4Urttp2GQDXOjEufHOrtFq3zJxPDCUtt4X
epPAenLLNhqErRDhfjZvwbwOKnTNa4FmAxCh4ZZcLl/HvEZjX+f84YSPYMsG0Gbv
5l+JENzf8epWJpfNvpL0BqL4gYV7aqup2jTGMUohNDq5r50NOiSngZWuF8pO/FIR
AwmeMhJMmOZv6fY3hETt23v0fPgnpcWbodIe9zPMbobnbIGQXhvqsfNqStlZSQgs
C1BTeBgi8vyRbLt2vrm8m77WKvkbL8eYjGtF7YbwkIwqS5zRmXeun6Y5ETjgP+8R
Ajqyra8opBTAHN5h0w0ZSAL+xIjZfQr2b/CJimczYDScnw0UO4p/2OniuZenfM/d
kxYf+BbAuHLa2wgEfKtRlphha/RJLy+3TkikgV6zGlziJ3wwH5vRnOppIKlk2xjG
+tfmABD58JY+CJ1NQZ1m2Zw80F9WEGG1paA9IX6Z9wj7Pq8EJBzgZJnjVK36Z6dE
5B9yMBN4k3GyWKJd3sgVavazb8qZgKTBgguAB6u++/soX3+oI8o/XGQE6P/XZn60
Py962J9nzxxkP3y1nwwC7Cbx+WkZvXEezrAe4uVhQMfVL1Mza32tSSN8oSnnumNA
+/TZDBn7wJPufStLiT6vKuITiUIBZsQXkTKRZbUF0RwBSU0WfoWrNsWsVNaYljxD
DaRHorO0iHBirgNhVfULFD9hZgP14ozYlAxb2SmxdVKf2EFRvnJWvv51Rnkp1boZ
oFmgtox0+fjpnUYpX3IOSEgVGnplKaZNQ6hRIQUnuNcjlradrJX6KaDhW/Z8Z92V
tPK+QXN8EpbrEsXsHdUuGRu5F/02uEXLZiY8fWy2jfR9GBS4IVkEwdCd59nEw+HN
d/D7d6SCSilKoVeRqpe/HEieGLgLmZEh5fGm2oi0DS+WW2nb6iCcpXr7DJUFnDDr
fghxOhDashli7RmYm0PtdfJ3ifEcwlwgiIIXGUu6ilUoFhSbdkho7zlYKYdrkA7T
ObqvO6MO492GaWt6+w0z62suMbXWmsxZtY1jNT5ESjsZyh3Z3Y41HR78kyUTQACI
cW+IpqHM23aqFtf3gzyyKyN0j+RezUvmzdcy60faHLABeXta6DeXS59xh+aooA3u
nY3J5zZaVsIiVPjGhYk7QZQcbw6hNIA9+SPIsh8cU8dvamDTYld6ZMX3nPymBw2t
1g4YR3yUVT73MuoWF7iYXEWXoKl9VpBXHi+2H1BmGavx0m9cRomhbwJBr7FYZ2z2
3vmiEhi/JgG4wOR+0N9VpKXLp0V1HJcWE16hdJp/oFCvWVHOhFaNaK27VmdEdwcI
jZDMFd9Xi1voceg2nCx+KPa+h8/1LhIi8joZiwTYmeyp2rLeaGnSz2/u4Tq2oMne
3PKKyxLrXSyvncbwO9kj85thtTvQMr9a51yc6QXySKks6RNikDXoa2kZnRxIAdIp
k/cGnZ9NtJnmjQZMaVlMvyaEo7R7SgauQ7G8DXOJmtVSttbKxDoQPTj2feXZtZTW
zBszPulISdiurNX6d0KgHuLKJhrX50q57aWrIGnPGeTIy2KD+S7pNsG6BsBrXSIw
mh4DqXfsqOQqCczsAZhG1AdPAFsXSfwfdYmhZ6rMLpo0eS8NrJdJxbO7Po9/0PPV
+47Tp9tLjeQWoCjzEZhLASwd9PiyvWiQUqeUfpDAFSGnMY5Rt1DvfU0k5By8h93q
VJsKiPauJZD9aRyyCvoGyJFtaIqmLweVVarNDLMHwkmoIhn2MNnf4waYbiBgMn81
/rZF/20sQ+BhjIOOtZ6xKUT7TkAixjneiXlhDt5t+YG5wRvxe+XW65Tu0drSH4zo
cThqWWsmfwDjPtPoMkwkLbgXE6UfIMAhLXzIJhC/wKqxMfrxZupRlwEnlQAUGFti
rpazpZYwZHkzZA5FeOhNsoP4uzQQyDLC7xCjepnyBsyE9FxWjUZa/OXGH0HXRXJv
rVqgSr6AdE/oNR8d5v/1/cDBK0Rlp+OPc6STqfR+BeZ3oTkx+jw63YcVMGkpND5y
nrqu7dklNyJJfPBufqDsst7vaUR45Kd5f+pJioWztGiFueqqZxAIAg8dC14Moi39
rXpGgroyeiDlbDljm5Ra96rsBJXx2ABy2IM+mB06weNPmYJ2QSgczJI95s769LGb
VxoDhaEGqUhFUNGYadTHQLS2XqsxzftEvDIn/btVLOZuDAppqGQ0mUSl1AbTXkkT
LDZAEJR0bTebWkos5LSlVqBrBCiD2TJXae6x3vtWOWXVfGVt6Msu9VkatAmA/ZoT
eSQdA8aWG+QLC+YTJjZHMsnOAJWIfij1aLYzfq2VtBDnLB41VFLw4+BTiK1Xg3xT
VCYu1c0bjqulHB0d1DvZlQv0+JXQqIZW/+lA7bn9N54k9Lf9IDQqh3+iHqevsV2H
z5EVL4lM9Q0uJ0uHsd7FL8qdXiimV1tSV0UrU3EM1l8oKev8XcxNu0bYQCRfE8lq
2a7MXbn3oNBCV3lW0vz+tx8OdnpGN1wau4OCEpjoUArqxcsZOfqwDAaDPTq5/fOK
qLBT1/n1AE7R9wlLHv9uGydQ/Zbi+e6XTZL2m6d8/4a6u/h+0pQLHLoc8tI5cmlW
/ndxYQrQ9TibyxKjkYAPbCAq/gib9HiRzIB73yza3GWBv+4FCKqIFhZ7GW24BiUM
2axyf8NPt3KpvVt1ngGwWctLFosp9AZGz8YkNizq1BmPZTtQFCOBh4z7yZVosbz2
bwZEldHSI1HzzlKEP2jaUbk/edPsTf//beu5RTHQi39EK41k5O5tBwSB5Azv1THB
Tdtx6MICbtt1ikeNge/6prlQVQTipYmVEoBSBc5ShJYRYHdZnclC/nu3qZ8hvNx3
Dp1sS0xFKGkkdeeYZ10qa5eYq5lPn1NcBGugCO0m5eLBzBIV9BUu6EyY5e5dxqSR
dIckCUxX1oYiWRGfFw83rTJnDfWsp3tXnG9OmsClPZRLewa/wsEhdlBY3TlLBROt
w0PmUTEX+L4LoKk9S62vykTnZgId+FiVZ6jNmm/6sxLmU1M07EulCddn/bUDdqoH
fmQypCWaLCaEBijnaU84gNdophSlnX0G+72CZqHxd9AAk2WK9pkM1/Q2ncTo4Ko7
Ol2YkuKIfUw7xK3yYCgm6J0KVUxKlwot1c9ZUMbse1jZ9fQPm0PbwT+XDsKZhuFC
ZNGiFh9sMZIU94+2Z5lxZk/OTlpuJyfbcJgYT7yPaGTFPvPUp2xazWiQygXoPon5
UpoHbI9TlzOUxxz8l9kftTLdg1/wh2pctIgN3OzwtKNKEvS+gGfsO/RkqGUsVu8J
C0Xpebs83ScgS0ogcR900DJiEFb6luP5fl4BrBvOXxUO3w3LGSULj0YwKjz7D63I
2IiiahgpkewMS1/Gf7upcXEl5ASXedLo6iJZGMgOB27uRU3F4FkibTKnodec4/aE
3X1HXNf7G8Y8lKfuw+FyJWRGADS5TTewCdZ3qIzkgI9U002VGvOV4UhEFfE4LQqe
3x0+cjh37Kwz87q49OObAa72JZvMSmgX/uwHdR+UiqyFiZ6UsYYnrJrhowPGq/EQ
7tPcLpZVa0aarkm4B7Nt0e0u6JsuLQawPO+Spc7tJE0yWmrpJJX5u1OPWh6eW0+Y
rj2LUgXVuBDfHxUZzjeyL3XY8qge9ajOOiHqwepZHfGGzAHaF1BGMtpedPeTAwLw
wyynui4cY5KvG1dDZqFwzMMIY6c/rmgY5z6tdfeWFBtsvAUEBzTuUX3QNSbgJpH5
luvrMgE7u1SRtIFJRbubMprDZ12rCq8E4CfmP1tHLGnAor6q7mkWO9zWuiX2RvLM
UDaECm9d+rzI6MUSQ3XQuOgxXEx9+fLjCXlLRNWpJFLYVW/jSQBeGR9bdVVZfmAQ
INDyzPfrbgooJCpzBPFJlmE+cbUOyRl8LmMw3gZl/Dz7ctOh9YrnFk2bSmSKWKm4
D8niiJvp/hMH7hTrpwZj2WGC8JVtqEZjHDp5RJzt1s8BAdyr1qfXmeEJ8CSrsPxE
zGNYHF2kjueayRul4tLxTqaGZ466WX4HSmP5RCiVxoBHkW023C4cLB7Z1+Dvq1wJ
AduF0Dq7OGmSxDl2SdEQ7ZZYXEAHNZbqxWg3NEchH3c2sVjAgCYH70YBMbUSSgRg
o9YUb7pe/rCBBwJGLI9NQIhyz5JtQUl9kSrDnrMhHcy1JiMmKZ+OQNu5EiPhWv+i
HuV6vQn12X2qyHnIDrBvdE4yAlzfqyCI+AjrqsjdLmKWk/EdwNlufoyY2tkyf/0a
E/TsHKTqt2TsruU6K1msba/AA1ah8PDhmixLS0o/tQiNwpfDgxAsyQO/cD/gvcjb
2JMt8Gx1RbsLq1t+K2hHmUqEU850pThSSqr1vDlhM66FTyM8fTcFqHj4tM0z183/
IBYtxD+c/LU5XL9iE5zohsnFhrw4xEcCfc9lOAdCC2nC8LSwcH0KTB+wLqHxoxMA
DY6FEjMZP94Lg+NFZqroUKpiNNYA+mjPu967qNOFeBryMqzgb3wopf3OiCRCHVvL
liNHl6FjhdbzvzeU/KklzSVuuJO2BtZZ3OtGYAvpA84HDQKJ3AKaujdDoCyTH17f
f9MHClEwqug3QPKwvqnJon9DAU4ktYJgodVJaS48K+SWJdgCJdQbywtg2P7SE2Hv
pHOaHrojxzn5T6WtmjPLeRO/MwwCCjbBOHmdI6bynIsQCDfix255Jp7ruGHrDJ8s
fptCdDBkzuo+agaYcALCxHSfNqATWsb7BDkSnNevmSDI+Zn3Zo4LO+s8ER/3sxgm
6zSaOQ1/th+jhLUi38u50dqvjQlpvcPBpxFXRQuxBxu9LgN2b5/PNN+YSOICqqlE
YGcDMiKWx944J1JAXcjihIi5waDpaDVmT+suQeB7B2RgfM+QAo0qXwU1w8jICdDJ
WVu4Qi/Ocx9OyOKGKOOadkNVVhKUt+qedIxnZbR4isVuUR1W065T2E1hrBm8y7Al
v3b8Jn4V/SbeNQNQ01QP8fvWN0yT9nsInW7xr9AIXf/UdmfPdjWJMXeXgIaN0KJg
tuf4swbKDvn/LrzX/k1OkLPcdFiA5zjWuB1f3Uq5+AX0p0nVRPwTYqHyj4ZsZacj
gfcjuqiGcu1dMvPllO7Xjt6pyR3Jn4Iv32dxH6OB59R1IGkQ86bRNmIrL+UzZTm/
JFiWnfdlAlXU3ImtUDk6iQZfdbb8YDJIl2VswynP8H4gk+jQtYBQyG/b9akXGwOG
i1iSsl5x/z7YLs1yMip4fBP8w2xTXR8moXjdauUQRqYTBgxJS9s12lT8jYPrgtOd
iNq2Xfjol4iV+w2rU80zt5jsUHNw0vIQjXKvafFeFbLG6q7pZygkHEnqU635yjmU
BUjhQjC/iBoiuC+HzGe+i4IOiVu/3j6aak7Ngf/1j4czej5jXBlUzcaL+gFaGEvJ
dGc5IYj3U3Zz+MpRsW3v4Sqk/WEfBOsHt0GVMej0bVM30x80uhf4EH8NaxXOw0wl
ylXA7MacK/rQiEtEFrch23Iieq9C2iemDUcgSk+rSNXnTphOzG8HUuZaYzfVo6+2
svFvXHJ5p6Akjj/cbCWG4OfwTSa6LmDBJC7SHOsEsQPIW5G1DPClO0NRT0Wo6x0R
NHXzBEnIkjY787mX1Mitl4I/my43jD0uz3qD3845a5+VH6kRixPjI9Mu0Mc62Kws
jxbRAEbfj0zjbeGMVUmfyKdo2q5BJc8HV+wSSP2zSXVyEUVHsRgEqeDSJw9ZsGGj
YxWa1ULEPixI2YxHPZbwIbNw+DIsDHIQyOyk/tXr0sMf4U+y3TaMtWdN+tDshjW2
/w25F1RHftrpZ3RRInoClUvQdYXX4xkxyxbpLY6ELl+Fyco1Gr93mJrpqp4VWBRE
kv6pGrxfK5SGodirDe2qzSBpFCMExjE0O7IvNQZqaNzba2Bm4eryux8bYsnfNkQ0
KjfjJoo+NvcNIEQgfXdLqmqsj9z5n6g+LPba5zenDxuyC8gRRtw9XCVQ+4AfxZjG
rpDQdrb8myScnaKJm569y6Sk3KgcFCEWCadcCnvZgLGTqZ1kmZpEPfVJabz8xhkM
GdG+B0OPIy1uzfQ5H1Rjel5c0dYL0JOsZDF5Z7SqebgkBsDtkr8/leHxJrYZRvOK
NYYCo8pv+e3qGlyyFh9MEOMs8omYTsegQVJxfFrviTrBeNgEzxJhD+S8llcAh7yh
CMool/EW5I5LNVZVnjqJGvyE6uJruTSSY/ESC+x9JHnLDoe+9ioKQYWcBkW3QWY9
9oKETgfJ2aGhkEh+LmQvsmuYiffFfLLXmtCfqrylXrFD5rI3A1GuRgfI9ruT6OgE
iifyYlgkl51/c8dbTcN53eAIv8KtrgmFC/tq8odlilyvMNwI2LlGTgZvLg2eWDRv
B3yxgwV39kHAn0IuZ6SBOlFDU46e5g7kI58C2YTAfqlZH4vVdolnsFTnbYVNBSqB
9RkmwpcV1DQK6fDhqMIRo/DMJdCNgXP4B1u/Z4rqVZpZzqGhhGxViepo9pYAhFwP
drU77Ctocmhc7rVms/YXeV7Ofh2eVumeSNjq5PTyCbXhNpz+pVGvK+EbRaAlLfax
D56BFfBU/uYIfO+p2IcNU/GV+WiuptAOWattx6TzD4DtjfrXsHvTKNhKL/eXxmzs
W9/v0FkjJWHqCTx8xathzYDP/1V9Emr1Uwis35e8pLCDZYGEM1fgx/PRPfU05of0
fRzOfZsIjB11Be5H1tkccdf8sFbJ9BPec+M8G8vkPNXuFGFTvmu+l0wB4Ab0Z5AW
yy7046lq+GhO7TEvTHi/xjEusLSf1eeRnMdCGrMsuiEZhSyXOnxO7TpQc8/pQqeh
ybmfu0nhR1haH/QJe8lLXDpiPTLTeHMikFivbCwwQ/yxQ92E/E2g+i56ld5cOB5j
sULP9ERAghc+qdwQSLuK2/P1P5KA72NkFLNEp8cbCSWjJ1ecQ0iyemQlTG6WUgbO
2kdG/vu9TycjtqAMZbnFA63PsVTSAOiq4XxDNIGoL4nYcwVvuWISAU6+K6jHeCeK
J9Nip69MYtRoysOy3IzymePrKHXD78qx8Dj9a1QPMQnzYGWiaAU8TUxk0ULgr3tW
sh6vxTZB7OSGEiUmNMDorbol4wwr35jspD+x0kLkqYc2LCf0fVGu6BUvwk5fuFby
31UzcpxUnvtMTfl1C8EUNbwgaB3yey69/03Mcr9tmfEwriT4tPqlkFXdpAhmdKDQ
5Bxj1Rz9Tkab9uzCNXcZ+zJe4Defe6L3oCmjb0E8lijNfPeHVOYI4pIAOr/n13H3
guw6caJxzCDINBd3R2s4c93FKCdpEff8dOVq3vaUhITiACCtv+9IjOe9hFQeTvr5
guSG4xap+YMGu4cBCYHlRY4i63ZzPOEU+s/zZ9HftKA3kj+2I/y5DpWhyPh79k8z
cPXd56gC4L1SOSAfzyujbx0kXya6WTyCPB/zE/g3oZMcGTKmTH5Pe+zyU30Tf4tW
PNkzhiN+9RqivRZNZXvX5blMYl4k0IxuiBEBA9zRebYCOLYGOXzYcyBYxkCiO5PV
p6vpG+DiMJsizRkrECqW0cuLqUodFmRD78IZm+Uz7hS/5kT/ms65lp+5TP3dWjTo
wI5q6mt3tfLPZeRRwRIxTRqHIDpelLGLXeWdc2OxEB+q9kANPO8TJdx9CHSTdsdc
CcnbQh/U87I+SfqW6nCpF1ZEQD8X1C2RVWvj71AvLQO+0uH+DbcM6WNBvGrhVsdM
mdR6u9vtrVwIQyadV2/UGdhru/EcDNOViG0FtArk/n23H3prRcbRWn6WKjPLeqep
zFP1Ud9+qgJ5bbHKdN3atTnE/WZmJFPv2zB+Oku45X5Ev6wr491eL/a59UAv7Dep
y7/HGKZHSn2TlhkqEedNg7AUP2Lmn0wAJNty6xs6M0SjN8d8uhT3fU89Qr3+4bEI
AgZt0V4KgpZuBRmhW+wbuWFy/rrSQC1Gi4a5GREPW+JhtZirCqPyD6bd93UAPSh5
OT47bIeBsHyQK8wr9/o16AE5MsKHvffAPN2VurJzq43iqynpri6YIaly7XgVZo5g
5rPwLtpIyGrAkzkg1oIy1ZPOpKoo04pAoOAhWC1WsZ3rkLF91TMGEWpi2Cw1y/ff
kCttIkFaNY+16RiG9f4hFauF8CGw72iwqg9ekXFZ3KJmTyikAV0tJ2FOG8pnFQDb
kAWw0pU+itLJ42NaCXrzefQD5DxVe2zkUuBefGAMvHFsCoQKDuL66TYkKf2UrVId
ARhi5Ce6fDfjCCe5OUL5dt+KFOps7yBJolCZXI4uXMhgZNR5Z/rmX1fXPUInhOHK
GVOqia57rolypg9++tE+UQ5ACUUN9gm/gsDpsPe1RCdOOsQxexnCvV0fRgsIesFq
Tik6jYkxGIPuJRO8pvu83hisCfaZTLX6TulD8M8NT/AShGKfpf3dVUxfD36Hj4WV
WGIKx5hGOEPGssTYqhneEpCXid+Kv9U/7Ff0Kw/Nj0luv1pIVgqNwWR10E+KOQ+I
TnfPassSiH99MTaoW1f4aS2RyfYVrkbUp28eSULyyO2czjU8ZXK+35ilMPlQrXJd
hBggcFqGT81QWaV6w9wFu8TIlojV8E3qHJRHUdPBIKpfLg/YIBzIEM1X9cMuoGGb
ATpSb5pC6OH4smzC7NjJQOReIlTEj50Bmik7mzPAi00p6HcoHv+AaRrWOEljKX3W
nCZQQUOWu3nR/h+rikBxOwWl790WF/dUl7JW/Dj5/LLcTiV2lrhjJEryINlYu82d
9It8843LLb9HXBLboESSttE69D+ehjxVRUBspaj0q2TpMQA16pqGeEdMwrW0TpeJ
VBTBbkiFzEXnnw1KY+LU7agGP1ut4xDFen3/PgHqoHItlrJbXY+9VLqVEDo0bl6m
03VRvGjxyHZYQVB/nEHUjtoWf8Ug3AUYFJTNIbatLG8lAs4ZS/ZZs/6AyiVc18Jd
oCn2wz1KUGiqZCRbw0dDAkVqeq20mIKD/wqggVVqaYtrdZhHtBLMhCzGEQV3b7fX
m4kVBr9ESf59jlIIWWRE7r74609Rlj5KD7c5I8QH8RwrGzpfwV41/BAVT4tzo2QN
J3x/J97OswvExNAS3gryXBo3jtnzYZKZrwh+wZsXT0tGzO4XF75qMq9zFqSYs9dD
exQkUCMVGu9TMiOOLO6xipXYDn58MU7kC9KyslxCMDBh0BvJdoAnzxZdSE9tM5NH
nl1wCW/wCYqjar5PMM5/0+fDJf+2I1Kse4TEpyvy5PYUehbm9uS8TNE89shJjInO
6DwdDhgvksnO/ZCkqzmqsZc8XAe+guvc/ptvr2HRFEfHCJjPvIegbP7HhRY94PmI
If+vZqhoE3uwmFGyHBG7WJV2yCAuXO8U8VoG0e+6dksNE83UggLJJGW26BVBXlnz
H7VNwouIoGpK8Uz47HwCn93oYlhWmDNUUybIGr2jWxmAb+ezC8EsIGsxg61laYQD
2bxABT8P+zObrOy/lJTHMXb3CpNyqhOv+tS9d5fe85ognDB5bI7mlTEHckeHDPPn
+Pg3NMuZ/kcC3VTV10mTcDL2y7l1eAtDwolcr75cbr0GTMuyFXAAGXqaXP/1MnIt
vQQ/yagzA11UKMtEwHmpN/oY/nq9c8e9PFSSBnCXoJ4BKDo7+rPK9TohmpB+gDWj
FBDCDQ746A/8FozjrMnrZT3AvHimK9xUfX11O4HZqa+3qrw/2Pq+w2tu0mgJD6Py
14/EpC7a1ef3I7vSw2SWhx5pXdRW+a8F7Gb2apJjFIPZgngYq2xrl5krSSd0g/HM
3FSrUY7+YbhiI7ymvCJnYPhgtKhf6N1hojrX2s8V3XWXoURgjuyZDrzbs1OtcPWp
4+gj6owW/LWfg5v7rFKLADBOyVp17EdR7GLkXDbj6mhFuRt6wTXowECF9h3fjtOF
cizZcnxzXzFtDlk7s35VDPx7FWK4AyHtJbq4dPDXlutjHGnPkziXWmSdZgL5cqR8
B8/45dgQET1XwccklcSr7qR93qHuBafvKx+W8RZea75DRV9TuTvdfpjJsTQQ8qOF
0eo520zDIsSF/imSBldP3151OWb2e4uJTcg3zzcI6blu6BTJZpBsAyZals77g4o9
bJmLWXzzObxEim3H1BanL7TkHvS+KvayrRHqQbWsQyxlrHAOxObhJ6f2FvbpnsNK
xzkCP0e6tuV8n9rXwBNuvISQBB8OYTpB7W9g8Ws89t5lJENUcO4mPdGybs0L3k+w
o8B5vxcKa844S9FJtWpjUMYf90ZjIhIY0j7iNYsomh+eI13biSoJIJkVbvdlZZrR
xjeh1fBrGiLU2QRas31nNy65i2iag3/fsgWvL6fhWK6J6XlnaBk4D90Dt1xt4N1P
dBcK9qe3loQ8d6ZKdRNff9vkFUIGSWo8WLGiD+RwDOFssCTubTQYGoU5kpKGFtkW
eubgAgqYhh5FNKGV0VMIL6O433XIoO8Dd1G22lVnpJKyf7MyG9cyMNaeM2n7GE6y
KBYohy6jq8byd4evvr41VkTYREZpSxKJFUvgxvmP7ihzP9BvHQ/A/ZVhd7bAFKZb
dr5GKuMjQ484+MT2EBkFWojy79yUa+HppVciN6P/DbiuBwvdV1NDGFQaVQ4VJJ74
51V4f5dffEWDGK86rXAm3icDBtnEy5I0yTwtMELzxVyd05m2E+pgTlN7CvAR4ORo
POI+SJKFhxIVT7BxJMKXL8D82ZZVxQ+0o5BWWJIG7KPuZVIr4EU1aA8XGj3J3QM2
VJiGsL8tYhgij2eAKFrJvcus5r7BPXJ0wps7rbXOWuXB/O8tZyvKHFhM62ymCBNg
9mRoFDJK1QBVAyqGIY6UEZbkUqNpLIPo9X6DMdo4lhPEmOW3B6aAYVevTfDcaBl4
4femoFCuVifVWCyE+MDJDWI2PuEeLtPmnsNu1gt9HTMw721adwUwYv95b88cqbVk
sUes8VrqDiN3eNiQnFvFhxsDdo5nGnlkr6kItI6zeJtm/UqKo82F2TiFzcQYHmf5
nkYgUHp+CDzANlZVp93lJIysyfifNbgsN2h5i3PANZFcpl/39eAhSUSQ+wloSZmj
AN/my+D5DIMtpcG7K2c1Pf/RpmUO32xe2r7ftSnK94EwXstwnvZu0BWpKVwIzM93
aAKWtocKBMKa+J6zMgtRY2HjVdaDt18ZBx+rnkDPElfSqfOj8tOVRlsW0DF6pzCG
TTcTvgQQvs31NcW1it5BGOGNlRHBHar6hQWKO4nPatdIfL0hcpSOKUycKibuDVh+
A5EGlwk5XG0/9baRHJ/TvfoNpYDkznJybVSpsog/7jmwyvO8w9lrvNJ8ZlvmpuHQ
Kml8Bd2Hr1JRmBfLyDAMhjXEXiLTaqGw0f+AjfyvRNltAxxFwAfFTto4qOOI/Gw4
5LFhis/GZ9PIXEKtPxsRZ9rIyx7C/rm1R7/A55re1aMFQpESRQO0BAkuISUYigwT
tWhkWY8oVts6kw2qmIaFRSYmlAr2EdjplnsuixVNz82bEXANUIu81yLOEgCyd0LW
3ALHJnA/Jt8Nvz+bDB5BYEGTJKSY8tfnltODSQ83l34eUfrLXH1AN/Wx0Cql+qwZ
7L0YufBJbYbPfrL23hR5gkdDQSfs1QiVGetaJvrL7BoZAae2hNfzl7i9/ujUFkQk
j/Y2wa7bFVtK7+LaJnE+VHU85NQBapFaBAwo+DD41vHZ7AgRZYB5ajRTZzkKzyep
7k7Upqz1jmBZGdRsTqFjuuuYYbUsk+kIAH8kC2pG3axje0KfdrPNP6MXY5WrBLem
20uC4XfNMw7zrmOPt+nP/uQzBmiPsq8jTzIftfoGT0EeiSMsQRuaYK5gksd6maU0
CFPP6p81YLZVjFMyXL6UJImYBULVKCYfzhxMSDsObL345lIMPhT3Xe2wZUHVEhzD
shD3j8tG6QTLP89H7RvxcqS0Tr+q2C5Ls04ztcDBT48+xZXutJOuG6JjNzv1BAFA
OWGBUoiFEEYkGqHHfAbaNNcIFoUGhoGBQqBzKN/EV+R1EEW1+Kac1flQxxoPNy6r
xJzLNK8J2t18WxGESrBMTotHNUAK584jXKdPcvFBvZzPqU/hfSB90OGHgz9p38/r
oCDIm2rQt4sUpH4ZNBqVTB3SKwcDRHBddcH2G2daipy9kTbiNUAG9J28K/aCVVif
+sGQq389Tg+nKyiA/INoQCSWYAJa04whqi66cX9UpaAoUrEqBi0kanoGPYKnpRr9
S2l3zfdtIKYNwBeDJRX0NQ+eQ0VszVQIdBMTyD7gCIbWjdN5P/5l+Wneg7yOZflE
QUEJCkSQiBB1symp6UORWVIC8Mpnd1lpxYPnYk6dMwk+BV2VhztTjeZxdNqYmrGF
+bmfLOu6Ly9Za09Zg4jLGSuL50yP4dFIWefUG+jqCNSVpbPWoIVbwWYaQx4jFNjc
FZGWJTzr1lRgflLcwxxas5SF6rCTK8M+ySt87mO2k0PNAdeSVSDv0LgzkMsaWA6u
+pgq68QzXF5IpeXuADieDcnB4A+XROlAetdNpGG7XvDkWuwGsa2QLyw7yMULAujE
YrvjtKgEp6qRMEqbkWOWMHn1vbye2z5As0BNolXwKwA6E9sKf5W6dqCWcmF8apPt
UViXgTAeWVtqz0NTsU4fWjg4ApqDA5x/TRWVzklO3GI69SrKXtb1OF0WGYX1SB1J
rJilwdnxWiWDegP5C5UK8UPy1I6A2f8kOecQtSPhI03r79Svr9v7vT8fdUaSR0zs
rffvje9gc6A4kU03P8519KsnMngnv+fcQklifSQiA3LvfDnPkB22LbbeCk9QY4gp
eyxscSlIQtAWq3/sVTo5uzQAzIGJ62gVqr6Ge2CHKtEQfV/dfgYgyxDF1kflGudC
4rcj+MPYDGjMuaw0yePZg1x+moxTam+xjNLnXyQZum9Iyx0YRDwLynKUO1eyIG/E
2N1gZMifePN1h/mljiUs7IIkePF8amLnfdsoKPyMRtuQoqyaQJlAIGzdwwYH/OX7
D7/AIHRsjuyXlVYyUEl6kGdsU1Oy5ffJru76/3keCjSve13ILC1pw2iqnjWGQDBL
PD1ip1JyCcsuPaJcCXY2R4GDXiCiShOB2FZhKxfOodbpcs4mVvhMNTKArYffFM4b
/Q/GU19wXC/4Gc+S2WcvZZE3IDVeKU1+/5oeFBwCyiv8PBNChelzjVX5jt0S5koP
X0svZ5rY6g1UUfm0279loMJnj5Lb1aUYcAJ2+lFnbExeKoskq4d6JISNYWrAKAf0
mWCc9j6zaYG9yL8g1ntKdZtG7TXf9WG2tFST11/B28RmFaOsWoOZIBikdMSc5Q+G
3Vme/OXhaAJfblLyL2d0ceqDNTi8tcP2uZB6sSdB8/udvEuCXw/lOMkET7PbqCUk
GAmJ0/489aQD6lUz0WAHe8Diki7pHHIkvMojXuzMNFLQzXk+l1dLhplTDsIiMgev
Sg3WDZTKPfmbDfwTTkRVb+paC8jKa/VpUhgBVvCXEUyzjJBJYi9f04V58t7yEgHN
7fE1/PMEBTXxL3BbEXPnhy8ohf++h+SaorOazTYrhIzJQzhANIkx0ljRUVom5zuC
SeZ9mAH8ZJpBPzttrQGZ3t0mnpU4fGW477F93xt5aFqB9FYc0//wjGy8alJEs28H
CLPKUy7f4ibObV4e3O+X/82gQYm8Cm7pBpKwWOu1l6qtqUG0fHLiKs9ZQLmOGFbz
U9EOpK/zalgoeNJSfVq30i3zJsk/WYELZgrI6nN1g4mUgIdhT1B73spIV2kWBv4M
Zf6Qb48LSc9de6G1vtVD/LSgPudJ6D/IbRcvh4+bASZpwla6MRmsIOHpLxAw8gcx
6xmur1cxxAqLvkDUJOmLRFJnGfYO9y/G1QAmOYhQil85qwTuzBP2H/Y7P/TOPvzd
St+wmIfvIKD2oAfUQK6x9L/rLP9dakrMJdOZ/GJMlIhjGb8ewYWJFk7rZjMTEdqu
DO3F9mZJ3BPX8byFOB44GRAwTwWzIB4lj3WI3dvWDPhxLOSYp6FYT0ZkGJNTkRK+
B4AZUeqzQ9XhWkiG3lY3a/eDnoYMtwnFbPBNwDbtDVu76PZtv7yt0+CswVlW/75U
+Oc55VQYRffPwUKpxLHqYNsyKMfzmJ0tycszKQFQLJ3cNoanAAIMXkWghnbzaw9m
0yhxYS45q59Mph0AZDVdDGV7+2y/jdvG8b4AMyem1KgLD7zu84n2iXqx+a/V48LQ
/V5YCZTK7IVuIfD9W0vJZhkbu+OCVJ4lFrpK64hBz1rf7+FcHqLJW50K1zyAgfKC
F7rBKpdRu57KUtQsCWq74tgCQyZ3IV5KSKXeLe2jbFhochGFaQc7XioGOLk17ZXd
ffPYBJObG+hmsraoQC+gI7u6h8yZzQ+wICTzWOfIAKDqnmeJzbiHpg6OkAzeCgKE
rwec/a0pebNpTG1HFS7cj3hbhLQfgp1KbFfWaf1AGVNAbU6scnbLlnzFeg84HKT9
VUxLgT1XCZRHPhl07++dvbdhK21myUeznTwdwUYsnCeY01/jtzZNKcEsAZj50zfR
WiiBQP7VtEaM2vqCWYtPnqcUU1dWE/hrCs3ihdi6OFBxLfibxgwQCdMBfbGGb4T6
bVH/BiotRQetmt4TDEFyUd+IOZAgpiVzsAvmvzU5ITHBW8Q1NnKxsqfcisorB5+f
5YPHI4oYqKQmo3HlygxPcLM9D7u9xFJC2yfzKU2B0ZZSNkXpCt6pX2L165C02o2s
JHI8ehXirYvwWrmL/c9sinKMUSc/33Mzbh8ilGXn6FX1q0GurpGuUZuG4wAwr718
XU04AMofWamgs3Rf44kYFHAs1741NvGK7rPyGTSMJ5QVoxdXgAfq2+6ROr99btgA
a3U+7HfVzsQ8VNAKChBuvwNlUwvZ5rtc/wTAuLcUqybevhaHjJI0Kxxj5R2PtHPS
o6CDLj95EHFTOrQ1FYH1El71XHDpJ74MbIj2aTJuBTuPTi3xs6EhwOQUc8n9D1NJ
KefENpDHGtnjdIkG/jkeIeqPJ5z1X+8lkHDuEYl1WgX+eTgW9/zQkkWG5kepkPHB
MMiz1M6z2ekN/NskpbgicHQzLN/IuQoBhU/gcfqbSMGhNVIvXzdM8jfDFKoWbIj1
jCbwidzcB8oYUvHx8GqyvECgU84uT7f3dn/j4T7lDBK3JPUWHgfVPFnCt87Bt8Cm
eKQbbBrBsFHVGT50nRr91WAH+LjYCxVycRUtMwVI+awsHV0sMqGnIY86qrgKWvGt
18YFxadT6YM11ilEAWz5I9H8N7AkxFemAGuuHGImBs4ZNX2qogAikA+DpWKzpCte
MZBLHMzFFnFc5HsTxO0/RGT62yeeXneUKM79R8++CuiJaLE3Kq/zz85exZPT35Me
KeRg5HLUA8XwG1/zWOKgoTuuFpboDmnp8bbIqCIwbFRwQX54i52s/OTFBqFS2iLy
FppWGMgG+93u86mH45iOgdDdEpopjX4t3azsm1iPRN5z8/3X3GNJ8l9pqQdNTga3
+XXyvZKiSYTkQVL1Xss/q3Zp77Fv4lwknimgCoNxqW6oj+92pq771e1+2SgRcJ7j
sQ7HJ7P/N35lwkRRgM4LNegZM0S+d+QcDFZJ3eTIFc65gsHV3huJ3DHiB022QU0J
Pj4x6AxxCmtfZ/d8jHghWx8gU9mHi74UyuC8CU7WWk7eso5pMR11w3zTyxQpRJth
hSRiCcGR2dfCuXCbXPEfjLS6Ck3yQJe+oDsoteVvTVD9IGDF1UrP1DfzI5VND8Ml
GOBYD6W8YHSLVU7bFXLuCq96x30XWqPtlOqa+cdg422LM1j40wIbsCykDqpi4gmK
707cnPruejcmyY79oRe+p1ANbofxSRFm6coJr8YA6GOo2gwnv0Ez4FRqxvpjoddB
UUuLNDUlaesozMfVG/J8zWtqrVqzS2gny9UOgMgyluYVXSwMy2PpA3htep8/CTtn
+ApmKxO2OmS7kOtL5PgrVW7ILU2YwotoMHIWfoulPyQjS7ukrEippeRoHinwmD59
4aywYe6XlqCqZhehbfwVZ/3EhDTfS5GldDlBkYEI7YrlOVBPk6CsfmFPGCMpsyzv
Y0nHXVTVc9rQ+rYkl92GarzSsq9NKsSFBvZ1jxSCvKLeVkk9Uh3ZeEfYbFSxkBjJ
6qRIFBUDVkBtqo+x+W2UVZWfAHaR6N7IMvgCATZbl5otNNpmVY9ioqqmMMPxxlUO
dDTeiX+gM+eodWtrnxBOk/brkkB1gdBQcit5SjsZO7NFK78Xi6V7ZVx3seroRQPL
xFvHwLB6vm0tpyS/DAussTl7TBPk4mZ2jjkS+lTZTmjsqEQjpM3mNc5le0O93UR1
0glFWb17B4i0AGj9DmARLS1nPiVsvCoOcGJRO6yoBfp35/hgTJVLL65FzcfjuGz1
DrwbosiuaWqPECPcZktRfdOgi4FiXV6sooI20Xt8GYbf76W7TTUpOUgVKnhrfUdS
qaZFY3pwv/KzHMwhIq+kxj/K/MMkbxKiSeB3OLoVu1FjBNmo0zkg+0gT1l/Jpfmw
C+zIlsbr07Ba5hT7EfrNWm+iZsk8C7eDwYlKnHjr79c3BeZ8iI6fGnBdVyrlEyWi
Ev5CTpmsGcbnsFqkTP49R07uziYN1hZFD9S3Pxisa6VdLlJvJJvhOZfs4HizZopW
q38RgxoBw2s8R2iM0JBQ8u//XBQldY8Bqy7vZk35BfKw+ab0rEVgY/SRh4CpI1Lf
IJDVm1nc3mAgkZP9gj/xZrT1G/QZXPF6qrKPTPrmi8qAdAf78C0ip+wufD3FmP1w
thqTZY1ABFkvGDE0EjIhRPT3MR1/xGvQyljLqoFok/h/k9W26o9KuOwTF+tgKftM
VH4rQ8OnhcJPUuzoMHFPcIVTkQKHmOhTWGpBZdjxsfcMOY6Iu9buaIHsmPirhCIv
G+3MpP8fYhE9hSHpcZZQQ84qC3JJ5dIRMHYnaonLANWhau759li7ch0ki6VO1CGB
PB9xyWyrr1l94tHsUOGRpzZk15M71sQweWG/0im8SiHYryZ0hXq9MrmTQOCMeFC+
fZjI8WFz5VAhbXrbpAFwHoZEvgVfJVgctiv1A38xlqFYBvvecbBbxs5l1c3cFdGM
CM0IDSaSQuDczqCzjj99Gcq32C1MXS0wRzX+8gK6mUJO6fqpQDMvZExIAV4xCctd
87m70/vk678svktyZz6Ch3K1UB8d5DolqTSLppTNPWdhy799c2DP5D7RuSAbV5f2
IA/Pzyso6QWUCeG4FjPm+qiEiPTBXFL2FGZ2sLT3KJxhsrudvpYNqBzHA2DRVi5U
p/0JOxNKAmgyvkSd0U7d1HK5r7u2TKVWFiaZYgd2nkgEiOHXjCL9lym/Mrc4J0vX
Uts5aYu3EJgZeMy3AUSZBLiro8ZAMH1XF5iV4bigmnOy5zlA+OtFng1FFplA444v
E8VqcjHmyczWkzAAA9sCFNTPy7T0PTzs/AeW1qLV1o2RZw7hydNYE39U96noq4/r
OmLItYNneIbnbCmVrRtgkUpjfba0aRSXVQX2lKqcI1U/yj1IaEDSuBIZTSQJ6siF
IBwT78waRWTuVrjxAtQz6XJcZS6KFCQzp/VUCqfnXK5OYXM6zFobVIIUSIzauf8z
jp+jnwJhgGlJ8OTQff1sFs0GG71nWVwlnOPm0a7i+iI5ieE0w0oPt5vpH6C2OZ/I
VtVypYGL4PGhkM7LC3yytXYgyE2AhTmAY10Zu5WWCz2rsmqx5M/P62Erqutxkutz
UJpB8IBMFcx1+04SnGcP0iCNC2B3Uo5+rD9MO10/BUQ4ONx+bwWXFsVMoJneVrPU
Z0sILYpHXNg2XCJHk2hod9CwAKSfVxBO3f6vjy/R6V20IfWOGe+uJz0A4OM3gf8v
wjQBsH8A9Whlhrix/3gdDZVnG8iYq9w7znwhEDbUFJtVTxKAoW015caG/ght+BBy
ON7Nbh5sPMQm9XMh2xLNPEFzQNv47PSkgL6BrfOxQbtJzuxLplIwhDlSFIDAEyrc
RwChP03Gn2xLCkQoHaHV6SrEmkfHS7pB+Z/sJ4DZx6IgBmMWD8dIm+goKExZLpLL
bFg/NgabkOYnIhrjrt2aXQZWa0ndCsDLt4XJFQCYmAgoFVZV1W76fw0EPzMCQOrD
0JF+rwzrlLDLa59feFopvaDjnzCUJTXRcFsXnQt6LfZTPXBKXIfQdIdI7d59E1tN
wzJ/IKJmj816Sk7Nc0HRH8534oJcDWr0vBIA+GkaiPkd+LSl+wQ7MHFxZo+kxvEV
Jmtjj+sbK6gKwuO6Mi5vFcNSNASngZGEfPZqN0l+Tj6EGT3CXrBXP+bOpLyB6E/W
YLxyNQl5G66hG/0KxKQhgErGA+UQsLTVqz6T8bovmTHOvupbmy6JziotoTSCKhRk
i0HiuL5+hP95C8fBw5bkHoltYxmxewH6e32NCmq4juPlS1VAXX8c+hwWDXUhIryl
CmVZ9bNXv2jmbshBFBKAX7zMe2j4b81e7e1wMrg5AmCMD6uf8etT16abAzzlrqRK
lVNKlD4uXseI1ZlF5yDTQGN5LYYqdgcbN0v7l6bXRM83IFCOcWPCATugEbpLYktR
Fcy4xeVJF1Og86ukkOi9RshjAWPt63+79+3V5Xm13Wi+l6mkDicfFwGA8N7qndmI
a76mGlm2XCXcx3y/ogtCkjUnY7Mm4ofxKRSkAzPhFjpGtFLWMoGtPyVFFaXVYjyK
QSfGLDU+YoGRRCPFMFPiIJROI1AqN8wCvlG213ed0qdA2CxM9m/qnjYbdS8rb/Il
6DZ3ruBzHlJi+UnUomKX7/8aSWbJtBz+ZO8Ma3OUMTCQX/UllPnGjzVpmzD7oNP9
ZL7+bPhmMItlPHrOcAJ4pg2WVMzPoou5sC2LOXaUH7qE/M85EVdWrGBOvug6Gb8P
SfY/bYhDnrM7jX9pbei0u8pJgWMaXSKMtKOjqXlXdMkwg8PA8HQ4TaV95CVD4KE2
/rXE9Vgvr4J9F8JmqWFz7+zI3ph31JyaZXoyBSn6D9MSUTBi0tcyQnQzIe61FwVT
K9B5hcSrpW7RpLfKRG+ejcD1pdHlXINp50Y2w7E5LIy1QfCgOo+VMBz4B3wikbFt
mqGT81HaGdi+32himMYXcm4F76V/iz0/HVNKRY0eJujBbHpzWWOZUfFedUzmy7BU
DqfwRvVeva8DsdQVXTXNP5Qk6AabDNczWPVNGQI9yTYbYvSkDJUyZ0U9aelpBg/y
rfzDjncHePcPc70ICxRNvoi3VmM8iZlFtNr0RJoNXj9IaYz5tSIoEEwlqCB18KSp
CfnbWez/v3C0Y1w6VwhtDPtkXZAvZ5UUOOgg4v4on5ghepg8XD3oTE5pYupShc65
iVzCTSRIWu3Cf9QQJu/3HZKe71dewgxjPD0v0HhKuvUKm/4yehUcv37Gr62myjqo
w+JhiL9pGxnOB3LAJeF704mqA34PSfxcsv2TlcZhsghWnryWfqwUOlH0N3tF+3S9
4Un0hmEb+pYZplfKYDuohcy6qWif+8qhr2VGgNBOl8dMKGYIg/sDTc0IdeTcUc65
FKlLRGcBLzIUMYPPVdn9ykS9HTodrFsD+5Ea6anGcLJUZPB8Tnje4eOKdeu96tqK
KeCSJ6h0qzsWIOBnymPKsdIpE7k33R5P2GFH/ugZw/UXwmbsdBHRwkGid46K0atl
hpFOE6jByDwwIhPDfl2vWGGhY7+EFoz5O+BgEO/hX1EfAYiPzBm0Yt7mAAmMYYf+
Bq1WhBo4LQviEvQ7BZ7KwCHzgt58xDJXMeUaj7lTuqx1A7ZDz3T+1j7pR9o3CVKq
3iZL9zcECZAZViiyv/yE9j8X+Az8vJc4dlcR4xYgPXSRZRwzNAIW53vmm1GYjIxu
2o+hSUsidABoGP2mnouQIwTCz6xE9ahI4n7XRyiTuMkAQJ/935CBLR08wFiJ8t4P
8lzRe2DQ8XDRNk2sU5BA29neBIAaHYDynLL7tQxx+yG8Xj/PI67dSfxhZyq1QlyI
2Y04g4bzaEKIDAG64+pLGk3bMomS+2hli2lQCen7Sy6FSy17+9IdlC7rXdbjfqlW
E5OHnplCpOt4FjkdHIIqdrAiWJje9q+UvwlHxlC6fCGqKypZw9vpK8M8Rekn/dJP
6/EzgRl9gV/3HYPQXXweH2PcM2T9amYuvyPpcghscUF/cIL2oUxyndUCOofyli6Q
8qut9JkS0g1OOrVstlLxMgjD3Trk1zc5GcY6QNv3gNhMHBhQzIkAg3F/F2I27Fz8
NIVsZY7Hn8jiNxQO3BX1xRisZAQ+T2yeakBE/GUtokBM8FlgDhwWSP7ar/oWB1fY
ETlbMsKyN50uB/Q+gev3xs+1TjZOYqi4/NZsantSFX320CtMvj7uXvKJ41f3Ik4c
RYsRA23QY2sgADlIlpVwE5oUFnUQLxLoTS5vVFITcmJ9T7cKcNku97NNBVN/SFov
JIfE7/ZA1Knpcyc+4f8rXRDiF6cAcqmdUTsHfW+jDNW0Orm0/qdYftdqFcuPVK1s
diwxbmV+Ua84eYa6NTTJxkDSpZDPEF341Y0NUQvNOuNLnGRcuU6CCCfJr4wiuNMq
n5XqgNR0HdOh6dsy9GjDVjau++bZ+cxSkFsiwa7x5RPiCZsyAiftmYa4jr6cMb6b
yzSKp+zMxDfEkhwzm1b2Mh+/2N8UoSxd0uB2UJnLRt1muaTkynOPjtIiKGN3cara
nv6aa7NIUF3HjWJW1wlxH1Z3Q5R9EOnsoT58rMfG3mk50oGpaPlyQ6EkV1IhKy8p
E4nuOevcEEGT/qQ5Mq0ggbmOYGsVZP2g6WA/RwD2BJaQ/mzr5bVeC0RNfD3nMszO
2fNRvxUbg2fxA+qOPrfQ88cCL+QK0vt5xYNPghmYaW3eopdhvIHDKC796mICbCXG
fVXgdJ/f+tDozse0FFhe54tC3qgurchQZj5xUNeoGHfCahD68iMjTSC9Dgbv9eLS
Qj7/PDmdU2FQcgfZ3IVUadTIIF9iEp9cM51WGlIyAhQ811gh/wA3DThoyguycQZm
GDw4IfhvJa7Fps9bVVNnGsZjUFcB1ke5h/rgHDST+0m7BabkY6DSFEbwUWuxh7NM
3f4bCTyr6ULBQQROwvJzWVFkSg8cwnWCanG5bX+i+MPPp5Fae4iz9DsSP1r9x8zA
1A90ovPTDKh55VgCtPLt09vSsBOWRSdT1D6KwdGIA6QlMOA+3IrUY2Dt0KU58bfh
bjuC4bhvJLQUwRoXnWKIb6evBHHCtDLyPIo9QjIM0qkT0N9aZKDuUlpyQSEOhmRU
rPTNztFwBrkyyxUenPsy+nvl4TI16FLpW1wgkYP1QSR2Fi6ekdaVEmkvmywQCpKf
qu7NrMKAdaljfLxUHK0dp1LYg0GGlBwpkenes21tOmte0DsiOI/X38WGGVszEVFb
HA/OIjD68LvsdMLS10xPUVIoAJIuD2fIr1CbJ2kWj98LhJDCPWzL9EYHQwABRX+R
ER0wqmTuZ4A0voRE4MSYegbZN/ANuFFqznHleaKv925o9phgiayT7sS+jeZY4XxO

--pragma protect end_data_block
--pragma protect digest_block
/hDZLLC3iO6+8CshKvGJ3cua7k0=
--pragma protect end_digest_block
--pragma protect end_protected
