-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Bz4UPMbS+BboD9VQcBsdFuwbsu/q2ZKYLWZJ4nLUxkQalWGZIn2wYPNAih9v61e1
ci7XnqlM6L+8h63mP5EfquaQHMJCr+PZDf9j0I7bC2ziNRCAfLxAWgshGuKXAC2r
FJwqBqoGmZaR4OyZXZRnOTR2SyK5Su+2xeUNdpa4epyOWLm1e3Sv+A==
--pragma protect end_key_block
--pragma protect digest_block
P5nogXsvsKr59xXWSE0XIXxpi/Y=
--pragma protect end_digest_block
--pragma protect data_block
qYV/FYT6KsJJ++TequS9pJtZaW5+8ocPfB2n2yoil4dMBx2LjIpr9jbFYW6fIbZz
/Z6QwIF+TQPx6Tv/DV9FIAzGW+5+6wcB4pvA6duYFLslUMwkkbQV6hMY/t3jJXxh
1P0XbuM6QyIlXa1Fc51AtkskXo9Zsk+QoJywbqwsRDGOCctnQXn28ZnvbN4ukxaj
I/X0iTzqgJ9zm+qipN9P6UJJ4xrTlmDGj8NQwZK7reoc4uGSy7DenKa8aD4iRuL5
UugbvVKvft5XbAeHe9ZnTaPJakWC7NIdnUmvXoBup1k9q4/2/hAcjtKXg3F9VfMt
QC0wGDKS7BIMjTFgZSXLVERuExCxgcpwzL5WFTruwOGxPus4sPwDd+7w5OXMXMZM
wyzelTE6KuhZiFB5JQgDxvtYd9CueKbWf3xqxHaf3rjMef8kcPBNpZGxxN09W3uU
2mtXTMEm5JEFe/gdkT8NuOKb7BwQeqMeSkavJpJ113+6cMvXcc4JGYzogDKqeXR6
Wu4XDVeq9BaWrDF+sZXU5NukCdViKMi5+WtqghHnJXE9SLszmGQ5gNjdNZbCyJaG
PwauGTf+VhQD2sOrAvxJ0eycK/S4J2d2XQRuVXBozcptKxp6Ljf4bc9jJGr0x4Sx
zrkaMZfR6YnRkYxIWl/u1eGKl45rU5j+zI4QZ3iD8NcuMKxv2VJFpSoSTAGuMAdS
9TtDNRYs/AcwRF5FPZV4sparTc9PTCBr2euFZEqOn7Tq4RHfO6wZwd0kn2XuyIxk
VeDT83DpxxQo5YUq8p9rcgDj7yrcAs3aKmfdP+kObsmMr0II7Ajk42bX4EfPjSCR
Vws8CABZkw+/KT968wSxQQ9jfu/6ZzFvlE0Gc/JxXRxLo7bq4sBKU8q+XoemfFWB
Mk6udaCzMwcnrxgcoBxYtJeRJ83ciUuT0I34B8pXu3wk3pk4tBi0h9wXW1Kuit4b
2uoYohGllVRtrSsnXttvTS0rJ+Oiv3AQINNo0YLFnZ4CgXWHkU7E8kg9RDZ3d83a
uWRSaHCB5Ta1bKa2qG7LO7wdCLuidcDTrtuMDP+d1Ik2jcFG8xTcWwuLXjGgRX+4
q2ulBrxnBdmkqYlTVFAio5tcG1YnRcLY26/mU0MfW/Jb266d3YkzySfXIPpPHK5h
SLBRcBDkCicwaormg5bhcGXMOGBMf3MjHJJWwV+n/zrpu6H3HwhUYJ1p/beFN0eh
AQ3p0R7/82RJ1x394tIUkvx8/GyHnwGAFqatVf05ZpAicv69RSkoJMvkTklr3yrG
ol6N8Ya4z7kFfdtncaKyTJxm3FqsS2CLDXEUKvLQnRi+f/fp1UA4z3BF8V4YQZOn
Eb0VKnaU+xki0Kd5l8OPqo8fzxoFEzk9IhPoasOVv3qWxD9/1S1geCknZqAPdi0x
XapSSTtPxCe1711Nh9eSMUGmJG4iTK/9xrrNIsTs7XQ2DGDiXM98C47MrV/FGAzE
JNg8FdHY846jYJ4npW5ew3TWdG6H+cW/ARfHK75S0cR7XRkNq6lZ8I5PPrmeIwDO
IByTw/N0xT7IHbcwf01UbczK5aiZZQ9i6Q8xEzzTAWo1zpi9btv5wY+K/zw/2hg8
ZyGzaJXvgiSTtYF4j7bjLEutrLcqRY32w5GSgxeSVxtsYt1yGbsFUh2E6Z4NLQRj
yqL+kqWhwPRv+EiLnctSHTcD+zI1aGyLAaAuXEcQZ4NeIPf/yx4aQgShAPzmsxGO
Crx/2MOezyO52qhOdzUX0caRS3aJYgkxzwrQCBXH2MToUJM/YgpFyCthRPjsPGAq
9q7KVX5jECGTg2vKJ6ZmhSCnWBytzX3pOWz3pENL9qRN25tTqBlJJIUT0NPGaYJP
8WNf9FYHeB1fI5NuoHFjaAMynegNfwWGJTw8rEXd0OqsJscK+87PghNDZzkmU52E
VNHq1TIfSEsvC56hKpLkN6HjJwZ3ApMqCbwYmZ0XESNqQD/Tv/leZG7fPUmcnML3
DxmwwGQU6Flv+UgZe2AzzR/Q7/LMoUCkzXO8JP4RPTlms6ur0NunlmB3InV/bJEs
EI+BkCLXZd4e8m2mPzfbU+bDm7hmzp2R7Ix5kUEWqvKbjYHcVgOzxZXXNy86SpiT
O6+WSI/x0AQL04aTepwRn/PUTOf9ogMqw2j0knm4gDuBLSsmrMnsdtJq9jVZziYA
50M7MdedyMXWXipJo5INZFfxrFwq/MMgIV+06I38filddViqpcFGCWmEvB+q+dFa
JJnBHhTT3sM5DXU7lrYWgKMx/UuI0gjY3eZle6cVS3XRmipw34jyJey1ukVMpQR4
r8GaJh9ZIniwsX31XMmOLnYcVdeIf4gYqVBqTRPBiere+6NaNObWI9c8t0rGcOrt
a80iF3nn/FhFVrbPdHpm3YbY4C/UqoI0T88JIt2bdNxwfBm5MWJ83ot63j3UbVuG
C3wlTm0tpZ1GwOcB1PLScno4VqwgVP8i4Pu7wUqb6JTRf9ZYbUaJr7jznUsWIide
FmGq8LAE58knNIK0ZO3v5+sAQ0AFPHIejnwwr8SC04NWD4X7w/hkaCcnAaTMM2KQ
l65960T0iVE8dnfivFwGjQdi18eYh/NdnvknP7iMWd0T+D6yGdAHHN8yxvLzr1/Z
rjS2BtwfgaExXnMq4BVuUUDomnjbCDAJNEmBI6rbz5IPHZe2vyxEr7htHc11vfgU
iH7sLGybC5iqm+E90cEtvDIlbfCrF3mxp9DQc+K+R6ly7rKK1Ym0xFUhw+yF//Wl
8fGO6wuZY22aZI0feFW6iMZf45YMv6jizRInee+aw6DYezA46uVxC/SwgMrvapzG
lt7V5OiohcIO+mxvzcbP0Q/zvICyrCdZFhANkozeR9r6AcANdTZW9qEiBFVy1Mzf
LtXlJLp4hyMM04yqT2uQE/tPzC/OAZbVhnHe0/hlY+x0aDupZa7GmcL0i07if+08
kn5RdN+KUranWi0jDryEVLxkUkR/xXSvXB0gv5c4bnU8ImidVBl7pHY/7vr7MdQ8
zhQRfw+XypKO7jSwdO0aqeTJTJM8wWYeWTxoHOYdgDOcRBH378yln01op5dlhwZr
rruzh/JBM1CXsdyHPjfch3+Nz4xyTV4korypqYkCiWoNZU4AxfFQoU/SCBjXJvfA
eKqHn+GgIuAVd88WmxB+WcU4l0HsbQSEgzOQFUlqO0WbtMbZG11YnFN3WBBjJ7XC
QBsBAlrwfxJUfwkwXxjkX5jJenkcDpFpwU7CiiX+F9Qxm1JouxN5Dkb9EDEkmzjX
5UdfWPFZIM4yyj1fJPTKVDGlmz6Z06iLFKcdUSg3C+l2Q2KnSSuv8Foon6vUb+6I
2gVESftTbvUYw4jIf+JQHE3IuQBcgiuBE77ZpRldF2EXk4AvAIiYGp81xkFjTaiR
J7HkX1uYTzo9no1yjGWLt1NpM0tI75AUv9itvjscNE+GdhP6Pjq61DzmWmMcxb6B
yZ7/6M1KWsKrSigLoKUs0ympcLcqW9uHjHXrnG3GsEXTKXJsfJLqOrVUp8HxqU+v
OU1ripjc095fIMM5+JtjoUCcOm3uisF3H3WGVhtbm57hNTM9iNIgZfAC5GXYn4Pb
ZNXsUZvLpaid3nRZOTQYr+pDSwXKr1u4DKJNMFW746GPoAlZKXHZbg0VigjRO5jk
3J7U0tTK3hOZyZ0ZLiRtsMo/BzKE9uWtGjt/B+C45zh+GmSHGIKUu4yiInzc+tNL
4cDjAeq6Pu3BzgBizJdI3bHZTy8CS4mYLLEE/4HIULU1TbItfp9BUTwTg7pSMKGd
5TWH129KWkFRj1dITzNSnu+p9lBlDZ1AmaiwgVivZluxAoCgLsdoDada4TFdz4LV
t0HfXtxPZLLrwVyYx3uFcbZWGvHvuILQR7u7ehLUF9/8m8moJlEG82tWbR+gWifW
cfZ/r7usWMgNP5SF/klVDqiuyqu6HCBi51BqqNMkP/GrQ3yRdZjjKmVarVfpupd9
AoSpvnT35eLgqLUw9aA/IMXMqreyjRRpdAixq5Ep+RiMR49q8xKvodjJoHRohCw6
TuiQLm2lZInMaYeIFlCZrMuRHRxnCm8/XQrXmaa4ugQJJfR2IY+n788buJBlmHLY
kR7zmX34OQAYGcNVHD7HaR+BfExYhAnTjMdrt4tlDD0lkTkwVYHaZdgGsANbUbLt
UsWHrGGGckA3Tyr/gxJkJNuotS5rBv8DSvKi9/eWfbi4OJ7g7J0MY4mOaDsHVYgs
WpDfXL8V1Ciy9wBL+zrytkQjhwD6X25Cnbr9+oZ0ZNsZKER0LoT+tIV3uCt1/PZ4
QFM8puuFjToECKnGRa5NhvbIgljxXOnxFFEreEIdEUoDhtr6Yj+7S2bKHUQXD2J2
QLGj+6LFVkubn07DF3Ay7QcsWWEs3mMEW2zzxfKD3S85oBWBrCGf87n64ZjkBhvp
YQsWTKsq7BBqFLioVsfTvtnghdCyRP6Xt8/b/P9/d/RgQhHOFYrGO+xLpJfzE52q
IXnY8BVdjR2ki9dIdQLcKVAQ5bofgSACbJEgPIG2nqLFW/f07jbRUIc6fTaQ7Xis
eIPKS5j0TjRZDeZVtduirsZukABwNUZT7H7QoDH/Qp/MPN3kWp27nRuMvrRfzSAM
zGtW4NsAX1qFPlSITDi3YHQI+KtdUzNW4+sgl+zhJ6hY5gt8nIOzZumCVE5ip0nv
WP0mhjbNXjvKAPLjikx5gDw45UBFUw1ck5hCwU773mA8ghCEWM9DKm/M8/7dULMw
yqmfNa+dH9kGZf5y8XwG+w2PQgwqK3VEkr/QUPdLG7gTFAmiVt2XZ0cnmc74AuQg
CT9sc+3qQ+w8dY4zGK4UjJsv7za7Xkzv3Y65MsnU9AKSpSATfZ4iYGBxr4cZqp1P
vh9aGmtucRb+1ymXzCxauAiaacNHImb4cgRGgWMuEy0MgEQYzzIvmLn7sZkgXhBs
sV7NlSD46E8oubTILJUpkXHRMEv93N8mMD96QZC3gzVWYc6Zi6ZxZaXq+GqTtt/X
/u7vBpnNe+CUviqspbmLsJVIqjMqotkPDzQcAYTbTeqn/uDwtQIm9YF2Lq6IvUc4
bA1V98lrt0PzwBuc++abeK2CMSVToh+bzGxGZaINg9U4J+USRVdTOjHNwrWoR+9e
zDJAPR35VqP6P04A1Uc2K/ua/r9203wtHKM/y9xygc6tmG60AM2VI9wBjs7UbtBc
Y8Xr9Gd0nBFbpYSBVQQqkSb9C4sia7jkpmsxO7eHZLw9eXAYRWEPTYk2Cs+MjA4y
Ra77HMUJxitz3bEfcouY90Ai/XNcslOjRS0QhHAL+OdAFxlZcP57GvqOQH7ZUpXv
rwbHgfDV4fnbjth/sl1d/McQJ7dYbNIUghNs4my/dSl29v2uxyGGh5UPpOcbpuUr
UxbuAYjeB9pMJ3x73HValbyp9UiQ0IsZNRwNGCAEdeFUVX+FqSJldk7Ap8tYN7c2
1iTQh88d7lFa1JLXJOkQKYu/s0qATbNmYMMUpsPLX4HNKG2pfd7YSj50WpVH51Gn
UGwHc8E6srOMiMq1vjmeyDlTh9UUtWSZJRZueMSYQeHpcsh8JYrvmSTs/6aWAG3Q
wQa0/kSROawTn9TZxH91JTSYkyb56LHTsDvHLbKqzHYaIpOz8Py22C2IV5guNUac
OeQmolxiBo84OpaSuoCanghbglZBDQv9druWAwr3n4gESF5vjAOaHzRNYXp/gb7v
Y57p3kUP8wsMSULpqPrWAJ5YJ9BsEoAhm3GPvjMVmEl+ORtNjI9iF1oepc7PyBjO
eAk17tAb/8iDCjguS335/4CyMmfEPR/IDBxD4vSU9OOgGJOLJIgXVaeTZtOHIowp
/+DnZ9/gfkiIyMCKyCBO9DHbSbO2YmX4bHWHF2oPUuGZ+41Tmen5t+MrjS763vxQ
nZLaqBz3jjpkAp8/5z/nIe77S1WNagWY+DBR/uR8SvAVV77uCwvwYHHwJm39+2lb
0ndP0rdQvTsUZEncF+fndkspKhNyybYGW1o5cEEtEhfz4x2PzwnOsb48u1lUyvv5
F+XJOm1TuijulZ0K7nTsw/RlfOTO22U7DK4zIv05sow+Wx5RAqO63ILceCZjjXp0
oWVqjPhS+UGomJvi5S6I5t6aio0gnp5Xtvgg4TdysHm0uTojr35nF21apwfMsSrs
UF2tuOL2jT5hY1XsSaIiEx2MsqbW8EXyimqB87mIkoIfgzxSrkVVBWeacV34PT8e
yIhh8ov+nJx8h8MoBBW9wrv3izVSAHDSp/9TZHdC1ficoh0cKzQgjWCVPMRdwYh+
3ldwGtB6wzztlFhSGmx6a3l0uuwTd5au+dRZjDW8Fl28zs+ewKyqoA/zb+mQ+S1y
zgtj/l1aoVayf5cetzULbyZ9SSi9bdEqLxzkbVg8V5CiUSAHevjIIzzYOUApH3Nc
ple9nYYbBRTfEzGjc8BRHfVeDE4a7g2RcM7fiPvtxGAeuZ/OOzfOqZZb5rzSm0V4
r+Em5mji8qGeHlmezc/uX+wuEsTE7t9iQxTVChv7xzP3kGyf20LsGHJ/I5ULnoBZ
f2Fi5G4elHsb8sX4lGx90UDdO5KBuUOfVoC6b4Kbf/0/yDKrBxNpr8wT2CfaYD1+
BLBHeweKbgBN+8/4ej7L1ZSm8o2i9gBvGsN4nS0xatoFFiB/jBoHv9/abbxA22dc
R/T5gLYEtJVpu7Fxh2nsMFlMQGKFEC19/t6P2m+SKMdWu03MaxbnXIYFV7IH4bzh
HMo9Rww758ZBUMaminuf5kMqRaDmK+2mc8oRBOsl5/4a+j3SDns5jeZAuYK8ToPn
qcPQIIQcLPwvu5dTK98AloL2IzQpOPRgtLLIYjfonZhWwH/IBpcvqgpvBzq3M3wS
qbQwut0fEL0Zq4bfbVEX7Gi+WCDwpaFImIf7pxC17B2CY3MYp3n0M6SZ//YKkRm+
imgrxcSJZW8M38ul2w6Z8yAGe11Zr4KyM+55VDbUxTWG4PwH18lLoXY9HUuxKVn/
9Cf2hknR5FQ9p0bU1htdggD9DoV1stC90ex5+BXXtAjVTNRpPWFihXRdiQmlIxsU
dkvhIurQxtqLzIf7w58Ml8xy738hKK0CaLsUmbR5gv14IJRXz+QLH+mPLyZeLxyu
Y1IXd4PP9SAvDmCAAzd89Y2WDhz3sFnyMmteI8/wYPP69Ao9uHLVehaS4M2Ezwvj
rYa70XcONJSZRUNkFLXFId9KnN+pfgVVIdRSD1HPwsPYllPtlAGv+Oa9jehRrj/O
qfoK77vQNcXu7pMPgDLKuuerNxX3nLkGfaLqwb4Se6sm7AyPr1ANKKgZQb1vMnFn
hZmIiLueeOu+L+srF+0OLGtsN17ACjQgJGxf0zV9lsJtWz+yf6bv+KzATSuNed5c
K5+RPKItGDpn4ahCtWvCrb2J3D10UG1Zl9rd/T4ij8O3phD20w6xX2EzbM7f6NC9
e2ov9hSdamQI/yPjyUt3ujUA0q39E1EhYNNruYMX43zzBsk0LPR/TxqldLQhL7t+
eEx/+VGgd4O7oGBEvinkpxk8hewYhssQRqudRJxWiWs+rR6oCLOHnbydIm1mR8Of
j8ZcW7VY4TBwzEkvLOCMfL5j14rkJCAUreH+UqMl96U5g2pPK/+ug3l1nEtNqOPt
qCrp/lw9qflFr/ZVCARWggveaO7aGEjYqns+SbmHr459UeL70biDlr1X+yE3xMpF
aFNekdhGNYs4Z8w0lhnDe6zOnqqnTWqhX9TI6OwXDsS3PD+iyQLYcDYIfpqRLVol
XnFROtBv/ycy3Q6aAU+voHuVaoFPE9mcOFMQX6UPLohwzaeieCkmKYkE9Z6ps0J5
/RV9JxKKS5lTFFPwa7ZsP0a+8fL2muRXWF55D+bFts2km11IpF1Ua9rK82PsG+pQ
6scJ6ct/Qyvxaw2gN4TX09i79vVOB2wJgwa/C5aa5yNnMGJVo1LVrxXv/1yoiV0h
e4qQW3Uy0HKGwQyvBDbZDWmxD5iZW6xPvn+FACqLe97W2y6ODUygHuR76btPhogD
TlXD2t0Du3nc0uOCwxUp968UrszrqOKxhzFnecovZGLk14XfXNAluushHt3hBsD8
m9B+zTXKY6KqoU/VlcPDWbKm1xWtp0WYamWmzcxpNISGwijdqwcXmwgDL9TpbkiA
NoD1Zrey0wlvJGkW1kAK3MaMNqSvvnpbkWUgIGh38eLYzXVFVGStl9gd4nzOhRny
XFnxB9++EzBilr5hEsi/TL6mcE67B4buJFXY3d90RN5avlzYz2AKg3wGf7SdaOgp
JGAtmofmStdgFV3VOxRXMtTzN0RYRQkFNMQE/qXelIMeWKTQmVMLBcWg4YkTTQNg
szt9Jd1kn5cKWt/jRrErqK7YVaskbpAYceHQR8F9aiNTjprxMb3+hQZDrmxeEkXr
Zso93ijAMqfuKmTS8x0aI0cD2LWsTWHdFGhtHqRumQfYjH3Cd3gYWaIUM2OMNe17
up41W14DIqCEdZQxw72qcRw4FNxS/IjitWN7afduC02sTX7sg157QcxUiO9vBMw1
rrBGH3lzXBhTaxTk7KetZg3IDATntbE0EMC7PZpwkOMW80UhggasRA8uIGr7R0jz
z3M03UkWQ1QQK8duyC4XjzvSfTbxCpBI8P95YzWthkx/S7u4H3VWxH+OTMVLpBBP
DirtTxCE5R630LsOykaeioRIglx6dnIjU9vGFybu+pIHUr8aNew0BqDRsu9QYfuU
tlL2J/Oav3nzMDGABct+vr5CMbAr89eRs0P+W/Xgb8JibqFWdJUZK30Wcj+k0TdI
LLHxIuXEQXzos1LU/jXXIZCzuALLRGmddttXkkpHBAXqP2uflT690Lby18COFuLP
w7HveZYfghr+aJh5Dsah+WfYMR2XHuv67nrxXNAKuMY0l9RuXJyzcAwRekcUW+cr
cZpoDZolSkkT4Ja1Q2x1cmlz9lnJqVDz9MvJyIbdWqH9RLUY4/0uHA9KuMsWYGNG
lDj7IgyndDGugkx5vxuPtffodmQXQ/Y5b7tMHHmtHDZo/bf9SrDqiA66rPgENzxS
J+B0FhaVWBmhjuEp/6Ir6MF/AXY9acKw0QMUh6NqXX1G4RCVt/4DMhVt+IvH9L4/
sAa4x90yuhI1JL+DhQfB5wKZQlAaVJUw0P7QsiRcwiYmuR+mTubhMCwBUAotCXJN
xhaMWZfHx2Ab91uQpFl1hIMoPW3R6qmdgmvd4b1nwyOLMRBH0G7+QNFxj2QxxhIm
1zuOOtWsw1GvQdGpV9NZzOfuFwmobfypp1bRp4P9P46Nnrg8RaBohrZXptNMuKA6
U46cET7+PhIbRB0HaJWwzyHcpPMs9rYtewc3TjcZthfXOt6xf60CNv0e3iBr/SDh
PdNtDsbghvBLmKpDaG4UKiw1JZFYIXZTegkZNQy+jR6Ac09SsYpUd5RI8o/t8mg3
bdV8QvCsBBucWCT06IWWTsAawrJVma8aikSS0HHOixSZ8UJwga6BNChS39ArAVOw
8xy7PwswpsiX0HJdMQiXBR37RvZabYeh6FDmw3NiAQlBad5jcN+Xntqg0RnA961Y
oMWGOHFNJGYcOJKm9/GJj9+2mbQpS01Jtak9wpGw/sWOLSNuvJULRQ8UFR/G44bY
CV+5mA4rVoPqEoJUo8cWXRunmIiI6TE4kqdlwDthdZOV7fPOsBJyeT8mNs9rDwuM
jEADB89HNd3Zx5g48FI6sW9jN2I/31x4Hxa6Oq3XN8zMwLjvJ9cZKRWmL/OCU8bI
CN5k0G1LszN0Ucecf2TF0OwSx0R5H+x7hPfyu9nvrUxZR3EFSoD3EddHAbc2U5ac
MpDYO908Ba0g/HtiTchH+pGhnr3SqQb9//9u2AEs7BqwgPZwDEa8DotFxw+a3oou
OCW3lDHJdJFWoVcAIU/OLIogblCht9tFcxttLVD7gdYKvub3t9gTBe24MgxYucPv
xBhvUA6z+3MqRtI4qOy5p8DlPhYvr51f04x8RHq5Els9G8ffyfUvGNX1t9f8OUKu
dmirR6ewMa9YFH1mOkj0QY+HpNYOrdpl6JGawTB1EA3ePi+N6PkCziKGlX/mGnGH
WG2nxa+6FKeKWaURWrTxE1RjgQRBoAXEDBRZmA15wsgBCdE6gxTGYX3VjfPtnjHn
zgo7I6tVaygkUsorRuxQFo7AUIEq8Xo5uIjfMDdxrBgmy3zzSt6UbWu7dN3Z+Lvv
WLo/fNbPG+0fYXMStaDqkG1uHFgW7Z7HOJ1L+vXzJGZixzeAgNp7eIQdU16YZSRh
SlKN6iFt2LTF2VX11oXDPQTR+BAoRS7nvdKAqR0D80RlaLRMSkBA+8/jvjfcZn4B
8RrV0CjZfRXkAkZR6ESy+ogGxgntqo4sTMLnrGUGMcxwqEkvbCSwYX4VWRUah0F3
yJJybKVTmBCOl0K8mS/s+A9sVqY1fKmVpnyJ4Up7n64ViAxV4tWkd9GTirMqpttY
Dz7S46JNY6bERpwqKVkY7Cf40yWU1KNAADxpNdY1k8+9V2Bv+sQ+afC9a5/16HQm
qFc1zkisNd6Wlu93bln0lc6qlXDuGiOwbO4WksDjHtA8FErIP+TBJ/9UjXikjFzP
tGyelbfN45GAovd5RBI3hrrOpDEZscLx7rzIPFcZulUFdOmPhua3kdFhU6aAUGN4
IdEprO/ye2On03fyItbhU/GiPnAytiWJfpXbW9SVRbZU+MTuP8ka3GJvl4kV5z7c
KY7mb5MQ2AhqFWq5D/5lD2t0AkBMxpm4UXvLZOxtn6a54OJqkqVwzutWxdoXfmax
lp1OlJ993G8zIBYh9UyWM6Gec0ZdnqfFMpgp5YfOKSV3WlmZCptiwGdqxw5PMK9f
TFJ05xxPntmA7n49E76Nxt1fknYzOwAqhoYkaouQ/uY5qCmWLfaakIzAbcqKNGT/
eaIYcbeGte6Cy+MCVjqNqXsq9q4c4N2HcxkFwhOwzBlTK9t9SEXcPBryT6WEmX5Q
qxCOtYRDTKzquCAsLtyjHHgb4hbk5J6RAz1Pb84RBdbKMrAc68JzjcfFe4LtAfMn
F80aJBOcRLzKAjvIWI5DoZLRxU1aOVKaAtVVXLrBZ3KHN9T61akY3eIfemoChLIV
/jT5M9m4EH7Cw5GiTyXUYOVBmAr2+OIMp/RRztLBKioR4xbKABEpIdWVGVho1Xbc
n2EsV/aE4NCsuyNkCWzuuPdJgEhxUy537qAzeKCjfL94d7twx0kztljXxodMgMHm
XMo6RfVC3VCiG/8HWjal4tpcKwa5L2qocVk9yoOzBJ2cLaJ5UhWegtfCCflUuVwI
TIMxr6mzpgXCUJWk5uacHPG6C78Noujcm5zz9z3Wa9iJsyupKlmD5QH7/xy6os6z
gVrB83zgcjVJ+kQupocjEIZ9b+rPG73XW64ctCefMmbMCJREyHX3fNfme/sxqAE+
w7fbuWweKTrZsOYwz9hPgy4/BhiugCObcMOVdmLJLCm5grtH+Jge5nOv1CtBzRC3
t20vRdPv5WT7yUlDkVxDn17/qrivrchIfl2qQ7GfM/vi2oKmdsnD9REIPL+BMcuu
gglVov90tUqyldJ+dtpoiKdrylKN4r04QrJsK4KODJ8YelgxwAYn1/QEbTu+irIZ
qaDyGuHoKWzuh5FY+WXjfxdPrV10xWGAxvgiGJbHlyZKfqy+i7bokO2mmy/ihAYV
QsV+0doIyUz4IWidML34I7iDELB2OajbS51KsrdnE2b0jFLQTadrU7oPndIam/IX
JgpfZ9jYxyqFpms1ug5sjSDuxv+uW5/dR7QiFtZ4GThJZsyEPWToc7AL9LW35NMP
vrSUgwxziQCwmULskaqW3DWtGgbtrMW50sWGtudu4JqfrEcDE0BhEa7s4DXXFLQ8
ydjFVaxgbtLtGfbXXKK+4Bnlr75Zr6jMYh498eDy0N/SHukWq6KRPfkYzP5D2fH1
uxJW3gHJKcgrd5TRciNx1nWa1TiIXPCo684ndI2xLUCjhgugtjfhpANHzC0TuYYf
o0kQjY2hazihbVthf86BdRH/rYR9A3CMNqL2DiMjjiwcRxY2TCvLddi99/i0asEa
FmVG9IWEB/mbet9Vsb5QQxcV1YRXsmNVo60QGOXLy32oMt6o+IbQo9MUCcrWFNen
jALTpUzm29zIcBU5M4tzXSEfKPvIXvoUKUaeN3eYf0hhEDdI3WYLX6a36MyM4F26
LjXjTE3T5QAn7Ho8TP9gftNYYHntoIdeheNSkTrgyAkfzOEJBxa/KaW79E2Eby7M
MAXQJ9WJD4yeEAPMnfKlkFP1MmMjwcM2+4sUHOnzXhUVG8WQd2AAno4dxQK7S9K2
X1GB5ia7AYToThOAvRRTtxIDNc5KPG1dVB3oPSNBGl2qzSddP4che20x1dr3C52/
pa+fxnyOzWhAZGJSw9iFgh3b7SaCO4ygPsxj3u9H0QJ6Tl6XITC9rUPMeYfBgufN
uQrDKB0lRgNpyD7lcUJ6OrmlRHixcCEP+J4Yt8AgN3NvFQkxCodjbid442/X4Puy
3I7pyE/8rPDn8pQCky7nWMe8qlaB8QO9vd2Tk4Qr5eXsrhrnS7JkbXwtTIKVbJo8
1bw+73N2An+mOfhtF3taR3X+9peTtXtDWTzzj5k1j0+ugXQ91cFK1bVQgSW162d6
4z9kvEPxQmOmyszuaHGj1SPWgR+ohbhfPy8MHiqLd2s6aMDN57ARM7jpwzI0hyif
a0zqWnO4mDxpl/IUdx23Y2aT7rmtuhrlLO4x6c3D5QZ2TX6kQ87I8Y/RrWvClZuv
8EUUDYSKUZ5LNix+mvQcANo4xvgAHvGf1WdUOb2pSlVpxrxP53AoNJtI+SHFZhSU
zezX+WyYa+gQt6kzEGgaJ59DPbhhz3ly+OYSkZf9mQ5RLKcpsGDYeEHTAKUGIbzA
IgBK2wy7uz1wNkwV6KgdhlvU+8U5iWtQOn0r4lCdDtien3S4CLLRZLomedo52Skx
UVWRw7Z//eGq2k4emdNHVuVO0tRkBcK0ZBtG+NQDVVlNM3VyBUvkxxp/NK24a1M2
YuJ/f72oWVLHzhebIBwPGI/OIF3Kus0hYFAm/Nm/BEv2WJJhY31ct0MFdxct7Sxv
CXIO8qew4/9JksczeSBCNkUTHfYhNzNdTPvuTULgsCVkmhFPXYkJGGfbhbvY/hAi
8nBMHeBtw2BW3xzU+Q0ySldC2dc5cM/sHnoovrBRkaeI2JU5JNGLy7Ez1lMi4QdS
ZkIpKdLN1RjFfHkxz1GgRR1b/pFxABJGc3KUZ1e7JEYgJr5RInQtta/Tom8aB+ZA
N/aXy4ktC50ei2bdj8fkA+G0XCpaFtclxFPf0G5Ljy1RNzOYvqy+pU9mSMHXMnSD
zikLl1xdjbncpC5apYGsx7XJ4j0rojuebxEOC+ZvFdkrEqrPg8e52NOnrnqwCeZA
Vdgr53h9EmU0YZoYhQIMtMjozfIspO+l46qG5XMBn5TrZBX4Udrvdfd6P6Zh+wla
2XTB+vHl7DkeGra/TT2r2j+w9Fvw5S7Wvuyl4jdtmNzE5XG1pm6yhRsrnzW39DkZ
tRu6Q1rceyZvmtH+nYMDdAUrgXYClNVoFAMhPpi/EBYXnxybO/kmlwp9XmIgYsW+
TECThTAnOE/zVbA+Jc+8EEyjc/NBrGu1PKstfl2tY8d8RTgh4l0A5VJ46yWW5D8z
zIkPd6O2o5YVMBK/W1KQntX4OJeU1P2gmIGvEB3X4VN0kcSOTmXn9RUi00tQbfTi
EffhsWX0LT6UT6HXwGBEzl9ryssSMyqGGELMrSI/CCVQEBulRzhQ2oZDeeAd7OzS
E4vSVK89XEPvEBEF7Vsxv/XmSN2sNkZbhO+WI/AEDZ94ztAFwEaiELC5zNXoOEb8
yVl+1eEKcisllCqh5ONRZ3SRY75iBtRp4MzS8QsG+3l2o4OAVvmylb2JE53EsjIX
xlxmIwiHNA4P6ir6ZtHTbZQOud7XMwszpO5dRSzNerz2VuJ8JeFfFhXqMNv6icjC
Ktfhrh68yTsbPD6KhnmLDDDVfocFhx4Znvacq0eF9bwy1qI32YphP5LD9UryOF3t
jIFzpTnR/cuIRqk1LGeSmD9IKpKkqrMO8nSzSCmuDqK8lKRHNDLoHXtucdwVoDgN
Ni3OIr6HMQDfrMZW3FE2VmxWiLHtI6mZV9Qsbysou0m/woMqf3bc7ZQZN4SvYTl5
5HntFiHvmBc1n0+CeOrFbPbBFVeC4TWemUoZrj9GiZYTiniY7KANl8EUWwVh6yYV
SyS4/Ogvl+jKNIIuqFGC1s2c1Wbvlx5Ou5k1Yn3M+zfUSx5J/GEL0eex/iZPuJE+
B8OnvB8qw+6Eaa3gUS4OLLvQEdUyfYHxBAr9pZp1ZfDBygYbTu854U6kBY7Hl4mq
xsHnrlw9wTlLKyw7Ug97gTR4dUhvHuzphwbQ3uwYdKQXmI+9RGhAwPrqwkFrkmLw
Tar/RPqVwN9uh2Dw0ljWzyWVT7cRZffAYGIpKPfggUCxTCEIOAIRqBpX3NEPAxhp
qUIC3Q/nMpz4vjbXh8gubfQKNIEAH7IFx7i1KijZahforN1SN6Bq+LBXgsyq+Act
2x9iLwVRTEjDQRCjdMx40PA9UNh7ZvlEpLXC4v5fNRohsCRkZ4TxLvn1Om9ANQr7
H54IOkl9HGyFwJ8dLDGXgzKUxcPam2k4OAE0Wv1ZrVrYIyX9+TUKSCIvVhUuSJY+
GgQbUzjxCWCRRjpeWhYsHhLCUtCPtg5tOOZuWQoaRQp9rJUn1e1rK4MKhcRDw7g2
7yEyoNiVTyR7qJqHd9MAG1VKUNDXDeoRNEMV1+NQoyq9VYMJsyshU9S+snwlnVxV
2T2YVgti1iJPYU0s3Ix3ifOBQ0nBr/uCMMvu4aAsBRFllXNxU+fMU558OeawN/WF
Nz9laEEwSYhtWK83nHPZ2gzxkqwVv5YQ8YGpFj0aUcvMAFyckrouJ1rftDxBPcrN
6YvzwgwmYuyLwtxBN/Q07WR6Yzw0DPOUoL0qyGViefFZEtrTJhCwSJdwdw7RrL19
3JHyrkg26VFeWjchC5sRSzDy7oi/DLiXgsHcxHDOrCyKWm2khNObxgWnLvLjKLPV
PDKLGFjjANy1LeZil3gWmaM520uwtgzxvf37Ioht8Sx3Q764lhvqKKIuXD9XrZMX
qMSdsSxkS092/ezWplm0Id01+eDWKxJz3b0ay1tsUrY0288ibMvrjBfhL+Sxrx/L
SVhvzQQDk7rw3XQM0BTDU+TDYTZ/QxFlMMn6DNIXg5lOTgXss7/NY8i/iECyV8+0
480yO5qmnGFxlsEVqZQxP9+w22y6IsAC4maCOvaDG9ZepinF07WJcKffLtBm7g2U
1AMJVnvUlsDqgvFJmHeWZo5Wp08JTvWzmd5I9NWnYdafYwJIgXPBE1JxRp9CVjvW
dh4o809jdTAKS+OepYRANERLAHg1QHRiVKaxA8SoxoNbD9Z8f5/hhsdtKliEfbbt
mvZ0f17AKAywBGCYmSbI4nu4PVfFRzCINhUAepv9FU0KrfUfWGNkajF/ULKT5nsv
R9n2W4P6BdoxUrtR07rYsq+b5XdxX2lgG/UR2DxhkmMD+wTwQytB4K8XupSq2cr/
EHQVZuPT3i1Pe7ibvm6Of/4SkXTh3KU3gOUdQ/Whd2ZbD/pJTqz5/cQGk67unckB
aRM258/F4ZSudLJMm9886Q9VhHZ2m9Pa8G0vyr5/QdPU9gQU9XRD3oKjOcH8Rsfo
M4qlA5HgzOyxuYZaHaw/zeAUVHbRUg1TMmeULW6QRpsbPNqJxJcR6D7Ez838ABNm
Q1kdVKpzIMzEp+EPabTJQ/g6idLynd5mcIHM21XYAZqBJ5zpONaOTYYHXwlUJdWe
7KXjGV2MjwOVZeIq9wlUtu2vKjDXVqO0c7NNWhQxAb3JuvL2JwAG1MDXdXLFySlW
jnPUwBrhiwWQm7rmfzEaEvMRJq/HjYuS3VGrKdTTHP0cRtdZWq/bXO+LqD2QVPGQ
9+7krceR3dVnQvMHOeQmpNNTgayqUbevrheb5WDYNLxbBFKegFbKgotd9v0iNdi6
LCunGyIxHN7wK940F+A5jeLMmEt5h/rz4uadb1P/z/fJORvQnQ4/+YOQx7WGweDd
4vqCQ33Asozn4KvMzKDJ4oV/vHtoZxDLT2nJVDnZ/nQHGktt594eQnk6WRPFMoqO
lY3JQ3Gedeay+/2jwE9/yumfG3VvOsk/HLaTCuPDz3oYuxnykhlc2cPGM3g+XZx8
lZvOp4wqik+JQsnrr1emUomD7/30DDMb4PkEiTd/yVgnLtT86VRY0cGm6khyuoyW
Pe9/QYXDdJ+lbe1OY+K2q6BPoUP1tcjdt8fG9LtSflrsnO5HcDmBeugz9zcBiDq1
OysMnMcTw1wFfuyZpaNvKYCkudpx3N2hPzNnwJ3ZibqtLfMrexsVrRrRmbluIUT9
tPGEFln+yh6BQaRr5SHUgc4sbBfjslC1xSgg3yMV2ZZx1ed/GPXnmneGIhRZ0LrF
aM3Xi+dHQsYQXICFmbzwULeLV/JYBf2/zPuTU0c+iBzJlJN6Lvrl1SeUtzzP4N25
piPizXAt31Qj0HEZ8+TTagDJFo6dXeTDVJTalmcD2fQTtFjCMDBlgjJDAKzR28/T
jsTfGlsK/V72c4kQitpL9m+lUO6ckANFjvQHpIJL0b1T6LbTyJG4T5qknctX3sBj
DS3rRXLx5R8Y4pCiIMh5hhRkqt/zoDSIBbDzBNmK68wkxmnGMzrbG/YPgx3dVYtO
uN7IukcG6ZlJuurO+YkJoU5MHvzLFjuSJwxXmduqAFDpDWMRZcjErmN8Gw1YNqQC
X1NnhA2Dt/iQQtiT9Z6vVwLN2NWhrKcinaHbrn8SB21bB0jmfm6vP7HsGMwysos6
RmgeC3+noSDXvA02uhRFlExpDrmHGFlg13dyMKU3UJpL36FUbKKGj8sCWBw7Tw8c
zu6YCjpWMY+Eql+7VCXmG9j2HQnZ/W7TaFPd9FEf4dR57RPru1sk1sGyt1gcua7f
bZFU0RgWFtWolx0+vovNmUi7oYDPVjF47a3oTtxRoBIbbaypQcieBTrqD8uZcwpA
+1DBcHhgJwbWTCD8ggf0NX/BeIe5Mf0dbwbt+dvxtQnpK87MZ1rZ2Vywk+TtPPoc
I/6onzyGHjllr6Sld3EA8Hv1UCP0rphrTIAiABfaLVyBLOxp3zXfySaYxexMJcOc
ThVaG/nJVLJ/4JRU6V5c9BVRbFTedT/hpPjVNw7+/U0oWbFGTQhutE4TUjFEgIJn
xNmUIygdjlQNf1U9PZwwdWfNalVS5tZnzsN87l8ivwT/VYUzhJNypY+hEcv1LUdt
tBk3ebR+2S4ke9aDFspjm8k+jSFm/uadJ7X+LNhno2O3NKPiNGioM2D4L7OSK+EL
mheK7W9qWJhPPlxO6u1zgia8k0lkvMw6cU+Q5iISTa+yUZjPSkpKZqVL867foKuE
gl4DJewotedUC8zvbTkbRAcfrMokYGKXzyQsHwz1vajxfS8mgFUNcESnIwJUbMiY
3l/t8HKaBaKE2smgdM4l/shAJzaigov6Eh/A6cgO/8UIMFNZuh5g3Wz48mr9/4sc
dadF9DQQY6BlYN/UjZhnVHTPvDQ/OviVQBijydnC06wn0qUfXByAbDwSJpsDABCa
HG3QbCxb03NrkajZEE5YOpGf2GqpzwjArQ5hEMerxjzFmNxeAKiYIkkRyXef4PKA
TRZdETSf3u6LdM+IwwPtBfsi1wfMawE6F/LS3E3dZA2Eyo4PFIzA+dMytB73OS2V
e8AT/faQWqHr85pH22VbMk5fA8cVhGzWrZeDjz2EtLErApjlB3dXdKLCpZ1ZElPT
dz/QXkp2RFmLkuNaQCI4W7duUXVrD20cYZEXLkJjhwiUBF2z0+xRVZaCZRjM4GxC
mxDjcFFHQMz/nhQe6hiYcxTw75InCGGWCyR5HaPREsMq7YTkSjtgYWslREvbkyam
pvB57cdCPRnZCvzguIuTgffRe0mRJ40DbxEw+pE+Dd1diKfQ/chib9vHQ/yWqgqK
yZCKeCNYH8ztXVHAi3YZW1u9QZQ0wsFx7lsEFJr1hzq3000pSr6cbi4CTtQwZCxV
VyP+croUANuG7LXc47gsXGlVmAf7LdBG0ebCRJVYOTlsqsElnm+LXezLkzdI8YMq
qYWJNMGWDgUStQBnNzBOVKWF/8gw6QnO9OXQTznVbfPVM3pIF2FVpPJQq/zbdK+1
wF7VZIfHpJgU9xwKPWBR4K5HFD7mqNSdrL+kWAMsN0zifaY2V1F8jeD0hzs8tZw9
LT/9b6BOTaMp9LenGrZaeXtSulzH43jJxv8J3QGT0svB8fkNpjIxUC8F1wWauhVY
MrXcrRLIePHBBO+vB/Cpx9ejW7Du214MBKrJbVEPXjI0i4vVs8h6Lpd6QLOH1/H5
g7dtm03+wAmtITjJ/dcdQHXVFtWJqGdmMYLZZXzIOG+BB3MaRNM1QUk0xjPC3vAi
5Refzm/4Yn85p/M3HUme8Im4brm/AMCXUp7Gg0T1JQu3FW63rxs6O3ImAvlFP6qA
2jR0ZTrETDLeOsGR2R/CRrgmslzNChRCfstJOXcpeKhJBMYLBr9yKRGpX17cJWYF
itK+MqjvFnIRJykV33C4KI09nrxUnR7nm9H1fctDm67Vhp2AsRH61M+iZ8bqm2h/
lfJjRjMew//xMvY1snlGgUB4I4kIsAbbLBHX9xdrUE8WjxlCVLeY8XMkPCrjRchn
HsuMAqKWxZimR9Qz+0zDPf3bH0LswUtxXgESmBBF7KugSKN85PVbubYVDpeMk9+b
O3gW9ZZZrVeKknQHBKJPSztOyr9ArcHoMBaWyQoFdiwh1x2llKg0znvX8LQPlL1R
97JQYMHbHhuxnn6q00Xso2Jz5BDEc93RfUUKciU+jWNUE2h4zyINbpg3virV8SZg
U6XFjUolb05dfC/rCWe6hunJ1kdkAXE7tLKbzrMfmXV9W/mIxElZYu9y/fclLCIa
QBNLyZF18SzP9YA0vqqkFifLJdKMeJFEZnr1SyvNsG7W/8JYL7Eq+LG4K2TwOCaj
RlXVA/wjIl8WDOHbxHxWa+kVaz22v3/DDcJn0mmf6lvLqqQvKx9otNtRrdpKdm1n
kXoFNEPXhk+i5LQLmsFdt1ObeWwT/24YsZpxvHEroo0sbXrdo4FnK5KHWLYpV6E3
Rvdof2goO9VZ6dXCwmve2WMHBiCyPIThMvpqGnXX0FEVjH551nFKAeHDVepiRhmK
Vn4C0wknqoKgpJOUSc4cCrRYw0Tj4quEQPpkEyZxtQhdNC2hF3QqXGnZOEcvuiOB
a5cZVvmUvV8SND7QRcTZ2GAyu96GGA6l59TVDv1Ijx/wA+Cj+cBBvQZBM7z25LaE
is3wm1rc6zHIlCIceckFKCOggtMtwvHU5W2mA82L0fR9Sf5X66JTNehE94UHIFz1
SV9gp++XmY35Yzs0Iv9TVU/qYgitUHphLWICCKYSMr3QqtZig8hrzFMzRf6F+Jwn
a4OYUj206vgdNwlZ/BaoI6iIrbncXH3E//v4yW0IzkERRcgeVvhUFUNjOqhqm3+M
hX1gF1apP+SPo882cg8FSA6LPl+rUUZ40hia++PvHCtNEwZWkNnxxeKRRP89eMv7
jwOoigbiKD8pJvHVlPlHXhproQnAtIsmwUoMtsenc9kbRgP0GGxG8Ulf5QksDVmv
hFw2+L/n5CD/AYADxu3XNi39Y6TZxaE8ubrP7UixsWiF4xpXuOZUcqWZC30kfubF
vF/tPAIkBdnwWVvFuhS8s6gZU32jSz5qmEOmCW9tcAjwMX92kOgZ7xrRfvwpgUla
vC+NAeesagBiKo8zleeF0kj6q+MIH9Hzc8tcSYPTD7/HKeMerBT57As7ZeQErWFf
q6Pd5gTrC8j4n+VeUgrUwdy9+h33smEi/3W9auRwXD+toaFp441SPXPO0MZB3vSP
4Jjk2JrWqbd61/ScSYV6CGwXeWTyTnh3ck8Ecg/YnzXE3maqQ5D2djqrcCaK4hJw
Je1t4Uo7LI2NPXDcIRh5eYSmxK7SRTyeObCH5sETwqgVpbE0Lwc+zyuqI7iiaeam
IppurViTp5oFET2/NZX5knmmfHDjKUI5K9NiQs2Quw6r/Qv936dTMoOb2WzhF2bD
0CIrQspi8Xk4oxIa75p72f2D5hAEDOFJNBU931ZsiqMppz4L01gqFNBTD+uLA2ti
QzHUpCv5HxHN+KaC51NgjAaKUKiPYPyhmxok4izTZO5l6adrtKVuksD/XfRBCguR
4fwGHFECXnjF0aTrsfOY2OQIXqFnwinPl2bQFLD50BZ3qq01fUt4C2xSgxhr/bKV
OW5Q4yN6I3iUNH5W+gK3hK+gD50O4wdOYxC0ilL+dWkKvly1F6Q1ABCQ+mZ6GUiN
iYgWWG/0ihu2nzF0aD2RvRDuotzJMcx3v+xzl0kofXtWEqdHWqEcJOC4VP/iYkzo
+R1CKDdL1ql5hYAnrhqPfrW0ZQluRQ7nF+aa7M1JtN7T6wbA/xlFKjCt9jlo6yZs
J3s/tV8p4txrf0AXeS+lZsIYtk407+SQLoNmSgh54vdE7ASDFtH+qjQuWiEUDzPy
oE1KajGadLF6DA98LyNJ7uFX/gLMG3XLz/iY+GJVZ4Hj1sdAhSpg/DhN0Asaog/I
Rd9odfmsDlxW87nP1viusV0uF1LTrp6CujVEGsxR/8JGOKnrv0p7NZzdfLFErlkV
vOyTohFOVXo5V/b5x3pzuD9/jQBU4RQxVPLD9tPH3DNIW1YaeLyg+FYCwCMUMseq
3mh3D78LsahoZFYwMe4b5v2BYGYS2CRHsoNSGRXl7UG1Te3TlLQBUrJBpbOrtnTU
mF6wcV5tAeJ8kdEw+iRmZ2qQCACSzCZixQO3qx5vxjXI+Fue7UVH+sz6ozwVmWkM
4svtDcQ+yw7I5eWStHBpceNTqAz99WB+te9UVJq+sE19BV43kziPc2ongDzAKSd4
HXyemqEJFXsaWKS+5FKWZxzkYi+PXYfMHC+1Zr6tEILGaO+2s+lL9HVZMSfG6131
rO2NBeW4HusWsdkwCsTQcnDEcv6GnhKIoAg8E5gTIRSUD1gu37A3r3srGescKnZp
iSmgR2sOADjUReI3xNRj9HENBkfq2cWlfj9/PBOul76b9c619QioxDHhDqz+6LXF
+gcG2sF+U38LurkCgMgyeyMRaYUTLhZXsP6Ogx0Ij5Gx5yGNEsDkjh7SaqvLOSog
71/bJ+4al49hN9naGxwW/IeFN024NZf948rz/hgKZmnxvK5FA7vTKx54Lndr09MK
ZdhpWix9V3/JoC6YRHLlaVQErDBgvcob6zibGrxgWb5a2Y3Usbfr0rHsSLOS6uNS
7rQLae+CVvbMJPccLp1OH3Pdn81ZS7CJfFxBB7A5DjjRA0lUddcgg34M4nURA5/B
VYIK7qYla81FAWrDxVK0Q4YLTvsixGD+4EGtvQwyP4SHjVPzWOavMDNfN43Pcri5
2twKdu4KD2mtnfkrQONyXrd7eyE7vS/yAD5OS8rKrXVpSUTapZyWXsQeSDP8rL/J
og7VB6zsJniBpDjq/0DPUXlEHTjk9JdlPInBXOicHhH7Q/Fyd1NsX4xncWgoz3bz
84AkGtrbaGKlYm3cqiJsVpwnGQZkaZlXEINDnjccO9O5O1ydlNVMWThDXQ2ZUu1o
KzngUyZBmk6ggBF3ju60uWweECP3q3apX90n+4o5YUVF7nnqb6Wnf5LYv4BwLC5f
FXc6FjWyGwSmJccOxS1Dgaucjk/x//Wbj+DmFczOSgcLZusec2A8JAx0fn27k6G3
YECNBDNhamMLI2tzprUb1WsHEhvwrWCvUGG7Cb9nWsOeaKwecLNVzNMPUThd9PqE
brxRRIv5pWUnoTf9e3STIZezJIlC6rMAJn+xlz+QiNvonDv0NdtxZEQ5a/3RoKB9
QwCftxSTcE2LjiNqEPEQzSURYxBdB7cPzkQ5uwGFgN8BjSLCJruCQDSgyMlKCQRk
IUrKPPs+ErX98YW0iHr3vH0NaKGz8pYXkR7bDBZ18LIjqRdo7B1IHo68pYSaPYwD
E9ZusBgKhc+xRo0kLpKdAhKRIVEFFh0/D0UyrVPhC7+DMPcYYhZmI5EAGjw7YScg
N1zzueW2bkPpb//420TV/Km1fFel7EyDHVl2bFHTmR28ZJgtxaJGTGiJPdkxPdgi
8SWNAI53hQC7quxFzCkHPouQvKUp9y7X6t6do30tfd6t3ZZLMfEuzgQpumSE64q+
LVDO0Dx+5bjGsFLKOa4tmbqqRTCv8Xiz2/cxGd7pbtJer91Qw4YrkZ1v0WZl4kwX
c0w/06/AiRz6soGq2RmzfH0/PDp7ksdRt1kKR98+cjmN0843Wc7N/HsLDIJ1vVEW
9RaoX7H9CS4NYpBBM7H6SUjtFCwBNhqkuSXTlPMjEVJxEfk8Yp1O7Y99CnKXtTE3
CI5hLIjT1EeIjH1QZ0d55fw1MLl3mEhEXN5p2PgsNFeaK5LApzSTKt0ie6Eqggla
C07A9KJ1XmGuH6mIEfezcA2RLTVHuj+82wcbNtaVgTM94p/17vUauPBQJW8u9uus
3U27CTvK0ks2cEM/EanNvjHXQMtMBxAMeezKMCX29cxbycUbjB2s28ijJ6mxIIR7
D+6GNDsRFXtN/WaP5vCbhFDfVrKD5uTtooR+nJ7ssYr91RftdtXU2mIRoDtuFnE9
SAi17w4mmnWIRwqxMdVjD+SOyBD2QZdhGjqSEmaOgmVXaS4wKyTKa35L3ye8lfUB
D69YfU3h2890/1Z1I5iYbR9P+F60ukATV9s9Qtxwd4/DupZ8s4C8Bx4YebDrQ1x5
u7np0PJxGw1B8F3WnMOIFuH76/o59wLehabaF6CjdKPaiMTLCBTBs0Vlp54Tzh5m
H+dS5F+78fxG82EzY8ZM8SfggFyVJFe7e6YC/uVoRF7Xn5YFnTBNVfwwMwL4U+ey
Wjy3A5Lf1iK1VoMeAuYdV1K8/PMHGJQdn7vlTeaUtq07omTfJ/tNXQOgLh8IPlv/
fYk1Pw2rZ7FU7/tXlAn11NQwNRO739ByU8EHYTX1z6S8rMcWetcpwD7DDCwz1lyf
MPsW1wt3StzaG3Oi7KefAfrHejdu1+qT44jrNC2MlwM3cBiAk1s8PEHvW+DhidKa
wqLTatkCdoJAKNVYy8XFBWuGYW+iPvw2wWUlUHCnWCXRY/+JjBMzsUoHE6Gaezfm
o0RBkRMop2CL2+j4JX4IIWh1Nx/2ytFui6hNjdmVEIo53p0yrnQ1PDC38eU85cKc
3xOWTW+J4lVlz+LxZedzFGKDdXmN9LGpeDVyjKrjl8G1cZzs2bAIBK+8yQZEOa/h
aSM6bbHCYmumwT8116gius3HB7ZIlgqbB077dhZ3j7Ybl8Y0XDwWe3QHCMsDRAm/
qOSTPrFXbjpnISwX306x7f50SXC3BTQsWv0uWPRGVMcT9y9if3AqFZ6ZbUL1o0F6
zVkOT0Fvukw+9nOcLJGZkheTZz05JLHjfX8ErdzC0YOYTlfMVL0ihXaIgzv0rHlH
U1TVSkmxxlQvbN35cT/p5CrqSztb+E0nQ3XAhQvHISu/mHzIM8iqk3gHgWyagbZ5
32ckdPRrMvY78bXrii/6Pmu28oYzfjrxrnnK4qJo2l/Tc0B6s07hAmMypzWJwNoi
FUvNKPuQQetG7ojrluZ+GHcS4OzelpQ/2g1Jao1hvyN8x5GXbIaVtVIaHFJZgteo
VdmGP5qx7cPB4QIY7PKyuIBsp8hS7OWX46yn+vc30ePdl0wINAxgqCM9GSUrn+rg
h/gXwfdzm38bT0kmgB/3cdYmJX+rOni3AQ/W7FZrtgBGsQ03tN7dGQC8GNoEiZy6
feM6WTTEa0WRMcV1LcbynTjWKP+691X1ZAzUc1W64OTq5B0X2uYKlpLkBGkyDAY4
Sp1d4MPbskX+aAq4D0eWY0Lda9V1c42iOGY7ZmJH4ZVEbrwndlP9pCtcBdLf5+6g
em6RrKuuj3Lz9+nx6QTmPXDirdKjMMBSt9+EzhtTkx/V+v3oZeQMWpBwYVXoYUo6
wB2yK3KfFUvAysPqcutcPTr00MgdFJPT8dxt7T4NR6xZ/Ql+cBwpoxbO5Bu+zSus
nFCM38r/z+OEg6V3FmwSES2PVAjzDotZk9JMUm2ASNqWwttcp53pxVrq2X4sPEXd
BlvvOfvMPvfZ6tS2ePsRFO+foRRAzPn52XdN4iNHo+PoysABVdAepvi2tG6KXTdh
NtUMDUUXBPiXpywsJVqxf7juOmnfZSIT0kSLPO8njxegIjMb+qIgEH1YyPII8lGX
XL7LzxBHHkg+14+4C0lYgU205KJq10uVOfcRQgXnM94JtxF+syl1LHMIHm35I6bB
YYMZlTXSctviUCgvofBs4BB7X5e3DDF/Tizb1H97vmmJJR1fxNu9Cq3G4jG3E9rq
Dgk+7ofzT2l7HHXIBwKdA7whDYQftVPZdd0sqnifwUsEEEh/1RYVKeLpkUL71DH6
hJCLvC8A3dkyQmNH1H8SSuS/+mDGbJL4sWp1sAsI6ZKSLfYp842+/zvqg4vnmmvd
9Mi8FFkb54lJvU2h/qmFal/RfJIYBPpkJBh03weZjKK6jQc0BnbHyLJqrKzzlkaA
vkwdh8Yd08/iXrH7pmiJXeedmJ0zSfdSeAuV+2I5+svy4Yv1uLAkoqDblCREmcg/
hwNYfMq/PoFCnue1lrgduqyz/4pPU8CNOkIPSlImfGnmYxZwbkL4ZeopcHtXqeq2
tnoYKYGBgN+iPgNsWp4/cQ3X2iNzxUvhOEtIereM3LvhcdjJ19/5CKZocimQdPPb
XzM1Yhm+CojN5uwmW4EEuHGttfBdm04WoxzYIt5DxO0E3XodxkWYiHWdpHGkt0Dp
QoZ0k+PQeWRpVe5fLPuQ1/5TxTeRzG91WNGhKE5E+qaoSfR1pzQSFk/P748agbwd
4S+6KPwokYUPgoib+vzp4Icdx+vYLIQ62ULijuFruvTdSzMeYBz/UUboyQ7AUV6m
KRkbrdXwZyzMVPvh0Ui1zCHbmZBSnacj5q+RdVULOVMy4EGegUtd9rGEAAnWSfrq
Ibqf8XyWDwDYFzmaWfRu7LXzfSX2UIxqD2ccSn3ie4OGoGZ1vLUhkeY93NgtCP+g
+QlNP7ckp/kPRdSg7VA98SpKtroNwUAm/iVSqWy9+Vuu2z4xDKTUghMZCTQm7OAv
wSg4elojP0dychf6P+opae03PkYDDzSNq5DpBwV2BN9JoV7Nk5IGlD4gYcq1gN6e
BP1zEZ8lvp+6jFahrlAkOx9UdtqpuafKjC+vtyfGtDhGzYKVifFVlmmFB2Jz73hn
ZbngWqCaLANH8t9Xudycd1tQzsc36Y4bxfY+2qnB7K4kpNC1uNqzGZ5811SwKCJw
exQkg4alACJMKtzQW8x3jC9iMMgi173U8eHx6h1EXBqWFmJGpZL4dLKPMIQWd4ki
bcyUyk7rExUjmB6Vt2VjQhnSibCwQjeJ6hegn7dAV5N6pe6WjUvErkcVprHzAwKC
OXCO5eZ3OGRG2FU4sfrzFYboBC1WNbOqp2wirIFCcmigwVgcfHXsEx8KUgYizfD7
Q2tBMp1Irjx5K4JWAm+Kn9jbVGErrkxlrX3x7jM7RmWuL+wkozkiWVcjZHeYuyHS
T3Ki1i5Fk4vOlpKXw7ec7x7ed4fwKK0F01PHj/DF03WY18dkgFOlUdJyiSYZmqcN
RJ/ZtENQ9IGUNIKPDJOdY+bV5/v5806KoJWKwDBG9yKPnm1CO7L2er/IqoBovYuA
w1gxW0HUOIjES5kXtlrbycr5wBD9EmilRGTPit15n0keT10XOYgYX3qjWpvrXBbV
pZR6puuiVE6yQUhtg1gDJ0wu0Nb0NldTbex/ZtR0TAmHV2WpQv1S2xEmuDZDl8NS
vutP4oe1teZT8Oez2+yvCaHq3AbNVZ4e0++h6JWFUbAaNtLd9I19s0LFGh5KoUSd
4pOSPfaL/gN7LYn4phavtpaeBCNJ25yTI3jBLO9bVsb6RO0TFtX8NEKHFnjY0oXw
fv369nBwY/b0ACOgo6plcZq1H0wUvLjj/vM4+Kn4IPGTRjTgSk3XClqUhCPYQqpN
KJ6Tu4GmWjz87a6WB5yK7W0jmM6A4IBJ4hVqvzX0tQV9EjCslzuu9XGmoAlo/+ur
uUPlIlcfiFBaaR3uT7dO7ooW/Cg4x6rqe2mSBkNzhSHQN05/zWTooLBCpbze6/lH
jrB6JhBo7KrdS866KwlZTpFaV7VD5ijdJ4SaBsVh7rjKC6nz6m2jj9UUMfQlxu4p
NmxpbZ6jwQSoe87wR5en9BBXWhQLuTA06YB4M0XRKLACAU8nX9ir9V38s/Wk3Krr
jt8jk5E9iEzxrFJ9wLi2E7Wg0OAng3Az62Yo2EnuIshqabXSFv3lyDglzJB1bTxz
udKXJQq1c0goGyRiBymyHdqopGIseIhlHDFZEhqWGDkI/AtAp8aUv0bOeItNpqqz
yXDsgyqno0NfpPITpFYWvNFn7/ZdeaFJVpTDwtgb2+N3gU9MptYByBVo8liwK38H
4WA4E4+npWmwr0VoLJVwaOUCtNgOjHMm6aCMsw02JxqczgKb5Ygi4iYKsuNuqvDY
FMr6DN1x10cYXkwkD9VrpLR2Rkfu3b+NwQHyIVkIoSS+ooefCjvLPLKc4DX+nDqH
Q5v6tbqJLc1gHiWGKYUGRyKKQs0+tM1DegbzVIDbNTIYf5iZfoNIpx4bTwAV0T9w
M0cDEFPp/9t9inQxZ2i4Vw9p+wAosQG3ymbO0ucC5z475UebXAj+xl2gpfZmcUm+
k0v2yJ5GI8awMhAo7QCkQ/rExsJg0qcW7ifsZt3T4kaSmEupupmlpTGGS9Y9PzyF
XXrbNg0cKCN4vhSrdIqeJMxUuxDWDUptUssIE/yPYoeNprI8QmGBKJEPiTbfJtGd
utbo1hA4/x8TdR9pni/eF5bCXvyObo+0sYxL4sR1papxHm9M8PdjEGDozccytsJx
bDDoS2pfJYALdEBkPlhI8lUVAgkpC3OSTvYCZ9W+NPc27vNxq4rNFsQKrjy6zFKj
ducNTLo2BKpkekvYe4KaLd9NBHN7iZvAyOCtnCu8J67FnfNL3qNVfAQvipnHUo4x
11qnZR7kJyNVaYG1goX1NDfPqGA9p7rsFpElwrjP+h040asU04m2aTFO9mTsDzJB
bsP58uokHn98VSt9phVFtXg6T3jBNtyQSYOgFlVAhLMCXsK76ZdJrW5Pqc0JCpFM
uCX2ikJGF9BL0YSR+FjpU9hLr79HNHzDVGmNl+Rtr0G1oAUsrzlcuuD7Yj4yvO3m
rk4XqjTWrXj5cKqoe1Sa4JqvdiPI+Z1ovzHNs7PIdBMHmZLjcY7UEm+S3Cl2bVYn
ifGIQ0DF4sFOhm3muH7rKmiA2UxwF7S590TrBfdto0gUBpKWzJiYC2aSlUIwN5t0
UA7qVHGL4ZyudC/KYLQf8U4kVu0+0TMkUkjgnwBTXKtTka3BXxfS77fl+1GWtmUB
MllWesRcUUMCA3HC/gm2oct/9HqeS3rwi/k4Ui4O3FJImcVbHJQCDIad++GMmd1s
yKdrOWffZ4AIW63J3jtORTxl+2z29ZvbJl12PhbxThFzgqB+OzWaLPpte6b4jfwB
ZvRlczLrqWAPuRn8l8qnCSxEtsnyGxA+LiY/oblIOa2hAPneZX4Lst+0RPFvPxJg
rM4uppjE2gJQSRK49jsZjaTu1oX+RLKkkJHQWeTghFScX2WbdG6U7b/q0wpCTLYy
a9wFuboIl5VBg6EK+Fy2K8S5N5Jeg5HJbeMdgccQVXyGPU1RIz8G0j5cbrECJzBg
R14XkW5FdcT9E8Epeljb+PiiVNZTdA+oStvhHYH4c2dneyARqCisRGJS09lLtYAa
IWO37UChKKdSrvzldDGrtfEuHNnk/q3A1Lx0jzfOgxjWkdz7bOjLSdLW/OO5C6R9
q/B5HjbhwLesCuHiKvQQpZrLlAZeaDXM3v+EjVU4F+Dsz5rCelBx5QT6yI1QG8lf
umxilRQeENVwwOrbdKjZGg42KcMcZTS7BzsEDfIgGmA7USv6JWNprPLuwVFrodbQ
djob28LPo5d1SLixT3rcfkOrVQZTvh2o7A0eQwzrlC18FUI3sOTKUdhEDbUq7L8+
dM3ftzXPNDJiI3QfMTg1NkCCu3nAPuraGmXZE8kkynkpkJXs92YVS9JtrdAG0t6p
hASY0hdD1yRjXM27ihuSoRaf2EWh/PpyD91OC/4uORV1sktZ5P7d4XbQrsYhHJv8
ImoHXDYObykEwx9j/99+AlH151zsX+/f7k533Q47Hg1f6+Fyg2bKpfkE0I97dHiE
5b3QNfCq8XiRH6zIKPObmASRsDuUnXOoxpxptWwp+Ub/LqPmoqdAqbR01My8QBtr
DALKTljghqyphnYK1irY3yHVjBWuia8plNYGch46DPqcHP7L9IVxBrZqeQ0tQjZI
JxDthui5YawS3KkSArCIXJN7clwQl2YADWyRvJlDyDZ47TMFiTVfw7A9L6R5KUpe
sAKaKUMdu3no0UKvzcudJDchn+fX3bnOFqLXPUCNkUiWlEoY8BBLRKfcei5WMz4k
zd3HpUvqj2qJXWNmkGTXsu20LtQMffLFbxbRofht8POzxNqmphY6NPzI+HbF5lEC
TB0+gPiqSH5TnnG6/gOPKEOb+ynjagVAKSVw48r7vrzP/EnnahcSbH9xSC5H0/E9
4SGxnwyWqd6iKqt6ZjH2YtYoGY6dfs7M9COkssc6Xgh2h/M7cDBMnaSE0HJW28er
EXdHuxW0FnXlahcDCQFSx6RDZsjFspAftd5XrAwU9xz8zp2vuz/RYDT78vEyfarc
odOj7rqu5TWLopY12BjwcLQm/9bqbz8hiJl9H9fTe+/X3wCfdCfAYn1+FoEnWQKV
mw84lbMZVvQ9OrrNJ4obFfN4Gdj8J7awH4wmWMDsaWuyBjRuJHQ0K3S2nsgmpf6n
wIcKl/aTL4JMrFfOX//reyJih92Zj7KjiePQC1AC3F4rdD22IUgcIDwdpBqKSSSR
QL/tw5m6198QahXwKlAQEpiHPz6OwMN+TExJhZ+o9dUyRYAUJyicg/8NKZKI2SnN
rrtSOZeO+bLNw978gX9vYIiMPTpI5IYT1/T+SOjWE3qErX+pUJglL/h0r4A+TXyG
BsypQvMWjRERYE1pkavxE6A92JEOQ+sQVndlZChIvKL/7h4hNjk1DWijAi/ePJty
ujOwki1STh4lagBwJA2eoKhNLLr8rTcVeRHXPg+XOPYxUCCZUDPJTXN1vBL2+76d
x7ztoMbKHw6fRJ+dJo9A3epxxX/VTQFZD9UznJX/czs/8Nsdycjqag9Bvrd8u9Kt
QbtbR+HkreRepYLTJhBzmra+Yv4c2io4de5ymLu0ja5y7Wvyzu++tZDQ/8CrhaU6
I2saNsQpTM171PjdQr0daqPfeIxK+KCy9qW/p7O9wi5X+6kcD7umfjYX86MW9Ieb
tZKgkE88rkhs3X2vATHD9U+V5IAaR35qb4poN3CDkBNQkX/IeDmcmskfrFb8dRKm
7jF1fY7H84ojntKbKMhSBBALm3Q4XxRnu6GGVaGBDsy3zkvCY1mNuRi9i45ZMQiq
pdwB40s4oMAMOkoO/3ye3/imSP7xEUc0m7SPNd7m3C2KG3k5LPUfluzaJRjIqPQD
2eE3zxatBymOGTDsFbmUpGikxyWsoDwIfNlkPV9aY1ewbZJcOQxRnM12kGlqICj+
prhPNFT72D+GLm0V6BJrIbBbyYqiXhC0mJkgFGIbMjVbSIKCU3+QEDpDdMLRr/1d
Wx5khfuo/5VgkGkntoLVy6HLIijIn4cY5bn7KgyxyFAhS9IivrSm934ihGutxuHm
k9bEDoVOZdQ/WpAuPU5dBBf3iaCK8CARd5UgYkD49v5wwgqYb1coG86QkOhR763V
A1qw+gGvDLXgfF7ZSP2qxvb0eFht+kTWqjlwr7G+J5xYtO5zTG7iwfB6Rp7uSFC2
s4Uh9Kpfg8a5ywKUqXy4+A6c/xhAJOm35UCkzs2jANWFMcPxfuFnRZdiHfPsf66U
SUOpAP6id5r2Pe2oXcUGkgiCSMzweUxIkvXRr9tc35AVw+KpFOjUbSw7/+rDe5mo
rZkL5A6jgBbgPGhGdFHYEE5Yb+Kz4IbyI9uBVGnGMC49RZo1QzzgGz9hlnD5Eifg
RcUHI+mGt1RTmd9VaTZvmwge6YAaKASrVoacvBuq0+1ouI956PQgA9jznBznP88Z
nOfmp+X5kFw7KFMWo5RgeqzltLsDRaL2vO2fCFsZklcbBtp1eMHfzkG/TcjXPX+R
zqeymwHs6QDy3Vm7cPx7s8NOtPYj5y8qPWX6KrNyU6D5WrcvhasZlOaF+0WT7z6+
hbcZ6uDbsxJz7Vgl7JhlKeghc/k2HR2E2vEnKxW/c1TwxeYcjaseRaVm9YB54DVn
FEK/qQtaCjhmvBu9CKNCR/NoIRUN7BhCwWdYuF5j9AvHPU9YKvK2WF9I/hPfA4U7
uarDEQ3fQp5EfE+1LOjVPeCViB9M2Q+kSv7LN//Xgqi7kSHXFsoslydxx16x5k1s
TdgBVuFGa9ypdoy8YsE4e/IbwtWYdm7r2lTZiPvgJGTOR0vpTs3aAgYHwhBq6FiA
Zh4uH8v2f5t9wgJjeivRlS5/GbY/KezUR8U4a1+bC/2VoqLLK4TtHGwQuvmaKB+y
7peKYd64BpCbv9b1utCDiOmdZ0WikRYICtFxWOHI4ggfTXh5zdEYaK7to4NPcuxL
J3m7n0es+NMKLAyLl6qPJaytbT5BczhWl8Pd8EIHl9kS4TLjY8qoIIGEhFiZz278
QxmBoA6bBPsPO/3BfX76DHEYP/CaSdPaMRJtIEO3yHsmWqvJOhCcUo6P0h96LUVx
hOcOEXptUfFwaN9pXMDzU9zu+LL9XlqJFaUmH1fhlrWnXRAWUSxJmD7J3zcOLJuG
PgOPg9rScuWqrFeEDyHjSIVcJIdFo1hvPhFX1ABOYdBhA7MrtK9FWzVOgNCuVfAY
6Qu/4GZEHr4bTul7Bod8fyEU4UaqLzk9RGkVJ/9aB+g0KIJmYjqYMAcwmWKbzkxG
cHBYiDPzxPI8ru/gBRljaNT9wbJVf+gkmlJ1q82xmkqcNFcLZjXfptIvqJqyrdKg
hK+Jdw9n8/CMlRzrMpd0lzcMnEIY8ZA6pIweNKTcNru4vgHM50ZTISe2f5Q02Dq3
sBTvc4lp95oj6FSd30XjpoTqZ3zfXX4CJDdK93gMoYZJ9Xq3UVaPoTtsdIfqXnff
d6ErRhvsGF0sJyF9c3DWhCOVnDWU20t8Q2YOvUk7X6cSnUHBlaJMQ1XiYL2PJJ6F
UYQ1V1F3dU2sxL2whj+eIEfetaJHn73I2KO6h7Kzzzq2GhqBFA5NijrhDchE+BYJ
hDylMQHkm9ZawhA1Oyevr18vvPwyo+UN6jnIPTIBSH1zgVM+Hs/m9Ji/fnA8qqVO
UFw/ddu3BkHv71bC7ScdJ3aN9XL470iDFxBQbFS2F9RC1Xtk6LiH1PMT6e5geO92
W2Zl2W3Kkx2xnkAzxO8Ge4HIA2p90qIcoqPNBQCW/wZyqWmQxmV4Nhk5ynuo5OUE
dhWNC7Kabd0lDVfrvDtoLKhbfWQ8C2BfccJIlTdfIu/D+WXV/62AurpIJOmc+XHe
K+aIfCSkCaI0lr2GKVYOXChNoqR45fpHdtrqrCNoI2mVbGdXVtEXQrIHIOvnCEQG
ugq2R9KdIUL4g3efScrOCUYq9KG+URuvZVNewkTZ2tGXZla+E/sRK/vd5c8ygciH
dXWDXuFpNc1fZcOSzOphjN6WnnFaYQCkb8zAalFTwNnLMFxkAkQzRPVmmaZ6S42W
Vgk59yTyTFVkO9rnRC8k/HruaB7hu1576tNB1nTMVCiEN/4BOoZzZCOK0cl0NBZa
c3/a8shZ4PKH62X0zkYCKw06jWPOM7smrwY7d8Yj7NQxx9Tjh2eE6PxGwxt0qLPW
amIt8/ZmTf2Wn/NY6aubpwPtzLnVsqP7gsBR5v3hZs9OoOqrvdPMWMinT2B0mUCx
gOgrVWY+/V0JhdznBGkYRBcWqPNg59/9cPI96//0XZy8ulODuMCJq4qBAY8URIZz
Ts60qtpPUnPBTbMRTUHCe/+OQGNNvLy8BenVGNl8xE7idqhVDILR1SoYEWNKZ3KV
US8RtXPbpfBSMuvrPsyz/18xHbeJJpEom992GRNn9HlIJ4XHqfmXrNpZxhCcqE8Y
agrOSH2PvENSzJB3ejZQrj+/5UpvQpuvE1TuiNM7LS+KZ7/F5OMkfTlkFx1MK5Ps
zF0m0xF4HKmbC8UGeVnNiKu6ym8UspjT6mLzRg/cSLnZKAS0ESyRkzNzZPwZqiV/
x0VyewNJ3t1eJy1eC8V4ZlNaK1KgP0+0kU1WchmG64B+5msd3Nti+mtiunYY29r1
E39sEUi3LMyL1F05jER9ddZBEZ63TPuAVz1ilmgX5ixAm0Ws5myYia7OrGA6lVNE
7AwEmDLguEavoFeRYKW84UhdRlovWzf9xMx8t+dLL6AaFB39pyKWXr4QErXyxOSV
0X2wKDKxKJMPztBchknjxlUYLRvtNzR7+0R3bJpCB7wz1IqyA4HFKnegE/qG7iLL
2w1qjqzpLh8Ao4+XgGvXTbP2gXkuv6m1NUDHMwKPJ+DYduW/eg5h+69VEQWN/8A1
vCK+dZiOZvILr1QmDiwY+MZvY90c8gC/wXqvj3NZUKfhFr1bsPM/ImvN/VBC91aA
yREJIQUVUmjHkxejC/TtydQ5em4ABNoA30Vx2bbdAN0ANiVVTuNOD6jxD80GMqBW
v00bPYsOGG72MRQMWZKlstRXbhC0pI9HhPfGDpqriNf6nJbVFjL1JXpSAhGe93S+
X6ZDIGjLyJwu+hP3UFnPkoLMgM13LSr5grv92KLXJEag/6vtELpYZbbfvrG5wMtV
anDKrpFdhoFE1eGGyOCi/hlKf5O56HJKQxE5FnTGFXuisXvPsguiQVMrJI36gbyZ
RoBvh5P03MeHmnHoR6e7PMfpD12IJcE7JhDRsB7GilF6KGJb+s3oobiDkaZOr9Al
SYFuAvU5AwtF/pUwVFh251h7DU9sdnmwzd48WCl0cX9uIfsNnJb0KsXFOBpZSNKJ
XlTHIeCpezGNuyiKl/YrC9KA+A7YaE7ybCldoHYun7ZY5ZpWgQepSXk14fVHXm9k
r8W/VHuCzjDUaCpiC1ssqwkkwKNE4PRX8dOIrW5PzblOol3dtz0BTniiq/rhTNIq
f1L/AcBhwX4ikQ+GcHO5W2SzFL2BJbMfxy7woEApCpomYvSWCXzdYzVfOzFeWaU4
H3+nzxLDe4MC5uO94unkW59epMAM93xhZe7mIubkPUkzdL61vLZDhvxJVUhmVKzF
ULcPBMB1mVpLwJ2ZA5tTKSg+Yo0+LKrKQWTGUSGVJcW0P15p0CaweYGlPP4b5MTi
59EVKv6h94ZMlETuL46ifpBPVGOdCfWwAbHWjxCdKcOxl9zlfNB9Rpb9PfAMqbaL
ljuhr8J8Daaw5LYqAIVyL5DdYQUZdQ6NSmjjOXQGy4olxYdh0bm4iHwH3T3IFXxh
R8uQLpehX1Ni/BKoJuOgAFmw6IcXffonCBCv9qg51FO+aAGSMQUd7gsDmaAkpP0G
MVLyC1UyiDfTNmpnquNdR2gOYADRiBi+kcAapk3tJr0h4E0pZ2GfYzxe4sJP+/3n
s1iSOiC/Tck2aRPSTg7CMRrDUAW4+0YxbusBRzC/jZlI4DgRkvGVgKdmT7fONorD
NMSiLDEL3semP1qxlrXp+9pEffjDLlnI3biOsQQNxt5LgbF8dtvaKaY80TiIAyqJ
xFRD3sejhxNKJgzxm8Y4aszM3g2MMbs5MMlEFs5SuWHmODWFv/pZj4yQ5FvgFzEZ
n3GIkBsUhWZJTIJvwdSl2YmqF9zM95rnkiSJ2TFhhTk0z4hQWyGMnLPecuPF7e71
sxLyZGYhltHt6Ayzanm6bQmKzy/LsQf9jDRomlLuQN9eh/BdqRW88QfVAPYdtTJs
Q1sGvx9/TXKQajQ4KTzDXM1EtYwIs+4Mb5yqieUWH8VMQHKvPPwKS3AvSaVW3s6B
Phu0mHNusB9MmR8js3ddACJbBeGCgip8dlK5QzIaf8E9I3O8jZ7xeE6a+kmLHWxS
CKG+YRsq2gfLZAa6rbgvcjcL/bgQm/3BRwgA+rJDd1jrxnFT6CJR5DQauGcRyPmL
Xl8Uryoej733oKijNgZJnJZS6xybj6dbklZTXhW7ukh5hsqLcFpx5bcQ5ndLqEGO
S/H5yKsvx3MrRTYPqjt/bs2yUH15+XLveYyWUpxC8adFtphazdpwnHKnrvuikO36
2KyGR8hTOUyim635CoFcRbyv7HpsZjxX6D31YYRKjo7OTLB52p0Rj/xqkbUZWmp9
yergnhwbn+onnbCUAwHdWo/O2qixiXgqjzOXaOezdzIrPoS3eFoIvX4PJqFFoisN
Q4nX/iF97+THzUSYJJRCDX3Y+Wja1yR2JZYV05H0Jelg/6FYYJxpEwqDRWaw4PEw
Jq0z40QiFAugQxlEJUFRuFeKS9NQm0Nc8ETqR0Ae2QY6VF5w/l4rwRd5JkN6rP0L
WFW7yPJXGPizUwPudaVPYMCH4qc/Y30js18IERw225LAjhYmEMv9jS75v697VYRe
5TD5NDixia+IVVv7RYneOS8FJTfeq/K9ojekZ/BN00us+8SVwuU8vMp7JZp5+Jfz
UxxJcH4Yy9MhkBUJGMFYS6O82QYaaWmlmESuPEHL9vG00x02XoVHfyx6GFH/pUWk
b7M6ndMxcjZ55CDIPgYCnS1tuX5SyeFwsVtSclAfbBDx3XSFEdtvus0bgXYNh9Gz
MFIeOqOb+iwk801h4QtH40ReYSvS1fsOQZKQL8WNaLeFmGOgmdAlFdYjF+2Djwa0
eTNyn5a/rZRfrJgFBGPlUtpikzst24rfADQjcmT+6go9OKEzSfSw/5yjDDMfYxPs
DuZyf6K/xedZ9KmCzHVSDn66qwu6nnDmdxC8CNwAW6M4zOT8IGRLQfu7Swkm+1UV
2RZW1K7qqxCwHerqPMvOvOpABZmLS8PJoIOHkMmPEqtNdr4e748Vm62ss1EpsYSb
/T2mpqUNfFIn2unZJ7d2ePLlejHPpDYFU7E15pwo1oHvekKlOQYb3it6t8YpVg8o
YthK4E7dMek8zmOqjIFOIthFYmW/Zs3qJExoeXhe/mZzrk2OGnGGev4v4uq7CHhF
na0fi/0Kdxm/mezu9POU7gXZePiaUupZCh8TlV+t4jxbBs8ZqoEi3X9NLkX0EirL
/ralMukJTg38vWhBeQA4rg5c7HisS1oD+UeARY/lvoV5TTMhb8FJfzoL7bb5nC49
95q/zJPhflmMfZLW5OX2Nyt3FyGUDQPiVnrbAH9xhd+Rnz2rRG9R1/Bn4zHow6rv
dakE/s3pJHGrpLZR5h1XoeW7iE87hnjrLXkSg7GypG0anH/RXv+N01hmwrt84420
SRtOXIS34SxCjSJnz6XgckNV+HwMpa18VV38TF7dh6A5CMATzIULVWFOUCRp5ga8
NVDlrl9Ro9n0cI9UMY5PfWzor2QCwZaCQImdqHCqoAsiSNVXvuwplckchiRuquBI
e7u0BFe7B2Hmu/5unYV+mh9t7J2zmij3u/yLfDuYKNlOSC5/TiU8xI1LC+MoC4A+
H6RTQVH1erb8Me0g8/FsDLUjMmz4J5YpTPw/Qhv/WbgM/w/x/5uCtw1JU4GTbTl0
oM9OKxM1Ytl0NBGg09Ch40QEFLrL20qu3PNV0n+6RHgOgMaJ+u768n6ciZSD5/qA
C4Q52vkivpc6UZkMrG4fQiSgzkZ43+WnIc2Mo+4N1p3EPEGhIB+GWxBQ6pSk+TxO
JJwMO1t+QurXU7NwghwHcgzzwhEbfzQRVRkbesZyr+r/PmTCU/uhKdw/GppA2sQ7
Lv5206iBfqiQS55pAZTfMmQ6GWNYwEATbD+h4CACPAIA8whzXsbxU5rDA+U9162N
buGbdTV4EHxl9/qDTHG40nW3CthM2LzFuPiOxM9UGtCZ+Zy0y44vjW5fE/r7FFMO
ZD3KoARgJ79v4yocLp5PVKgZxjDH/SVSW5pzPj5PJQbsr+rXXc587bWkH5GrfyD2
Ie8zWYLnan3QCa1wdV6tVg6c6152d2CoBclA9Q2kzgZh7Bus0Trzb9cO4NG4xijd
MbnPyBcqa91p56xsMMjSjC9uFz9Fcu+ZvnUtdCCgBufYPaSewERlVmFOm8uMkHOV
GLl8LmhP2Vdj4+0GoQIn5t9rthzJEFWFctiQKQcGnM/xVwGzENjhwBhjWHptG3wY
ai0jDT9DhK5J3khvhgCeLWQ82l9K27/SlZyrxeJbimo6SF7nbHJ00j0JP+O4qw3j
eLkuGmU3cfSTqNDUk8hsnAAtUZGv5BdweeGiKoWb6bS3G2NtP5bhQJGpt8Ksxwnp
buMrI4E6MWL7+ESjDQp5BXs7H9wk0e9Tt3cWZ959FltA5cste1KTGViJo+Gm+1Xu
HS/2PvG34ajhQn0iDxObHKCxXEhzneUJKIJHkqdRh1Avyb5QSU2ZUddM6lHL9cr0
oQifpxxGK0k3wmYCRLXdV7SWGe/lQPKUl1hyNaT7bZZkmVRDIVuVED3E/1fujeZP
hbYgU6Ud8XG73npnDHfFJ296wGQVQWqS/3KfkokrDaRQO3Ho07RSgIP+ZcyICE4A
G5nk/HZ4LweOdcZ0tgPgjh7x4aj+4CAQptFal5vhd9XZBF87a4J8dYjInSUciCv7
NGQoyXeLBCby0AXffXEsgF1k/H8NKqsMA2BSluj72dmGHxZEMys0RHbQHmg1akNi
6oDBs6mOaETmMfNY8hEk6OZ+9yFqqETRTfQdH5BlgbrY28d6YEJhC2QMyZGjRsz3
S2QTXhiHl4tJvcpTxKqTqYgNmnQmgqgcZuoHom2WsF1eHjZ7JmoLjbqqsgNc+mMU
cVznbE61UpZZK303m1LFQBaL0wZ2IM4JqChp4sCOsSQDUDRpO/KbHxzElchZE23W
yZtS1Uv2vP8Yci7B47nZBUAf8y0rSZmiZ0uJLgvEGRcNy7Z4Xe0HxBRsjn7LQ6MV
o5yAyYp3APZN5lwnMJHJ7KI01XXf66DZQmIN5WDGxhatyehQ01ntLALpPS6seM0B
cfpGEJRC5qtAlc+Dr2K100QZMZJCU4ft4lJ0A4bUjwBAAan3/sqBhCUrHq+wmCBX
x9rx2zHjMYXf4l5vp+Q4elbHVJrEzifbnyvrmJvprIlDdmnMOxQnWkFuN8iQyX/5
Pn6fQBn5zPHv1/75psLNA11bWtR7l4OnWt0ZA3Jknibay26LofGjBH+kfgq8Csp1
QLFpCgGeGanzdqgRytD5cXKe/EKl/w1L3uJuysJtx4iRUmmORs5pNlak4ycdoMtS
0Zht0QbkBwOGRLsobPYzLpt8biIlgdkbUs2Y43SfZXyX55wcJO7c8O/Y4r02VrVn
IqL01ZNr7FEU0/FMDzmB8NT+spp1s8H41nJEjK1OW1ow8/j3JJEQ7q25YOIm9363
iRs8cpoGEPUICY2oro2kua7jZKA3ewsR+UMWkV1QcHA11WN1N81H2J0y5rvcoqST
Rrn9DWBrjNCxzIEM/7nzSjAQccvPJ5SWChDIJpXAWdKbPaDkA1JYYBXnY74ZYqEO
zcdDbR/dybW1ZWQD/M4eH9fGoaCVm5UTHYyNA+K68pT3KWiqtiZQ638v+FPmHuER
b5V+BYlSsu6TQMbHjE4ix1hrZI7ShkZC1TgM4AdrE9GIgo4UM8x8weFqZJC/eq6v
Amvn2ya9DJ5NwrN3QeZb8ClQjplSCzutLNix/u9NUqoKLipsnX2aN4pVjSLwPbzz
gaTcDBvGB2pIitLyUYXORrvbnATpM/EWea/iAQwksPm7TKwm9ZtgNNKQUFXBNV/X
dObZMNQbBNMgtdVELh270By7QFQIYH+62oOZ6LMTJ06Adtz34d7HhcAe1PpKfd2N
wpsncUqavODJOXquRlPq1HH56kgfykap0yBhB96FSEyZEpKyjhKciaWvne/9bza6
/epCSTuEYakyzJ0r347Bgt3xNzSDWl7ZVVVDwHaLrl/Mc2KfkH/hzl/pQJZx7IL4
3RD0xT2TVtxypxdyfxNLVAImoizrZ3zGaG51fDcgSLsgwcnrPq4TfaRWnCTFvXeJ
kEN+xdw6snVsY3nMruW9AYJZJfTNzCGoA/Xdev4IwpWtcYoXuF7NUdtUvJ5VFYT9
AkMMVa+jaZNrl9f/6hUXElfl8K3g34J3kDhtiSosSCqRgAsbLt/2rGYRueVMcfXz
Cik1ooKrOgovh8leHfkswDNmfV5t57k4dqT18uww/Fuw1TQE/L6UB+xdZHP/dns7
qrKbtYTRSa0M9lsE3/7vM08TGJ3gNXHFOuXpbantV556ZHiXIyeUhWaawmUVPVmW
Zu1KRZ4Hs70utm7y5MYGiJdVVqoAxz7oZXKKecRFxoM+xYlkEnv+L6Xz0xuGfDAF
EBeySmxDA5+wKHZRZqZwjiMIQXBafkqXPsYam8VGKlf0ZJYNJaboxq5KBpRDfa7r
5/nOT5ihI8Ibz0b4kJcWLGsFODG6CEWFBabOYoal+8uLqKjmJVFBKM4DLIPzfTph
O2pR3X8OlLnbNX5BOlLxzJQpAX6fm+t8w5UAXaw4mU3USR8rdBR0YoofEB9YjwRT
XfVmuD4kJeK3TV+dXdXTsxBtNSA0nG9m/oAIqyE6zrKp1tnR8ouzsP4bf9p+LXEh
ZW+2xl3TUUpm7V0yvTSCgdar1MvoTw5CEdLbz2B5z4vBFVaTO/p4PlZZ/G5JCGNW
+mGIvNxmme6FFrw8OphgmKBHQp4FaF6OtEVYhLcl5FDa/8jx4L3Sb9+fzrLAEmeJ
EedoeGsJkWa4a5LjYaMOlUshl+MChF7aJTuhdYq3bhWPFDQmhbsQkpifdHzP/hWF
gRT2Tq2On/p7h82aU3lfoQ3ut3XdCaCE5d0iIeRhJlZ2dBXT91RyiZOlqnlJr1H/
5YEO2SGh3Lf8iA+m8cZUhzn0DPLiODbdielbrwJPwv5pj3Jh6BHj7raNSilEeP07
qupD1TAAzzSVHfmP1ronB99CVmhNEwitjuq+Wblj0p9LvgMKkqaeBCk6A6yuA19Z
Co9oHXVr5fOLI5mfT8HpbC+seDny31nnh6fVRm0KXnz7sJji7wurs7Ccx4UUfMPW
s5BfSI1cWoW3CXDkQBWrtauLY5g8xCv+HbqxAZ3AzbTYDlbwVVQj6qOJkGNgwjyW
FzvMocE1qoZ1KNWkW1nkYsDP/4GMQyJaql/G5GFjjbJd0WdFeCg5A9KXM1/Tg77C
XbRgdBALQACRMDPtE48JhmehOZKJNt9iC9JH8LFzVLO8+v193nCQtse+A0C0wsDf
ECaq7xFiJyH2ESUXdnsGgIYpSUooMyNOHkJIH+WOzZ4hQedqT4LJK8iu2ZWPzGlr
9qUeuZWTl9q8IoytYetdvdWLCOI94fbe9saVV6QEWuiE2nErHTPk1gwb4xaKNfem
LdLALEqVBUEXOLeu95EiqIg0xOrGVkGT2FuWLBJIkIqPUcW4TSOUMgVxHCLLfOXJ
oKq2KNHlIdlmjHURimpvYQe5KSjA1Wn+CNd+WGBSYzZepTiLsCNHJIuFuaEBKGqC
QdQYApNiO1E8t7nAT79M+uKYCyP2t8w9Tvm+t2j9sWws9bgtit3B0WbILvRnfw+S
HJr+9ybr2rpBB7kvzut6tzyH8jlrwYHDeUHWMiNNZCv9zkhd+221rx3M5ck3rX6a
p7cNnUePYkM8nqzCgPrxOq+ElYuA6EvJFAmBm6wlmEWc9iOFesAeAl2apBcqnAnR
Un2AFRuLY9ZnklxKtunpyS2wMTcWciwZwUb/4re6/+i3783kZl6Ed2SNDIY5WpZO
vZjkIHbybbYP8C0i1Bj5qyR0pmkPwZwtc4CFhkl1OPZZlBFAfMaFLVJqvz6IGFV/
UaKcM/58+CKYGMLnaJj66/lPAg6g3o9T9/h5lMsyPAej8lAAOE1o3GWCQ8q9PTWL
AliOJPwzZZT6LqYTF4Y+rMThv2JV7r0f18QUdt/77vYvPQ30M73dMnZ1RIejR+1r
5b+u9Kp47LSihkaA7oTztYy8xwk7T/XtXcUz/S+Sud8pFPLUs5QXhkyXRrBIVNcl
23hiDdnUCbU8TFre5MoNG1NWCja2xV/As7DdL3+X7MLHD+LiI4K5Ng4EFeMr7Ani
/k0mgLZVoUvm7TSeyxc7HHugINkeVe10oQ6yM3ZRDkDMteh6kDvp3PeRbpFSkb/q
zPEzx8ATtlYybbKwpBo+6pZIvbqgSFx/xmdCC9dC8ZSojUwqU668pfEqcVldoNJm
aDXNabvxVARqfXxFLqbSAsew5j6O4fi0uCB2dvCBczmdhL4c/onX2D1vZOAxbGqH
5jVPGxd6t2f2qwGybc6T6cud0y79lQjFx7xjhjP1qu7dyg+QRSPJpoF4Lph9x7Xx
Dkk6Y3ORb4VDLlx91/Mvenr8EEYqERoQA///v8v3dR1+Ff6xpVcJkSEdOcgEsgUG
5IdzsKLd3SJJnBCWFzb6imDotBofATraj/vquznW8oT7WE3rYwLqq8U93rlUE5o7
1qBs/ikA1/ryjZqWHxDOIIX3GkQOaFtpVLy31dbuggA5i2SEcKdZxm65a/yjyOGG
ix8wvCXE1G11fsZBTLTmJz0P/z63f2kutvKMS9joq7rtpCORl9QQuqbkxWso2D38
8H6w3vhXh+OfEP2jOHsV3evgF/8Tr+2MnJ19wZmFJFynqdfvUAvhAdHlDZYOZivJ
Xd8cIUp2ou3vO6NPlTXLXA2V4J4x0jRPTp4ROuWXfTyJPbTP9Ao8ZxYTzTNvyTqg
dlKKujqa5QKSCUjutKbDFgzYRtVAxJAa33yGf1Ivx+iTPAJvVrD3F3mS2ht1HYXJ
LUlrHA1Y6AhyRH4G/GjAYoXyrRidmPqqfr36BDsBmmjSJegOPI6fEMVQj1Uyur62
tpklk9+pIIWKu9ZYMpihRCW6BB4aftHuxrZcGxAcKK5BfBupCVah1vw3goWJnYB2
i5IDqcEr1zlPTYGN4VxZFeNXpFUmoGuYkiLvNWuXV3U6uaXRcEgp8lqDDD0F7ZP6
7+kAJB0aciOtBoMjdwCpGJJTANEOylorXeqnc5YE+V7TB70sDl/vR9hPlCQALaJR
eAS5Zovay2mYHs6LZdtJ721EN8cdrUvZ7aVR15QVB9/tCCNOJSDezNv5hGEH4QZP
1n1dL60R1Z/sPX8ARUaW+i2V2qTgqkyXrQYlfnoZKQcAFvppuH0sAZBFMpqV4eLT
jV+Au9G1R1XdRATLeE5MwcXYuUCHm5UMSXBJFmNyEs0iMHndrtPNvTDUcqHYCx9W
QlIO2lrEtdpEvv9+tHm0NlJq8k4oHNaK6QHT6QbPAFjp7EXTP4qGp8xzHKz9vjm9
Jx3C4laecV6V6o9K7d3J/JPq4vYhsvDs4cJfCzngGmbr1fIiFlZ3g5Y301udZfi9
Ac+J+yva75+N2qWWWPY5LyUqI8DFIVkzNECd4k8uvT0mtDMr1XuMD0Dx3dVZMxb0
wCpqlAqB7rYot5FMb5eJLuoxkVBrY7UMWCN0tHZ/JhEv7Ww6H46fu9L9v55YbF2x
EEOGL0lKgCzxN7AS7nxKJTpyxXvt/nLMXOjaIRfPPvrIGLtKZWI6TPf1rEFjbZCh
X1hESniVdi7jXCX5gvl//yVnlrSD01ngE3fHUJqNePV2NBINghwb0g5nY68YrxUA
qyzfUtO52zuvJ6nbzRxjrfQIzIIJ9OFwMApYtfzaXq9J5XqfsNfLnmmaCd6eYZaR
Kjk/JhBGduXfEOjcPoL41GW7AlhsubE8s/aOCbOFUKkqNQ2gcY8epzDY2uUKoAVY
R2FZMYLU/hJjGX5IEed+IM/8AgYj9ziIttupawffacF/gqB3VeASlLisUy+LIz/X
oZNomG2HAGIMkk/z/Pbi2iU9H0lfCfnmf9bB7TYmq1Z+zxVYJMWClYauF3cMkuBx
G2remu1Q8D6cfvnLdICe2VDeAD82M/Sbz4y8XV+4bVBo3MJP3AF5sTaY71IXkXSu
gOlfAXj14Cr/wZxm3+q/bFEl9Xxy/CT5FVlnYZXDFYzLJ//zOljMH1n+blsP0quq
k5ZpJcB4jD53xoHHlOpBNCBbJXCah11IPG8VCWbr+Yyk+HQvH5MvELe9OvElzUbT
xzvCHh7jJM8LVbhil6Hzz/zR2nNijDVDac6634ODGja9VQB4yZfS3Y9QOLViXSgl
HzJJ58lJaGZO4usItMrzC2ZnFouFm3JBnFt7Wcy3UOOayN4qLXKhpoAU3sQtxvRe
WYgZJeoqs5zKVhsTZxCCOn4d2OjiAhQJixEuq0phMZ0BNudINDmPncBLGqs3lXXa
QKi0v79+n4s+3tIemrEuPgJlPkal5pYCyoFXv2aosPtGxpJWvGhx/1BQnYUiSuNN
N4WYjqHgpjOz5MFmRTr4+LaJGs1wcOZkJ8j00bRrivu3igNfi76AuY+JA4LQVsx0
6MBLbDAiAyybAKsoTCP9/RAMV8ZeDacukYS1VnlK6jrmC+UKURE4cR47/If3MFxz
kKmVTGM5maTPhXnrZcjHUE7WAO3JoGa8eNdLc/TrjNRZNa7kTDKqt5kMi1Ndwh/l
o07jF+cGtmrzT0iifHVsrgN45sN1jP6geT6d+y3xLIFarBsUkLGpZ+8TDlGaOvBA
myFJpGlZuVVn7Kmu/7GFZDC1LW3dsnK7Gwrk0mYEcYTh5c8wgXq32IuhVqduVOiw
2KBTdnY4MdRgdbTGUaQUtF4ZhfnKOHTQ+0AdYaBWK+X0YB1cVJ5p39w1vX74qiUf
76X5JB4W8ad0YqgxZ4k4R0Fe02sLmIWL9g5fFG36rBaLnfzcWyrjfbqvDN4U+fl5
+ChGz26ITPfrWsPacM+9iVdE8Xx9W3mOW6wvXpYFh2juAjdsAKMZLZFR/komXgLk
i8SMpLSPwl0A93Ikq/hg/HGg6XnxK8JUK6mhM6DuXuciMBuydodSKNgBjsQGLUGs
qiOFp0MmcKNKTuoZ4Pzqt8kZE/Ln6Gpt9ZMgqUNhe5zx44EeAzMIbpvcZcnqu/eg
5pKKjiKmsIc0lC11o13TNAevcHJPKos16LiSP5D+NOc/3vOEsai6ZmIA6TpZKye5
jen9nbqLC47pYC3HFbavEcLJAR8onn7pvavClOhNUplgmCs710RcSkjCVmfjngX8
xoiHHKsOKBC9LR8GMNdbw9lekzbwOnKsahYjZS4O6Fwt3cTEHYh1Luz1i0H2UMWY
uCCca97GmANYMnjpL6Sn2svkyjloGoNEyDb9VCUXCOazP/DAaXZaPUyJWF0zCSgL
acOCirxAUbtH1079jCOKUW4DfAM6codWba3zCbixwulFt70ShmU8DNgMTv3LTI8n
vjRcgW7yhOVcFHaZ3aK7rWaq+p7hvkuxY9MIom41T7lj/NDTRM7PU9Id+w7qN77c
M9KiXl52zmUQ70wTzQXeqqFdBpg9UwnEhcs74FA3kIqYZIA4DSxhV74GLI21ccFR
UMndCHTTa8A9HdY+eA1w5enEIzP4dcXBhvm08i658dAy3iRJI7mrE4i21lz3A1Fr
7lYB2XWA2q50OQ+y9g5hszmh7Cw8L9lZBaCUdU+E3yd2ODX9MZExeCVITZSR5FxA
CtV5ue+cX6B4Lw47rt4T64e8wGVzIKReQlrVvM/yGVfE79DvIslCCy1rkP3yelmq
KqyFbhxxowQ1awEZ/IoI/XRm79VX7JUfs7gUlu+aNFZ4KAQXOOZbKWfBa+wtnqfT
5gvZXwc+1UIpFVn6cg9/guLLPE5bVJEe00xKketZbK9xamHy7EIHOmmgs5ea050q
OZt6cDFSNrbaHIv0KGQ9dS6W+/1JCvOmuwE8g0tEBq9v+vCSnM6XcC4avaWLj5cL
e9CJ3UlUbxDtH4iOvFTlHiAMUwDsqd2NEji8uRPp8uv73i2zhm+a3kLgt+8PGg2r
Z5m61ole5JLGx8AcZXtJ9+P5xujCK8/HDH3dovBN1V33ZyV0DWpxCPbUa6Y7rMOW
achpBjUsFtZMMXTrIDkWiJHT4meTqKWUEx5yRMxfd22qFj6QAE8Tw74ivEj9lqA7
yAQHA3/pVtnZAfXyYPZk2bNAGpHTHFh3hdlEqRrII3LcABB/yjoU4+yHIRSXRKFi
delMBSunOD0O4ITFt2lNtNMVVgwlHAj0Z3aSZjAezjOxNKqm5PbX2+4byGpcVARG
tgqGyzUleugFctN77LXDnEFQlqlJCJTvKIMzDeI5bwMKvGcsStwNGGXy1c94GsLF
NtY0Wgl76hCgOR8NB0/0HF+Ayuv6ZlDLkZFLSWjIF5MpNpdRq+8L9v6QAz5Xc8r7
A0FnqpT0dV4PeWnYpU9bnuJJlEY7piIfSz/PM9cebH2/q0Ojkh26KEpHWxzaxdYM
a5wMie4ZsmSTkrNuRUk7jtBuxqeJGKSxhOtRm94m9EIwmpuSVCMT4zUHLWA6kE3G
dXx3oL7F425vzvwgA2+pOXXwgffeZZXQ0bk5gT+PRpLRbJviPct1ARMu25jyUIxi
Dwa1KwkwuWbYtbjxiyNsB1QIyrnrvPjJqkte3Ia/PpCV5otDDEhsDEIY3HDDuHHo
1MarluM3Hx4vM0Dym1eYSVwH+ttEVWYrftI6DuEavbwapYEKM7h2oK16uo6jmhtx
WTTluBt2BKLVl+58t5tUB+zbtZfu+T9T477gg698Tf7jqE4BOpEoCzPf7p3sPuLM
9eQrWH1Z6XHFnsM0GxEnd8vj4YM/KMfC8w6vrQBy8qO7o/OI6FJ+zX7BrzENPAF4
GTOmfMC8KMiDf/61aAOPdpo2qAgHxnF4h/84NXK305FOGgbXKWkIXkuCT1VvpK4Q
9E/YckyERtEJtbi9QH8UMBkVzrmOqOMg9K1sm40cNES94lUN/L8rQiF1UheLd5zE
ve6hjvmfL7R5lCxL95bhLUkMOx8n33RZEb4OelpZ6EhVPaisTi+FvTD1jS0WJCvl
suUJp56xqy8vM190QwlaeaIFG1TJRaV+cLYf7Uf4lGnRuquo4HNNyW1Wre1oQ/7E
wiPmICcEAPcj6RDO8pHj9j34hm48OPRnyoaMRrA9BewzkG4S+B833p8uB8NUAStD
7P2sPFDjKAty/ww75LBMjlz8CD2/bZGAri3Xs3J/r1SkZzJ94ls0abWea6PMPeGV
yFyqZaaZz5zmWpHoQG1DHHi5JDr4bzq4QdoMohpomMGcbdTpn2u1w/BRrzughJOE
/KgfaiF4D/+AB9V6VUzyickR1CMmw8U78UYNHJ2lqu76tmWpqw40FYg8oQkUHB0d
w31DAaHkEL/Wp3KP1NpURZPYnivVHG41TZ2FtLABIaqQMmJ1NBKIwYRJ8EMb+JKU
9tFju32RyGmlaQ4Fe0FqJiVZebt9M5verFmsML45Bf3OsjGVAoYfc+fQJlnY9PyS
PMYXxyhumPYhpJ0ZULBQG67Cg0ETK0X7wXxogzoubjhfOqdrwiqe+sMwopV+mTLV
t1yTkS3PnEzzP/R4gVQXovJPHWosutorgdauWP2Fc/VofsiG5LjhWRoE3WPciDjC
Mj3z4BLpQzoICg9++IK7wz5Gh+W8eXDh7hrH4Zrfq69m0EY8EDjYbkvtA3jD4bub
SCjZCYXng7E6bF5Dl41oHQrwFTtSx0ASgHMy/j6/7evtCx9tUpEOAsJm51Ia0yEC
Vf9Yf4/3T72rur9XnTXRgcp3lDRP90kW/vrqtepQramk6oqExgRJu368/cltA4b7
unLTtak+feg83Ij8n12lTahj9d+VJasZve6EF5KaT5uql3HeDOKzEOnQZ76+gzag
/FNl3TM10+gpa2UafuFzPIFJgNILU90lWxODDr8umce9fEkQ1SXzvlfHpT2wGghU
wcxGfphkBCZ4SlZzvAab4f2Epw/tQVkH6Clh3xIr7zcliW7r2Ai3OVMjkxBJjL/1
LPzjyuvIQEOXI22BbuvX0/K/rc8rEkSZ9ODA+0NePxGb3HR13qXI9YsyymJHGEjv
zKFL71C4Olf86rONDHdy9FngJMQBvj3PT+ZqlVmTCLbHgSn2cxQ2qufDoCfPw268
UMjLDbnayxK8ua7hG2+d2vBpbnPTAENTP5wnMAl/w/xYiKzt3Z+l3i039fiRE2h7
kYIC4fHiacPsk9fFtNXvq7LxGUFmkA1hFNy36oh5tKocGX5V5iDQNEK1YS1ZBfgK
6WnyVFNl0ghwZX/OsAxOrVqQWdvAgwV83iLZRjUotMM1Np+ZZc4FgZPUVy1/EjkR
Qb0Y5+RL1Z59oJU6M5jg3B1rV7tbtFHqBB+EVJduf3ZCUEe0rq6oYc81xVCQ9bXS
MFr0wnuJIubSJo4LUfcFIpJzCAiO7ZSSFgjHtthM36jGUNTvqL0uUhT9B7bPtHEO
qfnNOkKZViof8MySAldI2Qj/JmT4GsH02ZlwuescZMvLMeReGpg87DXH5Dsi/r3b
TMhkqcuZUXcRg9l1uJztGzRcNrE9TYzueP5duitr00lx03f9Jt14/fay89j+mqyG
OT9ClVBU8UopCjKJD7w+ZDWidWBXN0oi3OmbDeQcuj/Ca30qbKQpeZLX69S4vDni
jlK3/po/25wnqW98pNEOq5UL1hFz4shaeCYwVTonIkYXNRWW4dysRmIULBt4VFVd
Wpfyl1jF6/8ueRJHup2bYW7+L4P2kEoMAhBAP8XCiDIXo9zwLchFw45/ihxJdVyl
s+HdCFz7ocHC3aw2EGLT1GupW9Xq+UFH9hVMxu5PpBmsDbbtXE1AE1P4/MBCR2xj
fGaT2hF35NYNrILVZU6h8QqjlUBr39CLtsBDangqNotGQyWoOKfAdlISJKvKsph1
fd4MpTRo2nNPP7i8gf+ku3YM9ZvlqlpTlYVxIGIcJJIVXnhNEmGRr5nv89y6e73Q
kKvSo2UqtYCYK5/VcAIwYT9FPZoP6PCu8Oatqf0SSzZJeeZZRmzdFhIm7KxYcMbY
TgYeozcaGQ4JcYJQkmAB6LOml39Uwwe0IYvBi/uuxvDzoU1RRJRL/6LtiI25EPaS
dmQleRFn6B9tDNtYjUxOdH9MLEIylJCatYQVbO+Bj/Siz0xf4EXwXewENZyWKMKd
zlmOBt//Tw1yxl26H3Hof0dYwQrKYJyS0YVjcgWMU7IGwt4VHKiw/hcs7f2Y50Bz
sqFpQd+tZA2evEvYlaLH3a7qDimU7C8DTxMcQqEnSmn8Lg9eP3w21FNVy/iQh2UT
jiuOdBADvy/+RsNNzxtfrnJgPv+N7ilVmw5JpQfnWq6DhN1nuE/lhTLJPV7hy7Gu
PdNxFg8YTR7rKYA61dn9Ru6G45L8nRuXzOQe1+qMYTki3UxbIfVlLZ5kk9hEJgKQ
1WMTjfJODkWK1jCpawCruonxI13cj4xesgSGUsBfTwg/NR7ZmLiz1YqzNQ9TgAbA
vdgXXGtZh8+EirKMTOCtb1Rn7ejKNsYZBfEG39LJ4wGZeSuHjmvi+1bJ3OTh2AuX
1Tc2YmQthCGBUCkuSkX+irzFRTnTStZmIipJbG5G5oVUE/lcGcW1USnnjn2dj9dX
NprhuTidWyvlzwa+0DL5IXEmuTSAvTA58xdbhfqwCToF0YxJEJKC7078Zh5QPE1h
fyvUtbSWpyemxbLRM0SDvKiRVYnucYV02fh4sin8itjLaWuK4LtrokFDbARU/wYk
MAsb7kavn/x8OAgXtC18pQVZZTiyMjveMcqAORTHMLaGg7xZZHbp4UQMPV6B4qt8
YoRkCAZURW6/SqZhmsWxPsdAx/HbbfiTJFEymP25srWhWFTtdKcvzhtA1yvqS/O7
Rb3nK8OtIOTn7NPnchxVB9deNynSHVMdmz7RKitqN+R4rZWOHP9s0AJvft4TCSIh
eLg7/feS07DA0NaBNsyKjz0r2LSTJAFzcwjvjv15bstPrfWbwwKHPkx8t5S2f2Ua
2Dgf105MBf89AYG2HoRamvyPCjhvra20+J3APlOFhhc1Q5e3Hzc7dzWFEtQZ+rfE
V8l5glK1jaRemBn4DQQWtubDHAP487oi8u3i/Afz6cT+SxxJWLc9I6kSsTGwxFdq
PkoJfffiYI3x0qKkYwC03lFM7E4pl5HOhRdhnCkN8pg6BhfGG/76CHCeGJKsjKQb
5YPOREugD+N3XsTxm/FirDSJGHKyn0U6PpmX7YhextDHnxXY/FXHxquj2r2boS7Y
NfXgwqUYWmYMMq00o4LKw0xkNvvvVPA2C550yZQiohK7AMKj5nS/4YIPBhGXNErO
0HR51CrfVmjrrzkaMDwzcz6qxQff6EcoRSgXIuM4LYLTQPERV6dNesZfDys/KRRD
f8RViYxac2kh1ENtehoyiG2IbAgH/doA4k9bids466UXa48bwd81h/FNTvW80WUA
KRESunWXTYdIvSw+aWBItGx/6YJbzxt4s7S81aqfSEptjTFHtzeHhKs3a8QLQ4t6
hiV1HoD9nrT4HLSmbGM+cBIv6ru9ghOY9+aGNdQdJZj/ZUC0s4pH2z65ABvuxkcq
N0FCmlcfgUeR+NkWPbdZ4l6nvA30ekLaz5U1unhkmFrcqImqHUtgoKWhFb6T/71q
K2THMWjQSrao+UW+lgSYovfm8BHJrRtQBPjZAjSoR2ffhU2N59QUNRjQHIdLf1MJ
NMcnliJibeX8+O877Pg3p+7z0qv9manH5SoAcO6Mi/sIrw0fXMWZTpgXRnZWgNJd
eDf+WTQCIMjSNcvWG7aU7QkOl4aKyaQUjPuZLghQ++FHansmOGmXY8u8voprCTEA
KhASDNF3vykJRw5Hl3wCSjG/r4KSgzc/Th683ijT74LnRr4mvn2GMbSM8SOOQb2/
9NYl6YczJueOZBkLh4Y6vqMH70kGXXUFOTjK/Fkq/HH3Bsb/vwDG34GhtOzjK8Ma
wqOgTnkr5Kku3ZEYzpDREH3+D7HDq1VzUA8nL7x4DgfdxLGABevx3QdvGMBLJBma
BvIuhWjKlPTKZ6RrHFtNX7W4DdgJUg42aDks2aRt+4TaUmGEMeGRrP8TysVY1WWX
3/FWgwmtPeqc47GP5ddk0ifamSqfuMY4ilLxw8lKmqlQYQWQtlRlq9EbaLWCejtC
TB+KWp4IUuEx2dJ6AVECK6UD3ltwkhYYo8fAVs3BrbfFGhXz8QldgU9jNpS0mCZU
uWLMsJPkvE6rPPngSoDerAFpCy5uM/LwqCAKh1ktVcGpWgSzTGtEfz1C1i5u0lTU
tCaNHv++V3Q5/G8wTyqZN7luiaIH4pAVQbVdsqLGdoPhZ734ZmiPyLjTm0xRtStl
Thg8xlOfzoKV1nOaGnCGywMu70elYQTvuwHT1zGq1l09K7G1X0aw6hxfQsPl0Pif
L4TDuplyxeBVTBO+tGSR+pIkIaIo5wYDj08dSieajZv0sK8W2mbqPbCBooUrIYrY
+QZcwPQkBcyp8hvV4cRXAFM1YDG20UlUCP77Ku4d7EeoZ2+E27O87aJw+T5clZuu
ryr3H/wjuI2Cvjv4JxjQNNCIXydDxAd7+cIyguavFfd5ZqLb7c8Gf8a+qEJHKz7Q
gnsGFjrepLNLnh90DGXJn4/5v5lsDUyJvi+S/BKmcVp620fUm4lewY/StxmZ/v9x
j/cgKK9D8vWjkSGTQme0K18D/EevK2gF+juIbqq33QoZThoul2aQCglPFdWEuLic
bKeRktnAaJsj09PLlBnqbJoaENWTIlKFSGogDkv/QB/Ow25FQoz5m8sdhuFfJEst
m9LKyMPWossdvomjrd1po0XNiANVuuCwkFnonC/tCCFiYL6qZXntDtjcYWpyA+4N
D1fIrfWH0ZVquphkX1HoP+Hn0OPkhwcj2CIAdlBtq2076CY0E6EQBTspTbJLlPv3
pRj/aL13Ex0Nj5d16nabkaC59meGfJSAMb6z9VtqTOoHQ/lBZTUgVHL2zWNvOL9Y
98XgWWm/2uM36nzjmpuMs9+FHbxe+Gyp4YF9bi9tnj9YVVr7/QMjHBVr2vcg7TfP
6MDHZ8GNEYjdwcQg9Vf6k5jkAUQplvFWe1QBS86XnAPclTyns40LYd5XukHWf6Ny
vgKhihRmh6AM9EhkfTFloJEb+Sj1+OkEc0yMT454HAUzuLvId0v6v/IRgrbyx+vw
ZPo1tcmksrs4Da3IaHNWsym+HwYdhX/c4apNYGM6J02TedGPdVAE/PLA4S1i9h1G
jKdmuhHII/530U7j15/iigovjpt0skcULQVcZv47qGkqFUIC0wMQCoV58X10pfJk
PTdF8+pPmerKp44Dc7ZOibKMgoY0YFZ5/YpI8VUt1j+lcvJGhccMIxUqPN2cuucD
Czbo50HzzunA7SUj3r7N7m4uxw7SkJucBgaX2JUeKsoxZoK8xJpRnnRHZjVsaWEb
wP+Osyx2PIsK65gLUrGM7SLi+Iwuu2uCzuzBa0eytGFAxgZBTPeCrUSylbwqhIdE
wk1zNtPT80OREo/mpteolSzQTWAAI9niQqG/p3FHsspM+MedXlrJojlp1y4mWTmh
Qs2BqCaixgHOW5F1aRdbNsU+DjF6Y/Jj+BcUUj0LtZsHtpoUK5BzK/IJx4ZQ8CjQ
Oyn2zc0YlwYw/4SLgkKTS/d3yRRyWLIpHJFL654BH88nhAikmNrLrbjGW1poALIF
yq+515L/Pwr+z6nrX9mWqxsLIk/rSnGv/P5NRbjhrmpYUPQQ9kHr9MiNmoPCIFLy
l9PpkO5kEbNijmlY+zP/YtdO7TvZd7/CAs4iSJRg1dFcVQbv5AbJnTG5p1FMzCig
HNSfzdWriEolPLWGGete+XxWILj5kQwBz3K0Xd8zvinp8czyEJv71UoOBHHN7CmH
8fwPMv2CRILFDVEeZtfFwqr8GhuW08nsAmeIvet+iDbbQvOmxyAn7ixDpYskbjFu
fTKvJtIVOCIaiCpjNaHFPPORO88f9lPwMB5g0YfuvJGqSXpTED1ap46P4mBh9hB+
1PXjPq3hCqq15/keV/W6+yMM4mY1LNvcc8LfmaUmRne3GUlrIsHgfXSxcz2Zjqn1
kKe4v7DUMoE5o6JcjZJUsazqMAXWre94aUE1Y4O3G79StS56V+1kOld601yT1I5h
njirz1dUnH+vW7PUIQGIyOk1+RLpKrEGsnMo7Laci8Bj1+xOmlY/mz03RzMZVXuu
QgpwixziYk3f82hcmD2D45YZYwE8Y8yojSuosrNfn3gmu2BQW6kWKAj3ZZo0kcjq
zN3FUxIPeuiHeUtU7rJIbLkg9RoZ0NrNKuLZURlma7LG6yWqEOw5MhIs5vLvMySI
oMye2n/OITD4+2XJM0nrpAOwQtpEixrm8pjGWvYOzSGvWCWCwY3O/Rmas9S93vLI
inZUH6mlJ2O6mR/cyjuLWuRR2e3vaITmaTiuxCHCSZ7Dg7xo7XtZzcBfHmMHehOY
JFFLpZBXb2tS4B8vHjslgGwgUgvv6e3CLXn19f5TtnFryJjjuJSzMm+pEbMB46/N
zwlclg8Zo7tqqixGX+A6RejM5Z2ceuy3Wc9FbYA4tV/wK4k30VAClwcS/NDBF9sZ
AyTTLblLYMMveH6FkTZ24t8zZiCSn2aYO785L+LCCEYEBP+ZqtsFR+mXN5sFh9Pq
RPBxS2SpHVejRgXvMWK/JRJz+h1IkPTNbxdpXi5Sf7yI7Te9FoEQ0Xd8YuQmdnWf
pb3WCBI3VEAXYXPjNvh4YbWOm5DFgYETXOfCw2dAcyRtEXg1lbGWBjixL2x4lMAL
D+uYaERS3i9EAswVxJ7gGk6xQvf26z5dc4KHHzDckYwVNAbiG0e446kUqXAoB9TZ
muZAsoNx3tmzuEmDxrOrnoxsMyJavxvGYTP9BMdB8eFTCfYX7rGikKPOUXTDCrQi
OZP9KhvxI9ZiHqKOJGSDgpQ0xXNDrCputbLY7AGxZvhXMY8f+aVMpHnnoOP5Uf3D
1Thz+nwPvjMTEmwICDOCG4Rr+YmVt9WSU8UPGdiJrS0kbtJGg/gckfhg0TBFwQ8B
KV6iakRh6jGzlKqAjslefHozl91GHOtUj0n/+HZoRU+N4c9XaFHTOu5tH3FSVLXa
jDd1LE8wee7cCFpt+NQJ8sZY6Y895HTLNLquxmFhugPrtioIjbzrBUtfkCITQDoN
RlvdYYOAxDPVWe/xwHPalYckPATUpDzixjLJiCFT9LBeerIDQK2AV+Q3RHTMjhnt
sYxPFjUCkk2UHiFxxV9a82CmQJuu16Jm33jVKGX28HX1tcWVHDhYkuRkpnOrrOUx
j2PcT4jinTgpWRgUaKwnLn1f53R8GgB4BKepjoJnC4vAzdSt6O88mDFYNKx0lAoV
8XP/7xC4wd+sKigY7AT0eUzRCTQ4/bLzHwnIzxhh8YZVhmg7nNWKphSIscritF87
+JMxx1qLaxnA57Le6l1wRYqqvBvXaGZupwvNMc+eVMCGztoCahHLTS9BbZjv52J2
qi2EaaFyO2JjAVDRIJrpB3jlirDkUQ97tV2La0LuAMgsYirAMKEYj5SupBMXUtKX
G4UmXmvDSp6hMdcP1IQ1MIxgiWbv8FEGwI2qoLx4/2ClD8tVT1nfhQPK4mPBCPxi
/7qXUJ7CTBdX6fhpFhdJGSDPKhYsXjFsev5cAGUlnAZWdhQq5dUrQr3m87OLetgs
73iQMLqsR/ecwTR+hevmXCyFflkSFNVO6jOBRkalkCVR2IwKrPGwQnqa7ns0P/gG
STLmUlAYekzUlVP3G8IKZ8lRtmWz4LlPSWrwTVxxHujQUaublGW168yIux4RxpNW
tHN9KtEnnjBBbysHRDMiGIxLd5LAPQdhONm5d+AXvBt0DQgituEyq4DWGScSWEIH
G/2Im7rID7Tm/HyVb8Zv0fMPLLB43Ngs9tyLfa5Okf1gEp8e5nyFRZpJ6W/9wUY2
VbkL9zBPd7n7u6B2x7fIK+SURI14/RcA/AVEgFbeeNqrSuFDu6AiETMH+co8GYBQ
7jgV1YQGXlCkOV+fwR+oqdKymk2USneeK2nT2WlR5HbN2BGNLqgfzpUwsblxYl29
bQSgnKQi9mPTp2kEPhxAlPLIpm2njGcUJLeyqNT7/m9e6To9NYZ9eDq7XE/MvdLv
cvwVtQz9V2HQjxf0AmcOASxsr/dpyG94AGh6ohwKT/0zrSkXvnhirBwhVz0ncFbs
cfzQ6EgmLlTeZ6LWZB7Cj7dsYnom6Cgyi/0opFhb8Mz1v2G1hO6kQEPUkMZBNv1S
WTrJvyK3hglFzgnXgENGNDm/fmMKcmc1USMiCRr7CoetL0t/ONhD4ybshYtzYI4T
tiGIQHxKDh7iHRZryeDxli0qk5doTFlW2K21hJXikkWHK/sHlScjNbcClbC5IKH9
rh7fPacUsoPcQ5O1ZxAPlKKrU5jezfH0OK9b2BVTUWlrm0nSgWisJ+wYyKeWdPew
VpMUSxt436aM4cYqUWWgOV6XFvd8BLMjD5Bi3KevI6jd806CCg0wcIgOev0LN3+T
rj2SRgs3MLygoLFmitAl4apwmJ2tYQvbQs8ClHYk44XPtMHm1vT0cp0bfbTMsRPH
pWx8ylLh2HX2SVgqi7NpgiTpt+Hq/sR09ZoYWd5454ctxwqqDyp9BJATde20BsGE
iQtzAHg0a3IRML3qfYMxo17zpIUYV8nv/nn4+qXWpUva5L/7AOE6ouWx3bobdkTp
fTV0QnvNrKG1heV1g3Uhj7T+9EzfSUOw8FjUlJ2z6ddJr6xJ12RH6UPslsImCBaI
kcy5aU/7NYnRSCsxKpaU0y7By4XsKJUEEZ3PjboZuaEwjZkDlS6t2n19n6Z11Xhu
AXLI0a93n0btQEoaUJc1dwBYKiGtJooSjXH5LYJAW6Kw4ZCx1TK7LD9h5wq3k+GT
27i3JBIK6l/ZmDTmNnY4qYLp/Zhl4YYXEINz5wvOF1eetwxuNz6weqDQ3amjSkwb
4Xv0oukH060011bPa6wpmU8wLRWxE0mClh5JRVdY1DR5Zvl0Vva4btSdZTCVu/Us
0EiKDW0AQL47btLgXg2lTcDHDBSd8dRrXyMl41zG0zSdAZ7gfWcuGoIyqT4OYN6Q
Z26AdVdzn4FlvrltAqoo+GKBkIgHmUev4GmAU+cqn4MHznTTBSq/hmJep3uw53gY
Br0YA57jxXZFTLB7nPBYcCtTAHiwcI6JFZdwifhlL1oGLQpkMAz9Qn/zw57o6NRT
zTYlfwAOsaOkMHre4AW7kXDrQMEM+q5ahcNFoVgdoOfYvOgcIE5Nfl0fekpDGUvH
NuYy36/+XIKvi4ozywu0rt1JblsjH6kE9HK7XUduZvMe6jNR4u/yI9hXjOXzG0tS
+fgdXQpnf2TwvZ1/iUmOvD7q7McJsr1+VApISvnNH4w3itdNXyG6kn9juqazoiXj
6craQ9x6idY3c5t/3t79REHp535KrON8gSCadKn6vMtSI2kV2sMJZ0pw3pxUYCeX
nwHO2Keq/RSXbf1q3N4E3pnTMcjXuZnMyK4We+t4X9bphT00n24FGQteh2zyPBh5
7BbcW54qjYab/fcRJj/yPBw4HzjsP+BpbsBMLDb49XoXkUgzm6Gagx+x/eBXS+3d
G10OZyqyM0zOTGPR5kO6RqFV5XCr1GpQqhrhDtkDqf+BQDuYpwcJKKcMYAlCfDnL
ze7YobsOw0hDVcmrginkD+pEtI3tCz5ASJwUWxwztlPuVPS9ONiRvQWZYxYRYecb
pOT1W+rzJ09zB/fWhtsrHeVwC3CZDiwX0LWNVLinJ0IM5HBpUG7DYbTewSTltQFs
DqinT2uH9LuW8eDXUhAtjnA+kLREK3/LHj/iyMghrzvxVOKxFKK3nM7/pllR6OYC
nyl8jQy4rvBf9BS/5dDYYCwkhPGBlmFhzMQVWhweIvxB1c7RObwYd1lDNfkzfGIs
KJhpUSSceU/EMfg0OQe5ThRICtxOjxnhbrbBsITnqDLvNLnP8tkE2EyrNHpIV95X
5SgbaU0Nsfx0yy8TndFVGX+abbpnMSmol1U9HMsRN1S/8a6PMK8VnHUkNsW8YA0I
WgT42Yts3z7J7J55jKVmjx1qrLRVDpXCcRxCGhgAXGTF8g6vuCPbS4jpNKG+0560
QZPOnMTdb6IL5WAoe610gjG5NbwupRv+PkI0cSKfPJnsB0vBXc9L6zclcjvsuNcd
tvQw7Yb6agqoAYn7L6lvgFYK03Qm4fAokvzQZPtbgNQSFE1dZuJjs5nOurS+Ogbk
O5v3/z2vELZvLBXa0qFmN/yZC6gFnVcE6SbIqNLsDtCWaHZww/b3XkWm7eedH3fA
rm/sYkYT7bnkN0zZ44Q7JT+4e9JBITexn/eh/y+NeP1BMJ9NFS0is4ftKRjVYqkw
QYIUnvQ6Z6EWcy4Lt0IOKeFiO8pmCP+rGORmd7cfY9qMmjgj3K0qDM7aSU2tB+3z
PaugWq5abeQc2/mQtUbnHSNcCxJLzv4oPoGz09xnELHSberveD/3sBYjZI4irPxV
tr6JOlIC0wMhYuKPOtBFld16jceTl5XBMA/YRHcvh/y/9R9+Mx8Kwy20vvBqE4MD
KUd1v9saPTfEkHkBKvp0OcJhnge3apBJQFHXES9G3BX97fSUpmuaCW5oClpqvwDz
+FortFvofC5c44TNAo6d0MuJxEGea0a0tEl2a6jvaGFieCOqvqVHjN9KhDVyCDkp
VnNbVPyKHGv3OJJSvjRc1hiNjlLUETswQ6/bZv1U3jzfxD0qSQeFGY/Unv45eLdv
2+yhlZOc+mO73dQP/n5zC+exkwvXLyFRtS86JUAqbKNappoy/ic74AQJ+pe1BFmS
Qlkw7pVOVte9798NTbVVI2L5ADrOKwgyObBRVd0ZJ847f36/4ZjrnffGL89UcNdy
51PyYaQWk7ZDJ8H+E305MTVNdS9xpUqHbkSbaEZMyEy8E25iDOdywfVfqhGQsIk6
ZncAJ40/E4Fke8w7ViW+z4SMq98j6ugpwqyLcAkeKOTE+daThJwHpJiITbFpiFHG
6S53GZAH3OuhNioPM8HcdCiVmm9tgQw8bos24eaQi55/lqm/wiFp+f6IFj6FEToR
8ZGbDJjtKcUSJXEo9sxo0UdDmkYwZizFdt4HgClWCBtjaY/Fsw+PMbBQdGi2tDVa
V5HlFohPk/LyhjkQiJTYTMVFxP6tjZldiKqa4MyliOjgY7GGbdRVVmZw9ty/RMHo
koJpTYwPmbZOZnJ37epx4QA/agHyhOl9MNSWxiyst/ufMAPLk76QGZhLehRr7gOg
B0J3I/agySCBrB5K+gWE3xTy15N3xi5pBQYOXYIWfRHjZQgiQazeugcLAxl4AfHt
ibWYAbR9NeP66QV+YONO4WX2xYCFMwT+lGTONWtVV/K3CkObDrr3H3kUL/5T6Las
tJCXEJgDUIhJz5sRQpkGX+RM2kCjtiwauADoLOod35GfS0yuUYzVLkmyl4XGD8or
eZRzxSuFGQud8KRb2Dn8IICREuZe2jbxlzRxMgvb9dLVM7FqAJStLPkscNBNpK0A
JXsH9s7haeOK0DgC2ADwje9vHJEBucHveo0xbJ37H+5bKH8HpBVi5lpNgtnkRsZm
sVGuNLdZkQBS8fADEQqokElWjhqzYn4YnApb1f2dJderNIPjatAuq2Liva+CbN9Y
4/cbc8kYnX/GBo8Q7pnFKTR9Xorin+cQGLlfCwvC+1Ly5qgCndWtNdbDdtKhlg2c
D8hCAvfcPuPWfGQiB5wnKyCjruvoUviudo0Tt7uIni8zsJJWo9Ym8ytPrvgeMurD
IwQ6zLbW81VNeFUtjkcYD90ydzqv/f+Ez1VmB6Z9DPEQvkoWg7M63ISzHY++HptM
ZTs110miS7aMHB+uGKjE09fzuI5RPOb+tSlMf+OSMr5dvxERPUeeIzoDOz5pSVt9
pYPjUJWsXLTA+ugkWMt0x6rMX8d8nSlw168pZaaLwq39NiJmIrzyGoPcrWSAgAEi
MWyzHOii0+6L3oHpZWKjDF0Hm6n/jS1Xrh9ggq2LeLi+oqg/ik+uFJQtjVMdelUi
0+Fb+tq8LC/n1i8rh1nyXymqXQakmka07N3B4v9GGODuHg58fq4u9cvnogCii0Hq
PJXC04nRtLR2EBtw7dM/97TphS8Srj3JRMsMgC8jwf/XGsfEcJT7ERV5bjz2pc9L
c8vv4AIlbslGMbeP/XwHxxOb4CLyLBlz1NwWQTAwwPTHJN382fRbf7UYuEk15pC+
7mE8As1MfBHeYEWM4WNwSsx2TsHP45KJaV+sJ57ySyLspWhjRVLswt1dEuG4eNNH
VKUhDUlIdYlF86fCl1AvskYaNpIyX3BxpP6wmQeUqWI2tExUZp2mXgTNWASm610n
gPso0VRNtzaQjyxsRcKhvAtQSK1GrurXg6BViPkRRhuu56c4sWXP5XO15B/QaoxM
ISM99WFhzdPGMaZRqaxKzpJdnkCSSMkaJL6aDbpW1QIICBBl+4eV1y19NL0bdoLx
AzoCnhwoDBjzRJlp1BEewQH5z6fZYhJeKAwrWotacCBQanos9V0hveSrRxEj6nLz
DmUF90wVNpRny9B6yVkHpRfXPI/RRY0jL462TxZulLHRWQF/4L2haiLqHSmLGvkZ
p8IE4vNx6H2KvezWdTnxbdm6Xy04YYRTwf1cl/a7kOrORBanwReNHpl8wKzkaOZN
kV6062ZD+l5vBTR9f9zktCYfZDeGOBvZEk50Rwe0b/qHG/YduRACj7tKl0+JTnf0
on/s+ZzOVOYq5vWdKXwdnvVpSHddnQlH0GWVCZEUmS+3KjO8158OTLa08tlVBYXg
5ad02h6C5zn0cOfBqXG4Jx2RbjpU9KCC9u5axPnh9ct1HYYRU3LmTuI1/DHfr/JW
Tvxlmg85Bq+I71WWjOkflk8+MR7lTuRGpOPNA6jvdmLhL5av6PGje0QLUqZk9FWD
fpOC6Nyz9ML+13fniF6XBJtfLRnLQ1NEetslPBR4949QIV7RAp1U1JrAiM4RV+FS
Vv3ljjzs4L+NcLgD4lYPu93Ml1SVH/tMQNg3jzrEoeIqcSV81dwRw0VfCoA8y3zM
H1eOIDsk+QVvRGmwIKj/dhOItPwCHkBv5vmd85ZSzTKBoF/FKKgl7JU2EPrmRCZ3
KxaMeA3dIpm5rBQcA4GoxFU2LsnEUB8fb3MacUfmu6SSdDTJs9+ISl8DpKS6O5x/
Wl6ekix08YzYIE18q5qRa03lTIc6skpU1Il1oWeTwg87QHa1TYY5J1AsRnnQRheF
vwOGw1khb/eALnK30Zp0ixy6svI0/TgwIbnRmgNz4otCT2A3DR6tGPF9Nhyg7R+q
2HbDsSkPUSPsINqaRQ+DPikroWiAXxqjB3bmPqo/yuweWlGrHnToBTKLfbdsrGeU
Wx5mi3UR6wJncPCKs0/jVcNcY/0VjwX0RYrob+yhFykcxYjDiC+BKu/IKuhcwu6u
TNR4iekSBGsADoapNhSunSwDOkjaEXcraDh2sExt7F+XUPQ8zpt8/rLxYwoAM84F
1Q9IWmpz6wdxfRO9lyoR1SQnKKgD0OuwzEKj9uk8hM0uPBwPVCFofi8RSyXVoADd
S3x7SXkoQiW8ycIKZ7R6S4yiGcfWv6Y28h/0Y9sd1/tQaVsnxZILZytWsXiVDfMT
ptLwh135v+t9z0pSwKexJra2U0zML/abBY2bji03089lVkUfne6NdqO2xPtNQc1P
yaNoo9gUNWQGpwR7Up520ASs8E2PHby9PVDwIqDLIMO5L1LFJ/7pja/RATFwHqMB
j4jlOU4GrPUlxG3p1VgnqCXZXds9ji2EBMDTT62FcxUSK6CA25pTO20DNTRR4BzG
i4dAJh2I2NbUsbwjWcyoJpgC9BObYEXXEaDcyDPrTeC6VdyZUztINTkFnda7se1k
tcdeowDuh5aKbjBkM447NXjV3f2BO5S6Tjxp6U9TX1vf2leo1Xo/XQ2e23AhgDAp
B8V3pgETzAVy+FNrpgsKenLaAA11UlN9vLi454VOYrMRJ1/VP4E1g1bSZC0RBB7S
Tb92420Q5QU+eTMHFXJD5NxzxIS0UZC7cYdLAGd3QUEQkMFKJD3pMagBC+fZ8dbm
z0PufDRtBxO/kwKuxv04yXbTKDQpg6CiwQ8hXtxwb1M0CTU/NhzjIOZgWMcXJjpM
ttd+hW8Bpfh04HhljtSJJ8rHH7gCLyRs1P8EOCw1ZoNZJAOX5aefYS9euqJyVqRo
65GBgepydfmBxkDX0FxvCIdcD9J1ynrMmwP2BpCKiQZ8+GSEdHyc410Eho/Jftiz
NGZCj//9IHDrquIRKQSawQ7JRTphrKPZ+akXteeq+sG5Z91TefDCYfKgqNG/bR8S
rQM3cctTMjoSM+nModowDAtYQzSrchLnt9GQT7OQGC9NDskv3rRF1ij1ejs8OVdD
Z6CIe5arPumBxgd0r9XvobVHmicckF/c2zSn3EWlUxIgj5hX39nZAjb9hklUvGE1
IQbImjC4LHAQiyhzmRfm49auaZMZR9lbFoWkPymhNEaSlFpCAeHa20gyRtLqu1NE
BcEwOjfycY+f3zuiCNpoQFSEI8+RFBclt2G34cfNUaNL4VjQVxhs2AZAdXXc2jJt
ExygSIRpei/CuqSayAC9pfIKfacwcfSRA0HExK8qEFYHmJSlpFpXs+GoRs9p44oZ
Ja9KKe0/Zg5dMW2HFPrRqDs6IDq1zYR65sB/so+EcDnc1CHORv1Gs7o5YzKvvAb3
3Nb6OAlPm/RlPKNOuNJzQE81U+63LrzEatjKpFCKSjcNx53HTJK7XGs4RuyIEmD6
iuOuShyIWIk16umMJJoCqy+PKP8uQLSVnKes6Xs13RK0t+DDdZXiZHGR1dj/VnJp
sLOceA46ozucT/gOFFSIEYeLRl16RdhcTR4FfDmGrpFEHDrWZtJkxro+V/zUBT0x
TP7ylIaJ7DxVMwD3ED6sLTXd8Af247aJFrOkkrLpN35HZw7EDfacBkZKkmyo7o5I
/f7qcVOYCIVCyswR4M6XXEgB9w1tGC+P/6m3NJRyOj15FNirX2nLs08J+4i9akzU
GrdI6JhtPyuW0SvlpdnsJUiA8FFJmgOJ7aYybqWE1XhYLAqfVP37BRMt9e+/MuXY
j32JX29VeaPCXwrqkNM5attVQZcbBGkUa7TDVMJgNtHLM0Xy7D97SDeDoHyg3MAj
E9VF/OBGmrv/StBKJXojSIggGQV9icxI5PlzQVufQJnw/M0gYo+8a5absSJ/SFR+
D8gULfniXngUwNhh2gDG8fgHnPg03SV1OhHl9/4flR4r9Qu9mOc2vQWqbCC0BMLI
V6d6+Eavv6fbs6L4pnHCjT7CI2GKKP7yXqZj/xsC4NM51q92ov2W4uvhB41eW/+I
ODO1pYN5sMwEB8AhiM5Vg6uLH39ZVFztjhsT4maSWnTXTLklv82zPBthl8VTu5oi
VO3Hcb5S1etRLDxNqFAcP7Y8+w3XIsKySb0/+km+PpnN6Zzmuy0v7yRZfOzyNZL6
oJdu7hxD7h6ORRR2wpTSL0m5Qjfi/UIk6xHBDReH8f0ncCBkMDKZyGNXTk7tsufc
0JOolkzcGOrCFnVGwSVhB9fxIVo3RaMl4QTZslDy6aKR0sw9LzAAHksb2cnXIhRo
SmFVMvc3cymqhEtVWWd0RNoFvFlKJ5slrVuhD+ZKr58cO9oPxTbhfhaIs2fC8JTt
06zbH1I8Ei0QDDArN3+2evmStEoEjITzIdd9x290yzZfkfgcmA6Pxf6pG1jQEtlN
0mrxhTiFgcJlcvzstW6fW7Vyxiivcgb8K6UkFGqpaNsI9fvjDB73XffP91LdRulD
v6jwlVFCjiXDJ0AWbSIVewq6ny1q92zDn9gn49j9IPryLaXqKw6nd+HunibKwIaj
n/wN+O+Eye/6VR4DAOXuN9mGDTcZSoj1vzGHohuqR55a6Txen3GwW5HtiznbGBzL
SF5wq37BxkrC2TCrIuxoHvzHVGIx6cEFhnwC9CtUA5GbRiNoKgZ6x/K7qTllZiOg
VFPr/qzWrqo9zR7xU5ZPsYviFSGX5mfQMV1zVpiIfcAt45Jh9aEQ1PtlJqr6FLv+
bV0bebDDea+vSXy+n9BbjFf8uqv4ltDaFBNEFj57hnv7TOHSYQWWN49znA3EgsF6
H9tDUo7ywucsH+8ysseAj1NPmbmnZ/1TWnbg43CoD0Y0AD5jgAdffFiIZfFPLVl+
5dPgoHuEnCpqbPM2K+9Vcyln0Yvkk1HIJobjHLI2Z+Aa0nLaLQv0+glK4smyuP7z
zoeQ+Rs9tQqihXkXrAwL+x4xTBIm3QLeL2GBb38ynwYpZabTP6tWAORjHlU51Vmz
8xFrIDNFRyqoEZnbsC6LosdicO2SXbkDP6/eFubbKDgs5ZimIhVM6vPrk90uARgm
XQIeNjZDAIcoOcHxcDH2xYy94gumNmp2/LTi27N4QeakcU0RSuspoJm8Hi09VuvQ
Ellg9ii9mcto3UFSnjGN1/9rce5uz0P7HzvR1O6UBELKfAj+HV2ry9ZNU+9iYa3i
8aGe+FnuKE0pUXYqblkpqxUbTwshqJ2YRMApABDa7KNKxe3YOj3n9pmvkPJW8GxC
yXWSlPkAAcI9qbkKAkeAAqcsvAAaIl3509nWT4ZDWFwEMTN3pL4NlaOrj9WzRjgW
3aoErsJXlFCSu+NN/840br/4gic39zrGCrYELMWye0aFbxnYlms4jKQdp8q0mFT5
3Khe3w6eireu9ODRILmNmXVta0Zx+LOsi8aZhJdHHUsGegdZhXi+bV24Z5JcHCdd
YG7Tjznx5FoFU/r1hWRvuALsgcsVKgOyIVxEM+W30FVqtHgkpPOjZMH7k6X9HhVr
eR3rq/bSKx63uuY+fed6JdmWRb4ZZTMVMWgA2PmNYpMpBZL8IUL8xattI5FwIw5J
N6OL1wCSW6rsPYHJPcS/oot4IZtdM/kUnDP4jJwYdfVhR0MoDhuMoe3ieGp6HQrB
c4d/6Drk6r24UQ2+he4L/p5mYjMzN2LSl+Y0ahikZUID4yC2d2ySrcZ7DPp1sOeq
b3euhvVoeesu8U5bbR4iHBdRJjEjC0AtD86joUCgFrDMoqsTsVCy1gLTBxEZE1ko
3sC8T2+tdB3ujL3btYYGu+/L82XCJ+5DBUx9wiWVFJyMshJW/Yr1ex7AUOTgcC6K
S2D1vsTq42/q8YMuY6WMz9sLM/GmtrS68l4wc8HEP1PPo/YS0Z+PfMiR6P+54bFN
b52Sv5UmRP6H4DAUCKVH3tO64MZKjtqhDtAIruHNX30y0ZsE7K06NVOkzQEgtGiD
dogWjSdkKoqX1PTxCfUa1sAGQjud7abxEu9TPfpeWufoGdCkGqOcRN9NWxP5TGph
L4ix0RWf8G9aJdnao/C1OLXViqHBC9a5L/8gqvfY+UhLVhP2n5wfcVOkFm49kq+Z
TSO+liiDjMZgO2r/PcrXytWDr08pmGkB1NjDy5dmA349L4Zbc6bMbFpowP895tM0
FolA/4N4qJLqtONYxCeSpmxYR+WadoSB6QIfPMb6a0sG2fM5cuv2O+f8M8M79bth
T1GTRDqvkiAyml64G6ifDecA/16sRCZ1CEnfdW7gNZ06VXyR83IOug2MJDbBLVeF
DwX6hp2BXabnjsw565qxxWIxacBptOm7dim6Ap3WDOCIFcqCuVol8fz2JK2GGuYR
/h85ouRhPwG8023DxLsNwtCG3ECasMxgDq7emTlohCvCHIvVGOBIXz4Rpu6x4Z1A
xTug3uUQ5adpvtIJRRDFgjBBTxGv6Mzqnu+bg3e615uIlE3MxD63kikA5rAx8/ll
Z9mKmg5uiCWqyT1Q8qpHYqnQqgYlhqOGc8YbcWwMn6YKZZm4xRYZBK+F6uyuBuBh
MncEAXUS0audIh/hGDvOqQJL3tjMJlqkq8u0pidb10VZ6nVHLzieiSOVPaHGFC0r
4cpX+ojt5afLehKaCsiu+BIjujKMUNCaLwqKpBCLEu2/lTzjsfGIrmbt1JLFNqRd
MF5oiPkGVLGxnCI0qujyo07JvRbQAvcoWTZTZ8A+WatywKsBQJFulTYXANb1/8VZ
rw6x/cO4Q6FbNOxRDE3w4pM+nI60A8zxBcEbj/Bod4BMLxkmjzZBCjoDBp/A2n9i
1iYE+GMXtytvGAPbcOAgYvgqvK3chcMr0MCq60O3/ZvMflsgIbqso7CCnJ+unJrk
CSmz5hXBrpF6gEcc3MgPcpgVyfxnWyIgwrbecaZnzP+HJ30SPvey+isc8QKDmOx8
T5D5oJ3GxAturjkTP3fWbhoDlIJBkCcOBEAuP0eolGCJMMdo3RmyG/53r2qBoSSN
UHjyUpMUTppUkw3ygW0RH5fPXUzYYYW5tYxtuAAClVyGDogkvZpu9/2aSgeSM/Gz
8wQn9t8aTnOfjI2CbgPyRV1YDRWN1gx3JpysLubpqZiZ1xoaM/TcL4IPke10KJv0
VnoIA5wZSh94mhu/ZJi5HyfY4/4zP5gGCZYvWp8SsSd9ni/ZylNS5wM559ARxtJ7
fdkfMuI2nFAZmdDmNIJzTUTzc6PAE6XBMQnZCvVyENm3oClKBtcJwP9UzgaDBzmJ
izRk33hMNO4QiVV3wqrnMWJUPUnai3twN1AdfmbFFCmXqykK6ApbUZTHwf64h0Fm
3EsqcI2SQq2iO/fflOAOwSCeJYsgP+/6cfMYLdha+9cR1Pg8D1D7YYRxc3nKUbsm
7+IT9k6zTQ+IDy5HkdeQDDxk7U1qWvo5IK7Lt0YnW7MrM0x3w+l6VAAtcR2Tkrs0
PuYYVtU/WsKuDAjZYFTMnl/46XbjAftpUQfe+53D5CoE2bks4g74pQRrv9ZVcW4D
q06hZV2/DntUACyS6HuBYRTy2XoCfmEiikiNtk8thsXQ1zPe9GyaT0F0HJvBK0YK
KcS/Nwnr3cNPbCUW2pEy5mRHDvbr8bYQ/rUoxvSyydy0dyfS8bzIeuY7QiXiBWmx
96PsuQpl55xzrR8KvEMmheAQT6NPa29W01GHw99LFH6Wj+uO7CtY9sTZ7MpoLysv
DOVV+7a7OApd2zz7utj4/Av7JTI24eRdoR3X0OkulDLNWXIuD6AI6mT5any6X0Fm
mOLV8EdpLj9Zy55aJIt2OjsY0IyKbIbG5HQboplmXmE8JNg/qN3srfSe4Gh1czfG
pYVadxXVZ4BTmH7GY+s5Cq16VOAdbOiTUZyt+XqnqZ4vzHYKeMDuffHLcaKT4h7H
2Cx32rADYjC27NTQDxh6had4O3HV62Rb2xW+cKuyWTREXyNSacCrothrAQmLk2BV
VMqSa3avVqBeMT71fzq9/yt8bHKuYzh2gyCjgt7IkpXdjg3qnlHu5vSdqYwZldY/
aKar64CI9rclPcqS5t6n6Z3V8dxfa6dKIzJ/xg1wYS+Vr1AoKiHZiwWxwBnhfkIu
cc+KnoMhUgwk3OH16CECv7sJ7M9/8InANCqIpf9gGmNuxLYZeWVsd+JJxOcnnYIQ
vJ/CHl1f+TzMx31FA9jcLKXN3jsIglwUKxFHYDINrf57R8LuJJmzpAbu2xpPi8aT
fiay3IqmpxsgAH94ejaf7twJw9kqm/1+1PI9byKYTigR2NFRL7OWNA+UbyKF0JuN
ma0fJLVlcXEN8XDbNg0vLqFDEilKEvnxCZ4+ZuLOiZCTvO8ap1lzWwVLXZ7PQn/B
hqHudhePSkn//jZ4HyYYSESjfCBmcZKkyv2QVs3O1W/3TUyQDP5zE17o3qCSh+kO
phbcZKNlE9Y5INuag0OtChvrsIFFW1WdBx2HZdrC05pffnEzfLjVpttVyXVpfqF1
0jJDFUmhCTxA39+IJlJ/GOS9holAvuSkSCe1jN0CihfQkrLPi1QgMTjubId3uUVg
+d1bSXhrJSbcT6aF4gmdp3Ex7UT/NN9tZ4PjeO8XM6ednY6OOu+e7lBqjhkPcvKw
PAm5IxmVXCadGjFELUzG7M0S2Wl+5ug7KqEu1k9jKKgRgCyAFQBURqFGOzzAZQU+
b8g2S3FwRB9uj7ZoI1FQscBUCkRgXzVOSuRnOpyxloTSMDaf3kvH0xNVvWM8Lwan
iKkmRJRGu6RJiQb+dYvyeddya2ZdEt1eoiPG8CX1y7QzLpBEIJvzO0fPh2YaDVyV
IA6UxXnc/927CFB4SWYtbUs7DH5ADoEKryQMFwBmsXu3T2h7cOGbLa2r/hZZNj9e
9hx0ap439XPnt1HjeL3K5jHLhiyul/fBExFdykj0LLXr4Zb5v34O0Y6jHh8lRdzK
lbYN1KhumRag5Aj2ZVgKcG+Ehqiv1GpzuQ6yINxUtO+244VnzS/ac6MlBmngL9s5
v1xfH8ZSOJWH3TzBFry4vOne+y3Sb1E0M5BesTW6DLFKyfFa4P5W5yCn2QHvb6vS
sNbLP0kWVxjE9VSllAIGvzTM/67QV611bEgDb4sw1YwgTV7LnoCQastnWRPY0to6
wZdsqMk/1RvRNLxqTfUnxWpn7p7YN5UrgUaBNtsSPk/2ODIm2u3v32Z1c/weLYTD
LOmsRhB/H1MqtrG1xhgrjlmAo4gGmMj19nPz/qUn0rCpCCrh0zrmDv0ovpVhWiQW
7VfmNr0SuDoK3v4y5riSsnr1/PcO/f0rXWEuugzRyrjiwCmcFaOSk+IwmiOG1/gW
9EmqjdYcZl4D7wo8sWJliRbzfKBNbU6R9BcqkABpzabyPtoVWFXxxdslaiCCa7T2
Q35v2qWZjVQTT87xFtucz1EZHNaUTaGDl5gZWbLU+/x+O7CMOqcU+KqrOfhuo4Jc
4qfcAkeSJYiP7zzFJX5JdKoUfBGzuoyPNPhERV6m8FzbChCJr+XIb0/sVOuOkofJ
eyQfGrwz5LSBRn9msyPoeZg4OBmVqqollRjD7na+IrukdRCSKH9lIJUu7As4qd8I
JdQxGnjRC6JfJ0Nu65pd9mCp6QqZ7MlBBANJEmM84L15pVm5xdMHD+mNQ6NdcrgW
3C7WTFTiYfOD2Za6VjOkToxTfT4LqfgtXp0ej84GXe11ZAy7/h6dSfjxBMSFOJFV
qVw7Lqha9sarG6WvpA0WrBSSk3ejJUiln4TEudoHcGHxsDWvjUwtR0Fl9LQaVqO1
PRzDoWif946ncCvfqmI0ccrzJrwfxZyHAK8TPhKFCOopYZR3YHVhXrF4EXgJ+hTt
05hmo0kd7ROtiBoDrK96EDiIci/oqUEayEFeMq7zBdk1V8fGGeo0Rzh42OkybcwA
Qn88EWE1opHwRKUXBPxAEY8Yfg6Y2yBunPysuTVrZiN1l2InXKqMuKMoe/+/OfZW
oNlfcba4F+D3Z3J+AEYbjs0YC44EKMaItB7SEKon+vlkzUcnV/yX+J/+2ES0tmWT
5LSLN2yFE5k9AxhNCi+nTO6ITAB/cVsRbhMRbCr98a31Lw+xuUg6zQFcQbRwlnFG
zVYq9CAAB+kDutarGU9dojCFxboVQc5GzSexI3CH2FrIDBDtW7tbIs4iMO3sR7+X
3d2CTP26d1sInjeJfejxdKVkpR0VmoeCmEul8e8PNNFXSy/ZAAN7+eJi3+a0RpUT
PnSR0SLHlM5XWM5TIUkRI2C53Sek3m5WOrAMkRPHEDO83BzBPiqpPMFSUNuO17ZH
cOMs7vwcdLF0HX8sYbkRt1SkqZnri7dPea3ZDXCs962+6ONKLkCfeQZO7C6CIdyo
yYvbeVZ84nQDKewuKbxe29qc3xF+T5GHbgSzaFIsXtBK88q8+TD6kCx2f7AYXerB
HOaUbM3T4ilaBQf5IAnNrpwfJo2lIuvlVu/kOfjAGaFE3bGYKiEFJE1+QA/pgPHy
yJYVTkT2GhBiqaUHSJCYHMbtuZ2nM42/HPtWjgdh/UPnCl+i55SXaHnKENu//B2p
8NXsr9BZwlyNMxtboSmBHPahkwKllTB5Aa8bcBPYATgXFXLumigIlded5kqf95A5
Z9C6pn3JyCTZyDa6gxtZ0iTX/daBNSOC4dOQrfxeg+h3N9hF9Xzo6N06hMilA7eC
cfMrvI7B+xTnhoph/CY4tT6LNIrg1c2IBar5z0iCAqgNed5O0Jg9xVclQH33vaH6
XVdI8dBQJMcKa5szL3i1OCxetOLUXW+U0eKHvagMYcGYCI7uKSf0FqDSYU3S0lkK
udsYVyUU9jGTNJG/OlRHUtVqmfacqwOJexYdX7Qla3lR0PxjVtlGwhXBj2ok2956
fJ+ZDhD12X6NpbuOuafrhglin43fqVlkv++dyYhUnvNwZLYh4qmYkemZKBVQ3ZRo
ODT8pBYLAQTWP+xsrazW1/Pwlk2T1RKMmgBTgIbDzoPPFJW2la1lhJkYOak65Jmy
j4GfK3P9Plpb98wMiCTZWh2GLOGoE3ts7vCzbMhS8tJQ4spA+sWW0aTJ5E87NY2v
3cerf+BAWd04zaNcZ/9m446U9EUInRF/HF3hE4YOZR5kqsC6CFcd55qd55vgAIyS
9CguJR306VDarWOOUWLVClgIkhTQGvljlNYk6qCMt9GjyYAw6LiO02vwEAYjkRgv
Myeac9JhAoUcxZsfvUH76yuLcSx+uJFGbdjDrfQTJQwqE/ECaBmgBDT8Kz5gGFVL
R6pDFjK00vJyRrW+toT6jcuMxOznI3aMSlobj1KyHu9ghBI3VZ0Lz3leI731NjfQ
lj/t+q5GFqS4NhxAFpFMTN91Um1fL+DtE4MqLnCsH8J86a6I+JPah8BT6RCI6q7E
e5io1YDoxbmhFcJR9iHbPTGKCb7+PYq6tLCJ5bhmLXvePN6dZj3nuRdiPBHfGwQb
vn+ghyun2kWgVtqxsw6TWxkOj+IZVi1StLnWvVvex6PH49B6j6OBpTuOQbpElhvm
ND52iZ8iFo4baLoRuoaERFtu65xNEww0VN5aW0uI7ZTzrNMELG/mEN4mdHt20LI0
1vJ1P1v+VjaojEF/oo3Beaof3nFNL2+KpWq7PDZt2wyqTK6V8L8LDvg6cJQ3C+xh
/PC9uXYzanujPzuGHjWgYvvUbJfvrrYquUbfXTzclzVuo5740ua63JWoLHWuJMMc
WMF1r87K8zw+4zzWSNM+FW0g+5IM1kjE04Gl73eqZQDD5NTcpBXkn3XwYHvQIvT3
nzG4ev8gCf+ehA32OMMzer/givW3/MQhx+YDDwHVq4EkTko4IZ2+BhwnPPo9QuQu
GKVVRdW9IK1b6B0V0aODgUilE2OHCaGqkfC7O31+8osOQbnohsoAC8dvRxmAWUOY
Er7Wba/68mnLfw4c2H9xif3RUwfJmcFUWBCxGqZg433CLx2O7l9bnQalKVVrgs6i
8spvf0RUo07IcS45zzAGeldn+IJK/i7J4guOHiBLQqmWZt8MjuAT2zBp/T1HAztL
vGsgzHNsqrYGEZddqnVuHlhfZbJIJy2+zGYKMT7BGdhyXavR2fugZLAwCG3vCC70
s2dQ+NTCOS8dKbpVL60b7HvqvQIoe0FDOtJhjvhWkVL3xg6l7VHFeTxKneE7GruF
+se3qx/87YOjxj0PusXo9MMwwKog8emhGL1EBSMTJR4iQ5JUi54HyVFAlv8vLGn9
yRXcOIBV1CKvezk/XQKj35vpx0W+3Dul/XuglMrc9+E0DoYGF82CBzA1oal/kiEg
dLSEYQwlc7Kbvd3fzIM/h1sYzCMm46EuvYuJ24s/Pet0Qe2rTZBmB4JMslI4t5yv
2a1dk5JgxR0AOGPezc/+zhqX7s8N8e3tFVgxNvyo1rDDtVnHMG4ihftUxoLw309D
uhRDuw6g209QkY0UUL8Q6j0GtwTv1odIkHWs1kMSAtQTvKrXzfW313EVa5JKBYNP
AhdLSNqA+LFSnFEF9SzsvJ8gKTboVeFp/ZiV1b+bA2or8+YIAscxgoDsRmOCLTBU
gGcaIFYtxRPbeF6mvDuv/tKp74FSTRXkeh0In1RKcj7w6GiwM61++1SEIJVnEQjq
p8J2Rbake21MD4Z9MZ+W9OUxsciQwNcop954SRzJNnm+kwuE74jLbBvVUeyfNway
oA368VJco7CLdtPFNGOsPwHdBWveduy3h4PFYRX8T87Ra+nvf4c4jrqcJGHSsAHu
KRCw4pLGNe8nBVvj31JgiSgxqjw/82YIVrlvZiVlbjBfNsghjqQm63OnvWQfMakK
1GIOMqfbQ/cXuDISar7cgwm7Htx0I+H//ocjFmtYsY+t5RsEgnHirKfuXUdYasBu
8ZPs1+pRwu99l/Cm44sepTipjxl/g74oi3SiyXbVyYP4qspcvOPhz0EBL0yWKx7C
A7ERoFKIM6KSPKnJmIzzDaoxNYUQ6EEqE8IYgo+UECaPYG6mEAWJBTjEtLZKoSkc
zkcwACnIxMyAF+6V3K6OphpVY4sxakf6Ik03Fs+PSigaIN/rXpdFMJ26tVoJiczn
xL6VB1TRKp53a0P2HAr7E9zp+zsgwFwV47X2Qu0DVBow/0s9eYHDhgOAS7EJJR1g
OlXsXMogL+Md8ZMkymP2jzIdjmDgYRwS/hoWpt2XY42Pnu3pnI95M2KGrcmOEwBA
d1obcY0DXNTU4HUKssc3/S2rfeJS0cvD7oIAlg3peqvZrVO1qyqxU9OZ67t6sv6X
3b/2dDlJcB9vbZVAImaWN7/BZHIzG6XbOd3UiuJDSDuKGPsuisId7i+yJq4SAx1E
RfqRZrLHR7nEu5z7LPBUzYRIolJnOKelFeiBkM+BdIcKEUGwxihL/3zsqEpXLgIv
bRyaQUillKyq5egND5vW4GqxOkxYuvjrB3dnrWekPsDB/YB56XOSlnDS2Cn0q5s9
ZCJVlHxPDLn2CatOXYZpBrH6lem1RduLgZghF1iTrCHNgiZgadtumR+1570bBCzq
ERrNcCGrnXRhuaKnMNDpOWDFqxcM/ifyFcj+Vz3Y8XO2F5RzDDpXxrskMZFlNBDv
32A+uDZxAPDIquLLv+32Cjsch7MR10mHtWkNQ2sIrFTkqfEDAg3yGJTZGT6PYCh3
AT9X5YyZZRV/eueHshYMAX+mso9aH0VHzQ3DQhxjc9qLg2ueRbk0mlpQvXi13Y76
vMmkoeuZ00kiPDGbni2LoiTJMir+hm6PFBZZ8Pju/7PxLMez756bCyjtOPX//PTU
erEU/aWpOxa5cXUVLfKL/kGb1Cel45MujRCiDUs7HRdiDERhWAbueHE7CCfv7pj8
FZrXvRr5z6SXxAAUawjJnprVVCSK6pXH32qE/fDALYk7SDSA7vrOxYESd3VdjdHb
DEQGcghq6O2UTaJUQ0oXljbl0Bhqf43bCN7bHECRQuW43bqWNgADtdegvIlK+ibL
SUkICdXV8N5duMPt2OcNNGUMF81VQvLhyiLUKDMaorzgRAAM/xj+CWL8Xg/Hoy/X
qO6p5Wged3YQPPyN4n2Bi4M19p3LmZOGcep3bmAscuAfKhTdFmNp280Kpe0YMUhl
MMDQFAb6NXTdJvEAoMuIP4vaP9vjHXIzhoEcCbYTq0LCkSYljT2JOxSvMXh5Rr4I
GFlnYC1mwtpIA8z2cvMKmTn7K2Q0wO6xm+NMNPAFkkzxaSv9OLRyojZYbiQTQAf7
8xMViaFXromfhrDht2xWNkWM4QacgaH42uc3Dv4lcK9K3Wbi9g/5QCoKUtouqjxy
mgPEA59OOMvFfzmow1VbRwfD8Dsz4Bo8XzZmOwvCKsZ5Avcsjxq8QB6Yrv5+sE1q
TSIBLe1AwCTNzlx4YIReXf1DMScQMI/lwSmiLJ8pIGzeavu6wfgerOaMfe4CTPrv
GwXwf/usA4TjAnaOAS5smyKio91ErP0kHRUvrZUw6XtJEjFB9jskZ/GIpbgW4lrM
V2r5r3psoMnwiLQ4pyhxPI15PjzIdD4i/67NpvUZvZY9qqjD5BRwg6J1g5r+Hd0D
IDdDDWr5fWFCkQfB4Ug+4maErkBQ6jbRrN9280jJNjg+lbGJZ4EZpbep6wwbzLRw
iRK8bsP0p1JPpQzvWWuE7EezDvl0n8FaQeuUyA8x3I84x6GabALh7uizEQN2+XL4
7CkvycY9FhqtxjLmxwOY5hajqIsQiHC1I/h+HmF2MI19vSLumW2+82sfQ+dUMdXj
1OfDE5XMl+WQcPeHESDbJEW66eMtUap7DYj0AGWT7b0HYi0YcmWt9/VJvGk0MCsb
vffJCPY3imWJbBvSqs38mRv7cgWCAD87SQttu4hG/k0Vjg1ZKDcBXO/uEpEh6/RZ
3M8wixip2yN+9BW5TUno+ni5En4b9ejpJHQaMLd720y8wBU7PTUWFDLGykyHiH9n
kNl0AWFoff3Kmm1LaAMPYUDpMsuV7XwAPLawSf/lJhBSJDBBICdRD/ZzjF5KH+ID
nYCHEtcnGgFCmlxdMDu8KFDMfWzCyKo37edqn/aCxRSX90o1FkAeUVePtKBmbPAm
xc1DR9yXRxycuphLgS0GqnTkA/q0eUgnG8TaqOv813r1mJnqnhuDLtqiTdDG4ym1
EHKGAZwLwu88SIMuVncj/bGb2jeXaeUL8dMGPEO2tjlj/T2b5nxBHoVnpTG6/aQp
S+7qnVUIzhE4YXyw5P5tThhuOiYwFGL5JNa4qjV6a4Me7MJZ0lal1dlEMcPLQOTk
BNttV7qCpM0MvnEuPKIvKoFeieRX8/7wIFWYLTRfkCT7GXa4moxtDMUdLKf0+52D
q9DF63xJPfV+FRu3m33YeNjQ+vq+jq7TiOSMrEhiPE9aJNiFfuO80JneKzyP7TvV
xfQEs6IbspDy8NNgDudXoh2a51IBxwAh5clM7mlDmN3Cr7bhgE+PhrhMaFv42mn5
ulfLAQHC5tHcNh56B+5g+0yfQ/gQPu0AOP1/pzUt6uYhK+O2yjbrhaov5NfNpZRB
OUtwJ28A/DG/rPw6la15Z2/03umOVehYZCesJv+8tkz4OELDPHmxPmnDfDSS1f8o
ELSovFOrEiUnvadaSDK5fkBePgNrIWZB/jphFZSeLLTG7quLltxrEQucqZqf7I4y
3GJ1kxus4fHv3y+MuICzt4gFhM6Lma4IvbMrJNfwYcUUFfnwjavE9PwadqSPU4AA
SlfFn6X/5vZNguwkWPW+YmWGbrCGlqRaxShSJ3RMikjzH9i7MXOalcTgNM+2Dm0x
Nro2MEyo7uC8DYfhUzD8t1QW+rcD8S4e6YtBHx2HYL/vQjb08p2/tWIPCNisrXK0
HFZo51LNLdJFRC7eWyifmW8lj7Wr+D/MvGl5fmN7nDoteAKejVf3ge4zkCNi2VmW
0xTh5fBP/Rh77HbsTa0KGoWpdsHHh9sRovkZubzNpxTir1RAoe1qFP4tK9dscpGK
A6/quxYJXJmcu1Tj6YmNuvjd+Wq0vIfJUgLyl69cr9ksp2hCefb3cApPotC5ij9s
zs/9mHr8l6hc7bEYdsDAg0aoRRNgPYybw/mQYZl5JCyGB/tv9j93uQDQrKbCnVVC
9WRmjnqDZScR5XZDnAg+B6jDjPpwa9cQlhwfAjT0TH/fWN5z4RKCiXyHtJmjmCf3
+/vYgTZlFg1GmwZCh+HRY4xHN6aaf1eMATLUNCDg9NbiK9KAcAZwAyjmxb64wQCh
r8pSE84+8+jZvHfnYwksIxSaiLuR+eHdNxAa4k+SmMPa9Z/+A+2NTuZrP191A0+b
OfoX8rZC0rlcBjgtBOxS0UgoxsNKyaGspnD3kyaweQ0EE1NnvhUqlhIgSexQ5UUF
T0r7ufym/Byj3aOs1sMDmmWJ5eqeUXkU+4PTWfGdbgmJkfvkJF8t4D1kGU8n20Io
+2xEyWAhyaWKotuuPVtRY/aH05Imd5kn9cfltbVb/nYVoePT+dLxHEZdTZHUbrfj
0IxpPJQUs/gnr1vmG/fJWl1JJZMs3YDO8UMoUolSSb4/LAjYW072giz0q9/AXHLQ
0SpwVftLQZsXClIMIRTNyzZM8CtrQ/2TVXSa2wZqjFNEp4/+jomsEKrDCgAYMQHo
iitFjBl1VJAJOGVH9/xSao4g9KZczBPwx4lk+gfr3WohqKqP/AXIpycQHPVxWyTG
DZnu5z5cK1iUx3mUdwYj5Zup4QMhkX38BUZUbP/BmrPIF2YMYxmelJ2u+SMYCWJs
WaEKWpsCNNiyhRbbsQtet3uC0uLxrv5q6agwNfZWtGkWOXsG83VLVe7yBKCcMYJu
/NELHcK2P3Mfkhej0FGdQO2/71PRs/rnZWyKaRJ37GTIQGTj4fxoKrxfs53xS9lu
7326ouwQ515S3+YnvvWrM5396QF022+tyXr+GmD8DSME06aW8UPavAe8y80m/sY4
+ZIMagaXV1cQUJfjBog4fcTXitphvPtHYRNxj4arywZQJxSdr4Wd+Diwma9lX5ab
uNo8xfgSLrOcPmNtrkeXTmsTLi7fy8fG3ccm8EVMECM9doTQ9foQIKqBxu7Ev5xO
l8Yu1HK8WtD9rEcNscsCSw==
--pragma protect end_data_block
--pragma protect digest_block
LVXSJnjpT6hiTDVYD4xrVzytIaA=
--pragma protect end_digest_block
--pragma protect end_protected
