-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fyJaDm0321uRUfSfHt4QhRD9t0m6BRhmumeRjjT2pljSbylMUQ4Ns0uwFU/t2FzG
C0DOkpOPllKrgtnYEbQUAiyjtHvWUhGpEYO/Pcywlk/EbqUB84xq062+45BKCaFP
QPoIUvRPnPKiq5npgPw851ExOCbiPV4RQwnnfQ5kEB0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7417)

`protect DATA_BLOCK
rvWFK5lp40Przm2JhMq7nXDIH239DuvKeMKnplFJrzrPQJB3DE4RRZSnb4UUm7Cm
7QyMdlw5REE/IQWlofDjXOQ9K1LUpbj/0BwKgvnWc/3TJ4hizowHANwK3eqwcesA
RsYhvNfsrqe+D7y9KYhKCSVDIq893rELbBCAq0+M+yBuQsUPg1XmnXWv1D6ed+kQ
MTOtbSkRYY5h4uQKbeVdqu6N8cPfS8AzxcT2vjCi8+rrm0Zfvp6lK1IZtz/Y/gOS
mV0pH3mBN0I7RnP48nZmfkvUAwRPSBh25wmzoBnwjjvqCPhbqSOzwIwFporiZXis
Et0QsmZDpiWmXQgVaERmSjFvsT/Ydydt4szLUqxq2CnjHTSSyTCn5h8ZbW+agEqB
8Zkf9qgpBuaz5gfohu7PXd+GsXl3Veb3MxZ5DuOHVGYXhnroIdIGgX0ZVn12O3bw
uwPxCSIOwyvo57VI5nT1/noJOIwS9phDCeiRuR6UiAunX5TGd6YUy0kOxYYithS3
YfmmACJp3y/HqHggF+duGhv42g4sVe5cdgfvD5F2IzEmjyyVLewA6EqajpQ1JjYo
hgNS4dB+Eed488AXiJ1Q1krME6FpYMnziw3Cr5UjKEnWqwHG3KJbIF0/dfo8BmtC
fv8MYOyOtN9XVdm42wl5TvPhdkSHNHKvZJboDVWBeHek97LC+tBea3GcxTOwR/Cx
dul5dVcTu7zxDJY2DxY/xRNS5YdYOdtOQLEgcFbo9XqUb5+v3jajH+h65b8gdV9P
8+hC87ZhHQr2Js04GQfPV0lIX5AhZ2zS+EDVr4C1DLhJKbKEClyImzFRQRI0z9ZW
omniZ9/R7KkAeI8AQud8b77ySCS3joGTI6ZVpgqV9/IRo6UFWV7vXsJrxUjKM7tI
QjrhFUzlApy5ONexVUPwEMt9HuGXu04nITWovWXwQcAftU9Uj9NGxH5CLasrBaUY
+5THK14wagUh2+57jH45baPkypLyMTuGk7R8+54w5rZDSewXBtpd+kT5lrNX4ALo
ECfSQc/ScF5jRaULpbEGdUJWvTFpXaXmkwVE3Md5J/HTtP7WvPoIGuFmK1tWUvho
CADFZJhYMx/bRTmirPWBEPZfekr3TEwpmG8MnJ/lYrvZjcw2NhrJNrSM2OBNMsD8
e3ayHVdKLX1hMDQUknGa/yq2IlcZgXeIMEMwH5fvqk3zcAvMA8AGNNF5PMz7uoSa
BjDHmlalZs5BFOYJRP+WDPQigE64hfnXdY3WB8j0UqdR0oKWDID1qbKpj7mEBYSc
rmgfsg//dxX4nstkiFA4QsMgQAcsspkfhhV2MEpgYxmsbCBzgIwqRftw1iLwR6yc
WOv+uxl8QSQSGoXiNLZ9v4hF2flFRn5cTJqvSK3dgslH+otEB01cNnGPi1tiQ8wa
g4aEFUTUSXpcUAYbCsRYUaNlu6xLa/VXtOPLfSRjCPJFHBy/EqM5FUBwmEe4bgej
pxNaWboCAivKaSaTnTpiqzks8xMyB8wfQdJk3GrnmHyZ7HAwdOpxmg+hBZVYwVB5
rpQjfnu2fa5wsPPYL1VQtjAxPPrYgi8kj2gHQXVNrSZbwZUliFXUYmROlAxUi/6m
1ghbNFUQtQlEwyeOCW7TLecMi+6cgdb1EQHYdnsHiGcmGoOxHMUBR7p5XSoklHwl
T45M2coH1TWpbLSE1yJjmOBgj/DM9axn2AoRthpYxMy5SvKupUil4iTPJclxVuVD
yQsif2T8mPKiRRKfHCmZ1ciZ9VIL6naVBCZmiZmU0s8p17XeJUz/ACoEqn5Fluyz
Eh5qHePw4tl1LzNH2kB9Sf9Azy9oi4+Otf21FEZzm8P1FUIeWLWHXOdUjDqZ8Qqo
k1170SF/qKYLVyxx4W50BfjIUcmBaMDxiXjXde1mbwHCJmRdUKYMQFpRnuRJAQbY
SiWP2BTSTSty+3l3kaA572OQmCTW5cyfoe21UkOdeOY9CRZDqvEept6HgLBLyBev
B32I/PshJMAJ98BBxlHXPuW4fzienZnFPty5N5nhkxt1mzBeilyIkscSPEoQT+57
wLkczMnth1GLa36RpHa3l/7RQsaDRap5w3ggFRDEElo3qvyHLNBzN6C3DXQHCBPJ
hE6jKH0PdSi9FCtfk+kRLh8YsUXX23eCyhLQCinpJb0dBmWHBwbzYZfKc21Z9T2/
LfLQzHDhWpo2/RygQBj1aul5troIPVRrvS8jqS3LohpuIGJoa01HMooptV5DtJYZ
aCZpaPpEV8iOD7cDSCrpkO/5+rwC8UkyPC79+RNGG2QEpgYti88EXHYUKK86YXhN
Du3Lc77IoBcDwBHyHgeWqxC80qTJ7AuOrsXmtfDEkcS01vGwqOYFQrUbMmpMMbC9
xf8pxvPX68SHTVnDQy2uNt228nVFYdjRA4NKEO3HdJ6YsXssBxTcy0DcRlLFCt3h
rY88LolLwbAGP4o9e5TxJo/tkbC/itDGHDCcghQm0N6oFpgxr7pAUi+tJemvby0/
4KlqUk6ba51qf4sa7HeIJJSUYGoMxWIQz1Mhe+Nmpg3yjc4njQXOrLcGlfyCCBoi
w45OpefQrN9uycpAh+nL+9BoBQgUcmGhYsom6cVo6r9UMcieR0z5rcezJzqp0Ok8
d6czmuHfR/A1Gt4ujUMDwSaf0ZwLw3WQ0WFqcRdtIy6ZOY7Ux6j4eznG5Ckd2qLp
SWsXkhBbGfRwnZlJZFeYzrzOwSLLeaQ7Vt2Cpuz5hm9jabcF+6GppttTbSfhgyIh
zAzN+l0fygllJlEn/F4/bdEXp0MViC9h5X207tB5UrFmG4Ly4k+406U2zmFHefzU
OTf7F2Ee3ZRStTrMxZ2bRJHsorj4ZhSLFOQNlx7SOC/SNwezpTfj0mLGHmRWyZHy
Rr+bvnRtjfa7Fzrgm7q6qgoNX8UNCT5R9AgF6jAJgVYpBHXLBYiKyP8wtmYJlkeV
JCMtCjuDVH61+CHcreJo6bc/ie2Iu0F6cRE8qZifcwm9unEpDRfIB/+FwWaOmy6N
7nbR6EFl2Z/6kTZ9PHumT0k8wZXFAXA7//TZ0adO8K4Djkaev0JM/gcT5GqbSqzX
jhfOmXexNiOr9ooXTdiaGlkyeC9spiuRZeTo9QpUTODVkxXbAaTi50owoVAMx/Sx
9ItKA0TGLnZ50iVrz/Gv30vNDihHBoeim/PoSthdI1fe2avl7viZbQiASTd0eU4+
xvkNMwSJsMJW+Y6DLdy2Or5lmFA2LBdlBBcMzQpU1jGdzJxP3eXudePP+8NJ9nQ+
hNMfiRsGM/nHYFQklokjcpKnu5yeSs4cteSbiv0CZfFASqYtxD5Y3gLHYJovC+Ox
42KEzrKcRJgCheIYhA3keGjzc16eRtMM8qQYoJmRw2AsXU20HPc8/qpmKNR6+YAr
W8Cciw9z8TpW4CGDmySmG8dChCVg67AugyRuy7NM9rZHmk90y9ZP2sYN0nNNdGMh
4VVtp531DAu16oI3Qqh//zmlM3UNo1NMgcx5Chn48PSTWPz0TZJhLco0/dpv6g9N
coDl8eS53FO1ciovlAUsUqLZtXr9YHyNS2gnwMSpp6w8A2eeVQjJF+Fi3cZlYaqq
s593QG1PR4Mtupd5xQxaOlrkUyieJutMdi+P+XDkAsp1L43xRtS/FgWgPjmWrB8I
aE1DuL8JR90t2t7xh8zZNEF0/unxDNW3Bg2nXhLtECSrkG8Q8xJtPUMGhwz7AlZb
CQblVXpro0cYqxPXHJyDq2KjRIyD2YqNUfFCiSR03ZROviDfxbWm0gGb8xz5DTGb
piokOahjxE4NcPsz0dLY/K2LI90KpUkGtj7odb5jKThi/6frqkvU5LY4bfT02iDf
riEvNtOFrSe9ACyzO20OIzMcLE9jpswddgoMNTBU6vWmVPsQtKZKIKGrsnbsSArF
rcoEwgNESPMn3Vz+9rLxz+EDxxf/FVubBADNXXokl6UKcHY649ieZR8p+9rBPiV4
3MOut5u0XYx98wNsqA9qDfAtnZBpj7HQSlEyDA8ngQcjDWA1+rN2p0/lsU4uAX+C
o3UNjfula0pR79tBkaCOsA9I5CMwS+F9S1EZu9J36gyP4R4Clv6VKamGraoI79FY
qLWB56qUa/poYrrtlfnH5LcrRbbtGU1nlk0ziDjWEkqIf1yz1Xk2EMbnI4EhohyS
w2tCEAB5xXPbRZnNT0N2aOFtmI4V2XchT8NX5bjN0O8pYu7fgkCQiNST1V24wEvc
OFtnH3jS+ElgDTtP3/vV4bbRDySHGCSIGdIPCgVOnzIkk3RI4qaFjVCgbAmzslUn
m6/peoemsu8f1RmoVX0gi6Gfa41SKM01JEfqOMazTKK/drxKpitHJ9slqXaNkxwR
lfqNNsYSwgI5yGsGIcXK75991j0H2drJ9klsdPRbPoZwGqQpIquUfFUYPQn/6JRW
vjfE1A/oJgT7iKVEJu1+1hMjeJFapReVlY/TTEq8StohWna+tqcKqBNDF7iLwFsa
Tpelk5NW2PvQNApBEmCc1crqgiyBFZXQx6CYqTE77KOtS8qKz64YplRjUa2EVnzt
8wkCya5RN9v7BrMmQvEujvdK+ccTNUnzHN02HWvwemwoiK5RPtE4Wf6OV21x6mA3
iaTaw5xbn4o14NCR4/VKV5eT7/cF3KcuFmPrkjieegBuzTh7yWCEthwmYheuEc5R
PuwrT5bxS3YC2+3ofpcDa4HJZQMUpKGcmX3YhV8l/SHthuWM3HtlrhgIhp4l5AIJ
8F/qyGKePISJv/ej6IfvHX4CUMGfZCx8lPFdtv7Kq03qPDvjqShFMTk8R5be+TR4
ivcn8xF5YE4YBVzkBwL38xmt7dhu+nLVIOXF4Zyh9JsgXnPtCJIa2y0HmGzysUbJ
doUqGhXAXn8jPbGDW+Fm9xBhJzoA1R1oLQvy8/Bgs4e8RRRGlqn331cb+wHilTqR
cw6Hz6cD/gaJ7UutzR7Qr8yGHWIJW8oJCjsW9eijS7PqqgJXaQYpulHzBbbELU5u
0RjkyhxIAHhEGsD2Gx0nRnm0OrCuctgvoI1jZM1WqUNXWCJUlXlEmWVFL1ov+kNV
pCpOoDH2a4KYkkfb+iLrkCZGWy30OZ+1Y2srm+k8AdalSVElRmjqOsFcKMWpTjpG
mNp3jBw7zOtAOnRt+m/CC0P384UQ24XHRRSFDs20ZHzrx1b3sJ0pu5f3IBA8D+un
EDFnucpp0TvyS7CDDbZy2Jt/2vBkeyo881U7IfVh32dEWqtUPjnPlOlSOMBtZI26
bg1DvIUFrCgtwyvDSvIJs/r1V0KntKrOjDEcLL4j23+lD/snmCMDBLxElxc4TKRK
u13kAwwyCFrOlmrmYHk10/qvhzyE+2m45KehqurlRqMPc1HoMrRVfTSGexZpXMFD
am17NJahfknDUGIbNZC0jMzixT7JfmVjzW95EZLPRV2xKMWWIYi1ucafagTd558d
k5sTgXHuLYlXrMvsX6moNaK0FlqS0kI+3OBQwWmKrwiKyR3Ipxau84498c5qjbmY
uwMtlnHtDP9K1mTiA8sbPQKYlPNTrnTYHSWILqhluNCZIMQf3ez59GRLv6ckMsDY
pbsM4uaL7JDaYMo/SkG0IwuF36HOj42jaKnEM7Dg0z+PTeqc3WHN69e0/qES8dMn
SSQka14ICjQDfRztNQRKo0UO+RiITY/xct75Rn8YrAntTaZM8vG56qVDz/7poXo4
+yLfi2qMeoEzc9wh3D41G+QyfrBcNJ9kEi5sNlkJLht+2L+HV+ow8pYvHJ8qBqcE
xOI77+QrfV56ZL3EffJKwTR03OA9/xDiklCEk69nSVPkmr8WXYqTJr4bQkdQhC1w
ZZxcaoRiY/SsApaYu6Hko7MyKctSa/m16s8LiEIdJXBGDbrXj2qsTwHwBuVcadwB
Cos4Mjs/4GuFQQVOQ2Cy9525G1X05TIKigS2ahz6PuZf8BvSw0vDQrOStLEAu1rb
JrdJXG+mvWFu4MSFFqqRYgPQCJvuP6qcEJroABWsrZqjIAWyIJ8IUTyshzG/gR+J
RLnZLy1iZpq3OnLTaqFXJS4/7fqYYW1pSV1A5QQuirNL42KxVjfWA83o5CEclSbQ
KPB8G+3RZ084g2m++sRBcU1oOsSxwq8XPT0ace/Vkgu5xcRK4TjtLET3JWt4kmRy
o0KABIu9bsOdj/ebkhZCBKqDfrorL6eoLeLgqOjx1mrqLwF4Wry2fGpzhCiif134
9UcUTE4aU+QCqXt9WUIMYJwO7068JgbEYl6InyAIQnJnh3Y3a35wSHiNzRmJ4NHn
EgHNqatgcC+Z9PJPztwAVDLlP6lBwkUUtzLBhTyJEgXetnZvqwH/l9syLJxSlt/0
3YYt4sp2p4Luiu0aik5PjLCBXSScZ4B/u2nh67sBqiG/J6EsxHAQSM6McWpLhTdE
wMNUhcYLYPi+pTVqgi9zDW35va8SumRP/4NP8ZrfYKShwwFzAA+CKsM+vD8e6i6b
otCZgtDOMnAWiPyEciOzGkkkuLKOTP2b7o/Vo1dc9R0FSVrLXt3/D34Hz+xkQWz6
JGAPvZ8H8XOw42BWnwbF2kMfLHUL7nLVfqgOKdxnAOb3HTJMhwNjhiC7TM10y+tG
mbPsssIPWFeuIx9dfpmojzzTT5eg3hoRD3ODfThijx0CxWmwNO83z652G6CLi9KE
bsXpSMaFCLE6oTfiZOJYaEpN62WUmcK7Np75cnAqj3tO/L80Fnvo6LmFDguYL4U4
tH+mIguHawP+mCAya/LJXMav+4dhHHOPJq9MzpEpGzRuq9XuXCM7+wPv2YSc4jIJ
8KY6BbGbQL3znwERT0o7dagGd8iLjtWbA3eUNdyJJ2mVhno1hBHna253ZW9aBMza
vFQ2s1icYH0gNhuciodGHY7gXpei2scwYsnly5xhPBf+8HG669yRebKO8RfXgbxa
aWXpNkeljqRt1knPG9A+kw2ID65ou8MD5dfoe3ozVQWG4mdaP8lmO0sjeGtJdAwH
0DK/Jj7xN2+8jNnbg6qz0dtycEvYq4NqfvxrbXA61XPwSpxS3c8FjOVkiu2uIx46
p63t9rGmTb/1kxisEhQJJFWV5pwLI6E7wKlq4g6kToIIEY9dQAwuj06rvUpQ82cH
B5TQzBgW2f9BUDyjK3eIwV/JQ9UdEBl0FbailrK/6KTU3x4m9mwEHTCYW+mGL3DS
ackThE40G4b8KBulsJUXOvThVjF9WYrXwLVbZA1FL6+LScYbNHs+g3vZlvV3uXpv
19NN+2AzYE4MZ3Z7JeHMwH068bKGDXYDXXYspHDrQqY+R4H7WFtqXkuhVxNb/FW3
22rShWR4q4zDFMfqKMgyN2cSG+TsLpAZTGts9fYx57PXhO1pm6rISSNUfathcLAR
j+rCZWNDZMqtprCdfiVeGKVmut5mDhPhk3J5SERfdxSGJCpJugXogeURyPVsqSM7
tY+WFp2tpuQui+vraUuIOiA13+DJLFscNTbnTjJWXahCUc18paUwpdxF2vb0SFQN
UbVVwv1x5td/SqndwunbHVGeEuWTI/AXrTK0Lo2KBycn9yDcLdwAPIPqVpHVW01K
jPMd7BG1wR+MmPPjjV1nzaa9i1jn0Gxm1tUgKK/lem7Yyp6vyofSisixsVzHVHtV
P53ehgm9gOnwMdPfDSwpyobd0B+LF6+afETyUCzyipbrLmn4+bWOw+n3DzwZOYwA
eoER/BbRHNvH2nXvnZrkVdvfT825yZGOfX0OvYd/AOCRFb9vxr7nr9R8QLIvECi4
rgkhC+n09MOnrdpDeBQlUcLNbCmjq4R215IehEUmsG3QP5sa8TkHqhfzZWS31Pfw
8hNd3sNdEAIEkvaDG0cuiNjmFYAER/QFIll9LWJdWdjeVsiW3jM2NUZ/0bq23o+u
jtY8LAv0IcCXK5BZirhiNyO68YGCKN7g5vTwOfMsQJZdyFNtUFq1FK3FfmXInEug
PGPBfUZSTTtmqRCb5YV2vfhSeBRC/DhTPevL4sYkRDiZj3VN5qFhJLbZTcNifXYC
0ifWNihhl9woXDgflX0g3pzddA+qVd2iLmqRc3VXUhQoxsEqVjPIVWT0ZJEf866g
tw8k0xnICTQptKlx05RM4D3897nITNBOdkxqZOP87/W3hMw7D3kzvd8ZcBYaVpv2
2KeG7qnVb4CaWn9G5itQvqDxHQEceCRxh7A93S5ne+StxFefYEUJ3RDr1X7pjlMZ
cne7ag1EWDRluRCjjmugkSOgGgr0ybJI5OPXcTmLZ7wZHEi/efaETGyo53ghX/G8
a+x4ys52L1eW8v1TokbTzrI5/ARxiUOIgf1okwo0gUFsJw03s0FOy+cWCZqtzLXJ
5qegXyJcuTeDDnKi9ajPryNzt1CYcP9Ojbbg+pYg1p7n+fx08D0UAENegb/SrF+v
+C1+ul/cVVirnh1a0tt0HzqJq9EpC+gGDGmQ1HMOzlOcD/91Yr/eqARg10tGZjXH
hj4lGc8zcopVOqrpdv2aMK0VUkE6VfG65TUAIkRI3/MxUjzZEELbwP3sgnmPHw9J
RQ49DbxYGZWnncc3CUaZ9d4hUqDTo0sugAgf/af0KAAGA/ChVgklGQ3gWTUQu/FK
53BEpE3fcXs8EcoVl3UCRjmlOnOK6K0MmlCt4olxzxnZjlwPtK9SjSYiSXWehDQI
r81q3dB3mWYR6Ow5Q2ShvNeTbhnObK1STToLo8YxWLTmM1NtmAuP2GylCaFn0Ig7
5CUZ10kmkjenZxIJenEnefQigf/UGHtEJABREFE0S2iOao8d56bM9I6FY5cQtI56
tNEql/MnZ6QYeCaKTFv0FHdDO1gLihTKZDJ5m0M8fHiP+2e3nXWo0WY4ZTWIq+ba
ZOhvMImLMCVOMarL8q+1XNzpO3wc4f78TKzgdqWWflDvaiZq42c2KX3wlL/u8uaM
ZJnGGowsaA8oQkl14awf8Um6tuQsLFQGNvN2Z/m18W1bOTlJHw+anoo5YmW7P3f9
FJbmHk3lu+9aKuuDNf2Jt0n9F3su9b9UYjWbb9z8aLNCK5AZ0TSo7WKRtd/+3Ufi
nMaAXqr6BnzU5VmRDc3NbQhG5GnGJ8WMJ+lHCckbRT+B93CIC8Lq3MYPd6Er263e
s74d1BtRHR49PbZmYDGvclNpKeZlBvrWKbT2e0fgRMg0lAGZ4iv4xn3IfvBX/5tP
knlUzeu7u3kGKNLAPnqXizhXYe9HmOD6WdoTKxON9suY5eEZHVoNDYFw8vICu6Vk
TXfHp/xeHXUQyoUp09lJ5qZkS+tkF157DKBRRkR5cFUyW//z2bEImFm5mQJXWxBb
QA6Qu9QMmhY6YU7av+QCbg5UXAPvFkAHIdSlZMcUaXVcjCjrdbSiyn9BD1ppdYrl
q19wYn+80gBfPOWXsNsAzRddh8Z+qID3gCR/2Hfi57ORvaL6n2uCa7rwdQbBpyKg
tVvWhidNJWlUnblroUArl610Xyh26GWq61TQ1qChNDxh78VlaMIxodsaqqE6Gd+s
VC/1gBn8NL/Ib+ioELph1tiBOav5yC/9TSJEBdyoyf9TU/I1+A3ghIM5n9UFquKJ
AtaabkYg3lDCRWVlyZoBgRnB+9uwM6epcMl/SamF/IAQnmc59S2wN29DIxlmw/j3
Go3oS2a++N+ZuQ9GFi7DKpvPDtD2I56MXce/+sFLIvSDAo6Mzeb89Mr/FkrtDCen
ZuH+y4J9yIBl7uX83MBjSdvkd/7aPOcgdrEBCWq2N0X0N/CXGqsrsFhAEWSOCLUJ
gZNMK7pYQc+BeysVinIKt0N6qtIjv2vuEm+Qn7Mtw/DpOxHHyQ1GIfH59YhRSLge
f/t5BPy0knLGdUuJbBXR0MEIzxhQZVH/Z9ijRYG4Nq16/j9efkMTEXvZ87Aly0WF
HHzBnQ4WTZ42EaScmK7rJ52x++szl4SNUXlZ+5RWRCgjon/SyaIOa1KeQmmhINQE
`protect END_PROTECTED