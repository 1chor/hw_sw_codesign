-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dMhRIDFnQs0OIlu4vMJL2rQfbBmcseEK+b+XdaWCaBIAqrgblbsWsJ6ANKjqrxS8Va1DRZL3VVRJ
4qRUJLsfqyHMUvG65+Vqwf2MQ2GXhwaiuhrhe/eqY6UcZMvxAlHjv0qNGCGlIbuD24Fb4JYgeUia
23WEpt01uXQfpGxNgJrr27q5V76SIkqt0eN8xZSqGhI1fnJl6r4B6Vek91mcaPr/T6+JpAwdk2ZU
wxh8ZvJMjXWBPKYIrw2qgJyWdxGy+DggBLMht07bbLXLnTpjXghaE1hyBJ/WrPV5mINQOgs4Kbpx
VCNrNEgl/dgChm89vMwvt8+ySi+NPHuyM7Eq9Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26384)
`protect data_block
iuBPnCK2w2fw6ji34MWrrOvaIZ2JDcikaNxpbMALEJIKD0V/zm+eQ3yRsrkVRp4p2MMQnAIADPRk
Pr8xYWYMcCgDDw24ccarFL3VLToKxxwNTlCGjgM2I8Sp3QHuWnacUdvHeYhHbX1rzAKcrzbsMyxw
T6zp21UOf50d/4Y8pLZv1p795DRigiBd3v+jIMWuBDznAcmR+VLGSdeTVKMdlPodwnam4Stx2Sk6
Ay2aEm/LjMQ6aUPRjjK8SXF2mkN3opa3qqT0Nda7WlLdEFD7R2D01IUkXlFGcaS7wqNPECAiK4Ox
MdUkagWp8BJaskkmk9d8L0OQpNMv4M4GVjXDHChT2zMZ3z4b5JDaxR0NaWNmubmvT5SZe0lVVz57
h/gwTvhj6LXqWa3+S9UdmC8WINcg1g4JddgGWi71Qk+jZmzxJnx6xZhnF8VKUwtbqG/Cg3B8J6p4
3aClS8jn4M+tp/N8suKllwHHKsBAx4g1UVfLEk4iAyLRS1uF2mPQf4JnJttyAMRgIH1nU2i5dEBW
9Uq9L+jq8s48KX4KWRSKJ8JrzJ1J+eb8ZUlW1qd17D2Kk6gAD44b7KxOg/zy6IFXXrvU2+gVjMOJ
M+5biVQspnCROPKmpAWPJchDk8zdf3zE7DcsTnoGgdrxVLAwExlaNMawI0k1/kdyD4R4HY7lhvnL
KooZw7DMvNjsV165vfvqQKs4gpvJoYkX8NlALOyoxgD9fdtdqg9K2F6oanca0Ns8JGsn2yV4wplM
e537dml7GLg0iqSbW1DV3fi7OCHdJSAQKEMv5cJ7ioi9gllTOKJWb7/ENCRbBWbAQ6fx60isoCtd
y//9LJIb4s9hQICifzC17xvP32zOgK45fySbzMcSb7B+LZV+0RSLsTx+T8t657TVafPaEs/D1w1d
bMvl8j/y8d43j/MyuxXqtF6hY3dKiJFr1v7d6tuq03IfKLJi2vEsbc9uuEkkjVnZyAVGfb0FNRGK
LxtuRV7lr2+CQ1dD8J+cdFVog2TR28e25EERDEY0VoDJAM8MTunpxBVHJVHyM7LLjwYwRHC9a9t1
LfcrodAaQUKX/6gedmDxk4bsHyppF8ih8pshu3goFC1xLAIOmWyzcPgdg/hrokjPiBhFvfaMSqP9
116hl8k/mbID33qbDOI1A90niGarcjNB0v5LNvZcWQ6+bvGgSTsXmvM/zKjx7M7oifXegqMPLJ2l
/BZqN+K3cpX02Ed1vUs1juAhCDejLVJ+RaLq0wOX75GCI0u2etyJw7sWbx3ZKqcfWucNvqwbTr9O
VXRaayZO8etYCAaZ2P6ZmEidNwx8Z6AHnFWz4zzia3Tzy2DZH1/C7uRYkx/ldacEzBUIxc6Bj8p9
9mW1Qs/bTXiBU3Rs4WSSwy3T7FLdGKp7hWL07pE1T8YVAeMu1g7c4feiY3YaTUzT2qaV2IdaPWB0
+Nj8syhqQsmMKWPhOjBQefmvAW+BALgFldE/6Xw77VQO2cALIPvDCkwrVTIjvsXJeEehpOMrmCby
k4viYfyJ4I3h84DkTsCaIGpzKKFr/zxn4UrNVH5Zh4hukuGqWJYr90s0aGsUw7bKnpAOMa/MXd++
9+9Oq4tGla7Pfi4ZjXO+NGBghFbmxkCN0JtLPu/MbSgiUlWFKL0ttpKiLnJRLFJWvmmfejlOZdrD
hRdrLd3AjpbSpQeelyll8LPfGKHez69EqAHEzZvln7uyTAeAHnXOCzpyFSj0aevynVLFalzmSCLL
9WMddkMBYa9A09VETz2YgXvrtLkFtego4XTEwKd8kjr9vfOEMMy/UqHLSekYpX2VAW+bqFpx56aB
WHID2Deu2AsuMd00ka2c0NDuCoglmfm/F6QsqKcFq1yv/XRkCKrkpaP1Nkyecp4/Q7OreZpN/xeL
lvZzTm5hSNWTLnR8wokczLYH+9KmQ1DoGa9nSUGfCEX6K+Qm05DSPPjPsnG46IMJ0NYqFZ9C6cYB
43cd7YY5pTfWynV/jLKs3pOIe9PZalcaKMY7Mxz9vG9vnMCoHnfiwUdgYdYe7yfDPuY7/FAyS2H6
BNhM2/N/BicUAPmE/4JNAdm5+ZMK1X6cfD3+p66Zg3YK0fd68H3oKc+rx6BNX1uq38SnL1stO3A/
8BdofD2mlxmKfI5n3gsAWDzeOLi+Izd0cpClWNVUhmIA+zu7UyDppl3faCgMTh4R2mDMXzglTlfA
2hEwiHZ+Pbp2gCiOQHoz2rMquGaAqq6Fkvf+EkPJMhDBqynn9N6buxJt3ONDsO7qwbwVeXKig9Lk
8xtJY03VA3x0n0rONexygL/P8HBg2mps5U9zPv9uQgvuhR3RKMWIiVkYRQGBUYvLl6WB9fSQ+tfK
AqLui0AwZhT+oADjKr/o27ADvt0wFaVZi+vZL3PjhvFiFCxj0eHcfTgkveUOFB6IqHQpHsbJx/J3
opYkfW6Jg3Sq11gxI62hirNCsIUdwJt2/NBiigZmM6XKmlfWwuvbGh7/YT+s+2inYV3N9C7rHiw8
HgIOFz8jwm+eH5csi8v+lP7bZqn45GXygrXjZ2SbC75Fmz6Ktf7qN39IxR9DzsxsYKFZPP3A/5m7
GazGUGRgi+OdE+W3K0gRo51G72ULfzytB89DmxaBX7me7c65XubmDBTmt5tPzNO+Grn78Cbivsu2
WMDtn94PMkQop9lRZhdNCPp8XROZCMlggvwQ+ZSze2tyfnh24GjR/VJpP36mKXRjiJ/QILCDhfyy
5JMfHz3Nc0sATI3wLY+JKjW6/Gbl/oD0ZHGBcMSZsVVARFM2jrP6GmGFfkiAJAfuDksr9T/SX3uS
3k+hNtamUbySmlNDGYEwL42K0GzdcVjuiEHTLviNvPBn+JuJdMuDaY67A2GW/3TVgxvHC93uLiLI
ldY3YouqYc1ZYh8U8XOehPJAfnBTyaNFbQS9VyObh2IiimCZXB3kw1H3P9rYs6w14q6ioNGVeEC4
klMm8LJ8cBCmhy6Dh0LrpEJnsYcVdEwRM3Baoo2XDYwTBex2wt/x1vMeTLlrrwlswkRyWcOdXDHt
pd9XHrFVfHHQNZ4UjYXtRpB7D+1algwpmp96cEoSbtIRn5XOfJZU7fDy4Pv2N48jjoZzfbZrVJvp
yhuq1Nx523PNP02Ub1++6c2Zo5x5mZiyn49O4B08cF53Wutx+5adJ/kq2e6NldapxW1kFyGQBV14
VS9VANYGee7qRfotb4eRMX3hs9HtY53DAy9OHymq3go+bZXfRCORFXjqejoJRc3AiaxENI/BYKL7
znvwY9LIhYSNCdqZ4vqDYkeHmsJgLjnu7kvxjetA8/P6BZyk5n/5j5NHtQv0OOuXQPMW6ZfbpwcD
7tXQzDtCOZ9oUXeX6mzOOClMQeszBqSsMJGYSVJ1wX5OTnuyHvqd29hrohx7UvBfn3lhyO5DRABk
P3KZ5CE1c3GwmtfD0GqET/M3In3F/4EcMuIATPIKifmUYAZso3uV21RKTAqXvs+H4WPgZiP8ntWM
nW5hcTcHVmgwppB26E9Cr2bspiht5iOj07+yYGRWzcaWD32X9qhocnJ0F6/BeIEeapaDZ+Lm87kh
hKkr4PkkmhYEzec/thx/TFlGb4VL+qz4l8zif9iXYEOMRu60fRcHxEqU/YaZ/TFAjdBK/5SS8EVU
PYRL7agQ7eK4XoR7L2ps8c+aPDlLrLhJCb6J3IQE4Hh3/GKMuuW+AoNLdgqbhFpBwvHU+iMacRRd
YNofyiALV4GqKAXOtZmfrqxYl+cm9FDjvcPeVa2ZeYKjuZ+4ff/ABUKTGoe8doHN+y58a4z7yTXW
wKLhqfWbAxj+2gm2lmayhkRZCO7z7MiE7uGBWqZGpR/jEJJd1qZZrQcZhKt9AoSE6fTKOddfJIIU
BBC9cbSM4ejSAkg+ioLrjpb8L/QLXYkSD5qqs4gFCpMPzCkpSr0lonOWt11NBgXGUiYFcDkRTN8a
It+Z6YzcSD/BpZ1mO3slhWuRam3IPy2wE+UmMXy+seYnWfUGa2LPBakIM6upWgKt5+m7cSamP/BD
DqmF0N5jaJW5oK7kOeX5Gzmbuxv9Ub0FC2k+IIfFSu3BDccRyc9ztba2C0DIOZ6DPERlZG4XXBUf
YbRWqBZnJu2UBX/616fv1CO2LLIPbtCr1hBHXF3uaW2dCdnHhNamT7FzqzmfxcovRSOWFfj3U8l+
6fyftY7lSUnyeMqWM02tGnNMGoOVS/rkBdBjFot9nH8wWmSa8AQ2equVO3ySRMgpdhf4ta84eAqY
0D0c0lEUnx2vVPkN/bkGbjO2o1nHSknsbnpPjJWLnV99nRhC0z9+admyKHXCWVmeHnUooX3AGoHE
IRpYO+5GVyiMf4RySaMS4qbXT9e4Lzg6VC80ahwyqOkeR6NcAdI3Wdqnf2q1zXsA6jjWjYjL73po
HrwiY7gQXBTiY1ub+JNVDvkSFQ8/q6he8T0BR4dfs/QoR1EO3pzv0g3jCdWBd2DrzzO/VrQbWqGv
WbnXp6h4cq/ti+UZZ4iBgDIGRSOI02U0fbqfD+nH3vGwmrNov08LxVxiOlqmphCCe3cTXguBr16S
M3qUF3fVL4D70dTxSFYoYLeAexKKq8TBzy+QT2YzdQvhP/2YjMXsLCUQm+6+0XHVNS6mebrBJwu0
Hz0EyRNVMCnOPQimA6ybiTN33uhN6qk3yxA35eHiJ+dVI0vyNigdebhUzyxOU051rG3CKrKE67ug
xw5yKyc2oygI4siM25BcIGiLJd+936SXGJ6SIbCUxRQBjlYa8XhnuOcMAinUbImKZcHVBcfTAnBq
SBKFZHv2gwFsC7l5khcLjwImozEfDDt5g05NnXFG7fUFSR7pzxjMh/qZwSQTzcp9GDpV1jypyw2M
+4YDCutdqzTI5p8aHuui7L5phubObMGCnypv0RhQ9rODucmQ/dq9t4752/3nj4qIoR3YJ1xyWyfq
Z7qfctITiJGpdoaHpij7o69gEGZwxTxsznWRAOOKCAijY7AP9ktyaSKXrgITCsdRhIog5lB8hDYL
3XOs0V6itRV9pDxYLbRao3SrO6yJwvO6EQ07cSuZvr5QBjqwWXx8nHoCfulYfHstWXgZC8FicMag
gQmGSXzzr/Rt/3Zy7tBkchfxYa4MxwpBid5zza8iDTRMRMER+QVXtqPz1Gf/wOFxctonnaMcqczM
TB6yHBRdbsoJwBzMKnhy9IPiC1WPu5bzNFXDlp+fp7G3Y8E7ftAYW+Oim+dsyhWBoQdLOTIEaMzb
08Vl8/nNvQmQ99OdHTIkHvpW1JyX4XHy+O33B6YNqpW2Oa0Ya3UovjqMLeRgbsn9xbFUXautalqb
NFQOk4QCiJX+SoGOUBmeYGxZu9D1zSZTCsyDd6NjIzRvRK2au4qnHEJ/mcQC/mFUzGmS7vL05k/M
s5JLuLpIxe6hyPueZsSrHilwS0mM3TUtaqQZqAbpa/qrs448c7G9zKWShv2UgIWspLTyVeRCbgeR
zeHGra8dIbB0nDUl0FsDL3z34uqTu0CmprIeNftITebAnrsSFIBpgCtfz5T2ef/e0FJ5qGGssuXu
cz//i7e9beCmPFwMgTC2A5CzI4p5edYKf3FgwQvuhjyXw2AWsk175EsHfr05rrAGF2EDpSDDENaf
emgo1VKxoEFXgL/BQJ1rgYUkIFtbSS+sTYKum17aRQiIV/H9m8T5wAXk4mCl9OgijdZ1vvvTd4Na
sWdFD80/BYejsl5pG70DSI/O+/N/Et9LrY2k68HAfEK8CVxMYqDeyEdek1RMQG9aGuJkQciNLf76
2coQIRd4SVN3nAjLCJGJc/CW2hjkCJ+BaBGnjjNaxLS9EaTsSCcilCc1z+BLChdW63txFdFY2qmY
m9+WkzfEihoaBr0oTfh6xNTCH89QNXi8ZYb9iI1ozpBDIiCvLm5vZp8dhRc+yNBsSFEUA+ZFhXMG
BaMpNB3f5FEx6VXuec1eaevZUa9DZsHizABgD5/KtupPE7KSKy1z6h9YgS67SzyqKudnpdYUOs6d
zWWy++nEQEiGF52aWbtgRiDBiWvsq9tOFpkfcP2zWO5MI8EweV33mtLbDsnxoNfVez54u0luP0me
k6UAw18uAuE0fy+pW8aHBN/e5kuXDoTj4k0VPWDpsSLfF8Gu3bsbXX5ATBFI4VXKQI7A1/XqpIB9
8q5fmsLyZjzu+bE7xwiHItGTKxU+XRNlMy+gtJPoiiOnUY1xu/h7GP0nzvqHyKf0aV0GtC16+hat
2Ho1eT0ajyeXWgF9HvRlzotpmCP4IPAd5QQ6jcrRKHC3YWHCXxtxRquPgsQeWPHb39jDDLh4UMLg
3qgzjPQnK4SA7dNSAg6gjxODfDvGAXAoCDe+U5UGf59tc8+gq1TNPnabdpGxFnVXXOXNL8IUvCWU
bCmYPzPxzj9gR2ha3q7et4/xQoNH5Sn8kcHRg1g1GnNoXyHCKS38X5dSJcykapYFmuSWFvpmzaYX
TXMOTjwLWYhv9hO+HczIKPzMiXN/mvy2jAp0QEH7cCUO7QuBQ/eu1zDdQCx4ckSnrOwwV4hA/J27
+PD5+c8+wyW+OL+dwWNok2haarhhLqpy3JPtWXpepg+sV9R+asc9D3fVCG7U2qHs92bvy9ouunDE
Ru4LfsfgSo2pEAd3c81lCB/POpBO6eXVkSz76miKjB4GVgC2Oe+pyoLvtQd7oTApT+4+v+nPm9KW
SmJsuAG5F6D2XZQ87xMa4iqo7lIIcm6XgKIt5QGu1mmVFqd6OcJjhBg3dXG7Q+HYF1UoYCvIDrw+
YCLK3L43MEul1SUU/KvCB7PRHEVmSIXw7q78CG2xCMM5e8eSHxybEOMI5grN4uIc6hh3saLLQSyX
buV0zbC1yaH4iQCU+VqRrqXHLpEtd8mgkXNvGgH9NOF3nqixmarRExrCopp75hQcpt+X1X25PQ+n
ZW+8/vXVsg+uUIFlCEeieSyTu2cn5vXeurqeLj+yHp7TTnOEx5VGwNGMt72v0NuwKQqRUi+SBIkq
BW/HTOzC+aonYzypF4GpV78t+py4ukWx2kBDxnKW5XeMYWYL7yVHfk2PhdH1t/hIEzXvf4N+ILbp
g3wChY/KhClYIdUkUVZQXpKkr5m3TL/0/EzaYJEXmukuhoeD/SSJ2U0zVi6/24mfTbQk/Yr9plQr
aiBaNppAO/VMkXEDZ/afavk8zyiE482uScxCSZ22u0+TcNKknQtF59wfexPmi1f5Dx4Lf4IJskmX
3exg7ulQWj41D08M449zFHaStlB1X1+KadDifsLvAQXVc3HwZwgw7Ody/FsUZS/9yjxoOGrUYWSI
ZkjlT7FIWwQjvio89gdZ+8LIfDG0g0HyLuP/LamN1awAFRJfMlr63RK4oy8oFpyoHuS+QJ3MuMGC
aI/YgfDHZ7TJqki84JDMtJ6b//ep97mXG57SvR9BrvqcWlTql0LYq7TUQkSfzEl8qMYdfK8dJzdM
EO9d3jwlIbtuYd2G6SxCfq7R7sOuEEfDZ3w4OiN/RRcXxAxLayo2VGjvT7QVJE8O70JwpANCFxIF
j/jHfUTip+YTw/FfJXAN3GLrp6QRUl3KJyAJQeW3ke2x2pQ1hAyIiuCxfQCX5uAeFGsDQvgUPT7T
rjzRYEhxbAH0/juzpTdSaW3998f1UoiSIlfKQ8xcwDnFL8hqAQCiB4EadfCCdFO3TVfN5dDmVn2L
1+pzskvmdh1zG538BN86U4KaKHU4Cj0RZBYIOVokWw2AUlui2xsZ6LP67B4n2HCU8OAqHpgJwxMT
cq2L6UTXexPFev8HaKQ+8h9jDINIHTJv9KiwV0NSVi/lPFSx5Xx7K9ViVd0sfXANvPAjloYRhHz6
w8zz89Q3SL7LMGboH+bPtYGYse36IYM2T5o2OpTSD+AnWa+dbxtZPfoYoEevc/VgwqRJ6jvkUvZj
RDNp4uH3vVgriWZdYWNkd95MpthZwUlYVgZBe01JJYSDBp+aAOkmvimLkePaLeYtkaKs0i2FoyAD
Rr2mFkMPNbeFyifjOfG0aoQNAPNS24Nh3WcI8IuedLpTj3Fupb/YAPxu0fhlPKNUikImwBpJHR2W
LojSWStOlwDp/9u1f0nocsjiTG9jyBjK/vcNINFwl0cgZbNKg/ysnX6Htv50aKLI5KcfZn1NBuQz
n1kKhUP7nH4lozfTCPrXts+/mwEbGMzQtevwgndEFzdYgBh30GF7B+q0LxIb+Uglk3fA6TBrYnfh
/T9Lg1mdllHivKqXvxhgisKOXbBonLs3OocDIpXsEE4hGXx131J5c95mO0HNPHWDqKMCAe7ahzEe
tfZDq9zcqV5pzpV/TMn4VsoOwZCX4AXPacJuMX79zBsfcXSPz6wgeIGqad1I2Mvp+fMzWZzVIbMN
q27qmJcYc7CggozVTZCx89DhMJP7QdmGNP0h/W1NCo29PdfuBnfoIuyjc6y120VwpsNLnIUTdAHD
YTQNSqgVon94LircZX1nrqJLT+0CokJcLkT/IKGX/3aYUND2X3REt3RrghXb8NRF4zL88cVjlfQb
d9J4qlCxKWQBGfLx7OjuHNw5DH9mYiBUus3mPimCFT1MnwOBURYakAJRNGrkVrBuiePNzdlbWLWk
J74yyKEpNKeaiHLU9+oCT5/HWkIFx0IJrKHT2XkzxeOVcyFP0y3fSkitHjiEcb9DCkF1NSWAJD4x
FmhUhsLEuk04nBJxDvdaYqxTjDY9sV5cEZ02xCBdYADOvz96uF+5mSHraUG/znVh2FcoNHkIq9h+
OAdlxi3rcohqOGKPhzqQFeVJYDQJKHqjWhYvp6iJzr+it76cjaDWrjjeJQ0ArgYMpnoTMlkfm8cv
YamUYd2V29pXGan+hHCkbyiuviU28MMK7SKhLL+/2TxHZmAIXVkC7Eu7wVhAtNrKnEvrtsxvNAG/
aq4A0BHdizCmkBrUQ5REogqGAmonMgddxQhecJMKWiqi43lcyu1K42KyCuLEerDobbBERA84z8Iv
2mzwc/AEwXQaYKnDOtK6N9G2atfdqDHfWkPM7mWMQaJxp/IdagctMm+l8Q8Xs5sUWeMteuBBy5p+
Q1ovRRZ6aYgK3gu4wWaXq0Z4UO+I6AUstucrBy8e0brOKz8zz821VHGc9zMsjp42sTIckEbDXZg2
nxo6iu9W1d7Go/kfjAbZ7Z/zr9AhPtoupqEYsL641n1wd+CyHeWz3bQTOmYfdviWEiSOFzNVybEd
eCmJBBadTRHSMjy0GClUKxnZHzOJ8QeQCSgsiEMO61DcDwp2EcIEdWcT/c0MDg5eyXT5aj8FLk2W
ZImtMCcQMvaTOMhVB7KfIFcLFXyOyVpTHFfJHKFkyCQcuq4ryvtbcZIf/GGdgdLkryk8yPlnVhfj
bpRFbHX/LX3tbIosErsnUy1bbhx+F+WPTAZZeAW7HB+FbtB1TMPuOnfXT96BHe9LcGHQa96xszf0
J6QEnYuLABDwuxKgAamZ8ldol4jxFmzc8aM5j3h66cUR36z0gsOl3SCPuvJ8IsCstDbZzU9EWSYv
P0E435EPEwS9yI4sxYjsqFAWLGwAMNp735B8P87mTgPSrylsJLRqfzVrbXZzoGcgcZomiP7AGuXt
I84CLxrqkYzUvAIM3TCyGAB5+3R/0GegzUkSiavo01H4ivjgKBtABf1Md8B43+ogLSs7W3fm258H
w0uMEl0dfC4pBqMqf4gluscOxsB/OpyNIwv7ru3v1/osrs5ppImYra80vBY1u9jzIDxn6vrLevvI
lp5fdgTBWraPWyI+DO545c6eSBeowOfTaEjm3Ok3qwsEk32NpNhl/rohZzlK2Vnq0JESOFPlbqdg
zKmYDpw7dxvxe19hTtbeLZauOHaTd+QXdS/vG/quxlk2Y46qSxIlBSFSU+Ls4yMeLcnHDy1l51KG
q5KY+IS2X+AZftvY10nEGKj7N7A0sGA2Wp0R0i8Ef6QrGXZcgf/SihPPVQrzIg+yycWkPiiBn17C
Fr9Ks7RMrHiGzzzcxcKAxl/LGE6/fG0KYvl1aTih+ONnWsTFYitElfHkecwfSimL2QIA+SDCf3u6
ntbqL2o6QReeL+AJ51S7ifpTOYD9O+o4gJiBzZk0MX8i/pb3bPgyuLyaNQHJtCIQrnsScapM82vI
A0Fejq4j9nJBCvIlFzcGJE1vO0edS0/yxEjFONhGQIub4kKRRYKwLqIPmJ5LxhTP+jYDPll2Bf3s
Q4onHxKVL107mB95lLCYK5NIpdDwQBh9d4hJBNzFJVTdQXpQIJmSskAHu+72Ug/3J2RZs75IrgmW
pTp0SNuPJym8GxPN/cQkEki4RFILgRoWQe3LVhO1f2mpWC0NCwZ5clFL0UfGJOEGreLAPyMjMqJL
bgdrtqC88sSlhLgF41p7GgEfHI+7E3LYQuIh3sNhEsZ3+iu262wMDdiV9H+pJYWwjrlS/Bc9q0Jo
RkbXIBaCgilwAfI30bGeEeOuC0qm6YDeO8DdBk/TcKBg6cmWd8NQtKmf++Ledi3FrOquWlQA+gU3
xoR3WTIlUZniVNKgvRcMrDUwUGq5WCiMLEd7I+H8Dp9DpOffOmEXAbcdCPxo0/8VcSKCru7PfHCn
jNshAHo35LHhfjhh9zhfaiv1GCyeXN2ihtQ0wr4cWNqaBn9pCqfG/doy+9edBYRVJAGkUFTbXpTc
gd5TrI0gWiS/U5Kk+yEjBdRlGgRY9kk/r1tPXTDChFUG4QMq31Dv84E4VdKPYE42iIB6e+1N3o4t
SgC4qX3ebmJ5t2liedlhvmqskiBLW69k6HZ2AMFlwyq9XzxyNi5nW57hKYUgMyY/8I+EjOcjMQjb
xL47mMmTwt7KUngtrBoLsvcEtEMIZ+EqPKoofpKpKDbqSVT08AI5ifeHdYHvHNyfNDGb7jo0rDcZ
SuFMVYM8LuT7F64/67llGawdTO0DMXNzzTSIkq6PUddHOpZQ5Ok7Lm4JPA2Si1YpgONJ01J5ZSUw
fjO8dRcFxwZS7tSKAvT53aVSybsHDRLsSZDih1Qs0RHNR/F8KlUSP2xz+DSKcai7QhEUI8XYckyi
x5Vyimt0OqsttLifMfRRguGik4whsscpQe3sf2/1PaDd87ev+opB18SNTei1MX27zK/A/h60wlep
tmKeVs33H4UZnie18l5Xdx5jKWpacn496OIP3XJsMHys140ZowcSWKriAh+zPdgHU4mUq84AlWzc
Atr+tMcy+XzVLC9xMsGwqBa5UUOIyPW3hrgYiHFjKEe02si5KDzfbVdLmexctTyxxt6xy0FDyRaI
KgiyrB0x4m8hOUDkJN2wYSYqO2LcLsxbV93qLrCKwWnes8XCY5d/mJTT7GlyuNYEj0UzePVjigO/
FMAl2oA+64ejrkfNqZqLBbvEmA8QXsAFgWyraLjKNabW3jk0mc4WH0fKvaUtbMmq3+vGUKZYrBwQ
9USUfCtwK0FYqUa4QHpM316TdgHT6E+lyHgXWQX1KkCwukwnTgrIFSAs6kEsictFRgkjagEE7k2M
fDcMOcSOHl1qRiV49wpO/czfjlm6chX570JvJbsiLqSMnkrkMKIT9/zTvUUdslg54ZZZrUXLemUI
d3eyaBnNudmN6SytxKgEwnjJZTcjFgS1TQdD0keYAfoIImbEHv+IYSjNXf75BLBKUw++wdLDR6eb
ElW3Krlm2RTNYJTcNS+nQAr6sTZWl6iEoihrG6fRqE2JmrdphiJNLZbIel7iYxTe8kN4nf/n1G3r
XpNcxzzftz5i1EhhGDl4pKwOGKJUdHo5qEjlFQDdnj/hgNflmt8mH+9GCNVlS23eofFzFPhx+Zdg
UNMQE0AzvipSZ02uaO2ekbXfzbNbCCiu+hOn0BM/MZjCO5KELAXl8sxVbeTImMBfDvrEOlvRicPN
Z+tVJLVyCpz9eyrgNYYYroCAcSwT9oMweNtxVBcUXtjM+nNTw/+YYgQ0tFrYK1hsYrNW7ZJIwOrE
Cs0/TFRQOBhN94oAUDu+oKpw2thSyby4V9lKIw2ZGQF3opKAbmevDV3tLF1DUfl+DQ3mFX7Pd3te
P9MqPn45WcvN8BBlNE3MGYEgsSnfl7Up9TT5nFTYPJHI9FtvPV/c+uDc9LtXJSkKtwVRyBsLBiQh
iMjKGU/+PfIbPCnEwLPVP8cTKK1/HPfmkUF6EzL9kmsZfJ9ok1f+EjdwYjhqIbwrcTRI2Tz9MxWy
WRkBwaQAVQV+6T8Fj0OC34V4JykRA4Eg6J5qWrJlT6J1Xzb/YJ02BkgN4lkFl5IT9xlo0o9kAVNV
jwZ6v5AMheG/PRh+PoOOjW4B7OFKrXRdNuAAYBBfik+oe28IwY8THZoZpypQ7/2G+pDjBzDo7rXW
SPyhyW71l2o67m1qAxRAssEDqtZIgFkwfhw2eWJCi/uaL/r0nCznDy86f34w0zI0vG0/1HsXtR6m
oEVit0Pl73Vt3/DKIdCTELi/OfmHDm+NDqnQuxDdVr7Zm9wrf52nPvcO+STbXcS2ovcqRSAspsOL
GqXyDpEBmGZx0IJToaoUogRssky1GhTWG7rkDZEVMAn+xNPA6SuqtoHHQQGrfsUEQXrFUpIjXw7n
dY3eNdkrhZsUBIIQgp5c5nGzM41RoZowrkcirVCsN544CJd6R2ny/s+2fyIo5QcNj0LH7JAyxAKX
xfGxf5QeIJ1jEI+XeoWp33r9GxzkpxGQqxVyIOcT1/FhGsn/zUFCBpv3gO5sk2s1FFnvma0wV7Bh
3oIAP79TbCMaxzrmC5X5Zgk9mbd1SFErNeAQMrZDyZ8otGDDLBibieudpZ27vVHhP85wSV1ZbTTA
84JOJlwxVixxb4mXjVXIWr3gXYoBDGhiuVRvAN8S76OwcOViFeNZXINBHHDwaQzBRtUWGjdW1g5Q
xnwNks/yKMbLnbZ0h6C/YKYXjvurIVxntQLILJPKKOW1ekOZn2yz8iGf+nWnpGddXymwvfz5KVDa
Eig6FvI9NfueEUwov8Wi+9qqLnxiIthjrQD78MoDkeIrk0igVMoT7jnYHqKc75/aoVf56gcHpHEH
O2BoVO+jnCymiBd2T8TP4okKIPDBpLENjlL46fDkbY2bpEyZuAIX81TVz7Gy9FQTQPhdjyqvfhi1
IC5PUDc5Pm8RYrvIq2taJYzDnbKUqSqwwh/AKjOX+MR7F61WIJ9BCwP2AMdHoAPx2KUbXTp30jTs
R4CK9hSj97CzN4ov7z0E2QYvlQoKRCNttntXeKXHaeXIcOzVktoOUxMZ+qjnC/NoIwhAeeWVLzbz
9Ld94Iiib5131qeJPHIImEQFK6VNy248noTfPj91TQ/LdCs4+S1fnhrzF+I/7ahmDXksK3LgKQ/l
zgNHD/gQWs/yAIcwpLbe34ECEQEhVYytlBDh0cc2v7lOZjlP01hw/XH9h0sVWYZtvgzYJGjY830B
pXw1xtDaAL1xNAvnten89ph0Bv9lgoLUzXqyHsMwOMCB9HIxNbDNEtCdyp98q8a7fVpzCzYwAkGw
J+7WIgPO6cg2/i8jlYB1b6rqqlzgTnucQEamobCo6tkz3UMBa7BWbDDQeCKqwfdXzttORqq42aQd
EHfQQUCT85/OLHrFNz/7Ftt4pqaLv7A7if8VGNEoSnROBrH/4xM73hQPf7pFEIqGzGMjqmkBLdxO
0FC2Xm3MK+GHWW5UzDntb5bqRGgQkeMVvx8FayMOHcLwabdLEeTG6IjNFG/q9adKKzHphNrnM0JP
3Z0HY1rdGlOQSvgLxSb2noSG11HdYnwsUgdR+46VGnWJ+srbZExIg1flxy6L0feZlkWvvz6euQWL
QSCRCnZTL2S8JUo4n8he2n6JvcPdVIzUfE+psX2xW808wIj/oZsDJ8ntYdkXfGC+vVnBBQBOJKrc
V+VA05tZApq3dCarmRFJKqGpIJpbR4HBLHtU1PzJwWdnKO3nzqwUvumbeQbMGkDruDA+qYGHSrXS
NqzdtQLlTFWBg6dlrAVStzOOKCDDdke3yaiDyrL2x4SMJTLsYyttFUCle59HZWVsRtdM/eOnzN9g
xV79e6U3pwXzXgt1/qoRISOoWjbIR1UhfRK4zl5u4Y4ZccyIenZyh1wOK5n6lYE3/74AqcNb49zI
6zr0baCYicGP+ipw+X98hR+xpUmlCEdUznKhsauY3b5Ss2eE6pSP3i2jB4SxLkQ694WFX9846013
ASrjJ3cmS/nalXBwiIqz2iB0J0Gpe1xuvrgQQJ1dDNcEi1wnDZBnRaojqv6+yXBretpKH2Z9n5zb
xJxhsRlMYi07IhpPQCZo0bZaDCTGQroT3dP1BnC9hBV3+C9eFkNlYopUKgl56ajSt4Lx+8EUbPsH
bTg3aPOZjNZjQ6950izRj07UrnwHePDXa4oaY3a3qHNsNHk8Sj292Op7xT3+JEOWuu7Y/Bv/qByT
cfX8Ez+gCFf9Pd/rGHjRTCiOASPr3qFy3vg4f6ojsLxgyHDMt6y28T+cAnYPmAdkXtzU5bVYXROW
+QBNGtAKhXC6S2wRTTgt0/gLOJsjgQfQicj/G1jkbjMeuK+ZfVljuGuXQXY07SKUWk6a/ezebIyK
2aiG+U4YQaI2L+9n4gw1+H0CB2xBkbkAVk4hzWNXAS9kJHVEottwC3cYy4p83IYPtk+0x9QozGaq
ibFwIQqUHI54tihXyZ6qwYllLzSjH1CYDwHVtIaFfwodwESf8PEfrqZJRNfZgRKBruFY2EJ3h43X
4ylb/ipjC1lSGyFxBSs97HtBlSxSyLkcRsQKYpGr2nbUjPEJufnU1nD4oHOyzomDaLzYYO+t8Hv4
TsGaudrx+Byvnn3LpGb5K4SxRIBm8t/uboTCahlVAXFPRRFcWtwj0YmdTrMW9xlfrZuCCCpgxyrK
Ybivj7miOr1rNmUqHls5t1PZ+3ZXsYv8HwqMyCPk+Ur2P/7ggWWryc9eUChD+pA68Df47V4lU1nc
OAqjT9lr0HmbuTO2DVb2KsMw/859/HTvqnCJ49wv3PfQdm2/xcmdWxWBYpMfeFki7mflZMrC80Cv
JUZdVmxtcrVOZM/BD2CuRWtq0sSQHH2REfgCDWMOQY2KWrJzNdmnUHzNiQrZehhlgIPjNp8TdCIk
c9pwl8wLM5ziT0KWXWDbrTwzJiVSg5j3a+de9KdAVMab7WM9X5U+OFSiWg+VkFh4irwlnbKoP81S
mrxM2yuzBmHofLIpgu3DItWiSmn3tVmy0KIRXUSqwQCtv684m/QNoy082G+Lb6uN6xnXrTlRnU9n
NJWmJkmehpAzzkknaUUizGzcDDvozAulvgznAjlK60CiZVy0VUlmzEBQPv7qPxKgx96hRm1O9wc4
PFomvLm5n0t767Ke4kzm6XotFrfZsiQbCp6sjkWehGaTZio5jOZagTvOshqQPwhdK3s8gvNqn1/z
YerB4oSNWuqZP2hntjRjZAhNfhilGQK8f/YF7QwbH+LzC+2TBsppbq04PzIujtGyqP9oBzHi8zkd
SVaBPtSt6uNQcGzRXFchN2kGozlkp0dnA3/hls+6M6akXPpBAWQs6vDN6gJ+MsRCpTsQHrOo7oQt
+ZKyIXZWosA8o8ZlSdWzs3wh0/X+Jvoq7IU3e1ED/kaoCqKTUeXyWqV4GV9R0JAkTylcF/XfVUbo
WVwPHjXOMmJK9cslwd1vI6aoUk3wkiQ/8uxus4Tf9mekXTrcUZxcXAvrpzf5pMpbVNzNzc/X8N8r
VVqt9ZGRk2ZBe7Vt5JN7H76xV2TDznD0OIWkBN6/UKfvyOQZ4Hoxc6Zs3/ACGR5RYOB0SGXWY8Gy
A+hO7scLsQCue77fqojHIBs6ZU8Y73Tz+dIkMARzPG3LyxFyHpX5BPbhXP8IFZBiO+qgRbV8wXRr
S1GJA8dkt7QujS9GBg4tFucyYCgDfNJpeSJHiN3Jh66oeU1CihRIAKBE4yfGQYrLyFbmIJaZoDx+
uKs+1JPC5SzFQ97NHPth3DS+Ea6tHLYmEnsrcs501RSGpV1t+8FrelMwBTVa+JiP39qw3hPY0Fou
ygUuG4VfMCzAcJMcOOvU3WNrnd4cDPwZFex9J28Z6Rl0ldc8eem5Swg2OOuje/1U8krMwARwTeiH
vvSdbGIJ5UixbsWowZ0IWwTcjYjBuJXQEYzpnM73MTOnMrBI7MzWhEEd/OCtODm9/IgjimVz2A4y
y0W/7PESRWrnDkD0P/lnwQ/Gnfaube0uLjI8x1ZRERBRuy9Z6I7yVdPHPmuaAJflSl/tvOElFO5c
u6B1AVsjn2ZXqtKJxK3+iLf7oLMQnYPCfsDbPbHbn15U0ODbY4iBQblau9c1duwplFrwgXD93BY/
1pUgOi+SuKvCuMNiegbN4VUw/a5iifA4eAldKNvl1vFj25ZRlSdt4fC3y5atwzeivMP7z2CLrQet
MK4xX9k0Zj/yHL0O1B0E6ldfcwBNhSSm2RFlQ9m20EAHhTtKuXrsx3TnSEzkR+CJv8vshz5tz7g+
c6U54z8IyuM8t5gAMcnRWco7o4ICXWW9R15i2MvWZwpnnDLuHR39I/wHUrVLcDXBouzcqmy9IBVm
PV/QOja95eR2W/4Tvvt0tcZvg46AH+0fkNtHrLvZ3gD4oF72Sm2i4pjulhdxcUqX7IkybwgI6P4T
U63sUOd9asq23gamSukwATh4+808onSKp93RflJSKQmCJwi8qYm3dC6g9jryp4l0ZLIvGMphJ8PH
i5BEaLpsVCA5r6RZUeophgUOsqtbdwe5QMu87RlVm2RrWcK/fNiZXe4BPmp01hNvb1TZKow0tJfn
JZNqMsuMleS4FjCKWFtJGvrASJqtBn2pw6vckwewqrMMkEEqtMtnJ11ye4qEUpaw0mXsLn3kYUpm
qO0KdjtTLEw0CtNe1IIzPeL5AB4o1Tbt8H9Ye+EDdGNChrqZUSjLG40+m3D9uh8AWPjsUXrJrkM0
chLFOKBsi0cLoJGHF3F1O3CGkW3gTbVx4WLUJtR6D+PSgYNN7UP6f+OTMwg/IOcF8foLNqPbmnm4
j+kMs1O/9qGTMSgAR6cj6swqbzk4fndEbK6xzW24AaEaocVM4XIIhLXu/Pvrl93gXhI0smTyIYAS
66RP6WABLfVcsxrYhyCKXQSQxg4aaon+96hbn+lg3ByIa5c8DecElkd1Hz+4SuptyelrMGOfNn/Y
J/jB8uyLIvUvH8vXAFCaqzAf39v5K62oIfobY1TqK8ohqvsg8afJeZ0u87NCpxVSEahFvm5unOw1
0/1sIfRupVXwBlJ5U8oTNgdBwjx4uVMQJBPDPhytfq3Cj3OWg9Du4ibiSm0bQ3I18tM1rwiY/WJ3
wZ+uc45nkmUyetJu1tN/LnqQP/LBb2x75KxAhI50SVaqXbMqUCwJjY4WQWDpjatoL+qWFn7bGP+7
gO+0Aod+pxplxJ5Y0L3OOabgDHrWJvzNZW7xU2i01DIpDlS8PJOsvL8L0YPUee9q4rLeDLVQqC6h
9SYGFVitSYI8VjUEv6eA2tC2kzi9YUDXJG5AIfFD0cKa7Mup4lwH2tFDQqjd5yreEDc0rkfi0VA5
41WXYwptoP/8tKXwlGtaMQFUc724MQjd1XIzKi75xAsTLJpCllzW8z6NoF+kUZ9nQ/N2KI8a6ehy
Jhy2tM7heuo+6O/OyF1E6Qm56GS3jrn4QyIz+B4/7ykeS5qQizzKlRYoH3H5lyJ8v86y/rXhZX+w
8fipm63XJ1G+KPq1ZAJL2XKL7LVq/Di2XYOu8osLPCv5tQiIQ+7R3SNHOaS2OazuGDTuujONaoR0
iR6rydG1WdToCv8QsPKlxggpOUmk381FrID+K5+ut0rskKoJ9lNUItcA5+7eYvwOL9z3lnWClH0I
xNBn5bo5TbtReh8pFszyyjnQ2dwaCat776s8tslN/0hYBKNTTIQTbYclXZkhni4ewoQoTdp2yYHP
H3M5eyEVDolH4AT80b82N0thckvUKV0N+H7OOSQk2wTLsR/k4PBPUzr9o/WXj0qfd3nF2yV3aWjf
7HppxnWj317PFAl/M9+jPvSywwPhKncU88Fo8ApllZGP5T0UWIs3VsAfqCdFxAhnVmNx4wcxMVCL
c4qFdN2wney4tuswFd5rA/9SecCKBugrJvYmPJrFO8RE0VvBxcxdWyWQFKuQ2QIOsLbQduQVXIlL
7KIf6q2jUn0iHalHf3eb24deg7oiYjb7KPNwj+jIKTEmmH/d52OiJgL6/sAHitoyZ3w1dsa3AzJu
XX08vB3TDZOD6FrnWrhY4C+InfclIBmnda1/U9eLwfijjgqaX/wexwlaeLL0vrPMyNTfF6Z9DDoP
S19ydMc1XobKn7ub4mc3S6fAOeog/xsHDsfsOhn+hxn3WId/K8pt3N34YHVQqW622TpQxdJPI3ft
B+T9QOEYoj0ToPTSC62A74DDRqcSmfdFP0LxAUDy9Yooa407F+BO142UC4evT7TpLUprPohEp32s
wUstOCXnr/XkaZBP/qyQpsXIpd+52cj4Wk/tfpDMJ13FW+m4qWXj3OWCzdA8NkpdkjYQI8H3A1dF
Mwi6xRB6JhqguUuppf1FUGH79d8pxyPIPrJP2DrVVzGClte5AYuOBTfqXCh9WqWfk3qEHbNA+D6U
N7RtUnQJCRyqGzOq21bHCRUC/fHt8tHsG4KVvne4OZkIGwADQ9dQ0C8/YybF6TocKwv2sRoWs8p6
TGMjf5rW1MwHDgKyJ98R2hwNh2S3yhDyml1k60odN9Pqj+s5LcdR6JnNRjZOwpNamWfKxXHuW1pu
+goUKTRdgVvh/CO88WLGf2cjrKgdD5LdDemB1mDLuGUYA6jIJRubR3aMjE1X+gnOgeuHOHLl1MGT
jG7szd6pv15u6JhaXxTaFE7/UtT3G2+EefKDJ5Z6PHFP6DmVx/NJTeSrymQLhPN5vk30JU2d2PwB
103iEGmiy5tUBq8Wop71TZARUk/GJuNAalFSNh7mu7uVYudJ93YzIlfB/DVXpbsuk3OtrXp4s33d
HQq0JVo1Ym/gkzecNHp6BL9nMwMv7zMBqirGzaK5g4AING1YutPspDOgWekBtrIuZ8qYnndL9WyB
v0HKhgXbahUol9Zk3obHI5CtqW6T8jklkHip/C87Gpt3gnUCI7dKSHfXkM6DVAf5R7GS5agte2SJ
oQETT/3gOnbfgTIV0ZUOTZmvIrBUvu6zTD/OODADDs9uTrUQ73jVrdaw+umGSuHyYvPCZjoKljzr
ESC68yWZcolgw20e1NiZRJyeRmrnk3TYgCQW6Cn0CFrAdeFh7w8//mnmI1ZTyVmJ1jS21akwwGg5
LN5o80/+IycDrFux6OsB4SDnv2MKwsjFK0uFwOs48jAxvZkgKqrro7oKqBg7MiHEVRmhKy8vug/a
+oC80B8MANV9F+AdMOAaHQ9X3yonzbmCye+KC0V3FeMY8qOg5JDZ8nlZTtCRfWRMvhb/JBCInL+z
YEf/vv3QceD/A1CQAne3dM8epG1yhFdxG0yq053sPUuI1qqBOojbB8Qv0hIWzegB0IDi195BHkpY
6EOxI8WR59/T48uThZ+Ewpo0jpi9ChkaPlkTySAjY5tLiuxTsW2AxxpgMVsW2AJn34W3gmbfJo4r
pikJnxQsBflofN3J/GgKTWbDPc3WGd2oZDjVkjgl8M7xMCpOp/YND1QNc8FaUICNaumu7yiNPMJR
Ylc1CkmrHUnU9itAyjD9snIRXGvIG3+pFdqSUXo8Nkkc6Wz8yJMcLJukqXcPGnRJy3cUf/0womlg
W4Rtef6ux1tcePW0gymlX2XEnIIvZXc+UMzUuTeu4wdcnGsFVB29KTa6c9xaCWG4fgaYDSG0BMsz
0g8Sxzl7Sw9J6LE8goHx5PNTTARz1lj49eB5lQnDzCOHMVz4oJdx6h7I1vVSeuMWtXMtGD2X054P
bxSspyDucMJr4n3uCOZ+HUyHqvnHupVC1k2DAJTPi2eFOOUuACiJrR8333feEKOAXPwyDX3hTEBJ
CkG7gIuqhNsRsNijbRYJxQLdrPFyOhf2ZgOeTqLc9ZIaKjWl6HU9XfrSek2JIFqye3ZLifQtjCSq
TiDUtt6xtZIguHWRKEdPIqgvin8LtrnUY9cOUPfQqQU1u92v/XBoZuquH/BzGVALka3FOyWUDvyX
tv9O73ihyZwXTMnIXNkEI1/SfuW4/YAlJCKCGF2F4d2dEQ/RGTqZ7WY3CGj7p6MPpGfaRytBS4iE
e9ou8jYx4fxMextXtiEfnZajCY90QiKlANtlhm8b5CmFe8LyS4HsRPuNRPWgXkqjV8I0OX6uXiBw
Ng1scA9YWP7JlkSfdmkVaMwhtVtTYG1pP9i1aLSmpzHIq6lQo4sAENMSbS4npJkCMGEiGrHGYRi7
BigOCITGpOa573aALm5gyzHjL9aej1M6TQkfPzrH/8+CTYMi27RiMXV5LNN8jJD/JWAU30pSpaMG
9/L56tCtobbXeI+I08zadwd6luGFytZm92Z9U64KXwrOnQrtpPOaCvmNIb5lKL7nBWMDq8g3+Y20
cZ+26VJEDwq0srj7GLI1wk13mdJQXv2hbX+mab+rhifWzgHyiBfqBa9SlDuH2MIn0N8IYFNxHPby
2owFB6sAWmx6BnQXNmZjM8ukbMRjG7zAdgTSc5mTlz0L5oZaiqueWEc4cvBiJoRJQohkv/GruV0u
/3IOoIy1aFiQqrDUWUtao6fT8rdDEXLuZaiafY2ymjB74Tfu28WxaFL20U/tr9yiqu7LxImwWTyt
K8umM2q8Arigku1dl/HOV/5a/8YBZa/bc7g7NajsPSaKcE2XqT7SDm6WWqZN8pYUp6C/5EezZjc2
Od8VgfIxaUiKuNjGvg2viX31G7gnCRxe9lKLiJf43p9JfrYx03W6DaIUc04/zF2GPbczJtPMVVsD
bBXnBojN7IX1/jfXYMw9n2PQrcJGATNjRYgTGGoByCeUllaBl3CjYyqsG9EvXNVD7PRr12TQ+RjM
0HuxuPTCf1luw3SlYOm73pTnX+38+H/ugxu1QWIFEVMB4y38rEcpW9mID63EPMCy/760cP9V1Fd6
ByhICn4QB8iZNg7UDHR2KT4lIgbQ1vvkmkzz8JEGjsi/pS+qNHmUAKCj8vQM0Ju1MOO/r5HwzPeA
4ziSHwgxHDuwAX1SKPSOkGBz0cHtTDA31QQUky7nW5wFac0jk+hnWHUfZbPoQhLIgwv+PqLF+KBu
KTj+fzBoPo1k5urwke0rLg0gneonk03EaTK2h/ju7SZRtwlGZadN5vHw2hFZSuAYTo7klIrV9pm5
UE4s+HLtwzHBXtru6V9KMcBtF7b191vMwK8wn2pwHZ3fC5cnfF+95UsdTkU0Abjf1+lr1DgbxDJa
9PCh8ySZORvsUrN95j1nET4bXmdra1yHEZT5AtTf+mEnDckugyzCb0XNhzSCGiWvCbIhFKLP+4x9
HoWI/qndd19y6Zh6qhErdDtEW/RIALiAEINCX/OYXOIeBIty9pLA5XnbdVpKbiOrMmm1qthy5Tm4
M+ES+y2tvSKdy9M2XSm8eZvKWFcV8mOYPmYzg33hjeIFxFFv5BnIaT23VUZNrUdcDOV71bFdHI3G
yWS7pDqsk1J/8mQMrpI6/mgCqFMK7J280ip/NT/ZWX5nmv+ZwgeF474miKpr6EHgZZj/MlZH9Do4
OKlSo6L+mrmo2QLNc8LCcjgSc8H4Fw/8y7cdVze/eGPe/vuwEMpZS2y6o446eXgRlYk5MWSBeLuh
+hakI32jgExPAVvFs9Cq7OHNZq4WjJen3H0S2Sal5STItK0UFkTRWbRSEIvJqahPKSuqe0Hd3XlI
rcc9Am8kNtk96k9ZLIDK6DV47xorrc+T4I/XSdktYZPqRHmnIm3tzuY6fCSTOW7f68Ux0n8m0Nso
GGmC1aNQkKwDCG8X8lbHq4vWqPwXIuTOkQlHSsjQj9IBgv3drNa4q7+d+qPPvfFKKq+A0X6NrleZ
Ol7WxwCGU260wlorbm1G1TgieKuQMTQ7ilIiH0YxHYnOIjNbCExeCoNvpPaj4jjZibU3hs13oK2D
Np0Ueo5cVGk454gnJ69yM/cCAMfu/R3/dko+SJ0+wt8RXH3cYTRTXuowkH8PAbvbvbVNp/KcGUe0
g2m2UseLxFFKKxRdIh+GvPbMXdKJLZll612EfchXbEcai1hEM764sqFeHoLp/nQxC/FBdgLBsgV3
JO8C/JiYfZfJA2qWqjINIJDOPGwA1IYHE2uHWFsLFDqNb59mGyeZzUujGhoWSZ38/za0UmxjA0fl
tg2kWZIHxLYTqg1dMtAnq/kUWifIBiNsdbMDVnhVYHq3lp1Pz7Nt8M0ZNh3/JARxVfP9qFuMmxLR
PS4fnZdCB6S23Zou0CKv/kU9j3Ald/wzvHBGFYaXNYZ+FdlI9uuDR/426ZjqVJrTYgAH49iaUwkB
+Clt/f21BRsJ5HjR9MxmkLtUm8c0fAUmWwcPrgoyw34QoKqOOf3HfhGAvO9wPhB+Ol0xexq9LNa2
FoAjOc9AmLM4y3IwLQAsS6YKFTv6n/VLy72DsYStLm3M5RWTAuJRew6gL/xfyltL5NrY5K9FBjVq
rnvqT51dADl95iUirT57m9njXa8uH+bgluuUtyWlHjFFMk1lSfdcxZzM9IyN14l94gmXfkV51Qi5
eyoRmy9lwZeF+Jj3+CcfpitLgMDs9P6g9slFKRlQoJkWanlRnW42ROpF7BflTU2rf8nKxAzFupqR
5Bo1mM2IublbG1b5mKW7OQPAskPnu6OdGzsSJrRihWw5lJseFKrlGAclhrb45fRqRocyz9cDpj05
EkKSWyFbS31mIr2o31CHpb0ssT5jenbd5voFE04Ky7Mw7Hyqwhne9Jdb8Lgh/i7jxke5mexR0tjp
U3PDh6rBpvzDUkuIkaQMWQdrEcHKga0VqkV8pd8LhHRXghCKOUblv59Z4pTmx5/KAqym3ptvJIE6
oMlmzTv5AzoitfrmlGe3Wws06HlILrCSCzMSkjgzAuvjfITJUWSzCR1oP12nsaNa6hRAw35vpalt
sUEsdrNUYZXioIQtXEYIqHu0cHmOhsAbjOd8olOoazMqGSqh5qT/Oj6yKC0O8aidpkSK6C8Npdrx
XDUIeMiFUgP6RJEqWsIuayfLJ9grnwamsgsrNUHOOaAk9omlAElVuVKT15xCTbmdRhGoY/m0FIOc
XG6ZRei4I9gIpdsOZTyWCqgPVzx7eYNCI/SLqTL/i0fQrxkFdyGb7jDqCYqylE3j78R/V2gNLczH
HisQroqXPZvkIBpXU/TYnhPHEJWQyHSOrTvCzFoHriGPykfOFlDibXP3LSR/naAcao+fPoNKKtlh
TqWcfjuoiuFe7c4Ffp2Y1gHMAIvI/eZiTkSYDgXFt6kVq6wDvUfYlh9OJwKtP0ZDAyaBasGvuv4a
rvUUkyuChSqkMn6XJNwNnQ+/6vRQTyISY/Vd3z2o0DEiRy9bGLYUMplHH2sViHLpWJkd0gMa6Xx6
6WCRqKLTcJVYvEW9dPxjh7WMs2B+I5RAsPYhkChL4KNBJujvIhGv/hHrqe8pyPqAsjatn+hygcXM
QNY70G6nYpZcdByRkxmnrJgAgUsVklQEkPVJeX+s5FWGYp5/7DmRmmVFnvzEWslIHrTJylzilmno
+zkMtSdt2VdyL3u8sxl8q/fzp/Q5c+hkrsy9FWPh/WBqD99Rg41GYaQWaIboaawclqEj6gM8r019
gYdUa1kSvo26Ox/WufhNb8DFAqhIvRZCaPG/fXDLcbVMaAaI5bzLHYI0d6V8vMxIoFJv0lajdiBO
9EXjdb7oXYXCYmYPmNx/tGAWl5h74g9rZjqLCJfIEnSl2wub0u0ffKnpb3My2o8SBYiwYmpw3HBm
n53Se3NduvibjFdXS0PN4TJH3fMPIHXC+KO6FebNCghZ2XriT1AbUAjvESy3tDKVx6Hs5DuGV8jz
47Y71s3Y1OFtqVz0qlGzAtOOP5Ije3+mGnP/zpjOLhn6YZwD1XnplmXpJcJWzHqCXyMYVmpqDcxU
NuYHy3hjU/zVZK7F/addqNqLCZpH0dSmbvs5xB7jtEVPH/o5m6zZAov+dtezZvIhjBNsCov6uOEI
5x/4XQKX4d1ssrOASjKZrSsnuxzU7G2wg3/hGMEBF164NOqQWa+AyfRUnJPzi+CAYk8jB83V7UoJ
iub8Db+eVi4hqIAphCf+PZ67z5Ovi+XgJFmhkinhvA3JimNm1f6M4F1N7BfZjceujVkbTVOR45KK
4HfAcfGXEfO+MGcx1VvB1Lr8gQ8dLOlyNSHZnZkUBFhHXdG+LyI5MPBRcJsOmQficsaaL4IZMRxx
mqAv8jLolCeeKO6hJ2Axq05kjHSfaHQqDv1xX8L4yhBM4aZIy5GOicnW0e97mzOqU7naw+ValDk4
Ek6xISTDfYX4W7kfBl29ghjy2RznX52LUx4w4KeMQYUYCcEnDigDI1RNaxG3jfmtrd50vvVnnuFD
YL2EcWbm/lwhQIKxGdQkLpzABW0I4O3iXAZmlXXR2w9dvmqk2Q15qceHvIdcFRH15cPy7rJVIhsm
SUZe8aCfyNpeqfhW/NWsAtJIcwNXIKtgfhk+AwetW2wEnrUmT+ADjAXkgXTonMKOiMA6qsWs8PpA
aSDmdGCr26vrvICyb4nJZCLv0o51w7aN+hdsY3b3yFkM7lbYVB9OhDrKufyuNc+adzeVUW69U6ZQ
AoqmmCET6TX06Xj7yaKxWpTn7fR3wHf45be0EP0YYJjc1lC5USPdGkQr4ODizPlqsNETjzIfPUth
xSVg6YQJwncrn3B0o54UJmKDhNchNT9ZVzpnCUXwGZQqOjC3kzZXdk/sf3HUDYhnMPhgb1OF8Gqp
PG+qu6EZKVTDn3LwPtyPkck4G6A4eGfWfpvqj56gt0O83FC4JJJHRba4YYwsm+P1X2OW46vzxDEt
kudhd5c9SOsE+jOowktzRIdPqS20zNJoeOa0SGJkx01DtERxEN2Ccuzk9H70H6XwufBzmcY0pmnp
QexxOCMdSqY92TDjOpA5fSI1InJrrc2ee0gCBtE0xQ4eIlC7yXbUmIbEuSVbL69jOFnqm7OhATkB
wuzgOFS8wctd1zxCq1jv2p7gxoL90+Ldboo9GDQ27go3VDl3CybGovfg4dEbVNV9NbyrRXqY9NtU
q3VylWTZveAW9MYmr/6Z0lg8+9Jq8gbjxglx/QqBblKYIs9cbzRvlOjt4/zTwMbBWETf4UNlHkqh
0Q1h6YYj9h+65Bspo55xCA2TTsToAThGBm5+EgRlihwqtdK5y87UU4wsgJusA+KyW8vMivuKg1+/
SRyEV+FFJSlk+z81kg3/aL/dmiY7pqie69VPK7JUP/+zuOtJ5i7uLR3V2yBxs2il/rTOPS0Z7UXA
GTYSs/l3EdWNH9EfPuED0OWqBcVnbeEg6LcJl7wQm5EecrG4C8yW5i+6bCBDwNTEJ/xHfr0dWULH
JeAJXgeFLLKu3LlKZLSVP3Nsm0QV1YGVqSpzvMgeDYha3uNh/1AWIQT83tRE6kGlgPvgQ/y2QlhG
YgS4N6Gcxn5s29cOMV+21N5q1Kc9i1VdB1jjs2TMZYawp8dLNkk4iXTlG6SbTEu9zojNT4jOQ328
LQVRuPql2pIgr+9XkgKs0tMTJmmhiO+AYYctj9bi6c3LfA838KJ9f0unanP0SWO0GSV3GNRVrkM0
Z+zO6TW0fesAlRFv0q1Rs/+I/OZPNvuURntLRstvR7iFfsQ/unzdWlCaRba1Re2EkXfAzB+vH3hE
PbIm7nbrCHSsAl+JHnOb4ShhHPwNRX0UAvOgp0di6PdbfZIMPZnfrw8Q0WEjAeVKAotJX9sFlydf
OVjMraLCymK6nqPst/QcPwDus4ElimIiTP8JhYEd+Q4hCcBaCPRqjqLx4zvH9mAGmD/9CTWgAyd7
96jNriWiIROf3f4oWS+JYKDtinaCHDx/wNRLX2FkzPlt8Wdbp0i126TBUL+C6mYov2NXkVaF/c2x
aABcEvA8vCCG02Z1jpwBWF01Po5ZJN1fUh6Tv5tCRwlZINCRJvLuTMAcf9mN6bZ+paagdBTNEnFY
Xz+pUIUzVQCsJ0O6C70PubKccYiDsKBLLqFInG5nY8/2M4PSZ2vwXd8tQYWkIVsF4lepmdD9zDhD
DC46dBM0WpseEvxbhPG7DXjQ2PrTxOvtUA7zbkx/Ep10uJ/T+HDCr3BqDk4qlQmrA0OtZ/DtfvM7
jRxn8V4NNeRt7DYG6fh6rFClD0Bp6CVVRR9VN5oCG8cDiWnJarJDA/RxajqYhrKqTov/jZblOnQq
RV+e+vY/KVRiAeImjLwOPbtZOJrbWjGfiX3zwNsX8/jw4+BYyBmtn+NIb1hvUDsI47KLwAI/DLmt
FHWFpnWxLUG/UpbLxWWuNEbqUEITKlEUdPGBqxKutd7olO63MsQcFstGYgECKTd8vmX30mp6aKY5
ABA6NOH0KTaKBhi6+MxHVsR6EjHum+hKkobwkkmYVZVUxdYEp45h+UZzi0y61uL37XzHnuuLjGz7
3IUVLVOztGASxYDy6xr4O1m63hXIPPfb83N29J4MSaQ4O+E6jucvlq0ZRc3inrHeXRtoDeFzN+0d
SgsW/FzHf5+hCX/QT6EnXCY8labXmEZIk0MUWiEE7QoaZCxS8hL51XBuGZO91XxKkIwwgQFbiubQ
hFjQKgsVwiyRJCZ/tWBekvJ5j3Ob5MH6Dg7236VesYmj0zoQzu1311mYbVA4IixC3jAsDVNWfwu2
6KbyVzKj0Jdoix6WgODdS9NMrephV7YxT7QeDGUXH2TX/fpP2eJmXwmgi3vuyi4EcnMON2jpztFQ
f7PGZzrSzbgQGIIH5WXGj4P4o3NQwrrTXZhyumlukZHT35aenEMnwXOAoxxksGuPiMSIag426fIi
JSOqmpZB1vN7vXP4OlEDoH9w1cW401lqRZp2Yb1GJQ7AcuOWKNKyHovz2a4penW20AAoYBRIzjNQ
pwy4VFKJmwRhfifTVaoL0/fhwzXeCNKeCDulzw0dAdf7Vj6NfjlYV+C+KQW5Brsm5m41NjnJOWYj
pdsN3NUPEVCo9qevr9d+FMMGyogCuZXMJ1QwK4hQLBLsjlagjRO0RPvJTjywYLM1hweWvlHoJIbT
OqShQlwe2pLo/FcF1MH2CjYepkFtwuan2nlAU0xStcEChEdLDBSQDTuGNJuf9Lpga1KhB6sQbrVf
TnlFZk4S4FV6fBC8zuUck+zj0/LlCE0i4BemZg2bZA/2c6r+GDr5C5GSXnyHqyniVmp4pYDiQqmU
vPE4rubcgDMeVbi1eEjSYJjjVa9T9nvgiTIg0SuL0XpjHIAEKJB3PLgZju6wEJr/my39DsfODNcp
UqABZ/Cbutjm6IhVkGqEzwbp4194S6RGQOKk3lzN4WQXyx58PL/5pPSPpSEcqS8qlkHhBtgo2SRv
Eug5yHkkPilfif37MbOCQ+AUXrMkPGFH0vUljEjODOfs/F4NezvxP79BWKT7efDpvXSgR7/NlO8N
loa+C4/RYMeG8CAc2XjHsL4d9ZPdToCAz9HCmfQPf1OOmQz6ehbJnWubKbf6Jf+3+MtsyRFgEuOW
LuR/2ETOpPKLcxPUgd71uvrhCtca3hctPT1mY3tk5YqrVkDR8PvSAnKrFTl6/uZnVw2pq74JQ5uO
4L7XV0R5lh/syG4QE+kXwF2dQ80VDbWSD25ak78wDER5RnF9Vwltkgg7Qks0pNdgwTkiOEil7lCl
J/sP1mSqrFG5h3xvU/tQ+D27mVJ9xK4xIZUL30i0M2V/Y0MGX+QtHL9ZHuLmXqJeKLd92vSmsx6W
Z3x+t45uwZuy7aFGIXXDGLWsRIg+yg0muIjC/iUv2suToDNwgF+o+GHPUZi4EwbodZfkeR+vtuUh
ms8YQ8K2rG6DNdcb0BoLIvDeC8y22EtQa1MgVKWfEEzm8TjHNl3HZkyQpKHv4e//M4EqeVYpkVRl
hjKxgKOUJ07B1MLugjyz4hD75iY8qBQAEK5mLwEHMnfWkDcXJVRIyxPG07ysHeSDMhGbZNl2C1VF
+EfRY0Rv8q30VXqaoG9xpO5hX3XL3DA+m2VGYDQ4D04PwERo8V/UcQACASOrOBp0tatbloiOKyeN
o8OAcL8lez2wM3nkVVWLdBfxrgbyMc5NjhA4bzdVxcSt8BnkZtX4adHCHufID99rC/qM91XARqLE
7zYa1eMoZHEiI4vSJVtjUdTM2Duk6fBR0cgr9yIjEwO2WmMTzaIgzwk0DdbHFdqOX6UVu9rSuB1D
dUpKc88DtP/Do0mdf1AUU9wRGGaNtGw034Rwmea8luKaFFs9Mmt1M9hXR4XMubq4EJFssVa5Xl7R
Nm7McLwW0pw79JBVD3r7/CiH8OnCtvFvrLkVfkD2+xxQThTZhs3f6puZD5sUD1SyR5SNeNPqjV1L
FVsMiw192FYf6OJmNYpWxGsZPmYIOMqtwLNPmvZdjsVNjrOh3i5Yc/PBlxaqHPo8KnWZmy+7YhvE
kt4IZd8AHpjaNpDvzj30tD+rM/Exr3oIisz0Km2SgxYtjeCiBDEjlJTQZ3hGVTRHBAv1jFTb21v1
gccwbihZI3pFfSemz8n1T5+dH7N5xkBR906EPcdEouPlqQL/BEJZ/49UL1AMvb5EqBB/D4Phn79L
vXCQsuLh1GljbiOmZpOagDWcolaaC4sBLqJLojwwj8GkrATTMmyRPl4eG5RZOPWvQIiTWz1Fvc8P
gPY+lNUzke3AjbaWvulSgk6TeVvsLiSvzQRiuZZFWcSU0IBjg5XvVUt4ikFSo0K8EFznQXnz4icV
XWc/QNTT6v3LCW9ooUPocBF8fjeMOP6qrYNvMEvTPCAn0Ck+6F7TZS0/JGRR2KOYS1Bvlan9Xa28
utj5p8C23oEdN7ufS+JUdMYaVkssdefLnWm9fslFcgVQe2ARRT6iBQmAHRyNUG2c0F/5ZMeazWw2
W0SvbrNkehrh4iZIwVs7kLQe8gYYHbaA8D/Gb8X79D0b0mtRN23MVhd9UidF+aUfHiDIuew0Og4P
+5db+S+c6ls0SkdB4TqDTsoKnjbKy1M9/QrPSG3IS3owTDp8ezanAMfnHRZNIku36uBbi7zIpJd6
RSGCrQm8GyOPE7CK6ofYG1y814hpcAN8zvE4cU1bBig2IyqXuIYkHXVWBPBw8SaB9ZO791FiiSem
s1ZdsVPZmIi88211pXow+e5uRRPk2aUEfpaYqzCUMoQDaHHIhmGyD7xCPR8LSD1dMsaOCaGoP6as
aWeBWUAyqi94PXZpt8qt4GWCXvagjJKyEbos/nsBg8+KYhV1mIHpKRjOx4/2vckEkjptR22Xunjq
5BLYipAzq4GdPFInFkRzEn+KOO6ZFnzruT6NkIkgXPT6BCcDjiSUtw2MXyxPyteIdxNMgfJGvAmO
NZKOIN+81I5TDXFsCQ/2UklqbVw9vx5vPD5J2JHrkiWRDReAApRphzsnpnLKBybb6fsRlYwOoE9v
KfHKjUymbRqp9oL9HWhF9QWLbg1D8RDUosKzzYEoOYzQWioIu8KrgK6BPV6AIDyv/dRBq+qJSddo
C9olQRlo1OZxXZdFn5Rc43c0FRPv6KQryR1NO+spwiM8IkVLcfPWJwC3olM/6D6fLCkOEWWMufAl
8YiuwXfFlwOzCjGFtDF30renJ3J6GyZv1J7OIHzv9eyo8s2ijuNy2QiCFeFiOHA+R/Jur3YOuCTO
DXzZKL1kTgLFJaS9xNaA4vKxTMwFkmUd00LMSvA6qNvi+Dabrokn2hYCavDgXY/sTNlnEg5uehRA
5jCnXo12PWKDjre4rJLPpvq4oaULd8BSQ8QNhmKt8aNZQopr0roJFME4oQRjmf0GxgWE2q4Qf2qg
rtpXVKrR5z8oLPk0op3A92IryIgmo0GQAgTEepsRFDKC2OrU7dB0VKOWYFXALylV7bJhy7ushL1z
aqncE0Z4OqDvHKeDpnZDlZ7oa9uAVunn+pwfxnpw3kf3Yjub0es8koCLbNMMCfla8VTHvKEq5pi2
xOkvBWmlJQvsxTlDMIEQeVxBSETbFOsHnEdxpoE7vtzoBehfIbiOeCFwEwU3FRyIq0V0Mm0iw6V/
W2btAkBagha0bs4KRXMf7b3MYkovKu44wAHBhTPZblN8QbaenwZCSWGkwODOsYu4y3HH6kVlGkIa
N+5RwWZ0myGqAhCqJZG/4OofO9LBLetKmZkfiQmO129aXAnKShGgI0aL2HoODEdsXVMs1Jbiu5bW
RL4D0Wdfp80nDr2eqYI+J83pUZwfSX/CcCTNdm8X6i0WCoS5Zi0w2ARd3l8/pURaQPMQB2AUdql0
S5r/+8aZaQr/m+GAy3oUTGD2rvp1rPdknrOAW6or2DTr3CXcK4G8i6sUq4MfVivLWWcPR+sOag/t
E1trmuAblznMz65pejRuVjOV8eg03M6JZ6mCrM6mk7comjY9VXDV56nlDxk4VyFPSDkKdPEfY0KH
6aVYlnHhCif911HaPgiMvEuQKU1PCylKAllkk9KanFr1O8nik/WQkeRpfhS3yD5JY11rGktmZx0P
DoTItTN/SrQlaw2PE+nomTpnZLcJo3y3K8C/PGAXYEx4ky+J82hLprnPONLEDeP0jsVvesO/VM+o
GyY7GBHilLr36Hv5R9/FMlVdxtNFA6sWP3GYY631PZsdb0F5xDFRWpKQh7fzMF55dC+FRyxSJM0z
fAzFOU0NMcQrk5zAVdRKihqoErHp0SF2anftgDBEFbKFklgVZb6gqMGwunN1JLDqcjZNqhVbkAgA
6T6o+P3i90NcXMdXHEQO45JxXadrTKdimeWx3n6vorNJ0SFA1ttvvCudVQVw5vTyhigE86GepVI5
LsI0kZROSTkkTX/Km+GgPBQB1xb12a+/bqS3793tiisrn1TLnefpiV0vnYmGdFy5BW4dG17XDMel
O+PKhF2H5CXURDEmVeKDjuE3KP/X+VZyiecvfsb8PZ0VlsqwHcA471ntxgaN05k9lnMEIIwLdJ76
Ll4XEMSMiqGNTXVmi074g1okVvmLWQkfaqNCrUfTK7N+K7+3zSKj0K8irUxgSxgKgRXQmlI8Vrpy
CfwyKNZU+JFrWCNQJxWLBflBxSrg1rGCtTIpf330FB1wDFtu5TkVJVSsF9zJLDYTZv8X28at8ett
D7geG9shlmiC1F/amVMEJxcAE0+/7012zB7jUB83j7zQJh68gdPeGwZ1+nVLDXluoXKhCiNvOAKk
r5P1mga64hOXPNGiVG2nRZqEWGAfbYIACSiPrlsZ2aGV7L5/7q/GjATQfEZef0G7zG8DCVwGlYKD
lhuhpjEnKbIm1d0J3Zg2SM/MnfIqYmip+XJzIiVLL8cnFg19jxHEg/wMTFQWn55WOMW7wrlmt2wS
+agqakr3oe7UPGqVcNP5NQg9buyTuK5gLeJl3RKov8Ll2ggP9avAUYG2dtAk/RrCYljkYaNsNFE2
OXPkPfW2XMrZuL0VKB1GfGFfd577VSSaO7OHAvf8V1ls1MUg1lt8TFuxqTikebVqquPRDehEnoQw
cUxsNj05NpuaIBpI2zA4v+50gH0kUV/nVfk1QfyHp9icrO9JOsi2A+bBh3EYnPIHP/mBtzRleZys
IkTh+JgDdcui7Nh6m2INI/whhFrYUwy7ie3FnU67ZXkOeaBbbR5PqWcMGEAp7TYh+N06f5FQAC1q
4GSFe1fcgmNJ3MWbe7isXgH+L792iHYbM8Bt5zE37hnCMCDICP75S6SKgO4s9jbVzvnzopXkHD/d
nzJBwpUyusPZw23Yy/8x9O91ivfUKOFql96ohSd67w13Rb7lrHQUJSyt5pYrzQyY9CVpB9pHuejq
RbyXex7TdrUi7fAkZdKrSTFf0nnKc5EHEiYArfBFawTxx//vAm8MPHge6ab2oHuvfL0gvNdZZSlb
SdB1Yoxi7b+jnjQaAhnrGzO5L/xJ0B6uDxRjR3HgyBUylmhAI7htfcCAL7hdsKgLNN6PevvclWi3
dRtFmRaxZfnXEYTcYj3kIAnvidZjpByMlAh0qWbXO7NP6LOA6spCumzI11OwqpN+CZuI+bevplSh
joL2DpVi57SlyllWKf1Dc0SRsfUcfk/fbr1gXda+BPT6LVNKXteKAPgSsoSesrdwTsCzsM9K55JJ
vSFClS93E3N1iOMvBYJZd2QgeQ0cfCNaWJT/yaN0HNQywNj9mB1kFoy0bF8zPoWDFuDSOYKsERwX
OJR/ZvmqFCypkPICAY7QIfut9LIAuJDL8X7lHJQtbf2ZzNJTIO7Ia6eUoIy31OwQK4jZbmU1x5f3
ri4vLlu4IFzR6NBagPugUBEZzi/fS5dQxryBClKED1cUh/uS8Bz0RQDBa1ktWvH8Cm1rKAptyegp
pUpf4wchq/BQQW+xF04AZ+iDwGn7uqz71NAU9gleKFeCPnwTQGsAQlEaXRcXzNHA4rBcgmTKl2qs
qSwzJinoRGWS719SAw3D+b/rI5yPhJB7MXdajIUNN8EdffAbVIxPfSuxewdsBo7qR62Lzxjrg66j
co456SvlqenaVP/duIblVF37hvZgglpwDkaNEU3QxX1up6HYprGSBFKFgI+re74u9M604vWRag+m
Y5Yh72phg+8dIuYFZHG25wy/VESGJYKP353iuQ7E/tU3lv9vVMiIoUNzoZr/XMPUrVRjFKbEMuCa
vls0S2Wuhdy1dSjTajDHe7fiXBPg4lE8ewr8LVLzq9zcaEkx4yl+hef/sR4cbI8UR52URkZjgOoa
PcDQ4rBLwRiUG/wBN4pOSVEw9QCeaHeZiXn2srgvGp6MAVZ7rIiRDYKWJcy0JvfhSRLfznMrz3eK
0geBs45GHGjrcYpy2ejLwMVGVhRwVKB0gJyA9XEhhfssXKRyyuopQ5Gj/TBAcqqsVlqcU1bKcnl8
9dYIJljf2kE7b0gqSSkXqKEa04ed0MxFb+dEXQZELSTP1BtLPl4Y7fq6zEbsRPB7nd3xLo7Sk0nH
bZ6MoRwkeDJZIqQk46O9LEOCreJd7J1hZT6OIM99dtGsiuTlyUaWI5p/V4ZvRtgHHFEoK0YwHvRE
qK6G/TBmriIXKh4GTbI4bo2wD9UqbM6ozFJhWpMpqbnXbPz0Xiyar3AN9/oljY3Oecja422HV4NL
+twFLo1Yu+CaGQtVT+qFHBV9rhiaeAaIKlw7igbOJ6Z+yjGtOBMm/eV42EmNRDxx8lQg5QqggDuT
ICzrFAFWU3fb3Kg69wV1XQ1USpRU7IbawkWC5HmXmmU1ugqk7EATlg6nRSZX4tPg5Y5AIv9sm+KF
XQ1HhES62SdBCdSs65P+rabjf/GcMQEY79G+GGa1BoNQzNTjEKDUo8OgaPesYhvh0HohGGYGud4D
IUV27PBmvhDRL4WK3z2KmLu58ybJw4ONBsvPTETH5ZMSmeBfP2pDpDT9XyBigKKKy/7TlAqnNRy0
xnSbXCucRHuojebF6Jpw9jQTBGXJtpZWGzHQknwKx/Ihx9aCfrKKaVSgTAi7EfVWE16hS6SreizS
cUyUwa31gBY7LcESdsUW96VQBHs7eunnYTdlZYdIvZTu+w8xWu7RxXvQHhbi94kP3MxEvEko62HI
NAtLpjrV8N+bZFq4c5/de7GhM9G3/9V0oP77IkWFmOJQC1TRVdqov2klwIxa38q3NFmBQpJVbG/v
3nFhZSGbfQx5R7VmTTTstEGaXc3cc3+nbGa2RtnzN3AURrmK3cuX1FEcAM71IBumbkrxH1qsU74S
PS4rk1E+NcMZRONJQcA+F1fDDR5uBO7HZSQRv5DL3o0fHIInVX2ojTCzdd6ZFw8QbqomrVwVHw53
/Jbv0hJ3lHHmzMCrHKkR8iKmo4dN5KKkZF3j/Iocok+26NXzBSmLrOr4icglIsnzSqJNhBK1p3DJ
wAxTY4JIV2caL5bwtveakOBBocg80cLzql1XdgwIem5wzmtXwjC2LSwN+pPZEpn1WEUbLBc+JFLA
tYemg1gBzZq8ci6sS32spLSMdITIhQNEfhu4wn0ahthvG3ftSKMSml/2dS40c8mjNqCUBbebnCZS
trm7GW4J+7+Rf51wtqAQ5uOKS8tZSwsRSf1q8uWZfMAPRmTJfCxQ9kPF+YNhjVhFURfHg+cZvuCW
nOltYYNOy/M6OSyRmH1nJ585+UYZ+l8LdUGHNi26kgN1GldlxUiGyWUe6hIJRBTOQxZV1alwlC/S
ALHHchycE8zb2bySX+2Z6Yh4KDn1pMEiOF13cfHAN9bOIheEIIEG9HBbt8Waa2Ymad6//6BB4J9P
H1URWiYhqydPRYKolYTcc15sdf684bPwr9Y7oxeT4lo8LIcMbBA55Yrfcce/czO3XmsoljZ/wXAp
F+Nerqj0cQBVmOqrv+klUN/uQmuHqh1nmPlJ2Xdd+a6KUx/Z6ydFZ+qhVo+0rR3gYnFKuIrDI8M/
cx9wmVnM4EeHp7HdT9yoYTa6/nVe5TS+6VBsIJahFMHNlTX4twoX37GPI2TSzBpAlAHVuLiXSi+R
r3I1OJRvWdrkeEBORb+Jb5/NLOqae/JX1F3igsh7L3iX5mXpVaEd0lHXIj2N7GyvyNqYjTFpA6Tg
D5DgRAIAeaukhXKUogqSONPqVSjB7sPoVq/m/h1wJpRUJzURwahEw7AEQZzYI1d41blFsELkThW/
qV+08aGuIfulTCvNvx22DYqRtraZMp0Om+tbSYspFeQQP0iBw4sk/6lroMbNS7cJKnwbuWy62hna
Lji46EIsB8EWTF6f9vFamiB5lHFcVTgwhPu92jAhxulaDn3ewRIIKwO7ScLVRO0pCbblmm9kD6qX
F7ZZv2Y0Bc398/rRaOU84j4QLURg9i70TwmMMnReyib0n5iYwEBGeugTMwj/hbaoby97dbPoTAtc
W7HwEZzJBNwS0pSgNB9BzPYR9iRj9+gfK9D06sW+YQOy0WK25Rnr/vXYjx9lv6MDkBNGQy7ohulf
z9cdjEXRjsP7OSMFsjpnCa5dDq/hNW6aJRcju++MOwhh/z4ztWwXnvuI6PrSl63iF25dMGBRRWaP
2PBnvSpb1KoCgf6pZr8IYpoJcl51gG66ECAmmNIEUzpzBJH3OoxchQfF8h8Mm0urQUYck7uJi0HK
p2M2/D5TuMTybncheLGLKxXs83RJMSQljRK8SVqMc9F2K3xs42Mb08Q7Rxs9FTnFCM4TAxH+aTR3
RVWstSZ9dCiaypVkrh7UQJFN5hh4AL3XFYODMQR2JGGa++pljm7ZUFOxLpHJMQ2vuhM=
`protect end_protected
