-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
LIR3TtS28gXxIrvWpnJfvP7FRWzgsVjfBx9bMQd3iWgs+ppUSMIFRUlMVe8Qfxwe
G3U0Ld+hA/Mt02MMPF7CtuL1xG8WYYERjNSCHJDbV2Rboj3mDa8qSrz34WkUtOCp
lqWHPcWOQcGWF0t1JKjZQ35PJxr7rbMxXuWTJoLIGxg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 17472)
`protect data_block
yrXycFovkl6fY7qlcwI2X5Po6VU7wOndXuQgXlXpJDFetxAYwqd2SRfs6fdkvcfS
udByMECx3xDYZMi3J9Oz3vDHp9kXI1majNXVpPV8QF/7CyJf7aThCa3nmhgHoeDh
alLFS5KLTygm2cO4QBsIz5zwjlZZiYpDcqrFC+IgMVjrkOXTfewxudB2CC0vxFOF
lPyLJ+6AIz5k13bFgPDnuBn2ZCa0wkatIvmkWe6TSqCZjzkb5pZrvxQCZFL672pp
bi3MUEEUtEs3vr1ofrKUPC7o0fcdjQ3j8dgFg7/Ei2lwSei9igLE0oYaWVzorCq9
SH4Sih6YQ08w2euQoJ07uosOSyw66uekdNEoLft0GSMr6pj7nzfm7jOn0CNi3Bya
bpa9I7a0TbOO0UTADWNuAWaEtQFqkBdR6z8xv3TvWpZ9JeClmPFMgZhqq4DAw/N5
/Dovc76HECA3ePVKtg/KsAD9w1TFK2MrkU8j/L3IXv8EKnnZHVnfOIsa1m9l76G/
SzhQ73mbEgvzCZrbPOBu+hX0ccABG702QUp0YSshvsgkLIEg4IpvpUBdVIKtVSUJ
wscFUoRxiMPyGFD1lgD5+rcFS2dCA3PEYuaWKWjeZBa31QUsfzqzQqyhuGPaQ1LQ
3+CUrb+On6bZa5pgjRVtA+oTQiGrJX179uIBtdCMqcFyxXFRwPyiGacdJZJV/Dib
49VG+FEqD+3IJQXhNXqjh1nnxmsJs+JlgpIo5tctPKNkS+HU+8cbWWPZZKMDoMpu
l9n/psA+wqaMmwKSVkJt0Ps79SNHR1WpUy0t60TgJl2+sDD4MJw6zzDRjzzvTb4f
1DSTi4KKnEQIs3XWmuYO3WLdnfNvl5DtCsYy7Asf8oQ96xS4OHNQ/e6/U6QuQ9/Y
Lu+ChYqeSrQoOsSvsZxeLmgQEs5gQVfYSXJYqdCWfpP9gpzapP6vtrBVSg/BspUh
4DbJaG2uznKrcY66mlWwvxmfQbWqKAE62CuqJEnxbJohb19q3G97I2vI04G9vmVO
505FE/xbYv5UmyjAb6PtLZPG8phdamdRr4Bh6rsugjV598q2vkeqiPIoaPvVuGOY
y49Ev8WIOIoaPhlzo3JRcJeefCUIOQBpe1Ucnk3W2tvuXFmioXRH+Wtnw5snXfzk
xigVy6RwyXaFrZo6mvMMF6DHqeT0i3y9gn4ovnpzMQ3LZX504miT82JPM2B7fnuf
6HHzlKP5OBom6uyQDC2zAgEmMp2Kh3/gW63B1Kpp3FLVVOSIWxn8NooKs53m6Szf
OfQxLh3HAKDBCeKz89d0mS5JyPiQ/UV6rmW3qNQZp3g4gxA9eeKyhqWp1J0F108f
S2jhueXBbbLftcXs0YAqFnfCAeSqzJSUG2TvPCScCz7Fks+XOfYHRqvOaSkEf++Q
72QlzCEMfysGTlwlPH4aUcBtq0+nriLdOQ5I+u+kYiXNlboCG1jkX+zI0zWUw++m
hvTWW2o+uiTxfxbu4SyLPMjrbiFkcT/voJKnSDxGJlAWDjet1nHT9o+OTjHqRXPg
3NQcqG6fF3LGgylpY9R33eeeMpjBGR1VWizAW/ZAJyaHXJaMz/WCQGfvLFG5HNY8
eKI+ofHHfG2X2uW5SAm9mzWJD0kqTKQaU1QCUyoINNMWL7JC8AhctYiymXazQ1Cw
ePKlLIJ4fyEGAd9ma5gT1uu9Xx8Akl9/IANYCE7gIP6mQc3noiNFZ4/0iFU5fZBr
ViymZ+nmNj4GjYk989fUoL8EGMojwBrp/bP8OfaG0eEOsxcPxqALx1G67tyR7BNJ
HylA1rRFhy38R/wapfoa/bKJtwSokfLTXnF/JCsZdk9dsQWIm+yOgJBNgOseLE2l
vXzfv0e+vOBO+fFM+WrtNNFalhnk0d0jTHgcKOU1YFazn1gzsxlCKrUYLI1g+xLb
vNwsamJcmMBiKzaIrTp8r40WIP5Q7AnFsd5MoVJN04TTY9I1LpSoB+MwlBPmbcbG
NSzv7I8UqIdpgFnAMnG3zqOwDmXifVF4o7L1Euxy0kBYTR1LCTx7r7FWQ7afHMsN
yWH/cMKYF+fi5IGE+9xel/S1911LAmp0H+Pd1Xn7p3FFUi1Dvqo27WjVLjL+RnRc
q2VBozTjj0jpdKAXWjf0yR0M78i8HvuKkxa8ZVfvQz2VkmVEXSI+Oue5NMjtsIHq
UOyQqhUrRFvcfFr63Jf1TfUbGb+Z5jtz4FPASL65zo42oveXfJa9xlV7J4Rjkoh/
SMUotItvJpjd1cOx3E3FhGJ5NH9emSt9PqilCKD2Anz4YPjIAICEluxyXQ+YpfRr
vg7PLqlyu+CE2M/Sd9Hts3cdKuBGVBvOM4+12eye7MiPbVepykXwCQPWMSs45j9/
ex48UqWXWft3lrbH1YGGml9OiO3znfYr4fT370BYuvSGYw2ZVeJ7RN2x51Q27yo1
XK9MwpaiaZkz1MQnbNDgrqYD4r1WcdT2Cy7uLodwhvo8byx2cI/ppP7sSlm/rD7J
PtLs65zXAVnhRMZj6MPMa39c+dZ9ANNl1ggdI69ovi9vPimpQtNhZgMNDXEnLeZK
8noyuJSyh5kBrsf+fzZGw09SKKBMC5L9pQ30CWtSJWua4rkRG3M52ABs7fYhCwHi
UKZJAkDwBSwggyFjNMJRF6gRvKy2Xyk88MXIsVeKPhD0udGxLHsj0lthDMq0/+9H
j8jq/lSPfxJy4xb6WNKKu0/Vt5BiVOIquh2E/2DA2RykU4wWfPqn5E4nv3YZ4JpY
Qhtm7bw5DAepNKFjNLi9VgFfyGTKj+JpEtBaa4mNNhd2F9sukv5mk5bK32jvlPeo
cXj/0P7t9zZxKr2QPchDG7PHEYuEMVK6DaF2Lx14n3ofO+WjhGeihzYTrPlULcyf
0YBCAEGXwXyRXDYH/Eb4lH4u8jTwX6cVIdAkDM9t0CxFxLQpnYKzSjEUOD332XgH
r8GPECzGU32I2V8UmtRghIGWf+e5iGfX185W7BcR4kAx5akiPoaU59oZMsw1XtBU
MLkZXIA3TP+XDdexTk5fLmKGL/5XkGeneu6D9WJSov+tKtNbWfPN5xdG/wAAPmkX
omas9W629LtIuO4O4iVkDbACS7wn8FNtHqvhiCDO9pca/Hp4vZhtYMxcNN2wx6TR
G2rLkjsbVrPbZlBxNSmTicR7rkJivSD6hK7xlGAKL7wJ9XDIfAwemXunAF6RAKRT
yUMEnO/Xzw78zLTp56/KNUaMLhYhwq/QaFCJ/6nfixP9MUC0l3lQbiENosTo+SEC
a4iVdBugbnbVZoiKeEd7Y1k7t684cZxfimwR+VR7tKnZLkVUZPWYEnlRh4WwvvzJ
G6pYz/Yj3eW8zJxUyj0Niu5zw7fLsOvjphrTWuJv2qUiPdMz4GvPyCXHlksgLSE0
q+tGeW8KRw/uxhzoW1hq+xBnxjVcJxanzj30zq7faZpmMt5VLldfIc0C21X9Jlwg
jRkh5dtBSuNzioRMPpNPpNyeQoPhgjZHKs/W5H6dngpd4Uv9rJwKlgLzCC/T/y26
dTGCgryatWNXwOl9JqO5KBkxcRJpBUzK8QEXfHaXmCoFliHeNg+2EgM4Byv6sKHk
1j72tg53JDZyD929TfqxPsc4sSyjOJg51R/4M1foU1h8stL64iZfj3TkrdABjWph
Ahqs5sSCEycnvPj8xTmWblBI+1j6vWTZnZBoYd6KiYK/EPNGPwucU40LdTiEQHSI
mQ3+BRlKxr8Jxf/j8AQrl72PLd4aLdp1wMTuOYqiCmRzRxDhSpmHVyDCfxOQyrnl
jVBfEze7us4mHptcxlrzAWrBxfjbTsF5iU1W6U2ENIuEZtUWd6iEXhhz2PpIbcZX
wEMvcRL6G601NfYXAoy4eMmkC3xio7gGiw+2wn0Tbqe8yXNCWB3g9jJlqJPg8Lz8
c+nO1QqECrjpK+rk/CwhAzkuF/IWPjw+eSkyEPmJsKdvtcDw/GdYY1lSvdBctGTX
yX+w24SMPZeU8xw/4eTtDKjE1XDS/7kQHX9EtqxsgPg8VFyK4hyuPDaw3vjl+/2x
12zocaDZX1wM8MRdJdouMycHz0pe1Hx9OTbkAAvabjLsplobKE7sb0Zo4iENudRR
k/RHs7YK2BZFGZ4Tiztu/mqd30RnI+Mj7iJ4GNXU3uWEVs1Gti3g4erJsVI4/na0
t6lJ/Pph+xupq/fLK/9YbOt3BKuQ/kynDQMy+FEqkCwI6BmEBcJXb39b0GoMLAmy
yr2psr1+intu8gHYKEsAyjhmErwUsJH5oeKkxicXWQgv2xK5ruYHN7wu4cO1SKD5
2BgPUFtWfgmH+8OViV8D3XGkw4bocktSoRc7miyZInmQGkMGzzkRzuxALKV7WXNY
8a9+JdxCo/+M/Un/R90BwpFbQkQ56CtASUuu0gVWGGTBIgugCKAFDlRnj8KjQ29B
xXiCij7F6Um/1KryGPhQEk/yjkz1DukNsJ7F1XEYHgZhIbDiLW5PbnFFx8wDM7fa
2sNsYN6zQijYMx9P3FhDI6nTzYOsaSQouduiojeaOzp46XTonid88SQE1agqMfVe
VGksVCHrAYWtvzCBRRJaASZkqYiZv5M3YnaHCEWe6/OBcvH6Dq0jXj1Yx+rhSbkn
uexL3Mff2k/FOcZcKKOeU/jqfX0lkKouvCuwLZnkskPbr++Re0MhIOjjHnmQc5Nq
VtEiURbUzxQB2lIL/EpHSbJAh6QScxEhRE8w6jOPtY77oSy4x/86WeHI6K/AgivD
COkq6CVeStAiELu/OA8Fi3aAxvb7KpHyq1x+u6x5Gih24mTWkx60G6Hd53CoBpEJ
OF4JBV43H866RSP79THJqwndkPDa0PcpPGEM0YdlVXAtnuhdV06dmS0P/Y8zlRK3
jcK70bS9CWo+dbBdN6qe53Q5RuYgxYtfrgAoflz2YXeKAGhut680RTmMwER9CwUX
pKBqcHELBmc9MDqLX+Sh4/N1LQkVDAteTMt0h7E23CLZ+5Kdpq7mmCdafPWQm6TO
HDk6evwRqdRfxW4BeHEl/wXpxxsO+DqkRHaXtIwsESiBG6q+UcKZlQVV2FXZxr8p
55nxOu64m/Ws3+Sqoe7W+g4aO32W0EcrSHv8L1T3tYCEbO0nAcUZRwRn5snDVii/
yxb7crL1DlVosMXWNiqqmTPo62Ap8rjyGn1ZnJvLKCPwuGacEGafH8j0uQBGca16
wCqO7TeVamqRqOt9rOkHcKB5EXlORqgDlaCW3Pu4YZkY5TGbQyRjZD5+PDsNyyaU
oealjAzjNjPuqMbXSNfWVFRryYKRetzBnPPtCul1QA1XNGNuDh4tFsa8FA2cNcpf
XKQiy3zO830oOeTI6lMo4ET4se6q/I8EM94lxzZIw4sFXPlpsNl9ufiHL1U2Dj2i
AfHR/f9uj3wStjMTli28jXQbw0ie099qtnLEVEb3WB00zkIJ9Hu0hrIhHD2jhwbI
B0cEaJEW+sDewJDF3YlMS3AdxhLz15OeQYTz5kB2DvafQVP5DQZe8s32aAiU8Pot
tpXZyzz6QuMpE0DcAzZWCVkVpcJI/f3qBIhszixh1A0bJF1vOxvQCt4oHXXt1Gby
rx9VbpEby93et6O+oiQylwHzfc+zRL+Fs6Z8ddHDj/xZUFKkglhUPFS2BG88d2I8
J1dLNnO1yV0evRhmMu6n5XfBaGpq83yTxLeepkYvBC8KybiZeW3gV9qE6v4ZJpa8
fhhf8hhsn56OKoTZFQ39V3RJ/hNumeFrqhG+SFNwAtmFXeP8EstmYtz04H68dnSS
QmnW8O2SGprxpWMrUKUGbq47Ej4a92ormFgRG+FIiSkYC1CqsMoJs0oQdcnEcy3c
s3NKRKncZCDw0swzEuDNq4SgVIzWZpXm3T074noLsu3KpMRfPtlVGifN+PRs0BYN
IhGpBctB11a6K1WNEGBBz5mLrLaEaXlZ5BuIE/toJCrdCnef6b2PIK7HZMCoKUHz
jF/OTsGH9ar5QgUr/7bA5BLJKrHuliXHdcjoa/SJYgcfa9UDfJ8tAjZwqPvk9erW
2gRP1b4kFJSM2Igt32o3dTaB9ISR/Ge/aQyMQMIER7JbZHsmrT65xZTkAVxMujQA
IVpBa3WRCc/wJU0d6/cIuvOrAQKD7GzwGzQI9JRe8pFafiUesdz/c7dGhnclzbxj
WCYpMBTstEfzB7tK2YhXCEW2yCR0+GDrKdJDYgxbWR0EpLkfUDtNWlWr9NSS81FT
jJlmDzFdFvE6fKPnRca/JNGseRBMbgOrizhkT+sCyWbd/pfKPDmsfmXXZUq+Q1ez
wt8pdCxG7OSHUAq11DdX9pkAom0464ZELCuRbt6DW36eXBb2trzTUutz5vEtE7Q7
79RE1IzKWPLeh8i2UXJ4vayBiSA57l2rlSQ678NSm5+hobHV0JEajbOZG0ULqeL3
tGXhw+bcM7/e78Iyp5+4ftelk6X4n8fz+8jmJqGP7bjAEI1b0345yoVAwATA+PWl
ispsBlpQDj+8DWxUYvccm+mjJWHrVPBQjtRdT4e31AYjHkLB+P/ezJ2M4FRRdfxK
np5NkrUBMgDeoIOhjGz+51lmont+qCDjP/KfSOXcoehaMDfAw/+5JMyDprZlvkka
WbDa3arRa4SZzO//xBjfHG0bQhMh/paLfSqUqsf+fzFAYyqY6pzDcT4Bi/ndRsfl
4I6QVLvKxYnce2CGQKR8E0bJ4yFVNUwWWONHbHc5qg8yDuBXbb/d+YuPI5rc7kXC
G5uQHmzAcB8uwcDK/Y1V8vWbiaPawcKZDRevNUY+K3RBT2BMfTskUveC/fs7Llha
DG/7fuV5DhYSkNIytLBM9lk2G94uTW68RqU2S4ID3xtNrQYoHbkP6rZsEhsbmxd9
GY91Wp5z/zipgPmLxhx7HHili950puIbo8HAtkU6p9Rh0DcMFlId5gIeHsblxjek
qSqAUFYyTTmsbSB+kGmHw6BI1r2t/+bPpw42GZJK/Rk7qYQwfFghd24E7g3HQVdh
GQg6tP9oKNdyYPPNt4qIXvAOm/p5A3VHqULYaXe7AVusfnb/Si1rZupvg+FgPS0T
uY3CKvxisiC9AMY/eDUIz7vmmEFXc57IlLaGrE8+bzymiG95f9e0fvBjds+KH6Un
jvlSzR/7fzul1ZVLQ5yczfzVswTe1JmYXB0wQSdVazRAollfsAEGIGM1nWktFMNJ
GQaDTQIQ+BdE+NdbrR8JeTy7/F8ew1CYWR9GEcWeq2NlTiVfptfme/vow10FGkQp
mmqPuQioqsXEy2bY1lrSatR2I5YKTAsEVtTKQeRR/tc4rE3Qt6gGUh+29hVxRg60
81GWeOe1xEzTcmhp09798jt1BjIAOCjVubWQCDmriRcyTHcpwvaoD16MxsuGuoeY
tD+t8aH7sIe30H8nAZr3u6ukXJDmH1skeHuDIiBr/x96IT9d6fNDe6fF7H+I0wV9
oamsHqtFW0ElJK2G7ZHdtPAbeQuimWEPmnpTM8ylRuCdPBbEFim/JY9kOKUOuI2N
swK1lzKgM7IsXuoX3tRa0l+/bJ9xlAEvj2uKCtcjHfC6yyn665jB/xuPm7AJjRGT
zaHMBO8YA7MdGcd7d9AEX7GmxAbbpaV+gNeXzypRhNbKtO+jVLctWjcJthoJ35K3
W3ap1EPDsVlhmVNaHXe/WRXX1sA8Ng5Qd6MO6pxhqQH92ZTBPK+/+y9koiEh6nYT
+iDDg1kVTIGWWJQ3kdwLtZPuAMBS4oZZkkTUMn47eLLR2n4wXz5MfmTXfWOwPsx1
m4JpcBpYr2we3OMfBC4iT9mZ+uiAoFtCe9WXufWOMIEj29jC2aVdWJ08hSgygOqL
ULVnXoOsxYpjh09pJhYG1DpocA9aPD4pt0pfjSXWDyU2UmpOrYtVoFiOun8NFFgS
h9+BfXjosmdWb8pW+YAxtAKcW8r4lqczuKIsr/aq2gsampqUNT4voLWXO9UYvB61
aeXpGT4PHOe1ROhnUgFZh+Q12YjXqj79oAb2cZ+yPuNiAo8VmMNN3elYNF8Fc0UA
vAwidAagKg+RPLMZ+tHj7b1CiD12PV+FuTvbOX33/O68kgy3DnbLjQ/hec49rJBW
pp+9/t7ijFwCEH3BaYOfiuAYb2xs7krIaAomtf7eQdFkUfivLCe9fbvsxt0shJDt
HJu3Stxr5MwGqzNODCkuNxPOE+LWsFf5QrdMLKz+AhIAjQsPfCnaxLOn7FdxGErq
N1qWGmzzttG2eu+MxuQAcwNjXN3/Sk6qwdLdsBH1cLO7u9s5fZxzZKI3t4piJgKL
Gas1XqyLNjj6Nrna5/tdScmsMvyzRANMRSUuSq9xn55PvefZqDf0PJ4t8F9WjJUq
/zcb0VU+ckherAo3mukDDL5oL/DLhHeMtDHlriUIgRQoJ2p8cbC2ypccZle7TuAM
4nn68SWJruCgSXWddAzXo15Y9ieX4emtPT9j8s4UD6UM73cAJ6Hz228fP5e76uIO
up8ZbgxyICMAlaRjeEJ+4GF8ugKmhPLgbvQxVvkpJbTnBfKWAvuZ+CIAw+uoc0yG
cc68nFsHxtmjzeV+nHsuHVPxlUfiIdKz8GutEajdvPZnpxSMA+q82bmLuWtsrlkg
uUCJEjCsWChxK0BIkgnIQexuDZZuOs1emmLUzsyTFbeltq/G9UncSg20d/3uYDfh
dkdTavE6Suk7vpr55NWW2ZGgSLE3FLXEK0Y1gBJv9Km1Gyo9ckV5FA4BbLO/NQAW
UEpY/CWTH4MOdbVAYOS0x3VTUUL+uCKKVGK4xGINsYRPflCorEJlkjTvknI/Y3qC
rMy4Tv7ssTNiVSve9QVuI1GOJVtybigDSSsF90w5KESZJoUDplbX6dqWL1fRb9MZ
FCZiACulaM078PfLvQWOSCF1toJ1apJvatQEzFm/K9/WF8dbeoU7m9SPFkip0iST
SPVndQziUyJQ4pzi111rhAbWBVDGTmOq09eQF+RTYb2kNqXAruIIzUC6WhzLhZeK
UXEtecxHeKYC5JXI/OYat/YwZzgoyyXarbQaAYmnnKl43nuOt0ZJK4q+rg76EYJ2
89rvRVZFW063P2LrHHlCf+qXe87JU9xzijTFAkC6zuPh91b24qXiA7C3jpRU8CoE
QQpSYyytx0iTloH4RIn89U7dcOqbcSG+WWt+aZRq7LIYHtqPLvVcQ8WjftG0iL5i
L+HRdL9FbWXPb4ty802JxJ5v3T+KlNa8CJfbAIMjaf+qAy6y8J24bEJm7IxasVTV
s1CaNNhPD4bCfKgS4AyKJL05PjpkjTxUaYZJwxi0v/0HsVwojax5jnh6if1A0ZvN
H1lcXS+AZljMyKOy5qTGSekWGTpQuDuOEWHgjmgPOn8VW7EuFufe5hXug8mJGNZE
jfXSseCgaKL20q2hGLIN5PwFM9b/NrecBIzeS3LESYIsGRt7ZSciIhD6r8ARWh8L
EPgE0wGLv4pZ4/ov5QkYZ7n+akofhYd/E2Q6NnfqoqHpOybDsdH7k9JhjvC8uIxj
cc6fUxdovIozZrJ5eT4nDAbVYT3qmS4HcW6/pgwCP4wUxgk4YqRyYkM45qw3LUs5
SpsYpecmfhN8LL8obNd4krzgc/B18soU0UvkoeyV07It6Hgae9DrqDBN583jLU1S
SYpxYV/dbtskiu6mtM+fyka1OjwJAjTJL88sEDotHHJxLj+YFYMjHVIMXsv7xLrr
9JHcub+/4dqAC1VOLyYHWjOu8DPoJ6qkdrWVWpert6TO+9Lad2Ol+ja3Rb0p3Ne+
yS9+NYuFeqf83fdriv2C/KccGf8bumfxZdrisP6numEp56F5/2hQ05m+HE8PODlp
yp46N8d1rg515BSbt8qQcIaH0+IovuXXzza89rqRdsRuI9zFRy0xi2Q57YjejEhy
wNoVQNUz9rQ+R3xRx0104ErJjvVewK/Je96Mb2wcwIAC2s+oc9ToRO5RACRoYgI9
uJmaI6sTsnjIlSd2ydCzFF3N50jJpD7f3EeSuAW4DrlbCgHNqHJxw/KOVY89nbXh
GHC38nOfn1ig5WnUyJkQDuClhXgyqRc9U+pVJF5d3QEje6owZdE7NYObWn7D+XZQ
8cg76fkGWydEklYJRAV//zOSlZXFw5HbegwOFR5UyYvhRtXC8wWsU7Ccjh4n6BNY
Xx8wDNUtG9ZfMy1/dajXnMzolth+RNKEmxWOdgNyhn/DO1zG8Gogtj7RvG8OAlQN
Py+ZlHThjxCYEdrHI0xp+861UL1coOcVs0xitm1DPWpu9/mjjgzqzFCY6eqo18ax
rim9avmnLty8wp/KwB3ZZCUkqioYGXpcUrDknRb8sC+O4EMUxrd2xhPCww+Ayx5D
TkkG+cFC9C27GToRDZdo2oIrYTZmXRG2XysrBB2I/xybOBPPdMEvSvc9GK3Tp6Rq
wwYK/odalzG2mt4wOm7f1kSlL6NWTMX+7NuF0U4Wua0RrJ5znMuDjN8/uao03Xt0
DJ9u7/RLQTX/YMNOwJDobQfKVmDiDRbIoaULed6FqSV2xTv+zMEgnyEZYWZ4W3XG
hPkuFExDlZpiJ/Jlta0RWpl3ubK0q4Sbm655NwvZNCg2KdSkeYD6/tsMVRFDh6UW
sfQqNDy21N9azDEoDpmnrVh+795oBt5RmDcsVMMY8cm5pUry/xC3L/lROFXFH6gS
eJ/wfTs8K73FPtPYOWmpLqo9EUu4hH4M1ddFnO73N/kZ3MhhBXAKIV73Xt7irKq+
h1Pqq25FuURaMVy6lP75BiQ39qj+bOhH9Mw60O7pgWyEQ9V76DgM+I3XDTpUw+Ub
SB+RwirEA3GPRe6syOo+SUjo5qVgAv1icHeAMIl0y7GrQeAiYoG4SztN+JHQFrqe
nkY38H0AAdjNUSneOw6BXPvxnQXDiciBQwfpIadlOm9AowQZGDU1Q6YB2XQjncRt
jn2j0+KbzshN0s2qy3Ns36zfAG6non1eRPpZntXbN4cSjhBfz5Ms7r1hGpU2cgZk
wMXD5cNJyUen/WzU3qa4sVLUpCTQnm5GA5fpA6AjvrRwpj/ZEvnG3HjNvm9aW7FZ
EZCBUIeYvZB/tKy22MUGjUczgZb3XkSqvnjr9uW2KNY5SEB9S+QO7/QarbnLWBJG
aYmKUsVFonTrnXxxQef1wBSAAAQLJ4scG9CUs0kHTrYipF+FrTSFok2NTR/4+eW3
cEUIaglpSG3Ukml77UTzXsMm/RSoDy9zK4L796kHpQYx9lIOVybxT1qIb20oZUZ6
xQEFLMhXA7AWXqogE0wgHzcS19gfULEkeEu4AHZo8tmIEHTG3fcJwQZjg+AOLtwT
Vrk8wvz1wKZnSxiYVh1AVQhBR3tJvvYrpaFDnKwmqCkBwCKrQ6jiwsIXiNWBlmOr
YPcD72kSTK7IQqHIOZCd9XGHSR0nUqDUVEL1P2+4CJWEDTfb7HwBxBefngqgwLJn
o5XpOBVqLpKutQvt3hauWaBXCC2yR+DHXUKTLZAJk6wEjPuMNS0v6BTFlcBtZe7k
SbB/VpWemQG8BQbaytK8uRmwPjnsgSq0g9Z91x9jGyLMnCcERr0ee8aMhYOHquXA
cWJDYGQdUmo03QG4DEPv5HI6CV8wg46COFUXlW5RSKSFz21LLqq4t5uGdilex2sW
PE0p6cZi73tl0UPmd4lwn2gQizRr1564HO4QOIPTPSC2aoGTI6vLy8PCBhKyXXjd
oUZCiQ4tUN9YD27wuAP0Fp+qS29yNZqtsjFQhYBBDmNoTfVTF6Yr96lgFzJdjrop
jmJBcKfT87gH18H7RJfHwS/xYrTSY16Xz4VQ8LCGuaJ/oaM9rCNA2d9fGxXConVp
+0H533DE5hxkpIrAxPF0jUK31/6OFcOmOFkNCqVtLp8gEvahKeMHJKOL9qThgaDf
BXZdC8Qc6QJd28Kh+XdJHVgaHsd1hOugzi37CLSp8sgR8mdImuVNF5s0eATPmD3f
+Qs9Z1DunQNrRZE1ezz9gyZBDpaG96wOMhLS0q0PDrLoFMCFrkxrIkrr4WUEpMqL
8ulWiGES9W4K9E6tANGel1f+D6g5CZ4HDPzOExxTpQvBHmcmtu/6noouT1WRMWOq
gVdVDFqsqqen+wssXxj6jvj1ktQXe4zgUuLQeJwBaNlFTIylkS3xl5WwFfs2jfUD
/vd+310oQUj6DD6UooXPLNjzmVwiHEQ1GbmotjzJ/EhuQLn6uk6TpzSu7+vtkM1/
zbszZJMK3b6O/0qHSe4TOiUB9TZo8rPQ081Y4PwI1PlFOyg9PuucYrI9LU447D7W
SuReqCltNRJ0oxz/W6TwM+aV6hTFCcXNsjyoaO0kgyrWQWoZtfI66v7OWlOPgmaG
dSY+ZCjCOlBSEKo1iwMhc0VtknPfZqvGHJO4n+Mwg7pFFu+rzkCiDrgbwb4Y/DZn
K+opMmNltyiyOvKqZqYN5qH3G5y/dtAqRCdTHJxZgjMTHAhJn3GVclJxM4vgr5Lo
0yU9yj4VbV9PclVIM0pde5UPHhVmMlMa7NDP8eqEYBa3CgK74xK5uQ3esq6ToZEr
l/7nJoT+SGXVIbpvW6xO3wp/XM2TeC/f/0zZIXxnm691+Dowxid1m4UpgqYb54Y0
jyLipenf0BSdW6y4r9856jfAlr6nZRXpjkI2Lt8yr8FH+umWDLprV14x/6xGAixf
7wQu8FxUIRFJoBI6sLM+ungGQR+jsQMcxJecKV+sGJWN78vIlGFjDfb/FpAKiTBX
XxeKYoAKvTEfcffMwu0Z/iEcq28bGG6n80DWPVdsSWKurBEHSsCkuGWWZI+flzqe
crl/Lo1+9LG6c0EnsHr6iauFldHiuMrzM74cow0CR3/Avm0DkyGBlScSnEkfWdzU
WsR3sIS8CVcJNk6WYUvbZn5oI4/XFtTpHgytZaiFG6M660NQY5ODUjkXJ2uqwNyg
hhRTlyZ+fDY1qcBvD7YkLIoBkPCSPzgPjrI/AARXXD9XUgetSJN3mLPlGlSkzjNE
4lt6rn4lBTQtn7EkCpeOU0bGvivGKmqtil5hkVdicWPaId9ZzQD8KVD9apVkQwdg
hhZOnKNRDo0Bbpzz4vwK+hC1l51x/lqCF/xKc8zg6uBhEOINNEhH20kHQBkbZztU
vp9TPrFBPSHzaaTQRGM26FGuUy/xI//w0G1ZlwJDjnVdeOY9Yhh1ChuF89N95YF1
aDlKDIp1Z0SxaxsCCjZsXuT6zCSMuehIOZt27B/pOX2WCYSDZG61Z44/6TN7oK43
tIOt+JYttb47DAWbRbiLLFPJy7P0hBx94b2OyDFdTc0TrwqO+9KmrFkHUJr+uOHd
J6wuCcmL1GQgbhjSaMOOv6xlOC8e/8B6A4zsYr0KnyzkwCiiOETnPUzLjcpm0EMQ
AgdB59rom0t1gzhtR+Pp+mYfUbT52r01wamkZhCFHScjOWJpPrFD43F05QIu6VfQ
PuoMRqypnNbCAemps9u6D6UpoGH5tQGVxQ8X1Jtqk+iXiZ5dOGjwc3ErtECBvhYo
SbJ5jp7YiP7LFHWhhkh9ejbIvrfow5/Cfd7OFFyNfDR46os8T/89VVZ1eokviiNt
sUqlTl/y7jiL21M6N6neKat+gkoPSeaZthUrXw5ngJsAtn+wWKpqN8QRWG/9nA3n
M3J24IezzHnks+IgAuNt7Z+yDkJ13yAS7u7iAs333M+qvY57mn4EUE8HaigzRwyb
fxgqT8KXk2bzyg1R1iDli7A6pTvmaxlOMZP5qCWIqZBFZ0pI6iFjRIeLwxWqLQ/u
1h823jWlUHGs357KfKIPHe0nCiQCUZIoul2mFVHyIgJPa6Oiti3QJ9d3jZde/m5c
VMLpqhkx+S2q7YanpVom4lJ17fSiUjjfwxrXn3oH98v1vl0+TqLogw4Z068G0oki
J3MTmw4Hdl75PKVob4krRdHM7T9c7jQwZytU7ep/9RS1WuYt/mpmcwPVDpNkXpvS
WguYWQLaSiylicF3cYu51CHOZrdfkx9w/EwIosqet1IQp+jZQSVx0SGDY5jXK1by
xUKZnTiDR5S/VprvR9mkALhjQ4x9DLk66+TMFszU6sUBVNh8H6StyhM3iZ4JEnf5
fJ7RcYjKSMX/LJUkZOfgF6cm2mN6gQYqCqfaOYqPsgcHUHrhKv7cqyb6PGdKE5CK
1JhkXrj4HbErddeCRSnSmK//JbTjZFqk0LzYwgR1P2mO+dG1lUJ6EvTeMYmahotO
kpdlPtfgZYtJS8MMdQxM2SVDjZXYgkVDXxP1buCnrHJdcqakqqd+wRde9OYdXEzy
t7exo5b4/zrh5mvgzQp36Gv/NhD5Nk45FZVW+prQ1I8EjOxnd3B2kgNFPX3MWxVs
uD72n3/fjtiM3VXN9Z4OGVPHl+xUBQpfMOqKWAb+0o0+imgHMPS4iiwhKsJEvSym
4JoToj0PbDPefQ9FxgihsikdJIIYlIIaLk7E1K9unaqEkT2CV/ktQzS4SxMPk7Kw
u6dVwAml0LsxXCg45AoByHfEvBabEd/XyLQc/xcMjP4yS5FIhbpRoj5yFG9QpRo0
QGkjxoKfFQfz2J6pTl/cG5IdO4inIRGoaiIWWqrrtDzXOYlsnmc/6s+rAIoMJzma
wz0E09SG+aLGJaHPpnyBOZDcS9WhXjB9UNXBPpYiQ1O8hCxCPp5KoF0NjEfOde9R
wHh+3UI9gnXywjDp3EYgcNJIqStd70Dwxx6GNeWPXr3qoyhJriwsamjjHluN0zix
8NU8LPYgqGIk0GlMu8SVOFoQKmvbb2uCgksFhxAISG4mnMbfE0csvypNhaIVFUu0
3532CpHozXrNQF3jGniB02C11Wy4Hah468t9Q6wuvxxPstRA4Cqhiz6UrfjPK7ru
lhgr5CuzPodDzIoD24V0Egmm7o7xJqNtJF0EYHYJYdG4I0jBFgMtSpk0z4gxoMpt
maSI+lRfDsDYOOeVIFI84VQ3goCS0HIepnJEAAA6r8DySYD9zFdQFEWqOxnD63xw
1DyX3FOmnNH9RfhwC/WfBcgwCfa4EFDzavqtrSXioSuvOieOEdtmuMuICO8CnQpb
okT+gtV72JRAdadomgPIWUVxU2FQ5w0zaZoynkkkXgZqfM6HFBh3xRN7CTQLPSpQ
CmYjtAFdXyZ0x2VXS3P37YEZiIqvdj4nSb/SaY9qK2sWvZ9N/yFYKfwI0siUZNEL
zQauFGbQ4q5kzB6Pucwu+34T+2Zdkpb0sFk6Vurk1AEKfM+6OGkSfHgbXyvNc6OZ
th+JIM0xcolE80bfqoHsBKqbf1qpX+Rd+thCgSJDx6TsTURxfePxiYkLeuxtmYj+
U+EvQxAAdbMDKQ07l7IU6xUwNvn53G4zAUWcrW9ZwePGVFl/9enrAutvxk+Dk82t
Jjzq6J1mjU2A1PdG7+uM7LJek+3n1bAu5A6ejwByXkgNg30si9MAG836ZNmgvGtT
uTUcafXvwOo6ZO2jFxlA5eERmxcONJo7UlVVpi88IRJr7Lc9goiFYpgZAcG5y5hF
PJrfB8v6a33x5V6O865AIw9tx2Jcc1ag0Ao5YExac3nJ7/aBQz2NErHSsG8+4SD1
Hy196lVuFCHCgqDkAM5H5I9C/8g2JwshFOmN3Dn3RoYu/aK6AMbw1z/W4sVoULay
vxhomIjn+CFQm1wVKH2n60mDbK93Suimcd7RevJKTWIY30ANT3PSZt+upTmbdHhm
37JcHckWbVyrlNWg8FWCPO1wEet8WNUyxdp72PorkUAC7u6nMvC8b8zAdEySmckj
+jGLYRdx7ylofXphmwOBarXewhfPIh5FDvjnTmriqSHmK2CApJZ+Fir4yUPaRjJk
BC6FJnVc7T3i7NE3vbEjoJ7LpL5cmCnA+fgX+zPczcNeeGEQvBicuJPlS5ae8yny
MWIvnpXwKlcNPHTEd8bGKFihNOHi4/0oLvjlnPMuyHRRU6n+wlgqAo44tKeP68J7
TrOsRyVk1whXzT+b8H/KegQqcW4+qz8FOmLjVQdFd59iStw9LcDBPOTdz3QmQOJ9
NyE3uVKXztGHgC0AZuy1MQ41Kru/TlXyafu1lPbvcB5zj6UpTPp2v4BLqEwGvsNX
+GPYdeVl1gd+sGC7/x738SQUhshPgcXpfPKqBdNZsepXXPOk9QBt2aHiHpzByX29
7DYV1hmEVNR7UIZhcUq3tsCAtBkSEa2jKA76OcErL1tA2Te/UJTUHYSMM1pBdXj6
582DJfI6OfH7Kqbmb1gAgcl89GBclcqJ9S/c8qqLsBREzpXXQcaLyUhSGNiFqU0+
t8xTAehq/57uk/DD4GWQVfciest3FmZjwR4WUxiGFUS7KD3vl5Q6uM+sKKt2zwNb
/s40impzbOg+9Ur+iLehyGht+MkNzdXCyq9Q919XUokupZBICospXGqkffOG6dIK
4q8Ay68yW1osxfCso1vkgCUvYWy1r3m1nFvrHU4Y9tqkRKC+z7X4TH0oYMthUjjG
pnNOWIyfE0m6HJgIm7ohnWU13lNIPwEyyWLRxC+yXdl/U1giIgEI4maIWPlXnmh9
X/Fq4yOx2OK+Skee5/rwg5jkW94MNIGDrk7lOwQlbOwfOP5Itd8/ZBstEotNjExV
QsRK7OGw4hDTLhDL5RVcjTZPiLDNnvUmK8JGj6ute6FTkXJD+LN502sjmS7jjkbD
JFUijp70MG90xzNzYvwA/OyC3bglcQynizwAIBaLl/Luoeg7/zP/LD8ZaX3Upf/i
p+63ipk+lFnooDidkoG4Tngy7/H6NEIRvKwXccncEFtBmHoOvInH0iKkYAw4+9Pa
1vGX+Od1U1ncl3UYjPSZGQpAliHTBJThuGI6246+MyWPRYJpTwL7AiBUejmuQ4GN
gvHU5JYmpvcVweERM8FaoMgvnMk0vhvMfDf+qm1ou83j8cuO6dZuBTLetEz/MPqs
80sWGZeDOtv22iIVSHBwjG8YIN4cLvBy8kxFpRPvV34Ixuyo0MYftga88pcRCQRH
t6/bjJ0x5DcomDVKB7drwYKyuM9Ts+QY6l03G2xtyM16Ly2wh6anfHLfcAahbnwy
TEfncowOqTsa1MgHwzUbWs3Q0F7b2c9N7Q+u8CImdhgp7q2P4PLw8Fz//wxbS2/X
2tvqwxJHwngPHmTq+dJDCNqx2mrzj6xRnouR2qvTPz16tBtlRn359I7c8XZutuHj
EAuPE7iJApKbaJfbAh14GBXEXFe/HKcPc+lHSRkfxXVW4AwboHKuVEh4ggE83BkI
IQGbRCcUSGlfpZrbaK6oa/i5fNRGyJknBPdwqx1UUVx3ZNZHly0BtgkBeZ/7+q+y
zZvi3knLYXmVL8oA/IseuESe8WQVJgjJwEdDst+pRDJ6RnwFO2l63ocfioK4S3oa
TNbdScU/w7aS+ymdGWiZOatc7sKpwHidPtvJd9a4GZya9p0vPxgOhR8TCzAWEvcK
1k+LM06mETtw/wzyradCZnsWZuTxrZL/f93/QB+tj102QR1zvvHFBR0ielmrV489
SzVIlq+pTBNmy6xEsl0/3lSy2KX/DIoF5bwON+H2bHK+QCIXQuNJTn6wsb9Ncg78
ByaQ/rUPnobXl5uHh+ZIF/vveokaXnKz3CeRwJOei1ixc1Pr3Fh/bFBpglV4K4Wm
RBXxJ5g6iziq8h/eR6qyBmaP54OejbhO2KAcH7Evsc8ph2W/xQfbz0ewaMDPWMQc
vQzQW6xMz45J4Dk/jka9ORQ6D698Ry8nFM7nowOcoR5sX3Xn0qLkualjpDUmE5gX
ETSfMbwmO07I86Ln49ki7bex0nXXikYpnSi1mzsI/dOCb7roda2plMzrbId4vBN2
gSDXeqqVuqhbqGezuFcDR3BSMSC+pZmi+cZi7xX1/zvezry8UuKuCNmMAXifBH5y
e9XmKDtU3x8LuVUVx04gI1JGUwv0hyfj5QEzUy7B6d6A/x+aCj6Gx67pNvzL2UVS
ohSNccsRrrowYIPO8lOXy8/ECxFNX83PVJ6uNkH0ZkrjYHzfAm6/Vdn05EIazmKS
nZ2geSeHYwWWxP08spayGxIBiTbs17+Hphpg2BN1Nnm1VQNBOUbM2QiGqthCRHPa
kZyKqiTJwQ3spN9L9EUWug05DNjWKdw2xpHqaXI8cgGbhvn+9EEU5zlEbJ5yVMJ5
BfKxGj72r6wHCFCXX2Ej+ku099amhAYm48rR+yYHdiFzP8rnl5DJj96MwkdJkboB
ba+uUfOzqVgAOsqLvTkusLKhXONirt0t1Q7TrISQCizc1k7S3WuAaPvjlDEyN1p2
twFzD+eS1HXmSG5r94Q7ZLO+uU++8AhxlUi0oSLcpoqoOm4Izxxy+ek7AURFeIc9
2gCrMpC7p/40jvq1ZtaneUGUiq9XGrTcqvaJTFVeb+nhHAR+arW3UUFByVAiqXUU
4s2L26W/0/Kbep82564LaBEDNt0zVXHh104FSQM2ea3U2XJv6DGJBM7Kdvoa3Kla
OlC+HUObiJYm99agH2xMcsIqzTwgJyzQ1rKE084CWVAwfAW8e1sNLn3UCqAj+iYw
+EPQJqlr0fcly6XHQyLCZqqshdHLhBg9V86CfNFkZIuvwRSvgZeakhiwHwodHDwT
/3pQ+fXcMcZauyqnE9x4e9Mgs4uQ5tBR8LKxCw5KPzsYhrr/PuNm9zpCxEQK3Vpn
DNkHxcErIAFavHz8TberUOgtY8Y1FANsOb9IUHL0MxgmZHWSENpAFOTMjWTOGlOP
rOMibyBEbNf3tOzzeZLEvBte56Y9UYJSrzzEm/CEjq9X9mBM/b9O4kmucYR29TNT
XHMbKowk7BaNqQTsnIjREswm7GElquTqjtsTwPLKYGBTCgJHl0QcgLLMeDHEjGiP
J12PA8Zy7YF5hxARoeJyahMNdd06T3Iimrs0huIGricvmwKZmmmNXe7oOlfHpJcU
ryul2bdDaBOg2KQktuGN7m2T89YXpEVf03h5D9HEM93q5Cqm7yzMyCOqjourClfM
sQk8LP5Iw56IWBkZrQN7l0xnImC0JYlUMAPUE7Jhv4c2RLr6tJf93LP5IimoajwE
FRXcw7qzsgM5xZ8+E3+rqEQCzSvgITIqL/hQKF9ZkjjqNJyXmH2JkfjFCu+DpWmE
A28aiGoAN4OpEPdEEPDtyTMWa5G7GseYQDAuxgaE8KsW6qeTRn+ugzI25332y7IA
3zeZUnEtMBnhI8ECVpss1AGkYb3pGB5CLd8Tgken7oBFDvgAClT5dbpkveJ4qDbk
3tMVtiNugojUqVvlwDTqwxo4A4PLeF9f2mvgJfJDcMILLhU41rlWyXfXkfg9XkGJ
c3fP6UQoMwspmwPUkuDLOxIOUe5UbsAXfLY18kEVFdzQUK+YX3mD9QqeZ/OYifQV
4ArCiGdBcbhfW/aMZuZvl2XmpRe6sHt71H8CWNBWJOO16KfO8WktBrqTONcYxZ7c
P3MMOLuun+yFHC6DlxKQEtDRdAJGrfe9km1khbQugkYDCi6xzkVJ0TH3FtfviG9e
rFu9/E48bsA9MbALYbw7sTiB5A0RLvMAJkBTSNC+Y+xZxXXpKXgmINwIUuUtu/bO
KvX4GkgYERwNoFZdpfQYHeIcSkuHtPvDEZ/KesUr6847z0vY1mJgl9rOMG41e96L
YCBNYXni0bt5xZHJ2j8/YONg0TPmpY3ula7cx/isDBK2k4Zg2aTgBaJCRCv8BE6E
Dir1pSVo1eTUomZXYZxvP3+/6K5Beh2mZ246DHS0g4z37g44sgB8UYgzXP1p7U57
SUBZcPDulcz6e8e4FO3QZu5MSm62/9atarRkcrivRJIPiFcn4DC8CbBf3+Fp9Zyk
hCE+ebZu5J2p5DKZ39aGzHr9lF2xVgsvLbdnpfTnBUp+ShsROZ+FFNJYI0MeohGw
0+/Bb8toahgorrQkd5SqP1r5Ct+5hlMdKXL3Z/oj7e855imYhCvekbhhqkFmkn9f
RPPbbZqSM4V331y2DZxRUnK5+A/f4iJ3bXCMZQyTdKDoh1GzqifIL8yWvRHJM7iM
/yRNhbiJCK9riay6qNkEEpexi3hml1/AOZ56QPY7MVLJq4S8IiaUWW74fc6y7DgD
j+dXBQL3xVmrsK9o1mk9YMIH+wceKrqPvVOSyob6xrbJS/a3MrABd84a9aYamcU2
+DQZhLRSqVpO4Z/JDrIx/4qxW0+oA5l6jWI4YQyq/iUkaP4W4lQU49OzBXbzHXLA
w0p3YvaMXcDdqGtQ95Xr0L2kf7cdRjnCnWjB9Dlq9zSb+4X6cbg9tE05QJAnmx0u
h1v74cs5fpWufDgk7dYZaVGxavx4c1mk6PhrzvhkSAw9Th3fHUdAXLCaJDZE4Fvr
MrISXYBC5mOzeKZltnd6TC93PYnio2OdZQsXtncJC8xdF4C1onGcjFeT+jVTZQ5l
YstymUD01gbiD8bBFq4r/OnHUpf4FC17m77fOusp9pvYKkznWlxpP+HChoac8zCR
ShCJM20VUCcqblnsSk5ldIMR0PgfEDEZzVZTJ5Nb+8e/ULr6Yibsi+x9koEvo1Uv
vMM/JTZ2rjp7B1lusHwbjTw2lLe4P7KtOvJ8lj3MEh8pkyLsW5+Njxfd9QkkLjSn
OThFYCP3bQP/MySGj57drZCHcsZgocHPOwHi8uvZ8SILCpIHCeECcpLdAZSZgFBG
O9PjjLK+P1J3LZRZguVxo/px5abYMjdbKGkUNO7BV8qB8YU/tMoFyLmg1vCRuJFF
9fM/oRhzzMTTqEKTxCWZM3f7MHC0CMZCDYPFKvpS91JYCn03XkXpFnxHZS73NqQF
iW89hPBBl5kbJGrPvf79u86JLR19D+9wtVWn7fZAgm5XdhB82IYJ1/2SRNE0ysIh
RjaV7MXKfBy3w9Pc1ISHhITa1bhg7wwg+PCbJ0qJ9uOAho0BztGMto5o5hXn0bMC
6Cu1oDdRhOaaaGAFt5ZKMn2KAZfe+fQKx/vvJtzqbHCEsx38Whs4M1zpW8BbisiC
5uxpFdk0EwikumtEAcxz+ennxGgVRSyJogZ4NzRDgjPGhUIqYb8iqrYaIGryffg3
g+ictNB646JzDnU9MynvXHyQiQe/6Y2bjzNmT9XtcHlNeRfR06iMTnKti1zVuajo
Z5mg0B1arpSIMhAu21fEu5xYHn7C98fo0ry3zTb10YrNmVZ7c05ADL45oVOVwdxE
1MDMSUzhXYIPArUozj6T5d+MQEZATgK9stRxj4U8mk3boAtvaijOujQIZipLP9zV
7Z9s9lIssmeSJ9SmuewthqVnXBPjl/Dl4+YecTHmcY7kBpAY8XmJvvgGs2XWSUr7
RpYBQNeHFciryN3OQaib39HuOtQUS+SHH0XKP2a7JC/RjMK5ae+di9x93+CFzvCe
PNwOuTW7Cp7WJjVHStXcLTH5IP33xT4r7leiq++kRtNXeuQ+9HQqH26sWKKt0NKr
O/mB9qHBWRkXxnyBKKCdSb5jW9uG12dvDRZM/vmV7dUOXR2TqDNxZDOeIwL4dnOh
PnyibZAIJWMu3gw3fvIHZSfEiCrH1H4i8VbTwHvewR6uDSm9wyDtoYYdxm8UQo2I
JeSMrcmS1+wiKz1QqVwqwJCK6JJ/THU4zPTF5UNI+N64E96unjjNJNQhpTgELMmf
2zfFHETzfDypMiFZLsI+PNCTf65cNyKmmCPKnLnJySTUWr+cClmVvd6jNBf0hWF2
9M/13oUzgkqEyec522twREo0m2/8wBvVqxt2Vag0bnLuyIGPjhCN/azD2tE10f60
w9C6HWxg8y7sP6n6iFWmZW56Pzghmb29ErBGw/f+CrnX09symBPbzW602wditXly
EOD1OaIVjlhbaARLxoqlXIExq+RWenMRRrECddtmQNemh+O5yYNzmkrOyGpY+9br
/cjT2+gqNaqQretSc8nt6UohPcIme5uv+fCHlfbg0NuAoOAn7H7y3zsaTa059A17
jfvwXZv85Ogf1gGOc6fp81Rpm+BJmRkHaiVT/XgVkVa8f/eEnght++xeQIkdsqK6
EfdO7z6z0Ir8+XuDGgyxzXEalVfjF7f+GIOk8qYb9ntd3fljIOfXq3fA0GXzcaGi
hP0qtYrbMbMAfvtAa0FiO2HT2Ydnle7Sbjt/vDeck0wsZ5FVT2WEqkW4+7APnFra
yBoViyEXvpHvyzgw8q94limMkVNEGl5rPKX/qLjoWCGpoLi60+Z7nZjNYj7YpoFM
n4/XDkNgYXMNi275vi1aXcF+sZdF5+IJey3JyEyn80KNZdSlGunzZWfvGf4iy7Wi
qqQZQZ+5h9aFcCfvPyq/oJwHhdqaiJydpIJlx522+hDZZAJkki6PIObpVtOt2i+W
MJy28bVjHpvLZXCK1SFfQqmqYoYrnLSAHV68VfW12SWiiNxEq5dv40BkuYqI2whm
Fpnn5dOgYOW96/NOLL+H46vBOA7cgqk7fCMRxbO5ATTS7A1XdFRC21CGSnh8RIzg
K2cpzu1HhAIJb7GMvrizM1w0ZvaAZSCo9CMf2F3r9y9kFV1JlhFF/xid1YoLWJyW
Mhqu+tuT9JUztmsww83xPzOhm7XBJFtk1kVLLuzbntkuHT/af/gKcMWYuhheI4RZ
lF/qjcqbR3kTmWtVsjdgdrCRlED4+Cun8dS8rsmvhRNO/VWom2/n/fDFeqp6x5U2
AQKCGg/W6psDok6kYmb6ip68POmeIJwhGbY5wBfWp9HecLFO/24OvIKtZxDlQmi4
5jBDIQAv0nH5f7eP8oTRbdttODnq1ZNDTMJF6JSDdkYmnVNltuotficoKoDeyucx
L2b90QHtd29iCVuPdcpLgQXMpG5eoCUcPW0cEWjLaE7GLJMzaW1cWQPaKYE1XXyV
j5kNj2NlFD7sNlpYANQhCWRE8CbeIz1l8ceMNYHAxjurTARhF8m7pxXiGWhGROx/
IsPWErob7nZ1xBCiZf+h2JJ/4Z7pKOLaeDYFoAwxxtnAXOgSMa/gldiBTnQreUUi
skHYfT155LIn+pHercWbUp9KYaGWB0sDtzrDNDmruOMJF9alA9LPapRNWBXE6z51
oIRDyXSBhtTphuUvryPYOABZP+KIcyo2cWYimbRd4Uzkc15xocr4bxrUwKdjxxkY
B5G/yz/AGrz8OnTBbHBZ5eCUgyOAXAb+UU5/Y0H5K9Kkt3cHL5CKF8UKG1faNweq
94HDbiMhFZzEToSUnXhXHKtA2tOc9NqMZK1fdAN1B//nrFnoMtpCjjbGP9eGuVlV
UG56FE5n58KHCqGdW56SqSWdsLz1lHQ3pAgmzxyyPeA3FnkNztjgNYTjWV8cBOJL
VD0chMtX/lrA6cdDBaFFxX+aEwqqcUQWBD4COK225lolVZRIig9gZFVj1EUwLoSI
42w41weoAkH6x8JWSSNjrPwpZxfzvxM3khEdeM/ZdpMNcADEaLqnLqtX+9sO9sOu
`protect end_protected
