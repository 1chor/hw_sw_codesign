-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
FBDG4eFNNKuSjP2HqtCgKPGzSHGXTQVxcHMU13xwbWEtUHgl6m2ZzEb10PEQb7I2
89QF3ICZLFogz0QAM/L+IW46NxgU0eu7e7OlH9IocVxsbdl+EkLsMip8f3yc4dvx
lxGqdQ/sl03Z7FfwxS78RSh5/N7YC46QysKY/lgxjys=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 70943)

`protect DATA_BLOCK
mVSOrBvYr0qepRQfkIY6rL8P5HQAANAHFQtwwE7cIa9kHyZdmQxLFXoSypvF/Tq8
GJhg2yWKE96oCIN41ti3bwW00A4G4zCuBnI8w1g12HXA51FoHW4lKgca+5rcD+DK
3D0sm/zNYfJB0IUk3aClFHi2QUIl2ALyjsEXume5JPW3eD/HnGki6XjJ0f5FwViI
/QqRclITxEbOZiUI7RXnbomunELkg+MzV/wjIrH0UhZVWltUS2r1qVHOMhHQRrmw
ARO0Ep4Kqd8MlpNZ68IOQW75ZoragrDnTlFzNQbppFmvbzyxth7tDjm0Px6LRMic
/VZwp+sS4Sd6urPKUANJeO0tRTbO/RQ8ZTAqGQAmJuZUctfbh35rmUBbaMoDn0kx
TxKOw8aH226HEGAXShjwKEmer3lFCnwDavUwETYy4nzemf9VIGcTtQKtRLWBfxTq
MLUQtIu9ZAZ7gOPjhkVqdH5UwtDhI+fDrh3S9ARY5GF4MR2HqXgk+WoEfLNLqo8R
wJGGbWV3BTgFhpJFWgu/7/s1og27MEUVmwo7mDCsTTelS3+32VHajFxJEYwbjyYJ
HJDs7Iuwy/HfWoshpjNt57ZGmb/US9JZT76qugaIa22oqKnOYwrvtYy/Svn3V5eg
aop5IM3xlOamJ8bLbjAXXsnid3u0qY+nBxoTsHtKnBPM9aA7ugLIeQM37iTzJzAs
NPkYTOc6EhTxWYvGj9thLAhrZ//SfNLcFa2uqKncxD4YwGXXgQHRWeMEs9IrbnFH
RL75xI6JRJdI+VT9e+IlmtLhiPTVN8T4ZVQbpUd8gv8M5n3JNZ5i8WzSq3sD3AMw
C5Pl5jOFsogn9Zlgx4fdFW4emI7LEyeCMlhHmOJIrUCAUQ9Oc5rrPdBSRtUNxAnS
lUJHBwsGw7nRGX6y0+05k/0+0bO7x6BZXFYmY7bqnyAgE9xojVwOD+PII7ILOXv7
lLqo7K2ItBRlIq3r28P3FF2VUHPgkCVcFsyqrlBLbXyt0xs5y3TobnGU8w+QvAVp
vrGPOVaF55cjTnZdCNiRBIf7I8Ft4jia2vHpjvMoUF9kTEhLCq1MkeNZETN9V6b3
M+nR/qQhSZskGAj6Zq6DZHRVFK4FSCTFHWC7ETsHUNLMxSIN24xTN/CSGg5hoN9q
AlmQ1tfekdEK2ETQwkUxy05kqGqfg5ZCZIrQUDCqGgDj1HjgewlqW3wu7cmYG9Eo
uJwL0cB4K2iDO2iZiLDf+Tj7siJ5dBOGG2Vu+AJvIxXUiUKaS5a0mtPET8+aJ5l1
GzjZWYTSSo858S4uBiYdHh8tiudJ95gh5k+p4lTcBGaJepjN0tlrJ/tWvwxQv/+O
RHNBA3PNpl/chsVifiwN553X5k6vmZV040iUYhIpKiyj8FIfRirhYnyiqAnwd7mr
lcaoVbQFfKLbsJpy9kUE10shcYDj5lDECYUPjwwE1y3YAKQZ0eOa1J3XsAcwqW2r
SPQCKBKHmxUT5nBOdjCceS7wi+2souWpfincHKWBfp+AYVuK0iGINJEnQrwwOi9z
RtMvFUk8Zy6hNhjpK605I6PujGkjGqsfWqLItjjYxn4r8rss7sHkYQBYu8ijQ0UF
CDdGyVGig18m54f/Dt+pnepcUAGun3P8vhL1o/xES++5PBvvIkAw9kmJqFMUTQTY
b5J3XOnCVTJLfdO9djGB9RVRhHmP5vfh3Ori4h77rwUey9sASHBt2AuDeF6cHu+V
CkII32XWmFxqOPOLRBoZJZj3koddjod76kVDdFUU7WnhyUuc1w4J0l9p40Jtr8Ab
ILlamViCLcoRZ4jvD2kePutaTZrJc5GKg+4xHHawvXezOwc3xOYuR7X2H1K+28GT
sSQ0EpcJ6En8Ec+wP3kKIs77K62Z4GMqCnMOpEaVB7QZuJrYj6AGfMIAoPGNcgMS
zJYGK3POfghWPiPxWiOjRZFvSvEt4HoFo7HgcJpRISM8kG6EVP27dtLeuBUBT3M6
Iz0RrWxZyZ03pr79atD7ey95SIn8J2Os31jt84ZsYNHSurPMJCTlPXlHAOLjRdQs
WN8ifqO7hQ+72H4gCgWkTmnSrpxqo4RPemion84xeXE0OGP8orwtkFEBCkwJz/Wm
cmeEKlmU49HtzSHGTcG6sdwDS3yrwSRnYFqj1t0RYRnoIwmKH0f3TmYqhasA4idi
7AsUxq3AzNVSY0D7+1TQW6SrFH1DLX4omS52S/yFXHgR693POlj1mfCMIdWItYs7
dKNzEtyvxwwTYf9Zbcpi7iVNmsfCoyTTOOSB25T6+7rBgGgVzNa5BdDB9gBAwwHs
hHUdCioITiZnkV+zbs3/TC+LvYZ03re/xwLvxv6YyVFKKLhczzgxQYLK3bbcpF0p
SWiyvMeFSw1bviQsPJyh4gXxWidMcPzEHLsVKKx0RFJXQ5x3iI00MDj4sedsT8XK
kc0GZsOAA4jSy56Ew54YcuOgcLMxX8ddTN1veifHNIZqne3oWDmpThl8BRM28Gt1
xiLwn+o+15B8IRkYHi1EBkui/Op9su+bbtoUUZAtf6uVzxvm+L3bfPXbrFw+cmfA
JrhBFruXLxbz1tIgwbi93+lCFlFYtjgAmHcl3n4OSmuBpgq0CaxwG4Jh+5BDprF1
4Qxzruu47S0UMQkJBGf/rnTDAtU9J0TvwsxFwAJP4GwhHAobJjSETzLwmNSmBRLJ
KysrWCfT9c1t0ERxxGw6woA8CNqNuEDqxXJc9c7xvAX2nlmpHE5giY1VTcWK04Yx
XkBHzIOgxge0C4w7Ub1BIkv/kOdowU310g8S1g8UCp/oWGMl3mz9GDQem9i+k5CJ
gfj2o0sPKCZCZdRgax2hh2GiDMUKE7++VoS00k7bMNJDoGTmhiiIqL4Ef26mZ7wB
3tLC6D9HZH0tZKOAaaGz/JH5TuibWYMVGk90jTrcb0f598V24MWdrkvPz8tfwDWX
fb51i524wGG3uO8I3F8OqNVUNaEn5VFswqiZfvMIdTqCo/uV5i23EuEEX+im5BMw
hrqrRaD52GcviuK+J/SSlxZ7OPFkTC7u9drUnX8+fYoe5w2nB98AcwRjW7CQPpKM
9ZoO5q2zSTGuRsagiqRbtJtpAaRKWusFCN4eCrwsXxUhqtIpCRKHfRpx6glfoyoI
ikKPKJnQGA4EDUoHn8qeQVL++E+EOsgMYNciQqapLJsw3rTQr1H0KIj5y5/d7w5o
MvTT16iPTCF5DwpfpfRwLm5FzxRyrwIOZ0+PAEwMuQq9Ul7+1JIPTsTkbM3LpB23
S48PxseeMwmT0LNPqZpRxCM943PrZcdN8gxcT/eEdCDi/imXqUVDdLBwnD59QFxR
oUq0NzeiyHea+OU9ySKzu5aETpY7yqtN+nd9dVIwTtO1zL0itkcO0Z+o4gahNyUS
NmdwrkcqdTAZFu0QmLlvoU51H8q64xKMykahQAu8GvV28j9xeACxrsl9fes/cYDr
zKuU7523PCVq23qzj7OcnUuY0ooUMP3SxH6FO9KKw4Do0K8ekhtGJ7tbAVF4aOni
DntCTL5FoOviBgG0fXLI3dcViU+UeKNqDtSJKj8tYLzFxebD0hPUmeZcb9raK1SR
f8RWXQH52oPeCLcCW5OwPCF0F6LuLHbFxt/FX8erPTeku1/PH/T417ky0pjdwRgp
O5dl9ngpjE9m4hlqKGZ9clGPTuOX7BHunCxB85VSpX4QieXA7VELtHt4rNATKfRv
iwuFHdz1bnIpjL6bKClKCO5y1KuWP67oLNXl0flw3l0KRokkEZN7faiSR7ZNFrJm
FUmhKGPTXedsX5x/kpmphHClDmWmikjAQ/caYydMBxJ7OJHGH8SlytTx1OOqnp7B
LyAJejWKoOpwbZnpaXDJnmtxG9uAAzaJt2SIabaTsGUueGPlf4XSHj1uv7NsI8a5
AET5rIH8cz9q7AsBBcGim1YxaRX8DolyyygooYpVx5HrQErNymI4L5cOxPN2L883
2eVGcL8RBukkmjD/aI10y5nUxFI9znNsBWJrxWQKZzZOsRnCWE+pPc+79CcNLocW
UcIb3bqirPUhiuBBRGUh3dm+jk99XGliV8FkJLgRklUQKXGrH8zvPyhGAhsh5AMZ
wCo7LeFOFx5akHZSkOgDaNpwBu+spFGwxHX5NMLJtFdgb6ArUYd/uMVpd5jMvVlR
Z7avc8RUk26LHcVvU+V5CrBn2gTx/r0OWHJYzcrJysGOkrHxUtTAYkaX256DUVu6
q8MoGCHbqpyryMQhLOWUeW6OnapE3XZwRDc/eLll6wXXx572Ni/E6KUs+VPBggwn
5Ms4Vvv8ZZs4phf8CxI0f8AZkNpFKYnUEJresxmLHxeCwdidN9tqBv+lTHPLnFB8
pH/JEtqauGjbAzgD93wdfXwX1plycy+hw3mgdxQ9AQS+Zbul3ACWRThLjde+vDde
Jm2hp9xSH8vS2o4NcEKOK3zNByg7tyRnC0t9UaVJrKUcOqzZeu8jbvj//qJKIaod
dgNTM63E0wNjvmSwx0wR8njFKvFUDesSpuyC0TgWaziU7vI56RfuVIY+nu1oTwDW
XRbZZYpkd4SVDlfqEQhhzwwt0GSjkPYYscfTuOl9o0lQqTtAMFUW45cBqmxq1xNC
EheaLN778n9I+YEBvee3d5XRWS7CTBFroXJFXL4b29ivqHp7sKIB2XFvle8oJ9zt
rstnIPHZYlIloFeYb75we8+SkTPhuFHIw2L03n9VkXZ+cUrfMCSvubKZ69dAihgD
tezcBYT2T71Hw7cCGU5X+bTtfum3sihcFvdOabMwQl/sceadxM4x02xQ0Q7EFx1M
OWqZfa8lX8dQn6M/cOISQQX+QbHLcHh7fq1iWHzXr/E8r5c7P3zcFpxtBIrQ+wfr
MRfsRJOAa79WGLQU2ScxuzvXdBQtHYqxORUyp9a72/EE8o5yopNRdoWq5MYdpjW4
6VayX42v3WZsgN+LV6UvkA3yERrv88d+QMHRW67ClhGVNZCYPG/DHV/X87kvGKxn
m6GwF5x2x5TXmmQ/DRIuG1/lDDACOG0OEdZpLBrOynTxDca/fjzHvG1Bq7QToIGC
8yXuOCwxM+6UAZ1G2xW+MTOGyS1qj3dAA4B4QYZntAcqd32bZsvUVpihFweJ06nf
OiZvgVJIGnsiGL1Hsk+f/A+WJMqE86JaB2K/F8upO3kM6Z93LSj1BykXDKXloesh
tYti7sxQglXOf5LOJ5yU/LWs2JTpLc4JKjFB9oocvS4YVLNeeix9rpFVdC42tQAL
pNPW9c2rIx8aqwDB7H+leW2W3OGV4NY4Dcnv/k99/utwpnfED27ivHB6r/osWyPC
yCYJszXV+QGp7uuHXcp9U3DlPJ8NH+hidOSVgnxsb+hn0IjiKqTzzH7gm/G7PpQj
hM3UBiDjc01yW0zOFkW7BqJkeCscE3oMwnIqgqYnCISt6OcvzcXX14W4oaJ2mSvW
REDCGX9Ij3RRowQVSB4iTFjXfL8m7rx/8RuYboDrYvUmYAQPBnMkdVN239Zjt943
WZ3Y72hRy4fjd0qrpONSlyyH0QJyVes+SIyhlgjg7yLK+WQBNw3x4DhZoeM2Lv5j
VfkEprOjJac299p3vvabv8o72pK5uFcuIs1kuk0s0LVtzeZv4j5iQJwMCbytyDyD
7NuLquRHDliDKUlvn8YqLWX4dSpqDG2mue0rcwEsU+1PaYX5xDXhDQu+JyaHKon/
Lb7lHAA/V06LEfsdZMpWmVQ/G8vlnNc7HLX5R/ap8bLcWKsF9sU8LZLMmP4fPSyC
AxB2919zTpZkwJpwbAmJANsSCM6PrLkxlbPgCWXeFiZb/VtZg96ImVpvjJIrKfjm
+20Sn4DTOwI2tFt779Sgp6oQzNyPQz0oUBZP8L38vgBjNe2t3B/KflmHrG+0Ru7m
IcaHXXGHItjEhuG1q5TNWs+Jvsr6m9I67wm6VAjlS9SeElqqoZLA7T2mdyLxGPim
ArqnJpthUGKqmhROIK9M3uIoDLjnAexY/DnkDVJ/SmQ6PVFlDCZe/9t5oeuvhRtT
U2XNKwcTbjVabbVvBCerriGQA5CrM2LfVhisS+taEIx68//IgW3HccEplLKbuesw
qRGgwCrImW7I46REhJYcGvO5XzefcVx4Etj5MnudUAuxHm7p1oDgoGW+3cGbhiD3
dIXE3jeKt0JEPjUOAYBURi7epY873PXw/ohY/rNR8LI0P9ZE+8Ds+6wfDfSY8Cwf
doMJstoI3BCXJ9yWGm6YPE1oLxsNw/ODy/ad4+JWAgs77vhfZ/hsYZaS2FtLqb5X
lpoGf/nAMkq2K4LUki15mC30jNAkWMc7wEodBBeIm7EjxK7dB2td+cw0+KowM4Yc
f2Sq0aTZ25GaSt3DzAd0+N81NCISOJlDVH8CvVxyR8NWycsxS3/EE2vaFgC5HOgV
USBYF1tocAEyw7Q5ZEIVUPetj2VRuLjTqVp/MYqXkVl6XZe7NrV4FMvcOlcsbuea
wHTXvDjTum3pESA9bR1/6OHqbXxoQtVZctUsMR8zJhoRNiL3zij1lVJKikLVXqqj
dqS55HKKtx91miCtmhha8ZZb7GxIi8yTEyOHxegZrJ0DYsWdDJgn5zuSkkd80mjr
vCQSCoFaX17EpcwGHCmmxppqvCccoEbqme4TNxSGk6Ctg2m3oFi3Clnv57T8i2uY
S40+dP/+duIh+yvzHQkRgVofYjMctH4YJpy6R/ob137DPSScUu3cYUQuUzem4pVn
ULjpH5ni9aTc2rgzupXtH1kg8O04RNPuEzOZ8NE1x/7T8a79crCpztPXdJR5NIGq
uiz6JERXxTwJPFKsxwvgVyQ9nT3reXYJBqsRURVC+FPaU7+ytbssuYzNAxsKtTQf
1c4ieh6GrqdCe2hdOAJHMtWxyQn0IUs7bM9RA/OEBBxq3r4yWogTwxDtLQyOKxEE
gS+TJt+GSI5cmqDI0s/mRPm4p+TkmoY7WwME2jGttWHFKzFVQyXQKcwfqFay1mfh
1foM9Q6rVCus3BWu35hW1cOCGfYlr1RYEbECH/dx792+8AO5mXMLoBiLQ6HF+tEB
fSedSrYb6mk7XaM1c2WV6oe2U6xMH1jJUDX3kGKnT3Pxoff5HD4l22s+I5Ze4hkC
MCAmqMXdU/yqVsIYOtf2brDb3FncGepIcgo1vUmfM5QZrYn5dI3lYA88kvBHb3Ku
vRhTMkYUU33M65LFAUMdW0rFeVLGVGAJbZn9x7Ae38WSiNuX5Rry2aJl1p9GKUKe
HRiQsBG5IlVYTS31cNqVpxyDRxjxPWh0DtSDIEEDZFwvpq4buloUkCpr6sLZ94T4
cQO9zVM0Ra3Ht0+6jl6TiFE1jjJdwHiFiVfEevwGp1vvnMYypnflkBVZ4J2/NR/S
LrSMqb4TqwfORgvFkKe12ng106o1Uc3wZLCDsIY36reiGp8cI3PlwoZk1hhmLJmW
sY1QZc2+1ecS95ouh0Xd3xG84gzKJYZBnwO8J954pjm3WVjN7jj/61DRjtPzoEW6
KlhXdRAaWGFS3rXafEJR1AF2OLm5vA+c+IkzHrzMYAP4bsbcIx+KVoUIKsTbKcyn
+n2VFmZR4vM8d+vAJe6psE8J5uSaH/wLiyS4OoTZB8EbawK5D1dTO2TVA8NFUuSb
CkSPERFmoi2jxwuep1tcWetDtxk1KEOLW/0YS7y7dFSi0ibBtmLrIciLGRb7KO4y
aPLYJUwANb/fb/ch4UfyvNYCo5lfhRXpMI04S8CzFBK3UsaBzNyREGKCO9IX5OW4
k7bpIAZnIiDyODfbfEakxgGaOwen/VvIekXSYoJ9a61hPbhhtgby2fgqIK27vIj+
m9auzdsl8sMHei1p+01Wx7fNstT06p5tOo1cJVrO21ILRF97uthY1PbrzX6cqsyR
BQtb2gSJs0IK5s8eDeFyfLWpv/RLhjoa5LYGNhtKsTRGC5Yjasz0GBIZkvy0sKJa
uHt9k5zy8NO/z7gg8nn/XJBaVvqONsdNZRbiGdOzGzQ3KKNzxr9T0Eq859mTxTpF
gkAHKQGLs9Pad5MnApShWI5Amb3eZkhwXmQVZpb9uV7RQ8NOT0Nrdk5cKDwZGRNw
gGO8yWilbdAlF+RKlfCVO6ysyv/sNxr7fweZyGqBmis2JTLz7S0FcfgBSVAsalG9
umuoA6vbVI32ZNabq81YEJAhUGiurn6JdixvU/vynSc9FdzlC2okvlPJ0+lEbVbY
nNV3iMUg+D/6LvEiEpSatzga6TgmxoffYzdUnhB4LTGHoLVH7pSGTy/ZtUlca5+r
7zlf3V4c++rXpFy8rrUOFjnFu81QspvE2XdD/v5Vud4/R0hhG4JeNl0vKAhulmgr
ht8BnF5ik38Kr+bCA03ox9hutKzfhow1/PPKDu7QsFEDOgTl2rmH9LKU+tZ/ksHt
JwbBbVdQmzkpJXGe3Ol+YLH3OtNq95dTRgylidhXiKzihRJPyts14QUl4Xm9KF8S
A/HzrwOid2ag9yk1wY0gLJvF2J6Z0URtlyAHgy94RwDHtuMNjz+BRz01enU1mgH6
8CDUqgyIKAlb348yi2XkRRbLRmo2+UbCNNKhHnn/nG5cWg+n7cxbuPoTN2wy+iDN
f93jt15qtWvmzIrJQ1RahAUOw0G9EGQt/+ZbclLJb3A8LOlkptZu8n1jydCYBa5N
P9SdO3Xl2wly5UMYhXJkn7VAAB1vHTetj5eMEwxCqI7AfGostLEwkSyaGCK30esY
RPpcp0F8l1c2x/KQsZ7O+7GFTfUZ2nINX0XLLnZDZH9V6RVHuAW+r3644UcXzjky
KaHZ7dInSvLd50f/yKgWU0WeTMvOmIguY6V2mAsNkpUB5iU2tlJ6NhvOtfTmRt2B
XkTjhWc22zaXDfD0yf88KeMSalLiHiqDJ75xugNEqQQuOXoXpAWAgHVtOQ0Esx29
i6QwK91Nzdn7R7dHd3ipC9zbOPJwi5/lsQMSoGIEvaEv7Mj5DgS69gHWu0mkfopM
2z41eszEfIhr070eqW+zpb6mBiL1H2uDd4u0sJ4+0dxkG6QYd1foXpR8AAPsXSeR
ph/l65lcWchVBZ9vTPKq4GxF3cHNvbukCz1XcAdT5rR3tKL0CjNiDzesP2E7WSp6
phOvN0Gu4Kos0Tav+BQPq1HsAUvlylBD1Ri8HQEHLZrLqCtQrRehwUyT3qkb4YGs
Z9CJucNwYVReFWNqv9gLJUsecBalT3Q679G0/K1qcLwDUMgBev+Ay3hlJnmwcTLQ
pI8NV03xwGsCI5t+f+Iomo0VkGfKsyjjDgbroPCT0K7iC+KOLzhAoRlW+WrGh0kc
ZKp77IPCv+LIN+cD6UdOCuazvv73GrjUZB/Xqe+LHrv/1Oxi50w3FMoRUcmjeNEW
YVLhvLwMwkWZHpjMo+Ja4hBqA0kEFuhImHPw/UcRJxnxERN0SHS7G1Ivwi15g1nU
xz0T82VS1Ufup0VxG76FgdvTeRJApESlsVHJ4Jj24e4aQE/Rys+wWFRCWzgs2TG/
GjlEMcQeVq2XHSOIiFUOatefcGq1vRNk6jDVAG3eLhSrAC9ZitYVJBGcfu+nS3pr
6szXBKPi8BS1Uc/fgiWbbx0p3KUoqqhAxYQ+QfnCJcp68/4MnyIAR2z99WMljEgK
KwWvi35PAdzbE7zGJIUp1/rZh4j587He8Vr/6vlz8MFqS4ZzudjRYyOMsO1hspT9
3WI0wqOPdBRSVxuFQrq6Qy8ao1QIbTjMnsETE83vvNOBzz8LcT8DW3ohRRtpWSOn
95yb109O0iwwlh+SmA0EpWiETvokrPSohVhaStnMWFfZAGUlSuCyrUMDkt343r+l
BCL0zr91XZxR0NdrWEg2fxmBb9pjU5G99yY82fNsHBT1x9bPalWiNp7augeiPH4a
EfNeZiCGKg7QYiklCPdh7rJJNW9wgTIk8rE8sqEiiCtZJOVos24z3O4fxFlwTZ14
xJGugyPHgY8cSPwjFl4aDJw9Az099foIcAkjr9VfUxSc4ndliI2UV5DlKdsQRz2V
GQh7CwMcOSjHRpZAj4nrhIJsnM+XFBFscok299CSf/cq5vqQGe1ZMt2q/7oZ4dE/
bmeeVx+AVdCJ/O3rJLs0H8myrZKJbDpcXDuOWD6jN7AUKVRE/zV0YqiTBvEy+cWe
ccjiaDU48GRGJAKdl4bSQXepS8PbGYFyHm7RSD2lIZzp1LKhwy5sMMNWv80hgjOL
D2NngIDnT0lLjJzfroFYv7zJHD9ZrKlW2qoIO6+JXnDUqU/k3eV0M8SBxE1iyEFK
oJoVGT0vhXVhYf14/Bv9t9fJaayPXv4c5MfcQcmb0Z0HQPbOV/7kI5DpkSFiNUY+
oTaGMoebxJjPg7PiDGdJ0AAWpQyt3uQl6yJH35VIMQ85PkTEYUCCtcbAP/d0+m6v
0AmmZRW7ZtSnxjAHZ0+/mL0XLltxwKjnVip0xKzT5gz0zCC1EQc1w7o0Cr6sO3On
Yuk1TqIb8RoWFSXRsBkfn63BLFZpeR3z+bRTus4iRPbeIN0YrChi294ldj9VWmj+
nAojiuUt3kP9M+X2UFO8YxsUxG5eevr2lhTofOwzT1u3/SExisZsc7iIV6nE4lkH
DcDg2/1zBDMv1sp5tv1L5VhmuHx/kM/+Pur13I6RkZYt3HvVaUeWoB8pLl8r8Mei
++Dm3Afh0CAZwmhtoxttMXEraIMqm8NWgXJMTdL00ipyB6TbP4RmVtT62Or1oaEK
OVO5L3jhCppUzexOvKzalq4ZYK/jRH15Su224e54+kR5vhkVbpV6OJYstlX448PA
A6KCoXpUP7eqWxXvoe0IAF2Foc4qe1uEameKBGyfEqOpqYYLknzFwEsuW/XLMtK3
yMhybo3jpk2fXDHlomFdZ4FQSgwA/DnrM5DHb1PcIRJYSDNJmO1LHS8uqu7bG2xA
D+tAUftv37RbvL7VKiooHc7tMJswZWWa+GHhEc+R/xQrGujmw/5forVu/k6aeik5
XfLpJHwHv0OQzHMhNqDsqhwx6L23E6v2vbDdgQe91ClSoXdkcpI8OBkAcikY+H9U
s7RmOtc4H+/hbg8zK6DBz8GJu+lYoH8jzCyzBccwFffz0Gs+ytYjRum79htqcuWM
rHNINsOXS8GuOtprF0natYrcrAjWXqOkUqywsxFfRZFCI3pEaEnl1J5GF4eRrDrJ
uJML0TOkEgU7nm0utRyNkzElBmnFb6DzO2H06R0S0ggxjDfUOq3AusqfYbWWp2X+
HXOHDLYUDNOhIlbp35pj7xuT4xX6TpxeNdQY+b0duGVEUbyw4Ikbzgjdx6iUftor
yN3rFCPGje/0WTLFk2YqmaUAnnqJF6x975ZCeiGktH/6lYbwjiRW9tEgEQhq99NZ
gTDMasXlivL3YwrSaJLwXr2RUm9y2y8DHi6Q4W6imtGumoUSXkJwog1jUjouN8ot
x1/03vreov5NxW2NxLGHqzFPbHbbIG7PhrbG/I9gQTH5xMieea8N/mutwmtDqYip
AyR+hl9aPuLRa8JPh6SOELOgVVOfnlDMNJ9s8LwfZd/gV4BfTeTIyl4p+64AlXeh
bY7IE5tN9ZQWVaUlCxZ/5CopiFUxglol7aWNF571JH4Qwz18KPtq0MKdtw5J6uFu
CNah2awpk2wcS9HlEeMJb9WsAumtgmp2D8XTn/DqyIiqN+HDj3ozP28jd+qxPnQY
KES9teiyRaUGlb+b7YmqV829TN78yUNCn1eAl8kfvfsekrzTpyuvN2cjakOKNDa4
eokYTq9GOQuJSzSUooJQ6c3RYdiZIruDWthPA8lRN9uAO4t5L6gIbpIdGFpW6jbb
8FPRuoaAXxJZ3TO2w3yCS248Ben8WlDiQ+T/v1aWmFySwbLT7/M9xFgMVT7qOMb4
OodOwR13zOebabAsCUXOsVaWuB7oME5ZE3fZ8M4mWoKDNRWw2f3W8I0WIelJiCxL
oH9FdTH62z6tL8FeViDIxyBk3oG3OcEQ71d4U3GyFndY8mCEobU2lgynvecVAPPY
SosG4iyvZJ0vIleMYYoE3aoLbgbLdMENqOU76dAAaN7Qocs70/Y4GzBV8XPnTzWb
3sdeso/jGXU5pLyleKS4SCvSgrTm3543BpVchRxugHmdagtW0PBr5yFsrzqdAF0n
c+W5UNlDVVMWqU1B93akLZAwVGcHoc76tk2EmdQnu5dWahA9xqeqlTe4jeXN47SV
LniodK50u3PsKtyAZhzm1V79/eDMcU8xvZR8KyJUvTAxCDw/WL5F/+e44OpI9Mw3
ig3usUjxkU4ftEhW9BkmJJOeN2xBRXBSDeHVi90igIKgIMD7r2133C0kZhl/Qwym
QdygWiTgUqXvGNdeu+002V+RZej8xGxgiSHV9Vz9D1ocdbnR3SzggkYuIcuWGmcB
D5+q6rWUBIMFehREnuOo2/8vJts3FOhLL4LUjvhdTkasHNOXW4K7/OAtSVda85ME
3CC7Ju3fk7C+dhYZCQM3UEbuJTmkMUgu4iYmx6fuSAPfyW8upVxSKe6jMdOpAoi7
6KO6DZMhUUe7XKIB4R34Uema4mh7e5lU2LNXl8VqjkUZNVLQgGJylCcNcGbsDdWJ
fhwCxfHWiahf0/92n19MUtyHxKgFWzbbpJbUFQBJUNmArDiCvZ34QSk5pXB4QSyk
9xL6140vvv/ok1VWVShpAkcBmG+4FKdrOvr5htj5Gq7H1FRNUaU/Hjulg9cAU51t
bjVfDIY9fslVavtRaW0m/04ocwGWEWFRMcuHnnlWhk6IrUEcWpVhgZA0B3Dc8CYk
BNkVZgYDcje9DYckvOYZIiqVfTPen7sWoJ5NztuoZmJ9Te9gq0hEfpJlmCMgQ264
kHb8vADBUbQ1SLFwvXwFx+XB4IEI+UJbGdKlfkQ7EjE5ygF9Xk+OoJSUzDY7PjhH
ZGsLTFNy/AME0tCAkFq1xix2mcEA8spxy4CFYtZHmFkh9POjgCba99FnWcTs89s8
x1rDYDY/PCZcvKWthOJIjuz72I/bSwRyXrqnQJQbS4mSmtoQaMD8YsTnpV7BybQH
mroUVt8Gt5uU5xNeuzm3/HdNIXOKgeoV/+DbgWsRHG197qWk6tLiOo0EYJac2zl0
9brbGLPFNpH2p+J8fOrUsXCZeOnS/O1jJ3hmgCu2aLqHh9EwBDdP5jTh7hc8NFVJ
jPSlJ16wn7MVArTvm3QhJjax/XtNiRBsoPWgNJQgDIwaLx4SJTuZBZ0Z4QL5Qdqi
lZTCMNWaTLHpYPjSKSFeO8DoblAGOOcjT3+LR3jaXc7TRNYtAShI7NtihsuIw4h1
bdgk/nWDF/66NKfw/ElPDv/pcdZw0PSexOO0NxWj3uotLtJTQCGebSVfR4NZL6jk
qweCDtM5cCwkI3N3ycEqOXFhrbr6TR9sVuHA8o6xYp+8/aoBAclQqqOXUW3xV5WT
LEwdJHmH2qn7AxK+s2Qp4MD5NCiT2OrCGZrsMFr5zCcf+Ip/vTfLlMjyokUiP8EG
HLsc+bcD3KcA79DMUHpxY8gUr1G1/V4vRiUNskoTuOaanKLGuFTsfeOs6+5dwvV2
t/QpM8AtqwHspunA7QCy+prK27yWuv61+eWaFX2wdFbuedLqwFZoZyKsC9N5/fk4
Zv7+jdXF9/LDGtef9Ly31xqRlk8eAYgtxOYRSBuda7EeW3ZUGXHU4iwJatF6H+gD
A8IM8qJ0S8YhsKEJH+6weTr1qDJjy5g2LKdQrpQjEG2WvPaydkOw0nB+vhvAAteM
xNTGoHFlPN+YWcQCWwEOjlamU67LthdGlHtApmvZ/sB6yImza6MKI0fYhYGwxsjC
ofL6SrgiPBD5zXCiNLmc6RBHlzZvKAimncGXWRdr/plVR5pILDi3RU9sm52XXg3V
PD4a9RPvAyv7pUfl7HtDgHK7CGKGJw87drEn7hM4QR1FG82ii82D68WTzg+TWRyi
uvNC0Qbx2KP/aQ00K+6NIEb8+5Oyg6QLILPA4ppx8fTLbDshZzIxh1cxCirHL5UD
mOhV0IMOLXv7iXGzuZlZIBnDhFR1k+hAkET6+2UYnT5t1JMt37KzvlYiZYM0m/3V
DmWgzCPOP3hsK4/v7WjbWBwJ4CuRgbOu3LI/JX8x5eayHH6AA1lvbF7oeD/0fWFR
oAO+8NH4eguQt6gsGBxIdKP7gI6HSDFrdcR9rra8mpTfYR8rM+OyLn69ebm1DR9w
HdmmLynFr4TIAyGgksWDqzpVHTfE62uN5Obzia8IIKrW4UyYCSuI8Sm9iMtGBZDZ
vvgp2MEmqHV7HxMZyHKos7YR8j9yviAUpFyHWTuOD2u1HSI+XDjb/B7h9qum1a8m
6GVYfmjYYcDD3hcGvF5DaaRPCWulwMXzfBK5DliVZ/zi1iNl8xNkiKmBA4pkBJwL
bwCJE26536Gg+D7f3cEGqDVe0JM4dG6IhX0e7ewxWrOfZOaJ2oPYWlXMt8DyBVEa
1zcrtICoIOmsTv9yEnL7LK49w8UhA8r5Wr7mnns1WkbHeegYhilPWpkhabnViKtz
cDElw/JTAOXsonkgiwOYZZxnwVje+GyYuIrfSMgP2MFuJS8E6241MMoqmFJ2TQ+F
D0mDZiXsbxlYzV4v5lCR3ThqoNhr7r5C5+VCOR0ggD2dyJPx7hApGRToieMUC3l7
egPmfBWmasBDHU12zJ1j4GUp++3vhFMTYRprwDyV6sE6as2ZiyQXJi39vldWo2ZH
UP/+fUYDgiaVH8/41j+XCiJHKZ5RVX7VexywuRPFhlsCSHKNXm/yeWfffSLEU7KK
1wRIuSHWtxZFDM/nYGeHSsQudB+vZhdperfiDRqOah3bNMa3sFZM24REIuMQVTKe
LQry2354ydw5r080q77XRbBvoRaMeSHVYI4Z1V8+sSbSmppjXDbA3TRA40Riqfeg
E8sUG4Xzt/I9WnBABvcqZVfqnw/nDQ9y0xnvSIvHsHU8ly2OBBNuRzjspHeDfTIy
icgoT4k36W4SAuqokqqjEIAENWcAtmajrj/QVkM5CGzt5ThDKFo1BtkDpuoMPTh1
zKa1ZQLf07PRkiGXxw8GvHbSnomPfJfx8FaU/NHP+yrgMCTEdrPQa+B+U8vw7SIh
P4fGv+JbOPAv1KDWwdsRTJQhaPYAgKLoAFgDy8hQmCMu5y4Gm/ib+gR9pto3LZNZ
edJjCA9uDv1zqkTRma1BYM7IoAhveRJ8WKes9e1Giuy2uuu0tJja1so0OT4ugHYO
oYWV8gzzKtcQVI+ZSt5Z/Wzcx1fbIRi3/HVjbsHcfaovmAD0LT8h3LC0zMRtJmGS
ZgZTbmRg1ysJBjxduCSZvtzi/U9zMPfIMb/7U0tKyoU5bdUgi7drGSKcAueAa8s8
6VYT/nlIlgtjRZjUe/jp2/RDuVDKXYH9Iad7CdqCORXkJyjlrV1eEmd3KwZWI0E3
eAPwlpQKMpc1nbZptdwBw6Kx0lBGDlTo8zBJURauUxYX4hUvJ8mVo8iBa/ATh4qc
Bk+iw9DOgf2bI9UX7dZD0t85zP6c55KxcVHfII8o8T/2bHVxkaO0bbOVnx2b0YKg
TCaIGapqcp3ZIzACrBBbg+pIfPzi0TQiY9ej+h/ITToeUjkt2QWcV4rgPXmu+PvZ
MoqOcJboarKp0ovRTHBlLJH9rWbra2C/+Gg6D0jUKES1IFn8dtzP5D28WbWlYrCt
GtjcmUqInZhcIKAzpkt3NeAKaWTU+zDTQUEJNyU6mJyn2Okovk/yHtbufzUQxoGA
ZldbKbxDOq2zVWvb5tURMcjLXGMppTIk4z4EFT/ZDb9YCsCbeozPuhtFhudYpH51
SwrtnKUL1hgEhhfyqiCZxL9v7mVBPPKunDHj4SMSzIRXLmND56XZNT0eSRkh1ElR
bm+fv80gNS/vDZbG5zpZuZ5zJk6I465q9uS6DabWlyYBmyQCV3HMavNGS8GFkWmQ
C6qhsNmrxQVZmJXVZ9csA/Mzz5NrECJ99+wgBAPoytoe+aUuUa6U2z6A4/wEX6jG
1va3Nkn/xp6MwiBjro8j6Hn/3SGUa3TqtEKm6hyVZD+KB2cIHSRemy3zaD4d1Ttp
1xg9NJtuu8k+e04s5M8n11OTEBPyZRex7k/75uCu9YerIOgNEbZN+AANOdAL/Ifj
qGGt4CjcWkmVYOgUM9JTjpz53CF6ogMFmZocYYWzge7BSy+Fffjqwari2GA2I+q2
0jtxPrfCsHGqEQKl8dMtgSdPanbbIoU5YwY728byyYsPZVMmKg9+tjasimDiIoBz
rt6lcV27sp9ktVPc8XAcjlLz//0g9GOpuQc/LZrpRp6yrvb5ui1Ug9sEllCy7Sla
bS8a6mSWprwBrHD0RdBFVyrvFE5KMHDAE3VAvn7axnLjSn3egggAEkeLdF2wl2cG
hkvi7F5CJMbGdydDtHEBncNOGWlZge4OAdzDKReEY87vkX2bfMMjurbtzMgSlZps
FfaKDAa0XfRwI0Hks2btYnx092Pzb4vdiZen6x4WInfORgViZGG5w3YFlh9W478u
Qh77usodlSn8rxjgh1zLZaxXs+FX6SbIzCL/8zD6SKy1ZwIZJkz6DHjTJCGchGAD
C1XUoGrVBcv0oh6iT8btCuEGCjcLCmt8jFDVlqELby4olqRigrwxVQkTHdqa8nkj
pal3DDeitbpwjXmH0WGwgdi4P1nr+y6LKSqxylHp+tOh5+eGorRHufPUo1rHpPj9
XyqgX4E5NXJYqQyEwjFw4w6C4bJBxq6I/CEFkkOcwNFCWTkCZmttSuQC4huSUs43
KZ8kwXmBS/6W5o+E3EIUS5CtVXUBIovy88TZQmuAu5sa4fIx/nw3wGhsmgNxICNl
NuxdCx1zq/0xlPE8o4ihttHZ8CDewfLIb+iUKG9To8sFmNYo3sGXiRLgh6VByYQc
jQRNweR83644Vfeu9xxnSztNDVxNma+YCX/gXq/UtCgUwm4ts9OF61M1nMinQKO9
maqSjLCHKW6J+ND8AxGkx94S6U9SR474aC7Ya0j+vS92CuhlOdjnGjMV4L1YSRLY
qkfNO7YVbmvaA+2mTwLx0DNDuAi3GsJt6ihbaN8M2vb43X8HshGocer3oCEX0z96
+69iq+fP5dWcI/87jUL5k06e5dKD7X4jIUwGs+E9ouLfRUrqrrBoidPx7BT/iQYp
rQenPEv9+j2p+l1YReq5thGeobjHFzSJn1u4+gD3xiw/EvyWTa2vOQ5xaZQOCqpN
gaokhFrI6o6d9pxC1QStfv4urGkFDyK00xv6tHG9opAMyUr1eRoK/Hh68yznQxjy
1WrX15aYSe8+JPMNoPNAJObKmTpqrCXeS12dRjzNqRn1VWR979PNXPUp+hbVNQnj
6z6rmh0/0cC0kTDGDPCHjI19jP7HSI5bVN5No8XvINeN6t3tUsE2vL0DH7xW9Cpq
u5JQw0o3j2RyGQvQLcur2215m7ZVGBPMQNRGpW05lKoFe0GapGCdCOsBeZCmMrFp
LiuXVn5cwQrJj/W/N8U3Z5qW/MtDkmL6kyB7bSbz8VS9Ccr+rse5jvNN9HbSAPc1
u8+ZMIMslRv+aAXaQu4R6RXB3/qptC5jbxThNIBsXNf6k39RezRedATlKJDHZmpc
YP/JVneAPRSfaYd//UlPERDaqZKnSnMWzwW4Q2IvGPbtEXp+KHdOSRp3UulBVkDC
9Ii4rSpgLYdAPkBVV15WzQjdetQ1Pm0O1KudsoCIk9g/p17xisAUcnKNKdrCxR7/
snsVe0d0jnSZ5Ijpwgao06f63QpfALiKYMasWHaZvObTqiQeCODQCKHUe+K6CypN
Ou26KJm5SHkr16WyikL8R3WtgsRZNbWo2z7hLYvtWi5E//gsKs74WLcuDOdzmfAI
RH8av0xLG7uh7YgTKR/2pYPfvK/z4xKry2hcyd92qPOrXi2fhjUHupfPcDZ7izRM
mnOqylB6JUsaIlzJefasEixz5MM+MLoLStJBmtcHDTjBV1sf9/NA1m2G4kbV2BtF
Te+lto27vbJ79CY55J5RQWTTdN9RaTA0jUQNB2ok/EjRwOe2hT2XZY4ZzL8SIgJS
dsOmu4Fd9sBQg3ZLi55kTNtiJ5mlc5oYEvnk5GhN7Mq1yLCUxhBKusagiK2/Lrvq
4YyQWx2ZRQm0yTx2M4vBhzZNYHkxJ906ZdZBEP1tF+kuKFiG5mgMm0WUZRNaOgTs
9qY2EHXUGn3lbBXap8q5WqXasdRtoktWW1WfQE88OtaJN6NJx5GND1qZXmTbncRi
hRejVW+A269g3op6iuIxNDjz5se0+z5p8NdLLsy1z5HUP7McSzviFV/Z/obNFuE/
KZrQ9HJBdnvhHiRSKr8VN2rc28uZXQO5wh4mnfYEAr0mdyGB8T6DJ47NiErEy/xK
PsS4oYEAJLnQMjyjKywPKPNMAOm5DtE+fgtUczfOFviKK5JVfZeX7A3R+uuNzxQr
uhaHDPrYXpv11LkkUHP5H39J7qBW0t+m85y5MQQy0k+DTZZKyBAV5OiKlL44HRlr
004iwNM8nfAmRfROlhcL8bZUuIFWwkB43zOeT0j8bO2RTr5RfppgUgcWcuCmhZaH
eN6GTEgkFut9VkJG3nUicwgTE5Hveg0HFX7T+O91iMbrbUvQg08QORhBrsOLiovn
zXF9u1dI/lVMybkEQPfEY54nUMYOxUdBfU69i5Q44P7lyF8xki+ZjAdFhCvTWmYw
/m93I3nWPf+U8maw4Y4BlxRhOdlIuCm9Q2Zn41ew+D7OOLp21FONBDCPGzfeH0ds
st3gMHr1YDw1TXWBEdZ9t8p2err1C6d2PrQt/+jJ33cO7Xh6B8E/Hi0MoErU3I+h
/iUYiIR/aZhXML868tgACuulvuaIRlfFbZ6IkefjNiNxj6R/2MBR2x7LfjSzd2mV
uIN03Ew6EDeSqMn0wYPSJoFrIrTiI69EzETVVQgTDu9HzsUnPwVxqcmCC7bhWnkn
7uTq9ZyA2ZJNTJ1zcDEtFTPj5gG6j3r4iPbV7Z4XzskrF290C28G07aktnes+w36
0der4MLIEw1ROhmsnIwJIR92Vb3fjOCmmsuxQEHoG+WQUU1S1wa5MOkuK1ddcDq4
VBb22sw4vgacEa/ARjMD6YAJYJr36M/mIM68N5uocYCFPn5+ySU8wvTvmOGehcrI
9aML2xoJ22pJSoEu9+rvE7EC+st453RN0vlw/XzFTuenmJryFdQv9sHl+GNTBJxN
iM8TMqJ9+O+m8pCMWqTVJ4poXyWqT7s1dB+/hCyrjDUhXcxxsNMWS8iVeirsevmJ
mkk2WgmdDIMYjhJ/5ofssF5XimnIyJVDJhTSJeE2MLm+WeTKWECcMWNDGvVeo/Tt
wsnN3609ilzXCQ4/RLKegN3vM+01hNu34S0LkccRICwmuBcgeltlMCn3rnCI3QcM
C2DxKhocX8iZWraHLyaukVUPAV3Xp+lO7Kj/dDaeiBYbVPyQCiY55bdKt161cNRa
xjpu3e4WbQyInxIdudI0VjsE5EW17iDbxHnhGV+FuQNyAhPDionZivpPg5ZJqA/P
+FnSNsWUGVAr412/aMfRmMRXxEqXirhUBu+mPwBko5wgJXyvPwZJgJcENxCls0P+
nAhu9hpdIbNgGbxBrZDZgkRL/FZkikAHNTwM4tkr3hd8JbE7CbuWBobHAmTdnrrZ
z2aZ8MC0A7REAP1R/SolMNmGJhxnCiacRakTDuiVgIwr8OIp+f+d92kHFURPks6I
gQfJelpjR6fBMYL+WNtCH19E/+x/3UZgcnHh5sHwa5xF/5iN4rN26qFXQzDF6AIl
RA/9ypB7/AAhoGd86A6nVd/1rSkIj4RulOyoh9Jwdd0H6SHSC6WoLKuIU1IGFky9
Mjq0F/g7vUJh8U8VmabbWidvnifOaoTY0HrT6zojwO2ZKslFL819E77vZBL2q/YI
+9ZwSbWXW2ihJHdd0rXXHnfzUkHyBbvtsJU2TPFkMACR8rVWeUwkVhAudEWMXD0P
YiN9zRK2sOqpPK32dvcvG86c9JLNZ+Ive6oq3V0Id12KIfZiC9weEl6+AFiXXyGU
4EXAOhFwjX+82EpA77G3+gveWtwe0lLV/bS4vRvaGashyiavzgrDbNwDA6P3IB/F
z8gtHorqHC3jwEFFYTo+gBxR5V7Hje8hsjnShIX+nJAeQQYyi1GxOLJgGi8AU17G
/jZ+d0hb+OhRpSxTASa1WHS32Qx5iWdDL6OH51gcJkijMRmbetPLP1Iws0Xck47I
Ep8Ya79jGeu1gtpUYaaSsA+FkhywioeUN2K6bu7Spq95OzZSGdBDTg2QrXqdG/ZM
2CuRmHWP57r9kWKFU6n1wIzL5414l+pF34FMjmUTJSTN6en/2I8GTBziIpr2XsX1
ZEmqc2F9fLFnwHrQY46z8HjnLGsm7DgYYYgoqqPlJMp9HY7KrMrgvBwXyAgTwUDM
qDsqu6N7Bq+THVG99mEx3bbWIaOs30tE5lhHP++fcqmOjZQGzb2gO6btE2u3QUro
/26j3Ek7wj79uN846ifgVY7mKuVDmYwERlqSUSlljq22jMmUHVZsmpcydmRteBzd
jIIERgosVmZfP9XF/qFVAUazdJ3TJ0LS3h10oCivDXdlXyR8WzQMp56BROO1PZvz
7mt5gBK5Uzp16jRZfdPkwVvA0pHzg1KdzAgRHiLjw6QIWrE1jj2VXzGJ4HbQCxsw
sCen7+uzqPiMzyx/QrZOVC/odYyWlm3F8bviBaWiLDqKCclwQV6LqGUXjuL4sJiU
TzBHyjQhI6C9r5/vVm1fcnJid8FXLHFo1Azn6u5ORUHPjgyzBCWp15OFESpoJrDk
nr7nhc0EiQx+47+t/3UHjnsQVRbNX1OUeaGVTtb+KVjA7iwfPkxCZ8MhDvtcmCR1
vyXXONiOMr428iABHEmAiR30m0/ddBjxhIAiNINPMVEULgbvpeEVtEMcszUkw689
w0uZO1oMij8N947qnaUiSZHu/ECZiwTd6txLJhXAI/95z4oPTbEEGFvCt8KzBakN
+SuWbH7krHAycta8bK59UXR3aC6LLpHbfBs6x/lspMqtptMvXoFboCOo7H7+SY0q
ePEOIM8wyzzLMxV4gdDuGB121k6DlunCe13gN1LuQ7vGmtxD45Ld2QcvEoU7vbo3
06sumpXNGP/QBMnOUSl6z2HVopKRBeikdGQPfsBZtvdF/3fQyaB6+B578cTIv+jr
CBVv5u/oed3yGwkZGwMc6OiDKhNqYVsf5vRBahmmYw5ikT2AISZh+cvZvW69VukI
CofA0hCUHIbsok1A1BKB8ZuAKC1zA5OhoPfY22C/j6oY+GKcn5VU3iQv5QI4fSnF
RwTTYGAkY+Qoq3XkmNzpZ9CjHpx9tqkPZ2j9nWJpmCTfWosyoQR7cUEvNcm+1mlA
HiTGiuwL/FeQIB4XfR8tX7c/WUKGPDDZOvo+hz4oFVJbye06CYSC7ZdwpzM/2z6D
wzjLeJb8yCWkY5ZxjiczK0kmZk51W7GoY2TDTBwtVNZI1dIgkE666tN0BRL99v00
qcIswdWBgDg+TfxfGQE5+9ighJC9qSi2SRYIK/NxMPe36T+G8DCb+GWtUpR/caVQ
OOwTtVZnP/3k9gtRwoHwizE4bQ4OWAGJfRTt+mB6ES8fo+cyh3Xm2ua6KzMwvdT0
ZEINtyswgn453k/JbfSC7bl4p9/QgYwmT9xw3eutM2tMqbmfPB3QV1uX+K6oj4vh
F1UNPKb5TF4bJcm2aGPUr5dM0qOn9z8Ugrh+mwGlzNV2KAQF8jgedWtEhecVjaT/
wvOurrlTe/hkQPBp1Sjg9TBRTLksS27NKPaM3JGLyi9PktVdFYHV6IAS7G7ZhZ1X
X2xQauE0kcSauixoJecSmTRnDJqbwxmA7g3H6dbgla+tol93lJZ+IV26rjNT2wu5
tJCB0y56ouZINAWuPWi8FqdmDNbEGimXx57SO4wfxZF3MZyQj/4EvSevzg+5lq1u
6NJ+WssqSC71z16eLkXCSC7itS/5xb3bx3dxVGyihVX7ldWLD+9yYCrYO98B2WDc
IjX/UwOrVIPeihJfFGERAVkI7EPbFhUOyLPUM+JaIFSI6l5RzlMfEHLS+G1DaTga
Ryvir1GRPw7hSnGDPcB55IQnRrl73Wk3i1yVcq3IJBcpoLNzSV7XqNYOIyVFe0bH
oThHKktm6AOBChcOE/ADRQjgtTok2ukczvnl4UfQXPShIvAw1HtIqzVkHW7xhN6s
pZ52E/sBV9kFinXesiWdl8Z4f8mmNHECp9RqCyz/uK6sE14ZpehywB9aQP43wpP6
MyfgstiF8n5D3c/n/p7gzWQjSbCr/xlTpjKZtYn7nZAPj9xVjb298o2kQGRTXkUL
u4p7lowBMhVKo7Z04j6nXvGCkWeraDjzK5cUqxe0p6OBC3gvC1uLTsEzTI27GwZ3
OTh0NE0DvC6JcjqK2O0rbpZHvGmdEPqvWOZn7PzP+adbL5XLNqGpmZM/eu0d+A0l
s9EzHqrQYE+zNRs+4KF4kmknD1XaTEbJcFotX9dJiiIYRSIyJITI2c1fwHf6HbbN
Od+bNq8FiOV39wEJKrupqlDFCA+pAiaGkX0bhh6/yCIXKHtwCqQikUhQ6IOKY7I2
RrZJKlYOp5aA09CwvL1ZfvW2fRa7/SK4Qki4Pd9/nnqxv42VKBEFTEj67vq8lL+/
/CqWKVXbBsrJhHPhJEKHu3m3MLN10fvIF+RgnUpYN2Zqmy7u4PzATT3+PmOLB7Gf
5J6CBWg8FMlM3mtb/KDa5d1JbsTyLKYp3aQxHyuElV4LAyRMl0yDsAGncMesgS1o
AjuD8KAWcGvl3MDT2t5SjyBsj8xZxcTpBbGhiNH9iWh9H5M7+2OL+MO8wYtIcE4U
jhz7G3lQxIeSYmPARMAidNHgsTepGm22voFYTcW0dzzypCy/IaEtXndtf/JC80d6
Aq6iqhKCZ82KGg1HikiTtG/9tAFzhgvy4YMnf0PamS4T5MBtMEqf3fe0CFozj6MG
qPQjCmN48t+OvQfeKxc3ZR1AG1lk41VNHCekIj+UDgYkhuMO5HcnaXYfeXDjMdv3
d8yYeaHHuM0/SD+JSBjm+zLkab6wYEVbHS3xTbV4BinYNLIwLyH1loy0fkRG+XYk
Qo/gMQCE+zh1Z2fnaeOCus5ZC8l2tXYf6Kja5AcHSqTNj1rSD5Dlhr95QHU/bmF+
5JNny9zhGdYGL5qAY1EhMbnjUKskAx/M+6W1sYg7rwBJswNUYHer0xd3H0gopzcg
3B+IpeYLbVOMPFJO+SO9DphPJAlHfSCeXWKaOCYOV+rrD1R/LhNqB40/0VDwjhiD
QmxjH0GCR6kT/ouRsTS9o3Hl1SokMJDPDr4FgnepyeAkUOjYp7OlmSK1mrKQJwO1
e0jX6rgGKbaqMapRDDNVsu6fxQyi8AgZQELmBFz6xNp5iVFRuEC71mJ63C8baGpy
/iHNjxiRdjSgU5pRXlpUNfzHPvJjBBK6WKXqs6Mt7I4+WIExgPUGXN7473GHGGg4
LEndUYjDyvvhBXtmXV3n0SmCdBQc+xGRuQdJ86PQg1y4xKmlfEK+COR82afM130v
Sj2tuJqYyfu4LVrw+ub4YLRUEob9fKSobCPtTRmiJRXLBwKdDx4y4Aa3Cr2BrKVF
W7NYOFLu9rNxl+p/1XI5zppZP4+zfHRKB7Ug6IxXhNEE6LFUo5ZhCJJFznU+6B/Q
hQ2zaafVaYcecUCXB8hMLl7QmR5pRjP8dWuxyLFqYSyorzVz6uQWNM2meXXTEroL
Ew9Srn4N0Zf+apewXDB8MlYO9LomPwFOA/sDDGjR5C1mZbtBe2/vgZxJRtV1JZu0
XJ43/r6oqnyqewMXqxg2j4tNc24zw9wz5+lGfxksZZMtMyjT5klM2U+edGP5YbdZ
h61eYZX+YGPpowQPLyKqAztTlc4nX1Kj6sVeLUNYcbF8v6q4AHxlLtuTfM/5uAyr
/GpvG3zdY+wKQFWFwyhB8eZtDhneRBfr/Gl62baBvIkxXbc12piG4VIGJEWd4YcS
Tc3bcwddjqJw0512NDBsg2y7CH94xgsSo+7peruqWSMYePBdvfTIKXSAF8Xrk1bz
raV5jPrCNK1a/OnNMkLJfgLferRQakBjx1bs63/a4fXmbjKwkHCHMiKZBWowp5xa
0thzAJPTJQc+ZfUJHl2/sSrtWuDcNHCcA5SYYneSIGyBduIOwiZa4ywvtISYTuCm
3Pj5rjl8tWZ+Nlnwvzg0VeqVt23ednNv5ZgmRlhtSmTiYRC5jEV6kRl0MdrWfVAA
vmh7nU1hBSBiMwPBiAlsMUr4lb7K81L0BBbwtC3WDqmHawffC3yMD5qp+P1cslML
fQAx8ZVeWgn/+C/yesBUrQqcty5o019dQI16YncnTfUwWqVmWjXTGjHwXMK5GEG6
LxmV1bcwXlVvl/juzk8eEGAGkQWUF+ZjPWO5xIj9kY//Mf1H6uOJpKb0OrcNzheD
fegl033D19/a8xV+O8GP+rvv4t9LpeF6JYgZfaNoeexZS3F51e5bXvPnoflAVCln
UoEk+QNt5ucKR5TrVy5Wu5yNskiEsQx7TyJA7CUmdzdfoUjrhGexF9Ph5ISSeYqW
X7ag4EK7NlGcWBInZsoKKIugpSr7cgdrebyiVExUWEd67Fj+bTSRWaMHakcMWChM
8Ma7zk7hNrqGaqE+Juk/JA4/vcdFL5CMrtPboV4ypWI6I+7n0kxALvlcS4D8K9Oi
/Ac7GHBxqoimQq8uyMGkr9jwiBmFPyFQent7rTTbxlHY21p9lvdY6qiV72r+Q/iM
JQI2wfF/JKPxCUbmfSam1h56p/IPow20+8lFjfW5wSUwNqGk8JjAMbXa0Vmuknfc
M2784jPxezs0C1XrZK/dUpRyV2uKnbG2ZG4DeTMI18pSOQiezvQ/lU91hUoF6Tvj
akEniD8vPTMIe4s9gK2pZK7QTlslZTmSiE63XT0chF/NuCIgZJ4fXpksV2eulk9d
aBfgy2Zi0nCE4Tbq9AWE3gAmyVVIK3QCY+UfrkfDX4Ljj1eXISETHwKaeP7s2d77
rS+rwH7sxqYU5I5vxuAfuucd/dBGKnnkrLjTQ7iSt2pleCx68lQ/kZBjZYWHjdA3
RVvaHMfhHUQzTLa1L23BMgbo+zlhJui3PUVj0+xnTznHhGi8f1+K3mmNpkPQSb9K
YDWLg8h70DSgpv89Fz1ZmBUg8l2O905Mdoh0EPZ/WW5H/J2pNPsIgV2GFTk/yH0o
uT+QmMSqwid0+HHK9E3da3IQIQ5tBT0QqZFd4shjpT/j/SFDwQWhH/6P6bXK2yxm
UEtOVtWceE9xRdX58iZBYzGr5bjZWJAP2cFCCR0yqYuL8+pJPpzLgfAn4UmPmyOb
WvGOolrq9fiGThvYqjSAefFChoQNTv4LGzL3Kx7JlmqB1q3+TB7BhONbUIScmwPt
5H0hZwS/6yT4HEdvxNMINjBk/NCET02OqpaYrBhC2whBm+nZftUGa4f3x+jiTB6d
y1k8lpebRhGzO81Fj57cuLRHZEDYFQ9ZhGUP26NJe+x9IjDpjH29u/3NT5Cig4dA
Y6YVBK2VpoCPTorhCYqdhaSgEZFBST5AxDy3vU1jwBf4JLdYq6tqVa+bJi3enhPk
Q3xhs3RXikhTfZr1mOT9ZLct1zuky0ie9TUJ9JFb431UFQ2eaTadMuoARZg8j7NS
KuvYzRsndNOUKL35vNCAMGwC1Bw9LKQDUMKFWxcLitrV2a3457KSDNQB33JtdP4r
Hg7cV5ymDjYcOfhzSvpGGS1AF3scYIOlU6ttpLdjKWuO6+CVYar1fZj8LonSzYFK
WmzOR/11iYvESOXZ8HkEhBtm6jZbyY0JxBHxsacGH2qJliYGYB0c2r4Kv9bJOaKo
+GTgXuzBA7wIcG5yypiVeEdusat4Vg7gzXwh+u87rTjDjtlGvGVMotp6r/2bdypK
qhTLfTAQ+8P1VilRv1Si14osRrlAfal7wumALgal2xU/cRnitGJExP0XrKO30bOS
q2Z4tItmRONMRncyRGLxFeB75SBikssZIdoCNiB5DZ46u8evekxP5WI/MuW8XvV4
BE8jpsc/yJWIbaC8tHrsQfd4qnSq8W8r4T6pQ4l8hA7deRLx2icP8kOMGSCQzStM
PrBN/pWMm3OgKKFSJDNKJWqZUvZ+zxiIx3OlVYyvIdFVLba//SpLlgPzlbPwmWJg
mHvdYIEHPfEgEHR0qaxEKkKj545P7epHLqWdzkLzo4gfNQbDrE7bi4xaGwR4Tme1
Vm6w7+4cRQNbTpkhlBVNVOIbFUC/MuhpCskGATAqKWSNX40ZWEdS06zGuWFmCOoh
lfA46EYj76XvOjofLNETmz4GCeiFgjetWig7+PGN3M9IbNNcjMX5ivMqQZR8aVC5
rHoTXVHRv7L3mxhVEUYJFZTYDuwwZYRkfE5nPxJIrUUVdt2LUyJWuGd5Gz1BNfwP
ViRs78XX/oKn2txg9TcFRbASSh1eJ6Yy0OikeUDMYSdad8xK5QExk4OjRLx2JCtI
SjA/jQ8yVLk5M0aTCMvM9ImELvrteh8zldN2Rp+EDU2zWX2H3aYyZj6EfQo5OV2q
RUv3G5xsuOb8DFyQGshR8qH9TxP1YcuHjbs+h7puD3eBKOl0ncHg6d6mZraH9yjk
nh5mhISZrk1g4SuBDzCzKI1hNrhtyD4E1Ke9aVng9lyxDH/UkiNbkaiOydW/xnFX
FLkpFKHiB2qE2br3lj0nVqfv8jm9h6RW6BWPTKPh+uQnBs7GmrxgtGNmkX2uuxiw
jcoZY+IDsng5R0WaCgnTCYAglcI6whbJfpq8MCibFqH9xsu7jCIOouLhBa0XpkeM
xDyQCrw24kcLuoxGHwytf/22Lk/loQLC8Jos/1Ka7p6D8KdsC4G2Y8+anWJRwznW
0QhwwQR/xeBfCEXnnfL8Piu62qFSd6Mn6v3ISLh8yB9ao3cfsjiWzdD4bUH8s5J6
pK207fbxMtY7n6SWes2iYc0v4EoLLe2YnlvTCbOs1RpfhzoJfbxr0rp7BmfGrad3
r7YSotZ4y7Ne3oO/SlNZtlL8YL7TDpaZQhNjbwfhOTBjslvBWtlBsv3NV4K427QZ
M63fdqbid+goYjB/I8rZ9V0i2YPi75GGW7rSX69yu2SOla6Buh0h9vYcmPIDyfKw
aHd2WE9x5SGCuK6/ij4gtJl/BKJWZAqBu9kNoueTIrXOVa7KnUjm9Uoh5pTCrixR
tDBA8WgbMFU1fnxS51yi0g0sT2JNdwWzVhA0+zn/Q03MjSOGRBFUNeqfdQA7sGNT
4P540E/J5H9X6Sm2E/iDWugvGEcjo0ohQg715PbaH3WSx0sjzCPoyoo5lMVdOTM9
1FQwUSyuoU0vfr8aJ1k/Njxzv9/Eh5Fy7I5MLJCqH5ejFRRRCMPUl18bUO4qaPGm
aw3/03ldHVZWSb7UkKkNGTNdv5+XYgC7t3eizBBWYSWyh37+C4bUAuYD/ih3eJIk
ttSIe5wEuOzNTpVonVffI8uxCgggXMvLVofAo7Qi0YzAfF/rr+ILqyczduCCcJyS
0JEv60rfqoJx2Sb635CmCBJHhhpSzU0ApnFsgNC6DIxo9JEv49hjPO2VZr9FfI0T
1Y6JtySdu5xjEhuM5mdnSMq7yOYdRtbovEZFzpE0EusP2YbdrWZLCFrC/JAfplVe
qIr1vVmLykO20xVNg7Hk25HqsC2NwweZPR2UHF1+XM27bkncPrxJbHiIa4i5vZ//
1Q1hoNIhDPzK8Dmc45bsSHSq0/rz7fP2vGTbf077oPQQH0ubj1aaKvzwQa4L7ZjN
wDIurnDllOJKYME/ZzCwmvnrIZcjy69vGrVaHjXF1a/kfp7VDHB0rYeHSlSO1Afx
SH5d/HiNSldeOmPsGf9cRQ/i/gJeOeLitp/2GLAZ2IH97zRQZesCrxHzy6SQBdg+
J4MFfek74gbIH5a1BdVsYRIqTZM4bNgzJTX3GWFHyNm36YO5z4AtV+nquDpun6Mo
M3LmWJikD2BxzlGXOS9BQCA0ImhXrz1OSSWHEwAapONCuPJ6zZLmJ9SU6yZgdcMG
Pr0DKF9DLugQVtJl0z6Y9N/WVGM3Q8FQKMf2Jo9MZNtes2RN9MLRUH+KJY8DZaR8
89xoBFDANqIgeQS9jr5ejC3mKJmHY5Dd3kBHHq94uZS6t8Dmrog2lMsUpQdDxaCB
UqqROFEao8L0BYJxrXzWGrm8yS2AEJg/hd+QTpUSWUjVojK3KZNeq10FGMBRbZFK
wWtfscBoBtFg+dYbneCFc6VZBWI91tiLr8Wa6QMU5HMEjYEmcpjQ23A2pHQC3Z/L
y2r2wGzo5SIfyGQ/hszsYSMdTH7Heoax73OG3GVSLF7kydeiOdZl1GNO65JVyWfh
zFUC7obOiLECpafLx7t1wqd8gk4YgH2l8q86Lhph9iBCA/hcmRmSQ8Re5136rUy5
p6OF7r/SY053XbaMoJeHBJh3lkMITzSy1dVMXLiIgQG5o7QvKkyv9ma5d12dPI2f
vx+z0yapJJv6n5ANpwQgcuQdcK5MO/xWi6xhejJjXSvGe89CxpicUuShkxy7br/W
7NFbVYVF9ftr2G8rS9OhdMoL8dU0CdrYISpKHUlUSajn7TyeKEE8Vb8f4402ohHK
TL4NiMO0f0HCl4TTv5s4+fEgOmaIShQiF3jZxjgLwRecFFvG7Tvml4pN4dmgjANQ
HCpaMXqT3xHrhXsXPODhO9Tm8xJTQxQ9VR+3AxQfqj+SxSufPUU6fGDHkBffgUcJ
aHJi1hxPPfuOnOF6UNhreJcjJf24U8gEREMCqZbzJZi91M7ndCgfK8LkPxEvQrWz
bq5SqAQ1Dk4z6ZarDMo6lytcFdRuJ6Ne05I3SHYG8tp7WVxBYI2cgKAN6Y0h767x
iBvoBbfCUaLxBKjYKaWl8S71b8DLZbLvaPrOzCz9L9L91XOyC1E5w270nYkFO1+F
jIA76MNSutMMvNDeSZeyZE+JMwjB9J5RVj32Z8IwofYm9A7aE/X3UwePK17Nj7LY
q7nMHAnr8u+0V12M16pLXf6jUz8d1Mw6gc4ZE6mCGpZyADIomP9RUUWgXGtaYrJ8
QzIsJKLFBJmlb3iQezKxSI0h+fkmjNrSud7GA1vdX0pgNaGuYyed44mNhsIJp0VC
6BpWmJ64z7Bgz8Et2+ScCg4Rb0REZhXUdKA8iZpXKN915kxhtZI7rwt2mfeDgh9f
5QLAcgh67huXDOuo/hGGpNapArIc8adm5KV+CaTxltU5/kTNr/G7FC+02mH66qOv
iGS+ZEQgwFwg9+Ex8/p84EJ9ULUL7tSmT2JXNO0UgU6eNjeajijnFA5YCoE8Nmkd
bj1jnuIbVsek4VkcazjNrv7mkRq2cD1OSlYpN29RVOm7KYr3aLCsMI/XbMxUuyQx
j/G7E5xRKxbTrPYLtj/+4zFVVtd74k1y8XaouHcfalxQHq4yhL0wDIax7FYdiODf
ypEXdqVoaajGRd+TuPHndQSwLHDeYD1ZG1/xo18JLbibcK2YfrViwFsRsqSgwlSi
QPsUcrWheT/IAHn/AZDL8UQqb1jKcEQYoyWZVu1GBemES0pEbaHrNDWstXdLYQMd
Ahc/QalFQCD23Ffi+N2PLGR4+VeupQ0w9Yp+kPELiJZ0mNMXMtp3Asxm/nT4lS4l
jcokd5KoSrUcaW3uvjdkSyzxZjB1nrX+adU/j+u5noATzfxYtDrXj/seaoHFeCeb
vl/lK0z2BSf2Ahj9Vwact3n54f/SZPds8zux88LOhy5tmqDHC6ZQ2UZ3EZNIzTAP
lnksxPHPDkroaE0RGhdmmMFFu2nCDumK+5xy16R5uCNjg4lYHDFJwrlTZtnk+XXm
oC2EnxMDZ8abAH59DbTOukkEVFYDJH8ClPcHdDu2zdI7po1H2dVAOgCw/BRJbmO9
9r65nko5ssUwni6U/ndQayapDoOg3ueDkGo2jhDZtzpDCrRdpdd1939VS+5O5hrx
8aenYswQ/9jBKMnaeYGmgre9qI5MFfKzujbzGHrbfykB1Zkw6SDnWXA2FqH6EgKI
1mbgdMU8zqHnrJuvmuJiZeQs+KkiB5/OI5AcJiqqQTyP+IBZg6xqwrOw+ZL7yVzo
QQLQLoS5QZ8mICu0jEOFizucwrGeTVde9TG15Bhem/4f3T4/B711+3AXTCj68CHr
VglUzyedTrOk3uAvoBctcwDVfF87pESkNXBVwnfj9nnI06kJVtGW5VtAVDeZMbZX
E7STb33gER1wqWJ+UFop/+bBPdUWt9I9D6mQwGB7xnZ1T+JcNXyUgBhZSbWJYFiq
xtlN1aYCeLF7/aIyaqUey7nElA0ZfeW8BWZOHT5A/Engra2mBQKGyEWG1sY24amY
gsKVpbm7YlM8kImiLuF1d/VT9eIKXcWSc79iRf0tOdeeFAlQCWnf8IEIOJz/i/qd
ULGxBaZktwQttyO6GoV+9aqXVodEGpbRCmPG7RK46zP2y7pU1NyHpCP76F4xZH0I
pORydp0P4NPo0PYKfFznw1ph4rFeLNAeDS0rA1Iy75+m3MZjtJJm970DoNLrUmbM
uYJnISVK79gyq3fx6GMuXFzFudD5Na0SYFATaDOfE+48JH0kosaU1cUiV0XOV36T
2ce5cmFZl44OkjXXxq004HOO4i6dlQphK/1EkRb6rGGbsxg3dEMMaUJwo8j5dTgY
ueouHn0H/XPyjiXqalK/pOdIZjAS8YpygrHIlzLbGDJIswVXvyFIQafJYr4Ojj3r
rg8NO95hl7rFn3Be2L5x6Wf8TJ4KkTG7rR6KgtyAaBnE2av6acLR2CY2OhxJd6Tt
NeL+TsjN327QqfLaoW2YgUajvjME4rztlxIbkt6NZwGbzkBfxiI4k0eTZ3uBSHBJ
A3Iba69DMNjLvCf2nYW9bziEo5wxtNVMOFlk1VScwmP4N4R2ZvWRY7T3GVD2dhMx
PW34adyuiMfTcnJn02bXCU9PVBfR2LreVsig2rmoqZnZU772MkeiPajBl/Hjisfa
MsKoX6nnC+nRofCzSh/4eK6iFD1m999Hqob2pWGfEm0ufO2inPN00F5CSgmEPtHo
dKwAJ4p6BsipyXOGRgHQRdEMKKuChtudvwk5dC1BnZ8i4g5l3QDLZk0ZfF/ZTksK
xZBMg7HkwUwW+62wSSOJWJBoWPJksrvoev8QW3tfanEzF9Tr76HIpodt9byaYz+z
Smn7VR8lJ+3t58CYb7n4qX5fKvXj1Sv/ol6cnTJCjJPaunXbthIfLuuoOXBYbknq
MA9+oGUrpG4Eplep78WCFMHMp0LTQenRHjHFwztfeWIl3AXItRul8GaGS5XXYR1L
rKfKvUv6s24/uB+fBm0tTDns+nG6kETSGX/KiyfRaqH9bSeI3yVtoia76XkRWRPN
We7N5NDMTkOCesGpVE+rNoRByQ9wuRMRl7MYtwoIrFC2+LfMyn7hmon4EFzuZ92h
XSq8GWwYe5Rqd4dhsmZPoImhn2THR6xAO1cwjI5bpYkGqs5gTXWpTJ92N2Byk5TW
SkEI2xoHuJgnJNMNUeL0YuIDsRJ9FXY7skXgXtemtelLpEOpn6b9rYoVNfQuV10x
gNPXwsfWcVzv5vaioFKkg5/Wz5TcJniG0S5AcRCZjrOj9ipmkvEPZalxFYvw4SwD
owTCjsjqK3oGAMa0MNu8XHj6EvxNHpp3rZhwyGPt8wYSHNBwlvhCvYHdNIdmJAiD
aRM3nGKx4NJjcyEg7hC0SwdAX1AtsEX3fjevKb1vaP9XZi2A1+rnes52yrSANaYA
KPGlKlVcqxU5DdSc4f0OD70Z6SDkMEZdNn27u78uOLcBm2rGApMRim7k6rwjBxMm
+v2z2DeiMAgtrHL8egRUUJczb6OHj2yUc6ojcpiITsPq1QUpJuCkPJ6EYaaTIg6e
ru/7eSSlkoRaea7dEqdIwKaY5BvsswHEOvAaqvmMRvB0tARnIE6ZYa3Bm5XNkAtz
O9Hh5DpbwG6AcHLtIu51x0EwOMHLwapwZjL4+JiUT3ClN6af9jukjy3+aHvQ/V5r
K6DW3ZQ9lkWhC5F8k0G5de15OLpP+mPhrHE65CZFk5y9zr4VDc018udaoKpaikZS
5kO+L2qr/b3+lK8AirV+SPBgfSKKE2TwIji4tXMHWbX/jelca0WnylPZ73uSS++Q
RXy9bWPHH6Fqq+nws4L10I42BLWwKHsxXGN8Gic4/FDPLwEnZvL8ILcjXpWxpdNs
l4B9Ai/84YciAbVqWIeX7HH+buhZ7gztoS2wwiOyjfKgB17xzNAXmr6dHO73Z6/d
OWwOCpsgxyMRTvtVUDcca7bpOvQjzbxUIawuC0gGElrb2h042Tg33pmOeQPfOqgy
IpS7tvJge9JQXBqLQwie1prHYxfekjnZGLEV9zL+11RQvsvEL98exuZrYBVF+3ym
vmPJXuw00f7Zooyvj9R6ldeMce2sMQgi8rbgO8ECEsLfyDH55zMDBK0Zrs3YxNQS
TblEWJ0iCn6c6iIWOYAefR53xmNDyDOf9DqcmdGm6DaYxqHorbLyocdioEn5d0zH
yDoyEQQxZYz6rkID+SPLmMwVmpy/FcBenPEEmY6MH6YoUHHb8xGEnhOjo4AGIJ4W
c9fF1l5sttwTyYmOCI0BJlXZXG3SsKi7zvT3Tc+qMYy+80XmHRgHu9voIByTz3P1
y6OBLN8+Yfwcu+T331/fGY1G9oxLItTeuv7z7ffNM6NhXqxjhskKSXa3oX/tG2A/
sMvvW3Cdlpdp8u7WKEcYKefWmZFkiwJoHYbqM+FGw8AwEVp0hIfGfL2V5EmE8rcK
J/lo8yr+hkqNvOQj4czC4VA7plB1MUfy+avgvj0bFSPzzIcOX2Xo9vGM/mxRwNMN
dKV6swzt3Ox15kItV/mHD0yFh8Xhi5MkrTi7eKL0TWte9G0BaGBHWpGHTDnGJuxW
wpsKEXS4e+pymQ9jHqc2sTKGTcTduIHGZe235Yq0jjKfgo7xCwO8ZMzyH2aVQj0e
CoIAdPlwaUjKFCmUuJeSKd6qQxTbo4YexEH0An1VdVMzDvzXwx8a0+6lCOaU/ZQr
EraZGjnuWBjSBcVsIP3RWw098lsOd28kZEPYgF8jPfWJVWq+iaymPOhWQSvQvDdH
CwuLGtv0vQWfSf3dBzMuTlvDQmXcjjg+zIeS99hTbKRR4m5KLA75p+NMljFssM5K
r089Ow3zq9yx0diH9SN5aekAQtARcjvJY/SD5GwzGY8lhoEduFucuPBR8bamd2TX
3Qga29magSY/i7oCcoNuyD/SQpXUkdwjKLRGXOMfr+9pQWucexi4LXGGmuox/RAg
iIpS9CZm1FYJWG85tXhyzemp0cUFNQM+TY03/cCZ8Iw6ZEOZDxOCMa+OGUpsONBI
5Ot6FgAGRWpAlYJkkoF/LbyZKUBpPi2Ah3qjn+mVQZlQHMCO8/xNkxfGCNMiaART
tIB3qWMgtSoGRhdm0YZWEXJBUfh20Ra5jo6Mg8poePBPY3Wkd7SyD/WnEOtEllJA
IPrMKTO5edHKOoSQ7QpGirqudLPdJ+jBVqvoARQxzLGJS/KfwM0tQQPksrsaLmHF
zcmYIO+LFtbWCOCeexdaZ0m0yVpK80BpQ/HPwKzNeCOFqWRw+y5iWZL+G95tIWAx
alUo/ak8v8GPut7CoZLPH3O9WxD4he4khH24sQk+/bA0iXVG1+N7CMKIkMc6mT4k
TKi/iThwWJbInR2wXoATp6rSigk5jf1ICeh1Cu9pfOhyu1VXKpvgSbYwNPSdhz0Q
GnIq/W3cTrhHHZqktAmFrD9peXQ4HZ/b2bu7jdXbDYbCK1PdKjhtJDWp5qhOL7j8
TAP6WXb3KxImqAvYuW2rmo7GRovoXFnZDf3viorojUceUSRlmJGkIsSja0KK7edK
ZC76M683Fncr+Q0R/PuNET7h4d2K97VjIrcn+agRuZwTBFYTBD9kzkDAYdx1qVMj
vM1MqTugNOxYVOlyf2KIPvXV3i5aD91Dy+ruutuCw9LmgYESxAzozxdKq+Ibc3x0
xoirMfhNQot2rYoAmx+HKczVAhKzj5lQNREq7r4u96TmHAQCDf3hoKVDIJVCH05G
eqx3FVRe7E7eX4ZFgx1/Z1hN9trWuoV5aazpjw1Jl30MhVqCMpb7Pb8uOA2OlohH
qB1AC+kcpcAh+viGv/EoTcZnmxMLr4/m7wzGOaqssnSHkui1q5j5XpctPxSuJtHk
2sEHmvN+xtAynj0ODUdfA8YAOyHQDzMn0YJnUk8mVrypgKcl/14uZXWBGNxDJT1w
zOljJvk4T2FaQ/IlQKMzmsrZFo+V4HfrTCsK5iR/sHmW5D0sumcm73G87WYBKR7o
iNNTR+uWNArnCDu++eCrRsyF28BbDOcAArNDo0NG+ebUKMPegjpKapnjFHa3c2/O
2n/nneBb+xI1DBPJBBDsaCiwz48g1bM61FIPNt1R6yX80EiNaLg4lRiy89pmRZu3
0BvkDPPFT/yVUqvvrtS0AlOxDDVSLtFyLLZJqrX92sAtfgxYjh7MJQWRAEO5NB6s
Mh1e48ZTy46IAu9NslQ/RcWMUL15PKUxhOxkDlROTOLgT1756uNWjd2MuhSBiDnT
/+w3Jh8r1vuSQY+HWjvJDHLTDtY9skwxj/HjAFWYEgpHQM8Ntrx6CSlFO7aGRhYZ
NcOZXHQlt7qjhcI71ivt3vmKQNV3XErwYZnO7eWvuBJ9YV53wsJHlU+mgOy2FeFW
uEvFg/JjP+Oztd53x/WSHlF9Ns1Jwv8xVHqVfLXCcfL7DbAYTgtix5FD+7uQCzMa
2grsFEQsB3tvO4usGMk+W7C6VvEs0QZ02BFHEegU2mOmrqbNHZpCe/gl435gZ2TG
4GgkMxfsChvixtHgXjWWqoKxWKDMmmyC4+LskV+SQAdeywgeBkNrDRm+JXMdjz17
yVPJxCH/r3koWb73gddH/IiIFhkAqoTl8PTP2USfkFTq7IEG0mu9clQ2hI4Viz+Y
23S44Q62AVPsElz6eC5vLwbuek10v+J2Kyy1428RweJJB7Ggk8hvkBymI+ot4FmF
azBi2AFCtE6C7wVMCq8J3oMOYuch9pEeMX6/+NNpvL2tcVjiGk9wzssyi4A5s/yn
DAU5zaWSQbFhksh5b32NkZQI2/E2anHsrJAJf+4DU1gsMtvEL/prH0PfnfDCqqJ3
x6SVNkuqA4acN0uW36A1LCBuC7Ap/x6oIWIttRMxKilJ0x0tXawdb9ff0ceXdX3D
fc9jdpP2YhMMGqEgaxk1N8cO7b4D2DmPcH4U7EeOprq0Ml5UXqQ/Hi869g9jsbZA
z4GtFMbqVmr+F6Xk1hLlwmhNW4gblSCVi28GwAy1G3aI2moItKB4zgVoiZvZYUGn
E5niQfIHs4p3qQ9GCGz4qV9EE5uz/NiPJM0tJi1NLJ46nwIGgeZwj0euORY6axZs
0OWC7MCXjoAxVRyI/e7DARGgUuZjq8Z75VIziOMYhaZqIVzUV+l32++nfScIyKz3
bRUkUoaFQvws33oIL/vvXUY4BV2yc2qPcQNumCEOYXTiQpZKBJyGPEz4UMDmFdFS
HNk4kIbxFrTIyXwELt0SlSCW7eL14WEl2Tr5EuqG3Y3vF8B6//Yi3C54nimaN8J8
PvgPxVOu+hZvT0vAA33QMu/GQdMmVF3WCRpMvs1lb1qzbVILTjffTHtugvly5CuW
BdrZDXeLCxzqjQaKoaQ5IO1FNWVGTnjFz5fKtrWdfdJkGLlMh+1mKfdZJfHAfkW1
WfWgKsbCK/YglcocPlJvgYvMZRUwz4QnbKA9igZzm8RVTonaMBg6qWbfkbO9ttvf
AEWjVB1/59Qr0TtZcm2NbolJwOwmBhLQt7LA4Y+gvrJ1LmkDZZDtmEsIpiTlaYUy
F4OM9z/IyENcA3pFg2h9SNHLcaF7gkCO0vwpfxBkR7ct+hhuZWRyO4eRSJMNCsjy
QJgNxqFF4l6qguqJkj/Hu52M2SFaolbWq7PebQ9FtNZ1yX7cMUWKdzd4rIhj4P0D
fzcaCs3YjAillkT5ZJ50iNhyQtoorBEOWrzqZue8Ath4NlGBFcGogr3+IreLVf3E
ANPnnxiuFq5KyR8sz0YvHGJPXD96RbJmJwEUNf09S7IbohJ8LBT10V5I9gX2nlOW
J4mE0/mGFALaq8059DYngnFviWjhkDsTFiGaSugTC2tq+MLkK8AVOPkefDW4HG6h
nvJZUMP5qOmdjVaqv6lYLeyJkLGfFGGVx7yqSWQHk0m0czGcKQhq9Grw/XMw3Cn/
fASi+uTEhXqEyxKr1N81Edyw7jRb9uBA9pJrGb0jxdFXjTldc/NJaQJDYSHJa9/L
5xifJmHnhBEOKYITJc0TZ5F4D5Tam/Of6Y+EDIlpLnZLqsV7/0B8vIjPG5+Fbwb/
FnlNTEDbV8EtkdHmsJgTK4TIxOaFhGHfAo1GrYauECgpITYWYLdbsqRev5IgSXqd
J996KN1tjjkZQYtV3z9rXHNyj14BbloRlvE1Ont7sA97QzfwBhgmQ3D+sRwU4r9X
2Ecgh1zmVdr1DvBPAbPjPuqtKAySS3473fcM+wJFUnJdYCm6J865NVMNrJQR/6qs
S+ug8kqGTAVlmHLBuIx+vd6JYMJxCuNyuuaEupzipF9+i6dbEILwV8W3bxM2E29m
YK4qyYpvkimkjcHyuk4mFJ5B3Zm4UhcW7LURAJQcb2OpBJcmX8yzEvTuzrz+sNuX
rrQNG6Mk1AEIXCdSghM/iw7/R8B2msbl1ENuOOV6dHdIbvhDrltXsN5ZsDbrZ5zn
tHTrZAEXFPD6zHmDjcf7YUacFYVHTd4yepWulDCUmtm4sym1YS1vDPXHH83+Xa8c
9R7fQIVebS8N4v99KXL4O1JEuB8NjIhR81N48RXc9PygMFO1TF+9Dndqrw8lQ06p
MXpi8Ekw8UH5+FnJPZeXOTxoYQFxbHCck39AwF65I/l526UErFUO5JR1EXRJA0R+
14WMA66PFtFt+1LS6+kk+jI8EAM+BkCcbSmMEi5Droz9845u1tUZt6RJuubevrhQ
9WKYy2edZ8vTnDtow+6R3MdEJGSiM0ZWEei6Y05LPaBRTXKdhD1qW1dTxnWZELg6
BOweTpqkdrIa2q3b6LTVJM4KOhx90z6C3tzl9r2rawoPFgintVQQevG2NsF0p84u
HInjBd7jr/X65kyEVvzPjpq9HEUYjgOuIBWZigd9ZeBCymaepuYagZmEZkdzeGEf
9VJ6P3Z8I0ylAWDgFF/ST+GcOpzVVgzl4noZKSy6faIsOzDi/fEQcsZ8W+K60ADN
uUqJtYC8hgJhDEkiK7KO8dfiCM/FfCvz5R0cZcEMxj+3MrZG25FX51LsCnqNyv+6
mhzdJ0I8mGfzivBAUvPf/3VdGJevjYASZdCy8lcORSn3K2xLDv1yg6N3oo0yMHuJ
WRgmgbUmVVDoqSsBH25dOJuvAq65N/N8LLh38Frl5OwbdikqX8TcnLpe8K9LI9c3
smarymgwbrGvHvO4zr1Wm8PZxB9LUmcWjr3nLfuzFB8V4Ug14m9KWhFhex/A5Jch
YAj2SyWLGkCaiguth1IAkeYMgFdEcrlBwJkW8SG6tszuL6u35z7kzLKqwFnVbcld
dSz37czG97TfFQkKQBqaR1gio3YFXsBU219PfdXFrZNKnE5COX6bHccibU2+h+Gu
h6Yvz1HEyC9eFauu0XQ1JiAxAvFqdOCc/trq9Bh7phe+R+8iDFr9f/q8aKcb/bbx
9XNBYuQ+o594i7P2UnNpbjdUX99IKWBP5kIDYHKwWAhI19hyKTIdvJf2Jnd89IBD
j9InlLvAYkL8eYJKBNFVUx6DSe3RQi4yld8OixCbvEkZR7t8iZlgrLg7BormFwI1
HHK0ZrFoZ4vVBSaC5cQjZoXSpomTOsPpPfWY+wxwA8ftxinmoFs7ksqB9yu/xQWX
e0VL7bQP7ivKGOTESiaOSoWFYlpfgUwgrpr+M1nYJcL/9Tr7OJmuecMnKxiqn+In
g0UWTvRS+ZSR5sa3dPLGd5men6wa6fzdxMwumitL5vFlV1SQ47iAuuZErljJ/9ZI
6SzWBVOaCrx/cxgtzaahQalyIUnmEKU+x5NZQIQck+AW7S4I5Z6dbf5yNZ9nRuQl
XoSNlMUEx6trGi8Im7m0VdWAgpvgja4vh/+Kjvh46cZXEDL5qYDhZZxvoYXSQTX0
IH5MqPXPYI8haI2bIlQlmcBmTee5cSnHDKNkA2eTVvN5dE6OrPslKVWkEbiTch6r
Wz1PskQJjbwytRfiuFdhAk9hgdhR2uGZtJxPco3P2K5C7QsFXOn3/DYf5uWeIk51
g6daUyvLO/FCJ4Mx+fBcWZTeNpCifBOUWoOwa1IU7x64fDvnF+6a/g9/eLELRq29
WIHGGlgjCVt+K7w0a9D4tQUbqK9wxc5+Ld5l5d5nNYz7RQi7dmJveSXQkqwQo5ec
7ff0qa6iq8+yyQvbeysIVDPREYJTa0GiNE2YQiBUSsU9PQwMCp631hr3Gu9imr9X
DhoOg2mZU8RCC9aAhdRoUC9LStiT0fv5jSbAPRoZsB+vPlrihPdN1toF6EnIX6iB
ln/bBLQpeiqQNPwp8guapPCWe+Z1yVu3bdwEiwcE5eDWqUTVSukcL9BuMJwxeU7U
S5py/5sH/JOeydfDGO0Jo6/89ZO+3VlwFEDpnRtSofyeo7KIxiSg267ROlxwyIh8
Na8v2eCzueqRXt6N8n5ukRbUTpmHkqVPRaOYYWsduRqpDLEi1iNgC00pTwNfFqsL
UuT7+PKoSeBvEChbr5/c5G3dgnIBZKo69hLJ+aLTXfKi2PBNcH8yQIqg9coYSN8I
JkWS8R+DSVqmX6h2jhI18HoXknwIXPeaoBDd8sylZXViPyK8kEl9j/VKPpuMmw94
aZPVwqn9dWKs6mmkMQ2Amirh2qH0/9/gefapDws3JonSODmxevCEkcVv69Tob08j
N9qRXc1+OMi6R0u4RSuu8GvdagoOIL47eAVsuOgxBDp5pddLqBCYdY5iPhnwipTY
gbgiG3KWrpfQTycuOBz7WuCr8SJOT9bj6m3YVNKRKzbskn+s5LAmueiZQ4GJq0sr
pVQt6lqW43jpdFxSdXezFHDckoTu/po/G1C7vcPYX4i3Uj6oaWT88fPk8u6LCXwp
h/H26ftd/P7OODL3suJZ84Ea3hX0O6wVIagJJRUyjnCf+iPl1gbBhPkTf0JRScAY
yGF1sEb5B1giblxZl9ieaXG8hncdMXYe4Lz8DY0QC8102MiNR6tWIPn0RkSKqxcz
C+qcKdCgTp1NyJb8N9ekUchDiCvlrsjIuByw/3TGdS7EJrzNzAuQEqO6rMKUWtO7
aS60sOUlluId4J64UCNuWF3XI0n+xW7XQKT7eiNhEVUpHpeo1JCYQdaN4CaTNCR9
nCBttK2CrWDN85rtFuM+O6JiDZ7RonGWKSb80Gf1gCtJcHIzWiHn0eXFOzR2sdyd
bE2Mxdxw1yfOnEFjk+p4t4+IssCpkipCg1oWvLgCD9zbBlAqOCjYTzu5QDK+ql4J
FZ3DZaMHHiZHB/YxtQZipTEiCP7VyNnneMIT5DhhaD470A/lNp2t7ac2+YSqsWWu
c9r3p85Xrm9IZDhy40hWwsusigzEDLOLIWERjE/wbsSRwLZDjX3YOFniZJHgXPMo
xz3BTZQKosQPDH3DRQWHEGrN/UljvQqS5dHGWKFWDbWq/CjKaWJ2oKAXF3UsN2nq
Q+8b5RgLdNmZwEG8yWTdMJ9cge3sCxXtDMatZaMNL32ogcl4neS/A8bEiW5SSvKI
IzAeiM+uPq/YqBM6IGqFn/K7iRL5zxUvXViHoiA29HbgjAt8E4D59QMDnRSAMDZ8
sy2FNkw5/Qiqyusl226t0K0n7eM5Kg8DvbsKVB61nOSbHTstaXSKvVKzodHNaXeo
VG7qcQ0CeJfI6Uch6XXV9naa+VObLhrL1jXS2cqecNFd+eUu6d8MBVtGy97mxS1d
ksbEmTi8pjubae/M/HOTbTHGSDN5gJzyL4sV1oCIe1e4IW98eeAtVEL9mIozYn2s
dRHEKY42jm0mLzHJGtpxzlNbS44+5nD4iWKdfEuZbnE5twzpECREuW+dv/AdSnBp
oCr9Z/YOa2WKDuR4yX8pDD704k75+pDgYwgnEwNDnLhVgLGZqZkl/bgBhJXzKl5W
2SsoO2qu2f9+dSH5atbDITCcUWZuQC+w2QKaI6TBF5nxZkKKAboFJ2ed7OIWDi8T
ZSXUzJ3+vHQ40oKjNVTtqu7lthX2t79BaqhlbrIrYQlG2m3+wdRLjI7+VqvHWjKL
TZuEXEuPAdaJXlsk7yzspjqNJdgEv/4aaQO0EI08wGGjeaNKrgd4NqCn5KQAvDZL
Q9K3ZuA7Hz2PtvsoV3oXMHxs0j+7tNn2zO5/sxvzU7eIQ6Yg0yAJgfo1c4ezCnHx
K3wwjEt6uy5XkarT+vjSulq+15Eoc1zMGktXVOAR9qw7AQ2Zpl7O4mAiFZqPJznm
gJIe1VZuaMOpw6bEmXuxRZ5G/751nFovrQShwXDd03nwW/Mqb8pvbHkL/pgsz6p5
JOuLVw/vpKWfwO21C/j4JM3TSA1+ddZbsNeLmTGCfozJrZyT6kbNnaX7+Lo6XG9q
uU4qbwl8heB872qMvLuED/Y8nhthewoctFT5d49MFTEu0uRgLgT4Va+xofRlLUcC
eL5ENyA28P13YfYlEWjpsHqI2/21Byh19GPHdQlB4GEATbYKlAXPF46YIuZQ4MNd
98q7o+o5TigMdEl098feVbgfOq9r8ACddD/m6MrYCkLTRSYV5WYoXAyiKeDQMOuK
bqNGP22IOHZ0tuTaANardpdEU9XadZc7Yo1JKjZtsLNbCPCVO5fEweRJOTW6n3NE
5ExA4R9guhTlklieOkpPtjgVNlfJ2VH4fFfY8VLk+eLrctTtTFtPBBItukPVuJSh
k+flxwBu+rX4BcmnuWJlexsUWZLTmELL0CA29yzRWhbAZ6cTh0n+p3HKV4H2Ebgg
5WcP0CeMx0/ofa+Eq3BLvBRQyKnHnLT1UeTDGdYWRmCE5kbbl9srOJpUIVDrJTxD
C4RG7fg/cVLtPIZpaK6rMe5WlzrHkk0iQzn3TG6swU73dyhtsDnIOXM1QZenU0xC
ObVK+b+ojLjIjkZi6SzmC93vxYHTChso2DwZ72+yHlaDc4GFkJoQb6Pa/ZXVYuAL
ZGNXx5/+o2yOhp5+z6ACYoxxy78HtgUnc/lEp8/sqYzpaghGtyh00zkWIf2TgN1h
inFrwFBhtKNHuH8yPyPTkN7v3QBjbkH5LMfdvdqcMLRFEE8jUyaaaaxnhz1cts0u
XWAIMWUb3Pi/1eDTO+8jIyplAOXoxY3eaxLiQtNwrcNAZmDqBpVBwOXW8jLx1uta
iEaTaNpffTE5jjgpIVhVJThexGFZqjsiwm39qaVdENF1GdEMzJ5EcjZVrXVgcZ1P
T87C/cp3ale6A8QG3FnspVA9462Bth2qWPwgsvznFiwy0Sn7inf50EGqz1R79Wcq
kzLEtT76V2k1Wn6yPQ1codytBe7CTC9u4h50vEScJ+JeewbDKc3xc/5Mxmx1/sOq
vB0jgRJfWY4GuNPgBLCuvbmDGpJSwGwOf8+5vir4Z19C5sS+T26aMhTjiAAVaDop
5ShPaLJCw2H8gxpEhnMuU6AG3dx0hL1XLE9Fhofr2OzuGu0OEw0pHdanboc4Fi6/
OcXVeGC7H1j9RH98JrcAy1TDHl3dh3+NNp64c6swGMYxtjFubbcLbiesy2rQG/Mn
GebI1kn6dEqujYV6TbgPBbnwW7U45ZG5eZH7RdiWka3VEz7Arp59ac5WetjyuXmB
+aFU8peBcKG3HlTn1ehFCm8PG9uf7g3EYF0UyeH7HgnZeUQqY9dyE6kJ1mHa0jqU
cQh/lG82uJU5xInXbqYIxso7S7Ysu5VRWh3V/r1pQ0Fv/WMe1/hZ2kF5YHlTqnHQ
vwnEZn0Jy0EkWBAAB+C3OM+1mc1ppfyPMMudYP4U7cdV8A3lALk6jIslWHpimcNb
/DlPjFfz6I5g8a5fLEk/0lNvlXCqyIc3A38cl8a4+zFXk3SaFJFmXvMynp8m04cm
Vj/NuQHWkl96hH3EDJSmpEOJDHIBbX5C8uOHfBjh/5+uhL1BemlsawDROEsVxVFZ
qt72QzCj+7Y5W4mL7szhwXqtFJSpU9hmZ0EIrbjqaZLoDTauvEtC74qaak7w0PWp
1FlfMJw+sg6K1XMZEY51j2ftzaiMOYkxtnhtgrKlgks8UZ8tzK6qbmc6Qkt9YbBr
cIuzhWlbC/n2YPiaAAM0tLFgvyPdsrRRTGl+dblB0W5Pbr7oxNNGPIzh+hBV2Nij
CTGQ70Nw0IjY5ND5DfaqWlKv6VjnpPcUSrb5048baYeEw/rW3k61fLPwq9f6b2Gr
R+NoloK2cOX/6wiVwEgiqCP3cGOd9a03g8GPkt21ixFil0Beng7f2UHzZZ8sGEPs
RcjqBQlkwAhSaU3oxtpbs/Byf/hGaOiUySYJ/FBOpyM6tVVDShetUdBtf8ixNs4s
PBAoF1PPPm86IsKSg7+k/nfSh4Jmj62PDy0/+/a1QJubuWN0qQqCaZAkau506M9o
mjCFECK9GzJNzBVg3xS/5CyOcJv5/grW0h7HUtHtwaSO4wfwfUboI1AuPaTCLYLI
S1K1ptJmBuA4WWvcMywYupbbj8KBdd0FlLAK0u4aKliWSzc6LqWZGnHym81trY3U
ApmLH7ZoPw6+TZe7dtEhbLWd5J5YhRCFZQWyxMgUP12dYuPomm4vPFMh0/0IDn2s
R6EGd+A6KqMk9NKWajyEPapfDxCcFbOOtqViAn+fAOqmhOPIpin7gaavTxFWhz08
Lxrw1CbIHTYIYTYdqVzGCn1TY229dlc+coJmnUCC0ulODjbJUKEwh4HQAQUDA/r8
HlNlB0JBSEyrTIcSdiFUdqTM6helM8J2Av545a15cty29qZ6lnjI7fhFtDjcPtg9
5bTzkASkXJClZGH7ZzPjoSrdsZRd29k9sGjRdWOkNrpfAys2kUW6PL9zLDctEfk4
QYDJxYwpJoNJS4EnIfW18V6FyihhCx3f1CZBH+TFDSCO0STe0qhUZ94exFF2LvJv
skAXsBBxoOn5okrExX+zC5+OSuLlWYWo+PF3JhoTYyRbxgRa1grunlktgSg16Wjn
f8NX/Xtf1iKvaWrB/dvsK1vFJT7ZBqKvg1o6IWV5kTeqIswta/bsspFUWQKa1wo7
O8JJH03cm3cvznH5KTI1JUUvME0p5hV6UP+lDhsbWL1G74dBiFL2lfNQ183UYiHr
+aOj9ykAjy8t6ohQRVX80YC4EQu5Vgatg2TVFCsp8LUHHIq6paeT1tEHKSPOUZOo
nKn3/0CL+nA/fZIupQdnJ/g/PjVV+Bwk3tRFiw9OqDpIyRVb+mJLQOYoCUVCUN1z
5Q35Y4kdFxPEclKOBcb/XDeScv2BwARHU+ObEXcYPlRzZMjgjbq76pgnERIH/C0m
QPWNTZsmG4kS/DJi+f9TQYzXvjza/oXqju91Lu0faRDcwZ3USwMkm6XSdUdrzdwT
oa+BE1tLxC/hyn+c1taxl+xy6BMFvlRI9Wq82mnY6MLcUyNS+mG2b1auuQdlVRfJ
g+lXcAEyE3gpd4Y6t91MqWVFuV1CxUN+r0fu+uuqntEl05R1VDpHMJpSYA78Rzft
pL01KuLu91zTKtL+KCFzkriSJ0a/qRruY9HVlwtGrg1qHNDtpPvrmOPrCHFYd+/I
O/TfitgQ7r6aJWNiY+QJ1pmqSfiaBlPiZS2vQHrM/qjUUOVxDNNVjexhGZZKd39f
ozm6DrmKBxd94ti+Otpb8sYx1gT0fpFJkBK+JiOT+nfzt/3cCNMtnqt8PqXMIciW
XECD3Xs6K53NQPKRWAKoJM0ssOosbDpFLi+cprIlPdj6I8Dat67HMjRhOkyG/KPi
bwDQDMLuejVM0tRHUi0HQZsGpyne0tkXEA4vHMS5iBgvQH3cZxie0F6BnIHpN72K
Qua16+N5+eZvFMM/kmWaV7SPHqZDtACYOGSr+nHbLseJJ6D04bNTZTzlXDX+nMrf
5AYiZrhM37En4O+reLgkKysfetViERyxDT+06WVYd+ztjjdu0r9b6Id4vB0gKj3r
KHZTWam+dPBM+7Z2trAJwoKnXw3E5rSByTMY92eO3MfzI2xQeIsx5vM3RLvvfyls
Vpg2uNoyaHwwZ6WEamRCa/UKewGmGa8PjXa/uhpZ1nMBLBdFyRMsKk62Rms8qHDB
wL9k7ubVDY6GdbM95D8IIoMe3tuZC2Yri0SLb6V6bqfQGcpa4PI5bC2jzLXPv0Ss
Ug19Er6gqRYvl0JncjZqoAO4k0ysK8/GPzv8YsTAvelRd4SAxbe5UL4ktUT1P7SB
K92Utf+M0BV08+4dlIAvRqAzHKaUN/X6SgsLcerJ6mfEyup6SgbbKs5GQsKAa6Jy
0qotFwvrnALjOlfZF4S09MeN4yUN4ClvSmfAZ8qD9kSq0A7VELW5VmhyQkEypqHO
dUBO1D44XI72Lq/kI3QE403kK2/ZopnfLTpij/RAdF1Yy9MJSuDeq2NQFbGXFCr/
M+oK34+9iv8gWNzdTkJlnxrBKLc9oSFuXaj15VPVRDlzpUjmQpfI2Rkuw+ERDPBv
Ta/Kfbgva50khq4k932Yu6gNQbFmGITkRRdIySYRQVgIdFWjBrBNw01LtzLidfCh
teH4ssM/3r21ViioE4QG839nCvscsaBXkkt4WaMQuVcymDW9idl6t3xOGm2G1wbs
RN+p0RMEQxYLUHc9DDGuK+OhHMFLdEqVBzMhombpRZgRvBZgzbKtUoyvyoHp/xEH
bz5qHESLN1rA7VNm+0uhe7c2YgFSy5aaXnOyTiWIpvoPRDGZYAC//5Y6qmil2SHE
o7U86ZpkJ7HSgnoj28VvMsU5LxnWmxCD+UJHueb24HCxsxyHd7mt3ubIGm3OKZEx
f2FEaHqJDekyrzd5KeNNsT6iSgpedaPpbt/tUlopRgVTLZV46oc4BDW4cRmV0OdV
xeRYUlEpS2f6r65fNbYcTDktpmeQb3UQp+jE1A06gwm8HUtiPRVtdcqLKvVvSB2v
YJk4JpUeXj5l+rrhX6fLgcT6XnAYJ1Jh+VK2opB6HdvEg5zGb0JgqB2KvYYfBpZ9
F/lcVoLGd8MGnQYBAJJfXXNbIe0KjAWFrrmctgLwWgCzQsXI2m2GksyMjl9MmvbY
x31NI/WFwwGoF9drG7SFOLXI3nJ04ERi23HJrEd4tmY0NLB/AEpaqTEqB7oawOvM
ceT+ZBNP4WyLXWlodLRsJwy5S41Sjh2CU0ZDc4nq6W5CaKnZg1LvhC3IqT2GLGi2
Rz96quv6XJUEiY+S5/J7y4PZBG41s6hdYlMul+SeobfivjJeuGl6CLZNNRVSN8dQ
EYK5LbQPoHbHcObUTxKFQcASfHqYhaiORuLat+b0ZmFVZn+NYBGqzvYV9ADjJBfo
fNbGtl04tDpEaF9KH75bNbHwmmk5+KMH0zpI6ofIkKYjL+hrTz7sbgpBn3HbwUWv
ArkdICsb0pW80e02II4G5+ya9oH2ONUGqbx5JFeY/9vYSrVg0jA6o6FBQUkQs2LS
srRNUyRnHZYEjmXU5zaVeS0z2d9n4UDLWD/Rg60yd400sQF9XaYrxwEfCld5a0sE
eYyP4D6hYmJfgJIOWWdcpTp1Wpe1OtUBJ5L3HuBisJi5hX4SjkPwovPbEbGmywyF
2SAqnUeD9wHP76tQvZ/h8Ei1z27fevwwwZgdjGCqC5oRzeuYTfwxmNjnBZc2G3Fq
GluJEfoMxeFDOrpljcu1aecv9xbTGYRdULksDomaQvRDpTy39IqHubaG3e3GuIa4
gPGF1c6swXIVKpidwc95/An2FpGTud7M3RZKyBLYSwcuMm15iWAue4/znzK3j7h5
mopssaoIYqfzaFGO+/Z5CI39eWFAlYM/2jwjqMd1R4Ea9xPpUE8WcgTfa16Sx0C5
AJ02lynKUfwMI8CDeeF+4QXdlC3oN8UXZzdHP6UlTn8X5X8SQKlhf7rB5OchW2ba
D1v7PsLaCafk+y0tPdARv2boB9T1bhwCrVUjpI2IkTfnDH1a0iyiWhRSxvfu2TK7
YKAuXY6KgYXqauiPiCRw9lsx7yOtrmw4YqMzt7u9my5JotXgixmbXaQIMk781MqU
WcvD5QgnKioOC6o3MLCnED3h5RHdBryTGJEAXk2k1SxyYGkx8Pq7YFprTRFHS0QM
M8oBq+c6QknkQ8EtCP5VAf0pKOCG8IteNJOGndHmY5Wio3d+U2UuOUEpk7Pto5U1
qnYXFHDYQkkCNNY6uPha+aneOdLi4bbHLlw8LTeHD363W+xl+4cBr3Wv+VxQUXBD
CfQlu3yrh4TsMkfHTyoYFweI3AVeh8Yk9WmutDqitRaqMA0hgi8BKQYKH/U6sYsV
NUM9KV3VCWe97yDW9YUxW/tCPA61qLxhvharZ/Xzx2HOfCM5WLB4YcJxP/miMdIB
pXtIkaWlCbjGWpkWNi0N1lyiHAJUp71atvrDSzOBmEp0Xq2Na/swalee6F/mlMGG
5glaUIiP8SmHhJhY8jR0yP99ZcGmBxYVdYLQHCkZhbA06vN2NfO+nE9Y1ULtYTrv
Ibxq6uXutovoXkM+7JsrpZBz+u1vJH/tBQnqGHoBmaEshUYAEPQEgNOQkFtA7dbm
hpSwgoKtrWfpIMSrgp4RiFaNoG0GfWkgA3tdSwiJHhxeE7maqDLS/R16gdWJItqa
fVnGKg75+CZ8RmhGAevZNrmgg7tB0SaGsxfu4ZYTx+oQFFpOL2FmDcQgDR9dvtk9
gPS5JMBWYthvhewW63MX8qKKo7jY37oRjIQB9PL6sro6RY2+La3PbhcDHGmEf6Vp
OsrGUw63lsgnPP2crRlJV9cST470mRmVGaXalFfjmwlJZY5ei4Wsf0/f1cQEvux0
8qKkZIVJVfCHD5B6s84/C3G5w5war9GgcUNwEgeW+sKzPyvjqT/zw60I+y2BY6qX
ffHrzEvp9dHqyNPImjlZo/5dqicDMGl9FOa6gAsO4G+UqgTuM8ufyXnnXgdbH2oH
BQN3cC4zP2kNsy2Y/YaaCMrKqLbmYdXQhe+G4gB6Ej7gepUHkxBITmgw3wSc2+oa
Ke+OhsnevIJ8nfuPNc9jaDeSQnOzVOHIqOFbLHRUH+RqwTGGn6W26jPsNmz9HTo6
Cco1eJX0klGm622G9kX/irOR3FUJwDjpwdcF/WHp71j9zfPD8j3m3NKX8PN46QWj
aKmxylIByvTyRl3hDbfYRL3sDwtzPcBhKZirBn89IPgzLHGOzHcvPknjh1qUEm+4
/9K4++DkdKe7k8gfNo+f8N9srNTigSQVnrHg4bLFNAcNAgRpddXR+5//VJvjwTVF
4lLl4wq8rpj8pc4O7azy2VMlnUhF1Tn2C/8tMqFmjAxoNgr2SJ0d8GsvpN5vxW8n
jonwiLeR1uFDKq+GtfykYq96y16evYMDZnznP9iie4cNToTKIhpSKdLUzkYEtwrp
RsMexUlmoKYuif5xdX9Q4R6mS/7o70AwZ6GBhozvYYSvUQ1auFxnNORLOCxsD1hR
nSrneZIsO6ICRxs1sUl6tCUaFfIMlsWgc8XaBs7uCO5McygNHvExRiE34cvloEuP
XioL4pNadIQCEq8rKp/SMyXMhUU0KWFnzIqMyifJxy0FEXj+hX3/n9BrZhOCeMYN
8O+JloWho6JNUqP6jRQVNULCV6Hegm1Y6qKxEOdJRMocGmrRDYkM+JPBCF9+fBK1
0C5jBF+3oxdgn9UILEjUYujOeB9R4gBuFFFqcMFg8wyavbf98/aH5ByOVxfGUDmx
CFcbzTc5dNvU0kwovEvimbqWLEdkGMPeDxCGb7JCQLIzwklNZq75FFGrHD8CBvAT
QhdTB4UZ4wU2UblKZPDl5JyDWYHw/RGAJYTYNyGBxSSFhjFY4UixEEiuoCfJYdMf
vHSiA+D27dzlc8XY70c6kXZurNP53E6Ebv5sr7mb3eJlVacLVxFAxhTm29o/YSjD
fOKhoFryGis7zJZLYcTv1wJXHVt7rFApDNSUY7W3mGTj2sDBGSTDB714rc2c6nOB
VL4czLDEhkbzFgf9FHK9o2X1DVgvJQpI8+qTbaC3w0cnd/rIRtwwQho56oPGVoDs
3IgzjhmmgxsmFqylBQTrDmS+laMvAC80mgXOwgUw9ephSPUi7IPvKQdjNDigCNES
9WO3FYXyB+n2Z+Nn9cWXrO0IUuorfpGm110ZqdyeEmbMVPZKdu/KnGgXU8498Br7
4gNaeTy4f1hoYxyMUfKrytGPdrpF+1gBlvwq9WLdNXkyqfv04rkixZ+qRBOLX4Ce
BvhnPHtD30ePNsjVmmyxNOGKWEylZetySNetR65XbY9FXO1tX48KdAokUbHNKMcX
OMXI5Qt6aIdRDypBOt/xoQNIhrqpTbpQfVA16VfUim+aVCUxSzWIT+WzotoQSaYq
IY8nig3fbQw+CpKyLY/bagT0kW3KVk1DunQHFzgTq5mc6VMSEr1sRSXjlVqOeZEY
290jAcUMpwUmtYxqv271iSPchTpYx19EAvATQuLUjQ4UaP327GanbzGi+88sFScj
oQ2qCoRwozu6ICxeHH+rs2cxYbAmRsUXHMx4XMri+7ZAL8kA/2RvtCSqs8aJ78lK
1fdM5BkpRzh/bTCHqJmO31KECuhDpmldvs0hyhhY2pI/1xTPudI5Z+dX6wgt1VND
/aJynRPKwgOUuhz/C89C45P6sPTGraRZnTkeS6NipasPqYSLuRCpd0iqLd9HsTYB
flTAhVE0KI8Dn0I4UTdEdFkxm3m0yr3xCctmZ4wGvpv7q0U2S/B4gry/HuXqxbt6
FtiKRO67P70cAvlexnf9T5BWHL2SBW+3RvQ/YGqVc+TQ31pu2XOaYuWPizWpDhnF
2/gMpdV6LlIyS2G4sU4fWoTs5sxx8KXcrzkD2FjVX/8rXq52m8XtuReD8zNkKXBh
pjiLRhI8sXuUhkxsKOytNd51G0Mrgt4jjlQ5a1kw9hj27+Pg6XC/j8PBs5PiCv38
TF65yhOBidP5SZmN6S+VOILT59TSwFSBJOmmD6j/ES5UV4BGNBlvH+64HbBWdwLI
e7Bv1IgEgEk7hd+EixiWUjUqrulILqn9kgRZPL4UwxOOebeLDqBNbh1i++0AxW89
JwEKfKvTwU2gpRk5CXLMn29imkkydM+upx8f3c/8RW23iuucOWaPa0uC+i9RnYXI
Wf/owJrJl8VX5SQKIk8ij7p1QRIm4Dt0Eirc70qYJQ/kkOBVJgawQfkYB3puImlz
BtdedPetnY21s2ytbdNhqEQeJGQ+rTgawoeoc6Xjt3NuD0+MjBQczo+i/Q6xD7Uz
mauL4Bq75o1d/0DXhjcA+mD0r5T3o/D1SPZnJOIr7C8StrmzbD5UT8JzeuXm9xRQ
YUvjDQJN4kgQEtDt2FQ4ax/ZBJmKvdQ6DSdvfMYE9U7ejGswO4tikQlimieSi0jz
FGPZAvjl6bdlB3dFlT1h96nCgDuSSZCycuStxwKk5DRG5ZJv8mruEutsfktjM5PY
J5gDVG1IkxNViriTLnkuo2w/MHeq5+pf7fERj5sAaF6xQo1Yl7Z6GymMdzi7ROkh
gi/w6lFYuyXJnAJb1ZPpRepNaFjwNhl4U9GKFvAnGCu6E9lZtOrjr6Pd8PGKf3Zy
bTz5edkG9wjMnJ9SNGIF9wIFiSPYWPho7PTYm3+TT8hyZ30iaYbX57+ryvit/F6K
TKnuYI84Tkb4YbAfL1XefcomnPNAqnZCIR+SqPSJ12Mm/IoqznXGGSTfjc+fBO0Z
UfV1+mlO4XHBkSY0JkwD6fxPl7PbmrnBzjf3xUvz5Uahzpb+n56dX6KF3W9KoQ7W
lQ1Mwt5W0UaoD1pfVruAI7xJ6VuAtUpXEy9X12nhkJCNO6r0P837u+5eROu9ZncF
F6CfT009HRNovw74Eye4b5r0Khj0o0xgv28iloQvq7dLXA4PdkkosYpiwD5VNL+b
uuUi4P6zAmi7KUZ/Fut1TGErisWe37VXxjrUnpljtT5guZU763I+UYCbHy+a5P/L
6qd3NZubFOkWb/LXvWPi1cPcKsT7njrc9dLxyDZVtgtEjRLsr4Ch+gcPI/Orcaux
6lSBgP6zZ02t9wX9HTfO2PkOh5wnIcSeZjjzRm5GZSyaPB3f8xRTmVTkbRVESrZ2
1hcxktsUCoWfo7SluM2+PmqiJp1NH/U6Wn74h7TtwrU0YbKm4crrtr4+/SAMyxaV
6k2bRC0Ec6SSnwXJ3YWuKzzaU1zzenaGQzRzKXtWAjFyAhv/irlzJwVlgUs0f34r
M1AMgio6Nuo+pwAAeUYjEOUslvgQ8/WjR8Ay/NZVXYUnA4kS9eB9ukArS2CeezGN
osP2vX1I++X2bs340CG7PwpMLi3/aQZzVil8+rYWjDw6QCCal4obiWq3AANX4hIs
2Z7KzohyIsAaG5Ub1UzFLHtDEe5h+bK5wL2jlKWAewLhL6CdNmhNO3LABlTzkG/q
z0qDC0qCanxJW2sRUnmqfM/eKnJAcnzXhllSK5pDv+NCg+dtY1f6U6765lPaYUev
byI1BK4JcuWKWzSI+2fKZj0veIVrMK6sq8SJJ6pSKnHpKjC2lYT5Z147ou98wZOg
HaaCpF1j6AI/csQ6GGp7wwjiqfokC1c74+LiPoB+KLEIOLJbSO6RRbz7GMgmtMwu
HNGR8gw5yHN29fThmbG8YmghFLp0CjPzcbYTgYc5KQYgHVW/L94GdN3Lof/k7hPP
BbUJYdnPQTrUSHQmGL33lCEWYnj1Ws7ns2QoaKNV0UM49YcZru/Yf1IpXk5Q1eDH
kh8jgmnZiaBQTKTYhxAGcKkt4vLKteEDvZEG9LCZovn9G97PzgY7x+64hgvvzmNL
IAaE/ppnwO756KY/dMSJzbDPKnu8hK10IVSKXkdMfRA7kWhDXDarZLQDqbiUXdx3
HMDT1nhS91IFxqfxswuH1/6RPpXjkWqHobcqyEQCHl2M+z4X+0zEf76oqfJ9JZEX
tM4ZZJMjpWxHf6XZBRuueTZ2LhF+dmPRo5GWDL/nEng3ejDkJo1IduiU6aTbmmci
Y/BAUKkY93mRFbPHV+qXdSTZIenHD2iOHuB+T2D9eexHt/LCPzDQCjQ1S4avv6pI
CZQIgxJ78kDmFxbRMeE3YZUcZtBNMMhwPwo8QfdKRSK/dBeOzLnG34zd/adsw7yD
D9Wupi4jJjsNxvKyT8G6s3yebz10gn3hzlRB9hWQshlR12HW8mmLvJsIOtYrEb/W
yneb5fnUo9nsJ9LG0RyEt3lbtVpJPxSZH2fUp7V0WecZuIeWvCEUm6aNIev/+7+a
5AnW6bkHpqSP8MW0r7S/go3IKrYud+I9sJowtpNsFqNtRSOtCgm04ziRfOznGdNN
ExoKnSoPizhNctujkGnovLkh/+r8m9EESj0xzkDmAytnWmzDV7JR/kCPkuQJZgeq
UCy553iqAeiFK/dYwDvD22sKK0Zq2IIq8cWAW3UJOxAALqlDVqH8ifkPNC6e1ikn
gK/Ew66rmttGiGDZXpsCxvp+hoYgiB9O+2zGMnIgBrHmCpjDNg0lbqLuf4i1m8J+
KZad42sRILDtPAjOABuH48mUWe2/XpA6nto0qwdaLhPFBajNXrM0XUSoG+IF0DZq
apYycJ1DfVBlow6qVnPkSVrWtWCTx5coyzUiUqKsbGS3v/2EZ6c55zcQ50Am2NVq
mxiDAqtO+R13+Au3bUwPKk1srKkY/2khQRL8E5Kl5ZYTcq7skxEIhd1U7OgASbtN
+l87yWX9GgFZpd3DUfLOew4JgtZWsQYaWjUTJ87abd9qjEi+dU1+QNNLlZi87i9f
i6uwfBoIuacWJ34fHGk64D+UW43NkibErcvhA76lz/9RqsFhQONZaBOJIUBpeAFt
Va19+FjWaSVqZy3B9rZdS3neAJN9xsALR0VV3tLdqAPlxv5ymRNgX0N7yUe4hfkq
88/HZkUHOF9zxr2vq85d3KSWNg6bIbpYcDSihP4D+NkMDWLVL56qU0DKleY8UvIh
7kgn8SAdS8SKHmK9BeSoIXQAXrTzkdMLJqQ8RQRyPNbm+nBZB2SnFbou2sGIhsw+
s813xXQLSyKncehrO4VMm/yeZC67Dt2sd6ITBfR5bGr+B4WPaZcLtv+IrzVUVaWe
uUaensWH0xsJNf3NVjYNIUWVhIKMhtI+biIs6bkq55bF7zTPLx8P1WzBuZs80v2x
6obHvSc0IwKQwU0kRdMXH8z/yAlGFew0foIEtuMdikmXwLBEKRbkDk4AvRm6JnTR
RU0hOteq9o1RgNAUKtLWUUg3suI6JR4a1Qzyh9G+AUd6SZRnfSGLIFyenV8MEnxk
OB0yt6Fu7SPaa46xiPc4zAijuAb4jlsRzB1U0x9J8pWj7Fm2EtRptzxOKXmVK0ju
uH2fQXBMAJPY1x0kG/YsCEljFnMmFWOz2+anYkHeLx7UEbNb0y6ReLQ1orKhKXbF
J3A6X/KHOoC3sLY71ArH7+m/h0h7E0h2QXG5zcPWz9WhhW7sE3YTOj0dT2UvK1Yu
BpoH0ZpCmmNmBFcpo5KG3W9LP62c1obmqEGhzaR/lso0X0gsqPViRFF/43l6Kqgb
DqW8ILzBB9WqS/w91ac+puRbmMYAIUscl5/SMpVvSKrQwqNmmXv5jibTR7YosHN8
Uy4ve5wEubIlZ9BegkCEL5gKMm59ACl4I9HCk/LBY7VCCm7AhG+rBFeR8Rll+uV/
OiZdHdAB24amOFjVGPTh7o4WFRARReAGrgcogdmqRBLKbEamyyso5HUn2ebQCnw7
vrOnq7EMAnOxZJ3Z8YcLuXdUp7g42ClnRrwBgHz5EDmgAoYXvhvF1gFa1burbVQh
Uh27PRaknqyR/UYVyE9jVln7sQGeYC7YIzaSi7tuTS58HECMskQ2egtnoCYywgAz
bRdaC9DK719xnBhsaLXmCY7nxOyCMkuCPJiAyo24EfTfJKyiY2hIvLTZ84aRroEh
UcKPUyf3lQNYYOjWU5TGG1XFUyvjVA2TnyZSMqJyJWlHVy2yOTD0xDptw0n7CATE
ptBWaT4OEQM0bwzfsw8YvmeonqAn/QGXQFalbGXEMit0xHOe28UmnTYKn/qZ8M1j
3FNnMXw1KIqmqD+wS0527sjQzXPgq5T3REUeRIt3M7xd3jRkAWVpjkb3gXGIIs9w
uzFG5gPHkcof3guOOdJ1i1R7ZeJZaJzUv+udrLOwuogQJvsDcRrwUoCIv3RCzwl9
fApR1Pub/oflmbuhJCqidLPYL63U39wnDDu5zqUyKKmVl3N3m/iZ5xu/0FWrH+4o
Qk4M0Wm3ISiSS1YxsDlXedZhbbWODGyqSiNdhXHQ/UIfz3JMCHstQCKyS0QmSp7+
tyhpSGKwKJfnEghk320kY2OWfCDX05XLnGYN/1PgYcAEzCjVvpxvO6lt/Sm7B/3k
uy3XQBjeG2B/gy4pv4NKbaZh3We0sTKb/1FLn15J5WS9dAxR405LQh/uR++te0fs
uj3mxvOZsd6fBpTgJUri0M2NuatMcY5LHSi/yA5ymsxT3nJrM8BWkle53IHwYttY
7t2gBZjzl08SXeSiukAqQUAzbecLpksRRcnCjjsNg4zroaPvRU9Bda3aJZifU6vz
RNrWOmDb7W25dtd9wMErgTPUo27WdicN0qlWfjtyPPwNMXszrAAcii5ZqFaRG6A2
bWUSjpHzn2Ug73smQclgQTlZLqHMFls8Q/3H9jcr306moVq7nbQQiJakB1SsokSu
CZdzeCf6egVblNhUgdOCUrmFGZ3spQ7IU2Jzjh48N9kXKuNlRUcc4jlz1QTzB/qv
7f1N5xkzbtwPVwoapgUoyv0GfgLwg4A7ZJiTOK9Utcl6cy25NriGh283RMpHbivc
V9Tcdj+Ggf+oUaE3qWGw6u5if1OG/g3kWTeDc3O4ESE1YEV8u8WzozxflXou49FF
Zleun3rIqW27Vv7bBaTLfDvBwIKpJE7vRJwG/tN3MvFmChz6khoRvjg02pT6QpaO
3OOe/14CZ/jC/QMA8tLJ0FZOKJLw8zJD/J8Kw0aXbFA4RJveVFKdRoFh6ay2RtCj
euskQVV0I+zrouG22UQYoHB3snQk0Wj0jg5Kl3EZah0w3z0G0Haj3vC5kda+84qb
3QjMB723VEo8sgi6CVA+CBELCcGOHWEAELqAqjxK7ucDjeJHmth80A5UEiQjLyg5
VS2sB7ANfJWfYH3F41ZJVJgNvqxoY7wHfP/ZqGqDr90tgE0RkTh8plc/mkqMc1v5
+Y9rBPoTcHnsP4lUV7dL5lPTEKx1tQQqRtC6gvh8MKfvyg6KTxhpfeA0g3TmGpku
oBsFjA6I/XRtb5XVJz/bP2s+nk7hIHn4BUtWNJKs/HOu71WEiBYeZdGnhY3PVH8I
wq7JZGJ8Tn/WZF3wqGhAQA3XDu09ElmvMevprz3XDiKKusDunAHJjv975WD6ER7d
UphKquX9bWxJNXSzvWUFTqcycmeYWonEOshGftxLIecNa1fFt2MsxQznEBpeBIbh
I6doCMJH6zxL6xo47QwdHIfFyoFZDVjQs+lPTYvHJDNlTonc5SmvQBZ7IgL9/3PU
386JG2/nVN2Vfo0Vg3IFzAQZYYHz/gbdjLkhIHXN70ecTb9ZpNYXqwkcpKfnmDZ4
e1rPbPBg/OyyGjQKuQUaAds3Vkdnk86M0XPwKy2sOnQRJtNrOZj/xeloIug3mO4E
cUz6qUXLcRC02CZbBcdRxJfkITE7XuKbMZW4ljIa5u03jvx4WSbs5ACQl07XOdNd
LOBQTxtl5lBLLhpx7Wn7qT2ijq0+pVgcnsvwNz2FDvqafehxrJajDzwkeeEY4rRu
O1Sia7xUJ9wViAjnJ2d4o3kcL3vATcLR5Qd7UQOECJ7Dv1kiys+S1kclaOxGHE0h
Ie94cEFeyiQJLgzGawUXo5hvSQy7rGbtoGAWfMTm0w/PNC8VREcMQn6xJFklZkDs
ih/6MBChy18JVLvPlQ89gqZaOvzPZ/zOqHEMSPm8mHAfjto+BzZqwpP9l7elHU10
huJuj68n/V/w0UIhDyshJpy93Vn4oSk7iqOzcAPK3Lu5S8u+7jP4gUfCaM4gOvcL
rMuwnn9rnbjnY+VZoAlQVxctlyOhmcwSloBi8zvhgeMSzjv9fQRU24dtnr8Kmdk/
m+hfBR0nfwPo4VRJFzELasK+rl6Sj9ytPP8GRvbw3TaI8Qae3y3YUAFx3/ZeXYR2
iXwCqAJcvt/uTx7Vo1wqgTUUF6OFD8KssK4BN4qGlzr+AjDbg0R3IisfZfE6Visz
u9wpugJ7uv3AeUYdzRxWBfkAQw841eOmN0EgvxkVbJ8qD5ZS9c4QYbl0G6pORHol
OvvYJ7k7eVQc5mt6+xxrVi3UdKtELALa8u1KzpKxtjmtJFssnycbHRkW9umjLKp5
JFXViBPZN7hWy3qdo3tSJbKlzJiGDdmElnFPW46lyUGqd8euDeY9zyRXtgT/px8a
CNu5tjIZQDwCHUBEijRTvM+W5uyaYHrnyDmumqKg0ihtYesAZXKOo28hcYrKC8vx
T4U8XRy+HDOMqQI+Snfe4oF1HtITkLQKMk68SeAANa1XVtT85oTF40C7xyS+C4X6
nMmxentRVXNCQRXmx3F/cB+ZGyiQYeaf2YHUDHZ+mc9wvQnGamCMXPzMEhIw+70M
gvhS27z4WWlc1eM/TFV7JPEVRpKmbysmsfpucm7zBGAeTd3crWSSaGEl0HVo9YsM
wq5y7Nw3PVb5U5DmKG3vxhRpDeJPVGVTSzxvBinqqpHTurs5aXJNB/IMtEopBbDO
KyviuZg7fxRd2ACevGQOqBXRQ4AIKk7o5uHZeNUV2FnS9xD2XjA7yAFRNvzmnJrX
qsSuXlKUrG9tpk8c2mKR1IfhOGDPn2Q9z/XtsKVgrioPpaSdKMGstJiwtM2KwW8p
+nmlQ1ePnq/s6ILfmoBl7TNszAXmu1bOgd+KeX0SVt8xUH5gRZIjUhzIaVJEcesf
G0r+zb1qZO5sHGz0GUM+ozCXTxqKhhR6J7RnveB58IBLhSjtbRHqWUEiOKQ4BbuM
QBuT+Dzdl60KUeZX0pjrYj6UkhII0H+XdeyVPkWNmYFeIP+75J7bQv7bn4EYVKp+
Z4rUyUV9Z3l+xY9lTyt2fYCMTGqDsDNwzlMu7fTrRt+FPHyBVrOLrYT6rOqtJeMT
hBpMmHHevIeRQb3dE/H1PBsdCrKSkx3qL88HF6tGXYeJHJKZucsAN9lfdDzmFN+B
ERXTs6ZLf98MVt7jWnGI/psOHK7kxF07ABMIP/tdw8m3u6XeluDpAJzO6uzjiLv8
tkB/e+Q1phsNIdWD186oJ3YXYvizF3lqV0L+8/7+9kAXe5mlheHLLl4zL/8LDkBm
pbjmGoJ6YqNQSyYDY09TS5qLOdWIAPKIffJ8j6wiEFJNg+Jb0bKm0A73+TL8SBzh
4s8cvr/oi39ubt5svWIxCASJe/Iaa/T1VIaEKYREOvg6xkPk0UUWaCaORGlBbQ0p
sORKtUazljtrzZ4pBG22Mv+C5ls4srf7ppj4o6jDoT2jxcLjhcc7Ec6w6qORpsoQ
/LDntPnBgT4CWlF3lWK6kf2NcOYC1rrZQav9XBb3tdwKIqyuBWsl2urdlMxS/hj3
Hb8y9VU3fbenvuViDoyhk2TvAdmCMWA61cvjW0TXJsAveT8OzPqK9GsXb87bIcH8
qxqzVp0guwouh1O9QFvG80/Cet5Zw8NuFpWIsqSJM6a/Z0D60RSKREszBL7pcyxH
Qc9m00WihhnzJHFaALL0lrH0w3PdluKQHjiYvH4y1KKmC+4SdJyFYrq6aunLmNlQ
SKhbWQrqfZTNJvdsftFNCWtF7N1kV8AKd8W82mKeBgknq0CuerxNmn1MIciRNyL/
PLY36zwlxHpUsWJInLmMg+2xG5cO5dHFlXuaassuXrBEzBrCddSLNuFHMrcGyckT
B8PhUyh/ef/qYrAUhByLqagU9pjFLeRLW2IDckZZi69vpeFgcBpJMJMf8DTOiyk9
QWWRaZb/8X++L4SEOK1C3ZfwHKpdq1mhXARxp8BQmv7KRoeVmLGkO4z/UnGn4c1N
7AfIVaQrCks55h8JcoHm5Rvvqn+zg+arE7rWUE82sCRZ5LZCEHxaNkPyrLJj+dCN
S2/bjE9aUyIxFf6MHsy0+pmvpvPY6O0Op/NPC39fL2Zs5E9tKWNMVdDS6dPuaaZ6
34vJEblZXvAVx9stOslJIjaN6227jnBd2sXBzy8jbGJNHUK8hWgUgrwFLJk3MJ9b
sJMd5XhhipOG0H5U7UJKY2agWLXG+HzJJhc/EoWo85WLtVPzCBnr90z0KfRPFmSa
4rremA+Sy7GPAevJXd9CTGk132kI7PTShoq+nXurwQ9U1nSK8M4fpGk0A/QMqo2c
fyVgzYAeNYiJIvTL2SRllrqK04jwFxxBWMxXSiRPB4K9N4Vi0ha20OmnBLEDF+9I
nllsCleSqzcfjenJ2YB8+6nw3+Dr3aMPM4Xc2pkrM8YXBXnU5NGVybEjQ0k725Y7
oCC4mMxWBKKqayfvDDhDC6S0+kxOFvznC6n1I5lgqFndTc8SNzfK5pYZjvqc0ZLK
JL0xiadffAGcHUx4c6zTyKDFR4tcOiESoByahtJupjGWq6rRIX1kaY9CzZq2vSVo
iUInxjopvcIfJ8P54TXnhEvGKuxH19Tu+6GwvydQ7pQvbCaoLYxz0pm4B+EG+5EG
wLc0/S8VJX6nFcqjYREk4G7VY7QXh8W474owlcU3f3cUyI2fnzRKgfQSgBrR15Yn
NJ04o7NQVS2KJ5RuMO924tbOlScuZfXurViXpdPD/RFGSm1n56GleSLzf1yDoFT3
5iVQu6egnSkrxj0KpsidaIw9IDJdJJE1Jjvq6tp79IvGOkx/hCd5x/KQrF2jhKBD
AelCP74DnCIXu2h2o4nJKcxDaWNvm0XKkpTMR5rAsOyIzDL/AEzmBzVFtBeIN+x2
iUe/JbUWuKiqny19hvvTJG0Iq0r+eLf+/IC5rQRt3qAiezwm+/gI4FZ+R31SAFdi
8MleuOgjMgemww1aW1MUoV6KE4RAKmrLSUsoHCeCstudMmnUYYl4098xt49qjrzp
dZuIj6kR8O6WnTrv1fZDSaWxSMox0Tto2Dc4OPAE0J+kZf5mnMLVtM36fcUEcPXO
EMGYN0VNSLCcDMQMdizWW/SJanz0f11ET39b2pTe+yvuVMAq9gKpjUyI1TWph/oM
Wv/0Vb4olZpwPMmoWu3Zw8gfSTcvYGaNAsmgRc1YDVSdO79ueEzj7kazz0NCqx1H
S8yW34aslTYf2HxRmYe2BXBW7e1S+FIdMRixB1L7HUBBjfNPvq4xfA9z1eX2bqRB
1nDY/vYs6m4rddsTQdVsBlyjomckDC6vaTJzUcGitd+cD+C+34ALxzBX/cAjv7zW
AWHAVfpXsgk+JpuBcSQMWhke+CZBbFMiMwZkkgmaCGOENJPGZsc4v2strvBB9nrg
wNGOvOavkBO5Y1/d6XeK/kCopHTeBEPkKkzYqJIjUFEf8a8aemLekhlHKpuXDCsZ
D5iaW7wj2nfKvQ6gSpFqCQFC3Kj+cVp0Cv43CPezBpD5ppIMfamysRDXUROdtcR5
qDYRpG0oR1o24LngsC8DLWtGpuwANAxFW66hrWOpwLJaUHuC3/J0sDV9SDuYuPtW
vi0PzPJEtysrPD4INJePxqCI3sEY8z2fGMp1ISOuBNH4Pb+atTCXW/1iIbRdWFtI
HK3iaufUAlFV/8gv2Ip3X/S8ArxDfgQ+zbDgKCam2dhp8ugocyEefMm1aSEOu92H
j1GSTaWfGsR4aqj6t9FFKcQoiyYMI82/9ZEEDSSr7AWN52rzq3l6+HXwaoCuLyU+
OpP2lFVURCy+WcUbLWFAeTwq15Uh7epIi2H8ZmJCzqhYDJuELWbipzTSyru5hVND
kQqiGOiATuDDZPauwFkjaUxH+7wR+ZYnGxkxBNc3ejigOpMsiBTvNl51WvK5szfO
8RYNrvv+pBjeDudrJxoXgMyFStUW45i6uBKIpxrme+ISnHpyHZNz7+6wkQ7Wirm6
zaFHs57nXD18ZWzH0sZm+pFD7G8S95h31pJuCTeXMPC19QlQyd5JYAyUC7/DgMcK
9OxwliMqoYp54exsD99r1H2NV2yYIuMBAMYJrWde7MfQ99bofZWlZCKwDA6fFzib
6e3fyXwkgZ1CwTHAcLfzkRTksB3dAuP7GNN99W4n/WD3eAmg6MTCcw1C4zUPkxDP
BmaEr0+rnJgkyaRh0Z6kWqoILtQ/1b+nWOLiIox3PJDU2Q15xY0cdH4HADeKGiVd
d1z62BBQyf6ffZfuXX6hAufojU1SFRExRY6wbsAyCeG8RBhPlf7gVc3QjJg+6Krn
LRws+LlkOuIFaXLzfmE9gYscTlzgt6R6p7cvvc8PJLe4CppjDpf4LfjS6KIuDvPC
b1eSu4WgO3Vp8cVzfHWgw2sFPUcFRH2T4qoIjhMyIJUoXEe8EkjJJ1jVvB5QCS6R
DHCrcdwCf0zh0ZkOUedFZ2fLTCtrp+sidCXx92B2XGwQ84VLubMhw7FEn8iCMowt
YwYc+bmB0QSgTqNaXmco78r1kTl87vF2tkzhWRvczSAJwmBGQ/Mfxw0bbgrBy+mI
VylJgqAahvY1zSUqgt25319eCGzfpnT3fJxVNQositvUYcJUfmE410IhG0rHuyft
jKKeAR9Mjlw9KHSlwsPs7CC5BFacH/n6wrawVNIlYTqBWUktxEBWRhXxP43kjiv4
+dBUYBMEnPxZ/Gi/QuejI5nlEE+9SMJpeoBiyKXJyBSfIQu68ChZ404qAtAKW37z
ye/TwsxGDTBHD4ZKDXr+3+l7VmoRYsEu1z2ll9Z6dRikcIyadDKzNVZEaPwYX893
5dEZmeQ2b7QWtMW+VQS131+l3RseaJL9fhhS7gy6rP6Msu/26nUHZurns4FOYUPF
EdlI6rjazuwhnVO9w+7CdfeeJWabhMPQ9ylOV+FvastDvcbHdl+r7K9XRYrVKQey
ttpeZ6AcfVkq6DgwnC5EGZLSDg4un91dZEpTj7Xn7AGb7AEBi4uYiluEnYaBm5oB
d76Ze2ZV6L2cErGrSNRZbdCEIy+F8aJBMKRL3SuVbZFUxXjcEhqLfwVR2AU6kNxh
so9wfsvmFkkaeipTdmCICLBCnvZL/5dTVpn1Nm/chPopKEHkky8qzjNIAxA3m7aq
DkObu/kjSsvqH3x6RLOVG0qWANmf3svD1wTtL8U1XW0Qhfdx4b/7KaBbfVyFHxqZ
g05UYnm+uPuiedLlY2TbayklfjJirHP7YmkJS2RAp3+36pu8MjqKWMSayCt5ToXD
gglXdi89g2393WcamoR8EPFhidn+LYxHHxJ2phjFVLVxBE2sA0iSiibTgPoDkByA
izjmJJoThGVHYXgj2rUQm3zTPfQ6LeYl9+N5CflRq8FBa3syq6NBzSiq3u1K78VL
Is4XPKVjwF9KqF9Y5Wp0FqjIW1vq6vagr+IpYxwBfePCragv8AR/Lw5+7k7YXnSU
g6x2DXKlIr5+esBM1iqcDbh5NhVtXknuo1wAeQoXrl7vMRdQLFyNKS1d8wwe3Ai3
eDJYcStesTbmahFPdvvIz29iv2p7tIUyNpwhbLlDEzC6v3qod7m65NP4O8CG/A/J
uTVzCA5CUoNS98pUsgACaZA1/CWrUFxsPEAGq4eOgySjhRuMt0JHvGkAaC4pg7Ow
PQYtA+s+Fnj9l14oCOX9i22ss4cn14dvfhvsCqskQdp+mHq9DIPg+FhsY26cUsYz
S4FXZgHdCglW+Whd1t7rCpUTBj0dZT5aCGQMqzoNii5ZJYIfrOUjXZdfrrDh66wj
OFAYmfa2fa8sUrMzJ8N+d6zwBfuDQlucP82YQGvy0lWJ5UGKw7mphxzKibZoLCP2
zh2DgaS2NMCKJtAYZ6yrC052YupbWjFQ5CUmrh6YgKGbkpVofBhy/QLoRrcb3LmE
lfNM/mJOQE3TP2DNpc8NrEFYhWGO3grm236+sc79ix3ku7IeImijGYm1its8RgG9
taKBo/V/ZhFMyIv9VBwMVpSbWoneMoKVEJOj5cU0Bq+rHab8D7Fy9EpVDsBCBZhr
YC0esZNgMP03imC83mPykbkAHHO8i7r2pgjrcKIJPXWlmmXpE7w0pNMVFMxiLcgY
/Ptz44rfqkxDdQcRwZDIcnlQKIwfIgWMn+u7ULIWpvgjjkkRNguBN3p52ybEFCBy
LAJJbLjeCfTq4GKCjfUpOjQRkIm+6zUqvNROkYqF2fyl/EMYXgOt4jBir8FVVr0J
SBUCFRhcHp3WDfyect4LGl+bKTnZBTs5sc8BZyjkD0z1nTyyomUP1lklAJ7v7VLX
1jhStms8bzcaAYZp6hwp0NyvulLWmbX+vvJRz8AFo1173cO6OBGZfqzs8jh2t5aM
GJ2RK2hcAHjh6eRZkhNHo5/I2iLWpMEO3uhkf2UCBF4UJHpIuibhRGyGucOqoPZf
aLNrNMqlub8ZqPq7tD+fnBkxAvzRV4cU+JkM8lE7W2Vv5PBFdnAoS/mAtEadhPV/
k8xTb/YaVPSFH8K9F5nsm0se0gz3l7ZgBJwLGzYJHgdD+yrIoO5DAk7/dKXpfkyg
XkOJAmRRGD9dBAKuaWwfAP1fSz73ZCnUOyvXw0+8WtFZG2gJJj/xG9k9jup1jlTN
8SXeqWG+52v2//0/6q8dEMg4z2I2yH7O1+95Le/Qjh+JNjKfWjvYXJfvKiC29oCq
fMGIMBEoan7YMrWnwHOle5HjCPYqDeUnIdyL3ofa2gOJse8jOhIQA4zgi9Z1WUIu
LYVX3OGLGJ1LMwE/UikPV7JZltmx6lkA0OCDspnPTVHz636IyycY5iY02oF8Ij4a
7EgbakGd2ONmnnULzyQFG3e8wVLMOcznGyWtdcwi0QQ+RPWHZTdUcF1TrIH0O0aN
VVKG223Sbr0R6FA0sOa6kgAHB8XTarCu9IaBvtRo4ULlfJ13LHQZRgh1/CeoTRo8
ySpajOHFasi+mKLnOBoBrDHIDiloc++F3F06JT1apw9WxPl9ug7+JHBQqFIMIhrH
dURmUNsTtMvxM61A9JZrVAgOIloBStDnKCvOg/s98ZyZmQlQIygn92fMPZUlpwlI
KbknaBQ/Uee6hmgco/kS+t8zJdj+nUsnBZY8o8ZnAMKw44JBbas3uWxgz9yLlh3F
8nueEH2qHhY3R8RnBN7UGmc0F4zG8Z0vOj/vsJtsveNK/rXHngJcW9G4ZVpk/Yij
jsdLatE4jVadQIq6M4HM3JEnseUgpzeuIdScXoilxxDuXT7Pr1XognT+MuQ2/4s0
rJBuOMB0MW4K9L9CqcfPK9AxXV0hEA3BsNXqJIzD8awdj4nW6Ww8BbUrxTtrdQem
ynkv/SDG4ydeewzPeAz0SZfKR5zDcvmKKVNxP82IN/GFf/4DkvXLXV9Tqbx5QENW
5ig3617st1sv3VRO99YTAbqsmEClY2Kkj3lbeEaHaTAX8m08mYaUqTSK+/fo6Q4X
36zUcLfTOdcotCqlAyQqD4ygPu8+uSb2xos/62lxubSo9lDS+CSS7JhtDvtNjA8N
YG90j4tKlvTUNJ3UKju96J38NKPWJIlv6SkHrbiJ+Fd8/+mbk0AeK1MxSPAlhTm5
Ew4BBtg6bNjjaik2U0kl2g+Rm0jfuOKk0ppH2zbsZ152Z9J7lKauX7eW0HFECXIs
fc3i7lNe7N9KypFHj9YtgGK14bvjIwLM8gX0xOytbIsYRUB6G6gulmWbXVgRJsFX
K7WC9/FJQ9YLRLaMNJeeVTdCRmZZnIo+0dd8EO+Oza+k1pJo8/lf35oM21e5uYDT
q0ShTgP3xwtms6zZVh8P3tXKgq1OGOYVqd1zKk9UdDmK5slnbmAtJ46UPhDYx3tr
8ObQiSDzc89mWnTqjSAN9cKRdxEt4hIW6uZ7adED+Frsy0iHQkOCO3Gb6YML909w
beWvFDrpnE2MfyqXXR79XGnyWiHidU43fnl1BwxS4FE4dkkbbtIt0SAupHWNwDXB
AnkNMdlhuf4Pfd35CYzYVYehqa+vkpVtW8XdyNgssCk2np8P2O0K1sSXTLJ80YAO
yTAEkyCLtwUvRG8cHdKCDPLq2iTLkW9pfQXg81S5fgJIctKprE+An+KSGm6Xhsye
14lhQUrlFDj6lNvzfEYyqNj8+1ag+Tt/iEFUehakZ31U7+KQxJRNhf9dZAxIWysR
cbG8bXa15oDXAGjtJlY11Os+CdnEepSBs5sngdV6/YysX1pxLl7uhfG/bTKnlpra
uITE5DW98qZL7x5GYQLNpTFnAjnqo+fup25ETgtzdQPt0uRBshM2SaFvZrF1i9UF
cJnvPRLr8Auxo1ofRnfDQh2FyyKTO9RSaVm4DXv8abK2ogQlktW+zlqsMTduI2f2
XTQwwi8T36k8MQ2WgnWKqIHUi7Q7LmWiBMNHzEaPu5bGb6JSUShs1/wQfgdCcgqm
FZLf7zyPmYBfs7NpGUuxRgEHg7BbqeXeSLFXtID5ruVHYij1NhsZoDUzGv92FAjN
zj35B+BK/lXR4OL34oaD5ZCUn1/zx+m3dqDq1Thik3mIFqr3ArrwiuHV0dBdkel5
55vEjCRMOQucwdrKKzDkWw/2Bp0kBr3MvDUV/GtisVhDqBSK1qZC6wBI5dAvGjmt
9et+3OEl6Gm2ALEjYBnBgAbbfuHnW3e3c4Z4AskF3Sz1JXGjDcaSN8OzE/kPw+Yf
kDcliuNKWIwGIpuL7D6uc0phAvZW1oWp5Bq2XvsLZD5jwrIkVtyhr0mw8LL+PV+L
9VZXDQpI75jYBkyTDmH4Ikq8Z6n/qE4F85gzbTSBFm94tHWTHjukw4ujRVLR2Kfe
KM2yll6NnsY9NlC3sxChIajSc9wMIuNjoP8GqzJiN5tvcASDWElf4vdF09X+sJol
zBqZNRxamzAjUbeCBzKiBUlT1t0/55995AStGy3elEFu+qEL3s+O5o/sUoYTJ/9Z
zvNxT0R3SdFx9l5LbDjsPA3ChnzWHeXFZ4B19yvRswVyCg1GRlU/3+QLz9I99NCJ
nRZg/D2jAyiP66W70XuVkANJjAnbp8D5KQiVaJN2pGM2wsIfH4v8GuRiuWo5rVrO
uU+aI+EdU4qPk6kyWWmrAJt+DGSBX9xWG3/Tvan+GdOsUgVrVax2baj7ShzqpvlM
H/BSpG2AP/2A7gL7xRFdEIBnjr9gssBNm937JYdNCa1wDBxnZFJgQ/YkZ9+/0CtV
RVq6S/OPOhjEbslzYD6pLKEpl+fFi5JA/pkURSKVuRy6UeCAYrnDZSfEOZFBJCsw
9/lUQsiRH+YatcYaCfPyd13Ppq4FaEc//WoA+xI6yG10FpZesWyfq16dyIc+Tn82
M5VaqPVfsd6rntp+7M3SogcNWULkfs29PX9hr/7hrRc0BaH7rQnrj0EusgJoeKhU
K0z25ZXb/80/xOYazcXxTbthYhvgFPXaSN6hSZToswk/3WuTSeZaVaA8Ia1yJdYD
uZIeR5NRxcnJhkObyV1i/WxgheaWZMB2cWARJ9n7YN5+7bu5ETMnMWBl83Num5My
q/0b4C2+pGXq/lLHD5hCtD3MArm6hdewk9n3FHiLiASXXA4KQDE+CLWRdhjLT+yX
slUvG6FaReXuvEJNr7W83ylre9ai1hD6TVTXocXRe1C6SYpMNAvlN3V11c7x8zt9
OSNhyC9LLEQJcHIO2DiDXEvUBtje98Zw170lV38mp2Y4jH7/NcYgRBTBTD8vcxen
4l73AFUG0vKXIW57tb8XMQUkEYpS8X6RAm9DIiBmcOoLOSODz/r3I1YrxfL79SU+
0oOt1kyq058AcWPI5pbYDPSV1isrwt/uD1y08wS0Eb879xY/Qq/8FmusR3zQvfgr
sEPTuv4w4IDRUU7V9buGzs3kLwRYNPiTSDqEKkLOnrmnAfJJnKE1jJ+uscKi6a1H
oUpcAl72oYRy5RRuxFqvUKloKsySB1LUkxvgnkPq5OSDv1DShAPwGL/WPFku/BzV
dbM/7f+d9DgLUxwRPHhgi9lAglYdY2FlFaxsq7wfnpQdc+8g58qXvoAF4qGcrMh7
Axoxp2s7ilU0GDv0U/SmrAFQH6buZjy3ILSiQs2uENlyECFEjzQOUIltaWbkhBJQ
LNuFUG1EPjcaFuR18n/T/YU+wxKLKMA9es4m8qGMy/Xj1mudhP7paFkeitaNzJcE
uBAk6KU3+ULoe5HOAM2ViBUNs9YtpOpqiuOamM6Zz0D16sZrbXZQhZs0BUKngYKa
yhEcmSwo3T8VqetdEMg99L40SJjjm1m6GoBFvzoTBsQiIOoE2+gtNHbsK51sNaOv
Z/CaUVVVVm08kro3FTmw5BGOzIKSrIxpINFlEWwDf2MEbcOM3N5hlZAg08xE0qYH
HX5y9/QiVbRRlDs1OsZ7MxchOUk6PDiN34mgpBouKOVGmFB6Jx8XoW4wQGjvbDrN
6wvRjqz4GiMpOoYwxVCN2Dp0Kw5qI3nO5f/9mxY88hdNPLbCI1sMc4bnQAhVo9WX
1cpqlmJ1YR5igyrMj03gn9LqePnLB+dxOFDj0J6zlqgUTttZE4Wh34FGmVDNWJPB
VtXE3c5YkQRDdLL04SQKhWQnRDUJtknMlPmS3KOoG0hfzxn+C+2hJ/xWEd6Y5gQy
IjW4+S6Laf0K6GG6tTjW+2OP4xlIm8Q2fgf11KEKxtL/N/+fkKPJKiajUG2UBQav
UwROcG4CNImZxzUFvyKjQfFN9WRyNzpWHtT4SjLPW22Lp34ZmHgm+D6sdQ+sFH/g
grBABsCGuDRsambXIrYM+kEiAxEx4oxMqJQC1r0Z5jMaGHx2Y2XfQlwcn9DpOLu9
jD0Xby8ra7jVarSOtwEqhIfTJzjgFGBeTzzr4TucnBnr+fd1qRGoCgnRCOKZwQse
EeuJkodWprKTm4FQrTVicZIcKIl53JKIoGJYkSIF7fy2zIcyF7ErZ7ZWsXjpbnpU
OaS9cGRbBPQL2NrwKNDARWgeiSVwP7KC00x+lvwAPL5enLwU4S7fjrANYPRoehxF
fsgVFvsNrUjJyhI2cvDEMyBicWh+thPteEtLw2K44gAY7Y+7B7sihbMTWt2At3cp
AOlbJr23g20iURVW8EhvEeKlop+aiI+1pqBOAkEa6U6NplBs7poUO8X0YdBCFx86
YlvuV2RxIaoYpgF3SOVDKeImxdqbFhh/8XHHm86PTqzR5Swb47vtVitVyoc/RiYC
6u+zsS5SQc49hdbTuWoVxhLrnjwLyhbwZkraC3ntSJhyyJt8yCYD9FnxKsXktOtD
w9jkEEyNrSzcKGmxoIa6ksTXW7cYlViKws/5hSdQuj1gXLXUCuR8ROznyjcznnFL
4bCGz7unBc1Ig90xtC5UeHpgog7Cr3Liq8gbjjQyO7R1BFwDo9irfFotO1Hex0vE
z56LQ0nZ+/otMIpA+fuq4ZjoqFzFh+jrx8c7nU4Sg6kh+kPRKHXJgJrjE8maGTqK
Q63l8d5aGQcoAZgrRCS1zCnISIqOvKA/czRuP151lTx6HQCHNN/dFL+hPr7NsQqZ
p48wtnGcQPTDtukr+nrrdt9se2dwFax5wzhkg8QDkrwfiET4cvYNRE36UXVEMI3O
f2/2BH7RH0+yVG3cOZ/i70L5fLpacR6EpQnsIlXwsJIRzOIHRhC7pplkeLf+54La
CG0SYLCjdF8+Hf4Rg/MXQaLQfV22pH+3cE8m0KMnec4Lbp4J+iW5ei0BakoQEMLT
VcDJrS6nxuq/qaDPG0kb2ECNEMmX5uA6Mo644iS70Hn91WXFcglPoZBjARRaRhdw
e1x+NN22JPLYEF7nUwgiYcq/CHOkwRAylXgfpuGN2O0VQ/u0fMWyqDgU0I5nxsoJ
Mc8qcgaAz/M/nH/QTuVCXhw2eM8OyVQE6bRCjZNB3bcnQ6M7S9zIESf0s2uDD2y/
HwPW3wonDhSMtXeLcImL3tvz+Sh+KOtG1tp5BafoIa8JRZekbsvWIkZLm3lwSZCC
huw5ZLHLUQR8GZR6e1jhZUR4zyHozAlvoi+j6St3ROV35ODKKoGgow88SsmaGD2r
p8PS+M7q5xIS8Dwy+LCQRvgJs8r+kq69w1izJ6jORds8xPKiEYz/sP+nAkZ9ABmq
nnFhdsaucOj4aClI+LkQ2T/5o0ePLVoLfhRqW2jxhxLVJPxen1ijM7BuOyiy+V1/
99NzKxNVnAcYw+5E7glm5C40o/YizGLdID3zprQMgVEOFILLVNC0G9NdV9xg+Zuw
3yvIoewdRr9/j2fb4Xrrlk9YE1DXw665kvEriv9Hh2waMrLkIymtVztvjj7zjimr
rKffChSuo2TWjOzawhUTLUpkdcLTgpWOe3U2U+xMQZepAya8lEFjZFoKgNDzoTF/
mDQV3O24BMyOGrP2t4B4h0OtDeMbIuS0eqKAbv/di/IUEAAk0c7Gl+JzPhuJdJHJ
fLvsXccbTqp9cKUu58Nha4MNvvioz6XmPKwNkRFTTjD3ZzxWXGhJVdq6z8kaUpbU
CVEv+ZnZ/Xm08Ql7xr7wR3mJSy/TnQCLvx1NCt839MsK4ychH2MfilDhKtAaooxy
RGiouSguLq+MEIeHASP0G02glJgZW/DHZbOu8LQIwe1Wm4dPIKPu5I4+DrVC/VKl
KNcArVscvHVz0GQGVkCc3oRMYawrlm7y85JrXG2C2MzFvYOSZf74+5cLSZyGw1PH
MtwI/VZB8iPI9CwWaq+gZYHF/4M6eDdOBYSFLdbf8k3qCf6H1u4tL9NsTTvORgII
lhpG0XGAtBo2P9/auPKs7IlezRcxsRGfz4RHNU360uJ1iEh7nvEJvcOvPl2CUURM
z3gmRQOcJQ5ikyP4gkTjtsZ+vDpQUCO5nPkjJNfPYr4N1oeticQmyZr0sv8Von/3
BWPoe7RrnlHiRcudWULp82BD1KfBQ/G+z6Vz6MIrz5SVnkLkUFenXJCRxHVhMEX5
KNwQKMuY6XYP7tmVgRaUz6Qk8sZ5LK9iMOJ6ZQheTrbuyujevn/4PROZMWXxDk3b
vxV2Vry2YBAXFZLtAFAt/Z6VgcJlW2UG6v0vOgMX7QtK5DKuEakba/xGrLZXDvLA
uthAOXSrzstYbUsLA6UP0YsSpJPCoUB7LZqTGXSiVAc+s4fCVv6Je76+DrpElST4
OHW9sB6VBN4axEypxxY/WoVjydcke7zZZdyaZwVIsYpLv2hK0tu1dCW5fk6ZhEvL
tM9KXT3grsgx0eRggpehA49xzH7HBR5C79HZmvIx1zQs913N2ORCt6FiZEhhOTyS
+5hto6d7RYQNOlDHDRfaSd4pcQlihu6y/OvYMStCdkq3UXWUAi6cPUNe42zUnqWQ
OC8lxCwocxIDUaM8QhFSykZj525cfVRHMCvrNnbBxR998JHrF8ZiAXYvowX1JO0F
0PRiMFsSKmfQvf6ZTehYE/ii3YeYaIvJfGVeDVpMjMj/dCgf5acoOfSpjSapfYaX
vzdN1VH/7BDDnn+g57ciTw7is+9cE12kmHmPhbMWXydRB+CvydkRhSo34AvacqxZ
rqKaNCNNlfoJeKcREAuJdfXFaNg3Io/H8WovTuct+NJzIr7fI2gnKjr0gUnHx7JU
awhP5DQ+QPq8yIgPn+Kg3KV/8epg7hsEFyv/XJafX+eX/qVM+n4d2qeyia/k7T7Z
ToWOAF0DGN9MtoiXJucji+SDYUNVYcmMcAeCkjjXhEQeo6u74yOTs/llG0TAmXyE
piW4OzCsD3gJi+2EYbCWM9H5McGiWPo1bayXC7X+CshQa+sOl8+sZbfZDz0IfE8w
Q+A6CeWqn8i9lCT/wKKvxvzWp2pOLHxxRTWO4qklylno0fY9Hy3Pv375PLBUB2H4
WgmUIX94vYRYv1ZeNuyxuKbdRpoNLNVjPK0e+oSUHWPXGV6EL+Z0LN25QuMRDsdQ
oPCOBQAZWQ49xms4viGjQ7LtqF1w/RmzYOSvKQJfm9gVsf/rZ4YKr2iGaJD8nIWO
cyN180sQprCli71uH8ITjzhFo437etw5lidpT1CEsp4mD3tY3h0Hn30WMxIJj5kb
e4ufkTrQhFweGjTDRtg1c6M9PGImz/xHcawWvWebuke3viVkWkpfsehtkmVbfX3O
IqjfbBTVN3gn2Yu4IJNspf/90NVm3cWndImpAScHO7e91rCvCs4hUhJm0VVlk1nf
BUZ0y7TvcxXrBzZP6yQ1Ji5eWRPLlq5/me6BsWRt4rOduQLOvm6rk8SBiyE0av67
QIuumInnI5jbuYWacCFTfv+XsWwj1Z9gENKxYjRSAspFyD5A5P9Txt4djG1BXdIn
RLAGOYPwJK8VbHF2AR7eVnH/dym23tYINEXBvIh+0s3bNS+Xk+6nuGT8beGMwgxQ
LnY0EnnCasMusGafaWQZ2KcGyvFWxASxWUSSjaD3/lWu2iIK+5cZYJ5gEgF8Cpg3
hkSy9rTMpLpBh5ONuIVv0ZrnRzY21VaqnIdckDjz8kPL28ljBFarY0nUrjhP8K7s
nE2+YnS4GFX1w7v/w5CS1wZZ238Jrf07jHRv3E8LjVLOgaUkiVV6bP0cOdpvLWxn
BhRGL7Ws9z04sfcwyAKlHLRsCDwygujn7LOgDNeKEZLxo2GBXPscLjrElvL8v7m4
3tom80nF5i4dBu/ftsHBmwa0oPOpVz97fTb7v7WamiwQs6ucBL0/3Pkv93i8E6L6
bl7ChmIB29W8Oib4DOgPqajUdOlcMACbdgPa+cy4KV8B3RlvA7LjFrI8BGO3/CzH
Ah395GnIM2dTyo9todHh7O/eyh+Ryj1eb9EnK+pqQdgapf7k7tiOCae2KrGzS4X1
8sK599OhCiKOeTBaU9ee4qtwg4zPv877YyI3KckKUlhDlcxVl2aFlID20p7FWX6d
KY7UsAUQWOze/gArBz4avCnGEUwSQefwLACJACDgWhrMaCnG2mGJcnDmhGmUlJ71
5lJHRaihDR7VrzRpSrrfgpK5SIwWSiT+nNlPSPm5GwHfd6qADxRC/68/qmiIZ04k
bHSzMx6vBOZL0DW/FrzqychvYJ2uZ2JOJUCLebV9+6rh6Nux6rGDIMGKR7GT9gYL
5pST2J4JKCA4Ba8EhP+ZKTvSnZVUiiHtd8IHgAQeM5VwNydfARtRkd0MYwDvxqST
RDNeoEBsREiPO8mRAGrssl1RebTKvYa53SPLfnMVOa+8gTJ/EPlVvsyFRvkQOfva
+gN27I/qZRdcLrvL7F2re/Pln0RYhWTvabl3EIIFPjrMguZXbQ/LfyVOhB62rIE9
n/ruqXZ47LJoH6uykyYG0nkp9yQYYbrHNHNecviu/1EhTy1ZBG+bGV7+8AhbCM2O
fK5NApXx4UqmCc37q9CCZeJTpcBSAxQlEx6VL1VWZPkMjKEju3SBAjmKDNghfmH7
XwIccuJt0siqGVfLOikssdAI0f0TGqxEu7p0Kt2ncezwCYOeLDlBW/mIJg3yKPRh
I0mW+KIQEyPgEEJpm/eTHarJJUPCWGaRFOcpbGL4VGKdmcNMnLd5H2escmVAO1eA
xnUXvv0q3oAVNOUbvcHDJJjkVaBdqSDbsQzD+5s97bHoHana9OeNlyDCkiKWjiHA
uGZMJiC8U+Wh5Q/jQ2X3rSHIjbFMRI/yIThFJXJrgafG7LuggZJ544UzgEKixZn9
QZsHCFb1Lan8dw10HWAN/D6WeFlD6pyekxCmjhSMrBMLs0sFknslYCnFffyrvwsx
y4a2IFBqLhbiLHvTP09oYtC5FC5QFRVMKWvRzfbj25S6fqwAmOIrO6ltxd9+wYtB
5cH963+/sVIAVDRdDi0xnALzPEgDyT7pOG71yrnkB3YfMUc7T8QL8BDakiUwlUjr
yTyVzQnOiG3Huqc0MOk+zaWlTpIeF/IkXTq6g6SeDMwC4HASj4ICK1g7XUiP2jxQ
YEzzGsgkXnm19rLQVMY6Tzs1laoNv+mDQ1iHEYayG6PrPDzCi7CBfDl/COh27hZ/
kD9UvqyKE7vGoX4IapF1nzDFIDwEthynO3loyeuVF22s4STovBVaXc3NdFGjTKZW
vv4NcsVvzfEaqbjbOYxeeznQskn+qE+vAVD5n0WenF0MqvyCaKT8/gHMIaBgjQrR
BrlmlF3w4hmYG6E8oEIi9Kr+KdguhfTOhfitJvjbbyE4t0i7w6SNq4giZj4pWr9Y
zPBMMNVeIYGlOgqx4WQ6UmebOxZDJAuipQqYJzlLcMYkn2c5EJ6CRJwR+b3xlu3B
oPoUw6msajQojk+nClLr72h6DNe0lihcgCQDn4IeWcdeOk+GPEnXkCaXAonFdVs8
uUHRiWRP5I4zbnGQOrcpfHEVN559A0WOWzXafqSvpSHExkgk6StRTfipD8gAcWrM
+boHSkxSlbH0mJjK5r5/Q5PUmsXr2hOtlUVLaozlG9bceiZxV/NSZqNwAB3ECG+C
Nr/72nO016t1/tgEiWPB4eEBhglR4FSDg3muDDIxtL9fO3on9NxyftQbEllQ+NoN
GG1f9wjguflVThTeMcGW2Z5QREZQBx+wP5emApa3FWGYPlp0QcS+qFlXMvneNDwB
pDwe5oH7RMKTupowNms2JLd/acLKe7ifirWiMFdrUmqLUGZIZWAkh72IOBWyurSL
1bEn6bhRUn0NTLE1fc7cA3G9HLohiPHBZCRL8JO2u8EDLzsNcOk+gE3iX9IBlQDO
E5yqKQrFXhF04TTSIhFvZOBrLDha6eFb4HQbfRTf/IdAJzfMqysIus2AFQWHqWUh
WG0udf+z8M2wUV0cihYuq9aHJyB3Tl0otrR7lQvmfTktY1IgSRJlPALAhR9rwKV9
bCzXeFjqVU/PZ/UEsTKIyaJjhnJyPRcLZTcVlO7MWxFwitqj1w2osF/HArKM8WFt
YQ0oktABQA9sO0Eigj/fMDvwr0znblMthdTivO/UvFRWu9/nNmfrTeFu2mS6WsWw
TLJZR1JXfuysdLIg91A+55AA/2gPZ4drmFYvkFGYYjeYR1U+gAAaL92GY20xJLlV
sEv8UpFljWkrWKuNgdKgWd7XNbq+CC9AIq8XYIo1HN9hQOOSMLvSaRgAdrcRXtH7
7PJJu2qGjQ9lpCmhiNO+f8C5JgyiPOG4HdOZJwWGAKKWF7FDksdM3t7AW/RtiLbP
7GX9R9JGjyZz1eINARm817EuabodBY9K8DxVEcuUjjgloD53FthmF7/wlFOv1CcX
b+dAD3xlS8yKBBC0A3JUqBvNtGvunUuDeh+t87nAY5wrUHh8uzQeQ5kpUL1cDZaZ
eKjZCll3Hg75ppEV+3V/kflJqrrk5tdX3VYF2/qmFxacdlKXmSjLBpJWYvrrLt3Z
xn9CkwF72QfJ0eek5pCvPg4stVZAh38Ll8fU5tuJ3q5sn+dovfkiNg4AK8vrYpNC
eniuXXscJUQdVGo2nf15kvjdASH/kzNtpTu8Iv58X/Pmj/YhW04tWiBjN+p4M11q
HL1og2SO8SYUGzTzX0G73w1KHbm6KHiYgjiDwlXZcs9yvbRhg/d4ii/XhVBIv7iK
D2D7vxSZgjI+ZityK7+b+MvaZEsKt2WdGSToRE63VHrqykqaY5CQZP7x4YBlMC6H
6fqim4FR3j17w86R6TTpG5Q5+ofnWLktStqwWfXnYUhge6WRQPtygGy6L3lzrDKc
kPHiPQ3EuFprqlzyiIBoL9ob0+rDwAuj8OUxrpmOfs0RZDfZen4myXnLB3GYaoo7
mguqt/nLs4DgYCXSoAdRJnrGe4SSYLP6EXmwEBIdZAtEPcskHWIZe/HAzalbKNQX
wX1u6VW+uFdXA+pYz6tCdoucQLx3tg0aomBy1kgyDn//p2KjHrhM4G8C7sS6rTaj
4FyugnJ864BKypCaQ1dkgc8uAZU9vJ/WMF5mqhmtRWM5A3fHQlml1hHkffwPhvGQ
6al2bAvFcweffc3kvzxTdj25OUy7yxE5fp826zoDs0K92mdmg6GtpzIrJY8W1EQD
ktUpy7IDUOvJASaUphovmwprmJO0ko9lv/44VhpyzGkgmSdPSdBfbuou83X90vOz
IcMZzpphIKozHfoBM7o5XnbsIE78+Wpsree0obLXXd82kh42Es2AksurXLhOWy3F
v38wT44yP5QRtgcvEsh/HqDkeGJqVakVQh15/wPiGdf+ov/N34/5eRxv/N/N2mY2
VG4zcT8wrjQjpRcg+fHdeag57iuzDRWfH0hZAUyAoiArwFQVYKfDoaCH28OPdUT0
zegCwCli4D4qjf6uLMWrV1na0VxyVE388Jo6UPrX8NRoboSW9b9UX6IX0fvCW0yC
KGHnwv68l0fGWFPLBvE47ocrCEAv11Bj6hbtXuET24k2DV0INaYEUmyhVijQ7B5n
xKVzqjtbQXudTYBISKJIJzkGLqPrir27f3HivKYpgEpZwYj3GyzDWZxVx0nqseBF
Pxa3Dn3oLIJegvHuT+aWV1NUSDW+msxzPbRzve7ERzYY1RI3y8ddQap+4xESKH4G
I0LeO5t0GxP6JmPcIfvD79s7hwJog32q+SJgD8kkC5SlV2yAo/NILbt2zxxTRxcS
R96MKzizavjjpM88L4j/531u7ZnJCCJalhhYlqCNGYdQfQ8AxCLuH3EDKC16CyEO
ahobBNtOduADXRbDJX9M3xZlm58gL1hMNCFVOD+ycH6FysuF5iiFMwPQVLf1hyBi
xp557p+uxZ6HWB0iE4RMLNANLXK6/scIJ/N8rxt74EIVAET09rejG3z05PFVATid
92qmc/sg+7UYoleTWvUOEvUPpNFEsWfzeVcshl4EyJpoFlIwIu6M0oukOrhQtKVz
DhgVljwoQROsMJFR1a8Os9CWSuQogrDsZFBuCmJmC8zV8v1wqOLWWO8yWYTnKtvy
kk9WvCGa+roZbdAXjADzgeU2QDVawz7pPYKzUpXqvskru9Ac1JufjJNKJsjw0khB
X98DPwqVMdYhglF4BPPlajICn2sv86xCodZ0x+JmZoBRgh2eL/U8duljEv3l4eIN
bRrTxIfIeEk3fGvMwg9ZihrUUGhdbETJkYJSkU5eJmfEJs9OlEwCIq7OZ9JWSX0j
xJKcw0OLQOJ1SHfpIT8BGiXsusDzJAA7o2L8yZdysMapFYVAGnEyT3yvJdPG3v7+
7BDCi8Az5zPp3D5tfLwAMjAjjZfHVuK0K8XGzAvBGVx9iHVimlIptl0fu80GncOe
KOrWintFxojZsVM6ol2Y//qr3dPpSBFucNIdio7dzj/jgl/eKuojBARtLxc3eot1
tVhGfs7ySqNUmTCB6hyZxdq4OUPB6Gh3CIE1BSzRqEycm3zJBAgvIoGDtjfdgqA+
wJlyhnZu49VPus5GRBumYQXdR90Lwrco2f3mIA2VXd/JI93+2RfELH2eEDQ0Tes7
h/8C9FAdUPyr+WdjOoxDNHhLWhhqOoJS3rSwfjwDrKtAtUgLklelQdRr/nLF+ShK
EsL6dccFup5hw97Sll6AFZVhr6CakuopHK7gwkBaeOf84R/cGYsifyIPNYIt2tZd
Vs1dKkx31eKyqEipsV13cNF/GBHK6U5riwkQJlMZlqyX+85+Mr8DdwtJjIcHcKw8
LyzNG/6PwaFKu5ZYROrq4UXJ7zZ3jnDHB3bWffAWn7g8+rMfC5YfQdVZYWJtl+kA
QY7BNLXNCp8A2usz6s/V40vUP+rQ/BVwQ6UVU5mF8uROZUbn4bGOhaZRzpYsYMz4
oC6xBeFFUN6R1Y2SR7B7PwgHC+Koh3bJ3ZXHApdVjFfQp04OGXzbhTlr3kx4ymt/
ve3y1uqMnr4LnAzdi6Hs8j0Bk1VqfRYGJPmL+zpCk6/jVFKASkxrjQpKV84dZhA8
fsGWop90OOU6RRxDgpiYMSIAykeR8sO4T0CkTUSZF942xdcv3GCanhFDjq3Y48yY
pam5LBICPdzVRz2MCIaRKTpn2mTEK1paHVWnahFgVq0tGclLo+wtWA/FTAqQ777O
byIsKieiNMct8GHzzTu8Nbcl61Qp6NPMKy2AalPUlTVCgTDYSJDmQnRl5Ty79HHC
fGO7otHeqNtyBYkH4o7it12m0Noo4XK8ftEf9sm/awc15l0g9GishVZ89RI3C4K1
wsRgMw4r/JpxyA7xJTEYxcOineZXkfxzShuoVPAJxLcHwBtc3jsrxbPL/dh2BEfc
xqT0x3ngei3J2mAMBxJX2gLWfaFvSirxoZj6teVWJf+ZLjl5hwYFj8GWiPhsEgEY
mNsl4LvPhBko10mf7nkWic/urLUDTFIVwND8h1P0DsIVSQV/b+hCa8adcf8/Kxy1
7H7HNqPNJOdWPFqnV9A947XbOckCkhVOubkp2fkhNHnwgj0TJJpLk7nd87kP0jVx
TDrPFgC0u78TK8ZihjNXBdliFZj3cpfOJ6ZiTUuUujXU/9D21KSw99WTKvcOCQIs
oUGy2GBtAaSHk/IACGXqYZ279dfOJyt5+yEOCf8/hOdoEoayWRXOOlKbjeLFvLDV
2gVrfXrWJkYN3w2Ij1TgEf/EpiE0ahpRw55mLMZf1ktQT/gYR+R1hMTL6vo9HBL2
Qvfh+fiz8FJ0syX5iMd0GGhM7hnISSDvki3guiGafkdwIjdHrRx/JYjN5cy+AJQJ
YEpA77HFvJsMeIuJ9UovJL9NHW6frDdP0wd1bWYzJRfLIB1ZlhsgkZCEoLCojDEh
PsAgPnHUV3tOVFVFIe66NKNc3X1w1b0gDUnpSDQeE/hyd25q1we85ql2q5hOZO//
CMbPcjsaiIFGlezdZ1mxezrmnSn41IWoPVGPGzKBgwKkzyTe+omuENVyrtvPvGWd
iZiW1uzjiRUEIl7XqfswjSv4Q6QAypO0J833v02rY24lbMba5fjHu+tWWcMWJFCK
A1m3OLvU8nHG5leDStQQ74jQ3I1qoQ7Kh+R5WunKrj73pXnHLg2JldGFdts4wMeK
G79JaihdT7Juwp0hK+9RjQJupW1PNQXO51R35wZjy7Gp4xMy0wOwFsywkEzjSlCX
Bt+62PDVAnJXZ95xtLX8pCRYyBbG3NyaXb37YhQUVVGqmxILjLLKTwwAMaXJiOjG
GSW4MmkiKDMeWM7+jqTkXNCjmrQrojI4KPjS4y1ulUrCLCpfoR82KzsMwVmiSGBW
q5JOBnQ9jXt2TBEreebTgIcqLWLR0CQCHyKX+WR6CqwiwSdLMdS7jlsN+qq5OmYb
Akp0kdTZgAWHX/hRjocXfWSB+NZboYnAx/Z8v3t2W7+hgsIZwSKMQALf3qdVFZUd
rMgNIv2qUVeeGNmGhScLUss8LqQjc/+Zdq9HOQ4ADWkjGIurNVOnA2ojNUcfsOL0
1tdHTfyuxDZb0WvN+VMPmuZcZGueuTtt+bTynLfw6Mltq72xhrZvEMbUriFruJ0t
7W7chVgOK4M8kL7tMZ5ZbNXPAipTiSgTykUEVmHLSPku0qxWGpPi6XVyneuDhdP/
Ip0DnyrKQ1cUQftLLDDQAjqGsbFZC397zQJwCL34TNuBQwE27mvuk+LtvKUjZSKx
I8+zBJi31GalgAiZ328b9WeJrA4OmhMdV2VBDuFAmvM0T7N3sGb9Ixrv0ksjMC0t
UHPv/wLu6rkbjA/o7zEvarA+wtV93cuUdBHM3Y5QLRBci+qx0b3EJ7iJBjGAXkBQ
EKxUG/gIPBFgGtahSkhvlwWmrsiMEwmquiHJqaSdoH/bpF+liJTk27D0A8v3NRmW
NNf+Ln7Nx1W7nBgh0Dup6tWRjEd9zjJBJUDcdcGlMzRPHSv90d4EQqcPkU+yfTxa
V+IfFRZkx8g+enKYVLw9MFNdL9G4Y44y0HwfiS6dEJ7vnbJ3CcKtuZ2cepdQUR1B
SEVqph9GPU1Pq0QWTUDvc8QDvPOz/t0hvattK3VQ351EsZGVT1TC8GGVEHprmtJV
4XfAKTHdK0TwoUR1ADNuEoUz1CcB80riXanOsAk5np749JenqDjx1U4QO37NLKcF
0Br62KYE+spAe0CcmZ4Z0WTT7X7TExR3L9BBrqV71Mg7ALj0PogsR1ESL3dw602L
dvzw47kUKBo3c+pL1sBwVRTLJ3vWS3sCNPMIs2fBz5Ssrcf6qWUP3h5Yj1DjOyni
0D5jtEDGw8IFt8fVF3PEXdKJBhj82zdlEki7NJDO8bKcBrcITlstX9qF+1bl9qF3
GyOE1IFUXVTnhoQOAVGuNBJWbfZjbuZ9BERShY51lTwCYbiMswjypyLHeyLYf3KX
zopB1QhoFbJxPYF4ywWuYEE/G8NmaBqrJGgwYnsQFIsju62UD5+Kc0Qj76etG8li
LaIGosLBtUxTOGNp3woYkOiGRb5JUzPDEbp4tMVeV98KqCBBo4EL0f8WvFM/fuT4
Kl8Yqxz4l9hqsKbxjTC5Tbm3F0IoSZ3GbT3d+/Ta16zlYxpUvZJrj96TyftJBzRY
YDTCXeb04j86pCjj9QLEUjvawJB4i3KR1z/bQGfTeip7XqcAjcDPTE4tPas8Zsut
DeP51PIcD1F86nEQgzWJ9jPl1kuxuI1N6K6RSqMzayJUwfdA38Oe4bmH2KAOwyN6
ctKZ7W2yX3ajuAMawYOHiAC9spKvU+1u4kX6LXVqc1pm5X6Enwdckoounqqdlm2m
wexsEhHyCDgAC3LXSxO2gjMLfu1+dddFAV2lbdQhNW2yyxjaQp2fcpHzrvgYha9x
uDCvL/XOHdsWY2MvmtpBDaBHiCZtXooEowyvgbDC6BiuKYOLlf6tYv/19b0Kdv9y
Ntpv/CdLB5l2zX5972X+rjGz1AS7GVcB5eTxygZY3kHfAOgvfu0GVv77L3mKgCDn
s4HGBYLWKSQJiye2egQLAoy7AZ3W+PiNgeJqMNdl46GPumMi8t3AlAHsDMZWyn1H
C3faPORLqcadz+sCFIVlbnaUzq5b7vjE797mJvBvzN8GztlV4M2EprIUfejZuNLR
bVtw9F5+A10BqaQFZoCemLRm9Hs3ezqib0YlyYnFj7vX1tajS+C7IihE2Nwt/dHI
xxm6Ia5ejSILvfURqLxd3TM6U64RtniZAKEfo2aYHvKbzAUmusNCx5tjlteZsr9B
98qbEsZFxMF6dF4VX490WZsfCYIi3P3X39iMr0bqO1NbeoIKzEohucMmkRhw8GWs
iQtClVMYUGUK0mSdi7u67P6I+vdvohTNilWlW0B9o7CkqnEwudoWm6pnYL3Nw0mI
AhPwf7cic5C0JfD6fvf+m97NyuXmkYxub4lo33eVgz7I+V4kP3ZDa8dEbLwO9VcB
GcOZg1aRXYZArv71jIj90QlFKOG4UfT4DX4BE9Pz+jxL0oY2hpnCIaSgzhkIKu2X
rECUc/HnoTrr7AOI6dh4TLcALMyyQuvODNrmgl72xnqGOtphfeW+nYDUV663ZSx3
2nv9HSRA6IoeZBLwjqtcwNKx5+ODuHEedq1cdJdOUFvXiVQ0ZJKqR0aNUNo7i5SM
hIiTKlmMNmDjiWcgSSWtKlwK3CWabVlBRWDX3ma6d8mhFiXPjI69qNR5JbqoRaIY
eDM4A42sNli47wEbkebQoVmf2nT+tl1maBez3j6UZtdEKbtyBbJPIhgDmE1e2c1/
yfOY5Y+xhjQFaeTb6gw3dx6sfdrMd/3gANlEaLFIE35m8l0a4FgpgrcJnkxtEYJe
A1VMLSKnSW36CGsSVJQA9GOaM4puSTcD1TNoNvCeduimRlwbbZIQHkPbmoEi6KHA
WuHlMiRw6V8kAY405E31bDHZWJX/hazfFHCkBoL+h7wgRxAV1qdkvMq+0zpWt0+q
tgAr/PWuVOsaJBBKuLzDgQb/BOyJw9rQXAtBnVWxVTXGawPiAR1tdicUckQ8wubJ
WyCRSCo6pBs0ValZip82BpK+W6DQprXaT8Fw4gOBprweIHQQjjAiVJHTChYgzOxq
ti7vY6TGVwPbNcYQ0FN6EhzvervIs1S2Cqjz3DFHp2M/83+HmyqEEOOgVKZYylWK
CAkyyqWiJocCsin92Otmw9eZ/wTnAkmligUK+XlaE+oE3VWE40kMe3witH2Jt1IW
hRZ8bebRwmPZYFJvQzp6WpRCRGrYlOYGMNEtpu7235Gr7GMqj83PAnt2MJcaud27
9wzbp2RwjhrrWCuW4QUN+uE6d2t4SWuaNpL3qSdDsswKsmEnesANwvajHs2DmN/H
Kud9R7V9Ic7nZmm2d5YmryOf8VMz7WkQa584grIkknTe7gLYohE3kLhrLHANSv5b
4YuQsiA/CA/HeQWr6BKY5+TYg3CMABiPAljrPua7MzwzikhI/c3rLZZ2CNbUlNOQ
HVxQWrl0lBSa9sEq5e1hX3iBtpGpnPt++CCTO6/q5DkL/nH1F8NBt6DXirfgtrCC
wdNB2spMjRm11Xxu4/OIi0V48nuQoUejNhYC3yv6IXL7hBHkgQ28Iqa/8FY5hZB3
khpRYSCh2mAJLFGpt0GfFcipJ6/02qcZeJDfqazGkM4FU1oeqYvqe6tvX2QYFVeo
o5zn+j8z8WLFy4klt+ZUnWnyRO/bOj7yFT5/Ou/7DbDo0pz4eyIViw9MCxEPDeYZ
CsJUCgUs+N867CWQmqfM51CPtoVMZc54TYrlNLvkeuJVeofsok7D3zBul6ZmadEv
vO7gHlIHTT8amqbzNqgyy61g813pmHnciVg9Ymhml63L7s5dq5N1dUyQLfmCzD5u
0Gsnwa95UpmsgEFQno5vezSjdfkRkHjcT9F+O1eeClPAkNl/QexvGXLumk04vFXM
oSe/z/T6KNA0XPiW3m5iGLNHwggT649EWG5NKIb4e1nVaZSBs239uXx6qq+oTWEi
wuxoHuWSMh47xnXe+u9UY3Rb688g116xnIYv0PPHJdXlgEiOBcTZ3YHZ6lh+s540
B3A6VWv87Ou5aheQUUokGFY6WAKH/HqMwbYYFkbVuOV0jKWG9+fvAwWR7k/LmKEv
6HpUULA5Oj2iVEyKRHIUC9AhztMzTsL5VPQUK5uCLk3wRzoPyPn4Po6ylqJ78sSw
sHLwlvTVWR0qZvUC2a9A5SwrTljn5xVV3Nm6DF3h2P/RLcsDKGtqza+A5mOtvv0b
Wu1xxCa/Iyy9TrYWIc3g8yO6TxTEvak6+JwPNlVZlRIWBQztVf6sLESEvcSKm4tR
85HSiQJ5xH1qV94+5IFYua81wuB7/3/8t66jb8EZUpGegD85HhQXs2K8mOmXb7YB
kjP33lPLB2FdALFXOBeGI6jHmVBNxc0L00/T8DNF73PSuXH4Kycd9n29ubQ7z/xU
syvQvBlr4Yt8X2/tDkz0gMLB6qH42vEuMnxVpZsUu76WSiEV8XlmnHHeFwpvLiq7
4vsd/ZerbBe1UrQUhiNqRcsaDJ87ds2H+Yijz0LzjGosf1Lal6SGswtH2E2TS5kt
51XwqNviXiuxHy0SP3CUdS3yMg74Mz4TZJGJvuLeKdf/B7MVcMKA4SGv0xouSvPW
RWVkqKDB+yXmBcLd36IT2U6XwOOxmbDDfykBQCMOVnsL5T5CQbdxgQiWQXGhcxao
5+F4/UFbkLGf70jPPQpu+6zRmSUWq/AWjAsH7k6mWmOBASw8a6jAB3HmoQAbX9Lg
LvgtUfire5jZvPxXyNWKCXEKEvesYqLx2Rm0QKgmz/k6NN3PnUjn1soiEke2o9uW
nWawPUn/JRUQkxhTHOGePizVGJCMTtaoka/3klLNL8chFgTxoun85At5STKSI9RI
IQTchAHmNYtCJEUiRne+VHaggLfr1seXOXqCGxIKWGL+RWzhHP+e62gB/Nq2lchy
gQe1KQC3UQdsbtf0Bn7bZBGytHSW7CnBD7XRaeshCr8tict1bStbjV8LTA1YQw0Z
aO4UJBKUORtg8ihZl4W1YoQL9GI1Ap38pmOxpNfOTbI0xhOWtAr+c5iAhDDztZ7t
QKw6dyAYaelwyGrlw7JHj9lAIHmgzrDy7KpA29lo4Gvk1SXOcuA1XIEzVOblV4MC
XJyj0Q7M/x2syMSkwOJsFnHmUOYcahs8WG5EQQgW60zVl1w6R3CCgtNMQRUidOfD
nR+PDrbsGPzh5kITPbIHwjvp+DsgOCJ/1l0yWLooRBMvYn7YULr7H9h5vxeNYUw/
Smo9r4UD+o/Q7v0jslKljAf5LXeZaw0H5IbNaXBFaGuIcHF5f1i5JaxHeBXb+aQb
nmWY4GGpBM/0smQKGpnb6HcEkXZHAwC+r02GTd6V0iGaU7yg8nd+dg2voeIGGoT9
Hk6vtjj9L60ql2DpDvNiR+rtknMFC8uUApBLLRDJvG8Ks0drZ964XkJUQv7wyhhw
stZCcgO8nuQ+O+q45HjFWZ86Sras8SnZupWSIFpSOQca2d2CkkAVy39en2pGkCd1
yXsDzsMJhA7L0adG15I4KoXRTGHmpsldRpG0Y76e+coO9JoWB00qztkqHDLNv3Wr
clswjM+KPsNjC4iU1XcdYzBgVEHEZxKyHPGsMYYZNawug+2V8tVYR0cVm55PKIWf
DpXJpWgUq+EkA17+h2fc3IzN7dx79b5/0YLi/AlVZToMtsEYLp74BoEH6OQoeqrn
QYqE7LWpllMgqW1ER2012OIgytIOBWuEcunpiHjLEvt6ZPCOHkfPT41wl3GPOAX4
9uD44xZl1o+kV6NekK3d35HXbk/eSHbheIEqJbJ4JwO3fDr1qUCj8nkE7V35wdKI
5RZQY6ur08/1iz4YKq6FHLaukA/OWIKaOeG/i7Vhtei+lU5l+uDhEYag2D4lkoKQ
kP4USc0sK9Xj/6uJqK+7f2v3D2TbnwfDBDwRsb45d89i+ahESQFD+MblgZsbORJw
1TO0hphywJXESXOCKHbHisXOsog236GmcBn7HFLSixUe0kVXnROi5IFnxFlJ/A5K
kLFpgwScV6B9LlZ0iEeNFLVHJmP87wxPkKOt8xiJL62i+SMJCUggDTI/ulOpzi+w
Rp8llrZnMUcBQ3z7M5TRyJ5I0gpQR/pA7n0Xv1+9ZWUyQhxKZh0OUHBCmgymJ8zy
1Zwedsqt9nQE9gWY2quZgx8TpIiJjJP1+U60icwQII2RrMOeRTOjq3/osJ67RK7C
VWxM7XoDvi624wJVZ1+tbDg2GIp0zrl5T0mrTmk3hGqzLNS7GgoU1Esdira9QFFH
UMpBkMrWMLNLRzTrCd2hx4L/2EgPSS8BA+kV7wy0K9Cvp7UVR4Wyvp/3s8uQ36KE
hDDUK62tPUufIHL+43pjvtYYH+d75kx71h9j+vz1IBq5kNh9q1VvLHuBxcNDcDeA
CtckkjNxNTF5Z0TNJuQ1WJTgRbSOUw9cyjtEzf02pgyXSBb2uwB0wIrjgj1zTEX2
7OX12F2+NO3n+Qu+2hC3EJHwO9TzHDfGWwXJhXnFx8CZ8fh/PGQUcXxnt/mJbgw6
Y5jzzTdMNYavpplLy52HgD+Wrzf2huULN7VumPxjHaTohVHEgolTMW5an3h3fVsh
ao8NEqO2MQpTCguGNNquXJUGjm5D0SBON3KzslUknnAObKB3pVeLtMF6GnYjl/l6
F8OgTxT8582KS3sfCBR1+kvOIgUctDwoEX/yDVhRhZl2jXYOq3MbfTItFSgQZrZr
sVYbosOUNVDgFb5kMxE5yq+a8fUH6uAGGxHq3FCE/sHKscfSRuaDU3Tvo65g8MJG
GOYVyJnIjtfgN6UTFXpFzWmG1ncCoFkYriRF6R+x0dV9FtlstHq5Rr7eUFN2IPLk
Uxt9nnbzcb3YjnyxzAywAoYT7x7Wb5rMUEYVnvK6oT5gIGEeKE5rD/uihV2CTtpQ
dRhvpjs1yZpRW/zG6R9OiyaRmYY8a7wQITY62LOaxcrUR09yK96+K4Jj+Gv1j5ST
hHEL+lvShE+QFp5H9jV1+Wa1JbBO35cZnIWeuHEDD5Dqq1GP1KfmdNv2c2yKdTE3
uFrDjLMPwc26eC8TjUrNGMJDzTUjanos7u+GnjbQpdbDupH8USfsXg+awdWXD6Wu
AOgYvydqN1O1+JVmYY+NFAEb42roDdMcIwGor6VAQXcSJSeVPC5QCYehr5d/+hMq
XUc6vrQsWkmBsEa8oJsBQADfa4hpPMvWsKuFVbQX4tcMg+P5lJ55YGeDF9yPp4pE
+oz0RDbVUkg73PEa2mZW6TLdzEyToFBEVhM7ttmrm66pyBdAZGwYyHtLKSjezFhX
oyLpv4p3KegGMnTchkLlV/wV27to0lRVAEs0l+j8pzWgeGAFVES52cNif4jUhtaS
Ds6WEz/AFkmIQdcbewofGzmOO6A6qJaVWyPVSs9ZC0stbjq0yPDSAIs+1ZzuCJhi
x9Qnn04lZ5jk+GhZhXIsqbmXRs0hMLRWvn2t0aeiawtdb2Eas36ESSAnbUxWIxeW
AZflxShjx2pVn0pdV/5EugzzPye7o7Ezmg57eY60aNiadoYons9h8T+CMZu33Pyo
Zr0NkBH/vazlTqotp4PM9FUF1ONuz7rs4g3WqyVTPHxky9BC7xSP4035mlSE9xEe
kVjPwfPDLX+oCLJkbP9vjwIOsxvNSOlt1jmSLT+9b8Jr8K3OiQhlYRlBHJe6tOJ3
EmHU+ZLvX6tRCd3Kr+ivC1HWdl4Xe+tX40xFEraFq7nwwGdP2sEB7hcMdEVWTHnG
VshpoyVkc5cPhosTZfUTJCNf4DUjYqj6Sup0N1tJWMwncFKMvxw7MqDu8uK5M/6e
EPBBWgacJ6JgVfjmf1dRXdaMaNkeqZcGdOI9bR3jpuS0zZP4dFF0q4k18rUqetuR
qqRwyVz7QWCZIlMOoNtSqdnWDjJ0d+7YcaWmPnphFiSZFKVGkNc3SmF42yEYEckf
i6An1v1ZXfzH/5Fh3AYYTialqWIjKry8uPWkXNAQYUaWeq1iNTGKPQexbNvNbZe1
H1A0jV7i4cmRz3dEW0IsMud9uxmfKv9U9DOGwe0ncJ/Jtc/BOHHBzllDxY6Ciu3v
7GMKL1m7heSQube+L90zhOxJLp1SdtI6ZMbNQTWXKWAjpIwFQT+oF2OYMFkpWzSL
YbTFD6QcvHEm/y0VgQCWNP7VXofOfDwrLP6gbtx3NLqbF47Ng+zEeRbod41GIrx8
EvDShHR9Lt3NEj7iS9FD+Fw6fWvQHwx7nsYXX9IJI6oTaWJueGX0Xi6yCtJGS0m7
XcIRs9SmFc6+xbDQxW0DCVYAXb7q5cGRa7DyDYdy1x0dDuFaX/UMUzCMoWgr8lJf
MKFl6ZAy857jmGTif8rBVEKZ7/jklrkWeJdy0JkDhzckuebZIiuAnIi/2r3YxvPt
8i8BioIu352qL7Rwu80Yb/juW0a9Dlim6z4chw+3edesE6j4CxR4u9hj07eGCKTW
vcSff4WLkD+1BNXf3Gy926VUY6jN6v7jsaa3QCD/1JYd+zeqt8HeFC1tIlSNRhoK
zkXg0b6pge8fjo2F61guaf6FC/42dciXpHdXwlmlXveEk0OsWIPpopGM2juIhGDs
qKTlm0NFiXGrNp+rfQAMZdy2wDykpc8KzjCqG9JwORA7TA2IZqTB3wJDeqycN6Rt
DQJZE37tBbYW8qmnGX6oK+iz5QVNSfPgYtoreD7OjccMfKX1M1SDZfFOtbOo14tX
8tU0z12032Fh1tNv8VHtzFgQ//HczmHSqPqQxDoBvjbLddzo+Z9cAxkVhAcnaEMw
AMWguf/7rBcr8R0ET5GAPEP+5AWzruMrTMmPtYid3bT8YS7NaZcvGj4TEd7JNWhc
X1WsQAZWgi8o0XC9CvRW8qDym7/n1zmm6eKosFdC/pUe56W6p3mKOojy9YWDH7yB
Z/mXJi//VyiePKXm3PKfMAuYALZdNnF0zk7tNi2D7mBKCvNq/EDwzlTZVUh8nXFL
b8xndWBrvyQ/dFINLPgrIUs+TrsjylpGWkvWTa7bcQ4i7it9dA7xc7a84qsgC8vt
3yfRV8hGg/yyBv89v9XjZJysMSreZRREonF+Ryw8/0RhzxmEpGxp6iQIyJwffFhq
V5F+1tRpGdo8Cex6cvf0KaKoTWEeWaALUwCfmIeouFU8gjbMlGZZ0lNYvRqVMMes
25ev87Tx5yKwDVZeh5XAm1ZFhX8RSdN6cbmoWvgSqmVbyEbGsLkMc0rKhZYdvCw3
hlytSDqkQRJjVT7LBlHHKsEcNezGMbSALeVxh101NYMHi51Ngr1rDcMQFWIX4FWj
RRnrQ90yePlPp8EwaJY7sAxxMMs4+GlDfkKmeyZIfBHDfFw4e5fBF/wwDRYGGjAr
RljsMl0X+l/trxSVysTjTfkN1vABlA0jmB3lZYSYPOMRSgn3CdViF6HjVsbSO8tS
ydYUee40s9pNiIMDm457yoi6b1WMYpMS6GUEazPq0HYVSTQgTj2pF87OFDOa8QdO
fwuWUYI1TIqtt41sywwbRQkD5OK0jU9vIXJUEnms0IeBEziL4TZ/LUHnBlGZNOVm
Gooa8NJ9PTP1Cis/fUQCs3kCs7xLDpEFrJU5Cko9PlMfop9HPQ8LJPGh5VmC79cC
6Z+pCTNywuwbONg2XZZ35L003qOvmsWjkMscYoICs+2MnpTWnbbZQi+a1vBwTNHI
clhi2Zk5iqaEe1mzOrgKoWxUHaG3T7f3njg5hWFfeuAVuHDouvVvyUi/iEM+M/+l
BEUWwtXDNHh3IGS0QjR+m7DvECo5OxVMjFvJPPJIwTzpYHbM1rAPcM9y0b/d92vq
gH1C6S4B+4rdBGrYXvx04lIx03dA/W1CJKsjEBb36ZOz75bd2StmAiy3ckL4JUcH
XLFb8wJJ0kbgevGOBRIFm1j6Wff6+6I1dHfDbj2evHUEvowsV/AuNYRqNgKkEciy
LJ5Xw2852ZIxCn+OY412lGmPbnLYMz1xX3eJgIhTx8V2jpaGEdDXFm1ukQwuUvNc
fo2PKjIGmZEI50kXiVvb6AafgKFU7Yw/nzsyXiIAsMXmUMXb/fAj7m1Ho2TsAIth
XXCff/ksAkz0+QtILK1uunpPZ2ZXIlin4burXM/XpsnJYqzsAK/8sdAd0B7mfkH3
cIzOUGqtn9JIU4qlA7gbcHJIk3yQNtCCbn8HtuSo2/rSloIEJ2c1bqpnv5Q7Wrf2
zbERFDq0Xcxljwtkj8j1V4m4VsBMOZT7+2WJHjBpJEavi9OAm7KGA38KxGZJao86
iU/O7vT2gV/8Ypoc9jIwEEGUl2zyiXpA6GFYWXFV13KfoVVy/xV1Y+EB58dGdfew
EBdsZMcAPYS2hxz/A/GaNwSxdweC+PndkE7+kpBELGLFrfhKVVhTYgY8LMncYnGR
RzsaRWo0ya+NIiCwIGIGfZ34NI/nKQ4zzESOI3GOEvVO7RB4IqgnatUJgnf2NqTX
Z6y4ThNWguDjHGo1lwbC2bvRvjcOoRN9KCsfAYt8kFGwABJ6Tt7e5XWPkwt/I9Kq
k5bGMUl1tJz5+fkjM+doR8hRapXFBFnyX6JhEYS5Y45YOhrdadoxeLsyt7Sh+rVR
fY7KoalSDu8TdJfZpRhXPvRnzp7m+B8RSL/4Lla2rj1OBsHI2qTC9cFay8oeF/63
z07LoVrjmCr8qWtI3k2/26S42bkaT0DVCQUEjts2Gp361sLeOPzM08h0k2CiL8pe
zID0c0mYzVTXVZ3PmMR/Xcz1+NgQBhb9wwBz8Yc3pc2VIQVkqICF/PQb+GbNYP1e
9lruvnzX95SHMS4Vj90zxCVbYBpCkKVAFfEvLCy9LCmpWIPSd7RnWNlMmXfLfRLF
FLg3tFqvzutyNV6sOvhxOMf0AXFl8DFDfCW5iQfmpgbOlIR6AQKqZFY0Ngcjx/K4
IoeN45AIwjNtYwX4gWGmTh6i7IPimu8vpifxJYZ+RoHsnHBEqbg/E1aIuNjX6WzV
3h7bsujESevm5RM5FrUiGgXu5dbReJZGuo02QZzcdonoCndLJOu8zm+aYYDYAH51
VrIDSQuzbnCsGSW+49AjVv3tljtkUY1AaT9htFWL+lzo396WTzsPBfaGYR5tr4+n
r6JKm0Zjzn0XTCdks+vLYn6BkLIhOHPJmRzjB9l9J0zum4jxPGcvIeTm4zIRJB+/
ifm2uo1JjheU7R5ARq+EV6w0gp1DZpCT66q6VohxZTX5IqK1RZJaY7SMkGf26O6l
nVeQofuIts2R3eWbjg66eFGs2xNSx+nI/KmHr2YfYA/jgNgcgd5j9gxpO/dybI3w
OQxuefy6C+xmPxPGgQex+4+pZGGACHzxFSAcuHjP8NB/QXtKtotSb9p4QGBm4vcf
prHtLSuPmUZ8KgwX2su3Yge6b6igeTE82kha8jnp26K5LqDgm7mUeKqGjOLF0uvR
QChG+N6jEbmBaXzelHMBGElM0k0XI6s7N0XVaSKiTk5TSejKC7fm3wkS21ulepi7
P5v+dMB9Rm27rurtxstUtwK8hxi+U+qKo48yG7gq6TipoeO3/2MoqUm5MR4f06Gv
PsblAM0NBxOPf45xtdDP2nVxyPuYbKR12CI54jcNBcuxbjnADWfQ1LujKrl353P8
3J6MdKn4D/Pd9wT4TdqKUxNKlQ0yU3AE6WDEcwMoa1WOl8tKRfUCoTdITJ3W7ZPa
vFBIp7EqdWshxAxY2dgyqjH7I8/YtBonpkfRQvcBFtjQcuG4+sx/RvV4/fOuWN2O
TRjpU+6uIOmwuJl44zK4y2x3/eiKh9Y7LM3ETG+i7g5fvmJj+PYn05CpxdGZUEK7
3VcQmnu9Olw87Ytj2QxzLpE99/Yigz9GrAeabc7tPyh6byhs+YVUJIEaJ3e1BOvC
k1BDuX85kH3Hfd0G5Mywldk3qPt1dt1J+rNFH2OtG3MOlk8zDDCNBnB5n5e1gqcv
aZCIs4Y3xXz8ndt/k49pz19/soogwuOoltw8/K1l6BuJPLl1EHmkZ4s6thlvFeSx
LWB6luN22FulEUaMALOw/ISvDvVCFls4MbsMSVi5hYaImD5BotBimsgbJllLqvpD
RDCeQwCX1MOun/m8/OH3xmAjMXdDgzD+Hq/gNCWO92u5wWNKU60WwHfJ/tJu2vvK
tVrdv9pcO5ANwZCCf5qHsjz0GtOJzKuXttwnRctEKG+sCgqLfao05Swg4eYZxT9C
FjlAMwT3VJWDPFLIMxHWwRjNP9XkAFtS9Qc2o/ByK9h/ICpcwA3m0TH3+LgbBSXC
lGQoAom5Nn16Sy6GhBxLP4RMNSy/1N57TEPfFPywecF529BamvP1iip2kXBIfEoQ
rxwprLExe1FfxGNlnH9s3YzLqkul9F6tF5PQz5h7raOBS3fnpMSQRwrBMFzDBsap
QUcSfuFeA5Vzz5VdWYuc4l8zEUXv6l3PH474dsjLxgI/p1+/mbYze1VLGFF2VSWx
I69pSp5FrdYA+ktcm75E/i3gAo62x0bnPIwO1jxqNHfTbl6/0K77rDh7AvGWsDTK
tN7DqexYDFFLpiA1aZReHfNS6N8hJJHwLOzNAgKTVXQ0EWbuZgWAP/XPiDrDvqSb
u2wN8CdHogfRCINmdxtdLcmnYaCoOIrFXTNy/zFM7dESy+ay1UMBgnfC+F8EwaqX
mbEO5ndkpUqFe4Vx8jlv0KC9xl6j9TJXK/HeCq16GuxPBcK0LUrKyHRik9lcGapu
GXrlRWscgkZRqOnEjzXrmCn6U37UgAJ6cMhZ5smCefr3c66G0f+hydtVYpKUKvRE
ngalJqbKZHQmRwjSK/VvD3WYCl0VLOdTlm9qDUywZM615uVR04GcRD64ZLe1s22c
NstcrdB9eaN0XPEU8oLsZKtb87VkvqgSUYvpvHbITDkaeJSmWDnFS6gdnARXec2x
uelpIVRtQDSoztfpogm8Qgw181h1UMtrDwjDkNKHMM1ypl4+oE4Mr6LxZxHQjFcl
TxqJ09FrvmZLeL5lLSF9szTCnxuol44URw6YjAN2lNKy7CvmuBOIK5i7OLpaybBp
YHWxJF5NTQdh/OK49wWpChFTyvEbdvMq7rUuo/GN1UU2rfbQ4ErYEsUIjKLy2nm5
I7TeTMNOBDLPFu91EIqit6//kYDonwIyOdok8WEZepPR48gNdoiFRWNh1e8pdTiB
kH/jGa1M3U5bbgKSr3UsMuCNG65wC+L7rQlATP5Qgil2KVy+oNA8XVEykhZk9bP/
XiloGrDwVzB+q+H4GPONdv0fUnytwM3ZqE2+DgO8hh59O4DE1FbmZPMzivaxWOX+
PtmrcWLvDwq2XW8ZumM5DeO/t1BWnZ7dAuuIPmGPVgBxnp1v5nsQjghOS+QnFLkh
8x2Qw7cIxXoQHrK4UWap9C5pkHEN1AdOphYvC+wsBNvAznD3HtlsstJlt03YDAgL
lDovEvHGdnxRBjKgFqSnsKsE1dsCnWU9dzXSVn1tNCtY0VouhaoCM98QmgJNOIQ9
0NShtd+uONaOMCcl/HEVyRg2pxhWLl5t0bJ1Akdk6zYHAMr2W0RI/Tm5l5DGADsD
8fHTniNMwXTfkUD1RIztXqN/Lpz452RtWoMlaWGzckCVAb4KLEsAbMJD1WY0ZKk4
XXXdMJUOBZ7LFeT2GR7xrtvCLsZLAcpNot+M2AhNfN5Yz5RHRjEtTittg6IM7Onb
qr2HxXq0zC+5tR6f5G/hbM80A8TMo+nxDlBDBmD0L2b43IFasFS4rw7vChMGIZEi
kamEbekhcp62QblkI+81C9DjB+IW4AvAu96WHyN+nStDc3/h/dBkgsZLHh+zA5wN
Inv39OIpz7EbNauIZPePy2NX33qsrCwEpJmNWYQ8GnGeq+Urcwxis01R0NIDETn5
iNGKIKmv3i5cEIK5wttMqgN9S8fwAmMbeuy8XI/deUZKM8t5fROe5g34+AvEs1Z1
8L4BL/u3lXKvMXTlt4xXIcLC0o7cO7y/pk4ARnGo9CkAQXbrPBRMsQPvAwFSy/FG
9oC5PDxka1RJtNkRPB6rCeY8crvdT2NycyL3VBK1NwNz+w9IlfCgkq/FdE+FFhbu
Dv6AWIM/tyVcSc+skbC1uhRgdAKzauZuI9ENtz0Ny9hLjpezpGadKRRqWRXc/5zM
rHqMVKUJLGsA2UoUL+wcrPy+21xU/uzFgdsEHcNFgzv3S//Ng4Y2zrHijzpA57ba
GjWMEJedxtv3g9v+FQxLvKWyE19/u/JAcomVoJYtsOUVaXuLSKYI9uUD5SajSchu
be/3e1RG0PkUGykh3qDeW11nXbw0s/XJ1hpgiylRLF5tw+wzXXeCN1wwkgpHExo8
2cZXAmQQj/WLRHa1hScHdAQCkHE1ffQRZ4w74FVz5U4IA5tUBVXSvk2sjl0v3cov
XmCe0BWVnCRRS8IVFpJ+mSU2nNBxIOLOrnGwA5uPvYrIt+O/OrxNhtEA9maOu+s1
ZConDmVP6g3ypOot4oRi7MLUoqU6pEuT6LAkBEceuLgAlK5j9PLh6BvtSg8Zu3HN
K8pCS6YGVPDRXOCmI6lnGr/i71UY4sthx3I34h5r+PEWxFJOLaGKLwcVpSkEcQ6P
njuSydeIdj71wt8aNXabbUePup2tk0kIqbOTd9RfJXNef1iNHV0hKQyicABPKhSk
O7bGY9yfNugNbDcchiYxk5P0156F1nvCVWhDJ83YAk4Jq1yDLhvOSsLgrlksZXRR
rxBrV+EkhVLkllR1jm40YEQ0ldga9dldGnbJ8RVC7TPLRy2XsHhj9WGFgHMK9J/k
sjhXoRhz8wj/zdokxS0wByV/mzVZIHp+Payi0/sKx0EMcJm+FzCDtUK92JkIkze0
lIj9DvhEEw+zon8gblBZ+JzqB9QXsY4a6A9O6QUq+KlMRe4dA3L46aXPK8kviAVM
FvCWcxtgAYvU2l01GUnSadPnBqqNURphspE1n03TvcVNhczUS36ZvAAB+C2/ZTpM
ZcIfsz8nB/XpoDfolPjGmtsqxuyYSK7oUSBU6IHAtBYh3i7adtVPI9Nk10eCl2q+
Ik/jkQSVTb3AZcMMTsEH7rlTUzr9MTWv3xfKCqHa/bp/nCpG3Aswvbflb2ixGMxC
vuyqQYeFyROxV5Kwk7G+WK4bzIUCEFtcVUK8ubXJCsraVoHba5TPpHBLpQEdj0/B
+KECI0d+UA5IBzFgoPYalqIHaea2Tt6sWAhw1A0dOrzodf5QOpeSJ0yWficE2u25
aHQYQ+u+cUOcOoD5WDTG4zACJLt7Qhe1n+IXi3AXDshNv8SHZGlvmRzrPpgyaswZ
+FDMYX11DdDKK1pI35WIULfpIvqpuE+GqpGsOb6yQj+4CzpntvXsjAW80E/9L5p4
FXygmmlRqafpREpt3Qa+Hbzmkz/q7PzCzLTdYZzn4/7nPw/DnLQr6l8x5fsotsF+
N9WxgBdBQb+TmRTa+M7SNmBvY51vMGcUqERJyTcs0638l3axQkA9MERihgVC6E9O
Inu+Vk1QZcsmj1S0N5iLv7/Hy+xCuL6rJZZ7F8x2IS3omeeb+cmG19L4sg6mT5s1
IsVM0NddiSqCXlirui/bwuV/pW3JbDg0enqKdEzP5yMx9BuFDiql4QiZ9T7HJD8G
g2dZ/ZUqHwSG21U9k5upX8sK+aiLVP+FlUnJ1vOEeXVhiEb7FMExbuVu2/EA2q9g
Q8M6dirANaUL6BdxLjTZW7x7vvsMSuiITcf7d2YwWp/PnDWSseNRXYsYSThPEkaG
3RPqKiqaZ7c5Aq/gN19TcvKkOOLmdlerP7HYM2LkiCBsJzZXfSHw9q0BmL2gmuV+
UjzXafN8dItoZYB1nkM6nknerbXx3j77ZrpDX7RFJrhq5V5CTCetwcMXLE8UkQOn
xdygXIMSA8718Sk0oHaDFEkWtNG57yqVJLPayP3IwHHK5skHokHV6XqyRqvE5fee
UroAjChJVDO/6r7RJXQP3qcX4N76K12RxEdo2Jd3zfOwApnpMnoN0i4bR9nxrAB6
Ydl1hFiUNI8tFKZ6yMU7L00uceT1OxMva9fHsKwqYIUiKX0YVPFWx4YCnxKfNm1i
BWbebubv8HCKAeJ/iY7UrLh7HxNkKZ76pEjYUcBRBY2aseR8jS/zy0cHfUQFy8mU
20Qd9pLGc18/7E/PEmuRUqyMLSBqDxLm4srPIHBaIDT4X+RSIfwtyr0nCvdkF+0y
qHMih6+VQcq48ewqJaHBZ0G2fCOERogSA6AVa05+J78Gktdglu+zQHGBPlYDqKi7
BtlphfLNQVGCmaHYzzJm4s0zhw1OezUc/GrvkQgtPihkFUp7DYgP0VJMQ3bYvQ4i
0q16yQN5tnLsWn7GAfpA2sAnhi7P2DYTIocAW7tQpzjCQy7RWO7LAS2e0uSuyUYh
4SjniIrD85nS1mg7IgPYHdc4xiWjg1hQeEnR8XvTumk1ZCSRxnNHPbLQxwGnlpFC
YaILDwVLCEvOtil++JOugFS3E7B9kG54YQlvMWt0Jzg+c/HpIy0qnR0z6Ja5/GzW
uTPjCJ5bJaCs4dl13IKdhgM+kIU9nCpKJwN8Z6aMa71lf5DOOBdkSx16S7LgLmgb
Sn1TTLlHn67T7rAL9sHrWQp5TsSCFSNHl+mnpj8U3ao3WWtBeE6pXuqQbstjuINn
jeFIGLylRyZh8e+SSBUMeXEC7GrRqww1f8TvNeTNRrqRmCSn+YyRuYVS3LOOMOTj
1xG3UbTVl0IOkxkFcBc4bfzj5hkRQF7dP05u2mxmEQUEi00vqU+KEvZvX5z5pD3X
XYA7baJ60ii3eGrRVla28k+fabTeOTeV2+Sm4CFk0HMDhCwo/66/tJzpYJT5d3D8
qX0HVg6r/V+0C/cV15stfjM4loizHZOedtXuPHBFeJ6P6tpIWu5OUnt3eW6raj4x
9sgg5wY4FpCwoxy3l7QMWH6hT3FW+lUT7cGLLAeeOMi7yaQI7s8grjduzmjfL918
eu2FeEX/Nj1iG4irLPVija2fWudUA56t2VxBSgJAR8SDT1zyNDPSzAB9rdE6kHTw
yEQruLoFmwaGRy0DX9s6kh3HpvumnCMHE21RAh5zoiv4ETJoIROePjH9e+G7/0bB
4HZzi2Sn2eXiIM2BUcVGHCtKPliW7uhb24Ggtb3/ptP4xtNJd4UtJurM2h2M9fjD
QjuY4Bt/hHw7NiMSSRsfQOQOfi+MHLaba/ZjefeV+DiwXe+IVXV/qoKCBIXWTZJm
oZtm6ZVY664bqWUkzrFQK2oEY9BiZT24W5H7v+2zngl2ZKbHtRfzx/4wTpEgXVoB
NM7XQf+shYqkpv2JGJPsHNCw6wgeYremIbeFKtLDVL/P+TcYkmexH6a2KsLbgA/h
j91uUGGoXg2NPpirZnTbgvr0fj5+Sxm/oCt/aV3ppclaxGt7fGTGO10tj5KbMihh
Jw9GCaESrjaD0p7ZhthKSVEFuDtcWiZNmIcJOnytNyfrmf7buFN+qayFwqfETQST
Mt17+/t1p17HOJPJFA3V3QYHUy0pl3SBFv/bNKLp2JMRGrzpHwLQhTYdaNb6D1a/
bv7l+gAhWrQJd4y0iikgU7smjwHL0JYryQRP1LaxFehZ+38XNjTccW6B3r987fLn
JorTA6+JLHJLsa2vO9Au37D+uicP1jLamIyDyNztbkoJ0B4de62DkiLtsXK1tnK2
NfpA2lnfJ+8xPEQ012JnTj6mbikEXteJXHdpxLofG3JJFp6fe/Y5F9q7BfrQrq+G
FSBpkjr7lxCej8EEmvJv0DiZz3r0Inj362NxRCQkLCB9fVpEN+AU144EkxQkiokY
fmzKdd8T8X+q/EmgSB40gxBeMm2Of7PwTpMzC3K3Fa/ZZDy5vsAv/a/XSTsWtK/t
45Izvt5NC+HbMjwXIaBw378oImMWyZG7+U5nqRQYg3HTyBwZijgl0MyDDtp/FbOb
WrmFxALfAOw1YPcjOaw0N2XewJtuvM+NWSWMo10Up2ORydBrx4+UkDnW345rI7hi
CahlutKTg932gnIgTHFDcd3edCidMghaUrkEK3/4CZdPpVgXQ1k/WlrwvoLoauYj
le5T8I40ZyXVd+Yt8aJRzXpUC0PW0JpXRrnDPXNCwWgEPu03gfncB3UQDXqgg4C+
rIpnc5fusOCSZoE3/eCP6/EF3JUuQiPOegQ3Skh6n3v+k2sPQ8dLu6N2zlZYEib7
oAkzVppYzNn2Hdcsu/YSiULWZUy26iG0Xe3e+0wwlrH4RuUlf9gbCx8Yk64qFrOL
MAtolIge4Ecp51t8sGCiF/8HdPkIK7GBsqa7/7tQ7ptqeESE+DR9gifneBSZzPkI
y48zvOTBFlplhl4QZf8E0CVLvoDMhwOu8NOFWMvpydBSNM5dEVK0P4oig/QA1y3m
VQPh+PWwnHOEJknDIwPTQg0+Nt7K0lOUV/FiwiZLS9QkKagrCSIkTZR1QsNYGukI
5tnrYdzDdOnypdmSNlOqt49KbIrSKW4oeCZBVV2IHH6tR9mLUQnXdMTIEVkOxVD2
n7i3xrr970sbASDAVcwihEVsgZo89yc7V5JFPyMeBem2F6sstdH+SP3sYrg5kOOz
3y7RLrmfDfqBu8EOu3eTIXi/W/jxhEKAEVJeMxRJ1iIahTnkxEl3MDNj6k9WVGKL
vFv62wVF0Q4Ke+MuTbT5YKm3lf57wSv3HF+BQMGXAzlmldD5B4M4rpvEfD6KP/qY
G6nUEpmON5fKAiHVmqUYUtY6g798yItnrxKz/uzBB/DFEtQKYHhioqdoH+/a2EfV
cZ5G+oHwFiyXOdqbRQMuF28GOP5IxOhvVJHvwe+z3W8GjCevr7Cp44oeASRCvPva
bfz1u/ROoyXSzjbvkiIWd0w3YMEFmB0ox8b/TW9Wj22etaLOywcGrUUd+RtU0qzS
kbcK6+L3WXjppUbw3saVkHypUVltcCQXN+vVQ8Z0OSyMehd8My23Zys3u+rzWzz0
FUsQJxS3vTxNwGswwNjnfw==
`protect END_PROTECTED