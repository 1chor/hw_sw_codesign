-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
oa/GlL2zBaKJftExQV/KwPuElAkE087D9fLBb0JQnQcAXWjcvB8b8LsaRLeZQr4u
YixPTN7cYHbUUog+RnOMsztKpys5HdMtJWKLdB3ajVGFz4u4jwmF+JK/U0cpzWwi
nbQnIM6Vl4GHrOAcKGe8YVR8K/bwlc8o7Fnf0D+SRk0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10308)

`protect DATA_BLOCK
yWyYGfZOtcUOUKcnCQ8K7H0F+vEeypmhGPxHp9kbXdMAgu66T/ZgCfTtWMZUdjDo
yT1hVldja5vMf+UE34nLT3FojA9F7mYdMpfkkKopLwrh/dzMLweDbdcjL+tcAWij
2q2Z62ugfM0hnv/t6ijddP/R9yJu3vezZDNS4JEORRQ+Duo0F3lF3t4uGxz71Kkx
qJNNi/eBjKayX/oRuk57YmcoAUS/djFBXof9Wu6WP/MXqd1Qt3vRx+9ET7ngjNMq
XC8HvMDna5F6KSIkjLoEr+RBgMF4uI10WaBk0kPWr2fX6eDad0aMD4hm6UJq8cf2
V0yCeFHswElM0IknmSMVUMI6DIyjFnQyYbqE6Lg49hEJPb7QW3Jfvrzn+ncpw/fr
Je1t14ajrqNv7v1kQHJg5uMvGwoNHZ0I+/oryIwIJuYh5ur3lI8mfgZKH5nZOEk9
N/0vcqVF1V13IWynoNMHCrjC1TT8s0aQ3U3LmClVXzI7bdF4DT4RIZM2TZhHHNAa
ol15Xc201NWHBerjhEovEzv8XTdMdhKM3Eotirwudchq7LqWGN9Lcy4D98g7zaxn
qWkjdABcdF3ZMsWfci1sGeFWQOO9bGldzU+1IuQApwMOMjD63Df8OkcBuPfLNyws
t1NZDKptGkodK7s/qTXA3ccY5fF+OokvpBQaGNGggkMkuXGqffoj9WVKWR2zm2sE
Z0Lh5SD0BdNC2qR3G0X0GRpdP9l9oC+mRwRu+W9RuWg0tejECJv3CafV/FaS0Fja
opg+vbIoC6bbBaU+Jkl09aeDE1XhVhcVFqX9ScvK/Zkex9aKHa36gBRLSyIaAYrV
mafhs/mR1nDK1d3X9BcUSJZ/0MROJdbmvmu/+o61RRc4XysGwY7dRhjbqU7iEWpz
VGBZ9GuF6dRLtgqulDCKObvgHdvR6aKUTTW3sQwzha53KcnEzGDILD27uXI1gAYK
I6KiqNZUIk0V4Hbx722P0F+0eCh1msbJFkeMGTtuDXpZ7HCrmGwDzXUiio19KohK
7dIGjzWY4isB2d2eiXVkVs6g5H1Oq5j5OtpWewWGLPkp4drAQNqajcy8WwH0JAjy
LGOBWVUoBjO6JIhCi7fNwAHa5vjG4pdy05ZSwJrrJROJ9LAgkCoz0X9sdWxFFnog
ASdby71iElha8PgAaIZgA/qUs9Ag+zON6oqQt10jB2v+QmCTkcZDQoyNF01ZDoGQ
Cg3hfTD93ojmey8aEiKHua0Mym8Uppbkau2ASYjbr1fn8J5xcDH8S/dMInfMjCmG
U703sNJGBkfdaMvBJmJ3UdQazJX7WklYOn/cDVeJUaTHWEqsbI6OvptcN7TEACw4
7ZSnzNO0J3c1pbTwBZR0k7sgtjD8k0+vQV1i5j9WQRACj66pc5pSngeCrhafYz4M
5smogysOsRmiSqpphLuR72xRd7r8Gr89wbMA1RBJzXcZirpKESSsEvr6glHX7asZ
ASPvf62jONXNCFKm/jGMclkK8ZScdT1aBoYclW4F2ZlS2PHwwqf2vpfizwaJ5NN6
HC47lJDrM8tcfaEUG69wkPiYQxDavb8Llxxr0kp1rf8gDVd0y1W6E5zBOwZWnP8C
pTf+y3zfCmtW2wVbpHHax/uL2jNr1QEozb7o1zNHvpmu5opqLJNsxd4vHCQzrFlx
skjlvr5+XOHExmqGced/SB/eihyjM43ZyvSKwUrmf4XaGqnfdbImWdPqA2RJpjhD
W8cZWfcEcsEXzxs9/B0J98U+n8Hyq3T4zAdf2U7w7TWzMp3SyOnSdRpRXt/CKqsL
QYz9zrwmdhkQ5QQMMEusAmrgMdZcYv9BeFQEvmlR6ZejQirs7ZrFyv8tLLYjFU18
gcmzcE0rxADTCDd4ig4+q1m2Qc+U25PJ+M3/27bRZxPFXb/fUvAZeLsUMFZtX/8r
IFA4PuWjpMGdu+Rx7I6iZOcGiIQ1wk3y5p7BnSFNHbPkpTaQ6U2Jj44//+E2oOYL
+fczXgcEyYPl1PkTm/PledGa0XFPRxk3uHmlC/OdsfvadN7tOqqXF/fLGnO9Q/uu
Hgu+ZgJUHGsyjgGWVqsr5tH7dribf+aaBShFO5cyPLZgfZFVCQ51EpXAqGFreXoF
R/EPdyN6M4M0uCoEx5OTtDbmqlNbxmJXe77Up6z/sAzlw9BBxfnQI/PECFIiKJ8b
myxkiKqQmiKG2zdjFaNO5csqVoZbo1YWIBCwZFqqFteARPTbkEeR6wErrVU2nnt3
9YGaiZFMq5/K5+TTI6fMKgIDsG7Ejc9cBaizPatsaMlFsOM/TBGPxsUejLlJW314
rmi2gxQ3j63Rgbw31AMFTwa2Le7nnL7d0gxeN2NvE413hUxXn5gOPD9ZjDsW9PHr
PDoDuVeNXI0d5yFMD9DZC7a0XCTVpYH/T540RE+aMV2faGZr0rkC6Cuy8coPaG8L
lLKdjORtoqHxTcvBhDP+OfltKOi3iAfiQ09duSG0HyPA/01QHJJbYYgh4X5hbwmF
CKLsdMZHw579vj3oXVRoz5ezXBu5yTyWD/ZDjeSPKVirbdngFdwFZALGKs9VW6o9
lFveCUJbylxYfSR/fNMSCKq8u/h77f9mURzSVjS8xXcq1qI10qVbBtVtLDCm3K3m
2RzRUDmogVBpgiXzIqpruelpbSjFwzYkG7cibSqb/rhkJEfwWWcRxURutVkMALQG
nJyYl/rXQkywJCrh9TBlNzAs8exRr2Rd7/+qSrcH5Zyoy67BI75z4pG8u+pIJV85
V2kA3rszI7KROGNGSGlsKFFPmy3tOBeP3PIruv7mK7LrBxq2tTzAyre91YnDJ8yu
9aidwYVvsVbtxat0btWPNtlFHDFU6uCxx9AJTWu2IXaZ9oCfz9/8weslQ1vyiX9k
r8PZ5/pELNQeuH7oZ455dE45OmCctRvLxIXgVRwyTbkRC+YZz2Wzvf87v22tQzcq
p/l7xHJLmXS2bqdSLZRLBZB0NIcPj5nq3nlO0GZHPlgNx1MV+t/L50H7z5IaOKKG
oez/aylLG35PcFXyf2+ZU+aiIJ5RCZbnSVgFx8Ip0ur8yNpxzvy266OMZ3vCu5R4
zViiyPagovNrTOW0m2D9luVcb+1cuS16u7DrtZilCoPHeFOXahhslLjfgGtyMMQx
5f25z8JqehFTzfADAHfetq0DENzcTjzwpZiG9R2CsBnOpCEBLGXbl2rJgetpORVQ
+UbxZIUhLQEQN4uzmbIUwcEqALt1LZJ2JxFBH0xUWp8dtonX5TUknUY3c/kmussi
v7XmSXFUKD7Xn6oB3Y+WNM80iV2WKICm7iSCl4AjQ9G78OfE+EWp5Seu+pDrpTrg
yTRVW0wzrYoVbVvcG+0v+xzRbgVEa6te/2OLwXG614l+t1JoHFxF5tr++Wzgq4aq
5EZp6XNRv+QGHlEnhJmc3DglmTCIHDRaqadMsw912Kao5cWnJ6Oe0PRz2fhfpbxy
VI9SRGqOty4pXt66OoVAiNj+3yL0w9PB36bsECkjR+zdHETGYyYR+ZW4Wp+FGLd/
bf/mJNjeugOT9LCeDy8sXld+T/EXdHM5zvfOaRAwVJyYgExUPI0WjsrTq1FGwNlJ
QkkrvgHZX5CNJ+5Hk8PuhWOVIk5j68y6Rjz5/M/O+kgnOCvMyqMf6Za6gW5W6VUb
OQMDnDVFKSr7bqtn56Jf0+raGVMiVCoki0A5LHKW5vTEzCpgCrcsdXM7Krjk5pbP
ItzBl2jpHBsbOSYhDOOwSLBtEDplxxKlhJE7qCURMRficgNvNA83gt6YqX3BEOHz
cTPTY9pk/e/a1DsIdW4H1yKneOKqPFjiWKpHbsftpyNk+/oHQlF7N1rAOGXPTWNv
9RFNz/1TEkAYzDARETVQmj3hIy/O+FOaNDrMCm/J6CG5IwXCrgbNrdLB7KzB5lYC
5WNHwqlQpFCwNka0z818xMXSymOsEnNAWaKEDJWht6B8wej5V4VKV+Wm7MJVaHJg
DyueK14ovkcyB8atwqA3Pbty3C/izMZy4C9rYItXRly7H/EsqKarVzyDktNRrItj
bxGgr1/XWDUXe03LS/y6gWtYWzetOD9s9d1QnFRvVCbnJXGO3HA2QWZuszUo3XIP
KDebW/S9AiPVl1ytAGpC8vxMYyxeCnuOzpEUYog40ttkteboq6gY/7WdbF+oRdqC
jXzgBkZTFx33YqKuiznOA9y+bYUWAVnaHHrAb+pQTPUIiTjWAfLThhIDfktRifi3
GMK3N2g4mqkK1aqdoLfDOmbi5mdL7Y3EdywYdWVrG/VqhMYDh21y5f1YPCvWG9OY
P/pcLkl2RgZQD9AiGIhWRqj+hoENb+HTAwY69umcq5lsw99fiUb4V75O4Mu6vR2W
MK6/08kNJEzJqJWVu0z/ae2HRrhQ9up1VMy39T/+aihs7QYYlwDLu2P2dkCPQ3PP
OBXH3O7VH9p5/IjEOYr+9/RcZnCDq78snjyzaNzMeKl1MN5AJPlIPUCzyry2pS7g
q1NAklQ+iDOupGD8yErvELCPwiY01SwZm1resPASGEwz9Si9fzPoRVVnACiWHimK
ZRRwe6ur3l6YU8B/e6v8rvEWlijfCS5yUv1t4XJBD1f+KPw803dpQ3hSaZFWlzJg
pOIM/spLq0HrmPzR+onajseVfMhc/Ivb2GRm6SQ39NPP6gN6HdGR5osYzaqtClAR
IVZQOIWebv/4RvUjQHtjukUiT0Zp3v1TJ5/tKQZgTrsgDSJnDR9V+wUhlYOQlDQn
S45ibUF7NzsdCah22CaK6I8aBy1d6XNJI3HHZJrG9wHVNgrPNcAKo6eemKOBFIFR
dOP+zH9azN4abkHQAss+fLVUG9vRfQ9c5sc+/fX+8yHCqJPyOylQ8hxjkvU0B02D
Fsy9Hbc9RnRcosi3LvjD5TiZm/XSmwZHreiwNgWL5dj20EUWlooWGOOj3VCGhQ98
vv8832Fo+0nfeNj71rBjGDBCDELPEMpJOe2AmZ2AtrmY6dFkUKTBlp1t6AS0tcqe
IIV689owFKrL+XZvEbBIXMw47oRBp0pa+jBK9obFG5n3aa+S51RNTILKZIoNQVjr
gZNCHaKXu1QQiqBrkWw1zwompzYW66xHxj4xjRv6kvilZS7yN1IDwSBMGBIyXmHT
L1vbCF3duf99S1ZFBw8lAFAlv0qjtEOHA7/SVpxdOQrUI0WIEgRUdBUCIdeolye/
p+N4nWfORwFLdK2P4ph5WIkJJyaskbw0eYoEEziFIrL/J7xqDJR5ozneSOBu7V6+
xE7ZO6EAzE5GQatFE2KtREKmIYHsRBMnGGqTd06bsDjEW8CeifYrTmKkvuKWCmnI
gUcC/HA7fTkRJT5cBSCsbl3oBaAPwHjMQBNikPbbD1u3PsULWDsHmD8ha+fZhsbW
repTbiq7bF5mSj3PorBCAEe92uDSnw5r0wRhYdj5+VDY0yp4fDxnUpiiZ98KoD0e
Bons+wsvJk4v4UP31CLoyc8yXh1OD1++PUv8Bgw9hy9s/+YHrdONBjnqiH6C/fkW
1VS5yjb3m1XRx5T/QVmkl4rEdLJl63MX9xNzGmlIqniOR3Td4V5sw3dkgI2rMNu8
qDqjrCxGNxXvLPM9S/pzyhJVgmyPPTS3TbjVTvaNlQmEs6GpKOjXCNrUY4ssLzl4
ncvlJm4VZdEB4QMYpvKS9Ut8sMO4OZ+4nT5LS6oYRlt1rwIQg0GF70dj/x6ZXu4i
fB8BPYpQrzaFeqOSNrRliIRIM72P7Vjxgq7bQTMOJdSlyAnMJfrIuJaR8kfVHCIK
fm7bIYOp+wvbvsUQc6/v+nRvfxZwyusuMsNYldP3mdgsgVjaR+hH0m9/w0ijutg6
rv42uywPm4QuTsCy0zG5Kzf+Ck9v351c7wb5PgjRe7tqG9xqvtr9Vl6/iSwJ599M
34jOWXjOJI/cSiwBHCAeqNuaBnBlNioPdWz/MfGXEBO73l9MtKSkfJeYhn8xQhUu
gkVYGxTMcpF6PT0LOyBLtjbHna3IlRbyp76cL/RPXlnTswkPwT9DTbijTygRXzr1
SuLfCqt5vYteFwMFQxYsKt2k9prz3QLDbZbKcPCQkS3RZtuGb9PgNZtiotDglFRy
S1FXqmBdwcr+gL4NCEctXxNjEUav18qAgsVXiAmvFUq98rU32KGDfhjk+SeMQU6X
iPcXjp2bMmI9+FxuBm2XMOUmn2fHJ2wDuqBWIybEL8jUvj7QuYdVVESSD2/ZXDTl
/cbxKf26JPelzef3r6OkFpTe0MHZiVwdwquU/Bq9f/sysBwh6lYxYcjkO92cs31h
gwEz29INnB4kT/eaBi1jRD014feYCPvo75MFlJ61x4lURCy5yYevhZbVm0wvtiwx
qAqhNQ8FjydR9JdaQDSjX3f3mk4WFvGnaxdUDj5JoGaCbO/u/TjkVQCc4GdTynCl
zWf1+JOye6nDNW6/OtZcRcr7q5h1wMl6dHpufDYVFYcOGkagq5Ysobz1ZzcycwBL
QD4TwkblzS4eZOwH2mqKV5/l/wwTULtknRGbPVgQO9ZHmmcFrj1/iC86mTUbgPut
aqe9XaNqhl73u1ldjGYPITOuZiVBL7ZiG/EEUHN1gmB5z/HTw3k07vrN4z4Nb95v
tW13CzabPOhS2PuGj9qetY6OKUp6uNKhvRiqWDb3GEKMLnl0KAdqqKZm6zaEof+s
PCYtsxEjQzX6s40crgy5qwHf2vE0ZIHRUIt6AJXgz1N4lcFF4D7HRxJg+VoY0fuo
Fq1i3WmQ7Lvi5Da17WiFA6PQyQWrEuMKI4A7F/X6A8c4pKFNvQ+gHS2XOUJA/00K
6x2NCDiH9IxpfF0Yg1Y+SOmAPFjLnbmCrYrfIEIsLNuMGqx+WklI4AJbB9NX+NK4
tOSAoef6KicWxZb89DS6J0GLKheyVVFNPhocsaqx066sh7cOQuYAvKRq2qks4XWV
ZdbbKbmbMBHvn76LQDOscji69wgAhQ4zE6NfiqlURIr2yfPjMXKT9yjj5kQhxJ3x
yuqyoRHn9Petx8nLE32NrSennPgLv6uZdZKz8AAwPS+ZwNDYZquGpA65w1B+RMu1
7J3x0bOh5l8LIPRDt8suCZy88r31m+6GYPD81NCy8gVJkpH+xoAOxOC1hGJYUz0z
hL8xLanOVDssAg+iQUK33ZgOrYU1xrI82Xp3IzLmCQ08xrFWF767uPLXGOoFENFe
tvrvCkvRPNyQjXzKQTP4pXjcz//U9sl+hN1gOU7t2XWE6zuEupZ9DSzL2jVDm+sV
6OIDp0KWehiNuH7XQjq5tgPPSx42ojq+MEYAQrH39ZaJxXEdt/pzrq87Qq6lD5gA
qvAMCJzefe0BB1QxKxxpQI2C+7vVd1hD9gsbndIEv6X2e0L2eBKPAtAIgOMVUGJs
p682Vtv4qXn82DV4HWtMl4dNovcCI58E/cOCvRkbT5kYJsYswdhtSPTi8oj22bvg
z8mNNcgxg/5bIEH7a7iSKrejcMgLEhyPYfMRTm3WycWhdiSvdVNdVAtTpkOjN84W
/392C6VAXfJJR0rqZ4/drzgOLYptXRQgBmAJo+vnDxCRAsbSIQguGtIc1Stc9QJT
nVC/EeWAqIq6RqS0USIvT0nFSOSN2U2yOch/qP0wk7Rsp9NA6pFh8rck7KuBJ4Dx
taidV8TkslkC2PU9L+lrK6Ub2mmmVPHiwyF2oetxrqSjYRymMqznWFWJnQ1PLXDZ
fsCQ40O7Jjv1NqUtuSvNKfB0KeWsWUGp3ieOmXrh6EgBbCyq4nqmYuuMSjlJ7gU5
HgmHJ4LyFAcV1+Vxdkb2ewyXc0AJ83eBR/WC88E+6S5j9cnT1j9QNXBFgTlDQnfJ
5gSEj8IegTQ50kloGusd0Ec6XMzRLo6Ep8nVPxMqz6C4IgckqEAigayqF760vO+g
znv6MBaxgce+XS27qIJAWM5R7tsbdQtRpVi6/DNwOKzRQl5sHOrAuBI6Plrdcdow
T9qRuextcmOxA7+Q+pb3MAGq9uLgBm4lpU13ZHirvhNWyRZTNA/plOYzltmeG9Cg
6uiURnjlEfrxHLmYLc31xJ7jpHn/h19qhTyfpXbLLfdAYUw8KSNH3JFkJhdr7BaM
OUfopuXPXawuLNPeYn3vukDYMApOnmxFQSfhkWJr67194/N1YmD5Br/35ktnl6Vy
Psl4m9ElbNt4aqBUP0+DTNtHD+RNgA2Nidze742Ucaw00e8qq7LGAP3c9CqcmM8D
AWfTvfgZDKOlKxnQFiwq1TjhyEi+lEWjR/n5rQBDwXow7dGZq3p8K0iBdaBCuVi6
AZn+Z0op/eiyuzhD8bsKqUxfWnTl3uiRvxxsg98DAypiVBZKK+K9PttJCIzC3JuZ
+sdHyglkhV2nNcm2EbTY2beACXUPZftR4axGecfFOZF0NJQy88QjbrLrNf01uORm
Yh9OzMeBYJapfguJHdG0T80c6m3+3y+8HmcdAxfKtXY4BtvxlQuIjtt88LEropq7
OUqZUv1taahTxfYlqSr1iHtSSg0S+Kea/qasZZPe4N/gB0DC8Q+8ZnCfB43beCAP
7DncyYYoyJFwvtzhTFSLjFrhHL5evH2fgJMGKrcPpLUaRb2tOZIykT52CliViK9e
RTAARsOWj/Ll4eg+XPo/MCyHDzNSjDIBH4jv0AtuBY+pfYtXd8Xp6ViG0RQaivIq
X1osNKY2mhilhiHs1fwqnYtwZYxKljCDsdg8syq6KtSmYN7DWII70Dn8JpR1jK8k
+UxhkgtgBiFPO4nztaXSrLAVgDYuAanPgZA2RwSNqAS7d75SXg7qMeBLvM9q91wU
MvFT8asrCLfeFxEcuElf/orRYWmJgjox4y5VZSBlQU+DHRsGyXmGccYO/RmXmDqt
efyyyOYTb0Np61R/SihmXkHfjBHN0ikwLl9AW2Sye3T+CMpmVecrlNdLYxvEG8kp
X6GEuwN1GoyDPXqFWbu03EH/LyTZZkx4xLFdD7eDXwaHRvCwmEKiW8neG4qvyUHt
0O30FZs8Hh5G5w3tgTIpyjkS0F7R1E5u44K5NpYoB2+csh0gWXpeuMFTjJyPGSh1
BzSLUF0xB5qFTNqIC0r38slWzJjNUbWuk+XxXS1sXdBmIDUCUR1LZbJFm076kOz7
n0kK5zlrM0eQi0LiVnohaA/v9TjOlUcSsBkkwKvWdAGVQCQ83YYfdMMYZIqm2ijD
7J9U3kSr/vrQM5IKBr/acJOpgOKy9yYLCDUk4cxZ9OznmZz9OSPBp+5GJ/ixaVkS
tl6nAOuqQYe/ll4DCISTCMCRKNWQ2KRjayXNRqNPUBbUhhgGtAZa/CiT8LSznyPS
KZGahOG3zeJTWczx4QbDGDIVHesbD0bjiZfWCk+odO8NfUIjz9//uAzEt5st8vfn
bA+UvEkxAdR3M5PLWTkaZUIqZ0t7hHJ+zRbfdYo+gtRDtreYx95wG+1ojIEyOvEs
Ngzmur3pnm5h8/TKZKj4DB15U+5zW/bwAlgjhpH4uPDhoHX/wEKQkWcAz0Bs+Wao
K0+IztqdvBmUUA89QSYAxJddebw5Otfmcia8b91QjCRvDnIZYc/2EqvEp+qMbb1s
i8inaLq0mFyfgNtaHH79HubYuNDOYiwFNgEeJ+ihD2IcSr8WABH/C+8RHUmW4LMv
9C93T6cs7S48NzR0tiWYBLkGq7bejNcaIFknuxxSNBbUafKsGD9i/cYWtXhalJYL
ehUTYM563dM6tP8ZRj0WFSmWMbiKLYegdiQU3chNzj12w1zeKLr805lTmdG6TYGb
JKp95HzB5+3z0hkB3XbYBADTAskl/QghBJGwkr7x3kAc1TE2hyV5yQr/bqtcpLTr
k0krRUnKcnvNxVpvACe9a6BE7lxagh0I+6QKuVHS97q8t8Zkg4uyrkQqjc/u/ULa
JblTiV2TWCErJSWWJ304ZmaWfZoWxiOzJMjh3N9KCDgBXXeFtKYxS83PfdFP+8Da
Pwb+ShjpyDbcZ1D2NrlTLcvWYjeCu6cj+8WTERa5yc/9O9vIHMEWrsJ+SVAmPGQQ
nDYU0r4Me1PPS2u3hZmSmgKnC5lzIf+EoJPOoYh2avYyLQRgIfWxvLr8bXTCd9dC
wh9UiuXzyhH1Pw73J67RYL+HSdiysFYUwXGPCDGfQ8q+tyH0qm879d7b5CQynbWT
IKxmnOAtfFdSPedkxdU9qMiOhr0B0ijAEEfLDSZ3qkiXysk1aqXeFLLnsO7rif+v
IMIYo/2AuU/Y8QbUZubLwtWrI6B0hiGokmgupMnlovUfiXluaWmaybTF3GcR/O7x
qMXp8YwSACpLY8Rhc0xKqPsZrYxdwYstLb5/YDI/uYHWTg3w7+ter5hFuzlefqeO
QsJgYIKFIotk1y9S/s6nsqbhnw1ISkYYmJqY2QP9TP7FFg232KzjliZGV1IGS3YH
3SGx8LdYXZbxWSg5nEFIvzPcyIw3ni2pWF0OatHRAFiWtPVTG0igMvZqp/8nU8rN
GJi+6wtZ9SiKbnHoRLK/+NS9Zvbm9Q2MxtnduR7CaPSzSUzGz8BYV8VjJmqV6/uO
MhvRQ21wddDoaNwmQFuVAm0o8PSL103/0piOX27KOuBZJbQbqOGvze7ltmLl0NDf
R+Cy+/YHduWlh6BWqljZahuMSOI2o0SUhXm23NqXDvERWe7lC5/+X4zZeeD+cLg8
x8+ntGsQ05YZMbnDmJDSGwDD02B9aDrgyGmMz4CWwcJC5IhlD4W6Y99V9VCjvKl1
qkrM7XHceMhSu6Z675g1DlnE9Zz9tkKjr7F8oEW1qPp4XOcvUTACLaazcz2Nu+7i
7H0kqNwYq9TfypnTMK0b8DNO4kgVJ936xmtjk2jOpl3iPGJdpG02udw3mVTZ1E1x
Vf3rMTHla0w6iC2OOngv3G5oF94xgU2SRX6s3GRKJWCmy6nAR1YhVhYA//DqICVQ
FCeudd2m9TzHaFJ+qpICykot6sDINjtk1ZOQZUd2XPMMXest0hNfqTKJWpxxsXRc
y0t+3rgtttPR64yy4i59lD+nWMvTdzQZZ3c8pYkeuGr9Xwtt7IKT1Y4LsOzzqE2v
DWtNqZZc2hMn3U52t6tqj3ZYwZdaYWu3wR1BzYKIQPzPE5MDaAbfFF5s1HV1ujp3
hovylqMkPATp5yD3ecAGzHZ8HuvO5wr3QD0RRbAdh2P7BIGK+sBZlasftP4rakQD
cihC1V/LiO7ILFw98bnupS+fU5nbNvdol3HwlyTpWVBAUpf05RnSQSSGwe8AjOOC
RLKCq7bfbcA9tfnR7b5ifuN4UUS60NLKcsjDTDlBn8HP/X0UnT1lYkA0qapVOnZB
0Rd/sGav6cAOui+spy+iCBTN8U/yWb/lOJ1KI0N3dcaOhc65phfPsCblcPmAe2oH
QL1heCiOR+rEl/rJcwxAFObT2cyXbd2dh9YLXfSJVM9o66iVlcqDelyn6FIlrVQ0
mSpLMRFa9lbRbj18sNIuLAP6SIV1LyfvPnsMCIkri0Sz9f8xVBidQ665P/zI/m0a
0PrWJQmz5lncPwfIQDxDUm0EwXDqQ9h0dQYqUsmf5hTabKq0AAqR+eLLU13uXieD
PGWAVbdTGc0B4vsg0Ns0ujND+HwFNVwTAtW8kqmDjiljYZoSU/OxjIsmgc4eqtnb
5ewdpSA4JSw5jA0/T1zJXCuignznW7s4sYRiJgr37qo989JjRPbK5JPKZsikykuv
8J7inqGE/Qo/QPfWCsWVihrhjB2citwY5ru8OmmF+4QNs+2PZpIkX7H3ASyvfYuv
fqcn34IK3XuOJJtV9Wy03e5NjjSPW2fCLZ8XwHTrQITmrulefDZsUSh1KSv+gO8h
5ZY79lOF+Wi3VZAtbx6JDKsFjCX6ZWuIAHNeyUCh4xiqH1262vbtRE/7QrxQmVwT
Tr1MM1Au6mThfzX4u7InwnQHevSVmlYXutyaLRnOlyfshDRrDWdPT4uTzRLD9Njw
H3aVOaDGB+wvuRMGb9ye84Fwh4srLxN4NjEOj+dKK6C1RdH6RnUa9yOBWsy1btw9
Id3VR2hF/zeyBigzRBBMCsNhc0fjb14JPz/CfZ/zPz7AX5l6V1v5egzMfYWZnIz1
aVroQhGFDEzCVuzBbj9vmgn0XG1WBtP/xjvLan74fNSbr4fUFEo7FHiylPUVVEOV
jddNDnyLs00FxW/MxVwfBrlVB39ksCa/Q6nOqpIpGw3ffhtkCN6lUXCL+bSKVGwL
Y0heSSNaubSMKprqz8gqd/RqreP/nv9OJom37i3cZaIUBMCEjiX5YEe6FEKa5ifY
d3Z4kv0iVuhe9LUhL2uGtg1j77H6YfIf7h8xfIr2uifVJcHk+BYo8W1e5bsf0z+V
r3Jjf99OdqhiiZxJRWnhHDvTuHq7JHsJEQYsTbEbQO1COKo9VDLYYb/H+VOBOMH0
gtaefs2ZwmOm96SZlqLJGJ3SZjPp7eMVfEapXbDF4SsJup3fm+d2Ys507hiI1aXY
nuTCbobH8CVVkd867AOeJpvVWssLJKb6srZf855PA4L4/012lLiocevXkF9opJM8
YwJ94rMrIS++mon+fKaJ2JbXjhIAOhEHvhv43FZgsBJnIkEoq3D1ZqsHERx0wybx
ZbLeaQbDbjtavnSgH1UqRTub0VdrjDKTyOWdjcbxeyFQctkK4wwfRWVNZa0BUi/Q
PcEL5XW2T+LFJ6AIy6EZ6i1BB6kyPWBLao/l72cXUI2nf15byfBJL/GcIis8wsJ9
dmMbnmqi1djPB8bKGohzkVR9KSmaIukOSGesUj+9edYepBGsIYvQAm3EAqpMTn5M
IaoTZa2UsJ24/IlFtbn/QmcQSNi+VQTtnNTO5qNXynfVUGIeN0Y/P9MrFaH1dNrK
u5YQ7DUyJpbH68kMyblsxbyKXsuOj2uFV8CGvkhy0DCXF2Sm5olfMCBTP15vI32c
rsAVZ24pOM49i6sqlb4cXWzzCNIlOBV5O4k3eCg4fun7xDXjBKMVccM5zt/drIYx
dRb7/TkueiPRGv4sBpKHvdm4f4pVu7JKFYsOdXPf2vSqipOASDmtHSH2Ar9JIU9O
o48/gNQUU/VezUe3KxDdVCTtiFNAyRC+SBIGnz6JBR7i0pQXPWqeKN+gabuO2/RG
oe+Eq4FTn289hbeoodPtiWOU9RMjlUk6QJiaMtIyO3IxfEp4iCTKpa0rjwvU8+TM
4t1rKHoQQJAYCAvc7JR3lsCLpebFmu71V3RnnqxGjmdQZgQF8hVNm0hghgafOO8D
sKb3EtdeHFtD7BJT20NAzTZK71lKOa37LAN6GgA6dk1l6qL0ktc3O26BokGrm/tr
SqOv5KdStIFRMgX+NirOIqdVXUpuBkbddsZM7W6hdQl5DFzLQ1tkV1UQe1c0F78a
VU19/++VXqnDGdaVgxsHgUluiR679xEVO+FNjeGvHi6y9e7iAnueicZp8+Q14nXj
tg3Uhn1toVstkt2QqFUqAOtKHLfSpIfthcU6Q/TrTYRlsjPvkI72t8/1Q85wAwPj
ZiHTD0gv99kbFi3DHuYPAbk77i5vB7jd3Jv3r9jHoxUHiBy1jMhWBTcHT/6i5SqO
sZkWjkNFjOj3qaXtKZrNkiPniqlc41a52MhQIGCW9e5dupzQPaTOgCsaJgCEN72N
4LO9gBLdkMIuMzAv7ppdTvPNTW3BiSIxWGMxBeBdx7hDXDQZrmGExIL3+v7BQq30
OROszSKWumfuPIK0cA7Vd65sBBTNx90ObBfXUkMDmk3D0KThzog9V/Wiep1JOtXO
09U2nXqTTyMvk0b4XnR2KRE06IZSAZ77h8g0asbKgQSvQ8Gxgz7M6ilwdLgizIbQ
4l0y+jzUnnrCUGeYNVI0Dg==
`protect END_PROTECTED