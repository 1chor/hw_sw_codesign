-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tdc2E/CCVsh8r14RFe8CC96Zb2ppFv261BohhpDB11dJuWQelP7lfmcWTo3eoKXE
q2YL7l15Fr7OmxLxKMSI3ogoFYkRPWh7fIhkxo7qZp3/OMzMT9iQ03gq4PRtDUNf
Qeq8RA5Xgbxk4rz9P0qa46jygYqbnQphEQsvhZ3Yv5E=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8624)
`protect data_block
ySmSyigJDJuWpts9dClnE+WRy7f5qV/hrcv+UhT1mUxc7vltK/O9bDi4P9lCvaVk
Ovgh3QR3KSpMaLqEy3g7N/zsDbT5NFE7RlSwEqmo6/vezfN9EyYu1pZz9AWdKpjJ
lok/K62NjPkFOd/2CsT18fHpQHxnA6JL3DHs6Wh47mWnyggprGVMxXpfydBmzEEq
gz8W+miLPmAB6o+8b2b6J4DzxANdUtZpmwpy1wADRElM4gCt49fFHKhIIeht4WuA
R4FHmU2Pab1ukEuGswjmteKEmVBNVAh/Qb8n0e0d5twr9bzoO3FQ+7MIUSXVvR6K
vdAp0nbj7YLRB1L4Ll81hQDkofNdXUjQQn6kRtJ6u5ekaGPOVGyAS/7q1UUO6vI2
QyVFEpLKEF49BQ/ieVq4JfBsI1SMnSkatkYhQLoiCdEEwowoH9IvzJbDWoqxAXNK
nuB0VqrlZnEuKA1BBEuBY6NnHOt3lMLJm93BQYPto5n2LEXtkvUoC3HPW/Ww5j5S
ElFTw3/TV13YJuXdjOTYdE5slTH2KEyDCxNW3/6ihbymZnBbwwZ4qYMDocqbkK19
M2sWAMbsnvKEUl1REjqZccEpqI4YPwlX4JuSVu0Ahil5y8L3sVrPqgmUUNq7bnnb
GXAIiuaxD5sCgbo9BQQQkHqAK4btPjijLQaPnulLQN5GGlnhBzwO0G/q3RR0e1U4
cIeCXAGaU5IayGAFUuHf0/YCA8fSyrkc/7VLJ3fSpwb0Ggo3UsTuIxvgZMUt8ZVm
UnHrljMVnrjVwc5ybVqrIup9r71RWOA7nZ4SqFBpIpU/t3vLGaHaoOMVdNeWxcvL
2ajL3lyHOngveooBqyn/EK9QHutC8CtOQOjHYMIrKy1haFKlwvm94xkmBovN8EF3
5AMK3EYs4H+GViLkxwWHOF/TgWgqKgnJmaCnxpau7MCvGo7Q/KgcpDQPAouMtpPr
zGD7p/cfT4hSp+0sdnULH/3Isr0vTq7R30xIB9X08lc9Y404NS1tIrcjGIjsoqHR
eu3+mF9fFVDXAILQknitJxFZ0i+ITB5DGGamLVZZcAbEE4JK+iSABYRpRtU5JLMN
NdpBJOkYcr/FJitGXHPFFBqAnuf/YJ/9ifYQFujtKtcAeoh3xhLdlrTLqbWDYzJD
p/SFZkfTPX7JvaKlSEvmnieNzZaNHWZWbCBjGQYOD27OpT0D6LyAD1qgpyybHLUI
BlJh8izFwBEWT2XhFWMAUlART2LRswOOVlBH95mE1xODCtZFqLLf3W/zjuN5blQi
DNqSD1Z0XyD2g1f+RFpaJZyiN5VyxNFqPp3Ti2fkaDkswDjkvnTFoAaReexS9WqH
F/d1KAdHsR7hhww8df1AibXdAAhryQvn4K97W7MmGsHCd+0DsjuhpRY3sdMgHwCR
JfINuGltSdF73ZN++b8f9X1UI9Y7pg/Hc5cGEsqrXfnIWsEMBXJ1x6GIkkqfYpfd
n/QtUH8hWY+79w4S9Qt+FVC4g9ZasI/8ndoWLgzoS5FbyDO/tqYi6KzcX4GFXTlX
tUM2L1JQyXjIjPmvUFO/jSaVBWpt2HGYbI6aegEy/Jze6pTp6kwYdWZG7/bQ53L9
HZL1tlvNZtoO4sZS8x4g3KTfI7oZeO2Bin9/AbHN3oVerD0fwhtzJhFD3WHQFEEu
zriI+5jcbTgVuEjAeWb4hUqbUK/PAsME2qClxJ9m5SNXA+fpqE8OlZWKi5jM9LQe
EXXJy+6RWz2ObkR2M9TPf7wT/4HBEBjwKnfOR/FqJV9YKrg8PyHgfuQMkdB22UQ3
2JBrR2kA2HWa6XvaX98xSNwstjnm09gy+wKfAdgE9v1DLhcpzksPUgJV/eRbPbDe
n1iF1jKYZDVvxBxGvR9UAG575z8A3a43grMLqSiJMgfsru/rxWtsVIb3YU//Vhy4
6+ZxbUYHE1hYGgSuJjikIpRjCc6qm/BpFfpOXVTHID5FX+2WVx9m8We6HZKwfqas
0vdZizHONGK6oTAVsWqP2Ux/2YlgCyI/EqY9+vNC20fGrw6fyk9Npn7TzUPXEBI2
ElOwrQB/magx2pJ6Mn9W4DdvIKwukha+6vGkwOdxjTpKsp8KgnmpgpmzXbpyQ4ml
blva6098UL6TNJRKvjGGaT/KdANZQF3uCmyex4xXh3QJx8fg63gOdf1npnDHPyJ6
TMFam/tcg7/KUrlSVhOQNhAJCp7gRKMrcKUL/6CFblY6yGlvVkkR1nqJp8viJ5tC
P6l4JBDcDSfBCfAoWtFg70DJ4mFouTVjORUfWbKw37WAdDbKSWYQZW+abaGDzdOg
2GjA8oHor+V0Gp+PNYENlAaMoDtKZixGj3/PZUhkuhrxRT5BZ7Pf7XhWv9GN18jC
WTV5SPdL1gLLUxkknrmmDWCcbFjfvhOUD7NY45nIp6HJA1qC85Xc4YrNiTgH1RFA
9bFXV1irgIWU7KW8mSaDyKwmQgxQAmlegAMEd61N6U2x1J2EwxqGQDEaB1gIMBba
noEhSgD69vyJxqxLXkHeU8N25K9RTov2KJmev2gv8AiY3U9/DhFP0C0o/3FJB0Lv
yezo2v9EclB5CQORI52+szoPVBZhpFnHO/RBQCOBs9lzTkjErPNpSkBBWGM1qOZR
Nmg82GsrIeRfB59HCdvV/so+NxvvLEL+Y951WteHArBWEh05Gm5HkR0F/dUC8tWW
hbAulpKb1hSNpci4uvZkoXluYxc7k32db6y3NAjkpqnD5BNfK0m2+ecp31gW1TOi
a7KsVudhbO1bWKsKkfvn3ufiMQy1ZRHtMXvePO43mGc8Vmw4Xkvy49Ee1zjyvtHR
Owxxla7K38HdpiZipEaxU5lFFVRijNXr/VkTwp8XrNI/BV123ovnXjz3GdpD/tvP
nrO65eRahAruhUADreHcoAAuCH/Nu97bjZp5HJnw8Cy1z7z+w0CQQtroURb4yoCk
GD1gYXIKLv91KZh/tPh4CwbT2GUm75QLsDdzim3aPHn2JdRhf9+/XF0n/5XtGO4C
v0F/nWj+G4i766KIm0tMTT43EHltcLj7KkBKWvHJb6sLVnQhOKaAreCqvjK6/auI
09xOhndewbZNuAs4tnaroHD+8dUhDdEHwFT7ZdRRBJ7X88Nmy4vrifhTwCpijZH1
1PsJ1hjsnSNQVHeda3EuR6N1luucvw9py4s6KXCThcR38iYKJehcQcyaekL5ZkPh
HwvjGEFRpC0tLYSpE8rx2r667c+BUsSjF1NIF24/s6SKuKuX0Hz/Y5WWtsv2pGXv
3PXeJiKA1AxtGJ1uRM7uwkFxyM9iYDBvGh1ACG+oqEOBIty+/Iw3XRBXnE25E6en
AL3Cb3lK6jEM0U8gHR1I1brTl60WBzBQ4tvfKoHYdtg4cijkO4BPJ6iXsTT7E7oC
bfnXLmUbvvyT8yjy5TQnMnqN/zatDPeJxPSST4MuvvoM3t3CFPagz3gm5GsZ7ZVJ
WRQaGQSmLzhAFRd4S17STQfoe42sGKgPWjP9ru4dcaYG1xGFje+sO/gOtu7vzPKa
o7IjTFxVjZ/aChjRc88bOsxV0nmU696LoYBNou+RL3O63ixJOQdzwocrsGMA8lHr
yNUK+sDn2QlPqqdGmDbQNTG5aY8FO7JduadLtBPl+rv5NSx5wR3Weo0JTlBJRtLj
IoHe0MCdhbO1b03Kdxix0e65L3Srq8STWkWxZhpGcM1CzN+mxQKVsJ89NPkkh2Rq
8Rjk31TeOTqhzVFlgR/qHQWssrswmq2qbBlL0q+UiqOwlQXZjoPdEAwYkJoHI9Bz
pBlu2hK51tklyAYQlzSgXmcKoJQ9YYOku4XE0/W3bHG46yYCCwEBDonvUe7YsH7z
NwJzGskntZqAAN5NatN/zT+IbOGRjLUpxp+tfbJGUOMU2pdtuFmgixLn1usW4cGQ
SxmPpFmPdF7wyG2sXh4tOp4wJ28YIuFFld/cJmTb2mDVGfJm/KiZlKpQCc0uTdC+
i6vPpZoBK7x7DTaQYT2+ezrY9AxtjZtcwCsQcBNrrLKnp002bL2ed4dlKyxzcTmy
BwZ1G5Ap9h3zRsRiOQmZciR7lCv8XO90D0Q0bJBXSYy7p/z+yyi3MjoU+SYOCsp5
2Npr4S9szqUdifGw8QSxU156n1ZCWn/urAVHuz3JjUiMwyV8BiZPHq0Kb8h8io1T
7tCcYCd/lIQJD3rdY5sd/ngsw8u/0+6JynzcON6kM6+KI9Ph8CSbEN1Xpk14128m
lmkozGvI4YVvaD9QRJqP2dJ+HZcpQRn+eHFIIdQ0JuciKcI14shIUu/Rh5qIeI+W
IWuJpi2vKGshl0oeuADVbDUQXbW7HZ7u8ac7CIvsKDwjsRqh0qkUaZfAxMj9zQ5E
JTtDllLzb0oe9K53alTvQNkxIUtKQ4sc9+hi6qM9EYoUxjpWlK0mB3eQGoeBKLBB
OyQ2Jy2ufsjNtWLvILYzh5Ybf3Udfeg5zkbzMliLyzXIwfaeoajuvYqsgBzjb9xY
7qNfpMBzroohyo86ndSIZAXQJqh2wD7rliQEe5MQuxNH5P7JqMVrjZdpvv3JG8mH
dXyRw9IdjZL94i9ZZ94kg2MWLsVo6LcwzxrOefOS+IgbcpZyVExOgnD2FkVKZ1Ht
PQk5x9sjwFRqykBAE/YAE9wnEVwWsba0RHw6dbsBd+H+u3N3gh2TURBIs/WzrVc8
8rdCuL4e8sfS2Sc6dn6cH4VvXdd1ezEcYjk9v3kQBPkRRG1ReXXEaAtmwBcY3QcV
MWglx6sTs+4RTyO62nIq+gzMLzZlv0Kje+CfXa2s1ky0YfiCx9CyhCkNGriUGe1q
SfDjAuL98Z0SScjLbL5aNiZZpiWudEnhFvllrjTZBxaUJFWp25F35t3uK2VFbK8e
SzpMNqNzIrR6Cj4esDvkl2EzJlPvwk/FV9SblVHlh7M+IsID7Q9Z0drjFxrxKIip
sh5NZBAEMlw0yAtECZAN5vvcC0fFh7BbmEYizHE08dueSDSESVDmvSTfSwlCUoXS
ft53lT/JYyqJS2hCdy77fl1UVUxtbBExmslmN4vH80lXjtYVzyVaZqNikPAA2WRr
AO7f+N3r14yyANc4TwWnei/b5dEEZbiO8udWd5lBlolX+7wQhzb3cNqIzn1XdgLm
tF7druqv+6pcZuqbTaDTW+pxNY7uKI/9jJDkjm1PiuKAuwvQdINm0Vw46FAPayoe
vI7cpRi+I9tQdH8lsPIejJmKgegVhd++o33B5fY9JBtS95LXN7hRafT+wVyLiyRH
eDmGX3XsERWlRb/OamEHEwM39LFL7ttpYduOgDmlHiSUKD8Gvatn6XsqlGzFvkrE
XwG/sccss+QyzQaoxOJX+wwRcYezPQclOQgwR7cyaV7QnRPRtL8IwGwW1N5bFNRq
IFeoU8F85m4nRsJHMHAM0QHagBwqvyvUN7NemNyNr5Lx+uN+aToigYSB3BM/oLYp
y93ZdK0uWTa3D1E1cY/iRFZKwwPKA2px5F+WHjQR58iSZy/mNQqkDUWGIwPgxzbI
TmkFJ9gi2wf0+3eXvT0NtghXrOChVcduWi32gl5I4RF1pEkLfp4v+AzYbPrgbUDh
7WAsSIIMhbP6b1TS4Z+wBNaFJrh2FgjaNpFEltrssJ90RTTeOvrbw5mLnarpFnGD
n0oqyBy6iUMC3L/3enwaxRzL9Na/yeH2ypN+1yfsS1+pcm6cYvxdD/oESHW8/qod
ANWTl7d6asTspKvuAFnRyOxJNQR0gCczW2L+W/89r9MoG4Qi9mCZSDzL0T/4BlVS
wkInuTs0gmsDwkw0YfotIRnvy6257M8kMyNmM6OeWlQ1gpw5MPLVXb4QK+VLyghb
wFCr6V8guu/7i7SURnlhffx4t/iQjGl6RWg7OgOMDFz+3byd7a1Ya8Nbe9zPi7dM
tJqndlOw1+hYkg5V8vQIAA4A1iKxLTETmWXllvO6Hox2mPM37Ujn0uXKqqhRnEqQ
Vd/iqoOjMQ37Y+AE4tX3sVeV8hDndH/2q1fPz676sGa1T6vFynmvEcLEihZAxY5E
pD7wDme7z3vaY9+DQmVPrJF+qFw+qg0Y+zbiJ+m3X0Q0P8miurgvtIdwBnaIB9rd
VrOwWskXWC8xgJsqT6zf3RggDZTrVa0BFMOoUGypJQ2oA0G4rrlUC7wcZrkNCK+r
Q9hCXFaZ3lRvvUEUFhQcFNYGP8H2o2DP1K4o8hq4zySQyHfI6s1ctERnAt/YMM7F
Kqsm69oZEgqdD65w/5USFd/jgP+sunjtwNNTBmUFskwYQOiXtUVVvFU/w0DPCyXe
3JbY1qouYAon44fn4E/Ue2ahI/rsVWfmBZ/xU4jv9tXMDslb1+PhrLU0QEKF6G+b
9mpEUoirAKicXcfs+5hHVXNClk8nAG8S+HwsnahTwYBVEwIiUMCwip0SviKlKtSp
HrMCJvnHuDkznu7zMrFWHxjPh2uFOUwgVZ6nC4IMw1ZP7dLxOSUleRqF9D1Gp+ys
aEVCh6T/LAN3+7bIXoKwuiFmBdpgfGJ8EXLF4rxxRMExtDRbBPvSk8BNrE1KeEFF
6hpur7k0BY0v05H1qIINXvDdGztEjbd22SayQls0qKvw3tAW8q61gPwoxPKbLM5S
AlHIEqVONFDqtTRb3GQ7wLD5oyzkzLYCr0CjhIdkNO8awZRzfFtkhA4H26N6ixr3
R6mDgyNeAr8I04iiAkNASeO67G2eTSDN2f4ofOLQ2WWdmTJetNcfxlZM2lmxREsM
aqPErRBsH4gmkUli+1a/WH/Vg4sfTcGx5N+xrxoRmO4f2x3vatP3vK2Ezl8Imyyk
EERBvFVDFnj58Y1HkInBwjZSfDA4d5uYmzc/JlNTtVUhlHs0i44CoJDp5JdJ86Qx
lWunwf7uZNO+7ewNbllZRscoR3CBr4WR/k79rH1fKzUfYGCqwv104Nf7b9XQ8/1j
8+eSn8vK5PKjJbtHxPSWCgvAU5VP6uBmSumWYuwYcvBfXHtjbX/zyBfz6l/zUwen
8orAsWpc+5ZTtwdkeP0ubyp2iQDK5uq0FSTVjBGP8XmVx7pKxzhvu+T8+Dsvf3uy
YXuKRkYeovgJwAoEIhD2yY+cwdUTev65mpzUhSJ0RLmP1yCyjLV5GSSeCIu7ByO0
Gz5K0TQIed2RkWwPkUkV7QGY3PW0KhJgmWu/CopDrVmFHqoRvuRk8d+hmJI0A3NK
yXg8SEoV02MWJyqKYQlhibKN6owsETGAPz6TUhZh5BcsfDOmJ5FplXYdfPTU00y2
B/mhibX6qB7/772uw00AecqNp5RA1Nu/gSBGBI80btWGx0QX0/2SSyDnneHGdRbX
bFkwOMVdRU3yqlmyzI59B6OwGSrNeOqyhzQBXlCWK1FvNomq9R+n0UWNaosMyjAX
rymqqrWL/lnVOurfD7VJ56RrtBBF0qwlqhf0ovJu6jTs+0z2yVK6BgG2cEPMsb6x
NKqIrYcToqh4biiQDBBZN3MP/pTshYx6wYzA6RVaOZ51zBpTgsppqJE3lACChQSu
XLGJToBsJDyPxVJE+l5X9+fz9reOh8i0pTqQCmIaTQsXBYFNcKA5DFpd9v3Jn4Fw
2Yg494UfsY05B2lhtd3tVNIy0M0/ciuMf88MAc7T2qEtn7Iyuy+tHZCwfUC5qTjN
5bF5iYaYic8EyPnKuT1hpS4PLGsnD6fx46jwikHww/K26N3q0rCD120nOl5JkWz/
7KSEjXyWxQtWv8ZLzY0zsJppUgmb4t9ihGtgLPB7lK0kkxVSE7W90/xN4yAP+tht
jazzNiYbpt8TaWAzaVn7Egi5EhfaVDl9gZZIHI04CqALDEdpTfiGZtKzyhOMWYoU
6BgUOCilBLG9wniMdN82FAfrw1MSoDAP4+NhK0RTI01maswfSbMb1IVp6OCFB3Hi
e5T7I5Qw18Rfga7KBLq6w2RhVk8afZ4jbqD/t0KHZyLrjg4oAz5PaXSldbx2iJSP
pYYDJ+JOV6mPh/XTe6FUfL1xgcCiWXzm865XVbpAbkrZOuQaS6stL3weSHx6sOg6
w6Bj/+hf/MUn0t81ny88GuZNTDrG8gkYLY64xWz5k7+2MCW7bV7eqCmCKcEMMT3I
0BD9Np5rt3RDfqrBQVGgJmc5RHs0YWrWh1Dl7pbL+hrcf861vHaZzyiP2ZeGr+Ur
V5a7mSMnWo6Qlrniv0f82yf5tudiTDDGQU25puE1pD1y7A/+eHvGy5oU6fLQmr3v
+jhH8u7I9pxhkQGymTrq9/Y2KuFcVGRYQUjVnfkZF1bPNMbXq9MCLmLqxLNjnbGH
r7QK3v6S9CcxhUWQkBEuafzEbIUJPgKFVa1U9Rm/J5RvgvoVb0lUr5MCEsHc5zOj
wqZLMm627E1Hob+HeKaYRN9fAqtG+lb7lIydfDPA9BIitTbEwkqwTkwaggljSp2d
unxidoUDExtgsNQC6ebXx8h+rnucHTRwAG0NNgmyIFHp35zv7xgT1jyYSK8WomUH
xXlI3Udp78ik0lIyclejwtxoUbRETgHcPM0Fo5H/WYErY49C/E2FEn+EUAvBLgZT
UIYGydCOfCR5QKcLafN0qmlQJP103+2DdiqWll1/3B5ofRrgZcdSmzhKgesQnvsL
uS2jd1C+PciSQ+bbQGiy7QujyheLYZU4GECVw3mCB7LST0L0Fr9H0hW3uIRsOoFz
/aZgzGsNSywKrKgd6WP31MxClFNpMCIOx5ri5YJRplAypjb1vZ+UvGyBB5ar1MD7
kyimVQgEIRQvXLFnL85sL+N5gm3J2GN8GaECI/ZaT+vNC9zyoDdY2AVgos+Y5+Bb
cneg/AW+qpGrvxfnH+G8LTC2aqLXtkSadmd3nJjc9W9TNHOnqpFqlNhL78i/+0cl
oe8buhX/P8KsY2qRWGNAWKK3pLlm4xPowNIySYsebaoF3nCMVnrjDqJPTohq9uVM
0Zd82TdID9QtPtvjkMmZRA8SBlxUuo1YZQa4w2bcFS9vaI1Np174g5jEVFUjOQxX
DxPvQwdpZW2mraatMMT9aYDERuq2KHD+rMDYanS0rpw7Stt1sOA0PNgQqhf4JKuU
Hi6JPe2k1BDPG5n0o2c6rN/J01nJDkqkd3UNpovh4o4n0h05xmAbFDvmCXnzypwb
Ei9ehI7z2LTYHMaOLHXH8PMvfWmEG6YQuH0SDbN8USatMKU47MKRBu/C4pJjuScu
61zJzP3izbAC51/acfDk2PTNHiX5+fKJkxEwXB1gfaVq95VmIHcyEU0d1PH+bZrK
XR0CNCpjPmHbSudhLf1kpCHgepYsDTcgaZEfqW04kdCFhsXr+LPVqBzzZ2yOJYv3
t7i2Kl2R0U8HgJi/6DbAGkMtrw6vO1c57T28QxtAwFEHMkXx2wmKk+P61JjXXRk0
Jsf1woBVBlMFTVYMvqaEYzZpB0ixpLKQpH8GMrbCT47cwhOe3ISdvWYwHgpna+VM
dNkSmcAV6duWgWZ3cTOWcY7A4NzCu2Ivj4/PCGKeFgmWnF4O9wPBn92MyHxM7SaA
s+5xUaqQBkKB8xDvs6w06QiqREOaiFhTV9jPssxTaGrhV/O81KMU1vthac7TmOeA
CwH4fJ6f6zV26vwj1Y4Ne3qsEcjCkbhe8wNV2v2BvySK6hMPF2m0WdPJpHVrnwuY
a4SEbqjgsmdHgaNtouaS2/07LzcysOPCDCdO7XMgqsWvCOQp6Ko50HovPZe24dJE
AiJ4I5onwN8stDdk8Ue0dnNW+38TCdK9y/1WiRymDeL9PGRJuyOkhWrusYtvtuWH
q1m+QFXGso7pU5muZSmuDVp/wyjPb6dxTL7Db4cCu1sy9S+Wg7j7LLn5gpWP+K/D
9xyLCZy4eIdSFxSyEezqI4tW8yZw05BjB+/VEuLnDgYs4ocdcdq5l9UqEwTY5tzl
yu1xKvqINkMn99BsuO4a0QVWiuoDkA219uPu18t3rOznsnTOgIkmj2qRNR582e3S
bL/dvcBdcT+6xvuyGpcaxFfhyW5w7P4I/OYTxGxKJd8zhEO9a95gPz1NkQ43QCVi
fiw/xboxCocQCehuxmkvEbj7OhQe1MOThh7Weyu3KhEsJVLSJVDVdXzZiMaDSJut
DMb+r9euhwZpzfmmQZRcmZTWHNJf/xZ9guMMQXLpkRmo4J44ljCdb3YXboB/qsVt
Gp+hO6Lq6LgVp8RhrLVL2bjcwfmoABFlgZY3EMk/ov8E/arpF8icch7IpoIus9Au
lCL6wfBgQ3rXulLwABgwum61mMCr0wLgUCDnyml+KwmHKCYqv5AcGFzeGPy49IP1
q6lGyKb7sU83mtTndXrB/RL2yKP/jkxCVaEG4GkzcyaYNVdH41MHQv+9fProFDdc
0ItkNzl/QekYNTW60rWcxvywnHwWWftyJy9lj8ggiUuMDhVYn25n8+zC+WvIFOIq
rMRmkv8PegLQ4fNRFsU4DMKQyq4EGBPuAYeKVY7VGGq1r6/hmd5HMoPO9Zemf9Df
sOJ85oyNFefg3c7RnFNnwgc+d7N34+oLBtVKrytnBe+SBz+do9VTjijl4aiYXWIW
Mp7hd/sUdu7dYGmXcJIF8v/yrCkm3+d8eypuLURqLRchDS4h0/mmbLsTEAY/2/+y
QzA9cIGTlBejqxnCnjqx69W9rxOpu7Fkp8UEfq883oSOhGqEbXT4KbLYTTW9iIbK
YbAVjvNR6o54x1sl5AT5K6+Zo6jRrF6lPNIrRmOLtCRq90G22VfpNnvHpvCIWFx5
2EPseaZ/jYyGJs/nnGc8CWTHS97qVMksz7ezWz47RNJFLMFoPJmgMLkq1cmBwvYC
T59MvWj8sFeIxU4uEPg36ZidvC1YhRlc9+PHtDzLj9IlZW5UDAmshDXz/jwrLBUM
gpN+19US07HfD5f0iXNT9GEERZ7awJltVtrgoXUd4qtAocT4A+uShZAd6LqDrQLm
9p9xZYNoXfx0d35glsq371jyyVHhfbj+fOgOuU7dG0ZfUmHbAlwuh1xgpFauQOif
bnADiOa5kxRUjfVpQgykqXLJlr/xuBgT7VKqtu4pEGzT4YGr4Z+TU9k7wODqKyov
s00r0WLtcsl3I7n/wwW/vMiKNpARuFkbcd5bXMPihAj61YuTDQTROdbTyls2IZs+
GqAnyLqNn+kX8ajojz0T6cpF3emeRBhbEQMVi8cHnY1MBlbn90MeqjfzNWxLQ0Ik
CFBHVVkEN7tCZJT6yxd3toFfECw7/vZ0WgWGLSu+3g4WYR3v5WgLsWgVXOjuAc8H
E8loJoGAo4CzaQQF4nspkSG3/8HEQ2RU4ryWR7+1nyK3VRplpBR6xxVvkU+Xb1EF
g8b1OAHgfvhTw6SUQbBNd49blqqoEA6noA6ZFeMGYUKBOwHkYwSf8AUy8LsCo8Ho
mr/FRYW8CwKui2G6r+8v12sMcLmuzF36w87LbAPwv64K+CS8juCa9inLKBe8snxh
w1H9LP6CGsynrg6wVsvtzzO3nq83SLxn+6N+sUDIlL9coKwF+UEeKPzMcV8GrNY4
+nBI/N2HQdsKO5vn3pG2ipi/o3781aLFQLKAKZKxtIA=
`protect end_protected
