-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sS4wnvlWjEn5mc7PS8qQ+EwONNZAQalwhOdfnYdyggfN+2aaXzN6VRwCVMuguJ4/ANQFdJS9YBD6
zjjTvUbVoIlyFHlkoKsndcuzrzAS/4Xv1uTruiUsewyfwvLdXVySs3n208nb0KqLvrgOuhdifAWu
Eeqzy/opVG8KG9DJyhaGvv4Ho4vwvn7II2u3ijVGqNj4HBqUO/MteMDij6/tcRD4Vn2Roa9evtjp
VlXf1w3C/nSVu4muWJmQaYuC/JC7l4a6cmCvQ5uw645Y2+SnrRwGQtFFVnEMNNB7RaoL1YZ4H+Rj
m1cEdVM/2167a5SLuIG2OYN8ce5fP4lBntbAMQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7536)
`protect data_block
Yd1Fgo5JBiaM1JehVzdx1TNZNXSalFde4Gwm7/8a7VP1GMIPDmyUlo/I9eBxAMofHYDGLNwCNqoH
cJg7wfhDYEkTap28bnj/lKX8MXiAtaOeUT5LnZqd3UcKHy9NEYorVs6P7ArjqEqDA4l9cF4rR5kP
4iIPBcnGF/KhOD80N4qxR11QJIgMVs5FAEjS9m+LvoBVpVwIKZaiePcd1xc82tTBbu0ScL29LpQz
/GimMGH3ATwvHKc9y+T/vk1NtyQUpPx5mKcBpOc+V0+Rh/GqTkuArLrJna+ZSFlcKTtPT8ZB26vV
k8NmE7YnNzUgUgsYwVtMM8xmwH9Pr2auN5mNsfG38UWjx/RTrvlCQAD7wtlN9aZr/JRDz/gtj60f
EwZc9OWeg7u0aq7NnyjXewz9moVnhuwKZi1sji5UfX3NfpZnTAru2XXSTTyftld8qZzn1ZNOkDCQ
FrKxLnZSJ4+h4Pl9s1AwOeeCnX3gxPzYAOoLWYTL+uFndCVmGd0KiCGHbHZTx6k2iM6aFT741xPA
T6XYZ7T2O2Eu8jiBtNrNp/3JCAwCA/0V5Mo8RrMb1NE3xEa5GDvuIxkFEYFT+0qXOmX1nUDdA3l8
VDK3USinq/If4ISim0Fm0wYHaUXlrnfXu66z7gYZbcGWWBLoEdggpCef4CKvmXSmh3iIPc0MfnzC
IHXSqG2S8OzG2kAWf1VVtWp8dJI4WRKSzX6J9UmdMPVZjbadq309b6XFZiz9QsnrmYJLVTrwIC6r
pQ6HmGNlXCcVCklW7X/r4mhOu6aGFfng+6J0U+Mcwl39p6YP8qItt34CzaZuNZbjuanHrLLc0BTi
Li+yFHMcV3ALd8U8+qo9SJIVcjvV0rghua6ThxZ9UX0QmRWJ0x271lXiAluE7hdGwRJCMwrEbkpa
GNiHMds31WvRzD4HeDQEuSLV1w5u+ju8iu67wo2uvclUJAIfwBSAla16SkFUIop2gOqoivXKDvC3
oC62rSRWmWllrHXG+zPmWCZKm1pqJILU8dS00CnqqcGkCRjjB4SzamM8g6pLF1/qxeVFhAwvxwU2
dZcb/VZEsMbPMQeKuqTZcNBRbPYoBQl9npp3Cx/bSfM9UK09ztpD2RxTgKjWRurJeoTlz4//c6MK
tezclX7IvqpsI7zWHrPWDPzrvOZSrSXJWtNv2bjfR05OTi7+V9DgwTmJTxANbsIpqew4Sxsc0p85
hIqbKJNkImK2sBvkNSMnh3x/LKLIDm4zx4598+VQSqHwfgKiubUlAz3s19nYToFNS4bt1tzYBKEq
GDf6tg7218nBf97V4kXy3wk+60y3QBRLBcm9U46qrfnwqIUQ6jtXHeHssA00M7AWHR8AVkimlj3U
+aEdtyaI5L1iWW/lG3a3OptFnpNA+cXWBFDV+ihfKEVBBmDtkSUlXTPktRWAbHiLGGDkDdYzNK+m
bdoWq/e7SPwi3jY31/wEAE+dgJZL1EIRyHQDe++0MeGuwGL4wTzo8zuNKFEYwuCv5qXAndiNc5mn
lUWVBMFZscVsYqjgB4LN9gp3cEYPWlzPraDYfMjJXqh37SmZxLiE8thoU2/a5IQTjWdTasVjqT/9
JKFYAoTQlxsxVi6m1xTj885KhEkgq3/8OBXgH/W+OJyufT8/J5FbGvPdfP0NWk8IQvERVngEUhiR
d+PJjDoZCGiYpwDA9Y2LoQDc4wXC1x1RPNVLRNK6Jt6SF7RmcklaVOyUviZnB2O3oDMHToly7r4j
zB504x9LM/aNViZZHA2A725EJRcRd67YG+FdhpoXQbZCrS+qxN6+jTHKCXRrLPgw0HzA168MOVTK
AMbjDt+Pouvx5ihJ3FSuM++KC0dkWoe6NXXjUl+hGNl41tVy0dm/W2TirlaFaqx14oH42sEcFtun
PEtA53U5r+1UFwnPCdMU0KqH2btD/jKIHvkTk8P49GNoUbVgJmfTXOxCb3a/xvug/4KQvQbiuCpD
UVF79oX2evgam0EJ5xy75OH9YrPoo3ypvKbuZ0WExC2Y1gynBHoLNVlcZR6+FtQyZMFTWG6X15Nn
rnjKOoe73MQR4RL9o/F33+hzzxui0Xak5bjzb6VNBPGNNuWOMabqKOFqCu28NeCcbLwk94ai3E9u
105MxhErX9uqJKNlFw0cal7iu7A4mUIN56YBxao2A5Z0h99ocJysoC1OT1A3ufLO5ZXK+r2z2dCz
Qo2nCEXRx0Qm0cBNSYQnc7bN6CcG6xEnY8oYfuQy6cBwgdUJ3NwY1aIfTkCUjwbe5XgUDvowTTFZ
n0R8wJYNvukekLHVDptxqyZUK59P12plcViN1WrjDsEqdQC93K/dG0qCVtxfpSZW2GoDeAnvIiy5
CLrrP15Mb7gVQhhTl/c1ababpmAXX9uZctTx63iplgweW9hOiU53y8+mZWPcItJohS02eYyONgGz
lqdNtBaFKDP+t4aZvPo0OY1MFwztrtCi32od6X16ZFKHscLNU6Gi2oQt/J+7IPlqDPQ9hwMROFAu
PbLoOQREV9m2FM8QD4VDhwgPgfLXZeqt0l61kPO1Sd++45k363XFC4yfOerz4vxj+msHeth9+Pay
Ll8X9X026sny8m9gezGXvSAQRyhJE8ITBkt9ewsDoMshedZcLKhRGGmWCN08q7GdB7F+kbjajHlL
Q3h3UcBHuW5bWIIunWu3cTKfzSxCBl7fBjX7y4bQspg0eA5O+L8bbXNwSXv32w6UV229MsQkzsFQ
+1W6Yk+hAp04Ny6xinq7mbi6zErExAarMD9k2orRq6tKS7FebxuxqPSxUZ5/hZ7ksYv2fEvkO3ay
yGhq/+ZBjDeKyNqu+71rxpV11PlOzGyPBX+9atJpyLWM68yPKi6trQn4w7NmNB6bt9DZOOs1dqBq
xJnKwfgVjZjkEaiTuRHSoXVTQNp6CpgwwTfGzq4ozP1Oz0Xa/ftr9kXnVBp6gSeHQd1Qp04iVDfs
+RCtlBt1iPl6rc251RdtqT9ZA+sjQpuvmPuRjTUQaZ7C12AUVjbir7pmjU7GXyxP/oo0/EsCwatY
DbNk5pkQrR3iLQyNgY7gIIYU9I3ZKMNljsYE9vuuMbvpfHja4nCb/QphAX+i5OMO6I4fWMQbRbeR
yD8Owq+OpOE3PAPK3jsv7qFKMbVJ5ACdgydqWAAZpeNCSbU/0zS595UsLddHmamU9dVhTRx/DMP1
x0e2orwyiIHQ8ZKO2yZpTSTdcP+g0JcVEUTfkrZQ34mvkIbsKM6+uFNRggfOvjlMe0Uxj9S2zzY6
YjoF7SjO1gIDYaI2Lpq4AI2EZZbTfFc6/HYNcp0jiGMpt2edPyZeqpfWYm+ZQKAT+hpeQxU1bSdg
1Fob4fDDETxwnqykQUs7IuhQ4dq5Gjqw+Rs3yqHiGgFHesrBqXmAGk505icaiodrJZRNQ6uxwCNw
IZCPI3685sh5vqggdk3tiMFdiJG77+AURfbI0Xh5P8yt5+ZzSQAv0iqA5HUHs6bWn+Pna7LTMX9H
oK8gOjnhYyhXqKoB1sWj3D7LJCqmSiqvjjHMvsNCbFNED9An39sUqiJ3r1g/AZ2qGyfGvcpapqCq
oEdVBzBMQrTB4YYmbUyg2z4cmpsTTI7ALnigXIc9nQi7hknpXBdTo6bBomrV9fx3Ek3qZ/LgjE5V
dIAUmm6eMKpTWgrhu19SGPbqXrJ37vheq5ui/etFsMhmS1NBRNk+gdoIRuMbnrnRRiO2UfXkoeDG
uEIyY0uDm4fFfx1ocsRmwmHqYGD6dtTIWYQ6Ki7w+AUpZGtk8/M6m/tfnMxlwxZcpH1WMygXehnl
zlQPrwEEZagmYLOvG35DLfrNdMrVy6a26LB1PV3entQVd2g3bSTTsCYcEXQjaBaR9+elLtkoz78u
Ul569Sz6Pi/4aIIcYFpJzP5lrVwdjJ/Ajil3m8QO72Ve0GN4ov5PsUunjZjK5WaEeKL+WZB+7E5R
RkshmKcTl3U1L7wbyb717WSi3D1mfYV3eiSJd5uXeL13gLVWXGR+ulUee8/0FFJXwc0d3X+n6dCh
i6KDuvIGChO5Zt/0YeSYpbeBwfDD4DwtPr42tq2ctHlNkHvdirXSYhella8nJ1ZGjyfjVUl0oYlT
c2btjq+WukExP3tAkfsl9VS0B51eHCeDE+Z/AsgY3E1II3qivk/ET+UF2yVA4ziRBYuRxGee+IA9
UHYu2vQgEcqWNOMYes9hqjeSsU3/uVEFH0b+vL1Qi2Qzb3NHaOmY+Fck1QJrw8iRNQR0HtDK8aTP
g0KwEVn4t7gmGaq283OZQIyltzV8W/N9sP2u4cxVgoaBJ/uZzyUWp7cgfHFXM4Rsj9o9ozGyXhXp
kOGhrIi8/0/9Q/WkaCO54HJ84P23Y6XM5pPxF33P4ezK5/lQEVHvFufRIEeFHGbHlYiEVSVVt7nq
cnZN7BIieEVkJc48690lDIJvGsvpQtviOACiE1JGTiPGOz2KspBW74K+6LLj7UuyFEWLaucBlv9a
C6Ti4lmHyW65gHd2/36xZPOJ5Q4JFPs70QUyXKEu6mNcTBIXXEvCI+/HdBdQwEZdrjyTtnKALgsq
i7wuI00unAo2DPcigpEGmaqMu/DPjTJnZm7oIPPyZo/wIsbUhlvyu6suHTMCbn68NmHjmewM9eu+
kVyQnfkUORnCT0P+lGIqPIJe0BFw9AqoYy5e0ds4DPg+wmYW0VNLuyEHRPJQ+V/6ZRnQogy3FTHw
4p8Zs/prwi9rlkpZkt7w6jtoYzo2FGU85lmTMYqt3xb1VkFbCkCRI4iIG4dSux2d37SaQP32RyZ5
N0BiB5wlvF14z/3jtDekZodLZDd4+7X0zHDs5vyJK/NOKlupxYZ/u5ekLbhTsFwESMSNi0P0cyO1
8fcldx62op6x6Nh8j+3lHCj2IZw0/MDNAC+W7YmZ3t7qGwIZlHHD76TVi7v+PF9Q1C/QncrQem8d
BZ1e3YguYBjcp7KG+wHEzZsCmiCZWoNDpxLqyZ8UtPTwI14RzXCvAmhvs4W8XqPef5Yaa5qmISBn
xvkRapWqfWxeLy1kWeeS8oUrcVcIxuKbzB4N1OoWRk77MXv2acKm90V9deJisChH+Mlq3jWBr5Wd
FSbjIJRL0Dhtma38fv4rPq10QMwDn9Y5m6yTt12KQSB6qGoTbDaAbb+/2gOen7VHOaGkCemwKw9y
Kuh6aqSL7kyoy18AeJSN0jDto74GTQ2oRjxkMA8RyCGIbrc8xt3LMOIgZ2LAscAIroiyOHj4Q7WR
C40xOYdIM2gz/IzirrE1SbkcuvjDGYbg6/HytU0c5eBKZ7PKVlawMEraf5V7J0KPAwaTHwkJP3o4
S9dPYrzh2Bs6O+A4DY3ZXZkdcDiB17xG/mXc2Zqok7JyYEZ9JFHUcRpuVSXZ0AmrfgeZYK4tQwYe
RE+D338bYjYcVKOhygUWt4V1fQNzjrs8FV5zr2E4PfiaBwFh3Oxm2Utx2cGEdxDMp0V95tZFrhqH
4Xgf38Kdfz5V0PSEAN/O/TX0tXpSmy5M55B/VS2AursG2wK0jky1Zm/z9rLDbeAtQ2NgbVxNd9X7
3H7fvYygw8hV000WOUAXwFNWYu8LJi+B3JaxsKW1DTANL4J7vmvMtYSKVFJ4mZRLqS5bOvfqVq4a
2/Rcft/ttF6HiZOXliRa9jX6FNIFUCxCg6pvKDJgrkJHhfRsqE9F+GoeCZztlcf1RadpXnx4Qjqr
bGV/NoROUC9q0+1qNVp68AZZU2oCZyI9LN/PdfHNQJbDSMwztjn9XXkiS4LcYxmydunv05ERW9oh
Pdzgj58GlyYAPuv2fTfsETcPbLEdshW3SdfYw/GJKHgIExZ6/U3MTw4GaBSDzFcT16wt/CpmQ5f9
fwytBxSrusYezwWC2k+kiV+FvHSFN7XXNEpKWBSEa4EWsIwOW/F7NvO93McIZmfaInXId5rcEJv4
9f0UWs3cuK66LUYeSqTc3k+IKqx294wt4u4SH57T9mush9U6+250MSR5M2eg3egdYHnw3F5L8vDv
jUjJXUpHedfe6I4/sL9OHADxT8pmlRMlLw6eyLV7dCip7GtQOCf4OjKeot2JmANEsWCxod+dbtxD
oJxaG2i6blAXN2euU4ZqivElmuohXO1WCeES2KyQrSIqaSvBh361FQA8/Bk74LOLYlH6YITcIR/e
kYrlXWL0TfuTh7zPjMjTGHgSj3AdGfyHiYJLRi4CX0DjHJXkW0IL+gT/VZJDaAZM+LeIlntqQB6C
v8EAf3MUPMSRBkHQZ4NpV9H8velcxUqGYsH2DgC+rSlz1xhhaF+xDJObzPJEpmwwxlPUqeE5mYr3
y05qv0FRKIGeTIZG4/4W/0A0/yTOId8M9tt6ZQh1GkLix9flJif4zFetDS5fZOoSCmdffZLvCqzA
0F+bg2LmKLR0t0S9UpTKtGsVJIFXWymhNNS57to8Beja4OE63dIu4WlQUGgi4v1IQnYDS9/BbBVd
rRRAAl2EM1hhYid2c+dIc2i8nCIYQTfn/RiidkCsUs6yEZAw3YHIEjrj5r9kiNPecAJOENy/PmL2
uz+ULxr0a7tF4CZf6842wf3Rgb7BEs4AX/4Z1i2BuchQWx9XBu/UdEAKVdwIP5FDTvtU7vI8W2+4
6GZeb0Av1tUj692gHYCM2c6WxgWcB6gMwe91y9pm/iIDLItz/1mg2CFaBY7U2VEaRRvSz4kwHuS7
PLYEwi7W3JIGRNtKWH551qtuSfmEAYi8V2DiGtjcclXvnBlwXdGN4hav7hmxPpXVswFPDPoZaWD7
cKDyrTFOuzK0w+y8/02VoelRYfQ1NJo0lxBdWHKw2adPy0nXy6vR6ImWZbNPVqWfdyooI1GWrjBG
wMyqIsErJLyju/tiwvsqVJfXI6kk1tzxUPRUrButqmaRYv5OtQr6Z+kNPsLE2WiQV+onu+ZHJUzp
YllAnAD3usIcTFsvgP3kqRj5xCHrB3UZkwA9zdTW6RLXcPCffABNH0flLTInSBn+xah3s8N9rgfo
avOMQ4NfFE3vdLkk2WQoFZUISxE9JQgJ1xJTf2KdQdEJ2GbdoHFKB8oIgzLI0wiQwz6i8rfp0ZRL
px5PBFl1Prv1CdfkHCcdReMOXMuawR+832edgixkhcRVgBEmiqdi3RSdu2IvRnYTw/zzC2gGXHcr
5CgQUOjA2UmdrVys1vf4BZ8RO85zrFUTOFh4GNvf39L4S6UJ+6nCGCaWGSmPOyB1YNqRUy2sd6nw
875hQTlTxaRiIt22aLIcEZGBFKNeXbXV2PyxHJ+hKA7js5adtGIgUr1ZnJ9wi/fhKCzYspYxRm1T
abNzamDIBRLY/9FNGbs2hkzajIB8/qDfMxpVGmwOu65uLPBqN01CSpH4FclpFw/KKEsECMB17TLu
csVqeTYQy1QqjGqSMmwy0+wtwyMs79OvXiTrqGj5obwlZoG7TtOE1YkyYOsvkrn6V2jnw8GAlPTV
ZKzaW660dRhfWQDlXtislsBqlGAgL424bED+nlyaPf8ZztYDHnN8x0TGqoJ5dRNFOhKB+rOtTBrn
MGikExngrmYUoHykWmT2KUUUsJQdk2vFfONNnBUU6JCXVCfdipFY49HJkvtX/Ac9b7IILPNyUiFg
/8xyp9KSG8+ZnW0WIm+OQZIYheFBQB9+mZstRFD/Mndd9g/ApbCcwuNfH2qFoZIZchxrtmaO6w67
Gj15muBAaqm8dRRuwPIw3HOwqbD8BGrkFd2zTi6rMUdrAUCXXFWMyjnrQJDtKJmbIQ7VtPqF6m1x
dYovOr0eXMNtd9lc/8fe0/8grhwS59h9FHg8D/W2rMqAcbsfo4uMq/Ho281VeKUvTGXqvc65dGe9
YWAYMSzqFX9uKa1+cYZCZ4qSIEEQXGtnWaje3r212fBbo5jcBlTdf4+kfIpREm1qrOmc4SNlf4Ub
zBLYJOiE8UGEBz7W8Io8cDG1rsRem0yHKDDqobb3tiyq9KQnJ2tMefUOPQ5N6h6qBzCzDvZEZaob
RCja12vL+UsdTE/5f8sPfLlgtzo8JG6wR82H6gczejFe0msHtz9/xQQ6dpdrRKIKdi3UNf9l+BQs
4GLHWYxbs8vO4/npOL5nppCPBFTt0tt2p6U88g8RHj8QEX51V85YTpusQotDfJ1ehN1zpGO/LrvC
BRKk6EJOO1Yq77015ChRTF3ZM7+Ff79K0N9JyUdw2WNIyRbNnGgYKDzx5wqf/QItOPxNZ2jVApqy
bvR527jwCda3kyV0Yty8R4uJy3wj/jUOsteTYsW2HYeyZT4QZdRtpC3Z7kywC921ub/W59Qq1GmL
6fG9xmvxHYBYdMmuhxAI7WrHgfVcaaP3dBGib5FPMPjqAH5g91Ms8m6ojo8Py9NRwqjCaxiWYs10
twXwfNLYM26BYheHccGwD/YAEZEbJVTbp79WjgAklseEFs4RH1mVcFObk9xKkNByiLVR7t0+8cYd
cOLyTOdH9FeJSI2yDhTHecN7OHOQ9YIIpWH0pAWaC+YhYfDxv3fRc26qOY43lNzdvDkJfr6Chr5C
M5WMATo4HCX067U6dgDc0Fpd0DUnMxkoD7q58P2Zm6EbPWrRPJ+Ik+D1OV+GGVpNsiiMIWh/SKgt
OoImmNNVMA4SmxKicgPQh425NHijNOotk2Vi5u42nuWR+p05OMuIpjJhC1lbr/LxwIkkA2KOSxsM
W4gk6LIv0bJQ+80DMiEO9KF55hqJ8zLWkIgD53iCOzxbTZz6sxsVICijTCHHw01wHLm6wE+7g0jt
0EdavudF41DynzfPYV1ZadfuUejfavWUWyqTn5tGkvd3JfxNnz6DXovmg8aO3wlUVN+AY+4bqVuN
az67xK22S3d/cc5q0lQnUvmxYBT1EBb1+GvU5odBF1TtsIvZIYazgqwfamwob0ivcLl5rSTfM4Af
arLKkZGF3KKzFU5GaG4BbCj9UziJCac4WEiSChJzapFxGC++Rd4EI5SuK6brKr3akWWFkC9l7CgO
934A/87VKkW1nNN3B/ThzOZMWLQbuJFWHfFsLfIO1s3S41zT1AhnIKpinvlPD9k3RmegLUqKak5p
mQ+RicmXodyHEfDO6UToy3twBgScDoRw+D8G3mqGOyFfBMye03GJsxAHvKo9L58pZ2P8o3u/G8Io
cf7M1DkGVsjFEhQeNmCKUHE0gWj2Fn85eVN8JG3aha4z6yBKM2KK70JlwLVOPPI4zoomUobGj9D4
h8vf47XQG9X28cf0LymsTwX+TU/lui/oJfczG+DA2wKUKGagq30eRpGcJ0HmJhvu2VRaicwfKGc0
bb2i+ycl2C9OkHceqKki7cqC6wK2Eq2+gcJjAP/LBmYBrLloixenWRrbMmo+s7FMGP6koMv/X5bP
CEo7GxN8LlOEokezjfjSwjOhy6bMMBrLAHEzD1h+uNoAHJAhKkxjl0TOXrMhYJWFMfrDJ3JsS5My
Ojbv3jCpIdvcV9+L7vEKtCcjo1Xak4m2879dDljQVYbFxdjtFsyclnNatu6p65QnPFWYxvhKKlPo
gBl6kYDtVUJ8F0EW95Beax5a5gFK8it5XreLuvjLg5TWGQtS3yParphmfdnrUrZaL02k7BmxKvhy
D+BRTlMMLOsa6i/T0XD49Xvan/MINfQ9T3iBbVgpa+zCcATYb1Qd3/ID1B4ujtLZExeNi/ux6mRm
/G6DodP3puhSdtPd2Q0rvE/JuH7aQ6u+P5cvEGtVryW9QlewXr2jeYE6dxXW07+gxJpvqys+5vk2
TApMb69d8TE7T82F4kN7f16lLB/au5vrYJMWYKqlLdKIwHjqCx4lMPgnO52NtVJ8rOUkhH/MqocD
2UkiNNwgqy3mlBswna0EtjE3oASCdnRlZnQBfJXMkXBUURBlXn8yW15HGaWHFTdxCQmO4rw70vle
g2n+N2CpLIOFutaWJqcp4SnD1U3N0rgHTh33VP79cAGaY+zuXh6ycmNllLL43+KIuh86+DSceJ/D
599VXd78I5qUfa1zopVRDXuXgg1qEt+0btcRrFNj3XVTwsP5SL9ztfZtjl/akjUiyfiH9VZxDQzB
ntDZC0QKMQ6upIWC
`protect end_protected
