-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lw7o2fhj69MvEx0VqMUVez+le1hN3zwtL/3zr9cKveYDHHNVH7kmgzGfCoJdV+efzHyhutA3KzpC
bK7h5H0Uf58oUOK7edM8NTdFQmcmdAnx4epHWwFmLBK4BkJyZSD3JErl7mVCtWBXf93Ecqi5gHo0
A+xAUzn0XsLwDeWKj0pEY0L5aTETc65QKHmb+XiQdx0OJRUdeWGMsO7EnNMUSp+6/AiURdZNOU87
qYo5xj9XDQN2+jT//ushGVK1p29jEIl/UDQqYvpS+FzP5DBwKa6enDU7LbwvGA4xgbjYkJJHJMje
pa9aN7BYb1fEh1iH86W1fcp2OFJD4X4l9SDb3A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9536)
`protect data_block
gI/559LjKHJ0KindsSYchNzWsXin9ydFDj+ErHfMxyfz1tZ5gt7A578RqnPO8LOoyNmQTVne/LMO
V0oCnw9Vzd8JJQayCBXsO0wHMoRXQgfLUroTtaxcCnQMGnjRz2IiES2BrVb+qM4OjaoEGoYJlJse
Kp8wQ62QdJAtY7iNBsBe1wDsbi+4YOkwsZeSwySJrZygM2pNRMOaj2CyttScW4SOnBiZc/9SF/Sg
EBh423p1HWvUz33IGC7JcWUs8pYmMhrm7QcYZ12Q5RTIf0jzhDIgGxR0rHabNDCNgaNk7Ur4uzBQ
+Ch1+r0Hx2mzj/vpM8lrRkabXTecuVLL/UuKRGKTva2YqMw8xRMrVn5zMc0GwwL9GfYps+C5Wr9I
EAjbJQL90DGtMkPhQpd5WVP+I3EJ4UuvhTxjIrHDP+xG6sWEobFe/VvycgIGh7tJ2wuZ0gZSRTe0
bIwOVpMWe6y/JvzmFMAGd6WjFEt9+inGNwhP/Fq/5AagjdqLtEAXBSmtt5faLWS68ryvLaNM9jFS
0TWSXsIHvEazNf9U8n9naq3Bs4WzCuTgYqRMKM8HIC1klbIGoXA6BdoHMt6qQuPw00VB1EOwMCs3
ivYCvB46u906SW4YEUDEPiI5EJQFJO2VWE8dr7n5wQmRq18alWh72dYswMW75hxsfrLNiLI5i6OS
JNlJyZ02OHjgnNxy8LEjLNlQAztH7rjVHR4xPaeWUGGO/tptorPzL095cJmRUvSedGC/gwBkLKXV
NmP4s+qwRPLGnLioVJ4YcAjDrOmeRFl0scsrzB+p2fDmYxpyMY33UP3IUFvYdXaNbvC2hw6LbNKd
2KhDjf4GOrL3vSl/B5WYW61SumB0ik4GJkQySMJVEEGtd6beqx1Ozl5ukPrTVFWc8AnGIPX4hgVg
Y499GfmW9a5rF0G3LJsYX+lWzJBCOtjzJR7BOPlfi+73hN2Pa/eILLRZuFOWd8Plsln5znCKfRcS
jvlyS/USqooYvv8PwmqjG880guvWntEZVeSdw7SLr8P6atJRo8scVjr0aZAElEF4WGj869Q5ft+X
FR+z+PdnHtoXHtjjGCvctoC67mfhc/nettSqPMc42vr1Domov6BDe+WSQ9mhAUI/HqRqvc5d8U6m
GqHMbNXfkX8h8z9AYl1WE9gzm64SAbhwRH9LDGnaKcowk3cvWOXn5MOruVcPayKvP0S6vYW4cARl
20vULf9w/xdJQWBTuG4E84iw5jLWgaAu62M1DRUlKn5gSg2cVvB3u/uJTX7aS+ntkjOZ61RrZswe
j0I7BcijbwwGbUC1mKtDGmocQLya1HTfp1FwluKbeXgqsTqNnzscYJouhM+EG63H6x64HjIFq3s/
xAl30rQHbQP7R8pVCxXhC8Vnkj0eNLeCBP8amhVbQCWaAfriurC5MLw/2na62HY7OkKs1zlooIgO
vHirFiP+trNbBCAzs7S0f7hFCc9prKmqSvA85WLjyYW+T8EMZ5hf0Dwm89iWjJ4ftgOC/PulKJyK
gotHQT+gHf/UwG1xhW11k7wQ/ZeaR4O276S2UnNjqK9fIIUeT/EXTVFEts3GqG9jNkB/EvBbD7CH
4d7Mdsyy+y1k5zAgyMW9OAEvDV/mKsg3lOUPmqhICtSlWMVcEpB8F+0f6ybW23RNHA2EmJ/VTub5
+aMkNG9W87vyC++3SnPA7vuaFPyMVf0o8Z1Ms+bqKaKhSSLzJG08jMtrZqQ0qKY6yL0eQHBLXMus
zqX+bItAOxcaQlEU14IsknjF/58cPVlr3xkxMr2gG9GEjguXfT9y3LQdbMjZxzg0e/boAkIpoIYD
UF3gtCgkRaDfJ4NFaTnOXtGw6Z+XQWp5WC6RjgoWgaeJ0/GnhOnhtxOT1p4ONK0plqvyIY6Fma8I
DxF1qK5GLIr4oiSK7r88UY8jPSaHVh9TwPbArHQkmg3w0XCawAvoue2+kJHYQzfKUeDJBYvhwI7x
xlxgcy3WSwcfMjzHl/m3S8uowuFn58ohwPwf7KGG1mVHh1fz30PCyHZ0sf/E6yV3zPcJ/JaNalBt
nkUk4qB+4cMuyub9O8g82zNjqtOg2O0Is6nkC8mbR9G+Lqi+GyNehMXJVGcWk1ujXAdDGtTyasnm
nUrK6S9AcUcWcU6IqIEfJxlwRJsOTIJ0Es19VC0ttjlNbd8Zzfz1TTGPRR4YNWT+qDBm26+B856o
6agYQP3M10UtbsCVvwsYr69OQVSrs9JFRS+elfpf4bXMPKYGVL4IQMA4XMByU4dE3I7vVa27iabx
NVjX9UKVk1+F5ngDkSUMumEdHfy8bIzUgcVVWI3ZSppmrXw395TCUVCJOsE3x6pUzQj+Ts1zXU/a
fzeDVLmYCZHKTFjnX8AfV+jdUWh8o3nMbxHi/izD9HjJQ2bZCgcYF827QQkuV4HAk+zMkBrhilfg
Y0x/gqc6QGbhzOPFbUSVyOkAwD50BJTG/PBgVdAHGyQ7Dl3XSE+NEUKAGukUbvEj6EuD+DAzXBZz
IfaGwx4Na2n+AhdoZYW7cFquhrB3MFeu2C6lu1zAh5yR35PD6Z7msIcIOvNtGfLisWEwNsHovxP8
XuI4O8m/QoE9Rp8ad4MhveRcXuPrkHZo9oCHHPWFI9s9vI0pJ0Vr4RSlaOqo8LaAnkjF+kPkrCsv
8oJMjg/6niE/PFP9z1cjmkVrBEfrlE9knKPkhhhAOUNu0QLd61WFFgCJf5Hq7a4ykDYCgTNU5S+g
NNjT+emlR5REOnSQeFZUG47P94t6zBi+PCrGD6UEtRvF/lM9/+mrnIWcodrsTXr/7kxtsGXInrB6
Hiz9ciSesjn6IsatcnNnAklsfKrGEX0BPIDUH9DOdv+4ZNRvxw/uXgBHpXKGVoZP1SQQ99lZrgOV
jMAF2oSJRZXJgL3URYIgU9Fqhe3cKp4enTyV8r5ppRONTcgrq97sg7AYtwtiFsGVvvGOzLU+y3V0
MXqpZprQLQv7/vkXbRHwf/TzvbSA2O+dXrr+zXacJIbOHCbkjyT0phBtvmS0DC48sdqdBqJBXUQP
E10Q1Txz4V1sarT9WK/I3lhUeSyN36oUoOqZ4GwmZmQe7RRmTgIxrLi731CKRZ7a5JIohUP3K/Nm
MvDQvHjnfiWvrIGMNqYis+sdRPESq3KqOAPSNqyCUi2grkNSWIVKg6cfsPgY+QSNRUWfFrRIIJ5z
MGMrzFJQMZmIfHCvhOGLdNqR1rNyUWqSjVlv37nlom/lzRewzzx8jUBU3WIgvSFgxQy59PIWh4uM
rA2+uDBKpD0KHj8AMe5uoEc4BGVEHdwCTKBQFvKRVdyBoCYeIcU+rbKBVkRmf2djE59Vml3ax6z1
AcH7N1nFCgnqX61SHVAj8LFJWcKAJ8PlN+GJpyIDNVyhgQAtMQzsx8rM9XCjEb11AHIf/MKK0s89
U3YiBm6oeRhXuTjFgDpONN8zbyn+4JG3Qiw4tOrAP06Y8HErqHEvh9aJscNmybgjgQ5QsOrqxWwq
pMAyV/Q5ngUxxBEWwgeK225kdt1ZfZlQ0yMJV15hLZQUbfuvsi6DPrXTqFvCbWYppNj1hWbhQesc
6jsgq3om9FdgaTPwCpI3850rMg47H5QgYvcMEaKEaDiO99dGwBCQ9NJ3y4J71U2JyMM8mrAJBQCr
8xi8AxP5yP8Vh3OM5deZqP4P3qAPJLjubC911FlvJYJz+JycKWvCCVGeoi6cUmhsTkAAvZesl8X8
f2KbpArVYP8032SgysZQd3SWP/vybWahe+fHSwJ3EbaQmBbCVoFO/i6rv5l975ykLKwzKjJL7yfe
O5e1UWjBSpLRw2R0jmFgBXkBpWnk/g/A6bg1CsGkkz1vSyQFmOiyTih7WRVgjtWm4uNI1/iqljKN
Ki64NaqAyVdDYt58/iAZPE4cPYnmRGjWTiFoqX91i59MxIntFfNTGmdhsU97DiopZsLPnZSdUIHn
kL33lvvFx7/fPbkM5UW0xQF5Cmd1BcThDpTtU20ObIVEQJ1QOaFyazrGxRq64kmMZV1jGKZUzJVf
nOEJc00CG8Ba/Fd8CeIRKHH8yS7LcDZz/cgBiavbfDEpSBGgqk4hEWWQmfRCbRzTVIGWYfQI8Phm
/KNruEMwSRMxzIRs79NBmcZgSDSn9jKLiLHRTzvkz/k9BiK/2opNHancuMlNubR3AOVckr2Ws6qR
MCdQMa+Ta+OCAZm0VtSt7E6NUGiZPB7dFltgjvKNZXRyombmwQPn25tkUV+1V8lLXmdUwQF2aQ22
erAWAdHymuW/drXjOUS3DFuya3Og6EIeYLhCiw4XkRkmotfGg65nxxEY1JpTbKElm9hTA22ilHKd
HZi6ACLJq8zhCiZLerxMoP+p3e8ocEx112bqkS1E5fHUqX+g3DIUZw3pqPXdjAtNoUnfqmQNmp1J
BsQ97Ad9PG81C+RBjgC1w58jDcH+NIhJ+NiALMgzQA0WvkDk/9blHVawLj/yk5VdQ94tbZwE7IgE
G7Ebxat4ymUYGUMEOPIU9CTUubs4NU+SyP+iQ8gxgf5z3PUs6tJxmX2R7zTmZAmo969A53VZlTJs
z/cx6Zu2QaFjBmIvoHnC34Pn/6oEFL72lPaaR3JYRsBpj9a1rCy5mMqwp2DPwwu+etH56sGT5pEP
xv9z7YEbBZ7+osRP3hA37xPlOI9JuzKw4rMbm8rtimSAXmfI/380L8arYIOASxxlgmM2POHVaKhx
/0q/Blgicy1xBwRJZgGGALC/QeiH+5berS7MfebUimWC+JtdtKJdNw8GelfHsITyMGhT3jkC+64i
ODROlodZdkpMa+yW46AlT0KnmJMhNJ/38hq00usCNS6qUBxCRMidBnZr3dZFwp0MDRilE0T8u5sk
FMY1xFpq/Um5H+CKl1nuJLJINCMJg6mD9U7u1J7ofcFoQ0mTmWonbXleK9Y7+hKAvkho2QpuNQ6Z
aLYoywwG/mNEwFoQrYCmuUxOzOVYJbWiyaEg0pqAgpIM9AZPG2Dgqop7iZpWavdG2e0Jw4z58s4E
scyJU+Pn6qbqd8ImcSBQ08BV+eshOQQTUjyZyipBexB97vyglKB4V7JJvcqDJlLNeMcp8eYNTkL2
xaMiLkZ+SINQFbu0Gd2OY+h8HCwVSPhmJw+utJBoRQPQsHstOepxPvBV0unbiff2K3etJ7ov6KNl
8cP8LmbPe+8kQzOvOzjZqcX2DryN5QlIvnXWe/EjDgeeHyU1Al6rtykAwe6toFEHcVobFl3WfDGW
HwGviWgxVokSL7zyybO9xq4Pod5NftYDittb4vMr8PkJ93EceYGGFJF98JbjpxTz8/3NYUlp/IGW
Cz6NsnrAqG6Hxoottcq7I972LMQnE9YvV4Xqp7a0ank+lSGT9/a6OyQjrpvCvhsvs1JviB8IFnN2
G1X5bH7BVi88xgK4fJwIcTRiZO6o/35DXBSVOJph9wIg6L9b1zOwtysGi/NjY/s5yPQI75jMzj+m
wnd1E8Yq7BOYw/LicsOAPloWBwwyOMN+sXIgajT/550WWsHEZGYf3kgQKWxidU9Gl5QDTDnmI4VT
7AZ7wrqt/7z9WuyK/BEU22Sa6n3wXON2U6/yTN4vSxVFluf/rcZdoTo1nofrHOchYkxqTC59y8vy
YsBs9QkBac/27swbW4KFHuTFtTp+A0fGFa6actqk6m0jFxcVn9vGb3tqypIT4xr9wZjIajB7cl5M
NVMuzyzg0yPI2RmYEObDPfHupRY1LSziWuiOIe/Y0eZ7c0ngWc0RoIR0kYPVgyZFdPXkzt5mYgiK
n7iBJV4gaPavT8TbhnB5dpF1MsmcVNnFXpazXPvXi+KLi2FhhtaC6KzCdiExMiHPcTujkclyuWpO
NyUxxyag8RAEM71iVOZiOGwnWIF/OvoDggr//mkESWbl4B7yGkyAdVk5zA9mHq2lG3aN+fgpWYV+
4iMQoCNSZCbtVmIIf4ajRST4UYmIcwXYxX3Qr+R37jr5FqkQ+ruq+7orNTY72VnE2JWvwpHI9ooZ
QTD8MOXsT5oIsq218lFP4WmNdRIaR1TWWwMJ/BpwGenTDbcNhjlUQLJjf5o+oazDrsXU0AOIZh1P
ZP54T8sBx6kwPUOuhm71L2/fn8w1bNKQc8PAKXRwA79xWDjZ8td3DkOGelgbA4nNtxAHBU3N+ifw
OiTmtazTXPBDr0L/aD4s6qGZGBftv7m7wyzs072le/fIq96S+p9BPfGfPu37nUllIrTkaapkYDpD
Rr2PWfBcQsfl/c6fZ3q1gaCMZ3/NUySK4aCa8fojZ4veGkbqSzWS+i/DV1+Q9Du7OzjAlYjO5Jf1
HVCv+CwQ9jkQPkCAjgk1soxacPBKr7qZdmcAd4QPIjJWpv1x2MB1Bd2PZMlP5P4Xd55Yx9es3eX2
Ka8gnTSDJ7bG42V6XqjWHsC5o6mcMvrrL6TGdimJsQV/VGU/L3HUio1/w57DWW99y6rZTW+bOdx4
yxCvnufpsCnWEqrvmZ/DVxVwKraC6lRj5EuFG44vm0UcrxTu4fgDeUZWgyQlLYDbakBc6dREuSB5
p3c1NpgI2RMyRsS/FEfCDImxuRfrCmzR5jomIhhmHzEpSvFCFvGnRtdcLEYQq/+a0G05aebJXIGF
NccqjeoS12aA8s0UQ9NZu4mrOIQq1XV5O2YCbanwjom4tGdac2/65wMoqaxaooA15WEHr6jnTkDF
X9ZdnksPYHOIt84wV0mGD7Re+Z58/9Tqv3xaZun78/I/o9O14uTCEkjgoUQuQdAwHvkPO5WotukW
yRcLWmCUGWysoVCaTfCYyE4fFFnzyMpLyZ2d3ATf2StIZ1LAStpvHLsI0H+4NeDl/w6z4X0eHca6
QphY1IS4K44DQIe5vggizmsB9LIxIx7xThhNIEX82SO71BO1eQsQXhKz27T4oCePvqfZpq+nGiS6
XXXbP3kSBSepIVx2utGq+gK8eQNCUgrpy5zSibzO4HVcCM9OxpjCzRnaLrmi3qKAoe9YX6gDJCE0
ooZoCfWxWkfv4atdtie9vvW6MJfXAMdTpbzTb3QctaYxfS1SfY6dmM6hlK/H+dd4B5I7qz2pr88H
/bInxouRLo6BvQvnMoZaesbYzwNnyvQtpiKFiiaR7sMw4UpCz0OP+XDj+WBZC1jfUZmSCQU0BZQD
XXmmoGW3Wv8ASFSHNd68qVO7zR01L8DWgBL/jcsEcYuBQ7m2nbjWU56UT3z18ON0B18d3/Z9wedB
H8P3M9sJm+/uVxLohO3agk0yuz7E/aGBRFzuuGk4ZBfWMQUJSIBV3CZ3tFD5/gRi3jzTLhmx+rW8
4boVqHHQqZKBfPsOT3qakMEZ+444/sQO7At90nuyqRQiltwZUo7JQeYiPADeSAf12RCXn2qETyHj
0otzE+Fr8GQKIlH7d9+ej/Tv6VZCehrWbwNEJPVPoJtSnc1PG1tnFaDz4EPCs+0iSpZBK+JjXXIz
S6MBuHhIG/8GZvvi63dRhrxKan6zYoTzabZ/YqnqBHF7qwhqsk2vnDSrGNpm16rJjhmPiQ2dL4N4
T84O6OekuzZc2t9k2KY+4IM93k47CAloTv653z/rTKdv92iwsbSengPMiTg5THaKWbLx7XpLn/H1
Z6gyE8ysskNwGHtNPDIKKzSqlyZYfpjr/6BF1gHwW3kmEJzWu6GFZxTcUWgSFaJJlf0C0Czyj2LM
KmJR4OH0ges47Gxd2wk3vG3YnHdhNWcGnbVay75+Pj8O9nQagSmKbttpOeEwhLjDixaqKLrh+LfP
LyviSBmrLqmp55V/U/Qc5ONiqbnvC9CrjB35q8UokODZxMnYM2VcthCzNT8psB5CX51rN2URKW6z
IoF23W5Fu/H7WQoWPLb2fQiZmS78dVaWUU6pTWypgIxZaoSMgUe1ndt/8R4ECkla2Uc8Jb+tN6gN
A3dB8FYJzc3yRmvJLQKGrQmgF5z3vZU20ktOQKY9nJ5alLYF97i1v7dmNMcSdoR+d+tj7L1/l1tV
V0WUr+EJeQ1nmnQXnDAO286C4XQ+4juFM/az2+hbJ0kQaZDbmTztnnXECDnsFkEBvKHNuHTkHM0p
+ha07Ck32Ctb5txNyKN3DRZZyQuvD/AR0XfPimOoHn5PPypwpUnvG96aqdfxkyZsKae2Hqs6rU2Y
TB7Dwl3sPqV646nDlNaiYA27Jd8i3YfspXvaYSYtv4uAa6JPDfdi6mB7uXte/8gH5yOblkLYTOOk
APwHplwUnVIkmZi9PrSI6P5JdnmlLMlfwID8DissmW0MPHK7LmHe+J7cRvzKQyeh9oLBNmIdpf7i
5Aixb2RfBP+AkKW3spoWG0o1YwVSxVOfB8ntOD/kgHxHQH3HW1cIYJ7PoQUVw7VpwJAaRlHAcq4/
yC9CkoJyL4/wy+uvMZAg9oMYqtaq4GdS8pV/g+M2FlLHlEpXV7yCle445QILXd8qIO7sXIo5rTCt
4j4E2l7SHH7KMY7X+iB7QKaPqhm/CgnoVtZFgichaCquc98e60XdUiUBMhbSIZUuj3TC5bb614Z0
D5k+qQLUUmpoAX/VLU9qP3iW++NvBUA4wX4jmfXGVTawUr2B4VwwU6gnRm4bdUsfRoSrmSzAKly0
JPZKIQxy2DGWhrS9r13fgv/WZdPM7xSwg/vYyhrIiJzOTMSKtxqj3lLi3oa/70dOlMHa7mXqoso/
VYFnlYThgMVvXF+qWTKGaKuErAF4VbT9BQkIk17gx0G4b9J5AvQ4+R+GAx8VVj76tqG41s5GtR8s
obk5J+yRGGHh56LdSJ05f9hXBFNQW8CtlL7qqxAwHINf6KbfFytbH1HakYIXshReIcfqxq9sLJNK
jy5V+sqNKbQw6IG08CrbFJwpKScUw6b2CwKd9fifirKPHt2wMraTmiZf4MhTYypf8Bz2qdvQR3sf
w4l/niVLRnAmYzbJeBZHWzKW5QvHWKFGjcGthi1tVOkFcuhqg7QhexAxpwJc6Ni+d5J+yCqfjfYE
3/7+rl5v5SdL7b1zReUDyAXCRV7CeaDa2ZNJxd1EjJ/0Xkdrp0nCCnPe4qLdwMBWCrGGQhf66P8z
Jw7RcoBWD+iWciW9l75BOLZBCgcVU3+qwfSOVzAMvD9qGlAThp5swvI01X2qiK5mQEHbv0mVbFnr
SH2vHh1bASjZstIl51q5p/HZW9UcSiZgRsOmiX+J9BlCn7cmWc6TXB1NLWHhTgqlImxEmQ4sMyUC
24Xxjw0utxB8IbU5cRj0P18f9FYg5rbzTNtLGNUqLmsDpWbSARlWPL8blHK3CWYvrUU4kpJW7BAu
LnatzN3Fnmu8R9bva2E94GXio89qrz6ORN2ZulfBUE81y1iqMDSa93/AzMyuCxbOu0Xozh2vtzz3
JU4nIg6vK6TbR5t3ZXOQGtXKVs9OIUKsxybUJ04stL2IKjq0n7B1xjnZw9oV/Np3WVqANJk9kp4K
qEBskUAwtAEIrc1XYcmsZuUYQutada2SSkabpYQjfSUQWtrgEkMrKTsREHC5OJM8SOQlSz+L5RdA
FZzCNDrDEcFQfSNZVMgiNgel48imDbmIsuDaC2CPwhfO7kqqZrSZmnG5ERNU2RrXGIol0T5Z9a03
K3pUAmryrMH5kYQyaqaM4sI1OW4/5onhrRCcUtlWt+TDJ6DErmOA1OsypOZ6njx4wZSYdfK0KMLM
PTTOWx8BBhwfCCWjZveiRvNJKrj8zDUNfOGyBqtLepUrMSQNVQqwb3exxksJDAiuVM5rNn7dmiil
QU/7avr1om7CB+EQGKXHALO/xfK9dTn+UEyoUxHW2VMe4T+OCqQRI7kIS1rtftICjFWDJvxNpaaW
sPTGiUifFi5jePPNwHUAPLXcHaIIuzU2UCeDgy7LAapyWd4LJK1cyHS6/uzI/shqqn1amYGXVCEt
hqd4iNulGTbeDpR+PdxFAX0923cR9qRyx/bafSn6SOK/rB210zCO0mvBeEk9ZVJMcbsQQBbs04iy
excgMkmdnr28WbOBLnhlHb3t7U/uwPK8NATcCWcqhPFqcDsxF1DqpvJsDnM10/5o5TZHPzR5CibU
wbWbwEeGC6SWu07CfCZj9NwWMJAJALvsE/bXRflA1sOunpw5RpwcRcf81h4J9p0WHiaoMN/xe389
UG9GeioQxPlvjYCtoV3M5UQhyE9EdWopzUMngHpNtY79q1+9wi5FR9UmalFUbWZRc9nKu1mLdO3A
zV8I/b0+Pk3oAZt5mnZtsYgtwcrjTPjIU0f4+boZX1jAkQrMiuN7mw8qHrKHTUSIIdBITYR2H4tZ
1NJxMOtZqRAAXRhpgLzrRsYtK/x/Ok6H7eRDhlFGXbzW+8KiLTDzLvydG8pgQuHpL5goO18VQGql
PEjK+v/2IV935l8QUZB+CAeIrpcIwstpnZ5a98G+YcJPOoQC9IZ+uskma2f2995D5loXHm++MDeG
LwfGNeALB1y7PQHzSPNcER4uLUtO6U/HQaifJQKyli+j4culeZEWdbqQ1KgOUz2uaafdsFeulrDI
1knSrRziZpEfIy1AScux6rLRhTJJpnXNyV2/BB9oU+b2OZyEapP78kn8ZG5Z4qMMUV9SVKaMgWHY
jBZWX5mFDw503FaXTbOXYiNx2/yeash2xnEHT+MKvZj4huPIal1/FIMKy501p3vO32EuFB4pTAG0
Uq+d5RLEGLgc1h9xV98//ioRDhnLqfi8yqX27mk3FXbvWP7UCbNLwiqxh9FP08xvMMScjMr9wj05
xaG17jSLu+i8xniCR+zIa3ir7nwF3Ft6+5f+dd1eQHmSsEUJAH9FEfcDiRn4RNDkAh9//3ahMoIX
Qr63VNUw/QhO6pYyYA9g3Rj3+Du0H4rGmceui6SL73dVe1uf9u9QfzFzYPW6A8AtYjH1nHKZnOQt
vtfpyDOLLraoyDME0Aix7luB470khqOcrJH3+U2aGbL91OhF9qAtJ0X7huW8nH56jM4QGwPk2UtN
Cmmdqr9ojsiSMYESdxv0Kk7V/NmkyiwQ3ZEu9T96/RkXWXw1RS9a1vyzkEJC01gCxhH11z8dMpz9
mQ+78Jg5kdQUyFXE3+KaoWXRseLhMK43OxUc0S74cwGLeb1ev+mGFylpleeVl9+YFao6X5IVdAaG
OCa9cJbAKmSQzPlFe9zdYMjDqOn+sj/xkMq0WkU/a5h6af07qcno8lg6JhEzqpbZxThxaEJX+DDd
rfCKrNBvVeSyPj03G1qf5MsD80yPj+MhUNXigimUuwQuUL4E7lPPkIyGzSbInHfBodOX+t0r/fBU
UmgY0X2Jd8iLorg3qPhQl6HeYCQnEUgIQafqDYq+ZErQTtE1shVQvjRPZzuGkFfaPo5laWO6+eIV
UM3vYMX7PGg190FclR1563DoGm1B5a1IlYVejc5EUBp13OkKA7PvZWo85Y+weKFh3V534ndGQqqb
szSgBdNF97p02vkgIFo5p8f3nnf4q8PY4B0oLwTO59j8F/ENVYja1fOAU1OhAVPMgo/qkrNggerk
cL6P7j+fsnoTh6iZ8pvsxkh0NE1m16PNmpcpHCxgQPxup+kSeR1e+ZWY7/2u15l0d66YDGe6Sr2X
FLvCFECePtr+UqiXZUCgci0NzYjbuQjv2fN4WmNZPISeiiO1qD1tpNIBu0ppMsRqZzx42LAlgPPv
GU5lspXfHON4rxsGAQAdOD47bJHtGObPM59Srch3hNeShEtzVx/+moYlIrhfF37w43jM00eR7dFJ
C6zzoEYV9KtrnMkyK0Z5PhdbOFZ3US4CeHZFSAvLnVQTMoaR+Zk67IRoInRpr6SYU9GIQAWfuPZM
LQipNx1bWioyEfzIne5x0UMKIGWV8qhWRqTrOezRwc30vZSiEJJxppTHaJg7PMgehLDJEfk9Epgv
e/LCAPh+EUX911d7evfQPw/goD2vcsaao4q9yZ9Aa9fqTeEwYbnwvQBOqFI0y9vvot5opFTvRJgh
mVcfRMNmojay8UbWObJ8OrRIm9RJRMHL6roAuHs8OtuMCwxe/ow3ytCsC/7cYJ1NJzOTIGSmkNiK
EJZzsqhuSxiyyO6UPi8B7YJ9nkvnfR8zHNpuMd6jfdVy+bmyDAWZhzZkAZNsfYj11K4Iw+831wkq
jtIl/6rBAwHWZzPF/MpQf6VUE/POqnWiTVcltfkaeoMfi4y+JBzmh85kTA09/3NUNUsFiMhMuA/w
tLUkwuWGHTQH/6Qq0Z2XprCTa0lpk/mxMHZiLR5n96jpSb8bLiA0WzEKNyRCD6PLcBbFYoxMhH0D
xm/cMko2k3XHdjellQtMzUw40432rVw1IAfyQrVbWJutHE7P6QqegDOxfQG/+JI9ucLTrbOKjiX0
uEFQFL8lICAznCuMGGw7pd1YkXsFAb2QVlyc4kVurILPohehitDwa72gAFfkEcYgo7Vmwvcdoqd5
bUWp5m2EhIKWf7t7PxgcIAIl+VsfpRhqXLeltVg9VTGYmPTK8pG0cwgzYDnv9aZdzLfaF8lcBOi/
AJNVk2uopUYulQDmZwtdYu2IDzZXIdQXBYqGFrnvUBql4GiF2LMEz/v8PnvFExYzmIrZc8P3/S/S
DHGdCkz4kQvqxmKGTjdUF/iU/AQfBSd6So/y78UqnO5N7TcByNQBoq2JDyzARVn9CMcRfea0mX6v
ZFIrqDgz+Y3gXl8VcV1MUp223ycMHfRSnNC+6EzZRdS+5Hzb5RIPCEBPuKdSRaXR00MlgazB0eh4
/r/HT0Q2jWOdj1xZA57nPhc=
`protect end_protected
