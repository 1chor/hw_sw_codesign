-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
+O4Q9E2wl9xBapEtw8J4R2SFgnxayS1wvHccsnYry7HMbcV9o/BmohQKgIjAEiK7
k8FZM8YMTZOSLLBNAVn7Z0f5FKFNcn37AIlyJZ0L8t1dhH8vKw6ZJflxZ0eCca28
8i3BgfemKFD5soHhFaRyFuu2oeWVFP//eARKRiql0bL+xX9k4Wr9cQ==
--pragma protect end_key_block
--pragma protect digest_block
e7UN/sKqszVUOEovPDfmWD3vMlY=
--pragma protect end_digest_block
--pragma protect data_block
7PMl6g02yGQuaoLLiVWCQHSr6Krj7Kdp9KlW9LKEye+D+BrJUeTPI9PuIzueS9wD
rvcC1qdL0DsEmF533ndoJr7EliL+dov9LOtdyL5qwq4yIqFO5a0hxQmGhTwbzvSk
oa3DChBRL+9uKbl++Md/6Pu5Uz9aNZfp7mwPU2nLBX3yOCs1isVa3XZn++exeZXw
x1lct9EdQjuSuEWiaKpia489KgeVmCKhjf3/QRo07flpNZy8DnHF8sCwUkM4/JZS
IXPtaV+eonbm2jaYtY85r9iHNZ+FfRpgPP6eK3IDlcQ68mHba+PZDFr07j4u6pJW
SuT2a5rQ67ImlUrvmME1QqE3HFOiHktoKb13oIqR1lneBwVRmGZj8Ib4U1wh6Gch
a/jE9MikH0LJwLHQKFxVwlUmp4LjP5mwkcfVXT7Vw5LKxLt0fIXKh9kwH5upSShL
bKhkLGd8bV8O7tWOxzvkRs4Yp3W1Kvd4///Uu/EsmIY75NWnHO84lTfVFkVd6iuZ
2mQkP0g9WKkAN/W3Dk3eOr2TIy+n0PgKY2zQTUQSdlvym9opshxn/LRRpNSKaZ32
HIknIaLe+VyR4aBCd2UDJEMsTTw3CRTYw9LD4oD8zqGiH5KOtJ5TlVwAOApPcyEG
/ha3aXZ6Bjx5IWanlYIU+Uvbnlu6R4LJiFU6xSXHDdxECHCMG3opUcus9cJNMQgp
yEVbGsWTnkqEpN2jpd2UuSWQXxH3rsF/BicSUYOzVy5b3vrJFgJ8asrbITa/NOWP
dPIO3tzYbDefSLQstKiIrsP5h2ACTD9d9SHgOzAnriQBnaJ9KW2bj4ElSMb3tZQB
hvZK/772TbiqCORbM4s3jL7ADZyAeWutx+svySxSxCf0DAsqG3UejLg2htyEc1vw
EfzrzzblgQhD3G8SZASKa6YtqTAum5Q4ORrWX70ZzJqPcAK8zNLiiwy8MSML0Z1S
5HTcI7WSRt9i20OdujtVqGT/lSeakmb56pVHVxT5D0/VVz0XvMGUH6a0bDEjyklR
xmVhgm8GP+eSGqNNofzNCW4G8RyjGD7/ft2VbEiSvXElO+48RtxfGr9LSG2IhlyP
TKvlZThXgbfF+5emTLalgeokntd2l5ed566j2ETJoiUrusyYqTxrGz6fvwWRuDhS
OB/aEXVCVeJRAIDNmVICuf3sW6M6K4YBUVt9TO8zyFSgefNFEXQ2PC+d4bGM12t5
Vx+q9D9DmYjyznmGYFUanN8xYlon4LETa7kG1+Cnpy5EmLvuLJjh8p0Q+MRDenlW
GmJwDiGs96cuH8boj19T0D58aX9IsoGkRfVS6sQHqaxrQWN5TZgmpKkBf9n3R5e4
nmLxEe221k+tSpM8OE8iA3zsfA5DFmRTgEEZaE/g1CAOT7MP75rQrjeHPoPUtVcH
cG87hWQrb86tZUecqxs4vAZ9Txmn9yQ5114IkTYD+TBz3RkAKwrBW1ERnpqJhTMi
tK8Aoi+dP9e4hNrJ0HPgMNSepJiWojB6cTVF9T8jZwl6aiXr6rDnVF3DE3H17CQ3
IkvzSX9o6GZOsBhNulxEkwQgJADalUxKJtaT70rXlaPFp7RI8gK6gtG/esykMbrv
1yYdYHiHOZtfbaCWnHUfQ5uKQY0p+I63SUU2/HMh+KlgjhmV68F8U1LK9Uy9pa+O
E6MtOKLNgZm2+22faFvSFdi5qphPqWlwE45tWvRcWw6VVYaL0nhSU6dA+JtteET0
0lOc7y/Dutjt3AbUQBHbe5eJd83TAqV+b4LOyvaeL+MD7x4nbumKHOYJlRbMtP0x
w2tfjyqxCAloQ82UKll1AypP8Z+L526KeFE5CVlRUwSOVp3ivGKbQXuCvUxk4Nag
V6YLOkpRpQ5sNVGGwASpV6Nu0lRLmgHv4cVQ+dm1Bow+Y+XgqwdxxP1EhDoL51BH
KIG/DnCsQUX6S1cqJE26Cn8H7gyB1qMI1pah3hiIku+zA5dlazf+qDqQJ/GljqzY
1FoZeMn1mtnyIhhZDmZLJGti52cuXWH59Va5h+WJKsMCAY2x/FT02tftrd+nnl6V
RQfyCXoxWskHg1yiLEzcYSh0Jqh1ZqChwivB85rzfDu0ioa5SWNAoXJhk5AIhuXA
Nj2KBLTzSUkvcJPoGhZeqiOsvWTMrlEn7Muj+Ex16+rZcF+XHiyIc/9i1D/I5JtO
I5gnTO0FWJzaJMN4xf72h3i5uqrRHqf0KZCCOLJL2RW5Xqe91BbDvz52axwRhdB+
uJik7SWCPSrBfS6amWFjUpGnA5ZC2iaxKupHuefsTSs2RN94Q+ZXz0BbpW8CPLt1
N1cF2aodI4nFwcm6S9oilKpitDXi7xUaQpSXXFLiClD4q0p7XdRv77O4NVfr1Aoz
j93mEtDPn5yejZ3CEbx2VOMnOQQztZBWD6BdQKyjs9y2S+KnlfxBqoMz4KkYO/eu
hqx+DVdwMB0xaO42m85eyDXVy1emxQvoGzADd47a28T+XJqinyrm0qpUXbwXAle/
4kWmeEzO8mjGoRo1FT9i4WLiA/GDrySFmMNPeKn6nEUNuyBT1DWIF3wDXxBUC+4e
etfIjGlnu5QwCsmbpm1uUS0Xr0ftIlpagXxg7plpdPzY+xuh8Hzd30XncRE7lZU0
pJC265zVNgANW19cj3W5WkFAidgVyTT7cVdbljqeT1Rz6dMMtIVTryFI0GuAeq8F
0SHkMyQOPX4TQJjwaxqWEZvmXLWBDsNMh9v9fkEBp0SlEWIdHK4D7KkXOYzW3s9x
nMEzz2CYPEKjt9JY2SGqYHuXn0b3+/T6RRFINU4D6LW9aiqNGwFrFUhfEJInWZ5K
aEA1MA3HFiDtt5kVDc8Gty3XDDB894Tj/qH9jZC+/REMNvjSLXEnbKR7zi9ifk/Y
WIf2XhKUsaO4ldSTDvkg+h8OxhjJKAqJlUcy9duYHVrZtglQOhQVo31CLgtA/vhA
QTry05ab7CIZ8SPWzsqm++tkqtsL8d5Ye2p6ecf7ogc2fJXYJE2uQ1KSUVJHnz0D
LXDqrNxiXjP8EdisKtBIDPpCPvmqL3X+0LtbeFWhno6eiudL4ErWiHjyH1efDEAY
CWhipgvlNkYKS9b+h3GI+DmJNJW/irR84xxt6qFeonid8LnO1AS8sdbQcleKXq+c
ieajf108X6xUHH9w7hCrarP59CtMONXsmBl28XS1ov1HOGI1Le1LzKyVP0gr0I3z
b2u4IQ4CKpqfGhSjr7kyBYzcIDieAulhWmtbt0djze+QT4Z7BjqmJAkR8qjLW5ga
xyFANRRNFaXGUmJIs6Na8jbNCTZABoIJvMg1Jz1dDJv+e+37GDk/B1W94jJwF1S7
7R+5qfJhBUpSA7v7hS+bTMogFJJLmnyb2bTTrJ6JTJmQsJHT84oFr3YsRRmrICNM
ttYPDVMHIBb4VtCXnJId+8acM/r8Jsldphx3kAWZmys0nnTPQ3Fs/hZ2sGKxQKBq
w1f3i2OekYe4GXNuQ50Sj+bs8wbBf6U/j9v96tv0/0zBx4XNKsPkFfw1SEmb6mSz
AcRQmEOMXWFA7/gacqIFI80bu5EEjh6oaHbmP+SkOvJYu+B92G/MyAFrSQW3aBCq
YzQH70WZoUoqZRD6Ub4xt1ueMofpZYUnPchiTlXFUGJ/XHRbmOJpYpME5tMhuy1s
YQRddEoZy3HeX+IjTqhfNttuQSnpFadNunw13LsUWnk21MhELtp6keHPSAs137yJ
O34E5xJ3oAiPpqbc6EdHTH+q42b0i7wEnreoVgZt80lW82lQxneoIBJZhSOrXKaf
JWKpt4yuYKeWekXcQyRp0va5hZ6QIc0gJ58cgN6Qk1Lt+1YR3tJoX4Wv//Wza1Zi
jBrcgKpmYV1QBg28Q72MLq6DgBr0qgrTHx9HN/2QnPoH/E/tOrtype3WsWINDWO2
6lBTT1uEMsvZ4s7ZaxAmdKoVfbupJHU5U492XDMGUYpEt2b3xbpJZ4RS1Tsu3KDJ
njsJI/h6blOM5b/RZt18MVTYuBH4xGtjshTMlFS6kOjCwKhmv1EFtpD8U+J9zTTe
E53MYxIbOLGvjaOscgzSO4eHmQXJV6yGAiZceAspUCNjmW38d77A9qZiEzt+jvZ1
TU8duHXOukIGGlzDHpGcQ2K8Igo2tn6Iy5s+HkzFwP7RYGit7rR9puFKuAHH0out
ycUJLKI7mr2UeTleLEcIrppMbH6627fgCPIP1rkAgUbV3Zq5aT0wMOVahBMt2gOx
BE/ATPAOFB2zrS5uZrAPyx1/5Tr1wTzKMa5wMW15N9rMp2ItTqp0P7lRQuDHOZ9C
KkM9ULkz9tpBrIRq4POzW/SrCA61nmNE+7i889AypSDUe+JANONbiIosvbbKtBMO
f+KciCD4yzAOKPlwwgtqpC7wMlUmxP0tscFmMyBpURQoj5a1s9VtvsB9Ht8QG+Od
dSoBwnb9frEtlOoTcpLdKvZpfFmxJQDiPtnwGXy8SP4t5Ew22KNc57D4jcihY5ag
V7jw0kRHUfqfU7sogXr94sIbnplWSpC5yA9SNAoLRQas/XFMKd4DCKvd4rj9gLIq
FHBaTEkLUaNf8UC0yw9qMt55g1dxTz4QBB164sZkYrsXikA8yQC2ZyWFPa/a/qQH
chxBhB2Iw3yV8Q0f9A287e0io0Y2DP2ZdwtF2MCJe8HNVl/5P3K3KXLyVQcc1max
ixIiEpcnZQ01IQjY7wVRV98+ok3LC2oFZbSkluTHMDrbVLdtHjsoCu+57trIGsIw
tygQbj+3fEOtRoj4DDM3ejGkPHcEiVdOqh9OmvzrGDIi0mnSY69Acfp5VoMssgu8
dZ3svEKPKX3wmvTVtabdNKQ90Z7d8dCg0QKs+65wfdGOIz9fxPyzhF8t1mBgkY+R
jVmjjLcntQt+U4LGoRD2vnBASVfiUlB7nY8nZwHFxFl4zWWXNI+14uDCcjBoT88S
OcmMiTQwoqyDl063GEXXVVRUsOPIVVb5Q16837EgC6Hxb1P2KH1YVyejDDPNMoDg
tBwcs470a7Yv4u0lmp4ktglimfGeAnYCCp7hqE1QL0UqkCarEeawUnlhdS7ufGaM
wYOlIwcyR6p9ETtFNhX7NxUh75gNYDEI9qxtuBvLHj/IIyV80/KHoy7jZ0XABNuf
PVZPT5NUw18Zjik1vI/7ztCtEZi9l4DIZKErxqbEhARJ3CrLSqRnNYpgFFko0mXR
IgfiRpEJ3GMsXCl7nImkDTbvbUFg7u1BCttNb5MbQ4pnNr5mQ8OdUK2PQJZ/I+I3
3ErrdEnhFq7FBwvlQMaZXpfES66hQk8efHd7wo3c0NQQhJwniarzKHi+RYFbVajC
6IhizKjwrqSh+EXvdsoRsbU62PO9jwbb5/4ViRuHyhqdXJ3skFVaQ86FiJGv0L3o
kAFiWGHRj7JY7DOFx58KBcUjE8SOJip9/RZy4kY/0Y2k9RM1vW2l+pE2BEM6DLWT
+NizlUbkMPgSwQEvJjumuBM6UmI/YrTTvPPfODaj0QdTBh/a6/Fr5fz/ofvsktB8
1g5W0uwOr1IpLpT6U6mffimqMCSTW8slBOfMbhz5Hmd4XXEsUraFjCCSbx3yEMHy
W8ia2oDWvXDuY3tlQP76kg0u2/fLCg12f7+C0hGRuBbzUwJRtaUq6KyYu13mVciF
rqO2lKb0m/+92Bp7kvpTWptt1H4aSCsrcuRpsFFKLH1ZIeBRGi23yPPSH7K/k10S
sU2d1GX3Cx6j/clrnap3lXig9ziN7Uq6wd+c5m75ZoXAgf2stqTPRWWNg/Hh1IYH
rOVm+NMovAxbqy3in7AWWG6xWGvWFzA0ga9J4T6U7Cb/tyj3E/TcCUQvzKtl94zd
xpAT/TFcVPxowy+IZFM80ojgFiqDEZt2tSkrhRMdAX4MDsQ9UOIKwYHcQG8adPZW
jQspaDkiyssheKSRTcnG0jvS1zB/moXH8FYi3TH53hphVRf4SobRlHlDWlzUj5yd
V7YZ80Ir41iZAsp5s2/lm/9YoyygyEFNBa5Cqto2fLbaay2uW2vyl8JdAajNFAa0
LPXKoBZ6eJ6Po5+tRM3JBimn0Eo4l+v9y02VdlIinN+r8hweIqnG0ppWwJHqOLyy
ePvZ4G4lfK8yOB8sWl0lpNBXDfQ39tcAnHBjkMNJhY/jXjYQZaKhAbogp8z9yiKE
T8a0nzPibwcmEU7wuOa4QKkJoKNU15sbo8ONSxtmipUqGxvKcDW6HxSxmz6zxVEg
jyIhPeOCBkIjuGlH30tXy3nPuRJcek0g3Z/9tSDntvDVyE9NhJUlmq9ofJFRw5gD
vSNOOs9NXsmVAcvNWgu4sr8uPS+Jt/38StWXFVPyBBYbWqyMgtjzYEX0Q5vJL6fp
h17ywnAQI9F4BMU4oU7Jda5rU9H940oOLQe2V2oNTMNPEzyiMl9gk1j3C3McfoJw
LdOo5sHbiWkpV0hEQZEgb09NPjXZLFBqQtp7pG/1Wv+vxi5OFkpbpLHPE4Ev1/GY
6wW6AblNz7svnuWDT1pBlGA9u1+Gp3yuo+NRrPdiHHseuj/a3ug9rLqxk46SveGs
07ejj/KP6i9KoSkI0Jeb4fu7ttqwDR7TlVfOEl+M0/G5ETd4rZVP9SZ6KodhK6gb
LZP2++AYkTO/pIu6MqZpu14yjF3np0ESDsiv61iM3Ukr0PUNsfGjzp5Y5MUdgKCh
0fy/FeFeneiYOtWtmO2r3hHjlxU3OHvvHbdwrvEVYTijUfzG1Rw7jv+T3A+DmAlI
uyQen6icQft8xa6X7p1cUy/fp7iXqr1hO4cGjGl8EyxegbLGjqzWvP3QSMTgPVH1
lfFFIse1asqPQPCf5AWdeHhHc8eTpLQ9dJBs9IcGcQnOhl99qEW9jVirnKMZWOL7
RwI6/lJAOvd1mIBDFaFXJP8sOZg4X8L5scLMiwot79mKVQNlYXNPDYRhm9U1u9XN
9QMmjVoeAKLoULUH9lb8YCQOlJheurcN11UPwW/SfuhkNyM/Mj622GxYdbmHoy1D
Eyw554jTOP19mQtapwVtypWaot3xFdxLrcIoCTVUPsTXTAMIA6KkfCi2EYaknSA1
VPHb3DP3D1lW1A5jD6ts1XEAqp9+6FM86rkbPZMEFAZP+xUO2QrVF89v+Vgef+UQ
QjHd+30qtazEWetChcSmr8dcUbXxuZZYoL800YBcj7IFPK2Epb7dZl1lZ4vxyJ4T
9XlMnWoJjQSWwcX93HXYT9Awtp0uF2PPNVRh3FssbymNqOXBpSRa8D97ZZ+T5+Xe
popPZ9mewBZd7AuM8yWcZ04j1HTz7zMMTDae23FvdHcVVdnU02pxADMGeR3rxYgX
LPXl3M09ZkNhpvoS5wNwIMfYDT6unwOkoA99Y9yDELIheCUYNCIgxidJ5CIqjqS4
8D4b1qy9w64C5adzrMELJ50Cuu6d6k43cts+pFF76i82le+yPEAtlXcWdz+pV/iO
FVY5SXNfb0BiOBZKPqbxvRGJORVvK+Ns7vapImzHG1FdynCHlOgRsQWeQzfJWBRE
LfFxLQzwF+gEQe/NgxZMYqBm/RUik1nZgckkZyh0P/r3fAz1DLwqfmUH6PNG87D5
RPIIPqBu84bIO/J8JSgf4NJIz4f1bZfh4aPilzaXWfZT+bvHFQcF1aKhSyZDeKiG
pZ0bPhRrWZSTJHtFStnfCcDRacWshrq3bwVtaD2NwQpbVHmaLSEgC4cqGPoD9qcu
B1f+jAt67t9g3d0XiZIiQTO7nWR2Wpx9S9PNOgCci1y5CCvUCHTitXS3dbS0p5gG
nXAWgRrWG4PKjcscT6RMjd5mC+OdkTC3iMMAtTsk4OPWOjCVu5hd6Txjpj5hWckQ
ftfchfQHSySVob3g5yi/OMn7dphm00fOKHFxZgUXGH1268wqD925D90xR83zLzTA
D7e2XI+etoQhNXbBHMJeJ0Bqb+72WqGqbZ0vARX4rLcpC4W1t8wdeh3uAc/CyDzZ
4/ehkefvYSpNYW280MdzDjKvb8XTl0GT0STjvFBQZ2y3mHaVzjTndD9wifvxYXDG
ufJ5oSXyo9FLRZCTFHyGC0xeSh0J67tnlx0bgbbmPpp+QvILxWOhmPh1T/t6GKkb
6cZhnQ48mJvQxxFhgdvDk4lOdBeLzcb9AddQjZ0N+RZFE7aZxYFbhIVJtFZmso54
y6l9qtEpTg7rsgz97eQPlsVu+gBm/4f9WlJTzhiBt5GhSWzKtjbEXOljRpL2oGkq
FWvAqDVXUSLlQpIm2syPSIqEvtzVrWrHp+6QR6Qa4xKuZLC9J/AOND5wS3+OlMTM
/mUkOJ3YLjBbt1EvHuK85Ix7kLn2P3jciri6poTeDC0h6lzLFTLbqp9yHsaGr/eA
UJy66PxoyamiP9Gio5put5sjFn06P0Bhf5Dub4Fa7SkCO0DZ+4/UI6kkJ9aYetzy
4xeUczj75qA34Za2+aVr7MG6C89wN45pn32ngvd32PkQ6VbdJBjzry62KOO1MV6f
MTLnJEUZVPOLt/j5DSs3Hui7RJwDthz8DCshV2r7H4pPH+oI6XgJ/n6dy3yLy1cj
ZiZ/jpQSgLm2aQNMEh6MxtKXPmvwW1Da6zhMOA/IX+xgkHstjah8vqTRXt0+3Avk
5mjEzRTMyKlpt9WYm629IbDQY3F6NVES6IQ+T3pDgf5cD+69/zLHJ46rIszHV359
5ki1Rmrl2snHaegiu040Ncvy30P07TCcudy8Kq5f3zzVzFnvvgPbm1XIJQpOXoBN
SQip1xDacLNFcwFsRUbU3pVBWJ3NviFlFYiGfcN45VgtVFNyVaGYeIlkc03M+krr
KywXWkVEUJp8kcxke6c+J3OgX/sgbpyYMonabdSoZIKqG2Da6dqsYgfZI3/1ZTPl
7Kmy5TlSc5xajC23ZKRABcuAf9FqnouEDkoLHspmVBVde9FLAK8Qu6fSOD0aWjFm
uUt+yKgoIT0u/Vo1m1RZ+SZRr6q1z+fbPOW7M5AUm+8Lbo1rgDy1DVfuzCwYJAeN
fIU+9lkjb+HsghAG0U97tdcmr7RW867f4QMs5nKMvKteblnXwOPnxU2PMuVXk6Y/
yOHTyyLrHNVim0nrHb53t07snGDWwq08XTE6iiae4OuJ4kn47dgrXzucP/AURbyV
YqWd1WwEqLtjgjSmvZdBP7hPbzc+AArezTlK8kxxWJT08G2ZsfSBUaJrhAxX5051
Ms/AdoqLaEqELoW/LxissgVFy2kl5cETBWP4TtgllTjw9ShokfY77cipAO7MiRvk
wnhZwp8iOI8zwqgXaakdIlgeciqsE6kkgWopolMxBR4Mdah5nvCehtKHcpy4w2v4
ew/dNoetMfoaT1kPXqxqRjSjGhxILm6JUm3Ciy5TrLuwLhAhwMk+InVB2DGvhlsE
bbaOBhLHegH/zofAZC8WA3hQEH2XtsLyyQtFC7NYmmkGRXniocQYwCJLbd83DiK2
NyV5jpLdo99u21OSnnYPa4KE6174FIeBWH4fLKQRWg5KvSMIsLMLbCViGzK5RR3r
R1z0G57fAczLzZH+hSbVTqXmHrBuOZlWhd40Gm/BeUs+mwqMToTTLCgvq4nV9UCJ
e7jJYgmdZjLbCyKEd7yFdK3WVzg8lFniT1J5rwrhFe7tbBtBKjGrfuND/Lc1xWqY
fr3QLgiFcRw77xD0bl8D8z9ut5lmHr9fd+SB3okMWCOvYWIeCGJJvfnc9T4AJPH/
1obeDep+imz3XBmtbgL9mx6EUtVl8t2SrsCif/1z7XMA4TvWaRFRXeQSR7Hca+ne
IxPHHtqFWhm6wUs8u+NLbbsAs8eyfN3dVVUlamGys6apoQ8Npf8cUgW11CBGdIQq
T/A/vKFte7toEE8moaOV7J/zZM261D2rc7y+9OeM+/a+ibHWqw531U0gFKWCB8HH
mE2IJnT9kiBK6I/R/TFzLTl5g82fQ4YqVjJuAzzhZVpodPTVsU+3b3t+pPm7MHVv
62ObR9b1uVVlWmp83G9n7M0f5LampivjAsUDADnqdYSJfBhppdXiotm9oNkA/c/W
qN3MztFqLHE6DgjkqozOzmsWvMJ0WM6lQlg8hADvcfN12+9QpUmrXMirZ3OQxQ3q
cG5W9NkiXQYGcUWZh07zrMSQ/a/zO6FqdIQihJZL6c8+tJc9zOqgC2MSMO/gn5n8
JkEKO+DvXXNwtmD9k7iYZnSsOY4BPupQbzL0nzzXfc1Rs/XBqQ6IAK0fdbk/eW4n
cB9bzl9WZA+tP2fn1UZhLAk7GXEWC+XfAaQwKZEQan8T6G6cPCdVSemkhP0bv2EV

--pragma protect end_data_block
--pragma protect digest_block
+9cFSSd4iThAsq9mV/WMKzMjU1Y=
--pragma protect end_digest_block
--pragma protect end_protected
