-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
XYKITBhNjItmaTX3NnobSDqGs0iuBAdG1GIYWJuo4qb156oxqOfGcxh4YcQHmb2Z
exlYskHCoFuGlC8z4uBj15EhB1O0soXe9Mz9J3je8ixNtrIAqehn4rpo9VE9TLk+
dOtn5QOaRmlB1mXshOw198tKlBL+sPM/jEIJ11tdKncu3le3UJ7kRA==
--pragma protect end_key_block
--pragma protect digest_block
2v2MONBF2klvhWCvKEzkjELPK80=
--pragma protect end_digest_block
--pragma protect data_block
nSHAL1exsY1pbbWjjgNj0EhJTGeOITCJ9dxIVDNV6XpQz/tXOzVwZyEYvtVhgSz8
6YXRn7W0BGs2vhQN0CYalT3ldGn3LWXyVIrsiV36pzG8X5yweiusmv2G7B5OlR3h
LKEPXXalBhhTJJy1F0X8X8YlKSJTLtZSnIUnf346C5fxCR+xT9Y4rAfS++H5vTtA
KNM540hOI6jmf5BpPpFU8dm3iJB6tktnVxbGohJdVTbOter8No8xkSLy84o0SwbZ
Fx1+XPKg0zMEWN+dAfnNYOyBtPy8OwospG3+kI5ufTwHF67qdh3bv9Xma6idCYOh
U653NJ0a7DhNvVyQHY9/uCPnvz2aSpTGLgWDXvw3ZCM7LSBSS7/adXFy6l3VxkYf
gDAdUVHTbYreqrxmkfttsEYsGLnRMLt3Y9RN0kCJADjbmow9tA1sfGQQLYjHhakh
cSBKFBY8329eS995+7P/Eg/YxQrzDOlPzeSpL38ux/0NKQdz5z08cF5lIcp67Tl1
byU9CJGmiF6gQsUWbpLc0nwXzW18V7oOlinl0T6vlA2GUegs+rxtx4oLxpLvDJgb
2RdE3nk8YvEW+Ct0mwC7QYm42tCAvIQSdF2NZRJtAWYq5cCuTBHza8alLsfYaYHu
OvffsLXdgHJ4P48aGccgOZ590A7u7XW4HYzRr+xPmxeRGyh9gPg9KX7cNB3Wm8qv
qxYGmluqAI3HHPu+Mcv9LPG5k9K9zjTiEjw42Yc0l8yH4smuAMntRrDKwBLXjV9D
3vnkBQkB9HlNzXToUuP0JTxL60sJktZr35eEhK+BNdhvBhCZhHCYi9cdGytgCPQ8
9ebOwND8ZnGphEx2v2ClXlvtdwK6rmYYMM2T5/BOlXdJamqRP89xpf1oiwqvkBe5
8DQt74Q44HFHq9Mj77kGXk2jvTCgM4Ck83KP9K+VZpu9p4BVayJ8gzuJzz1j0bga
A7eoGzz/dyDYlqXM4Ayxu4cW7vTkIbwEgHELZaoaI5qrVzpJsT0oQ7CyAZ7MnyB4
OXBivVc1rF2B6fbfpy7mMlIn5vEDRxjbXIDBX8MaTRJp2HhlBHz7KTN8/wVLpend
sTE/vHUQSA+FacPHqBDu0yyiAf7UwS+vpLtJ8f+yTM20xuj0F1UYfUv+2SMFIz/k
gv2QANHqEfUOm3PLncRvqffqY/CF37npUlVl1j38b2p+T5dH0yPHAWlqpggWaaZH
m/ExSK5Mqv1nYWDvKxu/kFUlLaOPTCZaLWDZkNmE+hqQ9d4aU2DEPAIFtRI/4C3X
Z2Z31/770aPteSYJ2DiTFrk5tfOBqtsUAmC7AQtHki+t46bptJGhQcCbTvQUmfNL
WYm/koEvED6DMv5aR4KMWbhKid+Ek7PCCVx/WKeOx+Mqn7dFURmlKP6/CwZaSXp7
cQKtOXb0nwmxJ5bD+iB+9sjlCxkiCsMHETq+OKzsxF5er/eVK01HCt9LJJqsCxiU
sGcB1KnRW1jOqiwSnDcOQK2pBAJaWz9hJ6miCJXp+GLs9iQ1x1emcs4SICXbSgYj
s7AYqwfCrD2bDraQoa2TD/c4DzLXrqWXlMDB0/tcapwgMsbI7Hv810BuIQhIwvYO
wFD6cIlhxrH2V3cFrPXtlau7VCokogz46OfKTAYl3ZLJ+5xGCoTOrIQM4Fhdti/1
93waDfI4R3YgGLvBJTFw9ef1BS+i2eVC8xeynNks9Ox6RuPthkwKCH4n6hMEaFqO
uoumvyg2ODIP2tjYgL6nRrH2T7/wf9F1iIuYwAoZXd+S80VLTNdds1JWbRtx6MzI
SacHIknecLAVRwY7/qnxkbsonH3xgPRQVvAIL0xbZ6gak7ZvsF9k5WfhMkm95cqa
BO0opZCEbmOR0zUSUhFZo7O2MeBScRb0yV/+ZuZdQjTnQ9vOmGHc+2jEEd7Yjyp2
9PhHbhMyIVMwGDSdiDIwQXjKXltVfRp3BuIQ6Leav+qjZniCrM5jQ0V0Uybs/5Nr
l+KXPPmlb6J7d7uVJWaW/tyZk1aqJVBMdUuu9EltD2kO4CfrNgSSqOvLVj+pttj9
RT7Yxgx+b0wGRyIPnJK0cSyInRxlFg6axYVWWuJ2cCkmyo0IFrQgNq3FCzsWqVaP
8mOFFT1yAqvGMq1JrZkKnifmOXOV+88ntaLgfyNoA8kewq8sDkhMb0bPuygpFcJb
DsusfO0N2Am/Lb7119xAVr+eJ0jzS88zArwJQpGZ3xXAkhK+eeYa5FtoNly9Hiqz
6/cnoUhG+Z88iBgEzu1rd5keYTnCe21y+WsMVtfNK4OEB1q2Fymng90zVM4Xy8nE
odgobe5/BS1YDk+96y+E+9GnAqLNTxfbPU4YsBci8x2vCGFYK5LUe+DfsIsXUyn0
wrliB6LGbi216PaFKXK9A/qJeYxJ/zyg/Q8XCZ5giWb6CjeVoISx9PvdwWlKVyXE
ST9qYdQ2lr0ip3MtKs+1KYN4yzjWWRpx+NilJr0sIyD44QurMpmfX+3P4b4+WR00
XM+/3LmkWpCzT2WO11xo4s7Keko+8knMJ7Cz4cX16NBe2hFALhNbR+vfEsmsABVr
Z0xdIvHFx1L5lGDeBt/QzmWGg/5HKaRWQTfnf2cL47jWfq1FllKYUhSq07kP+jul
qIGwCwxoAaHZQnwKE0WrOmWX3x8vRNN/RrOWZ5bzlO8ecAibPYGHf3f8NY8mIn1n
7x4afiTrAAN4z5eSu9INiaLzL0FYBK2PagtVf9SjLjyQhONuoscYK7YzPWgAWgGP
gYyzdlnFdqRhy6plnBjKpxeVerkpFH9Lm01Sa6rQb5/f9Kf7CmwqK8dse9KcMnzK
vtANWwp99G/qMU27y3W3hwx56nCH0KiN63UYpEVTTpNzoXMRd88oN07AQHy2GFqO
DnAsRIbJ40AXuGs9uTQLmbuzRAS1yssjtEYrgExMIF+25h48LamkN6XR3NimN5UX
Q0OpemJipMUA+pcIXkmFduuOu4YczPe8tDcH0vRe15Abtwisz3Uv7opi6MuxHI8f
KyUETfBG11rFNtxGtum1qLXpD9vrcKSz9lwbLebF4XViA4uRMrxrDA8c5RCpvRG/
d/WffdWFcJ4V3Kg1LmcAJ7LdqjlylX1pkykr9p7gXuCsADYrBaxClAvWJgZJWxTy
BXs0z4oyn4hXGC1gI51RqA2f+HqlOxgCY3xFsh+uCpyRLaz5dkxF0v2Kvzft85Bd
TM0BPOE+yfNdgF+99iZtAMtcE5L9gQYYblnMdwLvJpwV3e8QX1ZUBr3kE5EUA+x9
SR9SCW5HTsRWJgqydRwcWeHcHJb/qyoTOkrKirv+jXnQ9WOtAnV+InR8bfBbm+4h
ROImNzyIwhD+5x2+fPse44nNcAWepY6aCZy1uBdtHpXq2uJVDNK+laZRmFjJe8VO
uT8C5Hnh5racqfDpPktADVrNrbfiNiWqvSUyBIxJh8N8A412lgE+FO1qkTmT/liv
JNgFr6tQnyykXCtoRaXKr8jfEeOcOsHsXfoZU3Xc3Jy9RjipWx+8Vdn6NmuNdhO0
2HQaqFsfd6FWA3OeMyclo5xlG43So+axYSir/BXgJDd2cBDVK5ZHWiwPuDflrIjC
zQ9i4jMOGtrNJumv2fAxO3uCW295S+wJvcPxKnslMlu/kBY9/kGA3NgnjuMOk1pQ
aIsFZh39DI2Vz2kqhkKLPR9mL+IGbzE2GImMz79Ba8jhKWw0iFEVUc5TxmEx2WBm
wmAlpwM6DtFxAReuYo/v0m1U9QYCZd3OGG3oDzK71if48eF2jus/ejC025VV4i4r
vWKGmVqC3Opg0qrHXLlwPF6NOBsyuDnIVSyAYPbdUKQSf9iAT47zLCGZt8xBeGkg
aWezvaPjaRRq+2ybZh2MI9R+jIUGwrBe76FGZRBEAksxGGxHRHERQ6rBmmWrVjyN
U3BxNPRiF9olw2fhoilfydKlVn9TzPlGZBtywZp+VDRuqP2ePSHVK7BGDaplWIQB
pa3CjJxRKgXWraKoGkcpAQW0BlAQto4cp0+fzpbXrAquvZAkZDvzg+mbXOoS/V7P
rPyPI+s7PMxeagpAfV6dUWnfuukRDW9hNX/u0vBgJUFJNWRh6IPyR5nc87zKdXsM
UoXJ9r4B1+dqS6mCFY9OIAStmDYysxp3Eus02K4+/n6830FpJKVLwZD41vtail5g
QxB1HsJbrawdGAiV5vLrgnAl3jGw7/YsvX9c6mYMqt2ZjXPKPQQDP2NMRS+Lc9Lc
GGDqn9o0JPckeJmv4LSsxcg2xFtJphSFFOJhw/7gs0Uxd5otwb9pexB8d8Y2YOGe
kbLaPcL2dKK2gstj71YQkNvNDuw+4cAUIWY8TEKhWMO6+WbP8bW3ThlgNPbDDloO
MgblLEHzDMB5s4ni3Kinyp0nlMxNOIj5sn9HZRa90GlyH2nTpIItC4rCjcp8agI7
UG8B9dIsOK38YmgNh4Kgtj6rS5ygsp0YQ+cOG1hZzpvlNpd0y70Re8MWhKwosAnY
zXwDLL9gdvmgsC6YbQrc3PqCl92qF9S9QibcdcPytTbSFkyN0NElsCpLCinPA8Me
ZtyRgxHJHk8PCebgRnYDQcj3kgfKfpRrcznjgiKJxOVo/dPc8KIfRXdZG2O76hM5
1UmGKgNlMzpmUDv/b/h5dkOrYeG5086kpvx8u37Of3Ywp4a1L0VRuOcLDevBtJPM
i4Dt5swlk5n7N4Si2DRwz2wftK1rsKURo6xp8SOdYaTfnApRx5V7obd2aEhkWRwr
RLrDzum/08Emh3oq8K+9CnUAVESP2n1UVc2sCJE0woNt0ICx52Tgt0je1oPaMKlM
d8HLeYaVJSUhSNNiFV1QJ+3kBQkoSDGy2wCFST5JRMwfsu3iR0fY7oYLMzP3HP1S
nlIjCBUNud9IWltPIR4P4efG+P9a08kSDGxwPV9JujYtY58y2jUsXbYDtUpLZ/3s
e53IwW/vdHAYZwJ3h9AwgU8SAUOeYUdzt68z0vctp+16/BvHTOXNoBFGHcbGbN0W
upnQqcA3YpjiF/R8JJ2p/XtRKBEgJW43UfadDSbU98wwTiExZcvJRs4E+8OPOYCc
1Xq6+KvU4yAonbhuvQqpecVyT07c+y1Xr68GoelBAPoV/pDmWOujcibqopGRU6Sw
2kzWtth9aSYi9Pg4x13/s/jzz14G8zWhlROh+OOf374VRZZcArUJ9/YbW4RbOfxC
cHMpVLNOjBxQqHcYHye/2hYycynE2KLq2rQ3SqQ8vXlzo6IxUMegMLM6fDLcncl3
zMGi2FtBGXLbx43e9mVPsapbQ4Jakm9ZliQvOJXZUdWIt+ConkDEwGzd6Lal4x72
GB4pT1JgmuaDqreR9JxkORmwEbEC4Zr8Yn5YbH0uOQ+hjmY894nWAR8rWC4vchqm
I8b0TmLvZgv0BpMsWVYkCtIAOa3JMy0XNErQpso3jfESaojYO9n1bQTbrvelcceS
5ZuohKNpsZjAhgN4V2nX8LE09YLTKfAELuVhhtsvXUll/1VGRmy5tML9we1psGD7
oJq34wXdYu9jHb+idFEuIywLFJZIk6qTMary8trt8b592CPFSUY1x2mTVciEtRHN
B9vf5LgLkGKMmuqMUG5A4DdV/DbVga4pRWVDuLhbh0MUyP/ZRSS995ouh/NdNSGp
OAzMruMmFMfR8946IJiHo+RSPzdQYE4iTP0Z8cG/giL+ZVvn/3lmGOsn7dfB6Y3f
w2ylpPyEcMDq/sWc/gK71/9muXBeYqduEwGnMqOWB6NvEiZ1l4uHBubfxK/Pqk7t
2Bef/9wO1gsJCpX9QU4oaMv8h5js+6bZSx/3z+naA/bMNvOGCPoa+lyOr6v/ItuL
czOCw9KQ5TouxYqYJ4vFjqLTj9KheFaj1n95AFCgMNHZ3nbZ1w3WWEpljXSOa763
T7Wq7DxxtClSwnqjUtG9Ng3ZOO6tTgs+8hc4LC4vHP/NydAmF02bi9NG/lSNIXT9
bdNKhgdbhwzJgZz+yalEPXnHbYNIza/cZVfPd/wAbGzv7ariehHfBceCKlm+2xL9
/Q0q92pgdU70JxhD983jzJMYi3I7+QDC20dY2Po5rqlmLeabeRdQijLw9l0fkVuF
rgbd+aKaG1OI8xvpRjcdzuoIWrdsDsqNls4Fal4QhhRlppMM+RWAMtF2V1JTvMRn
td19DZYWJOoxBJWUXCyTJqRhK2ikZoyti7a2GmhtkVaNC3jgHDClleVTe5Iy6PZf
NEZ4WjokwDPZakTsrpvZyJBb4dH6fTBFhywLnsyEN0nQMrzDgXrLtE/QcURSQFhB
HKH1vO6pAsGtY2BgAND+PHnPzTKS96vAyplYMdu8UEjrE5LTmSZb8gxVQxH5rlP1
NhvDfQO8L1yrmPhnmWwNmk37O1RlfHFustR9RiVqZoG4R7+cEqg+liQm9SVQjNsC
RO7E31ZeG7wUmGgj7zbPiuju4AHO4kuaqmPPChQY2aeqmEfnTG6/xgIOly+nx4r6
56iJMFUngI2HO9aQe5oR2831nlL9IQ0DN8NJJArhmBmVo1EP+2qZJgUFEKoruUaX
MeWHNP8CA1auuEYolN6ccjMUWqpn7tNeW5CQCj5QoZFZsRNFC/lOtKY71fCp8imu
4e/+mhkpXRq9vxB5Mfe0ho2jVQUHxEXn2nOPTO3bRYvvnZHw2pOCkkV8KhsPSRzI
PPrMSjxeHuv3PoUkxDD9aA5XDyQ32Jf4BBKi+xUwLyarF5TS/mlaijyAiHgE4qMw
iSANLlpuRAiqAtsBgXngTizBHqt2F+uAaqd46YilpqNS3LReBKm01I3caiJYdM2D
PC5ocJ31YRhAxcZ88kpuzOSGng3W7/ySNumM2OCv5ISuIjfJCbnPZW9lTQ9ieUIE
VpdLpuZtQTYh36y5NmIdSFowjB3TGa4H/c9sc/jjyax4CnrsVFepJ5FFQl8PrRFL
Mh8OpJ9EOneBO1QF2Y0ApekbR2tlXyiZUM99HKGmKak5GpNSury29fzAcAfzx2q3
gAr+jxKYTmjY6LnH1y1vdAyBQ7e6A6FiOPPcmQCeUJUset90nG41PaR3QmZD//mk
O6f4uaFn4qz4fsarf6TnVUsn/Q8Of3KVnGGVZUrMP3auIrthn8HwEqr+me5Jy4fb
n4yCr/Ub/IZa4m//9fjMoXHMW1OlbOQsWN8ai3i2fl5i3pG/Y7Cw8iwKNA68Zo+5
W6T+sgijkATceDjN9VTttDKka0p48RReGtoMVlaMsDK6NPMNerA1KDt+GHdKsgks
3r4g12ybVffBu0Y7aOjVjMch941Oevgpi/xYLlQuxL3j9ORUWc5ilIf+Ee4wAiMV
XLKf0euOQnoCrU/eDmSQFTAlULTj37mj37ZPmvvqs0oPntmj/XXgkBBrp3iv1TRa
DkirY6OUOx9qgrKGVFP8SO1y2vKsZZWly9GMfYXEgGkqss1xTr5znoMOG1/txk6O
mMJ/+ZTpabCtJM930IZg5YYNd4pu1o446V/VkSK93uy2tjp1fYFf45uXl8cmOlBz
WTFVGrVl7vJoTpfPX/bfTVPve2tgxjobYT76/o5Xjp6QuTywDxDFDhH1Dn5MwEBx
hrH/JVkAk06ZAZjTdUE0+RE6LKCM1D84NxxxQYs2IrtD34qaAd9diIfdG13pnvoo
MFeupgBIHrOilezXez+kgHVpDiJ/MkgB7fVlooR68esfhFWxpsepzP1qhdjNU8Px
lAObGKRaFhRZASs0IS2epHJQ525RGIxKLbCwKlBbeagFBVZmJO1SbKViB1Lno3a0
Wb2BQCGFZQCW1s4YyM3FFTB5cCNpPRUlqVYA0N0nKe+snRcUtG9sKsjo9bOl/N9d
Hul+g+QFvIHRig5mTfJYtf2iMcZEHPFpbJC68OMfZ4R9/N3bMwLVvaXWju5Ly/HO
IPLSilQU/SiimJBWPRj5GW3QcxwT/Fet1G89viG+dlLqbV5l9fgM1x/TbL2LzlgO
eRc1WhMToyvg3++d7kRCxPDjeDhq8qWhEP0gFdACJtbPITaTA4kLfmIAB3kAIcm7
2+1fsjVhl6ecPJweUaoAd6IvWnA6M5Ib6KFriHxXAoz1ZBetf0v2eJ6p21LzhCcX
jLMgzj9cTwYhcDPAnrL+CJLbQ+OfvweOAzHXxj5d/5CgAfSflUwogmVwNGCD9Ong
vRp+m0pGuB5i12avtQKbsYPDuTEyxU0vWvVOra0qMN/tSJ+V3FCBjX6YMsdETKtn
xt9vLNw1/9ffPq+FysC1a2Usnwt5LRDfjvKfo2F4dRuJ/j0jmFvCKOSh0WlDQ+X3
lfaFLkh6Rzl0nL1xtJhpVb/nsTgx/MS8xu4VRFY6UqViv8+LX9WePmV8t4vx8Tgo
NuifPWAN0N6xOE56yc+uwuXrj+SfBzO1Qbfcs546LJBgoFAW1Euc/fp5LOkm/t+D
DVM820A5jmxNdGBOt3muWS0VJacZT+XcgC4Tp7EjQK37s101q47w96lAWLFmaYlT
UPwq6dtebqoHoQzF0OSvUq5DnjB/+adDXKBlO1XG2f5iFGvUNb7i/YQbAVr0v9ye
TpsA+RUUOn/5FEqazqdUPVzDnZVYlXISvwsDNZuespd81O/id3evm7A9hYwxxKWk
AfvbWvqNxk9APJoFrQONQre0Jh17NP4Uw1RamztflIKAVkiMbDXdVsEJiUVcnkHo
eBaqnnpMpdzE1ACX72gfv5gqxsvIoQyWp7ZE0Bo7eGnYbCX3Oe+Q4/S78lbRNvuY
jiskA4ZRfS7YOjpVv3o4HFETqYFZuiHOrutbul82Od1QXhD/oTS7/jgbwOQbJKxs
f/IWu7gOTM/tZLZIds+UQGlx/YkQD79iDgO8rAjtDbEqIKpsxUVyLgAoSHoFiDS1
C7HGnXtqbr5laI5Ku14S7r19UjMMlTwLcgNRfg/vB8x8R4dKdT1YJSNLU0UPWkSq
+CVrost9OlnA//CJKYgbB9cW14lGwf9+BF+UJUkT6O19E78w6MUJV3skwqnM5gA7
KAbujkTw43B+YiytNUDFRj76cDg2hdmw1l1yebUloIE0+Yej2khJAozwrsZx94gy
r43sPQIf2g6Yv7TEs7BvIT8BaDrmu9d0fOz8Mmm51QzZaqVztvZTqrAaJhX9DsG6
cTOsqINe+MYlndsGP0ljRjLxV1vz5JZQ4ZO2VOTPwgYxWuNg6c6ckf+N0lVLYVO8
CMvPoDEoalX5R9MzVnIrNT+SWQHY1QFD16LPpsGPXwFU8/fpj3DBVhamCisxCGFz
1cf1IthwE/G2uP1WZ/ai7XYY07MBBcXgmwp9Pi6TmgpGBsip+yGAi9X1PdLFd+qV
hFoTD8WXmEH9zYUuAd9pgpn7uszVAkJViGNj41JtyUjPN798Q3h4KWxy1RdyAb5u
PFAaBZUz5K+/wNhi184zhUxQiwaV9913pSivmkW8gy7QkqM5+gpcFCKgtGreegJ4
ufTvPF3TCd/wIVTWw54WtVZ8O/FD+hdMKn70EMP3biUCQrQFKOjQQoeMjIVYOWl4
JcHLfe1WlPdISEg+MWiNQdAWNijf2/Dfpld/yS7mnnJcjBi3tB/c1tIT1vSXAMdT
ZZPNuxc0bQRlVH3CQl2RG6hiLC9vhcEYDim196UTZLGlVcDhKpcWnqoovTsvogkH
zbAdbIk9edfbM5acfs5erqiuJBPHE84K7niC/Bx+JFRv+K88wzDqU9iMyXx2rZFB
KnqFOLoh9H2nh9C+8gmmcWHRBYSk2SPgvaGVAIgP2FkTeztD4ANbszsXhkkZ5Jdz
AUzWM9AFcjk7xs31gFm+ov4zNt+oegLP4yBX76Fw8yxXMRwWDOG/uuA9hKGEsBWJ
J12/QJ7xp86k0ibbsD+xjhMGURdo9Nk8m/UczpPd47BB3RF6G/A+VBtCCx2yPvOc
spMnghiLwrcUFVPeIfg/gz/ITxf0qb/lfmxb9VPSI3KQjloeXdP6UkICnysTVxPl
M21Lwed+RHIjHvW0US/mxj8njzpf4thYHiKHZWMnYsRSvokfokHOMHdO0uuvvW72
MI9Dy8VGn8xZ+uw0GLD43Dxc/T5QT6SIFJPdF1BgTEw1ffyBGKRlo4WIvJfJ3fXW
intbgDZ8ZnO7skrX3sz8MhDvmZRnNtGpM9gSeS1Ajlw9JQDWuSJ9R1Jxm9U2sE10
mfhakhZdfDCGQB5C1rsNLHPyW+aOhdlz81kAJzLqxa9bQLGzTxaJp3Z+EE9m2MTF
d1wK1knh+7NTNPO55oZP/pKq+oCH869GmkueXwBlJiUpyfJraoBvBuhmF3uaLJP6
UwcbMMiHfFD06bxx2LympD4yTksXjssAJcaakuAeTK3yBMQSTqBlLeLZP5WVN74c
VvXKCuG4IOuvEXUqZR/5Gv0bs9oA3maKxGyzYlnz789xo3bNTSuLMbVm83zCe5CS
tybPNXgeGiA39baaRVUkMJ4QhyT6ZtP4AhZnNM9vjGL2G5NaSH3KBDUdyegdyTzZ
ysPcbomgQ/D9bervo1wwqClxGYBEEIS72dyslnrSCLJxMH/Cj3/D9b4nCBnnKHet
9XdC9tKe2a2W9klgrgZUe4P4kxJkOUJZBbwDbxXRzomPW8Rln01DKTQXgOPBvLwQ
olVUMKNMx4f/1eLHflhYG8Xy7fp7J9IeyqnR8Lbgd/9yaZFqelCUWrVej91Ez3p3
+gnKTQr1h2/KKqiAK5woP6dmMJzdgfBsKjvnJGztGhW5LnM6q7Wi8mQu03uNBwKV
4+WR5Gn7qmMTcEsbKiitBlJ+t/qrsAWW0Ygp/rcC8VhzVL9r+yOPr+CIv0aO99Tm
yDbvc5QGIXwvk0ATjRco2Sir7AtmGbt38zrCUU4FFvtwW6ogEdyx6OG7bujLnUQ7
Y9+QMDS/VEv62LYJ0/8QL2nWskzMiY2usF3WrFH9rovrkrsp8JUDezNL245f8Tfg
BrdD5lGC7ZBLKeF2jJzf9UsGAv2iocbNJyjCfdcFgqtLtnepG4CFGVOhmVt4cyEh
kskutZf+A0eIT81RZYi4IUPj9UeObdvOjRcwLWrRb+4u0GT4MYtCNPSu1t+F7jeT
pRDACqTenMCkQ+U0Peuzl6/hAgMlN2OistUz8z10+BF1hOWbqsYcyfWbg9A0VCy7
BszO0FZ6tjLvfH0U16a1Da5dlaFPI8eRFDc1VIH5IZEPQ1j7q1pvlCy/9UJmFPZE
uIjW29BmtTXniKoooHFrXEtG+o864MBoaUx6FoPK+TZK3bKfmxEnT/20sFybSEfx
5efsTlZ3AWZO6CG5b+d02Hat85qEaBp5BeS10T0APnma7/Lrz2lGSCtABbEhtiL/
akn8CTkDGurHh4O97Fp30BQJuKQB6Y0HiETSt83o9tQN9sPK4PTIodgUWh6lISSs
01YYKpS1JcF2DWzUu8x+SblRGKfCctevxk8+h8oVT4yMxseZIlZJJ/zUG6Dc3TJj
IAPmkdRExJyPeExcckofc5Bw/WobmxMlY4LgMThzu+ipCGGa0eoXMQvAxCdMR5HE
7EIW/kyowH21VJxHW+VtRaABHMAh3tVaAh9qn566Jp0MNLEfZ4D5z0XynHuUWWVn
Md2znLrB2cCA3XDFi16NhTDyLGQaElpH1PrsYUVS5iJ4xMIV3evaFAjunrl+ncTF
onaCQpxc2uuBf0WhPMkAYzfcK3oIYIsMaBAA6oh1GWX3Ufiaa2laeatpEM24k4oQ
NlBGnQcQONAg8aOSPTqujrEDQhAjI9YUrHSq99vCEihbJG6qMz5OgSFXJtiqAG96
Om4Bl3WMGzkS/o6uFPiHZmG0TZaSEkiu9GPiQYZBqVPCiG3g1UdFsss2ngzrzQLf
GV8w8GXDwVtlyB8GDmefiHmTAqB8VW6IY6csudsiApg=
--pragma protect end_data_block
--pragma protect digest_block
yE0SXLbqDKzt0sCztJINPlyhUKQ=
--pragma protect end_digest_block
--pragma protect end_protected
