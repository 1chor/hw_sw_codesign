-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
AaLEccod7ooqb7/2sQg0m0vaMI6fTPdXcEJ2IPHEH0tNZJvOMAOc4j3KjB5uOiIW
qGLeW/s6MXH2QcZbwaAXkn0vHntTpUPw3TxfbVN8Y7G2KnuPnpe9QJO1DQO4SnE3
i8INP9kevEePISWrUWeDVevT3jQSpncYlihQV5FeCxA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7536)
`protect data_block
dVYKQp7qoENK8L7l5qPXVmk/VZy4VZri8j7VEB+xNIllfBnYzPArYROnn4GSZfSn
up4wYIMAJvWxYwCpkpPYTViV/Nm1TkRDuiM/77u+pQt5xUg/UnS8r97Omm2X/opb
4vM1kGlCEy4URwaQwsJ1/p8Q570wOIOLkZ/psQhcERgxHqkCTIEmHsFyK82f4QEY
IP8AGsdnlNoOd+55hAklWtmQZkq4DYCv08SRFiFpYOmJGt2z1X4PvjbPmUxbOs7g
I5kWax9Q8PQdanrSiqJtl+1Fw3y0ePMJf02jtRXt39wERAvgKt/0vY3Fs1wGJ3UQ
rGeuaD+ZEHUCkvfWEDmrjzyuN/JBM1UpedxwDa2nsdztFTwx9MhdxIbqm2LQRDLo
2QMgdp2U0UDPuF2+tHMnyteGsaFUYqk98lJrQ24WIDgwpV0LKCSKprLzc636Mxjw
9+nx7L5T832HXMSDL3UnS9S9PB+ti7ZaV0841QbeyhSZYinyVlPi6szCKk72yPTS
EEkOSK+FmLFZ2JBn+s0dANKuEwBWqn5lDRyLSfy/7UzSIoTt3U/Ny9I35fGGRres
Ak7/zkqkjTq9ByMhNFNllu/YCtf4x4P4MEbqEWDp/x1H4TO+mjOaNHCO0BPajkp3
JIdlKc+/4pj77/3usMXt/gHd+r1bNXGs8ULivLZBq9KjgWQdhUOgD7DblI2r5NLr
ezA/hUDeD3bsIpqXVB7X7h5BL1IQ+iwhuuItOblcuLdPw0+X9H0JjhoxoZbXQpBp
zhWmI7b9eZLqFADVHCSQGOz6I2nuD9inchmViXNHXgWg3wusGQJYxLxgeQMLpqyh
fvWb5jobeD9GLKeKyDjnflykvT3MZxcwnvPyIPcFvuYiN3pRKNYvwSjEdAwKW/uC
5o+xn+LJ18ex+sTz0secGPgLtHBdFKNMluSs4ci01zc7P+jyehtjXPM1x/tYVwrI
x19D321D/tiPlrohv95rWDU+u19hUHS2e/ufkTKfIKnH8h1PGS5Umwf/egPkYle+
9aLMRIzo6OgMcq8B8Uapn23UPNt38I4xmVwgpEemoSc5O5t0Mj4yJvRncEP16ObT
KiT024khf4xSG/i4kP9pJZ12y+QVBksn+wZVe6Rz0MSHy/u59YKfv3T8OfwwXsP6
u6xKN/6iW1D22w36LLctckZVIdEgjbv7deqgWQU663rZJ3cmonij0vZyHIyLIR27
ToIz3Qxi6rD1/XU51krKmlEfKNQUCMFb417Rvg1HvJzwiv2CxrEwfXMqLGE9jH9v
mZilPWwynkfToVORmP9IZUGB8s94t9WunZb7UF6cS+UzjvpUQ8V4URM4R9TKzeFZ
uaYdt1WPQit+GPGFjTYMpFe1aLtbpsBmybBUeYTvtgny6jj/lUb6egUeFZjnJXTL
9KRou/jgCV/FK1uLvpiazD6wXJdDX3+N5YQ03lGVR/ycejYzq7aK3jjzgOWosyvv
CBOs1ZUHWawxwW6k42mUeCLeZ/1TG2DnoQciBxlv1/mHEVFEg+TBTF72A3Vugpdq
07grgnHLp6NhpRWagoAvWbORpPt+Bjx9bvHP4zyh4l16pswcKAZQPgMY9I5iI37J
g27LvV9piCvuLVwN/dhXChV1ib4tpU+51e2tLfHaD9YJ9HeA4fxU4BmFbAnIlsRX
V2gzsDV9eD7NC8uWYl55R+OBYbR60mFRp6xHwfkp4YYzrXKbdOvPwTD6gJCAD56t
UCORm7ebgiO/9w+F4hIoWoo3CBXQOW0dAtVZSmQGAVnZG1/JYcoZ6zOUlZRInujV
ADJMnmQXPJDvhgkvKSNCp0vplLPCzetsVDDgLfEpHNQZvp8NEfPnFxhr7nMIG9TT
UFBUPwU3tOtW2AQ4s/jt/bESAGgn4U3J25HjObM8FIqDdsKVi8msJBPJ6lZjXE8J
Svb7qUjA02PdGY4BUhIyWtMeXudVSeqf899mvuH9kXymXrrqVM8EciJ/72Sfeis8
bi/DYBqm0KS4OLGKjbqNsu5wN7SRPHDewRNxW2QxLluUYbaEhTClpv+8xvPocNyQ
PA10Vh+AZ29J8UslBOJhJRB9vOl4cLLfgBmO/o1l6DdQFU9e2zDlCNMyHWvwfALP
o0Tqn+4IrWPXpyZkPKfQRiM5IbqKVv16/irF/Y1sp1Jy1pBYhY5yASBH+/XTQ3Md
hLaAd3bn+X2hWYAJlMNWE1EzU3jZh1Huev4x423apCWyXB6fMrbfzUWTrUEpjluT
vPMPYOI/WcBDEDg8W2ZGlgMC3qSmwhFnwG41SyL49u7G3RDHkOMtN1WYO58Zq3CH
eEtJ05VKKnkQnMD6giQNg7cR0+KEBbggGF0WTSYebD9FjdLBLWt6ECIqh5qj4Apv
AELve7gm8/sN70NzwPeTi36v9qgzGbKvlNgQHVfmdfzFFRxG1T6261CCmJ6LBQao
IPEiUfrQz+orMP2YVlGpR67d2ARlIrog7qICRLvjfvfGicvrIntGlu7wmkpmnCzX
k7rVLf1axpHkGJDdYRrw5GznMlz9iGvY/snSaIsmHsXty+hyP0ZNYlv6dYxWQsxS
bFW+wHUYe4NnpvVHIy6pFF+Q05jLwbquE82OGL0mKb44b1u2vMbfjZyApXdU4tCu
SBJjD28EgJduK63gM+8gLcqp/S701j5NM2wQ1RldQ/zmNdMlmGksYJDICIhtVJlB
utf2XHw+4UK8vq5jmpen6wW52xm+us1EhWXESbAzEvb0jAnuoSOm1SEHVV1BboHw
Pjw4sBRuDP5TIBjHpzhaBgmYnP+UNKEBY4i33jOuM8dqyt6TotLvL2tn0sn2pTIR
hWgc2c1szHPqriYUPZ48JZfeHOCCIZJNaB+L/JKOhkYEIr2eAZjDDQj6YRhc7Z7/
ND/7iGCSKS2Yb9wgnOP30/fsVshYsPJgJwy+RzKn8h26Tk+eLLrOQJtRejR71QEl
Zkx7lTY8VtbtD1tTCoURO0w04RKoyr3SkRBbS/SEWjzYtD/XzFgpgw0YXBoS7ZE7
zoRg1rC7GXMKxezH4aTX+Z+i9Qt7EcQ1INSNyqqsK5fAZ1M0+0qZb/FGyWX2qzwV
S0IDIY5wwRY5a8izMbrOAcqf3mEoiFEN7kAV94noWYVxojD0O69wL9NC4tU3pRn4
n+D1R2vPDnJmRrgxGi3yvY7AWwYTgvoYK70x3N4M7DbT6uvgCRgpk2tJzPRm877e
jKWNYSw9iuD6oSGJ1iYz6PTy4qia3GCDQdo/ABLXt2U8QO07RP7LQ0ZRzT7MEEM5
sqAUF0/7P2QLZEu8taFZm0bmxprd8FCe865c/LAF5CXE8Vo39T9txVXjNoPJIweJ
BT2PBFsxYogUWSrkRNKBdAESffjV1KHuBt6GWVMwBe685+LEcCFeK55hnX2PxJV8
+4/czBcYhBx8ReC0Y5HA0YOh6mFKqQzwo+PKalU44TOmiqNkkPtYAY5KOu1hyPm5
qPjGSs728raXdZ4XOSIAxCLbVApEtMQ5/kJ6Sni+oe9oLCUZUGmiDikiuel8A6yd
EeBqrAAe5NYfOaRomr7CNCjoeuyE+6ufYjyXx9nxSqZ5DVv8+o4l/4SwAAilL/KQ
MA+9t0oqbinDjZp63Ee9mqWZ47QQnIvOMUDOjSCrP0s8V2uiwIbVmVMCYbo0Gz5Y
heOYAx4/iJbNuHgFxz6783zFpuVGlaWQtunAP1wUE5M9yKgvlCZ1AZSm6JHeIJjY
4xmSL7z8phky8Xo51ZsoVIrWwFMYtyC1ReUXr6pgIUDZyfoMG+r/xRNO+mg+fvfe
LH678Hh68XOTX3RdPl040hi8wVfAhbqvmoKgMLkQXOqkE5i9Kxb0h/J4VQYZU6cs
ZLXlmOIoCC0LnOGtiSW0Ug5uxroggH7iy/aDxHco+wFlGAJ+cMfkBLmtQU50gniQ
wyL9fpPssC8RJCSAUQy0RcTlRL7rZ7A1dHuqbM+AyMAgSws0o34CkIcHEloyskuf
Bk5ddlqQYFhzV9S0RsQ2GI8E3vsP6l+MGt8UFD3cw1K7HbRB322nGhaU7BnOu39T
PQl7EXyYzsDZqBDbQ8ZJF3BXuabV53cttboTJlv9WbXOUNNlDrXcQlsQQgTqR3SZ
Ll2Lu1dh8CQiSH2zicDeeqrxy3MLkUQEgaEbtyopb4hXaGwF4v2hDUpEfvczYdYU
B2U+fAMiSJu9LADV1izm0IEM1aKzjoWsaGs6DFJPsubIR91UqCi4gQK8HEPWVDdA
UN6PNjcxKXDn2XIXJOO++bLt0CDXLy7+ngoufhDlHyKqvJZnPYNLwt9Y3/pkbv/P
FdUuHpCDHbQt2fdQTNcbj8FRG+KTHCMzN8rw9+bvnewr8xqBp50Ms7OJZISoEaAs
wLmp7gp2jyluQT+t/DVef47YtcIu/WXAiqcQoiLZavtwn7ixZRXQsEp6vFF9K6lB
yT72rE4w2mtoeG/3DZKNQMZoSxYBeb+LYnq+CsTvrJDCH3GwpM0yqeF/AwDwiFjE
P86fakTgmq3FnHBZ9j8gbbqYSPxDJkYuyMkkIPu/LMPeK+8tRDrqbky7bT+zTk/1
W+wuTbKgnRyiTeYEXG+LgzetPd0i7pafaVv58keO3mmsXWlhI3Kb/MLHFm/Pwnoy
Org7henfXHEkReUVUVqeZ5Ca/88uzfHh2Ot0y5jEEmh3YMh7WELS8pFKYysISTL2
oA6wwkxRFtoOscmj9ERvgCSLJw3MnQEcLzcgpZGsv7cOpCOVFpVWDJBPMxWEb5nf
P0kWT8+Fe1CWv63ZYszdSSf837djgeMKvNge58a0hSAICv6RP698ZojyKqConwmm
6lTDFMpr1cOXUvHDISb3ZkE/rjLpq02BxUm+6IFIvcdQJu1zxESg6u3I8SwKQdjw
llelmycE4B8if/8l+i9Ke0/IyDcuLNV42M/b3WniHcymIsnDTPpTAlSbZ59MTW/j
0u1WiTDB8UXRCIIpXLtDRO6tQ64T9Ae8Z3cd4JdGZLGaFRGU/ZPLfp6zXD1tV6Xp
CS9P2gJ+OGfxY+7nojEWR9WDLyh5oxziv2eBGivUhwatYPydBpyEQbBng72iDlK8
LoezCfHrnKSWB6SkXb/H/6lpsfjkk143TA1sePSZpmYDV9H+5VZbnZddDtdFRKJE
9TBZn6yDKMrjN1osDbuMHZDORJdTJmxRmTjQxHpyEfMo4NdzcllgJVbgwt8NXrlZ
sXo/O1JkaGDOtzV2afE6x8PYlU1iBkKmvTpNZDB9yanbp8VQcSRbLQwBSJ9KHozy
VMwaVsZUkj3r4A3MpfNlCjKxqVVuePDIIuNra88mrTpYhZdCWN/YQitBiDIfN26L
Td0p15s+aYYKzZcybkCcoTh4fGySAdMs/+0Y/LAR1G6kPUJ9FDkgLZUbeNvLkPnn
C4KcMbLjdqrrqsQvOkkny04MUaaYGpdPkyrM9d/cAkNUaFFDOl6S1cCP1E54Op2d
hRmOlUH1fD6BETe+nRQfXsAy2jYe5CIZfe/XcfaopaXB3qr7V/Z5RgSPWrO3fGhS
RzDjXpCLxsgx4NiYQ0Ky692hfI1l+gC3TL+4f3REain/X9KxcTh6WwWgDTGjoWlz
RXZiuCtjhTF3S2gh0/XK5fvtlWtOLUBkZgDmS7iOLszxRHfs5CFNlscAwTEsoIc2
+qhom6QqIQLxJ+Lfk84JRPZxd4CRnTsY2+FLN7vNZDnpsydmydEpemxvRgwHgou1
v0c8W6uLBDpHFCx/99w6UsqFD9OJZgqgxzG5qO5SrJrBSA3el0ok2lnzOZGwQGGC
hC1OFZ2WmjtAx7hctu6OmtRpdxHmQEE2k1phz20WjLYimGJdcDe+qXKoyMtzEq5Q
+8EEmMpletoDhLY6l7R6OCT7bxl9HtsyZROkR1HVUI8A2Ob12XlFaB0ydV3UaCcI
a8f4Y87oOqjo94npJPT548PaY4Cqd8/4JoiQkdhdp44eulGwmQyWyGhcphJhU842
DUneSpsqK7HIh6OYEaYUI8fwy1NEXOhm8SB2tflFSl2un7e7sFqJXB3KbkMis3x/
VoKGbXmAOmABfN6YtWM45WIEuZQ1yGZkAca7RxOUXmcBM3DZti9/4RKEAYnnHj1b
udwrFbNfoC3JUMk3Qlz2GWBOfVMiudIZ54mF+8vV/k/gWALRQ2dTST1sEUQTYow9
y9AfLwz4u/IICPpfzaklffUOlNJJ5bjadrQCBuQ/n0LU2hnNjuQ/wXnRhy7+Bees
uPkBgsOlXFLks8PXYMA1VbnnO0jatLHrBKRq6g56kUK/s0+y8IFRUCdAGHUQHy7c
Zy7PwM3zQWOeuWyW3gjLNbEov0uLC5Mk2YwN/fQ/bW0pICbaRuIpg+vp2LLbSoxu
fATZThbd9TtLjCnIPYowEaq01Dhab9qg1Wn/Ym0pIqVnd+nCLHSQbqiylGvF9H/4
5GjH04zSwhlqfF+slcaKRswMbxbkX+UQVPMxMf0bPIowvQQE1YkNoUi3WhtSgk74
2tkJFYm7uvJOXDEtaMDArEv5d1Nu+i2x+VR4OFOq5hhmM23gR/tEsZlPAsjT7WDb
rKraZbhNpjJn7XLyz2bwu24QBrGmvg3y/amO9AbDKJE41TzVuSMsFbD5IqfEKX2e
McKjDPLO8evYdtjlMc4S7tcW/jp99gIh2fLXQDoeVC9SoR9f8fjSuuJAO39pDlWt
vUh3XT47wgpR5lbZDGITq0heD7z9wfV2Dj+f2cAdbk8YU2Bt87+OC9+pZYBzSA1R
JKxtlXaA33nv2pkktdVVy0TvPGXSB3jKM672AdKQgTsoSq3mZglBTTGMU+mEZ5ZN
IPRF/uwaI0sr8ZxyPI2qi1zdfWdtzTymGdjS+3p/Kp/yoAkNYnouxlP3t0NY4IhS
WH2ePT9HIQPh/++9YbtQ6nFSanFvAW6QhqEIcaq4vPwpsbao6tKEsmwm+PHdgUY6
+nBW0eedm/W2CRoFv2glbPfGb6JUOs0zUZ2FZsYmepOYSQW86sEqnatVwHmAYm7t
mm7iTFSOpD6bes3eUVsA1wjhOp+Bq+Bk3UAEDy3zgfhh9jGsOp+6YEzR7XAXpHqD
TlRGSKuX36Q0NaOMjut2RdeixZPGtDO3jvasNuVfgRYCe3hCe6yEUSm7/VJdDYKA
lYBNiSXgi4ruusddjSM2rO/pSHitYk5mmzKRc4phPyXGv3MRpawtXW8/fIs50BuN
UCXa0UGxhWLLdgAdPrITTy0qzN3TOToSf+wwIa0oPxtZdhekfgcR/Hc+7aVxvs7S
rhhsD6IH3Zi3rFJ14oPnImMNd5IDFz8VEVzT0gI83Rx0SvwQJpDbkbxBdj0Gcu4y
6fBfDJAYOIgIo10AzYuVrtDf6sXHxM+7dJ6PQybHbBL7g2dMDvpUK2FqRaLoOtHJ
AC1IlqeSqkL+EQqBc3Xjs+WpGqmS3dG1Yr8HBvQbwJj04U81ZN324pwVaT9ZOO1I
FqOi/BJdnd+IUF4AhlpVasziZ5DP6G4x49pw/3hFffh0F4/fBnW/9uJl/01VcTMw
tR196swqq0WWyjGU63pcRHNn3Ca0eQsQ0CfFkKH6Zn+e8Fw5kdbs3WhChls0Dsfx
qRPMl3uVb9LkNCiVc8FwcFrAsMJAnQ28LKUo7RG75O8E3ctH6ICd4RdENqMcSJqb
X4iOFqQ8BhbbhOpLRQejB+h9SaB6Jqg3oF/GYMUFaVWvNCsTV4kATLVVVvLceLL2
BrJPlKfNJsD/SuAu7F8TitfBTfvur2rrJU4uAZA47zVZMZYcT+KSfiYw0zJCqv1X
ogyiJ8rbz/JEoYYztUAGI8faCz04m140/qdij30AS4uTazSy+AbRT6BH/1VNyXlB
y/930AmA6+5CV+B6ckD+8VFsukg2FGsnX6dDfzYP/WYTTFGir7lxDlyDZK0b0844
lvmA0V+FAMm/2RB+NaA/h02CpR0UPzTRs2CtZi73ul/RHvBWWqk/P9Iin9cClLPa
GazviugQYmvUlq7YqBvM+aaCdpMCEZAzJSdPgrCgWkWwA/4w3jw88AW1HZApWr7o
d7tbkeLtOnw/tDCZsUhjKNrVfoz3vD31kZhaEa6hlGmN+iu1+4r3gQhQeWNGI6/w
ennBtX6wWWebwxj+SPdoJ5cLfyGN3gsApl/ei9zpnTCx2at9u30ihWijWmKvVjNW
IBO3qnOX/pN85nYbW+txTxlyxSgT245hRRBspLkoMH2YsN8pHyX658dlKRlkJCCU
p4QUIOD1z4nX2mjcKfbip9kuUYF1vsB0PS8G8LX93yDQ7q+mYPWC938GiqPYc2dQ
oBKP2L0lMmSb5JQ7RZVPqdCrQ90TfEgP+COzAusQl/3ECnCpojI9pfl5J6BTHnTT
QMa2ch+O5Gqmn0N6mGjziZs2lTWlqXCgRZiCXMoUNcwmxJLx+8AIuaQ+VcrBEiS2
qOk9PLhoh+NupXKNuRh1eoOYKUKFnhB5+QiGT6W4ut+LMxKyCQdmIcRU4Nbl5A8F
iH4a2wDdUkPjMg3jgafYj7jl5+oOoD54ug99S/c2Bul3JEtH6eCfXUWAp9ix6lGi
YogvOnQVFG7M32LKdg0FFkueOufcQgoqS/WxMFuJ8teSRm+jp9JJM1GaYUWJmDvn
T3flNF7Yp3d6peIvmoZNRum1GPCnt/K+3f0cwtKtc/x8OTZioTmNmiNvLv0dysqn
CKGxsohNMxt3HVo3NjxRFuWlZM1wXDAMNNiyJ8i8UoP4s1gMiWncHBH59aIWuey1
tEGbyUbaIpV/PrPTI6yurNcGBo0KEyRIeqFpns5i6KB0ipevnxEQXfcfhZ5UHmq7
g6kX5q+O/bMPYnb1VOHJxSIv3jm4qbDBnKOUzVlHF0YKBqcE9JqQQHiG/qK0bLJU
788dZ7My+Wi1GUbIXnuRjsMjOytzDGnxZ2tqIXjkq79x5w43ee8OrIbX+SYRWExR
DCCcdD5YlT7GEHdjFrpT2eufyDb+8+7k/mpCO6pVxr595gueDl4Iy3rpSX3T3Qm7
4y88CL1IJBv0fh+WUxDff1uKm56cuPzSQrH6LuKIhKbbChCeq+9cWBfmHMx4tUwR
wD2LPF1nzBmKCme8QTpZSJEKfz1q/Skdjib7jcfVRAiOtiPcMvI7ThBkwEL2Vz3G
vmIszPtFIfjSP31zVwn/nV3FHEMsB+dqfz6odTsWLdibOKbnayqNdVTAgggsCAak
ONMWLvcKI4yZ7XK13YFHtMIQISUTQZZR/DQv8R8hNIxGhaK55pG+93vSouPoYjIR
xDX/Y8/UWc5YHCfY7wwhPAOiqUTGxFtBNj1yx+/ytY9QnzUiMJXxVEE4xQ0Nuuza
9JUhlylx6N9i8ZIcfYnamPJRFPdrWnQ8pcjjPtd7q0JblrP77A43q5sgj1eijBJ3
UDa8nlLEiG0j/FnrK/Nx/TLmIl/r2kw7tiN0HtEAY2RNthaUDi1/7IqIVKuYEE8c
W8qGSNdzml3aJ7rVXDjOAzzKHGqBGRAkky5iLktmVPpFYjCz85Od3pWrWAtKB2BF
TGg7v4KnPM1HcbwVTwrQuWyy86sHT8bVXpIpBISaMP6jFnI2uG+Y7QGoKHZvCi7Z
SZOtVm9P6i2N3MJT8WIJ7DOs14Xh4qawmfb93F2SVwOobwsmEwS35PG9PrGyzXsq
nKZTkMTxtBigvs94hnt7EgiIYn0bnFoERYIjRd5P6cnFt6J6yrRDnfH05ht9Ob6P
N11IoUa8szIoO9mzSIutf0v4I87PWdkLqDXTcXxhtBwYRgM2C0fKWDzIoMAxs4kD
vzI6RAWF8oGceuIM4DrdgQJKq8xiewU/6MddalVqhL3NV1sk83y3od4V5xKskCs/
kk5fL7Nd1PVR5xSYYF5hYfeHvMOZoEI4eNJF8UN5Yb/lLeupItOscvO1b4lyV6DV
vu737lYHu9zpq7tCXgi1HWg2JXKBt9XvUF/y0RApr60pk2CfIwL2Kfv/U0xWSm0h
hOYWxlYuBogFr0a2ic1KFj7Kcg9dUV+ZUB1BJI/656FcdhtTpqopmVwHUP6OEmyi
hu1/ThJguNEPKG/l9ZBJpvx8HK90Auelb41dMPmK3oyOY2tVjJKXvCbfPdFgx/Vt
`protect end_protected
