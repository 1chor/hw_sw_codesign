-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fQZyjUBIfTAhFVmfQAmsyfvyp3Hj10/YwIeFYWKee5huyR8XW6RJp/PWODDBNVT/oGvXmaTEQDfr
f/N1w5NYHzrDAB0WSry5CI/AiST6FkxbKkqhmdEtBQoDmDrDNRBfI/kGPZsSqMznsD4SDtZJ+scm
95IZz8GNtFbhldKSiNQluI/MxdX+gEdUgrlvAPyh+B7i43z6NkAtsXSWCnxW4evnLkilydnOhgK8
9CnTxJhoVYpifuJlLgr2qoW8bTZOE3ww3IPetqOyaQKY475qOTN7r8xxcU8OL/jbqIvzMijFEpPz
SbshgSEs5udhxULJGiI5N32SNZ5Vaxha9czRwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20256)
`protect data_block
HhjSj9O8Z8/t8jk6N2MWlm8NGlFGLajsRTroRLlUTYuLzCs2Y+3N7KO5eE3qvwrO6V5GSiQOmyy8
qBcO+uKL5aGFa2leDll223zNxXlBfodoMFocNxMgbmbiFnT25nfDS79hZH+5rD3tEJ/g41e4Y2ub
cWTssrVJdY/lJw8KOp7pT1oAZcxxK85vkhAU3YqohR5Pd9I2SX0rb0bQg6BursxPiNwqvPrDyqHR
/1Q3Cl+te3NtWt/AAGgSDO9tTvKy5SRwYDMrR47EwmfulcJeMp+EYpCptXf21RdXVt3bFZH8vqJk
45j+2Y+k1amwfUpEKcpeWZBXhQc3FgAiVzOmP52jSYZNEPQbgvu6UCD143kxzsoXyF2mViE1da8D
an1IHn1l/hddVhCeEoRV0nNx/LktUVo9tyPYfsWFHx6Ls67NAe9wtOXBWFb3i6oSb5HOcyO+W7v8
/7fmTF/aQmE2hzi5P9Tbjvqblsr1ANvJtLEdEIQqjOVEOTsawMcSaqqyz/15lQCutGl36Jaxm0f0
5v/R7huVSDyYcN0id7jpIrLKL6/AeFkjDrYNuacfoFIVeRYywQqGlDzFkbC2x20X6LWxlom1UePy
z6Q/e8GGkW5Xl/ejIuvhIGlj+CtTY1j9yUfvEciWIvRc8F8Mv0DQoFOi8PQ9pzx2Y+DFB+PqYY48
9uThEablNTXBVZQolHslaDGOGVdlmiVi7l8iimYugWiK/LZic6Us6H21is/FqMnKcTVApZ5Wp8jc
GFUKM4iF+VA47kw0n5STEPmV3kmvGY0sa8wvcSvjmuwQZmAyT/8i/Vlc3PjbCTMjo1ejhejIW4zJ
SmKU8+xYl9HtyRGgd8tO+fF7mDwog8dODe1QMRz7jdcu0W2hoUOoxfYAk+EAnZ6DjzUwUug1AICX
JxeoxlI4bBtSaHYkGo5TSFeQCE6PYIMPIgHYYeXH2t1GdpfU9Cfhf3t2XhtNqaTvujioov4Qjlo/
A28xWVRw1lE5ATy87i9/pBYNu8vjlCoC6LwPjssirmlfN50ss3218el8Z0CBVnzBG86bZv9iDyTB
R8szAm2Cy3HZKSITrHyPRjE0LMUa49hef7vdGAaHvajpSmzAURpaA0LLMMk8nJzrj6r1mgmhT//2
lQFfz3ebpcdgI3dvEtWx87J2cqL0RsD6Y0UNDAUw7jsbxXDOJzjtIin6o2DC8HPl3GjZwx6ICoTC
H79POJPym+pec/a4RGW3FvIQQo49ar61XG+E3omESEs+QZu33y8eF18CTLC/5cJ3J/FcsoGJ2NV8
Z1JdujdI/abHB16NksXyPo35HlkZlMaZU7aPJfgS3caQj7W79MqeVvh74pkz7NMUsWb7XqaIkj60
0glD+AHvxil7ggCX7FZO/paifDp4kekvbigG4tlr1swSeJ/lyU6sERfO25zhRAeJ5/YcO9F+sooo
6NTs8LsKhFmK782qsWkPCKhyQp3zaIEaBb06rb0364TfMoGX2LT59FqewHq2u4PPFFs1v8kWyqZg
xMOQUYkDhbvtGccp0ac0bmrs47Dzj0P3iBMhsArjdsoSsBJdYcu56xGW5DshES4DNguwLdcnAX0+
kGz0pYii+X822vnOH9Uzz/eymDnyaI1OaGxEly1f/2JTTGU7mPCNXmzQfIR8EJOGdob0tXINJHfi
TgW8TQnpajk7909XQpTtjK5oZb88EqzPLi//3rXlYlZmV0tq7/JaoUJsvbxRiXxq0Yc6bI8NvsBg
e3kBo/jh+jZVRdzJ+c+/c6Yr8sYWZpvxa2LZZlOQMcWh3MIih/h6rbLsNAtiJO3DXycDmt2CQTvh
gd4BeIniyuQcQk7dClWqK41sWOVWk0oCAO5SgzrjKHE3xP1oUYxK4KekalEDL8IkvoTFMMshVEWx
/KDVC5/3bWCCVskRlXDetWjBjCrn0ulhX1JAkOO1MwNU3XhPSxk9GATOvkeFm1+y1HdS+LDG6Jvc
ZIi79BhxDwPrWOBjaLXg8U6E2J5ykUjuVHWuHEbtri93F7uv+rU8CyJsK+Ru1wAB8CtZpux8UQMG
PKXwRd5uhwQP4aXiNCaWmCdaB/5e+/v+7atzY338s7T5m+M8aPam8KQvVSxTmqjOP+5uEgzqvP5q
kIcq9nCZtjtTCdneUhZ0kiBYd54HSuxCnssN2VmFiIlu3L4ydEoP1fgQMqoN4AevjIoCKT/8lZNO
zKil5ndkOu5IKskHJ2l2P5FeBWDW1vojW4lVJtUy4OYqLoK7V7oJ/yK5Q6bRht/znEFaPWD0hlhJ
qMw09+AdX70rYEpeGrIH4p0iintX6uh8I4egEUX+j5HiHT8t2Du8oRGYnPyTiuOjbCRrMYdaw3tS
JLzHlQ0quJ8InWa5Tc+OsC0JdG+oGok05h/g1ye+ngOYFdKs8KZoRYXmHHl1Vjn2HP8p5yve/Tzv
IDWKgE55aaOInJUf+QOYmC77lxxYudOYHAtfF1nq6WW7/uqvGaaFZbhpe/1T+fzJ6m7zA+FrKagp
QE9YEZnTV1HDpENCPK1ut2n8zF0t+0EPKqoXx8eKzBEg4buxX7V3AnoWvHUpcd+GtWpXL/7HpX84
NI3d0hEG+ESG5d4dWlBlRpy6uLI4j2SJ/uQbqsuvGZY46wOjiie1imT1CuE8JtfhVEBLoHmdIuga
1X3V/viXqoAtXsE6YfJtmc2QQaHkUBUdyqAqvfGnQ23N+I/mRq1400hrRSsPYC7Gz8k4atqE780j
EqwkNjxOg2eFRMQQQmRoDO5XEtVd9aB/WTxO0sgu0+qBJKatEzH4Gg9HaYTlrPbt2MnHyUByR1Ux
UaiMsIw4LqzTQxAdI0iXIwDYt/BHFBgmY3bNkER43FymtZ2G/pEHE6SNHLgt1TYoixcuCiDNciWF
MxLuc+oCt5X1NbHMgTYpnbpjA84U8e4uyubHd/LAI4a9dxqjqKYrMaldfQrbZu9rJ8lVIIPRGlZK
aidjePMKBuOErx63G2PwxemGqj5ys/Nzk5zANc+gKSvUMhWw7pRFkrTHaKFxD3jjnuwZlBvJo3Ym
CSX9B7gUtEl24jlq35lTYapPQeESwJ4/WfA+WBHmOML81tG+7Az1pWsju3L5/ba7k8zSwhGcpgQb
BG0a7Jc+YTBBl/Tx4R9Q9270p0aqsIEiRE9dh48VsCiVO2GvhQjx74H/lpZ2IfUAX/ejPQwn9Nk4
+mmwKwxD+iURd/3DmblYVU3kNntxe8f3KOizZOW/FuoX2jlxhbdOY5cbco2JiP0NRIBat+hr988a
K78Yn7faAysYfwpY6S3MYlSi5oJHJb0jUS26O3sF13R0vVZfT+WbK0vyu79oNexp3ixG+YBbgV5+
FSVEadP4nI9ymDMXLls3lPJ7s9RkI4z2NZC0czkjLw3oPh1Pl+fo/aG3V5aWqBuzpPipumsN2h37
wwOHvQGu0ENhtO0nwUHzZEqlJHOZI9qOIfVbqQRG8MHxLEG+sWwajsk/K6GvgmtlgrlCXPEfUB+R
DCFBzxq+DpGPnMw1V5NqJnmJlDdSFV5MRWoaOH+Eu8s40H3VDW4vqKMowLtWZeFPWUn+7lInCooh
EX08lQ/cmpSSJYW+WCiuKXRS64wZ/+GSgprlwg//V8kEhwY9FFN2nHSaSiOeVaDtzkOX3kSq/Lxi
V7wFNXNgPCUD4Y5rDS1Le9Zl+4pt3dA10Gthfol6Y7b49LppG1iMwk9rx1aEMpUCPeWXmz1+dnRv
ZwRMdPjC89JYHQWrO8e0a/SwbBHKE2wYy6SeDXZEgH8mh66Um+6B+qUlQaOEFzOn6ZPSSGh+Ptnr
hVMcdly7ecD96m3NbAQxyGzZRIh8Qsj1tQ34WyAw914zOfUhjRZgN6IQUSUMHOLa7u1bSvLd2h2m
vKFcI8NbkZf16LPn4/6/9Nt8v74qb3NOMQ2ams9N3wWiouXJ7jhbhIJbmgMEqDQXWMreHw2Xfwit
b8RunbryTDJ//v2R4j0ecaqjnxFBNDtleril68Niw49aHYq/ZosRAMFAoJXQGhiQ5/vvhG+mwSBX
jJzgtbgEvKAvyO1xJhZGZSEJWYGGxeE3lAVzzUs8AVzVjbRsGq6P4oAq6FRe7c4TgOqKMEeA68GX
azKTfXvE7T3DkiG6UXZXroguRcfa1+Xinj828KbbbfrhuuPyIOiwP9Kiw4TVk3DeURmSHiwR7KC4
/2oc7xbnS+1uhshQhwzp0o5uAIYr3WWUm3LB5f/FMB+iAxmCJFW1EIXR+Ld3ZLlM3WIh+LruX5zK
Dms5pOStMuAzuwFxoRbeQmfJPEknBQLAlsYN3X9mrn3PhMREJHaRH064PU6j+KcuKARUypm22H1n
XEMk25S9+YlPh2A/5U7cFl5xlFljL6PLhfVReoRk8UX2/HnzqpfmGflZ0icUrqnDnlzmUYt52yM9
ZnHJPPM4BPv8aAAAhEXtGAq9NjSUz2j8scJPzFGOvlof+HuurNk5+eRVQ0T71R5HMm6NHnNpOktd
jIYInhhFSVgF1RQMWtNfjFgtT65Gfiw6kEbzymXKzUuo+y+VNrfNhS+O9P2Oav4XKBq60yLuP9Dp
UmdGM+T4gs5w/06Po5sgbMpRaBnsSYZB5yAGzdffOmxIwvVXBaoMcnPG/XHeOZexM53R9hmBI/MT
dp+db6b6fpH89dmO/9m7SzpuOrn2/bAJV49ljTEfXt9qHl2OoXLiuAxDVi9SYoBF140ibVRJVl3e
H4D7vx04YJnFoqAn+eKCc7kE+lLHMbJHFl0Quil4aFu7MozlGZXuwNAGTaPo5/j3ypU3cBvJ0V74
URln198ovBVi+AalUhCa81dxxP47AGxYN5LUfvpBKFMM34wxZXttfJdeUSf0iZCsOZCatFLNFsgZ
P+nO7QKIJ5wn5RDJHxrp8/Uvsw8dvuTMAq6lXuzYFZKhfRjh4cpmsFAKM1BsONUmtEPyrlFcIi10
9PKCX3u1upN3MyEEbXCTUVYRSF29zb04uzdpaYu1MS7VrRAvWfODqgemBX9kgTX6k2BmDksssEOe
M17cB0gULL5TUBiFkGbsyELV2FJ+2LMAWLCZ1pLole8ydBVRJqsCFuATQBxwGU5r/PGSbgt3CSjt
wDeelWpTaOSwEa85VJEkwHSJglJ6dzALzsB3OU8qg5BkrNa1sa5sT13BShHZpQNWRMJe3Z5Mzhie
ySiedX+GuGpigKdZ4OOtEd7HSZDfBkv8Crmo1MG8YAuuWpptk9l8f+MgDIaU4DbZ5A+TKBdmNIoT
qod6gHc6F7mO8kgi9IdrsLwGVe1pnXR73zr9zktSGz6bA79IuTW6/5OP+Y8s2zCSe/b3/J56gb6N
Ersc2BurzJZTbaChmDBTXb1rpGwtPfJivD7pWoBTVKLL1vIVMAP0kWfy62qGvWsx6vIUxOTj05bO
g7SQGHetG9cK1CMf6ybw3O4oY/8gVAYv/Hu+wanMfclHtrCRVf2r3WFs2zDaJnU03Y7/TTl6pGS3
WPVDTH21bSmn1JUu+kUmXM7RA1cFh8wyDvT6etUDbqHMO+daQrLKDhsaUw4HBdRyDgU13c/bG5Ho
B3MkwN4PrVmmuGNbHwyOPAzwlE78l+C1hnXOMjyoWfT/Lxm/FO2hY2yPg9oeMe0piajUGAqTXcHc
NSXHOIFLB62JoJTL2hDmagINFf/XScpE//ZX4FSjhOXJXtKHfts4zd6cTGSC3vbOw9FnUBosKAUn
fCQrzgMeOd1Wm3XIHVN5XuGypZlpvuGAtUYk3IhhID4YXLRhqwrwTk89bIO6rnP6RuGn4LkJEvj4
AIx6jmcIKvg7hB1oeGRRi6MguRXOAM1xq/l63qnz5iF0m9zGPhYgEV/RJLsZUEOVbYKvQTdmfBmf
R12AVJm7tQLB8RJuO4n7uyes03wRHBAcFA0g6ZsPL2kkB2576zXmpC2D1tiiqQ56O1C/7ja1Ii7k
U1WMJN6zJC9IE4x1YXUfxgSfTcXbFlWQzJkFNXiNYczAVmn+CfTcQxb/QRKUKKkM0YJuZtMmAc8i
ccg3YY9Dm5F2rTRWXg0q+px6ugA0Wa6PimWPjV1Q0zENYB76imVrAoEG1K669mKl3IA/f9OVRCba
xeRHOKhVCTjc5aLMpfBmoRBC5imSwWs9nLtGhNu55o5SLh4nXJ0MuTRAJiH3vMuj84D87s2QcUrD
VGHNmCdvRW0wWUREEp2QBnPnQBFXhGRdzp/Hlbly91qSNFoXQ/FsKeOUJIGxvDFvhhJyq7zx6WmO
hN/yBqkrqflgzDcGLBVVbN/mG6ur9wma8hafAJr9qM/JFFpBb8W7C3X4/dm+Who4EcYXxlYBq3RU
qxeBAu7jDQu0LSCfntlxZhqbNS7sOSgTjtj+gTomr5vyurvqtSBlGH3mSDzBxhhOuPd1/d+lgeZz
IHU6cg8pwKPOlCqwFVKN3CS6oQIEKCeNaPFmvPZmDjSXRK+Zr/kQDmA33QQ7gQ2gj87kc5tdf4wK
NBNucFGcdwpZiOZWz21HE6aOe0V2K/mRXeoiQSvObLk9UBVJRhCOP1YxNPZwlU8tCsYRexm6b60P
eaHaLW4AJfHt4LUh7cSfn7tzV4uNFFQY7EWECE3Dr6UF2UQCklQ2uWe7Di//qHQkEaP3zymZ0Bea
FiOE4/P7r6PRcyLnNBW7qkkJOMORsJ1NV04u8tZ8rGOUJJmrflr7dibIkJ7WHSEcLBwPQIlz8DR4
81Evv41WRRqWzOhJcuEWPUD81E/2RV/kj51V1pCfYMASEmk9H5SCCVn67pthK3WUHtojgptydZgh
MXX6nhRfzCalW8Ba8AaRjLmJt0NoykhwPpyEs7Bq1L0jSAq/R2tcfAZFvnXEeWtFTd3/tgnuoDZG
Wy/LlRvo2CITo90kpnAAAs9Tz1FhQD580ClwSBwlSZWBPBBqee57ZjaKmpc64pvPe2o/1MlEL0Xs
k2UdlVSJQa2pabQJAJbpYXI6VGxlTg5toVsqzZHvqk04exLS9gWZ5zrVipBbKCGS0XQGH0xskfVC
NJI/3hMueU0ie1Q12ZG3BK/qrWeeu/JepGZXyjf25XpxHIQ0ZsPWcz3Vdtn9Cqw8ukMG8CFWYVQG
J2cDw41RY3oiRBBstLzG4jn3KpNxBckAjVbG2fuk5NVy0b/AjnFW3t3UC5zVTbQpUhRCO8NZBLfk
lBieq5VoIVr2j/F5P42MWMIxgCZgzJox32f98JraK7pu8EhOPac6kj2DN64CHgDnMjYfcQw92nZ8
jglGq33yt1yvl22izwU0CbV1c0QtKVmiL43lqIFWf07QXzT3f3zqxhyagpWckJXa8LjM+qScHIEx
EUYnMeKZKrUNpeTb47NqjZnEmS/RDrIHiUDnxJaFHwP8PqkpU5lui1pX29nng00FxwWuDeNJAdrf
gayLAA+exrYsH+GzK1QQyhN7zQOfpSKPYu+OQ+9wRpOXn6oYTmjLrbuAw6CSTxDRI4o5o8vCIqOO
Op0GzwjTrJ4nKl25L+WOphIAXpqD3HB5wN8Uu4aYy1Em99i8eC7Wrs2CHylfoZjTjIp0IBUEKxYc
g+cPh871sC6BHOzWzF3mciqNie+LamruO3fnwjWpcOFwsB/kmtUyksdYii7ls8rremvPWcWcUTkP
hx0SvCCrguDe3S1UMNRlaHgKeH2zvYAhCwMKDwgc0J9RtTt1WmJXzNh214qNR7vTC+eOH6lTDrOk
HXx2JXxxXKsH2iwnu8xUo7S0rRV4o6DwflwCzauJmCenxs/apEas+iCVcvYQDte2YLCC1Wa1OQa6
6+pBDaoWyYaiMdeCOvorohIOhHlSrICPfYtI6bYGPFZDWdHgEzKkSVbmILt0utLP8+jdOqGLeCeg
1CmE5yhmP6XDnMcKoGCKFw5tyxzjf1oCRK3Zl0g3ceP4oTcOcHm5xaArsRcQVW8Osos48kagpXIp
jKP9qIfyEReKmnMBgp5UnSJRAPz9YWJ0fOZaSBM2eAnc26ORV2TL6zrBzJEH2G5GzagfMboPoeJh
la245v3mU7S8En55fDTtfw0JgoNxao5ui+EjmD9ZC4MNK/CeLmyrhMuCas8+Am1R3eJEII0LDZWK
ObcBTRFyb74vD6ZYOOsSPpVWorBSSpPaX+Nkf4m1pe0rKZwJqe1ZsrOiQAYtGvxf+HSBXu7RUUJ0
aGCS7camrkCnzzACDwzS2pS1Ecwt0sOoSRPxfZkjoD4o5sXSeU8BUZg3de1hFZrstOnIryBJJWC+
WDY0eQYYgfOwHKQqNC5umj8T1tlGaSBUY16dXqONwUAnJ0bnwsqfgO3QjCIUI0NxsGzgo1Rubglq
ez74XDUcU1Ea0j2YC2ByqEqC1xqKhGw0orFXh7h9Attspf8+e/hTG9k2rSn0qi8gDem0k3Tz3YDm
IHAnqgiLJjxMnAmxOlKDblNKZWcs3cQW6BrL9tG8QxSY04CDjOGTAV8aw+9yj4Cknm33WdU6WHMm
92MiX1hAZTJuTwRpMlmqwTWQO98oT1/Xd1cMa0FptXKPkGNrDqJ41hKTsyyU6TZmrpN5kD8wu5Ru
aDUyWatNd9fUNqOI4MUSfEiQeyxaJHGj5+0KfQ16Ahbj/IyGGIyt+CsRPPgD+dXR39Qtp4r3AOsI
jxIo3lNM250Sj6X4yrpancexYyYuP+wYXRlrYXm18A/iIL4QqbfV6drBJkxIgPMPoEIjVu2XPW3N
j5jcJce4WGlSmp1XGuzqhJybc5Vy+21SVCHiwhoGcShWr/ZOGxv1G4hW0UzRhawK8jULBhe48j8n
06nucizoxx3EkAY9f/ALRvatN6t81Dp0Pj1bSodq91hlaQPymHCad1Z2vi5rWZjWCW6vlN0B5BjZ
STphLSX0AFA0HxqiehZOtfDW9WespCdew0/q0c3btjfCzal7pIaIjhk/bzoPU18PelGekP9kTWhN
SsiZzGsUqdV6M3alEGWoNJEWNC8Rc/cAWpfOtp3cxCNdufurbpiyfuLa1imnAgkM4EHt11MoDILD
51zzP2mqalRfYb0xABRSKWOBUX4mvjI4LhYC30d6imcEX+Qbabk5S7EiHKIOrYLxp7O60GMTeXH6
ILt5sagW0Fxg3PY2pPXVFrZqzHOEhUqvB2xBOU8hdS2ipgwBH4uAfto12T69JVLw9sVqcXXio/FK
t31n/y4hCD5FyA88UqZcVKWsCst9K4+P1yHO7VXVmbeF3kbYaVF2HK55pQ7T4dRsbkf1HqNjcnT9
MEQnpa7bk+hylZezMLOW9G5svneOCn7TqInPucT7ztBFdpjY1Lv6Z+EF82okFjO+7BV6HJS/Tcnj
gOSzGTrRecK6zvXYyhmUfXp2kv3i5UxbuQ2psbcljE1CV0bdT8/YyVINPgp2w8eSuabsT5xOvYYc
KiKFxMoFVddpFUGTdRx2Jv6RYhl5yHxMNbP73N2ScQ2AhU3H14HgN8jONI/WH0mZjXav/ccgAIfn
pkY5gRHcivSnBCjdw4CzY05m5KGS+uQhM5Gx/HQwDiovHAbrBc3buGcafT6UkXRYiK3v+6yMiTft
VRX3ZKYZ2Tv9RWyEwzXQqzVcuewlqZA7qJxSv0Lkg6eXRKRXbmCbwIy6OSYx/2jh4F15hH45Da81
CjEBQFqM8zu8Om1AtDvQnX4RClgLyIQAZI4IFstmkmQZ5LXxGn2FWyEmmpFifU1O3WMMy2Hz3QEh
Hxb4g6E1Tdzgz4b3uTCXMxqnBf+XF4x/poRoUDo8Cy2HL/V47c3Y3nXKnEaUwhA3Gx5aT5NEOVF3
EM6e+VT8vhSSUyCF6kbJ/KCqybwvzboYrVQiuDpMn1FZLdVuAYjEPcqYX1jn8M9ITAQs16UGxaLk
mAq5mWiOC+asz5+YGC2rCtQnsHf79bWeqqZEMPlp4ygvFOlWztHIp2e2K0KrXoFPwKFd6IjbZhig
L2x9rCV+tZMzooFKPmP6Xek6aDWwdsJ9FYJSuvX5IH00Heai14rLJMQrC+MbdXpg/KMjUmizkukE
0lKrbXZACl7NTZLIOehQEj/GsputmGOaAbCwgixIxG+yUDCo10JkG3oR58DIVmZkvEt1Jdcq3oKw
wi0X5p7rZOlLsvqzLpK2FVcCCyerjCAMP34SRZGzg6EXCPVnsIx+OIVx/R8CHBzSOtw1GWAibXgo
iMKRwZHIpyH8TujMLx4mZuuwRNwzNzJOcytutnNLed3kHjMnfSZAv68tC3yaC3S/KTY/q2b4d5T1
LJL0Is6cucKxQCPptyNZ2oUTyUjtkaKo1QvR9ugeQncwkk7Xy/q2VidTGG3tLB4FWEFBeOw4kZph
oSQ2NhYXmhGMOAfUKmWx/n6SU89A8kGc25fz092jFf15i4ht17fuqVXmtSvLteyWmFeBDJJIHBx8
RulmWNOwCO0c1lFmaSKmBORTVHeBPyHidVnJsB7ul2lbEYB2Mgd8yddlAFoapCn7JrZOjktQ9Aec
sbJSEPeRp3PDv5aIU2kZynUHyoGp1qJIUZvOlXqQrAkato7nPAsSJ6fy8OhCgO99uPBAgI/E6DEq
o2VpmFSY0/1kGyXsqG3TxT+274OpwQ1W2AcmiP99uWvNe8ZgkloYPE1HJa0qQR10Vac4hcjn06NW
3zSSiDKU6Osh781gNMuZk+Atwb3+L3yrH18CHnabnqHfk0CeBiJX1944k4AUDLoC5VgESq0UFxBX
394nyTAWTm19m/0j4KpJIugrsosRSenmChQLoNjWt6m4E3ofWKW1znU4IN4bYTRSegKDB/1lDL4e
9PbtJPJRflXo5WHiqtnASeF/5K+qESiOHRZf8WXnNrjunzX8M/45/mwISj3/fx1poBKif0ubjEPc
uNj13sgt2JkUQ/UvVJsjW5sio2+WGGSUUu5iYwPrafSdN9FHEwGTZvRBvac0c5j97gMSb2qlJoat
h6+PDlMz+7qjWFhLgrvLhOhYPaDjvn/oRRadcpDIRCMlQa6IqRAjp8Aru6WlrrUoA8OeotI1y5K2
7mr7CQ5fT1x8cxvr0RTglcGYny+JyZJ6c7ltARieYllnHZjL7ORUeAROX2AtIVlwoeplkzR7cHiw
SPVpdGdgXqGY+nLcxb7ekZFLzwyfBVHYxKY56F2MZrBSNwTFxOhbIWi+lLmIvsPdCAyXwtX8+Dsv
q7qLFtxICw14NlKmqHZ3HUY1ygqvufSq03rdDkgId/602iTMpKMBj23Xpp6HQI+A35HzAjVcRfzZ
aX+ERZJuxsSA82wAKsY2jvS0ftfW+RT8fRHMJMvctGsIyTgbC6pBXDdx2Zx7dcvybSru7oDBaIta
T8F4erpi4XqTuHx5nDHdxuvWjm11ebCB2AnrcFheCUzuLYSNwhbTxc8WSA/8B9ZE7dvIikdnHVwL
Qafeoracn423/Mtt1uuRSrIZeeX7eFDtmBTIVzHWFjkEJABMYJWz0pIvwO/CWbnQtA95h+C0E7zW
zYm5lfzTA1J2fE2qR6fmSMHi/N0S9+/MtOTaLcQq9mlyG2TeYtH5q4rkL8lf46j8n7hxO4tBBbiA
Nyz8fLkjg7amdQHoBbDZuP/Iw3+0kQASfD0ZH3Gup/Jxq999VzMvTRMdtKjzz8LBAS4QGATBAP7C
cK/Zjqtv6IXhGJYD4QfEVeKfSkCIIFq/sV98XptMh+7SqDihpTFKjnCY5T4LpvoT0MOmGXeHey5E
PhpxN8Pe8rJEQkZYgIE/KYVvnOHJlD2pw4D6dHm36y/66jV2gMAvO//ULHUSPWBfu2uqHOoOEa4C
IboNLZ5XOaVP1BLtFLGVTaI2uAA3UyFtczlkMKFKlTXJ+sbTLD6i0AzOSKCjbBvH9QhdPouxC+7n
REiANvyiEuA5ZqPsdEXSyipQ1AMP0/FywBLoKsW60XpY4CFobbQH0Ow6JiwbXh6gWIk/0Mf7PxmV
80GhxFHjNj5zpET49xi1h/SijxsH59/J0ymu+ekAKxUIyQ0HKeMgO0fMSS7E+DL0bnMDE7g2fuMm
/M7RcXuE3kMPaxJyr2O/R8IzBQJUylceoOkdDyVPdumYRIwqKuVHJ3kYzBAwY07mpwTDBT9zj/ZJ
frOXGly1ZLqCz4G/ssZEZwlP3V7Duj0QxA/U+ty0tJJ5yQZk6F/BdwJUiVUPcgzOxa8XOk/hOmkP
chWM2YIbjXDCPhqhdLmFyC0jRUXcX3jhl8XhvW+Jsnp1oFoHXdCY6gBJ6Cjounpj562D4xTzidRO
ABXnCjlbIVK5SmVjN58zrrXBZBuVewgG6nI4TEKHppJFbyFRsR7CUGPwJfyp/ZolEobc2FAhBoUR
v0OPUeBSYSDMlgErcLrdgMHyScuVurXQ8ydlxLscVTknNBXddEBX0F8ETcxQQYkh5W/m/iZ11YxK
EMqTjHBz7qtGT20rUvLGqIrcuqENfkVEvrhdAP9t1SKLAc+Zx1iVZrnWw1cgWbR9QJypi9D/X0zc
H5h1g3COC9xE9atMrxa1ost9sCvL1wJEd44IGQJ6MwuDCw3QNPEP1h5jM4lUMjFoseSsw1mdQv+p
0DEJ2jalLwUhaNODyZct25tCmf1RJ0LrtenPdDEgf1qEhCg81YYANLZqnFBkbaZISIc7hoUXvjMc
b6pbmJO2PXZlQpbFsKI8aC45Lp9s8lzXtnfteWOPdPPNwwanyHD3G9s/Nyal49mIOeDavkweVXEu
qOHjgKMXQIoS5+zOgMSdO1mTt0bIB6NKD/ZoNo3Nt7nF7u3L/5v7o3yBc5UnSjmUrd4weOAPQJqG
9rlwSttEBw6yw1TCMJzFzyKl01TpsZ6HSbhruniDySm30bfC2sGo3zsCzssC/eqLjeuDtoa2i3S7
sBvCeRcMc3JdahAmuQn7tucv4TIk+bpAHhVFBKWgjaxZmAeVS1JRFN19u0+s4hC8ETCnu9+LDki6
uMPKQVcMMEh4B1VGcFX8sXCL7wSQXigWdstcBnSXhEG+J0MCrRXyvCehUep/NLaMJB+/QZ7Ds1lI
ZfJbR0jobuxH0bUyXq6Y6WedbcuV3sw5h2w0q1bBjDlXEleCEorna+Rb/QaPPt68hzGQdOOVUSuP
NGJVwyZAfeQWDXzrCNCem2lowQ/BTDtMxCgXiBDpUynE+EGYDJgBqRQUQ6zhd/+qhLaN1cqwe/V3
Pnjb2t9pIci4PbHOjDHmtKZvJRE8kbUsjY75+r68yYfMY8TjyJk7u8C/FMFlg4WDOcjII+focsIC
mylywHTjelg44FT4JsZQgD2He0c5stxvcePYjiSY+zNV2RoEQk/WBT75Tqk9tARK50lsVxhVlTuW
0YCisxhoiWF1SjmAhSFeBKTruitsIILGNI3I3tYVXdvvvqJMAlCfwDUe1keeStm3X8XC8VaEmsdH
7AwgmvWCTGTkZ/E9TkihqeH6Zn03/b5jPH5uB3eK9vH7qFgfZ7pA+V3EmjooAXG1qulbJxYMex3G
3VEkq7eUFGCwJ72VvUmEwdjnYLTLndJ5/AUpt++UPggP865a7b3Tk2oQvQ+ajbOKluDDYnX6owli
XXKczk7ptUMVRpasDeExNOWj1Uk3NgvzJuH/qfJ/LEgW7y4FeVl8IMOqL0OAIVYYopBd5WBpPCre
G0LjnxBHt0mQjXcSuFfktbQgn5I5G4fRCjdIrjqmUACuPIuBMSa+pVJNbP9Ysu0meUzfS0KnI1r0
3ixdY+a5m071ljHeda0j4UcAn+OAwP1soZ3QQ+i06S3TXsq/jjfr6rVJVHuzHkKkPqrB0XlYArQx
IG3drf6nC5F2HtYZoA4aNTUOVwPNTLBCQULKH8mgZ3uduUyo7Gr3i6UJYqFypWNZy8baPlFil5ox
LtyYOrypIOravDpRvvzV8sHXir8SLT3y4bLhRYiWzfdcEpAVQLNcjr0qZ5T+vd0166S8FfwQD2Lz
RJXq8dnXI+ZfwXTvHUC/CUUY+D1KFFzPE8qyOV5AoNw31wIv12Gx7kge/+OEkP5tsGFXXkLBXddT
wFl9kb2qVWKu3QoaQqfspp+8JGfD7ry3C8YNSlUFcRsg8/NcOgWstc+WDPkZWiKLK46kwMpLCl8H
5DDZRsleiR2zGlxLV/I49X416otmhdaRUZCkEAMWeJOhdYtHwcX3xznNQglcsxKPPyBB5iR2goEq
/DRmLM+GQEu2oap7j+Mx8gOwCMDCVz+c1EDSK45n0EPRAnSfJpPjo0DtLJbjF4vLnafk01irVd6n
qScZOpp3g3K+HnUeEzga7bT8mASXy1pIiAE5n3P5kr1PxBNoJi4bFDeKW26+nX26vtVpZXKoz+kh
KZ++FSMUrFxb9IipPGSgYaCzWp56AAlSiGTTJRYeD1BK680i0g48AOXY8lbo5zlKJgllDQvOHovV
tedGkbq0BWwav1xkOK/tpdyLarqiezqgvRtAj5W5qMApxcwWJagThhtZoneBIooIfi/Veurchruv
XYNNg7nX6Lwd8Mja0djqKe8+IZNhsrCuQHIwLo2gpGG67wwpyHN5z2ZjPs6W7/Omwbc6o7m3LKPd
+ZluardNHz+jXK3wN1j4sbG6Tp9EfCVap196lKGqeHKfQuF6i/pPFYSf3h0p05DBP5NFsu/PCovf
Wtc+ddWU73l/TlikKyWCJdznh2aspL0NwSyHR+HENWFR4FTIrIRSMxEWAL3b6SZhrIQkHsFgvBHT
K3oPqNU5I30eaPqcapcM6q+IaWh2nCTl/mOiSsBNEA50aabiKf/06w4aaPStSq8G/IhPy29s9pZF
KIKt+kYz4AXAQNqBocKGeB3oiH/MYxTlKbaiqXcVOPQwVqvLNWxte5yZVm4VOJ97bLJgC3pCyka5
rmSz/nwETadhLjTFhM8jXZrUpJwUdGRVcCbLhYhZ3mtH7pvU1dyMQv/+HlYUrTYTaeEngZdIYxkU
wuCJyPoYtFueMhjQ/vudmLHDP2Gyz+06buhKcN5ki+FKAbsIxP7n9+Xfxe126UikhPDGkEwiJpI+
qyfIZa7e3L7gLbUPQFRiLZr+w2Ksg5bsTVX49UUwa+xBD66Ja7sfxbPD9kaXshH257H4ifNPmXsv
8p9yEGypKOUwrrK3q89cM2KlDZ7a/ROuxVSirUas8NDifpxRE3pU2z/QzJm+1j6ETWXdOhSsJSSJ
d47Oug6sSo7lHJKWfW1MexCcCE7m6hastlmSi5+VZ0hp5OmM5o1MiqwyKjcWylEJE8pQxAeTwmlc
hXWYNPLCJ0EpYITPsbbOeVpkXsIfKS8ovsibEy2BUCrFS3Dh7b6BnSwM88spqi0uThHKah7pjQe8
pKqozSvgAaTAOl82exnirgtX6O+wv1HJu8K4z4JznWI0gUO8QeQc7bRZQyRqQRBd8pne7Uaat3VD
EQ7BUblg0WWYZ5zdupMdla4Dr7mj0hJU6wnlO34KMzhTZWPboitsqjWQi+OwSfA1KShrxCxMnFw5
ZRDpQtTCOTBAH76TM+TGdKwf8llXIyXSLsfxE3w+ompQYPi1CqvU7wa2+ZEEFDXYcprm+s29txwX
hw/awe3GiuclXrkWSslrIeVXY6wc+jTUa/WcyWmpA+/JYHh6hBnnWWCegE7iC/Ao7G+GB9pXFKyP
bFDwM1XGCgxYq4a0t9cQFbQXkHeYqMeC6GpQRsGeTvyi0NpUQPeVKqlzs3w6fXuwXk16yvY3Zuaq
tkQ9nbbUMDMh6LTXg3xqt2OwJDjRD4mAtHyegdbP+vGtVis8/9JzT6rTSvYf9D3Ud1cJVEe2AaqV
jLPupGIJPz3nOkAw/QNkHO87MuUWD9fhSqHucsWHhqlJ852/zbS/9seUY5ZK3fkv/ZYaV0JuVsqK
cAKsKg5na092I0v7l7EHgFc6zltp+wVVGFSSLlBPKJvPA3guFWf5fRb5RaVqeJxSdEDDpxGmi0l4
B0cMYKxp72eF/4V48E7iBdx6jiG9CZ5ZwMyoYCc8kbllvonR0e3Mb4HjHWK1CLU1TZejig7WefKy
fMgthrcg6ZoJfPbgHSe+ZiSmShxwZRbY+BNiotv9OXZWg0SEVpgdxp2SA0SV5GHQhIJ2k0xrr+AT
Rru29APK5jRVFURQg7hnL8GeAtll1luhiKMIHxTUgqnkRu/k9HxJEWdajDZrgOCEyWEzb+n/eoXk
OX5Wd3dEHM8M5wXAgFs4IRgX5vNiO50eVXeZqbLD3HI3KhpvOIW0ex+nyrppR7B6WF5YGc+XsbMd
khoBdZ3xW67LRhnPQ+GR2XL8+Y8TLlZ2DxP1ZwShuOlLi8XcNanYDARRE+qAYJ2RfmECBwpTEe+1
OHCKMHjShhtC/b0yUF2cLscfLjasyQq12xRFcHqWoibj36LwKPOmRxOTkMKKPXu0yzxCrcplND43
78d0C5PTQXCPHP34ERKIAYF94000j+aiKwf01Am4wBR3Oodl5p3siMwfFtIGP9Y1GokGdpn/WKLY
QrVqxvReVJ2LppC4eKtRClEpcg1J5s9etxtK+vvGC6il3N2hZLmlaJugIgZ9XShOMgjw4+un+WiV
CCb1xmYcqnntouKh17TRbtwRzvplNVTlE58a7EVnK4wV0OZElZdu2dZGg9Um37l92v886NtyoVmF
ZG47IMZ1OW2PHsaWx8BtVjCkXjB5iZDRhDko3W4/6oayxWCqMvHDMCMxRtQh1nnhshvALCphzRBi
GuqkdwY8HAA1CMmy38an/+Y2Jq+owgJOOwcXtHfgNNcEUpYwvuQTdpi7A7mtLw/hpzf7Eu/n6/49
ZUNQhoR/GPtg/plFG6Z3sJeOHiLxhaYZG6Kg/7o1O0k5uNuZ2fv8aEltZokvqmqKXHvy3fyqbybr
IZRcjTfn3Z21UGzL2HUiAKUJVDTjEFifJjvipxcy11sQy9MDKjROtF9gfctEwuwReBdYybUl1kif
Ak36h76w2JcDlIpDI0sYCTZHI3WIZv7JMpph//k8GilH2gj04RNL22nMmUdRAJ9lvYGk8TLgC2xA
Ys8FkJSYH78+FG8vYLscBp3u6REgBEqkctQURbBUabq7DU3NRQ811U/EqLIwglr21CCABXmjPU3c
rmqt74ccEuCnF6ThmxPLXBLKNjGChszwUZ/H9iq7I+6pSPnZr6cIZpDn6pC0UcghIvEAhxpoAizi
W/+tVEunB2VeK7k5yDGMfZJ1yJJBMA5iA16jtcplkjr1bZwzBFkCLyfhygHSGtDYTcQD/lr+kgdM
AN5PyiLcfYKnXSn6VzBr715JgdTDa/YSbl2Ns/ZV0IwoB1TgSdVnIk4mEiXhR8QMklfUg8s59bg5
wCsCOMD0X2xzp0dz36Xl0P/ad8vB2Xu1Y7Ax+xq1C7jtuvCJVOXpmRnDltvDSx9jGkFTNXMNQM1C
GzeARJSw6Upye581NbUIFQNfNZgyGELHYDqG45RPo8FXkCLQKT59qLZsOmKD46uk3aeJ5XsbYnnY
/wWD+4EEOwCoVGmXlvTI+WXYN1Y8Mn6a45H8sTDxmc1noMWeB3kl5ffuRApkHUT9iGMt1UJuNnno
Xwn8S2rQ2FDt+WGOvqHTfCd/dKEOjoXOFiny7akCpdF12CNH/L6m6R7B9MeY80vvzIbehO7S4Cyg
qt6hN82AOfsm0HUvHtywj5dzQb8NTUWRdCt+iWJy1+KgNC3OkoLnLW0dYCnmcJiagDi58npFXrkN
5FLAtIYpa3DL7dBgaAUB85nKQVk8G1GHy7OlHm9k7r+1RNvbmoQfqlPWxj4mErOX4pp9xylgx+Fy
QYYP2KXSRCr4YJ+GdV5IyqYxPAePT264vX+kzE4GZ/YWQaLpV6nVC6wWfMm4FAp3d6qq8bl0tHM3
RWunMDN98unFpQOG7O14M0Gqwe7H1AUK8uRyU4jqyuZoT/gslEFMCsysmYQImXs9EQlgoUVbWeJH
S7MMRPnd+U2VRdVjQne18ZJVMiYXfIEDdP2qh72Mt9wEv55JZiSx5SbG27q2lHOMbYR4Qbi9nNJ9
8HfmLfmrACHkrKTBOt9kYAvYMrDjYf4e8uFcAAcqceTdHF6MRXga1aMACLhSYQfN3aJoLMUmXtjo
228i15ScBTsXuwBqLTPst/NjSjA3fUJChmsdEJdrgb6YTtb4UboJfGuKfz+yTNv3zpHX5ZUiySRD
VFKBygoKstYKjPPjvZuWLcwDlh2l7ReM3SyniQ9ETvEHgDH2j2Y5FwSFD3t5Ostl8+6jZul6qNgg
dIwykAlxJxO2pbx9TTo+hkD9N3JfIAJHTeqdn0xp5u3OR1NxDyICCdNfQ99KI/UDFGyFE83bHce6
EDdBes6r2I8mRvK+doFF8iAK+EIlbqBtEbhkFe9c4IXPM6Z/jWYEa/05B7c1MHXuuruUe0mZxfzs
f+MrvHd1yriNHC1TQZKzajkYWzUKDKwvYkgsICTxlFjvMOulJBbI1PZv5FTw3zpJHzf7PNA25lbp
jIQrjrJiX6pHhsTczSODLflW3Ujt3dfgPB1dantaFPhwraG612lYwiVFPYkr/+u+fqj6iuCSfJOk
D/ikfdzCcUhiDZOlzLyUEBC2vgRH1piTiHuKbt9Ug4Z/mozP745sAXZCk1UF9fOk14ibEYqdEVOE
BjXqKanJwi/YEkH722IYFTLBlC5SRorLAUsWO1enknXoywIXrq0E2muZWFAq3ElVyh3m5qnxQ/If
YRWPfDJysh74Fk+6vQHXD4Rmg81lsD5DU8kHdDx9IBvYx3IdPmbVweXILMNBzNOFPLG5beuwhJOZ
zqae0LIu6d0CTwTr/ddeCtCsFUi0bpGANnRff9UUiDtgrLB1ewNYwFW7+XiYXWo2yNGr+hhPxhKS
hIZeED38epAO55/mdTW68zAsgYbdCq0QnEuwDRsGNFosh/dNZFFJRwL5qBrGYNm+9FyafjVoxEUw
JC2eI/aUZA+7+UFOyBNysVfEZRPEbnOd9xH5BgWEykVUhEQ3HTn910+a3kTqtCIi/hIXE+XiONB/
pqzV/TZLSKRnNPPilv42niI4Mnhy/HTcjuyE2594aDNzxZQ/z0XwjmALSfsikhscITy5Hr5ziRsg
5FWES1e3LhW39+/rqWaqAEwMVLNIxXQytEcVMKO01RJOiV1YD0udZredGSrRKyb3N3RNJ9PzJk0e
R067vbXdeYM05J99dSaKlp/bNBIVplXMM+iGT3X4r+Cx6+wC+SX/CpJQzit40mX+/WLBW1UUu4r3
CngPHmmWHsNfe4Wx9z53N6u7L9Sf1ptM495yJvGdXuajCOiOWM0MP/6f187I0wRHoPvRuf/v0+TB
BDVWWAwaLBoGBwTuc1UQArxVB742fLIsrzyOrfcu8aTSeMswpxGJn7Jx/A4Mpg8Gxw+wWeAH+qaA
BUkOFOX5TBuvhw99NID+G88Ey2Q/tDPdVfwPLFDe5AJMErGC7b897EusotEcZzi0qv7aNH8sQNmC
pVustmWjKiI2Lt3N93uv37PIWH5y2H4HY86GgQwnvQ3Dz4MfcmlzYpS7L6utMj2kh4jgDOpf+71r
0CuxiqsXIvlz5AvJLs9KqrT4dNGuH+HQCETBfJXYaGD7vjrjL52Q915swCziG6SoLHrOqxTlBIox
bTXV29sdUiS18cFlCYpGMxnQZlN9MbUl5FMzqkrdRePda5PKfoKJHwGCFsrM/Cyp5k4gtRQfg8sk
+AU85s5oXaS1NRtN+lpnc9zPteriDAA/xscDPyObnF0y6JVkBnVZ3asNbLJWm/GgX00VJN9XyC+X
XiXbvjz2y4SerswwsDnIg0LMJSK0vBL5TXCm3j8+UoHuW+O02clAI+Lhh4Lwq4WszUoTlY5FmjP1
s//ACoW354/x3WHNl75gHBoBgSvqKLqBrjEv1KF5Lq6bCoJm6MP2ByClLRGzbePsX55C8a/DI4WU
NGPzmf8kM1YwEEk+Z3NWrcTcHq8IIJgkEGYVIjLpROcxwSWozGBV1h30nLUimJA7pYMFEBYH3UKo
+vy7TtFVA9SRyBoNs5EVEotIREcuIkMWqr/u+beXZ7hcipzp0Hy4DTuLSibvors5/aIy560dGZ/9
B/sv7R3Odb6Wsxkm6nu8guDhasxctqjxFpRAUI/v1ceSr1eIJ39fLE1JpzAjpSjNHsAcHSJ4WgOq
drnzc+KF1dCzR8/OZyS/6S0grfarx5r8e5FiNsMzJXQTpoen0smTdLXDSnWfbQayzdoqyZuXbLXY
dYlCfVvUvHf92C0TCo63GbA+z3ecbGdjERkNaLjDM6Kr1RRziGlCDEFuDKUt8/E6sdGskFO2O35b
9yIPWOFiAewWIhpPlQHODyNjhAXB4iZedxR9f4hV2OTiFvncDVOtOeOCzn2+3OAt8UXRdMtMFnnO
JWW6R51ub7JZQBlkLBcLoUz8U7XgcZiG6U9JLia9WQeUj/v6YMes1ppk3/4gcvFlo5+PfbnyewdK
75iZE3KmG9V/nW6muIoeOYwV1caadM4zaZirKo/ss6MnBY2V8eCpcZH6gmMzve4YuF/rjouBD6B0
kB5euYIvjg8hK+twHlsxUyA5n677NqDJWBfI2YYhBCCTrc3uuvD1NjZE6Cz5B8BfIHtEtf9ZN5fw
xug90/ZJUsIKSONRGH1FOu9+G6e38c4jP/5JO4/8jN0NtjCPy9cp6LLoyVF0ETEwynJj/zDErED7
mO++RVGq0r3Ein29hEU39PdAZPHfp6dssdjq7Ff/KsGzHerd+Dvrcp3e+8xzryKQg5fskCxMVQrT
OKbeqlZw4ZOSr2EkzXYAATUGDVkFlvTKTqVg1uuvxlmfmaEeLOUA7ZLJd0RUTVvMAbUrCcGg0Gd7
TD1TXO4cU7bvf5NnhEw3/uGe/7vMZ2ivrTSy0fMukw6cxQtNYpn44lI2vXCQnptTnfFNDkAci5yu
e1kiDiBLeR5VT9KBlzFJR+B4Z4IsNzjgfq3w1VSqz2ScZalyRAqZ5OiAAD7zUjo+mM0+HvauMPWL
Uf5sIILWZdabwdPrurg4oAn2j8X9DYh4HvXug8+okp7S/rLuiy7tAnMhtYSI5p2o6PHsWhf1t4gF
QHOTlCDd62cXUtl5CmDB0qQq3kz4IXLCtcEkNBR4+G6F5IHv1KT5bVevnY/k/yraQcAgHk6b78eB
Y1kpAVPnJPmSKU41V4qZlw8tz1XXc3ozNz5Yc9bS8Xj0PGA1wj1zILW5l2tGWvapI/JrtozXKzUu
Bepwy8Z1mdPvB9AvnRoZ7gmPZ7BwAwDiAb0UbCuKWHzs+QH5KT33l1xPsGBbqn5VOM87lJfua1VL
YcIa6xavhYjcvf5xJYOQNZoOtchVR3xCvDdPso7OE6LSImv75YVW+EDmBoGzHrxOMpOcJe9MDsN+
66S1xBRaOfSoUc+6wwWQ9xeV7KlML6lDXryG0Dj8w/sAvKw1PLeeDjzuo95Ib4sMbGGmvG6NJTxl
X7O81ixggT7lR20bgsG5lf3QPw0BFk3Wr18tbVk8isogsdbOHfdTjPU7ua+im930Pas6QKUUbNmv
YOAlXDujUBiAibGkyTRHB+tIFNpAfFeck/e2UGXRl3hu2FWz5YVg9V0ErgeicjxjnNnYs9miC8k0
u5w8ofoLOJzx0EqTTP3gaOANiel7gjfsal/he4yA8fdh+czj+Ez6TZjTm6iH17LFhKghT4RP01AT
QafOhJ1nKvrlsSKX7wfkLOx3+S9WdA+Dl8zc0gsmEUoM2mA8GptVJwUbjV/euQTo/hEony+LxrSw
SA+j5EqFUntR61jFiC7u4D9vsRzeJ/GSkV9+vswuvjvFjtC8S9iYHfJmsqdEwas+TSRMlhKvnUY3
s/wh56H7QwB7E14IV7+fbgo8OWhKNyXZ+NOtbiwrNImDgqQ/OcD+nDqv7aSa3z3zOWUznDtVcA41
F9fnjH7QNbxrpeOFwD6oSaWyXYWLD2b7/RldD9Appe80YD+kjFHOr19iALhAtYu4NMawXhUgsxkt
y7Iwt/pG+gEpYXoYP6oU9ppwXhlIjPJfusbQR4q/V5u6EOffsMsC/3MtXhwjEzRgdIrPk2aHl28Q
MLOr02jQW238w19Ae2ZTNRPsJ9KkD4T0CHyJ/zFTAdSPhSsA+RoMKgQEcPCbltxos3easwwNZ2V5
9WAuU0t7cYwNKuDC3mIwwaF31u+klb2LuZBLjERrLun/VnRlBprMk9UfITbb8ymAoF1mY7Tw0cTx
Cu7ZotnaWe/exoDT4kNBmubgX5HqPYkhJD41MO3scaCDhX6CFPHK/HN4qCIQ5OprWMRbILvwC64O
dd3mHD91zEDb/+BeAN4/kESSVY3sBhTdtd/zj6xZ2jkm6xXM6vxceDfc+lkRLLEv2tcIuSEqiyX1
AWe0FtxQZWMfC5YqB0+i5MblLZVgTNtdfrQlx1IygZ0qPBAW5OQVIjcpR+p/pJOvJAsLJuJmmxK3
CjeAwAtIaWHdwANS0yqfu4bc/xozDx+TQ7GRZzRBxFMozcRsp9RMAKDiAhNgIYHo1TSxa/CnGmEW
IQ+MCFD1rm+bIulpzoi2ezig9J3DyfUkWtfNCyIfHaV+NiyNlIpyrBbBL5Hi8n5csMwn5XIUsWTT
QKy9XKVKmF8TSV2e89/7zaHXQVDXvD3cYa2QC8hSox4NPIigdSjdrloKtzvf0nBOMAs9QlvDLemp
+YiFd/MIKGUnVPmAP8U5RRUSEQFx/KY09jJKOY1/Ah9zHxceN83a6Hc3QqbOPwsTD3nuiLUo4wEv
AWXaWwoZVU7AixGlMq/cJxRtuk9/naJ5GmNVX6RkD7JktosJpnzORdLHiMopmUu49+XED/xvJkE/
SFq/+dv6fVq2lRQrpa6v0Mj82O6K5rsn13y1UX8xLrMvpXW1T+CkjMovxnC2Y1/ZXGy8diQ1pYJe
y9LT1JHwMWjUu2+pcR/D7BFwj7Opko/Fx9Fm1U5OlECz/CyVygoUTzU9wYq8WFtMCCsQxA+llRGR
O5HRdSTBMyYZXLKmeyO2rqQb/lPejYtKdd9z/8L25s5buVgoJfRpZa/1db3YBlzOqiwk74j7yJ1v
70nm46Q2ZqQdoeSfHkgtl7Lm+0Z9grssTpac69xWbUjCPzFeMj9p7ZA/ySn60bPjMGV+ASyIeYYY
uo3N4R0f53idaQHughAYXrkl/rI45RFptzgo4TRsCC2pdccprZb0l/ma3a06FOqJrUfB+TGyIMeR
KZaK4X3UYkJAz2nimjtW7waHnMm4ConUOxHJbTIgtqqSz7RYEPifX0VfyJUghi5uqjB3KcqgQuRW
LkLlwVX3Cnf86zmchnxNRY8nN5pYtK71selGETLKz32GZohbtfr/SIpBu/kFvQxlCIyzzKC4SSCR
h2fwLEosiNT7yr8DtjLaEQn687DqJksX+6pJLkCOijhNvk+1Ay84nSZLVnnEqAk27tvP+kCFbf6k
5x4/JWi/Di9DeLsoPhsxCSVyJ0+A9yOwceWlLTBq2TZm/00XqDgThpsUBMQBB+Au1md/iI1gsYTb
hlfgqmU+PMuv8J/73ixxBwteQS+BN3z8MP++lNqpwgDH7eT0c59XC8S7lOpebhgg/3tKN4hPoj5C
Wrnd+r6WWitxDpKuWrvvQ8ExLh9QFpAwDmTCcsQiXZOtO/5s87WSIVpa1gpzgaXAkWCm/uXec03G
paEQDrg6hQ+4ekDpRpy+JfBMBp0IcqKETNdjJU5Iv6No9dROL2CCND950DgAzRJ+jywDLJKNvXXi
0oDhmz6+2z7PfcSqL+aOPScKWbLaNpLSI6bes8l5Ut0aa8ONaH3PVJIQ5SoUdCKtQ8gg4pvGlqIw
bxpIx2EhxgkbE6s9COp1pKLtpsK9g51uMOwEouc8lBhA1bWpjMebK01A04xFONhO78DRDahy3pvz
mIZR90PvA2d3IAgZHvp5cLDKF0uBLKgC+D0CEhRqET4Bdy8d9O541PZhk27/RL75CowMJGmEhFc8
M38BxYAvIqA+sE7FGIFuxCL7j5BU5UBik3LpfDR+hfpJja41rURuhF5dgFAuqATMyAKSuELV3Ill
e6mCHm2ffx1TCXwfxJUjfN03KnwAfnuKKE0+pFF62BCTqewYAblonHBxaR9MafYKNCt9hjLFwCKZ
szIGmh85pVEiLcBdxZ436MuAzmk3uxmxiJyWd/T8Jhl20+ujUi3tIxB5ejWgI2mJWdBYIL9Jp77G
RpLplMzO8f2pVUQXxWjrf+fnETSUhUuAQ5dzsr5fKyM/a066EtVIyu0ptws/CXF2Ov28raDShfbp
cdrHjq6odfl8I0GPU8ZPPyG1d23nX3a2Tc0ToWFdSuJzGyxMd/ASKhGrn6/ZEMMggx37/lfVem0V
Flh8dWJbbzpf2f7vtU72gtB3WZ6SKZ9fsF88dWB4mqDz9PE0B4hDO7Tbkg4ye1eKcrAJ3+qk1mCg
SYH7JZKMgIggUy4H+gVFZzMxaEhbxP/nZLjgc/xOlscJoF15mhbxenwFRIHIq7sIiv34Cmw+NONW
QxQqGXO31pyeEgdjdeyXUfcpJz0kUV3J3aVIrdFIRpjqs8u8At+KLRcnbDYqczV4KpnLv6A7QjA1
VJtWu7Mt4buneu6gaHJSvv8tc0Vo3Bm9tSWEzsfqxrDxJE7cmhHmM11+UZBOiZtlYHL4XZ068BG1
up+JCUIMqKvDmiyFPqxoILkRZrEKWj3L2qNF2j+rjjuUKhQsNqPat2qad42S2WC1iWWMKfKy6ttx
FDV9O3QJwJU+uf+uI/fBOnsC7IPHhpXbCHZNmT9JJsxEtv0zrYrtSRjiL64jZpTBJAMIsF7dLjjQ
WOplkImxnANCCTyCYNPP4+ZIuDUfcLKRm+1VsDbZUFIf1HvI8VRI7IzufA9KM7pVoss1SLrYt8fX
JbiT8gx4YNdhOFL1Zr6/WHEZARjM/aaGforB+CkM7iFBwIe5Ogc7hSumK84Q4RzAnNSCg90QfnVF
5PYYsoJFfp1asGIscEIgFH2T/hRPoxx44l0tBf7ZCKHWBbyH5icfQZtAiJpTwjvAA1cc+Cee+ohj
4puldeZ4R8+7KbyxS5AuUqiXlIYVfRKZv3gVjiHDPDPEYRJnYQSkqX0ElNzJmAvowqT8EPPhgIVI
/hIP/ShM5VZ/mXFxiiANSSlT8HRSd+crqevH2DjI17tvRXWvPqbPCeN+GMiicFfM9qCAA/1BWGcI
7vv5LsPsyT+GloKKYDgTjM5F0ZksyY/cauOFeqCHWsmRGmHZ4a7iMfpfjKJMB1cpuhwhhOJIu8aa
AaY80GU+k+5kfMER8LttFvDD4tNUjfjho7eqh4IORCCDiUeGdT20ySlWFwcrzyKsQZXgVPx/VU2Y
UgZ1YixfLTkPrNB5o/zhShamxY1Yt5P/TSgFKMOmU0EKC2+fkY75RO9lw6LEuOTWxclOyUliuk1g
zGGmkTiZlA4wuAu2EwkcK5gOp/xvYI412/4XRzo9oCIzI1FWB+80g4O4w82SBBBgKcAWnNzjrTsn
6DYljMlC1nCbgKDF7Pjg1elciLqnZVX6uF+g01yeru8ig1as0GjZdarjJrr3PoCncRYjzbkNd23e
HjL50iBziIlWXG/pB6Ak6ssPmK70oIavysmeAv1MHVxsmUTQ8Wl6PaJbxtMz/K0Y0uh8uGOH+R+a
UgCxE7PzUIQchMZK5QYB5pi4jWI+BoGUj0/FhiuBqxd8LWjtELbMEzBAD6SRzIDP7JhDL2sJ/Ihi
kjBeXpnFuO6SpEdB1iHCaL3gB1N0s1Ar+esoC+UDnUvB1e0/XqfkO/nsFfINoh9oT193JApttQhP
Gyb6hIC28sAOE9xSPvx/SwEMYzfO1zimFfs8Xf1/PvrYOA3HX6OvQFtBl4DU3803uV2Qp7En7z/V
I79M4D0MGXwCk83zSqkLyBSOJW/wDhuHgLO1EW6gpJOsvyl6R5I6DQiXMkGbMTXBPvzGlu3cW1Lf
qsXUadAihRILS1mVBlBstdbgu28/rdECMIHicmM/1lTlyTjsGuKZ4uYEL3vpUinZkeoumS468ysR
mJcJNlnjjOMEeU3HV+C1Zq5YMq5XQFDONEim4CVYJ+gT14PSMEatxADCXJbth5hHf41q6zn+Mek7
IqNYWpI9BJ1NQy9LFv8TvjBkC+esVmiYOEoxsS/RiV6wh0YAgxO0BvjWnIqenAAqulvIJEWbHt62
rrb+jV/18D5Pu4XEuLroCtr3sIwiIbUurZ2e7rEkPCbhr5oew75DOY5hf4uUT12yIx1tiEtJ70Ym
Rdc9Wu8uvBZfK0+MGTRULw9U7odGX+KMrFhpQgEv3uMz9aDlcgagHyV3YRNvb0QdKCNSVqt45kwF
oc+JfJ01LoHao29Mb+zeztT2hJAMybDvMAQiJ99WOocbmtqTDoeSG9pgqITzEB2o8KCKNF9rRx+0
D9hOlaEXfDKYfVJlRYLHK444tPuisjl4vgqPOfTizgeArqGMTR5I72clR0dz373sXMpsVMkhvBrN
QLG4EljJgHpLnNkhKPQLX65sU72XK9M86w+G2VxqKekNvLzMWLNVXeZywqJmEYq4kHD45ve5qJke
B3mI87bd+8FzqwAosZsm+JeEl4xx+NAe5zM6GagzJoHkVO3B7/AAVibs1u89fjgsrLUpQgEN929B
y+FL+knHpraCd0mRUZgmIkEItuzCPnqonaC+2DbvYN+1AGRMg8X6LAR2y6IViUxBQMWgYFM/2X/G
5KTd+8/+eVb7rVUC8Oo4PSttUbVCyxcqXoJ15SoBLHCXnLE6SXB+zqKSVDhO5ILIu5OA1ibg+qu8
ZxnAEp9qHseqKzeEpI8VnH5CG7aZ98bxKq1V0i1rzjB/86RILeBEhADId0dE+GQZ99fdC60UWGiB
rBt/XJvIVAvbLDs/BYySNhtALiwM59fPy8fOzD91uVKbRd543lM6VtZor4NoEvLMVz8KJli03Kdw
2WTj1EBnCNLezuxd09ajys44qWa3h5RCUFFgvij/Wa9osuxU63Qcuu+I8gcgKAVxDRW7ZwKTMSZM
cKSZqJ/hleqo6kyc3Vo7oo15R0TM7IWqNwJJh1fFN0YNy/FHUM6/hpV0dtx3+IB+JHva9tqErPfX
2F8SqJ+dmT8WUoQlhlJN4Fbc/oN5N0HFzUMLxhA4Ls8UF13bmiSiIe4/5vDOeyoOYIZgx8uQfsxe
hdCkLU8Mn9ETK7DAG5OJ58enKPP2
`protect end_protected
