-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
b8UbOn5IVGBop5lQalizQVQEiz28l1p/SYOvxtPMHzm/Ma+auhr1oJTYKssR5piHpD2WELknELbR
ku022uICSa5QgxSqTijECSryR/fH6ZmHqfP7g7DtBAImf2eTDv918YZeEkhA5RfF97PiFA6wYssw
mjN9QJVyTxi6oYMdObEuWhhd4C5S0/hbqUG1+VJx4+Ab+3clYndFRoRQdEYVg5u0KDjGHSytIjcb
mzqpeAaNPIedvpvq00Q/2lcEYeVeqQdUChNsXkPVIguTq9rSxahnw9G0pQJGvrKWIIfVoiXzhZoN
IgSPml2OuQF9VYC+76sEXbXA63ikJKh6QbMAlg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 69584)
`protect data_block
luO37HiRpV88FwgKKj+4zW8E2304DlKZBqdVKIWz4obzn3ojTRE6m9XU+YymrKDfKAkahthm19cr
UxVT2HVhBjzb+t2ZkjP28hFwEsLKAupAEczB9nOLLrlP4s70IB4AzG/Fn8cDrf65KD6fPVCq/LJS
QcGt9qaCrulq+DKNBBhbCd8F8sZyTBUFYHEllTGZyqfhFPcAgb+0/CKtgrorA8ccbh1VAhh94rmX
7SQTUf37vSygQEK6c4VUQawRURyHWfHob/NNw/9L3zXlplg1X7R/Y3QW/W/9y+Uur3gaDjVW/T3m
GHV8flt5MEZeS5WZbqS+krzdTUAMsUNUgrmJir1hEKG3+6VA/tMKXYXWPekI/SoPGTdhOBuZkbv8
W0b4vNw6GkZhjRWh+6/mhmOzXR/sydKkXaDG7cA/Mds/jTyO7E0KbRoBVrZ/Jtfl29XnCM82bV3C
50qiHaMs8Xy1ijY8Q5deNWDpXizIHwwxyMCshUtft19J4ykhudLiuq8pUHJvLAODTc9hNY2AwktS
vqpVI49voPL+hwrX7i8zwU34d/2x7GU4zY0yiE7asazmf0qo7ZehYuQHDhO/2EM4rGlbEpOqrOp9
MeSU++UQaG5bqOVZt3Aem6b3yVMsdU9P9Og4ZulplT43pNZd32V8KvyDTOwpQpc8yHIWRUew4EsN
tnrzaLLmbDdmtOksJkz8CmHo3U9qofddGezTrfr+BRa36gMykSeuCdzho5A5daY2sBpzOV5/wxOu
7U389wZdFWe4wTKusUWc2CPpTRJLm/2Uf/af67heCQwdiTx89kW2BDaSChmv1A8FcX086jGK9jLx
B6Heo3JoUz+kxR14M4AjjmomOGUAhFtfeaA4OXVVImABqa04XtEEBcGXyq5/65CLMaAzoUAIHWsL
FzcI0yufTnmOCsSPOiaCbsCujDUv7eni9EO8z4t1qo1PkQYrIMukzbahpRzqqVUzD0BJbXocEJAV
+mHcfZlDCw+Af928fxLdWoM5oDnsvPK5zCYVLhU1+Z+UueiZOpA401lO0+JfdHOJ2Yvh2glgKW9W
ADq4X/pZbmCAOPDw20ohNdU+MJPth+vc0UauHxF87aEg++LqgobLzxyE12CN2RwxWxsfigne0JhK
DVUJW+EhJWL/n18FeaKSMgs1GZMBB61wyQjUuetNQYup1UmcRBjSXU6GpniZBIPlDZzTUeVIG15d
3i7OcV+jhwQUEyqUxDPlPg/Q6aZgaB0yA9kIXmmR2wNPNbcv2HXnOunhDB74DWsVxbM0K3T7b/4K
aVvVzvUzwnS6MNWOaRURyw1PsVxFoY77P1rV17Nd5NOWeS6T+uIVIN2niMVidPGoR0hL8YJyBtkV
0b41XkSlGQh2KK5Ip+KhjB1rQUZoawt8e7l+9ehRIRTM2+BA0oNlmHghOLuAF4crvoMFUejinf+m
dwN7iLTlaRZf36g0ODxOjerYYpl8hGBKam11WOTUFvDwbq3aMqDFI7Or3mCv6oa3xtBDWn3Hnqlb
P4uQBEq+0DXCgsmDZxuJTe/pNMH/ldwv4ixmFeGQ8b19mIKr2PWAD+lk09wVkAIuJny7hEqCfSkI
ZMm38P6CjuYFMZQdgtIpJ2Y2s7sZwTkG7H41sMjds3PesvgZsIOtEa6QIrYKGxKlgAMVq1vU9Vaf
CDeP45F0vfxurX46kVDKOs49QqNZnkN7cvzW38ukwWlXTgB+ZItza4s4FvE8YgbbeUip6ZFmYA3Y
E/HPw27odatNF0raTEIBEeY437d4DmowFDaoEK/totFWbGLNoE/8qcl9NUyngoiyYjvOImtPhusn
gmPBqrW86kmfLHwZGBeR3i8s4zGieiDmmR/vo7lFi9T35KgKmsXu/e8xG4KgXAZH51XOYqy18S31
3koNFu7/twUC7EOdLgcZtHukuT27lnKO8Qtd0LKLwZ47ZhCaAgQaRBHQAIb0M4LEb4na7UmfDy4O
Ml9SEfSSYog7BJgGg3cgXsAnaAIBs0L5MWThcbFz3l+sYpuhahhC+6UZmRp0Xk9w8/N3hs9g5Kqn
Uil2g5Z5/Ml7A0RLuIUNuVz44QP69RLNTUnjUfNOCuMcu0Mb3kin2wBhCAH+iAb6w2tyfah2Qg0J
jKqw78c0KmaEwIZOEHSSk/I6esS+j0B+yAM+aF+Oj06fqosGc0esF3xkI88lnNfoVtBM1NqmCOIY
et/RroyyhL6NRZPoX8H478pusJ/SwVPIZpdtn+Tn7rBqSDNf0nYp0nmRMmp/wIzPMveLI6lGUvJj
CvBjp0LkBFey8i1XYztcEREy/aAm18QNEkRhkC7HnhgJWdPpdP6oCgkSy9wBbZhafNBjVdoH9JsN
VYTCVt56l2GR6j4pKPPaHlOfl76j7+FPx2ZaoGZjL2qfp8gnBFN2VQe/QHGY4MjzoUg3kQCB4FLE
0zlA/pnnfnmai3xmx/MK4ox35GmSfGmmjikGZIH8RBTs7VF+77uTMlTjd//Wjo86aUB5l4pdXXWD
ugum+itrrcJFRzIwe0AVqIUF59Mz2gC0Ei10jCH+EiO9aX/L36POdSaw39C5FfgH8mO5rnC7UGo4
0jKqJ/JT6CSv6WmfUivEGivdt0CAZQp32kEVNS3PV3olR+Fr+D6xL6NjZjCt1ZnOtUWn5OkRUU3n
qavcgB8oe5DHRADYvo2clBhLLT6XFC4cltTuC05ps1L9nj4IPmW9N1yrEc36RrMyDOcjRJ8+v523
6I40p0hwUr38xemNe+2CBem9+ym2BMRKDXCF+mdxS8iatKQKOJiD4WZbcHyOAw6Jn0B9qZEElrR2
CL1Spg75VWod0h0seBI4mSfh5doEXrOepA9LY+VSWANrg5Ak6SKg0P8hl8BY0aHqgp4yRyb5J6LR
jv2+fwlzjNosgdH8Os+RXqbBUjNnqBAKZ7p6P4l5Q5aTsR/9EDKNM9Wc6ql47Sn7XSKmYic7TZZa
YevluWXaXP/WardNL2bgNCYGulXgE5snFEpi0zSlUn+Etmz7HXmBlyqSb/DH8p+77qVpEvQ+6n7F
CHu7KQkk/KpJeEAvnSbdyP8bn0xGhQ/jrEoMtxXO2/Q5PIhOqZw6n6obpPs+zNWCH8fMnQBjytwn
BclhSS6hk4Hz6PL7A4nw7kf4IE2llkHRNs1mgNhrR4l8Us1OMdvFao8/bNGwiRCflelrWKW7deiA
cyvKz7IRT+Lq0UtPyMsVS7qaerGfPrUy/Z2PXLDMkm18HQMOQ9bDX/r510Iblkj9FFDSf46W+kKJ
3Ma737Cqd01ol6oD/3weGL4mURDnFcN2ApYbYM7BuL0jdqTTXyaCriyKy3cgP4orn27knFKXwbis
F6ocrmBAAMiBdnaTYE9UX47ZtJW75z5iZzCxPIEe6VJ6v7zcwvbTW9TgKi/fDfU3/nkFrHqFwoYK
Nb+qZle310hSg6xxabAHresuHa2glupr8DGlCk70Dz1HuV1slzlQdZE6ubFrrfIGrKePaqCFJQ6P
99wdmMqv+fJeEFLQrj5V0/8l+7dfJpJa92c/Ii0ds3MEn2BILASSBW5NC+hun00Sn59Zu6mW72Kd
x9/ywEYYMxp1EViD7DJA9qsPqAXrL26yVx7nr2A34iMrYUkJlgU2KL25bTwOHGFDX/QJmW4g681R
t6h0pnjgplfqN9zky+Eixxa412JxZOpNikM+bhh/WA5NKc4dl3bglzzN94PmUCVAgcvNKkB+i7ji
blmdlGtZlStZGs3BA8KeY0i5+7OW2tAKf8F3NnAADEaP0Bur6PDVKycJTMryNRkhSdsb5omPNEiI
Id1G+524CaXpQD33dui5+CY++jEk0ZsWBs91Mf98iB9GToT8qrbom6JQgb/x00ps7H9jOvDP3XsI
xddA1OF86KSmC551A96zx5vSf0GGg+6hkmJd9n/l9Q88x6H+JeSV21vAN0lUNb9/1a93XJgO3Ku/
DOC4+Xjbht1vHLWuKcVBV2mbjH8KeszDIgxapkAULkA12VzNLL4IQiSfjZ+4Tb/b7l/685OfPiNV
WJcCKwj5/9dd8DkjfX0QDfUquEBvLzqFbZScR8B0BOA2TC+ytcX8psRQGu4hK/YD7mx/XZ6J3m47
7dLP97JoVGJrmqO6T8YP19bMiUoi+XYRXHLBu/4KzUz16VWxnBzZIxU+sOY2PcGqlw2QpKq/UWS9
g+oOpJ4Baa2D1bP1NEzn55tmrCWcREG+fVZczF6vNfDT2Uz53/eMkogjVqBIMEpGDEgAVLbuig4D
iGKGs8uJMi3KfZc2IJAHrvvpp+vj5hsyZZxjydsv9tFlrczWH7WHB1uYoexndMVLi48hi9CYPchy
vPiEtk9K84zAgBqVkkQTuYFei2AuYer76Y13xXkLq/R/eTrZWVbCvfxntojQdwBt1cg8ZOM6oFR+
DWFe9aLdr/g37b1qxDogKErlT41xuH4SDQ7MPUyfJk/MVndY1+rwkbD0Nr1T8+wvKNJ5XA1/obu4
r0iZ8olBlDY+MmBbuooXdrUSwtHz+z6wLnIbSLMwqWsFB7dEpXVLmbZlQWk64kpDtMc53Z4S2uuq
qdHuK+TeSY/ZA8t04azxL2Y0KRtwe2mU0bY9R/93T0iJQqVo++nw80TfSCxH3Zypf+DatDzSqJnS
aB2f/Ldf8k+ZOREiHREuV0/V9Yq9u2yHj/jCDCkeDM23zjhScBOfYdDAddhYOBVBnasCIFbjTRo0
B+bT6Z/p7rwnqvRzZhgv4YVd6sPlAcm8PiK6pcUv13vxJij1ZNaNCmAx6Jwtek/vRv066AHsI7ls
xEOu/ePpyTDxGNeHnozLXJ+Blpz4YMD84X0ieVkGWZ8O4ErjHSfH+0QR/ZY+e5etRgcQS4m5Uf58
7hGlvw/wr+qtC4vBjn8TVN9CTjOMFlMwaOouPE3x0up/vK91Z3ygHTwNB3WX+vEMe30QyZE4dgdp
GidjbT0rXe+a/JIA6jmcVPisVrYvhws6A1Vk8KD1d+Ol2WtsKYjG6YZuXL7kn463ol5LxAVQo0sQ
KZHlKWWMMeMFdlT/4gFYV+2cchsPQ8VulBwY8g++gIH6bgesJTILzQAuTOTBK2W2UBK5tbdEnM2t
FMrv/Ivu5IpKSoJS6AUyI0Gx0ogFRcGzFuu0BtKj5W4jfILLr815RHaP9PJMc6Ix2yI23Dab3v8m
P8kMEkn5Yr3dH6fm4JtMaE+Y4aNjNLsYkEIqs8fRRfXDqTgjIXG3/2W4rbMbK8XzjnTTit4Km0lr
RG7KVHPNg2z/5ldOHM+6AbdUNgsA+hrLI1wm+9P2p18tjEo7oxBg9IogPXvqPN2jxxKC7qAszJmk
odUnVeAmk+5a0nU3f4GitpnMwcE2+DN+qCxH9zHDnZGjOnk8pdgFJVtI3oa00UNYUoiomVqmKcLx
r0fMtKEpEkHtx9MnalUIfFbaLxRsFjhenEXauKjyLNKEjqhf+U09PLc66CcmSh6/bdlDDfifI13i
6dBjhv2P5mquO9w47P0/vnhHvwfACYQfKrOMA9BdS1JZ4dJVrhD88ZHXJzOapFz14U3ciZ4rvOLH
evdpqjE4uWruSWf6kt4dSljFxi2NS+i6l+cAs1OvLeo0VjMQDjXZpXCgo4bCMXjHCGTznrjyxnwt
jmvcpMMbp4wPpC2p9SMgUTgKkXn7uQD2s8oy3ibpWtE05qf5AYfhrnu4U/4ZF/BmHfaXNLhPyWwI
g4n3dZI9F98mlO1tOfi/o7SJaJAhczZpvG/FTsapIPL6WvwOp7OLT/E+ZxW1CycqELHOwHYGBk9k
0gay1TZA5ujGelTIuat6y7buCIxDzvFwo6nlpucIXiUr0aVpxcNe2Pel+N7RkfU2Weth2tndGUCH
9iQ4uHm7TK2mBdp7/6AsLj69E+cPsELfex71DA5XhJ4BXyHK2RuG9c5qbliPvzGY8Bo9vfNj9Ccq
fcCm56JtJJy0aJi2WjPpDSNnMaDcq5ME/DmPeisa9M4ZqyDqo7sA/UO0xVbs8v6qTatCy0YXDhmR
ZqNJDSo53X33mNbvCqgKGY7UariiZPl/LEy5wY4ao5EkcfWCxWajyCAuEyhmohAQT9CNxnhb2+rz
rSp4LYtVVAsET9XAJ61Q1EXByc7KHG6ALThFRaa1nK93IHs2/SLXA+fwh0oTGYt2otttgoso6ckx
wytobJ/m4VnxBeslGzMJuO/sToE5xqajFap8JFdN3uMLMO9NEeSR4OjyKK4VYeD5kgF+o2zYHo7V
uuGbsnMWD3fcl/5UTIwhY6q5Z8T78Yg4TSwxuI1jqrXL5grVD9lEI0aV37f9FA05X1uep9fNGHV9
c63gI8VyGw6oMdbsunYIbtnW9BKhRtUXWpLwBS/zI9ncfO+nN7vBLDds6piu/KVtAPsSOe1pH84I
WPu4sTYXPrOgt3F+ehUr4knxN+ZKhIncmmQv2Gf0FH2W23BdSttWEyAQkNnpHsKmuV4dXIOtkGhw
lVpXznnLoVT8swgqSM8ZC7lI/xSWhF+fmkDmGpZeAiEP7qXI/wWNfT9Z44Hhd1UuAL69YIvbDwgU
yy1zg0uotogWdRIuCP6oe7c2a+gFNN//xOdA3hoLKZ3JzFzWTIS/2o6pAPbFNE7zD1Z9521uYj9I
0d4MeqXtPXH+RFlRTHYVhwmYOTWTc27zEMVICP8dPCYJR48vGpixJ+9H52ioskk76cpmHO85Hh8o
O0BOwB/vVC2BWF6y9KQMy44T5vSDwDHEMgGRH7H6KVbfPk+vFw8VlvkOktXeaw5U5ppdbxwcwHHu
ivAGu+kLgFv/k6iNJDGhFbezFG2fFv1P4X0xWXgEFEyKQw3/JaAzZkOEWvzKnQEaeS5GSTdb6vmK
NOXscneQdhAFcWpw1I2TGyhis3v1gfCRwF+y8cTAeEQaQwDinaoyQGolo9J0FT4BOYkpOUGgr/cp
9MWFWiGIvU/XpTAwobMi0ZRhsjnRqx/ztLsJEkI6bQZiaB9NQzQfXmbfw2zlseViczZuxbsNo174
vz7us1vsWjfBRBuaIpeQxzfowRjVqZseWGiYmIMAuEP5n32Xy4ztWV+UzYuf55N2MRA5q++nGc+9
ho5hmopUdldNVFO9IwDZphlnPsEivyheJGxUM0L0GPXYjTMBZHYmTv/E3XvYStw9QSQFq3M5WfcA
k0sZrOk7UYgqp5eaVr691dRl97HQN0taOyuVgZVZI37Op43/1aOWPCTHPNN0Y9spZZgHSLU8QU1u
UKX9IPnjjY/eEBXHD/ij9DeNgv+SzwcfQgTDLkd/1K2zMk3yDnXTRYnNImd8hv9t8QxHu9BXEomG
uCNd/uw3fZ9IVit+IsEF3rH0ZiZ1Q5VNs9weOIAeUqw62JcByWP2YHhnXc22C9oUYRgtMSiq8oEy
bR9TABBPSLYCFr1tACwkWKREw3yM9u6qcFqPPoF/6X1jn0gvyb0lbZjuraOsS1ewmF3RzYIpaff5
uDtUDtrxqw+pIRGo/h5nCyjRWElTo62xzsX6eaX9LyQVafrRP/BZLH/Xpky1vyhuKvltTUjLEoEi
zqPnMYQomeWOuk2b7Ki86oTFSHlDHE/bvPGtc/ENnnZhGVYtw4OwbHfHuj3fqtUwLSsHJcvOzQ67
T45VaCFHB94v6kSGWDVhEDmp6s2EDdZdD8HbL7+wxlUsMkNqbaRipcZ19b5ugpPyegpqgqIBqap9
oDycjuR3iqtAS1q1TzUW1RHX0WcQEqanZNxYy9yh5dDiOHkt3t5pv7pUuuedO0wi3XBFNycwPFRB
iI2OsPlZcRENzCoI7K4jtIxitfD7HIebILOxDN5qaBF80jzqscqA8nawpKv36MHollAZfbzzf4oR
Q0zqGEeQiALmd8cCwolazqKOT1wzTc1sB4m2NCy/e7RfEZIFWHvrCTmhxnMBhCCDmlefwidM8o+Z
e9ecy5zd97yqMEEIX2cmSbr98cOBt9HzD94kt/KuLxC8bOD8TaOq82cT6TFLqkz9ots8w6vY3nxp
ORQ/xfRWln9MPZYjC52mRMRv5XEHi+i1jl+EjBQMWiBWgFewXv9d+lc404epqyj4jt/dhnHOO/fW
vYLqtAGYvO/6hWNkUHwT1/esFCXu65w4ehqzgPfC3e+ylbWjoEEkqr6LiQzacZU2ni/9EXYu0AQ2
KWHQybfuxPdb39lkTrkYciYG+FuVzP0ndYSXF/0W4e3jQgyRIEXW87MOasQOu28FlyM9U6BsSFKp
sp1gRUfXLQCN5aJmAHRZRk9d+n1uVSNdkzs1eq+CpvHj9YZUnKnESWTeeeFPcI4HCXhNP67QR9m2
u4krPFf8MQejFs5a3PCo4AS1W76YYYJkP/61JuVC+co1euGmDjvqEu7KeW0HpTQnTB/6IwfBSBth
jFIww/HVa20YdqKmrBramkokyX7Kao7sX2uKI32NaG9QcGhiWGUFBdG5IB+jPREJzjUBBDqShNpX
upCneAi7zPUj8kTma57Z+BOHKSWydaQi/M0J6q46IQBiEATL/KSgmHfdKKcD73ikK+8IPeKQCrVo
PCNnjYxHDuECOO+UxgA3IxGNE8DS0SWNOERvWbh8bbxbSgPvCuoXgoLYXNadgWJX696TCDiSBr5r
NeTiCcplVryB1JBZ40yZkuhFzgzNdUPNhH7+rqX7U+8gdZfW7/Vm2KAAl+hbg62W7RsYKGJ4MDEI
Uz6n6X26mCYvOBbSN1bWoB9RU8MrfjTpm/JET4Muly5hkDqAb+bX8nvuLWD70UiWqxHkU7rAmREv
ZJLvStd5AwWQHeUepFDCQMYz3QAa6gvN3Lj85ADkpc83GfQiAleRRfNxp3EPIKv+VM3au9CSDZOx
rjdWpwvFHPgSXEV2L6bj7jOOKQPT44gVDoB0LOJrzbZO4ZIx8gMqIBbFPh/cAmi5kL3IPUzn5FsR
4tELAIvheBN0cz2WFa4VaDtjwsOPq4v8Ew9SjNcLKewSRe9KV7RrNDW7/UjKwZH8zVaCgev8zeD6
Kim56/ljThuBOmqStPBsae3jI33aSPAkXJk101UlX+2Hlp4Jz8qZPZJwMtIXxvFELEN5wXAJ1/bT
sflI164oB4qwN/oJbgqjaweFT+JK2W5r1WU1Po8niMvnJF+lZiMYhPPUBmGGwC/Gnzz2FeYmUcOT
m+LRHwge18nRxf6PBLLmdpLE03Wiz6cTDsFu83+m5LiA9+l2ha+eQpU/EODvOdl+kNWfJiAfCmgm
abrW5iiPX6yXubse4kH9eP9vzH3FkzXkRR+VC+USt2he077MH6n/xtqGokDwc5K4Xm0gDgO/WMwH
/qHaiDdp8AsmlBM99I90Ip59/8YD+GtopJ86V/nms+XZEPS0Id2isStqnsTwGb6lDb4+ohL6y0y+
jeGmWp14cizHKoMONnC09DjUgRBeYxMqo0YrOfwhuXeaPVAMPMU6P+UV4hKZMkZlfUrf4teOQAFZ
CtXNsLj+6FE57LMM2NtDY4YED9s3Qr/sr9QomOhHDozvtooKzqYVYeZcMqPER4/Uz5Dle0PlZ8+q
RkyTXR0gxkWatQnsjSWUyGjUWEpBi82DHFzuCd1IC2krGDs4mRHIuAaImWPWLCaV0xh/UVm6YsfM
zBK0Db++W3gCjVym01zdh0JsPEhLYBppanyqMtZpK23x2yoCRSPwOjFfUG5E77YFyBkH8HrXcskV
FjQ2xuPcurGL+ayd4a6QLBSYJri4cE8n3dxZax9Wrm98lIONmUK4ryczKZtTNolkii19VfnLsTel
JZWvoUxyoS1AjlgLItagiXs8z8cXIgWDYgbWmw2Y0s99ldGwmxcp+ypsV7vXiCpyO6I6iHEPXELi
B+/cPT3juwslUEK1E1Dts1k68//w7e1NJOsKZWa2gZ2Ge1Zk7Pr5dm5ac2EQ+dOS6LylWrsYO9/U
vVTojlLGvDa5IpODjVJjPCB8HIY/Q6yDNEeBQrEbvzqLiU1NmC/oM6jhblzPTrnhGfrkDJgJug4h
ZnIsbUCo2WVGJUcCwKPXQSNOivcbk6EmzjHruDPDBJ86KI3uwi22Um0ecAcVrP0+Y3vq3H1pKAIR
ZXAfXySW3nKgpVJ665ESmC5kq5T2yp7siwwNcFesTBxPI41J2I9chAlImcQGfbacKRU1TDIypy1q
yc6dHqY6GIsznR9Ejzvp90SvZpG67bmxbiGXBM2RJVGC6l+BhmAsF2oUgVAqYf/rD+9MUqb0EnBo
hnhgkHNDnHkWq4AytvqUuAz9RJXTJEZqgU3DKUflGB+SKnOhSf3O3GA6/swq/jWrTD0g3z1AUqPJ
5vHqLWLbPnC0uQXKLR9TNZ8BgiKWIJxJYEK5t2A4LN92UTpbaobMgvglejXMpBiTY/v76A+wfJ2p
jISQhm/axGdll6v/IEG5ujiaaeDI7CwIOUNtXcbP+ztEX4A2xl6PTWVKdHMzNJh1fd5iIoyBpc3o
VVEC1QXGqtIX0zR+Oi2FiXEd0Q2cKe38DL8Y5mZGuzUmkVP8pm0sMevVL1Qxe3rKUoSTIA7xKsgK
1lGHWrBZI5jyH2GRx/MtkZHrlzoVdLBRfe2SeQl0G6vp1gq8qY/Z/coAE61zHMWS6p2e7VA+Ns6B
5vFVfEketabRPCbb5uCViO+0zqIiNImgr5u7zAzGfB2cvXwd6dXFUehUTMP7slPrc6ah9BDeVHaW
BGaNmUksTcHQ6Lq4flo0A+MZT5ZQm6HcEG4l6L+a8LwghLOiD78RXl3NX4aGKhhNtYXdjT3AZe/d
4fWKPZKxbTZ6I901qWF1oXLLAcpxbFCzcRjmSgjxCcw+aft8kOZsgiBskS/bjY01zW6pFVK/3mRJ
3Hdel7vbbZiTXrKsH0v97GTZ11dkSY6RtajVhWbI3jsu7gD6LVdF5Zu3yJ2O9cC19oGQY4kjBCP9
3LTiJ0eRu1k34kg+TR3MneF7TiJUOVpRS53Rp2rT7kHCIQMKirv+pNHWwfk4HGmA71Rv0fKkhb4O
P20pVJJefpvgRECMRE/tPK8zDMnzB7ihFhcgNwPGY1LwH3XT1Iskvfi11DVLMQt9mvIqOSYDjq2t
DQwdPd5HwKfJpTR03TatOoUXyzlQEZRWiTD/wPqxeSypkcOe5UdH3ATszhrnqGklbv9tCwCWaGNZ
P2ijLsEIYOnAiDVbIslr6zCPd8V5wtQCks0G4Ce46b4i0VBh4maA6aI+h+udsH6G2SaZRHjCKoxX
dTtn0zYaNvzSI++w7eDfGhYMOgEguHIRlXgJFfhJS3RQ4ZlDgL8oV4f+RUiE1m4Wg1+e5z0HfjDS
lMdicmEfvMFtdA4LRcjrnkPnMh435zOXs5RHDqFLm0D/uvJcn++lof4ZyiT5VrrhZC1xffWibXyx
t+lJ+KO3ShIvHGkZiqGfX4J94GD7QNl0jFSm73bG+nLf94kJklCI+1kYnUtRcsHatS5/O8UJ+R6/
Cx2R1iV6yEuyqxuzo1hI66jWPgMkZDkI4wVX+AL2Ou/M4JeL1Oi0nxEvbh86UAYeR29qbI3QH2L7
Iu8M/aU6CrqQoBvprCUOeKiz8Yx6PlIS8IwxMgs/SOXMMTnHbVKLvOxkjwVF7JzJkG0DzN89jPBx
cjMXwDkiallhDwQKfR1CLWtWiHBNlfmnxadftc7/99J26g6NzY7ZwhpP1FfwBproS7DmEbQe/QDf
xSJDG/9GxUgN2rbvfFDcXgIVVyROzSXLVFwdJ49iVEPQxh943+6OnS68jyC5k/nP45sAyPUPc45m
Cfwx5qbl+zAspNe2b2PZByfcDdElkv3OAYiMD7P2CDPBrHmiGX7C6GXsd/UXf5nqj1qhMuzwwudm
9VJq+K6E8P0RWCG1YqM9S1xi10OXSIRXAHLYXrN/JtVVuQ6V+X19+J35gSudgzzx9ndY5u1Xzz/r
BeyowEeJKH4DPBmkq9qMEf8IQcCF7Nd9SZwbz8b7oaeAoesHDkj9Fd8DV4b4IHPxmtn3otB2aMC+
c+kkflx7eKmBWmI1jCqvx4HMyb3Kcifbrja3L9EAHb08kLY8Uyz735uFXxOQX5gaZRzaRDn70NNx
UZ90zAyv0u9WUdNJkUObZ1Y/nH2hENMJ12rHm6fwjNCRz0tjNoRXgxjamCVagUTAGuc4TEU6rdh3
0mIcjeuEfXPrpnQunZ+s+W1w6muogDuQLd8vwriu31I9y1zQlGzXyXcg5JcBvWpPnL5GGl9bNpBW
1STWq/6Zv25ktDIXIcw+fguvP5BeI6ugxd95YO044dmQUcQDZJofyPJU8XIc0oMygNNhMX0E2wms
oanLl/OVCgYc3RVaii9AJC1ALEk+vDFX+L79mFhFSctLIWEL6UlE8QdRxF4N76E9QDyhfWIKh2Qp
d1u5cykvmrZIbkpgzIKx9XANEQBhCaNk8LfHrsjvuIgkvxnyRgc7/A511eDnWYim06/PRZ5VEEGK
DxHiZsIfEQZN6GIGpPpql9goecCEG7eJHgQuwiRIFlf2si8Sxi8SDQ7EPNO1+8DKK7RAr4Fh/rmR
dzyvNgV4MSJTG02uaCtA2ERXz+yyKqQRzfQEUQpUziaDLGbJrSSnJQHaNHOBkQJlL7nT9rW1noMf
zz2RaQ5hkNoeffQdzAwNMWWFeGbuTFgts5gp+82350SMimeYcEo3rN6l0fmnclNs/SbWP8Khs1YR
pnpctq3xdYHWdqtzZYkRqIuilf+D66wSQmwDP7AZgHRqmPYwzIRyM+dBeGyniFTlK/ZMxt/chCiV
a0btnB+wddk//LK+6hliQYwoE+RYU+hcN/E//fZE6Nrv9iIJ5I1rwOOKTBDuuYz91wrlHRaW2kaT
C3M7aCcoa2IGEKIjqoAgEH0UXnSkwRcYcf9m/r3RQ6K7moFeyokm/Kn1MMO/NCYtW5sRPrKy8UGs
1lbbrd7ZpcpLJi9Af9lNa42rYss7oY/M6hmWf3d3SSyDp3scs/0w2taxvEZCnt7Uy3GIYdhGwXC+
VReRvWE5UooZDbOuL7Y5X01SJR/pICiAnZWvKgvgs1ZKkp+qaNfBf6mGMZqwvP278VN8DiEWg1fi
sGmMeZ7uU0MZcGUrlmUAH/JPN5lIPdg8NEoLlEu2xAFbUPtAZmg938rPVUnFqnLas/i9GPqhSO3/
09H0QDkgAol1U2rYbirTW3+H1wg6XghLwh/25h9TVXbcXQT3aQzZZNx4cKFi/yH5f7vjVeCyNPzE
utbL5WHQQ2D0iiHfxvBd4QFFwWGdeRxRU7IdfDBsrCSQ9H9aWPQqwqzs/CnDEnmB7nBzSoBOXuDR
Z+c1BYabBKIj18mTUpsyVeMNsgcbEMVKJtIo9RgGA77x9t40Iw/5MxVfNm+6Eed5VtwobUqG6+DI
CrNLIQp2rjo869AkuViOH2pQ/DxX/TQ1S1P3q8bS9oKUIyzDkPxvRZ2s9DGXfmMWVXh/LOw75cwQ
PS3KqGbyIcIlEM68RU/eKay5vnPkDVKZzs9p9z+US41GSo2yCF3/7H0c3WXulXEIuyLttoq3TpVj
zGfL1Hvll7nDcr/KufoDe2Uv+pMdu/mAZ+wmTBGWqFvt9TAYsaS3SZWMMJAVB0MxFc+lQqDqzRbq
/1dGWSx52m465RYAaMMBYhJTW7e1L2QK/jkPDkvAsaoRYVqCR2tk2M9cyFdndXkkRStCSvhYwjJU
mRJMAH88DNbHLApud3+TGgpjChroyRy0qa8shT4E1kguqJUEhFxmLP5gSYc1/O6N1l62L/o5lsq9
QGlH6bv1lRPjz6pnryVX1j8rXskGETh7HSdQI03IcVpPPSutnTW6TMuHJWxuIjAtGtcX417O0zD8
QETtCJkQ0W3Ztz73Epi06N/EYovBZAOjJGhRbYC/+i4g0AzEKa5NANWbjxtywsVY3g1zWM6tq0d+
kUoIo53vrMRO3G1dBlp4vMBwhuoEEOZk8eK9GPCN8tMnSP7RBuu0S7Ov4jXVad3BX7+5JeC2PJj9
JnSXUXgfZbhKowVF1c4UQwwSSEuYv051J8y7Hx/1FxHPX1KsaooMlcnErELpT73CUbM6qiy4HcmZ
Fa8GPFxz+N/qhoS9GPqCvuVCuGkO/otTlO8LUfCF543hc6QA4ehReVkhem24A58iDJacqDWkW0D+
fXFCT0TnMxwoMI1HNXTxDFkfGkFWP1RVckS5zs83V1G0fqkCONoKSRx8xBDgGeA4fH+p+ar9zplo
m6wE5aGAGIMCS0lIE271VSkHXDhogh+Gy9mx9dze6iCW0FdFZQaenVVwisyZ2xn+G1X1We90AdE5
wv/rWi6AoAACPsJRUX3BQoMUq977NlBIXyAt0WIeu3Lc9fI/nqlqwfC1VeWoDdEziKc83sXf0BOX
ejq1lxxhpCAxL4UYySIFSG4RqSJOHEoECbqAPr3PSW7B6WoHe3QuetAaowhnojjDgdMMgNDnlQCM
cdUDXp+MVrvDAUJlcSdNDltkEcs8EypKgo6slVfm/WlOewDaav0SJ9HeZbwJ3PSPgihu787vart+
7eWOML5YtUAIKFdcSucbfzLqJJNVRsQC9bB23Ipivj3WFxF/8IunHK8fThHauWXvOM3icPRvQEMs
MlHF0GPEqzHe+1phUEW4xz3MMGDte1UQoUZum5RoWs8waWXejjcwmIleEVVh/jp/mQVWkbZGEgpH
ruQjr7u+Ikgi1zDFUdFHpCZ3vSdiKgEags5opP2W13hZYR74Q1uiPNIDsvbAFWmIiGjSyYcXhIRA
YwziCOREzeQBsNDmI7kLWGh062AuLB3WFYclEuEuksQv8Y59YNBosG/AniI96OFZcrmLIwEiaKt6
ge5kpKlxJ9H/33hyo1FlLaC3DF82i+O5v2OZdsBQ/DD9bOG04m9psvTuFoOn7W8Jo/zsmZN4MvFQ
KnJJjUHTICR4hY2kNe5PF5pbWK7kOK3CKBW3XK8DHwGA6xEEedpZpi1nryRyXzZ6415wEK9ZW7kM
Rna/GCDHxzXzV1LwAsnZNXusTp6vhpotdN0srLFvqClliANV6LNADUCQFsLkNiI5cqjrrfODPN44
55IONQRJHS0ploEWd5+caOLso0LUiDp61pd6lFf5bwVuvyM261FPcNjlD/2/hd+csXOGnBQPbgoD
Q7J97GdY026pD4otKm7JUE5QNn7MBF3uAvcZJdl1V+RVe00FDwQM7kJU2Lyl7HPcxG+jxega2sRN
jR2rEoOT4c2IyvklnvwfVaSM6X0FmGpkixM5plQtz0lr8f97k71Yxfy3NbKelWj5dYjPSCWZ9kEZ
p3BZcSUEScfXDbm1maEGPe38zZirtbpYz8e9s2nBhQ+kW7Kq9AJwJXNFNrFWsi/AMHxYqTj0Y37J
w6NbrUgJ3Ps44kPIwMsmZbmahYplMc0ilX8RPmTTNu5wr3moBSx4RLlG9ryLpDMqxU7iYKsRSeUf
6W8fs8H9pkz7pjZtK5BYof7xwizZwe0fKrfM7KIX+/f3yYjH7Y+gUoLSmvGNR9kbbFbX4qp3M+Jl
W4RrsjOGebjPQerGwmjeZLap6TvYsOUFAqtFJdiFCufycQFivhMyIBi72c2nbfdBbZdDjSN7bofL
abNNSfvVxzQRXsUusjmkp8mzpgW2aeaC5RW7yU75uX2a4fJBfZ+Gy4wdLuyNDmtsKkklK25ztMTS
+o9dNB0+0XIwcjLQRDo2MTJ2YA5Il1H772gsBuRkdD884QGsXuCkq/vYNHmPRPdkGK95De24khSd
JTH0p3YiZ0qbCCoAdHfI4HRZ4RWHhgjs2RSMWD64NcKBsnd8DF/V3nkSaNiMc0mxuOsZjxL9KjAh
bc0OIqI4rE/rQQKGeScdNfhz3nsYxyPegR5BChfQynnAihoXQBJkZFXDPkhau2Rtpb6x9K67k0gJ
89c6wtSfhHShhtolTvyvqua/oEKlmFzhuSqfMAejkZudVmpT3SLkkr2XNa3M92uMfQFMQ/MCGIY8
H+FdAwf+Ic2Kt4dNNuDeRD4SQtgo2J1n1RrWuMhSrA3/1obze78BFUhlZIaalBcRhZ88NGEg48qQ
EZD6Vefxw8J/8M4ZEfAMI+9ABMFkdiUr1pNNs4Ty5GjKz1TuJ0HMW6MOI3JIQ28Fmtp4VmlBsy4K
QPR9D9fJfnD4Z85qtxizkwglCZlkuSaXK7jYvLqPfZABJonHma6W3DrS/lI30e+NGkLmZcn1PZcn
7mmTltSk+ItsNNTs8DnhxwE2Bhxw4klK4bQo4A24P0/QhEES4OqsSJRbhodYOWxJZIwoo/b+WhWQ
st8aolKx4ESipmuVE1ewukqD2Uhi6oIgx8Wdrwko23bY73pE7/8m0gmMEfogUHKqe6IKo1JlkucO
me7ql/bQD54yo0QG9eNRbQsC3lNcrmHc4woL4SH5/LRHFJ+ySmFLWeHfzIazPOKvi3fYOGLiEwOZ
zuAshcLt/1hiy8vAJ8JMu1ju1sQ3K6HTW3z1l3FZ2K6NL85MvbENRFJ8OpjT7acInW+mwV24llXz
e2AndIlTrOxlN4QKUTzjp+EVceCbiEp2IYXkgXrLFV7rCNOK2xYvG9Vgb5LHLmyQn/QMmNxF4V/D
blutvditebP5+5BGtQcwH/72uo7CN3wOYwHSJKCSaf2nsoiQhrolbMgz+AA9AijutoR9f8v3kg0o
7U9VrcgHp/zRaFrX/QxCU9LlzCrQfRjJe4/KrOnUlSTxNqb3cFf4jzWWyHG3IY15OetOALAgjqvu
H/JwJKw2TQ0jL2Q7lvACyy1uWI2pihW/FrkZV+hhyoarwbkVstzPGU0QEQbopGeLjFFY0Mzvm7pn
kwvOeFzyZxSDUPMidbs5zfGyRIVGjZjEuz/RJBYJ5Gfx1K1Oh2w1FKalRRQnJIT57VKQ0eg08l2S
enyyhuXGz6NGtdBzG8BQv4xaE3TG18TZUlYM2DkLws/EiGub0f4PeLLXsIMVIJwNNtAcyqzU60Ka
+uWDiqu9fdarbdSsAA2Kfs3yov7jLJarasMi52FxKhbRsl2XrDVyQTziLbz4FnWk+MWAzNCjfHMV
tcByQm9l6l6/vPNjXQiPH+izuJ+E5PK1/8V89cwNEWKHoqmMfruw0B7NKrD53baTgHxiJIA2vPIv
C1ReNyRzKVBX4ImZeZtTJ5otZ8ZG1pWNKzIlTdxGGdgBCsI/T81dMJl5ubt/WM+hUy5ei9lvx7PQ
1XDdjan92D/NkJmM3dkIFArHHE1arKPqBpcVGQ+0Dt1sUoCDbkj/mlLCEDIWJGGZ42C/OgLjqmDF
UjGEp46yW/S0kbg/n1bel6BZWdnHtDhpV/tinYW07vFI2JHlo7Rk9NG0f2LBHi3aBN0lvo1CYi0Q
ItEanhet8Vupu0TsWSpTQek4vkw2FKmC0sDOB4hFCssa8M0Awn4EWtfOXUWRP4piQ6hlKKRPWH3y
jCxRRTxqRmAm4zi6JbhlgWPOl9cPPUdKR0WOCEqijajTIzLJroG5cAIOwo5zbmCf8Yl9pxPo0zzX
3fmlqiFKYRYDScAFcbgjgd3UfGx06AVOy26i6yPwoHA3pqPWRbUXi2XOQzuo1jeHhpDM9bUj9FE5
Oc4LgcABYLWljW2ff8+DjOmizig3Hu2xIhO5vCx0puyxEB+KsjrZ69kasscSE/qUhyCn/jKhwOaq
ITzaU157lpvL7SP3Hm+XVZ2BUac2K2hMjBFXzRoWjBzXJugvSZxzOAj3Gy0NQ3gFICbuTPRcfRQQ
swsFeEjOICHOvsk6P3dIk91LZSFt0STfb8y14vW06Cmu7BGS/B0Rnw86Xl9hL8YndLk6j9KMTiOD
JACL9MSGfZFZ6iGJS7477FYV9iBfZRalfvw9g2IHTsKTOS+KkgdCksoTm7n2/TqU32Q6sdJMXscM
eApXecDRk5A8alyKhv9eTA+ZtEnbr2Kvfa5rtzEzY0Cjqzjj5CIq1vOhjBgyoUN3QcYx5FUejRan
/qy9/8V0GmloxGew4mH006dOfEbgkFLcCCgIL+M6/i4Dk67DKXsVoqJI9I4V/RKUYafQ6gGE8OKb
eMMrgCOPjgCVHL18+7IBXH7Im/+bwuU8a6EfBYfYjSOe3V7UO6VrvcZlKE1DhRn11OzqKqYSDcuk
kgY3f+8yyTBb+eOvu0lEGfXRk1QguTOg880xXJRAsV9eDLO+TCxySqmeeih01L96bN4C4Den5prG
aEUQWxpKTMeXv2FWwjVkb7w4dSs3ldGHAoO4i+xDgks3MgDoUOwAOx1/RxoMozdkWk3UU+KIM2Lb
z0Vp6sOs8m5ApJwZXJDYPEW9AJI+7rLgnCm1e5G4QPq5Waxv/oowz94CNzQYS/FisXUJCdHxptey
7ZBlKQE3deesLrlT/EjS6g/hak1ZJk6A1vKbYK+Du1+j5Kv87kIhsKM3XJkBnOipDqMiWge0QsjJ
G1AWIfYqtw0zU3fULErQyU/kcTGfTbaFBUUZQC7jlX7B21iZRC8GYQ58Oh1RJeJCuFJXkY+soPP1
JSABtjjnSsSh2hjp/ttAjBhTn87B0Wv8qD38e2iFkKZ88moolfqqTka1OGm0DeVSwMzVOI7M38dk
UETFqodbZn9A/YfgM8iOqZgsIzBUiViDcOKJ9mT9i4WOtVsuHTRo0QgZVHA8vlKtSjN92xWcIhvB
ut4g8plpC1pkcG/cDL/HUlOZF2vV5kO1J2y/yDaMoUE7hcWuS2dEDcX8+dyQDaU+UvKYrnLNTgHs
YqnRW+R2gE0mGU3/qDu26arMxv+aRhp4/9UOZh/Jb1Jd9A9BWExs3he5jiK0wVQPAw3Bv3tmAifb
H1TJuTglDR1UdGGZTtyFR4QDJmCzT903aGq7R/6COXyBz0sfm8k0JHErERPhdusgatqVj3TPNaTi
vJ/8ZKSnqj4XLCf5x5itn3vhAt0ImHuQ/xHlUiDVq4mj8PkXEIRbcdj13CyskxMbvFtghMp3b1S1
z8eHEeCm03++OkQM+Z4FV3JIR1EJ4D523LmLsPsDx0zrD93VG62CCVWPmtryOBVqTmX37EN4C6fp
Uw71QuRWQ18k4Gp644BmCF/Fqv+qSdd+C2rxF/+oVdOpD8Z3GNrVV7VVTVtr5cGMCd9VUfRFUY57
NI3Q0YMkEiqzj7Q6fhDvfRL8J2Fp57dFjO0u21Xp/54RdFqVJUkssnZyFOBySWQPE8HZK25s5/K7
CyT8ZDhrQ65UTiOFUZiJL21KMSRssUVNWz78D+QFSyNGof1u3U9mkBE0ZZVry5ZLpAt4pOmb5Qww
Bz8Xt/Ncdjs50GWgDxitUvQZ9T7C5+eOTczcrQSxWStwuelrl5IVdw2dp0ErC+QYqXcq7rDEL2IM
BxcM7/WDxgfUTuSWkZ8y66+dKYb8Cf28VYwEN0ihdXf6rsloY0Gs/W3gSM8NXE6F/fSEjE5JHN9+
/66FgXlFxev7efCRqtVDzqoHts/k5bkBpsi1o2aGSUNqN6XQa7jNgza/9Xkq2wysv2mK8Sdx6iSn
WtdvCs4KZdwdn8xWq3JGkoiMijM4HXfW8oEEYH+9CiTQ2lztAb4l0ViLCScDYUhJYwDsNGMFBqjx
+Ms6VTTRsQNc4ezON99NI5qXw1s3RIb5h1XvvGpDpiVeOEKWhS7xLv8l28IfEaCYW/vsIcWL89ls
LpwYSRkW5fE1q9+i9hC/gmihKmu4FdQcsc4a6viIabV8jdkzJjmpmm5Wkv1e7hKjk4EnZG77kDVZ
KvboZvr9usA+LIt+qZsKYsDFEvrr3MrHoKqIlh10MSJ6suFST+XI3qpdvWP9u5FcoS5XqMdhr7RC
y9yjkXRKFeE467ib+hAqHVk3sRlI+WDaLNf4du+fBkJD0HBw53+0YX/HUvFq1KH6mH8HhUIClgTf
6iVi4MtFSfoweuzpDR2luVE2M9Jm2MYgJfwH59XyMt1ifoXZDpzt8EHeOODa8sjC+E/OegEcOC7g
CHMiJvuTYyrU0HZrT8bNSCnpgR3jBij+XxRukfvaps/eXcJus9SRP1HfDU0XxZm7Zb9PnyawJWn5
sDZ0XaG26KzHxgdmyQMzvIVvl7bKNg80ErA9YeWuGvzzjEuptw1rfEmNr+jGFZf1dQ7qx+aEniY0
8kcnoPAAv3EGoQpMSyaiazZzCeHBADVcfxGDQcAzoW3OBVAAEeBs9+AlogGHL88oV+/3i5Ux1OwQ
+AIbLnzL/4DONl1GtD/OCG9PjM5gguvm0Cp5MLlEZpE5WyCbk0dN8pw72mfxFqoPMI21f1+vrW3M
uJ2K0ouuf1ZqXdISq6Y7wPZ4llzfCFbSGjz6/cF/eZYB7Ng24yylim/yz2HiGrcxSBvedB8e4Mwt
e6gLBa91TJjBOVmPKbvKX7VvkFv8fVtcnhvzrZZX2UIVsgQK5NHezo8w9sLNJ/svNVb7gl8XoFzo
q89YNodXj+u96aJpiHMwEnz3ZwtPSnSGAuq3dYeJc2Z+ALUu/WyXBp+Rdm//bzspECz7nl7UdLJf
JNpW8GkTylrjIenGdlW0aBH/GJ0jZ385CCvmtEl4yzLD2p/ZtbEL6uxsEcc0qzgKQYspGC/WcpCq
bPnb1HaooxqroyCR7EKXqwozxwFST3qrx2VOKVjCuZPRN8MYL1CnCIzx4U71hm7yQhY7/lO6sUmf
yeQ71ykHEdISYKl4uncqxhIkre1wj3KPt9ONkT+x/ieMfKUVRl/j13Um5+2GZviGwxF92tEkHEmy
NLEDvkkXNTXtgrKkVyo52UBgdhtGK/1w80eznHv043pzgUjw5GcGzf6hDiOb6xvavLTph+PNPTxa
UDdpnC48ZL6031oVU+vk8a5Z2mqoWP1qK9eJxOkArlE36ZTdRooLExByRkLF+m7wNxKbxJ4JlrBj
5ckNhHr7HZhilt5hVOMW5JI+ApQwHAYxKEoYu8Kb26Qpu+U0TekZHaLks0pp5AhQcf7nmYkvYctX
ac8Ptgt6XFEaPDzXiT1OF5PsX/11WXqmMb5JKttSAEDH6R71bkV21unMtFmTC/tMLVPY8bsMhRdj
2Q1d4GwbwyS1sJQ1cGc+g/MBb7d80YVsMGLT5iO2tQpq34e4mQACGq+NkfXO4h2APED0rmq8U6/k
TQlN3eoAzeQ06ELut74jGtfrZldDGknXx9xiqrnQwuv4HSs7WSCprPmEbYpJAwfv8BCwIm7CoSb6
UaPJUY5n2lfFxjgIEzuseQkJUN2Lfm6o4Kcd+jR1Pw8hoMF6/gOe+NxBX6LuCLaqCmWVUNO/Kvcd
wlNu8as+E4uRZSRnIjRfbEXk6KSSrLcurqYAdr/zEWC0z1K8zKpK2r46lbslXZ0GHq55HmhU8JV3
hr3GSnQMvhNu5zqGuwa12qizWc0pPR4OzF3Qg0Uuhyrds+lovtZfDO3AB58ZmNo6gVdKH9zgvgK7
ey/oWKnhEeHOibXAoKO704Ve5EiiOLAIzZtp1TB8F2ReDhPrzq6vpw556rcnXn6DIfSR9AKU3Na/
8MuXaXCDib01mYWhkJ7ePNCB2nn7R041smADJpTKGhhV0Y4hZ4KnHUFunKCfxDG6IwonJkvrdje9
QqylUxN/TEFProZ7VF7WYQITEj+4RWZb+7cRAZu6JC/uktl8PM3C/J9op53cemBmgs4q6dlLhhWY
HKd1JLCErg+ee/7kAn0BEhyR3QNAK5DKHp8h0ukqYpYJIBOIpVCmHe45mrJmTl+aCMX9hNEeq9x6
Qy7gY5K1VIQgMo/32CugqAEDHg/9jkKZn/ZKUfOfj6CC7eLiIJzKvxrScz30sqAOxr4V4LUjBroV
G1vfdqHQR054ZHehPtM5As3SA89YlWGEhgGQyBkzh4aL8mg0jErQuzbQm+lkev99lCkrka4de7jp
NVVXTj0QYCNEXzk4v+8F292ZMV7pNKnlGwpGMuviyadvgONGxyknwdtmnB72PDSUpHM3qNys5E9h
Wyj3ySE2qSvLQ848cVvoiH9Fl4CSnSXHsx9ksj90JbSb1shrxrca4OIM3wb5gzmBmlIxXzZSSAXF
rgkVtk/bb5n9t8IIMJyV41lgd+FXyagafWrAQlcKYE4OJkWBEY4C946S6Rkd4syMCM3KHpe0Qstl
ztDesj/RieGVO+VYnHkzYzFRCl92SdbbQHFpLxoQpIxQyox9r+btGSNqperXDKVkWs9HTvmdqRkb
hx4QFUyVIoXHAwNoJBFi2hTXqqX8Nh8enJge3UJWh7Ep/LexDcxf30LZgigKfbv0xmTfSLyjVhnS
PM0K2s18Q39b1UxR9kDbMWQlWDEjPZl9Mcwwf7ic5N1jRdwwj+gAP3cRbSSAedZWoP8npGfsUNMK
6CqQq1VpqXUSL2ykdPHyY6aX4DJUgoXlSQw0L481iP7P4dfqCwnY6fk+ta7SLr/GuCTWul4TDw6s
CFQm9W0fHp6mGPfTIzUt/JI98WQ/7SwOgxy7Wb+gjknfO1GQwOc7PFe5bbEjk9nn6S6Hx+tZwqef
XNEpDAfSw8rslEPLFKpcBIQVmoJnmESQrzIoWPtUoW0DwpwwLI6/R9wSLQcOz6KwcWtXF76sXrNe
Q7r5JgbfnbmxOxAZouT8C2xXElKVZbVrCEJRinCqkzUoO7mD/yCtA4Y8UM80MEPECAwViiUD18qN
WPC5kLVaM7b4uXkKhbNszTIFcfOzHutkO8RHQacA2HMf6k0l693VIyZUoCUQyrP1XDWPHGLx7Av8
tT6mgZ6HfF/1sXbirCExWrxRtxO1z+lMB0iKVtWdy3WGWjB5sEckPsj3P8nNvc7ij2Nr6o3ycuHQ
Jk4F+3YJ7osVAUpFY7IkaCPR1W+Kgal+T5b4luFfHhepTbTlMuYTMcNJDZQqsVe5k8y12a9NIoaP
qBF+tYEaGHGYy6JDvHotlbLzfnpZMoOkgCVPhgRbgPNTyTY0pRoiofE+hg1OcV8cxHxDb6n1Lh9W
mxC86INEwAsUpCs0ydU79tpXqiqXRlnZe6Cc2tYPtjOlqMHH79eY2f3FZoWEIxR6I44AT5kymErf
rqQk2pvxd6+N0HtnrCD19gfIMbRVH7qHMM6iCwwHRF9D1D+gLgTJ6ToJ8yZjxw8rjQpm/VazYEWQ
bGPDtZFxrrfFaMXaW46+qtPZ5xWQrr+yCMdXqm9AYmZX80lezKki+1URw/vBBWCyBTyXIo4X7TEs
MNcuHHEq8VIPZouSUEaMysly2B9ofP+r8pq7Ah3CTvFMc99BpjAvFUqloVLNpycF1BZOO4bN0H8F
qJnoNcAjJAqT9o5X6iidQ9qkO8ezjgRzr2pzd+A/sO2FAdw5OICpxm+ND1pPMmlbG3IJO75hbqMO
SWLxrP6WYWzmdqcwu1stfd/lae3l0pmnYqCuqeWLS73IHjMiRD8MJGbcAMBRTKTcki+X6oNrkUNA
882LpqRfu4zSe5ck6UWOpRvh+Ywa/inutUI08ejiYsbFBLR6t0BphQDMgn2KG7YMbaaZthRzf9TB
1y4KskWWeptWexRc9Zfo8jlw+X64pRWVNPoM8Ea+lxe9pfe7lWgSsgGPz5tDkwmKeymmhPm4C0XF
1Ja1yc0FIqHW8RV48HDarFThN8AC4NfnQ8ToR8LwVG8KRypiU3kv7O8WMhWMAO3p4Vzsv6QYx7c+
mcGvp6jQEbI+E3huV1bWYygeLkIDsb5qeYJwwtRNczZUzo6Fn2N5V6W6Jq7+wwLQD7RThLJYavhD
r0g+8dOdiAM7suDMcGxx6D/2gHA7xzl7NSi39i0rAeVAsuKQ+/aK/zXoEsckXN3PJ/bEvasox6T1
fQ0tDhbAVz0Hoik50HOK1ZUWdnTVup6I3BJLO4DppSXvCgTonqN75WknmJs3PPjuuicSSgf9vWTF
oxjf98Cr0hmTg1lqN3pCPSWS778tapRa2wlFnHyPxMCIWZovLkXwhCfKTzaKZfKtRuAaribH/k4r
v6gD6Ikslw0eA7YVEfPDM0P4f6D0m4rrrdr94kXHRU1coYnMHRlwjr6xxLAH89Q0IDe26VT4TVKi
XPhHLF6ORwoDqbMZ5ED9xqCLVCMHXtFmmxpQQT4xWpA0UDfECXIS+QxHvQmrOUd1KwOFXaMVvOcZ
xzPWqQfbstaiEKncw2oxc9Kmx9ZnlGrqJumUM8b6rnwGbhqA89bOHysLGbvwR4qTs7+av9eBM3ke
tMO1dpVzFT43ftO5jNMCmlm9Tj2/hm0U240OKE8Ggia7hPywxaP4M6tBkyNatbzRHQFxU4Axdd6d
oRe8r7JixuuSkaDc6741qHz/RK+N0GpxJny2KPtLoErYhB5zqLU+JtbbyKbskIcxvykJ6ddrdNna
6QACJNRZQix01KiDsSa8Kos4QHX2GOMm5L/wG99y6/EXACPeulSk3XCF7HtRpg9xwlBNokiID6dk
k697VdcEJuwI0c4aa5MQ+DSidktv8E79t0gsYasMZRj1dUXj90w3HZGXwdEFX94h2DHHYtE5UCRd
Vip7B8A0bkUnzf0Ld+RfZxAeqZVDsXpIGRmCRC3b9khdWe1yy+OT5Zug5yzFGzVF0cP41My77sqU
08Nujqkk/6LyuXBwORFobOPiesdRto+98O+MsqyamaWPvhEYngIWXkGxxmdUKDKD+7zxrMVlzWRW
i3gdtuEUGfDo7mFJikZmI2DEuaTYL5N+jd8j1x0jiY2DzqPkuzCMPZmiK8r1BWvbdwdVIGE3fvV/
uT9U1kNVxAcaNdnie5GMuZ6nwKXwOaKZIS70+Cw1ERz3jXVlIsbwBYNPvjLSs4En31fBVNhmJ1eA
uFsXgrg9LKYZOXKrbfM41U6bfmFGNGAvzVMwo+bedsuzkNnswTkYFSQ1ILEO/EFBkmzpspUztjja
JlzorUCdWQGYTpB/Y0+GxfZNuHCGR5TFr/gw5UMazQrb0LJphEJbryFT4UZ4Qjij+kpEfG57bc49
qwdMZUw1WdDYIYOQ4q44z3gK0HqcoRNyANTq1UNiS0d6P1wjt7POPl1n3r0kkxSGg5itPgr52ob2
MwIsQF5aylHeL2FnLixa5MmOB0IBKTyP4jJOwARmNNqbdaX3rv5eFXR5/UhD/Ih9fFcAui22JYK4
xMeZoZ1W1cDzmqwke+bkKwcVCtObG5bFGevgxZtsLPdHSQ5MfubktH+la2+nNP7hBccNf1px5cZp
eURAE2e9hWV5sqP/yfccxdO/O/VN1aBaXvo1dtk5Jfc1eth9jYQBU0eLbnBQ9sNKykXHo8Qzibe7
oQ4oEWGrTQ4c/ARH+5VNZ/iMUKeQP/Vsw3G1yT0deqK3/MNicda/SNiGDuxi3X0GqT2d11ez9gdN
GPkXqoAh9k1Kk5C1OFjUUoV1yBJhgv7SBL4s3X8lwY3CHZ2HAqIhQhWgrlYsZTCkmDMmr9xkqHbu
1HksIQdNMLDN5xsvsEYN1APA4mEbDMcSdoF3xYPf85HhzUkGbUetRAYvtHzkw6xPl3x447mnOCdS
BwQ+hufLY3zvEXd5jTY0IQfCR6wdF+AOBCxyyJoMukuzRdpXEL4SueR3+xQgUrqGWVKzlu8XhBwt
8By+q9jOjGGPyo9UNgjm/UAeEuSr4aqI51jKX69kY4pvGJRBAdVowFD52I8/mboUihv7uapUvtAK
Tc09pJzb0U5bQzVt46JqEZV/k5cyFFytdoLTgL0bZbz8zSqr+F28u/+RbJTlZObenCRfmHfHLnHJ
fcKMVBg9PSinEWcziAnOHpk0WthM1I4six0CmCLtAVXQJ7f17LEpvuhjNqRqGOxR3evvP0qw13AW
ZZE7WKUEuJtZEg+uUIcbVS6hN7cmWKpUV+YX2wQhyU3kPb/oWdEiKUV3QqSGERTnTSsLvy1bSi8+
ZUCHiJ9shUOg8V71VTRXTe0njLeyB7fyLgcyClA9LcJKlaLvseW6/oPpUde4cb+pDneJWkXSe4wX
wLgE0mlqZwKvIp2hRHjmIDCPsIUGo4mm0I/cSi7P96qAsQh17i2vsqCYL6IMjbULaHOgmARDIKMD
5Rps76rVFj/j+WtfIftGgpF/il2RKiqhw5Iz6hlmU1GfYQCb8haQ04EUv0WWu1WQax+vRGG4HSe5
uiOmO+iaQ6MsDOBdScIMOFibL7dKMGm92n/zmsH+Q7oIOyhX4561pHM/SfmkwDx8REhYOkEF0HC/
ahKb8zBDBH3pUqVKIE/dpqD7e18gRG/Giw1yz1Xb5nHevMGzMnibLV2egkOe3XAg0jZihm3ZnQSs
f52RjNQqpBWFNoC8xH8+Li6Lyot7Dd64d2bGer7K3H2BajRGoMgMNcw6M/imqnki2M9e/Q+unxYn
nCyxVM2AFJ7ICOQKgOZ2R8ZuoZMKnvfyuI9s179t9HgvfaDP5A1Jy0ym8yspRU70Ci3dq+K3vphV
I7lhD8ww2Dwp8TtyUFUIIX8ck2cStRa3CL9TvEskIVAoWM0kG+jumj5adrpjXMUCNcz7BH4p27pF
B5zXPHYeWoPt4LZdlPoAmMP8Q0Ax9YVz6VjTkVMTQH+8HhzcJI/3EdqUZo+LX/9rPhLeb+ZSKbcj
5tyYjBkn163YPhBqjhtSPdpUOH9jk52HsLaJN+W2bC531w0AF3IAy7Wdoddk5kQrNP0fpiJfFzmG
koaUuJH6Z5XWKCgXjPaSKfH96W7vCWw/LqOxNYv5781f6l79dF7Z8MrCNglM631VdCrY6d1E6Qhi
15WIfqtdaMNss/v42NZZc+7Q6l1H0rzwRq58rW138Df3alSqYkmE6YuSUMNqe2ZyMDQ7WY0rQCm1
JcBCWKkoRChbCGDwUmx9VfgEAu+2MMG0m1l/hbTKGXpc5mUhTc7oC7fIqI0CE2x3TH9EhnWlBgGF
4UGBoFSpLnjSkIZFzhih4lPq5ZHZxLAn8Z/pjoqqQjfYK8VA2FLqV8akulLBa7HcVhUP9cRrFFdP
/zeGC3tuIPITomJczXuR7HyLExM6Y4aNe3WiVD+kM+Kx5i1DcGeCxK2fCY7ruCDOmV0gn44lDWRu
gxlawtzUouVUmmBvmB+n3pZvvitKpwVnOMc7ag4681mgnrDj7T/8jbm2zOrB/MSy70VdUrrg3+Sq
Agsg8bKhh3eHohwJ8tlWZKTfniqwcoXhntTOhmv/iggTMl3dp9Aqx3/GxQpmNPVVU8cY6XGonthC
0f5TJfQE5g3YtPcDg4tR5ZbEK5PtygqcG7aDnqljQfwx2DM7BHPKP6rS6ske3g6BjUBL0wwrmuvw
LdDUF1DotkwYoQt18VV5PZHZ2Gpt2kUtBxoSP1HEenkrhP9Ijf5zlbc5yYRZevcF3h0TevCH9pbz
lesetyhU9Li9Fpm2K+Jq1PNs1854gXbLeBciBy9xzS8GZzqqtgZe4ARY5YPzMX58LAeHwfadSAOS
T0UGgtsIEO2ymxeq76nVUcRMlVjj44QCLI+nz0d6sT5h2xcieRrEAuwiZpnvQpsvJWA4e69pOLqX
gguHvuBsw+cdWugIEAEL3fj9wqI+KXNb/0fHTYN3tv0uL+IOzAwcAAyM1aj4SO+FIMKs3ejqc+9J
XX/MAkhPHTGBqXWr08Bbygpkzg9jd6Q6BJTr25JRtq70m0wBu6eJQrzLjrIRu/62zLLsrXirIapf
zUUnLo7mKoo14y9vrS4crD8fJWEcCHLmL6lRRjteqUDK/pQav6/KYAIIZdfD2w23d0bBhQAhw1/m
mJwBQscw0z5i/n0q7HumbHs4UKr0b1sY1tI7Is+uFMVQGPOBtCyad5zoSpgcMf0NgOIO32o30bRk
csrsz7jluPplShMqljBK1CubhM1eOyiwJbuk6BEP9j8g6L82XT+wLPop5WrBApD/KO7FvpAyIXCP
QTbgpwG1igFXLNA4cJBt6eyqbikY3nJ7A+/LdVZwuIsNddoF40eZBKe7Z6BfWflqdpXn05zvaV4H
88ur2cqbV1seaDXE+tUcLInYsd7V/xfcq2lOBs1dQsqqMGzjyotKaiIqpX5JP5Z/6xDvHjOZnpm/
zv/0d5yULCIe2JBAIyuH1pa1y7naLcCpJnWGcgdOiJbR8DLxNYvQ3HqSESTX3ij6yHIOKMiP9Fuy
BIsPkRdwoikX31dlD0r/wZU/C132WDDBhjpA3UlO5mp00WPRXn/eCyB+sFplfr60tf3D6eUojUgJ
zxgJ1PZeAXPM7zhYBOJWBq6k/3D00oS2YJBdM9l5IQghFZFkmxTh9YtqE4KHMlAgVCp/NW8Co05h
AhtkFtdo2X7gYXNHc7dPoH13Y9GNKxLMXmAisX1hBo5C8eZ61HwlAn2ygqG2f9Stozwlw3F33qrU
PtMJ+S/eZRbwpnQ1Qy6OM7bxDmMghY9wSNLd1X2d5qMkSTVYJegE3OcAt38EqdsQ18kNiNDPow6S
plvQP4akk1H0rCChoDphktKAkYqpypYE/q/n2yTDUsPyQIFgkEWbLzbysoIsmYiuTgrp6UA2SWVK
7lwGolkOpjcExK/Y0It71f5P7D9784hn8aLVIJmnWZODSJ1EL5dlOPNgiGUM4t6LpMeOC5yB325h
+x1t5WDhOdF5j8mjFxcpOD6Vi3juaKjbBLErd89XmGM7sbNXIQ1N7VHoAaCrEG23e9jISulwfixg
mB38jymLqjGF/payvmST6frM9Zv21LPcz2uiD8QamuJS7ih8fM4EVyGyvX0yQwuFtDesc1s8F+yn
Wya/lAQtv0nqQkmqVzcfHxBqC7TbmGlwCWcQqZ5VmdIx+6HWwORv4JXJZlekJFnnfPZ7QZnPRHao
98q+DjCZHoKFM5/QN+neHS990iMbuL0MfkrXEkOa2juYHKpV8cP8W990Orm23TaPl3J1EykBkPzd
j95Tvnnfk/UV3obWjVDgrA07XwzWjPWbLQNvLUZ+qA7CZCkWlmzNYkQwiySubMMNWsspOq4yl1ba
nMZP+4xTR0Dl5BqrQ4WU1BJv+BkZYOsQdk5x3hQapxxqo6tNeFmeAUDmkGg+laCIeAdrb/Pn5Ogr
E639JBtjn6MrGBg0y/3RNUUXG6eD1FgdHtFA0CUf/J1j3dxBXEquECN61e21EyGtWcKRgQSGfptl
R+FuYtwV2ZRwvF7AShTcYdK5chMdbS/wRrApBZAyYDYdZLYVZSb4xJmBdHTI754EoKUprZAkASIB
m1j3lTOHqyzyM76HeArO5gBqCybaf+62FslvEt4AD3Z6tCkGieWx2Mkd/bUEDq1f+nMiORncGeEn
SM0cqtfQ0uGwDFevYutMXDLu3y0vuJwmPRTr/H1TVUzwVCOPRDFVRgw28jZewq6wxm/jX4NpdtJO
uQ1hSnj9ioJFQ66vcvZ1LX3+Rj3lKjZieVsehfras8+HVIzouzYU58zZyS8axaeIkbajaP6TZX0l
Qtdd/GZEQrn5lmJJUcj4VGxrj1540BAplrLXXltof6LEDS8KOtMwZCFoxf6mlA9kf2GsCIc8BDMQ
17fwUEAf9AL2cQcgLamt6whQizrZX50jDktLesykzQMoQYcJiulg9O1nvVf6yWEccpUtKVeG5L6c
zspBgKc/2yr7VdcMBD+v8Vnzf4nWnNTLczYyhqVUQyHxcd9QEwXyr8h6wHg7I4xdw7EOVoaQiRD1
PdvKqgCoyXIRfqCF2YyWMAv1K2lPU1JUHufTpGKlquM+VKA5R1BX4b8EIFl5bmIvTEczWfChi1XR
5b7oNlESH4/pZnSyUvvNPoMFSGnnMC64zYWy3x0PbuBsK5Ss3eIW7TT2onvO22vW25j7s/ai5jAh
zedxCVm69PxDSttkk7YS20Zl07C8TwkaiHw6ada5eT/Zz4iRR1howH65UxXe+VcSKyvUFadTqsGx
KBLF9HH4yeEVJT9Bbb+KE39O62WECxSF1GMOfxYcem+4pdjvODh5Tv+HYPUTquQIpjCGXlKYfLvx
FyRpdBWFEvWMzPepnl8OvOcPheR3AgAZGD8IfS8BXjkiUKlUroMMZZ+SAtMMzFSTF16murgAB8Wo
EG35Xoe/G6Ls/mOzD1RIfSwCAZaE9erbazYq63ik1EcyEN1nBWJEhMVnb4iepGyXT58uLeZMPDLV
i6dZI9879QcrOvPQ/rwaptIZs6pfc+3a9kcf1bvw5Z2qa6DEUOjiG4v0HryQSxiaiWyU6DVOiUkN
xHcNbrgvGTfjAv2GU3QWR5Ub03H5ft9dFnf4nKE8zJOqgwmycgqBLsCxW1rylb3hXEK3tqfQpFiP
BdS3ORP2RBH8U//FjnCOlYG4x3DchquTBgNglCt1VXdNZegcaCdhyZX1uor4BvoA0IyS1B0AwnCW
nb+GW+srqeYpZ/AzplU4ZI9Yl/ccGPxyzOMttrVn5vCKG1yiyAEB/4A29VTQMowJWxesymRAcppy
yx8fUkGphUCuwImkDyNI93fB6iamZq/oMMDxAiLWTlMH3peJBdzsEdDTdgIwSSqWVJYRZjf/mJLR
ygpeUgBZGMuC2IqOEeO/4D2fNzHEAI2M3xkfYxLeHTeHWyadcF1VG/JSpKZ8/us1xSnQY6rY+ECM
v036HoVMQmSNlB3fOEB5PdExGqb/lAte10WbpA8gk+OMBFX38h65X4QYfritS8e1YgF3V6hTIypH
6IFvd33XtJbVEHhyu4QTF8O6/YQTbwMS4ypy6L/569GzNx3DJfcE3R3y9qPg9ragG8MsrNUnz8BU
SNzgVzE83PWbTyhLiOzaPFs6jaOBNivFwwgd6+MUW8edjhNpn9bBRWZH3buPi6zAoT92jTryF0bH
/hgpVKUXmSqyEoAOVXOMH1zmIWmXy/0NdCjIEfH9Xe3Ct5m1+MDECSubmtBpR/1GtAPUgr8x0b82
yoEaY6etCtbyb+cOUPnHJ67fYQOmLvxdF3viqGkRwwPeTnX5XDwMmBSZ3niEiS4oBM09lLTI7CAu
Sj5ZiLt3ZZFD0DzzOI9XKc72/m7VqAe3V31CLarmtxKDX6pYSEjR2zj/J68dXNJjtawUaO+8VauL
OItY3xklOB0uCtdbh2+I38aWdx6uqHMjKT8BuKDg6Ri7ZYgC4Cb9anJf9dblaB3PPOAyvKjuZgny
jRuiLPM1jAlk4L4F4H1rt3orFcXG/osimLBt3gQeUuuF8YlTbaA3R8bzagin5tPmG7yW4C7ENbN5
CCmYFzxvZtRwB79tTrsqaDeJfRTNqgzFmF1TFLB4V3EOoPHbwxw7MokPnLnUs78sQlFfWZc43XII
Rr2Psd/WYu3Yugj0d9/Z2NTAdfOL58tqFwV6S1EEEw78D6r4tSYl/8N+gah/jhSpUln1EifxJr16
Ven3gQhLy9HqdVp34ybRhQqpt1dv6NHUqbs7B7Mw6z0YWljNCsvYBnv398i2lz8UYIkJUEubZvak
hBMbUCyrKl0GOKk2/gz8VjhEHcY/HMrbfUZzpVSZd1hOr7EdGWIupf1wEOd3c625wRqW2sxWwiMr
sRI9TyEvURLnJOgn0XGrMotgKoDOVhhrZH23B7i9GUOgc0+ts3STa963ku1LKtsxiN0izTVgPjQF
YVLjuf0+EQv5BrryC0U7CCISjpS3TDZXQTIVNWdjdHGkgEjrUS7ooiAVwpQp4eQeptsabspT4F9e
fucKTGlvtlB26w+jVJD2R/mtT8hv+EsExftU4iF4SJUDF7fQq4ui9Ym/7ZFjR0ytDw4AZnV85e5R
10PBmHjZ0b5M3Hy5nm9g1rDLhuGBIkb0Kz2rG3RBbnbt2KoZEHE2tWFaYrc225AbggtkOcwDoSSI
kubeR5YhfZA4RfKr6B6Ew+mw1sDFwxPRc7gO3HNc9oT6QtjxXwFgEjR+RfuSiujyF4y15nUcvYnM
k6SE34iNgaro7RxEB0WFBFW4W1KnxY9ajT0SG/Bz1p2jmDj4z4CorvaQMj+qBwEQpsQPRMdthJex
w+Pe0Kvp4moIxOoL+ORCLumthSB8QbzOQsCRABIxpVO6b0xqmyV/o4qkW8xtR3bfLVmSAu8b6BZd
XgnNMvtiq+iKuxpVG65yln6LjKTdOIqESDTPRlzBHZPIArdV0WhlGkavM5jg48FQx9pTZ+spWdWv
eswEi1IwsMUrsbZSs5ZWp3ljjxgX8XliH4VWbh4xNX4XCor7hpP4ACdDvbQDxfGDEHOaVRSm34sx
nmrcDc74w0U8hXLec/pg7cB8HJjfO8qTtk4uZIrK3QD65efsLFEQ2WXIglOnX0j07bFQadLyeI+v
TlPkUHk6RB9G5Vad5K6UxYX4AqTRNo9Di0fMjpRYZcJ08uLMjgVBHzQ5Cv4sAegeim6wethSP4R3
nV8XEUC07psfNsLN7TB5q7UAVLQlivpCafAha1l4y6ruu4VmuD6oeLEaE9h5J5YWj1PzyiK+kdJn
p2qMVemwYm66+n7qcbniJFHH5JuXU6JlWKPGi/d8Q41DKgvJuxUnmpliuf+tLAvBASZfMVAmElQl
ZVKJvVF5hTsf3Wpyxq/jvkVX0k+JbTKggdUsBfeR4LqWKacM8qCJ4A6wjwZ/TLwTEz21pbmx8AcJ
URsJewjf0p4VQyuspcNPU0yqXUKbXS8Cye4HbLVeeiV51p3xvz8ltRiN/libczKqMQ3YEkTgFKpx
RGMonABx5gTxqdcU6kWhg6/5HhP4vnuESKsKn1LEckoNwQnQIcHb3NioAaXJPb/+1VCUryQXFULx
VdBVCPN2THAl8xhiio6Tlhx4lR/HAElX4Qr9l6EVNmoFjSAEQTaMmenf7ZaJ4VVkGpBgsMvMxgPs
nHlfV+XMkUdRPfvy8ASjm5YJrcmCU0lRC4dDsPf669fkxIHsQliIK4Oa8XuTSU+Sn6qi1yNNXqVf
qVedK74sGrXNxd2TTz+tHPw52005twzmLpbQGbC1fToi3qwkFXL+yVnHFPAANZ6r716ZBYIbNlUW
qUzasFxCn8nS7WHn44g7Q/ex3SLQvMcdMbFDuXKc++UaN9kzt6kNCxcnF678JzjaLCIw3Q+JcvhN
af758ASKpjVX7KoK4vspxN3tVmsTsWTGAIRdDGaqBPMiS8uWmG4zUurcMfwgVx1tuoX+7ikrszEi
VoOVr7qAPq/hHIDglOn3UL1+0fboCIHOe059n9zM520h71jul51QBs+AAEu3rou5/yn87a1sfsSp
ykwgmsoHvAO3qUTCzCdOL31Y8EZFhRCgeaF+wnm/xDcOemkOtMOJqIYqA+D4rWiNyDB3h9GVT6LU
+fPpK/wny/yqsS5Tp8l/h4eeQMcX8s3HszzsnUSLr6aOPoStjNuaK4KecKsZMZ3C4VDJi4T6c56X
pfyVTEpcWaTGUM4A8VBYsU7S687ZFNz9Nu8onLh+NFKlwqjOplBintGJgf/YijXFPC0qBKFa8NeW
Y5CjtaU4AYZkwVaU7k4TkoRIiM/9C1UiKu6DNgtEbau8Jo2n+fD+rvzithu55JHmfgA+6kPpYCOJ
e/6+DntDk1EumPRn0SpH2TmmhqmEHGChsLzGGHY3FL+S5weql7Bkewc6WTafO8zYeORXms+mEs2l
4kVOdVGtyl3ikij4z4GwXnMLd6/uru9lxceVjdONNh8ywXMleYfLq4xJW30iuvEHYfCTXSrHEegX
e6oa+sT5Ke0+qfsudQIL8MuAGDJYYifrQa0I2CpzKaEWiNM5OS1noW3IXCAJ54vjho7TAirUE9H8
qTMi1q1cBqJsNkq+ddhk6p7jgbEEmp6jLvX8A1etpyc7tZcyne1fBFEF8IwgiHe3vr9R6iWn7g5u
0hNJiAsHKR+juz2Jz2Tp+CFHlo2NO7M6QDVsU5IGtU2y6p7G676fzHeVTQ843UTpas/2GzJCQ+fr
+NIrv99bIyfxXVODa3MySPBg9qWlxXlLwzInPWv29tkkIcnfElHMj6DHDTSipYqV/HnMphsPyBzK
QOhRfI8yja4O6QKEqRLmiwRic6ClM3z1OardhAZZqd8eVoqUlxpPus3MjMKbBUYx2Xf1wZYr7IZV
o9wqVnveKyg2K2lS0FOUv/yY7BTuR+RfrO2ItYrtZTvivwQKkF8l+Clmzm7tpZbuWIq7sgsdC69c
zeGtSMpsyxHlaizJ6aoTNUw/gf/uW9rUTgirIJZRQPUMWpTgxSHyrwuH75rlEHJxdYhK7wFUvzVk
IKZ79OX1nNvoVEdXXrGIOqp7jGdl9Zq/HXqROJ1gos8sFUVZKeFKPE9idHsfYqXVWNPUH/IYY7Uy
DRzsqcgSuHmzZCmLNzvRuC37SFN4VCD5x4hi15t+QVRulZvmtfgHHSbvIGFDMYA4Amh/nHwhJMaM
LrnE7aOyZEfcxJoVaZxID+B/AcWhWaRf2dYmJEZG+YqIFYcITw4eZpgweU24Mz0vpxCP/FeDUjpu
2ZGj1id2WCFheS10j+qSFcLILhOWyaQlOiiQ3vjFaYDxg07b7kBiZh+jsEBjPolpE5Qs0nKjFRul
EJCx57gNpXTY9BvbBbXdmvNnNTSRuCS3bQaD/5qq0n93m6nB/ImBlUx16VfdQME05UtolCngs/Oo
k0oG4OmKfuwkCoKh0B0CAToysub6c7gCCzwtDrC+yHRnxfCa17qxh3LS3LfjfEltNEB04cEqyxEB
EHWr/sjhjdoKtyYgbErnW3O4GwuP35vN4spEfe6NYNfjlLIfDJaRId4lp7OZFYB6g2xPl5eWEomW
ORmq+UFClpAyh+/RRvr90uE+xlNmmn56BiJlDNKFMVOdHjYFkNIdvkYaWK4/lYA9xgD72veDK0Fc
ePUM5RalTKtBOHrtxiH/CGBwsdtn+crj0az+J6ZjDSwSN9N3pf1fnzNhyvl+KVNtFQasw09ZVg+m
bf+ffhL/GpY7E+zUx1G+8DRMCC3SLnz4+0JuqjgsoepqFv6XaoVGbDSvb65fBzjyubMDHd6WxqSZ
J5sMI9y0l+Q165xI8y7g5eLFhB0rzdaw2LO7gFIEUl4a+bvtePsuE+CJw3UHQDXLIHhwcC70aZIk
zW7O6zKDF6YZkZrcyrOTqU+mrR7LONJLdBtebyFsSPGY81wGmKflCesBvnA6bS1jxy+57JvRobe8
pzimIqeRTfbKta8ngVDcBVWMku2UOwT15mTPnoeDWJH72Jwp6ZY/wYcYALK9mMJCkVxlkjJHhu2b
yoOzRqjy9Oo02mIGDdyTtlBK3hQxTuLVDSWsFGe7H0B1j8e6CaYkdAbIWJUhipgd1V6KnU9LpBiW
554QEvSaOkYKOhRJgJ1pDXvlS8zWamgtYLof9WRgqrXqGjKrAKhOdrCOG2RuuUlblkGlfg0FNIns
xHm3sx/P0YWddHDJj4qN0uLpGtsuV3nhgTg8d66gjmjtFN3sSCr6JyXR2KtxGtvAkG9KhqxDHDxE
XgM6c5ydwtDf9wJpasWj68agA7Eg+NeaDkJ7HJZrJKjHwMOg0C5hqmLija3iS8tyO/Kh2qeJCl/5
d3lkzu7mbptlNcbn5ldlVkbiwnr3tax5YFoySTQqcOb+EBHE09nLUZI3dNSoPfOjI09GzChLQqZg
7EbJQ9z+Zk4FJLgH3k4Wp6XqmzGTk8qeJoBkEY1cdWceQE60UWqrlVrHJSCaTgv4oEzOJK2DY+Si
xosTIykFDTsVHoVOkIF0zABJ5RQJ19UXGFAKGXlXziths3PtBfX8uiHyBgFPfXpKky/CKr4w649l
76TKLQaaInjzo6ghIjXiC9a0MYIE5L+0KgfBTmVOPNxR5KJpJwNoExdEDIUwLgNmGs80cEwns8y8
GzmT9dEC5uhfhb3chk+wsaCHuqO2Al+Xf31cM3MA9HVtuNr0cowgMNoMZOxMqpEF1H23t4WwAfas
Kj+HiwAWHRlSdjbpzBg0NA9pEUluaKrDe1p3j68OdHfMKrNCjeuFqKgHi2s1UiWNJx+4C2VYnQf9
LVZGMzJy/lvsENhDpU2SZL1ER1IbiVirl//zJCxligQGCJYJjqU8H3LjdW0sA6GkEAkVSJjc3TeP
2rPaWc2CoEOXG7XJ3rc4eG+QoCkCuYoNjLePVuRyG7pohIQJJeWQHYSpsQ3/reeX7mF/OTsmNGBE
+KUbbEWXeubjkXYzaONqFbbOXeQtZWy/miEEqotaS6KiWsIc36WUnAupO+VFauaUlkfV3dUrNMUk
kAW7dbnNHSCIsVkM5BRSl0DAWuHiC3Plyn8OOkgpMVi1eXeuiu/JdyX5bYlQv0YEMXdxj75CImuj
OjVNUPO113kj6cMo5/HCWTpHgQAck6Jcqz0BTA+pFMdR9xl6nAk/MDQHFT4kPj1NltMYQIloolO4
FngO+a7wZpDmWfPWVcKsXwGvHn75nam+P1lou5cS/JDeAl12t6eLtBXyY4bOPxGfVygkL0cegh6v
EKqsg5rRGSi+CyunpIC1wpiSiUxiY0OgtH6HMaKqi50beiDE3H+iOSFJ5x+JVoaIcb2F1ZQiuEX7
lDMXeCDJy6uruqk5bEgA8Bf4UcQhaOjALRqHQSvnDBHWp8/rOge9PPbvTsdZRc/+nYouiLCOh5Dn
j4sjLgidVrrm/gjMNcEypO+vCF/aJpi1WBf7JEtmsiPSuIVibUCFgFoQek3FvHLsAX5z/IueZTjF
A3ID3Ef6Ky1R48f03a0POrEp6TkgMXRwNrotIfkJbK0cgolBDgrqlhSsKjVBp5rvWdu5NZw6y19y
i4aeow5RGtxRb1W4Z6FwSX/70ixbhnu5VAXCUCxTutttzpWj53XtKn2fkCslgHv4iD5MqM9W3cgz
lb+ZZuDUfqnMlzDLT4brN3A/dwLgxwXEiJN5rdtUcmFXbf3Y/NfD2IYzKljXqClzl8kGT52Q9pKO
3mt7eMbmYakHZkIjjofOCa234dstQaMtprieE192AfknsTWDftYny+TDK6xYSGeP6ikDBoaSNRnb
uhyBJp+eQjNVuaseCZ/0Q7j1vx1DC2/MqfbsaIpM+Qs2WxTFSmFRKHWgzU29hKSRzAHXTZuhYI8B
PCabAbgMICy/uBvMaUNJbxR3LdJ2iawFf5mECLB98K7XA98yky67zgsWNUmdAMMRbHuwsaaO32HC
hjdbTjbgeW/BcMTZTwCCXPNS5nb5TVQF8+YjFaio4i1tE6NEe2pUJwVSKRO3qxiIJgjabUAWAtYw
Sbqbm8G6zhoaaDxmR5XBWu8kjpz5R1FZOxZggdu7ksV+5tEEZM8GeHQtpkN3VtCjzACmbAzbNLxo
HnJ31jnxnw1FR/yJWnUlq3RCBVlF0jdzuL2kRWkpC3aq7AXbLNPaonYcgDfvodDwZ/IU6Xut93kC
anMZ2RJ+gZjDJsc+inR3EK7KQt6unQiKRF26LZ3wT20TmcCdTaCKqruWEjVm1KvwS5nsGzJ+5CGZ
TvdTlBPiFiycznghTujfXOYkK8fgSZEzJgUM46g1ci6sp2EKiZBEUdHdOGWICN8ySjab+YLeHfOu
sxD/90xbVWaORtiVtpKCrOaMBS6iWvH1pGKDwdus97AB8mYSGGvHIUeQxbf9mec+4bH9NOeCtwTY
eVWr1eHh4SHFC/t0EnubBGD2FadO2nvQ0ew39xg8bq809zVcMyM+O0sUyYZ8TeI8oBG/08hXz/Jn
67mM1VqKsvlq+QhgS+wgIFlEU1/gjZ9iu7vmrlTUVse/NSGYwOlY5K8EHrciPQL4djMXi2PcWrcp
qaVmQ6wL4Ou5nFKXoS6lmt1eDouTbaIPrQJ6DFpkyUdtzuAH8kISN2Dh2R9bTIHSfa3lTvKgcMZq
0cKybDz2us5RpMxE6tpA78ueDs4M9nym3sl7zXEVlw1RuwvrI5gilUquh3IBUHQqZcyLEPA4WoJl
BNIsw+Vliz475t0ibk8e0KvG7fLhAJ8V4OY1ZrW+9lujBBX0/WflNEetUP4v57GEhcCSg4Ute51H
kYNrA+CNpG0fhX5C6s9xndt/wlAxKBX/jg898na9ojzqDpeLf3vuPj8hTCpkKIrGF2AIeWuiFchF
4giOyM0vyMOdKiSDAz5MhQ8MeeGVvrz0S2+vTuaoJMZHJshPFQ70F1J2vw9OeBgLPQCkJG82zQmS
cQfnH34D37ca6GqIxTVGFZcFPpVLX3GQZ5IXlfDcLJCZy3dok0955i7p2Pl/wXNf/IMFRSte1iOb
q53Mft8RecCNZbaDP3RGJbWZpoapoARCIu0+31WfIhWvesCrwaPzuVo5kDVxPB9yog0qAz/k/5fV
9oNq2Fw3a1lb9BA54EdsJTiq9Ndvt+3TwUZydIshX3YTUQMgL1/w8wFQzOQ+KPWyeB989bNffHGZ
9/qiCeqhL5nOmS6RtUd9i6DW1YJD3u+/m/U8zQ/UInVO30RQKbsxiPZ/WRT+GGkKI9S02RB2iX/F
r1PuASsmTpbLaK5Ym3dodmc+wtZ/5oqiVpkXlNwM2wl9Mmvfb8m7UhiJSYJr3CBHjDkQey9GsI0q
DOZBfXRroxUu0hr5xVf9VAAaODTYte1E/+lcMdTCzP2hRibTttbFIdNXh9QKljsqgy+jBDC8T/eb
fldIWNrha37Gmluhmf+ZpMDkHMWaMlXC9PyESV9fcRkKlrgI9JpgxGq+O6rkomHTZacuEpejKr0t
j3Lb54OLZltkSlKcycJukIhzdSUyVG7pdJYh9dtccFs31pYY6JkGORlhD3qtHMJaYo/MNEH1TvcU
qfPhSEbiJynQwyWDEMvEjt2OR9jEw1VezJM9vfck6zRja0Nt7+drzLcAMygkrQzQTbXa2EJjHJEI
HXOUzAuhlIzCRI1D+lj4GnluKTKwrsoOy4K2CiFaoiAqT/Y163DuOZAFK916aGETMC4c8wlkrTzg
2TT5Ma3h1cUNio+70CoLBnYahthoSd6d/usnQrTrb1Q6H5si0iNoP45+NHVsZoWIduXDZztDd3gr
eBQD4C9K6tR00EF1dfilCMmkpDP9tt/2EwBPVY5ZkdOeUdCr6ntFoMev3doDQ0VWGs+l+h0b8oXX
VCsX/NeHI5ujnOjiR2IPN38WD+gveyNAuX1EZ1d/NqdDMxchvhik74TRJ/U2zA6VQNZpZZrLRS8y
pyBk2vL+GCAOtCRiXPukjLkoDvdxlPQSChaZ2f6UEF5E9qsF9HoNN2BR6xg6cWRzPysSkhOEEbFR
DHmrHxSs76IOHqE37XPPeyC/mEMvAp6rKw9XVoy9VOarSJlsKy6knMD6ph6lUDTA74jfPSa95mkV
YXXrJD9Pk/tXwivzOo3+/kewobVKGjMV6WHlgt1hkh2DgM84N2dyFUPOasWGXxechJ7qxkSH63bA
pfMgCXjocuMb5HaehNq7YJCLjctQKZoGzuJUS8GDNXWL/qLi1Z4v3trBXjoWdEX8Bp8ap/eoP/Xt
LjFhweQ4SunJxpg0jM7Kc6z566aswOQ9vMu8OQ+RLXv5fasy/QWkkkPU8NlsjW+Vns/YxERrst+s
HuAVetixuBOaLpA5dQkAfTj7qpK3g2rCO1zjZCYWL1xSh1975XuyEWJi8F55+s2iLeIRtGDRqX6Q
gEk48RYPHqBG1wEOlTVRGnlYjVygUn5ufdoqT/LaFDtwt+DZfT7AGA416Clw/5ppMTkoo7tU4mG4
lrLXiGiSRPY63Z7BmXh/As7YNJb5TUhIzSYXPUQBXo/SbGMXZ4z6tnyAZshn+Ej4BamjnOpSM+TX
eIrB41I8+IQ9hwEbnBbs45ojpYdvEmmWF/G7d+LT/myx7FE5eGzv846Z7lMosWxOqKDYnXTI3nhk
oVLpqL+yzHFvyw4vPbJ5Cgd9o8B/gnB9U01SApljVuFOuStuv0KHTuP/K2kudz1jJiov++xTw0/+
N+gg1D4gFhmKlSMZGMddRS5TnruYqcVdTftaW6DjBYm5CA/gPDmuJWdQAGxuReX9ceHJN4hWRNN/
2noqmuMTXcI4TE3iEseM5K7zw9nzEFPu0tnXq7VLct7b9NxyfrRRFPF207FufmNK0WfCqrkF1ekV
OIE1UfZusTBBKKLmt4vGMIdCl2ZrFjF9gpFm6Ws/nFVcWt80habjh11l8UBDPWnyBmsdiRzbrIjo
8OfE1OCjqc/VWSVyN8LUnmsrWRyshxSo7Vr2kVhTWPMvawPEjPEuUiZdQ71cToN+CqdhW0LMx27D
dNzQb6eouYW+jzhMeRwddCWqcbVNL+9c1aI5+M9RMtQa/1pKz/Zk9OcarqDafavXjF+JIHMgWZj/
vTt1imzdtx5XYfxrDUHhOaGIaoqk7OLyxNXY+Rmtyu2128PQVX31g1t1M1atN81meifRyW5dY8l2
x8FMUdrkptTVNs6FMJmqhi/hD1VdvBdPwWGFQ05wRYT1fxLES43IOYkrfdesL83xx1nVusQTAgbS
1HJ+VwmSKic/IuyYRCwM2vVLSjIEBjefpgKE3K0j7cN/v3wL+RNmBkAueF8JycFzDw7QUyK+TRL9
pyJ5ckQM7kampF00E9cyrjUBNXNQD2wLF2zxZu886LWTY0DqntKDFzKe7JqOQ/T224VSH/en+xQo
Fefj72QFJhogu+xBBtjwCJqodSObKzW1LfufQkHXrUJn2JWuRI1EkDhcdNqVk8n7pZm9BxF7p2Jf
ovzJDe+JbiiXKmP91zVA+8X+kAlb0gcG6EWkSELe9IX7zs1+yV5jsa4sruWu8ZFIxw17G/4+DmGO
RnnUNL5g2RU0+aJJ9OcuL9oN+sZK9PT8euhqK/xC5f0gU1EHHKA2Ka8z5nF6+5BtP7qbulXuth8m
kkUPYtdnlYmBEZnVofbcZQmgDx0abTYBGw1eTfCys5ehGtm7jZrqaJi3dcuC+cCHZkcWKTulrTTe
zarhw2/NVXt4wbI0C0172qZsaLc1QV0Op+Df5PG0E692gO8Uos4Jo+OvwIpkGzUfuPuzAnWzzVph
ORxRtKrqIDemTw3wDqbbQXyDdr3YfmOOOS52g2nx7tKxmj8HG1UJRj7dnfbS99UjmxOJMQW1NuVk
kSocjnoL8pSFdopgXDl23NJE5lL6Vsu2o5jpQHfONq4uu+lWe4jQ/trs7OpxGSVmeLM+Cfr9Pfhy
aGmANSe3fXLFT53VwAkEBHH9zZHUdO6Y6yGlWFLrWsUDJWIOUW74ZzhcsAdm+x0ZyjcNTb5ptEfY
SymbnWlrQYUqvANypFsiFrbgrSekMoUztMgvCGVlZ2trsNqgF4nw6tH+ZhVh0vBVhjS8FjlPooHR
1qESSnkfqTh8mJiUchW/gjK86gRWEsvkEEonZTbWx17A2/mYYq3xXPIiOqYzze+NT+A3N+zvHQH+
e1VlE9cSbDbBeGI4HcU/YGCOdROQTn9v/f2KOSfLfBSfKhX95qVkerTo5u5OyhtnM3B1blhMwOn8
E3X8iOi2agPkr1W87zf2oE2OV2/gDHVBn7AxHRAjkmiwev/tAC/d3DXmi0Fvqn5HiW5rCeBox27r
l4FqH+xYEYRhu7xA9zsAfWSqgMtt4/7/oZ8coLk0LmmQcORr4vMsZtgY1OmmsD3cMd4+ycYeaRB9
h4R5aPyPAIWqgavkErCGjBJ4KASfkNhw0YjqOJFcsqpg0lpATIhPYapDVIos9rV6Y/ccBDr3Xydm
3u7ooTe7D4/ssqrLTZIgnMVRsnhT9rrFO0t03kCyBUnwD1MIRVn443phl4K9D01QQHouSSaG/4ud
ArjYzyT90F/xfOCsyKa9YNsqxovYGHDwUSalnmTdMRSKyaUyb+2PtGTHW+8ctYsv+aStcxVQr5v4
68s9hNaq8ROVBPmaIglxty6XJIiXVya0Vrup4nXNKfJJTNq4fVCg1NAVOR1J8CcW7f8K2RTWkVTF
4Hpxfd+eHu06bbrp48p0ALMgXHfvHbCLmIXJZ8RQWAQm2xOPRWVH1fmCzL8FaXfcJ+VPdosg8nQL
/kpm/wNrkXmHV2iypesko5ozuoEA9mNyLqqV9K21yiXFI/QLZwllIFpx9v+PcmiM+BjxFeZ6eK96
PF3MLFUYutvxTlwfUtxH+K/Gqov5b8qViIGNVFeMy7ocew3gT6u95V1wEjBDyx7QAIgXedq6EZh+
V2LuKDEBf+2RyCdIafY1JseotdckRHYgjm+B+2djg5cVHAd6aNJhcbYbKvySPQ39BbsSpUYAmEyN
US3/B/AilhPqrSCU5+g4x09IEwjlTI4GKiGzrVQdSIobfAms8kORg5Q/PgxyVXl/IhuyiMR7TZDH
2rnkNDD6QTgXdkEcFPCAZlafT/Z08XgkEuw0fNX9mezdwFK8/3cEBwdosL3tiWLkpQjhW3X/717t
loS363Q5nWGTqSRb8+k6t7EipXlaBniKaH035dRxvY1cctIryXgM4HwHbuJs1mi92MzpEQVp6JUZ
6pfdxYxl8C8nkuqmdmhlooo9HUdPtt4JnPzKTJ489kVATCIrJLwbHxtUFRHUfw94Svy7DOFHgdf6
FGsAnPXXKQieN5CmGmtmKTIDEfeLzKmFyPXPMP4D7k64cfaOtEUtclCzWaSuUCw+y550zFiMv2l/
XOPiF3ldADF83WnO7m8anmuD6+agoC7CUz8/Pig7DsT46YEMM6+PFtDqnSedHlkw/o5q7+1ynwF+
kJmV4l89PyHXuwhPSKQS0j7nmyFJiXZf/+QpuU5uwzCowHKwxZ7aEzd6Qpgq9AQ5l8e0jLgIzJ3x
+Kqw/pwX2p40QfQMLEJnQARQbsWNjXhS5oCJ45ZALvDTl6N01/RV4NO71ep78MYuh99L89WL3cip
NGQIhgD8joK/+pVMePk4FPXJS96A1BYYx3ksJGEa3f06h90mhRl4CpGIots73NXJQCWwHmlh6xb+
QXOi3BNEnomkmh91Zg8Fj593q2NUA3kwl2mYeB2LbsElpmnoPBEp7BQlcVVbljLKrfZp+Uu17AdA
BUMKiSE9dlyD9I6BQgubv/++icVmOHUKq2H49QEen1GhwfPfuwyXsuxpI5QL3RcBeRonljKufwpv
NHE1bbyybEn4QXfAxE3XyDh3OxEhR5DpKLDQ6l6YSWaZY5wDofJ0a/q2e8ah8n4jfGHnjab9EFxo
MnjaiGCgCPhPcwy3GSNmxYbuubC/YYuVUfhnDsTH3hguUXOj4THBIJgST4wauAqHJ3UxxpwMSyME
5IfawoY+h6QYLaXwJ86GkxIQoxRCZ/ZFFCHm6QWmKBfc81rBZrUd1z8ISmLlwBl1GxjTDPdsCAdz
70izUKscam2fSg/8lxPrGfEiY/WktU/e4jiEFIXxldu5im3WmI94skolaYsESIx0j4GCNhHspp3r
9h+TzFXQ7PlIZb3m4j4vCUy7a5iO9UDN82noaMMgxTUSV4qWc+Yxl0YEi3jd3JytrB6KVqQ8+3pi
rPWtWsBpqL9tWmYgJNek+1QUGb9HYadoe1SH1DhYShBYthvxwGNtl8c2MJhX0Hjcw47ZBivgxWWw
oIogiPL6oVI2GYRMOZKdXZxJZg356GXQVIOzTKXWJ6vUmCUV+42RB84COyb1HS+8e7wC9KxgXhgP
qlnW+Ij5iXbCIqhHNtLMdBClIZCivhuUZIzunEZv6XbTCk3lwxRWl15Om3Ok3pNjRgUzo9iehj/c
q4C5flvGCYtsOtxAEc8xTRF8cK3JghR+CwzNmdxH91+NB4Qp+XsL3xnCGFcFjvxGPm+Vu51bobcK
osgurlqlx5XDWU55UpiZkbx2Ekf1ySi+SNqFBByVeuHSvMy1vOjT42Ez4P4x+wl5j+TzxWgRL9Qm
3rXynj9sX26X+VR4c6eZ0j89NYdafZpUOp2j71x8nw18sKd7WGA5tGfTDjPs/d9RDJNufZUDWayl
VSoGI96kPwbiuaCkMF7SaqpwaN47UiQ62On5rWetHOHDX2bgtvChmtME+5ztFnFi4t8l0SiuCr2b
HzILsadtpwTwMfkr/dwqzbCZhvCods9/6Q8xWK1hR9aJHgcyeBUYWUp6L3HWwSfOyGDnnIPa3bfo
vswsHk4IXSFv0v3y/RGFd7IdibfxXu7MxmB37eW80zdpNkAbI7LJp6Wb25XVxmeBNKaZHceB7ru6
/6Sl/Nvyauw3H7zvAVueBB7+Mz95dvkD2HfpMGyML9ppC2CC2udOZckhO2Ihk1opbbplZ0KUXl5B
fBmAV2jLkdIYvK3ze02GdeiqxJkrdjiT2HHO+4lTfDUxYZvMxWIzS7wgbfvxdvAYi6YAusSQ38yU
KhLZNMQFxJzcvga75DFOQca+3X8+XONqwbFVPLB0gCukwrzAIrKkkTbhU6kQ3lz4VrOBpHmZ2kZl
eccnYvlXBL0U2cD2EP27roDPcfe7wXe0dRXtBwQYCjJIRHlp1eSKRgvk6FuH8cbrq7JilcQFDwYe
IDFZgXtiP9s2s3qVivmQ6ei6EBKpsNXFGwrDIB9+ljvXld0igG/vsp1nzR3cftfyV4Hi9G90lYTx
Gnaz9SJjS3F+7mAue6ZbF9HCLuUkjZ0kEF+eGlHuI+ySA0EyUzi3PBVDpFXTDZ+ABoQOG4XXT/3h
2VFRiAkO5nmMhdH1rzUgQ7ncxZjppDKQm3CV/7873nv6PxTvlJG94ZjG/EuOHFA9gMEDKabz6C34
xMGjZ7KmSHD7oPBeS36LSjUjXDjyTeIh8CyxKLZLsta6GsRHaD8jzvs5S1Tpto6ortCFR/pmVnY+
7qtoVnW4U3kxbVz6xsOHwcSgkjO4yR9ZXAVL+6safuGQpk/THQwgtRQHi+fxagWzVsy1tyG+FqQy
cu/eYhA2vyK3+Z+8CIFl+ctHkyTcJoDwFyDEfJUURZ6CoWLDqrnCWmYiXrB+9/KyzhkxaWX4utHu
w/4fWHVHBuvWMoizzIjrPP9AtSkcSnfbKzE0Iu0xn5KvK2k1v15uFwUzSdzvULhonqju1Tew7qye
kntLJj3nR6WgIeYEI4+I9ADg9qLMMq4q15wKtH0YALSZU7LsWt2zshO7ia8uRlLjVeFln0x6pyWG
Jz7gsdKDLXiueEzPcOrEdeI4PPqH7tEoDFuBICiGp3hHc49EkItNj1RMcNuIHfRJPoMp7TjTaVgp
EAtbK3YmiIZEWi/cNoGpIuqQbwr2LHq+W8BBT2n+qHyu2y06tlaAVDfoKSEEx+kXrkLjJDN8yY/x
2rrg+ugC97rtBtrucVjNN5mbh3+jw1YHUucnDM/80lhiOaqhGbVLE9fNz6Mnz6SAoawKIlF0jWns
qTdlzwGDyOOxUrCVE4nr/rMmcpr4WZ75olgLxjUstEAYvjiMwbzbbRsogqEHb9dcJEiesqn5b57K
q4AYkCH2MZYWgo6yNqrlQtjnl20FBJZfQOmfUKYmtxs745NgiuJwHkLEsKCxnpgL6S/ja3m5gFZA
FpFQaQSTD2R2qs240QNn71soxz8iGEwushDC6eJ+qL7qc8+6b3ytjkCotbYl4exHUnvh1EJJ39Pp
itw9PRZpAv6F5w+V0jA7B0z8rBzymFaKW7t7e4e0/gdI58LljZP+62ylUZ1CVvlypJ5OGgqv2tEe
SmnYnx5EpZsmBgu40jNVc+6Xn3pHt6/hu0bJuhwr2PTFxVhVQBVODLl+jb1wgeBIywxp8d3oG0oR
/lgsM9QXB0amUvAzoKLqlnQFe1CFevXx4o1xMoUOvp2U45FaSolsJNssdm3qNOZTdPyYUz7QXlSQ
c5jjZ4lS4bk2VG7OT2LoYSAHgAbglkdHAvUNGNLZ+8yOYYAKVNwvE9gSab5kxOWNQfodW94Ty6gM
sAtot+eLqKH5igOQlwucLocB4PalXvEjqVBMfWjMsdRd80QESPL70s4Yymdjql+wu0kmt2QI9lsG
4t7Y/prZLnHijszv7auxwMt29RZyflLBKxUyumWRAiIASeoQi9RkEhwiismyVHxxiRVIM4/pDwwD
22gkBDE2BhrPP8VYgo9ildsikXlKzrD2LFbLugCccH3qCNZhh5463o2QV1VecLeQs0ZbwJnYt4cy
8q0J34KSz/3y/PGrH9j1z7HyhyI7WyaEN/3rLazv0qIfph51X+EzAgNz9XPzy2k+YnKdyu1hnkag
Hr2opntOgDTsEwrRDQclw/n6qznqGsa/8O51lYF2lkcdomszhIq+RZVpuFJQO9I3qoLJDtHZ2pAG
UWUCRXERhdv6pr5xRstsmAlmkhLMOQ1Ydsj7mSjuavr02Tr7H/Qt6P/Kbebf0smzkJsjaCT5Sdjh
uLBwN646fajcizEJwy4c8Y0nO9VQ8XpxeIhxHGjcVfj3NIoBTJdU8lbx7iwjT/JPNP1kOfnvIK/R
lp37vMqFIN6E+Jcd1xZu9GRmh49d5q6YHnXFuy3FNLwry/I7Zok9jB75ainwsSvwk07H6nNhznAK
Axf/9UWxDxZE+8GvHOKFNFIfwq93kY7/k+X9UpOqDADvvbRwXM5pA1ehMURqgTIh7mAro2Ki/xuW
xlK02qJkK7G4pOk1AnznJqo1BUFlIaEuDXUbUgBuiAR6TdDNAupQrXUxrzupb6AbOk6uRb0phhJQ
0OFHSbXpdpqL8OkbNRJsydpOPnALuRSBPMa+NKDdy0siUOgnPylqyEt2sM1vMrsx+zfepYS3sR72
5+sh6UK0CVDGYOS/vZWA5H9X06gvnUivU6o6CK+lK3WwzwCKj4VmdbVe2ZSS7PFvMqMgkDFnQImw
1LhDpa03UU8KbEQPLk73cJPcipgE/jvXe7crvqaJ7jiDNDdaj2xaghSeCKew++ZmFzWps1yUwo6D
XoALYYa0LDUgjpa+Eme+1LRt5WwxCq6bjYcnbCbkat42AVUJD4yfrQEfixr4rdyK6YzmUOIJA9Ln
cONFYo+R0+ku6/RJ7tOkthOXOpDuARabzYYIEMUUfoqcXPEbnRJAShgl1HL2EXLPMl61nj8ASZPf
GBp/0IOMXd9qJGjw5iHFoLNgapAGeBWHHaifQAFAX/Wi++A3kI6GLlayeHeM1erk/n6KuQPVCY4F
OdEQNT5GbOYVp9Q/+4xxx8n2kpiV+zVjFs42Pkgsq+K9I/VPmTKo614W40Zatp6/OdOpK4UA0KnX
xtvyVrUAMpVPGWdSRGLArSA6NGeTvBUb8/PUJIMYZ0ARlmWMjeW+vUjTQYOLiPiKohTC9Ql1iNE9
Y2UIFfgPAA6B1Ws0j/5DOpmyCTR6QkEmkbRP4ZWVjIdZZ80R5gzRUdG5kt9+xb0+4NPNUtGnJZIL
2ehofapi7kKiBcWPNpRCUiS3lUGbgmtbenkoXcUnVryrGkIltzAtEKlfP9riSg/mvPKcnAN7w+wN
Za0iZzyoONFFPmES2bjF+EUtPI78V9O2Og/Py/VwHfRfD//95eDQGOOBzKG5J8KP6AlJuW5WMbDA
xADcb1ueAQc+n5PErOD6dbfA3zziks+SNHvfOwWT5nx32NadEjGYq9e1TPdhU0t86VdMSaGYcBPf
7Dx42ELuG2ymksDv+JZgwoXtEsW36aul0dJdolxfYMm86YNRx/DSdBEOFYWbQs/0n6tOZTLeBpno
w79zOyD7gAsYPpyXCR17NnylbWC8V0ZydxYGGZakTnDrtcDtotJLujGC0hmqG9kKRJuyH9XzNBlU
b3R0fjz4hYB4jQck3eXhs4cnalUEJ1U2SRCnPohw1HzUDrDb4BJOMHujmcv3sdFp6WPM8kbWxLJI
n4wtY/Ez472/uFFfsR/YAk1/2HdW0w/pDMmcQPR4xwdG5E4Cc2/SXIiNk9GgGjwjnW+n4hQDw4X7
zHb/APpuIzvIjFGr9k+LwcDWp0/mrvzex4bRVG3JNE8633nv6tHdd0+CitV2Jnd5SyXfpSt+O3sX
oq5XeDjLeRcCCcWgSchaCoKErslgOIVmwZSt1LKiCRlg/L+GPJrtvPZfmu5e395pv+QqJPiTj1wg
gvzoJ4C2yytL/aFPQ/XOHbzPf8U4FSMpgjBwOFd5/NX+vN053/1dqRtAkYkyjqOZzbWddc3/ViZx
SCECYivNQZ2GPMBPe1MCIGybvhNPiLVdBmNG2XI2VkFP0L6Ppdu14pwLsRhjmb8DcCaSQoMPErHN
0BH1QT1/a6H2rfKxi0TqUtIMuFEMg61lxXrQ1qQu5uRXzkFzD46KsyruNlHSGcaoW/flph796X9W
311r6CezUzprEJco7zXJK7mMqzZpYhS8uQ63vtqcEybBe/DOLfIcxMdzNFba+VjXdaOPRkcyiJKb
ZYShInsXZB4Ab0gLt114zrzqFKZNs1+h8ZfgAvEgIkV6cW/XoDnto5RSe8VEfAnr9R9G7V6hh3e+
O4pA3dmprutJK5A6cqyG7L1hH9Zb75yzPwjea2Z/9JuDpmo+nNUbCuOMCtlJinlHzKt8sjkkhU0I
aND2ffQ1o2/I9i8oWuf4ZO+u9AoSJRqa/A/vrkqqaYO6HxSK+qRlhTtxWtEHU1NiSDyCs8Q+O4bj
mCA9q2b3u0YCXvOlg5IZwpekXDUjYSVl60zubfCWb8IU8x2XZ8c40rs9AqRFnJFg9nuV2Xlza+wW
PzT5eAwM4c+CDXDjMd8xOKskFVGtchYV+Kzec9Au7NlVpURZvGnF2Zn4ulVVCGjIIHBPSlzxIxLG
RF9GGtwX20k3iq39/9CUX+erTXNqMENV6PqBPx6h855QO7qckoriQWGeipcHqsdzXF4a6IBhMBqS
piLm5pqYi0XBj6r90rxuhN+HoMZ0D64OdNx4dz+hzEMP6HNEVuGg2o/jRRQHnijTqMbk2c2ZinCs
m+31lHWbTZMfH7SthxEcO+/vHcxqY2fssf7ERzJEspF+joHDxbYTqPGAQjSChYyttj+SoEZOW5Iu
b4erXlZiU/RoFUXzRYtZ6ddyWginmV6VK3WiHNU5s5Owwh3c76B7i6MEEUAbM+7kwy/PbPz2mT4o
mDSzDAEuingEHGfUthcK3zxxgw4vKhx2E8h6X5A9dpe+sg29TGO3dcYSs5AntKwpmY+BdHJ50Sz6
j6SjshISaMgRiUaCXsVB87bd/QQVjJX7oNblYYT+z5jTxtGYOgoiD9WvlelZXnPRoQvyLx2Jw/XP
+Fyz7Nq/bJh/xOxVWLlOopfo97QdB+pnkPxrFXp9yFnR77qDZhJHgxJNqKeP+Cn3XuzJZxXCJ/Ca
Povf7nuLIyPWXeza+LtpZ2nIuTUEX6OMs876y9nrsN8dWOLTAbIrabm3qSbHgiC56rsiIk1g3vb+
WzDfFH4pvkQIcMDprj81rSdNo2MhGmigImzpHAiex0g7fcXNSPVJT1N+9s4Fvb3jpOvPo9CoQ4mp
+4smwV/UGNO29iN+Z5qKMTsdQqN6ad2jCSDKWT8w0Q9ZffS1wW7digYoMf2RzxswnRGBVER5YrIQ
4AGTVK9DsuOLK3jUmHFx0sglP24JLzemAcU8CI23gClXiaKJufkIWOuHesVwODmIjKtPGzYeuFHw
faaZa5gfTMZfmKg3uQ4YptFx0fy484ro0eMQEq6R3kGbmYwh4ZRzmrfhwS1rHbbV75FsrYsRMvEk
zpzIcHSIGQAwc2CqNR0rujRSFy6p/iCr52youCRjWP7/fQy7dOb4u8ycefKUTe2OunXbR+j3yyPg
W6VXCSSc1ME7q+GUPUzSmn1wOLmopuI95qfrz1ez5HFlLy1/Lep5lX+ajA0Q6jKg3PSxd73X0NIS
/KNk6V9Hqn7/FkSIfgRN2BrcGjsozgL7R8gXjPdArstcEuR2cF1fHOWYmMvdJbPdQu1kKupKDwds
P8eAoTXCnidDVx5NhDmqnE9mCOXCGiBNE5fHXzNB2kscoAl36H+cBmGL3uGQCZmu4thuZRfbToK3
Ja/LERoKNG3uMsS0lrXTik8ulONm2uFrbPPJF4T+XnsrzujwZvfGsKfX724KwlOXd1uKB9FtNQaP
aX/gc9E2Q2yKgSF2ulkOWdKQSTgZN7CE5K3Twmq0mKPvtK1we8fX0qFee4hlu1AlDAESk501EXpU
Egy2o/sounHvUSdgPPWPI/c6Op/AyvBvac8zt301EyqxZEAZ0leJzh97UQzy3qLu4ddI9wEF7O4F
L7Hg7kzHCb99WSGjGgXzN8x8VmLVwl18w8vv0rSEhOC92c2wJXXAo1EO7ghFLGLoPKXMw7exGSkR
e7D+yppWOAwqrLOed8r+OwV+X1W08MQwvjVnc4WFh+1ny+8sSgzyYU7hVNTC9i4FYs9VVboCuOme
SsEoTTpmGfQcVnerezbDRyN/OC8xSqAeMFGxTzw2s38d2d4ragaTp7simG7S43Ar0Duq79NhczwO
wrrsUSVtV3k2r4/qbscgljZR0UZME50g8TK0hhFpetccTbHWuIAzjoXzvgYz5JZF0IaKPqnJFbE5
A+iyZtkLdfVgi7OthdEhF1aFNXFeA7dJtDmxxrukFfEPyXjQFi0TEeUieKWRTBbyjejdiuFUVVvv
Vbrr245V1NHS6G4RzeRwVvXDZSSGsVZILq9fHCC2gDTyrbiICOWbVSKea5hEDl60mxQLAzA4yikF
/TO0VPG1t2iTIpRTawBbPGpJksrTORyP89Y+A+4DGQRGVcIH/Yup+a9ZCAXf0zMTngUvb1+ye0yX
toKFliBRVMYKPW+j5m1iue6hjxPiVW/52QSR9oISNErP0Ir1qC1ZpJyvVAA3cOCVmZPxDr6kFO8V
+/yqDm2nP2p13vCwnyCsgu/aP+zFAqibPx/GPmqQhzS95h1A3ewl7Q0285z9FUD3SNKKDPdyI+Vq
eBw51+LY6qYIIhFF7HqakWrmk8zw48Fohzzi19ijc9EGs14sm4IXhK3jc+qvZn79KeZeKxMPF55n
bqteBZXlZVKc5/3o/9Q2ZpSpzlnk/PoQbWCZE/CtkvWzHurjDnvc/HHNTnwIsw7LqLg26y0h56bp
A0Rz6WzPes4ONz5Ue5QqpNCH4pjrAAtLWd1vsSiEzT70xKc3M/QUR6DkxewOnVwVI2A3f1n/OvDM
ilV9CXvAmuti+CIDvSXENfHoP8jAbzDQAyienn4fg5HFytRZLQFbQsjxk6RsK90w9txn8LjnRWwJ
AeG7cnX+Ua4DinkzB1t+ZiKnMG/xsdCvPSJrVFvCB9R7eQw6Gb0KFOi5SDpwgnkPVWDZ8D3pLzBi
epftcuYzjGcaKNItsVonFNNzBQLKnYxO9sis8OKCuSMOjab/xU3Akj/uFRG8jcZdTJ6DQGk/mCQ7
H3P5dx4Fe/NAF3OwsNrBmWD+rv6PH2zeZBr1FPGi8bV/Byt59adKYDs9AQoCK1VVUaAp+QcPwEza
ADqE7HfYj/DuVH7bujnkBHjaJGpft0HTiGWVNIy9ku/hgz3KH4aibT6lrM84tYNQYA1nDuH2/Wk2
ECYZlCrHx7k5mPP9aR2md9bPz/meNrhlkamHdnJZXzo5VERebEAImI4yIMBFmzZL6EL2vXBLHZ61
HTzkxWOI6ccnTPRnkplwipaYmgzJs71wKsF2rPEN9Lt5bJDnwYipL/uHjcZY/vzzUJnIjxhC2978
5Epxhp/NH++w2Dc9j0ozYnZB4z+nIxLC9cmMk+2CFV8oNXLxHsYkxMQoigG97TF0EMR24IFZIEFq
t0ikwHeWjHKXmK14NfMNDmWef9yjbEQ8W4H2Ofi8iQWYBRECqFGdUHfI4HP9+Bew0tBsoQTiidir
de1FGI/2bj2ZA5xd0WzxJb0vLc5KFAjB5rG5XvDQYSo0eKxOtHc9NHPoX0nYoYrDy1AnxxZGNOFm
Xq1v5ypP52lgvCpljOC9g0pOp6FhANuOFE9G/Sdv7luYQ7hyyamTszBd9wtgLkd7Pten5KCf+o2J
4luR2Mpl6TzzcnbHdtQjTTzAIWei23MWSVoKglxIoG0gLavtDELqiksFUC/+XFA17/a8XeVJDuWP
DWJTQHjh84KQV33ufIMoop2Eol3bS2f1yk37/cuo2UABd2BTAyEiwmFI7ZfQwss4PGsIKhtQZObZ
q8SmnwEb74NZ37mwM1zCd32oaz6LwFNf9K0SyOyDg8BiRtsILS1L1tgDJ7Fn2UE079o/HRqbG1Pe
oKalkCrAtBkAuti+yflRGCJlse8ty8c0rRiW8rGOc9z9683yEFbHF/Usnb7bEtOLvFfWI5DGWnVe
1WA2NHgC7CKuZCyUwJjNFaxu9rIs2L0RhTrYIB1OHaOevruRsFhKJHXpGbkDim2rOy5XXgrRfB9c
wLjH/6K7JzFbTjt1d94/erQV0bxYuOXvDZC+BccrUiYhOdxGpTa2DUzY65ap5QucNXwQA+bz3C72
OCypa1N1BCmJsBu422qHufK+u6U1oTvOUbt7Pu4UjBKZZ+E5trzsraZe6uWqkYkjw1iFavu1wbcR
EMZb2mlR4tG7sSEO2ePY/V5T6hobc/B74u7hnAN28oFQkSAne7mIX/2rzYzeTCjnTj+yUnuG07+T
2h9dCG6DRJf/PnilazyfSx6TBTis0r7rDES0cpMu9X04qJrV4R5mQOVWy0PNEx2cxUzcOPtDzgJg
xMpsB+UXZXsxwZIF6D6Ne013hrGzBQfhzSn+2LHThhLdAj+BrcWwZtiAzALdqQNzUAwmR6awSJvB
OCAUuROCifSlyzRUC0GpgRrI7qIftt13HcJKe+MDhLS2dmwoHN0o3sUAXZr4S1z6xvbatVPAJsS6
BvqJsXRHz6oDiYBpdMJlXRO5Qy2DBrFTJ6oRjxYKFGfCPfkcaTg5SU8UFpce/GpaAm+OiZ8d34gj
jWd6YpkozoTvh0nSGZxTmyler5yvahVksgOdW/miS3f4OM3UA9v5RzdNnNHp6jWHwnbLJ+65lbwC
KFY1rLaSMolXQvLTiH19VQnAo6G/vjDl0sm0PbJIEMCiieDtF/4t9XqmVjKxObCDiMzUh7DCJMuR
63lukZ/mwjoQ+zDtb+g1mzFd8oqJlQ3YtiBDjXt3PLwh2+elcGCG5sqVOMcpGlI6zVknlDDuZ4C2
CroDCX/eKxVCEjKcZUFbZVMpmrQ4/C1IVtk6dUhefLyttfCKld33lOZYz5Ecj6slnD3E82PweE37
Zy47AhxyHAKeCL1uLwblUmZ2hFWztL/YUXnNRXzqOZIBsnqAwwUM9i2i3DkfWmUjLpYIyj/YWtJ3
EPb1GgPZx7w+AkIwUMVnp/5y9rri+9WQ7/qIgm5pqs7k/aWdMahQHWIv3bWAvBzi8PdSuLEYSwjO
JFyxrD1NHPD7a+KJUB9PWU7jRXq97L0J3pGbWOX0bt1CwqkGOW7qtdUgprptPYDIXAKNegJH3jyF
O0N2WsttNpzY//UCRIPPp9L8/nuiU0OqknAEznvNn+MHogxlCB+oDGOVp4qQklVCLC7HY18QFTYP
bRZvRJtdNJ6LVmaNyNdfV+Hrt7mqrYaXDynogv6Q/fxuXKSzTM2kwJ2EncbNtZ1lTBaXg/KmnQcA
iitfjb+UgqYR44BIiNalcLNElEjq/gyxZUA88XEfDnf3/fFumIYio9rCBDR8qC/G0CbFklNbQNBZ
CQzu9domWOcXDZijtZgMnWmikIsR9cyppcGtVKHd4Fdqd6p6WUa3cDrgbQB4S8sTkM2DOYTWRY+a
Fkj+2XGSTo3j8x+8KThPSx0apA94xxa8apknrhJQvOSt8OPVCdpdl1ig9XYDpP407R78bFVzhRKa
Ok0RevPDbqUg4fPZ6pCLmMmA14ArApRyZC+TmmsoHYbJ0OudigftGd9YdjMWK/PysB7dePuhp1bG
YEiKlmqEKteHT2eGartI0sn/EazXkHz7jigpr+9t+G07SxDCmXLrP5wgswZSUk6NOFxyUY2DMWFN
Bz3TaKhLROO2G+igztS6jAicqTHQxhuwLtJGZ8tCguZi3+22CvK0csiyA7WBrxqHgzvY4KTbhzaA
J6lMYO46f87FaWB7pu6KOJ6GQLc6Q48KGr46A0EQxMOEkW8hoZ4Oau3OuJW5KXxQJRVV89IQfEnv
BMK6czlXj48jGOdCNW0m66C4VQxkGV3Ubqj/YkP/HzcObD8UEdQr7B/z8eRl942M6pkUThkaeS9W
C463fM/LgLrWqEFuj3kZ0V+X2eVD9Dw+zUtsAE68yrRFm+IcB2+P1yg/2y0a/DYp9nQhtbGDIRIO
gm9oBpsZQn68xmM6oSJD6FO0WZmoCL0GZAo94N1TzB9mD8DXQqF4fy+MV0BvXanmHgCUJ6zfDTEy
OvBvmmRPYeu+8WrtbyViRohufiNdfLg79RjhSbVG/E1O8VoBxMbOjrKUBg8r+7e8etmrTHS023fq
ozM5zKbk88IDC6VnzIaHamxebrxoIh0yTVwjlt80XkC1t1JBLmqAx6FLjlTpdzxiSzBdo7AqPRg0
rLVSS0smjy6RVPQmbzQ4KU9TW8LukxEuHPY0Xwdu0WjGBjuxY0Pb9ICN5arWxOiwUCoGwXuZKqFZ
OjgWHEEEh03YnfDQbgZFBMM4J/w6vewLfhdsbNN/YQViqnQYDDAALbv1WNUQfpRhK3NnhQVW/Ynz
B8s7yfHVTNvjpNgbzIOu7LTozB2dkwXs0H8ulZeDehkLP5AR4gdet/cU52dd1IOiKVAoaxoE9qW8
7mHajvApo1taEYOnvBH/cmt7CjY+iEiwCToVNqT9NQ21Hqr82v+idVT4ozdJ183M6jkHfk41KQgo
tc7B6PqRb6K334wtJ+I0rE/UQ9dAfaKJf3HOf7TOw9ece0YexPfYdVupRdxRQsYrUDYzAJeI/hv+
v9b99OtE8ACeXRVY+j2ZOrlx+DzidVDxgjfkQSvEybLieaOIjNYTYrn0daiIlfQ6lbMFBNupBJsX
/89C/VsLCB6DBaW8NyeW0uckDhFJ6OmaSDWZ19VOJVgKiWzJxVzHZtkvGVXVBki2fSxIcxa032ag
w6gMTHr2BUabswV5Xbxycf9vxrk5GaRbK7tyCCwPcShWloc5+bbWcZUbtcKqF3RUVeT9HNDz+l/s
dHe+qjkcznUPMAX5dFds7bnGnUMuqmfuw9oIaNU5QF7O/uyUkhe357wL5zybcb7yaJ4VX09qK2Xi
csMCmw+FIFJF7JhCovwk2jckH21SmeHgPkv+ncBrXTV53Ugf80Ho351VyCqNYMhXLplzArLU9pmK
myI3RMGFYh0pIgau1k9vNEsLYqgJ8u4nunYM3mKjShFhDPRkU4itjTET6XKMqnBdWajppqJlhbEZ
awMCT1hKF64c7G1uKIzk+sSKocfsOo/FbaCVrpSsZty0C+lzi7EN69a2GQ+0SEqL34X8kug5GsLT
uflam4eC1I9WbZ/ku4n33wagD2fyr9DrbeErepYMtukFcEI7K+MdjSxR9koDun5vllUEfvV9hNod
i6iGHkp2zefMe52m29Kz3alRj4jCaEoqaYvjdCZj6y5A23lJA3F/k1Lx2d/5OXkKPQUM0U1IX/Lg
nLMZAJowVHwuSjQqiZf9lmYeiRehGxY0n+id1aHP+z4nTtV0/iEzYUNkMZX7YiQefdatVxg39a57
nc24XOuxdNB/lmTrG1dftwi2/KMn3jkiqC7qHgx2L6OovEoRCtHrJDe37+F+93o/3BSfn1g+R2Iv
VWh3tfRfwJwS6Ot9pDTedj0i3taR8h9NybBTfBwR62XyRYg9Ot9VpDiMFsphgeLHBMDi8RAcf4Mw
MVwZRFWLT0LZpWZ1mdx/XnTRlbiipGC6Ij4HdlqK1nLU47sEKv+UhuFzo5SszCf/eh8f9mmbkKnU
0enAG0DxAlwrW4qqvFv1veFJkZSjOHNQ2ismQA3mEuWerSxakFHnlCJsRtNlYJ2aHu46F/ylsMnp
/UOuBvQtIGiB+Wyayrpuo3AGvnILocTB8i0mfPZbnsevYh8V/+g5P7bwjLSAuXVSU64PEIAeynNF
QDrT0Yv3F9/kJWccx0ydIjKMSKsmcwrL7F4slJz/RqC4yzNPOMai/gjXmb1cK2aSng7HJnd24xVK
DqKVMI1dIP5EWHxSK2fefdeHrHZf25rvcs7o2H7/4884OWIL23GPV3/Yu24UR45gzCSShj8j9MAQ
/1UsTbjd2ii0UqcLD8MK5DCUMTaDL4LA95y4UgD2gB6pPlOhlI55M2VFF6CWmSp5W+Xmzs6qs5hI
ePGQYsUa1cRAbTCdHGJ6E0E/wB9t1jLOJfE5lFWc5jy6tZgPvF5mCYSZGdzo2n5TPUJo8vTtc8YW
bvQUIwiF0dvdyFkbhXAA/w45Reft3WTdguuLSr3EpqLU//tuaWkMfTvUUwjhs8yQEoEwt+uIbI8v
dVaFPqI7O1Fm1kSIScLKXgYXVlpOTZRH+enFU0FMKvzFGlwZZCy8MxJwnbwTIeSfhmwt10ZpywmC
TT418x9aUhb1R9MyPPoifAxqXND50QPoSUouMVgEatC/YpXMfoMhDhAQzHlBQqr7EStOAzpVEk1/
9Fv/KyKr36A8WUUh1n29c1dUnQe3F77JEhS7ZbFAxunmdyjGxf5G7/xOgbwkxoG1OuQDYax8k75i
BOXGu2M4kyoqsS4izBcCLKqkc3mHMQzsM02r0mqsud82zMBev5zz5GZnVj9Dkx70cwm0/OMuwdXC
Uxq8c7rES0dWg/ge8x5qq/uTCskjDJDnRa9xkWMxn1YMbA/zBiyj9ubpyGndp7oLV3yr5wnQM7U0
6YIB/tiHR6OohkAJ44vHitTtAYeVghtBFbWn2JeOaG2hS8/gNd0ltazdGROwYvnthcG58PhaP7nW
bICO2TQiQRKvoKwyXyPlbZr0IgKJNsIsBjUGHQWZLFYqB9YBzRX7/jVX3lY/6JLLbiXKsotldBQH
4tM9t8mbagn/73kpzg9soO5lfcweFlvxXlWc1zxQ48DEd37PA3iDsJmWMiW7I7Kk9iL0w9+4MRql
ldrvadb0GYI0Uwbx97ufloGuT1XCy4mb//jPiixBen8wGT+SDqnIpDi6ciZF0BxqBYG0Z0Uojo9Q
oMwXAT18GFEWol8H+yGu0iIIt5kam1kllYvnzqjHBAO9utT3yZqOFrl6WNTqWnDmuX/kP83w7WG0
i+Wbov834/v+E0qrRhDfjaaOFbl/H/vtk9ahxlL4uokY7wQrBVFS0k9M6+333Fa5DM1IyIvgYSiP
ZezSd3kcNfGNcPNsPWTcwK96YQH7QIDgOFvA9IrkuJlZZXJWPUz+O+Vn6KNtckpYUdIBUlZec0SM
8AmbWOkm78ClyXpP5P1B/9V/7IjP3TPcVnmIqGVdebal3QrugzZQcE8ubk2NSt/3DjrS3NgMJXFr
kffmQYAM4t6TxsoRwq7f3KC7b6qk8C8Wuh/dhIBuGJHD9yBzRV2dctIA3+qFyk8FcDJP87pihT9x
rT0NEtKfYZem8JJAjBi5k1Yv6KQFswf8GVvMIhfD4GZTd1n4wp7AqiYIhArK7Fg40wIOXhoG+Eut
r88Y5cLUnKZZM3r+uo92xw2lyvUSKmOdN1/R1AghVMDTJ/KehGXdbyXr2O7wtIaaD/FeKygb4EcN
UdMo+ZxlFX5AssaiyoVizDoCc/Vu4xJRAT7P06vEmLPedonwZdXTzTCIMcl7BWtV3/WujYnWkKtP
90xW//6aHptQU8mx6Yh57YGfe1zvEQOUlz9pyUnu4mGZ2Nz6+TMaHtAJdfG+k5rBaXGp2TwuAsDY
TODwQ1zG7CaylQaSKDb35d+WhyLBqTfbhkr0gEpDIDIITz0CIaNFuMDwvM5kHxCllBUPRTjmxyaN
KwedtVopjGjfvSPHk7vHT0nRLMs+ktDvBmStVhbGgHHK/F/IBaGLwKWIgnxCmxHaa7d1qu5ym3u9
9IFvDOeDGi0SW1DLS+wkC/kyVFsqBX+Abk+XoYfRl4BIGGJQq87YlNyIkQ0F8AvMR+vppoDNdCzZ
rxJI7FWAIFvDuS1iaN64tpEgLyATex8PiJtWJ7vNsUOngp+SdeCOEFQ3NLqBVsPF84NsmavDTxhv
ShCetRLOu1yI9N6yHf/7ui86s3eCF6e+IICd5rsvnx4Cv4x4eCAgq/7WcVl0e5lCHXEnLnFMdxVZ
qptWQrMFHFMV8qc1ZaG26s6eE8fink6KbODS0vGoOUBXo+IhJY5ekRIKQJTM1cYJIoafWCok79VG
6eR3woS+IpVDRx8ti0j5zCPRRZCzkHZdCZ9RXPTtUWtHneY5mUeVMwUDNBxgwjxUVlew2OIaiq6b
77Jxikqcxew5tMXKIaKJsdH3lQf1YE2WIx0C8jcABdHhXTpvODxWOIoyyuFpTh6fo23mvMCH/D7k
BtoWvP7wiMgXoP3mZxuGWB07LKK9/6bHI8avTEElObD7h1vx+/xxRcyqlisur48Ixq72CEVfAqOz
vtswIBG305Jv2SjuVhn+lOPRru2ZftEXNJjdxa7G5JE/R83+K9hSSzKkXHrB7KiEcGt688x5lHwJ
6XVMQBhsIP0AoAQMt1kOy+rc3m7G/+TOpE8DOK7eJ7SyiSntIzHIH5iS7znH/8sxDjcxap6Z66yH
dGF+JJ/bPADc+mk1LV98iQa+tA3Eg+Lzwo1nmgQ3rKNbhIjDYuG9H46b5hgcTuH5olsp0CQ3No49
NrPkDxjT0EtzJshMeiCsSoZF2QVvkzNhHkBxPlwfg9Kh0irEse+iO7SskY3dEKCn45YVPOg20Crx
5jd29+bmj/Pk4wH0SUWIrz1WdFxHAzs1p+kF9gPIqZx5WPVrw+WyOwobYxg4zl8/O0gd5fTVvnlB
cj/fkZ8JL39S/LyXO3PaiY+ScyjovxmJQGH2yqhsJMDF3e75q1KrlJRDDwj4jhDhffNdxDEb3gVN
vVWfT8aVHsptfOdHijpj0WWjA2JY4auKxAKTqVd8NJWBC9yR8iCIAtH4kYN2WIgM/YI4PpqBZzOR
pXDFeEinvLwTqFo8yOXEtWcIrneZkQltp5EkF1RV8sH4BXGbVAuJYkDot1onn7uAHe01QjX0TXsX
le+v/FSTy1TlhO80M7rDDIK0TBvBufYVFzCjqZhn9T8sYaeG28TINSntZ9Enr51d8G55NSShGXuo
haREMNsodOTK0G0YLy2zPYCCXSvu3dEQhrw1Cs0sCO8cXefKcYvKjPoXEiJI8uohof8Izq/FU08m
92lIa1MkMcIzSUGDGc6mnuVaxKvEZ0KCzOn9ZBpl6IuWIwPis3eAZ1rDir/YNCxgpHr1700ugACU
H3WvGunm+5hMrE72cin5s2wvuTv352MU7a310YUq+qhMCxByYPb//DiUAlixDOoiU/MvZcOWgAFs
+keAu063wXDx9/B/h7/cr8y2EHaj0H+4/8IgGeZRKaIt3FKNZ5+vKThn2b4eD75F2xTWBHDL247I
i2uWGofaCk0FO3MrgF4aIGpuSSdFhRd8wbgqifjvOo3cc9wgl7H8BLNvc9xsspc/NYW5NNRQuWWh
t6PZguNGV3w5kWxqy7nGEaaSUxYxENIV0MVe7lAHB3Qg9cEcKi4Lbyu4yfMa/KjQUShjlNaC3dD2
bSngGGvLRHv40ymA1jEtqdhMXT9PiKGQZv6QclT+tejl/beYMT38wKh+C6jipeDuWFueznXa4u2z
OIJvHXLEeYQi5jEiljNlXMAK1UVxDr5wNv73KaZVjo/4ItP++kQK9vzjhYzvtzX9yuuYFlh4ARp2
cuPHx3aGUxjJ5vY4yXMWsvLKBszMDHEENapqLDvVEZL/Ae5S/8TZIdcX0xquW/OReoECDqJcDKQS
cMWsht3VC1tZrGzXqFiu0uFsR1dUGjizXk+ZBT4xgCguHYlLxkF8Jv3KdCOIEMHEzXnFe2SiTUb8
JVxYmfABMYzHJDVIS7ygSRf1DBtbCoEtI94HBY/rPOcTbdfgHwFgFl7d4vZnAUrfyg+g7WkJnePh
PbzGSL4I9DKVGJsUA4HEOnXtK60vLx1ecwyMQRlaGzup0XF1L++xo1J6wK8hA4iYdzPC4t9+dwGv
WaxfT9nKbrJWjKLlrnKClY6L3mnfiyjz9EMfgdr2Ui9bgaHZoh7X4JG00Nrwc/eFEQizS/TX2Dsz
t+AZLnAifAxkRaMwXgp9WFvdfw/Bh+6VKN2IKAeSKlhoqn3H5TZGMNWmXC48KQFK5d+rWW8cwf4k
fn6sVJLPJEytjwC4FsvMvyD39ATZ6PIvtsNfhev1+J1s5MxODisS9bG/LT4voe2fFjhz9zscozQW
X/lDAthWr2qHHwm9gPi2ailZhtBFVzxNy9HOcTjOft1R7yn4KOvMSqFGUXfvt1tQhS2v3lB5ai51
qHWLfAkxzrXBO9ohsFZI/qxHHFlUM70Hk02A3SAMNmie0mQb355mOYNfgcXMwUx4oCoZ4FD9CYaa
m/gtzl9L8XLauDJ82+Z51l4neYp9FDwxA0EnIK+RYWMy15gwczUjzwqiNdJS7wYC67/ars1LILVr
8PoXwP+r/dUBhI93lrsZc5ddBynbO75XoABLNhU92BbcdRDshydn5OpmWOJrYBIkOmME6Yp5K1W2
3ckhjEFH4/4YAZ8b3/zhFSEzzmRpNfjTK+atcLUnO5mfiNFANY/d+xC+qVKGGAo2V2HbRFUfbwoi
ziKCQmAJd5g/MEtFLzASpyieQR6reO+IkAwSdZH92Vr2MEd6LhkuhqfgLPMoqFHQtH3gIHSi84lM
Mf1IhDHNvnWNw6Zt/zxR4qo7FQf6ieO0ykJm00+XuM/zMDl7Jn7tYTWddwbrts+/aPSO+k9g4hSu
FIS21GIEBO/f73mwiRj9ktCaoOKX2i7GGt8lszzN03Y1eGzHH9xB/IER2Mww6HwO6IcHv3jPH2wD
THiOwSXJCBLQGmEnSIH/zjh8MTKVuKZ6Nnj0jx/IGRIKEzS0vRNjXwSgHN2wLwqTrp0vSRtBd45b
nG9HKgGGVIFhnucNEm2VPMBbm4w77gks9ufcjWig6YL4ug3V/kFYts28sNFGpzDqYiBJMn5U9OfF
XigT4U+29BjmnpXuhgXWFM0gBU9NfIHD/ii45UeFYg+dIIu1bMO+ellS8JDTvqGd3BPEeavrTFip
kGIEGZuRFJFoAk7lTLxrzDJ/1pr87Wg2A+JX+/zBwRMVQ+gaCvLdMC85tkhibTmiJTPzjJ842B0y
fGiqXjbjcKVMMdw1Fxm7fTUr2mZl5QlUYntF2Lf33jnD1cVuVDDHUOeZJE1QOm1t0uoX/7wEdVey
LUrViRH5N0cWA8yfK76dOv9IEAGt8Vyi7tTYSkNYI/VOjO/GL+QxPjYqP8OZhxy33qTHravQetzB
j+k6vLQitnMRe+yAcVZkbu+qKc6m5+1LOf91PbpZcH+pVZnsT+Zi8wwpU/j4FSPpd23EHhOQDJfx
mhyXpE9+dJu0N98ljV/KNI/GRWbTAyuh2YtDVPUW3nFucvAQQtTaGKHlR4ILZrfQKL6RBUdYtE/R
/fR/PjAN8XqRRuc/CylbJns50YU4pBzZ0h1icl3IXOISSrVAPQZIM1hdDeqeQqCFkYBgBUPyrDNG
ZKjLxxBEEXKBMhOFZLPgZho3AU6rg/O7in109a6nTipbJpBk6yPwqRG8FJoc5vgHTERrHxDV1XHa
fhsXDA/i2qBjQuAVVD/zVQbH0m5HAK6MiB+B95GLJGxnAyEcyLr5xIrC/270pV+PDnHguQ0NS4F/
i5MtL4arm7j1EBDuZX3qhLHCS7dDaxYdQ59dGtskVrpx9oluVk42YDW7ztuDcLQWozB6YsWBNNWO
qtwYpXRPgCoLdTzYV7uAT4kr5/HVZ33jfrbu1vidiwrOeVI27AOw2qRL93Qz0nKbPoaF2AWYak/S
U+qrVxboMFMVi+WxkdYf3gjbetKCiWPFsf8Gy0qd7KihH7p9Z4uIqML60ABU6Dr38gfH5ia89ZpS
pI2zQRiJOu2OsCHUrNajKb5F377yxfF4461O10MB2WYaaLz2O20o5qP5t1u93D5crMKQEqrStpsf
N1lm9VoOQhjBym9I7AIRB9Tzq1Bz0KvABEH8YIkVvj+VCheeD/jRq01ZSk8sRONFc+VmzTiXTuma
/gfiDmMVCpyuvWkG8IwnFjfUU2xSkKdK2AjqaD2MnbsHtHVmxnVNVEKbNB20MUUBv7HLsf57wr0w
EFHlquXZ/RNzWIULPwrWhh8BXNw7jHYnfzYwdEHE4pXwqZiDUXxyqcdwfy7oAhJ/ub8yZJzeFirp
CIhwNmmeVyaKTqLK0tm9LTlZp3r3jK51QHQe8TbGPGvX1441l9TFL4pzzFONRK1de7n67qqbLtF6
oUyW0RCvImVxgT91DDsvVe2PYLiHwcfdXJdy60UjmMKrRfazm/TJ+I4UGSIPpGE3ddDRilUk+6qT
6I8jgIR8ZTaTqfzLku+OXFFOt6ehTAOqVHVnn8SlMre7mMMtYU4/JF2RvLu8lHAICd7d7vH3sCiQ
w8BZf2T7vouZV4KwqwJeLTa3oxGruVuga7q6wsApOLEXHOsLESVgngC7+hxsslDYlCpEi7Z4vnTG
PSOr9Z+vkZWPWx1XMootKYR9+tYAbI99grzm8vWYaX7OK+8v26eg73EB896c64A1YCz9JbEaDzW6
Om7BZCme5QijJblzoYo6AwIktKvFMgK/y6dgBY6Dml4LIe4anQHLrJIXix2J3zPCxUgPMlq/kCwq
5nNmkOXAGDv2U0kK4OtvwsqDXWQMrNVFcbA+ZiLMsczvXQ8/dFVi+HB1BzNFa95aCjnAZbLiSEvC
0e/5cbgAuPEWc+Q7DjURUUqv9MklK0AGDh3KbX+tDIVWjKKNiDhpM13YKr2+lJnemYXoJWM84Hg4
G/V1I7plbdUb+xY3TZxR3mAJy1nglwpqehq+b82QJc73OEuzwp0GI7vn2XuaLEUMvdrs527VpAKs
Qri1Mv+gvOziUVYNhK8SRqAOAljVImSVXr63J6ynfpKp02zycgAfGbWIDXaEQOB2hoDHbMJuUTVX
haamBq7/EMrDmq06TfKaQDlMvWTVW42ZWe0tnGcqEYHCTU5OaGsQashsd7tjs20Dse2Yq2kA4OXi
2/sRJkSPFK7GAFcXvQ0nTbXSpugnBssUIhVxxEsO7tm6pmimHFKE+SynsiJ2FqPi4cqMU+fnGke/
S1okBM283YDEDtLrdQ3/UenSgUGUQF/D213TvXKRflCzEol7viUAJLtFIq2PWy1mF9ErYQvvzAih
9D6+/H+8AX1Rkn9l9nwUGx1duZ9DZsHrJeUNFQmN7rpoGv9+LB3u1rLu/kbgtzoHJq/UU2/TggqG
AVp5SQjrXE1zW3OCR2jLinm2mHjazRNzw/qUZAvEAOygWDR2hco+ZjHM4Mbxrq7b6Z8d88Cc3Jto
+VhyfVodW2i4qlZvJNr6nN1csecFhL1kOpo5zCR54jXbvKueOQlBcD6BdhSy+Dv1K0XTeLMa5TnT
i9Rd+f4O8TpRZtFUJeOv4CavJTdpIP+DAP/Da8p+2IIoQfMJz6jzqNYLLgphZMNoOuAdakM68HAa
grUK5+9tpdNjXLqt/M6EFEnBvqM3cDXDnR9uuh7wkHDlhSiV8ZOgXje5lSrRgdDkP2dHm8IOVZ54
49H5fOA0OEsvFeqYJoKm52dmRZoG3HqWAFNJnL9OJYE6ufUYXE0Up9u9dfIN7b0374kWUUCkwaLj
k0ybSwYR5NmXcVpvfs6R668kUo6bNwmgIyf+BQ4qHUvfGN2awR5ENXFx1YuawHIa6RTmw8FIqu2b
LZXbcfqvHPWBfPhSWDlHk/dR2DuroNRiUlkbDP6kp40MAM1rEZYFwREYdFSbpANH5/WLk2MYeSp1
tSNpWpC3aRAbasCONkbvAnKclBrvrJKeh6AH7JwiPTRJm2oUgJvgq4Zv26Ow5oDmZeajVEn4s4U0
2VVnje73H/0zUdZ4ARppn4XAPWw30zeZVSD2hyv3WZUYo4LTnlpo4NCHrg/xWSKfIQ55wXJQqvae
vWMhZMKoRhE1CEBmow2VAB2rwh8xPPmqtZinnSIqexpuMm6KXae0vGH39Q0cR0JVOSu/MCXbbeBv
WyZTRsWD3zCfkiwA3YjPSICWgqykaF4nR5UJveXYurYvHfmalL9/EmcFrmgFYHXHVfcJDJhggwt0
FEArYsE+FQgloQlrWryV9CGxF+oVASjjQ+k1PCB8vaHJQ0C9XRo6D8i0JOZPD1RF2ukFzVu/GNTj
WWlKhBoPwu4ImXhHO/S6+T7tCKiVP3LD+FDu+Xv43OCxngaBCchcUCrAzf0dIJ0D8neBeNn9xQ4P
pkKzk8dY786LZGInHHxfSr80MZXCe5bOMUYD9RAoav/N6PE7mlGqLST1UOVJ9jQa8zJLZB0h7Cgn
IWN/7/876WxtdP1a7wVM/2eY4WqxnkyhUwdiC5PwEJ7iB8CGCVFwo+Cp4YR1DpaODk2PU0nAxl/Q
RbhYXeELh2O3QFGDKS4c6EALjhYMSOHTuH5Q7cpjiWJz8PCCc2bE1CIKbqk9UB/f072vVQoE3UeO
X8JrqIwufe6RzzXTjIYd53cjATqQV1C3r+KlYP5EYvb2PvH1XpaJXIRVWDXf5nTr4EtT24S03UrW
XKdymJNXM3hNyhM3FYLcRpQ3Qm2XSxS9Ep328obRQ94GMFQWAkugCYHkY1UBD74nU27QaJ3DpZhy
r5kbMyHNJwu7Hr1mnpsXEC2ykH/ANCX4W2FbWCOUBQq8T6du245Uy/ACy3ocXqKhr5BqJZ522v+d
DOTbG4ppYUOpJmnA3IM8K4EGkgYj0gMIk40B7793kZlVD5IatmmrjzJGeNulYhzTm03+DM4h7ZaE
+hwcSD3eqByDrCcL1MuDn//XQPoBNzAofcDuchZSfz6j022NxIRJ16GFbnJ3kOY009mMDlBEchnP
gfNCePiNd+J9cUjEPIrOmxjxQ3na9FW5pNiyydD0msfDFn/b5R23CK1i/SgcT9JSL2pibwlfObz3
DsQVl6I7/d69jT4dsle+08JkWlWvzahvMHL36nJyB9QHPMU55cVycVravx6/yYyYp/Hyno4L6LyC
LtA8+munl22OptYEIpto4v+kVZulqejSGEuzaet8q3IuaCKAdJRLwvSk08EVhX+dhoDNiwWoFbg5
SAe8HZF0A7X2UkiLiLFbkfWbf2x1ZmQdcf+wCEy484KxdHvK63a6lvhot1VofHH9oXNn9Ri+CMfM
gIQhivzKDSP/oCAejxknK48DOWjFsC9iyhNDKDE0tNZeKVqG3AgHJDiEaobfsWlPRFaq7CE7CYHx
DT3GqyMP6/NQj0S2zr1bV7s/afpggE9CLzq9xv7nEzIA8W9KGQf694ZycxJdOtMqHzkzPgsAAIKO
Kbt558VoNjBcG1S22rtkqx92xu3ZdAGRvvVrTLTZwAvroDdFin7O2DGfPH3QJ/y881Prmvs2FBqC
8Z2cHkKzhxSpft89TH2vW8mOSrQSsdciG3dcIcqcEYfT0XTekjHaor0kSq/bDR7rYBfvD0yymMjY
Uq/Ef5jGaSlareD/XGumGPOJrA9mpFGVsVzSr18KpGZ+X+smAYNbT/CgNvSb2PYLU0MKN4Jo1jPr
dGoDtxn4kH6OhWGUdfqkJCXiPrzfkX9t6o/TkN2kZ4IfvgxQBChG1U2zESpAuU3Eik5rW3GFgS7F
ZUJ5IvyKJdVFqSjFRm5LX6MHbudJOcGt2/IyC0CJcFT1Qc0d4utrhHfnLnlBWaIFOL6JTsiRaHue
4oACLp1RB/Tbg9mz5/YOpWLffyYNWN/PbSs6dcupy3ykhWRh/+jgpT2JPXDsKiz3N2rZgszyXc3Z
srDzPYAOpU3qtMK4aeWbKKxfoSlDSCLJil0slCqYqUE5wuDlsg9i/Kzg/c2cMDEAbJU5yl9a3oZM
Uogce2PuyrcEIxwouo8n9YlS+XDnjTEXT57krTQtFgYLw+VKM8sNMm70yVP4xcNm+QceHd0jkrCQ
pgHMY1hbXu+NWGEFqiMhgGzJt7OZJbq6gR7IC6L/XnhbUPMpAdFBMDrVtW23NiBpo5g5LqigC2s2
1+pI1GNwhH+F+xsCUR+Cv74fuIFliicT1ioMZxrOuJL5iYRAUfgD7mzWw7hn7Gc0A2YWwCao2imC
b+Mv+RjrS2gOGRB5glk3GZZJpjL+8bn/ttTgydFFSTJ3a/RGRcT3ro0nL/pPUz8wnXog5hszgJUU
fdhojY10AZ6gDuz7H22gJyEHOhzWa9/qB1FE+goJTbRp/tDI4xnYl6aF/oU4xvm9Soh4IxY1BqdG
r5NP0ZIY9mzQIn0YCIUHpGCkLafSOTl5y+9Npsm+XqaKt/pdDM28frSL2co6WuQVIJkYvJJDtW2X
Ur3f35KwmXYKE1Odigth0bfZUz42ywm1i7biMQwdnOWD/UckPQZq6nP8X6inJJOIfHJgWVUgdzSm
Plc8qTxbV469XnGUTtNJFh4t9qDzX1znwtbT7Jh6s/EQtesVeDsgx9NqTfiVSwNuSlYW+ToJxOvq
BIVrEv4zqOG3XiBtthu7eSWmf0z2Xuf4QOvTw5c70aBPgx0CPpLS51prAeLI0AfnhEM/QcLyJsI6
JwnzkDE7kTscMSDX8av04O3YWRnTN4WUgLGeTDoO1Ow04VEP8VVLsngs1GFWfJvAT4Q6WTP5dwlH
v2R8G+W2oM07v9LnHSfRiz0ZiT5fVfI3LHs16kLzOqtdhelA/rZT8tBzM9ZCrKSO+T62iHRbVRgV
6pz4OqH7CiQO3ET0HCerYAGB+5iYCPCsnCZ9rByTFasKebC3sv8T0FeVkH2dtl90B+rvyxvLR3nF
48b41YfBSpE2awTvaBrzKzKuwDq95wanud2ETXJoZOapEAmPJsA0LylwGtodJw0QuJjSCR3eIl4u
su/JV0qSUJOl2qClrxEUE65ffmAMsi5xobJaB0YOwrg9SgyIxyLdlZrqWBo9csFj7Hi6/GtiMCeM
42T469LpOAb/p+UQvRlsuMRtHY3tbIUVyAuj9NpoQ95VM5j6ijunk2mpO6Ge6AxdC3j/WxlZ45Mt
+ZCNtgxBhlfCzd1/8lPIrYJT/kR8SuUrSkb0qZR5U85L440g2kjy8sFFTWVWnr/+nvM9tXlCBWfH
qUTIgak6r5wVX110fInI2OJxXJHDme7ystnRWT5VgxRjhfSPn8/gmho9TcJyOHz8taRJdGYV/b/E
cDMXabkI28bbO5n8i4FrfyKjSYoc93hhfQURh5aZW7Cj6Fn/LVRbq4znUqFMoTKDlikchVRi7jlE
th0rbcYBJlO8K7Ig7STwl5psce2nxa8Cst0awfOjp4OpR1dsHsZEsJ+lThe3lSIJmqb3yhU52Tt5
th8nxkxUHrfRkFZhI7Ytv0ChFpeU+WVT3COlAe3PwJK7K6fUG+xc2DJebwAAsX9cnLeDlAifJ288
5Wij4M4OGf9q8lWA3nY7fCGHY72nFHa3Lbg+RR6kM2oq7dBBqiealyHttSMatsmOSvLkCE4RPHKR
pNeydJSlCLuh+p8pwlTYDCQv6zRRjR7/VAqM2pBNPNCy3151++icQ9aAvAMO7rlMgIIzGH2c0C0z
OpWTQaSgj2k3UC2+bZRVkEcML5+mdDlyG700Z/TyMjOkwUwi+1NKNQ4bQeGLxql8xj0bsRDNo/7B
4K6zmmm7ZhJk9DURlrLl90l3PJ7FUANWkTsFLYfqYs1Yov+rGfmsUb3nDhwe9uege/rJVZFPrV72
hhF+LsIjzStPzgCFVH84+sqMzhJI4U9kvwZXP6O8I+I67XktnP7rkLLnA719NsrSgBYptnRSC7vc
d16vkxYD/gs6qd72RdkvprczFRLoEfnjbNvQ4xOxj8QTyeCGkHG2BgU+HYmDNILd/br4+FLz6Rkv
sRPPWQw/80IOljf2pD83sbbfhMjQ7mi8S6wGvm6MeOdJmDgiIuUkbpLhZCUaJMAdPJtVHAU6tkU0
C1Up4Ve+N5hFQLGMKUFS7wMT054+cy/DeljVC+Nrh1lvQBRUI9tA4p70U71HvDlP8TsMeSxxC2RP
B3yyBFNIRHuot84PQmQIe1YHnMBNPEKitPjT0qGBlED/XB5KUh5Vxmk4/bjAUIEebLiWi76gb6Oq
sztvXsdV/selyrO1cBYKx2w2NN7yabrwH5kbWWl+1Ydj5X7i9S97iMmIPZuXtmDR/oUegAPmZTdu
wk9WJkqBnOtQG2p2SkNfhWZAUquKGo1lGt68ra5twmGCenjO//CvuOKwM0Fr2lK8q1TYiipH1HQp
Vq4JkWYWoWefrstdloFEQyQ9Q4bsApsRBic2jo/8+6LrrWmGLL9TiNUY2C/0C6Pvh7uQFV6I5vzr
hmvqi1JA4vIM6Wk+MD3fk8cbhQx4YrTeZhlya1SYvZ/zd826dtN8Ei7PVYqrJH6+nsC09wbKeVpu
Qau+fHZRSgZrhH1lmo/Cg1qo4wHBA1eYOOXS+Qi1oDvxVkq9YJi5/VoV3Mzs2FPekMSRJixeXggU
nLhqol6tgYzq5OOMilaN28vumJDTJGhwQcpbBlcHcRctJ9ASyVyGQuOUkxffRKAyK6D0J3vnLPkK
WaaQSBPzLo3MVffNeIR7JEUmUpZS3cfTfgFPLyygvbGlQlzoWkdyMrkh3BlrY6TGgPO37Vi2Eev8
NcRAmKG/zNy8ihiXI9+qmBGEeI9uP+V4Ie9muIRyiYgxVtyJASFQiAKMb/uqh/xzK/0ouYAKA9JJ
ehq6sFcrc2rOlKbVJpBdhtvQ2F9oXMoU/QwbhoXk7kBHRZZ/Vf2+3iMDEOlN3HY5wESGU5P0Z7Gn
J+YH0ZK6n6KnxN5S6BhLFrHBnzR+6LBRpIGnb9NPLG5viR5I8IEdoMuyTC9y5W8puvlg2O36QiXE
jfN8AQ8klTuq0X4NEOAR2TuKbKWMFLQ9f5HTc+Ub6PQTYyTRRJpq02CGWfCnlM2rQyEmhP7VBiPm
0eeqL4R8hhqpYcXfOicFXBViSPSZaN11DMQZqAv36T9gGn52LYVbp3Iobr+tsRCA7oKaHRwKJ9Ix
yy5MZZgGz5BirtAE35z7Tanb7Ji3LwjqBug0OH3vxOpGSIusx0i1OhpmI/gevc9lDpRwQWDnhBvp
P5OZlRLMmsSu1JwYenHE7qTeG1O1rLlWslbE0V1VhjMG7eNLi5N0Lo01sadJ3NMyu4Ts1EHsqH92
9BtaVOLonSmZET61yCDmLZBBeCmxw+hqrheVE9SAB+tIv1rS2ezQl8o/1B8hvO4F0wWA1sZxWz0I
t75fPJFNMkqwmbsFv2vzybrfMawZaek6clUSnGWUDsFy7CdeJFFAPqUFrcICgUZlMuUcrlQGSsJa
GAjEfQumjD7jAqYwf2yqey2hScoeBK9VMVKx6LRKw8VxU/lGIXO97OImaXwRmrBX6qC2nAEWtLWR
iDFAU1MEAAkLPvAadBsTuqIufLWwc1YsM4xuCI3GpW0MTqo1ejrZBI+kjEV4VXvMSXJhMlke2BfG
VocqvQTmeMc/hobcwjiggpg3YJMbuhHjspe4hyH+qQHhrLaDRmtZ8Qsz6KzVUsstM8oOznfLJPe8
XLWBoZzwAd+tHmSrtkpqrTCI5UsKlf44WWuGbfsXkOeISK9Nqr1pL6rKUQqzpVjILLPY0pMh/oDR
WtXEoyDux4Ffzf8GUaBQTiEi1v1UrkY9ym4khTjC0ueuf1dmdmJYIRc1oGtlDYl8aLwnOnmyshfV
UvqJVdLV3Z+rdDnolXEqrPP5wX8WM2XElLm70eTf4lYPvhL2PfdxCYcKMFM0n3G4TUuFKFybmN0E
kk/K+Ox1xOPwqwIzIzXRpYFoUXk9rrNgMyB9Fs4m4QizWK7aAKflYBSuFVz0ZobZo4q65UauyQmN
HkZf94NmZDd+p2C0kPi66n0wyd+Xr1/BwQZu4DAZk6K3Gs2m3wsHWI+srHxQDf1SoeG+tLt9pwse
+hyUyGUttmDhm1V9i761SJyLQB8I8PVhOoiSsusfUGDd/VL3ltK0pEVAs/e5Y+A9cHWsuPsuRvik
AfHorEgjKBffeihxHfc1D9CCMIG1vcoOGHAaxR3rSKF3v5fM7QLDNY5dljH9xtg5l4n7gVSMBCT5
h908IGzMJlnIQz+/YAhuUolwztF3mT9vnrggxP54mnWS+FCf9pY/H704rPTItqYfPtzX7kRPGftv
v7eJz89gldKmicy33LjAszb5Hs+e/gLFgCxPPNlfvwKOl1IVHAFDhSGYVHAo+auok5pEP0y7bl6D
W4laP6jG4oHO5mrtdwN25T2Jq3F3GkXA1su1mjZzrMu6bWveBPfUImdAFDZShuhCG00yLh6mx01/
hQyI1/6WfZ4oQsTj8YW110CAQXkPQZB3blLcjAuksdGfP5j1IUNF4hvSTC2xrIiVecLAtfepG1vi
VnWv1sKmcL2EnTf1pONHzStiGPLKB58HS2wZV0mSAHgSAazbjeCTZUPVSPNmxN/A2k3UNvCR+wNz
smX1aCK1H5/IE97TWAi5ogtyMCiU50KcTApImsjFBL+toWj9/ARrrj7FK/67KEybKiU6HZOoudDO
gvXyqATJuxi/ZmsIeB3TnE6G6zeKhSXTfGxkYq85D2oE4ir/6b3ZLgfYZvd8EmVpO0ooWLedpCkN
w8k0OALxhxauE/kpQg1rLAIVIp6evdyPmEH4n0uLAmI0vCG+ORNkwko4Gxj4CygV3oOpgLxkg8P4
uUgAb401OPRv+NVH/bi4lHHafqiV0v31D5o3fXkoDF6ahlJjUSrUSbeDQsq2iHyxzXfnE3lEBFOr
Pb51BGTLwiisLXrME/NGD7xVHM230X6rd5PERSjPojqHokBe9nj7UasDHW3Kjn/Q/K4ptlfT32jk
Lm2koBuvlIKxmwHTLMHVs2oJgMWaSV7S0wg4sVZdU71HtQWBNOVYwnXRIn6CWaWxYvLPfYBIT9VU
mLZZTgDp0UQKr86nPF30aKH7foGobbatAsAuk39l1VFqtdITKpi6lWXOpXbb/VFRS8NN5u0QCUaE
8hkT6Nbz0PkZWAS12D3wsKRXPdDNt/hmjz+uhrzB0GC4IUnI0XbznkUdfe4olB0RBiraZIgxahaN
RgpnfIb/viVRI4pWtDqq8bFkI30GL/v5lV46mamBJkJe6MhcnEAc0c+RCrvLcONuiF4aF2sr/21l
fhcQcbRJ3N5oF4Kq8CppnWHo6M8sRg5wd0LkFtU4mpTh/qdm8aefURAF77OAFycxbOIT2uu2JJvh
On2vP6A/Rb/EdVwwID/tmLse73Qz0pCRoY2uZRSN0elLBVW6iBtHMSbNzCkq7UBG6caGxlUNrpMS
BxxPmaogg+Qt1D1+8Tqir+kVWFNbtGq2H5u+M8gZGBcELldOn4W04HVATyz/B/cHi7mEFii4mF87
OWXZ7acTVfhpJS9f2NdsZGB9GM5mc52n/W5Us3CI9SurM73uPXUnFc9Z5XxWzWt97fPXjl+fGPVP
PJDcrtqJs9FOAxiSCdpIKajA/9+kMkvbL17qfK7yBLUBWIh1/jLyKhHm6dVk99PGPJR9d0JhqlLz
m0LDyo7iM+k0d6X0olz+hdhp4XJM+cflb3Ti3shbZKZs0YwhWp2/cCTYGQu+LH4Ih/NK/GSLRsOy
ulStWCns+DflCsDHbIZYawVy0g26bkG1E/5hGLnLzOFNCkIxvFEsSKoyRdosdLWpHmUZUGQvluNP
XjUL/vMljlvkuNnrqYF7Dv1220cjr7I3Ca3nLFExFhYrZ8qPx0xqgGNMyRTSe1d5JRSpUvBXBcHa
6E8C/fcdrpU5amJwj1FhaaIX22hBLLvPwTQ1A+2ctvrKfLeZOmh6OudqVfVEKopiydila/5drST6
mkyR95BjUU/I6ylhh9ZAIpI5FL//QHHNYL0Z7mXZpUf/GcRaMlr8XJtkCVZCVhaiCHjhHyxqIJbE
jkOdDg7466k4MapX3eI0GnOE8wBLjLlEOsPfh/UbwbdddI83VVnA4qRWxdtTsVoXqfiV1b1o4+wV
jxEOLxLqjRtcIDU4oXC8YpRiFflg4tSoNSbGS3CqCuVr9GbQ7YVqRhh9joBNK0J80D1dVPNDzoew
PA2JALDS3M7lpxOafJw2EE21eV2oKEsCPX4eC7nF1a3XdlxfS4WMdpI6B8EhGkF/uToDB2Jakx9I
6erM5waLs8arA7k2O6CTesSRbYfXUHdxYUxjfYX0bjmpKN5XfRDeDqqNs/MBCMjcKYxVGyAcooL+
a+gux5z8MgFQTn/R+SOwDAyq/71/+DM3iH9MWU8RtptWM6qFP5lfhtp5XRwY83an9bLQ15sTENMl
jOKZKy0UotXlTQzTqedckfGZMqXb3tPN292hwQonBiJGI2tlyhkfRZTI82GH1OV0XUSzuXKklzQ9
CTNlCipRaxl/gb3r6yMlb9XrQAM7Waafouknpp1JulGOl7DIOqHH0T5rqYrjr9rGQI2aMx2j2wIs
O/7fGeYKbDDtVHhejhr/VW29y3jddCgnSFnHrvufEHlWc8NueBoLn7a8fyhfa3ll0epS0SMdoIiY
GyeiMlwyzFXXx82kI4YokOh0H+Ykzz8kNoahgOhiZEHAnE0ZbgSfyqA4M9WOmD9ylrHRaarDlOZv
w9HxWoPBKIIy/wgSq+5/nx3j11ddRA6BZ04VGNz5kjuBNx+DTXOjlvJwCxD7/VtQwjn2hBx361ds
Fwz7Oy4Oqf1rKqbCq95ai/1coCmJbZjDyyOpYKayafKYX373u+o/asWBVGcNC79gFXQ4BIhGy2Ru
xDxYG3kQDAus6AsVqrJ8gTYDQ2/fzfzTDAvKs1WZlm9ea64n3UZt+5WEfE62Jr7xr+eazsUY46a3
PnImCt45PY4VXjHO061GqHqPyPq8DVrD6OMP8Dj2SVwiEp1KA2RtspX6hiZ6iun2oiOOxji24qdM
oaA0CVMkmutS7m08pmHzQhDuMgqmCotRBGMAf/wE2Qvvdh9vZrJq/zr3ODiIdnfcIS1R7B2yFu0c
VWtZ2w6pQmudnypgDasIgNOd7YA7w64pUI35QI+tuT3NoAz1p+26CYbmh70WnQfOEtxmpYfoyN1a
TdFCv0ZLK/pDyJd3OtDPiAuuK0K4nHlifR9TqxwuNS4QEeOB/jvx/ub1G9hE0l3BDeorI0w3QCbj
94PyqVtRB+IKZIYTlRORI5PNzrzwjUBIl9JcXK5r2K0+iPXz6NdIP7ZQNjdee6b01Y2muIVWjA0v
QiJs4NI5Mdns9lhbGNDAMg7cvqiMPiBZ3pkC2/YgGDHEdYw3BEGdmx/aN5YOVYKpX/l1OtnqkuWi
zRgL01rRX8NPyNQ4l7jvnuHC0TghxjMW54s5o5pC+yK8jEM3YJFHMG7Mlz7A1nuQiY5zHNhyUSTc
GaoQ3E/2zmvXSS9P+W/vNvwHX8hDURJc4jfdd/fIdh5Efe+5CYjoJCjZvwlzFljhFHgjYIacnqMg
1FsKFpw541XSY4gPtu1dWxj2yhfGqyx4ApDWpxktN78BB4F+LBqIzeccUYGGJUMYFNJP77EKQ26x
A8u47czUWHWtDI4zbwiojc3Ig2fagp+S+jIFpkAIcB4WtCF/oY5WVCl3IP2rlAHO5+mO93Leu0Q2
Kc53Vzctc1bW15G781xDlbIhwNxvkYOUuxhafO5yvIkHMU/TGttj4W9auOtK6H4f1PBTsMj90wme
PcYkvyPhAExmZIAqr7xSxMN2nHYpKgbVxwUdYfaiM78d58GEkHidQLlf0dofgmIClyI4jMyLu6jL
sa+RAIUo2O9m0ut4/8NtnGMfJpOdlNeGrt8nGQ1Nxx81BZekrxtDG+5B8lmbtBKaaJ0WjAa4JBE0
qYYWr/jMpCUVsiO/VcA3wNmfq2txtyp8TKrEkt5TINsxpZrcm045y5WHU2rOPoeZ5zwdiyPu7q96
DrsMdaMY9mtFZ1z0AMJBo/QB7I/zf3AlJbuTjYa9LPJh2U5SHaUHXWEfMAZ7u/hSTrF60I0hLjc6
MY1+ELtFgOSJn0Uf6t8hLMBGAa8VlcgqoBRlyG6pIjastR6bLIutg/iek08mDoqaUHcrSikyAMUW
isRDWfUn13PcR6gNFbUBnyKMpB3+w0dYYRUlw24rvSyf92djlHol2InvvkNyxrT7BhqSPlcIh3pR
ir11xIhc+lhw3mdGGHEi3gnXDg7hMcF07KueSlaAFsfG8ySgeoeGJC5JHbADTpymHhgl/QvYcauB
FTq/weKjy2wOvCYdqUqZAZ3S6EUZmGpmprg3RrdCFEMBm5tl+2r+GagJuBSepI/SHGuYmbsTcyOH
ZmXzXd6c2maFXuuHlkzN566W9OgujuhmAu/EGBJZ0BzQUx0QE2xAAKCQ2As4CeYZe0FR6kohge2k
Y2v/kafRg0VYlAKyrhrjqMJnm6wb3ZCnvgTfTmn5SEpIc2IPqdiKeYJeJ9Fr6ghBCsTRSfeaGcpF
aTX/l4t/VHFALcA76C6kNFSYES4BZbRibJ1D5pHN7uO645t2fMwquFCisjexRoYX7jmPf+fPrRcr
Mqu6JCzDpmsBhkAljlW5ZYYLBi+8GpbQh6YjCyvG9lY5YGFk3HvcFyr9y6EO8xkevwOnDbC/IftQ
w8dsyKWG/VD9R5w+23gP89FaIOL6v9TtM/KDWkXb7bLix3tRJmvmxI7UuIW2ZQvFm8sYB2IRx+2K
Bnx8HJ1TX7bmgSG7+J62oodfl48dg/Adcwo9JpZqgJBK6MBKyfFpAHz4Xkuk/rnZmUcz9cBFLHxh
dthcutRFAkeF020KkVeP0BihVxbUX3f3U+Z92pTojCJZsVrR9Af6iujaNuub0sbPT/4kSz3dM7pW
dBbx6LwhQvGJdn5vT2X4On9m9C3FHU3M3kU8CamI3IjVTJcjLeyU0+x9FV2BmsK5HWXBNruUDeXl
pto19BbkNbAYbXouIgsPMHuNgaM571aFai00HieMF8TXez0B44xROIu49cmkgWuq83+gEkMK2X9Q
z/+PPonDNZDUrHDY9o3Bvryg0dvjc+j4ugpXwDkHur6AqgHGs1/ImdJIcRAp8fU+Q/83K93KVrjA
e7YESlAhi4d7lPI6vQtQ13J3VHSkRIPTwJh7FQCkvYstC6p0DeDoVhoCTNERrpIeX5p/dFIB9pus
G+5vTqcKP5B1BwXm0nQW8+ZCA7BuldlKpXpQAD0oaQ0yQe7WWXPWPXTpNKmD9nswbtk4mGsyX2Jq
gaTkucWITx+FKOek2yStAvjwlWXwhLjaDBosBxjEuORJNFz0IZBc35K8hnsYJNGBpfpZPrv1yLNe
D2ogO4o/ZYqQP3yEjG6mi8Wib/lz0n/r8jWnkK6iAP73vZ5DSEBEFsbXcLsPzRoxY7z+D7BGpRSA
RYFCwOYcKhoAIbbjpslgOBjhuGfaaqCnm8yP6k1cWt2f0OsJcDmj9jTicDtnUKPeYmB0VAqBkDqD
aBYDGuz6A7xYn3JerjNJLn85h94Y5jwGzn5agoooGW7k2PaDxlv20/j63WqIPAHx3ZwtF1X3goJs
LN0vttAZu8R80GLqnhnVecR8kb21lCe3XdN/KaU7JnjG6F6D6eRz0xWu+uauHC9AY1dNS78wozdC
Alv6kJ0uz6pYALSzjf3ca3dEQ8/4UTzmoV5jZETgKXFk7ys+Hy+55gysWiDWxN4pDeLRW2RqgO9l
m6mVVwNTrK2UJQp+QHtbrurNGi6Q3f0ORGzUfZ4AmLdSE2NaorSACQjUyfgm026GFeb+ViriGpbl
g9cw4Zdh4BNUu56/g81m+uMJN70ovVOdlQQUxbSfixpYKFUKHAZYQveF/GvLuClciAWeibXCP3YI
yRTfaT6Y4tzpv0FpAk9mNitmUBRvvN1S/63Bmqgnu3dIEnoBQj2ikkT6N/QIfVpZOzobqzC3TNej
cp/E5UMCI2Qac3XlQ7qUHDFvqkJmHd9gIAs5zenyAzFRknboumBDO9hwBXnZryxYogRIi625OVcu
2cCMSL11rmJM8zsxL2owiRfBGx1YKq5p82dMdNU4XILm+bW0miqAicXYRZk4GHWPQVRBEICQfwXD
pDh6Q3G1h/3O4wTGsPuZ6YFCZCJPFXIYfhAADlJY/AH3Ogcq4Ka0hY5WNpBjOb+ZJGHw+ukkN5R9
Ui1xqEcqspP7B2crwV7KOYVh2fzHWvd3O7hc0Y01AuQqrTWVVY6uBkL5ukc5Ho5TKHSlKVZpGyuM
xYn51SmHObkMKOnFlfGjLyjbdxzG4dLq4ICGfOMtswix2sRrS2wVOBLRcr7F1lFl1QEgQpA0hN9V
gYTU8O2O0Boy9rzb/5QXp1avxnu2c++uj3nCo42R0U9BoKY9IpV/pSd95ivA5QYmfactcoDNfImy
2A6jlx4kLbexQbwW+Z391Vjmwa5LrH6jaWO/jZ2UWbf9HIP5pv+wGlFy925MpugqPfdTTC7mg2+9
gUrjBR1OOJlRkjWHf45ESXan6xHWF083VphWkY1f+1hLdlYquwBDxkDDfj5CnGYYfF8ot/kTwLQu
FcvhNeuaferuUxAwydxmvqMWRwngfVTFplZIvBxO6yNSZO5gdHWCW3+CFtb+1sMb++NFcnXhCpf+
QEyRzwmEh8wne6p79BtZ1AqQQEUOaqCwczrOHIKXaZ7Qim6zGrR6NRM2uy8f7hscHsuhosPOea+j
Hkiw4C+vqaJBV9nExBmXFlsLq8QilBGZi+Y8er5+xyAggj9eIX61M66eEyo/tBeZM2QWLUWEmBs3
zMOe3P2gjN4eYtyUA4vWA0oyaE/G52UKS++UcnNjJR7/GxdgsVYJ5Hh8RXZ66iGn5fxmwY+TIHzB
5+9tDwv9sgXVsxLXjxlK0Ey0HrFIvpCXaKLR7eRs/87ZMFQgFJrRw89gZNVzxBJBcrLpKyebmwUW
2V5/0nO2qhM5IgbD1oQYeESLi4SW2+xBbNzM4AsNUv/S/6sUkeN32noN6/ITXjtYty9MMdcQzIOZ
6kyUnHGpB35LLoNeSXMtuLANHj5YJyRDzs20authN53MREDVd5QJ6t+r0V3mcsI1tY0VNAOSKrqK
lcRGTPQEGwydn77kcFdXEx3Z5BGNqe37hxNG10fkdKaUqx4tVIc7fYaQrbsbldFctqil0KD6+OBU
0M/3upP2WXnR70wDzyoRUfHfdVWqdeCNS8V+++jAdGpK4wl9FVnMAcSdH3VDqcX6gxtEN/dTcMJf
3JFY2KElS02pmZ4EKCC3qzKd4zAN5/oeBz0s67PYNNal0jrq+NoT4RQc5anqHVCxC9GoB/M2LuMf
9JVqV3qC9u7DcttBt/Mr2x5aE5ScrKJxHQcKKraBBw5jBdYwTnGjCRSVjcHk/tbsLUFjY6cOC2Yz
lBzLrW1f9ycTV0p3RchfAfRjV/kNhbtVeQF4uRIDwr52YvCIr/T2t2luU3MBkoObc5o+B6G2p4U3
C4+oq5Ij7/1tFEXlSMtwuCOR00hwr50tKdPY1fdQ0m5yZy+7ARwsItVmXr1K86GNeU/o62Hv40OJ
9t0DF1whcOfv+N49SNoMTf/JtneYfVjo4lcWz81OWkCXJETbVLbMr/G2vpqY3BwK7LVC+EZiEcjl
XxAJyvweYIfXeZvQv8xlolGvYMI7nh8QSMU4KTYPdwVGipILhNi93KEGDqqT+c2aQ4HD44wouv7R
Bt0ikAffWM2IGYps6ZKWiq4tWmXAhfVPaocXSfnSDJcScJdlcV/sqIN943G+K6kwyrQLIPc/0OUj
75TmEFmEmKJg960pw5gt5B95oA7vPOuQpHa+vE5HL6nPjlK6Mggx2dXpMWFHTIIboqfkUouIiuyc
wlI14tyYG0j5XyBO9NbMsC5FdXckhbA8wFeOoal7Mzj3AyUHu72CWuC9gSt4WbktwLajN0AEo7Q/
PTdlF8tP7AqoaXCcrmL69I99MDLD0ERg7k/dtcu8p+tkEsJcJxjXAsr7PFXj458IOhGLr8cutxJG
uaoA419BOFvIoTur/UGH56rm3iGttyKs8KZUQBPiEQdhUkVpE2ENq6EIIzV1NYKQVuYec8hSeXyN
CfZLlRhp40Z/1kOl29XhTjA+0tBvoEQzuKZOjTmjcTNinSV/3UdvYpKqVEVHxO86rsV4FHWrKhuM
GyQhaHpjXfhmtNlEVWJ5AX3LN+5k6Y65/deEa2UyTMyX4dqBtMydIP6Y1GvfDVCNDd+RHmkW6uIG
g42gIO/2/jvbXIJDCTkdp90NzzofQWJbjDCN+Sdhl5ZXHIEnw1yIZ4qboqs1lZW24JtRATb67duD
OhhCBDLSXtXBhbXipvd7+3L6ZFEGzDNjVsf+wqDIh9RToP4Jy3cpX/R5U9lGFG2S13PSiIRetVqX
QvcWT5WkZH4rtluA0cZvyd3USHIBCBb07E7H18sbU7rNWylBWO+rgDKrR7OAnNzFRgjMaxfB1GzP
VVrMGD0uOGKf/egmGxDnGFjgrvzUwqe+SjiV8gv55iFAhkax7S+Bfch6QVp4e3vCm6IaqrbQXjqM
r5Lf3INuVzDFnWjyS9rWV2sIu9gW8F496TgTgLUNWqKB9Q9mcqbwF3LkjelHIihH/7wXzPDS/TkI
eJkqbKFHUYCaLXYNrx682yK/tkF9k85GNp0qTHAwPfn20KVjIm1CObQRJ8YX6oFwXde2TFBgQfMy
F6V+5KH23aECEmZXwH44qG+6BReq3vyATwLK+9Uyo3s0w46HpgCZW7J7WPhkpeQV7PwHxR2IhM6b
ANi5f7N0m8eNofJGyWjOZETgJcFlL8HP2pq59HsH5NQEt7fYg8nWq6r5eKq03ZMsI+HgyowseivY
XF78DUWs3Kxc3xic2mQ5VY3SLXPlFR9H2d79nE1AYlXDsBLR8nF/p5xH+0yvifGp8EEIFRjlHV49
qeCcjRDujDi1ezMm6Qq04VadG+iODI975n9LWmsVRDqOdQqlqEuIsP1I/NzNqBdUPBaSjDv1Mpqo
vlYEvSRWivqOmoXOohGLMEOS3ZVnl6nYqFAGP1+3mn3ggwB4Ig64m40F9qceNnLthGSv4NRAsFGt
R/ahrk1RRe1q24TlqVmAK4Ojfgy6e7XlUpf9yIxX3xukwdhPxL54RWhYTcpSDwIzh8+Ka1bRxcqZ
vImxs1BhOctdAE4MKQ1TrD3Iwf7zZVi/sRaIeYqqwZKuIUAJ7ZOJgfq3jBfRvShtchDVlkvJdgRf
XeKRY+xQfZhaQrtTiMQIyYMi9eoHmAqOxprEiHyKs9h0ethgYx9hUlNpCdReK/7jxry4bQ8hlrxQ
Da69wK4xmWI7tclwuVrtCN/M4aKWSabFKGSf/7yNDn3rrL9UOKV7vgR43X8YZsqpQ65hx5CML1Q3
QfLlehUNozJpGl55cA0guQ24/U9qP2f7/9Lr5oiIxx0lQUvsQyKK3S+IbmG7kZ9iBT1DQsj9hr6k
AUrk6aSqiz/30qQXRNUtrPgd3e6EHLtRHPEmXw7EwryInPKdLFO5rDbeu4fKn8SL6HukvoVGvp2R
8CqYrMCOUtKhRdj2yxlWYicem3IPYWTaZ63x4z8AHWXkt7lIeMMwvhfsiyQGAP7g6lAGUXGJPn/V
THcBaUZC1k6YBnUTI+DIOWa6EkV5xJMrkWLmxiCLMLnl4ePxjxUeZsrOVFO/jnjpG1/CkRUOPkOl
0AdEsoIL3fF24sSArcNwzPHrTLAE9pL3q6IcQtll+LC35tu8MFqusdLMQ9/ipgmhE2cLVMOyvf/6
pIPbAH95jZ33zcnywtYQB3a6eSpS0ndQkRoFLXdbDzXr5YcFAfAf6nIW8k465K6IcuafXliqtgA0
GLeEJOwdkkv1uR1HUoWvRW7jQD3lBrJEHoCmYyv2YcXb3lMsyzaWIoP1Eg6+Il+/4mcINgJVfucr
oxSUL2rj0BVRjZyT23nwrvonQ1YmxQ0Q1n5IbrsX9eXWq9NqBoXBwkqvJjjNiZ0KZyHgUj40LrZr
x/8Rj/7V/x6xMx4ZPfo69Qv87a2Cywvpq/afGijMw7Z7ko2AuVeY4+BJPJqGVh3RMK/PA5sqgTHM
Jjqs9uEXv+kFIb2pn8zaYOIvSn9z1FchsQ4/v3yJ9xuZCMxqeIA9NRXGBrSsJch9wgeB5ZU9vWAi
ykzXi1zxEqzbUXAy32N3lP9iZDpcM456OlvDti+tiiJ8J5NNL2Px4/y3TMtwuMgGhijhXkzerGpc
i2Y1YiyzkqwflBlvlRWgLzf1UAVceBto54GW/xbeYCvj0awkmJYgTDEboQeu6mCJGWYT8qtrjGdj
SZWmHlCYaJ1BHBtQTpbeIP4AUhAnHP9TH9QgaKIm8incBrMI+gcuhtnd/5ZU5HgX8UHLeD5bF3Hr
V++fLCv4G+YsJFjvm+/XXr6TEwWDOx8ba/IO+YQfJbER7btqDnjilYHGDaB7SZyciUaCats7YwnK
wIS2I32JnWYONwvp+e8VGTWoClTG1CN2RJtmIwhl44RBmNYJtWjKpvMFFGMKi6L2PkbPiCaE+x0v
NRXp5EtxplSAKSyR9eC7RjqQqCKVJPJWTK211lE9Kna99yCnJg7a2x/rwQdGGrE+/1/+5EY0HS7m
b4ZBFVKYQ4GkuDsLvsIodNdIhVxm26I/EvTxa8aXoD1WfkXI0BHhZW76Ed5pD4qLEzFa9VwQbpPD
jNzzdMsqJi/PT2ar8SyXId5A6UQlN8Lj0QOrLi+o03U5Oh9OJhcTuyAArCaNIrTAgQRCitVShxTH
9JnXr0U/25CTOf0eAAXMtCXwUF/Dxk77AHz8rT8hPxG4jrYe4hkDKm79xMJBKCBCudElqwuWERTY
qRxw9x2ueNw2WFs8ZyQgZdGUH1GGigjzU78ipii20bL28Yx0dj/XHHNANHCoCEsGPfcYvLQexmVw
Iv26P/V+r6N+Q0XEIRMTeLfEtUNd3ReNru9lcW3kip0NTP9oCXzM76KgWk/tPmozxxCIyCoV2QfN
HMzktf1HVznHP9FSzbzh0nTpQG8jrwKvDq/R5sCYg/O04R4GQEM9a26dFJPWDFuuMQoBtvgSzBHE
C1kaOygdyx+7My2rMT5Ue58/53iMVWsFhvad/4xZJf38kM4B1XOTb9za1XsG3w/D1q4NcQ2nbETn
tExC9DXgiTDV70UuvJKZCXQuySIYv9v22gnsP6Ns2IpxZuFnWzluifyUFGxW3OD/XytGFeGD5ZsI
5FUVEXZuDRrfaIgNp5Mj5F8pR7Xmnlj5HEHn6EfbB6/ALZznJwLcaXje8H0E5Knflvbf+ha1auWF
UYjH4IAAOKC0l4ZI9CwMLuKtj9ijiOiF4X8zu5M9VS6PCQ0ylsxLVH0F56ziMjA9H3zVm0gpOLs6
IaOdQcTd+S7aLgT8oksVPPsCU3M8kBulLc9eKEp+4MIpKjtR04Z9M1+FJ2SCOqmyKUKCC4s0MDrK
EyK5wXYog7n4/OVn7Qa972PXsPNTv5ainsWeiF7LDuMTMbaaL+sDV3XigtoRoUAH6sxIhpsKRst/
AhfvD1PkWOJqw7zCCNDgL6NWevp7c4l2JOeUVUhbQHo235KJHu+BIKKPJAwxqPbGVo9SaFevZkLH
soOYSbq3RVJmxHVvP8LBTC4ZFiI5vgS1XwCgq0aUq/sTYVllFL0snU9kXQJEL0yNQFJcJiYJs3w6
Ik17BsXtNxtAAC+AgurO1v9hXlRtQum6Me8ZrwDx/GdkToc+YhQZ8JM7Pxg2TdzDe2vnLRmkH5ao
51kU1GxWLUiG4+n0G5Z7HunOEvXskSY7Gfjz1VejjlrxFk+OQYjx6qnRDjN0oRt1KRh7TvvV/B4p
PRua0lPR23dxcIpKjJQ8XrO4GmYeQmo2SFz/i9M+tY8CO2fm4zajRcpKUAa/Rdqzx3Uw8qSS4J/C
AhQ65FvxyUDXUlHIMaBMsIJultgizdbOYtQKgiVI6vYIA7Q7YFyqwDwHFJfyxh4rgqKQZTidaN9J
/BEmiQitzNyeoXGg/ILZGkR1dEhdYYQqpe4kpx3ILB9nLVhidsBkOGNl4q/fNYFe9i2YyZt8t9Hl
rpWS0/CcghQrk0w4ZeNAK+ZVPcb4xtmMlvmXeP1gGoYdvAK5Dj2bJlp31lHkyVxspfoXxcQ5b6rq
OJDZqaSaC2/chfmxtyedhKpIeq8k+Bq/voZncTQyrP/4/g0Q/QIyl7Juszxlsu2HmD8jfGNyLl/t
X0IuwJCZTKIMxcZ9YGz/tNUC6GGGUdBRBT35upHGPn9rD9siFV8JS+O6XJetGP2YddZruBkMX8/y
RiR9uXsEL5+nF1NoJlRHgRkgc7sGA+1/NbF/YSruIgNHys2Ryk3v9QieZxm/qIpmf8QR2P4GlIRl
CnVAa/v0Zc9T54C/WGDL/IQ+nX+VpZIX4ojyCaNYo5MdjI8Lo+nfYJ7gizMdUun0QxGTb1K32jqi
Sv6easNcyzBxUkEmpj1Sa2F4LMfQeEz9DZDUukOQlIdAGPxgqV2k3B2JZTh135ezwHjiTAFL8qO7
RJ2UdbyPJP9WZnaVDlcYfOGVRQw38t3RSPytZodjOYU8e/HqTBVjlJIDHRjYg3Yi0x9OItYw3zxI
SCn7uk5+QhgxvSoaa/21JPYRgRqH7yw+q/KmVGLc1sCwMKfPkH317Sv/BWq9EckB3YHqiMT+LDh/
MLJoQm3ErEZuxJllMXsMPUqAysW3aq6y9b3j0O9+tmlGN17vL2e+OizlV3grGlfz3CbenpOYh7f8
te6tyMW7Mrp4iAO2TKQ4vYCeplbvxR1tqVJeelp3ear5Ds28H7wsG3Na5XTfVVK5yhrZJNBWyPVT
2yI3KAkvHC2hwcZzDVX+z/mGEciNCZLYDZTHB6zkm7GJiYR9WxC0y0XFM6tDegEOOhEWGuULILxI
8WcZpovqo9nm5PnGlFlOOVeFV0CTKdeRtrHIokByXKP2VR+WN4g2ISnjG6MlkvAxO9bdWk8ztw9u
sfJrC37uIREmvT6K6M0o0yk+SDakOP0B0K7EchcFI3PeY0iV09s7qFtdKCExQTJAF63OfdSevMXP
5GYwhJCV3mx0XKEFxOV85m2zVQyMZhQ4sIzuCyqLT6Pv61PQ/8r8E4H21Ke+0RSh1dpw3yydWH1R
s7SdIJPlMIGsOobKSQp589BEOmL8Fs+lm3RSRT7g2oLhFPSgrubMvpFr0W5WJpt5jG39K62xh/Gy
NNQKcddyoV2YrML3BgjtEewfI40YoSQGZ5h6pXnm3oDa132vGfYrZNEzVHT4vyFiiDT2IpAf/XQY
Zamhit72J6TfrGzImppNCGjjE4RU96DE5n2yVrstS9sw1vSGmhmgU2Xy5uxnpeUuylmibrk9TaGz
xKNzR/nF8zGdfi1tQ2gVa3PacYvF2yYWPR7ttRr2lQJU7D9D19jO08cokifZRznS2XPN1T2DLfBa
lzovCqhLIg643QGd6DZdgEq+3DpUbHTUSn4Iq+hhBH+otZgR6jc0FjAIYnd1i5fPiklW2jU0TU/5
Innao+mWGvdZQPTaxugJVrpQkMiFFeZk3iwY9sBJHJmRatsP8Y/BY0iyBsVqSCtuFbs//eCLg3BC
SkXXj3JHP365OiB+wCaBiPupbQsr5bl2bIG2V2Z3zwPNT1X8LnSHFQehIwkFSHTXe2SEHsisIml7
/nxvl7ZF7lcSeer/FDyUropU1NlImbf24kS2Pk00eeRgFQusxXecFnXTfFP/7Vuoy9PBC8HyzNxJ
cUNzmyklW9VGtfPFl+q5PuenJS4I3AViJepSOZ08gtT+/jTBFUb0slPcKVWcb69C2cP1iVZthMd8
JRqe9cLdlgaM2LzmLdMuFQ31KkyzIjlMV8wiaAJhsG/fax43O2NbXxZtDeuil5LUHPO21xENjGBM
D62JKszizdT66Ro8ZW1oK5G8Nsv9rkDRqBGR0EaAZaUZooDhOxWJLinGmr23IJFBVX7UEVWf+e8e
xgCUCXnH3c0lOpGd7sxedOU7kaEtJq4HV4aQcICd8LAuSp/nYkTh1YfuoGbTjTEPR95TPZerNbNh
9hg2ytVaa9OTGERBjnoUlP+IlKJInON13XNmCpUi9JtAzZyCoV1y4LHppaS05n8zuIdHHfh8PY/p
SqeZENlNryJnO619I5XZv+SWK8dFsUOp44ZhKInpsQqXHE25IdI4Ctfl6tevbIwm+h+voXebXQbv
tpN4NuaEvU/pvx8+F0AmnCOw+csvP7/ACvvQIch/GwbpvhgTzM6ByzBzLcsNqC9dQS/536zHBp1p
T/gJZlOZmWfiJT8qsD6WVTpK9idMR11mpvokSFYyJqFs6X+YFY+i5oKbcxWQeYUwz3rn6HLctcju
PHSWfqKTOG4Ry46A8c0CNZx6t2zmrb7D9jMMRWEjjcsV2XoPApMxuBw6G+oSgrLavfDAv5zb3vH5
+kWaVphtHSyudPIq+KHhY89kR7kRjrmuQgVBla3EwFGKIPjqCtSG5jBQJRrGw6W/bh4ti+8Y4BEw
n4ChZHxu29hvB37/V0e4udbc1/LLLXy2efahWz5RsgnXgjacD5x+lE1irEa+K7MGLDEWMJ02iQ80
iaXq2OeSJYob+FuZLXQ1DoOz04fkQT7KzWJWeW1/7WwjU3PaZZkSXZMDdjuIM7F/eVKQYRhL3bWZ
DZAq81hT4m61VQmmK5J5jjA/6KpIGXhj0athy1Oze64Z9+W4663/OnhXoztikTOqA6dUpmZ/u+R9
Wuo8kEpe7wdfaebwV1eE5Xl3OiMMcC1uGn5lkvi7TMIH4qGNPsFuouJdml2Q45V/nkacvPLCu9WL
vtkagGO8iExrI9hFrWpGGPsrygMSSj8QznPW/KWEUQh88u1mzEqyUv78oy4i9rjCCHquXlrb3kNu
k32yZSHKkZYGDmPIt2yesp3psmr2NX7fSblkb3buv7fCG7VbWCzt4m8EQbAEoe2jtKLNW1ZfvD/S
gXcw5USUsW0zzvLkhBAsyvmBd0kWSjBTL33zeLEW//5fJXqJDeY/yfKY7CUwJDBF/Jx2IjJX4AOM
JpCfk+tpu4MaPwzeNVJ+Knwns8I+IOJlk0ry9Ktq9Q4dVwCe5IpB/xBCOJEPK3me4okYOR9La3DK
uFlAg5J+mjtW3wK+Ot9sevo9D36P5GtVW7jH4mJngcfynG3Kpul6E56v3K2LT54Mln6ofT4c5Rpb
4FxkMOYglCztjkMnza2rzrG5EEH1tR7zbNpMvD6m21uKQupgt77GExzsMeuWplu9pIMZbuhTKNSt
/4/wfpCGtRKVdZPxeO++SphF0RNK+miNIH0Xq4nUphW4zyNa3EFdkxxxsIFdO5apydsSQ5AxC7K4
v2hG1ZNhjzltkDmApmBXxAeElmnirZkPr3HDD37i72SpiRwGRBo0e2ELQznogMgx9P3MZ0S8UNkZ
XcWBAS/3V6IwySTSL4CVO0briXBMlHtB5ZWX0LB0y+2RHomBU1ewNfoDhX5R7EUYIijmBCkHnMG0
rArDChfs9w2XskDp2/guneg3ruyqr39UktscI/7d3W/e3eqf9LXydLyZV5NtYSuQnkEdxSK5jjnM
+JG99MjGnzmGo9Rg8xJOyV/1JcCuJQ1pUO3ulMzqZi5N7QNZxO4esLmeUxRnH7jCjJCUCuVN297j
ElwO1MeOuo8gfGPzOpkOE0TTHU4BgDdtMSbewvTOPsJwMvLIt9OaUzlfpJG0QzfDjh8ufGVbgo5m
MYGnyCBq2asHw7yKwQaNYxyfDheBsts1hDUl2RUmBMmOSMz6qunmgTv0Jp4AbmWlDlkZD/UPQT07
NeNTxB8h/07P/o6MvsiYL/zDNsnHoXjaEPp6Kb0Omje9GvzTSIwIe+b6E1YbeA0Dhwd92nYSRxfz
gTPCilkIQl/q/A90y1otlHkt4OmwhdqFrldZWVKRwurIX3LEAqE+jLNmIFkyqIIEBpLa/bGjHK9L
sLDyPV1H245EXTeEfFywwKWfTZmAX0dRI1+q74EFo+Oe8c3+EH5A2l06PlKS23RWETxg55l1FGA4
QnZBbvMIDQ/6OVfVTK7hYry38L3JmcoxKnoeh+Gf3OYd1/ZouO2Z0fm0GCsuhaNmbbP5uibG4KUd
Qa6rB+8S87FLNp5q+GAQjoHc2Z3yCRgj4KGLBnhIHlX/AsNl3wW3H4/m2ouukOHbN23ksOoGBtyA
+Tm0N26WXGCI5+lg793RLO9XI6ux3nuq7lS6dcF9PXdtfk6/xU4M2sDFGQ9/lliCnGlKOLMIa0sV
fh5d/Sdz6xIlr5cvxRVRrUw9j/mHZqjyHfjS3JjtbmMrF+dMH0+ylpB2INbVX2KL6nrtuOL1dbV+
nCigNuw7mizyJZwfhj5Y9deEM+O70pJk0+L8LfdAEYk8fg39YTN99+2IgHTUypxiz3KPAJFLAnY8
EoxX1FRF7opwvaPkyu8ADuDzLRG0U9EKDPTg+1gLRBTlMp/ZSImXFzlVuoweUUd7DLn/H9lnZGyL
C7/VaVyAfle2jgKELegBWZ9oHBUCYUMTGCNXgqmlpbqkZvvOhfWmcS75wwEEcQma4DRfAR4mfN7r
Xv/nnqRC9+DcPOkuvYEFoCkKO3NnoxC1NZ7Tvq8O/KNrjL5LDfFBcnxrW7mAJtKgismoOtlxORu9
VLsPtOXjHWDbaVV+uTDxn7SxCPWOR/4m8B8YJ4nMd9CBE4Q+rnZyrkOn/j3sRKXjUQMrfYppr6j9
mOE9KwOx/TT5wbjrMl0QMM3jSwSqiomzvQ12Kmf+/91xcPFH/P6zyJEES6Agc/3uNVvWcsmnrJaT
u9SgSCPDaOslBEnV2jsWDF5KSRb/1q7vDytwhrAuEvedqjPZo7VfPoSZgZRHZSjwsoecJFlGn3TF
Ocz+jS+b9LDc0DGsTyUTqYX47u63NBWGOixT5Wxx9nQlygb7KNu+djErffqN7dHY/L5wlmI3ff0x
W/KwUofGcMgcPQtNaTuqxwE0IzaftzUfFd8oTDOK9IxK63ERViFNQmKf7FZ5GVxvcwKrLITF1S/n
Z3w0wCeyUQjDV4dQxQ1oTOVG9jiDm8aXh5EmWY+lkmVkWC9oeAoCbtgSx4ggTrViyGfMlRaV2rW8
bnUVGyseXlBDijNyT9f9dE2hs7CGutuKR8e2Q5O4kw5HJadZc/30NPDFaINxE1gn410S0SyhJdWM
UsE3n4inxDpguK4uPCcdw/wlt3+Ax2W355lZcWmVHm3UgQtW86NKeYITyh9wrF60Y9mWFiHmphTL
EereSW2PnglxMeAvYTdeBa9g6HGUV1uOJMQhSfgsT0N/1tEPh7Z+n8mLH9ECX/uuFRbxHRM9jYIL
eP1RYiXtUIpiROuSrwKJ1SBMdgUmm3yW83Qd5u9f1OG3m9w9aLxQFbtHHodDYhfGvla9b7Strc+5
rQBZm8qYGN9OC0mX4S1IJDTGRu/HVozVkuaOIV+G8eKHhYTACiuqpLgCUMCLGMntqGe1/jKtj+Jl
ad6aNiyCg3DCfMgHNmD1Nw9HWXvYH0U9ShLNKrQp3AvyjSO1CGclM092BS5GJ0p1YH0aoqdiUL8/
RYpT6XJ2KNaldS1gbJn2USWJv2pwyCw35y2Pp4+B1rf+ad6DaobK0UMQzj/H0LYkvdJXqouuhveG
oRUTq+Np3fFM5Q5tW1csC7C9kaQhzorcZ4TOvV4kvQRAPnocieObO0e5+fPD8PFgrhwBRikX13CB
YqdeLlpQnGfckptleu5Ffcs6ydZ6VJsAtOWzcOba+leY1Jr3o57rk8szruoNP/MRM3SwqlzbxeeJ
GDMwD0IyxxCppctXkUJ/hew+c8nwHaJ4mW6sbvtXgAfMDpI0WXoQeH2eIzyefF1Hl13rIqJGapws
GlzCOsXruWBEHkyMBRhZE/35B8CmjPW5NQj+zyTgfpart/Nlq7vdkVNDcSj8puHZ2KuViTfOd465
Fy7+qSruN4xRYxKGT/59+LOO8FrUq7kaWacwNWt1H66ZQi1kk1zv9Lk8UoHwuShkofzUHeeidNCu
njgdMNm+lmtv9zEIY0jzswKzwKKnI+HpE71NbJbAV3NT+MoNtzt7QVZSlzci1ZMHWQ0DPNHHutDQ
+0INOl9cXxbI8FCInO9YJ+Sllf+ILb/Md0w2unzgZWaKwS6Jb3zp+xcZ1HntbBq5c6tjrZ5Wdm4a
ED8fSUxqOqU6yk9WezSIm6clgkpsEoJEY/cFMEZy7LYwMPshTe5buUi8vTGqI3fvwbEzMn1fswds
ZIscdn0KjQpdY+cCWTUbwnrSgGPnV8Wuj7SVjgSRAQ5VGP0w8+8Au0p85BznsVk3DK1C7WxO+BPW
sh45Lk8irH+kbyi0CyUCiIW9p3PNGPtS7U35m21ZpdTNrJOCU4XEuB7Okw8OL4y3a84q85V2PYuh
jttzEt1QNH4oNdvvTTKdi5N1WJxHoqZH1GTHVwgC8ldoo00YbC/x8iHreGmfPvyBzjbDQJnt/lBt
D+xSkL7tu3TVRRkXMyC3wsv1eA7jzy8cRJJbtWAzshpxNjyJTu5iuLblnlPR71wHGQRjVqKVqvzl
Tx57BJzUj51Obz83XxZm9wQhdxDYUYiuJtVgwCIUo+8WoF6r0ObaUPPgYfpU9T20cj1Larfxf2EB
kEzXSyhs+sAZW6egzpt/iymGqzxpaNiSgY2nqObtYJ9xH8rIR1JWcchkmcOqbR176ZjFtU+LJrTR
31tY6B2Ybz2qAOLmtEtaGCJOFjZH7Lq96N8SxH2Ah3agA9PdSOxTKzZuVn+3oZCTBQm+CE1b2gFA
fk4cQYvnSH70c5fuzL9vNd1J90wkjOdReMotNaMonTFgRhhV3hP85TG2VCtKO6oxzpC9mjLkBA8o
9T0m1oR6Qwz4h8pMsOmnzFQFt3b1teDp2lauM9AJKA+MvZdP1fVxPmowVGshemBHyOhWoVWfsyRU
lkMasfkoRSyfH7O1SnzJg1dfit61Ze2LarYr3dAyAmYLtq0GAI9qVQC1eKFPM0Iu5c8+z8tEAEl0
jQTyfF282PX5va3tEaNe2vNX3yTRqwhCtJqgnvfRia6RKgdCpp9KOzGv6nNOxoe3Oyg1FXAB51PB
T4eCE04IIGxBKwonN9EFEtmtsx94ilWqRfivn/tJezk0trcYFjYs7gQu6VQ1UCFXtVnM4srLkZog
8D7lojBbyYYhiwTSp7iRml8tD3Oia0fJflzVkNPqvvVoYNmGTlRoxR2rIekEkbRCnsofUtLD4Kty
SdwyPDjcRT1HciPyJQ6oOT3KeGKtHYHgWqzWDQgEwBaSqYxYOG0hZIcaTMRgXUKqTtJ6M33C/VZb
DqDRM7yqW2zAoR6JRqxGaVybLln1Ft633BNlRu6MXr7/gopbiyH7bl2l1/aHFndMiqLo4W9Ymtgi
8/WduZSxDXmXOfvAGlt3Ysl3GjzJyXAv5UXp7UrXhcM4tt0aDaIxbD3la6ABzPnF0lOp3U5MSSpf
QTJOHFH7xby/6s3WOGs4IyL0+K9ayXJg07+Ee1ErVTZn76VhYGMiT/PWNDXpVHo8hLv/NCkw42UO
VgsN5JmK1aHcLxH6WrOAop4Nplbbqpe4jSvjxkD/E8p58xf0fo9HOPK/2QWY56XPgmHcUZTS6J9B
Qhc/oSqZIIvvLTpHfMEd5vDCbv3UHZN8bOBgk+bx6PMP8Q431UGhqh6sRpaKlap7SIib/J9epDla
GJ9xIDmMP5lvsPlxo3BJhfW6xvWxjGUBuswzBV5lxKIl9liYKxLw5A3sTBC+jGWRun4GjtkVx61Y
P1W01sLBttwJOtyudbX0RPex7eyPP058C9KCDfnpCgQIuUZ6qV4bAseKwZbYfa4cOve27niWoFFo
41etLgkU9zJuocSM7tnRQ+32eLI7BAc5NUlF7LLFJ+2r87yKT1AqjMUEe7xGP5qnUUOWfkFx0Kzx
70PrBbtXVI3nYcSMrvFnklT4ZO8mMdoJJtOHZrVIgIUSsTewo19A9VFYQxFd105diO/G1mWFOalg
mjfNR5fHW/dWQgf/Ed85mg/Nag6WBxClHQo0ToW53w68oxxp9cRi/G262wu/8lsdbV+A+KDZ1kfn
GVAG1sl00aJcx1h9fOpJQ2fN8HXVHGTUUFD6fI3JDR3yhw5D1jx92fjTjlvVKh31Dc2Ao5S5Pwvh
54DvtFyonh8jnArAn3nz8yARAIywpCeHZ/TznRqeL3qH0uDpJFRYvo+oDlEA2qcs74GoYL9ebfRV
Wn8nssUnLtR1v2nBCPjHvJpH/UwemrjRSwq7L83Gy8V15+Y4UozgTfJp/pyYrENLVgerkpVx8iJF
N9F1d9yno4Ru1Zjy9qLcCYiQz6Kq/FN40w5mp1bwZO23YMqfn4zujCekEVzT8q1d6fRGcJl9MPQS
bzWaAJi2LRBSFgS9iRMKwPk7/hHdLoNrtTDgr1sLGUqZAj79cSdk8Hvt+ddHcAlNkUCQoYPR4EI3
sPWHfXRKiRQxd3UGVxL3zKpmWH3Aj5g16ZStPA7YA+qVosWxCITtznvFKJVtC6QPu3jytGY2D9DI
GF3RQxH7B/Q4nARmLQsio6xhSRIqwfjZVD4d0xcSKXZXogKG0v/IeDCdb+qaGQLZDzALC/i0Wrbn
bumTbRVO0AZ3q/dc2HR3JrkXxBYVgpXgWw69Q5Yb5teFytxGxNNgESooL9L8Ay4S8PV/0JARnZlf
ZIPVxc5dpOEpTxCKLTWBc223BGG0x9cc4HXXfGWRi/w0hJ+f+R6/gUIaHK8/5w0G7T/zfEDaJ1bR
mLtE+fNbyHIURx3HeKndMG5HNoecn33A1WyxW/D/rf0xQz2iGpTujtzuEJQ2BC9LBk/mJOvfOBY+
681QBQmcTJB3QSBgHXKmNjWgeKmtUQqQZPH27hMMgF3jKOJOzQa9mKxtSpkb5Ij7JXVh826f4rNT
5a2nchhvJoZ6wNHExmj1aBtYT1O+JTeplM2m/SdaJ1h3PXOrt7RsjVNzQ6rfbQXoacS7wDJdC/Tc
qNiiaQ5IVBcVWFtT2lQYSkUUzkb3dY4O+G1pIDaM6KdZveYStVv+8ANLnjO9Nd5tJ4PnXq+AkVkk
8bP8n6h2jkls8iuNM+1ENNjfB6WpGgd9B4qaqFckvMF+b0MQkXSFexXuk9A5pqNMKBt2WyQkXSB2
mvaqLU/5H5yZ94kNNCTF+ODGlT60KvgGmb1nuJrFIaaQPcYJy8mLnMzXIJtHzTcprf857x5DHCt1
kAuY2KYgVn2Ide26W7ls5Hul/z1BZBw8vYv8LPz0+BybvHiC/2WMX60vyxA9e9UKzJwttgZF9vp3
m6u7GvuvPBoGRHig5vzst5XtFchm6w+zpMzplEhgYUHLctLJRIJvuP1w0OfMADAiwrusEsSVInKT
P+aANSF7MpEi7R8ifYrwsYvLb5/ZTHg2pDe6eVAV/9jZz0EDq0sFpsLnBCm6cbmasOn5QZXQ6l79
mzlIFtXOFZ0m3rhof5qkZebY4FmZzfMHfh9kac7OC1Xp7S4Q6V8t/S22ae3zm3kjAcHz0Bp+X0FD
jI0UipKMnqQIKeJCrNz645EvgmYn3Ln5OvFF+WABT1QOoA2lZzWEtI5sfo5wbrjgGU/2sB/Mifmc
poQZ+SGkF6jBeaPKumm3XlT8p0rHEvTj4I8nLl8b/wm2t49KuLbj8WwvvKtkOvcA8GzKISwcyW8L
wRrXhUsCY0R1x+k6y5LCJoG23/FluzvwEsvazMJQ1ZI+igVzOXevCNkzc5UwmZhCy9KuMOZu2roN
k46byURCu0NonxASUMKCB2iL7GRZuaP8R9k5S3XoLwje1sm3idQAel6yHfnb0ufO2Jd9r6nRBL5C
Vm4Rq4oXj/sYVzd/fCmFybP9EH7LCgKbxF1VVcdBUmcBInMuDlRBFQc3xprCkVudQIghDJnRMHLt
cW7TQWlNKjSykVRSgTDACsi3f5n0amR4V+D44/BtXzZAx/HkrRM5CFEH5JWw7Vszpqbn+uaVOZkm
gIC2pbSTWKGkPBVWheD+t4rgzxn+fxBG/3613NKTTl2QMwQEwpg0/VQh2KbpDVudgJuCWvLIb4Hv
GFdGD4lcpyTL9zWY8ZYgv+uq75sfQsDq0wk105YQczJydZUdl/p/TjOL1+cNsXMODbydi3lFw0/3
LZjtuP6bvobAC9waQx5f5jw3MbXmN2p2rD+v6sPwVSI7WG27FMR2qBQLB/JzxtcM8Zd6MNF4mBXg
YIRqbdyXIWiqNtUtvdAaoxal332ksl2EqxNpsI5ozUlxQWr7gDuK4IjibEtKgKixs1aZzXE0fkpR
cAn19sHlYbMSsOqSYnInzeN0PT9bii0fB8hEergxEkvR4okSntHiPDWe77KuQacADkDY3DTWt65P
P1wt+tsrH8KqAYyTLSp+/3fxgMgq30R2iVYpmKdfBx0AYdpi4J1kZ+vLAC+rCF4h8N9KzfrXXxk7
eheqhhUwBedQJ4CcMP3POEdJUgrGT5VR01NORflAFaOzjjt2/saSISZyiMqYzAGvywpw02ozKZnw
eECa87Oidl3ptWSx03Mo5+/2DYANljEJSSsntfeE2p2sCffZ0KZCJqqA6XePbbKPMjPXvLIPGmp+
GgrVvMb15dWi1FRha2UotAmnNy2Q8VvVclh7eVW5K7sYmG3yOOMs0zLhDqX974CmPv5OrXg4rd13
GUIT/UJrEavH1h2S02afrlsrkjaqib7vrY0RU9VJ8Vf4VYZyCLBVEfjKwllAN8xiNpl8Kz55h4yJ
6HxagikI72pQ5R2hMH1LUvtss1b8ErsOLIJTcWckSy17KNdj7vi8zXUQbSIPAzJ5R3GFTKJZq1m/
YI95Q/KVMKnHIeiy96n493cf6i7uE0Coh890F37Yy2JA3cRNmU8Ik9qAbRPngX4U4UZE9X51Fpyg
1d2m+Kf0RkO/CSgilqTvHAjhGTEFvlFDWmTN01T1SHmuRXyD487vXCk2nd8ZAwAkO8VmdENTmxV5
6veVcQ8SVT9FjsUexI2aPA5cf0EtWyqRoPCJu+Z5uYKe3W1+YtfbPqlVxCVSpi8vxjrH/WBfauuP
T+nBPWtPRWjIUEx5QdPdHc3eubtzk2YqS+ZyWgGot5+7aG2sbGhscnuZGf6BE/q7miIvGQ8kkKT9
xqpiiiTTny6HeHKKuWV37QuepDbxtZVumfqIh450HoVj2dFTLn+3mzlv7BGXAufdvDXGO/JkRz/J
fKxEOW5+ILDjoMHKDqKa9mJxBihC+mnDCKNmj6I6rcwnAYLqd59/u8QugQqsa8wZbdN9O3VNWzji
HDYgdUfrtGedC+MxqIQx3QeE1jRkOmkZcYlYBQpjOjo2GAz6V+JVDoHa+SB1a/rElMKtzMLzdIEi
QTsVItnAabfEP36uzJbel8S04R0AAKwVMRYkN5o7u6N4Dyd0aDe0CqI/Iw4X44lRtILaeSTWM8UX
gir0g240jnvL1NDzcT3VNDGqSwghr1wvv1sx7jJqHrmICpIqj84P80VHBlMUT6bARIzUgEAq7QwR
AjxIx8+guvhOTILhjgBrV/i9qsNzEDW9kKPQG9qSl6AtLVFvsFRDYh/C0GQ=
`protect end_protected
