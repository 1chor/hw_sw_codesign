-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Y/M5oRsKwmAJpvpYxQBtXhFj4jJu5YkOw2KNnNud77BeIVJGXgdSOgXev5NFlwGm
LIbow9ofLkAbh3eCRAU8/8PaJfUAGNERiAX9/wQHAm4WNvrYcfgySaxtL32MeLsg
OXWuiQrKdo1tWuFFCMfs2fkBTZA4/6sF33QC/na45I4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 12464)

`protect DATA_BLOCK
WB7sANuUtXEvud5zKtmA5xq2PGbQLzsPgGcxxAHvbVy4/K+7aKaMzap+Bn5c21/Z
uVBvuQuE23WivUUVreyXyUTaW1QnP6r/zUQFGIxSHFsqb+W45yRkj+sGACgyAIsq
XvE/LwOcQxJolC3KGAxIYJEueK3gp/ajQTuKKB9Y/g7hKRRV2fVHvjnviBT5usjN
chMCeGhLskeo5RJ1vlIO1IFcaQ3b1elfiowzZbkrc0V2UuE/2fJtVKKYHF/8NK8G
0/ylGEBVrvm3MWr8dEoO2JFCvN+Bmv6qOvmjxUd6kla5yd7jwAVCXOgTrfuEcH2v
Iokwj3GsW2jANW2WiFIQfNSN/i3yU8ygfLFQz5XoxYoequ3W29AlmcFsiro/qPKN
GzsdpksC/9zLzHe6rhZYA8Zu2kV3yZQd55ELsKKg8lkiKaknz63T/3a+q4bwDFO2
lP0vPHVDPcm6Kqz3Ds2wPh2I3xHJ8xlLWOm89zPJMqtfhsLPUGZlxg7DUf3R7yRn
G0NPknioafwWi7l3Emhy681jRTTIgYbt0RQS3uYVpvhzGOl2+rTXxdhtuCm2zZWn
j6up8jjm43W6FFf38MqBw0klwbviNCEwlSVZBGySZHCkxQWQRrtUQLLR+wAJuhx3
M5yPepJpNh9REPx+H7ZW7+vxoetDXjbJAkHitfh4hNvjoAtNvwevzjXbc6Rq+MeS
Lu/AgHTnMdGnPHwzs/ljYsX4/GaVv85iR626VHRLYzgE7OlY8FqJHMtWpQzxbD2z
XIVr7QeMtoNNiw15RR/zkLOun8SQ5FO67Xu7KWeZ3U5Mh+SVHP/kh5p0rq2S+66p
/1P63Sv+JhcEHZ7nDNF08C5vtFhWMqlS3O+OOk5X3GBriyJfhaGTIxgYlPCALV0p
eRes0xGC3W0Q/MFJfWTbRLJ53PLdQQ9bcB8Zq/4ef//l9mb5vKDbw0SSzXndtqfv
DWtysOXzoARhonD1gs1uziSnEIMp7vDqcbnBkIUzNFrRBWnnxPw1nPwyw4fcGlcI
qS+0zyK0e19bJ5n4b0LlfAMAJK9OAS4QVRS1SNEFZDis3eFc0BfX5QAFg4giKcZ8
6qEeroisiqbxnrAG8TqcqX1DN3Fb+jF6s4P3pt6iaaNPxHrCvMUqHS17GasoeVXd
UfVjHY9BxMia5g5IqYvY+NMngcNtA0StknehL3ymCKaJDbr5mWRo7M+bYwcwqPOq
ogIjL4wkgyCQAToQpJQgFQ8BFFGYDDhAeiHwyhM+VWwHkkW0S+wnXdJ90v2R9+6h
GYwtAmmgl57Q6W9Jzj7jHPxXzmNHdvQNUyM6CE4hISZCwmoen67Gci3IxiAF2pNI
P1W741ydN/Yk/3tq4dBFM1IEMdBaQd4zRxoK0k1Zy+c8+FnKYqVB5rzJ1u0fDksK
OO3z9BzlQYtTFawcc2SenT1q4+IC2U9wEisw/2J7t6kcCxBDvybzjx5/5xB/dGzL
UzZnnhUb6GiMoCY1fflbUW4llhfrJE/sm/Qh02DmZNGed1cjcaMjPsrbHoanuKnr
y3sIhuyEbN6MhDFKcFB6rPQvW7Qq/3hNO3yVN7LEeiMzyq1ynVnoQudRt2VVK2NX
HhMoia+pfgpvWldRmU6vsDoQRh7f2cg1iUqTgrvAbORPe0OBdsCC+AwTfWjrsyXE
QwFdhSolodIomT8AenZo0NMdqSakKnLwrLPkADoIthomhLVwM+fbShPL3iROb+Cc
41cmhXNPrTyVRQbWgLKp9M786pWnK8Q1ngKDJSKiuVZ2rQqAERrk7beZGJijxczc
gXmOMisVIXRu2yR7/zJoTF6qPgQ2uUW3p5MPs0R5oJUvDR/NrCR7DyajsIYCEY/1
XTcGqnYqzFkq12KRBosPsFHhn7G29o2vYJ0WiK7we+HxNVYV79N5zUuVqtiiRH49
Rhm8TyZJJVs+fHHwyj8+1sjWmARtAiMKPcRZNTEdJGp4ezlerUSk1TuWVIHVF92B
rlDuXSzmxHPUZMzKjZzxz0gXrVSX2NlYlWVRiuNrC3ZmAxCFM8qHVaQc7P1XHwG7
19Qe9Q0AUoECvRsG7hjm+RX8yAesb4WC5yWWH+YN/FEDswx8iwyEg2v1Lc/DpaNX
n0IPaqB8R+LAq+Agq27fOQ4ajnNXLoyKnNeskcU/hDBQybCD2vkTNQTbqJbcMDiv
nxifJtVBZRukS9/mdld0K4UOzIscwXTxDHYQP6GRMPqNXDLHkmmmjErj49CT+98R
PTsYKFe5pg3/AFfoLX82bmOLdNJXs3ZSOBC9hxOOE5o/mtsJCX/I0vX4Y+e2icT6
eHmjdDxoA3tbUcrDJodX+aceARrqp0hzeqHHo9LxoJT8c+Pokr9lq5kHv7MGIZjB
cA7+lg7k05/Ock8AUJK6e8+Ssa5NrarvuGQIE3JY15yvM4DugAfCDbhxgO+4UAWJ
hHMEDR66YCiococ/drwhM6c/+q8e9AMiWFJqDZzRUMupiXoOfThrrwBmSdfK64yA
RihGwQdY+vAV5LtBNMSARIWo1TjskA8PctI0gNIYxcwGXSJzc0stYwRvKgzNZZh/
+XrkdqSoMWRKlYUkR0J8qYO5XeV9z1qZ+QSaLBs34p7wzcxEcMcis0miaH0J5NWs
2jb/+/1r7sy9R8fxCPoT3Ld+Vh/Lk6R4hzSLk9LrStxXB9+Lwofz98omV446IXSP
FkYwqJmCpUa9FAseAhHTgyWcTrVZpVvKO80QdC4nnoLjo/blWCk0gzT1x3j+JJQk
+yYv02DEgkJk52S5VtEt3PnBSNA346wcdsOs/mb5W/SZWE1KfEQ+kUwcMW2oJ0Rl
1A9sn3FZaeibuJl+Asg/HK9P1ShSkYeKikN1YwN3TIKrjC4yUedVAUUHCwer5nCz
QVldeDJabrg6FKHPepxIlRGu5GeBdjgnCuitvtBGDe2nDWvsziTih4cQOiPE84IK
lGhrVPZr3ygPsnW5sTRbcRolI89p3sdOgpbtrxP3c90fxemk1CrcM025YZTa5Bc8
uOMoB+Hd6p8YMDOqMEDu2b+oUt3BvlX5KWC5wvQ+W32Jc7vRlUhEbhb1HFskUMi8
cTW1ijlpz7Vvawfmqs4OH/62YgTY3ilAi3CJR++iqE0YTpoLofQePy067+0u2n2F
R3v57llxZMGu4QDs6kRjGOvDm6+tV9t4eEcOpfqNg/QLUIlkZHWQtWN/0+CtUUMc
IGz3E4iEaqUQ6Q7jor2lyQpmO5zoFHKhQDePHHpFm3n451mx3nmOoGQoE5kjV1x1
cuW4cOAd7eTGuCKrCJUjUaNXrCvDZGA9bE8WO5+vBqjRkKaSyu/7Trb4enZBeufT
oLX22/vtrvjPzWQNZBl46O3PJHcuimXxyeAVFltCnsAKsGxr7veORNoFXkp7/kNd
wsfsbp8igsWr1HZvQ1K3MTXljv5NoTGMYqrm8M2q33POZlOlZh01qf8b17IKg7sH
+nkHotcE54RnJY1KruDUSjFHCjouSxz6OGmi+aXfiKJ3f1NN2qGcxOQSlVjgyPBs
DqNQ+rSyOzyrfbcryVrCpjoW0qayJr4HJLFUcSVXcPyIZjO8ZR87YI/Z4mQFIwv0
RYLO7+N9nXNILsrK8YCnR2hI4UTNfqiI77hpuXMeOKe3orSHdNmcEFKdJBqpxtmT
zXbFVFWb1tyL5Ly3A3FRF4DSdJqomowh6cbv+Nwzvcp/b/aB32vhrm5FRoGajY4L
gXeBZdqrHci1JDcmQRifuOZ5RTd3GnQgccCnjRAnTLGx3pEuki05rtrtLO5OJOwr
y+X8XfQ7bJmmr13fgiYdY1iNHj7pVGziHirl2Lvfqsi3yIPh8C9YPr20bXwXZ8RR
PKHJz4wJVPpXIhETv6qLmvYwdtTAlVYM1PIlMRN8Qxa9G2hDpZHiP6WdxXomaEDJ
L8MFtXmeruqAzexwa0Hi/xIQvHpgYmfuxYFVXNltyRUutbkqcGGLIYXfYMgJz2r3
aWozZSnSUXObrS6OdSAvSe21oUL5ySE7ULnXBpuot7FAJy2hlCo0mjptrCcKBPsl
ZF9PJja+uj+nyfjeIYst7aRsDJX78yLkEEqvJ2BXvyvmaeU/U5Ltbst8iX6ptr0j
uM2WuGcPnGQDNRmlv8FaGBwf6onsmmJd5EWgYFqE+h2SjsfzVV4OPyAiAKLOMrbX
rlfdVvpRT9ESP16CHPNlEsyqnCyMTzvH/8159KNWwLe3Xbz9aiXenOWqBpNUOUd3
861nf4FTq3eMRGoZrO+OzmF//WMLseFNAHm1tQPWoqrFsLYCZX484SKHFs0H+47j
p7Htve6XjAMfI96PkYFIA9l4Xz8LeGNxxAH39WA5z4ZIrrAh5kW7bV/VDtfJsv/l
9mIGa5vK3kkDBGzzMcoimkpAGZsnNDsIc8ro1XA+gVxsPZ2qsuNmI1YAMPaM/MjR
hgwE146r+L3gvrBSOF1WvNzeFdpZbkl2KVMsA7LgQEwquOv+KgCSxdxgZ75Qx2C1
imXcQahouwLcgzZSURDUIBv7c6kUttiUnmlxHBSUKydrN3HcjX9LtyWthqXaxqc1
wh0aK+DFRJOv8W53TAGDvkJSqekOy1rO3/hp3bDy2K3YFkgaWMQ1K2pYhFD8EIFJ
FLLeSb6pGL+88gOn9hEVmb09xS3Vuepy2xplScMWYJEZofYNpAfUrRzhCObxJQ0b
6GBbQem6/ech6Pio4YPRi7Fvi+/zsvkBqWmwSRGiZvmiIzZFVlnpXqCWTsQxHVHx
8aHlCMJFEelMTgtRohgXKBakdtMVhvSZ012xqKqOd6DsUfKqCdePgn+zfTSEzjck
Zt0s4fh4EJWn8Lp77S8UudabR06gObtRH749QCBQd5S+2uzvX1Ham4AqohjhhgVs
bX4ZsbbMOvutg5lO7LQmack0tco/LtWkmo4RYkWiMGDkinPCz2zJo8qIJj/UWM/b
+YiQJX2KPsMkVg7dQkJiHGhIjIr9j2218mUxKH67NT59IxVd+gJLU3Uuhqhzep+Q
m8sDFJKDCxfdwVbTdS7d9ViynNW83dcPZkYy+kRm2swB90McjAzJmviaudG0R9rV
FB8cPOcSpv/OVQWM16L0RAel/dK4ZXAOn8l1kJxWlT/BTW0J7OS7ytHhbFesZinK
reOR5DlYuzTN4EhepdVUWVyxB/Jwb/3YJenV2myRUNMgwEZWwsgLDhXqhm9BERdk
kudjGr81OV8xioZUnQ1dyuGDXMm6qcUlYTVOKp6Dtx/A+i2Ka9YyNg+Qc3I71YUt
BOtBbTt0X5+W3V1XaPvj9QekUJ+Yatg5C9uv5i0XTd30paxIjyVctFEJ0rwaQSTM
0coiCuabfg886YdRyB/N75IzTKkjAk2HHdTV/6UD5qwK/LSKnphonRNsiAEADfHS
5T3pagJ6XYkCjMO/dsoymL/ZfYI2aC5cvmPezXy95oCOrGVYYSvRHCBw9xqCD+DH
jLTccyW9OKHgAyRFWsRl7WWAlmF0eNa2XZiz4NXM/ARgDSGU5k85/Qk0dmMatt/h
SdnJ5al/pOPkcumqRsd5yJ/AdKKFlzfelPQaYN1yr5BZQ639zEN2lWTUlHN09ohm
94oEQFgTsRG5SKiQyr4T89eo9fosB/lzKvT9akHXO53sAdh5YM6TqKlVCETw4J5c
NnzzvKS2EcQI8+wT/qI/hTdNkiskK69fqTd+xFGEP2Ml/qe07TO30VgcNlBv6KAd
gE1F9YeN5d5MKmnfvh1ri6k5GB9pfP2FtmHc8kCj1iP4EudlApqMTAnamr6g4SF7
0W7nQbPaf0Tcme6cD0hTAH5u/o09vcEmvOZqRIrfuApIqZkWG+4WHYVK7BMLKrpV
34XRaMQ3xPyM/Hjxc6EeRe6OmDztp1cHbr1C5giz7RvZ/yaqiZPEichbtNI0xUFM
JZ+VvBez/vTDTZ1o6JUGdVfGY3OSo5SupaPezeEpTbdF1v+FELlT5B+2TCiODoda
rjnPU6cWskLj7OTmnFUR+aZ9T/QvMk3Ex0nnUbG2CVDy6CNduyScLKriad0x2xSI
tL1A1PPQMLP7B9l3E0b+sHiZZEKXzDPuIZfAlmyF+kp8jULU/mhv0JqYbJvbF1/z
oA+j4jsq2c8QZwUsjfMh5yEF8mJjMbxJnX1Fr4m0tX7zG2FbaCRX3qmhViKDJ909
2yqqeQHtMcrgqhlbanbt0WY9xTkJKmLws/LOwTmEHg4vfADBoxY8O2H4XQdgvZB9
gGrswuHQP4tOM++VzRFkt0hRDPyOwiTSqA2E/wnkb1TBZALC8uKe1Jhnfz2Jgsg0
kOj0smY4sg+QQ3Nc343+ZS5wJyBZdmrL0EdgLWmAIUzvAWSEVjtikRwsrTLU1G4J
BK0q8XR3l+zhTE5akJORn/xBByVlQwqDT2OHDFPKNuyJKan+QM1R8sN6BE6pnZOA
lHRNnMb7ZreVp7NgRzMj0P0yi+t/oyAfrrkkfhjqhj4JGJnFwPiOJ3ftAtXhwe2Y
wF6lybtZ1xriMREBd9GzWSKMlyJzn6NcPIU/nbo+URHdupjkaTJbCJ+FKkbVfylD
381WJM90qFlP1/CSE9I+HkqdTxFJ3BA762JnxYq0EZra29sU1rxXMutMLxsIXb4P
JoAsCS03YX+KQnalzq0MAAUy2pVFAu1u6nlFCv0+NzUtQovrQlUwMIu1MFaC4AtA
kx3SOfZGaDdfclSoTD2XJKAOCo6q2FNsg+pLgszGXJXIARk4DTi9Lftg4PtpDYD3
/7P/jCzene44NPQ6IK6oxRJRrdYUeLtxB3xxDApk8zrZK50vedptLlioT12pHLxF
tlLHAWtRk56zFy+W9AYcSjQdHJFvoEhHLWxCk9lnQMqfooFpOQF2NAnvnTeyek7+
nq7Zr1WzcC5neuDU9/4dwiU+BL048RcHbE6lmTMhDiE1JH/JP+GHpzjp9laz9wl0
v9diRQezgv49GP1nfCHW5Emorcii67xIe7tvIzNTWG59itKoqRODFUGj9GIuuIPL
jo4Zxyju19Nh433aIGaPiwkBVu1uIkSX/4zfigyUoTsDGzs9qA4HKBfH38PTOika
xVDqsxtNACl1FSpkqZmlIuE6de8V6XY8bKtdiwD/wDd7DAdFCEO0NKEnCGCVSKLP
DJz4E1hjDZtwwEARPgAjh+MbwifH1TghggEGjt6ueovnhvHMyNbUtbfko2h8Yak0
nen+krdOg7fFiT6neMazTCruHGrSQ4wwh/tBcQyW5jrjpVoP9VTik7oPq2GZ847n
tKrXfgYxhZ7JVhNercE9pjdTxsf8D+pEi96WfKMsoKbAyRh6zDlavwDpccT8w2iG
LI/sgo72967E2Frd5g7iZMsyODMRJjZ6XrBRaT+7TLdmLj6ZBBKhlZF/CDs4cZcl
IS6/by7x9bmPsh8hpGphCC3cZJlfSwWzafzRtWyzIzH1qcB4wKWtAu40AGMKY8LJ
KVfXVRdEGqO4u3d4bolWkaut0J6f8ev9Jj8NJL7YS+0WThwtjeX+oQEUny/ubIJu
P9juKWwrQDDG/6oCQDQcbc8R4SP8ERU2Fs+d6Cx0PjFNGd5SasZIVHeF0f46wpKq
Qu5oe8hqaiMnPa+CKrx6VwBnwQxQXVEredPfy/PoeoDcu2nUahCgu1zBxSXBZgaj
riiAQ/ENJ1ikBM+Ie4FYY+lAuKMiMkmSrEfxo2Lb7YFlijOphslfbt5QvbN2aoz/
PjtzHepnr/bXPlbxeSNeHh/4lNVtQAcu7OM+tXhvwsQdbe2D8JDYOh5a5A/yrxJa
ijNfvJ7lbIx45pnZZSlkxrsRr8KiUuGabSUGh1ng/ggUcQZ05w7fPCTwJa2S5oIM
AigLAf0FtoNiDAKT8GjuwrqjW0Ja7A7TieU599urvkvQF8F+Y1l9/BLyTEDpBtVu
7SV5cz/foDcMPjfXOySZon7zkv0qlwiabcq9q4Ea8QHlFOrPE6D23vbmDBsQ653b
o7GBfH8Y3Rin/HjAiab+CypFcY5skXT4fxpsieNBaBrlVdIvD2xcz3pikUcsyBDN
GVVnj/09OOMo4t2VpLalRmynn8YmQHt3ZY07LVsmu+owZQDfbmykqAmKALq4u8C0
JXlkmGsiOgQiZreEU749Wi/wHpYgW17m+wE0eQ8rFznTSObxXKWbQ5qoDqMcsOVk
imFKr+/h49R5uEzsRQum7e42YYK3aHfxuelACzE80Ds4ym0+hYKmnFjMTAbEqs8u
rL1lqkgKn4Q4v4ZnQ4lJsvX8E6QpzrYLiKP4tlUevyuGn/4nzuwvYAEUguzkwWBV
TaxHrAn9HfkCB5vnPXs2iA10r5f3of3vbq6s6o6YV5wFRODR5GPYXecqfEoKUiBA
o3hABWjdm5fvrpYjG1WAwU9/kVZosIAulTpnz28QSTclwAl8lQ2dzl6SxCnxM5yA
g6Tdg2n4Jm/4YpkmFFlVd1IAsjQ5Mg5lb4JEaCGvpyU98f1vbIu8rSozbQ5GRoYn
rpk0GS4KEiOCxtU+U0tMo1XH/ygauB+vaG8D/4A3lxq2o+JKf4Bm/wI/PNU7YqsC
r031ZAhU/L9/zc8P8j10GW5ggMf36Pj+YdiQlict2QGea5s+jO3JzsFe2yqwCUWQ
xCQgFZWLTt4M/URX5prwJQU703By4whahjkr8dQ1hYxuCwAmpYXS9/ZXKDEyMiPv
UyOPYsVKJMlMqBxk7yBHVsyt/5m+cxWnA2+VQ7gXh3SwMEZbkOubec9dd2Xlu1RL
4hMQbxTauFeXUZCq/4mFA2817HQfPia2roffwL/+xDlyQtQEbiK3d/ckvtFiaPXK
1ElcUGAZuNv+J6kP1JUw6OVVni8tW+nn2XKuqdAuDCHp26UVxqRMgmu/60R0FBJb
H9s1ntjyusOCux/nueBBD/BCj9trLYTIJEEMFqxRRSQIfVxUtmN4skTuWL/R+vMl
Dq2ev7/sUQJwNgxF+IfymfsV0U3J52xQDkjaeomlVj6Luf7HF3C9VN0+rmOHaB15
lcbG/1Sd0vpBJMiHsESKjQ+LHGoAq/HxRpQwvNfAlxeZ6lwgJZAFr2dvH/Q/JjlX
465xiZvX/C2jOTWeqSorXUAALaV8tQjVf+6IA3dUY/Nxq0v5UTeDyg6pqqDgcxgd
aISIb4lUqzGL4mSX8W9hvgfdp82RBfTEwiR+O5YSfio3+ViSSB0LRQKcTMwwzFUa
XoNNjYdvKk3J3sW0bJknaBFHx7+X6DX9hqmLc3z0+yzTW4tSgaxhSfG9sl4X5nX0
QBkY5T+RKXCAec8bnJKff7kvEOmEMrc16U+BQkPFNDdcUwWuuSLJwoitro2FNt/7
8mF0Iw2IDQ66byp63JmVPpGBqjigyilzFa1H0d0YGUrpiam/mLG4Yoe3gwy0XPBS
sS3i3Ll2j+C6kpun4qPbGxhqnNvNDA812XoLTBXwkBTgNcVdmGCdkNN37WV9Ojeg
tA7ha7p2PCGvWlvC1o1HVMR/WinmBEc+UOZie8cZZczXSrbfJglMR7JRIaLbwFkF
FOjsNRubmvhVRLr62e7rprcBpBniwL1k4IPazAVlci8XpRI/PlsH18mdQAsD7kqT
92JiUWM8e3NYvbMNGxssfrWVF+nL4Z7qAq3xWTuw29YXEL9gnvJh9rh/hdCEXqmg
5FvZhSyC4tbE74Ml6HWTDTJaKP4CA+XX1oCx1qcfBThvLopQjFfDrG8q7RfhrrgW
XKkEVJU1D2DxH2J0lEvxAoOTW5UvaNIeVcgCqbyJlPQPHATGscgyg3USla/txKTL
YCM10IfuSOjB4v43L3w5N+H+ciRvi5CHILtMA08xV5Uwnt9zUcvOVtG64X4iVdAc
dm/ffDHfevQmauxrRol6kQVlZdAckRFemXD2Ib/SorTsntNByorRs4E+z6Am8Hnp
7UFIfZi6hbbCARtvlePr63uOufl9IwW5nwVnL6viwZxc3aNO7diU2zeQViNlF5Bv
iKN5lVsYpIr35hJnXhjv5r2nR+VtG30+aQkbEJCGgxSRKI3/i8TbOfu+1lmlBrAB
J+fWN3ydY49q64rIt6SZNjhzo8ZrEjJsJS8FD7gpsV8d1RPR9hEh3m9zP0+I/Vct
bc6A0xdBK7a+5kTNlzThYuQCAVMaMSL7anFsdD2S7g+Je+dhOJSnBKHiPo7R3sLi
xompLHwl6vJg4OJD0P8znLccso4pBG8v3CXfSKgk6jFdxz61ihHnQzP3MHsTuMsH
GhrNmpMtVdRpsLuhjg4Ji+0CYNnSH3vQsTw+Gy3C+klOt/MpCH6DWDpVNnpv2OtF
hS+cAKJbQXxFY4zI+0AOBFUx/NHcn3IefXBxK7zdVMlFDVACtM6BI3tCE42jUqdM
C9X1oQXyHRvG1DBv6PrE5bJJ7ZVDiUk2WtUBMlMpMEC+psV5LAs7kgq7YDyXMQ8X
fLVSXyAxbsAV6Z4XuToFTrdwZKZpagIbbVT5a/B+Y0d5GJqJCTBOXUVKrjS91G4Y
j1507/09pXtzNgRi0PnwXhBVgNDoQBpknEj07icFysUN3YQmYHiRdBNwCG4lDbme
a1yfhyzQnmFCkLQCjOljOJULbGGkfaXIJv9OHny75Wf5HPfrriBHoKPDQNKrE/fU
C/fV8C8A1s1zIWJH1CWcFfmL0kBXGuSJOid5vdMB0LNEV9fa0kLvJ2++w2hcnXmi
3KAhyo2lJPPWG6CnvbCnW/i3iI50h3N54aDFtdvNL3PrL5iJSczKjIL6dZkHTy0s
vm+AazyDPk9whHo7JV8Jer7Yuqy77JFyShupXJtFPaGFwDCJ0K24t5O6SiN8hx9d
l+Z3Idb3pbtIdOEKXDVem9YlLZ2k3A2C9e8ESA3v1qOYl8PEB7qiFfDMS3Ocn+Fr
EyeU6+868+iPRZEEcMsh/eZ+GNZRG/zaPnt8PqTqlehtxKzOJ6Qb9tvtXHAkd+UN
G0eOi4seldfZRXOslUvz+x8X6D3wziGdg/hd/hew3iQ2awfaMkAO1eHfZYM1NQjc
INGkkXPX3qtpFMIIaA7mVQHfPpZ/Gqy08LbUNcuVnrGqXbamLQO9jkU+oLhOSR7Z
YbF3ZALjrw5rokcZTvXEbD5Od041T1/vh1f7HpJS+UWZVNEntoCm5+raFGSQXRAQ
QDQNPpTuSKLy8Zp77NagO3pLfF+auHuLsOO3Fsmq7vM6Ts46dyeyZs0MRN4MWlme
RI6hfKTLTqzv1c6DDnaurSelVifKtkUxXrKCID7pbBn+TvmkbUFcpDoNK23sMMPA
Kr3uf1Vr2uT4iPq37HzwtZYqkgJEmEoewQ72bF7y8vropARXiNURViHt/zN7DLfn
jTMsbn3yYsTEMvj+tXaPXK1P3QWr2deBJsdrDBqoTaTUutzBg9RlAQGpT47/yvry
bZnv3BJgtneV7iyw2cXrO7Qcojc+ZUXgCiADQqKG/BkroZuT1po4UZgW+Y0YEoIu
W2WTyQMmrM1AjKLj8OiWT3OLzp/f1bvZUBrAkrbllmh9o0L+SFrRBaO5Efd51DaN
wiBEuU9zt3MumR08uFMaa9OQzdgkhqXx6B+6hVCcCJstDF0TmJz7qed06t24UHqU
FlOpNoRdSxFIk3b6oyWeSnvJjukA3h9zh0BfutAOHu+CbB528VAK8HjbUGLnVXdc
d5DugQjeHgVwDu798q3BVwXYccEeF2gmJQYxhXwt4zcTWebbIScnIhTwIRPvw5gs
LWiMNQNLqYdtbyYoxHaAJMERjuNA5otqU3ErFKMfIWA6ksAnCSGealfXZ+/VOszE
CF1PXyhP1A1QKEifRY2YehQOTkWedoTfSfLp1FMTlYilgBVxHUJ6o3g8+R6jwAd6
relY9rmdFk16tfXUcEAh656BkTmGhPJSwHh8EKLE3n7az38ihUZWGDgSqxlnpUZy
UJTM61zknwNWdElC1yZ4M74l6+wxDe+aOLzM3Azh4L5l8MPEtIoaKLc8xGlFu0aK
hdzCmyEqbT2mKP9SY9m5gQhTLSABrGs2CXy1JSBNBc1zo8RkM/wGQbB3XfyzuueU
SJAFX4K1cs7dtFRXmDDHs4JrQ8t2ReRYRwfUsqs2+U5gHWEAFK3uiZ9ckOB0jERd
Ae5io3IBXU99stBIDfMH7e+ffxQWYAbPoclloDrhFb9vKL2KLz1Imj4PGMY7OUqd
AEAv36PwGh0wJNYYEeDUg0g3h1uJR4XRAA6JnyFocE7PjyQlJo6tYXQ5cQ4Z10oC
niNMmTK/PzqZuz8fpFMGz6mVkztaLuS3+nvtaOMuiqQHqqsNSZX8NXQlFdA9sg4m
UtmFubbcmZDs2GktNA6vxMcAKQ8xnMLapWAgHRXyOxr0Z+U0UiXXMDQfkF+Oe0kq
MA94Zk8Sv5AmFm2pOx1t0JacuIr573uOBz3TLvIG3A5by+tNinEZf8LrEdAISDEf
ZojWCZKVnByxxNQVPYZE9MFi+Ub1JS47pmi0FgVjJrdWiot7rCEr9GMaFONWtCMu
7TkqKCb5XBSFeh4CAGBpTup37mw80kk7/6hb8Fc2mU09BZrLV96l+AlsaMVeUfRr
/wK/1IQRKb7cP9dSrunjXUDkpno8NbxVb/gGFZJFLbOzL1za0aAKHYw/07Q0zuAw
RBKW0zBHk3OZK9vwAeymXZpbzIz17JowqAfl3HGMDHR7R95PEUz7FzsCZuu0fIGZ
gLK6D08yyBtignHY0DEO8eBloRDAztMyBAJpEfmiFv+RqDYOl9W8k83ajYVPw2T9
/95YjfkjrRnsjFj49T4qypXFifVDYMNC5RMJjwA7JKTWagQvVQfvjmOiqZ6ypEWk
HGgvCcLzcyDVkdxRWW+ikYINRP11VKouTTDGdUyWKPjR7uuap1wPSOI1jtO2cpmV
TePeufp96UB6FdGZoOnr/Jxa0MJfrMF5Tb8KKWUb069dN+56id+vEPIXxEAHKuHQ
NfiBS+tbgAjDayDPYA4+sbn0N6QsQCT+HRzJIA+6pKm4OgBGzC1XUCyxeppx0bIu
imF+sq44QfuWRkmiWaPJzxRoVjOsTN0OU6vSbbZPKRqRDQdEc7P8bbU9u4CH4MpF
F5VqfkeXVurr62C41d7oHqwmFil3tab/PxuJAR1yDzBNvY6kMLs1jhzJtZcTWF29
LbAMhSH/9uWQEpKGnbh5wZ90kuRw/1w8hEwOMlaA/V7vqqF+jdoMrC2pc9NNr9nd
GNKOsIHMZqp2bhnXlLVW0GNKKOuZRXE5g3aiO4xVrIgpbfV4yoz4+dVwZGIluY1I
MV5OpvKpASMGLT0y4EO/wOECDtA5SD4kKMEyFOFQ7l+6fcxiOSa/peQ0nyKktUNV
Nq2BKijREmIwRYFjXex0W/zgLC5l2AyGkTPKWp3mpPzb25M1H2g2IEPl2+r1YyHh
nLPy2dsR5mYvexCScLF8Mexz6L0uopV7AcfXjHIsV0bbVnRBTrVHP7m0aMC9NaJa
Y6cEIT2Huyr6sgJylZXIC/qjIHegjgAf00uPGSwBnPeEfZfxjQjYDxdEOrlPDUV+
u4kpvEdDwn2wP979cgZ3O88QbzYueOqEEDt3xFFY7x2SuG6hGXy77uR6liZnK/uD
Zf820cWCVbH39VY6GBTtezlbeVcIl6wU1OgcJFDfr8fXAPDrzoEYz9MEmv1EcTcq
J0xZnNK4pDa9dB7qgCfT0lxOPf8YYOMiTKhOvNSCSfpy/VD0aSvsYA3q0I11rluj
eEkbG4tENgGC4uMONnyaT3LXUFGwoYaWqXWS61FY8uuUBrpg5zslPgi6C5UCsSZR
Xc7+Nsd88C5j/DorsJzKnd1DM+Rck564uc9k1K+HN9iOB1ZIBPDWxtNIjIwE6Qnd
NhX55Jjax+0E1SYHFm/rSLKC3KTbzbLqJMtjzOAspAYcQfoc177Vut4M67ak3vN0
5qv4FH0pIX+OTgZGpKzmZtwm+VA3dIp9kV4Zk4bcHiej+vuLZNP26N3/653wQ1Jj
J6JLS3cN99jIHChslLAfxcnyVvcgTGHSmO5NRu922MTLD+XajOxgyL9cgDnNTFVf
qXYsZK7WusJ7QCKNcQbifwA/1v8khiQXbL5hjgXZMUGEP/VWpvs/TtuVE9jX63fo
RNMH6PV9NAKdCQk8abinD5MIejtXNDtK35Ti24G/spe1Q+eaMrAERVccdVJzPrk5
DPed4nM4kZiwe1DPrfU6tx0iXIGuLDWbCnbFC059U4gYI/BZcXNt4MdD+iyb+rD7
AstsTM8A2ojbq38dTVU+Qz3tOWv05OUCL/K25f1VqRJP12o+Ok2MkhM1FKTXLGso
GN5qTD6IdVW2AiWLfzhh/Ujs9fyuuUjstiM3+9Aa4YRVYHdHLPHccCYkbdouIDj0
P8Q2RopUIAIx+TG3Sov5lqZC3F+lvOrNKkibtiYj33fOW7kyHPQJb0k87q3z4XcT
GmWs/bdSkzTJEiKRixcuduJPZWvT2ne3ZYM1+XiG1K+BGmpiG+Zf5ttF0+aphl1C
LG3PAs1I4GnD/UrepTALlqDnCi1UThGtUcSjL9mM8PZg8kw+wKO8xYjpdOl0qpW7
B8WmHyRF1CDw5KGKZPPt/csihQvSgNzNF1SWIHkls9VBS9NDg18NyCXn0WS8FAz5
i6HdAgsKMzNkQMu5iM8OYCSbS1su23SNKn26M1mkGRxDte4RwSEs5vres8lbRKTl
/1Z/81Y/xnJ4CIJR00agFTNnSdY8Wup74kxUJrKlnqaN3NPla5kvpLim3bdBXeZZ
0SzGt+mN6Zi2b4qKGlNtz6PT7W5odhEB6EOR+Z4BViXjTus2F04GQrH6+mEujPvF
PBJh8fk/4jnH6mUf+EqEOrR4yEPfaeXRXU7oMPS2OnH8+uX4j+Dq8TDKtTUgX5+W
Yc1eR4xQ8/jOl+vMb234VUQJ0Ugw3eqA5V3OeO3u6IZDg8SMwDFdR/EjsxYbsBkl
ojoHsaDVfAw702kU9EsE11BDguX2rPiF6xBButbXWkdLxQ+fQ+woCyx5nnHWc9a3
WabsDqLUVWTiE+pdXstkusQ//kO6L1pyiWfbXpF/v+6R0EjQYVPASqkqPfSrqYRP
q1efkMpNNgjp741oncY3IvXO+PMULoPz28roEt/tEjV72R8GAdOtt6b4hoyWhEAo
MF7iA1pkYIr5N9IBuiHch3xmplI9kEu68EINOH4w9qT52VWnHp40aiy/CSCh0TCM
4n+XAf0BakdkCK4X5RRSxBuyl7YLWqc6avu2t4Bhr236E4QEL9IiqpKRjmcF7lN2
bWLG/v0pbzOzpvo2ZVRMVIDO1w/9UHOm30Yp2YPJWDrZcHa0VM/NALkQXTg4LLgJ
3uVhNyWxtXDrQp5+BEi3++Rqhov0tve49XFwodBw8d5rW0LvrnxUrdcyCwCoPhP8
vuCcXJ69QNkp8a4jB5ltE+sGGWVxgsPQ9KoTlmnZDa1o1UzOM0OO1YqFchW0xgGJ
xopTGsew75by8h24OTleN3vSXPnwD8DhJ+dsOB0hHjZYK9cebjVUY74iqUCHFEy+
IwP1axtLfG4lV6ijJggXguCtbV8mFFqDo6/eWaI9tgfdrlYLm41Z5fmEx5ajlQwQ
vEGGzsKajydyPDZHdamvml5DpuM+862iagwdr7/kAGo/fh5Ao6R3X6y+yUQJq4hY
xyU2cjw5mZoGHo2esX/ioF7LLStiIpnE8Kp3fZtssXLQwQbfYTpk6TAXjPSDEcva
KotWngy/Z403LKwvwN6eXktaQzEJHsi+8dtuAiFr01KzWzvXpUaNvzBcTlq+fQ3R
EmXgQ9ei7UwieLeWs6oL3F5TdCE2FazjZnUk4rc2hLj3KOJ7+9iiMTwzmPZBYj5E
7r8EXUAKRp6GEpM0o03efwDCVL9yunhQg5OsMMUBmnI8ikz7mQsDvcNInk5QGKJT
/Gu0EFCODqGE4tBqo3yEv38HA743cA969PoPkRthHJkg60l0OU7ImdM/XBIZGNkv
7WqWRAQQ/D/G4ILWIEZZJuZRR2x3iB4rueMVs0qeW8lEK63oHJwvnNQn7k8WCuWF
y9Z8goX/olGlGak/S+MNPNJS/5viUVGi2Y7hEdxRJWKwhvqc9djfF5xYorI1ZiNR
WxCySH5kZp9i5VdvAAkwuKKEUdfKSIcqUIv890JZU20OdKsri8J1zWssyzQ2x4+P
p6SdeK76YzEMiY6fw1ZBUdm2/o5ZfR1h2qCP9QTkoAHd2nRtqtM0oiIDRUGVU3q8
sSRr8nwgvRsRVB2lJ+BaCHc5+wZ6Wcs/Afg2cvNDZZOJFtw4a9ePLOxMKmN1pdDp
zBPbQH0k6aVmC52CLWexHexUuw/WeDWxDP+LH4MVQMzbl7w1ljx0tNE5iL2PD7kx
j3V7n5GxIeHaTHwPKKRMAg2tX9FuYWfO/rZIQQ4gxys2NFoVdTH7OP9/z+6g3Ja3
L9ILnbMQ8MccHgOhPg0/yExnhQ7ArEJFAWjybk1G/vj8iykKHAo3kcOiplrn4sqh
90Vauhi3Z94RgYnlc3NDHt3IUDVXy4nBSxdW8jchmPbsN1BL2yAUzd1ILxw3ceOG
3SGNkWeXZ0QnJT3iuTlhhZgCoBXHN6HsftnN9jaasHBQ22i1FR8chjyRHdug88gG
IGNX5/wUhb7+KDWRLc77SuKPjXMpH+GgQNahOzRFcQ5TRXaFtyy+nvnZwavixgI7
NyDzv5ROOOjkgihsbkGbQdPLc3jw52DleweV2Zv/OdS6rjcYgPEftJ4PekrrQDpd
c0oxKN/zFCX14WAKaOdgjQ==
`protect END_PROTECTED