-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
mLnXsP+D+oVRyZrMEGrLV44afmLBbvRzYgoj4pWI5B5B4sLEQ59Tst7gyS3DG8Q6
ZVnknQgJ4Pcfb66RI7r8DYQZp2k14ViH+o4mx40Nkp5lwr6XCZtNEdVCNfWKJPHj
W7l9xhEybIvFvoS5jhjRjeYZXxP3BqMy6URUyRWbqbo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6427)

`protect DATA_BLOCK
8y2NTXJBMYou5J+VL2j96jGwL+QO2NzxuJXaIw6irTgEi1ac+qDwgxOpchDZV3V0
eLWMDJcz2PquuE8IvXhiuWUdUiajcMjnnSkR7beoQR7EB0RppHaoEZGjShmVfZbK
qECUy78VqR58R6G8mYNctOxmohXm66IeCNtCl9yhXzOi/CAeZIvhjK8eMKn4e2tF
Dr1+408qAiOIi0ZasT5en9zLmzz5NWaHT0DzSYdXO43q0TqA8FdjvYcV892p5/Qo
YlsT5HFNEpTBLuWDFinKWcu/G0K/d/H2Qe3MOxs1MJg+VrWik63D2R4lFeDEwxEN
c5wdGW8NLzU8yTyVodW3ESfe/WcniPMwJ72G4ufZyCe7Rj+iuozYKnvRkr0hRAgJ
f8P+swlBv6g2CPzp1KgFblm4PU9CPyNOzr0XrTZ6lmRH+Ni2/8OrNKLLT4oqPJTM
3B4epXSo33Hx7rW98ARzDn7I9NaVr4nzZY4ujWhoqUv1bCeZuM+7/QtXdmBBeRZh
XJIFxxsQRwheiBFE691PJp8PSdGTOgi/xCUmyXeai2U03SLExfv8V5RDGWaelnmO
32YM3gAKHo22oSC9K0UM+Wc6AxYfYwbldokq2PQl1rLj/9cJnnRKJexOeREt799d
EaIbpgXJsSZMh1HOaoaNQ2EqNyWRIs8DAyLePlVaDoESN5V43hbHZR4b2hnGgWFp
sZoxjQOyv6/AQrYgx6DT8UStKfFnrjw+JAcazgvUPiX133q8X5aJQcrdi3OwllEw
2yTy6nJIQq2+yiJT6JmsdoRgzHrayYUnYTVm5IJICAk929F15CRcLEeGDP0yWTZd
+peO9jqFvGHYQmChyWmaILcj74VxN64Phuw4iiPXEi4OnVApfP7IMJXK6EMjqNkS
Ydk4MaPoLTFK4EyKgm8p7AEgWIo1o98quZxdINIHQHrZzZW5p61/tGdv2IaPZ0PA
iB/axQWSewrTjq/WZoM6uTXjkcjOS7HO3syF6BTw9e3A75h9n5ny1/IE1wGZ7SMy
GTUM9v15TqQE7e0TV8BeTnm8DpLp6Q3svsnBOzGkNRy0ubWzNZzknnVRJyKdkz6H
7V77wI6RC6D2l+t10l0UVv7xI6sesazLqEeQqLvuJ9cxBFktZgm0DtaX0EYyhBd2
63vQGu0grQVPSqarxVhFPaplUG/mTk4u1GEqyhjpEInaq73lBhuq+eHPkSSXc6pX
0YuwGsJZW9nzgsTApvlEY3dlZ3FMRd5lrqgw+67fsAaRRhfabHWRuJsdaylxNKjp
IUgq5MzVyHZbXJUDWHvG39+irUs2/oUHP4MdznG5e6xMrx9mdcoysdkprYs6lM3i
uJdN0hxhG/mlpgTvgBUNKlciMKW1Qp6gfIW5rjx3CqNVEl2aOrRFc+um8jvx1g8x
ieQ9mWf9Z9b1BPqCOdIwGLfAbDhhrRPnAQmxyI80AwwNu+AzJ1TvHMvf9/likOov
hHZYG+s1wAv4gySWecb0aVPXicGPl0fnJ41gImRo2v5zI7GoSlxyAMNIqsSsK+CU
mf/ScAsKPoweDTMtkM5PHYTk0CI0S4YEmT/ixsJzR4tBuvEPdnkliWDRqffsY1We
PSUhXaNxDqaBo5R9oRZNfUn6zXv2sYs8NQHrUHfdlMQf7Qu5VSrCbPNIWDWzFO9F
WFWyvUY3JzzFwxm7VGoHi0L1fpPdlLBlBOQUbJBqQ25WLg83DcTKEEJ/c+5v6xa2
11xwVWOOzEMh/wE3vVT0IpgnT9lrj08/K1IjBqMYy2T2dSGrnQJra+0J/HqEsrZs
z1qeF/qCNdY1KpY9oEI818sGA3eSppQcnfjbqNKLjwlxTbtSu4TR4LnB20e0WmbL
sF7mv5fQMfWltmBWWS9FNVieOpJbXecvgl4dptOcON87RAUa5mMRi1UjFKSqx2dH
M79BjtT/DIb9su8KP8BSBS85e1kJ1ZepL4f3F/Db+35IeXe2EfXpXj3jPCoZzF6P
+M/gtUTfXJu2ycbJKPhRWrUl4wQ7oEz5oFg6/pLRIRpNkQQWiFtwfKnORazVlOPQ
1N4FC+ZBWy67jmsChZUt71PMbVzzpuO1iFzUxCMhfdTnoT7b+OoM78GOIU+I6q/K
HOTZsNQ85YWE4Bvzi8ntt1O9w4PGW75HxhRr7NU300ZdXVv4lnljs4/2ORAs9/7M
q9WD6W8A258jnmXoqS5204wbeDS0RNT5BurjUwW5F+s++SPAlTZPbGtmlWCn28bM
tMv20aL862L4g3JzEG2nADGyLa6cRI69ZstbsDANESIjzELejfUwAU4sEWhHeXNa
mMEmF0F1eXK52dR9CJ/8cs53fOcghnyyitmOLCvqftuEarKIXsyFltLpTuKtgcxg
hU7gxV+QwvVtQWLENAf3Ha+IeZmhc9pM8vzaj1lmW0LlMT/T8gnEjwFeC5yT3lZ8
7d/d2NTvtqEEL992jd5t+7TINSBAv29Vv2DrggUZ3xH0jcYXoXRnJtpsSG6jq7rL
yc0fkks86+ZMGP3og65ExejsfheX1/iWRD7GYTY0zEERX4vtPGTdkKUhLvWLTiKv
7qjAojc/CpmT9fLMk2JRzzdfucEslNtHx0QAiPIlPYcNDypHFJd8ljvKM9S2VAVq
4m3N3r3ZE2xB45SBsKVeFDsOndYt4n+0w8XueuKF7yljqEjHw3MuPpWxSDP363QQ
bkRah3DYNc6yyJDXvqdqENXq0O8F3J6jVA/x15rfo+D9GsaRTTCV3V+A3dSjs7MP
UnOOePW2eS8jiYVOBwrwor4ohjydSVJzMufC67ANaxBKn8dDQl7zuKLLUE2Huvz4
2V6FnhN+Ja+1Qy8ej8UBMFe/i9uR/z0Vrp80VgCc4dbSaLOXP6JmQFiho7Wsdkzw
yS0PP/g6NsFAHXaC2gReGLxV+B5XLTq6Yeh3rbiYZ5HVPh5YO68B1YFjI5nZa2MO
1UPsUSYcAueCzf99sLDgNKrvzhI4YZc1FMZ/8v/ZdOksjUK/tz53BMGSa7BNwt76
yNUZddznz49aNOWMrThwQ1zkSOAe+E3MYUpMn8HQs3GG2XTotnZy7ZGrykbSsi4q
IrtZr0v59jGill9IaPLauLPfF6+eNgVSK9b0AdpbZJJYoE2y5LT+s7kFfAj3Vce4
w/bLchADdBWqhXe4uGqARGv7wbQCZbLzDVPlrtbiKW+1CsQ2xAVUg04gI26JTwSG
Sx/fHFN2dJbw5cTfFfQaQTzxHDm8aBbymSLHN7CiqLNPd3tgnS3gn0517JbUw88h
za0/nYP8ECVLUrQVjhVXqE5DEERU5tuTAlUHn9U0mUBeGL2cEISaBmU1csxj20SF
iNHEpah7Rtf8kiNQfIMGjxYBSZd39nfi4VhdsYrcr4YRFSkSTiZMMgmmy/Ak1sUg
F3naGIbwk5KDHC7CK6GsqgiPjwDcpVqX+OYQMT1O63mZE2atk8AlUm4lyU5QRnE0
Z04ECC5PRLEv68NrDoAmNPpmea4DimqHWr4kh0uPG1P5UOkMYaR4YDkB1mdgNKAC
bEZ2T1TUNtKNG4mRwhlhnpNpyYZTJDEiYZPlJadCFTxATISVf/R3qWR52Y6fYC5o
r+F4zeOwz/bVfrTr1RAMztAty+VL2NwVQ2q9+8DDO0+gAu+JirsrQaNwUz/PE/NW
y0eJ8Hsg1Qj8Six3rYBlX+4VC3QxaNzp7gPsQbqVS09cPDYFpuvJEl5NFu/Ap8Pf
rlZSxE6cfKFTzPcqh6LcwdItDE8VDkNxgY051LM6WV5ntBlfNGPlTTIwrDWXr5jw
B0+g0MwiWb9i8WEXPJw/AcEKCgHaCJlI1TB/LScsYlBlQylhYaEEGxlSBaJZ7+05
J6j/fRbPFA+WRR89sI6SOFfoaVgKKaYRHAE9uVvIL3qiiLa54kG9IDS3dVoWalFF
sAEEhGtN/REZeVhFqTpFfp2yfCYnjOSfqQpvCzap0SmfcN31Ya2EVCCUfO/ARtqL
KlIRd3XWVvu0TMB+PJCTqLpMaJXcRWVsr4AZ22ppOJdztz+vRwXhxVTXQewGZyIr
I47zfcgCVQpIIR1px1uahescK+LidII2r0GzA5S14mkJZFqcj7XYyTIX5zgAF9SZ
a9f0vPRtBsKO/SaeB8Lh+pECZSwFlDqiiLSCq4d2pIXhHi7PyMS/D6kr3k/aNNVn
90W4GupvUXrlUMTGlB0Je7A1sPzk1JLzOmWeh/CRsJw/yAlozP+afjT5Eg0s0Uny
PUXC07QeNGrg26yx3zwvYrJQuBFIVEIODEBvsUZDYiULQm6j/FhrTpD/cjO+zbc2
pmQbAcoIP2/7EPAvkzsxfEMzP67KxiH5nGPMZU0f1ggqhWLiP+GGAl9TOntzGwS6
nN37qZb4XrekXv+lBOaE0EIUAHQHhQJpinEzjkOxbxkknaV2IesLTxAROBro8IxH
xsRgNq77I2ovqr/xdGJ6pG78EgfGjYk1kXS4sCiKUaXLNy8MDi5m/KpHBvyHuY9Q
+JPA2vPGgLgbLeJis9xDihG+XUz3tsJ/EZ9+vbvxiwYKYh7fcgn14efvKMLKZUcc
hkBZK85WKlJ6niNVHRbkO4MwS2hdW6sb9g46MfaQoYudDno5MdndGYKZI8oC4feI
o8uqJYkm43eKO8SehXBcBe8EMngAy4aABWVvoSzHbsJQ8eZYy4cmrdzeUzjpeIVH
MGYv7qGXPl9kYdaUOVpVBnEsBnbDpIgrYMRBM75zXikHkHn0kMnViqJt/SOGJMyA
DXq5cYiSSAUW8M42psAv+A76kkKWVhhtzq9iDodMQYZv5TDz6o2Ub/CSKWi2/+aX
GJA0AsOLuW1eVQQKY+w2aU0K/q7X8ZTgKXv9l+ZtyQelnkggyMIRXcLQHGfAVcUH
EE6HGzOs3k9OkPkeDOdKYfqJ+ONJVisx1jZWQxhGbnpvpxtrH603bvqDdDizaLuY
ui+EE30sL7ohjNnn0OGuicj6hjJU3WYezCgdHWA71IGmcFz/jQ/i2WeQ8yb1bgwh
sD1Ey//IOR1ExQaz81NckvQYzE4PXChfDVCrUV1NhfQ3aNL4Pk7an4ZJtoU4+oN0
ji5aXgG9PlVt6GJioTWUFvB8b1PFf5ag65GKlv0NA0nINGhaJS6WBVJyoEiQE96t
5bKfVaWD4lIUohFm6nyB21GdEL+xeceuF+xHpRY9qDiQi1HoH7S1ArulCL5w9q5P
MYhsjiT9z5g3bTjRFHUWjnF+vwxCEnWAqpm7bTzT9DSmzV1xmlgSjXduzW48PKd1
8H+8AHIponGGDt2GPv0rAeqnWku8vA/MHsibfE+OFDKQGX0+7OJx3s2iXmU2WIlo
dXq1A/z52vrr1oCA8I1V6gEHzvaRmMfk9bCa/q8JXaC6DNClGeAn7rj9UMwgYRhy
cChSAlTURbeIQcLpoJRwqSOu2Oz3RIrmrGbNrCfT79L2Oy+Jndb2uQp9crjQBsEE
DKV0bt/LXK+ytUp6wlucNUed+DTgovc+gDDu6uSptOdevS0KxZiq2h2YOcWnFb1K
YN76nfeDf/wiA41TbPQrvplFj4WYE8pLiQuvNbuJV3osOQoLqyosvG9bTaKMvZ9Q
C115Epv0lr6a+ehNecibiohOJgWittUnBMPkdMiypMdIDb1fszA1qnsMWWfRY3UI
xHJOTuJQxGmWk/a9JlVN0igDHQpccyLuc+ZhoxSR2WvJBUhP0JBE5qxzwcCCYIed
lanYjgr3LW6eTJCVoC0QHRKIGxATTL2OyK37cinpgXYeEjHqh6u2nIsYIDGeFzZO
/bF3a1jkR8BZbSiYt64u6wR8R/wGVuSuqWfau25F7aDpqmvBl5CM7Y3ya76Uoe4z
q7z4yPc4asZi4S2Om9pg5RNMz9tumvOSxrxNmlCyvZBSg51lPgJXJnvMMSMZA3lf
UcEuzknSSpzarYDDQvck0oGOIZiKnIqtAaeG6AS2URvRlTfz9V0EaaTHe71gEy4k
XF0w8nRRhgNIQ6j+mZAEVsnlNs/jyI6mPKtc3bmV/oga/3hl5MyDsCp78Gn2uD8j
ELWmV55F3SC/YmkD4ALbl7f1C9h9wsd1yVnOsHsPfrK0egmV0S5TixOI90ZXDYYG
gUd7N2vYfgcUQST3oSIIjVoNHQfXWaO2zf3lpsnmY78Rt/zCzhdtiyr5KSaFzwPQ
yX5ng/cbElVl2p/35uIBlkXu4mB2IZZzAFxHeNo8X2YHECaJi2XMeZ/oOB7spO7t
hUg6+/rQx3zpOHlnuPmVWslMyJuZHn0N/3Ki6w+q5dxvjyimLly2xhCeGt0OetA2
9FhCTrKRi6//a6Uf17Kf1lqReq52/itzED9LVtxUN7k3EqgMRMCH+OKAyEJqOnGi
sjUsJXrZ/XqfXi1FRrWBNVPLZH1h6c/2iAITPrCZU+CJTd0Li1Eoo8kJuPhxGzKe
tr/0DtwSpvAypXrkInGIn2wrBn5G4Qi2tDVJ212vFI8Wb6pYIvvV1N/bWDmhbifx
h/CPPcTyRmIiQ6TBZMfX7JJD254m6pRrG1gDzZpLK3WXoq38OzDS9bjwN50nOiJL
g4J7QJIL8Pr0tmEm9yFwrXCdCObn56p+dG/nB09Un2h0L4OgZ8+QYuYzlH/cjbYm
k1dPeYlO581MRo+J3I2ezRHc0acehq7ybDof2lX1cUvaVbkJ365ibvDKrlFxVge0
wqYrdMi/LpuENA8JHhVuwaR/l/lQgFaobzfaZZv/as2ROu8znGtDJk6ccszflcrr
9BhtN7Cewd45f7LSRJ03vd9Oewhx+hW90hawDTjqPwJ7enVUlOdq/shtkc1LhBVX
gRL9nC6UXUB13hOeXrjAOC3eCCGuUJc/dRuobNrptoiYbhQlZrwyYlVAoRjHNQ3E
wubWxy3oYaqhoCv39JmUUW7WV9fPRInTxapA/SiO6jDbPRoRK5LtDnmi16YsuRZ/
tScrBKRfdKFzwY/R7Fj0vA44tzkmySzJZYjCYvvyxQsPZmEHz5Azx6riUyfFlyon
sGWbhEypIdAChwTNMjMhUn5ItCOTEcIF/ZiADNxufM3VWuX5pd+uQ4K59M7/Y8Yh
krb7rVTkbMNhe8m35bknT49Nu0YKTCMEuEFSPTFUJje2iM92uwb7nbXzvCvlqxTm
FDJ1SjB2Sj9mWgVznwaj2G59a/nS+NQtZ/cqBKn5SzSTyvh4+jSOgK1zmk103WBd
cx3cJRZsG5hWzQhj9xE5vhSlP/7ZsXd+H02BmCKYPjW0jNTOFb2/2JJf/XRlXKsT
V5s2FmnAz8cxbQMfcux71Roz2oWMP1IvwH+jPCx8p1flMl+Ss7L66hbzgtU+bwrI
5t/3sTcstP+2SdVwPaXHo0VuPkxav5jfZdcRlHznXFxQk2AEOXBfHgpiHTmfMfEA
cUHCVu+jQLz4S7s94jdN+WCCmd69CpA+AS5ry9/6SBn/ZYF2WFYLPMz0jG/h5XwL
qqXKdqT0zWEc5IjuLtVRZ7XcPwimBPDEppprODmo3hH35Gek1ocg2E3OhBe8gwr3
HUbdjnWePSggLudslZroQYrYkMZv/jenjDzynEJsRpyuNSbgM8c5+/cMpVmlhK14
GuKyFoL9SjqD6Ap9HhD1mo1YB7ndPyY0DnrcZjvwIecKEnMAPSdcpo/gpyxoD8P4
31sMi0e4s8tqOc1+GWNASvxVV6iHbkp3KtqGXHReGSKUBneRIBx2jSyQ9FnaqZ67
Gyf4yxk8fa62BgK/xE8tD5PWhFkm8SqGiXxs2NmCn4KOTBB9mT++UGvS80FM3ezi
Guxa4KyZtYG1Nc+pWDh6wNpHeDOUn6n/pTsegMWveW6Q2MYCyu68Adzu46OVHZgD
rsI6N8ekKJ2jZEN2CHUqOZys/VsvD0S9VFhoXiJZYiwGBMLyi1nmG25XIMCixg9u
uj+2y1L1jHAxLkZTdKiRxf8taN8c23pmiAuJGxkGwQ2X64U4pdsHsgfsQqwoNplb
pKCpjFEAjPePhp5XNtGQe1AxZhfAwTMbaJprXGZuHS4zRKMtFCnSM6xyA3uhtCvF
eb+p+alS1qgHSXBKyxByLAgUxH/xBIFDwYieNd7qDzBLySOLizyIaPEfsvgADcuf
zw7hwalNomPkzG3J3ch8RbjuWGEluXKkE5BczO660YoRrxzJxGIkLSQOg3Hq5lEg
o/RDmYNjedHX4JmmwtnsmVbiNXPhGUY0VcahlXKbyH9Qwj6eYkXx6/3Qp1UY5PKG
yTyvw1a9QFg0Z5xG/j3y924KY15ClPvcKj3bELMgYYRnaDP8XmoCwoiyhmx+zl8m
AjKJ2NwKNUoONBLgtIOz2BcygBUholpgbfq8YUnZtSrzpudYz/dM1lEoNIpdVvdO
BdWBbTtCwXYlu8SfBOkznnByIbbj1Ey4+kgTcsukaqnQ82lSqnNLYnimpwHrZVux
q7a0tlPka9/0041+9niWwlRyXq3o038UGFLU7mnLoJgx3G/JbhJbI7L0Jv5SYtB+
nBCWdz0YAB7wCjB7MiE02rnZpw9SaFYLh3j5PUTXHpGOw7QUzmDWG6ptsXv1ojix
BywWwXbxD0zlOUbMQADLl3vET6KYcR/3Uq/BvCYWCdQulv5gnao/A0tU1EH4nyfK
kPFFybhm17n8OLTd+wuDSw==
`protect END_PROTECTED