-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
3g/KnsmYL4Rw9KBZBuLKYVyo3mQVRA5ncqSoqFyCbgVtFfY4gNe97gBP6y1Mi7Hn
4/SWAFm9j3IsC5vlBidbd2cwSG0jvt5Ym3klVhtn1N9qtRH4Yo1jow8Jmkb+lLVY
Bobkbuqj6vxkjtRhtYljhxu7pAZZaOiqPEInUeNvga8bw+1F5NaLyw==
--pragma protect end_key_block
--pragma protect digest_block
rUptM4WeAaQFoDmPPcrkV0k09oU=
--pragma protect end_digest_block
--pragma protect data_block
sNzMjyf0tZTDIfGMxGJwCxz/9SgQU+ctzDivjzNXFPCjO9wKWLNoT6qiNXXksZbK
3d3XSd14kNsczaBYy2qb1wsn9Z9lA+2Ulwxde5ijSFSyRFY/yUOsVluIB7q/RIGg
vU/NkkSOFkQsbib3Y1wXhYc33Ieh65mIe1Luj61LRJ99KhRugDN36qH+P/TvYBOz
m/iyiA1KngVE4mZmVV+05zQRPg4wul9sQeVvppl3/dZ2TUlBGynmDpNToNTgGky7
dXM3gDpPKiNq0MRaMPNN1TW+rewlqSVlslEeIm+xipZIaOVlYyQgxBR9ggghQlne
VfEf014+nn05LPpI8LlxOzwBmFjlBgHKiaPQf4AWXdHBNapxMt9EkdVw3+zqLvp9
sMhmzpeAoA9xFAODDgFDHc5wWb7QQa/cqzVESNm6nDuj58Z8plQSRKKtTmuklEUD
AABth5QKUJg5I1VIMpYQXqpimvc9WixTIih6/oRvfkM/3PPew0KtihFpgFKaqwrv
D9Vh1lOwAwiFLuGL7uBnrDy5SNkaTlghSsFtJZs1+Npy2Hq1JD3CeKiCKr7TRbAC
Xadee0QaTZ8tRvkR6yoTFeV5E5xdjYOSBPby/OAXY6DqHTgVVkpE72x629PVsw6d
Vy50EYkSjfrUwkWNrAA0Zd1W6ukI/v4WHvNhSpbYBoopo2CqLhJzN8wYJJy/oNmq
pBtWvf90A2Bxq+EQ8iEnC95ppd9Qg7/hZ/RtE+29ODSb+qAHBWa+em3t84K4gHby
NNNzBOuMKW7KkDU7l5yoRikRh+vngiUw64ysTmEbWw/JgSztV4GC4MEC4JQe+7jK
7LW7leLNTc92yf2zahm51UcmlrsrurFw6QJrAOh5NzLu/jItIVPzIKORCdpueJRp
6WGAS3A7TbyPHxBoycJCTF6HAjAu9Yd2H9f+bfKdZGS3nOxppARZ/HKLyZNvMhnm
PU79s1me0zlmr9fPP2DB/v9BO3RipY1jGUeYX0jDnwB1HJWvOaJLaOCHEb6WA/Ds
rqevJYhSS/MQijmLCLIXh6qQI9ad43GJ4SfdcJmXOVXQrLfRVSJmUgj9MY10NA5+
mnYl3gGbmSouS16XhE8oPa38XKUV+dk/2IDpSTNlx6AOEoEpBXrbKXdar4V/l/wZ
E2Y8eqWjJYNoSflH/Bkfw+pNcOTmbfF4M+ljQQyrR1em/lqTxe3+6PSJ7yyXeMqX
ERg0zczVUs0/f7O5n6zcgH71RTHuUhGE+uvsWjQXQJgPni9883QvdtvN9k44ZObu
MAibgQm1XyxcLNPR4Gc4jWUQLdeh1/C1jtuT7hnR34kO8NOc2DMKmQSsUU3r2ouh
+0w4dhLmzR7TgGdt/8mZgLsqN678pCIATS4NQW19ZOTNtPPCj9nHIR9g0bcoxj64
FOVMT/MZ8nly0GX9z6TriH0spGfnR8DKBUY1rpm1tudoWy3K+UjaiB9YbM77gUFh
Fy9J1Z1eVQBsf7jADIzcVNG9CXrT4/kvD/dboRVGuWgpn3kHYiD+z3me6DG9643M
qrfh68Y2EmBx4wacYB77BZeala7GKL21ozOyBsP2WxR1ljGonxX2PbifKTCzBhdd
oJTlJzaiexDpJWSLDo9MVu3Ax35zdfz1k4sFgcrmNs/a9SFkeHAvOyeCn3ROgnyW
IE+5bMQao5+UZQ61B39wsT2QP2x9XHoKRcG8TtSHauaPyGRxgp3+UmbLV15K5jqd
oi4DVdCUzh+Yo69UU6RZZcD5jXtEBh+xmmEkIXAvU6YBYh18u4aL7PpROsJxpl2I
4/dcF4fh3gCcgqg5qKd39dG3v9zVlVwPrrOrd7J7pZIX0kI/Yocfb9kuUwNZXshN
Qwn8kpk8elh7AdZl3tUzxS53Af66miZ1SMm6ysv1vqm10uxajf7QLuCC4yo9mkcD
DnNQLVUVpTEaERVCP8sQfpuSYlvl4hzuDG7kViBjbNk1z926W3EPf1vm3C6vJd4w
Xw/GQZDDsdP12T6hxv8A+x3SzpsXj4NtRwWhAgn6C0NkWo0qKifdp0lRfxrhajNO
O+H7WoSp/f31KgaHaQcRA6faku8QhQUhpdrpggtySaNhtbMGYtPeTWWlm9ee5EYl
7Jr/SRqq0ZfcRvAAfxYPhXJFf4KrBXjN/6CXxiujnPnWsXg3OpQwepBOzYHZ5zZv
G/SSdbneuZTk63Y0+E9Y8DyGd73I/zMwi4tjzH+2DUVvLM2ibEdSJ/PI5Jq9+7js
hsyysFZBu2AVzh1NGUV6SfHvFuq+IPlhXC8CGqd8c3feZG1e+6O31QUs570SaTtc
nFZvzxeN6dzeUY4tAFsddDaN9Ro5zHJcvP3h39mM+Fz3Wmr1WlszdsY77xPx4QWu
HvdWi/VzSbrorYysAX2m8opxYP3o9vHL61lKGCzHrv2SNv8rd+Im9AeMain7jsZh
X+tFMwt2Oyi+8wtyyMW5V2/lqkQLnZ31yzYj7uXdNR1EL5X0vUCpjgq6FzTBQnf2
3wRjv3nVp+4H0ZiHllMbX6mddZy9uiyQKqH5AaoqLshkIoaev+iaunFhYp8kWal7
syRNgMwV8621Sw2HKinr+Lv9dHe1zUmk+PP1KhIxViMnscFM4QWPnkzAkNk4Zt2f
YGjQ5H2v1Syi01O9wlJR8nLzNKxitXTkgZMf/k7aV9Q8oYXS1l8w4Inc/eyaU2pb
kdydJJzwzHifVDJ6/eAUVEg3wFUfRMyuPfddlepVy67fzhZbKKKgEcUvpJgCx5JE
2ymcAjL++t5OtdLMIj1zZQbzboMjasoeZ5+VbVZyw6bitHsK/JqLV0CdTQm6AAM9
U3RlTQNoJmGngUo1Q2JL2KEerAuBNAiNYlWUFWlYv56NlOlA3xuiGDc/XJyVJKWL
qTtGNV8CuZ6LUR1xDoA7f5cbC1RAwST/1KDqV/LF6coPkY4gd/rfazXFudzJgj5W
fHkoVAQE3Dt1olTa6doA2HHpFa7xiNtF90laYtpXoqm9L31bZGk45Cx2kLmSfhG2
dMFdGij0t8tmCPOu8MXAnmknwwwyduwb8wxaKowO08688cUDvOU0ldVMu6jea9f1
LGLNBZuvxi5rNwisD8HjRQubukInLcnQ614Br9RU0YzV6584qChlL/v98YgaT8eW
KJVFvL+rOYDCELQtAK6NfFmEqGgps1DgQHb1EXI8A1FjKrKF2JjeEva477bvsWNS
dV5087y1eldZXgvWh8mc8Od32hDbUEHURk/l3HUT2kajjqWV1t6hSYMjGJPLDJq1
VLN5yd7lrurCZXKwNyWdG9zYlfC/7kRfijlyA63LKfAjZEkszH4YP2YFIk5aHpjX
BV8OiOWpUTwMxN1qa1NSw0GH6l9j8gLBRlkFcULq0fhHQV/+4VH09DpvTEo7Oayv
YcN0BBhWRc28yXTGNre+GIKwB7VJEpljSsldXHC+oEeRMNjuykibJ9JNvcC6WCtV
BastcluQ/g+5XcMt4XdhiyeSM/6Ng5LedNQ8VFMNQQ4D6dqACtXtNoXGnnL9OtZr
p+olrIKl3qnoYvtImvNOTsJWHLVMZdg5nHYM3J1gbg3kb0NF0ac+2MKKVfUNd/4q
WEh0SrIJ+OGrSssl5J24KltzcirMTke6kGJVgXK6LX0+ij497LoJuuCz4hZU2cPl
BtWaM+PBt6/fHCrg+4s7uRcQLQ1pK7+RJ2ss7DAg197XvWO2mdDmAcbD8FhbkSd1
yS1PeSJWlHhM8dMPKzXK0nZ09AAsiORBpBNYs/hEt9AQnZiEGds4hFzL1wJhNkRJ
ycV2/3bwaqrwB+vzWJAcEMGsaVcUb2diCa0DFdCV3bh742hM62UaBpuU8/03uM9w
hveROcbbsK4PjC36ML82xfS01FQI94BWIPVfEYaWsxtuvNkMRmd9aW7WuPG7k52S
iiTSql3bJ1f2AGn0IRRkMv8/aBi0IUr5cZhq/ZZ8LRH5KFQ5j3y1GmxXnVFG3jUL
Ptfsz/HUYvW18Gq80VYFEsLk5zsWxq1ok3Aols4LG+iA8WzqBEafMjTBUwv2v/I/
gN59PghIUlPeVQfEKvyCTmEnkQVz9IUjQ2gXO5KMbTh3EVFl8hHua7tG6+0F0mzZ
qaWMLpUzc6J3esPngCJ6a9JbFwMGH/ymAE5KQeI/X6oSVeS2XCtMQ44pu+EBeeHA
SCIMF4f2NQ52z/DkoQ0la/KgV+yijp2YFpYM5GM/aCvsEO8a6EpuUsKFYt9RXV67
+Jzl/zetPptBXUWPU4kenkpKIM2gMJaJWGNhEU9K+VwPFLiUFV/97/zRcy/PnNxW
h+VB/K/hC3CBdW6qb7ZUiruLNcF+CWtYKf2atWJVt8LLu2xkbaFZ6MSTjseEZMtM
ofR81RoxkXHBIAjq8Es2KZX95OaJSI85ZIRfXYWwCW/yB7pJek8Pa08IQ54iAByC
0isUzZwA0GJL3BXD/6TmF9ikqjWTRKq7f31nb4MYvCnicnUmOxRKk+wyMM+raNOp
sIl0opX7Nu0KeNdCan6RboqY+AMqdXCMLz05sQR+m1u15iDIE4zwNTvY/9rjJa76
r1MctNwgLi3bVbceN6zIDIM1ImwEViaKxaxtkOwv9iRvy2/ez850mSd2fpid/swF
jxdXrU8ympM3hxUMKuKW+6QQ4lAd+kRiFxzXPOmXdEf+P6NqJCE5VY/tFT9m23wL
Yax6VjWvjNYBZQOLRwBsIhcwF+A1mPwWz/xGeSyi2aYmjGCCtvoS6WKLchiIbsWC
RsprrdlHOp8yRZrj3NrgCNaM3GJwRpmzSeJkUqHTZ7ZGQtiHhOpwHfismCS4X2RB
ziPwHcYMoMVPND+/k+2uYgw1pPLjdstG36jHo21dwdYcHviN9BddCC55SXfTbKXs
KGN9OyPznCencjBYe3knskja6yTHofzzYdOZNrahhGCNOgQCv73bLgk9HxlGQtuY
OsmRi8Y/M9PLH81Ls9O49smgwYe+q+62IB3q9maYn9nA9dRGyNQ/F8bXYZ0BkwP+
O+DzrFnKwroJcKyGL8Xhg5RE6EzezGXUIyXuMe3TbYCmKfFOwkI7Tcxp1xxQH85T
xeizgWlOJ+eK7+Kgcjt2gBe2H2ywqUOYKnGT30GjbaQ2jviph7ambt2kWVbmzghk
K93AT19471axsyguB6NL24OTODETv8PiWdpjCkBCzad87VRBm/jH8Z+hzxATJslJ
lUWkcy/9igAC3EfMxvYoWkT7xeIou/m7Ol46E1yXfTfnAwLFNQkv4yuSVCQyLjwB
4OzxA37Md5nm3dv4COFEkyBHQ/EhyuMjJvsS+lq54Dz1LdG6T5+/pvpyHsQQcqv5
eGF1pTe+Be0UMBG2D386n4rb2LVWUUsfZmKnm6seARkYmK/bmzpeWGBx1QMv25o2
0anGWV5tTkz5++l0cmgRduvZqdsIulTVC9FyUtbL+I8+/Xtcccm+fMeXjeNPFrCM
/FGz+lDZUmaDnS5N6Q9VnBUVoFcBC0lBnVYWN2F2EGinf/1LhOL6saPoYc3VG3Gm
bhNcRk+D3vVIqKO3J/tib4FDSddx0EMjw6gbXGoNudwjD5wqCpxdQP6omyMV9Ja9
dfnqb1d3E3zw1By3sOSv79GFZHKvGLjDUYiuYavzv4Lg1QMCwdECqlTUUhJjKaue
LIi0ocUQxrKn1LTf9GgAsb111cjEPU2Q9xN1Uy6kr3FH1VSJxnBorsgPL1owCFKR
dCU5NWndtLZ8K2qx58ZIEwvlFS8qEe8C9DD0ZF4YhvbGEXBUGyxMZJCzWmxSiRS5
FqnyYr1BLe8TD9jJ5n8nxJozWRO/4PdNM/quW7Cbdjb5ilj3Lxbrao0UPP3lVSaJ
lqxFONrjolla6DZRbhT+xhtFNqM09uzoj6IM1D/+GplJN1ogGk3+EelftG3CdHI9
27j1id7i4/J1MPJ0a0WN6AkxRrAUwYtC4doFQFuP7YM7a+zNteYJkeDWd4YDlx0P
wdzqNwUoB+MCbeCMQBpzfi4behWysaJs8eD9bDly6of4ArwCZa1r0v9Re7+un3hL
JyZtzettCQxY2vZJleQpI18Fad1siNHXNq8fM8mdwulMIF1dfXXpjZSkTAF07PEJ
NSayqTiyiPPQ3BF4iel+MDG5+fp4E3ad91KVy4YcGbHjKtyv5D5nh9xImLheWPs9
2X9cpluxdle8xUJ/l2dz6KqEhI4pbgKt1HVm/FNjjk4mZrBbbjsn+oTIsgXit6ou
LKFv4SiTM4yN+y8oUiT9gKQkOU/5fDEYy7/4BCfbjbRBS8zpRvsEc2u8sl45KNV4
W4TIvVvDQash0yiAY00XsjNVxg5dv7KjS5uhJWCAnNCF2ScnqgHsPyjPvSBf7LN/
ZTfm6MaQ1cqOoViAllin1KXzZecdc+3rrUyw/4NaenuSl7dRcLpac086cXV4iEYK
hjjTsarDLWwQb9Qhllk8E7Bsv3rFmhkoUohVZ7wGQ2RwpqUYlqMFs5HbyDixjdYy
GLeyLWJkUR2uEXWW+NyYOXo1dSTfsodnkko3a+OXRQWKwluiacKMmg1hpfsYl5J6
mmbtvIZeorKyVRZ/YmS5Dm8diL+2YydogcH4V08DmG4VxASyn9/fSz5R6SN5t9JM
pp5TUGYohFySJ8sCqdeg0g0Fp0vl2K8mrRMgACfe//IkXzbqDYcgDJLnTQL7zmjF
HBA51gXjw6xbwzRzW1QWcnX/10Hf2vORzRKX4U5qB4FrrRR/4Wp0JoHOpEBv1mz8
sfSEpTRjCtSF8srhXvjrp43/Rpao1WXUy/U2N/1YcUjV7qDq1tfpMdsfnzCR4M8D
NGW/dlH3eVf0CY0/sCdMILoKjjM46egDUg5yD8CHZcBvLLde6IyPoRZ18ZZOZaLA
8ESKsM7U67qW3F0urMFu2UVtuJOEI0GGytWTwQkBjiJt59WnF8Z9aNhtKzRtg5E/
g/dxIPFMotEb21PVBV5jb0v+vvOnyLgj4XnK9bgjlndTMiliGKocrJxfwkt0Glsk
iEwZKnuE0VD9rMceFluCZxUB8U3Poi/91hFtD28F5YPsEjKas+O9VPpi0okFOgj7
eCE4DHYTI1jqa0ASX8hJQ43e8yP/feSa3wv9izRL8AgyOmZ6DX9SJxBtMs8gmvdg
lFWXE7NG899SlBElU+Vw9FmcUfHh44rwVnk4fdaf93X/Y8LW9m5rsMUOEJ4JEtV3
fxVkX41/IUsE+fvsqYGjueTIU7sTBasv6NbJY09NIKxau8sLQdGGYotnOjWZbQeR
fFY50IofgInnSNgpwcH6OqiJbEck1udfC91Eqb3n+6r7n2auM3kD7k1XhVI0bbmx
YSEz8fku9dU1ypJQEqCrXxA5al+jpYX54YoJkKY4Mh3vXNWn3L6j8qMJSz2rT4hN
JT3GsCsAmWFRrgahRQvb1SoSYw8XXcGlKBk1VjsipKRfZLEnyCHJ/xExJlfNXojZ
v/4OEtdAiW27aPpjpXzTF5Lr+YUaP8PQVYe75Bn/67Tvlje8rXW6DZgSMLdj6vb2
ii89vzevKC/u2tJ6dyxVuUEkPni3cVVhdQY98R16SaWZrevo/OXEVYeRsWAIoI9y
Ts8bFNQ7req4WuxCt/iAX2CeUW/29tR9J9xCrIP1KCOLYrNQ0tZLAjdd3YW6GYTs
HfP672hz4KcGt2geC6vpPukVA9v12kRuMYrnWtfLapHUJUVD2wdoWELO5Xwpwfa0
8lZPqspwYBBiOgtErm5Fr3BCTS3K8DOrfGz1oZmdq+H13y9/p9FsBRJm9vVl3M0g
HRbGNALokMb2x7UTLQTB/KD77hsUFjxIDeLjj6yvfcHa2LDWSDQXdu8neBiWqeKn
Hvglj0EspUZv+KfqMx8D5oNx9Fa+3OVDDaV0DNTcapDzvwLDlHbijHrrsubltEii
wCsuB9CWrXlbIkAvSrC+3ie87Tx9yAfPXJpNCWgkas158ZwqtssCIjMQxyx/wK1Y
wdHnRGzbSJpBNjudXYNLG42tw6CqI5Th6cdo/WHG/xBpHIr7/K/hJZQiwMFUFyWQ
fi+RB8AOSlvJwD7sEoI86hzftU6dWp/pZ11WVCi76JdDj8qgRjXCPiqWrTO9Mt/+
VT3IHSm7eFzZwVtfns0L7dnL1e6QzFhtRRoTJd2ifEYWiNzDWAy/tXo6Sn7DfNfL
ui9WyMLAql7ND3XndEhmKJZrjWaNBWLQuTUqC8DlF/pDOJmPmtTWOLLUXTzkfGjS
mFzmWdA/JdWBFl3g96rNJ0cF5fc5rEcMhwvVIPspBYkdllD1q4AvVvxdR7rIHge6
PBweWCwodJdcjE4xzyphWSzoTVHvEpT9rJquZoLSuCn1ywtJYJ2KfMAy1wCSs+IV
qpgwI2vQQ2Tf/bDxPx29x20x1Nskq+NMTpfKp40gPtDBoyNR+46goiYLVi1xNhy0
xKelp3/Cj+q3Zi1A9hTV1v3FpEMrK62AQm5QVl536cZ3884PcAqdz8/HfCPPYQL4
H1aEoSB+tuNeFhsIADpMVg5o0iqIw2pcVFROYLusuCj18SX5RsuPZ4BrLt8eV9jm
cbvpf72QG8RA+yATSVhaUc2ZP+80nDen8l5eNL2pc3X9yvhx2q3nXPfV2H0bFYd7
PEZ0JGPefmUhOmal7zofixED6LWnzjdF02yOU4KgK2qODGal2wQN82zyoQ5Jbegm
OxD+2yTdLtoMkexAuZ+ABrJmrvbbnqC1EO+7g8OPhSKRRn7MpnlMna7pu3sMoSv9
GB8YH0c2YslLZKOQlg2J93RFcIvhSoUw0moudJ1f9gGTpCyYI/4igSkLLkzVqeuF
bKU3vOvmZRd9vRnKNA5TpRbcABVbEMmZdNaL2mDdKUR8iKTFYvRn082nQDaBIfaq
a3yclzOp+aFWR6t50GBUFUMrXGtT2WovDnu05jjxXDIpDhSEl81UqjsHClJMLYvF
N0OQb/7mro5qA12rA+W9sTVozLo66gepkbcHmy+AHKR6QsVlvOITjebnddFeLuby
0rKNf59AZyJ2xnSzo4MydFZsivfeZYS7I3dL/YM6yW+uOqyom+kbOrqmumU2IZW3
ZsgTEtsgV/YGttNqzue8C+gmKujg7yCq108cYC9gIilMZwo4CsbhqtjXWRE774Gs
b8v+TB5S7HEAPuuTr2KAnyVH4bufwI/M5rbUqZvObMoqvmho4Awr8rAhCg9rH2Tj
VIYLkuYdJn6YQmxhrwsvqSYUV7ccs/ArHORUoHBLQGxtAB5d61aUpvihknIGrYaq
9hpqBn4OwL1RyaPMqdHzoQH/SgrNRfalBjIiK69iBe4QZVIXZFtsDw6qrfD8yjVS
Wk4gA6mTtsxU2UC3efNLltUsYrhkGGGWgUW7s4fq1VMCHhu44H9LfuFpFhW7N19B
k5+MjLXhYgtoaJcIr2m0oI96IZSz/y6pID9F9UXJNpH/rwpuNLCZEc34s36YPR3S
I9Bz6MSXk77dvHI0iiqIqHnk+UNQUfvhj0w39RkuCdjNm7DVtRdGNZOQAURyxpvu
ZmG6QLBPomasqWaapdNzVnyMHrgHOFymmPjRI9xb+fAVUjKxi7mDNjmkZFse17cC
E359jPvotAlaosN9Eg2CH9HZRWc6A1cjZUNDloxlP1KBD4Ctgo+lsznDWULV16OF
JS+B0JE+6/WwU33nC1frWvQODQtdcAYO+aUG3709r+Sa9U9dkjvB4DmXEkYyThIO
6oXeNMtKlfrQK7kLc+CZFZ27bG29t1HkR7glOIb2i7oAaRhTv8D6NammLBySTIWY
4l4DyuLCuWSlERe3t+/Cp+hFG1hTc1zY9hg/it9Ul4Bdqpg2RhJYVf0nKT+sPmDX
YNNGAXLaynGdH8Lc6HWQIIJ6KOrLnvBjuLqOUQuZO1Bdr2yPtK/n2FTXhWYwcD1H
RjQ2wbuXXShc4bn6GJse5JAFuqXJHbuqruFltEtf7xXiirEUycqqDwkBV8ciZDhs
CHw18/o9bk/bVtabh57blTfUcp1+ZmGYl/XoWhzY50of+r+Qmle71X5H+tt2VLRg
g979xP6bkLybTOvIOLMGxcGyIldxWj1PAHZOpP3GGGnJzB383fHrJNyMk8tF9L8L
3HelkPxoD0+oAy3C5lIDBLVbayJCFCOCwSPTwzNt4kLRyCoNUwXXqf+Z5KbVkg7F
a8PUg71fAt5KRu8N+TJLD+vlyPN75GLIlcHs3H8ZPdVN5b9BOasz8hVJhiaJFMwn
dM4Sh8JuB4AItaxU8NJlm9SWvs7/hqGgyNQi4mrRs1n0bGnaMN37a8TdwTamxX24
EX2uCvTkDJzHk1/+XHN6UHKEr3agnyJc7oIbQovvj+pi9mW9zW3ZMndIoCws8qBV
6LBq7+T4cY4UrJEUbd6+JWukVvq9X+4+XHEireRQ8xptIuPVr5RYDZvveNtbkx1S
YlALvth4OSrpz2dSsiBNJeIbnHPaxqYO7WYScO7Ms2jKKfqax9rNPHgAI1K5fLC4
mEa/aXA8zw5yUCgRKlzlyvkAS6SbOIBjQ+vdCmEFf/awHp9d/poTT3/l+wbBooKv
6p7QY6ARAicvc9P1qm+GOVJRNZiox4zLgLv+fUW33e+3r6o2+axs2MqhD9D31OLx
HzpS4IfSCKgx2gNklG8Qk6GmpKa6fAts40UdLDJ/RYXqnPrVHobYp8oUgIrNwpuM
rKDVQ/AjH56hzT99yF0XFSdLIF2Hl7a5gW832JYnhHKmJMn9C25xtfQ8y1bbIwjw
Xw867M+W4Q3+NO0D2WFlN5PJC6+Res0/FFYtevQ+SB78mFfRPysK92PZXMNjdIYZ
fC/5dlGRNXocEeeCdvLiOHZPEAa9VVRwcsWu6BlI1UZ23oc8B2ES/oZMG3BYcRAQ
WtVli8aH3GMzSRWh3QvD7u7XTxkfT3oOZViCER1qIsQhuBf5q+VYVjH2DM20sSqZ
+cVKJhBObSXZWWp/gj8/Thq9hmAgGRTNBWCEFL1cF/jUhPR1jDrrJlXQtNpwTbqa
raoTAh2BIzXN4Dq3rKigZKQ/sXXUy/ULPWpbUh7THetrYorBHQKhdlqLwAvjTXlh
KYAkpnjHOPIzTCU98R1bmJGd6HAyoIChCjfdiqyzgBMGEBVmuFWuUGMj41jzxgPs
qP4I2EvbKZggO+FH9Y/gh03heNnrly4dUCE2sNnt98W7vLt3ke0zpYRLuRJzssrn
zZCwPgSW29c7jP6NtvS9RYPLUqwgIrfu63z1vhGW0mCddmq1Kql9nhVdLyAWUsuH
sAZhpXJ3UpQEfb/ohShzl5rT0zzZrHXY293lEjapNFGUgrx+QLcCtZBnDKjMoPG3
w9rX/K/54QLHx1DLH+0zYQqid52WmDI5bVYfeNHRb9f88hI7Pz7xRkFQ4QoXNuNW
obPoKzUvoS1yinVPg9tNDN2T7L20/4sA1PZbkO1i2jnJit6Y175CLrpHvsrjRglN
10ttjC3mfrGff/x3M4J87b9+3HZS5JciSsItc2vePWqNxM43MSg8q3XEs9qVLhgu
yYPVlxOiNXbTxXQxX3K1r8ovvv067aiqXpCeybimH8msyFJzWM8oPizyUJDRWpRO
dIB4bEzBl++Q+GMax25dRN2av2Cgxl+tcTq8AnMKYYUIOn4twl1nfb9+2CAh9TWq
RffVk2DN7BonZrVzgB4p+jlAXbC7oe75av/k65neJKLFHxNgtkNiQDFkVfPyHtQf
ZP2p64Rw4kA2i/fmYxL84dn+ReoYY9VbzxVRHDWGLGxs5bmVTPhXFUV62fBUMO46
ppRJkeFWfQouoWLnLPl4/z9cHxpcpYVGXNfR37h750AbW1fALBbXUdTd6YfZJ8Gg
A+8zWJmkVB/kiAArk9HFHfuhjUC9f4DmYhHDAEXQ790zD3e9AjYgDqNpwTTdgMCh
BhPolfa9/N5ltbjoRZGlxhI4e7MgwtWqK8KvkYJGQTeD4LJGFn7F1SVOU1UCOB5A

--pragma protect end_data_block
--pragma protect digest_block
uoktxhI2XSSDUQw1Q4efWeJK2Jc=
--pragma protect end_digest_block
--pragma protect end_protected
