-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
MsfVL1TfKEsWD1N2M31kb75y8R8BggKIlXCIM0kCFDbwsJOeMcWA4KKujFeA39Ou
4TYlas8J0zFLQ4EkZxX5RCCt352Hwkah4CdhLYSXu2XtgtjlrRti3Gxhm3WdmabM
QMM1/wY43FJSqT+e3K8gXDxJm2cqjQqgvl9w9jbOYdAdiujCdRAejw==
--pragma protect end_key_block
--pragma protect digest_block
RlvdG4zwBJoyCXq842oZ5O+MYPM=
--pragma protect end_digest_block
--pragma protect data_block
Q2uSbU3a7jdbwF+Nf/ZGS8jKuVVjkiWn+64nJDmRLYUyOIHtZH5rr3wY08UF0ksU
Zxhjv5yj0AnLkce8lCYZijj7Is1Oep4EmJ72sklGeka7bR5osHKD9A1Km3rFxh0P
7LfziorDo2R+ttA1edWSYW56/Qp4WNmjSVR+M5U7cYTQ0WsbLrzASa+50uXbAXTm
IycVHKba1F80fMM+c9DiWJ36zc3l7NTHldEPHGy7psCTqQHh6Ig0Y6E2hrOTE0ZD
qVNJmZ5GHHrIxdFuj0mMwChpWVfuUYziyAMJaFfIE8YIYd0Irgm6fODl9bDdYcCQ
RK7mitnyyrn4W/2AODdmbj79YPhVbWZocBpDdMxzfkh+ibyBEe7uxQkjiQS8zkVB
NJOfw8a3J4rQcYVF0chGPqbXqVeFrRuaz74HGuBOkvsCc5BpsS9l238B+JAmziVh
3wZJdSUFm7HiT8jbdahjpvt7DPb2EJvXfYjzaat7r+fYGGGoTVRO2lPSI+EpqRXu
EnvIcWhO6DQxnKazqCb7I54Bb4sXfMlvxPCgBDnKRhxrHdu9t8bBn3sSV3P1rZDO
5Td6GzkHDDG5LA0m10dir0Gez2/ahYYYiu9n0JN7nFk5z2CrIZ1tL+IR10FTztxw
myno3UT+eJtfczkx1Ak9EOSr9kYTmFenJVZwJY5Oyt9L4zF9Gfn9xu+sFkuycJ3h
J/p8k7wtpo8tvZsNFI96WfOlc9HR6DotXoq9UKz0Z2B5InXplROFw6Yn3l9pSTkp
u0unVCAUW3frsdtHN+LFmabABXTMNrFi5A7QQxXodusgJ3gX56MVJiUeLXzDCc6/
vA3HWBIP2ZmzyWHcZR/hK6qaAIyDMGNc+VxkF/ZVDz9Ayqv/Tlq82xEs/Hb2E8a3
F/TN8T7dEixysJOAxGwLzlSZrK0aKPrp89f1EQguPdefIyYlM6qQ5dxMPcDlPX8r
OezNA2WWXMdpyV+n4XxkMDqWBRpvWqyGJR9YEigN93W/apqyaxbfocxhy7TmjAtk
ShmIgwCR4kX0qW/9DeBkIn2CXWZ4Qc66omisYK9NOdG6bLurU5ox6ykCS/zfvbKK
qOqxC6Aj9OhsxxtHtWvozbk3c1KU+OHJBDW6ft10o1XNVT3Q8YKJuWdv6r4T5Kju
4CftmP0kWqe3ykPWtCkrvmkIG5izbfDwtCrhoGvdZa6WRjBeLyKFDZZtt9LwZ2p3
ZdnuyZZY7S/EqPb20b2MzeqOo/orEqEvU8nQijrQ5edMfDD2fcvcyCuklxm0XzQq
17BL9LpKbd528HvQAGWGLcTuJbw+/vO/Ebvx+sL5KWLFsW4F9VRFd0pYLEO+seQa
AJcP314MoHOUTEjtJ8EZkDLi/FP4e16Tfi/aijErrVH/RcMHrPqoHt7DY+TuvFxL
jiGyKQ2/LoZgMU9+8+ROUPKLtjsPRUTAUDSHZiOHxywBcqokUJEiTCxgD2tHF0F8
dBMC2SHfsP31Mp8nUoqL3fbCqk0JWgRqDyIfLI8qCbGYBE+wB8cAVcXucTIstOb/
k8Wot6vSv+eGD11q72HRBvkZ/IOzWWUtqwCR1fxtvnnrR2ic71HiyJqtDUcm7QTK
ZSFEA6odYNlv7yzPYEiyQ8kzK3067En+Ko8/SappVxlD3exf9Ve7it+SvH1zspsi
5Y7tY+6KXvKJ2a6YeCsXA1ecsRXQiS8KqPjVOA46F442QoyCjEmLBHcJqfTkwilf
/5+ySw7tHSYgkAco25p4X5uVD4NXv6jzgBgsceKqsxKCwrGHujiVXf/KdRQ7EdHZ
iCr3X5V5Gl9IV7ShkmAM7++StY7g83p189/QN5YBQmf5VuEZjJckXPSjIX9QHlkg
GpJH8fdMnMeLy7nLuC8xV2VF6PIu5ujXrS1TECSUP4Kut/yGGPT4YHgDOO4JqQ11
8ldUJ+f1Umh5pDMMGRfj5MYMYJHB6NJVNwCuAkqdARL2ex5lSbKYpWIrk+nzeW7u
XDLtBJtePQMahJOUInzGGqVPGuG/InoD44SjqzMXgT5p0zCl2SOtSWqV/eGi4Roh
KJRaKzqwYu7YYGsmrfvR9NvypVnyIZZj30LAIeB4t0YpUfNAEoBGokhA6xr2L5lz
Vt4iG96Mo6uRlm44UnwI2N4UHnTO16QqzuyDdbkZLYnyhYfWpSfaBQpPpN7P0RDC
hrnM/dKMhc1bJUeMFAGLS5N0EHr9ktgdDFfFEW2Sz5hXyHQRTzI/S8F651SpfaZY
A+pemxfK2I9UEOosVSyaXWqiyWCAUzPyVhfbG8NAQJ2QjdzaMrB/S6syGUAYuk+x
/v5to3bEpwzBrxi0p5dUcLKdQQMhKSwsxzSdl34N19RAfe6J6tFaGxGxpZUHz26S
93uzS0iTzuP20TSF1mHsqLt84kATlcc8N5dQiOSNwg8Pkle672yid2RQ2fPyOtLj
1COConJDdcUhfEunqlnr35FG/4EJlv4VhAmc2kqUfVswIggd4S5Lo/jjqLAexjXT
sdmvXxqsQoD1Btq3GbqGk5G3KtDFG/8/d6CQyCJoI6UqWRUInNJ6U+vmoPjQdxo9
X6z0aj7FhaQ4DuX3CH9Ocb4x6oLdxfUtshr38nkKGTvEcVHstQzpq2GKm8axgMYk
YPFDW2YYFtfyE5MmzDWSUVpTP82rys1T5FhzEH0kzguh5ahiq+seK4X5Rvs+fhLy
GRmn4tudqTDRzEAVXolRqMsBCcWUTA52Tlq1BuELU8vWyjxPh+d11OpYcO4KC6hs
cWikiz/u0jNoJ10VjNeLG9kRVip65dDUvWkJrutoPqez6MbaCJZWD6/JUrzx3j4h
Tv1Q98LlV304+UwToymR2sjcqwn+uYRa/Gm2uhxYCAFFjJXx6h6rQMrnxuKzpn4h
7UzwaXMRcIV6jHp7IQOHMqxDcs96v1Q2AwuWXca/a2NfKXzWJiDmaPtu8e026aAA
xR1/xjSdhsrSbVjSMraQfkdTBzME7sP7RWmsTCKVSKBAkr2i0sNUCbWH4Hm1fETp
YYA2W1bywWUFcEygZwJd8P3WysPhmQ2PEhBwr5WS3ZDy1G6/GSoOn1UDuGj2O9ov
ja2TpNYkJNYdWcweKJor//zom0ocqNVBIBpU5mKqLUo2GOJjhbVMLjWF9apQz+uQ
RCoZAUdvnC8k422E7uanZMY3kT9fBuFTwlE4KhmuXWuhkJHqI0KWHr22QbMt3Igy
fbAYhruNygctRLgLutiYQxPFE/lKu4cVivHZ49ifbdPX01bnIwg/ks6HfQ8VQ69o
c5CeOOmjamcvig6mTWMjDyHkNI1vfhDouTyFeacrbiFBmAMznc1ZKx2xFrhgqNGJ
CIIBr0CWdCcOxPGF4xkVI/XjKIgQEO9iRLF1JK2A7R5nrZ7ktd4BjOPrAbOE+0Dp
Dg3s/wBCO5VTUvT4iKj8Pkfg5d/l7khhgeAXz2MIR9kp3srd2eWQ1EjpiKKupOIY
fILxiR4ozPpbN7QbSBy33l/J32wfu0QcMwcuTOAWrtFsny48tHBam3gadqkLA17U
Jju9q4VMf89JEehi1Zpz5NlYIQV2s26/MXYj24yhBVl63bT54pDHX6iU3PeRYzLN
G4v11iviExvHYax2baNmTPV7/wa9XPOi/I8bMNH8QqjeaYPFmlKmeZnoZgSk+rpJ
YLDa1G+2nDuisqi/ZuYrAW0xwLPmgJZIVufkGU1AsHzTfLrqVCfaMe++TsGQzE85
3x7QLOvxADJKTHVS4pwSzeTSCgOYi2lfDHbWB9bhdy6YGSIU6rs9zZb6T1pYwl15
7zSjrXLP6TevWs2wKrQv2G2+9fwmurqUBhpKZ02ulZYJjYndMzp3objRmlzt47Hc
2KEbMuAdKl2FuiKNHxZraBd8P5SI4/xdym1+yTPs5QXN+cjTSwleEeCWi67Ne6zL
vd5E2+ESk5uu+7gUIUG20IDsoqq9HdQClADZxivEO8q43wUsr+kAWte77PzIbKd0
DoniaK2AKNXDyQGrQ9v5YrgbZXGm6QaSGziTDUjXg1/jr9eFsqiwrd+huyC4JDxj
lt0/ryx6X8+cCky0Y64hR9Oa2rups4hcUfWcjLnIfeh+QK85S6Rfk2XRmhWovnMJ
AIBjtT/xFyhXOLSauzeQz/z5+9EkZO0mwL9u1BUpJF9vrx7UcZHfsBjKU6xGLKBX
fvM74QHH6VjDN78kUKmXjIqKCdIQzVLBZmFSEnXMXNUgj/+dwHIbb88qCZgihWPj
e/3oBP+CEi6o5Hl4M4vz4XeJH7RtELeChuvO9tvaraFF1NudNHe7IJK0hoFYn46T
UgrXywOb9haupzC8RmjDxDq6Ex3h+FEuFQ58LWRBP4HWWIbdftjbKLJIDXww0KRv
1VN41e9PnYBj15OinuTUd91PMuO9KM1XDm5qDdE4tVc8Mtm4ekRAXNvelbw3U0Ss
9HqJnLonpoWqfeeG0ngMwRQHddpZYhO4hXJT3Tm0YFuySGjreQzmxQJaNHHnvBse
yoJRY0YbRDFqLYJ0gDBNFVFl5Vo3RzBVaoQueBJZSbanvjkY5goIacV68x+aASUS
0fFfPc5iMIHFyQnTn+ZxWaF9ggHWlvgW41s5xKRF6+9ixTsxtspo1HXAjZSiZlyl
Ol71po4lwg1yKr6J6uLIqBTZSj0biRQUy1FWTzOs/tY3jIpy6k6pvIgNf4hRWrW7
Tt+WsuCc/Tf8OuyJztNtsGIYpzFqGyvws5VBmA5BCIJTnis0/wL6SMaWloMj0Cuj
gqJ7yzdOmLrnt8DxrBsJV57J9zMpDM525uAhvMXDGptrCOw/eBE6OYYrK1JLyiAM
Mjx8jyWVYGh8esnyXNmd+dAxNH1wbgy4Gx7FGwIbsNmSpa9LGPw5JyO0xxNzLMUz
dbE3e8ThVV0eS5AKZUyzCkDRJyjYM9ddSiXB9scBTwQQ48pGEJtj7h2jUCe0xy0X
PN9/RKdUyhFJZySKoKxRBPI5sHOPedlvOmHdIGXyRegh38S7+UQg8AIev6QQ+kAU
pO6XsTaxx5axnxa436JUhg7Zs7CG1k95A24n2/PBeb9fs8Kcnmy8YJm1Nlaz8LzJ
r5SOVMLbUh1oXRMPR+tilWsDr/GpkQ5QrMhBsCqGjV3ubOHIXn5Tv2MaeRWtlW4v
ubOFVhbHXC9KNDKDJsXmo+ypz0+b7CDHuy+sfmNFo47vDMhQBZ7sv0sPQWT2avbp
md2D0CjVloOqtI/HUVqL8pO2t3F11nzVol6S1PO1I61r6glgUYC2+0+6ra+J7h/S
hmWG/dqiNjWzBCA15JpbnsEgl0ljE7PZRYuc5OV6CHpUHhrLYnpXk/UJMTMwfpF9
i1QAkCqydyc1GSOpMcoD/L0iEqZ+XCyuVqJ2o9nQ6ZrDnJOuBFNYnyUln/JV/ate
qEtBknpYm17gycW0AU00CTRkHvMXZkrTuikqvdjy/kEuV5yydx09TZRhOqvER2I8
ltsO/CQSmdXK1tNsJGRKWUInBUQfyYo6xx1QHWXmCNoE/iDYlI9YOPin5BABXd+W
ljgqT8ru8GuFnlsMhNT4vcSMCVztu1YGPlZDOlsykSBF+EwjpCerk162EnQ0tv/H
QKIGfATztUO9HXw70JRm361iErs7yNa58cTCefNLwOiOv22TuFs6QrPTnB8o7jPC
KPVUFQk5CsJxMbTjiQ3g6DUz7DbiiQeXSdtsKBzzhlVpAOPjUWLm1AxB9sjRDLdM
nxWK7dAlLEqSee+2e0JOsYsQL1eGB+SYo5wjtiyqPWsHJdESg7CXSp2iuIL+TqXk
AKlFMbipWFdlWYowdSG5JZYF7NpjWRZ/sHiKHRczKKUodgbFVFLaNTOcAQpoZOio
ut8J76WuJtRrBLN6N0xNIhu5fQcKAdIbjvsWJYmHWYgkEuxC/GNRujbtFVl/BEN9
n8fSSPbn7z0u6eeZj6svNJojLoGOk7+ZeItNVVGq+f69vEAqhWbLiJRthNQuoPu1
Q0WOVDJeIYJ4hODOhDgfHlmzB/MIT4sVccpYgrgG9RnDvgLAfSvs8h+0XI4Uz7/s
BYYsI3RdIXC1Oh5hf8TUcdQrawXSysxEKJXnb3B7d9Cj9YVBxFXWi9ipfVM+1YeP
MvX4W5U0antwiBsvpEDYQ4LATMo4/Z+DLLO+LBF05y1XVksETIBiv7l+Tpel3lZb
dOQGF91/sCprjwvtBCDUxL+//q1Vx+UV3FuKjciKwuApYisZDn0KWDQWQ+dfC0zF
MfoxUe3nr5akPBBXo0P6QSdY0G9GRgs1VF11ZePdXHApCBtoumK0RAgYpdRhQQLS
foDCse1xsN+nvon/8I/3NFec+nAL/bRk7AAFVCDuHu1kFFILL2s58YBygIyqp/e4
XkFShhZgZKchOtCnFjCXpzvzCyw4tlxJXwGK9OneHDW5rZJ8YGoGM80AZ0pzx4MF
qCu9HADWDzmFvkj5Lfc7u3iiZUtcxkEaSxfsI4z8dmGGoZZVZrDc3YExIB1N591N
z+PsogYjcl5bd5Worda2d8afnpYT4No3DvchQrJlSRKTK9B+69FIVPzcIMLnxj2i
oE0Gqso0CeC1B0Pul1fqi8zCAnz1I5krhNqZNW7VUTZ3elW7Gs7RcemRyN7qXD3n
Ni/8znh33tMMPEduXt94UPZzUiRcULO/m8js9cb6t0O0iVMvo1GwyYxiNp1LT2Yo
H47DJAgqUeSh18yFX87W7bizasDW96z3hxGQYVn2342s9N6ukizZGaHsBRsDLTey
zovwvuQO+up/QMPXTUBRtnwfISDGtRCH1KAm76CGLiLUNPJ9dbZYptUtAjabAaUf
cJLIeTGrkGnr3KO26gRdMIlAOoSPFpCgu6Whk4diLVTs1QtxhZti3aefatZRMQwD
wk/K24+fM6/eWjG2OBPmtR0nEaqZfvFyU5l3WxIY5vgY0DNEQgOxki1nDEOf6NbO
HRbONTFHqy4ZGCLiy7hqU/qiJWlx64yTwqihiY4VMiiSs/9QyxBaBWjTfPjpOiyw
d0Eg/i+jzmVwOh9dxLOFuxKfPMXdyG2C7fpj1EHmmIuRyUmEN/327AkEw4zti/8z
R1+6Ch0O4nFO0kPc1rUeXnAnQRUDQgmxugOQKZv4dtfzfR1091L7PvDBdRDJRHHg
hx58iQGrZvDjemW7RseXn6vjPjHCpctRd3VYPNwLNu3k6fY6eVUfdIQYP88kifvf
SVB9PAaQ2lK1xYYlGazQkFBDeFkzvD4+83z2ikgPnDleGk/Sbv7ncVqNgXtEj0vH
0gdIzZpcU8cZN/AQ7TLrgkNEZuv3kJQ1M6QmIIio/GLE2eR0ypmUZ5Mv4KMPqZoo
1cA50kowqmJ598w907b54iu5XFEf1a+l5QPdlGcsUHbI5H5sWTxJNCh9BvFfQzqi
xZpUwFGWvoBpKyPWfTPzF1ZqKeyzoXRU/uZ7mFcuw5SmZWkPUvwI+XtMrx40HZdw
/nzFwvgsAG4n9t/EKCD0CKcsuofRF8m6DAXz7K4J+/9/J5fcv3DKz3xdUFWwQ7pe
mIzgno7WXIK4S1BiOhen1kzy/Ptx362eiI5uB5NxKrhVaYG229Fz3oOp3js6F5LT
SZ/S7W9y/jFRDqkFgKbCkJt2xaU/QAn89s2gFm0mIBJPCwAJNkfQDqmVXOP20fgH
0KjI51Xl2FTLvXDbw0W+eBOyG0Lid6geENlSbq6IMWoZTs1XrJX9bbFttvckrHOi
aInshW5MgbqJvRMRIYrFFbC2ZFiKhV1FituwRuittBjgoYuFKTdIvuwY3dIkC601
k23U265R3naWZO/wRUe+NvD7ylXN64Ips89az1MlXfs5yOKNKbyDxUmBPWApBiER
k2xAqO/VA7Wx+an0eJ8lFq3frLiDARM4hGXCtIgD9GnLBfa52OkGwx23AA27Nc71
Ptix03XtB1ppx4WrbbQFoZz9fOCHD0aFRX+itWSmfgsOg3D3aFWVO0V2CuUA21a4
bChmWUyW2fBmTG+8XIl22mxCzB/P4lSUTQZJIHHRURAgqndAVmMdKu8xXNgObrcg
8xPz6gcOnCdbk1Ybg6Pi8DROa+nxO2wWq6LFJbKEw3hmVafrQ36V0SkUQAT0hymy
jfkvRvijuKHAtKuOG0DsDGLfszLsNkOUd5JMSgJGM9VihS14cRVr7KNgUGQboG8i
8x7cQ2fn49iM62iaOK1uIsnnnGsrr00Z8dPK8XRwYptxVFj+zDVSVpZSh2MiNYg5
tIcleSZF0VKN/VYEhm92bGQKbsh9yQD4VxpUR2y7cuAwspItW50vCuBZfTqlVk1J
MdR7bD3/ft1U7gJwRAnOwl6q54NJAhW9MUJGEOjORLAChwRDyD2d7C7/Gvk8KWyH
QbNuteyX7TdquIsliayGGM9ZifePVJpLKPmcLJwo3K9+mmx0LJ9PM/EXwMk+/rsz
lho3cM6O+edSlqbf+Wq23otLuIWV2Ny0uwtWDdAeIFavZNctRvRKxWoEdLMKqojh
woBYd9CJfS8CXxT82HemY8Cb7oagq0wDT90qtf/QQux6kGAyejTVMOLLT4XTmOwH
KoIUN6YwGB/HEnf8ldfJUAA5F5HAuNh9mQ87/965fLuFlJ0DjyAw75Xnf7e0STnK
Z1bZDLBq5rvnhPW8hWfW/Am6G2Mzpr/bfRBmRmOdswMTus7gO32KsNK4LzEsTgKP
D7bmeBCm9t6w55w7cGf6nba1LC+TAB9kw9mEJXggS5j2PG6rXUMp9ySK2nZEl+Kq
hVyra/LMvVG7L6M7CWuPBMD0Ldc69/QP8a8sV3JnDIkqzk52YRwExl1RINnd7cwo
SFJbqFZsai9M1aU9zlHJJRpRv98aPFpj6rXuk5gZmSvnrTp6VzrJWfd+GvmPVuRE
juQIrRgf5Wh0VcL6MLq9LiTYHkE7+5+rK3uAZTCaWc5SpGemny6ezqQKXQ5d0hOi
lIgTN68cGKRH9xUNktbAiofPi9TT2n4li03T0m0W9P1cdayeryNbJhGfAQsU4ygF
lfKTm4SN7HUbGRGJfrKX4+eJOb7943lRa0IgkPViMrD0b5L78HeU72Jl2cuq2yGF
6d1ZFmJOAFbGNdfznUEXdbkZdtiSuT7zgkSaPQxbisJQKYjYstv/cmlbqJlW2U9z
hBEfaj6oz7a5W0ZTBklyHSKGANGpj4KFJk47lqzrRlwL8SQzIkmu42m59nsRcXXN
uA27Vkj8D+WLgFq7P/KyqsvvgR8gwdnnwXNEQ6DJBh5AOlSa3mErQu/TPn/oL3yC
B/N1Vxv89v0keKne1pziGRqF/gO4F87nFiY+efepLXB2QdKGTUQHtbcJph/xbJRV
rqz7RvhU0Yoer7Ce+/YUtzoZOYlWc4sgmb3/6HuShoPzmU6KxmqjziG5gi5384Xn
XiK5OGPcmIFXowP+8eV9l6+/1aTiUyCM4OKR8+mFNX53Ld/BDFSjchJ5ioaKW+a1
Z68jmuHdAjv+xRDJXc0eILslR3G0oPKawWMIG4A4rFfxrz1Elo+f3CrGR3tsr0wX
/8kvqxR509S1t55DV+qyT4pge3AZ/Og/gbObKk4ytG/SK1YqasBmOyNDjQz4FvKJ
z29ykvQeqV90Li5pWpoARE2qYa0BuKaWjgOWsJHJ4J0tSdTLdkM82pK4kWqtJq5c
R7w0b6aYgcAJKPnK3CI9lWS6WVyFAC69j/uMapYXHMSvSxZ3jKy28ByW427ti4Am
/Aem3Pc77tX3DWCEUIJlY/TUJ7sagvwoaMA+NE2cMS8sGR5VsUn5Xak0hOL3/UPe
/rwkACHasjjm445o5wE6DVAKFDjk65bPqO7hR69SduzuaYWF6i3Aumzvp2WV6eNO
VSrVoBOsGIsB64SbvG43KkQq1CHcA52p05XEa1kiTIorvZeDJynNunbwh8EUWfCj
LakfjTpbcy2Y4XjZZIdEwzrdWDzQxvWWj037a8Dup5Fj2vSqg8H34g1sa/Nd4+x5
sD+NwfHseRnjlPuzCWNIp6pLzqfdw++zGlJp/DNTmRlQ+Wmvi2MAn/5Vow0S3Qz9
pUTvb/IjwxDtAgs6FqeJb4PNPgr0kU+oK/72pEmYGHK6VCfSIjxmIx3v6ZchTrRo
mOlGUinCQlUdvlem7ED28uNo3/vrKGZiZjljkF1A5g+S0wwt9YgEpONt1hs6GEJX
ADW1adU5NZ1Hk1VCrIsgjaLxhAOL4AUYX9ZQpWsP9ulUFAReX1OOj0s6SuVqVhtP
WtoMRn3G4nbxbsgCtTh1CqFUlD6e/qM+f1qUKSZ8AKh5mOU50iBfmjTJA8IpCm7j
YABKvTMBR7FjS2y9JKz4nzjAaOmrxxKOcdbT8LNTeH52NSqEOVozl0WylzfjTrKn
46sEXdHjZAK2pemJNDy5wcL514FoVRVDGOc+JD0Cm4PO30RUz9ynkLahvOXa5pIc
B3j7q/NEA99OjS721gZZfm3OTmHEUOT07p28j3XGTszfINMtzIX77Ju9dwa8wky0
lXHnknVyFH+s80MoUbvt+7253ex9o5FdnmCRDQAnyCT/eKL9ffZLdzHEsEUWyBa3
QdyzamtNP1BGgIKlL0yOMhyKsxnbgqp/NpTdYoTP2K6k92ASOMs6t4ytFA9kdd5/
spJHPrB2Lmjpa6egoOjaSIQkIhxM5+ZknTiHrhJB8MkvYx2gPbU3dF4xEKe7b2B/
tquM4dMGOfe7EZlyBq9ZUR1S7N8uLjH4z06PfOZ2riI/jvzOyYmgYG78aF/mzyF8
UJeQyoFJTxT079vkY7BidDa7jYjKjHwBQcAtzSTCrAcXE2HSw8xu8EN2NVVdTFmM
EluvqEcWrvhFs9rFOifhlpB23pCY1kg7OXiea5EI7PDEX/Wf5ybJiT5aSwCxr3q0
tnb4DLPnwpql73CKAqlE/tpUd9dV3jDOIXv6G4bD6setEpzoB9egYPCz5k9/KlK+
7XkKp5y5pM2DlhnckMc/WOUC/PcQXVsPwPf67EX7CXjMhUBOFSN0LaYhNS3BK0RQ
H9dE/dgaS9Z29pdDs+9roUtVUpdBRnw4dpoYt+/pbPRjSMJFMrwWdeHnnXfCfmIt
34wtRX/ozb23eT4b+XfVZXy21INADDjXx1+lfjr1Vo8Gh5Fp/UU41hBSfFAQ4SSd
8P7fjtAPH4nrHcjYHsWpcqxT5zadFeto/oTJ4AncrGzojKYdGe7FClzmrTuL/NlI
WmGkVve/ONmnEts7YprY/F800rnu0wA3aqNSThJ3YxWqPDVAGhGJ19xtyqFyjhMz
Zg1ajHFPPgqxOssN7uLhRUH0WDoiLZKCpFGydsDtBfqAGh4Xr3jsONw5IAlVrD5b
WpKuFtbEx/oS62+x/h1wNRQ/FruKx5oynEZ7KbdZMRA2ZnLtnsyiiyNcY6fZkXRp
Avv2lCVh8UJDi56RbHy6/Vpn/BIJgokgOpKCo1ApvmZbNK6H7rSAma3g925seHA7
46Gw2dhPDifLXkfkIwQoOOcdp0RqSlGdii9KLZAVjq0thOAlt9LHxCn13GuRjD0t
tniWHpTjGe9juQcjpXG4MHDUyuvVjTASKM4o2B6pUV7Kie+zLhN9IPZ8FsYXdJuT
YsAQIjTUytnopttd8W8f4+/X9nFxlKJYna76ocPJrypt28Dbjgnk9cSEphqDdIF1
Q/8Q/9/ptxpF6GhBHYHc8LaqR9H1VAnWzoLxux4rE8udAuMo6pNQp8wBdaXhkt+X
16yHzmTKseMjl6MNH6NK6o9HISmjmV6cPOyhDk9n/RqIOw6k2KL5uQidqfEyYM5I
u/uHpv5in9tTrFE2EhXjeIPs5l6DU+zb0QpFjwRMbXmnpfM1G0mNL4OGVGrY/Att
LK/9eXr8/pQjZ6fGfibX0itZF4By0FrOmovgSEjVHM8GsVXxAMS9ExWR5Y8SUfEn
jI64rzheoIR+gIWwmGRavvGFynehShh/CQli285xCPujPTdU/1b1+DPJmQ8Bn40P
MfqlxZopeKsqrBnwb+k99kHDCxrq/WJNofDchAf/8y9QcQNtdc2l59Cd09L2SFx/
ZRqycSDW8pX6SLA/KRYpWyugI84SpNzCMKCpLuUNgW8Pid1oCMVF1R16x/q6N/Oe
zkzZb+6rft1G09F9ykwAMwSbpaG+LGQVsBL4rfWbH1SXakszX3Ok0o7sdctjJJIK
9q6ffKmEioJFogIKG5mYUdCnqEOP679kc/F+lT4TW/4096epT+NN0fJsRsXlJzPP
Uabs2H6CvQxD26jJCqY3lQC8ftbZvt/09DS5nC6/WGN1rQoQlzaTvEjsYi/+yXyW
ic56XKpLFCWLPlF6ySc8PARX2F5hc7rs1gOSQIEFX2y5cqB9g2HExQtsBC4LTwTq
fKt92gs+rgnjKAgfjTVH7U+Tsu7P4+8SD28u+01JkRu5Rb2T7tI0PeKOgylnDN8d
LGoyDWrJfkAclIGHhNKcDmEAyke3FOIhDOKc3hVj5V19gVNTiwAJXcn8bGnUw61U
qzx0x1IHoRBrJm0+1h55hS/BekZAM+hEGpvNJ02eS90DvWJIRQ2+I8xEiIM+LYNt
Dk5GzNBTZTx480LTjzMi+6chze61TsXnH/5po4xGxutOPlJsskiX6vbzf28mtNci
z0PQ64tRCg8VVC2eyqV2stERjb6iQEWdM6AEGMPmJFvBfdWZH8vlAkLCp1mmUDLx
AZut2nKxIUgGiYsI4dOI4jQLGfHDrIZLcGOkgYYmh6we6pXuLunvegTco6LVTj0q
eYsutNO8ZCridQtMGPPACT0yBnQKyz1ztSKBdf7mpAUbPadd7I/OTRL/U+VHYvut
1BjsmoAsHSw92s836SHMODMwX60p6VF9ojjbVKXbjGa+qTtIiCZ+dkBboW9bvC0g
VBYNTTTvHYNrqU6UJdzZpUMt9zn9ZbtxvIgO/+xeymRzBJ6FMMSKu1/V22xNMjhb
gY1JIVuGN6u72rTsERLJltOtPYO/1uAlkDEVYKMmcG+UDXNLwkdifgOxrwzTo0lz
hArO8f/JtZbXDha8ZVu9cDQyWjcQa0gDagJbktXuoHj4cgR+dtWRcm5aS9SpjlyB
D+2jVzp/ZlzGa0jI2rmc7TYxoJiv4gItydRoizBuwv9HVjNI3DCAQl2YtbxbLTtP
aOtXs9t7TshwbK2Z5KeP3ZewOZ795N3atX7RTFXrqnrDrlxLEEIK8uSmeFenj5jC
Wg3phK8GFCLaojk35IOg4qkGK5UzfLbBqBMVzANkhSYKHEeZtnQ4G4pfZslJj2Tp
rCLuMs6Bo2951RljfEMTjTzjnHhtDir1c8CkhHleTu5r1KR1AymB+FJpbVx3+pLi
H7C522hVmDPKtnvZ8F8G1KwaljFw4av9RluXYUJCyj10R1DmW7UBfCyJ2uw6c37D
7zRqCBZkW4+PRc0tb1ZPZpkNBSGQQXeQdwer5UywUfMZS2A1igSPxXXxFJiyy7LV
Md3W4ek2vKl9p6Xm2ovBGSaXyJnpixbUfiEg0hpu1/c/++8E2NT4nQKajLfGdMlw
h7Z2pJ3/lRzAdZAmXU9y7riKZpty4esmLtxVbZy8GB0nC4dj1NCnKyHI33fVqFua
ngZpOR4sna8xuisr7GZZJBJledC76udNvVhd/iu89VRqpzuIjkMJYcRvSFMJXUZH
WzA4rt4QFFGXV5V4n044KFJGonw2yA6tg+iX8GQVxXPxTLXa2WcS35g3QzgAe737
pV2EkJcct6QTu7FtZNxZckFAokZfvTmTrvdfT5LXU3MFvcry77qvkH5tElF4uUjx
hdGW8waewAb+OIWhgpuey3zPY+RjGdKa9jwGd1rGF1DAaBRJ6Wabs7RTNO/zkXBS
y4l2h0Ih5qtY23/UC/V2kSw/Cz0xiwcD7jFF44gYi0/V+YZYckSum/gL5enOBJNU
r28HI3giVuEmI+irQz3uuX8z8WSGCp5enINKT/nkXbu7TO1laEWPrwUs/gU1dJNj
0FW5nIA0TKg7Kax7bnnVs4SqM+vQnoXiEvdeZeVg/Zsx0scUOGgVzVT/yssxiUL4
XMSEEsmy0anybVP6K4jc4YBu5AHvL7Ck2MwEfu8KmCrrR6wDz7Fjy7pVVaJWmTXC
Hf9+EF5qFYoS1Gp417CGTkFbve1kJ5v+WzUvJruBKJ4Zh3zGDnjkNn3CjsVkryxQ
oTfwALO2Iq+pdZxLqBF67EBVXroa7zP3LmdspClnr6EFal61OLdDekPJJNZ2XqB6
WO5hpz2M/Yd2z3ETCoq7vMpUlCnGZXZVyI+QJ08suqwEHkYCc5NQTEBnrvRJobxY
WsW0S7t/uyswA+SxhEf+OPvdno2aRDkJ4OgP8PTOFuUTGyqq7eD3C/FBjwfOT6Gm
e067IKWONR5hordgtWmo08XrozEBx/SfrdgswqjOdIUSoFT+WM/k4ZpLUBw3T423
UP7DfDcaSIJnRZQ41Rs5O8M0ca4V5npm+AKrlhy4FWVcieN84/MiEPXKLCNVP9Nv
ms7MCsCEuWwBTAVfXMPqSP0cdtWE0iU56vv5g9fh5l8F4kKqI0/2E9M/8MFbMWY3
ZiTdov78x/sG9EOvq/M/gRN0L8pM86Dfv/swt3Vi52dhKe/HOOqg5ZNNTPpvMV8c
WAW4ithA70A/RnIHJxty5pQ+JCZEBNzEpsdK93I+xY96pdwh3qVO8F3UVxsqg1qu
WSOMyPNTTFltU6I6ppJeY7GrCkA0TWsJ4xM997B/kMWZdv01tDihrXdO/2Gic6xO
dz1fiUP74yaEAjgqChBhWrw0+p2tvwlVvdVQBYOMWdjFi7iK/6O9Aoj8JgNJXCfC
UOy3ZsgHbbCVTA4PU6Mzu+iNw0LJBD7KnTLrR6HAdF+jny5g0vWRS7+rUt6Nqm02
MknIGpvpPF6B+3VgjTsvDtAYbNKGiuNE+KQi6XRXQ7yxApzNeo95gxZXqR5+ioiN
LxVuLRXN6OnWJoJLvEMuZAkk9bWT4oOQZX8GhsGaiz7PTKFag9bgNfIc0xqHCY1r
6S3h3E5JJQXqmoQc4Pa4LdqmC0LaegkllMAnafQqbkt2fz+BVm5zSX3N5FWCHxh1
OGkHnET+8Zvh2HbpNtn2M+ONRr9pKXy9jefwCt0Vawts1P1Ez5DQ8W6kWB1nyqzM
CHSxknRA27TjhMwgfGkbtJHUscVxSN6qbeVe3ffRvKwakU+awkbN6tKE/X4XnCnV
eiev/BQz3VMK4n+PGO3JuAVsdRHXh/lQLq1+7JCstYUgiAd/IK0FWkpOe+3BU7oX
ufs+ZtEoBQ5OQNq1+A8HARECD/kpNFDW4IrRpVDSzW7wTJtLef8f7iXJK77ZLZo0
ye+jNJbYG2Xs3DoEcrvgdRVjycl01rxDjYapii9Q7vuHl/qvYHmrFTTeaNKsJRWd
mYgmfGBokjw0mR6HdsTIGtnzggx+Mr9G9fswBHWW1kAy1YEiZdJBHsaIlEVBk7N4
UbBeX7OnKn1c8cZt1zydMgviYMPgGrFdrAwL6zjB8BxV9XyS4smAvBGTeADn0Fm/
NySnnYHiy6uGihfjnPyOyQPB3Y9LWC9tgrmYJVfY5PNukgvDt3w2bX+SkEW02WNO
RHdzOikomSsNT+mhSOw4QO9IvififOxAgilRqFxUN1PXSyHwOdI+uVlxYyQtMvIN
0pgVnuoDKR5ybebIaQRjFkIfrSIzYlcJ0yvwlIEBlWCpeU/Gl4cIuIp2TjX5dRF0
zBgl+QYWd/+u+DHdBW44242ZglO6RlaJLXnZbBiRBr4qFbCl209VBrP5W01IH9hv
V9Ms+5HO29L33POmI1+QNeBCkx55FwsOwRz2KjqaenqKPlxb35ZuGwohYDihgTeQ
lGcEC8XD3ciMv09/vY1QR9AQlvDvMrM4wYLrLh4iVyvSEinI7TBFOZpTkNmtZ25k
fbAK3d4hrKDJww2sZSZwhpz9JXqS0+r15cX4zJRLkACUSSZFJcLCx1de2vw+wZKV
D5JlRNrrNZJ1SNrskckwfqlPbP2yEroXcIrrNADrAhg44ArEOOteqm1EMH2gjEvb
F9cmLhDmW7lVO9rOxoRn2B/jtPg81wN5EjiVWA0GY2sW+DlUVsFwQe5vxOHIuHuE
dusZxh9SZsx8MP4x5XlGO+bgU3UOtxbFN+hCNCihnlhxb5Pq9bWcPMJ4gqcbb8Af
FTWHcSzH5agJE+7Hc1cJa69MPbT993FdwYjMJVD8yyCCm15g4vi48GVfE3Z2V/Ms
8gt2uBHiVymvpTa+NVsrPCZUfXrMbSx5BJsPMDiQp3PilDN2xcPt8jJMbhcZWt3/
ZIsr//i89DbGGGYzVbY9ggaqM1aSDRlc500qXJNBK2j7Bt/e49wQtlL4w8O0dA+n
G0s+XKvAPwqWPxY0krTnvp3/hHawzD3745K8wnOP4f41KJDQlEfex4kN7Brv+lHn
Lu622nNUpc0/4wHPAFRbt4jcBifkOsEyPiHpqI6i/GYJH/OAW6EHEvQlL3/T8W/L
okUOEGCe7jf7SQEbI/EpW1FkKWHx8rMI/Wm1SQbN/uQjJ28DHegp1x5D9zyjEdwf
DShrpD2qYD3eKqBpvjlmznKH7MAa7oTBlUZzmOSOqUvvu4oQRXF+9JlE1z9GSJZO
7qXMxAx3rqpXoaG0fcmDDHRwk7Inf9BTPOSjf/Y7VMYT2tBEjNX+qb1PRxKgZ7aH
wXWWsxjx/9tevaLo1zM+jY4AHFRXW7xax+1A3FxVsalsCf0XivzLnS9bZk2LLMjr
822nK0Hbt6r+Xh4u8+/Y3ByQGSlQ1qNYrXmX6qp3h0qLTbk95aidscWHxXj318MF
MzAV+5urcu/w10FSQseXLkALM2tj90P+nr0Anebgui1gkIgF3I7zkHUTgTC+Yh3n
mPXuoM0bE0XqIBrdUGYJ4Z7LNbXyf3aN+3gvnGh6N8xzVl724X3gZCl77r/c4eYl
DHKwHZL+19Rfyf20NWWFrfT6f8HtNlqcIwPvV0dLirwcYHBz3B8pgYv7eXek4FUY
lSsIZR5aIOY+4Xw+Jgjge6kE3x5Ysd4/nKbMd5iEqzctoxwX0zaUnsFjYXPxkhx0
7Plz4xF0vcrX4hzGMSs6fBJp0I0IBsKQMsW9mOekij/zxUUFVMso3SO88eIV9VFq
J86JDFyM1FhlgWgpzVwyVSDJrKfQDIM865C2pCMY88NefH2tSR6NcQvHE2OC4ex2
1k0FwY4AZrPWl6B76GAUispJMWroVaTx5OOMAkGM11eZ/QsNlMpp4EF2aFKuNJXA
SkrFetJfgBFby2XYO9x6TYdQ5J8jHTOF/Bbe3S4Dr7c3wjvZRA71S1lCHLt1M1SO
WuBJov08pll3Z+bHzyoXRqFc6zT950t76hmdw0XqAjwr4ouhBfo35fZBWGXQYFkS
tloCU8ZYMGQmYIpil++M3xpQA5LlXar1KLp6I25Em1UQUuXVT+mwf0i+DR9r8y6J
kuo8xE8tBQopx1FmA0XQhj483ZOqrBZMRNm5ApYO921Qc29b73pRAY1bMWCsJkRf
KvNG3eVYCGYkw3lumec+gNYJMzjiEICRCCO3t1R5mDUJT8HMebCcnCl7JIyh5mt2
uEBKmefbZoWIRwjr+dG4PQc7olzK28QsgYbGDMGyE3sY0Vv6CJuychUymOV5o4+P
vHpO83EqI6lfjf7IrnTM/NeT+Y/5kgmIBAzWZoBjbqNJBR+jQS02aqucBAubEkE6
G3dK1eEl2sVuTZz+2FuCMbSuAUrVe+cYNk6OSvi7RC1y7Vw4Yc+w6upiz7HryHUr
tcRdvAXFE4crDB4NphVday5GR0I60kGhyWBp2O9aGOEpTFypfYvSqXAhczjUowjq
dPj92gGnsaof+G6HqKYG7uec9JgVhaULme+pqcoJRvbgghKMLlACDl4uFyPZE8R1
TqAPgflqP9IpEW1RlUDsEWTDkUh+8LJio2vL+b+zC2hET9sVJ2Qx17r04OJqpkLI
jYSw6NJMTWzMh/f2ma4TjzhrTZXkJ0OA9iqBGHvaOoiZT18XdWQYEkP2pp/+TunG
MmRI3jMHOdQr6j9dzgk5p0G6mrbfqVlHx60oQhABUi3CxTZARatO33sKeSWkfCw1
l3wq0MDGceIVPz1D/XLWwuRYOHL8oXAs06zz1oA2TfMmpHNz2eT31woZfyNmD6qV
qQX1hhI8qw4XCEz/JgTFizEFLeVaaBY6uEILxQ5uVzNusuQcbFwopThBEL1qSWBj
l4jmgm5IptdHcbAhBept2apvWdS7Wvl+TyN3oi+viaL17K1AISODo8sjWsjbtMmV
MyvMHvuosJhzI+bi1Zk2PtsW6uQSrnxh2Fj/vo0S2mPyGVaguiK6ooVe4JU1XYcQ
Pti+e7w/2EHz4sfY/IBEfzITVvouEyDkc60hfK0WoJZKe5NEwrmcHacCkuWd5EkS
vAEnEKicMRbjM2rkFM6wbeBoIKIbSx6JNm2PpMXUC1er6hc9g7CKp7vSfUipYA/h
aNYOKy4EbdyJuQ+B3p8sn06mBVptBUtdhP1rF5WoxF3nXqr9ypJOtU8MCtzJJX/l
hnuHCKOjZtYTnDj26L4JViFIfE+PFlowOMacngUDsqIL7dsuEmy2tPBYVRr+AmWq
3BF0TPw7jsMGxOEnSkpfVNueQUdGFENXD+PMXMyJXK/Oxwa8+z9Wc9X/Le5B5jao
N1z4AcNhsS+7lHPTPLnwB91J4XqDXc+0yla2Rw60dbasLU7AP/iYM/s+0gDhIStV
LVnWXHjuai9BOv2aqUssQlM/OpQ9cxHKCS30WYgL4v0/VaoAQN0J0kxIor0RUCV9
cdjK8X0Eu8xeQzUufAqYebJ54MZK++MqYOsYEFMBKIRLqrYopS8IdYnNaG5uRTio
FBX3eHW3TrrBBRVF+dBzhyreqVZRIHfDc454v0gpIPaKZnRXpEvffDulz4wvVH2c
RKgjlJ9JXy57ECbpiHWqnqWHuAN5k8LoM8Grcdjq23syXWpWPRzlZMExQ2a8LuHC
oUPygvN2CJm2dY6+jN5GhfF2zuf29YlpZbHpNxK2O1FgHh8xR0chkAnSNBfzS0B5
0ARGxW8hBoKtKqpAqiKU3MBM5Rqvykj+OObJbyWjseYhfAwCsBekUTSZn0eRlDSO
1ipD2DLlFxrXJsVmM31kgMIy/PX5hjN5gSBvZCJ7GBdxhigrNJSOEo86gs0lKmHA
GAOX+uSCn9BemKCE2qsl5TXvsPyFIGLW804zZYUfjz89vE5AVhxbpt4dXvOIm6bd
4+kAyvUouQEPeWhszns6cVf7Zc8kdZcSVdBOTHoDDK/v69nKaj+8/uYmC7SA/Q+j
U7hG8LqZSTL+JMp6umiul8GtB3M2pN2y0t1rfd3rfxjHCwCPodSCdV+YkC9+Kzy9
PlkWsJeLDYEHj0IT0cZAvLmWfwklLgoWB/+Z6WYfb/iIlrFXveaOtmR+AvXdeQ9G
cdwVk81rRXhfb2WakopiaJuA7oTwKOvggFRSKz9WdhdDx59jkQfXfJgCiKS1Fdbg
CmJA7uCY/lRGd73zP/Lhl+Orb2VfbAi9SF6ch+17xdBFUyzdN9KyV8T1ycGGsrli
VxqwAggc+6S4uTPPCeNgkPTfYyq7D+FVsVfvmPrGrvBrPmp/0t7AISduX0Kh17s1
yY5sRshyfDPx7witV1afUPDN2jl/aLeRVsYn+JOrO/zUnv7Sz5HYGL6u4EgCKVDe
pFSlB0zpWRIfNtIM9AHDI981MDBhvmXqz/X4KINytOhul02D2wKS0lrqjkTapubf
vlZevYzeJ8HtSq9flWyfHzjDbNcwZH2F3JSlIdGW6MwzwO4mdIXsc0N/Gr593Oal
gD++E4/BU+aRQT8DbD8+aceUumkiwev9n9tWzdqhGRNgcH6W2DvXiZ/a8nlePfU+
2KO7S1D4M5DpXa2xUs4RMDqGRKTpQpKzDUezruaJzVOmqsKsq4bdkfo0ANaq/9KE
UUgGszLTY3MXPMrj9XglZeWvu0OqD2jeMMQtdIh5H9MdHJLBodoBPTo/oQm36ZI+
skuplWjGw+qS9TQh3t/u5WJLuAa/BoaZwr6SH0mAoIko1BSUBU7RmLiczP1elz3j
9kMg356j2687xMTC5HwWIO0R6v1nVxT+i9liPkmKdSQslyJCMgJOdBLYFp3ItDVj
iCRH2u5bune5UNI9dV49ncNWS1xm/zCqkF/ktMpptxF2jJcCKRKBWXBlCZ1wW3TR
EHwuyDrUzSVpSqeVtYhoxkBVTAY10VJ4/2TH4gqCcB0tU3gMfhShAkQmi5ojHs8R
snZyyyy5xqHYg+7JTN0xMhaw7qz10imjdv0WPylcx9U+M5oNNLE14TjIrxl937sh
FHov8WhYkddumPjZcjE+E67owEoGmvmYw9RsNeyh/3LCHhAHVpmKw+wqeCPRmH+X
sL4dRpGs3TcLfIVg57KE36CpiYS2rK4ExYTWjuPNZ7j4kIQEeR9AdPms9kYpi5YN
S+/XtWjHHmIupEfBBpGM4ylS6biJ8GE8XHiCftXpYnQR6CuybbfwB1vB0XoutHAR
gqthjyNcMdi+fuaCj6AGpFc3K7lY2WS+NJceN+KrIpawIr5m0Qh7nRpyPDjfWEdy
ygDT/w9S6EdzIBc+54QphzSrkKZriNjLCldSX1rW++o0rMbAq4Bygodn1N1xd60f
sqWyxlVkRI9IBLWN9glZmXeMjBe4A3gMGENkG+CzW3aQDyFly4muMqRYu2ru6Xvk
QdG8+ku6JaBvWq92R83woY1ysGAPeKt4INlYaGQ4QLYDh8aSGawbFgbgXXtexoIm
lC8rMsM1PRfPIoNZY0+dF8byJIXayiYJLFLA4x9XIL23MIVXQEUQMuyK2NrtLKUY
iCksn7vXIE8B7tnoTPeuMXLj+sugPlQN6aSM4hF/K+Z+4uWjmiSbohYmWQOH9Am+
aS/jEbZU6WlW7ofzMu/xAEzikcZDZTY+9gpYA7VUGV04Gg8qSw3D0IZ25uWDryDX
8CXHG7Z2zb1GIXd9zZseEipiExv6abelTSZFTkyEHVBlI8TBNlaUFaum/bvAuMht
tu0Lo55LWwXF1yRHtBjC4IGGMwJ624xDBycHPYXB0JDSUyQPk+l8b9KVl7oV0afi
08KazsZQHw0NL10ub9gWWxIkoBoqaNq+Ltyr3z9zQeokqR51aSHiTAflVZDeuezH
97HjEUuLABl3u2x9vRsHCVEHz9fE23Hd/pHvLf1gFewPh2fm8TiSf/cXUxarrgwg
LTnC0s6iHKAtlcfPWJH2vtvSnCgb/c/Q014quW1EXtcbV13LFAIEQRGZp5cVuVyI
EyCOaG08Z1ZtW4m2MHIg0jm8pU8eMNmHGfh1Vr0VXkUtqX9f7D2rsaS52d5Gw0wu
e+VUKlmrqo9KmgNG4oBcyTSaJTdctO8kBVKhBY2sjYhiMcb/NDhI1BXcVCRgucMn
bkjJmSuR81ZUf84+IzGJmUKyYCb1G0NkFk5kMH6mMnqTfMyBraQDlerNHBS5mvKD
Tb0nZzgB3Vh7UsvVlRoXoqQcZkr1K/ADoR3sPn97l1lSx9Zz8R0GkPuzHHKms71p
crMT968vf2KJr9A6m/GAfQKEjBK+0jAm8IytIg9C+9mWJ0D8UyAcTQaDjPfohIZl
st2Iwg6iY8KhaNNg+iS/eVYS1FqE+7SPHYtZC91l/bnlmIrbiSm3OfGAvoMluYgv
0gztBFv6XK/NNc4Pw5g/4QHpMuDNUhTfDlpsOeIiMciMawABqsYB7n9atKJvyH+s
zpA+HY8p2oED46+MWCB9bGE7cDZ4GXU2F7Dtj7KeGot7upNCNyd8mVMP/dCFkeB1
MlVM58Wk0rWX8gTsK/j2+pvG/SHTQGAdRJYo2Q87D0jVJUEdgso34FqIigwARirV
iLmcTzK/7+bo3BRfFTgeRPxzMf+C+but1w6olwgFzhKGONHOWCh5QGIKR4wVt0FV
u9ng+Z4PnBj0f8Bw8GVcRQLRimjemfw1hk6CO+TAoon2cVc657Wtdmdb39hOAjOd
zFk/IgENtVop6X/1FWKaqQF64ymbho1CI2G6f7eStdSyfDTP9AKweblop77a3wtA
qRFk4N+b5Dgo7Wwty7MOgtHb9z0bW6ynVeQ/8aVw+/2PNlX85HpXGTRUF1W5bLO+
VM03ytDOg1K99vcyok6gOEc26825qps4AOYAtbHMuUIFwsoR/XNZHNI2F06a1Wu/
O9jsmh/KfiGrti0ucgAQBuQZKpwJGjEKyZ+6dhTLZ8boKC+mkAtQggXObVZN2zDk
6SOd/0Gze3RWP5LYM+O3vb43cqBRkiYih/Wtpf6rRN5iEErXOCBZq9+CbqaSMnnH
KHo1/4nKjG+LwU7I7LYv0JVrS85+91jHZ8Sypa0WjdsGMjNoBBhLHqJtO/NjFdne
v7+8yWI+ymR5J1FGFERl/W6/KrimA5qdhWjnNFsQGY6ZFDP2ck2IsASWGOVZjRCs
29I+V1rGfCqyVNgAsAE7isBIRLhX+B8+l1e8zpezKRIySGokirvzI0SZdCyiQexW
KM/fdMVfBtjIdTWBiyD/AgFLP9aiTCSWvAhjG300/aL5obT2/raCt3xA8C+CYkr2
rWlpx+T8mSApkG2gkG1Z6GaUi6WTXsAOukDiVGQCPxVj45Me/8x4jyzJode1o313
HtfUPM+HwX1emJlF4RnfYrrXVEEDB82x36mXFy2LozgoEghyxhWWF8g4iNfeZ46Z
PLCSGb0vLCMVSxSmaJpmmC+FhuuxWN7kE5tYC2pwvHZFkmF6akeCJGh2288omfh+
UoepJWMJBpEJacCv3wjoczzoOFlq/a8q0S+MaJ7Qie3dyO5dimC47/zVfQe8AaAi
ElegqEQeHZEvI/auEIzXOMxwMMHs/UUYUor1Z5Up/4jwLvDsybTXggJJDPgcEloo
xHe8egc6SBcDMSye7tYxFjWgGcdM1J4473PXkFKiGk2kE/iutsnBO2rcILp7BF0C
ACTIk1kQhXpMFykwGYClrEkZ5Tam38asdObaqzJq2kvz6NTwIcAz6/lDeq2s6cx8
yYEbjdf/eH+rRD6xqF0cCL37hcBq/m9HRT02qX6eut7Ka228qMR/hue/tDoSosed
ceIkcmbvEyMFH8rL5M9alTxdu8X493ooqldUs1NKpIyEMltCRjOf0G1GnwUddFQY
PKE4qbReasfbc4kYOqDMFeI2bc4oYrBB5yePv4oxSy5AWWGtbX05zgeUDuNiuUvJ
ayLLYupVXB+EGkCDYhty1kVlgBk1IBBvyu38TuVtS13l4dO8/PTUXojpBtwvlSM/
aR3ZCm7qZW4XX9B3Bkz7loe9Vi5OPInHqPMtSK7pr8PuiyF9HS4YtmXQ1bATy+6L
IaAOHupjsOD/vlZfcIpxhl5FGpuWCorDP2KHi8EAHFN9VAZT2F+jhv1FyLCKDZ6I
YZSiFH7iOgX6CbLDXOeTsVpj0kx3hzZMnMf/d5ot9cInyAY4/AtXjWGMsAte2g2S
RDmiM+bTZlmUDpP4Glmvs7Mi0Y7tMkFXrcFCtkDAcQ/EK2p7CyY1XzOQ4SB3yLyw
CWqky84VHtsJSfZRGH2743tJdbGJOb9Cq54Jm4iOwBY8Na72EQGsbV2Dxhu7oDAO
sEvHVo9v5VnD6RDGeJlBrB561s+9W6pe1tHnGngV8h5aGSz95QF01P7p+sr9UgeQ
52Fg8Ppzcd/P+yHaS4XMMmM577aR0DOBMG28Soq1RlWuLDCchbgmkOXcsLRDUICr
M1VpmSXlt1QJgmr0CmSPxVEFcS/4/ylL+790Q67I8XmPHyANrQhqzCnq6nEJwsOn
5VJIChMhJyYVXeyp5yc5iOHkRBRfIpGhfOqAoLICVO0DCD43JFtxkSZTUIfHxcwQ
2fps7VWSUoaBMMOSDOOWRAGJj4SzUAS/gmNFegOvmClSTlY4Ck06UOZjI63A4yho
V6dwUP86fs1Fh+dF0qAjQ/nit2K/2e+MZbSrOOgB+G7leU62nhn1bjNlln7uzw8/
JydabbFNzHUFHB6ANfP7ITFsXouSLn3XL+wvk7ozcp1vspbXm++1C7uhvqR4UP8E
+i9bRa3nlXGHP2lQp/9pc20g6xB5wofjG+4VzflSdO7DbJNblyAIJR75yAdjOw6t
JxothtklFkn6a/sHFFvH13r/BYQqQr+AI0uoqmW5SlmmfbBPkauUDFx3Y0efGPYg
flK4vsE7jLlebgHCj7AbnE8pv6Z6qix9f7bPEdPW41luGi7dsmUez8sh7YKSU0gr
q/Dv3onsHS3JfmfpNLM/CX+yLjRPwwmBPyQk/amzTCOhMAZPpI6S0jmR5F5zuV06
RBUlS547+mWohPF6bUvwkCBBdgoLulYkO+dXV59V0BQt4wJkNdn7YFsAYXY+4mK8
wrKsOBthD1V5WtxU+qCiZh5zfCrMQ8NM1k0dI5IBMQcaIX41oVKmdEMUYpY9nssB
fq6tx40rdgVhVofbYkETNn45xAnhU+toUB5ylnZ9ostBlGCY5kv2/YjTsdYTwvMl
72PRcRDvCtIn21IHCyj5BverpPBZDvM+ZYinsMsV0LAVFYrTBSdxjPxMO8T5Fqb8
q7Ep45Xy+Xht40oK8UIrjl4b2drk2lrO1RaXQ1aAqrEjBNTYYSPiyK/p49lLq8Qx
fQXjbripk+4TmCipQACg8PNaVufYitHuSDPvN82coskP74G41eeydtSVQkzPRWqx
d/uICI6lk2gWGUrPBavbczMYsZdYP0hOMvFQ3Xf9gOsCjH/1oOHghuTOo1wgAYl5
VUBhjCC/wW7uOwz4h78i1QOtwOEtF7fO5oiLnaBDCTiaPjHvRkDO3EVFPBtbdqyD
cP7S93ECXxJsP19g5ioYmKWpdL9czaGJVe2SS/cVAL6JSuJuMAap3AoUCkJ1I8mu
ARv/Mbe+eIoDtwwD5Nq2K0qp+cnonS4uB4lpEgt4c3GOXcUrU79kiV+5bpJG5fhr
3bgzEWd1jqy4IbfbT4Q/w1nrnTQEG/BUYSTbHr+C6Guy+04XzJOuLwjscBkAYb5T
dHDkcqnMEcVzqPQubYWLVC4qVeFm7uGDHuE1C2UIZ5qVxSx3J1D2NeuKOFVZvkjK
u1hl0m9QMF5X+ccMlEyeOzWGBu9yZuYLB/6iuMNIdH9vbluqO9TQkizCcDyzvhhW
JFU1Cq7xPRKJT3B6djSERorEmJMsl2VRDPtijN8tB7ZCsOOA1laXUuZ9Li+nVxke
PuxTxkytWQPKfKpYlqaYbhLQk9atD5vGFAkq/KULfYfl8NV1esmpPMmR/3NSaOYw
ji+6c3X7+CqR89K42921+ie9YAlexme1r4SbDVFOGDpxeZl4B1CyXQyYFJUvLPTD
BVn8VP6COS5Z4oHJGGfI/msbkOAAELSwfTy4+UL4x2X/awrDSKP+HuiaC5QjTdaP
37La6qRcWd485+Gj7QGKOHVA9uDCc3s7zKmRHoPnwDZS8tOB/+iDHh6u9KUwpuO2
HKrA8+1KLm8YsGUR1e8o+/yswUCA/vdpD97RRg+qSFjjYjAkuM++XLTYEGVSme+m
QldYSEF2TtbYMkWuSosJ9vcnC0IjhEb84zTMqgiUYTsIv+PPTGPZvKzAGnY4E8gq
sx/dUExc7mSQ+r3mhG6ttYGcMthMSYJrBuuQdFcJCwasleUydu2gMsbLpLAWRgjZ
TmvF99KoZeATzqFhfC3apM+a67YmEpfTpJ1J1AiqJIAXEqu8szHhvn4AWxvqyOWf
zfQgapzoo2QoqM00M5pbBmqS0gvqx1Yu6pqxjTvdKtSfu8X2yWKGre0fg5xEVZvb
BPpJJXYDmWXPrDoaCVa0BZjqnXmRYMgd6VHOr/LwYCyVqwRfQo3XcTaZumzC7g6P
V9+tGYReuc3YZNcu0eYm9QvyxHfvUB++W0/LgMrRI/igbqI4xxeAMfVsW4bSdFhl
e6JTtQwb6LdA0KP/MU1ayzp4nzkwdOaC+3OY7u9D/z9eqtddV2ziuH5JuLCH9xKE
b/3zFM2rKxhUXrc3fBZwpYhdbBEcJAs44aPmxF6zXyB4d/ewJx0twHVPo9SigXNr
lCzZ2XNrz9sEotA2lj70ErZl5OFbaTsJyL9QHQmVdG0qptfH6+MhAPIZO+nKZTLh
ej1sm3uRLkkELz5sDT7Uw8O/Rej8nwujeQ31sbhDRkxUAguoHo4x0w+5MiJ2EH32
jVjJ4HI4MW6wr/zb0JnpsawkCvbaLOB29NdygfREJTlr/xynn3lmqKF004RbuCyK
uE9H+9W9sGI0scDLOx8yOMcOp0rMUSi5FGGgldJfmTcRFUtt8CrDazDCREIpiVNU
+BK7CKra4mjgM9yQhP51WX5p9TPB3gXPNP5XMazWu7ZcIIw+QesY6d+Sc6ljQj1i
xl2ivOUri2iWZlnRmW8L7wy0Aj4hI5fSkg2sTIY3oKPB5Vjy73HMNH9t+JuaulpU
hbDZvpvdhlmNbpJ9nQEOWQVy8jz8UnH6HxNUq3sWWDH4rWsTXT3oJhxNMuHnQDl0
TiqyT2UXWn58BcU59IeqoGaNsfIx8iRdZTZppwcGuwBX+Z8QwfBqQSIRS6QgZAzw
Z8K32CCNW5qTxv07GQ7DqKkVN0cWGR/ytXCgsd0esPn7i9GdisIjkew+eMIH6w+h
E2l723rR0mHuoeTOQaWtL1J0UWl7lnbb+3OHMLt62yM7k0dqjfaTGVEOhNMRy+c4
C/Sygr4d4WH5jFnnwrrS4eEYYYXGMo98deeqOPZX5nfn1gz3JmsMtnOTFE1V5NlK
IXNJektaLjaq6yfJMJD7FkM8LNGweL3RxVYa75MxlJmMPTkOjLqqxHHFGiJ9Cppd
I/z1PuFqLB5Ue2JG2KVoJQLfHvWA8sHuloo70F6H8hbBo6YuFppMun1ul9VqtmOp
fQEQpyRm+FL0n7G1vWUJO1pNbYKv+CPbNlKEpcn/c62ra0cQxmFIRwceG721t6IU
N5E7WCNUx6t96TMtzEGEKeePAKMnRnnK9cD3WDZvuDIbMdYr4FHSfTkdg/UXqx4U
7c/dLEnNA1H/DRTTNO1QbYqQc6XviOt4RhiYO1KPqDGT0pm7XOKsfSoBuzzSpyDi
0en/YhPMmwcTICGdicA/zf7+CYXo4oSupaUqEjaX7OMHeV9FLdhwnFzp/8atRLjU
ru82lacGMXIPVAi63Ov8vAVLTj15EBaSq+hcmFVaA3KfWEzA1X9tQKUJWAvHuw1J
JdAbDWRLvPZyUn6OdtCGe3iG5WWyCWMA9fUn1O3AgH8jL19iWVKJFB9C5JYvfLYe
7ldsjkM8uS3QvGDp3KYh82ldiI5o7db+nTegk8vTQ18pGa43Hx0sTZxXSjEHhUWP
LCCJnerRKqrE2+kgCn28u0VCORTXlzSzBGOdIvwDNsnp0v3zsWkrvL56x/FB/7j+
3osVwowF8vp/dSy4l6AuNEArPpJ/ty0xBodY4bI7T1BZOEKxBb9JMv6XeDiw1UEl
w/cpQdcxFZHk/CLPCrRqYGkxk1rxra0uo7gyIUO55FT8FFzk9YKdhDGfAFlDqTwg
nGeBfj95s/yhMmTxqO8Op37INbRccLXYJ2PlCLWqvSOrMp7TSK/md6DVOFAy6/u6
mRxl5Y7b2o4crrzil/uklN2EkxWTBS2+UyRgOBtbnf3NGhrxZRKa24l7sEQk/AJK
8bMmvc+gjhUWLcsyT2E/i25G1iwZA9b2lA2dw7dQ1+8xsDFPfvYgNbV2ndsXF+RU
mmxKUt6/LaQlSabuQP3jOpXkq8+XdkYZdgMP6g6RFD/bRl6HxpLTAEq8Oq+/pM2f
H/9kWDxd7wW396Z/E7zjz1Jhh90rAJh0BkuuCKSw8fY9IM4dSPdmiQe1WBHfx6aq
EQqiEof065AU650wYn7OBrVoY4Lb0OnSW4cqZIo6buLSDUcYArVEZXTuVATBaOGA
2uWpG5YYGOhnPnf1U09il/aHZPG1lqeVnf39yGkuG12tYZH3Qb87vCgZcUMm9op7
C4571ZBj0EWKR88filMmY6RRQuSsWLlsWwwPaXeppBjDwjtBZ03Wj+j7ve3GQV7K
PjdvWZIk0WwHl+9GBm/bjlTUyFOU1d6fSLTIu1wjerMBnOlbxhjgcrZVA03rghyN
zzZRNOS8YuosYCyvGYiOuKpiPCPgQSIEwZVYNkLzA1wNoU1yejTOI8iWwnteCHhZ
bK3KzdNrA2kgpG3vsjS8BUlmRvIkFEpW04z3ZmOhYW1M5CwWUYXtpeShnq+lYzoB
w6OQ6hwOOPsjlbRnSCTPCnGgzjHeNLvqrEj1assu9IwCYAJ4MbE+vQM69i0eNc/D
0/CQbShKTQWSFi4oYW1lLm/a0hVmjrLiC50mtLyR+2Blwv+cuQqhHAFlR+6f99GM
wc0OWnIYFMeXWqG9JeBxjludbI8KS1YyVJnCxcrTyWJKiJb4EEy7HFWlroD+rhKg
mPLkxmvKZ1vL/L8hjNgiBXaq7YAIEfq0zmMmJRSrpWxs/OsglI1C8BKGqwxVGSLd
XDRXgvVr+KtixdZkTpHnLrLjUymfvww+l92N3hi9w7sPz78huMGrIL2RLHdP0/Vm
LJZ4yIMxALW73KtPnavPA1JAdmoROJpg1jB8gxLVHWglUgS+EmEALV9F1pE4bZFt
GZ3mKMVHlEsqnlN498DdHPIKccSFEWjkeO+yckJqsqmIf6/v7co+pAlDryj1nEbl
8rriFk9i+gydbW8z+HEMZeIiMj7ykJb4h340rx9ocPbjNNZOBE9pM7IVEW587KS5
Rc30UGOi7npwWlv1LwnXIr48YfHf5EvbpFTLcjP3BX2QFzfHy5Il4LUTpPi3kWjv
7BzDY/sTWYq8uIYo7RXzBeRUHDD4bj7OQrfpVKx9GOT8X5Id64xJtDClkp9ZQxg0
uU8V95uJFrPnO1UYsLFkiTgkqqBufYaEI38Sx+grGMA2vk8sUIZGkb6tET7o7Iua
F8/SIip/JIw0uYFX7dZmThCE2JDqE9rnJApYMQp/GO/buCYJX40vKFSwCMHjI9zm
ayK2taMa7DT4MIkgIRBL169C2guKpEx/azULCij3gpjGKHvL1a+JG1Y2qxJlIbAd
B2NLXK2LvLfym0+kw3HYuNi8rbeX6pJBDjVwdRIPb+FKACPprkcnOn7t0hYd6pjh
idSTcoNNKvLGBvmrqnhrqbXSLa14YL3dgJfZ2Y9xtcdxffnVwGQRzQpt+7b+LLRN
fSfjcxb3rJI4exDnlWh/zv2iU+Ph39oAX+9g0lw8lRGcPBfi9Ux716olBEFW4iIT
6ltPvgnkIlLW+Gh2NHJmPwuFSBU6HE+Yz3DwajjM7mHKgNx3gFzn53QmRrAJU2kh
X0iAYVQdkxqACD0MrS9+lgbMRKJIvJ23y+kFCIk7/8fSYNLHYLAZgTwvqWfFM2Af
Mgjty/FcXJRIWaSaiM9mP6qwLGT9sv9EB9CWTGX4DcHS8yDFMH1Yec/HhE3Nucjy
IFEsMlfchsTjhEKH/w9ryAo9jRHoFdmkCkx35Kqsb07F8HF1H2IvJKB8XJG94tM2
uBVCg5FJgfRLrWpg+mI85IficCafh5zUmLZ8qMYYPzzH86bFUQJ181OUr9QzY3Tj
AOV4VxOdIUHEyp0vI6KhBxv3pGaO28rUbbgRbSZ21Kc+2W5HYeTB+nk+5E6CyPhH
ePeRfxsOOyVJe9E0srMiTZmWK1IvmF5c70+PzbDuExuFRy2SWK+y0lP7YgFJ1qrr
x6w+VhP37ZHw/OiHe7oFg0vrRv7fBSQosPm695Fjg8zY5/PZL0v5pcNZDK21OviD
oISB/YcIY/UwRnh3jwLsLyLnzl7ovUEr9I6XZ+rT6iqVwb7B96LJ4lgyjKnLCGLx
stjb1CT2xF/LM42g8QlFU2jSSOlpyIX7JBy6p9qi75gURmj6u3WtXBxq/VMBPJz7
ttw0S4oQVC+kxgFDd3TH5MrfDFBiLUjFmMYENUjQ2DT75Z/4W2avVPLWIpxCrOXx
tvRXZQ4ZwIlCyCLN3pAi/81oTHFUBjOJxvVv+PnhmfZc6q4XB7Nvll7Fae7tFu29
uYf63fVrGNCtx2FsCFT6+bs7wdTrpeTAbuuD34U8Rdezymw5GHmlnAAzZeyL3R7m
XqslRWckEGvStiSfg3U+we0ZugA3lABWadSjTLaPtEJdyQBGYiSjelVaLawm1b1p
9/xied9NNdY29ufWt/VcVQAtqfT4pLAICa+qGp0iCcwvTwTg55jLdmYq6BjM8glb
ibrbJ7PrkR+q9Aez+2OBwE2bwZXvyV9wtOVctBG3Y4GibrZQflUSqT+ORt4kpyiY
v75C/0OFI3xsPPvFcCfZn6Xe96oxNdbcBDQnG4aWgN0VclGTKpaQIiVGenOEsGPe
6NBQ1J1gnviYAH7Zq3JENKd2hlQ+hvV3ERw11wFGkYolWNPOtzKbEbxwVYT5X3tX
faUZv1m4303Ii5YpeO9DnVxlWx6wFgzrMecXT9SbyGV837bDfUYMZoP2AbCVmzMk
2r09EqQI4IFtTiCQdqDMhr2IKz2xJ6s0sbty2uhORtgBBmV+eErrinUt5olnT5jE
6glmeZHxMYEecMCcxpblTOLCr24BW/jPo0I5uu+0NOqKG/RsMV9YlPnt0h7vdXof
Rjg13JULEbdsD8njOGb7DdKgh6118BEdklpG9lWzbVllBEKgMqYqqI1gJMOEIj9c
o30aCyhGBCSU9MvqCLnoEHvLhqEQvQjidYFoPC1se/ydfWCC40IZfu/STo+4i7EJ
eyRtPQ7krXPAy57F7UWq8gWQ6vfy/fwiJAMc9Z5DJD+kMb/LlREyl2AczWoonqEI
mIZE8ytylmQKk0NRxLz4Oz99tqYm5iEYuq0sBtO8/hR5ZE7+OFoPp5k5hyqtsV9r
43iPx8rAgJnBvk0aPD4+l0McZ5SbYHz8oRmbqeJQDz1KuhHDsF940CH3UzywuQwP
OeaT1s4N0R7R6wDDJJrMWAHqBiGZHvZb+PidaY55qQpmfe1dkcOon8xC3QuTjDAQ
Xwd5PhC+JDwUAJMWtetJwjQVSduLNkWHa4PgtcifYw1QxAZOGdfJZ3Tl6Ngwgya4
6Tb/ZrsnczCzI7DZx3d6R940Lv4FW4K534Cz/nscmxLsY+7fZ+e+z2USgEr7lqlS
L2L7tueCta+Uc1mKa9uceFaBBhwTLZeaFGkueSK7VQbOqAwhfXfbfL0mrkFT7j6a
qnGFjT4pNd8c4k6RDLT4L/w/r57EaDGPKmjfuoEzCz6hIOCnac0i/UKEC04d3wKK
2uaZUW0cpxCrTB5KHC2dBIqbgks/HVDF6EF8NUamKZI41328tm/CF+C83OG/QxDR
LgyH8TxL+y+U+f5kwyiXylHCRlhFQ65t8H91Zx9vvsNnG8jTdZnvW+IWEdaSNCR1
kvLV8bt24/gSNd2PwglikPbYWsNy07rbfFpsg5jywEyTrEW/zmbizcaId7iLs7y5
G4FCsSI1Er9ASy4v9RphLoAyK/b+ztqTVjkK3EilRrIBzaIS2YzJpayse5WkzYRf
MAtZHRGzyVcXr2dFC/DGf6rpHKnaP/OXEmwSyAS9FJCFHhyqaOYv5HzUOkexdz3g
tEjS6si+hRAs8KwPoqXmLNvyZpeJzsz4qD1RjdRCM73iNoJJw7adVc1DZ9lv1T/E
3gARaBKPNX4izM/qxm5FKfo2Xg5BQqLzq3v07Bj+GVHNnOZXFpyiDlQdxfpPL6SE
/uXDYXZCz9rh2p/irIOdak4ImcJQvA6wjcJON4ojbwt+nLotFK1wocPa958mzVxT
oHb868i6ni4qn5rfjlfkpEkujpTguHep3hM7laMonZnEno+ZOd5J0+lC1nz8jGAb
deviPCPF6h4VmZlkJGut67WPvuI+7C6riJ6a29xkAXRfvRa+2ncatasP6koOWBGI
qK0pseNqUDv8GL2/NKRdZ7W+F+3kFnxO1sdTme7BYMCb5osyRE4J53gh80XZWuxd
+8LBsyBt+PNXR9JyNXRHmgYrD5AJCvGA695SJiZMWUXgbAD8JQY7lI6l+rMpOwPS
FI6lSgJaz8+7lOFLUSjurfkUmajhrrZ/9NlpouA1WFF3L6OHGHuV4ljKwe2rf5w1
gzIc4M3LVcxJSAW796cJx3GPhq7uxlq0m048T/kDGLDP0IlU2Dia6Jt/EoItucF/
Ml2J73tkjlkL1nUG0wvYYO93IqsqDpbcAbL/Zb1hyxz29pKht8/TOiLzIuG/kzVL
vzySWyCHhFY0oeL0pBUW63bHVg0XRZneHftF5t3fi5ii6AV/ITU249grd++hKChR
n0twg/iyM3UaCPl71GyVvNMSkV9JT+2VOzQqa3+dQ9/fBR5WHgmiCJ8/c7q7E1XQ
V9cORX91I0cAsEZS+zyKr0rUJdpl614L2B5Fcd0pvostbnSSSiVTzja35Q+DOKTb
Befo1govROZGs+KvlmzRkADF9+T+h2EzarMtGYm7VCxZtQ04xmRcPZeWLOzE4arB
uVZFQDDOutFgiQ0rxVoaffrs/QezPKQ7cZRjQQda3WuATSAZLQGUjJwYnwjDDG9K
zxQyOYUgAsfLAfU0LBdCou6ALeqpY2WAZ+mu+cnWNpuDOvL9zoYzZCqIAwkUI7ZS
dNqaxcgUHiqKQIHlJkpnNFyUeINRdzSjPcl6xyrHUhdY30JUXY8++w74mAKMJqUu
LAy8qTSp2Ul3t0YrKdz81a4p5wYlZKHPfpRDtAHNbjTBKHP3rsloYWGpH7tW7hgO
z0yv7V6u4ceBHXHgPQPBwOF1CAsj8+JAvryfnpau+vOmK7v3Z/544ZO4ECN4GFsK
T4+8lsQKDSDeGZtEAkp0hKYeLT35ntVK7z59pjCGs0dCT61Ryyb7TC9ff5E9sDrg
9+/uM6xuCzjiGIcPLEELjyyO726tRDn2k1yS74ajbAOUc1AAvukwXiSwvdH52a3f
F2nMKKV59lzxjXxyodElv4zZHY+RPx+DD7HMD3fnVhUt9iQAqDmczRcVwvMnrCv6
Bc/66xmtgHih2kSHG9dGoBm3WDGrYP6vjJmr3+V7b6JAhpr6V147I9TqGdO6jS7M
8CZ3ppsL1CPNDG/WIFS+tEE3VntzDOUVupvDYbX/tJ/F3wrzkNEC75aBkAgNay5G
vIHzSZWvRrsbVuBUG1zfUsT8fMnP/lDTLLlx9eJlxPn0kqJ5Q+coeuX3/Rv6qYmj
qLTIifKR1DgeTv74RSiDCpf/GeniEghO3PeBiUnwYARM2D48ZiOmVnmrnjVnMUUL
kfWvZHi7akhtbxPYVMHtYPDRq24p2eIaLONvChnPnk+idS7NZISxoDrZlpb2CNFU
geUuMo/qDbGTEJY/D/ptyHeDIzD1ctodOXiGiJxfIA2cWhXtubsgYVctCrJ4bBZu
OxCs94pFO8hk0D/Z4juGqWowaAX5OizFEtJ6oDmTTAzYy2NFXPtJvqsyqsPBc0lr
mI+NFXLqKg7icz8xfNiLyrV37e1Nb/HM6QOWVIC+tuYVam+j1RVuSHACqnasWDMr
fEmEnwYIOj+q3X76lKwlAf6UBsqda6uoFLYvKArf9G48YyusxVxLTNfK0xYh8N2p
x0vmNytw/kCGwTcBDl3iQAsIPMQpKFXytfgg9XUU2n68ZnKNSA86ODwRQbFVAf8L
q9W8IOmMN4YR3cLT4RpW5ADxlZpCgLe6P76KaWlgq6ABfTlNVeiFNMh4GhZcbinQ
+dx3QYzThFLzz6BmAIhQu5QbPMfW4v4axd8GyxhZoZHMfufck306J2HazOEYQFkF
Chn5Wv0+gnHhRluilOUaWSv/JJCnY2WoCq5zs6I6jeELAhJXuyX1Vb+Z3RNCdMT5
idvA1X9w4B0l6EWWUxFs9P+Wt6TldmFZXvObwKbMSz3octUfFIJJsiYNllWzKHiq
ughPDj8yLxumqJKquF1/EQMF7jmwY1GnsXLOF3vKixBvx1OP71tWv9z0aDj+QF5Z
v4B7P3By1dRtalWoWz1GgNYgmpaz/sra1PdCAtgEGyimb61dKQNiA+3a8sv19VHd
oeiQLNnzqOi9HKrY/JwFlyQ8UCBxviddqimMEN2x5HxKigzTGBihYRrcNG0c62Vo
m8HcNKuXn4DWPXsuJVnk3gjZzjhISjgb4S+XBc8CBUhOOpSNotlGMYxiBlTWLIpf
5/b5EfZ/Jx9EDPbt65q/l3EZbB+tTmTQWmN/V3TQDGpVsbySAQwJC9EFNGirAOpC
VtcDAGvAf2hNBATrhDE4o3NVTMDQpRgm1s+iVQ/CBa/L9wi8WgucGatGelGaf4pC
7nx3TcKUOr03/Ybtmho4sjCn3TFpLW3LO8w8Hoq3l3b9xWu9ZbFbIcF6uQvQpcaa
W5sj3mAljd8NLQztCYBXUrUiatuTmYm5dUfUzHxoMDgYzfUAbNkaNlViStXzVR1O
1fW7Xwtk6cSlV4w3TpwiFWqMhuukmhCuzJY+DY5SWuDYIur2bTt+/dc7nw/cStMB
ltNQFToDndt00glZpUD3bVflyRUnqxDmdayZsc066OJLT2EBii9hv2q3pVXMH1XY
hmu0/1Q8D7B2QVOMO6yOT2YDtM0hw0w6f60Z3TswqxumDdHFakb0RffCuclLULu6
Qpd4dm3RKFXusjzAictlMjtWZqnZD2N6bL8/OrAPN4NZDGr5PjBtAPL0GKJCUaJ9
gSktzQa7QpaQrrWTBHAiOuvdS2a+INOcIrkzKhPChfdHrvkTikUH3DJs6E/2VwWG
mwjCccvVLxoWPhf60IdLEBLYpLqKVWOStp2iKQB4y3qsBO78hFldHrW24Mxzwwil
Id9ft2Kw3zYiYhReEOPymkvFxWs3u4hrigv+mRYBcH7/qUKklGMIriMMsqb5VRu7
ER5H6qV+tJUmy/yY/fGVhv0UpkWL7tCAjgUDSOUYcdsqfXuY7proXOgKtkNk+Th6
TwUVffxqoWaRZXlk1PJJWBI4OlMAiAHo9Ls94gYZmKu4yb4RXp+uWvCcGaHw2z9F
zoy1lTUj9yH+CWauwmmJaA4YMr3Ct5/l9BJpbdmsHFxRJKJ/wDnNtVb18DxC2wfw
1m3V80RZWO5Kg/WETiM5y9j78ueGSApRbHGvoGagzrygG+ugEnMmwPKHM+gNgbSG
IQJ3Kh06F04u282Du0lDHtytcRyBncw0zfrt1+YTKsef+OXXoFd+UjCKwsMivxjs
3KOdx/gWp2b0x9t7F60YnRx2g1YNsEmMbA9slxrqPmachC3f21/wUJhExwt1TDVl
qPJ3LR4Kp5VfbWjuQZZbv9frpEXYQChHd7QJDeMr+hemPeHO0B/xB6C3c9q/RR3q
0Gd/qIv1LtOqJQrhEzquKMhjUMkczY2MucnAP9febGRfJ+7KRhk17zBONQ8ilo23
pdJEwoBArXH9ACVggt+4xk4lDkSqJ9BBYI76ja/GgY3yu2Ful5TKZ9mfTl7g1nHN
7/+EsA0Jtlrn1y1eduM/Ei9oABOk6KphWETM6y25cbWuhGqt/gOsliIA0E3KxCqS
v/8uB17QQtR9LI+nv+JgS3wulUy6BfMaDD6eIW56YjcQYDnGff53ugHeiIwSkBqj
PnOYJceVrMlEysGvsQAsDpeQTf8TKDJMaq5xmrPnC8DF6AlfOsnO7rOb6Xg84zUb
5I/Pvp8aoI+16/MxpbD3rFARt3IOV9BHgZzWUY2MVJ/oH/9+kpVsBHwsuKh/gygU
KvN51pK5nO7L3VFof7bWipcdf8wuzYNmaBZ9Zm9lfdI/f1P78Lk1Rg/ig3YNFGJT
xR4t/FFfMNRYUCpRFigSf+RARO+dYrdi4OExs+c4kzfjNJevM7l1B2fiFBgfcuor
hjnnnDol4IT/PAJUw0G8bkGAVkV3U8ZHl96yEr0WbaFPEScMdmhofrVK88S7mXB3
+UQGgt2fHm/wq5gY66n2JllZd2jJBndqiYN/eXTMcsOhiDVNRPRhzQwL9g/gNdrH
Ha82HLwsti3AQ1Z8eu3IMM+HIrbozOf4XneFv5z7HoTEdrxZfVbAKm6t4fqo6+JS
dSbZHLTLD2qPDOzKSRuKRCff0BD8IANbP8Xg4jG48gFNWPhP1r5FKbk49GVYjl0v
Xjs6fQqqRT7BdYzjZVoO4K11lQbOBfqlp1dfmAle95wlMwoN61KgxVM3FHJ7YD36
jW71Cg2PTLIPSBTDaXYNKCgi1Kzma8j+HCK07XRTq6gpptFBLmPL7JCR/rlJs5Yr
2e+5slTo8V9rPO4dm/ZUI8sa9khV8xCmah/xYllUsJpWGxQIF1LGAkH+a5yDfiyz
dPCwZtE7U7+oeuYdsdZqW5NVGPtpFJYSaaQ5f8FTcATqENZDy0DF9/glvj99yniu
ZxuQpDVag6BLRxeqN/q+ceg9SxRYTZ6xJHbYht7fX0qrXGz9MBzxCcpZJvdTFIpE
orcZkd4gG4xnFjEZXk5CE5Drg0vTTtnTvRsG7I9gPRvcQxYGYyLOPBKhYrAzUPv/
n5LuCctwO6wKqYYPgfgqkgdAYmSsaCqhdW2NO4+6CB8vuybmyzWs5wX8sJFsX6fb
zId13QQlIfVHwy2nWUk78r0mYFeHZiXBBckjgpD+NuY5nZfi3wyu3QlSi3amEBhu
XoD3KwjUgiRKPdF7+5B/gjxeLxP0bdsSrBD2Zxpupsv+WmjLY+u4xfU+vd+pOQMq
uARbt0hs9yVk9PfLxfPXnjip/mB8JhdJ2eM7n7UFSu3T8xda3XNuDKjGp5y3wLzq
0lS2+8vFml0DyQ0TA7Hj/o5xgBzgLk8ByEKPjgF61+vlWe1m1HSFU+P4nYGJVCWE
Hjb7S2rvg8hCyhLwWMbSprTE95aXra27R0lAASafxKLoFaave0lXDst/L9t6d3CY
GNnqCQQoPzmViv9LtFdPWQ+7MQrFG+AhC+viGpMBFGNw6G7pA/DUf1VsHKXHrMYT
YxDEceHE7lb483m19Fn7jIqsUcpKcwpAvH1rU7QnuA/7X4T+N3+rICFNDcl/uIel
qUsquTBtabYXZ2RDAf+Fm7BnxLmL7SAXcDRK6Oly0hWpO0kyWNzMAXivf9uMhTEC
IY/nGGcLo7RGpr+qg7TKaF/hOqkBgs6RM0d4MSbCq5lZ49tgxU0S5nkpPgRA8D8M
c+2B8j+modvBAFscX4msB5lbndtxHTgK3J6Sexr9zPSkF/XDbhlPrUVxQALCG+Br
+xGQSUY8yJCRtMJJnkW9bHF/Afcca3H065kNX7mpJOX3Q74syVmeW/3DOVURr1b8
MOxQXllfjZA9l4UBK5cOJxDRtQC5ixSE+NujtRekAAWwiioRISzx/C5C64K63RbD
LUg84zzOEqBnzjJCDYmqSLdzIDZ9Srb75w9XVegqD9OOJtgtvWNLn2djCjyVHSRO
M6G5MInQTQO8VUrJ739lOfTK6GlqJ+pzmoXCMFY+DKuNXqJTa6Vr8vlVxZuv3Hpb
tAXFUQia9ZXl6UhnJwkU8Lcatf8J+QSuKtPq2dLqdzs3JEkW1ax0N37d+ujqeuST
kHfGlssDjD7EG3mN4MwM4W7yXZzgj1Km7z8LPFEEnFSY1gTmbwYl0M+qd+lqXSFL
/WzgvJ1RpsbrxhL9pn7xD+wL6PfpllOFraG7oe51SmwvG+F/x4w7JnKznSKZeEwH
eH1v7rOACK5+mfly7uliszf6bM7aNEpA6GNPJiu8TnONAZ0O12cPgd9QWnlERvUT
+UlrdfMV42q1083unCzF3wz26Icm3Mg6nai3DGMnrOVKzoHOl+pbwbEQWAXb9VCJ
lCQQu9FB6QNOM6dQ1TMbgix3jhiKQah3h+omImEgpTISWdnrEC5D/b4nA5zpPLMM
X6eBIXi9AvLrfal/xfYN/D1UTvDOMGwpFUyxauKP4GKTxBQk9yuiNGskE26nUZQe
Jk5aRL+132+XgoYe9eRZsBVXZHwZpiQqlxQpYL5b6nEBHGd5txUe9RciV7Uz0iju
QOd15oDrtKQWR2vwKqfRiUoewp6rlgpzrUVuUTMTu4EAn/J/wK97UwY5YIzYbMQN
pkXFuaYt+VkKenJVjs5UvM3Kscyz1IqLm0GuQXYtwBCZsLIP/FG1L5ZUDrFIJ8gq
iEIJXW0I8zP6GSHPLh6IHqRfspGJpLWaEW+URZxx+3L+J1chnfKhKaTxDKHcghO0
ioa+3FgL3tTvD6M6uRaoxYNv3y5N8SkNwdTL9jxH6A4LnZ97txGdFOy/d2ptIOQ4
4ayynTnvxV1pDTW8+rvOfZkgrtU3Zs0m6kjNgcIaVWLX3DI412LfQx9Wf2YeL0os
IG5A2KqNQqt0Je3cY6R8T3AS2CMXk8lz0u9TIDp4nUuK3Dwx0oPpsOinFUR2CMnE
ehxZnbHrCHdFJ9LuCAP1GckEPqKZe2K3xB1NcSaETmIged6FUStVkunvdp61mOxE
wgNQ3NBS2iXJsZXkt1T9j6Fej5G4PjzERD2T5mgnJGVZlL3nFilptYKGxITxz+yJ
cs6spjD4tEz9l6pREfQwuN82fsgtkCXXIGycqa/5By9Al9snv0HHM4EXV9IzUlk1
gST8dP5eREKxS5tf2wZ8DtHUUa1zxsAw8Y4No1tsqLmsFiP3OBqv0YLocscxTGY7
EZhHrhcZosiuFh52QgGp8vopHbQFQSrmzQGfHPeTTEuYScFjE7Q9DxDoayFfMkWx
WJ4wCfaTPvNvVRnpdy1fYqvnSyWNRmxuRFY75OfgiIXZGw23bqwBE1+ozDA61m71
q5ClXA5UUiA0lOWIrjqLcpBthm8sW+Kl79dwQbbStD7Y41k3XLA0lj8vwauUk3PR
46jIYNP6e3oMfdL8FV51ZQBVhS5DUyKYKzJPnv1r03aaFUAUQS8XMdjHBum23qsx
Stn88XFMWzIYhRzPm5opGwyfx803zfI8+kJV6s8dQkd/sp3FiQB0ExtZtRiSOFWm
9X01Gv7NjqixFNsSRuVOuNU9RtF6e/rK5bSco1cP9XjFyssiyXdgPcKukskX6oHH
dQO2LQxDxBCkGFs5qSOHxUKcR7sKjmCwNHIGXh8gnuL2ewFhTaH1jGbd69itMm5n
zr9KTYLDemTGGnhRvLxrIzz+npLjsWEFPAMMYldUdrDQNjwVDttIKDk7gAWPaVs+
LkS/S/g47vx1pTr6rBMs5oUv1pQXiICmDKu0aIAyBNb3AT5w1SXiVZ80qMZIqXS0
F0a+DAXXzVQjbO7CAqtZBzLU4BYI4gMZz6QrXJI/1Hbcr/xbXG5RtPuJ/EAoMGwd
BiakwFYl/HOIu/jGERz/IbYmXQbJ4A6GS0a5it2ctoSwAd2CMrqgM0lfmqw1RLan
8XUEgGu6cOZjuiYxPNwmRT5zo2NgNKjbjmjL0U1nHck1qomyRTXNAqXnJbLEt+UI
jg5wp7kJDsRoi2ZoRNoshntHqlURt9CQHwdHHRmEc805k9Q5EKQON825Pl5sAR4i
zPGMhtDf3D5FB68QY3X1XKaCAmRvSrHHkx7EbVASm71jNgpxV8tvyMmTtG5LUpf6
on5G38Jd37XmoyGG9BoJucjslPLQSAjftkA/f9Mn7z3DVvD+sUJQRjgnJKq20FIS
A1DRhkXUh8IA4Ql8SgTn4ADm/tM44DnLS/D5E79SQkU1dYZxJBadMtDJ4ScLBdvz
b4WHEU1smQnutRmHkg7Ksx3IcK940ECSYlJLLNySsxzpWEHyQx65J9k49zuGyA28
YLjA3NoH2/lclDoykphWbD81F70xEJhEbIKsPN+avqi0vf7y25Z38ZaYhDX7DtJ/
8thu6fzjkpg/ISvlK1bYEd7Wu8iyd2JqemL2tsByGC8=
--pragma protect end_data_block
--pragma protect digest_block
W/gDp+WRoLMDAWC6vmoJGUTrEEQ=
--pragma protect end_digest_block
--pragma protect end_protected
