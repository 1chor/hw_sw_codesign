-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
U2M4lMp8xLAgd4GXXas/tQd4uvfhhTYmNe1xtv4442uypsnOXMyUlwDFx3Nv60GA
blrzfoVbANKuLYZcqUEP4CLInh77UHseUhAAixiKofoRC09QiH8BHS3RbGMnyAij
diiP3ADacGFVVTzmiHzlbJl6LZS6BRIxuPnjqYqp1/M=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6077)

`protect DATA_BLOCK
q37Yuqy5nrYlrFAAC9C5BK1tVTmHbT7e+vE89ERG1VXN+9kotjv01uN1ydISk31i
T+gJG+Y6o1B13izkAyAdbpF+/Q0qAmlPDBaing4tqe7iXA5XOz3e7QL3krQp6sos
gxl3HfwHtd3vRCIrEQyXZONgw5UFYxRZy/hztKByojj436uwg82JucvRdjKLaoNX
3ZhjwygMBi1qgwjNF60VsbjV8E1jhbSvhaCcFGebC4FHHFMKWDGS6URs+dzeZyC+
YtQZUWtoPQAcv8BPpUCqDDbPFWuYeabrqb4dhI8b897CBLeELy2GkqdjbDuZuVaE
S8EHjwmfEhX1uyWRkbJQ2oZvTtVYIEZNp8kWc+58xUAvdobRVsinhnACHwOYdD/F
sR2Pew7H6QmxAiJef9yGXc7IxTyupkW1UtHuxya+TKqXO0lnaZqVRmopdNPpAUf1
wtAl/MgvaeDxYKL83OIRnuJCMu2JQVidsxi2GZyiPbjHX4YL7V72UapAtE3jGh+A
VIV9kqQMHJxlo1kicQDC7CtZueE2SKif+SsPS4Sujqjt2FGm6lEphNwOJxic+X5i
9YJsPy9biFQY5739XvCUaIaSfkx9lNG+BRjzsgWX19llg+SsyoOYs0NI6ht7Ioas
r+xHsYDdfoAyAqPEBO99OBajw6yJfZmtis48cZvgUEsxIjwxbNghg8a6d8uBQ1YA
y/JvPPRrA4nuMY6SN6OsG4Rsp6pQWgAu76dTgg0jawEihYzK/oXi1j0NLHGypTTx
WvBtesTOK+AGUT7HRgdiklyAzn/lyJ3+Cvo355m9KjN5RmDJ9q+bNPURsk6UPjvJ
O9I3PRgSSUcIAVCX/IIp2Z46G9VwVosOaMw8qMIhmm4Yap3WoZn38+a1g7lzrJoR
JxX+H/2hsRigcAbKr41ec7VQFP3KaJvOulQyjJxuKxJ379vAvqSnc/er5UnsnlHN
nCKrQxCETQbuQl08hGIg9yihyCF7C8kffx2lK3tA0KzCsterzHjDUNLz0CuFXFAG
fWHB9MGteh0DAc0K4ZHAVmKvjmSyfdrK7qSCiXdTVYpyEHCqGaeYbemdCUdsSZVN
Vlw93BaenAfdZqk3MQX9nhDWB2lXe972YD+p+Z7Yq7OrWQKS98RYZBuP0hXuiXoK
oMAR7rb6dWd5KiD9ZkbdCGFYi7+uKqJ46H+5gTuB5j3SaiGE9gRU3SzEaE8veV55
bjDqLFCueauM6tq/1tf+lDht7vb7VKsSkMrL3Q8vEIJDqAHmklNakub/Cjr4LKxX
2GPKeSyewUbsWucRFcqSzTFJ7vimsYq0RsccUwCI/5+iQhhs9yDW3+62jhep0uei
itq23ApHh835EmwARRbFaZgWMNUX1e8ItaJzug5FY1FPj7AfoEHYcQ7trhuTrzNY
5bTOxqqxf5lSUkFGPFcO4SzjCWykb1LREKE6pul9feLdoWlNlN6wTNaOCmdlKvQ6
vVt1nRt/XgEqFdRXlTNKV4hCSUM+Irm6Iuz8MN8bjQwkgtwnN/0LR++ExV/EsN7b
cQlLD4A5xn1aALyTJYJHn7eg6PBl/kF+zx678+853fYMjJTuwf21joes0c8uS7sC
BH9tqUw6vMXZKi1ytHD88X3P52sy7k4tGRn0RWlaq3b+OF5J9tmopu9mbNYpiNlq
u2WyjVuoG09ylrmEbVTJHSQk2E2YPI92SO3o4NLTpSh0+XzmmBFTe/L2FL6wpWU8
Tdc16VEY718vi2Tv9J/9THn3AmPGkNzPCzIa3ZTfkpwHS1H65nk/4hpq7Q/sXuE9
d1WNsYE+rtpFE2mgNeazZaN3VT17JinmOYC0jqV+fWBFGiKKlP4zJESGDOzXkbkD
fop9a90AIisp6TvvsskEjDinvB2vMHxw1Re9CUwBf/15Gt/U2ys8fgIlkEtOR7N8
QprQif6r3p+Wqqa3lUrcLPz25EgE0I9QUxeZMVqmpQtBdue273eZUteM+T3ywncq
A8TF5nEG4r7nycDten/k7r0Lk7bdVOexUY7cqBz7Mw/EEWclvnEBfeRtBfgGExEW
JQIlfCZ+fyO8mXbPYBhbrlmS+hS0/SLUY7DN4WO32kmqe46LaZv/k5cSqo6BvEXW
mmZfkMvbc8zgdMQzGB8QFGvGQEe811+LbMzM75P2XG/zMfa+JXSGeMY0+TzT/1oh
I0s1LYPi8qyb2jQxCXJ+QBddSGFI+/tsvUkKg+6Hjoy2gRj/UkdQXc+a+FO7gK+w
mtfsfIlkFDC3vSTmS3ibUfCzaB2Qn9jh7N190aoKpI8L0qsIjAimW2GtpnrkYH7p
+R3NNuMgvcb3XMfqll20HsdaZ3K+4gC8b2Nm+5cyXyDnmDqe7Q0EZvoRgHydLrG2
49OWCWW21kTCak8XkpsiIczUSI2gvupOYOqLXVMDSHVOHpKWBN/U9OSEfQ4RHcKL
sUr6sLBo0LDL/fBBogG6AHeL2vJjvbGEBViVtyCf6AngZAbugWfWylVhnhbndiOk
Advv2i6RUswiEn+/ccw6yQs5K0AhyJrBdWCqORn6B6q5Q/12YGH0tlx2lLwTcqmc
4mKwr3FqbNQkjfdt87V1TGv+jz3A0OaYkS8HTlvJs4mG9bIFQ00XM0Oz2YRK6aWx
Kj/xXvqCPXhCWxOoOyMqqtStR0AobsSmV3UQvVWnsd+NlwUU4DCqw/bZ9fu4Cz1p
P5EfxB4DEUjO+4OSpqNzzSHx/qrExeBO7idIzOVznPDqQgyO3kQq3MEerTkWIpWd
uEo2B3vhi/2joaiJO3MCRBw2CRt0aj0nJlU3Xbxx0y3pRCMi3QM5VXpiJcWgQPYA
mLhxxm6ZdDKGLYoKCaMIabauI73sEaFLC5m1nFIrug0EwfIi3xoXpy1Tpvm0qKQK
5dGiJMDv7AHUR9rLNulrg3ZT8b6Wr47uiJ4O5kzch6PzQMp5CdCyFuS+VU85BiZb
J1HWP94sH2/Eu02zVLzGx57hx1b6ylzxhgY6Er1zIhHleSFTX7q/ZkXMLAn7WiIX
AxiXUedayFphy0Ju7O516ap+rlrTzqrXtth1MHHbG798BieLjnEDxsmJlce1kWwF
UsoE1GIoJ4r/iyEqg9dW+vS3XjaskHpSqTgO9bBEEKaDUaNjHq6Ml79WuiDrfkxN
CmpsDNH1eJbLzR6dLe9zqHCeVnM5Isn7s7eXC3FzfoFF3UWx6TX1WJF75qNXqIOT
k2MG/fYCKP2rjxQUakpq/g63PERMkMTfB+FgXGuax1m590j9Jr+0DllLbBGANXqO
BW3ARHR5iiIvVpZcfBv6DIvn6vnYzkprj2yMHaHWqE3UVSrWm6Rxb9VO6ausGTwz
vzqTUmJ47WnBbcsKpJWDEGIXlSfvpQ+IaDmK8tXmT/JpCZnY85s6Cvm7mrYTSCXZ
5oEsRhh3zVquMqvny9VBxUepC/KLIkvUBTDO/r3BjMF86eNpPEV9vX+2BknhN2FW
8bxld+DASPXBqeknHtY0axhaKRyXCCjSpx2BP3qOj9r86JhmADkRj6fcDvBjIu0r
r+Z5rUprTRHHRj8Pr9SGuBETLqJKzGeOcchMFizbDkKqVSu61JbW9nud7nccisxu
vDGe4QEJMQAtPIaXPdyxVw+LPtcpNJXUxAHsz58wFBnsZvUcbZZFj4OYfvhpzi5Q
CNh0n4T0FZ71yRIZ5nx1k/4Nxh54+VK35GPMkwvRoKgSVjf/UPDDm8M5B6etFlXs
gAZM9f0+/HAiTJrmhaL8p/DeTEURWkdqF/Yb9GRUTOK8zZwv8iLIzbzd8S+p5e9D
DjNAStbHhM9mZinEPs0LHNSqExQkO2broIRmj1mF5PdREbQ9sYD2eZfwLNZiWy6o
ZJA4xmVYguUo6Fa0l5hqeJG2mXKV/SLeHTL17Q/giTjf1+Hy1PLqcfpg3MwgkTax
PhmI60TMieHz2QVhmC1gc88k849VCKAfsLAzwZld/t09HWtlJk7plRE9Az0/akBt
Vac+QhF2vANhN4FeZtFd0/9mSsvF2dPWMHog47niRww+ISyGXA8MDrzxZbLm5LFY
YsHPJW468DASdGHAi3QW5CsHpfS2xDmUdGnOxsxnaW56gFvJLyKN/nD7puFoDxe8
HNDX4JYSj9XAXaMAz/EQWXqkQR+wMzFnta3z0ifqHoDdMCkm2o3xXsDK7H2L+jlD
vLz+6iKx48W8BUDgCRJmtoB19VDwb9idquPYD1yNjRDV2LRRG3K+Z1+oUrAB4LI/
DIOiMKwtxlxTmV5hw4J+AyMKSUdEeHwxF3fwsJ6CSMgJDCogAe9/6VnixuXQF37P
E26rCXFowsAU4MmIfqXOeNi7zdvZ37mrWBHRVw6sosilSl7Wou048LiHy/cBW1R1
MNHBWtxcrnio+GSZbTJwyFH/8mlOai0Af2mzweLJm0jYz0B1EgDbH1VcILe280mp
8cHmr4WG66eQj6VVhUuMHs515tZ9A+YAMVbxcDwxk1KaxLuwPzwv0hjwFedsRQqG
HLFYeuPim8GbTAyU2HKstT2wEWZ/mRheT5KkkJXWwcf9hI1bOYznfHP8+WnydbhK
7+Br6Inyen5sDnwfMW38NyaazhyLImUMopLey3suqrXaepafdKF+9ghVYOuftLxN
9Okp3BXOEDtqpx1A9hDGDra2fEqv9pHDhOjl37zR9mnVTZ4aO+RzCyqYQ1yBNXy0
gN+jgv1mZu1N8RH67pdnzs8MnYx6gxQWOEuM/Ltfb0J/bShB+eH3MqKPS/Flr7i2
zL2JVO4pvEhe4ne0KMg96YE2513m0y9ZIpfSyj7fWwDRnFu5nYayT0KrhwY8C5/x
o6H/fcCvwkdKWh8TKwib3XUvGXx+DKkqCL5hzvAEY7QdLEk92mC/KAVqhjVb+0Er
G3O2wYT4MWKk05Bvpv/Kqmk3Hrm4wq42pUoisH6rwpf4Sie+sJJ0M4Uy0dygqAHG
E6Mg+Fe4eS3soDGorIgCZVSOCL+2orNa3AdAr3BEJjX85w375LZe/1YBtMpbQ4SC
bCs2kWWAozM8wPew51gnAIrAmxxxtXIqbe8b0Zrfd5K91UhBX2ulGjGy4qTAqPC5
N82TMYjDk4ot1NpcUFjq/SlG45ves6t06LhGw+62apbFZUxYDBqBBkzCIwfIxijp
/abwO0twR5quzSAHJJxILulxbfREpbEXF155e8i/TYYupjJm932j98V14JhY/VzC
Dcq/UWeW1MFkY12a2S3/KXZPu/6+vHOq5SqIOL/OmX/UqI5Ps6LuLY/7DiqIJj4r
g4qdGsE7CkR9W5EZ8Yai5vcBOpie3qyW0c17IqbodQ+kmj2o/XD+4/7UEC1EgjPf
/dUj6VIKk0TD5sqJwBge1d7IyCkq91HQtVppauPDjFCrYMK6M9YzkdI1tvG6hEhV
E1+N+87Cws7Ry9MvSqNkrdw2/BoN3Q/WzrIsni0e0ncykidzVINkVirBRdvTa3Ar
X05PzcS3sbyupojEMxqenOJHENO7IqBiQYQrjA+eGGFn3mssaJfKqVX15rycpPU5
qomnSGWMu7THgWvXNS4qUjlvNyP6jAuTULV+iGoljXoJl5C9M1iVH/k0Om5+2VE9
P4vFd/2tch8vEkjXQHTZwhOg7ZEZNTcnoyHF5AjycwEsezYbbqX6TkidwbkdYsSl
QPzy8Wdigqr6ZoMGa0YTu2I9xpjeOXaXieW1jqEkGllZyxTav55CuLIfIzTAHITK
WrDWyJyhYkoAILNuomeRUhFf9VopYnzOxX4BcACnHEbPoqU0e4IQPcX4uw/HuHVR
RyARp2seIExJZOTuNauNxiaB3S+mNosmS6uLm2I/g1g7MMi4bPh8ApmXO5GSZmK6
T/HCIjB4t+9vU4c3/YZSY1+t7uhA2INXuy53sDjKxTolGNPioml09jxyN3czvobN
hcogHGZ5wus6AMNkPM6x8RAX26JS+H2Xx/6Yrfd3yRqQAYs6cgwt13T9RHhW9U0k
7q0We2ehPpxCs8AD9j4ACbJFOq8apjLerkz/nOGQ0Aa8N56VmSx9guxKbrYoGd6D
JPudpO0vHXUe5SGKUFtHAFrbAA8WN5kJInZFJ2Mwv86Nn5fwvgBbcRxj67Trezqp
RR36Ba1TO9nv8Cta1ahF4Iwz8fVB61kdad8JHXdjvDkGyLQjELz6r/KmF6XwmKeC
N0fM1iNFD63/AVJ6czlH5HSrOn6VhwkqUlnER7ONawnV3yOLq9azJgb4Wpl6Bn9+
f8c+Mj/6Isg6ql4LBwdrlBbgBwO8JLhnTwBo/hKkuNx8SMy5KRIvokdoVCBrUUfZ
qwkdhHybpgWsIjM6jk7L3qij7gxddXRKW5m/CeMBfvgbeikZRATXxK4DmMwfY2Mz
OQ/d5wX/2o6FlqbxAIl4Aqb8iXHSx5tGMtd9iVc3F0n3xtXXlxe2HgNaQn391HVx
Wb0qoWTkbqb5WcvtSYWe3nY5klXyydeIZ75k5uWvoxqfH27kopDFhsVUpsxL2hGO
YWFKY4cbp5ZcjH8JW2F6QNEBugORbrxrZmxPV9Acjp0lbLp61BQlFlwDAOFrkEu7
QmI/uuVQNFUHLis4HM7lE4343rv3eUQkcEtGccJZk9WDnrJfNn1y4ZOY0lIW8moy
SUpmDltwUuCKs6/f9Q3O9XzAGqos+5GtCY+z1iu9om/00o/UgbJ7wn7uODo73n4Z
rE0OqLxw+qe2VJCyVNrW/jXakOU0vILcMwJ0O5PWA9+BDydmhXv3z7N6nzIX3eqV
EjCQJS/M09kcdKOjgJsJilrEiBouvkCBlpXLU2v7Vi+8CQimeKD99dGo3KaE4aCz
WzmvVId6DJlII6tV94NqePzPcJb+qkW/QE0QUOtrQ+mTPkscuvIvnfAmlW5Er4Eg
BU0xA0fM0rgHfZRuepAT6kVZuN9JVU/qNI9asxBksRGgRCUjaSrD+/8iW/2WPHsM
IHVlLPs+E3Mn6DDGMr2OBz1bkd3MgjUIqm4T1TxCOhK8Vjiujq+lhRSki5Giy1OR
IuKi4RZ0TYYjzNTzyGvxHzrKtCT3HCINNABe+TFhNinxG+uQTPa7LF/mRGJNSQnS
Hq30xZRI+uvfwXDD/OSWJ+xeSbuBZi6+s0JCJOYhHuWPnR0L45Gm/GJCvV1jhCNH
DLZyzHJC+Op5KuAvVXt7rn9SbsRHL1gHWtD+IVIon+pmLaeuOhbBfgFdW9QLMo6Z
uaMOT7EmbJ3Od94DBi1+hR2v+Xe3jgiPj0XLRJ87P5meH0LpCwgyUo9ayDTVhAZL
A5fn/cCA924SHi0RsNQe9Qt1DnVNinT0he2iO9354bd6EL26pd2Rv+BCgLSeiD6U
xWvri74wPlPvFvzo4kt2sfklpeXYiqP+O6f87qBw9o3NPHqWqQnHvx1J1Ah6vIK+
0g6amt7Mx5vEx5tIvflunx5z5TwWYGY7ZSCVWHg9Fi9Jv1OJRLv+sjHqmSaIi01b
Irw3TDEpIJ2/kVs6KfPJwv5Pd+fO/HkNmQooq8NdISRk/FydZZFqsu+Yyk5GGXuD
mvvvhZ5YNiB78oOaNRdqoI+X/8nFpI+Earua82kl9jP9P+GZeZzoFrod15/bRl3X
gAsSlMSaZ55e8dNlpi+v9fTqqgelPkxSPsT5nNkjwxb/9n+wJ+ftK2pCYgzlgB5p
HWDeOqZHARj19Sidq6U8S53Xgcdo9nHKeuKmwz9PGUPvK5Kb0PhuyJalYG+/xNhw
+9Pzuu8oKKGYTbEzmZgkoejcW8Nb4iRYxGsyAVm40vuVOJdE5ouLnFknrxYYZr0k
tZxuSF1S02sMMCRguPvsfUSDkAH1GnUijlyV2xJiASIs+RXi1uzFG1PioJd2oZ01
Lc+9H0erhtHGQw3cvLUS36Ok1ZFq1Gn4fmzk14nO1Aqyh+gjM7l05tU4q5u1BEnX
NEv9iGIu8pbggCnIIK8CqUwgNe+kdj6yy/YUipy4Euqw3aPQxDDAbygn7a8DlEzJ
pBgx2U3rP0DHJobe9HQIgQ/JmLbBqwWd559OoxsyrIptak5d3sT8kj4B7VKJo+Pi
ivM/qbHjecViXkp/bAYqCd62lE/AQuoBxI7PYnsuKUMVR7LXIEwLDwg7nlZPlUR/
8uOhZXnjOBOIB0uGgh6F1AKrJFxWywet52ZhD3iOaWiSqqAYq+srUg7VCUSD4R1N
`protect END_PROTECTED