-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Op8ijMpdKGeyvArzK48XEXHpplIOgjnTmLLUDRAE6K2z+uOvu+pjy7rOHv1+cwaL
WAbDp+LFFnYv9NXfKPCLKsKVzIVjrOdrxsChIn7U0vBE1hOmbCr84q9s+F6ye++/
s8IK5KIX/BYY+HbhVsrrrYIUK2f/hp5SpWTwc53cCZs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 84722)

`protect DATA_BLOCK
yed4DtG6ELhWMbYmU5Gfy1/y8gbX8LCzqZxXKJOAteh2vP6lGLCMTLlIgt9+oarB
nHRAolr4Twmxm+bQqq/xGTc5DYa/9suWcdIRbn7pVkOTs40uj9CUuWnfyMR1wJaW
OKF9Vi1DRMb966DrRreX0amoJJikH/1JY21wro2BPb1wXFEq+s19ulUQtaWANE/B
46+nr4O808U71WDoM6fxWifXGKS9o4SAn6WV0orh6mmvZ5S7Xh5ZBzEuHXmnTJYi
CLBnzuHUvJ930YqDfmlIGO269E5HZH2ygUgNKK+qknOvoxP0MLmlTedxJOg07dX8
OMTVTTN3uRtzXAxIHVv40ZyR/shOUlsXrmoxYtcZbd1oPRnYpA0COF6jNQpTWIG4
C9EqEta/HlriIiKVbAahGv/X2vFLi3ekuUy+4+J43r09Hpt/rb9OJbYb1k/h8xNY
9OfRBUzMpPM4i1LdFtqNkOForeiPu1bVB17YCpXYV3DMBXMiGZJPTo+Xa6C9Uz9l
F/q1IcTaXzzgCwvbc/z91osXtQIBx7nqA2WXgKfg09HteXPZYiMxea7R8NxdNtQh
whLPz6ztCEe6EMli3VKp+FLczvorEoU7BnCKTYw7USV5WLP6LY4fjOecGQsCFC0c
BlyQz3grZzLAM/tukpupfTkdnltYk6QZNIMFQv7UCF/TrvoRVJoHYDuM0RLepMvj
WwmW5Exo+MhmL6yhEoZVD/4FgTyZNdJF+LRDWrn3E8Vm4xptKBQ1XYojsDwFJro0
UZtd7qs2hQjd3So5S+cs46QIIE31oyYotieN3R8PYJUThO/P5KgqQExPn2b//Yws
8GPbVeaYEOLkaFm6DopDbmyLvCsH8tEZN/45e2RtMjMSVLUw2Yp1NwzEsKmxmlUP
keUsPY1pUaezmXNoBUOv076NzUewfVoLB36a/phZzTM7N9PVW/QHEXVPu82nhEGt
fnDkQgjzVm+/xNddzRetuijxEL+JLmG6dGqaBQWIGOQbqTQCG1hLI7MI9QnGcMgi
y10xBuZvLAIlBauUOFadSkHMa7+7klYp2xn7eNtMPPMkM+2I6x8Z9HxxlrQ+DBtd
N0CbNETN7nggcb8U/q5CvBAvDZ/xMc4jeZy7Hgysbv2K5tnTC18n+lgzGKzDcYRB
jbO0wGfI4GuP3DixEpGY81eYFnENHbB2QlCaVrbLMrlmBQo9Gbwyc2N5sIsHxFXW
eBvmR3OStXXQTWkYsFQTVTif+GYAxhHWLRMR/1Dyw5nx5zxv2aXLejN2YXquQzBs
1ZZefZrkg6T6PH+PLuajHoGml+zDUJqkmaaBuxXdlW/OPnnnAxtEfVOFTCaKBm3o
qaiJHMpl796nKNxiI5K3K6RTW5K5Q0e/AUfS9Bx/ihNv07LRO7E2n+6T/5r0GOW4
VA2+MsoDPqg6t+tuzxqv9mgBVfrznd7EzhA6uLFUyhSmxScqCTucwEpLv06Rb/tr
u+W1rfAHtxfHf2t+TDFK5mudKbOUrrL8ZAI7yPlWuqFVZh34b15YiW2ZyJXZHy5n
CSUooijF/aFSPGbAeCpiNxRBnlF32yJ6HC3iYx3LqDqWQGjlqTlce+T19hne8i7H
teq5qTgfZqed2D43yhLAItx+NWK3KbeHypX64J0kCBtg48HWspqGEEyYF27gDC6u
q0RlGHGBpEwCjyUB9oy/JW8Uhvlacwf58XswoANAAnJIyjMyikITaLAzgW1xReFv
P1+VfkTcV3pKo5Lmf22pEZtvZoaq3SzTz76Y8HnvTfzvPVm6Qv6mOji9gINJX9vj
vcHGT2ZgFDda5/nE4OHRpNdHEBGa3UKPy69bNLbnERQo7gYU5YYgPS1YvqW5Susm
UezXHqevGLsiu+MV6v3tVAkFEVsE8lwtYUMHrcm42B7J+lW7TqR88WAmwPm176MI
HjIsA+aZAzmgQEfN6k0IMfqyUEO2AuTNe/tT/wslNRCXxg7kwIsW3KSv56Xcfjcg
OEtGl0wUvKz+NPFeb2xKw7y753HROud4EQ1y8OoUY1w0U82LWn9rstVN8BrNfroH
ZYSObiZ6tQMnNDa8cnD/Uz+nZHp9IKmZK6QyNFcgKqpa7hscywqz57frmraVqzeZ
43avi2QX09SlkS26QgRhf7u3fMobNviGkzTJ9LwrNy6MKsVk8tEXENUl2HMf742C
HEUR/k668e/zoyObyGOACPNd0i/0pgzk6y3xCZHgZo9eZ4lF/9ES52HcJgvMsMNh
EWaEvPdJNnuzPQDCnzfnOA4Ch/mFIKOvQmzudKvZXwXQFCdW3kcwZLonYFbQ5LBn
lrXwJbTQsYF4pFozM9BlXlrI6VgSp6zxePqXRmNjKmexKzT7Iwqn6JYJvP4Z9gir
ht8Nov5DSKpHWW6WGXSBk953OFDxUWnXiMfcTwXpSG61oHlg/dQL+vG748JEDyaW
bJbh1+OWepm/zBP/ndniBzpTtPW0xPBGb1cvCbgRV8/c+jKrn4GTo2l6xbJyYW/5
XPEoJFAUliVuRbaLB9u3S2w/JBzXwaJgwh0Rm0xpmyPx3EyNjsLDp8xWnBlk4jFU
bowGjmyPQaMyeBW+77tyWaTDNsPvPi02UFhXMamsFbvwT3QUDac1FDRiz20M5kcX
lX5cxeEN0maKphQujTLsamH9sKd6ysaHWAzxluyfqw5R+HB9yf9x/WCxy4j9RDfi
0PFOjL0FCl8GICLckKaix6XcoYpMcRWhwb2hhVG1PqTeP8iLZvzGOxcMaNvkfCYZ
z/LeArTT3U1WNRavNRLY3XUwRJZMcZXvFhB2fMU+nIqsHqM03tx+RdkKPWrmXUTT
b7GHaQHmH1kKbyqHEBnM7+sNxs+2XKoO4PqxEIrnQdLmPec/iS6G0wQ4K0rMpo3E
+mhAHn+rOexmIwfY5CHSvhZT8yV02NjqqzgGKhA4bx+82IcU1qae9jcO2nABw4DS
QNtKPstUMmFKAOQzTa5dMqSIE+YFbWZslKnRNqJ+tudNgR/nZ1gOHXKsQc1cs8T+
lsC8j0YzfbCf/Z+3doM6igFkAWS0d2qz7zaeRJtOQYeiRb/i7Jw15yJYrqlkkU59
dNR1s/9ecx7AJ2KHr4PVBHTUICFa9zIiOhbTaVt4fsyboq8sjslZiLE9dlt1L+Kc
OpF4IA0rkyxldyCOOCwJTJi+Ai6Jnwv/oGBFkE6pDuqKs5IZ9xiT+oGCMfTr8ID4
8VtFtDHfnm7PI6PPyDEYLAvTImWgQRu5si1eI6azLibeQf1Wnd+NjXjcbY5xRvF/
KFWrk8LHTYSStyulhAm2R6hXJExIPCAj7lCjzm+hsZUMWSccRr2jSIgmHS+YMwnQ
wRKvGkIRrM3xMnyJy55x6EBP1ditH3538ScF9IlvRYbgy0PgH2aMJP+BAXbvRZqC
84XZtG+i7Kc5oVGkvrDcuZ9amfJRyCdkUi1n5jks/MJhsO3J6P6C7BcZQyBuKhch
MYZO84Vf8d3ZPzZvnP6y6kp42lw9BzT5RIU57TSe1r+rD8OGaoyAHDYoKDs/rRXo
e018zEMrcfPqzSO/R2IrTbx5GLMMSGVhnRhQBNQOuXttH3yIUDJvGKyAp24jOGnk
5piUDSWVJKKxALNYU1iLqeyZk9zngYUeQ1VkM8QAJT6MTZAWNMFBEX10/pmDb2/2
RflKy8Q8dcJGq4rRazjYLE55v0HOV3E2gD4OA/S7KKF7QhD7lu4XF4IDCzSZ79fH
A5GB7CsldTjTlp/mgoXSWwPqE0/J6q0iiDV2dMdw6pypuvkRq1nLGO9V64E2Hqpp
9X8N35s2KXCTNTjZIkxyYLXGp1hwThcs2s5k8y/ndPexWfIK0faI3RrBWA541J9E
HRydLyr325l7wCEF/55Ng6VTp2n05eaeeXECABIsxBcSGETRV7DQ1TCB4RvcTdSg
h4kyeAGmNNsNl6/F3LbXpz/l/0Q+Mr6tRs3SsblD9ivrn2Rd17H3+rVqZTCGrLuF
M6BX0LsKS9HOaKQpOovPa9gTEmX909gvrQUIXFgFUUR8O+iVNOGRGXif9JB+Q0om
affufmDQMllQkLiMlMC9mzUynqPm/8laHsWCq0081riWmmAzz6kHagnjqcJEL5wh
fMi8BsBHgvOQVwHrG9QTQHSlpUFLbJ1ndX3NqejWp6p0zx84TM7ERLWHUV7qa+MO
lhaj4sMsd02EJySqvIyTkRstDtnZusBPBc1tFhOFJojJ7/fnqoAqtXyQzSN8/d73
nEUyMXI9SnJe4hP2tQ4yni9gSoeEjS8oX1OyrHKVJWg1LOMRhnVXadIDiD5jwgrs
WcG17VmvipTwcV8suia0ztlRQlao5l6q4L3fN5FZgqmgkePovaJ3l0PqB/QeXkL6
B2kyN5SMabx1m/NFT++mHKbakg2ItgeNYuGYAxchlGJMhp6dWDpSK7pC1YMyJx09
IY25oYnOVPwfcWJFmPn5lElwWf/EQcWCMmV5Gz0altF8GERgjdDTU39vN29SiFT7
GE9EuRtciceW4ddP/KK2dqpkmO5kRPYUxQIyU+A0xQJHV2GvKl8luM2UiVesA6pJ
dBo1cSzJYPVMq1fc90CezWWJ2fkEHaLM31WLbAdUTdq6/ZikhKFrzp5wfn23buaO
xn52lbzXAEck2uWxjqFOapyo7/LjvFCuFhJN6HBow2nKPScAjieZLRY9PJTzgQNy
Lel7bybseeuFAPZvPIJiesmap9UjCgz4Lyk3Ct5y4lj9z/lIIkIGyRYTnY8Uu+pX
CeMClv3z7Cc1OCps4H/FQPMASCYFZi0RAz6A12e0hGi2BKz4Vy84H5v4IlC0wNmi
beOUBhXNDx5e5mA9iAwqL4apeILqQwGuylclijMUj1qn2gF0Q2IqLR+nXfRj7Sb8
bMMLzJ52nuOWQrhEg6UoPKLkzonQng7LiZ+PLnedybvDWvDIh7n1GbUP6ETQem3c
qf6UUrWrnApWclu23zlq0g9J/OsAXVQbG4WNna18GnPZkCIBaa4tqmGu91DEp6rV
tdxGnEnV/aXbq3LAFaRs4O637tcrmjpz8YHZPGKQG5e7+Do3tDt7WRNnPbiQ8nFB
QnwhZDxS3POhXXr5PVn4j/tD7qpzZZErlj3bxrAMbt5mJzQyV4dPbpBoMfSJQG32
0CR0dycbXek4ZnBaLlZrIzbPFCnZadsyICdOGHVVwQXHIS50To3mwVDMi1XxH4iI
yG/CNv7RlTBpgoxznyPWyBkupBJiArvuNrb0RPwVB33upbx5tzZADomzjh8ekwUV
0c+yi4/E0+OgF5U5a9SjHvGE4kZ9KRyjtMTboJJG1znZal1vaEsgc3qP0BzXsejN
HSX5FwXSGM3M6PGnsyejRliNu3slLQpcP5DjuLUSlZq2U8f8zX3tELAxQZ9JeppS
mrHoKe2i6K1PUBwXyaSdn/ZFAlux6DnL9YnP4vAvYH3RnwDlMrMKGjIrbpLN9Gg3
zq1KHXMv1AhnU1jz+m8Xq441lNB+xjUC/hfHm6Fdr2QrRr+I2R5IL/SgPoWJoic4
HwpVYDl/QLAhtixDPGxzksCGd7G/jf6EKpsoUjQKOivOLMVw9G5KMCWdsXtrYZqj
PmMUg6czRe9ZQs3nkPeI5swKPdHtLwOEPwsYbFC1Dta0zKxC4joxY3AImuv1BTsf
xR7e+gTfW8hq7SBsA3TjUnzVxKz+gFj+2QQSfBVqcVb2QK5vz5N2QDrw67jEO1rQ
D+qRVk9IH4P52j9Ff75K6V+d1wIt8szr0mS7zXeYJmlf5sUJRIXiXQ0rFgqn/pOS
CbMQQ+BiOUq+Uz3Uy5jSQU9/KTj22G1muDb8aGxb3ADWAF1HAIZ2b9GX+57H6IR7
0neDKP2159NBQiEHv6/2cX24rpjv6rMrlxJlG1Vi0S5m4VMdK6eg5W61L39jGbh9
pm22S4jpSDRUpV+7ZRHg0XVTV8bq6buaA1aaTpEKu3+U+i40x2wt6nsIxlXFe0sA
valj3GQ1OYRhKW+cso4u83j+IeYZSia/sHpTykDEO0Y/FfBy0ibi4JAgiyhg1yb7
ZNrWUgnsYzu0QaUEmGoAhKV3uGzemIbI0kZo6juC6gnPRNXAE4jinarg9v7zMuq4
aH4r5UtsvTAG82yQ7vVFDW9/ld8dCSdzgaM2mNJs+cQF54z5jSYsewB3ituyEzXx
DVsS64g4cOD6TQSdV861SdrzlugkCDkUNKcfXKa7Jm22FmQnOxadflX8YAZJePOq
Sfo0lC7D5V/cmFMO5lbvIm+Qw4ifds9cR2hnv5yG115yB2axm1pAKVVpQJgrvHHF
Pxo65U1MOzN7Jgmfn1H5/joSSY0tRAmuq5FnJyZzkbVYDo4/ofp5F9SFopoaJEVt
vKK2aOEDYBRid3r1DbUiqB9e1QChSGUjScvIj5OKxeWm8nlHcxBPeFG72RSk3GoL
2Pf6iuutfiCrmE9u6rG1YAyAhlyeKmlXvfR1tAZPbAY3hII/4Hg+deLMp/1O+noj
fRSZjH86xkNQ24ObFsWcBpYvuhwM5hasJmPLKXiOoVRI4OIjX0CLjujPzIhYFkXk
EakhUqyAXFqLkbA4ZGx/+AXybV9S6G3e128/f3W2ENfIcSgLaBEbUjZ5ZeypIztQ
YMsbQ5nogjyUEo6eeXKlVWOh1vQ/oU+sYKdbZY0a/yFkmpPpNMUu8nLNE9jawYaf
CPAvlOrUPxUAjuQBz+VY71olLN6tin0mu5bZD60sXBGwJnffF5SFYiV7uAX/9h8G
9J2JM1cyBJLbVFpIAxrDxLmrJuZf6P00znynQDBevKn61SrERnPjqUuprJTlVPq9
67zt+PmNus02wA807lcfQwRUyc/6YFSDCRSAzYNQwauYWEyATADEIeFxBHZMhqjx
lJIwCD2xWYnsZaC502fpAm2v+2paJF5u17zY8RagPsmvGSROIK5RcqvNFxjz/Fnl
vKTYBn6wlbfjQ/c8NW6o1Vu54QPeJvUymYzkcxZ4fAKzc5RAq+8iF+/1Pv0rni9o
12DdAfuOP6b1wSFV0wqJqMOF8VnT7qA3+tMqDydeOTVp9JsHb2BipacLin+9NDyC
YdF3rkSW0njvDZZqPKL4o3dS+HrsiAFIKwXI4BudBS4Ca/riJ4w0N0JRTbRZq4ab
EV3DTnt6iWrfLpw/fUElmsAQiR6ImHzvwoGEM2ReIumhyETd2jDgZ1r3yS4F+lnG
7LiVl/7b0L4b+JlyxyrOj7Sr//MoA80E9jOfRPrV7XIIl46lMYk1Ab5DSe/uzry7
vR0w9oIjKsETSTrx9nlw176900RqePXe/SPvUM8POQkjG3wF1ayUhiLSd6b7rIlH
EVqcsfQ/sBGgKHsercdUGivLXQoBY+WXFe1k/5O3PSoHzsJBGgawQGKKu4vd9Si7
xHWw+witOjHoSTaGUZ8UAh1P+3vPWw0NBHqCFJFW/DZMMSNjoyBUdgZOC/PkjJ3U
gN5VovAIs4rLtKW9l/jIJO94sRvyxsxys3+oamdRSgQrfe4oOKswDZVjaNKw2xKr
mDVisSiwIppmFdDtW8rV2CXVFW/xL0TN5Glmr5LqJBvGibnfrjfe3otbqQS9+T3B
ZgUgNedkc3I8ewcoBtvPYNWuGb3T2Jla+jP3Ybbg76gaaDohSMhF2mw2rTKUK0TK
l3EXxUPxMf9G+f/pEet1YDoB83j+NggrqT1pXTh+aHGYX9HvqKqM1bS1omFet+GT
r597xcJ3G3vJdGxUYGfvEl4Us9bkIIqI/3hLjgL3dbG2EpSmA8id6uvX6NGk8CTh
Ui3ID0RMnBGRQWiZ1b4yBTFIyOxPJlm66n4Dgb+zZSwni683Lx6tVrulQTar4LSI
IvV0SPmtP/WcL1ixY4RXEA8FsPMoaZF1agj8go8TlIlb4Qy8jAF2Q4c2Q2xsIeha
CL3vlPaG/Pu58cweL7J309f0pGJ+OWfl2m8XJ4h1FtZUMi6+NQsKucjhWkIkBQDP
2kQkvafR4ycX0Dcf2aTMW9Oc+0CJfnWoYvmYIcH+wzefuJPl0g9i2HP9mqCVLK4N
Ts7Ly0hngtuUx6QCfIWFxMnFjcx3SeR/Z4+ALvn3WevZ2WaHZ5ooRw8THpxfmK9N
b9zTCaK320OaicwnjbVMBFSBw6czjILnciy+fG5VCSFU+E+pKzWPuZKKKSDtpr1l
yPePoOzZ/qAEzybtxThE/tIAYXGi4YvXn4cUwGC5XWlM/FqObXFuXidpz3cJoBaV
CEW6GBhWuLiM5BobbwecMgD+VCjBF5KQd+ptOMgaJnj2i/Xd5hTjRYmo0UZeYTbY
wtbAd7Bi6+LPqQVWJMmz3OSM7JPu/Wdo1qYAwBtlWefIchoNTWvNppBgbroMHbJk
N5MpdWqLLJaICQ6a0uUxIqQAmyn02HqJzgYPrVirpirgMTkW/5cSGoVN7r//W9uG
jW0/3WnFnxF+3PxDIcMrD60+1/vRl10ZedYLDSucCH05ewYD7MaayG5ySoi6gX9f
FgLaTwXtN3ycy06vs5UqPeJ0T8lcRBVnejPs69qulkpwSlScTLKR4tFT7BfvFUFA
maVMU4MkXss5z+BcmzI/NSeEc20yAJKpDaBx9FzBNNwXu6GRU1kG3A3rYVNyYMcz
ZGHuBWzfsbGNleOfv8bi1ISSwjQovwji81Yd0MPymz/MjER6zE6Qk9jrNNf38hqM
Q5TFsObiWYO1bpWMq/rIvadiRPqnYLqig6KgNcd1cOmJ8rDawpbx81GcwlnSmyCt
rL2cku7Bzx+RqmUKl+Vjle4QCngtaL/dOd7v9ObXpW9XOhtXtb+aGkicwBLkD1kc
Da7Zhc+g2CXEJntmrv00jfS/79e58Jnyg6imksxl4St7rqpqCwwyqymHdfybb1ZP
9hI/2kHzeGhc1HTiz0yu7HJrKi2NVAdQEzwJHiRa4IjUTuNUeRv498gQbJrp0Exu
lqJiW8nha8V7+9oatp1MMIsHpSzRwzQDuWdN3H/lq94Zp6rRTiyA+LvhVOmeNssS
u/Hja/1scHnTGUh8M7NUdcdarVdQcWcaNSqSxNT7D79rnR1Fe5oqW2yOc8f+cXXW
iMFrdXcIdPBOGirMo0IxQttRjxr3FLd6DWIYA8yzuoG2b1XFJYSbUWq6oXGwDOvP
ZEiLGDHMpeaGvvwMhSC7UehKIA3UyCU7bCNDKK8CQxOTspZiUXfKSu70SUeIDO9E
fRSHsP2J1EbR/wD47b/V9y2MQPFEaPY4AbpSjmy0fPmXtKZIKWwfuK8XCjP4uPo3
CCnMMLVV+/EX3K4YvGj0Mr4baWQiSbvLKnIXOU1ioPGT6oTWJj5922abMx12LuME
ibiZyNhC5tCKDChihdCgNAuLcJNBKs2m2vGmf5ey9+HAve4kPSFmG6eGFv5qsZOf
hF9sg+aCLsy/QtPMaYp3pw3ZNAq3p5/Z4yo8S+R26WRzaDRoe2FB9ks68qWCCZZW
DCKAOqmngfF+zymqc/N4lhtzurduvay58XH8CI9PI3e/QMeFlfRDsvAHsIb5kPeh
ekLBRCLqtqGh/Ap8iHjhTJ83PPsQ/WpmivkcMndUbQ+HmCSVbjppW6TZ3ltIiFuR
O3qB42d0sbmfzh/beA2/x4bSgv8FMXkniwyQgdPXlDxZW73+A1CV1V6JWkaBB4oJ
8Ge/jLv2HIuiF3juJF7gwh1HYM49W7junQvKBsdkXKSVdKYKeX2zTO/RbwAep+Zh
f3EBwnvUOu34/UsXz4MrGON3XlGdxlpPF5Eox4guCz6Nn9Z2Le086sZwvapq+LeR
id6RHJeo7/Sz2HzAjiJAv2sn6azxvs6sHqbzBPXuI2kcJnXNUaW1eHbpxyy1TBzm
i6XvmOoeYlKkuDESqpKiI6lyssfbYz3BJ668/Lwtu4ejzLAWX2wwkzWU9KNYcjnj
kYEhkTTHThmLRNxwCY6MjJ4SjlW+MkVltw/bfYt1MS5agCphYBcCcUNDoysLee4P
RAAPvdg6ejyUy6R3l8Ad7IVubbBRnF2L/xTxdiGocE7tY1nrKRcPe6ACkRYN0CjA
14wC6u3b8Nu8vnpm4Z5Z6Qe4MP2ZhApPb2b/nCcCmbCc43A9WCz7pQGx/zyP8t2I
+eRxgd8nWBCU7SlUYxDX1Ssj8ygdlrvoMOqcAm+/7dOMxQDTtyOirkLkrT42mIR2
mkUzS25dbBrwJ77yUbjXTcnZiBFYp6vWCkwS3I5okU8obCHs47/cvRE3oNQmYlcA
UBdrlSkiM7eHq2vrjsePF5F7idunBfu7GmvLo7cSs3kRuols45tf8Fsq6S40wMkq
nH4IWyxlJVM0lRvvOPDqcOOss9tp6RZqpZS+o5FvIGDUythr2iQ+M5AO5bKwL167
K1b//SEm1zCTA8+INe/5OGvU7O3ie/l3BNVay8rfv1nqDJKDOlG2zCqlJgBzBx1Q
bSRAdtKco62Uq94sRGmaLFXTUfMdoEkLF4HjYNXsUfOOgrJBqHB/4YWcx5YdiNS+
N44hW0twyJkJym9H7KRUQgaT2uuYS4rdA47IKebKeXwLOo6kTyXguSJpSAcXeJ/Y
tgI0Ld7ZuNmBp1/WAdb/3j/eRE481YhkAs8yXfCOcb/3kKpF1RS7RGXBKW/I4gQH
B6fq0NRvNQiy6If7yTr0fV8mETa97Xbh2lJzFxRaqHI+rE9twFYcFydcXj8XtqfJ
jnPuBok56tg+RKo2lNLrUIo+E2I0Gt05Y/TeDy/X53ops89pSkNwSHTXgjBqSTyl
aYLAeQWoss6wRG1ROROc0mHxjnqLTmeUiRuF7/QuwDpBhtjNlYU2juQPrUB/ZFvW
qHIwW2jPU0gQlIYdCGaI398pubwW9LK0sQSSKpg/dSWAWsrgg0VUtXH9Hmc+isia
U2rQUnwoK4DhRTXX0h6cpz8i9Yk+qmVviZMxMEoNOhagHovxpbQEnq2AUbIJLrQm
1BNG9k/U9AEI+Nrg1ADlbZ40NXa5b1xMvaJTMac2e82B4FlUY7ZeZ4kvyl/DTmfU
k+edNG6WxYrU5kcYeQ5Zye/nRJfqzpeVqIz+rzhfjuW2L9lTB9Tu4kdjVx0Iea54
z+4trVqVoXQ6hCy5q/PoP7F4Qs58lihzk0OrCLDrHLlp3+5r3BxX99S8b6Nlk5xq
Fet18e6O6y+vHn8KmvI7UchKE9njo1Rt/5+R8ZrL6Gwt0jQzE4xS0jik6hr9w18b
IXaKfVF27y4FxEjxzO1SFQ2WjIvdYe+4AQs597WjdVLhKDMIv4pevO2ANeMuAevs
h3wxT/5uPCUYsp7+TzqjeNBhC+1mhT7kR4ERo6VYBYev6AofU44RZafRrH63rjDW
YyiXIGlpu4c/yyz05KBPv8uyPhm5IUQEq2H3nMoa79zSKuIQpmjQOS4fHcIsKHzy
d0HWpf2L34mLMZ/Z4yOhBZkJeK+sRPpKxA+QUUU5xTZNShdi1w5M954aM+nlyAi1
WhEEPdnDaHgIDuTShvWAoYc5rGnhpG+aNvj2KI+upoZn2N5So2t9GKeKn7sEbUSq
YfqVG/tA2rjM4gu/lHHy5g4xdZDapqqv3O7nQ7QptaoaKW0fnL9YuUEQKsos7PCE
X7a+xbl8BCqwn2dQi+pWc/559xAHwYu2HmiBtrRXi7koe6cl8Lu8aF9MsFZem5kf
b8+Sfey4L1YiKLYS5OXw740bVIFInlizX82q+xY0kl5zerhx4WJCHYlUxFcAkS3o
A/93mQRW0GG05BafUDYdyrQu1jwX4cEMQiIoldOVxlaxE9TFe5QikPKnRiClpHJu
yS4m8+0rmuu00kaTamhjWCK9XR2d71o7GqPs/XS1Tvw7p94mkVSc4D5I1/7WgUay
hSDpSv1uZN2JiR3GTDo/7+yxx1flKLEC+00dL3pMRLS0gvYEIOSnXC3qA6N+Nt4f
lpkhPm19Nrypm0oycmEtaf6+P+UOhs1hAU3Xs+EfYCg3STZWqcB+NeW0XSvc5frk
UDVj0SL/6t2/KPVK8zHZHUSo+pufa77E3UTvXca9fJsh7mFPYYtisuxDZW6XYXyr
PNQhfZzYdjRTQ0tOQygevveCzVhNhHc1bqtI9S2Bnj9dBEegd/eNHKJAkFZVqJeV
miN3K2R4bJc/oB2lyi8KumrKWr+lheCN7591LiH76Vlfr5L3pOWSvmMYoKDHvaDZ
P2HMDZM98l1cqU7z4ld04JrbMT8MfH+wpyDmIqUCVEKw37HkmEqr9+K27Jwrr99Z
/smSOm0XuJE6cIUMDUkGRD20LSWdTH4GeT6sVp4GnRk2CdzGg/4x/z6Hpt1+vj53
ePcC33e6Fph03h/fDtWDuUWiIkDepaZEuHhw+ZlIG3CIFMbfJZ2DCFbAv0HeCUs3
lAW5iSzXTe1r1UQcaGSa3XikEFmri1Ya590YkLv8B2stDMGfrG1hGnuiijsmqknA
2Z3OYHXCfyor4CR7+KMHKOQlNM9OD0wraaPw4wyS1YlQdcjGJpdCUBd8EgEPfqz2
8EvCOm7OrcspmSPmPgQO6PPpY3uFTps+/2bbiBINMIfZRMC2wHgZkcRupHHUvYXc
ZQ1+zBCHv48qp1gN/mBLyqxqFDVyb2ZaMez1mSQNkEgJYkz8gbEDZz7Azaq5pN6O
krkfccHZ0BX319Ta55uzBdwxIqQmXO7Dqp3PeCvCmv5rz8PfEF+BZm2CpeXxdV4h
F8r8tjiDL0DURshNVWsjNIitnyo4Xz8e4BPdTyh+2ebtUprIafVHIiVZpAd4QHSp
QXEMeieN5S0I0yWVpnr9DK36kwm8+0HHaXhIg0LsXKCdrTmmhuo1ojaI/WODBgw3
EUneDXB1SNxyY65hwWHMSsu7EmWV2agwgRJSruuaEfeMLNpsvrdKQLvnnRr1odnh
tyy+564mbk+/VMc/04Vo2YRUWnrHkoqPOqT9BZt34v8FD1YWSZGtfrf8aGWPz+7P
LdqF1hhWL3eRJ070EAXqRYZ0A6djFzATEd8uZ413kkaf0iJaD5KJZtm2tBmucU1Z
i1yizpp527WrakrbFs4erztpfkO24XyRYRRF6NBUDETLcLjQxavEerEAFYr8yzQs
TaV3V5Yn35U/kM2TJutPTFJ8H3I+j1RJqV0lGc1wRyW6kDBTbfPtnW4PPDV4M7MX
tN3MucRsm18gimGPj5FEIX8HjOoYIZdp85aX68RZyb3DwPdY7OesN002Gb/Uqlkt
BgHns9d0pzU/poM0R+C5vNsN4vbN9qVkbsQK9Gi1nbPPkszzJpihzCKWoxqBJhZ8
0K36+aImaol6cVI6DZtLFCtMyp8lpPbAWlUGlM8m6OClrcpyx3VNnthAMtmpgVZ/
ru3xgAluuAVnYMV+o3o3SW7CIeVAmpxJeB10bE+9UylS21jWI7oV+KugCXcTSWxS
jc9Q4/C4HcSfPqUCFrY9xsm+t54x54GfDJp2ngjD9aOGeKuGeu1F3V2+dqkwXevX
bPFdb3S8HhmX5fdlBrVCKDvUABVKPuSE3l8LrEgRH+rEkzPHpBjuAKbt6Txx7vSt
bnMeZVS/EZm+IeDOdRHzsv/C1CHIPEdg7YbbcDdDUDt4KgcmGxin4hAPynG85rDP
lYAMTdzZMeFpVFOeu0NaYNROadsr1EoVRCKB8/ArCrIFUNcmbzDlG5UKLfIZv3WU
mNrFjzQ+w4Lt/J8oNx6v+B4l8YOXgj86mgKCZ9uJ2Qv2ERnHewxrt0AqGuJnvBJS
il7MkjtPi67kpq0eSh5xzMYxSAg6tABYfxq2rR0xCxAIwyuhnCJfYTpZ1176CHGC
KonCQkMaH2i0I1ONmqm2NZPYiewbbcvkuIptmRx9Vu9Zwj3Biz6kPq4miI0cQsqU
TXn9CPXkLLY9uUXTgq5ppBKaxqdzlrb5tc7P7JAXwfgZ2YGY98WNicmtfvehCTOu
QpPlRiFr53zWIBknjhTMuw3BhOAaacbKRqKDFY0Pwp5M5Y5eI7HSnDPTEp/guI4x
XgIzBy7A/TNaF//97MT3l4JkG1lTtJHJcj7+ScZtOBTbjnPhowjpXQ5DYngUT33y
yWsm9hQqXHAE8F0liP5MT16km4ouNpM9/yytjanJ25SPGlwEgu7hqgmmK7+gyWmb
0v6PmwqalxS2y/2E/Q0SxTBhIebiYN357Pgf0UUwAHDoJ2DKo3a6B0ZTeD9sP3nR
17VVqz4lqWrhsgebLzyTN81Phw0j8nnM6M5qdXlnZ4HAr3LnCL2Wav9hC5WMLFB+
OJb8GIsKjb5xDXYD48q5lTqzEPANQoRTmI4Fmm5woTLW5mOSuEVbXpaqgdi17Oyo
pD4rvrA9VEyrBzMGd/c6OvuCBlbxGzXGhDjpCrJQtZuFAlbviFY7wTurHZ+zkqOY
6PaSRMjKsTDFlxcOytbKDt3+Khp1ViiT7rPlXUWoADSedvBDp63/VmA+Fubu9LaR
GhF2tI4HfnL9TIH77gOI4NC4WeyK/dO80X4pUQI4abXb1dDjSiiam6hq1I/V+iMe
Is9au/L1y4iM5Es+Qlx3cQ7uuVc906BRU+pOjgvpMRZufZ5B32kiTXLQftgsxnJC
1Oz5DblMZWAKbKKj1pQF0aoJMyu0nLYP4z1l/aJ+DOK6VYGQCZQefK1DMEn46s2o
bAlBIXi30lyiKLrOUrXKWvjY13aiSWD+z8VkYqQWkuZCsjTsqNPUZVEfhMVPoTEe
Ps1riA+UZ9pdX9Z22OglTxrxYBk8QL1iKd/gazFawy+dUIRsVs6U8832zfeYNdoq
cBSj1QzHziwWK92Y5oc2PrhEOyj/AoUizY+G7KBBjT8/fJOzT6sMQ6AgqVkPOQzU
V3bL5lgVWiccl5GKE2o2fmWHaxhq1aiNeetV9ZWimT6GJo5GI+a7hFkbEAcx782d
qPtC22CbZOYTGQT3KxjmZmbLSeyxvqVs6QCkM8LBrHzX9B8unKx46e90k3mbTFdO
pYy6GSBbDcEJzVJYtj2e9upERXOsao6PZVy/AcaQzy9ok2/vrTEbUE4BWK4oEWjU
iwe29+D72gEF8iXyqopsBH92BdDC9AttY0CNopbS+Tcdil1/JJ3UF2IUDR1gExHX
A+WdigQpGLAAEsawC0gDZDPQ/V4cN2CDXvtEub2pVmPilw24GEtCHT3/uL3Cb1A4
+5/5KQE3aApWAUgM/UUvis7TRv/HUTp+MPzFo6JL0LRrpxXpW1U2gRUAwLjRzqbu
A/Hl5Jeqb9iNb48e9hy8ci4LcTlN1Ms2S/cI16C4r4rMOhfMtuVCltfU8s1NPCtS
6vUTfI7LLPjQm3DOl7fPeIhupdAjX+xqkOho8O2F2kaKXCa1QCTYj7Bj2kX8+dhh
mUKzTmef/PJaMYnUfvR7fjQq+fO0oNgRKtFSAsYss502yMY/d9eeqMjXqFqj4Hkz
/OSnA/CMWEImnb1D7F/R+Q+EbDPwhGOG/edgS9U7s8odu+jy+eWjIEfxoLUq01R8
lzRg6Hg/uFsgmuw5rClX0A7Eg7YNmKPWbQXEkjvodj53LBsYuHk9dVxlghXUwREz
ndH+iaJlDDXCyvzDC2zm6gDJnplhNObHkx9k3ii5QtfScBHFd6w9HDkzCI641g07
tNzLlFlY6eb4X96kH4qFIyd3NT2+J/xLUF9Mlgx1agFKL8v+WmyueqWHxxUuXMBW
9yhSEPERuxpFS9gG0ojssM1WZW22XCPxUvO+fNJfNN2sII2boutGAP0WeOyDfvom
JgmsxLG04VaR7X3s0kS6rHZjlRemK2jKqJb5U8efVxuy8P9oMAdit/SWC3FGaZPV
EQKf4Y9mkNRiXF76iO4zceL6AM210efb9lIio6rrUq4pMuKLYfhZmWwAGddt9ykJ
BqwCp9HKb0VRYZWDWABXZGKV7/Hq9rB34N95Ell+FfnPD/8Ki6LbEXoTcKGcywy9
gIBBvjq28U3GUBsN2wL4X9O2e09zw+PUUxMqHVv9JQFVvUItudiaFF7fjKg8/QYI
ycdT8+Jyh4iX+uWTZxs0AOxHKPHMtypydkV8HrBhj6v3QOHikumD3o2Ns15rb7Nh
LFWsT9cm7TNJs/yvIrYrJsO9cNBtDUWXMqIVmdqgWdGj+VOduH45RKcc3QLd4yXr
Kex2yRY+HCkhN6YFaUrxYronGE/Myk6IlJi0qnLqeb9ZGaHmPyTORZtU8gjTBylo
IfNt7p2vNfGlzbrJqsycNf90WCHmkiyQ2Cwke/dKydHAKlAT8c+rJa0RqQAR4DjP
UaSgXnjGIVayNAmoNoI8ZmUQ57n7DzD9G6Af6J8dvzJN+hxzF42YIO1DedtT4djp
4JiSr5y/XKzGali7NqHjPAdh/ZdOy84sEjwX/w+PWp7sOYDFZ9HOSCJWtI1B8ANK
USt8jRO/Sn+2xwR8L0jG3LZq3huS4P98dkHQe9U0aM0J+lXFidalV8VZgGViIn6D
S1Cnjvv5OAJEeaNAsAcVBXr/mwm/fxrXHMIcWvf5u3sePWOHX9Uh0I4TeEU1jRIw
UWHkrpJnnok/2Ehrt+fzfXXvm4NeT+d1IKmrVs00BJXuVh21d5sX2vY6DPURJXoM
Nvm+d4MAXpL1D9onoX9t+lAGh662m0hU6tJ5Zi0aocBP8DWyyeLabJWbYbK5Oo4P
FSBmMmWgtTgYM96NTtDPyl+ztGqtfRWtJizsHsUUqF9mGAYDSxrUnZ/geTa+NmBI
C5m1ZJ1BUilOxwi6Jz1fXSTkRXWVRjNp/yYhEr9MOR29RPsctgmspz9oUaKodT65
pL7ofwycrcndXOfijj8XyOEpfopkJPNhSbbqvk29tQQ3O2G4R60gC4aaJwHjRCEZ
0HgoAa6ZVuBdAj5d6uA9h+WKGD9if8a0ULiVUOZnf0NbiXuNFV/5rHhd8ynrJbZX
7N0NemVbd65Yths6FIaXT/9fXuyfrLK1RVwJ9iBuhrYkjitARUDUlZq2VhCSiYbE
cEseHte2mxC6pTfF0VYo/KwDYLtFPAAo4DCkcTPD0lpcZSmDyfVWGgG8unAukrW9
CmU8ImOj2ykn1ovRSlPXnyC2ZTqyiT0tNTLAy4iIK1S7eFS5KhoSkbPEQknX9pA1
p3HDAYpuktGXHq+QwXF9My1SXu+7y6bANjXz8BHWXYZeTf/F8K56NGHLvW4U2nOY
jNWY8XDApMe/Npiv99kDxNo4WEP1gBzgx+gAi2pIItSAHEhM1UjDRVms89uMZdH7
6BoscHGa6M77Wmu1EiK1aqWfKzyWnU/OlrTY0dHf0tFLWWvaga/THONXRxn5la4Y
w5PGOlH8gpGkParZEngbiR5z6uZy4qHhRyuHI6eGNEUtjsyXL+hdLZDDRu/uqBZZ
oJ4RUgG5PreltYyc+UuoPZkGiaPOGtdIi9+48oML2yON4xaZq50OkQcJQBvg3UMl
54bghH1iANu2OsJnTsDG6r1ZzeR90DS4JzOPzLAciaZCtFpf192/Li5ti/CPM/7+
nGI+Z/4xrg4LLSsnB27MHmM9Sdwy+m8VclJKmOK6X26u8RFO44pe1IV+EStr6IwA
Eu3PXDZiFGdS9FqhY9WGzVdbB9S3kH4WJK+cM+qiaMQiotoFpDuQzcq6fE1Fup5E
T6fw1R1ZkyMM559JlQXP3MuPD+MeQoo4O+X6g7zZi2FAOcB7njkyqAlnfeAE2+Qm
vGLIVPGUhnXzWLqMe7vJPlLNMUZIgRoL+nU+n+ipO4Ak1rhr8j4QNqslHFKR5t1v
ILBs8DI2aACJL9iHYRLl4l7l/7fEL6wpT5K5mhb12yB8+hbtY8jtHzxpIU54lOHb
4ARlBTm87IrJ7rroaTV4qoafAVocAcOMgZCQoJk+TF8q97gcXYc4ekR8ECgtF0Jl
qOuiAMWfUZc5yCfOjzf/GTWQQLA/gIEYZzNiCYZ7LZKybDwkSZW/D/MtoPQs7kTP
RFQ/E5UdluSYPHFaI/sxhI742YzgBqZPwsUnXGI3WycTvAjGMsPwV+6Ui4GPDT1x
jgA+7ejHPWJLkXsJa+wt+QquHPkEvSDa51XaC8JDsMOQiOq6O6qnFnL2AdAkQaLW
qeDHjed+uzWRiwWvV8gC0vlljVDZgL3U/lpp2gDxp0Pgr/XVfYcJVX7FrxvpF1Fo
tKopLWevrmZOVkVXyNzTrPVTRKHEl4kbZ754tJ1Y0cy8Xtvj0MOFpzSDVTaae8mn
D96Z76mUjbcB7P2+vgVYndGtSh7uAUHU2vl+03oiJSVmU6c+kVFYB2GwM6dcaXho
gaTnRv7EWhuTpSoxVnIs0NTqV8vdMJKIhmfvRWBeE038asLHPPI7gb32Amo/5oio
XFE1dpVP7Uc5CKpjl2q4mxUyVqWideNdL59JvzJFarbqUPqP6AJ3lvnht4DXuH6r
I/sEWvg+KxfVRct8SpMbIMhi8/s7HIvCnblgB1ND++1CP9pRpoj8irihwXEmjlZA
N+Kx/OxOHFTZu1JNaT604en5p1kzjwjCV6Nvq+KJDkRY6Z1ZhRSZjK994JV+0enS
GC+lYMdhgdnD/j7NF0wV/KbBM8dGumr/AzTRRk/VWu0AlaSKCvwGU4rXp0BRyfGE
xt8mMnHa3OV+54QSkHBSeMCL6SNoBXInotQIabcidhSmz3i/GKrciASTvwYFowkQ
MAhIvi3Rrr9lpflc1fmHJc95THUgWw8lU0wF6hoajNgDJ+UyWzeVe3wfpGYWXlPe
F5WKjC2srhkBv8KfZnuzid3/rVMHRxvoGqGM2CYYcCL42EUxZdjlL+FsuQHeVvmw
soastVRBcFy/dv/yR1fYBd0FVkzKX2CgaupOW+BjVmibL06FuykLnrgcApxDrrGN
MH1bUT9pO2ah18x4sjKAqL0G/PWmEEMLET4fZWwJMJzolTs34IyZW7fHFxsBGEla
J8ffV7Wpn6yk8eLS+gx2ccrWYhuCWhc9KziWjgKiNHmb4gMYg3NvzxPXn/0EYkcF
zQgdFflLSLX6p5EvymK+fywp+FvAIkoDoyu1dlgdS24LYxZWhYxQWk61EFEbmQHp
sSP/T2ekOtYJIy+arckVCpKrMKsWyARX5IefCfSEz2fZWOiBI22Ik4aNAjyp7rmY
sHRqd5lViEWNqwcOVAvXqZVDxW5zi+IdcU1EQS0GqNwJtNp/QhSejs2I71vj1EPH
fghPmBzDgXhmPZ/oIP3/nOtHEi+ez9e1MAOV7IZD8bz8skJiOBP9Ld66jfFIMDd+
I7NpEANAxi8J1HF1YdDvoFBPk6ipyWu4YTRHM/TbpIi19ZT372KmSpj++T4bMSEU
Q8IHQH87cWBc9Bnc3yJTVGBZhSXJ3hWk5RlrNVkpLfXJ80ww9KOw9ec3hoN8tr1l
WA0Wxf9/sEe3wmg78fhyoGRaAABrqpBNmyZcYOBU+q3i0f2wL48gmu6jOq0KuIhw
kglOIDe23sFnB1sUymdtIHcuvS/Kg4FT6oNMqWkanvQelBgC/hIlrQDdbqWMLlEP
1qjm3BuA7AujZYKtQtNx73BTEVqoZmYNLbYWDeMfY6WOAu5HOZaR/hZpCp7gx0sx
PgEHaM/hfJOn7y0Kb+hVjyxXZvdU8O+HvnSDeL+ukL3uo6etCSE/EMUNx7HuOvO5
AkREH3MBR70dofEmIM3+BxWT4pVt3xfz711BTbjrrtDFYgtN+dsiKsiEMUfNDCEd
LT+lsao9QlimCCaJWzj7Z4HeU3fGuvg7bMd9V2rrV8AlYxjHw50gscWJRVxw6/Pp
LQPrDusgfTveXpzxFmxUcnNQI95bLoUwFqQVZKI53Doznr3JQ4eov8bHjczLgnaF
ajjn2U3kbEr3dqqUgvsOa7GlyXigfm/EDgZGXhMZ/KKsOUApAMUoeMHHKa7IcNci
Mz/UjrmR/Caqrz+JaI6OgdMdoYs2lxnHmurSaphXgsmkhkGo/Mmnv93Hp+bHbuMr
XCbv4avc8XM8tt8tth9H+UBoxgp8WHI18QCUQuijEUPWR6/IpTUEU5NHad+FHRNg
PSitHsyXX3+VhvZ85/5vJh2sD+OwCg8ZW5WhDOwn3PtW2YkgY4Gtf4o5PT3i+ZuM
8xEc216LNHzk73aBaheqSmtAjmQ1JgLJC/KXLFXMkVCm//RZXfI45adeRZzDcqxG
PFfpY2wi0/rg9OqjDYT1dpX8Ew20dEl5qHkiC8ojNVJPu9W50q4suwbVOTUKDTAI
xlcIxYUKs2/Cv74gW4NwocZr4NDrQQTUusXe5M7KdgQUO+rAsphHN1vw5u7gjipt
tZtUDxU7mFCdqwbFMDK2AY8v/wrhyUB/yw412nhNrqjv6cWwLvyQ13v57PX4NY3g
7z7UJsy3OlAb3dfDBl5LAEm41Zo4f7CcGqLNBvKvHn0evdNX4WwjgxCHu7Ki5LDo
+SOFTjP1EMGz7397lrwzxRSu0Apydy6L+2/o76wvLCE2qBHmeqbVyiA4BQW4uBGz
g3FQItswRqeQjXxgRijEnWSNTf+o+MrqEE9194yD7lET1hPR4OpJPRyBqdhhkJe6
Dc8D76UT+8feRHFwlboZw35OYdLOpk7VSn0qMHcEvOutR5nyq7OKGmEacP2QQ4Sz
CtWo9khh4CHJl14mjHqgrKBa7XtWZzkFjyuISOzlAkGa3BEuXJi63vfLUuS10C+K
y1+8L6O1+RMVpCBHw0YgWNej2MKAuUMGTB9iFf9WOQa3e0NKrj1wWy9uPr56zHZU
reDM4ceUoBUA0HjfuhShWKU8h7K+DGjLHs6EQD+hFeYsK+73mxzWt+RiplLQHDIa
/vsCplHZNbwzofVm6npwt7hVq4JAIOzhOASaovGI1fklu3rI4E+qLAXY3/fSrWBT
a9XvFaTjOenvsIuobi8Z1dfQNwbiAeP0TUT1jx9Fr4mfASrN+NQoqafbUVPVnGvW
yWSL9hRqTlWoPQdyoLuk2Op+hTrhTX43Bwbd4H4PHm50hbg9TM/Dr0mo1v7ybGbG
fP6oZY4HXcGldKhInbtWFJTBBJ2iW6NlsBFc2y+Hf732nWu7hJprr8lGxQJyYVid
87xepwFE+ANXSa4LvQSOhsasB0bQcWrV3RxRYww++/TcwAomeppKWg24qB4tCL+t
fT/ns74WaafH/u7VZYme8xsWqCIHIQVG8EmTOIULabgp/2jXoWyeaqT3RoZ6hRmD
yDzZLUIad6QUE3lCGEjzYWpVCol1RmECw21Dj8XaLm/GglSGRA/BecsKz95z9u0y
oUIBUYZ6dfryVw+5Rqqj3hVArEyMPeceLDlCodvA/1ZQAtXGEpE/rymJm7iDVuXP
0VFs0IvGp2eOBOZ4MYSNW23AuJli9ukmqgKv6V8/2vr8TTR9Zc37ZFE0jQxa05Uj
sUiQLEVPoY0GMWuUeRH+DcElNesSwvb+a1XMnkYVGKB8XDll9lTjWe3GnrHD92k5
IocnCOYqONWyxgAQL5CCVaw/ZKkVGFJV+Ucbzopi/O+Je0q/EpaS7WbRCYu5Zr/f
XsMHoj3H4ToAtAcfHcL+Pl4DUOw4rreuSv87tsjNKK2tpPzFN7CAshfZNPbOOxOZ
oHb4Ows9zM9JPkivP4cPiCiDwLMhFEF5D8Qzv+Mans9AypyYwmebkX8ovoGsTIql
y+qu/+MciCseZ0pzQSdkmQ+DHvPrByQoO9ATdeerrT9IULxSqicMgocbOM1QYjds
8SpgEKJXhSxPxUCkHnxpkrmvq/9lEirxOfSDcKNwzlb5hNojfAh9a43PucxDfhqB
UP6CmxscgYEjG9ihcJMajSkCoyU7ja7iCbQsA7lPxnTVMin9hGjV9FegjSSfjVbY
zvsT9OXQpAu+5wwgMn+4bdyS7DdAz7JX4fY49mCGFTFVdjKPXGceNDPqMmseqtWi
POVLHKIgJWRd9DgexRtyAW9U4lUYancsmViryaggqg7z317ijSG39MbPUtHJ9F9O
3fENUL3XuKgHT6WSQ9dtNlHCSWkTZwJHBQ73HEaPbzIPtJCDOQADW/hYLWyrCuIZ
8awPwYNqpk/uu0GzARjYDYiXmpa3gWBCDsDcLn5FkWtUnrbQ72IhkIQlRxbSfU23
lvypYiqWzY9VQ/bXavxMmWMN8+cT/RZCKjpgK0dCgPBbTbJy8tBnNyZHm/vMImFa
drxs0KKFhuITjzUj3t7iXFimPlkVEfccOYc5oLc3i/SezSFync6K/jW0yaRyKR1s
r+OGcSBVWeo4801bnDOd9EY+FGi6h9Itixkub20jWl9/1NBL8cwqTXlxDMbV6Vyq
HDv8uOGbZHF30sjANfmto3L09nrXD+emEhACcjhfT46uKO/PkBqRwMiPiWVEb5dh
S55tLd8SJWx+iilqG5D58JAKV1vA7OBkLoXR3YNIdHXiev1KclqHpAI/Vubytio6
RxGoo3SCvcvzfCuuIbNoxQgv9yaRsNSvF8+3zxXwuFu1xNQIrsq7cqmFDn8HliSU
NcJm+o2D5hFrp5COGqfr9LDBQfcJVnDmwMTdAOZbopcGUbcFdFnKbtr4p4kPbVkS
YJFzTYLCTzS8Z1zTx6MOxEe1YJxmd6sxv9/m7xWakvcY7wgnUWyAq+aTm/zDsg5W
HYo6AQ07u55QWZKMYnsHlPl0Lh9FKSHgcsdgFHAEHu3jq/J7HBR6JMyBmvgxq+DF
Pr18n01E8uDsO0W5Kv4AOggnjuCtME7B96bGSKKZuCuIiG/qT3Xd6OO5eACa15Er
zSDUVSdVdn0ENwRea8VoZuGtBwZbWvlwkPhxEKZ87+XiKkv4T0fYfx/z86lkYm90
3is0TDflmo1uli7XwFnQC14ffCiHFEfWW0s5wHKXkc1XpDyLcbRmlkVVYxU77Oen
bcHZQFLW2d/mjyOf6JItE9OWuY+iQ2c76ihq0L7hLHvzeY3nEWDMhBsIdCWRRx9P
RipgVLDD2yzsSUUbY6cNUBu5ACregDFKAysXMCqLZ//2eZ6J/xIDCYma6AMlDVpk
+J4/cZQ/ewImHqJwvShTA8KsnbRZrjqOMxalnXI5TinsYUsHvjFxYEKLnGWp02hY
tr5/rThF4y4tpIUqYZX44PDbr0nM12qe4O3zInD/5yJ3+IQ7gXx/Krb+mVmXDGkM
vCQChTD9ftrmj+2+aMPwPkQ5xQK63yyqiGxBMRg9lc3Jnp2XOgXIWSu3ZWcMdlzf
gfVGZWYMdvq2o7M6TGCN2dcKvdEjeoGqH5nM9cfTIKlFUlo73jrbVtxutjExyFv4
WDVCUEoTEaY0UTDNd3R3IXRfRerMGyVu3+9Q5rKSBOrtuLIJ/dxdF1Z4odoj6GYC
YWW/76dvoMDygbamnMSCqGl3CtPG+ucptStkjZ3Q3vWs+8y8HVZ8xfLqI+hQnpm6
/nTTuM0BsEKxHbKg/bNchekkwqA9FGkJRyL8HPclcqBCrLYMyeT7QCY12NM18Xge
9ghs66m1V/gMjaxlWECwsiPxdnl1pPhE2wP/y3d8JktT7WkTjVO5zUj60pPZL2X1
T3KkgZpqPbCEtMgzr50vhkybBn3m4NaFUbTI2oF+02Unj2bP5pPbhDFYIpx3hV6e
sfHK9rNtn6IIGT9/p+X29tAQxPX6jvgeZcsswqrcZPnPwqduu/6Y2KnYqcGxqSOP
cx1ZBtftGuM+aObgT4H18iT+ON40xFZekej0PYvv3Ee5Pr8Oh51xzVSouYGkQscz
6Uzxl7OPaRjNUOK9WwHMDiGC9FDWs0IJ3JeTUqry+0pp8fS0k66ZsKaE3+N4WshX
NCl+EIyAk5kjdNWBCpPf3V1HixKFU2pBbM782n7rhaJiF3XtJXyVC5dQDPqz4OYt
gsQO+Sp2/RbFEBZnM7Wx57xy+ZhkQW5vmgF1Yq7FqAeATTEik2l5uZ6lzzIjBCfw
pqVus9HQpQE1CI024mllPxJ3sPuZPNlRwpXv3OQb1GR4+Ck0Aat4aUa0n+5zXakp
Lwxmp7tzBsQgd/XRT8SUycqmZEZmZSbcDr5QvVL7hB8AmVOJzRfiTimBORDHIc2x
jrseGqjJtS3b8JC14SosbJ7L3dUK1h30/PkArCv/aNrqnZQMHeWDMPf68pmSHhjc
smFcfdOVcEgE4CpZkOij7b/5VlBS2GVhLTay1c1yDFhG0cqw+yhZ/6kboq+XtURn
YLwhBnZNm1+k/dgqqA3+QcPZ8ry5zIBYmRMMWseBHYAdSfmUm8FmWqu+iS5b3fre
ApQVpzVDuJMTb8B4FqlUlJCBDyBwc+Q/GzFZeQ/Sp48A0GWn0tBw/4e+dT4QQBVQ
A3jfGfyI2UQYIJzcVzf8VI48yzHqbB/KbwSqkTyo8tpTnLaHe8cs4jCMESTFhfb4
z5mEaFpjcy6htKuATtET/eoFXXlAHSmLzXpZZmlvV6z0iSkZE1lghtdR6KyM1iNf
36KrFdY+lnqbaXxYzxd+faHR/i7brsesROx95daMA/eT9RrvQKqq2iX0TIDPQ5PE
x2iXVHZJxWARQxd8SWHFH77T6uTgPyI2X47qbYSY55Xc1bdS/D2I9zP7ELt/c5n7
fH7FVk/u09sgfptl0QWlpZOwTKNSl0V4m8rj6VD5E5Qb5A7MGEPJcIiLYDhTPJu8
l/9bGytxeHWvn09sU8byyytp5CNUMUMDYNuJIWL1NqqsKHApHsdhJ4C0yMgsAUoh
A9nVQ0T+4THjdnq2AbZQxjOVIxm8VTHOAh9OEx5Gu24ZChRGnse/TXz3piBc6KlP
WHB/4WTAFqAmNyAJ57vJLz53eOFAlBjHd5nUxBnJLeCJb+mCM2qR0/CZz+Z6ynnQ
sgleV2HzA8UQqkit2ABkBFo03Yds54u6eIQ0VofIJ3DCkeDbNWmqTQxhfVNYkG34
ZqKaUnsBNO148Qg2BT6gptro7IMK9wUq1eZqm8IQ4Ol+BRGtzY7WDRwMJ94PaHgd
WU9FvLdPrIg0bVrg05e0jiSKFpTS844+1dZLaJL88xPhmo2Hh+7ScwFHdFvjcUai
OZemFlCuRuA2KdHeVHY/COWkd22UVXrZWtkMfFfy2fO+YFeMSd8WXNXGPY9iPQfV
jsPrBbIxvJl6n7mES3q7dYTlIiLjbxkAgj1ot/n2qmnO/4n709hIe3Uhzqar9OCz
RbySynhJzjWSrha+NqHMFbOdizvMOm0xTjNrcGBCFfSAoXzYWU5TLxnz08MaykT2
w30e3dNlGmHBdHr4RwHUEy3sIvVADetzr4tDYS+puw2VIs/MEBDpAL8Y91KeEyi2
IRj7WO3iNERrWyq+CHw5qhtt0U4L87bGDAs9Rii30oEVlTcNs2Hqzx1gqD7BH9in
S7ytLzlEql1ssVInk7/nyQbpk/DWar6s3ZMG9+TbsHaAM5hiRbFRGhLUG/ukDj2G
il1/w9L38GThgTVoCGeXFQL6tzGmUEjTDhP8csAVr7O9Ln86ist3KJHgeMbbUlGg
BFNI6fLKAbJ5Dqkl35m7jBKz9EvzdeIkoS5xO0QjS0f7Uiki2/tl1LF22KdOvODz
n15qNOWh1FswXkPvtUnlHWXFR2Vruk7gipLVqwNQA+38h9NR0mMsLB1LXicnlQku
PUHiMOvOqQX9srBh6RgWWJ6zrv7nYBrkeIsmEsUmsa4BFUHfYdu9Mp1WHruhNR/t
M+0SnNGws9EMAZC164RdtivvbPNJiK0BgzYep+ZlB3J/VQnrtVBLObjNiV0L12fL
6YWG8e8YUoAAmqmd3I2HeU8ODb4mhOAVJ8Moy+xz4iTh/Nu5KMU7TQIa1kvHm3TK
GKXstFrJSwapIafet06zWInbRX7aLl+Vd2drzleQF/p4ws+r+rryF8MP5cmNFfdi
cTGZGHHrLaRXnBsWDg4BMFC2A2bZJfE4vz1mZvG/OgjwMylh7r2Nk1znnBfvTeUC
MhtEG1YMa+AKennI8Pc7gSEiW1eXPMaRnap0Z5ROAFdFQInG6kXb4J6hl2PcV2zo
VPHV6rSSkBTaRVUlqttyE0+bT6FU+Y1XNr/9TJY7VG8RTMmeZl3S0mbiFvC7sBwB
y0aECDjWI+uMeVYkC0be2N/ZmgoZEQmT8yAKrZYjXE4U8IB3CSY0VcXZuTcsSazq
WlecWDQcw97E34Oik9ryDt8VCvSCMpagsP7hhHQRQruSGX0VBrEnV8zdh0atTB+/
jb0f42+IyjzEwWLylFyaROtUB3ITRtLLJmXqOC2W1D2xQuwWyzWECviubfTYSVjo
Tx18gW+Ft5k5AsS04dfB4HCRScbCrRh7p4s1FWJ3iHYZ0yAi42JR03uFk2FLwVcJ
UQZO8lKZyprmfYj7loj9qsROgvmFMxeWbGMuhQl8OEIVA8o/HY5eWLj0frTQn1C2
/a76/eNLQPIbtHlSzXkuauImYr3gTfH/aobLTot5J9ay96O9gi+MZuLmZmN/9HoQ
Li0audKoEQxn16uK2dAvmEBldK/YqA9IcA7Wfwu+ka/nU510Alq+p9sqBJ0SP3/C
9z/t+K2b0MaLBFstzmeQp0IZyv6vcKESV66g8y/wy8fts3BaPOvKi4WjAyMiKEyN
K+7td10YUVAozYYSh6J2+0IBCEI01nNBnQSd301r2czibmWKacmSwt4ZM3bbRZRx
MjiZMq6iDLhH8IklX8d8l/EFNtmDGEIm/L/TyCxyRQOyXaFvaaYXDOFLTEV+KCCr
enG3CfJkugYtjnvtAgN46vk/O78ESaSxIbPKybZDc+P3N526cCflrb5XPRrBiOrn
NbRA3JI8IHWjFaTmEWm7sMOWd/fh3BJGrMlYVdqkAYt1c6jOphTyXNbJZ9cF0OMp
iKBYNM5E4SYVr33WGm4ZAl1/snv/eocY4k1cvSozqn3juBdpHXLnIrAJNydFk+Lz
hd0Px5Y/LmPSVd0+7BNMchD9lOOjIYriX/3H9IX89hBDv9kJ3nbp24iA4rrf70Zh
olRNGwQLvIK0IlLtum/oVsvsKAe50sPJbVP9v/RTvKi4WcKhZKc7Fz3gE0rXhZIY
OrruxX/gwnptkJNCD6JdqakufDJZipXd96mG+/c13zKEafqssvZxi0IX8KvQuKA9
da+WGfvtglrb88gw48Gf3JfSIO1STa8H+lwx8JAHWiqzbJC1f0FMlNjyJ37NVAAG
oN+2YrCu6gec9CZS2EaUFO1XGT3Oz2OBOqK4+4QWjJiwbVJm0Tj4M+sB4HbVuBE0
TOiKlU6FsP53RWdjeenV1b85ZOyjJXOhgsGdTXs2Lfg0WGfJzJhntqkt7qz+u7iL
OIeHTC2swGpLz5/blxozc2ol7+53LwMt0zGKMbtzinWhLgsOYVGvj01pYSSlwc0K
zCd4bJZIpSBvop8KIpPYsrd1uH7/3Kt0UcLzdPjQvUdR4Q/Whqg0nh7InxNC/nI6
LLKIMkkd/4Tcx6hO6U9d/m2uZ0rRKxdzbs/qlUOjBz7gNrVGpvY8UOTWNdPv+Oag
UXAHUisXq2nOVCGaoRRYn08fjt9pFUzLVPkueKHicx5KESJg1iDFVdsA56R2/9Dz
re/b8LPmYYAA4vtkydRk8HsFFU3kFA9d7bnKdRqEnDgiROmMpIazoTO55sUFVEtJ
Ro9ut4U/ckxlhlu0a9IBfxOe5g71z6yRJFWLYqTZRO1SKjQo+uGDqAbR89YGoppX
9RxNTFyD59q74Hkr32VTf5dqypqszPujnd1PNROerzuiwqpCyCgfGYMnvYGJ4bTQ
2uIy5roZYHW5+nzSHW0k2AQtD8QP0hOdjPMfV35/VYrEVbzWOoyro4SbDsZh9p5D
ZMdK8wF1IVjCL0FaEK1cBE67l10D/oXPBdqCUW8XqmG8n8bqjzO9cXTclDTJboBc
y6y8xG1fWIICWl96fB3GOYitGhywJqUM+CFd08/503+q3AAYMuB9WzTUZibD1FYw
AJfoiRveHjmUhvq/tVEOecJWgooEhi42WaWYHTLkA6INOPqmWGEQW5mjerokTkex
iYiMztbhd9kSlOVsMYhR6AyPWaDuhuogj0R1wsJi9d/JHAFCtsdhbrWrz29iR5xv
0u9f01eeQm9jXYNTsMxc1oqFdWDUprMVK5Qcw9CDUlrTkm8pVvceyUDIws6FPo3o
SzGdu8LQNaQ4JTg3VHQf/oVLMwTlYQSx6ZGZek4cUSEpb+QTCrBVkDZYWl8kRdeN
XcpjgD1yJ7ST6z8+iL1P2/vJ4Ai9Z7eV6st6xSAsJZJgwSFZlKWAQtB/ovjQUu5E
ldqkCEaci0PSgnW72xNvrC/ZjhXqkE5OzXYuoDTtARS2ZTx2ybq/1OcQXj8Rgxyo
Yh0WoSfloIK8P1V+Nohlo6quv8Q9gYkI4FtykUGSsMwDMtl5ayxVKup6GqcdaFGg
JPuLhm7x2rw5gmkIs8/iKXUevez/P8TN5KmvgKlSltKCwiW206FtTmUf/ru4WFC2
MskWwYReCyKvHvAY4hYr4t8qoO69Gciy3Cwai/6rV9+Ujbuct0rqTo9+D1ptgau1
3bfagxCtoikr8o/qyNU1lcwaou4oYRGa6PBvsO7QjkqHOEjDmmZ1KwiJb8hzDMjv
ilL09V/WRcBFct4k5aspQcWW1KCFSSwiawgixQvsOJakJ34jWVJAc0wlrN6Tz5c+
fYlNgq0jkC7R4NCz+99/tp5fyrccVdC/livw8TUb1U8AjRGgQd/CBMH7wv/5wWqG
ETm0+6ap6Gr99Hto8F02yfOywtmsEokF8GTM0swJneDTF9MCBadsIY21YFp54Pjg
ITNwEUm9c6iJbls1Yr1thEu/Pk4NR4jaFK2sXdu5PvYR3ynrvBC7SxhUKnMfZgYc
Vzwt1HrSXooxNlhjh3p5yhMYLAEE+Pzbr2Kjkrr7ICWdeSfexhCE0Ma7fWkxqxjH
Th4MGORSpQzIp9heGvZrvQoqFF7tOniuol5vaRHR1e9vl49W+vH/uPVxH042/N+K
RysJQ7RjRSvahoHQu98AGdddmQjyscZu4/rz4DnVlwUfYdsCJOndnnrqvwzGOHPr
dlVcJHMNvtuvRFcBFPFZhLtRF3pi8kjeFXRGScwUmE3VEuiZE7i94Zdm9z1NoCm3
4gIt17RMJ0J5+ZYgwQ5MwJXPXR9ttzcjipCHudqpTxzIrU4zCKy45UEuw8fkwKge
N2BhWTbOnGL/KwgS7/3VEIGbV31irFYxfnBluCtFxJdLCxyCbX/558wE4mumeUTT
6tet3a3bPaQ76rMIQ9elLLt1V5ZD6f/KrZ/Femfo7JU4P0U1O8FuVce9/XAYw8rN
IvCQZiMMVczj07UXYUtMRs2PbjbesaFi2s9hebZoF3S7f3yK2jK/Xvzp3mLJIkpx
q8la8RB2LkxBR+toGg/RF5s0gRdjNAJMnKZ2ZIMRGij2wmzgsPd+AWbCQKO1nfSY
aLK+9CiEu0J4560vZ6ruHu8SmTpAyeGJjBibfWMkfQssGVa+fxBAmSoxVXHnmV37
/Upd/+fjW1YUMWabqAvkYSZviWWW2VfKxGMWfqUEDQTZHQg8lKSOeeWsMjuayIdR
1tNHJrdLD78Gsv0IO/WNod1b3rKrxIrfLl5xf4PVuVNRZoOqMkl7av0XuskgK6JJ
XDKpnnMjCMOt/y8UINkSXXrPXliujpYPKwgl6KGhThYUjN5SqD5QO+OAjyPS4VYj
7g3YYTBQ8eM0Du8+11hVRu0hsC7Gv8OtbPxy71MuJ7F3DHuLHYDTehh9txUarYXq
+V6deFPoSfNsHNZ5BvDE8F9OBk7tE6MhKHDzUTfv2feCPLsApara6p5yWsliq1BP
6CBNZEpaHITxJcAePqBLe+lT+KNDae2zCizLwifwfGhztY5ajEV9i377k8em6ams
iKLu15OtLFEyJGeG31oUQYvRZoasS34DxIEytJl5rIJQDRZh38v/aqAtO4st5Q39
XH+fet+BXnL1QcEFZWv1ZbiR0gvjB4IzdZiQCXrfEDhAaqki0b+EOTFHAa7yCgmU
18+AzMhvTE/wez71/OkBPVhiDQo+fFC4NiniVywMcPGYZ+cecwTltOTyBh4sDoYC
8d8OhdYJG9By6jFsyk7oP+me6x8/41t6CF50U+B8OT1BgmAEwY4HTvfqIjhMHyDQ
wySQoV9o5Y87tAdAXFJo5hr++F1DWP1GJteTVyRsuv9c3+1fUBnLZG/we21C6vBb
ahSmM+qIm48jf95OA4i3RLV0eYPSjS94sh1K01EOAC+kKKeCLbhGRomtOlIk/TZE
GmQ+h04n31mAjByBQKuUAdtf1WXwoYxZW4cfhswttCPQhYuKLUTTZAu8RyJ4/2qY
iwK2dYS0XGWhuuK8Tot0pCEcqgp/kYrHChAZOh6RjgMXAUjz11wCY9slyXXRZyA1
K6ednsLGF9TztF5+31SCtIctj5yHec88UOc5zMbW/wLq1SLUEBTjys39TYT8rHO7
Lv6yoefBeB/6qq2faiNgHLx3ik97rAH9J4E4NdVEiWbzfGcbKDP1uWx58ddD0+7h
mYZXj9eebX1sTipQwJkPUgaN0V/ZtzQS8JEsfBZN+p/w/RB+ef6cdKfvXJOOKffE
FN1Xw6NQWN60g5UkjL0BXKlp8Z7o91zRBDpgRTDHbSY52bRPNI2Kdu1Rksx54kQT
L5TixJ/pTuud+fRW+nUonPbP9Xdtdu6mQDPIIbjNbpXEEGMJyiusJajcS9SKeU6Q
zQpgDAXZgI5UioeJmZLb/kzO9fWMF+d6+7h6hA1pEbXNPkb3M7Xu2RUB8R9ckCJR
mlAtWG5XLV3rnBKU4LiZvtURnxUvXSMG90g8eL3P1E/GDLs9nOWylEaOgpmToU5z
CIiluKLTpbMHr8otCUyj2c8PK7xtjgu40Vwc4Sytia6V9rHh90+CDzuIHSwE3E2T
Lf7iOgHszSxiwtkxFtreaizGxcpTZvQcFXoAxyb5UaQm9j1Txufpda5D0MMOrlw5
t/HPdcypNJOTxB/Vo6DHq3mA06l2/nNblDih5s2FEw/mICz8bmLjMd0MxMpESS+Y
yZDstIFG9MsL8f6HMmgHSApls3b1OEU7KTiBSY37jC9FGxfzQGVNcsA0pWjMujtP
GvIuVbqf1uoOUIpRcQTJSCZaXiTlJVlsyEdqfZvcXHtTEyG64dV5C0p+oopsovQB
oVo4GPDLvTbklGI7z2blqarbmmpltsQVBqTG2mvG3t5g2SHmIEHrCWxZvfJuwDp7
HblmD2zYvMxBt3XJvxlZd3WGEu+ctjOFTjA5N0XnjFreWQcAdgMjQVvRMiBlK6+5
6dxIJXuAFQeCkRjQkOwC85z5itYUhR78yYCwX6z7BRZU3iJTetQ5MuYAb4bfI/6P
QZGKJDNkhWagCRH3e8xXyYioyqn6DKhc/eerCsL1xt88T+IC+xu/6XaJylXJOqaP
Fe2ZfHkKTT83fMFANHR1fha/XBxCdkOkgEN275bp10hHjhzeb4M0KaSMXlQPl+Q2
7kj6iaVCcL6N2KKq3gIkIYvYRK+BuokxGq3YwvoeQ+mPEe6Ujkg9yAgstZvWyMSZ
0oB2sJqwCWvzrpOryz3xP0qa12R52Sqb1fYMuzVlPGi5kUmvmLDuvm4vmZsRq4NI
X+e7bzcp19OTnS5vMEPQKrcpBeZJAsrcWNIK4LWq/lPuL/Op5IbJrCWDTUeQT3PJ
vFQFfZE3HDB2RQ9vSoVxsFCIaTV7Na8eFvzPQIlRyVbuy4BK1un9GC9TkGlpRpvh
sQB7KBHcM0gRqnREvd4Np6Y9kCdojXc/x0HE8M0jBetRac49PLAzatwbRopqo+jD
HWgkdpNa+I0U0eS3kECSJSeD2DL6ekmiQ9H2JbHlSDwxkRtqI5YlLIbcp/LUzDLR
kwbKR0JffeepeNpMysK58uCZm8I1YIqKjpNbYgaQeICrmh8yzQKFxSjVHbFbj0+k
l86JtxAzv93dppSZMpWLR6Ht/rOjMmRm4BSb+Vr5uHHA545jaqzKOI5ByLi1lcbH
ETGusa5SFvcI3QTnhblVee3cNqx0wiBfB1snOz6rdatGxRyXsE5PeWO/SENN/C0n
rIN2G7dggBDLvQ3eTpXsHCWy1i2sHoDMNJwhDf6lbEXltIcMP6U2+ItL9YSoSou1
uyVE3OYL1Sc7bb0N6Q/9i1PQXywXbUIGPbvqN0AgzpnwFWWcpiPnzj18/jHjtTKt
OTmIRMhorQpmGzKmcNqXWemeApaI+QL6s4xQb/WfXtM6W+O1fMZDufU6C3Y5Fia6
m5KUpeAUjLlFQsWsB8oBQDhkxqRhzPChKb+S6LKuPtdWOqimqSw4Jn+IpGvszl6J
eHnqMQViJwABXRpj8Ws8zHaNtUmRfSSJmirG7EqSueuISXc+AvPa680Rd5gsc6Pv
5IjSshNJGb47slwru6aWbuxhVUWlkXQBUNW+J7pu+zdIUefHPY+Hqcy94LfzvLGe
ktLRDqWyjbVJIPpPK8nLicx17BC1O4+9HBaZEceZ1a+KFNh4tYpwwPShvyNYav3J
IaNviMHWbC9xoPixqlhFDCNTV5atiUcN1SmJwA211m+sRS+PeEMHi8CRoIRD2fD/
BEbcSKFFe5Gb+OjobUCSOkZdufNKqK+kRTEfFq9V5P2+jQDjE3v4HdWvLOpx4DPy
bmLCpJptS7kyNbSF1FycnEna4Tpt8wpeaIT6WD7I9rmLwBV0umIBXcbcJLhVt97S
QtaLbpHUVPn4c+OzzZS/djmF20OfTHN7TwIGKdKdn02SSdCZMi+ivnQid3N+heX/
+yFkv1aCd6Qf2SOzMIHlWxQRryAfLJhPRImoPGWHAiPdWuCNm3O2uMJT0LEWJI7+
gaV4FDU7043BQCiO+ZCoh6Fetu2BvVQb/QaHLP1XpvIslU6SPCkfk/xrSBUeBqGL
dWuD6fO9pAc0d1VoQzZY1t5Oaisk0/M9/56v0byIsNQ2xc5Z7EheFryZHeCGf8f5
SsLzaR4WHry/EyBdZTJH+B4YcYXw8YRQHtT5LFc8FyfOByidSADWE0FzLzmJsfz9
VWx4gPWzshOMHmEqJMNZJUaElC1BgxChkqnAbpZriOrZmf2AVhOrGKiVKKxTkOSU
btCJS7+FBTaxGuHLwaUoeC5QXvHqpor9AdLU7HrJR8prf90EWB+41E071O2AyexJ
W1JsCNNSsVncB/UUCd3478wE/U6wpwwb5Sf2riG+0ZV+tDT9lPPLWtfiBdJLRNgk
wB8EuYcu2kWcZvGrtuS5BtDtuzdFnFCUy+sqaTJnGyLmmc996/Edj8qcZbBmpIRs
hcYdGIdRwJtWUt5Ja2SrJzqC8lKK+cFhDEi4+55PNzosxVPYuAvzoHNes4jS8zEL
43dsadyoHTAmA0Dvb8F4u7DrX3c9nMINKzERRMyiACIVGCjCh8n/Etbq93vpHcNX
A08M2fDfE5mkZVYWWeQnnjg9H6tloW2qFfgCFogek5MAElYPmOytypUxEYRpKxHt
27tCdHuVBQbVpKRendeJd+8ZRRuhtHtYjRtq2Wnrm3dhtVg9SgSF9SG/kA2eJZ97
pgz0inoZLeT4wGJWVfUZQiDGbp4dwWQY4vf6J7i7wK/4YX2W16NX5TAfEYDVLPrX
6lz3X2bLy7+hu4lzGNI3M8LK8WcjK67Kz9gvkN+Cfb6inKNKimFopdiZOioEtune
vDrUDJsOWoxAsZnNM0QRa8vuGxM7AZ6wDXztTLJoqFxk5KPiklCxUjYuwxFr/Vd0
S8tT2PLMgMLFTZys4KR7PpOjQRlUQn8f0zIROWoNu6TcfOoUY+wUjVMkPHn+xJoD
MplpnP02pDuZKfBMD/wbqEX5M/Nhy9o55/pz0hJxpMyW8QP0NC8KaZE3DYhS7g59
QQOqfrEm6RffK4+YWSOlBnPu9FRvNffovlW7X/nqvPs5yZz9kRaaz9geDmGG5Qp0
AE7KrYd6d9tGWdSQW/tUc4bt6WJVM4VkOGPzmNJvhOaIYuOOkF79RQLhFobmcsr/
XL6uBIfHHkoZ2GD0DqRGKdyXmzBFyk8sMwRk6K3meCoPJ0WwSyIFCmxbqrQrS4Yp
GvQvfjf5YuII/g52o2z3S4zg4PAf0VCqX+dR1DaNFntU2Gyx1ToiQarTR+dN6RaE
2vvWG6gnHDXyPDtWCKH2Ibigx0GzYcsvuAfQcOlSpJCqVGaDPajxzVbzjAf06pf3
h2FxbMFaBXBxGQ24Ff6TK2LIOqUdYB5D7DrZFCr+cGb5kiTTBKxveTpvsaQps73n
0N7+CaFSr9WvnVCYH2Iqwj72LhtrHWuyvjevMcKmrTv6ryv6ZUpTZWe3RBMXlt0a
cn458uPUKXS8a4X3GnQcKCDpT73omgUIwdc90mqwkk48HlAXIz4FgaLx7EAfz/jJ
kFUAJC9tNwbb/iyF1DYav+FkosPUJHffimko/zns5qPupOfQ/HzpVEzycyYLa2Bf
5LhRjw94Pui8nS/BzDDTneoUcwhi6DB1X7P6D27E34UgyVHl328JPxfVnP/q831k
XqK87VOEH9U6cU2F/WGCmHSRfLGey3p6AWPb4A4TttiFq/gr4V4H+Lazi//s7Krr
UUUsKGewkxqIrfPMvRlH7qP2/3kUmMovF7RA9GXrUx66du9Zk4kupkvUcn9em6kW
H+F9uy5jakYNVX+1x5AIkP2760MMfuzCx8uwzFE+a4qZFPeLfI79JxZsDmSIM+D1
JQX6acgPPeIMvsJy8f+1aou4l/w4nr+lno/t3n5f47Z3bjJUgrtMgpF6eTgtlAkN
qYWqOlcG10z9/kzuSFvfNeugavePhoSp3j+8Lw51zspIYlCPQecRzxHwH5LXpZxr
f3MUJo6O1wJ2eTX4Ifr9zCjwE7KU8CwHOv41w7DPokWdxfnbVc4WQcvgvRRhPKN7
oNwqXRnZKDTeOah/uHs+gTW9W6+jIlbMZUfdMo58hyno74/mQ0NxNGmOQJvDF/N0
OefDWBSVG/8gWY1aYXjdu8DKP8ZB2ywTQkLpRFNuzZI1uYIjj+Gt3nLPrW6c8oBm
2vG+h4eFft8nQI5ax4wO9v8SrLCzmw39Et7E5NNMhqFnNXaf2ZSE/HjodgjQC0ll
5oh8xNFRZHBBaO73h1tKrA6/SmJ1/YVkN99DvDAxHInF5qLLdwuEQpb+4OJq0Csv
kldtGByEByM4ACgisVkdqvKOEljzbZ215MqQzE90+/bBHN6JtibIKvokYMoCn6ea
cLmwQGsmVaixl6+m720VZCoC7WncjH7cKsoxzIBCm1mcn05vXtktwNYO4o+zmnBC
B+vcN8sxxiawqO/wVY+QFKmiDmOgeAqfU/e5ovnDMehIqWV3CvxuQv7PTncVM1SA
7h3iLKugZuxS6uhe+IoOE3r/4KxgQzt0a8eRfMqNRU9N2YZzDO6i79wkMEvkjpBj
cXqPZ//sYrF90pwdmM7b86sjgwBtykHLAup6KlgqHubAZOAl+EKnf4gfXKWAVTdt
RGj0jkNL4PvGMaXPYkakqwla7118+IEdzX+hPDVrdZIc8O1t47e3vquTN3yx/QDr
HUJ0MrMOADUU6iUIvRj5IHo1/WBTT2RtCqM/R276pIVZf69nQ13m9Fi14BCMlCtd
bX8nw+uoCnXl7olEec2z5Xz+kpNtqyE5skzTsw0+y6jP4BWFAXqWXmEg4uzuvD+G
2dvbLNEmziOL+PBTxO3oUzXq1TVOhiYWdfgke1bobDfDU6SALWHrSW/fw9rRoNUt
kl7csJI1hnojHmW8nhe4DCw9pMwHkmKW9jD2l7K4Qk4kssmrqMOcDO56LQtH8Mpy
Y7Baoc/5jKdQHANwj0FeWgKKykesAyAW1qvLcvnXKIqkc0DH8PHRgHWtlFB4f/Cp
7vvqJ7DBSIwEmVxpP5KDnoVZMksruUKZ+ytdH/WDjVo0Md29UPo/vmKi9Qn2J2YC
i2edi6jHATlnCyHUiyWzQkfz7GQqF3qOV5g1PUWEVdt8JG+pBO8Ryh9LJBMh9780
szONWvBCmD6rPdDd9frWHdMqqaEOrLdT3paeJDySx2X75pyFrRDNApFXrwh/YeZD
EGF8W1VxtzKdjZbJvqfIy3UAsyH45+qYOGUBwEs7VkQS0pmzjD5WDapVzolWAMS3
eoPv/wnQT9wvn7tW3IwXwF5yKQ02b6Zfyj8sCK9UViHwy6zd9J5l/40r8Lqdmuan
ysVjpVV7ZNymIvOP/4ujLRXnFwVJrocmmO+JaNLD/y3QlLYMlAK895uIuGiL6Nmu
jztVEO0JBWajebd634cEXgq6aBU5xA2AULg1YgcdOtKtfVsWqIwSqoueHiXZ/CbE
yQGbnG+3/UlmmUgrdfRjefBBE8z1AElXJQmqpnkdPyBaZh4Nh5hrbm97ygNUUbJy
eKdktZcWoq7UthSh0VmByPl6Mme8Sr4iwIzDVxS//RPbKio7EEeA+xfSn0NPvohm
nqLE7aSrJLi8ZrDmLilgW4/FO237YLm01vQks+3qtGXP5fCftUh10MNlRRmOvn+d
R3emMNweBCchf7XYbVCW2RUxog3Edl5fAlBKNFZ0Dvx+Wg9zUx0xsAn15O+qR0AE
Gq+kyaJE+V7pXmYdHUVz8Blqi01S/i9jpEWoQRzIcPiSwMw8fNwAE4p7oZxskOTh
Wbh2juu1uxPL5oxznT61oYaIXe9k8bCZ3A4InQj+t2jCDp33R4U0TWmK01nEVnkh
kJudWVjvQ7OPVA4VQjmKmqf+tfnJVKJaJob3hU3TARnHGNKv+ecEEpS+mF7tQqUf
UNB3MuFuq/+M4+FKC6ehFkFaTBDpiYi+DefBCnXbT3SwMJfczqau7fjoWrRJlH8N
dB4GVCHjimKF6keHg23sf1LcNlSgWwAXs9C1IoQTKDlivytYC99M6yh6DFjdolSk
I5EBiv6bN0RjXyh2cCApX2h6/SfnSZuc1VtP6tgtp3PbczpuYI8vN6+ehFrjzVND
PwPAYpA3j5XN3JYTv1kzAtIx2Np56zZ2dhLVH/ba905+k1N+dygOq3sn5wckRyy0
43kf2JLbH3agFuixnndI0fBQdNVu5NnyiSgtc2U5evlXgcrbzys9w57iib9gPuvm
k5DKlwQ0PkwPArHgn1NifZJB9OgV95tO+Q68S76TFGKuB6VUk4/NaWv8/Jj9Pip4
ObN5KaKYBPrX2i5QBuf86O5XLFC28NJg5lE25IEcQuJmwmQd74tzN4J+CSqYoHIC
wYQ0lXteLFIyBb9y6nMUYAL9Ygbtv9IPAdb3YnxAWb0xM7eH0GxyCQ8uZykgGoAb
hQlLschZaqY33pXzNP8LqWyi1f5OiwTsgyPD9KF60adPQZZeH9XnbF5bHEsqLlK0
La61zI48y3SgzHpsQ/cz+KcgBnkakFHFj629wTY/zzSRcpm6BTVBUgyoNgnAaMk+
aQnEzPDlUag9byFx1P04toibf8Rc+DNISAnVMgreLRK3RPAZeUoL67ibwPjifp8k
I6+Qw8QtXBM9cOfrBqPznet6p+lnmdv7PI1zvozUunpcK4YT/T5U3PuxihSSp6jX
Q71XiWkvdPGPV4wShYGQY38mSZvhrPyxbsS4Tb26T59iRfQ7rmqloXmkPTIaTtmQ
kzea07u96Tdp4o0qK6IGrctfU7tw3wpS83NPfrj5CKHrXobQpB1+CREN+TIckmpe
6dVbt9PH/nX2P5iIs2DzZnt3PaZ/RmtHxrc2kgL1mZxXs/vQdFcYmnqCeV4renlG
aRT1ZjzMTuBrcLmZz70kkckUSC2yvzEo4+ttXpVnFznGUnCFGOKT7XOMjzgz1uJK
8np9cozKbocEE3VgOYNbogmlD6ifLhkTJhdXGc4X6v7q63FIUV3krluRKA6JZE/E
eAaa8H9/eTTLqEsMsoT7jYPQ7KnDK01Degq/ajVbBYhpJZbWhhmdEswOaDh3S+oT
+uB97iPIB3r5l+4+xJNiofUj1yYcHGvj8/0Q/jpdDe+z9GMr7mDxP4lkuLahB6G0
uQXOxh1G6xMBUUvWMkYPV5PHGzRvPapn4it/C3JJz4Kb7wZaA+C8S0MAjXLaaAEJ
9djaz6H0FYIWAp9ZWF29nSm3mT1rCXYyAsF/FCEZMYD6GJF/XL5JkEKR1MQHbxNq
cy2YD794XqOGYvT45UVSZaKzYIz0/HptHLPAAiYwstb6/EVtmtBN4DDuWcqlIFsq
8q6dl78HEYIlPFMLVsqGzQC+0lrFLvUDPCZ5yfrXlFNK/jSNXgdPLXGE0dsSS3ed
iuJRHyAcU3a/bvvU8t4k6FZbA4sVOK+OSoJC+ttweW5m1bv9WvdOwEN6Y0VkGIRQ
ntev2PZkgzekAGqtBZeNG1G+nYuAWodn6WhwIMHJ5NJHDkWMEA9qwnllstIUReiM
hmW8Fpz5uVRSNz5onVzRueWfedqwHQMB5QEqY2QqA7UC+FXPEA7DY3TMsrwPQ9vO
MOxGI/nn94bJp8AaRT/sphooqZVpwQy9d/J5rOOTzCRebHvRMSijb59tJp1wIEU0
WwJb7sL03D3aR0UF4ct86HjWxuhehC+VD69mnVshVEPYDKENP+dwyZM/OTnqQ/QB
+BemlssOu5FKg4diaXkXjKdDC2LlyaJ9jbhSGkLwOv0OiLZ1vXzZ5DSPz7moOG34
jMmkbqCAbAfx6VJr+uS4KdSd4IxWqUGwMjrATFwBkqALCStv0ZSn+GreOy1b3odT
RdHfz7RnEYY9M0KfK1DeizE0uz7dHF0ehOSw4xs3osDaEbwFbkrw+Lm6Ke3BtI9S
wI9SyouYAL9yfkFkJUPoD7ylBvC6lztc2uEIJQlC48pOk6DLohAF8pYyW7MPIFXD
6mVOGZybnRd06rMR7ZEm/vuN9NCttdXt1WHDWbaGxY8+MbZIJ1CKMGU/3cYpRSbc
u9gOgvP/efxa6AJmTUTtXyxFWomKcpIAmvuSpKQvVGaCBFl9RaNt5hrg8BFDInWv
3NpzfAjiuq6M4IdRR3zSVtDoqBLaHYDIUk/LHvEaWDbURroxqIo/ES65LkFnRtBk
as4rucUXRtefMqwRtbfdWhK6Vd7ZPLvWeKHzmBlWNQvuFnElgnvQ9HsJKV+oH84n
MyZxhZ37j2wP8waQ9jn02q8IlQCCq8H8E2zae6xfo4+lIXTmPXYSqc1MiuEsgbjE
PoPXtl1IK/Cp61HKh457lXWYY8gKHgxypWKJxv9SG3rU/nZfkjpzT33e0/a1mzyG
VcMC5m+mlpXrqOodYSepV4yPl6/74egLWRu4kW3q52zxwrUXflt8v+gcIE7O3FT/
SDWSlHyBLv8S8LK5WDkhwkoRl94Y3NtlO0meFGPUj8LgzqdWnWa6/QCFKZ3sn+Y2
VTD0UuU876/8aVOEZiLaSA1VyPYNYWlS8pnDZ93AcHyfyNQyDL7k/tDUQ6FAFlfP
lURjd6lfTgzqbTHKpEpldVGtr/C8GXsQ8ud6Y/Ua/SqOkvmtZk0VwjsRU45LLB9u
uyb9k7n7Dd89tWB7DiU6jsOA/EHZ+tDGQWr1OF/2udlkC/fv4D+hxFglBxL9fhfu
6bCQyc+EAF884WsWCXX2GzoNE1idsrjvMQTdC4He/4kXeXxOECnM/zezYnShlSKa
JDIeymVKFkJUfDlnh6xo1fiEtSOnhlTLy96dU18X2a5n8PYKOg5fvbLVF9lejCGg
1K90yAURyGCe8La1TijQONRKy+gubI4Kzdd6pJ6irWbceTBSWkkTkxi0dUEoqAxG
CDCdcuGEgY4rGdDq043oASKqjzNAE7yaH8ZMZIDV3qyv6dr8a3oKiHQfiZI5WU6B
P+xvWn2Uk2ItuAeiNT+9EqZOcuZTuI0ALP2vgGK2thXjloEwHeKjN4gzMw+007rD
CijyKxkejXar5vq68ViRCenXEVN8kC13XPpDa8CzrlxlLsVmXsS+Q+GjfD05Pd2c
IuTfo4Sy+44Az6eKAZJ/zO9vJ6b5aeyqOUxXoBheYmbw2jRyrqkmaBkkPsRpph1T
zPtnsUW3hmZeHToypCYKUVBIkaSprJMDqTEHrjwHsZECdqpqGSj12fhV/XMQk9jm
ebyOwlmPyu5GZ8R67Torr9Inzz5Z1ClIqYCJ/XWj1t5h8F/TGwA3qQyMjaK+OUA0
FEkSozgqwfxuNiBDaiE1YsNzjtozxexBgQaNZXmgDzbJUdCX0t16zjczfRbyR0wm
WBhEPiQuxgDbBVklmy0Of2SEQmjtcNeqlHqU6h4v926RWaXhGH0yRsuRaUG3YhC7
8vo+bSt7ReuEBLn1lTu5iAJDcidpJn+rnpgQbwOEv/SyHTIi1J55N4vdGy7LB8mV
oyH+HajsyIo6cz0apXp+08r2JOYdpdo1WBfoKU1/N7Tu/wQjVFf8dnVLnxaBQqwI
/o/bAWT7fn74uoWx2iyPvPNsOK27vASyOThCIKPmV/tUIPwNqXAK0ryPH2XbHWe2
DexaD/rVIeqMqAeVUYBGXNKkidpZae5b4TrjpzkftKI/SNglNQD5iYmV7zBCdEGh
CTzapcEkxJtgqVjhhExgpSN/CmF3yfChB6ke634YBlAzd+LfZHlKZnt5E9O0eAoU
w5Y8AOnT46QJD5CPk2wjx2oYk9yvqejVK8rwKyLLUnqYYtlgYYq5NT58KATS+jXr
/l8i+RetUxyNBPWkNFojO0krXCj0JtNWnHFrTpEh3Ige72vtXBhwgPF+Wku1wHud
EC3kGRCI9lS5rPu36yQXaXHTxPbulAKnsrzZQGK9Cw6C4RdhG5GKlCf+SAW0thOD
0Ytu+bxUHleh7yMDrqP+jByG8EVwGJUMDuSFVq1jxOsHuZP6QuzYzWxlA+JdvM4H
ydQFe3RV4e7bhaWPFvRaNhi6iqJ41WJXNCuxcWDjrQV2/4IkgfaRJc4gp02j4hsd
3DWCfu/8jtb6+8XYROCpNM07IK7OrfjSyrXDRfZDMLvErV6J7lRfO1xcGpBdL/X4
XJWzkCRb7YXr+Vi7ByaEuENnyz1wQDRODLcy+yCCHYh5qdp0EsHzMF9p/7WzhESc
ryv7+lsfRRkpoCB+YBDVZtva3rJ/4egRdX1yOJKXhuGTF/b16pSMPrXciJVkUSxp
xMojuTODPQpULGCCFwqrxRAZMEDUR1ai2pIcFiSvz36qLTlmOD93jC59KqNJCQDi
vIAN1Sl1F6uk31zBr3inVT5z1ygAhi5L5TC3O/jwMo+/bUuYapG27IEHsUmmcUAB
7+jbMP2Wc2x0jk1NGMn8KIEBJYTD0bMuA4g1vE49o94ZjbnY1edfNAyl+9N6vsDN
lgXO86YSQaBE1lpnLZB1Nlxv78uoSIlRjAqMyO2gUq7At6o18KhFYVKhElqK/C3z
0MnSs3oKUGwLHdLWbknUf5fa8PRe261Cgz3H2zCfcfMDmXUR5zWGEOg1OdOnW+tu
Mh7VImgwRiC3uPG9CcIqoXISD1YwMVMziMJTkCkPFq0WaUNtui4H8KR131BkTnsQ
XQnmzNGMuuMoNZSC03VD7RCCyBrbRU/r1g5s5hVeaBpMmqQYt4M+qtdrKB97B2Jr
sLT6QvbXB6kuSE9FEN9ilvQJUhlqwwy7J7yQXaCE5NdGSdkiCynxfTMkeevdi5/P
IGG+u7AZ4YqUH25XVwENqj27lNPWkVAnXWtpKAPhMQ1qtLYO455Kisy/iB7mmR9i
AA2FJPhlNTHaKRyrLhkBzE1llBXFPpFFzzE1BxXRkLau7EOq8FWHQzP9lnw1qGGw
Iv3qXvtd5vl9STdmfPil11T7V0YC8GBlcLiYjyzi1O9t3a5+IpNGyOw+W+Rhqgdx
ajS/vIwfnplBzzqsrz9+U5gZiL2nEEsCx7bivlmkvK9OsmXkvfWKh5r4p2dMpQ6o
VeSWsjp6xKiuNeMjCq9K1Doec3hMVqOipWtxWS9+U7n4hNqTaS5/l9Nc5dbh0zVf
MWQ/8Gda0C7NYPlklhakkVSg4sleeu0qgbMZOslx8tt6g95Be+U8cE8HJuowIk4/
cgyfqiy+Y0RZhIiNpmB0WFj1rSWT06ivgTXIzbVwIkp44bXhv/K/b6TYe/kmCcs1
1bETW82cRxwxdkjWQnXMxJdqiYehHmSiEIzaCqNR73wvWFoTXEPLtZU4wMpV9tbx
3zDmcGPjwFCmpWHFe2jgbftcY0i6jBOC57Sz/dmu2hec/1Hb4GBjJPiMsT2vCLOF
Fs9ueFZ0x8tIPxnbxg3atM9S+56qXSQLRYCqqtBKhAWwN8TbeXBP/2nFUSUA4VvF
dXQIPNu+GTUKku0qaY49CGniLXxJfkxrzhPghUtOIGh5KA3ANq7i4eNpNLMa4dpU
DWMH1xhVzitZM0tjHqm/8S3hED5iYaH6+Vhw1WsDWpX3vlrGjkMJIem9Y9ugFdmD
8U0txB6KDuFTkZqm3CbfjzqXOi/CSXDM/FBCox5X9ZISFzfF6bpknG0DtwV04gw5
Xs88r8B5TA/D+ZCPwKJDj3zbmsQyTyH9/gUicSnKc9Dotq+CBgyYTmGx2tIjPXSJ
cQvV6rofPBAYlQX41ZuI3+hI1I/od3iziU8GBa3T0E34o5ojC28qz3yK3bHmhWZT
jdzRuRENbqwtDU0w5Uewb3R0jt4NfVodvRxzcafynwYfAChUPTTA8EsjM2ij51K3
CzWNhSTnDLElC2v5Rhhshio7uKabSBnDu/dAIJqCwR56pU7qSTb3w0t3ZeYL5MtN
fzWmYALKZYcs6J060cxpwoEs4SWkfgQB4iGRk+EduYAZ/njEu1pqGN+642Z1McD/
2U9/tBt/iOI6ChnfZhoRPqA6BTdlxbJAKjFX3U/7i+hnRAUovji8n5LC5XUIqQ8l
4uiRTOXBKfvRI4h291eRBFo3SDePURuR9NdzAYU/eAnscBvRB832yaejzm3gjl2m
HlaK5m4Qf339R1Zfu3O/b/SRcZyj9Jg0tMuZbwohiyGRvDq07Wb6YeAVjLqSFJJl
yujxjd58DNmKR18ssYHaM3zW2hDmIIHk7YVTwBLWWmc/CCLiVyqfTH60ComfUV0p
4x5rh00vfYmAZ56LdjKgHTW0xrt84Nt7lf0zAuuH3v1wU+T40mraQBUegYPpCyeN
P1B/K/hHm2LeaLHQcOQTAUAD34PnQ1iEPYVboPM38XEaFfpS2ZIj1JORSK5N55WQ
JbV3QOrvpM68EQ3bD4Rr1ASQt6TPZuES2DaIvlYCoJJOIf1Z7KAqTu0rUw6ct1Qs
xrC3ciZFyqnOnDEyfqhandwc9rvM07v3yuzYu6kt5YJprPxix7N/DYQG112OdEp1
6r+6xP4WGbLnIhU8UiIYyd9wmIon1Cud3QWqxfuT6o0/QNLWCqr/BkFCIhHWwnDU
C8Hf2y+WCKMU+hJ4RxucaCp7t+aqfgMa6lNFoyDkl76u7D+BpG/O/f70CKBgwyK9
2wemoKcJGL+GGjalugp6rJiOwQFv5UzBCEwb8schHg0irKoyTKl3TGX0/WCdh6uI
AWE92Qa/t6LCwvcVOb8Hw2Lz8XrDfcHrA/m7E1RG3uGcA6Ew1LCiCNAByNQcrvpo
2Z/3PraGG0751PLv+adAbC+RGitjl7wEsIq1eynXN0nB3JRnYp8ydyCUcMdVYuKb
Z6wm9iosKdpj1y8m7ACq2sGq6GxUbA4ZS8vHY8xiIT6IprEwpBksMyydpfanY1+x
TV+xIujwpd61ORogdM8NIrh//gYZ11zu9O/2PiVww4YzuUFEZMIjBvttXw+UnSVe
BMRVKkOmQ+53fr5GJDlOQ3+OgXuykI250JDf3+NqbDcARo+PzpXy9E43jGuc3vkm
RcvRErg5kEZpdjFp8c0x6zbjsPwpPiRvxGjHvFtt86gN8LpXMpcBIy2jDKc/SHnp
AT38C/tlNAXR5HRE/tbNC6qEXvf+qe6JssF3zD2DhYo3lvtFK2bfL2pycqcoABw1
6LY5aRCdfwuq0WJH86/y08oHwDs+dlsClKdMt4pzlEcWPDrxvU5tUEUIAsUDc/Dk
M8hxMou9QEAkpaKgd093XHSGZxL4bB/OPkxmgtZ0XgFSsQK06NSNDELWm0wLx8e9
uackCDRPWa0BB6f4AeRfUCk2mS65nnldmrfmA55JeFTqwfNP34ryjXpBeQGTK4Jl
ghZwBxpn3VHMAP/blizXsDw8SMb13MAWkQyUab0Jl1+6ottROZ0nqPS6S+FIXQ66
J+6dro4rdNrcVl9QEnKbyOqzRWvK0E4lR4lo71TJqx0v5BuJLwWwB4bDydosJxpB
Z7nPPVCXYvJy7/lldjT4Hn/447Yoq307pTs1fIDdKYwffdcDItSE/p+uYOf+MTA6
JSk/7xPh0tAOJEbqVW38Zloki6Bl0O7uQvW507QaRDZ+DBDSyiTktv+Svj1S8eBH
iCuPMamuAC6k1tqoW8VJ9w9VNZLatoDZu2tPVq4Wu0xCEjz5orzijQTpra/JiVCs
I2Q88EyTAYhsWnF9752ZC4c+9gFFIwSlWiVqoWJrSxTVrZndgfmULByP2UJFgWm4
Vqx7eQuBmBbEex/FcRHBQBSYhPZg+MQN5yo+iAtj4GXHX2EIMV+TWXMa1pucVcqg
guKjyR15j6V8R0bIeEBZoEDfzuAvGoiG0IwE47N70AeJgjxeBzV4n6yDRQcrtwVY
B1u/sYLcqzBp/mK4fz1yBCJv7beUWGvGaOHVy3BDSnPbF5Kr8YOMaV1sBqhjywe9
DIBxzbEOVCr56QmuBLHtlYd4KnAseRWwGL1PghgbkjaonpkQS7zdly+sMdfeJm3K
/S1UtAQSQZnvmS6oABqSZYj0l/UKfP66nRrpmeI3IIjjcrwZvVnxMVEyZlQ4cGQR
RakYnRvQGdiqYkh/vXFz2t9mamXmUEl3saCAq/xnyTwjWJezGoPl0DoDTN/hj0Fs
AC7VZmGAehC+t4CBrz7m1AnWJnmwIR9p1K0MCezvCJUi60eLzVftnHumXOlF91oN
PBMqsxp4PeLhbeSaEelgfDBSeCaByYQHFNfR95NDxgt48emVrnTIMaKAqsXPZUun
Xm7hIkFBES1k66GHrbktPP9mJVx19xs4DXVO6AjGEBAJvlvf79qjFSvP+OJb/WGv
p6ZyALrGH/tE6JNUmwP+KJ2S/ew9LjDT7ygj1OmibyWO9rbkiaYxRs6ygXl2Axoy
HrZEBHojlTHP3+PiKRQYuUpaXXGCmI65NuoaEazK8QG02oGDcb6uG6eIt1dhJlkg
zVwm3iH2vZgOA7lT9f72MnxdFkLGAmvWj7Dg9tVqp3WWUlXM4lqz7lL2n/vZrHue
40mfnb5cX4oY79HQdvBQqDn8pwSb0dzgqo/ycOkHE7OxflecnkcONIailB8wRGGg
+CePrd4IMMCOCu8FmsmNI8NwGTb2O77Zbwx6s93hS7jit3rcBxemmcHA3+tnRv1V
DvvXEasJJ70fIoHBURruShNHPvhUGIRE3Yg3YVjpOVHIxO5RFlAgegrHl8kXt8kT
6Dw+lCfYc6W7nlmaxAhJwj4CDY58Vspy2Bfw+VlAUtlm7OhTVKblSBFMKNsfzwVj
dDitLAnvN5xItaQ9w28O9XHnjTdtFMjIAn3/2m1k0oQFe2knCGGjYtQkumJS1Dp4
+4quQ7tKoOAzDcxsdNnTGEyPEHf7RTfKAAQvCTFBJD4xpox7ssjtvchzQjpl9b9b
QwQ2bTt2ZvwtJNnWJn39Y0Kyo7H5vOm6Qg9+xnAwoAPk8+DidAOL/s46MphSu3ez
2s2KCr4y4DpYv/f8gaMDSQcI94dFYtA3UPVWNTMc+gWpYIWWG2C1hDRhUkS/oDjC
LG9G5REykOmK09xZi06I0fiRr9Gyvis0O2qgBW1tfQiQ8FHwkezX3F6JsaAUs5yN
uM3ovJp7FbCoyMTbZs+/mk/veLnYU2ovFfJ2MFPqRMC6tJXr+n7rD2MxtCR0whzV
Nrzj+X/RrK6TqnKlI81crAKYwQENTEUUBRV6nFROEHvJ+HbN4dmSjHqJQ6WdfeZS
ZtyIOuLAE6rH1jNR2hlYtQ+c5shNxmj2ahUdTMA6rQyG/EFJc7jJS4JNbj7UYp28
qxCsLy5ZDE25FSgApiqH82FvkAcxm+PZC2nwtE1gkHK2jTjySi0RTnpBhENe0RsZ
hEk2ElPFmDV7IHAh4pQSwy8f+/vTxnYCzmqrfbko+doA7t3GdRM1kQmgNvWAT+RS
qDyS61yUfoPJRNZnBfj/fFX2PbXRlegOD2ukyZV8C7L0kYuvlo9CJCyT5Z//3yPc
qBaPFtYf4XXMCLe/mmmGT7dIp7JtAiJxAmuAgXU/xN9vOFLfGHWFOZmw1D63K0za
Po+saYFW0JOA2UnkKRxOo4oRiS2WNBooM25myz61YxJ7VfStvAXLfZtED9HPOQ/P
n1bSyF3R1OHjzLnm02gy413AnIhxRK0rETj93R5/2tmpyAfQ9ICKV2Pe53WmM/Yo
IN1uT6WVMHQed6uzZ9ihHvxu9D9vl1FDItiKhjqIElSmUpQSBrZl66QqrYaC4tk8
lhtiHEG/Ou2+Oy85KQ81Z3YX2W1ay1EM/VUiwm8YOyvEYDPcfcYnn76n10+h1mZs
CK/uPUtOmiXcCdDSTc5RrthQ7jVv7DJ/TTNsCjeI4H/U0To7TjV1aktiypu4AoYE
KpjR6MWcYSihHh+dxHFY0OCh0AD0TZrk/Pd9Sz2P4EnZjt6IhOumFgXxiP2x8YLz
vEP4GETbGU6MAMkvfjYJDw+WGdUcyYMoIRD7e/8b2No0FNu6f9ovWGBXYn0La2TL
Pq66edtIGmfOb6ePnfK9MvEm6omx4JgLOOX/Su/38TGzYV0+1JiaJdPxHrx8nrgO
7GoQcChHc+J6ZCvPPTJ9fU18QMQSHv2qQlTkOJBFpQWE41oiaiijm0FG/kjuVQzx
iDYofkAVVEETBid5RRsdkaRsCu8aezMJrmi0Ux8+qFYkzh/zBH+gSQUkXeyBJF6t
c1g7x9GZZeuIBk7/C5ImLQ8XZ5REseppCRmTJeyuYoZv23pGPjC7wQrnYYlI6Hh9
p9eUhuSC7V9lwcLOD0WNjyIaxUUk0SQMZ40batTHU13btBRVBDOOrdVn81gL1M+Q
1nBI6qqaiCikhqHcfXurpk5DhfZ06LGwLoDEgMW5IpFfBCblyTx4qr3Ip79CBZzE
kV1zG8Rdx5s/0UUcXS2OX9dku/L2SupOyvP0ip3DR18S+Hm3pSRQOc6for3R/md6
1ov+c1aQulQubJyYaTaiAsetOCWDS3HU5OPupp2oSh1ZP8PH7zcH7Vn9neBD1O7u
7LmAbQefSuN2MStpZLENdacQhik/dg6X4lSmwscc4OpDKXuzWV7/ae+gjI82O4Jl
NdqJFJJVFBzwtM5UQaihC8md2upCw2kQwIwAzw5Yh/2cAwoL83KVh54/jMd1gMdu
bw/VB8o+DKwr3N1CVsQzOR5KBckLS6tdlFAJyNrCwbCItqJf7JoD6rLW10EGI8vU
NU4ynG5R1AmqqU3xO0YFxJyXfsiY+tOXQfcMrvL2C7tJBfMIGxqXl57RI6kfhf6+
9Jez9ato+YhYOgOlCQpRuYxmB9IAjCNTK+GeTej0OAjj5qQKb3misXge8gmljU95
1pZtoM3VuKR1CmnQHvQXC8EzcmVKKxOMKRwegZe/g5kVjRHggIbB/JkJ4N1vn+0n
ReVRZ4nXA6t9rN5DpG3+tbOSxZbbW7GXIAuY5QwbUUMSB5oPnDe9zYagev9veuBH
0B3w0zwVC7ll1SW7dOLjRxo5NCNokhks68IFgbmoo1R7a2k3u60uOCN6BBKmjMvc
DpVRFV6iL4QnumfAPH3ZtGCQf84bJT3CIjbtwmEWiCJ3LIUbj368NPe/WzKyzLWS
7CoGsBjRShlfLmjfK89T85/9poaNUK+DZNdB9UsiSdb13lwioYI/GLMbzfPkUZxO
XNk31DOemAn9EOPSjrCPMCAj4+PYvSf4LTh0Sj+BYyRRNkQxJk2Nq7OUbN3yT5Z3
s9V2bWFKEJ4zQRKIqQyB/1X/3UpeeQY5QEH4nB2wN35F6BPZWGaX8ytE9R2pLcDT
V9PHzmYhqvn1z1em1XQRDFdjzmIV+aPgbiUlAHJAHb1VcrjIVHnfnIYpz1mFIB7a
+rheu30V5Jhxs7lOiEpz+ijPzPRR/3pqjmOlq4Jhe+e+0wHkC1GR1o9D7+wwtxcv
mnmJe5OrXhOZKufIHnhUwdmKp2QV39ZD8D81FfVG3DeJXW7WIGHUswXlPegXd605
du/v1gLD8sMtZQACsMZFdboR7vKuiWYFsScXWtAqkThRUYZAABVPSRuCxE951U8j
xQ1xVZrU6KtJ6YesU3bqYrGLziOmnN5LKONnQgueVrPgwShU7P58UQx7lLg8zHi3
zCH47zGexa4TtF2VWUTXSSWsj+zqMQ5ihdmSNIP4XZD/RdijdFtSue/uJbWbQ4oE
qb8HkdQthhJ84KavJY8hHiJgU7uTf5nVuDYq6sNK7GpYrI+ig/81y9UIXY7jLXLM
unYwn4YpUDBbnR+UybEOrfV7fDu2uHHt9siTS9gVVKKxtw0DWRj2cPwDvS3LqzDp
q1bqPHnbTffG9lsIipa1RGSpwmiBJw2GmIl1i9TaZTDURDTLYDlK7/kl7CxGre8v
BbvA2h3ggKMkrs2grsFRGQQRqPNdvIAgTEl5LjHeRNEpRjYvR/a8MJY8M5o4VKod
moCr+3q9CMlglxk8cU2U8iMR+mLvoBbmoLaUv07IkWGIDNoFDyljEn6Dwy1gGtA6
SGO0VBU0c6jtO3eVGyvaTFdGUJ3cuNXD9NNkI3+L1RK+XstTuL9f9IAv8JzkMbci
I59sJE2BoXSpR5m+D7oktirMJDGWgmoC2eV2GDqo3lFMj3wXsgO5O8mgU4L+diXZ
83vLU4Y78bEXemK96/46/i3Smdrk2RfIiF7uXLXCp9T+kDMu6McsC3wIP/Ba26Nr
2qcI/lAR1C1s09XHI2p7Y7LoQOi6U2ggEyZf/3fdN9uRya+ffE5xvqRf55KqcGlz
YYtK9WsRPXMUOfmio+PlQpcI0Z7wkKFkC8HUjZF8n+R28eC9XU6UqudtiEzT6Paf
UWyYdOK7YyIm4kHAST82Z+75xmBw6JnbTTl6Un2AQGv67LUBYVSVn4RRSgnye2S0
0zCeUZkNjxZyRb1ltYNNejMKXMpZACJ8C8sMpGu9r+UxZMzAMqPCelx4u/5aBZo7
H9GwXaRTm1F8TkuO+ghQsFQkC8yG0w3cYN4n/SCbeBMy92x5Av1D1DAVuowKTxuR
4/sCXoyyDSfSdG7LBybAgSAdMrZKe9Y0CAHmQCGfrOkmnpNnIsLR/0oGqwgj+Jwt
PblEpC3iT7CFo6xMHZ8sQcdl6Ai2FlVawlJNXHXrkze/i06RWjz7xA1sKbzXg74/
HuS6h3ADkj2LLh//wwcrnpbv8Z/yVrWtwypWiAbhd5jlVazKKt4xemOlaOHtICQ4
kevR2XWszBMUh7w20x8sRP4SJPg5iXDRoUJ9X+gMU0SmqsVvNVB+oee4B8A9aurG
7lZY4Se9lCa+aRW8TQ9zaXi0+bbRnG8cWyfieAHdTMtoK1xstgACftqb9f5aXiSs
ZT0/v912XrBAUEI2SUq0/btOqlQHiMw0Fn7uUYsLOhHmpV3Hb+CZd1/0BXogDbuc
L2lczwhhTeqIsK1ajhxsV5FJshwSnaUAiIw+L75qcunYpTl1S5G2I2pgYDw71SBI
canzN03cVvhzl9GKg0uvePASEXoxh4QykjTEvlf7n3cN7eLK0LGoGIy9gq7lvhLQ
VkBlwRgxuk0MIgwqpEitB5X0P/oldTiAgCBhOyTdNWgL9VPwtRqW69C0XTIGJkLT
4v2zyIWXnge+rpCmNy96EzhZO7nU4+G5VunS7g5L/Ur2r8qdlM58rrPTfmnD0loC
WewdzUCWrPFUrixSyJBg/iVllR1UqEaGWFwuHBcWJoaBSgL3sjbqZpQ3XpjuSSBM
1ydBd6gmVVGQ5zh0vKBoW5dl9SMp0FY2NM+LEwOiO+MlY+zZ9+BMkOmDqp0aEKLB
UP2MFem21opndzliSbU5SkRBeyKWhmghVIk4bNGFLRgGrGfpgkdcO2V7OTGv7Ey5
lspULBZ7Lr20ACzCh3G4fL1w7qr6WlFamBufzp8+beZ3mvydNFNy1NabyvhV++ZF
I7UHR4b/b33+q6ZX7j0RUBuhcQVlNDBNCUo/rTCuUxQaSAn2/Qec2no4uE6pcISd
to0eAD7v2/OGsZsXUCn1+G3UFEaSGAEvnEVE6v5IGkYE0hQLZF1gIt0N20/JcNpN
kLegKC8qjSzdWfsV9fAAUlnpq5MmDcVn0sevedu+ShT166ktklQRkRSjAlCZ+sIT
JbAUUFxlroLY4VmanMdbpUIrQl+hVesIf5mjD7X3r4ltIriendhXK2u/ImI4kVFd
qDz0Hjr3Db0nhz/jOaVMHfOqmIQwYxcf+m6LpBd6+T0ktpi5Hsuh+8YyIWCq84Mb
LeP7SkQZferfD6XFn08g9CpBeMA5r3EAOLGzxlAQmCgmMkdTUVZ9VsrtftxZYiBy
2pdQ/irjIQHkVL2Em7Q7ganz2tZrugPVEv3R/6gh8+54FcWVeLuNazJl/G9GN6Xw
Y85ZS9FwWLDJl8C2fkdkHzAqoboiPo1NgJaQubkqGJTltezDeGrZgqTszdA4BAfl
vCIXvfUM+mbN8/Ad18K0A1f1NfTysNtz+BzsPdemT9t2LLC0R3o/H7oPt8l26zS6
uHWTx97e+ad+d4UpwHqjr/rZAC5ltAHpCt/Tu1ZMHeGIjeP7HkCkb98MmSjOa0hP
rclh7Xuy3dhSpeGx5kohbOZsy2dGZ0fHs+AVB6myqvXw26MxMPFUoOtATyxFIDDA
nQLLPxJ5wrvCXDoQU4G5uzOXViwRKvg1q2shnXXpCxCZj1wzrhAWPrp7PJfXW6hF
gdCQTIcR+Ht4UbL4toAJUC4lIQM1vxgCJWwdvoMy9gsMNlFiQj3iF67HYhqjmu1Q
9oupq30KIdvWKdb0IoXMN2o2x5RWXuqfQBa3BuUdL63NIJEm3MSh9Hm1/9tAAshY
Mm9gz5lqEyv/9kPUcG804iVuBPkBbFIfOsYMk/d0HuQzLEPiOyb1syTgmV6DvXTZ
xefjCE2msOOhLccO2acoRpWOHlUOpEUSmfpENLaxdlcGeRlqrBqwoE2653LhAdTr
Bmv/eqPrqy600zSlKNafzPaDaKaJE+guy2unkq5tMgW0ZYt8p0B3nDZWp+kuhsFO
vs7u+DFSWLFtNUVqa08qtPpr7H5/Gkyt3xBL+A+6HgjwNcpLzwl1+n/wfDCSZhR3
oux28czOZpMFhjzGaQpakHXeqnw2ih4G61r89vdAaR0D7MauFBVGf3odSO0oiF9a
YN7SUDCjX3d5f/GTYTlIxosiaLn2/v9i2BBBUTX1JYoyPrJDedh1TqTylDftzF76
R/vCuScvt5igOSuz9Vz3Tpb8bbQE5jLBywPtVi+GOjXdQjACp0FyFW/dCVs3FBgP
c2KJW+amodVvjS7s5ULUUZl0l9MGt0rjNVFKbyjnyOOZ+HO1z26KaoPwa14nbMBQ
vwe8tiCHmX/ToBZgRlS2vMu+zh6AtuUSP1+HnQvQNcZM8B1kWeJl8MDkpqDL0eCO
cftzpW6w85PdIfbN6Ha1YCl3K2olwPrsGaHjuqdfnxFOp8/W2RtiBJl7Oj65koWX
0+bBXPFMwI/I6fj8pNuq4P/zSgJUdqNzQeqZoQoz0fPoFHO7lLXLAtyx1PXCilvF
oJVdkBiUMe/2azKptx37lCBU9KTtvxCn3RXpJIKd0UbqfMlw1Wdv9Wgwzoxw4FOC
8Nrp1t/+5A2iXN06JT9AUvuLCIuoSCrJA4L77XegUJ9LkHvwyIjZU9hWW7aS3OMI
kfpfeHhyEn2U47SRplrEkwWknColGRTWVsETrLQQCKNn0XH+6xpzEE+nH1w+YJwv
IgMhvwOotpJi/B/E1kp0eIXn5tNyYPKdHvD61OL1JmwtYaX1BS0AXXx0OvOCV+Vg
mazvKOdND0nkkZ4hlSHrI1j1qnBQuwjEmcpNYNloTgQZu0AP0xsJ4wnAUgCpk1wK
NoS3mb6e+xeMk4uNszmeVs/NN0hL3cY5sZYuvD3s76BwMY75YunTjIZCav3Orzhj
Dh2Pe0UK3UEd6KKSYpxz0huORKHUs+/mFxS0/pIhqzlI2vDCsk/ZpxjMppswc9Je
WGo4N8xXbtvMD2lYrXUnb+61aSM116LxqeDiFX6VxJO0WLG+gjkXH0rhc321DrCY
SunQE1SyntIfj2PdDWne/oad0LoB6tvGoK8fqJyje6ijk0CFMLBt8PT/FjqPcS7O
rkQnz6iJJLHGRXqZEIAdqE3CZYYiXs7pQ4KDD3IEYjfJ5rHpO1jg+zKyLlMboips
phhe8Nph+qqIrlu4gtwcVBGVF1gxMNthJjupz20eGosWtXsr9AYu8n+JQta72z5n
mKrrG5zlsNtL0GRpZLTJr/zJRPIc6KcCjj7V+P9kw7Yp4vLkE5rk6LoXgo8kgdC6
rHU68l//zTXxP7rnum1HyKudGPgAnSTlqmEbYA6vXtoIDmeH9R/p4ROeChcKifOv
F5kyQr83VdQQiiIw5aQfl5X1BgpaMMovN5MYVHcCPC0dwAz0Eszy9wlHYqaYObqm
Ao4shP0nWGjYig6aqOrcncGDG6/WRjAtw9gA3vHG+bN6mSsEy/5F+NG7621vl2UD
DEZJvn/eLwYYNdxApOeZTy6tSBOsaEX4NSr0V4Hcni0dIrSlXn71x6a8te6E1EF1
O9GaRmri0AzMTsGDLHGo36iYfhFcpfUANIwvEjuUlm2QfT64/fEDSlv9mOyyByU9
LYhLxcp7qiTupZpCVaT/mw6I81dGlcwhLLkVQ/b+uj1snaqUgw+zGsxF49lZ6AaZ
hxNEUAz+wiDrNkW9fseBzXANvH0jwPVd+Rmgt+Jv7J1qCMXYkpkg7YT5WXpWR07/
83z4jjjHsdhSQapuZgjY46IMVVFru/8oJLbhb2Gt6CmLvk93WGgtuXJ6aIQ1uS8F
lkn6FkFJi+PlXCKS2KrYKY+yBxNYjBvpifXLvLryVt0GeYUKvAobaUfc/UcQjIUc
aedv9RLa8Gu+L8lyaqkIKd8nKTAaXljzr0EURyqmUPdrWtl5W9KweZIToHZk2pzp
weGNtYiZBzADQJplcDLJdceUnaOJygm0RnvzibZAVVKdqVXVFek0k0O/ZDDkvXfi
Fbbj+MWl8Kc8jFV3JYTAi43S0MLe3Xpawns1fx1IpOnRFXaQfs+F0tEtRyQroySY
YTH7h8L3u6v/x0D+4S7cRviX2VOOYAVDqeypTJclPv239J+w/y31eK1EGqzDsOeB
vyTxGTXeWQff345B06GIL9Eoao0sFPooWYmC+DBiew3YlGC9rZBwDtl5677Fl3uO
PRKn7CxmFYXUm3p1k4g8RjJ1Hx35QcWISrrOBB+4Csp/pkU3PZG6Wh+t6vvkPxb5
OiP+39PoajE7Ohm7Lny2WBvtuDWhXwq2NNAq8vMGj5FaV46C5/z2tnsZz4NVWINj
vUx9Ey+X4NObObpqwO9rVqVPkwkWavfQ6jD99nEUsuJ9Nr4DUWJxLC2heP/Oqzf8
gjWqtW/QYByJw1eWwwAkGcTWpB5xxPeidlo+6xQLYwAXddsXj58Q8SQ29dExOWFF
3WdpMyiglD8qFf0AWZLKZ0H1AP+QOmo6xQjMIGlNcPsZVTfy6ARO8W1fcSM5DiEy
e6SLS1T5SThd099cHDnHDXurxDrkJdUNMnELWQaH/xfUexKkvukZfMsyKU1nH6iY
MUp33oqwg/e7WOu5xEEd6pwIBR41h6bENI5Cwzg5yZFhMKNcWXfRYbDeowY4eP+e
P+4Zd6a+mEEap9Sbm0ZEfg8uQ1GTITVyGYa+xL+/O8NbbhREIYXh+rh+P1NqZl7M
bxCU1OYgyUInROq4L7c/Tu3CRi82BgGwpDV4NGhvxY/ITY/rkmfUB2e+FCqnomWV
WH6fUadb6HFNLjrP2eiV3npCzaW++uNm4ePF9eNwyIzBnnjAkITVml2FMu9Zwjc9
gez3D4tbdzyarAi814bKsApmdPF8wNvPr7aOsYl6RuBjWKP3P7/wb+zpEoEdBjdh
p3eN0jJMd5gY7fHzLA1FOSeC+dPJvdDEkOCA5IiHp9NPNQyqgkxPNhVVUeYTq1K0
AGWqCZVZQWgEThbwqK6dzZi8l5voGd3NGKZawdpSNYtZl0BbXP4u7bWV3K2G5LrE
FmiFZSJ8JntUXG5lE5/FRPvo+RNxIiP7+YptpE1uGSbnsCST+zrwbF+YMikKNqUb
e3RaDN7ThzLIkUXBCVaGhW8+hTV0o82MVAbNjak8/+zTPRtiVTz1qNIMERxnIdHC
trePu6Bbse6nyuPAjYYKsz5mdmdVOv/zn8HVN5DvN/lxV/IPUjVpBG3d9p7F+zUV
JxkwXSrne5Hn6ej47Y5i3VY5BB8X2QZZ5MWCrOjGVtVbfib5Gyplwa45tI/7ulVz
qz2WzhPG9ieuA1ReWhpGDgdfdPC6dVGzu8CvkufkjpeckgMzzBAEHaHRVp09Fzce
/x/h0LZwtpDU0QP9EwIFyz5+VPjRKjLEQIOlJlUKYRMq2fjb3bAZGwwyUdKYPOLy
siHFU+f2tfcl7Stzqz3plaXQdJQOuXJ4UAMU8G9FrxGkDoo8PHUiBfySmzGFJh/d
WgnPWDv1FY4+6vKtNLlXSIdWAbelWsjvNNnLKpjwbru5Ve4bvpVWs7ZUCWHh3PbZ
eesaNiH3LHF/8hf6v46gRkxGP4RpU+Fwr4DASlkfadFftDmXyKGsm+yXbhtrKm48
v2tByapfxle5+ltzRmaAuwSE1qquYsL/P0wQJSotOTPHUnWuZVzoyjwmWhqH/4Ak
QzP/pxP00Ac39YrGCHLI7m4ZxdqhekIiL8ZAaGIo+RkmDO8x3EAYaHBP/kosBtRa
DlxZnWZ2Lt4mgPuAKhXiAmUnP+0ZAW7gpLRYjTxyFuJdCAaghG3lUyibKG54CqtA
+oTlZJUa1h3w5oywErJFdbvv7IVHuCizwLOlqQOkk6PqdVnrkCYus4dRpKu2sXKn
43foraNdSQaCMRCanxmdELOtyCTppuocImtbQWbvXGk8v5bGKwgpjpWQP9tyrB59
6elTEdkoR5/TyD0Kn7gWqVcDLcIiq/lhBrShlUXZdSbaQVeAotwqxLCVCmEj3/EB
saxjOzm7L3gsOCh4jkCCJLiu4qHE5YXOMp8M7CXgm4VHW9kyqgOp7JOicETAAODH
couweBtyEq4GkW4L/ALGYHtyWysQIlgbxZnmyHK3oxu+T1a4gmHHFLjL9ITqcfxd
sEYsYcxu9BG89ys9KGgdNyO3vw+kgBN6dn1t/ABxiw0rh009ovLy1iLM9pdQZu8H
r/oBD8ihmFDqd9+nvIkAhAPRcFCkVqMD8SQnYmeEpwIVw2uCAgJ1nx3HYrGsCouW
2PXLdzDVegVs0Sfe0QV5AkJq7PwHCVcKUU3UMltAnLL6OP/+sC3Jayj6xmieVrjw
dTYCqknh22dOpSiuQeAa40EjoAwuzi3DWDe8gZsM4845Yh6ypJ+ZYaC1POz7TUJo
d77Ts6kUQOFyeC//mFHlrxR/iU9AOmilYqomBJCpLe+mkmwJuxGglmDA1o0N+oGV
qDA+OS9I5JQRj1X3sfi0fqjz7UIR3EydHHwDe3gW/rYrV/I5X+JeXiKzk6uQS4oq
FaCzFHbfvJRmxm5LFxDePBwNu+4EdzBe4uubOfpKLVsj/cjHzHfyhXzPlpB+p6mM
kO7v73AM6pJc1vTBuqTTtfg6+YnUf5/8t7luQcs3YlTXYWTF33N0caCzJ+wFiPIN
3ptGg2uuZB9k/TpivMNE1w4oCL50KQXleSp8Hpib5MZH+vfpPJL9nDwh1N8bL945
zBQ5AXQ3l0HRhe5i3KnX1a8GeVFAifC6IFYYzQGurolF/q+QfS0IDxlf7VP3LqiN
ew36v1q2H9VEMpPU2kKUMTFrI7rKRrBAdBKTcLKxG01zFaBhnYi32cZHz4Ez805s
iD8n9GmFIKCUq1VicTd/liin6JeTgBa98e5VNbOJE28k7Vqt4NOvyx+GtMzDnHdB
zerIsriTHCmHbuBc70hXgTJAAM0n93fu2bTX1W5USRLPqfPt2K0lVQI8HNi4Kb+W
XlLB024eDOHde+edKj/V3koo7orzfegQS1v2vsrdnrG5sPJHDt2o6siZ9oawE1CZ
+gHh30z5t79ceTGZtoLUJu3qDu5NQP1v5xiS2+IpgslDNOa/rd2PF/jAxTnmTK6u
dJ5hU9JjWmmjUM3HI+iUW48kw5Lc0j1fFb84p+RBX8q01giOlsa7UBKFnLPnSoyI
jip+gVRRl9LxIBo27HDDYNRbYnFiyytKtWBtZKBgHluiCxnQAfGw85rm6EwJLVwo
W4zV3lKRAELL04e44HXMXM5A4Yz4yN3iH5w4rZGUn5mItkigD9LkUABHsyPF4zlS
NmtM/IYFwbyXlLUZ17Q2C9S6NeqGErx4mVTkBcfM+Ccd2OYmsuDqs/gNj+1HUPE0
UT3ZSgc2lj3ThYozwI1z/RgZrEv8jW3HJkdNxWXutTM8V4pISFT1eQDvQxgbZQSr
jcHMgkr/01RjbZ63bzxfhqITO+TTUDtIJySuWtRp5UyfMBzC0ueSxxTRqEsG5zIk
IDPCe/nr5pSxMXk1koR4UdxRE7P96trkTcZ45NuSSJOeevC884awy0IFNZbYrML8
yqfbJwKUw0ReL+U9rtf7X4l3oeSOq9waoNBHjABfHOqPssd7+eiXzlYlFiu3YIpH
nIBz2EEzCxHPYND51z7/pPW+LDRAyD9xgwXyUvwyntjmCwwXV3jJkVUWfXLAtdHP
3Zig5LsgoXBuKL9ENwuDiRa2XjAMpd9DoRSzGKyfjRZCqVgXkDynO6SQSwz5vlEk
WgR6Y4RSJ67RGwvj4E2NYk8vYdaRicCHXDMX3L8t45tNm5QYpcRMWCC/dPTD/OU1
UqsQuVC+mN+/O9MHxxCWyVQpqTWu1BgfbH8PLCcFNxZm7Je9ALuj7ZPdDAgzUrmJ
ci1AjC1C6hVdPIyjbUOBH6Cpnkpj7S59yPSiOdUYcuvd9ax7HDPY055+ChfdzeDw
dP+7M+qlHo9+Q5xk7prRklFnbBPy6G1vUTV0ZiGLi554aZpIJuPgQEZOzLlXx+Z8
EA6KsjB4q7hO4sWyV+rj9viANR7qVWUIR3YiCbd4ZZtNeviYaaIeAkiXUVDHkVEu
f/76qxvuo7TcXyzi1Mb8UB1nwKUAeYBLFktvpmXo/KHilCwYNPhb33+RkNn7/ehm
kkAvs9P4Yr+nL1xYCeDY+km2wQFLaSFNn2gil6phtEV6wTeMIkWjRMBkjPI4vC32
UM35f4FSKnUvkSlfLY54g7QpAJGlq0Js4p49q1di3ERtzyVJ68I1WYAH3xr4dDvs
hN87gMjEyl1Sc6NgWYu7NKb9xKy3PG8JWCz4paip4/E7EbzN6Fbg4p3lHjQOceiv
npWzWmWeK6JduMumrINgceekpMsQ+45zFrXfwOYvQrX/AgXnLZp55bokTfPnXbjP
S97rem+jWod3U8oOPhdfnw/q9qx0yvSz04u2nI0xeS7mxczmZDsanqDfpeLA8F3r
h5l37xCXME144DgkwYkPeUJD4CObvpkdFCfuArZIcQaJdnc2h/RDQG+RrKX6B0mW
t/qWDiT0fKztQ3uqMN9z7gqIjs7YaerXwOJcoP7kIiQvDoq0oCC9+QVPEPekUu87
bjnEXq1ey/tNI93wvgHXCIWj0CKcp8FOUarLNdWX6zVfj9VFXjuY7p1e8UAp3AC7
mWHChaWxa8YZ3BqWrCfG6sdRVwwvOLftWo1C3u/IDYaHyu0WOjThLM+VTLWqTxti
eKTHPgUUT1fK35N2f2yfpUI3H+nHqrJGJglYLduBC5cpZ2eKZir7Y0PEOAzSj0yL
hiJjxi/IZjvuc9eZzENgNkli1hR5mEGPz2BRCE9JDJgyU/MnwazhccGa6GSiGzmr
UuUxh6jKz9QqJHRJRhPvlLS26OfjZvpkDOi9+1jYBDRbf2UM83Iw6IPcqCZ3qVYe
GqycAVE6Tpy55JJ2YZY+vQGd42fMS0y7pGxzWzlygV2J+dX7nuMj3m/OV5xBWz1b
caZS4++Ngy1DoKlKzODeVwb6zV/Cc2RZzMqCzEdHc0vDOt5HnODAIMOHtM3f9VDw
0+OrFtAb1KuAQw2cREbTCfG2BDlHSlLMwzQ8vXa6WMBhxdIZG+Q0c8Ut2aEVC3D/
RdMkaJzEKRSuhkzYUlh97zdSHfLdxcrF32xl2MdyBjm76X7TM1gwuEyjCKNtRIHK
dgk3Iv8eBrXk0z4Nl5fq3zXKdXyn4Motlsgs+rOlpCf+jYZrHDaT+BUzKu5wR9II
A/98ZoAQ8VoYAYTypF4ROec+sVhe5QdPQDjBsGY6Ie1XJg3JUkR1h3hh4iemnqXH
jO0zgiLDOVWaNu0MvrS411EHfJyq/YAj8a01acbECiIfCueLIQkQCwNC1YwY6V5B
cdPcjVdH9RTIuDNGOicWGC4/oLmR7vgOHjRlhUjKsghD4y5sDYaPchAJjp4bvpa8
cmM8zaQh87YKQSUGxPRCxpMI2m1UqskdsZB86ZGIr6t08MLiUwEroFbuLIMcL5VM
ygJjDvRsX3i3YSw6W9xK2y4omWndhLsWLSXoCFWRcOjVPuDvuC9cIP8EnSh7P39n
9vXzPVHMpgGROwxxQHAbHiNH1ZyO936qD2U4uCah6RC7SA5yCi/Qc5decXt7JOe5
HX0I9UjM54qWsl/sBmIVsmlZSkh5VjoWTTKhaHUt/2L7drj+XO5JTa3dMKZqvfl3
km+KwHLrAgObXe5h4oJgaB5YHVAx2iGfDpLPHDz14KrNozVnbvcyln+8l6ad2sDf
KsOfNIRFubUnc4PnEueMwD36l7BPvn+sWxnJEX4i+mzt40l/NDMlXwdCjejNxQ2n
riZMipv4EsyMNiR9Z0naafPizXeAEGh/8ow4bIJJJSEshT5d5huvxa3hzTAIfZJl
Qc2j2swfns+NXEmoKv28q7Um+BWrn4jtU63Wa9WoVOtkI6P9pedFPcTPsuSTed08
jY61CpzgPVf9ivifIagMcoJzd2mMxNrJYwxVV9Uzyc11QnoOZO1ReLgd+4qCV7Rx
tfFF4UftO+LNl4liO1YDe8NW1EKbsKA2OzyYNvptHIME551G58NxF4Zg/sV18DTJ
goRJBuyiQY4NdMrpWS4JY6KGwtARc68z2blk8p73M/LPSk1z0jeby99lBDbbI2co
htyG+Nawjx6BplwHKiZ4O+QI4/b19NymIEGr1QBuRHs72bXy/V/D+398AuwOUK4e
LMqwUY+5RYli7IeSbX2+kyslziff08qoBotVlByHepwkO5KFLxFTMHpAYaM2BpWC
0HVANtUbfIQ6a+noOrYiGefgGpUR6vmOvOJdfFB18nWs5SYdtr0+xOE45DYh6f2L
7QvGWUaABUkrlo9PF+oEy0Pq202V58VGtflbxb6foWwMB+1RwB5YuJwTQIr0q2/q
hly0+uGGhrchl0wPMFJ1tmzuOs9sMD5cpI2J/jRa746P0BgiE41RiDtJdoB/ZRVZ
hEYowrFUvwD6g+VXRkw/i3Lda509+IbTkdYess4a/h8wwn4N7QPXRZuV6QjMaGoy
jN7aqA/eUDcUgeS/GxN6ZPt0NSVV7V3manM2jSnPBnOLMtUG8z+2gTFgFQYnDOrP
o7hGn4vXaSOF0TQZzq0HZRED+rbSx4P64Fg9F4A6AW8YB9fpp3Yk4CaFdwovgojo
2UcH2rn1BNyAvePTyPKB9bsne38ZljjA+psLyxYQ3Z8RcYVZtW1k8HvFR91hLFMK
6uxxYhVu0daCcdoEp3YuTguWbHhAqJjZ/0KeLSy+pO68fx4Xswo/xwOmUSFbYgTC
Ww4eCrVXLJZjH2HrHmIuReaY5Tpuw155A+tP8kRRN9GMhuxSWQkuOVJVnKAJK2CB
Rd7OX0bmZMTlA75aGsCZ1+4TWorUqx/j5GbEzqAhhUxjRCcyCnn/gWjfdzaqgJbM
qsOdO6dpmxt973cGKpFvIIv39YJaa7EMNKUkfByKmUAN1spAvVPa6y7Zts/hlzkD
G6rQI11hNbcevZuAqUwXq3p4LOCShzU3x5ajbszy4A4A9T8UhKVsdfb5cqiWLSqp
abB5LDS4HnoWNHnQJplM5gHh0FLgu5wrApaoF/uU6i/cMWZBs1scErcgFVwqNA+s
L/SvHkrtSmoLxcFP4VmyuP8K5ycY3ZlFls80LBubiBC+lc4nUw1k/dAKL8b/0XtG
EYYtMuBPnJN4ctnqRtqnMSVhsb9HFGbO0ck98Ym7Fx4/Bb7BGN22ckVOz4q/AXLE
3n7eYIaZliR54vspOcpEXeGgmXMgCvvMjNT2cJ/pw3Obj67kRliaKm8k/Y5+CEa6
4UQn2tXLy3JOh57GMmSVH8XGD5rbwoHdT0NZOtZhAvxvhLXf5jd4WKTYglQgG7OS
plTrf4D4JrucIPgC1sxp34YctOQaCjvKzl/lIXVId6vUsB40yT0tUQTywYAdHSWE
SLhgRaaM2Sdtg6o6teozZr7EZFhVtGEmPK68lKQvC/HZbjzm9bQ/srfHKPhPvaC2
ZXykF5cX7iOhzGt0hjX5cVMZ874rysq+vMZFbX0gDkY8/6oNtWPggHwzc7ZOCce9
IbmN5vl+T8poIUzt3rE+4I3VuP57aY5DOj+lltGftii3prqRBmjxEKnmsXd7Etdi
LWgHdIxtQzCewfKjweqAg6WJClGAbUlFV1quu5+PEWCT9GeQYF/MqVn7NF0L3Vey
6TNuFfx6br536Xiw2peyp3I64TstTXgvkwfJFYjBh7xUvdOQzHKUySfNI8UTJbAH
f8M6svJx0GD7hXQg6XwCfLS+kesN8s34668AyWANN2KvytnEGZHWCi09mlM6Gmey
hLSUXJ2hRA+Ap02JQ8t4FIdUZriTgxEHGBbKXn9PBgUlLzbSVemyGrdMccY01rav
W6qzgVkKqfMdYIYp3OM2EfgXa9l1pZXrVqsS6dwcQ5w8HiOuYQl/NUQFdTx4PlrY
4gNy3JY51rpy+DC6j4jDq8vhvkccI3/35LvJq+CZ9Jpxa209LVacpwl7ctQn0lW2
li7OCJECqUoVxTUvabXvfyaZ0KtfZ2cUzUO2+jTIU1aF18JmhFNRTTia2n1RRN8n
boessrt/oYrdSn7WccQMly2rEf6wQa7L9ou42MxfXiQMckVKZt+CVLniVOVICH0B
OQ0XRN+d/vNV9Q2nxZcTL6PwJfvGyCt5JFPkvNPFg0INHFu3xUxtqkE+Z73fVfA3
e4vhdreTyW8HwXnMzxRYiV5U7XRkRtUA00+ZZfI4iq/gf3/Oek6SqFzxcdfi7BuC
EvJSFzVBqx97zwsAw8hy1t7TXnt7IQ3END2rkcbxa8/AIvFmiGQrKKW5fq/XUxkh
cUY797x1fBTaUdfG8GwKTSn3CAu8e4KSGhp+8gVUOpvFtdKT7yV9IVg6vgxEvVPd
U+XTIEJceKvKywQYLH5dCsS80PL1New1WUGW+8fXfL2OvmAZjYREZnkM8W4Jll6H
Sol9/NnN7mZoUgSuxFr4nS7KXwLFGytYRYZvU2ITRkI73LHVhTaeEzg05u00EdTe
Qd/xciJFEfxTUzXmpE+ASbI8ydehlPY5lQhesHStkVL+B7a5DU1LfszJdGHSUUFe
ZgYUBVPfjAsHoMwgFwi53HY1/fs7beCrbPTgwJbhXP3OqcYPrn3tQ5qwJvinPSZZ
bcsch61Xd1E1VSFTyIyurufqS9696Hii/mW6sjNUfIBMfjwTDVwGUL3Uif2442An
77JASWaZCEZzjyg8ozNc/9ae/PwCtMjL60itNHe9lUPK0hG29zm8fj9v1abLQKMm
k2lOgwJxvvxkaXTstC0nDhVMbawvkGtYt54Ck+GA26lEtrSF1s5wI354Id9hxHZF
5UExEiBxDaz/H2fGQed0eknzNtp74q4kOOw1bqCX++pb/6dKIlpmFLvf6+3nzKyH
tcn8jytmE7sBAwz6l4Ud8HK/81Lu8l2ER7hWWZIehpxB53nedZSYWOIStkrJyCjh
gKgf0QoKT/Y7S682JT1P9B8HT2cuDUPidYI5tLEG/CEVElQTRxcZFdAwnmwlJzg5
I5cTK7j/nfFX4ZKni5NWgIZGa6pL4JWYTjc9G4CL1ssNx9bOC209Iej2TppAzJyZ
qUIEFBq8nOLdpHDXyn8vX6PIL+rWMBvzjQc5v1ZdVEzgaV6vahDNLO9qm64h6oRS
R49+9s9Z5tWQXGGAG42CFuJymfHOZ2L2G/D2q/e6ejF1dwvptjsR+Lv3OSlAyliM
lQx3ShSgwvjz54OzmhHfxhK0nAI2etma0AnCaGvBfkdfD5ezLUF4HI01gIWyrAbf
1EptBjiwlUtZTnSy5fATQQlF1IP6HzIl0yn2NDEG1Ai133zJiofVscsMsYk5xStX
dcoHr8unFMeVX4Ij9fbuhdbuE/02lxZbrJ4prBKgAxdUELmX4mrBPfHqMR0JzvVM
eldtKTKz/FQPTH5C2JTHaet0cUg8YdygAtqARQ4/4a9Bt9YhtTj03B/AvriGlSuz
VFNsQu/1lK+Aj+lJxD3VpY+AoR+SQSlXMh1ikvf5CFHix8aj5a8q5WPhILDdGY3b
8qmFZNn3ZqQjVte2mXvdiZhg6D3pHrnwbIVURfsk1LzIBQJDD7j4NMtXSHXzdhIO
RfzO5j4PTdoA2yU+M/fPqTpj7cHL3QJu9IuWFP3k1hqA+euZc4DeWrL0+FoDfP4E
PoW2h3ppiK1sm54qWHPB7mfsgFx5YP/2HV2Eo4jomgGOtGxh8/zFb+aAHumX+LOK
m60mZCSZK+fcnSJ9fgxvBdwkIlC7RfwTwulp3R6G7jYK3N/KPI6ML9oZj2YEoCzB
UYtm8nlaDkkkcBIURKxX3/BzXPHpEfHYgGZp+Ww7VWOwIACq+VO9o5IBHPqSlc7Y
bQorIrR6RKUdU9EMu8k7VGHT8LSv7j1gidbbanrS97rdP+AzQFzl9tn29KKGE9M9
8jzs+kApr7XCBtYkzm2xYpqRkFnhlrF30QC8JrwjG+t0juAJThiiVZYQnPYiHjJj
KdzPE5pe2rYai9VY9EobXRo+DnP1Df8Qb4eDKy4C7K795t2RkV40J3RpZu+72Anf
rFynSRiSKWWxaMUayVX2Op2wXuqGUQRbttMwxbwEFxjCf7xAGJjJ1fgoRxqPHp1O
agTuCO9MgD3fwzaFfI268wnFd/jKhyIyLnNJgjSoRcUElwRh+0boM8KrCLo0SlrI
g2nnYW0rvJhk7itA9bxkZYvfSH9Wk9RxZuuMx9u0YLxx3xDDxSMjQbD8Qd/iYQlV
18LWU0Z5LTZJKFmbyXuMbUfiZf3NomLOUADE13DP3Vc6fUwOIyTZ2PQrxKbisRqc
mtBo60bzHplPoyzeQjmVN1Ue9u2fsOis67mTAfY484hbRXOfgFuxPvb01ysnAdcP
vEpzVvurrflvp2889+8YKS7E3tsTyA4p3luJGP/V4wT21B30NYZIlSp55GTwA0Me
o5c6QLXmmjpZ9RZh86UjUeBc1kezk7AE1L4UzsKtVMsmsE/AfHuQfGNPUmwS79DP
sBbsMIq8MqE342q1biQnF17sW6Ww61Ev5l4WJ1FI8TKR1OBC6/xhJFBbJNtkgfNK
q0teFhiE6CbIM/qY+n+fVDboHIxGnjNuL6d8DJmCeWpjrcx843CNfASS3Y4tFd5J
aIuHpQN49YLhqyJowmvpZtCaN9gyro5ZfJpHB+yB5kzmUjGtVBz9afD96bmwM6dE
/DhJqahudfd9VoIvgbRXIEtgIANGWQhUTIvWuKTfLd1HUs80Gf2cKuF/9V2xGHKI
VD8w/PqmHTUCLyKofXhT8RedFOWCMt/pCVD8ePYxUOUQYWDefn5VQGCXTMEnqXr4
/hyT18Oo3uVBBqbqSEPclVd6rKZzxMkLul65pDIBpO3S1VYcJnxAD6RklDKcuZI2
j24TbqeXctFZCw9wtRSd0+cS05FoX2nlDaIkcPGjvjhJwsDIFP3CXtoz9b1fYH7G
0AE1tktiMyPaC/RS7O1asPeJC+R0q6BlQN6XH3XweeA7sAIzNUAq/XGnaVkJOj2N
T3TIcGiegwRNOKIeqaFyyakvRhn1npguPgGMVcBvwpn9fzv/luk4o4hGBVQ2yLcN
0d9Os+FsMquEgcYpWZQVq8stY0FhWQSsM1+BRMfjZ2uneJbtUGI85C5Z9C3XaeqA
f5nxJuwvvNPR3gTGQgTXvJ9GLVSKHQ1gShWu9ElQqj5JNUjBuxCMUfyBx8lJ0bmo
vFqJJfTIoqvoGFBp2Ujp0seJ3tTREvWk12+OQtuZfD/8ZsW/5p70XvJpmMJ4A0Dh
u52exKqNf0VFV4PrskpHN33HIZ927E5iySRJIpXZfU59ElNlX8xoBok7Nw9M7kKc
Xyclo2GJnSKamwGNdx/C9qwr7Y4teMvK1AJ1yxsgSleQ/4xFkeck+nsGRWfyYrnE
+6DslnkMs0k6fhZqoSWb9zZ9y0TbSPkuLE+/ah9jUbvxV99wgeCKQVu1YOF/rnyI
q0m0CYjT25cyp61+T8WswZ35oD6ln8Pk+EFdhtP0qfaY4sROa2hplSSwjzwj70+g
XqwyXGOqgT8raO2gzPFIqBiNWQbo/lr28KZUSd4soQbOyahuYs1q2+xDcSwpy3uR
b5/6HByxwTEIl03wdkw1Za3tp4qcv/KgbVmM/E8q7tFSvD77ZtPdUwYUT5h2vfJv
6TaIsGD/3unb1qJk3lczqB2iu3t28tceAWvHj+aNVZLCg9kqZPv/HyqS810ADu4c
S3vUMphqci8FYlTAU2i4MyMkXo2ywGZ1YgpV942cjGYGbP3Bio61H3s0uUCUbCQQ
r5XK0oam0TY+cNWnAJwjCQbG9FBNwZXIFmNiptPndEeDfKTrY2bGvxezs4Y/OBNT
DNmijO2bkoePmWzaEyxY4gOdTQvYP469AG5rYdn6Uml09wdJDcGMNhS1tGcfxPoF
XdBExCrCJugFmkvucYxvfUc91p/wTH0mixq/PKHrtlsdzKGKL11qaKCpjssbjGmG
B9D85+T49jaQFw29/e8MVmYsjMtxPIqpHT/8prWZ/FTKxovUWejzMDQ8cCsCiRgf
ArftJz/FOMUHR7r2atvoqISscNQRVKnPAJ2fsOTXcNrxy9sVaPwqeTnNXgO+vhwp
gKLq3kLFEBVaNZq+ti9z4pnVm7o6iiD07SCJds0w0JtJH9zqfd2Ppez0xYXT+Mzo
HZLKooC0cRx8Lh3vcLXeNp0/4+JD0TqPX9gtJFzsNlnaXNJTRiHMozCla598h2QT
GBUynmGyiliX347r4i7tC2J7onsow3BDRtDJ0eIzjGcwvdsdj4l7QKUWBTjkmZp1
iggzT++ncoTpq3UREWy5BRARbieZhpbn8Xzt9Q3nphptKLmhTibZ4BM+btztV+mw
uGnJ3KcDw4PJMelkvtgYJzpxzyDv/77RHZRSzgy6LehQMyg7OXEX1iwD7R3Sj8Mw
EhaVChAubF2IALuawOXjjU4qhYtVIDE/UqmWeFkTheibZmUF3pbnJzzsx4pOoTp9
lIIn90oa0ELK9KYj3zCXfN2Tnm1idtngvKMx/k6vnHMlfpNMhOy6t61LS6mioSA7
T8iOFtXi7hJ1Eq9VNSpX0jDNCPWwLkVsm2/eCLJ5WXWN4qblaXwMLSQeRfq8WKsn
tvoTiQxJqmQLvr6bBY9tFf8uXP9tdKimzrrj4kDBDJVGVFyoIJHl47V1YXQcjM9h
RG4iN0/C5mNO9g1SKf17xknNJo7QXjC/kyyp0vOUJmJ0r1Nf6y2BvKIjBWe7HJfl
XABw0YShUey3JclsIHwKiouyiadJWBTthoNXWWjobR4AVdMokYe5vfmNyLEUVCEH
JdiB8+iTiWI8UgnP4+QCmhQx91Okka72jp71mGcnZuyW26HpsweFkPCnFOh85/2Z
mDGgXGf9DCZNjaXa/joUP0toyoIVWEcoLfWySeQ2eq80D5HIeaprdN8jp7HVvg2x
uiFt4Z5uX2BBtzEVgwWVc+NzxJcVCMzb/jqSm0XmuUq8kHsvaBydXrbBZURs4YoO
OqFKumBo0Q9iLVB3zufMQXtgWt9IQU2Cq5pxZwf19TJQAFwQbTvQRhp/bZBb75LB
y3y4NFjruXQJUJ2b8QzvaI3c8MqakUqk2Xw5CmYA651ewL2/yvk0es1zo19r4hVL
Q9Lmtnc8OFa+sfXFMYP+PohPLrGXt+cSVXMV4/qD4lP56hWvpYwsWDTvPFW9DNbD
8jUEYjXYiDx+ah1RFHiOnxGu2uCjIwQTnwqc6PTim9403TW8hKQgQKkutDqhXWmy
jfckni/BLcRT7QMB/1KdDt0/HVF8AsvJDe+kFQgPTxIHErQaRckzuF+WG0Q1SYah
aZfMahraXvALEuqSLBAYdQzjEJQ59Sp4B0jhL3Yij2CUmymIpBBuRYDGCMKXFNdX
ZTOWW55+4g7tVaMea3FEX59DFnHQXnaTr5lOQb3K0zbCs5UIElXyK76zf/2wywsY
WgnXXSqUOC0PVJP7XEtxvnMoaBgn+lkt2wyEgv+UDwBEnafObAbBzcy96Gveq2qO
u17UXQdw5n3GID+gflwQhFvm02AlA5zfOaHdL3FONgoNpmcFPIBAzKSVGJULBDHz
8d8qyjuzaWsUN7ysix+koQPzU2KjNX9YxQW7wHLsVL8MX60k08Fu418HReO94EPt
749snbyjDXMDkn+30hl5zbb/3lmYTK8gMm4/KDMGn9GV0nXY+W1BlKnMGk5eW2Yv
0PD3lifMlJAGmaBxanmdgGYlbKIzZzGb3ornPqtZbwGgcHze3JZbu50JGp/C/RTW
2oWjEGuHDXElbCbZJY51l44IHtZnLVHjtp28HNsiRNy4sypKgh13OSnZQwczyqKz
yVu1CNlBmSRlF2iQHY6TeQ9zZSK265ZVrq+zymz3i/p58wKRo5mFF5GnMslOP3JQ
uV5JnUef6kyz30jFubd0IvTqym9IqA6esT8SwwhZfE7vFu9GIWuUyaTaGMPggaA7
8LafzWJoM63kLYapFZNEJZBauO/tmbQjpmI3CnLA6O/+QoMN+JYK81kD48Axg0az
0Qo9oKLD7DKxU1QkvxlzUXnQ76FFhD5ozsfLfOTvk6XYzBBIAW0Ap4ua3pinAeTA
o7MoUpOJRRMEJ4OacWZpOmSXwbMaa3YYRSbILPyQVPIYoFJJshARtN5HdC3CH6zn
pmCqIi2YLyUNfUWW4gjGImFZmgdAXMbTovpKJgRvKQHWy79EoTLDG/cC+XOzqC29
Aeb0LHalaI/wx7kQK2E/S7tczaOKQ/jobwVaV+x/mjosGm1Uc/oglDGCNtgZHZh6
tFvBm2s30WlZ/nRCPT1Glw6R2ktAbi3U6G0PM2o0bVXtTe+q/4KB4pMcmyuSAN+u
32hTQIMgmS6Nfm6py/REq9cYKm7Vy3qqYi2uG/ZcqPuuzD90sOYnU7BILaUnJasS
NhohkdrR0K/F0sx09vV56KE+Z6TJ/s8ukVxrsn5dT7AFWqBGKfvmPKYNQGvb7c2E
LHEDBIYf76OHWxk+UfC8kNsC/2VMsytzDThkIEdju8Ugurw38kHIfVU3cQXCVJWk
kpQ9DsU25YsKVCfEO1q96/3YRJ7TtWPIi/n1iQ12/UDuRxvXx6QHo89r6jf8ukiw
T+uOdzar+mULiSdF6NT3KF2Nea6d3T6/fkURLpjd3MzWrVi9oxyKU7cDGSiwFLE5
KAe78n6Gk7znmPebHl+3fXfIUamvfj82TERtsOdVoDUfq5VFaUchuguLhC5ih51X
sa98yPW6Rfsvv3fmilc6Tq4BT7IcxxsghFIkMdilXVhJCC+fvhHjQ3aT7p8Hm0tA
fufD8ly0ZdHdQ5IIxyLGq57edH1mJBRYC5uhQ/IpwiVNxDnOAAcwShyHKKL2TRiS
2MeRUfr+Uv0MAEVIhV2fZ4k9vnBCKIVYB+/1sXoXYzq+Q9XNqiKAWiJc5C5EODQ4
pAxWgeQ5mAcghmm4kDl7BcPXLUnJcX7OQuXZ2ZKdjBfXPYuNFo/orR+/mBOX1TJK
H+MvF5va86lYNTy0Ec2cy+WURrlEuF50dnBooyahRjL3zQp+tFhqa1uC5RQBMRkG
U/wK4KtJuf8mkmQ/NLBT/DSK9krY5t3mJ6kSEwnQ26s4B5LZSuukMhcAY8Z+HAWS
QJ2WfhbOX0Ta99WH85BRF7FHUb4VlAQv3jK7/A/dHJtZbLkxw3fTKAwHz7q70ONC
toOu7t6PGnuRuA+0QrQi6RHPpQvzkn6/w8wd1T3G0pqEaz+bZLwOFn+Fp6aZtPkD
gdcUBht714U4xRYe5SRxmNSvqsdGHrmIIfb8jzEP8E7bAMSkanHS50QxYRRZIgbZ
TgKocvksmcZrzwVrs/bK4VdtOdcRSl4Pgj17i/mgzo5tbKWsb9hblmcbc2DXk2y/
dP73aS7VhFZqM01Mfsgry4Ynivj9ubTk8Z6cSn+9oguOKsnY45Xkh5vSQwUGAbxb
wuxy7O9kiG/5hB7CkAlUfj7JW/5u3l5ISb34hWcHAHohSL76wqYUjyctBGI25wyj
VxiAB2TebRaVc36uftfe7Iyg94klBw+dUqsbz/TxNhsVDrAH81rESyG9cvIbKX6C
qwPty8vnOOSVM870ODC6fCoEXsA5qkP55V3Z2MS4O7gCAFZlZ0K/x/PaCyMC2A9x
31Hg4NXYkB7cwzaou6CYFUNHdunvzE1HSS+8EV3CdkabJ0h2kDKq/H72iHTmLVcD
cGHlfR+4XO3kVpq6PQkhSCC8JRlU1hfMWarEvPnz3fbn5BOZuAJRl5Q4fHaRpY7T
qibwRK5UgHVlWUEHD5wQosyu4OGgM04/T9n13XCxTHj+W0Ht3GIXqlqipKW11Iuu
YDETPUrc023U2jlHtIwbNJ0+JxdeMm5zsc+GzeDM+HbodNpUk54du2VimpV8kqf5
tk10ca87n2JQtys/lfocm1fSRV5L0ZnN6mbKzSaiVGvCV4pQa2RwiNSrpR8TzqMo
O/Yrw9VO9VCuyCjr49cOHgOkPmU/9I1oPDT2Ef8kDgi3QR8cxzeA5Aih//aYj8Uu
WZRb+xXD37wZsJHuXB/c9Na9laE9TeE9jTj4fFDLkyQpJrZeTeigxuliXtRiSZqt
TsZeiyjnU7HYA/Y9WH9p7tY4KCndo4gCLsQZ/iV4TZPt1H8K8MJWXfg7zIn90fJI
iZzh2rc7J/2of/TEjduPiNzi5cUwCfIQduO/DR83KX6bwtsBLfiZasUTkVmUJxMo
bdjweJMAG0d1Fe4Ja/iCdZr+8w6svos4wk4FM+MZPgvrwuhHmRvPdgwVHUW4rP2H
+s+oXjWpuP8xlp28mx/Sqj5VAlUzwOVJ+HhktP7LZ3tcqChc2gXPxpvCc6x1aa2r
VZIsEirypOeiZzMLbchk6ajb69YcwdPzCycmr3FCRjoOCe4HAgJCm2BRJD77iHDj
+wFFp/9OrK217FmLW8pZeqSwpacNdizEJ59D+dYqGb+USaf69+l5JYexzeXcTgOP
JShxz8ja1/N7/+zN/he1YpjjF16/CHFa2NY/w365WO384UzYFPFmCVVMnYSpCGQ1
LXwzfpjfDGMN1/tqTmAM5SErZfo70+mYzKn33vC0txwvK0o1qJ9RDLtalbJm+He3
kVjfpNXaylE4lUebiO9buVSdIKplmcupTDJtNJbZRdWn3LAcUgoJajfLsM1Fs2ar
rPRM6jDjikvsxUG9HF13+CEq3ul2f96afY59Z9zPFC+qDnQs8bZZVecH98mNd4Xr
dpXtNRtxEz1qeTdDkNmFXiBK8djfzCWlxpUcWvUEePdREEw8gjbB3ZnH8sdcjaqa
mvMTDwW0j9WA48FImt533ZuvIU+Zz8rk7useNuNiStQjlDCsD27nXgLqivUCS+wb
EoOXEwJIHk9O5KIfvd8207IdS2XDj3mwJEJpkWtOSvKSOZgB4hjpLJUpwonAgHqB
XBiwtc8++WFytBmqg4QsrxrxJFwofxnVFa8U1zePOLVMxq82NuzeDLzlIq+Tk7vg
ITlbnFFR0saGobyH/J8LypL+2u9yJTWNOH+apmRGsyZ/sCRrFmD6B7+ahp6vOyd5
9pe6wikoCJDVKE8qTKZRL47MuVQmcwlHmjs2TQSVgNP5pI7Hc2gdn2phEEBv5S4O
rhH8O2rln+VkcWon9oeDT38H1+utsgjcdkMVCQHC4vPe9Q65QYDFC++Hgfzb68rx
wK158jz78Gn4wkGhU80D+yTZPI0rQkNSSSP/3w3LobHyP3wcGH2dPvI08/Giqg0m
+iKTdlJ5XyVjb5FUA4jxDWAh05KVtn6XFug4fxGrr7rN9JY8bYe8vaT2nQII5Xfv
tBWGe5xQlgAYawebQMJZFzQReKsk5kCWCzFY8+0pVmToa2C/kW1LFQwf84NiFrGg
tYFp12YBWKu4BsPfvob8JvQYdYAc+6qTm5fYjwBwSeINETe8d5jU+grQlSV6wf0N
1WeBUzZzeuUVwX1iv7MMUoTC19VRWBKj85QwNziV8WfjzFNEYFWybGYugLoSIrcF
bG/1Lhr2rme5amFDJxIgDVDAC2wuuvH4WNBzhOyP5Wq/anFGQvbooN7JY0KSpSEm
6laC9iw7HxXZHXU3QAGZj//tXIW5YkewYPiaCfjiHOTE/38WKinE3LHEp4Wrr+xY
LrgiD0HS7xd/wmMKz5UXJlfRiyW6PeqA4OHTw1O9SnmFUb5ccr/3OmMvPDIu3a19
hmEtod7q+tH1MDFcYXFlbqUDEGLtw9yHqYOqLK+8XNdyUY/vV2Ri8PrDeDXmPqiz
l9IqnSLKgYECFFlH1l4R3qGUXGMd3RcHaxMBM32sjf/VzggLn0DwgiF7F4Q1Ozv6
M/B8NRfMlgxE1x+HZHdPy5wsuoD1U7bdF4mDSn+ijfT8xC7CAsH1Kc5rvacP/ses
bqzUxcfgJYtWJBYRzw6MQcIkcWHqb9ADNk8gYRc1FLh4xsd2FaRAyBCz+y8D++m0
Kb99A4gCMMzx73JPH+t278ppUYRZJpwFE8pIjoWowWK2/u+kIXwqE8/5sIGOZJkg
5biNk22IO01H+jI+Cwg+++TpQ1RYldBvlPZ6O2Qykj85tKuTGKW/IO1HbqzLFe00
P0qsywNx6IR1uKayIiqTwN7XEEXaOpD900pYBlLyzvFsEjv329nqbxHENxwq+bUp
uG0ap2f0SzfSHvI7pTPaGVqin6Fd5z8rWWUpIQQ0hxVRnE9kX1nDgb5aho1X56HU
lrwpQ/uKXJ/QJDMR+ua52dK9b2QKFx2wGdShnV0G/Ipdgvo0c+OPw2ifjw+UBiIz
rBWObjTnh3CJ/vzi9ZRMgFOb1RyuOQLdcOH+mjot+BryfwkhF7Fre7rogHafba0X
/BU5rqFGWqsM9/HT1ZJ1u0O7b4rkmv6qqI9G9nzHjqOpwIiA0Y5kTPbaGaPPDrq7
UmfyB6wi1P8i5CSoL2dPUxzIZq+XqmKKzxga/+9D9loXycOwDWEzBHGEPb0Y67DG
9VubeTUdh0n6V26TuVT5KKFHUUYu4d7BxoYI58+KutyEZzHhMwxaAxloMUkIK+jk
C89RaLxx8G+gBD8g0FF3H8EWtlEMU0aa0rnqIIO5L9wouLwoOGUUVmiyGLgJPM0D
MvfWLiu65NeDQ5CSMDOCjEDAyVyPlJStuTtZSKLyH1GOV+tYq7bv0mpauO6EbxrE
c5yCfAZoKLFAXVFgyoHypms1SyCq9KJ674Rgdo69eU4IqRMP/dpppfN8YekFRleK
oZPYv4/BRzoXALuTMRIkmaVtP4l8sDw8IDdN6baHSXVHXuXxDuBiZ/2PLTulhMCf
seiiJH2LEhAbqb3cIFa10rIO0+IHA9R2D2piBcOwYC7lfYp7EMX79tknTI4APkWr
ZpCVeuTsyEyhGf0M+WXJv5xI98AXUySq0Nu1oZcNVE+edm0ViP1W9kcDcO8E5Ndy
x56qxVPuHUQMRIghsQVd980pIsP+gYbyMijlC6KGSa+aU9wdhtYc82xdHX05KhvC
kTFxoNo/DJCEgMpJULw7+hKBXSmqnDIDbaBjOWptHgOlrHMuE2Jf/cs8dJrH2nYA
9/JEll8LzC9xp2+7HV3jzR9F4IT+lF5Y3rVbaYQQhz7twgz+RBgf8UWNRo6FLego
w+3JyajyHLabP2S37RUnI2vUT9S66iA3IGL5AGZE6pvNQOFJ9E45i75zX6ouKZrV
s/3VarRkAD63q2vALfGRirSxPWByXb8e02FbiaECcXN1/AH7D46rKqQYyWNp19EE
VDcb7F1ZMau97MdDPRXuZszo2tKtqnFev9PdcBCrwhlM08Fir6vySW4WtrvwCmNl
6gghaukLozxXc2SlhTJgnDRiip3H/FQmim0sOeCjDmAJdBJDqKdUZVRWlD+rt5Z/
o3UbV9+BIF/FQUA29AhJdUhjt2SVFuCd0nq9WFeWH7ThXWpYh8dAr9TkVHi53BNS
HDIaLRi3u8AlBe0R0Dp6zcnGLFGIs+B6yT+yAA5HWOU11G8oPFvzi4na6D04I72U
bqRfbCKZYd+bsx/pRtVEH+Jj9E4l1qY1NMsfSOS56jA86mJyxqgiOseLpXQ0nCPq
KrsPgMkHel4YqGTP5J2GC6IjOqWsjopCu2/cKz4BBsWZY6nn7ZeCBfFdLtHBgwE9
sTkvI16qay+cbuaZILRVLNQGro2Xk9XecYIBaVx9oD6xI8o7K/MUpYwxlhTPcQa/
5x6tKH4VxySswyA2vx521lPDZxdQ5l0uhrvjNh+clbqwYmdR/KO/fyI3s3uomWhv
1zZZ+6/A8QvH/DuhJLEzzKzSJ4LO5okjbcPQepzPnIJNko5YRx7+0saWXBDVAn9c
H73hErZEzjg6Z3hFwmmD3X1EBALvkLPSgUrf04VVt6S2anSbnycIvhm/v65ANGrd
Uev6JWL5p8l019t8H/wBx6q9Ik5vi8IDqpJW2sKy21rFZKF8ssH/yjhT2OSXqiF4
mXVxBZji6OsP6m9frLp7WU7STmUtT5h9XXD0dVRRNlCrCU9uS7GcKrIvLh2I2WhC
0OsDHJnWKOD4Qw5wSFiUNErvECUINGChYs3Y19fH9ol8Iv0EKDXHBAsaDF/ZGeVt
w2puItKwuBR8Fkx3bygNIexHhcqEc7t2w/5nGfYdqcCc3eVXPZHKkNPGQNMCOnhA
tgS9iUw6sqXsCszmCSfCXYBGGPKMWR0ywBGFIoj4jIlz/PopkTLmAtgCCV+T8qU/
3TXnK4qVkqU2O3kmS8eF8fNVLfEuOcTcW+9ib81tr349jySKQvzhs7oYwiQy8J6r
JJmDVCPrliw91VyQrjeBB+bOsqeRn2j7Q397klL2uyvywtDBkxWfX7sKH478UCix
vuK1lsPyUF4yD/eOq+ArjroOFP/1Ct5eRqVdWzJXRGxwZIXgaJlK9HozB73R1KxC
rn7A//DfixXQNEPE2M8zjdV1Q4OePr1dEEhdHKlJ3v1lYwzGQTItXQ+3NMaNdrMU
w43ZY3nBrVA9DljpvlQv0xLsdPn4ygeWsfLywLLlRuUJM6pjIbPyGSj1Dbcpl2Sf
FwMhXUeTVWGd/LzOV4GKYN/kpru+upD+spwWQxy5NtIPuZnvPYtBV2E+rZXddk3P
DfHyQDKe3BUXjCTt3EJkClOBbmEzf9z3nlLzpli7YDnOFeVqlDHB5gV/WbCgqgpL
0jl+Dzv6JCZy7HMGmYrwh0KvzQslzIXvj6eRl3dD1ZvodS/12RqilyY85a7psF1s
x/j+Z5w4QkVimYzQtlykeGLGrHzb8+SxwXclZp+ooZb9UqkY4IdvKty2N8+tQ+sT
YMkJ1yVFXA58kFTmGI9SFUUhWtoXtibdcoOqi5bYr+Wht09yjC/D3MehiTxIjQQ8
VH7gp7xd150HeKWkNC2ul9XDmN7KVoYcBXxjCAFS/AmroekhBFU6O5BRYxjK7+D7
qtF6CIQjO+IMyNrrZissJ3mItLKpTJbPqigunKgz2ZRutA0ScOraQ4B8zmTh0egR
s5qK0G7yh9gL2YgvyuTcHxDc7gLOplcNo7zJ/iSWRtOz2k5Ucu7m7E6zDduEEEWI
yfqRO00ylQFHgnMY8/HZBFFOrtXLPj45FECUf7+USBxu6Q0Qc/ilLYfCcZeZIAZi
FclgFnv/c7414aUUKOrm1n8CDxJMdU72E62zNbXuaMuKLeMeKR0qVQmYzV6uSYQI
UjaFIFrRpURx6d65Llf1AgPsUXz6LNrRU2ZFggZDmuJRBJm4HRIwDgtJkjNpX02c
nVa38TFjanaSaYLYPW0Y/xJhDjmrZ639dZlEwizMv8v5AvqgQluxMVBbvItB3yRX
S2ITVlrE5bZ26cdKYylE0WGdtWC+fbPM7eFmcABjUb9QtnaQ5NZH/LADbKfjvMHy
uNPlYlDcNSykEP8qEhJCwYMvwbkqaI0vB9PIRJzQ+g0H+TbogZMko4wKv6tRuJyA
QRlphQpdTykOIPZro2gy3aw+dEWgeCjhld5rTctQC0GuHRVRL+O4v/Y8gxtu0NLE
82zgQcThw7bC+bOGm9ud65Ybjh2+iDO8xF2rLJ+s+SKLOBeC0JJKKqUqnkAEaMt3
+nxHkw+QX3z2gL4fZBR9T1yyLnc9Lh+l+x9So4rlWwpUcyJfuN2bzQCPI7nhgkgD
UvpzHGrnvB1+cbN+CU2xbyBCpErKV3S7ws0pVZRM0vD0o849HeaiQdLKDdy9qpO9
ozFNkngIaGoXMhMDFj7KDSLfE3GuIEcAAMOx4pf4AtgDOaTMFpA/9hUncT1gTI00
ZVK5fsMjVlNm7+ilA5rffVOIkGC/YI5gfO9xNix6z/U6IIzPyBGGjijVvUAaKkt9
wCPIpCjY1jtXLV1GdOSR3d8pPzvC5qldYit95auprieJXZYjVngOXm8UkH5CFpbw
RiEff0xoztlfPdvt+8ragjeoGEORMTIZsqr+d86izhggYHlPz8Ikc7tSghHiKVUB
n1+tz246Tm6B/8xl7XnkcBky933vRG6KXuYW20MYY58xe+gmYE9JjYOAW8OJRDV/
oUZ1bZ3NOB5fBFvIem0aoswdHwKncbCmezhD2cSP1sKVLTR+wkpXmvRiC60zcVMj
gXGxavIcTtV+6OYxWOqkddlEbI1lQo4VKyZgzl7cNeU3naxHx2RYBZmsj5jUFuTq
dqRkQ/ne1x58U0+f3VfJt/8ejfXZAkU2w5OwwCn1SLlc71kcR9MCTDIm9SX10sP5
SzhWfyDjeXD9LrIM2QrNoTHJsB8qrAvlSSv5XRjjhDYq2kMqCQtGQVVm5YMNHewa
spBmXVVn1qx3VylEcdwEa7I/nyYeEB9BOW3bbXETVf4iOx48xzX/a/ccFhGsaOQ+
pTT2Daqwsq50CSMyOW66Ar3pBBh5LbvsGKQRFKzMnbENG0A8fcqr+0hbto627hel
KPv3VmVHPtk9Z5THW29KGLe0PIAfhA8JzvK/bv3HtiLGGbuzJSKZRj5OoitCmUg/
YYdZqxhcnQ/6YPlsKTZ45hY0jDixmv8dON6IED5vO2zykVEcKBIGMPdNoChQBYIe
74da3aqYAvX6aD/FAQ3lYffjbJpkX3K1o8ggz2iQYc7RStGlQOVEWpZYC2d0dw4O
8L8+7xA9biG4kY1VZKFT3Cbn4B3m2+nhPKHZWy3YEmjrTeq6beewy9QhRShTDH98
+SB0cv0fkVcJ9B1I30AIE019j6WslJvHxbcR9TCitJRjd8CAkSZGlMehQDDt/xvu
UOd3q0+CJElXHvRC+npXKxBwNjgh7EFRgMsEWZkTB3dTyF41lHBzUhlTDLMex2Yy
fdCXw35rXaNFhHlgQse1o9jeS9tXZIlQ/mrZ5iHJGgdkh+c8swDqvqhl00Z7eM0j
C1RnmHzIj13cbeY85gtsXSA7pxz1KSskoYCmY+fw2H+S6jkykNOrE1rcZ9OAcezY
78u4mnLuo4UBkt6rGgcrJm7u7bFmBsnFFEM7y3GlUPdOu1sjedNf0xRje6r60Hdr
oRk7F3uB9IapfFXWQFDac7+yadsw1xSuA/6LRZktD8ORFMnGQECX/kPJT4m9tpfu
8+YuRmifuGZ7+ivQfhOfAfLisy/GHYKUwgRdU7exBkItfEkyRVk4AhE1hA+XFV3M
rsMM8nUdxq3nwZVNn3g3Ug3PUoeo3+LwAPjmUyAGr4qrBK9tLKjni+tKzKVrZbLT
gkBfuOTxzCrIvtgyP5/13y0nTlUuawfJ6mCJqveQKOQSx6B7csTGSjEGoZduQhwB
M2FQeN3MUnLnUmZ/PkvEyo+gvSlAc9hlnpGfmNbQsyz/Z4eS2r5u2SfBYHwD/eqC
pl1kAU3igBpviF/hvH5G8xLG/4KLDKwRHRpxl5BOgKJqQdl/60sDyOPO2H4n79bo
BsATfEjvVOGXIPUvN41rd+YwfA4BUo/kb01byf0gJQLuJug9RL9uRf/iCJkjg4qm
c/oc8QywI6YBjcp8+VcBalmwoQ4auQiFHWKVXYveUnNqxZfpk3CmpOjKH60dmHTU
xEtlP36v3GDTR8Vj3otla+8eSnIbX6Ab4gy5pGRprxIsRO8UdtM3Jad6sKO/OnFx
ZeNkr65dztHAsFy+A2ig7t2Jo4VJOq6aLYTIXKW1VaVZkugEPpD5kXl6ZZJ1ndd1
VRTQj1aW3YmXCPuMqCZJ+EF3wFKcs8HI3/OX/NsG37LBa3jv+IPAFsMrLUtOsFRk
zXVxNBgkRKiu+NX9SZDVnID71essF0U0mdg9KmJLrTqJ5IYAyGxz3Ni+yMjwUj/P
LKstT0CIh7FPaHdeiwpktNsAgR4DsxdBlZNEYNWJMMuZ1duK6h5fJt4yE41oOFCY
MfD34Q/HAOqCX/0qXIz9h4PZ7fUQvyE4/lANIUruraP7+3r8+txgMG/mG/7YpBJ9
ed+cPokFuVg+jibaFWAFdJL08hC18U5yyFVke09jNR4fh91LTGhNlTCflm8DTP0P
7L4l+9UQudSn9FKQuNQY+dtgTU3Ot7y82r8qCSM0SCRiy6falL7wzNk6hhFpX0jB
qxxvKjDI7PgM0IijVrZcGsstvX8q2cLIa2pdCwqQ7/RZTCgQ+H9ZquUAb2tFN6J8
gADgSpuB2ZoWHiF4wKzVLq3hXlSHxZCFJ13UaFNP9GIuNb+b1hzT93htkfl07T5v
n2uCG4khtmZwFYMewaW5PGdIRt7ow9hciIWJaigHDHwtsiYndYF2VZrvuhfkJgZs
kHsfYaQBwHFpO10XdjSc34fQ2L3TVHgWSI8TCQ92xNncv1e3YfF3PHiR/X7mX/LG
rUp/f8QB3E0Zby/LKCvV3r0nmlXz57ETkW9oFXwg6vxwjDFpBb2VYbLfNAG9Einu
0+0Xg399SOSuWItwSpBHGyyN26XnKMs5ZVHJOoiUEPNpd8vOOT/Pt/+lJKJjaLtC
ypO8YgfvCHobSyRDox63HKDchGWgHrMWvOFYquMj5r61H9aExnhesPXcX+8wG1p8
ZaBc3kjhwVABH9JuErIQ3H3qkpxo2m0r3cJ9aj2GVj4KF4TFOTBogoABxnmRkY+k
rp7idy/6CMhtBa/XZjGHQafEZ1sxwvvDt5/4sheE1QLKwhbv31pjeGiAG9bEb1SL
3xiR7JuYGV3FVztrwpYb5qw3TOWWkJ4kRvuso4Fl0f3TBVRpfoJQgy6fUpHpAJiG
x1Fq0TDEW/c0/lLYnWY03/5a0jmi1W/99nyQdInmmYmHQ0hc0NX56hx0S27JD1mR
tHr9XDHveRvdp7jp+Z2QKcOvLw7k4JZbr62Tix5WD+6bF06wowi0HOhi817IolAJ
c2ipSfhcT7CHHohWSTKemlrujKR1uXIL0XzQx0t7dT9WyxBkYJvzrOZVwPhvw52P
9+WHl03lUAG3IGmobG/4hkNXwq8hQv3ps00MgOVDIIcbGhL/LIn4xTRV5KELZgsM
gejbxd4M/C5zwJWCq5ECOwhmaOsXKvkV1B32q/QALj1ll71/6vy2m6uuPWWYNJhz
DBBSY70Um+u11ZWfyUMQqtUOdrhpe0L2MDSV9OpN9CAQmXncylocvag3UggkRxeN
jOkB2NjoxtW/W4RQT+dcB+6vRpg4L3ChwIekhZVR8m6fJp3poVrO1VNDbCVbgDuR
taDy1LLlrAADh1RHfnIbJ/ofa7iipD88HUPpxJI7/WOAqnx4SnkAzW5+QB95opb2
eRlXJjAapI4iZ3EbC/MjNda4eKLA03/rfI7HAf8K2OB/L2liSLuaesEGyTXbB/d4
AqomWEml6P3ArFC5J6Q2oUzDzt/HlMeWhtGQYRq2d+chVghihc/CipHvscYg/RYx
zvJKFWMTc/5Y2NPVkZ1gAHl4t6VFMYZiWVq4Io4ioAEzhT0SP9+RKFMyWcxeKLMx
97hZ7QIN0FRaOWLTEWZ0S3nxLyZ4eEwVzqlkdSIH0AmxLI0lgigng4nJP8LNcH4I
ndvOZYv1n7OYZLirsbEDCSvqebGO5mgUWyWQIcsHq07cWOGVVfc+dF2dpJON+chR
wIGGUDHn7z3Uz/cNrmNw7PKu1Q/OpUvMaF2znO16TrgI54UznGf6ZRCQZSO6AUhe
+WmoiMDztrOYcnMsv8Yj7AiHtHRlPnfStZ7JKaherwT9lLyA70bqhPGHwGAjmast
CJQCYBxMrITgbSEzueLDRAUNi8Az5ix8ww1Y8cAAiZer1q7/Tpk9+d0iyS+q4JbH
zfs3FGQvh5C+oeb5ho7cY5okezP/zfkn+BGXHMiiFDaomP4mj1qrBCIvn0smmudE
gJeSKkBIpD2yhB07ERJVQTdMvrT6y+PHVFDweTUZPx0N0aZOqaz11D2lYbg8yQN2
l6toJtPydvVnIu3yYfAGK0n01ag1N4U8t8kLrWsY8KVWSVX+bPYCpRtO3lVEl1Ij
eWRidN4TQ2pCaX4fuT8940YgeVrLwfdgOxWyICh9Ebeos/QXyK4TcKp7ZcO2W+bM
Kq6eLbTmSZyHS1CK31GzO1HF6gg4W9JHcxRNyhHLxJ/v2yIDkrlVABNmv/RTROGy
eLXBQL4nhCRhEz59vP25oHbqL5a/udqi35lHt8+4eWLTewZPo8zUcMVSVGxWHt21
dRhxocOMW1hgHxRCpHhpAu6YKy7yMR0KSaW6ASMisSQzzxb9fjbmZw6JKcyNs3vi
mWxY0dCz2EzRqbItcQDw3RwuWc1MsxVOiKEZZtpah+rhtmVn/qXC/+pMSuLa2UuM
z6ZpreqyVn7t7zA/y2YkDRBc+S+LW5KRpT63ke+7cefsea/wC6rIvd5HV24AyefX
Kp/BX+9j3pJ6bk6jctnRES2bWLiPv4z7uS8t1Jk+WYYUnLB5aPGX/SXNe5fMHbad
g1MMS6Odq9933odo0vok1IGTOsi19GggCKrzLbl4ZXKybZRTNWCW9v69us4GkxE1
wVNPmCAOFROPra4fXFTa+jPzxYS9VYx38g5CsamWQEYWmB/nAqtrSSfhs9bWQF33
dNiQuAYUpSu6etpTMiVRnVuxpjRH5Awf8crm5tUt25tdIMELdZ+Xf+Kju/z+Y6Me
n+TuIvrej0iN793aWYBnEgLOtI/4ut2m1V3SpD6NfUXzA3HEMnGaJgGZLGkowvkR
yNnY+yaID6yXBDYZO4wfNb92shZhsfLvp1hokj1FtMKTeoMlfx7fSde0hXB8FTFW
PIchxgewjENbdcHyhRoXMHd5oRQD3iRJaaoAR43n++qrnqDN277vS7P/c+U6s/C3
0DbsXwDNclNC5Ih8bCRHA6IlamCeVkLQQ4Q83d/TFxHzJ9piSLM5tvNW9SqDkrb1
8/F01he11OoCPjoibS1ytTjGVkfBmMMSk0eeel1/Td1ii0clVfNPOjflIsXK4iau
MnbJplybYkPBE8ew3AV6zF1TTlxm/IjyDw8Y3rFQz/4mxuXI9qsiaMnP9qTqn9EJ
bAKmmpZPkgu856R+UtQdnojkbR/mhg2E6/tToBTAOVkuLmKBTE2HF0MphZJG0A2I
1dBFMQaUtuCRetD7Ku3UgRYphKyBbykpG11JWTDTlrV70XQWS8pVz6KgVJRfhK1r
VE5N71VBlIMsFG5TGrBbR2H9ZJQ6usfWvNFZl/1qTsg02niJm/Fwz1iIGd1expaI
Icw+bIWF79XgWmaGQgjWYVXUf1X1w2so1EZV2/uobEQNL0TMPKjCkoDucAqEOduJ
Thor1an5RoBSVDhO8v2ug7QjnA70+BjHnCqbTOblJMsqevWNafAXGNpnoSCSch7p
qZ55uZm+NZqw9zlkkTOCYZRWmzt66I+a+gHHaZ1cb3kuK6SeAVDqzi5w2E9DWumD
Ag1o5pOSq5W9nHEVCMbNPLianw2IMeJWrWzGxBd1ovCz0vXwlStwyUIpMCgrrRly
9YJKn8rQmTqFeFHOxyecgEMvlOnCGmf0UwXLg6hf0Egnjq8KdLMUN7LB3nKc6b/q
pH8h04HlbJyRPYJ8rn1+hOIukzLOwRQL7vJ2XR/EDr/MKJIWW346YkF0lV5/GGhr
pO9/5LxGnl0z0e/d1+lEwxWXHyGe5R0ak6S/6WEE6RDPyVzUc30HhVjPrv+lUGpi
m9eiLlAr5UKE0UzRAL4NKpyn2BspPubZTIc7HQNksN+LQmAo0vbgUbhkdA8Y8ba1
cTsJSyBYfFiFuN01+OEuOlAipffGaBvN3evW7PlMb2s07rErxmd/Jj9a9bXL1zfP
F6CtcIA6SK+HK2NN7gQBK5E8J0a/TZo+JBwnmNZD2ZHGbitXVQcQPuxibKTdZ8GF
s0sO9kSIYdAcaOpkr2dARLgrKang7LwFN2w1qpyM+dXwmH9ugPl9vsNMuS9hOG1b
SL2RqknfM6nq4C7BqjoXVKgICm+W0cXvgyckOuQ+PrmoLgJPeXHTiUi9qJZycAyB
h8mSuhEIZIYbh404GbpMHia+HEqySX/If9ZOpq7cmdS6glM1/CGTedTQtc+R1Y2d
brwXTAqCYN1vKAuJy04owvHgRmCqURv9fJChUjOrhVMS7yRHsdF+i5iyfTLkbsWk
UcT4NrSO4YoSp3QJKejtBPfrxuSCYZpQjhSX4ivThW/lb8u3ftNfwBVNdCYTNfaM
3P8Y/1/9ctitTGKWqd6ckyZKWkmIRG/Al0P09lJXpbcx2qrke488ZcJ0EYWrP0L9
S9t3kpKKng0dkjn1oAQOl4qNCXyChbVyIYjgZ93F9/OnM2n7uU7OX8kgal7SW9kn
MQRPRrC2iwo7ELuDMftBMgAp6kn1pXQJOmf4cg97E+wRggcRPgLKpYbJrkxcG+VW
AnXV6u4wpWgR/iSdH2LN0LUmDc2+XF0CtmONBLK3YfO4kObHve2Qd1VlunJAu3h4
2GgEcuTRNVGqHhucxTPj9PC0DmAcKym88ZXFdovjFKdtvZFA6oTc4vcu1TXKHA2A
FR7YTrVhvFGSZD0ksAtea3iN6CxKe3w8dyLe1sqii7PPEDfhTqGdLMfIxpn0LOc8
9AYpvK+m3eAf/mZYs7oJVpDTNl4wSX4UrRg9DFA6XWhQqKKnPTTC+TZ9eGbyoHSy
kQ7tA66zonZ07ID3iKkvcAvdm6Qru22vQJAYvM22rnZcKe2LBp6kmmAeM1IWTmCg
M/6+/QqWhD42vCO4KA6IZd/+GgrdxYeFYMfvMKfZiLlpYcnhWwTkdle7O+dT0FAK
5XHXPKbkwYihYdqVOaTE6QXouKpv7fPQQXzEJURPpibrc+uhYybI3J885ro83bcn
+KYylyAlaTpVAmfgmRzYb26D1owio4TgOvjLDEbdq852E1tBw+FAtQICdixKpfBH
2vRANejR8PBoIuqile/ip9Tj7CbxnZQzXY5vBwapm0vQpM3G1ygzV6PzrcyfzwI/
aXfFGTzH50yPnU0Wfc+wJGtEx5nNOkGiUQA3Vsu97C3u74Xs41lI7AefXNfDMcr6
7eR4VEexYuwUttBcjYRv7IFpsBwFkteiEEM3iVwH0z1Om4CzqlWc7vdul9myWUoO
T4Ot9i+WJW3Un5sp4UTnSqtuobPTP384MnSPHpzNk+EGiqoMsMvTJ5dBiabV+s0f
uUvxA/oriYfihFemZ+aJldYUNWT5D+ixbsfZ6DAuXVF6WG4w2e4KDZ+kWOW9LZ5j
mLf3eP1ZOVx5NEJrCaYmc5CBPTgUnXB7m0fk/xD4so3G+jYlgY56H9hIK3YO8CKW
96+BFUCM0AoZCRWjhX+/yh1Dy7N7HPxR6b80DAhTRQkb+8tKiBl+GBTPEMagHnAJ
rcK2gghMma1cktSppqtQqUSzPPNWisl2DUr1CmTaiI44Rx6xfoeE8DiaMxVNljix
FKPXBlEoN4TyHit+pgGZf/e5qN0jvi6rGmb2kyLDw0FN7R8KcUmhfIJRy717Eohr
ESbh9gazqjUCgXaUx3G+BeNa2kEdNRNdCwpDMKcbruQVS/wlukZ1b/S8pcCRaPTp
ekLjdsBjteISTePsykRGplPlVa8n4PfobIkrUINT8myVO87/OpTOx6KOSac6/9n+
r5NQQ7u5WecRufDI9frwyQjiwd/hYbiXCQKNAJwa0KX3CVNyw+wMCIkKeKMYl2fA
mdzaF0KSiKRmwwHWBDcKCffbFAQ2CBMD/04CdFiVxO33uZGWR6VmIeZN13be/alH
RuDAbbbZqCO+aJ7hNbgbQEx0zuLNOvFd9Lsk5Ix6zrVygHOWKOZBqQpct126uAsy
gn0v3dngrigf+gIYIRcj/g7vdc793qTo5EfQHfN68Lmv8a/OVHQ9/bSQz66F+4F2
XlC2uTnGlv3Ya7ehC2KXaUBvKmIckrkoiUCk3cOJ555ScXrnR7AQzPYDaPRIXEFq
6UILlylttS77eESmx3TVdL1n9kxAZesVVGB58TYxLghxpG5ugkmS/tqBdVCStdHz
qJ40UzH1JoRFQvnr21Wx+546vcu754vHlMJ2zpeciNhUNDkKJHTdZXzX2qZ9seEk
fI1x2dg5+87gSyqPZ5p2m5Dviiru8Wq/e/D+FvtQLoLQldMIGuKmTomj3D6zNRiH
QtbdAX3JgrDqTkz4yxfMpcQ5/Pv/324AiUb5iJ1a3lxskY3UMfln6EJrxDFWdF5Z
t+i18hXqVddyXuQKuDIHMyZ2p63WdHu0QmJpZA/DfObNkW00dt1XVX5eg3S6sFkO
xoGYYyZ3chdUcG3Kv1yUtNWK0XiHMsCCJqxnvLK63xCTgjrdhd9W52cRNXbnBE9G
37exV+Cy1DvWRQpknxbrrqde58C45kn/o32JAr9CEjKPSuSQk+OZdrrac3K/A/tQ
nZmy3nWAqouFddn3HcH9tSt69U/g0cBFmhfMbTf8IhyXrd0DoGsl5HVpRLgQ6kQ4
piiq8+NIXsv0ECwKALJHpyUe4HXKu4aHH8vkEvwFrmcBe2oNoyBasCIbCSTp/KST
Ye2BBOfaAXdVV4AWn/9fZGv8q2yTPS0Ew/74LKQvlfGRxFQB5wMa+6LV2WCutLIu
BRznGv1sBEmukr0fB+FBde6MnXXC7V5VKKQxYvrdC4TawUyrbMHVxZaOG1kDoBAm
ReQy7bHXA8pPDG+4y/s1roKzSMHW01iLZN1zwat9Z+PngZykJX8RdmA9PnpHAkN5
6+lZX4I+w3U+hL1fLJ8g7ATKEPVjU1Yk+ybdIgmjr7So65TKOALtzR/Fqlw8QwW7
LFvsLd0u7aU3q8FHSef++Y6GpU0T/kQ77+fWX0YWb58IU7htcZXFDFB1GLWuQfj7
DF9A9IMq7LUA52hdbRkUciLowIkjj4QHw5tT/wQ5n9ASjoEI1lTSWKjvV+z8ybNm
D2S5uSJ7uEM7yojanH33255K90EHstOyvhj/sqTsgv57cEaF1rHPvLyiQV58POxO
/UcRH5u6WwdiVcpArWhjAYEM7Wd8jCppFtfKOCTfk7WSQGPfDm9X8UGxy4m632Ne
dSTEuWWZF0+pIHn/YpYMONTTbRWvivymSU4ka723sjz2fpzYafRL0nr3/V+uD1MM
JyDOmfyFnns14iueYmCYz3yYIVMTZa0O7IUpMe4y71UkuBBWoelTOG3S7c3GRYmo
8MmyFAHUhUEKRfBrhYzMRwxb8Tn3Bg71h5S3hezmLHao1yjHQH+CoR7BZAMmXyqZ
YRR25aWaalOgqRQgxs9326Qn+DYAbRmJJJRBaY599a6LASlcndwuhlwccjzhEwQY
WvWsXol1yMuG4/SMOBBvxRJSSQ7+t/+mxn7sxtooZG0wJYWGg81GOud4c6JRcFHg
5u9o5Fsh77oCoZPxODKuZ41QWZMHK7D4Rfd8obT4xzeJvFz/SuaL8wIUBlRZschE
qzCjNlzfu/2osgrVNb9Y6LupmhI7TfXiRF3nCYJErNSoDsvlg1urU2dKHXwAHIk/
2+NRbnbckZ/IkOKPB7jzd67/0VxHzrPztEctFYbssN3RUvKjc5uQ0LcZkZAr09TX
FavIl6vTa8swY3aULZzqU5bsTQa7KnwUSlZkt4UJChhC6uT4l01XSJuli3FIWbfO
5efpBZzOQQ57esZ1TrEVZShktihaFnYanqw4yEK2Jm0/n09e0Ibjou4abLgepzsv
0OfZW9Tg4igTOaiNPbYbsISHNhTbdPUhOnSKJkJwxxPLB8nuO+4Nd0+rx2k9F6V2
4hCAxMCHp9Kw1286iDpLHWaBngq9DyKZLpeH4acxj/H+AD8FsCqEXpgx3Yf+sz3E
YoTcMrPpmP7XEyRvEMhZBO7IACszSSxD0zTEXWugKHIAGl98CizcxPR6wF+O5VSK
9n1a/jtpff9Vctby9G/ei6GR5bvmswHFG3mD1nSH0kfyNmgPy1lxpZbpQFq1KOIu
OYh2oSQsG78NBKl7MlOt/l8VfxWS3pnjTAabpX9OiRlL/YJUihjVn2SmnMPQNne6
eNvuhk0ZCg1rtczMlkm0srWpbAdRI2YvuhFYn9WTPgXoyOZB0STKvqbRoI4PS1tU
ox+7hzvoB3Uld2RsA4VtKAjBGK6msoa/xjocWhKNi0VuM/Vfe6Ticetyhs1ihpYw
VMNEYiRJM22ngVfMelS89vpty9nI9czhVIb5JEwpsIRGLCpVD/y1MxwsvA4OyYVg
mal91aut1jP7g5En1AhQI//8Xp4GAJhRNp4Yoqt/TRSxWjo/iZaRdifE6ALWeDq8
ZLUdKA13sGGRZRswVnHFUKqkS+DCLbA2GiMXiH58zcbGWNw2tzrjsnHeogc+ErB9
K3UdhlfmRhs/Cr6mH+cWcpW49YKMj9BqWSLl4uWl2nKRMNBFUNWXAEz6KlIkUEfB
RkaeHpcCwtMjxahFJkO95fKNjb7/NgwhiunSpGvOusnS7G6xyeGoeOcBIOQPrdEa
wCPPI5dLcfGJYNrNN1iBBYYmeWQPDokrT+3LsgKQgcWZMXfuibz1tq9TY0Ql0EFx
ly+GRe4hTTz/wSuRKN4RLHxN2Mm+HbAYFCKWiiULO6rQPcVPxJPXtwSKD4HEKOWe
QDo+APQS8RfhHpTRghQvq/Gdko0M3Vdrebr9Skl+q6Zlcv7gUkHkwC7mBC0A8WRe
1DV3Vt6FKL3uYkGbq98r2jmBG8xz0F1sZyG6F3XS8I+FUsx30N5NwwfdZnXtvSov
Vc++90iyBa/McQEcFqdXLUsJYnkUVfTtp8k14NmoIJpO8RANf3iojXaDIDqHVUZD
gZW20K+6mb3mMN/EvgvgKEoA6LYxQNurv4+LoVQ3CiEwQ4CJdnjoq5p0aYwP5I1Q
VlmK5yABpb/9s2Wzh9Cpd+HxfGDnnW6qlIfzI4vnAx18KDWpHgmOkl5u8/DRLRQQ
syyG8VZFIATsVDHaYR5tRI5NNz5ywNNeyo/VGMONjAye3Jxy/ZPKvIeahgm15jSI
Uvv8QQR4/kf3WkrI9XUMQuf47d4EkJEnNKSB0aT2okgDNG9qsw8vUhCgPf2t5t45
TNqWHZci5/QXGbWYHFHt8N6XA+XbHKxGUZqlGL6C+cugODg3hBlgqiXEF6rBdmIF
QSI481Nj5C6a0BFi27EF4k99hnygwAyNRGuJ7wSzGMPrJ4ai1kGePrjIJ7ZxixMC
DyzRllaN3SVJUZF5eeFDjjTV8pQXNXg/80Ol0a1yTBd8E8WBNc2b/TZWzTy9l6LR
md6cgg6j8CzP2VT96778GigemQonzWpeL5TeWSO3isd11r1nVlbSGqWUxHX0UiZg
QGAETUbpocuYaCVhYur8egIT2cBxGDk9X3G15BnbGpGv8qjxIOCA1ES/3BvNRI3G
GLxIE8W70fEcwpIynfCeU5fHLoTBsPnqO++7JyeJ8jkMTN7adTr3VlBYUghjDE6n
y/Lvd1+FpOhUojY3rEUvL4TROgbZpGhVk7JQc3FzXLSKvuccHdRkEBFi2tMj8xt4
jOm9gdq7J/hdbZnok4FROgTyMCawPVloVKbIbpZ3A0nVDrp5MWJEF4vMP6PDkv/x
Pqa7rgjoEhdm1ZY++vvpeI1Edr0yKxp4V68MZPo5pE9nk408Vk9WBHDugDLX5jxT
bAzooo7gi88TUDTXFyJwwEEr1z2ahScza2rEvUDH1bnN5fEmy2HN/ZfKyEPfTdOu
ptpfvor4qLdRIvqKXOaw9oCMMxprUYJ7UIV0OnbiNW3Rs1/XoAePJeVi2ebR64T6
LGHYOnLaKBt6b/EtfstlFLfojhBvbU2yEm7nzNVRvkG9AmNE7ogbzFbjj/zEuKN2
EeUrGcWCnW1bdcP0GZnilq88vKG13emkvfPtuQLEEygaTYwS/zdtryZWgD5hr4Eo
u1j7ocbL0aXxRSoKj1hPtkPzY0nf4XWvOp1XgZgiszdwSOEcYNY0S1zBA09+WlCG
d1NRcdryWtHW1gz7sh9rmP+J2loObljOkfuBUQcK6u4vojRR9yUSput9plyY4ZK7
UjcDAKfZJIgBdMPHxSA7v3cPciUwIuTfyYRDL3VsBji8eXL+BboacVT3rUamB7BC
jpyYyw6j5BJJ3zPlIbV8pbUmqDWJGeIIvcaJH1oa6Sjwiu3BIjncty1Z+DdOWWXO
I4pdjSOPvEXX0qMEeX2RV3U/rUYmGQMCL9XgiGCOGnks2Pfe+71LQinOelrxvlDS
g/wkM081j2875vJkjfvV2Dg3TEV7V4jumBt5v8bg6yvVAtUuAT+AOMyJr6YT6r5U
WDhzSF/KnLHgqgowhDGRT5X7HzKYA0f389cqd1xEF/XdyLl3xK6YrOJafgZdf//K
fGnk/lznbccdPSUdYjolj0VSosjbAunfk6JQlf5QQrkZRfiDn0w93pYDo2ANxhRQ
gZiDaRE3YcPtjWt8qrZA8KEvTRO9BSX5Mi+aaK4/sXdguag+82pEtfQnACpn+g5e
6ZOTEULe0XtP/TmWxSQpyplRMyT6TI/P9TEVAOwrmji1+/bQnd73+6ttXvuT73KA
/snYtwdo3ak4f3/DtAoZltgHnsBVvRxZMpOPNdO7sKUbUP0weP/hrHqe8eWuPkqL
NN8wgJ1yz5N4L3jhJp/XpLZ45BWcYrSEbWHR22nst2DM5mo47ijH2nZ0jc/Z190W
HFlh8aat48wMsDVmR7BLvObU+hhAQgL6FobfcUZHQDjIY4oZ4g+baH++V9nYc94t
Zsx9jAQQERFOuX80gYLGV9jbqCsHhcAXfHHHrwjO7kmrjkWN5IeL0QNYb+zWTGKX
JUwwnKoo5EQ+X6xRmnVd/4q6ZFB92w5H46DB+LplNtcVVjQmU/qgGKdb4ueBxGIM
zGlt2+xuujPKzI+Z3N01dFCNl9MT9x+5EvO40Pwbqj4wVqClbpYOWH99OPJaUN4D
M6CEvTMgRgIuxBiZFWygcMoEVth6kMMX0J+VwIiCMxYWT24o0/TWpOqFLa5xgLCx
qLQNcCIQOUqt+5HaWj4bKxWVdv0r5iygKUfggKRQ7lyxw9ts+83xYnAXVY8whfhe
XTcphIPg9KyCBkyZCq9T5VW2HwKRzvP9B2g/jcVGOWBGDms7cp6DokCvVWAWZIk1
Zi6JVPnYCqB152mZFYQtqt/SmDXRo82BSsmUDu0iRhncay1ZvwhHVNXrLlMMnemk
fTm/4TE5wh1pTRH3YbfLgZS1EESd0qXVBXbBBmFHDMrnIFrzFwina3zpQHqaNvQl
MqRJqC+46QqXhoXXMtKfqzCdNJ7eKaltpQRQ4UL7NeFZfdwjyeJ/4oNg2IOg4d64
YOYbbL16AvxxS90btM35pbHuo6Oyyy6nKDb0QV3Og3ZG6Rsq/+/3Xt5PS6PzqF8L
CYw5xD1QMglfqCVU35tAygm4SAQ0kgGA6uL1P5S2D/TkvHoSi+WDjqb83Ympd7Q4
YQGPelLR79kff+7OxEpU0BAuvDS3mAcaick89hY9g5jcPNErxKbEj9z1+M3PHOPO
b8elBkhZWbtcRDT+euQiMSwUQL0f84m5rGiUEXvQY/RaYtGa4Ru1EQm2Rq9bEUnc
U6BcggWljUzKpB7V1GJfIxyucUtDPTtyg53Tz3dQ1lyQ4cUaY+Lg8xs3G6wD/NXt
RqMSpvcjldePoq0Wco3upnWz+/ajyfdDAn+QfsEl8DhCpAA+y7kA4tXKNxkL2GrQ
tQGi/AoUp2EfXsobmLNKq5FsQIzvZq+uvA/PB2+xG+/M607IPjpfp+NMwBRYl/Fa
IB57yyHxpz0bglIEpAxr90MZO2sjKCmRkKnUG9lOp82j7dEPFyq4u2yfYQ1shQA5
tb5YUgRUPDvNKBvePUpB0ynWylRsj+Nh5rHqJD9nYETzBK+BFm0BR8HzeVfdfJqW
cfO+erU4/twy6LAntzIU5lpX9ooJIAvQ9+5QJed8soJ1xSCbX1K1RtgUs8pan6QL
ztzUuz9DwJM81/IFMzdUjh5NFe+rcLXcQNLoj2QNl5E7sKx+c8jsD1O5X8ddO5He
VNF+DQ+BxpNvVNLl21yYw6Qz74R7nRCkVq/AhATyUEie7GuG5tq039FpK1selDol
d8SmzlsFeIxiLWRxkvHvaFHMA0X4tnJdpoowpxQe6TYDbJVLJLZOs1FYWI61a2WN
PuhkaAuGh1tdZ3Z0HTMeWf9l8wGvAstWa97YmZkcQa+iiEPHmaH4OLdypBBsIbZ6
z+BjpZsUQiNnWp23hChgDoGOvRdaFrNaM6fZpCxD9NyCiuMKkDr3doBrgL06RF7d
incVSU2Zz01bXGLnXp5nxjJdFyBtQjkdAP38w51lWZtRTOZXmi82xtipB+ULX5YI
mGkhfdamNwijwDi+iaslVN33zi2KrG/6uLPTlEhbQ55OIpCxdAfCnDDLlcZT9Qwx
fV7aoWIaFN7TDJV2HVYofEMYxIprGKq6IDceyNu0yEKaFAGogSWTqzxkuYdS0Box
DBDlh7LQ6n7eeu24PWtlJ7dQnuU6XMVCEvsqVBJrPCaVfJnqZ6/C6FMqoY9XBh6Y
RzjPL15b1i5fEVlHMEW2VAC/47791psLHV9NrRv8PC/j5o4txqHAJoNYuINIv9oK
M4EUP7FCtl00b8Qwdf8jYBWR9xry0LdndTQW5pWRr3MXBiABHSjKVweKRzAtsooy
O4l5uKNNkbu5PBk/ogBS8JFkwUhS48tAiRtl+7lNxl320IKcIw6Qqxo3wkvdFEbz
YuZJ31P1ui+XLwUaXzddRXv4RHNiUq2mE18pVfqijPe/etOX/PUeYzv/71pQhnTM
w2Jy5bVjmnumoCmIpag62H1cdLjL2Nl5ikJGYuz4Xqn9Fl53SN2e4OzHB8PXvhkp
4J9ZGkA5jXYwuLkJOCP4aF8lxacutPgVwjYwB+Byr0HXC+UfM7cBTwNZz7XNQjx1
Qu9HUGD8B5QkK1CpNohSfgOMTmPvU/CNMjNMY6oVhcb66TYW+LYWci9KjVprjg+V
jxjubGO1PO95CLO4UXR5i+eNEBaXqas4QV/aIknfoQG5H5TMUSkWbCMBqB333qlw
LmB8iIrsw/J1ZgYiDAUa9/LB/IlnbqHO6dSBULt8WCdX0B+Cso3AtYGnYUSFD8cE
ullCf+pDOEMdmE1QbiAkHW5mH+s9YXl9+2BoL82sve77Di+N3Z+59Q/DlkXT/HtI
25yFAn51TOJlGN6kxLHzU8QKyxVZ5ByAi8tHKRojzR7+naAxIheUSbnSsoSX5Kvk
MJzE9V1m7oGjnskyNqqQ+uAcvilmwUcU2twD5DvDmLIbEacvDlQbkWQkvRCT2SzF
g5d/ZP1c4x657CPG05oJrtDmYIG28o54mbQlT6infoXOTaOct2LBxIRudyswQXz7
ycnwE9DgJzKHJ+iyDZ4SLKme5Gz34fiMQN4GbiQg6lbJB/ZSNI9xxwpa8km5R9rs
IZ3TpBxi85StGxLIRYCug4KpLW0UW3ifT/nok6lCkhLWld3gdOS1t1M+wWnBwJxi
1WEdjn9GwhlllbGubZsFn1bmKl7bxByFDOhdu8qQLhe8ot1yp6m5MDl9aNLdLUHA
E2B1x+2+yuUo7yQ7dpYZVMD1DIwp2YP+AQl4jjdQTKM303PLbS+D06qRjGVl172h
sDCiP5a02FcynijsPnToYjMRtpS6vda1WXRiq6vugqWH/zzpv3qRalQyxeDYi8vY
8NnnqywKg+I2aHpNJn8VJOdFg2O+MeLm+Ad34yHUiCJ35ssBBwMwdNR4H8/Ws4kA
8GUsU2e075yPHfk04PtvpjYgc9kdLj/cGq6Pe5IUKcdRaS+uJKkh7HYoF78CyXr9
KFU3kiEnHJoLJQQgXzTuCMl2LdIeGsKDslQ9FSrdE2EmhDZzdnz8zGbkW2BcblYd
Ql2otcB+C4/ANeCGZcW+i6mVs76IT7gwUCTJw7iQr1K7iYVLOb1INuxAeNiGAsd/
efmSnEh27RgBePAgwGEbcKYBC06PsAd0/dYt4qbM5On3uL7DPnFriaFRX1cMY8C2
TW1OA1oOioxlL4lYtj4WYQICBfRjWrEGYHQ6AyZ/4U2r1kWFVs388MCJ2xlwENcU
XY3N/IvCRg6ynaUQbxGV7mI5IHV50G3xu0+cbRqC02bk0v4/R9+7MGoX+iEUEGXv
RAe73r7wWxpxCDMmiuP/acS/PVVkFIKGXvcBJ4lTHyY+BvJdBXCzl26W3Q5lq5Gf
Nabi6lTbi2/uZ9HWLxJSMJGlax4S0/c74ppBhxymyX3ytbuc8ZOYVmKiipQ95s6Z
AByJnekG+MzxsFwcoQzlTVsErJp/p4HCkjuYGfjSFi7FI2kL+CVfiGuM8ql/Mp5K
uMcdO7yaphfQEuaA4ao+71TSwz1/zHBaRRX74M1VmROiNOCLbtAnF1PsbOet3rJ/
SFSfCSQOO/Y21PEycsgFZ09kJqz85onDc0TePS7k1u/vjz8LYpDDLuCcbcRAnMFy
x9oMMgRe8hdpkgg+u2E03b5qqOOmu2XA9rXdeGc55caO3mCbpYEztDEktyfL5ANp
OwSdCPAzsSXvteotFQcFceFTEvHyEPz3nFUr1uV7D7Nsw6N0sx8cHR3mi0tgjf51
IvsuevAxvBmSnWeh+hfu0H/e9rfmEDMbsL2apw05MjjWBsXOdB+V0w1AazNCeY0+
9cqxFz2blcpv4sNYLOaRSx7EA0AI0YwK0W44USKKfitTxckamhRsl5N4eOCrkkvK
jMDPEWQl29ovFFrWd7LY8lqBsytbfBnsFqKmuCEGqdqX3vsG1cvOMyY3gKG2kMNY
I8xB73MqOG70+GQa+I0vxsOaV32csmVRHKwECTVzv3UUgNBmzHwP+QJXsHb838UN
W2mwxm6wuTq/3+sEriTpakSgFuIf4joxwUp206lO+YWD+mvGMGsZoZ/DZGDc0raF
Hq+M83ORlBcUXQhvonpDOT6jqZ6iy4ToL/8wH/PrAFdHrHFAL7b+aPj+L9YDtFFe
CPHBD9Xmog+BESXC8tO8mkOGg8Y0HXsPbThicYHTcawaRQEjIGaofJfNVTVULSw9
GKBoHmJRAPL6LlaVv6fXv7uAnj4xXxPJGVBV0VUEOXCeRZlVHtp6rEw2dkyEQQLM
8/2/t4Qifaj8Wsy3Sz9KMy0SbPTPVNsvjAO1zv138lhiJTQIQk6PqSB3E8eOAb+d
OKo1yNkFahoy+VWb0trBaEpKiAc8CRv6gnS3M1d9Crofs5V5G/gm/szjf0AFmDhP
S5GVA3umx4y6AinZsk8MYEVXiJqCPb0FkUqrYRgb1TKud8aw10fPaJIaBMkY8Kmd
Z+CE7zuaaAItEKtPxJ5hi1d7isfbzzJ6hROtAJUgY17bDGr+vmroZWsMUmHXPbBJ
5+gdn6cyC+IZkWw4VSSDDyy6vQrV/p/G9X9Qk+Sn/f7DkMWNtB6V26glJkT3yuXv
1QHHqY/b9DB87TJYNun+bptBzkwqQqdgW1nTMy8D3hfp5Vhx3c+79EBi9eWJFSjh
hsQOKxb+c5z7mmHSSUBxnZ21Jsb5udikdUYwJPeRsk4E8YsVDf1+5L87j8HCkbYf
nSC+U6GGvKhEWE0LF9Fe8Rq3Rq7o7pXQhfq8ldOTJXjNX8fIkSZ15+pQMnqUN9G9
eKIWFD9y0H1ZRbtbb17hc1CU5K9ZXt2a2EHRcIiKCdHp7nvUz7LBH2CsDfK7/W7k
IZtasX40pmqVHXy3qCnqBKAzb9dh0ClVtckpu42fLz166SMUbesA3X2KFbIQ/1gJ
FZ3eWe5wp+9i2l1eaMzFDIj1eLpbj/qL++RdlgBRPpHTd5iC64elz7Y51C6c/Z+l
+Q03NAhQob1PozfL7EKJTfBnHbPaKExjt+/MWAyqmHUMov6dGMAW0kFu5GFCzwNu
xeBXlcj4qrj6kiWGzlxknuSxoeqhtQ0Es04OGS26eS6qjkTiuZybjZOzEFh7ul9n
8W3J9PR6v3xz/wsrcPRhSm8UaHupQsHdjhoSRTrnVoVwWaBFg7WBA5QtSB2MBvob
zD0iSFOxx13zn6MOsYSiNMY8l2fANFzqNNFwf2dMzbljM6m6eUeEUJDS1A59eglK
Dr/s5r4CXnZXK0lPVcy4co2MVa/Sj2hBJqFTc9US4XNU0kk8/N/Q9bYFDLI7uc0l
ZTxYa62sgufDeycErgV/Z9UIt021yBYODp0U9E+0k8idnsLWz8tsNKu4PZuM4OS8
mIGoOThfm7mCkB0pK9MOPOr1WzoCRceqKPzJZPmzObHisFsooNCoYjxjiL35N6LH
b9LZqXN54ZgbKzLCXMCVhYPlGqqz2F7e94ThfueFBqbkilyy/h6Rjfv2WBc1JJpS
qufRNAz5nnUmHU0XW1BWiQtX76Ca2QSodVG4/pX4hPpnhCvgigtxAXapjLLgVbv4
HaRmYvElZHJCXfduEj//Mrwjl+JjUO8zxjuhr2d1IeHgL1H4mTbzhTUTONzwkrKs
pO1G2D7qgbHEKHdw6VZjBk4jnMe1Z5sRwriKCeNjnI3KgX7BrbTSf/Ks28S9qbyi
y64kUQJ0IdZ9/lV4c6v6p/9yGcOyqZGzuFB1tMgGrW37+iDTmufA9EEBuZwShl1s
tqKVEAWBtUG/HAZTFgI2pRHi5jtKY3RkWhk/ut9RTi9MhL8KPOkCTSLw1y/b7gkT
5Tuqf2pcOydTganOnThX0OeUJzPb6x419k2YI10rcoqAsvF7/88KzWZZJsaa12pL
wFozObt7RQvu+SG6NC9Z8FYACIBwKpQWzG6nuNR/01jzv8o8ehSK69RUxgJ+/1dx
a7IS4040wpxznvf+n9Syh52lVhE1u4afQwNI1t+v5P4B9ilImoL+aGBG7m+x2KM2
nia2L+06Tqq/P4qZn/8D+n5WaEVcZ6M8fjYSiojF/ePp3jQj1kUilJTQ1DrcPEOy
Bkvs4nK5rqjauVoLEPShMf03qCVn3oDApxB1VOiHdUhHK177Bg8ylaUbxaohciBb
0D7R38jQTpe91utePipkh9bAan5x5182VP4ewDbfN+4Uf3LuB/Cgc65HGTY72yTh
TRn1blIVL5TaV4BbaDTtSe7JCLP/MObbwLQmXD3Cv7HBweddjUm3lJI2ybjyMCEN
qrNsOjtrt21JswP3wcExaMpYY5siqvWQgfarSPhpyHelL5nBoNfnSReIi7ekyxB0
ESgE/yrxtMjn6GAMn4D7doidsXXpLgWz8hY670TjmTFG2jsPoxV0zRFt3hyFCPO4
f7txHt9S3D8P/36JhPQcKcSIiFVSZUo3F2nw+FTrd/W3mIWyZPY5v/a7UeAbVpMX
OJNNDjTZLtgYYoCb0Vv+lz35moDnho+5Kea39+JT3CVstYk67JOz2yKrMBrRHD16
QBz4OvloBRVMi/uzrDy/hdY1Q/6VqHxqugbdAeCNHCvp7Fpo9mo+WowIha/g0rRG
p1yqU3GAszuRUwgp2Twe+2HDOPRBy8yzcywTcgHv3UYzeXhXeKuSEuV2sO96xIjM
IAeL9xruZxpU0/BNrHAvTTLCSTsiXx9u0NTVmswMXY10qkrZevzhZaEaNdvlsDPi
zL6Qsc/MeU/lVBTtgXv0z1MW6r9yAlpwKhqpv6baK/zgvLY5BG0EuSXD+tTaSnSR
9ZsKAOGRJ5VIaC5zLzX+fuUPwUaNkP8eY3QYTjof1CLdL7eQP1dIcNbbr94ER0J5
7kFY3brEO/f+T6AeeFNCUzvHlgFiNu2gueMNoY/0HoCB0mndVCp8oKKJJIrzJJaz
0E+cQyGpxp+5QULNiVgCgS9+hNK1bTWjhIg5AHEmCEYzpivkWVuKnJ6FVUNG2VI7
DVbZIce+0J/ilmvFRBuW+pKFwSkGCjRaAAcjY/M5ZjUUaSAoApITLi4xHTmxoW5p
cxuZnnT428+vm+1/EoHxvLO7RQwObMnAr6EkGknqkE46zj0tpxvxq8ERi/54whhQ
EeWdUTt2xhp8pe4ME7Hl44J7/Aa+74Sf3AmYKDwZRX2BXF6uS9qVOoLcbRv3F0bO
hBBOisS9CNzUkPdVf7bPwTxv9BwSXEhNmUKjtZ/pwFvKCgAnTlY2gKYS7ApRH3wS
jijSCwWf7PrirWlVH2Yd9iLgw09rUDZzGiCcV7tV0y2sXrCJREHU9SA/M78k4eNz
7loR/eKg0hyHV+oGbLGVn7m2kfW6uCfJKHfxAg9mYELLyhXo7NyivWh5P7I2pAUT
PkqGZrd5nlA+EOT0yYUaEPoWZ6x0pJDr8yKlJuqE36u8DzyoWlUw39AWypYzZ2dx
RrRMHjkbt/RfVf3cq4iSJYNasfKMa9xMuiIdP8pDraT9EukYv6Qu6o3YayX1/C4q
8NnNSwrA5Q4Oc21EYyrwlv7JGlXow4E23h+2HkkaxsHH7suOCXrTY521IPI4+/M8
0xn6xAW/UxzW6d1As5hj7c8J1HVaOHOhovHyabK1TIdoa7aDl4MUYyVVMbrh/edw
mQypPySzLtkKJVmlUHHtTdz0djZp5PYUyHw/UaFZEQWBoexTQfih/HzW+OvrltfE
fN0L1Innl1ir2ScxleYAIQmH4AKbASGkvTOMT40GrmC6FW9qIo8ky5nlwQF/Z88I
iPZb/OM98caZtXlDlK0PObzZvCC9hEEUoD0XX6jgrtzDkSEog/8xN3xHU9kDFrEz
jrgcjPpa/7+AmEM05MX50Lb/qcsMN3rcA9FQEAuP9TnyGC6lo/cFpIc0KBvE4QVt
NbY57XRbC4ZRoSgMQervCA3o7SVj+vWdrl+rstwBOaEw2fL+KkMt8EMpyru3k6MG
0BaWKjGzdccQWSvzoIbMI1R3x/bmtwkz7gcVYqbH+U0BSLbL91+jBtrZGnz+mUfo
6+cOqlBVBGqmqpfT4mtjZM5Ei4PsZdrgqpxmlYSZIWNtDMTGYNc/lWR8J/pLz6/t
IKNqjnnl9w7A1nsUiuvprmE8NMVGaZTkRfJS1gAq4h5t0RBvckACVZxYWM09SBJy
FErKBo6ZaNkOTb2wpNDbO1jokiwUQCpDastlnMO4zrbP7S1AGoNof/4qBuOKUEg4
EKgLhTQAMZPZ76bdOpUGNfzGhbKMjqu0f7StJ33VBrZons+8qKvg50SEjV17EYRa
EeHBcyF11YleHp9gk/OzBbTfFoL0C0nMnsFHzZB3AwNOBJOFsW82ZPY2738AA1DW
htIPRtoshTh3MwKKybXyzDpQKGm2xY2eegdC7wkRolmsymYq9Cep4IddR1VvmN9u
IICy/KwEW139f82UBE4QWMPVqifgZbye7sNVejC41f9qLM+O/JBtgtHtfWnV3pl4
OiPrS9Ait35aznjbbkmGUx3eUBl0nIoyd6riZzXUC1T7cR5QuyoUST0ePC6c9nuk
KFfKMcc65VUiRahO9hhQ2UG+yn1LHR7CSAI7Qnsnx+3jXLjInsCHu2KsAIzQ+1Ot
sbyD0Zuxx6omDbzcm1GVRwWbzE+H0973wewiOCCsq0+90SImXFoEZVXVAxeOqYXY
OI2DJC7YtHZpBT1e4J0MIwHmakjEab8SSEPsaqzEk1NXWcxCbVQe43eGGBJ5e4xi
A7BRzVHziKdFWnsRZV47zixTsfHe80qx+b0wZLzfzVmYlNYN9hFKyi/sBe4+1Toy
coZuBlZIfGQyiI/qKTcVHOoO2UQGe85ogDlELtk3Gosq1vtLOv5pXi6phLmudP4V
YoP6IdUxKZO6tlm02USrQKbODPB0OC7t5cW54eR4yQBJn3WIrrJ+tfuwdVu8IM5Y
vcc/WPz9E7DNDNmDoUsAn6q+7ZQYitnptoDjgpAr3V8ZkF9gCsH4QwH9u1pKvdIx
0npWMebMdZDQfwIVhUeZ1vj4pXBhdMb4K2OEBNahgRwUDk3LIM+LK9S1XtUqG8LR
0tbhjGozgSP5k7gVFMzPyVNh/GLslLTGUbDxz/eXXE6xV5j6kmx8gAM98UG3XYEy
QxBk4zW3YD85HDh5YbCRoG99y8FJzlTsDd+jQHdC2Y80WJgHd3hJVXvSTYBJQ7XO
Bm9nEz9xwgVjy6bcVZ80GCoPqipfoR7KUemoLlo9eW6cQ6F+JeJUZ/TDi8kf7CCa
HvgDWJITwxwN9MFL13Lj0hdk/ctc1m8FAsx3tUyqqOxEE4iAPwsV5Oi9FBjxscGe
KH9imX6B0Aq1JycRsUTKhn0dFO99QlC7comY+qyRjxayZj2bRMCrm/zhDUbCSpmO
aJ31DUZHnXTlVA/45a1VFWGUgBnis+dDSA/q0axLNmLxRu/SD4YelDXLjvW/fS6J
XXzMVq6cHVkcwNQ8JB8lhO4xrd+9VLbf6kfaACPYjiwB8U/mM+HCgarQYCH2/YYN
7VOaCBQMirDkeFrMZw8b6PvACB0xBKWZg6d8H/2rhlwg5UJI2wlQ5OIaCxUECmpD
ohSgDMHyuctfDMkYnanleH9fuTeqz9a+zmVUwnQTY2rWqYz+5xMCLdyC+CYhGM9f
HJjROjRo2dgrjsZX1pGeBb+wO8Au+jrm5wb0T1xtVQpdMM+nbeVdg6lWqyJ0Qu0t
uD7ec0vxBk6hyZqB9DnKiYjLQOvNweFxZmxCBLDKz3RXyp88iotW96ebCWl2Hen7
hsRdmkkT9hIUt6iZkNn3UuXvIxJ3riIUOBK/kESfc3EH9EwLn5L1X/9sUaLBgnKc
Pup6SlAhr27XxYrmsoAnD6tHMIBrB6WHKCtC0YiU37xCyWvcCpyXrGZvgum/QbGH
/XV6LVZFKuQVJzk/5tw9ls5d0XLkwcnQWe9sffL21O4QKBe85Des25FsGmlbke85
LyTC3AnsFczl1NoaPmeuvQn/0lt+JtyF1mEBfL+L5QJeDP6l/Do3g2YD2AY6dTkS
8/vWSITjmHQjqPpLLPPJkoJLAURe1PpNvdEwKRY+0eQfQja614NdezlbsdhQOq3X
036MDYnysnyaSc6Wk1oJSdDw2m20j56kj1CvhwDqlPlSZPepMIsRa0vH0diqVqS/
70BemzWco5FWbjyDU6Z/2OGzaAwaai6B7RBZot4D+hr5S2uw40Irz2Cwuj7jrUDs
Xnfc0HIlg9n3nnHbdu70J9e2ExOQQbwbenXxE7zjo/TUAXHF0roDcoyYG2hjubbj
w3+GGv2A+1QlMyvH6PRG1QaYHMF/7TlSaNiFOhYniBKvMsRbmGPS9dPT9BRSzWY9
FOUVqsZFFtL2vd5aOasyi0KP0saEja765mRL8d4ca/5HcGGp74TTYgWiQf7mdu3Q
AWkRrrSZNlyK3hizgqTVnuub+l8KiVtSovRIWvjIVI4TJ5WNuL2lXTWhFU8zgLAi
FvtF60zoq6kanVXKnl12E0TGpQqIpxv0UOpbH/q8WWiViD6H0M8Y8G4i0ZurJ/Sl
Wk0lj6w4c/KuDqYAds4kZvIOT1xOFCl4qQsKBivmLHQ9nZGg6xkhMSZSTeRad30R
sVoSeSRwgQbS/up9XCjJsChMOg/Qxo25Df/B0FTNBiXzxxEwgefoDNWvwDo+N426
MFRmXZFI7lh4koXI15DDfb2379UVMsVrIgBxofD+mghL0EsTHyezSE8tX8xc4iYu
TTxKqCl30UNnJxHFmCs/zgG3e8cAoyZwMud8pVHmHdasTEgB8pI8nmSh4iYYnrqE
hoOdz1b5B1xQGZY8mFn74/j/Uyf9GSS6CyDLeTZMR23vY0XnhzwVfpQv2caUHpb4
ptQPqT1RZwDicCstJiP46sd1XPMl1lgMokQcBtwZim8rYQjXY0sayK/vW4VXDEjR
+sq5e8JccBlY4YQPeQbH58V2heQGcd/laSPLdUqpEepHtx9NLyNOI1vL0MexC1zG
BlL6G1Qvs3EpEV7Xazxe/A++aiQazirEr9tCZIqIehxbL5AVJPiJ83Mn3/5+g+DF
ZHFBSJITgPO8LOOPNtZ1mx8xM0Rcu0Nem4tSPZ5sdXMW+9Rfvr1CMo+JuG3FtX6C
SbUiKDZPutiWAyMunwdzYe+L7bwcAzzrlQc9Pr1WrpBoH4Fv/67ZSPLkiGfZDa2Z
G6ODXFbmMgTOPI9wlEOS4lv2ZRfzpRict7+ijygwsARDxQovNKLfsegKUAAIzrOw
HKA5mz6y+hgW85khCYDKnQ09LyyphagOHZnbmQr6LztTvaSON+HPGuhssOgjzy+1
VnqbmE9wLPsPANtdnNyZH6zRjIF9Mv6Mx5iABXmn/AW1aiMmFCsafLxv6CSsGNZ7
bgGSRK15qqNfPU+z/99jjD1MJqFyLnHkRH1kismCx2BIK7q18ULpvWcfymuRKLO0
WfoK6eJHvFgwPhck4mVzWhZ7lH6ryJWyP56on8msEiAH0a+M0vrAkCkzoz7L/906
D6UBU6YU9/6+nd5jjJm+xvkksPMEt6GjJ3Cz0UvuQzkMygt1t8umMsCX/x8UaWuR
Q7H6Ywp8poI5Alxz5vT7ZdsS3mgXSNGQs8b9rm9WNCKaKJn7y4mBGa8nFlGzqvdE
V6dT5qr53IAyx7egXG3uSTEm2MdctH8Bk1gsGC/3s6BHgUtTQMdnY93/guWit19o
GTaEbChWdtibe2Pxu+14lIUlrImXmDN3ES+28+CY3ql9XIzmOPperwvHVSeGM510
0st8a6w8sYXngHolXbbgr7OHhtyyLT0X9si0uig/XtObXnDcveCcKWybbEFqu9K2
fuibXlfEVA5vYQCOoaJeTvBDqAB2uoevKdq/Mbn1b1PC06OHfwJ9wkvQmf35rNOj
C86LoqdTtwMDuCoIt/qdDpqn24wD86UMRWK9WpzeFwsROA8LoY8tl/Ic5Oc0OXTl
oFAZw7P1Jh94UMldii4CMgHX6FViB0vVFqzHXcmCkPl8ifuYlbFs8FLQb2RAVej4
BKY0YJEbW7ZCCWFwAXGyEOmaV/gPynONO1LQmwdurqTsh5bwaiTdsrWtLL2Fa8eE
HnjA5eY7tHerrT0B6ZYyFAMdysoU61+TNn7BUefDnq3MDs08sV8kHR2CWqSMj+iO
w8KNt/fE6US9L7ro5TSclzGbb+phb45AtrKU6Bvs4WjZCcCIoWUgj7MpK1BH8+Gy
FPQzYNEvi2sfprF+R78oN7VWfpOTsiu3wTUxF1CMUkGIK9eVOVLfZWjvRHb3VHyH
t21Pa+XrIKIx7gGE9ozbFLJGh6x+E/8QWhk6l/AORAmQQpmMK3JtlqdRL4xVZp3U
tWsdCtrDQcLyK3AEhoUJrYMmcgNMwK0XtL0dvqz4IxkZEo/rvRqcxInRCaiiZm1s
0U8offtiUyK2qrwHumyeOTBQHbZba4WJ3AAB5Kznoq9XuECFM8FDSk6qk1Vz/Fr3
eD3D4EAzb+e8CMxQ9jJeWZOl6xMVyugPrNxaDDef6hc7vhQpgzBo7PHZxJC8O3X7
Ot6eOE3HB6EzbV+nAhF2/BXmviiWclJtXpZevZluPvUrL0sCmtTRUW7mIcEIgqkY
+SgQU4fuy7zVUcU0/5nW94Gewi9YbrM+eWbL+FpMu43FuZPJXLSi+Ai5ectUyd4j
qBM+GNpUPJe9R088nBA3VYnpB6VVl6wxZRKzqTPaO3pK3he/F6y36nVYfnoBT2Zj
LWVzlfYsBVh4Iz1GJM9Ox/GsVNG2LH8lbE54tMKhkzBZDZ+fT8T/QJiPRVxVKOTD
rTar6M90cMgRvWUt4MsdRdnrsF0IoJKAxiEhK+hqceWHlVayfBiSyNdx0YL2Jeba
u0hSmE6k24k5DNW9PaGx35rUY0l6K0v3hBDGrSkF+GYC1Q+YmlsA6S+CCFusXOCN
ta7j705IEstlcNnTf+odLnKx9mPjprMMGZTzuHfaBi+/A3LtxugCpwb5USgvyuEC
bYBUpnsRQazS35tVgKLLDg41AMEL1GKrKnMZzo83WU3XNgQNTpEBrNzb4kOezoUZ
KJg4g1oeEs4w8DzRyxPhl0a918kaDrvygyi8ZplCmQQ4RJMzIh3Jn4S+YYAKtHax
ZdFwngKLz/fKmSyY+ENwDQnD+5eIIrXn976m7CJjy4dxyF1JJbX6Ho5vNhlOlCHr
nZ3F9TlRiZVIWgCsd3LcpgDF80OM8gDh4p5lt+T0bBpfvAJkbSfnMfpvmcAajGQT
q/3Rlrp4tPzrZqvjgBoQzLlQWvGGXPwXqg08FkQr3T0faQ+nDhCdlb+ZoDuNM5Ta
LWuH1mRfKkYBbr3c+E3Ob3t3tl5AvkrCAXg3hD23/xtbs+CjDl+aLJO9aroDseE8
8s4jOkCpAqU2MYyeBdCkK646JK1G8cStcENDFuhbw0Wmg4SuBJdUOBWzF0sJqlh7
PYLmWGs26qFvFnRHMkzGQvfAuR7rLpMdED/R6gkSxsH9bABlR4wqgEh03+dNwDoK
VVlg3XuYD35Vv2o+2y7zK6aEO4EFfpftQQFtgaFqdOVNp3xRGvgRijn0o9u0gSs/
/whriF7mqPrG8QoBDn55+jqa4pRCwZJYmJkm2PYb/KsAHTiQU8qekTISq62dI6YB
KBrEbmmm5ZXJ2xaRQJFGbpWJ5duAR7qlXvd5XDFsKlD2pA4YshglNg0mgYeNG0BX
yn/5dSzu7RXLCjmJlVVjTcufjmTYg0bQ+AsyD36/Mzim/1QPWcAaIJuOAH/8hsuP
MRkyeultP4Sg7koRN8XAmM70ge+uR6QRxT6De/Vxc9WsGCqgistG0qqDLFRWYKw2
sPoRSyGuazluGB8txxmzAdf8cF3lKLp1HiXIPeYC9A72MpyUiFQQNdsFGSqcmHCt
QtLNCN6QKoS93j9uZbzzPyk56pgZdHXhgWLii2X11z92SoKGfURt9g+5Bn/uzUo2
k35xVcERpWrVwds0w0hsNbFgEgF0g1jynuv1GfKp5XKhuwV/Nz07KHolAlGrSvkn
ZJmUU5+F2RRgsFEbZ1jyvxggabHSCarJ7qmVr9uaEY3cjonm8RbTFWjdURR0zK44
Kcf//kAw8uaZEYUK/56N5QYFRRl+gAOxMOsANJhDgCG8RinGhW4MZDhOwigbPk94
OmwsB6ey+OVdsq8l3cD789rKa0e+wiFJX0z9v+oQgYfF3Dh7NnuZYc5Tg4gSEzlu
BbM4Y7K2zFRAg52PrHgKPBJzLkY6q5xkHGPixG3p/5JasXOXfUSprVF4aoyzenaA
GCQsN5Lk2MrD0HQhDzCRbAFgsvRwypwojKn8MFBeEhtwO6oSwU3/EXelDtUVa0LJ
5k53j/PtnJv2WQSy3ntyTd/Q441CyinJIZjddM9Bk9QYmuPY9TogPrNiNBFKVRuB
vUawihOE+SP26JS8rwvATpFBY7qTlli2cjMiS6gf8es3MOgZfWskzcYRPeUDVLRo
luyuDpjYZKKY5wDBRb9OLaleHKH5xFuP3nCn1JANfvDH5Q5nyB5lNzjT5P3Q3EAC
0tObobdAIQYT0JU9RNsLJEMLyDDeXyx+9UpZItVX3avE+BlVGCVMvcLHnlaECzSZ
Y2z74jOEvTIDfToUc1feoSQJMUblh523ljjEROTaJuaADUlvxGWqTvDzQAD/LlRJ
Xs+hnb3OP1PL/PP+mFutCLGJXtQsZhon456uKSTK5EnDmktKVxK/ih9Tex0x1qL6
BTgqN+NvFf35+jR2R0Mth2V3F0MqL/rm9Yn4ZSozv1vWWYmwV/xfPdlO9kX+PTk7
HSIRBtu6HL3k6trq7TkvqXyAekpGTK1TI44v+BqLPmYBMdmLhazxilL2SxcP1vkB
sN/73bu7210ME69mLMhnvRs1ANSDdbAt0zaphaS5tAuQP4lvgJ/R4PgRBiOJV4jK
IlXp2rIsHCfwvq8RkwCLIJMmWDY8HotqMPL9a4LXt56DXK3qTm9YJ/LwqeVvUrV6
CPInP91epV5sfMGtKVdLSagbwq8+ODB4ReTGmrybb8zQ6iT3KrVIsKsIUlnCAnWf
QdHZ36tPo78Y81RI/sZAdkd2QWBWBmC9/QnUjHdlpCGFYcxdQ3Yhp/waFwQ7CJeV
mdSFx711CXN90Zngh45ER5Z4KeYzUG6dMFMoYNs2jjjD1E4anMCFqpVWD3ZJ1KBf
9XqgDBhpNlRHl68qMDyAvcAtHwiJREY+1DElDrFImpxIDR5H0q1eGCjPHvGpz3YE
6Y3Bi5nyohNzH0SEwtt/NGhSH6KMXT/4gaXsnmylPv9lExDkkalTwEpJZEQ74FWk
OBWythBPaXXKZQRwj80GVOKskVJVZ1GHBTny/URIrN1bykMH8VQnxcTLJ17rnrYW
2Vbw+DC9m1J5R5bzQwwt0LWZnj4hCpOoK26GJMUzQXPVa3te+lqJiXSuKlQxpgDn
C/yOJ72WblL7DyZ5d3P6U4r+FoBDb50huZ4SlJyl3TVLnXolmVb6QZMwua8AtQa3
/+FN2UqAfrXBRoxVL+LuzneUcAmTCFrnNW5dHZ8VJg64a0Oxd2S0phqsgU4qEKlE
izbDaNL94uwZVc1bmZg/6NLJewcwM4vShhSlyz1zwOk00jMnlcmcYPzQEBi6L+5w
47bJR5NSeqR40vEGPaehwZ0xUw4igS8ZlVVMrFyuUGZX8z6CQebMj9Q38YV8NynT
EP98Af2GPsgUHZxlQqiHw/nyDZxu1OpPeSA6yacH9ccW262nODIUx5UX84LSP6zX
auavGuSYD3A7IRgm2MhIy+2Kv71ggw5lv92TElCojkR1VQAhi++6dpFo2tkI3thN
0JBOZ2CNu1a0OAgooA+ZedwZSxpuLxskXsVvDrvpRNdI8TCMxe4ZXhblcPyPpoWj
ItwABFcAVhDaw356ynQE4p5lPrN/q6wbAM7iVj9a3NpGgZnLww7YgxbgQzjj8vPZ
fnJptgn6Ho33XDYTPlZs7FILnTqgt0t03p4VygMwbCnVNSYSFaoytvzphcJZSvZA
Jb5MP2lh1SvEv4v5cTlPji4UMABKSHhImK4UGpX0B0XlhfmNw+xC6IJLua7K8EUM
JV6F23WCx0rId9vA8j+Mj+Q9RPVGW2EneM3BAVGSZJhENjY5SFJKamfM00rfflg8
DMfN3bXFhOXHyKoHk22Az9AFaz861oVMFEvgqXs3kiQjAkSoVxq7HcCEN0q7v9F+
S3NF6uxl2XB6hbUKuOlRGzG6OPRauwSvMgx4J9fFEH6Z0sY/e2Mdl2XAy//LoXAk
S3ZAr85MuPdEjzaFMxLnlH/0TKUx/znGvYikmwdZJzQjszwidcF5+Hkzvpg2u3yG
L6rpILkhdjkwKluOMmbkEvn72bYqcnZh9PiBvzYLXtlsfkAvk0su2bNxoCB/9l9h
nPCV4DdcGxT4DVRtw/UK4r77xaCsCTzsQ1UVkSGrV9B7PrZLPcI68aintPz66zVD
m2XlluA+bfxRjB6I+CrZYIcDWGGRZuwDqCmFpaqBN6WzKoaYnb0G9MXzMckfYDMj
eSaEC5wG2G0A6B5pvVeZzDyfmPkUHEvNosbbfymagx8pBzcdEUfUnH87QEbVT/SL
eKVSi6NVVTW7XvpMhHbmj68wKrNbQWiPP4A2nBDEO5WxBH+gdJK8bCTL2cp3cHLp
ju3PzS+VQp9XNkboJFdkS0v3hsoEpNVXzbhAaLJRA2yY6pSMu/KLAuLK0Hovi1gy
FYZGv+gf3iwCi4mM7/n/NWCE6McRGepTjxzOq3LJ6ZZuv6Uzhjzf5OSIX8XkG0X+
UeYu6LNThrxixv7g9zNQk0TFoVTFV6cANNU4mUf5iUfA/g8eXVQ05MVAnYyPOMDZ
XLNrMmJitWHtz6JpDpPS8LVXhTkmQWp5QxsYDp+CNxw3NnEPqYdyeFnoi93TXBJp
hn5IpZ54EjkR77LBiB8Ij/90zuUgML5r66FgvyTU2zZ3pRrpe9oHaqQkXcOkMguA
53wj1VryZPGbPaNIQSBt8lgeGa7t8fvD6+c1gXpTZBQGmDK8kTiAQWgnr4fs4Tu7
vpEQjeHFGGQqNACTQKQ9605rPYxk0vjj/Keh8MHWOEykuiZc4wtHActPvpyegG0H
tfrQy7sTlhMThEDFRqeZb45GMIaGYuOtGMsY5IUscvLCTavpjjwke5IvzkyP8i+u
NxALPYORl2WJEkGQ4Tur2Si4R68zgxZPf//d0kNfwJ4Qv9AdDR2CK1TQudli1gjr
qxe4UOTf5PRWl1zmugtdwVyV29uOVAu2m3ZZvDoxfEpT/f2Ny9IriCny61ptdz5t
8rEoHFOYVomoSKKdeYHTTjrX0fRM0hb1I6XNhqBMJvpi/Br/+dALo1TaIqCguO7j
RYLDkb6yFcnnrFRJC7uy11KKz37YvmmRFeTtlBgBjh+hR/Jkr5ZlSZYHVeMVAALV
2hL+eCRzE/IWG1/C8PorpdOak+XDXaEqtFhPdeiKFlhAljcHwf+IiDFUEvyDKBQQ
dPfUb6O0z4MViqL+9wFCCtrC+Ztdwk7yd1YjhUWRT/PIsEvLpfcoZYlcm0YImRD2
c+SoOP78WCYdUCSXZQ9/UqrexPJwJs7XZJRdbohWDyxT2t9VOoVPBGjKQb9KPzC2
O5MVDisOPpP9vuetN7fQsu+R1to6KsEHijR0DEk4ss827wEOx4lUnhrR1GrCylNI
BEBpFaUMTsMyYOKHyuj66SDRnNyuJ9g+4Uoz80WfAWrjqwqNWeE44ZLEw0rlLsUn
0fjIF+iP1V6NdiPDposxCsm6O4bbqbnKWqe9U9PU4CAkoP2bmrYLvisxs0PcoqrH
v334cA+NuyjqglxPBWyVy/RTN56V8rSVd4jnrA1VdwxwJZuJRxOTqFLt2zHF5cg4
wpbDvg/Abvto+x+MrhaZ+ENeRU6DOUOXJ+nykpkMyFLkeWpssTyuK6Z5JiLJE97D
coWjo996+DCDD0SCl5jgkfJKU42czt7I9mSvmmNshbS3H9wvIpDo6u3RrfUh+0PF
biaNWAB66IZgrdKPS8q59UVVt9ZxPAAs4Yg6uXAyJbZZ8HQdZAL3Qe599+PCq4GV
YMn7NAmzQS0OG97bV4mMxIXajhbPRGrFdH4w0ybTyVAARIqWoCbauymdYtl2VNYz
15xXwqOokfo/ueGRVItu9jsyC5HhNTzKaNoMsiae96Xfq1t85HmV7vf93G+HPBeV
ZpUg+jUgYFaTMr3YLjUpyNemYAEhfVZ4JQKyHaeR+Wla3ELnlHEDpHGBwX/vOoVj
cSb4i4gVwV+bSaqNKGWiQimY5Mx7biIqiDUPK2FYi16//X2GgwCiXgPufV0iyrVE
xSUw73IxO77vzXSb/glP7GFEe5W1Tuj/ciOxUHxjVnBuhIkIOLh2k83gF50LIAyC
RE5KK4NncG+tuThE6gL/9Jy5ytw25R2U/J5RbQ23voYUJJob8zbykQrYQyMOjvjR
O3dLEZYWm5w16C0wJ2zLb0D3jraklmHGhjdMrskIR9ZFl5an37UrY13O4tu3YB7J
Qp+sX6+TGrq15zLwuCEWUgf1K51vVo70KyDv7MP5QR/tozEsp7QyCAq8nfSbP9TV
UfUz5aGsihElS0QY6FVMtlSR4fihyf1mf+ygJ5gZTPuVD38iH+pj90dKMwuqTukO
xYFMFjUhtR6hX57Bv+YhKtuPBnKmKMnYOzxqJXM2dsks2vmWHmzT9k0D/AqnOHXP
vFEFJcIB6SOXo0moTZw6CmCtZM/vvhVhKitGdX+9JPsRwLlqa6bq/kWy5HCmIN6/
LbRwWJQ7Nxov6Y0ZimalNBDknPqD/sCpVEV7a9FXow2ofdPu7lRkDKNi2KEfBRC5
yMBR6rY2sQHDIA4ezg15PqfJzjreELFFWm43poTtwDyp/5yi0byH5muGg//zh2rV
E2NypTFNfa/mzgpEbdpHW0EKa/DNLCD53ekKbQaMDckhoaWXF4ro6z3s2L5wqNOm
lEQLszPB3w+Ev2g0ZI1djm2oJrGtgOhqwvMXkFzupLZxkWEi9C5WpBZYmZOUJ+DQ
ue1Gov4qAGOPSEIR9zXU6Iel5vRiz+Q2rvYsAX2AbPPsfyP+rQleyM/a2NrIupuN
7UZRboBn7m0BE8/s3UokfCenQbZzHP8Sn+G5Od0EjY3S6kxL1qiHHq1eme593BwP
TrDUt72cdccPkV1sjb1GDjQTtWwcn/lsMovkB+jJbg9GZ1Y+xbZdvfAc28AC5Utp
S/of0CTc7vlyPLPAaG3nFxZZqSjI9fc3arWjncjkf4rrGWvFyu1YbHn8EhRjBT9Q
Acb9H7frd9DHhxy9Wny/pl+hGDXICt7hDAOdiAeF8zlwNq+erGunzTT92gGZWz1u
FsmhRof+BTwF8eNfTT0Qa/qOk1ITaz1s/NE5KcevmVcxQ5vyktwLB8kQS6f0vokI
GJ11wyVOMrJNUK/B1Ag9H+e/Fx4FPLNLgj2wAhGmM0ardAUvUXPz/pKR2pzOKdWY
vd8DBjdzCFK0guUpQprbZQbZxWA2adfpKXsDZYBj4GfJRUBGllfKVbXuw4iqRQwp
gsj85qjz2yWrAejGlA2LEAZjKXf7t8+0RjJ8Ebmw9ouRAre9UdulBP5XI02JcHgA
KSUIo4ZYt0+XyDKOK5CQ25Dw2EStNf+TuCoA0UD1Ha+hxiSYvZaw+i7VaoKmFIG4
Lmk5VlNmp+/PvBAwKi04Xd9lRiafgsQeflFwBNLCixgttN6lBiXHT7a/aZKbMCKZ
1yxbITNR/AqQVCC68jTR4To1Do6zuDahZ7+5WRUnAUEBnY0hxC886r3mQApwmTv1
EBo0+3m/Ywmg+ykE4LPy5dcBHUonf0F9uxrlb4uDvweW3HWOTgKirqeigd/uFwB0
0RoyUwzEVsp9iad/5nisuOQ3eGRcQanhbvMba1BDjQj1RZ9KI05j0s12nsb3dml7
3Pidp0MSElbYfiDk+Vz9KKB+SawN0yiXo1QSTgwNgeUByp2Ud8tnVPHV2YxuqsCT
y8FnlSoAWV6yJ5nzFau5PG7WPFSMHih99yrXkvrQIgQaJEXwMIvXtTSdVrEUZ4SL
49GqCHgt64p+J8aFp5Mi4rAietu3T/BscJaFJm0Ygd3JFCCxzf8kN/RguOklTzTQ
q1+XynfY5AvVSejHnt3QWF+y8YtBZaHXQtldXHzEDDC5AGJAebG3P9X2aTgq76CJ
QmFZCnCyWBumNTcQ6pZ9nG8L1+6CfKSn7zVv/X8/AiJEWe7J5ODVZTf3HZMWX082
H18YyJejOTRg8CxGElkREeql6UT2gmnsoD6Fm9TpM+5rxhraaiqxBcU5kgkdec3B
nFt3/Q77nK+3gm4RShxcLsXESuFGH+m6Zi7+8vtbd0psb9FJr3AU1Wu2Eb9f2r8e
9PESYaB0NsAulAkHhqSC0Nhhyh/4mb6xnhnJyYkgq56nVVoLfyQsPai9nz3oLRMK
HV9H/H3HFzXNubkGLGEYY5kiqsOrnIrAae6eocF4Wj1O98s9kbEGBt2ROhyAMI/o
Sz2HoYLtjqdBVGqFyudKnQvC8YgQsCtLIEHe+7WIb080FgB7gCt0M/XiRVL9GFfa
B+nVP1HbvPeXO74oIncfw8Y7FqF2zYO8IsYi4XjOBsV4wtCYqGPHQ43Pb6Xgkckr
VkuFlmidykcyK782SmOiPGfDW4ci1pQXQgUhKg06bKrcD4nMfEJGKai4Z2p7CW3r
EJpnXZG3ykVxmQ9v59whrFBjVFL5FP+uiPiFoWovMrQ0ZqLhd+xrMAe8Fm9ZSaAa
v0CejyIgR+j7OKCYNaHXBAH2pVjZOTCA+4/dNWGDxrjCv7qxPw3niYbtHygHkBth
N2phe5JvlFOpss99FxZdzXx5Jqhj6R5frzpJMr3Gs6ZxgEjHZO0GQglSIRDF8kaV
hMaKK5x6ryhJ5ejMlm5S+BZPd2g3Z4j+dRfXp7F32fPJnk3kkfda1+YAtJTeV96i
o5GKIPVaGlt7HN7Ireq6sHHLF3VDBpafYW7WMMp8TIApO3Xj+Ja+R+eIY5dAdvYj
KlYXejkZkVAX5+lEFVfstL0NUBzfnccL1XTl+k9I+M8xAl0isM8jszooafzdcM4t
1NFgVP0c0A3gBi71eERM+0GwH/fNlsMrMRgw4l3vyZL3n2g0Sl2eiXY+lLL2wUda
PKqTNjXKtsyB9EBFKKwECj4hYdyoaXTGEgxvsJd07XRmIU7ldcWayNNA0WhvNx0S
0brEv7aA40/Lg8c1pCAoGK8UZsspC82qkkcbo3nPh64s5IVoPEN0A+x4qMR3oBj3
7fWy6T40GxziWX40deyace5y/ALAlpX/eL+IxYqfaLXi+udVXX727WuDYm7MQkaD
CgJeaMYV+TKFrZLAGjrgbabicKhbJ+cTE0ozFjtOvv2I+6fNl/LLjKfVFdxC59TF
3SOWRo+OD1AaIQ76SsjP/0M/k9rUSHTzcRCwZpzBLVKKqBkMHWxkE6x1qjswsjA5
nJxutUDuh96G6m4mmg3fad3GtJnw5uV/rwSQIR3VpGcMDaTyye3ls0rp5dpYkr22
kUpms/xk2/FLg4miwYqsvjh58Vq3SLF/960Csc7YjCNjcbyCftI/mhTIt25xOBKl
M5MH85X28+G7fz0jk4QGLgdMufVDvBsK6ga9dl7ntv6DNZe2y94ng8YVSHrgQGfs
gdVC1d/suAVRtxgwCcaL2GsPcBij6ah7kTV+aE1N5c5T2L979xQq7cXpPJH5kzYv
w6gUG7ECSi+l8IVdec5lDn21JG1Bmm33QeNfvz6QLeJeqwyJcyEtAuHWcwrBmvlm
PJncozNfxU2LVCFIshRWdW4wqGgmtAuX6+31dSMxWhBrpVK5bspUkPHfFc23X7DI
ASd7rRLb8/a+fOfSY64XMAb0+vDkpN6UJ5csc8Acyi34+9I10VuFBzXIMjpMeXsO
z63j7uSpcI5IrInFLEPCtAynYHkOiFD/GpE2b0pVIV247qExqxEXlxBFGXJlDOiT
nBScCbx0KRgdwTVaLoMYeMuQYtl7NX1RjfwlMMKn6T9CRfuMhyACHYqY+4VgVN6w
br91lj3Bcp/CyWA7nyvTn9i8Oq4NyelupPYccMFUQvczzRYGkrXoRxo0rN9ITGsA
1Utr53b126cladRa6b7AFdSOcsvowGPUmxMqyn7FMYeJq2fLcdnx+e1PVuJdDs5P
DqrQLQUYpLHDCHon0XIC08+Gzy7QRkOww3QhWXgQda7l9xps2+09Hsit/ejNIQS6
pc4tGjgRzBi1+YSJFh0l/bWlhoDCievucXcL0+ByW5Z3PCMwDj6Ue3L61u8yOyrN
3htq5MKJ/wl6z6nwFOYMxd4o2R34UTwrw+a6QWSpjiOpmYqVC0E9cHiX1PNYqOb9
Bd4sKRPOl2xWrJ1bQZa3uqvblHKOhjxJ+SfubljW4fRdgnzyDLX5Lczfru6xAfLS
eyIySDas77+HAHC/Vg9McoeG9ZXYZTLbNtRoBmgZ8dAXUYQTf9EfT9oemglLOm/I
huF7wT/GMln8fEmR3l0b/WJw4Xe5TuyTZzefMVlLQDXg4yCgei+jKSBR/wFBBkjh
f/USPkQqUQ6/1YtSHmY/zXy4i/doc2LD4XIyBCnLmTMU/pqrIy4mcGBOgSwM5k74
k+R/9NRdvuh8zOWNfl/o5CtyCPfTD4BBrOphQJsnz2Fkt4lpxVCUsA1ZfAXWS4Ep
aVrEJbOm2LZzHbd/N42Iw0Qi32J0Ysw4ay5lX2nnvZRFV+GEGTgT5nznHvCnvqkn
ZtUfWawRibQfif3zgYybnh9gEhRsO2Pnql114udFCiyGmrl8wtWiHcz+GEPnO9Zb
UBB08gK8fFfFrgDxh+3l6s/7uYuBI3F52vDaxOQCINjwpILO3KAbI2bb8R8VoeMe
BRis0TqZApODACSnnsc/JuW7zHvD07FkgOPyU6Aw77pPF4T3fue3dZ5zQjn5Oxre
pBOoL9lKo+l7XHglRzCuEdo3nalW+VVZ6PrzQEhCfacz87ApfTMlaY5ng4pJuaPf
/zBZStsUKrAs0ha81IRrQwUSEp8NyEQNvwmNruKJZl2phImZbh7+iX4Xd4Xc9P72
xXzEre6Gl1k/PAz75lnUA3nIGn5Zzdk4zVmD5nAwY8FVcFjq663LVcyaOhHQaCuk
KJRUd/kX87n0V/kjMb0cVhvMcUaGPAvHgJKwX75ohSMVFAbNrDyXUE5re2yuZy3J
ycaf400Rxv4I7MG6apRaE9MSH1ImO1+qBaLB8ODAHJWS100FLbNJydYa0Vz8W4hC
z7NTrtNTLSC3/5OMaPOix8yIS6+rZBJb1IKtkKXl0OWBHbBvNJP40SHg6/vDJADv
JUkCh1R3K5ZsxM7M/CEFt8NQyBPA9LbCsZQX7UsutOXBDSOjZeh6W0oflXOI4DW+
zVSmRg0kSOW+R3IwEhKgD8EdYVznO2HcMwi4zrf7B1MEORhYwgLXAN+faG0I62yj
B5y/PP0yDMploatEnTaYvwIvmDP6/WkU7cYjJCE7D0UENbPp/yZTHyRPJ5L4Ykct
Gcr/nJiRa4zjoUVaCF8k9hsi7xwrzI3UE1L3OMjNZEu61huzTXi9po3gsxng228o
yEtxeUp5tuo5fva5qmzaMy0kSb3uwnudq000TAJ6Mwr+seCD7HkRFUXjfN6Jdn2W
bTimCv/s3wPXoSv/srnR3h9jt57FqqrMdMUS9001J3cVE63TSaDoU6FBRR4VObfg
4NwtR6n8QizunKDpuCi+v8OzkNf8IUFNWvmY4isPkvI4kyTcvVl7pHopEMozIyZa
5mW+eclB+xCqujX18cDAAjgPR9jY3YsnVfIXZ0kCcSMLakLo4wb8HJCfhR519kSY
Q1nUgY3NQrSRz66xOHWlj0O47uzTaiAgWG/n8+d5qPRhbeIvIzXmwCg1/m5tRl/f
3ufwkvTWa948fN5CDQoaoy9WHQNp1GFyLbdzkReEXoJDAMXPMVOp8t80R9zs6Lgb
arzk/Obuxfhp961yTzfVoEAe+/MRL+r2a9dFMTd0gmx3HIHzkIZX7VwSd7NwiRqe
igGgnjanLtE5lK7KjsH31IjMs9sRWmEsIclj7pjC1zad96qx2FN5HQAXiMRim4zE
2FdMbx/WciaM4KVMjcXlOXaSq6NQ+aN44GwhjxlMEAcDOhMxFiS/N7vP0iKUrQui
t05uoXLyeF0oXzU3CFRZ5CVG8cAoigzbDCgjNOEheXFmPRVPbrRhVhb+WFewS1iV
ImRfeHjl9/qsSIDwo7fea8i2Yj/xTdHG4QggrPEYMBrVC3Hj38uCjuPejBcDmpLf
V6WoP7dTPi7hXVTI+wnF629cBtddL38/3VN8qWFN6J+MzrUvjMaCIH9zCPoM/2lj
k9XX0vQ5NjwCYsc2m6rmNM2VE0oNMeUUx+HcxLCOkKgB584gcnNIqd9iN6uFk527
xBWg4oOzDofLiXcvlU6hlrwO6IYCXVSeSDHdiYIdgOiDKul8Mn8pQADB/AmSCBLx
S6C85TxGtdjqomE/omIoCXI7fv3vjf0m3wf5hi78Bnb7W3D7ZjnyrHq9mveRheLV
SkFznBUycsXsquxOI7CWFfoZf3dDR/8vKP0AtQ2T4KoCdWVPdC8yw4Ft5NvG2c9e
Vba0Y63jDc+BbtW+85PLVEtK9q3/i3R9Iyo63naT3KRLhEo9DHFzYr9hB2tW79S+
WUSxlrb+wFUsbzPWsuCoZFW5GMUTHVOU5SPBBDiQTDCU/qiAp9jZhm8zXIajaDm2
gKGbTEaWwf+MjQmV3UQEZJkXIhFaP/3g/9y8y4GehxJWOhmJ67rPhupMgXvRe0ht
T9ih5zTBfVD27jGhlQvk7KED/sO1r4m0tU1qlDo76HAmutUot5eYAiRHDqqynoDY
7B+6tc5Ar+ZmiZNO1Oftjy6Djb3iLS0pM4khl3pzw5zinJUUy7Ca3RT68K49u7h2
976I83FsL5FBgSZSugEUNxuEsUYw4ll7ISOX0VHP9teJAVErDBcorDjAIpVrqhPG
z9J5KHIfg209E5etB6/+pxD0eM67QWnuVewfa1LXbKo+ieDX2R0YmPPBf/m+2Wtn
YqYLlDrtwSTI607QH9OK+exNkDiYDPg2h2lWt/YxDOJzEckJisV6NWnFsZmZa+Sl
9+oVcZEH5ZTO6svoBg3x0dZdgrqJB4WATYg+Dd5pNSGWfy02Xzb0XWkyr2RtQj37
H2X8bajHaZ/STp0TVA4zhtqg5jxBGfSlur8wIJlH5itedqgzrB2VJIF+AgcY09wp
ktQmSnWRyDcZjsmgubr1F1U1Occb1eqMs9i6Af5jL5r5fCD/MtGvOltb7Zrs4f72
Z9lZBwjNCLOlziZ2XknbV65AuNdpg5mo/V0CAHqls+SRgwPgIH9HK2XihLp4l0nU
fcgbHtM/dJTNJCsP1fbOXbKIm4fpHghrr8IvhmgglggpSDgoPYVFYDASS8/cqNKg
CMyXyEAt2yXPm1N5JEmWzXN1UYKrygdOWbOW9bDkqKFLuXzJB29fFQvae6Zb9yEo
EGx375Vbtfc3mzFdJVS4uTDzTelBAMPHUkbDUSFZMNmS0rgQSCG0H7+jTvvQmDsU
MKUVazMpSvvfASYYKi5vRJe9OhxjPhcVfmzaQDBE4zUuuzTYFusHqfgPY0MSWxOD
ahQ3/qi8fXOGr3+FRiDOVLtOl9AE6Yt3Sjg3AdWTjbPMPAANc4ElLpM/l85WKOG9
461AevJYOclqzPrD8lwnfuaWh0FiVN2z28aau0YQ/TldMfo54dG9M+jUpevBrCV6
AO4OtKkWVhAMZkSnK7SC9vd+IUhqxGGUtL++s6raog7R+btWD2km2SIDdCW7CJY7
K7ef4RRnQz8j65H2z8FP9WtyqwbetIFlJs1KMULKT+Y=
`protect END_PROTECTED