-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
28ad2lOYPy04p8/GU/J8PkTZGCmECxTNmNWIzLfS3Vnyrdcw9YOpSaSGgyZ9j549
gze+1HZ2Z84JMXYdOta0Us6FuZZNGFuYCim3M782roPFFss9kxsCYNAnDvrmJzkJ
Tc9hwdWgjaZ2Cpl8lUlJoLcOKk/ziL/FtFPFZRUkWvQRyh/wAci1Pw==
--pragma protect end_key_block
--pragma protect digest_block
hj1GiZfKNnwIHyiQnvchGBFr0ko=
--pragma protect end_digest_block
--pragma protect data_block
Wp58RmbMx0MZ8vU/sHidPv0xx6bhMKtNF0KpZ3S93X+kgPHZj4XcgBUcHT9qK1fH
/7dmcd2mChJDHhUPvGDr3guInVavvx6gjsAhV1QNIcBvHlQx5hlfafaY808VZTcG
Rz+YryEQeK5s+XYUZqk8BTHjyKLO6MskyIV2addz+BFzajv3yRYzyN/0BNMGVWAW
SdMm8XWcGNIaAGHImhmA+4Qd2gX2S+UQ0lU8TGXXgPzJtfe8q4mxArXlLv8V1B6G
PzyvSkOQdoD9r3IRwyFkijTCRPGrIAEIgZlPVhF4Fu7N2CeKXIx7mAHleujYrzv6
IHhQMXzvBhTkXl/joJaTTfnsG8ZxP1lmCJ7aYFEaIZHBwRXpo7yPjvo18g1r3tDz
mk0bYM4VUCV9SFRTIwGaANOpyFbGzv19z1DOdgjRDwHJQP4qgSNbknj98Wvact0L
cp7I94iMY3vSR56eSk8IxIN3Uj4LrytmsBJGneIGFUUvGfRyVUsk25196OPd1qyy
5lf2zzt4oQjbbz9uPzRlZ2qbHtuMYWdNGil0KoA0A3OsmI/OUol0BPYKY6kNLb3L
8ukmWeOER65eyJMn6aMFmDZFJW67a+lDNRCgKmmbYl1JTUBU3mEsSa9DwAjvYYae
wXo/VbuvDrmRWPyuuzj8CYmz7Pymm6jKQ1Dm9x91s3OThUA3s210lWucGTZGAC3X
Y1PcKCfYkaLhbEZpAAV4Fj2Y1sFwGaoWV6MnI+OsFEGmCzfX3p8tLRJ4bc78IPWz
YVlGBpaE9QN/AowxHuHYmK7CU4BjQR3P7axKKUCkU40d9uKAV8BkgcAgxEpTAx28
a/nYzo8l545Jab27BjGWYrKQ0+fJZIV7oy7jDkS/GZfCE/2VNNl1WingnrY6map5
OKloOMMtDIUY6ih0FylrwBc0WEaLImfzHZ9y881QgeRfYbwr6cwdNHlwK5W0+pzM
AgM/yY+R3YxzeJU2A0QNTJlOGYv8pHIYj+Yc07jfk/9BVbjCPo551pTsTgeJ4xuA
+HfIk/exHkiphdCvsQHZsA2R6kdIEx401yWEvLkOHEJdoKb6NWmKRN0ucmG4brTL
VQpMtf9qNV4NIGsMt5CQqkN2VC+neEWO1an7F7GXWwMd3ReNPHDc4AI4eh7wsiL3
OuJUhv0xUGPHsFaC+nb9XmH+D65VERXHnFyC80GXE9LoucrXziUGDVTY2DwjU/Ha
LV4728i55ZQfWBS3G3Lcw5KBHP7/v0KDYbCAsCrHPvH1NBsbkAy1TO7nWIsL+MH3
9i5vzhScLAjuTsbFnbS4PRhR5SFM9O/np4ztPDH3u7FhTRSVfnscwQYzqEQ7NsCZ
iO3qNLX36tOpMdWuHOZvX9RWWQws7NgOSM4BzeqnsEPk9wLxVScI+KUJKhqGrPyd
HRNc/6USFc50FX6FmbMkcaYSpCXPgzkm39Idt+uA37ooHNKKA9BozACsfO3iqMZp
RqA/NWhm8WS2UblklY4ZIFT0QPF2QuOuc5043Rj2ke8MfSm88fsZE0PFt7XxIHSB
1QKcJQEUDDnoUVutFEXplDsqaWYvr5Xi+/Y1BqTc7IESSjvWhdyjevZsYr27QO7S
rL6g1Y60EV+hLh6ZXI8OfzuLQfFJ4lCbbDgca3PKquSYGk/A5WFvgjH4w/9LtsGn
NLEngCK1X3Cvj9y04mf3WJFGN93a15rUf9xyDfea0hW19ULyC1BtuJ+CKw5BD0sy
GVkM+Ha8Em6ChZENCqmqFi2QvGCIYBfLwsTtBvWkMXrg2K3aZLb7BZrZlVnsOw55
/hbVk6GCw8o+YQpigZyn6o1WQOfDJBjNFkW3ckpY4oOt9eP+NHDZIgy8t/EvB6S/
So4r90xauewOq75Sx24AzTgqA5eHzdZ8mwrVGCLLSAs2qh1TrvS/K7ze1tFBgE3F
7GHhT0LFo0mmkDz8ggByxeXbiZc9AFYJgle/i7VHCbeJ9DTSauYplOw4h4oiwccj
fiA6NYQwx8pIjA/hdeJ6ZfYUO9IwXo4wb484EY++QdNojQ9VPcFuAxcDynWseOKt
KHpxY4fXYDeGXJsFDC47xoLGzF5K3+UuE9ROia8wjI+DPe0a18iB4nhFisd4PUUm
i8u9f8HNgtKl0gza3X/2OmMjqSIfToxttrGx9iDbDQ/qWb6LHtX+HdtqKhP8oLai
SBkAJkDYUtPnNdZq2r89Iyuqxf9cXpq4RNv4ZqI3L66f8hnTUj8+Av7UGG/aueyQ
lDqv17JKwG7r9wd7Ym717Z8jz9MOwTnwUg4HGT3EsbVIuttynb0SxXdZ+saJLmX3
FQDos0qzbbTMrgeGUmzmw5PQLVGpgfnYDdGP2s9DQcBNSHN9fWO89aSgmiNXIGoJ
vjwLWmh7N6JFjjov1QgeJlOn8+5STRnFvmgTn+Pum2P9r5dFvFTyYYNQ7sZUGZjn
spofxBTmq3rGhNDX8EWpe+jzN87IIE5WNK4XjezFEkpwQIjIocjgtt1NyQfsdyVE
temB5K/Dh3a1Ae4u8Kf44vIt1P2t77W4lj1zFk18AjzY/TIiF9kAzY+568bj0vaw
l9xHOTY4Rh8+jTGGqADUVzGbl5Sv1LkVfutNwix9d9znwiwUmXbB2bfLvE/89qcX
y1Gdordnu3lfnV2hDPt+6xCtMnDZ0eh2NsjtmCZFj1/fcGC+BjGSDPzJRbqE9m4N
PM0VWxz/H9ex6IYpPXiXSWrRqDXAIncvIZ0GgVpTlmWLm7xm+4xdzLVqxD+0OqbY
rq6xyul4UoQ2AgxZXK2OWK2G/ploZR3F87GrVJ1K7xxECBQpuaU3IZNJL+BGnj34
ktM1X/9/26Hk1A74InBh82rZylaEdryVWTIapZ4KWb2RaghzQVhdmUTQ4zlnFRob
N4sqec5oaqJZ2/sV5XCzqfcmobK5O6XTAYLIugksSmZAnTE54JoGI4ZPbnpPUZ77
1CCUqxNlLAk8lOpJ3qrY0shY7WRNUEi6LR0s+9V9pjsq7jYeU1h3EQhvIgtsxW0w
mfh0186OVQMGi4M2yF/4BSubJtBfMAuNupK5cUXsFa2TWDS7hjUJXyQoQQCiOr8m
wyBYixSER8CcDb5tuekIt1f8gdhOx8FR+3I+474IYoRPF0i8CH3geRVARp5voGx0
zDdOZi4WF+REx1nVZXa+uxhimxTT9GoGG6XtmlJ52WYHQyLdUQSindNm/4erkiJP
1eyRFJs1Fw3NH/WGgROnYueCFFxjm2jwlAT8bcB4Oexnt/amu9roZs7fV6CNhxx1
F2hpkVhCdEc5JX3xFi1kgNrcYELOZIDf8MC5U4adUg63kPtF/XWSZfax5ts3kAkl
+IEqOpROezGAUe5XzIBbzI0q/d2LSOUYhmtoemMhuMthgOc78FzoyjCgSXihm7zQ
OBEBcyjLypheefntbdt0X1gar33aYgr8ybOk/5Vldz7VK9TfEpD4VtyGoEjRJnnJ
vvRUgaQIn82mso0Ni0gQ06l0Y8fWutlCHnjHJQymxZOe1extvzDhQ70GVlYNV08H
UeIr08uimLzeUEKW0QebqXs+X95cpEjzwRON3cEfGW0GKYBOmDmGZb4nhKaLcskQ
j3l7hp8g9/nvwg7oZXcGf4AucNNK3+hzkGrf3Fv77bBoVCIn3xxNc5pga7SEEmsZ
e9YtUCoBJo05qCRvkV4ZyQKdxQchI4dT0DAH0miRk6tCPE0WbK76lLSpJWkTETtt
t25OEHYWWCsOow0dVFCApzuK9x0nXC+Ea77Afy6iGzAWZVCSYhwHMNZYUEKiOSd7
FG5ZqomsQ4fjUWoVb6iQzrxRlWkMYuKPBH9j0821I6Npi4AvCmzOLbEekNXLK00R
kWu94MhSgzqd+IV3R8j/ZOxo/WryzwxYKTX/1XwNalVKW4F1Avq5EcvZBBSajZaR
9kW3LBlDii4NgS/zewVkJQCxbxVxJiDjvtOQXUxVRmylYirk3SN4Dm+a4HbRE/Ot
X+Rth/3L23PrT7+hnwjZyKI5TM5C9w8vJ/DyLpvJpq6rBSvHmTLpyc1XVrrHZH40
YLC8RaCmR1lsA2GvN0OzrqQfM3fSVM0D/JgWl9NeJVRdAKkh+IhpUVkT+uzgg9v7
LuXzxlGnc1kVj3E3OVrFruT949L4FPkaf3OpyPLRfCsoVWeJ3Is62rxc7i0NxAiW
l6pMggCPNT5zZq7/fl+Oek46+nldOPjQhVBlyxDm245m1wiQV5Bi7nnkdsDi6Cf3
9a9eNKaWE5aV1cZ8zdXggsrhgdu+tuf4YDdS/227A6KkmJAaPB+z6w608qHNul10
ZEGhPuRSzZL4SHHK+nkGVGOOaRi2W46ItraeN7B6EvEbcyScu/V9CCJ37bRFsETx
0LDViN6U8BxkX+044ngXOHKIz+vqsa5/x+ZdYkE3CYzdfk6anzbBrkb/Q1Frk6Kx
jJ80LcGHLCRn7kNiQvc1gpmpKXlEC0FrHv8wEpbjnwTxwFlJ4vzmu843g6V1dQVh
7HDYUW89CvzCm2gb4G7uJ+8XCliGsVv9bOTKj5SBeqxrhybQOECuh3YFhM0EO0nT
ICQS8qshrhhchbssTwOq/2v55VDOnjCxmMUkbQCC6qNii6Gw1Q/lhPcx+DNUnfev
oAr9z9a9BLUYurJIFx3kBmNqCigg5ObUKPNfPWk+GlQLIprf2KZCg+Za1jDjJd8Q
jsOdKtXa2q6Q2acO8D2yV+O5ns9Qk9BUxNJzIwwtVv5Ar1tZ8aA1/SWVvllUIBpN
Y47RjWqr7dvMNTCptALNaInTHe3j4Zno+XrOPX4QbZVe7CSf65qzGtNPPuBO6V2I
rKUn/fksOiMguSoe3x1JOPQ8gYQ/G7OjS6fFw3ysLvLl5jEG2KyP4lY+pFAD3wEO
yISOZKmWkoE3pSRYPnz6/5Z9d7kJFoWDH0yw+dIjn7gq9LStHRXJOS7rKe/foEYF
pA3AHPGJ/HDiO7KspmZn7Zz8zLOejbrvBkf2q63+/01Feh47mLenJuflwf6kbHHH
0ouLcjiOn+dJD4AqNert2SxAuA59ZMGWM9/6wdwzG8BQ+yJFwgdpq1BON82hpacf
5Zt2LqnDOlRI8oDbweLU1V3L/0FPPjQgLdphz4OJbqMTiuiSyBbQ6Wln3qqC8unQ
ZfANQ6kAisCOZh4V+36Dshh5y/FjjuX3YUBW5C954LBMV4wn9qSEIjejD27KCgvX
yX1jvill5UgNaPSOFnCywJKXMEn+TeiloftlKrhT4TNn0oqcfA76lYnQ4ah6JbJC
KRy+tozA5V6H6MJaYIZH//hX4eXaec4M6fnKMgMCngJVseT/Yu9b354OreeK7FKl
BXRItuCNuixcVvGtMMyQK8OgK0K0qtCsZFFysPdTuYHZ2AHYjzmxVSFChd7p0uhC
5l/t7wXdsLp91/gGmA7ezje7HVkuxaRLPtmTqppQR6FllDajf7VvZFHhZaq/IFe5
lMF+dPyoW91eHUBTOBjnjuQoIPezSPFDvrUcy48ggmbmZMFrbP/QeQP1tYEwXqBT
6OZAo717HBXDKanzEY1Clr+ljNTkuOjKCcXORaH2hLyG1gFDCl1a5cncpYqYzW+J
/hryx5aubThoLmRhS9S3ouAEnLtL4AwqXEAeYUaN4lxXiHLkwl+2eYG7ltOM4xXY
WA7DMNSiYnWMgKp13cN824xKY5eW22I4U8DgArOPynUPUl+CzK6c98sQrdOCUSRU
JcPicWzijPNYG8rKmKNEk3ZaUPG6FBhob+vnZbCaPb771VV0NZhGeNXQSMaDZntv
IGCTGJj+SspIIrtwwKZpJxhxpB+oMGvvFPAM4SgqjeihQd7K4ougI67V0IkTOrL3
cHBe2pW8E1Lw9ptDaCJqXr3dSQvW1tINq/11pASrlzMmhPVgua9c0skTjLYfJlDL
JQrY/jbcN4QR1iis5TsuwlInX4YrnHeMSlHOO+EoqTQb0BYHUGfWH2g9id1L1qYr
TDnzjAo5zlqKlsbtqEA8oeA/mcFK5NsCU+njV29jZSAz55Dc8wB+LDIAg0BRC8Mb
PFCcUtLJfluwH0yEuQotWpAnko9uCa66hqKmjJUv/jAlVKLACDOwrYl6WGkUlz/X
5B+rUXAEz90TDcD0tB4FZVmP020ARuoqrV+9X8yLJSIrAbH+sWFq0Vaww0TW27rg
SSiIOkUO4mOWiOjiZlRuTZTx8la7viV8t1xHoiQPA2fT9A+fNIQCb6h0KKjdeHc2
9fX39yscRnaA1y48jM2dqGCHWSfInIDT7vOFB9O3IeD1sde6njr+UnMcbbLkh68J
Arwur6C4GTgHR53n8gCDni5LdNDKGqExj3rxawWzv46Xe/ozAvcimNDraXN8s2tH
0N8s/EoDGQcMwO1eoHQBNC1KBCIX0uxF0UxvHP9USG+vbMayi1rx/0fcm7i3ryU1
Hv87gEl/MGXwO2aRorewsQeP8BXC+3vqEQee44hlvLpN9odkkrtmsVikxOJJFiGa
gAPLtA/HopwunXS+nocBPZfnstlhg8s9X9uqHuPjP64nk9G0fI4UaQPqacNZH3tC
Saj/hKnSmIKyEde3qQg65f50wXqZGI1UnSuG+yZ685NaL9Ii3PJyjRBNA6O3AiS8
CH0d5hU0KQz5PEwRp2rHaTK35qT1g5C04amijFmB3kK3MUmBrynVJEdXg/GNsE4J
JAy/ALCfjvyJ0pORLsTGy6uKaXapDLCSDoqtgAGr/aFY2yTdTR8e38szUBhzzLc0
Z9b3GMqbp8SIp9tZgwVKA+wCeobHO+AXXvyzsrRZBA6WQHkkB+VRL/40WP64sJ+M
A5JsGUz+maQXtgkkfbJ3ZE+4K/4GFWS+I9CUNrvEIzgL2M3GzWQbpqTu+GZQV0mm
KjDyyDbXHgBessRrznMIrW20XZDyV1oOaktaQVt29q1SGcvcc4+6OisyNzrqh9/8
MkRK0OP+CMr4f6TzwdF2tShHnqMCglU3mNFxOXOdgVNg07zzukUdDT+ARd/vgDLy
YNo96LnywaiRVyoyOAbuzhCn81VG+jllsqJgWzMS8YQn2sQv0Y+J+SSJriynwRAg
Ech1b4DG/2J9/iXk67n5blWcbf/fHVVwNIWi4qk8uua1yuSw8pzdj5lEwb9hyinW
+1jGsL+QdOjVPoAMIjCGBsQ/dHz9XGSfwwhkXrp7o328jyXcS+l1qduCiekeRAsK
zL9PT3Em0TJpfLNFj/ymI0H03bb0sHA65Vk4og0t6gZQ3QDFfaM4LryziC5ccv59
hCQTucI+9LdxD9QGquWixE2+cRF3Yh21/6Bfl1jAJae27SZFjkwJuLONy6CD8SnH
Hs4Hh5uoQroUrWgzHmfOTxE90z2DVg316sGkNDgABVj1K04DhFfDRpGZ7CTtHp+D
epW2O/sXpIAbIFSIU2CINncJPavcf4lPJncOwj3EkQHwIPKIzW2BTt45QiTk+Qm8
OouKSOdHfjTZ0gFP9aW+F5nTyl15WLZalKkSDAOuuzG5feE6c9hn2B4WwiO/5jJe
KWJs0h/Fu1aILsHA+FW76P5/6NtIKk9eMBu+mrZJjfRhGOIPe1E0G/8Fo3yfhheo
HEaKa/M8RgSMHAG2kc3i0c9SMpb4vfULcZg3WEq0pMMCiLwV2kDroUzgJinx8siC
8VKosDzdGf80GVRTSfe3okvS2fzVdktv4Cr6RiA+FRm2plw2XuFS5y3ucOY6hsOb
Typnmasy+69Dutz078HZUnqI2DuP9Ipn42BuGdZPpso6UygKKuSC5bnRxNfRQW3K
hpEETqf2YA/bR+YHaphbfFBrXX0mzSGwSwWYcY4uxjsIEO87T1omLbmuFKS+MuIZ
kwGpiaPLQjZBLdbtELsbPrxMfH85b2Copq58TEK2s+c3EcFkrEIhSd/nUwpu9CP1
gfWih4sRcXtmxZB+dtZSLo3aGwUOMhtLtFszyeNdvamhK7ErdZCf32qR4gefxrfo
YQ3uK0DNtmxjNIyDr3hB0hXRVbG8+Iu+PYPD4r/9l+rXpw5UOUEPloTKbP8yqgWd
1OvNclma6KLL6wGZ6Jw8pLiL9CjZJ9b6XZ9riyZZqXahLnSV3ohJJG+jwOk9Kouo
ao3GXcJIcr8DxSxLqmMhq5Aj6L6q0pxwYjZ+JCQKKfy8gQrjo/aff3m5TSQLfiF/
aoXh+9aZFA0+joPNFZGooO27g74ycXbzsdY/H29mOixq2K+VRNF3a6FKNX9CgiWK
Y4OWEDFOk0bvfmBtm62/fahRtrF20+xezcE8v1SRJxYcd5zYiAtfP/nWyzax5zOx
t8R/4oUxv0CjvezRmpwNXbFr3Lo9xLUrkUNcbXIa13o3xT4kPEqdoJhks+sKKCgV
dBQ/5ayHvtg/RFaW7KzvhgN+mgUyTJGpV2DBJmIjiHdROGMytmV7XOUeW8rynfVp
TBUJArTlenJAykVg1+L3kro1DC7NCjQFscken8/3Ij49kOXZXM+tyDhdyy3DKJCM
b/0IdApbRj+csw1GvNWD7JQbRzAGsFAL7WqvCwRF4hn+iVWhrcgJOEAJAa5MS638
YypcU6jpd2vf3RvOGAUmNJgY4NcnQtifUtKkYVUqpFrT8pZi0AraIr0YZTKsXKoo
3tBQOn/SaXZvEf6Xy1T5PjiCs6eKdBIUSPFx3ZnGGEScYiv5vyK358K/oUE9NT1k
n7IdfAK/GMVeBVLTKPGJuTXiFECXIgn6i/L7fewnCONyLPUaXLJ4huN26JetzK1U
OZJ0tA5JBwaD+kx3y+VV5/ZppgF76Roz8qB4FJbq/+2G7HXtCACTB8DKDDq7a74y
OldXTEn7pRGcntLhV33GFCi1rIk7qIO1Bvpl6AkElqeGQuRNw5Fbw9ZHP3wgPwya
fJRU9mZmiqqpzvbzQAqzzmcLQK55vRRv89DF8lxqWDBo7gkXlxJKatD+LLYcoefM
coXEHBFCLjZ6YixQZYyO8U3r7OS+QeIHf/9G2ecYU8AVdE2OMBArrphcAfRMO4o6
mzHN6w8lIIyJN9tsesEgMqaUtHfXEmfPcE+wuvvhCtDgi5dsNBC57BE0AtXdzuZT
KiPuEiQ/0syc4IOI1FFL1JYpBTsilpMzrWrbYlbQIq9Z6HQl9A3rDCcH+WnczuwC
C1f0vSWSIQXrukVx8mF0rCP4WmW8klIP9qjKZq3WebmV1f5vsOqI6DqrwtUHA3/Z
/4VoGw0nEMrsCkFnKpGkiJJWHQjmoB8+osGjvo7w9zNLevAM4qFe2lHPeee3UtlB
Z9no2S+uKZXDggfb4v6tgI7azdCZqpOysoiXNk/LKLluNBwh3rAiiVOjlaAZZEqz
E2H/GDi1ZI1wXYNkEKoEnezdB7/0A7RHtsEp9Jqkwkzpe0vafGOscjoOkA7vZHde
GO5pRgwm6TBvCgqggSPwK1LZ5QvaYU6Uld2oZK07Al52RObabYtRXuxi+oyf8Joh
qRd88jthMETmSMRczYpsK0SfThwAj4RpjQn34219ulPHEBHdhBpKKQaAFXkdJ6yj
8T1xuhFxU+Qu9JhLYUMEo9bS+ctdxvYffcM9hpRLml6bxOf010hx8Jw5vy3Mghjh
OFJLHWJdSQEQkd+Tsbq0n4BpN+2shRK55cv0VSLbAiq18JG4awKD5pPwcTkf4KCs
H9PdQp7TW+OSahIP7MvWKDKrV6omyPkoEA7mMYlsSFm0CD4xNfkdcXQJ5TanEsIy
MuFdUUzCtCcz6Ks/dVQpYfOVLuEmqJuWh3UcfRe/+X7C8rDm1MOTcBYAegseCL99
28zjJlnwtQgSCD7s7snDuHOZbrBHPzGHFXml03Nf1IZC+6puPkNzZEJNDyUeDSFX
XdG8xaqFmadnGrbcSo24F+YvageC52xLbOCTj0LEranEIlxk16TotIobvyq75rwE
ePr8zfMCwrdTBtyhVU0xXxAOujmlw5Z5tjjsPaKfzhI3322Vb+2eu+3PiXvGWdGi
2nLrT/SxiZwwrDa8VVABWvbtyeWONf3zBsDdfoiuNtCz2Rd3RVqD28dDSZi+Fh9w
to+qcZtj54x6S+TVNSBJ/7HBu5pct/QQqR16bE01IaoFD7+a3QtdRuAEJxa13wIJ
Fzi2SV43FyQvGGLcqCLoS1Ixd5kxSPGJKBFVO+7/AtY+2fiKRa0j3+4prlza5w/B
1sRA1RHIXucrudY6x9PylmH5lbQkd9HJNcQIoiERbvOAyZ82so9gFU22fDEGIvw9
fGl5LWIs3q3J8Rh3KijPfiEKwPAWHeT6Ci/emD76syAcjUnl1MYoKy7EqFJtZy3T
tI5FDwU/jw7zvDjknS/fpFd4Wgea73xme1N4c9NhrLVroovbBYqWsRF2nUBrbrAK
EtM5XytkyjtagghqNFjCoFaeVrqw35qG+wuQFHKxPcA7pNhNy2DLfRYYOKNOfjyV
w0T0AssxhZ7kc4BOmHeLyO+6CK1TbPtiSAjw2TWPneNSpJ1tD0t7euEoRrASOEIh
P/RHipB4uPokuKHNHNFr9ghqkO2zqTVkhx0MNFtkEDvF+XqCeKCJ+Gxq3AhxEK1o
WsORKVoUKVxqwZXzviw2tnMJhVsO98IqtCa2MPejxw8pr77bL1YbHrfYwQM4rzHx
411163oywBv5O+AGep/JtSBpkFYEqgo4tx1gvy3HyByN8LeRRuBS7k8AjClqPzLt
Tvr8Hsl8O9C1N1MOQHvXmEJPuD1VwGIFeh31HM0e8OGEnTLrJQVfOfu/TuRIcakV
v9EXiT711dqDbg7imtHpL/VWgsb5rl96potZ+4oUSLYyC2dOz7cXTi2O7GcJIGJe
dqoUWMmAu72EhkPlFd16z+3lYgGVmqh7SrXyMQWZslOc3bwJk6g0opzkWCDZzrEP
/OsM+PmR75cZZ8YoYIheK8NiHKpHUvj1bC2hAA0VyHyndZ93kWCi7NhOA54b/ce2
5fAfpdFaHxtN0u0d+0hfPD00GD93neHzSpjNLidRv0mRKJLF/k5VuMXsyOd2LT/L
+osRaffVewFOzCjQWNKQCk7jMnlFJZzau6BDl6qEmBftLGe1e8NabbgTGTBvHQCs
0z4m7Zgr6I92TWGw9FaiMmVorzxOFNlZV7YfwkGTy0wyvuLXoiyn5rQ5ke65bEkP
AHFLEeCBNVYYkw2j/DCJq2TuN6H1UFEgI77/nCpDRQGAUNjMveFSRLf/uSDDqvgk
luf9Fb+/dWJnV7/KjyZIk3xjVa3cZUcCDctRHEbR22c/g+OUPNnMe7P8A99f2l/n
xZmbT4JJ44CefhByrv1xm7Hku/qkho/HGsEw3jxCPZzYmYk1bpXm/x0F0QcR1yM+
r7voM45d4HEub4HglYPoW0VYToBqfOBkH/kc6pR3EcjMTt4CMvA3WHfHEY1Kwom6
FGpnYBx5v8Aiyr6tQTzM3UoaTzKswnOtTO+9moWnxa1qu/KcPtKlAreohwM6GH+M
PyxScszDyEHZD3oQdiU1ACxbAbOTj4ZYLr2jVnMdYl04fiIhnh937t+Kz6cVIb53
Mt6Oc2b68tA9PjfpoAUptYR7kisgNbcktD2Njpxx2Ayj2lvXgRwZ8ifWj3YfEPPp
chr4FLDttYbAzACd6xTFL3Bfv+TPtrZ28ENWaPFJlHLNkaHPbNkK/ScED58ugdrX
5jj+zNdU2r1ZXxyHxsF2Ms2mGJgV0w5ICJ1JEbT8+FAiUnsVk4QdxQ9C4b8C9PXl
sHoEkp5a4VZz3YnPaY3eQDk9blXz/CgPbmVkAsjhZr89JBPdqHcAaQNfxfGEllGo
8ZmCdyVCJ/ebQgMJfHxf0cdMloeiPXV6MXrn4r72zZeNIVZEvJHDskTleVkzHnlS
QVv3BHKOJcHOpaD3rog9B33jDqYc1YCwEwv8lO9jicKICDwEkFaosmqo5X0BU7qt
azoBu7w+3FBMbUf38KZ9/WofIPtrn2xsTqXK7HE241JygvWYeqah17k3AQaB9Z1t
HVw+WAD4s0T7D3RXfyQ3zYAYDMpCuvLSZhOtAgUV/+BqEGvzkqcQhOSughgTs+rg
gq8lG3MMWCVaBshKr4m/WFwDaSSlstJIPVGp6aAI+nJVTaEJUm3DfiNr3dvbLjSJ
gcIK9e2ILnwiNxjC/TFfXedVW7qImjCHxfx8qFbyZknbxS2mDcPdL0xpxObPgTQV
aj0VjWMZWjYLh8gJ7MRQQv95KFIIplWp4i0sDg81eNAV8JgtOGKiqiv8eEp5kDK4
gb8tn+Q4SkmrLqkuXPrPy1o30zHCDU97E6fxp+RFi79NKX7CCN4BXSmljeVK8p8Y
SxhVUnDCztLf5JDRwCgkpMTKXKNQupuPBvT4j5ycRFvmHyWDNrmhaAxhwnZApZWC
GN2w8HVeNRtOCGMwtjPvyUuHAuGoZ8tHjVCctPLyolE+n0eyFiQgDVNl7CQJFznU
9FWOVxygHQ6iTclru6z6w2AHkR3BUN7Tjfp8/3WBsgmDYUKAg1afMyclBW+h0u/h
IJ+fazf8Q9xWNKAdBnaxv9oWjfevoc+XFfS8b8gTVVkjrnIcu91PX05c6TgHIjuF
TQtmp0r+nN6XvFgsM1Fld1ouRy0157PCYoil3MB+pbtuDSepHBTkIbgQigl0MQvU
amiFGDlBu1DBnJXIhxsMpZzwFHCQMfQVt/KGXJtdLWvwkzn18XiQhBOISt3+hw+x
DZCo30DDfoiMwOX0vGcnP/yskrzWfJtH/cdEg7fXGg8zhhCL32nKWX4vFGr+PA+u
jQIwnmI+oGP7AmlFN4Eqi24Z80o4Ew7wvWb+RRaduW5dTUy30dEiLsiPgN0SSddg
l03rUhj9rLLIwXLsMv8XH76bC5NZTnRkzWBUYjm+BacAnwUHI6DQqwwB0qG+HIFW
0dHeGd3NRj6LmbcBkp+l09e31fsrEOGeo4S/XkR6O1a1rB5UC9hjB1Hd5dLdRX4U
8V/Ftgzg70UT8zkdsvYwzKB8wBJQgSHET89Tw64d86rPHp/r6vWr5LLseaVlsJrQ
/xdySg2dK4lxB7AEZoaHrKP3s5Vji2HWt4AZXga+C03GKDLk/cPF2pX+XtXO4c4m
/68njCv5ujy08GrQH2bmUIinSITAaI14vXvSpHZ5jaMYYoeDzYyaimzjEfeSMLNn
jKDgG0bUiJcxdrw3XROuq0s9qMwA0T1Jqtknt3RJ9SHK78Cz7vuIGdhHJcr6K7zh
ioVdrbNtFk8rdov3zczqpqyoh7A88YMdLjzOHxumoZ+m9tkL3TzZzyENXrYIzXe7
npXctIXv1H+wFrHVCtZP5S3klaegnYniSgGL1Q8czVtrEge78T4Rs+0yZsKBhGsE
BeDrdqT23+sPOfXZLLorwel2myIegi/z+cg7iNAafmkhvSYQTcjZ6eeaNBCK7/67
8aIJGC4fQOgiXxNK5dm7wGfkbS9oRJbbVlzC49McVySNV2dhGmN5Vl60+hAN3+7q
3B/w50CEMHm1XZeHqhzOMQgHvuJfau7WnauNXOxyG6DuP3S1wVEiG0Hv482Zmui9
zLr/IyhjlsZVj8tc6xW0d4xT/vNAJuQgmDQfTgjuEGoiboBgOCfvj7nd/MNTl7JQ
whH/KkQAISvcUAoAjOQ6ZVqmImRwK144tcSCJMKgAG6PDIWmB2H0QJ4/YkASvEH1
94qGowoWYX5RG8oQFb6OZ+iOPVkI6TFTBCWbKmGFig8mvikEJaecWQWomL9EzbBw
l06Ugr4lMx/73JymvWeN5z5csm2l3k7zVKT5xPrd+8hTbXovG9BvgniwF6Qo0/62
Imr1VEwGBBEzSeNsYqeEyI2Hsl/5MEbgk/dd4/Qyyi9T/kk6SY9vbSMJs6TZUJ3I
7BdZPMEX97BnvYzufZaRlqeMtcZplRyrCWhOfcVbB4UVhic0SLhnRKpSBM3XRYd+
0XIP4qzEHA8eqJGOfh3hPtnt46iEmfrRkiiqBb/BOedYXleNt0kHNshVd/7712dl
EkPdOpug1vVjeAd/PZK7EBgjPd7/zoAIlWzFKCCKbij56/2RXOnGFj3HJACt0Vs/
6gmajl1WWu7m8+Udfi84rDfAXByPZ44tTXS6vsyjseij94SJZqJfQwRKCuJRO6ek
3umZW7xNMuheqf20XgPcE9BkVMGtjS7j37L8T6IqKOgaERI7uCMeufvxbQEATYye
OaCETx1EkxJJ6lJJbOWe5bnQE9o2WrtNSGT/o/oRG+SJDlrIhJ3SOUXMpDj4mjUH
CMm0mwgWoE7TIDgd243MHbL1GlRefzCNyl0j6kSyLw05SyALWDd+6TtC0/d7iL7L
MX9j35EKHOaEr4vHoJgWJZdcq09Sd81diKGi1LlCGJvJA1XbDTx1JLe0+uzNgELz
+4tZenK9s05TbQJGMDfO3ocfTAKepHZ8+3/Eztdi2b30ru0rW/s98TnO1mPvd59f
19IVWznk8bSiiTsR6e0n4e5id/bzOO5RSm25FJ6tYKoH2Q0UVq/TIJ/ii1RtTE+j
3bPN1Hvxs+7xJipVwlBce7r5aN3ZTaIejBA14TWqP3ayzJuQIvwips/DqiWViTAl
OrmPReCphNhUqRqk6HeTlnHtuGBWGClO/1WYRS6JdYKOV4S9Jz+yi3UiYNbhelaw
DjgpkhoiTPLA3dnbpqH9IDy8+1NmoKjvjKkNESEdUOCppGe2T4vFv3yUyGlHVHB3
F+1QE3qJkMKxZmPEX2W08ILEu44gIQIWokY81je/0dFb4SIfcoI0lHfooCOz45Xt
dn/XNIUnBlSQ/uV7K9UcSqSl0C032d2EUftPtRqMsLwhAimD8L1+zkQPgFqSCkiZ
tOIjmsvCWlOztKGGXk2ZgZFZBL48xeN6MU1pPbghniDZFpf01TGu7L8hLOjujqg7
EAH1Bh2BBzaQhu+SDtHfNAl2qPxoHA+57REGUl/7sO/AwyTCcj+lYk4Uv4CWZs45
9RNwFLROdnr99csuSvkP5FfFyCIgl1g6vhQY/yCAKy14a6vcEgOe9BZ77W/s2wlU
NQdDjeXzJE5CVonvjny51hfK0sgXfkE2kXs2PHx/jaNYRe2dVPtqKDPq3Kw37EjU
CPrJDSfKu6EN5xugimwhhupPsiJ/5WZJhosIqJXqvKhh6Z2HsHK4h6wGd7/4IiB1
WCkVEAOVc9gZ0Gjz6YD9B2jD9NYYnij7dRJeaETEJ2capKy/yevjH0FU0IeKU4n7
CAo/uawDrYc3DX0WgnQJJ5KT69rXCDN+rG3tAfrFcstuT3wEPs+d6TqPwISGrJdl
qqFTB5i/RwhrjqykMbL3uXIHCilOhuWpYotFatRkQ3zT2ICeckhsqYwQe6sT0bGg
YCsQi7fnjINGYDNgRysICs9zK1EQ2rfXsplrfwBR75n4nClZFUylbb8+G1b1bAjC
2HiVX5KvYbp3n91GbeVez+PWtnrEqzO/1jriKT82uR+cm4XCYKD9obw1ZlwplSZb
TnAtBz3jGpztlPsyQerrNFFsHV6KXK7Xw46XmQPgDoI3XT2IeAs+3zQpRVmNL3EJ
JBCLsIOYKW+UyBO81Lvn5fLUDd9Wtn/+U9PsUHTPmZodmXdlkOc+A6c6VTBxbpbo
kVGSawq/1k5bULjrlrewJmTQEkds+QNXiOzUjZR2pTWKMJMPvH3Za+xpnQ7o+L5x
9brEeAEcdd3wz1RF5p+RGDbgFFyMwKRW5QCggiMO/QxIQSPXGl3SVBRa2BRsnPxz
zbunmR0ELGVp3lp4PtHzojumuBFW6oGsgDo8+3ScJlfZsfQay2AYZAnvTw7WxcLY
To9D3pXb90R8KiwllBa1woKCQd9tJTVhi83yf/dl5PihmgPJrDpuQatbppnNB/os
B3HuFxGEBOdzEGj0POAptO3tMeZTtM/LmtU3nNDf76Bz/adYUzyeBaVyCknDofzM
hE3tN1/jEm9oprpD+AUskHHwC0f7F8DiXLDxCkB78b1gzQ1cjlnS2shmfMwXevXb
X0PEzHFqOAEiPDuPuj6twxx/5XXDR94B8YJH8FmO4VNFt5sG8/8ZlAsg5YPFNVTn
oUA0tVha1+uFR8q0Cp8PFnnYmXibpepxhk3umnSVdi8mKu85m1g5H6ZcJLdSerIU
7uG4L8JC7bmbxn0sK0dSxfdfGlP6d9J4vz+oKp0+h6OxiraDrjg2Xi13rU34A2K4
YvlY+eq1jfYK506LVQ/BbnE7hncTeHzTY8H0co/CYLOFFvFHkGao8D69guKwXCy7
N7NrlTE/4/O8ArnEigjnh1e0Pz/GsxFFQkl74nYToqLy74qtgZrtnePxmn5O92IP
ClKlDUuQa7OSMWwlWYA7VfYtgwrKadSiNu7k9453jNpv4pGFp7T5pfKYOLWijgFQ
BwQy5mYgqQm3ebyyVkarWZMu26Isb5o6NWU55813TBTO2xOiR/+x6KgjsQGNyhd4
ZEHgoer4IsQZK53HuLuKI8R13NCkuFM/7NvhGXCvamsKH0M1vHkbJzSpcaat7age
VTyzRZQQqFV7JeVm8JvliMUcVrjaSlxZ3tg9NGjM7EBEa3cg3ibklI43bWsYP1+m
gnW7v7E8ZgBwIK+TlAt2kEhEn5f4eY9Hab2NgLM6YFOENjI8EYb7lD0aF2hYdUEP
G85HzFoVOOujUJgP3s1u7UGrU7vBCfMAlzBWDESbgT6rl1qApw4OstG1r3Ummry0
6kZKId+eA0uTjV8tzgaiKLWarFI4zbWqkicsL3wa2sPR1KKmDlq1YuRV13WC9eHM
G1x8A1HRia7XV4/37eSksPd1lHIkRCINSeifFBMHIwrGanA8bPnBNIokmyuoYG+S
ASkTU5pERiHNb0IrPlOpvLqsnifbBzeIP9q8sYvlRd89jCdIFdHriZrIljI07Ktm
lnZO4ZFybegrd6cJCnf1FhjD1s6Q0JQxv7n+mVD/hgNnl1ZaOpJRILwfyIXSuQOL
9tX3bQw4FabVan/X3BdxQ9SZQQJGXzKEziH3haB6RVUhn3oO1uR+xdTUAauFB1rZ
LfwwYebFLtZQMU7AMEe2O+VnB33hBnmK3D0mbOgUOcfzbxFUhpj4gTWjvQETHBed
8ySP6qQ4r62mULw232cySRcM5JCbxoPxucV//3VL4Gr0noXURPDlxPjVbXI50OR2
WxtlPBMD0O+h+MxeHLPGZX1dwpczgbwT4nWM8XmP9c7aMr/I/R89Qb8qrkUZjJ38
ONM/OiG/07gMQqGk8m8QNmdV0lkqus8kjn4iuvj+dCHsY8u1EZXGGrByDAcq0ckw
rXO0gFRJT5hW2iIfTMj0RlahI+nCjm217QMDv8a2MFzu4rfmw9LSxelwIpOh/I2n
v3l/H0IprKU5NulU9uCakux4z7fos6ruuGiSpD3digjdaib6jlv7n9B9r/yrl7cY
8kT+j36GuhP24SWy5vAl1I/QizK6bazQrHf3P/69hJfVvn55OtMZprQRKJNPa62X
tPjWM/ggYiD3VqB6ZVaS6t6yHFXeW0WkTqKwIR5U6k5SmhagXgjhOFM4IJUsW1nF
qswmgxlUvFmff/AiAL0ejd0yhp7/O0anr+FIK7MVO3z6iUdTQ4kmoYE9Ay/vMhDM
m44OPtZWxuP5tCQGRW3U5+epLL/cZJNExwzPHy09lWfMKawYv0Lor7CQlqzRZqIt
16yQknYPRh78AJ5i7IfXzRd+2MIyfswDCnIGcOE0jvfJxITYGNAFMJX3HaNTKszd
ls/UgJ57ywaRJbkL7hnGOOkBTi+f/LRJbMb7FgACLC3hqavFkx5AzIITF0KyAsuE
xAZo62X4XqIDy4m1iOH9ZMR6+x8FSEkNZVaUySuz0uSVTXhHhZB1Xi/txCDw2a23
e51Si9YRfoIZHpuDePkOS3/HlTZ44IC3a5M3l21R+EaiOqN2tk0GNWufMVpY1pia
NHdQKAoFeNUmnNejv93TAsECumNbxYjYM7UUQNepcLUHOd43ZYm4JeG6eWil208i
gaPHCsugd6gVPyTQ0/qeqMCNylbMNNEiE8LFxXRwmd8A3H1qoTAUiIPvNdjjyffU
Ua3h7Y/aEgh/oo+Zj6/zcNtoHsPka8LX1ZfSBGXFspW2UNgHr9Q0ybbMNUrVxRpI
DQplYP0DsA3Om9tLyMT3thRZg1FMMaNpegGbiPHMStVy1/PobYhXj9v91b7LxydP
o4LHXRyUUqzCUihpJjjU5X+fzYWMnFxDVknV3uCz0OxN2NkqOrcj08Y4n07qM7pj
GCoU9d2UwhWIDJ2UEZImtdZkQ32P2yziWE70k9nMfi0iqQomHW77o9e2z2uANbbT
lBIc85AkgXWHerUwtfDYYjvfmI/V769bTtnWKrjKLNLvLd46JZzcMa9m2cyl4ubm
uj0Vw0fvYm2bXTBEIPXE5GiKkP4p4xSs+94Aghtwd3jbELwxJ/VuXEZVOPtQbBWg
WWT9Rap9ZPwHB2RaJpqPnnO85myGkGxUOOnHAu1LZ4UxFDFsqfenSOLNYpU6WV1x
WR441lVxoyAEDX4ZhHQxvzzjNUwqvJVR9PWLiOlKu68fKNYJ0/FzG6P7WwuS0and
W+fRBaeuRDPaqipe2lr1kthJJ0cNZQf33ZddlPt5K8C3tijzGFVCJLijKM2zImtx
m8wc6flUYI27tVQMqQGKtsRnmgSXx2KzlSZ5gL2nF6P/noIHsleFT+F2csC0DnBY
hPHvxP7nytzoFk1+bsdkM8r+El80c47Qg7QcuNmzm5QYtfA7KyRRtVgNu7O7uFVF
C6wlVaeECt9/075YqI2MZAyu7MYHRS2cHHWbYI6HSeQuDey/CeNlCH2oF7NlTI6d
Tt/yJgglL4yiyOmXXw5cXRfs7AQN/+0YweM1wxODLjlKczXevzQLhSkidRE+8Ia9
jTgrWvNwv+Ikl0K0mC8xrV/mcSTE6SkIOxUxj467fBSGXXVJogSfdzOvsCRzI3Y3
srKA+luUhcs1MuUSoIRr3lFxhZrw7/fkCcLEq8uacs9tqgCIS7FR7ZeLaeRdlKYJ
x4uJc8qqlm8y50hXq+jqiXhCoQoerOfVls2hFal9OgCeNgwzU7P1ZlQjKVQHnthe
swBirwpqFJVUyYJIBivyZVL+jHiZKTzC4TD4uCvFgNUvS0iRRX4oEt4HGtbECMeo
mXUPUOn2lOh6FsnSX9EQBXcvrCxTDFYGZTpMfxXx47yzgi61JV464ehwF5OW5yGm
q5dgfzFTMEeqOjC1BKeaj5mRw/sGmahVaDcv4Rxh9CaZnFzMC+3MMQtRzR55pVp3
YUBuuHrhQt684b4bjP3NeSgiOu5DNv4p6OSzgp1Pwpwe39raSK8bq7BA1uIVt8HW
bPXoVQ+mF8PU+Bfc4tARnuY4OE92757jRKpCOqDPAiMTQ+KWTTpr7FGtgeKd4h2/
GA3rcjkxbiqCtLq3rF8Z7obq087V/uDV0ZelBvC/6VNMAv2CY3BCpdBqJJJ0fvfZ
3/MWoOTCZW/pXtk52AnVGqw/TAjY6vdVfkFjJiENVkcHA4/PuCSC6lMLEWNsiBg9
N1WjhS0ZWU0IOGQgvodO2nxNYZ27LLKqL30YI7KA5Ov+hTlw7A3z8la6gEriiyP9
DGynpS/9X7B1LZClqYAq0XR65XmULhf++f6kicqbsEXq4d4q1l9JPftXxekVrr3T
k1Pnt0x45z9pbKuwHFsncZIKZ9blk0vrzpoRtnXD4Mi9Ts7JSwwoGYjg+xh9+hCP
rvGMvtlIxYfZj1ySjgeul4zqdFeZsQa3vvQiesBWIQSJ+291/7nsLI/PZmVqHRy7
jLiFT+Z733ZI689fyHrpXG08jK2bUXMjDchq5+mu1FqUUZ7ZNC8gOIdi0spqNeUq
s5ic8SxbxGeIOKuqiYZHi6upjAI37rb6Uco29xXK9prmywie+tpxiG4ZT69exUwq
eoRjCUUibG2YATVHuhKFEG9NGOHBAIOXl18rbYeBs7cSOMQL19BiDb8VLgO8TIYw
lRDeFVguE5nSg8hb6k6aiB1xCxJyCdFiXgcYehc8Ds292fTs51qVPtYzY/HlETX+
AM0y1VPPdf0APoHc3cO87zKKW9BCGgbONMN2CaEvHcyJqlG36TpnUHNNPgWtJjoJ
rDkSvPH3GV19t5bsklq6ZxSDt0PUa8bMrh4qmZfh9ei7tONOMyfmGijsNiU+jjfn
LpDy7bogeP7tcBvupH7EnW/QW3UZeUdfMNjH42N6WcIWz3DXfIDjibIZHgV2L8OE
XrUKtN6TcuTKwCEm+064amBsuKPLUwcQTxjeH/ZvWZNCM6qFaoXytil3/DtrcN2c
RaRYn9f+ztxHb5Bkp2rae0ghe4vG/H7XVXfsUnRXuCONUBmCVbaoT1KdbndwCQgK
gz/DoYywQ39mt17U6+tVmHrD4+/Q89+RObC2/vxcW3yS9FZ1oW0msqdiOzLnP2fg
sXv+bGtj74AQhqgDNKuyJjA/sAybjcO6l8o3k1w+kbGrO5WU8G/fbek7EMqLKKhK
WYlGoEd+WUzRhIV/3LGdZd2FsVM8HQvMCdfCv1EyCPNRIX9rrGgj7zhnLk85E0sL
y8mShmNIa4IvrbahBhLDACvAEqc0tGWmY0qVh+k6BJZa4M7yxpeZGEoaVTrgvXCU
/n1UKaY8D7vKI+lrFAIYutNDHlinOlucxVRC9Msp10yokGXVn5Mh8bYmOwvtY0dd
CCMnLahJSwtbY/yEXr5Ros6dwIeSrAsfSdzWgjR6eiE4UjeSBuFVzsVNYZ+6As+a
+BnMr2SEETHBilRuCTr7K46kWt3uDILWTl+rd+uMfmTeummxE5d954cIk1tqNsaO
2o+xhh0/LXfCV3y+QmILpQzONmHwv8Rr08SrSMkqe1qrH/UfdFReWeR2d4L/PWwh
dToMQ//5bkrNOkizDXkrSH5E6CXavkKJSlXCFXmUctATeWr1k/MLDSvXNHymafFU
oibyfhlO0rejpuLc4eSTKmcIiuJEfdIZPrKTGvYM+yDzKQowcGxILB+LQzk/ucb4
8BxzOAt+xDY7B8VQ5gQf1MPYuVfsLZzkWeKBM1HnA6vWqEr8pptp0HZuuTyhehyI
QLsJKVG2VXU9g8Gdwi9abEcKxX5TbrPv7dv9iE2Zt7YuZYxQVpJK+c4fKneqDvdW
s8QXdpBaQkNb56cS/nLT9GjkI7E2DlU/SzvsU1VvrjS0Gw2f5YM2Ft6wXYUhkqZ4
tLSFLQklRGrAOhZufjagNYs6CavTtM2QAcIR0b6+RusBuAMiHNR+vDFgRjQSnv2M
+PpIVROYcvkhf1ZWQACkXRPlolVmdkZubFsXphbhprtlQesBaKTcuI5KX8DuXZY1
HKEVtyfLKINSlmccKM04lYpfPQsVW7zDfoeNFazB5ctRJMvx+3PjWThdEKWPxjr9
qBdBQ94/yadKwnp+zoo7U29AJ46OohkFZqI2RbutvVPzAhI5590GEbcqgQ8Wi+7A
LjU+nroNjtzFzM1w6zxUBWqEXG+ZBowvwU0tMD2T7yxuF0hDq4msCvaRcj1C6E8h
CDvV+1fsVuEgr6Hl93AqC2VwvEPNC+wHzEczuM0EdccNy7C6VdyqCKkki4nQ6O6v
RgD1zPItrs+VFb9Ltt69ysf+H1+WlWbuTMJ4/rctng9sRfWTxmahlT1JL3311d1k
q4OfVTrm21z9Cy+x0uXKthPCpI5EyApJXQOu+VW49HJPd62OAg+3jehLGs4+SnE9
78bqu3JqrNVV7CWr72oY/nzdk9C9B961scKJLveOs7QiVUiLPpZ8OB1A63xGr1Y2
ZFc5dPKBUaFjD4NRlM76FhbelKdzcxeosCMpXQarPNwAJYbaDgKnudIJwsRodR5I
mlsvdwiSpNuK9uItcyqWVDYSI+veC+/irRWbrCb5FoyrJ2nRZKLlNqu+Ii1UmqFL
JgZCnYVOHGa+kNSqW++nADkJJHl02qLoq7rHxNWcs4AxfTrZr5FUhLdpG1X2HtQw
/PN93s44sgBc6W5DptUfJZAl8Y9mAmDUg6Edm8n6DQ7T/7+UqlLsVjJz9O+ls23p
K1fRYxqlP2tmJ/0UEV7Xhw66El5SFYE/zzfbLNA+eLji/giGn5f8D2Dl0eV+apQ4
7oD7I7U8NdBcHEWPdrG+wtGoVX+cxlMgqvHqdAE2m6vvK/jbZSNlMXXReuDgGAJK
E48f6MzfE81cAVIBkYKtNN1pwBdFfV+k07s1BPaItSJgAUllR8EtcyFr8r/9ZmgM
wWMfgqdUvIEQs899r5O5oLlhQBUdEKsyy5OeLNwC40FqLkdipQwcp0Lwpm7Bg2u2
wE2EE4n0licT23eHYosLwPTBJGCmp3hoF0J1MBjXhJOAjZYryb9bATQnTtf2uMcS
P76hu1m8tdh8SZbDHvwJ6w7Shoo+I5hxc/4E/173OuMe+TUqfl63wXxy9uEZ3vxG
lSmBSLBtJv54m65OPhigbd8lxe01GXUkNpPBFNzqynNU5CFeqpLXOGiPGYxRNM12
EXgyhanXOSKrb4UxHkzF/8PHNlqtftcLWAn0QfGN7Jv6JvM/PeOR4NCRZpflYXdY
V/ys4sIG7832+Y9b6PWoZC8EX78BDXfedpoM8BwMtnB/fiiJtvyVXO34fDzC/5IT
9tJ8RPADMeyXMXyq3rlezcFP6pymMPwl/Zq1i8zCgRAaKxOX9FpSaeXnfv0v5FCo
a/geTgYh8L95Kvz3JPK5cWSVTJvUXoV46prHFthZ620rMjoDlTz7cuUM99jAsg8c
gb+6K/ycZCdpuTU1AxNUzLa0QGOrceIrG68iRuWt7mr9UOETiewBZTRlb2+H/jcC
vUPCq+1NpeK9uT3oZf3SnHmkcyE6Vm1jtDDpvy7UqxNdm858fG9mw7jLEHPEyIow
Z1VITOr8q2nUUbMLJQk1TAEz/35Ea586U3jtjstg1rIYqujDQiWr0bXvc4vVITFT
d3w+lsj3hpK9meiY/BzuIEvni2LBEpdS51HTaUsjBM25f/UUEvF5lsV9q831+0uZ
vxgu0Prc8Uy4GaypnzL550W9OaxuuihqwC82cs1g6yQd6mOa4dn/bcSlnMfGE5+V
JWADmMostfVhXz3OVISCT+0ZpsDz+9Gynlvd22CWDjRt5XybAT6emfROWVF7zEFy
98gYogfoo1dp5IMPbjFVTAUttUK6UL2TzEYz+NG4NkgQ8AXTRJD9trYdIApsX/9G
EEdUF4jfjXx5+Rs2TGXedhfAqHM6OtCwq/Jp9zwxO2NAGQMycTJHSIkoF1GZvCiQ
ZpLgOMV5V3z62tRP3Sz5pC4SPYNHr2jlghNt96sm090O4LjBCVhtaBH87j41l/P/
AQZ9fuuwQLJIRB7gk6+5paa61xzuR/xJKCu58focLrGaOLDEgL281Xd5hVq1qmtN
Qq+EVnrH77cx+2ShA59feZFIjUe1YCDEP+v8gdnNrrm8VRyBoqrcgErcOm+a64XT
dPIXkA3qkYhNf32mn7KAx7SVzjqCapv4kwaaF1de4t28hxpR0YOTnOnB5VLJ91kG
olzHKNV36jgcP23nmo5OKCun4LBhXJilJtMH6ZT1BmJKLau2esUvAZENoISHc4aK
iwJN4CJCEKjnf3dJ7YpWngP/6XEpGCe2aDhoQnEMzbGzmbojcya/uGGlgjtep/R8
Eq+vqBupF6D/zJJ0GzlAn5nTXoWOCfUY0Fis8RKJIsMNsHZcHPVK6qKvswzvXIi/
QhLziu1IqSpjdKWy5lV2QfqZiNnlWD0zpKUGLL0bvyUtLamgOk20ck6YtqAYF1to
TFtUnshpVNkON/6Ellba7i3MoS13TaVrcnCwwAr3qp5w62CDq65NChWNmoc+ACsW
a6calcUY41IVFebthnt1Eyx+d9XVtzosGNTzGxIrs1N0/DmOw1V66z7LI/Eb+Gfz
vTDNOb0tmyiIfEm9a5Uyof43eWkkE00TscUWImD+WVAM1OkvidoGk1/usv58sAdr
GtsjUn55S2Ypa/Tv/rnqCzRRT3dq+fsxJmx5FiEqCu31FuH6fLdIWP6fK+uiHFIz
kwlkBAIMbMbgHOKa14W+QGMs8WII4AmC36YCJoCtRZ7JvlObWUg7qOva+jm62iiX
mI/mLAVQn6ICb+hb9MbbB6odlUlTgqYWPVufjg7OIL+g9xEMWepbdxzexfUeqFta
CU3Xlk+bk0PT8JYOTMRyVuYMJpaLbScNBLUVJ1UX8WXTKfV4aXyAq0UblxbO8ifD
xmMBl8ZrLcy+A5uwumBYoI8H8fDNmJEBIWUAFud42JqTbBFqCVMs5bl9jzkOtNgL
N23l67OYzvdP6Y6sOH0hFo6mLBZXpfzRbL2YkALHGkBPYJk/qESXhusHCtqRYq0Z
gh4HV6lur8gH8oWTy71M/9Pjju4fa/MBnmsoaqF6LxNKzC3vPtX1KS6ZI+p/EK2O
mHYaH11eyGfPqzEqlPouUTOfir9BywqFtVVdeeVKtjdlUSeXS3mbRgR7qkuBKvla
4I9vRNsJg8x3FsPsULNqY6vWFTMyWA/XqqAIQpICXJpbxFZMkv388W2DrHspzS20
C+bAsZJUjj4+FlEWFMtCslDYLe0EGDenFV4e1/im1YvkJUX9TdBrqKZVUf3w8/Jg
iOiyWaaefzowp5IqWz9T9z98i5FwbkxkGqFd1pALgnFN5Tn27dvBlukwlGcC2mpY
zO8+q8M425YgglaLXHkue2PAogtwPv56rIZuSA+q9np2CWuoOTDEZ9JxhddhLOOx
sUMb/KcgxsPOLNqGkHAcBXNFRKhO3zBhiKUQVQAYfaFAZmbFUDYq2J1T70u1hGAE
dYenIDDl5JX7iVMHcRvnYuAH5fmOGyTe33tnDjhSwBXwCCd4POqVzbXEFwFEpfCp
ZYvPkrseCZmJPfGUMXtX0VSIVzGApyrithZwhv+iA72T/oILhuFjAnl+YIVlGhs5
1QLpVOusNR2QoRmhU2KEYS1QXx/OdDzkuooamdnNg2ugT53BjZvlTNeOTw7Ibyb0
tUHAuuWSpcwjzXx/wmyk2AhdhS5uVyhNxbW3daaZhdvms3QhY5HcUAUvDWGV7nze
dAXusOQqaIwBwFG+rvt+RwlcYmHHkPaTQj4sOL1hYxfOWLH9ccj4iBTokaIoz/WZ
QN2bxFnyeaNgDkUUJAUCfrw0wRw5xNUVTlOm2uPkD8ErWRf8SLsHso85jznQnl4t
1xwQxe8Z5EUBVVcbE6nfzUw9unoOC6SClv8LtG1tK+mFS0DYJ7uY1NsjZJqoW9yu
J2WJQSzp55V3Vk5zhvdZDuicG15yVRSxeTLhvqp83tjD4cuUzSxWrgqQLk6onGAk
5hbD/el8qPU63XYmGmOy1ELNgHutuUvv6fVCtPFdzE2bQneFgcCe//lHcFi9Lshq
boBOfsAhro37NZEncqus4IY5/8u9FW1BFWd6UYX0Mig3rH9KX0IUQt5SlaqB4lI1
IV5TivcODaEhtyOy/8B9z4BslzXEXbxCnOi+XQ/3OlWOPiPsHkCY0hBB/66bucLU
qg9Rc0rS/UuQcylGQ/H4MbhrHqarRnMD4t753WgkWudm3FVetQcqtq2zWxl6vOKp
scRe8CQ+j7cLtM3MGJUR5bBMgEDzGuyruubj90oWofPbSveb5G0uJSYC/b3VQXWG
odZybSNHB6njamXO9PtC2Y9AX1rEaLt2/CT9vimcCusbzJ5W5vJfJpfYCw9/Sv8g
sQ6e6aMKppbf0x5MeknThZ7Ny8YfHIYXVsEd2ZqeU0OtPRKx6jJEQjmhTIelR/YJ
tHZxNL6JF9byA3imjXUv1yK892SItVmNKENs9GfzAI/uu3+A+F6tNyMzNCCMl+Dy
e9voC9sDC9Ymxn5S3MWR8nP1Gow9yMlI1VgEnHcIaN6qGSh6zKxCqftxded3W9O1
dIufzWrIo3KjNdf1lMBgvGGNhF3BSDb/+XVWYoOJaaL0qHJK/pve/G6u4iqoGY5+
W3ETdAcpm3Z8eDAoWjWIVNbCsqFIoNJ2QgaczP+rGrFxqL3ftY7ANPrOEEC3lQzy
tpPYthYpDDhBihTa92HUgH0Qps/fI+SkMs5fOJIevn1eJZ9hxwIQBvBRERlCVjxs
o4p7CbTwtDXpJvDXYqovN9/OIYEBepeZeA8s4iOGGR6oNRWZ/knv6Y0R14aZrykB
ml7Cu2duRDVSDjJbBVhn0fltBGtg9/AfEjIn3gkqIChtAMGL9a/vMnwhUJ/PwoPD
RMZwYmlbruD2L2La/UplTHFDdJopDxywIjJmHC1Uf3JqVDK9q5qFTAvPSL4MTh5O
uSRbo4gcaHfcocciPT0FdKwLyvkL6mgLncDL4MCKlorovtTwNDSKBbW2ilXLkvnR
nwzexBrgdcCeESOqOX3ZN6DFDB4e8I9w2kRMn/QcTb9RuyMSFjB4BrrpiqykC3aP
q6Q8IHUSpjbLqdT3flnFQvI1m3GSTHWbWtEdia5Rn6X36jSHYQwMKW1HhZvMZPgO
Zqa4zkRQK2i7sILfgaK+80DH4ne0dCt4k+X4p8GewFXcos6FPvYLIh5YQ14gnLfK
LY2td6N7wWg9PNsVYWRlJZeI08znRm5HvQ7k7NfexE0j3oAgEpOcFEVHerm+7GHJ
UeYCLfZQPBe4wVYtCn61N3ePmBiRmFhr4FJrn5nFE/jrWICDnnrCxW2Gepj9DL3f
F2dGM6JVz2ISuZah60OEMu8GnF2AUC58T/pdMvc7WVVFKU34hz42htupk4yz+IH9
klO1OJ5MretFoQt1HNcBWp63fIeaF8mmehLpiDOr8Lk7Q4IcJnLWfVKc37wqCFET
X0m7rCWFcd/mfDrLF6TV+OWmLYsVsal6PuXQTqEWvKZ47qfaEjwq7nt05oIw/X2s
oLpdY3OgefLpGNMfvfBfit+BL+Els/crij6RdE2WndBYPgLSQSDQmoMB8e980C5x
vBcw3eIwa/morrLmadafFvL9bniLqMifFUH5uhm2SOpi6L9Ov3xBWcDhjVeAmxoo
6VXDH6Yf4Xo5bxZ8dS0wtMdKImAwFmYf3bltuDzK5YQHWBafm4hW8mtqTzxhVxCI
j4aV/QRcAxcA4NHBWrJZ5EqTNvDGcEa1ZAsEYBDA2bSeGin1hSA+KBzc4GUC5Hhq
kLwetG2kRchy8Cy7oIwKSK9R1wpdRdMSEO6PoCSf8vfJ30aK0+0H3/Byjd9ziKUf
Gt7hXXediU8oaIWnGT/3gs/XgezHQsIJ6hKKMhZY+zeG6ZvczF1mPLvXh9HNivVR
NwgrbNNpalR7UJjkqTwaRVzOiNq69OSaBRdBaF16TINtfiDQs73TvaqNWxMYJqA1
ovaSYqhpKEct6efvzbBJWpm8tGOISpvxFQcmF8IPRgBvxydSfJHci0betRzG7+PY
3dCxf4lswvKwut2HBcoo44xpGaNr44AjsP7BKEo7pzwx47wnHiP80gqiyGjXKKPG
GqfDTuC0uOI0t6rl5VR239ZyXXDKW5ZcT3CwzUajA/0DqRrF0vhuCdguAdUluRAZ
7h+VxJ+OTmPBVFQHxymDStU3LJbCxY2wub8Qh2ba0c9CC1laHY1r6jndBxgNyd7B
Dm/3a27RPvXCvmN987lx6HXrsCiPWB37LPUjod0zYr3QORnLdQfbomZnp+d5yP4+
hMxJ02OuBgT7nH8n5GhU0UvGdRT0qT9M6czdhlm8Pu+O20cdqBsjXmeQVRujIDgR
+rzVZU4tUkYTNdqG12k4+6mgaZpi8OOu78/ZcP0mJClI1IpkhefbRrAGqp17Wgpo
MYWW+CnxTdlR+aZvjoQ0ptgr6/f87Sixx6iRPSTsjgMLR/UYIkxqcsN2tCPMIFS4
Dq7BSi+CftOvFGyqDe8sC30+ELJz5rLLc9Pam7tQ36Z17oX6K4AmFM10GuPrI2Pm
8dnD4NZkkY7gMxvMmEHC9dnIBPDurg15dNpqm51lz/cMDoUPpHeDHqcrKVrb2oRi
6JGHWgNb3DMBpsowNBnx3zkLG4ShQByxNFYnKH35e9tNDtuobzu5KdA+bcdB+5zS
YjvNaG+/nmKxm0ekC7iWXbAqlHtDkDYLg/GkiH3YKHICqeBIQ81XTUXqpSY6aZvZ
IzZ3+/eGcxYtOY2qyArwwo2hWecUJjP/dCVEgGrmqYdJCO0NeDFCrF1vfWAyZLZw
+YRyvVEhlpUDi7PbdmR0pbLsGiEUH0x8AkUWcgONwMulVSI9kAtspzZi6lsKTP6a
R0KWqIKeOYsl7eEowoiXdb21XdKpur8x55+mHilkMnUK5mUmhcJnO345vOdr4ki4
Wc9RwaihmNtBt0puv8DdIgu7wtTtZtt56XELRzOMKFZFTCpHudrvBmP7tpkka0sY
9AAHHLIJ/J5CVWKrF7lcs0GUcbfdB9NNX2KQ/Nr4yvm0yNZOXhdTHIfYa8oXgDXy
q7SWDoSMIeNFg09FQfLvpbojDhp2QHedy+Xg8cKjB8h6U1267dEcnIIHSmAen1EW
Ru6wc7g2KTMLQRR2LljgXaKzmoxDFH907qiIlEv0sRMhBhlhg4+BRmpOWVaoz7pd
JZ5EMA+wMY5uJ31tDHng9u+Anri6bsEP1b0C23YdGTznDvVFY0JZxeuw5nYTZjMI
80or18pXRZP1/eENBVw3Y7wodCp4fD/tn54hbE4GJ1snpVBwKSZRofeWeUClUg7Q
2vm58SEXf1kcuZy0pv3buqwywaAGgr45h3Q92XYAY7STTjZ+IGhA+4KkXJSy2xjW
SIdDw08aIIXnQBGdgE5L7dxuHCAP2byO6OutokysM6r1Uslz2zZQGVHW2snU8JDj
W512luf6uL/sg2EaoYherPVSE6G02K50VyP1TCTGolGK6MNVC7obQEU8KBkCtsdZ
KA2WcDYgpPYDC2a22nasFUj1tkqaoZEZKLjeUvXVKJqQTQ5RPd/S7ojUqyT0veOa
Ypv0osXl5aJnIpnmG5OAF66mcJAHygDscsa+322/5mV2ENEEWCkU3eTG/QPfxJuP
XCVCojmihSo48/M1ka9lEYry4+o+MSbl4tZ5xQDpvkCekEZr+HrotHjOO7O8h8op
/qq8ffejML6wigJ6787swDV0s7obwCL6qm7NlJzLA91pkN8uKhwhcMLg38KyWa1P
03ITOLSJT292DREGnkOlwHUaHCn8KX5G3V8jeapx14QbBA1dtjvW2hUnzBpSn0nw
+HIhIq9khdBEvs1lxxhG/Q1bolDrBhEoG6iSNQ9CprHfiW7lDtvWOnGtz0tarlfh
qTOP4FM2MqCEG0C2YlmWlfIH0yaEDLezoHCLb2oN41HZNn7bYWEPxAGbP4IxHIUt
Od26vJeKebq1K6CiWkhoKlIrZoy0k1XITJLAw852c20qvYo+lfhUc26ffgepsc2B
DwhfD2SFUnlqgs/O5jCDAlkvc1bMR5pHjt63t+y8PPRi98iNwx0KxLlvGSP4rjqq
RMVRimAcBunK4uvJYjzG18aOZvAfpgr9StqbE60ahrqUrZXFruPzfOfhAogh5Bi9
tlj1w203ZbKVHgomRmuF9ZXtzizVdLlLT/EZw86TGackDx3+dJVo/3jHWSYM3eIb
Rqgtp3eHHHfCEkXMqMqw1aByDz7MEQX7ViVkTs4f7+VKQJxlZgtmlrsTBdD21hNn
tlc1itRocgQ7hh9IeKw9dHJPwM65IkTvRkQSv4ow0GIHgsHVvz8gMlHhOXPjulmq
rvE78bVJtt07P7zyGarjSQY+ZKc7J82vxA6Ao/34A12yQzhh4OhH5G0R4W2VO7zI
EijD5x931bdowJCGz+48734OIDJxrIMpyU6cab0YYB6o4SiUabgnz6WHAWaaRRbc
kI3ny+sR7ce2oROVOJQQ0m/XaXuYFZ0l6eI+GpjMx1E6GH04a8YycvzS01h6BFXp
Qg4L6PKbO7eHDirdl2VQSeydAly61D6i8a1VfiwmAFWR0DPDO013zj6wWt2SzZDU
zmQ0K10gBO/syj5MtsHQWCeLfK4bJwuDxB5IJIFlbsowtkqpvqNRiUOdaPcML8JP
ZNbCndGw/r3myy7TuAy6Vf/JlCe2QxnHgXg9Ahfs+Urkevq8HDavPPSJX/zYSkrM
4RZir45/5V9hytQLUUUabSyMq1QIQuSf4T4T5gkwLNhZWLwC38r5SD5CAeYsaCcu
Gf0nbq0KrqOIQjRuSMsA9rKp5qua6nLzOqLwxQcRp1FE0D2yp4dj+moNdZPiLk4f
EFnNK/IjRjoXlWiKrYNRYX8B+M1pr1uSAClTbmrxoPfpEe3FLo3K/WdeQabn3DlT
euqORXVKMSEeGwweQ3UiK0IjkPF/KdpS1MG5XIMWoBMNjKw0HbxNH0kLewjZFvru
N3GX7Vt+EBawi7z0d6XXX2o6UJzxdocBShxUmdRAoXouo+YJ+Q9PpvDfKig/eanu
G/4RrCy8m45DRNWn5W1FrpjFDQLZRwVLP1GGIM5sWbOFyyibN0o+EyydwpRmS2l/
fc4weKhMWULfCK2W1+BvsfmSmBS6A1VwQ5M9VYa2gBkdXZeR7eDsg+19dM8UYmOs
PALJzTHkrwALuaCjI/9v93gAepUzMSgwlZKSywQcRF4awJ7pWTkNbhf5snFLuXZ6
aMeeF+aRviMLpqsnMLJ0hPZSScvLO3ia9ddaL9H7/MfufjOBzpJpfoXWKHa7Z7uP
RY1zmcPJFh9/dlX0G/Zp+IWJL2IIrbyB5q2pm321QSYnRSTt091o9VB8r2PnzrPc
c9sWRt2spSmLRT7DicPDjGpOXfhHeRVRHf49/qoiA5CTMHR6OkoplveLEEc9jHZD
wyQbDR5yhPEAatDlu3G2DxuJSPgdMBeZd5GFZdpCsa30IkYS+qYLTaEWt21m8IWv
v/SLtJGgCdez0gEb3vXttuSYT+ZhryKn5Cyf5YoOIAyFSkDAgOOhIkNlux76BYfn
9Q8dbEBW0VhLCYU5dWOWvsE8kh1dz6ztLMUG/wQDqof0Jf0zKdvVPHFQMtYkhOmT
kXWGWs0+jBzIXUmrOT34ssx/D9CRfc6FIXg1onKMeUzzk3t0wq/Up1YgW1yOgD9y
EJOE6lp6/m5BHsA98fnp3f7qcH+KT4XB0CpaGsSJimMmgPfZMrUxg+0PH7AbeKpk
WM6Or/477eyfAud7Gflarsza05fPW0qrQSvEH7OglxG9IN4WF79z3vRHjCvwMg/t
a90pv9p7f8f0rRlzDpD2gi9fh8YWAE8hjUmV1dOnHPO+hTPGs8bii8yFJxzWXvEV
eiheizGtqx2nk+vJRfzKS+6qjdeXzxBhLUXk25gnZVtSTEklWPcRjbfsDf+PxgyC
DkJi5o/1NRVoR47WbH8FRgEA3rB2R4SsVBQcJVPkZblDvIpsBznkVUJIK8d02V6i
Jo9XijZKDW6yBDn0m0EyYjLNc2oR9NTGukSw3q1bfF62IjK+fAWWsS2farx1qmrU
SFUETd2LU8VunB+23Nku9S2LK8eHfdM1j4g9c0IPrwB74eBwTSsXPQDk9Kzn1P8l
Oq0XhxZBcEnmrquOwTVot6Opcvms3pTH0Zr2px/RsQeC0Fw0yGjVJr+BTdItF6fR
3JTnIlMYa2YinpC8e1JvvPfhkL4K4hvQVVWEZkCTP4+A5y3/mmKpEgDCD3rmMMIX
vwMGci5L5CR8y5YAPXUBgrjvQVjXvLL0njKo1S1SM0cat+3GDTLuyRwcoiBtN3eA
tlgNIk7rjn8BXXw7L2jRoxGhbAYGq/tq6ne7UTXL/vctabFx068Qv0cXXfKi0uC+
q19jfofIpRsNOOXnCKJ+MhRTJj/8PPTwafHu4BfrMwogZYPKWOAyDDmpmly6GzOd
P4zR/ZvnFYtuL77N3XUGIR1RhGz0B7zHueGrDxQ0jITRC+ywuiVYa5aY1WJvCMwP
4ygnGK5JzTyeqhpMlcj8emA3coQHc8F0g+X+wYuAIV2eRGViuvlFy32A+toWPQd8
BACKmHOSstbWTTI7UsFk4Pz2QQYy+lgCO3LDTpiNsvCT5ynucVqAjPgo/f3RnMH1
Rqalcd/v7u6Jpxb45VrEKBLzH/dZeTKRXSuYJt1UnjX4wNB7it7ef/ZQerMO2peT
fLjfOyAgPhWwuEqL/6JkGUBLnW8RCKN9PHE8dQ4xiXdt23H/flNPQUYqQcoQXOrH
dinUUGye1JzRq7rYrwhY7aQOSrmMIJCRD5nS/cjRKPyELSIH1KbxNTqZfx9r2t77
9DMLoIR7vz0BbMxPeMVDwPXIivoLemhxM1lXUO/7nGHcoj+ECt84LFL43LZScpKA
/iCqvIfh6yyFPxwQQoXRTQjTt7y1hzIvZBwsVhQIk/Bp3SL2fczYMG78Sz98aRGa
85ZW/75hr8MftuNiY+jrb0j6KAwuglxs44qP8zOjWCNjPPtLALRQYM7XphpmWHCf
KhHlcQLrwYNveJuTMtDgFdyalFfh1FbIMrRRoEUhIA6IjtKDiK8TlXYP1ln8zb9q
fT+UEhsS44QvjEltIGELJKewDoCrLfOrrCQVEW6+Mu3zcifBA7GaCCx04zmgD+vT
ILKBmbWgjzyWRWRBa2rtxaZMmQNX6OQ9Pha4ifKDQPWr12VOgPYBeAUxK60V8xpB
5luceV8piJk7D9krjIUPwdyTsV6YArcBDMd4fVp1Ke1pwAkaAXd8aG1zZFv3lJRd
MOhQ8ZGWvOR30eo2VhfODL4qMeDHjqKF5c0dMpCVbYDmcaiVSJZLW7V9wI8KmjqZ
yPVH5ulAOzNfipg1amQHReHjAl2gWoBDOzxnyRofwQeXPYnrNqNsRy0gpn1Yrt2u
T9yElOcVD0AspYeg/2LLMTIOXjop5GuELHWc7y+tT0z0YjnQJkewvraSDSVq/iR3
SBVg95dLzzy69Ej7oIdV2qr4tsnzg2Sb7i8tq2MdjW6p4E/uv7ZmHuo57DaRBn3D
M0JBss88RkExSDPz9eLVaVAHLBG0JIGVFXprsmnduhNteZ8lyWlhHL55lyvCiQ/t
Wzua8mM0oEH/PIA9Xq00B+t19tHOlEP/vPuTgNL2nKGSq9X0Pt9rM63xMHt2xt/e
66NAyf3N0z3xdCZ/RYOBc1W+rSx8oo49zK5PvwTvsb1F4Bbk5htnPzg3QPmQRTlx
4s9XKG/y3UyUYTZRSHiyNtpZcFeBGu4QULCJgyvw6em05yiNo2nEUOumAXawL4Ws
jTfXcRyXoTYo9/NjmPnnUrh9EdIsYOfmyGdO9E4uAe/Xs4OcDHB7+662GUOEgk3Y
ovmlZLlQRA8ZoXHglRzQ7g7KEAnngsVyZCwop0atALC1n7YlnRbDlIJFN1OyxA8z
mVz7YQ26YJibgIGDCr8TPA3PHPiBiMBz9vchbb9RdVlBQxGxnLC6eAHtGYQzpG7/
5xRjJs1wjIP30CUTrZGT1J2dgrUGIHbiz4I1QUJ4KJTUAgOsGULgDAnyhHggR4FE
nNbSZ9Y/t9W349LqPtMDZZ2cE3HAuiE7zORPo5lWp9buuwMsefBLyjmJBgBMUkrl
0WDQTqmd6RRulc/36nKTo7bJ2QOEMhMQop8KA3jEBOuM/bgdN6dxFu4tJ1VfYjGc
RLALwW34JwfTDIRxbHXStS11lDmHlznv6IXZadPVWQLExGGiJI4Mk9/UwKbeyDqo
mLhx/wUmyozitDH04MVtxAdygToa8ylTmWfrV+gfbdOHcxtLDd20Vn4l+YPkP83V
J1qPo7FE8lDyPMSnYp2uAMjjYRCfyJ5KnsNmMo/0bSUWElVkUT1G5mOb5c7OKJZy
2Yeu53OLx/NwgJ1IhNbWWU7nVm4fUlrc+Sy/chsX22HFJlm0vaSM5tA8F1nbqZAi
0dzXCj8G2p2JYI1dIqJOi9s3t3px73KWgyy19ykGPUTUnZsM4/px65LwNWnSZxVm
gAzDwn9AWDnxgIMsaNycxI6HAdt2LnORFmy+sGqxI7vdUC60jZJBXXukKuyOtvYI
4h92x6K2TBkZ1i+3uwRe8gXCdnvodj4f01BJZ6+iwTvho7ySZiLxKsOIk9jOGivE
zuwThTf4WpcPVIM2j4U1VYxUaYp6hpNdX53wSyTbvJW1Qed00RTkFozMjXOGA9L7
hrKgvCsfE9aMOVRgPfDTAPm9J+ult9Hhbu+W4GPcM8M+7lbn2ryqhBnwC15O5EHw
eloNjbvXqr9rXfSxylCp8AmNZAd5GbIGTHMFvye2lgvJ2+1YgvmcMDEaV0pe3Fje
iPIpi8ImYqQjzijXlr7Yy60Ua7+rxALC8VN0FLn+XQ7QjHQ1ZQ7i2QHfjDHr8frh
Yrk2nU0yh7jhTZVy4AIuf415bWLHnxN25a2nT19h47ZRq3SGdG2eZFJpD5CHn9AF
JI94BYn6+0Eubh0OBwxc06FLEyMqGgZRv309QEL7U/kB2PxLJ21hYK/zBXcpw7aN
n9do4urnptG+3CacZ+LCDFLhbi5J71p7+O4nTVP81mtGwYSVS0gKDKGiQnVL1eU/
P+OB8J2npTFfZ7j2dBQZxgiMoojCf/coO4itBu40vzRbBSTJ43khW1BqeDyiSIts
cOmCUJEqBPy7mC4cQhFYSxDNj5i0QLKQSxUYa/SXWwvTItcNEFWBbW5K5tjV0mQ5
INmPcsCrDz6ZbLGLr73CttzKfK3BlRKN3aYF6dAz1O5b1mX3HHykPP8gII7Qplb7
6me90K6lgzRVb6ZV20KzdhIEgbxmRgNRp7Ab+xZwksdqU4gUlhi9SpiVl3EV1kwi
64SwqmfZpxMvC7N2uMd88TBaxdZpTRNke+A/WewluDdmmZkpyOWri7KCDlcvCKbt
mzbwHoR1oeDaAQIrn+bvkPV6u+Ad9Pma6FMKTRK8OSOrV06wyFAwuJ/W+ku4e+Dn
NHJovwUh2Ngbr2j/uVdbHX6IKdpXOEiieY/youe7WegQB7lxxMEvI9bbkaN7TSiH
dF+LHaDtRqrVCxHrSDudq7nmdLtoCeCFIGTykdvFOJYwVD/7Ny2/GyfDBLej4JvU
GlxQhMowZ2PtRwEDKrOzrB2Xt9qyqmtNR/muVBGPRpcBLjITj4y8QjtP75MYylbc
6Lyk189fPEPrDnHBtsMvt6hHrQRBUT4eVRuZLFgAWqNxX1kBWO/zoVTBfKwyPXO7
fR6NVccIM74niMIXQWpJmQWIPlEJBmXn4iyjGK5b5KPZY154lGnIW3TF26Sjy1kX
8hz8UL4PjjOCwNNCjHoRLPNQDzea9LXg9Kwh6Hn6on9ISvZ/Q3gaiEp2GILaXx0p
O9AfeFGumpU7/Bn3n1uTdp8n0bQmpZFoKlTsP9qIEbNh4ld2u9K9bzr0B/zSiNDM
Wa/X3D3IxTNBlpnNLWTbakvl4VeP3cukUp+Z3XlJ4Y5vHfG3D2dLt7Gl0g0Uw+gc
GgqDWqJi9Arl45SZzwjuvomKAUOvwmTfICEimylec02Eb93NlU/+Pjgmfa5a+1gK
zVzTAz+gmy1CRblc0VoYWP9sdWjPlxLUvZZ0EsMgA4Qn9gE/JBXhm644hTl3HtyA
wEjefbGV5ljAG8CJoqpZJCoas18C8Y7q6Q8hfUbwI9FLvE4dtWr67S+rXO4pqay3
1wd0c1B4tPl0KMF2tkwKvhrNkQf4GtOJ7asaqwybtU9cmdz3sAsHuE1KF+IPHqJi
cofvsjWM5q0eWQEkkBhkSZZsT7KbrBMmqeTYf5J9luDqQa84I0+tyzs1QC4ybpJ9
mhaHoHOU0Q6t+BK6wrcqcohPNkKE7zgLWWui+yQVkL28TBoo6RGUdgKgmg2MYKPc
t72OB/mnJ47sT/7SNWi9yEJrqJYLoeQRR+UfIVSK9kpdoz44hVy+a8PHgMQWWNn/
AB797FURHv8Ha+nD3i66VPfVf6R8RnGXFtNADQHSOamhmVdEc+2jt1evvDBJnOK/
0yVTqcE4VgoEZvvxNepW/aKFl85ew9yVEeDYBeJun35fcwIKU+Ob5tMfywxh8V/h
geXqfql2SRlRjtlQlw6XQAn0zisdeYyfOGlyVEf/PXnFjaR4AmLN0Yohu59iSaKO
GEyNsLNDT0V0mCj+7PL5zZh9zDFVM697oBXfefa6nwTib5S/hdkfceEjZNaC4U9r
zc8d8fj728adbAlpnSOMdKttrtf+E5O0rFHGTuS8NFxiI1miTSzR1Z2KNTnVzbwD
K2h1HDpz+45jbZkQ1EIO+Ae/SdPCrleKBvf2+21nApnepOJ1MFwWuhU5q4o8m1ys
cTHth+SKedBl0o8gLDfisnqtTofFWxYqyuTLaz6AxN5vCa6U89xiFglj08QiqHWE
IFMi9cKUFjQMyHZWGCC9JKe/YACRMKD3B34wJ2ytSMJXewXmYR7sZhEBEF6k8grL
bgd/nGrUAwYDaGPo4F9Gu1iA56JdEhuXoTIbXW9HT6JiNUOnc5R2skPwV1RPVrPO
IFLNQYoQXKunvMYi1aDRcgPntQDsd6N3VofuE5pkXsFzRH49ypf1aavSxVUrHrRG
YF3NWG9RbXJJtJU2q4XPSICHtP2BAd6tGk8GXzcGHzHTfdfcAKmNGZ6VS3z9pbRs
M/5nT0mUTycSMMUSKmxY+svdBLHFYY0DmwGVDRiW0GWAz6R2cb+jFieJD6RmgA2h
P5CMtVsoS0HgOhgWtmlL9ezTxCs2BLSWKyUHvtzqM8adaIZ+WofCJ1IpdOcy0gI7
fDZ/jXwTcdqABwixpJn12AE93IGtvaodKUpaEwdXdVz3F9lyx350rcoO2IiugprK
iav9nARbTZuIm5G/F8Q1gGt2dnR8dv07134St0vyR81BTof7zGN2i/WmBs0MWq/W
CLvh+BGwYvzxZT5a54HPlKJ9xZv/fcRrCCehY5+zlaAQAsTubE808mMnI4kmJlRS
nv7NgUFQIkdwlCxss4Tq5HUkCtbQ7XUycPUYjgJ9nKJGQAiUipkbAqxIIJeEUbO3
vDbdVj+mrIuJMFypxS7YOh0eUU6LgmR3rTP3Fuik66S0n3+caRcj7JDRyI7Y4e9n
HqSpU2ERoW2ZJhcvznaf7TZUJOctm+FNsUjHfblI+UFRNdgnvw8ZuNXuv9/Pu/jo
i7JWtrxIxI8E2cUv4P4Hg/NXJqhLVAt6ANFd1Bk43IkMEhARhd1hM5IHe9gMgn3J
HHgL3FKp0/ZpiwpkscdNKr6yKezeBDYLwF59YQbb0QZH1Ys1weVO0hRaTaCjmHVb
xOl4aFUOrg5Mt8dLSUMXFdHURr234OcS4/LR8K/02ObO/fbrNMKMp3pAS3kh/BCN
bMZJQt5Qg2zj+x0fKf7rOZNHexAz3AmzEO8EoDlkeNNCU4ahjiggA7oIvRg7QT+A
jj8IEuBxESD3qquoktP8tj2j7U13MAVi3nwppzW8qbUzTJE8OpbUvF7RpAPm3LGF
QXFODI+e+xFfT76X14ozOwbEmUx3Xdp/rzNbAE9UYc2QaY9cfqQpQ+XGoEsLYtgw
KpGZGW6opb4sA8ou8y43rzW55BZo5IeUseuc+Os2d0ah/qiIQWAfa4rSygUXq4Gc
HM3vHU7UgxFkx/IZVJ4jFsL/RhNbu38Kmfu/a2mqsdMXPaGQQJJeG9m/bbVpwm8Z
A7rhlsLN55+/+BrzTktOjFW7yZBqI7mAGLAX6ELW5MS3XSSb3rNcp697UeFQXojq
ylPmjul85ACDK49309RVVnQdCqd3ryw9KrAuEiTXH5FfOxH6CsapuTWXxqJCTN1B
+I1e0KwuobeegR0YGeBkAXbpvcregRG8YABsbegY6AjZDdK4if27AmrXGhQDLHtr
KOScfrKwNcOqm+4NSNmjFzhMm43GNAV5ClJCZkMIUok3rtYORcm1jP1aKf93MEOG
qQpTICoV2ymq1wFuteel7+P0MaWDLqASCtEFGIiIV0EjMUASKdJbi6P4snPDYLoo
iyk1v5yd/L7Kd7xg7xGc4KbNFkNWSlTlpBQtDyorKhNa7n9j9MGev7NH7KejNqGN
Umnt637f+DjjEooEWj5JKKpZTFglqK3mp0exXhu0DychypUM+rHVJyWV84uiYqr/
1D1+k4pjlvE1AM+aGuc1EUvDDlWQtxgvGiyZwo/Lh78q91GW6qd3HeT0imB6s77V
Lo6I9rcnzxFPLzH/FJC0LkWPmwBdYV2OHUxZ+kwBUFmoEKVCKcdGopeSigXg/eNd
lobjvGTnL/Cwm9RYDIOfzwOeI/DtGWJVOxofdZUgTAjSuEQTwY1BIZrsNwxrAFt7
RG9XfM/xnpOJqa3UPV4Goy1Q+a4z48wuIw7DwyGf4JwddcFeNO7QWtM3Zm5Nf64X
BgrLk5swIApaz1g++KJ6FPWR+XynNrwzh1YAlMNhPudQUyQ2/mt1W79dAuoAqRCs
VUaCGBfJekAoNRlw6BQST0r26OirnfzMP48RES/oqmNiRDxNdawBiRVvkpV+o5XY
p2yUIarDydgY1RIDYVzl01o7Mt9VBTcZt37j0s+uKvRD+tqTyT2m9MPB2d82QtgV
3RvpolbAdtRLzcttZOCzoXi+c1u46OfM+sFPobR81IR+Rh9ZU9eHminqp1Q42tBk
hI2XbWimnpEcyK74z8671Nuwt0c0ZrDi3lt+omG/YPVHYKXmz1LipN1FuGh65MCi
u4MPhgFpoi+8OstCa3WcPEwOLGG/9PLRNdtVf0pu1iRcsTrqxle5tYGqXN75zY1o
b2AAPtLknpNmxM0sKtEFPiiULwDnsOVxgzjucalXZyt4I6DRTCNA838Q1SXr3/JG
9yU62HNREwPyBxX+1z6k9Mykjg6nZVBarMsYsP0z1e5uYTafgb2De3VnrQ/2gTwK
ap58UJIIMp74uk4mT9YOo4huWZzJPHJ5GSVFPpQWoEXtbX3x6jyoF/yzUM3uRw7q
Mpx83bJfO3i38/DWyQXTPwxa6ID+Q08Je/spOfbLSnX9U8b5/wPu67Ia6taSKBrj
ONQ16QM6JsoRcYkf+AwY7uPOO5pNAHRVgMllKvnQgXMAJX7/bSqwdyDiadbKurjf
wb8VGHMbstLbu5I6mM/5xQMyzffQkKifJ6pNWD+fHy/C2//h/7Vf7//piWmNdHE4
yymhWh5XwAaifIpdZyBvceOiNr7YMhK566s9fhs4aVEL4+LfBzEvIyGeSfO5DQwx
24q2d5f5h+2XK29d+NgrB14SGs60uVq5rk9drew8rfKjGchLyNx+uTHGN2K8W/JD
qalJkHlC8PaZJRM/2lP+FszltXixDSAhrQtTUOUTlJ6TLgB26gsLmEjyUDDkFWux
BGSji8C9s6GsuRuQfxZ1qK1DvYyHYERiDl7W4E1V+Sg2SY0+hkKevpLxAlKtA0hR
goDh2/JCtqmqrVAHxPPrm3dPQ6qi67iqkC2mSenXkmmvy8XBj3IMQ3X4nE8NWVz1
cvX1fbJ3dcdN/c1L+0s7RTUXd3xBOHy1/Od/mm/dxhTZxwWvIm20lxfwRGILyDGh
5qUoFbaPP5eVXFDMp5JAe5egUYppvaBUpmKB0OH4bzde4y8HyNYq2jLeQoS45h/+
CBRtxpMpdsteQh3aKzYeESkLdR0TmBBWszXwnuO+Nr4LUw74h2y9D8CXzWTbEBUI
ZO0IqLIOLo8ILGqtgcf8h5bB/31KMMyp2bozzV5m5G7mamJUXTUJvfSe1HdbUibL
rQ+2sZl8POtco1kLbGaN/HAwKpdzSg1CLTGXngjsopuufkq/G6KhNhnqdWs1rgRw
R7OH9PPMUSiuT8Bw3+aER+3yxmsRmo15Sw+HWlEGDsm2/Y68C2vz5I0W63IjVGVl
riaLXD72YzDMXYR9JxPmOxcwKbbdxXaUFw4dOicXyZhADgXJ4HJ+6sQt+aqkiPF3
cEF7Hxrmd+zX+lVYN8a195I9YUJHBbJcgebfu5alndzdJ5irsHdMdVcqrx2QejBC
QxFYxk2eo0/x3IhE0AiBAHvAMHQzO/u/SrQ/YX73ZWFXlAGGg4gGPOCjzAf9X4Jr
EaLdlfO495nBcy+ck/cXXL+a5gdNUYYLqXqiPx1DRZkIjAzQ/msUJEVx6snXR1W+
vL0CHahNWwpcmbWWovDRCHL/JfhOfpaDwRqVrZThAoE6RKn+4Ik3v/6FoiqFBvyV
xzjlZevrEZcx9xh1xfopUgqz7w/Q0NSsIReoAhwk3t4AcLJYkdSv/RxmMI6+ewDK
6/BsPg5FIMe4DYhMtOe74MMV07rjdReRn2UBvX4S/y2H+aKV/Sglqo8j5dXHhLOz
kJPaLFSPd9V9OUEvSFXntGjx5zl34c73hltT2XgisNooIJzuy6GPBNIHxzYoeJq8
ua2H41+0n9VBc5mnT4SGhRSBAjxjr9R7LTki3+flJr0TS2WZP0SeBLEBbXVv8Pwa
ZCgCSHAZmcvwm6e/SmJASDvWIHj/7uREeepCHThhCLbSMWw0Wu1NmFxpGq2RTWqy
KldtUdN7haLrV8+YubpteZlZnxVYO7tcNyP3qucmTDOGzTLm5TBIXNeGPu1ra2bc
F9Z5yY0wCxoEJnkPuMiV/YDS5S6elolopA6xCJ4aTGr8bEdp/oxnUQmbQErpdW3A
XQXaBLk3zQKHJa78gJgtMlDxOITphn+Ov1QlhMic/Mr0qCF7qNoUPkGFEBqruPCs
0gDjUDRucUmJaKLZpzVX9yWfoMWpmtCI885F0UzwZEfbsAhISgG1OuNymRFeFD7r
k5Vb9SpH9JfcBoxn+257azyBdVo/H+++b8KojdxmiwPNXGd9apzGjH/MMl8hFhid
Sijffn6xz3BH11wyaNWuDL7aiuTJ49ifrYreOhxe06qIt3Gi6H8cV4RQU5OR/ViC
wuuXqZX0lDAk3NM92xBdDbpbBThb0PE90lCwRaDZKqZ3XELxGZAcmKJWZExa9uoK
dRsNmar/2HkqVhdtD3tW6H4yu2T+uBXArafVP9lxYF4+xN6/g09AiTsFm3+gI7dU
Sf7Dr+U3xHByQKCv+H886MO+y9wZvKEq7U4490F7mgX4qHI9aGonkxwnp7voQ1+t
kQlQag6F4/eBSu9PDSxKgpbZa2eqCGvaHfJ3N40/z72whkiagXas15NGdx1br5Zj
tK9LeBM2/4ckh1ZjuoyntABup7QdcRpnQiTMH3EJqENZPmSxMxZRHRFDQ+YGR/P0
/+Z2GIVUVPKf6HWPZ3ruPKbrZPlxRrLps+Utt6R3AkLvylaILrJgm4aa997GSr4M
GHsHPRZjWBpa1d2VX5HTkP3OzFxU9ADUFvAS4Bc/EJYTr7St4HA65F92407q8ihE
36Jl9Rqh2Lr0sWQiq9yn59je4v2J+wTB1JFomq0mcLpPgc3f+5Zl/22G6rSaM9i6
i7lrIhsKXS/O9OFQRZBHKAn31sl+ESOOUleazjZAvdrAg9JUksdPTpATjvn18UlU
FurXTpMl/1ExlbFrN9r/PEdq1ArbGN8toCZfKLnqG3U60vSwtIrgvj7ZFN+m/1He
kAp/G7Q7LLxvKRaqz+bqILszuJkK1hpGyvo4GZsToAbNVVx59JdCUnvqii1Bckls
3GVI72L2m0SfAtgPPkPciOsE8sns+O7A448VmRzNe9ezFvv59CNO6Ux4/zoimqWw
QcO7IT9OAcdbCL69tqP/TS6+tjKPSBiMqjaq8rCvqdRloFUe/b/7naxkeOedjIOo
szpccUO3bnyopVHPDcbfZkrrM0ul1koKdfYK8kVuI87Ie+/QQRKMT0xkJhdawmlK
zSH5S6fNG8EvGKHtHlEifmGM1Udlv53wnlTuSvveL+AgKW8GB9yjAlKapJAQyEwU
zCRCFV0K/Ga8/mdC1jcT5BKEGVp7pClxXdjrunVQbtu7KpGAprRP+pmcVhT7Vrye
RzBpGVYzbT6VyWVJOImE345EOl0Pj88j4AtQK1TdoLNPvYsUoqJDXkptuiVsSQIo
GQzcUNeLCGqIGiPe7cMkyXHnJJZV/ydgCdo98WkhV/tKapfuqS36OWOK/tlEySI7
6l7wRT2/nWNTv398vbde2bOjIRrwaj1I7GyCLs3LTzL3jv4x61btL6WkR4EMZ1oC
nri8NSms7aBWaFS+yoNubYjw3CoSZOg2f+UXz67kyDLHDygEV6Nfvni/fPmi6kvC
h+mC8gW1AJMYqg6iYxZsL7R8J8H7KkcrngDl5qm86cUB9Mkb0g5HlKMCna+MiF+J
OJ1mERDGuKmL6my393gCBJ4K2H95I6hmf7RTReyvNOsdt6ky/zocMvyC8sEhKpdc
u7sqHVJCX1HdUx2/re4b/l7Cefc6u9Z2D6Hbxd5+B8VHWibNiFjiuOKyQO40x7Nl
cdajFXoXl38QJGXyxhfj1qfE/PV2H34nvbab9YF5vemDRIyrJmnP6iqYZdlU4FYX
idtU1xv7mskEcOB/IvKKQhgfgcWeqJozzUAIduYTFrne2uudlug93R28u1O7QEKz
il6b0zseQn+Tjv40en8gx/ujZ+W9KNvfYXxIt0UUvL+eBRaYScNZruqKyGwB/rtN
nCjm7AIWT6lhGKggaTgU+HdtxNwbgOp3bgnknNT/GUZfxo77YqXnfu12b4tqM9Ei
tMYMd1KS61LrKxQS2fei1tsQWmdaNjQ3wtf6FMehKAnvHeyjj4KwJGhRCfe2K0rX
aCArhgp2BcHaeTRz0P//mtQTBbCgT//ND6E/jl4i94SPKvIrWZszyJmU8pz3Kdm6
NLfpNqzXtkp21kCTQjoTdZ6YWCEbgUsmCGU+HJbIyFl6BTvh1LdHqOb4WhuvGGcj
otbSymVUT7Pyik3Z25BuuQm7nfW6CYEP5QdHz0ZxjWPsNl+OR5kbgB4vN4dipEt4
SwpyLBhr3pvBQ4DE+kHLVh8bj3r/2wc9HZ+n9tXjsEoY5I7sbyK5iOA238bW5b+X
ogmXMGwYqObksnJ2MssGxocNeu3q9R3CsysISGmPe1r5T16UMyxILEUeEsjdm1bE
cUJA9v/RpQ3D+08aEThsKcXJ0Pz9gg5p+l9azNkDT4q5iZed7cmG4QUuXofY5TX1
OO82RWagN5ENAt13iG5yDdOHIFqxtW57kSHc21WxiCoP/fGwV6p9CDapMu4HOJtu
+ezxBlvZvYZX4SekQz86/99wF9lV1y0DqY7PR24wgXyN/6eVNSzyWv21zcE+qoXX
gsUri8663Zl3WQ0ZHY2S/8inlcOdt5Ll9uIKr2na7DtseVtYyjRSk1ZVDruXK+N/
Tc4rwYm9VqpmzL8rF4x4Ptx/PXqfKuHy6G+UhsxTYk86gH++KQCS7tO4MHt024yh
AWuu/DSodtxS4/yjocp7QfyWHqwHCayq/U2bQIyQnk8efD1ftDryTeRhj/aZGApO
krmOzuuuVQDpb+lhwOLx+Jbf/57oHkB0JGyO4IlzSIDvR/vOohwV/kc6QZKNGdXh
w2rcYkrehqQeCsmn8KgYbxM/QdBxfF+Cy7pdumZkjIZmXFDI9lgRNq/bfJq5CG7Y
0lICKVIFycAWaISa6B6Q+OGg2BRu2J5owcSGRknMs2oY0I3I9n7ISDajPhYw9w3B
I5oStNd+2EeaH5DekWv3NfVyA0r6u/rDXkfgTxd/z3KRxrGh6ZbeTL8+yE8s888s
WGSGMbTh6rzQYzKVuyHz7zGD1pRJsQMPtqpwDEFxyBOTlQtjWHRGMNucvK26TDKt
jFGZExc5qJnvQT9vOhdZamfR174DfO923Ur3X5MCadOKCPpuIW0D5hIPm7zuJ4Za
/+KkZa6khREe9vG00fZeQ2s6UZhalIVehkl4NeABjR17Apbld451o4jW66MHW4qQ
vK69Ohu7czuAxDsn45cs6LKiatWkSzrhUTma4qytfz4TWQOh0yUZ9dMwyQcHLw5c
NGHCfd2g6/hwgrufPGgXcZpa8If4ATmekrqqflqKkkmN0rZqzPstDRV1+QbcHxir
2qgTNeUmnUTd0I6ygGgCAl9BEkyajmGP0NNryEWDgeOfz05ZiLj1v+mVW7301lK/
kofkeUutuC5ogxdLiu1ofpKMksP4St8Cn486QYgtSjxhD1Z2AxlLhhFhwzbcDa4x
SvleTX/BzAVh2XIaZMfI4efdYpIJKWhPQMwKAqWqR+CUPOshGlajNxjOq4FpcLIe
CrYUGtxbOOIjxrm3pI/wYmAN84dj/HAqbhXrB6AhMuFUKAnyTJpvJp30S6EkdVwm
N203gTcAWY/kUY/ru6stH18E08ZVx4XaJLokTpyDWVe/zzIWmcIO5IrjWmQqk12n
N3iYxsXLd2UJFM4TJGjVw17NUGNzEh3DdLMf/WfXXQOYxfNJXugT7Oosm0LiCeU/
aDDlp9YU4KNBUeEKUbBETLkhXW/3PsRuDJYmfWyMc2AlryqGwNsUEismKEoynODf
U3Npnm4DFmXn143uSxPm6oJaVdpyHz3ZMKtAM8/TthcHIYvfa8vYyXEB0R/JOTBD
WCprSUhWbH6XGiQA+ODMFoCElBF9lAMrkSQdyzbDZdh/hha9A0USRPxy58CtJnbj
kNjqMTiXMyEIXH9QjAbb2uXwLvY3C3NmqNGkOE61z1Xz4Er1P+0tXHHJ45tirUAT
UBeKkGgJQcvEngfSNX5eLLuQkFHfkha1i5v8tIs8KJx2x/KgLN2z9NKVD0kwzrZn
PzDAbLgdsh6KhVDyI422d0cUWGHIvz69YxLpmWnEZhn0v7y+y0Ym6wpXPsAHKepe
sazl4KcC2fbev+ce0PgxQAtxeX0XBL9AhJgTJ9P7k2HmU0AwK3jl/AaBIr83jCnd
wy6k9und/yq5alhnA9rYquP0r0/1D3kI4BtO/tuywzzGmpHg1TyRCwiiNsL+ix+h
PbDeaCmq/wyWG0tTMsnTS143St4/I2Sh+WrGL2IjC/kx4rbc3HdJNfhs0+0vkSP6
nXWK0IiWC67a0QQJuLT6gHy2/ECahOyQOnlpSMuEGaSk0rV/s1IpyaBdpBSWwh2H
6nUUEfulNo6iogv+WtwK2d+bxtjbfprPlsyxj5CB4gjHi8+Ze9xpr/t8lLNYVQWk
jv/Ir6xRfRArrSwZYJV7SJo605pkcLrPbor/1PkZ5jstwREACmwTs5Mel2Ua2OMk
gUazRNu0/nEBal7LXaHgAqEa771Kv7iXf7ztKFVgkeA5TCMfbLNtm78QCChWtzfT
q1T88M9LbiE7W7DS/t7l+lS1fj9kxLr497SspZWJi9Wcf6GU1GrtyilaDs3odltp
ILU0+4qtbjF0jxUroRcGpJu/WlgOD3A1m+leSCqc55lJur/+cFQg/OsXYn/jJ47Q
tqkrM4QmsOGSyLvN4SeqH+euzWtpMw5CCo+9K0uzruLnwjJyuT/XbFFiS4HoZ5zL
lB+b73eZ2/o9+5Nq0u9zHrcHKw2S5lG7+cuxuWkXvxI1FTL8Te9kd1yES3STyv+w
/UdRo61rDtrL9l84JMqZIHQK+wYOKj4yJWMYAEap2oBRDDnQtFacIhezoBKPuSM8
iCjv+cldu9R/artQQxfK30KD2Q6QJT7VnI0LI+NM6StsGeDmOpfBb8fotadNzO13
52YReriF0MAc+ckasUPau/MIhklvo6C6N7AaGMeglOA8yIbsZq/bMip0OBQn/vrB
wi5oFZhiG1KCaXEuZMX7wbd5CFAALJNlUU4QzSh9nBL8sWZUpYdX6tAX49c5xuPF
mL9rLwCxG0mY8fGtDa8XorLNfHDxSv4taUngPONlHTDqr6g8rPxDHZ4dD//bDWVC
xY8bsQsB0TBBE5wXQCLxs3jBtOBygvi2Adh6BZNJzTYw8URTS1eQ2ZJGSdadq29W
tRbDYpD/hb0BuC4MYIZeOQpK0yPcfY5klxgdvLebAN7d6gTL2NYvW9jLIXwHbbfC
gKbQR8LuMMI9xgH2bpfM/Gl6ITNLvHKgR4bcy6N0fFYMnpYF2CVsaCoMoCMm1Uqs
+r7JohBtK5+V1yjBr/uNoApGAepJDuMjz/w2zlCEauf2z0dULkFP6MHp6POxzxfH
KeVkbmCi7JPPWYU96Ay9bSHkluGo+1GZk/8KqJf0xXlkv4sajZ5AyOEHscQUIoXB
WMa+vQMvIx9Cpn67SxgHolC06ts05cRUjSqsPx8k81Y5dmq+FfN1GX/DQcBpCoqj
Bb8zQ55fZHEUC4eBw0VzEt4Sc8tcnj7gAe50fufNtzVV05afgc9mj1aeiSrp+eoG
BUfJtAB7HkrehNF0K8E3k04bgQVyTV1BRVkhTc4KaFCtk6nWzkkzij1UZEDm4IUM
qz/SndRgSycXndDfZvrldf2uRS31BndoOC2Zb/nT5801DFWXpFvIdM2HzvNQvm2j
Z+rSU9VnWaAmQjaDuFA5CCV5g1miaHBmDvysx/tkHjaHrckOYIgZKOgVMNlPqnyB
g6UhgsSrVYO1t9o0sR5wjdDZAQOu34M2q3zrgKDqaejQfSSNipSgmCCcZapYgB+K
k+IVE78PXt4xiPJJVPTXDyG4PIln92w5SwMoPeqDgs+HPLNpKPhC3tWV0pAfUust
FY5VnbevJNuSVbuwRsrkko0zXA1lSZObCnfk4qdodFgtywwdpW6LfdXg7sCba1Rw
nY1SHnWziOpsDCJxFztHq9iU7mSzuaVVK1z3u8bFh9p8VdSC29oj1eDBiGgjj788
B9pZLQu4WnWa8UVeXKNpmHBAp3w+XU5VAjF+miZ4h5Rifoxhi9PPkIfXPGrtM6Dk
i1JQ/KfZPIHuFMXkc5VIKLxMON6DjrjlbNIN/nQoquLCcKdQW8ZnTKxSuGuFp5ec
IVmQBrJpYaWUavCaV06x4jwcPcqjVgYtY5NbkrnrFktt13h/tKoyr/P8VZkwtdb2
0A/WHhNhT4kPLqRm06zQLqt4bATP6mPcjcvFbroHYV1La4GPH2Aj+hyL0w2aZcmd
1pzcako1fjEAgzqCjARvxrh1KHiPv8pmUEU4jU4xVX/004gwPdrkcou8gPP/dueo
rYTrciikztTghW1tE5eNfHOcGjUgasp+p4TQ00uOBQi16bPqqojzJ4sHd3ALP17S
DhAU4W23IcMtMykuEV5FSjJo86QcEdCueRJznabL+B8rxvNQUz+Q7Bm3+Fk58XDN
UeO7N/5zKMRVxZ5CGj0UBteAPeU1MOodrCQXJCcwZJVqaWRK6xqpy+NOehZbx0LZ
B59xGuOleLDIbPOz1XOt5MIdJ3bKEnmCqWeYtJkkP4SPjVIGpBtxkFsWDSX+5ftT
LIXnT/qfLXn2clH46IzXlNpHK1y0TPzsd4gyyZvRjGn98ekaoaryvur2rspsYJNi
QfqnzErBp0oan8CLBWfawJaRbuSuY71xZG7Ar9c2VYiaKtjXxQIDv+AkKSO0N/x8
CWw8EGMGowRJNUtoM1pqYARd96YqfAaftriCS9nVnh7Nfhab/XVbrwkfzHYqhcAB
6vjnjphNC0dJyD8azosW+egGth5AyNiwOa/09V/MjEdG+I3BNwPPksoD9Ja5xo6l
+TZCZCgD8Z+gmS/mPnrC7R7vJ81p0zWGTC391WAJu1LbYcVOrOOyA6LkuwrXMums
tqltV/8bDv96zaHnxPc+XfhnXNyTufZInri2ZjkFc5htBZqGWEVejQD/FAUGHjXH
FduR6UPE1SMmNL1SjqNEjrr9gTuPl2fncIw3kgcTwluDpVaOR0BK/07uMKr27AjF
aucIlrjvvDfQ89Ova6RtSGZERxFGpI8O04Cnlvic6uYy7uFq8wGPsld7WyhPZfkI
7O7Qbh1OU3ig8tYmvZnYhl7RNwajnKPYNozSDHhjjPp1A+0bO8D8hZYDMcindWSC
CL6BWAXLK4SHCPrqLS6kyPHRpGKI99xQOoJVuIoLMwJ3Kq4Z4xJOFmyqGSMDVHWd
GySqpATh0905yX9MmOSTreX93kZDWnRVsRIaI1rDv0lYTsvR8G8Ix2HvhcewqVjI
h0gcqOGcFvLLW7YP9m0EGg6mUkoxcvQypf3ZgxpsAwkxsSTOID0Jh+Vex/kR3d+B
scSjT5b2kJx0ZuOM5hdpdpwHws0tMq1qEUY0SsQf6A6VcPyNYEbZniMzOBYAAsA1
lNq+NYZjU57VZWI2iGE9KcZ73uoRaPI1s31gNp5SFuHj/WmpW8sPcFvrLRshmEnc
G8qn0VTSQnUigilGcHHwaijsz9611j5YM8p/SQK3MbDCSfb62FMQvzREzPxoOPHD
0/8mlMTKORLmdZrWf3qjV2WoNBtFadYodYKc2oCwzE1ZXNE4XE2osGTO+poH6PzE
cmT/8u7jI2kZwdfSvHPIW/XL0tRB4P+sKJHWArExX1RCYk/w5UpQML31FKw2nKCN
L+N3OmRDxlnrStyjziKDifqvZzDYRnI0OfCYAHIlew38hsx1/OE5RhJjJaqdbbto
7DWFrKBTiTCkiU8CeRQaUg2oXcfSHwcuEPPXGS5SLzwi9EvZZAXiuiLSjq8bUTlT
IXsavTqoV1pv1iGZoyxvGgpNsKvZV6x4+XsRwgn3pSbXburKZ5wIHMO58wAK7vRu
nP5SOHmzoWRrcA8SKa1wOYokqqc3Dbot6Lh6IR/rKWEVmt8z5Iwo1bT0BT4dJ00h
1ifJ91SWV8f3K0uRUMiJhAWiSBFSIC99jRjksx79Wuy7q6IMKmPjZQeb8y4+PRh1
d3XI609Wk3msL4FRfCgZyw5e6/hgdhqII2zXVXMDuvUN/55PIggY7dlpXzpVB/E0
OefHycCJKLGiu5QIcUKNoKFd9W71OYD2+N9iBITZuUfZN+665qje+rtAKZQ7lino
gJjVUSPI7F3jRCFVb9EYdGhxR0IzUL6CNypsURLdH2TQgmrCgBl22kAJyz5/nBQe
Wa1fKOVwzNSSe9GXDrz4paM36Xy4hiH/w4oMYWefdQaYcO5wC+pXPtTvs2C6EBRx
mJan0GwXf2IxvOWMBw8m3D2pj0Hcj8xm+bmxz9SYvkOF6klhn8eVtlPJ+LhBjLC9
evg9elkARjwVTrL/4+HIv7aSKmRW1TtjJlL0ocUj+J4pSsKD9ShhI4tLcJ49C5/P
QjkQaa/tgln56sAsUo6Ri0kj/vyo0NmHkvKdaAo5f9tbMvlOf41BuUwn1jMxBvap
Buk3w/0LtaxoLE9VgYjNP4PB7ZZTqC5n4684GqUhHHrw0hLSjhLhAcFK4SaXQ025
XLTtg2X62ZuGfIeGUZGDEayPry5DSCGfHa1nRkfeMFgnJvbJbv/DVxWJFYpXldk8
XPM3Vbhvf6sIwtYHR8oYEbJtPFy+S0eKD/Cu18g5rFtVyKZiieXHglTtET6G4Iid
ZaZUvF6wFSNSW720pE+x1txpl49+w3VV8W6iQC7iIQhAg4F7FJivt1FNdGKcdFDO
dUtSU7HE9QOuO+/gkJA1qlVc8DtcL/hFf/gq+AeQ9TPrTnxuysv31KA4KrvnE3w2
yjyTwANwVOW0inMotn/rTN4Rmkc+FJWHWYyG+LjyIq8xyTRHpFt1wBIrNJVvjWCR
7T38HPQ6Fu2aCiGfAifw6FbecNQNgoRwbcu7GNPS8I2YtA/IAvkR0AKgzuW9pt+Z
1JAxWA200QIBX/eTjf6asO9WQJfuCcv05W1oTEMU/9XFG66B4yNWTU/LKnbqlD85
0DgJ/Pg8nZs+W08AVJn4t/ZKFG+QSvXfGRB932XQ+vOOpg4RH9GP1feF6Rc53e23
v+s8/yWrYdGXnimJ3VG8N+OdGykrc+B9ok/fY1tBmPncOcdqKP+yumICZaLyoUll
e9kCh+xk7+rGwMQxDC/SETemnN72slg/RQ7FS4mIl6Q5ltS4/of6C8G4d6Foee12
Q+ZiAi1J1ucOgI0VaRLX5r41cvKob7OxYOkfkUBJMenFF01m2j0VCmTfHDnA84rl
CgurbV09g44H6/hwRw1VG1RB2iNo2V5r6vsJSzgf+jGxfcEeME144e3qJuqMNUK7
4+GAwaMdowiMqMH57LqDHG8OARrOjXv7UVIiMe/T68JpAQ8zW8VZqBw6ra86nSQe
du3kmljHbXWBCHrdY0xobe5e65insHVr1mjsogaLXkV7koCR+yNnrX6YOtMTI4ja
T1mlob08FOgsSZid/Icwfu4XeHsKMFjHh9WMVtQBhwvByQmawxz1RPZFkBk5GUOZ
1TxMAOvqNvtfPYmDKQzKPBKmRBDgsRYiUUzwDvnmLTJMDf/zQN0AZoloOr4Z2inF
dnLadl2J6hAdwLCBMcvSzOXr2SE9seh7CgNTIpkSpwCWrrPnQwvnaAR7fMBIKspO
E107qwFe8nCcGaQVoTUF2fEmw0VQadTbOxnQeFZ5RSq3eqc3csT7eug8rG4Ufe2g
fy4lABm55E9QP8QZxFgaJZfsCEgwUvPgugDdm5eoBnN6op1L4MNn2KeU3eJD2+hq
o20uYxMoEQHNCn/sqD+ML3gymBWYSoWbWQo0s+rewzmqXtaU76gesstsVTFjpBLq
CdM6TdDcmnju0d1OeDe0hOGPHYwNHHWCbWkA4CEaWxG8gwYPaih5fDqQJv8jLSGJ
RT2d76GTIb5StPbgbIjT2yfri1LFmt1UEEOiSPmxn4w10MEz7uwKXL6Y7gfDDjWE
HxwudFRLt8ywsvtdeMIhZMc6sLpbb9RuI7KD7qA4mrpWWy61Y69XeLaxGDP6M2aX
VTIGm6xVJ7IgJuIc5+oGCsY4wA36W+/BmnxOLTQ+Zx6GW45YlvIP+Pl+KdU2NlIf
NA9RFZLKh3DM31Nyw9g8u39bAPeP6VOLXnMjP50kAUEgWTwTzhSPpdcmgBr1AvLT
1c7kob7a4vsRRtt7BD4ccPt6KjyfhTmwtsJxWhba1OxAOvU6ieBmluFF21Bl1U2q
PZ79sbhlwtgOWzKp32u2zrHQ0S6RBacqCFsU7xvWybXZe/ff55IF9xv9Z19zzkIp
u/AfW1IujzRKLBP+IW18pvMQzumhwy3Mz388V4WlvXhTjzuwRvcbRkuF6oq7aDKL
Y7XuHF0bCYG035KuHxKkhHpXqctpQSJCahEibcrbWTjgm/7MqKXuP26UXWZsvtn5
khrfbbL+PS2KJYtw1ap25H8NDP6DLwjIgmVX24V8UMJHIe5Wta11MOKeRhJUuVJF
/U7rnxjnLNmNnJdyzjMLRYlzbkCi9Q3BtwidkXem/0LjVgTTsU/9Q92UUj5vP/pH
3LeyhZ4bmKmeAvYmmWxynEkW5vCruQ9lRkGJrjs5twlKtHVarbLsQUFUYO4sDakc
2frjRdp+ucmnO9R+f0JrdyTChpnHiaiuVsXQ9KRUqlJENBy8i9XSPv5D9bqZuUWV
nHSZ1GGadTwJD32SKmP9kbRBRsPafNBK7JkGtL7OTnELi/j061MZo/HKl1xNMYlh
6se29W18hufXHHZ+ikokLB/bxVotxyyAtjnFaS7UbiPeP7ATknSh+dtIcyLonjnB
QF6i6vSlnUmWdnoZ+7hDH/GY0MgqcYnNH2PL2gfT33BJIpE5l/941a6Uz1rtqpir
21T+W09z/84DI+Go8J8fwAVEDnXkOkg75mI2Flh0m+hhLRnS97/UhoXitJf2bhfn
UYFv0qE+kRk6vQnaH1TcuzeauwzYMAtwqY49g3jQXwTm5v3rNCwNv6DcUE2bdVsh
De/vWZsitsD/YGdAoeaVsWcpiEb7mMZhi+V4q8e6A6IhTtYANdk6uKpUtLTuncOi
b3b5/l4BtU8OkB4+jsYWKmK1tfpfakN23b+DZJeW+iNyhRvsHxQsb2h4OCLN63hX
YM/46CbkTfi39STPN7JKG3SfeqDQ5G2KSc98wakD0CvD4AwwghIj19DNNR9FKfqb
ZCYoCXArjDxdKM6MRAf2j9hk9nvOHyql6bDtS9spBptS7VkMmEkscJH692xl8MKT
Sw9LuTQpayc/Q+mOLLTqzZLjJKlRtJOs0vvk0jhWtRv8i1OEkCz49NcyNYDkxd1M
ghYK79nyTYXKuiLtG7NilDGIxMQGN7yUi2TyymnKUibnec2YyogjdwoZUPe0o0rs
5fTmYwAWAUI2sZipNcDcaUZRnpmgtPrIsZs0ik9twYl4Ka7+NsG/PEE1g8iLzejN
Co83fFma2WAt75bfzyHDInaqp7ciK+LM4SW7ys96EfcKzfgj/NNw1IzJ5AFA5NOs
re21fFk0Evjw7rKrqclScxaSuZUsrB0gIVYZw0h//xxknrDOcXo7WhJSNNJhqNND
8Wusx7Txxy2GNaFw8XksIjThovskY4DHr3E+iVKhnm3/1YH/6aCOasTJSy2AF9vx
sYtM/VcDkh+uHin7zuDaeJl6I3/Zm1ImKBUOZxg9pI6aWiV8+bFbSD5p7YaSGO6f
HaCNo7vYosPvQYBVknM/GlN0UZ/8LiRaLExfe6XjUDVn4qRqQLtqGYnBlAcfezPl
d2egj0Qe8Zmx6VMT6oQ7aP20WzMl/h26orXMwGE5yaN6mSfw+CmrXFTeyha1uUC+
IxriKen7k7uCXkJjOcWj+V57Ed8rulMyq3PPkm3JItX6/Orv1cwlW7S06k+PySXC
hPmVccjey6mrAR0ovOQKukbCuFhNGcxJZnMC5tY2p0qgA34TTuyz2AzzNp3XsVPu
LNtYARL4z0FtN2d/Do9Jk2j/HqTzXwi1JWFF+/J5E28I9CaiyFKBcfwMzuTG7RMs
rEs7oIMl3X/CMZduuB+EL0LuZrZNMVGbKMxOlOtF8aGsHvuIS5Y7NBMsW2xJmly1
sEfIYy/GjMg8ZP87YDvYl7lUNnECfMkOa4eB1WqOyz5fOmmhmD4Ehk7pFo1lN/Kt
Os7t2obC48MzKO9itUrkhZD9ihRBuQr0fp+PAlbuvfExNyp6YiamYSvuz1aAMEvc
NyaTgBrVraV3GjmrQl6VqwXSltRaZPWX1M3jMYGtn4tql1AzhM425l9TihNV9yBK
7LFosvH8VSfsN4hlnyfRYcFLoXYDYfMCyVmOTzY3tX863tZlXBPoiEXlvyA+Tl5u
zLaLpJcO2HraLvZXlYwlUUAbyxYM8ScegAtk3HAVLmJyCkMjeVae3L8ifcW7Wrrp
4JPNNiLqHWLa3vVs0HgG820mzKwDVK0jucQqaTYAeL/jQfsgcExJNYvUOtdtSaDA
oMXpJGfJhOBwS73qdB3z6deTnbGcpXvlddwYbuZM14jp7JXjsX7dJoNDRN1VpSFP
JHTB5dh5gwD5/wvbPuWpy/SbXI1ujmDtNZqXS+Xo8dNhG8W+R8hIWZCSDJCHrAv+
ig0ZhmkOdVz6yjYDfHbPQvg+8v8cFIzcKK6Aim2gCE8i/Sr3wcqGs7QADFZ1DuEH
cJx8UsFB0FoG2R4UtgZoS7rbxIQc7Mj4+JkiAAzzfSnW3tPJKSWLLFpEpxnUTKsD
FXYLcxAn0bKx9dlFZXWu0Y7eQ8rgBu2q5b/Agkt3eVGX2+bY4GIvfhZbiVJhaQmQ
gp6ggge+zWtJqgZjSSJv9Mfb56Mb+fHKiRKNLG1eCmkTEPX1J/9KV5dPcfFYX0fY
U3tkg+RQKbICagVHkVXixlKimhLn+4LbyovsniQ9jgV9IybaBc3yQlk5zo/isf5B
bYP50NwtBai5ryrntjV7EgPeqt1W3pBiVetPTZSRtt6n8D9CZhEcu4bhixIRDnKD
3YT0t6Mgl7tura7r71IMC/W5anLjKbiyDyL4bvugaG2w7zBT6AZnOR65mcROWy03
nCvwCqSKVzwbE29b2gvGeJBeBqDOyeURDDmKV3MYaL9CxBRdeiKxnF6yHtc9MfMO
IPtqEvwkhZSEIyTBGg4MvSnhqdQVv2JAtKeQL87hgRkPoIQ4Vq2Z4LvzlMnu+01w
DxFxORrC97t9gAP39Ry4U1HZy5i35tBHMTVZgJm8EV6qNUBUa2BnhAW1G9U801pt
Irfom6gPW9/byCTPM00J2P2RrH0l0gHWZdIdhRTvgKIquNqS8o2XwCBvQ/A5r2/z
hSh8NHolJ0hDCRzuKThQCz5p0Il/vPbxBeoMfDMgyY4vXnnmH7NFdz5GqRXIGF+I
H9hslzZgOHfH0DtgmbRb5Erx05pglfvgYrj5k+MfQCV8y47m2aA31hRCgsmcaR1L
HwZSLsb01uhj1xJ72iZswRgCC229HdF8rsmwfTPfYUsTPMe769vz3iv/QTw+V4rA
diFo0KHxa5/dVmeCaxg8pBThd/YVphff0tJ4lJLrr7688J/Q1K9s/wqmVzu82h2H
qj1wqDMpGHRpELFZhQ/EZjd8n9ui8rzJePOKdy2CBNS06dDu1X4eN2v+0jwfiFj2
RAIQq5vz0ROy0JGYxSbzhoWl1fVHVrmeiVrsn3Ci6O+0ydcGMdcl9I9JBdiWdQbV
kut38HzajKvRwkZ1vMxBwyR+PRYugbHWMYTP1/EqYZP+zgt/VfidGVKZxA+dHqDT
SnX7dw0j1mGUpfSW+c0WJZ90LJK4Oqt8vvqIAmAA4k5XoIcsLnTzgoTcvWRgj/bk
dEav2JQIgo7ODjJdO4/vJ1MUSq5Za/cEJAP5u2BIKHNtZamVQmTn1lDJbj2wjipo
JY1xpK827s69XC+x2itlGxrdAZZ2yhz57rNpEBBG8shdjSoZeiaarD4E5z6VR5LC
3eh07FdmsZcx4EVxrU+NKATo9fNY9WE5b8Sju2gcEwXCmNoJInmw7t9DI0K5zNG8
LW3h523BLnO+Ui+DxWm2WwCewjP+7zwCbvI133g4/XE17IOX77xAaVKt/RsIseoD
+Fwpnv1QXYPCZrGTbKbnyhGFAXhmOOrSRvxnOvUtWsUDVCwNyBZm+qpIkn227GGD
BsxynOII7PfrsnfY0TgDO9SDJ9q6eCsfazIqryUyF8YeVFxU3wLPHuw2FOWwLMMr
KA2M4MiQkn2H85ETL8UnMMxGsziyhxKS5golV86r2ECZ5hyPnsfhBtLN2KgHyX6V
0buhHwBJaIMlWefSaE6cA2kgKdj185miUHZl6XYPbeMZt6KmXhvhJXGx9oUFpmAM
3hI5Cb6k1qDc0Z2/vfwwSesvE+/qdq9C3o4muAo9fd9pE4MVkBRJp4dx3SlAt6F3
fNdRQX68qlUJVYpd1FHjHi2vG/bNtOp2k8/MGXnhTifOu/Z+D+ZUyiq9LSbuZnxi
Eq1aGUsCsKW+3BqqD00RFqo36DKmAnA7dsOdJNg+Ta8E0sEdTXz+8pr0b+kp/0hs
/j6o9memobLcS+exl3isbM3FvxGcrEa71XBTZrxThBRuRrE4M9V9bx51PSsR/K54
5f9ZiNOfpUQbEd+4G7NgLYk63L2ITZU3rTvnA90Zi7RvqrdMUi7v6tdFRMeIFYAG
NAu4YCRLZ0fO191b/9+gCGQL78cCR+mx3iD+xRy+GASrZzCmssO3Ujj7iIRWN96x
GWXjVajpk5I5/2cSCcw3jS5TWgaqxxrhqdyANaMrCe/7ZibSgQF5czgO05YGun3M
bA3DXwOynsQqKadvD0H9broGhEHcWg0U8LfmY2aHxBdYq0IKfgzE3P4FxGT9KDwQ
Cn4bpXm24BfzfsPCoo5YaBmaaBI4oCnLBID3atIiXT5U6X0pLuqAfVA730ffHORL
OmWhle8X9pPX9qd+skzpoEGRR37KJ+E8iVTq1msK8hw2ErPaEZjfK/dw73veLKJ5
jOhd9V/hf14hI4EHIsEQKv5SpcVcOljQMQJce75Q8WIy7eVBwyBWv3ltl1nCcdA0
jGe7fmzqyWwWf27jUZTJwqMWsWjo68mBQmQSNmHdjFNlPNnx8ejVSrg1ix1BtBH6
U3PA+lMyUw/27BI9mjBF88Xs1aS1TnEzpTcka0qql8+4zayg0TUVfOhI1dyxNzgi
cisCcNorcgYItlR/YovrXKpHgto88R7VqrYR51dbGeoEJC8HMXDX+42raGNRlwtv
c4SF7xbGjitYGXN6GC7feFXbzNqGCb2FQvLEQFsKDv+E3Wm6keOI8SYC2yio6WIL
kCRF/0hJtOk1khyjFOOzr4TZQjN+b9kJJgxvY2USDgOgfwsuuOFUIi3dZh/89hib
NVN2Fm1ZvuUABJyyPlAl9X/BVb11VMW2FSMT3CCiUeW0zB1nh45CZSbV2yYXRbll
45M2NAbBUCtuROi2a09D+0lXRbHOMSp/xh8lQXrNIpQeQQLB/18l349h8bKfPljb
cpwsvaN/Pmoyq93Ca9WiHMtYtFsSpBGoJ2vTUAZpZnWhrYHjrkhmfPlGWiJLfuL9
/wgH2p+TJs7nQCDdDEqPPrL7/1IWUxb+CHp/F+qZaHltxniJckBJf5nHVWXCo+yy
ueDKMHmIuX9M6JkdY4oyEr3WyDeIwVVQRt4ynbvrKgEokMxYXSqewLn6kH+wcrag
xNyLVHAxhm23cMS2ikdz9fwWbuwC4nPeKPEJ9J3Je1++B6kOLldeEyXhBGL06A/i
s+5uzUuvEPPEY6t9zdyukm35s7RPUJtcwcIQ0xZqJNMN3XGdlkKxYZh+ifjB3lqI
BoTHIihKMkrSQ/0gtcey5YcbMbJlv/NflSZHhCtp4cC4qT5p2Eoao3UzQ3e6wG9N
4gjVWyfGxCU+84EDdI+s1yyWibmm9h5ud0GfHZSexsnFtikwp5rYrLuv+CIsFHxF
5tBb9YAT0Z/q0jZZPFwRqb9TtD3nyspENA+c0qlgn4gnYsX/as+80tUiOy0PD+jF
bZeCipmL8UAA+p8Si5ACCU9+1+YmCu/2lOWPmFIw1FWl9I08t98Hm7I1pb9Y6jT3
8Zu2UlhNSNu7aw5x77qEkoJ8R1jGZzPxWIEkrDmADRaFlNGxKn8gXOHKK/OqlN2p
Sl/SCQUfbQ//JJgsCLHbMNNcu+riundA58eK97k/fy1kQ+e6kbjUhTuvZ66W5AAM
Sc6icw9sV+8DheG1tqGRZaD4H/GF2Xs9xZXoP8JWQrpQsyP+csZjCelfXPAKFQVU
WiOZIX6KvkRmPnQinp0AQ0aAcjYbp8NCI6wf6hqWXiFChX68YAUXBhFzK2oNsb/Q
HGFoeOLj7y6fGHCZhIIzs+m53+nEiA33i3tV6KoaT7H4gD+/ikEA6mIy7EwASOgA
cgrm02jPwHNPKUxlilrAlrUwTNN6Nt+q1EHJoFXcmn3F4UgJSNHO4Im7U0PcziT+
1867LjUFOmF6Splu8wnMgSklndvXvGyH7vMK6W/oFhVINcteW59dle93a+7fRU4c
hEM0ejAdetvibIyHmq5JdGfA1K+IigI7u1QGW2YnsM8V7xN2Zm6wllNQGaU/Z32u
Lc21NUz6b9VOANZ4FCIAsy/ZTcCV47yrTQ56Qp+082qhFm/Vo6KcovV35tYnI5pt
BOP8cPLDqoDjhpd2Zf004rizQfGzIiO9R0bZnOyz1urnA52XdTTld5jbF+MZN3jv
9eXVmaeBC2IJ3HxDgsGEI4csxPClkTMYYt7EtRHPOklNdf9pJttjGec2h5LUoaDL
fqtZXpvWtuHhEBNnuWI87vBCWB5UFlbiu4TfDBnl3SPeJCsfN2WlaHQMF+33oUjD
EEajJEK8iLBwo8Lu+5L5la5f5DU7zn4RkveR1QYf4Eo+8rxFcOGxaQVmGi0Gx6/L
JU4FXR4XRSyXVNw1mndgiKWYTmqlT7XTNp0DjG60en37Infcg1OIpkxDXud3qBIC
ll/jyg7mp0B/nWwOq8jFileeD4VY3LxuJoYJVCuaCCQvahDUuqJfodNFB9Y9ogMr
wwV6BCNemZCiJOX/Jshec5R6AT8m7sezXgPfJELQdeI+rcBl5hmBLHt9ETFvmLgO
0KQm317/PYabvikfJ4pQjZIqObe4sk/odxlGvuSAjkooN9ZNlJhaVE9nleBkEcnm
w8NYOHCMKNh4GaU0j+FyT2HmbwrBpbFdQu8E6jaZK3eISu4uLB83HfkyCN3tK+nL
28xj/9P2t6mzRgEQSXQ8SUidwHw/AMV3wndkX6+dljAd6loLivDvtPm4lAzCTZMF
bDXARF3EREKfcYcXIUhSA4FZdRiKLyU4DptEum05KOmzi7k4YyGAkqv2/Eay9agt
X8d1ty5IRnuMWho3GlKAAsEhA5NiuDX0CW88f78qywffGQQMs3+O8nAuIH5ZbFNo
RgFsuXsG9v4VYlOLdjQronY0oweIDAM1Iv52QDnTF35aiswFiGqd580hjaVlYQUB
Zfn+m2ByoigigU0bzXWfHwYqIKv9G/tGodfvhqVM7sxaikzAgNKt2mvoNcv10GwP
G7e5CbdsKJmATHaEPKUCthyg631OaZAP8sPrtEA43cXtB9eiJn4QwVoQ1rKEzxFo
5wljMjWGSghskhy44Nv/svhD3fJmjb5eTNxEn2BfCIald/J/T8WyYmogu8xhuWpw
npObwMqsNV+5U6ncoCbC8NyX7hzRHcsu6nMH2CSiRqBQ5FbWsU05ukG8YPLJiTCx
oMgXYbYKZas14qpDZaFxDkqWOatBs3lpxbCD73d970E1b4LFHtlJ09JfFFvg1Dho
L9YueyxI1bnhFxCBy0s8gN3vhk0MXUAn6MDAfvHCLfA8H05gqkoGw1yEDbDScZIo
Plz+E4OU8Yvtks9kMYlCcyTVZTOcWWdG+owCgiw5oPg7gZX/WWNWTuB0TypDFl+C
XALQvApiza1Eev5VBANWqOxGkju4GMtPxkgNPsm0PZD5T7rrnfDH11kKN/YRWYYY
oYB4Pc7a7KEVvoY0VmqMcGqf/05jWrxsTQ4MHKXMw21i5SHo+egM6Daq14aIxUMR
RqZU2mlS/KmPSIldJQ9y/b6maH6JxkxQEJm1QTZb7ZLwmN02fD6cMCG+eAePCfgo
UT1gHauITJEiHo8li6Lt/0pkoHs0VaXtrYmo/c5RznQ66xH2epye9iyW0n3cScu9
tUYlwKS/4rRrFyQDCisngosqy6RVBx296DoNazzrxcBOr26UrEV+eCo1R+xYumzT
wNmXrFrSr7zI+Am+ZRCs+7wXo/hxWZB3mReJxR/gIwgfuQshgIDHEebH783iwjkn
LtOHnqWicWWJdjdXwZzm2Wq2bRhRFgldjdgRx/zkl0J67WLx2Ywu64Q/Ocizi6CZ
VBrf5cDJ7miqcGwdgV0FAcnqtmuz64Hau4f7WuLhq7tgcQIvls5SDfJiqAkTkdmn
uBOrH6F7KC5ZpxwEMlFU3a2q6r+8pPxtH9gZsMpRjG2zU3xVOLGPcDcHV3alPhm4
u8ZbW7GWoa2mjqd7pp7zfYPkuMG+iCgPjmOzhw5RVpZ31z5Z8DQJy7n5Pr+K8cLE
BtUe4uY4mK0HvyB1YAkJoOMLWRutDz0LzuvIpKWtN+xTQRLxOlMp1hHw1YkDenrS
twD54QshqbMQMwPUq+7MMjc3Y/zb9qDFpOaj0FYhnkQzqRTFd3p0kMY18zFsRR/C
gZW62u6kxVXeaDBeEkS/lOo6usRB1dtTI/qfeFYI/dqd4hBTnUeBkUzXdUEuwkIn
c8nwiXafgMwdlZrXxR9xv+FTQBuHPLQ7a/xLbXIjZoREDMn24s+KhasbKso7iGIe
0wKRacPpDIh7Z9hsI3QPa/2pCNJOfMKpGZvnGEBW+bIin3QGRa5kFwg+FCoLSCak
F73+L/k1f53ps9lsW6JaBTsl8wGJ+zdmaWsaDUD7CmJtgZ/tfPHrNPikzn2s2K20
ONNh8iLsCBNGKCcsuNjT5wMF7s4uUdJ/wf6hvGZX4R9MCOn/19GTv8CFro3WktSV
YRWOJPzZV3kQTqn6cvDhvPXVO+7UP9Q+XxHiidJxLR9mx+eRxw5KTq/riinKvvFa
HqAvtJZlSq1cF03zRNonXoxg/2xa6YZmOSHyM7/6lWrB0tyRvxTArBKgAFvaVB6z
OKVHrpiuWz8ViULOs/KyA8GJUl+u+Q1tZmTNb1plai5pt5cbXNuoURc4zvBAjRzb
sPzi2LpxVICjdDY2zTkwiVFURMeQ5jIUl/svmmU2MoPBNJKlIiSkgBwkcj2efHn2
AwGUtTVA5ykKSDgAL6s6/FjSt4KIBF6sZNbZN3RINmrIW1aBHMiEdiGRWoMjr19E
HwqfRJifrnA5rKkGDdTB4X1M/CNWTzOg0r6PiJNlX9+rYkFfeL8+JN3Q5AZSOQ84
eQBpP0UtAvVzRIKxVjn1yx+7+sjeZDuDr7EBQL3GXxFtqyK8E59ZFOtQ45Lb+bqb
TT/vw9gpqJhq8Ow8rU7QAADKQ6kWd3dIvlFx0XYuxOt56qExWX18W7bb91Z8nyac
0VSAGBhECmv3BgTR+iDXmAQ20FEzF47zk9LW4lVeItjWY22vKyD6oSapA8yULvtQ
4spFlusXIoe4GLZ7ZMcAtI7eufVYo5v0/zil4wpZhf6PWwrL/fWgAaSXuP07m/zg
/J3qDI83Z9IKk4Yk2jkTDxZShQ75m86Snsh0lKr+usY98COgScUxo4w3qLU232JV
tg6U5ZlNMQz2leE1E//ypF7mlJYN4NLMgZbCtkVih8hPgKLa7ovCljOAk4WeijEl
wWiAh3C1l3wBrGNJDqmbvo8/3Zw3Q/yHPzzBTRBfyIacdPp/GK4RuppFdysZj+WH
j+WkNCZ+18/bUC6Dfnq4kNf2x5YcX6jm5VJGNQYOizbOs1enSGGhA/wcdaVxV/aH
Qyy3RlmmnzW5JHImEk2Ak1l3SJwu08aBhvSYIvdof+lQfo8GUKWD0WDLQGhkaZUp
VM7qDkJ/hl4KKT5yJvfIz6ileOG4ileDi3/dWy/Oxip6CT9Rk32NlzkLq02tj0Q2
DSJVzH2eNZfsu/QSNHyxZdv96RulJgxHdzIAf6AVsaUjD6+Ft37q5w+W0eVjskYX
WJGnSEm5b4FD1rMq8bZ8YTs3SMp9tZamVvK3lX1Z2vKfUGHqH1D8Xy2PcSpM+wQe
vwBMznUPUn/e8NsuVjXHeVYHEQnbTXAGGUDAFZWHzZmuLG4uYGXiQlsIeRLDJzKz
3fb8HAIsNCUWYpHC7KqQ1D2rXzBJNj+NKCP8QTsT4pVu1zcVRSsmgkHynrZt3FBf
vj5VoyhBXqRiC0cYcXMGhLYysRIXGmcDD1NEEDMlynLf69qIH43uJf7AF9iHVRgE
/SY57DdxgoGKGFZ7c/PBa2m3Q4LDotVfm50ZxlJ4E/eEvPJry0JyqlCMADSf1jLm
QLeOSUGYJPK3AImzYSlrsgZiTpWKjsVvpmmEL0pv2qCOunSf3XIzdoY25cgoeBse
p3IVIu/OA054sXZ1MffheOPgU6wAZRIXk/xp3ewXEvCJ/EQKdf4M0mtbeQOZMv7f
IgAOjpDHSZKdAEpKnIsYiQ9hzueolNFKk2c+fAE5G1aZXZRUaWWSzO5RUF5ze0vR
EaFr50HYgAx7az0xa+PNOsaVFe9N4bOTqeg/qraw+66NQXJiLacnKWFLOh4Y/C+h
9EL4LjnJWlPT8XoZUEMOJiSsuG1UPQ6a9pDb6yjb9smEZY+hC7VvR6LUaysOn6F4
Ym0c1L4XBEIcvNDWk9ncAqbmS2XXjdjmaqyrleHtTiJ/CvzSVf8gVHVV+DMI12RC
zVVsvivLY/pWGBUxJ1cTvRZJMUmK0YshAHZ+qHMOdGnYY43cUlMnj5Y80gbjAA5n
t6ivmbP1LhyQVTksHHsIn/QtsvhcVPjr7cBO66eE3hG3C+Kak1GzXQinwvZjqpx3
G/rJN9miqSgHTv1gG/Ma7ui+uNtj+4+8rAq0ztjUFNf86ZeWQvPrv1UYFgfyRWee
OYSjCfG1ekPVV6g/BvmcvgtkXOzKPrach2JL2wMZ0M7bXk68oM+Ygp5HWrOhwAYx
Sc13x9Tkl+u3cr6cm5K8eHpbLRu8oOhqPzF75hgDCmNnnE1drp7kOIOsS1V0TYon
esNeUxpUMIvayWIVI0yREOPQKBM/qvbtO2eet3ymauoQDUR7sIhiOSy9BD81RYRe
MksrgNHWD6uUgLy4nx6rjIwA8bEHDerUMriAgfe6Rr9NnchdiJFsS21Hh40FCyx8
YHN4u685zbQM9e/RtkJ5Nvn0kccZvkxHvqnm7LiekVZ7J5GmtpHQSozztr9xnhy4
IfVQ/CIkpvQL1yBaRmOWQL9Kxc49r0o7NNGHZkST8qfAxXO0AsDTy7J51leHrqVn
q9Ac70t0he6SfbajK+n/poNl1A5Fepi5upvuzPQbneC/lx8Wnhepx1XqKQzbzOox
Pi3nKjCvmjtTbV4LNxIBenYZ+DsH3e9Wx8FsoVAh2ZyQRqraTv1yB3Z18paKtIjQ
axytTO2GL6m+JmcnAxCO8h0Hqa3lW6LaySJsCYhvlatsOpTkxN3y3ZGMm/O593hz
VVudlhg7+y0iJE+2BvUKvxqo2+ChpyLDc93vG4cA/0AsmTonFCgqrynALhSSzk+R
OIlUhIFbVHWGKKypORS3HAQhAWPrlV9nDF486T2cVLcCV4v/Li/H3EMtbpMIusqO
dRvJz6dSY2nka68z1Z1o9ZtVMuyF7DgWmXiLhmptB6UG3o0Cmk1svme0+l9t9QLx
tfVW7E10J37n7uD5FBHMiJe3rWLdcKnWaFjnC16JLUa4B6+IqQCxSg1UchkOhi2K
31QGTESiS9SxCCkS2HVjH67Wu2ANbz2B0rZ6kmIPcy520IqyUsRxJ8Ax2ANvfUTQ
lhp+d9tstYjiHpUudgwrf31KENCpBikizbHG13dyWDEj1hpsZa+qQQ4d6AFD6uia
gpcZx8YzcXVlFMxgmrVZ4a77E8AckJwTFAmwxdPOWiTBxhzRrU6eyhlPRrHP0vVa
JiZFoa2TsoGKHHl6rKhDgunMvVd+PWXxGj0e6aXGe5dfTulE7PVAB1VMhJgwEC4R
ooGvIjq8gAFJANeB5gOItGEzKG5N5sojQh15sJ5RPrI3ubRYZWPU2NpjcxPnsOZh
caPtYH4QC2Jmh4VMZe5JSub/WJKN97iGJ5HSqkmq8/sXgskKZZ7Iyg879fHcHfuy
OKp7tmQAQrJrs70P+UKO5CISVz1lKmM+Byr5m+NgJnTwQBeEgORYMgJcWqu+kdu/
m/O/f32GC6evSjoIBuZmWgTWVG5j4GRCCnrzsNJ9VvZay+5A5cPBj0bzu0t7dYbl
sjNI88HLb7j1eeHU1rldy0vViRYrQ3GSiUgTL1Nt3cI25Df336egtZV314VPBMyK
+83sDYNNA+A2NWcvHNM/BhEhvBm88qo3s2k+ajmdkjLNMiJk81qIw2LngbjiRDS4
qRLDKP6e/tfLZzf6rn48Yw1GJYpxW7pX4u/eaCVevcgmBFtsJxCuFWQ9EWMnO3YP
QOypDmBK5O8vxPGmUUiAG1MckMrdzA7L6F9E+LTY9AGH8HaLWWWx49b2E+KQDmR5
RkUstq+63AHPL/qJzea1SFhZDxc2zZuznO9YvOddlE873FvSu/PZiwDSvwvMWg09
/P5Iof5vKIG3TvbXDhZnguziKcMQdYiF5heYbAsXYIh9qWqKeg2PxWgCp65Pz76J
k89T4s16107R4lFyKgQsBlBpCooZ6AaHS+tTcaj+FAPPDi9sF2F4G3s6kiXwuhl8
8Y0dNSqKMTGs2437xeZrHOVXcrG5k+wTvNVy81ZjSJQpNrlcqXZLmk21o6wvDcqZ
cS+ycFz4NiJ/2qzCOmO8BvqNQxjmX8vsVYxvuZ9Zv7uhZxIZ8zM5d1gW6vrUl2Ms
HuA/aB3gzmZuoX+nFd2aYa2oMEsMc5ghBRpjYkIxc45LD4tSHOokL19Ydu3xWkha
DK80RHt0kGbWGfEjSRNmY4a2+yI3i1a1tEvKWzQCo36y1vtg2AWXZv458WwEzIjy
gpeDU8fgZrK46+wZr2M/i0VDdpcKNWhgErBX9K/dZet5LfYj/t+PaQr61xNjMmp+
VIEs5aKf2b/SRSw4UmU15ZSHsE+adUvXccC5xIstRjA4YW0dnM7lUl895aZ8CP9V
bCXhscwrSSkJuDF7+aip4isf2uCpCExE82tcgebZHT6ZWdD6OBo/ncqte4Y0Ey7F
jeKuZaWuQYrAP7R9YYHsC+uWFUKCOXVDDh4Fg08mgJhiz/c3lG5qRICPy1+2gyD7
cvjE17EJInYVw8GV462W88rT51I2+odUld+HrgGraoszehw1LUp1m2mKIDpFvO2S
o1RkTf5alAA3ufYtFASnXTtEreasIGhLriYbhuSUfyfeQUgyZlXqCebS2q+bPgJz
Uiq9mp9kjaiRjA2VTK6r+71dTBhUu3smmFWJDjGx3BLUwxWYRstnsnv2wf6puISH
Zr3j3+cKvLl/93T3JQKG25453VZYGOjIotUm80Q1HER6Nflx9kfRzGt3VTGfYKJq
YpOy3Jc0UcP/ltCMMRUQQumLh3MIDJj+XnTiTfSl4JOJa4F8GzcaoKLWd4/RRBsy
wAJMHBh/JNhmkoX3eILN8p9pjX9ZTeYOtKGZ2lfA90H8D9Dxl5NgaN/IcuIKNGFp
S9Mofa2zOJwHtnzuu76/K85llsRoN0Hbx/aYq61FRBeh6BM4tegGW7ftgEqlBCFy
YSFM7E/Ryn91syGM59DzBLX1o5/h3Awupu3C3Upnwa5lC11f6Z8aiKJ21rfe1Tzx
QV6tFbWr16r09Tls0ZPjDDKs0rOVWG4l/AiUwM96hzDIvP8oaj25g5aadfODk+dg
2u1UZLeHp+6tRJfjJGgDfnm5I4b9t5ecPkKTTUj3nMo49MiRxNcVESwsCGDrC+3Z
y9s6ufQviLHa4jdQSz9OvvFrhBhhImVfI3wnmqQhto/GlnouC3WwWbI/Ycj80VT+
73yatJ5+dQ4L99ZYf8vv0fBX2E5BQGLPCF4QYh9AqhBGG8ynAbcKjzWzFj0EzCME
LB3NIxpoKHrSRYbPR5++WndVy1O4+DZbPtqWqd5SKByElDM+DKiPzqkx17wp4ErM
cCsYuleW7Hb/foopBfBjI+BoqTsTnd/VuRWxYMK9HzGO+nlsBQca7DDqgeMqwle1
DBCdVsENgmjfbvTn6umo5yEuGrB7UnQDoMgA6AufSM1M/1Azm5raRqG0ux7NDlLe
T+LCAbHAO6ummJGZ+4yUMqFAUAZYFBhOVvefNITd0DJjpZG76tdZaLK5h1kdKghA
27N/oBdnsIuoVAUmnEzIMs/aaU3P0hbMxY7hoLOUrOEOWZv4poJClGATrna5WD/8
/X0USpO40t7jnqm2Tm3h0GyOGLVlUS9jgXqkfAsfmlJfvQFgKnm4oeTuPt1E8oqC
uVkuqgT+v2iUby9vvfWYZc/uBvL7kIUgMgnxsQQ0mHTGoOzKPFP2pMAWanoMqzY5
yI4K+ipd2+uSh6ZUAMb+g6FsFwkprshOjhZlSGRfz6zxf6u6tiwgyCn/Ydgiy5++
gv99AxOzwzwXd08KqhzQp4SWIreZl75+4L/bnqeif6Z4fHHJ3tYz8oytkGuCRPaS
HOMpjs3aGp2SeCYj1wtauMSCZj30kSzKRNAonvP+The2VSk5cCdGl52lG6EerK4M
TQT4PZFqhYPv/OoxKIC1AxHp2AGbzUHwqJMa9Gaa7iNxUYaaLL+udKU1EWCuNqOz
5PQ43PFI0GoX+PzbbcTMKn0vNYfAVITWp6AdaapVVZnNO+A2CrqRP81y322eqOdJ
p+4AFt5nUT/uXPsJF/wUwfXNgUauUmWRQPTIIspkVkeJU2kT3C/VwGlpG8j93G5E
jmZeR5RJlQny0ap3nZ8Ud0FrPQwXZzrYoqZl4JqgXqSQ1oXTAk8neqaWENwQLD75
UiWghRI23B9FR4h50vTBUr9i5I/8PduoHYciSd00DhoYmWEuJL29u7cfLx9yyp6v
Y0rpEyQ4I1LpAna5m9//aH3g8DzoIwd5IuLMmxABZE560MCFr/SNz1YafN5FUR1F
FuMXxI5xLseeS2jByYdYUI6F8EP9YXCpRFKVNocJgJqhsftGHSZzfdUuuOhbTNy0
ZBcamZzrLD2RdWejdN0fAtshGpwMZogOlXiOahkkAZbIIch5PpfpUUy089D6BkEe
3Ww85ONmKLgGrtmvt6n4AghrqtTlPpUiIz84CciuWNxKoRBNLn9TXCxvg9i+lceB
xTG/c/+MziEeZBWtI8tlmlGwP3IX/NxBi0trB9aDMSWnUmNHoNfFcfkEbebRdD7N
NGbDlhgEVQQlJ7cXTuVgRby1a/Y8DCzIsYKigWBmDnCiyOkulsdsqbtzq++f7u3n
XR/q039Ie0oBriJTPmNWw20S8wYP+C56Oosk8lBM0ap2y76Ja1H6sy1qcEiH41j6
wDZkR7tE8KCZjBT4gttw4g3+v1ScOOXzbkpaVvZ/bKIsQoE0wk/04mwidCwgol2F
4IA0I2fjMoYmnrkHReBIbiu/YARgnoTfDSNSZY+uFO9NM3EwuHKVtFfoSXOm5CGw
Bu7zwH0rQwGgMkPj78PdmqVehrJt3F0m0NyhSUlZUkiQCGNANrMIKAIyRjMvfHfM
/eRmqOA0C80yYvrc3TaXHrBZAkZeEz0Qx+WPQHgFjtoR9AD5a5EaHK1wv72F9NEy
nFivZxcXxCrOaVdJU0m0kp/C+XB5QFH3OHNoohg+hARpaVeyQjpMYoJxknMzvHg6
Yoj/MgTZQKkCTrwgMScdMEWIAbC6VjeVei05pPBP1LA8dNDq0Ubetf02Mhihp+J7
C452hl6bvmcbhA/YPGc3PN848VdKm6AdJeVMV2NckK+6C3B7NufQfGx4mpgmolVV
Th+mDq1IDr04VNVVf0QO5CjXHL0WgOsYQAHxeV7FUuFH5n2QBHBFFa5XuLJktIX2
BirgP6THewhrlFN0jX0LTfmdxTYbuhxD3tIOcD556t2EdspGPQvUs2216dwSIacq
COL3WM6MpTZatrYu06h7Y8Q8b19PGtcq4S9Jo5DBi4/vVWmeUEQUbjdxonFdupiz
uX20if9UFrco+rZNgJbal857pb5frZFxEO5QnwtZOb0x1eMMOiHHMwEXRTby3cdD
jpRt1qNM/wAtE69Uj2p8HozetuMcmwgrEdwduuRdBZ4JZbMsS4R4JFg2OdjAlwzi
mgYTdHc4Cv7O/POnRD9AZ+oZRpBQalB/tYFrtspNi33CwCkhgxKIYtPjS70bxlrp
fcExbAR9BN89L+zlGy46B6uTlArn+/KL8yDS742QTlcHyvfI4lDaj+YyecK9Ndq6
eEUrjnU2sM5F6nVH/v6InEEq2RbS4sjSJPV4ieJ+TbtRCXsZbq8N4mf0S69O8Syz
5bweLIXSlBjBRcU66sgiqIT6oXblYgEkkTXkcy66tDspFnELfaq8JhEKuUlXSEiu
/LagG5Zo+EshSk1SJhy7uJ4wea184rHClO5QDYIIS7Vp1HxQjFDEGAiMtQvTGjTq
kscojkuQiYO63+hnFaLIHaisod8oA+xO/T4L2fAbkjWs4tgDbgs/5bWVd4SKtMUq
EFmKKAYggG1vTDJ648l95mqPm4dkGQ3Ac5fWTFaNcwo5Hlo9CP77amzgW6cp5SMZ
w/CvTFBE1eLWY9ZTFgyOhqz0TvrxA37gnrUMQrC6LIi2LIXfyqvw2zHoW1yLCDvf
3ATiwS0xO3jFhJOCmqbM1oMuhKmeKGFPneo698l6mk7azSWLapnlf+nvuuEy3jvA
0GMz2mUruGA13xHQzxHVGm4h1v+ctC0L8yx/unkrC05MFhgmK0wFLzeFyPn/HdUo
cPw+TIFaWomzAGY4Ofx3/blZCclTRfpqqnBAHSSF+It2La8EGtjMmyljhPO1PveH
FMUOd/RnBHhLrfV0fUvZdJU+nfbCvhsXxV2kuruY/KwJHpIsKPIASzW6UuqH86et
vu4sleZdO+FfsBbq6gTxfEHxsbvMCRKFEJ+2fU9LELrTxP+9otXFP1dPCkrOHXef
2RO7ztGwW+wLwNigWqnq15JiSr2SGIIM4eQZMm1iIvItv8iY/Kn8N5ZpaHC6gmmA
jnOks+fC/NYSae2JNblW7gmlLpm8X2pG1m1tMtMKSOAAWOPeR+WqQkOMvoCNQ65A
UGxzhoL+j7YVKaV7kWJGJy2kaurO9o2qK3JpDpIohfi+S/LMqrEGN5gRhCI7tLSU
72ioKUevxUIpdsbSkE8aUEdZX25pJxosRj+Vp4AwrudkgVzjFAuq/w+J8Rxdx2/T
IRsqKGDbyO03KzOjGl6rGJeDo3vWJI8ZT5TEWGx4RRETh7mypzfDnu6uA+Ydj+Oo
OwCzXafDrmYVEBvFEncfdlVJwnoSqycj3GN4hefQ/SYf9jKnIiRcjnh4xE92CeMh
dsYn9XHuef6tICMy2PHRv5ppGtc0dD7mAoYUOrvZZ7NnLqYFho/ZW2R9xHW/faVF
4HRGVBWJrq6k4yrojvs8sEtqktDXEyg+49aO4+2J6dXZI6sksaWejhXWRWEPH5ER
Qv/FI4vnx7b6Br3x7TwVbnyZM4pBStqSyyfuIdknp3KctHEt8fuX79KheFmnwbiJ
sr4P/ibET7MQ0zt5HZ44mKOEkbUVXUq2p4E5KqtFpxtMIQDeuqFzoNo5QGGjtTPt
TmomPOeCvKuYe4wGJi3cHJvLv0W2Ol8bSRl4vbzqjRvNNOB29lItNjrajTVlQjpO
9I2krtsjfry+foK7vUegn5Bmjmvak84r4nW6lFcG6kGIBpi6Rm7TwZWDMkcJO9Jj
YXEdNRtyHwPj5opkxFJkd+cjYpT8R+fEkdPIg8Ulh4yx0bVi03qWpJplYjgT8kr6
CHmNLZWWjyMW95Owdd7xSuDJf+RrBy9aD3U3lpxzPqUIS+hzz7YJ4JQGk2stddU0
BbTBomT12uoj8yl9E8jQeglTVzWpMiMTDVO3xeOE4GSpOc/7CQp0Y0R/Ol9QSrm2
lq17zTuBwzRNvvfa4fiHPlvh8IBkhgxbED3TcaokcPe1wDktw9oulf82oyxDc1z3
Kl2+dAggIn4pv8TCyNAkYM7e3eleheH/klzKeELtBjRyP12MrBzG7AXch+91Cltv
qAO9tvTpFd4D9TUPRET/0TUjEncoYhF2IcwexFGaGHgHi2qwfeVU8CXZT7GNnAtg
m5Lzm0T9UMkkf/sBX2WuXay0ypvSAUxz9Oi/71MErNtRAXn/94y4LIGWqVvy+xvl
C04sga0NFeYxgueAtJX+WgUiZXnvKRN87e8IBJ13bXoUZb75ntZllDwh1H7DlAi3
zAMG/sx6cOb5Y0D7eL/0i0r/BBNBWxfMggzaqCaWDAXqDkPfC83LCeTUMnw6ltlw
kS/FReqtaeSnfWxZcJQEYkse95WBfw23IowwXQ5tJjFGDHWNhexw6zwh+aCSTCp9
AOKWqyx8Vz7cpl5mfhDaOVobTFKdZXEwjwaN+6Kj3kG1idnRNgQ6tHkEFu5jv8jS
A71dcU17knX24MViLcDzjJnPoqVMoysdXJqU5BxB08Km57d+x7lVaWSlQmLMLAPK
5lXzFdAp0QJnWoRupekw/ZnIPyCpdrcwO+AQoXmJLz3U4NFSitMD6h2WoWs6FStS
78q1fY+YhqqujlsNUdSaZuL/ip6+Xh871xnYLB07QHTwp4tBPuggysmzS3JiThHK
CsrE52Ww5XY6+nam4FNwP0jLGtCoXQqoh7nCf7oq+4Lau6t/1MSut6HOLrZCQ8Ai
ahg1VIhvWVMGyn3MQhXv+mrL31/vaj8n8UoyqzUxDdGGd2Ajco8Nj88lXoWL+mb0
Qjr4UGsvhYyJA0+VhzPy+2wQQ6lrxOIw7/d1jJp4Yb1h30YmKrwKMairECvK92gm
LGIml/6tkYWSdFfjVQ/fas1OLxZEsXTgl+iK3sBB3k9vzsf5Cg3vx6iQrD0+4foT
bWf/VjDENX+S1Kwq4P9RwIc3/4mOoDm+mMwkxcykHDBA6VZevFB4adkB5z1QZDYU
ljNCPA7Vv2LFJ4S60MtMc6oKcuF0tH5H2tMzFQpBvEzB9KeQGlOfBY1XoNkyU4Mc
ft+wSfJ+ZRyo+6axGuaOO2dTBuu/aCtlynzWe464p0s4qNGsNaO1yByZUxvdrl53
5ga84Fpc6wOMJoI5ePqvhpaV0IxRRW55gnPrIWLDWIaouSomdidXmH2N30bUinc+
PmA2B6vcPJ9LYQn4w5pUhUNUmp5E9I5O/nUWI7UxLlW4OX13LiEYSlb9CPdE8uMC
5enH80eRkDBjobrQlNY7U5Zvr3jv/twACYg8i5FqtW0fFT9AQEcwPofjtqhZlHtM
VaEubqB/XU51Kz6JGSe9G/Dr+5gKoM1Kkk4KNu5JMNAiOmBJOS1Oq7tdRaD9hRJc
2TNsGP0GikRRQYhRdavXh+6dzeCF8ZeC9GkigJ691Xis0eo7/093dCpO9GMINS0a
2iPU62wlYkNQrFC8QU9YbO4GQNsq2zNVWpn4Hr7ogS6EuAopdT2+GFIeJIPXbIEj
Fn3EMGXdaclfnR20EDFM1fidF0Xy7xqu4nEdFJjTcBHh/NjgGHTMGCL5sH+UBTUL
Fn/x0/1Qv4DRscrJB9aAzs0EN2gGovoXp6beGbHX/kbY9S6pzaVMremn16ONksqr
NW+u4kDLZxhpNUNpeDs3DtTgZEILrwK7tHvQ+YFBv07QaqzPs4/IOtN0a7/3SzG+
p695oxeB4kYMf4LV9xYNi0uY2e21vrXYmjvu0HL62mYTPZgbaoq0DVN5Jv29E5mO
shiB9kHJWbis59p0cCQeYLvRugwz6d0QoJ0ueHgXnzITg9e1pQPoRKlkqqhWyyPa
Y7EctHTGugUPV3Sgf5rHYHLoiPae1PHWcSVyi3AMXoO2Hc/Qh6q80F4ST0tu518L
moylJWmYMgp44NLONeDDFQOMOo18VakMDF1Yrl1bQAZe9cZoy+4lXEa4SjVdDo74
5ytvwN5jJtAdjWD37CKbSFYb3z7OOJVwU2SyAR5XuUHRnCqQUVsB1iCx4MriVIaf
hdpa0Ry7H3g2Keajvrw4sHpXn1to6QiWmmNlOqHZ4muP9xJynlx+qg7kKiKnKWB4
ebUpRS6asL9mfzpiDbUoM+ypjouPMTucFnVAeaOf3Lds3RzWxK+IG+II4aSP7kQp
K3BQIJx46mFkBUEd407mUxZZ/VKPrSSVx7D7AzkEv1nv+lVoQw8z1vo+85eCEQqI
9lXG4PGuiJELvgNbHNpaTt7ShWL+45CTUGvMOYZFbLaL5vfALiBMcDrTBoJbtJV1
TApIghMvlo0lDHMu65oheToYmaxSDBNVetAVcdD52P6fgbKaI0+sT/qhNwVmxVQW
2ZH8+NpFyhl6tX6nRkrkDBkSTZSezwGtH2X4nJe0PCLkEiuxM+Ei76bj3zVDT5N+
ewQ0SbrJXx89vmYLa5i37MYVfu2qSzYww+gQIMnf9IcYntMGGeNd+hv6y0svmv2/
14+qKWK4L6gDYdnQIj/nTBLeq4QBURTvJ1AJxmqLuIkKE6AHu8Hj+KZlL6R0wB4s
t0aqk2jdyCldJsL/ow94Se0Ru1s8mvRecW7s+ArrbCXS6QfXALZpGg6VrAWeWzIW
cGrvvwxy8ojcQhpvDw2AviiAIo3Pj1jW+r+yf0DoVMvaaD7nt04h6Rb5prEktZhc
+TQbt23LTLRjXmmXFAv+fcZQHUhlgm9neFNCTNTpu94eovaoy61IY1EihvorjnJ0
FuYcOE9JyvhoMYvXmf/WRWjiB6TdDyX6hX2wskyhCcPyNworGc4h7Pktb/V+Aau3
B4MNoMg1ifttzhr/KZ3uO/bt9iqtj5w7OCwRAWw2o50z71G37D1EjfE9tjdVuHB4
7+G8h5BML0f7JVqi7k1X4KenP35pEKLEJsBxT6MNp+wrzuEvYnxAy/SO0LnXKGLY
/Cua6720pxqedHOmaRAsizDjVrr46RR15EVJiJKmdUo1YVSDpkrNc8Po1Wpfp9KU
d6yCe1+uwiPWc5XyqDH2LAbTxh2TJaqtNq1j4fzCliOW6j9AD6+JnB6JYYvMl3VA
ivkHAYdQpCVM9MrZh/r6gquN+M5mLxAga/pwrjvZB4ydqLrl8EMCOxSRUE3EHTOq
eWdHM23wa+CE8qXWAcB/XQGPNrgvBwQrDo3Mb8+5h8qm+MU3xS8+p4r0tJKNHGtT
7o40EL7GkeA2Yp8Htk30KDBGzzeJZfmqBdd/VDjUWabc4qmC9u4RKNwSlc/l5W79
FIOgfe+h/1u2cCwjVG+Kvy3TGKYWBamvRDdnVF1j6lHLiuPTlkzwmbpktG5aYLZV
kPpenR9HriaV0FwPfo493MebVgBM95z44NRp1p5EhtvwI0TbkAV44Q+EBaTQ/R2P
caFsdN93Xs1FWxAbfGl42rLPkhYWg06DumguTJbi76okO9LEh7w3TQfIqZMKHIS6
mviXuFPswkPym5l3aqTDwg1Xmvc9Mkm64SylVZ3vsfAin4OOG01b8eiwMu43OsFU
gF8fJ3oJeK+bl7f85ed0BYwtxdzi8dEDAMCNHh3jhXYLdPQ0l0NG6Mr9xdfoDA12
kkxTDeZsS26SmoDHcCNYqKrpHRFq0RfcrO8gbAZ+BH805OtmARi0fgbKz19zwueW
cyvIBeEa/am3SGk8wWN3T3lr/8gvkrNGOiQIQkZ16yhJ0t1tw5P/fhk9RMQpiSME
zjPCf5XSvT9pw0cBpL8s8Bo8X4MSBCCqUDinL+ddYhtq7YvVOFJKJyER/GA7NpkN
3+1JXVt3/6ek52JE3/5mYmVVedWqaiuYsQGe3ijZRMfPJlsHHczo0BjsR6KMqAa2
BytHOOpLUeLLd6Tmxnqmmr4zzcaYsNu9jrijWaiMVZEclcenUCNGTgBxCKKagRxT
n1h87mqbLAK1B1naDUqYJN5dYhRZP4EK7MTuaneQob7512GnrAaC+VWk3oCKAHjH
VJDwI13biV/pukcfAwRzB2cgkIooifpmmFPOcPy45Cz2HvvZ1dq2h9lLvX1vG3qU
ruQiegIZAOTsreywmIOnxfK/SkkRuA/lxuhcMuZWqZnz1DOhEVpmAdmDpn8Cs1wb
Kg265aM+HZiEXQutAJ4mJBiFAGKup4KYbzXKZ4c1SpO7BXiDCd0XHVyDOikhNV7O
JNHtJjcPlgRLWyao+30ytN5wmaDj65dcefy0FNPiic9GyUYlWPv9j7diDzZch3Je
NubrefSW+g+N5XeLjhK/cfOR+57Y48EgAA8FhpLeaCFkKWGx2DeHp6TExy/cYi3M
GTik1rZNIlqxtLRI5zFrDYuGzan5r5yZXW/9rgUoi7zeGt+8/Hex5H2LLpMYKMjR
And3fqq8XPey87eT7sVl5ZaWaLpuTL7fY/azOC13UsMnBeReAtNZNzpeiWEZMaC9
YPwBxd7449WW9YhfGTZzO9qoZR5qZ58UT6972j1113b/fDHkX/DnIoBOv70X9M9S
DWpuNuJmLyzhpo1af+NUn0gXjUCXqd1dw5BiyQeQHDkhDhUjm8Of4yEw+nttTAzy
fnIdfBYlfWIwRx4N89q3MVrRiXitzyYksxTFsd6fx2a7FvLArU933Eaau07b46pj
QWUAZRj6zsVDo3Dju3qK8/qk+eWM2ZRzHSe7iad4ZNiCmmeCOHmNZtTxDMQ6x7FL
unEq3f+DLpCBmIIj81euqVsUnap4Dip2KIxVkhFSc4wJVdR4BuvP1SAodBnhz54U
3R7coOL3FmE9lX7wWvPMW8qSxBq7ZQck+fzYTYcV4U7kAm01LwznumuWBHEhKBV8
j+9sOr0JpdqjfueK81sQOGgpSw2YXpWoi1ezbkIUpm2sDqO8YrkM4XsUGuqWyyIZ
xd2zYI4vKLTelFBR9fPA3HWlpwBxCCoPRrcMNZNM+Zuuh1zg95ov/cfb0PyUA6jX
e1jw8/9Grw/ULXq6y8drFjcV3Q3AD8r2EDyR1I0SN8eBARoJh7QX4azUceDr6qux
dsD77UfEr5HNWfbSQ/536q1YAh4NW9sj4MwGaQ7ZesSv34gDssUjCzCrvHWyz1tx
dgWI9AKfJmT0juSDWwHqrhhkxRp/QDppre545VvOGHDWsScH6V8qEtn+IINlAkCf
Wb2P3uktV4SEtwLNdYdc3p26nq41MZAdICESeeUxeJWqDhEs//L4vSUlztCho77x
k+cvVcDeG4ZyWjQ8yuAjr/53RacX0EhlZ6GSs91nqpgCJYl6EcFf/wN1kIrgtLlB
WD2aFG+wT/zG51oPrz5nYI5ijqnFVjU7Jxvsfv55fh8bZD0weWAtu4yYlp8CaDXJ
hZZ0SATMLLBV16LmBRz5DXTDLSgnXissITRF5jujeyg/5vVGHWxAIOzLzb9VGAf7
EI8b+IebzajARWALhVcFoQI/JGo4AqnrHjx3kUJSIn0Wo/jqGXxCqryRbIa8XOf7
6XZtEpXJNNtuuJIKxPqOezxbVURBOas8tHfOicGN0os0u5pV6vYEkn9Ur9TlHMwU
yqfqrtrqbnbFRjYVOGJ32BPfhIbxbHcT8v6evPOwb4wwolDI4FikjM+gJi4DdAvg
G+SSdG5uT3wsFi8OMds/B/4mQPc6/5/vMv1IBgeFWefU7h/l24DfK2fwdk2I2CMB
FH+pIqC+DYpcW/NW8y6PzmvUwgNIJEoSYT2f29sHOexoNVFtEsUAr0OMbs39CYPz
w+MMcEEfBTlvyMxVDNid4NTQtGRKwzzCBYnLr6XcjPp9qiT0FXwnho6+i7mhylkc
YWj2zM40IwDYwwLukUMxtOW4HNgPCcKz+Eq8GauwBmlQsJm62d7zJdwcMmg4m6zc
McshUE+zAiKfd0yKQySjIj1golPCdhirZbHBMmCqnARWovqseNwEtBfYAcL7EZM9
+Ij90V1rGPwN0Rr6GZ7J0Fyhfy/ItwHF4jelwEQZFI3d30USyhRkotswajhArJk0
PbLVn1n22DJYeIffx/g8T0Ivt5t1z9ZvykQT9iNEuZN04adKn7KXK3C/O8HeKCz/
qFpo3+0F/lK51gHS2InULajmKBcOcCSy/b0DA8uA4VBfWZNonDXrkSdNfykPXkdn
6+PNY0XBaQgHqlFbxe+0iLVeEj86ysrdVZ/Hr/W6HR7ZC6OKri1jKsPDYBiA73cW
QvGybjpyg8Jebg1AifVnT2KPN+Xv1h1SuiU/Ii6HVw4NOOhtMH0zH+zDFm9PUngX
tCTqIGz5lW9D+7H4kbuYNZUqT6Oec3gPBkDQVZpoWTRWbax2rjWzWBoKC8KKgTAh
YbH2uS8JbyNPWIWciiHPyQvr7zvFQZcVmCSz/F4y9fdsY2GMgYAehZvOkGGIyBKk
mkckT9OhMul9CAafpCbXzEta9Du6F6sFJSiRI8e2onf/DN5nfmFB+Sw6T1QZe+YR
UqUUwRpEIRk0SwSCjsm7uUUZiVxxhVGlQiMwFVwcTuyKAEgqY9KvOg/pJgWNfdmu
Y6/IukAze8GVbpFY8Ut3mBF+liJO7b3CDkEI++uTqtQgssGGulVJtiR+D5CupLz9
AjWuH4tgI47jpviuxGCQ3HEcpGDpCDsnaJZWBjsW/P+YF4P78wk6T++1Trn4rSOH
lxY5BQjRzdj6/ScP767seaUrfILuwqUsYjkI7oPKipD5yJO+QjksUq7TXXz9h//x
cwV+7UDNquUyrnQzSEQsISJcL/ZTPtjsnwzTyWAJy0K6Atx20Fswel3oylUpvmrI
SnPUC20QO2e4JMEd21tz9MVaKsVM6JRHCNRmJqtQiecFoRjct1msa5k290yxlGsd
356YjyqUO3Pai4Ry5inH19oQ4nOaQiv9BtzhEMJKZWbDmp/R3+2Jkp3z4ulHPdVO
kqYVfQVZVOHEurxZ1L1eLSm2kbeNPF4ULUienqQDH3EBCLoka8Ykelr6Rj4aY8rf
TW0mTrraKZe4J4ZYHI4lY2D4o+6B+wUlQOyWE5rpBe2Asv4FKrv4gsoQFrbY7Ygv
reiT5J+aCWOcvsGHb4GHO5azX/AEkVTxCDzqFBR+2y6/xqlToggSEtADviFvpSkj
K7oJ1ZU3ru9Z21tbHPFhRXSSmoQracEb0VsCIWPcFe2NZDvWHBGgYXHf52eEZelU
SskW0rT1miWUg7mq1LRH0wTTDoFCeivnHOErGm2PDcoiFxXqawcSEWyHPdllMOCj
vujxfizIM//FpZ5uG9go+R7W+PWrYXfEYHA5dMnYCcvhSTHfHgB8C3WT2yG6JbRX
DVOmc5uQ+DEfg0Crdl4X8jsopCgwXYy64+D2be8Xs4MdC9TZm8HnbMK/du8c/OMb
SdsA9mhZIWwOWCkQT9bUP5eiohExAJtmLs1h/c0xBKZW3Co9GkDAxi9JqaZ5z+ZA
qeTdO/kdQWpEvTplPe4npUj1vmupIYoWwEhspsxnZO96asmvMD8qGT9hxnMiw4R+
VrQMZ//gIDwOHF6jZc4qpOJOcwHyBkZ+eL+LaWWYBmDyM+fiVyrcABB51H+LQL+u
KeqcJcUrveVrrp3t9Djt8diDgLCluMDlikI7gr0jjR+SO+WWawpptINZwsEGX3WJ
OOR6fujLwq1wlnPHXZ54EtZLIOs+13WDCntOHzeNmqZ4RC41xAOJWuO6UeMx/T+q
eRyKCyDCBAmKt4F+ExwAJWYhOULuzLhQwvMKBWIv4TPhA+a00+/YafxwGhnX0Ldw
WCTlGSPrTxB5Q3ieK5DYU2LW70+jzvrcZe72f/suJyfchKLiMuaBul9K/Exe6pxt
kQsB8MdSgqh7OzlhMRv+oi01qm0KL+hj5hwT9zDcvC2TsZtL59mybXYfVAOp9FR1
ZKRERc01AWVObwmPColAfiIWOleiXk42CP+i20PSmVfvHr3ZzEDQxGtsLHzVleaw
PxNCYUvfRCcnQRuI1SbpK0mY84gHxL0p6j2fbmtnsYTNyJ/+t9+d+rmtNf6zM9qA
jZ0aLHMijplkpRXRICLyytBL58+mUNP3X9I89eG3mtQVEVGVsN7TdErBTfa4QWRc
UFq2vSq2gnFugIAzzqdJx7PleX7cKnc3pdapBeJOwNvLGzEOy0EMx753vjbT9Ibv
TO/dl8bIOMdYgNVnGLndMk/BDM8q4wwOlTuNCKTJosStNHbCHnB/1kgoKqZL6lMS
ujoIpdB1TX4rgLmqQyOUlC8wc4nkLlCzHsV+X96AiDH5/vDkFhTx9Il3Bkrku11a
1dBeMhffPdR3Pz3omJyEkH7W/7QfFdpqIUxhjFBjL3bjWBaeQMe8/I03lEgUJBZj
79Bnb8QZHOG2IwEKFKvwOV/r88rdsv27xSyncVRWRBBCMWQGDXEGIeYTpd6Z1GrQ
51NfFZ4OAShm4tdv1x//K+U/LUX+s9x5wvJNfbdACy1/zsXSC48bhOiG+btgPsSI
PVgVxUf8iOxhxB+q4fhKUxCfgmGkJtmDKs09QoAD2GpekXCx+1GEaqh5k3QDTGYB
lFFeDx1Fl7XnUrhmOQNZ5iGa2jgYFnDB++DKvpiGHrZnHc7NjG7FaY17azJXh43d
UehbEFX9mgjiaV3f2DNDRV/SIeJ3BUNFHvjho8lKh8qPaGwMdZv5kj4sxLj2YgSJ
V+Yl0Z3saEf2GYtlN2YL132K9L/ljcTfBQwdwjJu6PtqVMexIrLGUtSs0aieOU/j
4/93NWzANMzCEkAG5SgzpvadondzRPlweettCCS+6aY/H6VEKT4/+fhNESCwAfhT
ecuKuyEMVtyVRiSseyJog+aR+R4OEsrxDg+nHsC4BzxSvt8RjA3JNUa2CwZy8gXi
wXmlz7h7C/XT7cec52dlKDyjpp3ZxaIZ4YekkRzptMBVXzvbh7aGDomShO/fMS99
zjRwxJXBBu3gHfd4STG03wxBR9vLtFnOHMoj2FH/8Q4bjuYEb6OjJxQOTPJLoatX
tj9ZbX03EiPRt6vsn28V2Tbzan78D6LEMYcg0fRUVfRM1ttZZ/kYlUuEqTyt4EkD
M9iASJ7UDrDPwMNz4oQRg1Y5uNzy2oJN/n1G/WpjLobMduG1697BXCR/iaEctWKx
DgR74ITDjfAN8S2ooR9on9bmHRToeFJ8q/Xeca3Arpabz1Ccz5mK3mA34F6mDcUy
pc7voB0KL1AzGDlWnDlMv0G2fcXXCLDwazchRTnibrRqdXFf336fFgFgo9XiRW4s
ff2m/kgWdpCmkQrgz/40NdX4Ab2WvCwtAWQ6vM5n70fKz5iV+VDlxT21SrkYht29
6YA+NjdafFQWhRVWyBDd6I8KYxoJldOV2yKCjynhLEpEonR87iBCzYx3SlaFSEXp
2u0yHmrA9rSB7hrFyk2WUwIo06HvE3QswPf2mh9jc9OKwW08s9LFlQ+JbpYvL5TR
qQRY/La67iWLH+GUA4zFbZNOc2LQZb6mmXq2YObzoL/0b1bD2I2zVXjrmULse0KX
ERNFQRRM0oay+sLCxrMrqXdFbBRTYeJ6V+AJZSmY5MIMqVbYb4tDYyKtDi27ahIC
uW3Y8B1cHvolyBSR3DGWl44pVMyfA5Oa29rSXoVWq6YwaBefHtZ2CAub8N6GEBn7
DrM61Cwy/FoPNy54dNKby1XSW3iEBP8VFDdJsPX7fXCUiAkDB8Q9I52OVekWx0ev
mBNk3ukOBLukmSKnn97bnlao6lX3+L23yL+mfE7YrUPxCbvcnUH+DvcPQuTgbGDv
3wsHSEZBxe6RvJu/eX0Q70+N+4DLyEoyaXABch2eQBikl8IVaZwjyK5yHA7VrQGo
Mrsb5lxKUXsVaNnY5UGcQds2OFefPEjgNtq7GEjnSeqBfWEEJfIe2QLmHnkVg2Bs
4qg1n1REeTco0KLx3XyQ/Hnl325IwEYaeRaZe1ulBIiJ+KuhiO/iCtNTCRGtQG+A
13um+xBDQgnItW6BGLLT2O+/v8kJ/qGpuDMRfMhCy14KAfo/Vr5UkxnY8Nn3Y9Ao
uGD5O58m5O0WegL7DWCmsYm5eDWUUosY3j40NhKRiaY1gUeNou2+e5PF4rU0XsxC
wL6UGfcXnVPSwh7BYOojfaVLRQa8kFxgRIaEQQ2OgN4gakcLjMgMNU80T/exH5d/
JztV/yBcBsiH/+2Hyq0CRUXtUYUn0LZ4gQSDqyDmfhLvOXZYrD0sBCVJKdQu19Kv
buuoWktPxYqoLtZrpFAFv6cKKG9BHF7HfhiCqKsQTy8hR8kN3g//5T6dRvyJIRef
uIyPr1nUQRgsO3iAkhVW+omp7ZE9YG7KWpH47vGNxGRJsljFgf/AArLgpZgaitBX
LH6vRwwavff09MeqsSUFP/ondmBWAM9uimWJ2fA/n+b+IrTpfRjghcD7xn1P4vxQ
gvYOi1mN6j8Mky4keO8P9y6IT5w+Cr5Vr94KaNCmfmc+eUC0rZbhlFno4QP+p8Rm
bDaKHYWd02O5fKqwAlAbsL+qskedTIa32Oq8XKnITkVqusiuwSWAs5whwqKRgbRe
QO+hYtKIcOn+W/KD0wSB+C9mH/y35DQ46tq+zTstCwrjV72zN+LCYxOCIJrBwKf/
jiapno98jECOOCSI2tz1E2l7+bj3YTbzoZzLQEJpiTK/bxSxjm59+tH/kCxjAEYd
mM5i66qVIrOztwvjQSKoYy0QqseCZIxxSCq7H3qf5N1a+J0n91K0LB3TO6s923vg
OnQHgNiMkbUavgbk4D5a1FYnjVCKt4yj5YwPpyreDsxVBDNK4esVBAnXsexADxXp
vZQz1aCgVvnicO1uSBv9mknKomfB/q/E6IpJ4wlCpCX/nNNw5RFjxksZ3ocns2dK
vyvGWORo5VDTN7M4F+FbArlVPGyQn+hwGM0VxvBCViB0sQSHobgRMtbfXO7zDiHY
ZTg/RAJz85OCBek+x5Slc06/OG6G0/bl4WFQGEE//kUqZarUZoiLLNLt5HFq5bjY
GQwawvepinR0VdtRjDJ7oUizKDiHcYEi5iHKhtIWIgqnKPOoZqc+71g9FPrtFjTj
UNOHF0unbsUqbThJPRZAKcapxpLUGK3jWCIw63aWiuUzWoRt5iCMAyBOmNv6B6Wx
3woZLHEPec1WCLOjt3N9VOvSGRFeCfMOQQ/JieSkrP+4CXMaOkl39JCMjTyFkIMe
ZO48hjqPDwVyQjq/75Do6MMAp60DOG3sMcFMcmOUe+m1o3hJmQ8Fb4wSLCtF6IJx
ydAmD4zyAyAIPTHCs0kPftCdrT+APzzVRoE4Ls4mdYwpDjqztdny9DXhv3IniWkP
ekn/eBLyDrZUFZJ7OBannDArzcBET+pnrLNjA3/u4z4A4QJkZy+RTNjcl3szdYAc
yCBZ09XKETA0rMCa4KUADQY+rEX6AUfUXbnIfPXlcQ5H0mWZ1CY6bwkV03bBA6pm
jz25PFaGbHz2oDUqfCTApoBbGLjF8Dx6cf42clNDjD2Bs9tZbULCrA6ziKeJPhSS
xleq+flvY1EtCXc84kB6lM8wvCBhFxEahjg2dKrg+cvJgyq9xSOkoi35FyvbGJJ/
qwOBz6Gv2RFcJ68nhXlcc5hmDpOXgRllQNbjqzPVJa/8Giv2Be0BvisVQocTGBsE
Gl35UWEF46+gJBkX51i/ps29U8eRmTFBK87e79KLLvvZ/uCSAHNaZaKvFNMyBBrp
WDsLhYOyw9Nwi4eZXeBsvC00Wjeo7bK6iNgZ3X/4ei/tJLLuaL3VeP6Et4zY+bAu
gnqmP3aDXjAbThHZNgYvL8kyj8vD6nuKgXjZEAUg/cOQ4m0KC0RoUMeUuTUrmo6y
krDDJOiBLZP9aIl9FSXYX928QfwCmRslDO4/wA1dZdBFOah6Iz2n3WRJsVGbd2mX
0Dxbu+vI6c5ClZmRjHlRL+a9rg2G8s1CBMWCkObTAI8FbCqAFTIFEeSJp9QvAR8o
u0giS4IMOCgp4sM4xmcpmFo7fAHxjkIZPaFI60r3LKvsptIPJaCmALElHqAfL09E
v6pvHQOmIRlaJ0HXQyAbLYWremPX8qqDsGoVvwuqKZ/v87h9es/MLmFN4JLGtXSV
y4mNE1yASgM+owXbzLqifSuou0qJuv+tSgrGkVuhceXyzCQkZAg4tNApWLB4eQw9
m8nfmDBbDBtUhHvkH8Y6m2llHVGadJMt7+obnbHYEMmJho8fzh85fCpZINHH/bW6
6ZetjhHVPknDj7k8TRQG2WFUGjzvjw2rc2Xi9jCQIxEYNkk3zeKZmxi6s+q1mFor
6DFd5ZiFXUpd4eFsHAbMjbpgOzvGdCT9wAsH3ZEbFgFtneBrVbtBp4CrBMwsBUIj
skkTTz50952c3TUQkY0c2GqBSUDclxh5xLwz9ZICXdzbEFIoKdPfu5wo6w9MSpyj
d9twADeutkiOrMajXY7ceceM5ZauXa5lold4EogSwM5BIJxkBrHe6h/2uEZzjzf+
Oomc6vLApbikZnQcp/J4u3zbdIDG8TT+/DSKFIXI0g6sqhWv1KPzzkcMVUL3nsW5
w4VtxK4FfyMWWTvr45pfxdYGgoZCnFrrBWvipi5c6P29zRFmj+T7uHEIyXPrEk2D
aX2hM6AMy6+Oywhzx5DUn88N/0CZDuSUUQCwgJ+vdCiir50K63FZbhWqzt0CB10k
IzwGGbh9XrbvsDSIbve2eP8zC4JHaEQkFJZWuDAp3gXClltk56kqqj98ENKwyt46
R/d5F31fM1brWPKyJ9/TwLkTqUXZqZi1K0lesQ+HxSsCzFb2HjhrX/xucxA2nyh2
AxWtepbYYNX2tA0LsWFD0xB54/bMZFjnrlJt5PTl7BpLwdkOQZ46+r66grWW1Rv9
xWcWJKzeYvq+YPIRCJvLScSZwAUvVbMQyHmksuPvaIape19ftRhkCpWW4prrHvFX
glhqwafcBEkuqcIlF2vQlbNPQxaClOvM/jFo2T9mmF+IvDUTW75xhmuar1+6+X9Q
0gjKqL9pKqrx/kuTn6QKvNaBXGy8LxZIFDQeXTXlTSlmo0T4zXx4WCRDBMOZTyjx
lAnkX9crC8oPwFS0AfFrxh3TqUj/IxX67IwR5+WJ87CYoPvwXupDcUnOWuons2ZF
crEm3nLMbaF40CICEzu5HzfTwOMgeGe4R/pkrwBf1CXHTOENimfoj3ea8e06Xjyi
7RRHzduCZZVHJnlC6pYoF38yPt7KD5nrRCnSV1RSlSrZzUvEUtuypHxTeKOiTSzk
Cj55DfrvkHZ0pTiYlyehDfOu+32YeqFGfF2FkaO5o2EkrJVziVbrX4NGLedjaBwy
OMCuyW1LmgY8PJHvUWdr83lPS3T7z9qqFB8Ros1PYUhF15hH4YFzQJafZdM2LR8/
TqfmGu12sPTzm5bmDDjRJwvCLwvcEbQW0eVABiZrZmCCLXzFqFc7MBqK0CO6EIds
npZRKXXzNQDnh79mz7e2JDQKQZOshmVCQVNr2Cp7dJT+GjSfODqvGL2K15zWpKBC
jGFJIScjIAKoFXvPDho5kmPQU8ES3JbruqwpFjRUPLr0HSgDd5voJSpCEZbaw1+1
QUzTF8N2INyM4XzJWXVamxM0JhFpYYZleXJRg3z3XwdTv6OWOJAqvWZf+e/fsczx
bdML0FllH+0fv+wW3X9Hkxx5Vn62iPkIVNjk5i7aptSC5LSwM7xf5oRxC718ZNVV
hCj9FvWFsW9EXlt2Ajx4zkUnVdY+QuEN9AVejfrfwAvbIK1paNyHQ+pi2q3IHc7x
1/TNdoiHvM5QqMjVkZmK5D8bZav7no9E9ZAdeKgHptjt8vcnyau292LcfVOJ9Dz+
UCicPyqZMrhdmg42uP9sZiwhYC9CvMGgwNrEXw2/uZTC6pYV+lPsLcnEi5vJ3y9u
JBsD/+ERPQzXq1IERAcKuWQbSIZ4vNeHjaDOKvdtBJeM7nUsh9q7QGURHrLG/gYp
WwEFW6HaR/g0uCZNp/3L8Mu3IOebPdJbAkpF4PkfAi0i+k5f3EH9XDDBu14TqzCd
GuQNC8/psE1skfDLfa2gbvMqCJ3Jj1xHDl+Mtxdm0AwybcLSDBVMXFJwwFuE9s7F
t1tzXO5g1NkJctNSLMugBnzEFylal/jbp+rIs8pCxXaMLSb/1AY+veRLzAAhjIc7
r7NVYq8iJ91zbdMZOaX8dNez9jRAUxQ395oK5iIxyo3oarg+gE3bqwVZz2MOj44D
FrqbPqwcbTJGeMFWxAbUiIjqkihO5786SvdNVZzxD0ccNeFa3aU9R1EoMVoYbos7
uIiS2KdyePS2Go1lLjchvBE5pfVhjje5ktO0IwpHIjKKdhnpNWZK3IYCRIza6/Xv
nH1OXJBl26ScBSTiZr3BEbjOGmt0MqdCpZI95ytcECLVuE6Rq25aW14zMoewd/S9
5gk8qzFn+rO7EuUcwVhyerknvqQsyKCEN6wegIwk8W1eGGkfpQbcVGYJjQpd5OhW
g2xKQTTF6RyeV3jYhsSi15J/2Ch86s9BWQxKGEckWVhTRDTy/U3xtUqnvJscXxLR
zL44yYtP0o9nCs89nBA+dvikCO77HuuL1AjGmNlwlM0Z20uSyvWsl127jLq0PrZG
waMmnxW/T44jHEqCMwbnxz8jwk4cTGcjUyC5oAazcHU9qSxr5Ac40rTR2xgTCWdY
35gQzikrpB2XiWfwocEl7Qz80SF1kDg8HaPwiRrR7qq1EEQ91Y57txgTzqvVmRDP
aQI96KyVPCyeuFhbIPZhz5dXt5o4io/XXQM6eefeoCibowYrtUM5ufTsGXJQ03ab
JpMUQLUzn8LTR006Ub3ART6TPSdcMIh6JAK+ASRI1K1in26JeAcXQN+UWxLINU0i
f3nApMe2YMhIj8ll+gf6WH2SYzXnS51ODi9h6XyMq+4Jg4uYnERenbSQKRJmSVvY
h7t+F6JsN68TfCtW9zJ9Pb7F5aanLMPxA1Eh7O4bq5FkaS/YhsW0aWtMe1nCnkHS
fdRbcqHvZ60gFtoepz6BHYq9GCbTxgg1cYz1hibwnLSedRRHniXEXP1IkbJunTsi
d3P3aQFJFxa1NAOet3yKdIYBDiZTTkID982vV5BtTu/CrfP/HVEMAXM6bBxYFNzm
xKfm9P1oQ09tnCPXrtcNmnXH2Rtj4UFSdTuASxoWjIo7ttb2c76xI+j/MG+ijKfu
dLVlaypeJn2FxsYLoaqLQjDRbAHrTstOI/J4jkKSr30IOUYAfOWh3RXZHshzkCzI
3fx3YIXL1GNi3+X/Vf9rq782qnj+py+VygNJW6/wbXoRsJADe029LflE+Z6yRvWd
buMHqVd6ksey9bDXZmPBQw64CN3wYAD5rP5cGnkKO94tj6A1Gfqg05Z7IhwdK+Di
L6uWBt9BlMyoVjO+khkwoz50xGjUJ8GX3c1Xk+74pH7dgGxwBuhp6uk4srx5v2qh
fUif7oWlBjorPdEju7wSDAhvMjmyE2l6wW150wrKTz9SEM4Zk+/b+IDdmNqFgtu/
8ACpMHTOeosiM0/Avql2N98YRMfnv+5Al+90qmzr+saoLD6dsemo47fQoOZgo2/5
9Ea+2whwXGBpRv6vvdJcrZ9SLF/L/q57ZwRDNkTE4h0DBm68U0LI2q2buj/blpRg
OBdH98kITngRxb97nzJv+/QGBaCDZ8dEHj56NT/vMHLYTfLHe4W/i8ay2GkvaHQY
hT/L4Gv2NHMVh41bPLhQ1KrbUs4+eUmL3ig3C/ugiA+fSDSXPYD2B4rWGdI71zD6
8Zw0gLGEYGxwZKy7AeK9sLVLzdnhK4wIV6JA5WxzcfA9yPER+nFBAeMKIXYQ6Hun
O6iBCsSGzYF/IVZk73qbx1QZJJHRsW6GbMprt2L0urr5CG8ayCZba267d/5ROGA3
4PVOyEFKlF+83KmObbDYwzCCpSR04tKTq+E5e8a9GdYQhkl4AdwoeqvqvBUww3JO
W4qDIOt6Kb15mAjkBfObDa1SLXoPigFLZbj7DctKqLynR8rpERHpYw31orHS8znR
+8juDkdsU76qCzFh1/GGwByV/dIepg9ox7n9MLCqD4sFpWSwXXJD7ZAYtxHhO7og
8r59iIqZZexQ/fscrL/30pWGPjKKlvM/1jDD3MQZeLb4Tvx5i1G9wXCdtRe+mXOI
e+Vm2Oke7jHTHMrbCpR7CmowKLLOwNtia+zOABIcs806CVuzj6jDxpobbp6f9hbu
F4V22Meu/+84ERkn4kX1ntthYCiBphXxvcKLOI9MhEB42sr+H9zowPRtbyfahW7d
fbpjZM1lMqz8qFwkG9u+XSrkeBCQJJal2dJ02wqMaQ+37sGp6UcVln25EBOp/+gK
uzKvqxErMPI7cm/1bCKGlqbuT3QHQeMfUAHmbxlvvZ9qQsFcj3cbbu9UqT0KNdzY
M6pBeKuGBJWPtEW+BDuHPXDF6jHdozHl8fJQzsYlmtcjcPscGa/w9i+Rmvw64jhq
GNnszHec5MrZgk8iz14YieM32JXgRhdgNDmr3GS72FTleDlCwp/bP+TegQYROyrL
2qgMR5fLOp2a5BLmNIm7YMLor6+YNbd4NvwLwMjtTrR/A2c84vS6+p41vk2c8Hhd
cZ5E4/QlJQzy3hCBCI9WvFgS/anRE4pKKdS7wSbfD8zrPOjhKypNUFV6kgGcyUrq
EDVWM8lcsGF2qjVCcw0SFus0GDlNry7gC8rAXja84tRZISTBg341805sEXu1QyXU
eDnz6XujlQ1R0mzTTN8St2rnHDEDYiNStWfbo0FY6+eDnrjiKMFaN4ONjF6wvYb8
W47BaH/trIR2Q3fkG4F2jcEZXTe5/8/jfspSl/TImvBhwcqXlLYix8Dw0chpPN3x
ICbaLKV3fBvRFFiODIuDMHQTIpy7kEfnxlMZAEI1+he+UpnVjuFMAVGhkGwj7lhN
++cGKtuacgI8PRfd3X3w5RmIdhbuOSWNK749x/oLjTFlib3rvx8rnGRfFfW8y1A+
yBd3yEpgkxIx+THniQbNsNv3E1uufegSttfdRUxwx8i4buZkjvF6+JSMMVXRFXrI
vqtYEiqc1akezbw7J3UgEwJdcs4awd42Vrb7lbG04JG1Jo3zuc6YUTXSIfZyYUfB
UZCSH7EEhtRwwrfBgtVdp1y2AuU73Sga4cwPrgg4OZZp9xmNyJ1E5N5vzKVZpuG+
j15e4ClcPPb25AKdyCZO5ERh9x5onl4cX12aKglyrvj8xRdXg4+TTdrD2Lto1t9d
vmdJ2QLoOEmhf6ITpyB0otbjzXXD823DU3CVm2x0wYshVKpTKdUd+aJONNlGAD2E
3am8IIpCwhREO+k2xmrMUyKD6YY2QmZ1pzJwU5WCXKGGCBg00oMgLSGDBoip7fFX
EGdQW/L3m3gLe5QzMlIfUjdtE01Q0Gr6NRpJ/gg6QIfO3I7V1u5m5vCihmy5QERi
cR3AhY1cogZUURglarJCnI0Pv4nkHBsK0ZB0gDbny1Xf0ZZv8YMGRdd3fGEdECax
WnF4G3TI/YeJ+5cxtn3WEKbR9LTQKMdy5bG4WSVio375zSJbMlmsA5GR1lwm0Tqt
2432AbW+BNjFMmSKuaW+OgpLXu3DWlwg9+EySsQ5CtXfMsCnCwDarnEhI9gjoD0W
ZhbTfd9ouyBMXk30JPchiqHtL8snuyiH5QQ/7QP/AYhT7zC+6L17HNCSnD1qiMYf
2XDWP/VB0ms10+00Gj0PbR4uuHAZynRbcP1iCNkua9CEI14jeFitRKRy+wbg4Pef
6DdD+wF4F3htDQQcsaV6OXSbTolUiGKps1Bluxbhg0ajIs2rV/4CtO2ZuNXzgqnB
khOVqB+uxY2slVUdNxMsvb1uG4QLOr5iDq4KkuN55OKzjVO1Al0PI88abFcbUaij
eraWPW9+0hd3oSowh2V2tWxHOT7GUyIFgGxkSLxjAurA5u9/xUffJ/0Pm1rCMQ8q
s4HXkvoJCzjn55iFnbg/UYSzLXtLJjBAQb9zDgFzbWZdlfHkzWZHrdWrpMLMRd6P
ohYMuo6Ar6oElhrPnbHjArXKjfoDvhwarswnJYoJa8V2WFo7ArPmHx60lgkYRaIb
7MEnZ3oejHXm49XkJtCI5EBXEpiDidZmSZ7aBTah/IRgU6Mibb8IHqjVp/p4b9Jh
R0LGrrkaLDTiNTRX65LOX2IpOxHJBNg+iPeNt4oHDugQrLqqA2Uy8pQEOQ6xWaGO
R93mhgrMHw2vqC1+HDSd7hknfOHdvfnv0P40MVTWtJznhObOYgXl6yWQsJa/9ZFw
X7n0zqJbzk0ZWNwDE2LwwCqUc9nvPBUyurKS7nQJIwR1puC6iJ1lBqgfoU9icLV9
f0i1Bxu8/G0j3Rn6MgEHjg9VmC1eDYF7HqzRBtYrjidmxkqZ9o2LhqqNdYIT/jgJ
QptsS/MBvAWA5BFCGB1gMpXK0+nZi/3JdgIxxubtN0OdJwbhuAbPCqSj/9K0ucuX
wr1rCLajcvrcIcZaGTb3wofzCAN7KpfQvrX0tsdTiqHLQ8yYYPd4pvszeLkfjpNO
JUukE2cBIjujeWdcrxHPQG/q8cMq9ykrylMo6cUrHc5BABC3cQpl+SZgeDQ12qlA
VusnroalgDSZVLy/NZ8BkJ7uMP6dkJnZY3cpB3lJ60dxc344j8MEkEbXf4rJANun
oHAF8v/tWY1eCt1rgkGko9uMBJ8NKtxRIrkQosy1QifpGYeFE1GWQwAtCL+da7Eg
IDKuLqx12lbc2OmQR6sdk3bdcWqUm0GVbgmD9sMhZVcSB81l4fQauRO21JD+tS+5
y/922xUMQNvTy390AfQ2Ut52BjwZF7bM6TeJecW3KwRmRxUFGgOGpXWloMesVm7S
RMqPJiin5/gYrV8TWexzRbUOrzbpsDjmayxZF51CL4uKoT54CLlKVvIMWgRlwu9g
q63ItHrEJ0ylbcmrVlIDLvLRGOF90PTWuiUQS8Jo/8dmFcg7RGlfIfEuST4hLMb+
SPD1La18RAz9IjS0RaF1s0KC0P+RkyJJobbEpI56SzuodFuiz0jNDP7Cve0BfYPV
UV/tEsiEKM2GulXDhfQn/8IS4V87IVBGV5wDcxt1uv7srbdcBTz4hmY7CrnEszOW
i/aCVA+z7ez8Hw06P4vUQ6dy5MLTmYWrnrfKmTMlUJ8JNH2kftaDQB0istf7NAeq
y6e+S2M4rXhopZkXepqZvaNWVITB/aoERT9wF6xJ6UEamdmCLDsWgQOWrr1uG8PE
4+z9AuSznioQCS41JpmOvc5htAgl3r4fqLEISd/rrEblXD+sIhZagF93BdUKbaNF
LUa72E+VwrlzSUuyGHGxdEJOmbJgzEsmNaV4K1KX1NDo07uqx/7K4y8NlAwBiuOy
mvuUGh1tfo3oRfzrxArp4n7Ls9feV7aYM/raR0/F6tFN6YPcFTg7/hRIsWP9UnPL
SZVYCzvUe2h7qkOpJIW+3GBpquAfmR6Ra+EnG2Dx2iJTrvc2pId3HjRIkf3XkuMi
6W5yjarZxGcqnGU3lJkUgBfzHQYjx8UtaM4gYXNIWavy1jW6YFGsVwb6j0/ydp1K
zFDzIUyZ1QjriIlhuFClFOKpUA2ynlgtEkevvuPvTgdkLhUdjPppoQKbKX4UC5xk
y0urC33muyxA5HXXOL7aDVPlUNJ70Z/Z7vzOhEzLACdMLJjLJA5l1RtINAWI7JHP
FOweNRSOhnJZvzvx2MgZc2zynUJUCsaK40fSh1/i8iDPfEVAzkqHDmkggZ++Ulcu
yFnFE5IMVqbljCDgwGBhKPfRASMV+HGjI1JasZgi7957FrJYp0Nq2zAsJc8jemQp
OxvkHsDRdzkp3pElQndB79uoA6iS4RVLdjjYMr4OFN0fs0acyLONz/tLR82ncUE+
9NR+Ai+eaBsFifEaI9EWHM/uaih4+KpCIdJ2Fsb+cknhnqkQqnI+5YTAtIrZQboi
/0SMFKN7TqeCKDu91WZGNyTzsJQoe00IutaJaEOTi1ngB7HTZ2RHabQP9cMwNyi0
QjyxTT9KYc6kAZj8j54NPjvLGHV5ISHd0BOYfjg/HzUWHZN3hmd/7+mdZnye42XO
JQ49RDef6bYQkmZ5Lmqf8NOTFzydW95Q/ChPzrNsUpTl/GG1Ypv1kYxhCEqMUc/6
rHj0DocFCsrmRdni+v7W+CAyEA/bjRUEZB0eQI/ZIuXMjsL8DIkTnYjQWwqxlIER
WTYzI133x75M99ulD9inan3xwiDgteSewfo3LtIeiGPP0XTpc+YvdQQhdbTPLssY
OYkZC5oaW6X4WhW2RLDTtuIQ6l/iQgR+9vJTgvV8hFioqrh8Q1tDqFho0VdwYbQW
HMb4BFeH21jcis+gi6EV/KAirHPpa/f5gXbH4rQQapoH5oRNDvr/l+awvqIeqp/H
NxsTpf87bYI/OUJXas6jQfKv9wcWwWDcU8l2Jm+zvrtJIyxX5R/NkY1rz5XFtxGa
i7+4rOzy6IyG3+h8DayJcgPkgWQdzZEGM1cLNL3ilRO9lVkpgwlHHovAU1+JrG/X
r/NaIBf5baOphJFcvLz1SF9A8sLfAKtid2OF+sV3FW17VDOd8VoMudwmsL0zfEHE
UBvM2hvH0geAUU1OJay8Jf0UPurrwvL+52CrxaPW2KjegBBxl3/kkTw7ztyt8MlQ
t9L3miA35OhY4/g7Jw95CQJVdCU770k9gvTQp3OSUU4mboapZFYrBRVxAXcRjQTk
qHeCBSbcDrMUDzHiL84pkB+42MMHnfMG4K7ZimzukMGnK5etUa/BP6FsHR8eLzK5
plNm+btms/LTjNp8no9+9kbICoub65vFhTwRGLjWcbC7fzP7wbBV1pPlzLzKJx7G
kVPiKTaur4kv8hJiAaNtD6ej7j1dvJH6+7nv253gef+VSeufSA/yBG6GCsVN7nap
WBy0ZD4gZGp1CdwsAlDxGNHg1rxVoJ6hQnygruD34FtR7ZVAo8tIJeseAhmrHS4t
cOXvV2O3wGZj/18G9vYk/oRANWXuOGN+Nc59cWpJ0eVyovSNW8ZkJXvC9IBFNczu
Tv0LzdqqcxDElB2PSQrxDZPp2wZpJ2VmRN0oKuRKCBUSqDBjwZZyDSydnnjKJR3F
yNyvmjPldQO4VfUGPdbzG3TIRb0YA2vB2rYB7zQqAN/lNZJkO37y0PPSABDFTxMf
rQfmS1khVj8s2jk1VL5fnEmldXlNEfohiD4VkJAgaWXqd7dXWONaiU4l3z1E9Kon
p+WSKsW+jrjoZkdSpf0ZSMu5rvmkMeeWgyDm+tdu/Ux8jFXJdD0Pne+QAlAFhpjr
tq9WCERT8ItW2oGDGX8F+q1sKOmuxqDBPpUMwdS/Y3yj7sQ4T13Ysmlzv9eVZsyV
mCZdafHlCu9PxWoO3GQv4ZvJYeGuWY9XDOaw85Nz3NnMSd7Mr1lCFHpfqnM7Sq3X
Uf0xMtBf/RrKfE90C3nyd9fR9At1QPZHJvUsYGkmD6UbYIOk5YH5iw3bogVZRTdf
0oDKqerzyt3pIC4LVEhL5+eMMMrToBvheoeAuXBTN1OjJ64BMQOmwQzkAvgF03tn
4oc8HfOVtNGPWv1yZGhIMP693rQxS0ry/NFhDRVf61huDW7nmRspXE+Sx2DIdmLP
qibQD2VP9WL/3CiR+9NkUt8gA9mcW4ww3rg16OZFsOyPKut9P/vA2l6eUmWs1GUK
otkHjpejdo4o4UM68LreyVOMSy5IEDPsMwhKc/Kc+v/gd0G9IsNgellb+IMxT1T2
cN9T4bhP3Ksp9R0MAwRrUxKmggth3Ami7UmRleBk4Uc7U2zOg+JrLphoGYGRqR2+
gYuy3vw1yyNAV3iyJytNQw0yxe1TU686fyuKaCM/dYXAZYGDCa8NVHjGUPr+uL+0
sPcfzK7SJ0PA2dYSvsAUTaw+f79XtuLHZymt+6dkZX9O7duqfVhmnZ1fxxfOfIeM
DrjPGA7NWUiyJDYn0TJ19oYc25nlTEQSQEzO2kpfNcoMlJDfy0EfO8QnsYPTPJ7k
u/GAYbWK1XfdcQH44ighLbcEW7nucHIWzFKIveihq48cIRzh2P+mSuxo+3a/RVg9
1oI5pb8laj72fwGDy7AsJC0TvIrMjpeFTicZ+WQcivG4MlPLi9shMHk+hDMUfBKO
4z9jUSLAMEvIOSnuWGjkFafLzPp61lpfoS1wfV1+eUQVQ4fVKmMOCvnORkZoO1mD
GLnGQfPDRpR6/whb5wAmCwYqZvlaErU0oyVyLgJPl4oUoErzOgHhvrvN4aODHsgN
5phM8h5sUgI6QWGGjQ45neqoJYblPJ+dXyYX04cMfDHfaagYYHKnD1JTByrUOxuE
EMkc7jwFTUCQ9X3H4KKnq6FB3V3FgHwHLXmCPlQVLrW/oXgbC1wUt+2u8wfIw77g
LnpU4PqCP49j5csd4QapaqYSPZdmKzzzMS1qTSZTtx4FD6js19rxaTm2bOMi91Q7
HoRN2JOZZ5aUejf48iULDu4ppKPRYyRCmsq3j2FcW+Um6pGWTQk+pgC082srGKUH
6xGJVJ9qbqo3ZZZCAAwJsonjwtOP2WjGmXY4AJ74ZJ72KhcIP21OBQ0tnb+C7Ts3
ovtK36pKC1VFznJFlpoTHSOBI/1K5uWZ8SdluGXL2Td9WlGsL+TNo9TLMqV++hNM
uUXomvOUWfppt7DAyTigByzwvvNS6FAJfwbtVGLq/AJBImewKwzZTovvMtw7tUmW
nJoFxzT3fFA9Ml3/P8d2HrCc9Yeoi0K6EGsLsaFtYFlsRJeoozETozv9mN/ed7mR
rsffu9yfle+NvnXQxM6tuJvTuhydrWtYZRr6YAcOI3U04CQ6O8Abo+IkCICjCkAI
7hH/v/rBsLqMC3CVjHJt3ZEI3A3Wr97OCKpRvqdQdwvSJUeJe14Pk7lOjlc+P8Y1
0/6Hx/fNNvhfmnYjneEA+z/nQ1P0k5WTruWyyA1Be/cMd3vNVEoZ+EW1DnbwgcEZ
1q1E3hX2Fo3ZfntzTxn4wSBmhN11KCAdAFodAalsXVm/515TCauI4DgQhYsx4+vH
IdsOosC9zR/jVtqZspFkXs0IilOGS9BPS2/a8AV/EWX/KEzR/6vkFb/HrjDTsCaf
4MnwQcdzQlMZeOX27qeUZyMqLPXaUCzLr/Pu9vtjSXVvOMLsORjRud8p6LxTddjj
uUEyjnAC30czUshg376Ds2YhH7HQz+3xMVq6fMIap0fVlZAuQk8+JGWT5BQ0OAkL
XFdlmDYEOeHACSia4hyzh7ZWHUCDzERwRankFtog5hbdJfLtMwBI3s1DyTfmtqSi
ujR5R9qNVHdy09gBZzZPoMC2JCs1JoX1MR9opaqXIwIv2rN1RhSXP1NNgDKBzimq
QGo9xUn5U0bxHmlGfFUZ0ZaTjV6yubhYdFyXCHnOWNReK+q8vUSOxjFEORmF0NZT
R1ozfNblVAkwxmik5cuPQbxy/6CQgzS7CfhVbsS9M8+BC4VY3vYJqTKKpJHSZft+
wmeUeKKqUbLJzER1OLJ40lkRNS0WvH/FYIXHW1ElDfkZiPthPQvF+bjSFIXnb6vq
Btd7H+ZfPSz6mQMX+inCggUw7zkGDszv1RQxkjlu94n2C2aZUPcRkrjA2mMwL1GV
TPiJWUUOua+NzzpX2JQrv2pbRqd2RKsfxD1fa8/2aft0S0Y+woU5EGUKPmJo9mm5
9i5wdwA0KlNzaBuudH1DtgQ9KLQ67jpDvZWXd1nijQ9uwOYJHw73aUCZPJQpVCjp
i56eayfT2kr2FSUSjI5sDaTKSjXU29730VmXQ05rA6tCqELcSOddtezdu4SjTNZA
+DfqqPy4+3sput06QhzcbdXgRQ5xuKeKOsaQKYWNJa1CPhlX3Tjff4iFQXtMNvJd
WaXnyU7z2uWAr58gchIbNYr8PiKWTAmCUkBEjq64XfcgIcOHPFGsPGN9tcTON2Fa
5MZKFKngee2PUvVzPYoa5f+mEdwzQWYQ59fUjHfp8c6XXPHR5L1RRHmgPjPDeWqe
avjGT5K07OQj7coN3XVhM+Nszo6yK9hCBZJ9j23wGnycQvyobBvNztjDnNC7SxjM
ZKebxJgKJXBnZfYnxPRhTABa29t8LYeoNxcbZJokF9UalGlPEaq6uNfX11+JCk9u
v9/5CpJEG3/5wohNboFtiKZiif7gW/9lNdXqHY7NJwYzscKJcLthS6mlzBKAl7An
R+4HsETU++5pJDWgbB5QP4u8Zo0JX6tkL79ja9DMqN5vNEvUvl2YbgSC6DJ4gow3
W/jAhkTspAWBv4Wzs4Wn/Ws+ImGteV55a3dqzbBGeCrifpuZ5DFAlS0rm658LQFz
Uy7RKe8hx7GvJ+ey6NoLymzZw8Pkl0eB/RTX1jWz0nqzu//9MpaAuvwdIcdFP/5l
2kvMF6G4bqQ8NgzLU3sU4Tm7MF9VcQhfE3MWFWIKkmKEdLArdYN1B8UUG8UjGbmU
5hLJd5vT7ioJCHHahgsFzxJqh0PCIcPnbOrndxKyJrEx/wF5vy34eaaJ1AO0Me6e
R9BpMY/DUk+GpVQtO1+S17YUScpubZtHMXD6GR9Bp0voLu2ylkDpoiYniGWAVYmh
Kg91jMVV8+0ij2RfO5zNblgjFzs98+T9RqF7MUVtR0c91CPU/fXhTDSK7JM5DkKE
rxXK+ZSkOLKiCSSL0kNQH+DvpoF8A0d344fKm/3fYpSPLK7JyxZv3EDByWKpVNNZ
oqobDdhL244WOVoe99deEQJRV6L1JQlTDJdxEvUGKpA0VFmqh+EKX4HdHHVEBIe1
/B7k/mXTFH2F/eRzosDEclIdHv6Ru1/JUmsvuIZwHH5gvMGOEosKTH+4HsSsxgg9
/5c5Wb/NiVd3T18/1oVGvgd8RVVUn3T2yDxCPY4GJ1tbjwE19GU/GsVTXzbffnD7
5uJDQPH/FhLoTKbXAns4GKYPS9ogrmo0K51lGpO6c+7qLJ7iDp8EA8HyiRC1hdly
RbmdFaUEm+7yXNl8N0deJnPjdrX3jolE35hl32Xs8/shQHfSWxizMm+oXI8LLCv3
c+zd9Ql+oYHbPL3kuSFTHjPm0DO7o6M3dPNFKp/5Wxz+6tcwaDkAMQ10Ny18Fg98
5stxx2CS0cVGdSQg6uExm2m2jHjY/L/AfFhiwq63Qp/sEK7SEAXpMyytW7lJ6ruW
njRU56jq3EFdqjpxvJGCmVTwQZVY/2pO5KJwzlPkIuyD94vyHtuE8nmEGcebilq/
PHYNKbgpMhFoR00bm7XNkRoDypRyXuKtfXqCgfoyr9F6rv5ElGUFniz/CKMX/uxf
fIXH8bJ4U8L+LT7lm4MYt4shuLk60nUXtxtQIT6oPrt0DIJ1XYeyNi/AeX4cvC8d
70GEtspGFaSUml56P71+Xe58EGo4yfC+9Odx7AWV0g+JAIUqyLyJlHeqamPIhqYH
ckppr83NxV+xRX64XZhPQjPGEjFJ8nD0azYLt/sKK+Lem8UJy+USONBc4OsMhidY
vefjWGcmIsk5e3bEiG/25GNL7QqfRF7N25ntYPIM9Amp/U/k9Zso542FP2wju/s+
jwiNxCM415TivR+Y6UbuTIqwauTFNCK6KVrh/AzoZC8B2gG6cZ99cLQZyOaZ5Xoz
R5+ygUG7Lsk+jDFGtoZUUBI2QJOlTlYhIg9g680JbVCZ5X9RnLCHgq3BjUDZo++l
eLfxdK9OfwahLeudI8ea8Kwe0FNN7dPr5ayGkolqLuVW3/jlh3QfoXF7KuoKYh4u
WEsMkm0vYH31yk3Sl/sWqCB1/DlUBPaklRkGHL9wuogEFnShqbcWVXEGzwRBDYMl
E9FuXqSlLsL9vZmEkYbXDQFGABEGL8UOSo2kdHld9mDhLONEkJQZuP3l58mqrC6c
T7CNxHGJ4Vff2EPyJ/iS9IV0AqHlr70YLIq6hL7YnAvhf+wjgvusB55Yt697Qxji
40AqKf1Mn8qaiMwIPguZMlHtEqAjdaj2MOR4mws4YT59QBIwm1X02JsdBRqmo+qk
cc6NvCaRHM4rkym0nSjMdux0CRMzai76GzbAAPy9FCJ61K8SgejMVCx/VtFdgJcv
XSY9VU4heca2BN6KqMh7e8OL+dPNAKlJbyF9tIo8EGMrRyLioNxz3QzgesAQVuzW
2m0rCzq846ONXl5NX8ggknXScB5uDOl0svPW8WF5drkPgz6+ZkPOH+jA57FBDPjb
3l0yOxvPUgV3ElrFRiEiCl5ofYRxT8eQGkpBOiPkmv0S78ntVL69fwnHLhGNL2QS
G3l+qq1fBYWDSNf3dGIikDg/dh4iT+VkcpsUjnqBdJrfotvTh/PbcRDhomLO0PHk
elJ8EooR30pS3m9eE59se+ktm04HxfS/WMD4cvOShradZ4u2eBzJE9dbc7wOjg99
KNQ6XwpPkHPM7T5Rd0MQz3t4LnEXZkQJ+NUxIJ9ckQKa+Cj/AZGJ+WqE+jMHKvx7
R3wZvZGy0UAFgbHnMETBx+uaa5vO6H0DuzCzqmHoYjh29JgV41upMgjLizV4IeS4
ELp0xGwNu6EoNeGLAuBSb70m3L4ZxJr7wiJrXWKlWc51+dqFmURm6uskomK81J4K
kQgvZBLQ6HGJS8VDabqH0Tgz+TLNGi9gjh8rRg7LS7eD1MubREAFbPad2BJ8fVrV
PFwpwuf+OYDaeu89ENnY2Fshx1DKhtom8ttlSGHYKxNt2QwaxnxaOPdrn22Mq13E
5gdXDB3zdU0S5QgaWSLPVcHQNdxgtpZ7/HFFhXOPMctz4XEXU8KoAnn34M1/L9fl
F906s+gLMgVzupEsJifrmgmlZezgBzpT5tAIs6ruJYKScIVmaKAnq3EiRmDN+Xg/
InNxlsp5GgJegl072N77FmXmbq1wswP1ECT0LcTJhNdVfvZo6C2vmEGymStnaB6q
2r4ZKvl9D8ITTN2yUMJ7jBj/pCr77Fke8c9mzr3dlFdjjHruR0JNkLoPIKEgD5DC
duNScNbO4rpIOYjcxoqCTopGH3hm1qiTW89hG9JWQ8p3luETTK/+Kb9H5Oab8c0X
9sUWpCvGwtzcOB/ZWwKTsdYNsCDa2IqHoKJxXR96O2c5vgtDalNsumA7PJ4WoR4g
78xWM6W16ddpcyFBO9IOuhXWXinJypyCVoNdBZ5b6uIGIZr5lzAPyrjyY6TwGnzC
wc9BNT+TbXzvtlTr3sv7Y/brbGxHiowT1pJaips+z5SgHKlscmImggM5FyWvxNCs
H/61EKO6cO4lcxMymox8Wk2s9QVCNAS5qgvJR6e50Dp3puGTZyYWpqpOYlevBaC/
kqwjY6h3PJw3td3NfX458VmdGrj2zAr9qhXMLpvx7dBCCghn9MlDZPA/tu4QJy4V
i8ff+KZP1GTC5b69cwLaJ08NjF/sjh6O+eOsDtsa6fdddY108ywrFse0FWKQaW6d
GxLX5Al0/1N+k/VeFvSGsZi/BcMER/l/7hTzisZ9YDyFXD8JogY39QM57lLNgxwm
uNinoO3IW32KIDnw0md/h7glUyKycM4Mc9ErUOy6IaTIsfKXcKetCQuyHQFAU84a
KYS6Mq9C+0zQbVgOCwZ3n9/6H6eCWbWJWdDLJHYdvxkJwzioq929vR+06haUpxUo
j/xdZZsVcHxBzAakn6CQfutKeZHyK27r6z09rU61SgNfUVTcohBqZuSin+MgoSvr
5rd07OynjmA8Lzzeu9/8emg+5CXz/qLNkLNBVZF25g45iioNpy95soWZYV9vxyBq
8BYrtY9b8c4Rg5babjL/sCCHmqtmG8H1Vmvry25ZeHo+dhkiz1fSoYGtaAhNckU8
gJ+SSvDRo/sNnzyJO9MNh9YW6AcoiSvH506utDSgBC/jim5LPGGsa0w5q/xjzb+t
BaSY6umsYo7GC3rB8wdM4O7VXKMCWra2Sc6zPzuqv8i+PRP2ttsAqNDJ0FrWG01o
6n2zjDC5tpWVhoMvP1umAK2dPhGrgmJ9S6M6xB5bp+yk65gckucn4KL2ngQMSLfY
phXtKLpWcSAgGfcN9drKyDc6GvF6faBraEGr9mRQgXpFP7W1dX1a2W9E5ouEarYX
x3h8c6io7+Eks3eIRoieN4lOJn5OxRaM0gwtr6PyHQp1/BMZ6B+ZjtBp/kZ+Slu0
HK74f7jAilSU+qxY2iPdVloTd7YvKGePrCl9WQxl/5/vVLnpzLkHilDVPS3RbKok
rXugBGSsAwi2mXoxQVAQpoMeZkUnxwMugI9WJJui4Uf9mMfvCXyq0xnZgH1aqdef
OyH1g0rSQdvGzPay129FVz8N807w1CnH77+Wh8Thfs3t0eO6SCHqsYwNznmpv1N2
LNI0F6jzoXPx5ztDEJyJSoYjO4HW36rDdWHcFPEpxTiqy4FnOW/ygzxGx7GaWS2a
FMfnkh2/3wwKYqnMMM6BVGdUtH3I23UTSgeiRwDVqixOZBejs7wnl58KjoJAfoGr
qyJjVYe38FV/kNEnCkDjcrJf8d9Vqo+F4MVPCcGMJqpe708vCchOyAMxBEox6txP
N7+L3uRsEJKNGsHb0PBFuv8mAVooCRDfJzr2UaZkTjLv9fe+cN3PUqP1elFbAxZl
O8v+QTDOFEJ3oGejmSc/jw9Za9SiotUhnX7VVO2F4tHlpxHTB75p2vYwzXX7xuP1
GxxrN4ugcUVpiMg/yJLIG8Ik27JGrZQ4PKq2BIYL/sbRM32KP99qeGrxJCAStaO7
HuEP59Eo0pApQF8I8dPwQoB0sGtb14yiPwtZWi+FYhoMk2lnxpbpnLwZ8JtMt1gz
9mpJJXOqEmlLp6+WKJ+aAZRPefSrFcnS2yBddfo75x0u/h2XZ7qBVzAX3P+mXCGf
qONcN9/uy4q3ljNCdm0Jw/kWdJXsLc7c4tUKRb8+B7FnCKxUGjfBCM/adsunMJ9y
5z2OM2cKGIk7ZRdOKjL6/2HI+XuHavYhk/sLhDtvPY5CNUed/9Sn9xxjjox5MXkc
Zfix5GQkKCiOAIcjv+JmQPMjKpUxuduAMdiFI0uEw1gDzaYO8cLO/FwTUmdx4nIL
6heJ5uH13KfRFAR3dtjr9SACUrkODz9xkDnqFFC0IXmMPfF6fGlDpBIjIFzI+afs
Kiv5oD7nulmvn2o/6kwlhep2YESQYU7tmJ1z9GR58Eo3eZrTWpgAIonDE4ixqGj7
vOE1tSE3QPw/0RZzfx2OBWZkmwjh5jwZ/VKxhFSN75FIdkzbXo/2nNJKgBhD36AY
SyZq9PfagDXbO3ebsoFBxnzqrI9af/TrX6eRAFM4IrVu1YsjICaJeXmpry1AiTC1
iUegKdPD9QmaICpKHb7VQY8QIYiNGpXroYj0Hb1EGtB10tv78KTEPttzZBkH39Tw
wJLX0a8LR+tSdZNXK8BjC94pO2lRO9O+FQoU85QISMAOF/aIVPTrhOZjb87eyltQ
SbNj5Cb8GDtWr1zoLwtAmhapEl9NDLXX3Rfx4qbr5nS71ay3BHesZIeFABB8FqMj
hbMP/MkpbdIOaI170Z+2zt/1YBAhT30juXYRqbKO122USBTBHMxXNlMr+7cq7425
lACO22OD4HdqHNz3SKhedn9AjyYERnekUpH1f02wBIFlfEK+bAF3RQQoH7LAT7qz
1YEMPWCH3IQhXtEjPNIoAmjnHmhCc7Ak7DbmBLZdR/DpxVZuF0xPpS6Sz0daEygo
uSYunst/X2laRNeaVB0L8jyC3ZksXrtgi6E0aTVQfeL2mQ2h1mjoc8P6wGb7T7E2
O/MbCN0gzNlV3GcSyxYYYmD2Us5QFk7M6ItaTG7uYExHKd/7tjbSsdHDhaxmaaCr
sM3asSEQd+OazBq6DoNw1u+uD1vge6gojgjXUzrgiHUUUaHMboCyUwpi625EbDrc
kha/UrksOMpmKms2GJF8AaAcKTx8fG7bKJeVoyGTji05OoHiGHnQLRUzinoy7/FA
NfQMEVXv0KI/0ag3zfmudgOpLXQFw56ZMm1rIcwht92edYEI+sMrgvpYYdXKVR+p
Gw4L0/T+RtvKXhsLeZdnJBszl9detEN/ASYUZUFMIjDPTELFgRVE/TtTDyS86PAS
2sQwi3lGR0n2t428EqUIp5U48i3iFG/CCEw/qpnhuRscP2rVo2+a9ua5VC6YZ1QG
Ga2M5u1VU3K0xXcVZyQu48brgArwLqAPJVC5RHBNzfIKhlBZLOptaetH0PSaYwLO
I1ipko1kMQz1jcUreJ1QHEqAPUavaZhBRtT1p+qRfiEDUl4QxDrMUZPX/3r8eGIp
A8ny7iwik/U7CR63yt/usu66zB6yXkLtetqzxWBuUo0a7kbWubUX0h3WJib8dabs
j+wC2pDNDFTI40vD/3GJvVhPTroXUj3WzS+84TRnS5Qk4DUbNs6e59vyqf70KTv5
fj6vVK1qB5XkiOV/4ihYNAD+D2aHUC6dQN0hcEQ92bqI27c9LZ5A6xkvl42E/SWw
J3Lq3YI+/c1v842VB9Xk1wOSzeJrkKzRMAIChcahwsmWX8+WrXxLAcEr2lZq0pb5
ZJkWTY2G5WvfOHclCi8F9uE2e2SCMgH5MMXbWg5zyvEA+lovFA2pm0of2Njtdd7m
GHNuYPpXYGQsQi+krj5kL9dhxKtOSch1QV6uiIbngVlHiGIjphr6APx4RDJRkofJ
xkuDVe6y4Mu4wXUqJWn0v0tEPMF1670P7rXHgG3IZza7oavb8gd20AlM0r6eVloJ
b4uew31QLRpD3hTBID3NBput8NmQxrbDtlOJeEx/k+JxYU8kI14Kq+b+FEHvdDOp
0KG07wUuQL7afaA3OvDSDv70lRCdC5zjIZ/+uDbqDtIDNAuqthzELTHUjZovjF2k
PyeL2i/ORUPwNdSQFLwSWg8r1K1oWdPHcimQmj0CT95dMJY3hAl4ImED/S0W+3jp
tVWBgvXZOJqd09Oq02YM/IJtRQFcVSE0hlRUeZRlUaXaDN4M88EBgVs6iOyrZ90E
qihToiTtQzk6WznpX4pJvlvRhV5gjaoKkw+2HGHCxssXV/ce/1A+6oBdN3W778YF
BkFjekIwVIvgRnbieLyEZPjB8NLXEb7SIGWbS66t9R5wpcXQjHhIeyMB+VlfmLz2
pDZNnAdlt/w1exyQsfeRgYq80iuyXko+xK614bWCH/AFaFK0NNZXBVYpOD4xrvDG
+EdCi1jwsC+JS8pbLNBhjLdbSflLzD2MdJdwn7c+9/zxGAnHFn4UeKL7gIwW6jlc
dK8P4GKTcQEefmkP0BMlb2IDyONVgt4diAyPlXJv4NRjDU5zgLtlynw/aynSY4Ga
pI+4Ch3mKK9R7CKN2No7myqBtoexxyfF0Mvblo1XBW67vJmRuVl/8o1RTYlv0qDo
WMN5dZ1LNj00jOSFAMlXxKP1XssEQzjppBCgIJ5zUnGtylDbem+CXVDmAp1GjLEw
Ul0UkegaXdCe6uVxy2z1xt8trrpzDXS1KEy2cUiACWwUggtD+puQWMC9lvlVdZaT
BF/vDoGS8yBsFwXstBcLSmci431sXfav4TxRFUjlsQDeIfi7kOFx7Tml/lqpgSVV
oRa4LeuV3HDblBRFVEG8A7kXZKptIxUv0nkCclFVTC5EspZRe2dkLj6xVdwBE9gE
Ww+qnB25uctkJsALSFU6/MlqbUzwiFXbvB0gGA9U490iihb84OyLgGADMotQNPPf
OORKYObmaL4mUqCkFn4Wp5vpDtDOUTnzYSHZxDEYDQjRDfwGrJbeyIbXSc/E2B7d
YNz9tRu38yBm5BAn2cV13dgNafsAw6gMr8JK12dhWz0DYzzX0+sQ7lKPSP+v/8Vd
cJCu+sn1dLvRaQuFQR8Ka/fp0nD8qWCDhMRTM+uQQuwlQLyIBvf02JGpYpGbnZan
llHle3mHyRv6sJwCB8x6jkb5dJ3uMm0bqnA+SpHLY3wAPWz5WTy7h8OHkxTg3mb7
03PKVc8zlzHV7LifsXDSDC3UtaNRSHimd19J6/VgSXEKbwFCcAin/Epo8X5uZU5B
YVW2wGT0D3klimj6Tt2FRq+pWgsK3eoO8jD2cssTU1D2KW02vQHWbYxahfanRmvW
bz8EnTvf+fP0ggzjOgZmIvEL+Nm4FvEWNtOCS0yOA5yh28Re/vrY+Ez9WNPBQktk
1JfITDSnthYIWmt6LPg3BrYydu5R2G0BHEVLkM15mkZbiPRgVUpOH07DyTjRZg90
VFXbn2YVonkm5pNgj0+n2cvlWNFoc3AdMryQg/KczVgm8shIrsoDFXPal7wuPqlJ
qFLz4YUm6N+D3C9PmipxNhSNy3HD1d29Mkds4lUfDZOvYv6+27MAArNvaE4HhYUF
j4AYs4Lp3ercNsOfjNfM6K9So4dr1MdeZQYgnoruZauINNfSSCzwC15V6SPmIYyl
on5eYv7wtGZbvCM1qEsdcDbe0qpC2lOmTZpy5miCqju/iqorJll4B/gafe2avSUZ
XidkQXSk7uS8bCprAYOP77K4fhGWd/yKHglJrQAV1epAx44mMDQbQrX5nseVM4ZR
0OnbsoGT80u1/SKJC5dJlKZYo6tmKWF17A5SPtw7h8CMJp9CscnCcIJCE5b6517F
0YzwypEPscK327c0rRFkP0cldX7QX5aQTz27KC/OAzNIAPidyC2XLvQMjL7r1t3D
d3xbwLiO3xUam5h+Q5kTyYS9bwXoeBTLKfXhnvQr1yg9DG8/4cwSh/ga56SlVZZT
87zT7y7GtGiBU1nYIY7Wf4BFPWlRR27DLzDUYD1YN0TiBlYW559PH0w6INZO1okQ
1QwTh5A8orHJJk9EmAly6/uHQrgdVqHi0oko833FwXggxT/1/mbGgSWCP+hfw1Ni
GROJHind59YaDa7HlHi+9OaCMBnbQmUCAuBLhrOP6RbFmuXm7xOUiPJ2MdIo9bpC
zHt1Ju61roeAG3Jdtw2uGhNU8Dnkf63FO6+j9Y87mG/LDgt1u4iptbSWpnq3AWi8
xNha792LONpgem4HQlLdGetdlRRM6fUV5j/oryyS+1cwR9LhF5ZcO15o0d1b3DJs
LDIaeJuJAbIDqEv97XVByMTrnoIrKQqJnFx2w5soUHjTKZlzc81jOIIiSySTOQUB
oFxA9lMotQ2J0Vjb5ZlSOp3KdSw4Ux02GaY7GoUidmXuzsQghguk+TOmwYQbJ0P8
PZvkzYQ1qiHFggFcNfXlrJPuQkIoCnAvSr3MX+ymoDtMbpAKLQf/7buxLC8g5aR4
TT0m8gfuzho3a1R5d/2fiRDu1zJvHXxvQ/UjYlZJBp4q+v888KJdPQN+WlTe59lh
7/rCtywDahMK/b28ZFCoP9FArWAmwX4TNO6Z1mAwT/4OKw2B3/tv2Cr9WR1HJyM+
+2LSBFQ6k4V2DXafnFYNINhzsoC77PRWwE5uzrrd+BgqUHPi2z0atc+lTQE+fmFz
AfkgZVh2sxQ0qcoWLAjqpw3WHLZP5DIHbQBXwPFR4iMRv7rNxZ3cWh6Ij91qClP5
e0nEXdETlpAjYTCk4v0mGNBV59cOObBNEuYJYFQFSUv1o8QtrNddutOXs16fiGVO
vXeU+C5j1EowaZcpdzvLyti0KoP00/W4pRSXnq/lFTlpa7/3ttFNJ2AWQdK/Xaia
o42cAlAEs9on6/JOv7D/VU/yEw/bcJWOnLMjuzPQQkx2f23wFKyFXH9tUIaFh1b0
qb3CBP1DSzeCe1zlDZbNq4if3KvMTsypiNbyWDDrSXMISG3Io2SnbV5XKCmqWtI0
f6ccnCBZpJx7fv84B7q8xqoeEeQ9uoiQtuLIaOl19jPEuE9X/TziDPnnJuv5u+6q
VBBy0oJxrrgOnIT4BnqlRFqT6HWWYtXzli7KYRrAiU3rsop/lcegCVmGRQ/y1D8k
gnuXexO8kyuNznf52KdsJDAWONayenVYgXXy3Aa69ZANbEJSu5Lp7M682qSWKKRN
ZlpqmfpN4Rdv2bavwc9KdTo8KBW6YRaJ09v9z9aGd4mO7QhqJlatH7zH9I5PCwIR
7b0gw2C2KQKNFggekvAlXcEsfcHg5F2Dz8xlCc93DfFxEz9EpziksbXf38I7c4jx
s3xc5Hi26bPDTUxF4n7onpMzHg4oJBDzBHwnxTLNxX+NaUNNqhQjGAhwIFzuTn5C
NE6WLUAz1MTsQ9f9pgTUORoFgHztObZMq1yl+BJhSxTDbQZ7ICHnZMpCHRS7std1
8elnCU3BLklWZWtPW4Bk5EJhSgrHZeIvCN18IKuKnmTsUioMTLWumM3XugLq9Oiq
re2NObTQvwNv6t0qRId942Z6g1ji2ZatxwNEc0YPpnpAJSJSZJmq95CwQAy5QuT3
i3aamuAGevtLtMrPdfb4oSq9Yq57Br3CBMZsDX5Je6VtFyYyKgPBdaEdTED66C36
4iYTY/ogfItkIn4MDMVatuy99HDr4PaEO96pN3f7G9YYUGZBnT9mkX8p33QGu2ak
aWWaXodVVV8eCiWHJnCwIq/80wBIHqq/nYqpSvc+vE/I1ZGOGonTxKM/AuXHz9k8
/eCwHxiW35xdsvEKCW0jsv8/eYcozaqwxE6oOKWBQ8LkuyVqH87Lz+ndVu0GgkLP
LT3Xs/BdFJID+YNu+rjq/atMlThmfJ21+2JkeQa2zs4x4RizAf+V1kyjOCv8ddqQ
0z78EWNRKmgnZz0TF3QJ7mshcuv7hGns+CCXoAno8GrT3IakJxPJIo+yuwlQX0os
aJVNPoNoADEC3mFqthA8L9ehsXGSZuI9zZLjKCkJMrihPfdUqTgnbGnAEjy8BKhp
AjBHwFBrn8n2Y97BM9qaRXZ1xEkaQbVwEMsUEr8SpW2T9NBlLdXJWgEkePaf3q+G
t6SSLakfp/y9s31BNrLmNO0O/YDyYKDPujyluxGP9y1l9D0OcqFG+jrzPefNqKCO
hb/WdEVjznnk2dg+tfcD4KSGb2c7JdSA4eowt61VjiOrUuQtOLvn3sHtoWhXvwSI
UA/J17y+1KXYcuWRet36OzUkJ0alHd5RV2L9VsmjORpYhYgsRXKy6RaVJlfEPZvR
WxWoloISX1diQKqqnDX87ijjG9aAxKGxvMmlbB69Wlpb7aE3jebM77EASzVmWFMu
ncO8OWpiikm6HsZBSsII6S8IQoRZd7DmJq8HMggKTnhLkmH6rDBvL2gqLr2ukkYF
qcFn1x6zXKX1e2q1aF0T+D5uKKplsmyivUFFlAOcu8cTqVAVlFuHeHCaKoKpsguT
hdtQV2Ni8VMorG5kWuBx3afe9d2KDm0t6U4ktiLbgUH+E3flrWzjq/X3P01nlXZl
JPu2361qeWNxFv+vflGZ2CGb3hGErmzh52NwDzDQQnZuRTM66B1LM3aRq4ojXMA1
eu4SS9vMI8cnZ8NtqVczK0TMeVijJtZljbRFpApG5sJgLZxyGTLBe2h5d51wyumy
IB822uzfXIbvtgEhr0geZf4G1JDaMns7irrUtByq4ZhHeQP006Ib21Hc8RMs+Poz
9Zq449vEjN/OI9gDXRFCxkfk5WvR7EUKUmhp16YUfqQaxkunF5aKStThGIZwst9T
2AfLLGr39ry3R+2F4Ctl+5Duprf+NKle4XD+umTh9t2ArfHnZ8ztAdx2jTNxxfVg
XcOJuR0awFtx2HhziRenYeMeV7g9V+gH/mnC/1Oh3kifOOrbsIOYyca0JkoVG5o5
mX/oLcwArphI901jIk9JlDoP0E9xw816izyPuvmRWhkTnyFt+fWH3OxA8DDhXXII
3/ckjVsuYlSaso7PjyIyaQsPnRBSkroJVHSQgiu7OanUL5I9ybeAdTHFnRGhgTn8
2s4+QedTt0kL+sSMhj45pE75LaDpKnpZhuH+qeZXTB7Br0JOiBKjddtkAchynMCt
WbXbVGbmp6DhKaq1j3G+8v6guxhgTslkH2q5GrjKxZNJxuiQ5rQdswqv/TEvfge4
SL2euLriz8R3Y2JtO6kR6xccUP5n8W/gDiTlmTaoVVNF/6hKC/bUEw7ECQAfr1jF
KyqsNJ+6OTNDMZD2dIk/76Hc+5YJNANfXyTQ7Hi4FTSV5dXorZfj6wlfnPgW2YOU
aw5DEcDtDXYo39ZiShV9q00BnMQnuTuCfm4hmS3NDfn5MulP8HR1kLiLlXDW2bQH
XHAACV5AjEQ0uvynDGpGexwwcfdF+i4QiVcCFG40IRHSxgi9sSCvMXkuT0bUZmE9
u6BPrl39onlz6NtuNwKjTmljYm0Lh5VjVj2S/dY14PEHC/giBro9dL1xzKVgtFQh
tBL4SwZ8nKtCSgP8tpinAI2aXJGjg/ixG0WSvuXBg78SJ70tSz/xHnCeLAmUcBz1
R/W2goZ+NRVR1Gwll09teeUQxB8eDdf3fpSZps2ucF3cOFElosIhwYmH7nIvzL/5
m7RSN6DdjrMkWMvjbo8t0kKnyAJQT8+jsxSZt0X8Kvh0cic93M4xBh1eZO2Y0aJ5
O2TJynhoa9nSv40XL5Kjx6emrHZLtsh8QW8Rtljy2806oDOmpQA7byJtYGfpBHo7
ilRNByWhxW34s0YU5MrSg8VyPmORuSw2UGSx87ZrP3Kcog1+gW8pHya/wtwG02+z
7SJSTILK13nwqpIA8Oz18SJlrsiNATXlayrxfYHagd3905nzzD7GMK2wL0XRhwWF
xqvKJNqERnKkzAGLbsgdDKYZZtghYsLwr7pTa2eUt6INL496JzNX0c0IhVIBiH5Z
+MiEGEGfFUGc5UK13PzEfzLVDxEd/TqTUvNR9fRSF1p9SwEK0/pJqkb/yXaAv6hc
uuxFItzJfFg0i92CFxSwp45NPy+I/y0hJOLLNrUASRvyAMwOznKdPRSZmu4qmL2p
+l3Brid81ZEOxlct7y5wl6FSK4ZeXep7i9trz3XKpzwJ2yH19tN4JAP8jyf9UzX4
I1P/cpGqI49MzcDbje4GjM5bFkW1pypxDSLPqa0JMHFGJO+hGTQkItLmXvdoVkqG
XW8VEXlsPZomdXAniryLBZ1HGNZ82Dca+8XB3fT0G/5R/dQfWC9Yk6HdNqVPJptN
BZ8N8OuUFbnIBXmJCyRM4KN2TjzF5PLn4CNnFEDYbu6ZANnSNIk/QmCIDpOQ+E/X
w7A0SSEvghgtlEuFZ0Kl3eewdtLsnmrEUr8LPvR9Mm3nigAG4BbBCOG9jcRaBPr6
G47XNoysEpOWVJVYbMaCKTtY/wE+eTpaa7HpDr2vt4spE+fKCDg8sv+vJN5jXMjg
bd/S1LsM9CdzYWy34pIWXFDmbmuBhYd0Q8wFJLgiblxqaoybWLYUnMZKy7FT3Wk8
mjrqg8DrfRIBuybfLBaA0sLXQHYHdKqJxQ20noIpXZF5UQsIeIfZ1z7OzobY/MLe
RMft+kRlPNF2yU8xFeo6MXYh0lvEMBJL0xtrHnEYzt+TxnDM9sQYI/oROwX/+YKP
2PnTBx1cec4G35Z9dkxdcy3He6CjCv+2NzpVz81Lu4bjQmoN5fevaKYj+XBsul9P
7UHEmoWD7Z+M9ccBvJnUZeP6THV/cLHfRLp8GzgtF2I05lA9OcB3Bu7mltwHU/IQ
CWjHPXIV8WUVGphTssKDAE+RHTDsgF1QO9Fy22qQPn5QfWiqRq+MdzmLMrk3T4BT
I/ju+gWHNTeZCoDt2xr+maMMaj3y0ZAFZnNFwMk6YzWwOL5/52GaHFRJlGQuC4Q/
9X+39t6OkiINxpL6im4NJoKsVntnVhMsrILHStG+rFi/bvMQFVQ80Z7rbE1Wnrrb
ttnK08rZmpA9jRPiOBExRHjk4en5l3+N7tuzz3llsmNYE+qc1eGVU3NeCU/Vu12+
DLWIKN9UU+HdQxIslZUNY+kMu69O4TbHbiGvt8yeB4zS/OMRBdhDEyamA4IkaPAC
8NlnFEBRE5KODLrYncflSNVEXiI6QtaNAuFwfT/mtzhEHALk+VVJOXi9g0L1njdk
epmUlshpTG75CDluo75IJzMrSenCTEe5fAZ8C4xM5y32zETF6I0LmbwUJNIouNqH
9QQHO3ivIgaRcZCuD93qInPK12iQrpjO+8PpVrkNc6uNEzl5rkCKYCyljt4imRdm
jTT9i/Qw6uPndKzEWPKwIVgUMTrCzakdaogIU2svxt2qrZtYal/MgGU1EhvztAXm
+KwL2pZLEpfxl+cdV1vgSbteQp/taaA+k+kb3+8u44aD7XNde7/XwkbfNoGLTjcA
L7lxvaP6WUy9Yx1+Gze5hXxFX3TBbvrcCZd8rJtreBYOYOUlvhCn8x7q9ZwBkIk4
F7qn0Xk76y3hBchz6qqphchWj0F+QGjnw6lz3CFWV6184fWoW1vsJWMB6jjLXMU5
d5vyNnHx0kd9FgRkjs2xQdHdzBopyPAC+WxKK8229tWWvTJe1d+1Rk0CD/QNQrQM
QS1j81Y+1T6N2flkT1QZZvgHRhshhfFoRzl1CITbSLeXAx3KzEZmItMY4YV2Z5cl
qEjMQPWzVNVCPX90JOQQRnw2XrdB0OixnaPxr2uk+lcjlODdONhrRmMF7v2dVXVS
uTWGKmDNogVlDVHvYBSBtkBLsS7r3Yrmv4BkOU6qFyz6MAysDHjqLfJGLDKpv4hY
MgbeIPxUQPXOkzIZ/4K1nfIVPBW2KB2f+ZH3LBzm3kLHvm483Oy3Q4FJwtwMZPhv
HlUMlBFqVultYoYDtozr/yG8FflNi7gsecxck27I885Lreq2F4gV7f2BcVCoh0o/
KEQc8zZi1IVm6o+PD6w9EbjDKAy7sAtHOt+S1q8fKpktBgFaLqDeFyJyL68G2p5t
Oa2ujszxLFxNnv8ykvkfTy+qMrqKH9F9+1LnUUSjjsvXfH/jebP0FS6h5DRXhc8J
Ekba1Rr/tiMDiku6Qzm7/6sOwkOMDpQ01DYaXnQBn9s/JYq1fk5gglXQRvrnIcwd
cRfM7/ukHBQhaiQehm24/XmR6QC3mDJPHi1Ccqhvo1YYJB/oKURFrTBSb6XK1ywL
NOjGSBUjUp09IdLRpr29pgCJE3U1zcKbAL4IvlhmZC6iek11Q+2G7BLSnAikxghD
tBaCmDf0vbJ+RGayhUdfbc2evwOe/9u5yd74jOGNnazsbIx5t69jQhp1sCvhxbDS
/FOC6wQheX4kT/IaO5UpXvMFyT/Vx55TTOGnrM7kcheTkUntmtaTyc668e8qs+Au
qwUQeqOstGJnPXIimieXR7ZKUp2GmUvw7/Gb2MoOId02R6/NV4xYGKtRSChQ9FHy
JbRbizhPzg1uIPvmsHLCoXFnhdvhWE0d/byIgXhdkMjkeMYZBHSi9Mw2gweMWL4S
s7kYsAIT5N2XSwkliorlHH/TsDCXnNiXfd8QxXr8rc6LZbZevPKABud7opH6yt6E
4KVAWfDPCN0mZmBlG3mYxDSuUxc7Up0IlPy4Q3weWMcISXU/OwqpftxnCSSH3vZC
IQ9wa9mnGcuoPxHkv7H5qwSw6ZJkZFxrlvB274vzKNv4lOIcnX2dGRm4ej3W5MnM
fwaieYXKqoJ8AymHxIT2r16CNi2rSQ4Ha55bFUWvzq0UeZy0Qrwd62FOP3/+fg6Z
lubufRF6dH06y3MZd+xfhuomXs2hZLMK2UdGl/ki6BYgsrZvXYT4m7JKS/AfysLu
CvhnkhteXPXqksM38IVxYBWbQQdMQaDOZef6GW061bvGaVl1fU62+Jm6gOCG0edQ
K4GoyC4zZcrYE+i+070k9oTFm8syzwWguJlBZEoQjsFxA0iq8lrJTKMM7GxxninU
KprLvVDnEXHYCS1Ke+ErQWmAubBvMoW4dfXaI/5exyQVlCkFcW2cLq2LIwGzXEjZ
CU+K6c9ujET7BOTkZLO3hwNghZeBopRT4eWUaxtAKQzV51nmh/9BOsc1AZEd3OMr
LE/xLfx/ySg6x1C92tKqHc7Pz0CIkG4Zwc/o5tUutvONnIVIpis67oPXRD2wo0LK
l4JUsXupqXui+3yh2VeZKMYi9OzLxF6Ejma1dCoVBLqZ0ZZ1wXDV4gJi7ix/GmFY
654L4NfthNz9wV2AxydCCL0rNxgQu9p7ZtUnuJJwINCYuM8mfmXoKzUoGQIp6DtE
tSK8qP1hJK2n1OfkyxD1sOCk/LTtLURQlk0+c3GqCOX4fNMdmF03A4TSQL4VBMEf
6PX1VqIe9MISF62isa1ZaV+X/Lypt7FDkFh9e+B+hQDFsE4QbwDu89KVP4TfjJ0E
tt+c2MarRN0rEHJ4i8SxVi43bm1I2X8X5zYIVw+SAhct+BygaoDA/x4O+viUg8jq
0gM5oeU6IUn10zeieeSHQpgEqWdC1hGFqURiftB3ecmX0Jl71d/L3BdT/KKJSFtx
u3l69IccjW0H5yHbqpAvZutDIR6dU+auEFZ83gYNTWvQWVoBIwhY/riqf/sdjQUE
s27nPt2T+0CP+qNoEc+sNW/M1u8QNORvq+kSGy0RsjTDxxRKxRMETKuQZnc01qWN
Xg7uhcxNDzYHP9vBRC+jU5crTC7qYyjfIy1flqor4tnLYcXlJJj5akjKO3rJvxNB
l/7jUz18xdRJYN9eqeL37A2HmrH3SToqTRUBYBy9mTKrKTPaoK8ikCyA6oboga6w
f4SP0X/t/f/sgZXRu/gXK7LUwsUHT6743cgLzZi2RAkqps7lnITWBUx0oRILP9U3
cdkAzwZs6P/LcCWbuXLm2uWyWLgdMj6hJetvPpZy1ilREbbGeDKvxf8CvBJV5diV
h9eaCJfPaEq7TQ88gLIv1CmR2glugMROJEFiBBd9yfp7+TVAFq+YvLVCpt6svRpi
wCPI7CpQKpC6IxVKS6uYrKl4Rfz+39J05Yatl+M1O2K9v/9lDG3FzSxTaBGF7R0v
uVqkf23lRcBlkR+fKBbDj+E++f3gVi8vu0m8nQKNuhLtfiqfytBA7LOnTZrWSnd/
HKjiuvhetvSy8YhNM+7s25BUCN2kjYzsX51BC1Lsz1h97ct/0Ns7QHKz9V1M6Jtp
oWEJ23rJLkQggYj6bmdwAaHxFE5Gip9KdpcVhYTSuSMzbzjRATUkFKCswNfjIOuZ
ysVLAh2gbm6Q/RKGqow7YDgQpzDvSIjxDogLcKrHlhmS+rTxIu7NT8bzYwqJsmM5
UpodjQ3lsHIBzXVWB49DDyAHinwtJ3wByFK88B4WRlFlJ82GU87jyGajYIJtwXr8
hiD9selALNkpGuijgEM5Awq0VcOxA1tZixwEY+za4gvnc+NRqgeQ3CswV2WLxlv/
aOOMHCkYxgFu/ZedXNsoIIR6wUGPdXlpvZRQg0o8/gqWpqxJUs+OJzdI2ZDhgviS
/61MvT4N0s+6pa+1/BpswYZtNmKpfaJcOGcHOCSQ03lMDv/vftAoNvc8SqTnXleR
dVMMmiwdK158SWundhoFuZKrEuHB+soxDcZXbLeS74uI9MpVzs5lob9J0kMorGwH
arQyjHtRlbBPHXWMXHZ3Tq1cmVhiKKRnHb9cKG3w/b3SGjmcFcqfASyfoWo2BJ6k
hCtBoq5TpgQT2xyKUsUrEp35+sKYymFU3VCdDlxrs1BqYyv6nCOkPApcvfgM65G2
Y/hAN9H8Guatz10bnOCfjErGwSO467o5tQzvlHfXHQeBa4/Gl5raTbhHjlUrdNNA
8vfPkqO5NxsY6ECkcc/WqudNJ8Npfyp2VGKk1KyzIrap4/107JCIwd384+IVYfWM
w4lQmnIXHAxZEoNmlX08j4+Pzp/c7N1q9/77D9AsJI3YWtQyschq44BrPTQn9RRf
gXztF5jbLaStVTNTqsIkTOmedUL2dlk3DWsM+OLXeytfCr3cuAQizaqlYhXikJMP
uZuvasz08FrfOIotM64xp3sBclu9/YiR6Rm/Exdw3cr39J/FHKL93UJNyaYVUwg3
fKarVHhVnwgJHml3t08H89NkWfINrijh0EAKMH12J1omHzSKKmm9vz9opy4LuZfo
laprKWByOShNx9hangZncmUQ/VwdYjNN+kIu9+Gg8r0PjuBDe348UBgWV6Vy+xET
89nVvHT3Pv/uYJ8Q/rjjmjxY92AA9fzDtaj5qaYFKs0b3xZyQq2l/KcBDBxESubG
AD1ODoJVIAoJNdaShYZH3mfjUBF9XcpWJbmcwY5O4mPeeFUAM9ZDO6L68iXC063+
t62sKNFFpr4LlSNBgceTzPzaKpksU/uyHpD89Qr3kwHhO156QHcLF3Q1vmYEGpah
VbnLJ34QY9BlNhmUzlEAHRa1ftLNjJoRr0WglLnCGv9Xoxqvnqir8eiI0mxFEZKM
7IJhZMMi3prXA3XudUrTbKdAR7h4QjMO1cixtmFvf1m7apedP3u5D+ZGg3uPsZuB
1HZ952ne7ZTY45mlmptdArusV3AoNyz8FYdwNMtux+Mxj+7B3uKBaQDbOO5QGqmg
27JKe93wQEVwWXymv+j2gC6JNAa/ofjwdQsoSd1whWQuIj20sB8tvVaHqXo6oyp5
3nabOlfwzVvRr6xOxnxOlkWopV2Y/YSrpNUDVCw2BiNo3VgdXTCnDuIwwuDco8uk
9ObG4wpgJjglFCJpEBl6jsPrk3cJuGWEkQY5i6lV71cBh3uaFuD34IiHMC3b4QDs
R0r7ilKjCzIMIuPVfPNqin07EEeTg+gGv9GBk/fuSkJA3FWhCKKzIcban3mUPdRK
viiHF0wyw3ezXZOvxgjSnhvcjQsvAJ4ZLv0jVIo+qs6zVwnGk+Drh6xyc7emqC8a
9KwmE8wQEI5diVnmLbEzpK8k/qD7O8zwLJ96EtJFx/CndlnUDTZp8KUvwTPPg/ry
ycqv1cqwT3wq6Tw4ykqvmQ139HzCtAbW8K6yBbPObKfe3uV2Y4ZL5vJOjUunLj7X
OiNhG02NGH7roFKzZkzBcfxmrxhjracQdSAN1L2AHABUOVCjDPG9Rmjglm7UJc3h
YPcgUa9/5W1ymDK9GULbq0CBaIQMtawdQRciYCO5L48H3H+Xs2pQJCyMiPZKILtG
C1X9y306BVkq92R5Y41P9Q84HaZuYgBIJRn/EmVOa4E4CCUB/MEbkAKf7cuPfdAQ
wEenXoustg7Qislc7E3x9pNB68VDZvDoER1iKQzBCGDrTI2jm2h/uHMc5N3XZWCu
yAcuftgNb03vyzIkvNS8wbnHNA/p2g9ULdhFHuw866+Gyu+CMS5IrT+0CmMIxPtR
o+LW8cXnOwc76z9JyfQyjaEUBzbBUSpkPCEU7IFb+YkQv/Wqkv6R6LDzAjh39rIz
h0a+R5bq1ITDa3O9I1yBLtmZ8KYE2eXfq+5GDKN66lKiHyVM7qBKoi2K0KCUEEOe
dHGobc0/eeTYpLuf4VFS6gOeHD9mc/qHh9EL/8n7Fu6WZVWESy5DqUBE1Azd0ihm
SqsSih3mF2fHOvCtkAY6FQC3OJAiSw9pvBK/IdmUsAhxQFW3SOQrLBd69K4DIfw8
h7QCD75AV2bqgmbei6QIjhOukxzPA0/v9hBOLHtXiuSxNwDIehcFsiA6E+2agMlx
cQmuNr8Q3DHP0/fM/frr5GppF0p/o0b0SPDuCatVUBg9cTYzyAKqwpFX4TZBbwrx
7v/Q36SCdPn0wJVLZjOzmrZtJut04IQnCDVhY02YtucbQ4/nUIA8oI86y9++xjc6
EkukPscWKQKsj0K5MKczFOX5IhjhL19pWFgX95arHMJkQAgjxqAshbJClviM+VdH
N7KqpW0DF33/EslVwPaEjCGn0p+cnfM+zyGOvpdvt2XMcCj4VY9RrjfosfRu6pQ/
cxbEj54z7gyzar4xeXz7e7bmxx3Zj7kH1py9AiUapd53DnjHglIftv65vKa5g9Qc
WZie30+aqeWKyNAhoOsUygt4h2y3N7ZUAqdTheSlzA5ujDz+bJumLE14Yy+mdJjT
VM5HgtQWzmukCBrU0AqAdUjAaHktBZXUg/HljZkBZSvlYm4iR+qe6D05y/O9HcUz
Y3xf1KIFCQ3Yqsdv78U6AIF8i+0JDx/tWJfbo6tsriOZ0Xg3oppewV74Vmz/YELY
RUfWU7swdX0RK7aMDlTY6VtigQ577j0WH3e2MxQEEzpgZWJj91AGaJC/qyhEq/OM
JHAAOKm1zlNRR/ZGHajDPy1hCyepZ+kzhZiLX6H88nNgmD5eWXOD/xa3JPaDpPyE
cbDl6X3qRctCuX/JHhhMjzfyxNkcYWG+KWmyQX8cVrMi5Klw9zvuHHWwBG1ZM9Ra
L19gPtpgyOiKeYnz9L4kga9SIQz+oOVxTZn8RdOkt3RKBgJ6FPrmeUXpX/mtdd55
Fa8mR9yFv0rHkgd0cam4/+26vAVn6H1Z6fllsIDvIdwoKmENk5YkL9T1xaQwZe/j
jNgLXdy6GxEzh+bPhJQsB6f2Phg1Hk4QkpjCxXDRdYbBvN7TZi1rR5PtYglE3ahy
69egOLpWthioQHi85Vy6pHx4y87RvmRO17RKdKNxGMLmWIp1OI8IqQMFKPdq916j
fEQe5PCES9mH4iAjYSBt2kgs12lCcxOocy425dnD3fE6PvFNaFN04Ls1mL8z/sae
AEudIkAO2JX4Ih/oVv1VksY1Z7eKPkA1tlSeuh/r5SsS1mjFq4GxdSZN85dlYKDg
LmbjMxOrpl3lIfLoDHsf/hQytNAMl3rGCbPaMR8BkXo4NRG0EQTz25+fkv1tABf8
zdBFG6oa4KiZZOXeO66fM1jciR7Xs4Vb0Bt8akFsF6qxWlbl0FjB15FVUn/e6FpD
Pd1w+NYLNoR16fuR20iV4sNs2eFh8SRhgxpmZrp8TtA4lW+ar5m1woRMlJ3o6OhB
OSCcpFuOrZfS1hlLpcRjlOgbLGL3tGSfaESYkqdZMDBPgYJOV02EIs5W2DCkBStX
VznDuJZYIGFGG3UpZibhWlZ7g5uuhdF0pNhSCu/SlSPMoU8K1yxQne6lO7Mg3nzf
um5JjqcO4bkKsivgFOdrPG1rrXJ03NtkA4R6/4S5ZldTC8iC5peJomd8ZoRvKl50
hO9qXNlMpNt/mNxSQoyWpag/vfIIkqMoNlHBDKyyynKma0SvdgmJ5lXwZVzLRBtq
dRKSHVIQWG149h+8Rk0v3yqUjJM2m4NcsFJt/+iQlJoteC/V/KWtBxYznubbgTeO
EHzn07cd2O0dFGRJ0x4ywXiITVXfmIWxvVzle/r+9Qz2Z0cM0lAXPVdDh4+Xjp21
a/kyZlwLBpU75fA92NKxobL7J+PmXiKF0cKIEWzvYjpMUkXh99To2/JHdfQ39hji
ZodyKhBwtdfOsYxEsPGN1jvBaH5bc7rBDsvufg+d9AHINdDhATMyqfz/ax2PWBSK
3KEYeLyCS/spDmfg4W6pB3482RoIDDgAkLIJtvKlHti5W7hI3nhnXO/ZNroKYjSa
DJwSeXYDtWWTX6pWONuroFd6QQaczd28yo5ewa2RqyDjzzFlX3zhGxUoL0tGG2cW
aESOFwyAjw19nYKPo2eqwjSRh+xneTI/M8SmXFo9wXc7SPlv7ocO7KNqxY5+jKTX
IDQtGxBXZytPPWuz3/EkhKxQ7nJqBwAc/4P9qBuAZVpXfiKjaQAUEBbjJ1jUtU8T
t+i6DmzdzqrjnMjCdOtXr7xc/tqGZPfzuu5klybaUYdfatS9+Vsx6jrNN7/znrr4
v5NRuQbzCWEzLoIdOoaKP1yeAcMHdxZ4fnH1hcT4M36BbknqLl7r5JsevYTZeRb+
l5Sp2s8S4oz3raUpVOGbObEgCiB9fuSsWw58h0+tkVtJLbz9SOysRVP7Wrfmr2KI
Uy7pP0oZEBjq7hykda4n+zHmiEfso+RmnnsSzmaMOiN8qgCKTpDv5mArpXiRwM3N
1h/NnC9HaZXZ/Z2HkvpDWmKJkKACEXrXcnydjLhM/KVXXL+5fLmmEM5lmLsBiaGW
BnCH5K6TRXN2jwVYUQg4VNfZle0VCr/n9J75IN0lE9j+cm56UhIfP975+vmUqb1c
phGFUFzEHlAZQafA5QZ6uMo9dw7in6qy3zl+tL0rBy7QBFIObqw8qbR+uyA+4OyE
4sp6Z3xy4nILOv2Az2Lvr42uxBFOMcbp5UNa6Xgs9sheE4qRmiPyQ98ue+x95k51
lXKw1epVfJIoN9SDiEAT/98XtRRhtsOUkN3yuS7Kt73HGP+K99n0wuR+Nzdz4hVr
YU0kfb1AKt0IWCOgo0Avx5LSKariJfxsqpeGh5Hy4RgblzwJnxANAi9yMbsH+k5B
ihHNxpfkL8QaYjXR/doKA7uDZ2gMk5uNjoSoqolQpKm/pnmwssJ+MgKITnSxYtCU
dlH3pHztM5g67UJDKia2Zbmt8MnGkwM7PRfS+be7grWyzT7D9FQqoMu9li//nesC
AM8jF1b4E4Mqo19g8mbu/0QyhSC6m+9gAodZO2lpS+02nTVL4Lo60DdWwcwnhz4g
JQQZEOeAYDUCqPKzLoGVYksDO1NEWynHfnNoakLl9HREGpJzgfWhV5WnEg8dWRP6
X7BOhWZTXTPJtY4o/ZsjEuFt3yJe3Ax1D986AniegXSL0nSA052wV33ayj2R7quD
EdEyHCW9oFgw+yRZ37R+YA3mjEzMwbka0kXruBjBAeT/M5aUNr1r67OvXdTO7M9f
f4qrXpx5ms5XvGP5gNz3a35f5DpPRtYdF+KNeFWv4X0Q7JQTQrNn6jpR5WymTgeJ
u/O+HHkwUAm7iO6WXA4cKgR0JliAYlJglPjuGt/n+HChvMZIQxpSX5QxbBGpRrEm
X0lwVREccblEUuPuY7IE9rhUy3t/82LbIVQxlfh4r7TrwjZaQIhPGwcjxAh8hNwJ
ClbLm8fUbVh5f9PgOp+2vOa2wAafCU8O1EZ5kPS1DfyIkF/WM+tIFxKbshdIahDq
hzAyx1XutpelNtUns3y0kYZdGsL4bIO5RglzZxbTCOkYyuQWplQE0L06SoeSV/b8
cOwSAB3BQwo34tFcFYwD3wdpsvIIUCmIA04smr1r58n3x6sangjk3pkwkg2bqe+y
29ZRyayDyv1KmFQ183V+jOq5Moc9rzSiZcO90GXOlQm1Wh+60D88pJAW0tzpuOWS
q1jtlDS+YRFyio+b5egEZ262CkEgnBkxpVWVjywyk9PZ55NSG3a+6v/lMqg4FQ8c
f2hYIdSHJ13zXnqBwHy86pMC9AMyhN6bTNIk9l/twReVxSoRf/NyQozyV2MiDSOk
K6bZe3LREUUywoQBDB0IsOLCi0Wm78tqGmIQFg6IBCiidZifuqn8r1OvgHiWyNhh
DnllrOIL7P4aW7MGWOZBe28+ZQo25VN+DLZ6IrND1tTGyJmcO72o6FiVtHosS5RY
AL98S6ewTCSShrq38+6ih19WU63D9dhoOZ6Ls5y/jwfm7hBGZuo9bU74zBOpU6Fg
K9/6HbtuHNaDZfWs/uLIDB40mh3RgmHziz6TG+YxnIM2iLIy7vFBoXBA2N4INofI
z0ZpqiX066ihxBxu3xjmGNAycN21Ze2wlhezpWBd0esP9bUcbOyMV/OIcxbue/0c
oj2Ltqi1JvxCAx/e2qBdvbowzrkq2GmN3GIJ98/BzyE0k+lVxC/uO6yleIv/974a
DUr52pFJeRbPCC2DPtMx7o6Ej1dOJQrQ4M6upvC+3aZKX+TR58B4eOjYpXgb8z+7
bNI06eN6c6dxl/iEW3ywv1s+SSfAoFDTr5i3K2pMZw76rG4xLF9w3fjBsMNUBmMo
3wGNkk90Zeq9yLFLBRKbr38VOjE5BbPsut2tvuDpkS3Wp/E1lxw5IhCxNYU2Gcmt
DAfVScM5vQg4a8gd2uDgNedum8jGGnCfJSN9P1S8oA166Cd6U5tyXaf19NUvdK7P
BfYHvyjNrM2Qr+OhxkjBLKv4du79PFwRbPMaDF+oqPOBKfQfD/kvqD1uBXn2zNZS
jXrvx0l/ZcCeUGbzf/aJ1Kq99Oup/+lQFPpjpUikXZkBbijEv0nW62p3ULFY7TVB
IOPtQZQx5Pvi/nufloQkFUXhYqCq/kz80uq5v8gT0rhkBwfv2LQJAurFu2crOawg
BOvnlaFJsAovMqI+Q73/EGYF1wF2gt1iwF40VmzXLofTWleqX0W/TROFlON64sMW
8IXFWruRk+nFYfkzHrV3eSOPqk2mlIvuKPmlttVDK3uZslkzMPYTxCGW0MSlh0S0
IxytnE6jU6jxJ+F9ADUL/D2A2nBz0xZX4nLlF3QDHkG4fB75EAZ9hU9YaIyUFdfN
3S2NgJgq4J4tDZIJDpngu5L2RGyxYMMeazCQjx0qSJsQ7PXlh0I7SuINbAFAavrV
Py3HcxPFtq6mzyaY+3WoVOaxszDKxqnePsb/YrxuzWwywFrOLSg4FirkDbulqB4N
1vWHi87y05GrELoK0TI1rvi6tD8xM3T1i1fdpEO6BH8UfF+chL1GJoasfel9qqvV
Ak1GQuYPe6VwX+iGqBhS7xEu4MHlJ01Vpbq2jfdC5jkvkqRIfBWBu43eqBDSI2wP
2G7JHGR1KSFgU6b+yr1x3/R/jJuO8ahwtQVVIOQpEXwZrluEeHUyoIt5j+hYponH
SKst0+g2WaE9CAJhMOXXWCAenaDW9e4n5OgJ1LOhSmKetpvVfaA5y/1rBeNIUZmo
sU1Fse21YK/JOifSAsNvJ5htxt2CHUux8d/lnU+ol4G7LTxaP6HsW1FyqjxD9g5m
5PB2mxYo9NNzJk0x6hOvHOfoY+zr0eUrb/hrUlSJwrR1FQ3wqLWTsO15uBB3GQij
VLsSOWD4R8NpAhWashEcUEo04j4uGpAM2VRDINgDpXl6GlnfK5suzha6I4wkzCeC
MpFdOumif3zfzDa6Hsugsxug7QqMA/vPqbN8tL1FG1cZ6+/DsynZOYzYRcwQChcc
ml+UuNqCj1MN6f6lJBLXqCr6246QrzXln1sz6pFyaxdoWhL2u3wnW1wrzu2Hkd/a
KQSBawhCVRDsoKkySuGTircXFUG0T4LAp2OOtU5XvMVWOVg6vPCAL0OyZZ63gd8s
xZ1fQW9I3OPLfcox8EB+gfpKQjW/ZjGmj0LKsi0LgZ6BJarD2bi2mUUCVYZn5IWj
vNAptVvGhpG/NyjeoZ5nH0iXOu5NImdXLd25siTf23UabktH6hS4W5D5Q9GhQp4g
4My4+2sEHSSZdbagiz0qpWrw4u4ZSC9pNLC791yUyjLf2ZiWUeLCa7zO2m+6Mg/6
NPI4fPBEo5XZvsqAP34pP3NX4hAn2I7OJNfpqD36qHgvSbUYOOgVKNkODLR4VBzW
Vsxo3sXfJbg2ojCCrKwBpnjfJzDdmOeVsbUudV/liHyk8rajecr1e/k/VH0cxzCZ
O19KyPCGjM23cxw9xa0+Z3NUcW5JUNpeEnQT9e0McEDy453U0vQ2qreJJdU2ttqB
wdGFMbwjpBxDBfSmivBBbZnt5x558IrIwOi8Ak90f7X7ZlgsvNFXLWX2IZqVKKGf
FaUEPuHhYMolJOmRxUcn7qtZ2hzEIORu7GIyPrQHZsmTJoznd+RpQ9YNvxHoXxgY
Xt5Quq7iusD1SnGaAOtkgp0ykQJEfLRPG1wA/hRHb3eY6/atb9bkIDsXF90eV34g
s3iZzeTtxW1ARdwt0SU3F3Wy1jMY6sUfs2bP1sO3VeVs/lMGNMT4C0l1AeruQGFI
25rP4+vfvAUgVXklrBgo+b6F+EOz+fMnwbuVXkMvAKAVq2nYdAEwUrcJf6FQ3QS5
Pd7qh1fWOecer1kFR8b+a8c01x7lSGUnsyM7Jr28rt9kenyF7eVhdCzx/copHpf+
kamjB3Burj8kZDDdE1QZmOXnAQ4y1OyjnD4F0OLdMpQ6175iQXjFPQ46NYuBg9qE
wdRUIC62COwA7IUhGy/UvktnZC7PjO/I5iwQaPgeKHAaqS3jyJmN0fugJ7HSrnst
2FU92xuDthLSZrlXzRXBZAi7kLKSQ0/kZpmySVq3q83nP9mDnMOcPgpFcSEKDrrl
567eCbgKmDCVPTe0kcxteUQkPPiSVZq2lie5pX1Gv02Pp6ntOuTtVDlUFBf/Fkkj
aw1Pb3jz+8bKBrVHEMX9r2bfWRTbxZcPTUEs+VjD4Z+wgexWl89cvJcrlZ6d7eOH
MLpdNKeSpime0J0EsOohTChkgSJ+UbEsTrgegL925qXzni33Pfn2DXAyc3VD70hi
MlC3ACOP6xuIE8meSk9MeUO11ZhmXLXiIu2p6sG4zSXAS91I9yVBmZAafoYcMw5K
ktt1OiHS/xkYu9VrRGMJfZU5ZULBifcV5RxLpqYm8cd6tA6PYYU2CiZy7RhR20iy
QXMuR7DjGJRTc9w9bPOLPyT94h9KUpXR3jcOwYLXLset2BhAc7T7qlFdgB4WIRIE
P2t3NMY25JRsQYvyDUwovpcsFv8ef7mmnBImeCMz+dZJbM0fnTRapCY9YiuhToin
0C0niRZsF3gUAgxU3m3IViNfLJ25SGB1djEl39+9D32dbU/+D5OEsqYkgtiOHlRp
NqcpTwBZ03H76Jcog2ZAlTNOLdngGRG1UgaqDyBimck1S5jS3gMcOXQId8q995ZS
shySwqvDkI/DU6QJ0in03F+cbmO8SgNCIbQkp9KhgojxlQ3b7WbJeBq1s6SML2sv
zeWuDR/lAR2+jmPeTa76V5Yo+4APoRx5Y8Ka2Jo90FwfyZQ8FyIZ8VKLbRibmnOB
TYgM0vsaDEzqncxHJTn+jlQXQLjjPWQvrvz3lgxihGN8bJjxEdMN2I9UdOsvMoQ5
Gzd5inWHt40QbjQP+rWylt71cQTNLsYY9T98hLbT6D75Zi6k9wwuV8V3kd10PaXM
IwZYZ3rnTla3qQ9TBYnBEu6Gt9nOcI8ciQffK2MwUY87lRGpDu6zGEQOvrwqZ7Z+
np4c/RhKiyYJQQrT3L0dXtt9gO6gJJJYQs5AhUyUrDsWqgPo0GI3YssMDBRgZbBK
0jpSSTmvCHABpJA8BpE5h8TRf5N0d59wUmsQ087CMwAJoGqjrUsfjQQx842Bs00A
pGN5kyHBkxaa9QT0dJ7VL7bvk9Jt6IGrPDzPNil+vxvPY4E0UCgbrgVJs5wP7z30
b+8NxjeS9ziGtRMUyjAZY5WnllRq16kn6Mee85j/VPBvDDGV1IgC6PU8MsE8C61J
L4SxEGW4JPM0DL6ptv1TjKfjM2m6G1Io1r+rvhe6OnTox42Uf7jH6skeDMOuz6OE
+GrHfr4k6p5Gnn91f5DhqTqbn72xKUBsHGP4R8Q3KXYjNN45aBMYk9GJvuf3Nwm3
qw7l9ugaMH8AcWMu5eMek25bXBjzqqZWcOM9QpkQdL3J1qdL5k0L+nHpxW2Gi62x
44xor/e6t80UEyW4igr1Rw4c2EeMHccDzs5wALMmPOnu9WXNNsDYtekUdkDP6nk+
seCMQvCjj6rs809i7abtDi1IJkDvPx2g0HhbO76z2NGEYPcvTVs5PgZiF1lPHXho
2OsC9OCekiBrhQs6slZLmIiJ03bGLeptLpr4SHdCydM++LR+yTndif1nn5u9edH9
rVp31oy/AngSZG+PBXzgCVVPsBofgefGQV5q9DDF3jI2vOMSG4ibxIEFR3dwqhT0
ihWIJPwEaoxcz5XvRO77jYsjkey6PpDgJx+LqCvCKX2EMIQrYng57osYix5Mlc1t
xG/OtGWUdNdQRVPcvHIrBbBD8JF94/FntWwvj/cB0FYbsJ+H6VAlybywGJOBmY1k
RxzUt6tVrLgXQkXUTI+PuhmrpWLDuqrMaTrlFnEG7dd56sz9hJA7efrfR+4vBlAo
yXhzM+kEzAn0NKGAKwfXuzoNU9HDD/N/5hoLejxY5bF8Vw7Ntch2XE/6+B/OijOh
/TH6MKiDdiGrS38n4jWEBL/u80BgOxO6H+SV3DZnNPFesWODxnUkbXtw2R6CrK8k
cwlge9+5HoTfe1dv2fUTnijuE6laS3qORy9ZtpfQMA2O5+mx2HECE4p/+Vv6DaBT
EByIIxqdCXi4P7p578VZPv2lCpBpDEC1oPb3quViNUszQUkmK7wVwnZqAVyG3OBx
69far8ML47yeQ+sUUnWhbR+nNl2KpZRMFe8WfoaeiqsiXsvrUexRvu6yViLQcCiJ
wH4UL8NLUmtv0euvaHHOW8Zi+mQ5IzP6HIAu+O+EfWpSH0q5TkHzJbW1nzMRKgQd
+Gz08dCGQ8c2qFDB8A+eIBJ/9SfZg4CGyQg5CrdAYjjpM2tGXSR0KGd+KOaM/UD8
153jo6Y2sq0tbofFKlUp6xDw0wVr/lnx7hHZ1csztRNggyQZ5uIrKm9SNOuc04we
cXx3VaTSi747TMFmMkO+6LRUuVmwQiiNDxiwSU3pNUYTGTUdL0HdKMzdFFFYST6z
VLwEYIoZj770MjPpAcuNjV8nhFe+VBfnHSnEP+fVsxcDSa6vd5sGEc1m0tHEO4As
klzsqSz0qygrmgDz3nWoTqtkfRxSrMbPEXuww6Hr3M1+ShON8usFVyid/+EBi8t6
qHqli4nRJrWssjsH14Z6kKO8v0jq2oANdxSVSroSf1F9VMSxaZmyLkN5PYeM2m+h
MFRrEm9g1ynuAODY4IRs+kJ9OK9Kg+WM6XIOD6xJqjYPPFfE5Hcv/Y0rwasvV/Eq
NCQE82Tj3F8QP0VnWJ1vMRY5wlV5MqGJANFLs4SmbVHD2UZ2wBeMJKyPENVOKh/Z
X3E2MBIU0qRPtHlLdwUK75c5z2NcInxvoe6j4XXHFoodc5Eg+m/p/jViR39Zb9ex
KGDpWg+UEYizUcXXJ3QbTVy6XmoEHZsstT/v0/Kn36Pn2kzq3VcAL7+VkVAI2W4A
uwuPqYn3ioYQN+WuGIpPwtENTTwRj/ExztbaPv7BNok5lpO/ofDDr0l2NZvURM3r
7H+D0xHCyLki9ARIC/Ut/qf9cBap7WkS9JRKmNZBKtRdo6joO/uwmgH3qI56U8JV
sB5uhof36fDkARV4BNfiTeNDCw4X1/ysa26Hi7hZ9YQjKTVatKmRpRRvIwrdr/IE
n4u51w/i4YmCATRxhxWteRl06mSc4ccihvWLQh+wlPIaKOHRD8BW0HbdBUwHw7Dj
4UtHgSCm077ta12ebzx0URgujIeFQs1Sf6tf/pJIk94PGtu31z1MQm2GvAiON5I3
x8I7y0tGwRs85/qgFnSFq+ehLi40WEp5Ld5q/vnPAM9HTAdqHhSvG9RCX4mYi9Bt
S69sNcWJSAqeOivHEnszMTncNZj/1yfT6orA7a7Da8DxG7QYwUDtYhR1Dokrb0g2
0b0FLaoYvYa6Mchn7iCEJwvEXQDjieuXl0XbfcxfqTbbesw0gtQ0xOpR/+gP79Gv
xRD00QoVkkLp5y+72DzofBKsCf9WRnLtUy/PIHrE8eF90kk1c7WazR3EXGSzXYTr
sK8QaQmB4MVzyCvWXH8Ea2tIUpMiYA7cS1ZboSP7M63DX7kbwuPZtJK9Tnkv8OTW
na+XRAXRttrhbyfJcRUzbe6YopMcSdL92idtuzbmIhqRas/Mdp7Et6h2GS67iJJE
TL72yV2ikuq/7PRaTDuyUlHjn46hq1Qv/D//6fqNUimxHWDw849BUfXZQfT+Mk43
RujaRsbQCSvFff/lY59NkKbeQ0QIKtdcI6D4enOIHLKDfMR8DeKcmRr9ZcCiwdE1
lG313gb+pB/3QUMlEnFhAvVwwTxDjGUXpgdj4KwWGzaRL9CgK+Bi9R8dtCLwYngW
/YMDHOzROegdcpzWDFK0SYTaaowgbi9FcOoa84dPJya100dAfk4wJp/uc0I2k7pm
IQHkd6vjfrCW56eSCQVsWUDpCa4sHlYQKQhMg+z2j4RmXHKlxhgx7cmyK1vQrO2t
mwu03rDVboPgG9Y8hSMx/GFtnjmIdyQx5wL+Ya9RDpt2RDLKK+9f7tWvLP3X0vxT
o7CxUCjURnM2rK5IXbfC1T1NJ5h84V5RjeiKKtGVGDlQGtOah1h0prACp5IedYgu
PAaj6YWtt4lCtBzNp549ww6TkpKoKcgmBGQV3YbinI08HCNKoisAmVaNVqylBFkC
x0KDYhySr9eJ1DpsAA1GpmA+OPlasSeQasM1JYG0IFg5FaZlafAcnt9xq6lEwNCs
Kr1qOoU6NsUOp+pU36dVqtDAxOXIWYcxECQQKGYTVNb3BEldAoJM7uJ7bbufeusx
/DGqk42Q8PuZPvTwftHkYfF9LFYIDad0QDYQ5BsMBHeMmEobCCo+Bpzn3z4OvpY8
0NV3KyASduIOpDeI4jmhkFx/i5woNhe45pQSBDcZOnabe1LliHRf6wiIDcb3Qdxm
32lie+kXMvmFTxHYsEA4qONtgK1Ovz8dLTlkcfo1Ev8/075wiTrIlyOAkQJCG1Gm
gKBAvVCH7IcrlMo/IuaNUSh4t4FfvsVW6VXNQGRyyJZpox729B6iG0tweNaWT97U
fPog/yR8F+R5QVLW+4rEKJ8W6fbvOToYm20GPmoXao/oMtam3lDNXOsiNtHPm0Vf
S3cCx3duo/ahKEXBiXohLLySDrL+m6iBE9mLhSPI1eeDxSX8ZOOXY1yc1jUmhK9o
dCOqWxP3j2Z0095auSEhgt18xywtJPbBzSQgKRijPNGRvwwGtelU2C1q2K7mDYhz
p1v649xFJg4NgLul5AevU5F+U1vy6KCnS/sZJMX4qDBFLD3ABj2gm6w7k0VRWQKE
ro6lHF+ztzAhzV4O4MzML57y/HMtOrT1hcKDKrzlnet67GLB1KhVfSIpfu15w0VJ
46crRxfaVwAsCno/xw65RSW2SpXcKAVgae9rTk4lkITAcpBaLpSpnTEu0JvsYCFV
bUHL/X98FOGEkLdAfrV3GKrrvzJGgnoj322fIxL/h/YNg1pisdjb74Spe3ZzGd0e
BH9S2sw7PJzJf/QptmWXkGh/mpBbxaTg53YD32oDU2IXv8HUkrQN9YIrb8CvcNWr
OvC8QnBYmgDxolF2+7rVtOXhFcWwUHubTnM3Ge9ZTB7EVw1sJXCKTKWpP5Cme4Vb
Iy2dp7i0y7YinYP34lg4lf503OrMiwNw39kcw1hqXbEKp5oqQzFMzroEZ7bUhtES
YINbV9II1ULVVtmbh80SgvycbFWkN25A+mB+76a0Luvxfv2KXhN1Tb30Is+hAAFI
DxYV48r2OLw3JhW4UiMfN+T5FzTk2YRvc7LHee/qS1HTE6l+Lv6rUtHEJ3VsS7sy
RdJpI5A01NNWN3m5VoMwueVJWcw9JLICBKKaDl+/kxq572tEnj9BQMoM9niTr3Xi
yPpMFfOgNejVMVLfaAJ5xds3/oYmv6RsSi001C1YlYD6WNCmfnNG5O3rcBVob0Z/
wHdCnANWucf/HUd74xVUw5IOH0FZOanueF/2U7fcLQMwMsIWJuCWOzYZLk4/Gayu
euBRQYphTX41Y5tpDnVlvO8K54qXc95a1gt5zN01RnJTPhsfO+bXvBwgiBbu7n8i
wcfe7xOGrzGOM34DGbKdiaMBSprgSz2nSWbwAV40vyOlqx9G+R5xnQBR+zjydBHp
NmyXuifZETRYAjcRUwCibM9lllQMAWCPaY7kWEuFs5XU29vl0ONkxd55ab9POhQC
xth4m646N1dkmOCRyoOEtVMtwlR16L5LgI1GkY+GFNSwqmqM3dGIYuDIzfv4UBWi
fgtj5uI3Qsd9NVoiGJ/dTaexjYNMMK3Pf3gVqYztdnHbf9QzzNInNf+sgpqjmxgd
OY4GdR54mYCWWPg4rlsbWZ8G8uauph9nj2peqoxqHTUWBWZ555Jd0dLsXfy8LikC
1FMtIod/XoI9eQ/kdkLNq7IDwbwnsS/THM72KYqPalvw1ANnewKva9HU8La3i5t6
tRRfbs/Eii2YV56e1uL+B1r6lgh+iLUjC5mfZVPp/KyoIgaMTm3NUkilWTG1tpQ6
UQ6110LZuGxzZ/fofkTIJ0ttZ3NfUoLVazzbbjOg2jj2rjZoaEzIXmSw95/WO9+v
bHmHFxhWXUwRjfwdDap8WzM/ybb/oc+CnbL2L/UXv5cOwO61lmkN7U3GWuE3smfn
7VIet87W5713EHyEsA2Har2zyq9IBKGQGovL/Z1LHpM6zZcnPtRlmybJ4iP2jDyV
dsHUsDa4P856jaGQp/LpNB2XMo92lH2gAsUrWnPjfDNeF4V2YD3eQFDX/ipNesS8
AQZwRmA9NYQXC3FqQqPv5yVCBJKEeUUQGHmpzR5Jo6F0LOSax9Ad2KQXKRRRTTKE
GANkTi/ZS0jMEPhqNBd/IT8P/WNa3oWV0Pc1qxrrCf77EFwvSy6a8FwpYugjzGkW
TwtpjmmOujShFXEIuEC19bC+qZadjs0ZB/E/Yv5vRmpOl+kAPqxJjaNR17S47kmj
4Wl7CVS6tec47sKTfm3BHp7H5U+SqapAfjscFdS2qXo+8Dt5Ozzmjmia8GpN+w/M
LYksoA/DwwWXBrQx0KxxaXOj4evZRzbEt3HeiaS/nUC+WGwtvq15qSL5I+0wbNGY
AYKf0NG/l0l6Us4D1AOXJBAWm91fu8Aw56X9HjlJ/f7BbJ5sLp37e3LRJ1LDGQSx
p16VcPezfTyJwEf4PPQ4ttZUoWC9f2gLMS1FGnpmJuhIT66Dt57VkMCUj8J0PNkr
0xzdUTfa3A+q9MvveqUQIPl/4mtJycayX8xiU+tPpVoAiS9rqigu8/wzO7IJqT1k
uERaJLg75VrQVdU5BC67Yx9FiheS7k0NJHivCI8HoYZlN4VJs3yHRKGVGsaMspu+
2TqpBzm7h+r+RAuxeQt4Y9UXUfCmLjD+AqHelaDDWk8AhDa/7X/QHloDc9bLScLf
a4FAncK3xKsjQd2hUaizNd8+562pp0TlxSguAIHTy1wKndVj56fuV66k6A1dGdTl
2w1WRdi5KE127v6waZ8rXERF1ANl9WCvVmOSfUCQeCVpO1wLDZoVHPVMKPenOnV3
Z56dxuaS7rks33732DHtvIdd7IYA1E0e9Kmfu53O11NdEGnnNwVBX9/NWk2Ocxl3
57NeHj6wnqwf8HYL8atORc++xDE5Mdk2y2ex+VDPiKT46nk1H8JVf/KpbgAwIWuN
zA0uXMHRz+9FqxdpjvDTO5EqulJQlZi3GU3+dNcLh2vJDy+sj9IWMRGodc/FebiG
+cNCrEKjzeXXYMHnc1PLVcJJRJzE8gHHkCGHyVglpXXnsXPUmUR4xW7jvt458P0T
nJKi9NlNbx+9xrivsNKVhQ9NaRxnf5KhdTmYgrgC27OiJpZAbpojL/mbN7BoNyLI
MRBxmB0g6osnetq5Cc5gOBvuA9LB2C+MrWe8AxKXgtOxrNQnEiyrrEIBDkBaq42z
PXcozbsR/Cq6u/XqKG3GKUdpoUawiPrmbU37WUO/w95wPKTQgFJjZYPgrf0LfseL
JlyaZX5WGjYlOebvWGsUJn2WJQ9NPGeS2AHEgF+wVIRL7py64k4Vd27gYdBbUyCj
hu7Vk3lN36aVm/cytjUOJO+WYQxcOor5K6uo2Dpqi1FruQCM8zQP/cQo3rADeuro
kpiO+g4yZ0kU79n5wfW7bgC7utiTiP555IZGTYhYI2cowJKrgktgV5NUp+9o0AWH
fPf3JhaefjA3IbFoefKdw6TRYxN16Nz2z9m2d9nQzHvIBls8WBB7OEsh0KIZJEtp
gV0kF/KMgLJsHvDAU1xkTvPLGIgedoI2iE0mVZJCEdA//zh73T3Yq7sxdkeW8yDm
KZ6d95qWiK/FuxN0IAFqaLxQ6vGH4Vd6g4NPF5gc9BkIzgcbx84osHR3d85zUISm
Yr+7apCbe5Z4D3h8ikoQ6KWPVbKYOrQ/aTBBQR6Fwztv5uAujH1kssSf9CROYF5a
9Zl8mQNNZ9mC6bz6dPxVy7v3Bg5SiHnEsEMxXoq5dgOIxDX3ZhtxE6tr5BRWCcxw
TIbsjg9ANWRBw4larKYoM3DVeWAyp9YG/nXtpopF9Q0KY8x2EFg/4aGD/uSVk0S+
7g/KfyhAtn3N0hywh8MHQrVxWM7WKY9xugW13MZZmS33KDGDIEkh4LRIQd/Ah4s6
E4SL2rCMRnGItJrzEtxuNWScXUqCIWC31H8UE0n/WHvRXQFV1YxARv5y08HUw/Rr
CbK4Fc4jlqFO2nmsZXwNLvBfrV102nQAuUWtpclmGIiQFe7v7JMiPMBU0y2swX2A
BUXlNoD9gLkFXjw+szGbdQovnGdtUrcW6PTrOq7n6gOzpA3jAHZCApzKQ28v99/d
y59dblyU8yTktJipr76bsfE1K7Otj4xbY+7pgGrkDZ+qT11TgVtPLNHjguhrzlUI
1VgJ2crnbQwYh4L3NBN5UFSgCEhdPbrCV2ko/D4ngntK8PTTaJ19bbuRNMdU0q+B
UT1aA1A7Z9g93FvttdhMJ0JJ+Ov9/UP4LWW01BWbv4JchhkvWgsAq0PwU6h6N6j1
NLS2f5nwMGDD/kSqBiMz40/G6jBgpqg0RvQUAdxpPi+44snkDzfgBDvOkjgOMMRG
1vfdhfGWMBkNEwg1zllLODjw5dwfSvf7h9RVt7canlx6QUyrkcFbO5UmJhnmknn/
YPQSEKWSRPSOxNZWDGQUU7QZLD11Dd+2uv7iSqCsIyMnE9GMu4ecE8dgWfrVZH6h
ZF3AgnkfbG/a5rhmWb70n2cA1sVgc1+yZ8UcxlnTzwiGoOb1bKX6+xSJiCKZUg6B
zourU4TdHpPGJhyr4rKTpC2MneZ+wLiaSJTO0DAtpGuTycR0g9TewFPYd/HHbUgD
Z+HhRQWlhPjcfNgv2gZNKdtEIKC4D7W1rZGB2r7GJLGupct3qcTH4RNzZyskCQds
nvcSxKF3pB+CIvyMB3uilTUS8oI25Wece1PemwYwE0O1xiAf0MKpCub4/5q+YdIr
CmAWUViT9BxK/qqH9UKx7J6KXylCnzEO+dQSzmSNLY926bZlEV6d1z3kjLfxV5fm
PEr/MjXe/qQk5ZcwuqZq9Npp3XjluWRdZXZUXULHFSbyh/PMrCXylZhO7p4BwhV7
oYYCZhiyPmD9I+YBq+bZCoJMUzquPdZHnYa409jwCqPAvRvuNBCE0NM7J/XUbkMS
uZ8qBNsR8p673pmP3LdcF7ypd9EXDQO/D7oA9AgAFOAdhRHUjzxNupbNPoYm4Ibm
M/Zns3br0920TSgHah5uoY6agHeNNvkOxqGQJKdnbDxksuECaCjVKjh3A0ntvMNx
QLp6eoKoy356ZgbDBG4Fn6iXVPIGv8dp/52LsBXwYtCwtieRzzHi9sCqxVSzJvnI
baKhJqXA4BYO+fN4t/S3LRaTQIp4ihvLjfd4FYRndSaJzIKi8v7kA7xd3IBGuFZr
qn2QbHYUuyaiM334xhgHyuEytb15qyKOkVawNPC9wYouGH2FJt/r6o9ndjn90zxU
HnQJaeDwSKRHAJq5Z4r66SZW3G8cMK84Iu1d2kkIAZRHmaZRjMRD+rLRdFuGJjdb
puiUmjfqUw8U27+RoxsKP8SYtC1u/wN7hDKo1d0R1dmOUdS/Ul9/eMMlj9z0KFA0
WdQ9RDyiJaXHo80koyGYCOOi2OK5zv6J3SdWznM9i0IOt/vIoRziqDvVzB6Tasg4
Mvdijd4NArWuPSgkWgnKqEzpjMIzEPT31SwPOrR3ab9bkZAX0V22trtkLQv3gSfY
ogTRm/KWQu/3jQnCTNlaNouJ8r6jBQmLTHicFUSzCTITPuuk71Eqp22kgIVZC6x+
vcsjBt3Mj9Ao0fGm8cPxwjxc9GkYRoRz5tjwAdu6FCwpMXybxktWu1GPwzQCIwa0
KakX5VokyRimYOOfitGHBal5MhaxRjIqYMUxnmjshGWMhCUEJWC0+0FuYCUb83Br
VoVS/g7ke1/iGNL7+szYy2fcIpYf1xmImxNnia/MosCu8vgLklpH30z3rJSHapc4
sTbE0A9scmGjjs0E5/NGvuarc2mIzvp0m53Py1BkQE3uxtOkSdHvndCp+Byx6S16
eiZgCXgogPfi3rUP7MngRR++6FWKki84pr7CmG/3KEw1Mh4KCTYfLfJq9TlTm3WH
Ht1OxvfJFyPTvyBWBPlTNV9s669gHB+M4BCV4YA51IofIGok5gDi1mEeZcyqeqTq
BhjPogb5qfFYJbxSckeFF3GW0rIP5NeyCiDyskbOJRuRvQ4Q+t3C1E0MPY3pRmfe
tLApPWMCBdPKnxou99gjNsj8Ggj2MBEpm1gQgbTemBSail8y84sF6p6dMj/PkXRr
Cl4Yk6NulPtyrvnkPsjPvz9nUR3wmO81n69mDDtwAHDF7bb27Gz3Cyj7RuseYSj7
YdukN5dcpjtA4u0XYWXryM+kGXBX5GaqGc4yShyzCPvcvMMJwLl+XLr8tQrG3q5/
uN+1DNMa0Iu1d9ZBx+HdfoZFnFMrlSg+n3PLDu3sg5vUxH9puTPgwdc++9UljFYN
/ER0HQj2SX5/kua2cln5/bJWGKklbV5Wc3KXgTIdLiefRBvlLQqUJOBd54lfyQhR
nnOsUUEJYx8H3oVOusQ9g7aY/OLcBsqgHVYvPyhnAnlRZTES37wms0V7nDuk219o
2EoEYXIV8rGeKr2li07lCN9CC6gV8iKdmph9z+GSIS6RlIpxIxVIx9nTyVePMeRs
7tO6hL+fOajTio7IGbSM18v+J0s44/7tUTdq3S/8z+1ijE/KhAGpmOoXdw816cMj
v1Oi/r/tT5NFACFpKZiLqiuejh9y097yR4KsB0TspBvQW3qLXCmxjDHiFxnKLtxE
Pk/SHM4jYD4Fu7oMnZqROGrlUavxj1g6RAX+XYHpI/N6j4TlGd82NjIXqTdY6hbz
LTYlrzjoL11Jy1iRzDfGbmS6nw1eF2OHX7fFt1+4NiugiFKiqN75FIDaZIuhbHWY
Mrvj5+A69fUp/gV+wkRCYR8ypYnS30tWNxyYxKw7hrQvtrDIX+lX4hMvHtsSYl2d
MLuHmSrw6jgp3phjKZ9CW5tGNp2oGPw7yKoZFq/ozMoe4vvSCafX5aTBdQTcDYR7
GsLECqGO1GVj7rBxuczU7ZFxw3wvcPPbbQn0xFJKIN/CggK+fNY//ZLISJKiV7oQ
52fqlrIRxTev9ihDBlEq6RpISJ5pGlm41WNjwayrN76PK30qrNA8ANSAR7xbxfDM
ZZjSs20H0VaSA34IIsCIhQ+hYKndPboLm5cTxod6q7OHf9WzCJTFzFoAdw+hCZCE
mVbAsnJGoq1wLtgUdtID8Z5HKrsYLexlITylZYAa9CkcdpvMpJA66dz2MRbfC06F
kmjwhyssjqcpbWNaVruLtyzxHCpeSONLZrm8q+Uj32vfL5ZHXKENYV0Cdk239LBC
PjXuTEAcxbBExMKcvcUfSoQNA2UUnID/5p+/0KpDvLyut4JwvBIpfKAZjbvBjZVL
V7vbFrxoA2T7Di/ik+IdD1Td1Uag6Y32ljWqL9GZxESU7cnt0C92WIiqKjlbG+30
zsv3i+n4UdVeu4F4LpkY3L6BZCTcsRCQ9msTmkV2uz4ZY6fUKJg29Ck6c2tpF2eg
wu086e2+jbZh2K1IK+VFWwnPJqD47Pgwenlix8nA+HDLx7bz9C5dXIQugq3e2/o2
Us3nqAPrIkhpLUUApV2lVZVMNj7MO6dLayQN3K6C0OnK7xRA22WW/M5P0AUa/FV/
jcwbLSqKiuC2V/iFDubNLNiLkDpjhM6w14uYFpZC60fDyc+29D21JLMc1ZSv6rdW
wszNTdxhNCsyEjMcJaNjjPCF4RFm6+FU+WwLnHpDPwNYX/ryTKQds2Bfr0MJlPbE
BF61dbuojPZ5zZyy/xvVuZ7n1jtPOyGN+oZF+IR9zBz9csPghvwUkfGk7F8kIYFd
1gK5PqdHaOUjF1m3EfIs5Q+3dk6fDpHYtZH8uE8l7uyq/cGIxhsRiKNdC+4gzhGH
Yk1Vbda587RTKsKMmHBzCwoS8jpMgM30pE+9GS0AmKlQ5IqmJwn9FIyyOCyNm7bB
Ag65/aQgIDYgvqpkMJNrkzbVckVgTYoFFY7oaW6BSLlgxXGvEb7h9DKeV0Sqhph/
z8GxSdmBw/ZK5uWIaI/wMA4WfkNvoeUTmn8jXMgE2pMdvgkG3stfDPwO6/z/YUqs
cSsRmQa22QUSu/ZuVcSmj9KshcGaJOlYck9HHmnItCShatyHXmJm1p0Uj7+Sc5wk
McOAcnptA+/BoKceXOyQHThqN3sxIeypWiC1vvAxC3wXMjDZJM3ASsN7WaS/bXwH
QTDS/HKQq1TRU1oGYthJ6xm4Q4sgTcI1WnhLIGRIgoTJBTjRMcTbzrLrtGARBHI/
MUN9cRBVnm1sOiNn+3+R4y2UXzL/xzee5tJ2m6qmitPFJqW/Sz9W+h0ddUwPrveg
md6nKU6ClL6mOGqeWfUQa8g7OqALDC0UVplnIAZSkED6ruVbsIsVkJBKu9NrbyEA
NfPcGbx2akkASxB78SuAFHhSTCe/e76/tPEaWFue88gvBlpDaUsQi834ST1DewmT
ptWMluWT1+xyg6I32WJcwqNVeOrjfgsYeAmDCsdmqY5bgz9EXtUl353PZmYb1W18
eWPYcO5xNp2DQ8YQ3qRDpbMu/K6jzW1Ot9a6xw3W6a579VNUbZuC49whbzQbZzzC
vK5LrcGwcpXVnc/UvEm4G3mSwA+oFsjF2YUJVgiGF5ffSXkN801kmp2ssyPYwDXv
zyOguuz/sltx1fgnIeXHyhnwOLXEX7l1ZH6vJHQCFmz75k9LONuTETkSXO6PK2DI
i9tA5TASekWcqD8wDsxZS50YRvxK4hLkMlwBA+GgfmDPObXX2rbZHtNfhJECbQ5T
MR51TuC1Y/AAKA5TBEznoasRfbcJmScjKH/Kd9AoaZMPsOqq/CCo8Fe/SazNDTHi
5kqiwaH9yhywrAA/cEWxrnayzLZOIBiWIIU4NAV2p3PP0Cd6PZye8b8zwKRlHL4m
5bknUNyw8js7mcsgEqJk1+nFbtIg184th2qen1gwW2JmwIfVarrImKKNTbvra6i4
InqIBy+y68klGB6qe3h2RuDRjIku0/vAE1J3YVbzsI+/yH/WUw33BlFPZkoG0yjp
1ET8ouUPPZ2GpijbfpGezQiRxMUX3VXcoT9sU4XRAmU/QwhBvWFWBjziAOYIJMTA
yc65Xb+P8TBKNN/LrXzerjKvVBRgnvOVqNfOZE9opInqCL1PNcWUvHtoehMkjB4m
auygrau3ytoZccX/TVJaisVBEC6OfeX55BZ2QQ7aWJ3AriHbya/Uaf7MD0KmrZdh
GkpMOvRNOBXPFZYwMtbfOciuX/Bl6y1Bn4hHfMAC2C2/HuYE2S9THcL3K36zveMs
8O/6Ts8eMkCc0E8q4BQ9suvZdrfaPMpk1jxxa9XelMYTbLabIlfLvPdQGV/z3DS9
XAsIWAF5eDtOme8EM9fN4G3QB8pWmOBpbtVVE8tAmXAPrHREv5H85mSvfKG+GeCL
dq7o3vx9TDl6LQJ1VmaGe80+742EcHDQ86VDeKwrZYhVwM7lKvIe1FjgVlooyNtv
2EKbJ4wEuhVZ8F11zbevKuOBMgIJ0765U8WKPQgDTSAVUhVvIkUGDiSQc9u7DPnS
BQ9+EtFy7z96yblE7Miu0fqT3jssuPVrtfOfMMd5P1WfY60xsrP9ElLg+xXxS7LT
gx4SvbDelugCSe0ppG0aZyQHp5FtpH5WDtoIOGap9NQWYWnhoSqz5VLJBvLBuvDF
NILobArf9d0dM8bhhTKQi9M/N5ecvfaJKnnb62zbJzOOJ6bLY7v3ieCs2M+slMAD
jMlc3xknXsYBAu3tfhsJpPQVAyrf3PXDk5k2ijg9xH5oednIx0FLRsvTTVuzsQll
BBESurjrBag9878hfIqbrD2CYU70Ckbo8PGhcv5WCSW+TdZ1x58tz7LniPHacsmv
GmmgqukBqga0QqQ2bY94JnyBMmiT1SlZnFuAVLRy2AVnjPG2yGAib+EzIeEg2sPR
46jlMXrROw8hSNXsztKd/bydGQGnT8SDWd63zXIMkNo0ihZp9asCK5NxPWYlrOzo
yeJ8slrHdzkhsA6zhTt2AKhbj8KC8tOof3gmxTHlW0NEknSmLoNfzZ/u1cU+eRpe
GWIXINhkHDMfdO1HWKYDmChJfCMs1mh0t5EjUBhPUEih8wMbVsQuuMqkZsUqCM04
embRyxWQ7h5OIblTXUYQkxaspSeCng7TasRaIE8/KqjyPozdAsMt1MW+k9mFhTHN
tRF8FtlW/zWWKG8acDVb0X/qTKb9IaqvvznkLaJBOH1yp9n0c5GeFKiLBEWQQKnw
Gjmr5bwacvxOWrjcewqf+rRWN/UthyDTHCjs2Bg6TCop/Z2GRcgJrI/0F0Kf1sMg
XDzWmLZJvxjlHJc2rosiHytunABv4bb60FmOt0DJZ1TlezcrfXNQn8Px09W73q54
l5JO7e/LE9KVmzoLViy2YmrCkA1UM0w+ZVWfl0oNkrJAZPpfIPL/88WQ8AUpSyLp
rtJvUIiYg9n5738IB5TdY3md3kwnAl65APrb6atsvgFLWtKD9sGFbnBY13v1nWiZ
CFA48XQ8rVZIznxJb1PTx+/1/owQ36Ao5vrwm2hMvCnpgoBfhm3KEY2+JKil9u9f
oRWpMyl+TSHYd+dDclm1qbFab/t0VIWfXAz9sdYFu8oeaAYovkIbkN1luhG3KLsY
6qHvMjQ8n7a/CasNQ5xFiD6snMFcv2rEIEc8yZ7Mnt0DFMaWdNj4W1JcDLpNRQY+
Mdt5JE/hnDjiLTrD9Wq4M3Z6Fw1TvXh8l+sEkT4zHGp0r0lQmbU/gSetiFSyIeQe
Fgx+c4J5Or9m2odapt1le1N3xKsipRNNZzfr7QZLoXqaOWn1xPSMO74NjAlUuB7c
Al7C5JW5vd1l0HiVM+HOcCFrtX/eHfRq4P0Qk6BZWK5MeDlQx4e/rxphEysCMuBt
A5S+O87TZcYTXs6dotfep0TeqSJ4kP9sm8eeuCt8WyajtoeanD/xuA6fv10SptaE
jqPLOgZxGXW9VQDWsuQxJFPPSgAS8o16JZbaI9t8ROEVc9fkBaXW7iqC61ZcUTz/
QxKwHcmMg87AkGqbF/f4SE1vUMWoWPe/qV/m5aLKbdqTWMl83I45dg7BYcriMq7y
eEoWSBDDUXfQTLHGlNJ9ldAcqLqXGDMeUzeIv2aC1MZUVz9lT0vLaoJSD27lFv9/
3aqQ4ZhrjlO68eJpdZEja+w4LNqfT+RwE7xWSP596YLqA0l1sW9ETP2rGM/FwdvP
ih6I6fbZVAMv1lF+YbS5nVVB350GeJuR+dj73nrSPBXRno0NTas1bcr88H0HbSBl
ZqdmSWyq8DHohealmJ6m4R7bREGZ35f0Fy+X+HBx9BaeLAiCN+B/QuOtJcavg7ca
mQHVpBDUEifpEF9tHFv7DT+4nHR5O6wNU87y+6EIkqQUjnP/UHrVZRsb9dsvgwrb
Uw4R/cILRuE5ia/enodhwt4HSs8wcj5bMsVBwzraHBIqnXlRaAeyCH3gGdLcjp5w
Op6FO1NYG9w0Zd7sjXQOVclMPsHA9U+6ukMfhnTMQX01LruZcvy27/8QdMCPD2Xv
3od4GO4QGgYXZRYf+xaH+wD+m6L0Car3rHuBGC1VnkB24eUrZ728PvT66MYBfoJp
jCIUqfX2W36IO/XPjDdONJKYadnNtmbxBr9cMgwGQxnVycpWdILEX8R4Mnejj4ix
Oj1cH1CTjRHrv2JVRrqRLELp+5NrXKb2pLODtlYk81uTK8yAuHmx/SWREIHDT9E8
ZeX7LDW5lzrosV3vPMCwcloBLQYA88JqxseHt3J0PPzW/OfXS1zru0yK99tEcffG
zLLu/nsBXh1ucKIK2MHZ9nhkXivjrR3g6yXrCcJ2Tr7gXGb5iK4ISufdpe+TyLUM
BZ9jy1C6u4+rYQgx4FGqDU4HTRewjQCkE7MVtBu82/6ZH8DQfZMrLQF98pbdRg3F
v8Zn1Pe723sGQvbx0mHbj0HO8kci9khun+R3n8y2zmEyTw7AXa6Lq1q3GOnCNYSW
X6fQQJWbLfLoP1iLI0aNrvBPIP/G/Aj83p5LACNA0JhwZQjdSBmISkNvUXrY8Ugy
I2bwSUli10pZg//H+Nw1VG6gLMyEB6/5yeltduelM16h5DJ8L3SmUgKgwmvBTaXz
DzaiUB6cFv28c9MryA690sYWvvKhHvUMcYr7iiRgtlsB1mpPvTj5FdDjI5QXm+nR
EPiUG7C8smkmSgp51+KeYY5lrWTuO2KDCkexwq17ObsHwM7Ps003X2B971+8TX08
rOQSsMn1V7HZLqaStYRyygA/ftVdmOzOXSvWfMkuJe5X307xBbWTX6gkvE++6Cxs
WzKy5xy23jaCDdhhWrm0JLqLLF+Ezx8MeqRRXSwLNSqmeUazmFD9mFugYqRk2/4z
Ta87PJJVd/z6zdaknDh1gMOtdSqEUOavS3kpsC50Q8VEm8ekuyhupj1aC5t5gIgi
AM0/85+Xd2Gg+CWqMPba/t/G4uqBFWVkx8fys5D+t5d6h2b6cOZsXql9JDINgZnc
7upgQLC7ej79GXie8Lz9YEbF12BPFnvgqxeCbw47vrUbgdGjGCmvxnGKL5YuPyGg
rRwlEOaj6JaL4CHvbz6UY7qnUFZk44VLma8rwor9G8bIajpZTSCRgtH3j1CzRPaj
/5FkFsd0BVOCXc5z34MJlof6NSYnh/CqA6RArJQKX+SKOnujqUd3ps/bJO6wJI7X
YRtupsvJghfh+QtX6mseHunvvYESGgZP1GwJWmJZpQbSTpg7xp1iJeDelml/tQ81
SK783fhQaPVYAdD7/1kxztOzqwFDiA6yTBTwGzpghcpgrhFFLbd5vbJeeHDbjrCg
YdIDBJdyv/BZ2BSJJkSMCvOTXDE8X/NsjypS63PKCAxM5qFCcj6o1EEy5K5aXnz+
0Dpn5BXHPzfzlN61g4aFg2NBVfT11+nqG/fJdyQq9rlBPP3KCd2xnpO3fU9/Jw/f
J+7S/JEIT+XRpG3hX0kOu9zMO9MwtlczFuKfMw2N0jnhxonJxFqt9dH9l4xUBkDl
a9dyTDD6TXCmzVWlPvfkCNIS9O0XdyzIbWTUsb2QFCPT2tcxTDZZvkZ/Bm1zqQEg
0U1cpjxWslaFcbG/AZ+EjBH1L3wCFMb8B7PDPi48wAZsBhLl/bLR5faz2febFpug
kE3x0YP+TNyQ+W/cfxL5JpNYpcBggz0pq68WZLtZAP4KLTVK6CUrf1Q9uiL8ISvu
9VVRsPbtVzYg768g5Cx954LY90LOK7UgsFmpIs9cJuvS4oiYI/nEF5jvAKCAUDPF
WMbI3wp7UiZkvFSms/fobWSMCkufB6zmS3pylm451URZHebeFtKRC82VIEUQYTgF
0yaqq3dOtjoVQLuM15JdbJkTkx1YRAlrOifDjFMm/b5qY1LeHtoZtYsou8/egdfz
spaVMgMn07s2/p+VYHtHUXXf6FYBlQYKM+8iZa6nYboy4mGta+iqKc+55kSflIOw
iUG2KPqxXKFAH1VMsYI8mTU9Enr0M58bjn22L3T/aDizNTIM6l9gTdcuPpCp4jLK
FwbObKVrOh4Q5Rgbef5EDDN27b5cL0zRsXBlgbLX5bDY6I606R5MON6zOD3eqHqE
KQOE929P9cCOgX/2c2QX72pYFO0uz9TbWJnRHwVrK1RYFx7/6LFTBBNNujsXsxIo
I8hN19jxmu7ta2LbDJBRz0xiO/+uLb0Fmwli2vmDm3siq0s5URTuReaNOSA7jNBc
KHsL9Mjp4dzooHO4PxC413jnS0a99qG/CJSIRzM8NoR4Jt7dK7lLHVsWOXK7qtCp
yTWM1z6y0m38zUbyk1vuF9lLejONbWKSvhBAPussKGbU68HvwymLH4/GxI8ZeOAy
3ihjFfeervLGs//02p2yoEnJ2vWtcZZne08kWkUQjIxjsmmg5+dny2FzirOQ0I7R
/aXMHOual3aTyqGg7sKV/loAH7DiEiMLjIhNwuhkGpGPIPxpHfhpA68+Ao5h3CQy
wOkr89Wpbx6sptInuq4g7sJKcQzzxj9680Ne+kdUy0wVPGD7r9Udn/vrA+X8iGE6
cLhBqKqT8d4kXVIcKRkZb8UzDAHf2yzRW81fBeBdwekGhNev0WQ9WT3iHWzLjodB
SdZ/Yr+NbU5iuNmRsSgjh1qREMNbBmQlwSGakepBLujZjzIY9tWfEMiqX5SzImzZ
nby3Hc83cJXDeWUyk+DPWMokVm4dCm2NfHsEPXlL69hptEvY+KBKT2isHj9Afzge
7zTH0VvSRBRuVDrvBrtAEX/mdL1Ql9QG8bw3irfwwwxmsuZHjVTo29Azk9Ri51Kd
VZkrFoVXpEBXgmPaRJZWcPA1pzQo/8U25s2Lnv22qgPB0SbOCUCbLVjpE3vJuvEn
Qg0hKUR/Bhf5GisfKN3jafRpBqTFXFm2l+fjqSaZyWONjI/9M1mfuSlI1z7T96sT
cgDdLgv0QLYTSECYBRcGBiTrsMKGyU+PgBFEE40GKWjCls0VsK36OZQWgVh4huxT
o3UrJqtnyZCNHeockoe6PNtLeH8XdtIcT2LsXJ+iRUk7KDoUgSnJrJJffI8sg7u6
JU3uc/UkOuVWEFMFvccA3SGxaxzxhnnzvPrIt4cbXntBiO68gwlRICwsKSMqkDbI
pD71FetTc5ImkRkv9eH7xOpr6OovtT3V5NXs0MMAui/XZengytkSfQUXXXGI6J7A
cUyR4kQBuUgo6kBzZk/QDlmXZsxhtOTBLZTjhyh5PUFcBuIBKJB6o3libF3Va0dj
AkXAyMu4B17hGxemcy13AQOvNIm8Hh1taFrkwPR/hO7flD1mrKQBWqpxivgOFBN+
VlIimCPuJseo7NFQwhxwAXYpPClUlExis0GWhjGrBRfvmSTLIpGHQhhSZ8XEgsqJ
n5TifvGT8orytzGRXh7H5OdeHTXa9naio3XIrC+6NgshXh9N47s5MEjqHFGn/Qbd
TY8GHa8yDZeayyd4jEiHYguSGnSTFg0LVR6oBEJhmvTetnhF50dpaTenQ64N0Qct
E3Mev+bBA9/IbVPrwb89WX0+Rr5vpZYylFPoBxQKmbRlxdqxFTZpUBWuywfClYgB
O4w57dqJuqqajkdgK6yC+e5xM/uCcHoEyDP5CbcLL+wy0gGnQdPkAkTVNpRbLRRq
nyQBZzKS5EpT5/vGsPGmwo5oxFngQ20okS8FuHP6WwAIcOgVmU3y7lpqr5ZkZQ/F
z4zHWSkZyi1Kpr8XmjeQrVS2NTwnZYG8NP9DFfGs2EGmjeWW2RWjVht7NsIo2zxk
0xKbY5VzjEUr9aCWF2teTMusAUHHESERQQDL7X2UraIF7eLPDRvxRaZVIVvxP1Oj
276LEoeDrJWf8ACypmstpn41ECHF3ygonX36Sjq401nJ1agdeAvSU02ybSofa78F
SBf6fkMfnBtXBRpCgqozjswsGdxUCfcsO2bzMu1oqxJnls9weDA7/T2ppOGJ+jVV
pTS8rKYV5a/roRo7RToH2sYj+FLj44EPrfv6tHJUcbyXqT325FigMfQAwFRcgBkg
bRXLL3QnwWvU9XjcfdbfBmsJ/CLGEExdm2PMYhCXenQeIXHlrmvpNcvcn/8SKFYR
78gJpDXlQRuxscaBFb7odEreLDw+px5zQaVPu/Gi9kIhlgMnAQCifuckh2Ey8coE
lGJabpm6oViLeeukFFzaMtBJFnOWSOyh3J2yz1ykPr1HodoMojds3uUZZ+/zY8YU
WAYGxFyh/3yVofLXryfmGDsGy5SAMYeHBarhs0lT9YrDCLVt9HR5ShXtQaRhNpdb
XIV6qnHvycFWuICn7MCgDZzncwqbBp9zycckpe+PCFKlEZD8gaTzIe8SUJOGtYKw
NsdbSV/Odkhqhum/VcNfG58xnpwLSGwZvmPVWElRXIqFoCuK9DNZy6Em9GY3YHio
cm1rrZi4RDnB1lvKBo2nmbNqVyTi6yRIG/Oe481P4mu73BNWiBU3aln2/0K7XTPI
rGqE/hiYRn/SXNZ5hZse34cqLWV1tDExeOLXFWevjh8u55a2tTeBrpslzFXkAFAT
N8CRjShK6sXd9Oh0cEfHDVoBdmEu66SMIk6RYN+GbXRtKvwYq8eFw+t7hxbhJAoH
fEeahBBYEIzQtGN5s7k/P3NGPxcel40huMu12ac9GB9W4KRIba3s8LK8bBKkRk/Q
CCxcxifHrBAJiE5IUVEPWrS3NRwqpk7/xVx+HmFAK82j90c99oV6/PXADBe9yT6B
TnBATms0SP7fvP0mOW6mNrASu+jLknpletJERvVH5cqnYXOoroRG4EqiVsPTWgl0
j1ExKnVH8jnBksPfbLAWq/Y5XNtMvtpU92jgUNdHb84t1COkphG3qbbBnArhaW19
7Y/tF4WyFuCPHHBXqg3Q36PKcs65FZSJxS8d6RdWo7Yee9TQ9zwuuztW5Yf1XoAG
PcCgVW2dz1o+Hxs6hha2XnbctMFkg9oFa6Q6zQjo/hwjnR3b8zvJ97LB0t2RZfJY
b0aVqDcFC3dxe89w3g6/jXqZWfE2C3xMhWjHXkH2/snpF752t/XgWBhU89hTJzO4
VTWYwNuBnIkBjDZiPQjeFpMXCbUDvxnCVyJ4uUeTO7c090emnl1KKQZJF0G0sI2B
0NuvrxNVMM+S9vDgjLCBddOVyr/8dpm2xtEZzS6DpQ5B5ptmCR6oke4BpAkgBrZQ
1eeEmbP/QcKlAtPmUH+DrI9zXrZetZUs1NWjJxT2/38Y5IZPMJc+rwcry3u2oqkm
oaJrKpkqufZmoXeE3uLhIF3JUVRuoRDUSR/HbEt3NMFizaDE67kZxbKF/t17Qa5i
0xE/dXisKJRBFPeujDcShACFtzvLJa64fzRv7JX3fyOYBld3SzmTL0N+YeuBEqbX
glAQTi8bDkruBpq/dunoLl82rXaTaSjgrGNx8HBqAEjjxyslxweHtd7wRYfRCUC8
puu9ZlSZtfnHtpyCtudv0Tj1sMQuaRJGGmobuiZtU4lbC6o9BCE3xA7Cdi0ZWpeD
39g/3jcoRU41oyid2CXWFR0hz5qHvgHn/cJXSXsIqm0QxNaGLW4irlueyXwQbv4Y
b/9MqUpXqq9+wv7VJtLs/+iS92QRf3rtSjqWrfZixknn2KfS/JZX7Y2XzKKbKBKJ
2p8hVULcaBAYg8z5cHRc2IX7xIrT+HKiSj2fdopC+aCAfgJ3uSmlo3QZ+iUQai5U
IX8w4/Ebw5ZIB139TZ1f3LiaCqIisxa5DTdkR0fckYEVqGF+IfIrbh9qlmTweFDT
Olf2vHqi3YmP8vNXUZWE7V6UiZyRGaJOAuAcrIpbodwIFXRmauCOKaYY8faIoGVM
ALnWYaF4FwHiCWhyawt1/UYUKsWy6Hr2SnqyXvIICaexM1PLS3eHddI7pqU+3gkp
0Tny6abwDhDg42fZiMK+a82xuBLSpKyV8k4nobhCLGEAPZxCVRLKkhEQeL4Qjf9z
3EJNH4rYb9dwpuQQocBHjqCKxOG9c142TJC36lQUI+Cb9yRF6coOWTOcNpCZlgkq
WrpwDaMXg1fJaxs5NcE5H5RTQZgmVayS61Aa00gHfza1gZm67VEbh/GjWyGRTHg+
Fma4XnoETc9aQQe/qF36dZj/cf+LQfER3M2d3ceDTyraWUUol6tgxjX6zExaTJmC
6Eu+VoISdkro1WFuFKuJQuiLCXe2lz7p8wH5HxGK9+DFID2W/N8VgE9eq1DFX1kS
3Jr0Hca9AzLBNMQD1NjmbTuLLqhwSFiOp+KOnNcs/Z6atjzv+Ynw89O/PZIsZnxb
SRvXfINXWlRr+/GDWis5oMWL8IzytKnue9/24Zw8HcrLC1EhHzHzlTfbXPgWQegG
CuSY414Kz54FkMar2H2sqdExFMY5ZuTnXPXPBpPpCie7zvPz4RbCD8Ws2HqyBR5Q
Ohq/1SSZ0+lmuHgaFiYlWOg3J70YaVI57+Uc5TahpR+/PbHvv9LRhP3HE6YJ02oy
ikO9TDA6vlZ2vkZtWbUdB8nwX4msig3dtA8z+/+YDcaZ9LsamAkdZeFinatjPvg/
CThS2+RKkIExLiK3uwnTcOx+NdZo+ADnCLWogLxFkFV4nBnYm3KtAzqbt263ZVDG
0XSSPdSNj3iLIeaWCTQfxs0S9f3hjYYVDymJt6BohpeD8BNNU4NvSVtySlbtw3rc
6O3loa39kiJTQh7TfQlPWDMznh2mILOfnHSiR5Hmy9pbOHHVf02y95vowreNpNrD
bDurD0d3CC7fynwdT8JYHfKMs0mQEFZmEj8kUVzjdmMtrV2z/iY2nZTAowlxKRpn
Wb+Q4pWlnl1Tb7Xd64h3X6scmWoUp5Qo0GnAI6PlrxBxNmo1nvouHFIbvbYRttWN
esHcP7OthPFLe2Q1ESLFFjYXpgKLrePIjyJNsGtxtBdAz/wxtosCJKlh0xWSqFPa
9sgxoEwuq+tWBaSpwCwK0JqU3g7z9HIPOnGUqzHoFKvg/UGzpGluTaoKLOLQm8dv
XLNUUh6a+ZD670bSi/dbVLY5Vu2/uhV6E3fbrMF6yIIOn+wRWBwBEkpUUD0J8+Mg
qI+23COf2yIMU+/k8wm9JfV9Kvb/B0PjNVNxxWp9zYqUF8+GEcXqAEevfXBwfMQ5
B30eo8cyz7hWQQLmx7XWTwttCNA+z3gVMah6miBTP9ugp6g0MvvB0wIZgPhY20Ek
8lypZNaWjvxaTfmWTOcVFGRfAc+kcTtbBRDmN5Ks1fB4nqvgspnTHdWe9aX0oG74
Va4cFIlwdX8YTRAonDr8hyzXH1GjGWUldjbJZRb27/ciZsK9hCTRRxquEBZCaJYD
zcqPa0Wcc7mSvPXbQI9iUOLz9FglbsYIBKLtmUoMogVpBNL+8bLTh7IN9UDalyS1
dAkDUbGy92H8zfSqtGUbHQOxqw3gkWhgP8+UXY3qLOrBuPQ1zejkxNKjt8ib783/
FOBpLSeK/9rphZbIAPBf2d/NY8VXJgdHgIJ9mIv7g1PlUhk8lY227t5SyrpG2368
CdZ4iIcqMNZJ7rEaTyk/DhghrP0r3htylBPdx5grscIkMhJHaGsx9UMb9Du/t1tV
T5aqXNZ7OaWQCGg7l3FEus/AT9hOggUHxS/O/TpQIzOuP04ftybFOA116fX3+x+6
JtcvoGzGXnQZ5tsU7feUH0r/2a+1wmV1UbZJp0H0ol0/0ogM4ElKeRx2y6ILJrxl
4VMHtRxp6wVnF1LHYnCwNQqbgNzkgtI1e47QgagKARTF1wXQSJ9zqyenQHLK/TMS
P+02OT+cNm9mMfhh7SuZgklsDYMkti8RPkU1X9YlwkcJvIUigq5sTeLWYkajoMM8
+3EVdZQkp4/9cFS3warstqPV+S2CWrfHyJIy1yzU5YRWy2PlA3wYarnCQS4CuqEe
FOrtP/IjIoS17jBkkjH0llnRYzy98ZGbH2daLc0i/eHqKUclKkFvXASluj2Swr8C
Af1MvCpzAhFAZmIISw6OM1cGsfRb1/zTwbd9ggAazfxHMrIroUA8EkwEVGJaak3+
MQgju9CFxvMmU99S5mG//huCg989s3SJsPGDnXK5ZzaVs0gMlBGEZexCuLC9fy8Z
d7ffAknAAYPeXPnU8H6d0MInBibuE7hbA6R9onkgQXn6X0qorwHOFDdBlEcfvwFr
j7zUD1t7TJm3Ag7keS6t/6cs2tWyXupKikj5xrc4LYh8Bo2j2KfLRYsAgM++Ogt4
srvileFTk+aWUEBApPVSLjh/PYsPBiS02pix6SLuGOG0gIMuvSgwTN5Az/RhNwt+
6TzMqJKSMi9Thy7lR+vrP5foVsVasbbpJHjFllWXLlmWb2pGfpjcduL3pYGbwBDd
uDOMGo7pkwQ7QyS9ZzYeDvP+NtR3xu8G5uQtX1ra+y7sdModEYB/yhyNV9GsX326
opC3pUpS653mmlrZKRNKNhEyIXiRhzuWEQu6H3d0+WEu7evIlBg/GG0vGq7ZoMSQ
Ab8F7XaaF+cDhrpcQxJ14S43UzOqnfVv89rsS5FV9XyNKy255ZvIvoA9MY5O+/M0
NsW5xEvigp2pfGZrMpfqqaZdz/3+Mga6vPjfE33wuN3gSSdqBigY1PwRa/Lfsh7f
Xs0nMJs7TPKYb9peJeVRf1mO35qk+1Yx8dS592NQadM0owB+Lr8wvm5DcoGyrrEh
6+r+kKznlY30vrzoOYl1c8k53t7uGZo9kw2qjvgtOpNY68MBLKI76A7UWzL6iVdH
m0Dz2KHLCIf9asCT0Ks07es7mucik5Vd6UzsE+WzmFv3Sl0M652w3c5k2ZrnRVGM
7tzBADB8Z53yYQ8E1fDlU90iewVcF6p74563hLlvXtxvAokstSgn/jVjsUQHae+v
CU/0aFSRT03jhofrlx6QwePnCnfXagS8BPox66Hd8Q82Kp8BuriS4IQsNmJiMM1r
WCJcKcvCW1O8jEZTpU5LFBFkKZ28+YAgRNc1VPN1icLjXod/TsolU2PnOhwYmImo
J4glYjarTC3WXQv1J0CEQnizXrFQvoJgGgFUMt5ty5QJ+zStHD/W2tSDPDcfdPm3
RhJFoNIkENcIehLAVuQUb4u2ZEx8KqFDqQUMUTA/OOLBzja2vxjXy0AfHrQ4zoaL
zrVx8KDT6lfY9jys4sK4EG8GWFvFOP+Gq6dthOFzURaIPF5WvQKQqaQPD3RN0MDy
nV5dt/2BhLASmBfvLJcNoa6moo0O5qsBBpxMn2cH5X6KUcNuFv/TV3kpW4R6jzdF
VhPfSVgno4rVuaGA52vkR52gCijl/5G+nEmtOBir1FFgx4ukreuPVBgDl5KIIAwy
WbopK8ZisGRbC+0n6hzE1mSmxvUeeDmWaMsmVywjfZH8hkGseR81kZ3fAWCNC9Yr
scXq6QyHPqbF9DKbpHNvSCWM/U/0eThECqmAgUdKsKnb2UJ77qRcIsC9vLmJAW1t
IvfKD8KFEt6G2nIPAi4HrEgZTyJfS6qzUgTRi514KJQCeBBVQsZEPHydo8ifoWeG
Bfkd4c3z6DBB+7qnZGOfoi4M8Jcm1cWHpfk5ev0rHGexUg9rQEPso2+KxYbLgzCH
Paw3KezTcbD8v/SNEB3TdDerC1nvjJH3wXFphfe0mzfRxoQmiasPRPbWepkyGY+v
AbW0hjypTcH4nphQBjtpaBABhu/nb4XWi64tTc0mUYZeQLXIPZ3+CF6V+pir6Itm
16NnwiTdH5D6KFq3faIbtSEOOW3u1xGR1u34Kjd5QMPgp0zxbjsyzoFVVCySayvC
KA5WvMZihfqvVo+F/ZCCPod5ekkQ+lpPmVtrgMylwIVEVncyQV+nmxx4NlRezPJS
vjQ5icM7iabrh9RpjDO7B59hZwY8l5+vCxUYoQ9tGWrXRUFeQywPDqacIJIEoYdg
kruFur9p6HuCohrad9aNKONjHF3kTw/IUT53A0mDZN2+s73Z93NLjQCA/m+hVHfc
WJMFCy++BvL3l9jC63JWHXOlE0es3d3+ogqSeHDn1LRUogYXApgNm7oSpwLHS8IZ
xJeMTWM3wuZd5P1NQkIphsTmCJo3SRicU+l+oVFWO6vArJ7C85ynyX4sHuK6dxoX
Qtn+qWOU5/UsNVJF3Z9RhGCkWXcWjf+XC5hQBFiWImJhLR1KxVdaCCfq0nXyM9+J
tUGn7jMlvl3ZcQkOffDqJXgeFXt7LGGVeJ+JruXW2gNQWp+AdRTQg+MfZippjqET
0g95uCh7nj0o+VW8YQKQAlP4rsz/MUzOhZEoKuw2qJnw2E18bGVhxPHSrV42qzB1
cPHvfXv4PnvYbPYGaq4DVDYrsrt00tdBj1NuXQojfGBDY6j6IIhZsSQxTPiETz4v
Z2EbnRo/8pMEWiYII97g8a0VZU0b00x1gSgDOu/D1pGBlmRlmt/Uljq/Aw3dNN+S
HHP1+1VZ8UR5Uea1wkt2Trr5xzj0D8WCkcQHm3vOdap+pHI7GcZ/xJsTz8nUKNVu
laJVHnPuO/Hc7eNJASxDQNQGPVg8q94zfkC/uIJCHgknCRK+0BUBSjI5WrNc0vgT
1yNPbsEOP44PyyBx1A1aYx94+zIkE313kO75UDYqXeBDgZDWoAgI7Ye7hTzCaZgz
jsDOXzQ6Ohy8TTP34QiL6epV1Ew2W4bYMdeliQZ0AA3bR4lgA5IFrB+Amopdk/uD
QeLmWGL8KBX6oAUygGkvN0F7dIJN+HVGZxlO2cQMJ8xwNwR+ZRmeKixPK9HhIPF1
DDks9F46OEgFJgSIPAYvM475TOZoIGXg6pogiLK1/TuToNgC+YHP65UkqK3XejJT
HohRBkZyX17Fkh3dh0dtI2Dw1z7TsKjS5uk2MOMGm0emjKhFQBWU71ZbnTKgPPTa
M9NFOuzADj7G+y/SThqtgCDveBlhpFhzbHzxzq2JhaZ0NEIi6kyPy1fbE0+72Rgs
XQVnpeL/r3BeZsL8e1M7Ksd29UKJv00qGZ6fTffbAYFQckNCg5e1/Lbc+qW2q/JF
9mHes+v0MEe/nZXY/ygAGUVkar6TuRUKiN37glmbMMxc39o12IPt+Rce4HDMaMU8
fCDB+KT+yXFOBWoJO4Qc0cneU1TOo0X8VMe/R1NtkhFRwA7AvcYEUBvB3m8XgIiz
KGCwcPZHg2R+fLeG2muFEcM0yX8Z4o/5iHV57xjPcI7jS3N/Ou8n7BwBRlDmq2UI
t7vyEJGFCuSFG/IY4L0HRE/mpFOd1Bfj4SoYS2/1Jr6HFtbCM5jlsd9jegFoZEfs
oU2xyBM358EG1Gw4i0hgmdzVxb0ibIIrUM6uXoTc/heQ6nqUwq67aDOKoSyBhVaw
PvkNjn+bNjdMPcJRNfBMs0K7oHawhQQkeW+lAcr48+fZa3PGGNLt0DzoUN7CCf01
g/zVvjtyHscwPX1+8xhYM84GAYG+YgqKi1yix6MFESvzHolGxOfonbJ5gElIDgP/
d5lfBayDOBK1GpsKM00c9d2ySADC/xW0wNHZg4R5nmG+mWj+Z+x+5zgz38zRmYgG
yqsEon/ax1Ccm1GkKrykMMw3puw2wxTPVeCYhHZmIARaPTSb7/KqxWDR4g5HT8JS
SEl3csHDdYSWz714TK6LEb67XX29ckm4F5ToyLg2BabjmAj4gvLF8kuhCsSqS0au
3wbNnl1y/ERkGBhR+bqKt6+qz/p3BPZAjyo5qCLoCK4HlTOSNfAGsoZHMNzoykJ7
U9nTsmAyCkqvvjgstcHtGDbQG6I6Q8j9VRKqBhH9tPnBsWAaqZMMhPHo5+OwgXbm
vXc94nzY1u+9rdIM1D2HrlxI/G3typgWtyPVYxjc6LxQlKedEA/9USVBjfhEuwPg
AH0Aye5xf1/pDZcBYmF9OIuFq8YZ/6kqwvpYJ8fm7VgmjQNse8jRiOSJAOrdq7lI
vqzm3RUKi+6qd7LldpuUnhF3KjMJ5N/CCBWL1ywfroAQYjnzR8FEZbOEn3SICnZ7
KedONPWcFHRkPn74Yc71O2ARhj2r2i9OvGSkkGrpPjXiin5K2BhsH0uqQr+UN4AJ
9IaEKI7gc8Cfo7nywMpU3PKz5U9Lar2Oav87QBOoRDsL+Z8lcDvftWRUyAlQoRE5
ES9dljDu3jg4z+4guRZbzNDywE0u/1Qx7pBTyvbAd1YiOENhfGeCW9PtWtTB5JkJ
RwGlCltkqxlYAxWtpSIe0+HNdfACGM6Qll52+uAYSseZ91LcLWGFJLU/IJ/M/mI/
dSpoY0HZIgGoidw7hUy8IykuwQ1LZ+3qTdDBXFTq4msC2JBs5/sRmD++C9vKj4nT
3shpDnmuEM/btxaWMWZLjMF2uCP4PbuU8jAMkogFIO1FVDLE/tpFTrX6D9Ml6FXC
pQkZAzmMOJAWtoHtB2sCMB9GSNYgimXNY2vC35HG03JM9DvhTWdU9YYYwIRY4JcS
z7dZvMyeM8yioWqL4/yG3AozDvIPV0eYcQZtrUmWO7GwFfLNDdGcxBOHTvuS/Pbv
w78dQ8XPOmAzc57rFQE/pr3K33QvhSZhPLnrpDFqe7d4RdYNS/40+qpbd8PHIF79
cfwrYJm9kyZfwLTpal0JvnHnl+eeb4/MjMesUdIMQPEtNPEbaiwgN/+keV/ReaEQ
QYcQaHlBjBr3jDrpBULySM4/FYAHQFlXMG/QA1sxiJxvFRbj5WtkP8oDFdLQg8FO
w8FI3WntHlbAWNNWpMCaNeO04iCag0CgibujcFKlCyOP8m4yMT99CUlvIwYvGqZ3
6wNwU4XxWo6alW76m+ktz1rf2ayOMPdl4Lc/iJ0T9erPtO6+gALgiiiFVIH8hicF
H4Xa17gpm1wrqEVY9GDV7EAZxh6girPPJLjO05P0RYI6OGinvaMaWjcINMOw9fm5
lTNxRpMm2Rsyb9feb0Rvux/PYgocMJim7ms9Iw0lnEkXl3CWRIjg3unQRdjG7GID
/qiaSFlUTqsIHqB/VrYCy/aIHR+M4Y5vN2O/6L7RB0iGliOeDJO5gh4whgYTbvOr
XQkqqokVlCqBmlwZVrJejSUeWipeNvlbNf7b6d3LqVEQRyyAFNzfjmpXvfZKImpv
gW5RVuLDFkRfvp7LThzCYqFgf/VlEjSLkPrFXno8uda9XB0hBnGccZKVsYsOJ8Un
wfrEQN+nxJYYrZof3EynWwoF5qWzCrtPzrMyg6t68fP3yd4dz7NUH3yw/PUHaw0S
VJv+0Xb14Tgv4KenLS4s484je8pYBd50nqDVH0WyFDfWyQCZs0ExSJImyLU/swpr
7skPeP+JPA5WCRgdnrOLWADqWfI3fESfsSRj7LN7VDe1GqFNO1HxbWcHuCFO5b5q
YgOU155+h/NUV2lDevwDOziy4YkroDHKYmx5TRRjf4ia/drL0KtKhg4ZPBDaPy57
gWmhn4lsxQJtObtTvVH30RNBBuccIAeNYr8qP8MsCveJVqst/IQbPstqnKfdoeDr
XYmH0kB2wZCkzYxWkCtHeR6UHykVOb185q7nKEO+4XXp1uE8s9qbP6xqKyr/bhC9
nCz3sdA2UCpSJJtMXbPipDk6Uzy62d2CEuGaS7F+8dbM0yY91wC532COGCoaZOmk
Spn+wVJUhBE5bIrgOhByfwuQasoZtVo0woo3+2xOdUaXInf+QOnFt0B6vc0c35TB
a+WOBVqsU4AejRk88anwkI7eEHJEt3XSLCIkE6ThRBFeGWFjcO2hSUUCaAr7tNH7
9Dz/EIMuBKOCbFTf0Vhz9ZtxXDt8OD+omjz5F9EuNzlvyC1xYQfJhlT0wZjiTvEm
QwH8DZRE97FLgjn16Vd/Wh/HAQ8IrsJSRYDPQBPzelbVFKIw8MIDmP7HRq5j5wfw
ZhNm8Z71a0Q+lSlcBQUoj8Yk9s6IBdYVxstsWmy29LM9enqzrtWCM/9EvmlvWJsX
NOAew+F8kJt1aNKYQvXN6/8AisDy8k2Dyd99HprgLyh/DdlTPOxZHLOzxwhISk8l
/3oJorDgK4VGuHfveYJ9jPO6zIBwPOw4/Zse72R1lK7hlqeBZwnllo2O1yOzYXPt
5Lxy4M4FrK6bn9v8e+zrSDd/U2VNh4gJCOjG2XMlpHEZRMFPZ+FEsKW5bQkcf7t4
dZnPOv0w31KKsE3mCy+wRxkou3JSMVKNOe2lXq1qHdnBXTymxemBvPMx+yF3lGFw
qCW2lu91ek8UiKLUwrln8dib8UNT1Or/IpBo/S4SsyqV8H7Xtpzfc1RS+yeDMxGc
uhJBjA7m3RD0zF+2IU8JS8qIZm/1J/iGSiXxR5MsvHV7JivIaPUvMWYkEX4PfZP0
ZE0BX1Qqszg9VOLVvtHgNg/p/Zf5ukrkjXpps6/EK/m1s1sIAxkCgnwOQaLuBmlo
mjAazHflUpsw4qwGLtD8xZ1Bw0KWgnOOEJfffFlzFjZwJAgwp4Q1lIhuxlfy2rvL
ijTS71orJ8p8/B9Lq8pOXR9dKSyR3QbDXno/dDureIEWrGqdIRch3ZvzoCPnphvn
6vf9IQ/So4wbBzzpAQx5Kwk5flSKWPKSI1SNgAJpNzZSu2S2SlHzKr7b3v5waJQb
wa55Qehsq61NUvPmjitQ1NN+ICzOStLx8SAeg727/YjJKx0GxHU5Xl5Wim9kiAca
Jk9T5XokyI5H+kGqPuDdPtnr3yImlKhyXFcF5f8T8xGDAZbpqPa6uSsl1ODm7AW2
BC2KbFtxZUQ0NjVI/5E0KPCT52Kn9zkGnGQPr5XP9QdJbJkcfjmESy/hbNhsaCtj
AEOMj/0KQIQ1pnmFsZ4/aAWtm097/fEcGZkdtO4fX7RW4VOrvqhENCg4zzxDqzfO
or4u7sj/ONwEVZLqzLG6vBPETvU4gk3B6oTSQDhdMc97J5fpUv16Z/SpC6F+/nBM
7EAoj3nCI0ZXHYZ4wdzMwgZ+ViIh+WIVAP4BYc8WeAb2SvYDnAlWTQyf2zZA1ecY
raKQa3K2wdzIi09PVcIj6pvFriMv2xxxplMi04HlNvaqqnUoOD3NuCxKMNvcMAOb
4h78CVMN8qtfRJBgEgXbU8OYqlCuBjrgEZPd73i8ypZmA2p25arg0E5p/rmHb+tv
159wUm9Ez5cSNzLqknzDoEby7jy55KKRAmlNbj2AhJe6QUacko6E+RTsLux4LhW/
UH5KWJeW9CYCpLL/O84VpbnlzMo+sNHl4NfoCOp4useG3TVKhGI8PMWkq2kf8hT7
LMcxXfUCCKYLKLngcaNlDu0aiQOiloWiM2zpj9e+HXtzJRTpuF0JIBwWIV1OoGeb
n81RiNygWbZwBf0LetWoFbB1ooE1bmV25aIJU1UBidoaWGRYglubasv9ziK34pEi
BFmfQz7nOy9h4ts99+E7G8S3PEVagKJ2HvsIwkFXLP/evasIJaxgLKXxNTbHXQQg
Zmei8NirO5ivVnSSB9L1XZNJIHqN09O9LjEd5/hJTgKjxHY1tgaq/ye/g/D/6O53
2gUSP6nOVPYctgYNuTc1aKLngQLEMmWzAfhRc0KLF+aCEXzyS6mIagt44IH3BlV0
CNMu8ntrh7gg61UiOLe0sXsQoQ+6gfwjZaoFDeFSX5wdRdo/VR3tbNWDkiObb8PR
u6DqTaZHfWWbDXjVIYnoHkqpv9WO2SEh2vpVNRbkvKoJTST5HRCHWPN3JsRZGKJ8
lDAvexODIa25dwc3NmLcZOkxywOuuFSwqMMtxFpEyvzH8EMFOyEPmf90kdgLhZSV
a7Dj6zVXkCSuEGuryfgvD8x8zRZoh6wHoa089r04xhavOWNjjLAIcwtXq89bDmiw
xjH/2/DFCdYtskYCotVB67Gtpl5lLZ9eH7Rr3YLZEAP+7t5rSf/ERfovFleFQyX9
gNw9mnn8gz/EAn5+Uc/KPq1tAejgTknvLnHhrayxQrb+cLCrFGgj/4Vpo6rJk/BE
jbyf5WjrZp9TZInzgxNhPlknHkkhW6PBDZ4TXim/AwYgMRO+apND+dj1zL0f3Y7C
U4NinxsYSbc4JpylfZDN2yT+yHhMOhtySVkssyzMpb8/ZxYiyg+5Q1EvnT9ZfIZI
7paEqyBR+cMkqHa4Wz76Mq3QifIELiyJsXfMpuNFXwl3IpQbpLGUHb7xiVaConhC
qmiFN0qZZBsOmvmMuAkFJFFje8MpAE2xnMyAQXDsmEJJsGcSndEtTgqfPz3BtpAi
4ghYDabpNCv+4y8TpNq7qapFeNfEUgpZsgV++ILnq6bIrvhOiNPit/P9KfCrXNqx
OytktTjJ0MDm0F0K6XW6qpyXlfr3q4QcFGBK0unxXpObs1skE7XYpYtqp8AU3aZQ
Oc3jxsxCcdc1+jHn27HZqJOo1mIusFdgDE9yim9nEtsZOG7iy/4Rl0Y145rPDLd7
uyIiJylU3zE8wmJpSJEOqFr0uTNXr1YNVlhrYsasLMGrkP+2CgH/hAeYV5RrNnLH
71NxUl/cuNxD78hqWd2ApExdYfb86vqqCA9WMZHNVoK4oxqVum435ujSbaTgcOUO
UUANyQvkZo/Y605fFTnMXwWNy3U4AqM7rX2VlYijh2fJ277OCJ3Bp5Z1XgsZtRjU
zLIXXJqc2kfMs/TGb5ymXujYVSTfaKmFeg9zBdd6XiRGBsB3r5bm6qPiLNrWB4u4
do0jnyK2gqIm38yhJt5gOziBhq1TL3LxRWr0xEiRE16Nw0dkdkKakyxDfNHu4PDg
bRGIAdIwB3ZK86adZSdLUQTnflCm5DqFOrle6rV6YXKOEHp00XqTVD5CgEJN+BNL
g4gefUbetrk5xcXHK10lfe62OujIBGBbJRIIiw+QwfeDEfaWonPPuO90dIWAsEgy
Zwo6kLesBN5bM34FDcwFW/N0xj/nWeKUIPgrVn2LzMYXLY3FUNg8Z05aiGIr/8Kz
nkunTkfrN52WyKQWKRN9nZBScleE9mkrm/ssTC9Nk25YLxaz7puLKxERzg3Q4v3I
bvWABYfJ8+kdbd8ejVLRx7Ojl5kamui6eWGF2m1l9pA1kOvsSM2yID1EZsR4CV0M
bPkViV0QGg1EUbfjWvejtGRvjAviC6mM7o5nmzqah2RE5Afn2TrEI8BCwL8Q2Tea
DpOaVWxdLaKImzRYp1Dkww2wRlcScLF3MuM8JqjXrPbeOwgebHvhIOMWlN9JkWlz
eZdUW+S1pnr5XZzxydU7HsvhwOXBZinOKqRhmAMESZqc3V11dpX93bz1AzLnMDl4
k+4mcjigRiYSoBWx26eCG3bmURAg/jgNQWXQY/PPrWc0jYl2Sy4nh6DqUv5epXSR
Q98k7tfkmQmXmIFEsgNz4u83M8irVZDnzORBecVrg58QPaaJmG3Kkdz/Mj2Y1vbC
XaoBKXyMibaKIBXVviZZtu4NC3t+azj2QagYnT5W+722pGcNBfxMTWw6uCJtweSk
dJI49dDGtbYAz9wu1IJK0dU19jD7yt7xUAKvDeE5/EjO0xKDnb/kbx3tcSLtUvaw
DBe19oO+esyVrHqGDcAdkPbF2hy2+Zp6S0zKzCQVQWeXxiTsMvJ6zWnDniGQeGZn
tQMsYmA/mrTRZRfMJTZlpTGlp+PlGfpuebp3ZdQZ24hQ47Q90YP+uu9AS7WWQ6GW
iQChY6xpDw7ief/5A1QBcfx+1nb1rwcC8dU1FO8T+YzZnB7vjL8nQcsAbFl5XTk7
zg4c5zgJMV0DA7vPgD5ZSkLErcdB/WPXetCsvo/scPL1/sKgxNcF102T5zKZBGF/
5bku1759wpWHDmt1MBlAxe/MRTXZ0tcZqXBHdEtrHS54jv7459Sl16GMHFXvRYqw
je1IMODw5j4mU9BlndBJQG8uDobs6Y0kEXEnz997RGWTOpgSr5vxF8ZaC7eGrHBG
YedmunMB+z+O2Q7OB4At7FS8bci5T2p5UlbCA+AAhSEOgGe0UKHZkgr//rYSDDBg
83qOWP+UDm27t0LMUB5H24FvJH6ZYK4+DBXM4Y/joNBZddPPast4FLZs9Z5/WOmg
ymoVMbT6c12usr9CWLaYVr9esaSpptMOtJHotkV2cDXj2SyxVb41z3Gsq8gf8vJN
C0IEwZwOSssctyLvEva9wqzB2TX400KSKxKUwYWADevp1WPAv8U4zkq6h3J2+2RY
OpGWz6YnkEWz2E7L+EvkluSquwg5f/v31chq62Yl241PEHEOex5kyKW9IscwVkAD
ndbHXpqOjpHLFIENCk5AbFUo3SX6T4HnNaQ5LBqPp+Vq/B6ouDUx+XopR6MkxTzX
bUjC4+8lvtw/y+jUy/BqQEFXaYNBM9t645kCGKCr8sTo79bQ2xaU7GQp6cTXsPfs
P2rN/qW9kxCcamrQIzM7JptUN20kPjke510DonQ3rex4JyoemCqdYBNHkCLdrhjp
vbnb5XyB2XtQEy5WbeQgxfNCsAwdjawuvX4G/skxuj3ff951D9r94cGhfNtAZpTi
D5XOunO6ORcYmmFbezkCcCIrZw/IE4ct/vmDD/8mY6Dh+xvtXqMg7xWvru0sZ88x
4xCHZOekp/tpYo/Qpde+bbFmmMZFwo2bn4YM9LXyQbtSe/0wTIi6vkR72pbzph9W
50iRTesYC1cfNWlRkJlapiWV1XPnTJu9p7DseQy9seeQ0i6QxGGWdll6oNPbS8mk
koaEJ5VDeDC3sILVlyJKVWn1VDhB1+h/cKROGw3J2L3EPEruDeK6C5yLIQcg5fo8
3/ODOHQwSJesm6Ob0KBq717We03kyE18kN8GLrJ65KFRuVx4xYIhHiBge223CG6L
+FU13AGFDl0dUYkYEB/LkahleCPeBm697zg4rw+B9blNugtAIBmkJ0Yx8cbv2HxG
uUi8Ygu9NzT+OHSg9TUrsWe7mX5Xsqy1a8qv5jeZso7nyLIIXyIaBquFCDDGDLGV
sJhBAocOSbc7jsVS7rxo9AmSoCflq9Pl5FmxZzVk9hQyoeXpYnUkK+mwb/6/BljT
gs4gJ0PMvHfvfsWqyv/g6wwpouC/sf/KIOH54AgP8YAjs72xPgKWqs2eAfgrlNnm
1+H3X5TuUDNbRvxJtrCd5lKUdp0z6S+luXdhh4T/E9fcLBWP9l1k8yjCwNORneCB
giztp9vf3FMDgX6f4dh3SaESBkdPglrR8oq5l8rjsPi4+FLjT/FtzVs7J+tGO1zS
YHyepMO/26T3WSagOflM9NxgJNbLMhepUoyxlFmgCJ/gi1tadejCPSXEX2n2Ckry
of5Oq4EIx7XwS37CeqaTB0z6ExrjfNEElPLkUes+R8wtLdJIcvCn9UOUaQAr18p8
9fzGRgWo6CxOUXhOrXWt3fEwk335BzF5i+IOMSB2NuemCNBHUsd280m9f9voaZJH
JgUaIYtGScE9BjBn/JqCoT3Mw6dOVehX96SudGhYRLPUgX2J8Dz1i/bjyyF1K3jZ
MniQ38Xes+vS7gn9qDLTpu8WkQCIc+GVcBM4LbQCAgGlei1ipF76nqJR4rBs8myn
OxLeXNWxxfx0AOx6LYu/sBKjuhWEZJt+U2BEYDdatDWnfjEMwrnP0WLIf67WZy2t
1fWARRn0KLxe9PGao8Z9MWcioVQyPfrt/mBh7nSCwTY3yLmYVq6ylsB8z2CXJue+
CI+bmSLUpfid9HdGke3jLwoLGosVj9DVw9SttDxRjhlS+7ocnNNf4/Px1NnQ4Hdb
8gjO1WoWxG7m30It+pZgNOkXJMd7Tf6QCzKILYIil6yyFNJrabWjEgNc6EeaemJo
2F2KBj3OdNtAMoNncksHHDgJUifwKuylkIiHcsd+0V7ddYZefLwlXxg6uJfqeaN3
rXAVfjuyhzQAK0nzMFNqmu3JRi4KEC0Y9dubW9LjkBpH4E1TpqHU+6NHHCaY3iJt
isjZ1+/dZUHS5FJ4HWTxF+ggcARf0RFt2uAdpYwKrnQ+QzQCHEK3fiZs51a1JpgV
tfymFa2/BS80NSNK3RIJVNUhu5ev9+MPs1hmdkzDrZygqs4Kg8BR68vUmGGmisQg
8Q67M1kZSLHRFaQ7e4WeLbVcsuI2Pchaf6ZmR3XC+PpS7C9z1qY5m5kvKZ2mxraq
lq9kTUgxEf+WzYqTja48MZ0JsYQbSbSvUwbqQH+6vQc/VL7Z+u04V36Tc9v3rqda
x18VWgt20Wd+28PeJNOFV1Vd1FEOf/Ff927HYXhTaWq0/54UbK/1KZYrOPp7ZFPY
TNTsPm5N+ii7r9+rud4e93GeZaE/u5qed7B4HGh5xJbC2WqN0lfSPZGCsFj9cJVW
NSVZf/MOSgZ6xBLaIpufRwABKazoD7OaL212ZI5LVqDekaXkJyE2vZRXqL+B2L3o
LP38BHM052/5BxTWHEnQNbmoeFE/ZO0EoJJKliKjkDyDPcrfpZXAC0wZXp433U1M
74hziEhtI4ItaJXMrTiyHPVPhN1Akzfy2LynqBT05hEX82o84YwzN8hTF3LIS0iS
dxO5+VxgX4O/LPMnLmA34T6Y+ZLKDjZGdJ82l7BBJt+UbYf3+CESE5056NE43PX2
L4ZWaapRxmmIlWbSgpd5dtGBPPxL/gODACJDF4jPuBoW3vbQlFx2p5LDs10JnQ8t
MMXJPuNxB+QwAmMmEI+lJziF5o5J2D/MzK0TwGE7xmaxn6P+4pbt/3LKvgTzcmhH
CVyojpHfiOVnVsgL8kOwIYqwC0ESEYg6Qh9zT7zqeeCKR+3piJ7FBlP+47sm0KTK
o93YAEcgOoHQdKpdXB72864STj0+9QLRlT+RrLdR9UQ9YpQSjYHgtuVYA0lSCAar
UTc31zaYeWULVwiLL8Qw9MKIONktymnwpepmJi5Vwsm/kSFCW1yYPwML9qIFchA/
diB0qtfHE8krjvh+SD42I7ToVbRWhkCNY853ZDCF7Y3weKq7t/WAVcpgV7locYt2
PuTMCMPLDvsSXemOWm7N0tgXpuiHNJ0bjndUOjYGHtrUdCV4bbuuSYnmd+I4/FCj
gUrGxW6+WcfoO61ithTVHlDZv8tJpGA2JUceX9O2MU6c0wz6hF7i/n9XtG5bysFT
qFS2w75MP55UK7sHz/IA/9lrkc1B681T7V05FroAesatwgXD3DQ38q/kWp9cqNQw
HkWO4y63GihrGE+DxP2nTvOf6rWuHExAdebRFBg2sOLFNZvNgsLBz8PZ64o4WhYz
Ybh4cWuQhJGjGsuB4FC5kcHR50h5jTq+ek7GW6ZwUgBCVz12vfHTLnOQKwB9h4xx
hQCdLSUjMVU8Tv64pym6WlNsIKydePaf/H3BZdgsR6PCY+/4/x/l9bbhcnoIB2kd
zG9rVbcnx5GZ1VxSIeVXavfBjI2Is6nDHrlaJIOhzU2CmnzIWlwb2CfnW1992ev9
Gg2rIjItp7q3PML02GQ8v+7qrXv7mV+wDTfLf+RXH4fXQmGujcBF6gVv4qRyC5iq
oewu37m9oFTFv2E4mFgLQiO5RxX3/ILh1UA4gz6hpfH51FdGSBGJBX2DFOc74wsR
PX1X0NpWCkLbdXteIw70V0vDzFddjBJGjkBX9mwtrQakE0H3NnRl9EexAx8YpdCb
UP+r9ZkhpKxnV4IocFwGbytz+pGLbHPIxmhf7DUcqxoSrGJamJ8u2YN3x7QGyyLZ
xBB+1D7kuFJseDzOOfRs3Cd6EhaTjqxjlJnAnHf4AEeT1y62Tql/NZeTAFbj4m+S
Ukgo4W4//kmhP9Lbj9xXPntPNJzOemJRmwtoteGOiFto/u0HNcnjgfCa4AqlU16o
1tkVI6Q4c1ucyRSIy4UFnj0yD+mB6omujUJBIfI6/Q8kYvho+NCbh0+m7qhZG2Ug
yh2j/JCJZUUJtSDuY8DeZV/NcB1BUxP8JfjfLJHGj2d2+RrFhGODDyhaPgcuNrSI
UO15spRYbBVOCdvALrPd5MV+y6RyAUCtIEtLrmvB3zp4sJsv0g/PXLN8D3UUeuFB
UNxAeZB/eJJj4kM7OCyXTjGROIdes5r/m70DxUZqRV41wIlebWO0yP8K7OMNXUb2
DSDvX9HyCLSkpP+idPUBxZLgRkua/5iYBcQYoa7/fPS5+YDyeJ3mhjLvXfyRz11G
9VoWm3otbWBmzBAE0tO+NPiQmyMoFOTTZEKflGAEvBvCXUgA9OUyhQPi75FwMhBD
KIu78S/2TaZnyHQxjy5/XPWdRDHtR73faFr+/D5kD1djAHkg/g2ZZAjWHZpN4TIb
MiEsNoDgF+5orlM0PcQM7lBCqODvgp/c/1WOThL17IgZnsoIpENqDdGk7VEnm35u
V/XL6P/vRXBiqUhqq1qYjon9+qNYob5cCcoKfAD0Xq2m59Qlm8LrGL851vdzsCO5
kg+d/mCaalt4SD37V4j0d5Rp55lmTjBKQ/PqopEn8KwfS4n3Cmgof3hTfF/yr3xW
KdRZIhlMp+TcGz8XP5fleqU+Pofmm2J0puAh8Hxgo38qjEdAQb3VSA5zAFuX0eXq
iwND6zGoUzrRxLfVyzSbylHBlnB0wYS0pL9xyns2wNZn72zWTiry+Xx7uRbZuDnz
hlx1Ci3dqyztLwrDMWLdCETtSa9Thl/NvXvUF1q3Yt2mDAff9PcnJJ8WuA8fRiBH
x6fODgeO6zQsyWRcCow/iAkmK8yT/WK3RDPouE1PTmdm3K2ez6li1zPBpcAGas8R
ZZdnqaRLBS9VqE5grrgMDeXFmMpCa3uKY4gzfP3gjmz9KYgQyXgaSv2b2GkI12Zq
ErNHDs6rP+uX+yIzHjsQqUA+FgA5rOzEYoOrkzdSqYsCx/nPOH0hp1UEelJTYdL8
m+UFRw1AswjC/0P3rDskFo9NRQiiZpT8y9J18XfPkMfN6u8D4C4yH7weuaNhsYCE
7W+AFRVowx0CKV6JPaq+FajcXuTKQItlSgOcCuYhEKtNziowncEELwX8TJy4BAip
a+vd6PINzvum9MNJGLAt1e0Im9b42RruWqnL8lvzV81sluWqbl5HvE/Vp/5uFf30
e5ivUwnYC/Ax/0KftDSvUXOvv4rwNpl+gx6eHauHtPPo23IVEqfEAX+lHxEakogU
tM4lgqSahWY/IGqzRmR24LFtgRf3pQ1J3IVHXcU2EY6VgyDWtolqksLlEUHfj98a
70p5JGyOulZepC1MJPs5Se80gKu0hAzDKdYyd4TaxiuQdHLgWjU4C4YMAD9luD/r
QkgPpq3Yk4Y+nwtl0CukWdEg1whMy5dRtGh767IJLdMAOO1Xd3xNNqa9DVY340Ch
HGEQXL0B+5dGQxdakmE4YLGe+htFMv9P8V6stv0a/p7dglnLzHFo1qR7rHEzUyZs
8fQyF1gSAb6kXUzN/W+pl9DBKhKY5WbtQJfMoo2TbIpG0oJ0o4xq/5cz9WcaNwlo
hqS7do9xeszfQHS0cAefn1X8UpC1o+j2tWr1wfyaRpgdUXiiF08cYLnow6LN/u1f
AX4y7WCpbesC0wsTagfIxIbNO92M2J/WILDfu+Un/OrqThcX40gnkoj9Tddg3ha7
2fezFbmVcu/vNq8gXYm6Az4u1cFEl3VlBw0erbRpSM6uCzjL3hztWqYHO2bQqWHP
dFJPBuieFVEkpQt/Gjabc9hutwIowxE7ArrZLvwd8TIIFdbIWWLN/RiWOUG78/cs
VC58jFIVWK0LSMoeQAQ8jebcx1SWZFdLYpOCJDoMSrsTPbhxCwz00fV26L/CHADW
l+Xszan2oDVcJjnCiRnnBe6HYtTJW/MGbX+6w8+qdjGkKfo43sFPUhntR9/ehaDi
xyNhmLV161x0GC9HQQRCxXbE/Ay5LhPDsNbPj9gTczBO9nX9PhIKIG0fEFQYhNcm
fUfLb7KbwrwOj2oiO25UGbrdB/I3JuFbLzGPS4rAoKUK6K0oLYZKaJOt0iWqPt8H
3At9BYYHT1C601QiNsb2PQhYLbsDI2o/RUrkuflIbXbtitVwaKlyxoETMpmPD679
4jT4DpmEivfZQ9CFf7nWTaurBxfY1sau2RDSHmDJT3t0BVX8k5rBHy6UgqLqeACk
Z+/cSYqM4bW8qK9Rg3Bi+7D80k1S0zuFeLvobhjaVnrR80vbIiIBDgk8lqMrtbt+
VSvpA9iANiNay6RHp4QW15JLnN55RcrgzgEfe0ihxk1rHXFvIfTdrp2SfdaaCm0j
5GTSW3krU8OGJPFODlMqsiQLdIc+VXYgKZz2TeoYJtzM/49/eoBDHZ6GZTqx2avf
G909by2ZPlgPxwijRDo1cKtOMyDpKcvJXcem6kAqZ/65v+7j6iDAvhVtJv8+hA7W
2g0RepurtK1Q37DOgn7pf6mVhIcAFxj+ZfP4dUClXSQiSR5IUhHH+RYZtyhuGEQh
ceLTAFSxU0RdIsATbhXlYhwkj+w2UPMe66xqvZyTes0J7nDqHbhedZSOSh1lvLNN
0B7dZ83/NeqSqz785fR8HIEWHiqZQj22QzElOwaCvwpvG8UOePX68Mwg+7PakBRB
+UhxiZUudapC0vGQMvWZjYXdfEXVT3qb48zC7KjsNOwOXesq+AFh3IVsPiwOwU/2
foWV1IVLTmQcx1kTShcprNVRA2mwBsCT9pfljdAe/cp5EdqCy8a0C66wQlDoB2eL
tf9eMZUbRb58+JolirRZbdhMX8/jExBzPzMkeHDi1mkaNxiAHT83Rculm4I6C6AI
QQpR+EZcmPmcVCpA/QUH21Aq3Ks85eilZLf6Mv09Jfrsr8919iT+GYi/6Pb7kKaB
0ydIQvam56ojW7UeU8xF2xlKdR6iYv1Gp73pz//Bybih1ngXhZrTvyPfPg7SL9f7
+Tv1P6m/lauMPTJi3Eot/xnEHXuzDkSTQUME2k/0wr0HowlZRKBUdDaAOQaKwUQa
hiLkItw/o4rPSayiGtRAwOkT1r48MlC8bCWUSxR1umCCivGi6+ejfSlhBwDS9Mzn
dN1wU9RGcSchSo5SxsHnyUk30sOz2BFWjrzpkocyCdHg4b3FMlKxjeZy7Snyhgin
2/Bf99ggi23j/1aD4C6JVtWtYisqJNxLIIfwFeNB9PbKe3+GqD4KSOAPyH75b2fc
+PBcCXbgA/ZzTEHE/dFXNuKO9JfxftCAp6Xjg4y0LEWIVhgDUvrEL9wfA+0cL6Y2
VbFbKNVzcjqJDOCYryIWDrDd3Zt7klnrBv3ykD1jcQ9vDH57J9xNP8yUhSa/Caye
w/avDvjYS3ISKux7t4qhlw9/s9VHjtgngmaXS/NJoe1mNFiZsztNaiLiXfIyD2bO
sCgGMPLdmeUoW0x42oC5Jf/ZnoHKq/HGkG9LWrC+GUv/Z3N2xqw7Jflcyw6WsjFb
6x6u0a9R3UkEAr4YZz9Tl/WBOUGJCV740IVQPNZRP06Ur9+htIGQBQ8lbEE+KJjU
ZDBIL1osHCGvEsTI3KEkeVpXFBZaQQ68YTfBqe1Fom8MAkTjWqWLtbx8IYdddFpI
mopyRt5ozo2FrtlyvfCXTN7AMRwegn+FjctjXNO48Kd+A+XRa2iC/gSBZUhAR73W
+Njx+dN+rqRaENefGUanQd5A/vi0/WLomietpXooxqUb7o60ZxOc5K/Gr1EUUgrd
b2NEKRj+ZKQiVO1/b0lsIRcvBIIilXEnFTior1CHYlagh/XGbOuPYJkPhx5iksIg
raxx46GnnngPPmAFIS9GB38aWSBBq62QJty2wz9qrxQruwhSMt4eofgIznSsXDQ6
cvItSemQVwxceiSavCYFRPPrbpWW2DJJTfn/185bPJ9H9fZxijtspc8pP7yJO2b/
8bRspTY0l4xLoKUq9sO7waeudCZ22/lGFE0noTae19LmQluSTgiZFjXlTBt8CPJT
M0aTIklesc9SytF4MaB+rR/zIb2E0L5+cf32uzK5LtIpHIOSU7HZLJ1KVDvKqVJx
Plx8iXunpg+sCsHQHW92EhhZ8ffZgCuESwEKSoUSVpIPDm185CE1B1VkYgP62UFQ
/YJtgnsXhTqftZQWT4ueAT/YjeIHxB4gIbBhPjXScX4D/eHLFwTNVyAlozT6zQB2
Mz4jTi6ksTHDkn1YUDHnqss9dhgQ8oVTuiqnvh5E+kenbcLXsDqtiowy7EP+ETR1
b3Vt5U4V+BkAHyWxQXJO/YNg8F7Lhl/GmIXVYuTEvvnwV2IQbrfJXU1PAeGkt/HX
vjPZW3cEqdjPT+76KuawY7leVNVXqvKI2ka2TTbcAM92MG7VZ4bAjkVKPJ1LwTlC
SaEiDVEKaokjsqZQ+iwyng8QlQQOjDsybG3suonzcb0pqYcPH8ewRIIzykmcbgLv
ErMCk0mzq5pDOLRyidDkO+YjOah7MQwKKDhOsVt3wQpOdyhLHNS4OYDwM/IZ+9XM
QJ605VRIeDJszIbthCL5mHG2Puh8VFIxroMymeYAYgx/gEs7NDuMn22gOAiUQMJt
uYs/A4RpAYXS/c7N/1koPDDWpNkA6YOOCyhDUGiGXxhE2m6tDfPXtCbAoD2Jwfsr
wBjtSGjdqXW/0P0SAUNylD29zELYgHxv0FMyRZQi+dDGhciMk/pTzBYszblqFdtI
AIQwhQjHXMa0S9ux4F5aGGlsJHl3gZ67xn9740cQRoKKVszLSRdsHmtVJUmAMiF4
KpEQL0UcjNf26LhuQ5Nh5vj5X0vz5eZJxJWJVRgEYI1hFKYlGS0tF3WgWm9GsoIR
8cQYTuutyC5uRs4lj9PJQeb5XQGxVjj2lCyu0lyx/7XQ9W2jJoZA0gtNKmav8+/i
FVTUVNzDCrtcDHTrEe9rXRa2lS0By1jlkhHGC+SnOOJ9hbGmp31gFvdpbOxJd2Dn
yljcIkr7zMfP1Oo0STDI0vSIyX/VaEbhVcx+I1C214vSDxN04MFPgKdqgkIgfTyC
XW/braXPEv3QXRcbzrlLJYFR9dcXo2e0fUXsrqH4XA/LQkgeZbNeuGx2/92EUS7m
qANkvfGSdHJfqP7hZt5epphF+pIEdeA0RJr3gGW2hqynp/EWnz3IpXEJeFnyFeV9
amLKCX9CRJWtAZZ4vKWtCY5P/jVtMd+Vw/GiF31X3rzeHkEnlJy9o1CMU8k3hpdH
FAtSwGyq9B5H1J3zRhS2Hbz6DUbHuTD1JCZvrOf6WMOMyS1oyitYbnMZ3CyfmA4p
af+HlTpOgCSWppSYm3fMC0ZpIkh3mrutYjCS8TJOeZ7Si0iDNyHtg6fExLuPYv/g
Tj+Gc/4FWt8rIi+3Nj5Vyxe/RmRErbMOd2fWP9L8lmH3jykv5m4Q2DAyKHwsbGR/
Gwx+bz2SqSGANGgV+XkG+N3+1z9BPSWZ1Wv+7yawtmRW3EbbYZlCEqevEYK9Rb0R
63q2ZvfmNyf0vvdBsrxgNYAY5273icQJOUi7gmH79/QtQP/7yFxomg2oYKerSYVq
pyVejJEtstlTeb6puLgsb2ZNg6lR9tXgmwnP7MOh13Ja1c5Pa5YGHaFaF2T4dCeX
rHZsHND7k/BLXzmhHDVgtJ8s00B7SuW7K18pd2j7pkGF424LeWm43ovaY4OyqLSJ
XC/jRGEyf3zFkwMB5As/pSQ5M/vbwXBAUZtCEvOwGbURTyl+ah6MPYbCr9OukJVh
WmTeaYfstDZ3xJeJuoM/Da2sxMIcr5m1c4djVJHX7FaR3L2XaE0SIggdf9148SWB
lUnk4Kq8XTeDmaa/pSKtk8calbdoyxGM9mzZcXS0ZWLvqTmpHmE8LRAX4fWOWwkG
k1cscQWvjkhiJyRa3bnCHpBNKWnvMzST5GZ+lUcm+eeQzbu3DdBaeri8WZIoZf2u
eqt225mxI2skxvKsdzs25I3CiO3TOaWq+cXmUYuc73Y4Ry8/hj7Q2L37j4KMbLy6
UDCg+CMZLhjnPRwI8By5edN6yLjIZhwR0Re76HM1/9oHzQ3Vzz95TxeUCkTdOGAQ
9KA5Ii9XuYCfAxJ07astkXigZb3TGzTSpIvkSxhacW3/SI61gDvbpmQl7KsP8LZj
eMvkvm+nr2P4WS3BzR4llTSoXSlYm2v3zGdfgGYuqFLojXhr22hMttQX65R74XU0
3Pp279NZkuwHnM0qvToBWTe54jpS98t6cGvBeWqhhCj/2xPf76DulvPZ3nAiFwNM
ptvfTBmz14btaMsOp3biBcRlMOjqDlYGDM1ei+cpnu7qEeiEPXrcSYFFkBV/VD4W
NM9ZWDhfcPSTKeIBkGTzEOYT70zsAYRcvRh64cfGyeRf9no70zT/g/tfDXebdnK7
4yqu/GN1FLA1Li2SatzjOsx9eT9I7SiRbE9VkbnE4lztqa0o8yFULdKlDYUwc2Rf
Ld3z3vaRCSJssRzQ5xABFY9BjRmWN8R67MpFsOKcK6y8LvEOAqAZjX6s2DpJL0Py
IMkL15gfXoj4qLNs/4aZKNCjDhu3fvl1IvYnVQzjOJEqaB8YhgP2Vpi3tQNWCvH5
HfxXIw1ApSexNBknxSHQC2dut3LT3cZJtCwJRWxMLNfPQAqyPLqJhI/TwPougSdk
lK614ggfjWQSLQkKOMmbMSi7XJcdD2bZqfx5HAkhn5yj1r5jDQNrDeic5Rb/a3Kx
lBVOf+RoK7DEadGdSygMRLu5mDCPqNUnrOdjbIG0xPstzbFS4OH7j5U3wsKtvb+G
j+2dFsD8KNLaeTzk8AV20C0RZeVtE3Vl7cNRaqTcONG2rteF82I+j5zt76UaAUbQ
vOVziEIi4xd903OPeaX83gIbnvFgjrl8p8z6seSi1WGbSIj6F7YCbBLGHyFQQ4/w
m5bpdco89CcXi/aoU/yga2hq8ykMKcAZKbdY3XSju/A3TsILna0c0S+H3aq5kW2D
ZyICsAod4kq6BS0IqnK+dOpedb/pv+m3cmBRHBskYOdCODeK8djoi1Vf7BIn4Nso
fZS1dYjJnqBzoptmBPzZOVuVCdxHgblzkRWbZqbrWEm6z0QPkk8TWeN+XstymdNf
Cq9KXIwAi8TtuWr5z1QBrDMef5Ho3HNOMA/uS4/EBkaSPcwgXLpTe1SLRoJ5vSrh
/R4+B5yOShNfYJ50mkMYchGd4ekIjXssZWKyxNNjpn39EsQiCb6YiSa0q1xgjx12
8b4fzGl5CNwSHHqWKxqiUcMHOcIpAT5RHJdruMVywqzvclKCmdYq9NRx4BGElrXA
o7VCP31n1d+7Jcp/0EbIwWwDpETMKhntZe8iZ7ZL5xbs+Zjtq4n9hLnTZ3uxPgwI
46l6sxopGDfSSqy2vFbGsz/rLuxPv2GfwqlzGc7C6btbfEUlkh2uX3W3dQbXIo1q
/qL6QXjse7J8XGR4c6Z/VWtCy5AENT0W9kup/2i4RBCzUh+dbhFu4illvv59lHZw
4KLXSmh7EpoRWNbLlQ9v7Ju/js1Lzs1iMvvEc9hhyneugcmm6USS/xwVSIKULb5U
yrSPrM2W+VFHVNmozennPRkG+p4qYKJSUUAGRSrjJxo45NwJbVlys1PTlngtNFOz
bbpXK5knjtMhdETDbkebOb8dPoSMXA9ta36F/GXjNeX99U9hwLoBD1rZwBdxmKRP
2XLnNoME8h/rr3sptyh/nH0fJvegrYj5/BNKrj+TMi7DrUB3pAfo5HVT+B7bqrhu
pow2wxYnzSHsLr5VrQbK73iOhUQh+MY3z4cldGpEeWatigCdqTDqg5u3VDuaqsqi
yqiFDv4yRGzgNQNm/8ivxXLgeLUWKGfA7hn3kBCEk3goGVMD2b7VLxE+K/gYvaUF
NmJdjMZMgz0q2ABOphYELNz3CIsnQIz1H+FoACws9+fbHBEfq7vTnozj+kLKGPJH
mGcPCjwD3i/7IhGu2AjH68gH5Jbhgm8YKyztkcDUVNWgapF7zr2jCGgStVzPU2tf
SxjcbcmTxGTnG5OYQ/9ecwu0Db9RR20M3WrbJl4p55CIoNGwb5M/trbe+b2ZYf5f
HwGAwWKamq7pmBNJiZkFdFeSl2JgjBi56WR/ctMUxJyapyAycsrc160aLz2IVDiq
QUX4vCYUy3PA/XCp0wEPmQZ50uGPJqtoYMX1SU9IAVs=
--pragma protect end_data_block
--pragma protect digest_block
cOJ1O+qmVR9IMaFR+vduhsMjyCw=
--pragma protect end_digest_block
--pragma protect end_protected
