-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
BSN1Ilf2lRwh9Iy1Yjl+Qf1eROQfI+9IWh84rrrFI5fm2lzBzhdfEvYsvTLAJStP
ndoDgk0u5bkaie2A5TDgQw/xvR/+/7+27WE1EDLpbIvzNXS6L4M38zpgkAj8oejH
yvpBPSg6EHwwzGoiqM9S9HJ7sxt3fotiU6kl87OYBDo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10471)

`protect DATA_BLOCK
NnserQOlD5HN+i96wfo1QTGptCR+46U9SiSR5FkGjgGOQQLVZ/SbYOFq9l5MtdKb
/aGgfGYBarZHb6+daiQh/jt6J0yR1iAP73/fYOGx/e0rZFPU41umtB08zw4V/EB2
YVkXNUzLYJ8SqAHIZL5dE2dFOLvcQP4W6W3tAZ54b1HYGdzX4fIuAFbCt5rnYf2w
C10yQSc967hK5AeGm78UKmqyqDj4QKCkKLRHLPOSR8kqKN4ATdqCZTEqBeR57fRy
VJMz90bKPveWpHdIfcUhI9gc0/yZbWogMcE7hZn/H1TlNYI15vgoD0rDOK3dr2pq
ejmPVzf/yfVY64lwV2GYefCiAwmigUXbd8Flss/r/yOVESOdFzkKSHkNZplC5dcn
XfUAVENyjytcJK5dKbD0DK4Brakr/fnXZejPHgkxcoQwwy+Kcno+wz6bKsKj/tVu
PZq+apLcGUFcamfFy8buvF0Fw4x6s8AplEXNnDuqZ2kO4dVfdG7h6T43DTbB9YoD
H/QANW/aFqnLvQbW+tvlazwv/8ML/etsKOCPgsAFB7xOm8O8iSVQk0M2l3pIeLhK
6/dVdupex1GbUhVJZG2ephsiCjF0FDPE77kiA5rGgRYKamndA/AhNIUar5ylGAoM
BdJzuQ+95AAZSEi6UoFVxb3hZEL5b/hYREsXIOuqP3SvI4ea4+6mIblnCYGnBCEY
zAPtrzq9b+OcPl7mJ7A/uN+frzFvSbLckKpzdkEWrfba88TjHcueIGZKuvygovkj
DYnW4uQbdHu3/k8eDLfTPNcZa+hqjRdJ3k1QcDECxGpHV+SGA3o6Nnq2jgIdpJar
TPKpj7AYoJpNuoOmVOJ+pE03ESHEME9gBhBHU0x9+BfX1cpjCvmaFa4/kNGYmTRI
PE0E83xPpFLug36SfAf40HbrbPYQ8Pqh88BqjL9/mrwEEfu079DWg57FsFSDJt1f
QVVdrh5U5prqoGYgBPpTcaLPS8bi0p69oaDz+YOJY0Zl7Z39cxFaec0vAMYuZGMY
u8wJX9buGeBDLckxvo/q20dDsyGmlW/gXJLqpP+gFrPBQiq5KqvdCa14umE4KBwc
A6B24PSMwe0cVZj4SbmlhLRTE7Gqvx4tDKgEKiEqhfeMYLXLzXlBTT6Bu1EB9T0y
TwrcvK3I5cDLfU2bGjXISxiCC43vG3j/hyCbk7ydwzR/stUq6rjufeg4mjvewTVZ
LMP6DA60067PgPKzwvO0axKaqq+QEPQovxO+avld/4SNRp/7jIqkKMm99F1rxbMt
PT/E9U9HEFuE4tU1m1zgGzQKVgYpBYYhxcKKF/hCk5fRbwv7J/YSYEvrvC8AzXoE
nt/BZBHDwzMNGWV+mDni1G/jwhMBLPFAJsKuLGDg8ROuiXtmcFjLA9Rcu4WUKkV3
Y5OlsNZUynV8gR4aHGjLdFKlQpgq1jS+N6Mb8gqNkZXIGs9Z25V3WtIVTxx8GL3c
aGQKD80sM8rlM5MxUAeCNeBRv0Nv9cymTmSSMEivcmhVILRYXzDfRc8Su5zNJm2W
UVYYX+VydlUKB2AAlG27Kkyi1G7qmNhefnmmEvHA3TuoQkF0A7s1WBS03gyX7cX5
v9Cy41EZtoBR61vdLUK02GLMCrixTJD1sYhioeWQZ0IvALD8WS4BLnIFuf8Koekw
96L6ohw1Hzht5XZicdmwmlUMUKDcpWeb5uSUaORLcfsmZ0ZmGBB20j5MX03fEgSk
6WzRMARwTbAiQybwAoxG01NzQb28GnWwGuN8BnimOHjfgflz3uO82nRGACJBl0Ys
r7Phkppd0j8mdymLCR9jQ6dx+oC8MiSQUqgnYb8nc1faHBPPCVlMRJGxNYVjcgod
ebKgr3DnuDccfXB96i5v8h8DdcjScUv12x0oONAawWD3zoJpfVM57I4iMZf4yFnS
Mrmx7TldpE86+/e3j9rtvRwdOMrpf0dwO0lWwWf4DJpeELF60yQ+8P4+5COyjGSx
+znWsm0jbC2mTumwKpexjifBV+wodHfHChDBpck2d2AHdK5+Jy37xNoeHpxOpR2Z
ImwQjzvqZXgxPQXmBhlnDm42tUsyLRTC1Tp7lGE6WLZYo87l6AYMbGefks9DnSud
r+EVutGsUMc1S7dcEou8paEtgaU/iRaioM/yGK/0qzrYbE8sJwqVyHkcGmdCk2eV
d0RMWB9AGJjToC4uNo66WJPdFA6Tt+JAfvBT0HUSowQ+kdcAVTJrmdUQfswJ1Exv
95GGXi7wLoAM64UuexDssIO83d9S/pWAnAVZe5xfqKHe3nlPieVY+Gf+2rp4pk5V
33Tqw7uFAaZ7VmWp79Ewp3ICs00vTWz/vNhluWp2VPVPDQSQMn/x8xaTOvLvyXjV
PB83WJgHGx/SQVm47qMzRZ6CmdQ48BCEK4bvVWis9WrGC1XdvgY7RLFVN9dCa2ZV
YcBBrFsvDSpA1eKtF6aBDFHSQ+dKtAV20BJvv1NEuvn4lWyqgqsIgIpZvL8sZQK4
KRUJnJ1UUty9b6SCgBPsFMi0Z71N8UsxCYuAdsz5GLzMMf/D30JMwxFDAt/9CRPC
bvB73ff7PC71M2+jrSHRmwkcAKhJJZx61vyThHXTUaZ74bEVcPyAlep7bg3VxZM8
RBxnueGgz7pZRt2Hh3L2jKEAvhm7SyxAc8f44sA2weEVcgkeq3X38NYpR5/yYFIL
c67WrU7ad77RoPcfM9sN6jjv8BKcF2uh5HGn8Qdl5LZLywYaTMIATb6ms1wrFJN2
ocBLQu8fjLOnBHZFvIFbdSdwBJwxyNVc2Mhxm92N5sDphRg5cBsqnr+IcvCccPs5
DLskA1U1WE1K8+zMrtXNK3/bfikiK2kkfRkk5Aa5DDKPQJBizGnLjCBYs6cLO4N2
qBlr/NibnkxtLW5zBMrQnidMybf60m6fmQBbk03+shsWmKEeZM3ET9JTjCptF91M
zc2c+eVP1mOp2DN8MXdcXm0UEJFXOKfLcfCQZz6ACHAYPRdzL9iIr6QLpRvkWuGd
lRLdvVKYM++2h1sir482SZQtwdHjrz3mDSAeCLQzxHN1ijOK1hUTTvc2f5heTLF5
cOGYWc2RziZfHmnxAn8IWO/BdXaA6nAOYYQxDb7dGIdsnACrcRM2okcz/hF0rc3X
eSdH/wwAYJaBgGn6ghuuD5vedemtwp0v/wKdBxCkvB1tGS2KRyOJiHhx+8/LSCRK
Ds54yUb0jPYUCwPlExkYKXiGW/hkRzkHuJq7jBH7hoqusuW1xnwRs9YyA0ddjY1n
tdS07TmXNu/M637ruglZESyb/aV/lZlSMk3Z72ZIZefpqR4+ZGxJ28YPjvQVyYxT
C9aKtbdw7YbQ0V1Dtxzsbgmc2IqIDlWa94z9H3qXVbpQUeOlHGT/PO2bie7efFCN
ttIbiWE1reeqjZpRCvP+MzzcswyKEZGSy08jJFiUe6Jbq3bT83Fx8jmUHcOdHKdg
ZWUW+NtoZKqO6E3h+ym7N2kIuDsyY2An4Xi122fcYa+NzAtMqKJg3qezodJTVBB0
xaWYW4Ug5SRntVCfGFyOAtG/rqf2tFd20GZvW8dtWOcwfWe0so+cuyt0ZB8xl07T
8Y7EpjMXgfxPfXG1GymrFzqYAsGko8ZMMbWgBqPT1FBBhtg+LtnxHkB2JsCb2MLT
RjdIjBdI6Wc0VWxnY1s8Z4vZg4v61IxZDtX8D3ox9IKcUyh39E/YcULgEoJlnNB9
B19WB7MENfe986G8JsHWnHq++AoJRQ+VJpvO3CeVK8fRiy9Z9+F5nSvw3DwizRe1
rvaVpqee55gMLETfBeSgJg3JnYhzZFeqRa/5BGkPLRoYfjOFzSr77VYCPCc/vJdn
b7pANvPtPWVEihlK5YReSa+7XBrSfC3K/LU9JOQUE2B1ah3wD9RUDRWKZ5x/qT5h
C7zYymVbFP54kMPOBDGhw1RbZTMYmd93sRXG5XQNtukYyNKNM6RMp5pYi21ATAg0
P5FIqrFGoA3q0KzqdzAQ2+xQGfTSuckELaLJi0FVgbu9J3mAB4ZXUgKSthPd9gMn
NZ8au8YGBYKpXBlh7BHMGeGZr/uki8CRb2SGq87fnCxOOMkB9WE0+cTrAQSQag7h
Z4yOfyR4l2Phk17y2YoP+7Gk/SqcE3tYa0vLT2zFlVviHgzIq3o4jep5UyywPATJ
8ZurJMRTYZ8lxMElo9OFwiVDNufnGt8rcVnctsXEG9NZlgInP4qS6/kbtochMeXR
pSVlrNrV0ChfyXOMLdtzq6qd/eS49witEdNTii+muICt1vU91zmhq9oZAUeOORaz
+MTnm+m3JnTal4SLW+QHh/e1qysSDJEJYeSmpiWHljOWATWAxC6YlUTGf1yDenJj
Zwqo116sScvdhosVgYZbABEq/ybWOpZoCOquQ5TDCVkatJuP6/jgoyYL88duPcj2
U0q1DzaTQEvfG3/aagbKSTGOvghXm1xOTr/lw8kBIkC7BP+J/DOALBOdCwv6WWQD
Q+7eyXQFGpMob6R21BjDcIx8LOdaAX+2BqexI/J/7Ag6KUaF895OeUXgnqJov51U
WvCMDPPqZhLSVi8Gt3agy73G5N3bnpC1SdueAu0TGAK7x2idda9vxha0R+IoTTF9
K/cYljzubF3X1lwshnjQHvD02aOYxHyozGKydbKEKfV9P1H1p68uQxkbat/oknxf
GUKJ9f4GIsfFfLRjr6JrnozVZXee5o/8SAGyHhtaqmLZbYGdWWHpFN/bcRkSNDlZ
/Uvs+n8jZt2c5I5TkuS3sMi+I9kaOtRlZhEWxdgZmaRXvGC9Xkkzk4ir5/eN3pEf
cIOIJwQs97k4nyJ38n3eUEq/2e9VoES7gZEN3TNiF/2RuiiFGH+rehiwTTkWvQR7
Y5KhJpUbkn3h1KQZUlMSncvZDTHm++yLZRXXrcTvdyFeKsQjEq9XXvCaDEFJHRuC
GvYqy20KgyR31vv79J1Rdwxbg1uGrm5YaHl080JXOg2U90z9duxHB8gMqgLtvx5Y
npGafY76bh2rsE2vw427vVhEMKsMtN1j0q/BKJeMyvtQHi1vcDxvYPgqPH9td73q
nUpT05RPNRUXQwqnUiBmlt1elIemcH0UB7quCgd0PMaI/pDeU1IZzj1F82AnhoSa
xss0Ge7ki/a6lsjNZHgL94yGdG+Xvzm4U5FyAKDENeWVOD2khnHexkMhxZwr0AqM
Q5C/s7S+lF0/NUggTCtKz7ojOo5zhlBwbKMY4fTyapatC0lQJBWK2G5jX6TGnvG9
cQMIQKm1PYF6+ZH/YgrzNplnF6FbbHOLciCodgWp9Sb5K/QoRAAo7+I6EsFhfWgg
97VJ/EhTyWIxJObkSIwBp8m743XIqp+J/t99MmsxycbVH2baxqcKJcTZ26j7daUy
ICrCVnDon5QWIHfKs+4P43Iveb9cW/u6SvEy9iUvgwXkyC0P4t7j25Q9kr2BpV20
7+/YredAjOxVylNNF51rffnjIeMQp2BiY5Bpl86wF+khOBoh6+Cuae3LJzW2iE7y
VSQHs+CAZSwQFTUcclXLka40Y1s/zDe8H+R4bnkSoIxjcK2CXCdGfsNFr6S7/Hex
9vRjZ2jJXS79s9bXiZhnwjn+t2QTj2LLenlOIyroOc77AbCy3tCcpJ8LQp+Dpk0H
K/5utpjPLxnQxEl5OZyizi0ZbvnIGbp9mJUa5KT6MYTy4R/JB3ITwt93Nk4HC84+
8CnbM4kRz3Zj9PRg8mGyTrHk5msebTkuK2DLF9pmFb58uNG+VHd1BMSXei54BlaN
ivannpIh6pSk7OD/Qv1w9HJTX5PG2nXWkmy+bA5da8e55SeF6SkjV4hGCt40E2IR
x80bmSIiwugxt4KfuG44+h2Rq4GNexXwoGoeba00nh7vE45yPCYFzq4bBpsiUD3s
NdDnxujWtbj7hgNSUW1I9ZKGys7RDiXPTnZdSsiPNL3wciO/5VpFAXnzDzpYWZJi
2u1kMtsaj4e0XeluGf8bx1f6xezxjbinPTa/9u5wRI/RqARkps9lsPO7nIoZr7pM
aYSgLHh6ZVh3934EMxYZAw6NQR3CCxvDfIHlfZjqmjF7dNmdsBD9cR4y+h7XDpZ5
U2lmJQTuL+IuuY39WpuzmcADChv/PN5Pu8/ebmBaDynDZTZJY2+gu661I3T771AF
4xmIKX2ZNNXMpGVN/PbpDDVGSjyNoddUP1BbwiBUlu+hcq1DZpdRMeo+cmM37LF/
H5XV5X7uUzyiP62AUKcH27iY1RQfr5Qpu/SYi90rRzvA7SRpugyoxOIefJF9UBzN
jdoMNAcYmyxHoettc3capVL1I6OI7kh/VzNMSJ/W5R5LklVsDgYf0pycAMh9urE/
mc4aFksqvQMYakbSGVSvIvMCWRq4YHomfPchGKb3jRgYNUDxZN1DOsKBFTKkWiJw
iO1FigVexWgir/nC5qpEqQzqlC5RQEg0MvpJB2q0EuZZZh3LNTbBjZa9Cumb3DDD
u65kMJ20o/yVWQATR//6i+Elq0vu4mDvi4xYxhkY+Z6kzGuWdQC56i3v2Xn1SEw3
t0hqqufG+o0jpPFHQNEvZfV18cw9cm1Dcr8xAeplMpylmE3cCGm9MGK/Z7pxle7N
RZdFLZKDQvzhbOkrrCgSPvp325OgXTVki17A0XV1gRExLTVD0zDTHe+kpLhtl42M
UeroPGj4BMh+E9pKFolK0iY7BZCChpJ4iOv5DnMK+RZc/PwXF3BSXtYYDq/Y5/z0
RiO5zYhcmyWjjjZE81s7oAizDGQKwgniZBO7t56T66QJxk3Fg/GQuDUbaMvAIIu/
bhjoR0Q7EosNTikTiY0Y+sIm5oeop7lCqMxMQsOTs9Pu9L84xWL/7lq1rDOw/6cM
d2J+C7sAk3koPxQfR0ezp3B/l2lrtitJV6pFzAKKShEtJGqLV6tgYxgZ5frTvbhI
go/S1h0JLdY92/I6tCwZf+VJh8Erd4pRkI6yRg4XAw9EoW7xzM7N/pNP7nTb9yn7
BZzmpToxgxOJ42B7uIX1ZrkkezUH4VamBkaAjpSfYtHzezmRMzA6eea5YQLJ5NU2
dbdhLvq5DMkOpdsUj+x/q732f6MFQAu2Jhl8cZjW9aFu6eo7kgH2pC6qVPzC9liU
mnliqZX7a04+HxQ2TidePPDQcU8E36x6L+vNnK59plLhgI7sjU70ORgEhOBF0h29
G/nRle67698G0ifsWDrDyFv8+oWdiL63B5t0fXHnNpPQht96oNmzyjEVnO5Zprwj
JwbpDNoj20DeEcdUJscTIqdB6V9YN+xLrGD6IfZQ4xawfINyVEUh757qcJ96Plgz
Nk9MORii/f6iyrZ/cxVqgNzqkOBYyanGR1EnoMjd79V9P5mhQPij+Pcu1jYL5uVW
2tLXCANbWL7afRSTecfrmoS2Lyq3SIZKXqrBMR8X3trgYb/dPXv3lRKLvCh7e9DQ
0j1YJagSOosIW+Loy6IvPaioFFVy0d9N+qG5e8rp9JCiz3BnXoCpomQf/gVB081j
NXPXeoGSrwDSHhBuHYz/vrC5xvDUHwc2L4yUUQ11Fz3pkIYhnye7byNCKGnwh15u
qjy0TkNknoLZUg/tkbHxh8YPQFpmpkUS8wJOAPTABC5dPrKkGt+bFfFAPaXeMCDj
jNvS2UEc2LuGYby8EwMAU/dAj87wk7wSwuOBb7tv62hBVJet23bzCYzpWecDnwkR
i2ZnESaso6cB2QGyuMWLSk2B1e1hqucAz5QBSARlHalaHopcvzk3eFd15ch2ZNUe
yedamNaDjDKAn2AMIoPVQuaKI2UbuyFcbSE1clhxZqA1OgJLZ135jndwfTfGJt8N
Z+F/61zSnB8IZ20tD/JCYtWlMfvovRbOd/Wm/2XY0+VeWmqffqFvhdEqTYmQy38z
kiNzB/y7FdKkV8F49uwKzWP56EbPoaof1xTFwawGPsVVa003cEgNTjImxGqqubfO
+ekp/gVDAJf8WJVoCb9iBK2TrRBkMyiOAeNqLIuA0FONOKGGAaVK3InTg5Q3GLEA
s6I4+VYLYlRuKozpmcnhib6aFTP/2A3fiL7SGW31N1xrBxsowh+zENjKQ7pho9mY
7GOyQ/8bx2ygoGm6BzTqe3Y4OpEG+yPB6TMf7mPFxvMxBKGxb6y61YJt44jhcxzT
Op7vc0Dd1BkNxYnNPJbJns3Ypy2cmN5nraIqGffWO46xpfTpOLDh99v4aJu6dyAg
dcNi1sVyP69n+mJJ2ZJZzM0lSsKx/a0aRzdpR6qgubp91KxDzrIx7LuK5747eLlI
G70XPIxOpqjLsPaepyZts2ncGsWGKVj78i7TPBgziSBl2+7Ot9FbPQriC3fmeHRB
RhjdJtW0jXHDmbC+WgHnUXOcvpr2+NDp2L4JdS8rXOoeSEqktoZtz20BjQxcT1ll
t5u1rIo0jyOCfSl07Omn0mN3FauRjM6//mwBa9I5sttxRhOPlKLCy38by6g2NPsB
NcCN3wTyae7JKUS8nq33fsxXAslf4rb3qayLD4UCVyNF8TqM9ht5gvPgbN13KHQg
3+Iqf/myJFT1IUi8RTWlUeauQ7of9DSyNvOEJbnqhYNpD1QiLcbwULJ1hXoe59SK
hiaxPSsqR06HyGGauj1dmPJmuLYpfj1rneq3J7GJka9RRNwm5fFRKqXfC+PJHy0c
QSdaewWw4GD+MWqkPGa/D0OoGe0wN5k5RLaZRg7vzaxiAvOvOnjNe7PqYjq/6G5t
k/z7A5RyA7BgWRh++9x7TPy7aznnEjykscOG3i+XSV7yg9hK9CqkJFhnRs5/x/7f
+mHppBfM8x9bMk1/KDGWy/EUM1Ea0Vo8m3HC/DK3V4yrbX7AzyvLlopgSpOimcnn
xPDCF5d+BLv26Bm+18Cpdd15+o9JlNI0LGdGPHzOGEnspAE1B3/HveMO6LQHl1Lb
aK622iXixD8e8AXYXJBNEnW/5OJvXSzLzeHw5xirDWc25zJ/FM47+AezfV/1GMo1
RsdQMgvkfan3c6l8BG2+gopD4APNI18Th8nt/vmpZ29rQUR6JWf/KJkxnzX/T4tR
jSz0EVXQi0buwFxRkVDggICBcyL5AzLf4hK95V7vW+7nItXBytqrxEJGaP2iPFci
qStq2wTzXmSkK2I2Zc9Z7btMC+hochzTpbgr9RwwOqI22jvRtbW0bPCbEkVYx2Py
oGPinKFG27dhyiEI5UeQv6p3uXGf7WQr6MXjci3JMTdH3sfELivaSOSKFlOYWJG6
XVUEaSD/hAUsGq0ZAHXbVji+6y5lk2nivWxwejwhvViBU7GEghJ9rlVPnsj5nCMG
q5lzqyA6ApCZ/1l0CoPr/Gx7fIqbJsMoCtBAxUixjoicluAWq1G1kh5KfgDdxnHU
8RlpWV6dyHloai5hNqIgMMWzqWPsHBXeS/b/YCW5bFp219IuKMiHmLS3jesfang9
mL44ZCDra5AMuzCdcmegmiNJOVqzcZB+jlg86v8Fq3+NVSzzfvpDk+mcF7neglvt
JrVKLqeJ9Y1ZO7t0VmCtaS3AffQVC7lAApaG6UaZqynhHrCsUKkD/lKjoqaZdzKJ
LhRjqj187fyQzsUkiX+6MCjuYR2GI+Kxx9+iLrWVO0Ub88Xj+mQfUULBGRMsofcB
I3SYltI0UHzpvJoehN0N5qvheukXwnHYJexQPmpZ0q08rwRjJBhoujNAmBgr25PY
iKo4b+wmr6natW1MX/5hY2opMQLU654hEmJQd+MJDKuVWY75iVVsz7V/n8AfQENZ
FYXobeph24apaob2yJlDA0K8JyTI9g1QAmXvKjrYyFLDdLRUYSYggiHS/iSgeB05
rIv+4mihfrGYYbYYbUgFZufTaS1gir5BHBRNlJNUeluKOq6RsCn/wbkbvaiuxLRW
e/pQYYn7GRa30ZcZDXN+4k/Fm1jidw3iIKE5z5LMBnLieJdGhvGbQSP18bwA81wO
raV4hwb8EilNduy36orFNVa5LhmhhDK2QmGCQlOlnui7EllgyI0uNPJ7ugqwv0q4
9sE4QZdmqYMe2EbIIzEhwX2aMjpgeXtm1ix951A8PKcfhI6meENy+7zMeDVMsOCJ
hsaKnyPm+SQViKPwCgrgrx3BrQNZucvwEAraMmk3PewZHwWrlHVFG2Ko7gVttQjA
RS4qNVLV3o9rYuSvCurLReFMw2hMno4JcMAPy3RkHtb8AAhJOaBrwK8xsSO4w4h4
Q+QxUYNtLetn05EApRw8nNOpmZt38T+8seCzD67GFWePa8koBdi7gV0OHrh9abEa
GAcxrY8d3+/WIJRG1+0J6YLqw/9rkpCOG3667FV2n3VrNxnVkj1T9+a6WrpeixPn
LxbGU/0sx4xxyin3djvr0m1m8zuIuXmU8UXV9DF2cPVsCkR9hBEr0/gfb878+Z3x
cRnGcAMcpFgSXx/KXuV8Jei7vuc4cSmTRbOvLth5EC4t55DxR3QPZe+p/s+O530o
pw3+jnqyg0ZE5GsPHx/XTiTqZmBhbgm/ax6HQs+WXUksDWf56fuaou8Nu3rgteO9
Hzy06d2KgUWUpgbPoh8X8zwB//rnKqGdncQX/4+l370n8yqsJPvbDDuZlR8Vvq6+
p3pLlcB3pwefHeGU8y07ZWvPOmdpOI82Kb5yR1j4H/yHrlUkESV0Ct036BSdg4m3
wz1duZlfyzyrIokcR8qw3oDke5+YbK5k7v0S2gc4CyWZwgrIPLr2P4aaDlOw4tbP
LkBDQpv7CoYvpA0fWp+ERk1qExWDhWH3P5+XwUX+ALjjaasgzG1kaO6dyYKHR7HB
zZSC1K6+W7Y/10IVXrR2oVS5g7euCfWrib+XZeer1ZOaT+O1ZsYXE4LY8C7mhWzb
KCnnQhLyBcI/5HF89dmTSxSlLaPQbldgeaOiC6gCYZVwYQai7phlYKJ3k7Nij8bp
BUseCtCdTZgT6dg982G+y7LCa7TP7Z/gtp6oP9uN+c9F2FkxSODLCUov6xhHR7Dy
IXv4ihG6F0ZF8fTdx/qkPQf0LwO9PhrujHhnKlhmUGv3i3PQ62ft6BYpvrPv5z4K
JmxOlnnUSeLGXcD7QuyNsiGxuPr/BCZm/nuY0B92pDi+x+32Xz1dXcUh4voskr//
9Y7GhyNA9G4HMoyQCNRVQr+KScwbGYVia1FeYiBapvGtU6dybTn7dKOGZmFpWIHp
pU5/7D7W9yhnUaKr+3RN8bK1yEWhJ09cW35DuzMEXCmdaDwhkQ9co1mUzatJejnB
KMhHTk/BiYsqEN25WuRub72skv0G6/w31QmyXJ2D2ekej8DTD6/8Un+5qMwg31hh
0HXlhBNfqjN0AX3o3yKlsUCGAT8fEkoWKIYdAtyU20fRou1bg/wLWoW+r2Mb9gyX
N7Va3rn98I6DyJ8XguGR4x86dCIW8ciKjvdXCw6Y0mEaMzoohGWs9g+nJTaLMlBW
ARwxn+wK1xxXwzYHY8WYUsg1mSEnVHM/UhPdY5cfQ4pYoU4u3U5wAaWKCC3t4LQ+
WJyWIQn24sZCJugvtCi77NajURxrMV5/blYYWdmpvIqJJjIfr/CBDLPBwks/FwDy
AFzUdRlVoCb41RbacTup6Nx2kO+UGAG8pjgQpDMXFSoeei9hjYVOnltXBdIdUvoP
4sBLGCOkNlX9kPmKeqMMgHfTf9bU/k+TsOaMTqb2VRaGaEOr/JveC1MQ0XRji+6B
gudp2nBpzvVb7Kw78IGtRgQKwq2I5k4QMZdjD9UlVipOYy57q5FHzBoNIHOwmGYx
32pXysxP/6fHTysDHqZdlVXYw2SaZZeEsG08GdxLjJGs1irsY3hDztnBI6Kpu/ub
9NcGhHEQE47xvFTHJ1EXKi/8lNSKyH1MaER5BYKJJQuJrdkv0/PnLMs4z438XEy6
MaUb2noVvQZDKF1S4l3vv4xogpL/Z/LmfkCeuXO+Q52DVtnh5DSXHYIyHk3dEgxQ
Wp/++rsDhdIfvBV/9DOcw6O4qpJfIrBJCjYymvfjfAQloPFpSF01TNg5Kyovd/Dh
u9GsjePmnjHHvZC5LECAIRGx4RmdAdW1lC/NGsBUtB8BOPVghhocHvf0YMjWL5X7
X7xg7dsOnrQnhCNJJ3c1LFcU5MizkjaJJJWLhs1OkKgQ7ur4eBz7cNFiG7TtRqSu
RtKyBtVkGEnUXYL/pfCC8LVJpLMObOM4OxVGX+6E9KbxF3SyT+E4ZfadNJ3qwljY
tUcX6VJgQHoYFKStyrmoIcqUC+zKHdK6Y1wVljrw4GufBaK+7yRTTE4WZyzvBTHO
YSSuMk/RsPJlNRftBGSUgI3jLYLEcry94NBSZglKxvf4NmecLECah+MhietwCuX2
9tJgL0I75SC8kHRB/J+jxRgCycuPOSYTmqFOM6LLgubuJM9AJA4sb3Bd5qW2le2G
H+6lsyoc3dOOcKdIbY8BCOguwqUAKACG7PA3t3yIVj1xZv6t74c8oKMOnpPvcEQt
Ifevx9QUylHW2XXMjFk10tCVQIMiovFn/GLN7wL+aQELBxjNW4aq8Q/U1pCaH2Bg
ppcDtJrihByHOZuticVVuJfekd9lfhZY7nNBtMBWWaR5RI6ZtWVoE3529JCy/eha
wx33dc3IdY1posBovNV5TkFBYIf6eykurUoWSbsXdqU3WlfyzQLP136TTFovLr6G
DmTxswx0vbnmWzUWEfaqjVhtkIGU/fIKVkWCn6zpD6eZy4zbaFJ2sQo/zIanjwSq
99YeiUxrKhkP3Vm20xgHty7e6FRwdIfNastTl9dRKRe+7mjlW7cbKCYnZhf71xCH
CQ13Ww6cQiO1UIbfGYvlqxTVGt29awKB3Eq5XAjhqfIoadYve/9l5aOJL80mUg++
4h+bqO7x/gTefW3QuFYNw0eAenqpNvfWNLLOcnpVzivwaTsy6yySPLIjUlVXg5sX
9GuI/WZQaGIHZBBZE3k5FD9v657r4WMOtms3jovYml40lsG6Ity9Ikj9lJNTuKzF
X0cBZHg5h2E7X1aSdby8WdFEO7XqQijbNfTmxPBgviVoG13TbMrRLXtcmBpmJN//
tJaajfKvs/SegYXj+rGn9Y+zJ7TOynGNU4Vc/cRokWnH4TUsFLhO3snaepMmcG2J
m6Xdyh60sTl/Yybr6bK+raXzDBJoHZn4ohQ1GunLExB5dLe4ffXYNFu0L3TAtKZ6
dxB79WXQmvJz6yE+9bHHYTInNLq5o1VShsNI/0GiJU0WbBAThU/ceuE6ERkA32V1
c0vV3P8BSdM7WtWlCEqImQjGb1hCJqZ2BXRNQkebgYZ1qNNbMwpPk/5mdrpxXkgk
K17/tsotcjz3BpGbjqWwAnWGsXsoHyaGapfse4uE57LuiXxO0+2qZ6c28A4VexrI
aguNDcYvJkOnsB1HrvedyXmHOmVx5T9euArsMiY4Qc9b25KxacK8vI3WaQOmBHlQ
18YHTH8pC+gKZ3XbzIzukhjs7cVFreIgj8u9necY8xcALHS9kC8F++xuaCu46CA8
cin/UOFW4lVg0sD42I5CoWWXvMLExPuD7fh0BuXchvkSv92fWnYD3yKsVwLUC5dj
3HVNwXd55mVlx7NuAnJ9kvn9lkkxvHNqlw7+LrOqM3f84to+p2VCbc2bcq7PdAIG
8ZrE5QUnQjSXqZkjudqFSwibtaJBhJBpHbzLZzJSZHPeuALCPANm2gBy9EuXvUI6
AFp50o90qFi0N8SHxWCHqPv4SnRvKVlHqEoaAMSqkmQCcZfbwRPBVK8YipCLR3oJ
DaN4ng8lYemgNMamppquJM73AZzU3P64ILzwbT1TJmJskRpem4NTw19pVOJdSVz5
+yKaSa00VPdgrIouTKKC/S9yWZocEwNzgiVVW40TUmaW3FkgkvyJrvl7vImOPfbi
EhiPGPpdTnNaBs5Mm/3aRym2ScYQo9JZtFPE1DciGC6/ERJXykOdlOpnEAe1E0UR
DZadshdTF5rNzQPrWE+VunBb4x15+UrwCrXuEAL66UyCeznuFkjgMOfNI6cJwZr8
W0MizQGgco4Zs08v51cI2Ei8Mg/X6p4R8OFY3bcOjwQ=
`protect END_PROTECTED