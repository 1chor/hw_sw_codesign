-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
bcZ30W6Gj7ZhsDzYY5X5W0U+ksFi6GObwSWTuLyxUKgGDIS04QkeMgzzWLPfM4YU
5pZ/354+A2MNvkoi/IQ+arf0di7qm5v3Je9u9qdxTHdSvFKYsxcJBAxdBedIveB3
6B2MiShVxWfzF9H7BLlxPtkSsMWWzxoo1rScr+qFpraoJjjs/2fn3w==
--pragma protect end_key_block
--pragma protect digest_block
iFdFkefPDD05Q3N1IbcLScvITLc=
--pragma protect end_digest_block
--pragma protect data_block
sviH0IJCsvVl2h+0g8OE1yhcmOHoT1wKeFuuHSd77++HdaPPjVB2qCbJFb177uRY
+pi55oMznBFJFeJZg5LJaSIHUw52E75bunThOQvlrPHoDaYzRd7R2qGmFduX14D2
V/hOH6EoFTn+LdZG9v+KeeJEuWsyjdGpMSg+B32LdIitNJlI1ebfnxDaWL7GLl5K
dCOM4dYx5pCDc7/Iz2yHQ68+oLdbs6moqk5TxttnRBzhqLwbOo1pmKpX+HNcA1Aw
VFG8bIsv54LJGyXcLguRoZumpIy3C9sbHQlSGKWRcXOg2pwKFHSWy9p/XGcgJlz9
H4oL896rxBqNj2rp/fUdL3aBjbMDDOphjE7jmShUAJS4Fi5dGg7DaAqz331JtvMm
ZViEQY+wJRHVCzRFhQDoZYev6qU5wa3wVt8fe1r/bzYznWk5r7n1kksV8zNlhq2z
VO9A6ZYdB9hlJWWJICen0w4US3Ji0ay8tmxY4xMZYwGidIR9qbHpWhz+c30TMmla
So+M+eOdGT9Z6TCIg1EURwUWxRvhy4Zc8GQtjGKE2dqlJgO19yLfKGItILpyHbml
j+sZGRNLcl8kFwvnGeqB/AUk37OuFKGipHMMojXVQT3xCa09x8NWGk3uWsyzPxfE
Ng9fRaU9S8FVy5rh8e+cEHZUiJDmj3NmRg0EcUuAAvSKX/pz0kSy8w6ThyHP2oy0
uph1D7r9SVQ0CkRIVfL+H44fPPg+EEAnum6CnhTUXfCixiFmBdo0pfEvuFZvdDdo
FKTkcXKgeo38G/QjKYbcut9Wx8Y+v8rWTIPOBZbqTZVePmZzf5gMjxv8sqQVOyTm
SBuJvGzJXlav2o5OIKaB0wg+sRBaZagOzuySVIW3voi/dOV52EFA/XyELmxJqqrI
KRWPObJps2bjvh2wXeYMjZoPBTi/tTV17Cj0WTQk4+VYtYj0kzXN6bCwIbpuTDcB
uMLk73H6ja6pE7JRvgbFrEXDfr50dPw1Uy4odJvlivH3D4/smFPs4sKa2AjqukNh
IecRuEOGGWHEhsqAv5XBS1hPHmOQ50nuveaOoayLpkwcij9N2PfDbVJG5kmSuHEB
SGncMcgi9vi1JSFN3LUEZCjuv9sEPgiJExoSavi2qNGaLgyPydMZl7XuWlSNWgAJ
RL3pyJ5kk+UP24Xf7f2uqib5bo2s9Dw/ELtQveu9Lk8FYcFEcpnu9ZskED8SB3fB
h36SaJyNhKn9G6SJi+p90F6JVmGeZx/Zs53jgY0bsR7/gfTQW40qJ0PKogWh+Hti
zUzIsre7fdTZ2750gZM/0U38UU4M//saOzkb6f+fUAT69tV34R3ggAg59Fgr0v/z
Cxd0vyiE6tnixv2fpqcgKWZP+MK2uL/VbjfJEe4DkMChv/yeuXzX7nzu6HyIrQab
yYPPpeEHJhrkcoApiZ+lt0NsgRHfTLhzPP650BjJutNUAqBlcjce+e8u81KKbPuo
P3YIoG7NXgqBxLavclyNwevJgt859YWc3aSZeyjNZWUvkqzff/F7nvGol5Luy/48
ajz9ou1eT7sWhFWeOgM2YN9bx9MBQxFUQUanR3F34upipyUWdJUNS7tDpA7D2+CK
Q3meHPtFeSP8Rw+cb2ccWMelVKsOSeCp37pGEmDfq5TAn4FWyvUVBJ7N8bB7KzfB
cjcFvAJKihhsUwbwJDgSQ55RO8PVwSFC9OB4qRSj+j8a2U8fxq+gMz6m0bhx5Zg6
bN7Obb5AIPt8JcD4ijGS+MTmqkAj7Mo8RlYV3QIwK2n/3oBElBj+YjoVx7UJYqel
4JFE/Tu+ZEr78vGumvr9rnLtSK6VPQD/SRVvpJosKjgOwk/GR8oPhr+YZsHI8Pbw
mXQtrWS0JdAOAR1sA9aV4lvgNgPj7NV77YKAaLTgv668mmOO5Ajbw0do91nc+Rie
Aj2IoSJ4pl9+yQtwpeJGgAz2aunvk/wtnFSsb/29FcaRxKL6NrmWZxzNDjiqm8LO
3ZxunQBwJzWq4tL1L4QH8Gh4dXsI7R8aHs3YPE9qCv3xhGg/R/dsmXO6Ksyfpyfd
YedGhwDdZUTuRzmXRmolq6EDJRWiWNbsXk3j+frkPGa+ErFA7UBfnqgomABsD+9M
d65pgERD/KeM+DtgFfAIxuQWlQ+bcT4oYXb7SdOHLEtkpC77z6RxKqiQFMyrbzR3
YfM/8eBbs4TlLtISGglqmNx2EH0bDGuODRPKx9VHnlRWyT7gcF8ZKzD/lMHjySsF
J9QhiuA9QP2M40S3CR6xcpNbgAVOt9Xr5ZivCI6wZdrWqotGFU3Ivv2zHZ/K8HLd
IHuEAzOpYOvzeFpWE2SMPK6sAsI8slOZ9ldQlEw/+sm0JL1/cvJq1EdvqbJI6JwU
HOPViEWymUHt0JnmzJGHa+NPHunQGvSnAqDBskno0zNHUYiE2/pfqVNxT4GVs32A
sfF4t/0JIm8WYXZg3xLZ/4iMlpU7TaPX92dj+Mx0JcpZ+A45s84ZJvsshoDb7n+Y
8A10i6l6cwco4ZyX1FAgN2I33JRPxFCAlj1t4zVcFqxkC3dF/PNBPB987NmARQBN
BNwHt8hbtjcZpDfixxhf0rE06il+bRqb/B4igGuxMXYCBbiu7J15QA06rXBPUaPE
ibtJVOplyMewDXhNs6M9f3ZsY1p4hXIYruHIoFrVlhs8cw/Pb6mWYsf/DUCENvS6
jnfUP+/aDry3d7b/9zo/6sBFRjBi6nvZzFlJDAbCJaoTxXii7BvEJMpMAUt94RJK
hH9uc1aQp3H6jU42dDQulMwAgL53nFbSbXz//J4Mq7x67FdnUqBqz0K1bYKhoHJN
b0EKtYTZaCqIOwsrImUiBhBFA/7Y+pBu3qsyjJFSGpDcvjfZL7d8sHOCsyLHO4wA
DVOH5Z1BiDA67HHqKQHN4sgo/mBLmXWUKmk/FA+SrfwU+RwsGxjuX2EoDcnby7tH
yRMfrdGZSRtJMjp9CSL0oQYR08PWoMO9gPGXoVo/hFK0Cwq/ATCphl2A/uQc4Z1Y
v6hhE42oF43NC7nyEB8FmX2BT9dAhfosEW+kqPzjSxdr+6JaDEREMGtJ5UT8dQiz
W3qaZO9XUFa35vMWn6HsEQs0a1yB94vETco0LPSiMqoNsS1LvVnsRpKAWG1QuT4k
CFPlyFtD6jQgaEn10RONXdRg3gTONVM1BjRR+WxdvlxEMAh+Jsj5ixNn+G49d7WA
//883T9Pz/Ff8KL8YUwwZIax0rASW/clScWJKcqVxRhb2FCiBv/fEAgy8mBTxlC3
U0tD1DiFC/PhBvsTVDRqGaBiicIQ4wuCnUmJ/Cf6QTW5M6jyv0eYsn9fVDSKBNTi
vU9SQOfBbKRHJchSouTk7gk39AC335Gmj770eusT6O9lZqRhNMN6sONrujIyet4Q
Uhtv0J/Pz8QmjSvxRYRLlLuNpnawANf4+4hqlG5nLmat2yhxCrud+dvqWkPtRXzT
Z0sYqDqBfvCY+HYei6k0byCK5+G6tkhJAImbVBlJs8stIKoOqJ5xChtH0mML+NcX
0p5A5RxersPKBi1adplBdZxGD4YbDvlGh/s7j1P+z5LTZYX+eHfrWklHt85MN7Rq
Y9Lfa+C5pPo/MOFSBUhpfTeutB0z79lV/6BBPkqkkRJtW0kiGDXNBniQ8n2W5WhK
8kcl++/6kFeKMgHE0hNfHm2u+CGs+KcC3yOlLOx1TqImSOqUTGIY9Okjvf3+e0rl
f2W0beEnmn4D7WId98j9oxEHKxqxke+d/Xu8PIyHQTOm9o2G7eEcY6JZiyMWOUrr
yKZZsuZSzW83mAv25EzFuWTjIoqVrk7fL6OyO8FsQhZ5Mz42tq+9LnLFDsVd19Oq
8aBAEaB0kVZTZkCEIElKU+zOTx64AAPrl2kLXtILkeMyXhrlNGY9Nkc9ZgbeVGWM
ewNPMrzuh50ADnsaFGG2GzTnGbym4fxyucqPcrjPIVkIV8NArX0tqvs8/cJdkZNS
3QbmbNHYcRrQf6Oej4zyV6M6OGp/Z7HwgqOuXJgjQyk+rQN43nYpBe4FF8CHtSlK
EPt70xMcI1uKpf7OFF11ovL0cAxSUpvPJH5V+4pWV+mmnkCD6JWyxehZFMyq/jTu
D89ymMJEQlq2WsaW9lt/jG5N22TUC2lesqLwqsESHZSwUcvmDSvY5XTljIMcaVdH
VnP6mDqN2HgUHNueAdn7MD57qERAjythT16ebYbDAxKhq8hdVH+QRfSHsC5G4wDm
i+kRqnSg/XCWLywyE+IUCDPvXNOCKcjJBh8Szz5hVV+/Q5dgxNUfbmjQgyZxzNwn
5e8Y7jHtY6ftYKtnq3znHOFEnq23pmChDwpmV/TmW5Peuh1+NcYwyRPeQ36nAK/H
jRNsf58zyqVW1rqsgVf/q70gP6GK34Fzbz9bf8MSIW3bbZ4+HDtFGG44F1N1WFFl
/MTLOrGn2ZiFPxK3kfL9+AKNlUu2XmXFKUyTW7YcyuikELtt/Lq631m0RfKABD7Q
9Y77nZO8dCaKQLSgYRJ8D/n13K23LFA1nrUHqqW5k6fUQD2f0SjNNJvsNUEvwOJ1
gbVSyYvU69OU/5taR+qIR0rnCYkD4LR0f6+wY7v5kR2o+EWvsghghO+6kYXDHLkK
9u0PcohZLyYyCyDfCNAlcSMPwLfFKozm6W3Q2QMuC0LUBTBuFBhmBgBBzD/Lvv3Y
wsyrRKYgvyim8wYXjIUWtX6AkT55teXx85vdzowOczBLA4lmtBwH5LuGnPSXh2h2
ni4W/NEctlL6R3E1p0GQn0NZ0rPEcOtdzBEFgm/fenTEr0fJc3885V1y7bBrqK58
Hs1w3rkFYwhSVNpACUpd13a97UoaNVJ1FCrckcK+qAXxcy+uTFdp0Q+vcifbZINy
6jMJ0+RqS2nzh9vPAaYajQ8uJu8jMCceW8k4MHTRVmhW7ib1DNgbyrJYWE5dZ1nJ
5O13gscuwmDTgIYQqcYc13m/K7n0yq6MsZlEqgwpz0/C+zNx7+ZyJZZrKwwq/7pU
yqeqtve2/UkN1pFHcxVgFEAcDWCe7Uqr67337wEdv4K+JiYv8SL/IkvUVNgcsLPR
rcuVjYm6uplJHEECPxpbzIP3W2BXW2AC3C4D1NW6mN9DmXPSA62NsnkOPmuUPP1W
lP8xkIrGEntkvdjTtmBwo0N1XYE4DPRaoiHYrkoUYuD9A9TniH6zKJ5dmdjG+BrL
pQa3yGtwUZfPXJBVWkNf+4BZf9BAbTCEuZ1yLyloOsgZRbDdbN7rWuygpNNZr9p2
1mWda9GyFp5rie49pJMC0pSzLYEeCw44IffwuZZvZhL91LsrqxRNa/liKugdDYZz
3AvVld2+Mx1ZCMAoxZ4h0tPxUttVsySCcEdtsmq1xpILhGLiqHb/je1a8psiLi1J
qYigSKvofhAe5uWIwxC2LOfM2meInjzlUP8S74uj9wg0PDehSQVlRcSWpK+PRgFP
PPJoLVU/ArU9McWtxwPS4YdXeeMCI4/aE6F0JBC0T989tCGiw3oILItilQwZhBGF
BLtQh4xG0+/U7uKAKJ+hKY+iZ6kwSvvD4mt9lNbOUS/mfXjthETbo3WMN2dc8bol
biQy8Rr556QoQT3+Qsi0T7UzTjoZFOWxWku0UAhB4hQTONgo6OvmN8etTgYPkbXm
biXKrwWsvj4pr28pvsbvIx+Ael2reK0lWeWXhl9G/uKSxSW7tE7mF0bCrT1XnTyK
4M7otUyIv1RemhFSawqKA/olsxrQGTqYPik2OgB4eQkfH6k8Pm4NLQakLXkwgFsT
+ukGAip8GRLxykLh0F1Ks5J95tbrPd6uhxylof6c4CslrXPvgtOPS4eb3yGNgkUa
yMRjZ+OVlkgSl8WQnCgZoAeG+yc6scp47KDZp3zXHm/1HZQjGNfi7XAOtIKq6Rhd
qhoRgMcl8YQt5fsyd49MLWqGGSzlSRF3REmbcA4+aWEgH9rx4HR9N2cvKob+q2ZV
m/Megi+XIeR4Ha9wxqt0AYmnn1HbTH3czi3HlTyagH71C71DfMhXXwav/3yGtPIK
8M3Q1lnJfJfPaB/5h0h7yJxe569qASbopVdm6D0LFgndAfSe+2MeGx51YK5Usz9F
yg5SzSm9BvHFjU5UCEPRN3C5EYInWw0T4r9sbUhNuiqqbJLDocfshhhzXVQELfdR
8JCAxeIbEyca3738aSzvP2QgUSFHE3ZX5VXRjyZW3W12H6/sGKC/xgHqGbwlq6Pc
7d6RGghVkeFW7dz+MUa4K27dQPVHlkDx0Vj4ezKg256wjy5aMTAo5Fyn/NXSENOw
s9ug6zy4GmL7YDnDmwtWmfjO9W1VuEMv0cT7lLMmGnxWH+a711F9Fue4hheSTOAT
R89hmjDmId0EwfYnfwtbuDLjtmlxJXBbW+UQPflO44Vow0K5lpdQTWs/lFCiQIfS
v89XSk5M2nYvfOiuNjZuCn/JqSmWjIgeNFxWc23i8npFl1gohZDaE55M4pA3Ewyn
4CSOA1c5WnH5SiB2/TCF+IUpFCx+yCyME23cnePVXUubLMpuMI3lJa5jf9Mn7bwX
+QQK/uvNqwYUJVuSA8UOOPEvjjqb9tr5yjMUCrByMouRsLoaUsohmechnFE8avSB
5QZUJ+WHwSKOFlAzybEkXQnh/DM+osRKMr+jhoRAgLWBG6aRgDrBbAzupVLc9tOV
VfrjlEbVzlxaeNyEJ+P3DjRMjn93RfS2psY/gRSRomCxuPJyv5YE1/qWuy5vXdBK
igFxMj863RTafp7wru2cP0QFcs7byeAMvJ0IiPamOzLL2rWnnHXuc42e6F2iCQd/
tmYJV08r+pq3bA7igH9Dl8++a2XXumnk85kwAb6H5DRnoLg26q7d/KwtgTnkaJ6C
NYGrRrhZ+YF5idufc4qeWJ6ErOquB1UOqY5Hobzux7UtHz5yQHarWQYYaehHLqGI
xNdIMrE7yVBleDpZ+hEPbeZusK0CFFaF/wCBUAeUjbFjQLrg0YR63c00NaEh97qX
nSPd77e4TjYfLKJQ4CbRzSuMDcOLKHsVAlcLFGiTg0lHZwAoVvGww1Nx8VecSk/k
MGKiQ6l6QqiyuOoxAiYq+qSKgLIPH0zYAW+Wi6fBz85IS5w22gYofFkYwL1LR+ZL
aoCVxWVEoas/kPxQvmGFS5bVHFYI/taQmB3apAh0qNA0PcZt6xyooWHd+niIUvrD
ZmmzrWNBvd6UPd292SKUIPcJqbtxhPnkQ1TtZ8XIuHQCln/RGVD/rgTnuZ0ncnBn
rcRpDsF98TX2n2uR9mqoYqsfVn6EKWqI8lPKd4u06/7mfa4B95/yXwzNoS2HRBL8
l+Bmwlnn4n8nZ4Q0jAaltD+uvsDyma5CEC0Xz3dPxPxBsNqqpLShbzdmFXc56iSx
MzCaGV2kFhDUhwLbe2eA/DVsQIHBFC7GKbKsfDP4H90CKe28aiMuP6oId0k67MAn
JG66eAeKvOOfaVFhdMoU+3YPLiOqbOM/A5gIJNXz4nTAEtBMSgJgPrU6ZLgWNEwp
/6gG+N8rPHl+LdSMdDGSRd4ECkGY3u2WX2VdbdruQ8X5QqpnO3ghpNMtDqETz0YG
/7yj8BO5fNHL5sKRxoAKuelUHgiQN7WzvLO6G7Vec0axgjrqUTGP7S3hKvmLQmu7
8wKikoVe7iOD3kritJJ9moVc6D6nfYD/lrexGvkHr/w252OxKNlDWn8ZxFYn02q/
Sx9y0l2c/jVY+Y2ZDrtTQdWBlx8rhwQAdaN9DwZ7239rWtROeaEyrpvcBVC3kfsa
qoDf8EYaJqIS67xL2/ZLPTeBRlKceV8fxin8cXceh9b8FMRXdygGtJPnRGjiIHW5
+Up/4jDmCfa2YL+TI7v2IT89Bfn+kXZrE2yM6ssUd7NthLQOWy8yupQ9BxvlYKqX
Kw03V5v4uRyjFPrzr1RPx0TdGEwNfEKHZw2NBzqBZfd/c+m0PpjDRyYkEqXr5P1H
uIfQqbwfWSYdvm3E6kLVt6c20XHgiQ8SNIEzfh69BPwxsZ7kPxzOUR5i4BO/mP+B
JnWGicotmYhBvTU+PNrBVj8LCbUpPrvtSyTRBcc/Xgyb8kgt/e5/atbji1Vlvpqu
3+S116pkb0G5sTPo6EDdbi3TKt+QfeL3R4JLZjaz005gEGxZs7fUxraauBQNm/Wj
duXjRhbneeatp9Ea0EiDMkAVXmkZQLZSz3sd4mejHBfKXqOrLMaBw0AP5hYlYIRx
PHgQBXfZoLk78pZuwWPpo4Ok/SVVFuddEEs+vuEQKfMJIYceJuKhffB9gAPMQB0D
jG5u5DDs5gHSy9xxuYKv0zc2d1i4oikg3OFCwQ/KyeSqvXVz2NK7uKq1zeD9yCOz
RcNtg/W0x7YERM9jJtrYWn3sLL14dudEs4T4h9SIPp4l9rGPCnPc3MeiU1ewJ7XT
YJRYYMTH3Us8m1VrLU7ujxAmEtWSkdfCYqU2WfUzSnCY86X9hle/6SD0EqEh5Y+F
4XLJT+u8DA6p6ijw1ekBxnHeuXW5KpqYxLi+K2pdiSejTerCGWCcPNS3HU7hyDth
aTW1MYr9KUqpy4dfZbq4pnRJWBzwd+UQATLceofuK+KN0Bk6k2qCExfwDwzbzW0w
SgP5vBxIGfdTtW7TNDKMLKdESy/YGv4N8PgqtJ8BE8gD4qGAISuq1ifRC3pn9CJa
m/WaKR/3iRv04nLa9kjJ07VLEXSzJvO6xfE+etpVTuJKonnmXqTcmIBtA6wibOz1
w3i/R3YQE/boH6S0fXzgTRhwXw1CxJ9S3Jmh8Q8oW11/R/eYfNVhc3kReewtEWgA
JX6EgLvsV2cLElMnEgZ+dm5E/1hE80AvRk8aCpK1s/rp2lz1H+Z1OI+Bhb7FlHHl
l2g4gaddOvfBqOFer/sULxldJUM1AMiWSrPGnsDzyFpUWpqGxC7WatH0xrshOZJD
KMAI/ucCSj0blN+rT33eazl3VHnch0PRJgWD8sxjQ84+IhzCpRGG30RdqDGgIC8C
eGVIxcRF3Drurr4FsqAYfiSqvJRn7VAWM6/YN4Jd8HL+4cDyYPxB+tix5CZLmYWy
zPHBCx0hGOFdyre9x/A21nU6uYxW4Ov55p1OKWGfAqZt4BLx9u1CIm9ocTgmM7Uc
9MGdZN+S+i1JuDhKNaadU1mGWtyoEXhpGoEtTf/HrcWnNhdRSERiX3Asx7nFhG6K
DxJ3dk6wPCrPlSVUYsHM+A29EhAQfwz7ZPAeVcLdsoUxYaNOON3IKtFrnccAcw65
CI9NdToS00IEqJPz+SX3rzcQj1OdOxcvczODPQQyY+mliDTVPpYNFF0CI2Nr3R3s
qyubki2ERwNDS2bdYM0JMdkq+0CRwIkYKFD1fndGo2qab5fRdOf5cig1FeLHSfoV
rBMz5nBHQic/wwQYHPlB1WqKn56wmi1rSZeU0ja3NYVLdAJ5GuCoJvb6+8wy1moq
LQtHgxp9NfzUaPKoqkvBkuCOUuaK/ppDKElWdWivd6RGGsxFy6sRbByGtaiVQ0Dj
fxSL+cVnJApjc0mPPHnEaln0opLa30WpM8aphs8G2zFxTLcBstHDqGQtzoWzISph
xyuqAho9XxWxJu4csh0VP3ZZ1FEgU5BI8iXXwWKratvtXbKpZZbTAr2mATrCYE8s
o60evxrSd8GpT2loebRkn/D7ByoRgLlywzNkaR+O0vsoIi1+JgvgHfVxSayMLCWt
8sjGBqIM7Joj1zFbUCQxcVYtmevrAyJ29b9n8Nqa3Ir3BB/Urri9h8ktUBybkYgc
zfQ5V1SmrF3XGUK0le+98stg96UfzGG4aEaI/o4zSfAkO71DQp3FvNRJ7jV/E9nP
QwE/UzCH6LNwgdyMY+zi/iaz5yr2uiUZhQ5BUYi3h5LaEHzVtzdGa2Q3pd+s5XnC
wY5YjuXRmFSzQAFdA45wWv1bghiLBQV1eWmDqH+Ky6qHQ+TPhWocEiKEQ0k/i4fW
BCjffWDslFLxtQNd1CZLsVjwwzBYNNiqn5wQcudD2KF451zfWIIVg52nYKTRk/4T
FPwSaZmYRlTRoOtz2iUYjr2fHXb1a8GZBYV5y8kjoNZ4XBxWpa7UiiYdeIOQAcrK
3Cj8rjZaErU9ZtwdtRd2aS8dooFU2ztFC50ycKCPYBnYmVfkGH5P7CBVjIMmjwXj
20RAurcLRXOJA+6HaXZXiw5rf+xPod8cpxI02QBVlWTrL23mVNwa5A8x7WXxq5Pq
DbOM5BDdi18vg88ilQKITjADFaL1otUJdxXYE4ivIhlLuWMjTn9T9s5fb/0sZjUt
LB8v2EMKkH6/XTu/5EB6m4o/fZdD3RnHEsCc5Q3VVqg/1+dFNnIeGyLHCaWCCKpi
8MKXBDKBbHTgio4OvO5ZlbAoI41LHsAjgF8VGNw4Kvebj7D0K6fbJKzlF6nRMEGp
eQorpbpQz34iQtaQIYtPdQ/uhQmerCGcfDeq77uVu4GWOVUAF28AebCJo4perDlI
hh6nwrLv3lciSZ5XU5s48NUVinOp9WSJQLh0wnbWZhl2DZPZyoydXk3JkDj4QvnH
3lUW68auslSTYc881Q9W1XubZAe/TqpLC9luihpYlRai8Z55j/j2EQowH0/2vmFx
TZPVY+V+0E4B0bdbvmDsP9X48nUN28YCZzVYiS65Edjam5r8GMVwoWfrKjhPrZRg
ab5s3TqItHHiilg1y086+oUEDU0DNskdz9iM3z394OWNMseNjZHsJR0O4JtBqbUd
RNhPwSKi4qpPBeCIWN5q3Q9wAelnxSzcPHHitZFjyXLdd6reXRnWFX9BVTaFNqo/
bo86HzY4QfJmAduJn928beRkR7WezM/0OZ8FdLzMXEBPkChUscUUUzj/XMhngTkj
r7tdme0lTQdLKzMOhHPVsh0XDUoBSgzwnLXY/rfYD029ARaA9zwzmZH0gviedda4
9BRC1ug+Ij8jinWm2NHrEO0e6xS2OJ73S2/CF8wh3siaOpLD32/ArXdXuxcL5HHN
KYVWeqPuT9XbKC28hS9Xx4/Smun/Zb+jCNeyIjuZRdWqRQg9wgnh0yiDFH/jXDkx
swJeLjWjTdmkWi0rkJif2Qi7pKZCY+0RJITuvwxTbE2tMoCkJFy7KX4WgkuJLs5M
4YDXBeNGPvMoNQEmjdOhyk+jpNi21Oak9n89nZN20H9yX/wS5KLIGZ99qj9W/0dD
NyQ4BJAELVOuHpdyrrTPL3xpVKUp9UIKcbZIoE8l6qaLRyolXbTyUdjEp+Ld9Ybc
ROoxKhIrjEOIHsF7lAXuSCd7WsiK45FoRr1ikjNcfjq1Nwn9cHaS9CjH2A6LtRSz
miZZfL04s1vQJHVctbrKqfceG7JWBUMRxoW+/D1sD/J4ULR3V6vYgaVVNqT8cFWh
7UOHOjLL1d1JgI9SFiiJlJmn6etjkmOiE0e2P/ziDJtTnFFTi8fZIIQ+AazNsX/t
682pHEqCgSn84Oej7O7aXqD80gSqlZlmqoBlQtGe7NVZFCUNF1hedcWTjmzYAZF+
GLPMn6nv5AWybvnm3BEGW6Dl8FiA5HVMA6G8k1ZitBovUdtT9hlkqjxtF/nqGqJb
XV3yL1nTzzKnUT2GqpZbUwrqt3VSuMZd8FXRORWSn/2GmWX8UO5HycrLbz2gjTse
ZMSdWsXHFuEr7JI9/pSG3FAW2YyK4tqPvyoBES4FQ7XLDwCIC1LrcsHbYTFoXl70
PUzjkLP4i0aSp416jIQA8GtlOM2LGlyMih5KAQd1+nlKIQgWHMz5gzcpRFgpSsAs
s8EcaAQYf2X5RbuUJozFP9ppHgVz59tRKWWUO8WVbo+TB7VfRxq/VPTbFxxRjo4h
otMSGXtLU4oQ8WqAXIKaquvg+efRZe/z9tv2jMKx85YDJx3dLBTNHvD1LeP0cCSI
9N1bJtgbbIkvGp+PJKRqNYJrbe385WvtuRxHj+VwRmj9QXIyr/hIfjvk3FWwKJuV
Y0KrAT+UJyYaLtCO8Nz2y2RjvyDBSmW/2UBZtqn4drbq19S6JuG+qkoAJhE/O2Ek
mtqRXDFHoCoNjCI19upAZP5krTK1GY4jWTsusBo+FS2rvSr+YueFxtHRV2x++nc7
qQqITdHCmhsYDiM06QQpJqFHeJZmL1vzinUBnFTsKojwN4j8TnsAiKPq3h67F3oQ
7cPESj55Qh5zbmWHwRtwvQc4q5FtV11m8JMp7YYNFok7IC19fC4MhznDFbIgFx6y
bqY2Xhr65c8/8KwnIm2ADH8QZYPNU2xPQ9iUR7aAmJS79fM3Ix7tUIoduYkVgXOl
RXW+Zshfen3zTcNMHImUzlhCFHPky5Hyq0qgo7dLDSkOTmfhf4nPnCp3gmKtlvCN
Gw+N0fRf3RcAsPuGIpXP3tjm/lXbZDI88s4oTFBmtW8g8AeL1tDLtkxOy1zMWIER
TRBKVjpr06Sf1SDcG+dJxEp/iXhSgX4DMbVGvD7v9LNnsB9cemxdt0om4zh0+irY
cTxkJvtMg+PqeG8lWOtlzCQQS/ge9eXfi2IsrpAziIR94MrEPmsmR+bVTeTcFLPY
dwzJEqW5dh3ZNZeaodpXwXCO8r0Bd7BwgkDNdLMZrFUc8vo/isX9mhdUqSxxYUyd
OEVcd+SdbTVpw072Kx/jQIDXkujv4+A6LfzQ/okgz/VmreSDQwufrGf5ffNJKiHv
rOnr6nLUhBZQWhPwFSCsZU0rB4OS5DzOYWOI47LoLTZzQXeLkhWIdIpCIBMaZ+w3
yFH7NrG3ouaqzQJYoBqscQeZCJrDggRZ/vL4nqnftXnIMWuGyDELgR8/YbaBDqGV
vIgRzU+dUugACeih7SjXdzRJeBnTvEKmV3W4MTBGp1D437Fo31438w9rrcmx0PuU
CBChDrdM23jf3FjV+lGAOclFdghoYrA4nWqofDU/CetvRLWOaH5j/OswGoTVaoRS
KtlUI3oUj1qhX9WmnJUiRVeCblmFJFvI5iU08UKGhfl5HbaFOxiFSR2AGpqrTPa4
0f8PBD6p+KayiRtVVmvIm7O0XGWHrDx7R/bszfXyKj0DDQxggybjgafWNUgAvWfH
qNXNWcpdrSGj7em4KuKU9G7Xyi1KnTxasD94EeYy4XB6ReXJNj2npJr//RSWrTIX
J1cNiI8Ce5F35/p5MN9WMGHRo2OkWucgQXN9d9ZVnJSZo2LI9cS3AjBBjV+RKQUP
PKxIXVq1EB34x7lqUM/BMzCq/gZtw7nHbrPVhtweDcXrofo0PBcURa/gGCCvTXbQ
mCQhN41MwL2YGu8wMu9iZFuIe33yI75HKlfTediDWBhoHRWx1/QFQlQjawxawRLt
X4TPmDKLyxFufNWmZxyrGqyZESVZ7NVdlyMgbnm+iLDU/6jAmQlWyLtBXIHgxctN
RPG78M4gfy35lECUo0AvXCujnohYfSB35n6hVyUJhRHHkdaKVkQWPHoR2+pLwyDN
ycEdD/uHldvvMdpHQe6wZeT3KiH2sWN36UdWqW5Pr+OczWKi/7BfJd2QIsVa8cSj
ui1FfZMK5Mq1zXmxAM1I7ncd0j9tPTu6qFbcnhRs/psNVvpZN3iqc5gSIwct7JnR
yZeFksRphl5iZNX0BH7Oxjm4wTFzAC+c4OF40JiEHhLxUaXSrbqxjLR91zyudSzB
gqQA2XmbOKlH4gwmQSQq2qPxR8dBCM9yVZ5fdQVg8c9+zQ98DHcpDqz/PBUXN4vb
zrU4OM4qef/91Hw5CK3K1Vy7TO5G988UzHdsx852Dj8/7M6/hL0JdwDgcbY52Kln
biUByPl2AX20Rg3T/zuARUBaYaKIT20PRM/lkBPDRfIXdbSDDc17NnI6MISN+WFe
DhGLwrhL0Y3v95qh/1AYcDNqVPCETk87bfc8/F+y3woqquBDmgwime93xOFw18jU
ron1MeLa4il3SAiOT2ZduItYV2pAiHSV5F6o28T2f5U0UDOtXv+Z1ICNccxMBMix
u4X/IZoScv9YxOSb++j05HEDhQ3vtgwVlST7RBtSZM/3O5J6iwN3+BaXmFA/wiHg
/eHlBnaHMjtSWa/KDcsEUVsWd7pTK2QgUI+T6lWmmvHdFsvlyHsqGiMgJQzQwQ9Q
sEfbxrWB8GSWzYJE6s//WLpYL4xR8zcfLFOFlpCUZ3+/ItWlc0MTAN6Zn5VvUL8E
jjTkCpIzMIynWhuJDy7lEPv/WJZ3M8sOvwEWZdK22rEgaO1fWymdvwEnvd7tst5S
KuveCTTg3xdKCKefWYSfJNq4c5eobcOYR61caPkfkxpvPZ2QCrd5EzfzCXpbJLg3
+q703XKODCTL6hL6OlzbCyA49VlKF0WoR1Zvpi+9MbjG4Os7CKYMZdvEO+A1UtGX
f4Psx6gYnehx/Tk3iZyOPrAj4KjyvfCvIfa6J2vrwg107bS07oa8Yw/PTgaLAvRi
Hsxgl39HCC8DnCi4vjdx/YE097aQ2z1bFOOVlr+sbILWDMXZUrB7XD92GO4jS46h
Njp/G9xczYaf9u0spjYfwFnPZ4csjZuHnLv57WBny1BEkBI47o45cl//bH2pBdBJ
ZhFqiFGZYrwHvSFiIMDPxf40rLdGOepL1znaaMhzzPgidkulTgVmfJjF4dlju0Ob
FL/bilQZc8h/iJf7YPk4jmdRGwx6i5Nd1dQENLAJtZtBaQx9PhkN875+8XrE2zQ+
3/eF9tF8LtO6EvCThoXBvg61tWvpXU9ixQgudAJm9zWxL4RaXRFBawTjuD36PXdg
J0V51ShGtPOVzPjZ2k+hwloE/IEBkZQYby4pmOUXDnrSvR5mGjJMLlPjmZuRmdbv
nb/UhQhptoMSO8EudN2END3MWL4Yu8AjdFH0Ht8VUlKdx+XaNc4w0okpEXV3H3ym
U6a8a5BAzt5DpsWDk0fCULcRnxphgCySSsAB/69jaYGMqBSZja/UcDhR22pS0UG7
Q/MrXF1xQpI1fDn54l/XxxCqNHkVfZRQ6lDmq/jdZpFcj4pWHkTy0u2mLsIuDUBU
GnA/rY/GTiNX/uwr+DcrJd/VyWAxHgFC3kZzub4dRrYVBgl4BNaMCH3XuJwG9I68
36KIQrqc8xDiXETBscA4NpUcLDlpQuZjM8wYpT5xgnPWXHZfu1rV5m0EgAP5BjxN
v0HPt6Fj5+OcqwZhiyNakX0N+FFMXFF2ehWgxdXl2k06EfYQyx/Ok7pF/KIhPjXz
cTjZzoIWrPN1/ztOGb+8tVhr/MhKOj6TuuicwtUK0UEJISMqt79CJ8rhzJcfMr3l
3kXx2Eml4iip1cT4kbpOH769RcBa8YTCG7R+CFWyPAJbHf4f7SWxRnnphgy68ZpB
F54mfu/cZN2TBnw8bYOz26cOAgctxVoISmoFCaTGjE4/zw27oCGzIvahqc982bxy
md9Wi8ItKOJcOwDIbz6FAdatkCbndtKmL66Ici5MWXl0VyNlFxG/sf0+S20hGJIp
BIP9E09Qd0IITLjlk6E4uVuEtjTmPnjVL2ZhpLbyuIpUgZPCQO1OHx8MRmoFKlSf
EUkBlmKhRjVlF4O8CeGSzAj4kma5GrFRQZ2y1nhUBHb36V2OHwK32wggfy5KwJKJ
k6Iz4a0IMfAeDF5l8/govjo0ZjHOWiTZMHtOnKzJjJuM12tUU0AABULq4bmKJaZc
ggKSpmGdJk+WU+cvE4mckxzETYlyv3gRgSe9z0BVg2glT0RmeMi8Ixn7oc+BwNE9
3tnmwZXaommqvA+eX3JxbdUcGU3cNozp8AyR40cs89eCVp2r6FR7g6XbVen65HsO
1M57o05SMAH+R2H8xMJ2iBTydzboGSJvYNPpzsH5D873LRjKrxi39GlReVY2mN7R
Fe07VGXgI9qTkofcAgDaWouwK3/1arlaO8MONneL+hTX1wGZP0Gy07Smt2T9PSwu
Qi9+rRntbBVBKlmPDzWrWz7HIlvpgHD1NuX+yfO0/ywLFIlk+Q2Zx4GHl0IiHCVB
E58RTWdYLM9iT/audUyuZCNUwH2LzVF8snxhQwijmGsPj+9W73JbroQA/fYhwOx5
trF93TS1iao8Hryp+pQC6G07t1jk3guEHSzKnR2RSlxoDj6wZVoL3hL4d0B4PWiD
YYk9iKft1F3C5Ss3Wp4A91IS/tlvTb5tYD4SvgYFzDQ/2An0cATFlhbrYjlusRP5
PSNlEEFSGYdiucxUd5aB00dtYWm+SUD6dpPrKsgzgIbn5DjBPepYyTRyd9LjqJ5k
vCCSkOIgzSaPc6PtndBVhhNkoP/39QRBqYx4X9CWz+HUS2TboP9oadGZ8eNCgw9R
V0Dg5WTcjvZgyY9URmEvveEyoql6nk+JKUoRKcaLUU4diOYUkvS2On+LnDk1YJGP
gsNfQ+6PFsIvVMIgRmhINc8X+dNrerJmZsgn1Krnjy8jddhgwWbz4faihRIPiEzW
Xq1rOyxzd4vuSasMYr6g1t3/EC3nRMt7wrHloKQjvW4soBcXVtWcuXgV4CRJ5rGa
Ob4aov5Zo79Was4awTWB+1PrUblbaqtjh1/JgMCd/t4ysgwUOkTtLCJ3OmuJAFun
2tT1oyFgjus1lFNUrNQS6QeItTavGPs3JqPqJG4TcWMdzMrwFXFXefKkAj5LjsVP
7cxdsVVSITXazxX7V5tycJh0TL9Xweox7eNzhty8vG7/BMl6Mzb1sBSqFN1MH65l
JfBeqFrAfuo1Qz9QLx1rmAo3rERSQd7kI1cUpkVzHUr6qe8WCMQloLcGhI8yxn3Z
sVgvreStKnysY50IIIVUqyLSQp8gMGoL/MOcRp+MFc/yqCXIOACHnYByqUye+47u
ZWeeGBNSsAJaN3KiW6/Y6qsjkqYRw2KRubZUBW9bBLVm3rAzKwC678wcNvbMqMxx
+XddUIzs40l97DizV7TfKluG/a1FrndgriZW5YtR1q6R722kzhbb1+GF/mQtXhxg
PqBAh/hLKyUa3+CIaQOlhtGYLULfA4OCtx76iLhHkTP6e/zkHYSH4gdmHTqoExIm
L3ujuFNUOuiT4WpQaU5HzmvRcBjM3DfzXLYlvpq9FoxDeLd2GfPOOYfvSVT49BUx
54Hri/oH3kGFGY4QW4QH/qAcx+2Gkta47dqEVfcABRpyr+w1jOyZgTAVyzNqT6o8
jGtfy0TobW+nJ9SWCb5awhyQ1ZnRQ33E4OXT2j1CxWKCF0ebJg8E4wpXOGrEi3YK
0kv/BfwqpQyUXlLZswI24VlougxSO0KcXxv3dXZ0dUvJoCYrq/WeJroCutmWd2lR
9Rlt2fd0vqN1etqcf8IU/M5ToO6s5jwrJRxDihFCRPIW6oTQSwVnE4KgXz9l9z7W
PUIvWc60Qozd2NoNHy8dEx/fFwYD1fVWIY2PHjcc7usxPgKO/r2Uy0E0MxPtjWxf
2Uax8PURCeO97gQX7+x0sgX/ydFPb5iO9KWY6ncoNo5yLlWf6B44ss1oiXSM+0ik
cpCSiQjkSY/ihT22FaNnMRGBHUDvfmux4Tq+wISINCpIHgMzlgkIDRm5/kwOC0Hc
HB0AsCYMs4iS/cdzZ6NFNtA3LFE4mNTvl9+iy6jBLZR0D/A0oH0tuJppIyAtfQMY
r/inkyy+TkC6qc7QJDs+1anXvselTfSDGB7QLLNPvTsr1jEkNuF2+vdgNo3of2E2
S90uk2JZPhAS+O6vfNr6B4R1Cb0Afkd2+CtI+ie4fp6riaT/fsSwHX2oljLinYHt
TCUvvs3KWdSg7ajFfrm+vNaOXiJB8DtkxDXqbCRRpbjTNiW78WAsO3mt34yeofA1
tSI6daMx/A2q/HypIeahcBawx4lLefpsNJ98k6p9Y1vflr/hPLDZNs5/iFOuX7qW
hSJg8cFPZGofqRD0FnJDTChlGomAC/ArsFBg5TYMTd3ZdOSrv5raEVzfa5Woxu0Z
nEtoyUBxizLWS5aM+3dJgfVWFBenz1nPXLTvgyKoDPA06YIEdlFdPdNeOBtYISly
92NhgpGrs3ghdr9PRW5EFP1OOVTAlyxB0fDcirzmKkigfkJvJuQEZHhNj6K6ia16
NOMh0U50coDWZFdXam193MUBdamjBan18DOEkRCEp/HLrdd8ewUDaKU6iF/xqE4B
FE2YXOJYuNyZy/oxn4BtQlalvhVdXpzTsoeT7WA7H7USpJgysedY5s90MfzBauyl
+wy9u3I4l4EiqD2tczmY5uN/fKgreOJT9msEaTsQlukL2q9TmF/50ytKIOfThNiv
E0AEyj5C/NP57nMlFxWcDQTQWjWAlAuYJR4grgUi/EoBaqrHhJs5A9pfn29xnEdU
QonHtnzTjnOwzPQimnhTmMsvUPfslFoH8PHVWHJijanZ/t+q9cUROKE6eucMfyNC
hkLjJxDFVLMwCRCypymhH6dezgnWu9dvG1ZOMUZyf3fs5tZb+5pmYsR/OSflm4j3
jz+rpjpLPFGFfettCaf8k8JeOftU9z7VTyxivscfE7MkXITVoh6jCMClbVO8Gs4z
glOyrP9BD1LTA8DZzrf7TaWBKGEcloDlIM96sh5WdWEWJ3nE4mYP7Xth5ikVmX9c
QoPA7UiXkuJiriZeJKmlyU8l3CIQmEYQMW7jAy+knVHwj29FWM+0Udlu7w43XkO5
9PoFl+vkk3XXjteI4UcPewRCN/iUXF0exnXCNTkeWbeSiHLUeSTMSaEupoKqXMqs
LxAspBBeEqpbUgJnDVzq1nnif8yzfVGa9CsMhcX3BGB7x/YHvQTIfLjLK09Jz8sV
YsHoIXtbyLAEk4u8AqkS/SBiYIc+6T9nAif6n/cQO7ECfJgC+1/KCloYJdVg7MPX
uTv9x54iN4T1DXeG6jaPtcrFHSxi1nJcIBQqBsl4eVivOdR7FNJWWd2+Pbpcyq/T
MiV2oRVfnOdtfD1dvq+O3+yLE4Sg6UwNpsKsLIXAACL/qVD9bv1HV05sJtzxgUUV
PXLZiylBRQB6waLRsnnMkAJG4x5mGRjiiGbUrC06tIOEsAKrAUzh+H4Uvxpd5TBE
4iOae3tic/1laqf20kNooPREuXOrE9u8yeSRrhAt/BzDKzhLkCt7mSIRCaN4i6Ap
BJ6Zbeusk4Gykpk+M9wb1jYBUqnGItTtTSDFtE9Mhg1d44LbeL64hTC3akpW0WoH
oWPKUewFg8MFzHB3Xd+Pjct5kozkSsAlYGJWZvnetMQK+Ejv1JbxrjC3w2cxc3Og
YeGl6TsdW0okcnDtgIdwyr9xgX+sa7TVnTpPICwM81Fz96TOhomxY7NmOqhmJfJq
pGrairA38FGAKt/oqjHFF4jezWC78KKkj7tNLyh6K6iEJ5pKlu0PjfxJf4+GLEro
mc5cOmBUK+iA2FPgrk2Ap/BAGw7o0txhRoZyxf0Eg5ouxykHzVc57qDasYmcmHf+
UXeoCOd0rWl4cS5sjY2lygL2Trau4OOzk39klBZmfI40AnvRNpNURV+32CLUyEc9
aoaE+h6MNqVi4tDwy3v07g9WKhgUZ7rZ1UNxnJP5z/uhezcRfATt64dzaML5QtDt
3Awz0QuRZayh4aUxBwa4/4M0//aWs1/Xb8aUu87qILJfsqmXiSHjEYptSGui7KOZ
f59lkqZq3y88W2cbI6IFHjYSBr+wQD/vyvedXv7DLF8jhmbOFYMurFiQm3iFK4Yd
t34hHV7P/8JzPHMdmLMWkII9CUH6hGGplrcDZhonkwfr3T+8K5WpA6h5nz5P1riE
FlgZoF0wVMxkxZudwClS5yNgfkcbym0KqzSfkNJJVvW4LUwpaSTRFr8aUDV/mqdT
D34CMyuS9sn2ny1DZto11h+gOLyaTGqa/BEejClx5b94qG/2LSaJJRWOfYjw398u
9WPPLeostPE5JOcSZZf0WBUBtyi0dmf6QK7mYx82v6CtyBKf7cwpeIBp+MnPXX1F
Hp4ZkFvhsLRORxp8AHZ44tV0djBzayAqyj9UHHhdwEetC3zvBlstPZBb60d20krr
cddc8T0KSA/0EOpKZmpFVu0Keqy0kVCx/XsWa9jAwcUAM/VEqj61pBAkOrEhO6Tu
Wk/t92ve9wVWbvUtiLyYN0E52Mo4l95ZSdg8FDaqPJb41NFFy5PMnooqWyFY6syD
NyVRTLIGVdm6x9KaCbLaQhTrISWEs7Q1twdYd1jiivpoCG3vZy6mlrv0/BWtTLGZ
mzot/5CMoK7PEtb7JYnKJJ3Yq5u+FQysWtgWAqL3W1QviISUNqgnDCPo/slATJmS
szbSHs3zmx3/MkrXBaIP+6IouqDYllpQP6jgbEQyCk0eHxaiWn2DoXDYZmOZoyb0
VP/RfBeUz9upMV0qiSYXdePtRgntvkAm3OA4nAnZ1HOU7Z986fINP4oB89uxEcNn
M/vjSPVZ9coVssm3L9zq8880dPQsZ9TEQjOo66va8KSr0Wv+sRbZYNKQIetiC3cz
xPsQIoD0k2P+C/Zz3vD3P49uvDcVaCF4VS+UX4QPVqFUk5qt2l7yFEdCsZwu/d/Q
pPQOKzDjepZLISmXXa8L5CVJya2AEh+OkSCjNeLHx9CpT3udtaN+ay9NlgJrKWkS
Cj/MLG3fPJlacqJ9PIaunx4NETne+revRyKt2zFzFkcwKEEVvBhuuU2w+pzHf0X5
aWEEt0e2gZNySMPBMOJWKfBE2mRD/0Y2WYVxJA/Op3VqdQqtnLmya4gFeoJ++mxn
Wzg3CTAQR6aqxIY3IC03FMRzDFHMgAzXIpmwnBvBcdjINnGFiZnFieu0SAr5iTNi
YA5NgZoR/9P/HjSCitN1y5o43xsQPWFjDNnV0DAgb4qj2/4shARKtwU7oAArqyAN
/pXWdHMUdhuOl5hILVFd93A62LTrGmDfZT5xbCEhP4UhtroeI4yzFVq0Wf9PWW7E
+lXXQgElevvZ+N64T24L51f2nQvtT3qfIvw7e3xbUqNpcJN/3MVTAvLR9JKCQNhE
RKO2zx/1YFjv4W5epBziThOkUuszwVPUnxmO3NZ/OvZiib9CxonrUKxNJktwCv0U
BdfRfflPOsBG2IeLVsOw6DuZPeLUT3IWE4tfyuB4s//wZskrmchfjckAMkJjHpJ+
GcAKrYXJzwYe4nbBkhzY/cRXeAl6bj1BmzHk77eWOd0sBHBozvN5KJPqkBcOaveP
OkMb5qlcMeccSROK2KQTKveb8EDFdQR4H0Axv2fnJMovJhCN/ij/n9VQeSf6VeUD
F9BL67/E2QrZ5GPvBGetsbliFe9eZ0Eq6e2XPcdSQXypfeL1YGFGIUK7P2GMcLqA
pi1X5RZLY1ulhlZ0E17uQ3RcurKXPaEymKoJLX6eakhrZrMvAO7NfuGr2/ffTW8M
Fc+RuSbCg6mtJxQKrITzA34ub37Fkmqy/5pgIjnh1HSGysdBDVQ01v5Soo1SXpgX
qSgFVQlRSUg/A6mEbOE8rVIuWs/qf/5p1aDVc54ooGfCbksx8sN/XD7dgLRPmMtg
lSJ5H5qNslpxOnA10vlKPdaDEI9jwFc0c0YAIfUxDpgcd32P6PYiHvQR5GmLAWyg
em9wumYV8MCBy6c7CoeSzl6av+hjfakGqOeCfjtN/5BMup4TBabKDNZEKZnn49pZ
LXuIslyKQmbVUukSuAorPGvQEWuhDadQmGAZ+lgPDOFowwPGsRvIlp8Rx525/PZ7
x5OTQZSEaIiVVi+0KcgTjQZHp6R6Gk+U73JqiUngXkMblu7gzU9TogJSQIEufRXw
rxrpw9aHwvNYgpsxcgfSsGwApw69ZPMN4U0BcKhmkQAPdziP+aj9AHQrUOXu/LRC
Fn7GAJaKHGr88hH6u6sVBKgVkWI+LXgXUlTEF9yBjqW/Iw9S6WYnVMx+WE5pGTCi
7BVJ1FFwTpGkBBxd70RvdaxNBkSYw18cK/0YklrqvEYm0Rs9PqAfwzctM9C3LSHt
KTdzglr23Dk1Q4OVZEICLaaDLkdDCdt867ILOPWNr8ChAkJr2FxYQLLz7jP+jfj6
w/88pEvwsFbtgTKsGqa4nSnJNUTRZtMLw8bH3qYDL94ZgDNTqIRZTnLnf8011QGE
fhacw/SiDKMDmzzzAPj4hHlI7G+EQTH+n4awP6uUHVK2hglh9VMOX0vL7NKkfTMo
SnXRd7Px5reLlKTx0I41tWPWcFl+c4+vrhwTmtVxyZHuqXci/ErzjwQdlQlo6tX3
lFTK+7ECPGIEU1vpDJqXBBYkDBHAsVd9pgwuk0J0kw7EXZxjIA9+tfMyR5AEJ5SM
fB0+804SwPWICSqQWslf0we9JE5BASlsmpbO268pYvLAUXoo/ugb/NFEC8F6ZyVP
tqczhHIWsksEOHDblLyi4zd8kkfjC1MiC+erZRHacV1TlbzEFKybD6y6uDBG0TU0
m7BJAQ8852SDzqoVjphbQ9XS2g1fFK4qYu7fBrMO/JEboe9VGU2yzimNSi/wDyTN
kOP8uHDP78GKBq2gOxVlyzl+kTbqzAzgUX4vFGMCarZGIfbvI5fD7C8o1pkYD9G7
wDXefkKjyhof2N70xBgbA6a0RUK87El9wFkxsfR6LAfvsGst0qqSsQ5meZSXt8xv
QzjT7IPrSjc751gzhiylPpgQVnsBc22jF0SN3HgHzqcfAjrKGhlsVgBHapTbq0hU
/gR2MrbTaCcLFCUeTGrHn3Fiw/PHrfAcwxGRKDinBzeaLRK393Gur56r2oW3vAO4
C24Q8AMXSiUXScbkt8EoWjG3MtFsJH3L7DzJ+wNv0L+5MgLjGtmrnu0v4UYlU2iE
09vW/kKehlDHA/v2o3aIexOd4Iir4zRhilwAcgPRGSodxowvsQvCc9etgj4NKeSy
4KuiFzsaMZq9Rb7amsj3udGB+0RtqN9ELjGXDMyMS/iMW8S/l4gTNwwCI0hi7RGV
CY+4691XMgIOMe5iMlnKWKFGWtVePoHzDKKRAql1k5Gk1hYrR68kXIqwU8tylsfy
+27Nr9PkDPXSaIOKEAC9NZSGk1XmPaGczeZRn6BT2L2Xh62A3w8dr4cEU4od9KgJ
kQP2RoptttQvGi2qC2zZAuwAurU1RCqgY42AmdRlnv9vjJ8FOkqPsR4f1Wn9Kal0
mqyWVGbbaChYPj6zZ4JZCp561/ph1pGBRzPuLolbmWqQorOGbmhWbMPc05OUEefa
hycLpNG7jcQt5GN/uH+TDrIZa9DEgHYrxvJ/fc/N3MXB2a7mpfPFwNAN44XffZHY
fi1vSjUt4zIyxDhiFldh5lhn6bdDcONcnfY5Mb69LtR4cpLnj7E6gKtGFiSM162Y
+jY07bYy8adI9llHS/OSllwzSuDKkHlRdr3PDH9LsQIilZGmwjSAJCrBPBxfJeNG
Bfgd0vHUjqnXtqKXIgiDAeDQEj1acFOQVbtNvyhkKUzLAVIZt85/V++429CGIlT7
EgVXYXl0Gi4q6ZWBQy2sDwOWAgu+t8JxtT4vCMgEZKClrbnP8Z8LlTRCWyeE8Z5X
AOqA/om34JrhUC+IK29CCAFiel1AWuGL5cVkN6PuWnOAOyw7/y4CA+Tkc/NNVcwD
w0c5QOFhzNfnQTVsytB9q6gwXEYy2vUevEVaR2t4Epr4rPKDcTMfZtZtuPrDiRLZ
fj6NwNSReu/Ouquabmr1ozT2vrdOTkZnnPlwJ6uSOtbGUBsloREJOLHRIk05aAru
HkRF+LwX7xThfbsgLpc+lGv1CxgkDhbagxnRwYGvslEZJxZRhU7px7gqKPffWdpR
c9vKFv9NCO+9kAml80dd+ENUAghX7Dlygd1bjMc0VN4JNdlE+rwDbp6LjxRtZcGQ
+KBnRBbPT0/Mq1uroqHGxwZ92Ab7J7lEmlLBx+aXG5WEvk+tWHDQppsTqQth07bC
8az+KhVsdWgG4oiFT0r/cWn8KSAcRc1k4OZGlc9f0RpOy3mXBM516Q5IAsR+yrzA
2nQRgBV68HvB95hkjlgoH6bvbul84kPrIQ6ncU9LwlFbRbJebjj1xfTQMGIWAP5o
dTSTGBC6WBkL5V41vsuwYoNrPYHhQrF3DmRoXTI63K001OJbxH/kJ7G8AIdoA34p
IUhR2GhKIjxL9qrDuhkfgnfMcO89vPuctxa8fijb7pxpim+A8+JCRwW0sZh2DvDK
VUY/WGbwd+Fie/6TOrDsPXdPup4frWp4NZrm3J2/FwlHKG6myWV/g4JCLY57lic8
Wr5uNO6eoPQUH6j7fdp6WtV7plk7qSsD219y2KjW3H0X83rYL6alaN250VdXPj4F
VUrWN1u4a8xO/cpEkLhdcELg2kXvV1+O8MpG4nEqT/Sih8BFaf+dCr8p93MQo9DH
8xLD3OzahrvTDhsNeweNJxZMrBKLivk9Dhra65izTo6GPQRioHcvTouWlMH45nlV
3mJPzVuW70AGvOb6uLBbtyq0nmgEuT+rOtBzY+RSAxPY40L+d0XROallfX0tHXhB
SHZ9SLn+hT/PSSYZm7d3Ng44cmWCLyxadEtYy8p6KUo3Y+YfIYhVBKfmW91FVCCJ
Bfu1viPqsEVsOjc8yoSupbGdLekkc0STtC6ewpUqbfb923LXU2G73EaFgsQp9zb6
QB5hKRQaZMfvoR0pCMTN7WC1fhAoy/Ag6FT/UEyqwZU24GhKNTh6EquESX/KoLPc
lF07KMwdqLyQ5YmsMoTcMO4NavHp4j+8LIf16V9ZmAAe5KM8n4tJ1kx/gg5aiuKj
Y6KsEDyS4OTGZ14hM1vwZxmJoBMop/cm1JMlLjr4mrEDmHg174vjFJ7YmTGVSBeC
raFkKoIKcDb8xZpdw8bAzas89jVMl+7CoS7uDBI2/jszbOdJlaZ5ZFA4SOhmSxpb
mKKUieDSJirXxDnOjaLIOUdP/TwFLh+RG4qJEAz6IVnbazIKiKJO+hWE8p/+MWal
LrqeWmWGdRxvqVNV34Z+BFsvsuq7H7mt6VtgG4+KWzSaX0yiZMvh3QQOxLt2l+b8
ErF23qRLZ83MTTU7mbbY4BoMocHljOkXAYQ5YXOIFcp7WxldG5hkHOg74yCHXD7i
F9N+wxJVJRPqszi7EZ4Q2s4laFJjndJZ7zCyUezwvflE/HMl5fWeKPr/AYos3v8x
qwfRd0HN4pvJ/IivTt+rTjBy7s6zLv/0Foe61ip9Nv4EiCsVqnknTpdZbd4dqsAu
+EoFAqi8YaMEdj5mMbY55+5M2u+rFlVd9TDBsZT+EtR0Yo5C6qieHfW0yqLs/Svx
7GNXPhYvEgwhHtx+EZyj7iS1iAtNo7T/qQxfbbQheYrAECu7MRD/3U8ngTuyJNnt
P0zIGUg+aFlyZcUHfa+3l+PLgDVt73m2TKGXMNFq+AfV+T9gpgXkiMMe3O0bzm5X
7/ZAOxrEZdCpjxdgD21lCnI1K7/TRVEaoXVBfmibSaVh81bMfQd+SJr3FYPuFTOd
FJcO7kySCG8rhsT6fqEdIdFM5ImS8qIIRg1MYTAmbqvVFLQu2dEyA4lyTVS8hWZr
cidVje43Tndq2H1veeHtDdA1TGx6r1U6i2O6rzr21RSgOcq0kQWdn+9bkK/N31o8
YfjNNWb3ZhrpsQ3hQagnd7uvFDBUL+RETbtarsqjiSi8MeHci8zm7TLncAHZISUs
tS2rY5M0xrTNALvs2pklY5mml6Az77CoUJFjBD8FomFY0y6i0Gfp3Twe2lRixWK5
YYsRQtUWb5lRXx683JRcwTGetSPNewlOMyLyAjP3fabUsMky9Dr+JJWwJpaTfEWu
1LWcGRezLhK/Q46WHrRVSZL2WDCSKstN6f9stwTRqSIHJ7KM5OXdBBE8/ejnuPLl
aKPYAa4bF9KhSiypgsH7Y/GJgFDWowR5ZCD4+UDKaTcMouPV0crLRvpIW6IiDVG+
FJ/vR43S1QzqeG4zZZJNuOn4Uf8a3xX2idAwPKIL50dd4HVlRXksimiYHxx3fN3z
WZDrv81yWIiQFddX1zpvMILBkCyh/BRAxFDws1DzfU5Fpo9zyS+TsO7XEHwLsGDC
8CD4akcw5/sUUokpHXVTBhXXUxtDXFxlw1+iO23XcVnHl4XDXiMG2mG68Rpbbujb
C44yoJHN6tHRML/jcQ3JzefH26gjVgc2AUHxyW8748m/8mDTo+P4yizUK9W5zbdj
bgV27ZzgLKmilPZ0ViRzJkOVzN+FtsIB9ap4iILf8BXtwW7WN1n/P3FzvEU8DdEp
AOQS1eYMPCzE6cScNTvi9GrjscYSt+AXW3E9/YApvBrB3gz/sSMGKiDlv94TCnKe
qdklgtGArVaas4/vhecaqr5Yf7rhqWB9XjzUIMKatW1k6tDU11emH6RKrpt/MyXi
sr1AHDRge49wdzfUWpp3s5BW63Baa+ZkneleXV03wyBck556pwphbu2+EQ95GBYt
ii94xGUNUKeUfmPNU7PXHvT6X4b1R+bEPHS88VxEvMNgAD35gK2/BoxqO0WfgF0V
gsUkPKd7aQGtOjvvbOTgAVZN3yYLhrMKeg1y93/UiDK4FfnVGEvMED0MCq2XLA5E
Cdprk7LWxFvhKGcqExM9G7hcBTS2rYK+qr6pqzO5ey6R0M1T70fPGWC/aHeE8b9l
KWTOWKd8WQom2xiDTuCU7pynvVTCs6Q6tnn5pA3A1viliMLhmiRyfEtS1tYhlVwO
hRnwBTGvXie+EnrQKAkFeCW2Q8t+AnCQgc9tCLAPdDkLwz2y+nSnDjhkuq4KUvlc
C8jQm1O1GRD+7FtC8YL1d9ItKSepd6djA0S5/iiNrXX72/GlqU8Iul1AVq+NT77/
jPEftZoZ5O+EcYR1kM+hDo21EgWkWjYwbjtnE3rLRHXNBFOvUq0pwSCH8Ee2yXST
QBWKeUQgoWCSldhqp5hh/ZISK7+CqDSSecxfAqqIiI12DkgtbX+UZZd2CW/ud4fD
XUmX4mKxQP3YQuZ231cUz7rIvOexGfPegjV3NZpj0LOa2PqMs6f7Ugr6qfAFYRGw
22ZWGAIlXbIFwvXGfv05Bb+tt6ULy8e5MW0T8/BeIaRMnC9INupIigS3SwFN1BRZ
3V7w/TcKzFI5cPtOADPcLxTtUv/4Z/GqIBlibbsBCUR0LuD1ef/jPAY8/73OW1OW
Jxeow1jCfGHnUWsfsjmvOwwgp1UGdJbYooCThcQAh0oaPS9NgWFOMNcA9dLiX7OP
G0Oh8NfkRuGKjDq7rZGv3OntbN1DWnrUAA64H38V5F9JO1iRqJUBM532yPsE+Q8x
FWxl+vtsFcMmStTbmv79+68hh2Y5/DcgRMdQcyKmuYjBReaVvqqceszuJkkIUPvi
fUL9Ma/G8vEnVx5ADaUJ5wuvMAtTTmMV2zXc9Cd3JYx1B59xL1hX+80pn1t5Apno
QahPtR/aYoHVkA52l293d6cLW5736LTmVJ7MwqkecliMg9cypnyGADAyC2c4/UyD
RbdgCvRP8XnRYoIct245zBmT/4cO1q6H8qZuahTOdF+ORABRTWKd2tQI+yQpu73w
F8edpOX+nKXoPJbn6GCwiLDuyynZDIih+Nu+dxaMbyvXLm3lOCUAP56ZhBeJztNb
4qF0SR14SdUuPnLqSmCkjp8tgwJ2HZh8QOT6OXdC1bsvyaiK1QanurGBX8cRFc5R
Vm8Mh2Ol2pxlEuDuvxq+ljvqqVhhMepF8Fmd5A/2lw+i5xwGPMZviagQ5Fgvk7na
fiFoo5LbaTXy5r1if5lfMtSTVXNTVqa87NlFD8fRLkWHRBlKK5PnUZ2QxCE14X10
rCIp8c4i5zAu6PggVCrw/boOZ8NDX7T9iAkzqIFKN74bCnrlQVWuYH4xSAw75/mJ
YzJS167afVdOkicSsmLnbtqMV6gQW5uotx7xUYalYTyryw0teMCxiJ/rIfQu/4cM
qbCW+x3sX6lLCS1nzi6zHc3bu8FtGl14KtAMIWhipp+yVjBraWCtQKWpQNoVVCep
36BNfc1hE595oyEDHOx8Qf7+0VQkGHDoV3qHtHU59oJH14bTH4aFaPYrX4YsKCpK
5fNnG+fuI3RMRSTe+jtqGnX/V9tVR+jCMIWm3m456nxoY4wsYmDLCYlFXZdV3VGI
4NvAKYy6HJIFPqxzYIk3S9XpGEAWUtlySUP0hQJDOVOWaZyYXcfbn+mkQqOpKn0F
uJePywQJGlfeh8mZyKwcu+0crBZLHqELfOBjoyiEkfKwAxq10NjLcWGM3sfIwf61
lMTLZSueAt/8jgrmQcw6eEBpTWyq/8FBQztZLKsYTJznqpBbZPGBa7EWtqDYuub1
nIw2Afpc+LPMbrhNbT9GhqS4P/JhmFiVK5i4WrTkQoluKPS3nqrhRrmYMXLMyXKE
2TsTuReZOlYU16MBL/fRimnVrtnAKxDRxeWxtrIh03SXhh3dRzQTm1wN5qD94e3Z
5y+tXyUEsqpmEOzAGSwso7eBV8905WF7joYFtvfHRtlJ6AIIeFr53SEcMXf4Qsyd
w7008y/S4yfhAAR/UEFvfyn5RYoR9c/PQqTAC8zV+CKEvSvf1mMjYetDi8I6jj+m
ZjYXDDHnbApP+7u2FqR5bKO0gSUcEC4LPOb5vUyOl1vo4kkcu5lt0jRDsofht07b
lahRZod5HuKZESV8+PFCoKIBxqGfL0+eXMZYcmIo5K8UdkOINUV4mBGnAXoAEyNv
dYTmfxz4xda3Wcf8SIfp/7+evyeXHik+TNwod7o5Ww93+7guqncfXqVnpcXKNy5N
eaHya2fsS6N+AKqcccZGZHpVOjX4lX9sGPrpEeVty23wsvptlyhM8AQalkJo62vx
ZSsB0nkhvEPA+0h1iF5JAiBo6chMzrLH1R7BSOk24+IGtNMBf6WLBKeJ4X79cpcC
OOpKlQg+e/Ku3+Ad3sfh6vY/GsEnfx+zWDSYlIEKVu9MOVL1KHDNX3IILPSieAGU
wkP8es0oV3pZvWv25YSVEOhkaaWQ9s/UZuYpNtzYpZMQqcoWv+bRooMBP/OqIwvv
3XUySA1rnCoXR3fGdE8CUwXf43O9ZiXk6Rh6TOMnMhMcHKxqVILAII+Ahc7uFBqJ
traWJS7gVzB/fmMnGsuZ48jXMncPARx9+dz9NKDo+gji7Mjjk8DTgelnRDPP9gCS
iOWc5+7Gr1Rxh4Lto/p9HhR6DVI6wsq8qacGIwxtWfnEb+bDcM4IqhueX4wpDT+v
Rb6xPNGTKAZOIs+HwFAJxUO/+wfz7+KI2Fe7AvGbC9N0IHE0o8PcuqcjnQZPEbDX
mMwri1rxpdERYarTlyBHSuuSnxLqc22OBI6LJQt4o7dVIvaZLN5OjuALNWWpSdKF
afnVGUSBbnypiaHcDjAc1GoPOzTVWI5MboTIEeIEh4m3WjefyYFHEKwTGi4DExNW
0M1XOt5VEWZFUGcvIvAOSjr0UtM/aDiytknMNt1wxienHrMCzMu8lrK115qrMBw5
cNJD7gq/IraHLn0nRhND3NuAWs4nk7lRUpR8M2z63iKLwHYhFoAi+ol7JwHYRAmj
/q+N4EzRxPmUJRBgLK//qa9d7z4eMs8GZjfmwnLOopp8AKHqov/mYhir03RESRIG
Y/Q/nBuX6HGRvnh1rKh8PnVqbAWTgZoZVLB/kYDQ9afwQLHi1nmjKLBlesEV8Kuy
bG80adA04IlhyOXtZjwsGen9hUW7IxgbnzjLrEIvcaqRO/ZxNnRLxQrixjdZ4jE7
LQoaYAvSHnwlsA0aZK1vBR2TVCT8rQaaxzalhO10RkFlKJw8HzVM96k7E8UvwQoW
yWDNXrvWJSU8fp5wqpCosbZCZBGP7YFgbFvuqPd472I+zm72YslN3/uuMjrNkUbK
lQdz3q+aSjCz5fFyjX3gwwmBCOrJGTepOjSO8tfgbPN7s8WTFRCv1WiwWqDNjrnA
B1Y5znU7q0io9xnN0zcxQvj6oMgbUndSvvaqsKOjWrJBfYteZdhjgz3WWWVlv4cn
pbZtMb5J6dSTXaMbYCmgt+mc+i3Dj8gFtaDnTSBsYuvmX5+XUKjb8YGkctKRCkPU
BnhI4vGU9eiJRz7QyQqm3ut4H/EbV6cKKSDG3O8Ycbay6n4WonxK4pzm5QETqQQ7
F7UbCIL3SZCQT3+OG9ofOTSAfp5Ep2SCvsczA0MLclWzi+c9wAEfssWWpYicKUK0
z5Ojp0Btq8bImiWtxoBP/lkA5F84eTakKk/TO8pQ9s36W9aNLwbCb+FSqlISUVa9
ejFkphAk5Gssz6VgAw8xkQPnztvxJzgscN0wxpEViIoitfPskTbDDbGGFKL7xCSf
ddtFcZHvcJr9M6RyFL5IqWuDQ24X1xnAfD/qDodBZaJeaS/9OQRMDmupVf/kq0il
saf7XUELpX8+B6IdwLPxCjOB9ziTrxocTpiT/mNkcwS1rmKiiOkJCGRzRKokeaFV
SpJ4cCHOZQpClU3UBiNU5OFppw7tCFXCPZiUCo1i17p9jS8JxVQzWqsbEiyLTVqF
g6pKyAcCDJsq42Kj3dSiinvM6DRbvLx60GUud0mEOIlesCtpWL7H1ZoIR232abyA
jcyAJPSBNoUMjRNoN7D3crN/gDhWRK0SH9Nydpvt8Tl/01PlsZ2lRzCD7LhH1EKx
jNAVg2N3yvj30NzfSLhBXTg5dmsBP4vYFU/V39hFr3uSykU4MzP4RnXiMWggFjb9
abKDIiDLMWdRtDx8Kt17gksUiFBmvYptsZC2UH/T8kV9/NtiTQH7m6a/nUgZuU6l
TI67SbpwNI12UH+bykvy+CveQHEwop8uoYr0l1sy2HbZxV4BpZyN8H2J75rKAXy7
R/SIhMaG5ZIaCONAXh27cDknPmY2hVktgD+6zWyIev4bAPONqBSANGp+TlkMlHi/
ETqHA+PzLYXitPBG3teVgi+w5omNEU1leXj+GfUtiR8pfJTFuCbx4M5/Etb/OqNf
zzJfhsI9f4/B6hgdGxbq6qyMQjRYGF/tLeFf4Tb7njnU03MztQIupa3tlU/fotjU
G4XHpCebirzi3chP4Yr7LybjuyZyWtvsNQrYRRgvoMHsbvmtLloPcBaKSO8Q9hMz
EUCnAVNc1uANPVx+JzKn7jvDnqIVLjEdCXMNNQE4RPxbMhy8jEyTbjiYwA2Kpx/Z
61ePe1lg1OwigUyx0uww1Ff/7mfw46M5lUVXyddKTF9UP3Tk8Qg/wiaNoS5A+Z6y
G51VVs763rZVHcLmrhZENkOZFT71SDqrswAk+HlNkHoq/g/YfZAg6lnDQiK7aF3B
3JKafHuySUxm/MPiZsKqtIQKRsGhzBxVsmYkyx+Fs9HxJ1YS1OlUNedYLKKHiIH0
H09OCX3xvXaQlTOMqBuKGrbITi90VB+6PS28n/4cvVrZpOe5l/IxmEQ0pRWYfPco
aCOWfuNW7Tls5juQgmLcb9j4n17CmQ/M64x4zEs9GFzmPi+ryFl/SopeMd9S6WJ5
iMzFVtWgcRIcNMiJoPLjpr2RPW0cGDWJmC7FO24Ait3rozawCRi+T5IU03DmBIhI
AJH0S+gOdfax2vEY+QoBQ7VgHt8MGvuEW8LpGvk7yZ9ft+AQhHZoK+fbBrKBuayo
mnbCVvXS24NRfFvZ7UaRC6hkuvqyOjz31LLUpd2sscKpcZgLbV3wOcPuI7RCMgnW
OioqxZEP6VCRPv2eQa8jEYnhItkB9awbwIIDwndXmO5fc5KXf/x61/oGeLLGHG8O
nrXVTspbj2i+LHRM7+axBtzn4B5agbJCU0I//3i3eC2xV0rtMQK0V2NmLjGF7707
KrcVDZ0Zr8JCPRD4PM6IjMeb86XDW7IPf2V02i3KmizI00wfPO4R4O/haJ/9biZF
/D+cYi/eqy4m82waWRvUOvDEgZO92XdwFFbyoVToDFsPUh4k9JQzWuI+cjokO1vh
tuIH54Ci113BeJaBMmCmUuOd0Ts0lWqc4ggHkKnivOtIr/P0CF1evS6YElm/itwz
BxuNgZiPVwCM4lni1PWM8MhOlIFd9imVk0Oi8QC1QxwiEesW3rg2Er2YfyLPFlKN
dl7cDFvdXmB7rHcpCmx0BdVhcaVFnPggmBEYTYum4DN1v7Alv1w6Uc3oPWA2R8EZ
grVXKxmcQ4kD707qprQoe0fCD8PN+97OdeJeIQKQjU5gspHDN02bW3Yub5D3SjRm
I/EfKBFpQgfj4iJ4TBdpA5z/yC/3M4wfEA2ohGnPAYIs+ZgjNzeA8lOTRf0JlWfX
gexTKSOQYydhuCbqhXRyW4Ht6QK1qfq1gGyDZQHOhOVxvCwzD6VEH1XywcDWTM0r
gWfuhwC5suaFRMEpjK7u+2ntAhFlXI+J89YIBmIDuaTzyc1A7vLWY7KgbBQNihIb
wYPi7/lcKCIJjPup1xYM+cQWc8jrWeEsTg5gKlaUoS0Ud2IHN9pHXTjAKOaIou07
PJ18Rj31NssSEMqmxpW3hz3CpKoRVSNxEkaPAoM7CXCNRjx1hq53zm53PdMrcjCd
K1hmpIoCpb0T3uxGXkV66ZdaX1Ta7A+BXQA/Q0cQLaIV5UYcaX4wAlS8xReF3wUE
Ckmw7ABEw63gDf6kX3GbaO7oauTjV0D4TspGvPm3/YkoYiukTZldnPKBSPOA3blc
7k9Qpqat9hCmgczm9gY/N47+IULMOmvhkRp7qDmviaAPaCXE7T6PrD7IvP7aQsLu
HIWi6lcCxP1GMOeas2geNmo3g2tKvJw3+q8mMFy6zdA0NcUUNhDk2wqpL/oZPUXJ
zEVxKmuwRv0IE8/C+Ztdm74s0jcdMuvZXR9Lor7BW0utIUStMnyEV9JoNe+cKzgR
j+UEdRxWjejT0EOtb5mGNq2fseh4cec63eOtnY/T9cSkMO+1Jlx1FPQh0han9LOH
MBlGHTBP7UycBCgcHYwTaY+JqbOYCq87fnlOYIcYvyeam/TCeNZaWkz67MWok+6r
Cpt/61QqH3Jrdgn8CcUSliIs4tt6FlOJjV4wpeJKosmfHJaWmrMD9hHh16IqTR9u
r6/feAl1Md8ACyRU/qWySmZtrOn46YoSBm42i1PtBBkaRSfdNHN7aSGi9KdplOk5
/uuYnrlwvhD/4GTjbJgEe6TOUJqWUlGWEosQ32LVatpp3s8m5RDx7pnnLc1QaXxi
xp8iCRf8NPKf/P2PdRNrc0US6mYQlxRS5FLYKjXDtdcTEnuo18pXVexDhLBwZTXy
u93Uin0Mp99JiIoFi+hFBDDcmUgIV5t8DVs/w4W5z+bl3R6OGmO84MG9H+l9R5wf
NajIX9MentQkWQYEdBceWGCl2hVsQ23wI3Z1tPbBpxjF7hjBeuMf5uP4y6KkwpIP
zgsFsFJZC1huRD/LbVgCaaCTGVGrx1jtQlo9ZhKxpfdrwebw99S59maN41Hb8Wcw
b1N/xIN8Llk7pYCD759QcDX8xR6aCWMVPBoxD8v1NsD4ycQkcFdyxDmAYkyzivKR
VGBr5W5MmvcjqrtdY/NvDWvdc2kRTWzX6W4LW4jccw9fEAeh0kJhkplDkniVpWtL
oqduy8YJHF6QxjPd/BNWM4q5J025thZR5mxk8xucQ91Jqg3O5E7+GlLyMUdVusi8
/SEys+JzprGFFOIvzf00fjJKgmuwbWb2U7Lc57cwuTGPRpIqtMnHOo6PnfRfRsgl
U9j+s9Kq0TNOYxHA/tVOpjlp49oFwb2pVj1lQF6vTY/ygWcqc1kv5gSoveRufvc0
h/UGtGdqGZC3QeEql0Y6RsesLwxxQunlqnyq+SsJd7CJs01Pj3nDS6Kq1DJDZDf/
Yu8gSw4P6Vmb3WzgYd7L9Hy6w7CPKOYbwlEPxoGVD80ZOPqSV4+3rKlDvXpJEBt8
KAXnoI+egdgc+9vqouLbtO8THAiAkDSyW3vgMINPqqVE19S5dxD3Bq8dzEPEdm9N
DnntXi0rmp7THSIkhPLr5E4knuUi94j+mcAJDeg35ripe1xLJqmzOlQIbuhFTsDY
mWm4Xk7Es6EK0EIyVsF4tYMx2cANWspXN0oZFSlisNmOAXBiKYEdOjQjjIPESHi0
gQUYEoIfXFA+kCp6/cBQ0orSm9fjqKsgRDkawxDn5FJ8AjnrqH2URu5vBbwlX/fk
9RknuqaY8jxBan01MtDIDto37lm6sTY3SEfqMpwpN7Q+Ph/8V+vwOVOK1FHgNm5Z
dUn0z9gT2DOm4EAD0wS9PLneI+2LXq/D0HKjzfgIkcpmslnkYLR5iNWVJrONtyFW
1QR2zB8FdVOm2aFnhoiQ+U/QkLMeRN9mbwmsNG1a1F4jwXVw1oxmjgW8WIDESlmC
bE+eWR7wvfewEdteZBK2qtpUOaLnkwHtFfFefHgDgs0cdJhNr9cuLep1DswbFABO
zS+BI8o7kSWMSgvDHHTH2agc8EVB9BsDsJ1KrcMjQXEnLiTJn2o6ngyYqzbmMQNK
7ypfoAvdU8YUvgMMfD2+zZ7gWA/Cn3lg3b85K8l6W/SLlnqWJNPj+q/z9j60A6y6
JHmd3drgINCO2YJUM39EtEbpZ/vgQ3VeIGJjK+HRPJs8tbwL7fdmlaxGH0NEwEjR
jiKnbj4gnhYznCh4f6yEPCg+2sEdKiwJxTESkICflBIYHOidPe2r2VxqPNNXgSdb
cs6a46cj1Xwf0HE/AIfG0Cp4rrakx7bhdQqfGW698sfjiMmjfAh4AjKvq5O/6BVs
VDi8LywF1FmV5P+lXNeCCr8boZ6AtNKp6Y5VqL3mDlqU0oerFeTFDgFKcM9TB2Xk
IEn8HYFkDBypmBHAuXfGKVdYnP6Yj0IoSyYFNmFg7ovdwavZnvclo0BR/2wB/ive
IIwiZ7T69Iv89Ld6qlnJVflztfjHCdbj8acJfOS1JOpH/rms/XNAFdCKaMiuJKe6
YJ4+mz+nuJJ0tMIV7xfxxq4eE2dRVPOYaay8CoZE6hk2RM/7NQqFs8tcsPNoFctg
00AG7Po9NXRou72/JEHINfyxX3/9ZwOpHCmHwoAlH3fbLzyv1YFM55rHoIWJj1dd
HOrNYLfF36gPGORnU1cw1wgVZE07+VlLdsAYHoT07frpPGUarxTPGslx4x8ZquXS
RW8oalukcNDvBXlFs6DXI9i+OSiUGwNYhrJTijtxG0Pg7rlJY6eoQItyvIUR/I9t
YOiHvfZtMKAHJRU+ByZFNA5ITclrus6fh5k90paEm3wAk6RuSQ0I5UVLLWbAeSgD
ilPyLsavL4amz8reMufrpIjPq0cdb3u6bwFmTjf4ixFGet7j8BPSlZYPienhyI1r
qCjRlaCbwVX31EJEEHeiOrKI4b0tyDeptTn6EJEM/7OkMCOS6ZmSufv2vfh8SUFu
FhVGviHAhzj0tkfcjWLrBOuPTKbH0NUo0x3vYfVXTBrDaY29HYbA9wa5VTZ+Avs1
wQ8j5I6vLd1oDXvP/5NIR09eBbatJ9POhv4hh4tQK6PLnlKTFq4rwD3Cd674FP/e
ywpHyUHovAGpNMygIGr2GC9toPyGHOIsDEOSt4fKJpLESsG7PftKoc+b70qKJ29g
y9jld+kmozylDjSWjLkVqRYSlxipsUd2MiIuZpLDdYWu5avo+W9xYkYLSLW7E01N
OjROk28kH3FLCCANcBRs0FfN0v3Un6v0/cLOzt4moWMlH2B+BZOW5WIziKv5JUo2
1/Ui5PwquWHr8/wJLO9gHB+TqjFf1HTrDhtdM+sc3G9/ypQU03j5T05E+DBi952O
ME1rtH0+SPnQPwjJEyS2a/3Dz20buY0N5hoVDaSwqCIMSlG3wtKzxEWj7ugogDN1
qkgsXMRkJKIKfFVbT3SHWKv4c2jbWpRtF+8j8Mc26FOmW01THEyV7G8vfyYupqdz
S6Z4LOdolJOCTXM+UcMxFMt+sjVZYbt63jFXa6BtNNoUJOIHSE4GyZ7Gfh7n20g/
2jutQgQS/GwqQSYhFhDkufl/ch+hw+kDgmqq/OjuQN6GqmlUM+gco8VhTnHhMewz
xbmwN5JRLXB4YtdMN3I4v83DkfPubk4gbJrrbJ1CYNKp2RTz2lyVXLa3Cr7bA9y0
xOTAEQ4mHJt8JfqB7tuuE2nVmJEUettl3LRSHGu2zu1z3SPGPqi9lTrVAHo5iuOb
QHxE3IoJM1en30NmMTdHpBbE/POIy9JDx1pKrx9xd2le6uXygn9P3N/MECobG64Y
Dza5hAgMZavHtID3W8NbbJWrNIBZChcFwfAwT2um4RNm1B6bSuwLMCb8GXuJYJPi
lRucZMNyUrIRQBXZhGnawMkzT7YbJqDjGrlEqNvEBt3h9M245mn/sisjVGi+RR+E
Zx5awNpK59uQCt/+MO7CAlGwmoSVun93I4luNt9guPIJw8dnJYt3cfcMPEfFg+OD
kAfIECFy6Vq/OUq5gLpvD5mwcK0QkACXXS/SmyyW3c3qwe1dyekJnog0YYN2vMmv
Ksc0j/5Q+NyOgaVhcYrZPJcCkI678GQbNvMgmlH4+BxTXqBm3J+vOV4f9nLlulOw
4elSa6C2L1nMacIIE6QxwH6lCGu76SlpTpVl+sJoZX9ubbSCIPv122DyLj1vSCNb
0e/GilzE2gpoHBtH9CmsDuMyxt1AINir4T0A+PhzW8sUZq8ZYWUTtkdKDOuYamVe
A1H+nUPGUcqmkv+aR5eVG53ahEzUAwrNN6FGuFAiFrddMmKdW7xYDrkgxuLsHteR
mYq3bXKIdzJ4UQkDVblN4rPeazCJirQQrjOAebx/UO1GoNubIp+E9j3DDu94Id6s
mezkH3UxrVeRojbglrU+NR9/laUXOoS2jXQ79CX7LufcGeJwD3kjXkL0Ih6vK/fb
pbJ6FHGSukE3mG+jQLKGeSWRroPD0GMyzeNd9L6cH/OnlgR62hMHAEbFzlwh0p4C
OuEb8/7ZBOQ8Bs7RzZaUfrcfdSYkzHt1HkdIKn3r3uouuisu+ko+0cIJXnYiXnxc
gyGN4MEQvwz7LbxYL778V0YMExpUJCnEt60QnPAM6XaiEj8ea2tDts1yCpuQbv5x
l3UaB2xx5c0RrHs1L+UrBCnTbdoAl+dW+0r4je1L7YFJxiLAfA8dOB0gE94OsI2P
CYLXcNI6IsVOQf8qv4ibhS/bmeGqhxEVnp6QamloI2nfb9eWX1aNZj7Bl0Jnz38+
lIZapVrP3PHvOZ6UpM30dzpwOwbD4jgBg0pcn43OFRTsLsieQYFxhAc6Xx+7JDYm
HtJLRSW0PkYxjXz/TBXBoQaNeD6Do8WrhlS3HkVaVCfHAGFCB+vu7pt7c9KMqvnP
81bAIIyzJmqTL9rW6sIJ1liilBMIq9mAK7vXNpW9Hb4bH6Aycvcud8ER7FgguLJ3
3MPgLCS+NcPCnzLwVYLh8DMRWJ9FdT3HByizWXAka6xOkPMdIzm6S/ADSXHKrWRf
bYOJhwApQk2tgSyE9F3xCYAcSLRD9KUebQcdIRf6/nqzwlHzdYIwg/+2fmHOUnUG
Ol9k7WYzHeih40+11RvHwVTtmYXJV3WaZEXXJk52zmxXbTBproYLaMayCB5SSJ6W
EP9W4TnVmIukL+FOBkPhNAST5AoNj9T4MKSCuNzq4LBi4WRFYKXS/QnlF0L1ed1E
Txuf3onM4SaqFPIieXSm+UFbBMF/S1KeOwQixCHSGCd5By6v2Oktj0nJZ5tMVikI
SlO3Cd+Fm+2MnnkSN5ceuNrEIzOf3tSvTlqhBY6j0JP+u19y/0XLhLTOD8KBCzJL
CgMwFjiO39D+eEVakYYoz7F9vG1ailIbE0NQZDkU+lv2NRQWtbIM0vx+NYjDEOUx
qRkJ25xsh9cW3KZF0WVt38JHv5EHGVQN/7Y/cNwNVwUmyucH3U8HWYQ69/ITPv7E
NVlJt4Ct3lEJbKYwoenXmwVqxpV+qu+3y9lYhIjTxIMgmVJms6z5XuPyXVnIhsSI
cc/hf3UkeIqsdO+LhIgGTORJ9729kiCTQwziZJ6l8OKu0hL6glenrlQERFa1D+XT
tty51z/mS+n1N9hdpGejze4kQSmtP1h0hJaqTDLml+Hdk0IDe2d4qdUgUKH5wVCK
UwjuIs6d+cLV23QSwRiburH5Qhk0tnc/a7bpblrPziS9NSQQuC/PfhaZN+gJrEmQ
BQed/9ddjy+N+7JHtwo2WwuXlIOfHSu7eKPvGGw6/4Bhn9TvjmAFgkyiZ7nHkBne
vXFjDe7LKqKrrMYBoS9kYRHeCzHLYy0sZ5P5QMwk2wKkRVkel5bc2vQAJeiaRYhl
AWgKi9DC+X4CDde0DRm7zNRw8uei5FFhB4UzIdw69P4HlycUGsJ7lkDAELQiNuS9
j928CDwhNESs4uAOjQDIqrYmot4CAsNb796E9T0MmUvcvvUR0Snj6/vdiU5r9fUT
LighzpOmsGb17+IGGczNGdRheDm72borbFmrvd8TKannRTDU9Jz7NPcXSPBpm4j4
aX1gb4mFBEAde1xS0q3izD9LEl5IIBsjfNRWH6QCqYox3vv1+W849RKCjkB3sNJj
Wuo9R+VZs/Pjwz+5ju8lfcgKY/FJ1l9H6APefwemOd0Wb33SNV6f+TLfdlO0yF+A
4qNkqXn2z+WIRAN2vd57FvQyvMsfB9EzQC5HgEVQTQOZ8zNniVj3PUfuk8vGa1bz
nVim8PSlbtG1PgOCBrSaULpLzAoAx4kQGefuWV85tMCQE10SwSAsmyyhDGpzYWhu
HsH34y2tbvAvR357mJLl49oiTpbNMLnlYgTm2yvfi0Hz+FeRpiMNpklm1HXJCQmc
DDltBNHt9ZFYZXWpchgwiRr8C79b7aLEHuIlR6LPOwqlSMZrFBn/S+koGKmb5UO0
sFnS+b/05Pn3yKYHkow1RshcoJe26K/xpH5mnM8a7C3FRwAVjnV3LM9ZF7PkMLxu
9KNTCmHOw9WkV2IxR27Q2apFowhsqE6b1D0ewBE2whdNIg01uvoa6YshgGiD/d00
JAVJIhCGKb8LY5Id75zTrBbFX6bbyVpwrd8JtJ5GZeU9kEypFUHziEhtE2Y7N/La
knBO2jmTQaiJ6vsqVXYFpEa029N3wPwZNIYtuC/IsWt/C978zo3yJf6jOaPESZZ/
o6DCAdc+Qs6uMFTZttOTXZxvGvcr24U0Vn5WDjHfXzmyUsttbti6hwdJkKgA1mJc
DdAs6tAib04+d4Kw43kRz4iIQiwfZbssJUMBn6lW8SNGZU+9zbDUlE+I3NK12gD+
HXfViGkC9rh3tNLNcBN0iUF+P0kq0sAKXNSaGJt9Myt5FWGpniR9jLMtKMIi0y6F
rrA1OYHjmZSFU/P5+GJNHbv58FRudCj+punX5IXRwIbEv/vUSN6qr0Bxcn7cTsBx
yqdo1M2b69SJ+1SgB30iUUndbPh8lxSwzN5iwhmPWlmNUA5MJ8I0gQuYYkujtWVR
JoYv4wVeCW53etPyMvvNRFRS5NhfkHAUjYidZe25xr2H2cl7O1A34OqWz1KIRTp+
iHh6PqJvU/MQRERfbaljdlKyHzHZIHnrdwlqJlnC/e66j+wBaYq2c3U0GHvjuDj6
DU51GT6ppQNS7Ex0GVDfpWBaOYILs3bB7Une3pceNguaSK5i+u+oiBIXNJuQlj1l
BCS25MowQTbX5pXsbTb/Cu+b/AD3c/flMThBDH3A8zH20XSeT2RgVV7xwXNDW4KR
qBRODY/7Mm+/rHan6Bw7snpA54UcUk70X/QWEQ8wcGxRymbkP7d9/jiTrPo4OyuI
1d67QRWxgAaJOfsroKSNMf71SK+UVe/1NhlIucC5RWcvcUe9jAM7KdDJ6I2+XIWS
eLZKux56A0FRKfwGCYX7SvCEi4RX9VxQOKP6wH+NhkhMgoVsalTZAy3korAbLMgv
oMIeXXAnobMmlykbOQ6MEBQ8w6fwWETqudztk1AUCvzhx8DuxBQabeXJMWt69tiW
wK3mvKV0P7k4fyCA9P/QZNE6Bol1i9CZ9wtXGOc+F+vyCul7bdbwLMHYw4G3102P
+5wwko9KxxE5w8ty3zfY4tmBZRUZ33QdyT0cxgYME8HbwxQvICXLX0QKBrShOeY2
vrqHAoZuHd1t8uJx69yHVSq/Mk3y04DKHolni8Rm1lBRx4791Q0q31mEZ/z79a0m
R2LivVXwGCV7a5jcynbDtGuc71fAathgVtxRUFprOa4IgJVnqZ5MsCxY+FaprL1J
mxOcVbYC6jyOQeVtS9bejkA+uoPm47cCIJ+bMRGXFa+CCs0QD2c++8ifqNzWa/tD
bsxoR4iP0UWHYzM1V8DiAeYOnveXtYy5Nvaa5h8iWubmcasTqjGpu98h7yzRNRia
V9aw8um6DqN4DOpIfGZtZn0LhtLBaudvT8SGGCLH9UiNd3lM9GiWlDmBi+s55V/s
S+9UIpkUXSDKdERJSErUlseVYtpQzzGa7Ko11ij+sDKKfepF80AIVabAC4mzgRZ1
UTI39CBdEL9GmhQakCj8RmN8i5JNyxO2rhC4UagyX87QL2W+pmMmXrNZrTcPD1yZ
F15a6GwvfTlOYUV3ZGR5RBttnN/Ter49G43tAZBQ4h8oT3gG9CXD3MYVrxZLVgna
jukHT9Jnj9fDj7DKM5+GnR0QvPZ1vQYYOt75+/x3AASKKIpMHEt8HUj/TG9xmz57
5KpjbIcCyX7ZJeJ5rRMlOlrKRBuX9+phR8tmvjIsVPP8TV5JRoh3O1UyUkwbXeJm
bnz1hlyujaowZe9gV7/BW/NZOBMyY+/HAT7ndF4h25ZpbauuXnmx6x6YAhAS9ItM
BllZ5Cxpi683ujWW+i1O6UfSO3KC65unVeeFr9cRenHr/5B03wkwmPyfESKRXlzu
n/KBc8vljbxIX88R7GGMCX4Sb/sUeZF1mDvtOadK2T6WcSXzK2UOLV3mpY/9TRrr
ZwZAkJrLSDtS306v5mkxz1GTkmnRPVyWt/uEMWAFJballjEzNR0JEFOx41i0H29W
PWy2AIj2N90tRnJdAxExSFaxqsxOsazkZ4HBz4k0I3iCXhLe5pGyk/UxMeNrxCGW
WWEoLc7Im488SkAZFQxHkvy2GDNeV/3ieympKYewR/qEB6gu5laXPjxcruA0ThRU
GKT9Z0CKpIubQyDClmtmU9T+Kx0tLinmbVQEkEGXCAX6Sb+DgAzXtLugYP+Ylj7o
kviENbSG3QQwa9JxbzGYFZTaBiUu+fLaPjxbDjQoCy/ZJghX9VWmxGifkTrDL/k4
dXjT091ntmwsv32DCVdnncZ3+S89mBffX43F0jnMDbsTaZiU7QarrgqkVUXqOj4K
SF/xi2Q6//w8kl++R8MMCIOiyUbGp9S6qkfxBcgVEM7VFVTWVQrxwOgb5vlYFpo0
+eyCHxrkDbciua8aicVpgJHqZ+6BSTylgA54CYLDh97oj1K2lfrgtUpmbMt2tpwB
uT57BpHjT61g2o1mwo980s9989EGfvSofU+wXS4r/cD3nK7II6k1fyxK+8pPnkae
3hOnPrnPioPQuuqcqv8gm5I/7NTfM4YXFa6Z5P/Yu/GCM3mlZmZW8Rw4SUW65Ze6
FiH3sVSXGkYIxyh4RII1TNijDiqGuzkZr0jmNn5Q60L09TeLsEZue29gXkC4hbdu
c5oUwqko6RGpPQIgKu8dRflOp4K4fTlPvokMuGo1rbjmob/SkfcJEz1XE4yTZ1XE
G18wyA/I3C1RqY+9M+d2tVj7VH+AKO++MrnSvZgUAi+io8hv/WT/0LxtSDSqZMc9
ty1OJdKyGIc03Bfoo+Z/N4kaaej2hVBKZWtdL6//ZkxPLKai18xref54mHA7Yfqx
JOdjRwm31WDO1bSlPeRtzqHhjyF0iisnmro7kFFvZxhpXLsXn9/GxNoetGGMk4Kn
AnVqttPdx1q/Lb3kdar4rTQ44FdDXH6iNr7AWwZID+VFLIbgDWNZonWy5WYdZUOi
wxnx4RZWs0M+r78vjgouBEkBY1QZbgy7JMXOjT6paA9yhQBGlsRCbFJsE4NXr/7U
+xlrP59TkRLrOQsaz3qmYlVgcLHx9KbzcvPhAzrTALJFWGQwc9M4GzyKwQQAnFVq
d1LumXIUE2R6ZlE7NWqr/n7vtTSSe7XXkzmncDvd7/fw8NfgCnVK2kQ0nEM+E0sL
zFX5TV5qJIpS3iw44Of4BYUVB8s0qqkgV5qWLYr4igWF34zPjdpFQIPC9QGgOYyp
x6SWRynEuwMv8d0Rg/7HApEVA5tbnTwpC++GQlEGc9oq59bLZwcugieXcAx9b6Jd
zD632TrROiMkN7bdmInnxxzs7DB8vC6IxXLOWOktUwh70VM9BSPeXP4wdJtOfgYT
z+O77kS79P6PjvH7FvflIjA4tCipKwmMxpnVzvk8tT831t39pQcjpInjU2I0AxTx
mnPhJ2w1cl9UOKhc9VOlKU0cEtK19SHZbmifvlneV69BnO0ejLHEasA2hlR8utdF
W0bHBTBbWMyH/4O/kkwuKNndcyB9+4/Mgdpmg/eYoKmHWj9lelC69iS3uUc7GHap
BTfNA2Ah1UtSZCQ7uz8ZImS052lnhf5N+ZaI9EoUnnhBLKetxIFXm9ZSu5+twkIC
PNTPcWFr3HQ78FNq1oknc+uikh8M75UEwJW0rSo9jYqLLlrW6fCC2r3Tg0PmZ9+z
6XYzoM8IPju22HbgETE6I2o3mmLqRYtn5fs8zrDsRqxVl8me0U8fHy+md0AFRfOB
86Csf6li+STRPb8QELurdtqzo6L6+Fp+I3dVqq+CDBl55CRVRXdFtowLEQOE3bM0
LfZlsr1qP2GzHJnCsn/O5k4lYWxAXpVyJx54ksO3WBAM/cYEHcuZZFjb3ksJYVe6
4r09De/AO/AtJwV/G26WD4Qy1k+qF+TOrMZCZWSHdC5dXyHaYoHmgWYwqcUtbmWg
TLetyTOZLaeHowHTe/CnV7NX2xIQYbjerLwBI/JoHY0KNj3y2hu1w/iXN1ylyYP4
/91ETYAG3cS2Mhv4mSA+gJz1mIDC9Aws/gd+I8MMEQsue0HuxGag0cgentFujpHt
ciI71YinvPRO9k009YnC5D7VXS851RAQomizvexC1HOV5YtfeaLgIZEY4oMSZLGo
P1Bm3B9kSYS3iJjgI6pyQGZR0udUp/RB6lUAVNauS+/ogOfr42Fp+Z52vAMybmqp
cGjcYch+0QlMdJEAO96Vosu1wy82v57Q+yvfLgZsHrUgRm+gdd+LGrtvD64ejOkz
Y26HF79VnpPD5AS3KkSAjgXW5RpIuzA2AiiHRs1p9fU4f+8tTWGaEoL5RYc/84fF
bkZS57j9PM0T0lqu1AWPQjKxJ41kF16CZOke4Pb97lfM2dQidJX0ohF/fevNk0+w
8I/LgJeASSfTH9YRPmhC1xi6kFeMKHjA7d9CeWwomx0+MhADgTfW3HbxRAm7+j5w
LQipHtQQNw1HwUJnkp1HY2loYJr6wcbM7lSDwmd/CLgJmcmI3XZ+Ume2VhqEbIOA
byK5rnAxU7845bi4up0QpAonDm6bOAaTK1X7Wwc82iD0tc6qTG/Im0qXgfGkWCtZ
Qg912vrtd9c87OM5MCUHDe1awJmK5zgEgW1b9yXojGvbk5z1Jhe7ZbLueYHXY9V4
tTR40V9AJyyvhtE6ddUH7B3pnYC4AS6TYsNGoBFzI6szFcLa2a6QGA70YzxVxt+P
NpUJVWKse3dNfZKKeCQ2hbpbWfkV/Lr4rpIIt/nGzr7ZEWicQbyyH1nb+nFonLpt
/nQgWiY4CAn5VyNmHgDZXlZQpNf/lRf+5sOcP2Mw1Wv7IB1OIBQcPx4Rl3PlTx2j
A5npcB6eKLoC0iH36eJmH3a+hd0i81wwuUNf16fEMThgZFqCY6K3IZRIwWG+xFjY
p3uKgMVd0jmPmzXCIisx3SLVkxxtdrXn86pPkdHVJWR3ck2XIDnp/ObtZ43WO4CA
Iv3jhszlmE+u1klAIVvjKn+ccmCegqrtyCmDJO9xzoS6tDfUYkvxFsy0UhKS8nbV
soEL0Aq+CWBUg5GAALrdTh8H3H6UtMNbr6x0BDjP+IfOzGXkG7JZfFf2PpKFqbC+
BtXJyY7fkb5RjJRWR5pnuopccvOZoVapg+j+U+9q/i+YEnzsHctk15D6t3a7htuw
14XvJZizzvsO7vxQ92HkxW6O6j+o1rFAEsh0xUnezZ0GQ4uKuKPnqdnbhbnJ2rmp
DiDzMHH473pDbpytZZ6fGYqELf3fU1Uisrv/GstUrgxbIB8zSV9qnMTAMsr852dr
XNYocSI6aQZ8ofuUx4PxbPBEgUwIBCY7mPz8ABJoCfmcDXnq1tXRyD7OewojvZJu
3i9BXdeF6LlX33DF21y2RMMmb1PJ5O0vROiMgGV+/X+sSD54NOhSyXRoUhxJ5Zan
MEt7stGkJEl1AzCqGPiqLZhtqr4nFr2dlHAdhcTwO0K2/DZo09P+TAaDxxs/lZHE
7ITqug/yeHk1nM20/wzicUYNS95W6T7OaW5LvIJFHJrXyiXHu9soNczgM7sT7q5B
8WlyyChtgpYRshS0T21Xkq2A1/k1ExpZWQvyHJlhVwLlB7A5YeWwOc4K5a21eST1
TRrukvS3jB7PqDkzQm6Il+RPpRXDjEJcyQyVZxSIqCnGEueSgLyOtvBTv3RLrnLv
lHemFGLBqzUf3bb4JSkXXvB8RR5bthVSran1EXzpc9hvA+YMBoNl1Ou8WG4bB0jk
Usq6NWLwMKPBWcbm6i+CBe0hWTHP9b/xVTKFv2RnqHsTSFLXFoV4AEKfeyUDIoi+
8gElHVPgK3cXlNvgumvplzRSYIp4RU4mpUDXCdEJ2vye0/SCLIC5f/b397XnYnOc
5HTh3YIBCuzR1dpRu0ba6PQg4CE95Igd5bdiPPBzO3NxwGds6gaIuqttDKJfmjHM
j8Vyk6yLe4lw+sRpGZMjN8wwe6Wsug1B42Q5vyWXv7E0hTR5B56eLSCZJUKqrvuw
rDtw5CtBDHiooFs0Zs7CgrZSTy9McEZoYoIkRX09eTIxjbCI2NVwDI1xVR/z8PAq
8QaFR1lnUYyIwICBzCt0FvOuc/HQ54/17T5g4rPFKfMuwslHsy90RJzG3BDPaOF4
PgqkWUo/mxIdbhsWEOsBQXijlLB/w5Jo96W1XEYorc0ei9QJkwMLxZaExIv4wQbA
rRuVd29IFVkl6XfTnkKx8htpByzD35JDb8j/BfqCQ5U4a47O+Irj2XNijzkfQIYN
sr3Z55Klgp7+cKHfmXY00JmXZPvZxJOJ66j0u4TDf0AGpWWMJv7QhcQO5hFoBsMW
0StuZe/yHmqUBCYwrC+njjDi07ZQenEppY91JVm0y+EuLh1JnV4x98LdfeeG8zC1
Unlqe7Nq0sx3oUg4cxHan5Pc2/faF51kTsk/x1EYvS4Vu7RsStZk4RAo+2g1KxvQ
dWvCkYTASNzzpiBnoiMwNZIBXAc8+mYlamvuh4foKh4rqKktI1Rf3p1X5dSn9pJz
++Wbp9dPFORv0hzLyl/LqVBxAX/OkEbhJ5OCvvvLK1pxR4PC5uycfYe2ZNiwbLaA
z9bbK2gJdXincdVkvIK3NqjcUa25Y0+Wvd2qBaXJmLSkdE6Ggz0LssRggZId5CPV
z52r9inotN4KVrGYcfSqt1pNbgHB+gHup44WOw3XyulvntZSC0MpoID9xYIxQYep
HfJTDBszE/qmX/OVPdqBdvNf644lx0RHQAAbFZkDDqc+zh5ecKFgeOyJcjBdJHfo
kpJZoKeOL9StSOUfEznCugz68HR0c1yPC+mU1AyhOnqGg1oBp2FtjMYAYY7sNly3
PbH9jIaAKGVgXFsl9f9Tabjk6Hn1DXPJNXS81HWx4HV6hOxkLNxcKY+cW0FcygqT
OsVGyeYc+Aq5BNFStGCVyXyDaKPnaqFSJFx4IuRr9/OLiDlB8N9YYA1LZl4WYKVK
7/Wy8GpO0+AocUbXzvRXX90HwhwOxUjBQH2+WgEWJT7weNsarH9Io6YtdVAXtFjz
az2mXNk8nUeuUuQi9l+lZeK+f0LjFXpNO0g/DEwjEQ7+OBEF2e7yUIj8H8V9rfJg
tIsySc2JfEwAZRv7wEKyRHhWYjJ9KnsJFBs8HN36lqtTIOvBARTMo5N2dq9ddCiT
EMpxFay8+u3QNKaBN8M4xM/Z9PHSTq8BIR4caaJHBU2qASVa5OZLJmNW9h7zjfFa
CQltRh8Wra0OSEJptw4cyrsktGjaeCLUihPTpjOW2XYogLR5LlnaSFJ/XFXM6/8k
PMSH59RKtsoKT0nKiXwoGTxIC5OWrJ3IBo82MK3ZjdUS4GxhAgRaU8BDK2fMxxct
5KRvbGmiiGNKzOiB9tRJe04DgPLTOnKcl+UM62UaXm4Y0j3fxxL3VSaQuVH2+wbq
+SvDCw5OsVaMJeTxQp0pJUZ8LeMlTY3qJHruXTgR+EA/9T0RQ/NDpXQEiHWyPwKe
wQ/Jwwyes3Ubq/KtIWfmd4CyaT25vlHCyD2OgunWyG07vcGWoClvnG9ZxDlcOC8h
vIrYwYQiFmjrPP6C7bI/S8FE8M8UNHn3J+GcpO+6eoNIRJde0zGMJ0nVmpWFpLLF
FlgW4jP7aKOAuKZtoBFLRhJuu/bjgPMYmidjPbE4If2aLJHE2jlRVSt7G8ZJVGKe
Tn0CXFgsNelM9i6SPpdErpFayAKB7LIZslrGW1KRctCz6X1dMYUkdu1TXzKTP/Ax
0ur/qrbm7fV6bu/Qbre1DTsfsnI45yjZKBsJ2qWbnJc5yx4NgjzToTvkPbjzNYK0
o4xVzvHNFOw/DwtAYKiHqVcGHE5aVLUE+gWI8h+f+WFbbk270k6sbd/ufMBzU63F
YUZGNctDSP4q1Ct3CiNLbaOAtRGf9yfllU0b7835mKoFVz3yj9Uz0d6jLXiSTf4O
7CJJyzb81ET/Y7lWHY6rNP3OcOXZRNASGLoa2crcxKjj6eW6zyZXDUuopNiFJ7Fr
ionvUhRH/mh8NzMDFUdKQsH0qbhB6daI13UUQdU2NOkY0f2GBSsxRJzJVV67okOz
SuYctHUkjDwGdSZxo4txihoxF7VSH0QTEakV5t0e9PIjrEo4IrwRJOVgqfAYfGBo
81KPC6OxAkNuoYAhGvrVzSAF+2rG67ETZmQepoVnxPutkQbQLH/Hsi5Jsjvbyvac
MqUxXiKSU4EjdZZMaRh32YiPrT2ZJ4s/PtTCsnr+0WBgtlCm8J/G6gM244b4xH0y
WxisanSyeQtFdfYpX+krUL6NHRDYyUPS20glDr7xcXotIDfI1gHz5Agozq96t//s
8Ilu3mlYMeLvNrAQx5D0wDt0M6l9Hvx6mmLTyzvpMlnBrz2GejHjM74apDFCmBpk
itHQv3n4xcq+RxJXhxmGpzbtxw+XqYZLAJJVKuiu7BRU1kXQW2nn2XW+VdBhxS5y
RVCWXhOP2fL+ISApS/YH4NzNTbv1O3SEkk2Zy1XBPnqLH5Z1ns8p0XAELgZDzw/z
LuRiHTYFbaxr1Xkma+ynm8ix1ZwEaKlpFr+jOMUyLoXhPj5l9KcBEkWpj/tdQaBg
CVabl4f52MfFzM0naBOuUyj8i6gQNd+aoqL/Z0c2L+k9c6mQru+133Af1XQdswDV
QZzpSQq36Myhdg+wg/FuiUIc9ISb+ESXG2hyUp7Pecu0yi5oHYyanZhMHQp4XYO0
5LO5g0toIZ3hrDCDFOQnOXkLM3XWhAFX8d9p4INSJtqVn1hfDdPjlaZi+TH6zMJl
CVBsqnL5o9mgpfmjxTIA0lwwm3UHO7hXiFRoM10UjlIcBiDF4MCXEpqM9wVwWnIA
aNkKId/6LOfo93noiJceoEAytRwEPy8FJsuJo1T1pqy3O7EhSKk1BeCCqaK/439A
dHa9CGWchu/lSspFuJ9AlJBZb1GMpXxpfxOcG4Acqb+8Io7sBV1NGyE/XgdQjC0C
8xHUYM9ZzlRTixtvXThzrKotDdmfQFimNkx7hvXNtOxE8aM1jm80c4WU1nU44KH4
Nu2U5B9pdDim7hNmKaux0P7oZ/oiUY9koQqa618/HcvOGf6r1BzJG5yUaCXvri9T
DZum7lPw2fUiLiF2CZRT3qhUDdieI8e6lJDvSR56vEbOWxzuQ0GhAk6OoCbDkBxR
VUVmSJo30Zn2x+pbvgYFwXGiCSGonhwX+T5PEmztvHdLLZegYlill8GItnD+J6d3
IczJh5Xfm4b6rXEI9mGRyK+kXX3YeLyHYYncqglulJuFFsLK/rQqi1QD0W/AuzkW
Y23IPo5dJ0y8BaWjtljADWDg2V+hdPNeRbXTfmwJ13rSYjxZdV9+8fIDv621yUok
i+rDW0x9Lo5dBmB3eLfqfhfhq+V2UHb6upKTjSWNSDEjj9H/UxMhM69T13tiFLmD
2jcpGzJ2KeS/JRkd/sgdzghuDjgzOcC9Hck3S7b/tcLeqM3qNBRYC+pTw0EVMZ+q
z0FKxmAXFUPNZwQFgXKebFld+5lyUPBIFHE3UBuIp2AWhla1WDxAe++fRMZyQgxo
zbUjQvI8T3lR6HdMFtL8v2FyKkrG7z+UHOmz94c/bQoZ4SYkYff3QAv5d6hD1Oa0
UdIWSh8kp0BxH/rXE9OfaO9IouANmYd0maGumHE2rXgJgEJx/HAyhzZiajXMFmUd
OeKMYm3Bnih3lb5GnNu0TnXmtTOoLSx/qD1oH2AS+snfsbwGe+x8v5Dnyop8bt9v
/FcHiY6qnEJ7ygeV0y9l4Dynn5bN5LnzuFQAiLoZYYX6etRQN2+EhVY0NkDLdpwK
WUALI2XtudAXUGHceprhFAU0tNATBeOSsPWeP71DGPSnMlkJ4bDauGTCk5Frt8VA
h9IjqEj+VwUjINhPbV9sMmAYabqhifnG1OgHsXx8dtop82bAAqJ5apKNNSQGh71g
tHDy+2IDczOj6U8zGUITw6lh8FHZB28A/Z1vtuQVuyZslZzaNnSRwOZ9MxX94fdv
GXddDxQ+3Pwj6d1ZC1KGtTUe29A5uPbSi2US5+sx7i69RkOTUOC73zOK6ms6bonS
j7Nh8B18ePQRMCMCenr+FWgE3koO+RpLK+bYNFOgp+KhpGSyUerUKxBAk7IVL5QX
ZuIqs+51qZ6kS2Xb3osYeMyYcVk3xRzndsRlQFV4Klo6Wt4s9S8Ex0vzpHgN3AJ6
11stogigQFJZ9n3rGwsY3/u9Z1F7mVvf8w4KeE4VssYLYO7DHBm6mLYFmjEka2ij
Jgr+NQT86ZkYsEApBhf0tK6Zg7T7vqCy/KCe0AVZL7xzf9wZjRKXOEKZ9i2L/xG4
AvFTcD8vSnIoh/F+ldzUG7sybM7g5DGFSXrACTihBQLQiQWs6YKiJ2cOath+3qZs
KWhmTncu4AFAYA7NzVQwbhkDxAJ7/JyHySTfoZJ0szNSNHrS0Q3e1jCq2q+gX36k
3Bu2/4rFmhXJPQ0u4pJ4SHRwocHu/qw82lO5Vo3gMyYbpgsdoZkZTVbdgWDFOT8Q
zwt+XjcHNC1APPdnNxGsu0R7TIbCanwPtmZOp3t3ojhugQCKrl0z0MAliibC6sab
dgoxdjZ+W8S8ll4TRJFHFYMZ04ynA36pbdPhiooW9qjTJqPiSErFWFcAs9iv9+MG
fvPOA6htNx3ixZHWhue0a0D6lMwPHpq3ALhovV+WMT3N8uOnCtJh0IqsQDCMaJ2D
Pe4eUuC5utt0lzHK5St3KV7Y4bTeAb41xYJubOLLvQt67zokXvnr0AtfQm0lky2V
iu3D30UwjQpTamRfaz1CS0tkgclJYcHJc1FANg8Fzp3zWJmip31+quP6Srm93FSF
L2t5uNiwULiIpcZgqtpdiQbnbRANiaIR0dFWVyrY1l4aD8CCSdtpoKj4cxLvZ8tn
yjQ5weiXw1T1ejIzGMishcZGHN3RJidL3p+CKsSzJ9viTuzQoIehbRatHW0lJIJl
eUU5SLe0fC5PDf95MUySVH+JbHvmAejiYH/QRftjczCbz6LnvIPOieag6p7r3xDj
I+8Vy3SIlLp8e5TGoEr2i51HyDo3e7rGPbdB7g862/+G6toZWbmA9Wat924vxgiM
OnzivjAApBjMhjCjJqNujJcobzfMTasFp3dUzz3jR5Qj9Duqpc4NGBcM5oG1AVY5
dWjRFS17Omod1pLEp3kDgXkcHbxTLg3oFGJnB93bLGk7GbYuFZh3lS7kWe8mOp6p
43MVquxpiWClwQwoW4GofF5g3aWDqrb32HJPJOA2wYeMjcv5PmvnLhu4MVFESX/3
VRnUxFB1ndcT+tzkbCBKa+8Ofh7kGpcuJHibks04H1/3rNxoqUGWECoYrV4nRtWt
WWqi3J01yf32l+AKzx3tZWQRv1lcKJk9gtr6wSVbhmN1LWCZK61ZSzawyozD+Iir
Av7ySCkfNXSYmRajh27/PjMKbYzgbCePR96SsaaUhoF4KGf24KvyNpHTYN/KbzYW
3Uj/SyBjpcYZuxnYiV5Em94UggXkXLEbOWKzrdlnniNbgsUmfuysYJ7ILJ5Yq7fH
4ogduOpYhSNpisS0G9jG1htzVmDWH797Zf2/HBmq50kcsdmir7XBADKkZu6PK/CP
Oqqg8IM2xtzotP3xDSY5rUWxB1hUQtPTVKMjvok5ifP0/QHXJloco8Ammxpme2VC
bwRa7eMsUM4TEzJN5NLK9un9dHufGslW8dHdzxKiHcFAskut5LjE1crLiMaKDm1V
hqPaOXoHpKPaz7xTc2BTd85E3X4In6qwUkE53dDTURBQJAIqxI62TA9JszKbXFQ4
ZQ1jMVjMYbV8l9AhrBlZk41FCln2AOTH1WamsdflLFjBsuhorP1tWWUTPx4IVohN
Z04RxjWX6DsKC7oE8Ltwyx9I8c9PVo0vCjq3bTePTw4FuQBv3W+Xck5dTH5gLsRR
hqAqgAKXpmsIEKX/92KkcQY2dCgGiqd6rQijzEetNp7Xcx8G7kQ7wh5C/zqRB5j5
pXgGUof9qefHlaxeFbH7RfMWPRrToB8knAbBRW1r5JMrgbv2hfyOE6D5cx40uwe7
UybgDh6vHBMbgUmFc+I7XZEFWuzDHaRNiPHOM8l4C14Oh9p3ZsAVh/jmm+AAzeCj
YqBuyf4qdcLO66oc/TdiWPZe0jYRSowT2L1+cZRnTtHjpD+wgsBAzcXqwuUW2K1s
3RI9XfFqE94NvurAgQFpsrsrMJ9L71hEON3qZJHoNAlAbveY0+1dDEhKRgdxSV7Q
w6qKNnvfnTVAk+TQ055hbWxstRp2i82q/Pmt8p9KARrzd7Hqa/jWAhYDkL7eZrdT
NVSKItjkC6G0NUym8TfNh+v9xyaF5dxahboaO3GH2NWKBXSa7U0UDnj4h2f5vMk8
y0WJwGuzZOo9LgkiDtHCIHAwqVLnGzB6kJV9tFRzkZpTeyakn4+PpE3HL93/uI4f
LAMo17U/ABkDz+hwUpbu5WzFPqxbiiR1Sf6gDBS9ULaBhOQkZGwaSGUPQPM1TtwG
EoSjgIMiSDSWUj9WrplAjy7VT45ISmHAlI6R2dniI0T87W4UiNJ+L90m0K2QRl+0
4BV18VTKSANshq5DH42ZfsxxSEgjzqO/WY/mrgi1vyQ1qftl27x+qDDW4aySlKtH
XlQTsdMS92IRsolC0/yRf/G7g4XEsM/I2HBn9jmXqQKT+W4gkk9GCauFVyowtahh
fcTKg4BbHj2AarDc1cuMEIRgHX80kWLL3+Hb1YqaZtYZA3mPfgbXQTfvmfS4/A9B
8q8VL9j4soHnwgStw/BX16eN8tWqDnLa3PtF3m5oGJ4pF3PyVM8J2J3sxz5B7EUD
a9RC8Dn4ivutCNIr9v50Yrhi+XiY+SXoo2aDpvrkwNe8vekay+1w6P1mjaapdGG7
/AOxU280bCwNSmjM7OU52VEkTcvwbwf6yJuADAT+sVtJI+EUAHVImpEuVP+PHy9b
6e76UNSu2b9mdyQr/vVgVifiq/M85R6Kxde40cPNcFakRrkRtRtgDCFJxuVNhAwH
sq1BBqJDxN2kEYIwzayOmGtB+A6cWLnrcQTFw/ygoPxtAsjtCftOkOmaFVshFrVn
I63BHkEyWBVq12hFy9Rx1JFMJZ0ot0iww7sSY11BWWcOXp7J7sC/xZqSbwpb3Agc
MmA0YIT2Dn465e9UxGP6Bo1zkGbkBN/Gv7gVe0rqO1uFpYvVW4dU83EG1rLDRNRn
INEO7rcKMBDlX1zVQL/o7i0kazZj8h3ulBbT7eoEXN4/pdy1HlPGPAu3jEoWviDm
ao1FR2rJhHcMZS+gR1oqainwJsVqz59ktHk/5Cq1wVRiw5pAOxd+s59BZoxfOhom
cqH904z5g4BiiVeGh0m5FPgn3OWYMjXpDcEU7G0oivnoLTboiDMOTTRatrZ8It3s
Y1lM8GGiZMMBeCZzFhd/agtzV68njtvWqEYPyFzyxz42bndWZFMaFI/OIrThGrNH
aMq5/SyUB8oFEZ42GuAv4mi0EsmMAR1a4iMMoGEJehxJBmqzoEbdKj0KtcbgdkAT
evbgwfBj+WvhT7grTWbsCrI5f4f1ySSEa1XgsYPdrXXt76ZWl/LQRRWfJWXy2buN
uv0MRL7DeS9ZBkIY43AUTCXByheDhB4BywOurcOi5tRk1yScPwdYu32J37R5uuYz
HKSlXpaOAhQby7H6xMtQ5K9rx/YS+9k8MAPfUQKiK/7rg/v3VZxQj/vIaGgJWrzi
/PAk1iGotiqWgv+sNNNPoy46M5J84GtG94jF+8pqfYAs6zEpQbhOLo/Uqts/zMO7
sq3s99kQLTtaoGjVLsspY8ejSR6WxE/yFvC0EaV4IeRoheOMzORgBU9AtUA3AXj1
k4zWO8Mf+EFikyhvTLZ8XotHlKgJzOjgUo2M5ny+NWpsfx3qLxZWGGu6bn/jJplP
4L6V4rpEDcVebZK340BmXitbvPoNUfA0NxxfX3UG3hwIKhjcPdQo5TSx2DiB4Oj8
nyg7ZdaV1i6WmfjouKULMHoaqzjViL9A/YsAX65GkJWpvfVsOQcHK8oNX2h780q8
Hl/lDgS4vZkVOZ2KfxDYHxfaB+5+/QV7LfbdPplFaxZa3FsyZJVJkCTbhuuy41G2
IYr9jxN8xQ+YqJ+OX1yprya7oonRHb0S/11VW4768cXLPP4DhgiAf7qrjqm15Lvh
B+Z352e+VYl9bAF2LWbvvFkmFFmuLPUYtSYQleFB8PCsM0i/KRraRsGFNolid97j
AeSV4Hkn/EjxBY5VZ2huLaMbnvxBsE/q8upSSc8shX6drZU8qU5huwzkPTBx8c0e
EBot003WLmFRFst2oxViwxWchuoHAa0qw8593GwfJTn8GR9OJ50CxL8txwMmAMu3
OD8NFN+Rdn5O8IEhMGyxQ4/b3cN+BmiIKxzMcra61U1Q+lbHPggDI9wkuWwfXYkT
qdn7gO+X08kszE8aJCbTid7SOz8kXi3uVTpWbUNZQMcpUWkS5wnM1fN8Njr3kLG2
gS9zEE8EwIJtSQd5HYoG5jkcBQ7kCcSrzGp8yfG+WZhUjq8nsJGbTsfkZig0Sxml
yPneuef+zPTd7s+pN9XwhTbP94Rzk7wfpnmvdTpZNPTW9lkex7iS9mwNOpVnhUQI
dcxjSO1wTcK7RwTyWpLZ4vBLVYgsA1evCzXUpLjUCx+luBT/fSzuxb2MSywHO61L
tqhT6UQz8w8n6HABcwdJAMYulJM5nyOYqiyhCqDoUovQniTbbBLiajeE5NpQLlez
WZqTPdiZt0RNGwknlifpjeIeMkLRSXlIzGcim1XFbGhhGc96VnMuI/oEXPnT3CnQ
ZHg1ekIPvNNlx0zgn63m8lRSehmxgTUUyc+S9Z6PuD0n7oU0OAwQ1SzKbG+2x/wa
xbbP+RSh7GMXxWFfHRJiIOkKTdv90xyGhMSsofUqhLPpAOJ1FsKgqIWD8gwSk9LC
MGgJPRRY53klgRzuhbLKc30ao31FUMuzQB63k5mF0HKRIqNAguNdok6Ies8KJnZU
ydz29mAn/JxcfRE2r226eltqJmoRbA8kjMFaSBQG8tTjgu5iF1SuRfkZRBKYrJ7+
Pd+Ymhy1z0iCaTGqTkFbKiuU8Q0eWJ2S8jGFA4DU8FOnBSWKDxWD71IEvbchW4Lx
cEqU70Kkm8JCWEsO1oA6NL5K3uKW+h03bUnKBfrKlvUWxxD7hTIz8XDiOl2R6+0w
uiZpPg5x5J3CIvWkDRL5qArRZwqb/SRObiHScvyUAwePy45PAIDux9dUiI3RyIqm
S+36+PhrGw3q1zUOJ4cPA0RXiRG+Tzi3ut13T9o16taqZXMlipXeFOqK4uAUx8vv
zINaQqDn4hAyA4O5QxcveH+vh+9QGxG+85CVcoMmS7Jo/rUMhswKhyXCL0oGSFuI
+rJu5xCfDMPgB0YOlWcbIPbfAnSuVNiSBHSHbSJvyCfRp/i/ddC4ZPAlJAK6+Mk3
eWdAv4m0/nj2De+jo/QL6zmgZkQjmHeOPC2qUw3DWB1YOgaDKSFEd4le/WRCI9LM
bE0beeSFKF5ik82jssS4QRK0KqqIOiDc5XG6YKLgt8KWu5Yp7AWpUmn1MBje7XGs
Eor2nkTqI5WrJJ6vWnT6WuHUy4cdiGOZxrhu+k2ULWmSfQ9usWKqu0k40cjHADBN
R2EnGdvrXwu0hZqtSQSZVAnqM8qEOPjFntHe8WeQ2prY9YGaBD7qLQKDZ1uMWtKt
qpECjkkVuNbQfiEorP6x8mRuN0jCg0DBiyDe2mYZTq23snzmSlruMqIymBEhzdLM
p2AIrZ1NeHZO9YggpKt0jYvU7Vhg+wViJZHyI2S8t8g5Nzqc2huEogMUUctKG5W1
XNbzkYtHni74C8lk6dFZC9E7sXoFzygsfEGDIYGWQv2yFXfWG7o6ECl/rmGQZEvD
sFKitI1x20zYI7RG6Smz8m97TDkVpUCQwbtqsLhOof+9MRZOR50U3LNfTZcu9Gu9
0HTFZcJZn7T1Y+rgXHzSjkJz1MqO3rHY+aX2fuTapco9Q1VfYYeF2SKGdjsr3qI+
Y+eG3RLHGm82ZS4xHfmSOtwwvbtPwfFtwvK6kLk5fUBujrEkWt1DdnjgL8ZVWc4K
FSH4HU2S18o+OrShRwShHbP+dSPXUln6s9aAmRArTRo3EXFgQ4rRiFrQv/H54TRx
fraIJINN88BkliwqeriSeZxOjaJ1L5GMuqDDKOjVYPZGDshY7xwdukQjsvwsnLdQ
+sepRAkkkahvKu5jd8j3h7xHEnizSLx89oU26FV4A8GM18Orl9VaX8NoLXaf0JpI
Ka4uAytPHmsOHOxMIjEkzwAmO7FDPKiaRaMKUQlnV8Ohf0knEvWf45aY+ItXP/rP
Dp6xJB2NRvBO0zRingSpyCszyZTM62/UwqtIRfszVAslzU5rIkZPLRVFWbGCO3xF
TRd6i8pqi7rhNDFSI1TA27GTP/f2UdFHcldIHfXE+gM7cvcjFFL6Yo3n0dV3mtdN
DDZm7wgQzR9KL+9wI8Z+3sJ970FlZ7PrfNj0TN1swx7Qlza7rfIQVMpXZLrzZB2w
+RgRcUKO3KFJ2NaJkwRvIiz9KGGFOdyrZ8CFrb9Dn0vuDyKjcIcsVh2iHutHZ6iv
Jg1FhuSISkwhzvIYK7YPZJiwZhfQowfMScjQmLds5W2IFPyoAInXWFFkskCYC5qE
lbVNlSYTlqutG6rO/45VKKz3xq8AmCTizi2z3IuZaEGYqhYD+bK4O8KIhBKJO64Q
ph+/lXV2pwt2S2nL1atk1fdddMH2dS0SHbFXuqQNXbKcO6x0/5aToqN5hlKvMPg1
uDO8hmGbkIq51dGOfkBK22HOD9FCRLi4ZapiE+LWC1Lqdl/OnPTwhBKb2LXKiBJY
sErk10HiO1+fviwDB7dhHjPH5N90QD+dKXbxgpsRU9lsxOrmvuX+qOV93b9WTB5j
lxQfPTDb+p2eWa8lBG3lyiUzuB8hezjENodMRuTqRGCjREDjfbYn0UwybuurwsYv
lOTGvmpXC7DjuvRfJ06JJWQUp+C2jwaDLxacOpYwHABuao46bO1Crr4r/6ORvctS
fOMaYetz5rY+Ls6q59iDQ5umbuma6Lc8R2W/yw3bRYwQEWr5r51kWzLBTFn2abtQ
o6dZDFY+47bzVh6RY226lkdRsRN8A0q915lQzAWf5b+x+3IzL9N0eR0ZjgfVgb+a
5LS/0AzgnLjozX/oBjIHnULRxrcBQS98Z2EDbNmTuSxy7IJpA648Zcrxfw6THy/M
pf+hkdcd92ZGuEnyBcRIY5qPe/dYKRKlYZGTv+AtaMQJymqYeFJqqLdh1cBL1vop
UWj54Y9J3Qaa9POTJffaui89cmjfvKeOJsaBDIdxntPGDPlBiWCxT6GHeXEy+E5J
j67j5tOekmgqmgMZ8lxTx3Wmmm0L+TITn64a9NNUkf+y6/e/bnAExu7O9xhnHEl3
ObJJDTST+wdEKV75QnbJEDdFbIFo5PVQZqv09si3fwc1jepDh7dZUpR2FoLWy9PB
4lDAvzNrKPgC5Qs/0KrZ1CpXQzoiRVt/RkpR6UZy6CBobPao7yZmoFDUAmXMO1sE
CFwaIzLzSyMMXZnn2Kw9xicpAIHzutVvZFqna0vWHoH2gGaABENcqF9gkoAScR21
XvUnkS8VB5KsSr+CUC44/kQJqv4S9p5d8SfOYLyBJOY48TJaaiSiWaKyy7WBvmVU
ixhMUOimGOM8zatfAKcY+ovN9o6JjulByxvZtBO83lIx7FXc37OsUKy2dLPmxQPn
PHIVPcmOto3Cmtc4VlfK4LjeH40wTVO9dxDELUi45DUnuzG1qERsflL9fr+98Fmv
7Dqv3XG36HU6cVKHgmcadAgIVXsl2DItU4FA7y6PvzINyaIWSZKFSTT/2yf5nQ/n
cLPQx1Qxub6U48/DrkG+r7Uf3UbDAvwXNG2GCnSzF089PcgYZ9fbnsPlNyIU6dZF
rlYh+pKUBUxwfn9vO/qkffhOWdeF/Ynt4Ah5nJW1Rax+SLgaiBWJlWDGQhKexwm6
davVkBIMMWLJ7dAQhieO4TIMToqLODZSjo1tq88WxJpnFAPMbtuuJVkLtbkVzPlB
1lkhvmGVpAzwnnaL7/tqaGwrPNmMy960ALM76UKIKlZFiiAP+bCEIgqYBOH4kJft
R31MJJ4RBei0Kq3VMEdnfs24+r0Ouhz0loogFMR2kJJ9hECAyeY0cmyJnhPxkJ71
QfAl/idb11kMw5VojidQgKVBf7CkOEBpOil+u3k7wpkeBSyCTvsiMQvDu0KGvcRh
BOE7KoiQbbZq+V1rc+fYjnw3WwYQURZCgavR9FpqA9ygsUoACzigkIq45H2enEFR
pEYNHkoXMYanD0kZlyIRNuOQB3V7XAaMqJ4iykyY//Q2bim8+K7kJ2S7e3fQEv9N
WmfHUUuYPlQfnKSTgDTmyPEHLBo3fr3kjEPFmhw0H1bxIY+U7aBf1TFfNB8LBbSV
MvXtegN1INaMOf15UiI3A8GwgRaGH/AubBczcJl2N2iKNM3OqrSxNv3zgQG7/dz0
AHwb0UFcW5hPQ0p0MNNv9Z6Pzy24KuNeSk5Ifjmr+8hEyU7wc+ErKiNSFQvs1DEz
OjU8LCLaVAQuGYTdGLllcaz83aLmuIwSNhUj8/l5a5RMEb7GurSUdkW271Im9ELd
TmbTEVP86LkKOpXKQgu+//JDX5oufoN+xHmV+W8rTpOVhXJiDPXdb3eJmoz8k8NA
vnq6ApzLge2c4v7kr37FxxWO38GD/rKGM2ZvRRxX8P2FpkG+NFp3ye9VsPOi5hN0
Hj496B0KbJbI64tqWGlxz9XkyJfzMcCLS/EAHk23RSDq5H+1h+LzA4CVHUss64lW
FEuELrk2SI4DdaBul9SvW2mG9+wRy7okoVSf9/HceaNWAzp+ZzkQcxCXpK0z/mU1
uogc0jroaW+/K8KlBpPzJZuwekqpG6FyoSPoetk/uYIw8hO34Kv/Lp3mS4wM1tVX
5iMWYXs4bP58NliEFgKpAYupHwHlhyoSmwu18Au7byj7CqfIKvqiONvd2+ty4nov
UQ69ZGEGs5QEi4i5Qm1wfnnDCCZqsrIhCMXoXczy+23g4/g/Es0Kg1s84SrJqC/H
1yQ5MxXXFQCB6vcKkKTVDJoCsA9UAEg7GGZyO+xu+klm6nMUVXwsdcQRyGkpaZxo
ifeZxvdU51OR7xbPbGEuUKiAZ0FworGChuP456yT+Ri6dbpz0vkUDt8bqiOPKqey
iWiZluDn0/nbyzVijsTfaM34KNDM3iYzQzSq5AiuY7Vr5mSYlx8/TIKllbr+eg8a
VYW7UX8iCwCXTogSgTcodA36S5gS5vh7MwYoIsfUFZQJyk5dUpfrsBwaMJQnWu8E
uvmrgyWoAmLQolb/nkJJMXwskjPIdHMYopCMd+LeYRlkm20apkf/MgpgqQBqNgdP
lzai5YfLHEmWw6ZFLluRFQKQ6S5FCbd9P24y73mcVRHKB+Rbu0K6SJXPE1R5sqF3
jyjqmBTwHeM8ZVFCN3b20FUFzl0u2DMAH3HaFPcIt91ryw/0XAmLOEkllsq/UZQo
LoIUfBRvuwaeKvsrW6GW+DgD7lOlelFySeS929aKQsjOIczv0g/KDVemgtY+81Mt
FCm2BZXDE4hV/M2NVWXhgu3BvgNQO9ursoLyW0YFAH6WAfemPdNjwHtS6ienAn7L
4rz25lNMcNklgt6/pweElgkL+3U0voVM8M3gl+yfOtQnGTcRpuIvngUchgaj6Ahk
sjul50NCLzB+J2ty/mPe6p6GgsDeyKX3IWn+g8TRnBHQQPEr6R7Ka7VFiVLu6JdD
gMH5nwII80dBddgN8MD3hu1Ep9enoJ8vw0Za3aZBUij01tckdQLaSodrVEchhsRI
euUMS6ikk6Fc0GgLwMVIFdKPuXbPU9bPuVJqTOsjIbzPJWfK1wxDyu/avTca/ry4
CEYk74qwrztXPkNCloFAQWH/ZSAVcPF6OFtjLtNdVnMXQMLQDe2OkDqc8GWIAC2P
IPHTL4BSrhsz+a9owK8asoSC4i6tLuHOaOe5aabuC7YfFSZKxlDAhbGMGILJi7UU
6rrvhP5ZEHuPcymyoMIbogQ6bEG/EoJMNuEYRtq1a/EghINH255w/itmIRUHmGm1
TVZhMB2GsOL5BBoY9pE6joSpBSotULd7ZLAutewjlGEHUcWVdDkBLvT9ojxXfMJN
vZWsVKB33uA4jFeaml5iVTGDg3EhSwxJsAbKcIe0INv571ZRPuucVnZlVRJ9KjTV
aIWLyMMptIFipxE5sDLnVWoRUo5wmcGY2yZ/krcNIWGqbnd+fwgoP5fN8SrGSNsd
wPejSEH0jgGituSyaGs1+8wuo5zJ1orb+jDIGV8SeSC2a64KC5jfIXQdDj38sG0v
DgnBiBUWgy8IOqODgatYCgWH1KihGq/gOjYh2oN3940r4XACpC6uwNy+u9AtnTCy
WQNSaps5Y3TyMRpJtv8rwQNLlDe83yJ5JbYRtHOqEHHw1MH/zHbRqesfCw7TvMG1
cLKUkhvAS1bcZOsbwei/HKCrcAIKB9KmiH3hTNJRVxZ9swsP+hF65vlCk4mJZpj7
W6bJ+YN0IlNKletB3Xqxk6T1qu8gQGkTleYBSPyKbJiSxeX11BCdl1t4uJGh16nY
wTN8bUUE2JeYZos0hq4qxRdZFRilcZYewbFbJfiezPfMaUWahYc271X97s21A81+
JuM6Ob5PwbswjDz/o36S22/AjYAy9xS0/wBykpHv5Cv9uOxy2mdlWpq+BAip4GtT
n0cemy1SHFeSSxDXobQ7kqAD8aOGkDkkzNb2qMj1wm7nYHNGq4Lz1KrRD9VvUhwG
kIBkdpnICG5b8bfkgbI4pVAlGzdcspV9qvUTlQDHUBBWprtg3ze+yAZ5UEy+iNq5
g1RRRukxUU9otgxTnBKUWMbOaI/1I98lQvYZ/PIS+NRYFAKD3lpvpOFyE9iIhSfy
UnC+EDeXq9NbpF0R47oVgdpW2G27nJ5jQWmFtwD6iXdudW4wi1tDC3v5SkxQK2o2
25es6pAYGs9QoUnx0GGwd+5zAmcZRl3oQh1uh4dC687+4bP8nCy0TVnthXdGQSxj
CktNvgzevotIRMmuYLJZAnQgqzRa7pgGbocr5RKS3LNc9MuxdCG2DTjk59gC9GL7
Lb/ke1CjLR2YoYJ8bVgfDPHnG5s6TIBHk0n0FbVB53TPcFy4N7SrBZeFy+KFYRpo
0BZ9SFL1To+Lw1Ts98WTddaqtoTSqsKTVMm9cP/hUKO1gmTrj+GSXLqExMkGDIHf
ww8qC+zn8DwKKbAwyGwmTRwz0OoQbp0E8EqldIfklGxYeepyK+c3OX1sK1YDJEU9
14rRlPINLbB2gXyCqr6FVIywWQrl4xpIpVGZ6k1/YGQ2s1YOIkGwoloBa1VJQXjO
z6KVqa6bIaod2EzWLVjPepWXFfFYWX6dk7OssFb+IbrMKwDYtH8jPgaOh6EJpWkJ
pIno5TMeJyAoLuScVX7eyXigtlsn7YPuofGnNCJZnPfFwaLSCtBDEZtTxjKXNVxm
C5M+T+Cg0Gbi6dmQHJR2bl9JCyzwGRKlybGb4RVsdaurEHsnhRPG4hBGriPbwt4V
lrsn/CWFYtg+4UVfW6FOiNW3tOo0DWIdgIfTSFq0N5i75u7n57c/PIeS3822R0XQ
ePYmLtwl1U3b+jmFICzPXR7qY2htLXEdyk+Ss3pkXvyasd7lC+tiMH2X2F5BZu/j
SBdggd5xnLckNy5Aij7LbMMij6FHor9TGwrIvJPG1CUNNA8eq3s+rsSkwyH6Gfyj
8VpCKukgDTqgiSybGibCqwmi3BjMMTw8JAqtUH71zOyYAwVSL26xhBluI7E1mp6a
f2OV7XiqhTH4cskKAvn6cOKR42s061HCBzaE/yUEPObLOA0/FI658WVSDRBAPlHl
JxEpbb03IU9LxRJcubAoOHkOq8jIJArbqs94jLIKzWZz5XUYceCB9ZIuxEwCmihD
cl1+pfOaEYX5jbUNceEZEYlEV8OBcIvomjBM5KiBkRWPNgMUwx8TGMWkjYdJrfRu
IW7QzDINWu8LePwFfSI/xP7O0lGJLQabTmGS2KhTcgpElL42I1P28IR/wRmcDwuq
Dnuyr86ZmRBc2qFzCEkeCwAakelRNY7tadx8RTV0h3yJumYUabaAD2fOree8VSLx
2ImLKpij7AFZ5TBlz/As45sfQ+iaELv35gZBg9IaG1rKSa7sc/UmUs0yl3L/4Mej
rheo06/WqSClIk8dnmSbjFQgfWNWcaPre89Xv4Fn0qgvQjY4p20fa4NgATs1+P5H
bPTmmSdYdETiKcf2v17a6ayMWIvlDpJ45+dYHDjAu3uhSHJvPDgz/D/MddYHTg3I
wrxOpOPRY5sO/biP0a8K6G2PSoXzT3GT5dPh5a5gAWWoQxBsrwwXd7o4D3TLW8nd
nU/o/Jx3//nUSLBVXI0DYbSXqpNM805+dcFkP3CYkKH+/EWQyprfJUH+0RYpuYKE
Qp+d+kuRnOEp1PbPWfYwvJ422RTFix24v5zzrfpbq3cUIiB7pdl43kih3pWEDQs2
04NxXMlfhvaL/4EC+sfG+t6LNssJhUR9LG76dSbyBINJbQx7q5aEfK8C8Vu7rJiB
oi3UjXjyFa+G4FkG7ZxlrNOq/+30Zi22U9kUUc6GHNizXUaI03xWv/P8bcWX2UVf
R+K3DZJc3qIK2JhmYwmPQjwqiFC716S/coayO+Sz0mQ4Uy9pCe1Xk3Y74MOVu+a3
1cs861ty5TEzBYfNRECBxBDYepvMbWaMxZaFHZb7VtHkyUgG3jLtsiAitz7FgW+w
B8cZXoO/iUVilnJaIzm2JjgNXCAA/v6aw21VcSsbOmaJ82K5T8Wid9T/sKs/QmAn
uqoHz0v21lB9w794kMz2FXEIXNnpVfnLIGlNUREVVxZRHt8/IUQkJ9Im0Ygid709
UefG5DfWj12CJuZpduxX5wQyFGYEumu9uEEst6/Yc72X3LOt63tlp30nrarT8vWF
rv5WPSe9XGX3meplR7IRx3UyMRnCe//H48nlbl2uf9PTyuHZmsPCM4EEBS8wUBIN
TG+Lnwl3En/7sxSqH44wJrt2hy9RNvrs9M5oZbmcN8r9wnLIlL+2aZtbOtpff/gu
05lUs/wWAS3vt5ohSb8VePyhn7g2b2HT4JP59BJXjZC5aZsdxhGe6N/ZiYK5mvy8
548XCsQ2aOzZyyzkUHagJHJ159jolMV78bQYBB0y7UjXd4/iBSGdYuTHrOCXpt4s
RpZRmQbJYuT5Euz4ZVC3/xogIbT+jyS0vGVJ7/awGhZtejHIuo1vaS+8kkjt2dPW
CFuUL0FlkJzpZqB8vkhVc59l70b8N85ealHto4wHggUq4nZ+lb3E0942I9k7pqnp
pUFBqHYqSgI7Wsa5StCxQrIwUJDVCY4lG+8iOOLyP/e50uOdRO+4i0E9RANFCNHL
wpAGun8PhriaoY1Y1gUuaJLrJU7EFU9TIJ4xzWWPrMvMTlFk4Amf4BqCm9e9BxKs
dlpnIXbekK7srJVYqV2l4uwqd2RQXvbPN2FqIZ5TvvA7fX3AROyQdOhszFvrKC+S
1Y9gjFSHe6+oiW67twIGHZauUB5Ugmk3uXs9TRIh395z6QyVZiJgxb8RzUiOpERA
ADW18XX9J+gfC1/FiBqau0S9butALPnCEmKbxlFrpm7e54lyirl7CA/twjfNy21a
DRUtaB5Qd73IsQPDpitm322LdVvkLZJsfJ7WwR5AbZU4LrF4zhvTtMnwj9wgyvLk
WPile0B+sVtN0KeEwmjKHwG+crt1it85ZTntH4EiZN6GGqtp1j8v3jN9GsGJ8BIY
IRBl0qx5GbbudphH5Wup33r745AI5ld0gtC+VufQB6AJ1IQxJvyYALJMXXy6fC7d
68V9QZbBbyOHvlKfiE26z1iSH8q0xV24a5oRgW5KzL1EDjXb/L+c7Uw26G4PSqCe
oOe/WPPZrPxVHUf1H550YTYL8XQfW3iODmAm7sLRx0gfLX6cZdV3iLwRNrWRQGU5
iPuLTOP4ifE9VUwR4qa7LpwFEJEibQTAuHsDW2+5kY9H9rfWvTgZypPRON3f5Fp/
Vc3oTfpehhXwdoX4KKE+lCUX5UzdeqYFc/4wI6fz5PYzSZ66J1aLiVexPlgjsfb2
RBHQacaeWqyY//Yr+nuZhUNuL6OtJ6Wvpgyx7GV67By58IbGvMfLxNvTreYLchux
FXyNGSt0pCi75gB9K+ozEriz32G4BvzOetztiHupoqVCWSNlHuSqn12iNS2pt6J3
3l+zwgSBhJNSlXJY1NVWmDzXInmk6JRcVMpS/ma92psDevk3gisRWKMhkAjLHn0h
lhnpuUCAWpv/eEQi03eTSvS6cBbs5AgZ3BEWmU9OGeLK7dV9oSCuvwHBAVQHf3F1
yaohbqmFktcKSPeCLgLSbBpiEGygurGPuHmCxzFO4TrH90RcvWarECxF6nXIhmDU
viCppVrHMYsVGybmUHwhurL/ORLz/koobtGBqX727ikbxeeyhnmkyP0ogS7YmGmq
FVVNUqAZ5UDbh9zF6rtCEWtMZQR1iCHmgMK1FNn8Ax4Q+QbjZSZxlaKK9iuy3AtW
dLgPR1msRFJasZwjDayttUUzFyL+Yex68Lg4Bd/gUTNaeafhWaoO66Q4uZg1D0jL
INA3t5owJ5yN30rrQ6yPYuGXEpftSzfq4pZ70hYJRyNvQLDe4hHvA9mU6sipNS8O
xndx1pkg7+f2fjD7nuVWPsqtJsso93o4TpSR5aWm9CVSaWQZdXwKaYCAyRJxlfVC
PfpEMdo2xxmvSGRXYDLIuswFTrR0dzkOFq5bdIakth1bTwjWRPX1lL/I2km3lK4s
DHZYI9bCd7B40p3xto+fEGhSJLPvE9EEEkRnvxIj/DhKaNOE7xBDetto6GWa8YaN
Dl6R9LAE0UNrYAdyzgWD5bULgx9uj+ItwljBzl+wks07D82qSf1cIZOZVMigyEUe
3MvR5nkCQBAMQN6RE2L/w8rbZM7RxGjCjVHPddxufADcRvg2Pp3/kDyPdvxdVHyf
/rl/eYS7nrO0PVUJ9MKlE2mQQ5K9iM3Ueu83KP7GOwUCo8VsFj+ddZ8vMYOTTG7c
p3tzp3RAZ1OFYHfr67/LCxcyrCgJG0jIFV2Wm8WZojgXVWOyAOULNMcyTsnzhyvy
gIW7bfSZPjmznrp2yx8/4rRNSbs5PVRIFD+iRLfC/zjwJNs3pjkZThIwXhy6aGXo
ju4fZ8BxCfMw8ZKLlTxQJJOCxEl7KG4AZQY/qUEc8IG0bfypTEMui/YV82jZ0FOK
pNOd328/mZr0dZXUk4dTQqh14feayM6jakhVAg4YOH2bAt8AXf5USg6g4027XGjS
HFkm/uyftYyvHoWUYojSRBwaBkG1OJwFOu0ZoQ4FJfvhfo6c2bP/1MZIlu14qvdA
4SG7GGEM684w3Uz9tBBO9Ca4vnZ4Yra36vRsTqWug2NP02xuaqGrNzYUDJPAp8Dw
qX4r17QkoJbj3zwscPUhAJVGJRdeEKbqtW6KYupOJmsrhVvx4rXYEa3mKkAE2Fbu
cUL14wOP/INhO0MHv+e10zCjAhWj3rDC1JHxydjF95hTHshkBMJTRIqr0ALLGVcF
+ZRJ+l07hyt45C5kVD+v9i7gCjwsSZ6QQk/acafF+39wMIbXrRY8C4pVMmy5zYJB
U5a434bf1PUq9N7WKx5n7rU/pR7LjxF5nPXCFcUUcO3b5i08qzwrjVPPA3c+AcOJ
GF3tWFQqn+57nGn5LApj6AjjhWvnCbzSC1IijZUFbEpK0H2FDiGy8GC0FsurC4XU
t56zcEgKqvClaXcOnxEvsHxpCMhBZ/OOr1wOuAwlKB5s8/SJee+qiwlg7DDkr4sx
JMpH90cAjYSyUuSCkB0yKzdyAAH9E0EkzCzi6GE6amMgA8zaCQFEv6Hhkkb7bsNC
aaM4YVD1FTQ0+ukRN/ql6ygU4+RKPrxaV3DajbpbxTSVPnc3cu7Pi89Qs2dtSRzU
fRPtIFJW480bhGO7NrTgiPUYXAMkG/0ddjuASnKOkYKt7Py+62nGDdB/BswSL/Wz
FwcWqyCqH58Wp+2p/jmksQJssNeAJaRFopPISZs0CGtCDkzTBOyVKhQzQt5AwHlA
Sn4kstE21Qin+NvcQM7/7z29KbGhw/HFSEoFzfLdlGL7OQq1zJHu/vLMyu77lnia
KQ5iwvAG2WUDbWgvZ2hPCxb0Q7FM7ohpBhOl4ycrD+a3bxbgfrZh0eDBF+S9wtZh
G4MAIJBA2k3uhRoap0mZF/JeytN1dzieF8CCBTwSB6ji1ckPMgzQ8ec9OeoR/y9K
0KlPRkTEVzDxlOV0Th2U2mwJRQMAtk36VUq7QZ0uuRPdNigAk+vKu1jez/Fk4H0n
KyrMy9O9j0m8sI+XLhEtBjSucAzW1F9ILPV0NinEMdAp7IN0eaNjkZ9kdr4wvNJM
AaGmGxEOREkztW6/T6eaa6ePM6Qb+yMRaOEgCJhPSPjdKt1EoqcemfPlY+TQ6Xuz
kVdEVdWyq/+fHa+JCZ/PRX0mf/Ryr70HYj2WMUyV8JFTn17fomkPPFJLKkoBnvFa
TISoA23Hec1O2/qiTo92tyFOP3ocb9dMYZ7hQGYkNtqupDbfshlX8xLn7rZGcd9U
SOQ4bJYkVvIuFUgsa2pdaBeAmuNasV3oUyjy3m5DhSmlEm2mXFHkqVDJRpn9ujQC
0qjRDeFRtuB51MCxbARZqYH+jsyoxFGdKIDdUarQrsH9aonzFbJhd1v3jCv5MAcG
T9F/IMBdRx/6r0VhDMm30sCq0FtOgfnqI2uu9kO+c0B9CJO9ZpLe+1jiVRTO4Kgn
p+vSWWJL7R77IbC/eQCgtX2ShtToHGrF18a8Fjsgw4NCEftFocHlFqpnkcUMKJR5
0QDjDl4ybQiHIGEsQpp7cXnCsxyv3DWNB4/dPtnJX5jquluOgGV37pq+u/7r887j
M9oXfx4V3DvoAZ0OROyGko96k2Yu3Kj+E74JosGJ03+OG+TNfnt7YErd6YM0Jfeg
ubEkS1T8aY7Qrngp+xbotrAygM/hn47D5DS0NPnYTJWIeNI3aaS+AXclVbpIcej4
8ABMtzHZ1hve+4uWy2nW5UGWhOwqQaliDw+ieP31aa1aknwHfYH1WWGTTgqmUaYe
qWHmC00f6XfJtO4UVBdYbSIDmSFApkQ5ZanGjIr7C7yFqPnBWwWJWyc9XHvzHhEY
2i+N5gS9g0i5p3qiWpBWrxntg2c35WLXSjVRa+Hyn9QCG4QO6GwMA+R4GNsz8npD
/v/K9UkI9i39Cr1yQgjykJXzVSWHh0km1vBhMRVGig0V9QuaDMwTaFLHqKTxO7OV
mUPLx8pJYnEaV2bsDlPpeZVEXUirBCmKmxuDMwk5t5E2jd9+Jsx4u3NmSKJhMpP9
/TkUoaK8Ri7lDftgvONoFqmyeitOCrpScOi/sUlbmpF5sjXRPOCFxMzQDXC+PdU+
fMy2t5P3slFduaXTzKyfPJMj+QEnJRs+4Kql0C/gII6ea+WtsXI01cMmamEDaX93
VeDF7hJcXpw+eqKhHYzGtXg0pyQX6B90BArZml1FV1tAwxJvxeEjan1OP/kpsSN7
IoZIMLFEItkHRSC1VF9Fe8FBp7rthPkFiiui8RRomc4p8Dd2clEItnX8D5YzXDnD
VTJOzWKO+IxLZwHST3jOGK37kBcMpFJiioR7rV844J1zLT42hxPQEu69R5miyCxP
YkCMjjZlgK/WA9k1ZtEMtqVCL3ljaovIDY7wKndqYWsLyCK7DoizE2Y8YcWEK3jp
URty4FAYlxVrTzIeSBA8anuQVKmN8bnm1sHOrj9VAI5qici9qtUwNoJEy25Sp7u5
rWUXgZr0nUvkh/k6VmQrz+5Vztd6xYjMDmNAFRqeuBm1EluiGkF7rckdIp/w/Dmi
9ktPWmSQ8HpV8O7zeXcB6Mfrw8qTd/PzLm+BthB72MM/tPkQTx7ldVYsJ9o8NJXI
lDRejiguXoJAeGxTRbTYWfdtVeiyOfFgXwNP9SQW/XyQRKLBCKm1XNeIwdKE4yTS
s3gDxINrB/CGJ45sTxOFdqLQXfPCwg0BG2egpdZWBgxWwk2rh745tXrDd5N6fdPT
RjBWCIzWtUzCs2UAGNyU9EEB3PlTLbDLtLNWdAeGW1v/wqZc4HwxY2JUr6A3dKoa
Oi4L6Rfw9FQ3TP/cLVlKPDXICaKsGLG9XZoSmdOXi86w6pM+o/txmV4c5Fw5dS8K
4tHSF8klQahkfFLx8Wl7djGQtL7HviytTAlM8d0zhDbarv2qf8IFDFPkBRua6y7r
AI/dbFJ+8Ljln939+tkB8JyO8qcA+ZvsxPfdzEacyCcwZBo9WZIe8Sz1gmvLovoU
VTnumppPy5xdckX6qlyEDVmtgKG5CQsugy/pcQkN+GIQgbYUr31g/qST8/ofCtgw
o9Dp/neMceTs9pTLFaj78P7QH6ehkZkg9JYhrYlhCnBYMoYriMB+3PuwfntRwLQ8
azw2nQ0GjNtD1ZZQbTUM27FrEQKWbTbFNnwM7kLx3dsw9VTi8SXYNcBI+ItwP9x+
aZ34l6dFxilNgq6Xg5cp0yoC4ihBHp2wZfuXpE3CCmNJizyCuQrUupSOltVAi9HZ
UVgw/VlPbKSGq0ZSAvwUiDIMEPNeAhxvzW55JB2Vl9No3CWh+HRbBL/yv63Llc/3
kbzB3KSr5ZPfJp5UNuaioVNi6Pq20nNIE6kxsQfJtn8Nk1uyqxIkMGKmFDXy2uu8
DINSojna9A5ikGDOMRNWJzpaRuFkSQkY2XLlhRBZAobMkCNvInkNaXUf9r0siLjO
Ab7YQpF3ZQQdhOZ6Csrz1o5GjQnbfWE+ts0wRsFAPZ6TPGDF+0baT34JpiE5E4Xq
boeSo4Yi8UQ36nriJjWwhvlHKh2tBLIeDIUI8gVR728feu89aZt7EXEAyGnaeaFy
bAyJz9GxOZLfoPcBHECmn0Ij3ORsb95KBoCWg5kpPNk2dtkvLgNKAwfPcMPwuHp4
28jg7fw0oRuQT/ffB6lcOa78xE+Ow1a4nSOz4nHMKe1i4au5PvL+ZIM7X122kgqq
3rIlGcC8xkFKQFLBdoRkDwynalN2z0nVqVT9EATryxEjKZdsLQQea/FrO78FNl1j
3ba0aoUSKOhAtWW3/CzZ76nPe8O8SsqhGsm0sjmo8FGr6SDhFkKlnnsxxJS1k5h1
7+pBEORWEMH0ujEyQcFGTZdOAwaxb6jesqpuC4u2bai831mJ/q+l8HnZLbAiyiy6
muSqGVxeGnCSjSKI9R51wBqZa54Hv8N8sfX678CghR14x3sRuXN9bSn6T32fbi3T
tPARJP/m23YI4+loh50YxX+Oonhz2EW7t+q3W174vjfJEnz66waJgS/NBKPoMAG/
qIicNpml/rj/NADbePofJSb/tHAffG4S04uCGXlMQ2JarhBulVfU2Ukao3ZA7/8I
7C8n/69frgQ8l3wksl2gXqlGscVeIB5boZ9FaqVPCAk1w2XYvjd1FJlgB6UZL0lX
Y/oyORckXTGyTdlu0sK/9K/m1cAyViwaZ0NSpWVK0cYAFIn+JwgS+xCxfKvnNEcc
sn+gL8ZJKGo8CwsKre7gjuMd9cohbQxgxvvwQABw1eH1kHxYYuhZ7nnhOyQvfyOG
WSZRxRZVAfN2ahohK4kWI3jBs6I+W54yc/Bd47/UPSE5gBgMxqIsVmZvsRbTicsD
UJVg+uX7ovPWq6ZtYicd/ZzkDeR+N+5nsd6sF4sPIbZC1+bKWHDX6gNzdZvClHSN
fSu0WAbubHg2T5iPlaBRPLbRBFm9vPhMbgM5xO6JTLm6yM+QHZnTEuS+w95RPAFz
lwoijtCEuCUNtX+rHvHcaoReH9pGMURU9cizQCJR5uE1oT8ApqJ7Xp9070r05yGq
L1zVzE/XTpX+fYrD9j6onGbTXsG0so3dJLJ4FpoBcKL1QGhlXUCGQit4WZcpHpZR
MW3QDFdvrqt2FyB/o+UAPIcZfojIU2VJlPOwZSI3Nvr4nrZ/zRxmru+43Fs1OJX5
JBCuD/cBsXpycfZfEzNI/TYJ7enZ8agZL4Eu5XLY5e0L1hArd9f7CGgBmI+7vCgi
1VQub2D6pVqrg2ifI0/fpWsuE+fbqMGpk/o4c9KIjzMfRK+qqyFUOnINov0nZKLh
rLuSLnkQT3hbUsTd2oG8daTh6fbra/Di71H7EMHVDbUbhJUuFHiaF/pbDKCoI9FO
9XLRt38xHfka+Jl1CdZtg+l7km0ZaSCtA4MmPmi42mjovmjRg9v0c7j+EK5JA++K
1q1Hvs5PUGXK44pT2sK5WjEDExB7b2jCv27poqTxTmy0t8+GTEhe5HiAsAdTll5Q
MzhM/8anCwvjixXCAi/H2m/Wij5N5iKEzjrAgiXr/Aitt00qpK+AnmQS5Sj1wvE+
hv1Az8K+nEjEkrM2PEgWQEApSbiT5J84XilRlWt2MMFkON771pukB8igTKU+TUV9
fQm3mD6g+RO+05xA/MTCLpkdW8LHbgO5+jtiQOPkumlSsYVqAJYz84w1v54+0XT8
KEzzg6XD8VhH19sLTcw0yT+aQ70urQ0Uatn7mMNWylpg3XukQrgqqNfkGHQYrLdB
9HuXYU+Okn6m84z3u9zxi+UV6s8GVQBHSkm0b9De1zwqYEeb3EI0byXP6TxthlGP
Zf3LOlaaaJdybF1XMdgBSaLGzXTQfZQ6dpogjvpMJ6XFNvOGSK3O8wSa0ia76kUC
UYFDxVEcV/ef3f8iFhb/AiEGVdGbfV7LI3oPhbn2eeqxvk/+khGQDlEj9hA21WIH
ojLtHgaTSqSTnxHhyIZOFhmEsYgvPV9n5INlwe18cBybstkvFY5xQ+M13RWEWHyb
aO4UnQMEBg6sux+LqKDjKY+NS7TcN1yacuFsPEplAPUwm6N0okgdunuOUzQwDwNx
5o/U5Lng/IH6wvSwRjMXaISg6osPkP0q6PQkUKRqlpwpME3XNriLn8tHWEFSky0Z
B5DOa4sJ+OkpAWH+LsAGi4Kb8r8W24dxzJYe57qGVkXhvgcdvBCRApQkEgPk8b80
Cc/DvfgTLNVMzgNQ5NO2/LjD/TkaioGwwjO+/SsjNs0GcF4iVJYJtv5oKuYZEYLc
T1N03sFlqmZVGtc3Vft7g17NxYBqE0soZXCV5TClcP8gO4T/LuSP4UdSxJy7BA0u
1MZdkHj9qlpideT7QFcgVyuWVVFrDIySXhQbcmyP8mr+iaxtyVVddy/Q///oXuLq
q9YcMg+5msegKTV/7EMYp5925ZzsblzEy0o0TIRAKV+KtbwB85fAhgX9QvwFC1pQ
CG2JRXsfe01hWOEyvBOJrnWfgfr8vq4i2Oid4LUkZSBkAsFoLxYGBOSJr9CSq6Lr
wwlwBszQKR1OK2njqNiAm1mjhljVAURznrDd/jV549x8eSxGkOY9TcOBc5rE5bi2
K8HFOx1iwAegE9Vrzi8DDjlrZBdaijf4A8EjpmUEDniDWCs6VTjYFd0hLbVlIqRf
3Fh8fOurXzhjjW/C3wPQZ1Osye4Y3WLqSuvCZ6dLalJUEBxdTWdBfqAGmdHXnxYx
iJUQM6g9XaFSG4m1EQ2JnmorJUSyRZ+7+KvGS6Mpkv2ra9CwICEPC/rn5xm8zkUj
aqdP+ZHgDbQDb1avYR6STpquJo4z8Z2L3B5aQcHCig1dFwXrH9t0LbKK99IQewNR
O/ENoWFWT+VjDjyOrJCcHp7dGxHqvoxHKSvRcuprlqoQiRSCbWJHQ2zysFyY6RhY
BFxF2A+/FukactuIaHrA3KJbS/2LXay91GITOKROyeFzOUSW4QBxNlPpJUFOJWl7
EG1BPXazdhkjkrJIE1iWo5cPt9tId9afy+FN01cjSzDC2dL4X+wB+wGxxDIbfS19
9EryitGOcZQmNEdc3MpEVXYofZtfwTnhlC1segTRT34Zc6J2PskIZ10NHX8ai5hu
PY+X+njU8pWKuGoZc4VOVRTSj79uDuoVLN+o4Mne89Z7eeZ0H4dKb8IXOlmKbJh0
eOzSsZXCP+a9okaaf2eq+rakq0hKbbnT893VrDWo++23WCcJrL93s//M45JtV50C
FEbmYDdVzJ2nXT8ATLrS9K9QDtnzTeRiBqXfWwuGY7zi9ucBRSycmbYOq4JlYH9x
A/KrjtNrGCPTKW6fKw7GYgKhdCQI6ZvvJ8G3P0I0AshMMtrtEMkCXqkCRSZqqg6x
9YzenAhN1rqNyJQCZ1WkAwkZRRNv+GOYzQvrNOlm7DKTRv++Sok2I+qsLjN41Fia
DRMZKikpJt/Oz0c9CRWeF360uVP4Ieu2kB7Gn7jipvQy11MHg5to1TvS6a9UWa1T
AHpO5iWIDM8//1fGyOe4kzLPo6q+s72rpP2DhIchDuNGt5AdiKQGdfrVENliSm7Z
Ocff6oWMlzbxn9qqb9NrbzAD1ydAi2MO4heqi5CI9+G40nE68us/Us4moj3DLDVe
QmzhNfw0slPFsaosvDU8WStIRNgpdZ+sEFKy4McOo/E0VPmTEsOpVqQ7TeYjmqBB
Zjc+DTj0JpgVU/ZbJap8DziqztOvenEPVI5XjV7NQXDQewzTOyEOsOSl/UdItd8u
ZkIZHygWT0X4arOK90sgpzEJ0CERDJbCj4/VVKJujPF49wayeDk2RKcaVGRwhHRM
EZ3Tt/kMZA/zdkNj2eFTU/zEoTevc8U9AisKp6u7/wIQMtEah9B8NwFl1G6IFOkf
/B5XUFJViGktIQnVY5/CJxqdzc7Gc/vIJ2YIxYoGFJ3afridprNQPKE86vdPCSCX
2BX0V8twnLxSJ2pCaHcgThjnPYiEcTNjg52Mg03OX5poTiNrSv5IFE2HlQGAPC9N
gkydyJaYEboPVOZljcJQWc/XogwuDU30Rcpi0N4+9Zk2WTfuRfHuN0bALBuEXe4I
I4Uvap/6UyFHnMHMrGwtPqBArtyye49EsN+KiNKLFPDf/Qr9ll0rOu4JhJPWkp/r
n0C6dxN4nJcMtumHJ7OwzaLDEPqZ8LaHidfGRLyAZteyKxbWgqbAKGT/qT84LDnC
Mu9IHKfVcihKBVRqdwDYCGE3xAbSvI/YaVYZ39rilPzyNzEmOQb7ETkvX7H+YN+V
IbpeaN2kVfj1Vp4jQ+GgrOtbrVOjLUKLvUjMUjlcx9ckPGheGWMXt2o7wQh0RgHb
NP3veGA/9qWBx0z8FUTJEf/BkXemTkk9UxTkLm2AKkyOfT9+MKZQTeUw+O0qDinR
v9zOVA4kyVPwoDsiCzspdvk326v3QfIqsWFf7yI2vYt8PmgAlh9boPErdu+ItZ6J
eV0zHVExSsbX4jntP3qzpC0f5v+A7Y3GqjBpp0p9/7TlA8pBLBLcf8/r+Nj+vzZX
oFGn0h4N8gB2IfIU44cov927HXDeZhE5Ndtwo3mE6TcA+vVqKVLQ+/RpcfQlg1p3
Ro5a38JXcD2Gn1sTNA38g7aLHNi5dSAdphjbzqP/oavkmzFHZBCDnsuHb1wZFIYs
Gg6heEQq4By6O+65FpmZ8/drJXnPP2jzAyHiPWrsDTy8wHud5jV4hbcjPkkGu6Md
LG7Nfg+bxVhWbx70nIA3+VqGccwiofrhlzXdC8LYNlZa/ZWt4nwLnGiOUoJZs5QP
He+KCrD4GJpVbjD8Gvr20pd7cEqRpDtVLlpAjqFz78N2BGSLcU2N0j7I1ojO/25O
9aZ5jR69i+QGfv+Yfg4zlb48R32j/ro5RRbBlAX6ssAJbsN/gYro9xLfhreftmzI
kzu5Tl3JSj8Avp8W88m4ySfzO1qkD7ZaxjugRVO8IszhQ8F/YSGmITCcUo1dBk5G
fFyGjgIzxtsif9/9haPSsTvyOz+mNUSM669cJ8lCdLsISRQRg9GQys9dENMlMjeO
ON1FqluJ71teO86Nzq4jrhasb5sBg+rDQVMh+OcVp2zeLzwbtSrTwLsNhv0OEEox
yTQE3tWSIa4TgI+LnvjyajTJVkHyoKU0mpfxfK9VEpsbJ0jSeYKdSsOnAikVx+Ni
jnaukkqZJ8+iUvLfn9Xlcz/7lqxqjrYiv4Rclckfulw78fFIJTDEcRiGDKHad/ta
0u5VO0xzUK5iFw+nr18W+kMxg3ke3OkHCswxJmzbFpAwCuqlLkGktNb6VCw8TakG
gi3hL46S/3D1Z60Nsifgp6jlMi57apaLo/jhPjKn37vOsKf/jGmmWITKfMWshgh4
OKD1HKDIApbEYMXpO/0NKwr6/brj8o4KFDUE+f6jgRRZCRxkvRVRg+yCO8WzBkGp
5iCAPuYnADakOSX51xYifvZOQMDtxT/n2iGaDPusmDmDfZSQXFy9pBi8AwcdIRft
oRC1YGkyH8Mz65nIEZANWkEopdAm1TqMmzkQ1/ZrkeAw47qw0zK3WUPlos4It40f
Wiofix7gUDw7mWiA1bLVn74Ej8xDzeYuDzIGwb5+VNMjPLypPgNB3PPZcIhi4fiF
ZR/SHtsv4wU4BnkBWuZAKmzbn7CvzIF+PqTI3Eko5AXvpepAJoaswqud8sJbQFDv
BH+K+J6D0PQmrveTuP0bPGlR36bUaZAa4wF6NTLvmjsdTNA9Okr/McYtENlET5xu
p8BDEOsSNEyp1AXJwg0HJwUYPW0rpcz31fmUYVLQsyKIdOh0GfVPYWY4xQatlbLy
DCNFMnv9zO1pms3n83df48hceff16ej4oqigR7kQ9AA+AIZUx4ZPRpEXMYS+2/6D
TiaHdyKvBW9B+RHawgSPp4Xg3iBTevBEm4WNHDDqh2FxUrjUsr1pxfyQqlD8IIP4
cmxJoQeKQDL3yyVGdSneTPtz4LyovYjg8NlmS76R2WDznNbyYOY8PQ1XHqc4RyIc
QD0gNgOXWq6uqSUWVc7b5WqqWitHH3Ho3an/s/p+I9qv1ga7GLcp8pL7sXyEZ0Xs
c/axQ/tj4M0pcIgzAgXW59QzSVKNi1E07xj+742g2IBKrjcPxdtX+1QkTxTWlGbW
+8I0ZlLD1+QCgZSYAQV0B0IJhyOndLp+AlWbF+p0WNb+W2PQtoAVZEDktfD8xZtb
zMSDYkQJAgbvBqJrdGjXkplhk+Yj6L7YPz7p835p/0lIzHeLetVAbNrMbrgWuVf/
yJhqt30JCdmODNgQS+79SmbsHdFqS/ucsfwQjVT80FEUsItCEQGCXc+Ma1exYj2x
ciNhPc2XY6Q2EZc1uEO5Qm/EpV0EQogVMOjSkWFV1PLKqQVPw4FMl7n7yj0UWWln
5aZGVk+TIjX3NvCEUkmO+FWKlpJNxLPTTkJRCR8XT+8vnds7yxTrJfNxzfJ/s4s+
uBF3u8Qbhu01BuUKrNynwUNCR88aKtFiq7t+M/LK/3mij0SvRPjBwVF0/WFgftZd
VYXlzLletJ+8U/BKRqv9mGP9DjRmVsWhWX6/cJQDwqSboAEtMqOakPwo+Ixlqcwa
i9toO8tn4oYio0rWU9Jlw3nRTlyqti5HnfbKoatpWtBO1AjUdTxdbCXijr0PVts7
MNYJp1bCMxIKLKm0iGC1Jv+qk2N4ItP4brr5lFz1KON67jlkHZwIVmpsgK710RFk
QBFNy/cUQwY+xwbYL7QQRyHaeJHjo4k0YUxwo0b6i99cCyn/LgCnkmBYVEqPsp9H
uSa4DpMN8dJ5naQPFKHRuVm0bt1rJgUYikk7PAoUhluInSthY2H2k+VJj7u6+JEM
utlFkefQ6RoH7pj3I2ZExtzC1llZq5u/M09RuXrBL/DgvUMcvvQfR8X/4QufK8Oc
4Tk5kMNVBKH+dvxmahT+hcsw3dqUgs+lSwY3Ky1thz9bHUhN/I8h6dhhp5IHULdJ
Cv9I1Lu902zUf6+uWdPeapE1hhFUgMjBUrV0qg2UgmacW7kyB3MCkcI/ShQ0/nuY
15bu3/IKph4qIz1y+jEtPew8U6U+wsIKiS9MbkdWCqwu9XhVRy09dqpyB62aA9io
95FuShEZDrKm0m0cpkQNgFQvYa5veFIxaX2ElGHA+LbBpBYmItL0OulJwxpzPaRH
vZy1EkuuAmi29x0mr1E7IpPqYELFUw1LAeC9op9WIkLItDl1LWqm232ANxt868ZS
wDFvcXz7U69KYseSxjIqBK4c/OSw4PwbqoojbnkOiPTh4K8cIKP3edYsng3RMIuY
2LFfh9tcHljxyvdYqoPl7pWXjS+8QF1KQpEdlQ5N4+zApB+h6VlRLG1UDXq9aK0I
s1jfLi8Ei3Gm3viYxFkWXPjT9YgUTrIFmIqtpk93B6En3mCBTXgBLFpQbZyHcncC
6BwVq2UnLvRpbr/5dsL5u2a/aQ82hNXZTVSWNMJG9MXNml2aU5juWhETK8S+hl9e
B4m+XbpJLbTQFCstHrVq7XpCj0KzQg/J9MNC01RjPklqwfJJM3ZDkP+946xYyi2y
qUnhoTu2opxrB1mKCMWNM2vhrCc8kt5jJHOSdlTPVQO8QayZ/FicZoDqg84dnnCB
eIVHtUS0eJt45ApjMpWFU+GDcaAoGZ2pgsUOCcbs9IKB0+/1/qFfhRusq8MpCoHd
4Paru4peybptEjN+KdXrN93pS9kFhNGFF0qEkuK5lljn3hok5BrDb2YUO+jpQe+U
P46uwK6imArzsMcRgg/wX5/f+oyI8nev5IielLMcIE12iL4CME6xXnFnXFzpc+yV
VqCRgS7Q1X39SM6oOXFu6TRIrMoEjpts5m8szIYlbOonItAxD86g55JkAIFVvfqd
AxnBqTeNZ1BKGM4sZIlCKH608lgZurYErELVJrs/eh560umCANMe+q65Jl9QKVAh
3VURWRYNMh/Y5EKmGlAYZ+ZvPUX2QQeQ1v6TbatrA7euEibIee/wMH7xfqBuazS2
kiAg4RZ6YP/85UWxLRSaIvrMd5kVMH6+0YOuyqzRHoiRcnwEAIDXmsXrH3+LVFP3
pLpuoFoaZsK+QaZCiWV96HEVRKX4OT2abKwV7UndVzPlONWrpCEUs7IZPCJSSJO3
Ci02G2B6SQQ4gvIKR4u6LeV/yKiyc+vSK8K4geUjxQB5mxXajxpxH1GXrNDyQAXx
BPFlbz1rvdmdCP+lYwm2+7mVqJToFpqZ29bOrrUZEqtkmjQ74CvZnKDj761GGy51
M2gKHjUxoUecE2M8jeB/BO0shIi61Fb8L2W+Ds8YNWj8ETmuT/WOml/p6s1hANzy
/ngXdSIgTZP+3D/Ndl5teskWMJjDqmGgL89xo2oP6G950m1OBvxYRZzZ+Ke2366J
cenBrVIA1PVbg7pJ/RPHDLRIQ4Orns+j2HJPWPSTeYC98CwAt2hrTcf/V9UmPYqo
CFKlL3HCv2jItH1w8JnnF4DGT4QPjM3X/NiG3BBYckdJnEC9QgRqHbFWBKe2YtNv
JLmzsD7+cB/A1+lfzS5nqgvd/anVeCf1CKxMGEXhEgyqYicI29Ufktj2u2hM7MZw
+GDETkRgx7ISuRlpY4QG8elby2wvum14sl+krDdpkuYeh6BI40NPSE7Itv5uj2Y+
eBfLHAkhXDmKKIPMEkKA+5dyP+yvFPsFmyIWKIjAFUssxpHm+Nlfb5l/u1wcF9tj
08fRectK1zRueW8MeZ8/NLwhtx3mQTLlW9uCXyPnGP7Kz2V7mdQz1IQ2UF7xM9Nl
EP0ZILnTFH8v6Kcb/YrbaB3T6H90HsWd3AuAfJK5MnQ2UA90djZoj3PgVQT3oWIV
Fzd0S25xzm28jFdxdKdJRr+oX//gioj2w2SznWeV1UG9RVPgYSmZ81IR1cgq2Tx3
Ivwyc8n9cyoHvQlya6IGe0QunLbNOsvVPWh6vUJyWL+bcaVfD+YN4beCx7B1FHDo
Afqw6lLaY7pyP5mg4AwF7g+DyYEMUtls9rZlu6wI/3ZnEPWSkPdKuKeHYcBCWvFV
bs7XwGKbiuIXhCVjnwM4YVMJZe84KwFPfAG4lhfr1+bekKAMyfMO25ZdZqv7OJRU
/Wf/ThJOmjbyiYIq8VcXS1vbpmAichGy/dCBN11Po9BUS8mh3BLeTYJy2n2Bev7o
YCeRzYvAccSyL3T6EYy9qnx+uJT7sdacGvDEsdNvarKxqJJIP1kNuCJYd0Ynavvu
fqSTdkHuuhV7L5GoYi+2owdALZ2W4vTMFO1mycUqqyeeIhtATCoGYA9vaGdHwfV7
1KHQgqHMetvpTRgZxXyuXQLNPuf4n1Pm846rnPSmaO+ZrwPDZas0ovzumpavA3X1
DqwiPpWmtXvEc+7aLU6hnxnfyvPOhpEoB5vPIf+hEJf5jKpqo5R3ynfudGGvfEyU
Wewg0TRHA+aSb5lmDfbqtyWza6ckGPRZynzWof12A9vzN7LSLGCmTP/BattarAeo
cVEsJDvdhPG9IOkuXTlxw8zwjoA4GqVMc7WAvifbLQbGvK0uS28WaFKTI8O6W2bQ
fuiggFPpmR9j1XQemZUPGf3gh7+lgLwQ14eea38+VMZOue7j+Q3n7UXIq2sfMUn3
wzv4uYPDX6bVyXLFf9a/Ps/EjOEa9Uhd3AklEfEPzmi4x+1Hyp9G9owiB1tNmrLk
YQkzkh+dOwWLct153WhErA5v3qJtrrnazySRLUSrPkibsg22PW/I8z4I1/SBuxCT
UHDIMh+IzZsQxjT/gJp3ZFQcOW3k8cmB3IhkSZeiQFXgaoVEpNX47lYehdnj2inK
lqp7j6HKOrY+zGU8LCIrtp14L0WVSbdhD+JSNrsaUEXQ5jfNNnVUqALleU1mrbLj
SKTajgV7m4RzpYxKlxIvRar3VE8olUe5h6XEbqsCHMX896IytBAm6Qjqvh8qoK5q
zgXH6lCnVfiNJf91Vf244yEhSOFlOdZUcHck2akt8ZoUcJKe1IWrWPjofv+1j0nF
O34nm3tWKl4WHvUEV+fkukkrsMK0Vh7ecufS3fj0LvM8ANHjHbiRLQbd1YEb7nzs
ZVJR6gGa///i+QQnTuLiQaenZICuYLUeLwY3j7y1xaHMozrS5IldHFYzrY+4Lhqh
6OskkzlsBzqmI50XUCiJIAIj2dS2iaHKpUo+VKcid4nS7hAmZdj+oQIHdpYIIkyD
xgRRGPojjF5/KXn7rRxVEC4EtDrWxIDkhSJpeGL/ViWKWZiSeXtMARi7K6irhnBQ
CNI49W4bXRdydFLdeLwDvLT7jvCQddfQDMnV8j0eP00VRw/OTAyGQdVzmS2sPBcF
+av3UKyJEpbTB/OhfhOAQBO63dgsuQeT25mEYPF9+VqN+BSAC8TrIYWW8jivDJM7
zRNuRIhUqjz1u/Uc3cHUy4opjPHOMVuScVp0kUVShSskaKNziq/NQAgEJnmk+kDT
VHi9BK16SOWXPfxrV1IwxdkhsoQqNlYaZCEcwoZXqKqurhZDz4C7d4MMxgDj8vlo
y9ENKWIW2J8A/ejMqNS73Aq+bdUKtomMg4atgA4TaFD9kBIZ7SCi/kk9MrZGCz3A
+1d8LF0SPspT93yZfMvYEkEy2RTULEuUzaOYcsZg/qz1nBtT7WWgKmpq5YiFKq9n
PfH6HfSh9yFXhFOKB4Po6WDtSzbrKHXKmWVoOvcMR2O3F8QsEXkxfCMXUaD3uk4y
iF/yWg9Np7OISbhtqz+wS+HQ/O3zs8MOH+AU0sfkWrb8bHnqs/ubNukMYhHiZbTx
+7ZiENJ5dRkdIpbvqidx76+aQJr1pHsO/gXhCxbdinThENZ0nRWAxIpRzW2+Xf1b
4RfqGUas3sHEi6qxUE2gjr1tgQsn8c3d5zJ5KmWk5PbRqd4ukU/Tl36MmJA83Fxd
KfG31Bw2zIO/8YFGDR7MqnsU/qZ5tH2OjQxlJEZWWCDVNphIk+1yPI+AwMVdEZOd
fNf5mgLMu7xYpqTzhSOU1XZTxFwWI5Sj9rwIL/fIq3g9FdRHnPMBwnxV7NyMN1BC
ttrbyiI0ntJ/kfcGyB9PvUMH3tPjZU5SuxLvvUDBlp1f0TqYDZzIIuAyQdaSlmrv
Kmpep3ea5gxSnkQDvUbBaVLwH8AX6GvAo+f6nSaa8KuIfXVIhUgSUsJzU5auc8zS
DN1XTx3wk3QQs1vvuqusMJ3+5EAu4PHle4jhAU40csSp8DiGfnRDeqp4OpXtlBps
5q5i3oAsGZGMonaiLqomzktI46UJE2WohCDm8TBWmZygmcguf8ZpLIDn4aAXMfH+
Xmi13keElQjQ9T63NZoofjEr7O4vjkOb464wgEklO9BTBkfYJWh7g5fxDfsv0rZn
jWlWTIZPL54BhD+k4cL2xebithVAUb2mTkqa8D7p7Gy6Q/jVpAbf2wzbg0Xxvw6S
asQsLphFVw7E4QIjVpyZPPeBguBDtttxbfq+gcRLU0T9G4Q+JshEfIOMS27JHHJm
/vaA4bjnFhIqthls94YPp8G47mvaxtYIolOIiPXB3Ow5hMlULHiyNFw/CmvSbGeL
jFp1KQTKLDJz/Fgea46T8KiyWOQ7nBUOiu43e4jveMvWZsqBXigyKNB8tfrWGIVJ
N3Snwn9OhQ3c1gMKKXFX+9S7hV9B+XOuCxXe6Cu5gbdjNHba28yYV8Ql29Bvzi/r
P8La66NyVNf65wWXvvjohNglpUnIhc1ZopQ6J9k6XM2LIJEtk7j4/CNF4CpTKqxj
MRRaIsARnjr7NB0LKaR6NGaSDeYquwIbMw/Wwb4Yl55MVlcoDjsyoBkSuxP8e8dL
65U2bOsbs4q+Adi1qAGszoTikKc4RGMS/G6HEvBdrMLdTGIsp0K88ZTZCLG9e1ZH
HJpMFb/0P+80XvFEm8hEEdZZKri9jrK/S6aJnl+VHS9gX8BMyzve279CoHYE1Mmn
X3j4IaOyVQx6URFJ5CFKLMwbJANBoOdGxusLmV5ZKhQMMHfqOzIUPYw9seeheaoa
g+30Yt4t7cbuZ+kYlTSze7ewmwZPfPhZVjP6zZwtEd5iWYX5BAfxnx5008aX9L8s
XIeLjtU7T6sa0Ny0Yo1Zqu9BJqL7gWxoKgH80FigkDabIScdGtlHzYGMv1TYlQfZ
pphihVjCttI7ajyRMkjar5ufxI87ydoC7nx5AWueNuEtOrnJpz9flKWAqtjl0/Td
37dia3GiYO8FeI/m2Iq+JgzwiysylIv0Nno9uxZ07QL7qXu5wS1wO4e8CnynMJjk
KQ6okaLeG1gXnrd5X82izKJtiVbvypLRUyCvOgZcbQVjuvtVjNtXhliYHeKqRMAY
WJ43gfqSHNnvCChmd2Kxz73X0kgYn09nPafnS79FmzWs8dikj9GsZnTf2oZir6dX
AHZP3nuOCOMVSxBMayRNBLWLzphMwwZE9KJGvAQTNJ/vOWeWXAeCcAkB3ozry08k
NYJBG7m/hcYIJZKpy9AnLN2/J6TruA5ciwRrWIsCg3wi9OfI4/vk8f4HXJATeLpz
p+R4HifhD5HfUoeUmcGU00FLquaUWpoVxPtnDGtGJ6hQDc2cv3leAuPVOkh3RDoZ
cFfqRVDNoUzYr2DL3EXmCjQV6Elv5kNF7fSAek7OEPky487NxMpsLFT8JHhLNsAL
Oqnhebx3O2KYtR35Zg8uE2ZgxpDK1vcZTt0e+PkJsWTDifkwfoZSBlaAHXVvToPo
C5P0vE0bgS+rwF7IiFrxJrNCrHH5KlLNRzfqgr3FOJGNeKVW8ObwE5oAtlFenvyw
d61oEoQp2cXPMlgxMayEJCwkFDZJFj9/i1852Jswfig4mlGXKE/BrUuPE2RtUom1
9foOqwxqJkL3SoaBbmgmZE/RwCHGshRhbfm0veJVsVgsSOTLQANf+gVtZpiXUXe8
hC6IR/0zIdGJ9VX9KQOECoWCB4TU63n5xMwWcYUNQb9DIDrsLfjoy4zQuO63gzV5
aArE9G2JuMNfEeP74xeXae2hDebU6Jw2/Fb47hnQvN7+tiok2Z6WFGHBCqBcs5cs
yFHVCrC0X59gf5X9bfyqvJTjepQFeihwBWOeARuFDjUzIX6JuF2t+ED1867m8qaE
Gix5KcX7AgbpsO7kwpmV7wnw85SyHkevJy9yAKSPdCkRRKiPXuHsckT5jta19mLg
O2xCcCLxGWv8te2MP6rF+bepmdzBgDH22801sHqnA1bWuGvZL9sZyorhuG0SeQnx
PCxu7fr/DsCCtEzOIBbytrk+Hkg6UejSyhr656gLnmZ65BJppaPAbBKp6Fdom3Tp
oZ+/0Y9Pg1oH/57BtUqwweibPTvfzJr+h2UFBORfekyHq4yajeXkoPO2OHgpfCGm
DHpSx5twng+EMxqhATFheY+ihtg5yN8327hq17iRKol17d5u11+o1NATG2TsWY9D
WOh66jZLrmBLkFSKN1jaA9xXWeiNeMSf2EalF2zfFAOFrzdlQ8zs4c+TJnNfDNRe
UL9fVLeleH0pg4fBPFaIXHDjaVqJ++vHJvrmFagYNKib/Z8TCQCBJX91oXp/trut
lHWX2FBNaIIfgTyFpocOU+/Eln1fVKqBFdt8fGFtYZfAyjm2wrHRTYqOgHVVpKxg
AkUwb3386nt/y67QUwQwkzUIhrPRUzxGQoQI/2awf2rnNRxlIKVDA0v3fYkV/K4J
BzaX0yvmtXqZ1zz+lG/yPib2IvJOQkN6QIw3TR7nuGdmrHTVzAmAp+gGSITfUYCU
G6Y70qMdW+HzKwRWKeMLlmGBbwVtMbMR4oW2sa4nr3wc62z7/vkpM45/qmSvEpXn
BDsJ43elMj14KY6qJsy1tMsBr82+OGiJZMBgS0x1JKiLNitjwE5lS9LgGnMO9v6Q
pfp/V8VT7nDm0G4l1SCkhxNubXSbUNGl9cxh2pJXeEfybeM/n+yMRE8qaiMgCfgM
N2Z++KW1+bripZlBi5lrJwOrRDUAItT8WifoOOSEI7KpcLouF/LmfcSVR0C1OJw5
T+yHbll/enAU5w2GGADcdBFSyVQ0xuug4Ufw6RkTjGnovYOxlQpQ73hj1nCK41Ia
aYNsMXut1zJMqMtIuDLWC8q/9ZSBeP8AVONMa7WxSz0iR/vI3mmB2yKXBj0VUvLx
d2HmIxeqGIppTlfumAlByCUwn8S16shGn0t0EOMV9yc7fPiJF8+JylLXKqiDxO8F
9jE4DncDnCgZ6WaFSawL9FNNmTJhojxi1YFVPeV9ySo6vLVirYbNuIAkwy2q+O1V
AqBllKvAnNa4obnPPrHK5tFk0vmAqBvgKfa27l2SSu1hHTcp751H1JxHqVRzCqHa
TtGwWOUbhjafG2TLzSltcrRhlaU4LYgLGo1/q/HKoP7lf4Z6/zsTpfi/LLVMqCUT
Z9hyt5FBNiOPYTdAHO6y1fWoqMFLfjN6iwxsDqT0Nr0Qj+V3e0xbOTHM3f854aa8
JplxgX2n3BSh1gPvpcvdysr6+UJVaJ9zQ5qSgziR4SCOSzcP/M+L5uSMKtPrjbmQ
ae2IGlSpGBil+CAMe+fPXAffRAlBEiCe5ED78rlT7EARFTRzUekFwwC8UvM0Rq2U
eE87VOmh8tbuIRBcEt3W08U2th3MSgo93elIE/5ZFWTANy+A1o7PyawsyA3jFecZ
6v3oIRHxEn3VvadWurFikWVbUPRCmzy9OJrVWVBHOL1+dI77R13YuCrl5KNNeoqV
17T0PZ3D1z6OvAqjtXidJ9dEfTGd5cXHspHl98XJT+qW+vPv1pVjx9OXF0t8fzFI
U/NSGkNB2wuf0uufnqZSWSSdlBDsLyKSRN6QHJCjLGqrRUEolYUtwxqD7ULitXKu
OOQ2gE0m5NsrBvSR1QBw/oKdMCsKSaRn9rAvufbVs0nUkl1e7WltiTwpay6h2f3u
qQ0lDAWlMSyillRwSayPwwT81rNW7i77Rr9C/NuvME/JauJgAZVmAJ6ahba9dRlg
KV/KdfrqjeLyd1DkV2vB9sfA+Lw7TdINOM99Qfk2W6CNb6G61/klynlGpeNcxawC
hEf0gPdwIT/9PqKz4cQS5UXnBupHnzm+4WWT79kVHcC6+byvXkbOF529OoGf/h7f
18UBfyRqXI5eaKMw7uxlZWsSecEoud4RfGvoj9C5j8sRv32Vv1G1rU83yc9mHqTm
U8Lk5z75o43kEYUe8rcvUTOki/g1AWqcf75Z9yTvisjgxymhvN8g8foaSn2NGcL+
q8G0yDdG4Rt8SPGfufLhkpQWcXxgQhBGHAN0FWVxerf09zytDF2PICLRyhgmIrsn
Uw4BCJLTTIkY1YXceJN0ScRABBqw/XycJgKpR7V8sthvU0j7wyrcbm+Assziel+F
fuffxuhoVB2FNwAOMy/bDdOyyI4Wz9N963PgGGga/Yzl2JRVipO2HKBC6fwhEFve
XRAQ2xPGMmSRcdyKBGtX/SRvv7+JvdW+UIr7T7SVkRFTwHMVW0AZPR3JkEHdB0ML
HuqNzexE3tkKAdDwtnNH1oggHVDV6CBJLRGGqi0i9Q7av3hgu9oO+kzvRGYBkz5O
Zv3lOfn3xms8pXSmBU7djIHZPiAs325E7GkBs64oeDibEaTbZOJnUjRDe+zI4m1p
PMmojW5utT2Ex5bPUgndk6nYn7wrE6R3mmaiN+w73y3qVCzcx0ZImeL+qmoLof/A
8cCQF5TP9QiVreL3W12wtH92Z2LNcH7Em6nwLfXP/Zeh8HgraBOjBuWTq6hM2hM5
ISKOWbNrKEs53NKkDO8TSzkNISNfLsDfQtj6UyNKgpILK+kPlqaJNcXfv+UKA62g
WhmvnYu8CrviveDB8ovrQJCYsmchsVXHslrLZ/s1JK2b3xrndZbH1t5mJjNQ2QXj
GwKMALOdRDNSZswlnOKQJFkwHjjHAkjKidwmbFm4j5IK8acb/tSS0c+w/lyb9ZBL
JcKn30bHgYFQIMpAqYExj8fbnzfMeTfaGhlUwh7lcvTVTcJa/JjrEI2+HIR3U+4H
PQDpulAaboLlDol4CWD79j3mKMksaw6uUpL78pYbwOtd19DLkqGdJtN+l3iG2Q2h
J2In8JK8kaXTfeMuPF0wwtsNk/Ww430rnjlaE2W62dP1cyIFRN0fWG5CwKlycMI1
Muvfd80hTk+ZblxpggRw9sjY+QvGAeCxAnbjSJNls6XqgeiaS9PRuaeuZp7e5xBS
JcozQGtsiTrwtTY4jo2VfFw53jluS4g8vvbNYTO4wWoBb3j65Mr83K78Pn+UQ/Dw
vgLQDeWlaxLOEOqRcUKAoL8jkOWLtXIbvVd0Nn/Vnh2vAkoop94mZgdS6f2WjDu4
dvrieW+4GkUxK/UkXRgyxzyKG3JUehjwwhxb/o5yu0aXfsh7hCf67XAfZcGt7wQB
kBQayw8uo9ATaqF7BK3Nn97yxLinV6ffB/6VCAzgUt3EWzzmQnk8YcaEfBudqig+
hH4su4HhoJy8LJdv/meyjeslD3sYIo9nnAdRg40AJKzPBzk9dHmhgd/aQfigzWZF
cZYOQpZ6hdfTApZheKBYvTbFfefp4FCZszkyxwba+uyxgkAnq2mXFJnDOz0c/qSp
kYQmMLStmNHqIccTjNM/g7lwvAuiLVoVBNeplhofO08/EQN5Yt36OjmqE3TDYVCh
QfelAescEsW4yej4bFm0gpvvnAiSftvgW1KZMsmP0g2NGORqzKiAUnc+uACWQjjf
aK/NpQQ31s2HWDkiA/9zmQPRHtyAhXcOpUbc7fS88BHuX74npms2kucL/K4PFa2u
jZaANMqx/hXz43RkhJeuBGGiINVAqXq3a5Op2HVm+8GWp6MNjLLYlpQyZkNeVf37
h3k9J4/PHaXC4ZZuSsF+H0ziuYkiwlbT0j2n5wbbpafoJhfSDG0IYM/lept4R6dH
PLK9OO0tvHSip6RAzi/t6izj280At+cZ3PlXv+aBD2qaoDf0+OqexLZ3Gs20zRAz
wqFg2oj1U6vHp9c6AuCorw3vBuZ3LgZvUpCbjUwEuV18QCnyXZMwtthPUxr/KhY9
eLiUeYskfOdNAbF1f4zaC6bC/KDLyQgdbQFIX+YnE3+RoITlc8AYrpzlJ40R4n6r
Ix4WZsED53sEsRSJaXUP69z8/+MkfE4U9xTIYQ0a8scmfEGUqeutlGJG2PLbXrFT
/JTWLhGJrjXLeLDFk4kG+VdtbVKcHBUZF4jm5wqupHuJGIX0Ci2zhGG5pVwLSZbH
r8sf5MGo0S+/SoAgDwkt2kFxugml5CDMYumzD/XmjRQzoudgVRuSyh6yfNdc1/Yx
H5Y1Rv7xtsfTL1hXg8bvCZki4IBESqKd8BsqxTkCEXmz+F9pRkwC5++UbgHh388a
RWHhmOvtLyTAA23gQbjNrgzc5bEaFtf570CzpoAYsvBYXjKQ7c0pfDlllKIKrAly
4tShZF/AthFqOToRSnlpiUIoA6x3+LFNC48rbVz8eocJPp16G3809J+G5XVa2gF7
Oe0JnN+2yZ1thGeHfgtVG8rxrQMtqNaiUbrIGTNTPIjso7WE/naRfk08AGhB8f+0
yZBMm1uihASvQUCqVHi9pAYwciWrq6ggL86KUi3TtqaGPEg8m5LvBazgPOZB+vzv
Xat5adNertJt6myflSVEGpZ+aF00PjivNvM8vKqglGvzc0RoI/Y1W/Ldwvi0w72N
wH5Zs1uVP5jC/nqI50zp6850paI2OaEQ6U+sYuOLWSPJKl85YTrcu7/MhyXKFc8o
KSVl64OA/MzH8mkuQz8IGsLxGcoKgfnK1b5C4CzTbkuAUFVbKrMy1kO6HuAo7G1g
3VL1PmvhO3BYKokVm1GFkrXEYl2qgNFmBGLpwwY0lmgzv9FtFgt7vSDr0e9fKHCk
GF9C+TcAarR1uAW4KaewMjAOs7PSUJdco0Lv5ZpwlJskbocc2u9SjvzWRCL5Hahg
9i3aNI5UarP28Ubl7rwaomkGdfojXtGjk2sU828s3pmbAyqTtcuHdAdRFPTNhqWY
+1RsZBfyg/8eHyKKaIPAteE7Nyh6oanr2MI5YdMSGIhTDqBJe7cU68Uflj0DGJd2
cAUqddoihCkrqcSEm1sNc19DQk/bLxKg+qSBSQkkjhOBOpcRoIr8aAQn8gxJ0czc
mDajJQb8LvJon4lYB526CDabjiEYvq1Lf3DdypnMXFsFdFQUyBKvunpi5NMZLDDq
j02jnvKYoDquJHX7r6Tba1OyrnF//iy0fhk35hudSHeqcMD0bw8vUDeVD+JtYx8e
ZG5JGP3A8qur8yrrGPX1YhjK21gnrrWeQtcXA5OJaeyWkxFPvR6yo70ldVehyUkX
Jgog8axYJf0lBHdU4NOHrjia05wyxDdm0sMO3a0qtixTdu0ykfbQZzWMHhQgh+aC
W9horfwG1DMhBORd3blUlkncbD15d/lF1ozW5gJcQ2lo/1AV/t0j0zYyIKchVlYk
xAWp6oES1v91/2mdSwjyc6LTQC0CQvV43gCdSHXvyQ0F2Tce3jvdFPkNbR+3AOZU
hKPiPfBgKPnH0YHQZt5n3yxF1K4DqYS3zqC0bs32fALhribaPVI/dulEmkWAx8h5
3xiwcQA+gUWXZn2mIGJD5hmc1kQRSsjN4S3XBuhFkNLoXmA9KR+AfU1rSBG7lWMd
2u83nLVtRSL8T3HIkEXt0+IDthyAWs0172bp5AtgWmqGmD4Db3UguXsm2NKzmS7B
q8N1B514WWkwlESV8SqhMnFzUVYj7ImXwDKqFoAwjcxcJbQrK7EflGGOHHdWdwLz
EBYVypTQ5ZDUYlEt6r6I+mdjilJDbOsHWDdwraNQmTJaKUTZDyfQdPVBOO1HrdBa
36HN3MrcBnjPZw7ETNaPRCSGNrSMZbnxrgFtSrkCpgI5s14Sn1nY3UJhN+GQVQTG
hdOcReXl5qp28mjQnCKd7hnYFuOYggBZch8XMZp98pe1kMhRvl2yuxFLr0IHLGG+
1MdtH164+NrylCgHGDE2AMkHOi/uz70XO5av+Aqu/Ba1hhiyYn3L8lMgKilnC8EQ
YE/4UdZm8JpTQxKbdlSjejnyg7MO3aNDD/fuhYsL3Ws5NXfMXpOKiJ67Dgdp/70u
MUrsZKSlASLwngfZGZ12Ow+M4ym3UwtEGei3SclkyeDX/ixH0EEca4kQmQ+6Dj6L
LOSgkkTCVkxIEP7Hm7+MnQ+apVpukZzicpcpNzkX/1VOKTzJMmTmRC6n6+XooOmk
622JT1Oma0H3X4/EIaQ/BiYXgDowxos05xzwIzgRODz6jUUOm1AMM3TIqzFbIqA6
NpLkN0suZ1975/36aSGPbScClqyrHyITT+gYJYzq6UZcsAnQDcicB8mjoZX/xDes
PjodhqrqktiKgpJLGngnbGeFkMSE6ZSYVtYtJtlJ1VOJkMC55To4LdkqgvkXOF3u
jGuKJoXsB3zPINmFPoHKjeID+wq9uwOvlGK2N8GkDyLvGNSQRKZO2aFXXhgnT99P
CSF9r9yNo66ypwHky2SzOrHUSDELt2GiqCeor6OhWv4R6zIWB9L3Dv+xIDljAXMI
DQ6uDEKzW1hOn6KX1G9X7g8igLQEDi72MZBn4HnZwuTmmbbA4brDHx4OCyOfFU8h
vyyUXVP3oO7yzouf68h5c8jOLrGdeEmJdTuydErOO0I6ZaIdiGd7ujiwIFSvi48n
crWxJgR9oGz+Qn5VBfEtLbjyCGclEXljXJ7weiMoOf8ZlWNcM6ieiD3BAeXtZN5v
lbzF3GiMBbEGa2s5WAE1eduUtYEkfPKs6Btd2WgKI+919AvNOq9OiwK7mh6rRU+i
4+pm68FvHpuXKRSJfuBzzErU0EgadRA68+T2NECPby5XZ3ZIt8tW05balTjNlpfA
b2drEZC+0BghUtPi3uXaGIpnjZsFYsKu0PtNP25RxiwGytktI6oUa6idUDCb6BdP
zB8xbZjnOk+AqdEMeiwpfNi3YrQdP+OQJ/L8jS4BlkLeel2DWK9KroxxmMBnbThV
361uw08QOSBnkw/ckvUAkxTrSMnMBeJ70P5z6VeSXoWUlhf0HHaWP6iDwUeo/HAQ
j26ynH1Um5nXnIVppoMIFN3Abej+Nkl8N64YD1ePejwbVbHvBiItor8KgB+SPehs
n3pdTrR+MgV6HEh+X/nckHalTEiyjjTJdm/DDI7Gw5/t7rpH1QCCaSFCOgyt1sKL
t9pKBU2HiS6TQkjFclwEAzRw5GjtY6kWswastO3bNhrVUbgCua3QNkZWlVWmmeUP
U0m35vgauFYTqtfNRjYGytnK6Ks7QwMn6kVKrJd1pT1NCwcg1splz+ZYkEU0qFaN
WTIE7/IqmEWBuWyREprcsXLY5deOpEJOYQbNBINy+7Gj+Rh34CZF8uoDfPZvoY0Z
5HePdcqW8HgEUcnS4bwJ16jbLtRbYe/pJUzenuuXBRpAoZWkFaK+yak3nJ69489p
rtry8eOXQX1R1sLX4Wq81m+IrG64XlqLnyCq7RKJdUVeYBj5bmSS0YIxhJBPk0Q2
pvjMSwZa6Yu5h3MYvKJbVRETPZK5gn2DyjycGaUx7t/FtbgItHYErygelw2n/wts
Xc6e29ZyHkMZS3BAsoOf7wRh4jlP7vtws1B+6tvhCq08rA3Jt151zCp3lPoZuP8j
iNVqywJfMCdfLerYWVQSlGbSq0npt9CGSqPhrZj4Nv3hsoJKQ0ILHcz4km09dQ4x
wrtLgbSKpx7gyUQW9+FuVXVhfWMWG/aLYjYUxxSG+mLyEJVWPOeyz34GbASJvtxe
QVQesQCE7hbDXkpIIaZk8UrKp6VW4RYZYnE+lfl7qmMNyBWKwy1cN93FTWSHZCn/
ahJT6tYZ2aeeuR5NIJOXsr0pzAmCRoUT9AFnLKDC8RoC68/VQMfPPZDgxVH8X4M5
fd4emn/M9nLw9MyelDddi1uI5LcaOeEvWaPXd5/L8Jf/cjLLHWh81UcONhfsKCf2
ZMyecvVpoKB8aY6lnPQ5LCgZSTZG6q1xjRI7ymOSEBqLI+7roz9JrKiQUl+peKms
7MCGx6xjxEbrKGiVImmZv51br1BpOXdrsh2uuGAWpqS8+CKJnqv4DgrN7DEBSTWs
46veJ1wTHNbzl0VqthTEPzHcEZ2R1p4Dym5s2OkfTWVd/vsQydhah/S9QQupakIn
tSDf02RmgmVJXT85v5J8famOt/Lbk9qHS2EFQnsi0+eEjI6Lrs/qla8/ZTJOPSbh
SS7m0vE/PcEmlVDRJa0rVphyNxvVaJiCnPKUo1UPj2GVvNEcL0F8XBIvTJHWgxXI
UPiEuH7YkMve2ngXd2R7z/3HZF+A8jPWgKpNM3sSOvr5N39gMQnmpPpJm3gA0YPG
xnCgqkG7fymCln7chdfMIGV0NH21G4HKNGXzGZwlCP4OLRmdFKZxSkzU/9bIGJEX
lhgcB8/Wgdwy1CxciagpP06ncXQfsRjmFiAQXRDIdc0+YGj24+u+5BjnYQ/22pm0
CCoKIuiUIN5V3Xxre97aRtJYn3fddDgWEoyZ3tNZ/ZLcStvFHMqLQYi5Uj5+W1QL
Kp5BqMzTtNqEv0+YqlsdCOj+geYTqci61+UPoDIEDqABYhyupUe/AvIJdKJk0qaA
WdzOxtDGUi+UWO2XHfrBkLdhuqKlgHuCXlNSuLXhpogPVkQCl+U3AYrmTess/Ozg
cOtR5gpqYz16ASGc7PI6GQqDp8CobR4YEEarlCrsl0L7kM6NkuSx6dW9FCiANTlX
VZgFsbnFINIM+gOg3f/CxI+ZcAhuE1Y9NXtrVZDaT7n3ixDGYJUkxEBuWmzCth63
C/9h/kCfqyAOHmqtHzRSIMMmTJpo46dgAhpgaei9USWF9yoyC3GDBlVm4M2dM8rB
fZ4w00X8e1CVBu8g3IX6XX6Z9yhSMQR98REAkzjrX209mUDe0vQNT91zx0SumXdj
FZ7FyBkNa4LRTsd+3NnCGoiW35jprBD4HTkxnz2FSenYbTJbC8dpOLxhNq9+Zv5P
A+Q7mPZ4jLf/HxLQrdxxrHz1U1hnmTdvAK5YjLZpynlnxbtqRjGM6tF5SvX8mYLY
Ro7xKd8C9WJrsz013n+70A9YCZ/t4K4Oynve7lrMbDHLTekYd14RXfivE0nKF580
B5rY7ln0CM0+qi+XySR93ZmIF/fuUIovyKj1kHVRk0IvTU6q2J6o7L9QZPdf/P21
cYoYSbgqGCtMxJ+oFn2/43CVsJ2y7Gx3dhdm0k8DLX95aQwBQ5O4m6B0rbCpPHTp
AoFr/4qKqX1WgBVzEkI9Gub2t1sfzZMiP/s5sD+HmrXF+WegLCSiajxXlORyaq7g
2yAzSjtj9BWX3PRsBU78/LyAyH19yFmNKWJqg2hGtEnMneVsSOOEUjApWsG0VMWN
EXrof+51IyU6l/PzrwKdNsPfMc9YuCoe9lDzhXkCRLO6/9tSVG3SLdBNmD9GsyxC
rqrrhEjPwXHUfl/8ie1yljgkRZlZqxr6UhiNvdKGhNL0UirC0aVyvVw/i//4U5jE
VvRNW7TDAUiXe27GI0ed1ZbXVcCoXc69Wv/IO+zl2kC28orNVzW3OAbq0g4UjuB1
bIaDUv7iPP8lvXcTTzbZA/GYAe9FRbiiH11Iail+qtdku1kHp9ovkbzpQzBR4hUx
UqwExp9r0tobnRcYUn4EvhXBChBO/3xm7JQPAl7VbLMqoacrt76vwHepkZVH38G9
/Ms0IOcJbvANgbI4yiePXNGn02oqfrvgFisWyIgRhJxkbvFVr4+/++SM/l3xJu5V
KhFn2wSIUS2JlLBfW1TN1eucW/408ooidbul+TrrtuQLNRvdFkThVxKdkADPnuq+
VIeslk3o89CG9PexinkvPyOuna3mDHal0YBYkAV+1WUq27Z6kpyStk88k2YgHP2m
1YB0HJT6IYeXhvQEGBzl/wCzy687Q4XaaslrUVoUaIGL6EncLm7E09QDbhNw7+cM
uLXd5yMuh9B2FKWzxvp/ArKJ4bZrUo5xdz22qIxN5DElE7RdW3saE2B2a2fxG35U
Gd7vw4Npw6Q2e9wVes8gUE6yUhiab1eYDsh3iEynfRcCdqmeGvCQE5LJ9aYEc3Bk
o5qHvmicvPuwr/0JYu36bXd1baz+NpkPCxIqNzYjdPIazn83CHORmQCBmnDeoEbA
KR19P4tqj9ZIGQauuZplYVoJUqyRQO1RDrzNXF1YTvk9YfQK0FDBP8/mD9EWKA6G
hp2dAo7rwpGy6UayXRfoDZ0vZEzBhNtdqS6WvOM/wd2VwMB6nlESaj+Fvdrv0siq
aJ+P1XpSocFHJcUAl7/IFOg4Ezi1kHxWdK9QqwSMd/gyyWTfd7nW3skDEsCQjmuc
UDb/nLkFFTixoeC9JbznpWWgEm3jPwb5VnsHQ1NGbdv2BdOIvuwdQNTefy5tTu4g
Xq2iJ/O4/sYzvWLKiLeri4wwPiL7DlkpiBQtP+SqC3IDrzNt/ncrlL3C2/R9pduq
MHKEbXeC3OH0LW3EXrNBGm3dD3eFQ3MBIvNZLQz6cQarTagXR+3utR8nXAar/cpa
Z65UrmY3hxWlaENT9oQwjsG8wb1NIfKPShPHBBUxNa6xIuLr7z1TYql0CIxHKDDM
cNC0yf+OQPdTFuIwH1xL+Sjt0asaD35e0LsI/6biWqPu2hhqxlTMGJ2HRxfrboxa
s/E/IYY+rW+1kCoTDTqlkYh3txuc50P7s+RQLHthajjTtt2HYsoHi0KYNsMfeg9W
XK9pZsrhulnBClJFuIoPUXd8i7F0bFE2VJxaRhjkWKSSf9kT4tA6iYijf5S08jue
GYozRyj3YRIcBNQyfHfgg7S3gO/WGyoWQ5tjdg391oUvdTr33kY1hC99dhLrYNRb
5xNPIQCFJvJOn6vqqKZpwH+dIePDTr9Y8TTxHUxVg67EXqh/Hyw6VRbe8BZdZCHy
gUiplgexXSX3fzwPtyCa/B/EdR7u1QbF/7R1KTMmMJ/uLVskcA3TzK7nYmNreqxg
djioZ5mXPzq5ltg0jS0Wkeqqi+miEkWu6/PSRdG/25TOxUaGsced6NafN6AVcz9Z
Tm3iBcLCiujn6qLnjG2m8MnQtkzfogyCfcxc1+WJ8mm7bcdTpxMPoEbgVtAU1Bq0
sYOUfwiIZ6dnPLKLNn4Uqp4iQJ210BCkxoP0YpVh4WKmXTMlBbQkpZLiyZNs2Cg0
WBzCz0z/zMJub5dJ0hsHawneFZm49nXXEqMHiGDPSbxNsHWinP6N7/97HU5WvJ/Q
XAq2bIRIpTGadY8TuorG6vncSmduhjQ+D446VzEeaVZIUHiIXInOrmQEVoJMQpE3
UgIfGbpK9+8zb050KbDHmcAtjYZ7IcCZ3EC9IKOcqw+pv8Sv05PfEy8ipZdDw+TG
cs25PYqWYpueSF7pGcEdLeXNaNgyeslAwkQK/myAXdbmtc0xlFGhVBir2ybw9+6n
9LrlUNn/vCJTBd4zn7OE2Q+LTbWCeLnhft//DWiaYYZNR8RtKPFsc/8rpHZ4+KQ8
N2vSZkCL+lN3I4c83Np4akIpfa2tP1mJaO3s2/OyMm5/2h1g8IU7/h1eSsuieDbo
xAy38BnEEIoezOegHxs663P/mTQ9rwHY4lw+IWdqO8jjiMGLH7rDoEsJgeL8Kgcv
3h8Kbuf6itjO75W2tbhX77/p6foUNW/EQLMf4frSrXuKctL+e9o6Bixxngd6yG5r
R7ZscczBSF1gFhyhVZi401wp7THa9dmpF2EwOmDDpgltOMjbN/yYXg4hfpQqfK6Y
YCgnoJ2bbx/ZxZZLg81ETVoeFTlWeuJH++cDNN66x81OR5NZ6gKlNgb7ntAEMOU8
8EYQWc6OPaZB6c0MyaS3VMBurWpa+N11ifpYjC/hnk9JXlGZNhZWEf/SiRgg/bk9
SscksGJdbQXqeZ/EeLFI3Ihh+Yekoohz2oEVKJWOSMuEweiCEGbdVKrwnyGZ5v5E
w8sjv/qdUSEk16MmpgoASbVG9b11ziZweFGnFbzOFvR968clNDw/g1MV6zhRjUFP
iM69yQRfNZpXVyXgpYmPldTWBRFDvl3ayvHTXBM9COl1l70J2iXW5L+TrV++/p5z
5iGvRKHmDUcVlHnGlVTFHsTWEppI8Oz0ok0C8G5TjkbSf7TjKhqjbfE/A+XmTdZc
FmnQSIqcfnAWfNsQU5FMGbLpuiDTLqTCOuDZD12D7z76mgP2UJlFle/omRuJJP+g
cH4bng/FFT2yRXsV4KBj04fjmCJIlIQSuH05BVpEulok40o7y/FibLeN/oxWBo9k
ZjTSthLu7uEuva17JkeEp0UCcamQu6IvhqSceSFSb0cy1NtqBE/zDbZ88TEVqVGO
kzHXgZ4pJf2Mm4TFlvqmsN2pWTa4hyrxzQm/O5XfrtACbLuiOKSC/YaohtCrUcmI
OSY006AKAMwAfuAUxeqPWg/pNPOXZDhFw8LXJYyq+SV/ak22P6Vri8Jl+X8afZLI
Q9sQpe6KPn5HKjzX3kpL0MwATewVebBME+3DL33/tmeqVkZON3eG3mpI04LwkyWY
qp8j/fSuWC8PE254Zgw/Ai7Y+dWg67LccWnSCwhuAHrZBqHtkqc3fgRj42t+ic+o
HfNGSgBDJGxABiFpJT9srQZE5Ba+W1p7ktrT4IDV/3NTBemIGUiy4t7LHcamUN25
+XVmLoblucJkpFcscqqqtE5p85Jm67oS+t758i/vkCPKH5bfaxYFiV7H1oUHGBXf
Os2Kt7I6EPKYYLMiYkYFGJOaNkzxkU8ToOg8NGby0ks2ThTsw0Z+k6j04W6sxIAA
GTDoljhvyd4X8kluj98HF3SXI7LqNCVMfkK6Ra1U7B+c+taB6c8JTvDYLySU5c0p
4WU+4+EgvH6r+qZ5aJ5ICwFuOFgGK07Melg3nM4g3vFtvc+hW3My6MSl6SfBLJtl
uOJ9+jJV6mBLJo5htxsJ8DGGXWhk4v2s1RIx4rQARl7jmJ5MFR+WJ0s8GvTm6Gh6
YR8oLhOCedSeLn5hKXK0ExYn0h9fuhg9imQCD47wxDcHts6WTwoln4JkYzteB6bC
6AnKMo2qr85f9/lQC/ehLBlXQfGDxk3cqhOAZroXufgYamV0+fDPE4VGb69xN0aH
LYZ2nxk6p0b1ruf4dpJHLJtQy5jvz98oiT6RmmWA/57tZ4CFhNMGW+M2Wfnn2IDr
K4bdhaB0v6BKKsuZpuI2+6UNyZ+HbeBoa2RRHZT+SParwpopnlxNj4uFNzbt3sPX
xK8DEGMWAuiOY//I0tq4820dd0Ve4R0TKWomsYFiMZlB4gIQEjWQkAnpgT+/lGN4
dj6/W38Y6WepKSUjUzP00Z//iU9stWf81Bk8EseJUCLJjY6/+jEhAfS6FERaYemU
O421O/WIIxNjOdUIav8AsXyQ0xejpaCNwgVyQnX4ivwS6m8l+8CSJnBbihwVwc31
htnviMTRg8W1iSyUH35PuNhom+1r3mPX3TF29x76YBz6+9C1cF6/qJrFROrYLx3X
f1BX0d5BlTdVCM15P4631PKjTo+0bYPiAY98+zedZME0DKwKbl2S2dK4yjLwVQZP
fe304Wq/gJIL8eP9z40P7tWQlWwpaYJie2ocXF1q74IWQSQYTRzHPq6YothKvA5F
Ka/6lOY+gWx8e6LIwbAAHJJQ1jDYMsxlE6MbueSgNBmSQ89RnjUoxtPQ+vwBHoeN
sA/SKvGu6FupNfcImXdqjH9oWffbM9NQQ5H4dCT1Zq4RhOYL5UPXmEjM6KOSwGe9
GK8o3Z3g1ZwLFL02YCcgE7TqXyZ6aseVRxsgxn/cZvt6onKeZExzWec22xuOcxM1
U6piuNOILg//uTerlEzJGN7mU4qJz6RhuSCu5MKgiztebdlz7aWHZ/UYJvxhpYS4
bBTwEfDgfDg6HK51SrgfHiGGYqdBOHqg+pQ6mbTX8SiO6eroS+OcRrTNSb8kAKpp
VeVARjOhE3w1l12Tqm0E13tKC40F75GyrtDcV13lKcwB5NQHjvTEoDsS3hCJH1o7
Ur0wAITnHOM6YD7az1+o/7zckazGxZ7mBAlyy/Pqzrx9dSm56nQNbzkmFywxEBXf
LpBLpxjnQZIvTKwZrDko+NdsPIUziPx4yMiY3LIAaPLxOYN4Oxy5vV+LBgHd99fh
Tlb4IvJS/x9Lp9clxihNopfF3cYETYnqjB98RJsyFmcHg1aidh/VPLsBojimHU3S
GZsYkcdBc/ZX8yMQlnb9H9mI8efcMYnsaFNd88TdY1R7FI8EhNwqap/dmUocp+Ap
x5vBQUjmi6kbqGy71R+Q3oi0deUokKMbSfeQJyB7rYbXZ7mAP1ZvHcw8RT5SAjQF
+K9u4au8gFy6nHYr5Sqzkm/YUmc5SeH9CK4uparC0Qu7fUrVMa3Cq1yfW6oc/BHl
X9fEuM1j9AWEyrOb35YeBNTg2AloCYp2puwiqEg/YRLXvXLVgieLJ598aE2lAzuz
6DbCO2rXMUxv/gagr8EXx0MtA35kNty6/L+t4+lCB1tmwDYrFfhwQHzICBcc1Y2I
nRau7tMP/2eRFW0pKIv+LAFDtt8uDTHddSt6S9rfV40PWWiqLObKKSBW2fUoTwvM
XWO0Lg1t9bgfxFRgRZmn2QyGEywl/xn25C62o2HVnKIVCLuqLjiu0uvndwMgdqBb
yTKG38teqCVUTd95Hs/EWxJlwYvK0fQiDckPbji5A/tsAZ324/L7nIjFUH5P/heq
9pul+ZkPHGLYZrBCyS97YS+prxLd8TMrp/uZ/PYtrPziTqIlRUWF2k35DqeFmWtw
toYk3h7C6SFXwHSKJbxuIJKf/AkaXAdwD6iyD0CLbPwwR7vcBSB+FX0a5OY4pe+S
o4IHYKI6kFXl4/APFAZd3Wch9gWz82IqIRj/VUdXMeTfCHPuzSaL8lzPYzr3wtz6
d0LvRGzWNUv/fYmQTEriWZyHqA+7Z05/dN3i6QvmASd3LUBV3pQEHBjc1zkXvJjT
iwYYLnF7LL9zBE3CCS8BDmggUhEFuXbOKioiwdlZt4Y6gfqLPnRvs6Bt3RXHs8h2
ZPzU85kGSSGzJYZewKk+r4Vmx+C0RCl56B2PBQnlGPi54S6xc0j4liWsjZwSfbXw
nIGePltruaBfSIyg2WfoP9QprRtfNSHEL8RPbC/xAPkrvN1FKDV64im7Dwzljju7
5Mb7DVksc/jJ3LVOQVzwDoatrOcD6ock06UDqU2n5j0/uJlAwcbVl4uLyeTJRE14
Mn1tmVnKh4IdL4GJIlSaPFHyb0K7v8IKEP7nDTmOClSoWf90yjm+LZM6pHoxyd5y
KBkXMCC9qs3kTk4oygNs78t35brEPrsEeYKgu0aOIFOSXoXS6GuXTr2pt/6BMw7m
qF1vi6New/BtsEThQZNUQ+071YDZWz6L8z8QG2oiPbPGXpQJf9ERvv8YkbB8kk6z
+exgUJKkVoZgmEIJHihqYb0wh1bcRkHcPNpxpb/0fUtQEqzr32iVZkeZuyA7ErOP
UYcBgEfdNEoPDoMBEg+VYNSmnVLm0l4ubZFMXeTbyYdrve/KWvX4orCPYE5utYRL
cP+0Weib6OM0zjLUKDoc+guNQz1eAOJEq3y+Kuho9FNK9k7CvJsORhttl9Q5mVLN
zbad+xJaRL/a26gCU3EhTB5h2YMiIWKIDFp3fvP6uqJtpkyfyXw24mchjyilRMmn
mxZMIHc4ClOY+KkPaiIyXEpJ11WDzftfI//vm0PZIC5UetPfKWYjRV7+DuqtqL8V
jfBB0b6LPEtLFOfXOzHty8j59OR/ZTS5pBPxDSEzwOPkzFdWqpwCL6NvTrmUg13+
JYIT1Fth+grmUn3Depm9A7SCw8H6ocNno2vQr1Jg79GUefKPy7stABgKK7z8STls
nk8o2cd5MhZBATKTIsJ3EQnyOI5Sfe/dM/kgSiRI3fJgYCmlWD46hT+VDAy27KKr
atBZXivnECvXxRsnN74d4W5RFA9f+pRJ0okUddpTcyo5Ug/CsHtp5rIPHTTdzeIu
3xPHIgWmseX+4Q1Rc6ZOTTs5cQiPXQ7YI25ev9GTo1WTFVDRF9AT/7jhFGeHXNF4
Nbj9STxfehvNAEW9n3F8Dmyp/BtKXgsCPnhtOrE2nBaKChZIVRVG2rhTcDXcuoMc
6zUUmPfEDFxiDsc8S94pAiZIb4VwmB4ZrO9bm/VrzrgQcu2mk/rN9tEgmQ4k6GR0
Xjvg3udwATN9Nymf7rjKkQNN/o1vEgHT2yvt7IDxhGYDtEYXe2bKTgWqvqOeczYb
jOWWuErJ1lSmOVL5gm8ZXs1X4NbiCCbLqT9/8AZ0V2buqDxGkZ2lIx3901QwRiC6
rvRzXJkdOUbtqdGOMORyR5iCfvfCY/vtUaTh3eDczCbgoGhekHqUiszR8hFbvSH7
XCAEJqbs8Iis0qPApMbguv3LXAXzezyTxhgJau5PsQxyfej7xXYA2xTpiOuTyA6L
ffdD46+WGKHHtTGIKMANStAMlOhdqPdTvBj9G2fEH7MjgcpmoMWz1RLCCypuIgMg
rtARo5FWBv/4P+tRZHb4oF+JXwxPGvhA073kEcLHejhtZ3bJdWvWg/A5qKN0Gf9p
MKDI+L6Q1yUnGKL8x+M26mjHhoWA7pQJf8RWHVJqhGQV+VAU1aeSxF4TCCBUcKra
yoFZ60p0ZQFQ4g0Ovwpk/ZcjdYy6pj1XF4PvZ1CvpCVw1TwrFzvmtTd1NJNA1W22
259IAQzw2CHaWhoVmxTzg5xjUfa7RQZDZLRpj5F7fn9++DpF25pqfwR9OB5Bs9hx
l/cYCk/DgH+YRQk+ttCbLxQznrm0+EfOlA9dEhBEWvFrVypu0PP5kQD1PDuvZzhR
4FeKnHD23BVZlN2l+Oaf/irUNxc5IC6L8efRudQYwf9ZsrsE5oy5oq274aOIM/vv
HjZIYigPHhWYdcYlGQFfDKf4SMXS3JBXwH5F1vv9Li9w3pb4NTQ+CS1FF8XBhRXt
/kliyjZzs81t4hWEux0MfAOEPniS3ZqUYZ93yRnBECZ0bcZh52pZEH1kM8Y9BKnQ
Ry3hLjl17EYctfSWE7G3HbdaqezA0cSC/vF6nWQLgB5CKi9VLf1UVjvpcWQur2s6
BSkr+vAiK9h1o7mb+2xslqFVG0FE2KZ2X59y3v5c1lXECnc1H1jHRQqVa/Ow723T
WgNa1NdPmzMbjl5/DcnC4/JVy4ntaXfi0cdDCuz/I1TlcfcIY6fCKXPyR7PZWIfj
ZNKQwFXPSSPQgnXNJL3xC/8/CBgEB0BbFbupMVb4v+LSTaWjGlH+uGDGuZPc/En2
q0xSF0k3GoH7GFZBWhPi/9GQJG+zA0tgSskk09LcQ5rBmKcEEdSosWRIo9ukiiSw
/bHlZ7nw9M0jbU/CE6afM6/zvydh7Gu+SS5sWVU6kHQiouQyo4r7iehkztXpIoPm
LVGBI9op5gi3FvXykX8GCtOIZ3PaWlQ1C3nmDjk7Od2dymRFjzkAT7TWpxK5CxMR
sIbxG9S9HPPsG9ELaWHEk9d/7fP431oCgBDl6OgRygOtP/FhsqXNRoI9khWk9kqG
YaVBhRR+KgSd2qGW3OXhSwHAd10Ce8ApGriT2xn8hgYjYKGAgRNPpz7EgId+CfNF
jsiJ+usBoHTJ+AWx4UdQN1fRJXnoHBInKmuOBoqLfEBISYwC7x1cbEKmH336A9xA
U+rGPBAYFei70ozsWHiGVL68hY5lC1372p23TroneQtWiUYHEHryJwXkBt0rz65P
ajqNj74u21xaBlWDzeQvSuUu1+ltk2tO4YtPg/lW24WpYW9ibx8HXZKOh4p+4wnd
Uij8Q+GxClKEvlobGnljN0oSZy1ZqD0fSAU5ZFx3UrKAIT52QG84e6kRX6GjqnM6
y5xo0eIUXn0NQXgS2JeYetWP//eLYHiXBbrp3IPj8hvf2Yk2lZdXsZd1kKvbn8hp
JjEq5nKujqhO8IPmqhID7ieePHfT92mSorM/FX4bkH+E4L0pZ5R3KQ6CwMnG3k9j
5Isj6HnUjnEkDTTvY59ASeGn+ATgJVPQPbXLDMdB0nGCLswNNNQQT3e3zM/mn1pD
qafhAI5mm1spPijliiMJ31xNtFVxT5ft0bA+42Ki7+Vy0tcyuAeA3YUFrf4jAh7T
D5qptF4rkCa16M8YNVOCkh+t9us3nftf1/7BqwbB50oZ3HwepD9fujX+r69qxyAQ
DUwY3Y0D6ifXx4q7uFp6QBZpq1/MsOD4HEThMTKPDHJDvw9WTd/NO395Dd+A6iNn
T9Fhlw7zAemkXxeGC4qyeY9kFt7xoDdHo5i3U515ehbuvVRaP1ANzynAjCLNKcp1
b/ji6bl2PfrkbKdRyZqkalUB1BnbtDHpIGI3cm8Pi1sZQdZgdUe6IRFTVOZtUth6
qRLjrZlqxR9hjY5YCrVFI2C04a6X+m0+5XS9pPizlTdfhRo8LfR/ywOWiG4k2d/+
onDOlaMPWI5Y7xOTm+FowBslyNEWVSbtyPhY70mozQHTNi/d1no/D9cHuDc7uiEP
IFCOO9qymjnspH4lfBaqaYewS+0fjG5dPWVn/X4lKAyQ1gEAbsnRx7N9knakFQpn
FzAM1pYXlFTgJKteuRbCb1lL3x99hrsWMitMEXowUaXTNTtu17dwFUSfFkMY9mEu
2qYoZCEGQDeEt5tmfGOP6YA6svHu3YWZLpA1mA8R7ew1B9wFphDAvxj4VjMBkfS6
CbUchmCfosqDLObVysOWCztMBYCJpNGWKA3gGDNCD2Ce2UWccFnoEP5/VIPr0c+C
stCd6tsj6bHwAlZ5tTS2JagGbTwEDfogHaIJ480pmYcNkNGQGNVZi973SGIM5nkw
nQ3yYDOQK2YVSBajiAs2DMF/C35pegYRl7VlkR7X/jHIGW0zqhZm/lU52SRbetsp
0LbOo/YMTZiol0CVv8IKgJvq1IgfVRpFpMd+JvRJr4OddZO9zz3Oftfc2HvtmB2q
EURSK/ef95B0ePA/HGB5RVNreB7hoDreMGsUSPNkh7FsVZoE00PXoNCBZtXyHb++
FUUE9H7Gbj8PVGILNkyi+WcLCXzyjEAeAN/hZ95LgNUyOnHhujU/eNyZncWOdQ+u
Sq86PFqNBEIUH/fRrdvYKx/bZ2lAkbQiifsgAOvQMd7nHjgyzkGTfVCSKoZMddUm
szCRjGO6Tp8G3cXOJL72UmciR4ePVg6d0CTMuoKZfYJRJlMLBHoLu3lf89qIP2go
YvJo0urLCBfGStb3HrK3mOnTNCn31aoxU9iMaEmDIyaVK/BduTuHg2jAF55s0poc
J7Btlcm5Oa4VPgfSz+pawsUDe6yGfHz/LKFPGEejIRwDVx8SGWq/ucIrT2ODbeNE
RaplpMl7rZgjDYTAflRE5Hv5GD3dpiuqxLsxI7CbaEhvqorLkj9Hn6PfjADODtvd
mJxRiErAU4LNsLt9pGJqXOXgaMaQTdEIeHZifFB+NIulHD+xUamqCRKtkzT+hXTh
xGKQlyXoA43TNZzKYWVmwPyXmDDRS4MPbhZBqrO46WMKQCVAtZp2C2xOChIS/t3E
jO1DAcrL06SPm6VkAdrDZUqyT7TDl6de+IKSrhLR4dbzb1by7lAMkrXRmWAEn6DU
gAmdL6H+ZBscaPTsisqsTzQbK3DIK2I8x6mIMxb0ch+/VWU6lncuoN0oIH9KVWrs
AtXGLHwdH7by2gFfDe7qXouiHdzNgPpaJeQMh2ySHussbq67KUMCwXXRjbFM3Ji2
6S5mMtJ3WriCOXEcVzF9ZmRO7qkC8cTvt25uyJu5QuiLe7/wDPx7G8sqQ5PqXYal
CT7SS5p1D8nsSH6aTaOjAhvihquJObLMxenSg81h/T/2ibI7WTVKEuGV+PdoB9TE
nn+i/YKavyI6XYT1+bJBFbPtcDHSIP6gBfjPZ56a7eglA06Klwx4ytvOHO2nw6XX
bxowHs5dvAcBUaCSWGVdpeQgd1r0fYQ6xwjMORDzEHa0cTS4X4j640aY5kh2lIoF
sR+cpPeDkpebrj3ZFzIEv72POxzCigSTLwHgxth0+R65IfKqIhUfSyT0DCLUI+Sh
PfX0SSCH5x7SB8rqqOjBXOFRH6bzPKZEWlNrmltNbyf765pLj07zGrUv/r4gPk/f
+jWCcTztDe3NLiv/ovfUi175da8Kgqdxcwed30Wi+6RbgwhGuk133ZRc66LHDQFp
ahSJJVCXUzlxCXfv5+b6FAiVMjrDar0h1f3QplbYxEfJs9o7rQ/TxRdFqYG8Kjyq
zJDaUprj7OOAx8vte4nxgIYAvi4EiK1D/7yPE0wKxzA8uFM5QbXv9m3JIpX+zE9a
uxSndVBVJvjaDN6fStetQDzozZG6/vbnGTtTegwNCFdZUrEL+GeA1Iz2ke6rxuhg
XxTYW/Z7UM3ngAjDnl9arRAGiOTbKdvJzzKz7IalqyNTaaWJmWfrKoCkUW3j1Ciu
J2nSoCUptDiBy9zV85sGgfShRN5EtjVzzcrG43KeU0mZSvIRwhqGR5Azku88a4NT
zXUBVDzAQP1RPcnfzIpUhj7x5OQTmFzBg7doHP+c/sXjGTwF/wiKK5Rc80oL0G3u
rSTZ/fpSt+YV8b4VCCMJwkqHXsGfI13EhQJPO7orfrSUX/zdZBc5rtBp6/bzPeOB
BN3g1hBwqO8SeMcuM3JUqMxxlJ1lZdJ9UMr9hvtB21T9FfTwwF9alPAG31aCAc6G
mGuKeKZlZ+qATy9NRSXCcEy/+OyfkRR8Bdyj5Z1R4PvDYaZ4FVIVq/tVQfe0tnYI
NXGZEFZwGWDKmZViAEExF6Rc91g9f+8HE0qjt1ns97D20EDx/WEXrFQmw9+lMh4n
uTyXNQZlLcyu4lejOPg1l1JvrvBZ8NzevdJaxF5xfKCRSkREclnnXQzqq1degcMF
3oZi3wOJBkGIzX3gmQV5MQPACDTUp4XyA5hj+obsIzV0kSJm4/DqoSPNAxEb2Vxq
Ki40BBs05uflUjNMoB7lMiHZguiYc8hyhY999zfXSGnZEiy8uuyW5+0SRo4McauW
KhXyaNwdHXSy9hNQKpmnqZibN7x1KrR9ij3rpucEjUn1X+da3mKmFb5I0pbUnaXh
Ax7qDr/1gtEuWFou4UW0yItzfTzXVvVwhbc354gdJO2pjGSnEbppOd2GmLlQrhgB
ErcnVzdfQ4NAIDHdvuxHesq3KqsyByJMpaqI9eh9qYioC50XcBlzQ/hsU3frN0Nw
CARRu0dO94oiRgeI5AEV2bWofwTdopmusd+nBVz2DfiMRd6jRYquQcqeg2tOLTa9
h6F7Sp2dYzVA2ly170wedZcvwS52hBWmcfwdxIyJmfbdnGOV2Yw8wz/K/7EYxxGR
XK9JFg5iglilDBEHy+jpVGtxgW4ev9nfHvq5x7leOjQs9g9YgGpRtHYr6d5jyqVV
IOlYUMn+e11yR6OQgg/wdo6u9yLJm7I3fEGB9VwwlPCd8ehlN/lyv0pAZr4IVbcI
OwG7KWo5drbjVpr6C/bDYSaz9d95LzDrwim7BfYeoi1ZejtCkB0wTxj4uAHEAlMj
4og6P36faiUD43m40X/YDJBWavOfbM5VwozDHqDEGGJOLjTQ4qzJ7QTc1s+YdbU/
wmBU5W+6ePSrWi5pOqRAI46nWsU3Qzmo/8YLPxqKWISEfb/TIqtGgRK+ed4AKMvG
OiDbnbDjsJmuFTI2Z3OHWn3KFUKyb1QcN2/UmJ1pXxiWVBUZ47laYf85+4cDepUi
RsC0ACgz7vq/pQeoc9bHQp9dM5UmmKsb2fFZety5DovMhQDo6qXV6wmsY4SMUvIL
7JrGvIRtCmuy7Q+m/jdnpnNll/YIFAwzTVWLGB7zHij2R5OuGBh0TygMrRvpsWF8
Jjsh/tldaBQy3tmPeKT4npr7Q0o9bhF11xVezPX4Bl7LZhBzMcK+vvfWboSXFEeQ
JwbczeZfa2xufIi3UyrtwyHokuEu2/nJvPgIA2J8GLjiv1tx00zrmHv+0FOB2rtn
uq0h36BZ5LCt1/pniKLrra4NeBmGtZkZ9FpxYJvPFV7XZBNgNxtErsEa0v/LCXuG
B8uvcFsCuP0LgHq/Uoyi6DWCpmVVJhsVOme2atHyBkBt5bHKTFBne3D4u3lN/9eq
rLDqZ2rzQQtWE8VM1gJO2FLVylvhFpCJert6e0bGy+7L3eiMdsA+ZSPAmc4dGbBW
0PQXN1XPPGTEVJy0OdCVVj+zDpt83r7P9e4RzboVYqfnJRwj/CzF0usNELNezWU6
sJ50c7kF6awh75NVJ2Ta5ACXBzrGpf3KMwC8L/P+Q2okFsEe7q52w+x46SP5wkLz
7KA08Sy9asXmFgCFADaNs9Q0RXEatwgv9dntalQ4aE4JpA+IO5cn6hNo5DqJI9uw
j/H7BB3JMZbPFFnqcl0cqfDeW0lYGOHyYke/YMcCgt8UkWzz6ax3iUib6iSrcA8p
j3E4q+/omjkTL8gJJl4BAni+LbthJOnPMELSN0D223vU9CjoV/DGmBahC1mU1dY4
zLXxV4Z71UJKNKEg8BXWtDAnUOc5rIk9usnpMA/pETbJDA7eE92UThwCL+xikw2z
XJ8Z+8z5Rn/VqUCQXWDXHPmjFFtD8IZxAB1scAV+iWzDXRb88h+vpBbkGbLZSiz3
DUFWmyTY7HUvehTZIwtR0Gl0IyGQ3SJqYNoHT/a8gom3xPPPBcehTvYoSB2o8s9C
OEPYFB2/l9V23q4P7+4kFU9TOohXb0FDQHSXy/1yFO9chReEUjxXGOgGBWMyNW5k
fSQKdnOqaDLZkbmrEmgAl3xil4uVoLkQTi+1hsNtGBTsy/ZG2lm0zm4j4zEZFRLI
Lu+4dQAfs1lGXWPYzN0dT2Q2nWNoAsx440sVSTzSYOAs8lZ2K/v2Pn/DHsZY1Pno
Cn/0RSo66xymsYf4hSlwDUH5qxs5JUmIGnN31iu6gZUEthjvM2xOl7g4jlMwH7xH
N+dp45XQhuH2/tdG6KAWEO59PunX8sJfsO8t9ror6wgxj8wAEbTUDiipLX1RRWYD
JdDjEn7TorZoiBeCipQLEwBT84gXavh9/PfJU46/+fBabEeOpxzuFLYyXJ9V1VW/
6crwuocfp4FTOc+TwlJGCn2qz4PY/43EeyEC7s+I4zjmmbRynqK4cs3W3Zzznl5N
8M59BiuaB5fHabe4R33mNo0GOvyUiLUvdgoKEA4a6EEqN4rTEcCga+5dgy3lA8dY
LtLjrlJDLbT7NuUyA/Dll+DAnSAc3gAVCtXO/lkFd3ZOTXfsZFmaUp9HBRUFYNuq
zabPUoQo/kLrk3181EzoXCjeM3tiC09oNt5mM8cm9eNfatd/X6uT7ZcH5hBlGFUy
cpBXKTZNhU5NfzUqDQWxQrPw476U3jlBOb3SB168vr0frNVBUJAa3ZRvoBI9Ra1s
/m25CJs2icudqNdTJWfyopVsYIddmh5G0rWlascYVJm4Rn46zt19NnsKV3YdfmT2
5gbtedUyUJRfIsR8IGRDZGDSVyT62ONnUhI/4baIJ8+sHo2ysgOcmdNDy35mBnoC
p0r92qUJNls6mTFm93yto2NvAb2x0iouabtvhLaiX+hzPBP/UmEu2H0IKrzp4pRb
iBPkiUWUGKdKxmYfUfGuw4qEnTBD0ZVdpSrl7zF06klK5i3dDnc6+U2X0bjAadPi
kksK0QUp2OguW/6bn93LO5LRaJXItEw0SBGEiXmiAtMVyFO1o9LSGzxskS4r+7RG
Oh/14NjDIrsfGUay/4srvh8xFKAz6oLZGrivTgj65aozd02fhNzI7gAwgzDwS32T
8QL6Ht36SgoI7Aib26ZfFjzUx3R9eU6TUM0QCprAWbrGZlO1eVCNnTwdd32eEnFz
jlHZCLnIgZ/KGH3xGgRTZTfWpPLJTfPkX/zLc6ZZS/vv5vCXeYSaZZhp9q8RliVc
SOnVfA/dm5R+jUc6q143g4xGh8mRELKwBN4nLvWzeww4pk5xp4VXU//7a6yz+aBs
Zj/wBQOcTkxHxES4H7VZSlQxCig/tf5vyhEs9cAC1+7MPBb9wz7rWnX8gmRmqJ/s
Wwd4k77LN3gKfDpc8yiPEldXKTXSUHahUCHY0/4ZIxHC7EnJY82ZrPy1yORJGnMA
54RiT2SfRvN0LnLxOBv5nBt6vsveCI6IaK8Am3X8j0/a58BEbtUoEJsN5m6DU/jq
ImkRnZzdbd1sEtQpgcPnyqkDvMkRWRnb/SfWECpIoj0P2E18LjnrdJ80xUNK6WeO
1C+xoNUUs5ZtfF02SvnpgdK4vA1/ZdE0N33NHpQ6m/aoqwCf7tEHRIgLlMzhxu9Z
HI5qdsd1wBByZwK9dKDOzvuTHLse9jHVORLETh2IBvqL7ZzyUibhVuyXHSwzMtoq
TYyrw0jR50ZxQZm4bbdC0D8wM9/WJxty/VLE5DDJJ40VSl1Ps9fi2FWnWyB9pLeC
ECIaTeguyg4Zhm2qmbbc7pjybNEkzd0wMduKGkcK5+e1DP0aNKgZ6SfA98+XPtDB
LSw0IoC92FUeJ4w2K+c52R/NZ7odTAlneoJAEY3cINR9ufpInSO86/qsW49hnU1e
PmxsG1eXrQvfNo9vhbdZSS2/50mvmwaf89S/exQ1McDQto/6wqLIXhY5lYVZ54V1
8jGgRWuqmh+Svr6/KN+kq1k6tJiGGNCoCu3m5gQU3CHLqiw3Ra0qoQf908pT0oyH
f5qN0EHKswXyEIjFGd3rkGudNMQG9BBLckzmfzeHgguZbLJiqO1ncTr1WkU0muPG
6i9EGxe/pqBApozw+e3454Am1DtCzs6CXWiw8MH3NBd2pN/1y+m4tHBAn/kYI9ho
g3xJ9eAICpJG+Nk+qlavN+GEtR849PzKqx1jY41fL5JST7/BtJCtMSGStAJevbHj
AtQHHOuii1ml2S0hTU/kF+wktNvgn3EXnkImZsh0Vt7SP1xXMcq+cRYd7c7BpYxe
sKOVZexJIL1DN4DWpJb/n+zmLKGNzw7MZb39kt3i3K9Al5Z2wLarDL6MGT6Qy8OO
VxnpoyhhPkop6V+DoWGWfVZDw3Bdgux0Iq0/P0eBi8ChbAXLLbA5j6Hc0qSV3GMa
8BiWlrJVkeoUsopTGqoa0JqVV36/yJU6TY/7VxoSkvFGJ5/eTlNSKXHhC7RrDftC
nd56iOFEd/0ss6EGdDMdojyEdirbk1apE5+HRAR5ERJdpDH1FsuhtK02S6aKWZU9
9ZoFPy7uhSmZXlKedc4CZ4O1Q+JTVCMdGUeIEM4HB3H/68VCM8Eyk0A4Yt+8Te5N
e6t3gF7Y3flMC2eUh5OJaUhP2iVvHdfC3CAFgAiNqrNIII9v/a3aoPhPNOuK5V/z
NJh55hMlz5H4dCHJc2bwAzaxz3k+W+YgB5oWaqF2X+VApolz70ttwHY/4+Un9wAB
17T6bNkaJGJc3+NqT6st9aJi074egAvVNeUVU97wUqkSXuxPvVLZ4XTBWgH7ijlr
e0iQwsbbw15US/JQ7OmUMFTVK8VZoX/7FI+ynjKpAIOpE22VWZiCyZ3Qo4Byi8xr
29CzTPnWlw+4WSifyroPhWJQ+I/ud81MuL7P7OZscwc8MrQdMpCEMYLku1pOSPBF
v9/un12/FR0+VTeOK6R4OXdKrCiDgAh4jUQ+s7IoD0/Q17uf2wZncSNzvoHToNjj
p+7TGoIH18zlwigEwySohJAb+f2GBryat/xi1ybX+fvWinq1mudZDvLODNzQXdI6
ECdSZZqS+GaSdd9hE+ymFyfuEDDy6bWrsb0Q+WR9vekJ1lSZ2ocD0TsxXS7lHUs7
Wbq2pCYQtxukKuoxIff9jvANCsYntPLT0bytyqS7FsSq70qWpa1ENQc0KRNFzTkC
vAdUkuhjRzIOSf93jCQmvKuntnJ3Sr8lLhIfEv7GuOmYvY9H5RxD9p9XYY3avL9S
l/4Kmt1tcOIq5KNx0gkqUBBPZaRw8bsFyWumb7dlStdZkAvZ8QxKwhx2ZZNzTDcK
i4w6RYvRqooN4hxIwi4QcDewL+n5pE5QTyLS25EIbRI4y3xgHTje4b5IPtZSEqJ6
6zRkDlqOxU5HC+Hfo08Ji/QFb8OdQNEbeRWr1CdUOx0F0ReRbOkIozyG9zExiLvu
55aNITq+FZD9IRJswmjWWmzbaNVYn4hODqcXcOhMIzfvmUI8pubsgDoueAtIZMof
jiGWfTb4UqrWY50N+etUFAT0+LJSPY+e30HP0GjagmNsuMtXWPvgsed7sw53XVwg
xvG6nIOffutLdIxsOmw6l94IsrBbULc3BSNd4IuSWWoGHg4ZIwGyvQ2gaoHwdPbe
EonNoWXSOuugujHsrFZmAIqF7/EkJJIZX5edHxWMbD2Th7bW3TD5y+Au6xgpOCNT
SX+6qWseluqqgorMSjeZB/3gPj5B0YVoR0fgKFbo/6+meMJZK8U2T6Oz27NGdwyx
Sv5pfDlyeTqEmq9ZCuk916OdgU1BW1ijdm+EXt6/gQEsrERHW5VaoDRJjNx6OVLi
hUrGQHv5FuLutN0QtNyUDjOZGgvhqfA5b9s/D6DF+D6CH5LKCydyZT3WFCpbDWru
Swk+gdZtpC2XhL/eMN4Bk38oABKPt7B6PibIlY6lAsApX3kv8AQ999tCRY05DnpL
qNUSGgQrimLhqsE4ny8ybuYm4kGl2JFNg1/FX8SQqyUpFicB7z1Lr2vwf8KjlPOY
u7DIXWrgHN8Q4X5/S1Jpf5IUQqOLitcoNMoNRm8l830a/S788gYuOh21QRuc3mq+
WptzEnDgt/UYSdCTA761RXISSs9aVnrm5E6L1xmS8PHRB3auiglgeFkjmzOEODy3
MeZFSm3/n380cZVxEDJyV99wbNUHwjz5odS67kqRYL9CmcsaS8uJdKhRGVBKComi
NEjILDphz3i/rZ2jgdpBrD/dT5EGJqvzO/+72BxjSL8xRvr2yyl/lPmugJuL7KKL
7wHqPxqMFPH+dXPLxD9tM9BjjZhiqqGGW3g21fJUQz7+qfvj3xEDoJ3ODkRvN6Oz
sJ2llY9ryOyLFN9e1vKFaNGH2bI2Zfmrlq8V4n4V4RPkcMax1XvWUhfoz4ZAfDS1
fRUJXJzKftJ/KVROHISy1ELx64QSjD8CAW2kHviTFEa2nLMnPcjnXsi3n0URYwMK
smmuQTPAhZWwuaQdESCvQzfocxI+c4Cd3IBumORR8AQSx8BLaSBv6MZT56YZ0Wad
4smsJgp5/Ds4/jvaWWW7kiTi8nJ/zkpN53hBczmLLrwwL0a2aL6EiWuQ+HiwkSmU
W+EgOEbiWJYJDosQDfOyPfIrzVoKGvcU4EQYooA10mqlhISOD9E4Z9Nde9mWoCsN
1htR855sGikqLDjcpfHSPd6S4UFjiLx56Ynhp2YaCSRgwvnKFnLpRpPJE2fo6k5H
k/Pyw3fXaD6bAyQeNmwdC4DkD+u0F+s+pviIYH4WSA75fjXA8e8Q+8W0iJwESlCO
yY+rOi2HT6AokawdaFBb02/+5sSFH7BJZVK2jVUWFnd3vLDVC7hXisPCT8F9O176
bT3bwSIm98SZop7txIY/xleBPiyI5CeRmd6dzFeU8Z9VTw2NvBegJPOu7kCXSJ3S
k/JeYnOv+QYnNJFwDVC5Vxggp7IsTPdvFvfGnOoEGo24+L6rcBHnqJ7wN0IzBFX/
gy+DDDowpFddq6m+922yetinRD+QfEy6CLCIF/Mp9RGMDlhttlXc5atJgzgrCzdr
B8Yog2JsPy24Uvl6muOqZM/RVVI6Ot1+Xl/zFkwC2nggJ2FfKo6YpRVSJZN+r2aF
OIEH2GDTEzaGU91oSKG7jsSGt6MY0O4xMPcfdxewQaKQiYGw45AZFRou2XSrcCN7
X0L776wOSiAHLLLC/ZCBIK7++CPa52+HcbxXCj64gy6myMduTN6DFLiNjptEePFw
SoVgk6NARYpjoEz9bYljhcExOKgpAS75idKfWA0NqCvGe3vkFgnV+wJea+A1ened
spX5BLJSVSUQq9hs2bmrIFu+RO2xihHuMJuojbC55mWvWABv3ecdLePOlNa1a0gJ
SA+PQFR09rkAl0Pt8EMrMgfjl62TYirOByvjYUYC3UU9pvtlIcxJ69yDMrjQuISU
wvsJAPh2H82fF5nlNVGOQbO3efVeh+9yp/912ztgEshNkZGl3RRjga/LcLTbKl/f
9AL67ymtH0V/zgNg2KI9svqD4rfeCPK79hCmIwdxomAhR7a6cLSfRH0ccn8NSl1K
mvVL12IPZlowWm6lKy75o9B2/uJZHN5hh8c5uJ0YnKEvegdRl8tl7XH3XZ/7eeKm
CrgoCgM9CZpI7i9XW+vaY65o0QjsqQv1vYCE2czQo8lZWCnu6pwQdWKODaDflc4c
1OelAUw/P0cJxRIrukXsdfsWyZxEyWcoyGhupJyFHksM6yPBaSIcZhrxF85GcndI
/ltd+t9+8hYZ2jeSaAPOtbAGRi+bM0kG2YaDtRiCy3QZkP8coU4gV2jzbqP3EqVT
swterdG95fxoe0dBtbB1cI0gJe5l+wI29LKAgz0ZyU9c4Gy9zv8NIL93cU/KWYn4
t+v2O/WCK0ZeTGxlFoRum8YJemINbd+rWr+EKrVh5bz+vhr3XZTmfzGRD30f2X8D
1BWMVUheHEXGCL/zLhlv38mNpdyO5OMLaRGm85ac050CpjxfCJMl03dlpB60+Kq9
vXyPw/bWDlMXX+8dUVXwFKmEmoxKRNk1nLBlFr8VAVS3MoIn76tWgRRF81gH/vOh
Fee9hcVXR08E01v1MPmb+KrgnoyzgUdHdN7f+JQLK1IMoRhmtI2PcI6MH9LlZwHG
PHDnqfuE8JbmWr1PVICQSCDRuWLuPglbS6lFyhCjGAUf8d4fXJGksLzgKayKL7K3
lEqM5H0b/WZPU5vPT5DNLyj9imq6cBB7+RCS8NW9HzzJr7j+jBi8Gxg3YeE7ZIIx
Oh4xu8bphF9K+Y9ONrDrCs0TzFxcrFfTg6LVgBr8l0+ebeeI47kXsFpoeOB4O41+
hBS5pecanhctkiJJwLM4V/OG6ZCM9dP5sGhfCe/u+Q8HXJ/fZQJZGiQrSM2gsY+n
6/PxfhU45Sn0D4bdsbxy+ZwyLvV4v0k0R9JJMNYz4FiSyMdfGMboBay0HbVVUOE1
U0gePuZxyvkSDmpaaayM+pXXopGOhzd5+a/QL/rSjUanM6FNuwS/w4RzjOnREH2a
meTagp5sqz06Fslm+yfJZwBimpPvbRam0xkmQEDcZGLviUTW7KnoTpL/mmtzIgug
phcZPu5EWtVfxWgIYoImy93j9ouB4qMfef4qoXXZflwJ7/LcvbRkDhBkLnPgUDG7
2kVchftawL4MJfOAawKyYAxY6087T72IOcfrOY4gyurf6spLpmzpN19G5f3dH+mY
GpFQGAgQOb2nhxhBYJ4A6aYh2SCggltnFwI6jXsA6sf8r1U+QIE7Fy+YQ2aysVki
PwmQA1xgbJGmNF2X4DWx0DS7VezUI2icrsCiTOEIq4Qbca7kVIOuJM794jB8xDvV
m3A9WRCy1Xge3ReBgzZ/UyfunDWGi1JCkJV6ZpD51Zs+CJV1Ip+HDMFpMzRQTpRu
iFWrIc2UeWky1n/bsF5x5yVf5SEeFIf4aL2u+VlNIe1s4iJPc3FW2IsxymfpBlzE
PK7Ab9K8PDtcznf7PtcScSV/sp7wzPQ5jHSTZLaAdTFA/VBVoz4NYlnT6EfvfObr
c8RGlmMObMm7MIlzxojsvlK3CEsFW1UkoytwJ0N39z6novwVUfZM9lZDeRP6ORDX
vhYHpTbfh3uI8qkFk3Yn3MiAaQDkQ6MFzXIQ8K/bgiGFcTRjK9wChaihsenSWgKK
sJBbi54Jr10hyeip90HRJ9mlpW0GJ3CZ0QOuASiLQU3c86bw05nIq8rI0berxZcK
TGZ8uhdYCLf6ePGEUp0rkenNX0Ux70MP1/ZFmUaUwuZ33iHAcFMdKxbCz8Vj6rJW
iXolTDcIgLHGR1d2m76c/ZUpRrWorlt7j6j8Qt0+3EAzffJASD5SLNz5vMykoEOD
cvaQuUhOB3k0Z27KH8pyuwduw19KLCPieaBiOFddPxzTLUJNVNCbbGrFL34SuYcb
TBK1VP+xYXtunoAJoK64KGNiZIh8ejHoJiWjSgufEhrNOQumjVyRi6+ORv3dohwX
Qhs/BRSYjY0G5y0rEJAUk8EKs2Fni5vj+mSoZXFtw+iUFeQ4a4rK7ypyocLFL+pv
R0mBgMDu9rACu/1qx/xawkNr6Ng/3IOVYHkpYDnMUMlLAbvvlEDj76pSFUaesqet
tOmNFMmi0anGYQzSs9x1xJlBBnCue5XoUP79BG3KVgiFbv8FUyK2CZOFCGauM1Fe
py5wErh0FqOX6qlwSuH+m6QcrgzIRnJgHT9LWn8BrNBf/ksUW/jRwNZjmFghahbf
u/M8IUjLINm0YxKFoGH+6NUVtVUjRVxkvnJRu3fVMAAamUADXj+DPWAkTPdNMgU3
g2GIQuC157XihHrLIOEYGQMz3CZUWAhmYi5sXkPAHEZHauF2MenISlMir7wIupky
+1KoBVJPezlvNuyf+7uKAEejTAYIHob4rI7f0/DSXXx9wbsoFbexd0/ZALbnewXN
RCeWuykSHPmZyuFEfyIUZ08TgrxOk7by8VOoy9jlmVeQURzBxFJcmL81fjXk1tmv
95qGvLNKcLLXT9/oR5PdDrj1l/EsaRlJ2KeBULarb0mFMgeV3epjCYObLHLwyTfq
8PPmI3DdxT0AopaejZPBcYXnq9TXc7TJFlVEnhqoctszeGvde7+8Oc2TO1cWJIAK
4ZGg6IIOYDbkMx/0dnXn4lkXw3E7f+JUCqW8zYokLBqwDGhPhkwahXUpVnvGz6HA
5E8NFAYZBwqwP8Qau80rI8LK7cRF4uZ/OMQrVVFFW3GfYY3kYEuljeCTOuOf3V6P
WU8E3+SzO7BzmleTlY4+Cv8O0ErAJVBZPQ3IaWZHMRAy+hF/UAWDfooGT8bM1jG9
W99hQSbnoy9hLMXwUeg0Yj183/yKsVq3l4OQQpUmqLvZQ0mSdGokrrB5QdC35LGE
7Kw3XJ/5FSGFMlDOyPdWtUqs8C8kzLySfwofSKQ6D0BFIqM+dU13ls0Ut4Zgje1D
5MjK9C7lbQPBvX+0dHFRh8Dw0P4OQOOWzGydv2u2o+z/gOdU3ngVZc5u41vM4FX+
C4fIc3GB/RnGYyCbZWwOpvdKVaBAaUwZiRsTaxpXn/mYTFtrFz4wg0jQMKNY28Pt
EOjG8JszC35fHebTtBkaune8Ox9jaACZrOfvzarBYfLmDAm+iL/GQWCqAzrbXl+Z
ANsEWVDmJ1d709BVdA2UdaQ9DCr8i5Bq7qQDYwMfXgWk0JIDvSmsqCrXf2FkU8bb
366OAXuRDxvFw8feqxyIonBOH/RVOF+T7OR+B6tRW1YNZoq7gwM+mTqxcFELKQcG
G/hZWxlSxm3doQldJ1t2HTmVQPhjDHkWhjweQ41wOgXI8DkycEZausJgmvFtt+GM
ff9Dd3NGif1DB2sl2V7m4XYsQDUhG+cwfzqtoqHINPO244f5kS7iTO+TPd5kVWAB
cen4JTjtKhpCXC4QK+j8znCmPr5ApyUN/XBcEWJGrt7PMyljNs+UPnF1fZfrBmpF
YVX8EpwQNUfptMHNOhC8jCLmu+CTMGKZFLC/u5N8qVKY17v7wls7ifOrGdFg2r8y
URHm0QiIuHw/stZdQ9Vz/l/+E37EKONf2pjBlRTN+5cSZY5gKfUw8/UQcWjCTSTs
QeSSCI+X+77F6K7XdYGG298u83i/k2aYlBk3u/DGzox/qseUQNzkZ7PYONLzqd+r
CMIw4Zgc7UWu4V/kwDrvSxdq9O9O+5lP08GcTrQTj+oFKSQA6zZov6OaRPqBIlKG
YQBcwFuDiA2+FBskLPL8YySglIosACjDlVMap9S7RQyDatKg/V1+gEKt1WFo3ZhL
owmxfnTRfdgGV88eMUqWG6jAQZyBr3EqdIcviWpa+qsyzE2sFD86bvj1DaKuFo/m
pzt7n/62wQDppF0A/F2EkLqKVAALJjUQAx+6ffA9+DayJcoaM9ovwxYyWPAl8rBR
YK1mHIirogLotFx5/4/QWDmO635NQ1BqXhQqT78JBB0h6mri9oAnIpWQeAHqGFEW
77VL5bjc6ugFXGC8nje/x6slWLTTwe337kZiXXf+YgZetyzuT4R8ap10J9Qae6ZC
AiLXIyLjPrHY+YD+0u3QS0+Q5Zj6AqU1uzp1I+TPpMws27FgbXBgc1CpW1Kv+9mg
vs0MlMcO04MwUMcocfzlJGlQW01/2JpThJ1kQBlJ4lrs6HFhMrAdT4+hWeIyLWMt
w1q4MuZuCmG7ZcpN2QZdLpBcs4+5fD0MDTnSHM0XfvdM5WZrObvjy1M+EyrItuEj
XEjdQP6bw5ab2wCjwn+mTTIBioW5/BrrHPiM6vOkPckCeWhzNsAIhaUJrIZ990c3
gjobJG4R0CR06XbpHBFqPQKlY+IWPNZKIzALQ7wJh6ZONCH35A67MM2bUd0GweH7
XUC/sG+2L/DkMr0z10XRPINCz4cvs8dCucqkzJ6EICq61pXvxGhIavFwdEEg4Pn5
oBYsNsVFpRIX1/Y2bg0MPoegNlNH3eV1315K+50f2so6RqyhI90UBC3SlSNi117H
/bidLKmeU19HPb+D2WstN/DISjGwVhPq42pa1/F0s6N5YNqScTrYxg6/BrNBgdte
AGmVkRXnAoYohW0sP7bjm1PRf68Ui+kfPWM+IerwO4CWdtwzZR3SmdhY2SVIsOfn
NDW9rGb8imli4G2dcHSKw2nX314V53lA1ZIJS5hMma3fYTo3jLUcVcAxPhxe0ClW
ObtfZxcxy12tpqympa16q2RJagdcw33GmHluG5VQJWjNumzbjrEFaLcyJrTPisW7
Wj8iWvDfhToKnUpyNgeiue1SLs87Vq3GTWV6yDf/166yVA+6JolYrQdiUJ5BTlXr
yfzOle0e/t6YUf2oRICi//YpGA2N2cvnYdN49aWHK4BwztjxsRJhSMETupIA8FAG
GwKFrxsJjZln8yLjMoGfeOroh/Z6OmIHwM76LOZ3tT5qtUJdGx5F15EJY1wvZX+J
07dHEvm6A8lAD6T3Gi8aq3GHSqdPKxUWn2ur2t2iXsjZphtc4aV0QBoyWuKIh2Z5
wdN+Ywl3f67tA8CA+4ZvnKtoMhZM9py0Mq9/OAV8Ycx/Ha3J7RFuSsjoOGub0rlH
aRm5K/nZ7Y8B7ckiO9WG+S5l8vWUWrJFVAPzzDsItmvAb0E+rNH/NZaHtRR4rlbw
YBKNa3GxhtVldCfNI+D1QmEtIvV1gx0NZ+DHkmfYgYeFQOXhHt+rkN3kOK/jlnGG
ng8+3muKIqVZzulfGNHYer3Lokh47y7m4tekKfN1Bw/otSfrH0xb+ehR7G5O5xTo
ZQuQpCMZ4dlFujbCFUwD1rYs3z6sdN98UT5GB1cSocHsFMBmW3mVWbe+Ex7HzxQC
dn2ahk27tStf/cG4cbY6hzFbw8N8wZJ/zwYZ/h4vTtGHel1wvwWQO2jmJdK2RBbl
7N1bDuRhfnQCfF8IE6zSM+5FoDiPoXcw4CJO8nGMhEJQhxSnu0eONlWBovjSQXGE
kNbf0FWeKNLlY3tRgc9+51dRZCpDBW0FNM7fKdt56nNHQ56gc7unuHOLI9SQXCzQ
PnEkMQ+eyTBzTl3hPH0lceEW/I+g4Ei7q9QS+xj+me9st1zb4RsV+WPH5PJ/vvL2
DMc5SMFim2V0+ic4q3Sb02Uea8jk8AXBJrrPMXKNB6M1IvYjQeCN6qcT94qXPhZx
/C/VCdOeVK70uC6rk4D4cRO0XvilQkOBaHi2XWGlslz5Ph9Vfqu0RuVeP6AHX0ay
tf1mzvN/mC4+KN2JPgnolLg5Yh0DGaVVYoaLpH+Lgtpvjbh+cVdO3Am8lDBmxxPJ
XpMOe0q9PDQi6cmlch7+wX7J7SYYPEH0ldDjWuqLCi1WIY0cQpEZeDwTPeydHVKj
gBC8An27uqXKUhduljXp5Z0fMGk/sQZaB4nWjQ6mZ+2n2enQurpriYvK3MfS7rSh
alMc1CNVIHM+yd5NOFuH7V9Q97p/tvz8TBIWEaRZ37uBHc7rA81CkEAvbuGTEEGT
vPXNO4cr0ZLQB07ibjfFkk7F9htDYr779SLHQn/dbfItHaiilPbDihUs+N2VFjMG
y5c5xb+8b/RLtltooPquuNUmN6k+ouGxtjXy00gY9cd6iWH4CZx5wWyj57pTT/IH
Rf8MR6jPGa82N9Cw8GOUtuSne6Xg6MIRTUzYU9voJ/bm9YcfSec9rzdp1ASr1y2L
bLi8yt6xlDLHy6dCTYt4uW6NVg7DMSiiJolIz6bNNjgRzPhXMGRbQALz4AE3V2nZ
NyFYGXH+nqaT3SOUpaUG2QfRr9tpxPVbAu7EIHN1U4RzdBtvuTWYNid7LJ/3qXPs
44jfhIBHr65iriGvVMTVHt0MMyoygY+d2pmYtSzLdXsSTjvW5Ogocjy6ebQ5A8+P
Wuwta5xSc/iPyfHv5XUw+Avyow5QPjNuMHhfVYH074iNu7dOFHURpGqsh/tR+ZSu
cx5GBR/dBRyxUHUu9buNo1IRGF5SxjQ2GVi5h2pUVw8KuuixWmowc/E7hTHT2vG0
5mOx+33+6MFoGCIYIvujbrVIAEyc+sxnEEpYXR6W13GnsWS5uC3xhqTV2oHgOncj
U/59HuOo5YIynUy1qd54W44j8kI5NPH34p8KAuhtB+zSEl7WLVd1thNeJToFeJ3e
T1O+HyPJyfqEmZrtz0g4WhXQKJtCJ9dpr2fvN+S67s5A8nOjbwnEiiqHycPVwe46
RksqVMYxrPen5IR/2eqe5Dx1ML5j8Uf5jjY4kgWaVgH/JimN5GFHi/pJomWTBDZC
sQPY7/u2LzoTdsQLEcKVwQNY+yqch3vpElsEaaFClg+bA/fd7/GR0nsuV1bWPDXQ
k780EDFytQChN3oQncrvAKNKv5MSXCmHVgAIsOeFRnPu7REiIPikaoSAqkFoEB6U
KFlpf4pTYEvh11zOZajzKt71IVOEYE55Ai9qmyVAsieTvheT6co4VPsMG1V5U2Fy
hGkBx7V08Lq8u7t0KDAzYfPP7chk8oPZH+PmH2D3r9jzkKuMjDfORXpk3j6Y67YQ
jVpEc0TF8hihcXV9i4HS8UasDngt7wyj5yO/AXSom8aG708yA7tyc1MkX6uxeRx7
7CroOL76i39xXVOKuZ9blaXcZfXKw579791+wMEbUvrQWTGn0WcbWNx8YDYDvpri
ZEI0ISOmSkjojnBrGah+soiUrRUaVc0uwqYvUkwmNW8gnM8LdEIiXQ5OAVY54eNM
d5YyWTlJlPGBMpFGtwEOhNmWtLhV4w7CMAYlLomqvW3TjMLxLJbDcDvCKiz0dVyz
all+4xUUBk9fBQs7qf6UbuQGgiN8EC783QKniE2sO7ltGhMANPZ6ZGiI7wNQLIek
81kha7FM5dQYM0yGWNURmapcihpoonf4G8a6Uh1dnwoFW5evqZjNgXyB4qeDSGdM
9JR3kYR3WsZWmZbcnNK8Skv0UKWXAG+c/drGqSpxMwEYWieTcO7gRwY9FHJna9Po
eTJybyezAVKMqoZ+ZTqhLwqRPR7agJi04VAqFg/BXMtjxp8fkhUPIMELlyl/ixI8
/Ky4RDPrmno5dcjs7F9jD7Ik6Ezj0aUS513gUurq/2rV4RrYWZIDvyvGgPo1qOw5
rI4VazzYmkZ1MOhvJ/iuthVGMJZQiZ/tDPtHT1aa+lX0C8aIJWU1UEHnw+6fFyWd
l2SYYhtaVigUnh96oH65hPfttbWtqqlzcykAqI/wVd3rMNFA7ZCXVr1u4h20Up2T
3dlix5DsNwdkdhxTB3s7sJWt5evJDaxdkz7tuSdBvZfLdBEulCNdMMw2U+e1fay4
RhDODkaslbc6Q2viz2/uarFfMDXcHBHg24PpNlfFDIZ2nQd5yy5afngEBkCiB0ft
d/8fGGdV10gzQwfl/iOMRKh1CW8/dyiwpwfVVJhineJlRJbONiUIFpn6tnpkzjb1
fqz4+RwzRH49Y9wtaKIsjLCep+85bBaz946S+qRpYzRYOkQm/QfnwesMbk935JI3
C5qpFbjlX+nHqULS8q+SDCINTFf06YLz6STYXlhJEiqjtCsPNpdbGCuygaEmk5la
UVDhYs7JBPKbUFizRJbEXyOzbECXRaWlPYNXvJY1v9CiP5MvIVQEON0/5NQw7AlK
9QhbAUp1RBtTRVDnkOSTUPMzsMUyR/19rhzRSDhTCDT24nxEQ2o8IB2ypVdjav3d
S+8Bje+Sl3DQjx0iBDQ9EAIjMwvzB/LRC7co/klBqXNLu9aylBN7MJxMgyy8niFI
kdDpszGX48UmW2hZP9Q9W8Dhuk8OdR7+SlNu1Zg7fCadHwNcd6CfVbKfh5eHM0Co
7zoJcuTiWxixFU5LpJhc0Ibia3vcjJ5Q7fpWLnkbVeGVrSqn4YOsJR1CXNuXPbRM
SyxLkpluFVGqxlmxJ3ZcluKfHX46gcRIZONisBBae0FGtrG+YByA0Os89GFDhwMX
Rmf3zOpYzSt6xocNA0Ocy/EMsFpFXcxdRiiBI3XVLGPVZSURSvvT9h7PyDnIZJ2n
WwdPfBO47FWCfULteFSehCBzKUUIILtfv4vslLBxQu4dmT3gEqqVT+Cp8958el7G
/BNRF7cR7q/Eyt5Vo9rxb8vbRorZo+eKtn07ercyWzNwPCROOh2TuUzNd7+HRfVj
LG+ZX7bcj0Li9vjPXkuR7ZKQhwTBILMWqEpdh2qKmKTsJPlZVA5MO2318IPsyjeQ
sy0wqT42kr1XfmjQpYOYw+FZEvgs/kHKT7udnYCAgm/kwoG5iFh8ss68YTTO3X1M
8PErSEYJ1Ae8e+V0dZVJVD7StawEsOuK6O3HZmffGfmPpM0sRilZhWf2pXj9DPDB
hOgImoaZ2J1xlXi6MJzRJsqWn7U3jpx7QRAoptxafBqHR1HdzSwGps5ihtVmNGpc
yclhXLfo/uwtysHj52rgVzZvxXh5GS/qtstPbkJiCp9xsl6r2N/RImI+t6NxRpt5
Xu8F300k9uu+X1MsWWWRgv+yeT3wBqXPpg4M/vi487l0G1CnzRImDty33OfhSMsy
uG3SRr4PLdtDf/JA/OGpvJUSnIOli5kOhKYoFMloCZg+2vdsx2+ZyCAAyu/qVtWQ
8nWTO7Ld0w7jHVLKnnY7klB9QvO+XpniEaN5iX+vQDU1hCQ1HcAMYu1Y5uKDvw18
uxCCo4BavLMi7AgOx9HRLS9crU48a668eTMWJBdKWJWd+GjrbwlBjD/hf6lP7ioE
2Lxi8GOZx8XVeGtKs/ZdubJWAJWz5gT3ST2YNQ+UJyHBeO1Z/V6tXWmx7mghGf4L
Fxr4Yo0sS67oM0bDUamlBwKviR/Dix/KaT59+5+YRodlWYSMzgizRjvNquqNfNJ9
pVLEBoBA6WJEBsxdqbAhVzQqzcQ47xnHf0Qu0QSRes0FehxEyVkVzDUnhxe8h+k7
kNLFw3gHVWaZeJQNEFNwsYLbwWLrqspYHrnyl2Hvf0uSLuHMrCpMXHnzUPi99792
fmjvBpxPIoF3G8LcHbCXnTiae9M9kY7PyaI2R/9/0CWtfNfeQ9CovFYRdwszD0g1
yywO/ROCWs2EvQ8T98+tjygEJG9tWE4IJYwN5mbt042N3g/kfn+IQNAy2VnE60gC
oxOanUQkvzN1acYD61kaNN02DyVAOHw08m5Ta7DsOWaUseDLya/OFvUmdTie43w7
/dVN+1AFPz1GQnJeFcc3SbBNpQzOwuQarfe/3fU0nRPAoc1fOGtsdr1k9jVJmdNI
+J5+OJzPvN0Cb2XwvVwpaFb/VdOsveilSpK/1bOJ6eevrVH0/ninlJyjUtmBb3wM
jhATZULiGMQV4FKSzvNlBLCU7MPjUxA9F/LTdBFUW1NQbHJt2ggSdcRMlfr8xxuK
6Fj2sphg2oF5YXhYwCNRp4zrYjC6M/anTyH/32tq0DmjTQ6w7yMttJaejMvapzij
Q4JHnX6L8LyhpP8naGKEy4Fd8gZox3JWzHcIZeZCFsUUIjRP64J+SbO+Zhrj1au/
00rVNxt1gmclopr8mikoCY5KOp53sa8WxjRRMjRYVFU2813CPa3bkAHDnjLCUylX
Cd7Utim+ZzrPDZBZiNJOYU2oEOLRIlXkmZJklx92zxXBZ2IODHGRZRQC2YDum5i6
gJEZENl33uXlKladRnB2SZbm58ZaMsMljF0Wd7OImpMM5mSvHKJfx3+BK2sYDY5/
1BhlvxxPdlX/b76CbiQuO9jviZbSdulCRsUfOoMcR4dc6SetUQoXULfAKa960V80
/LjuEWS/yrmfqKgd3uidbHzQg3wQQ1yabAr+eswU6fh2LGYZVV1b4EnoIjHyB7Qa
oWuhmzd808CcBYVyEJQgti18wna6JHckJv6p6QoUdmvYXFlcXn8tBNukAKTLnC11
RBRgUBoakmOm2n+Nx19Wf7s/vVmNyGQSMGi6YfsGT99L3qVWaKvBBBlWRZHbVrkN
Z58rrFaKyJ4PvnW8CFb2FnrB3PIoyJqDaXJNCUoMtZCQPtCKAJqSn+KimaO6xSt/
w2xI8TnJTkCWZIHCoRwq3RlaTc4CX0WcfgmJVXQQKR3A94OyiiDgBkr4uQKgKb8H
oe3a8S2KraEZyjJIq4smzSHmnDunfdZcxmm68kKa4Ng4LCvW91xoW+meQ2zNonX5
HpJnoKZ44W32McIA23r1yctV6w6d490aNWOSSOERiHV3x8sk3sjAcx4lLbYUz170
Bh2wtpGKpqgsr0un08Krmv7EzQaaCgo6S1uJLMpm0LhhjrLEIxVjK+PQlV70SNza
NzXJl+FHIfvAkIyhXtepZX8C6pO7BIWiUyZHVJWBJbin91/4fWiIpcYLQS38Bw6C
CuZctQv8zqBsSOex+gyyxxJ3AegzDqPgR7dXWXTbSbRxe4BySsP6sM/uW6TR/psj
WbUZ+/HDQ0vA+cYu5SXAq/6N1fHScYClD9jdR3xk9RTZq6HhjzsLaVMVsdsDOcIn
Bf9U0cBInhJaWK9NZIGkWoP16PDZ/7grELTxJP6eFa4BBtty/2TvbDq1PBjcMzWd
We4x1y0SAw4XOMspboYq4ARpdWgX3wvHGs0YcW1JkPTjYy8LcWVC9qgLnjZZT1pi
iOnuczx1mkeBcVQ9I2laDD1M8vdfI+3I+Heq3vLAVru5nn3XFWZeGMk4hmJawOLj
YAFEp9GwS6/yF9zQreRGwhj63a3eFkcdxE62q52inD7fBOUTzOjqM8s4QCaswUGp
goi3aba9/9AhYXKsmtSwpL2YZAu2IFpGsZegGGpT+RrRDyNGf0GPZbKOftMIsxMb
e/lOc77vT4IWXgbAVnEBCwsgw3PYCepYqEii3FxGKmi+YFD08Zz8uIL+eQxlSyIr
F4/iHKtEcgqZ6eJyZHU1uw3Nqd0qGCqhTmrBFoGx7eNqg6TbckpSfCMS9oCzjBHq
Wviqqmp9wlhR/gz6x8FDD19ghQtzgStBdq8e4lIxPkaYqc2lt4jNYvjSmr5qof8f
+woNgsuKhZlsoohmg5zRpwQxyd/LVsJN5GrQ0XL9+AlCKb34oTl1N6+GecFav3qX
R2XAZLrw94p+KNaJrJhUqrJbCXrFmFd4S79T6+EM3CrzHOY+nsBWvVO5fN2rlnmA
1A2dPXw/AImPB3Y4ZhXxCZ37b4s6m43ullbVY3/STAGkI8rnhxFog6N9RNmfbw53
a2bkFnJ+V25T7sWMx4hEtaowrsHmqCByYJ1QqsYeop6O5zUG6QBYdofhlsOI8TS7
jvxEUdzFgnH+IsumZVNDgtcRML+jWEXIB/yAmdAWtsnjUe77egnhI91GGgp7F7Lg
jSTsXvA41I9KrU9nGlWVUIh/22tkJE9sKZkUTOWvfNNl4DaLpYDwpiFS7OO3AlJx
S5XpJd9IKGdyZwH+eeKKCKYJV0ubboAjgbp5RqckuMuwcUvIh1iqUIDhfkuTyGT7
30Ardv6R5iQoJPPmHZFfC5cFVFYY2KX7e3vnJ/9s5CrYrs+oJowirdpVDWNX4mX3
Dv3dJuFLjQ6AbBD1Kp+9ajT59a94F/7KUMEBnVroKMfTf63G/A4rAjkk7T+9k/Af
6MlefdEG3CmEJjYBd2bynPYTpABQNZoDoH4G7opDvi9lQ4ASBDYIiPTHLeYiLlkp
jj9L/tX2eyD/dCjyitfpr8Mhl+/6of1+LAUfD1z6aM4sDLo0Ljn1mXecIscxHiwp
f7AvzvpJxAsgZu9a6naUPD3zkRDiZ4LMHvuFUcq8iClvqXNIu0oq1v5ZsTvcytwC
aSZ8xsQ9ZJJMOf/HLMsUHwx7guFYh9ZjSrhxfwPWF3RP5MtjDqgtsYJEd5aM8CkU
M0CN9M28huZ0y7ktScl/83xwlHUyXZdvudaA06hDMbEA6lLUc5dR5iHVP/wxV9ZG
H62BbDutVxVIj9+pvmh/+HkO5sJN9sM2lj4gcqHN0kg73w7SLFIn5ktAp4i+uIwc
ms6mi4BY4eX1Y0cJdjMFd/DI729adOIoBc+3ks3ZIRlsW/iSULpGkqie7QCzLKWB
12vPjzyeBlo4z1Wq6r3ViegrnDRTEhhY7IUXEC/sPWkAnCSX+JHLHlDx/Yn6kBut
kwhmcPml2XaUxWP23NtznIEgDFVBx2i9iUZCavZePr5lW3cgzEwqzb64xhb44Eqy
dvdIG/qos2IyyC45bp+rLuz4KM3ntPVvJ1xj/yr68yOSa4+mENhPT7xI5DMjsPCP
R5mEK5z8hdNyk4uJZGc+BYvmNwtaxAXljGpA+lkSRTe24evd42ZHdUcN8vh+eEqB
hGyGyO8weYB1Xt6tBAflmUxUwZk43npoLoMU7ddRsB0E1k3JQ0xIoLea3QKmqeg2
5iBXWBxb9X9nLyJvo5W9jo+PP0NTVfXPkfJnSj+jrEGeBA2pkpPkzROif25kiUIM
WM8RkdJoa4yZVl425z/xw6DXJHKCl+eAOiSxAGrwEsxsmYEYSPdHVoXzw45PpJDw
Bd1mWLdAsoTJP+lAzHrkiBdisGhw7Y83CXKkIP/fdZjL+R4DGQoZevVZkHgq9rxj
k6kPWBbdXaBWrmW85QyXy3jOu2NV/mCqIoRb9+0mMgoiAlAQlLF6S/Se9AyTcZU+
TVk7lc61inC70OG5Oo6+Day9zb1LuDnxkhh6XVNLORBNqmghoe10xgve6cH4XA4E
QGiDkWMZBWiLWP/mVk8i8cRYCsct2ueCPujqHSGkQkyYUxK5JqSbew9mBqY3you7
9y8Ccm4F0sgJvWnks4mwEkfWm6iSudiMpUoz+bjtaauR5AIFvscgpw7AA8qNZeDM
XyId6nlDhe5vrC3gfIkdYu6DEZwfii5QYq9uezi9b5BQHyQtcEDFp/2VTXko0A1p
qeCnmI3yJlx47h1ZHssVj8DDOMG9Qq1906koj6hc5RfbeOmjBWFGIK94O64dqG6n
N//fXm7gjTdMAXstIMMdw42EDAGG878FqvYS1W4We+Hhl89Er6kwZOiQhkauweuo
7hLoPW1YsyygxmQIdmQrXDJD8EhalMiNXDEjD+KyczamlVzsnX7gs6KY/BYE/0QI
LUEc9y5RHwFNP+mZmqHm05BCU24OoEHNfA4v4/vLKpeXz8tTeoUzGfS1+6fNhb4N
7bfRTjQmfZqmplvR1eGlEuK7g9Q2RyFcKDuFNpJyJ+OwSaJGx/G5Lb7BkC4gjzQC
BafFzXi4h3qr+4iTcps40NXTdgIO9YjsgC4r+tkjmQA27yggKp+8yQByJ3TjLk+A
Ub0NxV29rC08imVmLpbuYr9Ls8r30mhYETvGDF83qp0uEzco83htUOOaOSFNdSTD
mOxAjX+ZH8i8HDstbNJ+uss9JUhZFdluC+sNsABd8Wp9C3bct+MDqCNL1fnqBPVp
HFj0tr4eoD8LQTnjpRaKsZKf58WfeieFcg6YfWE0KyUnecmW3JuExjJV+Ydg3kpn
zjtBV37BGPpyIIeIou17xoCk7CaXims09vax83FrK6s3fxRawd9MuudbvPG49LyC
FWb6QkLRzJh986hdKF2YVFU3pGgZiyB10bZgsMLq5jHRevEFwjsirQ0h8ps8I1zX
hI9tXJ5Jo6xQnV7RcJlyouCvI65l5Udg+LyFt1yWBnrR1ltQdxE1CR9LM7CPGnEN
16n1ilNtyoAirP82RfKJe57knON7TLkPVPnxypJaEpYougi7/byw4YAMSSoP7lGN
dW7KnQIXuc5DzQyvNWhFVOQimvHoUOMR8BChlJqnuZIBhyRiW/agDlOxsBNOgeAl
vOBL/3BVq4uMAQjnhcTOs3MlH7fjt9AqHFlPkiXtXLzaFoNpwCenRPwUfzz02hIi
gctHAhtIDLwLXkCejOBUROJKjGjV7zocx1tJeUipLWJDjrfagLSRK5E7i89UlNXu
bx3OGB175kHV8asV7de1SNOccyggKjouhXvAZSDfcqCHXIGsn8KFa8wGHEFTpaIa
OJAHShHy3rQDrejCEkszOVll+mZU3O0LVceroNaVibiv/UnMDjVv7ith4yZ+kBBw
V20nKkxxVk1in0H1PMynAJWBCcgRx0zP8OYAICObqLkBDkAAfABorFd0bfvbAIo6
MhuKUzjPikLhYh241VhSiOKI3Xc8Yv7foVkW+tspT4FJz6lfBq6CUrM1j8xWi8gb
DUXs0yHMrsosZ+X88E3KbdodEhbeW32E3YJzAhWGCQkDVYyiGlEW9DKa6fxjuvwd
6ooEUYFqJ5DHSt7nC8DGDhpLTSMutLuRiUZxbQXmC0qdpp4fSBxMPiWaxBshBIRo
0qr15RkHsu0GamXtfw/00bRmgO1Ssdxvhfqhqy5dJP9G2cjtExjSSpDHYBxmCkQu
81xVOQ/Eyi8/RQF1oUH4dmMznpl0pMc/FZKDmrUl7a66H1af7Ea7Ublr0zsswfu5
PF4odS2N7YBfvR8nABRBDdDXnsbeDpeHUdYqkgdat3BOL9mmiuw44UXwq5m1s8c0
WyPJtn2+OfzMEoS5mbcBMal+SzdLndDJ3rKIbX/S/JD7DTLsK6+OM5zy91uGC190
pnzPUhUoa5SbR40iK0PrOyk6XKPZzuQgw0IrrlfPTC6fDBCrw03VzZOMOablWLXm
s+qjmNIAnaP4CBFetwrOvQWbIYxjVi6ZhW3Paf7aPGlOKagUkU5+YsxdslmOeDw3
BCIu+grTRDEE4TeIwh9SxkupZmWLLUNEIHVXrH/PWynHfor1GULmImOw4Gwz0qiN
uDIUA7DLQtqmEKnH34KazY2HJzdyoZ0zAGGI8jc7Mz5KE6oRGmWJIfEY1nRxBDsx
MJGvC8Yu1LQWB+5Djg/W9Pha6LcuuUmDKL7c+zJcgq+w8S8eqypVqIk5dJ9pymZq
SiUCfeP/YsqMvMmtRNdS1UVCAbmX6B3IX9VWvnprOzoNnr7fpsmHVuU3vVNaQOrn
S3IPnXqZmSFSC8u6KdNuCRQtSI6r0hU7X97Nd/hRjj+PJ8/q+LsUXYomGleBtsjp
pPbXoOMDk/6WCh7EetyWYmKg0wcUllV45eGBsha77mF5TjIOuwn4tJLtg01YHh/r
M0U47N6Iinv+65IzxwJjly6wu8GTViJe3cR+tOl9HrMaUIavHkVB0kCqld0+FSjc
EeldzN5cgkCB1/yDBXifvrsjNUUWJ5hHeUxjYv8yyIyDHcKeiDrI55ppgFoNjer6
NT/IQ3XFQQ/12TpX5JjsqpbtlBJVThLqPa1MWebWU/tiQM+35DH7Iz3h2Vf6XBlP
UjcontBShmdqQskLOzMz40NUoc2zy7z4wDb9mxGLmfcZ+40gnjTsv9Pwmx9c3Hd/
1caZtUJZk2D+mZyzb1ho1MWlZkQJ/d5eKK4FeIU8XuV2lvOtS6xT1dMabQRyqgJm
TdbAQpC5DtVpxg5vECe/w21gvLamxsXdjhQTAcRXw4pGNda4wvNm7Sn1YKof8rnm
Z9zThc1OcuY+DbYpi47a98JqRSf3yW1rAEmSmRS9af21V8Yp2Ko1XcoZJ31LI9M2
p8XMbrosnDjRVg33ji7+RMPIYEFzS1g6W1DGjwbvyfMi6WGAIKtseIvdiaLt/xKq
HN9USRETSqxILvbVyII7+WcEHrYQmf9+y5YCk6wDrHYQ2aIsc7umzHAyOlQmsUcJ
LK8D4UUPbunouhOeDUNeKkAt8vMHScMLbRhGcgJ28PZI4sbQLQI2i8Tl81tNKG7o
jBDgx3jTBo0efponrD8VJV5uNSqquHNDHML0ta2uOwsNGadSvzQAM7OzCRPO+hzu
cWP2cLgGWvzxee11RM1jYr5ReJOKFNLdX7uVQJ4yVGb9Q5Dk3gX7wmXe1E7Cx/My
ybEFQltsX76XHu/ZBr+AseZzUf+CBGcrCQ7hFdadCEvBFeTAyKZP/v7ybCxMDnik
gR9M5mEOO5PgKCsKxpVCBGcFaDRyNxi2O5ogUF2ZRSb4yTIpE2/Ik6XpD/l3nYA1
EwOEiOQIq5iJxKqssg89DcnIcmChBIRIHusZGJIRzdC6PaGO/+kH6i9Vpina3SnV
faG3w/gzY8PxZrhoTINoWSVW5MJ0QFG4vZx7DvgBf+Dr5d9lW0oSpcKRFlOM+MwF
VmJrhmPjAr93T4h0Ce0KueRH2M3WYKsbJsRdlaniVL7NUSzBii9bwp0WWJHp7Lf8
j8/lRZKy8SPvx/fDO7aa/Cwnizc3e4oGvLWSXhuQgCXzvZjQwz8RI9a2/ghgHPuD
WQPV0285Qg8tfx5dum+5F2eLVCyThwhyjeaaMR5xrSUcFTPAjbMgJaBGrl5KdHxa
qjFyuYOpmmzzs99KBRYDfAWl0ac1TvJ4n4K/4A26V1BIS48ypRG2d3MTxVpI5t4t
JWwrbYkf7A5Ho8Cl/GznmcXSJQzNm3iKJOJIBACAToacjIDYOLcpm7tgHuQJr5cd
LQxiqI89xDdxDMl47GcXkQnlf8W2lCJ21Xt3ADddvUP6jZTb77SVQTNE8sz0/as4
c0+c+pV7iSi7/gNO/KOSO2WBo4E8Wjw4AS5pzMrm0TW1zLC7hZXsO4NFDkrnWy25
Flzn6xWycd9fjW3LHbTmFtLpdx+hisGzqqXo0Fw8t5rp7h2n7WORSuXOYn8pI837
c8JjzIgkOgRVe8kDOISFGXtGBPHoWYLfVpv12z6XZaokwQH0gYtFHlYh7tyYmvcX
nWSBZ2Pcl/zwZfX4Rzds1bzZReb/wRlqJzyLDI3X8Iq8No9PWKqO26/aq5vQY8Ur
eENre7D8ltaQowwtfwO8dYKeDCNg9ns5aYZc2wcDLD/LnftWEJHG50JeY9lqBf/F
zfpDxd6/vEsuzxXY0avoCAbhMWhGUbXCwsJ2CiOGvEdgSOF86dPGbykgDaexB+Yd
1NtfioziMzQwyhChAmwyx6LptsnOi4ybry5hXDKbSaDRcX2jwhi9xS46y2f4YLmW
mPy5aDwkZcNp854Z76ItZ3h85lHqRuRITWoK9fWs8EtKg6KP4oEG2RXXIONTgw5w
ThG/hCH8Pgaax0iiGTmMh46+9UGEO/3g1p2PoT5yqkuhmh15iEtJUoEgeAKLvfpo
BfSw10agFhhVQI9vb0HTTwBqyzke2uQTN/3V4mmXxxtVTn67wkfWu4nDwsidYThU
TvGgdjyDK03izhmsVo2n/3uP25bC4931v2LDENkVN3e8ijJGPjq78hTvDoVP36Xs
LQn8sU2WXuzkv7Su4Yc4hvXLisK3+drHOfuqiZLSOMPMVWSjyaX5lYu/lkBqyMhD
ShJwbTyfq6jKlidThHg8ivYb314bxxUu9Xivhoh7kRmqkbwYHRx6CYkoCl783viH
Qc0hdcua3GheuPPqpAvQSQkvrdcXnJNtFMcibKis7rMTOaTxaFon9U8TrgpkgN8p
3GYS/5A5Jfbzh4BVxLHUotoL3jIcmjCzaoK7fHkUn7SV/rBJMxWqkdOpOIYGwDG3
VXue/0pNmfsC9g7GJ0leAb/fH6uYwiGh3QrHioOuGgOtcKjkHV5Pvnhx2yu41wCg
/9y3/yOa2IFWmaxH1HIrGjp+5QpLunWiLQEizhjRmRAuO4GyxVupae+5DcTTCKLO
zz8pATFBnTVrNAx5a0ttIkiL/TmOzi5lIjRnIGYwL8Sfu7dn86Y8F8E2a5o4yBWW
ElIL+ghYdOHKg4ri1y5yi5rvclBEuuPblhY5i0acfN4Z0ZYMqNF8YCeCbDNkuJqq
f849NdydqDzI/oW6Q////2bDj/mB+eiNevbt72kEBfxAsEuOnDsbyeasGo1tiqn5
Yxk5oC3R34EEueLADb5Siu0esoZv46APPXZpINZFSZEAZtpY7FG4gOUTj58MoWfM
Cznyy5EqCLby5W9imyq4T/jLHetiEvJHjZ40d2E255uCq8RkTLRAZ43RBthnCL20
/d+DJ4RShwFIYpzdRXvmuvrSGzMqLnpevYAtzzKr5nAkL3lxGnOqz+Ea+Det5/O7
S9L+6BzdlNc5otM/qjrnUbDAjewP5cD61tcYINoy+OGv9/Yr2QPplVr5bxup/77T
X3NTB/5kyNJ42oUc9VS5mdmZJN3j7H0Shza/4nAfAIEi3EYOpk1WPOMo/8vU+z1N
dkGtsR/Hv1OZWpKkVSIDqUMQ5XNpPF0lEHde0U1MWyHbfXR1WnAUb6iDEYBusded
ckVsGhhzUzHTTGqBsaP5uAi1jhUUdjZU0arUedePYORfn/g/J8dntsCTdDnV0Lst
TzJ02fZrmkW0/8stC/AxGSvGcpdGvEBTPqFrKlYLG5koAoIt5JjC7qfl6+5pYjzG
7jGpu82dYqR7JZQOvylc6vSZI1ozMG9NBlWi9eZA6SmdCKZdqnQfI6xRCy+ZCP1n
Dty07h1bIFHGuTucbEkOmJyC0ewXc6wzcs3OsqmR19FAE/terZoTtWsBqSIOONRC
HtakIimemBMrXF6Ki2gpcFZ3eicFtOoatlX9Nm3/x91Lo/W0pzbvtsp0EB2y2U+L
/A7kfQcMozJnmwgFe2RDCffPpdKyHX/yQi5E1p+GRdSLxpw2JXldKgKcUF0zrKZL
SJONCQ9hr6TgbV1q3JkCLDah8g0FtaVPEgIK3OwKwplJgEQA1V2Zx7+JXbSejeum
jEleCznPQpQEf8tr3H4lTxAgaNYSJfJq/SlShKnLEWpHxiNTQsVPsvFSjuWrh2oA
JATNrTWcg3bPO+fCA+8hTqMAdllquzIxreMzDWqU+ViaPqtjJUP7C0VBfb/4toOM
UruKDpA3owNdEZTMNzwaDW85solIasbXxpSyyG/lzLluGP+DoDC86Q6+eEDaYwI1
Iu2wVzbFa/HY+4NF9G3aG1Ln8M6njIC4DukAunxyOFmcqSd9AL1YK7Lo+AfwseXV
JoBESZqKJz0IdeoPWCqY1RIG5GuKRWoe2rQdLtTs6VCogqO3xyoev/Le1QmklZJj
hcbb7FDJfo2xTZA97eUmuT5x//PWjUOYJ+QpT1h7nvvOF0I5xy36FYVCIQdrkCO+
+SovHpIkmy/vkLBSWD8erUGLJBV2F8Gn7Z6NjbbnbCOMI5T6YfqvT8Nw0zqfdKeZ
MlhtroWTd6XhTftG17SdlzPvptHFyGIAHz57YElT3ru7kiFQVRuF9wvGoxp5s9R2
W5E99kGlCJlMd5mTmSQS5UKFo5/nNT2+LtJcqt+vrPgFwhhlhQcJMsffsrMGzHAJ
V8Ml+xqn0NI7ZqqzoJTy4fHEy4iV3XOht9gKTVV4xt5psYcfLuSiYWfWhAxBf8Ph
NnkLMGIv0amWgBhOJMhYTbUdt4eSFkhzHi4wW+K34FxMdmPk7IcbHvgSfS+QHLTh
0x+SuWg3idqIMvxgTXOhNQz/U8odWMfg6BWujsuqhdcmYO9XxzD+VuWB+TYy6jOR
2djmRao51aMhJtif7CM7fofKBcE+Hf+6TLIGQ3R74Ex6TkFAMbP+H+U8xyVjGIn0
dlDak7+m/YT5nf8r2Q/YjirN3snLNHnfV0+31oNnsEIM7ka8X80amW+dGdQk2P32
EY0lZDmW2nZukf9Np9zeEiV4qB8LTYGDQmzaDuRQ2Xnck2FyWqBxlpuuqXc/4Wlg
P3gAFGFLY2rbgkVM35sodasul2B6cCUY/LX2vFdlVEW9cqw1K+fGOrPHdB2Zfo43
6g/lHu49kKMyKv7R3yA0HB7X3qFsbqk09XWxkxkPyXrFmmJRKcvBqwxJikvwltJ7
D1cxNBaOtR+5n03XHywebpQSkQ7Y/XgWRk9iVLvfJEzhTegqRmqdWrHRSm5FoyPk
Wote45zxCtAih/5xNHGhRoIhSJqsbDB7p8Y2xSd+Ke/PxS0XVmVRPIYpG8X5hZip
reyqYZhFvrgIaNnUxBMnPPMyRycEd9pv5eiod5JOEPLN6KXWSVapvk2hikuU4fje
QvyUbAXRkN5zWEvaqnwOBVdmUAShcB2HcoVRMZ3zARIe5nk76F40OHx37EBM8NfJ
5kbT1m8FG8bSVbGtG+b/OrBeoljFHDM3QsNOnjFubIGSI11mrn/d42V/xc7MORnQ
Id8evVLH918fK7WgVVXYzisR/ppBAMgc5Dg/vdrwFzmRbVq6TTBj+2qPA9tkprgC
Vi9hSge7nhLTExzMt4v0xD3oTWURHvg5yfwlyZ4JDYvYfenLQ5qPfFsT3AbEKA7C
HowSpKtGaba6Ul3AiVFMmld3gkryjFv0f6yKvy5g7eGQvd5uMff7V/49s/I/cTg6
bYyLSc8eeT8ZoI2b9yCg5F3a2PTj60KJMh6FyW4O8wWTPMQT4QeGRR4hLqUelob8
QMU2Q7TG6sk2anVao/UEWHpr7faokLt57jcHxY/aEJfW1rqZLrCYMXl2nttKQic1
tkt/L0LVstMi9nX6NPZK4P+KhEsd8nPxMlKlYy4IJNU0B7lKi4/NakE6q59RJB2x
AiljLQOZjEmTQi0eBVU4MrHcYTQ7tJOZ78Z06m235nvdv13GXSSGRDwCM09Z0gE8
vm8/fO/F9c1h8kkwucBf/f9y1qCG1eolNKFSurrcZwH3OB+WG+1rBfz9WfPFcbcR
OaAX5pR9d68dVlmDCYbK6EhxuKESrXje0rqG3AZfZ0GZsXiedWEvlFNU/K5YYiS2
HXd3AdiQ+aQn49aah7LbosS739g4tikWzfC4O/8ZMIuCyoaQERBmY2iKcubDDQoS
bQvuOjvVbj1ZAmVKUyej9leRbSCsOaTKLmfAj6XEUZ0+zDmlXmb8cgLJ/D8Cluty
Dee56SBub9weXL+Y/QorrjgYf4r5Ciq6QONT2OHTjDPXv8s7ToGui8kT6CMnpgwW
KsVzinOjyslU47bctOcFwL0ddEoGX9OLe2D8XLUMhPAJKObFylCW+vWqpEiV35XC
gr+SBewKOTeHxrtD/EjcyTqsJanMZx9yvtYSL5u3aKJGy5QOed9YuqQBpF1Jm6Lq
7UjAZDw5Ddxn6CNEF+xKjjxAIYrXfXkDODlF+SDbsylpMWB8fW+MuvNEZgEjawWu
fz+ALq4Tmv/8i0vjG0m5BRDaVE7P0mW7SMTxNHpdUkXi5tg1i6l3MdIxnhMKjY7h
gkiQE+WPm3NoCnqkeRM2vYlWqTxHFA/zBrAVFNP7ZYFqYmHCRmy1EHZ8hP6xT8Ma
F3E9vFVuzGH0bQXstKWmodq0S2QKwfOaE0eUtUC0ETZfTKU6FiNJS/HNIEP+bbU4
TqOVZMVLupKpuXpWTBGRYWPL8u4PtxKxUMIBvf4OP5HUQMf7va2uS+/nY2IoNIU/
O/RHGP/Bz+DoTk9MFcUIKmndKRR6IcCi1aMv/oJuAXjT20aFLJnJyy5kjJ3QMCLs
TlthGnsLaFn+USKEgGHy2xb3kX4gJuJhvVoClWjIm842Cp/JyNtc1SeoUFJRpABq
KuXepb6fEl+enIFvUHLh12w7hFBZRhpKHgeSS5aCB/hqRhoJyp3cSYollwN3gffD
U1zrgGvd6kVs0Wi3z+0vCulnptQqaH3/RhepaYMYE+sreE7Mo/yeCHa1hujzmHsZ
OCtIOa4R8hocXGGq1hC/gbZyrp2Cf5ZKj2tD1jlzFIvos7AG7qAo4iJOUmt/ulpi
zvTiNK+K1dK3FFmw31OKdgDWs9zIYQdRZXM7p8RIt6TC8mV55D+XJDfQ4YAUi5M8
JWRg6IdFxbsil+S+t7U7fSQmNqgn6HL+hwyRNNYXnbG+c8dM6YCcFfX6qnkfRObm
ZxaliCvbH6sjDrZgdWJDSrRvIRGRQzWBX864HCTqxyhFuKZdADum0uQeZBkV6Zqs
oX8OnifXmD3IGLl5myIdArMXLyZxagXdMU8wnOttYsefsYaszSZixnROEdPPGyN1
kZ0+4wMH+CTpKJvce+JRtR8ggEnI2MB2HGiL/lTv+gFxATpISiy/Xm4HtJTHL6bZ
iVTT8LW9KX266JQ2oe1hTrwGiFSjVCIqgewxuQbKSWZYAzN0aTKzLxwuKWh1Ior3
TnoVqQ2m7Qzf19bixGkHb+KaAD3LK3OGHXwytdooRcbvVORIRhxtugUrp5271+sn
L68kVfdoaEI4VuiWNwRfUb+F33KkzW4WfH/wEsznInL/6haByhZBYzOz4zO19syZ
UScd0RH2ARUtlrOIEcZq5WNSPZ8fhHLtA7dnFLLQfyemhQEs25Rm+/hKTz7gXbC+
w++X5q7IjwSDCkoC7eieM67L0PDFj4vZDKWcNMtD7SAXuRN+vumlx433f6d/lPAM
11PPntH7HW32EIgYrWUaCgwCerwToW8ls7tJU6XE9oZek7uHXDKV3OaipWi0gcPB
ccG+9FzL73GYcQSWm+mS9y0c7P3OVNTO2++z82Dg6NarLizS7Dv091kdU6ebbhl0
qz/lmjrH0PbqQ2hi0CqUrekzDQJ79cUizirN9mDFsT9ypBAcV6XMW9FJvnH9pqRN
H36R6EjKoh0ksPZHtLrDks6mcnqRx7Nog5czbP7JAMBJEqOtaGsaK9v/4gx2Iuy3
bvjMoGfkCPlrVl6ftp2mwNs14dd/10o2no82jIgAUTg9cJjDC6wvy4IvX7vkFNSj
HOnESa8X6HIfZv6TXfWmsX+o/tRm5oTlecMJeXcvqYqDBu85fYrnm/71ajdQxHwX
uvE/B7iNNFgpfsoen7McFrZM69JZZ4f0PI0DBWELM9fOnapOo9MI35cN0SMk6kD0
wtQQmemL3XptKejrIyTl0ajzlKj2weLfU4/cOfF5q2jBRjA0NHBzGqJLOUExbXyw
aT0aI+8SkB55knyFnZz6JTSvB3UgogLl88fcVTIjYLwzJm9tiV1qlTbfNFLdqIEQ
7rIU7PQR5wIlA1i803XWA3qj1tNeae8a6W25kAaMan0=
--pragma protect end_data_block
--pragma protect digest_block
fuviBSIgN6YcNYk0URh9X3zzm2o=
--pragma protect end_digest_block
--pragma protect end_protected
