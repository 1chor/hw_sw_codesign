-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Nwyrl58lQMIuaG4XxeXBwwy7C1zZE3IzAEsrQxm0njcOBDSeQk8UvN7nCaX838hM
QiXOJFGf1Mk36Tva16v3QSkkwCQC/SWEgE5RdcDcrEfCnsy3cEKSXtVbdHPX50u6
4KLGrDtFv2/J6h0GcvxlqhMEEyzYsukcdjovGnFYdIo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5120)
`protect data_block
ds5ANiQhbbkgjE0lne+1mAeN6QTy2G/lZyEdRS5/ob0zrPs2HUpo66LCWQ/Xg/ka
bifDb86gv8It0uqptOlDRjwFjX+VEJ+FJkR964gyMnepQ6gtg1X9ktJxpjwk6wNZ
H3dXzHfDvnF/jSW1l0VeAvCYZIZw71aQFk04Dub8kvLxzoacKZq6stIVLOG05YcA
9U/U66870DafAMT9GdwOMbAbcpMzDyUfAXGmVNQY84/oDzTXpEq0YlbbOwRCahbK
1dXDnKDxNtyR3yRJJBFabujJlNXyT2S/paiKWPGzNBidec1hTliZIpTAjMolbhoJ
8uvcHkMnDES2y//ytzp+1TDynG6W4HNgZQBJ3bi5Z4PFytn3YhWUrERrqpO+NbOn
BOn/xFAOxOYe/pF2lwpB0vkLod5AtF8w12ofzlj8SJnSyahvvmR/VKbCr1VLCKUz
+gXu19Guer3ykSRcv72taxsrA9F4p+jKwe+eX/kF58eBm9lQWLUp+sJMKyJRA+20
B5L8w1+1MOE6O0ehfxi6pJGXTf9YACi1fSdsYKs20MYeNqpBu/6Kcswal8pDFX+h
SXmHs/C7lv3hQWFSJd/XGai0TRZi8Me2A8rgvFTVL8xN3keu47r5Gpq8JBOKd19y
Vc/pMqvJdvBCGSKgsXw+duSC9e012DUyqOGtHpUDuUMA7LELGoZN9itI8I4mG0Y0
lvmzlkC0APr2V8z1VLw2VyY3g/DtacFwLzvkmWkfNQJxt9PK0rWDmDuFtl0MMtGk
cQnWh7tvuWLPrgz0vQC84fDPiqa0A52sSUlrkUMr574FAbFw7x4qr28ik6os3jn+
elBDvNsmcJlWq5u2072oA4UnXcy7KbpihWEJzgZeySRmetQcCi6se/GVhE+7Ko2A
q08SVOg6X5uXTYFnW/rqj0PorjNxkllzsHqihAhy8TX/xcPd5o1rT0W37uafjG1D
Ze+9Dp4GXllY7K8anZj3Hvzgrt9lALYX89ndEBGgOGexsUBqJpUxaqhx+vWnUYTU
YR0H43cUe5VBuQ4+q+crX0Ut+QDKRYpEnF7xlsJwBqzqWsTy9ox0tgfERF1F/arA
2p5XWoZqOeeGg3f2N3zRZcsBdw5a9B7J3+TD8R8ZAPejkF3uHjww7pji3TXIEq5L
VtnFEFoGDkrKu2cSLfMPYY37cC6m856YdHiOBWcw1n7tXUbb8eft10gPvn0pgO0o
PqDO+3M1qaYRv4vZmR7VbWZ6D59k4G99EUL5TpCBTA4wOzMQ1DLrDy/t2q+C9RvP
hfMhziTYJYrIj7opIdcFL4RoCKsYyMb9JcLp97iPWYcTt2LjhT60p1TWab2k/Lk/
nFcwiWgJkJMThTyFYE2qsXq7NHXrQG8SNtl+7D8EdWLUa3uzD5gP4n0Q4nmhg5X0
nKLWgq/V+E0T6yeAHAdx8/00/WmD3vbdhuHibvl3YcuVmcnJ7W315uPQPf9pfKpr
p6DF9PpWSuu87OClLzq2NPPAOFCqlq8X6rW+NsUm5Txp2851BpxEP8sB/nnjRsrf
uo74UKT5FgDxRH6XkS1JXTGMxUfWJwROQbLQvJzFjkrifxvhunnNIonIY18eVVhV
nonmyp/VCShhI2zM/F11RVk+e5+IraR7VsISX3OIF9UHLJeaB+Z0jv+AxlXlrZBd
ZfoxO+AEQCOApxi7r1wKISSlyPMZe5QUapx7G5z0z3zpNoGj5Uoo4s0UBnRhPTLK
hZqFpzBgbATw2nZM74UNTxJ7G0TDXYAMjDpUwj8i+z88+Mn+u5jJgqY1HDIUjO8f
ET5SD4N7B+p296Ndr47QN7xjUjcAJ/9QuD7CNWP9BzkpgSOG885jPOa7wEHwecm5
ROXUXgjDepkRFAsLeppUBIZew9gBgTtf3zB+abmuwCbEeP/iNDnLj7/EeSUfSP3W
VxUzHPiYPBq351uWQXOX4q7dNdqWCQECsCgMlfxWkg2EE/wGiXfKrxQMnQZSCUq3
+kGUQ/qYx+A+DAJPvD33ZgxS6gTzlBWzP6gEVMNcOa0SIMqdy9h1flApHQ55C4sy
HfYSlUMAZWLUyD4mrJBM7IW3DzI2w6n4eZbDEaYRoOK5myEOOftvES7Zpo7EfRZY
68wSiPlfEDnHcGyZ5Uzrk8OcZjQf3+eUj2xi0ON6iplHy1vlHzOWdyIboa0DMZea
/aAnFWREDxG37sgiKD2Ihx2VSa6q5kW1DxKh7Kk0xOpmHszH7R1xNniQ1SQ132Dz
NYE5EzYcGUeMnOzAelIw8HyFYsdt52nurzi+I8vIkhhDNxYcaFmqVXMATxlvRyVw
Eul7Pek06EhzJF16z6crTMtXIPH4LK2OLoKmJ+lNCdPgvFaYqmDcSdETNxEewpXx
ewhl49ZvJbhTDJN9fpkq6cf/CINsEBCdRimkYv7AeapA7JpOb0toNvDLrDA4QMt+
FpwLT/RozjQw4M4qBp70NscXfNABDs0SootjfTguA2Et2GYbM/THiefCX0wr9C9C
XR1BTp2NgKhLVUt53KKR19cCc8DoT3AThsP87EMtqqL0SVZNAd+GkAoVWxxFupeC
N38NVjOd2aXNHi7feqMZ4rJ9W2uboeHJZOuhmzOYqfuhXGwYdqaPTGHyuoTXU9ei
cHXDAeQ5wM0VPEgLjK1Xziv/r18cqNNsNaybP5wohwFh/hBHzfnd5REUqjbnurGN
CL6PzmN6BSNc/At9xyI+zeZZ/pp+AfZZlVLJ2lzlUUqq9Ml/1mQY4HjBGElH3tzo
l9unLW77NbbpOvKK4Q8MxpUxLeEwDUkswWi9cfvMkQsNAgeJ7b3VBib2v4Ia0SA/
EL6I0lFIc8u147EyFEJHN2Wp6iAfdIq+Fc2iFLopfXwbfjXyYuCW4B94UySwazf0
psrFLvwgPE6SOTYCl4ohKS0qHksOTPNI92XQtNX1b8x/Lpj1CFHo0o/1Wdw1r+z6
ZOjz++/erKbAHkuATAgjXsDAtAnYR/3hncNeyPhFU9Kzg8lp7iwYblpY52/mJgAl
dekYoWlK9VQzIrMXNHjZw+r406SxjpHXeN+dPObFIg/UhpYoP6b8Nh7YSUdAxDRF
LG02GIJ1DejytjpDDjgPmt0Eb/J/ind/JV4JM28V6EXtn+8JRo0A8EnI2fjCiLWd
/Sa2qPv377ZguRqGmmVSXxT6xHwM25WBYqnO8ZMThByvfEvX0XCirR2wBuFRRgJ+
5dLCLcqU90uUPw04VahB/CGgrsrn0Y3M5ENOAguWMHQugzZPQee1kyfmEngIbr2t
M3KJU0uR568XBo2ohAzVGKcmyuEhFgJ4/gatEbvnQ56gr4dkRYOttvecskItyVfX
e6NDTk+5UE+zb843x0ysaWpMP0Mj8qBGWKkYjmBUwPr1H1EidZsUrVBkxTmGedMM
bj9QFVKf/y3oSysPcoOlRyVdoVd4HRMtulZfuHLcqOhrje7rMpiXhCsJs7lGiTlV
LResDVz/EVXfJybUzXDpzSpA9TKGnPSq6eMAOBIq3hTN5M6ItYxQyyBfJwlfzDoQ
tzXNmDPFstrE+gSAuZbf57laBFoOy+wlOehSZszw7p2QZnvCpdpZ4iDsMgj+yldQ
zQvhwFGSKWyzcU58NSxpahnfRcAHvMBuD8FyAzKd+/WoQFJkQ27XuU1/gjeGJ+e8
b4kmkKl58r8oxzeBv2fCi9Gmc6bXvOnk1BgIH5Pb1ih27lQK2MGXIYPXojhORNNF
TVYvCO3/ZIj98xfwECCX+QWN3TalLE9+SGmAtUp0Unb1o2ft35i1PLqF4SBgaMyr
vYktNhamH27XN9Z52WkZHBSSsZvvunoLj0wkK1acqTU7wp7gsArg8M/cog7UQQeg
TC3XBbTLOHMf1HPyWWbgEldY7y3rq9XOTDlQEajmSRV2Ja13gbfqrxaPrFFzv6FZ
/YmaIAAhDMMESnCM/6yTbd7mmiJS9svBhpa27SFxmHyZhX6d0Dv52nRz2+x/4jpE
oYlN0BX3jGL1mW+yrCv69MT2uegmednVo873TEm5XU1VDFhvGvrJTqdceMYOt+Gh
M/Bn0OJVu1XtM7jXrZ58lAHHhIxqSuqIfWVogURag52EfSvAjdMQnLnfTCeXW7gh
/ijiaIH7wnxcFc5COG4HuYjKsJqbGfDKODTXdUQAg7rKjmYlLZkSjQ0l69Och+mF
F6zA1pKc1/Xotf3CsmVZXdFGHo4DO/izouvnW95m9kHYOyBUuYg2rtFotbePKK4q
ClhzRzgtFi4EzN1v5v2B2mwEiFaxs8XQHaj+aX3rRp6BHQWpNTqZHA/Y4IHSe0aB
+n2Ul3QalA4/kdpcxGrcOBGQRk79/ZJKJkv8zNqx0i93MP1UBaIMJTqju3sgMktk
mn3o6QfgsIqCS6B5AzGelxxQzTywr9xaxMiqtYmci2xi7MwTyFcbtyB6SyzjKTRD
wmrFI2rUS/LkmivP6t+AfVkWideX92tsSVOqW5WCF3Gwrg5Fok3opNZQ+qpcO3ZD
DJz7ZgKe5NjkkoFfM9U7heFiqvzKaoVKHGwrdKxecLi8o8fLeMyYFz1KHMrepKkA
aibsissCY5nxYJqutiVh1lVnj1LJfE5PE9T1n9+HA6+SnxUJkCX/q2sq3Qz/MNi5
BF34rIQbSwkUmJ6OAMPp86bsBubKA4xFOjA1GcgNzpn6SnACQ9V9MUwQhw4p+pu0
pnt1crbD7YJSj77L4PUrL4uY3GU/f01/nXsmfEXsy9/8ReNh1oLqWefXi+miXZrC
8RKU0iSOJvhVueIpGViViRMYKM+11R2T+a344Ive+MFLMOW75W5QQxllipmml+bw
AN1U5pWRD/T12RqQQ/II+Nzi5WAU2WELClF8EGzESj/uEZkSeCH9wE+YoDz7q8V8
3U56WXfOx4oJPbV+205unSSSoIKp8Sd0pMfbIfGQrnc3CITKLNjANxiA5e8iJ0gS
CvrLtwp0GLLTv3e1ghfQhekduxWhcmbUCX+LDzWnyl3kjYLqc4ziPWgPAJbRCs+2
xiuJ5KYbQbEqdz+Uw1rnprrWG/Ii9nNoYx+et+yr1fY/TVJdAIubyJ4Tj6wV+thI
KhyLtZmyN6qj343Fi6UdD2gfkGBGyN73SIVoajM1n+OPzM86kRFCUWjfQNGuEplO
g6E82yWe6zX6ijbzIa4Wq3rYl06Wu1bWRw7rVNBPyKx3emDoGbDl6+beq5+ErGNm
2qgqdgefTkzAdJyA3nzCco9qPfBoJzsNSp6sgPB6Vn+5XJ1DQ6dfCMXwYjs0n4eD
edrNCjAAvcN0rvTIt2NMAxBCGBOIvx37RGbM4JisjlwAbxCevQu4bqDXxePETMB5
TZoKi0IcZEH20wHADq94DHWwocjiAR0OPViNc3Bp6qmHqUuSA1Dk/8DRwIK9WXez
7pvdZont58KtGY0ftQOop7FfxQC4bYwi2xBjO+0BKPeG1v/zg/RiGFKz9tX/QIep
8zs/vFTj6z1V5IXAWCcfcNTD66jKnzSzgQ4xlCa/+ycWGJIm7wOtv+Owt1Q4ed0S
OtsRoBItuLuIzAZOi4xv9d6mEljiImdhpk6gCb2jPMucDKo4J0eu79QnfVTdGqJy
i2+1wOns/rrRl2R5S21U5Rk+31mqf6tXbB0l/ntFxgPXgn0JMCOY7LQb4nZ7I/AR
iFi2rxXpgdM2AasdVDwnhRDlxSoM7TfP+4w0bYMK7eHGx/bJbGSn8fkdKUI4s18b
eWQ1MW2eAxgf0Hfl2p/zoggzkU0IShytAzl1iKofWXEFSo+uH09RdDJV4crGOywP
bcJXgs6ZgwXaeiazMiJjlzuYlAyEaYyb3IoJaGkrw7+V2Kw1E0CBcuECHbraiUxb
IXpiShB8VnDzFklsTxYwZ8j3SBk+TMRZ18geT1vdljO42xGcdGSGb3trr1ayAo/j
f9cJWKKezW8clsl0B4KLXyAkOTsCxdC4q/qgzDDtON9EP4jNaS4pg3wHsfZnQ0Ek
UQJX2UlBpuOFfON8Ze6IiwWLDruvdhs+/YwC2oSMPBcmfXt1h4LrsiJ+LDYxrmWz
gGbqFuJb3FPHfCGIAvC1rJ9guxDZu/bW8Uhyw36h95bYBOKu1Qqj8wZ1ZfAtkppR
5uCHbqxeKkqtXamp0qLUq4Hv7y4+NSXw5hOIKlOef7G51LijIoulGBlkB1OGn2xQ
aSRI31igPbnmal+dBbf6kkKONKzLNBNqbv8aYJlT6KsTYAGLxJbtgfgb68qxDFt0
seWQbxeTQHkqm7u+bgc1KubaDFeK0nwLRoxow8yWo9AHeVHsYcGZ76jDUgS0ThiP
kSG3Je1fyAmBLSOKCIgjFu7ON/uNhv+ueIJPw4ihdg5vWPI5AiBQbe9kipMicAnJ
+Nus2zGfkfeGBWRXlkuvdC2O6KJ9oVUZwLdcANzeLrHFtjZAgOFRlHLAcdJVFl5r
gR5RH5K0v4CWLetgOMpRhRUiNV+36TbLmaCQcDVmh4TwV7/zBZmb3YnAlByI6FLe
ndsdqjtF7eYGmC6mGX4ewotK4fCWtWwTUWmxj3BT4D+bcO/lUL1r1kxLR9Y+Nh0Z
dh516rlHc37VWOIc9NL1R5kR3rYNWQQ5PMB9VpStTpOv2k/FsJpf0Q5/nbFKHLl8
uahdBEboHhh438gNap3HkAipPWLSVQYahXmYmPcahy3MOoAaesgnmmMWcZg0+948
G5XBJkiDNeEU9Lw0Vytdv/ohrCycVeFDJebmeRynBjcGr7R7PfLIGo6b5y7sZGo+
KupYYw9Ebm9o39j0DH5CUdmOI89IC5BmNtyO/czuArKRI8K7SoIfAJaq9kXbZUFp
G4RW1cJSd3SU3FqjSalcsM/asleP91MtBopoWkzRDT0=
`protect end_protected
