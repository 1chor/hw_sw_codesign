-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
g6MjY0lKFKoKMW7l0o4qYkA30N7Yv8SyIx2R6B/RQ7syCVtXVoVSUpnVtQUMFn3xgnOuW6ACNndm
xQ+dyXcm0uvf+r40R4OsVU5rxjxOD+GtI9HHHAi7g52lCp5SVJk1fayWzf7RAZyQmK03CSbUg+Yf
59LcWgGSI5vf91UKvj522MSv1qX5PbnyhgnS5wd54h1/UlRDupx6JshdeRZhPLlDTlLL5IgWUzfl
iFz0TRmy/ZcKjVeF3Qqgw5zDUtNt8xrgVgq6CEQLmLElpK6YetXXaaPP9GFEEemB1xn/EPxTV+ab
YFKiu3hj8YhfomiadNR4aKj0U5GKUtJrXnewkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12000)
`protect data_block
DPpUIbmLGy3mziHriOUbsa/h8fXAYotYqhit+VeBFakbFKxR13PlTa1dMwYRUnuSZtMP4t+HCKD2
3k/loJCaCBQw8QVe7ymmK5TwweFpUEvITxwtKt3Y4MNs//V/pTkVH6tmNKKcb05dRxJbmpc4u6bD
phJwDXk7XMj7jrQAqDUn4+BBSZWM1TV+ixxBuKVjpwlEWvlJFcmap2ivs2PonETVtQ58WsfR4Aby
p5qvHxwXhWhlUZ/jStIiuk/oMGn4qGTDM4tOPAPdog7wc8red8EaxpLOfyxz541P6QZZwZjx/dAk
9iXPhPAvDou/SOO9hnrKo6JcJfBe9Ggw49eWWgHFQ71agbojU7506iSkjwvaXSO4zEkNdwyHvFrR
GF7kqcfqORa+8BCvW8PSYYiBosNPboTukq4vWYA+nE12OPllLo0ld/yU605yUP0TgI3ycVUxC4VG
iBQfy03x2sYlc4yPUdGmEkwAkpnIVy5QQuR8JqS2d+bAMJskErRbWNCi1xXojnL0SKI35YUF6RIO
afaKTNI26D9pPVp+ilW5TxNnvELgk5mxqCJaTirP1CGWm0YTJhjA0Ny8+CbG4FpQuOGCP2lw/TmD
tY9g8whyVfZT5vtrKoUtEY3thnqf3rto8mSulQysMoafGGInKaLcbd9GjH5XixdhiYKC5pztSRfz
DezZMB8kMS65dik75RH9USS9uzEy9jtbWpN0hRTadj5UMrW9mnWALZjwm1hCt19EptWBkdwNFDVo
2s7l+M6kOxP888mEnZ9CtozD5y5d+BorJawENv665h1odkr7wmq019PpmWMmcdu5E6DBd4iKgzma
gSLTO2RJ//0AkquhOlZsR5vgQkFAUReE0670BmgHphS3R4HbqfZ8THuOMYgZnP4eUMg+oOxoHR7m
pOlvsd9UrorLW7DIeBp5OEvfpGTQOXEMXKUeLH6RwUeLMX5aA9Qm1DbBIbQTfMUDGrOnYd12hm3g
Y8mSKw3zLh7Ixxkm+Dv320HlNe1WDDbbKRoSXEhT/lELV0/43DX3NMU1In8XMvQ8bkOOHMHPT6Up
Qsg3/xuKoKHypBsRAGHhH58OWp1k5H2RUtc8vd0iaShsB2FDUcg8v1JNkz5FRDXM4y++RgYX43aG
cIg/PwVvTc0p0hwczyOH7f8D9nYrOiIftDbioPhcNFV47iPbK+GeIu1W8uo+X9NgArwZblcUX2UP
ps9emw482dWQuR0SoeRbpd1v/wLCtgyBPB1wXA7NZvznUsXxz932bJrjsM2HknZhoqdaIbIPoqaE
B4HBqPJxiNpUiyS2LpliiTxjv6xN3kV0HOK7LxsZJhR//L5bRac/DTOVgmt4uG5xklCpj5QwDZHs
oUYyJi+1DYVoOkAxN7/TEJALA14Bb2+dZtBpPOZSdTmscOe+ZPdyU+IDflbr+7ALN9jq85e+Qawb
NmmZmhbgNgRIKGk6UwOyvnehWItEeNLtjjzKORVoXImKkJmx2+9Wr8MlAHuRAyWHidRLSTXd5GPK
yXhLMLJsa5ocFySdqHr91tGQ3MOY9pLQFtcZOFXzKpaqsLCGW2hnYi4psMfmkvAiwTmrXFlI6kYc
CtYkurn9/9kUgb4Nf1k5KhtRgtgGGl0yswBqj9wQ/VA2To85nQOoWZ0SCiqEcM28rYLu0UXdNmVv
8PuZ/T589erQbSXHGhLdl39Y1PWpQwp4Zyt2SBFBckK9vz3Y1r/rMNp+zAwqYr6ASRNlHGu/7upc
ZUXAIcu0NxAcsI/x6dJi5347QM/z43yMNSxORypuu7rkL1eu9wjGFFA9yPh6Pdut2QM0iDSkw581
vkdZzCHQMfYaruRS8tL4Fi8T5CxBHTGJGk093uQAZMfPGyvUiYmD5Nd3OJDxVX/VLJfqfF0idA2S
lY2Wq3GDVljSKvE1mq83XjTjiOg8xA3WOJ8EWuLcELVLp1Hqd13a5aG3ypFoU4T4uuHjRnF+fHM7
a49KKx79UPFnkqTWcyINvwHKueeoj73OlwvP+OVhzvcrr90ymvdKO6LASUF26i0gkPvwsIY25MC1
Y6CfpFzTFvwGv5pTUOx5O/yKU9DQsI4MjX9pNgX1cvbteVratNW1pZWpePwiVLYhsDpRO/Z2osog
s4iIDFK1BjtQ6Sl+sAdGIKWxCTCFlPbQCQzbtxWi78b6QybQjUziXkcHXpz2Px0R/AL7SCLCIuZr
8Sk7luD3fbcu56qWnrKbB5BaW8Lo4dIJhlO1l/FQ1kRXCmgfJgAX+J+ZAW6hBb+rRJoiWCI/HRWQ
CKG5cRCFiT+eTBI3rg02hgyhSfm+2Q1m41TRASsDTQ2V9LUxQkzhPg6oROllaQ4WatXEJDIrGwEL
1PlLkInXqQcMN/hUlqc9KQaqZ7Wo/3OFk9KToarMcaypsIAXriGA72CPz/GrHzjyKu/qZrrYbxRV
4FgUTj1h7Mkn3tHetQvkzNUoMqmZOr6tQuBQfkUvSyfgAwzEPNLCIUmcJflNYm8vUGQ1AHGWVXpS
+NyPXCnDGjeXB5788EPkEzWIbFk+10T9uwAFk4qG7Qrm6pLRAWcEcV9SoM6kB2fWEcp2qEMJoOO1
7EJIPtVvF8jzZm2/8YYjwKCsK3bKwaEsmPG+4f/NQzZX3aFSNvkqVrwZ78iUTAgXd6XUBwoBKDpv
v7Q9UC+WI7Npv3UaZ7n9t6hQEFl622lHnnKSfOU6nN22aEhXZCTRmolml/7rd4Ce+40kzasB8n1L
5q/uTlej0RVa1mNgkopARIn77wAeStKMFjtteIsf2P8gL733YFoHyu2ZkZR+ndX/5sxxSAOqXzau
358c9U6jjhLu2c03Jv5jlbYiVtmM84O1ZMp0OCG3Llp+QiUFoaIvRGpLRh06ERKyWUguNu7BFS3N
guoMnurNrtsWZEc4uS0J0NcPWv+AsxWlgshaFkKutTdOYhI66IyubMD4ao2Ikr8abAU+FV7y/kK4
yOiAPuKHCJHSSoMyfK+VUCicpk9hMvgPfziNmRadx9mD637lMbwmHwp+cuT6X7Wr7DSvM2soRbUS
C5ZdlC0FyLEBmN+xyM3jl4gM5RFBOw3D3aA+IVaWqpIttU67f8xncmbgOkW1OHh3bUYMDBHZAGcr
ReI9+3nuzHzemiEkrcdRFVV9EIJ6ysju2Dkt3mzgLu+eofV2ZR2D+xk1hwkTyyszD2mhKKcN7vSe
Haxx0zcg83rzfaVkpBQGuZMS2SLdYVY6UILu6IWU4VuUi9+qOVzOn8TOgz1fxxdWyQ3/KOPsMXU3
q+0Eh3hfnKdhiXlH0sEeWtZjY319N3Y9KDqYcq7egJ8a9sw6rcF1pMqfL0QaHOcR5XMCHBsSA4Sq
Iub8f07xi+2fmCiwZMohuU3yw6ArBNy2KZq7Y5PDF6rds3LD++ntKG/h0hEbocCHo8kW18RfcNYf
alOM9nxj5Byvo8evfBNuIFeeO4CFxT/IVywEdaMVXkP9yt/CV0T9Car1CYEmL4fCxrJV4sgdOalc
m6P8YGeZgoZkBapiAw247H2QNk/Fh21IVOM+0hifwVvHugmjwNYhkYFx9gkwSjfHTcaVzj2Q16/6
v0vfExfTfnSs4gGRz2e1mMFRuTPWUHynmtMhMiy9RieHbhCftKQ85YfnVw9lormPEp9681A/Wpvq
OH/n0v49BAcqPeDGpIZqfn0B7FPv1IZY5LW74g7Eem8SEGkHSW4VR9f2HXXCaRJAEjQe50a8Kn9L
98ecSxJf2lTf0NPWxi4C3DZv737tvyLiEBbuS8DDzfCo74wOKX1eiO0/0i0Vh8rSXFh139XPQMXQ
/kOo81mkI2pRvN00g19f1LNXldBFy9XFAbWVwA5HHdoJRUq/6IsaiyW0FoYvcXYZw/8dLzZ5qlrf
lNSVu6G+La7VLUaPYCIXqofA5ZuLRyM5vsetBGJgm8PPRmH2ACkroGG8Hi/i2lBFFbBWklWJXYYV
vzCACzlBlWU6Wgm3g2I3NZXndwkbaqC4lcXKnWrFBZgPqneRSeLv490VGVPYFwgKR6QqVu2qYd8d
3MpqUYtn6IYXq1R8/pv0B9ECzlvQQXQEpK//EvP+0t++gQq+xVITsqIk4BJ0Q7NrMY4lRDCCiwPi
ccVNCBBnUb/tOEk1vmMHPzGb0RiUsXT1YCKvV/FFjYzRWuontSml355Uj5cjFasA1jhQKyfMFBoL
qFQOaCDmL0uccRdZEkaDbQn1V6wSrefuasT21z803IWola2m+Ptekj593ZG4IIyLGUWqfRcgNYTi
lROVHQwUiLOu1vr9bvwCbf047kaaJ2misD0ufYTdiNeAbbJam5P2durbVmzo15WQnEZoaMNKeMTP
vh82BcQFTn/Hmy+TWKpG2UAWfHD+o0Q6w1OihLzyv6Dct6nfWQwtNZRtdflFEI8bI/ZQoy4siOxz
QwAFywPQKpXBpJheBSsKSXNS2WzO9fjfGHjNgHKYuHpvfNm59lyodnW2o7HiWqjU/INB2rW5VgFs
lR3XWIkvdj19lkfFQjEo43s3GJ9z2GYwzj8r2c0K069bO1vHEnIteN0SAbeuyCPoR503Z2s1OElk
Rog4l6rBFmPzB9xjtKxMS0gt82/cREQWsKRJro/iDlSF2UC+KCNkJrAg7bhJqAjxzGRSt0ZhOUz9
F2TJjyN/YTMyKBRNP3AuCHyBjw/RXgx+78XMEWBPTjVkhKA4t8UCgwsu3Tbvv9n8b/gx2DI8OfU6
HldTvxPpmXCArAqZgce4SrovkMloLlbwL/c5EXJg1q/tuezSJ5Dmbl2sTnmwAjwO1r7xBfQ2x223
ux222wAZSYydZVnbVBBmVJ17XLy6ZeeOS7EGA4dwkftxfGFROCEL4eO17jmoP/B8CDGqbncqqz+8
tDmW0Dcf+Ktch5NZkMBng0O4CCOmMcExfRdNGEYqIlOJEW4Z51N2DJb+6GyIYP324w9mDb0Diqdw
KsGtyoRJtVp3qFTM+6IMVqyyUoF81HZIj8plRIUOJw/uX3OJyJk3BU6pPnfN+hVKUO9f64tUBt5U
GugUHlgthJ2DNkxV3N21z9cLZXO3gJY2byscS6FiiPbDTOG4U3I7g510ldtuYGPLjBk74rU7gVVy
ICVrRet7nwcs1zTsmKKfFdlNuXdK85TRWsQ0OUxcVKFkMl9XoxCaW1fbYLbEJNNyE3mX4VjVypXQ
4MRi77K8Y3s2b/k6GST+TggDeUNN9ZpfOAhvp9cV8jNN40jATiAYbEHe3Y2qFqe+L27hJZDbn2fk
1iZ+LrrU9oPFYQxQqHV3pffd9kZ9TPaEai0vIY8OGxsrMsbsC2V4JypIJKgLRgMD3lGnSPLKqIJY
YAjuUbBhOAAJcQG3Ge74zUnLq1+nIeTz/x5bFqJlNOMt3LRBZS1s07IL4F0TYXc+/cYYqIcWph+2
iqP7ADrBJdW9oto2UnJ5x5aYHBNN8iPQrLDiTlXmEnmdGwwgsAFbca9Adk0l5KFfc4EaEfSQX0Fj
59R0vfkr0mOX9EmCBrvOSn6EDwPkr9yhNbiTpo5Dt44E2yuZKvaaHaPUG/uk0agWy8l1dAet0xzA
OYD19cf9pQBZVmqFgZaQzfr8wZKXaIASN9bPvB0IPHz1XzAF+TBXkGT+KyZ9DLzBX1U6avQUJ86m
FWWpxcuBAXtHjVVBd6M1riCYFTZo+kidOxoyjUJJAv9mhatIJx8P/OAhzM+m2h+NKQw6jCoutqMG
yYWPvWk0p7fQ6LyEXlJWkh5Nxzzd0B5AITb8JckHj2Nk5dvcuO5io4lYPxioWWc53FqJ0B+7Xgxt
r9mkeDY5ReWWCFXKMO33tmNcW3JVIB5cavaf8ZRIFL/EHADy1h0dFFWKxwD1/YkUcaaNPwC/BiTs
mHMXeyZPRAmIza3EyDfXqAa9QyaxbNYu/ibWp1YFe+IHj+XpJfl/rC/v2HelLktc/tZCBn/XTF8M
dcBRM98Sz8A2wVptbb8a30zS2IzOZbzoqs82tak8pZgOIrIl3RqJBcV+rAFJ979SpMEhbUbQ8/Tf
snSe2rI+kxjXYBMvZ9gVRmgeezBdf3QVID9WpCFo2EeOx6oiexPMH203VmLs/typThs2ZUQ8d2PK
I3GAQMT3vfx0ijTt+k4y5ldbrEpD+J7JSaR59mGzCobNn1wrBGZfj12ePuPxmq/mBZwcYKIkGQgN
J5UMyj4AJd4d6/5W6ISqRncYJivHYNlRHetXnAok71/kFC8lAsXuZdJnD/1OOWfgg028dV0+QZvA
/Btjwv7dEwpUGvPH7L6TN0RaxcbfTc57IsG92mWi3eYex3l19IcvAfNC2OjCQQsePE0PDfXf5z/d
UJKXPE1haDwfS+VuwjN4WWqr1NPDGRHZ5dFS2T+aGTDUx7tqZivvtqG+iOz1yBOgLLXYUslJZTJB
iF92NTzoz0vG3TNzESsq6W6olcgBKUwxOqzAauANzPgdXFZD2tMBFfQlEv6lbsJZfYeJRN4rikAG
4uoVQRZaZslBlBwq0bfxA3HLI2uAPfHZif3PTu428zg+zso6MUkLHLX26ET1Qte77LsZ+0EM7Hsm
pe95WSlQJyUHybCECZ9Mk9ECPUB9rje4TrJFx9rT82VsigMNUtNSI5iXUvmGoHdexNyNQK+pebDc
a/XhmgRZTx/fOoXoMP6fWuGIEsgfOjTJWBXmxyksst9NSh/tWy8RPx6inJyEgaDpY3dRJaaeZDIQ
BzZxw/Oas6SeMbeKnkzJLqungh0D8LnO99SbbiAg/yd2uNphwGV0LQB9AtNEeJZcFe4MGqwluxES
NRUZ2n8itS+8k6DZUxn7t3kokZEMDOJ2dPx5ieiv3cLfZqStQYW06dqRQziWSj/K/m4KfqKJqme6
y578AxqKci8dD8AKwLDVJR0fyImIWHus0mfedr6+HzEh0GeUPXuHyb3uXa8OElotHftCqto4vzV7
IHEZ0raNebSLyq3DznyNlExIxzueqp2YkyXGWYM2G+T1ZG1A9M2sd2NnfVsvi0AtPk9tbZoBtW0O
yx9dBqHR+w8BPOSFAs8QipFasr4j+rukZ1w4cBjXJ7+OqQ+etYqZ2oeUByngjkzL4GJgYthV32qc
8DcBTLYdUzNWU1uCY4dQjHwwRf0BcIRT1UWEP7i93mfSVfJJLwWui8gQ93JzfTCY4vsB+nm5EA/J
JB2osOspKDG+El0zY70i53NMkwiFlm0kxtX06hpLjxgQZrtfk0AB/3HgxmaI2OsoHAW45Koy5UoN
xsWAn6XrwilRxvicPOJ+Fi/NFZl1+jBKqE2vD9irGGeBCSAL82GFs3G8w76nMUcH9iV9UN2H22xV
A2YcGwXstdpbOjEVc2rB9dIFkC1klevLTysYxIJHa1LK7TuR3qvyQrzXwcuFaYbK0EnyRMTY8EoK
NqGAtMjNGmHyuToHMEOdxgsK6gOGXkEA++/s6Rz+T7wMErUrl3WJFw8KL+eB+ZYIKpC27obUPPPG
AvVQNjkciKiud+gpI9aTErRJipFxhum+Xa2KK6FLIGmNpH+o3VayH3ndKA4FjEpl8jCK3GwvLvwH
zSb+RQAq3/nqVmkW0Q5U4GwbCGsWqI0x9sl31LClaRgny15fgVqYr3daqNFlI5uF76Hy+o/QTDbc
UyMJ+cR9J5YeBSFfU0dPu3u8zs86c2DxKpTdEnpOQyB7giVwtJglhyqUY0xM0C6M3hKyCgxx5GRS
Lm/eX5/j0U0sJ+0LoRWKp95mjlbt6Ta9JIgiIcDgffZZx/xNseY90ydCIHJdWXLJOyXZwOWDRwQg
/Oxlhkj1/VeEqcnQikhJFROAKQeCs8y0aSLc9kE22gj7/SpjDz48BRfklv/IQkrZ+Tpv2UxAVJEO
FuzlgzB8hVcsJznk1gRj48RTUoEWww1/FLwAeGHRjm3NUv4l2L/s6of3yCvffDi5wPU3VwyL4MQS
Kb3bWb4pv4tGlUO9xXUVYAu2gAJwJ1EsyKA4lGZgY/U2nJ4en9VLLKsacaBzEIAOSHbMnjj9i/Rw
WaDBnjJyDJM6ujV8hjFlOM8K66/V0FbbeAWr+tSncJbHA2HoucCC2mYS3kHqenhqP1239CedP7YB
BbBNuwQNs/v9kgDe/rPEGVyihUjstYBPVRziLJIE3L59UtNkfcBuE5C8jMZVKktWPihbHse76234
a4O+Rt/K6Y0k3s0bK7UNN7h4gdtqPVeLtRpoB1VVwT0mtA4mBpVVS4We7E/y/wNx3lVIPfrQNRuK
5pTpS897Oi2JDFRF99rOFElA1Apx3wLaIKXKboPWNQ8bZKcWSbmMg1Ru2BPKYKA36h/xgGsFeabA
R+w7EvhLOZ6o/Kg7JWbP5bfPSWqVZhwI3SCa62n3UYQ4wohye+lSlVE4AQs6ZRz7VhvHF7cW/bZs
mUGE6U5M2PZiVQV7I+a0e5hSxqouVjnBBipQlj7hzU8Wpx809MY0xeFQjjpR5l+vEjwWGov7Q4Wc
/LS0buxP9B2SPQSor90+Ynq3/Ns+9tDmo7gomb46tfK+xP4kUl68GMYyJ4hsFv9zdlQt6qxhItnz
cPN+uZBD+8m/F/GkUsz7XvOjxHvISrrws23WgurUgZEdcy4cTL2/HiGNFvMsbxZMHQvSDQNJc03H
tNg5vBKETPyND5FADM/gmZhCSxvGRGh+IaOtSpESTTKs9SP8ZYIKNO456SFacpRtW/04L1BCqbQZ
1GAw5ulqwKbFHubIkD6k9PS2b1Q5BnjEp0IhHt08eJKQV7Es4vSljmMaJ2gI6xN97gemiQXeBy3x
2YXaH05ndDELFUYciBIKoNEUoQv9j2kf29GLh2eDVhxA8jGWDR4lSsI6PpXR6LY3CHQbUNcmSLL7
0KK9JeOp6WltsIBvcz6NmhqUuGU67Ce2Zs48g8Veby0S5kF+u9QM0WRtzu0pcYbFCr3AtOuuXnk2
ztAo+KzSoCV1A3tJiKx544qpV/2fHegkXArgPK3H/nEFuYmGgBL87X+4JIL8VvDPBEJ+4eIwbHYK
xySjWWkk1WfAXKr/ltTZH9w0D9EWFF9sAC7XF0u4Ak5wehhOZu29FONuS/2ZFc+aiKwy00pRRRUX
ZRupVQaF2u+5gn2mjq1Q5bK1WTT8jDPRdcoSFu5XdETBnnOsXo2PXNE4Zzy+L4rlob2o0EMIXGDO
hV8VVhsZIP7YK81IEURMl9rwhPTPAai1dz2st26daN1UUMXeQF66zksBqfOs8hE6+MQr3KsVBumx
O+4rUQxa1+BPSF4kyWymbt8suj2MixnwkahOFTZllKxKEIGDF5O8rYYbqMW4mdrC7xSmTiz7gwr5
lYDKgrvGyZVos0gG2NiTQ2IHIGgLzsD1/xc+eBAdJFwZ5naEGa6pgFEIYa+xxezYU30ceLivJOOw
V0ySgJ4CqrjbIFf2A0piHu7Yb/wl+NQdRfwOSbJ78vSGhS+eTrViUR5R8fQanoVRMLbMnEM4rUIc
PWow8Pc2w7dDZIlvhFWfAvn2L7VvFi90OwQlg4qZlRp/oY31kODH27T94/7j4wf1tIgdSKu6+B7o
vWWUWcNhXbPKHp1Vxv51QdCk2NK8A0HGLw3ZCajSdUiBxXIMoZUpak39ENZB48cQeTpjcxAhzzOc
94KIY9GAGeT4mo7OJKCi7uPeUJC5cvh7wxki6NReXw1zxRwrcbr25HH00jAMIFCecBc5ebmNOPhy
/S88tiY4uXNCPOsuYAlWDfwgwd7VSlHapPGn8nrkVJnewrEal1QI+ATQX1BYv/NiszqmjRTp9ZrX
1MMv9eSccK9lOk/n4KbeJ6PV3pq45XFKk+IMnL3w1nOfQeC2k8WRlkzF0BkyJUxPvxOFd5FwMxXn
ds9VxQ68tgCwI95tWOvWj164Vc5KdGWYibIx1HOZXgUYoh5/4i+p/oIcAix6vaZJU7YrWDQq8HcH
kftQnKwMjfRfhfNvp9xtv81rDVkF80lAq/W9qYG7Ont/+tnpsfsZpStoyUSQyNimc3qb1l3QSxHx
ruqPKFQKqnJyuwLP6imBldmM8eQYwvb2YMe9a70qKAcuuQuF46xMbzJIvG/q7hVptcovxU0tfwd7
RHguIIBHMA2hxtNPJxhF4MLFx6ZjRVH0tw7iICh9QS6XrRcRddkQ8ACxdFEzCPCrK1nxWc1jL3yG
lMXPIrxz8acPyL8ExVqL8b/ZLsmV9NNprdykEgxevVG8WVj+EX9MJApDyEnLD46jAS6V4Nm08fQg
BNIG2ykXVgIGJTVvpN1Dn+MhIdnXBPf7u+8qRZrhZ57JLS3H2rLiD/FTtriSFJGNBCHSy66mOJpG
HPpjLiz6TpZ/eGoKIcHEUp5UC17Oo5UgCMsIqfWBCBLQ1fbmVKbYcD53GJUodTkPl2HsWcKw0yt6
H0w6GfJLjJD555VaKz2t7mKLuqqnZcOH8iHPA6msmtp86TwOcSxUAEFoy6vw9ga8+ZFUQuieD9EA
25fIc4GpDSOdk9zb4JDLF50OkWYk0j+7ArxkFEPOO4KDtKEnZM39t7iRKXX8Umblpzt1/yTEYIav
dnVGjXmfg+upFuD7CkpbONPHxWy1ZVIdHw6OYQZl/VdPlGAopv+gfWKeUUQfuVNRXcRG0iGtmal6
wFeDljtBoBW2/UJLnZouX1VEw/dPzDWJ+FYiIEakzsgMduIqbNYekbVlqEVtMwkRfuMozbmmnNVs
f1IFwYtlEXqf3L89ChoE0wZaVNWNwWl4Q6be4maOahPxChI2+O2rIa/CVb6AxGPEF/JMjmte9CnI
tan0kUVj0qHMKBqSTxz24hNo7xkfjHEO1nNqQBpJ4HgB07ecP3CbT+jV9BhdhjziiFnqrDM/3Om5
iyjxsM7ePrINqcMGnpb7XU5g+YVTJ1MPNsG7XdfwpiajT3P/r5BOt3I2N5kmHASVHOlmhLGhGctW
XXdcilQyTUxB0ZX1bq3qAPHXoMvEeUTs6qDroqpXb6IrBlIlDcf8eyUslFYbOKcY0sXCMqcofiQ5
KYV40wGt6rqPbjCvxINnUmbeqkezxKPZ2oYOl80xEKyhLzBkzsejJezDo6PNMgNmNbcerLm8AVMr
tz3GqaulBzdMKz8RzM7O8i9DnCBKB+n87HcQE0928OXpnLgJaPH9tsnRCUHXfGKQBNe/6PR9x5iB
dm3MG+8Etem8MVHCWZFbP/RFV/E5TZHvkSAKtTb1/TSCWwVjn3p6iuEuouaRHRD/qJsbkBG6vKOx
xojy+lhQNw+XRuomf/bNhX5oAHm6brjODWWEcdYfP0ILaxTGlRJZwL2Jb2iGigINSDj46v/qSaJk
/u8oTUz15V875HN3N/Xtj0IzgIXBOySfTMfWYVvWYsTP83xla+cYtqV3AJ0Ld23Df6TBPNWvwsak
M4Fy5FXZA2x+nBNNweqE+buOoFqHm8UQWYBcG7n1zebasTuaYL+1O0XpYbLsxCDzcRwJelIfSW77
pftu3EPndbWpLroA9JUMneYk6QgZvLKSZgnLDHjP8dMWAgO3173khi49uozNM9SJQ5HrnffWItGK
QVeRvLWkdIVBTK+Lq35AQ9OfRsMtS1qSZ4cGEdWITPyZOqeU5ejRjMmIBw+n0ivQnQ4Gm5+eyyML
lTcgz/is67gGc6jvMS2ni7W2acD2vp09kfGF2T/SSvNT86S3U3LeFBjG5lP6xL0AAwt3cYE28R7J
ptbwnFVbcDXb4ODR0NL0QWDJa6woOff9XvKPdi3ltWigL1XZqxalq67DMhtpGaObb/105fmJCUYm
U5/ZKu1Yvu5rvPcEICHP1admE+HeJ6b7y24vbe6jllKdo2YEOGzFYaA1lkl3HIX2kOJUvUNloI8M
IMWoTYQysseyDKqVHUkcdBkF6Xgf0wiR9zCwfWfngzQs9Vx9YLIgE/5lb07MKk83fKJNPYmBc06/
Kion01P7LSq/VDHSQiV1zPkt+K+25db88wr6YT4Ftih1/26NWOM4a/+OLwDE3y5QIxtjmbR+O6b9
GOQYKL3SDVJOP/KpTXbhCevrHsoV4w+An9dVZjJgL+DDKpxEpcASNG7C/Lfhl7hUua5hQ2N/1nwz
zuljpfVtK59aKFRtcvDATaIqdIKQsjiTnINo2Xz4Sk83hjdWCEyW4828McvrgaWi01CAVthBT01/
E6LVHw6VSUr8YNBr4JEirnkyQ08OV0hK7pwvd5BcbLBn4JAumXZZHhCA9umif/DZGEdXJAgTTojE
uM4I62U/7zwS8+Rmq1FaCYXGmNaVDd5sdut+S8xYw8YKdjLpxlZwChm0jZdPVvB9pVwF2MEZX+tr
3ItZ2O59vWW3X95gZdakTaL3u2H2yCbo+r/kpn0i6HD4xl5V6aqM1heCvja0GDl8yKZ+uA0gN2RF
ZU15IifWFekJ+WlZr3itQ5kRso4pmTR+EX2ToDn4Iu8AcuqCWea/FOX9JsQ2bbvyAlKYOCKjIIcM
snaswR3b0eL/Jvc8TET+aoM9yN9oGHhcgIhR4uKqd11mJDTU4WatV3W1E/gCajeCsGsEJbYwtZDM
rFy7HcjCE8LTvTz8VTThOi92BU+9k+f2E+DYfy1Ctf4OZEjRsjlMmDEbei6Ogu/WiNl+4cDqR15l
6Xd0+5QoXhr9ajQi/DTHheLd0PKpG0W4W8Oy6LEUMKGkGZsdpwmdufvKEIytH63F5gjz2aAdS+CD
p80diSykcIfw/AIxjLGmA/J/xFm2425Z/P48q5q/tc9NH8c98E8yPO+wPYwpRuWDcFLIvcxG9L3M
bzckE89oTyg/KO9KnN8/+CAL/YrbHY5VWxW9KiXaSSWDHntB/hhNl0kx3OdLh0cKeuXSYdf0E2Be
a8C3EaRkWyUOMO0IyTBBFEZZUBqxnR0j/ZMxM2EPMcD5IEtx4VTXEdPUit40ahjGNGCzr3GwGdTA
OOXdQtqDsEU2UKNsGccd1Y9WHKJMSRHEuJDWAD1Gvb2czsex6u7vULvK9O7cX//LPxQEkdQWiBzd
Yq05y7cTppqqAL+0U+806OzwliYRyMXyolZEFcGM+IeHRi5HKlEWsJaleRvJx4xdE8FJHvlf9eou
F923x+qVPxKd53PlxLkVjrjWXGVEUncn7rnutnNzhQoE2Ov3l5VJDApdsX7Kd2ZYqgZzqsWt4YUi
UjWw5ngEtLX1GtF1+TJGlLU5BEbVcn5Xif1k4dsIawxpoUjQ4SsKwMzxQaPvU1B17lDwE6dRPtRI
gtVyuGKhBZpxsW8T54ZJLZAqOGwOCJn440R4wzUoss/B7oOaRAl5TabGkJ89JCBdLkYty4rC5bxE
2SMGkydkranu5OQw5a0LxtHL6A6YPIVgaVBFp6p6L0ysj9xb1mafH0GBbM6tZRbTRSzjOCnK9anm
VCSlSkMANd9VBLWO82BLbLNQ/FhOwVtj6eYlDpPaX315YaZoP4YBtN4wnRZwHj7HqFHZK269cBts
gW23wngIcbeufq311F7OC9iRfoEK8smhUo/vThKjoop7s0rc+mYuByNxOETAfHAs/N1BLimchdwc
tIcONsxyM2K2l7cqvhw86wMTM4PJyqo4cOToqOQyPO24naHPi+Rv9mQ0/8riFTOQbbEaYlzsc1aq
YSKtjYfAsP3ksffNF84exorKEU+3cZsC14qruD/lccCHekvG9KEeitdsPOMLgHfFZwqNj1MGtFUM
74d0ZJi7tSrorsNwvDDEWt4DGR06maGEXdGUtfsLGKZiB5wFHSWcIf7QlDZg4pbMsgxCvgtMhun3
zqrlglapIetGoRubrt5y/bsAgvyXbxviPUFUOrSImdCTpVcPH76+GGd94MjQuaa6lR9aY9cTocSS
Dz53aAPcoGIBovpdlR2+f9eMq9GZ5WzYkDZbyHg4sTKb0TUwK4TEp7iiZ9c6FUjr7AZ8slFpUIuw
PFx5t/flunP1y9UtYPgk+4ugyDyxdV5vAlikG8dJTfMKQlmX+Oj2mUZx5crAsbSYgljq2gkjFXaK
JfEokzxxoqR0/DRLyVLiOOiczONz8P3hgxuYLsGemw8PPaXfxcqK80bpg5q+wE68g9ZUnWdKYHwx
X+9XEH1L8VY2gGOmxCBuWA/nOKRE9RImyPicD54pHNYR+Jh1D7D/TsMMB38uWrjJOZzrA1u3+jSJ
LoIEJ99Rq549wjw/rheT739blbLMK4nzFL1G6gqAcxg1vM7zEzR2+uGNtI0X3B/3A/8FsXtdR8VD
us7alttii93bI5FLqeRTchwnrxedxSqDRJs0Kz48OVe6mszyStGAJpsqp2EUjgcT5dNk0uv3TJM6
WuMz+bU4SF+3s5e0VJ86xKa5HRXZcR6pFCcmGBNsNR5niHW+O5prP8bRosOgUfUFEESTrBM68lAh
RnVS4Um72favKXg+N7t4AXrMKFsoCEAmWgq3FuiK4wzp6TEaeMVLlbJtwvPtxsdPdUJo4OSN4tun
2L23Z8e7kurCrvxcrM72Hv1TGIOa5pGSPH4GU3qonPnIQE10DREcyKhu+/sI1KGjjCX1lKB0FIP5
VPwRBGcnCuf5JCLhsZ3MhxBfPqRu8XciJeDGisx6FHpzYMMQYbqwSywMXveXIc77VbhZbw1WzJHj
kyXi531KcAFwia15yCVqAxGfdv9od5aSPj/vKo6zrE69d4wFByXL3cPoBqw3sSGix/c1xgIbSpaZ
rAhJXExbWPFu+D0C1NM9p4vutSH433ldIADaanKzZNjvs14B7a0m8RUeAH+cEXFcNwcmH1Bi8Cno
yLlx96XRO5dKR9IAfI6kbmV7804tGbaL9jBTCqnsYwceWXN/PmNtt1v1rlztnjQ+Jvxzvr73xGam
rf8VJiSG2bd2zvJoQottik557QA5FcEpaQ2q9d3AiE7rJJnnW7LQPTJW1Bvvl+XzSzY+uvajUG79
rTqcHYQsNF/xM0pBekfHvPozE2PixdfAHO9LiWD4A+Ylq4Aebbv5hwMzWZrkVygmWruN13/szCoX
kn9YamSKskka7ISJUMcJMSnV2zM70WiJdmZ3TqgMd3i8YTFEB3VQzQohbbANB2/Fa0agP/ixuzRX
r+Rik0HQjZf+Y7ORJzG5lowvBt6Uj5W4psUmETGVjbuSI5q9MspsrrrAK6BrWvwfDbGp9O+BZ8rW
0gVzpj+a/biXs44G62SN9QEalYM2gfB4DEfcxvraQXf9ZVJ8x9n6L748GNUpo8gv6rwtIWQzsBFc
MNBITniB2u6FZEdfK5s5B9bufFWeTuYRUmIknZVGo/xEo9ooWIC6V/EYd9RpCP52ZZ3wAHwksUOa
XPVNXZOPoenRod0CgkbQD5tuidvYFTlGFusL+ZFNHjPFofhxA4c0kRzR9FfdgaLcEvCfqp5Ba3+5
c7HTF7vCMQ0l/Afrg4xUuEyhE8+1Dn7F2Kqmd9ahMOL649GRI1i8CTQc8uMIq85GH3+ErnMn5NnS
9nHtsCKAgDDBhkAg635qHO2b+ve0apWhte5gNUdWO8NalIPQIldghRTiz5cbSln2ye72gV0I0Vb2
GN7PrhR3TcktKxPXdnbxdaEgvIQDpPDcRIJmt3YanXUomqLJ3rQ7T8MV9YocS+WVATxYFfGqQYrA
aRHEN1ormA/8KAoxz4kNrxLbN+17UM1KaZHWhBfkahP/WAOEsfhXE3DtAjZP301Uuz2kwxVI6Gfb
Oo4UCd59eYTRhSCEbhd51+qSwXbtYIgGh7O0TDqerPt/tfBQPfOCJiYW7aiQ20JB9D4MXDbocToN
WUOTNDkith+U/AAd65BUOtvi3oMfhv/XQMDWdHBDr1I5A50LBMMjvSmz3qgSIfoy+B7SqRnu77rp
4v0QdbS5Ykx0w7cuJJTE49VKsQXb2vKcpM7i+dHzszT+5BvLGljYItWalCYjcZepbZIXanzibAsS
5n0pqXsVABHghrflvjQ6MZhnIyyQVEfGqxUi/lsUX5PueKR+CKmWhjDX6U2ek1YQ1AbDqpi5V784
9olfk+jZMEOFCdcfxuTNkwIwjneJEGv2XKIR1vDg6T1xkTxuPiygeW3bPPKNBWh+RJLFUlWoKc4V
pxfE6f9g5/4HQQRS1xxLGOyH94Hrz1TthmxlEMbg
`protect end_protected
