----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 16.01.2019 19:03:49
-- Design Name: 
-- Module Name: fake_sram - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fake_sram is
    port (
        clk   : in std_logic;
        res_n : in std_logic;
        
        s_address   : in  std_logic_vector(31 downto 0);
        s_write     : in  std_logic;
        s_read      : in  std_logic;
        s_writedata : in  std_logic_vector(15 downto 0);
        s_readdata  : out std_logic_vector(15 downto 0);
        s_waitrequest : out std_logic
    );
end fake_sram;

architecture Behavioral of fake_sram is
begin

proc : process ( clk, res_n )

type block_ram_array_type is array( 172032 downto 0 ) of std_logic_vector( 15 downto 0 );
variable block_ram_array : block_ram_array_type := (others => (others => '0'));

variable fill_block_28 : std_logic := '0';

variable skip : std_logic := '1';

begin
    
    if res_n = '0' then
        
        --------------------
        --=41
        --------------------
-- 			           c_h(0)   	                      c_h(0)			         d_h(0)		        	    d_l(0)			       c_h(1)			     	  c_l(1)			     d_h(1)		    	        d_l(1)
        block_ram_array(167936) := x"028e";block_ram_array(167938) := x"ca00";block_ram_array(167940) := x"0000";block_ram_array(167942) := x"0000";block_ram_array(167944) := x"fadf";block_ram_array(167946) := x"4dd0";block_ram_array(167948) := x"fea5";block_ram_array(167950) := x"a310";block_ram_array(167952) := x"0046";block_ram_array(167954) := x"45b1";block_ram_array(167956) := x"0328";block_ram_array(167958) := x"199c";block_ram_array(167960) := x"fcd6";block_ram_array(167962) := x"f228";block_ram_array(167964) := x"ffc5";block_ram_array(167966) := x"d7c7";block_ram_array(167968) := x"ff39";block_ram_array(167970) := x"189b";block_ram_array(167972) := x"0503";block_ram_array(167974) := x"fd40";block_ram_array(167976) := x"ff81";block_ram_array(167978) := x"d320";block_ram_array(167980) := x"04e1";block_ram_array(167982) := x"9cb0";block_ram_array(167984) := x"09d6";block_ram_array(167986) := x"e790";block_ram_array(167988) := x"06a6";block_ram_array(167990) := x"7b28";block_ram_array(167992) := x"060c";block_ram_array(167994) := x"3810";block_ram_array(167996) := x"f677";block_ram_array(167998) := x"7ee0";block_ram_array(168000) := x"fcf7";block_ram_array(168002) := x"e730";block_ram_array(168004) := x"0065";block_ram_array(168006) := x"65f0";block_ram_array(168008) := x"0582";block_ram_array(168010) := x"03f0";block_ram_array(168012) := x"fc84";block_ram_array(168014) := x"4a08";block_ram_array(168016) := x"fb5f";block_ram_array(168018) := x"fa78";block_ram_array(168020) := x"fb37";block_ram_array(168022) := x"6ac0";block_ram_array(168024) := x"ff7d";block_ram_array(168026) := x"e6cc";block_ram_array(168028) := x"01dc";block_ram_array(168030) := x"9b58";block_ram_array(168032) := x"ffaa";block_ram_array(168034) := x"a650";block_ram_array(168036) := x"fdaf";block_ram_array(168038) := x"c610";block_ram_array(168040) := x"fe72";block_ram_array(168042) := x"8ab4";block_ram_array(168044) := x"0104";block_ram_array(168046) := x"c630";block_ram_array(168048) := x"0243";block_ram_array(168050) := x"4f6c";block_ram_array(168052) := x"fef4";block_ram_array(168054) := x"30e8";block_ram_array(168056) := x"fd49";block_ram_array(168058) := x"b118";block_ram_array(168060) := x"fbcf";block_ram_array(168062) := x"4740";block_ram_array(168064) := x"fb9b";block_ram_array(168066) := x"dff8";block_ram_array(168068) := x"0257";block_ram_array(168070) := x"fa64";block_ram_array(168072) := x"00f0";block_ram_array(168074) := x"53e0";block_ram_array(168076) := x"0200";block_ram_array(168078) := x"2440";block_ram_array(168080) := x"ff3f";block_ram_array(168082) := x"5e9f";block_ram_array(168084) := x"ffdc";block_ram_array(168086) := x"ae46";block_ram_array(168088) := x"ff95";block_ram_array(168090) := x"4813";block_ram_array(168092) := x"01a8";block_ram_array(168094) := x"2bc4";block_ram_array(168096) := x"00f5";block_ram_array(168098) := x"792a";block_ram_array(168100) := x"00bf";block_ram_array(168102) := x"62aa";block_ram_array(168104) := x"0030";block_ram_array(168106) := x"c158";block_ram_array(168108) := x"fffa";block_ram_array(168110) := x"a8db";block_ram_array(168112) := x"0098";block_ram_array(168114) := x"c2d2";block_ram_array(168116) := x"00a9";block_ram_array(168118) := x"5465";block_ram_array(168120) := x"0099";block_ram_array(168122) := x"e2cb";block_ram_array(168124) := x"ff20";block_ram_array(168126) := x"d5b9";block_ram_array(168128) := x"ff55";block_ram_array(168130) := x"fdd2";block_ram_array(168132) := x"001f";block_ram_array(168134) := x"1fd6";block_ram_array(168136) := x"ffdf";block_ram_array(168138) := x"bcf1";block_ram_array(168140) := x"0049";block_ram_array(168142) := x"4709";block_ram_array(168144) := x"008f";block_ram_array(168146) := x"aec2";block_ram_array(168148) := x"01ec";block_ram_array(168150) := x"dab8";block_ram_array(168152) := x"03a4";block_ram_array(168154) := x"44d0";block_ram_array(168156) := x"fe8f";block_ram_array(168158) := x"ec18";block_ram_array(168160) := x"fe60";block_ram_array(168162) := x"fa9c";block_ram_array(168164) := x"fc85";block_ram_array(168166) := x"32a8";block_ram_array(168168) := 
x"fe2e";block_ram_array(168170) := x"91ca";block_ram_array(168172) := x"007d";block_ram_array(168174) := x"3f03";block_ram_array(168176) := x"ff53";block_ram_array(168178) := x"a064";block_ram_array(168180) := x"0079";block_ram_array(168182) := x"d0d8";block_ram_array(168184) := x"003b";block_ram_array(168186) := x"cc37";block_ram_array(168188) := x"0071";block_ram_array(168190) := x"23a2";block_ram_array(168192) := x"ff57";block_ram_array(168194) := x"ef82";block_ram_array(168196) := x"ffb6";block_ram_array(168198) := x"df4f";block_ram_array(168200) := x"000e";block_ram_array(168202) := x"0ecb";block_ram_array(168204) := x"0115";block_ram_array(168206) := x"7a40";block_ram_array(168208) := x"009d";block_ram_array(168210) := x"0bd8";block_ram_array(168212) := x"ff9d";block_ram_array(168214) := x"7f44";block_ram_array(168216) := x"ffca";block_ram_array(168218) := x"8727";block_ram_array(168220) := x"ffba";block_ram_array(168222) := x"3985";block_ram_array(168224) := x"ff9b";block_ram_array(168226) := x"897b";block_ram_array(168228) := x"ffdb";block_ram_array(168230) := x"3f61";block_ram_array(168232) := x"ffd5";block_ram_array(168234) := x"5330";block_ram_array(168236) := x"004c";block_ram_array(168238) := x"57d0";block_ram_array(168240) := x"ffea";block_ram_array(168242) := x"fc83";block_ram_array(168244) := x"0005";block_ram_array(168246) := x"2144";block_ram_array(168248) := x"0016";block_ram_array(168250) := x"cfd0";block_ram_array(168252) := x"ffe1";block_ram_array(168254) := x"88be";block_ram_array(168256) := x"fef7";block_ram_array(168258) := x"6106";block_ram_array(168260) := x"ffcc";block_ram_array(168262) := x"b416";block_ram_array(168264) := x"000d";block_ram_array(168266) := x"73e9";block_ram_array(168268) := x"0171";block_ram_array(168270) := x"693e";block_ram_array(168272) := x"0095";block_ram_array(168274) := x"30ba";block_ram_array(168276) := x"ff83";block_ram_array(168278) := x"dc0e";block_ram_array(168280) := x"ff81";block_ram_array(168282) := x"15ed";block_ram_array(168284) := x"0086";block_ram_array(168286) := x"344a";block_ram_array(168288) := x"007c";block_ram_array(168290) := x"692c";block_ram_array(168292) := x"ffff";block_ram_array(168294) := x"940f";block_ram_array(168296) := x"ff98";block_ram_array(168298) := x"a0a0";block_ram_array(168300) := x"007a";block_ram_array(168302) := x"0d05";block_ram_array(168304) := x"0101";block_ram_array(168306) := x"3fc6";block_ram_array(168308) := x"003f";block_ram_array(168310) := x"b35e";block_ram_array(168312) := x"ffc4";block_ram_array(168314) := x"8264";block_ram_array(168316) := x"ff67";block_ram_array(168318) := x"99cd";block_ram_array(168320) := x"fff4";block_ram_array(168322) := x"d8dd";block_ram_array(168324) := x"008a";block_ram_array(168326) := x"c924";block_ram_array(168328) := x"0086";block_ram_array(168330) := x"678f";block_ram_array(168332) := x"0005";block_ram_array(168334) := x"52fd";block_ram_array(168336) := x"0037";block_ram_array(168338) := x"af5a";block_ram_array(168340) := x"ffa7";block_ram_array(168342) := x"9b70";block_ram_array(168344) := x"ffde";block_ram_array(168346) := x"16b0";block_ram_array(168348) := x"ffe3";block_ram_array(168350) := x"bf38";block_ram_array(168352) := x"0032";block_ram_array(168354) := x"89e9";block_ram_array(168356) := x"ffea";block_ram_array(168358) := x"c7bb";block_ram_array(168360) := x"ffc8";block_ram_array(168362) := x"59cb";block_ram_array(168364) := x"ffb3";block_ram_array(168366) := x"af06";block_ram_array(168368) := x"ffd8";block_ram_array(168370) := x"bead";block_ram_array(168372) := x"002c";block_ram_array(168374) := x"1276";block_ram_array(168376) := x"0001";block_ram_array(168378) := x"949c";block_ram_array(168380) := x"0008";block_ram_array(168382) := x"06b6";block_ram_array(168384) := x"0009";block_ram_array(168386) := x"3954";block_ram_array(168388) := x"0018";block_ram_array(168390) := x"fcf3";block_ram_array(168392) := x"000e";block_ram_array(168394) := x"e316";block_ram_array(168396) := x"fff3";block_ram_array(168398) := x"b40e";block_ram_array(168400) := x"fffe";block_ram_array(168402) := 
x"435c";block_ram_array(168404) := x"0006";block_ram_array(168406) := x"1db5";block_ram_array(168408) := x"0008";block_ram_array(168410) := x"699c";block_ram_array(168412) := x"fffa";block_ram_array(168414) := x"e5f0";block_ram_array(168416) := x"ffff";block_ram_array(168418) := x"c6f6";block_ram_array(168420) := x"0003";block_ram_array(168422) := x"5dc7";block_ram_array(168424) := x"0006";block_ram_array(168426) := x"e987";block_ram_array(168428) := x"fffc";block_ram_array(168430) := x"7f8e";block_ram_array(168432) := x"ffff";block_ram_array(168434) := x"faf3";block_ram_array(168436) := x"0001";block_ram_array(168438) := x"7ea9";block_ram_array(168440) := x"0006";block_ram_array(168442) := x"1a88";block_ram_array(168444) := x"fffd";block_ram_array(168446) := x"9a19";block_ram_array(168448) := x"0000";block_ram_array(168450) := x"047a";block_ram_array(168452) := x"0000";block_ram_array(168454) := x"07ef";block_ram_array(168456) := x"0005";block_ram_array(168458) := x"60cd";block_ram_array(168460) := x"fffe";block_ram_array(168462) := x"6646";block_ram_array(168464) := x"0000";block_ram_array(168466) := x"0b37";block_ram_array(168468) := x"fffe";block_ram_array(168470) := x"ec83";block_ram_array(168472) := x"0004";block_ram_array(168474) := x"a137";block_ram_array(168476) := x"fffe";block_ram_array(168478) := x"e9a9";block_ram_array(168480) := x"ffff";block_ram_array(168482) := x"f862";block_ram_array(168484) := x"fffe";block_ram_array(168486) := x"39a2";block_ram_array(168488) := x"0004";block_ram_array(168490) := x"1175";block_ram_array(168492) := x"ffff";block_ram_array(168494) := x"5656";block_ram_array(168496) := x"ffff";block_ram_array(168498) := x"ef14";block_ram_array(168500) := x"fffd";block_ram_array(168502) := x"a2ab";block_ram_array(168504) := x"0003";block_ram_array(168506) := x"86f1";block_ram_array(168508) := x"ffff";block_ram_array(168510) := x"9279";block_ram_array(168512) := x"ffff";block_ram_array(168514) := x"bd6f";block_ram_array(168516) := x"fffd";block_ram_array(168518) := x"2758";block_ram_array(168520) := x"0002";block_ram_array(168522) := x"f03e";block_ram_array(168524) := x"ffff";block_ram_array(168526) := x"e90c";block_ram_array(168528) := x"ffff";block_ram_array(168530) := x"ad78";block_ram_array(168532) := x"fffc";block_ram_array(168534) := x"e181";block_ram_array(168536) := x"0002";block_ram_array(168538) := x"7244";block_ram_array(168540) := x"0000";block_ram_array(168542) := x"1ea3";block_ram_array(168544) := x"ffff";block_ram_array(168546) := x"8f95";block_ram_array(168548) := x"fffc";block_ram_array(168550) := x"ad3c";block_ram_array(168552) := x"0001";block_ram_array(168554) := x"f995";block_ram_array(168556) := x"0000";block_ram_array(168558) := x"59c2";block_ram_array(168560) := x"ffff";block_ram_array(168562) := x"82b3";block_ram_array(168564) := x"fffc";block_ram_array(168566) := x"90d8";block_ram_array(168568) := x"0001";block_ram_array(168570) := x"89e5";block_ram_array(168572) := x"0000";block_ram_array(168574) := x"79dc";block_ram_array(168576) := x"ffff";block_ram_array(168578) := x"5afb";block_ram_array(168580) := x"fffc";block_ram_array(168582) := x"9016";block_ram_array(168584) := x"0001";block_ram_array(168586) := x"3cbe";block_ram_array(168588) := x"0000";block_ram_array(168590) := x"b42d";block_ram_array(168592) := x"ffff";block_ram_array(168594) := x"4c19";block_ram_array(168596) := x"fffc";block_ram_array(168598) := x"78fb";block_ram_array(168600) := x"0000";block_ram_array(168602) := x"d4a9";block_ram_array(168604) := x"0000";block_ram_array(168606) := x"de1f";block_ram_array(168608) := x"ffff";block_ram_array(168610) := x"339a";block_ram_array(168612) := x"fffc";block_ram_array(168614) := x"8302";block_ram_array(168616) := x"0000";block_ram_array(168618) := x"729f";block_ram_array(168620) := x"0001";block_ram_array(168622) := x"151b";block_ram_array(168624) := x"ffff";block_ram_array(168626) := x"283f";block_ram_array(168628) := x"fffc";block_ram_array(168630) := x"b087";block_ram_array(168632) := x"0000";block_ram_array(168634) := x"3b1c";block_ram_array(168636) := 
x"0001";block_ram_array(168638) := x"513a";block_ram_array(168640) := x"ffff";block_ram_array(168642) := x"3c2c";block_ram_array(168644) := x"fffc";block_ram_array(168646) := x"cf9c";block_ram_array(168648) := x"0000";block_ram_array(168650) := x"080f";block_ram_array(168652) := x"0001";block_ram_array(168654) := x"5e0e";block_ram_array(168656) := x"ffff";block_ram_array(168658) := x"195c";block_ram_array(168660) := x"fffc";block_ram_array(168662) := x"f1cc";block_ram_array(168664) := x"ffff";block_ram_array(168666) := x"dff6";block_ram_array(168668) := x"0001";block_ram_array(168670) := x"a665";block_ram_array(168672) := x"ffff";block_ram_array(168674) := x"2813";block_ram_array(168676) := x"fffd";block_ram_array(168678) := x"1103";block_ram_array(168680) := x"ffff";block_ram_array(168682) := x"bc63";block_ram_array(168684) := x"0001";block_ram_array(168686) := x"df03";block_ram_array(168688) := x"ffff";block_ram_array(168690) := x"495b";block_ram_array(168692) := x"fffd";block_ram_array(168694) := x"2f95";block_ram_array(168696) := x"ffff";block_ram_array(168698) := x"993e";block_ram_array(168700) := x"0002";block_ram_array(168702) := x"02a6";block_ram_array(168704) := x"ffff";block_ram_array(168706) := x"7194";block_ram_array(168708) := x"fffd";block_ram_array(168710) := x"56ab";block_ram_array(168712) := x"ffff";block_ram_array(168714) := x"8031";block_ram_array(168716) := x"0002";block_ram_array(168718) := x"0286";block_ram_array(168720) := x"ffff";block_ram_array(168722) := x"6867";block_ram_array(168724) := x"fffd";block_ram_array(168726) := x"8527";block_ram_array(168728) := x"ffff";block_ram_array(168730) := x"819e";block_ram_array(168732) := x"0002";block_ram_array(168734) := x"37f6";block_ram_array(168736) := x"ffff";block_ram_array(168738) := x"9117";block_ram_array(168740) := x"fffd";block_ram_array(168742) := x"9a4c";block_ram_array(168744) := x"ffff";block_ram_array(168746) := x"7c0a";block_ram_array(168748) := x"0002";block_ram_array(168750) := x"4e01";block_ram_array(168752) := x"ffff";block_ram_array(168754) := x"b4f6";block_ram_array(168756) := x"fffd";block_ram_array(168758) := x"a23b";block_ram_array(168760) := x"ffff";block_ram_array(168762) := x"560e";block_ram_array(168764) := x"0002";block_ram_array(168766) := x"5a3d";block_ram_array(168768) := x"ffff";block_ram_array(168770) := x"d1a8";block_ram_array(168772) := x"fffd";block_ram_array(168774) := x"dff7";block_ram_array(168776) := x"ffff";block_ram_array(168778) := x"73f3";block_ram_array(168780) := x"0002";block_ram_array(168782) := x"6a09";block_ram_array(168784) := x"ffff";block_ram_array(168786) := x"f855";block_ram_array(168788) := x"fffd";block_ram_array(168790) := x"e095";block_ram_array(168792) := x"ffff";block_ram_array(168794) := x"6ad2";block_ram_array(168796) := x"0002";block_ram_array(168798) := x"6830";block_ram_array(168800) := x"0000";block_ram_array(168802) := x"0e7e";block_ram_array(168804) := x"fffd";block_ram_array(168806) := x"f8f6";block_ram_array(168808) := x"ffff";block_ram_array(168810) := x"7da5";block_ram_array(168812) := x"0002";block_ram_array(168814) := x"6fa6";block_ram_array(168816) := x"0000";block_ram_array(168818) := x"24a9";block_ram_array(168820) := x"fffd";block_ram_array(168822) := x"e587";block_ram_array(168824) := x"ffff";block_ram_array(168826) := x"58ea";block_ram_array(168828) := x"0002";block_ram_array(168830) := x"861b";block_ram_array(168832) := x"0000";block_ram_array(168834) := x"5bcf";block_ram_array(168836) := x"fffe";block_ram_array(168838) := x"0636";block_ram_array(168840) := x"ffff";block_ram_array(168842) := x"5044";block_ram_array(168844) := x"0002";block_ram_array(168846) := x"75ad";block_ram_array(168848) := x"0000";block_ram_array(168850) := x"79cc";block_ram_array(168852) := x"fffe";block_ram_array(168854) := x"34b2";block_ram_array(168856) := x"ffff";block_ram_array(168858) := x"80d0";block_ram_array(168860) := x"0002";block_ram_array(168862) := x"6bb0";block_ram_array(168864) := x"0000";block_ram_array(168866) := x"985e";block_ram_array(168868) := x"fffe";block_ram_array(168870) := 
x"1347";block_ram_array(168872) := x"ffff";block_ram_array(168874) := x"67f7";block_ram_array(168876) := x"0002";block_ram_array(168878) := x"5a8b";block_ram_array(168880) := x"0000";block_ram_array(168882) := x"a6b4";block_ram_array(168884) := x"fffe";block_ram_array(168886) := x"22fe";block_ram_array(168888) := x"ffff";block_ram_array(168890) := x"6682";block_ram_array(168892) := x"0002";block_ram_array(168894) := x"663c";block_ram_array(168896) := x"0000";block_ram_array(168898) := x"e72f";block_ram_array(168900) := x"fffe";block_ram_array(168902) := x"30a4";block_ram_array(168904) := x"ffff";block_ram_array(168906) := x"75d0";block_ram_array(168908) := x"0002";block_ram_array(168910) := x"2c44";block_ram_array(168912) := x"0000";block_ram_array(168914) := x"e44a";block_ram_array(168916) := x"fffe";block_ram_array(168918) := x"1c76";block_ram_array(168920) := x"ffff";block_ram_array(168922) := x"5353";block_ram_array(168924) := x"0002";block_ram_array(168926) := x"1ab9";block_ram_array(168928) := x"0000";block_ram_array(168930) := x"e9ae";block_ram_array(168932) := x"fffe";block_ram_array(168934) := x"4e87";block_ram_array(168936) := x"ffff";block_ram_array(168938) := x"92ce";block_ram_array(168940) := x"0002";block_ram_array(168942) := x"1536";block_ram_array(168944) := x"0001";block_ram_array(168946) := x"03fb";block_ram_array(168948) := x"fffe";block_ram_array(168950) := x"0566";block_ram_array(168952) := x"ffff";block_ram_array(168954) := x"523a";block_ram_array(168956) := x"0001";block_ram_array(168958) := x"f642";block_ram_array(168960) := x"0001";block_ram_array(168962) := x"0400";block_ram_array(168964) := x"fffe";block_ram_array(168966) := x"2600";block_ram_array(168968) := x"ffff";block_ram_array(168970) := x"5677";block_ram_array(168972) := x"0001";block_ram_array(168974) := x"ee4e";block_ram_array(168976) := x"0001";block_ram_array(168978) := x"192d";block_ram_array(168980) := x"fffe";block_ram_array(168982) := x"21d0";block_ram_array(168984) := x"ffff";block_ram_array(168986) := x"47c9";block_ram_array(168988) := x"0001";block_ram_array(168990) := x"cd49";block_ram_array(168992) := x"0001";block_ram_array(168994) := x"0f92";block_ram_array(168996) := x"fffe";block_ram_array(168998) := x"299f";block_ram_array(169000) := x"ffff";block_ram_array(169002) := x"42b3";block_ram_array(169004) := x"0001";block_ram_array(169006) := x"ce31";block_ram_array(169008) := x"0001";block_ram_array(169010) := x"2b16";block_ram_array(169012) := x"fffe";block_ram_array(169014) := x"2a2a";block_ram_array(169016) := x"ffff";block_ram_array(169018) := x"3bf0";block_ram_array(169020) := x"0001";block_ram_array(169022) := x"a34c";block_ram_array(169024) := x"0001";block_ram_array(169026) := x"15e0";block_ram_array(169028) := x"fffe";block_ram_array(169030) := x"22bd";block_ram_array(169032) := x"ffff";block_ram_array(169034) := x"235e";block_ram_array(169036) := x"0001";block_ram_array(169038) := x"a474";block_ram_array(169040) := x"0001";block_ram_array(169042) := x"2004";block_ram_array(169044) := x"fffe";block_ram_array(169046) := x"303a";block_ram_array(169048) := x"ffff";block_ram_array(169050) := x"1bcf";block_ram_array(169052) := x"0001";block_ram_array(169054) := x"92fd";block_ram_array(169056) := x"0001";block_ram_array(169058) := x"213e";block_ram_array(169060) := x"fffe";block_ram_array(169062) := x"3095";block_ram_array(169064) := x"ffff";block_ram_array(169066) := x"04db";block_ram_array(169068) := x"0001";block_ram_array(169070) := x"7ff0";block_ram_array(169072) := x"0001";block_ram_array(169074) := x"154a";block_ram_array(169076) := x"fffe";block_ram_array(169078) := x"4560";block_ram_array(169080) := x"ffff";block_ram_array(169082) := x"0124";block_ram_array(169084) := x"0001";block_ram_array(169086) := x"817d";block_ram_array(169088) := x"0001";block_ram_array(169090) := x"1e3d";block_ram_array(169092) := x"fffe";block_ram_array(169094) := x"53c6";block_ram_array(169096) := x"ffff";block_ram_array(169098) := x"0c66";block_ram_array(169100) := x"0001";block_ram_array(169102) := x"7179";block_ram_array(169104) := 
x"0001";block_ram_array(169106) := x"19ea";block_ram_array(169108) := x"fffe";block_ram_array(169110) := x"3e65";block_ram_array(169112) := x"fffe";block_ram_array(169114) := x"eb42";block_ram_array(169116) := x"0001";block_ram_array(169118) := x"6739";block_ram_array(169120) := x"0001";block_ram_array(169122) := x"0f78";block_ram_array(169124) := x"fffe";block_ram_array(169126) := x"4a91";block_ram_array(169128) := x"fffe";block_ram_array(169130) := x"d187";block_ram_array(169132) := x"0001";block_ram_array(169134) := x"6d6a";block_ram_array(169136) := x"0001";block_ram_array(169138) := x"1737";block_ram_array(169140) := x"fffe";block_ram_array(169142) := x"6935";block_ram_array(169144) := x"fffe";block_ram_array(169146) := x"d59a";block_ram_array(169148) := x"0001";block_ram_array(169150) := x"677f";block_ram_array(169152) := x"0001";block_ram_array(169154) := x"1986";block_ram_array(169156) := x"fffe";block_ram_array(169158) := x"6d6f";block_ram_array(169160) := x"fffe";block_ram_array(169162) := x"c7e0";block_ram_array(169164) := x"0001";block_ram_array(169166) := x"63c1";block_ram_array(169168) := x"0001";block_ram_array(169170) := x"1ac5";block_ram_array(169172) := x"fffe";block_ram_array(169174) := x"7a77";block_ram_array(169176) := x"fffe";block_ram_array(169178) := x"b4fa";block_ram_array(169180) := x"0001";block_ram_array(169182) := x"6902";block_ram_array(169184) := x"0001";block_ram_array(169186) := x"3019";block_ram_array(169188) := x"fffe";block_ram_array(169190) := x"a19e";block_ram_array(169192) := x"fffe";block_ram_array(169194) := x"cedb";block_ram_array(169196) := x"0001";block_ram_array(169198) := x"542a";block_ram_array(169200) := x"0001";block_ram_array(169202) := x"31a6";block_ram_array(169204) := x"fffe";block_ram_array(169206) := x"993e";block_ram_array(169208) := x"fffe";block_ram_array(169210) := x"ca13";block_ram_array(169212) := x"0001";block_ram_array(169214) := x"416b";block_ram_array(169216) := x"0001";block_ram_array(169218) := x"2355";block_ram_array(169220) := x"fffe";block_ram_array(169222) := x"9546";block_ram_array(169224) := x"fffe";block_ram_array(169226) := x"b71c";block_ram_array(169228) := x"0001";block_ram_array(169230) := x"4303";block_ram_array(169232) := x"0001";block_ram_array(169234) := x"1aa3";block_ram_array(169236) := x"fffe";block_ram_array(169238) := x"9d2e";block_ram_array(169240) := x"fffe";block_ram_array(169242) := x"9818";block_ram_array(169244) := x"0001";block_ram_array(169246) := x"58ac";block_ram_array(169248) := x"0001";block_ram_array(169250) := x"3a1d";block_ram_array(169252) := x"fffe";block_ram_array(169254) := x"d05d";block_ram_array(169256) := x"fffe";block_ram_array(169258) := x"b687";block_ram_array(169260) := x"0001";block_ram_array(169262) := x"4527";block_ram_array(169264) := x"0001";block_ram_array(169266) := x"449d";block_ram_array(169268) := x"fffe";block_ram_array(169270) := x"ca71";block_ram_array(169272) := x"fffe";block_ram_array(169274) := x"adf5";block_ram_array(169276) := x"0001";block_ram_array(169278) := x"263d";block_ram_array(169280) := x"0001";block_ram_array(169282) := x"255f";block_ram_array(169284) := x"fffe";block_ram_array(169286) := x"d9a6";block_ram_array(169288) := x"fffe";block_ram_array(169290) := x"ac76";block_ram_array(169292) := x"0001";block_ram_array(169294) := x"41d6";block_ram_array(169296) := x"0001";block_ram_array(169298) := x"421d";block_ram_array(169300) := x"fffe";block_ram_array(169302) := x"f1b0";block_ram_array(169304) := x"fffe";block_ram_array(169306) := x"c43d";block_ram_array(169308) := x"0001";block_ram_array(169310) := x"2662";block_ram_array(169312) := x"0001";block_ram_array(169314) := x"29a0";block_ram_array(169316) := x"fffe";block_ram_array(169318) := x"eb98";block_ram_array(169320) := x"fffe";block_ram_array(169322) := x"cc58";block_ram_array(169324) := x"0001";block_ram_array(169326) := x"3d22";block_ram_array(169328) := x"0001";block_ram_array(169330) := x"2b9e";block_ram_array(169332) := x"fffe";block_ram_array(169334) := x"de04";block_ram_array(169336) := x"fffe";block_ram_array(169338) := 
x"c24f";block_ram_array(169340) := x"0001";block_ram_array(169342) := x"7333";block_ram_array(169344) := x"0001";block_ram_array(169346) := x"9800";block_ram_array(169348) := x"fffe";block_ram_array(169350) := x"d54b";block_ram_array(169352) := x"fffe";block_ram_array(169354) := x"9fce";block_ram_array(169356) := x"0001";block_ram_array(169358) := x"0f32";block_ram_array(169360) := x"0001";block_ram_array(169362) := x"7c93";block_ram_array(169364) := x"fffe";block_ram_array(169366) := x"ffa5";block_ram_array(169368) := x"fffe";block_ram_array(169370) := x"b730";block_ram_array(169372) := x"0000";block_ram_array(169374) := x"e0e5";block_ram_array(169376) := x"0001";block_ram_array(169378) := x"3181";block_ram_array(169380) := x"ffff";block_ram_array(169382) := x"05a6";block_ram_array(169384) := x"fffe";block_ram_array(169386) := x"da04";block_ram_array(169388) := x"0001";block_ram_array(169390) := x"2035";block_ram_array(169392) := x"0001";block_ram_array(169394) := x"440f";block_ram_array(169396) := x"fffe";block_ram_array(169398) := x"c53e";block_ram_array(169400) := x"fffe";block_ram_array(169402) := x"87e0";block_ram_array(169404) := x"0001";block_ram_array(169406) := x"5fe2";block_ram_array(169408) := x"0001";block_ram_array(169410) := x"dada";block_ram_array(169412) := x"ffff";block_ram_array(169414) := x"0942";block_ram_array(169416) := x"fffe";block_ram_array(169418) := x"a844";block_ram_array(169420) := x"0000";block_ram_array(169422) := x"b1ca";block_ram_array(169424) := x"0001";block_ram_array(169426) := x"6a2d";block_ram_array(169428) := x"ffff";block_ram_array(169430) := x"02cf";block_ram_array(169432) := x"fffe";block_ram_array(169434) := x"b013";block_ram_array(169436) := x"0000";block_ram_array(169438) := x"ce74";block_ram_array(169440) := x"0001";block_ram_array(169442) := x"5eb1";block_ram_array(169444) := x"fffe";block_ram_array(169446) := x"e344";block_ram_array(169448) := x"fffe";block_ram_array(169450) := x"7d49";block_ram_array(169452) := x"0000";block_ram_array(169454) := x"d8b9";block_ram_array(169456) := x"0001";block_ram_array(169458) := x"6a59";block_ram_array(169460) := x"fffe";block_ram_array(169462) := x"fca6";block_ram_array(169464) := x"fffe";block_ram_array(169466) := x"5efb";block_ram_array(169468) := x"0000";block_ram_array(169470) := x"b007";block_ram_array(169472) := x"0001";block_ram_array(169474) := x"0b85";block_ram_array(169476) := x"ffff";block_ram_array(169478) := x"23f0";block_ram_array(169480) := x"fffe";block_ram_array(169482) := x"3d13";block_ram_array(169484) := x"0001";block_ram_array(169486) := x"4ae2";block_ram_array(169488) := x"0001";block_ram_array(169490) := x"c137";block_ram_array(169492) := x"ffff";block_ram_array(169494) := x"a01b";block_ram_array(169496) := x"fffe";block_ram_array(169498) := x"d0e6";block_ram_array(169500) := x"0000";block_ram_array(169502) := x"bc26";block_ram_array(169504) := x"0001";block_ram_array(169506) := x"7eea";block_ram_array(169508) := x"ffff";block_ram_array(169510) := x"3c9a";block_ram_array(169512) := x"fffe";block_ram_array(169514) := x"b29e";block_ram_array(169516) := x"0000";block_ram_array(169518) := x"daee";block_ram_array(169520) := x"0001";block_ram_array(169522) := x"c5d3";block_ram_array(169524) := x"ffff";block_ram_array(169526) := x"1fca";block_ram_array(169528) := x"fffe";block_ram_array(169530) := x"652e";block_ram_array(169532) := x"0000";block_ram_array(169534) := x"589f";block_ram_array(169536) := x"0001";block_ram_array(169538) := x"3f92";block_ram_array(169540) := x"ffff";block_ram_array(169542) := x"8cfa";block_ram_array(169544) := x"fffe";block_ram_array(169546) := x"d4e6";block_ram_array(169548) := x"0000";block_ram_array(169550) := x"a64b";block_ram_array(169552) := x"0001";block_ram_array(169554) := x"4d14";block_ram_array(169556) := x"ffff";block_ram_array(169558) := x"30ac";block_ram_array(169560) := x"fffe";block_ram_array(169562) := x"8c63";block_ram_array(169564) := x"0000";block_ram_array(169566) := x"b658";block_ram_array(169568) := x"0001";block_ram_array(169570) := x"54a7";block_ram_array(169572) := 
x"ffff";block_ram_array(169574) := x"6f85";block_ram_array(169576) := x"fffe";block_ram_array(169578) := x"c634";block_ram_array(169580) := x"0000";block_ram_array(169582) := x"cb86";block_ram_array(169584) := x"0001";block_ram_array(169586) := x"85c4";block_ram_array(169588) := x"ffff";block_ram_array(169590) := x"435f";block_ram_array(169592) := x"fffe";block_ram_array(169594) := x"c155";block_ram_array(169596) := x"0000";block_ram_array(169598) := x"8bf4";block_ram_array(169600) := x"0001";block_ram_array(169602) := x"4318";block_ram_array(169604) := x"ffff";block_ram_array(169606) := x"0301";block_ram_array(169608) := x"fffe";block_ram_array(169610) := x"3c0b";block_ram_array(169612) := x"0000";block_ram_array(169614) := x"c797";block_ram_array(169616) := x"0001";block_ram_array(169618) := x"6086";block_ram_array(169620) := x"ffff";block_ram_array(169622) := x"9d7a";block_ram_array(169624) := x"fffe";block_ram_array(169626) := x"accc";block_ram_array(169628) := x"0000";block_ram_array(169630) := x"db0f";block_ram_array(169632) := x"0001";block_ram_array(169634) := x"7fed";block_ram_array(169636) := x"ffff";block_ram_array(169638) := x"7826";block_ram_array(169640) := x"fffe";block_ram_array(169642) := x"d27b";block_ram_array(169644) := x"0001";block_ram_array(169646) := x"0b5c";block_ram_array(169648) := x"0002";block_ram_array(169650) := x"3506";block_ram_array(169652) := x"ffff";block_ram_array(169654) := x"17eb";block_ram_array(169656) := x"fffe";block_ram_array(169658) := x"581e";block_ram_array(169660) := x"0000";block_ram_array(169662) := x"1132";block_ram_array(169664) := x"0001";block_ram_array(169666) := x"7746";block_ram_array(169668) := x"ffff";block_ram_array(169670) := x"7a32";block_ram_array(169672) := x"fffe";block_ram_array(169674) := x"7bc7";block_ram_array(169676) := x"0000";block_ram_array(169678) := x"4936";block_ram_array(169680) := x"0001";block_ram_array(169682) := x"4697";block_ram_array(169684) := x"ffff";block_ram_array(169686) := x"8fd6";block_ram_array(169688) := x"fffe";block_ram_array(169690) := x"a3c9";block_ram_array(169692) := x"0000";block_ram_array(169694) := x"93cf";block_ram_array(169696) := x"0001";block_ram_array(169698) := x"64f9";block_ram_array(169700) := x"ffff";block_ram_array(169702) := x"7d05";block_ram_array(169704) := x"fffe";block_ram_array(169706) := x"c14c";block_ram_array(169708) := x"0000";block_ram_array(169710) := x"c8aa";block_ram_array(169712) := x"0001";block_ram_array(169714) := x"e2ad";block_ram_array(169716) := x"ffff";block_ram_array(169718) := x"258e";block_ram_array(169720) := x"fffe";block_ram_array(169722) := x"4ba4";block_ram_array(169724) := x"0000";block_ram_array(169726) := x"425d";block_ram_array(169728) := x"0001";block_ram_array(169730) := x"9796";block_ram_array(169732) := x"ffff";block_ram_array(169734) := x"79ea";block_ram_array(169736) := x"fffe";block_ram_array(169738) := x"4ee9";block_ram_array(169740) := x"0000";block_ram_array(169742) := x"4a83";block_ram_array(169744) := x"0001";block_ram_array(169746) := x"87fe";block_ram_array(169748) := x"ffff";block_ram_array(169750) := x"bcc0";block_ram_array(169752) := x"fffe";block_ram_array(169754) := x"ad82";block_ram_array(169756) := x"0000";block_ram_array(169758) := x"570d";block_ram_array(169760) := x"0001";block_ram_array(169762) := x"a1cb";block_ram_array(169764) := x"ffff";block_ram_array(169766) := x"5718";block_ram_array(169768) := x"fffe";block_ram_array(169770) := x"400a";block_ram_array(169772) := x"0000";block_ram_array(169774) := x"194d";block_ram_array(169776) := x"0001";block_ram_array(169778) := x"3e49";block_ram_array(169780) := x"ffff";block_ram_array(169782) := x"bff0";block_ram_array(169784) := x"fffe";block_ram_array(169786) := x"8b16";block_ram_array(169788) := x"0000";block_ram_array(169790) := x"9bb7";block_ram_array(169792) := x"0001";block_ram_array(169794) := x"d6d6";block_ram_array(169796) := x"ffff";block_ram_array(169798) := x"9c2a";block_ram_array(169800) := x"fffe";block_ram_array(169802) := x"86a5";block_ram_array(169804) := x"0000";block_ram_array(169806) := 
x"0563";block_ram_array(169808) := x"0001";block_ram_array(169810) := x"62f1";block_ram_array(169812) := x"ffff";block_ram_array(169814) := x"8875";block_ram_array(169816) := x"fffe";block_ram_array(169818) := x"6423";block_ram_array(169820) := x"0000";block_ram_array(169822) := x"4d1a";block_ram_array(169824) := x"0001";block_ram_array(169826) := x"9040";block_ram_array(169828) := x"ffff";block_ram_array(169830) := x"aae2";block_ram_array(169832) := x"fffe";block_ram_array(169834) := x"8d73";block_ram_array(169836) := x"0000";block_ram_array(169838) := x"25d0";block_ram_array(169840) := x"0001";block_ram_array(169842) := x"6269";block_ram_array(169844) := x"ffff";block_ram_array(169846) := x"5261";block_ram_array(169848) := x"fffd";block_ram_array(169850) := x"f09e";block_ram_array(169852) := x"0000";block_ram_array(169854) := x"6635";block_ram_array(169856) := x"0001";block_ram_array(169858) := x"b708";block_ram_array(169860) := x"0000";block_ram_array(169862) := x"049c";block_ram_array(169864) := x"fffe";block_ram_array(169866) := x"723a";block_ram_array(169868) := x"0000";block_ram_array(169870) := x"1400";block_ram_array(169872) := x"0001";block_ram_array(169874) := x"7fcc";block_ram_array(169876) := x"ffff";block_ram_array(169878) := x"bbbb";block_ram_array(169880) := x"fffe";block_ram_array(169882) := x"2e01";block_ram_array(169884) := x"0000";block_ram_array(169886) := x"35b4";block_ram_array(169888) := x"0001";block_ram_array(169890) := x"9d1f";block_ram_array(169892) := x"0000";block_ram_array(169894) := x"1972";block_ram_array(169896) := x"fffe";block_ram_array(169898) := x"86e7";block_ram_array(169900) := x"0000";block_ram_array(169902) := x"2862";block_ram_array(169904) := x"0001";block_ram_array(169906) := x"b638";block_ram_array(169908) := x"ffff";block_ram_array(169910) := x"f250";block_ram_array(169912) := x"fffe";block_ram_array(169914) := x"9f30";block_ram_array(169916) := x"0000";block_ram_array(169918) := x"00fe";block_ram_array(169920) := x"0001";block_ram_array(169922) := x"c0e2";block_ram_array(169924) := x"ffff";block_ram_array(169926) := x"a8ee";block_ram_array(169928) := x"fffe";block_ram_array(169930) := x"415c";block_ram_array(169932) := x"ffff";block_ram_array(169934) := x"a9a0";block_ram_array(169936) := x"0001";block_ram_array(169938) := x"4a00";block_ram_array(169940) := x"ffff";block_ram_array(169942) := x"f318";block_ram_array(169944) := x"fffe";block_ram_array(169946) := x"5bec";block_ram_array(169948) := x"0000";block_ram_array(169950) := x"0af0";block_ram_array(169952) := x"0001";block_ram_array(169954) := x"9891";block_ram_array(169956) := x"ffff";block_ram_array(169958) := x"f7f4";block_ram_array(169960) := x"fffe";block_ram_array(169962) := x"5300";block_ram_array(169964) := x"ffff";block_ram_array(169966) := x"adfd";block_ram_array(169968) := x"0001";block_ram_array(169970) := x"30d6";block_ram_array(169972) := x"0000";block_ram_array(169974) := x"236c";block_ram_array(169976) := x"fffe";block_ram_array(169978) := x"8aa0";block_ram_array(169980) := x"ffff";block_ram_array(169982) := x"f29f";block_ram_array(169984) := x"0001";block_ram_array(169986) := x"3600";block_ram_array(169988) := x"0000";block_ram_array(169990) := x"0000";block_ram_array(169992) := x"fffe";block_ram_array(169994) := x"8aa0";block_ram_array(169996) := x"0000";block_ram_array(169998) := x"0d61";block_ram_array(170000) := x"0001";block_ram_array(170002) := x"30d6";block_ram_array(170004) := x"ffff";block_ram_array(170006) := x"dc94";block_ram_array(170008) := x"fffe";block_ram_array(170010) := x"5300";block_ram_array(170012) := x"0000";block_ram_array(170014) := x"5203";block_ram_array(170016) := x"0001";block_ram_array(170018) := x"9891";block_ram_array(170020) := x"0000";block_ram_array(170022) := x"080c";block_ram_array(170024) := x"fffe";block_ram_array(170026) := x"5bec";block_ram_array(170028) := x"ffff";block_ram_array(170030) := x"f510";block_ram_array(170032) := x"0001";block_ram_array(170034) := x"4a00";block_ram_array(170036) := x"0000";block_ram_array(170038) := x"0ce8";block_ram_array(170040) := 
x"fffe";block_ram_array(170042) := x"415c";block_ram_array(170044) := x"0000";block_ram_array(170046) := x"5660";block_ram_array(170048) := x"0001";block_ram_array(170050) := x"c0e2";block_ram_array(170052) := x"0000";block_ram_array(170054) := x"5712";block_ram_array(170056) := x"fffe";block_ram_array(170058) := x"9f30";block_ram_array(170060) := x"ffff";block_ram_array(170062) := x"ff02";block_ram_array(170064) := x"0001";block_ram_array(170066) := x"b638";block_ram_array(170068) := x"0000";block_ram_array(170070) := x"0db0";block_ram_array(170072) := x"fffe";block_ram_array(170074) := x"86e7";block_ram_array(170076) := x"ffff";block_ram_array(170078) := x"d79e";block_ram_array(170080) := x"0001";block_ram_array(170082) := x"9d1f";block_ram_array(170084) := x"ffff";block_ram_array(170086) := x"e68e";block_ram_array(170088) := x"fffe";block_ram_array(170090) := x"2e01";block_ram_array(170092) := x"ffff";block_ram_array(170094) := x"ca4c";block_ram_array(170096) := x"0001";block_ram_array(170098) := x"7fcc";block_ram_array(170100) := x"0000";block_ram_array(170102) := x"4445";block_ram_array(170104) := x"fffe";block_ram_array(170106) := x"723a";block_ram_array(170108) := x"ffff";block_ram_array(170110) := x"ec00";block_ram_array(170112) := x"0001";block_ram_array(170114) := x"b708";block_ram_array(170116) := x"ffff";block_ram_array(170118) := x"fb64";block_ram_array(170120) := x"fffd";block_ram_array(170122) := x"f09e";block_ram_array(170124) := x"ffff";block_ram_array(170126) := x"99cb";block_ram_array(170128) := x"0001";block_ram_array(170130) := x"6269";block_ram_array(170132) := x"0000";block_ram_array(170134) := x"ad9f";block_ram_array(170136) := x"fffe";block_ram_array(170138) := x"8d73";block_ram_array(170140) := x"ffff";block_ram_array(170142) := x"da30";block_ram_array(170144) := x"0001";block_ram_array(170146) := x"9040";block_ram_array(170148) := x"0000";block_ram_array(170150) := x"551e";block_ram_array(170152) := x"fffe";block_ram_array(170154) := x"6423";block_ram_array(170156) := x"ffff";block_ram_array(170158) := x"b2e6";block_ram_array(170160) := x"0001";block_ram_array(170162) := x"62f1";block_ram_array(170164) := x"0000";block_ram_array(170166) := x"778b";block_ram_array(170168) := x"fffe";block_ram_array(170170) := x"86a5";block_ram_array(170172) := x"ffff";block_ram_array(170174) := x"fa9d";block_ram_array(170176) := x"0001";block_ram_array(170178) := x"d6d6";block_ram_array(170180) := x"0000";block_ram_array(170182) := x"63d6";block_ram_array(170184) := x"fffe";block_ram_array(170186) := x"8b16";block_ram_array(170188) := x"ffff";block_ram_array(170190) := x"6449";block_ram_array(170192) := x"0001";block_ram_array(170194) := x"3e49";block_ram_array(170196) := x"0000";block_ram_array(170198) := x"4010";block_ram_array(170200) := x"fffe";block_ram_array(170202) := x"400a";block_ram_array(170204) := x"ffff";block_ram_array(170206) := x"e6b3";block_ram_array(170208) := x"0001";block_ram_array(170210) := x"a1cb";block_ram_array(170212) := x"0000";block_ram_array(170214) := x"a8e8";block_ram_array(170216) := x"fffe";block_ram_array(170218) := x"ad82";block_ram_array(170220) := x"ffff";block_ram_array(170222) := x"a8f3";block_ram_array(170224) := x"0001";block_ram_array(170226) := x"87fe";block_ram_array(170228) := x"0000";block_ram_array(170230) := x"4340";block_ram_array(170232) := x"fffe";block_ram_array(170234) := x"4ee9";block_ram_array(170236) := x"ffff";block_ram_array(170238) := x"b57d";block_ram_array(170240) := x"0001";block_ram_array(170242) := x"9796";block_ram_array(170244) := x"0000";block_ram_array(170246) := x"8616";block_ram_array(170248) := x"fffe";block_ram_array(170250) := x"4ba4";block_ram_array(170252) := x"ffff";block_ram_array(170254) := x"bda3";block_ram_array(170256) := x"0001";block_ram_array(170258) := x"e2ad";block_ram_array(170260) := x"0000";block_ram_array(170262) := x"da72";block_ram_array(170264) := x"fffe";block_ram_array(170266) := x"c14c";block_ram_array(170268) := x"ffff";block_ram_array(170270) := x"3756";block_ram_array(170272) := x"0001";block_ram_array(170274) := 
x"64f9";block_ram_array(170276) := x"0000";block_ram_array(170278) := x"82fb";block_ram_array(170280) := x"fffe";block_ram_array(170282) := x"a3c9";block_ram_array(170284) := x"ffff";block_ram_array(170286) := x"6c31";block_ram_array(170288) := x"0001";block_ram_array(170290) := x"4697";block_ram_array(170292) := x"0000";block_ram_array(170294) := x"702a";block_ram_array(170296) := x"fffe";block_ram_array(170298) := x"7bc7";block_ram_array(170300) := x"ffff";block_ram_array(170302) := x"b6ca";block_ram_array(170304) := x"0001";block_ram_array(170306) := x"7746";block_ram_array(170308) := x"0000";block_ram_array(170310) := x"85ce";block_ram_array(170312) := x"fffe";block_ram_array(170314) := x"581e";block_ram_array(170316) := x"ffff";block_ram_array(170318) := x"eece";block_ram_array(170320) := x"0002";block_ram_array(170322) := x"3506";block_ram_array(170324) := x"0000";block_ram_array(170326) := x"e815";block_ram_array(170328) := x"fffe";block_ram_array(170330) := x"d27b";block_ram_array(170332) := x"fffe";block_ram_array(170334) := x"f4a4";block_ram_array(170336) := x"0001";block_ram_array(170338) := x"7fed";block_ram_array(170340) := x"0000";block_ram_array(170342) := x"87da";block_ram_array(170344) := x"fffe";block_ram_array(170346) := x"accc";block_ram_array(170348) := x"ffff";block_ram_array(170350) := x"24f1";block_ram_array(170352) := x"0001";block_ram_array(170354) := x"6086";block_ram_array(170356) := x"0000";block_ram_array(170358) := x"6286";block_ram_array(170360) := x"fffe";block_ram_array(170362) := x"3c0b";block_ram_array(170364) := x"ffff";block_ram_array(170366) := x"3869";block_ram_array(170368) := x"0001";block_ram_array(170370) := x"4318";block_ram_array(170372) := x"0000";block_ram_array(170374) := x"fcff";block_ram_array(170376) := x"fffe";block_ram_array(170378) := x"c155";block_ram_array(170380) := x"ffff";block_ram_array(170382) := x"740c";block_ram_array(170384) := x"0001";block_ram_array(170386) := x"85c4";block_ram_array(170388) := x"0000";block_ram_array(170390) := x"bca1";block_ram_array(170392) := x"fffe";block_ram_array(170394) := x"c634";block_ram_array(170396) := x"ffff";block_ram_array(170398) := x"347a";block_ram_array(170400) := x"0001";block_ram_array(170402) := x"54a7";block_ram_array(170404) := x"0000";block_ram_array(170406) := x"907b";block_ram_array(170408) := x"fffe";block_ram_array(170410) := x"8c63";block_ram_array(170412) := x"ffff";block_ram_array(170414) := x"49a8";block_ram_array(170416) := x"0001";block_ram_array(170418) := x"4d14";block_ram_array(170420) := x"0000";block_ram_array(170422) := x"cf54";block_ram_array(170424) := x"fffe";block_ram_array(170426) := x"d4e6";block_ram_array(170428) := x"ffff";block_ram_array(170430) := x"59b5";block_ram_array(170432) := x"0001";block_ram_array(170434) := x"3f92";block_ram_array(170436) := x"0000";block_ram_array(170438) := x"7306";block_ram_array(170440) := x"fffe";block_ram_array(170442) := x"652e";block_ram_array(170444) := x"ffff";block_ram_array(170446) := x"a761";block_ram_array(170448) := x"0001";block_ram_array(170450) := x"c5d3";block_ram_array(170452) := x"0000";block_ram_array(170454) := x"e036";block_ram_array(170456) := x"fffe";block_ram_array(170458) := x"b29e";block_ram_array(170460) := x"ffff";block_ram_array(170462) := x"2512";block_ram_array(170464) := x"0001";block_ram_array(170466) := x"7eea";block_ram_array(170468) := x"0000";block_ram_array(170470) := x"c366";block_ram_array(170472) := x"fffe";block_ram_array(170474) := x"d0e6";block_ram_array(170476) := x"ffff";block_ram_array(170478) := x"43da";block_ram_array(170480) := x"0001";block_ram_array(170482) := x"c137";block_ram_array(170484) := x"0000";block_ram_array(170486) := x"5fe5";block_ram_array(170488) := x"fffe";block_ram_array(170490) := x"3d13";block_ram_array(170492) := x"fffe";block_ram_array(170494) := x"b51e";block_ram_array(170496) := x"0001";block_ram_array(170498) := x"0b85";block_ram_array(170500) := x"0000";block_ram_array(170502) := x"dc10";block_ram_array(170504) := x"fffe";block_ram_array(170506) := x"5efb";block_ram_array(170508) := 
x"ffff";block_ram_array(170510) := x"4ff9";block_ram_array(170512) := x"0001";block_ram_array(170514) := x"6a59";block_ram_array(170516) := x"0001";block_ram_array(170518) := x"035a";block_ram_array(170520) := x"fffe";block_ram_array(170522) := x"7d49";block_ram_array(170524) := x"ffff";block_ram_array(170526) := x"2747";block_ram_array(170528) := x"0001";block_ram_array(170530) := x"5eb1";block_ram_array(170532) := x"0001";block_ram_array(170534) := x"1cbc";block_ram_array(170536) := x"fffe";block_ram_array(170538) := x"b013";block_ram_array(170540) := x"ffff";block_ram_array(170542) := x"318c";block_ram_array(170544) := x"0001";block_ram_array(170546) := x"6a2d";block_ram_array(170548) := x"0000";block_ram_array(170550) := x"fd31";block_ram_array(170552) := x"fffe";block_ram_array(170554) := x"a844";block_ram_array(170556) := x"ffff";block_ram_array(170558) := x"4e36";block_ram_array(170560) := x"0001";block_ram_array(170562) := x"dada";block_ram_array(170564) := x"0000";block_ram_array(170566) := x"f6be";block_ram_array(170568) := x"fffe";block_ram_array(170570) := x"87e0";block_ram_array(170572) := x"fffe";block_ram_array(170574) := x"a01e";block_ram_array(170576) := x"0001";block_ram_array(170578) := x"440f";block_ram_array(170580) := x"0001";block_ram_array(170582) := x"3ac2";block_ram_array(170584) := x"fffe";block_ram_array(170586) := x"da04";block_ram_array(170588) := x"fffe";block_ram_array(170590) := x"dfcb";block_ram_array(170592) := x"0001";block_ram_array(170594) := x"3181";block_ram_array(170596) := x"0000";block_ram_array(170598) := x"fa5a";block_ram_array(170600) := x"fffe";block_ram_array(170602) := x"b730";block_ram_array(170604) := x"ffff";block_ram_array(170606) := x"1f1b";block_ram_array(170608) := x"0001";block_ram_array(170610) := x"7c93";block_ram_array(170612) := x"0001";block_ram_array(170614) := x"005b";block_ram_array(170616) := x"fffe";block_ram_array(170618) := x"9fce";block_ram_array(170620) := x"fffe";block_ram_array(170622) := x"f0ce";block_ram_array(170624) := x"0001";block_ram_array(170626) := x"9800";block_ram_array(170628) := x"0001";block_ram_array(170630) := x"2ab5";block_ram_array(170632) := x"fffe";block_ram_array(170634) := x"c24f";block_ram_array(170636) := x"fffe";block_ram_array(170638) := x"8ccd";block_ram_array(170640) := x"0001";block_ram_array(170642) := x"2b9e";block_ram_array(170644) := x"0001";block_ram_array(170646) := x"21fc";block_ram_array(170648) := x"fffe";block_ram_array(170650) := x"cc58";block_ram_array(170652) := x"fffe";block_ram_array(170654) := x"c2de";block_ram_array(170656) := x"0001";block_ram_array(170658) := x"29a0";block_ram_array(170660) := x"0001";block_ram_array(170662) := x"1468";block_ram_array(170664) := x"fffe";block_ram_array(170666) := x"c43d";block_ram_array(170668) := x"fffe";block_ram_array(170670) := x"d99e";block_ram_array(170672) := x"0001";block_ram_array(170674) := x"421d";block_ram_array(170676) := x"0001";block_ram_array(170678) := x"0e50";block_ram_array(170680) := x"fffe";block_ram_array(170682) := x"ac76";block_ram_array(170684) := x"fffe";block_ram_array(170686) := x"be2a";block_ram_array(170688) := x"0001";block_ram_array(170690) := x"255f";block_ram_array(170692) := x"0001";block_ram_array(170694) := x"265a";block_ram_array(170696) := x"fffe";block_ram_array(170698) := x"adf5";block_ram_array(170700) := x"fffe";block_ram_array(170702) := x"d9c3";block_ram_array(170704) := x"0001";block_ram_array(170706) := x"449d";block_ram_array(170708) := x"0001";block_ram_array(170710) := x"358f";block_ram_array(170712) := x"fffe";block_ram_array(170714) := x"b687";block_ram_array(170716) := x"fffe";block_ram_array(170718) := x"bad9";block_ram_array(170720) := x"0001";block_ram_array(170722) := x"3a1d";block_ram_array(170724) := x"0001";block_ram_array(170726) := x"2fa3";block_ram_array(170728) := x"fffe";block_ram_array(170730) := x"9818";block_ram_array(170732) := x"fffe";block_ram_array(170734) := x"a754";block_ram_array(170736) := x"0001";block_ram_array(170738) := x"1aa3";block_ram_array(170740) := x"0001";block_ram_array(170742) := 
x"62d2";block_ram_array(170744) := x"fffe";block_ram_array(170746) := x"b71c";block_ram_array(170748) := x"fffe";block_ram_array(170750) := x"bcfd";block_ram_array(170752) := x"0001";block_ram_array(170754) := x"2355";block_ram_array(170756) := x"0001";block_ram_array(170758) := x"6aba";block_ram_array(170760) := x"fffe";block_ram_array(170762) := x"ca13";block_ram_array(170764) := x"fffe";block_ram_array(170766) := x"be95";block_ram_array(170768) := x"0001";block_ram_array(170770) := x"31a6";block_ram_array(170772) := x"0001";block_ram_array(170774) := x"66c2";block_ram_array(170776) := x"fffe";block_ram_array(170778) := x"cedb";block_ram_array(170780) := x"fffe";block_ram_array(170782) := x"abd6";block_ram_array(170784) := x"0001";block_ram_array(170786) := x"3019";block_ram_array(170788) := x"0001";block_ram_array(170790) := x"5e62";block_ram_array(170792) := x"fffe";block_ram_array(170794) := x"b4fa";block_ram_array(170796) := x"fffe";block_ram_array(170798) := x"96fe";block_ram_array(170800) := x"0001";block_ram_array(170802) := x"1ac5";block_ram_array(170804) := x"0001";block_ram_array(170806) := x"8589";block_ram_array(170808) := x"fffe";block_ram_array(170810) := x"c7e0";block_ram_array(170812) := x"fffe";block_ram_array(170814) := x"9c3f";block_ram_array(170816) := x"0001";block_ram_array(170818) := x"1986";block_ram_array(170820) := x"0001";block_ram_array(170822) := x"9291";block_ram_array(170824) := x"fffe";block_ram_array(170826) := x"d59a";block_ram_array(170828) := x"fffe";block_ram_array(170830) := x"9881";block_ram_array(170832) := x"0001";block_ram_array(170834) := x"1737";block_ram_array(170836) := x"0001";block_ram_array(170838) := x"96cb";block_ram_array(170840) := x"fffe";block_ram_array(170842) := x"d187";block_ram_array(170844) := x"fffe";block_ram_array(170846) := x"9296";block_ram_array(170848) := x"0001";block_ram_array(170850) := x"0f78";block_ram_array(170852) := x"0001";block_ram_array(170854) := x"b56f";block_ram_array(170856) := x"fffe";block_ram_array(170858) := x"eb42";block_ram_array(170860) := x"fffe";block_ram_array(170862) := x"98c7";block_ram_array(170864) := x"0001";block_ram_array(170866) := x"19ea";block_ram_array(170868) := x"0001";block_ram_array(170870) := x"c19b";block_ram_array(170872) := x"ffff";block_ram_array(170874) := x"0c66";block_ram_array(170876) := x"fffe";block_ram_array(170878) := x"8e87";block_ram_array(170880) := x"0001";block_ram_array(170882) := x"1e3d";block_ram_array(170884) := x"0001";block_ram_array(170886) := x"ac3a";block_ram_array(170888) := x"ffff";block_ram_array(170890) := x"0124";block_ram_array(170892) := x"fffe";block_ram_array(170894) := x"7e83";block_ram_array(170896) := x"0001";block_ram_array(170898) := x"154a";block_ram_array(170900) := x"0001";block_ram_array(170902) := x"baa0";block_ram_array(170904) := x"ffff";block_ram_array(170906) := x"04db";block_ram_array(170908) := x"fffe";block_ram_array(170910) := x"8010";block_ram_array(170912) := x"0001";block_ram_array(170914) := x"213e";block_ram_array(170916) := x"0001";block_ram_array(170918) := x"cf6b";block_ram_array(170920) := x"ffff";block_ram_array(170922) := x"1bcf";block_ram_array(170924) := x"fffe";block_ram_array(170926) := x"6d03";block_ram_array(170928) := x"0001";block_ram_array(170930) := x"2004";block_ram_array(170932) := x"0001";block_ram_array(170934) := x"cfc6";block_ram_array(170936) := x"ffff";block_ram_array(170938) := x"235e";block_ram_array(170940) := x"fffe";block_ram_array(170942) := x"5b8c";block_ram_array(170944) := x"0001";block_ram_array(170946) := x"15e0";block_ram_array(170948) := x"0001";block_ram_array(170950) := x"dd43";block_ram_array(170952) := x"ffff";block_ram_array(170954) := x"3bf0";block_ram_array(170956) := x"fffe";block_ram_array(170958) := x"5cb4";block_ram_array(170960) := x"0001";block_ram_array(170962) := x"2b16";block_ram_array(170964) := x"0001";block_ram_array(170966) := x"d5d6";block_ram_array(170968) := x"ffff";block_ram_array(170970) := x"42b3";block_ram_array(170972) := x"fffe";block_ram_array(170974) := x"31cf";block_ram_array(170976) := 
x"0001";block_ram_array(170978) := x"0f92";block_ram_array(170980) := x"0001";block_ram_array(170982) := x"d661";block_ram_array(170984) := x"ffff";block_ram_array(170986) := x"47c9";block_ram_array(170988) := x"fffe";block_ram_array(170990) := x"32b7";block_ram_array(170992) := x"0001";block_ram_array(170994) := x"192d";block_ram_array(170996) := x"0001";block_ram_array(170998) := x"de30";block_ram_array(171000) := x"ffff";block_ram_array(171002) := x"5677";block_ram_array(171004) := x"fffe";block_ram_array(171006) := x"11b2";block_ram_array(171008) := x"0001";block_ram_array(171010) := x"0400";block_ram_array(171012) := x"0001";block_ram_array(171014) := x"da00";block_ram_array(171016) := x"ffff";block_ram_array(171018) := x"523a";block_ram_array(171020) := x"fffe";block_ram_array(171022) := x"09be";block_ram_array(171024) := x"0001";block_ram_array(171026) := x"03fb";block_ram_array(171028) := x"0001";block_ram_array(171030) := x"fa9a";block_ram_array(171032) := x"ffff";block_ram_array(171034) := x"92ce";block_ram_array(171036) := x"fffd";block_ram_array(171038) := x"eaca";block_ram_array(171040) := x"0000";block_ram_array(171042) := x"e9ae";block_ram_array(171044) := x"0001";block_ram_array(171046) := x"b179";block_ram_array(171048) := x"ffff";block_ram_array(171050) := x"5353";block_ram_array(171052) := x"fffd";block_ram_array(171054) := x"e547";block_ram_array(171056) := x"0000";block_ram_array(171058) := x"e44a";block_ram_array(171060) := x"0001";block_ram_array(171062) := x"e38a";block_ram_array(171064) := x"ffff";block_ram_array(171066) := x"75d0";block_ram_array(171068) := x"fffd";block_ram_array(171070) := x"d3bc";block_ram_array(171072) := x"0000";block_ram_array(171074) := x"e72f";block_ram_array(171076) := x"0001";block_ram_array(171078) := x"cf5c";block_ram_array(171080) := x"ffff";block_ram_array(171082) := x"6682";block_ram_array(171084) := x"fffd";block_ram_array(171086) := x"99c4";block_ram_array(171088) := x"0000";block_ram_array(171090) := x"a6b4";block_ram_array(171092) := x"0001";block_ram_array(171094) := x"dd02";block_ram_array(171096) := x"ffff";block_ram_array(171098) := x"67f7";block_ram_array(171100) := x"fffd";block_ram_array(171102) := x"a575";block_ram_array(171104) := x"0000";block_ram_array(171106) := x"985e";block_ram_array(171108) := x"0001";block_ram_array(171110) := x"ecb9";block_ram_array(171112) := x"ffff";block_ram_array(171114) := x"80d0";block_ram_array(171116) := x"fffd";block_ram_array(171118) := x"9450";block_ram_array(171120) := x"0000";block_ram_array(171122) := x"79cc";block_ram_array(171124) := x"0001";block_ram_array(171126) := x"cb4e";block_ram_array(171128) := x"ffff";block_ram_array(171130) := x"5044";block_ram_array(171132) := x"fffd";block_ram_array(171134) := x"8a53";block_ram_array(171136) := x"0000";block_ram_array(171138) := x"5bcf";block_ram_array(171140) := x"0001";block_ram_array(171142) := x"f9ca";block_ram_array(171144) := x"ffff";block_ram_array(171146) := x"58ea";block_ram_array(171148) := x"fffd";block_ram_array(171150) := x"79e5";block_ram_array(171152) := x"0000";block_ram_array(171154) := x"24a9";block_ram_array(171156) := x"0002";block_ram_array(171158) := x"1a79";block_ram_array(171160) := x"ffff";block_ram_array(171162) := x"7da5";block_ram_array(171164) := x"fffd";block_ram_array(171166) := x"905a";block_ram_array(171168) := x"0000";block_ram_array(171170) := x"0e7e";block_ram_array(171172) := x"0002";block_ram_array(171174) := x"070a";block_ram_array(171176) := x"ffff";block_ram_array(171178) := x"6ad2";block_ram_array(171180) := x"fffd";block_ram_array(171182) := x"97d0";block_ram_array(171184) := x"ffff";block_ram_array(171186) := x"f855";block_ram_array(171188) := x"0002";block_ram_array(171190) := x"1f6b";block_ram_array(171192) := x"ffff";block_ram_array(171194) := x"73f3";block_ram_array(171196) := x"fffd";block_ram_array(171198) := x"95f7";block_ram_array(171200) := x"ffff";block_ram_array(171202) := x"d1a8";block_ram_array(171204) := x"0002";block_ram_array(171206) := x"2009";block_ram_array(171208) := x"ffff";block_ram_array(171210) := 
x"560e";block_ram_array(171212) := x"fffd";block_ram_array(171214) := x"a5c3";block_ram_array(171216) := x"ffff";block_ram_array(171218) := x"b4f6";block_ram_array(171220) := x"0002";block_ram_array(171222) := x"5dc5";block_ram_array(171224) := x"ffff";block_ram_array(171226) := x"7c0a";block_ram_array(171228) := x"fffd";block_ram_array(171230) := x"b1ff";block_ram_array(171232) := x"ffff";block_ram_array(171234) := x"9117";block_ram_array(171236) := x"0002";block_ram_array(171238) := x"65b4";block_ram_array(171240) := x"ffff";block_ram_array(171242) := x"819e";block_ram_array(171244) := x"fffd";block_ram_array(171246) := x"c80a";block_ram_array(171248) := x"ffff";block_ram_array(171250) := x"6867";block_ram_array(171252) := x"0002";block_ram_array(171254) := x"7ad9";block_ram_array(171256) := x"ffff";block_ram_array(171258) := x"8031";block_ram_array(171260) := x"fffd";block_ram_array(171262) := x"fd7a";block_ram_array(171264) := x"ffff";block_ram_array(171266) := x"7194";block_ram_array(171268) := x"0002";block_ram_array(171270) := x"a955";block_ram_array(171272) := x"ffff";block_ram_array(171274) := x"993e";block_ram_array(171276) := x"fffd";block_ram_array(171278) := x"fd5a";block_ram_array(171280) := x"ffff";block_ram_array(171282) := x"495b";block_ram_array(171284) := x"0002";block_ram_array(171286) := x"d06b";block_ram_array(171288) := x"ffff";block_ram_array(171290) := x"bc63";block_ram_array(171292) := x"fffe";block_ram_array(171294) := x"20fd";block_ram_array(171296) := x"ffff";block_ram_array(171298) := x"2813";block_ram_array(171300) := x"0002";block_ram_array(171302) := x"eefd";block_ram_array(171304) := x"ffff";block_ram_array(171306) := x"dff6";block_ram_array(171308) := x"fffe";block_ram_array(171310) := x"599b";block_ram_array(171312) := x"ffff";block_ram_array(171314) := x"195c";block_ram_array(171316) := x"0003";block_ram_array(171318) := x"0e34";block_ram_array(171320) := x"0000";block_ram_array(171322) := x"080f";block_ram_array(171324) := x"fffe";block_ram_array(171326) := x"a1f2";block_ram_array(171328) := x"ffff";block_ram_array(171330) := x"3c2c";block_ram_array(171332) := x"0003";block_ram_array(171334) := x"3064";block_ram_array(171336) := x"0000";block_ram_array(171338) := x"3b1c";block_ram_array(171340) := x"fffe";block_ram_array(171342) := x"aec6";block_ram_array(171344) := x"ffff";block_ram_array(171346) := x"283f";block_ram_array(171348) := x"0003";block_ram_array(171350) := x"4f79";block_ram_array(171352) := x"0000";block_ram_array(171354) := x"729f";block_ram_array(171356) := x"fffe";block_ram_array(171358) := x"eae5";block_ram_array(171360) := x"ffff";block_ram_array(171362) := x"339a";block_ram_array(171364) := x"0003";block_ram_array(171366) := x"7cfe";block_ram_array(171368) := x"0000";block_ram_array(171370) := x"d4a9";block_ram_array(171372) := x"ffff";block_ram_array(171374) := x"21e1";block_ram_array(171376) := x"ffff";block_ram_array(171378) := x"4c19";block_ram_array(171380) := x"0003";block_ram_array(171382) := x"8705";block_ram_array(171384) := x"0001";block_ram_array(171386) := x"3cbe";block_ram_array(171388) := x"ffff";block_ram_array(171390) := x"4bd3";block_ram_array(171392) := x"ffff";block_ram_array(171394) := x"5afb";block_ram_array(171396) := x"0003";block_ram_array(171398) := x"6fea";block_ram_array(171400) := x"0001";block_ram_array(171402) := x"89e5";block_ram_array(171404) := x"ffff";block_ram_array(171406) := x"8624";block_ram_array(171408) := x"ffff";block_ram_array(171410) := x"82b3";block_ram_array(171412) := x"0003";block_ram_array(171414) := x"6f28";block_ram_array(171416) := x"0001";block_ram_array(171418) := x"f995";block_ram_array(171420) := x"ffff";block_ram_array(171422) := x"a63e";block_ram_array(171424) := x"ffff";block_ram_array(171426) := x"8f95";block_ram_array(171428) := x"0003";block_ram_array(171430) := x"52c4";block_ram_array(171432) := x"0002";block_ram_array(171434) := x"7244";block_ram_array(171436) := x"ffff";block_ram_array(171438) := x"e15d";block_ram_array(171440) := x"ffff";block_ram_array(171442) := x"ad78";block_ram_array(171444) := 
x"0003";block_ram_array(171446) := x"1e7f";block_ram_array(171448) := x"0002";block_ram_array(171450) := x"f03e";block_ram_array(171452) := x"0000";block_ram_array(171454) := x"16f4";block_ram_array(171456) := x"ffff";block_ram_array(171458) := x"bd6f";block_ram_array(171460) := x"0002";block_ram_array(171462) := x"d8a8";block_ram_array(171464) := x"0003";block_ram_array(171466) := x"86f1";block_ram_array(171468) := x"0000";block_ram_array(171470) := x"6d87";block_ram_array(171472) := x"ffff";block_ram_array(171474) := x"ef14";block_ram_array(171476) := x"0002";block_ram_array(171478) := x"5d55";block_ram_array(171480) := x"0004";block_ram_array(171482) := x"1175";block_ram_array(171484) := x"0000";block_ram_array(171486) := x"a9aa";block_ram_array(171488) := x"ffff";block_ram_array(171490) := x"f862";block_ram_array(171492) := x"0001";block_ram_array(171494) := x"c65e";block_ram_array(171496) := x"0004";block_ram_array(171498) := x"a137";block_ram_array(171500) := x"0001";block_ram_array(171502) := x"1657";block_ram_array(171504) := x"0000";block_ram_array(171506) := x"0b37";block_ram_array(171508) := x"0001";block_ram_array(171510) := x"137d";block_ram_array(171512) := x"0005";block_ram_array(171514) := x"60cd";block_ram_array(171516) := x"0001";block_ram_array(171518) := x"99ba";block_ram_array(171520) := x"0000";block_ram_array(171522) := x"047a";block_ram_array(171524) := x"ffff";block_ram_array(171526) := x"f811";block_ram_array(171528) := x"0006";block_ram_array(171530) := x"1a88";block_ram_array(171532) := x"0002";block_ram_array(171534) := x"65e7";block_ram_array(171536) := x"ffff";block_ram_array(171538) := x"faf3";block_ram_array(171540) := x"fffe";block_ram_array(171542) := x"8157";block_ram_array(171544) := x"0006";block_ram_array(171546) := x"e987";block_ram_array(171548) := x"0003";block_ram_array(171550) := x"8072";block_ram_array(171552) := x"ffff";block_ram_array(171554) := x"c6f6";block_ram_array(171556) := x"fffc";block_ram_array(171558) := x"a239";block_ram_array(171560) := x"0008";block_ram_array(171562) := x"699c";block_ram_array(171564) := x"0005";block_ram_array(171566) := x"1a10";block_ram_array(171568) := x"fffe";block_ram_array(171570) := x"435c";block_ram_array(171572) := x"fff9";block_ram_array(171574) := x"e24b";block_ram_array(171576) := x"000e";block_ram_array(171578) := x"e316";block_ram_array(171580) := x"000c";block_ram_array(171582) := x"4bf2";block_ram_array(171584) := x"0009";block_ram_array(171586) := x"3954";block_ram_array(171588) := x"ffe7";block_ram_array(171590) := x"030d";block_ram_array(171592) := x"0001";block_ram_array(171594) := x"949c";block_ram_array(171596) := x"fff7";block_ram_array(171598) := x"f94a";block_ram_array(171600) := x"ffd8";block_ram_array(171602) := x"bead";block_ram_array(171604) := x"ffd3";block_ram_array(171606) := x"ed8a";block_ram_array(171608) := x"ffc8";block_ram_array(171610) := x"59cb";block_ram_array(171612) := x"004c";block_ram_array(171614) := x"50fa";block_ram_array(171616) := x"0032";block_ram_array(171618) := x"89e9";block_ram_array(171620) := x"0015";block_ram_array(171622) := x"3845";block_ram_array(171624) := x"ffde";block_ram_array(171626) := x"16b0";block_ram_array(171628) := x"001c";block_ram_array(171630) := x"40c8";block_ram_array(171632) := x"0037";block_ram_array(171634) := x"af5a";block_ram_array(171636) := x"0058";block_ram_array(171638) := x"6490";block_ram_array(171640) := x"0086";block_ram_array(171642) := x"678f";block_ram_array(171644) := x"fffa";block_ram_array(171646) := x"ad03";block_ram_array(171648) := x"fff4";block_ram_array(171650) := x"d8dd";block_ram_array(171652) := x"ff75";block_ram_array(171654) := x"36dc";block_ram_array(171656) := x"ffc4";block_ram_array(171658) := x"8264";block_ram_array(171660) := x"0098";block_ram_array(171662) := x"6633";block_ram_array(171664) := x"0101";block_ram_array(171666) := x"3fc6";block_ram_array(171668) := x"ffc0";block_ram_array(171670) := x"4ca2";block_ram_array(171672) := x"ff98";block_ram_array(171674) := x"a0a0";block_ram_array(171676) := x"ff85";block_ram_array(171678) := 
x"f2fb";block_ram_array(171680) := x"007c";block_ram_array(171682) := x"692c";block_ram_array(171684) := x"0000";block_ram_array(171686) := x"6bf1";block_ram_array(171688) := x"ff81";block_ram_array(171690) := x"15ed";block_ram_array(171692) := x"ff79";block_ram_array(171694) := x"cbb6";block_ram_array(171696) := x"0095";block_ram_array(171698) := x"30ba";block_ram_array(171700) := x"007c";block_ram_array(171702) := x"23f2";block_ram_array(171704) := x"000d";block_ram_array(171706) := x"73e9";block_ram_array(171708) := x"fe8e";block_ram_array(171710) := x"96c2";block_ram_array(171712) := x"fef7";block_ram_array(171714) := x"6106";block_ram_array(171716) := x"0033";block_ram_array(171718) := x"4bea";block_ram_array(171720) := x"0016";block_ram_array(171722) := x"cfd0";block_ram_array(171724) := x"001e";block_ram_array(171726) := x"7742";block_ram_array(171728) := x"ffea";block_ram_array(171730) := x"fc83";block_ram_array(171732) := x"fffa";block_ram_array(171734) := x"debc";block_ram_array(171736) := x"ffd5";block_ram_array(171738) := x"5330";block_ram_array(171740) := x"ffb3";block_ram_array(171742) := x"a830";block_ram_array(171744) := x"ff9b";block_ram_array(171746) := x"897b";block_ram_array(171748) := x"0024";block_ram_array(171750) := x"c09f";block_ram_array(171752) := x"ffca";block_ram_array(171754) := x"8727";block_ram_array(171756) := x"0045";block_ram_array(171758) := x"c67b";block_ram_array(171760) := x"009d";block_ram_array(171762) := x"0bd8";block_ram_array(171764) := x"0062";block_ram_array(171766) := x"80bc";block_ram_array(171768) := x"000e";block_ram_array(171770) := x"0ecb";block_ram_array(171772) := x"feea";block_ram_array(171774) := x"85c0";block_ram_array(171776) := x"ff57";block_ram_array(171778) := x"ef82";block_ram_array(171780) := x"0049";block_ram_array(171782) := x"20b1";block_ram_array(171784) := x"003b";block_ram_array(171786) := x"cc37";block_ram_array(171788) := x"ff8e";block_ram_array(171790) := x"dc5e";block_ram_array(171792) := x"ff53";block_ram_array(171794) := x"a064";block_ram_array(171796) := x"ff86";block_ram_array(171798) := x"2f28";block_ram_array(171800) := x"fe2e";block_ram_array(171802) := x"91ca";block_ram_array(171804) := x"ff82";block_ram_array(171806) := x"c0fd";block_ram_array(171808) := x"fe60";block_ram_array(171810) := x"fa9c";block_ram_array(171812) := x"037a";block_ram_array(171814) := x"cd58";block_ram_array(171816) := x"03a4";block_ram_array(171818) := x"44d0";block_ram_array(171820) := x"0170";block_ram_array(171822) := x"13e8";block_ram_array(171824) := x"008f";block_ram_array(171826) := x"aec2";block_ram_array(171828) := x"fe13";block_ram_array(171830) := x"2548";block_ram_array(171832) := x"ffdf";block_ram_array(171834) := x"bcf1";block_ram_array(171836) := x"ffb6";block_ram_array(171838) := x"b8f7";block_ram_array(171840) := x"ff55";block_ram_array(171842) := x"fdd2";block_ram_array(171844) := x"ffe0";block_ram_array(171846) := x"e02a";block_ram_array(171848) := x"0099";block_ram_array(171850) := x"e2cb";block_ram_array(171852) := x"00df";block_ram_array(171854) := x"2a47";block_ram_array(171856) := x"0098";block_ram_array(171858) := x"c2d2";block_ram_array(171860) := x"ff56";block_ram_array(171862) := x"ab9b";block_ram_array(171864) := x"0030";block_ram_array(171866) := x"c158";block_ram_array(171868) := x"0005";block_ram_array(171870) := x"5725";block_ram_array(171872) := x"00f5";block_ram_array(171874) := x"792a";block_ram_array(171876) := x"ff40";block_ram_array(171878) := x"9d56";block_ram_array(171880) := x"ff95";block_ram_array(171882) := x"4813";block_ram_array(171884) := x"fe57";block_ram_array(171886) := x"d43c";block_ram_array(171888) := x"ff3f";block_ram_array(171890) := x"5e9f";block_ram_array(171892) := x"0023";block_ram_array(171894) := x"51ba";block_ram_array(171896) := x"00f0";block_ram_array(171898) := x"53e0";block_ram_array(171900) := x"fdff";block_ram_array(171902) := x"dbc0";block_ram_array(171904) := x"fb9b";block_ram_array(171906) := x"dff8";block_ram_array(171908) := x"fda8";block_ram_array(171910) := x"059c";block_ram_array(171912) := 
x"fd49";block_ram_array(171914) := x"b118";block_ram_array(171916) := x"0430";block_ram_array(171918) := x"b8c0";block_ram_array(171920) := x"0243";block_ram_array(171922) := x"4f6c";block_ram_array(171924) := x"010b";block_ram_array(171926) := x"cf18";block_ram_array(171928) := x"fe72";block_ram_array(171930) := x"8ab4";block_ram_array(171932) := x"fefb";block_ram_array(171934) := x"39d0";block_ram_array(171936) := x"ffaa";block_ram_array(171938) := x"a650";block_ram_array(171940) := x"0250";block_ram_array(171942) := x"39f0";block_ram_array(171944) := x"ff7d";block_ram_array(171946) := x"e6cc";block_ram_array(171948) := x"fe23";block_ram_array(171950) := x"64a8";block_ram_array(171952) := x"fb5f";block_ram_array(171954) := x"fa78";block_ram_array(171956) := x"04c8";block_ram_array(171958) := x"9540";block_ram_array(171960) := x"0582";block_ram_array(171962) := x"03f0";block_ram_array(171964) := x"037b";block_ram_array(171966) := x"b5f8";block_ram_array(171968) := x"fcf7";block_ram_array(171970) := x"e730";block_ram_array(171972) := x"ff9a";block_ram_array(171974) := x"9a10";block_ram_array(171976) := x"060c";block_ram_array(171978) := x"3810";block_ram_array(171980) := x"0988";block_ram_array(171982) := x"8120";block_ram_array(171984) := x"09d6";block_ram_array(171986) := x"e790";block_ram_array(171988) := x"f959";block_ram_array(171990) := x"84d8";block_ram_array(171992) := x"ff81";block_ram_array(171994) := x"d320";block_ram_array(171996) := x"fb1e";block_ram_array(171998) := x"6350";block_ram_array(172000) := x"ff39";block_ram_array(172002) := x"189b";block_ram_array(172004) := x"fafc";block_ram_array(172006) := x"02c0";block_ram_array(172008) := x"fcd6";block_ram_array(172010) := x"f228";block_ram_array(172012) := x"003a";block_ram_array(172014) := x"2839";block_ram_array(172016) := x"0046";block_ram_array(172018) := x"45b1";block_ram_array(172020) := x"fcd7";block_ram_array(172022) := x"e664";block_ram_array(172024) := x"fadf";block_ram_array(172026) := x"4dd0";block_ram_array(172028) := x"015a";block_ram_array(172030) := x"5cf0";
        --------------------
        --=0
        --------------------
-- 			      a_h(0)                        a_h(0)			  b_h(0)		        b_l(0)			      a_h(1)			     a_l(1)			    b_h(1)		    	   b_l(1)
        block_ram_array(0) := x"024d";block_ram_array(2) := x"7000";block_ram_array(4) := x"0000";block_ram_array(6) := x"0000";block_ram_array(8) := x"feb9";block_ram_array(10) := x"a290";block_ram_array(12) := x"fe79";block_ram_array(14) := x"a730";block_ram_array(16) := x"ffc7";block_ram_array(18) := x"7700";block_ram_array(20) := x"0120";block_ram_array(22) := x"8e58";block_ram_array(24) := x"0011";block_ram_array(26) := x"6d93";block_ram_array(28) := x"0000";block_ram_array(30) := x"f559";block_ram_array(32) := x"00e7";block_ram_array(34) := x"072d";block_ram_array(36) := x"0054";block_ram_array(38) := x"1984";block_ram_array(40) := x"ff90";block_ram_array(42) := x"690e";block_ram_array(44) := x"fe68";block_ram_array(46) := x"8f5c";block_ram_array(48) := x"fec1";block_ram_array(50) := x"4c08";block_ram_array(52) := x"0173";block_ram_array(54) := x"27e0";block_ram_array(56) := x"01c2";block_ram_array(58) := x"83be";block_ram_array(60) := x"0043";block_ram_array(62) := x"09ab";block_ram_array(64) := x"ff7e";block_ram_array(66) := x"6a30";block_ram_array(68) := x"fec1";block_ram_array(70) := x"9caa";block_ram_array(72) := x"ff91";block_ram_array(74) := x"9cb9";block_ram_array(76) := x"0083";block_ram_array(78) := x"7bab";block_ram_array(80) := x"ffd2";block_ram_array(82) := x"da51";block_ram_array(84) := x"001b";block_ram_array(86) := x"7afa";block_ram_array(88) := x"00bb";block_ram_array(90) := x"8d8c";block_ram_array(92) := x"00c2";block_ram_array(94) := x"7d1c";block_ram_array(96) := x"004b";block_ram_array(98) := x"cc6d";block_ram_array(100) := x"fe4b";block_ram_array(102) := x"1e10";block_ram_array(104) := x"fe45";block_ram_array(106) := x"c672";block_ram_array(108) := x"00ff";block_ram_array(110) := x"25c7";block_ram_array(112) := x"01a4";block_ram_array(114) := x"c740";block_ram_array(116) := x"007f";block_ram_array(118) := x"e8c4";block_ram_array(120) := x"ff70";block_ram_array(122) := x"95f2";block_ram_array(124) := x"ff31";block_ram_array(126) := x"b3b8";block_ram_array(128) := x"0061";block_ram_array(130) := x"9f7d";block_ram_array(132) := x"0022";block_ram_array(134) := x"3027";block_ram_array(136) := x"fee5";block_ram_array(138) := x"cf48";block_ram_array(140) := x"ffb7";block_ram_array(142) := x"7d9c";block_ram_array(144) := x"00f6";block_ram_array(146) := x"882b";block_ram_array(148) := x"0168";block_ram_array(150) := x"90a4";block_ram_array(152) := x"0062";block_ram_array(154) := x"7dde";block_ram_array(156) := x"fe42";block_ram_array(158) := x"2520";block_ram_array(160) := x"fec8";block_ram_array(162) := x"a102";block_ram_array(164) := x"00ae";block_ram_array(166) := x"5bf4";block_ram_array(168) := x"00af";block_ram_array(170) := x"c38a";block_ram_array(172) := x"0032";block_ram_array(174) := x"fc49";block_ram_array(176) := x"ffd5";block_ram_array(178) := x"9613";block_ram_array(180) := x"0019";block_ram_array(182) := x"27ab";block_ram_array(184) := x"00b7";block_ram_array(186) := x"83ee";block_ram_array(188) := x"ffa4";block_ram_array(190) := x"aa6d";block_ram_array(192) := x"fece";block_ram_array(194) := x"acb0";block_ram_array(196) := x"ff71";block_ram_array(198) := x"55e4";block_ram_array(200) := x"004f";block_ram_array(202) := x"78de";block_ram_array(204) := x"018d";block_ram_array(206) := x"b5a4";block_ram_array(208) := x"00fa";block_ram_array(210) := x"9408";block_ram_array(212) := x"fed9";block_ram_array(214) := x"5658";block_ram_array(216) := x"fef4";block_ram_array(218) := x"93c0";block_ram_array(220) := x"0011";block_ram_array(222) := x"c4a3";block_ram_array(224) := x"005d";block_ram_array(226) := x"ac98";block_ram_array(228) := x"0002";block_ram_array(230) := x"d084";block_ram_array(232) := x"ff5f";block_ram_array(234) := x"250c";block_ram_array(236) := x"009a";block_ram_array(238) := x"da42";block_ram_array(240) := x"01a7";block_ram_array(242) := x"ef18";block_ram_array(244) := x"ffd2";block_ram_array(246) := x"6eab";block_ram_array(248) := x"fe68";block_ram_array(250) := x"73be";block_ram_array(252) := x"feb4";block_ram_array(254) := x"28a0";block_ram_array(256) := x"0024";block_ram_
array(258) := x"2147";block_ram_array(260) := x"01dd";block_ram_array(262) := x"2950";block_ram_array(264) := x"00c2";block_ram_array(266) := x"98c4";block_ram_array(268) := x"ff1e";block_ram_array(270) := x"fed0";block_ram_array(272) := x"ffd7";block_ram_array(274) := x"7ba9";block_ram_array(276) := x"0025";block_ram_array(278) := x"47eb";block_ram_array(280) := x"ffb2";block_ram_array(282) := x"e761";block_ram_array(284) := x"ff28";block_ram_array(286) := x"f6b0";block_ram_array(288) := x"ff3e";block_ram_array(290) := x"c046";block_ram_array(292) := x"016f";block_ram_array(294) := x"26fa";block_ram_array(296) := x"01e9";block_ram_array(298) := x"7c84";block_ram_array(300) := x"ffb2";block_ram_array(302) := x"65a6";block_ram_array(304) := x"fec2";block_ram_array(306) := x"0d58";block_ram_array(308) := x"fea6";block_ram_array(310) := x"db44";block_ram_array(312) := x"ff99";block_ram_array(314) := x"c7a9";block_ram_array(316) := x"0154";block_ram_array(318) := x"d274";block_ram_array(320) := x"00b1";block_ram_array(322) := x"7f9a";block_ram_array(324) := x"ffea";block_ram_array(326) := x"7bdb";block_ram_array(328) := x"004c";block_ram_array(330) := x"f538";block_ram_array(332) := x"ffee";block_ram_array(334) := x"fc5a";block_ram_array(336) := x"ffb7";block_ram_array(338) := x"8166";block_ram_array(340) := x"fede";block_ram_array(342) := x"78ec";block_ram_array(344) := x"feb0";block_ram_array(346) := x"66b0";block_ram_array(348) := x"0162";block_ram_array(350) := x"fe1e";block_ram_array(352) := x"023a";block_ram_array(354) := x"6fb8";block_ram_array(356) := x"0041";block_ram_array(358) := x"26be";block_ram_array(360) := x"feec";block_ram_array(362) := x"a1f0";block_ram_array(364) := x"fe4e";block_ram_array(366) := x"089a";block_ram_array(368) := x"ffa5";block_ram_array(370) := x"0b97";block_ram_array(372) := x"012a";block_ram_array(374) := x"4ec8";block_ram_array(376) := x"000e";block_ram_array(378) := x"723b";block_ram_array(380) := x"ffec";block_ram_array(382) := x"3a4f";block_ram_array(384) := x"00e9";block_ram_array(386) := x"0dd6";block_ram_array(388) := x"0091";block_ram_array(390) := x"198e";block_ram_array(392) := x"ffb2";block_ram_array(394) := x"4dd4";block_ram_array(396) := x"fe1f";block_ram_array(398) := x"89ca";block_ram_array(400) := x"fe8c";block_ram_array(402) := x"2d76";block_ram_array(404) := x"01a4";block_ram_array(406) := x"9e4c";block_ram_array(408) := x"01ea";block_ram_array(410) := x"0f1a";block_ram_array(412) := x"0021";block_ram_array(414) := x"6967";block_ram_array(416) := x"ff61";block_ram_array(418) := x"864e";block_ram_array(420) := x"fef1";block_ram_array(422) := x"c3b0";block_ram_array(424) := x"ffc0";block_ram_array(426) := x"f7e2";block_ram_array(428) := x"0043";block_ram_array(430) := x"f2d7";block_ram_array(432) := x"ff89";block_ram_array(434) := x"8667";block_ram_array(436) := x"0050";block_ram_array(438) := x"8648";block_ram_array(440) := x"010c";block_ram_array(442) := x"f616";block_ram_array(444) := x"00a7";block_ram_array(446) := x"7bef";block_ram_array(448) := x"0004";block_ram_array(450) := x"f92f";block_ram_array(452) := x"fe53";block_ram_array(454) := x"52a6";block_ram_array(456) := x"fe81";block_ram_array(458) := x"2ac2";block_ram_array(460) := x"00fc";block_ram_array(462) := x"1030";block_ram_array(464) := x"016f";block_ram_array(466) := x"3b20";block_ram_array(468) := x"0081";block_ram_array(470) := x"9daa";block_ram_array(472) := x"ffa4";block_ram_array(474) := x"a316";block_ram_array(476) := x"ff33";block_ram_array(478) := x"2c21";block_ram_array(480) := x"0031";block_ram_array(482) := x"83a4";block_ram_array(484) := x"0015";block_ram_array(486) := x"ff8e";block_ram_array(488) := x"ff04";block_ram_array(490) := x"1d6d";block_ram_array(492) := x"ffce";block_ram_array(494) := x"6e9c";block_ram_array(496) := x"00f4";block_ram_array(498) := x"dc30";block_ram_array(500) := x"0158";block_ram_array(502) := x"af86";block_ram_array(504) := x"0055";block_ram_array(506) := x"222c";block_ram_array(508) := x"fe31";block_ram_array(510) := x"ca88";block_ram_array(512) := x"fec3";block_ram_
array(514) := x"af74";block_ram_array(516) := x"00dc";block_ram_array(518) := x"9aae";block_ram_array(520) := x"00cf";block_ram_array(522) := x"3d6b";block_ram_array(524) := x"0007";block_ram_array(526) := x"191b";block_ram_array(528) := x"ffb8";block_ram_array(530) := x"bcba";block_ram_array(532) := x"0036";block_ram_array(534) := x"1b16";block_ram_array(536) := x"00c3";block_ram_array(538) := x"1b14";block_ram_array(540) := x"ff76";block_ram_array(542) := x"3867";block_ram_array(544) := x"feab";block_ram_array(546) := x"cb96";block_ram_array(548) := x"ffc8";block_ram_array(550) := x"cdd4";block_ram_array(552) := x"00b3";block_ram_array(554) := x"653b";block_ram_array(556) := x"0138";block_ram_array(558) := x"2bec";block_ram_array(560) := x"0076";block_ram_array(562) := x"1659";block_ram_array(564) := x"fef0";block_ram_array(566) := x"7e60";block_ram_array(568) := x"ff54";block_ram_array(570) := x"9c60";block_ram_array(572) := x"002a";block_ram_array(574) := x"7b4f";block_ram_array(576) := x"0021";block_ram_array(578) := x"0f4d";block_ram_array(580) := x"fffe";block_ram_array(582) := x"2ae7";block_ram_array(584) := x"ffbc";block_ram_array(586) := x"950d";block_ram_array(588) := x"0087";block_ram_array(590) := x"4b79";block_ram_array(592) := x"011f";block_ram_array(594) := x"1312";block_ram_array(596) := x"ffb0";block_ram_array(598) := x"bf13";block_ram_array(600) := x"fec3";block_ram_array(602) := x"cee8";block_ram_array(604) := x"ff28";block_ram_array(606) := x"9401";block_ram_array(608) := x"0030";block_ram_array(610) := x"f991";block_ram_array(612) := x"016e";block_ram_array(614) := x"b030";block_ram_array(616) := x"0095";block_ram_array(618) := x"9044";block_ram_array(620) := x"ff33";block_ram_array(622) := x"997e";block_ram_array(624) := x"ffc5";block_ram_array(626) := x"9404";block_ram_array(628) := x"0038";block_ram_array(630) := x"da8b";block_ram_array(632) := x"ffe0";block_ram_array(634) := x"71f4";block_ram_array(636) := x"ff4f";block_ram_array(638) := x"62ac";block_ram_array(640) := x"ff60";block_ram_array(642) := x"7c13";block_ram_array(644) := x"012b";block_ram_array(646) := x"4612";block_ram_array(648) := x"0187";block_ram_array(650) := x"a9d0";block_ram_array(652) := x"ff96";block_ram_array(654) := x"9cab";block_ram_array(656) := x"fed7";block_ram_array(658) := x"8734";block_ram_array(660) := x"ff31";block_ram_array(662) := x"760a";block_ram_array(664) := x"0007";block_ram_array(666) := x"78a9";block_ram_array(668) := x"00e5";block_ram_array(670) := x"86e6";block_ram_array(672) := x"0037";block_ram_array(674) := x"1c79";block_ram_array(676) := x"ffe8";block_ram_array(678) := x"f33d";block_ram_array(680) := x"0070";block_ram_array(682) := x"a745";block_ram_array(684) := x"0000";block_ram_array(686) := x"aa7d";block_ram_array(688) := x"ff95";block_ram_array(690) := x"ac8a";block_ram_array(692) := x"ff28";block_ram_array(694) := x"7d73";block_ram_array(696) := x"ff4e";block_ram_array(698) := x"f55f";block_ram_array(700) := x"010a";block_ram_array(702) := x"54a2";block_ram_array(704) := x"0157";block_ram_array(706) := x"b4c8";block_ram_array(708) := x"000d";block_ram_array(710) := x"b590";block_ram_array(712) := x"ff65";block_ram_array(714) := x"4aea";block_ram_array(716) := x"fefc";block_ram_array(718) := x"b018";block_ram_array(720) := x"ffb2";block_ram_array(722) := x"8fff";block_ram_array(724) := x"00ab";block_ram_array(726) := x"3fbd";block_ram_array(728) := x"0011";block_ram_array(730) := x"c175";block_ram_array(732) := x"0000";block_ram_array(734) := x"9d6a";block_ram_array(736) := x"008b";block_ram_array(738) := x"89f2";block_ram_array(740) := x"0061";block_ram_array(742) := x"3633";block_ram_array(744) := x"ffe9";block_ram_array(746) := x"0994";block_ram_array(748) := x"fec2";block_ram_array(750) := x"566e";block_ram_array(752) := x"feef";block_ram_array(754) := x"838a";block_ram_array(756) := x"010a";block_ram_array(758) := x"1e78";block_ram_array(760) := x"014f";block_ram_array(762) := x"e446";block_ram_array(764) := x"001d";block_ram_array(766) := x"aed6";block_ram_array(768) := x"ff88";block_ram_
array(770) := x"47fe";block_ram_array(772) := x"ff5a";block_ram_array(774) := x"ff08";block_ram_array(776) := x"fffe";block_ram_array(778) := x"c929";block_ram_array(780) := x"001b";block_ram_array(782) := x"42ed";block_ram_array(784) := x"ff7d";block_ram_array(786) := x"58aa";block_ram_array(788) := x"002f";block_ram_array(790) := x"9756";block_ram_array(792) := x"00d4";block_ram_array(794) := x"5d8e";block_ram_array(796) := x"0082";block_ram_array(798) := x"f4c5";block_ram_array(800) := x"ffee";block_ram_array(802) := x"394c";block_ram_array(804) := x"fee0";block_ram_array(806) := x"6d44";block_ram_array(808) := x"ff2a";block_ram_array(810) := x"d7d7";block_ram_array(812) := x"009a";block_ram_array(814) := x"b4ae";block_ram_array(816) := x"00b2";block_ram_array(818) := x"55d4";block_ram_array(820) := x"004f";block_ram_array(822) := x"6540";block_ram_array(824) := x"fffa";block_ram_array(826) := x"9c1a";block_ram_array(828) := x"ff9d";block_ram_array(830) := x"1d6f";block_ram_array(832) := x"0003";block_ram_array(834) := x"f2b8";block_ram_array(836) := x"ffea";block_ram_array(838) := x"0290";block_ram_array(840) := x"ff75";block_ram_array(842) := x"d53c";block_ram_array(844) := x"fff0";block_ram_array(846) := x"eda6";block_ram_array(848) := x"0071";block_ram_array(850) := x"d039";block_ram_array(852) := x"00cd";block_ram_array(854) := x"659d";block_ram_array(856) := x"0065";block_ram_array(858) := x"0c59";block_ram_array(860) := x"ff01";block_ram_array(862) := x"0a70";block_ram_array(864) := x"ff21";block_ram_array(866) := x"4eee";block_ram_array(868) := x"0057";block_ram_array(870) := x"9bab";block_ram_array(872) := x"0086";block_ram_array(874) := x"35db";block_ram_array(876) := x"0028";block_ram_array(878) := x"71f6";block_ram_array(880) := x"ffc8";block_ram_array(882) := x"05d4";block_ram_array(884) := x"000d";block_ram_array(886) := x"4e8e";block_ram_array(888) := x"008d";block_ram_array(890) := x"e737";block_ram_array(892) := x"ffc6";block_ram_array(894) := x"b92f";block_ram_array(896) := x"ff26";block_ram_array(898) := x"fb4c";block_ram_array(900) := x"ffb7";block_ram_array(902) := x"e1bb";block_ram_array(904) := x"0064";block_ram_array(906) := x"0cd9";block_ram_array(908) := x"00d6";block_ram_array(910) := x"19f0";block_ram_array(912) := x"0048";block_ram_array(914) := x"6e18";block_ram_array(916) := x"ff5a";block_ram_array(918) := x"6920";block_ram_array(920) := x"ffac";block_ram_array(922) := x"1c35";block_ram_array(924) := x"001c";block_ram_array(926) := x"3a54";block_ram_array(928) := x"0001";block_ram_array(930) := x"e521";block_ram_array(932) := x"ffee";block_ram_array(934) := x"4a66";block_ram_array(936) := x"ffdd";block_ram_array(938) := x"1038";block_ram_array(940) := x"0059";block_ram_array(942) := x"15a8";block_ram_array(944) := x"0097";block_ram_array(946) := x"669c";block_ram_array(948) := x"ffdd";block_ram_array(950) := x"3e3c";block_ram_array(952) := x"ff78";block_ram_array(954) := x"9c5a";block_ram_array(956) := x"ff7d";block_ram_array(958) := x"ee45";block_ram_array(960) := x"ffe6";block_ram_array(962) := x"1dd7";block_ram_array(964) := x"00b5";block_ram_array(966) := x"bb25";block_ram_array(968) := x"0070";block_ram_array(970) := x"49eb";block_ram_array(972) := x"ffb7";block_ram_array(974) := x"244e";block_ram_array(976) := x"ffd0";block_ram_array(978) := x"031a";block_ram_array(980) := x"0008";block_ram_array(982) := x"fd45";block_ram_array(984) := x"0017";block_ram_array(986) := x"0ff9";block_ram_array(988) := x"ffad";block_ram_array(990) := x"6837";block_ram_array(992) := x"ff71";block_ram_array(994) := x"646e";block_ram_array(996) := x"006f";block_ram_array(998) := x"deb5";block_ram_array(1000) := x"00e5";block_ram_array(1002) := x"24cf";block_ram_array(1004) := x"001c";block_ram_array(1006) := x"e32f";block_ram_array(1008) := x"ff81";block_ram_array(1010) := x"7023";block_ram_array(1012) := x"ff52";block_ram_array(1014) := x"b413";block_ram_array(1016) := x"ffe9";block_ram_array(1018) := x"1cdc";block_ram_array(1020) := x"0087";block_ram_array(1022) := x"c9c0";block_ram_array(1024) := x"
0010";block_ram_array(1026) := x"3900";block_ram_array(1028) := x"ffe5";block_ram_array(1030) := x"6100";block_ram_array(1032) := x"0041";block_ram_array(1034) := x"54c7";block_ram_array(1036) := x"0036";block_ram_array(1038) := x"b894";block_ram_array(1040) := x"fff8";block_ram_array(1042) := x"07ff";block_ram_array(1044) := x"ff5f";block_ram_array(1046) := x"67b3";block_ram_array(1048) := x"ff69";block_ram_array(1050) := x"e8d5";block_ram_array(1052) := x"0077";block_ram_array(1054) := x"497d";block_ram_array(1056) := x"00aa";block_ram_array(1058) := x"e122";block_ram_array(1060) := x"003d";block_ram_array(1062) := x"8a9d";block_ram_array(1064) := x"ffea";block_ram_array(1066) := x"7bca";block_ram_array(1068) := x"ff73";block_ram_array(1070) := x"d363";block_ram_array(1072) := x"ffbc";block_ram_array(1074) := x"bcfd";block_ram_array(1076) := x"002b";block_ram_array(1078) := x"3725";block_ram_array(1080) := x"fff7";block_ram_array(1082) := x"974c";block_ram_array(1084) := x"0012";block_ram_array(1086) := x"735d";block_ram_array(1088) := x"0038";block_ram_array(1090) := x"23ce";block_ram_array(1092) := x"0050";block_ram_array(1094) := x"102f";block_ram_array(1096) := x"0045";block_ram_array(1098) := x"ed0b";block_ram_array(1100) := x"ff5f";block_ram_array(1102) := x"afc7";block_ram_array(1104) := x"ff30";block_ram_array(1106) := x"4d88";block_ram_array(1108) := x"0031";block_ram_array(1110) := x"453d";block_ram_array(1112) := x"009b";block_ram_array(1114) := x"9840";block_ram_array(1116) := x"0076";block_ram_array(1118) := x"59b6";block_ram_array(1120) := x"fff5";block_ram_array(1122) := x"e0b9";block_ram_array(1124) := x"ff86";block_ram_array(1126) := x"28c2";block_ram_array(1128) := x"fffc";block_ram_array(1130) := x"d3d6";block_ram_array(1132) := x"0012";block_ram_array(1134) := x"4249";block_ram_array(1136) := x"ffa5";block_ram_array(1138) := x"acec";block_ram_array(1140) := x"ffe2";block_ram_array(1142) := x"5952";block_ram_array(1144) := x"0046";block_ram_array(1146) := x"fa20";block_ram_array(1148) := x"009b";block_ram_array(1150) := x"6b68";block_ram_array(1152) := x"0057";block_ram_array(1154) := x"3c0f";block_ram_array(1156) := x"ff50";block_ram_array(1158) := x"ea78";block_ram_array(1160) := x"ff59";block_ram_array(1162) := x"2825";block_ram_array(1164) := x"001c";block_ram_array(1166) := x"bbc5";block_ram_array(1168) := x"0047";block_ram_array(1170) := x"d13b";block_ram_array(1172) := x"0050";block_ram_array(1174) := x"d7cc";block_ram_array(1176) := x"0014";block_ram_array(1178) := x"ae99";block_ram_array(1180) := x"ffe2";block_ram_array(1182) := x"51c7";block_ram_array(1184) := x"001c";block_ram_array(1186) := x"c09c";block_ram_array(1188) := x"ffdf";block_ram_array(1190) := x"424d";block_ram_array(1192) := x"ffa3";block_ram_array(1194) := x"6a9a";block_ram_array(1196) := x"ffd5";block_ram_array(1198) := x"de7e";block_ram_array(1200) := x"000a";block_ram_array(1202) := x"6b53";block_ram_array(1204) := x"0090";block_ram_array(1206) := x"20ff";block_ram_array(1208) := x"0080";block_ram_array(1210) := x"3d40";block_ram_array(1212) := x"ff9e";block_ram_array(1214) := x"ded3";block_ram_array(1216) := x"ff78";block_ram_array(1218) := x"89bc";block_ram_array(1220) := x"ffd9";block_ram_array(1222) := x"dca8";block_ram_array(1224) := x"0027";block_ram_array(1226) := x"8b29";block_ram_array(1228) := x"0049";block_ram_array(1230) := x"78df";block_ram_array(1232) := x"ffed";block_ram_array(1234) := x"2141";block_ram_array(1236) := x"fff5";block_ram_array(1238) := x"bc37";block_ram_array(1240) := x"0059";block_ram_array(1242) := x"88cb";block_ram_array(1244) := x"0010";block_ram_array(1246) := x"0d58";block_ram_array(1248) := x"ffa6";block_ram_array(1250) := x"ed57";block_ram_array(1252) := x"ff87";block_ram_array(1254) := x"a139";block_ram_array(1256) := x"ffe2";block_ram_array(1258) := x"91b4";block_ram_array(1260) := x"00a2";block_ram_array(1262) := x"9b79";block_ram_array(1264) := x"0070";block_ram_array(1266) := x"6a66";block_ram_array(1268) := x"ffb6";block_ram_array(1270) := x"a85e";block_ram_array(1272) := x"
ffba";block_ram_array(1274) := x"3dc5";block_ram_array(1276) := x"fff5";block_ram_array(1278) := x"b401";block_ram_array(1280) := x"0011";block_ram_array(1282) := x"fd6f";block_ram_array(1284) := x"fff2";block_ram_array(1286) := x"58b2";block_ram_array(1288) := x"ffc1";block_ram_array(1290) := x"18da";block_ram_array(1292) := x"002c";block_ram_array(1294) := x"8d3b";block_ram_array(1296) := x"0070";block_ram_array(1298) := x"769f";block_ram_array(1300) := x"001b";block_ram_array(1302) := x"1de7";block_ram_array(1304) := x"ffd0";block_ram_array(1306) := x"b24d";block_ram_array(1308) := x"ff8b";block_ram_array(1310) := x"1a3a";block_ram_array(1312) := x"ffc1";block_ram_array(1314) := x"e472";block_ram_array(1316) := x"005b";block_ram_array(1318) := x"d094";block_ram_array(1320) := x"0049";block_ram_array(1322) := x"c5a5";block_ram_array(1324) := x"fffe";block_ram_array(1326) := x"24ca";block_ram_array(1328) := x"ffee";block_ram_array(1330) := x"5f52";block_ram_array(1332) := x"fff4";block_ram_array(1334) := x"c79b";block_ram_array(1336) := x"001e";block_ram_array(1338) := x"96fa";block_ram_array(1340) := x"ffdb";block_ram_array(1342) := x"959a";block_ram_array(1344) := x"ff96";block_ram_array(1346) := x"7196";block_ram_array(1348) := x"0008";block_ram_array(1350) := x"8ef4";block_ram_array(1352) := x"0064";block_ram_array(1354) := x"6be1";block_ram_array(1356) := x"0063";block_ram_array(1358) := x"129d";block_ram_array(1360) := x"0007";block_ram_array(1362) := x"8e80";block_ram_array(1364) := x"ff75";block_ram_array(1366) := x"61bd";block_ram_array(1368) := x"ffb7";block_ram_array(1370) := x"1c26";block_ram_array(1372) := x"0040";block_ram_array(1374) := x"8a7e";block_ram_array(1376) := x"001e";block_ram_array(1378) := x"7242";block_ram_array(1380) := x"fff4";block_ram_array(1382) := x"469c";block_ram_array(1384) := x"fffc";block_ram_array(1386) := x"91b4";block_ram_array(1388) := x"0039";block_ram_array(1390) := x"940e";block_ram_array(1392) := x"004e";block_ram_array(1394) := x"5d43";block_ram_array(1396) := x"ffaa";block_ram_array(1398) := x"0922";block_ram_array(1400) := x"ff70";block_ram_array(1402) := x"74df";block_ram_array(1404) := x"fffc";block_ram_array(1406) := x"b865";block_ram_array(1408) := x"004e";block_ram_array(1410) := x"eb7f";block_ram_array(1412) := x"006b";block_ram_array(1414) := x"3eea";block_ram_array(1416) := x"001e";block_ram_array(1418) := x"276f";block_ram_array(1420) := x"ffa9";block_ram_array(1422) := x"3e54";block_ram_array(1424) := x"ffde";block_ram_array(1426) := x"2438";block_ram_array(1428) := x"0003";block_ram_array(1430) := x"9605";block_ram_array(1432) := x"ffe3";block_ram_array(1434) := x"9621";block_ram_array(1436) := x"fff5";block_ram_array(1438) := x"e037";block_ram_array(1440) := x"0002";block_ram_array(1442) := x"9a55";block_ram_array(1444) := x"0053";block_ram_array(1446) := x"db8c";block_ram_array(1448) := x"0067";block_ram_array(1450) := x"9ceb";block_ram_array(1452) := x"ffbe";block_ram_array(1454) := x"a623";block_ram_array(1456) := x"ff83";block_ram_array(1458) := x"0a3a";block_ram_array(1460) := x"ffc5";block_ram_array(1462) := x"f9af";block_ram_array(1464) := x"0014";block_ram_array(1466) := x"c27f";block_ram_array(1468) := x"0079";block_ram_array(1470) := x"7d03";block_ram_array(1472) := x"0035";block_ram_array(1474) := x"e17f";block_ram_array(1476) := x"ffc8";block_ram_array(1478) := x"89ab";block_ram_array(1480) := x"fff7";block_ram_array(1482) := x"a974";block_ram_array(1484) := x"ffff";block_ram_array(1486) := x"ab61";block_ram_array(1488) := x"ffdf";block_ram_array(1490) := x"29c3";block_ram_array(1492) := x"ffc6";block_ram_array(1494) := x"83a5";block_ram_array(1496) := x"ffd2";block_ram_array(1498) := x"33c5";block_ram_array(1500) := x"0074";block_ram_array(1502) := x"a185";block_ram_array(1504) := x"0090";block_ram_array(1506) := x"8292";block_ram_array(1508) := x"ffd3";block_ram_array(1510) := x"2468";block_ram_array(1512) := x"ff8e";block_ram_array(1514) := x"deee";block_ram_array(1516) := x"ffb3";block_ram_array(1518) := x"29d0";block_ram_array(1520) := x"
0006";block_ram_array(1522) := x"017f";block_ram_array(1524) := x"0057";block_ram_array(1526) := x"3485";block_ram_array(1528) := x"000e";block_ram_array(1530) := x"70cb";block_ram_array(1532) := x"fff4";block_ram_array(1534) := x"266a";block_ram_array(1536) := x"0031";block_ram_array(1538) := x"388c";block_ram_array(1540) := x"0008";block_ram_array(1542) := x"d8ae";block_ram_array(1544) := x"ffd5";block_ram_array(1546) := x"74d1";block_ram_array(1548) := x"ffa3";block_ram_array(1550) := x"fd78";block_ram_array(1552) := x"ffbf";block_ram_array(1554) := x"2f20";block_ram_array(1556) := x"006c";block_ram_array(1558) := x"2664";block_ram_array(1560) := x"007a";block_ram_array(1562) := x"9e3f";block_ram_array(1564) := x"fffb";block_ram_array(1566) := x"4185";block_ram_array(1568) := x"ffca";block_ram_array(1570) := x"55ea";block_ram_array(1572) := x"ffb1";block_ram_array(1574) := x"f765";block_ram_array(1576) := x"ffec";block_ram_array(1578) := x"1b67";block_ram_array(1580) := x"002b";block_ram_array(1582) := x"e6b5";block_ram_array(1584) := x"fff7";block_ram_array(1586) := x"c63c";block_ram_array(1588) := x"0005";block_ram_array(1590) := x"5e48";block_ram_array(1592) := x"0034";block_ram_array(1594) := x"224c";block_ram_array(1596) := x"0029";block_ram_array(1598) := x"c796";block_ram_array(1600) := x"0006";block_ram_array(1602) := x"8e52";block_ram_array(1604) := x"ff91";block_ram_array(1606) := x"ac5a";block_ram_array(1608) := x"ff96";block_ram_array(1610) := x"bf26";block_ram_array(1612) := x"0048";block_ram_array(1614) := x"561b";block_ram_array(1616) := x"006c";block_ram_array(1618) := x"4990";block_ram_array(1620) := x"001d";block_ram_array(1622) := x"30c3";block_ram_array(1624) := x"ffdd";block_ram_array(1626) := x"5571";block_ram_array(1628) := x"ffc6";block_ram_array(1630) := x"7436";block_ram_array(1632) := x"000f";block_ram_array(1634) := x"803a";block_ram_array(1636) := x"000b";block_ram_array(1638) := x"aa0b";block_ram_array(1640) := x"ffc0";block_ram_array(1642) := x"422e";block_ram_array(1644) := x"fff0";block_ram_array(1646) := x"5e27";block_ram_array(1648) := x"003a";block_ram_array(1650) := x"a55e";block_ram_array(1652) := x"005a";block_ram_array(1654) := x"6770";block_ram_array(1656) := x"0020";block_ram_array(1658) := x"2a22";block_ram_array(1660) := x"ff8c";block_ram_array(1662) := x"84ea";block_ram_array(1664) := x"ffa4";block_ram_array(1666) := x"e046";block_ram_array(1668) := x"0029";block_ram_array(1670) := x"ce16";block_ram_array(1672) := x"0034";block_ram_array(1674) := x"8b91";block_ram_array(1676) := x"0016";block_ram_array(1678) := x"f38b";block_ram_array(1680) := x"fff6";block_ram_array(1682) := x"21a5";block_ram_array(1684) := x"fffd";block_ram_array(1686) := x"4da6";block_ram_array(1688) := x"002b";block_ram_array(1690) := x"3223";block_ram_array(1692) := x"ffeb";block_ram_array(1694) := x"20da";block_ram_array(1696) := x"ffb3";block_ram_array(1698) := x"29dc";block_ram_array(1700) := x"ffdc";block_ram_array(1702) := x"17c1";block_ram_array(1704) := x"0012";block_ram_array(1706) := x"a678";block_ram_array(1708) := x"0065";block_ram_array(1710) := x"94fa";block_ram_array(1712) := x"0044";block_ram_array(1714) := x"f459";block_ram_array(1716) := x"ffb8";block_ram_array(1718) := x"132c";block_ram_array(1720) := x"ffb7";block_ram_array(1722) := x"7607";block_ram_array(1724) := x"fff9";block_ram_array(1726) := x"ad98";block_ram_array(1728) := x"0015";block_ram_array(1730) := x"6ef8";block_ram_array(1732) := x"0011";block_ram_array(1734) := x"7331";block_ram_array(1736) := x"ffe2";block_ram_array(1738) := x"3ad7";block_ram_array(1740) := x"0016";block_ram_array(1742) := x"21d1";block_ram_array(1744) := x"0058";block_ram_array(1746) := x"ce84";block_ram_array(1748) := x"0002";block_ram_array(1750) := x"c4a7";block_ram_array(1752) := x"ffb2";block_ram_array(1754) := x"92e5";block_ram_array(1756) := x"ffa4";block_ram_array(1758) := x"9047";block_ram_array(1760) := x"ffee";block_ram_array(1762) := x"4a92";block_ram_array(1764) := x"0074";block_ram_array(1766) := x"90fa";block_ram_array(1768) := x"
0045";block_ram_array(1770) := x"51b4";block_ram_array(1772) := x"ffd2";block_ram_array(1774) := x"03d8";block_ram_array(1776) := x"ffe2";block_ram_array(1778) := x"7bf4";block_ram_array(1780) := x"fffe";block_ram_array(1782) := x"d19d";block_ram_array(1784) := x"0005";block_ram_array(1786) := x"1c60";block_ram_array(1788) := x"ffe3";block_ram_array(1790) := x"b348";block_ram_array(1792) := x"ffd4";block_ram_array(1794) := x"054c";block_ram_array(1796) := x"0026";block_ram_array(1798) := x"b6f9";block_ram_array(1800) := x"003a";block_ram_array(1802) := x"d54c";block_ram_array(1804) := x"0007";block_ram_array(1806) := x"5764";block_ram_array(1808) := x"ffe9";block_ram_array(1810) := x"e375";block_ram_array(1812) := x"ffe0";block_ram_array(1814) := x"3b51";block_ram_array(1816) := x"fffd";block_ram_array(1818) := x"d6de";block_ram_array(1820) := x"000e";block_ram_array(1822) := x"1a66";block_ram_array(1824) := x"fffe";block_ram_array(1826) := x"b2c6";block_ram_array(1828) := x"0000";block_ram_array(1830) := x"76e8";block_ram_array(1832) := x"0006";block_ram_array(1834) := x"2d4b";block_ram_array(1836) := x"fffe";block_ram_array(1838) := x"ba0d";block_ram_array(1840) := x"fff9";block_ram_array(1842) := x"ac50";block_ram_array(1844) := x"0000";block_ram_array(1846) := x"b612";block_ram_array(1848) := x"0006";block_ram_array(1850) := x"7829";block_ram_array(1852) := x"fffe";block_ram_array(1854) := x"e918";block_ram_array(1856) := x"fff9";block_ram_array(1858) := x"572b";block_ram_array(1860) := x"0001";block_ram_array(1862) := x"016e";block_ram_array(1864) := x"0006";block_ram_array(1866) := x"d13a";block_ram_array(1868) := x"ffff";block_ram_array(1870) := x"00a7";block_ram_array(1872) := x"fff8";block_ram_array(1874) := x"bd63";block_ram_array(1876) := x"0000";block_ram_array(1878) := x"79e4";block_ram_array(1880) := x"0006";block_ram_array(1882) := x"e119";block_ram_array(1884) := x"0000";block_ram_array(1886) := x"9453";block_ram_array(1888) := x"fff9";block_ram_array(1890) := x"f41e";block_ram_array(1892) := x"ffff";block_ram_array(1894) := x"2ec6";block_ram_array(1896) := x"0005";block_ram_array(1898) := x"975b";block_ram_array(1900) := x"0001";block_ram_array(1902) := x"160f";block_ram_array(1904) := x"fffb";block_ram_array(1906) := x"3d5b";block_ram_array(1908) := x"fffe";block_ram_array(1910) := x"e4f1";block_ram_array(1912) := x"0004";block_ram_array(1914) := x"4ab6";block_ram_array(1916) := x"0001";block_ram_array(1918) := x"0f29";block_ram_array(1920) := x"fffc";block_ram_array(1922) := x"bb79";block_ram_array(1924) := x"ffff";block_ram_array(1926) := x"4496";block_ram_array(1928) := x"0003";block_ram_array(1930) := x"1dc6";block_ram_array(1932) := x"ffff";block_ram_array(1934) := x"bf59";block_ram_array(1936) := x"fffc";block_ram_array(1938) := x"edce";block_ram_array(1940) := x"0000";block_ram_array(1942) := x"b1ac";block_ram_array(1944) := x"0003";block_ram_array(1946) := x"6006";block_ram_array(1948) := x"fffe";block_ram_array(1950) := x"80d3";block_ram_array(1952) := x"fffc";block_ram_array(1954) := x"14c0";block_ram_array(1956) := x"0001";block_ram_array(1958) := x"a264";block_ram_array(1960) := x"0004";block_ram_array(1962) := x"566f";block_ram_array(1964) := x"fffe";block_ram_array(1966) := x"1774";block_ram_array(1968) := x"fffa";block_ram_array(1970) := x"ef0a";block_ram_array(1972) := x"0001";block_ram_array(1974) := x"d646";block_ram_array(1976) := x"0005";block_ram_array(1978) := x"b77a";block_ram_array(1980) := x"fffe";block_ram_array(1982) := x"97b1";block_ram_array(1984) := x"fffa";block_ram_array(1986) := x"169c";block_ram_array(1988) := x"0000";block_ram_array(1990) := x"a024";block_ram_array(1992) := x"0006";block_ram_array(1994) := x"050e";block_ram_array(1996) := x"ffff";block_ram_array(1998) := x"cf16";block_ram_array(2000) := x"fffa";block_ram_array(2002) := x"0ef3";block_ram_array(2004) := x"ffff";block_ram_array(2006) := x"1451";block_ram_array(2008) := x"0004";block_ram_array(2010) := x"e1b4";block_ram_array(2012) := x"0001";block_ram_array(2014) := x"4e36";block_ram_array(2016) := x"
fffb";block_ram_array(2018) := x"7ddf";block_ram_array(2020) := x"fffe";block_ram_array(2022) := x"c5e4";block_ram_array(2024) := x"0003";block_ram_array(2026) := x"e134";block_ram_array(2028) := x"0001";block_ram_array(2030) := x"57fe";block_ram_array(2032) := x"fffc";block_ram_array(2034) := x"ace2";block_ram_array(2036) := x"ffff";block_ram_array(2038) := x"08f7";block_ram_array(2040) := x"0003";block_ram_array(2042) := x"09f4";block_ram_array(2044) := x"0000";block_ram_array(2046) := x"7dbe";block_ram_array(2048) := x"fffd";block_ram_array(2050) := x"0600";block_ram_array(2052) := x"0000";block_ram_array(2054) := x"0000";block_ram_array(2056) := x"0003";block_ram_array(2058) := x"09f4";block_ram_array(2060) := x"ffff";block_ram_array(2062) := x"8242";block_ram_array(2064) := x"fffc";block_ram_array(2066) := x"ace2";block_ram_array(2068) := x"0000";block_ram_array(2070) := x"f709";block_ram_array(2072) := x"0003";block_ram_array(2074) := x"e134";block_ram_array(2076) := x"fffe";block_ram_array(2078) := x"a802";block_ram_array(2080) := x"fffb";block_ram_array(2082) := x"7ddf";block_ram_array(2084) := x"0001";block_ram_array(2086) := x"3a1c";block_ram_array(2088) := x"0004";block_ram_array(2090) := x"e1b4";block_ram_array(2092) := x"fffe";block_ram_array(2094) := x"b1ca";block_ram_array(2096) := x"fffa";block_ram_array(2098) := x"0ef3";block_ram_array(2100) := x"0000";block_ram_array(2102) := x"ebaf";block_ram_array(2104) := x"0006";block_ram_array(2106) := x"050e";block_ram_array(2108) := x"0000";block_ram_array(2110) := x"30ea";block_ram_array(2112) := x"fffa";block_ram_array(2114) := x"169c";block_ram_array(2116) := x"ffff";block_ram_array(2118) := x"5fdc";block_ram_array(2120) := x"0005";block_ram_array(2122) := x"b77a";block_ram_array(2124) := x"0001";block_ram_array(2126) := x"684f";block_ram_array(2128) := x"fffa";block_ram_array(2130) := x"ef0a";block_ram_array(2132) := x"fffe";block_ram_array(2134) := x"29ba";block_ram_array(2136) := x"0004";block_ram_array(2138) := x"566f";block_ram_array(2140) := x"0001";block_ram_array(2142) := x"e88c";block_ram_array(2144) := x"fffc";block_ram_array(2146) := x"14c0";block_ram_array(2148) := x"fffe";block_ram_array(2150) := x"5d9c";block_ram_array(2152) := x"0003";block_ram_array(2154) := x"6006";block_ram_array(2156) := x"0001";block_ram_array(2158) := x"7f2d";block_ram_array(2160) := x"fffc";block_ram_array(2162) := x"edce";block_ram_array(2164) := x"ffff";block_ram_array(2166) := x"4e54";block_ram_array(2168) := x"0003";block_ram_array(2170) := x"1dc6";block_ram_array(2172) := x"0000";block_ram_array(2174) := x"40a7";block_ram_array(2176) := x"fffc";block_ram_array(2178) := x"bb79";block_ram_array(2180) := x"0000";block_ram_array(2182) := x"bb6a";block_ram_array(2184) := x"0004";block_ram_array(2186) := x"4ab6";block_ram_array(2188) := x"fffe";block_ram_array(2190) := x"f0d7";block_ram_array(2192) := x"fffb";block_ram_array(2194) := x"3d5b";block_ram_array(2196) := x"0001";block_ram_array(2198) := x"1b0f";block_ram_array(2200) := x"0005";block_ram_array(2202) := x"975b";block_ram_array(2204) := x"fffe";block_ram_array(2206) := x"e9f1";block_ram_array(2208) := x"fff9";block_ram_array(2210) := x"f41e";block_ram_array(2212) := x"0000";block_ram_array(2214) := x"d13a";block_ram_array(2216) := x"0006";block_ram_array(2218) := x"e119";block_ram_array(2220) := x"ffff";block_ram_array(2222) := x"6bad";block_ram_array(2224) := x"fff8";block_ram_array(2226) := x"bd63";block_ram_array(2228) := x"ffff";block_ram_array(2230) := x"861c";block_ram_array(2232) := x"0006";block_ram_array(2234) := x"d13a";block_ram_array(2236) := x"0000";block_ram_array(2238) := x"ff59";block_ram_array(2240) := x"fff9";block_ram_array(2242) := x"572b";block_ram_array(2244) := x"fffe";block_ram_array(2246) := x"fe92";block_ram_array(2248) := x"0006";block_ram_array(2250) := x"7829";block_ram_array(2252) := x"0001";block_ram_array(2254) := x"16e8";block_ram_array(2256) := x"fff9";block_ram_array(2258) := x"ac50";block_ram_array(2260) := x"ffff";block_ram_array(2262) := x"49ee";block_ram_array(2264) := x"
0006";block_ram_array(2266) := x"2d4b";block_ram_array(2268) := x"0001";block_ram_array(2270) := x"45f3";block_ram_array(2272) := x"fffe";block_ram_array(2274) := x"b2c6";block_ram_array(2276) := x"ffff";block_ram_array(2278) := x"8918";block_ram_array(2280) := x"fffd";block_ram_array(2282) := x"d6de";block_ram_array(2284) := x"fff1";block_ram_array(2286) := x"e59a";block_ram_array(2288) := x"ffe9";block_ram_array(2290) := x"e375";block_ram_array(2292) := x"001f";block_ram_array(2294) := x"c4af";block_ram_array(2296) := x"003a";block_ram_array(2298) := x"d54c";block_ram_array(2300) := x"fff8";block_ram_array(2302) := x"a89c";block_ram_array(2304) := x"ffd4";block_ram_array(2306) := x"054c";block_ram_array(2308) := x"ffd9";block_ram_array(2310) := x"4907";block_ram_array(2312) := x"0005";block_ram_array(2314) := x"1c60";block_ram_array(2316) := x"001c";block_ram_array(2318) := x"4cb8";block_ram_array(2320) := x"ffe2";block_ram_array(2322) := x"7bf4";block_ram_array(2324) := x"0001";block_ram_array(2326) := x"2e63";block_ram_array(2328) := x"0045";block_ram_array(2330) := x"51b4";block_ram_array(2332) := x"002d";block_ram_array(2334) := x"fc28";block_ram_array(2336) := x"ffee";block_ram_array(2338) := x"4a92";block_ram_array(2340) := x"ff8b";block_ram_array(2342) := x"6f06";block_ram_array(2344) := x"ffb2";block_ram_array(2346) := x"92e5";block_ram_array(2348) := x"005b";block_ram_array(2350) := x"6fb9";block_ram_array(2352) := x"0058";block_ram_array(2354) := x"ce84";block_ram_array(2356) := x"fffd";block_ram_array(2358) := x"3b59";block_ram_array(2360) := x"ffe2";block_ram_array(2362) := x"3ad7";block_ram_array(2364) := x"ffe9";block_ram_array(2366) := x"de2f";block_ram_array(2368) := x"0015";block_ram_array(2370) := x"6ef8";block_ram_array(2372) := x"ffee";block_ram_array(2374) := x"8ccf";block_ram_array(2376) := x"ffb7";block_ram_array(2378) := x"7607";block_ram_array(2380) := x"0006";block_ram_array(2382) := x"5268";block_ram_array(2384) := x"0044";block_ram_array(2386) := x"f459";block_ram_array(2388) := x"0047";block_ram_array(2390) := x"ecd4";block_ram_array(2392) := x"0012";block_ram_array(2394) := x"a678";block_ram_array(2396) := x"ff9a";block_ram_array(2398) := x"6b06";block_ram_array(2400) := x"ffb3";block_ram_array(2402) := x"29dc";block_ram_array(2404) := x"0023";block_ram_array(2406) := x"e83f";block_ram_array(2408) := x"002b";block_ram_array(2410) := x"3223";block_ram_array(2412) := x"0014";block_ram_array(2414) := x"df26";block_ram_array(2416) := x"fff6";block_ram_array(2418) := x"21a5";block_ram_array(2420) := x"0002";block_ram_array(2422) := x"b25a";block_ram_array(2424) := x"0034";block_ram_array(2426) := x"8b91";block_ram_array(2428) := x"ffe9";block_ram_array(2430) := x"0c75";block_ram_array(2432) := x"ffa4";block_ram_array(2434) := x"e046";block_ram_array(2436) := x"ffd6";block_ram_array(2438) := x"31ea";block_ram_array(2440) := x"0020";block_ram_array(2442) := x"2a22";block_ram_array(2444) := x"0073";block_ram_array(2446) := x"7b16";block_ram_array(2448) := x"003a";block_ram_array(2450) := x"a55e";block_ram_array(2452) := x"ffa5";block_ram_array(2454) := x"9890";block_ram_array(2456) := x"ffc0";block_ram_array(2458) := x"422e";block_ram_array(2460) := x"000f";block_ram_array(2462) := x"a1d9";block_ram_array(2464) := x"000f";block_ram_array(2466) := x"803a";block_ram_array(2468) := x"fff4";block_ram_array(2470) := x"55f5";block_ram_array(2472) := x"ffdd";block_ram_array(2474) := x"5571";block_ram_array(2476) := x"0039";block_ram_array(2478) := x"8bca";block_ram_array(2480) := x"006c";block_ram_array(2482) := x"4990";block_ram_array(2484) := x"ffe2";block_ram_array(2486) := x"cf3d";block_ram_array(2488) := x"ff96";block_ram_array(2490) := x"bf26";block_ram_array(2492) := x"ffb7";block_ram_array(2494) := x"a9e5";block_ram_array(2496) := x"0006";block_ram_array(2498) := x"8e52";block_ram_array(2500) := x"006e";block_ram_array(2502) := x"53a6";block_ram_array(2504) := x"0034";block_ram_array(2506) := x"224c";block_ram_array(2508) := x"ffd6";block_ram_array(2510) := x"386a";block_ram_array(2512) := x"
fff7";block_ram_array(2514) := x"c63c";block_ram_array(2516) := x"fffa";block_ram_array(2518) := x"a1b8";block_ram_array(2520) := x"ffec";block_ram_array(2522) := x"1b67";block_ram_array(2524) := x"ffd4";block_ram_array(2526) := x"194b";block_ram_array(2528) := x"ffca";block_ram_array(2530) := x"55ea";block_ram_array(2532) := x"004e";block_ram_array(2534) := x"089b";block_ram_array(2536) := x"007a";block_ram_array(2538) := x"9e3f";block_ram_array(2540) := x"0004";block_ram_array(2542) := x"be7b";block_ram_array(2544) := x"ffbf";block_ram_array(2546) := x"2f20";block_ram_array(2548) := x"ff93";block_ram_array(2550) := x"d99c";block_ram_array(2552) := x"ffd5";block_ram_array(2554) := x"74d1";block_ram_array(2556) := x"005c";block_ram_array(2558) := x"0288";block_ram_array(2560) := x"0031";block_ram_array(2562) := x"388c";block_ram_array(2564) := x"fff7";block_ram_array(2566) := x"2752";block_ram_array(2568) := x"000e";block_ram_array(2570) := x"70cb";block_ram_array(2572) := x"000b";block_ram_array(2574) := x"d996";block_ram_array(2576) := x"0006";block_ram_array(2578) := x"017f";block_ram_array(2580) := x"ffa8";block_ram_array(2582) := x"cb7b";block_ram_array(2584) := x"ff8e";block_ram_array(2586) := x"deee";block_ram_array(2588) := x"004c";block_ram_array(2590) := x"d630";block_ram_array(2592) := x"0090";block_ram_array(2594) := x"8292";block_ram_array(2596) := x"002c";block_ram_array(2598) := x"db98";block_ram_array(2600) := x"ffd2";block_ram_array(2602) := x"33c5";block_ram_array(2604) := x"ff8b";block_ram_array(2606) := x"5e7b";block_ram_array(2608) := x"ffdf";block_ram_array(2610) := x"29c3";block_ram_array(2612) := x"0039";block_ram_array(2614) := x"7c5b";block_ram_array(2616) := x"fff7";block_ram_array(2618) := x"a974";block_ram_array(2620) := x"0000";block_ram_array(2622) := x"549f";block_ram_array(2624) := x"0035";block_ram_array(2626) := x"e17f";block_ram_array(2628) := x"0037";block_ram_array(2630) := x"7655";block_ram_array(2632) := x"0014";block_ram_array(2634) := x"c27f";block_ram_array(2636) := x"ff86";block_ram_array(2638) := x"82fd";block_ram_array(2640) := x"ff83";block_ram_array(2642) := x"0a3a";block_ram_array(2644) := x"003a";block_ram_array(2646) := x"0651";block_ram_array(2648) := x"0067";block_ram_array(2650) := x"9ceb";block_ram_array(2652) := x"0041";block_ram_array(2654) := x"59dd";block_ram_array(2656) := x"0002";block_ram_array(2658) := x"9a55";block_ram_array(2660) := x"ffac";block_ram_array(2662) := x"2474";block_ram_array(2664) := x"ffe3";block_ram_array(2666) := x"9621";block_ram_array(2668) := x"000a";block_ram_array(2670) := x"1fc9";block_ram_array(2672) := x"ffde";block_ram_array(2674) := x"2438";block_ram_array(2676) := x"fffc";block_ram_array(2678) := x"69fb";block_ram_array(2680) := x"001e";block_ram_array(2682) := x"276f";block_ram_array(2684) := x"0056";block_ram_array(2686) := x"c1ac";block_ram_array(2688) := x"004e";block_ram_array(2690) := x"eb7f";block_ram_array(2692) := x"ff94";block_ram_array(2694) := x"c116";block_ram_array(2696) := x"ff70";block_ram_array(2698) := x"74df";block_ram_array(2700) := x"0003";block_ram_array(2702) := x"479b";block_ram_array(2704) := x"004e";block_ram_array(2706) := x"5d43";block_ram_array(2708) := x"0055";block_ram_array(2710) := x"f6de";block_ram_array(2712) := x"fffc";block_ram_array(2714) := x"91b4";block_ram_array(2716) := x"ffc6";block_ram_array(2718) := x"6bf2";block_ram_array(2720) := x"001e";block_ram_array(2722) := x"7242";block_ram_array(2724) := x"000b";block_ram_array(2726) := x"b964";block_ram_array(2728) := x"ffb7";block_ram_array(2730) := x"1c26";block_ram_array(2732) := x"ffbf";block_ram_array(2734) := x"7582";block_ram_array(2736) := x"0007";block_ram_array(2738) := x"8e80";block_ram_array(2740) := x"008a";block_ram_array(2742) := x"9e43";block_ram_array(2744) := x"0064";block_ram_array(2746) := x"6be1";block_ram_array(2748) := x"ff9c";block_ram_array(2750) := x"ed63";block_ram_array(2752) := x"ff96";block_ram_array(2754) := x"7196";block_ram_array(2756) := x"fff7";block_ram_array(2758) := x"710c";block_ram_array(2760) := x"
001e";block_ram_array(2762) := x"96fa";block_ram_array(2764) := x"0024";block_ram_array(2766) := x"6a66";block_ram_array(2768) := x"ffee";block_ram_array(2770) := x"5f52";block_ram_array(2772) := x"000b";block_ram_array(2774) := x"3865";block_ram_array(2776) := x"0049";block_ram_array(2778) := x"c5a5";block_ram_array(2780) := x"0001";block_ram_array(2782) := x"db36";block_ram_array(2784) := x"ffc1";block_ram_array(2786) := x"e472";block_ram_array(2788) := x"ffa4";block_ram_array(2790) := x"2f6c";block_ram_array(2792) := x"ffd0";block_ram_array(2794) := x"b24d";block_ram_array(2796) := x"0074";block_ram_array(2798) := x"e5c6";block_ram_array(2800) := x"0070";block_ram_array(2802) := x"769f";block_ram_array(2804) := x"ffe4";block_ram_array(2806) := x"e219";block_ram_array(2808) := x"ffc1";block_ram_array(2810) := x"18da";block_ram_array(2812) := x"ffd3";block_ram_array(2814) := x"72c5";block_ram_array(2816) := x"0011";block_ram_array(2818) := x"fd6f";block_ram_array(2820) := x"000d";block_ram_array(2822) := x"a74e";block_ram_array(2824) := x"ffba";block_ram_array(2826) := x"3dc5";block_ram_array(2828) := x"000a";block_ram_array(2830) := x"4bff";block_ram_array(2832) := x"0070";block_ram_array(2834) := x"6a66";block_ram_array(2836) := x"0049";block_ram_array(2838) := x"57a2";block_ram_array(2840) := x"ffe2";block_ram_array(2842) := x"91b4";block_ram_array(2844) := x"ff5d";block_ram_array(2846) := x"6487";block_ram_array(2848) := x"ffa6";block_ram_array(2850) := x"ed57";block_ram_array(2852) := x"0078";block_ram_array(2854) := x"5ec7";block_ram_array(2856) := x"0059";block_ram_array(2858) := x"88cb";block_ram_array(2860) := x"ffef";block_ram_array(2862) := x"f2a8";block_ram_array(2864) := x"ffed";block_ram_array(2866) := x"2141";block_ram_array(2868) := x"000a";block_ram_array(2870) := x"43c9";block_ram_array(2872) := x"0027";block_ram_array(2874) := x"8b29";block_ram_array(2876) := x"ffb6";block_ram_array(2878) := x"8721";block_ram_array(2880) := x"ff78";block_ram_array(2882) := x"89bc";block_ram_array(2884) := x"0026";block_ram_array(2886) := x"2358";block_ram_array(2888) := x"0080";block_ram_array(2890) := x"3d40";block_ram_array(2892) := x"0061";block_ram_array(2894) := x"212d";block_ram_array(2896) := x"000a";block_ram_array(2898) := x"6b53";block_ram_array(2900) := x"ff6f";block_ram_array(2902) := x"df01";block_ram_array(2904) := x"ffa3";block_ram_array(2906) := x"6a9a";block_ram_array(2908) := x"002a";block_ram_array(2910) := x"2182";block_ram_array(2912) := x"001c";block_ram_array(2914) := x"c09c";block_ram_array(2916) := x"0020";block_ram_array(2918) := x"bdb3";block_ram_array(2920) := x"0014";block_ram_array(2922) := x"ae99";block_ram_array(2924) := x"001d";block_ram_array(2926) := x"ae39";block_ram_array(2928) := x"0047";block_ram_array(2930) := x"d13b";block_ram_array(2932) := x"ffaf";block_ram_array(2934) := x"2834";block_ram_array(2936) := x"ff59";block_ram_array(2938) := x"2825";block_ram_array(2940) := x"ffe3";block_ram_array(2942) := x"443b";block_ram_array(2944) := x"0057";block_ram_array(2946) := x"3c0f";block_ram_array(2948) := x"00af";block_ram_array(2950) := x"1588";block_ram_array(2952) := x"0046";block_ram_array(2954) := x"fa20";block_ram_array(2956) := x"ff64";block_ram_array(2958) := x"9498";block_ram_array(2960) := x"ffa5";block_ram_array(2962) := x"acec";block_ram_array(2964) := x"001d";block_ram_array(2966) := x"a6ae";block_ram_array(2968) := x"fffc";block_ram_array(2970) := x"d3d6";block_ram_array(2972) := x"ffed";block_ram_array(2974) := x"bdb7";block_ram_array(2976) := x"fff5";block_ram_array(2978) := x"e0b9";block_ram_array(2980) := x"0079";block_ram_array(2982) := x"d73e";block_ram_array(2984) := x"009b";block_ram_array(2986) := x"9840";block_ram_array(2988) := x"ff89";block_ram_array(2990) := x"a64a";block_ram_array(2992) := x"ff30";block_ram_array(2994) := x"4d88";block_ram_array(2996) := x"ffce";block_ram_array(2998) := x"bac3";block_ram_array(3000) := x"0045";block_ram_array(3002) := x"ed0b";block_ram_array(3004) := x"00a0";block_ram_array(3006) := x"5039";block_ram_array(3008) := x"
0038";block_ram_array(3010) := x"23ce";block_ram_array(3012) := x"ffaf";block_ram_array(3014) := x"efd1";block_ram_array(3016) := x"fff7";block_ram_array(3018) := x"974c";block_ram_array(3020) := x"ffed";block_ram_array(3022) := x"8ca3";block_ram_array(3024) := x"ffbc";block_ram_array(3026) := x"bcfd";block_ram_array(3028) := x"ffd4";block_ram_array(3030) := x"c8db";block_ram_array(3032) := x"ffea";block_ram_array(3034) := x"7bca";block_ram_array(3036) := x"008c";block_ram_array(3038) := x"2c9d";block_ram_array(3040) := x"00aa";block_ram_array(3042) := x"e122";block_ram_array(3044) := x"ffc2";block_ram_array(3046) := x"7563";block_ram_array(3048) := x"ff69";block_ram_array(3050) := x"e8d5";block_ram_array(3052) := x"ff88";block_ram_array(3054) := x"b683";block_ram_array(3056) := x"fff8";block_ram_array(3058) := x"07ff";block_ram_array(3060) := x"00a0";block_ram_array(3062) := x"984d";block_ram_array(3064) := x"0041";block_ram_array(3066) := x"54c7";block_ram_array(3068) := x"ffc9";block_ram_array(3070) := x"476c";block_ram_array(3072) := x"0010";block_ram_array(3074) := x"3900";block_ram_array(3076) := x"001a";block_ram_array(3078) := x"9f00";block_ram_array(3080) := x"ffe9";block_ram_array(3082) := x"1cdc";block_ram_array(3084) := x"ff78";block_ram_array(3086) := x"3640";block_ram_array(3088) := x"ff81";block_ram_array(3090) := x"7023";block_ram_array(3092) := x"00ad";block_ram_array(3094) := x"4bed";block_ram_array(3096) := x"00e5";block_ram_array(3098) := x"24cf";block_ram_array(3100) := x"ffe3";block_ram_array(3102) := x"1cd1";block_ram_array(3104) := x"ff71";block_ram_array(3106) := x"646e";block_ram_array(3108) := x"ff90";block_ram_array(3110) := x"214b";block_ram_array(3112) := x"0017";block_ram_array(3114) := x"0ff9";block_ram_array(3116) := x"0052";block_ram_array(3118) := x"97c9";block_ram_array(3120) := x"ffd0";block_ram_array(3122) := x"031a";block_ram_array(3124) := x"fff7";block_ram_array(3126) := x"02bb";block_ram_array(3128) := x"0070";block_ram_array(3130) := x"49eb";block_ram_array(3132) := x"0048";block_ram_array(3134) := x"dbb2";block_ram_array(3136) := x"ffe6";block_ram_array(3138) := x"1dd7";block_ram_array(3140) := x"ff4a";block_ram_array(3142) := x"44db";block_ram_array(3144) := x"ff78";block_ram_array(3146) := x"9c5a";block_ram_array(3148) := x"0082";block_ram_array(3150) := x"11bb";block_ram_array(3152) := x"0097";block_ram_array(3154) := x"669c";block_ram_array(3156) := x"0022";block_ram_array(3158) := x"c1c4";block_ram_array(3160) := x"ffdd";block_ram_array(3162) := x"1038";block_ram_array(3164) := x"ffa6";block_ram_array(3166) := x"ea58";block_ram_array(3168) := x"0001";block_ram_array(3170) := x"e521";block_ram_array(3172) := x"0011";block_ram_array(3174) := x"b59a";block_ram_array(3176) := x"ffac";block_ram_array(3178) := x"1c35";block_ram_array(3180) := x"ffe3";block_ram_array(3182) := x"c5ac";block_ram_array(3184) := x"0048";block_ram_array(3186) := x"6e18";block_ram_array(3188) := x"00a5";block_ram_array(3190) := x"96e0";block_ram_array(3192) := x"0064";block_ram_array(3194) := x"0cd9";block_ram_array(3196) := x"ff29";block_ram_array(3198) := x"e610";block_ram_array(3200) := x"ff26";block_ram_array(3202) := x"fb4c";block_ram_array(3204) := x"0048";block_ram_array(3206) := x"1e45";block_ram_array(3208) := x"008d";block_ram_array(3210) := x"e737";block_ram_array(3212) := x"0039";block_ram_array(3214) := x"46d1";block_ram_array(3216) := x"ffc8";block_ram_array(3218) := x"05d4";block_ram_array(3220) := x"fff2";block_ram_array(3222) := x"b172";block_ram_array(3224) := x"0086";block_ram_array(3226) := x"35db";block_ram_array(3228) := x"ffd7";block_ram_array(3230) := x"8e0a";block_ram_array(3232) := x"ff21";block_ram_array(3234) := x"4eee";block_ram_array(3236) := x"ffa8";block_ram_array(3238) := x"6455";block_ram_array(3240) := x"0065";block_ram_array(3242) := x"0c59";block_ram_array(3244) := x"00fe";block_ram_array(3246) := x"f590";block_ram_array(3248) := x"0071";block_ram_array(3250) := x"d039";block_ram_array(3252) := x"ff32";block_ram_array(3254) := x"9a63";block_ram_array(3256) := x"
ff75";block_ram_array(3258) := x"d53c";block_ram_array(3260) := x"000f";block_ram_array(3262) := x"125a";block_ram_array(3264) := x"0003";block_ram_array(3266) := x"f2b8";block_ram_array(3268) := x"0015";block_ram_array(3270) := x"fd70";block_ram_array(3272) := x"fffa";block_ram_array(3274) := x"9c1a";block_ram_array(3276) := x"0062";block_ram_array(3278) := x"e291";block_ram_array(3280) := x"00b2";block_ram_array(3282) := x"55d4";block_ram_array(3284) := x"ffb0";block_ram_array(3286) := x"9ac0";block_ram_array(3288) := x"ff2a";block_ram_array(3290) := x"d7d7";block_ram_array(3292) := x"ff65";block_ram_array(3294) := x"4b52";block_ram_array(3296) := x"ffee";block_ram_array(3298) := x"394c";block_ram_array(3300) := x"011f";block_ram_array(3302) := x"92bc";block_ram_array(3304) := x"00d4";block_ram_array(3306) := x"5d8e";block_ram_array(3308) := x"ff7d";block_ram_array(3310) := x"0b3b";block_ram_array(3312) := x"ff7d";block_ram_array(3314) := x"58aa";block_ram_array(3316) := x"ffd0";block_ram_array(3318) := x"68aa";block_ram_array(3320) := x"fffe";block_ram_array(3322) := x"c929";block_ram_array(3324) := x"ffe4";block_ram_array(3326) := x"bd13";block_ram_array(3328) := x"ff88";block_ram_array(3330) := x"47fe";block_ram_array(3332) := x"00a5";block_ram_array(3334) := x"00f8";block_ram_array(3336) := x"014f";block_ram_array(3338) := x"e446";block_ram_array(3340) := x"ffe2";block_ram_array(3342) := x"512a";block_ram_array(3344) := x"feef";block_ram_array(3346) := x"838a";block_ram_array(3348) := x"fef5";block_ram_array(3350) := x"e188";block_ram_array(3352) := x"ffe9";block_ram_array(3354) := x"0994";block_ram_array(3356) := x"013d";block_ram_array(3358) := x"a992";block_ram_array(3360) := x"008b";block_ram_array(3362) := x"89f2";block_ram_array(3364) := x"ff9e";block_ram_array(3366) := x"c9cd";block_ram_array(3368) := x"0011";block_ram_array(3370) := x"c175";block_ram_array(3372) := x"ffff";block_ram_array(3374) := x"6296";block_ram_array(3376) := x"ffb2";block_ram_array(3378) := x"8fff";block_ram_array(3380) := x"ff54";block_ram_array(3382) := x"c043";block_ram_array(3384) := x"ff65";block_ram_array(3386) := x"4aea";block_ram_array(3388) := x"0103";block_ram_array(3390) := x"4fe8";block_ram_array(3392) := x"0157";block_ram_array(3394) := x"b4c8";block_ram_array(3396) := x"fff2";block_ram_array(3398) := x"4a70";block_ram_array(3400) := x"ff4e";block_ram_array(3402) := x"f55f";block_ram_array(3404) := x"fef5";block_ram_array(3406) := x"ab5e";block_ram_array(3408) := x"ff95";block_ram_array(3410) := x"ac8a";block_ram_array(3412) := x"00d7";block_ram_array(3414) := x"828d";block_ram_array(3416) := x"0070";block_ram_array(3418) := x"a745";block_ram_array(3420) := x"ffff";block_ram_array(3422) := x"5583";block_ram_array(3424) := x"0037";block_ram_array(3426) := x"1c79";block_ram_array(3428) := x"0017";block_ram_array(3430) := x"0cc3";block_ram_array(3432) := x"0007";block_ram_array(3434) := x"78a9";block_ram_array(3436) := x"ff1a";block_ram_array(3438) := x"791a";block_ram_array(3440) := x"fed7";block_ram_array(3442) := x"8734";block_ram_array(3444) := x"00ce";block_ram_array(3446) := x"89f6";block_ram_array(3448) := x"0187";block_ram_array(3450) := x"a9d0";block_ram_array(3452) := x"0069";block_ram_array(3454) := x"6355";block_ram_array(3456) := x"ff60";block_ram_array(3458) := x"7c13";block_ram_array(3460) := x"fed4";block_ram_array(3462) := x"b9ee";block_ram_array(3464) := x"ffe0";block_ram_array(3466) := x"71f4";block_ram_array(3468) := x"00b0";block_ram_array(3470) := x"9d54";block_ram_array(3472) := x"ffc5";block_ram_array(3474) := x"9404";block_ram_array(3476) := x"ffc7";block_ram_array(3478) := x"2575";block_ram_array(3480) := x"0095";block_ram_array(3482) := x"9044";block_ram_array(3484) := x"00cc";block_ram_array(3486) := x"6682";block_ram_array(3488) := x"0030";block_ram_array(3490) := x"f991";block_ram_array(3492) := x"fe91";block_ram_array(3494) := x"4fd0";block_ram_array(3496) := x"fec3";block_ram_array(3498) := x"cee8";block_ram_array(3500) := x"00d7";block_ram_array(3502) := x"6bff";block_ram_array(3504) := x"
011f";block_ram_array(3506) := x"1312";block_ram_array(3508) := x"004f";block_ram_array(3510) := x"40ed";block_ram_array(3512) := x"ffbc";block_ram_array(3514) := x"950d";block_ram_array(3516) := x"ff78";block_ram_array(3518) := x"b487";block_ram_array(3520) := x"0021";block_ram_array(3522) := x"0f4d";block_ram_array(3524) := x"0001";block_ram_array(3526) := x"d519";block_ram_array(3528) := x"ff54";block_ram_array(3530) := x"9c60";block_ram_array(3532) := x"ffd5";block_ram_array(3534) := x"84b1";block_ram_array(3536) := x"0076";block_ram_array(3538) := x"1659";block_ram_array(3540) := x"010f";block_ram_array(3542) := x"81a0";block_ram_array(3544) := x"00b3";block_ram_array(3546) := x"653b";block_ram_array(3548) := x"fec7";block_ram_array(3550) := x"d414";block_ram_array(3552) := x"feab";block_ram_array(3554) := x"cb96";block_ram_array(3556) := x"0037";block_ram_array(3558) := x"322c";block_ram_array(3560) := x"00c3";block_ram_array(3562) := x"1b14";block_ram_array(3564) := x"0089";block_ram_array(3566) := x"c799";block_ram_array(3568) := x"ffb8";block_ram_array(3570) := x"bcba";block_ram_array(3572) := x"ffc9";block_ram_array(3574) := x"e4ea";block_ram_array(3576) := x"00cf";block_ram_array(3578) := x"3d6b";block_ram_array(3580) := x"fff8";block_ram_array(3582) := x"e6e5";block_ram_array(3584) := x"fec3";block_ram_array(3586) := x"af74";block_ram_array(3588) := x"ff23";block_ram_array(3590) := x"6552";block_ram_array(3592) := x"0055";block_ram_array(3594) := x"222c";block_ram_array(3596) := x"01ce";block_ram_array(3598) := x"3578";block_ram_array(3600) := x"00f4";block_ram_array(3602) := x"dc30";block_ram_array(3604) := x"fea7";block_ram_array(3606) := x"507a";block_ram_array(3608) := x"ff04";block_ram_array(3610) := x"1d6d";block_ram_array(3612) := x"0031";block_ram_array(3614) := x"9164";block_ram_array(3616) := x"0031";block_ram_array(3618) := x"83a4";block_ram_array(3620) := x"ffea";block_ram_array(3622) := x"0072";block_ram_array(3624) := x"ffa4";block_ram_array(3626) := x"a316";block_ram_array(3628) := x"00cc";block_ram_array(3630) := x"d3df";block_ram_array(3632) := x"016f";block_ram_array(3634) := x"3b20";block_ram_array(3636) := x"ff7e";block_ram_array(3638) := x"6256";block_ram_array(3640) := x"fe81";block_ram_array(3642) := x"2ac2";block_ram_array(3644) := x"ff03";block_ram_array(3646) := x"efd0";block_ram_array(3648) := x"0004";block_ram_array(3650) := x"f92f";block_ram_array(3652) := x"01ac";block_ram_array(3654) := x"ad5a";block_ram_array(3656) := x"010c";block_ram_array(3658) := x"f616";block_ram_array(3660) := x"ff58";block_ram_array(3662) := x"8411";block_ram_array(3664) := x"ff89";block_ram_array(3666) := x"8667";block_ram_array(3668) := x"ffaf";block_ram_array(3670) := x"79b8";block_ram_array(3672) := x"ffc0";block_ram_array(3674) := x"f7e2";block_ram_array(3676) := x"ffbc";block_ram_array(3678) := x"0d29";block_ram_array(3680) := x"ff61";block_ram_array(3682) := x"864e";block_ram_array(3684) := x"010e";block_ram_array(3686) := x"3c50";block_ram_array(3688) := x"01ea";block_ram_array(3690) := x"0f1a";block_ram_array(3692) := x"ffde";block_ram_array(3694) := x"9699";block_ram_array(3696) := x"fe8c";block_ram_array(3698) := x"2d76";block_ram_array(3700) := x"fe5b";block_ram_array(3702) := x"61b4";block_ram_array(3704) := x"ffb2";block_ram_array(3706) := x"4dd4";block_ram_array(3708) := x"01e0";block_ram_array(3710) := x"7636";block_ram_array(3712) := x"00e9";block_ram_array(3714) := x"0dd6";block_ram_array(3716) := x"ff6e";block_ram_array(3718) := x"e672";block_ram_array(3720) := x"000e";block_ram_array(3722) := x"723b";block_ram_array(3724) := x"0013";block_ram_array(3726) := x"c5b1";block_ram_array(3728) := x"ffa5";block_ram_array(3730) := x"0b97";block_ram_array(3732) := x"fed5";block_ram_array(3734) := x"b138";block_ram_array(3736) := x"feec";block_ram_array(3738) := x"a1f0";block_ram_array(3740) := x"01b1";block_ram_array(3742) := x"f766";block_ram_array(3744) := x"023a";block_ram_array(3746) := x"6fb8";block_ram_array(3748) := x"ffbe";block_ram_array(3750) := x"d942";block_ram_array(3752) := x"
feb0";block_ram_array(3754) := x"66b0";block_ram_array(3756) := x"fe9d";block_ram_array(3758) := x"01e2";block_ram_array(3760) := x"ffb7";block_ram_array(3762) := x"8166";block_ram_array(3764) := x"0121";block_ram_array(3766) := x"8714";block_ram_array(3768) := x"004c";block_ram_array(3770) := x"f538";block_ram_array(3772) := x"0011";block_ram_array(3774) := x"03a6";block_ram_array(3776) := x"00b1";block_ram_array(3778) := x"7f9a";block_ram_array(3780) := x"0015";block_ram_array(3782) := x"8425";block_ram_array(3784) := x"ff99";block_ram_array(3786) := x"c7a9";block_ram_array(3788) := x"feab";block_ram_array(3790) := x"2d8c";block_ram_array(3792) := x"fec2";block_ram_array(3794) := x"0d58";block_ram_array(3796) := x"0159";block_ram_array(3798) := x"24bc";block_ram_array(3800) := x"01e9";block_ram_array(3802) := x"7c84";block_ram_array(3804) := x"004d";block_ram_array(3806) := x"9a5a";block_ram_array(3808) := x"ff3e";block_ram_array(3810) := x"c046";block_ram_array(3812) := x"fe90";block_ram_array(3814) := x"d906";block_ram_array(3816) := x"ffb2";block_ram_array(3818) := x"e761";block_ram_array(3820) := x"00d7";block_ram_array(3822) := x"0950";block_ram_array(3824) := x"ffd7";block_ram_array(3826) := x"7ba9";block_ram_array(3828) := x"ffda";block_ram_array(3830) := x"b815";block_ram_array(3832) := x"00c2";block_ram_array(3834) := x"98c4";block_ram_array(3836) := x"00e1";block_ram_array(3838) := x"0130";block_ram_array(3840) := x"0024";block_ram_array(3842) := x"2147";block_ram_array(3844) := x"fe22";block_ram_array(3846) := x"d6b0";block_ram_array(3848) := x"fe68";block_ram_array(3850) := x"73be";block_ram_array(3852) := x"014b";block_ram_array(3854) := x"d760";block_ram_array(3856) := x"01a7";block_ram_array(3858) := x"ef18";block_ram_array(3860) := x"002d";block_ram_array(3862) := x"9155";block_ram_array(3864) := x"ff5f";block_ram_array(3866) := x"250c";block_ram_array(3868) := x"ff65";block_ram_array(3870) := x"25be";block_ram_array(3872) := x"005d";block_ram_array(3874) := x"ac98";block_ram_array(3876) := x"fffd";block_ram_array(3878) := x"2f7c";block_ram_array(3880) := x"fef4";block_ram_array(3882) := x"93c0";block_ram_array(3884) := x"ffee";block_ram_array(3886) := x"3b5d";block_ram_array(3888) := x"00fa";block_ram_array(3890) := x"9408";block_ram_array(3892) := x"0126";block_ram_array(3894) := x"a9a8";block_ram_array(3896) := x"004f";block_ram_array(3898) := x"78de";block_ram_array(3900) := x"fe72";block_ram_array(3902) := x"4a5c";block_ram_array(3904) := x"fece";block_ram_array(3906) := x"acb0";block_ram_array(3908) := x"008e";block_ram_array(3910) := x"aa1c";block_ram_array(3912) := x"00b7";block_ram_array(3914) := x"83ee";block_ram_array(3916) := x"005b";block_ram_array(3918) := x"5593";block_ram_array(3920) := x"ffd5";block_ram_array(3922) := x"9613";block_ram_array(3924) := x"ffe6";block_ram_array(3926) := x"d855";block_ram_array(3928) := x"00af";block_ram_array(3930) := x"c38a";block_ram_array(3932) := x"ffcd";block_ram_array(3934) := x"03b7";block_ram_array(3936) := x"fec8";block_ram_array(3938) := x"a102";block_ram_array(3940) := x"ff51";block_ram_array(3942) := x"a40c";block_ram_array(3944) := x"0062";block_ram_array(3946) := x"7dde";block_ram_array(3948) := x"01bd";block_ram_array(3950) := x"dae0";block_ram_array(3952) := x"00f6";block_ram_array(3954) := x"882b";block_ram_array(3956) := x"fe97";block_ram_array(3958) := x"6f5c";block_ram_array(3960) := x"fee5";block_ram_array(3962) := x"cf48";block_ram_array(3964) := x"0048";block_ram_array(3966) := x"8264";block_ram_array(3968) := x"0061";block_ram_array(3970) := x"9f7d";block_ram_array(3972) := x"ffdd";block_ram_array(3974) := x"cfd9";block_ram_array(3976) := x"ff70";block_ram_array(3978) := x"95f2";block_ram_array(3980) := x"00ce";block_ram_array(3982) := x"4c48";block_ram_array(3984) := x"01a4";block_ram_array(3986) := x"c740";block_ram_array(3988) := x"ff80";block_ram_array(3990) := x"173c";block_ram_array(3992) := x"fe45";block_ram_array(3994) := x"c672";block_ram_array(3996) := x"ff00";block_ram_array(3998) := x"da39";block_ram_array(4000) := x"
004b";block_ram_array(4002) := x"cc6d";block_ram_array(4004) := x"01b4";block_ram_array(4006) := x"e1f0";block_ram_array(4008) := x"00bb";block_ram_array(4010) := x"8d8c";block_ram_array(4012) := x"ff3d";block_ram_array(4014) := x"82e4";block_ram_array(4016) := x"ffd2";block_ram_array(4018) := x"da51";block_ram_array(4020) := x"ffe4";block_ram_array(4022) := x"8506";block_ram_array(4024) := x"ff91";block_ram_array(4026) := x"9cb9";block_ram_array(4028) := x"ff7c";block_ram_array(4030) := x"8455";block_ram_array(4032) := x"ff7e";block_ram_array(4034) := x"6a30";block_ram_array(4036) := x"013e";block_ram_array(4038) := x"6356";block_ram_array(4040) := x"01c2";block_ram_array(4042) := x"83be";block_ram_array(4044) := x"ffbc";block_ram_array(4046) := x"f655";block_ram_array(4048) := x"fec1";block_ram_array(4050) := x"4c08";block_ram_array(4052) := x"fe8c";block_ram_array(4054) := x"d820";block_ram_array(4056) := x"ff90";block_ram_array(4058) := x"690e";block_ram_array(4060) := x"0197";block_ram_array(4062) := x"70a4";block_ram_array(4064) := x"00e7";block_ram_array(4066) := x"072d";block_ram_array(4068) := x"ffab";block_ram_array(4070) := x"e67c";block_ram_array(4072) := x"0011";block_ram_array(4074) := x"6d93";block_ram_array(4076) := x"ffff";block_ram_array(4078) := x"0aa7";block_ram_array(4080) := x"ffc7";block_ram_array(4082) := x"7700";block_ram_array(4084) := x"fedf";block_ram_array(4086) := x"71a8";block_ram_array(4088) := x"feb9";block_ram_array(4090) := x"a290";block_ram_array(4092) := x"0186";block_ram_array(4094) := x"58d0";
        --------------------
        --=1
        --------------------
        block_ram_array(4096) := x"ff62";block_ram_array(4098) := x"5c00";block_ram_array(4100) := x"0000";block_ram_array(4102) := x"0000";block_ram_array(4104) := x"ffe1";block_ram_array(4106) := x"e677";block_ram_array(4108) := x"0007";block_ram_array(4110) := x"0854";block_ram_array(4112) := x"fedb";block_ram_array(4114) := x"e084";block_ram_array(4116) := x"000c";block_ram_array(4118) := x"2c90";block_ram_array(4120) := x"ffbe";block_ram_array(4122) := x"7053";block_ram_array(4124) := x"01b8";block_ram_array(4126) := x"88ee";block_ram_array(4128) := x"012b";block_ram_array(4130) := x"c338";block_ram_array(4132) := x"009a";block_ram_array(4134) := x"d2ea";block_ram_array(4136) := x"00a3";block_ram_array(4138) := x"e932";block_ram_array(4140) := x"ffe9";block_ram_array(4142) := x"bc5d";block_ram_array(4144) := x"007b";block_ram_array(4146) := x"e3a5";block_ram_array(4148) := x"ffdb";block_ram_array(4150) := x"8fb9";block_ram_array(4152) := x"009e";block_ram_array(4154) := x"202a";block_ram_array(4156) := x"ffe6";block_ram_array(4158) := x"c73e";block_ram_array(4160) := x"00cb";block_ram_array(4162) := x"83e8";block_ram_array(4164) := x"ff0a";block_ram_array(4166) := x"06fd";block_ram_array(4168) := x"ff85";block_ram_array(4170) := x"029e";block_ram_array(4172) := x"fe8c";block_ram_array(4174) := x"d05a";block_ram_array(4176) := x"fe8b";block_ram_array(4178) := x"924e";block_ram_array(4180) := x"ff9f";block_ram_array(4182) := x"0dfb";block_ram_array(4184) := x"ff4a";block_ram_array(4186) := x"73c2";block_ram_array(4188) := x"00dd";block_ram_array(4190) := x"983e";block_ram_array(4192) := x"0016";block_ram_array(4194) := x"5fb5";block_ram_array(4196) := x"0034";block_ram_array(4198) := x"72ae";block_ram_array(4200) := x"ff8b";block_ram_array(4202) := x"21e8";block_ram_array(4204) := x"0046";block_ram_array(4206) := x"a808";block_ram_array(4208) := x"ffd6";block_ram_array(4210) := x"8a59";block_ram_array(4212) := x"007c";block_ram_array(4214) := x"2d5c";block_ram_array(4216) := x"ffef";block_ram_array(4218) := x"a695";block_ram_array(4220) := x"0105";block_ram_array(4222) := x"c0cc";block_ram_array(4224) := x"0152";block_ram_array(4226) := x"9a94";block_ram_array(4228) := x"0085";block_ram_array(4230) := x"4e9b";block_ram_array(4232) := x"0087";block_ram_array(4234) := x"7fbe";block_ram_array(4236) := x"ff6a";block_ram_array(4238) := x"cbf0";block_ram_array(4240) := x"0067";block_ram_array(4242) := x"cdc9";block_ram_array(4244) := x"ffb9";block_ram_array(4246) := x"5117";block_ram_array(4248) := x"000e";block_ram_array(4250) := x"81fd";block_ram_array(4252) := x"ff9a";block_ram_array(4254) := x"3830";block_ram_array(4256) := x"00bf";block_ram_array(4258) := x"e531";block_ram_array(4260) := x"ff88";block_ram_array(4262) := x"4dec";block_ram_array(4264) := x"ff48";block_ram_array(4266) := x"c60c";block_ram_array(4268) := x"fe27";block_ram_array(4270) := x"65a4";block_ram_array(4272) := x"fe31";block_ram_array(4274) := x"3fe0";block_ram_array(4276) := x"005f";block_ram_array(4278) := x"1263";block_ram_array(4280) := x"ff93";block_ram_array(4282) := x"8e22";block_ram_array(4284) := x"00d6";block_ram_array(4286) := x"b0ca";block_ram_array(4288) := x"fff0";block_ram_array(4290) := x"778f";block_ram_array(4292) := x"00ce";block_ram_array(4294) := x"fd0f";block_ram_array(4296) := x"0048";block_ram_array(4298) := x"7922";block_ram_array(4300) := x"004b";block_ram_array(4302) := x"5e5c";block_ram_array(4304) := x"fff7";block_ram_array(4306) := x"c82c";block_ram_array(4308) := x"007e";block_ram_array(4310) := x"14d4";block_ram_array(4312) := x"008a";block_ram_array(4314) := x"dc30";block_ram_array(4316) := x"009d";block_ram_array(4318) := x"0c10";block_ram_array(4320) := x"0121";block_ram_array(4322) := x"d5ee";block_ram_array(4324) := x"0014";block_ram_array(4326) := x"bd05";block_ram_array(4328) := x"0075";block_ram_array(4330) := x"05d7";block_ram_array(4332) := x"fede";block_ram_array(4334) := x"371a";block_ram_array(4336) := x"ff97";block_ram_array(4338) := x"e80e";block_ram_array(4340) := x"ffd7";block_ram_array(4342) := x"
fd19";block_ram_array(4344) := x"0048";block_ram_array(4346) := x"b36b";block_ram_array(4348) := x"ff99";block_ram_array(4350) := x"21d9";block_ram_array(4352) := x"ffc0";block_ram_array(4354) := x"d64b";block_ram_array(4356) := x"ffb1";block_ram_array(4358) := x"beb5";block_ram_array(4360) := x"fff2";block_ram_array(4362) := x"fc98";block_ram_array(4364) := x"ff05";block_ram_array(4366) := x"c286";block_ram_array(4368) := x"fdf4";block_ram_array(4370) := x"0404";block_ram_array(4372) := x"ffe0";block_ram_array(4374) := x"5d1d";block_ram_array(4376) := x"ffc2";block_ram_array(4378) := x"7e4a";block_ram_array(4380) := x"01cb";block_ram_array(4382) := x"10f0";block_ram_array(4384) := x"0084";block_ram_array(4386) := x"d254";block_ram_array(4388) := x"0064";block_ram_array(4390) := x"712a";block_ram_array(4392) := x"004f";block_ram_array(4394) := x"c9dd";block_ram_array(4396) := x"0073";block_ram_array(4398) := x"69b0";block_ram_array(4400) := x"005d";block_ram_array(4402) := x"bd21";block_ram_array(4404) := x"0036";block_ram_array(4406) := x"90ff";block_ram_array(4408) := x"00c1";block_ram_array(4410) := x"f3de";block_ram_array(4412) := x"0056";block_ram_array(4414) := x"048c";block_ram_array(4416) := x"00e0";block_ram_array(4418) := x"df14";block_ram_array(4420) := x"ff54";block_ram_array(4422) := x"e7bf";block_ram_array(4424) := x"0003";block_ram_array(4426) := x"e515";block_ram_array(4428) := x"ff06";block_ram_array(4430) := x"a0e4";block_ram_array(4432) := x"ff43";block_ram_array(4434) := x"33f4";block_ram_array(4436) := x"ff77";block_ram_array(4438) := x"46e6";block_ram_array(4440) := x"ffa1";block_ram_array(4442) := x"d478";block_ram_array(4444) := x"005a";block_ram_array(4446) := x"b99b";block_ram_array(4448) := x"001f";block_ram_array(4450) := x"9068";block_ram_array(4452) := x"ffd4";block_ram_array(4454) := x"ef58";block_ram_array(4456) := x"ff95";block_ram_array(4458) := x"b524";block_ram_array(4460) := x"ff9c";block_ram_array(4462) := x"04c9";block_ram_array(4464) := x"feef";block_ram_array(4466) := x"c510";block_ram_array(4468) := x"0028";block_ram_array(4470) := x"2ddd";block_ram_array(4472) := x"ffb9";block_ram_array(4474) := x"cf11";block_ram_array(4476) := x"0173";block_ram_array(4478) := x"f518";block_ram_array(4480) := x"0100";block_ram_array(4482) := x"503e";block_ram_array(4484) := x"0079";block_ram_array(4486) := x"be69";block_ram_array(4488) := x"0054";block_ram_array(4490) := x"cbf8";block_ram_array(4492) := x"fff2";block_ram_array(4494) := x"622c";block_ram_array(4496) := x"0071";block_ram_array(4498) := x"42ef";block_ram_array(4500) := x"0008";block_ram_array(4502) := x"8f4b";block_ram_array(4504) := x"006f";block_ram_array(4506) := x"8f80";block_ram_array(4508) := x"0000";block_ram_array(4510) := x"9ee6";block_ram_array(4512) := x"00e6";block_ram_array(4514) := x"d429";block_ram_array(4516) := x"ff4b";block_ram_array(4518) := x"dc38";block_ram_array(4520) := x"ff52";block_ram_array(4522) := x"e40a";block_ram_array(4524) := x"fea1";block_ram_array(4526) := x"89ec";block_ram_array(4528) := x"fefb";block_ram_array(4530) := x"73c4";block_ram_array(4532) := x"004c";block_ram_array(4534) := x"8bf7";block_ram_array(4536) := x"ffc6";block_ram_array(4538) := x"4ea0";block_ram_array(4540) := x"0041";block_ram_array(4542) := x"0582";block_ram_array(4544) := x"ffd0";block_ram_array(4546) := x"3266";block_ram_array(4548) := x"0080";block_ram_array(4550) := x"141e";block_ram_array(4552) := x"0050";block_ram_array(4554) := x"1b12";block_ram_array(4556) := x"ffef";block_ram_array(4558) := x"622c";block_ram_array(4560) := x"ff49";block_ram_array(4562) := x"6abd";block_ram_array(4564) := x"0012";block_ram_array(4566) := x"95a8";block_ram_array(4568) := x"002f";block_ram_array(4570) := x"6756";block_ram_array(4572) := x"0124";block_ram_array(4574) := x"1d3a";block_ram_array(4576) := x"0103";block_ram_array(4578) := x"4468";block_ram_array(4580) := x"000e";block_ram_array(4582) := x"2401";block_ram_array(4584) := x"0039";block_ram_array(4586) := x"8079";block_ram_array(4588) := x"ff80";block_ram_array(4590) := x"
2ad2";block_ram_array(4592) := x"fffe";block_ram_array(4594) := x"b506";block_ram_array(4596) := x"0003";block_ram_array(4598) := x"a651";block_ram_array(4600) := x"0070";block_ram_array(4602) := x"29d7";block_ram_array(4604) := x"ffdb";block_ram_array(4606) := x"18c6";block_ram_array(4608) := x"0032";block_ram_array(4610) := x"c32f";block_ram_array(4612) := x"ff68";block_ram_array(4614) := x"b76c";block_ram_array(4616) := x"ff9a";block_ram_array(4618) := x"00ed";block_ram_array(4620) := x"ff1e";block_ram_array(4622) := x"4b71";block_ram_array(4624) := x"fea3";block_ram_array(4626) := x"9e48";block_ram_array(4628) := x"0028";block_ram_array(4630) := x"db4d";block_ram_array(4632) := x"0008";block_ram_array(4634) := x"d7b2";block_ram_array(4636) := x"0115";block_ram_array(4638) := x"4844";block_ram_array(4640) := x"0033";block_ram_array(4642) := x"fe3a";block_ram_array(4644) := x"0018";block_ram_array(4646) := x"17a3";block_ram_array(4648) := x"003c";block_ram_array(4650) := x"f6dc";block_ram_array(4652) := x"0066";block_ram_array(4654) := x"9376";block_ram_array(4656) := x"0021";block_ram_array(4658) := x"e1c3";block_ram_array(4660) := x"ffd3";block_ram_array(4662) := x"56c0";block_ram_array(4664) := x"0022";block_ram_array(4666) := x"6c5e";block_ram_array(4668) := x"0091";block_ram_array(4670) := x"7c20";block_ram_array(4672) := x"00d8";block_ram_array(4674) := x"ce02";block_ram_array(4676) := x"ffad";block_ram_array(4678) := x"dbc8";block_ram_array(4680) := x"ffe5";block_ram_array(4682) := x"e417";block_ram_array(4684) := x"ff72";block_ram_array(4686) := x"8ad8";block_ram_array(4688) := x"ffbf";block_ram_array(4690) := x"a973";block_ram_array(4692) := x"ffc6";block_ram_array(4694) := x"7911";block_ram_array(4696) := x"ffdd";block_ram_array(4698) := x"e2c3";block_ram_array(4700) := x"004b";block_ram_array(4702) := x"945b";block_ram_array(4704) := x"0078";block_ram_array(4706) := x"c700";block_ram_array(4708) := x"ffa1";block_ram_array(4710) := x"ecdc";block_ram_array(4712) := x"ff4d";block_ram_array(4714) := x"b625";block_ram_array(4716) := x"ff6d";block_ram_array(4718) := x"6135";block_ram_array(4720) := x"ff4e";block_ram_array(4722) := x"d0a0";block_ram_array(4724) := x"0079";block_ram_array(4726) := x"3bf8";block_ram_array(4728) := x"fffb";block_ram_array(4730) := x"fd02";block_ram_array(4732) := x"00ca";block_ram_array(4734) := x"f1de";block_ram_array(4736) := x"008d";block_ram_array(4738) := x"8a98";block_ram_array(4740) := x"0047";block_ram_array(4742) := x"7d01";block_ram_array(4744) := x"003b";block_ram_array(4746) := x"93cf";block_ram_array(4748) := x"0008";block_ram_array(4750) := x"b0c8";block_ram_array(4752) := x"0060";block_ram_array(4754) := x"3c7c";block_ram_array(4756) := x"ffe6";block_ram_array(4758) := x"aa4b";block_ram_array(4760) := x"000e";block_ram_array(4762) := x"1ddf";block_ram_array(4764) := x"fff9";block_ram_array(4766) := x"dbe3";block_ram_array(4768) := x"00a0";block_ram_array(4770) := x"345a";block_ram_array(4772) := x"ffb2";block_ram_array(4774) := x"c48a";block_ram_array(4776) := x"ff84";block_ram_array(4778) := x"7dd5";block_ram_array(4780) := x"ff2d";block_ram_array(4782) := x"a3f0";block_ram_array(4784) := x"ff8d";block_ram_array(4786) := x"849c";block_ram_array(4788) := x"004c";block_ram_array(4790) := x"7976";block_ram_array(4792) := x"ffd7";block_ram_array(4794) := x"5c38";block_ram_array(4796) := x"0013";block_ram_array(4798) := x"7894";block_ram_array(4800) := x"0023";block_ram_array(4802) := x"b2e6";block_ram_array(4804) := x"005d";block_ram_array(4806) := x"f6d7";block_ram_array(4808) := x"000e";block_ram_array(4810) := x"a3a1";block_ram_array(4812) := x"ff86";block_ram_array(4814) := x"7dd2";block_ram_array(4816) := x"ff4a";block_ram_array(4818) := x"0035";block_ram_array(4820) := x"005e";block_ram_array(4822) := x"c393";block_ram_array(4824) := x"0062";block_ram_array(4826) := x"12d1";block_ram_array(4828) := x"00b5";block_ram_array(4830) := x"586c";block_ram_array(4832) := x"0081";block_ram_array(4834) := x"7aca";block_ram_array(4836) := x"fff7";block_ram_array(4838) := x"
8485";block_ram_array(4840) := x"0030";block_ram_array(4842) := x"b22a";block_ram_array(4844) := x"ffd8";block_ram_array(4846) := x"237c";block_ram_array(4848) := x"0032";block_ram_array(4850) := x"7ced";block_ram_array(4852) := x"fff0";block_ram_array(4854) := x"51d0";block_ram_array(4856) := x"002f";block_ram_array(4858) := x"384f";block_ram_array(4860) := x"ffb8";block_ram_array(4862) := x"7a6b";block_ram_array(4864) := x"000b";block_ram_array(4866) := x"fc16";block_ram_array(4868) := x"ffb5";block_ram_array(4870) := x"5e60";block_ram_array(4872) := x"ffbd";block_ram_array(4874) := x"03fa";block_ram_array(4876) := x"ff75";block_ram_array(4878) := x"2258";block_ram_array(4880) := x"ff39";block_ram_array(4882) := x"25fc";block_ram_array(4884) := x"0028";block_ram_array(4886) := x"769e";block_ram_array(4888) := x"fff7";block_ram_array(4890) := x"6fd6";block_ram_array(4892) := x"0091";block_ram_array(4894) := x"766a";block_ram_array(4896) := x"002b";block_ram_array(4898) := x"4924";block_ram_array(4900) := x"003c";block_ram_array(4902) := x"0bf8";block_ram_array(4904) := x"003c";block_ram_array(4906) := x"24ff";block_ram_array(4908) := x"0002";block_ram_array(4910) := x"22d4";block_ram_array(4912) := x"ffd1";block_ram_array(4914) := x"919e";block_ram_array(4916) := x"0003";block_ram_array(4918) := x"c80c";block_ram_array(4920) := x"0041";block_ram_array(4922) := x"559c";block_ram_array(4924) := x"007c";block_ram_array(4926) := x"6c02";block_ram_array(4928) := x"008c";block_ram_array(4930) := x"7840";block_ram_array(4932) := x"ffc6";block_ram_array(4934) := x"c365";block_ram_array(4936) := x"0003";block_ram_array(4938) := x"1ba6";block_ram_array(4940) := x"ffb4";block_ram_array(4942) := x"224e";block_ram_array(4944) := x"0002";block_ram_array(4946) := x"23fc";block_ram_array(4948) := x"ffd9";block_ram_array(4950) := x"012d";block_ram_array(4952) := x"fffb";block_ram_array(4954) := x"9baf";block_ram_array(4956) := x"ffeb";block_ram_array(4958) := x"5fc4";block_ram_array(4960) := x"001a";block_ram_array(4962) := x"ed28";block_ram_array(4964) := x"ffb6";block_ram_array(4966) := x"9a8f";block_ram_array(4968) := x"ff85";block_ram_array(4970) := x"a2f6";block_ram_array(4972) := x"ffa4";block_ram_array(4974) := x"5369";block_ram_array(4976) := x"ff82";block_ram_array(4978) := x"b076";block_ram_array(4980) := x"0055";block_ram_array(4982) := x"bce0";block_ram_array(4984) := x"ffe9";block_ram_array(4986) := x"4907";block_ram_array(4988) := x"006d";block_ram_array(4990) := x"5aa8";block_ram_array(4992) := x"0035";block_ram_array(4994) := x"f717";block_ram_array(4996) := x"0073";block_ram_array(4998) := x"5b64";block_ram_array(5000) := x"006e";block_ram_array(5002) := x"ccbc";block_ram_array(5004) := x"0003";block_ram_array(5006) := x"9ea0";block_ram_array(5008) := x"000c";block_ram_array(5010) := x"8873";block_ram_array(5012) := x"ffe8";block_ram_array(5014) := x"1b44";block_ram_array(5016) := x"0036";block_ram_array(5018) := x"5327";block_ram_array(5020) := x"002d";block_ram_array(5022) := x"deae";block_ram_array(5024) := x"0079";block_ram_array(5026) := x"e8f4";block_ram_array(5028) := x"ffbd";block_ram_array(5030) := x"95f0";block_ram_array(5032) := x"ffdb";block_ram_array(5034) := x"676e";block_ram_array(5036) := x"ff79";block_ram_array(5038) := x"4273";block_ram_array(5040) := x"ffc2";block_ram_array(5042) := x"b007";block_ram_array(5044) := x"0008";block_ram_array(5046) := x"abdb";block_ram_array(5048) := x"fff9";block_ram_array(5050) := x"dc0c";block_ram_array(5052) := x"ffe5";block_ram_array(5054) := x"ea04";block_ram_array(5056) := x"ffe0";block_ram_array(5058) := x"d2a8";block_ram_array(5060) := x"0003";block_ram_array(5062) := x"91d6";block_ram_array(5064) := x"ffe3";block_ram_array(5066) := x"d6ee";block_ram_array(5068) := x"ffc6";block_ram_array(5070) := x"3bb0";block_ram_array(5072) := x"ff6b";block_ram_array(5074) := x"ae38";block_ram_array(5076) := x"003f";block_ram_array(5078) := x"b617";block_ram_array(5080) := x"0028";block_ram_array(5082) := x"fd7e";block_ram_array(5084) := x"008f";block_ram_array(5086) := x"
4d22";block_ram_array(5088) := x"002f";block_ram_array(5090) := x"086f";block_ram_array(5092) := x"002d";block_ram_array(5094) := x"e36e";block_ram_array(5096) := x"0068";block_ram_array(5098) := x"fd9b";block_ram_array(5100) := x"002e";block_ram_array(5102) := x"2472";block_ram_array(5104) := x"003c";block_ram_array(5106) := x"1907";block_ram_array(5108) := x"ffc5";block_ram_array(5110) := x"f3e9";block_ram_array(5112) := x"002b";block_ram_array(5114) := x"cd2e";block_ram_array(5116) := x"fffb";block_ram_array(5118) := x"ff42";block_ram_array(5120) := x"0042";block_ram_array(5122) := x"e100";block_ram_array(5124) := x"ffad";block_ram_array(5126) := x"bf00";block_ram_array(5128) := x"ffe4";block_ram_array(5130) := x"c8ad";block_ram_array(5132) := x"ff8e";block_ram_array(5134) := x"9cd0";block_ram_array(5136) := x"ff8a";block_ram_array(5138) := x"ec55";block_ram_array(5140) := x"ffd9";block_ram_array(5142) := x"7ad9";block_ram_array(5144) := x"ffd6";block_ram_array(5146) := x"1afb";block_ram_array(5148) := x"0046";block_ram_array(5150) := x"2b7b";block_ram_array(5152) := x"0003";block_ram_array(5154) := x"7205";block_ram_array(5156) := x"ffff";block_ram_array(5158) := x"34c7";block_ram_array(5160) := x"ffdc";block_ram_array(5162) := x"c777";block_ram_array(5164) := x"000b";block_ram_array(5166) := x"db9c";block_ram_array(5168) := x"ffcb";block_ram_array(5170) := x"0a45";block_ram_array(5172) := x"0027";block_ram_array(5174) := x"4756";block_ram_array(5176) := x"0012";block_ram_array(5178) := x"ca49";block_ram_array(5180) := x"0078";block_ram_array(5182) := x"4844";block_ram_array(5184) := x"0059";block_ram_array(5186) := x"a723";block_ram_array(5188) := x"0013";block_ram_array(5190) := x"45ee";block_ram_array(5192) := x"0037";block_ram_array(5194) := x"ef91";block_ram_array(5196) := x"0015";block_ram_array(5198) := x"7bb8";block_ram_array(5200) := x"0057";block_ram_array(5202) := x"f2bf";block_ram_array(5204) := x"ffca";block_ram_array(5206) := x"7a4e";block_ram_array(5208) := x"0002";block_ram_array(5210) := x"8b5c";block_ram_array(5212) := x"ffdb";block_ram_array(5214) := x"70bf";block_ram_array(5216) := x"0044";block_ram_array(5218) := x"fb95";block_ram_array(5220) := x"ffbd";block_ram_array(5222) := x"5852";block_ram_array(5224) := x"ffb9";block_ram_array(5226) := x"a92c";block_ram_array(5228) := x"ff84";block_ram_array(5230) := x"80bc";block_ram_array(5232) := x"ff9b";block_ram_array(5234) := x"eb6a";block_ram_array(5236) := x"0001";block_ram_array(5238) := x"6260";block_ram_array(5240) := x"ffb5";block_ram_array(5242) := x"7b05";block_ram_array(5244) := x"002b";block_ram_array(5246) := x"6702";block_ram_array(5248) := x"fffe";block_ram_array(5250) := x"8164";block_ram_array(5252) := x"0052";block_ram_array(5254) := x"d949";block_ram_array(5256) := x"0015";block_ram_array(5258) := x"d013";block_ram_array(5260) := x"000a";block_ram_array(5262) := x"69ff";block_ram_array(5264) := x"ffe5";block_ram_array(5266) := x"01de";block_ram_array(5268) := x"0027";block_ram_array(5270) := x"37ca";block_ram_array(5272) := x"0029";block_ram_array(5274) := x"848f";block_ram_array(5276) := x"0055";block_ram_array(5278) := x"1c0c";block_ram_array(5280) := x"0063";block_ram_array(5282) := x"d620";block_ram_array(5284) := x"0000";block_ram_array(5286) := x"816b";block_ram_array(5288) := x"001c";block_ram_array(5290) := x"4dae";block_ram_array(5292) := x"ffdb";block_ram_array(5294) := x"4dd3";block_ram_array(5296) := x"0033";block_ram_array(5298) := x"10fb";block_ram_array(5300) := x"fff2";block_ram_array(5302) := x"b9a8";block_ram_array(5304) := x"0014";block_ram_array(5306) := x"08c1";block_ram_array(5308) := x"ffb7";block_ram_array(5310) := x"956e";block_ram_array(5312) := x"fffd";block_ram_array(5314) := x"dfd4";block_ram_array(5316) := x"ffdc";block_ram_array(5318) := x"d555";block_ram_array(5320) := x"ffeb";block_ram_array(5322) := x"c7c3";block_ram_array(5324) := x"ffa2";block_ram_array(5326) := x"6c28";block_ram_array(5328) := x"ff7e";block_ram_array(5330) := x"5574";block_ram_array(5332) := x"ffef";block_ram_array(5334) := x"
f7de";block_ram_array(5336) := x"ffc8";block_ram_array(5338) := x"e1b1";block_ram_array(5340) := x"0050";block_ram_array(5342) := x"0439";block_ram_array(5344) := x"fff8";block_ram_array(5346) := x"2f87";block_ram_array(5348) := x"0045";block_ram_array(5350) := x"57dd";block_ram_array(5352) := x"0027";block_ram_array(5354) := x"5b53";block_ram_array(5356) := x"0037";block_ram_array(5358) := x"860a";block_ram_array(5360) := x"0015";block_ram_array(5362) := x"690f";block_ram_array(5364) := x"000e";block_ram_array(5366) := x"fb4a";block_ram_array(5368) := x"002b";block_ram_array(5370) := x"71d9";block_ram_array(5372) := x"0039";block_ram_array(5374) := x"49b9";block_ram_array(5376) := x"0062";block_ram_array(5378) := x"30d1";block_ram_array(5380) := x"ffeb";block_ram_array(5382) := x"049a";block_ram_array(5384) := x"0015";block_ram_array(5386) := x"4d34";block_ram_array(5388) := x"ffc1";block_ram_array(5390) := x"aedb";block_ram_array(5392) := x"0004";block_ram_array(5394) := x"cff8";block_ram_array(5396) := x"ffde";block_ram_array(5398) := x"4fb7";block_ram_array(5400) := x"fffc";block_ram_array(5402) := x"8893";block_ram_array(5404) := x"ffe0";block_ram_array(5406) := x"7c8f";block_ram_array(5408) := x"0000";block_ram_array(5410) := x"ff93";block_ram_array(5412) := x"ffdb";block_ram_array(5414) := x"7c1c";block_ram_array(5416) := x"ffd4";block_ram_array(5418) := x"db8f";block_ram_array(5420) := x"ffca";block_ram_array(5422) := x"8c28";block_ram_array(5424) := x"ffb0";block_ram_array(5426) := x"bfaf";block_ram_array(5428) := x"0001";block_ram_array(5430) := x"b7b3";block_ram_array(5432) := x"ffc6";block_ram_array(5434) := x"5c5e";block_ram_array(5436) := x"0039";block_ram_array(5438) := x"f1d2";block_ram_array(5440) := x"ffff";block_ram_array(5442) := x"ab1e";block_ram_array(5444) := x"0051";block_ram_array(5446) := x"1478";block_ram_array(5448) := x"002c";block_ram_array(5450) := x"e132";block_ram_array(5452) := x"0036";block_ram_array(5454) := x"62ba";block_ram_array(5456) := x"0033";block_ram_array(5458) := x"2963";block_ram_array(5460) := x"000d";block_ram_array(5462) := x"0825";block_ram_array(5464) := x"0023";block_ram_array(5466) := x"283b";block_ram_array(5468) := x"0014";block_ram_array(5470) := x"9cce";block_ram_array(5472) := x"0064";block_ram_array(5474) := x"1184";block_ram_array(5476) := x"fff2";block_ram_array(5478) := x"be78";block_ram_array(5480) := x"000b";block_ram_array(5482) := x"fc2d";block_ram_array(5484) := x"ff93";block_ram_array(5486) := x"add2";block_ram_array(5488) := x"ffda";block_ram_array(5490) := x"562b";block_ram_array(5492) := x"fff1";block_ram_array(5494) := x"a89a";block_ram_array(5496) := x"fff8";block_ram_array(5498) := x"e77d";block_ram_array(5500) := x"ffdb";block_ram_array(5502) := x"cd9e";block_ram_array(5504) := x"ffd9";block_ram_array(5506) := x"6017";block_ram_array(5508) := x"0003";block_ram_array(5510) := x"a43b";block_ram_array(5512) := x"fffd";block_ram_array(5514) := x"e5d5";block_ram_array(5516) := x"ffe7";block_ram_array(5518) := x"f743";block_ram_array(5520) := x"ffb1";block_ram_array(5522) := x"7d6f";block_ram_array(5524) := x"0004";block_ram_array(5526) := x"e9fb";block_ram_array(5528) := x"fff0";block_ram_array(5530) := x"99e7";block_ram_array(5532) := x"0043";block_ram_array(5534) := x"0f31";block_ram_array(5536) := x"0003";block_ram_array(5538) := x"490f";block_ram_array(5540) := x"002e";block_ram_array(5542) := x"df50";block_ram_array(5544) := x"0029";block_ram_array(5546) := x"7325";block_ram_array(5548) := x"0033";block_ram_array(5550) := x"1c4e";block_ram_array(5552) := x"0033";block_ram_array(5554) := x"6718";block_ram_array(5556) := x"000b";block_ram_array(5558) := x"766e";block_ram_array(5560) := x"0032";block_ram_array(5562) := x"9c34";block_ram_array(5564) := x"fffc";block_ram_array(5566) := x"0434";block_ram_array(5568) := x"0035";block_ram_array(5570) := x"7406";block_ram_array(5572) := x"ffe9";block_ram_array(5574) := x"c2d7";block_ram_array(5576) := x"0028";block_ram_array(5578) := x"a987";block_ram_array(5580) := x"ffaa";block_ram_array(5582) := x"
797c";block_ram_array(5584) := x"ffb6";block_ram_array(5586) := x"c5bb";block_ram_array(5588) := x"ffc0";block_ram_array(5590) := x"1fd8";block_ram_array(5592) := x"ffe0";block_ram_array(5594) := x"8dbf";block_ram_array(5596) := x"0016";block_ram_array(5598) := x"3cad";block_ram_array(5600) := x"ffe4";block_ram_array(5602) := x"86d6";block_ram_array(5604) := x"fff8";block_ram_array(5606) := x"20c2";block_ram_array(5608) := x"ffee";block_ram_array(5610) := x"e6c6";block_ram_array(5612) := x"0019";block_ram_array(5614) := x"babd";block_ram_array(5616) := x"ffe4";block_ram_array(5618) := x"3864";block_ram_array(5620) := x"0005";block_ram_array(5622) := x"6887";block_ram_array(5624) := x"fff8";block_ram_array(5626) := x"277f";block_ram_array(5628) := x"0043";block_ram_array(5630) := x"20df";block_ram_array(5632) := x"0024";block_ram_array(5634) := x"64d0";block_ram_array(5636) := x"0011";block_ram_array(5638) := x"d56c";block_ram_array(5640) := x"0012";block_ram_array(5642) := x"dfc5";block_ram_array(5644) := x"0020";block_ram_array(5646) := x"9999";block_ram_array(5648) := x"0039";block_ram_array(5650) := x"21dd";block_ram_array(5652) := x"fffd";block_ram_array(5654) := x"d692";block_ram_array(5656) := x"0014";block_ram_array(5658) := x"d91f";block_ram_array(5660) := x"fff6";block_ram_array(5662) := x"547e";block_ram_array(5664) := x"0036";block_ram_array(5666) := x"ef87";block_ram_array(5668) := x"ffeb";block_ram_array(5670) := x"3a68";block_ram_array(5672) := x"000b";block_ram_array(5674) := x"e18c";block_ram_array(5676) := x"ffb3";block_ram_array(5678) := x"4bf6";block_ram_array(5680) := x"ffcc";block_ram_array(5682) := x"c88f";block_ram_array(5684) := x"ffce";block_ram_array(5686) := x"a1fa";block_ram_array(5688) := x"ffc7";block_ram_array(5690) := x"38d2";block_ram_array(5692) := x"0008";block_ram_array(5694) := x"06f8";block_ram_array(5696) := x"ffe5";block_ram_array(5698) := x"4061";block_ram_array(5700) := x"001c";block_ram_array(5702) := x"cf86";block_ram_array(5704) := x"fff8";block_ram_array(5706) := x"3fff";block_ram_array(5708) := x"0020";block_ram_array(5710) := x"0ffa";block_ram_array(5712) := x"fffd";block_ram_array(5714) := x"4191";block_ram_array(5716) := x"0015";block_ram_array(5718) := x"1fc9";block_ram_array(5720) := x"0004";block_ram_array(5722) := x"51bc";block_ram_array(5724) := x"0034";block_ram_array(5726) := x"2ccb";block_ram_array(5728) := x"0041";block_ram_array(5730) := x"a047";block_ram_array(5732) := x"0011";block_ram_array(5734) := x"5137";block_ram_array(5736) := x"000d";block_ram_array(5738) := x"23c3";block_ram_array(5740) := x"ffe5";block_ram_array(5742) := x"77c3";block_ram_array(5744) := x"0016";block_ram_array(5746) := x"d0bb";block_ram_array(5748) := x"000e";block_ram_array(5750) := x"ab7a";block_ram_array(5752) := x"001e";block_ram_array(5754) := x"c5ce";block_ram_array(5756) := x"ffdf";block_ram_array(5758) := x"965d";block_ram_array(5760) := x"0000";block_ram_array(5762) := x"c116";block_ram_array(5764) := x"fff5";block_ram_array(5766) := x"6d94";block_ram_array(5768) := x"001d";block_ram_array(5770) := x"6fb2";block_ram_array(5772) := x"ffd7";block_ram_array(5774) := x"0380";block_ram_array(5776) := x"ffca";block_ram_array(5778) := x"3e28";block_ram_array(5780) := x"ffc9";block_ram_array(5782) := x"83b2";block_ram_array(5784) := x"ffce";block_ram_array(5786) := x"2c3e";block_ram_array(5788) := x"001b";block_ram_array(5790) := x"69b7";block_ram_array(5792) := x"ffec";block_ram_array(5794) := x"3730";block_ram_array(5796) := x"0018";block_ram_array(5798) := x"b33a";block_ram_array(5800) := x"fffa";block_ram_array(5802) := x"6911";block_ram_array(5804) := x"002c";block_ram_array(5806) := x"6c7d";block_ram_array(5808) := x"000f";block_ram_array(5810) := x"e48f";block_ram_array(5812) := x"0019";block_ram_array(5814) := x"575b";block_ram_array(5816) := x"0014";block_ram_array(5818) := x"432b";block_ram_array(5820) := x"0028";block_ram_array(5822) := x"d40b";block_ram_array(5824) := x"0042";block_ram_array(5826) := x"f603";block_ram_array(5828) := x"0006";block_ram_array(5830) := x"
a5f1";block_ram_array(5832) := x"001c";block_ram_array(5834) := x"db74";block_ram_array(5836) := x"ffd5";block_ram_array(5838) := x"d00e";block_ram_array(5840) := x"fffa";block_ram_array(5842) := x"eab4";block_ram_array(5844) := x"ffe8";block_ram_array(5846) := x"cecd";block_ram_array(5848) := x"0001";block_ram_array(5850) := x"aa74";block_ram_array(5852) := x"fff9";block_ram_array(5854) := x"e931";block_ram_array(5856) := x"0002";block_ram_array(5858) := x"dfd3";block_ram_array(5860) := x"ffef";block_ram_array(5862) := x"6de4";block_ram_array(5864) := x"fff9";block_ram_array(5866) := x"57c6";block_ram_array(5868) := x"fff5";block_ram_array(5870) := x"9531";block_ram_array(5872) := x"fff2";block_ram_array(5874) := x"6e45";block_ram_array(5876) := x"ffef";block_ram_array(5878) := x"d017";block_ram_array(5880) := x"ffe1";block_ram_array(5882) := x"d8c2";block_ram_array(5884) := x"000e";block_ram_array(5886) := x"0cf7";block_ram_array(5888) := x"0003";block_ram_array(5890) := x"a4cd";block_ram_array(5892) := x"0017";block_ram_array(5894) := x"94ee";block_ram_array(5896) := x"0003";block_ram_array(5898) := x"37d6";block_ram_array(5900) := x"000e";block_ram_array(5902) := x"1d12";block_ram_array(5904) := x"0010";block_ram_array(5906) := x"d686";block_ram_array(5908) := x"000b";block_ram_array(5910) := x"6b42";block_ram_array(5912) := x"0007";block_ram_array(5914) := x"8f4f";block_ram_array(5916) := x"0001";block_ram_array(5918) := x"081e";block_ram_array(5920) := x"000d";block_ram_array(5922) := x"9ef2";block_ram_array(5924) := x"0005";block_ram_array(5926) := x"0b81";block_ram_array(5928) := x"0007";block_ram_array(5930) := x"34e8";block_ram_array(5932) := x"fffb";block_ram_array(5934) := x"7382";block_ram_array(5936) := x"0006";block_ram_array(5938) := x"ec66";block_ram_array(5940) := x"0001";block_ram_array(5942) := x"de6e";block_ram_array(5944) := x"0005";block_ram_array(5946) := x"7fe2";block_ram_array(5948) := x"fffe";block_ram_array(5950) := x"3119";block_ram_array(5952) := x"0006";block_ram_array(5954) := x"bd74";block_ram_array(5956) := x"0001";block_ram_array(5958) := x"6844";block_ram_array(5960) := x"0005";block_ram_array(5962) := x"0502";block_ram_array(5964) := x"fffe";block_ram_array(5966) := x"48ba";block_ram_array(5968) := x"0006";block_ram_array(5970) := x"1e34";block_ram_array(5972) := x"0001";block_ram_array(5974) := x"158b";block_ram_array(5976) := x"0004";block_ram_array(5978) := x"c7a7";block_ram_array(5980) := x"fffe";block_ram_array(5982) := x"7d27";block_ram_array(5984) := x"0005";block_ram_array(5986) := x"b7f5";block_ram_array(5988) := x"0000";block_ram_array(5990) := x"d053";block_ram_array(5992) := x"0004";block_ram_array(5994) := x"84cb";block_ram_array(5996) := x"fffe";block_ram_array(5998) := x"a117";block_ram_array(6000) := x"0005";block_ram_array(6002) := x"6df9";block_ram_array(6004) := x"0000";block_ram_array(6006) := x"d522";block_ram_array(6008) := x"0004";block_ram_array(6010) := x"aa8a";block_ram_array(6012) := x"fffe";block_ram_array(6014) := x"a522";block_ram_array(6016) := x"0004";block_ram_array(6018) := x"f8f0";block_ram_array(6020) := x"0000";block_ram_array(6022) := x"6c6f";block_ram_array(6024) := x"0004";block_ram_array(6026) := x"52ed";block_ram_array(6028) := x"fffe";block_ram_array(6030) := x"f7d8";block_ram_array(6032) := x"0004";block_ram_array(6034) := x"db0c";block_ram_array(6036) := x"0000";block_ram_array(6038) := x"88ed";block_ram_array(6040) := x"0004";block_ram_array(6042) := x"5d9d";block_ram_array(6044) := x"ffff";block_ram_array(6046) := x"201b";block_ram_array(6048) := x"0004";block_ram_array(6050) := x"d4bf";block_ram_array(6052) := x"0000";block_ram_array(6054) := x"8d90";block_ram_array(6056) := x"0004";block_ram_array(6058) := x"a6c7";block_ram_array(6060) := x"fffe";block_ram_array(6062) := x"edb4";block_ram_array(6064) := x"0004";block_ram_array(6066) := x"21ce";block_ram_array(6068) := x"0000";block_ram_array(6070) := x"09cf";block_ram_array(6072) := x"0004";block_ram_array(6074) := x"40ec";block_ram_array(6076) := x"ffff";block_ram_array(6078) := x"
b946";block_ram_array(6080) := x"0004";block_ram_array(6082) := x"7d4a";block_ram_array(6084) := x"0000";block_ram_array(6086) := x"2823";block_ram_array(6088) := x"0004";block_ram_array(6090) := x"4d49";block_ram_array(6092) := x"ffff";block_ram_array(6094) := x"cb33";block_ram_array(6096) := x"0004";block_ram_array(6098) := x"ac93";block_ram_array(6100) := x"ffff";block_ram_array(6102) := x"f6f7";block_ram_array(6104) := x"0004";block_ram_array(6106) := x"024f";block_ram_array(6108) := x"ffff";block_ram_array(6110) := x"8dc4";block_ram_array(6112) := x"0004";block_ram_array(6114) := x"43e7";block_ram_array(6116) := x"0000";block_ram_array(6118) := x"335e";block_ram_array(6120) := x"0004";block_ram_array(6122) := x"0e6a";block_ram_array(6124) := x"0000";block_ram_array(6126) := x"0432";block_ram_array(6128) := x"0004";block_ram_array(6130) := x"83a4";block_ram_array(6132) := x"0000";block_ram_array(6134) := x"743d";block_ram_array(6136) := x"0004";block_ram_array(6138) := x"937e";block_ram_array(6140) := x"0000";block_ram_array(6142) := x"03e5";block_ram_array(6144) := x"0004";block_ram_array(6146) := x"9200";block_ram_array(6148) := x"0000";block_ram_array(6150) := x"0000";block_ram_array(6152) := x"0004";block_ram_array(6154) := x"937e";block_ram_array(6156) := x"ffff";block_ram_array(6158) := x"fc1b";block_ram_array(6160) := x"0004";block_ram_array(6162) := x"83a4";block_ram_array(6164) := x"ffff";block_ram_array(6166) := x"8bc3";block_ram_array(6168) := x"0004";block_ram_array(6170) := x"0e6a";block_ram_array(6172) := x"ffff";block_ram_array(6174) := x"fbce";block_ram_array(6176) := x"0004";block_ram_array(6178) := x"43e7";block_ram_array(6180) := x"ffff";block_ram_array(6182) := x"cca2";block_ram_array(6184) := x"0004";block_ram_array(6186) := x"024f";block_ram_array(6188) := x"0000";block_ram_array(6190) := x"723c";block_ram_array(6192) := x"0004";block_ram_array(6194) := x"ac93";block_ram_array(6196) := x"0000";block_ram_array(6198) := x"0909";block_ram_array(6200) := x"0004";block_ram_array(6202) := x"4d49";block_ram_array(6204) := x"0000";block_ram_array(6206) := x"34cd";block_ram_array(6208) := x"0004";block_ram_array(6210) := x"7d4a";block_ram_array(6212) := x"ffff";block_ram_array(6214) := x"d7dd";block_ram_array(6216) := x"0004";block_ram_array(6218) := x"40ec";block_ram_array(6220) := x"0000";block_ram_array(6222) := x"46ba";block_ram_array(6224) := x"0004";block_ram_array(6226) := x"21ce";block_ram_array(6228) := x"ffff";block_ram_array(6230) := x"f631";block_ram_array(6232) := x"0004";block_ram_array(6234) := x"a6c7";block_ram_array(6236) := x"0001";block_ram_array(6238) := x"124c";block_ram_array(6240) := x"0004";block_ram_array(6242) := x"d4bf";block_ram_array(6244) := x"ffff";block_ram_array(6246) := x"7270";block_ram_array(6248) := x"0004";block_ram_array(6250) := x"5d9d";block_ram_array(6252) := x"0000";block_ram_array(6254) := x"dfe5";block_ram_array(6256) := x"0004";block_ram_array(6258) := x"db0c";block_ram_array(6260) := x"ffff";block_ram_array(6262) := x"7713";block_ram_array(6264) := x"0004";block_ram_array(6266) := x"52ed";block_ram_array(6268) := x"0001";block_ram_array(6270) := x"0828";block_ram_array(6272) := x"0004";block_ram_array(6274) := x"f8f0";block_ram_array(6276) := x"ffff";block_ram_array(6278) := x"9391";block_ram_array(6280) := x"0004";block_ram_array(6282) := x"aa8a";block_ram_array(6284) := x"0001";block_ram_array(6286) := x"5ade";block_ram_array(6288) := x"0005";block_ram_array(6290) := x"6df9";block_ram_array(6292) := x"ffff";block_ram_array(6294) := x"2ade";block_ram_array(6296) := x"0004";block_ram_array(6298) := x"84cb";block_ram_array(6300) := x"0001";block_ram_array(6302) := x"5ee9";block_ram_array(6304) := x"0005";block_ram_array(6306) := x"b7f5";block_ram_array(6308) := x"ffff";block_ram_array(6310) := x"2fad";block_ram_array(6312) := x"0004";block_ram_array(6314) := x"c7a7";block_ram_array(6316) := x"0001";block_ram_array(6318) := x"82d9";block_ram_array(6320) := x"0006";block_ram_array(6322) := x"1e34";block_ram_array(6324) := x"fffe";block_ram_array(6326) := x"
ea75";block_ram_array(6328) := x"0005";block_ram_array(6330) := x"0502";block_ram_array(6332) := x"0001";block_ram_array(6334) := x"b746";block_ram_array(6336) := x"0006";block_ram_array(6338) := x"bd74";block_ram_array(6340) := x"fffe";block_ram_array(6342) := x"97bc";block_ram_array(6344) := x"0005";block_ram_array(6346) := x"7fe2";block_ram_array(6348) := x"0001";block_ram_array(6350) := x"cee7";block_ram_array(6352) := x"0006";block_ram_array(6354) := x"ec66";block_ram_array(6356) := x"fffe";block_ram_array(6358) := x"2192";block_ram_array(6360) := x"0007";block_ram_array(6362) := x"34e8";block_ram_array(6364) := x"0004";block_ram_array(6366) := x"8c7e";block_ram_array(6368) := x"000d";block_ram_array(6370) := x"9ef2";block_ram_array(6372) := x"fffa";block_ram_array(6374) := x"f47f";block_ram_array(6376) := x"0007";block_ram_array(6378) := x"8f4f";block_ram_array(6380) := x"fffe";block_ram_array(6382) := x"f7e2";block_ram_array(6384) := x"0010";block_ram_array(6386) := x"d686";block_ram_array(6388) := x"fff4";block_ram_array(6390) := x"94be";block_ram_array(6392) := x"0003";block_ram_array(6394) := x"37d6";block_ram_array(6396) := x"fff1";block_ram_array(6398) := x"e2ee";block_ram_array(6400) := x"0003";block_ram_array(6402) := x"a4cd";block_ram_array(6404) := x"ffe8";block_ram_array(6406) := x"6b12";block_ram_array(6408) := x"ffe1";block_ram_array(6410) := x"d8c2";block_ram_array(6412) := x"fff1";block_ram_array(6414) := x"f309";block_ram_array(6416) := x"fff2";block_ram_array(6418) := x"6e45";block_ram_array(6420) := x"0010";block_ram_array(6422) := x"2fe9";block_ram_array(6424) := x"fff9";block_ram_array(6426) := x"57c6";block_ram_array(6428) := x"000a";block_ram_array(6430) := x"6acf";block_ram_array(6432) := x"0002";block_ram_array(6434) := x"dfd3";block_ram_array(6436) := x"0010";block_ram_array(6438) := x"921c";block_ram_array(6440) := x"0001";block_ram_array(6442) := x"aa74";block_ram_array(6444) := x"0006";block_ram_array(6446) := x"16cf";block_ram_array(6448) := x"fffa";block_ram_array(6450) := x"eab4";block_ram_array(6452) := x"0017";block_ram_array(6454) := x"3133";block_ram_array(6456) := x"001c";block_ram_array(6458) := x"db74";block_ram_array(6460) := x"002a";block_ram_array(6462) := x"2ff2";block_ram_array(6464) := x"0042";block_ram_array(6466) := x"f603";block_ram_array(6468) := x"fff9";block_ram_array(6470) := x"5a0f";block_ram_array(6472) := x"0014";block_ram_array(6474) := x"432b";block_ram_array(6476) := x"ffd7";block_ram_array(6478) := x"2bf5";block_ram_array(6480) := x"000f";block_ram_array(6482) := x"e48f";block_ram_array(6484) := x"ffe6";block_ram_array(6486) := x"a8a5";block_ram_array(6488) := x"fffa";block_ram_array(6490) := x"6911";block_ram_array(6492) := x"ffd3";block_ram_array(6494) := x"9383";block_ram_array(6496) := x"ffec";block_ram_array(6498) := x"3730";block_ram_array(6500) := x"ffe7";block_ram_array(6502) := x"4cc6";block_ram_array(6504) := x"ffce";block_ram_array(6506) := x"2c3e";block_ram_array(6508) := x"ffe4";block_ram_array(6510) := x"9649";block_ram_array(6512) := x"ffca";block_ram_array(6514) := x"3e28";block_ram_array(6516) := x"0036";block_ram_array(6518) := x"7c4e";block_ram_array(6520) := x"001d";block_ram_array(6522) := x"6fb2";block_ram_array(6524) := x"0028";block_ram_array(6526) := x"fc80";block_ram_array(6528) := x"0000";block_ram_array(6530) := x"c116";block_ram_array(6532) := x"000a";block_ram_array(6534) := x"926c";block_ram_array(6536) := x"001e";block_ram_array(6538) := x"c5ce";block_ram_array(6540) := x"0020";block_ram_array(6542) := x"69a3";block_ram_array(6544) := x"0016";block_ram_array(6546) := x"d0bb";block_ram_array(6548) := x"fff1";block_ram_array(6550) := x"5486";block_ram_array(6552) := x"000d";block_ram_array(6554) := x"23c3";block_ram_array(6556) := x"001a";block_ram_array(6558) := x"883d";block_ram_array(6560) := x"0041";block_ram_array(6562) := x"a047";block_ram_array(6564) := x"ffee";block_ram_array(6566) := x"aec9";block_ram_array(6568) := x"0004";block_ram_array(6570) := x"51bc";block_ram_array(6572) := x"ffcb";block_ram_array(6574) := x"
d335";block_ram_array(6576) := x"fffd";block_ram_array(6578) := x"4191";block_ram_array(6580) := x"ffea";block_ram_array(6582) := x"e037";block_ram_array(6584) := x"fff8";block_ram_array(6586) := x"3fff";block_ram_array(6588) := x"ffdf";block_ram_array(6590) := x"f006";block_ram_array(6592) := x"ffe5";block_ram_array(6594) := x"4061";block_ram_array(6596) := x"ffe3";block_ram_array(6598) := x"307a";block_ram_array(6600) := x"ffc7";block_ram_array(6602) := x"38d2";block_ram_array(6604) := x"fff7";block_ram_array(6606) := x"f908";block_ram_array(6608) := x"ffcc";block_ram_array(6610) := x"c88f";block_ram_array(6612) := x"0031";block_ram_array(6614) := x"5e06";block_ram_array(6616) := x"000b";block_ram_array(6618) := x"e18c";block_ram_array(6620) := x"004c";block_ram_array(6622) := x"b40a";block_ram_array(6624) := x"0036";block_ram_array(6626) := x"ef87";block_ram_array(6628) := x"0014";block_ram_array(6630) := x"c598";block_ram_array(6632) := x"0014";block_ram_array(6634) := x"d91f";block_ram_array(6636) := x"0009";block_ram_array(6638) := x"ab82";block_ram_array(6640) := x"0039";block_ram_array(6642) := x"21dd";block_ram_array(6644) := x"0002";block_ram_array(6646) := x"296e";block_ram_array(6648) := x"0012";block_ram_array(6650) := x"dfc5";block_ram_array(6652) := x"ffdf";block_ram_array(6654) := x"6667";block_ram_array(6656) := x"0024";block_ram_array(6658) := x"64d0";block_ram_array(6660) := x"ffee";block_ram_array(6662) := x"2a94";block_ram_array(6664) := x"fff8";block_ram_array(6666) := x"277f";block_ram_array(6668) := x"ffbc";block_ram_array(6670) := x"df21";block_ram_array(6672) := x"ffe4";block_ram_array(6674) := x"3864";block_ram_array(6676) := x"fffa";block_ram_array(6678) := x"9779";block_ram_array(6680) := x"ffee";block_ram_array(6682) := x"e6c6";block_ram_array(6684) := x"ffe6";block_ram_array(6686) := x"4543";block_ram_array(6688) := x"ffe4";block_ram_array(6690) := x"86d6";block_ram_array(6692) := x"0007";block_ram_array(6694) := x"df3e";block_ram_array(6696) := x"ffe0";block_ram_array(6698) := x"8dbf";block_ram_array(6700) := x"ffe9";block_ram_array(6702) := x"c353";block_ram_array(6704) := x"ffb6";block_ram_array(6706) := x"c5bb";block_ram_array(6708) := x"003f";block_ram_array(6710) := x"e028";block_ram_array(6712) := x"0028";block_ram_array(6714) := x"a987";block_ram_array(6716) := x"0055";block_ram_array(6718) := x"8684";block_ram_array(6720) := x"0035";block_ram_array(6722) := x"7406";block_ram_array(6724) := x"0016";block_ram_array(6726) := x"3d29";block_ram_array(6728) := x"0032";block_ram_array(6730) := x"9c34";block_ram_array(6732) := x"0003";block_ram_array(6734) := x"fbcc";block_ram_array(6736) := x"0033";block_ram_array(6738) := x"6718";block_ram_array(6740) := x"fff4";block_ram_array(6742) := x"8992";block_ram_array(6744) := x"0029";block_ram_array(6746) := x"7325";block_ram_array(6748) := x"ffcc";block_ram_array(6750) := x"e3b2";block_ram_array(6752) := x"0003";block_ram_array(6754) := x"490f";block_ram_array(6756) := x"ffd1";block_ram_array(6758) := x"20b0";block_ram_array(6760) := x"fff0";block_ram_array(6762) := x"99e7";block_ram_array(6764) := x"ffbc";block_ram_array(6766) := x"f0cf";block_ram_array(6768) := x"ffb1";block_ram_array(6770) := x"7d6f";block_ram_array(6772) := x"fffb";block_ram_array(6774) := x"1605";block_ram_array(6776) := x"fffd";block_ram_array(6778) := x"e5d5";block_ram_array(6780) := x"0018";block_ram_array(6782) := x"08bd";block_ram_array(6784) := x"ffd9";block_ram_array(6786) := x"6017";block_ram_array(6788) := x"fffc";block_ram_array(6790) := x"5bc5";block_ram_array(6792) := x"fff8";block_ram_array(6794) := x"e77d";block_ram_array(6796) := x"0024";block_ram_array(6798) := x"3262";block_ram_array(6800) := x"ffda";block_ram_array(6802) := x"562b";block_ram_array(6804) := x"000e";block_ram_array(6806) := x"5766";block_ram_array(6808) := x"000b";block_ram_array(6810) := x"fc2d";block_ram_array(6812) := x"006c";block_ram_array(6814) := x"522e";block_ram_array(6816) := x"0064";block_ram_array(6818) := x"1184";block_ram_array(6820) := x"000d";block_ram_array(6822) := x"
4188";block_ram_array(6824) := x"0023";block_ram_array(6826) := x"283b";block_ram_array(6828) := x"ffeb";block_ram_array(6830) := x"6332";block_ram_array(6832) := x"0033";block_ram_array(6834) := x"2963";block_ram_array(6836) := x"fff2";block_ram_array(6838) := x"f7db";block_ram_array(6840) := x"002c";block_ram_array(6842) := x"e132";block_ram_array(6844) := x"ffc9";block_ram_array(6846) := x"9d46";block_ram_array(6848) := x"ffff";block_ram_array(6850) := x"ab1e";block_ram_array(6852) := x"ffae";block_ram_array(6854) := x"eb88";block_ram_array(6856) := x"ffc6";block_ram_array(6858) := x"5c5e";block_ram_array(6860) := x"ffc6";block_ram_array(6862) := x"0e2e";block_ram_array(6864) := x"ffb0";block_ram_array(6866) := x"bfaf";block_ram_array(6868) := x"fffe";block_ram_array(6870) := x"484d";block_ram_array(6872) := x"ffd4";block_ram_array(6874) := x"db8f";block_ram_array(6876) := x"0035";block_ram_array(6878) := x"73d8";block_ram_array(6880) := x"0000";block_ram_array(6882) := x"ff93";block_ram_array(6884) := x"0024";block_ram_array(6886) := x"83e4";block_ram_array(6888) := x"fffc";block_ram_array(6890) := x"8893";block_ram_array(6892) := x"001f";block_ram_array(6894) := x"8371";block_ram_array(6896) := x"0004";block_ram_array(6898) := x"cff8";block_ram_array(6900) := x"0021";block_ram_array(6902) := x"b049";block_ram_array(6904) := x"0015";block_ram_array(6906) := x"4d34";block_ram_array(6908) := x"003e";block_ram_array(6910) := x"5125";block_ram_array(6912) := x"0062";block_ram_array(6914) := x"30d1";block_ram_array(6916) := x"0014";block_ram_array(6918) := x"fb66";block_ram_array(6920) := x"002b";block_ram_array(6922) := x"71d9";block_ram_array(6924) := x"ffc6";block_ram_array(6926) := x"b647";block_ram_array(6928) := x"0015";block_ram_array(6930) := x"690f";block_ram_array(6932) := x"fff1";block_ram_array(6934) := x"04b6";block_ram_array(6936) := x"0027";block_ram_array(6938) := x"5b53";block_ram_array(6940) := x"ffc8";block_ram_array(6942) := x"79f6";block_ram_array(6944) := x"fff8";block_ram_array(6946) := x"2f87";block_ram_array(6948) := x"ffba";block_ram_array(6950) := x"a823";block_ram_array(6952) := x"ffc8";block_ram_array(6954) := x"e1b1";block_ram_array(6956) := x"ffaf";block_ram_array(6958) := x"fbc7";block_ram_array(6960) := x"ff7e";block_ram_array(6962) := x"5574";block_ram_array(6964) := x"0010";block_ram_array(6966) := x"0822";block_ram_array(6968) := x"ffeb";block_ram_array(6970) := x"c7c3";block_ram_array(6972) := x"005d";block_ram_array(6974) := x"93d8";block_ram_array(6976) := x"fffd";block_ram_array(6978) := x"dfd4";block_ram_array(6980) := x"0023";block_ram_array(6982) := x"2aab";block_ram_array(6984) := x"0014";block_ram_array(6986) := x"08c1";block_ram_array(6988) := x"0048";block_ram_array(6990) := x"6a92";block_ram_array(6992) := x"0033";block_ram_array(6994) := x"10fb";block_ram_array(6996) := x"000d";block_ram_array(6998) := x"4658";block_ram_array(7000) := x"001c";block_ram_array(7002) := x"4dae";block_ram_array(7004) := x"0024";block_ram_array(7006) := x"b22d";block_ram_array(7008) := x"0063";block_ram_array(7010) := x"d620";block_ram_array(7012) := x"ffff";block_ram_array(7014) := x"7e95";block_ram_array(7016) := x"0029";block_ram_array(7018) := x"848f";block_ram_array(7020) := x"ffaa";block_ram_array(7022) := x"e3f4";block_ram_array(7024) := x"ffe5";block_ram_array(7026) := x"01de";block_ram_array(7028) := x"ffd8";block_ram_array(7030) := x"c836";block_ram_array(7032) := x"0015";block_ram_array(7034) := x"d013";block_ram_array(7036) := x"fff5";block_ram_array(7038) := x"9601";block_ram_array(7040) := x"fffe";block_ram_array(7042) := x"8164";block_ram_array(7044) := x"ffad";block_ram_array(7046) := x"26b7";block_ram_array(7048) := x"ffb5";block_ram_array(7050) := x"7b05";block_ram_array(7052) := x"ffd4";block_ram_array(7054) := x"98fe";block_ram_array(7056) := x"ff9b";block_ram_array(7058) := x"eb6a";block_ram_array(7060) := x"fffe";block_ram_array(7062) := x"9da0";block_ram_array(7064) := x"ffb9";block_ram_array(7066) := x"a92c";block_ram_array(7068) := x"007b";block_ram_array(7070) := x"
7f44";block_ram_array(7072) := x"0044";block_ram_array(7074) := x"fb95";block_ram_array(7076) := x"0042";block_ram_array(7078) := x"a7ae";block_ram_array(7080) := x"0002";block_ram_array(7082) := x"8b5c";block_ram_array(7084) := x"0024";block_ram_array(7086) := x"8f41";block_ram_array(7088) := x"0057";block_ram_array(7090) := x"f2bf";block_ram_array(7092) := x"0035";block_ram_array(7094) := x"85b2";block_ram_array(7096) := x"0037";block_ram_array(7098) := x"ef91";block_ram_array(7100) := x"ffea";block_ram_array(7102) := x"8448";block_ram_array(7104) := x"0059";block_ram_array(7106) := x"a723";block_ram_array(7108) := x"ffec";block_ram_array(7110) := x"ba12";block_ram_array(7112) := x"0012";block_ram_array(7114) := x"ca49";block_ram_array(7116) := x"ff87";block_ram_array(7118) := x"b7bc";block_ram_array(7120) := x"ffcb";block_ram_array(7122) := x"0a45";block_ram_array(7124) := x"ffd8";block_ram_array(7126) := x"b8aa";block_ram_array(7128) := x"ffdc";block_ram_array(7130) := x"c777";block_ram_array(7132) := x"fff4";block_ram_array(7134) := x"2464";block_ram_array(7136) := x"0003";block_ram_array(7138) := x"7205";block_ram_array(7140) := x"0000";block_ram_array(7142) := x"cb39";block_ram_array(7144) := x"ffd6";block_ram_array(7146) := x"1afb";block_ram_array(7148) := x"ffb9";block_ram_array(7150) := x"d485";block_ram_array(7152) := x"ff8a";block_ram_array(7154) := x"ec55";block_ram_array(7156) := x"0026";block_ram_array(7158) := x"8527";block_ram_array(7160) := x"ffe4";block_ram_array(7162) := x"c8ad";block_ram_array(7164) := x"0071";block_ram_array(7166) := x"6330";block_ram_array(7168) := x"0042";block_ram_array(7170) := x"e100";block_ram_array(7172) := x"0052";block_ram_array(7174) := x"4100";block_ram_array(7176) := x"002b";block_ram_array(7178) := x"cd2e";block_ram_array(7180) := x"0004";block_ram_array(7182) := x"00be";block_ram_array(7184) := x"003c";block_ram_array(7186) := x"1907";block_ram_array(7188) := x"003a";block_ram_array(7190) := x"0c17";block_ram_array(7192) := x"0068";block_ram_array(7194) := x"fd9b";block_ram_array(7196) := x"ffd1";block_ram_array(7198) := x"db8e";block_ram_array(7200) := x"002f";block_ram_array(7202) := x"086f";block_ram_array(7204) := x"ffd2";block_ram_array(7206) := x"1c92";block_ram_array(7208) := x"0028";block_ram_array(7210) := x"fd7e";block_ram_array(7212) := x"ff70";block_ram_array(7214) := x"b2de";block_ram_array(7216) := x"ff6b";block_ram_array(7218) := x"ae38";block_ram_array(7220) := x"ffc0";block_ram_array(7222) := x"49e9";block_ram_array(7224) := x"ffe3";block_ram_array(7226) := x"d6ee";block_ram_array(7228) := x"0039";block_ram_array(7230) := x"c450";block_ram_array(7232) := x"ffe0";block_ram_array(7234) := x"d2a8";block_ram_array(7236) := x"fffc";block_ram_array(7238) := x"6e2a";block_ram_array(7240) := x"fff9";block_ram_array(7242) := x"dc0c";block_ram_array(7244) := x"001a";block_ram_array(7246) := x"15fc";block_ram_array(7248) := x"ffc2";block_ram_array(7250) := x"b007";block_ram_array(7252) := x"fff7";block_ram_array(7254) := x"5425";block_ram_array(7256) := x"ffdb";block_ram_array(7258) := x"676e";block_ram_array(7260) := x"0086";block_ram_array(7262) := x"bd8d";block_ram_array(7264) := x"0079";block_ram_array(7266) := x"e8f4";block_ram_array(7268) := x"0042";block_ram_array(7270) := x"6a10";block_ram_array(7272) := x"0036";block_ram_array(7274) := x"5327";block_ram_array(7276) := x"ffd2";block_ram_array(7278) := x"2152";block_ram_array(7280) := x"000c";block_ram_array(7282) := x"8873";block_ram_array(7284) := x"0017";block_ram_array(7286) := x"e4bc";block_ram_array(7288) := x"006e";block_ram_array(7290) := x"ccbc";block_ram_array(7292) := x"fffc";block_ram_array(7294) := x"6160";block_ram_array(7296) := x"0035";block_ram_array(7298) := x"f717";block_ram_array(7300) := x"ff8c";block_ram_array(7302) := x"a49c";block_ram_array(7304) := x"ffe9";block_ram_array(7306) := x"4907";block_ram_array(7308) := x"ff92";block_ram_array(7310) := x"a558";block_ram_array(7312) := x"ff82";block_ram_array(7314) := x"b076";block_ram_array(7316) := x"ffaa";block_ram_array(7318) := x"
4320";block_ram_array(7320) := x"ff85";block_ram_array(7322) := x"a2f6";block_ram_array(7324) := x"005b";block_ram_array(7326) := x"ac97";block_ram_array(7328) := x"001a";block_ram_array(7330) := x"ed28";block_ram_array(7332) := x"0049";block_ram_array(7334) := x"6571";block_ram_array(7336) := x"fffb";block_ram_array(7338) := x"9baf";block_ram_array(7340) := x"0014";block_ram_array(7342) := x"a03c";block_ram_array(7344) := x"0002";block_ram_array(7346) := x"23fc";block_ram_array(7348) := x"0026";block_ram_array(7350) := x"fed3";block_ram_array(7352) := x"0003";block_ram_array(7354) := x"1ba6";block_ram_array(7356) := x"004b";block_ram_array(7358) := x"ddb2";block_ram_array(7360) := x"008c";block_ram_array(7362) := x"7840";block_ram_array(7364) := x"0039";block_ram_array(7366) := x"3c9b";block_ram_array(7368) := x"0041";block_ram_array(7370) := x"559c";block_ram_array(7372) := x"ff83";block_ram_array(7374) := x"93fe";block_ram_array(7376) := x"ffd1";block_ram_array(7378) := x"919e";block_ram_array(7380) := x"fffc";block_ram_array(7382) := x"37f4";block_ram_array(7384) := x"003c";block_ram_array(7386) := x"24ff";block_ram_array(7388) := x"fffd";block_ram_array(7390) := x"dd2c";block_ram_array(7392) := x"002b";block_ram_array(7394) := x"4924";block_ram_array(7396) := x"ffc3";block_ram_array(7398) := x"f408";block_ram_array(7400) := x"fff7";block_ram_array(7402) := x"6fd6";block_ram_array(7404) := x"ff6e";block_ram_array(7406) := x"8996";block_ram_array(7408) := x"ff39";block_ram_array(7410) := x"25fc";block_ram_array(7412) := x"ffd7";block_ram_array(7414) := x"8962";block_ram_array(7416) := x"ffbd";block_ram_array(7418) := x"03fa";block_ram_array(7420) := x"008a";block_ram_array(7422) := x"dda8";block_ram_array(7424) := x"000b";block_ram_array(7426) := x"fc16";block_ram_array(7428) := x"004a";block_ram_array(7430) := x"a1a0";block_ram_array(7432) := x"002f";block_ram_array(7434) := x"384f";block_ram_array(7436) := x"0047";block_ram_array(7438) := x"8595";block_ram_array(7440) := x"0032";block_ram_array(7442) := x"7ced";block_ram_array(7444) := x"000f";block_ram_array(7446) := x"ae30";block_ram_array(7448) := x"0030";block_ram_array(7450) := x"b22a";block_ram_array(7452) := x"0027";block_ram_array(7454) := x"dc84";block_ram_array(7456) := x"0081";block_ram_array(7458) := x"7aca";block_ram_array(7460) := x"0008";block_ram_array(7462) := x"7b7b";block_ram_array(7464) := x"0062";block_ram_array(7466) := x"12d1";block_ram_array(7468) := x"ff4a";block_ram_array(7470) := x"a794";block_ram_array(7472) := x"ff4a";block_ram_array(7474) := x"0035";block_ram_array(7476) := x"ffa1";block_ram_array(7478) := x"3c6d";block_ram_array(7480) := x"000e";block_ram_array(7482) := x"a3a1";block_ram_array(7484) := x"0079";block_ram_array(7486) := x"822e";block_ram_array(7488) := x"0023";block_ram_array(7490) := x"b2e6";block_ram_array(7492) := x"ffa2";block_ram_array(7494) := x"0929";block_ram_array(7496) := x"ffd7";block_ram_array(7498) := x"5c38";block_ram_array(7500) := x"ffec";block_ram_array(7502) := x"876c";block_ram_array(7504) := x"ff8d";block_ram_array(7506) := x"849c";block_ram_array(7508) := x"ffb3";block_ram_array(7510) := x"868a";block_ram_array(7512) := x"ff84";block_ram_array(7514) := x"7dd5";block_ram_array(7516) := x"00d2";block_ram_array(7518) := x"5c10";block_ram_array(7520) := x"00a0";block_ram_array(7522) := x"345a";block_ram_array(7524) := x"004d";block_ram_array(7526) := x"3b76";block_ram_array(7528) := x"000e";block_ram_array(7530) := x"1ddf";block_ram_array(7532) := x"0006";block_ram_array(7534) := x"241d";block_ram_array(7536) := x"0060";block_ram_array(7538) := x"3c7c";block_ram_array(7540) := x"0019";block_ram_array(7542) := x"55b5";block_ram_array(7544) := x"003b";block_ram_array(7546) := x"93cf";block_ram_array(7548) := x"fff7";block_ram_array(7550) := x"4f38";block_ram_array(7552) := x"008d";block_ram_array(7554) := x"8a98";block_ram_array(7556) := x"ffb8";block_ram_array(7558) := x"82ff";block_ram_array(7560) := x"fffb";block_ram_array(7562) := x"fd02";block_ram_array(7564) := x"ff35";block_ram_array(7566) := x"
0e22";block_ram_array(7568) := x"ff4e";block_ram_array(7570) := x"d0a0";block_ram_array(7572) := x"ff86";block_ram_array(7574) := x"c408";block_ram_array(7576) := x"ff4d";block_ram_array(7578) := x"b625";block_ram_array(7580) := x"0092";block_ram_array(7582) := x"9ecb";block_ram_array(7584) := x"0078";block_ram_array(7586) := x"c700";block_ram_array(7588) := x"005e";block_ram_array(7590) := x"1324";block_ram_array(7592) := x"ffdd";block_ram_array(7594) := x"e2c3";block_ram_array(7596) := x"ffb4";block_ram_array(7598) := x"6ba5";block_ram_array(7600) := x"ffbf";block_ram_array(7602) := x"a973";block_ram_array(7604) := x"0039";block_ram_array(7606) := x"86ef";block_ram_array(7608) := x"ffe5";block_ram_array(7610) := x"e417";block_ram_array(7612) := x"008d";block_ram_array(7614) := x"7528";block_ram_array(7616) := x"00d8";block_ram_array(7618) := x"ce02";block_ram_array(7620) := x"0052";block_ram_array(7622) := x"2438";block_ram_array(7624) := x"0022";block_ram_array(7626) := x"6c5e";block_ram_array(7628) := x"ff6e";block_ram_array(7630) := x"83e0";block_ram_array(7632) := x"0021";block_ram_array(7634) := x"e1c3";block_ram_array(7636) := x"002c";block_ram_array(7638) := x"a940";block_ram_array(7640) := x"003c";block_ram_array(7642) := x"f6dc";block_ram_array(7644) := x"ff99";block_ram_array(7646) := x"6c8a";block_ram_array(7648) := x"0033";block_ram_array(7650) := x"fe3a";block_ram_array(7652) := x"ffe7";block_ram_array(7654) := x"e85d";block_ram_array(7656) := x"0008";block_ram_array(7658) := x"d7b2";block_ram_array(7660) := x"feea";block_ram_array(7662) := x"b7bc";block_ram_array(7664) := x"fea3";block_ram_array(7666) := x"9e48";block_ram_array(7668) := x"ffd7";block_ram_array(7670) := x"24b3";block_ram_array(7672) := x"ff9a";block_ram_array(7674) := x"00ed";block_ram_array(7676) := x"00e1";block_ram_array(7678) := x"b48f";block_ram_array(7680) := x"0032";block_ram_array(7682) := x"c32f";block_ram_array(7684) := x"0097";block_ram_array(7686) := x"4894";block_ram_array(7688) := x"0070";block_ram_array(7690) := x"29d7";block_ram_array(7692) := x"0024";block_ram_array(7694) := x"e73a";block_ram_array(7696) := x"fffe";block_ram_array(7698) := x"b506";block_ram_array(7700) := x"fffc";block_ram_array(7702) := x"59af";block_ram_array(7704) := x"0039";block_ram_array(7706) := x"8079";block_ram_array(7708) := x"007f";block_ram_array(7710) := x"d52e";block_ram_array(7712) := x"0103";block_ram_array(7714) := x"4468";block_ram_array(7716) := x"fff1";block_ram_array(7718) := x"dbff";block_ram_array(7720) := x"002f";block_ram_array(7722) := x"6756";block_ram_array(7724) := x"fedb";block_ram_array(7726) := x"e2c6";block_ram_array(7728) := x"ff49";block_ram_array(7730) := x"6abd";block_ram_array(7732) := x"ffed";block_ram_array(7734) := x"6a58";block_ram_array(7736) := x"0050";block_ram_array(7738) := x"1b12";block_ram_array(7740) := x"0010";block_ram_array(7742) := x"9dd4";block_ram_array(7744) := x"ffd0";block_ram_array(7746) := x"3266";block_ram_array(7748) := x"ff7f";block_ram_array(7750) := x"ebe2";block_ram_array(7752) := x"ffc6";block_ram_array(7754) := x"4ea0";block_ram_array(7756) := x"ffbe";block_ram_array(7758) := x"fa7e";block_ram_array(7760) := x"fefb";block_ram_array(7762) := x"73c4";block_ram_array(7764) := x"ffb3";block_ram_array(7766) := x"7409";block_ram_array(7768) := x"ff52";block_ram_array(7770) := x"e40a";block_ram_array(7772) := x"015e";block_ram_array(7774) := x"7614";block_ram_array(7776) := x"00e6";block_ram_array(7778) := x"d429";block_ram_array(7780) := x"00b4";block_ram_array(7782) := x"23c8";block_ram_array(7784) := x"006f";block_ram_array(7786) := x"8f80";block_ram_array(7788) := x"ffff";block_ram_array(7790) := x"611a";block_ram_array(7792) := x"0071";block_ram_array(7794) := x"42ef";block_ram_array(7796) := x"fff7";block_ram_array(7798) := x"70b5";block_ram_array(7800) := x"0054";block_ram_array(7802) := x"cbf8";block_ram_array(7804) := x"000d";block_ram_array(7806) := x"9dd4";block_ram_array(7808) := x"0100";block_ram_array(7810) := x"503e";block_ram_array(7812) := x"ff86";block_ram_array(7814) := x"
4197";block_ram_array(7816) := x"ffb9";block_ram_array(7818) := x"cf11";block_ram_array(7820) := x"fe8c";block_ram_array(7822) := x"0ae8";block_ram_array(7824) := x"feef";block_ram_array(7826) := x"c510";block_ram_array(7828) := x"ffd7";block_ram_array(7830) := x"d223";block_ram_array(7832) := x"ff95";block_ram_array(7834) := x"b524";block_ram_array(7836) := x"0063";block_ram_array(7838) := x"fb37";block_ram_array(7840) := x"001f";block_ram_array(7842) := x"9068";block_ram_array(7844) := x"002b";block_ram_array(7846) := x"10a8";block_ram_array(7848) := x"ffa1";block_ram_array(7850) := x"d478";block_ram_array(7852) := x"ffa5";block_ram_array(7854) := x"4665";block_ram_array(7856) := x"ff43";block_ram_array(7858) := x"33f4";block_ram_array(7860) := x"0088";block_ram_array(7862) := x"b91a";block_ram_array(7864) := x"0003";block_ram_array(7866) := x"e515";block_ram_array(7868) := x"00f9";block_ram_array(7870) := x"5f1c";block_ram_array(7872) := x"00e0";block_ram_array(7874) := x"df14";block_ram_array(7876) := x"00ab";block_ram_array(7878) := x"1841";block_ram_array(7880) := x"00c1";block_ram_array(7882) := x"f3de";block_ram_array(7884) := x"ffa9";block_ram_array(7886) := x"fb74";block_ram_array(7888) := x"005d";block_ram_array(7890) := x"bd21";block_ram_array(7892) := x"ffc9";block_ram_array(7894) := x"6f01";block_ram_array(7896) := x"004f";block_ram_array(7898) := x"c9dd";block_ram_array(7900) := x"ff8c";block_ram_array(7902) := x"9650";block_ram_array(7904) := x"0084";block_ram_array(7906) := x"d254";block_ram_array(7908) := x"ff9b";block_ram_array(7910) := x"8ed6";block_ram_array(7912) := x"ffc2";block_ram_array(7914) := x"7e4a";block_ram_array(7916) := x"fe34";block_ram_array(7918) := x"ef10";block_ram_array(7920) := x"fdf4";block_ram_array(7922) := x"0404";block_ram_array(7924) := x"001f";block_ram_array(7926) := x"a2e3";block_ram_array(7928) := x"fff2";block_ram_array(7930) := x"fc98";block_ram_array(7932) := x"00fa";block_ram_array(7934) := x"3d7a";block_ram_array(7936) := x"ffc0";block_ram_array(7938) := x"d64b";block_ram_array(7940) := x"004e";block_ram_array(7942) := x"414b";block_ram_array(7944) := x"0048";block_ram_array(7946) := x"b36b";block_ram_array(7948) := x"0066";block_ram_array(7950) := x"de27";block_ram_array(7952) := x"ff97";block_ram_array(7954) := x"e80e";block_ram_array(7956) := x"0028";block_ram_array(7958) := x"02e7";block_ram_array(7960) := x"0075";block_ram_array(7962) := x"05d7";block_ram_array(7964) := x"0121";block_ram_array(7966) := x"c8e6";block_ram_array(7968) := x"0121";block_ram_array(7970) := x"d5ee";block_ram_array(7972) := x"ffeb";block_ram_array(7974) := x"42fb";block_ram_array(7976) := x"008a";block_ram_array(7978) := x"dc30";block_ram_array(7980) := x"ff62";block_ram_array(7982) := x"f3f0";block_ram_array(7984) := x"fff7";block_ram_array(7986) := x"c82c";block_ram_array(7988) := x"ff81";block_ram_array(7990) := x"eb2c";block_ram_array(7992) := x"0048";block_ram_array(7994) := x"7922";block_ram_array(7996) := x"ffb4";block_ram_array(7998) := x"a1a4";block_ram_array(8000) := x"fff0";block_ram_array(8002) := x"778f";block_ram_array(8004) := x"ff31";block_ram_array(8006) := x"02f1";block_ram_array(8008) := x"ff93";block_ram_array(8010) := x"8e22";block_ram_array(8012) := x"ff29";block_ram_array(8014) := x"4f36";block_ram_array(8016) := x"fe31";block_ram_array(8018) := x"3fe0";block_ram_array(8020) := x"ffa0";block_ram_array(8022) := x"ed9d";block_ram_array(8024) := x"ff48";block_ram_array(8026) := x"c60c";block_ram_array(8028) := x"01d8";block_ram_array(8030) := x"9a5c";block_ram_array(8032) := x"00bf";block_ram_array(8034) := x"e531";block_ram_array(8036) := x"0077";block_ram_array(8038) := x"b214";block_ram_array(8040) := x"000e";block_ram_array(8042) := x"81fd";block_ram_array(8044) := x"0065";block_ram_array(8046) := x"c7d0";block_ram_array(8048) := x"0067";block_ram_array(8050) := x"cdc9";block_ram_array(8052) := x"0046";block_ram_array(8054) := x"aee9";block_ram_array(8056) := x"0087";block_ram_array(8058) := x"7fbe";block_ram_array(8060) := x"0095";block_ram_array(8062) := x"
3410";block_ram_array(8064) := x"0152";block_ram_array(8066) := x"9a94";block_ram_array(8068) := x"ff7a";block_ram_array(8070) := x"b165";block_ram_array(8072) := x"ffef";block_ram_array(8074) := x"a695";block_ram_array(8076) := x"fefa";block_ram_array(8078) := x"3f34";block_ram_array(8080) := x"ffd6";block_ram_array(8082) := x"8a59";block_ram_array(8084) := x"ff83";block_ram_array(8086) := x"d2a4";block_ram_array(8088) := x"ff8b";block_ram_array(8090) := x"21e8";block_ram_array(8092) := x"ffb9";block_ram_array(8094) := x"57f8";block_ram_array(8096) := x"0016";block_ram_array(8098) := x"5fb5";block_ram_array(8100) := x"ffcb";block_ram_array(8102) := x"8d52";block_ram_array(8104) := x"ff4a";block_ram_array(8106) := x"73c2";block_ram_array(8108) := x"ff22";block_ram_array(8110) := x"67c2";block_ram_array(8112) := x"fe8b";block_ram_array(8114) := x"924e";block_ram_array(8116) := x"0060";block_ram_array(8118) := x"f205";block_ram_array(8120) := x"ff85";block_ram_array(8122) := x"029e";block_ram_array(8124) := x"0173";block_ram_array(8126) := x"2fa6";block_ram_array(8128) := x"00cb";block_ram_array(8130) := x"83e8";block_ram_array(8132) := x"00f5";block_ram_array(8134) := x"f903";block_ram_array(8136) := x"009e";block_ram_array(8138) := x"202a";block_ram_array(8140) := x"0019";block_ram_array(8142) := x"38c2";block_ram_array(8144) := x"007b";block_ram_array(8146) := x"e3a5";block_ram_array(8148) := x"0024";block_ram_array(8150) := x"7047";block_ram_array(8152) := x"00a3";block_ram_array(8154) := x"e932";block_ram_array(8156) := x"0016";block_ram_array(8158) := x"43a3";block_ram_array(8160) := x"012b";block_ram_array(8162) := x"c338";block_ram_array(8164) := x"ff65";block_ram_array(8166) := x"2d16";block_ram_array(8168) := x"ffbe";block_ram_array(8170) := x"7053";block_ram_array(8172) := x"fe47";block_ram_array(8174) := x"7712";block_ram_array(8176) := x"fedb";block_ram_array(8178) := x"e084";block_ram_array(8180) := x"fff3";block_ram_array(8182) := x"d370";block_ram_array(8184) := x"ffe1";block_ram_array(8186) := x"e677";block_ram_array(8188) := x"fff8";block_ram_array(8190) := x"f7ac";
        
    elsif (clk'event and clk='1') then
        
        s_waitrequest <= '0';
        
        if s_read = '1' then
            
            if fill_block_28 = '1' then
                
                if skip = '1' then skip := '0';
                else
                
                --------------------
                --=28
                --------------------
                block_ram_array(114688) := x"001a";block_ram_array(114690) := x"e800";block_ram_array(114692) := x"0000";block_ram_array(114694) := x"0000";block_ram_array(114696) := x"f92e";block_ram_array(114698) := x"0240";block_ram_array(114700) := x"fc34";block_ram_array(114702) := x"7d88";block_ram_array(114704) := x"f7d7";block_ram_array(114706) := x"c620";block_ram_array(114708) := x"05b7";block_ram_array(114710) := x"4b50";block_ram_array(114712) := x"ffad";block_ram_array(114714) := x"3d9b";block_ram_array(114716) := x"0572";block_ram_array(114718) := x"fc60";block_ram_array(114720) := x"013a";block_ram_array(114722) := x"2068";block_ram_array(114724) := x"020a";block_ram_array(114726) := x"6600";block_ram_array(114728) := x"fd57";block_ram_array(114730) := x"98b0";block_ram_array(114732) := x"fc0a";block_ram_array(114734) := x"2b4c";block_ram_array(114736) := x"f77a";block_ram_array(114738) := x"f910";block_ram_array(114740) := x"05e2";block_ram_array(114742) := x"9ea0";block_ram_array(114744) := x"0182";block_ram_array(114746) := x"bf70";block_ram_array(114748) := x"042c";block_ram_array(114750) := x"a728";block_ram_array(114752) := x"fa07";block_ram_array(114754) := x"0750";block_ram_array(114756) := x"05cc";block_ram_array(114758) := x"1718";block_ram_array(114760) := x"0743";block_ram_array(114762) := x"3e18";block_ram_array(114764) := x"086c";block_ram_array(114766) := x"81a0";block_ram_array(114768) := x"008b";block_ram_array(114770) := x"f68a";block_ram_array(114772) := x"fdd0";block_ram_array(114774) := x"897c";block_ram_array(114776) := x"0217";block_ram_array(114778) := x"0c58";block_ram_array(114780) := x"05e8";block_ram_array(114782) := x"fd18";block_ram_array(114784) := x"03cb";block_ram_array(114786) := x"17f0";block_ram_array(114788) := x"fed1";block_ram_array(114790) := x"fe88";block_ram_array(114792) := x"0143";block_ram_array(114794) := x"2fb6";block_ram_array(114796) := x"002d";block_ram_array(114798) := x"8bc6";block_ram_array(114800) := x"fee7";block_ram_array(114802) := x"8f66";block_ram_array(114804) := x"ff74";block_ram_array(114806) := x"aef4";block_ram_array(114808) := x"0235";block_ram_array(114810) := x"b7b8";block_ram_array(114812) := x"03de";block_ram_array(114814) := x"f770";block_ram_array(114816) := x"01f4";block_ram_array(114818) := x"f0fc";block_ram_array(114820) := x"fcf4";block_ram_array(114822) := x"5c24";block_ram_array(114824) := x"fea8";block_ram_array(114826) := x"009e";block_ram_array(114828) := x"0271";block_ram_array(114830) := x"3064";block_ram_array(114832) := x"0366";block_ram_array(114834) := x"2bf0";block_ram_array(114836) := x"ff8e";block_ram_array(114838) := x"493a";block_ram_array(114840) := x"ff04";block_ram_array(114842) := x"5452";block_ram_array(114844) := x"ff04";block_ram_array(114846) := x"68da";block_ram_array(114848) := x"0069";block_ram_array(114850) := x"3b9a";block_ram_array(114852) := x"00c3";block_ram_array(114854) := x"a6ac";block_ram_array(114856) := x"000e";block_ram_array(114858) := x"5bf2";block_ram_array(114860) := x"003c";block_ram_array(114862) := x"0b59";block_ram_array(114864) := x"0059";block_ram_array(114866) := x"d692";block_ram_array(114868) := x"0108";block_ram_array(114870) := x"886c";block_ram_array(114872) := x"016e";block_ram_array(114874) := x"fc34";block_ram_array(114876) := x"00e5";block_ram_array(114878) := x"97fc";block_ram_array(114880) := x"01d2";block_ram_array(114882) := x"46c0";block_ram_array(114884) := x"ff8a";block_ram_array(114886) := x"5f3d";block_ram_array(114888) := x"0098";block_ram_array(114890) := x"6818";block_ram_array(114892) := x"fe69";block_ram_array(114894) := x"aec4";block_ram_array(114896) := x"ff0e";block_ram_array(114898) := x"1764";block_ram_array(114900) := x"ffb3";block_ram_array(114902) := x"a163";block_ram_array(114904) := x"008e";block_ram_array(114906) := x"4df6";block_ram_array(114908) := x"0064";block_ram_array(114910) := x"b71a";block_ram_array(114912) := x"ffe8";block_ram_array(114914) := x"0eee";block_ram_array(114916) := x"ff7d";block_ram_array(114918) := x"8738";block_ram_array(
114920) := x"ffe7";block_ram_array(114922) := x"2434";block_ram_array(114924) := x"005f";block_ram_array(114926) := x"15dd";block_ram_array(114928) := x"0097";block_ram_array(114930) := x"cec2";block_ram_array(114932) := x"0083";block_ram_array(114934) := x"6ed4";block_ram_array(114936) := x"00e0";block_ram_array(114938) := x"85de";block_ram_array(114940) := x"fed1";block_ram_array(114942) := x"9cc4";block_ram_array(114944) := x"fe77";block_ram_array(114946) := x"7f50";block_ram_array(114948) := x"0051";block_ram_array(114950) := x"6136";block_ram_array(114952) := x"01ec";block_ram_array(114954) := x"71ec";block_ram_array(114956) := x"0086";block_ram_array(114958) := x"3528";block_ram_array(114960) := x"fee5";block_ram_array(114962) := x"af70";block_ram_array(114964) := x"fe85";block_ram_array(114966) := x"b3dc";block_ram_array(114968) := x"0095";block_ram_array(114970) := x"f2e1";block_ram_array(114972) := x"0132";block_ram_array(114974) := x"7dca";block_ram_array(114976) := x"ffc5";block_ram_array(114978) := x"79ae";block_ram_array(114980) := x"feb0";block_ram_array(114982) := x"bc54";block_ram_array(114984) := x"001b";block_ram_array(114986) := x"a8eb";block_ram_array(114988) := x"00a2";block_ram_array(114990) := x"702f";block_ram_array(114992) := x"ff2d";block_ram_array(114994) := x"ebd6";block_ram_array(114996) := x"fecd";block_ram_array(114998) := x"9eac";block_ram_array(115000) := x"ffa6";block_ram_array(115002) := x"ddb7";block_ram_array(115004) := x"01b2";block_ram_array(115006) := x"7184";block_ram_array(115008) := x"006b";block_ram_array(115010) := x"713b";block_ram_array(115012) := x"ff10";block_ram_array(115014) := x"3854";block_ram_array(115016) := x"ff0b";block_ram_array(115018) := x"1014";block_ram_array(115020) := x"0103";block_ram_array(115022) := x"14e0";block_ram_array(115024) := x"007b";block_ram_array(115026) := x"b6dd";block_ram_array(115028) := x"0051";block_ram_array(115030) := x"0898";block_ram_array(115032) := x"0030";block_ram_array(115034) := x"a615";block_ram_array(115036) := x"00cc";block_ram_array(115038) := x"9510";block_ram_array(115040) := x"00b7";block_ram_array(115042) := x"cf1a";block_ram_array(115044) := x"ffb6";block_ram_array(115046) := x"dd5d";block_ram_array(115048) := x"0003";block_ram_array(115050) := x"8b36";block_ram_array(115052) := x"0033";block_ram_array(115054) := x"ee73";block_ram_array(115056) := x"003a";block_ram_array(115058) := x"4f03";block_ram_array(115060) := x"ffc2";block_ram_array(115062) := x"7f72";block_ram_array(115064) := x"0013";block_ram_array(115066) := x"5964";block_ram_array(115068) := x"006c";block_ram_array(115070) := x"7fc7";block_ram_array(115072) := x"0066";block_ram_array(115074) := x"ad43";block_ram_array(115076) := x"ffa6";block_ram_array(115078) := x"b330";block_ram_array(115080) := x"ffe1";block_ram_array(115082) := x"5fa9";block_ram_array(115084) := x"0025";block_ram_array(115086) := x"3749";block_ram_array(115088) := x"0021";block_ram_array(115090) := x"fd49";block_ram_array(115092) := x"fff7";block_ram_array(115094) := x"2d69";block_ram_array(115096) := x"0040";block_ram_array(115098) := x"fe67";block_ram_array(115100) := x"0048";block_ram_array(115102) := x"07ba";block_ram_array(115104) := x"0035";block_ram_array(115106) := x"0041";block_ram_array(115108) := x"ffaf";block_ram_array(115110) := x"8ec5";block_ram_array(115112) := x"0034";block_ram_array(115114) := x"6e1e";block_ram_array(115116) := x"0027";block_ram_array(115118) := x"a482";block_ram_array(115120) := x"000e";block_ram_array(115122) := x"256f";block_ram_array(115124) := x"ff81";block_ram_array(115126) := x"ef07";block_ram_array(115128) := x"fff4";block_ram_array(115130) := x"81d0";block_ram_array(115132) := x"003a";block_ram_array(115134) := x"c138";block_ram_array(115136) := x"0007";block_ram_array(115138) := x"daad";block_ram_array(115140) := x"ffa8";block_ram_array(115142) := x"f9cc";block_ram_array(115144) := x"fffa";block_ram_array(115146) := x"f3b9";block_ram_array(115148) := x"0049";block_ram_array(115150) := x"e4ad";block_ram_array(115152) := x"0011";block_ram_array(
115154) := x"7bed";block_ram_array(115156) := x"ffab";block_ram_array(115158) := x"9da6";block_ram_array(115160) := x"fff5";block_ram_array(115162) := x"df4e";block_ram_array(115164) := x"0047";block_ram_array(115166) := x"d8f5";block_ram_array(115168) := x"0013";block_ram_array(115170) := x"5d7d";block_ram_array(115172) := x"ffb1";block_ram_array(115174) := x"7cc4";block_ram_array(115176) := x"fff3";block_ram_array(115178) := x"4499";block_ram_array(115180) := x"0046";block_ram_array(115182) := x"1bbe";block_ram_array(115184) := x"0014";block_ram_array(115186) := x"13cd";block_ram_array(115188) := x"ffb6";block_ram_array(115190) := x"50da";block_ram_array(115192) := x"fff1";block_ram_array(115194) := x"9e6d";block_ram_array(115196) := x"0044";block_ram_array(115198) := x"90c0";block_ram_array(115200) := x"0014";block_ram_array(115202) := x"a46b";block_ram_array(115204) := x"ffba";block_ram_array(115206) := x"394e";block_ram_array(115208) := x"fff0";block_ram_array(115210) := x"4e6b";block_ram_array(115212) := x"0042";block_ram_array(115214) := x"f10f";block_ram_array(115216) := x"0015";block_ram_array(115218) := x"1ccf";block_ram_array(115220) := x"ffbd";block_ram_array(115222) := x"9cb6";block_ram_array(115224) := x"ffef";block_ram_array(115226) := x"4432";block_ram_array(115228) := x"0041";block_ram_array(115230) := x"4887";block_ram_array(115232) := x"0015";block_ram_array(115234) := x"9297";block_ram_array(115236) := x"ffc0";block_ram_array(115238) := x"90e7";block_ram_array(115240) := x"ffee";block_ram_array(115242) := x"6142";block_ram_array(115244) := x"003f";block_ram_array(115246) := x"8771";block_ram_array(115248) := x"0015";block_ram_array(115250) := x"ee98";block_ram_array(115252) := x"ffc3";block_ram_array(115254) := x"2c7f";block_ram_array(115256) := x"ffed";block_ram_array(115258) := x"85bb";block_ram_array(115260) := x"003d";block_ram_array(115262) := x"c596";block_ram_array(115264) := x"0016";block_ram_array(115266) := x"3243";block_ram_array(115268) := x"ffc5";block_ram_array(115270) := x"a7b8";block_ram_array(115272) := x"ffec";block_ram_array(115274) := x"dd8c";block_ram_array(115276) := x"003c";block_ram_array(115278) := x"1953";block_ram_array(115280) := x"0016";block_ram_array(115282) := x"7932";block_ram_array(115284) := x"ffc7";block_ram_array(115286) := x"dd38";block_ram_array(115288) := x"ffec";block_ram_array(115290) := x"4131";block_ram_array(115292) := x"003a";block_ram_array(115294) := x"6d24";block_ram_array(115296) := x"0016";block_ram_array(115298) := x"b383";block_ram_array(115300) := x"ffc9";block_ram_array(115302) := x"e35c";block_ram_array(115304) := x"ffeb";block_ram_array(115306) := x"a3c6";block_ram_array(115308) := x"0038";block_ram_array(115310) := x"ca92";block_ram_array(115312) := x"0016";block_ram_array(115314) := x"df78";block_ram_array(115316) := x"ffcb";block_ram_array(115318) := x"e110";block_ram_array(115320) := x"ffeb";block_ram_array(115322) := x"360c";block_ram_array(115324) := x"0037";block_ram_array(115326) := x"4174";block_ram_array(115328) := x"0017";block_ram_array(115330) := x"19b8";block_ram_array(115332) := x"ffcd";block_ram_array(115334) := x"9d18";block_ram_array(115336) := x"ffea";block_ram_array(115338) := x"b413";block_ram_array(115340) := x"0035";block_ram_array(115342) := x"aa2d";block_ram_array(115344) := x"0017";block_ram_array(115346) := x"334c";block_ram_array(115348) := x"ffcf";block_ram_array(115350) := x"5f98";block_ram_array(115352) := x"ffea";block_ram_array(115354) := x"6670";block_ram_array(115356) := x"0034";block_ram_array(115358) := x"326a";block_ram_array(115360) := x"0017";block_ram_array(115362) := x"4baf";block_ram_array(115364) := x"ffd0";block_ram_array(115366) := x"d7ce";block_ram_array(115368) := x"ffe9";block_ram_array(115370) := x"f0a8";block_ram_array(115372) := x"0032";block_ram_array(115374) := x"d371";block_ram_array(115376) := x"0017";block_ram_array(115378) := x"7799";block_ram_array(115380) := x"ffd2";block_ram_array(115382) := x"5fbc";block_ram_array(115384) := x"ffe9";block_ram_array(115386) := x"9531";block_ram_array(
115388) := x"0031";block_ram_array(115390) := x"6168";block_ram_array(115392) := x"0017";block_ram_array(115394) := x"7b09";block_ram_array(115396) := x"ffd3";block_ram_array(115398) := x"d616";block_ram_array(115400) := x"ffe9";block_ram_array(115402) := x"5069";block_ram_array(115404) := x"0030";block_ram_array(115406) := x"1fee";block_ram_array(115408) := x"0017";block_ram_array(115410) := x"936f";block_ram_array(115412) := x"ffd5";block_ram_array(115414) := x"2b7a";block_ram_array(115416) := x"ffe9";block_ram_array(115418) := x"1053";block_ram_array(115420) := x"002e";block_ram_array(115422) := x"eb72";block_ram_array(115424) := x"0017";block_ram_array(115426) := x"c7da";block_ram_array(115428) := x"ffd6";block_ram_array(115430) := x"6154";block_ram_array(115432) := x"ffe8";block_ram_array(115434) := x"bc68";block_ram_array(115436) := x"002d";block_ram_array(115438) := x"9072";block_ram_array(115440) := x"0017";block_ram_array(115442) := x"c98b";block_ram_array(115444) := x"ffd7";block_ram_array(115446) := x"a2f3";block_ram_array(115448) := x"ffe8";block_ram_array(115450) := x"83cf";block_ram_array(115452) := x"002c";block_ram_array(115454) := x"5c60";block_ram_array(115456) := x"0017";block_ram_array(115458) := x"c9d0";block_ram_array(115460) := x"ffd8";block_ram_array(115462) := x"c73d";block_ram_array(115464) := x"ffe8";block_ram_array(115466) := x"477c";block_ram_array(115468) := x"002b";block_ram_array(115470) := x"4814";block_ram_array(115472) := x"0017";block_ram_array(115474) := x"e92d";block_ram_array(115476) := x"ffd9";block_ram_array(115478) := x"e07d";block_ram_array(115480) := x"ffe8";block_ram_array(115482) := x"0c2e";block_ram_array(115484) := x"002a";block_ram_array(115486) := x"18fd";block_ram_array(115488) := x"0017";block_ram_array(115490) := x"e0cd";block_ram_array(115492) := x"ffda";block_ram_array(115494) := x"f32c";block_ram_array(115496) := x"ffe7";block_ram_array(115498) := x"d8b5";block_ram_array(115500) := x"0029";block_ram_array(115502) := x"1b82";block_ram_array(115504) := x"0018";block_ram_array(115506) := x"01f9";block_ram_array(115508) := x"ffdb";block_ram_array(115510) := x"fbc5";block_ram_array(115512) := x"ffe7";block_ram_array(115514) := x"b1ae";block_ram_array(115516) := x"0027";block_ram_array(115518) := x"f97a";block_ram_array(115520) := x"0017";block_ram_array(115522) := x"f3b0";block_ram_array(115524) := x"ffdc";block_ram_array(115526) := x"e8a6";block_ram_array(115528) := x"ffe7";block_ram_array(115530) := x"797b";block_ram_array(115532) := x"0027";block_ram_array(115534) := x"0861";block_ram_array(115536) := x"0017";block_ram_array(115538) := x"f943";block_ram_array(115540) := x"ffdd";block_ram_array(115542) := x"d6e9";block_ram_array(115544) := x"ffe7";block_ram_array(115546) := x"3772";block_ram_array(115548) := x"0026";block_ram_array(115550) := x"3091";block_ram_array(115552) := x"0018";block_ram_array(115554) := x"4494";block_ram_array(115556) := x"ffde";block_ram_array(115558) := x"e7f1";block_ram_array(115560) := x"ffe7";block_ram_array(115562) := x"3d3d";block_ram_array(115564) := x"0024";block_ram_array(115566) := x"e260";block_ram_array(115568) := x"0017";block_ram_array(115570) := x"ea82";block_ram_array(115572) := x"ffdf";block_ram_array(115574) := x"a1fd";block_ram_array(115576) := x"ffe6";block_ram_array(115578) := x"ff44";block_ram_array(115580) := x"0024";block_ram_array(115582) := x"47d0";block_ram_array(115584) := x"0018";block_ram_array(115586) := x"25ae";block_ram_array(115588) := x"ffe0";block_ram_array(115590) := x"84bb";block_ram_array(115592) := x"ffe6";block_ram_array(115594) := x"d628";block_ram_array(115596) := x"0023";block_ram_array(115598) := x"44f0";block_ram_array(115600) := x"0018";block_ram_array(115602) := x"191e";block_ram_array(115604) := x"ffe1";block_ram_array(115606) := x"70c9";block_ram_array(115608) := x"ffe6";block_ram_array(115610) := x"e3a8";block_ram_array(115612) := x"0022";block_ram_array(115614) := x"6ad3";block_ram_array(115616) := x"0018";block_ram_array(115618) := x"098a";block_ram_array(115620) := x"ffe2";block_ram_array(
115622) := x"059a";block_ram_array(115624) := x"ffe6";block_ram_array(115626) := x"956c";block_ram_array(115628) := x"0021";block_ram_array(115630) := x"bbe5";block_ram_array(115632) := x"0018";block_ram_array(115634) := x"32db";block_ram_array(115636) := x"ffe2";block_ram_array(115638) := x"f4c1";block_ram_array(115640) := x"ffe6";block_ram_array(115642) := x"b00a";block_ram_array(115644) := x"0020";block_ram_array(115646) := x"de42";block_ram_array(115648) := x"0018";block_ram_array(115650) := x"42ae";block_ram_array(115652) := x"ffe3";block_ram_array(115654) := x"6656";block_ram_array(115656) := x"ffe6";block_ram_array(115658) := x"4471";block_ram_array(115660) := x"001f";block_ram_array(115662) := x"fd21";block_ram_array(115664) := x"0018";block_ram_array(115666) := x"3244";block_ram_array(115668) := x"ffe4";block_ram_array(115670) := x"5590";block_ram_array(115672) := x"ffe6";block_ram_array(115674) := x"37aa";block_ram_array(115676) := x"001f";block_ram_array(115678) := x"418a";block_ram_array(115680) := x"0018";block_ram_array(115682) := x"2a9e";block_ram_array(115684) := x"ffe5";block_ram_array(115686) := x"227a";block_ram_array(115688) := x"ffe6";block_ram_array(115690) := x"5572";block_ram_array(115692) := x"001e";block_ram_array(115694) := x"a8d0";block_ram_array(115696) := x"0018";block_ram_array(115698) := x"6704";block_ram_array(115700) := x"ffe5";block_ram_array(115702) := x"8a82";block_ram_array(115704) := x"ffe5";block_ram_array(115706) := x"f8e7";block_ram_array(115708) := x"001d";block_ram_array(115710) := x"bbde";block_ram_array(115712) := x"0018";block_ram_array(115714) := x"4f00";block_ram_array(115716) := x"ffe6";block_ram_array(115718) := x"6900";block_ram_array(115720) := x"ffe6";block_ram_array(115722) := x"02b1";block_ram_array(115724) := x"001d";block_ram_array(115726) := x"1192";block_ram_array(115728) := x"0018";block_ram_array(115730) := x"5de8";block_ram_array(115732) := x"ffe6";block_ram_array(115734) := x"fec6";block_ram_array(115736) := x"ffe5";block_ram_array(115738) := x"ea0a";block_ram_array(115740) := x"001c";block_ram_array(115742) := x"5198";block_ram_array(115744) := x"0018";block_ram_array(115746) := x"5726";block_ram_array(115748) := x"ffe7";block_ram_array(115750) := x"9a30";block_ram_array(115752) := x"ffe5";block_ram_array(115754) := x"caa8";block_ram_array(115756) := x"001b";block_ram_array(115758) := x"a8ea";block_ram_array(115760) := x"0018";block_ram_array(115762) := x"5ffc";block_ram_array(115764) := x"ffe8";block_ram_array(115766) := x"44a8";block_ram_array(115768) := x"ffe5";block_ram_array(115770) := x"c4b1";block_ram_array(115772) := x"001a";block_ram_array(115774) := x"f7e1";block_ram_array(115776) := x"0018";block_ram_array(115778) := x"5eea";block_ram_array(115780) := x"ffe8";block_ram_array(115782) := x"d3e2";block_ram_array(115784) := x"ffe5";block_ram_array(115786) := x"ae3a";block_ram_array(115788) := x"001a";block_ram_array(115790) := x"51e2";block_ram_array(115792) := x"0018";block_ram_array(115794) := x"619b";block_ram_array(115796) := x"ffe9";block_ram_array(115798) := x"6aa1";block_ram_array(115800) := x"ffe5";block_ram_array(115802) := x"a178";block_ram_array(115804) := x"0019";block_ram_array(115806) := x"af61";block_ram_array(115808) := x"0018";block_ram_array(115810) := x"6754";block_ram_array(115812) := x"ffe9";block_ram_array(115814) := x"f229";block_ram_array(115816) := x"ffe5";block_ram_array(115818) := x"84f2";block_ram_array(115820) := x"0019";block_ram_array(115822) := x"0bb1";block_ram_array(115824) := x"0018";block_ram_array(115826) := x"693d";block_ram_array(115828) := x"ffea";block_ram_array(115830) := x"8841";block_ram_array(115832) := x"ffe5";block_ram_array(115834) := x"749c";block_ram_array(115836) := x"0018";block_ram_array(115838) := x"6ce8";block_ram_array(115840) := x"0018";block_ram_array(115842) := x"6d7c";block_ram_array(115844) := x"ffeb";block_ram_array(115846) := x"1c9b";block_ram_array(115848) := x"ffe5";block_ram_array(115850) := x"7174";block_ram_array(115852) := x"0017";block_ram_array(115854) := x"c7a0";block_ram_array(
115856) := x"0018";block_ram_array(115858) := x"5c36";block_ram_array(115860) := x"ffeb";block_ram_array(115862) := x"a1f1";block_ram_array(115864) := x"ffe5";block_ram_array(115866) := x"71a8";block_ram_array(115868) := x"0017";block_ram_array(115870) := x"4379";block_ram_array(115872) := x"0018";block_ram_array(115874) := x"67e0";block_ram_array(115876) := x"ffec";block_ram_array(115878) := x"0d27";block_ram_array(115880) := x"ffe5";block_ram_array(115882) := x"4e73";block_ram_array(115884) := x"0016";block_ram_array(115886) := x"afc3";block_ram_array(115888) := x"0018";block_ram_array(115890) := x"6ddb";block_ram_array(115892) := x"ffec";block_ram_array(115894) := x"96ca";block_ram_array(115896) := x"ffe5";block_ram_array(115898) := x"3d6f";block_ram_array(115900) := x"0016";block_ram_array(115902) := x"1c31";block_ram_array(115904) := x"0018";block_ram_array(115906) := x"6f32";block_ram_array(115908) := x"ffed";block_ram_array(115910) := x"1eea";block_ram_array(115912) := x"ffe5";block_ram_array(115914) := x"3bb8";block_ram_array(115916) := x"0015";block_ram_array(115918) := x"8eb1";block_ram_array(115920) := x"0018";block_ram_array(115922) := x"73b4";block_ram_array(115924) := x"ffed";block_ram_array(115926) := x"90f0";block_ram_array(115928) := x"ffe5";block_ram_array(115930) := x"2b2d";block_ram_array(115932) := x"0014";block_ram_array(115934) := x"fcf1";block_ram_array(115936) := x"0018";block_ram_array(115938) := x"68bf";block_ram_array(115940) := x"ffee";block_ram_array(115942) := x"0621";block_ram_array(115944) := x"ffe5";block_ram_array(115946) := x"1a53";block_ram_array(115948) := x"0014";block_ram_array(115950) := x"8929";block_ram_array(115952) := x"0018";block_ram_array(115954) := x"8224";block_ram_array(115956) := x"ffee";block_ram_array(115958) := x"719d";block_ram_array(115960) := x"ffe4";block_ram_array(115962) := x"e945";block_ram_array(115964) := x"0013";block_ram_array(115966) := x"f84a";block_ram_array(115968) := x"0018";block_ram_array(115970) := x"9582";block_ram_array(115972) := x"ffef";block_ram_array(115974) := x"18c2";block_ram_array(115976) := x"ffe5";block_ram_array(115978) := x"0280";block_ram_array(115980) := x"0013";block_ram_array(115982) := x"47e2";block_ram_array(115984) := x"0018";block_ram_array(115986) := x"63b3";block_ram_array(115988) := x"ffef";block_ram_array(115990) := x"84d9";block_ram_array(115992) := x"ffe5";block_ram_array(115994) := x"0887";block_ram_array(115996) := x"0012";block_ram_array(115998) := x"eabe";block_ram_array(116000) := x"0018";block_ram_array(116002) := x"7257";block_ram_array(116004) := x"ffef";block_ram_array(116006) := x"de90";block_ram_array(116008) := x"ffe4";block_ram_array(116010) := x"ef2c";block_ram_array(116012) := x"0012";block_ram_array(116014) := x"70d4";block_ram_array(116016) := x"0018";block_ram_array(116018) := x"8383";block_ram_array(116020) := x"fff0";block_ram_array(116022) := x"4b2d";block_ram_array(116024) := x"ffe4";block_ram_array(116026) := x"ccad";block_ram_array(116028) := x"0011";block_ram_array(116030) := x"df4d";block_ram_array(116032) := x"0018";block_ram_array(116034) := x"6f56";block_ram_array(116036) := x"fff0";block_ram_array(116038) := x"e526";block_ram_array(116040) := x"ffe4";block_ram_array(116042) := x"fc9c";block_ram_array(116044) := x"0011";block_ram_array(116046) := x"770d";block_ram_array(116048) := x"0018";block_ram_array(116050) := x"7aeb";block_ram_array(116052) := x"fff1";block_ram_array(116054) := x"11b3";block_ram_array(116056) := x"ffe4";block_ram_array(116058) := x"b79e";block_ram_array(116060) := x"0010";block_ram_array(116062) := x"ffaa";block_ram_array(116064) := x"0018";block_ram_array(116066) := x"848d";block_ram_array(116068) := x"fff1";block_ram_array(116070) := x"a21c";block_ram_array(116072) := x"ffe4";block_ram_array(116074) := x"a963";block_ram_array(116076) := x"0010";block_ram_array(116078) := x"8191";block_ram_array(116080) := x"0018";block_ram_array(116082) := x"7c43";block_ram_array(116084) := x"fff2";block_ram_array(116086) := x"3e69";block_ram_array(116088) := x"ffe4";block_ram_array(
116090) := x"e1e2";block_ram_array(116092) := x"0010";block_ram_array(116094) := x"2548";block_ram_array(116096) := x"0018";block_ram_array(116098) := x"a157";block_ram_array(116100) := x"fff2";block_ram_array(116102) := x"8842";block_ram_array(116104) := x"ffe4";block_ram_array(116106) := x"f62c";block_ram_array(116108) := x"000f";block_ram_array(116110) := x"a04e";block_ram_array(116112) := x"0018";block_ram_array(116114) := x"b3bc";block_ram_array(116116) := x"fff2";block_ram_array(116118) := x"b051";block_ram_array(116120) := x"ffe4";block_ram_array(116122) := x"ba3c";block_ram_array(116124) := x"000f";block_ram_array(116126) := x"1878";block_ram_array(116128) := x"0018";block_ram_array(116130) := x"c93a";block_ram_array(116132) := x"fff3";block_ram_array(116134) := x"2e8c";block_ram_array(116136) := x"ffe4";block_ram_array(116138) := x"c45c";block_ram_array(116140) := x"000e";block_ram_array(116142) := x"6154";block_ram_array(116144) := x"0018";block_ram_array(116146) := x"72c7";block_ram_array(116148) := x"fff3";block_ram_array(116150) := x"7598";block_ram_array(116152) := x"ffe4";block_ram_array(116154) := x"a0b5";block_ram_array(116156) := x"000e";block_ram_array(116158) := x"3ddc";block_ram_array(116160) := x"0018";block_ram_array(116162) := x"af2b";block_ram_array(116164) := x"fff3";block_ram_array(116166) := x"de13";block_ram_array(116168) := x"ffe4";block_ram_array(116170) := x"8f7c";block_ram_array(116172) := x"000d";block_ram_array(116174) := x"aade";block_ram_array(116176) := x"0018";block_ram_array(116178) := x"b64b";block_ram_array(116180) := x"fff4";block_ram_array(116182) := x"33ab";block_ram_array(116184) := x"ffe4";block_ram_array(116186) := x"47c0";block_ram_array(116188) := x"000d";block_ram_array(116190) := x"0204";block_ram_array(116192) := x"0018";block_ram_array(116194) := x"59ea";block_ram_array(116196) := x"fff4";block_ram_array(116198) := x"fff7";block_ram_array(116200) := x"ffe4";block_ram_array(116202) := x"abdd";block_ram_array(116204) := x"000c";block_ram_array(116206) := x"efb3";block_ram_array(116208) := x"0018";block_ram_array(116210) := x"9642";block_ram_array(116212) := x"fff5";block_ram_array(116214) := x"20f3";block_ram_array(116216) := x"ffe4";block_ram_array(116218) := x"9f2f";block_ram_array(116220) := x"000c";block_ram_array(116222) := x"6c67";block_ram_array(116224) := x"0018";block_ram_array(116226) := x"9794";block_ram_array(116228) := x"fff5";block_ram_array(116230) := x"674e";block_ram_array(116232) := x"ffe4";block_ram_array(116234) := x"8e43";block_ram_array(116236) := x"000b";block_ram_array(116238) := x"f6b6";block_ram_array(116240) := x"0018";block_ram_array(116242) := x"8c48";block_ram_array(116244) := x"fff5";block_ram_array(116246) := x"a7ab";block_ram_array(116248) := x"ffe4";block_ram_array(116250) := x"52bf";block_ram_array(116252) := x"000b";block_ram_array(116254) := x"8b6a";block_ram_array(116256) := x"0018";block_ram_array(116258) := x"610a";block_ram_array(116260) := x"fff6";block_ram_array(116262) := x"240c";block_ram_array(116264) := x"ffe4";block_ram_array(116266) := x"3318";block_ram_array(116268) := x"000b";block_ram_array(116270) := x"9168";block_ram_array(116272) := x"0019";block_ram_array(116274) := x"037f";block_ram_array(116276) := x"fff6";block_ram_array(116278) := x"ceca";block_ram_array(116280) := x"ffe4";block_ram_array(116282) := x"8fc8";block_ram_array(116284) := x"000a";block_ram_array(116286) := x"8ebd";block_ram_array(116288) := x"0018";block_ram_array(116290) := x"a0fe";block_ram_array(116292) := x"fff6";block_ram_array(116294) := x"d14f";block_ram_array(116296) := x"ffe4";block_ram_array(116298) := x"435c";block_ram_array(116300) := x"000a";block_ram_array(116302) := x"5948";block_ram_array(116304) := x"0018";block_ram_array(116306) := x"c446";block_ram_array(116308) := x"fff7";block_ram_array(116310) := x"64b9";block_ram_array(116312) := x"ffe4";block_ram_array(116314) := x"6a66";block_ram_array(116316) := x"0009";block_ram_array(116318) := x"e11a";block_ram_array(116320) := x"0018";block_ram_array(116322) := x"f2f9";block_ram_array(
116324) := x"fff7";block_ram_array(116326) := x"a2ee";block_ram_array(116328) := x"ffe4";block_ram_array(116330) := x"6261";block_ram_array(116332) := x"0008";block_ram_array(116334) := x"f4d3";block_ram_array(116336) := x"0018";block_ram_array(116338) := x"499d";block_ram_array(116340) := x"fff7";block_ram_array(116342) := x"de31";block_ram_array(116344) := x"ffe4";block_ram_array(116346) := x"2401";block_ram_array(116348) := x"0008";block_ram_array(116350) := x"fe7b";block_ram_array(116352) := x"0018";block_ram_array(116354) := x"51b6";block_ram_array(116356) := x"fff8";block_ram_array(116358) := x"6ae0";block_ram_array(116360) := x"ffe4";block_ram_array(116362) := x"2064";block_ram_array(116364) := x"0008";block_ram_array(116366) := x"c8a4";block_ram_array(116368) := x"0018";block_ram_array(116370) := x"5cf8";block_ram_array(116372) := x"fff9";block_ram_array(116374) := x"02c5";block_ram_array(116376) := x"ffe4";block_ram_array(116378) := x"757a";block_ram_array(116380) := x"0008";block_ram_array(116382) := x"aebd";block_ram_array(116384) := x"0018";block_ram_array(116386) := x"ecab";block_ram_array(116388) := x"fff9";block_ram_array(116390) := x"1b04";block_ram_array(116392) := x"ffe4";block_ram_array(116394) := x"530e";block_ram_array(116396) := x"0007";block_ram_array(116398) := x"9997";block_ram_array(116400) := x"0018";block_ram_array(116402) := x"237e";block_ram_array(116404) := x"fff9";block_ram_array(116406) := x"95dc";block_ram_array(116408) := x"ffe4";block_ram_array(116410) := x"953a";block_ram_array(116412) := x"0008";block_ram_array(116414) := x"1a70";block_ram_array(116416) := x"0019";block_ram_array(116418) := x"0e3c";block_ram_array(116420) := x"fff9";block_ram_array(116422) := x"93c1";block_ram_array(116424) := x"ffe4";block_ram_array(116426) := x"4b2b";block_ram_array(116428) := x"0006";block_ram_array(116430) := x"ef5d";block_ram_array(116432) := x"0018";block_ram_array(116434) := x"803d";block_ram_array(116436) := x"fffa";block_ram_array(116438) := x"05c3";block_ram_array(116440) := x"ffe4";block_ram_array(116442) := x"2e5d";block_ram_array(116444) := x"0006";block_ram_array(116446) := x"ea1f";block_ram_array(116448) := x"0018";block_ram_array(116450) := x"bdac";block_ram_array(116452) := x"fffa";block_ram_array(116454) := x"ae5c";block_ram_array(116456) := x"ffe4";block_ram_array(116458) := x"a409";block_ram_array(116460) := x"0006";block_ram_array(116462) := x"6976";block_ram_array(116464) := x"0018";block_ram_array(116466) := x"c32f";block_ram_array(116468) := x"fffa";block_ram_array(116470) := x"9a5a";block_ram_array(116472) := x"ffe4";block_ram_array(116474) := x"7beb";block_ram_array(116476) := x"0005";block_ram_array(116478) := x"e6d8";block_ram_array(116480) := x"0018";block_ram_array(116482) := x"995b";block_ram_array(116484) := x"fffa";block_ram_array(116486) := x"cabc";block_ram_array(116488) := x"ffe4";block_ram_array(116490) := x"3146";block_ram_array(116492) := x"0005";block_ram_array(116494) := x"b004";block_ram_array(116496) := x"0018";block_ram_array(116498) := x"cb2c";block_ram_array(116500) := x"fffb";block_ram_array(116502) := x"6182";block_ram_array(116504) := x"ffe4";block_ram_array(116506) := x"5197";block_ram_array(116508) := x"0005";block_ram_array(116510) := x"10f2";block_ram_array(116512) := x"0018";block_ram_array(116514) := x"88de";block_ram_array(116516) := x"fffb";block_ram_array(116518) := x"ca6e";block_ram_array(116520) := x"ffe4";block_ram_array(116522) := x"b081";block_ram_array(116524) := x"0004";block_ram_array(116526) := x"ebaa";block_ram_array(116528) := x"0018";block_ram_array(116530) := x"bd84";block_ram_array(116532) := x"fffb";block_ram_array(116534) := x"7a04";block_ram_array(116536) := x"ffe3";block_ram_array(116538) := x"f416";block_ram_array(116540) := x"0004";block_ram_array(116542) := x"55a7";block_ram_array(116544) := x"0018";block_ram_array(116546) := x"8615";block_ram_array(116548) := x"fffc";block_ram_array(116550) := x"713d";block_ram_array(116552) := x"ffe4";block_ram_array(116554) := x"729c";block_ram_array(116556) := x"0004";block_ram_array(
116558) := x"26f8";block_ram_array(116560) := x"0018";block_ram_array(116562) := x"adfb";block_ram_array(116564) := x"fffc";block_ram_array(116566) := x"5d69";block_ram_array(116568) := x"ffe4";block_ram_array(116570) := x"1ecd";block_ram_array(116572) := x"0003";block_ram_array(116574) := x"a215";block_ram_array(116576) := x"0018";block_ram_array(116578) := x"84bd";block_ram_array(116580) := x"fffc";block_ram_array(116582) := x"e3da";block_ram_array(116584) := x"ffe4";block_ram_array(116586) := x"25fc";block_ram_array(116588) := x"0003";block_ram_array(116590) := x"6e9f";block_ram_array(116592) := x"0018";block_ram_array(116594) := x"ab1e";block_ram_array(116596) := x"fffd";block_ram_array(116598) := x"59e6";block_ram_array(116600) := x"ffe4";block_ram_array(116602) := x"625a";block_ram_array(116604) := x"0002";block_ram_array(116606) := x"fc84";block_ram_array(116608) := x"0018";block_ram_array(116610) := x"b9d3";block_ram_array(116612) := x"fffd";block_ram_array(116614) := x"788c";block_ram_array(116616) := x"ffe4";block_ram_array(116618) := x"5d34";block_ram_array(116620) := x"0002";block_ram_array(116622) := x"7344";block_ram_array(116624) := x"0018";block_ram_array(116626) := x"9cb2";block_ram_array(116628) := x"fffd";block_ram_array(116630) := x"9110";block_ram_array(116632) := x"ffe3";block_ram_array(116634) := x"f8b8";block_ram_array(116636) := x"0001";block_ram_array(116638) := x"f74e";block_ram_array(116640) := x"0018";block_ram_array(116642) := x"4a38";block_ram_array(116644) := x"fffe";block_ram_array(116646) := x"49e9";block_ram_array(116648) := x"ffe4";block_ram_array(116650) := x"3e20";block_ram_array(116652) := x"0001";block_ram_array(116654) := x"e6d8";block_ram_array(116656) := x"0018";block_ram_array(116658) := x"6912";block_ram_array(116660) := x"fffe";block_ram_array(116662) := x"8dbc";block_ram_array(116664) := x"ffe4";block_ram_array(116666) := x"7078";block_ram_array(116668) := x"0001";block_ram_array(116670) := x"83e8";block_ram_array(116672) := x"0018";block_ram_array(116674) := x"5068";block_ram_array(116676) := x"fffe";block_ram_array(116678) := x"7528";block_ram_array(116680) := x"ffe3";block_ram_array(116682) := x"ec90";block_ram_array(116684) := x"0001";block_ram_array(116686) := x"5490";block_ram_array(116688) := x"0018";block_ram_array(116690) := x"67f0";block_ram_array(116692) := x"ffff";block_ram_array(116694) := x"384c";block_ram_array(116696) := x"ffe4";block_ram_array(116698) := x"2902";block_ram_array(116700) := x"0001";block_ram_array(116702) := x"1b4c";block_ram_array(116704) := x"0018";block_ram_array(116706) := x"c41b";block_ram_array(116708) := x"ffff";block_ram_array(116710) := x"829a";block_ram_array(116712) := x"ffe4";block_ram_array(116714) := x"2cdb";block_ram_array(116716) := x"0000";block_ram_array(116718) := x"4798";block_ram_array(116720) := x"0018";block_ram_array(116722) := x"5348";block_ram_array(116724) := x"ffff";block_ram_array(116726) := x"f950";block_ram_array(116728) := x"ffe4";block_ram_array(116730) := x"817c";block_ram_array(116732) := x"0000";block_ram_array(116734) := x"3d8a";block_ram_array(116736) := x"0018";block_ram_array(116738) := x"8200";block_ram_array(116740) := x"0000";block_ram_array(116742) := x"0000";block_ram_array(116744) := x"ffe4";block_ram_array(116746) := x"817c";block_ram_array(116748) := x"ffff";block_ram_array(116750) := x"c276";block_ram_array(116752) := x"0018";block_ram_array(116754) := x"5348";block_ram_array(116756) := x"0000";block_ram_array(116758) := x"06b0";block_ram_array(116760) := x"ffe4";block_ram_array(116762) := x"2cdb";block_ram_array(116764) := x"ffff";block_ram_array(116766) := x"b868";block_ram_array(116768) := x"0018";block_ram_array(116770) := x"c41b";block_ram_array(116772) := x"0000";block_ram_array(116774) := x"7d66";block_ram_array(116776) := x"ffe4";block_ram_array(116778) := x"2902";block_ram_array(116780) := x"fffe";block_ram_array(116782) := x"e4b4";block_ram_array(116784) := x"0018";block_ram_array(116786) := x"67f0";block_ram_array(116788) := x"0000";block_ram_array(116790) := x"c7b4";block_ram_array(
116792) := x"ffe3";block_ram_array(116794) := x"ec90";block_ram_array(116796) := x"fffe";block_ram_array(116798) := x"ab70";block_ram_array(116800) := x"0018";block_ram_array(116802) := x"5068";block_ram_array(116804) := x"0001";block_ram_array(116806) := x"8ad8";block_ram_array(116808) := x"ffe4";block_ram_array(116810) := x"7078";block_ram_array(116812) := x"fffe";block_ram_array(116814) := x"7c18";block_ram_array(116816) := x"0018";block_ram_array(116818) := x"6912";block_ram_array(116820) := x"0001";block_ram_array(116822) := x"7244";block_ram_array(116824) := x"ffe4";block_ram_array(116826) := x"3e20";block_ram_array(116828) := x"fffe";block_ram_array(116830) := x"1928";block_ram_array(116832) := x"0018";block_ram_array(116834) := x"4a38";block_ram_array(116836) := x"0001";block_ram_array(116838) := x"b617";block_ram_array(116840) := x"ffe3";block_ram_array(116842) := x"f8b8";block_ram_array(116844) := x"fffe";block_ram_array(116846) := x"08b2";block_ram_array(116848) := x"0018";block_ram_array(116850) := x"9cb2";block_ram_array(116852) := x"0002";block_ram_array(116854) := x"6ef0";block_ram_array(116856) := x"ffe4";block_ram_array(116858) := x"5d34";block_ram_array(116860) := x"fffd";block_ram_array(116862) := x"8cbc";block_ram_array(116864) := x"0018";block_ram_array(116866) := x"b9d3";block_ram_array(116868) := x"0002";block_ram_array(116870) := x"8774";block_ram_array(116872) := x"ffe4";block_ram_array(116874) := x"625a";block_ram_array(116876) := x"fffd";block_ram_array(116878) := x"037c";block_ram_array(116880) := x"0018";block_ram_array(116882) := x"ab1e";block_ram_array(116884) := x"0002";block_ram_array(116886) := x"a61a";block_ram_array(116888) := x"ffe4";block_ram_array(116890) := x"25fc";block_ram_array(116892) := x"fffc";block_ram_array(116894) := x"9161";block_ram_array(116896) := x"0018";block_ram_array(116898) := x"84bd";block_ram_array(116900) := x"0003";block_ram_array(116902) := x"1c26";block_ram_array(116904) := x"ffe4";block_ram_array(116906) := x"1ecd";block_ram_array(116908) := x"fffc";block_ram_array(116910) := x"5deb";block_ram_array(116912) := x"0018";block_ram_array(116914) := x"adfb";block_ram_array(116916) := x"0003";block_ram_array(116918) := x"a297";block_ram_array(116920) := x"ffe4";block_ram_array(116922) := x"729c";block_ram_array(116924) := x"fffb";block_ram_array(116926) := x"d908";block_ram_array(116928) := x"0018";block_ram_array(116930) := x"8615";block_ram_array(116932) := x"0003";block_ram_array(116934) := x"8ec3";block_ram_array(116936) := x"ffe3";block_ram_array(116938) := x"f416";block_ram_array(116940) := x"fffb";block_ram_array(116942) := x"aa59";block_ram_array(116944) := x"0018";block_ram_array(116946) := x"bd84";block_ram_array(116948) := x"0004";block_ram_array(116950) := x"85fc";block_ram_array(116952) := x"ffe4";block_ram_array(116954) := x"b081";block_ram_array(116956) := x"fffb";block_ram_array(116958) := x"1456";block_ram_array(116960) := x"0018";block_ram_array(116962) := x"88de";block_ram_array(116964) := x"0004";block_ram_array(116966) := x"3592";block_ram_array(116968) := x"ffe4";block_ram_array(116970) := x"5197";block_ram_array(116972) := x"fffa";block_ram_array(116974) := x"ef0e";block_ram_array(116976) := x"0018";block_ram_array(116978) := x"cb2c";block_ram_array(116980) := x"0004";block_ram_array(116982) := x"9e7e";block_ram_array(116984) := x"ffe4";block_ram_array(116986) := x"3146";block_ram_array(116988) := x"fffa";block_ram_array(116990) := x"4ffc";block_ram_array(116992) := x"0018";block_ram_array(116994) := x"995b";block_ram_array(116996) := x"0005";block_ram_array(116998) := x"3544";block_ram_array(117000) := x"ffe4";block_ram_array(117002) := x"7beb";block_ram_array(117004) := x"fffa";block_ram_array(117006) := x"1928";block_ram_array(117008) := x"0018";block_ram_array(117010) := x"c32f";block_ram_array(117012) := x"0005";block_ram_array(117014) := x"65a6";block_ram_array(117016) := x"ffe4";block_ram_array(117018) := x"a409";block_ram_array(117020) := x"fff9";block_ram_array(117022) := x"968a";block_ram_array(117024) := x"0018";block_ram_array(
117026) := x"bdac";block_ram_array(117028) := x"0005";block_ram_array(117030) := x"51a4";block_ram_array(117032) := x"ffe4";block_ram_array(117034) := x"2e5d";block_ram_array(117036) := x"fff9";block_ram_array(117038) := x"15e1";block_ram_array(117040) := x"0018";block_ram_array(117042) := x"803d";block_ram_array(117044) := x"0005";block_ram_array(117046) := x"fa3d";block_ram_array(117048) := x"ffe4";block_ram_array(117050) := x"4b2b";block_ram_array(117052) := x"fff9";block_ram_array(117054) := x"10a3";block_ram_array(117056) := x"0019";block_ram_array(117058) := x"0e3c";block_ram_array(117060) := x"0006";block_ram_array(117062) := x"6c3f";block_ram_array(117064) := x"ffe4";block_ram_array(117066) := x"953a";block_ram_array(117068) := x"fff7";block_ram_array(117070) := x"e590";block_ram_array(117072) := x"0018";block_ram_array(117074) := x"237e";block_ram_array(117076) := x"0006";block_ram_array(117078) := x"6a24";block_ram_array(117080) := x"ffe4";block_ram_array(117082) := x"530e";block_ram_array(117084) := x"fff8";block_ram_array(117086) := x"6669";block_ram_array(117088) := x"0018";block_ram_array(117090) := x"ecab";block_ram_array(117092) := x"0006";block_ram_array(117094) := x"e4fc";block_ram_array(117096) := x"ffe4";block_ram_array(117098) := x"757a";block_ram_array(117100) := x"fff7";block_ram_array(117102) := x"5143";block_ram_array(117104) := x"0018";block_ram_array(117106) := x"5cf8";block_ram_array(117108) := x"0006";block_ram_array(117110) := x"fd3b";block_ram_array(117112) := x"ffe4";block_ram_array(117114) := x"2064";block_ram_array(117116) := x"fff7";block_ram_array(117118) := x"375c";block_ram_array(117120) := x"0018";block_ram_array(117122) := x"51b6";block_ram_array(117124) := x"0007";block_ram_array(117126) := x"9520";block_ram_array(117128) := x"ffe4";block_ram_array(117130) := x"2401";block_ram_array(117132) := x"fff7";block_ram_array(117134) := x"0185";block_ram_array(117136) := x"0018";block_ram_array(117138) := x"499d";block_ram_array(117140) := x"0008";block_ram_array(117142) := x"21cf";block_ram_array(117144) := x"ffe4";block_ram_array(117146) := x"6261";block_ram_array(117148) := x"fff7";block_ram_array(117150) := x"0b2d";block_ram_array(117152) := x"0018";block_ram_array(117154) := x"f2f9";block_ram_array(117156) := x"0008";block_ram_array(117158) := x"5d12";block_ram_array(117160) := x"ffe4";block_ram_array(117162) := x"6a66";block_ram_array(117164) := x"fff6";block_ram_array(117166) := x"1ee6";block_ram_array(117168) := x"0018";block_ram_array(117170) := x"c446";block_ram_array(117172) := x"0008";block_ram_array(117174) := x"9b47";block_ram_array(117176) := x"ffe4";block_ram_array(117178) := x"435c";block_ram_array(117180) := x"fff5";block_ram_array(117182) := x"a6b8";block_ram_array(117184) := x"0018";block_ram_array(117186) := x"a0fe";block_ram_array(117188) := x"0009";block_ram_array(117190) := x"2eb1";block_ram_array(117192) := x"ffe4";block_ram_array(117194) := x"8fc8";block_ram_array(117196) := x"fff5";block_ram_array(117198) := x"7143";block_ram_array(117200) := x"0019";block_ram_array(117202) := x"037f";block_ram_array(117204) := x"0009";block_ram_array(117206) := x"3136";block_ram_array(117208) := x"ffe4";block_ram_array(117210) := x"3318";block_ram_array(117212) := x"fff4";block_ram_array(117214) := x"6e98";block_ram_array(117216) := x"0018";block_ram_array(117218) := x"610a";block_ram_array(117220) := x"0009";block_ram_array(117222) := x"dbf4";block_ram_array(117224) := x"ffe4";block_ram_array(117226) := x"52bf";block_ram_array(117228) := x"fff4";block_ram_array(117230) := x"7496";block_ram_array(117232) := x"0018";block_ram_array(117234) := x"8c48";block_ram_array(117236) := x"000a";block_ram_array(117238) := x"5855";block_ram_array(117240) := x"ffe4";block_ram_array(117242) := x"8e43";block_ram_array(117244) := x"fff4";block_ram_array(117246) := x"094a";block_ram_array(117248) := x"0018";block_ram_array(117250) := x"9794";block_ram_array(117252) := x"000a";block_ram_array(117254) := x"98b2";block_ram_array(117256) := x"ffe4";block_ram_array(117258) := x"9f2f";block_ram_array(
117260) := x"fff3";block_ram_array(117262) := x"9399";block_ram_array(117264) := x"0018";block_ram_array(117266) := x"9642";block_ram_array(117268) := x"000a";block_ram_array(117270) := x"df0d";block_ram_array(117272) := x"ffe4";block_ram_array(117274) := x"abdd";block_ram_array(117276) := x"fff3";block_ram_array(117278) := x"104d";block_ram_array(117280) := x"0018";block_ram_array(117282) := x"59ea";block_ram_array(117284) := x"000b";block_ram_array(117286) := x"0009";block_ram_array(117288) := x"ffe4";block_ram_array(117290) := x"47c0";block_ram_array(117292) := x"fff2";block_ram_array(117294) := x"fdfc";block_ram_array(117296) := x"0018";block_ram_array(117298) := x"b64b";block_ram_array(117300) := x"000b";block_ram_array(117302) := x"cc55";block_ram_array(117304) := x"ffe4";block_ram_array(117306) := x"8f7c";block_ram_array(117308) := x"fff2";block_ram_array(117310) := x"5522";block_ram_array(117312) := x"0018";block_ram_array(117314) := x"af2b";block_ram_array(117316) := x"000c";block_ram_array(117318) := x"21ed";block_ram_array(117320) := x"ffe4";block_ram_array(117322) := x"a0b5";block_ram_array(117324) := x"fff1";block_ram_array(117326) := x"c224";block_ram_array(117328) := x"0018";block_ram_array(117330) := x"72c7";block_ram_array(117332) := x"000c";block_ram_array(117334) := x"8a68";block_ram_array(117336) := x"ffe4";block_ram_array(117338) := x"c45c";block_ram_array(117340) := x"fff1";block_ram_array(117342) := x"9eac";block_ram_array(117344) := x"0018";block_ram_array(117346) := x"c93a";block_ram_array(117348) := x"000c";block_ram_array(117350) := x"d174";block_ram_array(117352) := x"ffe4";block_ram_array(117354) := x"ba3c";block_ram_array(117356) := x"fff0";block_ram_array(117358) := x"e788";block_ram_array(117360) := x"0018";block_ram_array(117362) := x"b3bc";block_ram_array(117364) := x"000d";block_ram_array(117366) := x"4faf";block_ram_array(117368) := x"ffe4";block_ram_array(117370) := x"f62c";block_ram_array(117372) := x"fff0";block_ram_array(117374) := x"5fb2";block_ram_array(117376) := x"0018";block_ram_array(117378) := x"a157";block_ram_array(117380) := x"000d";block_ram_array(117382) := x"77be";block_ram_array(117384) := x"ffe4";block_ram_array(117386) := x"e1e2";block_ram_array(117388) := x"ffef";block_ram_array(117390) := x"dab8";block_ram_array(117392) := x"0018";block_ram_array(117394) := x"7c43";block_ram_array(117396) := x"000d";block_ram_array(117398) := x"c197";block_ram_array(117400) := x"ffe4";block_ram_array(117402) := x"a963";block_ram_array(117404) := x"ffef";block_ram_array(117406) := x"7e6f";block_ram_array(117408) := x"0018";block_ram_array(117410) := x"848d";block_ram_array(117412) := x"000e";block_ram_array(117414) := x"5de4";block_ram_array(117416) := x"ffe4";block_ram_array(117418) := x"b79e";block_ram_array(117420) := x"ffef";block_ram_array(117422) := x"0056";block_ram_array(117424) := x"0018";block_ram_array(117426) := x"7aeb";block_ram_array(117428) := x"000e";block_ram_array(117430) := x"ee4d";block_ram_array(117432) := x"ffe4";block_ram_array(117434) := x"fc9c";block_ram_array(117436) := x"ffee";block_ram_array(117438) := x"88f3";block_ram_array(117440) := x"0018";block_ram_array(117442) := x"6f56";block_ram_array(117444) := x"000f";block_ram_array(117446) := x"1ada";block_ram_array(117448) := x"ffe4";block_ram_array(117450) := x"ccad";block_ram_array(117452) := x"ffee";block_ram_array(117454) := x"20b3";block_ram_array(117456) := x"0018";block_ram_array(117458) := x"8383";block_ram_array(117460) := x"000f";block_ram_array(117462) := x"b4d3";block_ram_array(117464) := x"ffe4";block_ram_array(117466) := x"ef2c";block_ram_array(117468) := x"ffed";block_ram_array(117470) := x"8f2c";block_ram_array(117472) := x"0018";block_ram_array(117474) := x"7257";block_ram_array(117476) := x"0010";block_ram_array(117478) := x"2170";block_ram_array(117480) := x"ffe5";block_ram_array(117482) := x"0887";block_ram_array(117484) := x"ffed";block_ram_array(117486) := x"1542";block_ram_array(117488) := x"0018";block_ram_array(117490) := x"63b3";block_ram_array(117492) := x"0010";block_ram_array(
117494) := x"7b27";block_ram_array(117496) := x"ffe5";block_ram_array(117498) := x"0280";block_ram_array(117500) := x"ffec";block_ram_array(117502) := x"b81e";block_ram_array(117504) := x"0018";block_ram_array(117506) := x"9582";block_ram_array(117508) := x"0010";block_ram_array(117510) := x"e73e";block_ram_array(117512) := x"ffe4";block_ram_array(117514) := x"e945";block_ram_array(117516) := x"ffec";block_ram_array(117518) := x"07b6";block_ram_array(117520) := x"0018";block_ram_array(117522) := x"8224";block_ram_array(117524) := x"0011";block_ram_array(117526) := x"8e63";block_ram_array(117528) := x"ffe5";block_ram_array(117530) := x"1a53";block_ram_array(117532) := x"ffeb";block_ram_array(117534) := x"76d7";block_ram_array(117536) := x"0018";block_ram_array(117538) := x"68bf";block_ram_array(117540) := x"0011";block_ram_array(117542) := x"f9df";block_ram_array(117544) := x"ffe5";block_ram_array(117546) := x"2b2d";block_ram_array(117548) := x"ffeb";block_ram_array(117550) := x"030f";block_ram_array(117552) := x"0018";block_ram_array(117554) := x"73b4";block_ram_array(117556) := x"0012";block_ram_array(117558) := x"6f10";block_ram_array(117560) := x"ffe5";block_ram_array(117562) := x"3bb8";block_ram_array(117564) := x"ffea";block_ram_array(117566) := x"714f";block_ram_array(117568) := x"0018";block_ram_array(117570) := x"6f32";block_ram_array(117572) := x"0012";block_ram_array(117574) := x"e116";block_ram_array(117576) := x"ffe5";block_ram_array(117578) := x"3d6f";block_ram_array(117580) := x"ffe9";block_ram_array(117582) := x"e3cf";block_ram_array(117584) := x"0018";block_ram_array(117586) := x"6ddb";block_ram_array(117588) := x"0013";block_ram_array(117590) := x"6936";block_ram_array(117592) := x"ffe5";block_ram_array(117594) := x"4e73";block_ram_array(117596) := x"ffe9";block_ram_array(117598) := x"503d";block_ram_array(117600) := x"0018";block_ram_array(117602) := x"67e0";block_ram_array(117604) := x"0013";block_ram_array(117606) := x"f2d9";block_ram_array(117608) := x"ffe5";block_ram_array(117610) := x"71a8";block_ram_array(117612) := x"ffe8";block_ram_array(117614) := x"bc87";block_ram_array(117616) := x"0018";block_ram_array(117618) := x"5c36";block_ram_array(117620) := x"0014";block_ram_array(117622) := x"5e0f";block_ram_array(117624) := x"ffe5";block_ram_array(117626) := x"7174";block_ram_array(117628) := x"ffe8";block_ram_array(117630) := x"3860";block_ram_array(117632) := x"0018";block_ram_array(117634) := x"6d7c";block_ram_array(117636) := x"0014";block_ram_array(117638) := x"e365";block_ram_array(117640) := x"ffe5";block_ram_array(117642) := x"749c";block_ram_array(117644) := x"ffe7";block_ram_array(117646) := x"9318";block_ram_array(117648) := x"0018";block_ram_array(117650) := x"693d";block_ram_array(117652) := x"0015";block_ram_array(117654) := x"77bf";block_ram_array(117656) := x"ffe5";block_ram_array(117658) := x"84f2";block_ram_array(117660) := x"ffe6";block_ram_array(117662) := x"f44f";block_ram_array(117664) := x"0018";block_ram_array(117666) := x"6754";block_ram_array(117668) := x"0016";block_ram_array(117670) := x"0dd7";block_ram_array(117672) := x"ffe5";block_ram_array(117674) := x"a178";block_ram_array(117676) := x"ffe6";block_ram_array(117678) := x"509f";block_ram_array(117680) := x"0018";block_ram_array(117682) := x"619b";block_ram_array(117684) := x"0016";block_ram_array(117686) := x"955f";block_ram_array(117688) := x"ffe5";block_ram_array(117690) := x"ae3a";block_ram_array(117692) := x"ffe5";block_ram_array(117694) := x"ae1e";block_ram_array(117696) := x"0018";block_ram_array(117698) := x"5eea";block_ram_array(117700) := x"0017";block_ram_array(117702) := x"2c1e";block_ram_array(117704) := x"ffe5";block_ram_array(117706) := x"c4b1";block_ram_array(117708) := x"ffe5";block_ram_array(117710) := x"081f";block_ram_array(117712) := x"0018";block_ram_array(117714) := x"5ffc";block_ram_array(117716) := x"0017";block_ram_array(117718) := x"bb58";block_ram_array(117720) := x"ffe5";block_ram_array(117722) := x"caa8";block_ram_array(117724) := x"ffe4";block_ram_array(117726) := x"5716";block_ram_array(
117728) := x"0018";block_ram_array(117730) := x"5726";block_ram_array(117732) := x"0018";block_ram_array(117734) := x"65d0";block_ram_array(117736) := x"ffe5";block_ram_array(117738) := x"ea0a";block_ram_array(117740) := x"ffe3";block_ram_array(117742) := x"ae68";block_ram_array(117744) := x"0018";block_ram_array(117746) := x"5de8";block_ram_array(117748) := x"0019";block_ram_array(117750) := x"013a";block_ram_array(117752) := x"ffe6";block_ram_array(117754) := x"02b1";block_ram_array(117756) := x"ffe2";block_ram_array(117758) := x"ee6e";block_ram_array(117760) := x"0018";block_ram_array(117762) := x"4f00";block_ram_array(117764) := x"0019";block_ram_array(117766) := x"9700";block_ram_array(117768) := x"ffe5";block_ram_array(117770) := x"f8e7";block_ram_array(117772) := x"ffe2";block_ram_array(117774) := x"4422";block_ram_array(117776) := x"0018";block_ram_array(117778) := x"6704";block_ram_array(117780) := x"001a";block_ram_array(117782) := x"757e";block_ram_array(117784) := x"ffe6";block_ram_array(117786) := x"5572";block_ram_array(117788) := x"ffe1";block_ram_array(117790) := x"5730";block_ram_array(117792) := x"0018";block_ram_array(117794) := x"2a9e";block_ram_array(117796) := x"001a";block_ram_array(117798) := x"dd86";block_ram_array(117800) := x"ffe6";block_ram_array(117802) := x"37aa";block_ram_array(117804) := x"ffe0";block_ram_array(117806) := x"be76";block_ram_array(117808) := x"0018";block_ram_array(117810) := x"3244";block_ram_array(117812) := x"001b";block_ram_array(117814) := x"aa70";block_ram_array(117816) := x"ffe6";block_ram_array(117818) := x"4471";block_ram_array(117820) := x"ffe0";block_ram_array(117822) := x"02df";block_ram_array(117824) := x"0018";block_ram_array(117826) := x"42ae";block_ram_array(117828) := x"001c";block_ram_array(117830) := x"99aa";block_ram_array(117832) := x"ffe6";block_ram_array(117834) := x"b00a";block_ram_array(117836) := x"ffdf";block_ram_array(117838) := x"21be";block_ram_array(117840) := x"0018";block_ram_array(117842) := x"32db";block_ram_array(117844) := x"001d";block_ram_array(117846) := x"0b3f";block_ram_array(117848) := x"ffe6";block_ram_array(117850) := x"956c";block_ram_array(117852) := x"ffde";block_ram_array(117854) := x"441b";block_ram_array(117856) := x"0018";block_ram_array(117858) := x"098a";block_ram_array(117860) := x"001d";block_ram_array(117862) := x"fa66";block_ram_array(117864) := x"ffe6";block_ram_array(117866) := x"e3a8";block_ram_array(117868) := x"ffdd";block_ram_array(117870) := x"952d";block_ram_array(117872) := x"0018";block_ram_array(117874) := x"191e";block_ram_array(117876) := x"001e";block_ram_array(117878) := x"8f37";block_ram_array(117880) := x"ffe6";block_ram_array(117882) := x"d628";block_ram_array(117884) := x"ffdc";block_ram_array(117886) := x"bb10";block_ram_array(117888) := x"0018";block_ram_array(117890) := x"25ae";block_ram_array(117892) := x"001f";block_ram_array(117894) := x"7b45";block_ram_array(117896) := x"ffe6";block_ram_array(117898) := x"ff44";block_ram_array(117900) := x"ffdb";block_ram_array(117902) := x"b830";block_ram_array(117904) := x"0017";block_ram_array(117906) := x"ea82";block_ram_array(117908) := x"0020";block_ram_array(117910) := x"5e03";block_ram_array(117912) := x"ffe7";block_ram_array(117914) := x"3d3d";block_ram_array(117916) := x"ffdb";block_ram_array(117918) := x"1da0";block_ram_array(117920) := x"0018";block_ram_array(117922) := x"4494";block_ram_array(117924) := x"0021";block_ram_array(117926) := x"180f";block_ram_array(117928) := x"ffe7";block_ram_array(117930) := x"3772";block_ram_array(117932) := x"ffd9";block_ram_array(117934) := x"cf6f";block_ram_array(117936) := x"0017";block_ram_array(117938) := x"f943";block_ram_array(117940) := x"0022";block_ram_array(117942) := x"2917";block_ram_array(117944) := x"ffe7";block_ram_array(117946) := x"797b";block_ram_array(117948) := x"ffd8";block_ram_array(117950) := x"f79f";block_ram_array(117952) := x"0017";block_ram_array(117954) := x"f3b0";block_ram_array(117956) := x"0023";block_ram_array(117958) := x"175a";block_ram_array(117960) := x"ffe7";block_ram_array(
117962) := x"b1ae";block_ram_array(117964) := x"ffd8";block_ram_array(117966) := x"0686";block_ram_array(117968) := x"0018";block_ram_array(117970) := x"01f9";block_ram_array(117972) := x"0024";block_ram_array(117974) := x"043b";block_ram_array(117976) := x"ffe7";block_ram_array(117978) := x"d8b5";block_ram_array(117980) := x"ffd6";block_ram_array(117982) := x"e47e";block_ram_array(117984) := x"0017";block_ram_array(117986) := x"e0cd";block_ram_array(117988) := x"0025";block_ram_array(117990) := x"0cd4";block_ram_array(117992) := x"ffe8";block_ram_array(117994) := x"0c2e";block_ram_array(117996) := x"ffd5";block_ram_array(117998) := x"e703";block_ram_array(118000) := x"0017";block_ram_array(118002) := x"e92d";block_ram_array(118004) := x"0026";block_ram_array(118006) := x"1f83";block_ram_array(118008) := x"ffe8";block_ram_array(118010) := x"477c";block_ram_array(118012) := x"ffd4";block_ram_array(118014) := x"b7ec";block_ram_array(118016) := x"0017";block_ram_array(118018) := x"c9d0";block_ram_array(118020) := x"0027";block_ram_array(118022) := x"38c3";block_ram_array(118024) := x"ffe8";block_ram_array(118026) := x"83cf";block_ram_array(118028) := x"ffd3";block_ram_array(118030) := x"a3a0";block_ram_array(118032) := x"0017";block_ram_array(118034) := x"c98b";block_ram_array(118036) := x"0028";block_ram_array(118038) := x"5d0d";block_ram_array(118040) := x"ffe8";block_ram_array(118042) := x"bc68";block_ram_array(118044) := x"ffd2";block_ram_array(118046) := x"6f8e";block_ram_array(118048) := x"0017";block_ram_array(118050) := x"c7da";block_ram_array(118052) := x"0029";block_ram_array(118054) := x"9eac";block_ram_array(118056) := x"ffe9";block_ram_array(118058) := x"1053";block_ram_array(118060) := x"ffd1";block_ram_array(118062) := x"148e";block_ram_array(118064) := x"0017";block_ram_array(118066) := x"936f";block_ram_array(118068) := x"002a";block_ram_array(118070) := x"d486";block_ram_array(118072) := x"ffe9";block_ram_array(118074) := x"5069";block_ram_array(118076) := x"ffcf";block_ram_array(118078) := x"e012";block_ram_array(118080) := x"0017";block_ram_array(118082) := x"7b09";block_ram_array(118084) := x"002c";block_ram_array(118086) := x"29ea";block_ram_array(118088) := x"ffe9";block_ram_array(118090) := x"9531";block_ram_array(118092) := x"ffce";block_ram_array(118094) := x"9e98";block_ram_array(118096) := x"0017";block_ram_array(118098) := x"7799";block_ram_array(118100) := x"002d";block_ram_array(118102) := x"a044";block_ram_array(118104) := x"ffe9";block_ram_array(118106) := x"f0a8";block_ram_array(118108) := x"ffcd";block_ram_array(118110) := x"2c8f";block_ram_array(118112) := x"0017";block_ram_array(118114) := x"4baf";block_ram_array(118116) := x"002f";block_ram_array(118118) := x"2832";block_ram_array(118120) := x"ffea";block_ram_array(118122) := x"6670";block_ram_array(118124) := x"ffcb";block_ram_array(118126) := x"cd96";block_ram_array(118128) := x"0017";block_ram_array(118130) := x"334c";block_ram_array(118132) := x"0030";block_ram_array(118134) := x"a068";block_ram_array(118136) := x"ffea";block_ram_array(118138) := x"b413";block_ram_array(118140) := x"ffca";block_ram_array(118142) := x"55d3";block_ram_array(118144) := x"0017";block_ram_array(118146) := x"19b8";block_ram_array(118148) := x"0032";block_ram_array(118150) := x"62e8";block_ram_array(118152) := x"ffeb";block_ram_array(118154) := x"360c";block_ram_array(118156) := x"ffc8";block_ram_array(118158) := x"be8c";block_ram_array(118160) := x"0016";block_ram_array(118162) := x"df78";block_ram_array(118164) := x"0034";block_ram_array(118166) := x"1ef0";block_ram_array(118168) := x"ffeb";block_ram_array(118170) := x"a3c6";block_ram_array(118172) := x"ffc7";block_ram_array(118174) := x"356e";block_ram_array(118176) := x"0016";block_ram_array(118178) := x"b383";block_ram_array(118180) := x"0036";block_ram_array(118182) := x"1ca4";block_ram_array(118184) := x"ffec";block_ram_array(118186) := x"4131";block_ram_array(118188) := x"ffc5";block_ram_array(118190) := x"92dc";block_ram_array(118192) := x"0016";block_ram_array(118194) := x"7932";block_ram_array(
118196) := x"0038";block_ram_array(118198) := x"22c8";block_ram_array(118200) := x"ffec";block_ram_array(118202) := x"dd8c";block_ram_array(118204) := x"ffc3";block_ram_array(118206) := x"e6ad";block_ram_array(118208) := x"0016";block_ram_array(118210) := x"3243";block_ram_array(118212) := x"003a";block_ram_array(118214) := x"5848";block_ram_array(118216) := x"ffed";block_ram_array(118218) := x"85bb";block_ram_array(118220) := x"ffc2";block_ram_array(118222) := x"3a6a";block_ram_array(118224) := x"0015";block_ram_array(118226) := x"ee98";block_ram_array(118228) := x"003c";block_ram_array(118230) := x"d381";block_ram_array(118232) := x"ffee";block_ram_array(118234) := x"6142";block_ram_array(118236) := x"ffc0";block_ram_array(118238) := x"788f";block_ram_array(118240) := x"0015";block_ram_array(118242) := x"9297";block_ram_array(118244) := x"003f";block_ram_array(118246) := x"6f19";block_ram_array(118248) := x"ffef";block_ram_array(118250) := x"4432";block_ram_array(118252) := x"ffbe";block_ram_array(118254) := x"b779";block_ram_array(118256) := x"0015";block_ram_array(118258) := x"1ccf";block_ram_array(118260) := x"0042";block_ram_array(118262) := x"634a";block_ram_array(118264) := x"fff0";block_ram_array(118266) := x"4e6b";block_ram_array(118268) := x"ffbd";block_ram_array(118270) := x"0ef1";block_ram_array(118272) := x"0014";block_ram_array(118274) := x"a46b";block_ram_array(118276) := x"0045";block_ram_array(118278) := x"c6b2";block_ram_array(118280) := x"fff1";block_ram_array(118282) := x"9e6d";block_ram_array(118284) := x"ffbb";block_ram_array(118286) := x"6f40";block_ram_array(118288) := x"0014";block_ram_array(118290) := x"13cd";block_ram_array(118292) := x"0049";block_ram_array(118294) := x"af26";block_ram_array(118296) := x"fff3";block_ram_array(118298) := x"4499";block_ram_array(118300) := x"ffb9";block_ram_array(118302) := x"e442";block_ram_array(118304) := x"0013";block_ram_array(118306) := x"5d7d";block_ram_array(118308) := x"004e";block_ram_array(118310) := x"833c";block_ram_array(118312) := x"fff5";block_ram_array(118314) := x"df4e";block_ram_array(118316) := x"ffb8";block_ram_array(118318) := x"270b";block_ram_array(118320) := x"0011";block_ram_array(118322) := x"7bed";block_ram_array(118324) := x"0054";block_ram_array(118326) := x"625a";block_ram_array(118328) := x"fffa";block_ram_array(118330) := x"f3b9";block_ram_array(118332) := x"ffb6";block_ram_array(118334) := x"1b53";block_ram_array(118336) := x"0007";block_ram_array(118338) := x"daad";block_ram_array(118340) := x"0057";block_ram_array(118342) := x"0634";block_ram_array(118344) := x"fff4";block_ram_array(118346) := x"81d0";block_ram_array(118348) := x"ffc5";block_ram_array(118350) := x"3ec8";block_ram_array(118352) := x"000e";block_ram_array(118354) := x"256f";block_ram_array(118356) := x"007e";block_ram_array(118358) := x"10f9";block_ram_array(118360) := x"0034";block_ram_array(118362) := x"6e1e";block_ram_array(118364) := x"ffd8";block_ram_array(118366) := x"5b7e";block_ram_array(118368) := x"0035";block_ram_array(118370) := x"0041";block_ram_array(118372) := x"0050";block_ram_array(118374) := x"713b";block_ram_array(118376) := x"0040";block_ram_array(118378) := x"fe67";block_ram_array(118380) := x"ffb7";block_ram_array(118382) := x"f846";block_ram_array(118384) := x"0021";block_ram_array(118386) := x"fd49";block_ram_array(118388) := x"0008";block_ram_array(118390) := x"d297";block_ram_array(118392) := x"ffe1";block_ram_array(118394) := x"5fa9";block_ram_array(118396) := x"ffda";block_ram_array(118398) := x"c8b7";block_ram_array(118400) := x"0066";block_ram_array(118402) := x"ad43";block_ram_array(118404) := x"0059";block_ram_array(118406) := x"4cd0";block_ram_array(118408) := x"0013";block_ram_array(118410) := x"5964";block_ram_array(118412) := x"ff93";block_ram_array(118414) := x"8039";block_ram_array(118416) := x"003a";block_ram_array(118418) := x"4f03";block_ram_array(118420) := x"003d";block_ram_array(118422) := x"808e";block_ram_array(118424) := x"0003";block_ram_array(118426) := x"8b36";block_ram_array(118428) := x"ffcc";block_ram_array(
118430) := x"118d";block_ram_array(118432) := x"00b7";block_ram_array(118434) := x"cf1a";block_ram_array(118436) := x"0049";block_ram_array(118438) := x"22a3";block_ram_array(118440) := x"0030";block_ram_array(118442) := x"a615";block_ram_array(118444) := x"ff33";block_ram_array(118446) := x"6af0";block_ram_array(118448) := x"007b";block_ram_array(118450) := x"b6dd";block_ram_array(118452) := x"ffae";block_ram_array(118454) := x"f768";block_ram_array(118456) := x"ff0b";block_ram_array(118458) := x"1014";block_ram_array(118460) := x"fefc";block_ram_array(118462) := x"eb20";block_ram_array(118464) := x"006b";block_ram_array(118466) := x"713b";block_ram_array(118468) := x"00ef";block_ram_array(118470) := x"c7ac";block_ram_array(118472) := x"ffa6";block_ram_array(118474) := x"ddb7";block_ram_array(118476) := x"fe4d";block_ram_array(118478) := x"8e7c";block_ram_array(118480) := x"ff2d";block_ram_array(118482) := x"ebd6";block_ram_array(118484) := x"0132";block_ram_array(118486) := x"6154";block_ram_array(118488) := x"001b";block_ram_array(118490) := x"a8eb";block_ram_array(118492) := x"ff5d";block_ram_array(118494) := x"8fd1";block_ram_array(118496) := x"ffc5";block_ram_array(118498) := x"79ae";block_ram_array(118500) := x"014f";block_ram_array(118502) := x"43ac";block_ram_array(118504) := x"0095";block_ram_array(118506) := x"f2e1";block_ram_array(118508) := x"fecd";block_ram_array(118510) := x"8236";block_ram_array(118512) := x"fee5";block_ram_array(118514) := x"af70";block_ram_array(118516) := x"017a";block_ram_array(118518) := x"4c24";block_ram_array(118520) := x"01ec";block_ram_array(118522) := x"71ec";block_ram_array(118524) := x"ff79";block_ram_array(118526) := x"cad8";block_ram_array(118528) := x"fe77";block_ram_array(118530) := x"7f50";block_ram_array(118532) := x"ffae";block_ram_array(118534) := x"9eca";block_ram_array(118536) := x"00e0";block_ram_array(118538) := x"85de";block_ram_array(118540) := x"012e";block_ram_array(118542) := x"633c";block_ram_array(118544) := x"0097";block_ram_array(118546) := x"cec2";block_ram_array(118548) := x"ff7c";block_ram_array(118550) := x"912c";block_ram_array(118552) := x"ffe7";block_ram_array(118554) := x"2434";block_ram_array(118556) := x"ffa0";block_ram_array(118558) := x"ea23";block_ram_array(118560) := x"ffe8";block_ram_array(118562) := x"0eee";block_ram_array(118564) := x"0082";block_ram_array(118566) := x"78c8";block_ram_array(118568) := x"008e";block_ram_array(118570) := x"4df6";block_ram_array(118572) := x"ff9b";block_ram_array(118574) := x"48e6";block_ram_array(118576) := x"ff0e";block_ram_array(118578) := x"1764";block_ram_array(118580) := x"004c";block_ram_array(118582) := x"5e9d";block_ram_array(118584) := x"0098";block_ram_array(118586) := x"6818";block_ram_array(118588) := x"0196";block_ram_array(118590) := x"513c";block_ram_array(118592) := x"01d2";block_ram_array(118594) := x"46c0";block_ram_array(118596) := x"0075";block_ram_array(118598) := x"a0c3";block_ram_array(118600) := x"016e";block_ram_array(118602) := x"fc34";block_ram_array(118604) := x"ff1a";block_ram_array(118606) := x"6804";block_ram_array(118608) := x"0059";block_ram_array(118610) := x"d692";block_ram_array(118612) := x"fef7";block_ram_array(118614) := x"7794";block_ram_array(118616) := x"000e";block_ram_array(118618) := x"5bf2";block_ram_array(118620) := x"ffc3";block_ram_array(118622) := x"f4a7";block_ram_array(118624) := x"0069";block_ram_array(118626) := x"3b9a";block_ram_array(118628) := x"ff3c";block_ram_array(118630) := x"5954";block_ram_array(118632) := x"ff04";block_ram_array(118634) := x"5452";block_ram_array(118636) := x"00fb";block_ram_array(118638) := x"9726";block_ram_array(118640) := x"0366";block_ram_array(118642) := x"2bf0";block_ram_array(118644) := x"0071";block_ram_array(118646) := x"b6c6";block_ram_array(118648) := x"fea8";block_ram_array(118650) := x"009e";block_ram_array(118652) := x"fd8e";block_ram_array(118654) := x"cf9c";block_ram_array(118656) := x"01f4";block_ram_array(118658) := x"f0fc";block_ram_array(118660) := x"030b";block_ram_array(118662) := x"a3dc";block_ram_array(
118664) := x"0235";block_ram_array(118666) := x"b7b8";block_ram_array(118668) := x"fc21";block_ram_array(118670) := x"0890";block_ram_array(118672) := x"fee7";block_ram_array(118674) := x"8f66";block_ram_array(118676) := x"008b";block_ram_array(118678) := x"510c";block_ram_array(118680) := x"0143";block_ram_array(118682) := x"2fb6";block_ram_array(118684) := x"ffd2";block_ram_array(118686) := x"743a";block_ram_array(118688) := x"03cb";block_ram_array(118690) := x"17f0";block_ram_array(118692) := x"012e";block_ram_array(118694) := x"0178";block_ram_array(118696) := x"0217";block_ram_array(118698) := x"0c58";block_ram_array(118700) := x"fa17";block_ram_array(118702) := x"02e8";block_ram_array(118704) := x"008b";block_ram_array(118706) := x"f68a";block_ram_array(118708) := x"022f";block_ram_array(118710) := x"7684";block_ram_array(118712) := x"0743";block_ram_array(118714) := x"3e18";block_ram_array(118716) := x"f793";block_ram_array(118718) := x"7e60";block_ram_array(118720) := x"fa07";block_ram_array(118722) := x"0750";block_ram_array(118724) := x"fa33";block_ram_array(118726) := x"e8e8";block_ram_array(118728) := x"0182";block_ram_array(118730) := x"bf70";block_ram_array(118732) := x"fbd3";block_ram_array(118734) := x"58d8";block_ram_array(118736) := x"f77a";block_ram_array(118738) := x"f910";block_ram_array(118740) := x"fa1d";block_ram_array(118742) := x"6160";block_ram_array(118744) := x"fd57";block_ram_array(118746) := x"98b0";block_ram_array(118748) := x"03f5";block_ram_array(118750) := x"d4b4";block_ram_array(118752) := x"013a";block_ram_array(118754) := x"2068";block_ram_array(118756) := x"fdf5";block_ram_array(118758) := x"9a00";block_ram_array(118760) := x"ffad";block_ram_array(118762) := x"3d9b";block_ram_array(118764) := x"fa8d";block_ram_array(118766) := x"03a0";block_ram_array(118768) := x"f7d7";block_ram_array(118770) := x"c620";block_ram_array(118772) := x"fa48";block_ram_array(118774) := x"b4b0";block_ram_array(118776) := x"f92e";block_ram_array(118778) := x"0240";block_ram_array(118780) := x"03cb";block_ram_array(118782) := x"8278";
                
                fill_block_28 := '0';
                
                end if;
                
            end if;
            
            --~ s_readdata( 1 downto 0 ) <= s_address( 15 downto 0 );
            
            --~ s_readdata <= (others=>'0');
            --~ s_readdata( 3 downto 0 ) <= s_address( 3 downto 0 );
            
            s_readdata <= block_ram_array( to_integer( unsigned( s_address ) ) );
            
            if ( to_integer( unsigned( s_address ) ) = 118782 ) then
                
                fill_block_28 := '1';
                
            end if;
            
        end if;
        
    end if;
    
end process;

end Behavioral;
