-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
W6OPY6nOG3MvvZtAMeTbSUM6OYbufvO4iIkAQGRHBuoL51gnDstcV5NzXfssJRi3
y5k8569KrH9zBkLE4ateRW+eWo1Wcf9NIPJpHErhY+WEvb++86jqZqpylK1woUg3
2fezG8BNRDqAHPKtZpNqMdnXTxPzZzejl3riF+4f9UMvogpgwsVgqg==
--pragma protect end_key_block
--pragma protect digest_block
OJwuyl9lXlbaGkYWkbLcwbB6v40=
--pragma protect end_digest_block
--pragma protect data_block
Epav+FGuRCwS5TGdC3tiLUw46kXnJIAz+hc1G01I9/mxoUyzBFMRHfvV2bxKUvYS
LDlmOGZikWkwGUsEqGCLzY3FgR+mDe7YTfFKH38C2+rcK7yfNLoUaVZNCui8a+Pq
k6rnMsktI1hpjnWiPI/AIXk3C9dmdcwerKb8Kq8pfHyB0aA8U3fDLNI+yYg0By2L
NeBJzXGWsHdKNiHHqk7pPy0hNtd0r9AntFEOFV/vMkSGb3qMkM2nZ1/y2UiscOZU
ZVa3P3AwsDFRn2Bf2liWl5UjIaBglcurTqym1fgbIBtR7sNUqkEU1PZpvcX57fI3
qwPfSkHC2gfunRtOTenwvRY8/wWk4QFHODVhTDCv1awMWtEFFKKY7A2XJVPQGUCn
0lR/1xerrwQd9d+58ccGZ3NQS37uEJAL9juSitOlYwfvFsvtOEL3bBsJ3APbNZUw
tkxnrUmUlKy94A6FGHaCsgTFvzkgmUaYVE4lRQ98aVpA0yvULQ2LS4Rdm+8XRZm/
TYjHJUw//YiTYm1zuClsKNwTv8nVZpkTvNPgIKNPJi4xpNjfePVach0HCWK5kpJS
FatINscs2AfGSAZEBW+oWcshA6euqG3w7BzD+MaOlmEj228DYvajibSHpCeDtq2C
EkJL6np9thLcvVFC5Rj8R+XlzJimGUQKdAP0ZSgPaXIENbCQbB2K/6ketZaMXg2s
8qFsgec8IWM8Lf7pcRLfy+KSonJ83qjDhQMHwENre9P+g3t9fLZjbGIvfnQ3Ng4j
2M5IFmGNG0gfz0HJr2ReR4I8tGPfsqlMHVnaBUKvNjT4sswYqx2SwrVYOnzE56cb
K0a5+Fj4RBX6R8aQTH5tsMHTe5ggkaUyZlC5IfTtG8An5ETH1ocbi49dRLBzj/il
1gLnv3qWwWB1qhfRCxHk3wWR5lN1pUAIEac4Llw3kSuS/OwE0AXTs+jvLOODq6U9
fJF7Rq//4ItWkfW86bigveVR0abVQyAcv5hppqkKBQnNlLPMFOdhR840SkzQ9eD1
K482nDxxz+Ohp/fO6/m6+7kT1T6RDERl6CybxP91i7mMrhrmEb/7Ru7CWFHiYS1S
RCfGP2JZZ97zV3wxlcZ1fIN7MCuH8Xq5Ny2l9ySZKP88fKA6JNaW5xWspBktp7Dm
N/qfhZLONROKHAlowY8daGk5vFtkI8X4LtTNIY9EBW1I9Ycxo7qLXUWich5pj80f
ldMzbUpYqsx4bz0vUUhbme+TXIsbM1ZBiOBB3JAHZH0Dkm6JUtUi3qN3HOQdreTR
Z8S6x8uJrxZFEfFgidL3lyvzRt3JycYWsbVDGdfMNrZn41u2yloKMZeQHrjMaNCe
uz2OPrxgsLEzMCz8iTgDdVbacMxQzsTagBZuY2RPK85ljcpzxE6s85+9/E3HWmWS
hJ0HwaZ/eZn0uNlc8Ep+ZJU+apzdT/LAtg6/L02R8ztQfLUvz8j9jmLpi1Jbrryv
0BVl8N6HKYD6gdZohGjlCjIRb9972+6K/t66rpOAB57bbhw9cRoRekXJNpKkP0sS
acIjvb4NMWGzeBcsu3oItq+KEiLghMxEUs9dL2W9SRkrjIbS780HUF4ASmZ+YyC7
v/ZM3dbqFIwSHrc1FuvvdBYNTO3VdywngonVRGycE3jiSxcBUVU1LM+i8JtPAyAz
1iEfSc0Rmdk46HtZBE5m+EOAG3DTR5uwhXEPa0X8NiUxoPzZYPwJ+hAgN7nAALIA
Dg5TN/m65kjmNWcFYgwLz7vb1xrikyCEThuWIMnSjBKqtYKceXXVIFQpcTEYioWO
JQMbspuzuBDcmmbEBS6Fj6Sq23s32wbkw9ojYcDlN6xyVVbDKNVWF8oSyC4tWJ0u
72yO34TLiBUJWqU/zZ5Yfv12jqAW0bOClg1vCglejSxvHv2rAzEVvS5YBFzBRy/2
zm6eQ3yJrPwwpC4q26qvlWZUEJz5n9AZU4m5pIlRFcPT7qLwy4IC/TBFyf9eq6c5
tcqWteIdPJsOwBClhp9JfjUdmcDjfF1ylxv/9W1iUzBao+JRemWmdXFBw/ookrjQ
bMjV5bcb61tZkOmWVylzw3SHyYe1iLg9ydMbvIjJIMMXoNa/R7oDdDw+bAmmGU4h
UEY7yvouI+Vlt+oRhxBPyJLev/2Tni8IE6JDlnIDlKxMo1fI6tvY2BqGhiS+VWky
+yDJz3mW4CRkiJRQDucqucAYHOH7i0wpIARMTXIlyvI6NKjHUhQDBLJ19V9otFWF
aDYXOI/mmUyrd6HBw76EMZeqJkhU9oiKL32Jp1RMFw8FR4f/VwyV5fFy0+c3aKSd
eRaxHmzXObWQ+fUSGNKMQ/dxv7Pfzbnz56mFZGK+f3FnVzv2NlNF5g1I2O+jWosv
pDsOPV0Xie5UR8bxYfD4vsrWl89/lRzRS+nN+lLBMHnzg4AkRcCzEiE5AwSx6hdB
gobsgoWtMlXZAfHHyJaCcbawin7DDLJvEWm0W/k0i95EHfwrq954OgOEt4KR/ezB
TImOKf4T/erofXlNo/lZlo00Tr53ozNvdqY8U0tVUJ/QRNeH32VBEs9sTS/GgHQk
yQpbpTk4mWQgTSMsWQfb64G6cmb12zJDNb2f2OVRxrWlc5P+IdMzZiTVb8jL7ir+
YSw5/O1Mu5KxGsGpcJKmqbglv3K0cfoJFMgJCFXpEDnxfhXlh3ID+gM8LqF+dfnj
Zxvph9FLwcA015yoN4rYrzp9ybsI5V8Tq4dtY2Q/Y4rir/2MzkyS115qOs9ptRtF
8t9pKXCteDAT7wDH+AoVcc/2vLyME65LDvPwzFp5ZcramkNZQmXiqAjHzzc5npLe
2scWflGDT3PLsohCvkPXrkQhzWmCpdX/nPPxDIC29JjnapQPUlDtAOL3oI8WJS8F
vhZrS0cRw77w4VNrZziP7QNaDbRoasWEnVB6lqmvWLGhRFnmoentmcPiO0Achb/b
abmLXiEzt+6cqClx2wJ9ZKvySD5/rlxKIXW3DvKomBWWLnRQh7uVNofiJdawGniU
PhLT+vA288l/ZMlrBb6+QmZThMqjUtFe72NAoADWYZVsbYdyc1ouuvPhXuCZRfMv
m9bzcbGRb0955uDqj5h/YuT7XmD261NaSxmFJGX1GY8UNtxiQUIQX/eZSNGvLDEt
0eQq5lhJxFVCN36nvr4tXxKl5SWIea57YW06/fMC5QzdzsAiqZ7ddwmLOvCGAuy1
tEn79K5YuFodQB5p2eaeMousExRyexhl0We4jpOujxXClht4G//775L5dn/TBsFu
+Pwa19pOcT1WBHtkFqSAgIZ7bn9h/2nvDwX7cXV8w6EjyBESWUaiXtlsPuLBj9H1
k4Wpeo1JHfGfuXBLrSEo+9QsbAJMJ/u1s4deJoWDOUuMELdsXXPce6JW5FQVWJNY
8Xsj11fX9e8fzYWHSMdyLexrQJkGUtRcC9XHqknfKkrEPKkUtZt44oMf2IsOsZ+u
yIC8lfuuN50rho1edfqhIapLL9OQK9kfP4sQ8vyOYqC4Scx9CI8CNFdT8eoXalds
hta5Jkg6lywU97dKpDtsTWMYi0RNua5/L3aii7v2J7OsnONjzy8JeXkyqXqJpcz/
dE8kR0vwjGPKyBT7BG2KtSteoh9drqBvGe8bLMUvnkGx0sEG+AHX3SHnBcMJSbT9
CcsxY1q0lliNxh5TG8rV03ghaDsECFDUPV5FVfTErEjHd4ORN2z+EV5ue79p2MOG
AktF3uuvn7L4NJIo8REVi3B7H0RWQz4q+24/FzpPEpDw7kBfDsJrDyFwtYvuQ2SH
VPinrLj9fvKK47+vZhxZmeYrgooK1k8zEbjB3CuhLkVVeHhke0f/9jW9hMRp3NGA
SQs210b/DYLHTvWz5PWCs++CRMGxMwXAPtN3BbiyyDd920sE//wQxba0fWyg6Phu
zqOwm1DeiPJAu+srLEnaOiRTNQJRRHVPHS8pYn4qCBRU9lQQ+gDau+tatCVhuUfz
Cbi40cPDXody2E1wBq9yq7s+Y5OyXulO3puZF02fxE1JJKA7sUM55O4D5Yc8Upfi
jHyat2tNX0tiy28pfyAxVUZ+zPDWBRwQR9JT3ujKYtINyym5RIOoCVV1q38NBMiA
F+iVj2ft5SxMRN8/HBJYd7ux7s2qTzdL4QCrqpDK8lOx58kTs76If80U1ONmFQeH
YbUu3yqxG7xTR+/QPHtJlYAB2OfEu2Jgfso3MbKETCaQeZEauzHDJaXcfv2TH0Ig
F9VEur/Ck4xT1pwnJVUM+1p32lxW0d1Wl7CTg8JnNKD6RsnaS8PI2yVCohUHoceF
uqCMQ++wQn0hAWBfWHrI2PaEhpI9JdJJXIPao9uDJLdWD4zniMUo29nSfbgSr69M
LsHO3eFM0YqKxwm3z00jSrigP+cBw/Odi+/mXY/XnkWIIx/QBoprXaJD+KfmP/vT
793zLZVWM1o/VmtOottglTBGD5v1GAwrtObatl8BbtHuABfg3Asa0hRyuDG3rofw
DRWCYdYtkXfQhvF43b3LPuLChOxiEIMi2ahkafG/WUAKfvuiybBgJEBwqTPdmZnj
y2mL0aK22sKIIXFtrw16MVUUGreiFhn6j7ev+bx0PQOjCGIy/D0mCl42w1QhLZ/i
VWNTi2f1X9MpqtJlzHKjAQQXuRYljXWSMtDQPQTs7Zc5Uv3gROnbCgkr/jvP2Q4x
nUf4Vq9n4FmE7HPQaCjHgC+95kwckD0uz03xqEc1di3Qm9wPL95lohaUKcJ2yO5j
kipdc/pQpHgOy2+Y6RpN90EUs2rZUy37vgoqxxKiaDXIyELg4I7rc4J30ZWVDOwZ
majl8QttRb0ic1FGm90bkDKfXitjzMQDL0gSpKrzvQVmmAtLP7HaJeEWpdw1l2uU
Wt020hgv3fmIJ4jgw9Eo/jYYA9k75d0lTNZRUGrp7exBGJh+MJoFEaCY8mjOzU/L
j/OWDOyjrl2bbVtlpwEUhqt9CU4tO4iioOXWlecKOr8KIvopo9oZFqhUBRX3xxI/
WHsioKzg4+lCcoSN0fl9M7MTyXPLarwCwQkTDOMTaRYHL7lx015FgNOmGXoNTYaW
2yFuDtf5uCAwg5V/3I9c+VUdK5RDNp/DsJvLyqlEMXWTsocc2p39xkDFEM2dDTBl
pdZPmf0+S0jsLP+Qa0wWzrzqDKQUaZImyAReF9z6QJm/NFDvuT2aOfezPBdiBho1
g4Rlv/7wLmCgSL8eesmsw8mrwJ2Yin1y++z9rF0VFP6OEOdiBwZqyyUduSqpbDMh
VYYPlkfgDBvBwxYEbjkpdCI2rs/v3mZUS04hV+LoCuAM01guUhBFaJ6fTQFfCjdZ
s6UlTnrkvk5aVylJLsmsM8YBxfUe2VzkHCQh/f9Ms+jzp2egTYiGuSd4MzG8R19T
5lITuVxLyxSLvpp1dz/2CXaYoUKYysILbax6iF0mrKh5Ac+V5RonVe7wVbUtsFgQ
2AG4/nXm7r4TiEIvvm2XLtCXTFWwiyZ1WENAMpqYawTDLDNciFDdR0YE+miBFtJt
cNl+80y/rM3hs1l0JQM0drXGtBJtpoSZkIA5gV26KYhhBjgnGvhoDpynz4SB5q5M
hHDEC/0M7gQQEMikByvXlojcOy8elYS94aDzLvdFKw+KqGUqZ5sOPHg7XzXsg6na
iQuWm5pjtky45utm+NFgZcpOVDzph3hdjjtSggJ128AFUb4WYXsQxDF9rq5OJElI
ZHgqFNOl23YAKg2UA12MXLkxbCD47qmcYgrQwIMxzAVD1T2sHN/m+HisLtnqahcV
NAat5AIGm06nixBK7EKLtgB18OQae28xud+f5fhMVFf7i6qzk47B1QSQLHyeSu06
ragUKZhWsqwrcwlEsYO6EZtQLm8BX0PTc/suttqXGiDC+/NJz1frybE0tLB9jrew
rLhZ9rCmYBKjKq3L9wOnbcN/fdY2QllPnuKRQW5ZAKeYDjud3wTcxUaXMqJExiqT
cfZYqEtX9NTodO1VDyh4o+58Y6zu4duj5cUDe0yjibeHu8ud2Zw/rCLETugi020q
+aE5iYBC+NmG3SRhh3qpHOZC4pv3y3BxH47ip+O54UDiAXp+Lph2z/9uagJ0/2uA
lwMGs6TXUnRY8pDRpDWucD32/qDrROiFHq6Duw4jvLjM0h7XJE4o3luCbgvBqeXI
15m223Xwn4T8s8coq1BTBAqh/i+BXAk0AI2qkcR8uY+pphShzHFjnOdhb7POKHo8
+SrmAwe+6EoudMM/BWv1s+24Nq4afdXB5YvoxH+csAZ7BRxx2gcusv7t9d6JY8Ex
Byv+1IzR89ZIDOzkWnGQkA70dz13ZIeszZ/KauzTYlvczHDKxLvcOz50C49mZI6q
ztwULHY7+fN7guKkS9wg6sJ6qXCGiymINtB+cwhSx7zVc8e4txiDBdY9rPWaLLmj
b4iZpbGZhF+GvA545YLjSyIUaOUmEtGLk7dESBOG1g3h409Npirh4ABinGz4kWI8
xkEjBCleA2EQkwiHUzZhiNP19znmJ4aXANgu5ISpfw+jl/uUQSTQcMUTaEJBjQc2
bpCB10K/Pf3cW3tpkBEAXhmSFbSH68wuWG9kZlGmHSUlJIpdfyurPkAbXiKnrHXi
LYlGoG0bshbaZFCDYqYzsAczfmgDKNyxBpTe29OCuHMVrhBWoikykwC0BqZl/q3V
I5QlhlTaoEPLzyuW1Fs2CQM3LYIDw6VoqK3COLOHSxHO/V2AIyjldeQZZKNJuoBz
80vddlme1Aydl9xJOToJOD/eZHriJHZH0bjif37K10F7o4SanRMYvgIec10Tr2mL
r4GfbZtrENoSnJbWDhC8VXBLoemyYmnbTd75Ugo/htOC83yb7R1mM5ZBvf2NRUUH
P7a03ouHFIyRIOXG9FYIgy/I5Pl+ET9cSqEiHqgStn88+3FY+NWyXC8cdHsu4lwu
pJy98wa4HIlIOaJQFRzEEfzfdmRGSIzNecZmIepkfJQi4BnF5BYgzcMM0AXOwaGM
JLpBm+g2/uba3zICJJwu6o4la03e/CDMBbeU0oBh9R2aLN/OBikeKevXWQUEx6U7
2kazJrG9TchSHXnoHmcXxIQYGOuF/Iy8yVwcp7xsmTRycu/9ya7+oZ1bxzJzBODz
xAD0aiJlJPlxHJTwncIspmiYYub5rrSftpy6iBSgvwM=
--pragma protect end_data_block
--pragma protect digest_block
FYTrYnbUnVbvDap2y+kYmNU2vuM=
--pragma protect end_digest_block
--pragma protect end_protected
