-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
a7/153Is3mW4ZwzGSvLyQD/NiLTbI4H+d9oPy24MbYIPyor82ZV7vFmtjNMWPSX5
j7x9unbCa1cVk4fd8h8Qy+p5nsEAieGsIb2J8Rjj50jiiTdcT3H6d4SRX+ItXjQO
TMpC3lFD/+6hKXWtoZ1xLJzIsKfpKDK+J6txRLbDfSo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9248)
`protect data_block
iofhD4+ZHw2/0ofGhDaprraNafNzxBlbglebtUAqC3h5A5Whr3NLcT/DvCoVnAA4
3I2D1P4pHa0yzOMorPOjE9vBLeopMqd+F8L6NytlyreItSIaMkR8qYVJDBXutRsD
c5FCIpPw6CejfC8JmRNjHBD5ZLLik/FBYo7i9WwsPCw/UKxgacmlaiXszSZFbNCG
iUF9FUbMOWXg9RSv6Lkn5g4motvyQJRWAduoD/8Z3VpkmF8V0YIRnf5AuvxuaHNJ
wcF0T+2MbetRa+fokOL6Y/b+UTrE2svkSjKAb6f9k1d50g+mBq6MqpMN6DepQsPQ
XwkD5hmxfnSZx7OtY+UEIFxAZhhVd86dc/DCJUKG8OKd3NONmRyKdW0M4XM+Vdze
QplchXXoroXEc7LaJF4XZwTA2/vnXUcB4oibm5l0ihdNmXo9gqgm9mDI0UaB4bo9
mom+AFGy1gaJsQ2kF/dHHrgNkizJ/hrDtdswC3h/m4O8WECwi8BT+vNEuJbyWuUT
NaIrSKtA5jLRaH9ZXxYk/C5gRs+dhpW89cTKnbgj/ZwiTlmZrSiWOW1bfw6k8Bwa
AVLWUlKsKgcI/Eq1keMJB6pb6f10+DpwptJbBPmK9meSvMAn7Abu9FX4rFPMNiwJ
PUWZKBbSQSkra7zahQSYdUOXnbkJK9++2B+PSNDa5fvy954fyIjzZ38NerokzuJY
fANR2mQUUDwcWHPjj6cxJdQCAiXyU1r9VCXXbP9gdP38I+JaSEBEqoI6GLWImBCP
/1JWAmvG+JcU1eZIlS2H6Sr3FNmqKbkwQh2sfZD2btmrKlcQkUxCsgzm7cdLsVn7
IhV3mJnG9aK3G7Hz9kIZ/PHVmrB66QDgvyq2GmECFBmpXGyssv/wYFcOxNubxR0J
YVV1L8RsaEr9irdSgFl4xbrataNkXGky0SCkl0g0JaEbtrD/o03zEy3i2MuDm2C7
tb6cSsJbZol9jdNXd6sjM863wPmrNJfqZm2nFtKboQ/L2giZYKJoMYUBBZDWs0DN
LOzynPRHRWp+IMAiSh03kTnfTm0K0FIiksBPHFywOkKU0Te+DqhOlDRrlv1euWyX
lhsputlkbqiATzEVp0gBhFvfsEIMYoOTt/Mk6sZamiS2tXLoWvNvc7ggfwpgHebL
rcMCq3RiRRrq+EESX9NlBjy+poA1eEwIsE+A6+lB9olUqKK5MEAvpyhhX71f6WGt
TOGvA3RgLwYKer7rQeDdmzXYgtqavjYZINtWC3RRsRxpzEYDIHU2MEMU9I7FuZSd
zW6K6eGSsZUu/XJhT4HnbTJiJFqZ84OsjPv9Jvq8uBx0d0XoUq83LFYLb6PUX23V
YTmEpYfWogp3XP9R37gkdJNtATJUbCFaAjH4T2RaWYxJex5IP+sHoPg2X8klhoff
ah25Rp96Irra9K4Ug1Y4zZ0hprdg8oznVfXggwdlVheaB1JLNnuz1JYQRoVTdjy8
FtlglJoAyJOPbNTTpHjZpvuvMVOZaU1W7cGo+Byqr/0j/iN6nfRbvDNrav5UD4ut
OOr8/OwKD3S3UI8ddW4PGdHGcXCV5CQvnKtXJDPfo8duYficMVTl+0leVzwGSOeu
f/w5Hl2UnW90hPgfrms7R9fqyLSvzB1cSJIpgDSypodLNwZXzP/cZ9Qk8BJAa3/i
DmVrxtTBGdQKn/9mA/S0UWX+YL7l0tj3v3SvJXgf4owEyeeYPPMwm4kIk3txu0CL
IR4z604A7sG+kukAo3YDEXcTsOrZQPVnilEdCPricr5Z1cVmZEJJhjVodJpZxkX5
RparT1AZvuKLJD1bVziJoeB9yZPVBf3zEghKzDMDcQrWZ0FGZB6+rmpefygRceLV
gUxn9XrK9U7a/Qtt06btMr8wbXgtkNKZwuUX36wYsFkSTs7z8xLt0jAwsP4JQEls
eTPFrCDdG2LCWc1Cb8dbTWPr/iARL6JOsdgpsd5NqtZdOkm12Ya3Gd52o6VP/JwN
VU2TaEkHC74T7oyQ6pG9mfLikBXLIZMLZGKe3eH+vGf0UlpcczMNVOKRN7WcdkSV
uq5ckvXraIEsFqVomrj0JENGi9y2XVEjnPXOjaHKWnFHwU0Kzd4KohnEneQ9MCn1
m6B4xcENw9TsS1YDJBDkPICwlvhDtzNZPPyHr5mW1eSD05+AL6MkI2B2qrDEY8i8
mlVkc0v2sOUqUI8RVep/MdSsfs1Cf8GYuMUdB11HFiYTnYzxcK3MLPU76zE3OD/8
RniuCmeQp5FDSeNosD7/dd6EHjXaCbn7MEPclZIo0q32ofgvAVvcQSZAKl2hnNCG
ZkHAcwpqld/cAPdpR/IRYsCjNEKR7FxxhonZjXnLQkQgvrUeCLgajgSlQiN5X/qC
Pg5LLlmU+IOFyODKN9IitVbh3hvgeq7zkNp8RWry4o5pKoF1bPFyzSyJJiddPzLl
e1lx5jXiKpNVTip15fOIS+SHfKE3Ltps1Td+v0Zt8xrwsBGvt+APf/Fd6ISgjs1C
KJNl4Nwz+ufN9cWL15l17XG31oke1MdLNYeWwqFWjq2b2WI9legkEO7qyfDVefX1
pJGr8fTdz59p/rjXKG/efhI7y5SKtiRiaOr7MnHU45FitpsWGVb/P0ZHzHcFIqbw
6zKbr1HeDusRC0Lr/y5NNS6WzjqValssWFwu9s4FbfnsBxj1tazt1NNC+BBZioqS
JGwYGBj/AJNaXgmwlrnhuCidF6frwL1X82UvVo/MoQd4A0pgEI8IlUT4/Lt/7dXt
4iEnxODOj4lPF1zxOaBrMoI7CL2Cf7POkfNlGIN5Zc8IaEa1In73npTh/L47uOtN
fandaPaqecDM5kZRLTJr2qjHhqPgn3bepJpgqmNjJQrpyKU9UMOEn70fhqUx+Z3B
lJNWzRP6qlkRO1H8T7hh4BJnyuOyRwmkh13RQwZ0m5+MIt/JgzIRTWb7p7PgvgyK
6WWXGwPlhp/ZGrkdgklue/y8UN3ewrYzqG3iAy66r9Aoup4Vp1gYMeEhjqw5khKq
Uj0dIXSVrLdzi6ucHGUHTkLdJ/Y3/BIU4i22c1zOtXx6X+413gmQtHfYGrf5Pw+A
hW4g8R9g5vd1BAqqwirbTQf3RDaOOGEOttzemgbSumyZXyLevSV+IML2Gad0Rl62
PbO/UnRpXmXTpBlC+HFp2A3IyFlITTGuvG7mmbKDo71HfnEYij5GFy5W0EXmctfl
uwEDezczFos9hCTkQEaxmU9ICeQle0SGNAAiihOoHVwkmd6lmSN4qFm5Wc6leLor
38RR0qT2qb2BJIXGhkivQ9DIAVuga5+neLpkCRwK4+V/oTCm0KqjHrgRYcIy4rGO
MDT+Wh5gGD5RK75CpDBDbd/X15vR6gm5SA8q1EAiW+iyy2wFUsWccDvclCDKLv2H
XkwKmJLGQEA0/1Kb4dpbMXd6nuXW3WGx5NfASMOg8L+0uHerBAjx4VAsHzSxSUoP
AN3BIgOUtDvXP4SBdYHYlfgIk8+wrMzd6W2IhwIlM1zkUsuJqAKD02ZxmXBq5J29
LIF7UsAp09RQSegL2mRAjFKB+CSD1PyaQIZjNhVXEFzdERqfmT0mfOwgCPja+SI0
k4o7NP6tmPGqX0VcfLbIYpeR3MHvF3P3x6+Gcon6gOzRUldb5OY5E7jOUfURXVFK
O1OeuWhoODmKPHn6nELbp4U9m7zJPdy7N9qF6rcTaDnYPmtn7R9stFAkkAxQOkx9
X5hgHUsfvfrA0jiL/g2cfPUNsv3g0AabZYFvD79Tk8oNXqayo0Aii8CGZMskzujm
uFJbw99XaVgFYEOP4EcB4bhWl4WSJUoWDfdH4ahP5GhrYlBb89nSLgTD9YWyT0Wj
M39uUMVMtZ2p8zFnYfCKsVLORiv+bpkpGjUsRbNcr83qQMtd2OgP1YPRrw8d6JY0
gxbQfOTfUtbVjzObWrHvxVEC5x4N4d+Mp5gPM8CNcrFf3cmgjYi+4r5p9sNBkuCG
kAdfe6s25pAvBPCjv4rxrWN2mnuaGsezRZLxIk2VhgIz1/IjQLNfT3LcxJPKwEEt
arONPa7Zx8h9jipaYYGoAu7e72Mfp0eyhm5iSy4eFYlG8Ep9M1mMX12pXGEzqxrB
Kg6lhlYSUpxZOddrz61B7U2fDPNt73UctPwveDjr9n5h9dT/Mh2kXmPM30bZPi14
chwsy5WbqtYlXY5VTlTfvDCrOysqrzHi2zXWLGh4Yqmw9m6drjS40DJWNkWgAx4T
RzQ6dg9A6LpZwB3pf0bGHGxw61J/f1rkPh3nosv2P3bWSo0AySch8nanNrKX5bXO
V7n0r5zt2e62C6H5VhKwfMqiyK/tYJSFJztW/H/elNh963EnIi8aWJwlrddTCtW3
wr8L02/oWoLjwOybiTjTv9uMnU4ReXUmh3NzqFv6jjTvHGLYu/RRh/rOxOYmbEr6
GfwLy4T4legSGK0VgmTxr5EuPjmdDuwCiyjhgJSXR4QQ7yLdau4PAlHo5lZ9BCQL
u/+1a7LjoqJa2mhK+v13EokaHgA9F8l1eyvyRIwIHgsVLX9QtusYFQop1DoEZes7
TSHL/ugrfvCULq4GnPsS++Qw57SJGjDm4kT7uuq9muiWbCsJeSHiJYgeKp1BRQ/0
N6YMhyy/D/qay5rp5mYp7VFDOlT+836qfVtqUil4MgEOASu2LarDwSBZ6cJmiIsd
bLqtGs1T57MaDCcFqZEUHl1G0ra9evTbG1MLUr+bhEduRKCOYcV80dOgVmxa5LIG
irlkoV5WrdEY3keTZdyU2+jFrcwBwA02NeVT1b6llC/Ydobxp7PPjQWMkzD46ynd
TG1b/kOJpNzL/i6e3sW4KbnyN66DbExcx7+nTXWgESL4bL1jnAgSS6EljFIEXRAO
tzb3376kxyCsk7x87npIzDVmEfp4K80AZvXkyffNmsCKIttHRYGdC/c4V55BdPA2
B9R1UF7+J2LxeNgOL+fDRpj2EcG1mtfPvAWlt2pqCBHgS+RoqBoL/pp/T/uvntIw
lHKDosFAfgqrW3Jl7T944dlO3c0TdfBl6Rd2egIFHpbmyyCsLtRwEy52FsXC15tY
VFhF///RB05hgybiTnPM3nD8JZX/7vLp/l+5AbbiiHAA/nSObRYWqAskB7fi4NTm
Cwh/f53m98RIbTbln/uHda5UlwZT8MjW8rE2KuPfUUoS2qp8xuerQs+rWuUmiaRC
mQu8lv2A5QHmhVCEUlzWBdT4xU827gsvf+cx9e5OF/E8FGnTItKLehJ3JWwsHKJo
LPn0YaWqzHRmZaLWRpnhB0HwYTssi8azSrERDpPBlSg+PerH2LPmXscbXrzxeDde
OtER9yNAZ0fg8rWwJKKOVfKcjVioBbTyeLGEERomR2cJgAHSHwsmkfquZ/GYZVpQ
+NqzsJoqbYq1y2ToUoyrYVV+MPTAFTZSy7iYmLGIxpvsO/sdXmODOxp81qjiMG7N
7E2kCza100Ke8IsqrOJ56Mncet/AaQS+OB805JuFNjzlQ8p7qMhsccMieiNvcxF0
uSVBfOpQOFvfLDWedXNlZgRx1AEz8KDAjemAE9gsUw2WkMuS7Mae9+haUhejjfty
YJ2a/htDS++1xQ8PhyIwrmcO6Jb2EoybThXIdyCQrMjzQfpCKWKqMNghXMbHOAVo
80BKA+mHdJaFY7TUUr1AOVLnncSjz72kHXez+E45gLZThd1m01F/wlTQrRaVUERF
F6YhJT7WcP5aksdpAnAdQ8xwOtrsR5ijW0VRnVIF91Sn63rGpKxg8uW0lHwaQitP
RvjvV6eNPAk9zUIv9K1k2icRVltSXyESt0C7uuJIzsejgr8onmtLoEOX5a6U/xyl
lu3X1BN0l7s3QLk4MGgOLsWlQ6MTjP/fz5cOQHVdjJ6CQB6fmVgjWSnl+vksBo6s
m1lSvG6cFF6twjoglqNWCxM/8npDAE93qrW1fBr+zzzZQ5vDRN2GFjmj0lmxmnim
1C15eKLNkHaZIptoJki5UEVLfLjI6IYndOrqErfIXp/quC/drsOU/rXP4CaNBEqs
TMrsbwmJTKilJb8S2FPIHTYgXkh6fvE9Yj/3lIT1y2rpjwaGKtD1SexIZHuN0rF9
jV/m7ahICo4ktcT5mvnl+ammbdZq0V3gC58mXxO7oCrscnkz613fCmmMh7UcRXDU
rCACcHsoCpAAlzBRmpazpH9yD8QGlFOB3txK+Gwe0y3PzvH1ic/RmKj1hGV8acSY
eneipGL57Cif3XWrGuo13Xie/2U9SIqNp5GXi5PgB5UggpwVxRRqmcebUKrSLu2/
or0sDMur5Abex4WDjNaPT/Ck+glkDMNr8MHNZVE7/+pdAwZ7MtkqTjPjS3Y0rBBS
Tqc8+qh29hiBqhF8CL83Ch2PDImQsuZdIxiAP55JeZndfkK2PbsZX3Kl8/wpZhnN
RcUUDUoyMjGptR7A5QUlpOSKox6/vTxsjw4ceOjJszA5JTQyY4TBwjtpd5p/OPZY
uCidTk5vStCwQdidOLqYY+nkgNnwnfjgZ/XWza0ueNrYNN0UYiLlXPb39viArWF2
5A206PGlrOc5EJJTtWT3+Iw//GY35UFnT2A5i7/rcXw2CIIvKnQo6WiyQ68L8CKh
V/sIU7T/FQhYJrFwvmyDWBreTcw9PM1lWbLB2Ceyw8YmIM44lEerf85ySS0eFUor
+rtHzlKGMVJkEAAmh8/jLrx3+PKKIudrk7S6pXL2VakktLLcJlNWq6pnarUUME0g
q1Tey8g0kiSSQ2u6qx85jlgH+DhU9wYw7ur+RqgmRMOx9KtDZXgLcpzImm/N9rnf
dONRVSZevj2BLYXORUrs8NQdrW1a+r14r9IFka68L+Loqc2SEy6MzaoL0rWmB3S7
sksnR+X1Tt2F4QtZLM06FUTVAW6P7hZWr4hoDbcNB+dGIwFDr460p2NETRMv+MII
bzfIiEtuOutaHyo63RsdmnhFZgQp4bGHDwDE//JIMqZokP9hY8UuwqEcbVXAyWoT
EfHtcQ5DLRw8yuSHr13McG2S/LW26iJBpsXjt98KKGiY2cudR6oV8PCEureZoVdf
kdWBjjRZJmHby6WNidTYCYuFW9xXDxUUpTdQXBiHDH7oTXJnuPiOtf33C5tOw1bg
XOJ23j7K1zZUm7JR4FzVFtIBxA4JIq19ow91fVGiiheyT3R6jnIAl2+4rV89nPqi
ioC4a1UwaKer0AZXe0V2XlewXd5uTKmrmH9xv6lH4+U0cc0xQOILRZdeLHhWsPrQ
BcliQNTdooFRRu5iBcG0f0ligGZGJKoGthla1eTKgm0SHzga8mlyFaR+5UbJgwcf
/OZNqs5+/AfcwSMRGA4fAeWftJAeu8/duDerfl78IXA6To4z4MudHl5+vkHoxSEN
927zno8UVko3wuEeK/CudmB/2sbL4zNQbNoLj+KKmKXZKVdWqCJ2QUJIDqyZN9fv
iNprPlQPDpn0nUU9A8Y3IgRPXeVKlIWNGU2T5umO+RrpxVE3rNVt6mBrghN7fKmh
f9scrAsgRG2D2xhcTyMvSqImIk/cx/xmSAzOAicCrivRAZBZbNfgF/4NtrnkZ9Ik
uGXVxQ0768l3B5m+gbMUPF5OnfPAkHj4padgEvQNV5v8nKSzF2atSh4kCJYNsDWz
/1di5gr/wyUaIeXrwJ7TvaG+7+jkUQ8vXxGI2ZEFwcr56OQFt7CFY4l5AfehGb8c
cj19UXynfZqXGJvAiSPPH0ZQVqJ7fkg4RRVqSYNN72LXLhcrlzbGsdXhPKTJ/4XZ
NKt1LEwJz7fNlN1RT4oaF6kU6ejSRXudTtEr/NGFRWiFeh1koPqZBu9/bAWY5nGz
xqyeU68DJq1ELDgFbJBKkN3bygAvlNCxvqmL/GRU9b1pW4B5VMBGI5N0XrkIqSkT
CRVJHpttJo0ExNs3AMQJPCuZuzKy487YMi9ouI7OuZFpTxNariDjkG5rU3clbV+N
ZZ9aAFwjIdtIi02WWDbCBDJpGMBeg5Gxxz0vjjq8EE0Q7yNTETb0cvahg6n4rWgt
figV0RhZKg8u0wtWpKn7WcRQ1qUIhZ8yPH/wKiyHWaZ0Wofcb2KmEEd10E7UYGAK
+Fr70JHUUvzfvwzWi374N7uh4dRlQGhstjxmXuTDG9S5s0xyrQqyXnJq/Of1HClt
flnnRJtqEW28T8ViuzsiGlXoR+9EuG2oR6xXFeg3G+jw8mXxN61vOyMWS1WuHe0d
FB7fz3jl32Bg2q7z1vzzfiZ+2c5xBEHUJ3pN/yNj0DK5oCeHZ7zB3QQc9xJjlONc
/uyp2JJp58voaVHttKTEDU7vdU5WrdnV8kApltPDBOzvUa06Y/BCV/pMsthxO+ie
w4snRYN5ULki0D2/LFKa1OadEkHPQMM5c2lfEit93B6Nfdf5cUNuLiSj2TiTgYo6
zelzBhvktLZEar9lI7HpVB7zRZgYs4cP86Q4nIwUF+oN66N5G3o5m0BzRIkbEVDs
5qc+Oz+ur6SMKUGNfI8uMeyDjZcgl8ejLZr6I5vSywIoM6pqGmzDJQaP4kXYJO0r
Bzt/uh3mmgSGawbsU2yT0/fmXGShA+CdiUhTmvbj6nQSPYNpVkplyhlj9HyeKdVu
hJklxhk8nVra4QcCl9h2TJZmM3E87sCxaWHVZ74DX0Tt7epcIlp3FNnnboPX09AP
th8JZN8Lprm/v8NVosV/7axXzv9SPDERpAN/q7/k3sFTF1Qhqnm6xH8U2W3B9ajB
c3Q2bZhufWJbJmSKqlgPAfBSFg1Z06xvUdyO4Jha3BeF5DvEyobCa6rm0I8FbtxF
qT5Py+kvxAkvxYHMO5DwU1WbpvkFOKbjl2kaDiYAY0d2bNGqxjujcFECfIvgIlCi
j8Ucq01Z5j+t6hGA0NlzlcSqW2B9JF390TS5m4EFAOuPTFQSFjDDopmQzk6smgNs
xtcf3MAzJ8hrOuQRuo7kXc2o5Gf5q26OrOmw+E1YWEd8XzUKdAHNTyMaywuOB9PK
oaEO93sDYBoureYLDSzV6q5h5xhctzxfZVyngAEM11qiUyekMEc2l2fiCmfIqb70
EYA8RcDdmwkekkH7pg8z0H9J7C4TEyM8dxbjOSWAxs2LeUyWyW9IKHpNxLopHAx6
OMSDQ247rovc+7HvPm0mnxhSE5rhvLIWkfon2sJ4g9ZQLuiL8M4UzycQT6RvEIIl
7YJgihZyvGyQP9118SuATsLyjx87nrAUpz4cC1NGR3QcB00YXaqk/Pat7dLoyY4v
07LO0OR8PDvS8EnmU5oNqM0Tq9J9RiLXpA+ig27Ve2Xc1QoNImFLflsN6+0B/tj/
HRE0nMAA+LBdNp68oHmBc6nZBeCrEHBEGz+gceREJRzSpbwHvni+v5ICfA9QCGhh
raQB6p7O41ojF4pKi6cbn3kFr3fzOanKxpEdYohZqn9rdu8PBcip19avF37YGTdR
whC8+xsX2+poUQFvjcl6e59KkPpz7AtonHQyo/PkYgLAzEwY7/X4fUS+HulBO82X
wC6nOVolpzfSjLLSMIFGjiWfefel7Tlz4dJbMLEaUjQiscOG1djiNAMTi/8xOTpV
Qgy0ZE5mk/dZ3MR/NcMNpFEGOYYf9ULRJOElny7pLk1D4+AS9nPqxorBnZWEea0U
RxxJ2EPmslfW7rmJXCRmCE3i1WHwcAA/mgrgCgrXOge9p+C9EOEBH/jZiiLWl3gf
PN5TN74EMx2u0W860lUKOU0EUp0QIby/vw2srPjK8X/xlc1etCRGJotb/2XALGJW
np6fVjR4cP1yyS2dLrplj0Xp9cA+k9jUs3fN7sh4wb18ttYrc2Tm9kbjvRhX17hC
JCfzRXJ4ZgnCxmH5+tVA4B07Y0mPgjXXpzeXamCwg7i2PKdgUGzD+yRPtGj2r+3o
OhU20cBWcHEBxSU/tyqvZETUw7nMYKrHgSylbhJMxM5OGXmyaRosWdvkskZRkBZx
FQEo5uvR6q/GosakMH/UnYjX8MrBxfCUCmKi2N7OG3PZwPPkVaeiJqutQX1bcELO
IJfD81wFhPWxcyMIMA77vobDespn7TSg6jM5s90WKQsK8U+jFPUQgBnbIRP8vw79
QJOpfvDfcj36/tehJMEr6lofpXfFSEJgdMlap9dQSryl7ONCE/xQmBTXMPOo/JF/
6fXcFbxRIysWRl6F8kHlncAIUQAhleQlyHv7ivGDQ2IhEXFRQVd5W+uCQopHetSv
a6KXYPSE1GSRfUy5yNtN0AobD0rvLHftv56REsnWK4j0YXisOYOS+d1mW+J3hFPn
eJwdfn5oED5KzsKy2LlR9fafNepX7S5d7ASNd8hH2hDZGsrLw3nVglBzFH5MmBS/
JxOVPJvhehvO7r8caU6cQm9DGPvrBGolUmARsEjyHfAIAwiL80uiU24zsx76g8aa
bXMp3IXCBMtNBuF38U5x5O/XXe+IJ0ByEtlQnb2gNb6oEorOkr/+0tzFwO4jLqnL
ZiXmhJ1gaqs0Rgublv4pzZkXFU4Dzo0IqnQdK8hqA1zYlVpZwo/iUL+cuzOesyMu
iuBZEO5wPTjBb19XPoWdTjH2vFxGNFMCQBAZIDX8dFdDpOE7tjbwQ4P7sOhwK6U1
k0IzV2cuCyzB2po1AAXWxUyrg3ks3sxhHsvcsK9T1Yuj6+S4lz0Kht7cyJ/Bv6Kz
Tn/U7prEF7uhm2XNdZCSWGc9LXLdRwFsBuNkPinE+jeTHdTpOxQdGuPlGNrm5lFp
txS95s/iGdhq3HKtUHQ76ERtlFJCeSqnLmMKUq5e1XYtiO6Jqzjge/YJG2MX088C
V66wx3f/TZz5wJJwxbuBU4WO2A+GJqkC48B1s0ZuzajVUH9EN2v0GLuHaYoYS2dI
OdgnzgS445woeqipbe1TkY9jjJ0fvwo2wgyv3olawoY7rtHmSjFJimzZ/lKe7Od7
aPh8NPz+sh8LqrARA3QLeQnH+EfSJy/gGSxWCtXYdNxd8v1dyQnQWwDXJX5EczQJ
vQxhp/lR0SZqHuOS4RtUZURWC0UudZf1Z+LI6B2s+Uk0xywyaedxwKUN4GUMAVTt
2N4/hsO1ojoXmOoyUOSybO+eAiWn5iRRY8HhpQaOxegQVZdlCQ+gWuIPCGNM1m2Q
PUv7MvDC5nRblTOYRlq1v+VsQgYaVtIkcVt6NZwZjILZNN8o9eRpgGtJ8rlbTsul
auqPw+MpWRI0UbyxUzPKxMc2VGdtKT73LJGkzAld7+VKWYUW9zM1AACpeQWSxLvA
UlXovXoJ5HpgagBVbfGZ2IXAXhxogZrImcgl2Tp5JEyxVwLSOHOjo5vy+F3nyEI5
RMzCNwWwUPbCWxU//DmfqhGQ+Lv5kpQbeP9+MGlIhl6hqLBgrcCfMLkmYgxBe+25
OWhRaNskjnTGGm6sAK8yVe9ZZPeYtIAvRJFJljIgt3tH60L9GYlip7XVgFZ1ujOb
dajpIs92qph77VQ0+XsqgGcyfWHYAk3+PCsVXv1+ZqAzgnO5i71Mhs/ra7NmPDl2
rIaoZ/fW86qgSDc6PdqPzCxJEXTv7j3rUuJr6WyTJH+aC6116lWrM0WZbFK5igZA
BRegdJGZbjaq3nL+ZYymRi9yWHqEFr6nJSTcTZAZkYUFYoDFxlAEQIfNEZjV9TJm
5f/42FomE31Vpdy6S1jGe+O2MD3CruCyfQ+zj31EKelSYWAjFQHeaM9YO8txyoyY
LzLrajGJ4bL0waySlwQt3vgHT4QNyJeaH6Gco114nT6stvMLAk5PTBMNcFzp7YGc
GOT1VL9w9SLJ/khGhbTUcsRpHh+slcTypIOwfU6UdlJp3T7wQEsAT2QM5bRV94K4
uy89pZ243w1OGBNY/bRgsNFgxz2aVuKqVMrqkstqx9/lfATy80zzUVAHaIGIgEUT
fMsRDkLVvDaKo222CMzz7HPCqypoDXLg+Og2cLZj87jjCoTC5yFNXANAdIkrp+RF
ealDYersm6j4nno8cxVvUbJdicyd/zQ23Qy6sUOTgnReaK0205OV9BHqoCCWgSW2
PbqkwjZhKUqv9FimElTdptTs2KluJDdmyyu8uV2oDa/BNjLAeqH6lBA/+ez/yIYM
aiuhzrGzo8gPVHbjJLC4lBv8LXmXONmwLw709oFS3GYIM+hUNYDhYnCvkK/eU3ZW
I8VRdVC4BL8b4SXmiiQw376xcjHviovJo/q2IfnnCYtZO5HyF2aoWWXmIvyUwPfa
d05/TYuyuic1pBsaEWzKVlGMsrbepAWoi6CxKM5qajB9fL1x6oKPEGNG36VyGTsm
bTiujjghYQ6FWfUNMAbLP/Xm1H3JG5CnGFUt4y8Z/+UwU0UcMfGMMqEaPIYG6lhb
b3d1J9lBIxwqGUgxOkaqcpnIG3UesDfjbnqn+K/DVj8=
`protect end_protected
