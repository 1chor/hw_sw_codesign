-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
JKlnwBTiTKPdVBpXhyAbY3Tf12Utd2rS8STpNOIH09tpGYsJXavPtFLLH37hQ0cM
GnfpsHCsGdOVMGtIdpvyLEdHYQ84PkF6divV/DsxpJCwGAs2HEtrnR71WkEGSjCw
pNUAaVkXCrv1Lew+yVwtaVIZrGdj3PxnKMWjK7l53RwpYydsnAfUng==
--pragma protect end_key_block
--pragma protect digest_block
hSv9TD2z8t/RoDyDw/9g5b/j2Mc=
--pragma protect end_digest_block
--pragma protect data_block
mp4v0QtIWyOhWGdgs2EDGV+piK3QGZW0dOrKqkyBXb/jDIjyqS+3fFSYTkPWs6cU
XIREpOWPRL5D3pNV8rghd0/Vb8Xih7417JLdRkiCvneoI7PITAYnuzZ8G10q6eWx
WIGzsXtgC85l8wd+Yx5sFvuXaVtS4bIRRa4VNZTNxh5WgPreQlkxIQr7ugyT0Q3u
3CUaTaaDJD8ohE29ivQbk3OzeDhTr/n+khFdk+cmehpxNGtXfVACBIFK/1NnsxAL
eTS90gEbLXQvuWB1pbomfkb0F8NWUdl0qi5UoCBFsopL/7YhB7ymzezKfoWG8MNf
GxPpN2t3q/71xkSqlT4RU7V98k1zRUkJXF5FvOJV9IkrUbM78RFi5Lq1lHHfxmVj
UNWiq/fjoCzBD85+mXHLjVbIXNkZQ+w0jN+tT1ndBE6cWnoRcCUVe+eANH+qAzPN
RVL9eKoO6OASGGPkFuDX2aMPTAr647VcduPd6OBevjfati8h3xFdT7euHGib4n4o
qe7ina22TUcFWxt9XzAp7aBfW9KoqEis4QX8oFEmX/mqjnsUa2/KCx+IHczmWFtQ
vRplbgCqskvHbStjyVRxFFZ4zlvKa7wyr/VhMx+w9ZgF6KEoKgwV8U5Y9EBpx3Z7
DSzv3fc8FiHG6NkwFoQT8A0zEoKeEtRjuuHM8kRt1pP/a5qR7OZGGgn6rMPCwF1E
6FUMCwhDSAv6C55gz8QmwAGpMFpt1vVMyoVx6fQm7rg+pyDc9ZfGb9U9S/2NoYXt
zl+OXzXXPp89WW0XfUTnIBJZ4pnH3VKLJZS/pYiBj9lk9fXBBjfiCSN+pz97gkPB
057VxPsZG2RcHRi+RIGmdCuqbAAlpOZnTf/LSAa4YZPCvsRZxc/NdphNMx9y6rga
Yq6IptzuzPQnM2hBVp56gRNLaM1wjB8l9h6egRmK677n+vmGd6ofXXmDZo3auyiY
N+K0Z/d2AHEKsZypoMswlYUL+uYZhjjInwNw8hbqXGje8ysq3G9DJfcA8iSiYnIY
9VUg+TN5XALyLySz9a5gKL4653IGzOmXbEZPmVvnwVEdHF/bePdkLRZGoRnfkoOp
m9Ywg+hgSJt4F2hPmMZWMsxte6e/ukzKIigTCoiIaMJ2cmv5o/AXI8VMrQM6DsSU
D655uJSJqkYpOV6xbrKqxzE8K3NvShDZ9uEWCDsPcQUJTLP0/ZMhiRU3EzNpcakG
9LjfcofNoEMvi7R2fN6GzeXgX1+8qaXsG4SVjW7UOZSH1JL9RQvvl0ds9X6+8Giz
sxxRV6Wu9bDMmMCQl9TOHPk6TjsM43P+2RYEN1RjXo4r81UwwROdL1/i26IlbnDX
07Jq51JgdosvVrroPRa+zZGEpvo3OtBeSkUg28agqeUoleF+DfXP4bOsYY22+6PK
BQ+hmlqPLO7Phmo5kklklLdZoTC0tKG4Az92dV+GpjYirxrOSgHj4jpUvK0YlDra
QwWg5s3vj5SeP6/iupV8cX8Esuw+Xltksb+2vB6g5Mc00WA08RdHhaKTpvI0sTYd
LUkovlvGklZGyddl2F7OSAmdIMF//3a8wq+rca5EgdceyAOMJuVU1MsFLYVaH/Tr
bUoE44anGoXMRHGzPsImfcPLgH/ZpJ3NRG3Ltf4eFQP1tP9TZN4GAsuizr1zQouV
scRpOdnNcVU3ndMw/acdnykUm6qbau9hK5jYw6U3PXbyznC72OO3QQRLr/QpV7Yo
cmtOochiH0tc5XI5OKq1U3xwx8u/nmY0IPmjGK+Fx0gd0xV5NB8qp1OlVQsiCMfD
Ea1Jk1uWYTA9xfVuHmM4yasGF83a6G08m0KkfauyZWJYounq3UlN+o9vaq5TTVjh
SrUUhh+GuX1Qbk+gWmm0kO02Z9Toy+evMxyfBnHnSp6U5vzpYwVZZWWSyVfnDP1e
lV8lSOaCMNJPjxyc0dwprcOKjUNPRG4rEtvsFg2gOCev3aGlFnXlkxJS6G4GRnvt
mxcbv85BWneHiNYQHoT49biqL0aaLtDkwhzno2SuAgJxxMg7RKiaMu1vfl7TnGfZ
X0WydWNmfSAE4gBIiefolD/cgbJrRpz1i9nPUGAC99AKgyPRRl5RQzhe+Cg97wMs
xv5oAK6UbSjNB9mvhg2p9O+PGZr7of/duh4IxPDT20soHwdXpd8SbBE8IhXT+85d
IolrOgCKzaiYOsLJ4ilnqqijvcikzHC/AsuVuKslOWkC4ikcVUO75UYdc6owIjpu
4dMkN4NDi+Q0hey7I/kEo9Hd8V+AfsCVr/U4QDgojOBektNWv0lR8fzKCqS+vtEU
UsNeuGdTLaAi6vJdSZo/HBhmHAdj7BjcS+xsRmehAUppLzYi2z6I6TKB1FnavtZF
7hz1t2KZS/wox8HNde1+92lZ5Rb1g8xDPAiL39xjPdAw/BpoXRuoeXQBDwkpUFLP
jvxFABPllMeiCaLu8+iZLg99cBrxixkFIv9ht2m4iuOBvCs/iHYQ3XAZzjQ12F6D
s6/a0hrBiLN4AQ+9HCnt0AATO2DXjuSxxfxPCD0Kt4T3CF1B/egdnZH6Kr9jxTH2
9lQReSHkv3UwELFmsl3Ze3GV3N01k/mxPgIruKnS2WA+l7/lD1JFu6n4LMQOJwGV
RZWILytfUeV0rlEPKByj3hxHPV0cFOJC6yRziAIi3pjsV6E0qwEy9KWc6u3Krdoh
brQ+/mbkM1B2Rr2z3DWAhSADQsdnpzpVQcbduUnAxtCcjRpxCSicQAqil7KNKw19
8oq9jpw0hED3CqunFP6u6FvnKr8NO+frdPIg19z7CHMeNpStkbXYl66iJ3aLodiq
Qp/uc/HGwrEz1dnmHgSMOWhmmO8GMy5ZWNBrOtVEBnxL6SvSghBZBM35w12Tec0p
LCOcdi5EZwVHjwn5KSZRrrQmTLDeUY/oJLGMe1jKC6Ig+gIujK3+4No+VN6J43qp
rMWrpO34Lem+KmMhsfR4+DGLdmFTbG8YHjgbdTzmzn6UMBzMbEoiMOGVMRVoDEtI
v6I2lmTBV0o63d7m0mIBtkAoBGbUW7HAVhSsOXmbG1Yvac6F9NiGHYTnzQw7+3HK
d7fHkFtdWiw5QYsU9a6te2GEyLJQhWBmObs+oZwq17aRicu6XjLePSO8nTmBZyCQ
MXUSkdayffpQFhBH0RP9Gro+fx0hA9WbD5SB4JoWTz/3lqkMpZbIf0TwWZ0C2jYT
mTze0ixNAhm8niI9BgbJpUgbTn+PsY86i1Odfgpvyz21FVvLqZnuJeO/ynlu9sv4
saFUorfnwHWFgA352Mylo2JIAqLcp4Cke3auMcwuMWWbYqZ3LBjxQKqGBwLUtkcV
tvROmdvQiVdUmG6kk5NsqMde0PgbKB53QLuF/nwweOoCZm2x6HS8G8CEILxVSfVD
UpeoGRUMjjNm1uPBO++QvL743pLiS6CkmXIz7kbRB385GYITccay8nVNmSOk3ucy
I2iSfamm/cXPL4vHhxTYDme/52w1K8DWQRBmKaweonaNSKtz8V9lU/a9gfJ4t7vp
fR2PUjsSSkuUNa8/DZ4CsZwuetPQ8IF+KQ1me8RKQ/LcNUWZM9RJtD5rCywSLc2d
R35SjyIXLhBHuC5Mrf+UmTd0TgspJQ+sBWBK2tAHDNS5W164bCxzBgYLnvw0xg/n
W+kP8mhMtywtgXFATiMTlVhgFdBtQeLN4FWN4exXoR/mBh1PSHsZj4CH/o8DHbcY
EbFIiXtkxlulGGKtG/F/ebu0B7AKlzih1s7id3FVaq5+uhUa/8DGUL6/JGl5WaiT
G36Ep34tpr+dCoS0B+wToKEV22v5XVJqI5VvFEtP24eu0J/axgTwabRT9A6wuNGU
EUjjLcAoNYF3a1iuYFCau5roISNYZd/oGy7DObddBL6MEapB4GbsYUONtQRaOf98
4qyYADwnXo7Kv70eqhGbmwCHVWhtXiKVmk7cDNY+dsLjyWX2gLpBR08/AjUTSPsV
N/nL8/MI4ssSTze6SKI1lyakog2rNRRVF+C4suObD2y5P4+vXVOLKR/AEjWRlDGn
0ACtxD+eqkRlnCgv8DyyBNEAWqaTwpeSJtWw/k+5iOEUH8MEUNv1WetgdBGSdWB+
s8+Bt6iN212eJSkuGIZXdlOOgLf1pCdTeJzABrdpvDRD4581HpnzLpaDfvKyGWW+
KmTWSKNJq+fOM2d5IQpfah3/1+/f0UefIFEliZDcFAZMzid/3dNoXyxxtM1/TvoS
mrXym1Mz8UoMwGDh9ew931FocO0bqlsXExMZYvq4h15neeGLdGS8/yNfHEJWaZmq
N8Qbndj50pd4LoA/94xeQFwt06Nrq+gPIS7I52eLXL7TujAvTKbMmvtufEAdnWsy
Y7zswS3NbixGAN4ZLYFqUgxR8oj+EJto/PUersgEqtwYGH5Co6ZFrZJ5aGhXs22T
XVotkTWW2OY5IvbeMY6ZWKCU2ls/sZOKUfSK+1VfLCFONWaRSI++D4K7lbgaBBj/
1NIcjAzr15wfWcVTSIFZ9K98HG97519znLbhZODCJcHatILNPERTaKiHCYWFpem2
h0G02OLF7uhhnlFsDadlEVXRiX0PuyTjClsTOZoDFX7T4mFtd+3cZHdgjx9Ulcxe
Imy+O3iFok4MyQ1wVqxBBahxxaF0CB+JTRM+Z1QX+14gQSAo7hJur/5Aa/Ugcj5L
PP5rfrZ0gnD/IA1YFofaVZjnJ5RnOnyV63kdkD0fd9UMyiNwbThICXXcxRSvU4B+
KpaY6wp4s+GeGuaOk8IqR8as8PtZf6+qKJAt8xjr5iPffFBIcLEGpORE+Hb9+dm3
TZ+cSorMP0mt2o2B7f4JHcQPEB3IbzAUvti8QLrodXtyAU1FCfswTEqCLT62bbty
ZiEiqPtxPY6cnGvSxwiFtgGClOvHfghQb6uVwOzdTh6DgI7EeO8Rlrzq5vadWlXn
N2cb/7D7/cs7AnnCHp7Xzj/BfsWjBp/gy5y2ETVttrxJMT5+VJGwxkv4o1Kf0C26
/GjDf/1Rq/nQUcxbDyzev9uAzfxxDeLkXOiAE76EpWDUO3oatlqNWl4kV4pyxoNO
W33AOLPi2pNBBx1+hE9JM8IGqryZG08lyOgOpN5qvSz2rNpfoVag+zzf6ym2m9PM
DWXTgC/3WmTF7T2UzL6IunL8ujIis3ZXh9Epc08Idu5k4NqGjBVr4y6JPoiTZlu0
8Cg/ftDi64eVMRu3vzFBkR35y65Ly5gxXoPRHZFn6T6d862UMUg14Fookt5RXYbb
D2MvFUA+Bl2pzSLbCIGmzfS/mXraGBUgXLGMntxmstHIgY3jOZXX3yGH1KiJ2fKO
mPRy8zgoFl/BQfhTIYoHm3cd9fK7i4Zi6zQ8g6cKLtflTTCVvWimDaPUbRexFYsR
dEbSVDTymsx8b474WBmDzTk6ZxTTYZYOxLDny6Vl/aWyWiko2EIvyRLlatkIKKjh
nu7pyDwngRSuM2bdxikwIpORpiyEYj5Bch1vcAia6w2jazcUs/fBDLTKPsc9ZmH0
Gl66G6Vni+mu3gD/OwFsoqagN0na0Uvgx7mU7GY3IU9IeOaqU3iGpizMZWe46sdv
NzZwsgtphzC3gBa7TNAxCiptF0RgTgWhABMsGbEcsRNV4rW28uQypB+ecs3V4aXg
M2/F+vpw/1yFMV8RTdYGKmrGMj2VQWQHeQtGRuY+cEXYMW/nvReDKfT5pVgDWzRn
H0NHLKxbsxAz5WbbmTGcAh7l6Cml/kE1MZt/pKu+UTqw69mz5sZjNQqPWkdCH4sm
h2d1tu6dsH74Xek9QOESIVoQmwmGdJzFHsdlyEibv7OKX8V0MyI6p1IrNaUB3Hw9
Uv6e3gcZiq0X06NPQT/X3jUWTA0POIx/bSBvwCFPX/xHLbGneArELLoZOYURVxTZ
hMFad/wKId+ggvZKlo9Jez8SH5qKoyTH7CEEkkMCWKFr1nbYsxWgZdalCToPgP9D
9EvJFKWea4UZ1ThCRtxLJ7ehKUei5Z78raAVmJJYxGN4IMixUSbSXkt6QpEErEnl
3oKw7cz7LKSqHL8DD+v6WamSsAGLCFRWUMueTgvNfAvd74yybfTP+T7exs7sGXh2
w/aDlT9lZDCixWTv+tX5QAVQxsZYYnezIEsw0/q++9gU8Ht2jYqZV+3gd9OGV/Ty
bVjTjAYY5bhrgUPvn0khmhWhg8uqr65si7nArFphoSFOF0JuSo2b63od9iZ0m7rO
dkLrhvf674wup9bDezJVmAunUecOjvbCn+d+dvtUVViCj9CzbMjQeHQ8u/SGiGNZ
cLcIv5feikEmVIWKWhzVvRazbS4I4Zpf2WnHyMomX3dFm1iH209QUazcHU1DQBU4
t/XqqG4fECiU1RwdttGskH3FQTq/jdpaONCfx/ZeYphkCD8i0TUtltK84l2rCokq
eAodEGopvHZT2b+nRbk4ahSegMs3xD2/LyDzi6x31vA02C8m3uFwwECAAx6jbeVV
leYSYcLZUIPJI9iJ38gmRQIrTQQz8xflVg7Whz8/SPQACsk9EbIzJXzj16Vq5ON8
3ITCUHiQNSEng4M1625VCY2t/uvXTABssNtSfGTkYfcZJGPs8H295O8ZbDm6V1jo
cZeTwz18AKIk/NTky0XJvm+s9HZSv8PczRVIzLA886uCtq5i1u5Xv9MPJ/Ktvt+n
AIwGsxNKjaJ7b1o7nwa8PStZYKn5f2LTRDG0QqTqd5IRCCcctZNXPkjqEMIzuFre
23FkcuCoO7X2UvMgiJ4GHeSH59DJ5XwltbACTt8yiPLKJj6XLU0lA+fDmbB0l1UK
Hz9DI2BWKHeSk6SXtTGpC5j1ytDPAH+2OfMwZrSNcsDKFrEOwrt/q60MVEotyaxt
5hI4fV+bmNsw+iqt36qN+6Msee+ltfWLjGnXhrocizNaWAe61a929nAb7E86ndEt
s6JS692+SfhGIPF6b0EpQk1XG1hSTpXOn6I3pLXlO29kAAV6z6kGqYPXuKdcMyis
phN3BCF1OSHnG+6iw/rDrdtNeMe12SYiUOUSu/y2p87QC6aYlf2B8orHTUQqyzXP
dPjItXX7fTzrvXgCPf06I2NSRfqV6TGPGFCBCO7lu1uobHhrc2CRahofXHMCO84y
tRuCzDswOdKhWGa9nYqdIQQQUOJgvZ5JZN1sjRQjHe4lJVciuzTBHD3zLNTY9Moe
9Tic84JjGTZg84ICS1fqFrkIVNsbIGOFOqXk+pMxiGpLxlO4bEFkzlRKRFnnmef7
aT7virX+7K4DbhcwnzumBI+P7V91TB2kUOKcRwEDCMZAg/xgZDld16HzElqBRsbS
asEUtuv9g3rwT5kjTyr0vLgYo1GvKJSM7FhzYAZS3Xgv7iZPn0Vcf/oJL1mnYAll
pUBld3IkUZmK7YDJwUphTzpEB8CSjIyxLSJvOzfMjF3QyNie81Km4LHk1Be6Dj6W
En54ASaCX1Hcoy3A2C6zY2zL6WVensmpPjOBXySwVYX74VfpxPwCYEQ9vOV7YipB
joVi6s/U8sJM+6KyBFegLolFneqU1iZi6XQB1ez7uHaRWfUnFlGUv26VJZq+m8MC
fCdpf7mXOx96DzcFvhjuAxWam6UX0LVzYYIaVBk9/l0fOJ/iSkhGLWrukvKlDBuZ
Cr2TGlUwEKSEtaisFLeV0bHQXWKbXFEj+gBjtF3IC0/I7rhTyf7eNp/61FLhnaWo
/N6NSNaT/4ng3l4x3C3qxKiws0Nn4FiKTtyeR1USvHen+lcZSZGS6/3vIVloIwtc
vPHyZR1KB4fODxr4uX8cHCELbVqLD0W+fqKOhHH2GTIcMgKy7heUEnPx/LsREKTo
ZTrCIscYNzyjhHhE0x2qXmc+IUnxqxHq2vse0gD2sPeDAlmJvEiHJ9B0NAr5rrAX
O9Z3Dv830U7QJwMpMvIAaL2htAOSREEJ+ttzFvGZ7zNLRqCESNUkjKTQD7CiULUN
v7G/j4LKkeHvz8JAMav9uQBQQLXm0ZxYk2UtucnkeBr87xYb1hoClnzyPYafuHKw
OOGqmfhuvp/p53LUSXFa5lfOLgKPGbUfmR/maFW1knj+Wxo7j3wHvcOqkOahCj/k
a8mt5D1HcKWd4XUPaSlMA/ifIKnKKCNA0z1MwFZe2vgjv+GGz6ejNQtfCN7yc2fv
7cbKQCPoNuot/1HuhEjmgGlQ+S9DYSOL5KoNMP6YwIx07OoWATa5tG6MXbHaIOp0
kR0p+LFeaSPG97LTqSsSwkxqAK0iDLD0vCl5DeG/Uo+ekxmjofEDNo5QQ3EkX60V
P9B8zlrydAwjbMaLj+bSRDGWUBFJqXlz1eSYMGGJKIE0rFr8nlyqTEriVCQAIyOm
zAImme5bMlcysfo0kU1rbDldXbmm+02xawg8Uu7jP7kBWycZfif3D1DjRTYIbmCD
7+V4tHcOUtfL+Ckk67JeOvwSeKlXTRT7Zdo3K03IiYJmD7uv+bfW8HLJnLEi24h4
jpzAWxoyDRch5atfJNzfBviao8aILBj+ZGG6ZObkRF1Xyxdwq7EG+6ipGaxByJly
vgtG2aTiclVCvySmMNo5f3fqWyyPoha5MIUV0Oe91xXGxYYtqYBwML9I2KIfttvC
vMxjsphZPPB+xISBldstk6ut8ArcCMIJbdmQbgj/JnKQEkVyPEFhF+AeR5hUhe8/
A4s/T7HIWIZSMjecmfYPh+jqOMsxdqQ8IkOXzNTW+21x7KLZVrp9RN6nxcaHMAbW
eq8A1My6qyGOF9/jH4XT4Oc28D9Mbw5W5qcVb/WOjpORWyRIlzgCNb9XQuOkkx3y
zAiqocEH89zrJMtT1dOU7Rcalje7sMYNmuXBZSiisi7jdy3WGC/oTH55eai1S/NF
A1aP2f1VCfVzzrBDUrXm7tDLxGqroDlEKNwrprRteaXdgwyFzqjoKKyzM20Gk8fw
2ht3hZGETKK8xwsvAE+t2AXJlgoyCvtwapQlNEpn2FVTgy8JWM8dL+goJHQib4Ro
D4v84aQ5GH9goGzhLm2kTIHEOLGaIA0XqzkqQtGe4/r7/3XHN7A8G/Wh/g7f1jcc
xlflxxenBMvjVDMhDM5caMGf2YKhC7M0T3ZlSJk05B8dcWTHMv0G+FMySwYmYq8i
0DbMIHJuGtS+4o2dt5j8X5AZ+SuuWZpluKaUNDUqZpJrEoFKAUP15hAiPQuSpdbR
MjZdc5ilxPjCSTTMg/w+rw1G3V9ogjwz18rDv4Kd+SI+rgGhA1mDt7k5LAx/DJS8
KYz5TMc1Ch9tke/C2QIpHQXx1zovYsiSbCPa9SQuHcF44d56UPvep+l9ZvhDTYUW
YWC2gf0DGvMrgWH5fS56sQb1m/e/VMuRRmnUyaZmrI1xgzuS2ODB0DKuzeHdqoIH
udFubaI7+Vxs1mCY6feYIufBFWN3NXY9tDQaYp4tMgbO7LFJ5TByTEkaoI/XDz7x
WXzzrEy+sGJgIBhq0U7uCEB32HpClF7niZ9UvfGO3mVoOTX0zgAwUVg19VVHgE9G
g56mxO1NK5Ire7R6E7riG5gBBp31rkBqR5RomOFhaxvz6K+bjLXgp8vx+mhni7Y/
MNayClK9zaYPGV65Ed5x9JgGB2LeO4fPv0VUZ97EgYn3CHAQV3iRb1yzP5G6Cm/y
QNFaTH+9Fy4Fc2NKtoKHmfFb0BZWnZXBGJtikTQkP4J44H3UFP1e5IFwntESR+2T
3f6FepaAwOyzLhzOQOG60NfwEE4nDeJvIyEmEM/L6SvC0q3zbLlg6d/ssA0YbpXo
kS1XZJ9U4NbctfMO9j+PEYHZyKAe29O1s8PXbs7Ltxp1Ka1/2oKeILW8uuKqnJRn
ZlqjyfGIGF3vtzVqSMMBspgayxxx0M3krCnVHLzQhMq7BMKvBHMAnvyTzphmLecy
L1r1p70IF/vR/1/ia6/lbGsHQ5n3QgWxjKdZOaozD6EkpGnJT7fGEIuCh+yT/JMq
D4TAIKxNRXEbevqsX/4lmEhFo1Y8FJZX/ZU90xmJ5naOzyiK7nq1fOj+bWu//zmM
qKIBWpawqWBGInm1FNfa2uD9Lyg9FVRdng71bPmqW0Sk8dDJb4hGBG4EjC433NjR
71b7H7pYG9wXD9bzcuRW4EF2hFFXhtu/jKdOWUhVtINAWhfE88SsLH2bORVFEbjc
1a1mMpmzd0Q58r7azQsn/gcTM2YwXQ3vbx2ceP89a++TniVshVEAqfvQCMI3kP7U
T/rKYbCjOvQyOsOlC6PzVtbPGdcIErExvWpFBwu0dwrJ0+1GzThx+WI8ha8uZVPk
0nwmqrmQA+LHd9skSXL5ktuwKJ/3KnvojgRfwtYbEo4DfeaYPfDxYYAse/mlWgms
pY9joirDqzbDsME6ZWkybx1nfWEvyo6xrynvcoiqeihgsV1VsEycPcvMltWbe8qK
DCtitubVs9/BndZMROKvISQ/TZA3zIXImSsyprsAZSfBxY9PnlvOrH9z9HIviAgz
MskgCW3lJMy43XNJaCqpow0Lw97nB4XwZLIRdm1hFGEmxLcLCmZD1Knvtdq+/Df5
jdZi7g6UEkkPsREaE65hNnRRhDPxcJRYcQnV6a+D7ZvLbwgbrYltR3XdIuIYF70b
rMvPrbe01WhW07g9G2Os2ahkfOJ3fmriC455IrxKLg9WCX4zmudouI4DNuX9/GOV
78ihAnJm/5z0mf8lAqxue837NLeyqAaQU1cgBud/hB1ibxSoOWqvr9NzLeh7yts5
Pvc+WVWKl3PmVc+XV3wsBVBvjFJSNPzvioIf5qSJZ0I+LUIuXCpmVdjsICw840Lp
zuX/878Zr2AkeiFCBT68WoHXRzOp2iJ6PlcErh6As6drNs2zKIRMfRiB4lKnr2VE
AfLSb/E4w77E+CQKhPCGNqW/LuMDZXP46TBIdowA3jTWo4IDOwmieGmHuErTk10D
R0UzVNJPJxLQxzjxCN0wskBgN3kCFrdfXg21izSW1oGZ0fd9Ze/5fTgPb6dHjXiy
NO51RGqsO77lHJwtRUx/fnER0XLJI99JcA4pEvfeZX689Nq5FQmCjQmmLJUMDFse
ouJ91mbVVeufeO+ObzM+DTe9ndX2WW65307DU8B0Q1ahqtUp1ON+v8CR+vccYEWi
SXAfBENxCkaLBF4gGnCPHmAvZ2gt4iVMedsnYtRm2HLGUICpV5pfJ1TtHt73hMbn
Eh5zkfTr3MF7m/x/L4qAclzSONfco7BUghsNAPb7tBXUlbcaf7dZ6y0c6Dx/+wFS
1xR8WYKRlTIJNvsKPclxXu8hx2pE/pbkgUnqmDNBEwZMBWKVq37AGdK28+LAst8Q
4PE2EOcNEfRJ/euDPY2BZcHAdyP8kSzeGaSonRTxFiZwzQE1MIk53wdj0/rczmMX
f3KswR66w8uNs8nXdPS+u28AFstTVDPlukRlzUWtjdUy3eV00zSkpulk6b2StIpE
MG7bS/O7MHeHKckv7xmW/1LZK/bnkr/tTgpP+Kws9vZcdNgBoWqSgxwnDPDmkXSO
12VUBTkub3VdYuzm5TQCJjM3HqcfryegbdfkM0/E1RQDt9jjd5U/xxcQ/uli9JpY
WPoEurBpRnNTy5zcHsaaUbb38QJpCZbpJ5ddOSmCghGb30pRpJ7nX/jei1P9zQQ2
+4VA7X42yRJFkew3gMxl0vC/P5paTvcHA1GFBPRLci3ED4haN4frUUJbfIuruD+L
xQYg+CfPCC3ZlglWiftWT6OwCi7l72dR86Z57PEvpJM8CYo0qVXt2/D6MOivU5o+
HTREmEAosum7cq4C0eTe/XBvx4fwAlKWB78aJnpfmPvbfFHhz+fPaoYRp4PXbwFB
7Oy3Fn51zYXMd34l1Ot6yzQTB0HzJ/4Ap+x5YEvKS2RgXq8ZnaYoNO2IyH5v9Zer
zKmY/aROBEHnmxxBdPonhlLF1PSAfGWGJs8T1J+/nlg6rczvmElULEyazqxRlDaG
AgjZvdZOTRpnSNXorsWoaxc1UwKQHOY9WQJjTN56C3MW8RPa0REHTykyu5tcKsRJ
YiGWCiTM3n7A8IQuI8PwhVHyinRKUzgSronzBKGeDWuaKjyGPaR/0ILClpYIo4LK
ApSfdjA0TJgl8Ol9yq8O32QyncEW7GZAfTv4THrDZyHjb9IOIe9917Rpy0Y7vA5v
/ZTUh2gfdVPAR8bBReUINb/PrBEaS01tKHUqqHSTYAS1Qvo8sSBsmrAEpt9q+La1
8LiIwbJhlz78xQbST7tNCUCKr9jorJkei9A0Q6Yk1Zi6UoceUm4BG/TZJycwui80
eR8CpN+UMmBw9va2aY44wpxeHaAmNI4LywINsB/RzPrKAJMBx7zwQ3IpNgGrPz4d
S3Fqo3dKjCT6F2fuDQkc8g+vpk2qJmE1v6TtcutA04LIGLT1JzRuGYqn0sL1ThkA
vfDg3oXaziPVDHLBrnifF68o92kBfvdyvA9ownreuew37JbDQkDmRNZGN8+1TguR
3Pjnie5fOLVaSIsnw6MB0hGtLascu6dzz2H7eFfv5LDMIIULxQ+eR4S+XkGpLRAX
c8IUkGq16/CMgdqyIGcJC9cFABWKGpUf2mMAKObEbiy1TWLOBxuAX/lmQ98TACmF
OEtTbHNmm6Qj+gXNltVlw+wOgMKBpiMYOxYrx/f71/CsDFhBr76jvkUpbftldV19
hemo//P8CXdM7+uR0cPMWKeyx1JWomy/Xv/Bwaxi09KjbCcWmz9b0WwwNowEyYrS
2wQDCYjvSSq9Ih43azfQPd1aU07yVNxv0wzK5rW8azF2Z2G8SxBaxS1z+GWabgPY
kgs/NywtX/qUUtwSrhU2dkJKMHCCyznvaSJxRiXJf3rtJlQh82uYhm6DVTkKHnxJ
HzCLZUejDN4qyam/aYtJOyU9Pr8zZZu3CkPscie/3EZRuUsxwJttuVRSn7jv/ABj
tC8tOjoMIOlcRFUY+zNwrjUI7QdoFvunvQje5xCpQXkEZROvcylv3fx2Xmx/edIt
RVtbzpE93O/2zRnCA3A1Y3zxMd9NehzesRefzCf0KqMtVgcwbLjlGstGk1Qzuxa0
HQ0yQOeXqXa8x0Ta+PUd0d3HAoKYeKsiZOuHEVuUQ59tBX6EirxWq2MYBvp8gJxK
PvxfmQLlG2j6j+p4p6b5L4gPuaC3Xj9t1jT4dtQCKYee86I5jvfPrri55inti31f
0riFivN8JTlTXcVO+4E2jN6u0WNg4ZvjToUZcha6ypZ77BkGY/YkmfsJPeLgNEsn
r91omDgyHgsXRaCltG8XGvpnv8qolE6REZAsAYeevxeO6NWlxK9iOJWqAqkqMYyY
L6kNM3SCq8ztfFPqA8jWqaz9W6QTPymATISKuX/GBOTeM/DHO6FhuwopFzGmBRQp
X7dVlIMvO0b/UAQV05PS9rDxhF09JEWIC9SneSNU1vbS7jePVo0Tc5SgU5eMtB34
R6o/E1zsY61MZPKDHQJLlrHUCfDgvcFHo8lK3U5lJWsJHlcAOZBGsp5EnGkuL9ME
uSe7xO/4t96AarZ7tCGlYli14C89e5mNuP5oy7Nc06YdGC46WBjWOn1jbzdjK41J
0h64Rgtk5NNsmF4DjKiTY04rTH/WHPXN+gZpVlktWxup5ifaLf02//+50fOC9Sog
S++hwM15HCbkXzw0WjLG9swcxNlGXro7HI8ynMn/TgrylpjSEil96vMPMdw9be5/
YMW1KZyD5MjB1jOFgfYJj+Een8Ld9Dvp5EmuIvFwSAwM0/sAKe0krqTkGvnT+fm4
hld4xQq5s6kihRCgllAhmzEGrqPLXp4oc7I2IZ17SkipETiqpzyf5IAQyDpZvrh9
x9MMcrD7aQQzxUbckpoPLTDVBLyCyxyndL0hWmpPYqJzM1HUNVTOPUHu1bEzd4zz
pl9Obgz3cigvYOkJNOHK/ERORC2TxFy2B4mQk9NMLS0cL4EMPVPIL9nUmxM0N4d+
PziJ8bsmF9PetsIr6hqQYmCBY20KwLiOPN/iGqu7pSyACWg8DdPtzTsoHwWVO/UQ
oKZ3KAC6ESNN+bdVZw32pHlhiofKEL++18kOGzbpc/611g/P6fSj4R2bkOMPFhOJ
D0zMgqftxMUbrd997GH2LdCo34erMlKKdeBmD40n1Azkl0zJc+LaKakF1yrRMIVv
oufl6Kh9VS4W6uAIrwdsHOsw2Pkz39voAqr+fNwwQJwVvjThWw8XUBfEWgKpVvdG
xnSYsCNx8tdSN4Aiuh4DM/vlq8KiL8oy50mUF2KCci5ZIwjgMBNl5MvWDw7dPPIY
wWHQclZAYPVqQ24i+yrWlPa8ldX0Thg1KYZfW2X4E7yY1qPxK4SF3/ZyPe6RnBhZ
a2H0q3zvORRCXBfDDmceMg6fuwYx0CT0eBV1WKQN3DqrADQL0/ArIio68z/anUe+
2TeO7todF8SjY+ycMxwMsPUmS7dTyXvuTGiZWNaEFoNr7T1lQiQPFp+nPYpvEYgh
Riiax9tdMPcnWnQt/hCemhjO11HyONTylB37ATWI0jy6rYoy2XIX7CCxTqPm0Qdf
w4HF7K66cDK1LSQ7fYkUwozpB0D741SYt8Yls6SQxmfZKBPb8vRWeuujJYHskAQa
/kzND9h7l5f4TQFszvFscZlWMMHqBrfBqD9vCA+dzRBFJVorEHy9wcXzli2pk9lP
hEIXDUL24Zg2tB9yVc+FkG1jmKWl5SA3Hl4VqVmJkFTqPynZRde0rWfIIYYzAbLm
m5hjCOgc1yv9lJRXt1jmKh2QxlM7Zyz+RwGekJSSMK34++eZ4VHsyz5c4ru87Kho
W+3M4nzwK6Kt9TnRB2HQBBbzfr4Eh7tcxyXhE7uumjywN1+/GIO8gBizzaLr7WBr
teR+C3Zga4zfHIiJZEMbp7GT/QuyykVVApYZISY9Av4R02JY+qcVe/LJACHtQ0RA
8gnlqR7SG+Zi9BZgt6/MRUJqRROVd+yoLpZxAx6+Nws6AMt42tFjysCGrkd/QeQz
Uo2WiprW9X+60FofQfFofd1Sr2I7FDK1yJDMTqzCCzTCNPgPKIEg3wtJQ+Sqb6sP
X+9J1Lj/maxb/Y+nVnpCAkDuJMRTAqwTzc+GDWgEbm1vNrREeR1a1VrnZ9F4enCh
wShnKDJ7Thw+hBC86eOUvj6czSc3UFPdj0q9eKbVVfhMKFwROVntuFrLUhaIf6Su
s/if4mOQkRGBkK5EMI45NIX+AM32jafnbYiLqf55rzkY/JIW8JhzcFKWVXIwBCTv
YqSumRdICHe2h1GvBWrbYcJ5VGE0Goxur4k9JFVTxUBBBhvp3PLTOnJAvBn+r/gi
t4/f0ZvGKJVZIX9TkladeN7dmTP2hh0wsvm907vIaPLTvIlK4h+FWRrfve8CRkjD
okGZn2kFM0hxvN0yHjf30wuDFgAYLGbnacmPw0cEpvhdD73vyEa311pqADOQEjfo
BXC2argQOm8tq9wEhCOejO2jrYYC2aBYpjWGJMLYwe4GoLceVeJipgVezqvhqaEN
+TMZBba398OJmza5SVrQV5i8vIIGLmgW7/rybv/vTbKifVGCBd9kh1HqlvLFONpM
S3h7h7NaSd45Vbfja2C1E4dguZKl6UKMDXrhYGIvxGFWgfqCupLkYcTQTzDvRfr+
P/8x3P5Sw1qSGM64kwA09VcfvHl40xPObd9UkriBMqLRiBH2XUPd/cUkAhWP1vG8
1S0dcmbBnqi9t0T3SU41kbmAI9+1WIfQlffeOZKgg7Ao9fzY3Ke0lx3bfV9c99Qd
5cDdtu8/wcovqxRa48wz6qVQx/6uBzKSOaI+PEFIU3kWjIW0eb7f2+v1/RIcmIg1
12RvHalVPqLaOf7LFUPZ6Siuo1s6p3nMxIfyOXF95Wj5hZn8mY7gUrQDAdNt4kTZ
9WJZ3NWM6I6DqbV9Ez9hLtsUDSxKw2sc+b2IxjVlFsL2fgCd2FHjD6bRoPZWEwTl
5iVnad6b8ARuGMUhw0HQekRpcY3YWTgMdbUDJrDMCqOeKwWUnGvDatrjHZcu8I8U
btG9pFYZ2FaVnnXYF7VmzQbdu1mOnbI9/nQiWZhMhOCqQKqoLOLUZ4H3rQG/beAS
BbwzDG3orgRDnilZG3OjVFFw+g1AzQXOyfBELfHpcHM2krjDsmzk297TzGGxm1Dl
3b86Lway8Hx49q3xITFBEjnQq65pjE83eMWPGdfCLQgx/Btsskemtg7Y2rMeRQRr
8zhzruHm7KK5f55JbS5pF9cxR/Rva5oE2L/hT0ScK4U+TMcDyY5fCd3U4VLIjlRh
8vhA+nGj0Cr09okB6CICIZprkcGOewlvEN0vIDG7KNpRZSHwsooCD2rS0pC3tI1z
lsyZc2OnEz5Heul1xuVg8owjE96bHqUgUEEqCma9HrGhDlHUFIdh0qrw1DwsumS0
m4XKjsc72R6KNJLJd+/Xdemev0XzbTmr9hR0LSRiy18/Nm1G4+QwvFQI+NK1dfC4
IIr7HnRQiF2y5NrF0EtP8veRzxt+XjDffKNrMRd7/WEg30n3AR9pd2cjKPo1zEuN
HkhOJYL61oUSmWBPt5QHRy3lOlHDvMMS0MnlRp5SepWYd18b40Xi/K98a2x+mYBj
5j0531rezmF/lleOv6MmET/3dhZKUQ/kCTLwJevriTMTUnR4BeNVSV0t2edWNBuP
UcuzRFxEgBUvave/3BxGS/ZzJSphLjNwewxBBpch6p8ChcCnFrEH4ByJ4X1N2vWx
kJ8cLoZLROS0uj3mG58xd9XcEyf4c8JIDX8Ii4ttfWqDLba5KEymrQLfQSB0ulKK
U5BTNj1E6a25ORZm32j9b3zf6XN7YMHhqvC/ZHr04CT6VCIUenOEZPKuCrDa5d10
MQ97et0jaGJ3FjEdaRXA0p3RFBbcMvUGwbVfsoigkF1bz2aMpNBBUVdHyIt0YWDO
VraYXVnHYBJw/uf7mEEApUUZYMndcnzZQ2g4B+94vGHdTdCPrc8J23KFGdlxK84O
1MROX0H0N7cupoCIw+jfTtG+BkGOIJsi0pklfi1K6ZP13LA6et9r3GaguI/9Kmb9
qKnoO8EKorWAJOSwtQXgFNV1997ok3dPZdB3Dz9laiCcANZfivBk3geXfEWXwUQY

--pragma protect end_data_block
--pragma protect digest_block
mirQDrZhHCIemPzESdVBWr1N07s=
--pragma protect end_digest_block
--pragma protect end_protected
