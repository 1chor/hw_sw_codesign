-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2NHhTXUYaVo3pk9nTpo3KG+iXJKWklci19XNoxm7O0KLu0E3W8hJa+w46yWrS4az
5epHbXZYH3bcU6YQDZX7Rv8hWOKPqRe94kmc/OCw92C727cNKISBKh8f0t6W9ScG
RxY2cAwcCXOU9K8Vmheg2wHXBkDsUsV8JKQlzhS91jg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 190112)
`protect data_block
YqMjZmn7aAMTyej33zo7taPImX+nJaKiNcp9+GEN3WpckkZEL58uUT4dsWb7LrQk
qEDLwqqm956JLxk8CJqVHFJb0NDGYo04SU5n0VXM5412xqqxSsESlekJYKNFB6IK
io0DXIbd1iAqThVAgdzwNfBMIccWGkJvnSm60mbA0pa36uSS91EjDRugGO5kjl7+
arHA/lLW3lJgOppELW7fqQuzxlT21uKP8a6BeAPwr1AsVfXU8KTgwR80Ywk3CIuq
zRN6ktxykKHA3ZDUstYs0h/4W8CCBxfhmQo/fL+WeH+02Tux6riLyaRUz0lHdCm1
jwP98hLbJmYEGnhrNQIcvwt9asEZRJ5nZd6Wfo1vJ5mdrkVXzH78165vtjLnc6+9
oWJ4HXTWTYsHRTQsxQ0rUGJXv1EyDan/Wpu4eSbcN5S+k2bCQChWWhL6GM6C+9rl
DH1P7b6GHbV6hBmCy711FjTWu3Iq5JbvpG6HOdwxcpKSUvwhYdKWBY0290tkwxLg
7lFbom3JbRq5rMoWiuf01ArcXaQqDscf3xDLdsSDObFu0eMue5N1d1HykKl3mcw+
z1Iayi1lV/rkFNzegK8oLjY5LwvLWq3J5ga+s8KAkZseVUZwH8PbiyklJYfoQ/SH
lhQcE11ws921cyu3gbfgi93JK1PxdQycVlLfwIxSsMlZgYoi+QEc3gusdWZxnwqZ
l1VZq4BfKS/eRkuFd0gYcYPO/bs5v/bzFF10OKMfz8/EalR9MUvlorinwbMOJ8UG
cPOzvUouFw4WQLMRKzyEqKURyyas+JngZZ3sNVPW5Zc8JaQyHtoFCK+N5kvoJdAi
nLYtCzEisxGB3Il/kzSee7ST0PX6UbD52WtNKM+UrxUuFKwLNTLvEKDs2QGbMDsX
evRgRGYNJRrPgi0G7wfTZpx8mxoUpYeFt7UR6BHpRXRsFKQsvPrIId385FhaCxpK
OjpW7pasrkQIuZ5KuxqVZEKOLaIk5isxf1EmtlONj2xIwzyuw68O5KAwbUX1+i0M
D8TUilEoUIhmsmYso9kipXA2wcXvsAK7s5IJ1iwDDI3fG1WmR9CeESxu0iBUCkD1
mjF7ib1jOLJVRx5bHxXRgD/7uSXwdvGo4qi0LJZEu9iH+I294wdltMzlYnN5nTFc
Jrwmf2WWuZEN3TMpb4A9wg+TozHoLTjwi7IqXQpolc83LyE9lK1AVoN7xNvd+t2X
4DmRccQrjWkfgAz+pvfISEB3/zFzzuvfwa6I5X0TnQ79uulDNbkRMFdT9OuP41lr
u7m2ptoYygJ1O5a7VCAYd4LjJwgJWxM9Z9Ml39bKr/62WigzK8zR2eTm/neSeVGZ
PBlztjtAEd0orh30HWqgYDOpt7dtJBHKsAooDAWhHM2/uI6+FFcrUsYpu0Qkvq9s
sDKHsiVt4ZLRB3vqm2laFFYn0iNosmpb5fGPU6HSCDa1jlsS5wRy4Uo1vGmoOEog
tkOW53szH05NL2Ekyanikjsx65+yBZKfK/v7wO+weg+e32xiHYpXBNvPRvTmZtSM
DFlNjM95/Muffufc/181SULitpAOuDP7cpQ5Fz7tmE3a+5Gcm8AtzSRs5jdSs0y+
1DGzNHI4JnAGr+K4ID+X2aJzNmsnfVq94oxQbM8m6wwd7CvoVrcXtMCX56kVBXNn
NvFKqxazEvqWaGJRucw6obf/K/8EkGR+zw2kU7uzN9lCwwcySpXHRTCULf7+IjH0
+rcwtpQxJzdI2JKBR9zqESOifgA5v8YJvY71/yS2M86i7IRw9X1LcgZe+ZO22Vgw
kqTOrKopmyJ/OHS0DILG5mDGt3uNlT8794lj1SxfKVh8iNXv6+ZCCI69LYggkszD
wVWDyon2v1GEtmX8UK2XZzIkF8dmw7HZsv24JlqOMh6VuEtg1iL/T9lvZ6y+/tt1
QRgS3hVVvg6NM2OWBF3mJFxTVavm9/66Fv97ESnAX/n9dawYq7J88N/1MNajnRMx
YYceLaKwf6vNuV/GlH09G1LSH4Ji+EUU6nWru+F8jX5oCmidVOT52DJbRURTb6G7
57cvlCCg3+Md4gLz7zMHawHs5TdeWAlQ5f6gbWBVjMX3bU8ItbUaAY/rAYuG66xU
OWGy7/Yr4+/a0QivHDjgs1RYE1aC+7vYMrvo2NAZey37rd9lANstChY04YgqCVXi
IDQpjhpAe1J8Lbp7yiDQbuQTowHj01uwg1NbIonA5Djc6YNOhI6CPImtm9ObF9a+
oEnHoeG/h0XOopPRh/bIfpg+C/IHjtTukvxSrpOkBVcfDkS/9LGarcAQ2TWgbaqE
XHGLX8CoCyXY3FuHbdOdGsgZo51DGf77///KVp4s646cUHzNRlkHUoUBIPxwPnCZ
tFaOlh+l+KH82wyWGhjNFJPSEikhPNsuKPNQQr0YHSPZEbY0ZHEg2cestcwomD0s
B0p9b7jJGkU1TnCANlxkZv3GCGgA3TzN8inRanZr4yG3/AJCrZ8KatFwh70Rrnkh
QnRuyl8Tik6O1eDB2+KR3vaf7myiixwrOh8Ae8XnSKv0LWzUJqNRVjnGxRl1Osvg
IFWHtuIZDDLdLfz6iMfxwcMVOeTC5x23Qz/LjzUBMivrfbY/xkICAB8RR8jNPcCs
00fagAOXMJTzCeRwM0xbFA/5UvVXGSvWPsStb9srl8TT2Xkfy9wgu3xjE74yl/FO
sxMIRtCT7SxI+1GEImGQJKRPVt+C7y67kpDp9qxaj5AY6eMS9rxxBb98qh3atppe
FpiC2zE3xu0LQasDzHbWabJparVPhfd4ziQGwqEd9i/oKaDs8hQsMKD73eKb6tKG
frFcBrjGVDQgF2t8lu5w5nN77JbxS4DO63FTOESJg7w+Hw9iAmk3t+kby/HQMQMP
StoC4N6NPGj9KFWK65nSxhad4k3o1iSbC6xFRY7V8oaUB4ix0F6i/UolqjHuyjIy
EbQBvWWV2CnJjVsl2PZTY5DI1QykuQxVNLl2BG86hKf2gsmk1z6lsilXenlw6tKW
IWZ9VNugx93ssimHHc9epDnNa87PfFYDXkTLEEQIRRd4eXMrIoD31K0a22Err/ob
lfqyprekv8vG73oCs8orqktlWbV2iLHWSWNxK1pkWYLvLwmDkuKiSQSxij7mfT+v
Lx6Sv7wNrXA+lqk99lws5H1j94YsoJq9V6ZGTwTS4sAROo/e5Ef6JBE5S2MW+VQN
6JHWHcs4/52sVJ3nMd0AD6bcZOXF5pQNvpiBox7MLDCwDQammXbwXR8bIjMmAwnu
98IzrPBDEWz/lD+TFgQhGNEOli0YlfW3gRBK5pjE2T17amfhEfuiUjX0c65Ydket
MMpCVJ5Kntvi06LChyA6SsOln2Dj7w+8P1KL3/C60I6ohH2sDAeC2VrYvVkv80MB
nOk6fuAt/rdyVMJjbaxwhCrakV2+9UWT6IRKHuacSnqnro8AMgk/s5mH4+eMqp0k
BV+X9M82LExYfmAiHtucEj4k71tBwze0YUcVI/ZdaAU3nJD+c/OcVLrE8BPI7fMp
6OZfkxrbXaTmzLy6iz6hCHYTdtbHnB4YnKlJnwTQ0MYB/yJjwtNk6RRnO8NkWv8W
kpc1SOAIFJYi0Cp1pPsogp51sBEnC6Qk3DFAyP3Ubic7BGrKlJ+7/Zp5TflnP5Ac
dSnvHo++pAoqKcvex/CRiV+4qR3LrduHkXQ5auZ1IPT7DxcqKFL/Y5ZNs8YbRnd3
MxZC5FxgvD7OV7dpAKp+V+yB4bbCwLgbCJ9ZyRfmjcpn9xfjzQKCZkEyyZpweJ0U
GX+u6W7sXYKqaKvn02cKKdtrVTJERaAa8ogA33HM1KSoVgM11VypiKHmJaO1R5P0
vnYluyirqgmcXJchxP4xbcE1VUWIue5arvkvXnSSx5NyrA3yMZicn3Vo0o6psIoW
9LksiPHzGkPsgOs2ZDWtlVHrOszjZfoE1w6aVPMJNFwl+fAh4hYR1rf8vr4yFDPc
XRv9MrNTb2SsKFi/H8C5vbpWguz7jmFuMrGPjwv6cXIq+OofT85Ms4DYxAIl5uu1
0BRI5gFp2vwlt9uy2f/Cnzrt4Rn33FbnTgOPIew1gNODH2S1bhWdf4ZAbUdSgRPq
Ff5jALRREGZINFVI144Sjct4tk4jqb9lKoR/URMyBkk8jXi2Hw89YRVo9Dk/m31/
Gp8vXyk93fHUubUyJXuQVFJE7ckritINwDtHkAEQjpV+9umMbkpF3vXH0P4VKK8A
YmryMusGP7Okq50WEgy7BP1PZSIBEU8Jo3JD3DZqdH6/RhRXF8ExuslkzwQn14NJ
GjHMvOmsvwGuDuev8+p6URQbE/L4F0sJvpqnCo10ZhpzA9HxSCkK6rCleAeGmNmp
RFpbzsYi7lgA6qmyyUJNsiGBF7VJroRZoHtSlv8O+rG3wHX87yEHDzMM0/S9Ks0K
1qraIPjjaYF5zJNsXeHpwanUSnX1Zr+AziXFGp3ni1G3GaVdCT7LOxPxKX+HfQXP
wCvIII8WL7LVklTpyefjOZiJtwR7NB+lsF7HwGWys0xRlOdYXSiTdkh9alWmhpYs
A9af8VcKG+k05LFqRoXbaMLsOv+mtPxBFRIhKcT3PbLciM++j+4mKx1bQ55Oijfv
4VC3buJKWpeV5qvQBUkxbJ93Sa/6ax5C4sRGH65bUhS7kxKG2rtDuaC2B8V4KZqZ
xm0T/nh95q0beLBCjHcULFBr+GgN15rwZLtiXkQu9XSPEscV3C2Zy7cUY2AkdIBy
Z+pXXEz2sWN7ufdQNJGeD0iApFdqfbjtzXt4l0CN5W8pa7ePOmfuW75woHtHgN8+
C7PtQ+xxqzu04BcbNpRNoZrgHQrivJnsaFzYO+4DwHjR2tURRjjxU7Xzy8FhYps6
6i1QXZOV7wYQeF9oaR7R/2/7sf4cEjyU4ka4d1SLPRDPEazG4hcyuGECntW8zts0
kPVUvPgYntS5KubmaJ7eB9xML5hUWHBwp0Z5AehDLa96XUFemaJKCn2fEqKH8hVQ
qrGfVxIgCfTM7PVHF/koUc3T42BEVTNxwKAvejfOY13mYnoAS5t0QR9HDw8LUKy0
gJGa1plSd33WppFrS9pzsfaH9nJwfrYphbLnSEIwF3Db0hA/HSwpGEnrnP9CHfgr
CtBZbSUp9BerxMu1zFSeOzTNMLElbeIuDuhslyKN0ayffUk2cN6oalaBe238VFTg
OCEvNA0kJqXVoDOqnUAVJJxvUkCuiGdVelsil4rTBauq1pY1EUB3Jqb1qQ/v2SMD
NKSSxNnYXoitw4URDtAo5QLu9HUFb4E+2/r3M0Ap+9zw73I+odsLlk5i9HYpP8+I
ePlG10kPHCHhkhxSw3gHy9MLUDD23jpOFOKvYNFxjWFrkv/EBmyxR7mTDDD1YnNQ
RqucmFdfgP7V9WXjHFppj934ZEhbBFxLdj77zor5QTZLrafCC7/qKnOgBti6C9A5
6ZX3n7MK5SFyNNhSu3s2KCMwDYqmDhUBndCNs+n+7rQ3fhpL4IkAl+XZjUEkbcHj
CwhYqNpNP/EXLMyw4qXH2GeJGunB8W31SbaPWrNKfon+c5ioLEyXwgJf9Y53HT6S
Bg4BVvZ4rELAmNl9ueh/D8u4/KaQjFhO7Iazr6v4HMqDTRbmzyFmN2ARnMQoXDx4
LM/EJfUO3lDVxkAdejFimDAVNrg/e60hJiryV+8w+jVuVVfUpKe78NxWh1Grt8nC
rjM0kBdMiAhqPdMR2TZEEynuFt7uB0/TVzNPFNoVXHOUf0IXXegioO4Bq1ScFgNR
2XbiZDEJ+y/1NsgsZ2Oj4SA2a4XMqo2xriiMtldSHxrgR6DOOxXgdBwGlZOgVMwa
n4R7z5tb/2fW4VjOKoTj2xlTSqFr6anyWGQ78laJhvG65U3eJuyu9RoDso6MEI3m
DjqJ/9ma82uoo3X7rZYZI7GRpWdOGqkkPUFNTL4RK422uZlvgXtSH9kVKPPnqWy+
bvWipWRyvabYNKL/s1l493n/ebJMJnWVOurWfooq23hsJugfRqmHlLLu9Akl3gMU
Y+RY82P2/FBMGMRHrsHGnc0UbQiYJ4vRjlKqi7wuY1n8VGitvzGX0AqzLFtMqOW3
Y15hk6nDYxx+wlYNjL73B5xa8YwJR8N+G5VluhSRomj0N5PF+26Mbh6EWdu158Fp
44BbOB2T2B84Ro6LlFbigm67TjfuwX+qZLDTyZuSEKzbrmMM06JzaAAIpJXx8ncO
Vt8VHz85NZXMPZJ4ZUkOnXLLyBGJhVd8bNI8aEeXF54CXLumQc5dqQPsL52sb9S8
Bc1+kmYdT+yt5gKnvsmnRbEKJ1TxjdmkZr5Et7qSZEY/BVekNL70QGEPpgehERLi
ccY8l3CePQtoJpY1xBcX+t44OleAe2h6ma+h8lUCgJopbRZVvwZ5vP9laMEESmyk
A7/w9c8CIZLQCi8enf2tVvnQEGmJZ9UtX3CMbtjQz7BsDtigVTNoN5W7/aJ3OZzY
6HVQgERdUOmnRbdw4cCgfdw+flFarsuEu+tJEqyo/d2oOXvXW2uTMs+NfApE1ujm
rYH184Ug0pLmMP1TLy6pKPwB42isLLjoy098tusQZj4hng7+zc32bq+au4XgXJ+g
RzR0X8PJRw3g9lAywDv3ac/FHiA78XOMPrJwuZxTrVimVGxb7vCXuVo6W2M4wCzY
g30uLp7kztSWqyWIZGcRaSyLcu+GpHYIy6olDiDkHBRuojaYAf1lqYME2gXAr7XM
mg35b6bh8F31XNOxGa71QavraXC4sflnvobwxxEhKUCdLPDv3PJ5zUlxk/EG6LZV
sRLGf/mgX6v5JJwtmGHc0orvNAa9h/F9tREOHdtP91z+i+lOGn7lAdD0FVwy06LN
2DFb0xzqfHSNsurbLl7LT4Yuvwmak4llvzHZPNnXkEd21QEErmuN3aX7FIP9NY3T
Dp7t/1J0zRE1OKzDO9SPdMvFNg+5nXh8SG0sZv2L6T4+gW0ylge9exaqiQBfsa1k
GmRtvgDz3NQCnR/meq2WFgEKK/tCeIBhdFQqcvJPvyx2EQ0gpcFzpsDpNntrUODD
9uPhNQzHo+D85jZ/uvPKO+bneF5LNtL6RFSq4yLpxbQyYcR2HK+Y/U1kP72876SN
UF1nGpw6no8UloUKYnPB9GCE1LyjUScujazYADZyfCgj+w/B6jYAQjZ5zEZVvewy
ar7I122BLQipFIim+1ia2xBOI96E0ehhLf0GKWCDlOIOHYuB2j+5Fvr+tRpZThky
sIVNuFl1gmbJuGxUQyDLGz4epNqA9esDi5Gf593xUBfwy1eHPA1S//zYbNyxu3iY
7MPQeF9YxPjq3ohFx0+txq/fdVbY+4kNZonxTx4UWVPzo8Ye5nyZpo0Ej9U72j3m
0eNjs8Jm/EI3hqRClw8qHoA/2bFsH25svyB6Mi+aJTlZmigM7LwpLeKAknUabnes
Yw06NBIUyloDHm1Q9tqMiaNJZBm6M49MOOqW2dTh1GmG4Hf6ZjhgUVrgswg1TUah
c/4kuSO19KwNXfn7UwTcnQLYW6nTo9j/t4Pcsf1y+5PzwTDyiaDrEYTXFgAsMtT3
O/eN6bWF4Rpfq36hj8XR6Ms4JBaX6efLS+cRV12Jidxm/gC6PUnD1cCuBaPgni8L
v8T8Y4i5va5In6EcopfvVQp9YSzLvxT8HsmBtBH2f90z4qkZMIvKcnvKsGNsSQS/
LVvJGhwlY0OyrDjmCROVpU9KNIAdBpufpEI/xhqfpYz7b0BJr1DjFW/XOHkWG8jb
RMuDalArHEw6VlZANhNWN+cwXraqrLVCRHQ/t3aunsPQhZzD2PW6Ed2sOrkSQXSJ
0YibZyMqToptssXo5Gd5Yze4jmLNIzCNBkmeq0lo0Uzf9W65UnTjMVb+u9p4zHFK
BXtRT0ByGCAcvvr1Y/4xojyIww7pM/eFiKArMtvj7rxp+6kcJtDVfU5aIFYxOk8u
j51vOOgRXEKwNx+qEvtkJffD0TBfDD5taN7aSoWdi1Dm4Wzy+vcdBi3MSQJuuiyK
LGHHuxTee72ss6fziWLo1Chr27FE6K+/it4VGi8qVJwSpgug9cugbu2Z7lZFMpEC
O0QwWeu/QSZFfhJvRutloNgX0XEzIkVPiV039bYG6dDZoozm/uEi46aTXhvTT11M
8yx5xyB3zN2KoyW0A46M8G/v6vYvIjukmIv+Qh3tw490GuBg0ImrIot8Ju4nzjLQ
E4rBRty3C87fDvV+zx7nR8erqfBK5JLxRAg3xT2fcPky3oqEphxqkcJ0XLI77Qsf
BgQ27fnlpKd4YcRhwIwlfYowxETWFVSn3ehE4xxdTapb6QkgrBW6xCEdKu5Nn1Uc
i5vfwS53PTblSpDNvX0PlJJS3fPgw60U2vgQUtWWr2eR22IkBN0BuHMeo47VEyIq
HiWvessDqvgrJvs5GAzQ42+83YFB4LjVzrfpMj4lrKSFRvXYcpMVVn/05UkblQIt
vaKsDZ5gJY4t+jHWDYz11ZmKuqH9Y6ZleVsACLnUQvFQlUdszutNVae1Z6b+n2/d
6vAQn5RYtKK5kdhRYkxQOyv1LRASwEKA0hgEUhRoejD+tMZl2MPdSHLgm2rC1x97
WwDhOgZFojbPi1rIuH80sewIjkj0ilh8xJRn0yNFu3Y7VJivcI8uk7eNcgrhp5hs
3lJgR7ZtLiqHBx7R8pTbXoFO/HZ5RdV20UYYU/8nf2gNx41dgI3OmH57XEvQCUme
7UA+mnxyqY4phAahdR71qAXfBQMCczV3EO2nzVip9r6BtyPNn1Q7/upqWIFh6WDj
GDYUybQkZHgM1bK+RfCeQL35PmUVcXLffGyDEoiXlmH5/ErVkQ9hmrQz5p0C+q64
l4yAesWsmVXbdCZDEU9FxbDaQRbzFz1cAgqj+NfBtwrGaxurideEeyzPmY3/T+9O
0je9+NO4xGLZaIvVJaf3PoG1i7sXllTBmZA2IEtIfBiQTFpEXc049sRNGU/NMY1A
E4doA3wY/EUWZDxq+i3UV7+ked5wTy+cqD6YvHjqLfjv3XghKIqmQPDsUUuWoXrv
LtLDBHEXAIOKHKyXq5fpllVSO08TSm2PTpbvarj97prhVsgXJrPgOxhrbw/wTfC7
+GdUohAylwlyIFtHwefne9LRBkCdiGm3d+AU/jTQGrC5Ymq+P2Uy8tkv0ThhbGm8
lLRpkPcCQZHQgvft8Ia6fwxxr/Kq1iVo/PPoX/Kf9ywFgEYx8epDV3ShbkBJzfIQ
usq0ZzO5H3RDfb5BPZ5eoh4DgUl8zkFZZ/+jI2q/NM6ex7I4IJSPl+1T04vnayok
AzVEhICJyT9hN65nfQAAGtQokwccZKgJwuMDprRxMXD58MtakCFIhPnXkAGRTC30
D/diPJnvdJmjqJRqYhuOVeEKFA5Ul+1keNsvCNTq/8pKMv9VHHPeTaPAjY15Noyn
9kZlXZLi+xV1um5O2bmCAgmI4NBmpIw0Uc57gL4M2P/D6cEir4DM0WUuv7xgAit3
/GVWiXS4nb8niN6dvhsNETW2XBFUCyIseVyoA/kP8f8ym61SFQM+3ek8UAj7/Ke0
kGl76EOVpvBK8f9jFLBQyAB6STUlyWuHXV3N5Yb8+g+jWd+dHgf+MXIP9s4qirU3
fKx5HM2MHcE2BUA/6eDnhNdV+Vo2IL76igdJSUvwk3wOWd5AtTi+vAcg3Em9irrr
B6+ND1Nuc6WeBYsYU5PRaeWiTVIzIvuDV+A8vnofdSty3ek+5ZNCMJCF9tjoqlb0
r75Gx5mg4t5QDG20bEq74aOoSwEP45X3r8OOTN24FyADasPldUNDsmkyPI7RSJAx
Eo/3KOE5k90NOg0yrQAMx3EnnPjjLEmGqJWVRCeDuof3S6TceSAPN5cZue8BpK60
k5LoRzHUMjvqqQQZGEbpBFwS/N8lVxhHn3HQ8bpKwfpgjUriAxnQ/cwNKRJBDJKm
X7b8z07qxIpmcMpSSF3irWvrl42VHrQWkaQxO36650FRHRy7/v9OVZBsm/P7jdvM
bQ2AYUZC/VAps1HGWpeTESY2oMZgyAqQPIDMpuLUB7yt7aBKWVmNAFK4rvDOKU9T
t21gkE7KvzB9ydLbZt91uR1y315pQO6OlfP9A2NCFD06I+ivtRAaBE6PNv9qAms3
N6zxCudb6q5eg4UosdzIAlFw1btnJuV9g/8hv4cknpLDhGT31evqrZKolS+r2PSr
UvxDP6eXNo6WSvyjWLYRidZVn+injSsXdz13bla5UyftaH58006iTeP7QAHv4Cy6
Q0hNG5JrlmNfmKrmH51O6IIfoBZDx511MUeW4r8nivWGKfK6Q/tthOleqD4VGt7A
zUTMBl7MbyjOwqTNE3azA20sHwmc8iwEw9c0cVxc5pGYmCLVT5R6T9nLFn1/sZZg
b17n6p3IGmfXi0Jyfq8ERVYnKSP3vd95LyPmosk9q9QeTsTq1ahQBaIGkfPwm+K+
fWY4rEtm2WXoH3Qmw61WnVx125+jqjFv0O2CLM+NWhMgI1QQhMYie/1XRtZ0Z4Nk
g/wwOQ0ZGheu0pc0X5CTVy/2ccjgdDVSgTdGS1T52IC7mN1mZn2LMz2UQhTWWc8q
zxFxjVij2O7pcIQSy9IzYA1v3XMO/FBfnHOPidwK47ifcd4xuPc5h+otV7c2GRur
qduFIbqENeqPRUvHPqdDmBXm3EGkd6wi5Qx7wdOavwTr8tVm8OSFGx6QmOTMF1Xl
K3lnxPdgGlriicQdNfBuaOz5cRtpKd+YyxSs+b7kHpVV94Mhur4+BFX/yYlT7FJi
PGnKOFbCkFIsfXHG6gLHAJst5Y4z0gN1qW+NBI1AWBnj9Ew/AmqnYnS6rp65FI1k
HaklEC/r0uOSffinhsPGsuk0djPWWMviBCBMxFzTrttQON7Fb/pANpzHIxohj+/1
ToEdYoHBgLFKdwAPzkhc9jSjemRTQQ44w3cwmihFCPf56RFigTO2k5AdfMcNaJAm
5vm33l9gnNwX+APrxx0HNy8ROFMo4NWXdnVjyiO8tOwkNlwfewKR7Brmybe84J1a
fiK6dAAnzclZDr8yJlfpcEebRFYt41VHGYXwh/pE6M9A0c0quBpsFvic0YrbJQ8T
Vay0J2yg7nOHSThj7yR1oAnATErr5Jn3sqxJexGq+I0W9FFoefyQb8BMD5pMkSfS
A726iFbEu9zC9K+sIn58J71jjjmOpIuJTZYpBUfUPG0nwD79pevWaJe3W+wwv1Ze
9UIFGVPnplI9okbf66/MrYu82HcrvGs20VpnM/zSbSr3AMub3yhPyZzoScC3dIQQ
PmFoLGCEm3T2Pp6qQuMEcd0TjuofISfo0q7M3HXSwaJd9ME7EmS5M5G/tTBoCVd7
Uq+wuT5vWMw6fh05GkQaUZz6B7fT94NfEWwPDqWjoRhBRzox30hv4IPsJnMLwbLQ
YsuCjLC7IDGfJvMJlhX4rO0Mg+ytTxl/bXgIDCi2HXlW56M8JVnFzPa9ESZvCwHR
t+x9+Be/JqfRqdpTmuxYU+3gUFe6Pewd8za7EpJtvF06e5ON9BZSe/uP8wmFepEQ
MOLIr7C+pwhqTLFimWWqF7GVLTusiwACet/ksh5+yPXEctfNNQMakIuTthFp/m3D
j8WWn5F+kJCinBvXwbeMFI3gNkZ0ZnIfh6egsP3u2eZeiSuLrD72CrCvttGn99AF
DS55MewKneNsTBlpDCSkSViRcjZcLcCkgU22W0TweOKZV3j26B5YoLtGgqParRmv
E2D20gxf2qEc1DNDz2URVheIENmKgSCbzv20gMwvJYgo+o2u4ydJUjTfpQ9ihz23
mnSRaf5KDi1dFT5unlzzrow057xvyr4dZ9Rws4UgU/iRacOlIvIS0CsAOD6hebuw
Q7l2GEPs80QEnYwOmatVaZbp4YVlgzqOD5p4bc2Y4sXusIEKKpmvZTNMhgtmlWPA
lJww8maj2drWp/yzzXT5Y1t1NfDpUhV9Jwp1omEbuPrU6DT20EP6JUbj+6v4dcxf
IHTQoiu5FMKwdvg5b0/pPzFTn1qjOhqso2bA5Io613zX2TqN+lH64xXCmE+5yhYY
8hlOlDwfv1GKhnFFDzH83yY2kM3vbzQysxN1XPIagfpXJVuhA6koHXjiEpOeKZtY
JVY6jtgVtVgJOJdGzn4oUPTqgLsVqsh9s7lyMoomQo50zZ8S+8ZVyLk+bfxJhiQU
H1bXSp7lg3Zv/PGME4dAiSlfMAhPTVxle+hch4FJ6AvzXyT348i/GhB8VOuBwB8i
O/+MnMYSUdH2N8M80ZOAicoXljPcuM3RVTGhtEp6iWcarz8DlPOFoqRoOLNnlK4A
pceAkbWhpf2X10JWmW0W5YkBPiKWReHLJkd6QsInFiPKTeH5L8p+sXn8eL0jmMa2
Hq/ZV8sr/PNEgJM2u5zWFv0qM7ZbMd5vhdtWL5otIaGl0HTEFoSoqmmqw3FUfjWj
1ceEed1vZa72JVj6cYoJBGuilAAfiqbvJ8ZtTxpu+tPdwTqJF1pyQo6vKHht4P9N
tHCr6AC+mgncfHFlSjaDnksTLr1awwRIr/RDbK0/Ife1SNJr0hQdzoY2o3p+9mn5
HxquHCAAy4IQNAeqAWlGv6vWM2cTgOIe9AT6jx6LnYeSsGPsmMghMDUvQ3VgHzUP
PTUrJVRLYThh9HsMIBhMiox2bDtc1Fi+xOxk28R00t0AfJdszhTP/2ghXy1i9bKa
nihPMlU1qiCz63i9TSVBUVW8AnkF5v7n6mBoBtzu88kPKJqavXLE/EJLFrZB0Uty
5zqZRG4Z+MPam9OW3e/Uo/LnCb8ZMOpULfttdMFJU8/ZdmBTHyME+vm9IQBBBANw
uWxWdE08T8GCJ+UDz4tNzmIvhSAVLwI8WLP1+D6X4X2it9CofEEXK9sMLQ2lhoZp
YP7ui1xsPXwplIe4YAC48NsOgFkYK8bgx0Ubtg9j/JpJgZykrkHXU/tG6iD3ZUkR
eiujEKyCiFBn4bQ2vkxoA3Q+e/QIrmUy+UyMCC34DDPhszI/BWz1FXkW/GuA1xy6
dr4QI/8VVeFV2U0ogZRx0nC+7MkPiZuhXk92A5/XoIKGmnipJf/l7OXOI+zYJltq
QsTnr2CCzbKmBkfT2/H3cPkR1RItKkYTgVjA+lQGPlwFBkx5RK4+kVjYKPvY179o
z47vo6BhG3yOmAW3su3QJhpJ/Co0bmminKHjYGpKWJAf+2rdM2U4wEj1jcvy7NpW
7bz5fLovAXruNGqfIfCXpDARXYWKioJbrxnUh1wl87QPMhD5uy30vQvQOf9ygSrF
D4vw6kkbbd/rCo6AN/J+cR0kk6JWedK8VRQ6u/8BFOcuoTn80oSH3b8qxpVF4Pjp
ZbbtzYLj/fvjWVJk7LXfk3rayf5ZoRsx/XjGELtZU3W9w+0av2mHP3zbYQ4JykR9
VZej3OXBcrtZp+ECJblglhvcaCh89S+ZW+G7Lr5URUrhMLeHzuffxwrTW/m7hWqH
xkus7JTN4tnxe5t6a3bLNuCFuYhfxGHU7F6+JPMETXoIYgHJmE72UrTfoAzvKVYA
yeVdfhlTxP71qc7VS21wfy7Ok5RobdZ8Sbw2fmjBTVzZ/1unkQha2fy3IXdti6Xs
llKVkqDb1ZoDTNYu0smo1DzAabB4P9cC7fPoTyP8jYxLYk+0GgNXlPfoBZVgk6uL
vbWM2uTapWjBAwkoZfIl46e/t7gIThMqHIOEwUKY2Nl2Gjn5iORjdOYzKD1U9XZ2
i024dNidCwGZ4Vk0kKnI3E4tHgt8gwGoZeUKp2ltPvYyHirhi+c+eTC3uL/JBZAe
1/7BDsD4NWl+FtqPiPGTbA/srJs5npZcTbzu+YDiI391IyL3RaBuG9cQA+23gLNX
IxMf/lrIri/IupHz+f8VhcuTA6D1r1ZdnlN00RWTVaGkBQwT2BwyDdjJ4juRkoLs
IBD4w4Daoclty9Jp90vSSrkDYaqWzdIjLTpKjciFs2IJYCYzH1ShAf+AQEqxhMDY
lKNYCDFNQjxxITyx/AOL9QeSfsNZwvkkknE6VwMTeue8Lu8xLM0ydeuzogIhw0RD
6WDKvKV6vrltYDeHIhsOqhzEhPsj6Q091CSRiwCX3h/dbuRvwBeS1Eub7j5GyV06
Mh560Q27iaDfqQqA3Ql7Px/sfnX1qW7mV27u/uRABULp6Se2TtkIqAnCuFOWRv2s
l33gQ2eUruMzds6Q7UDEaJH8qihOTIPdYCDMJH1V08MdjG40zGTLmyUMeIcjlh6b
8X2skdXmgqqBdC4/92qgctHugcEsluHC56bASkBioMlNWrk95AKjlYt/Bn+xzgX/
qIYolSIH3WPsEMmx4ibs/fqV/S+PWpYGJ7nIy7XB96YNGegAdTmweG1px5Pw4Cad
Tt43m2qAwqC+uVdONoJQeXGGVUpAH6Djp9H7lLfAARs0DaPR5MUXfXtW1XpF78ci
8UptWDvwiy4WkUO8fE6XEvKlt6YmhWSo4qP8TsUi3BrvMF9o8xrYRnArkxKW/7gZ
bn5Ub8IKAhAzIVdA4roIXmQCVs3oaF3R8MxqdQeDWC3jfeaFo6AvTDZty9xzLtm+
9ZyyGnykV0XHMwvpJEeG91RuOsXOSOsF6UPl7iaWM3Ipn/Fo7BWMkt+3yM/zPghN
qlEy6nBLJv8Qn8StHCKmVS1PwYtj035k60EI6Xayu+AtjVv6izU44yMZ0elcqR+Z
Hhusl0BIBiDgwh2wMVDf4TMqV124baiFV7JDK/Nk3XHGlFiWFW5soFmA1zMjP7nV
Vo5OKFAEG6bhftgrmyMYanGSAmPX6PhG3XrrV4e+lC1UFXFd5lD+ZNm/gu9k4cxV
MfhyE69S3TMhYJX64r+D9ZoTWFiqUSJ8o5G+tkQ53q6zjLCegDkvnuqq6jCEFIEw
hfnFR+7hKmP1d8N1S+qmTqWG8LsJu929o+SVg9ci/Mp7YYBYt/nUzYw3+6YruGt6
8jemtKmFN8GAn4uOTVxPnrX8LeCBKf341X0zjC3Y3nszwMv4Sg3vVN9cssGi+1gO
nJnpzdVlKE5RvtvVyIZ0jkXIUXMj8HeauvViu/AP0zgj7w1WhdsK/a6nDO7vbIti
VYL0I0Q35LSf3hoq8FOLPdccXu4bdBabwVdoaetd0kQwg1z/GVz4cedaf7PplNPT
9tt3OvxFJvM518Hn//g2Hi6xPWjqJe6/h6F8/hRslitdjaqzHLNW8P6fpoqwGliv
+eX80kIM5Z9MFU1KPlPTPH4PaA+gJG+tOeLjBc2Wr/J+a0DjC4V3R2QCaICuLULI
Yxr+njJfhYMRhIbWKSwf9VUbitx8nHFaSLvFcdrK7C8b5RlBz9bsbIHv6F4HzZTp
+EHdDp+WKgjH86dWCTn6bOXJ6R4krBC+QuiSg8qHmiqy3FCrCeLuJV8IkDCSwcRA
LKxfInGxterv/PJ441wErm6S28HBdjCeVgbT7KjEShzn8TPinMtLBaRSRbMLSDz9
c58E/Vsw8pzjg7qdcdFnNhtgKJZXcqAVAdrCU/ox/xcH1Wb7PNl8j6gmRRY0NrFS
mmPb9EeS1J0cOl5znVGgR9oFfZ1b0yhDy1diqyuiiZn2NGhMUDRwdayQfgzAYHl0
K1WkImXYsissL98QtwvmVrWfPikQwVoryewHMnboFqZe7vzYEk4SCoPTRSHveS7r
/LBbpQ4bcoGayJ1Vci5P3HKgpQ/CBbgqpQCL9ivTKV1MtZ2DEVREJahXk+KP8zCc
qQ5jUnBHtCwthUp7Z7NgqAZFKO3pA/W5gAajNpECvcotaebFH5uv2N5rTkxWqz1X
5f0ZL6mjwOQeYbPrPKyEiaDEzScLzIMmWsb6jj8tZF1hPh2qv11fw4LZCXOryKm7
+Wsm4pvp/x/Msj1vK3ouQddk/3kPCTwLO5Jo3ocUrww1/Cu9ZmuUqCKSQIQzvthz
Wu2SIsTLAwAEHSw2+tLTJL5V4VyVhxrA6QSH5dJwYjdZYI2dt2w067YpYZyj0lBZ
Q07gxAAJNd72bZ7SqgqbB7Z+qTL1IFTRyoqr5wBn3L4KgR2vQfS8/OyaOcwP2QhV
IGmtyGTcGnS+GhqDKXH10k19eTV9Yk3wlmkNNHsUtd/1h99BMQzVipnyPrybKxKy
5poHfUi0VlHiKprBXnO3Mgtn2sHe9bBAJeCtiOuwcRAVLzmJyVhukDW57AuUUbHb
N9dbRJ7UgnCjuoCMZsu+fk5h5N60kY/xTkQlEJsvAFaVB8Mm8puIlPmK1RGkGM3S
YXobKZU453UwvN0dp14MJXGSm6CVZdz5Yo7khqp9NJ+zgTrStBejoIVQ5fOfGLZo
5ERzDQq6O29VjwQ1gqgxU+szEVwTPFDncn1VE4SownaLJnq2cDxhz3/cdVqgsa2C
hzoi1yWqc137mb/92ydx21wmmrf7+lWkQleKU3VDSp8/FBaR96gf6ov2miBsbN1X
oi3/x6lnzXJ2W8n/Y9DEZxyrZ+BNQt8x/kydWizT/7SNApUxWgLDWKLyJJjEUDWn
P6mXACl+7YOacWKMXUyk5zszuH7UaQDFmwBTa//iIZyHBmJjrVrljfjmwyL7BW5/
7w3CQvbvXnBj9GChKWQ3r+ed9mErwFyeNKB9oTIXGWHaUEW/rT0MaUvMEEVatywG
KysGzJa6gjMre20gZiUdluwTv3EaPuBxSyMaFMiJNtArGV7I+C/HenUJteVCVRSJ
zb7om1LzQF6AQrTEaov3mp580UATRx5dSRPe0yOkWxrsukiiD3PuduGL2y0VXpQi
NZqpyt/jAWQAn/R1LCevunNEoUDqSQ3oPG5M9vE3TQ/lamraeadd+amvW2Zi+LcT
640IHhp6h0w8LecPEu1VDkHVwOM2bncR4Wcv2cnZ07Z+bWQUUZwhuvGTmffKhPO5
TJ1TnjWgbdov/nIfom/bxhlPZna8P6/DCo3Gb+hQO8cDP3a8ex6BbKikn8iVhmlO
tVgA7HrwOT56GNWl1xfCu/2+Pp05MANgWY/lsV+f+CV1afbjcCajin1fTcVq+D4W
hEQ+uHJOSffLFkHfrRd6OEAvAxNRSFYLhTyOaapBGAhcO9sl+LRKWghQfUR6dF92
1dgbIgh5JaxX+DaqYV9odZYecofE22WGJOoS+GU/zbTbKQTPpH7gpGh/NaFJ8Hp4
NDPo3fakW4NkwUA2+Bo4027arPrlpWRJUmkMmktyrLsOBR+lpHR4vPhGyD74HSvX
zvJ7RtxR8xh4iPqziMN1NImen66tkWF1B3txzyKjKVSCmcT+Jo9AySZ0+P6YI4c8
q9nQa068ZkG3ulH2SE7IAlLNKfoIp1CCUemSGZ71aMTlud8thqNJUTrPrcxSFlCP
NFr3EV175tk2M9f5xRAyKO3k8yG5vNK6ZohKaiSoZwrW6yrSQfaPvQlj91f4AwTF
R0fJ1AhqSvrqpj8d3mxmmj0yTdOGTljmcpVLlJ0uH9wh+EIhNp3wpVx8LHcSc1+p
xrHXz5YlLjc1Xv35x4wtei9eCa4DG8phwXGA8ErVlpC2lHpngN8MnCCU+BUYqUqr
dGtNzr7g0Ny/u1QC9fv8PPN4IbXBK1N4vpIvCY8KZuKGEF/wngg08iuUh5u4PMeT
I8wFf2gwKGLzTOgXYyOVbgdGjTgG6J3VA3eietOtn6Qphki8H9uM1wCa5bG0PKLI
j0mNU/dZ0BUnlB9AXbAa+eV+8RjoRkJbv432k9fuCXLOAJQowTRmU6So4idTVN60
XLe3EOhYQzNFN8FLshrkDjA/KiBWr6Kaz6cHtz7G9nuneQ+n5JPf/L0r98ORD2i0
7gYojME/4AWROtcCbaUJd1dxi9JTXdzScmyYcHu2RptRjNNLYRYkId3i8Amfo38z
hbctb83IWuSKxljexgKx61EVIVBYR4YbmSYcwevHCbhunguW/iY5XpS44PFaZDsm
NbYAKXJzRya9aMRO+07QFVgg0KJVwUe/LUgz8Ky1DdPkRekO8ipqDKrrcDY0pOPo
AYndWMD59WONEx41SSIGOhHSIBGDK5Xkz0c1S0QkpJTHNdC0wDw7ZR9PQIESdMrO
0QtiuNnsvziKwrSPERxAT6i3Zc6fcoJTYJfcW817hmSCQYBKiokQV8fa5R54lA9B
r3K4iH2aEbWflCZtZr7c64AInBhra8bEZUn+1mIJ+YrSgPrd6zREVvZouXAjiyY5
CexVB4g+kS6saeEiUjPPVxsK3X8TC1hauhcyfE//As2LZk4fUmfDQDocQduWKVFn
WOP52URdPEL/uqr9zxGHtzUkJVUB6fE/gk3laRb02U3GyNGQpE7h+oLg9sk27WC4
E/zlnko/xO2RmTnmnUqvirP4fKNn2HFczLRhjN0cMlOyTM3MaI9mZCkcEO4dFVsN
6w6vaGaNkidX85ROF4VrhAZcRg/7ex1UeDupPtu8rjydR0JUjcGq/P/RMcw7Gkjh
3H0hRMTiE0+n5duZdDMYahdFSkeJ+yJnrKwErwLtssfE+NDbENou/Zm7I5nhGImP
TCBTFx6jbtfgavG2hSk1QVzaB1CPWUHxey7BmL7sLZbH4Vz7MOT04zRM0LivnaWL
+7UVVzw61QREpsimL9G8PNmsxAgNOaLZJOvRr4k6siUJM7qRx3XDaS6aM4WRIL+R
vu090tvKrKaiDKCtji8tNlGwKG0qQba5K96qJL1yfbnxxPhryHBN3x8zGrC/emQ9
J8rOWL7XAC73sXOeb41deC5tl8G/WBfc3vsDsEYJt922K4yBxCb5ta/eUiuRLxap
5Rj7sfpFUNtLA7WF5vXLvtS6+vmxx2D5PCnlgU+2cnt43XvtoCNmh61iKCm5Un1T
6DSFe36/3P+WvKwF5iu982jKQCbwQln/TIZ+OXxYE//qPiLOhuDw8mvVnT8VFHda
yc7KgVLC/zi7270RZR2JMOrRrQO+1xZUA0h6LZFNiicpXpJ1D2jCO8SmpAvUP8cT
tJmdylhrEgBfum4gh0ulYs27/Bw5DA/CxYSDx9xJtzvVPt//EWhM3RdNg6Rmq43x
c5qa9iJu0jCt3BsrFRdFhaZrfyz6BFeoR4TyqgvKOrsnNQwWBAkoSXtQEw7U7pKX
gLLNp4RT2TiA8trKlcuAj32PiYvz1ZRoAsY8jY/gGcnhavFRBGNA/l+FwKzunk0t
RSVjsRttRM4/6sYOu7aRGcdc/b/FYDXKikjMOLc/WtHUiHNEblGWaItCOAzfa65g
80oiPcMx8jgrxaS9/jJ0xfuzku1jXXkrK+J7CjYRl7RIBMmTWabzN2Ctz7VvO/db
eruHDZYAw6p1s5IToDt16rfrULNxVXVQHmycJiAg8wvT1baUqihAbJd4keAJMJBJ
ymz+VcEzn0vigaoJeqRvM4UIpsmvDsuUZrBqPMhEuYsKI7Jf/IlgYSZ4SpmK66zc
Pkz7RUpg6KEl6/Lkw0Q8IAVlIhAft0P+XiOC8s58ViF+PUYzv3p2vBe8VFl824Eq
Zk61LByl/rjQ2rZj2p91Q92RSQyrtyqVnA1y+unXK7nDuKa7xyKgaXIt7Np0JDrG
KNopKjtyrG0OpdBFLVLgjLZUmNykV1j+6zHZcPfOr/yUKBlzMw8b1Wag/gzvLSCC
2KY+TsHDaE3MtLYg70fE3uOf/QbqMnQXL2xAwZknJniE3xH/Z+nOXGfJ5ygWh+mj
L99k2SDJfbRgZPK1hOm0c3egq+ydXWIVMgJrCmy+sQtAgJWilYhJ7MeIc/5HKsg/
QJl7rd7ndxelnY+LLgKVeyHKnpHLaeb2KDYwF3eUCtTWkUPvGvmHIO/I8ed4sITv
LLp+NljbaFJZI/rKN1AjxOEhTLspQLogN4bZVd1pB5RhKPPea/mlIUemryU+4gnf
wfNnTcna/B7hADTsJLi9+J3NGFBYuvioYU3LCLJtS4OfLlz82Uya4+nfXrYtYhtq
3pXefKlMkdMMII8nuFsQ5/6LncSLx2645OnubFNcubnqvy8EGrxGbsxarG6No07K
xxUQGwfP9saYV3gev1nOZrdP6hecLdC4bRpOqflGy04Id0Io6MJykjewxQU/KG2I
BArH69MJrB3FBrjQQcMLcG8S/1SVQT7n8PiqqS1RKsVbEdR71ZJRjDmd4oPIC6SK
H+KDrmbHqF9jFLB/0jecvaBA07yo8oQAgC4HzMrz5Q2hHEHDAAXV6b0fH00TZ0ff
D59L+yKkj9R9oLtSZF2QlrsBx+7OToZrEbce19NDLv3b72KMXQ9OaB2HoJ5a3ctv
vMsChH/5ZobkfMhjhVPCpVJEyJDwvMoykKkD9DA608pbDXMwETTXenrHD98DsdO7
i8CnPdZThAbflG76mnzUOA3EKuO3WB42PvGwkGnKT75shuZ0oRnfKlb5+SlkHRgJ
y60/8zhzO/veOg9vxL15i1UCiUzovRCBzcZTLinSNfrNMsLyaL5W/puqPJ8/qgZt
hf2escUK1FpMNjolZVjVeGt4/stC+HuBXCVF9wksiHF2Rp8jdKTT5ASf2fCDJFBG
Xgs5uvf61X5KkABK6mnv5f2/6NjdVUMS+mJc+aH9jFNA+0GMbEfArG3ny8f1D81E
kLsFnvWRq99sIa34AE3PT6x1F72LfiYMe/7kTkhER1ZIgf4h8OZAckKmVSRmv+1h
X9gcse/D/IjQSi1bxizcvei97yRIOI+EPt+7XjR30+N2WINUzo3ylA4zTKZMWLGq
qOYHq444FKGxf1EP9M5ry+h5QLXAFeM4A4kOogIcwZlMD5shfaBu2Tu39yek7sGd
pbeVfv7IQ+HQbDCJsa8HRAtO2IaRBtE2V6UKz3F6dgid2gIxoB+kTTp0vgCeNbEh
066fGDWWCkkCQlHm+XCpa75EvcIO9QV/tEsbpptAlzZKLYOdNKDA5+F11vwHvGxl
DfRiI5tQqcAy5+UfYok0tzQDq3JCwMbfYplbTDcyg8oEhC13R8vpSIcY7dgInXVO
6eNFr/tK5ZefeUohaWBJK9/5X6HiE3sWaTWhnPRzNc6xyXzUqSLL6zJxUNfkTZRx
4S1m++GfATsm6N3R2iw+D+46MFqtY7pGiwKXa+4C8NNvlY6akvz0Dj07vGtr4pPg
aJOjEeskNzFTFjK0HX9u7L22tuDzHsFe24bhooP6pelAJBVTOqV5r0ZAk9q14UuT
HLllruqnx109Q1ws/GIT43pm4Vw3IeC1uAjJlmXH1WxFh+NVxkqmONNBhdH4WgF7
N/OnjBFsOp+6KmuoJSX5JD3Alez4qKxYhIzotyRFAymTDeHRbCPCNC+h1SLR4xWQ
okzFTTl9eS+V7Mr0WdtJTSCIsZcStCsP3yoiji4lkHtGXwdz4/zR83RH7mRVusTC
iXHlrGWi7ygjJPSzLzE9q5PEMSd2zFdoDpL+ad+l3Af6dRnEd7+YKlVaNHZgzVsV
X4DUSEKW4HypVQ9cJ8wmZUjyMQ+f8h3/amZBGxC2dTaslXWziuWjyLLs7GgQxcj1
YyiNfYqJ9ioNq3EC2qXp5JDT07R660BEitrjJVeR4iJI8W7GlSYNPN1eDhGeMey/
QpyScrJGjubg+AhGaIwPQyE1O+wyElaJLetWDKLESULhKW7VBKNvva+KIPWYBVgy
XhI3izHWhzwVrbzHnDk+Zf9otl//L8Lzawhnm01ZFMEvvZvH4E+lSzBYhUarx7BF
NSSH32kCHVoPnINoQezxU2TU4LDGqjLlN4+Kiu1B7yBd8FIqZwRhq2dnbxW2/OPE
HxdUasnojsJ5aiVXmNi/+gbuOAXJBvIckjPDXsybABzrrXZtG0PDly/ieZxvKsVY
4fPGto+FdFJ6jXwg2ZZvfUKbvzU4s9k3Nd7hcO7RWkNIdfhFUluD1eQH9qc1obUB
cd7dAAhCApOOiTDSpWefVnaHS7/Pf5Omu0dVDfCrxq7k8LNpLcBLEhXq0lyztO0J
lPwjwLgrDtxMe7D47NGLwL48iNl9R+O+Ibok+fQnZ8BIx7xLLqeXK3wV8nK2zr2p
zwRWzuJxFJoxTGNW7VQZoGFcoHIbzIoBMc3sPs6+bfhvx4em04z7lGj16XbvpTGR
EZa8iLMNVdHQUtCrkSzSXJ3mVTe95HtD6miwvRPY2OcgiRTuoXLOBCaLQy+ggQXE
aVK1Afj8koceAajgEVsERNxBqXRwmxnJYQu+IfkuN6jS9gEyfTL7c2uYfREDdTvL
8UfWXoJ1sfpzmlQgn7Kt2IiHUDDkhRhrYr2XYDCM22dPq92+Dq7k+mDWHK0aMgKb
1rN1Lv+O7zSL++ih5Jhlflnk2ZLpWDBzPIvX+FEQpidOV7LEvQTf3t3QsWz9Baxc
nOer2war42/h6su1e6EEq0yuCqYZoWGRk5JvbCz19fWYstUYsQ4GJZGNd5Rk6AaZ
ro09+AQYygQLCOpyJkKyIrNZGUdgCjMSXLoS4iuRJ6suusOTXdzMDwwtFzuxEWZy
deOV1x1rJiZNXsV9y58L1xNlTdUkCPTAadtf02CM4E/oCz+RVBsDWqAplivdoF6L
dK3ODZGbxj8dz2ypmUWyLpP3nq5BNQNdQo5wkoEORHEiwo9QPaHcNn60/gFRBmeD
yfaXmrZGB+A0AWcGfntALo4+7OC7GwcNBGbLl0aqwVJQskqjZCnVZw3p69wyyCTP
pBwBneKcykDe7pdNCUJybzfq2SC1hD/ejXdvl9zQk6L5SheucQGtsRg19gCMBbDB
AZifSwXpVUqAB53znfyIzj+YB2K0ysSXNsHEt8QcRN4RXFi2nks6Qx2nzGf+iXZ7
Ym9vN2yX+ixKpbHR5nTPEQAx9Ujw3aOTJmcKbQB4MzEstg/giLgESxNq+GVNxlMV
KD/s38m6+8ykYJAJM29aNIa5JVPQ6tYwmMcZH8KKpBgtyXrFY5ztp+x8QkRPSbiP
sH+3EW94sO5OXqid9XXDvh9QyRZc+W7uhP09FJfv4vdfvsxtGb2d6rzV7STXZSTU
LChiiTvX1d3oMhAlXmds8Ud+4lR/uF9jnS1qEWWNgU9/dYHSOiehaL1+/A6Fjlnf
alrlManKyEQ+SA7vuQQVyypditkVS6DhEdpMXmwBB6yXoTl7DwEmESfqfU4iZLHv
WwwxZh/S39XbEmq+QmcwouXZQhvlKV0hMGVwI7QIUtB7aKeCtOzCD0tGuBVTTuYy
kFevnLX2jTK5d/n6dE/SFL7egXvxAle5m+L2UnIdfyuAL5LyZ1ED9GJfKUkOnxPI
7+rAk+uKr/pMr2VNsc+jbgK5jT4s8WtE7gRxMXbYctW8qjUBTISVWhbyljOI+aob
hVXyIEy9R1NsgXYjl9QFggFLr3zkDODnuqqHdCBzlMsypM8jQHTE8i+z6nnobbiE
UjpcZRRMqsXJn0riZR7qU1BBBFzJPUr1gwhaBsgIzJxXezYolvuqyiN3OQCnIVb8
RQHzMThfxzF7WuexmYMDksvvwzq5Q9OPZNO9z/9KF2djFn5Kj/nYVsAFkZj20YVQ
5IrfmiDS7A5KzWamtGdQPVyfug3Y/L9lQsJ5s+tqQT5J0BwKiA5QQQvxBy4u4ytT
n2vVB9zksCEWJqxbmRWprH2sxaXZw0kbgWqXhqxWFvp1CwLB9VHEFX+ZWSU9SV8X
PaOMWNMZoch0sepW3NILLmjEwheVqaY2+uyMnncfWyTaW1AYbkj7dU+4LW6iTW7u
mnNvh4na+Zyp8b4IUAWIrgeTllH0TwWcnkt2anE7sFrQeUtkU60Hw85Ksh+7bdZj
aWk3glBgG1wSycYAEsmt5UK9LnorFFEYRPnscwJtjFg/bN6QgEHzpKF1AOV8OThR
PHl7M0uTa5b3p6diI+t8pLblfW5f0E8z3W4eYTWe8PXCs8kBwHOrcZnd4spLex0Z
4FeO6kOlsRhBwUechh1kSMjXhCgRoOcFqLdDD9Tf8P+YYAobnBubW+siT+i3DsDA
QKciSunoiM7WIOwEyIra4EM/s3g1V92M/9ZNzt0eYtx8M326SDR0fKeQMQ/fiBEb
gV9woU89XfkJ0TgfR8zfzbF0ZoG2flF2brayYmsNoMaEwRuG8lDsEbqjqD5dxtPZ
Kbr/SlJ7RlCg+1MHuRL3fftiJ3ZKFtONcdi6OlqK0yvmPlcyIuL/PoRujqLkCFmB
1282JTbCe/4C+u2Uh1Ni4c/drYmin3b+IZajTW29lIOXQQjc67ZB+ND7gAzN5z4t
yndH5N6enZXshewAn/IIFjNy9IQ6qPNVWAzFtBQ5/xEly8k7JqPGFMmoMc7kBlXt
HokvU4IdVwnawCgPXKqPprgF9wbla1F/1FFtQJCmFtFcpBxYZzG3cY8z4g/qZzvG
wRi+Mls2w+1VsBrCRC+z4wZD4KbQy44UTda7cQNBBTweBNTyd+j01701XHWClPvi
iuCNxESLDh/KKPfg4piQplenFrgCvGJIY8xXP3MqBZNhIi1o3eUFlx+CRjG+waQg
V7zgr3L9Xl7QgR2urOTe2YO45FK6l3LnxuB4csAlYm59oPyaQ2xAkHMNw2JHEjHY
+J+NfogAO2XLVreI767TOKcu0hhU0MCC+H9KPOO5CsPgh832M34lRxlmhk4Iy01O
6Ezkye8AzCygmYWM4oxE0n+fCKh776oxs4eBttkYYS1sa8ilDoXTN3QSnNdARYOp
8iabyspaNdCjYHpDIgNO33fyMLXTr5PmJ9ZyBPvsi0iMgJh2MogcLv478FSM0UFE
RpKOgex7lLlCjZwrF9Qq9S/4giZxBwysc8ple9gGjWwPY+Mnag8eT0wQkNPFygQU
DYWCt28CiBnMOUclnjzZtY3r1UN9sFbTIN9ev9uxNim3BGeTqemaHs0hJVgeJfmM
eMaELkufIcmwd9RjcfRnS2xdVylzQ/9ffAjXvoLFDb8BSKCOf8lhlKv7ag513QUK
waIiwkJ/57xBJ0wRTCfyMUSOyAoT3PsGR2Pk+etysNy8oQlA9P6T+2FLCCsw12Ls
U+XqslHE9lznE6ZuFA9MO9wvG/p4fTsOR75xThg68j8UBu95suvb8qYrpqi4bzfp
VPz0r4LjvYHohxWRvd+E82F0oXoL820MQo4pwyJpDXT1DtnjPdcCfxYW9ZOWQ+nm
omE4tp4wqOmOwbtFo1M2b6a8hHAt+wgfkMZ8rDKCxywEDOqKPHOysp0LS8XWSeAg
mWz+cd2f7jeCrzu4jNG9LAplXeDEpem7PHjsPWJPpWyw8dk5Gsx7CnHxl9kI9fzG
AEnGKOVaS48WqkvzxxEGNjXG2NzjeIErGkXg3tq1cUY0K4W9kJ8DKPSrZAqxVurz
d4ip0XNV9OLKNcGbetnEVnTplyNxTMTBM49ieyXHGQ64yPIv7o98IbNNB3dulCtF
DDD9eQ2D5UhoFUUM4WyDCDtJB5ogV9jReRQfZLJ5QSZWsseIfYHQ2RpyqaBnuzb2
D+AVJ9HnIvVZi1/0TR+TWWdIL9MitrvYisiC2t8dU1N6gL74kkzgtHj40gmG1Ew1
yYmjIBGXNh1SBXc6slmCicAT37XpyQhs1woj+rsH2x6pz6a6HkYpL6ldWHvyLMTn
khF8XWTUoeR1uqo+k8PoPNlQoXwCiqrfzQuky1ieDoUWVssUjm9SAvru11yuWNCA
fp4nVNw00BIRGeppCsxkyrm3UplUHf1Posf52rRRY06BuvSwUzEkObBMFZKiFGjA
yn9dByxgaBMqShm6ttlyutyp9dBVJP5U5jQFC8DNG+553vXz2/8qjfNfExcAuU1f
6vmyzEENby1LnJUCN9F+cglCYnvJk/6iE3LZjkxYadTlsHCRpf1V34iI2pbaoU/T
2KC9jaB6KICKReTcCOniCcV6HeibBPrNDwKStsBKus5FVRzDCtXg9dhatDjrp4ij
2nocrE1CJm/YZ8TXVUYVdp4awS/TFppRIF8wvyN29T3/IqL4btmg367gLnfXidSJ
tQSPllZBl75rUi94cvPmfHw5GjZZMunGEAOSa1Q8rZxaj5B/q408N4unr+n3Pm9V
2+gP1ps43sAvSk/pMjz4sObRcRMKEzVv+RLeUem7n0/JQwArvI0tdFeqVVCqtGAu
hsiRPdu15wJb2XtK6fW0CSO0rUXTUxbWEAixMXLkLwAlioIGMxyByK/ce1pnMAf4
+b7JX2CIK9XlEYz5isAsv9Edg6TRJwieBry5Fdvkf5g6Eqv5Wb/WMSVTOJqOBa1e
MNxt5KRdf0zQBdX/18WonQE4JPFVTMzXoRhHKQEnhsFdVwG7QY0nwNNaanXAjMpN
RYEkfdYnf0fp9fVrtbI8bX/leIoEzOl4ysLob+YN0NRn2h3MzxiuZPU5pqOilP5F
s208V65uEW5L2gTmeTDc6Oo3/yfvaG0JLo7bbAjNGMFj4mYvW98gKwCkiutmm8kR
0Lx3sLi5s/2ir5M3azyf4viUGYuexfMNb1H5O2CufK6dQoqsrxygwP07Q4EnC40U
dKds1KDAogU92yScRmiy9bLYsWr+fwtIQw/BzreX0qxoeH6+14lZ6eYr/flJIrWF
kY9ujmi5PRYIiENgZzntka9imnm6GgrnWrLSiwB0jxso5sK6p5IlLujqSewzspwj
sP9nSjkpWJylZfdUwNPW6nIA5RS0N+HyvCSx0qtTwgi9SZNCHBHSiegg2bLvLRDh
CntsE3I0LyZCEHRknhr/WSfIZZFCxEdhE73BX6t5GeHqcXDMZPzKVaRW9hLtGt89
XQ2DEkd6sNn7//39Xt1UP2CrzdfWdt2jUNV2rSndcQVJdxDlOrRcn5NzHWO0qbA4
/xtCQMtJxBoDwB8F7XRABimb8vK49PkJmu3GQx5Cwudi5hV0nNXJjrjW8FPc7jLl
rIl4B2QpxXHE22LZxOBrBRUWrW864bVh05aqQVI/RjU7k/OyQ3GuL7AoPGOfmjca
RB0Y19ukVato8oS9+LBi6va8qcqBpHnkXQIweK4EghLyRu3bqU59IpsdSCUKBBw2
QueMNblInBNFY4eBMeaUsJsgOfoXyTZiRSudO0my4ouYyBsByN1xvf/sOQA0Xzlg
E5za7rnOKrkJXxfDjADiNJFO4ILcN6d++47D1V8kcY4kR8gNqb4F6P/HQyAjKP89
zHEqxCHRj7LlfTTzgUQml1RgcPjm8WM01Uk/qdyzYLRwPkMrBPDadm7IjSpWbirF
SfnZ9P0YS4f94OTQQz2inRfiynt7UEb+mNEpQu/qJ7MrZgPLR6MqJdLye47sWKSj
PB7Gehjl+jzSTm5XTF7ggXX6ZpGHD53t9Mkjoq2RG+5288MwvjVTNglrELIf9e2o
MI/bQ1BaVv/XAoggyTP0WS2pPQ6QTvtA1v9rYITQ/dgPd5TIqMLPkN68fuWHD2wB
ytEOyvnhj7jqk/5nODeuDD3TQw0FAwecs3486HOSsTvMjxmejiNI41YbEEQOqoMz
37u3OXCga2CtFtYPH926Kludsf7sp+WxW53Cp6y5I5p/gArAx4uiVABd8OIiIztt
ukObF0MAI0vv5QCb6rxkmAQ1VmawbMPkmhawWj6ID0ABcaVVkFBLxeOb8tR1XxG8
d8SmeJ8o6GIKVD5LZiE2l0XqFOyQ1M7kKW3WklmP7+O28GYyepI5FAESAJ/T7wGs
YbgKEBRCkIbOAkJJU8+b2/lxSVBIzB0VpgJHY3tKINmcmIg8DSudw5wSyBUiqE+z
kb2DUgVw8lYaLcilEfc6QY/p77GNeFeEyvXRDrK4NpX25U1LgPizEP33jCAwbkJi
wMSSJhdC3r3KA0tzbRmlG/SMIhG1IRIpTIKPecM7pevl5HGZH68OZ2W1fmLcye+Y
WEH/vShy63DK7KBBRZTdemyHjQsTcaIQkkf3lBcxKU+QXUpwsYeO1RhtC3yadF4C
qEVCMAFFWahsNfPu/cuXrTe5w+JRLbNOHjfXY93Y4uOm3uZ+KdsFKG9NQy8wFYsf
VHNrR2pcF68pQi6CeMHroFSIW2q7YXbKzxk5PMGRpMfAZI0zi0HuEN59FJb/7JC9
DJtY+VD9JoKYMpFNsUzvN2AAQAF8ytrv00vRM4hKONeXNWPS1ktskbObgIkfKibP
RR7C9FO2s+TEzgQehf0ST0EOzprJ4IPbJ5amZ6NZ1K9Kz9IezZQBvf0cYgJaqvV+
JqDWJ519rsgDZJhMgrXbHYFU0RH55Ii5/GUn3gvE4dw/pqgocx5k7xX2BEX+OqSS
xEvPfemVekIreV0+NzebvoCcEUG13HQd8bHU2wy+u9ZdrmlVjQnjtlmnXl9gWwPE
dlZi7QH+1gVPB2dx5GN01jSsjaB5GAd+TBugleHHBP3TglfJqmHi2PBXiPMhEnzX
hJg1s/eOAw24HUDdDoZASSGyOi/vKdHKcDUZPBpDsWCrUkF/8jnzRsUMuOtF6M49
3q9nDWYFgBqKt2fl9iLX3wjd6DAar6DDSONH44O4JYndj7tPpEtP92qX4JI/inW4
SwdNnrs58MRIf1UmiGx73sl0Y5B3yc74TiHBWoVmytYqCERHgWFCQUDcN3FQ7cDC
zrVYX42jsn3SKahwtderfZtYBwBZa8gTMxN0I08klGSfVJ52dcXcpmp/QaqJiXYh
nGNEueOLSFgKHejD9kXGGEtBINW78ct0cd234Iv04LKj4kAAJHtJYkg7nwPyDc/W
L5R3uUHHzSHUrdFKIoo9B75rpeC9kRqeb5sAtOL53MLg6gPtb4WMwGAgIwTNMvbN
Xoug1/UmmjkAts50nP7pgYS8MjS50m2V3+H5TdClZk8svngfIvoVDFBWaqkmtsZG
lbmMin1FRPwxQ/QLdNcmHjIP/igp1nXxpdBEiz0XkQnSkZor8UVqofbZ0vLznlXS
uhDYvqHHHoCvxhsj/0YTkZIuFBGSe7RfmwN+JrYzdsrt9QDxxq9otiYZzeFEroiv
UcS80bsqdP+l95ty9Tp6hjNFZRGz9ZnREfr3br16aAAe0n+HLqZLjyi9XgcbVtq8
6Fr/S6OmnW0ky1aDbqLupJRDAEfdppCgJoPjCBkYOEySlw3uNF+lzs2/TPNv40ox
WN9MwPUFG/fNPJWI2Fr3s9rLgRtdRet1s6Ix4uD8mReHDfFZms7mpxLvIPRk371G
5UdUNfpPUkhRyiM23RZWuleQu2XlREwbbqFjrG70zJtD5VhXcaSuZ43XVg9aFS/1
JISYvjCh2ePh5+iXvbYq85eUBlaOaCyrA2HY/06RQTp6ZxCzWtc1fI+RI6gqQhdk
+C+bqwvrC16On6v+mOJZ4ei3eMXHbx494SAQXOd+vBApc7K9QknshuV72NGx3p71
hMTq2kS0GpmtQ5IIh74NbAfaa1tm/70zIsLYCsHxzMPYcieW6zQVOdewwFPn8X1K
/pP1fPMEEHfe7oIeaIxs/FBzns13I2PZv2oVA7/fv9m4W4EVUyI/N8SARttyi0TZ
LxCz4xwCN92cRH2bFoyxw+OV6Bu2i8b/mp0qQVuF4tTp3C+D19kbSRMD/J0s6nwk
wHSfPFmFfHFHYOOs/zrCVr/GIxYcwMySHi3wb3RPw3gHoo99HiHOrWHQktGNGdsA
fE50cB35RtVgWlpEJTPIGfttkigmyUz+zk2wXis5+D7xQm+N9vWYAyaVqogHUWjN
aMe5hOWcfRdEIsOLfyEFOapVUt856OfR3FMyU/U0Au2FD6Qy5d+aRgP1R5pSMeoW
S7mcfoPGp3fG238EWxtzIB3vavLmBFZiwrqy/vcGWHFaBQ1+sY0V8a/22lOjCeVe
zumqIAQDtoWZIAQ8JvRIQ+GpMDJr8YC2cU6RUmAVXsWbix6yP+P0FgJwjDtjr0pr
9MpqbMFahuQtRCfy0AVKvFl6JWyBeLC9ajbo6Zf+dD5wpx4YYK2UrxU3GXoI/D8/
dU/ywf+pCXaEufZwKzA7UTX2hanBXYiyyGlSONxUdpDBlgNuh0t+00NBI2eu+wZj
Ucza5G8XcfO+Mu60oXbXTnYTmRO9iLPEUlbIwU8NJPD0QUm/1gmDwM2LeyoA+nV8
wZy5JAJuXtJQpQPXNqh9Uec8X8mOVTIJ8c3AXpbIrcouUGu7+nYYoVIqgRX3x4Bu
lVix3pXgQKVtPX6AECOa+SDSYg1Yoy2okT38bf9GxdD820Ywpa2bwSCRRVQA02uw
0ylwRWuGp+z7gc3EhJ9hJ2hPWwltDcZ2H2oc3NEs35EMxrTkTZcYU3kI3RxAcGzO
JxP3YFhYVEcjim4rxcEu39aGg2RXAhtXcNVAQHlctOWOL8tosnWKmjDnn4ba9BiM
B6rgSBjfoEEypKijcPxt2VSFAHSDN75zoAXAq3g8R0ZIUnuNMwpoCWrU092zmATW
mNlt+aP68JSTGmnPwNdCYNzMtBIXTozVcQ2EWB27u7CIA55zoQyJUikf0ZNwv5FP
G+Lj7KRomTyXo4OikTec5+X/xyf0fQeat/UVSQw0t3IodI+sXB2LpH+MhV6gH/5n
GR1ztyCkqSK0IPAXhe05DTSIExe2nN0W8EMAk+1yol3AGR3gFHcp7iDkdT9Y7TfL
YteLyKZ5RM19rJ8wTEYuxt85w0D4KjXXE2qlGnVTW5zsXPCLxiv5EYp1kQWDH60O
sLRxicCdgG3v2r70qp9gzz/4LjNXWxp70OZIyTm5RNmhkLqciP092m0TErl+h6G6
QF81rOeSLxAC2CpKOsNfKvqr6Jicl8EhK6KIN6KqLtSthoQrQyiCpcHO7IOxARJC
hHhYfViTKaf1vT3Fh+k1eQFAMcyaQObn2k9wmgU18wKmVm13vkLYO7twjUP56rqv
ZzsicYRi8wdl4BoRmiR6v29W0BzP8d3/aSmJwH3sdp87iXzXjn4Ox4aKHzwp7ROQ
fkyAN3I22m0/aytPV2GtRAeN90OWs6p+YIWmdcSvMFTm3qPKwV1IYsjbVqxGFCYl
dlX4ylKsEEjWrMQpkkhGhci40BFbvFCUOvT9mpknPsGLGSobYQOCAPTIs2p+pZwx
xD+Iv7q0FHSUmAZbTyJL80mOeJW3sLseWS0gDqUgXObUkOoFizm1HoNZCd5PZhT/
svyL/SMrn5sZwRCXpduZUS86VWBjlkmEsllAQFaZW7iiYqSIoL7V4516zmlanSdI
kpGDczYdn+IfCAxdFf28uHK2THwJbN3nIeVfjMq+K1gc4kcC2i5ylG+4gAV4uNGD
Gl/QrL+mvs4KFdkaX6oH3+tcXLR6w3FOwGTR/mE0+6+q3QSXgqpkKFi3reoLu4v+
vr27UeeOw+l694isWPmTZoc0JCTmj9Gv0axs3KjPGmfjBUdvRYpQZC9v6P1dfCre
6wposa/zPTEKiT9bWjhF0oU0TVs9zQbuFvUnDILZERAJpy1g7lZIyLY/Lzynf8hZ
LNz5tyZkPx2HJF2EcqPk3jE0PbOG71rroGrNUIpHzzlbY0ZKGfIGOxYcU0jJ5Kdj
G7hGV5+inwYFsXt6MsjLGRFn0rsFexEOUW1OAfId0YAz25rCznGHJ30vx/o5kpfQ
ZqyMX3rE8FTAbh3/f9vrjxIBBMMfS8iQOMiSALPpGf+Hv1jU12T9x1MhE5DEptj+
QmoIxazTDSnO9lczvVeu2baW+owK8LvJbZEi5rlJxC9wQ5+2izsXiS/ZUYmIhDoe
uLx7A/zDb8GGo0KkPpKDxNz0bk+l3BIGD6pXzZsyfJdMDXXLvNrYMHOG0Xxdjb+c
3SzaGwTusOKri1gpZMAkLDiYdp5jKwPM4mxzaepesEqF0PW8A196jK6//ddMy7jk
Fdfg+GikVDfx4l1dKGzXyoWXYN6xotmMfP95bhtKV4HXx8u/Yw+x1R7QylcKlgIT
CYI7sQodaP6x1AW54C1RaVbBATlHLSkfwlPFDMwFizyD3DDrdnyW67L+dbFJV203
BM8zIFuENVMDZSwek04u+noC6pWrj14NKo+DWGaKDSJ8ahD81DmuE5/ZtnKQx/dT
qgVCPXna5+LX+r4lwhXUcZTj1siCGrIYpNFyTkKk7bMiOrJxwg4uVj6Fzh5jCdBu
VcGcEIR65jxNL64HnOYrCAmioXomW5ixyXC8/O82s5zBUklSoS0fs/bSg5aS1lwk
PIl1ezrUZFlFLH3jhyjn3a3dcnswOj3TuiPJ2oXnGmEJWJWr2Lkhg5YKiNjYuxiU
gZJz+d5Hzniwb0l66+DRONlXKpEnETlMU26kG1WrNc25soVSMKOuHtWQDJsBj+oI
mIahGUtXRHQZXFDT2xeEGQlEx1AsixJKIJPcD/J6mmRKRjnblQexnNv8y+CVZX1s
yI0wPEpJqouvYB5toS2JHZVEWU0PyDJaybuHGviMYI4TfmBlHOQPyPu53r17esak
LZaR7fFVJChe7GoqyAEGHtXC0/L2ZqXKdF06thHZ+IcAQog9jEHOpirPrweY/IvM
s58ZvlEuY24YnNt6IhBXiIoTK4cMU4Q4hr1ypp8dxRZ9803xi7toFVfW7GcZiu/H
mb7Bpi2tymuuNK2b0bE7s4Z9onX0ydX5JgQU+CEgCpY4K03K0CcPB6jqR4XJI029
5ywGv9SpVbFmj7ACCxbkyOU8SCfleBc0grF8qD4dqqLZnqZOp7oMvqnTFH+vRH17
u4JK1pmJvV/tfZBePihl5UYtfeI+ezOV6m82gmI0FclBw90KS3nKA7ogFpWANyr9
++rxLQI/RsZnmj4+mcgiwBhBE/tsUHoCqZKtEnuUoamP05IAptVE5XaKVUE400vK
LAuzts+q0eLYIcYPdQwr/kblrxzizAxyqrl2l4DE6cWY3wdqtE84d8tTWuvNH5b5
/a1vkSsWu+kpLHo+yORQGlGO5nxv37/x+Csl6DcpN4NI5+B7YC2PYsiDvYnhIkua
IF68MOpT3+wQejv0X+eDW3lM3D7vpCLGAQ9OtNaYdC0oIxuADnlgtMPwaBrnx4RR
cA2FhJdLB5WchaPsOYr4tY9PhBaq9qMX/LNgYyuMOl6UxoMKtCFysSjsF6m+ymrk
DcL5jO3OHrfF6+9tq3E3df5MH+AtkQzYtrEc2XdmqAudXjpfNOlVb293Efixl3FC
b6iuOZmaGVBqeDduaZcZdrMb1HFC5iKQLhEyXjmehneosStZmWicRSVOkE0Ba06j
+IwUpxF/qMjThHxZovyileeBPg1zjkv+Gf+2rcxHggiSm6N/AAY9Enwb1NSPWPmW
Mar8X86dCOn68djdd3XssW5Y9I5RsIQPqbQHC0Z4PT4795qu/9chZP65JlcAd/fS
p0FYtftor2xfGr6PuiQhgHRUEUKrwZnmgTJkyV9KAReXnmt77JoWAvzxzYAMxpwV
Tq6P89SHq427c7cUVZK77HoEc7++5ynUD9qlAUNWNHxjWy1Rii403lCip5JO4zoV
g+zyEENYqehokNCkeEZO/iT5AIhOPMjH3ZhEi51+kx/4B9nP8dkJ0ytIhg41ImKm
wVQacar0sWCs5PsMDirvPTRbhisU8PLGIt7ejtU3xYQp7CAWPusvYvSFuBNEJ6Ry
40TzQ8Fw1Tz3DyrbOnexgd55rmM+x89lRq+a9NCf6sLYgqiA4sToeskZwm9d8U0h
c5VsMKY54T0T7kUK+dE+9QwbOHk4w8CicGM8HGAsdyeYF8AzgE9DlsTumNh7b0fR
eQw5ysjOhOtg9GuEz2QdzC+2QZGB3bzvuKyJDqxm05vG1EcsfTBr2CVjASFw/GOf
+9sI1Y5S04TNfDQS/2/lhRRsgouMi57dgg3+CRegQvRFX3j6kySSJ6O+ZgmZdxeb
BAPMHgQdQ6LrdPgsWPmKDTJC0ppdRWYr/qiXpVGVcZVobjVJOKQznzgPwzAPOTY3
NJy/VaBnGf9Qy14SzMRemCK3OmTiDzv5S7WcbzcIEBeEwG/3RTnWwWO7Rx6eYPD/
MKLGTLemhq3/JAwVSs0bdYaOZC0oy/bgUuwCduQ9eI0zshV6Kd2JZvBehex8DAAJ
FEHD5LAzQ8tOf3xcgg1pQd4Jgh5FItH2qZ5H8mabhU9lCD6skCw3oY8cbdjArJQq
x2kAI3W91F51BKADayRUUmBtbq97rkXEnckN/6Jj+PrhB757XyaJ68TmmH+w/WD5
Rqi4b6ArEmbkt7n38TzKgwKvoAvRPkfKiGliSxAU5rnX643L0oygNZ+683nBzsEg
YjjQ1+wjDKOafzTEjhZ2x1Fvcwb/QxjnlJML/l6OBxWAnBNDELOqqwSesciA6zpb
ygWFlZmR4idgyqKba9Kr4MeIDFdAYp0QA4BbBX96RlM+peIQeH1p6MEtlw5Wx4Ga
LoN3x7WGDPHt45truX4yltePa7VLTMdC7Kvg4/XFuYURy8ERPHblArDW+zBX1GFt
Hn+LZuNPnKfqEEj4hcPTJrGXKk6ilIMWP6bLhElTNi3O68lVsS5rMxJ6ZDKvgAUa
xCB700yZrlYZhNuiU5CG+20TGOdKOu0bblumRtT63n9WbIc789Pyj+JFR5yzoIOg
WVqn6IISmyFFP9shJWW9GVTWBX6de3aZpfyq2TEDh3rYDhJNEAi8QWCapdksL0rS
WD9VUNy59IJec211hptXIvmlT88jXTy1q6TLT5b5Huz8DPx0XxvXoNpZ/K9iNpcY
O03ud2pnIiFX4LkRpOspIDn/jpvxWM9T5PPB8sPCv15S4Hbmm/+yozf4wH/oJvq0
ukiZT8GMg3PY7FvRnvrBTyyezVNi0odSJ89JUvi59F9vWaY2JKIu8ASg+UBi1IsL
TC3W+idCllwkgag7KS28+PKcaa0PZGbl283DRHrC8KQy0Cy41UlEBarYfQsz6KtI
12GjKL5RmiMePRKqsoprXZ0/JrEbR2VKmh8tuv40tLkCKX/pa7wE36rq5vQK5Cro
DzXMM7o4cVdp34r6cjGXUUhqqR+znxF6pHGFyiczKxe/VvxgNjsMALwQzBEeRHBY
v9cyYpwqzXexrFeej93TG4gdojlL+8n9Spn/5thhafXrLRdv8YEN6p2RhXcy6bCa
bvofpP4tmaC+0ZaWCkJSnjjZTCRNjuAmPepGmiZ4h9m2vprAjqN0o7Uh44FcK/Ei
zJDlz78VoifALljALOW3AxiIGHOoexiMPMkdp9uv+BeVeLkCnv+8h4kBm2YUVLud
mhCrnCdytgWem85+E5B8jdSdTdfMPTRoUKdBkX4qCxJ9eEniMk5aJPs22cRnjJhy
7x9or7Mj5+5d3hdTJmiNEvCEO3pOfY7z8P4MPS9g5oOH6mXQIv9jb+rQurtZybBD
u/ZeDiFKWXfjlwVBqDiJZ00dykZ/fmss/eBxKimepBXKvwWKY6F799P7PdhxdP7i
Ep/OoLFTITHTzGA+NuTE/x0b/z0ISQCvzWvPVgEsriV1zBjmVSaCsNGN4lp+HWKM
PFsJJDMv3KMtP/ujp36yLuc4+PiZMk9e0GaDuMXYYSinn4MBDFKADlPQshmCcmPV
/0Pw/EF3pxNfWd8y26nyh0NdSDR4QXlZABtaNaMBlhUq6Q1m/lN2UzBK1B6xzn9N
s3RqIhcqp4J8z+3mEjHpm2YbXKAeR8Z6nPAWv61cUX/56fU1JBUfKy03sIJGdTe9
901oYM1md9Q81BgA6pmgIxRSKxRajvbxSbjocgvrA4c8V52/ZSpxIJVs1UYTFsrr
SI56VxaGjbggi/paJ4mXpCNUkZ/HrkjI02qvk0up/uasR/DpF5B306thkZRVvHNv
y6C0CoyOOF0xbF3xy8tOBThbbnafLHkaVGmJ0Qyelo3JoiO3utzde/QIPto6y1C8
eGs9LLTM6XUCGzJ9JSlmz1IKde3kMJyBpJJKzwYSB/QAE9FnVhj3MxEAO5T4s4Qd
s4zjjr5Vm+6pScrnE7E7mdZx7EzA4rcC1Ucm/dxz+nJhDxlOOOmxbay57tUi0kXp
o4ZxX8oUc7a4yHhzfvDXyRyuD/hVIQWC0ln/VQ8otFBfEqTvXhnmVyoMbCuTA6di
3iGGeLQN38nSDbXoviMr6pi9s+Gq/4Q5px0JLQpLZxM+kwgL7pI7Znf9+iOEgsUe
CjXqoxrRDs7VV4m0PYyBePtUHA+Z5sgNE5aMRT7omzudirDEttb9HDJwOFEz9VHA
a8sUSXiM1JxnJKWvzwlgocbgfPgGtcNlBYBOFWDdBZOQNFN7VRFz5Wo+vp3pY1ra
psk4dtBZrLHjzWRCVXNEJN78Gaa9SnOebIQnPxD6eBFCZuOuHVjTA1BdgML8WvpP
EyFFYBJ8TMf9z8VLcN6EJYVrm9xgH/EIgi2uHkl5Gv5bsGq98VqcwkUCxoWb19yy
oC4w56WaiVB97kQq9GvXuusEKEsm8yvGehGoLZaX1j58dtwCXfxwvB7I6GUa/b+O
HK53KCTqFrIAqlwt2wCm2pGAf9W9lEOMag1OSqi7TP20js9T61pJIOKxQqyoUQsI
e/vtYnAl5vfnmlb7eBtVZSAJKK2Ugl0jYXrYiTEsgyG4MC6T5RbOyZCWm/vd/gal
dZdRhHO+27N9pTBdxP7whRGvVpC8pygV72byYsactWaBcCQ9Zou1J0r6vnYV0r/3
4i1MleL1pJjEPEYfyFRk4eFGpdyqCNgnwTioFPgwSXqMxql+DHsAR8A6HAgvfE2B
Gt7Y+67GxpbAiVCpuA8QlD3oW+vCrngnBFrylYs/Xm//iPLBmD97FT5ndhJdWbpK
RpT/rXp6rWe72BKNHUckfQ/BLCtrrS6gyqY8rC8uSmGK/1kmbmrMt2Zt/qs4BZ/6
nR5HrzjckUKxaQrEm/G8KP4pfUu98xJEQmJlWd56S4lFE1RW3g9GTDL1ciigPGOt
ybkMZQUZXAI7CkJUAY9g2bbXWQmcTuayI8uTXC973YOD6oHNNHx+MDfz6uFXtdk9
td9C6DtvyATpk7yIf8cR29ebM8HOudD7sdaiM1U9E8l37nubjFMDd7kBSEZ666R6
EWwO+kSsNSHCy8JpOYDAozhQTcwgP+/YqcPQ6bdQi2qwV2wrc98GaiibGogJFGnb
3aO0wALx2QXQp/PBcNljeuF43GmRDWV6+7v+8gW1GnhJ4TlSt96HSq/wXwGnhZ5q
3+kgrYqqjju4XAQu+6dZEjCyHi6FWwFv0eQXRVyD3gz/wVd38ic8xtJX62n46gz4
0azFRJ/mKiLxFt6ebvp/3r3UoOTIO4q/z/OIdtIUaJ0mb3VmvLueKh/k6atX/p33
cTpQAwnK3imCZI/lA+AI/H1MujPDcfNmLH6Mqq/oaW6eAxsc6X6cBmt8H8STsG11
BLjJm/nHQtRHRE5rzlhY/lPzZH5pK1nPK4nnRkddQDXTPU6cR4myIrBVKvfwkYPH
Oqrk8f2z4yMFxRI8ZAHunCHwC44xS0AcewT2Vcl0SfZfxOWFKdcUG1/wkyuXqJCM
u4ChUp8HuNj9+y1eTOZG3Ih0AyydHkZPfhj1l1Fc5d+KHiie6+jjIvz4hG92JQgz
Wm7oFLJwf8kL7apCQLLzw3Dr8IpQ6fkaEZj7VNM3jJXpqSVJYmP92P7tMsyRkE7Z
Dwk7+vUpL0aNJSGmHzf5DDflBpAXhBd0TYaXOJuMRvHpN0alGHszq8Wm5KwuTehc
mtj0SUYKMJ5a6Ylq6D/KUxiLOJeRMD+wCltuj2CSEHKKtKG1E09TOMtUclgTV5fy
qIoZnJYB5qo5qROlsYo2edb/Ba4nzk33iXZsxs71+0HqROiKdAyWKVZpWrb/zGso
L7DhPJITBHOnRrnkUxLWb+M9upQqxFunh3adEG3qjs9TpKniYlJKnq3fL3MynTgl
xn5SkBvOOFDwpZ5li5l9BrVOHv6j8cVgAZmoTXEXKaB2rPHW1mnRWqbowCAqBoSS
UYrWLX8bYEFl11FVhZJOnPsqn7Uq58SPwXAIzdpseByd1q6/AcFnNe/XO7g2Fkzs
yigOt7mV+J5FJotEhIVUeOTLMoO0vFDKuB64+/U4gCUAVaCR6oPuK/RDxkZyfhcq
eG8PbpVHHFn1TWbawGD9Pd1whW6zUHoecPYJjshaZu6M5w4i1F6QbK1dxgZmwtwz
vvSj6jzbTQ5qHCGz23N4Z9R16AeDhrip+1uZYQ5u/bpt5u5iJ6IE7EZRY7kvRmTl
as8RfeOZUYzJ5iWufQxphUhPQqKsJRSxMy/yF6HtbgqlfF1K3alKS8AmbuycHbD8
cauwC+Pv5Mi+r1rJX4qDi921JXMOohTxq9Etb/LyvdU2GnD0DXpDECG29Jl/zWvW
803u+3px/uqap3F7wXUuU7JONs2nrKTJylEkzSp10vKjUI7kve6a6kid0eCQCk4k
XicO+BikKNY3MQdepgqqrM+mVa2OXBJYonPDis7pvEtek8iCYDvEjAnNl0AF5yQZ
QRSpMQzbcFUfYbdTjJ5AQMhqk8IdJKtjI64saPgbsL+KN49cO9EZoN4/E8wqFKeK
df/W5QhTpMfoLEXgm2ZaUMeOOsxS5NtjwJmXhlweY2SYZI1B6jvRrfEljA/d7aDC
acJCa1MIy5G2o1X6ndnx+TTfx9MHaA2zqferItqHg89mWPy/4yOcAQ58nFcJ1P4D
CF/xM4SeAiGyzCyLy1hRqOYoDDIYaEJbNrnpXQi1Oer+U8e1kH7PsNgVZESqN/m0
31OkAqGWs+3zCF96Tj6JGlKXgaV1FffZ6K1R/JUo8Wa4K/vojTJjX4XKdsgWYO8q
kAc0u8+ToZdv42oYnF+ebkXpOTbvtAxyNi0eD8AXwuTE5TXvcQggvoodnut1y1Cw
T19fpGdVlJDCCTChypxizhb0NbbClwSYOAjLsO0un95sKgqjrzwsRN9og3Hj2Neq
tbMC6IGLC3dcQ73sZg1Pglq5bfLvJ6k9ygwbVHeeTv/QHVDdYJnWeT0t/Rkgn8gq
q0HIsHsTbWI8ublFlpB62ERaX1RpLQpwKUSAlAy+C5xAy1HNAboxsAa8d8RUBIvf
Fo0UmKw28qoe8zdUBqx9bTI4KbwFXoPo0MI6LUUEwgbhuDumLwuaNzxUY9FHjtzi
faznm8kdjuS6d9eoGnyXJ0IF6qvQtVZY2lBzGPYVVidDshU5ZuOVpGLffQQIBnCe
oo/Vauw+dK7ZHY1jCh+1syYAmhwUMggnUnEW0AH8wcRNbBFFk4uZtAX7B9YYjaMo
yXlEP7xwE3h702XxaxTp02axXjeYuBLTH/TbdMzkG/uoIJm+3mufNB5gXxq3ItVd
qlwMPZccUqzOFzbGeToFh92TSRRxEj9qyYUowZ1Ndwj5Cs4K/C3VOy5Xhh8Q5pt4
6cUjbUo5OmMBsHpF+7Vrt5/CI3/83h0qPyscLxp4WnV4ldoMSfvJCxg4+ySpzME8
5oEzYg5TNo/urRGUipq6WpDgr5ZWPQr3naJPsD6fsBtnrHquoD99Cz8Un0kVO2SA
McRtxVvRURQTpBhLEXBCj7Q/JLBAnY1NyND20AFytLpnKSDLSuPsJMSCrGmhz0ly
TYi2lmBQilP86XR2KJLxXMTTEZ87O7FlyL+I+tguyOAXDE0zxbcmrzV8g+fQJgp3
1ScPyPEA+Oj2WEcdtG4PxHeYG2/fjnIUBmwgrnhMPwnvkzGe7Ye3APWBaKk5UbTz
g9RmYvad/f7YZkrtGlRdGCcKOJtUB0ph09R9cgkRucdTFV8RibL8qF3sMzjajtrG
Y06LqY/IBAGlvoSOn6zU5MHia8hruTuGXCI4dN6SH24Tg+ZVCJpmNk+x8pHV3eL+
96+SSXMQCjqaMX80b3z1VmOfniFxGBZO5cIrSHdfh4rp0icFNyEkVPMoe4EZoHnL
5fHYiwEavcD46lrZDqx1+WBbjodJT25haENpUlDp3Su5Voi6UPgjmtoHacnID/uq
3Xqw9xCynpumth1DE+7MD0/GkoNPBvsV1Lup9k+Yq2tyIh0SThlGy+xAAPT8azEU
97Klo8a8iIVmi8nr5E1Oq/eqT9jgdMMGCH6NVm9F9vhbNfnoGymhdBRSUvs3tacF
RejD8XVjP/KTkThH9Gar1570sVBwbN4LA9JUWTosXGUAczWwVvOrgsOKScPhzsSD
y7cHNosZsLMmv7KcM9h29QYK4KBupXb8NECPBHlsFnNJcqOyDKdE0lVQisAdm2Gw
yIbg+m/iISGm2sIXT0xJq+SE3dqY9H6a/wCTpfEuO0ufYb9agMTDtZIxM8dBf3kU
t2wfrUl6uLqIRu2b1ZoX53//hu/rdbW2n9UdxVGVhb4vePlaieFekzT4crTz0JIi
qEpxLSJtHSdmStTIxTnJxlVltSX2g8ltAzyh1WHwvJuZGBixU82d+bDU/32Y3+tB
lwSWuZk+t7lZqdhOmx3ntRramnbbzovLoT/TX5GZwiQsPkWDw+733W65wBah6Q34
zANvay3Biidtyj3TNI9eSiZoecjcgrYa6hYM913J6nBLsXGg7q3WyhA+moXsYNiF
lLlU5p8Zcpe2lC69oQGt/IE5+M0Xc7PpUjZWowrUgTyWAC2ulTwtSEnNoFQfghZa
MESlu4sEtq2yrRPLbyQe/DE4Dq+fUti2444czaT9sSZ7ED9ipioLaKFk9YLKXkZk
iu4gz7vye8jb81sE5FDgZb6UDQxG58AdWFEgwl6pjXO382xkdxcou3bpeMFn4Ejt
bdmkHag7Ggf+oXJWbe3ZNQWOnCNNa9m5igImP6GuDBajCpbKunt5satjzpvOnwHm
yGQDtjWGdWDYdgwsYHq6UknjXVIuEqieuSqEtsLGKopAXs0eiiyT00tBRWOnAEVS
Eh9W60SGJemXoLYspOamOiKwSNoe0zmrtaa6qy+6EUMxseKoQgHXfI1N6Nrojwu9
fxxl1HMGssjgZBExgxGaDxHEhjLJfgmu8gr3IUbNJP6vpUK5kI/uB/UZIQnylcBK
eEMs7JqSbCwkmfyFt7a2zBqsp0wj/R8FC+lykFtkaF1ZTTrIfdXu4E2Kmimc72Ni
Sojh+Jx1p5HKl49BTW8HwHrXcLnhxFVWA5IOxYjQWPfbFPKKq4iKd4gnoiH8IxZq
kuM9L+8q2yT9IVQjom5ugCLWk1FCRW4viqOqS04YvXa2ydrig0f0Y/OunN9MvgTW
fk8v6viPSBUv9EQxwYUQ2tnqId6bKG+dI4eoe8N95NK6DJtt2X73VVndjBARcbpe
jkIw4LihHcnxVP5PkjP3ocsloDdaWUfI2j9DrNEq4DHYY/ex7nIFnid05PQAaxnF
J87l62O069ryZUJoXFXFSGJ/6BWastOWV5jFOpQuTK+l7ndn126mfC6brcs6M+pm
qmCnA2jXNIWOewzXfZiqVJRkCfoATXRcuear/x4bPw1fcx+wByTTPDfaepnciHap
P0E0wTOZfJH9nzoNyGOJkm9s7CbBHut5sybkZjK2kuv7cra3ewTV7F1Ix5qIZr9j
+Cx0AOzUTPKdUEqzshJUuyi23qWyBRjjKC9SG9TsWGdCqarn81mEuUGdUncRVKWI
0lhxcg+nxMYd3MYRdxGYPyzRt8f5IKPU2qFjOqwg5/VZ8r67hKLXJfcQ0hoYY33I
Jl95hqdf33XhyOvdrNv1i9wo9UMMA28nkjXaLIFcKQNJ+jFB/Uq72bHu5AXP4ltn
53rFzP89xBNC8aOixo3Ulm5mz9vU+V5QUEUSwTXpvf1JGuAzlOuOe3YQHY7heK8b
JbNQYWydZARILGKYOMGkRKEupUvDrraM8eyRw5rqVkps8v+eiUeIUOQ43usoPp2o
tkluQ9XXrgK79dhDhdBKnbyl8PeEQIMX/DB/THmArxHxMvCQSwmMvnAztVq0Tewm
79MKQZFVZKHRsXw/OFGkpuZvitYWABjE0xSmgY8qLWnMifhx9UYlZWJq+JjolNy0
g1N3PIBLJYyaMnROFmpZ4id2Dkd9frQY+3VSWiKA9a1H8Ng50b4eFEF0x9/dWXCp
62Si4KCQkpMR0ScMoN33yF9qDvVYZt69W/Kt/r2+nF3i8MdUw5/4tO105lS8UNre
9Bzv3QCj0nORW9CdL6Qcf8fyP6VzZPCAX5Qf7OhVq/Q/12eD9E1ufyBcwcqPPvaE
KsWC3+HPcbIAFtOTyO6yqb1YXGEHOj7cUrCq1AhRf4VLyYrTd13OX0G8pu1pZ33l
O/2R7kwRw68W56MmwZk5pfI/tpS6D+fKw14lY6bEGUv6Ja/tkxpO2KoCwb9xE/0+
u5meQjhsl3LA1Y7ZKXdSod74WHsCnu6e5H2nRzQzuWUfuFuFRWQOqU4yHgYwAytq
58Dlnj4kM6p7rY58902GzdSglM1AUZJq0D1mZtve8HKXqRIzGQWroOy+gFt1T7zg
vj9xDiFcOdtqr6OOsVBgIBniFSBva2wfh60qbyB0JA2WapgPwyIGSlYH0nvWbH/E
xgRERn4Djr/0lQa/3xoDlCym7/1nos+Pq5Hbwl2Uu5OeGfPXX64AJozi5WGbljdw
m8CT5jyS+wZu51zp/6MI98QmoaHF5ufkf1POFYGueDkOoVl4ZV8F0l5cEL2bI8+B
83Jr4uJyvYMCrHR6D64u2NiChOWPuq3ZyjRgNP6B8lRFkoegziqM4r67aZxvS7/N
DoXMXfbj/8SnD+2mFfpbbAOu7zo1MmlGFa7C5fMXHMEor4gbJod0Ei/AYobnlNFN
tHbKPrbOyy9o3zIg4ZLRLdpEEclzuJhGyc9VC2L0HM08ZfffQaznhuanbqAKvZvx
Z4RCDM+uG9YXDuCkQnbT5hzE8kthuN12bpwzqeWkU0vjdnXnEqODgU7cdWVQyEs8
4AWn9zkSmZfxDhf+ACJ7y9b5WKiBmVmBG3o8wYpuYb0McWR+fcoTPzlLqaJGg7Td
bKomGhA273fONupguDjxHEhfQBhzscCpyjy/eWsv+wj6NDkcg/PRt5Yp8ksVHDUk
LuhcK3JIduUhM/HgFVs42RrLCQhigpQFBo1nEJ0iZoxM79T6IyoL/x/m+TT7oAxZ
SkLHV9bF+q7bZacwG9LugS3pBnnmUJUNibcOz14TYa/7S2vA27duF15VuQMZGJYd
HJ6LP/GwnZh6CPXvwe+Dm2Kg9aDk20WcwReqUTpwCRibrA0s/aDHJfm3YFYf2IH3
22FCmk0cT4Ud4Bfa4roqPVNiuMG6uYPyWvJRXahYJeNf9EHK4g4CwJRZ4ngB/B2K
tCFWTt4h08OtZJ+JukPf60hiz5gaT3izRp3PCq4gLIW4ldSmV3tAghVTRiwSsQBX
sPIyebpHxXzXeRVzqY5KBwTfUiC3PV/RJ6m/lAhrBx5XHh5/n/K1zK/2lmCEW2Ym
m4R+UIhoR1KYRENWTo55JcmgQP8ue6jHWf5TmOOx+9R3grNvIUvnBEaweelXvj2u
MRHjP4IljtUTXIAq8dZLSw5/iLgokO0xwDcj6V2zcOozorQq2dRVHE7gIdPqWO80
aBaDuZPNMUSM68ybxemCZbiPgdaNUL3/hpFKZXmGcBhVOmn73ePAla1NMD9GMFjA
gMRziHg/Sexf2KMQ9lGQQjOxX3xxWWNzfb0LJUbyQtXrMgVBA9+/CxQavob59+Gy
8nUVca1737WcrQB0tODFDxn8IphR5DP34+7F0Uo+qEin4N+evjoHq/Rkq6gZHRnf
SISRW0q+bjDczaFSVcY9spUlHN006PZ+ycytH3FTNgyaEk3hRS0KelNFrF5hEDaa
1lABGIQ8RE7a65xaMmQ1NCEeABSr1TPZ4o+emA1zoquiCnVO0nxfRAIrp4LL/RTi
5HEQV3XF/xOTGYPPP48RHZKOPXRu7h3XzSi2ehhOkB1YGM/nT0FEUPwTfc1AP2Tu
3gLjU5C36yDV8zqENc23pNngvtbRGLJ1KtkDvE762Vy8vZceMKVGVhqeSi0NkQyf
lrKzxkWaFNvRZZ9lI8TnEnWziqFrMDhZhjICoZasqf93B0GKu1bRTJCdjOaB/tdH
uv74siwIlNHnjPE9tyewMLcF18ayQMNKhwqeMUQwL00ppvMvjHcclt2yLh8UzfLJ
7Djsffj+8IYVjok48qoo9NJBidLOFY05KjRWvnCZiuPW5QHSlIechDdIPpnuBe87
mwngao/XkeL7B4Y3zTBp1B7rBlk0IQUY26lHYmQwvGIeNnL0i4WKKB3IRMq/LSEP
AQrsc7v2xiJhLPvXyqXzQMdD/BVJsZ+fKFuJpmXa3aXkegW4scUYoiuRJREMg/AU
nIy5SIIPw5QgGI5K1jCpgekqgysmjN5vdPqTgRDxEj6c8ESeLQ9K3XOhML396cg2
XLOFMjpyotgT6HfursmSMAIAJX10bmliLkGVSiyZw4nZ5mA7Hbkbcdc2S7cXeUcB
MHmRzKCAi4kkLgeIUQmK+qZvJstJlnDL2DoT3Hd6QUCWi3kWqVbhz3eajo5H7/Qa
DxLQDA0dSgORZowweKwlBu0fJhs1pKI1p8+1ywwTQqVSXJYR3+wiY+AOF/WroHYx
sQYXD8ORVK2NCjec5Xj/HC8YMRq3e+ukpkamuu+nDcZ3zfRtx1QfQUjPHO9Dvv97
F5Pt+3NVnMMa1Ag/YjJYRWOjGuZ+jLvtulg5vajazJZ8Ghq9++wJXyLGPDRyMPu8
KC7C5sBiQkfJn3Mh6MF9ffzJnX8vMQLnIovnBeL8vNGJKNGQZxuSowhE5NHTVOyT
0HgeOoL+Ci7xRNz33OPw7kEfoC/0TxJjZme497YYXX01XdZl9CDNJw2hbZHOtvnO
Xb+XLNTwiiHGrFfVZLagPOsy/foiaQL3AMtQ2IZJ8DkgXivP8/LBCAgHjk1ZdN6y
5wU9mZ2ffqwLtzTzVSsGgdi8ngNTEd2SqoZZdWWspp2Y3flQbGyfND/mk2r2KSb+
kykCiH4SCff1LjktpoQwI2lMntf1Nq1aDauX0t+XZCge8Gemmui5VTcordv90w73
g2jKOTa2AIlgxW+DBaDyulccN9SnA7i8qJ2CWp6hzGAZPTFNBoZqPgIOLMX6luIy
eiIwqxlX5rv3wKONezOLBiDRHb9epBLmZNQascOa3CX9mRr50AB15+qYJT2XtYSW
Gm7Il7qx3soxmnLqkQtI3P1mHVVO9yDiQPmoRyyNZOiMF2F3712DhjYIFYlEqKM6
YeLwIHpzzazeC2V8yt9lA3fZKyw0SmQ66nAuR0LGvg6y2OoIEoIRTawH8a73eADh
+j0rWFnWP1u4PlV1+h/S8BvwSgrNnCe8hCm1kWpdLg3QZlLAk2HRWCm83XGNmO+D
vucZwrHfbI2WbpjsKI8zC0Mr0kXdQnrcMVxH/+Ytne/euhyEsfZC1d/uEhO+AnLW
J5dt4RTH6jNEOqze2P0iKMeqe+w9Nx8te5/f5sKmpUjgImBZejBuaQw7fNGjql8/
Lp1PYdo4lYgBogsWJG6kfc1AEJclL7/+S9XjnO+FwS9oI3/3BchjtlCNQrdhqXR6
ArLIhi/SP/Taec5LvojhPd5BW9N2NrFq1C1eKrG1d2NxqZIJYIK3Cyq4ZlmTDVnE
oZ4arEv8P5sg76d6lotmWBNo/i++bKz0CduDKuebmUxdsRiPl5VWuFG/bP6StvV2
cD31UKZpR3iqo0LfsPsKzetRMtn/oZeaVPNN5jPRAUsFjNfOBMsHGUy/ThTbk3b/
kUwUM9yu6zJvKZWatRdzqDVvSEbHTTSA7b0Nvjrke0vQMq72ab0qm7JfVm5WXYC2
Tl0pG8nEUBFz4QyPz+pCR3DcO1u46cXMb1NR/53vD5RHvHDnvBXJZcScTS5Iw4hk
i/YVeXxb/PMED2p6dPb9P/CWwNI5okR6XtpCXG0AQEKZCVxNtrg7spGboR+StQya
aeziLGu1DStg5nhJgHvUQd+CN3tlzc74bc8cPSSweK4N7Oj8vaHakQTSXcfmfmqS
qpZx0SEuH752C8vGHRGOrvRN7wrTdktJBA4wCGTbHFaR5Kgw6s8NOR2zJH9TySRd
rYD8GGw4cBWjREa2mY8hB8Bx/DBYShtafOKebGQZKFt+E78vXjPuLojT2/fYFmrM
HZx9XbRF4AEoIuRD5YzVW+AgCRyjIiGlizinLN3WZsFUuh7nvQ5HnMmawl4DMi3c
9sIm0veyLSrTFRvS0BFa/mOfc0ZMJJrVCuXvo0OiJaT9mDJbGny0t/fN1e2v3EdC
Q77fweEUHuPY6VKTxVDVnxUF6s9qPnymOV49knKTLk2WsHbykcaDUzPoJuDdZl7a
Q7kqi+PwDkG0nzw7bvCc73QB90ExBUT0gI8Prs9n6lYwDowiIfXy3xzzO3m304O0
9k3rJDUSXhHYp9IVrKng8kC4sfztaDt2AmVh2EJ7gHJBZbZ24s/V+lZNNv1sn9DN
tcplNEot6jM+3OCec5/rZvh7MBBDI1WCUYiTkPWYCe8EbC+rzq3NCd2+CGK5budt
ZxUmgnpDgbsMB/U51KN5A6qR7xmkcbFYA7V6BZEjBd4WLEAJtoMvssSln/S7qcZ0
yvvpG+QbjAoKi5nOuNirFTgd1SirbVhcrgYYlgt2EWt8GLlMGVlQ0m2OJowMB+yn
8BmtsogV5UV27NuM1bEt2t85cJ9csxuV6UPk1AeKooeutPIR1Xpox/9Pe3Mu+3iq
VSRugW1dZ+ZEWl2vWEk5rd/bRhjBzSqnL7+exIgit/qK+kSyUlSsQDOMv1YpXXWt
eWeNXvkp4aKEAz4xQYTECxOvq+GQ668MH4c3fRJYzPMLp9XnnR+VbHMQBJ4voftI
NZDZXNMbY7+/v5kczuoP7AHjzThW3tUkVHMZd1cIfN/ia+D5W9jOnFaa2s7Bs88r
cmtDYtNBQ8W1+CvDVBVJKSiNxOSWzPoYugjIkkDPdA9PInH/riqK5WqxrQkcv7tr
btAQHm2kmlCmQRLdaXTykxKGtiWQocX3TjFRUGqVOv5v1gwh0OglU55SkrYiFrZZ
G1oVnUyfrXU8TDr0815ZHfMub5ISOIJP8p6U5wHYK/zTq1xvtYZxnGFNaaur+qt2
5DAxlq92GYcQQnzLs0Mm1wLVaWObFD6SKoOpWe2YAsphbc1efagsMGBsepXHGF+4
FyFcLIDgdhjGLRjytliUR1sJVbQWrAqm2TtG/fjyD45ik6CHKjypODF2efwZDY01
wezV9+V/GHm/TKE9fIuhejerfe/gBIww5csM5xH5IPXnYTdfrx0WxiIfTr+CIxBh
lR7On3hKWQn+tGpp7U5jpZrKZFl5b5U/I2T2dlC5Mlgqpy5nLR4O3xRAd0Bv4dgu
WIioBNjn8PnbBMrRXVDRST3immKVumnA4/wMTgYNEmpycQLEO7kiL0XP11/78ChA
5U6q3Zr1nrkEMhcz+8Jn75ghSUPF/M4UY8WLQwuKBPdrMx+RvJq8t0AbipO1Agxh
zQXPNCrm9FXiWp6HZ/kNaJHcV6tRW/cI9VNrcTmdwFVATgq5G9mJmHaD74r8kdoR
tiZ9SSJqb8rxcnUzNeva3rYuIk8RX8LaFolkhi+89tji8JboJfVgZ3JeyUhkD0ng
9s9/Ox+PpILb0TK6avwnP6zb+gbf7XHCw81WUvc9r0sVUAt8MX88/+7K6cUoJLrI
KDpXHeLFZS3yxSaJFYJDkYTlAQucGhYM/XSZpApNGReB4AostXQbsWBsLPO7xfJJ
qi/Zyxag+YAOcjizi4PkllU7WfUiIWVusLWIO+h7E3gGPxMlXyeXEbPmKG8Jzxl4
I1QCELWGAsQ8gg9wFsXOI6WeVj9NA9o46ZQADO0Q83SxJUHceOZE1a2VLFhusZrV
byVdR+blMV3OK7WhpVI1+LVZq30Nm4V3zRFwmvkzkzuq7+kN9R3nRcwPZvOuEk9z
j2lB0WPsG3CGRvS26t5OJTy1wagj6rmfd+cIkF4tvjxwSAl1ZaJ4lt4gGpcblZ8q
lF/hvBY73tyxBJMwa6lvOZjeSfuDyceyTO7wCbtEsXs8IhMdCoa4vq7+PF7Yg6tR
956bKpy0LHWq8/kJoboQ7uSheojGQ4IVRL5HkLyXueNHBXcvWOT1ifQ1HyiakFa8
s9JjT5ijMF8QyXeJJTq6BnNUiZ9DCTDjmULiPOTc/mfAy1j9HlSo4nv4Z71sj65O
QXD290fMUj8fGmjRiPFVw/v1E5vSOOEXxUe9ZGG8cvjNIiIB2QZEPqHuQl6qHHjQ
UW6cCAAKPkJ3nYfJHzNl188t25VG0ELVZOEpVNCwcnrwSrd0y9wdbHEVmro1e+LO
3kiYv8PGe1BwWi0J/B4fOCCN1DXl4pyGMfzti3LnU2SXBvEeUQnlE44ls3kBLQ6w
sjbEV9/zBSrMcTOO0f8rO27d+6YyUkjdWPOPe2pOZVLBAYS++6e58vfQb9VCpyv7
QfUxsnooh07Ep6KHDt6J4/D960uRHE/AKRpmAgji+/riq5byw+nOxJSUtjwqRlLH
0MY73pxRCGx5i1JtQ+clxxTGhFMyzyuV2u3/5wSs1iCzudeeC45lMRpfr8BRrMSX
5gdbgwb9C+YjC4fkPB0y3q22zd4vcBND2eFD7GlQGpR61WGWAwxKLM9+HPrFk4bi
W6j2agyy4ZHUrBy3DFTcj5RHalZ9KqCufEYJUOFoxxvU15NyYRrNk1eVRupA647R
YKvMKZX0AMvFPFfPQpY6gHAHeCP8EikV2XGFJoZlfsQ1gAgT9V9Y7tkRgXzClYdV
iD4Pv66Q+A1r4yxloTVtlj36n6U/RDwPhw4EeHibLzMEpSoP9ahjfyZ0ZGFqLTx1
1Z4zoDygH6CftlKRELnAAlm1RZFZXXtfqzQv2fj5yIYO/mY48e+c46b4h4Fq36bl
nqOQ6ARu/RZ/TwufaaaYEHtCilddSt+eP9eRqIiqE628zoxfQbcFOlu/JnEyJ82I
j35qHRbw5FNLw4HfMkpFLRx5OrB2/KJ5cTTsDXqRPVOQ5hM7YrqBsep/cdBn2LgC
3P+ftTgv/gqGnW+pYGnxuXQ9X3FbhkaJwtcgvs8mn0X3A6vQMnG1W0Osp5dSqcVu
buCdg9QNAOS8czQM+qOv9rubq9UwFWs2p6LIBUc6g8zFOpNoyCXDvLMNwBq8uNx+
UUNQqJM+SScmcL5M3H4U4RmCpkQuJj0cpDziO3cN2xEGnQNYj8aq0PlY2qxJinE5
67y5/8ga0UfLR29/j9ZlwaqD1i1KikMl2eEqpzgXSVQFy1Qii0O5VSFz9OAhgTbO
4Z3HD4In2r/BT1uY9d2GSrA96HyPm7U2thzZ4/l05qnVXtbWpn9fwqnNTsHvB3IG
wBwBMEsH9OuV/YyWOI8IP8wBGK8eUFnpBweD5nABQrouAKTMFQSNUcSWnvR0AgD8
8LpwsQTXHjY6uKJAHAa1XLo+a7c9Mu1SbMERdnwjTP7q4HkGBFaLkXJPviJ/Kkk+
87YqLcQi/GYKTNyvmmH8rTrzDiHq1PxcEt44m/PfwDWlX3p5IdUW5sSmQjMj4YDZ
KL3G/4ULAo7Lq/fA9banLWcUqx6xp/0Ljn3RY5cuvzBzmlbHmHtHAqmNPbJgqpfK
5jBDwiEE/Bt243iO8uLz78N/HAwN8peSIQg6RbPw8po/1+SGnMTNjquOvOVqj3kE
GgBChFdcK8MJkUhm4+hjqQ9Qv+5Sp86e34ztDkfeOJ9zInesbtnTtkZgOA55UWOB
gDuPUNiOUjzWVjibeRbgyEnsyFjJHoE7Hg+epoPiHtr0PMtcbhnAA9KpneTEcHC0
+FJWhZWLkB22ZUxXL2qh0zzMUYBLXxP0GiDd//aahYc12hGKb+PxwoqmCTCIHthL
IlM39NBjLBfERJ7ncUX1wJf0TKhibDEQlQ2E4gyw3+f5hV3Rty6CZTa9Ujc6mS6v
ajmsFNPZ/s4cWZ1SybgfXecPmt2U6xx5+x3SgELU6KQ9AZtgjyXfeXf2zvy0xhpV
DSPOuPj+CciuNktV/3gw7TYic/kojrKd/A35fsZMqvbAVgZJj/alhI5CzZD/S6a1
24oE8tq7KcTl2Pp7fZtxXV2kS3GUgRdlO0PHYF9vbAmMJ/U5hc7eIza8xcv3ES3s
TXJCJD5u5kzlu144kHIcYq9vMtzkDRmZW/hU9XGW3VX7pKKF9lI0UkMA0ouH60ud
VMAg0bVn72A7/sT48NtPLbdoblB2oKHsM9jKG0ll0AS2IqhuJy4hyt5W1yKEiwKc
aViXB/efsi5fUw5w6omsE2H3UogF/SDv/16ztawBKcJ+uvXu250laKknjst8Q1Qh
NMv+W5p4G7PIpmujbLvTBSk+Aci0T47214XO6RJB2bmY8Lwv6kA9r2CgGrvcgaNQ
zn0jPsVEQJuskIPpHSHV77FYipGrfEuKyrwd+d/0txVMEB4cEAdESpIpQkF4OJVD
eiZM6aay5Ay1oqNZysmgHeLWR2irhQ23lkLnZuby0lgPFkBvAhcGo9W8QKRtBL5r
faVycqOWdYSG15h+oBdWcJXB2yuvAuqZKc/0iQ1AxkEmByCEXaHJ45PX110OUr2m
ozs4Vyv4T9sadxgJADeLZmqfGrrzwaHXhK8fafR14TNvASPMn6JDgX5CLLlHKx8F
YCZhcNjP6qhVxlygmZVNH2jsb0+CyISnIO1bVW++fSDRda7wpF8n500CSgsOQqcs
0ZxyGeEAQS/KhKxFqM+H8bjQEOSkPA+Vn/lNFVGz1FUDtYd4UDHplTVBbu+UKFUI
hyrZdUepoSlAUvyNsQzOvNw62A0mpOJQsE55bCR9X/NcFdYbHTJvoQBFI5uirPps
B0dOeE3t1lZ9ciKOvHTEVjaQ4BuGTXsyqb2/hIEeYG5PcQmSLCpFFEOHaw4cI+A3
4amV3GoIT+hdhyx8jo0v40Sygu4IW9Di7/hpPyKx2RenoizMUtbzhtb4Ex2wnnCF
R7Hv0byB/NYH7XLIN5Pm05c5Fpp3VLRxxC5eTkELtlpIZRMXSe7wMOygPKk2CUM2
rcJrIrhOrCf5Cpw/jPe94RmxI/n2ysQwsA72ZwlA/u43rdYyHXaou3wN1DHXJWnv
gCGYOgfJH8K14+wshT7nzu1zLf2i56r64eIvMiC2p6g3hW/YsQqPt847kEKlXoKl
tJj1JRGBMT4JaK60scrskR98MVk4sjMxQpAIZ3FBVUtuD5BgEHyONyiGrFPZBNS4
0f3DHWUHzrHao8kKBK/BGxQEkS/Xvh3rUpzj4n9CCdTQBPXrURvUZPXEFRVefs7Z
SjIj105IIYOiE8H6zLnliLcMFGAHrlRZRLzdg2pZTfzfD60T/384CHm56ujWAqqR
8tn+pLuFtnjTE+LX2traMH3RUyjzncO+/HmSJTDFPUUMY7OEeZqs152K3RvQeTa5
Aa/GUXnanqUZZWXC7iuFqrhqhBTvcuepwu4qScMGbCfdIXRaIl7x0HJqK7bBhFbN
Oh5+NElNSglLgwcxhCGDqZHghbmdbaL/JLlifCmNPYU8pPY/f7620jD/20CPJdA+
/ccO22uWbX5B7ZLskecZvGT5EkpJ9vxQifp80+EzWfvVstMDdAIKxKL3C+0lFpo2
5nF5amCZh75iPxALDJweRtJkZA2h7F5qbWat5eMfr5xyVGj4rBKxA86hrweGgG2h
cnwhw3GuWr9+DepF1gB/C+6Izn3bpLAXAzwdYEvhyNQRBW6xF6MpgsmayB5klNPX
GScXtQNzghW7UrBgQ8Fj0APhSraa+dhvz2mfaUtmVEeXKUNhE31WTMhKRb5FGwFK
DnxoiLrHWQ7E5ostrwgO21XyFmLrE/GYDXTl6zrJ52X6UGilrfsdygGCJeZmmjQk
PSDs488870q4ShlRzT7RcjWve2xt7h22K5+BCZvJbsI0GifDuFrdzFI+Os0imUHi
qFb1lixiMNmCHEfKN9qUqd1Mw6vmYbhitHenKGQ2LF07GC8UrC/Wd/ZRp/2ArYZ0
Tz30TXwC2ErrapPTfIQEDhCdFSVfevPXmcrG6fz5e95ip7vfrFLLuNPB29GUL+MW
p4JI+5kv9Rkovhv0R1NiDFUw2WovjpdjZjv3ammKPUK/fH04BuHxh8Y04zDKoZYm
V0ssIKxJRDJD7o1OEUXXGYclARVhvktrWHn5BLzQqE7I2MU+86RsOZ/qGsmT9y6o
lqFeaWncvNYxPGiww3DQW9/mfzSzTUpaSSOHgOR//yXq3KV2oHyYvmisk2f7EG/R
LtgIE7dqIHct4MAuTJobIWT4DsaYUSZoQDnXEeNoyPMs2N/mFEnC1BeRZzv1xnhn
xroV308C+k+RqT/y6+x9QxUCT5R28lU4FV70SwGczv79BN7jmQQTiKeANgiuPVD5
0ss4Ixd5yTGltcmqIvQMZLyq2lKykLUpP8RpzEaxX0mJfCodpMNSPXt/9nJmL0t9
f784Ww/tQ8xPYhk5EvqaExmSgzCq2yB5Ff37eEvUQEYQP0DM1xMf5arYi7Rnq1TI
Ri5er6BQDfYCfIxn6/11bI9ljSp8AAX4LoGyFV+Bmm1F467/f6eS3mnsZ/SbGETX
Kep0tpA/CE/6+siPc/YXrEawuygRYWyuSjZ6BNnbHTEiuyuyohY7QYoExcNg6Qfj
RrSqFnzVDWpydxtUvM2GH9GQzO5l2eJvVKWiKsLxYuD8ECcsOWJ3Uw85xS93uORd
fFimqE1cQ+IxEA2Lxxlhn1twAbvf+mM+Nl38x0bNnpzBFbISE8bb4PFrkn9cbv8L
otlAWgBM2OHPHFKtbwKTKyfC8j0sQgW2/JKEq4Nt7PRRlCIe2b1slTEs2JpllC61
dYWVfWpokUlrLE/CPJ6t9Dx7KOjnirYJVTJc4NQRcuKi3c6vQQAoOAY3CuGmB++X
ZBc8+3kNqrmjyYlB7gWc/x0Cgfyxaqu0upupQM7beU6CA5DM7VkPjkFLnkX9FE3K
Z6RfEPz69FJA2IuPCVVzWOmKo6cbWaua7Ph6XfxUZtMDEksHz5ji7BWPkBAlGcfq
IDrM2LhVp/dwaL46AOR0X0SdKOlMvU9692tOXDBRQHE9XvNEEbCzykckhuvx4rPS
SrqpfCv4RtqaVXa313SkHdU6O7XDbNcswDWgMNyaG2jvxXOwjlW7VipvTaXIZzlu
mB+uiFmwxhfeSydjZ/fnRLC7C0oODPyjCxzcX52MIAD5kWFy0FR3p0PVhNJxhcfz
/vEXScksCiCps1nIaTXPE5gB2/26vfeTnDAh8vwcJng+4SnHu1QbPjDjESEAWmaP
jnwPPPqtqYtI8ZOZtcbjJliXG6ar7rEHydNT/LGgZVkqjq6hXPZL6Z6lfvCGxM5S
KcIHRhisV/9XoQ27jjP9j50/B3/m/rgTbAlXea/tN2YEoMmPCn04UAJauEsEDaev
XRv14O/ASBvi7JtatTU0bqplotymEZvIbjRncigX9BOWrjkhCUUk8pwdhaXVVeYC
8o5YKQ76y2QhuUbGmDtuXDAdjNdZ13PSlbT2rY2/TYAHG32Lcq9L+rebaKZ8Ah+w
pf/d5NWjp/wOIoQXrMdd3M2ILwxwSDpniGjY193VcRLLbNxSp9f64XGayq5Atj3V
8CsCNpMtkXxo6lzytyxtSEZJmu3FCf4GJb5L/SFLfRyguF6kGavvLDSR3h2TcSKP
errLGnN1ei2zOsyxbDVJWMkTh6tULIeSlfBeEb09blnciAO62Phr1vq6aStGY/Gy
JNpN7heHoISj5kezpkmueqqOC5JixhByoPDx1IBTU/YK0TKHoyTQtu9aNmdLU/Z3
3YyI4LqRrD1DyzqZlU1UZKxdKiJ2cAcImu2ooWDG8ccc2EGCAKe1uERoXb7/T1wH
VoXbvsq+RoIC05KQ7Q4O0uSPUJWNoFzkI6OweWquSKn9/YW7vdriVtgbYsnDjVFi
hQA/Dux4kt6HbXoTj1TmFh9bVoniTngvhASFcmFYj9LWw7fClRB72zmwATBsWuR5
x8LYunQYGayxSVUMhDlpK8Y49Xunar2N9JJMBh2gxADTIsuZiNGQoVuQgHp93axV
jX+YuPds1HAQlr9+El3TPEwvT/d6K1OZzdLhq5TDWrAvrulFgMV0b+rgNJR0TIfh
uVmA70my9UYrc+zkusxbBpE0uSDG/pKD3lcs3wBAftN0pa7gALmr+LYnjw9EGFET
WMQjAZoXMuLEgeVMSJeWbXX2ULefvT9XeSnPKQRDIvpNjk4uzKbTDkUl6Ih7SIRo
J/BEvvmALGH6i9i3keuWFwiZzWpOmG0v4yvnzECHqYCfYrh26+POKndej2teSrc+
312Yd5J9909xI0j05VMOlYiV59WvMo+ES3wCw54F5/ZtF6p7FzKnjvKSfXS8hC7+
9+W+MllnXG/UNUM7Noz3CaiNt5puQcy6BfvZvW25+SeG3Ixthrqcjb5DvQhUSWG2
5lTh4ZyD+F5JmcU/FSTukTZcVr37aLg1gZ9K5O8fQab0k9IOwb6sQUFtV3qSIy8x
6hnp8HCdlJ0JdcuDxn4d1BNLmEn6MfUeti1CChOZ2M8HGTAunEdkpXtjzZpWD1zJ
yzofm0ZwcI0bddrdO1NcALdMRIqc+o/nhTTsu3k19+Yo+ki1Ria5NTSmcYoWCUu8
n6Rv7etvgGHWcwOc7PqxiIqm4vDdosrksxG+baFR9srIZU4agpVdoGEyK95VVbXI
4E/PWTQ3BUW0x3o5KQDmbOhamSw3N+xQk86iShVhsLTdZlmqdPoV7aKV3LGsfJNn
/u6R7nKiyU9HsecbaCD5EOb61jpVUSDWS1mbcbyCv+uAys8dNqu4p49HnjIlYQqv
WLJIwdsT7Q4KDPXthfRdMJyzlK14KCO/ya6S8k7QxVFnsTO8Uvu8vD944E70yK99
k8QwBWmpnCSmBvuktqb8RICXOwkLIsGf5Z9UZPW9PU/cX5AWierBHuSOgiUj7gaG
TUzPQZpE3BMTrfjDr5/cibF3GpwxWyL+L89q2yJqXLbQTkFON27AWyCjbZJNIfYN
z0MWeuVAbYtUHCweIcPo0TFHJAk9MOft1eFB5d0dkj9yf4VKsbpLmjmJFHLTRoHS
c7Uzy6IHGeZ0sMOpc2ManiMvPL4KeqWv3AtKKtdznRdPcA3BII6UsPf/3moy3BIU
NmwcqrOsnI27TiEJPCFi0ONazVA7HtajCq/Q58TscSHeCjMYycY8XUcXp9hKkfI1
xokWJfUuv4Yzin37yaw3JJ+/QdSwvFgjQz4SI8+Z11ecUi8kcfd0zjDj4jQ3ZmYB
TiW95gDvgMxM1lkq3EHC1+fe/HZPQiKM1FqOTIk/70m9AUi/9kLYuA6cbgmKsinQ
M9+bY7nG8Og1NEJ9chxIdNF3lRKLbcFQzFsiD72eMHI6Oe8GYp5P+0CgU8JdlNZR
65sW7GtJRSL1X//uw3wf/zbfTC395D5/BhzdDzrXy5lcYF41btIUqKhg8O/cA3pU
RO00urjZoHkxbHoOteaHC1fc9aRHOyC5GZNXlzZ966axXsf+SWVey5vi5EyQZwqN
PJske98wNVorTdA0/R17oMIUAPAj6R81ohpkZpi1kTbDcPDHzqB0vKEeBH8NTxB+
eREm1foGEPNk82j89U+7zAHjMEjuYxpuBdipBJ2H0F7tnymeT/F37gZiBAPKhkl1
97aTv7KS2rvOjD3428jD36BQ0zWF79QXACtRH0WGksYy8oyPfxxqDVYDf0OUMtjL
oytMzdWV2+dDAkCDspVBvTld0EIe7SJs0IiQ5J4YaEUOVHTKslajZp9aK3gSjcTp
TNiZTTxhWayLl1gkxwZFYO+ZUGxdBQ06tCZri7t+vbTKu/YloRt05OZcpG70+yET
TBrGnXFxl0g9RYA+1Wi6fMRDNMd3uzKy5tlOy8zo4e7mXQU0zrgaSrhmwEoD2EFY
tLrzqI7kXUeAKtDHj+1an4qGnhH8eQuih3FiIItEYDbZ8Qeodg0usKWvew0DtQjd
lyVCiNw3tzHJygsRlP5j2giTlI1eBPBr/aMSufD8UWMFNOoUzwUHCXLibgd7ueC+
91YX6UrH3EE8uHGevOeXQoZpNUO/2L1vlbUowITKTghMcG3+lu40JVMHyYnZlDlo
VYDfv4geXxN2FjSVWoLynOeTxBRunkq/bfpR5Sxww0i8shXviXLXY4V2OJcJcGfE
eEEAUamLC+Ps84VXp/XxLNl/fo9rNvQQ+maYYpeKIAUYaFfDFhDNxvpkYkt3+ijY
yb2ePpJCLV/bL+0l6uO4kMKgu35GlXcR9/Qw1MfOj7f+LeHObYaEKjB88T0Np7ZT
2hwwFExaFk8JrgVB8LlGycdf8hVggW2cjmWCT9jgGFGvVMD0h9FCYjj//K6UAOyy
e+Mgwrx4G/IfsatWqOIpEPdwoM+8Utu8+Ba6v95xPa6cY0rrGQVCareyWKKFUlQc
kJ7FozNS4Msf19YKUwdY2asIUViRr1vnYv7dacddWfWOiD1J8Sh/hYCPrZMTKpx8
QuAJw0B1bMPA7U6VHwzbSVABuxvB5kmTcMYUfyec8z+XVp853nVSS27xu5Z5P3Fc
415iAIONwpD0rbupOaHd3GO/tzGcjN/ZNUoYmsihNOtD5ATRVsDdZujU8xGlRBQ7
Bwd52ZNDN8uV+l/n/v7a8ajSMLHpt+kLdAhpyiDpfQZYL26IU5BKcADCRl01YRB+
mByKEKFSxwXdxAuPOyD6qvSYovpvslUWhpFJ+5/OmpYcE14yHOaZaRpi2ZVZ0F3u
JG28GOOg2g9GD7NcDUW3aBjtM3FTxmBYuqm+i/aI6NYE1MkFP9B0DOsFbggw1D2X
Yc1IZ9Q0jCUIJDoLi03qObnXXVPWCo16no+cx+l8ZeomT2AT6BBbDiOSXLD4tfHN
3P4kzZQ4A6ez/8bx7HALrAqpJmAaRIbYCagSBn9qncS7FXRT8o51qZrA7NiVeMr0
jdviYmkgus05QY5GWknBcGFAjruojDNZcHEuGmzHIEWi6uBA80N3NIL9SFDPY54O
Y6Yvb/dgny770PNkDVpwGD6Y9R0nn0GSEHcaJOVAOvIDst9XVJQbjXhr0vOyBrAx
OsIocVjM7eV3vt7oqgdav/zNRRhwW08tgP+LTL03vMmAxRscVYFZf7B+Mv40YM5X
OPEgBghTrhxux7fppsJm9sHb+RTDYmv+VkiMaBRCD2gLnMFr8hl1eBf9+goi49+l
odPEGpKtPw4c2WVGMPW/vxpGX+h7si21xXfj7l4vTprYXovvMrGycNeT9g/ugqy8
PGnBv6Amz/P9BywzU9b8XNEd1if/RtC6xgc5DRPEJKZjO7S3/RLxxJzY2TDcbhGu
+uE43rMnfixmG3o+z+INpp0pDJzMZsu3ol8XhEDKenbs01tHWT8EC6AAOzp39iON
yKwqxXzD23Ie5QVh1iTIdjqmK1xZhFWg446f2YlHBhC5rHw59ieOoAerF/9q4I/V
48HFFA6OLl4qFMq9Mq2/dvtnlo32m5fBZvzKprP3g90KWbp2SWfKpAYMi3wFKxWe
ZYmIUnHFeGzB3tFLOEBbSoxw2zyvYdeWLjRcutmrw/0R2HXUHUFzYKIMnXEvnsBo
hYOgDJfZAHYm1758Iu9dIGVEPxWIdQEqYD8VWtQxIPAeBX3rAvc8JUq2KUJGj+2F
9sfT88ILikyCeKyxR+nn7kF/a0H/55huyZ6sA/mnK/FBjw/V11Z82w4XrM6Ut1Vq
c4e+B4u1Y4/xmzQ1OgKj3aZatzltrht3qRIF/1faCaXP1jFL7VYomAetHmB9zCqz
plG1Gz36D1/LTqD3A8bZdtphf3cQ9NxX/WhyIKRhCAiTyJrbWGSfYeEYN3U1Rdwo
jmfbev3Wk78QM5CfZ7poUOZMh38x+YjNFDXgjMTFBLI0f7ykQCIv3bvu0gM/IPb+
+y62GJuPAUCGjGRsYWkeiJAes8zXaS+IcSoo4qzjK3+PvfJ/DCwcccJNnfmrX97u
IrUpaQKjpi2GwBrsJvnGExVEA0N+ToV1aUIYmjtNXAFA5bbmawdVk02kgKm37zhv
a+FZAjc+CaUeff9xUxUGHiM8HUG1NlKIttOEFFB1hf+ki2LvEaclpXEVnYhAsQqS
z0cY7DzqKcCu2/4hCqPPIJlia4/LHDOr62pDzKbWdkG9Q5PXvBBHmpe/sdi1v5Hd
VA3nrlCPLPqaZFcF3/9MY2OE/+IX+n3uGhTjB6Z6yJM8va37MLOyxw5qeEY3g9HC
kae9L/W7UgttNdcrk1TJRt/+L7Wz5KxPpMdLSUzEGrIZ+YUVqB2BU2GMogepjhK1
rdN8niDPVI5t9mlO8ANtKv1b6HCLdoZkOBDFSC7jvBG8DTuUyJvuntPYhuTx3OMX
/kdyuHGvInNW3I7LMPJxuykFIiWhFJOvkQMs0dnCN9/Kz5iV0TZQ5K6hufBOjAIZ
YGi4lVnK2djA3TqKO/5vawbLAtEhD4iwMSZLq/Muf3WLaaV5EkcEqR9Y1uAAuwzB
+1Xoc63W8wZI7y0r7iqnDukZfzqOgxZ5NTmjthPgaSDIC3jGC9wiBofmRlN5S2bM
wORU3RBP/kgo9y1Rkbcx02qDPotHa1pm35hjn475Oj9lRaXW7ITFPDojumkGgP9e
2AXIYrbOnindPQFBDJYNoxmM7EJzogHBpEGCwgMqB/MaVpB5wpJvR1Max+L8yRyR
NmXovHcbKZOBU1TmBpeO0HMVu00+jLYjdHmmFt7xTrwrcF58DioF/4wg9BnZvKPD
CC6EQj8xMvGaltY0nXDf4h37dj3xhlysX0fRUcSPmIFG4+Daa7OtVGVFIygfEf3B
/n7bJ87rr30KCyU2KmFYTy0A9EQ3MAxpgBomEWom/Cx+UluVQotPf7qdU3CUv1rM
egvxUpzKzkOY64gAS8Y3GpVmMmh8tnctOjhldHsFq/HTDxJU2xIF5lrwFSXVwJ9H
rcraPuELMoajV3fvKo0Avg5mQ7Id9cM86OqiWNAfl701hNzwZnFw0UoHWbszpmhA
XFnqorXUZpWHXGITwvDQxc6WsM+7n6/3GOAmj0ZwNCJrA0UsxO/RdcvYuiq3SGEt
epv6xtpzNGIj9Db5WeTOpUr09xHaJNapjUmZ+tOgnCfzHH7NptzFFsmiPf3eqEw2
VbsMtaNf2bKh5pcAxDLwOVTPL35gfxY5vHfhAEMlKxPjDl8EbBOD/obk8Uhdl6Zz
+hKDUn3debYIMElZHBDjk3edgd6HUJGACE6X1j7mrtP2cNG9otaNXCJS7t4B7Akt
uaPyi74r2LH+bSSGAjPZSfBHifTxn7Lo53DuVQVZjEpUuthhblfYWXl7/PaQROlS
ycWZy+omZkLfKNBXyNyOdhdii7c2FPVi6S03lgSpyiuput3XjeUWAfG3gksHQFoU
xGjeJSNl/tVptzi7zf2+pTlYd/gAC9XKX5t1wrVfQCZGUaGjO1nJiyaHwOu8LjzD
9KzMMH9ylmriBv4BMQ2GOEFbyq34vT0TfUrI9ts3glXZ6FkxNoJbD836CUhU7KdB
4zbnAmowzzPsid2jL2SZGZKoMENHBr3a+O7/5zFrG4LJOfnRUQXaDQ2PN/gzDfrg
C3hZcD8Lyipn60PSZN6g/q0tEJ9bQbI4xppMQ/NbWSn6afx2yZ67vucAHip1j9cP
kx9ETW7+yE6MUe+YpFhMMhkw82gRFONYQ+yFmZBbha9cQbyfg94PVMFiX4L4wIWF
4oTYXmDsH0ghxgu4Ib+ixZWKuw8yJuyidGulDGlj0xLChsyhUoQw8VR6lmegzvqT
DccmnrjgUMjGE5ppHqjIVHhwrnLvQ+yniRUO8ZGeDYC12ugYS/3pDUHUsNn9GTns
FdOm5ceF3qRwjyLGOZ5d57y/aIYniqJIuyOUeOPQ7OFDopJMAfQ1/Hy95q7ec737
uEHAzFfppX3Hmr5XDp4GxKc4l3Z14Kc/RebbGjynTKOOdVn4Oag7C6Pdns2v5GmR
H0yUT/imMPrSWm9oaoMj0jno9glwCRgyJkOlCfBCh/863gP6lkxJIP/htpyliatd
x8qo6Xyi7hXsxVkBEqTnaDlc+Pj/3zdyEd6LIJj/kC6gNNJeBEYKCgWB4gpKCPX8
Ev0B9mIqI0VwFmUUrPfso9KlDclc+ub9hraaM0FC/QhUFV6Z3a1dzJyOc8FZxfQb
ApkoW8bXu7cwclCNDkfJWElQvJHMebyczjPnIkpVeUueFmtqmnpCu+CU1f306Xf7
DglsTajv6rpXrALYNG7j4LU4Wv/OULNTRYdbrAyLovC7LLCctW/obeUqN49TP64N
vYSDbnmyE/Y0GpX3JqPF2tcRFlvozkWqFf1Fg8XINi0gLNkra4KPAIQxm90uur4C
q619HvAqELqzIEqM8t83gmKcZZCQpfrzT5s8BHNUuE8suTTEULbkVXlfAZKgPSAk
be1V1tCuIq+uzNWYn4X1mS8lzneCh0kYJf3AWHXzybCIvRK8S9S1MQQse6XqhOa5
KV7OHwKD8ziJEP2GePlc83hnJX5AW2NpOaPGQ+qXqx3EW5c9vf4IvJCeLOYGramD
eYqT1zaLKpwbsmQYH9PFfXIXCVy0Xbgj4yMaZyt79ZxGuv1SyVXdfv7IneDzAKn7
6LVuC993gri3hJRJFlqMa0gA/C3SqaYuBSQo8BN5pF3QPWozfH/WRU70q7KnO9/L
A80vP1jhlrIjTfOfOox0zhDgijsSMQBJlFz9vxto7pP4chXGnl2Wi+NSDpPn963M
6pu2Eubl0eYqHiHioW4TU11A1sFlZc520tgUwgQ2pSbM0yJ6nAkScJ9/18lF5YwX
NkqPqyc8t+2EcXP2AltmNzlb8/jsQRHf4zXLLhiW0CmVpxCD94uyiOFKGddR6EVb
sPBBMWgpUssUIU0QwFCwfTlS03t2iB0XVdJZYYSnP8lGWec5z9OlqnHr0Goo7hmj
P/sD6DzuCHLncklshhAFh0IsFEA9deIuPeJqOpmrIOORvVk67/8DeCic/SWs+TLw
ILNm602aGkil856VLViatlW7fC9YRnqdFhfuoG9F+Cj56q6na1h+CIaxEYjko/hU
mmECIQFoPp+qv25ZtnSveEo+joxAwGY1AMIczOOi60TfikwOzSJvjBCNgykYREXX
mVPPA0251Um+I6hc1n/njai5C4vr8gkKIOuoijxDWTUq1zWKwFa6zu9Hy8C/rz+5
K22k5LCzQ+YSlltXjqzU6W+87h2WQysN79lsIiS/QfKaxYlw9xryCCAEYQG10Z9P
iISezfsSFowgiRSJ6ino0TXG22JGoZxadglmrG1+MhUOWguKelPQJWKxVHCba1IT
AMwX2nSCmweukP4/Lhna7R9Q08DZjXfnOSewAiv2x9Tss5zEmhXQlHgevesUCKKe
79CV2gNldYH2iUY8ZvXBK/1MW6ufIYfQKgFxzal1ggRYd68SEFKf7yfs7hbz27yV
LedtRcLvBw/lWIvGFtHm/T/8R/CDPFvlRvabc8BpuWaZIT5/teqwUD+M1Sw+Jpm0
5qErDxgdeCyNKRcjT3Qz0vWh/vqTJdQXNrEGKJ6y5g8cyVgue089ndt/OklDuPfP
oVxp6PBnOOL6syJAyc9S2rHwPQjAFOMArNR2fMYqQ0N4iNgCAW3Ofi1JLqdjuLd6
8dMK1iG7nxMcQ4EGuYdQcZBLW9RVuGbWxtxkpJMtcK4Dko0w7xjafVa+RNY+mmOJ
MY0Ywkix2jnvgx2jeegKfa4s3Jq+B/7S9G2zkejyG7cDu1XTHWVaXfN+urTz37Mb
k5wa6D2rU3R0oLwFB+I5XI64IoMX9VO6k1jvg1Y34eIvkzuu5Ifn/GA5gLFr9EER
dfapaJbY3cSebVO6WYsRKA5j0t5Ih4BBtyOxHnbRNbNNKoSg0MosZ0P7P/TMo+dq
/x3Z6VX/THOIXkBYtRlWS1OUcf9xu8nrF0JKemu7yPJBcU/lY3RKrD7jiFD7bx9k
DZGMYuw8rWMmgtojzWP+fJjcTuRtsZ07e64HuYmfcaLcmTlqyPV0ij3szUXZ9SaK
d1WzQjSWVyacaWRpY/TrQiOlrd1h10KAsGLaDqfGP02QJC94W9c/YFL0vheV04MG
I93fFwsHyUDdsg9Q5UmRxvBt0cpFNTPNQa1YRXCE9ZY+YqS2I6DyfWCVbW5XXDRB
snsmDD9e7EXmqEPkDAg8eJ0a/TKffM3nEKvATLlWX0CJoxDOHxKhQc/6yKHhU07F
MjnHoONhVVOH5tFrAkp3fGG67tbTSAzQGQccpar7X7/JAd3T5qOtd7Bnfj/9/KVl
8BHFzIL8zauunV3JwCKTlWvAC87ZWqctsKR2feGg3UWmj2BTgYiFqmLhQ+QVjcDd
HF3JP8lGRwvKU5QhFrli2qwdMRHq8LsfMsdVDBzThGte5EdzgjEGRf7wGeBBFouR
kSbIuS2Ml08RHlczurnKLGRoc2DulFm+xOsTTh35Y9K2DW39WqHammNQaG1gj8Vg
sZ7jr8rgJROg5lIqAEwru6y5itraX4Ap1aPr0DsiLGltBuifWAmtRhxmvQOSnuxm
tFUR36moZ6pHAvmt7KhmT1RQ3HGApLDDST19wXO/j7JR1mWlG7TNKmm3XVpBEmmQ
A+qv5rBETusPO4GiwMDVbDqgAwcF3lOJPBlWthyASC4KFGmB7iLrg6CSSJwnv2wv
lxuB6G8s9Ui059kFfQ0+nFGiWP0/7xAOSNeZUR2C8l/Yy2uuko1g5AD/KpUVC4K+
4wgWVJPWI+CJnE5n5KU5ceeSF5vyOfSgLp6T8NGfzO3r+yvXV5CXjDcikbEYW/Ge
COQt3QPsmJYDl1FR3TynWFGe26TAS63RuPQlvOoz4HaDo3Umd4ZXwwsIfU97oHZv
CmUJNIinPhxIADhvnYCMjPnlrLgTStFB/6PNVL3tIeWkGk4PHp5xrhXkP1/mbcbk
wTHyoKRQxpEzaPqBMgJ5oT2PuLHBBdBH2G6dE9vWvLeoEsqjFWgneP2E4/OiMceP
zOYhtB/OgMWXlykYHvlRG4rCY5Q7cDuxnOFDO8rhIW/8R1+mDhbw/z87aNMPkaXZ
KwwzxpPOLTodp72IyPrwZH/N4Gh3kytlSu1LGqrspLeBy+3m1DwxaZqGK15/AAuV
/VdIXkTlERYD9jbTGkzpupRHDXFSebUYsbgOwOotA54LvhyOGDmW3aNSh4+8WCJF
j7lgdf1/UbgxTj2GBtd9u9a0O3/xJIh53My/D/nAErOAat2s5WBxO0bqnhk3+RdK
TxGCSY+9afPGFyeZWxqSGdTIwTBs4UeI2rqTeXSktVGMKh9CTAecI9b+FV2CnTlj
7zg3eoQVDbZFaKcaj6HqKDyhUqPLiNZQurFf1m03KGEXHjWr1EiyImpGgI4GOvr2
HRu3b0RoytN91GSpJdzZeeWCZz7OKZOxyGxGQRVQt18Rc3WWAuUjC4o4sufDP1gL
P+YQJoillz8P6zRKvUSB4HosXfslWlr3u3C9TA2kAeE3hlHm9a5Bc4yK43MFpLMs
g5I4IqadQ3p1xaeCxpjdRLKpA+i59bnIIfUA7S9UzdWG3ftlr3YTlmtvQP2fvN2o
3KyC5CuVtzmIWOyyEboBb4r5U0cdef8nndmirc6hztVvQGt1poWDimqRnM+nkf+3
DuJjni7IaFoOghlGeih5ACRSEXHruTI7U8P7i1jQ4qWOTotpAX4+bDemo9128PtS
h7aSlLStQi7eLiNFfd9Mwvlsir1JyJZ7xPSNszRadVPLRD8Ac5ndKsdCslrj04bd
3UItHTVGhJKh6LvOSE4ane3cctsex5oO+6cWZ+W0jLNssvS2x5RWtmKAYUC/aSKW
t2jeM9zu7f/JUK0mX8MxN3aquHHafUWOjwHlVw1WgErEqePE58zmaeDHNom54Mii
+1ivxgzm9DsmuPvLOmOoTrG+bX+yQNygrTDVmgWd0LPKeSliUsZrnFTzegno0TOT
XMUTwUuHlAh/3ncH07V9Skv1bszxFGla7jknfFmWBEgRod5tYX25zYlmb8h2DzXm
HzgHjlAGO3jXvV838QshLlBhpta16KMzKGhq3IsmINTnUYAvROyRL4W+45kQ7wAB
vUQP+wGQqMHkSAsrKePi50JdR/XdxN+HQWSbeA/Bxf8vl1ugsDSI5xkQa5Xopylh
fJxuVH2OuBx4Y7nJNuAjmU66Ha92EDF+5+o/K0RU57UhMOmNEUOLgYElsSL6IPLi
6X41A0mw9Xje8ZLISQ/zWbjUAlxtLWCwn0MKFGOqUuKx9/mWr3cBcrSXOdW9Z4v1
qhCFdoOSLp52jQuSAKglOYy7Gr1orjBwgnefQsYfRLW6ouznjoOW+eIa2REelKQy
1SkSAQ0D/RtcziATkSdblq3eqeCFoz2ja5vElJ2OlYyG4n4pM1DqF/zN/3LCx8Kt
yBxajsrhCVMw2u2sphZfQb0VqVFzztwN3e0AVOzzEB7gMDqH+HkiABqaIVGZEaJ/
ZzQs/LSuogdNsmK+YkELUWsr9mLcunL3Dt5tCfNiNtYbPF8KHkuiyNAPZyLv+iDH
1YXFN4sLenaxPTNzuhOd6LEBxOEZA04f/HGcqO1wUoLEhof3OcktmF587W4EQt45
cUcMhDStgA7inrO+fSPjN/rPg0mlETb6kwjjfOs936AUHxeSAMmbfCdmyecqP91p
zngyZfRL6DKGnjAi2/fOvlfD51HbZ5NuTSR3ALV46wiJ2gPMfU9DMFgSv6soJtKt
YEAnw9Xv3T5JVKZuzUuMmzIIFyKhNLxBYZ3LNRlEU5UHH7ZC4vGC3PWIfetEJJn9
dpS0xZhwvBztDhcRr9LaQGaudPDB+NA+aSEKEhwPCd0q+fJEi+dlN5W3SW0Y9FKw
JUOsQqlTvFTdwJSPI7I+fi4i7ZZyy6seibkyoA2lToXjaNWe2Sno9/QLDa7YNTXP
anji1z5i34Ya3V6UJ2BWsMCDdJrOlqUzsCioC8GMIAifzYmcu+b/i7j4RInyvSWR
oivrIyJ0/YKCRM7b3C7NJSeDmRIGeN5OpLvAp4yFZBatmgjiduA+x/W3MNaK8PdY
r0Pdr9+eDAIE5VPVcKe/0KDlS/LkFqCpnRb2BXp75tAUbmwdfs5ajai9+7925WZe
S6qNcx7ZlLVkubC6SqH3gntFfbFWrgp/hsZ/2u3PIuBlgJB8D2xiLI7PLPYARkK5
3qzCha8V1HvNmjUQu3zSy5vEfr2U/sx//UO3lTpUltFiEJNNMfyWl6wtdfufO/Io
t2CHhrOQjWTJChqnsSJUT1j4BJcQUa2rsy7aLYH9A8/6In9UUXPdjYi4EG2x7SVw
q7KT/OF8vGQS1PT81JxnNOmLgpYBvRNo2+9CswFJVfjGVRu4ut+BW9rlq6TaeGn+
aMKpChrKgaVgwMp6+8AselDVNP/G4lATbqZKUzUYSWjiU8cGR1NeI6y0uwL16Szf
+kxWLEEQ/Q3hF9Ih3+anUirUEXBDlDovKZNTaiIVZ6K8Cb9cFkqt0bUdR15nfYLO
wdVH/JjHHxun9RXCkWRLgPvdlkR8sTnwsUfockbuvaKJ5X4C734g0w7aPlXsYuEV
0o8Dhg/ApU/kOck2EEoFtZo50C2HnadQHGQDNWCLB89u+6MOPrIIAm3g/T9ffW/O
vGunxkr1IujIILeehclzBWVlRmGQD7KiiuTsH5Zf+A7QFC2i7Qz7xqEnfG0/p0+L
wOWg5Lfgm8Ix5/Ed/AwJ1HfmLV4i4BTwNJUUw9ZjwpPlx7zNes/9k+z6EXlUWCD+
9udReKbvif+VEaG/5MnpVd4MkBAE3b9xTdUwUNo87RVMziJgzsvr9peMP6x9+aI/
jICn1p57VJs4o6cHC3hLHJUWL/15+F2Hku7XAf2vucc9SltaEofnE/Z9WyCJmxlf
gjIhdg5HMQRWWBuNeh3rFCEdngs2regQKepi1diflMZGUMPS/6xkw8Ojyvxg8k1i
z7avghnWI0pDhqktCA9hM6e71nhFI2gMJCOL26bgw4D14dZqg/WawhzE0CwVmzf9
Zsruvp+q5OoaN0N7scPNOlsSqW8fDs0u9sN4c1r9BF4Xt6uqtlNaLhCihYM3INZZ
ao1/u6s/tedk3dc8WwRnk4QcW9P7K2OejB2yCxNIadOTNujCwAH408TA59sm/Pbp
BNyPdwYNieVxr0EkSpvAMQ6HU5tWtXTrnYxyxO7NMn0tmYbP1S5iSRZ0gUIJtAn7
RwaxlvMkWoVrUbYBy5cBM5/EUTPltGOwnV3W8NCGhBp1Va4wUdttSxo/gh9SlYU1
AW0KWMCEELUs5RVJ/h2Ic0ZGHfMT5sRXWM2lsW5cd0qNzZK4eNYKI3SHn6z1JH+0
YMgnSSp6GjYSYwWIDBi7cLvuU3Xno5lNYP//6sZmHM0I3d8yyLWObhPfNMwgAh6Y
jeJHtjfl7UfcnKAt+6rQFbjbUgFjfDI9jpED7uyM89bNbn0cviGqm3UP1qvHT0nr
FvLBKaVnYLMk703l2EtVC5eQuiotiXAEH/sE1yJnb4u42wP3j6O7Nfm+Zc/ZtvbO
KR8/WTyDsHjQDIyUfIBSUKjq/ntBFKgQeLusWxPT4iabsLozUF1kCyH7ie7yNRrF
7JfBU7xDtc+ZuSSHNUikedQLkThIdX9g21x11IUW5eNt/Z1/02ljUDNMEiK63Uky
7hJxLfOZ0tDK+G1QRWsE5HEKxtear2ekPwY6gHkBvmQCgenmVT5899vR79QhV15t
JDmf9irnQi0xOxsBtCXKfTET4maWgTvSILB6Flkce1ANL/yiK16WtUeffUZ88/gR
4b2qCINA96l5E3/UcWGc1vQvbDYV5Zi8bgHh4iC+R8i553nKt5XlaN9PvpNAoEuE
BSdeMT4MgsZnpZ1isDz9w1PNwhEro7TtE7dGH7s13/FjRiHq4zWRVVxRIi9xj7L0
iK/gAuVUmQ17j7piIJpmnMId84txxQgucKbSVgNm1TiAZDXk7RZ8orGj4+qTfwvc
PT8W493tkidyipCzBgt/r4yOP3D8ZGTLgglSWZpiIdezhf3+ALCitVCl4TG8pyK7
LrzNZWLlGoP69+gLzyXFPXcP7zQrhoCwka1voWsk5V5/hSwFTn8UjDX6e4XzTfzX
aJonLqBtK8bJ4qLt+2CvEKSE6nDvHHjo4TfNloqhfs1lkOJJnPQ+OC5EjO8pROsc
7iYnOyVtBhSBw74AuAFQFc2NtibBbNfO1x02nMBSe0oyDFz8QVDo6z5k418DLhuM
S0Xx0NGUtZnJe+46c+xeV+OAzW6j0qKuoukhqJyzNt2OTgoEBEUza4pF0T3WmwZV
VmydGLi3XuN8mMkAv8KEgt+zytVISCNbzEg7mWxYEII7GYmqDbCX6bhpMoOWkFsi
hPs1aznJ+aR6ciluTB1bNehQSq8hsQWLwe6GUd0VGfKfzUpivYreJ5fIacuS1qyg
bTrNZ5B8f2ZaQvL6nVDPrjua0YwIyWvYnN3QC2uv4kUUw6Dnxgu2+66czGSFHG6P
EOv7nl6VKRj5iZ9ccOi5qWVqkEK9kMb50riPBGq4aWsNMMtNO4vH+5YnatrTW45P
duCYBBU4FWJQJy8Lw3kD1id3Sd6vUUeb8XkH9Y3jBHP7rwANhYmGJRJHMNif5VSw
MaLe3jI6ai5Jje93By8nlLVZvL5QT/vUHzQdPhvfrzbGJlV4imtWO0wxHRSyFUl3
0o0GwZbVZWZDXfYxakBddHnjmKS2JQBij2VkGiX8bQFLlG4ZoHWddP1CgFIMN+DM
XNtFwIKLM2YVVm2msPMWSBA3eY7AEJCTAJ/+tX2z44dH9J96cSMIOk8AzqmVze2Q
O790SU/dSrgqrHtC0m42KZNtVB9m9v935tPXHOhbx6+i9ZMIulFjVuox33D0clPw
sRuUu3nc2llTPGhiTsLLxzs5W+ugHlFoF+1Nh6nNe5nxkR9g/bsJczIVCBGJfC78
0fsuaHhs2B3EJ4gVsfcmJB2qcjgw7ZrHhmuw+/SxIMo2COloc/Gr/mjkBrfRLGXU
pN9eV6hLjHVChhPzXjlLWS32fbM68g/lb/d1WF0DNfITe1MdpSdortT7IS8l4Cmi
RTulC1R6mwl77xKmki8hwJfZUBiMh673ymgQ9ubXwDsrLfJieKFtT8fuVF+pMdcL
gdP8qiOABy6BYRS6acMH8R5+fO2Jya4rx/2bqcdbAsjqzSacsgefsSQtFgyVX1Kn
/m1VRcbdmUoSkWiXeLQ6SsS2g6yu3ghszr+fxNyR27TzKIZhSuWiP2erDfJNy29P
GZDI4nTeMtbZ9NS+ZaByozuZ+CjAihJrgJ9pFU22l38Xhmeyqh3F6QWfo1NeB/RZ
l1w1QbogJ7svt4AEyGu4wtX3AOuDd4VQUScXPC7VI0SYdjIsIgUrWSMTr6uYtGgv
ZkXrsua2KdiRHXWQjFbXnIJAmEGeVAUoclX6i2/jWVXuMFAuovZuvCh4zvD8fl8z
q+FvjNVBKKfzls9P+f0VhOgStElB7vTzCtd/mxJ5QqbGO7rwA6c6xuBjUCUAdlHN
VsRMYkpfn74MKJkEV6Vq+dVxIt20HnbgnoK+qcUaRClv3E0gR+CMtqbk3QsYWsaw
+W2doRPFFDi9DqQ20jiZ9Ed64KI+FCZ97ge2oso4FtFYvx+O7CESl7WoZHRoaT1O
p0AF2K6ZZzQohGNJpAJGSHqw+AKqmrxzFFiXFT7MkLUtlsfF6ux5paQlWzUr8fCd
gG9/svnAE2+aqkjonFanpyLMJcLhHsF3BGUXodmqLbk4CBeFDdB2l14Y4Qv10RGk
804O8v30iz4hLu+yInIMW8pW8pbFb0BmdpgzgSYjsXvec4/M10zGj4VvdTf0GrM6
Okq0JuxqxEWKsw8Tk3TaTI2Yyq0RTnFf7ua7YQxx9Z7UwT+KyvoTMGP5AQ7lxJIT
PN3b6CuMBvz9M/GPE1aDFZQuUqImS231esOb0KVQXj+2hCQtBJGXoxx9TEfAKyA5
vaCp+zPx/yln2VU+WMrBWDQOyoWLK7MZO+JqnV7RPqMx0HXytMB4joHt/J0mFeDa
Y+S/KeL4zCDjFPuWIf7oaOG3miECmTrHaJXCKzY1xp2ooHTdyLhkUtjDpL0Fc+TQ
dPwaqxezFhW4sLZUmFN7VJlpsNSA9ivZbz0twLXblIfNHSa9CgpqC8+v4no/0H57
Cbo/u9BiHaeuk/rFcq1fL5jLvy1GiY0136oPa2Y+C1wd/rjlq/pMP7PKvWRIBdMf
z4dUnk3Dm5HdHiAutRvbAG3y9OGT8EpUoMOBUXrR8m/DL47xllYHcQsB5aW+kg0Y
5L+hv8ISDPdmwNhdK5w+ZWbtI53CEjI9fw3BEn1du6eGmYWbJ+EeSSIfSHsgkev1
B6fsSyrp0KP9HW0DsPCF3vfcBneStqT8OXzlN0WbMdTurxqHSqBzn/RP8kWmIlPQ
ZyhwIsgZ3zvLMRexgtSxukgz9S6GxUwkjyG6woytDWoG9PpgyEJ8ge/nE/cvWDuN
JT8jZ+iLgZ0k3/MysyCOyy/Q+SfoWfcVEq+jQKTqh3kzS1TvzE022HZ0sqmrsXcq
NwC3tZSmHzI6lJbrdS2uD30/PXYrx8DX4PGouLHgIAGhIfajjxv+UwJkbjrjI/j0
jtqLeMWyieGjQMEbxMGWDCbtSKyNiawoVI9YP8d1zq6YnwNt2m6VWRlyznvK/ViZ
XiiVoUyl+p0KXYlvYsk3PHRiwttWNgaPNrQWtOUf9Gj7qXnPiGwHBhieB2b5vllt
GYp+0pr/oUrSYkdGSsTUs1YJSgdoTYGfW0T24gWd+zD4ooXXK8bwns9k1PhUCRXu
TbC4TEy4yF7ETo1BT/p1StNNAe7RjoKKbjOKqe+YX9K/a0jkvCxXMrfPWaEjNBGa
q1rCDlH3yzv1LzKYJTyOEd0MoKWpopyoV5IPcswa2HLwIviu8vlOcyfHXciTt5IC
NeIBL4kqk+hhuL+HfUUE/mZFAUBtj2M+lbi8TEq4cC7imFsr7VghINqoQrYKMxyv
UOfQPFZRVLJHFhjW2sAdEdHGFwIUrR5aiwZhRnhuYwDIkefCEJftfvB2CsGuDJgi
nWZxutLQSfMttDwNrB81lUDlLnOfsRuKY3SEj18EBvjJMiAN9auBGMs0+iDNv3KF
XVYcpQvSGBjQsOgqYF/MvNUlxxlRiAPetABmK0V6zuxMujc4NRF5AFrkIDK4LZ+q
xxlJ/tHZ0iODwtgsvX3O8Nu3cmS/yXs0gT3T7rnDxjaEh4AYVIWJ0yY8uOWi8Li7
ECGnfOP2Hhha2cLZB4inZWcr7mm3qjvWMXX703qXGA0ZbeoINi0AXfmgUSw8+sgC
G/1t3mt6gRRTUNqsl0KI/gmORlSV0SQKwEYkx/W09NTZE+sTRpV7JMUd4kZTZxiW
Enj0faNbrdT0ORD+2skooa5rKYVC1VpEjaiGPmaehnzZu5EQvxDxhH2EQ35KwBWe
kPlk6h2qeOmoZL+C6TtUJYOQ0F83RAhrk3E0PSYQ1QLjE3xkZ1zIZUyWhfOzuMqT
D4noVhSFeCavR/Lozysgjdqn419cp57wbeybHfXFD2+6Ze6Ul6Cek2S2/r1Bkyw4
kuk6E4GsmuHQq4wGX+lHnpByJxtn+ngvdT/DOagvZ0gmR7e6norU31pqEgVc7nXa
4PDJQGtYe0Ft4Rt40Bd9vstOlKH1EK6n/FaroN2FjaFUqQQ/nE0wZVL1Nsdk7hg5
/gwQQijBJKsc/SP+TaJTKr73H8FC2c+0h9pMNeLTUd79HrYRqAZqbkS30xc6/8rf
ZP2UA33nL2yGfOH2nDjxPp87tmNAoSuzkpDPDfv0Qmr6CsR8dkW0+2JuuKut9Jg1
s29H2YGu67rQLU6cmi0NfkJ6Tm5fcEvFPZqhzQQMDgYuJBpUtQJkzLYNTAQW1wKV
iAT67ECiExwXK0YLFrhVCSHOIhDoe1XgqktlVnDV+0WuSfTDt/MbNJ5CsaKbHDfo
raZQZKixFQhaxNDIPACXz+ihDb02JIdqZn1giIfQuSAGVi7OeuCGiAbkkr8puCan
qgAoqGTwbijAq2wIxztIEmRyQ2eB82nlBh+8yPejJYQ5XN7wYG1j8PVUnwaMPCGW
hPcnMSOSvzJdhWXNzeAmkI4QGP1miYaBAOMYhTnGTT2WnNzZJrAjBn2ep5eUkvUt
EncP0kgdZFSod7jAcyiA/DJvK2G+09FzEEM4W8FyQHYWe+Nu/Oeeu72wPQ8QMj4n
km3Q7OZfQw1deYwsJUOvxrNZCgW0+iWRyehvrfOSlwjo1HhUDj8YTAykfwvFmo4V
Rh81EkxRa89a+HnQecu1POoKXrHk1xBJjnXXD51So4UPHfrZMs4xHceynyBNnOF2
RuITxlkt9TjLGq95vRvOzzoeo3S7kdbmNjsYaeY/iW3qI1Kzf19DkC8dTAXeX+/0
9kIIs3Mv0ccOICNw0tI+FP8U6wt7QG4LPRl1ADiyLHAFjg9RNjjcbXJ0KC44hlnL
4zHNJ0Ml+UN7tgVR1InFbYq/1OkIh2eoPt3YZJH/jnF3e2nUmlKldute2e9dsZVX
yeyeH4mhm2y7BJp/MqkGp3CF7KUnxCwsc7UgmpOksoSy/wrqcQTynT2kzc/4wjEi
JFMHytpsLLKhIlrZ9Bd242Gzs7Z+29TmHWcHr2ARCcJZb51apRzyrUYR3aUHh4cg
CaBqCparaJCtv4KkkX6Gdc/ddGHZRow44fxpPaYzXGI30F7Wv1i0grKygdbEQCiW
JaewPb3DTSD5BScWw/60Wp2CyUESjxTTZEW3ZVG3QjagmHdRe6t55J3t5JrOMa/O
QW0Y6376zbxbO0cGnwKWgtiCh9mHn3iCiDuCiunuWM/neFX+xM9Bcv4Qg9ZiEWMX
UDFPXY/ChnQT/E23x4assgYtLb6NHWwbzEq0VN1a4+vUa90YHPdbI9cWMtHZ0YTu
ZL9WI3cHgLnMykHjkzxW8zPHdiLCgFCzN+xZgBPwdWxzTETxbkDnK7sDsf2V4xhc
yRFZwoH0AO1EOkz8Z9+aUjQ+llNCyzag2tcU5CSAy/yT+Db9ECQFwVin20fY6bNE
TiZv1uB0j0U0kW7wIQqldeioBzcXRE4ZREBgV4KVpcRj0xDfY8gr43gZ/fBM+6hy
UY+AFT8H94oY2R80yjA4PwGSluTVb1uJJMY52jTcbhzZ6a6FO85GOKRA54Hg+P9k
Ra0lKDaOAf7EIxz528+w5udLQos88DPpZOfRhXOLEB5KtWE0iKt6zKA4k806CCY1
NXrXQgXb7ubYOSlre4jVVYwbc4llq+1ZDiUeRdfkXBn9UqdGJQojUv6DkNR+5quG
OpTP0JTD7M33kQmX0SKBCuw6N4uFzCB9ZvnTnZwP5xCefFBRyZxONFm692dMicvf
yYPciVAUtGv2Mcit1kod7D6KnUnQktboWjI86UOlyVA9eQgpDmRjAUUBPFyXbzA5
wCyhF9p5lwkvWF3wVBzatJ5ssggSAYDM+uhckVHRV+vYmW+yP8MGLW1fDDdMYDsw
W6NqOz/6mDYc6JxMRk0hcS1MH6qpzKCHvRm7vF2bDbQwIiEfmMv0U4t1iB0icmEo
8wKY9jg2eS2iUwOOELZkmrvVfTSkH7Dzr+Mbbr990bqkGtjajv2aFQ5CyPAWNw0Y
MtmTWJ2AGif6sGGUUXZCnGrubkuCY/YdWOd+8uhgAykZCl+21QafsOYGNa4iL0O1
zhfQQSfLlsEP0Wr4AGLP54EAleB1jkr3MVmGZK6WLLri+HvMDgs4XgkxunFeRXUf
kcF8nHVcpd20B2hysyaoaoi9KvuaC9ItvE4U6gwqhl1KrAZTqey7z+3khpMR0M6w
n+KxEOlCgNsV7VcF7w/hLD27lSbSJFTTggrfYnFci/tHJvlLGn3ODC2n7+Bdm3Xm
LMyFQ2joT6hhtrtyT/2UJyF4UwLgcpsVhU6FcVw0o1/QCcKYkTqKJ9Azk5h94mX9
gt6Jl6VrnogmLLNMASOnJcvD8LHwCGq9xgHyiteZKA3AcsyahdQDDJqG1I69Zgbh
j+bSM+AG3e0nOY4U6ze37MNrhAi+qPARusNcTJEvpFZrHwTG/7F8W8Bva7TKDb8F
OzhiwklUnRX/qHjyJDlrxf+bdOjG0TMCYibw1sOUPxW166RpWO2MErmoqYO/fO12
Ox5o/kNZ1xw0jYAto7wU5Y/L7i7epHtb4fwr/tzznp3XcO8UpZfbGTrAzrPgRxEi
xmzajhwI2rlH/dzuSCuXFkUyRcjXaW5UglCB+SfKSRrq6amKotj99wa1mvPj9RwZ
14MlwUsvqMlNc+7YZ9gvpAL6T+B5a+KLzJfVslwZhed47dMWebXuXvSrsKeJz18t
ohxDZAafti9z4jC4rm8U3Jfi6jln3wBo9RQiDLYcWqJOCxLhB1uYmeeJfoSTm9r9
46cP3vJqhbQg+vmY9UZFirNpqm8AV50bZaB5NFV/gE8ZLJqOOEUeAhp+0tTdgAyz
mZ66rfCYsJVrtapZCBMRZ0ahQlgszhRqIpM0tL0o8+1biSp2LtOMrPPPk2/rnn/3
tRGKwCWnqabJe7U02Nw7D6IR22no9If2sEvdDM4cAkPinr7yR8Vl+CSUTO7Ym3aZ
nBsUUyC/VlOeJEaUX95QpYyNcnxnrdebwUstEwjnaA52VB/5KlHVgbr6gxlMasbR
+hGjPmgyrq3X1UPwdOJynis0TkEywTgvKla7wGn7QhWma96e4uWa2Dk5AXQpZmcY
NfbIE7J9SY2wupvpzlmI6E1X1yBkH+2C/o83/AFEeCUCC8JbX1VC8POpiUC9sQZu
xP7Z1jf1Y7JAHMOvpM8if+i4a+hTnxIqwwPezdU5LiXvqYNN5uXCUyBCWyOZE2Do
3aASumQLt6S8OWYLqLJaRNX/AvdatEl1YaqPUXi8dfVUtGDWOdWE0hrFk+zFGfnE
lucr/fq5s3uEQgSAh9oE/mFjh8KW3jeQwpqXQoq43DgmPrspDsT/OBbjDLjzwoU9
Fvvq0IuZ2iY7ikvIDgfN1icikaMmw7P3cgMIy3Yw2ex14TRzrDLclKxTFU+C6vmY
JqMzY4aYt11TI4aY+FdyFRbWq+ffXtqhITrJSe/yQ1zDSJlm+8EpixtjaVCRvZk2
rCUCoXVwj+cH4Zrv9p06CquNCqgBE7N7+5xs393jVfCZINv0x2yE70rnfd5yU29M
7hYvbqgKe7ln9UP3zSygr/rpbSdx8q+ySWwPBrfFoh6FMlDTk30logUxGFyRGKk3
Ht0p8oIsrKYb96ZTjHNeqH9DluaCWAqhTK0VKbVjUycFPZGeJQDrc5JbKuYvVQ5u
/clLL3/0F3MD/QlBihTuB4aRNejaW08EivNR5XxAKFYmHeNQb10M+MoavhMyOtBe
mC4rfD+oS+9MTBHOrdMS0aPfLieTQErpfct9QRtyx875jClPYz+/pj6ZX+jXniNB
mOEJjH6p8FWUjIKu6DFcR/J9EHQiHD/arBhvsDhW/+fQldsyNnzsZpbZEIGm04hw
czACkr/6PGXdAJ+fC9p9otAuQ8+0zOHhYTfAVT0Qq8qTie6KiLPw4nl3NzzXWNbZ
Od8/hp4FK8nD+jTHxdnqUo5/gtXmEQ7PWt4mey99NWFS7B4lJcDsFzrgluOL2Q3F
Xu+6Vdf1qEOn1nzcB+5+n7+PURkbHwlRCzZi8t22pOSdheeP0NkkHQx6EkPzk0Fl
k9icSzZt9BjODeL051AMeCHgYmj5TLW7mv/d1WAklAgC/6wqp8ujGqnC3FdeCguC
ILGO2at2Y66drixQA8ZG+Yibi+gX7r3KTWhQmskt08qELQ0G6Heb9Unn5ujAHRAu
fVEqGqES/vrASzVkfaN4vPFEd4aH/ktn+yx96g6bzOrzxoQsRWF7C83nLsWPxJIm
BnwDljXtA4JfLmI+HjIiUPQJVmB79Gcu7pfxwm2F2e43q5E+TmOnOnuG1Lyg6B3E
6DKeOp6pJiS4QAgW89HM6mZRkf//Ng2V+ifskWpCvkJ3JZhVei+DCLpYavvCSOnA
gznIuY4lETT3tgmu7BGLFFe+fTzWCU0kwAi5efvqaGvG57YW+1YPwSz8mhdRkAO9
sfroIB24emCK0P/wB9k/1AjHskzoPfmIEOm3D+somuWQKPPjG98qzQff48GtCYPM
1nOqK6mK3/thDhFth6xQWwHFbm8wSQWj6jmUAKQLIOsS5x1ccKJICW9dsah4DZS0
Z1iRYpOihzct6BHYt3Uv7YALneUoia+7/bQZwZeSAbz8I6pzOSFyNjYASBJ/IMpd
xXvEvoL69Z9Sm6jaV5ojNjxC7zOjOu+j5ujnU5FyiIERKU7HVedLg8j0MeBTFhk0
O0cJHFXW7FWo+jBWEiDtKFmgEhwdUijzRWJmZhddNEEiu74aFSaoiDh2PK7B6CTC
kX5uTfecJCS9i7V+MDseIPEzMYVtGrxr2XUFHNHO86fWH2kdo6IbmiUu5JGNUPx6
3CWDNRmKEeMN5SWW37OViYxDLGnOKkvc7TG2y31AfE2bRajRJmxLZHrSkMUxN9Fe
GtdCMVt2U+PCvsy/vJGB5fO3R57p7JFrUX2TzMIYGu1di0IfF8z7CQqmnFgUzyG8
VbawcDIJmqkKkC4UKhmNDnsYn7zYLRUCkXwLgeT4vqTwilnScqjXXytoxyoHNJ6v
qoBNAJozTdcvQtap+ot3KNTVijv8u3UtNLS/GBjbjzebVF3Q9ISsTV/NURLkc3pM
XpEEbov6S7mpHf8Z+q6YuRpydXt6Avnlr0dmtE/FG97HLJGji9fk6KpEPVP18gfT
+HFlUeKwkC+y52vr5/6lKQwDK8NxU30jRp+6RlHHgmtWkkt/rGRx6MTEisCKaMyy
1PS64/j0I6XuKjsBLAqf7NIgkwyLB1EX3UcwHQoRbd+gvviMo2zaChOxvphysBXF
RDWMYLSoMG1tgJRo8vZY5cnER45NsStYKk2b8LPaIY55g/og0XPN8SK/uZ+1yrKB
IHBOpRlDMxGAF8sv461R99DqmzoP/gbMXrV04/t7Um7E147EAspdfY3opBb9XTgz
l85TsCfvc6TJxpcwTimAdjNRkYK3xHnO2eeQV422jWbG9zgQrzKJAsdOsO56S0hz
68VaoAqhVqxMZfPOLWqOSkOZYBsyVjvpIDaSxcIRKdbkgkxhXDxrTPsozUY6kyu7
tmyAKVXvHnUF4znQNtJ4mA01APA/FYJs462Y+th+18vuq3WifjpWSf/nnBNCGUn/
0zOXv8HDYe3F3dNel1QRNT5WhnE+l4GGjQjwLtbqnBAdxFoFPKx7fSffyEWXBrfk
DqJ34LQlDvTXlVwcbPPYji+E+RM2s5xBMQvP9xqMP5vN3jZYmWGfrLvCwdVrm4IJ
3dYA9l3A3GR4g7DSc5ekCsk85y/YqY/E3HmIOiAbxOB94M4GH6pffQwgN4F2C/bj
t5n5Pom32kHb8EpR8pvtKKghSQcaeLho5UOihVeJaEo8lll1qP8Gf7n+WlxBzcyh
lJIqkEAzy+MBwA7L0b8h4yrgp4s9bW5/Ilp9aSpzB6SOrrKXyx+a0MItcKIJP2sn
OcvdkQ9eJWXWLPuJWOAfDJbYR0+jFm+BuOqyc13K3pEDh6qjnBqJ3Jo/xnCbX1pN
7EaGxU27WByE+5M73uFs5Mq0kOzzGhyv/Tu51QzmJIZTA4G9cCEX9Txvmfovk0iN
LtmHrZaQJ9J6CnfiEUnMhCXoPjH9XThhSWoGmLpmj3JxhbsnU1kPB+BMTccLX5Du
V3m0e2HoRtCs2LHXaIRsVq2ox4TRpLNuCNiyTCxNSqMfW08R3hr3gUIKLV/cjznt
6J8C0wzCEvHB8IRrfoYxDtilE5XRUrpCvqSd4fRhpB0g5fNjPjRaMcUboKsfxh4y
9ypCs8U8kgc60FjfI93u2sC6Jy3GW92sZVnoRK4QRZLSxX8C4Puv142ta+vI3jM+
ko9RrgAmSMuEfmrux8JjYJCA9zAwgUu0gVZNgkJgWkSBhHF/YGTbmehoxk5lC6vJ
O3VwGVEdoda61bjdXRkGPIkBVhCSQg40u8VUSYG7iXXTO8MocCP8RFh4XhjAvijB
oLGAceu0x/GHXLjZCsZvZLXoGjJdo/6zjjbh0Y1YtUWwRDecg+v2A1GG2u8NZs5p
TIH4g23bKQc7ehB80q/+qqiqRgS9EyQemHS1Zfc8d92qo67WHlz2oedX+9jl66xN
a2CB/gZS6RexHENHNfcg+2Yc11gnnk6deJ9tM9RHctCrMGMAiTDI234pBF+I2D1Z
Zju8zUrg8O/8szCDYHgiRHTyNE7s4mdgWYAViNSUcoXgtm4eiUR8tTKpYucJTp+x
0GON5IFdRK6zfObUXWRautm5MnTaJJG8bCJTlAA29lTDrOV143Wp44XLfep4Tz1M
8jRrQDeGaTCiyrFmdwWnBjg5GrubwL3yQ3VB9Lc9dgStrv/yLGE3twJua6lGL/g1
MLKx9nNiaD2c3VKXE4pXOp0s50zJpvFEsqSOolTuwMnqu9y5GWT8EmrBvmjkhu/B
a1jaRUy3LlPjoNr/NwPMd/8UlD8YKBktWDEApLeij7XfvUiCwIYOt1/6+Cc6pA0Z
W7UpXUbjkT7VJAsrFnzSsObMDAG55KNEJvOoluvNmmdbkgNJo/SgdZMqWz64czbE
3fL3XcHWf4nxu27ReTaHZHiN1cveyMw6IaUXgrRh7ubvpaIFutv+bugZLwhBy3ua
5MK+iZKXnrsYd2U+lgCU5nOaS7GZFUwOE+tCgczK81gU4y23fZkmtV4HzYqW2peR
vz5jfAIPXjgjjuR0yt6geMTzqT3fMkFBu1J7zPkWSXoHZur5MHL60xxEYwxYyEtD
6R+BAa+JOa8jr4+fD9Tx+tE8+oImn60LLHK62aZtQwEW66lCa/ZqUww5yTyjr/s+
sD7EKkNqKkymR78h/g4xEkCzN+WKR1yalQGhZ2kbWUrnOATf1IqafQ6MKTeUm4Bz
fAyYsCz0OLUI8O+Rv0Oub9s+n+ShqpBwbVx99oaKffb/3/cO2QYeX7oPQ1YOBJ7i
YwbKWjKw9a2tkzJIE8Ak06++PyPw+NvpWn57m7mHAAxkkeUuDSfLMSf43eFDXw/J
Z+bpWDzSYasjOJQrjrBxEw1dp1Lxe5YneubAwBUDrXCV5IW2zPJdUxJdqWW/G7ok
mJGkdp2cv36T6jZGdlQU1rAONbiD7w01RB+bUcwj9YpqaqKOUPwZEyhznAzVRX3O
R2HekJtY5dBk6p9+n+Swy4p1oTQBLOGeE3kf9qUkKZURVPg65hc5mxk5+qdNQwU0
TMe8nfB5fTzHtBg08q9AWOShHrKI7y5HOYs2HPJ4W0+BIt+4Wcxdavn7WckDOrcv
mHbYh1ZFDg3M32igguAMMifzbkaH+esml1O+OxaSQ2g1/f4dvrjEaoyxiJ1fPySe
kwYSVccfXfrpo8hSbs3PPnsvimF+87xO2BuF7ssvXuPqO9mDxoC0Twxop8xyBsUS
TKLQFrugpZM0mk1ObYiPqVMnOwhLyXp8VX1viOX2e0lSnvdVuielO/r6CnPipVVL
z0q+LY3/iYVZdQt2j9/PKOegqugV529bwec8iGxKCgPgN8fUR3eop4YajtpX0a2F
DIx4YWGr/iZKDqUCAtf31gpSED+WV0UJSdn/lZC+JBCPDD1yzGu27gzw2gPfTqae
k7DnDrq/MxxuHuFLAAuyj5Zg2+noxUg9wVUzFw4OrHpJvkUg4ot3H4h3bpeoYmbk
oTtlN5dSMWyRXXq8CgtCR3nC2ISAu9FKNuhBeJ/DNQJHSwwjlUXeeBFYUd/HmaUU
0Hl9UkzCyzBudZ9S/RN7TawIUrmCuxZDNu4wxPibAVGUazuD1zUzn2U6SCq2JcAM
nul0NUzX8qe2LbaNqhAdY/u/SDwpNVRSbBxC8hpIh95e+0ClIZBtJ55iwIvFFIAh
INQZG5dMUjxcS6zS+5wjZfYb+2+bDN/4oau2Xx3JoMGHoNPJK6GfFLUi1Dul+y2j
VPWGsK8bI4LgrjoYV3HHNImiCWnerIYqCqrfHYe0bWKaYxEwjY82NFibazx1fM9e
oLxWxrnDAu5aCOr8nKw9af4uS2XeBP5h/qJKSVR8bhBvcWX1jAx8af4Dzo+M9uWG
wp6HCnQvj5kTmwYKS+t7ksFEqZWetrC3HQEaBub8X0cgubOOXdRQ8POHAWEHCjXs
V6CABj8IdXuHMKS5zpoCTncv96yEl6+2eTLQHXtyMuIwnBM8DWF/5Nyjsp6f6AA9
f4QzrSIvXyjBIkFKvEDOM3yeq06rQn0jWcgcOEYUUfSUdKsDr5tVLPay6Ns2Clqp
dY1C0rF2fOmjBmKH4Dq9d0pR1WpcY+pvWAJLF6qrUHEPmsG8mFLzvGw9WsbmwZND
3i2clKaImnj5O5Tzuft2hqo5G7fR+eZwPlHBtWonP0B6UDu8B4murvAC1eoYfnnE
+DmT+Ki3iwuZdLmL3pV8S+/DQa/6Hi5FGyQhbt9d0UruOHKAaP8MeXsEMDePhjPT
kbUIsI4oxVMtkCg7gRLtbt8gi47TIHWnCXeiRuJN0IMF8r/e78pdfNgwLuz0g4z7
GmKI42QyOGkmSkikzNQh+vJkq/w/ussADDNWz2ATmuZRDiR4sPcpoYiJgbHa97Q0
cR11s4EaVkNXrSsdiZ5a+aIsQYIBiSzp7J+ljV6jMUKDPv02FNYRbl10+joEjYzh
t8/JjfM1Q1CTBDp9Hh4tJ3nvN9ltl2XUjuvajEZXpekoZhHLlpHqGhQ9LpgtGoEv
5f7mT8r5zq+zJtZRozfVSVmOceEwBLpLbj7XAGnd3hcXXG0HNsU36n6nl7dQISum
5fVgbkvhQpXJb6BpzqUA1VC9W40WEZG44irN8FPT97YNR1rgTjNcrMviX5YGxGxa
WpV9iuiXVDBDEIgjiDJzWSe/mznyPqJ+GcL6ira+Z+3gW2LtI4WZNcfzRI9zWNLa
1a4B9bE1iDWQ1KPKgfHf9GwJHk+6genFkplG6hd4IvA55XyqQZsKOzxxPU10he4o
VI0HYzHuD+i19nXhuz0LSHv6XrOtLaa4AtantwsKod40cra6UTNVzqffbVQd1vrF
Q8fCZFfGatNdrYGNOPZ6/12GhoOVhMEuDR1mqBSg9efh97Zk+yNVm12kQorozzMS
/bsBRUNDLLTvPrUa24ozSNcmov3GKFxO9oGHhd9o21WT4g+RdUChKwrSE/Ztiy1y
Y/hPLkSQCnXa/qGfazOz7T8MRCbDR5pxyFfWXyhYd8OwOEmuFYQT+tNivlK1j+WZ
pSgdfKiNEZ6HRc3Tso6UmmUyHlNBtphw5YhXRPBnfPhQ6WW8M55znOPNw1VsWSs+
tCDR9NSrh9GHfNkeiWT6VjxrgZS9ofgoKCflPLU1l89ikfOLiwoNYnGVCTWwYthk
H3O7A2biIP17gzjEJdgjMFhwAfDWozqoYFAxNC4lN6d8CLXSZ6Hh8MIRCaJ23Awj
qXq9mCtlDLuzfxwRVvk0qpAMJYOtuqgrMy5TfGsFfMSJxslcohN2lRdVCekQaJWu
pgq/l9MwzcfLtf7RTJVx+/Ou7u243XhYojcR4e640RHsp3q9Lv4dplau9cZOkXYw
e6ur9tuua8uUFmJX1DzkbhUubjRMxPNtZPPAevPandYRtgBJKiEuEvuumfliDAko
e1GAbPav0gBCx6bY88PpCheaaMNMPXdnoV8G7V+j9KyGYSucM50sUu77wqoLSeoQ
Snqod79QHXlZtBUOhmxGsQbV0wFHVPZPQxnMni8XHBPAAw8aBA6F/E6YD2jY9ecT
ED27JyAo+H2o/6yXell9exkb22xGpuYVjJklHiuRinh69ORlyUnI1YxPSbag3Wkz
Ia+YRqAilcgJliF0foYiEkz68OtE0Sh0U0VSAJFf3oq6ZWoUsXUwZ3VbM23oNcZ6
7O3JcLXETeCfjY5/RDZOP7q/vLicKtk44dWiE+8VPLsmmYElDfv6eFoEv4lOBui4
yusVplunp6nhDNJuZVRUwZPpHSGne2f1a+OCwfD/1Y/zaqsCWM5XDgb6ZsbpkjFO
hjF8XqUmEtrm4HATSIqeo5uk0brpK4Ht7BKuB65wph5DecWmiRjwUoPQpolYxxD7
rKf/9hHL52E7UWIcw/HapfjkgKUXvRUVjRYyyWLSApVvmi4edGqoDMmz+YYV7R21
1BQes5iIc4gA94GHqMP4h77LU/WiC6qws6LX/aMdKEO9Jc4//J4gs2HAnzpmYXUb
voLeCEPDE7GYATiXq7/KP/r2jNN4q8JtQZm0gHN010ii7TThrEp5k8ef48HJDREU
+7Jo8DjE5PR3RzByBG3oy54Qgjpcx2ovsX7gmzV6FEYFP6QcQFFkB8Vw7J2wusmO
kPLDBE9amA4hka06dCUGhad81wFc3iZx4ODiwQETdzW0GtaDTxsBKvof1qPFZCNH
aXg0uhKvtXxHxIPUm1SnT80dti+fNHwvpRKcw4YqOs1q5iLMiQIg+avbhtKtsnzT
PizszbbDiv0UpvGoexR2IwRFWZ6Njb9fF8znt42nG++AebbUfAl5m+Kw2seszLZi
IF+oW2h6rfpw7g1b4ccoiiPhD02gIMnkt2OFcm438WkEBgIHjobwHHNOOz/dy9nX
v+tY31eMaAvhsgLmsT0aEBK4i/sYL0Rn06Vp9XO7L054w7T5+Sw5YpRMiqM/iYLP
2Eh5OR19LNmM+uUq3fDNxCqP/djSlKd+kpBP/+vNcPzLd/fkgc4gwOYPRs7bjg4z
7bTIOg+adOtdNu4e/ppXKHAbFXMUtWaK/JppCfsUAhFbSlGN7W9VmCPATwmG7q6I
Y86mdHljeBOQj0Hr45IUfXe/9qg1hP7Oicr7F6y6g2mDVTOT4WYpP66pFtLPaLXT
9IzYBw8NhCwD28cU3ThZn7tZIZ9WQ8YzJvpjQLe9rZfmcPzxEjCIyvFHxNndxKFs
YRkeHuJRheuqxwaFBwtizQ4HDeG1g33o8ycCO71nqVVC7cARi7bhLs8+ka8lb9of
GYucwCAtDvC7i2QU3oVdH8XHoXuN3/uDrOmmUkgmnuZ6GGFSkVXroPaPMtL31fdH
KBVhSVFPnc5KzsuUlAaHNoy7sMd0h8VTwgnOC5TAEvNp3aZ32KFaK9ff038k6rCz
6QUZUV0EC/ILw67Kn7fve40eDYsVsTWo2JqJarcn/Rb7Sxz+nr0dvpF6Cc2KkZ+F
izNnuZV/NaxF9yk8OGeFQWTvEgXhKCPrq0zzJF7QZ/WWHdxLS7JQbb7EXSPS8v+G
q7GMntGl9ga7qYDjdgYYb5BsAoVlFoWdHae8YcmrzEzplwNPqnW2IJ6lnUVfHzMy
PNl7A8+vN2R4EJtVA/rdtfBVHOIonc2qmskVGc5JurIrcomfdndFN2wGbgN+05wl
LrSUokyMqVBmAXVMHDkVBr2wA2Sp8lYKUVAwiP+zKGxtI5cYUAJlbW3UU/eCC6NL
8QwSscooOU5P6FU6BKrHywLt5RhfMMKetvDaTl7c6gqdSh+VZHKswgr8oaJuis9c
38Ty/hd72JA948NaTpmSaMlwzqI/g833h1Qy840UUwJ0FoPkeGx4kPHxVLptS/CL
p6SqWedcewTZKkMJK3j4g3BjLubU/IEJTu/aZHj5rRx+AvGfvEaVaaN5odjOJqnd
gSRKPpchDrCB2xUmnXZDhbw2hA0sJD+X9nvATWqfL2cT9BH4D3jOG4KagyCJbe+9
91HVEQt6602OCK2TXGVy4qXd7bdDZH3Mh3AFmHeqv5Uyae8JJheZSXNEZK+/TS/h
D54crQTp3DOXdQn5mEAXN4otBmmvMtsYVxDs4u3OnQaQqpghVed9EfJ5mpZ68TYR
PP6unpFG09uTw6y4+11zcg79PgBO46UwTmOElG4M4zAq8DuWO8DIxHFJoR6RPjsP
C3jeG7y5e9YE2WZ9OumKGgIAjSCwGL+8bm7F+JU9kiKJYlTTh82lGo9Ueg71Irc5
KxqmO1ofyEOufFpjhan/P4pvrF5eIX/d9fZHRCizwBomFAbrYSOomLz4SypUhMUP
RtzrQ8xTqMKS0AZi10+K6pXC5N+rfzuVjFTFfoYROLOOu1rkkdPXf3ITtohfbijL
ZcAEFX2ov+4bb2kMvCRKsLGdwSSXJq6A9Yd/VlEv3g5H8ElYIx/wSCB02q9AU59E
DNfDRWi5bbGW3nXXtQuz6pWjyl4AQ/676C0GD74etNdF7odqtaGmszr8HUJQkNrv
VFJG+Uz4hbKvqbxKL45jNV2XGQgAXBKOsOGzeps5hzX7ecxXVuj5Kqa9vatYTfvG
wONLQiqStzKOViUa/A9Rz1QaTzDHKz43FDqWbOZHqYMm+LIYcHuly/6CQ7H2HCYz
zVnHsSiIYXd7a3IL9ce2x65gVNV/p6ymqb/3aFeungITMn41I5/40wSpnAR8aWHg
MCSutbt07Q3oYcoc+GQ6crP4tRWBv9hcLj+Yj7fkOtjTNEILJykIguN/RQV8nmpn
i+k+CIUDReFmvxfDKWstvYaIuRaeULY0dqn/5LkB8qgGBk1sJgzedQl5z8G3BQ81
zJ9U6zptNzCOBKeYYWu9IBHSLITnAHFY0U7Z0BvbYWDzzuk/x5xaEMJhrq1YRyE8
3sPFd+5ALd/4oB04nBSzpr+jgQ8KQjta6KM6peY918sU2Fei3S52+o0AWn0mG1Qf
aHYeFvsVIml4Z7R69WP7EGTgXkzn0xAbeVDlnfqNJy6cf1GY4BCb4Pz+D67UGGMQ
PnNYPSc8A7fvVoXAsX5TofjXt7Zh8+vssh0J9MvqIUE47qtESX72QETcJQYzX3OY
DXVCPG9cFrFPxBKSlq8/qjT9k/Ws3DCvcc9OxLqSlnhvccXSE1uvZnOcxk6W63sp
RgXQ7JBXLiK/9JMzaKgQrSZ1NbzEHp1ruTPOVWdSmAnum61bq7sDnIh0ieVjIc0C
+Bo3lqo/vGir/3wtvgu5jY11ZA2QgDnKaCBeIN6E1qB2+Xi9wKyRkHd0HkUQgJ28
NWN9leG+54jELO9GUmcMRW06r0+sPXGsi3UGNpVB1SwkS5ZDvlUsUXJqi64dwiMC
ZP3+2roMN783VCTpNqOg44FnE3MpbIpIkWfnP5RFRYCwUt1V36PIf2b1vMTfgo0A
jPxN8t7/G1PenfJYJ68CuukIXAsr1BrjMnlGZxV4uqxMbVsTJ7oCMfpzBk/Q/YKp
pVfFBoIBzhaP2QaT5LpEF5Jn1D7mt5AUckbpa3DU7VfsjyCsa1p8gyPFdBKrZ9CN
oKKxPGhtqhazL92sELPMiqgshGc5C9j4SM50stpAfbnMDMMxOO//K16bUiEOoi2G
DXD76P2jcrI6LVWkGQeF48nAJQj5laLlFOy7IYoRXO2D8fdBfW3o4zQCPkVvZ6qz
/fYKGITnCQRPsHJX+QPcgcs35IDknx3ikgxMI2BzjbSS0mWZbRSh6SiacwEOyOJs
fJUxXL7ej2cxkAwpojPSz9nzJqs2zKUgTR7FwAYiD8/r3066wr7vJCyOxLq+w7bJ
iGWJ4mBM3VOcyXdOjNIwWtdYohciEzOFPBa7zbPtFYldqJIEDkZgsQQpwJxHCW4U
I9gXnVs4MC9nbWMl7jUtIrbU/KKtfkkztbyD02L/VE1tnK/xx9fkjvKbMPT5gAXB
eLP4+QPTbeGmCsnzGMoA6MhCIGoGB/Mi6js27cXbFl9n8kDj57sMgUVHI1niXFlR
9bk1Wcn/JlM+Ft+1D/cavpJs5ANXnEqd2flcGQjKawj3mdY1tZnjn5Vb7pUqff66
sWtGaj1gDgWsGTBHufbEhNJrp1syRzVZhaKT2sajljpYNtWh0HqvXRyWvJ6z0q0W
eUGmfsXbUgtIaLFNAdCHMGn70xDSIiSckKYTeDQO1gJQF/ySrVcg9yxo0zj37gbo
UK5PIBqNePPEUu23eMivPmQ5z+H0gbGkNDmQKz1TNAtDreU4+ZRQU3+QylpMrgtX
xvGrrl27JCN3FsMS7Y9pb9o4kYSdEdFcM1lyPeX4KySFWgmqy4ZSAGOdinErM3/E
m376s1m94Sj2nCeLKGVYFvu10goDugr1g/Kdfa7yxIdB6mNN+H/TN0qJzkAVsKPi
W+/iBP1Nz1+K4BVgDwGyb/a2wseNUWrRA5AsxOmT0Vuf21kyWdOXQ2041RuD73dO
KN+Pw6p/OGoosA8Du5nnEX0g42x1nJdyN5Se8hu2WZzyGW+YpB7oHu5P1unMF7gD
/SOGVdXCou4mqo0+dAJnl3OAJnDXkYh6nuVWwNeN3e/CdaRSfVlyvc1qiWE5UhNp
ukzSo8mj7fZ6y3a4sk7DQ0lONAtVk/PesO9dKhnsQkyF+xXll3o1enwh1WNi0qj/
o9Cw+IoC8KLRXZna6d4BAAr4RESVQHBEP4qrfrDxIpvX1+J41m53W8Q11umDjaqH
bgxr9ccOArXUfi5GHX31vRPT+SlLOQNLrmH/CCXnkfVN54pzXC7XzZHOct77DpNE
FAZDU2Y4ztBeKa4KoT5CTq9lN92cOAvltMuvE9PhDnhJkaarG4KBap+nqYYqmLHa
02LT51MYPX3ymqL/88iE5ZQwZ7x5MzaAepjqCUmEobC+GsTxMfcUgHhL4XPGBtNg
ulELuLtlBtXcfkd9cZtZ97KxujmIlkHLeM3iD7LBnnPc8kc0PsWlNSGXVsovQ+EE
rBMDj7KmFPVHE8Nv10CWtcqQeEW7N4JlV7HT21x7om+75SH/UY03tn57qgZZZl+k
XecHX53tD6Xh/Vi3b5ld3hbX8KsWEBYZXIq453zeBXTRq7ukZ6a4wW+Hg1BsRpzH
XBUZi9bKLt/bA85W4IhR03UD7CNYGPNSM58YdKs3vhj5scVXDdrklqMB+v0XVdgB
doEKPAdbwZeIUCxamKSMnVb/ieFbWCy5Q7V3z7679tugRHsd6CAuxF9IIHM4c9nW
UL7OXxBGKGttOHcW/btSs3erztb/BJeeRtABUP4vBojqa0d+790WitPCjiFLiENg
+2UiF2wIP0O7w+xqecoDJ5ypMJ6Psd/2ATsMNfoViGW8woW2OjIRVBc1la7W6wBx
pPT2HL/tie43kLxQ3VhgfgpeS3R4UYDKRNa63QljHBxczrUy/iMJwSIkEKhlD/eR
N6JtoUfbM4CEpNnMKrdVzSLToDD8xUh+MlNHc5mHWjqWBAUAXPHvgH3KFyFBk16F
tapTVMAf9EjW2/jhVpgZ0bb02w8RDtlZEUr03gpQ8XVLgyoLpSGvVJzcRudv/dpj
LpjlJmd9TPKkG+NHUx+KCYN6UXpr/gnb/0qfbhyOJG8Z8ToyvG/07MakXHV/9dUj
s1qirQvg114q/9/wSPzxRxBW0pH5fjY5ZdhuqSB87yynxyDe4GS8/FZLqKGGX9GA
npH2tN5McSKK3HyhqnLwVm5/26T2Bk3tF85rrG389Q517As8Jk3Aimc1+aZT0rqP
dN1Eiy2O1dNj8KOpPLURY8Fsmnv8OU/AMJWtDwna1cWr2Bi87VrBPlL4zpRayvWi
LL57K0+Ut8R+BpBrc3Gfg/pS4GQ+LRUbTIKn7/ycJhwnVAm8A7wTqQL28oVSSxKZ
j41YZdsmgX2mshqSwxjoE4+oWCOkgyr5JsoeXT9epqHaeNCcc/33giKPaeA7Y7Hh
eavYw5oN2l6c6i/nRnoI32uxkOziVHbSp8fIZ+zpMkIN+jJCYNJVYOcpFg3szbWR
gD1YSQRzQnz67P0Ue03bFiiQyIEU9ZHEXr19YwMLTHMC1+E8k7FTWEkQwfWZpL1Z
o0lQ3bl6pCY/G5pfMZZ0WQ2P9mKw33I+Uq+IcIZKIyOwRxCurqsOmTa4bcKsyfoa
Nn8B2JLmdO6LoeK89L/MEGyXFbT/UEMeog61x7M2XS/ChBgjFp6Xo4qnqrgQ1aU9
FhsieUkKEY9hy06LEmCG4Kp/PG/k/+eZG7Lv87qPVasJtyyZTyZA4t+oPgl8nr7O
OgSn4VrohJZn1fUNsz3yb6wMpm4uoL3gLJgTbiVSyGo/DXiqm58syv4HIbqPucsM
vTGyUuxYJYTiljOYlM8XXlB5drokGZ3rju6sU0hJVo6yi5/6aFjCSWBjiTWJMoU4
l0qHS8650nWAy2LU7jgdd1SOPmj4I36SNuuv7vTultvEDj7Mgpo7oUySZtm6zkft
7AtnOVaULfyDCAUZ/lH2XTpg4s/3nrT788SgSc7Zs7ZthKjBh5A2uoZocZQelZNO
xxD7lMBPO5c6lf44Ty+XM/fMjssjWXRnb7OWgH7V5TGiAp/2E0yIWALuBh8VM9DU
TSfFnbQn59c703R7GZj69i3tfRPAjrrTMLRwhEtpnXrL+sTq2NDYrt0KNGO9bIzz
MlD1xyZ5mZSGsYCecjZwUm3aneQ41KCUyut+9T/c3HqeIY4sOVKxTaNvvxF6Hcbf
6Fb8etpKHhRrmC/JDbPVlZ7yg2UeGSMc/B9e2dBFQ3kKj/C7yUZ74XdNmVZ1pSor
ZFI9lmyqTQXyIS5p3fF0reVTduQ/ve28VCP/Lkm7lEWRzmZa6jf+hUh7UXeTG0Ut
jDK+G/56LYQDt7LL0kuKbq8p2JGNJ5+tsDjqb69v2N1vCatEfoPGAt8YV0ea890z
Jru+Flnp4gz4GmEdMoMZVycQI9fJQhroNbgn2DTd03hQz0ms5pAJqVL1+zJrbAb6
R/AZgkJKz1/GHDDqC2OlmHkifZfMVLfn/iaD9BBzfybYvsRTk96Z7N75rC55LolA
gOxsvSWlN92CVGZ5IfPWyMyZQYkfZvTjoBw/AYzdtLNEheNp8ve2qOe1M0AeRCno
2svXvXA4cKut+V9lYBwhnl1GvekVZWiRahKJ44AK82UKZ1f2h0AD8vHY8NxZcmOH
8s0dDv+S9MLq/E/NpzwmDnTT8qFSlrnoU0WLKHUj0e5WXzkZwufUZaSIHMIkquwx
xffwacqNIjU0/KxzZx6hHlqQKsPLOac/SgC9ODJDyR5jVw8SzDDrljLBrUzpSaFb
VMGCDa32pRBuj8NcEDCvLLe5yji8qWDwTB60QmAPrJtw4UMBfsIZsFreFsAX5cFa
ww25M9l4dswkUY+Lm+XuI8ztw4gkqcbhRk0OKgAEqiX4z1PGOy8rwNbJX8FzUtiG
/ZJCQ2vxWtnCK6+oW1ajKe86kYsQs2QyH63JMiRrO4PM+mrdfv5nW7x4/oNNs8a/
X0dLzlujlGlTwGS7xP1/NButASWsVpbkRPhOdS0u+mRt0UOYNguwTQOpfXH81aCd
GBJsBI1FVul4NPL2fDYF5HAEYLZAFJrRY4m/Z5xNWul6TgYRlYL6TR38x8xgC4pK
K9CxKyU2oQJURKs/BPwA8HQear2uHmaVm4kT5uc7Tpv+MyqEzmPn0LqGsJHnXYut
Ymnu9db+WUaaWBkLmxbZ5sd0i4V2/W3MjnXDnoMU5lgDRnqGaHvvT3lcRNUnhV94
YeXvNIFudziihqGjfwjKoLoVaja7KRZlT4ggBAQaDHleWHnIrAr8HhOoybq+aIfx
tcHYBljWFewb9y14MoE2F47jz+zFy5u/HUpunPE0BGB8PcjkKBrjUSVlV4B3aF4m
JFivxhvqDxI2dWFop6ATDp7ZQ7TVODOX113jxbcle9z66z/JU32FCoP5ivxiTLmx
A3G1CcnrfCosbV8x4CFxZNJLLcdcRsusxdhXauc/xBQMomNRM/4P9eqOfUp2+sOB
nHnvcFmQ51H+5w8yp+svmkBxZjrAyRptrrTaJXq0dar9h1uP8GRqKOFbfjz9aO6U
8JyXOjRZysjZ/bj3vs3fFEdZrDUyOkeFZSQd78WipBaVCZyhWgicrzqStzKXgkwX
RBbd11Z7xgFEFpA0pvdCR0tHJyc9LvzhWMEfWKGHzTA564QNjm50/L9AfwSdx9nO
zWpS6jDBZZ/qj2ljvfVg9yyJpZgoTgutl+727M/KgoDDJ8gCzeynOa3X0iYe2zn+
34a6A74RPIdKrAXH4CIjy63ghVc4KeBbnNIis3m3cuiOAJZH9/dTGIrKiqPhcn7N
ZItTPCFYsiF93wL14j1WnkFv8DdwzI2bQV5Wd6Cd8v3jco7pfcCUpUrcgUgif0uq
buFVEsh1VDpagPGF5f0L5yLzMiZ2VKDVeOljRrtqOeZOG/HTeLZREDa6awl0mKDF
0Mqs9vd0/0N4WnVO5fNB1qU2THWH4Pb5wZZ1lThV482FlTyuoArSaKzc2Z+rAsHQ
IcFhFNHXmJIVO6T4w+JL7Qds+p84HZo7HMZavYK0bLWaZyLx/Efi2lRBdvyi6ibS
GCPazRt2jLa92QpM0tBQLp+TkEGyXKLsdzG5bxH24yIxijoBcJWFWbQ4H0rdrSQi
VzxfUXrE81edWpI/9MFFa2QbtRNneBwLBb8Uxhs5gdJB/fX2ooQFrne4CCgyWtp4
MXtoUoBk4OLlhEjQwias7VYyqoWbboYaPXO4568rrkQK4WuOm8sPWAyJKF/Ybcsy
OnBuSUlPlS9JFwxMOTfuu5PS3yztV/Gy+GDq66dec/HX79BqJR6SQUZkeHjdIzhZ
FTH/Nhd2UMMceAp7DyQ+kaAhuxMUzzm5NXqzILDs+aa64WbAytOGSzb2w2Eb/bvG
WskdqMCp0MrE7mchzIQW55OHmnxRKuW93cDHb0Vbzvh/UEdsg8ME/RbkS/Roxfi9
+BKJ/u5IvKsWG1oPYG7KTmslNn0aceRwuyE07b2/vHnkPzhk3T3sq5P14rj/g56l
mVT+h9z1hSOo8N0rBrIDWxEE/MIwgNS8hmqPIuVuEcORsQ/nSfYnBP+ZT7Q3pZ8j
/AbWERcz3HUbCFp8I73AYcvykEb5M3G3qfY/8mAz9GcgJjqYJ6n7gojdLz97j07Z
OZhnooMuY799ZFB+FEphxyxibmza4QoC9HEAyNmWquhncbg6nrGVE/MVZyVtwUjS
2ULHOzlyH/VFMU/OBTnHxAxbyUERQ7pg+YY9SLI4tBU+F7NsjqvyVZCYZHaTAGYc
d8SlLbNel6aikfqRbmawoXW7fFK0laFbRdSTvRLnIbwiPqL+015Ou9HOa6JsyBKy
BawaT+cYA7vwIKOwclqau6HRjZ4DtdW4k/aBi/OHIAr8XlpfLBshib7HDGwarLEN
1yd9nvNb3mukUVJzjgMF+nb1RKfwePXKZFPNIBoKQf6GF7icceNyPFNwGkXDnN3t
vh85B9tSMfL77dWB5ojZsitXjbIf1ty2h5zE1U2yxaRVbYz09WVwAil9Hr0ZRPm2
of1gCi7Tiw8LU3kBTB2Da8Wt2j7pOKkF4PkEsb6+CHuQhUSKd2TZ3gfphFgJql6H
14fPQdS2q9/fWRj2bsl8YetQEqBv8hp84aTYCm5hTQsNJbH46kTF2NAqdWau4vVI
ioZWO5CXfG2KPupqN/XMH1DFrOoUveV8q3g5qpv0atUEY/am7ctKSs/VheRisrIY
sF/GLRlj9B9Jq07PgBpKMAyCYRhjQVd0IZZqpPn6NOUxqGqw0SwQ7YK+5yR3mAfw
RcIuokws9ruEMYk5d9QuX4CF/puYH2aT8lAFA7EUjIPlHHSLjB9gmvUJ3BZrVZkB
0HKzChYU+cHwW9I3NCZ0mbSpvlYYwOgJQHg8vy9UZWQtPhSmw/KdTRxLTaIxg2Pp
2Rz1Cb6owT9MmAfTUXyi7OQ8lH4tBCng4PlW7+5MkdiB/Rgvjn6sTZ1MN+4PrAGR
313u+ngFjm2pD10GVse8TrAzrAM+8h8jIPOrK5Lc/p1OvjKDD2P6ingcvvDuuPVz
7ayIWz2GGgcnng+auUgSr2leJMzBpJ6KgV1dw01YezOHttU45C1EjPs05RPDmvs+
M72u3aqoUoO3u7yrafatpySYXiAi+r/3SUNSTF+pnmZJobW17ZlE8Zb+zIIDjAE7
2I/tSUe8X9Zv2UwCfkJ51RCIeH4oEp7QSzr47XkK0MsLMRWCnFZBzWqR8EVhw7Eo
guLPim0vejy1ybOR+Z4+Y54JN+5I433WPRM46VMfj2dgiZKOLndkZBu74FVQvkiN
KW3a+4S4FAHgTFKriIqlaWNIR6xSSChm8bNmc93zgZcMWysR+6vj8guWtu6JZxsC
Nu3BSe3JNaPL44Lf0TgDwpS38q+y8+L0oAJZHuqBLctFkgqenEJQCrJlSTw/oKkB
9kL8v0CsUWvnW1EZVdsj7j8DdtqUBHlukrkoNlnza3hyfHMa/ll8mmdYOXl1nfOm
kwT/HZol7sxAeZPr8hZz96FaE01XeYDTBVky3MIaLrALgMU/JMdX2Is6qwnRC5wD
GuS41fexhoCjEdA3yFEkbqK57jFHCqUbf39TFAMT0Qgyywhvu6MOwjFmOaDDCJ1j
oEk3kQq6iiTrQVWyRQ31lqkUkLzFDzoI+wt20e93Mf1B1/utCcWSS3UbNlrnl3wO
zXJnf6NIMXa3FFz6HcgVh5UlpKIMKePBw2Uzc4wUzNS6oZ/HaFJmV0n0avBJxVmy
HRb5x30HpGbgsWo1S0j/hIsZJB2/RsCpZEQ5DqSApUhSTmU6o2Yv6ptMJHSAfW0n
JM6sfGHO9uy85c9kDGondn96O3pe0GxRz9rIQURbmcMgEpoxtaB7X+ZnoHiAzbWY
oDzvDpH9NvDuG5ct0JS2P2Zm8QYZI9JSzWEC4IgEdTfzRxPJBjgdVQ4/+0kf7Yaa
DVaWAN5p2kA7YGCBY5fLRUIpdIRsD8ttACxdILcHtlXaHIvNkFTR5uWX5zWM4ipY
7RuLB77zWL1wuc9vxfMroD0L0n8Q1evWuav6Km+RPvAxHncHq1FmWn4FnsN65GHn
U5MeAoFudmhzZtg0ERRAkR6Lz32nBCcR5jJ3CpfMvAceb2nuWatJfHh3VxcKfgMs
SdpTZMHXYQ0qqnMPh0I+wdRaRpVbRKjzdDI4JHZ7yUxaXzIEk3NCXiI0P4rVfQXH
SJzuXn1wyD+Ekt9xRuA1OmfGWHCAEUwErNDS1Dr7zDDsGtct2TyRdOd2puluGqSD
DbCtWBPvbAB3tDsM4Vr6JDkmP2JJbuOQfepdDJocIoXPrOMKBel7HW47bJknbgL8
WIQOw7R9cZxZN+UGKFBvijA+kPgeCA2LkNNZZcWoyv7gQvi9rcOBhqLeHg+AcMZB
Dv4qwhEOIkZbSKD1hNyFIi2uRY09xnfNkVUTLUgXXqjS+iRRc0twIOHpBrKaK9r3
8LMrmsJWPhC7znH9eDfRmDtF4KiXSmccTJEnknZ1SeAStiuXd+dLhrGfWhsJHnYG
BBoWyqqIzuDe76Q+zz+LIhG2839eZRVx3ZpyLs6+7caZ01LTk+1sLC+utXVEBWtf
qvV7xdyjoSPyQFs7M39faux8dhAwMwi7U1eb+mMFFrw0jzIWQc1izhGKYr9jCnhM
TBgxrUWOXX5N2zJZUUSp9mvKRzK3ktzskanCDjejGbAWnKryZXMvvcUGBygCEYwH
cHkeStXKyemkQYvZETCShRx2bGdFHpNVk5ZvhPdSlEytLB9zX5jYXWFHuNok6sfq
oGRBmqqF5HhFVxSc/K4OZ82tMrWc9sbxByUZ+e5P3qdfzjTQYC/qELS4sF7vCDjw
xBfvFZIac0ZFvZK+i3NV44JjiAIA3sU7v7zW5vTOPaWoKhwjuY7hBPMFBER3zjXM
+JWcBAefDcUewvoDnNBgpjciQTdF9NMcddgEpK3WhYHa4LY414EG6r9sKjMzM7oX
ZLSUBgGZZDUc6CiEZnuo4YaA0EPXLr7bFOe0GQ9WYeyBkb7Y2JmTiwXlrExZ8oFd
N37eGlKCZjIoU7QxSm6N1fjzimiWCYOOe/Wlqs8GCiKxDcyDMzPSOxtLM3LXNN4g
EUaji9zCB1/hkjhtFvXm2FN3+vbZZ91CrY3QdrYW2F7zIxz6ewmuj+gRM5a+B0Rr
34C/VJ00XwmFkpN2m+EySvtacI4KPO/wWfXaMNkTmNgBu8f1f6be3TMqhs2lgmY0
pKd/7AJoQU4+aV7sbAPNIQo85P0yFI58r0I38kbfWcLWUpYWq6rhvgI1Egmw9FT4
Fb+ncmFCC0RX98T2wE+gFFya0NGY0Kto8C/kKghxM7KIt4ql+nVS9GamooHXuq7p
F9pTI2wCyVv3sEjJHwYLxaZ8azVjSBjrv+X22yhrQeZMqb0TYka4Lgni/gk3tRPD
/NgbnlfYLXhQ731Ttqeuxetovh78xU5bEppmXGmS0za9+s2yQ6EA8htSXp8MFD/V
WTAK8ODV1VuiH8TSzZN5ztdVlrmYVE+jKBBeRmYk/WtE1/h8h/iASqIDk0KuKaVv
fDJY7vrrLdSuSCQRUaxmi9XDAl2zowIJ4LaoS9FPJSjJ/ucRyfGf8IGhu7BZ1Jy8
/FCDuW1Ub8VI9X1BJA9LORZ6+U/jUBuEFNksJ7t05uoBiUZEH2uUl+7JfB15fTuY
IKsubCmviiOMKOUSXeK76/Ec8jGbygQ6vZNMWL4vEaxaY/42DOzy9g3+j9ZFDPx7
Yhj3Tj3fjd05Gu7WMXSggTjPObJd7ZNx/30ZA6cdmqxusH0tc6fFHc/SzvDdLH17
Kzh1zvbWzcJVITGChmwXOr2USOsbM+H1+k8WpBYJEr8+A23B/85Ug7DumHCIHGWX
VpvzAAZXyhFQTKHb5wKBk7GGkgzfacrS9BS19srpX0gXZzxZQCj+fsqQSjI0HjnV
gKDu/Fy74v2LvGY06T155qrkoFkSzHDgZYW7JoZY9ueSvbv7ar6lI/govz8yJRLo
PiZ/6h0oFBYOMFkqa7o/5PNqWuxk00lQkm5fOhRJre0nGxG3QRiNy3Lq/qPAzcku
ppCjBSAjhd9+43qbCKRXAtWwJ8u1YXpQsjt+o+2m+sXxEdx4kb8x7T6BfmmxZ3jk
BIu9jjPjEHX5kDqjWqgUSUt3Kitvdc0aDCRxF9hrT9JefUxODPF70x+8IW4ftBV2
2anvI1xVk6/Z34cY45XShFmEJ0T/y9K3DlzbT9PUFPe6D3s++Iy4nevsTYBR1cYX
toBQ/bwwCeqSnaPwHZM4OXPffHu/01nG4QeydEUaANwOiFRy5kkfVPf5NObRwcOw
/qL9g1t6tFCwSlZi+gYyGopYoEC+cvJtVwVTNs99qQdeI4+LRYpGRAeoxhWjGjSU
tNM53W6/3qpfMZ6140mCjsYEV+XPPfnbzNhPJo08lJW5QrBlMzcO0uOWj4j5nmTO
C90iXNykSkG+zA6t3u+qmCfqwKlnCAhLnrix4x+oz+O8ZbSIsSQHjgUFyvJ41bcj
QCDcQh3yCpMCY0KWv1Ntf66OOnMI7Irw+jEp2pqbXxs/OuDGI5yUEArIYwYRTSV/
7jEfFPpmWL4nh5cVMf6xg2JGIELkwYuKXP9XOl3TDhAjZsv3iwBlanT0wshR4XMj
+isYruxxKHqpV0LGzGn3Id4SBna8EMlx9gbDv7qVpw5bBTggbzOBLVa71cKCYRvP
9f2izNBRATWXhsA/EUrnwZtH4MDmnfq1xiGHMj9RzGHcYUTKAs17/ZGy2z096Tq6
0lajNFlA+VEihSNCx2DqyDaB5+4QGoATY2YIPQQiaCxdu60j6x0dAwYutQ+5AzkM
6VGy0DSaQHyGEr6HjqpeL82zdYnWVxE91JuyUHtncesG++K4tFNqqLdp/3OaJdg7
uUDiv90Yl8+q5WbyUB09Rq43kZzSF5P/VRz48VpGE9CBZtb23Y9g5N1MRmH/USpW
kQF0ROoScHPWfv9QTYoyoAuEQEsra+G2wcYQ5O47uio1at/49LbnLNMpaMiZgMyt
ih/0kAPdD2vjVgVSvjic6f6mqoj0tRsczjTlQv0rlJiBKmJt/xHuLIsXJeUzydke
51waiQ/xW9I/g+dmhG55mDpXLIoriDnLTcWx5GHFpRJVl8KeOdmlp1JmXg1GZ9Yf
0OGJYvgdaI1/m+6HTK3P9HCEQwQrV1/qnTdDUEWPzkUyJhtVjzW52n14E179PtXS
VAgphF9Uo0mug1fH+VnQPdZD8sG6uiZiKhiYGJU5fg1L1/nfU5Wd9o9Df6o3bBM9
1naTxM9Kn++te8tijZhgdARhZA0DVNm5noXR14wz4c8wx6tobGn+ypGhSiqFi8s5
L3x+h54+FC+zz+qF1p3nCjjs3HDCnqN7XvkVyAwv5gKC335QhgxB/ujeCCUpoUKS
c9HUdqrNT5lqyCtUiG37LDaBLDUHS3LJMabUmHlFnSljWt6Z3I24lLF7ThJabtQP
9fX4ThRvgw9VKpgtxEDZ5VqAR+mAHEjDroMX4m+RlvaOXKDJ4bzjOpZlXVTcWJaS
p4nAKsU7qXg9R1ibq0Oh0DzhsAplODjuvnBkGuSNtYd6fpk/mGqLxVzLGedkrJd4
SSXuUS+f6GR8+HN0C75Giuk4Ibzw9JLvDrZ4Qb9Y18BPkFUWdw8vxbO3Vs4nCfim
2sZ4l83z1aLqEj4YKIVpo5Z5Ow0ZDNcKK5NSh7KE15UPKoyZxdxWMr2aUj8KayjY
V+gHjTK2n9BFDC30SwKVoCo7aVuTEAA9KLsHKbtG2F2ACBhfz4gUzDHSlQUyZzFn
Od81fVcfe96v89lyyMMxFjlz8xuNshXqiDO/rkASfkXrvmBKaDNeWrwSkvVtZyZC
n7go9aXMfZnogukeR2LlqBDtK5sea3SiBg/3zeYrMtgwvhYAoG4C8W5ZHZ6DZKDs
2q8xLAbNfaAE9IPSVX9NA2UqzZBG8Hd071D1VQj0jDswkt6MrtMpe8lof5moN2Os
T/jZCePrUVbSB51OATYME5aX3Ek8miYd9Xcm5YEldagDO+5iZQUuf1SQvjstsIeh
OoimM4nvluAzfnU4YlWZHjWeVMCWgwXClpOr6uOzaLcO+s7UpmHrz2LdJIBaKCbe
tY+FKW5sxkZGrG7eDs2L3twFUsSMTe1/c2YQ3a5Jx9c7FxFhCsnKjGmIshwQ69o6
YFSXVCS4TophxZDFXRpmlqcEvRFhwtsislT51H+LM9koRJfjaVuWF8p8rg8ZhM9F
1GAE1zOZpBMj7Pp/z9PYoZjCRzmezKrvf7wuRzzSxrofb2sjXgrsNkNoWwRcbBIC
/W1prPNBbeWF+YuUTcyW1Vk4QqMSbUCKvLBKqCpQ3dEXmaWZAsHUBXPCGCK/+7GM
B4CuuFdikFy6+51yaX0sSDUW354GQcON3tg+JwMoG9VHCiTyULJZhEqCiW9NlnD0
EQxIJTSbau4D6XjLcPIaIiwq5jGW9xh658sDOMRpATPz5uLcNH4TnakxOsCJlhua
Kd5inzQJv+TNAY1wMD2whojzvkOcF82k4H7cTP+h6SFamIiPx3lW9Yq7KfWSBFtI
tIbKbX6d9IAf68JVwY99VYxJpWkTFijXHFzAak32Q84DRhlrxiYOrZlVKeo/ds67
oyB+dMyc3Tn+wGG2bpDh6bI5LZKxTVM4kRDZd9IoQVVXKWgUHTQEtB4F7Ydvr7gA
EgGpAWrWnsq1HIet7AoKhbhacYJ2MRg6aXII+LZm3NvO0zs8Wza/4KGcQaymdqvF
CRF3QIETqFALIwVKoB3kH5U2HwQ8rAQoJKfgM0jgrM2Y7T4tDavKmmGIggUilHDY
aS6yzqXb+xU96QenJrzVc8hYX2WkqRTPg3jsY2M/8rSCQYsHLM3sT1bcSDTePA3r
1/rn+VGQW5vSmFl7vHLNGc8kPTdoaAaEfpcAICUVDQFxS/brfF3+6M2Ev08wK3n2
2uktidkL6xAiqo/Lulp2lyytgqWn+tE/hIQW5osCICEG8/nOaPmmRBydhzorU2gc
6YE04FW9AKEqU1sZuNkmtZeGm3HrTDI7rd84YelcES0g5JGBc4h7ayMysqm+eMOV
ejPpl5UrU1sxRPmsH1N6oRIBomiweZ3FeRMq6h7T/H95vlQ7JoyG+rX7xjEWLLV+
u1yRlSwjfXw2oybNJj16BgwBi8FOm7whXH7wNyLWMb2eKvf73TLXer96JpSK8O6E
cChrgx13WbSm6+dTn9EEjpYxPIS2/bk1fiynCzWnRgv8Tm7MX98iYnVe7vMXAf1e
1J1q+kb0ahiWVEy7N73VX1v3IsFt4IhP5nYRKsKJ812l5RKDeG2WnA71YHitpXgV
e0DW2vjaDTmgWIScMCIJYtTayq2l3u923Ye0J4y7IJzkemuQJb4qhP3hnreCtRwg
8CQL+wSQUp+yEOKalLWK8sXDg/GWMqVCUxr7/ZDEAds9Xwq2XVXD2EuHyfWBca8Y
N/C7+KOragomMEz0HbDtCurw0q5D60VJaCeFnybPMkHrA3D5hh56DIfJNH55qQ7+
Zk30z6t37h9JBfRaBynGjNmNmwQnXw3IcglaglyhwsWe7vlAfVCYUJvhXRrIP9Ks
U9fCLi246+7N6sIQEQiUiMS2ax2qFN9gfHniU9zk2MTR3l/0BUr2uPyPUlPkaUjh
f4LNmyYnKH/F3PMeqYqITnPk/xQoA76fqvBSfa8dnEfUsL4TIEX4so4PIJVJnTV9
tGphSzfa6/dlkjNwCU6uUmLE/8XZIkrNEjejIbEeiVH4dMD7337+QR/HrWo8fVwo
O7582KUCaVxWJNYh8Q91gfoHDcFv7lw0vBcfq2U1O67OSjZe/yZVZDN02gGjPG5M
ThWbkyKZRdhCP7WHxgXiVNmrCvehbX5WQFKfdUn3zkMNB9eiSW/yHWaerdAPijSw
ZO4nopJrITEGzF95fDz6ntQXOKn8MSL224BcWKFe3I3wtDgy6y9YOGViOKgNT9KH
mquaHl8tT1wFOg6oRG3BXKu5tXhr0n8Y5/AWp51mYF6KvDW0XhxHNwci0jWgJJm9
Zes40wN/7Cy3eXABtPfJ3abgig08dynhH90q6Pa38O8WrIN2S95K3BYSTOe2+/HW
hGzLY4ARs4knjQhGxHYzoC89wC8NDiD52QYEKEXP9XOxgMhjHYUYzRmLeIeB29IL
FbuMoOhcI6JBUYmjBXm9l4MRO1L3aMzZaFckjmbWsO50+krLrXi8jte8D0Fu+y+k
9i9qwhxxCRshuEZ2/+T7avXlfBGZSEH8t3VuNd5YsrJfAu1xlRnbWTOJepxKu9Bo
6gGOH6OjVij5u1WQ/QB+M1tmglRMQJPMGr1Ranwwgw8iTE2tB2gQYW+HzUbPunLm
V6jU7TpWJcOUzud6No1WD1mIl2m0w3Dyb3lrwlfwj+J1cFc2yoSpT4uTlEV+XVYo
2FMcC0QDL9d5bzVNWoIMrscNlgdIC5Px/AtqPkZmf3RlEdHGeLCMAVTw+VoeJMDo
27VSjO3qdLhM/WMLfSexfV+EMcyWfDQmjYCY2CyZFMLatJwLfvOKJAAVu7yVM8wl
H4JEQKgc3wHHvfjAZ1YjBWB/Wkbd2IMueeFe0veiDT5r9hD7iJZtjynfpSs7tMwS
2Yve673WMYEE6KqJJ8Rcl1HXNeEzr25Os184TxtwCwZJZ4tg8wWESNR/V49lvdZD
LKezvpairpVayWdCR8t+HWUZcqqGebs+XJGcsKp1sTuzhSpAgKTKxd/VeCBgZ1zP
lwF9v8mlALYv+4dpUe2mZSgN4MAEIigayERpM3iWU15q2XRcn7dD6p/EYBP3gq28
nUc67ez5f9DFyrul5lyMTqcQvpoSyk/ZuchfPZ1IfkESBs0xgoRGl+ABKvF25V21
Q4Sl1wYlZyei8NaQF0YMyl+1OBNtoVUPEs5X2aXavvDTpfoRmoQKth/S4XmUJrEM
Rdh3Sk9RWV/5R1mOgCyTYwk8m8bFOCpn8tOCtSVfhbblhL4FrfMYqhqdFOIArntv
sJ/0Em4ubtc9Etgs2/n3aYxGPQLoKr0Ivj/uBBRLDqnmXLWNG0n1XlgKJE8q+pdk
QSpQhI/QegrlyTr9TmqQF547K7Bng+fGK7+cPgXjiK5Lz/U581TeO9R7wiTT6XJL
ek+ScUKWwnTTGiHfuJskep8dsNNGVrnX7J8uEg41fWWxOrD+VKxpN9NnlRp+inSo
qqVgoLAl1Xw/YKFh90qS3/rHEZq4rokaS+KHx+U+tQ7/K+ZTmGkKft/KDd1LU0gl
jtNgduhwxohKXGEv7mnCZ7TxuSKgX2gvWRWU9BazExVa+zZJDTtcYdJ7rn/nCIn4
0lxbQSt2Im/o6iII8m83NGs9FA1RB2RnodGaefKGRoY26EEDltxHQ4YLzDo4KFdk
sC6OAicdySBcNOtA5GzXvMAyJ8Otpy3fHCkxWsHBpvvpu6XaDgjUsuHItZO9x3uG
vva5yjSAtBQObARqFq4H4rK+IuSaEcMvFtHdz0WdQg1pT3mnmftPVKBTtmJHHUi+
AAXCYseZ8EN8fglWan+m3yuF6umZKC1L24HAZmdfPvl5WZycFRWb9UUmfBmFTkEX
RHtVpxE6McZoUBCG7+qLUtT3nSd2bTg8TathNDscfvZ0VXy3sq+r6+JGsy9bcaSm
1IBr//+nmoVkqk3T2jwbWEM4kw5G+TXzW31y1DxodEERbEeWeD/Z9xF7l2zhDKB4
MN+501W+TrDwqBVUqiwmZt9Pa4jv/4OcpbNh9jYfPNLTZALthaeaeC+TBo2kMgmT
Q1aaqzuxbIsI0fruEQF3Yd3ufwTn0P9KfofNtwPJhItj8mWewKRiv3CeWseJNot1
pJlM9pQgYJhf6qsglIN4vzQUdrGjkscvqzj34JeSBDmB995I5tY38VgbnXEUjwqJ
CzrOO6PR9cZ0KLp8vqiwXhRcgXg8zdqe+WTvCWF1DRLE0mg+Iq6L+4qByWnr2ymF
+x10SS0zcN0yFWPTF7DnzHzzoRej++Kn4LGtAB/HJmcEPfO6RwIy4I6lj7BUpcLH
9d3Xc1d+0Z5l/ka/70HSBNPYhtH3CvE4Z1Iy/usNh23evoq2iuiBdQ52/FiOUPLD
SoAUUx3qCvSzbI/PFf/GbSdBB3Ww+4WCSQEwOzytZ7OKqgoudVeD2VVHjCzjEKJx
CZluXkgTuwc7HRXAYAjwfVwEGc27044gsKDGQocK0qOn72z+kJgIxIE+5QiwthiN
SMcYa3SSgAvR6y5OeYsLJQ4/Ly7VbmetjrB/pe/A3xYyTPuMdxnZfEUY/hEGnTcR
ScrUhs3VQrwPaRTFy948nNOISyxBtxA/CZQxAhrGL7hfey1Xro/cDdiIJzBrVl0M
5ogU5Kes4IrSqnUt6AlrUDxJesWRlzvTN4EpTBpiZV1vlpkRapywSmsuAYEvRvo+
kHnoy0BsXHTe2/qY3kUsVNRARtObTD5uLc+fBgFkTuscX/IBQgUKD10VXp2edQyl
HQHv3rfNYyO11KTfnLmmhlgYb0b2urAflVX0ugbO6jEddQR4ZkBQzrO9SF73T25p
Dk+n32/6Pd38Wv83lTDRb5k3KPPjcIVD6u30DA3FZ8heNqBVfRiCz0ZpCy5BcIau
1qS8l1Lja9kr0ovr/vWSSnS2WzQFjtSte4iz/78myud47gA8Mua20N/a3/UKuYOt
hj38CCRT13o+IwCuOydxYJm1szp0p6bYB0GkyTyJ2WNvGGBKjlK7FpBsomXV8SHp
2/QFQ2OqF8F6+dmlvSRLsnAsCWJ2uY/APpom1YBSqvnjAXX/SRfk2PNLlD1Q87Xw
kAmfRwxUPdzQdbR6YvUeLk7qgu290t5QJD6saYA75XVNcD/OVabEU/z7KrOyFIsg
KGjnHCPiofCG5NEiZlRODXfvpmWbzP48h2O40v+bjveVRrw774fBqjbIjIKziIFW
RxIvY6r5nVwqlqIQ5buQW0QINDGeEs5IAt66pnyjjgIJTf6PMf0xm/TDX4n5YA3f
fHYmZfgjlh8odDraY65Q0Z2pAhsisN8Z2V/ovAPE+GCbCLsb2McPiUvTKWmdCyRD
uoWJYR+ObNV3Zwb6KdAE4YIEfzFD1MBfKvK1sO9APW9CcmUsCaSBRB8m1RdXHIin
ZFziFHbipuIZTZQA4CGzBNfiyNiPKN3gS9LuiADYTOb6N14bpPDwt43myrMlUvWP
aZNtV/rwD1UX/en0WavP61NPvGl0/De8BEqYa0EX/6wY9FrdzftBkWYy8IDVGI67
AfgCIKPl/FU9DaTUZuXw8X2n0ZwzLJ/1gCiqeFvgX5s6ENgP7jKbjFmF1hMUqUjS
Y9o7R96YSN0lvtxOIqzX8CzvKVyO0hSnBHBJ5PBw89wuw16OaNXsvHyAAjuiWAdM
bl8/u56TF2AuWRy5iMNMgrk8jPzFBpuN4PvPcSpOUz6VCqtAIajxIHhZs0lzo7AB
evW7KMSHqKr3FK10u3Y1XAJoJWaaH2HVaMt/9qi1HsWzRu8g5zKIrjZdo30THUyP
emTG/Iwx4f2IncMal4MBKdvwN8EOKdO6wUa9EJ7UFKJXj4UmfwmNjv78aNYOufeg
e5crulU7MMUKWvgWIo3hZB58jQJnwAjkukHphYpB02z9QhAh1UUgms1A5gUjR8O/
qNZcTDhaWqkSDxcvS2D/J/5rO1sWd/CgXL3B46PgzF5XoM6RqWOnc0dQheJ/7BzT
uSsqSjvuHusOO3pKySn0UxTOmT1MQocRJmPeMt4Eyyi/iIEP6UcvT/GmdUPhHMWP
7jfjtqtHYNNHkEWxEAlGmCEP5GlJG74iX4TSCQgnqyZeeT7VLPO7OA5T41EZ9JPL
+unpwuYsaXZ3SLp8gF22WFd+GzfzkCVqphU5lQzwBfP88qywgQcIXkQORm8ikSeT
xhE8Af9SHuCgvsq4gD24RgbDIRUmwfkb3CPISubeuG5d/B8Ff8GEc7iDED0Kw+EU
yZY3rG5qGSEuuRrN+9eCjuhJgC21+nJ7NhqRadDF1R1kQG8vvuMaTtQNZDPkRQQj
VXdIMKcT7FjaT3hZ7g5WluN0xsTI2ARhEuhNqK/ReK/mw+y9VNr69DlE28yCZnHe
b8PoVQu8kkRtUlp7e6gmRVLBhgkafC4F+BMc+4Zf0Fp4f8hApnlemsYybHtKxh91
1U2zbbtfVyKHve/BaRViL8pwvejo0zuSYNst1rUabSVQe/8Bf4QGANl0KRs68FSJ
uo6PQuLID8B1tsyqH7bkQyKHhcJ9EK1VKCU8VWeI5y+aG6TdsEbUZndABMBRsur3
+F+01WRkrwKc8+R+MR5dooUG/Pqt56RiTS1HwBfYh6AGirc2gmYqCf+pu0dHQOmX
s17ABgKrYBGZWTG+8X+D6aPWmtWnFgySAIjoUUGl+vMi8JRnRuTOCs30UBp2Orla
MSYDW2ZPhlQchHdjZ6bid+pbkOF62E3nBenH+CJLzP/xkIoXn/7xS6Oz87NYwYrT
NVjBJGinDA8V1ZnIFFjLtYnW/SWWp/45tkx4qI6ihmVuGGhvxdn8fwDo/SnnY5Yo
PYJ9/6+dHOiOfGjn5mKHlur3pgfEQf5Zho0iEE/Uu60THDlvl5WoCPqz2Uln2zWg
zCI8Fyqfohh3U+JFvaR3DXa1z0GuLEHnYQAQms43tz1O4fD/XPkLEfw97eXRznxA
udkUKMM4B7IVhYM3nERJJyQU4oSGCQXBDvrNk1d9MfDaJzPeRezYtRjiH02d6l/B
xXhy8qMGflWjkK9TGrhWE4kAuA8Nkh8g5tl1j3ncrsEhPpqMoKXrBlDdh5R7yV+k
db1Z0x8+xDc4vSDUtMTJNUfG86QlFtvNVlaKf9nUmCgtnsOgPwPGYt+vOaZF9ZXk
WvuOcJxpj2dCII/wKbflHlkfwDU6jsicpDJJkoyf588lqiBrtlCqmZQzRahme/yo
tBG6OFejwcRtVAxJFzJuImsjQ0QUCnCebqMDIGqFH8WDWvqg/jtm2uFpthONwaNZ
whAawa/iNdfjvCP41QEqoiboxy/rlwxRHJ7aV3yXbOpQLBS8kb1osbVyrR6/41dZ
Yuvd+VHpP0VeLSqNoX8czxfgCmhQpPM5vw6nvCa98+Qv6pTnP2WMfRlHj1eOIhDr
TbOQZJGG1FW7UBdsBiTLghXnIRCCke258FNYUJEuDoGRPMwGO6QiORPqkacL1vnf
1rd/xzTZlPvS04CZEP5dyb1LiNAc020GzcD0DUBXROxSf79xDrM3jLVaZXMUHGiN
4fzufHlKdZYODyl18WiMN8BGrnuz450PFnX6Vy2+7ya2LXuXSCo+Q38HPF8oybl2
Y/5hCrMV+bdwgUUxAC+hB6lcMQJe2cf/nFIpKGMQ8IJTEvtHSCsvRJ+WHn8e0cj1
bXBi0Do5EGJyizNnhth3aEU9bWXfItpspeVefCB7n2uVVClqfvgDi+1XJRo9brUQ
xay9dp7f14hRpUWf8ooqPqDnsnhfSNdq0ECUR2+SQX7oDJN1DghOvhqVu7PUQD9P
CANP3dEmrqQ5Qjwo+Jgymkjs8On0+yxtbPQtUs3qMEi5DPbrIVbVzvd2nVowbgAH
cpj4dPKqOPFm6KejWvYNCvaDHOYGrIDD2mwGo8aChHvUAunWy7rSyd0rwJKTF7yY
eV07zd3pR2RIhjTPiDnqTxSFj3U0bRqyFify46CqdLlRbBMmWI/73vtu8F92mTm0
okZ4vuxB7kqVBj2SCvEn2+OgqAOiWlqpRHgeR3F8y7OON38ZqNnWGtCDjY24KiZw
m7avuZtq3y1A/I2SNwf6XBIrsQOCyRWf1LQPtWj363aqx9PS4IYO86HBnyLuBE26
rvxAQmxxdxgxIIcoMQhQE3UF2KHuhZVHSReuBNyk2rVdMUUQaHtVtZkOSqtscB0V
+j5aqSWcwSC3kZfNCEMnyRnzHk0pIghXluV5Z8+3NT3nSBphiaw603jDJEIbeyb4
94CAJWmjexcq+ZCloId9Dd8Ld8jfjLa2Y7EVJxRsZrWq/R48EKzHnU17Iq22cl7k
mWuz0OWe7mEs5U5jIRXt2P+yuiWMpCS/Vs4vTudzTM9l87xOAZueQcQqgKnJn6Z3
kHjZNiyUKqsIB+cILSpbT0PvoXbmcREULeUCSo5HyTWSSBARNMKum1ZAWJD1RGLL
WmgBrRtxXWNEP64zTpx8at1GmhDDBt+gctOLgwsnn+WyHxPqu8JARvtP0yiW27U6
CUFpqaRJZJXRaPBpcgmYyvnLZ9qf8yhA3IHjnrgNV8P/tNkS2SLd5WkpcuJOz6yU
xJyHqLkoUCcXGPbrUFYihMRuGD5r/e2GJADSGTwnKuTO74/qLH0fTHb8KCHkjKdS
2FhsaL8ioTVvwtfTQdaE4KE8pZlxhhe6eX/rS1mgwZ8KhrsMH9PI4fgKqcXiSO1c
JPhSYffjQqL57u8XARnL9EhIgTBubac/uOY5dlWEGBsn6BOl3CUSYmR+sIvXr0bf
61hXb6frTOU/pROPMY8DSknQDXKN/Z9vtVLji83qxFc1AFX8p/FcwqTk8bteShkQ
27WXMgaIswtFFAkRj0w8QNvRaON9GEfm+YX2kq9QxdcDbgzTx66a8icfMo9+c/WP
0TGh0TVHeBLvxv8+j79Escs1zEGBIrKHWIFIZRLiKbcJSe6Bg37wBgmRGPK7pDnZ
xi4y28vIuOr9Qekc86Vv8fF6kWSxe6rFKa7Q4j/x5LvH05ZCpenyqAMtUIQym4KW
W/7gMNlByPSsFROb5tqR1FESOSgMzyzh4ByBiuulgim46jIzCAHZ7lFPeROQHbUl
8Mos7mLxoarHc+BNZDptONmrtDEEhsBZiqtgwxrlLJL6/bE58Pj0XdID/0hZftCQ
6p6YhsIS/MbNwBYbV5dYBSk/a+sltujvDB8mlbdZDlaPBMBQZIIshnC1AraHzU7C
Jjh2dRzzxaaUWKKItErlcdLvcw7zBHiXsFwSumaIOBK69htWFv8QR9IGsNxQoOH9
Ce4ZbUQ4k2YixcaLYMJ5Y0dnIzEVWud6H6nPHx0SOueeik51Qv5/ZdLCcOMCf/d5
J/gOyMlWpYRLHkjUr5mDTxIfgJ/X6nJKCJBzPwKibmK0wpS5+XkxkHWesbAaH9H3
Sicta5t7kaYPn5EOiSsQ4Xjg4fkseHFPNhIpc+rbNEeJJDSiNnUK7wkQ12CcqQf2
d025/LkQUkBQYtZmCqlnNRNbArz0PstkKzaiUwUkbbVfSPFZpbKSXHSUc+uv80/M
hPbUCQ9HIKO7NaXWqf4lN7quqqPfMX4xIZF0YYPoFpvo5DZ3DhEh7cDUxvL2VEhI
E/3wgI4qFrZhr6O/6uvQ1+Kun2hgVskkBXO1r/dlw+N6GqU1ldm5acFpzgdbj2Bu
jVR3HWgHU0r6R3CaeY+58s2DVFkD1GMNy2kdn7bM3jynYmZsNXnSSLVgkc+XhVyH
T66mel6nDqmelV8Oux4O7+FnHo+qGUBPszlCIUNjtxvouF4tdxkq0RWDwwuPMDPb
txXHWlXdjV/i+MaxE6b3Ut9ErgOPov4OSq4/skR3AQO1/vUTnRhdJUhM5nKNXDMp
tFyEA9uzWIsm53aMQLtovd952EiULC8sSlXTBtDyxkoTCgT3NwGXAIiOiO6c2fnk
8ruW0OSjj83+gj0OCOS5qxTvTpoqhNY3CD8H2CHMpOk2WvKFYfahU6Lak8zU78/r
b6zlbderfNdGBqBRgTVxc+ekjPNMHQgzkXD0pq3MzJE5Gs5HL6jGgoZz4GpVdDcH
ImWDbNffzETOMAs1pDB/eCvEdAF/mdHkq9rKkcT5Lr16OjShl+AgYElv1Tod6Poh
oFPtg0KP9jpkcx1dPJw0e+FEIRMRVd7a913JuVBoHSAlHbrJHLKyLYe6jRneyLUF
ft0zgyQycXstnLoeCsFyUbNVY+zTIXxZwM5Vl98vjPq26LqAd8nB3W05OA009emy
ki836bAFwsS1prqV4Jhwrt5C/XX0x5Mv+flxpljze22mgaCsZKle8jYMNUXz73oA
VMYyljU9RbP+Ryme5FokaYI7srHboTAyW2PVPo0paZtnFe2BsIXwvz24PiOS9N9l
lmJVn9c4rWeaixlhoJ9jW/hHqZJEZtkAx7XLPfW/QjsEORX4zxX5LIfmMGpc+tIe
zCdT7nQuk5+gXg9jONhZGRQ4aSSCAUwzpLT6ohV6wJEYNMyFEDi+WkIK9vfm3oGR
DmzHs0QGDxbvAVj2w1bGaEaLdLg5Ld9u5ewSR37LtuFRDycDpJxSrUsT60rgupS6
znCGq+OFhhwEzUI247YPhoGFPkzZMnKt5zRKPu4lIUuKRByoRaWhTnR+2JXJrc2h
PM0SmDqlkL/SSPmsUEt2ugqgSt6mb0+nuHHfzLnzH49vGkQQX8oHpUmosYmnZwqB
c1bByP/QrTEadtan+I3UYbuQ03UtEKCgfVhFLN1dqmC6j0a4PQE2oj4hLcHruyo/
RGvPPwQ7yG+Ap7C+SfiIO7RN23YBd/b7RZDavM1oEoYUPmYpsy0i2CIgXs9MMNDS
J9xLwarRHz3N41/MmF4tuVqTmnP45U094pBf6X3GxNfFQoPd0qKfaoklBNmh4gTt
wWXOpM7/ctj4z7uFRqxuO2Vbp2JgHrRaqBAjzeLmIWuslPK9GC1AQmqp2hqrTwFq
ts25LLwKwIuIEQeLAdCqElW5TPKNQU4BPENAJhr0KwWY2dyqZL/q68Z7nFqrXYB+
vdsglAueLOA0FVGnpQzzXnxdiPL5KSLf+7eZyxO4OM834UG1NgWe6vb8XW5FT9RO
HvWpNvVTplS2jsA5nxm3xDR547Lku15OHfYGCAnylRtEIIKvKxujhvTkMLLbY9TK
zuAK4CADHe5yWEsxPfP7J388u4QX5w5AlUUFTJdz4jGnRg5ZxBAG+Wk8Gv8VUyCu
TdPYySkxmAWtjR7hIReIUgSeAOMfpHaJSV4FbHUX125tNFK7Ft7A4+ryUAAK3is+
w8EMmpE8jX1ZSNPBvUxYehR2yZjy8w4eQXPiOnwFVareSZrzy1jfDdbv1TV470dU
/BnDIVGjQmmgrn3UpTjDGJ4X5l+219P75QwcRqJrMEHVXAgXjmTA6hc1+dthv2m4
uNdJoEyRX/eHRqqt5pw/Hs568hgfoAzCnIMkKQdpFbWHAWzsfs88pFw4GWuR4D2N
KZeyzYYLYTR6VJUP3xl4xZABI9pWxiKwHIDxg7/Qb9wCUumNd9zk2bOYWbmdX0fc
h0j+KIeR+jRRPYAIVV65KkqOm8bciK2QrSlGa7xs3pDH0sPtlL1eb0gchLg537sa
zLwzoXtHRn2BoBE6nGzyr1RsAMvAymfn3ic5mwqJVIu/VasQFJO2GGUkg6v0Qhrw
LY+o6M+WHexqum+L8wUwQLcal+kZJaBxC25ie/5XdYDzRt5F0bbyemG5FnhzpvQz
FTiFqht4v/mnve79H2YvB2tamgc9nH3V54xaeQURv/A7B1un2qBV2ZnpXemZRFCa
WL/Aeao/9P/mJ6ZzHFTXrnWow5Uq59gPbHGvdsZQz++GwbfILBzQ1N3cTo+3hZi2
DU5mp4uvXbG5pIEzclkYV7fp6yekjBWWS83jmQ9C7R0yuY3AGIqKzH2m+LhpFIky
hjm3AAQ5uMGmCHNsVYuPG06ah8Bcl6Z3Nl3CZ4qtvI1s5a5iKTrmggKwzSBPX7L6
217Yam9pXBtT8ohTAdKPCPT3vuZgG/Bf5XG7HeILIko4wd76sWL82BB3m31qsB4X
oilP3lnfJFRaC/T+NxUXxHShYtPFmFbDQ/XXE8QIJsqgei5S4ubFVbgDq5JZW7Ir
/yCzl5BHbCt9XmnKSWc+pkX/75X84wZfcWRgFlAcV34Ol8vdrgZIZAqxXo6VMjfl
CbNRXOnt/oB5k7Igc8JpTws2NFEcJK9XDEoMBjD9uOERU54wKOwyBhuOGzSPpDAs
Qj7JN4mNDw8OTmyIfxmUDpz+0mKqspn9m/p5kxMaH9WX+YWxZ0CXFyhI4GzxTzeX
ZZZjlkKfQtKRQPFUNuRGJuZzcTDNxi8iD30zGpah/UGz9UassaweqFNIWhoyB4uX
rykup+Ad6AUaaCOySat1Ff4a2uQuregezW51tKb7DFxPMxx/qLH1cACaePuywj4t
5TywQpRlqUBQl4xkMHWuZN5Kv0qWaCxN7Af7Fi1/SEw00UtFu9rfiYJAXVq4AoPH
53RU7Sf9SUkekIubNdNL9/IRjXaMq9HpiEpug/DiOMbRbYzxFVB3Swpg5152txDx
3IPI5wb1UKpwqH9wHUQqSD93DnhJsMsu4IyFtToI8A6AZCfvwHzkza8nTw3wP4UF
oTyrLXhwY6LjqoA8NS9Hj01Tz5ie10yFX3jlB3ceNzCdq10YWevZwEgksS+jw5tT
ait7XgXffQMy5yFKuKn/TCqcMOkzHDdEsKo0TCRMY7QtZFVJik9GdhYLrxzaf7IH
ZGynoWxtH6INtlQH3IWokJNyGLs3cR9pOu5rKFIPdIJLMh+7YEn6yCHA8tYJnJOh
qCnjbbHIdby3QWADOg2LOnnaN8hJkStU2O+bdGPR/fT4aCndvoUnCfXlq6aVhosC
VYo+yWHQZ2N6KD7avnuNqcKoYO7FyiSNRgEFoOQBBQHyE3tH9mTg3GUJ64zQDlWk
AthOCSVdM22dF/pJnDVJbdAeanccWQ3KV4QVsduz67ya/gF9AUCDt7JmLlOEfw0U
wVkTJvOd86cDNgQSZDv0ipS+GgxzWWrvH5ksP7utQFjuRBVcTqB5JLxxr4bZqBLb
775AyvMd3C/33Uj9IBDjUxKRZoDksfunoxZdewnKQNTTaXWcHDdcmdqkx0Sqmo2v
ZBbnAhoQoIizBUJdNP/82g6WEqcNPwEPT3Z7LP0Tx889Bozji/luz0PurR8vZglH
bIAc946+c77DFpBfOvz7JW9Q7PRqxl1YP+2r9Mu8umbpHX7eKNFdCf9yd8E98RxA
qCnbpZdudsU4BEr3lMyHfFEw3mzKLwKBUuhVOIen7QKL0Xw4knFQnps6LmE/7P0m
5Fr66k6yH2hO1kf+HQv/xOptCUt+bi0ZKGnLKoLcyclOu5c7Qyr2z0KDw8XAygvv
mdsURKlObN6eecNoB4mOhUB4aUrHDcc1hM9Vl5I1k3vlF81WdyXYV8XCXRVKE+BP
cAXe1CfQ8MuUDbjBmXcaMEPhs6NYBwG9wtPcazIvM33jm3FHjp94RLiJNVrWA3uw
RfwngltkVDNHG3uq1t1fmBHEqzUnVq8HT+oZtauEzT3RJaep3JuaLHnW9PbNByEW
Etr7CFEl7MWEHpBDrIBTV7CkSUANVMivFFrT3fiP9sYaDmdyAWRUi/ru1OKiAxGs
VCViOj/TEZ591T5vVtwaI1vfZIO6+MamI+/qO+P60R5iEK3wzyScJD2fuALbE10K
iAHNJfWyPWbhW+/r6n64OPOu25WAKNbYaAQ4GTJ78QmEkC1+kcvl+RFzX+HUgE1M
XTOV7UJZq/KmWMeeNJv8GfP2EnGxGEGLlzblYKR4TIWn5NnjPB47zKwdZpf3T8dq
axop22rRhwTcnFvMFi5tXXxbOa7zcj39KJcb3++pfMk3MifVIb3aP+R5zfS3D2Xf
zlRJ09AffxxYvBFFtwNK0JjIe/NF3+Fcxris+QFyHjAirhjd3O5bhZLIF7A+KkfD
ZqrnRh8F7nOS2fcpi/ByQ35IvxGAETrNewG8C+nqeVeuCxqlHeBN4d/Ob2Owpgq7
aOmZy+8ktv/dwR5btTAVjkLfEdGYBrGqxHB7yMlfFM4/uAATznJhwkmx1N4Dq1ep
5tcx6Xia+8UolK/gQw0vo1TslaMoSzgwNt/wsQqD8VK6d+Fw4LP/dACfA2mKi81m
C7tIHq8kdvBjpsfEW2aykCqUEtaaQUJ5j96LyMUMWpi5c5cTS1OT2Xpin/z1Iduy
U3LK0U+sirU/RWjHB69+np/YPweFpsS+yoqSysCiMhlISVBJipeU0/hHn9uGfMXw
g39bYsyVc+U5DPa3g2W5kz9gJKMX+bOvp39CYK6za97F82MGqdaWcI0l2x1kEgqJ
wsbe/cfstGresqFNQ118v3plNfqlBsS/YWcgPLPn6UESFd4KlPnfIM5W/kWryWbE
ZZpeOhF3pFSKojqhlHLNqyYKzSa/kqpzqTLc4toxNVVUq+5gGcBUU7DxF87nwOw6
pYM90XjdMbitwQ0PdVnAOZw3wtPF8HttUjtSd/1xb846RmPfYgQmOI/W9Cpy5lkL
8Vs7L3r9h0XR//LQndk3suxiIOYmX3Rysb1CkUrATdKz6YCdaB5hzqJLcxMCmDXx
ans1AJjoPgNB6UWPIMnuzDJAIJLGzM4VpfjUqQJOTn2XNfKvhh5qlZN+Q0l2jrKh
z5uDZd0SfSQ7fz+foqOCacRE8jaNPWiIPtEUrRbgVR1bEqXzICJ5uKHVdb0zltht
Qf1QeOkSGrMa+FkmEOTm0rQQqnLrMlUeQOZ+OZBTfBiytEHMNpQdGLGyEXrwtWml
3+lQIGTtPS8xMz13LM9dZs0Lq8khXgNJIX7Dt30HDjz1CuW7ViECO5aa5oDlrcTv
j/CljAqLafuAH7Ud64rzUA94BMKK2bl+2HiWmM0c395/bNhs0RqHeI2y2syfs6+7
IOpJTbJezWTF6wWI0MVmjEsjMttfiYpobIrtEGOzcMLUbGK/q/dM7doXNrKyuSs+
Gsb3G8J+fbFXGIPIG5C68S7ZDUpNJSm2IqIT4glwQ/fibKMInzgOyZOuVLn2lPyy
OhP94tIFOYl47qct+CeqlTo5wJsX6gn1JKGNdNq9ZluJfb8ei/3wdn+jjaDB213f
6uaoaieeF7bYaHHrRyPcJ4HcCudfymjh8gXIlX975g7zFS/n7d1xQ6R6ybqWyHrw
C81+0+CWqFgPGuUtdmlAF8kPSZNQOri3WMq6rEOvdIvDNLH9xQPYThDssfPBDtGN
r1l7xuClSCGq1YZzJXEmy09NWALh0LQMni3z8zacJXAl50WAnL8vo2ssUf4rSMBk
mq6yMZpfkgxOFD6q3OcIJpTHafrJ69AMd5T7xnMphU3te84rvM3qaXdyMHHhzPwK
rwatSIFN4hOPSmwA1P8Ex+CP7BQcicJqCGa5DTAo8KwuD9C+Sk3KzbgqwiKKsyE1
y8fMeFQ/qWfG4Zb/OjxrpN91iSpW2u+ORvRxjBjUcWNeHWKTBYVezO1CdQ8iJjAi
aoPK/vsfzBq2UeNMDCWPo8zZCjfaa2YMEBMt+XuAjCrajqIuzRstJHdK9HfRScYJ
nUlwxfsldAG2u7pVEUTszLrvT8PeSEwfTWGen0tXxCZrfDPR2w9uBytD1nUUfgfj
1rkhKBFD0Kx1pfi/gmxaD4U6LcKhwgDaPih5wTLkIj4uxYEAqZr34S8onhAFmCfS
0ZfCRLFnHsLNxDA0EYu3gdis1GVqCGLKXi+XRZGJoknJWrMn8cisfwLh3b1X8cHD
y50yEfoTxohvdxxQqLcvjYceMDICUW0hYlXLdIpwhkYjT9FqsQz+liv0pF+Y9hWL
O5JPUQunWXR73QXfIPiivXzEBMNJEg9m1xOGB9aswFi5E2xg+4LjwpcTmMRD2TiG
1arC3G+TccOmrO+7JBoXK/PgUz1SJqQx/dqZx5039PZCC4azW1r58qb+IWEZeLuX
w9HzQ0qMX9/i8kltCew9Lr1h4xbCM1pveOVQP4kzW5/TMWjnStTVokJSaLuMZTHm
g3ToNmh1qxGAtCLrZwmNrgV3Q4x26hkknpesFiyocJ3UX7Bo/Y7Glq0zpDsgRf+t
lIIgL3tothMeUu1vJjQSZYeuVX4+2bR87bTD9BdY01siFXtBWsno6fAWpUKeshl/
9T5+7aci5a1TIgyoDgYeO4LtZqTzbtpTUmnDvapJHBdCVLICGsVkPbd/DKgBje39
+A7hlr45l3kMSGVqoEPEbjNJdu9Ad8M55y/+urrFp/LicUq4Vu8Rq8pcqpqqXTng
t1jKi/6SA4WG8bdRGasnTaL0YtkCWiEuOmoj1TXgf+8I6lYxx9HnVdsWhzJAVinW
O27rRSYwQAD3YDYPU9pIbkM8+w0PYUagmQ3hArcsWuie2wN+DdvMoMqKdgsQ+aSG
KzsubpJqNHk39kbcMf96nSbeD3/VZBdGkvJm1piyAhsI4HliyjE2rjksS+J7fbMY
ykoN7XOpeGSy7RItbs1sx44jFJKncuCnl4AOeEYlmYIgJjsEjTYUIoAqUK4uS24g
vJROx5CHho8Y/m1w9ok1OBUI5dg83mX2dd3EMtYWk0nAlPnYCeArPUgGypU5v6Xt
1ggN3Bp4NFHEoeQTU9hjG0HK/Jgd+NlQKT/GMzVAq1/v5u/IuxuigvUpg105nd+U
9/f4KfzQCUoALAy+efO19XtA4gVb3iSl6ZrkMB3qYWMnOX/o19ked6VaAJgir9zg
s2x7xjv+kIE1XEpiSBBGKWfeMLecoo8m+7zJiNFsdC2A25hgW+sMut2Pr9GR4Ov7
Md5TFSddcf0r32PeWB+QrQFwiBgHLD/MrObowa6JaMao7AK3qDg/oJTlqQ/DQ6Oa
lN+uFqSnuP6qZHoLjETNNnimH5Fc4CDoebJil3sy9mQcFpO9VmwQQPCLusfGx0zm
ZPObv+HCJ1HgWZQRXDB9cdKR9tSSnfNOonX4rTc8hN8eQ6TPQ19aGsSLi6HM3w9b
M6l3y8omv2DWUJ/+ZYtg+sRr2igyzMTQq+N7sDAtk1HX+aex91OWoBtrMOgJloCX
2VeOIwh91sMJ2U02DUSAA1c3DnaCxvcaRq4aI8dDzrANI9rQDmqmfCXbhooyz4Qr
6mOLsV6L5/RECuz8M3IfhbLrBSaHNIIVuJ4/eX/VJyMtLJKjMCGKbwmf7uGw3SnQ
iew/Ut5ALsEwoUnJnPf6c8ZuRqPcRFzE/wUEotldCvRO4tKa09lc6F4pPzEI+vqq
fjlnUYdzuf1vLki9fBLsWCLvR+t8qy2h6p31qZKuayWLmHIgdMSPkUjvt2dW2Ts8
Vc09YrsESzTYpnuVAcy4Qo4+aUF6WZE+teqQu5l9KAsaFtqKe5PTPQbU30X4MK9u
5cLPZMyey83A44VtD5tuMzJiQgDy5XPIbj7Ie3QdQmoYZFNudEyzEFVO/Da33STe
e3petOlgNqpa3LP2FpFKaLP9mFZ2c/G2e6nqWsTSR0E2Ry83sX/g8FlV0koi8cA4
Aj8r7DnU1LZmV3g22YF//mZlEgyPxwUjMViW3iW3j2JTFxTaWeZ6Voa5/xTle6xP
TVOglgUwxp858/gvvvaN3t0piwQ/jE2rA6HSJqwxF+H/k4UCKsrD4MDllJ7A01lS
Kpi0M2z7gCqx0LqHlN8QTgkuTPYgyAQIOG9MzqQr2b1xjVtM82u9+zbbyVJtx5bD
BLYwg3iOoCnBRsKtH7eQY/oftqnJauucQjbPQ9GbvZgL/PWfddiNFG1vHSyuN71D
wjNDG0Yfd5YsV/pKD5vNxAhKKsh1yaV4Ibiz2yx/vA5cZppMNew2BTC1khGOdf1G
lTUt/jlz46VBkfmP3/Nv4qYaeEj/F2wP8aygRMhMMPtyBlXj+rnV4ncmFv1MOMqv
d7w07fOJktyJ/iWdyk6hNrgcBWR8echxR6TYfrMQhoN55hb0ig3uPr9SGTUdytRS
+NkDLEwesoLAYR7GunmvZa+8SnSWW0oPM/ewtUsLZXYTKRAjfmphxU8EhvB8o37Q
G+gCjCVuqs4m4R1HkLhEDAzMm2r5EdVP+tPa1vEcgPxOaLwBQMDb7b2kG397hdKu
2DEfp+2UChVPBpvujiY/uGqBoOiYeKvcSHyqKmMC6uurRNoVpJx2SVdR87Ccqb0N
0lDeHNGh405iIo4bU0m/j7zI8AKLOGhNKqmyHGMfJe4sNSzZYV22ePP2NHf8l/YR
xAvIGS9WxmT4mBRdMgcTapiRBNShPfSXuPfpq8LOA41uuaOu0dbNQO2nGoOdeemW
7/XO/YLKBqq4Y+XEOi9C4a4+NM9Ev9f9ysLAPvTQWIi/bqwS51PyjxvLWdX0q0/B
b+jp5Ewpb9cGkK/eIPs8f9VSiPcvnNsPxYynTNZctbtnuaHiqtROeVsL2KnJ6H8K
8X+mQtmcQWgWNvq9a9DAXO9Qvj4nys7dKvi8bGgIztbtV0G0rS2zBgyBzgtU7PiW
R00D4B+5rc9pwYkkmRZjOfA5yqO/VowOBCWJXAxrM4TROF70EPLm+cigFzOqg8z4
0RsL3kYp6IIfvClNl7+BAY3ELc+lj++JHM5pE0b2TxOqxm1rxoPbfTH5oyXQeh6q
qwO1UUPxfH/hNY21fgeqQQUd50Suky6agtQXmtoZovm70HzlrmZTFWbZuoDSY/A9
2WK4vhBJHU1JrSt+E0+QjNeIre3WkjZBZMdzp6atK97m0t2BHS5j+3q8ec8NxboO
geBCetFC/yjwVwmmTQC5OMuamDJOVzubcX7fFdyfL4BU2qD5ibPbvnk905xtSVwx
uTqwpnwsaqyML396KZUJ5qt3Gg/NmwKTtUpXRl0idK7X49tvNfzTojmoJETFUWIi
AL76AR3cu56P1gNDVU2aiF2qqQ7us+z0OoBkhX3O/2yu7+BAJX8NaBARh8+Y53Jg
EQuo46BttD8OgM2OlbUxRbrAH3ZY9HwzVR4H/VMo2Bjg1wMYBq0YMvuvLR9gM74i
6R9ZbHHEoOjPwQKjA7Hfj6eLEg4lz7XMsyzT6K0FgDd0mC9K/D60vzlgvc2o/mcS
iyGTsk3bczmCv0GUYNo3aiyUBaDnYJUFQoTf+oYLiadnXcSYJY1xYNnp9lbR8zWR
JAPne8Kz2+VCaDJPXD2hTh4rfQmhdSNS8lF3FpffUagIRq1qR5sihHJVGHYqmiZa
qPufQgtkjxxOmwvcj2bMt1PHLkiMoFfEL4r9Tfd699f2ierOeIgohytVRChB9EGy
Wpc3rBRxf2bBd3IHLlHeP+HzBV34Wx6gM7d3ZM4AoxKgPL8trg1ABlknAfXG0rWp
UFQh64nEHCowpDuQmdGT34xaXXxVcMOplHRu4PFncGkSU+Wd2J4mikY2DzXzDhIE
JUHQst6yOcGfSi3R5vioYXCYRYQodYdzDmUzcBTROfSEUh2KA/GfC1cUzYQ4Ogaw
sh9RMzwQ7LcpXtjIBR27s13qSBhbGSbjun2iov/gwy8/LKGvCV+A8vHY/C436G/c
Uug5KAQwM07+1ZyL7ybLSDVLN71Di/hiBj7s445XdWtSIxM2bdSWw8JNx/AymS8U
tlpLMOvIqUvhQ/Q6fu47Jn8OnmmI76F1FUMRjl8jyppeHs1aUy3TTBe3cHFmWQW5
Ed5sd/UWMmBrqUjDoPkDnGRWk3+tomn7lo41/VhC461hPQ/3a9r+wHzdyxFdtfK7
u7DlsDy/SWW8ZCl+W7OO1q7E4uxo0pNrR1Jn9g1fWhbRv4/wgCIK/7TOn1xJ4Wky
o8W8qIdc/dI18eDnOyUlYI63k4t7adv3sCoTkogJ8qeGHk1kOficaqNSwlHB5QUU
0d0TrJx4/nDCyRp6HSzmIRpwhCdDJdKJBvGsXny6ShicGY+c5F+pP1QztkbF5NcS
9ntttpFupB5/ppL7L6NqGaZZ4+Kt39BylbvrsIqOaZC4XFQHFxdwOYwLA8wR9/BK
egeAwONl7sTzyhbgYRS/E2ZfTuPuMi0mOEO6SABm1OpX96BnD30iG4bQwrOSb3a0
/rZrf576jhMwFx0C0YJNB+9chFUUZWrPLfuNGqiOdU5jsFi6qrNWoIyj9ebW6gYB
I7JMmeRyDDQTvbi8olxt3XtCa+sHbTPIS874xfZgNbN64IgOv4P0+z0i185khTq4
DKYsJ0BbelcYcdeK5cKbBGILdZVKrVTZF/ZYbaQn1JKRKVnoxIA2fQYizNKbW+Xb
rzkFB1iSBgtPIcByiR10D4NqQbRGYoZmzHJ5AqQ5Jfx+h/hNzrkuihkaQXuFIgdd
O3ntbHootUxXX9oQlhhgAqXGxGDj6t/Bw6pfxzzdtXqtEPkKYuTw/deJZyhg3UjI
JOfLXMtCKOe7vKVTmlKcpO5lVxQCTTTQomrVBtA1Jcohp207lG4nbYeT4cAEXIhF
w6Z31WfnBbyUcW6phspEwDONvX6qQF2A2iBciMjceLw/fO46151gZ8vxu9OvlaJy
YKqrx7CE+qKgzARUNRtUaBG4b1mCrFATN53BYlNyaVwOfit4EIaj4xxWXaBHSwsI
tJU1c70WQ/QUun4kZBw133wqcoM0FHVWss4YUqZQYxO1a+IGM50UnYXFWKIn4ikI
9cf0wcrsyQXd3y8OdpV/zQhjEn2XmvYBMgYDtvfiLehf89dgKN+PumNBcT+WA8bW
2XmHDlbzdYBLyXPGtHPvXoG9xJ6kjyFL/J/pDfbZvGhSJjljtsC412RhHruu6cpd
iVJOuxVx24szOZf+4O1rlHUjSNmVc5njUhxqMkwoJIda3J+aY9s2PfN8w/YbJ4ms
7sJ4PttVqNnLErk3VqUzeU+mMAscauUZ/qRfwq4kfiXUDwA+fgDq7k2CpZ+FMWRY
xPbWayHSraX7RR28D8w1ARxXlNsX6ja8aQAWoJeYUNcLM+ly1ipUpmXyx3VXt4AQ
n/puVKZdtIU9kYsy8qm1BPwnOOSuGhUGVwQOXXaZgWrlKz9X7ZXjvn6f6Lb0VYAN
T3GTmB63wVDN442AUdZeoeUGzPLzf2rkXvkGqjmEA1ujqJ7nqG+16lXgndh+pfXC
tCxZF5WtW7l+7Vdw6604qeBCPRm5nyfn6RiJ5l8ctERp8RlVSY4wg2HWRtpsc5A8
EF60icajzyciixYpe+xTsGRao3Z4neHlTQCrX7xRXYqh5Zamkcn18NLa/cTEi3F8
Z54gJF9FDbS/4b5bJNCkTRRwXQlUp1oYuGntnRJvmM14jwuUQNk+0MDG/9ZkUIpA
x03rykkDgGWptpjrGVWWFkATKm7BPSsdj8avTs28bc5OK9AgM8k73CrZ4iT9o6jA
kd2+btyWu/GYCo2bAG+QUtqCBjopI0giuZqFyTonTxUS9wK03++3xXe7hqtfR0GP
oDyiTyVCO4Z+p+fOSAsY9cAQwpDr+jCTexUzRF0/plXY2BIkfaJeNIu+F/3h6xMZ
EjbEDmWx6IZ1zrVCA07Rs1Z/GDDdFpOzddkXRAhOHDIWGb44Mi5LmOwBZ7DLfKI6
wTlugcOdJNGqAB0qRI4sFbXDfSN8qR1XAuisiCMyTVakbHYmUqGAOLdVVNQqtjHv
ks6BkWO6M9NVExquXXG12in+nNiiSbFw3JW2sdmMpNT4LP4OGXViV/Tw4vdOjO/X
Zn2oG4/l+Y94Aasked1MwJZ/d2MhyDCleA+6pLH0Q205hejpbXqFYL9IKOhVF7Rl
fHfOB4TQivqwrCY7pWUNYs9zXhtiKPlk5/pt3i9hEabrYq4qnzUM7l1+dCO2jt8u
XdFCqUf3rJANEmIO9G/aBEKoD5Sy5zge43igyG2V5TF9atCtS8KpEbonlMJRqUGG
9CEm1QDTZa8J2dd9e2jWqaGI5BHUhc2z1TrkpRQwoUuJ071F3gDAK+xiS6aJ1Bnr
y9yGhrfjeU4fRZEspRBOU3jRW+hR4pLgimKbTp6vC9ERqX31/6Ok9jMjbCy7mtFZ
FvjmR2CG/dnFOaN+VETVSPYqJxtr+dP9cZ+0FfXtvH8k6on2RtrT8m7k1zppMH2b
7sAo5bvf0rA8aRtzavFbBRKMMpSpNIPiXce7mLOx7aNN79Vs/yBrApd78VeOTM6q
JL3VvsSDYzYsIfDEBR27iv11LJgqINT76o2gXisJiIT3ATv6D869TO6JOtrlUksq
E6UwZCA1CQo+3tx1Jufah12T6L50hrwBAKduGnvJ5qiXeN4fuyav+5+OtpOMfVu/
cfWEEytvos37km0OPgnlJmVkDbddmH+/xNEbQbrizyNW4O1woyfyO+g2rSoUz+4G
BwGCuHDB5WHW+WY4CrccoZSb9k86olODnxT2RmdFnr7iffNQsE1I4unrAJRkRUkU
0wm2CGrWqmXRIBOtMhDwFCXAKvj5KpVBUQ5QAXkjbghnoEf82dyUfud7NP9TFLXE
yWnYUmXHnSkwMURcfE8RjDGhvmsM2cC/dD1zLmvz6o2lgaaNXxZ23x5jvt4EZTR+
s0CrV/iju3eMSw6YbCn9vq1cPyKDivMYPS6HOKLOvtjExPhyEixhGIDKygpiacVW
Mnwj9a26UkmWer2IZvnBrpRokQ6LMn3Sh/x1WptIGM7N2wq7GhrQoNg39cliOg+p
MYmyqVAoLEGyrL1+IuchvXNLXQvyvkbV22dWFQ0J+LzLaHiHKPQndChrmPNIv5ET
L9HOJadtnsha+OqgHLlOjAKJ8OmCjLs82ZZOS56V7S1jxMRvOvXpne6XxVgPohCl
kPHKxq5EfdpiUcte9uOvaKLu1Soj+8w5G4A+RsHM7SoqRy5bXbAuWvW21dn9U8yp
rjbTrS/LMSyDjGIFFyTZFRAk2JLRcSRtPZs/YUuKL2le0I3avqW84XdoFHLNnA7p
sBXdYAeoZjTNc8EY1KofFE4/zHOA/RvYJEELB7v2WjeGVjibYzflMCRIzguWCS8D
dUDtfadnjWTWzafraZmPcGpL3G1DD3eCAW79OhNDTNDTMyOluipXJK3WHVVmguFu
oDFemSPTGj9Wlq2lBgclhp71n8HLG/TvqQMlLUwG3KVLis9K1dk8lBnnDuOca8pH
AnUOwDPlp4lHVmNm3YwWIy0sQD9Afz+XxAVLxVVncOfV4gxbe9Mki8TC36FzgZc2
tkLOb8+uSYLfTBA+OErOxIWjWm7C0IPc95NeyVEhELoW6ZVRN6sj9UAa/3laDWXq
zI8guKAyYTF5UUNa2eSSPeoEjyNouR9iZjTEewU7LSHmbAUQJej3tdxs7UwbL6ao
VU5QD8Xn6ChRQMNZCrTir/oK0h5pqfqShl61SYwGe3xcYYIEjURkV6GwE0UrhqHR
hfkh9oPwZi+1XZPwL+3Yd1FwwLknmiPjHdq2dv0YT+yuZ/zHuoxKxf2f29txwFIH
NPq/Qy3bBKY1wquxZclmUsgApj9o0baCw3FBdmT2ZAyN9/1khUsjtBIXYV1bi2xt
/YEJjsG/mmdWwNureJ200RI7YnOWhwJ5Zq5YbIPdOAyoQ1T9GEnR5n5kTDoxl69H
BNOR1HqTgeUE0cnxcXes8Kb7FaRC0tegM3PGYUtndaJUqdIDUL+OqtodvBEduyCb
tAlBYOfltQDwJsyf9eSvAq7z/WMs/VOfAy9DfdEAtgjNeWXDraggLTk4nUeo+XDu
Sx4OYmNbNtf8gIJsLT9uav7e4FlFP+98Li7N26YrdS48PL9N/CiE05Oo5OjrhW9g
YZCbUAHQMFjlxM2GRmEA+6RBlcwjV8YGhKZ/yEYBpR6+HXoNc2tqvKPlHwsyU3f2
MjruIjJ/Mq6J2YhH3kMaCXT5Zt1wbnM+Uwa5IyQQh+kXVviCOYju//f37uXuhOjs
tZRsW56N9vvnoBMgOjBnC6MfXXKvk7iaxCalb3CVioNInmKeGd45amJxrdq298yx
HRXZQlvSJwq3oMzqY5l7d3zeQHRkqS+EYL2xamkQrrW+5iRTy8NrGT7wR2AOiImk
C5SKvcD1Dtuu72Dh/jQdWIKeKyQVJ5S72lEvNMbJZvMrtNVp5WqXNBlLOTnbHj1d
dlyX37P2pn3V5SJUrLifeK+H148BMJUCpEVr1k2jE+un9axSkJ8F16unxrtYW4L3
aBEJ6nuri0lxG69Js9oyzDmMPUjyCuBuYw6MsOQoznmpwgfRTCbBa4MFe4ZQDb/D
qc2VRmJ58Dbp/TCfpO1U+LtFL5FJAtbYpfhFtAvRgRrAM3Qkzqjbl2tzs4T/AlIF
ODR4gipSl0s5rjP9M683RCbuFjjyFz2EDS/Df5eECsmpguCkv1Q+JBkJ/2PBD+I+
GFnOr7+Zr46UwCufmStwZ0zSiKr/xC7AW4lVrfi1Ina+yh7Gej1ZEuK/D+p6XolD
kV5R8dfIExzvSLnMFSRfKXQF9rwL4JagoO33CrdjgK8QBnq5rt3Lis7HowbH/V/U
X+6/N8Vad4tSew5AZ32zD9wXD+Y6kOhsfu6Ue0RvKdwfJqqweKUCC+ACGCEAaXbK
8E5Qp5NrsD2BIgvpj9DCrqWjG/IHNJDF2oUe/5pv4Jd8E4EK46Xfd47zEYVj+vnP
vu0Fv1hii4fnQjSZDxdxLdJGUpiDfKiRjiMozJSrkZowUMpj8DEUew4lDQDLpNO6
IiLtPV1IQ2Qqj0x1gN4efcHxrRN3omYF1nxPYhiM6DxWzONJhKD7OWmEJG851+ti
3TFQoqXwLiPPqR4I1okwbM1Rn/YunPiEFAvXz7aA+XmCnHrTfGz6nzFE3XvIDWee
wc+houRABAjYHnQWU8gLtFzV+nfbANXzLVog3HJCFya3tT9effcFGGwEyqx4Fgoy
Owa23XFCfXID1Mg64jQIKtidX39xddcfruIROf7tMoocij/6s0osrg/9YJdwowqO
mX5wOhzOOofcbOFHmkIwNLwZAB3p58nzGcs9SKP8Fs0xHaQ1rcz/F9zx7zckz9pw
9ibIGldz8aaSoaLFo1FHnGBeRH5xf+a2FhESOaMtM/8EQwpege1uDFdAmsOcn5Dq
lySuE1eldwsEfVGRpm7LOMJy4l3F6dhq/vb97P4nMQTeA2/NspgrxVV5xNnH9ilB
Ckv2wk2LmFOfca2V4n967R0D/lr6LibOQiOIIhFhlUuKzmKX35ilDeqP8u3qC3aX
cOrGVt3iFZPu1TGwsMi43bzgjp7uX1s0FKu3jotdqabrD0szaX/7VMPhA9U6PUbn
etXCeEP12yOlnGsTG3Y4LGbeLQSHb0su1UWO7f55A/wFN2LHzgFy5K9hM4T2Jg15
2qfo1MhCy4JXCpntAHiME9CIjIpgl2VeuGu7w6WtC6hqa4EmAKGfW34NouJ1x55c
Az6MDGr7cyhSExQq1PDgaCCq8wmfH2rDbx7nNJZhiFA78vFfzUBhqWNxWwmo8+55
NUO8NOWZZAwwh9MQK86itBmLO3V/nhQTmZcJYeEvOHaFodsiA5NRkNSKS2/9h3mW
sJigsFBDJfncS+sl+CFR+z1ZOc4IuqZBxxbi0CjXqoDv0oLaZzWBh0Ifa/TzSpaH
Led7wdvnvLlqngyShTKZxPMzSXon1ZLl6TPuOBDyvg4mLYlj9paEFXgd29U7YSBH
zGjPCXu1HHhVG97Os+l/aKj5Gsd29Iz7oqgzsQHuOEcKZdfgpD+1HghUD+zp3TcY
GCBNsVSUF6EPci9eip6JH0QbDy9TgxcT3a4rS43E/5+4tJmhRjKfbWMEBbjNEh32
KVI1tdE49Dly3BdYB3bkPZ6eg4gIYOdQaVysEr7vQ5ru0EDRXaF0Foen7asPPk51
RjgSPoFLDo7UgKiOq/c7UHg6nsv1NfPZRblPOEAOq5rDXgBrKI4rswQJi87Hxew+
2ALZS4ZeFuPPPE+sGYVQv+eQf37lOzSdWgMIbhwGKtMIbx8RJHP+wdNpGoq9+AnY
Od0t2oCY68+2VOxvaawsDG1TCKUp1g+3o6NSLRvT+r8fgxtxsqeHhzU8w+HasN9J
e1P68NIqAX6zk/HRtQXXS/8FL7k7KbSiPmkPxlIrlqBijKf0dKXYmZtqX8E+a/AF
0zLrNtNPY9p2dSIvEozy4wCndEg4Hx82f7smxsnlO/q04/+Heh3+b8zptOmK/4SZ
H2PZz0JekgcCSPXjoUCEl04PK2fKI1tM+E7ZnUXyBHwbfAUlnFRo4ZeaDkKWV14A
NcaSMMKZ44tZ8jU9jgztlfn001ngr4SJu8f9Fwn4IDKt0XWara80vsxQfPNGKJNc
5hgZ9qcURbZTd74JdvwBG3Zs/BS5JUN1B7Wwt2ETtvDncPVeFLpJ9YbMzCIzjCxv
1z8dxj5M8BP3B2OE7JXfFGgoDw5TBNrptj7pD6AEJrR5cikDVLR/tQt5x9leoaS5
J0QCLvlK0EdtykuCmRJf8UFrXOvWJz4nb2KZ6XuVhqN3PbWseSiykkXsCK4fPYdx
/VWlrHXeMxM0VKc1w/ftbnMMKaihHqgdGl6+v/AOHkr9/sKBOJPW2Xf1UqjlgFJd
kiM46zmgh91RM52+AfNNvy7Tkj3Pg8cAYP4I6mhK6cArQEPsQF44A3jAfFUuqb9p
kcl9DTfoa4X4rQnBP+41yxg5UEco2V0vthgd9LPg1L82ixpYli3ZtocYR1rrDqGD
/JBkmpiRRAZQ209w22Y4P3vgWO5xwjSkY7984rvaUd9C5+0QiCHUcOQ6tL+JCJ1C
PG8bUWWYoDGDoiuec4Y3GPYrdLkyWEpTk50XtrNj6E2Zcv5ylYmreYKkaHXd/OYw
1XrR0TXlnQZ2miESFM/8WO+6InD2YSlSkRdCnqNuHbAjW55FhNBYI2Iu3YLb7Ur3
8lTq8FXlDpu2Bu+FTWnj+GzfdVatCgkD0UG3H2uy2fh4ClIBvCNzf1LUMdR4jIbt
W40LotTv2R/kIR/a4PwiFSLM3oypAla54Dhndg8cC13A/GHYIcrVmVERIfyI7hy2
pF0wmfLqmHvl8HKED81ff47BSJXFui/DwKa2fmJXql8YJD7Te3A5zO32HEUzUDD4
YH3qRJuPoBsL4f0rbRf7TkfG9knrrYTApQaBfXsIk8X0wPrkC76ISHj4sVv4Tx4e
FkuIb4nt7IMPJBpB2nkxEkdacHQvJZBrSR5k0zsWhSQ1JC94rfXs+Uop2kLY1xDv
1KoAMm8i75usZpqfOdMU/J9FUOpx9c6qkv4k9YdqG5c9+hznTMJysbznW4MmWz1G
nY+yOmLWxJ37naBboxlNS/yaC5BgPcr3HZED2FYbu5lu4uoHUT56D2OCwCOsju/4
IyAU3s9/V3eUles0mscER6cCJQmVGDEfc2lCyMonIwK/cktRKuv6a9w8/dmjlHBg
2lg5JLPpH9/m2s5TCaRsssKerum2y7iFJ/5FLnjECS3XlvJFyXnlu8a+PC5ztDf2
x/C3rcffhzrjKIYC06GLmh9z3idtw+p5HuBhWqj1Pk0O53H+dPyMkKTDFTv767xy
z+BTepIUornndhAQlEaX4DjWLaiTjBCppY8PfzuyrpR34RGPKAZQivZ4Dl220WZy
zuTn6WiY8PZPzJKccc0+OwXExWKSuYq/LqANIB0fXT2X0ZrZRHAJ0lj/7kL68QPA
9M2SwPlwARRSikeLMDDS4uHos3cO4aaMTpc4CGGNaXgTE2gjvvzv9WgORhEo9RCW
/MdaaDCCjD3JRQN3pAz63XIO/+oKSxEYR3xYyuBcdRG1yuIf+qM9APqYOLAdp7q5
cbYaerChUvHucGyEwzpQYtxXicnvqqoyKFzP2/gcIHS/iPgAl2QlCTz0COsWYyha
TOBTYPw+DiO/JA2Z8d1Xyi5Fe/43U4fIF0ei8lbSjRbwqbyyeIRa1eynEwCTCCdP
oEOkQaXpJuN+w3czVSHl6dewRLJ+VzjLnhMA2uhsE0K+AWTNHYDl/ACgv8c+hFis
5eSWilBTyha2x1u7tXZe8WzWrb/Hs6+mVvObw6fl9/6r4YbOqHCvrSZsVcDogKnR
s2/T1Dth+JX6xjaxSD1aMywjtSHjGaAgBmyuPfA6u5E9YUpLvrQ/078EONhfoDik
SRp+xD+D070Tnk8bLVzeNv4Ky2vZA9J5rzQPPk6h+cSYfUMhFylbXpvsDx8qfyl3
Iz9oakYZjjaytJ4Pp6bADXO0rwsIijSfDgU25GxiW9f4O/wZknrhVByH6gpNUl2T
+JxrYwnjg2aQVHQIDJFS2K6yfZj1OzMIdpX+XVFzP+9BWuKad+EeR1+tTqq9vWPU
awedJHMvnvKqP4+p+OhCVtwwCOVUuOvJQBBX1Z+okCprlmecPPtldtDx94ggXNPH
qqP8m1Y6lPr/tyb/jKZws/rRYaXjXvUmuUr16Ta83xKS4Q7fCokcCta7N0Sw/XGF
d+BKLBwIMsy8O7RONUqe6MjNqmXJiSH6l530ek2eq1rC9+mMZRzzjK+JwOZJT0zj
j0mN6pR67FJ5ld3esTGg0ZBxb1B98le2C2k7BaZC0YYG5yiaIY6/Gwr7l574shld
jMQieQxNlaHShNSQDaYFmwdwtMPFkpEfUZDiKs3i7l/ToaD76DniSra5ETafYLDM
OXJoyzvxqZp23gZ9QNJKcoq1eMJWpG1WdClLZF6kbiT/BIjxA/s4O+3dmpkaW3+i
EbUaCUSW9vLVTPgv/D90crcfTrbByix7XLGAKoHoJJqsTSOyod6FyrPaltq76W0X
33XMzbDyu15ecvB5T0JJYRWmM973njJTfygytuz+I540zMK7KmJQOnfrVKSR4TrQ
j7i9NgzSNwmLsGQAh1LpKYAlRJqu/CIaL3OMABJviTTTwPmfu6RSfS/I88n/Vdh6
hUV+t27wGa4T5wzM9gdsz148jlgun6Cy/FYHpWGXwRigD5fz9wiQrH2yMa+jp38S
YZTSTZkcYnwG+jP4t2jHizivL1R0zB48PSY/P4N3k40j0ObwxBPtwmm1tuymblRm
R/+5ATJuqVTJGZhvD9qU588zc/TMaIxaniWfvKs6uBTbzvZSmuAihbJkaBKgyOeZ
lqsHV7ZtelDIQUfWOj7ovxIr2SljH8lsG5H3FxPVjV0xbcKN77kVN5qEEqoKj48g
ddZmv67CgbOft7Cf/QuiQTozngCURPbQY5e5abK1rGZnk60b7updua3bCzBo0qUZ
TQEF557vbIP8YUSaTzMM27EIPHZUhOceCRZrLkhtJq7XlqavNtXmD6QwtN+AxBTb
JfH6PQqOWdTBbsYkoXXFrDUavo/ere/X/gYQjaa8aUhPyBiWPTDffrD+RGqQODdx
eU2db4o3/QA2QRhQLkzQm9/z1jEM7yKfYDi05Rm0sghgCEiFMFAyBuZ+t3TxRBnj
66l2G6/pSz/vimTU33aJcP40BwwfIkcIukQoJ1NQlkGakBesjO5OH6xZNJELgiNX
dxHoyO+n1N+zC89nKxf/5PCu6SOhYfY8Du5TFrfSNhXGqvm0hHBhQcxXr5gYlnAP
Vw9vm/hrNBef+7wBgPbMJW9jWm/D98hpOCs7eggzZ3nIdJ3RYgiPlQM6CnISBXR1
3JtvLQ4DSqHINBYoi4wfxmmqBuDdRFuByyneTO0cTljZjq4BfEOFhQtplXVjdojX
7U+5Yt4RpipOM58ob3PtZvyGT82ZgSkx2n8UKEet0Juoejj9drdQwTjLnQ6279N5
VPy71WD+QMik9s5SfmIsudi9VrJiJnbDvq6Xy6synbspZqOui1vCw9tNiec4UenK
aVZUihiPjTdxDfs/aOURzIPWp95w0BQxTdQqhwdWZxaMxThNP187FvwMGsBF1I0e
KBNhBkypHT0nrAGl8OP2figpuxcTwwL+OqJSeuN8emfaSc6oUAGYouMaePGsp2Ya
BKJqY7cNkrg+MTlzRKh6voHWw4OX1a9qnKoDg5To19P9GYsDlJzV1xN9VrOQuijG
vgVAv5yFHomblhCVXC+K+3kCbFmIBpgHgX+OApGAYl5qWBhiFZctE0AiiAmg2W24
38bmF2tEPiiI5WUyslabOQPZPuMi04fZbYHVJ5BmUUJhRx7CAs5CzNI7AXoTHnAj
FXB1hBE2LJk7/hNI72m4Knw12nY2PaE7HXSISF0ANksXHyUB7Yh16dNtMX2yn8eA
rho+z/e/Qp5pGEVIg4nGkn7maCRTQUQ/r+5akf5P71GMkrtr/2rim8GpE6XMKC0I
KfciA5V+8q2dljjkhjJsE24SXqMR6kCZcMyz54xgRUNjnRZKCNsVyoYRevMjQfgW
eT5zfAnFxXW8qjYK7hHrQlNP59MHgcQpPcyIl6QfVgqrnrcLERFzHJH1Ad96Zv6I
Kv0hYcTN7uLlsSfC+aXCrMUk0VUwPPeeXD7KtipG24IjY5C4rpzfjGd8huN8zUAK
TJOYu6cdh+7KDLLwt+qx9kP6FcaKBmTZtdKK6N3ClO64xawJAw4GQmaWriuqJqSq
YVsdZoqobQQHNMAt88gK46IddMYs6mnWiIEKGGdy168DxppiEFKcrQljzCUPvw0D
hHtv9qRCurHkaRkgXkODTVcT1m08aykCqE4A9+ewoZhr7GAv/97ouQbYtWS2QQIN
pOjE2r98vBPeGmuq3IdCz3b2ozDiOYS/S+k0Q/if0mu8kTuowVCqNXeMK926VC/y
CmsiHtpPw3wHDVXM6TsmTxMHW1z72gAVTFqXV3gxNLhYIf+OkUmYeV9O4/8FucM0
CqiRzZiNkKypNLW3zsJhZa9CkMKRWJzHtsIGPpOd8CMellPX5e9IbqUt0kLcMLhR
uiM9Nsz5HYB04qtPHrK6JjGZWBk+wiW+7WOOAUqi4Q64k9nld7a64OrjWev+b6L4
rnhvQevYsjq9b69bcEZyJbPWrqk1Qz7hb5fiyITmvJI2lYdiyL0yZ/5EeUO+ej6d
3T2/0IouY0MrseZ01Mu/FEOrcw1TERtRRL0Kymp0AXiIHuxmm3oE/Oq4w9cV7RfS
gvK5FKmB52QFTVZ8OJ7Jhu7PTsZ8Ey/IEqEAonwc8zjQ0mWGrIfbCXgOC8S1Gdxf
b8zK3I00BdXycey4TxqdyZjFcviMHv7P+f+V+sqPlMOga9GMl3GN9rKLUdRoSPzt
vl01vG8Eo8ALmm9mAn7sFpk3fN3CFpUhV8K8EZMCwwK9o4PsfTrrxyxZrn98oAqh
5x6kvdEs8vl73UXZZVNhsGN59PXLr6SdvshOikV/BLvWkjml1HMej+K5PjnVLmeM
zq2JRymPIJFi7eo3ZCqJsted09tW/XBoRZcPjmqMVUjE6T3feDCYpZU2Kr6eewAl
gX7X4uL+BLLwJaBJLEnFNsUE8ntMUvPGhNhKrYUPaBk0zK1EEnNRfo11qvfIHmPu
9VKynoxfwcarL/GR/0waPXNJy5Cxiq3VrkbBEzCvT32MECG3vLXIpWEdVj9UY4DF
XQ8+5+sRKgordfJ0VJd+rxGDrlYcXPcXgca84zUPBXeyTIb1dMN3LD5+ru/rXNfO
wtolCHCe51kxlz/W8q7/gxLA7jtrKNX/dhTIycanYnRkeAcjSMozntmwj9qnAvFh
mj0b07omyk6eq60z9V5pnRf/Is9GD+ThjTetCr5T8IVH+hkIIX8YaE0ndu7XFWlN
59Dr4nPQFMWzaXDdN0cWATSdFvNKi6CP2xj9/+e99QXWpFOGb80HuLH8MT71WGcq
YmLTXNf9R8WkAJ0ZsmZeHwVRYIuDzLWAPMo5V21zK9Z1xxxkTQw+i2Eqz9L9/nwT
IoU0D/zk/xSSHpg9Ep2ZCbeMoYxaHnpUv45bXzKC/3O39ekus7Vm5UIXJ4gywGhH
J8S+BNhzrKCbSyQHaHRouZTJt56GIal8Eqi7tnPQjrNcyS5XspEb61WZB/tPpqbc
PY0kJegwulzEQjyomsAEHJ+QJ+nJacfV92S+CqUpnvH6pYJ4aVDmEkkKeRbpKdbd
t0UWnMAsEoTxj4RpKEcJl/eJHIehsz8vkGiCNvms0PjunbYrGRNdFDlWdrp5RdLr
f7B9ZB8u2CnX1CnInYfJAGEl32IvRWeK6IAz03LCTgw1UlSQq3W4aH+HSXrAGWPQ
enhowwYkoJ//KZIycpUX8etgVWtspYoTyQp+/cq2sMtnEE0HowYnU4vxTtRCysux
AwhKZoTjmFBRZmY+hZ7pE50HMOILBsPKZiXEFpVXq0dI4Aj55O6COsytHiF2Vx5y
6wSetnXG7egcL1O89tWxr4gto96qC8+Az8mC1C+bAevTxfzuskwSR1G0PN/L6vE6
69qFq91DAxpFFikxWV3N2ybM1jZtYwu7iMicyjvnsZLBVVS6Dk1t3WnVCDNNaEz2
rWE+IGQq+JnK1wPSR+u1LoUjSJcfKwdOf7rCVkfCjty+eGyNkDBAfoNR3GtIqPnT
oIEVt8WNrqMrLBPqXBYDjEau/6PQVZi3PLtfyWjVaV7KI6PeOQsefmoiBDs+YJ7d
6ZOGuYDuIJt6y0f8ZHXstfU74M+vVKzjAPKtxTqewSDqY7d87wZPeLX0+lzLGbkN
7xHwJUh+EEIue50EQRTLlCilvxXD9+5HGHhI/Qr432oNZmX6tY3chsHMYaFy6LAB
mmoOn+io2vlzyMRsuZpQ/SKU2r/57GayZaX0LtUZR+zGjDU9Hzfn2lQORJo2oqqP
7AKhOvi6d6KnIU5Bnd9us8frTHPupXkZY8T1IK9Mw3I0HqP1fdHK1PjQKA9v3jrq
BlofftEIclyU/9trafxoJ5Y0qNp1/ShyKmnu8vJOP10/lwxErh6qIj7TWaosBH5i
7WYSlk7Vb8T8Tke8hdGTiLe8pQ8lkaFs8uvN63pbn/gDWIL4n0t1v+UgVTCrsGCA
68FQ5E7RV7dhi/NEew8oV2XKVlCDcxLgkGAoktqKiWAdiEs6yLj48TncYorpWAS3
CdWbAJ24FHK2BFnu+e3ac3WFiVGGC4yk7i9fV5PE/5ldKbFWipHXyd1c0+fo5qGL
Hbg0Npig9ILuwAfMFQMcY+qhtzvrkSZGKOySu+f93Wo9z1bzzpwFAqc/kAj2GD82
plHOj0DzlBIjvN+eEWNNeHURmtJbAO53iZtE/0jegoYHY8OgpLiRbwZL+i/cgvV7
9eGz6a/zGTohZs1mpMsUZa5fWgVz20ZYHRKnoPEKOMWZcxL7Ea/WsR6ZZ3W6dN6+
hUJGRbB3dc9o9VjST5s1R5pp8hB6TAhs07UPYkNUXn7Q7pEQxk+XbfGSrWAh1+ta
iXEE22BU4pDnhi00jAEyuxtYXdPUtzT+RLWQnwqamKUBgtfhceeZaR1qNwrTI3LC
uwLEBiW9wfrtdMGriHnmXbgnxbYIib9CJbWTeeg5lb5az5cGY875k//T2LfRwHWc
Y6dxoTBrWWqgENoVPYF+dUxmKrXgYrKwDr2syDucoGsj3VC6blVIdA4tWUyhcM35
LVilMWd2QJpEhvh1Ieu4RaBtNfXoclAb8jPXF7NZvHxRuuirFAsx8l41R9XcCNzG
jhi8SkeGPK1Cq+8YeY3Xqgu5wmWtslASo2WHqe4p0ejwC1Zk4kUl7sZ+0fYEnaDr
g4UpnekXb5s1rXjZazEDV7RejL7fGdKqrFn69WzyTET1R3sfL6B5QQbBwf3SU1sP
hP8jS6vrXwbb1b4TIQXelUKxx18CyM3D0QCAauSUGG0thG5uru+lIcP1wY4lN7Ta
VysxD33weKrDMGiTfGeVLN4GRrK2CY2S9d6x7Zy20tCD8GrLmvxWJhYXisNVPHQJ
qdLCqalkeuTW3leqbe0iWpMjDTjgsKu1yVx0DJjoaK71tjPhAVPApWadOdmZZYMh
tu+KhVDJmvwvOt6zxrB20jmjMYcHPY3MAoENMqkhpOzse2vFyKAfNsheRZsZV8bw
U/zjAfUCQySJfUWjrQQLHwAlq+zuOOQFl5REdeOxZbN3lOevpemuqOAft5tQXrlC
PllqOl1FWCPwwj5OPLLOjOej5+4aa5JOuFzAI0+bYvGKs0syo9/++OCUHETEBlsc
L9+1VpZqKXj1dIzDeobs+146I1w5YuD7H/wiJ4dt92ztByWnEES5qtqv/5CNT7ER
b+OcMACBlfJtNtKbxlR8WNby4MfpGwE8GNGwxl5wlArfE3yZrZO/4/z5Oow2twM5
MBJ4uTUaEp/FaqrwKM1TRQVAB/x5kbx9SZdo2gYMFqfvZEWfJuQ9O7WuW5+zQCsi
lOhb4QSUNLQl2OHlEdVkiFp0kmrVG4015nJyMPsM32smsqZfbXqIEYgfrY7f4BNT
6Dzk/p7wTRLX8A+A+foke/jwRP3O9hmg8iB0Nf2idMbmipthplidRxaBUp8hcrq5
Y2p8pSQ0EkWv09a5UWHNB9LbQkESZ3Z6T9alM0nWV2h3vGXmqZxBdET4943l+uPI
RxVxKouDrskw15ce/5CyXYyO0JzvCBVqSuE4C/oib1NWOQxU35Bl9pn+nq32A1KC
mgYLXLoyvMBQwdAERIJ555OALnYKtL6ngouweUMe9i3aY4Waj97gQaKoJhheCJeE
AH9FwQmKBlD3HY64TlamOlsuKlHhHxRbew9V/ApiBthqVk+fRawVFuObsJhE+D7q
IDaXopJGSB9U2p3/yXYwGgxSpkxnnKSVO8FZno2tzr+pQ43/UwOqD+LvxaJWRpcw
I8F1XKqfxe75wAZoQSylu1JLQQ2ATQXPMrDJqaM79QOG/w32gtZhYnbOCCP/vdym
uHhCbXGI9Lr1pdigaP5mpzJfvPUu1VaBU/KcizdBGZlQZOzD5NJ4JKqu2sM398DI
SsUNV+tjkDHK2XBJ/PmYXYaLVbAu3ykJEklQWJmggCcDNPTLuZj1nqWbqJprovQU
XrY8kY68WKecGWRq3sT5z8MOy69qU2SIMxDK8mG7mNvWU3hxJ/IGo2E/lG42+irf
HkfwfacqNxG/aPFi7IPAo2m4ytLzY+2rj5uKGr/krNqUiIBXQg6Ux/ZjOUMvOOds
qlY7PZbx4K6h3GMLHgwWakv92VgxzO7Lv2E4oSa4nDV5Gr2TInKXi/rwLNU0o4Ws
6kCMlIWPRocb0NZuL5mDMKwmEOwVdLYEx4pJMVzVYSWdh1r///15TwKCNjrI4R1P
sAMm0YOM7hdm06gmGueVdSe4/ienumeGdYQjQv3j+lKCg5ssUbzn7sg/D8Qulz/A
FxdvDCdEdVNjPzPd1E2ByAtB/CorQZchf/ejuGrvDCjkOLk7k7xzPB10do4LYLms
m5E8DJg4+Y+46Qv7cBGpTtmJpi4zrgpZ8ITT7f/c9grWYUzhVHSkMSD5pvezMmd6
2ok4TYaCIDGUVRvleynzvhWnqYduR30XXhPElP/CGIXvHtgMJRguOhtEDrmrvUx1
Aqc+m+7Jx4pv3wnBglymish8lPoyCcvITG8jojJqdVtWhKoJK3Cb2f0OC4YTgaaV
joD+h2PtzMb8kul/IhmuC/2VADsN9rEOeSICK18YQYAIkhRT4d1JsZ3lOwD0qj8/
Mu11FgYysKUQTGPd3xE7jYjR9VFXyfH2Q16z8yHGwZW65vxrLQVWcAzvbWuLhEID
64e8iFbHt9OIfZ2ITxN1MiNXAmpHlKeCmXnpxh+dawrY8gNpwlD+9e8/lPRXaNuA
uX9KcMMBnXT+aGRNEMwcixI7pT+drLqRfuDeXt+7znOd2uVVo4F5cpDMtJrP8IP5
21Ft/6mxT62Aq7MmcjOd+nyicGmltGe+j2hKmf0rN6TzPIV1IAQyg2knuhPevhtp
kOrQIdoxCazcGjBFiJ4UWmdJUEFvGhPebgnvLZEtEzWhXXELJ7YfTg7FkBC0UUmv
8L5aw5bLMiX5DQ85K4Gx7bpxKqM/AYEdTE98gf0CmFcE7yo0BBo7GHt2fVy10Q1x
/sHSSiw3Q+1Qf16flnGF3VTFmh+1afc5HDAGY2D0nX+DfXH3bE1/wjOA6bSe8icG
Sjq5EmGY29vIAZ86UNCPPxC7v2Kr04PA9wVPhcaIVgglZpsgyJhgyA5h/seJG3HH
2BeQygXDAc6lvfPFVSDmQLscDvDL1UgNzAGtqhze6aT55U1UbtyS6g+MAaEbrGil
2bdvqI8fH76xKpJAE50zg8zQfEBRiBc2z5fIUbxs+OXsPRhJDZ4XZslKitRRTzVo
O39E2ebeP3CegB8sIYAwMoeaZ2Irs5LNdwCKGfrirULb+zkkrdtiiFQW7HJItHso
XsQ9nBJPQ41eztVorBaeWff7XoLU3eCTuAZ6D6jJLFbadLTxBpS+IxoSomImPQBL
tbJNWtj2VZpmccesP4k6e66shhgeK9xhkIfznkvtAvJAzrX8mfkMOdmK8puUnOSS
HVuwYJqNekSyu8l89RSJXGzRkdzdA66FogibgMv1+qDfs4M3bw/JeE1DFlFJ/B9t
UUn6KesGYdJxfy5JUf2UHtsKjbaXD1aZ/DIzTK2NW4lLqytQkgwkqI8eZn1awGXF
ObllvCkclw4/GYYGUL+VctOGVV9v+ZrZ5V5hCEpxUGkW8stepMALiAkW4Wu/QLQ+
SAaH/CydzZeiibSU56jPQImQz/20uJhHh1YZHPDsmP1Nh+86On/jQ4M//x1DJQNZ
LCkBj/XbssFWWgjBHaI9LHHg8knJpDZpNbk0HewAGA+aAmGlwp5qYpNoXypyh2DY
aKEFIor3Q/czW5jRuownc2Hig+lU1ZtpA2BtgbGkVRW7FzqyuRVBEfb+hreCrMuW
kVmB16D65EJGJdICVAx6Yr16HJxrZqzdJAk6GLrYuByECUx+hgMuUdEH3DLe0eht
AuBr5hbWyiD0+C6SOrA9CgqX+nd9BuRXY09jXkERrm9IfjnGAZ/WEmkR6kU6/pQd
KKnjru/HXpK3isL9f1T2WBtug9vRXxdbKTx/2f/b4pQ/M5sPGCOiUv7Df+5iGf7B
7rgl8vuWy54Gc4xfazu9j3Cje/KAGEgWbRKHS6v3/AEopPW6rxROq1Azk8jTX/w3
jYX+b3He1h2Mvw48kI41YrEFb94DIrAOa8pz7Gsu+/MrFKjS/JMdTNuK3+D8OTme
gKj8MHt9lXqwB2zD44Lx64TmnrLKpu/uVWm7dssBqz/LWZukqYYFbAAkczENxRAQ
eKwXgRI6lcBia8Y5uHI/Wl1dPRId0DIhjD7YIj2VJIl/FnnZLnWy0LbqH2Hhzbv7
I4cLYPGst+UQY3R7DvX7x/Q0jEZxS9rA9H7CJHctFDaTgl9ZKarl+IbFaFCLVWm9
a1B7iVAdl1avYuy9Haql5oitCqHRehCIYSJt16ccQD/of63PV/rcjVP7VRmj71QW
984FxVNKOTGRd4vX4uYsvXt/1nDOdF2VcGNurRB6rbT/i8vM+bgL5FM7OHP26sPc
WF0KGXDdcDQSeOHtbVCZ0JEkkFDnt+oS4a2os8xTNR9VQxEWNgr2IvElwK505EFs
3wK1JNfXxVA0Q98Fap3HbSYjNVzE0fTs6rqLJKrnFKTVnPZLL1Gfx6ttFSUDYxEv
nsXWgviN9IUsPbUkEGLbTG+jMioNra7k/dPlMq70Pq4qG00/lVq+kuyzrkGKpPIq
n22p69KdSIFQgamg+Q4Xy/SKIPoVDszPsxk615v7RGk0o4J4e2ckRFMB4a/2uO1x
1e7hydUWJ+Ot+7TxWMHl/+70sjC9Ag3w3wHvIZr/GWXAnbFfUUiqceroXcpbCMUW
wvFxM1WBegbxzKrwv9OgCEXZe9DPyH5+z21NoVcSkwWPPTfibq4PeG/itSnGLMTt
wcHS1EsYkeXx/6wcrCm5AokNV0KWz6YFzZRzvHQglqb1bzxn+98jJYE0Ovqr4bzV
Bxkl1wGyHmuROM8833q5DmErNNf4cqauLekdtowTwJ5kQ7BJI88GTdw4FLySuDtD
mfCK72x+vLkVTqa31X4w7BdmxI291x4fAEhp1ImrVO8mnfXknwT/QrXrxONZ8vRu
7+D+eZ2rmDKZS/NVnfOAJbbeXoz+BoYqKPopMi/mHmqdWCgZido1XNeifmxkPiLO
isMNtVaWUgcAvUpPojvL4uT99cmm2SUDWHlfkvBHMReUHfRILJu+1EsVysrba+ID
Ho9xEDABkVNdyHwlITrU5sevo24k9RIDTElndxY/hCxFir2kOxf32zvhil62aeQ+
RT+I9NEAssu/SzVkIMlx1ordREN9GOYqH4cbSywPe1235q5YAENNrxEV+U0aAgRd
LQzbOYN1EWvvPjXMR0fPSINR8vSKGO3lUENu05BGudozihN6u1jRSzPAHxxL3gCg
VUFcdc4t4nO1tPqhhxMlOzpiK4F3sAG4+jjBj/ewEpFvWJFnje3eRL60le5lFGqG
nkfp0B4GuaaxJhKgrYTDAJTffdCw/qRL1Rm/OHcGpatWAKHyun1q+uqjTX4M7HKK
mS1pijU/HLw37KdFQ3wPJkKt11s8Sz0u9g1StytCf4C5LTLx/lyhatzaNeIeRINK
5zItrP/8OoXe8NGQ5s3LUUjYu0QsfrqKIGtSIrrupqjKiWsdb26sobQ+tDzamLV2
Eyg8/6TSLmjrc7gTQR4nl9jjsnjZsfwgeAGkbFY9EF7cv77f4/HcXgs90wig2r9I
wVWMFKxhM/nzbXfhKQctVeBlz5kjMzXbGTqvyw0sqbzhfJWLNMuZf2nitE+ZPXgd
uXRtubFjCyEXMDJVkVTifJ5r0usmukbBBG7bT7e6RDI53PP7gHVrwernSkQNGM7x
s5KFV0HCHqhbsGWoIZ9xBZOrUBFohlf59gg3oSu9yR151qJjOYnUUtt7ee209KQZ
cNgs3NtnOOp6q0Wo8bu3Mdp6seBdKJCPQKJBjnqSNWyF/XipqG36kUdC7EjQZ8PT
ahIPXBU6/cyr1qjBWydGGY5s4P4+Ajd5/NdbWoMqN+GuxX8vkVHJlHuWkXOJKFTv
IsOUKxDF71+H6w6bCxk3q14qAmp32IHhz9COeA4ioNH7cnbuSBmYlcxpX8SDKNif
eSzzGGWG3I2MROEykfS5PdLo0Cn/U3IW+k76iZaIEdTjCzknhQO2fILenrV1oS3T
+v2aEcGblZyLbZvCPVniyvrJGHYnB4d1MVZ5UC82dRwMo4XRyHq1KT2fTod7agvz
xsGE7y8C/YAgGwfKPugylXyeOaxjQGiekM+HL9dCb2Vsy9exXNWWKv7tuwwGlumk
9fwPbLpxrAJ3l5qjQsV9RXk6GWaRQKqoV25/ZdH0KuCex72j0dyHLQPHRDLKNwrX
vQZAHP8pNx6DEHBF0EQRVvzN6EKMMObKXzeG2RXPE94PlG1y1tB2MqES48VOJp+/
c/r/Kcawuych+EOQBNMo63yj6OhjjcSC544quca4K0Z9W1m4B05/s7uGnlUYcUFn
aQOQ2x2yceBwt3TExGw8WoJGesEc8yJ4TzJKXSuO7bwiSwwWrRaVQtqiKW/LjWiA
UwFb5sq/17iUE/qCHPXNzA3HJkT6zmM84PHd11Nax2zqfvNhort7DfLygvjVW9Ya
LMzYSwJhSYKT6cCfELhIVkVOtGeo8BjjDkmXIhxnjYETZrMdqcdfeesnAJ1DtYeC
xQyuCfUE3ivYkojj0dxwWA1DmT2V4MzV6ym1jL4P1TXolop686saT2GO+Ihvaz5E
sym4Q6ZQNgUIAlOE3hH/eQ+NFsjQgh92orj67WqsXWC2DsXTm1k/9nQI2VjMw/+J
x9/elh1M3RkxvDNLDyFmlzjVHL/dRqN4wNyBAJSeWRmIbb3ukIKqrnHr+LQwQ6g0
ARC0hfU/5/kBHUh1pC8wn9TFofallaowf4AsnV7ABrSrKpTxl3rrE7iphONs+Nt3
/sMPZZORC3tk78FXozQ5wZ2CH4/2XsOyypMJXaVsDEpHXeOt5rCnBj7m4cX/LbNI
SxNuEciLTKji5dbepzBxFBLPL1BOZKv/VVFRz73UgLQUG+aHPqi1z+QxyQOLfEdu
dixnj7bJGGGe4himnfpZ3RSBuxTFUTnh0tnjxQ9Snjo9AHriHmRGtOs/FXFVm3VF
u0gIDtg3PQ+/uZ8P4w184Zm4mRkRF7XwznXN1g/6Iq/bvrhpoD0g0GiqscBCIi13
iINjDy5ZcLVd1nU01i5Ck8rvAF4nPPgPLl1dWgGvro70bnABxRWHkmo1Imx4Z0P5
LOyHPsaf4h3aLSU6xOuvu6cjxiLlRTCe+h/NlmhwDQRaSD7DHLt0Pl+Nyt5EgrzU
qmBD0KthJh+pxKeW5Jvk36zTBLuRt5Ddx3evOjXXA78DYydM+hRyN/np6Hucs5T7
V81WQXLG8Aw6RBskP5RMskMcrXEoxG4Yo0muJVV/qqxh5NgOHvrWW2vujIrk5hzR
ejvKclmukCgfqwveQ2oUOJMnGjOESC9kYACC+1TfGgqBAx1KaZqOFbLpc6yNp2/9
XQC9l7TVME++Xf5Zx6X6f3SuS72sfDguMWMHg06u5jZpPFnVrXoTVqBfIxbZl7b7
7LNFFbs61hcJ2/HZFfP/rWGeCoiB/WacsgUoet8eVvotRd8F1qM0dJ8b0m0v0Nio
8r8cQ/62+2Ost2LBTC69aL3OdpYrrdG4Lua4pjO080fh367bMWvtCz+hnTPpPEEn
GY7J/4TCnNNF4mDiCYck+rzgo7XL7RJavFutSEkPDJ6HCHTHbGrH9++AY/m4RsCG
Q1qoJjL2BI/Q0QLNcwpOUoFuyn/m4FcylgATjpJNLkKPuA9pb5s/tThNF2ewMOlk
uB9S4nzMJ3rBx3txpxxprxRxcVxFEGKUmISBX+HUuFAHggVk18y0yrKC9EBfwDhC
5LRWctLQ5QwlOEgQX+bcvyT0fUoJ9kSRmwgNQbi+qak2Aqs6cuqRxIZ0v8qXynXQ
BEnGcIBu6OFytYKXNX9pRPxYFbi056w+C4Q4wHYhtPcs/nT4BgDUEz7CwwBmATFs
0b57G20g/TRCFssC2jEDrI7WZ6mj0FS0j71KSuA2TWqVIKbFGeZCADJjCgfd672R
AmV4mbj85snXWsjQI+IPzYOjBdIL9ZiOzVVfRV3s/tWyQ49tkyuU/pgSFKyYWA3H
qpVKADVoF7bKqaSJ7WYJi+bz6QE0GmzB8FyRAFI092p0XfyvUwi42CJrBTYrPa67
CreehVyE5qoXt3MWYfCv2HRSB0aRZ5ZTIcPgjIflMhfp9pJyD8DtOg/CFXQ7RID6
9cUYTSYqkT2iGyCNJ/PGp54iH8Q9HenonIOkrR/ZltHwRBfPwBUKUta3DTIGIpIb
tGJN3/m+7q3DG2i/DPjm1VDHpGHpTG7atN2P794KRhabF1GOV1pN6cDdwhbSsGZq
A0b+vBWA8vSMzy2l4sQVih9UQTAvMMZQGt7mHUrhN0o1dS8mjcg8dkwNTFgXkG09
/jf30TTw2PYRGgwbG8KMJKrbxCg4F8Anm9u5oVtfK2gcP041p04vlpkOmwdxtL35
Xfy4Ef3z4j3r6YjNHvavSS/tLcwcmaFzH2wOyyCWIlA5YvgcaevvRKG+I0twcLdg
l+w+uf0GGLUpTcsh7e1AUq0Sxfug4EPP6qYQQke/fTphaFDbSuUJP4CHwt9JcjN0
YzB/UtUXfL3wxWZqAfM9rXVm4B9OFAKStplQrDR2YGy6+72eKLd0kOAoZrjhPWRW
LFhMa7rSyxY3TZQJQ1OxpnNczQ9H7t9ETsRXvyHf0QCL6TJxA7RX5/btviyWqNT+
kUvPTcyGHl0rYeMXsAHsT1WGoDzrbh52kMNhAAkiPXzkCeCz8o1mLRzQ/ZXZ0xO0
HJYaQQC48gVxCdu4OisBJqw4mj1AKSEqReC9NSAVPzJFExmRPE4GXX7xgWZQJM6t
GS6dTDrk0xBUP7rc2j18FpCjs64Uv7efalRiuh6M/a18SqvJdUkJJUc+00S8ZGgD
H8zEjllznc0ZXCAayAVPjzS8rLwUr+bAC9dHm8v0xeroBP6auZ5L7Vphh76H8V1/
B9zjcn2jauTtilNSlaJb2IsclT7D5YnnyBDdVsn+V1LO5VF6Su1ZH87VDBBSwlaY
/oO/Qasvnvw4hb72UeBG0Uc8S8QlOOxdbeJ3iOsNBEjKwwKK6aOLrpIKFVKFamWd
ueQGthjoj6Zbfzovu1fm8IydMNBHC1Cgen7hjLQF8ABmjYAnFS3lSiNpdrEtH2DH
Y8nqx0/LusfFdfVvqzd6oFaoixKFDYj5ZKyUwoIv2fmzRTItie69glUQeq3lSky9
6fUkxWsn11tR6PlJD/HH1NtS4Dx+KmA/1T1990epkaN+eeSz5RlCSms1/NiBDBEc
5lUVbl/I4cuHtkPqMZekwcLP4loaET1OjcAjis8KcrkuHwsOeUbd2Ykj6R3VJVMs
RVzHJxN1jsC3hCGdXsMrQgU/XvfNshWmZxy/deAJ1TBxpzWhhunwU4tPfnbfp+Tz
HsuuRzFyfGrm0TGCH06WYojnYBSEK2dJz4qS8QPW+FFdkk5Z5uHMjN7KN18tvxUB
Q2rED7/ukVC8S2899MOicTGmNBOYB3Wo2B23lzf0Eqk6UYd3LBRivsQ2Pt12lIdy
jtAs98rJp3QmM2UCKd1Hii8TkyoDAjo3D+BUce7/wNyWkl0E6DKP/zjmJ2t7dbMv
X734SKavQ0iXiuyrvUudBfHb974UHRKJiX04Gbe/TRvPWzm2pGJj+8+bwiSr/8qz
A8PuNO0St+stmfj8bfecQka7sFtQGeIt3ijiHx84ytXL65VJ0Xl9uz1rB980kP0K
+CVVeYBezJI/qxt0IMdP8cJxCZ2hm7lL5mAvuM3fqi63TrRrw8qweTJe6+lqH86N
csXBpEGQMS0g/qvh7SPHBxeaXwiYcFboIgtQ838RqVurmCkEJIhMfBz+kLNeg+PO
V42Mj/KmIgjHXa4ljlXu7Wi1+Yd+jyE79tAgYep0/drq0KJ9Hr9Tz6T7nxDc8daC
/p2BO+6AlOtXSDx+EfSyiWpFr68U2KCH2Rr1s+TGCM7r+4ModlPMkz047iT9V9UF
fSgVPqzlRako22ONUFYkW0+gKG6Ed/ujUrZI+gg3AY2iZoSAVPxVF4s3coUWAXWm
+PK5RXxhXh+wCilBtOD9NGJHXlpFUNH0LhTzQPNI+EyCq9k+fIWydVBkb0ORYNAq
Zxg08mv2vNXkPX4UzEXkrw02+s4zmNlLit2oCXlrup4lcdGBxV1oAccZ7zGprrYN
1hFLDCVeJsYTDUMQlCXxtaoT1iidz4WVCRdXS0Z7XO9Zgtn8kPYVHeKPzoEPaUwS
Aq2VzvkUW9v/atEQe7aAwdTcaB21Vsojp6veCanPHbuKVZm9neucnl+uaLMLc6MC
z/w/iHSaEfYKy+E+37sCsw5/t5qnErtvK4NTqFWsv9LRofXcTUmpiQc6TsgGmAH/
KRF07h/JggxUV/iO+fyZMhiMt0+OVxCOzF0kDCPF59Ty8tnMEf8ahjEB+zg36b91
oghSxERkHtitdwEhaix4AKpt33KLjoeag8g/S5Gd3CyKWTlIr2MePr2xGM7Myzu0
2DAmeTtYJ69gw1ln1xCc8Ylif/69Pa5N23Czzfdr7R5VgGBYfkiS5zkHYVxMjgLT
7pp8ajJvKXB8X8JcfU9u1z2cpbJS4FdarJjT/06bb78qDhSeixN2GLh1+fTnAmFu
SZd/Urhi9LJXLZ0M1D0IkMKBYXhjQcPdvGAqEAD9TDPncKqwhiU5yA9XDoH43p/v
kwUTWCnX8woomIUJc4pSOs1NQF8h+2dn4M6qDEP9WGvg33eSTH3C7odc8owaawEw
epmHsVvqUFsMPFu8Kd35hXn5PlGuBy4/hKG1/5NDJX2zjHgiImMswfgqImoik86N
f5SmAIKs6h03s/049ghdWs0rxXKDljExtxPalOoJQiz3WOrqMpLp3OtZnyLYp+bJ
GZwO3lK8DW8kvRfZ0pClQEz/k+vByT6LPkSCvLBB95m8Br2wFJE/c1H3G6YzItrU
EwNILsOrPoAAol7Ost2Ehqrg15urwArjveds3wbPzAA7YKvT5L/7/zm0xwgx8hAQ
+mCdG567m4Q/NxaPbIUZ3TubcOTAEljLt8MayOyQZ5uwJ5mldM7SPkevk4VKX+OH
vfJGfhD9+hXRuR+LCpRX1ymvnviAdSsFAkrS8pD4sqi6dRNGbs7JEihQDV6fOwox
HuWab1QUIo+wkuqLpT3j4djWw/Lm+g3zdIzIyUXXaa+zkL4xKy1FrFn4hQAG1GUC
rzwUzHUpUD5u8aBM2M7jaOZAGGzs5FdmFSS6WlLkkdJfi2qGqHivqULpYAk8A38/
Kk+4do0kVCH8pfh7CS+atnh+xFmzSqIVjbJW9MfVrmX1uibqJKcvDkoHqsI7xZuZ
dSczmP29HQwQbH9tzT4gqsdbuORcnnEF/zRJtmSuZfHWDzIHmnsebtrOcMJB4kLx
71y4tM73FTiBK7/8NmHcTDnpYkpT3x73klNOAzUmYl7BxokXc8Us+dduwrr0JsYx
ajz1Mlz5mbZ82XurR0itcUfGlhRgWNRhuarhQaifPFBfX/fZ6mPLugskS36YFho4
0vfjVYNQW8UBaiGG4eJuW7mhQemBrdub1Zrr8AO567XU5pttUEvFQ/F80h96DVbE
iZSJU+cpLHdDpNGmhFhLeNkSQfOOxXSyxeM2OvNjwxipUH+cbYneanhtmR3MuFNm
nD36kFwxzMtYMrHdgPKaEtBqbZI+5K9sD8Sgb9AqdhSbnmGLZPtDddFZDVXreaKX
ZOyfFflqIH0YNPIDTpgGzxHDQPXTkOdCQe6NlfKVBEQGdcn9FzoFobQwEDVGKChr
l0cLEm8/CaZTKXfCK32eCn5dmdGyUFQ1eJeDo8abMaHWkSUZdmOov0WZQyG1P9pT
aTikJtJu0Z92Jnrh6/31EaAKK/lICjlEOOhXSpwVZq1Dc2D0CQM8mqByw+maeti1
xUjn4uKnoUu4051FWUMcmq3HEjDz7vRHR21vDKL5woZh/dCYntMg8V6Rgl5eBRwj
KX8yA3oQUURPNRgMVsi2YeFYTsC0nph4nLOT5NHbDUJNAgvJ6Lr4KYCcGGGwVdFM
eoet13Mc9Ud8yeOe0+jLWbbyqmULDENyL8zwpV8KIQdGxBAWqbi2n31nAoo08dd7
3DBLZiK0OSA6IhIiWBjiSV64iP9h33/KPmxmMNhow1xkmYYJq+c4cm2nhx6oHh7b
d0YhwfByQbD4+NzKbFAGm+DEhjjd9GTlEDuVdOQKmqvOa3B457J1zzlSN+8b3oVV
S3QQSCgwj8xSBjSBmQ2ecZrDfjgdtfx24PpoMvbgupGN/nAgy9/O6cpDhNcpIieh
cAVyzVGiQFGfEQcBY/Hol/PpOLN0OZWS9QB/N8TxY602189HRY2sQPL2XoHC8Dja
zFmTdpUNvveh1g7TaWn4Te3OtJK+cOM0I2ewk6IQ2G5+C5QElLaBFyqkopYG8CBm
e0UnUuwyPZkqObSPquE2dgbKWaRGay+MVLXwDHt+W96DuKBv/b5uMNPTVsEdZxCw
FaP4QRCBw3tvWMJYKUR4u0GOx0dHo/91Kd//ElWMmuLESAa3zpWw+d+rqv14y0Zj
U244bJlJb4P4aVxeOqVrRDPm21xO42iLapUU8xk+38FJDPjAHJJHUoDbl8MM05N7
4VQkHlR9trmXozoyKZNHtuxymP7t4/9xdFXODHwJsgXPNSujE2o9GcQByU08OMwA
kwhQ+XeHon3FIfbSgzf4KHriDlGmdO1WWBiUsxz8qquwg2FGNGU+/UfQPA5p6zTq
7Gxku6f99accczeN1SZExazh7IzpypbYRpEd7FZYEQUWSCetVonUs5/N915FIlOR
91bvZGN5+RX8OVZtx0I7r5nt02aiCEnzTWYUsXJGn92hp1+i6iyRPSljfv8tNEFz
j2HnbGnGRa/SPjpcPdaF6eytWIL7GuJOL0EDUNmfRhAr21qgi5VUGdvr4X9t+iAy
6TMEgyMwA770yqqit9wmVCBcHglarW3w85YutFz6owu4YxIQag1DlGMEGBlJrbiN
95ZWZHOnmnRCU+ST+CUBbneNqRcmvng9FZ+/+iBFOx3kyoXKQeazqZd9sGXDjWy+
0SaUUQAuk044nr9wKCA+fp8KQ1lSv2JwL8rMTWguXtX82agN1YMMJdjOGCMVtqnf
gl3ra6tooCl08ZuGe/gW1vQybkIa4ZyX4W++Ckg8MNv30N0kd68+4jutCIclAmX3
kcvpYjBvSNupUFiJ4vaFSddPQaCocPv1kX82RgeVyES/0TsOOt9ByGCaYGb0GYka
f/xmEmDZJORRTfO93T3XvN1FOUpX4/wL/ZemiLYohhotKYQXJoNRvR02fx/TFLCX
/V5yy6HKQieHXm5/aXtzbjpr0F/760XMaDPfufw28m0/pGizoSOcZUTEyOiqIUp4
ylwKzQ9s/Y4ZqfV8ENNTwMb3Bb6VNSjbuEi00ZWpcmiU8NtAIH/Ro/Qkl+OiD8Fy
qx6IBmU8L6ETfGoi+g1Pt8B5w+APQ7cM5to9U8jQ5OEPEqjOj5dFxNcIDvyb1xZl
nDaehhPAmn2IOWELt6Zmjgn9QB7yrrD3DCKw0Wy82LvG/BGOsdbkwWCMEGdQmJqP
PlirkzmkCZD1snjCoqdd4RKrhqbEBrh2M5n4V/jQ2aKVyzZB5n3Fa/kg2ZGabrna
YM5tzDdi5VBrsQb0PtQ/TkmsTwP0yauZ/ord2d8AfazVSrGCBOfQaLODkAKy+Jwp
Jm/2HAdB1sUKaYhP9SeOLdjhk3YAvccDABhLeu1IqQgPECLy2rijWNsWqc4Vwww6
doOSGvVt8GE8v3xRKoXQ9VgCVapbkPtfm3Feep6jsiBGrWpJK36HpdZIX4xfRskB
aYY0mqdIHge+uS0R9v5BGenHCGCfJAh/nB9hk0aNjy08nWapvnxpsZfl04bIot9y
6OrPP00pCUtVx8As6NyLtDgY+MBHQghVoPSAS5sqA5a4tV341gii77tki9UcmJwV
WU75rEF1tPGF5nC7stxQ+2bjpsvR88M1Uw35mv80RiNX6mK6E2RNRYfxh1h9JHYf
gh62CcXyZOB9PVOMgKiJSGKPYCPAeq/p8CiAMI7Uqzfqq1rVRGvtusEkS0DBR34U
QjdkQW19+rmu1VhPYvlCtZ0gV+FTMpc1tilGVrCl1EVcDieFOI1WuIJy+nMx9Fdi
GV6fMB3n2rnq2lKG/Z/tKUGzHD9Z498zOqUMQN2XZfrQF5Q4lDMr4dy8HE8U00PE
o5i3Pob+lEN18hsTQtKBx/sneIL8lok/HAcizJcV4LlpAggyEVTClng0aEJvfLBp
yZyDBvrLDxurHrpcx28czsufTi+/j92GD8+yh06UH+aPA3tqjXJdcG6A82vOWOs9
F6v1PaVuTEFIhqJolj+IHFPKXvwUPP84rte1vZVx+Av8e/LTP4RYsmDkQgdbyXVZ
XUFqx7hLDpQjd7AF6fYoDKFpzQj1uV9A+8uO1CXKdU7mzCQMqrjhxaAgo0t8UiOH
TKYYq1pGv5F/++hCRkgozjvHWq+gXmHPpszQgVkTEFfwp5h57Ekq6JsxUqVTVK3V
VTxyxFFLhq+k1wx2+5fYGLEs3mHM32/aLiMDuu3gTOmwbAlpOmMhov+Ltifxs24V
t7IN21LOIzVOnyt/ZfDvgBi5bDrO+7qdgh84e3KdjpAWKboggAXqBcTEh5wspFaU
dshRNkjoIZKaZl6SA/2r0pWzMUWZaguxeJwufe9mX7tXeEGPYBjAzfhA7CNmjodS
qlGDFsl8umbmNv2VuM1rRllVeZ4LwujynJyyBBNWkVOSK8htCgfHIkLaZZW/Y6+A
odb017Q9VhMY5RppN5Rldvy83fbI7B80VAGTJwEmfdLtGoE1FtkSFg0+jl1pcYVr
Ohk2wVIo5hKKWhNSX+pfPOom8O6z/SvX55TzZTc12KAb3f4HJSLNuzIHbfU4WLjV
hvPS7u2shHF0Wh7NcNSMR7XoaBcG/gW83E1yVT3h6RK6SnvN9tp2XYsmCFNkxZY0
sDlrulJgNJyrBV5Gef/ufpcQ2tyzhDTrGr/T6bsy2ce0nu3nBLtUcaaM7DNsks1+
gSk9cTKARYFGhB+NR9a6WkOPYQoJyqlf0WHUzuseWVKoihtCNPbUfz4rdvypWWiA
9w0k7sf1cD0iHJyR0lkY9KI9ktWaIMedpjxlttA7W0KUOMBlwBQtQEwM9YltNXqZ
M2z39QKkolhhpq/ajO2rOuGRnefFDEMRN9MsMz7w14Ae7BXOdrEWWSuLRwKq10LW
3WEsNq2lqW0LhI56XolN3gVQdoI5MmGw2EbwvhjZ+HSyd05LujZc8SeVqZCikI4s
iXP3ibf9eVksfhAnfxsebHYpwYEmR989Ss4Zh7bcB6Zbt2STVyyh53Kp6NMoqv4G
eOVakRGC+TUsnKYDfuQBX15hgwcj0VgIVu9bMALw+EUQDFPmH5k/6kp+cpkSFX91
0sw8VRezMoVfAvDnPTKCZKegSfsLUaIGglMjv1z96fRRdP8dTJdNu3KDyqAmV4/m
4Cz2O2Di9jY4FqgwJyYQh8GB58njaD88iL7CiQZWMcaQv7DMuL0qcUsH/Po3q5d3
5UyH1nbJK8XBbZzqJD+Y8RYcaFEovNqm3HnsG1LxEtI42jpSkgGxRhelphjCljwJ
UDPTyRAHids/4pTngTRW+/8G4iv8OmJB38NU/gWtWgkTmztAqpWULMIAy8X7h6/y
2AgnoGhKLIKHkcPyuRdAqhuGoT93SzKlD/BFbnKnfxtSOWGOP/5sabZ1V2qJVMOZ
aBYbKtMeAF5onv9Z0/z5D4LK5kEbe9fGhd0iyaFzPlK09KKFKSt/3uaupJsZBHGk
Od4aweT/FxozilCZnhWsAHWg02m+t5rtx6JvETYog4Ie8ikriLQ0MdU70kaIdvWy
U8Nn/56r+Up2K7DFks5d6Z3jN6qoAfN7qjuA2H8ntO14Y3zJIvQV0hjMw+5LeLoW
vDWqhAHHlMmARYUaXJcgN9u1CLfEXEzWiHVZ3aYbHfxGVf3WpqXzrpX9N5Z0wFXK
3BfbnaHubMxTuZZ430gyTTs25A8NNf/2h8lRHnuGdvBPHFCJlmD3z+HhbW8p3POP
kNZeYu4gMLdMajZe4BUbBIdvygyzex20Qu2IIP7I1FXgqyfNUZrd5911ax5/zL6r
ZiKeD7kt2uiR+sd13Ukp8/Ns+rqhetsgY1mb2eMi9onHpqNcQUgYJZmrvyzHRnZX
fn1VZUaKM3idl/+KEVMrJGeyh4zoiTms1D4urjIxOPlmLICfyNzbyaRV8xdKT0vv
mUXwUubo6fku7x54jovTK3SC15QeeOkqpbQCyijI1NlT70QwmEbZiF7WzJSCwVoY
2icb8HiycPt2S2CW/ziORPvYwLRG+itbH4ade+iFFS8ErS5Dv/xsuVl2Sho2PLeT
JYBL+bII/LhbP+oz7OHHSpLIJn3hhAHWJIN3Y30I5tGFg5YcKluPQ+YepqlgphXU
7kIW9Kf3lppu204ha+vFqcP8o3cTENYNT7oYgO0WM9HrTweXTgMCidM7esSqX4rl
+K+R6EGxAJMweH8HNraNqTxsBCs+ixp2mddJxuFTP64WDhRxlTKbD5PyHkMbwxla
rXVOm45XSlq0+67ZM5vJomwothyrtNUMFnSqQGnMtBrhYlJr8GZYUwnNASrZQf94
lVhjnWz33ln51b6roZ/mccsonOcP8B57rxJgPW2wDnBAMtjh5N5MZow4UTdLX0CV
Q6wpxQHbLmvSdsQqwB5ng5DCs41C9WfgdPMkdKhXwOfpwBzzkKTx2SVb9dj17X3R
hr+C6Qqh6W604hh1+M6ExRE+KmRGtZx9TKhSIUHvdGZd2GlLm4PXmWGdgYk5zOwB
e8Forgc1my5e9QzWAS1dmGj/CXsVZWtuXoWTjS76Lrep9sibj3IUy0yJXximxDX3
rBx9ZOPczfzZWwgVoDlfW9Drqt+Ik7N3PvJ1NEiCwBWcPgMBEBcg1euXbbYCGVIu
LeDLAXVmKMukHafY2Wn8xK95fRSRMbrE1iCwO1VgUXviGIskMR+QupFlFSrpKogd
6o9BhycqHOk7K9VvVZDl/AQ32e/YADIXKMGO5cs/3o3YYaH3QDERIzDII7TL3bkB
TpQL9w52kWnABdkyrd+wYnrIJj4l9FhFogiGI1L8Own9AvUKpuaVGNfzHX6hY8w9
spQV6bKITaY2MeHD7A+aBUK+yR4EhHKdulvNRkve1dIb2Y1UGJi18mmUNTuBWPdP
/37OqVzhcJrAht4MwrYMyH/j+9aYJ0L4sDhHFjBd8D/I0cD5ew80ZYfnAYrdqw6D
Eguo0SoB3N8MQHtaxzXhNx2KZ+/bggksQNq54SLkq6J/4AxQvEc7mJ3j/nmfMUg/
JlDwte3B7pjvGInkC5F3qhxwFz8rjMfjaJZTcVGhrFE6+8b+s8F8qMlwE9mbh9cB
Hw24IOQam2V2WryNGENNL4afhyOr37UV0VDI3hFBmN8IMDTzpZ9GurKwnZMOOsUl
/uJjsGRXaKGKkOESR9KZpmvdvng6HWxsCcoCi8L/YZKefXiyGRKrscCxcsSGtgj6
iSH3gTNzesyiwR7LmBi9H1tOS51h0ix8B7rDbvnky6epKnRph9L5I1CQCe1St5AI
/icdM02YH2qjknD+JlBY1XNQV/6PDr/gzBamNJbxGXNXxFXb5GVL4QsBF2t8p2yb
67T3k7jO7NsNHVrh2Pq5Ng3p+FguvYPwC1UY3AZlfz6MsxPeuB9dzi8ayFvA8zWY
snYD3hVmzaHrp+3V2Qtpk1QH8IJ8GqESWnMUHiVq/ngVgpZxVZ1H4KFqck1WX3BN
1AGWU+sUd5xP/fuBfjHglePl4YCh//bldAvfeuxiLFJX+/lWpYAPeoqlxUXRjC6c
VuWopSev8iwh4yDt94TDPzADiaWjqMfWXAioGR9IrmMXJGebBL6/4zNZLyup0MyB
UdhVZ/fqDYLU9fqMZiPsisKTg61G2eN2GmHPcdt5PYNbfwMix0USGMA8aHCeMG8m
A371nM3GLXe+WcqFq7hPVrGMoEfpbbfZEfCF7f3NwTiak2ipl9cuANqBAzXRFCIY
Gv6iTGNwp4wQ3HA36MYxyMUTYGfWGNul0TRS5eSFThkmlCRUCwQ+FTdUnHQ3FAx4
9YsUcEJho0HaLaOPZG+aePsJzM+4Og83YOR2EL03WsiU7ZvWlHs47Kkzx5FGBUn7
4yx8CkB+MTUcx9YiVT16xSkjFQIEnfL2Y3oqX8Vs8/VCMhBZw5LYXyD4nbkeSK8l
4UDJ28DhcfHYiv0QfXPw+frzrzkBvYd9Xb918Nq6kL3LpZRnG7QLQbNaNlthcbfm
fN6UXpaHkLpmRqHxgPrcGXJr/89WUZu/ZtIMlLlNUjOARfyrVsLwH6uAEU/a6V6x
bEhkrGB/6L6Js42u46RYW9PKRcJeTel+dO6+JctfH/CZpKW/0lS00PgRyeOVcZYw
1pdRVuJoeA+T3/2aBipPC6piA/50olyrGHYwlRFSMjPpo/ZUMBav8CM+q5zsQnho
j+H+PLkJJ48taDW3+3cqkGi2LPovtHBOVERDgt6l43SMBoLfgtv6MqEcqUDNHz5E
rnGsg7f8dydEzP182dpnLmJlyBO8PVyCCYrf2SAoyguiewnGZJ/rhGib3H4w+mnj
IqXplJYKA2tnpRLCtc1kj82Gqam7D3q6DFQw7CqB3QF3GwWInY9htQHSZNe3BDwv
+JfbsyKMa2lz2jAAF+7M35E/HY6voiPf4dIHn6x7xNHWckG9ISHOagjO0qrDnxM/
rE1/oZkY5oZoCN5tqU3gxSQiOou0TXdDCdah89ibqcVmAnFzDpWlZyQDiI5eUEJX
x4k4n4PWn9sH42CVc/rlbr4YROKU0xIvaj2VIsIuZ/2NV3dSdi2CCLzYBHAswtHU
wsgKhO0fOvuHPcpPOVIPziWxeFJH/1f0lXottrrfaz9e7Z057SO5vmjoe1hb2bQv
yu1QusS3dCyCBcODAI9Oo+4JFp8i1UicVVBqFV6qy481/8uCROdwVX1mDx95Jq6p
q7kVz+wmJPFwcNA5iXx5s6S58qGLM2KWyuVJ4fQP05KxuM7+EvbErZr52H+LphzJ
RNTyCd6iqYhR0fLBUvu/t2JtG7/9mIwOtxCIQLQ0ZdsFpFOjGB7fCKRQQAhva5IG
jFQVMmy403xIwDS+b5igSeCwomSdKmOdyCpXTjr7RAeTDzLhB7+CA92xMvxR/HQ0
o0Q7UqaQk/eo50rBYKu42ZlNxOzNqOUzczTLnvadOPrTz98LLXjt2beI9YL04VTG
D+59miYmEuSxzALMN3JlqbGIMzOBTpUxwTV300TljRv1m5SMNCc7Lg43zFciR1p/
QbkEzS4dYB4RBB7PEEAYNc70LE1UfHvpaS9j76+ziirg01tQe1YrCZYthE1XXhzv
Qttnq93tfPim01inRN1ZpqBx60DjukbfFKIbmBUzjQLvF02XDByF1Riw0biikZB4
TDOIbaZtqgoLE5SmOFCTji6aRSDSC/Db0NoiMX5c3LNuXFV7dsSmoQD/MjSyV5nZ
F0ZBNaFxf2AON8GuIINx8WGFaM+JWq3SHWOJHQC/dHgbB1Qch5sjepEnPj/ss8R6
BbmdSqtOhmsdszxwp+kx/ckV/ENHQrH8jNl8BcAOi/cGDxDhaXrcXFtAeWwre9py
mH8s5GLTupd5PmwcAe3xUz2EgKka1Uug8P0Ymdlyg6P5W7edqQ5MwVh1dTgzcBjI
18z8aE2vLYdxs79NL3sdCX4sDqIlM1O3bsrJe5YIBBNNRr0JVzHrpu2/YN2bVK0B
7TEG79jDjHpVqiid+Vi0tFIMr7uInvzlH1MhhOBMoTmoWTgoz8ELk73EC+hIPD+n
91WsPF++elE4Zxz7HgrpeZQRqRk4k1xH0LGeGKNELxWqBlRfJUfT3cxHfLklHEan
VmGaODEMyS+LBBqyqJsCFcC8GhPBOCWjx0cdeC2KuDwyNtKMXB/YlC/fIrisbS5m
TGd+iuW/m07NwsRd+S4RYe+5iO+KqhMWu8W/ePT1mHhkctcgN3UEghszlSCMfGJK
3lGy7ddjkSYy1uUeHOC/zGbrYzBS9/TVh4kQBrmTzSmcopl7gBF20+uVgc1NpRNs
GcJKOUY7/NUKdpuNK21d8SxJSYU0RZXOoaucZiUhhEZgVnB2YO4I6bqpKh80ISP2
4WMYABsKSoKgf/85rtYI6oGQEl+FwPBmfBE6/LB+V3nuDU0llaI9LUFDBFdAFxDN
hArh4e0J8wk6T7Ao0Z3Wh9r1VmkAcFdyOSi/Z9N+4oT9SidgnAHzTF8PioQzVShb
Z83wVbUhpG8cxzYovY7IANZ8ThbBvhmEJ43UEuT1m/j4PgZDAooxwwn5IDPcDknE
echTLKdsBFrFel8prBa4ZrXxCBhFzMpyCpk8NMmi1Ldilyw4K1guIQy/GkYarjjh
Oa1vcq5LTQ+EGg8y5kFIBXUls8rV5E/TWURU9klCiw1MQzsyNhmFurffG+vAihMw
oY/LhvnbpY0jRz7i+JKFgutTFr1VkbqPLsPBQQ7xe0NX2X2eRLzj1Ws8RxcmIrju
LuEYIHcgJFETAOJ52O50Zsq3XzXyPGHQOjAULiS8SMqMuHlrUC9jkMZFk69lq49a
k9qiWkZmgvzpaDs19dLyyNNOESK1MlJjWOSX3ZQJHGtkorM/UBsAY2Y1joeMgF99
7Inh9YOyztC1b2V0fcOW0IZrkmULQlw06wKtpWuKsU76QdoyyQP9vei43gPaWAQ4
ljW08+cxP9BdXZuSz0TvAbk/frRqqCiF7j0BFZh3sfnndY7hcQGYqZ0wLLgisqGp
x1GNiCi7VvcvovY5sQxVFAJFtTM1EAOxoYY2uKoDeCxNqHx23O/maSoTyGBj25Q2
pItmNR/EK9YvyBTw/W8hknTxx50InP59KlEmDJTkQFk6KzBvauIp/SusUCpnuADq
QzxV4KgdAdgJzg6Bt8IOs7aDkUBwWky7xb9i27RbIuUmgQWulvGesXDPeYDpbSJD
LrJs6Nx1pHWplZ/KR4fHrRruEEeiSKAWP3m4MAg7x8sclNb9VNeyRUnlEhQ0Aok6
k+ZBIS34Fr+UWLZdqrL1IUKkCfiYG5cCplAeJQKNh/1uJtQt2225ozH2nXKvAgQZ
UmDA2ZkTtJ74CihbuSI1QINko7lsjzE/OgFJZhhVNL5TMfksnVSCHeDs5RCoDAcs
RnTH3pnEaGUyQfcBbTqW7eMBwpH789dI4e3vx2k2JSGGyO3tFvEbfHwMyEo7SgCV
eWERzIhlbOL2bOXI9LLGRgpr2MXB2M19vPGkrYzuA0zjNrlM6GYiSuq+HPSE0Yss
qOjDBEyZRSFwjxZTC/nafqqsDbIDQ+PWsMMnbz/CUP2x31k6HG0Zqfq9S7UfYbtZ
j1ahF5SVHGJJwCa6u+84TdWt7XY5SX/FKNqNwFq5DYzl0beC7kzgm+RJTPJeCs1E
fuY/6dUttN1HSzv8NbgWatnUcam9A2KMPjyjjtIYUDJil/FQtGYXPjogcRKqkCLy
ipuYHV81iJUhLY8od83nQ7hri6+EOWZ3epAHgviensGPHkTPd+PYVhtwQ6Y4Pg81
pqNwbIv95WnHhEHgzxfjJ054mqHE6UD94tDMiN1QNybWgzFNqsxs2VnXJUgFuBrP
kfCz+m2nwHCN5jxi8AJJWsqxklMOQv1mDpMiMF5kMxT/gBRpuwoxHypHmsZg2+wA
8X1uoNHLk/5XpCeqopISVxFBprbeCHOl/hLjduzFM9xNl2RD8j4rMLiM/5z0noWG
BewpDAbzjEGNJqkeGWlajKdYxchR7poqh9oTP8OdHks81CP4qz6EDZh9lLLahDks
nflwT011hKPnOp+Ll3wWK5GUMaDy180TZ/2LGRXZp8QQEOtoGdOyRQji2T7qIQzI
/uSpyyNzaSbSMZQoKAE4QPf8bMi+50MTSxOC80yKePFEv5dzcZDWwsPIq3D6D8ep
b4Gs8V1bx8oRzgwERe4OcxVtqer//k2vvLbA8DjgqtPp22XkYzj33QLUhJFvKXbA
rvhq8DofOjIuvUoIyLczt0yATHhGn2SiYMlcWggcYbcHr9YVsccnZElypAJbsswi
oEg/VGziRQxw4Eo8v9kJQphzHiF8DK3wK5hHFe+oY/0J1h03oBhfxjKPCuvHWpy1
gZ75NuwTFoV99o5KhMzIpX59qjaCX868knFgvq4eOagDfQ4xsJalRNk/XFW2aD8f
dGtoeWrGf1EdfB00SclvGer75N2PzZRnok3N/2Atnrk3wqL68xNkhdPkgrndIYkD
89YJuAH4qjRqy5HqeZxAhe0tUadr6a3PNi5yf8/F5o+J5sBHYPjmMs9w3nZ8Rs3A
46cpkHBO/3Y09X4BXcic9TFqYAn7sJKM9u7SwFxf9xIU3d5B35lc3NjAsguOFpDP
NuBCnXnMpcsZi6GkCwcbCjr90h7Eia0ZCPBDbs5lm7tOt6a2efwD7db1FKY8EwlF
/IjhctrHQ5vbT8vkejW+IaIsxmQFf2eVYdVT3Dq1tfCE1YBFZCyaT4BFlrnkibQZ
fst1TNI5VSo4B8ZRty1iLw1Mu8Jyefv41hZAwQlv2XphgDip0GS1gw+fFFKVT30O
i81AM0oAtJGYBuZ2T/Gx4Us/ij8DEwJxP6BpkJ2ttFDCIEvVts4kYL/r/R5sndPW
9nrBd6H9Nv04S1L4xMFo+dZZmULCjDYbAJwoifP8JAeNprPQ7nCOpECXHe8As984
fxiI3p2KJHlgZG2mTSlP3q4l730LJNZsZ63UurtWPLtKlUXYYcgW2tY4147pIaFo
sN7yMuW5lzjh9PmwPUSmNd9ytim1WpxuWhHrMUerAH0ARJHMdllKc+vOqPC5pIbu
TiAaVTiqnLzdRTOuup4w2lSLkOQYcUYe3drvUC6xKX0l3l5dIJH+Yb5XvpQNW3hy
g7RoSNjEdCR+c71r10FRf5Kf4HRPIM/aE9we59mu7e2LqwmT92YRbz9HFpB+UH0D
LL4u4ZQJap5usf37u3dkkstte487Gpc5m1URBjmpakJR/o4qOZq2Bu41eqJp9Dup
KUawiHGWmyO3ZH7LpMM62xqI5FEIt/i9bOeOwlz7G2Az7BWHcQ4fD3iHUg50wnAD
UBTmQzfphvAV27A+YB8dLsaB99zc679ZkabK84Q5sY6lEYOHnlrf9I82LKO6pchy
KDfhSAHztduZATwNaTC9lhJFAQua3ES/msI3/hhNTgepVkoc3rI8Uk+bHmlkA/1O
Ecw5GlYyL141l0ihczfW0ieFOmRt0pKakTJ9We4Wmj5sRmm24dGf+77ikkHkHqXi
2u1SfxoDB52l+uGlPtTD0rK09FRi7ZI5D2mSU0bUqPjPdXGHAAM//Qx+3RnQH1E2
mkVTYg75DIAFmrDD16T50zNbCHU/6U/TYQOWaFRFJJ7TW36fCQFE/r3O4tiDeVeh
xlilMGJS/4ylt7HgSUirvW+y5Z0frHvosf6soHPzHtWY31B5zJ3NJfA2sDSUVCSM
KJxT41HsonMbOOA0bioocBOuoBkipCUyWYkFHj5rMsfsXCRkZ0MuzX9RF33qmVCd
Z5vZ0t0+5s0AOJ9wFkRphhzENErxEo56bIr/AB3YN+cL0HRDg7fszoHE0L2n1PL8
xMr1FOwao3vQIsprRoRPWT2ohj33MeBI9CEIZ8v+BBFAmWDwgzNV4c8PsXUWx9pB
nJQFddooxQSDWPqrx7OpDOMRbxyW9Uby6EbDoQ8CtT1EaSgTT6mzDjATlZbD9n0z
Zh9yBKYfuUMhXdWFpX8mULbfGqv1bLtj1ci0Y34bFIH4muio3XF35hBkC33odCfn
Y+roVXu8XSGXkL6qYKFp9O7YgyqVjgASqo4VgUq9v1yqbyLaknuIDruh6JzBxG7f
/lnAqi20+/Nm/2IXC2kucFlgjb4uKFPuiqRcGWPata7Ho8DwtlPy7mRWkubCU1m5
cws/5w4Fe3fRHDDIi2eP1XY5ZhW1tFQUb5EnxJ2GbjylPX7Z4mKKNyv+l+O7BSDG
u5W7Wt0mjbAChct/1Avu4SMyhlK/nLIOc305vvct0G2ZKWOc5dTaAYzkQXyhz8bT
ajdao3/+6Tq/liToKi8tcRXBnadpVMAdFwJsLBznImxBf6xPjmK9HdKGuDHyK50r
LiiE/Bww1lZUS42QKT0WDsoH37iYfjkcUO0+7dI08s/FpLZfb3Z4jOZYOdrqPudV
rQK8+8boi/mrhGuk86nsl6jfsAFwZr4Uuack3Vhluzpa5XEWEvZ36pvNajX5LxPx
9hBUv93jr9u2VGcvckeflg+DQW8mtfw5J8U91sGQ23bEGeV/SlxZZBD6woGOh3EE
r1KMhWlb3TVio8Tbare9BPr10Kbjk53QHRICN5pAOxUbmnDy/d5JrJd5d7icZ3vY
ke593PcBQBQ27ayKEyFpvkCyIcdtc3YWlyuj53QV+gfd7X+y39qxqDeiiCRzzJkB
sOR7q03q6zQ/dd2XRGYM2J9gOHjrWTKtNDUzoBxGqCUOGoxPFMFXFZGfC7uWjJw5
QzJOidoM6OIaL6KjKIHIzI1cGLU3/xxmm6uXPAqpydZ4gHv44E/IqBTIS/Kuci7G
qbNCuuXfDApKmbDOz+okQ492KNjDVM/etsU2yM1u3Ae6bcN3vj4LZzmnbYJEcdPF
aOkw9rRoAdu+muJ1E+rorO/H20MNiYYKSoBBI5IJUrFOh6oIUgGOxcTOm3gpHmYV
zsFsDnuhr0xF10TaMxWc8XEvBtjRL64hGNO4iIRkL+/f4OnwzYCIeFaGJrqXMMOO
F+Cv1+JBXR7XXpLxNyx+CvB1Hj36xtDZmYlPo7+hTvnVR+OaMn15G/XWOltQvwgO
ZQSNUfqvFXocA/aiN1XlvCVPXJOuOXqu1FsZS36XZw3TAWc67d1GyyuX5zEXfAH3
tWTVlgDXaZ6HCEPTbyb9FVTlfyyj66b06i49Gq7mZbaAfQbQ67KUQv/MBn1WVq/o
dJXZDrIQShtiYDulvKzr04KYPbDnZp1WxzioQh77AlvpYsiNYw+x6BiCfcRGZnNC
ABoHg/Z26SdpsaPDArzVtB/bkVKyye7Yyj4JpJo0DJqBIpi+SFV3Y6sPz0Mcx20K
mHW7A8gG+DS6KY0ad0KeLhZJtWXGE69U4JcpTSDDiJ97FFXHRO1irDpfTGioFOyz
fTTAKPOV7u4NyyULCCg01hrD5CwH2sAXMpX8pls1FlCWNKlSMm6d2B4+/i0kGQRK
PRDHJvfVqhKE6vzYlhBc/XRzkL0AhvLfIhSQGOU6a4VLIvZUMIfqRG39GZRnVTkJ
pvhOSodpaS8fpvQts/AdBQKuOYzpVKQGFrU3zeawte12gqWpkYCZ4a90SylpJwvv
/lS5vKi2bFy5qkHQ7YvcDQahE8jfsd67j1P6TMQxaHcn9v/ZY3sldrShnHBB5MJz
RVK5SN2VAdh8t/IPp69ZsAb6fhLQBO9hXjnE2JVTTbWBEPM/xZ/38YRomRSOLmS2
BwDZPKQrm8614A+/b/gIeTeXDA+gD2ktUDUlBjNaNhxk6dlInMYs2gzKbKzr8/lF
EBoBZruhpSI9jXELwDJAU5+JuRWCSbR6uKez1CzvO1LcGc3VsYxu16qdVEfanG6m
lUSKV0WYotwUEmrTAsSFXI/0kHgvQgMwLqvi0XtfS9P/ySZbcElVHx+yci6u1aiA
N6bEbhRcW0hTN/dc9pRWkN5YWEdDPtfMWeXkf447VBrgO3ihYqxutsnAElkF1PHS
gy+lPlRQKOOGetNcwMicvuBP4fj4ppcciY/FYllsJA5FkKtzXCnwYzK7RSVj9HVP
u3I9zfRK7EKO89EAmdWl8rpr+1tRMeIq4UQcRXaZp3U5VBtZqZ6xT7Zl0yP/89Dg
MvS9R41o8G6slz4bNEnnHsN5Hdny31JH48aDerXqo90YTW6ErHlGpYI4tVAz9BXj
AW30+jOp+hWXW1GRHeNG6xwH06TjYpwZmFdzC6tHCO00WcPj3ijeeuA4KJ/XFkMF
wAh260+2P7i+Xp2jJFhpCZgdh1IG7XabOYlpSm0vmoP7Dxy1/K/9E96I0SDlETP0
AN2l/aOoBoMmuBMBFkuLJmcfHl0fd0SmKsSu+R8I7oBKDyQzvJp2UdnSkIxWVgz5
qt5fAQhEADybx1Yv8hJ/1vWGABofkeFfDIrXf6O/59xvmxdNJut43QHia94GH31P
LDhdQeZMc2p7eMhcAM/rjFrgAANihM8XpV3tHMzdEo9CsC5ciHVRP0Yo2pJ6qLpd
ETALc/rRlfZkfqUAj7ZLvoRR0mP/ofZOA7k3eiZ5vjPM23o/xq7k0baaJ3pBnTVl
tfhjVQtxi5xeZ7IcNr1xhbIyJ7SSMVGxfQhyDaMY7y4h+jIL5ga+0M7CUfFx54h1
ZOG5w9t+8xdFFp/tBeXS8ibjAEjZPxie6nlJmNweB98DkYi226rh53eRvo13CRFt
2+4neCQ6GT2HTsewSxvLQnCq7Nk2M+lmJtQXCc4ENNL0XD3tN5xr53GHo6uOcEyP
TqdJ1tJSluP2WD2hhpOimQEL1/fri5HDwwYDqdyGubOHW8wFCwYGy1drnLPpB9Sk
O5qFROkSKiOoPzdSiHojtAXr6eORuIwY8USPQLTMIdXMtK34Tn3GhNhFA0IWa5zg
2wM91Dxs3C4S5DUfyAF/tMSbPzjHlKSePSfBhSinys0cZRFAlVE/6fsb0Z/w2t0h
eDs/Gk5iM7N1feoI2PyTtConhlPwDmHKaq9ja2Ihhbvq+t1E5IPtfgDyGxolm2wE
vukJVEVdyWpsamJiWcUoDXQrjx2debKbFuIk2NukwEtSEnmV7cRcZHH7pl4Ojevc
tZoeBXtp1ztQi2fF4XGxtq15ejyH/3CRWS8OvNDgQkuvOJ1gS2EmfCUbKTAm+YkQ
9MLD1RzM9kI9Qw+3ZxqH+HG7WgMKrIQibwhYqhAAQEQc7nZObaARPESpwVRu9sGD
hX88ZObRvSRGifnvttuKhrBZrpITiOrNykdUl7WtWFiOL4NBBCZk94W1aOuR+7wG
LuObzlLkMm47XlbMmu651fa3Yno0R20ZowKxIEGqdF2GTN3h88VmMLkf1L2nR9FR
sQA19UD39p+4rRPFvkhOT8rQ5c95C3NMYERTYCyN6uAAozufOetcMW1ZLeOIlENr
VUvYsBkraX9ghmr9Nof2UYlxqB/7poZhWwtayBlUSW1tr6FNGKvOfGaGNU5CKsBg
Xt5fFzXT29tYuAcsXqglMwwvKcPMcRDpKU6PxCqEfyaRsESkh7k2RPrjUSLUQn4X
mUE9LW9x1htcmzr6NTjd+kXSoed3k55z48Ag1nGDwH7iMpXODKhQ27XVS5Kpd2PM
Ye9ApaIHkTLXYBJfZ8DrsK0TJdpHRldThMNccPCvWgkhS/65jssOHeoLdA1H51rK
cZEkK6jlBBH2gaSqXo7Hy3mICe9lT/nS9BzpRqDlSMkPvjjQ8TMwjzi/YxAHmpor
2bs1ySdngO/EYonpS3d83YXalEOHCoxc2j/m+EyewCdrXG69vFXurHNA96aLV0U8
QnoHWnRG8xiTSa8igPs6g+ZjEBYJHOryi3uP7Y18G15HQR/8JNyCRPDYXnKhn9o0
Lo8HY7TUyefeZD9jG2zDFapGx7fcj0ASgIvpqVXc3uMdyNVmd+J0Eje/nUuwWXNX
rBCmJS39KTc9sVJGDlzgzlmmYxyM0WkC2tiR0OYKycbwcttN7XseCVecMirNtsp4
jFtD0hmS+wF0hL9OE86Ai2rJYHdR0619E9tcRbXgY2le2P9bQhA9WLNrAwPUwi2B
CHIh65rN4nTLVDxf9SPMvjcgErabqIL+/+XJtUvwyI4jj9eNXks70VTlR0U/BG71
HUTIFq2h0Opf5ke8ElrerSds2Qa+IKeU/TRGNcOjPi9RPZ+nqWTHcq6pwPRf1C/b
zRHKVaK25NijGv8U/cgpH/cjqV0Y/WCoxqyrp+Y9ToaXIpii8jqZ9Yu9NZzsTOoS
Tjkd2hzdHnfyefypVCnWNEYPPBBqXaUmN0CCxtgoKqjfGJL7QkP3gFOju58ZxpBY
TqwIZDuNjykmG6nBQ5h64YKxTaN8rGrK989urivKcnRrNRX9p5GociOi3gpnHpaj
8YTZ0hATN5QFbnFYbBn+d7A7L4knfGHg792xqM08BqgcaKXJnQcy+TiT4LYE2e+D
Q/GIq9Cp6XSHp1MU8FGUqLDq0nq6GgwhiIs8YJhJ02zxzB61thx9FHHi39xZ3J3i
yh3GLkZUp/gb6ZpOG70Ch8SQ2jpk8t6KfwxhngdGFOlnnyC+b8Im5XldDBsKqG7Y
bq88wgJpK12qPISDJlPJ+yz7XJX9+4MbR3FqjRA+g4GXGVA5vQDDXHQc3dLHom7Y
lQvIulVnOHESVhug/XK6ckHeWIU7ywjQWQCGj/2NT3ZoFTLluwTkDf/Qma/sg2fL
dDUaOhBDRv9QeDwspbNq5DhRwBiKsMeHMe7ltVg+Cn31AhBvrjE6cjnskvvHEQVU
Lxe1NTkAsGyLsw5/Xiyw5xK4qjHiFZJ6RhSQ1XbbtJJLKFSGp+AuFvRpdCZx+cFE
oMrpOckFRBfAC7+B8HVKJRmGNQF/STGqo9/xIeNO0VmTDpLgoZj8qC3aPrugbeV2
4Ca8K4W7KOTKydw/j+RMhiBgiyE4yFXxhGI0/W0CWmgzQxoz47SvCeGWjUrLGmhA
Q15L1xJ7yfYUXmeDSj9glb0lg4cGQWXoE3IP15/15DhahNlvcUnZvP/pE7E3+3W2
sCb3XARouhkeEVajan3+TtihkKxJN+mr56EMsKLjr5Ga/ji1eoq+9bcvRtTTLcU7
WOG5fa9A0F6RsGFPMr4GuBIwl4HHWXXeC/jsW7KFB0JmXvePyOMPAMvenQVKw1DY
hKJsGKzDc9r4fENBabvQSfLxB1NTGLLhCVZJdFwpK5ndXu7kb5e8avSspBhlCeG7
/PEzGmjgLb2TbnGN0ZukiTX8KasjLuvU2OYPYsfej7Nw1lCwCVCzRiqmJ5fcJEW1
ZgYXufYxXhVxw6No+ynCeGLyhpCLCesi6jFSQLs3IxLbAGMBPycvwp2fTwWc77Eu
GTCbOsEomt6/Fk0HjV3uFFL7Bw0JIcnvbnxHLYcFUx4nVP6TPhEnNBpnnzK1eDDg
7eYXDnyRSC7tD3hlaA4Ck47Dwh92IPqcFsg07FF8WXCYwinIeXvF39isNCTFjxxb
4arBLQJYLwRB7okd7LlSc+kfhj8g3FzN9Q/DMzW4pKtCGjOVPbdIw53vii0MuVLJ
qRnTMvsKT+NlSjVK+3h3zcL3tc5OpEtMv+xLrbUFbQVtOXZiDNT23cRKUW5SuQ5C
IJRbVKXSsBhBs2TgYR+Zn6Tew3II3gqXjoM0n922p3LkM0jgXa74QRrkKVUPlU3s
84QTnjHh4XbigDiWXmXBQQbsliC4pPVSL2+KuI0mToJKzHCbMlxmWYjWF0sS7qqy
JXhrTtH9rp334t53g83l1FoyMS8SGRZmtTdZcuALFRQ3/Q5zbKYjErJocmaVrCFk
O1icS0kDnUWaKkKNpNpoJIu08qYHt8rOYMMy26sF2gon6x26jhATjX8VqFm+hfoV
pX2qTftza4MBNUgnUVvDuhpNUUzrKzeIpcenTCJPdrY9zKXg/WMKZnfg/ipm7dTx
7GolAz5lNK/WhP+nNvl6ZNPUMX6W/r8FL5FpeJLBMtUklPkOjQAUEb1RuXEf4tqx
AxdLJFIbzFxryVpHzZOW886d90FjNihjmz+YitrqJaCpIUtnR25p1rl1Pgi1TvM2
6w65CJujGXn5K9S6/dESq6HN2BgPbt+CbrjzqPUfUI8NmSeSOgWf3aKw1Cm0MIV3
6qJhf3i/LvS1nbqezTdpsnJqXP8fSFLTIKtciXTE7OgHj6UK1ckgqRKg7KCjX3Zb
Zx9tIUBi3kUzRLKgniHEyhHiplfPii7s5eidBhUA9+8Jxw5Y3fGKCu8peM/kgowP
EIoBlvR9YCs46ciioN10N2WiWCxUnG1tx4Ojh8fn0BHdEy788QXbFRHnRMJt0dij
sr8vq+zbWtnqeijAXRftqTAngjPsFGjJ25ejo0qyX+vEsLtV9xh8pjW90ql2+jBN
wdgWyKz2T+tvISgAOUHw9IrJgnMqBeQP9Qi02aL77sRfghZQYZK9HdYOmuSlx77k
l16FX9WJIzl7iTC76g62NsYqI2Oq7ex5HXtVWp38wwQssPX/AKwIiExlamqxYd4J
nyLxifMMenpQQqtsUMqcrxgThq/zMyrqQLPabY/PLQvHUuMGoc9+P+zKxUdAHrgY
cAfeiGfvnLAj2gE6PJg0Wqqi62oMu1HqN46hf/aZbSxuFuuXxrwprIbF2KUfnuzU
7lfzoLUPbxV987qsf2+BEgs1SecJ/X+Jp4ngFO9EofpLfOb7a2W8ELDPRxuG9Zqt
mEAsA+ECAe2MCAOueBLJYBZ/TvyiG9wupSz11FtqL+GaN/a7C9giZ6RULjBOu+gK
Zhf8hMZ+r97iJMzPFSs7DU5XQOAe0nO4ColB1vFQ26RsKY1OB5zYNb8grJQfarfW
+dd4fj6EYJ1IEhbqgSQgPoJRPUHZD9cX/MK6BDsNcTXp72J+CdzSMzPuDWCpyvN+
fx5rX2KCdVszQECNmfw3xZD0mnz/H0IdkI1hAdcBHcMtgxIXtE4ZvixhFTPLke6/
gAhoBkwu5qDgAw3cxD9MYkeRgDCUG8MDSYLEtQVaEuruupu1/zH/56E141bxgNRX
izJSHGjfJujsIoqZViV+0VoOzMgln0bHSj3IGU6BpYWR48Q4SKrtobp2aw525HAw
d2RDndoUTwzXoC5dPyucJBqBCsS/ts47wkfIB3lutLsL8tCkP2gAbVnZUNBi+EOn
7EHiv3RLpgLCiPzwluO7sTYq9rxrAw18gG8d10ANXKA1EFq2yGYmgdrkFv8XXUbt
JeUCEouJpjbqJnKQu9sbewXpjl6P6r3Bss8HtCxtNMPo8C15TT3q9ly/IcpmLMp/
QKIU5iJEjd0Or1tcSNEC+WcAjhaFqlT//O4gI/gfE4XqoH+sKIad5YXXo7MSj4CM
usYMHHqWxDQPuuVOKJ+qVX9XLJaa6nTLAEcxVKiyJ1PFIbVChQXli4AEq1C32lRh
FFZ75FZqE5gGpvXIE18oNFxKomQypyHt74krBkr4l3iynJ2f/g+4xO3AMUFP3pcF
HWeXk6eJ/UTqaL0sU/cSDL40Y8xeNAsfIaAInA3rvDmQ8uqf0BM95n3IuklqxJqj
OoJ/OWzMZZtRB4V2Trjfr8+oRwgQqMxYTAqRGqVaycCk42dk55DhD4zMLap4Nq68
DCoZoInbhXwXkw2sutyuhVfdG4NLPDPjzHQAs+Pn74qH99u4ZiY4RuSMxe1JNSAP
0SOCt0CEJl28p83Wpeu1lglTADX9/AGRE5FJWfpayjGUixng4NFRJG7ugHJA2kC2
oxhGn/wjfo3K/bCfO7BC34Ifnm611PWEPc1EnAbvdHlrXvrbwPIaFSVx8gBGoDSN
Owqt7f0sdcxXuEhvU9PTd79TiZhg4CW0wEqob8Me1MWw9LtzX4cFryWEIdDgYc9k
C9i2kOsUdzy+f+LWQHTyDEPXzUkbifnyO4TX1mwbY+2VAK7TcaHE+U04/BiAfTTg
flE1h/fQdqHX/KUKmXibbj96RJoNdxHU0PSvMy6fxIRyP+3fzVVzavv8Vwn+s5Dy
gX8EnAXkGUfJY8ujIp35MkzOj42/iJn3RjxPZCjfdvkiD7GBVhcXTfiXCbt/VHXb
a21Q6jHyAKZOGsdG7ib8PyWBZGWUaNo7qypcjY3ASKlr6CDlFJvaJrwuRcIAEC15
B+W382itMyPV7q+JaZeb632dBBGiQFd29uoTOYsD7R32hjMujMU4t/coYGS2F15a
g5RnY1ZfxQMbE9BORl5Kn+ZKKak9BoA0HunQZ0+1W2mIhE3dc1up9WF12fq/uZTd
+2LdcVniE35gQQStz8TrlDijKND4cEtNFzqnkiwdka4TdQHFEQZCSQn4XdZs+Zvn
nO4KSNPHS67apWM6jdlZcZrAS59alDfHyLBoaigGRnWFHxkKNcanqhkgDelrxT5e
LGGN8eoO3M4MMlXsetHpInCHnadY3cwSuW9W7GELqjl5M3X1PlKlJTOuhBLhnN+i
9xt5zVdA5znX1lZAKebn10UubE9mfEmDx0P2v+Zc0241beb+wjTczJr9es8wORnx
Z46KrViz8DjbRs/PyRN1OTuJhIfzYj8Z6eGHHLtPdDJUYagfDVmusGIEUrodQuRB
9zcCdW/7h3SG6sqF1E0D8kDRL/wvVfc49ddsuI4p8eDAZDXF2CkpvWJU+sVvoGbw
0nk3LLdcdBfdLeC4m3wXlYFoxVaoHco5+v5v1YlSTIN4WPmg8awJ75STsXp0Ap5f
ZiBQPNK3QREmd0IfpBYpz6yA3k/WHCuXsVMnsVHCUjwUFq6eNfeV+Yu+KaLO0FCw
Exz8P/k3YEqRv/JqAeux5c7W1bKsovQWzMCXDAwCGqVNYhSR9FM6N8FBQtWeqvie
k/Yqia2MLJPaV6rT6PYYTYEMVai9WluQk7CunyppdBdgbAtSd8BYh9lyQ6Tu9yXp
KOrJYirADm4xWP4E2l/nupU0EMgVtqqxsFfBh1duxJz6S/NQP2zzOyRv1DXVCcH+
hI/Y8bMoQ6GVGmXzQkRJdPjudHgshhI7o97uEDOeFtV3WV/w/VJozHBmJeoxDeNz
UvJfb93eyHnMq/4QxbZo/4bmKmRahOMmUcxuj+dJPB+f0KszqzX5V7SfittCXxcR
D6K6oRqnzxS13VrC9KAtdT44T4EYJrvdZ9AqM1amGGvDiKv9wszVeXKo9psFQBQ+
yWk1jyZ27HEmDuHE3NUBegz0lZEGqiXFGKcdAIJqdh1MkfOz1tQa08aOHnEAjvc3
P8xBotHZUiRay8hWHfyh/7UkXcgNEMc98yEUGbRwyxNmUHrgMKk8CkIR+nA0c0SG
m1BdgXsbgcyqXCFzVYHkO2MU6Ckwt0g0dU2lFlAjQ13JzHlKN97Kzltg2Yzn+8Ua
1RdzOp2RPdjE5H4WV6LMDmFVAHmhkWPF3bMMZbbIaN+rp/HuHMGwaabSRzG83N4W
ALQ+nQHpBw4+ERZgbdQOYuJ1419xZ6Lwow4mmpFpjaimffR28m0e2ONLQbqoqJY3
S5/CM68JLp3LjttV7l1DE2bnAD1cy7bORlmYoC03trEcYo1g9kGZFHfpTBi7JKvR
LVdhaVqYeuqTDxyNKW9UEd5JQutwdL9FFInPhr8BT6CdVX0BoUTIr+mUKStvN2Sh
MI0lxh2c9bqf2/KXXkRLaTw9tdtHIVedCFvUsg7wWESLBByVhQmajw6AmXWw+6b4
DaqlukFVXhdJPhvWG3Af2BmsDK35YXQvrlHMupgfPKdNR479LxnmWY6tPGlYWtR+
5KCZRyDX6fnp2qfUffVFggeyU2EFumXS16U7WLVc+YeTYLSU6CqZEDwgi94Xz/Ve
AaTY8UCmfliUrYHcJ1g3LXXm9WKLTXmP0hp1OAUmfCbPIM91YOa2wT8UiOzfi25S
QjuWamOMOgsPTuiywi+ApsbSX25bhnj5UI9nyT1Y68qUWzjOoX1r4VVee5OwD242
OQTgBYguhBQmIPMUwfbF/upaNOYItZMNXVTZBSjZ00a8eR2pl7wVxsbPHvIXyTdi
QFcbJro3egwNWMpTmNvFU7OSN7DleD+r1+n6nYm11+7X39wrW21GOBPf+lgIqlfi
qipw6DCUpOthkRVmGECz5IWLlh8MBbMUcaxY3+nBN6/6aUTcRVBX5vW5ntYCxDcg
8FU4QhcY/fujyRVNIHc4kWEA8MxDobqFmzss5ojQL8L1eJvbFltpiBvC1uruX7MV
tZ4Nco2oBHYbPndoP6Amd81AVQJsqlfF9a0FggCDDecJ0yS0A6TOeDo0AaaBX1Ui
F7VQ4HqlqZS33PQTqwE3RTVg6jiGxI5kLFNt4524kab7IaB6QQoB+YZ7KbLEMsTL
uvsa6LcswAOT5bFKPmOBmgZLvZZDIOuZx9pwlJbN6TwCdjgjxtCHiV4Hn+a4WUOc
SY/4TXZwJYva/3bkOm8288f7iCgMJj2+EziBm91c+OHsUT0sCUmnKdSr4fId1Zc+
hSu+ZAZUz+hH2ua6aBszy973CxRjA/kOFOFgfXOPhwCcCHcYeMQN4tVMzLKEtepx
HhTbRyY/srse91fEobTLT/mBAQ99OfixEcsbeAF7dQeTYtyxkqmfowbnFQPkiiGK
8bxXX2TgfkX9hjAiiCedRnz9l3jfStqnjKJfx+hgGok5oNcKqXz889BHlu+qiepX
0SQEyr1aAU8tPj3Q054LkFyrKH5/RM2WoD7Xjf3tCNrQf2aKs2vYhxnOXI8ZaJ59
s2VRz0TNQE9JsBikvnX6wEvAgxtBYIq31ujoacZAJj/8VDAboky+CcNiYjrYZbna
NruvWIcZGDbsEqvJdb+iCUutsZtMaa0erRS2+p9owzU83yK33Al6dgnqAx1EbATN
fl2eh4ZdA8MgloynJysGQ1UdqYZ/LSTUhuwH7tQXf+lLDqzlCjLEMpKUYEqbvqqR
pxF5e3Y1rCJB3HqYMC4JRKZgYrZ0yz5oObzoGkfyIM1JWiY35SeEXdthIvwV/mBO
IRHTL48JLO+/Sus43nIQJ+bntrEdsYd/pdughG5UYDW2hdhRPKK2shtv/hO62YIw
Tv9cOhHaoEbCzsWfQPmBjnVSe+tFyWEbq0ui8r46orp3Vwb9wxQUFQDtJ1tOmQOh
pOMqG+/BfuGlPm7YPwYOlhsyyXHSKsHAJTb63rzLRegqd5eXURLk6tMC6x8SEN9g
+9RS3F+nK7+omifqVUgh9Cp6HeltDaV6Iy9+HbW8U7SAxYHkx38kqsmHbtKihTpt
RDX6XwhPXEoQC8Ob1o1viyQ3GQsy2WIx91x3iUv28eqEEmI/Crzu6I6+TbLnM6+Z
Dm+cONQeqiFrNAmUpwuiYNMOPFAkPTyES+jCu/4pcRNTlmjpAHFp+BONXs6FLpIV
iuXANQSNqn0fBeiIsDFuh9VMetZZUvHozhp4odqzjlOwajqBVVOs/NZpfzc3+w/U
O/sZBHE/ZxxHsIjJRcMNVDvo/7rSMXvSYIYjt1IHEp2GCJM/aijynFwEjF55dgf8
Hm/panyRfl2RqsxWVq8fmCbwriU/ToL1rKvR5JLoyxIxzK3LU0FUgQrJt1Zyvlm6
1iw69jGngvBFP6OWf+uwT7BZTsRfs0P/Uyrw2qvHczSy5OtCml/NsquvcnnQEJnd
xElkGGgciMaglRR+DLb3mJyTkZgc8auvwh2RULIDEOteeuo56hZ2ZA1E3yLI9T8F
QlLODQma2h6UhXUzbsusHvMeHVyaTFj9OhQhzqcNzOVcMK5j5COU8cgASi+SlF8L
mtjAUyMFJCRkMB5JK3k9vi99mGOumZdpRqjVNbWmpVDMoZwsXfu/kzybDpx40BNC
CFJfwg/KGpk/DhINxVAnKWB1QnPzRPJXQ+7Bj+3KhfqL0j2MufphoiBhMJKtyiAy
jV7e6wwD8jcZdQE18eMSDKAaZgFal7u/pJSPZNNS2yUD+yZCrBPd+Ro1E41xWPBy
FCOpfLg4hgvcy3XhWTSaR5ugsiDt2gXTfK9UbsIFtX2NHS9KlLvFQ+5eQE7uLkwk
v9hrnWWnzAAdjJ23lwRPEx5dEOJOuMSSimiFlcOkywtobajjFouZtLNp+cXNToQ6
qlkiAR5uo2TVXeMVmjUw84trEerMcZCUXfcP+b7V5HnHqlNTZhBuNdPjXQoVmdZv
GeVrmPafl/xmZKyz1WXjfvjTM5xlNmhF0IREfiTjQw5cfZy1tarjlGvefqwfiZpn
OicbOK+A2U7GkfUVVZgO1P0eJgpB1wxwyTOehDvZQrVK+JMTy0ZPWvhUZqaDoSN2
gyXBLyeWLLZp5EyG9MjGA08M5X0R/AgSFqVhU90P2Qp5Cv50SAevRLWPUFXMWwVH
tg+F5VMy9JPs4xKXYO5PmFnfAs+AfVWkTseKSNzahZzkLw4eWyxPCxvwSyt34ZLV
U2Qnt5/92bU4AZXNsdWvRuqbGErApTPd0s4YBgGwClLeD/8aPu8sdPlCNQHTl4Em
Rd33LDNz6yJjlyYN6rwjaB9rRdnqOD2trJiE6rSGsxL7+ORVAu6dd9sX1WXtv5MX
NGp17X90KLHEMpCshT5lKl6kRglN2dxD3nC86QYl9qsEAtFjP8jBCp5kinHChxrv
rV6rnxrLuDpMSIZCpQf298SsU5SsVB3grefMXI6J/XX66kKq1OOeghvVb7S1jD/e
xII89Ngt1AbXfkidwWd08wFWiQxFIzsK/NwGaYIeK5b1BO7c9mnB7vTYv6XrucqN
Pc7MIXt4tEIMH4DkAMAzoKvMnABt0+PgJOS/9oPzbN5kT+7tDMglWAB7keGMSbSN
iLJZjwYgpja9urNp7pVoH7LLaaRP2PdZJTyMo78fzywidmpapa/mx5BV7w+QDocd
WdC3oqQCreY2JgNbNdccUuioUuik1zTjAy26DiU9XS/CsdDyR765hCpjxgNwYrZZ
9GfiyiOVP96Yr6P7OYtRaPhFUgVH/nfLK/p80ZYm3OHEIhGJSTyZEge+iD+HiSZ6
7fhb901J6la4c/n7R/qrdISnCTGTET1+GpiMBm0KbZ93q8MkWN236YER4UICxkMi
LwDNFIZz+Fr9LDkucs4nEXjYDoYhkG5mNhNlXHe+4Y+k7VE+etGXYF3jyqFEdehy
qZdWh5hLFc+iCXcCICYjLiUoU8/2mvYC8Z4Vf8DVvr7cJVGN21aDm+pSGuFVs1gM
O12u6ep/LoryHELGGQSUBBDoZamjhrw2A5xIsz5yoL0dfrxnbsMGB+GJPhouBRx7
Ic8fjnTt7szEsS2Dz3NiFaZsLonLy8Ls2sTSjIkZPXeTJzEWBM8esDP0dx5kGaYA
aSCodmzcy/XvGkBVbs21yMhe833lVxGmLadU4c8bbFVUjomCKVITMH3NyMkxcJHC
9bivVmQmJsApiuwOLqNtqTBtjLUA5Y8MTUBgIy60ZD3+m0t6JvM1wLj34+tcUWJn
V6EJ1XkSfiOliY1cuc8Ft0qFSI0TfeCqW2Lor3VYe9i+OzSsiJfPI8hrf6q27rsR
xdkOzCZG0jQ3MLJ3y744fuk/OvedBxV4P67PAQXAfGKoHHi7uPqcDttuI52kUU03
a3WG3xdKy/d183dQj6IKON28bRODvWLfcvIkSzBEQwN4kwwerqPl6uPVal48+pBZ
bYueAHSHC0sPxjrciF5bR/h9qoxJrhQefcJASGn/wnsUrDvTYbOA5KNEYHmY4YPA
sPhYx3IzkJlh4jsd86lNDX3jaY0wIz2Y3EpHwcOJtya8diVymoUphheg/MyN/9O1
g0COPcUlHpaAp4HpWz2Q0ag3z0stcvuFaR3wena4U/0SeLiikxcunTYe4g+rP8ih
33YAlElnU1ZK5pzqFDW6OPrexATIMtpBuoKATMLLneIj7nMK8yCisGmfLUwZfNMS
DTgGD8EXDyVyv+J9nNGp9v5DRqWk+hD8FADWIEszrT53pmecnefqYNnrE7ovbm+V
JCXm19bVQb8r959Z2fQ5EirmGiZcORLgtv5ydbyN83gTgmI/TuzZ21tghKwB0PW1
p9uKOXYx5YsgnZjrAfFbYzQSitl+xMVfyTYSseVfgztUftBAzu9lYSGEgT/ByBw3
qErL7pciYktzdIzkj4Nuc18sDlrNiLWtXMaQh0A+QAQDkTKPwQ6kX4UwAZHJuvCC
ygW28wNbUajFQ416ZQh7Oi3eV1A6NHgmfjwTU7bsI1WuWAQ2I5C9bUfBYxyoxB90
vCIQ3iIitMmztF7/zy3PfHviuQC6hEAQhFciwxdOB6NvmuMyASsNXhpn5CPKdzKN
DYC44Z/A1UhaX03vg9PkglUQFQpmXNlCqxsKsMr7/1tFSq/LC19XhdDxjHiK9lEG
AybpBaw304cYoBqWu+ivj65Gqf01i60ua4LDEe1qhhlC1MaVr0izafo9ifI08h7B
x3hSYdkWZhSTEoCHakOOKfvjVOXxnQipU0iqrXzywPh69oTePtUrbLNj758l509J
kiEDYn4WySSm44oSeVFP1/IwqlAw0SlakICLwcTMCeWYqWTIqP7pnM0gtlsoaNp5
eQ7oGTN2y4/osAwGfqw3iRogHPpFDO3Movhk9LDYAmYQL+WyWZBK4JJAY6yqQDXs
bUbTbQjMwbt6wCQrm/91L8A0utHOvoEhztDCDrZB8Tns9TLHxxpNM95K3W1NjYkK
8qeGy4HtYZSm+f6xgQNS63GrWbMnuHFQMXPNnVy4aY2QCfTpVXibTlre/TycZQos
Gd8K94qJo+hKjf7u28YYF8k42xwVlr6Bm4Hyn79DzHBtcdvrnOai6Oy7QR9jldWk
t1nGZnplVvbTCD7F2cs3HL7LvI4IEBlkdVyxgTUz2FwtMD3B6KPVQV5/1si7DeMt
bTM7cUuuNu4v1bzC/p51YluUBW8NiJsjY4J6HbEFCQvZgL87ezdN7KC7Fi/0Gphv
ToEmouNVQHQPjV+2IBQXlmo13VhgmBmaYowUb0fFD7WzclSLQs6raCJ2wmfuxirZ
CZaD9QQWsiIFqhmg58+K/C9H7e8taF32iD7toRARd4vxHwys0b2rkkkC9wTjv/8D
zej8iPc4+PxqemZuJELhjk7FKsoekRQVBDQx+ZUVeCJDad6WI8WSe8NeYkgl1sXc
/6Ystm3ZYItABM20Pj+GRY6wiFVFLsio/fVJBtR6JOzK62HwS4HAuIV+FZMaS9Rc
65iRMucduNZjIRvV6x+8iQk9L1iJNKW/0H7nggFFO/2/B+OPKTbnT0KAPxlcrrko
7V0pD93VHM7GF5yUwttucR+YWto4osxyUcbWm9H3TIxwc1l9Fd5MbNdC/9CDJpyB
8xnL11SmUU5ThCOMKIyVcv/zNiwCrR/ld9oygjJb/eJUYFptZBrjc0nadat0GVPo
6M/rfmU90LCeAlZYbwlAiJAFrBhmXLSZ3sOezcZ6NWnxPVjxL9MuBpc20U+a5X6y
Y+4FovQiSIH06rqTa3BTDP87rDmAQzaSC710SHTg1pNpJK0JF1YzuFnwRgWTaWkx
b6lfhacvADkzMG5H2+qvisNEpBErlbo2HIP4jUZPAdaEbFKTsjVx7wf5bM34Wsg8
cnRRmTwgXkru17boYOq6VchwdWgLdVYWju9q7TCsIHWLGSMDZEssy6zSxPf9JhbW
0mJJRkIGhT+9G8Nas23e811otAAHlPVfEuMtYTG4fjNgbbgCwwkaB9F9oo7YqCxn
Ki8jkntL6N37ikbPpWmwApKJ1W2YO4Pa7mZ3UgHDrSROBcb4GjVFpXzXt1/8uH73
AIVmeFWcJn04Z/BoEnkbhquD34n40OBH2mkPJW0YFwfuyxb6laruAa9s5FEQb1+D
cxqG6kyjzplz2uC4NTV6nzu2Ic+09qsHSGlmnMa9wohV6i1mnFIiZxjhZ4zOQg6x
5iIKpEmW5miWCSrIlku4xPsLPaw3xtDdKdQ/NoMsHAUbHRr9P2UIm7qGTmUZbQ1Y
9pcw20yb7YHQta2XgbfNDxNJwDVHIvr5OJL+QdyI5zliLGubkcWYcPZ69wwhWodY
/aE6wRNi2dtlieEghrvvAwTaFa8pdNB90QV53R1RkB6vDv8jkLOPefEfsm8lE7u/
r3vcv3kiloKQR171VVCRjHMR0mSCmX9FYiK+ZsMmoD9PSQ9uhhFg0AbCwXMpcOLC
ybWPL/J/N3aVTinvjDUZZmmvv1L5WwpRbftcPOFA5zl8njGwAT2gGvP+kGQ+5OKo
N/KXSIpx3lu6+/G+0aCrdxNoUlUQXnf1hc3N1zobCv9wAJzNbV8EaWGw9v2YkJNk
0rvkWKBALgGts9lN2DkbDwK2gaa3Kdj/I42c5JoAdZ4viS799qj1oGSTW5cw9HH5
I54CBfSiJF0RZy+baS5IWx0eyDlFNQs0nREuamPyTxaHtCVnICHrS46u9vLeEBBw
i8XM92Yzq8Aj+PV13aybj7URpFlwJ0U3p4Q5//jgtmIPXD+4kzUg9e9l+UM18GJE
busHV/TmYKm1M5a3A7vZgHDwRWQ6kF+wgQLZper2O39fEdNQE4zGHFEfYtWk0DL9
V3tLy7RKJCwCSZF+o0HJmb41sLfANDlgtJOTFuomMUT6zXFrM20YtpKJAF1DG7BO
Zlw4Hpm+ZymZ4kOdrFTXeBUnajScguZugFy72dF6/eSDbYhVX2KugWnFYjXcJJ8y
6q/4LjsMwM5VoA5HxshdxXkaeXGi/2ELcLPhViQ4v6BZt0CUdSx8CzFSpHU1so9u
x06be8HjBcaVbIhkkD9NjZZNCoB42ZMYBFbpX7bflfv+Ph5DUV+hh29rZW/V5V9t
FXJyp+x+Hl5LrmonR3Q6HlIawuCBiBEuVSOlK8+2S905c6Z/byCkEtFxDjX6EKB0
jfDzik4g5UmAFSWXTdPa3xbO/Q8YULd4kJaxoKoIG9hVnsdNOIs726Ud61aGpnPe
KYcLsfEQItxXVsjvf1dgvJCcN5Y+ZHY1t0+M35YVAuJSu9rV+3k8SdoK8aEi/UAT
ziCTxmjUuMay9kNVtIdXOKRh2bvv/y6bb88x1DrL6ms5cjbQiPJ+9566+xoyMiHC
sIE4ceenIbvzkguUkmZfAwMsTL6quc6QzB2XzJ90D64OWBkxJjson4GxF8uRqbk1
RYn6HT0omEixUKkXgwwCIpStRR8v3sF5DHc+j8S1E4aiPdrbWVWb8erAx4WfW/8f
/qeTVVEgQkGJ3enCEpkbl35CPUIrLMfWcb4TRLRVceMpERgvHwJfhE4h+sqjMzJy
kpnVFTZvFaREix5Y5kHDPaUj8FI+bH2Vq+zrGaNv01T0apDfO9ycCN4kHP/WoGJC
dpp7A8IQ90ShKxwsIaJdfvqWqAjxvCDYd3TQmWc6ex/KQSiRaB6/fqcCvbPPHaR4
g0LJpmJoAukW7HqIC9g/dbTBsvd7EoKlSJxV1roXcvjZOPIiUHQXio3gxHKh6yzk
9QCp42e1nqYRrhef0ipJolq/xt+1DV1JREkNL160H+SpclvAbaobuFpaz3EBrG5k
XfeQnJxOuL3MOIYnTXQrPJPs3O+BLmzbHaPZ0RryWqPJVmE8QJ3y0sEnUoCLghM+
S2aGLzav+W+flSjR2EuDHOAMLAyqDjjbNssBzoiM5Ppn+6Hli6OsIqUF0WVaYecT
X6NXiB+2XXrVHFYFwoz2kmX2oFMgLTvMhfAkhiZwkyPF/VZ9C9l7UFpxsRDknSpp
ZHKJzphMa9VmVX085TP2JJE2s41oUBL6ORYm/EcWdpwkfpdbfO1QonLzoY8oVFYr
ojcd8FPqcinXuHggcRZtKa1WVAZTzqPoq6vO2QE37Vbln9mYMUvSe1TFWZjVK7wM
Lhux9Mi4Asi7AqaxG9q+DwMacGypwtacBLmHG8+viBFyKOrTAvmsKjnvONYlH2ZK
3u3hIMgTh/DB3vddJKDanQ6S4O0I2WGzVrRPO0PWYRDhwkvkgXSkwBFvQyTzpx9T
xOiNN7eyMLkVwlkGMuFtn0P7XOi/z/2hmi9q+eKfafImrDGF6KTtk6oggwv29AgU
k+hERvc5v7xInXy0rAe18++UoETvUFghYgnlwKnu4bO3ASC30rX/tBaGIsWlwDw3
c044FQfYiNF6d/e1CZVOKjzTgTBqRSqWbRnBfd+8pkgV34YchLkvdK0b2dwY0tM0
JwGCWQjaNx7Iw59EN3FyhtD1hK+rJu1h8JK/sGSR3yUirZqkY/NiqjHt5djZA2+C
vBbEhG1st7EiS3Ry4d4XoKx+SUfi45jUfRbpozJJs8K4wRt1A9G0kLVWpADm1mL8
xe3xkq5+9FoQ0gLB/BwlU76/uu9ErSoV5Bsvk8m07cRsiIaSR055IiR/hU0ibQFo
TtKwS+kcjat5W5CjnIwK+sSCtlsLSieoXDZjfNfUsfzO/0dH4TzvZSBsd4w+/O+X
cL3+NdixbTBjnyMMfAiSUGTARdTo+yi5IvO2TmZuj1IGFtPD6vVE3aCfUOIjEB2B
Dwtmu4K1B0qBU8zSYcGj9yC4BP/EqowF8YXFSZuYEp4a8+z+hKZMQtKmzLQcCy4Y
GBPUY89E4MfC4XdZ/xeGnJ1xDUmZ6JdgU3n94gSn9tc3LO203Enf/oo+l7V5w6HI
MskqEgkCnzVKgONFHSa66jslWdvTQoiW2KoCflpG+oPrWaC8dQwFc7cCvr3WVbXh
2nFr8nvJSdBP6bGxZL15t7EQCwiRGfXH8uf0yqetbZUhr3rgT+2lo7O5Q+7rf2lw
kgigGHEhsTEygC8q14jjc4/U5vtUAqGEOEVM0xYqVfYmBmPFyQbsq9m7MMiY5oAr
GWaiOrngCbNvQ3eH562pRV1WHnAt1qCVxYeuUMV7Cbo79ZUOqFoXfnNmi5lgR6Hm
7c0MWStx4A60jcrCv9Xw96FAuKeTTZC/HnlGUZ1Njs4Cl0km6Ky3msBZ+MirLAYd
w/Oe+LptGt5uSDCrmPnN7chYkONrcrgqiGSBX6OEFpOBQW8KzuedYPZubzFsd0/e
c5wLycTWSb4ACJdsiXG2YNSFUmwad6SshUycgSgT+mPUY9LFVEyAQQZWUxZWGkJr
s8vTd4fzDJOwt3m1r5Y1ZDpm9ER/cVxhTkaggLZlX976y1CMorJE2oUCJ652K3k7
CbU+GETMwjySWGxjDc3wClLgTAlrfQpL2FnEuRwHCQJdGFLoL3eEEynfQXMSrvr8
i535hgKEjibG6xOYiNTBpoWYucLVK+qz0XWnN3wLHBaZxXjTlFHZytlu4IhLsUEi
ORd8sYV5hxkM3RiWU0KruNd9iMsn2u/YkeX9rLRHRr0P4oSiQ87UwuOodJUKTh7w
H21M6VtgumXk8h5P6LU19oHfoTcFi790R6RKgvmBi9DR8Du2/7dprVPmot7T3jhE
keLpEkvKVnk+DXCJIDvMV9IO+zZ00w1gT2YPc+mwsHCGJifhEYRmAbvt10pzTnYj
WrXB25AK7kmsENfomWvFaf3GCfI7Cma3FoFHZ6kQrdOeh8/JTDGFF1JPrytzVH2L
+75gg1Tyx443PcPfghnEUsl0NTMukeCRa2QSLdySB0ERhQl3t/CbtgrFUQjuEnnP
/NuX7BqKfWwoSxWIereTvimDPDRb3qk9dYspjjW1vk53eZfSK0L63S5dmCACo21A
ICfDSZBDaMPpfpAC10omGyrRhqKbj5w/SpHjDAXquEUXwuIUvVDWTtT0l99/Isab
UZ7oEvXVZnMXjiu8qvvga7eQjzeQOFfRFY9mTurhfavvpcPAcSOghq44AkpU5PW4
nWwUf63j/r6yBM5oj1z+Cu992H+b15Mxy9uY+JTXIYLM+WZRdLyl9wIdHVvBMTkv
7dkHM6gYCpbnjCx1IEJ9agYOh6k5UpDmo7tREjIWIf1c3bh3/xa5iTkzlAUf0Sn1
FDwEImYArDIEJWCJ/2G9NyApYhyntqnxs8I7l4KDognwqiVNRsxhUSQ5hJaclbq1
9rDJuGX50051W9Zv13rt69fDr2FgPsBYTr/3zY+rThJW/GGg3S/WCbLVL0lrIrbg
kSWlWnUcg63leI/SL3J5VLSVA0+iB/9KNwGqXGrWDznV8BgwV/3UoEJ5Pava7iAj
kJ1lpipfYGeKJkibNSLVN0/5DNLLMbAzZC04mEKDrJ3FWGGGboVLV8HU7uIbFN/x
cQxTUc6jdA2esqLNpqHnFgEPcGIuR1I+mqlZiMRIzTIIchN1MjYYeRONbOy6jH3T
RsJGbgL4OBpFJ0HCQyJBk9P0ugrzcdweVrDpvdiNZAjFP2KpWDA8EzdvoTKpShyk
4JKujdfV+QqV572F51u5408Ihcf6qMEbgYHghAgMdftiJHEm4pafJMNvB2Lx0KqG
w6nJ5G8pXPOFB0RWNGliZPioA8r+RsIpbCE9iM2SJBCEYid1iSPKaL+eWO1o7hZf
ZwePBUfqQOGsNKxtq1FH8puaXGcz7ZUNBnFEAzjYSm3rrDa9MCWPloNG3haENujY
GvZru64PTuoDyDgVpB/N0CxP1aLbPdxaDub0GjPZPvIs0RettQaOsnyloyQYzfXQ
4zztfkznhq2EsjCOpC00wcDWChRMgxnBzEP/0/ufuIoRoDqgM+zQgggk/+EnFxfd
87iWMiNDF2M4tmUVOICAANewGZe9ei2sZxN7yJ6P5qQWcODQQdibEAG9XSOOSvUr
5Y7s8og5qYaEFPMhYE2TZrk9ZzoOzLOzXG6rqz7iBF80gQ/hPGw1qwN34WcaA6bo
BpmJ6Tr3/YQN7dTmZrTzEyCZvSQ0U3RUwZmZ92cP0BW6mpwvhVlhGUx/Js1xP62P
MXYno809ddS/6GPenum2e8XcVCV9ZR/OaPABxnyzQj90GulWDnqoU2esHKla5ZEL
6s0XKzRErJj1cVYSaJUEmrbEu9bB+za4chRcN6Udbcgf6szbVQdxfPoUtV0kivQj
YhCzg0WKrth6pIwTe+7wEpLoUXXcGEqKJq8bar5IfjAvL4iLThjCp/q1jOru3brq
anq4US86jChKoFMjFDaK6grHWdYjp0UbhnqitzBBYu1rpAFiFTXOZxXyWeDTtsA3
SxfU4xOntsZgcoupDjx9akBPtO4RrBUXqPjWDzmORW5mjzt26Nk7lWDqBUuKBStI
KzpE+nmYV6UqYY1m7+A3yg66idPNK6gP0RLVzIFigN+JZitiCZ4PyIXJeZdGfe+c
SQybrTocXYeZ5yupwbulaBxQeUWKtG+1VRGA08WrsigV6CSu71OKbmTmHyM27nAk
cg08gnmYHkJm5+qwR4Zgz9xE6HkpomMd3HI3XvuuOYnkgxC0sv7GwLh9I7qgF/oJ
cGoNCl6tBpHMNAwo/05H5uKoiMaPfSFtqfW7+YPhWstHhaskPRh0zh6PVx/mBEmf
tyy0hdkd9nbVm2lwhSQqx0N+5aCOxx8K8iEViyUn9TVmHTNivDOox2PmuufPgLw7
iMSWOHFvSHco3/teuxGO/mGYBiXWrKEn6EEi/23AMCijzCC9s8qCVslQb9TKOQ0c
bwO0Updd0vSzAsLb6R4wzlv6DmZ1HbvJKO3Qo9VXleMi9G6He4YVp47ZzgBMxUg1
o53M1jbDV0nsEM70pJD5XkkivTtDR2WRdQpmAG8P30/XefVrISnQ1cVVTVMFpDHy
rvvF+SW1Ij0rmILn7TFx7K/fnWhIdDFB75k2XKG1tXtCeTAiLL0kCGm+kCftKtaQ
qae0RknjxFFzm10LhCY9yciRSlm7Uo+QOqof4sTRFM5lio31s+dG9Z21dNawZsnf
rwTJvhG3XZ8aj6t8RmYQeJivQ+yGwKKLEtm710WLOIsyi+fgzMzjyM1kMbbUYG2a
h/UokbQ15BfrEAg3Bg5eWYK+sXFkULdh6bXV8DX7FntmH60gUKMBrKo9USbYtJmH
S6fS/JfQSPxhWNVWthtgl9vuO3L6JnoLFg7rMOrVDxxwNgUkApHEPgpabzNX1UyL
jzTWbSewMb4oNhNhcpb7F01xtNGBaa1LhXzf2o1dVyumSF3v0nQbbrLWBzwDLXPR
OZ0EcxdbMwDS7wVoJ8Lr5tCYJenusISCXLJitMIoqKmWAoDfCBrEgfdmV4EjyWrv
GM28vDAStoyGayMuAE4vAYRLsLVHB1QcG92uhEimiZz+HmFVZv0ktiqbCeFQsclX
Tql5jpMbMWWDiPNSWc/CkPuWTEVoq5cxrYDVFTdMJTvUM0IdUcUtHqwsoWCWG8sk
3L7LqzSNbNsKBGpVwRW8zMmEDNJ/uoeWD0QL3SZQpny5gV1XSKwuFK4KUjU81CEA
00TCaHBdLn+7QI0pJ2jzQGCc3mVelU2z8O4PzVqM/52j4IJwhNIhnIPs/5pZb/dc
SyQ6h/DnmtfOJv1M5yfuelW6jwZciadkcbf0mr0mxkZtrw3fVW0sdjNQW1tIh93J
AeNU7FCzZTsOb5UXO8d2dhFy+QLp3QViKqAZkMUCtH1Q9Gagbuip6YI0dUy4TZeN
hjy2FIRWD3PxBC+Lvtgj+i6mC7v7S7qh2V+4svWFybF5KBKo9flOLC/4I3Mp/MAa
6DGdT7czvhZvZziXBHLVBPniIkr+cUXfxTi/7aRRP+DQsaqdfDeOckkFPHrtlS04
SOmpaOM0IG9OCKzsSR+S7Gx9yYW6o0c3JF9SALPqw3D9QuVPOtmjzxrXIQlUaOnk
m2NqTzzW8DJyEffANlS9qmzkIdDr/YVuE05R1JKalJypYVR2NoJNoolVVtmnhP8M
xwlHSCuuSlHY9Kv/SlfamBOmMB0yH4xQyFwEkjYxLcgCkUfA4uAPTYKFS5j7v6YW
Vvtfwcyi8DV2vBcmk3cZoJsQuedg/5k5MepbBABGxBF6ilrHI4dG1SFGk1ybzEn4
AdOsV2PA5NJClBVY6/83lQC//Ib5Q8gPyd3hVOOnqDFQYBpZ19tMkFMk6iknOHue
eAYI/Oc18GbGd8dgM+HCKQ2fNDj4b6RhzVb8eYbu6JleOJDzrXbQlGsTdPYB8taG
Zmmd8FpPLAtsWtEcPgaOCUZmjwGvUE9FBo+QovZEWUcwkXOTHyQNg7BD28qAEnnj
S+BpKGVW6r6jY5cNS/7DTAVYTYpY3m2UbirVLGIomruE2WLMSWbGDPoTdgBfqIih
yUGng9Tbrwop5bW9qkWy5MBD1SF1gIhSGoZCaHRsxJXoZb5lbQOM2u+wEZW0IXTe
Fpo9CMyqnVDPevJMM+ZjEJ56dW6TlCkQN8BT7XLdspI3xIybOsYUzYsgx1S3f0dl
g0I9MprOdoQKG6+JOFDkShcwFXOIXz9rBb12ey5H6T/09+zZpN+RnT7rHP4usaF3
k3HfwKZQWPHAuuTnr9xcRTrMQowUhd7N5QVJhK5Mt7vjjzsMvbDRoLo3OvcFP/IN
a88F+hKLCvFdLmSZd2GEpazGQERWTnLd86s9rgIqE1XffzuvpEwcmsfs6+Lxi3jQ
awF0nYyuiCrkRBTB1ltEtEkgHKTApUtjXNEnhNmLCdGGj0IBgJPl9o8GsaZbYSUU
RPyc6mZbwKOW9ki2tEvz0Tb5ZmbCY5SJIFOaIMsLNwQJ400jqW+XTZMd9hxaf/4+
1Q9ZPjR6SR3WYejgQaiDlnji8rZoJQPO0l1m+PFk6M6RPWYk0FSyUZ+viICRXOkE
nzhXH6+3gUTdl/8MJcxuEPZeganULI1+XhXOK4nbOPWs0kCNqGrRnKru/84HGMub
j94H4lXLu5IMuJLlE+7A/llEkOJm6s/uYNdwO6gY3P7DYsuhgZ3iNsNcnWZ1SEpd
1y0cJD8pHJPVPmK5bUb3VyRz22SXf8Upkmu4IVbDCWMrlqsOIOn/4uNa48qPsYGY
A0pACchuFIMyBu67MP83wZY5nhTN09WwggxvwAV5/X7saxVFuZ5R+DTATIoL4Xs2
AU4wDyAwb3xYH97sEXG2/Le47UOjKSzMTU4SZQwZ3att1M2jZakbbZqhEYCKpLel
ONyLr7OC+BhRMQDHlUarZ0ockIpYVuS9DYWohdMOnnoSdwjasJbSxnPBASwSTNGk
sVBy4sqN+vNewJkdP8pHGiUbLkq4mKY/YgqFzsUU4JdZQa4f2eikuHNrMFhqk22f
dA3mFJT7LS7FBIJBtgA8FROxP1iEFTaWrpTQkqSA9mcFJBDAoixhvMpWrGDqN2cb
VEKK2gRQRJbxKH8+GJe9MneCLjDvrgGR9oxJlRYqTfT0s4ATJ6A6bNmVs+w+I8Sh
V8LiRJD7RMwdck9CULSJpcGg7nqZwECAIcj5TePpi+D2bOdNF8zbh0z25eUbyfHo
7rr58zTJdO3Azdjs98sINeWMKjPNg2AEL8B3D3GaEHzgu+LSLZGO9phKL2zji/1u
l6uZ1LOIbUUqiw+TGr98tFnOQTnAioVZjJzTRxASsZZFJ/BGfMTXxwcJVUDFbm4n
rL45uHDsKUb+fnGhcXFjJLkvc18M4wCREhxrf5LZKoYSOjGu1lCUTL65YetHaHAZ
JD0h34thN5q19Ms+AkkdwuFxf9S5IIPygEIoW20dEUlFdKiRkYFF2nci2UPjePCn
HZ4mdo/OY4UsCugfjRiy0/OwLxtD5Rae0Xisf2tyaw73N90KKtS5QEn3RSUxPu9w
U7rM5BhjDPPqvvb1DhPxBr9vbU5kaLFfVIZTfOtgClvPgJidhvChLsM1SiMYXgGc
pLjYRnbUpuYzxZwRKMXbUVZoEc23rJm8CUbandUo6+REHvg5JCoViTzo/6RZIbGg
fyZ3C2BcgOKIi7Ek1u5aTdl5+fUhMzrdL9GN5gvO6Ej4DoIyriFlUdFpR2g+zNM4
cUb7SdOVgssx7CNFAdUAsOffUbKBwQIPuO1IuV/YY/tywBdP2ZmNUIRyZWSdMV4k
/+YFjOVykDBArnnhQuxaWzwmu1NvO1++Zj/nHYMQM43hHMWnY01+NcKRuCHjwJf+
RyvCXRcMWIgh1oh5vmHO1E20DUlp6L5N3VmxiR7XZjVZQi9X0VVRyL/PN9dPkl6C
SRcE9lSGuRcXlc3ZDBkk+aMKxzJ/FWTXBH4TDuIgs2GBJXKYLS2PXRLi1NRhmvjX
TB2aop+YoW9tWFIHU3T22Mi2U8q2UnQOCM/YICgei5nsTxtHotsMFfvZiSjqcClq
W0GZROCJU3MbB109KuTF80S1d7EOJfEkOYIcBaj0CFx/B4gZCIHlVQj9dpItK0v6
oAFNyX02xy/MH8pZjbvhWbZUzeoTRcrg7zIMIPPrNeXyFfyocOF1EnPyAI8j6Ljz
BjW8N4CDITUW39Nzr0hx1h1MMOmJVjRacyMxgdNV6mQSVPHRPraObDKxqGOfiMmH
ygZjCOvWbnoKTfi6VTHKNWUETs5beHGO6riO0TJqrB+tvmciiX8dxIrHwM8YQD9X
ffaqTZMAnlD+VE18OPSALQo8ratqEebOJWBx+3yZNIjXJc82MBPGXGigxO9KoDjI
t2ozu0//mgYyqdKciA3E8SF/QnIEUb2jKb2ONspTq4osSEf+2QDlrzOpsYF/zFZR
p4NAqc9r4SLKalZR65r9FjQif5PbQ5LS1f6wl5zWv3K4gIRi6JFRHWjAvt94L4sv
LMWuKTguW2w2PU4MCjpCjVn9tREYloFVqgkXDJhUbm0TSFGA2GRFu41SLQURwmSC
NzBBcg5K/bzanhQf1OnSh63G5mJLs/RFZHKrm5bz2wugCygUZ6gPc6s9RqkInuUG
LfBzmI6AQ0w1iF1PBmbq1SWBz6QbmH4hv2dCe5y/hWaremRHcgiU5FCWnrYkx8aO
0xdj7txi9ZNap5HiN77XN3i9v2mrBaDdTcHENNGUCmTtRZhZgB31DuoF6/AaMb38
XMwISwH06WaO13QAV6KFzEzqEO5amCKEZKSlZewC12Yu+XGRW3gFcMhvjzRqpigE
dt2XmxpSyR9juXAjHYzjv/T7VzjbiIr1WNwUy3xNKFtsZoPA4dKcq9VJUoyLDZvQ
5Qx+eLZfs0P5lFXLXlVyZgXf7oF9IYyAfEWRKcqDCjxl/xzH2A/TRoEoRmZoTM+h
93zCmBm734+WingVyfo+VE21xhWoNfMs4p4xtM99gTOoC2f7+0b2DukGF0ubrXVq
nj0XD2S9E9oqfWHV3Pyb3sEWQG5vNZGE5zU7g87mIVM9rcmGrNiU8UiwQKimZXsC
g6r8auSJq5YMHGysoGld6JRP2NBarxtesCfMPLjPMpwq6aE8jBoH70XfTL70znG0
7BohVsADV9V38Mjn0uYXBeGhW3Ybb1gACLUiQZooV4e5Ujt3hC9eqdcCiKhJyakc
/mMNG7c4DNge7hpp1I1CCvC85S5hyZ6VI0OduGjuEn5Ol1XYjaioEbpML1ujFYcl
3WEYg4hF1HfZdoyXj1kDBIrj1tpeZ3w05G8jsvqgGSAW/lqQrs+5Bd5ZZCxA/4Wn
qSuvkR4HpdzNGnBaG+1qtd+Xxutbp+GDdakMEGqMChUYw8QWBEbHMBlQokdYiReV
gyTTdpLCQPcuXn2Vfsb7ERCb+h62cZwyfHEYmkWiBKruChbYb8b0MK653Fk7Y70w
MILiDx9QrevVswC4qj53uggcQ9EW1cxjDjbqH+hPAnsIU6TnnPgW9nNKf+MCTKxc
YkGMlASG+T6XFRBV3GIJh4B85K4FFsaU9SDEi6kcLs/0VILRUTo94FViPtqgPTxF
dR9bjTTlSavSS3creJjB4Iq5RqYbDwjAagHFJ1tixaXPOjHbFBwW5NjQUrjAa8dk
7dCN8b8nmsjKsBJqqjXq3pPO2Ku7znN9cKtjGV68sk8zuj6PHtj3RjtOPnbjb9H2
i8o92rDsH4qf3tkejJlU7N5klECwBqjWjQ0dQbUpJKxmI4HvZxi/5a5CQuMF0YNj
2UBnhyHkC1A+FHH0XmYBwp8/0A8BwtPSifh2P+SDngnoOH/XksVgWqu8ZDExRzTf
QVanGNI5N0vZOOELRCIb13C6z7Lk27jyqWAhzPBdDk0HaOdiuw1hpGrVb79NFj0x
lPnpIMHOMWOlGjj1gOaVaVo8BMAhSySFp3CjRWrJrwB9ncymrMMfi5bCdCLcN4s1
d4hcEC4P9Ds3M8JantSVeyrdIASGbi+skDERf/shjD9dl6diz1yFoFApVYvxz/J2
1cGsoCUZGuL4mqY9TnDm+hSRPEKdmg1GUJ02lxnHUcVYZx2HI1an5Qf7HrCMbThL
dCbA3c9qTTESLiZI2JA6+qhE6BZD4qd0uwuJ+GLpJSHgHcyjaSjhfMpALp8vXo4f
2iNnk3tMVW9bPBcYUry3MY4EcB8cb96uYXLKfpIs16PPo68o0EoOyddxz5F1eiyX
tAhzVxNK2+j2f5T7kTGm/aGMZrDu5WptblqaMtvF+yhiYW6FwGbW0IIJ6x6yEo2F
7t5KXihKERv0UvquiGqIAKPA5kwMLCmp11XX2X+N6tJsTvtFQ1O6teV87Nyr9fEm
RKv5k38+A7HUa/mbF0l2RtFgEjduJqo5ak+ekFdBD7GtSJyITdbNSOBFNO39DeDv
Eou0U5Q6g79sbrHjUfx6uIcgoOTFQhMAmEghsNSHHRqRwvMIZ352vZ6U6ntz8TxE
d2MOzxjjTPSXcWzmkqZSzGy0MV63RhgInKcsiTd/2sXvmSQNi6gPVq/wzlMAuYf4
GCjPgCrSk4vNT4olfdiKJN0r5h0lGF5F/e4DYL0j+3MGP+y0wOyeY7nratIISDwD
33yVnHzMnaNSoFYA4iGiBGFNN42uP/BQpeON2DPuijBHY1vHX1WNWbXT6PkZcEED
r5os0yrsuUuhBkQ41b9zi7rv6dnMkXKVgHcIRVVLah+L+ZkZ2ZyN7tvKU+9fSiLY
bnrSeELeADWxYveaca6oIqUTRyGfXIYbjNHX1xulx8wrtTYlvkNCM53BljXY267+
s5g7BDsap+RmY8ZgHgarzVkaYkBQ97n9t0bnhXHGxWEVSGewHLtxDeq4wKuqmrQx
I59cxvFfbfxKwNKXRxvTlLg5pqfl7jGrPti6iE6UBJHQ1zGU+ugFO/+lniTghiaY
Q4S9MrxthmPb8RMNz1vaO5G7feQGr8KhUUt12VQf3VicqZPh7AaCchgFgN4tE4lJ
dTIXW/8B21h1V42FYa3+GsMwlIWdcf8XbvFwpLMt0AvI6nUY8X8EyEK08oU61y4H
Bmqzn3e/8oqu0YYdGnG2ifA5hMo9ZH7swqAmvOaC1OywjR9OyTQW/xPVyKLp4DlI
1bG7AOKqi5F5dPM5z3KhYCgYFnPgFtSrBG5Lux8fOpT0pCNEBnQ8S3L6OceGl55J
0DjrK6BSgAUFXMHZ+5VeyefTrmE0c7WjFC2q+D7bzG2nQtmhuYhMrsZYfh3wvaqZ
LVupb3q399fwe5f6l1I8KBUtfW1WojH1QTiMkgUHzLxUGWWbe/rR7fOM6+HEP558
6rTuYOCKn9RKLn92Ds5K33z5x/r9xa32ySszTykORcb2LEz/koC6PUXEcMhuzVnR
e2GU/dFgNj2P9HHmHTuAiVRntymEBP8fD638aTefvvnSvawEELkkmmKOkit8HxWG
PV+bKp+pP5FRfRoVzbiISsTl2eLKm/AAMEFmjkcGZAlFjt6xPw2M03ZY+d+vRR2C
DOolcz7wBDVL1Vl3pROlipCnpbzWiBoHoIW7fzSNQdn1g5n2EoTckFYpw40lCzCR
6VBKdOooARARkdK5ZLGV0F7Iv6qU6cLGHGEieDu2sJVhXuBGNRPM212y4R1g/vz+
RswErsiW46s9sgRbyUUDvHpUQuBMXZ3WII22+XYx02/tkIxVs8uaQXNyTDRsIVA3
fGJevI/2kV0hetTu7quYvu2xdz1lVmarCpcx7FGWvIJPonKl7J6yFOeKNjghGeYJ
1ja5ZKmCpIHsNsQGIZ+ah+sDMQjgNkvrx0cmBL2Rea0l26rNtmBQ6IZfHSYdEAXc
+NB9HDA+AdYpG43BzMR0Oj+PargM6wcAH8Kdi0I2AIb3Mc+0d/EuRzd+c+nW+bFE
35YZaibU6USWClaqdiTUY/bdfj8ln+qeunUzkT7jIr0wcbBp76XzSyGM66me4fM2
1mq7soNNe49HAM8q/qFg75m5mL5uDhn4KhCbiJxGopbGJlAn0754dNwyO5NDEz0o
Vegx1GIebOi1/cOCYcgR7L4HMLiJWb8bAOVyUVWYMyJOSpbMv5gGicPTDDnwoVBh
MCUzBWBfLMIU1SfOK7orl+VyVm7iBko+4Qb5Nk/s2jxsoN0qWDQJ53HPupc/kmUV
lrlObEhTk7ww+OuxWcPnb6sKETNGggwML+OpGOofmvtiyTkYYwG0IYlNCFj3Vg0I
cOqg/erWQXPoM85zrowx0iIskrY+by82sNnFruwSgP99/IXr6ydzeRLS2kGwKyhp
BaCybqA1OtE4XgcdVJASSsvnpplsAnrpiWK3PE25L2480c/VVIle6gE9cSkL0FrQ
2dVE8l76uoK5eBajjSzguheP6q3VGyG+3iqRbW3Gl93yyErf1OJoSBZVTdqIKNfP
PVMuVNu4QVVQf3Aa/RClqv2L9fLLtk8UuSzu3/5I1ga7nQ7WX1XqYdZ+HbfZgtDp
SLJm321SDGrtD+9pP7mhnoBF9VzhGexNtd4VxlYtGNrJegWr4j2JNAScRphCrx3O
Q82oZNWNa3vdXMOqiRAX7oIgE0n6KRk7S9BTu10LlMzPTDpBpqtB7BpKsV2vIKgu
420p+Jqf8YheeHXXq6ao1cf2JKB1caExoK7rApQaB1Sobnk98y78N50gajdH0eWy
Vz7tl6ueXW2v/rJdD9QxGZCpuaMFJIHW3pWE0y1A5OOyRjNI/kxp7nVNd9aAaoA+
qGy3+b76gj5sCUbLZsAmHGkpTnfZvAOeghAeVpo+r/qYnO3I8c+z34RwwpTkuVBH
uAmHzW3t25z4eHK0nVDCsOuZMcYo9cOm9VB0TVULwqRZ+YmutTSemIc+QQ6Ybx5W
eyVXQqQOv34O+JH74M9KTiCVCrjPOZJ6rtwqEFgJFFv1BXEO9C8XCjMXavxCmKvq
FelXC0ebY0yyeNyVhKTjPdW4q9xj9k4Vdj92kULrwpMAEcc/7+qCuuZyC/rqp2GR
mZEjzOHGkeMdsJxxTBR051pPesGL4dqbMZh9oWnY5EbfgcZrM7A2aWXphiy8PolD
eg8y5KgqAfbfOZ/2reI32B3AiZHsOItEGXwaejXrod3ccLMgQKiLXCaSAVGeoxLP
nEXheIKlMsmI5tmgF7yPOuizeJ4fUUG5nLYxBISsUhi5CyKMWKKiqJdkrxSsJGG/
yvXAh+DIFRomuy5h5uJ667wZD9M7AJL7tgeD6pimzuExDsm/nyBTwWFCiNza4C54
ggplIh+61VycSI1HtlqIawn97pFvhDNIeB26avjImWgMOZZCbkYE9hEN+YeSWWJL
zCTXcf9MONT6j/KVMC8jniLfoSdLkQ6weB5EQLllyUsb1+wwI/2idvlUkERSojxz
OxzX2qXiTLUnsLFGXVef/TSk9xbGjIdxus+z3soMrdwXeDzaDzP3Cb0PBaSO6M6H
tbPjLj5M+g8TTzImbNldiGc4X9/hZxJ9sSI07Kpu6UAr+1gpS8N1/AHDIhpLv0rC
19mHHYXK7mbc5pdIPBvgIgFeCiJg/tAEL24JjgQr1hH4pUfq5cXOae99TYb6Z/J1
fpG9EuZWKl3OLNBlSVLsc1ssItZJmJQYMEjFArCzS7EXreKRunCyXGbA0BH7pFkk
Uw5Reo1EjTWJXpErPIFE+ekYC9YMtRcjJEf7m8ywpMsBZ9sWTO8a+se0+iBwjx5a
k0w8hGicccXRD+dPbi9syY8mULxBFeSEkWbijl93vyiVW7h/UuRhGzbNa7pZVPso
hITPZMqABW1URng5z4e3Gx/+xO5F334JxSsNoJ4zg5PsMSE+Ip0ICnmAuGmf2TOc
uUsEEVmxgsHeSDNyxkcXDG1TNXz17i5zvjwMOc6oroAX+j9nT+rf3S+7zqoKBsle
YaffKTyYLnTXLSURku5nD9M2w4lRD7zKfYh6G6+LXX5s442N7xFkkYx8JQNQA8jP
WEiU7sl3spJ5eFLfQltqeuynw325myMfzFalabsNuwAHKm3d5JmNRprzUIqijQbo
Hx8sWU49pOSZqSJJCNBYPChXhGejYmPtdZ2H80gVxaHvM/zctlhsRVQJJ4QjAVOW
1i+Buw4X/xSJkJ4cvXt7lteJUBaBvh/SXnNWZSQRqrBNTqtKrjdgdu3QGVvcIzej
tOSDlnEAE6gXGtJ/Utl9zTekSytF2CLDSUHcG4zommEIj5+1rQmfXwJQVv6FFEWZ
dfUzTPJtwvFGW2hoD3zXq4R+04vYUdB+DrT8typInbcFW7jM14+32BNhjwDB+KJ6
0xRoZfQ3PSZyl74IHlqcIIbVY+EhFZyhPuRf3oFdcpzzNryPA1NLCkdOOApP/jOk
AASxdSnutH57ytLtvrj8uVeU2+tEJCWC3T23h128WV6TnJSUKz9aAmEZHy5qLzQ3
OqhavTKUD2zMrtPIJb1AlHjbJQ3yPhnvAVhAX59RLLVQ8TneZFwjs1obfakstIGw
S1IbLmdPI8c6xVfsN8yoatKst3FBcK+x2obLhnRiyhhIOY5465qS/F2Z3MZpmoyW
O7aiIz8U2QdxBJbCqv/q8nliWIAIgiYYlv1OQ6TglxAic1Dxu++Eys3BJ21IEiF8
iKh9s57PgDoPMCc6MvALGdpGGwpJ2KPxj7mhQAKFf+ssdo3owKGodGUdaRV3TwVR
8b2TgpMQU7E0T0DzG6UyNNELWknLskMxgLN4U7EeiNL2HZbxiWtjeyVfwK79XEft
aPyUu51qr/0y/aR6PfuIa0DlMJHT+v7SJBkZt+XJM1OPCqyLuQAw7oso9pN8dq4P
fitNV8CgdpeP2Z7WlWPP9cRZqlwvAJLio4b/anwmcMsr9D0lk8S20JvTHHS0vOUA
xvlMrjnsWSd9jcjW8qBgGU5yAOjzn2dTkc2IoSdNMdfMrVo+z0yJDDBA4cqUXaYA
MBCcLgwcUiKhT7OGgM6ZgbuYE/vIeMu0JmoETgroF43NK3qIRMjsyr8wuJtzuCfJ
n/L9BLioAXxWIwGiMzzfu0CDdLgWjQT/dcwz8nysTCWn6Dut3IGFXpubH5oxTr+V
3F5v73uik+hiUx4RF0LG5LvW9Cp3uB4jTxXUkfyRjPDEs+21q+BBbcKn0nEpke4d
lCah0nk2urZqMnXd5qZE2+p7NXzJwNeQ4rX3Xc8/Nkv/iIoqtPI/X0w7KwODza/1
qG3+tLaaqcVqZpxtwhNE/sqeHasnfVQd5Sk/wnLGjhj+SRGRg2Qzg4BXdYcT6uxy
0w2CCP8EHUgONcqI4iVMWwbdv2qV50kvDq8mKlDJDYSw9lGiccdrop3CcTL0lNP1
bjl9Sz6jnSuAd1kwgtDeyh4hv8sSoYcKtcKujBEUFwXH41l6gOC3aAgxaPzY034b
hf/3XAqjHXmxyaMgdacpNPKnChCpXJidfxuWZbawp5f+EZlCg0a/MwPL3PYYibu8
lRbJvdygBkwbA68BuZUH636PjXcMz8F+3vheQvxwZS07TjbvWiZUrU9HVyHpBeGg
ASp33ti7gXawB1s6jL9O6478VS96fT/pfuxnDPNE7mLQczIfvENGeEYOicXtQcpZ
2k9vHYVBKQzHf4NC8RlamrOh1sWZet9BpPsOuXSrsTdwZGCYzfbqrQgKVa5cqj9i
Il+Wf3BJJr3eu7iT4KM9lDL211TJX4M/lGBzBdmXnz/2Lp04Ne/z4o4MLDeWC3zt
0/txNUqiEHol9VsKIeF1Bwk6tmQHWyMi3c9WeNI9TP6ehJKXgXi1i9x8+X7SJyEV
oXYUJ/GmNIQnGUDsEIUGn94fb3ZbmDwNtTQ1LrubRDkdMGtCwszGdjDeOy4Ziozl
bpz0V/NXQWi9TzqhA3IuyGLp4rBp6Gypcu2/vvJQIag6SJnVgwjopbzIXne/9ckO
a064+NOqX/8TP3ujYPqzV/j33TADNAnQvw/s9uxrqDiiEm4jIVULOe5jAm0kJekX
M7NIsncEsh79KlJj7jwsF5xtmrPcCfXFaaeJUA6L2/GZ20WT4j9z5YclD28IyUOc
i4pkXqWwn/vKb0snv114QbEPsy7+qthrvnuQeGxTSYfJlZVcy7QDjSBGm6ou6YOh
IOpVxzk/uDGMsPKkMXryN7nw+Ndqg+oGi47sE0lgbCWDwcIamcHuERpbu0cNPMNT
E2o6pypY4XEDwGV/mygayOT8hh8XWJIJENDABVp9VgBGidwD8EYVo8IDOciHE4Qo
FOu22wADxzoinGnWLg8tGuSQbJ8oNuQ22dp1ZsoFg7nA/QEAWyWSI1HxIpdj7CIE
c/ejgyVspQ9qLNrizd/cUTHP6YNWojEFoJaEk9NATsLwzjRFMvRx+RCyTp6hx4zT
jG8KLmJkJdfDLYHVaLjQjPfi7/rn5lXzrFIWgNvX9k5W4SiEYUUAUXbSc0gKP3K+
JSA/9S8HBEMnZIVibCWGwwZlZNvylCGxmWY9CZctMb3TmPcQ0Wy7oF3yxYcjWBtm
h92RKTvFtXX0NfKi20GUcceIongI33+iD5gCAvQy0aC8JjswEZg89W6+1DfAXId0
YuxE3qgBJrM5rNyjeeHBoIdKP/bzEXvAko6Djb2w7ykW7QPnhFDxtGnktzF0Cv3+
O/Z2AekqwF6T6RqrRtU5qXUacRSbj6Bf7tjhFeWbDaYunsAXIck/kPkNd3Dqg9pV
cWdudhwaa00iIUsi2YO2Z8wnrOHXV/JFhi3QKf11MW8rZnQeU9OBV3/ed0WSNwq8
HetwotnZklDsIa5gDMzORBDsMQgCfHjKc5hJypME5yEEee6KybbEZOryTE/JNi9t
uR8LtqWP+f3U7HkjUsXxYhtMzBiiJ8WJWq1sIT+brwpwM9NSQ6JzBMbBZEEZAcOs
FUalGKhnLQ97genN8n2BkiboswyDQJt8J+bTI2VZRpGuY4xkdOXEe8FA/28scuEH
lbZQBAifJQ9xDu4pP7oe78ruT5q3ZiUorug7cRGXr6Pc2KBSlHa66WllEzSR6LYR
e3lAiXdk+/Pw7A4+h4ChKrHNkykDPo2F4V02iKA/VVcFVo3zNpj7yohVpYbqcNYb
ivd1z84roETVO71QroN2GjAcBWpIzraq8VMTkDeeftQ/ccxFDsGMG35RDYm9tVV1
g8ewPh/uF/s7lds9HSktV+JYYpPhqvQha7Atm1s1BwxtUkYau1J0hI/iQ2Aj0USG
0HzT4fZsrK28T5TeBX5kEdw24gyF+3Vp7KnrIAUNxNkz2pD5d0ApEV0qczuIWvg8
yi0h1TIRO3WvPBzGnfG+ikNkpihgot6QUzjl5c9syhla/sfRT/1dhAuorXQf20HI
m+JD4q71lpEuQbScYo5JRlvGl/3qnSMcyC1H9i8UKorDF1FnpvGes8lD+XSu5lL+
sjMfX14ApKt3hLr/wR7SE8S5wqzagjJ2OJn/YuVdsEMMquz6sP6j/E5dhLnxWncC
EPL8mpvmYurq1JIP+mpZlJiPBlgzyymEEKFGqmUVVckocasQVW2AX4YZ6jPnUvpL
688qynkDkHhtcJZvoswhh6oQHBRuPs7/1va4sdvNwOcJtL6rE/SQ9HcsZWM9k+Dv
B1KHZv5xURak/X3UzJrOyCDnNDjQ0y+98rk5iE/cntZ4J1aBU7EBKBveFpKUc5AV
eb4KkWXxktYo5GwEHOPjxrZ/Xf0SeyHs9vEB/wBerhQ14MebN1zhjiE3+IEnzIw9
9qvhV46SCfdD3LbnVh43w9FliqNGygBqt+Jcwnvgo/sJk2UzPiT1f5WfiVcTlhQq
/iJcA0FG2wLop5d4RSm/E+VLU5KHgysTnF3afHqL2U7H9ljGFlA44bZ42QcgloAE
BI+Kld6pTi3Sble/Z8iIXQXr3UAzHbmpoCINW1QH1R1NrbTldjpRk46Pwt/LxkB+
UPbAuoTBtCFDbOBYxFrma7G/vSvtpCGQRqkUnQX7NLZmvpMmK8xDglmgYi9ICa1e
fIdnhgHDWPH3R2kvsdHTO+vOM3qKHTaiyvJ/6VOWMZOfWnt36uEHKJnsInS3ofqZ
MK0xT9qytmqNAx33RkT5qgB7WnUkg/+r97ezQisVVz3ElWxGHnEWZmQnV2Xa9lqO
viX7pawhl++gWXwT20tZEipqKRuY5AzA/dbdc8QCQ44zydCcvlnZHhD3kd9qUpnL
2Wk0LjnE4SSFFJghRNIhT4zTe12Mz3wKYgs+Uh5MUrIAVZjMAq04ZQHTxMvNgY9P
/9O53HeBA2jBKsSTGX31J1thgOk6Vomih/kmFTv4mgro0mNZJgUJijmYvOF2ZqrO
PG89wgzoY22rglQgPVTc1PZrfqIJyFk2+trYeqEAxUf9u0l95HVKwXiFh7v0NJOF
o3Zk5z17WdukpHjyYWvY9eDjN3A7kJLq324Hfz2IPLo6DZZ8rVoj4lkkFVWAB93u
XkS5oHP4yccj0JmkxkFo0/H4L9/BY8AJZDGaav6Yu2qVrIBdaamb0llbjm1X4wQU
okWQTsYK/i8uKkUp7OYx6g65caESjR/krt6tr1WXKWgFifQbMJZiYu6iYtv1A0BE
qjGbh1S/cbnZ82oEN6hxhgyI76vgw08/1tadyp7xOaAMsZktgqWA2P8endaWnPb9
H8XMrnglaG3SOTc2irQ6lCZap9m4nkgNbnzkUwB7l+ozfzp9flWHBqNJLErLpvnt
53Gu1v+et1fVt1f/4H7kqCk+LrG7tpQnk3JPYQRZEPHGQNysFRSFQFXzArawzXs/
QDEfayiMyssArZJZyV30q3euKfU9FIOauuCZKOOiexHqWKVtxhP8fIhkIJyzkcpL
RohwDy9ENE8HqQIcNGA+mKZhzNAiT1nEH276ZV/twjw3ikr3DwrWOmhjPZqwOjYw
FL0E7whiDyosbtq+k3arnG0RCD+0RFrjHDaRibwW1MdxRTsMwprPhOQ7ZmiCgBJp
xAW/z2ycgXZS9ubcnVXmRJ3W2hM2W+rdOCKVN8BdB1VU/jgfpnq4pbdto0W9YleO
qrD9nrExj7GdymvLIU4iTA9YyrGoVbVaeI5GRqHvSvnmuzyBroHrt3Fq+/Zgh+UM
fFu/eow2pS9H3l+Jo5uDnbuuMuwtTgNsyAG+SHEpe65MAk/wHUC36BjYS8RwoQot
YOt8fSSNkyAzek+xiltzpFHP3OFq7sMPmIVhZ83FklI9m5+/Wn/VZI3l9I/XiHUE
UDI3naLpUnVbekYuAWdOFvp01cHTFlbqC3F1fnVlqotX72ed9swAit5nYjoLvYL8
OlUL/sndioLOhPIY9qeDwYIx4gAUfswkTeciqzhujDEuiGPSVM0b6IFT0rA7qEnZ
VrMD6XYJa49E+KgvO45bC381Fx0dDFMCMqI1S/H3994QDMtWRF3hFZ6/aZeBGMQd
l8LXUzLNUxEA9/jWj/ij1gFkZqTazpg3ykJVOdfMmojJfL18Zhmnn9XA8IuQrNQ4
xmavTQLv7giE21E0vPmy2IKhY1M/XVvN4tVGzscIrB4Og7JfUnjU6qhP9p79+vRd
VgtN0zuFO+OxG1GVRQqkpff5T7WBI2UknaP1rJL0iasS8WyMxVYZXwMsXaEQwkxo
uEd7NKWnVaH7ilrWWUpYJBRaBEkC7jUIucB8I4aXMxuz2nwkczNg3/7NkqBUIELS
x24HG7vBA1jjG0zgG8UUTvG51ep2C18+k5icFCaMRLR82rl5kBvu1Om7X5pwLT7a
yq7MMh2YAYaNX2zKcyvbwR3sXsxsFzsK6SaZGcYEAT5Y3GE+mAaEYr5F62oGk8q2
AWm+Tt/dOVsBnEVe7h6qPr1EKxEUUjYek0AAwgpW9eRj78M5xmHiLXN2sZyxBJht
GKNDnkkqtPE5NhiUcfToKrPf3vPhg1bWMcBoBpPBGjs5LFEPMsXM7ubATxLamn5r
L+YJ5ZSgSs31Ty8lj6PtVGza0XUw422VoVbYEncwUOZZW75l3MnbxVc7MkmRtJaS
DPfGmpWjUBdlKnce6zZgvHv7oJ92XqbMxmIwQKAYRhpHhOa3o+QBrdSx8yYSlo3P
Wzf+NRha6ABUPyxisjy9iei30gRK2pg+1FtpNIN981lUyj/5bwi8dEC028Jj8zqg
iXW8+TVX0mApG33nHvRThdDq6B9sq3nyrJhWbjNYtdceC/XCWFn45UVkV+EtDeec
L/cb6fi3wy1O3EDxF7PYOAwDfnSyQLayHr+H9wIgDbXAf3weJDopEDkkeYbVvNBz
Poc6N1CK2B+wz0sjbicUADrWXNtsrfmQULRwS16JQcvWuq4hEGKC1R1sQ+FmKMTO
K/s9TXTnHWOPX/hjpIv/VQ9+A6brBI65WQ5Qw/yXUrP9BvVhpahfW8WhrWmq8WdG
ciGzMA//yGTC3/L5MLcnkU9X4fy5tcUli3OK4HhtJaHzSwVt7uG2rP03VlNiNM1F
yoS8SCh7lRBIzImdT49LgayRW0250F9zKL10nnI9JhAwdqmAD58i2cNLm3ttiKUF
guDklhanVYaUN97wXptfaRDKal2e801LqDJ/EiQDkYEEGHqWbg4eOSBzwFl/g4Fu
zNdSpPoDGJwonvL0TGZa+kQb3m0M1olL0HziLibaBXejYk0auBQBnVUETt/3Ww4z
fHKwcTVWcJUuZ9D7k+rMvuLbC4i9HJs0pljCIkkVL6xjMXQ3MgRyCUM+xGP7qPrb
8ErhXG7Nib0Bi/PtwiAD5ckHdVnuZHI7UDXSRWXyMS5rq4QoLyK0d7nHQW/GX9dp
bYQoEmfxW03Jh6w3BbCIL0buDkqsdn1o8vCWiGBWMah5qv6MuNYnkRSawlJJAwIw
tuCMhtt5ih4k4mfG5HylPDdOJ1KHuTpOeRGswJp7Pap+gj7120ekJ51QmTLInaTv
gFWC34RyZqg/aEVJUuq2oxiM/VMQVf1HdmifVYzBDjsXE7rXW6qyyz0I3NG/EHDS
iG2j5EGZfTjcFSxQJ9j/G2q4XbDenkXVnMWdeiO+zERDqqonPxyH8ax1x/A4E39w
Q1k5WGi9ZhP1/Xcrg6V3sVFLfVEJOCp+PkKSsMJ5xd38gNbxv9ErEnVXd9mTuiBQ
40AhDxkxxSWkL+AHqyfwCdYb4g/nAFF4GWM3kBLk2Uf4RPMdzXiPVAkRqPjWHgjX
GsoksK2351zyMuL5oRueuUtmCMgJjc7bfZn4NpZcnkr3kwam0MR0GaC5Ta9KWnit
/6ZfXHF4ZAz8DL1X6QR2WU/OGKzWgyCY6wbhbNJzhsC6PLcttxGkPH49Q2CXjqb7
xFVMm98VGt7D2ps9umQ//2rv0n1NbgZUe7YIJAB6ywz/r2hbr8CtjiZ+H194VL6c
GttlAUkJCErKExIe2ZMWrLhUkJqapEIVwrEiP4yjttgjdv8COIxfjq727+Y1UklJ
1D49Z+PC0GqatK9vEq+UX7+Aa7R+TERvX/zWyH5KcjR2JYHzu5A8Hwq1gkuyZxLj
JkZUvtVLUDuoPwr6T3ylBMZRr5inqR0qVvgK29k5OfZElzMdfw3YERaJV5LlaS/p
mgzRec6RA5thxwuwDzx5u9+/cUEBS7PxGF4kf3zj6WYLtBSS+wnGGFNNnMMWbTXc
2UrljUVtV+FSFJxnMH5Ka/udKLtRo5saPj0oBjR5RG9ynDOJN/4nPwWZF4uzTio2
dLOpK8evPj038NtUyNrRycb4bjhD13Uz/a0yH5ZhoDtHaBeyOr+joloE8Kn31SIs
i/e4eDj0PXiNaegIUNHkRhj/ewWtDJovaThCQk7i9Q7bfYj7CGJqbZVVjQWcovAT
CxBKNMAY/WsfxTP26TMf5i8KdnFesRuRTTAkwUie+xjpBWOBYsfgyT0NACeVcqEQ
kxTUMuSACvHUXl4fE6knNcp19d2s5XCWukoi/TsqfQa8oWIoY7TlT29woOCqLzlL
37cX0MJzX9r6uUt3yy3k2i/b8moSAL1zQrqaxx2nh+J+0QSQn4MWzI7RLexb7jMo
JdcJOxEnpORakW+18kflapkYJnr4y0M0S1Q+Gn7EMle6mU9thp9/WJ9L1wvfz0hn
8fRomQZtWxK+ahNxCzG090571wdrKqpdnWSoEM4SZKosCc4iKsmDC6Q8l1veZwBs
BqarVs1AWWCvk7ntysv7lT0XQXgY9f9dRs1a5I3MRGZK9dgAX4IdOMjgrkB3auzh
h0zb/KTtDUiNjgJnSrcISre0cO0bExApy4W1Uz3HpkteX4tftUkx8iha1jwmCsBL
reYNTL/Pl0HZCH9amKdW1o4WPIb5/SzpQEBUXKosvaR5gNBBN/lUHQmFUsUaXP8D
fZ1bdtPAs4m/7TG5ZiofUh7O+rSprTNV8JIJIZQEOv0tVuSWKu6bXSxVxYL9CUy9
HjyKg6XLDSw7ZZZTIYJD0KM41VUrTOodzsTXyTqycYAnaKTvNLBx1fnGCL8TO+Ks
tUnKbAzML8VMY+A/zti+QgRVu/+7uAfJOtj0gI+C/SPMPuF720XvP76doRIpxwAS
Cc42tKx1dI4jbPa1lQCij3duE5cecehIG+j/pjEVvxVmKnhcZodxwffBU7RMv/BP
DX1CXk4NI0ZlBoMBkG5xQINyVbpHFTmiRVAyC1kiobqX4CCSDVSkbBgtDYtlLoRt
y1Z0CVcttLdPrSpi2VgS4aPzKNs3P3D04irJm23SrL0UJ9i1Wn7Pm8QfGPD2lofF
MFUH0RR+jsnPd/kcrIum3wOwbFwe0EDz2GxAgSJx4nw5tEKGwwXbmIQ4O2NE55xy
gbCe3Ik5w8dRNEPN0Y8m7u0PwE2z1GNrWEeG8f+DlKm1hnoCZUTW8yFcvzwbeaSA
/GzenVaA+D2DiX3gXj6PVqLl0gxY+bKggZtoFJh8VP7s3QXRxEVFJ+d2VsX/Mu8f
9lK1/AWksta2M2xS374yMg27S2ldQIe0H3CUNZhqzS4XKqTcGvFwRNhxHeIN0qBh
7vdx52nvD8M0RFShd9PI3TqwxX4ZZGQnP1+f3TA3+VeeYLJdMr8RbaV34qcwLd8S
G60LYjnfq+baf2TaWGkSHQd0Gk+fvueGClKsKw+5FVe3p64vXSkBQOMLEIc/7PnA
i6C/OiW+if3KpzOGb4MXgA8A0pEN714hgUNHTp4kgWBa5FFKSdRpkSKdNdH2XAgb
fXtjkC4rJRjZdOIyaC3rF7mL8S6lry5ZLiutt2ZNsEByBp2zb0zeO3oUO5IDfw4Q
lTCvp28fU3sfNLf6Q7YJc238S3103GQJlmRdd1DS5kLRksCdszzryDckuR2gXy4o
bn208PoBSal7kLJcdBn5jeivp2mHYoj8e9VIX2NWrh9mKopv9g/uEnOUyOWTS14R
Op6D2HnPZBsKbITd9WNdU2B0/1WRvE3rmn3KnVMoLzoKcQOK7Pxd95dBpiwWU25d
UjARjyPXNh5ayusFhua4h50gqLlbDzY/GMZkBuI5TMgBi5EyuYOKDonDzoPwxwZs
pxCAcylSBKjmadkodCGP+KhUYBFkFc7zOJOrReZcpg8/27FC1E0j7zutSSlpGHKE
G8y8qaPoMLGOqUItPW0C9SjbMoXSf4YueCMuPNIAY67YL1kzCrjDlj0dAcoPkszi
1zlniqOIkvrwwIcyxLWTyBiHge4PtSJurCpLRjVH0zAx3R8Pa25XATDggv3XBRRl
BMXr/QeNJ13EfAqn3T/rCPM/CXtMFPO+QHuMbEAIg5iAp+cOliUxB2Xb/oDd5qWF
VbjiSTYwrSmKjfl0TRPpSKmgtMlgl6wfPD9KMzd7cRlIBSjOZ5SCfvej7OmPqgmE
pCNmFKzEsjkPPXNThSR5sYe/WBOY9CcrYQeV37eskxOJp4FulAq5fvOrmHcIZjXX
u50CVRCffvUgCmgbyinB1hz+F1Bc2g1bCqhIT4wq1jKB5A1RSwJSOBnEWsrIIy2k
mHWjQewOkHl5obyjOH1e69LapioJ7E85OBTIX4qhuxDxKXv4ThV9UGTXioPvbs1U
H0NLZsIWwcky9lJ/8DEYVEqVSOypkxvIqRxhWYjVdgbaventcMS0Nr8VTdmtKSAy
Q1o8jyqNFt9mpnEx609k3gJWEx4mjUcLAPsCOLIur1ECMRiwe0DhNK4YXe36bV+L
mtIoigovIuV09rSR7B41qgBgeFKyhkRnsphIc+vw4RJA3it81X7aHHfjX4i2dZXJ
AXJWaE/8pD2U4O6rKVH+g+W41PDub4dHOACmX3wwtOtPnWM6sOhqOaFkQ6J/v3Gy
d91U94it8E77LLhngknrpY7/puS2+pnAZby3ZRNgWzZ778QzfRhs5f6/t+rxI+uf
nOGUxNIstUR0PdjFIYckj4OgGM8xapEz/4YKzsiek/bCgxTye8k5cFO/2NSWCTHn
FgCBLhVliLNXF5Mrvm3s2xYBc2MCVorlWqYRnb9wAou5GtqrdYRlcziF5iq2rBGG
4WF9dml/lQZbhnearz2GLnld3BnA/9OcS0gvv7Zf286ptOZodckI8ZI9wbqwXAcT
GjVOUF5X4fDAz01TwQinrmahDpDkCWmvH2kPwFAF5jGslgmXoOvdk1Foc4/TQC32
i1ui9cFw/ugaSrAGZdlNGuYQZozxtVcQDwEVk+9G7earvaes3rfVkkLN8WNrOD9E
QguSIoBshn/B0hF70334PoZT4qZH8iAGVvWsRlTaFJkt4Lw5r+sLAGGtnJUxaZzo
ALo7CcJpkKjz3OdCmgWLubMqV1J3SkzkQqM1A2q1VueRtK6B/eJqi84U+Y7OYR+w
TDvVla1BA0Pwt8bXclFEqOYgS1N72HiftCquZTKHGB4+bvMVrko99ZYsdQnSK1in
dS08vgnl1wNOJwJPRZElltXb3sRrBSNkCBPXYfU23KSbU6reD3QNnwOFrNLJdSQ5
pgEBrdhQkcWABIpNdfqzRNR1uGANa6EbrhDy9yIizzDIUgv+pijwvzNeENjxJFVg
XrT217B5N9srTy2m5wl1UYIst4cajN6dOWtYE4JXk75z2BxAqnWLEVxfh5gd+U2c
BI27BNgvYd1qJuQC8wJFwuE5slEXj3RGNxCEPYV8cy2z0JU0ILnRiwwFvbV+6Qx5
4s40WcH0cW4c0+AcNIPArBvM/CkD5PHrV62SPhH1gnlik8dJYxlBntXfCbH5m/AM
B+LA2L/JYDhjvnkdvUTpVG5AsamGNQRhDxKZT7Oty1NVuvhfDH8fh/XeFezNc82A
EkCnSg4V10fSvmLWBM05LvLyDq1J/qg1izlUwY36wZeZyrmPXKVNXhwayNjBXT6x
Uvwn+c06OEwev5Z5yNw1HGvp/GYEzK0v3OueM0NQRapbITGsvAmTCMoe5yNHV1Zk
4MY2Sm3yKtG+X9EGf8pRogq6fOqPNX6YXaHSlz0U6Ktz+Z/yVwrMEz9SjCejiy+L
pG2nfYZtEBstKsSCGK0wUBtBoQ+raJd0RKSZddQ8bhH2SKDXG4l+sZB8u8p/kRpZ
DHXaLEheu1NiPS21dlXz6PTE2mQtwQm+6Viw9zxhGMHbb0cHlMoHsVDHlMdgyKgm
FUMABcvTGUV64sd45BLReIRQxVnjqXKreNEgJ99WiMF+oUqWIXNsZI72LN7R7aL5
y+krbW1EoEUWxjbjXKlMXOUKAGefGz+RNc01c9Dzvxt9aULSQY+niUAGe9YrseyM
ONMV7CgMKCrnCrHX4dL9h65sSXUkr/7r47yiiu77zL6NEes3TQf97plWuHnJx2Du
ruMVZRj1hpoWFtUB53/GzVCKgN6x7g7m/rWVJpfzKTiH4800qToCM9DyJk3xoCRF
KAWTfMeAr7aBleGXgGUNYuLxn2IOS5n6TLhvs52/5PXUYYn7z+MEF/Fx943+EDAC
qSWliy8vk89if3rNxdh3k1QJuNR6SYWq85PaJK1qUXBP4sIO0c7vDKlGJKrq4X8L
K+GuHSgJ9JodIauxjRzqUw0jpNOfuhcBjc6alzleI9H/oprCGu7tMiFFIp2ZqJR0
Ow7SXtlk/PjRR/j7b7+XMOmz1TEIjoqFJ0i0VMKpleQhIDFY4PTanfnfE+bJ/5kI
mYQpLGiWUjzNplGn9Ih+2x/aJRfSA5exzoY1m5mGN0TOxjygrGmxypQSRtZdtERj
DsNHbF8jKW1H6w4KiAGiCkbHUaif5o4GuBRgobEYYqfuzexl3jI65xDP1aydrU6C
xY0CddpkZCyEfQVTQOxjaaFYYbIUx+E3B73o7RzGAhwmCaM69TXqLx51nICSp4c7
dWq2CzUFxFzvLViZ3qtnEz7yEaE74+RcktBekHFJ0RT+YYaVnlapB7eF2Waf+ypj
A2Wi0U8L1qvmOKOP/JLFLycQKBqKsvDFa50Ae8OyJr21xUPQm5rCl/UyL7AWlSlm
b+0x2CF7Qgf3lVX80czZwfTVm6HkreLWmGhxaCb3hAffEv7H2mw+jUXT65GlQWTw
zmsm6Wp+WkwLleyOFe0ihLLvBQw53lqbSB6cZqrVearh5hJk7pBmJILkUFRmfm2c
4m4C33C708MysruWSdhXRv+2YgJC3FkjJEYxEDXWVo1tYfI6THZa48rMg49TeHlT
ql2idUF2kqhp7cCCLfrRne7xeJLFupYMFj1Gbrs5nwtRtfFh+OgCwSlrjuu/cv/U
cgqt0HRddyXvaREVMTFJfnJ/x7Xxd9pMVlohEcEPY8xKOgZX/+3SYmag5DNvyIZx
ZkaQcKGBu6pE9+hb6Ov9WZRf194LYIFrAadAP3X97p7LeIvnw3i7w4KDV6F1ueou
7WtX5gKtyKUvgakWpejhB0oLup51orjgSzt6oim1oBcAJrKBRSt4Ieba09OoEFnE
vhh70kpJdEtf1nIA1kZsrKeocXCGDDzwO7xJHAxly8vnXicHHbs68l3bD9jl6iL6
VWmwULd406Mg7L8FeTrfztnfcTXrFPcm1REuzIPs1F8CzaHg+mEaXU/+dGUSXEpj
YwC2izIT60enloRLiBLpEkyOnlJyndTW+7y8W+gFj7eWnr3ZAaueB8netz23I6mP
g8mHfikLYzS+pUbBjWIq2h1HPW96bqy+9CzaCk/J3/d4uzFfjihwC+G1ZFwYKe3Z
Z8eS3W8hS8Qz/N12jeVMbBKshvpo53zyXsOyMLWzOkUF+HKym5YkDk0nLKpCK+qY
bVQ6UQlTkGEnUCthKLRSHHnz0l4BezrE1Tllz2rQsCvlwUjiLpHdpbC1BFsLQSwv
GjEw8KkpJgakUIDPIHZRnXyoadcXhvGfpCeag1jpOE00Y3VKEL6S0D09PBAnSNVq
pAA0MNstjRA9fDiiUnGJGvI6i+g5hpxxe9K1Y+gdtQVyWypwkFFXkMsf80wEMxoz
MroechoTOzo5oIMD5GT4mBhonF5E4yO8fEzEQVnPChSviyNRT52ahd4jEiFD64Zl
WUCmcb8l7ghmYRSy0z0WMNZBqbFPvDst7noI3apzDqWfB6wlo2k7CDJMRihsCPmb
a5mFVdGQernp39m8/hJyMhGou0t8M2wyF1EC05pbsLtyNkYIPcpdSLcHAEadur2S
dQdoT7+V1bdISS+WQVcnaoO6Zqy9aHOebJb+zP8akFcvT8eTr+xuQPYv2HYYUrcK
IY5Gl1uEdDNYeORqrfUYfhP1HDfbLw3GZEGDWbdF8uBYZ4d4mkzWCJxYTMeQXwm0
1w4gGCoJaSfFpqVcXrS+d5e5F1PPLDJnLvr/G/XdtWbCy9EQiV1wzFrVTGef0ap2
tUCbzB/kst/qUbjJY5PqrsrMmFbgbNZFYAGqxkDBm+q8jj8SLkH8b9zJWVRGA7MR
+HA3iFsU6gHqiSU0DGdFNOYKxA9lmrE8h1kIo6pcZaPTNOr2w+udSsWYYnqTQuSt
MmIIgaJB5AZhvbrp5/3JjLmmzs8H6bK5MXBFLuvRC+OuDT10guIc6JfQD+tNPtNm
n9N637nCoATc6a80Uuw2s9yXBeIHIrK7pbbdAjpu5JzgQg688MxLI9Kujt9CBPo2
nacMPeMMgFJrE9rvsYixyb3raC3nQ2XvNviB384+u19m6IM1H/Lt68pzMr7R8BA1
XiY8Q2FEiz2Lo2C8Mb+upaM9CFU8cIOIEgaKTTh3w3nVCG3RWR9QUiWbfMNW+pvJ
rtHhsEUw2U4roWsaO2iEW9YgkIlHhiMOGWxvbUL0iiidz+l6z2J/jUxTpioB0sMm
YGut17E25mZlxGOVVmTSZjeF7FCwAmWLz5EW6U/2FRbel9J+0+iNXfRIRNhi0g+s
2XuAiGplf8MlMZ6cFAeeov6OA8rH/mWowFI6znB15RQO2I6m9tDLPDurWEh6tS/8
YpcFklfXUp4IuTmXlU8stWqISutEG4eiE00ZK0ORaZfitDrHNud0HF6wPsYY7flo
xuTz1itr1Sd7YV2wwAfAVvd9FTE0q4pMUIuOBW1+/yUpjjFLwGcYB2zzHUBBBzve
MS4jB9u1D71kLZC9qC5m7yuci1jDVRoMCMWeJeN4uEA/i4pfePrmFBHuPQqacXqy
TQ5M/uOKf4mttZURImwrYB4sKCLBLIoENCHqOCoyPYVUuL07ruGW20gQXXMNZ5bF
XnJ0vg1ZsL4glyvju8DPj/v/UyKMCw36uYIJgU53gUKRJhgz7Z/70bX79ahnvjK4
1vjRYQlJKdz3EPojSxIg9Ovk1o7wUFULRMz42Yf8uUCmNTdrgnJ7OKv9cO3IjraL
ISG1yh0I5lu0gqGQgLi+1113RMtgVnpCKCJZCRrkQQBUTVhYmF+/oJxlSq6PxZ7P
pu34EiQ/RvEfntXdcvVdaVP8/WIQz72T5UAXSf0HC+dN3bFnc8Yrtr0CxGZAcerk
JTQxhrlc1dffl35EXf03Km2C13Zy8pU97VVRBbkGaGSLglGJWMmFjxwZDD5yYiTN
56XawWLqxwohLcep4xPB29pkk5Z1Rw/MCcvy3jmj/oolOoW25RlWq/tfSRedjhvQ
g/wpK/1OEuAA2CYPj2PWFVOQkXtzAKj4jHcwWiSTwBcElRK83zr9JsKXw49p1jke
uKrUscmeDnOcYII+k4+mecbObcQ3t6QlfWSTKIrln1E96vZpRscJkJe12PgqTnqL
u+RnjVo9aPd896jOt6SaejzHGGRmGbq1di1XtWuk7r7ThUae1hk7Ycm+MoTf43PP
TPClTAUFellS9UHV7ieAMohHGfH5pqItLXCZ4WGrIWdxSYqZpjjy8L7Pcs09GTUe
9UCiiA+tPlJ+wdxswRdPLqtm8Hci88fkcyqNsmnlIC9E/8+a5O+uJuZ5PwQ/i1o5
1lOZTMMd7oa0SZk82Cb7qPoibxD7GDn35vQtx5dYH46+0jmvKfHJIF+E5eEliwHO
UUduOcBp8o/g1SSKpJx28cBWNSsPMRx642pgQWl5J59K7lcI1hRjnGWo/nQ4uDAP
pD+iX3xO4HsRYNneF/c25OncNr/t2hdN47BemD3n/V5oaXRM+nR2HmhZuDua7rHD
i1HFiuxB8eW9QNoyoXRZgDcGSHhRP+MpVMpZu6rYh6qVxDc1pMTsqZxc29mKw2p7
ucv3YXyqtPtz7XMkJUUOMc3UR9PxIJqYqEQOoTMEO3XnwVluDjHySaqLbYDZfddb
QsDbsyvfM6kweScg1C3WYbQjbQPcg8GK6wisbTKThyMCrzslpuwt0DB9JgQEsA9G
jmW/w64vSuGlpuAL5RW5Efgfa7+6ori9KISx7GUL6FSoRiojeHZAxb9Xkw1Z/K8y
11sbS9ApcyMOjSMdXV/qX7D7pJ5BZcSSwd1QJJ+0h3dCWjI8PDT897C+RU3rcyZ6
afIyLv3pBPtk5vn4MujxGhjufUiJ/nKKUI6a1kc8Zw+8y9gLiyk3Y14ClRxwnaV5
xfBBe6RWg+YuoqE1sqTEufYzFPfMF+BcNO0lt2m/w12nns1ma52AuzF64p6SdDv7
NAftJ4RjPzFuo7yY2JgFU5axrHbLphmg9BAIJpq/0uUCDGwGFv11oN1SGhZDgmV8
hhAumC+U11McgPn5GY6bPnQPBf0nbeP5UXay5sPZhwdlNGsS6g/HWF1jHE0u4RCI
aoe8E2IRCaxzzpAOWOW103YebRBwFkgdk5Pl3Yddso71vFflGqEyk2huGjnvWB4i
4GDRqGFAKg+J5xAelyeYgA1EPv1vO69H8tzRzGFz6OIgvA+lwL4w6w/5NvY6Qv+W
JbOHzdziyhbkAIK8rol9K1squdJKwjIL2RazghcGqGgpP2qiYtaCDFn5bhG6mKrH
BVI7fyMPnstTqb3HC5SHvqz6ZEuTHfunYYEb/fSGl1L8hUJOnigDLwIkyhYA+sya
OiPle9obaxmXicbL/KScc2MnMNkJpIFloBDkv/Bzo51bOSTBVMeFz3BEemH0Y3Cv
gmc0bPUlGGdZ2yoLrtf/Qm8aF9jnztQjiNpSZZYwoXEp4UJm1qMy36yQ9RTlZ2gG
II2VyTbVxV6RRyQ1+e1RrD6mtxRughLLDHbzmDkeWsofVTa0JdduAOXNZAUnZQof
b692j9q0nnDfTIRQTlI3UGHjQwKqvm8QcyT0pr91BJ6Hqi2bduNOjAwZiJvNSZS4
+hESypE9p3d3QxBH7BBCKncarCE0CuC6gMp+R9yJxs86vxpZPAfZFZ+EkEs19k5M
55jZU0irOXes6u9gRuQ001wOMshdkd4tpQWtQQQyEpGaxGiLfur3B9krF1Xl1apq
Ok+2cpzdvNtY1030aiBeg2XZ11EPGerJgfQALh4EI4jjNhUWlcr7ECLXxesZavKN
m5Yxk/Mj7gpGN1NljQyBmus9i/7x+iCIxsQNxG1SYuDoxU+nzppWu2+Hn82fziRY
qWmBfLrayy/RqI868ZpSoT4qGinTaP8UJ6nXL8UVtRlpllLtdRuFMgUbBKnJnHHk
+2Pv54T1N1sjaEXqiwRyWQGR6VOCviKnfcN1dy3Vk2Gh9Y0CckWhz/ksguS4KETL
FpK/Ps5daFFXHD9GjwdN2ifs93PF++6d+iO1cF50J941OYSfmMKbbzeYBtPIdRUE
Ie355Hh08fXACGXv2NlpSEZJchRSvWqvWBJH5uXhuSN3dNCRe15ppEzqgmU2C136
cRSOIOogWaUhobtoFzb4imwDWXBbi+SJ12uwcSCmFqEg7CIaCwKJy4oaU8khUfcV
VM8wWxyvIgRpzsOPTkTd1E2hTClQGWSICkGRK5GwZLMg0f3S6wuu2f593mDn+e/N
drnlkQ5EoaMGjj0k8509LpkFVKyc0iHl9VPvqLBzufhUkzHmuwahsSW4leVaDy6P
vFC+B7e5jtNG0NDhrO+DIlJaYNcFEZ7IsgjXXlRq/MvJBrwNJch8Izn5EIhVtLP+
hQdYXpJss9BBNMb9iakdGr73IPfr0M8D/Rfx869zh8M9WXNFtmnFNdZnPVBTympZ
gyNFtI+EqMO9llfGC3CEbs9Pb/A6ti4xcUKjI9PM8gpMw8HqUQupnDgk3FJD7nlB
sHg74/drzuE4PttyTG13kL+9OsReqU5tnb9iJJuouoFawfhV+go/gto5AvtUxYIG
N9VK1LFEettjcr7KptHwUXWGVFM0jHyyT87BO+/gYCRsWNR2RhgsutERgzwT6Kzx
alXS4L348OoejjaZ4/u3ZhabuPyh4TNVkwF/jrkMyNdjyYnqNWNjMkzT6TM3yF5K
n432qBhkssEbL9KghbktV4VTTt0I8YWxbUc7oLkSqEthoI9QJ4HmdJn6VJcVrrMM
o4OA7uB3JwuYrjIx3mekF8AnlgIwa4qB9YBmdMZ6sAPiVttuZEsQUsa44aIwVwhR
YJ4yl+V6jU/2ogZB5CDb461yJsybbXWgsWt+ZAMB8rB5+pZ2/dRhAno2QGuJE7OD
3b8lR35/mPAYDpg9uN6+M8ObNyY+U14bAvFFnOL+025SJwnKLnVhADCvhZgPnTbq
HrEb9G14MZrdBrVs1A1MciaD3QFaxif8ez0Vl9Dq1Q/84BDTvNTVbiEWtVamBknL
vjDCYnD1ciu5SN/n5oGC5FTNiVKl4kpjt5cazobkLDWf6ogzRMksha1ivVxXJ/JI
Tckw+X/N8rLC5hHKTuOlU38BaTXLrI+lEMg1PVG7IEgrI6rW/rnpoXRYg+fgfyS6
nD5/sTP4EfvhRZU1X1nu9pmI94HX7XB2pkd0m7CLAsVeqCBNPlNllzT97eDciSbp
NfpF4hWFKxUu86tNqJJ1EDerrEAgVk3PwJsrcjNfcgvn2HbAGrJWV8CW8Y4E5x6f
4Q6Z3zFtXGvOcQyEOR3JIMuMUwu+d8tdySIq5tOP6EgIgTDVWaziXnyny3wYELWk
R1HFO9wvoayqH6uTdPIyspnDukA+zZPNVwncmpWg6m2NG6UklurD44mAACKZmp8Y
I67eDNnqyarxPwW4DYcABe2fr3AfbUHv6MXQhCiN1ZKnFX8Bpq2lEAHI3+9zRA+y
RLqkdo/emwG7wkWgSamYWWIPJ0ak/roq9FaukgAIIpQEpx31KXiQJHSU7xBWlPoY
nAQ7w1ZrL0frPVIOUmANUvHB9ui7PtRnlw7X6j1oL39I5jRzGRKAN50eyhCO08CW
OO/zHlPwKKXSABe/pT7KHkBVl4vYCdG2sDZtPaCyxfiBATUdq+FWL+vr2AARxz3r
mZpMdWvSXbY48NeJLnTNZEShwI+0AUreurUB5nyDvlUSo9DESHt6U+DXuI5E3VwT
lvxt90SD4ECKmWgZ9wMfqB+x9R6ihLgAXFzA+BmLvZGCwXF3fD6Nta49NQkHJeJN
i6gMOMpP+CzDLGpMU0DGIjJ7g0/TZLMiWPLIvghMZzkOWIr31xQxIPdPZWBDZxoI
NYlsYpwAfaKXRVUSgJ+ZTTEa/dvf3D4EhTkuSiba5QMWMFCQ6TpSWMcW+KMcn9Zy
f8Q8HgSr/377H8xNliUtxbHcibFxG/cbpScByA0RA52mw3acy8QyOP2ocfXtEvAe
//LXO/0HGAAM85XzBIHaAQEVnxvAF5XCdA8UR9cJf1B/PdkKiICbI6xSFfYtxE1x
rA1AQT4zbNTFQCfJlXnxLdxOYFJ4uCNg5oT41N1CDtTjvu0NcrhJKbUWzUwXvd6l
WYgRu3uRs+9rb1pGSp3ZDMzX2g6+FrkC+xD3RacxR+0pp5Job5QQEHsax5XzD3rA
DSc6fTMs9okxaMtQUdBQs/aOQIh4G66DuaInsTHRPi4iufXCcPlSVxPmDSVv4zKj
/JYndbqziK8GFoilnOH5VbGayywOwQtIjptRcLMPUyiRYSS5OAMR2i/R2qljfKj9
9iX3X/j8JZ6thDbGDewqhfmH0HmlusYOcl0/qa5SbMY+FzErEjwJO4JBZupT6ahz
KuqrtptO8lq3UWyaiPozksS9mX97R6buUYWd66YQtlJQUb8tllOq8kOlgchyPd+W
V/pMbfz4YQehPGKSAYnn81jCyAqAOhkCzoAzn3x2VaZVRiTmiyQULBmYrkg4A09a
9GQ2DpVYpkERwYWt9cnkwgTgmhI10Snp/io5Cf4ocECBsIBil9KwXqbxX+trn2xl
TTVALYIbiqjltGckZpAIPuE5ayBlYQHV/RJL2gESgG949Qa5MpBNg2S6iI8GsZD0
LsowANh4Kxc302pafroqb3G2HhIA78cv47aRLA3mn7BMwYRUzopn2Ak4PINAp4Y1
y/paDNE11TMvap0A5xpE+jOJT9E+4q1SplD+qBV3dG6+7706b2O8LkUyco23nSiO
fZrErs1tKR34jrbfu+zgMo2aJ6Kmwzfep5WehGQbRSK/NwaOl52zm7qVffhJ4FYo
RbUTNA3C4G2zPv/rXdfGu9ej04d0sIcIGoIbaodQ0goaBHYW6AUqRg5Mwdq9iOYn
LbNOof/lJGTMXhl4n96ZtuZEjyrtEO+s3OyhxvlY3IAlwSYryazX3WnW3LvtGhtM
MtEIcI2Okuxymmnc8uq0ImKjsxSeeV0KLHjfcB1nYnkKHjsaPl+uUbEuwdiZjKlA
88TXT78Q7eOvbYYFEh7Gf8gWzf+Iim16PcJ5fhteTFdJ5Qy2AZqI02TQ6Dh0conR
/hW5Og6/5igPolcjWZ+7hUpyQTWnLeXVoxrF9opKb4M1/Z97bcA7CnfbaB0XyAoR
yWHrCjyzRkLjE3jc5td5tttLC/JzjDSOumbVvlL2HvVc4cc/eeY3Qt2dZySo3Tjl
rfoonCWiBiyKMTxQbghNliDC+6BeJIHcEo7rSgunzllfmXJ4fd2ACAn0r+OwFRqT
0UR3dZusK3BvBXkM1DeB/H7wMOwQUaDhHQ4jF2G1qalDugrvWJDIRFMV2BUYYPUQ
mpifVtHsin4YQRPE6XDI+UcLEMkX2j3MRRK5XzwqMjG8dmfX2753PjkknN5aBkn3
7lOv2/PbbGrZGbIPvwWPfHLqsDqWtz1wvItkjcPduplDZvJa2bzrpqpGlkLYL/XA
pjCxFRF85F2LqYt3BrJLADk8kfUB2S03P6FXdhpYN5PluutuD0lt3GgZ779jER0u
bCUPrfFzX2ZkbBW18wqboFEiObVGN6WQubq3PuZ++EOq4DDIFNPQPngj1IwtbGzX
y95AbhnNU6dV2SokixwZtL0rOSMR54d94moPbZ2W3CFpg9trE09+c24ssLiLM78B
jd/2A/jd63jgghKNeC5hULVzKZ3UvVHy8eJmjAn28Us0Lb55GMAU/FtSLNDJYRz/
kQjKp4bnE0C8pNwjHMiYc1pXUROkM5/jq52Jz2gsBdMe3O6BbGLOJq7/MlxTZoga
QR499wwG/U9PwtnRFsS/gMhQZSp8Y95dSkzPT0VZdVur2QJqBk5rprZ3a7x5euc1
LJMxGPwI4vGftwvqejs36+LJMojRLqqwUj/EVNNLnigFwTw4AGzE1ZWGyJRpcNqa
l5mM11S8/nWhVCywKn2oU8t6gxe6AEsRTuWxlx7oqgA3NY4w6d3che/RIwwYtZhG
+nVb8y9+7U/JoofXHjS2JJMmJFIQ2E03sBB/wic9PL0T38Xloy+OLEk8tnCxeDe+
EaSSGykUx21Ckwz6CoVMk6MNuqc1us3YQk1wiMI4QL+7rAp8ASh4MYTTm4B1Qpsq
PK0GmI7rOeRyAB6m/6U8e3uPZWGuOc5G+s9jMxMPDrhBqLeIzWOJ/A/fE7m2Ulh5
DWhsxHA6OGtey152VMMtqWvplgBK8nX5WaJr7HP0OLy5/6uKRnKnOZ4wDOMUYtXf
cSWjD0a7QDaI0paLqr+ANkI6n8WDNRywE9iUzT2cKuYpfdpBO8edY+XQgP2k4XRq
E3meKo4CpgAS3vMLpQCExk8KOwEeuAawvXjvdqgCbNFPSd0UcQ4bjMEZI0qJ0r9J
VqXJ52QHmcANeIvJ3/sBHI6BqfijVggjkCQ+ikLcsqrXaeUkNt9Yojk/Bbbb7v5e
zSUO+VdAtmYq85l5g1JALolsR6Wm2AGNsEroEza3lGpV2CthmghWove9qZF34Pyz
7ra5JfHwydkLyjgrj5JGaHDasdgX5L6adIOPpWQ4U9hCJ2g6yMrO3X8GrqSD0VpH
BS9tbZIEtTnUinnZTzboZruo9XaO6C2+UKd/Tar5kChiQCGVLJCqxjHsGRZIXfPq
Sx7X1pz4BcWiavk2uXAed0yaosoN8ajl/XOcCDkDNUmRxdcruBMvBlhcTSlpMocR
3M/FBKQwCSj4r3DV2N5z9VlXrqGvp8R8d3A3f5JPw43yzaC7Hzht0M5jqMAVcPZ7
Ix2opwPOpe4N7BwW6jcXGEY4cxpDkDvhxuU8XhfIXJXIAGpAUHzepHqNHmiRIzrJ
kRxyTk6YIU0pnL+BL55WYohhVYtFSv3c/o7w9h6Zbo8jlb5jQ0e23Nidt0CYNJw4
mpE6n7SXXIkCQBiLoZGeEHkLgPM22CMl6v9jb4sQBnzXxxiDBhu3afo1eZAmYHhW
WkVwTyH4GM3PLjaavJA957+43T3jB2LQG6taQxQHOtIL9wv7HOb24REeFkYjM35h
ZqH8A406V9MNScNAKeqCyHcjSddi9UAB35Hgfu+LmlY7lQ2dibZ9HDgxUeGan0aD
OXzsohBD2f5t1mqhpX5lBFXy7+uGA8DOuhqeLrXZAS8L1YIKQyp3cWPSfdy6VaJA
aXVOh9LxYiWJhnHtq/hH6QnFztyysNiJxNoLFZh1uA1F8LprVf6+LNgIFfr9uVe3
WuWpXcymEZqy4tIwAQSjqOEbLRRykK7rj/J/7o0+VSWyCSr/85Opv/kfMKRxim9n
qrruY6w94VT950KXoQqe9EtfZV1hiwYncbcEub5SblCCja4wsU27P/72Ch+xjPDW
gwUdSJs5G8ccgaIo62ugaBJf/i3O5+feLQIzuSwUsyimFJ50HEM6Gx5tAIy+uzS5
ET2DAZhSHzYAYpt13TzN+TGGNc45aFyslptXo15XSmOzLjSg7aIJmpjecpuLDahu
o24qTFeY0t8kALoAUVX6ztHNdLAbNzBz+Oh+7zYZkJRL40xUCC37KY8oUSVS5TLQ
5xuays42l+9r8+uJgb+VxvCByupfQf/aVBI9Zj9XalvtzB0oUu2qTQTynNpQke8x
wT4yYRHwa2tXAxoT1+1xIOK0IGAPR0gf3Rv+GxE0IQnJMrC/p7Kv2LWZVOYRVZgV
twP3ye6vkVMtLbpoglEeqEV1w9Zq0t90/MTm1S5hwV9K7vahwQtYCDV1mbF1VJv4
czk0UEmnS450dJ/PaRKKUyIK04No4439/zZz/nmz83PeH70z1RWz5Gi0r1Ba++ze
Qoe//hzL78c2/jQ1cR67c7NExxv0K4ZoAwFYmc3MqbJX7449E+Y1hehCac33OAh8
t83pXzBpiVcCQX4YrT7SIHq/bs+OmHErds7AQuPuZZTR+leGscv3tloTMYe/4MN5
wsutxPc/Zi3pNcodtVrjd1Q3ArSggQ4StAk+knPWqnOa62+CPTzRdiflh0bkUHWE
i3pI2K6C39WDiB+HT/ISbueTwuOpN0S520AnDjcM+bs59golMW3RTRaBSuBVMhWD
BXxbA9EG26ZXQ5Y0WP9IuQO1HO1IVzIERfk6linABUBuFR/yLREvJezP7ToUGUe9
zlQzelt6wHN31yarKrQmLbXxfwzwVHEofPQX3y3C6sQmBjiT0GUvhKXCrM3WfVMr
v4MiQPKOBEzCodou+J8yZIaGPO5akj/dQvPoSgz+Lt86J7lBpLMRoegBEOzXAuFd
JCP7ANWRwuBYXpmJ/26ZOiHDN+0ZOZTbZYouF9rcYaRhNCbtBM5X9omZLfBfjQFV
IS4i4xP1dysxfXpEPTbdTvd5eo4/m2cRsK8Bf4cKncDUitfuAir7mEth+U0n8EO2
dhZIpEPGmYhZl3VIjyxQXysp9DGkJktPurzL05ru7/K7miPnyjJLyVtiPbdq2fbl
W6i40qnbVzSUSc12BgwmqjHrNvwhyyf8MOkNCsczvMirzg8vpVYKQmuo636HOrnD
qOoL5GsenXMKHnFvg2r7xFNdGlqEYNBI8RLxwn6o7e/hNaqS4XxrUpna5yz0C0kY
xFiGMrerQ9hK0H15eB2S4n+1qNE2SHQFfvp7/coTReOsXynSGyYuQikq4Yr4Cc2r
YJn7FsO8IiZVwqGfNLlsGUerTc20nudVrt+hyWQJw6OuxJB51E76d0cDCxpIH2ko
CCJm1UK8m+XIhqwWqFhbk0uIRukOLA1nENGDA9hfPiuSwzc1cNP2GPZJVsnbkGnf
8ShldT8phUNHdYIzQ+3mrTxMVLgVVxli68+7j/jlfMDWDC3V67tK8U7hvReudOI4
KWoNAEzI2hgdivYcIg6R4rjmB9mrnmFU85gpH7Ap3qQNOfgiAly+n0Ba19mkobpv
Kt51XPwrxl4E1qJ+AGAnGcLWqqo5v+g0wl0kfxHupNLlkUVBJXeZyV4+kBUyjA1o
U3x8Kdaj0XR1d3djSXCjvz9EWapgO9OVhAdv1Tb6Ctg9KS8I0gTU4v7mtpuxmti3
x5+X8xY48RLp4z0kQufY8xLDSc3EA2o7LcOJlzukxxXhFNHhmqGuuPqWdvQdZoRv
agGKR+nK9uN3W5BK2VoYASaESGdFeJGcHBxrteWEuVGWC+8OK4/pqdjlNb7owmh/
x/vFiG/HGWF7r/cO5gR9WS1MfWZ+KEdvxB2xk+DTxVFo+IC4ufQwbsuIgiwPdNHI
4zsmDsm/GKuOLMtFtkD24ad0eyTqwzJdwoWKzAIqI0Ki5CjtJNiw7lOd3hFezYH4
ndsZQz2OYsPYCeVZnETIMRp2ip3nTywPxp89SYOBNemnR3XHMifCAqWDLRap0pUJ
qpCJVPxhUGaxytukaxoNYY9qpl6aXeih+nquOL09w7Io5nESyqA4CC1FVCawnZJ2
EgT4zjFA440zx9H+fwyPd0Gjh8Toek2G5VHdn8tDJRSwe8CAebuyQEj3S8uxFi2B
+5pzysq+WggjArdQ+m8eU/lDVxiGdAbHL5ZW54WYNCZDf7R3jywl0BPAmH4IKUua
Velz8ACOOC5B5El59XHTcpYwGhaPhwk3FGEZ54gaNhb80ytV1NxGvyBqM4DIi/XP
bHvXsAjKYhTAjoKK1nIamEGQ6UVhuNsLIAOkbkVgzMXyxRzEy947KIeOCpposxqF
LlxAorjrcpC9TGYIoU5N/87ihNOFDgeAiX4hT/GgCxyVQKpMYdy/2r2HPpSNCuB8
dBzRI6X3fLJ6YLlEkNUx2kaLD3EzHln9BPZFBbwdUnaQ6gltva+SAqwGESPoGzlt
+Z26IFM90i2lzGkW0vjF7kIao+nfmSwnLFrBgNazIZbPw6fMtVYkUuZHQyUhFzle
R6nlGTHTHcjYdsjc4ll7qWzVWN/Fu0+s07PYaFLR1sHcVuatbr2STzwbGyuan7ZN
M+ZHNmYntGQ/tGd8urt/fm+VR0FNaZOQRa+4prjNlJhVXjtxYw0B0ssSK2yB2YV0
gGHPak5a09z5EGhnE56eXYJHQYtSO6HjVl45GRpnkkiw2+Cvf/YOI5/IQWmGuWX0
Iacl6ZKeRm7WWsu7yE0eAI89yikvSLOwcYpLgfqNbFmZdUi/96g5y3YAyH7b+nA7
o9CM6CJRUUH4grf9mh6ysjzmCOEryV52PTpzg/MNgnHbjhp++wldH69BB5sUUnqD
A6IyRhDL6MJ3u+I3MowCujcYK21UReylex+oFrtbLyzNMuLaa4R4CVcL8OYc2meZ
LlpXaEl009/FQtcQgLc/OwtRp8tKAiDQg+in95uja+SNEoLfKKKNVTbbpBv/h8sL
lHlss4l0x8FEVc0XdHWfNSKHO5n9rOuqD4vnnjmk5ZJUb1u9bRUMZwFvsjL7yz/3
za6MKtp8sm7816K4KrFaD7LlWhTv8yXK7Gd/U6qBnhLMho+SJ3Qhhq+B0AZq/k7L
PhWbYa004fLhJSbdmhzyZSOfV91HLYD4Res/ZPSdNKJ2CZaVSyEikmTHewPN/sUu
qzzRssEJ70rrAGCcKkgbVe3L7Q0DR9/jtzyjREfJopuqwO5Zix5wqqhEo/WLkTjG
PXbUom/52qgO982axkkKRLLdtwvLiMzWlPgVtWuhVIUDC/3nCOw22p5hVH6dh23K
l8ZOglfrtpkqOTMdo9V6CwG9InQzcQY2ljj5flMhPkjN6XnKoocEKHB+D2XfYHpc
F5YtvPkBS1eurqpiJbgKjOREjJMEkvBBP53PrF618zLgOHYyxiZ1MXBiK67negpi
yj3vJE7w8nwRT/y9bOI25+xGMkWwVsh0vxQSM5I9VSPztWrVMiUf7TzAxN5pW25H
zP2SB70JA99VS9gUHHoCCewVoI2hnOs2U+x/v+SNDdfv8g4sGq54Xd+ubrM6w1yW
o/pbEhg9ylf7W5nmvlfsHA960gxx0zxPeMYZkzzea216rLDUMGCufmjn3mgvGSi/
MMlLt6oMoz9lJi93nktfIlyrbNuSb7agBglbk1VhLsqArvNkZovOvPG5/5B5ikko
cRdikjd4v00acxp/otWGB0BY//cFNZ3hqHCLWPjI9624YIWEi1PaVjlyBENFK7iz
VZGllMTL/AUfgkHcKqyRKODwrBSMod3lR7ifa2+ot8wyzbdXHzv23Nant8lnNnYs
feRWmuyHv6YzfbRCGf9S60OoKXfguD+PfoIxXUQbDlVR+kBrLxcmKUArN9DtuqtH
TZnFWTAqgCtgLQGogOLpJc1QPJEQaCZKm2sI3PVxno+Pvmmju8rl8KFGjrPKFPOG
O8J/RQ6N4oUC76biI6QbjDLFqr9UKuAwt2gJdGps8dGs4+N8+12zDGFHDQYUXXFi
FE3tzfrv0m4f7upYoMydNLgt6SW86++SzbDaSLT49rnGfkW3HBo1e9QaPe0FK2a0
OfGpnMi84zNhNRTyUm3lhmKrKVpEzUzyZSuhqQ8+Kg407XgRyZQds2QILFzwjeFq
Z2ZksrG14EotPSjlt7AfgepoyKQ2QYRaUUnuVGx3vJGry2fc5+A9a2aLyY6osQG5
aH2tgt6WDofYiSy3V/S9DHd1c8Fp+jUgSV5TpaDKfwztK34AWwwClLvpkHgQM90Q
NZHTeHTXle8psPOrXqIisikp0WglD0736LzRU7CBPn3Y/riuNMfpRkZWjUQSf/PR
EdWEcptugG9ye7NkepEY0S3G3WSlc/iPual+e6+sscuG8x75EeaelR7z0lCeXC0M
CXjsPldtzm4rVYA7r3mQfD6WEyuPbna+0wleG5svzl8SELIw3TQLODIWBRvzanRT
OCbq31pYOalZZpVOqdh0dEVPFAZikyaXKcPYyIFpv1u6g/uFSF24KyGVv/ZJv5Bf
qe95qEUj4rrhZncFg10YFo/2ozAIIxXZxUdXm6NORhZ93iSVNh61QMLS44AzrT5n
XRUTCfMw1/p4bHvGo6EC+abBs/GfHzrTxaTHHhOzcF2xqx4BQCOi6SbBdxUEj68h
n1pDJxYLsDTri28tWQpowP6H1yRzzillwud1j+NSpAnm9gFO0/cVvBlRLxOrfJzI
BU/vet9xXWv9szNd+vQPxj5bVlxRsDbDc+RXPEALIa4b2n6I6shkRgNzfIAU7R8U
GA0ixgCSiSfR9dcBRnvJ7k+8BE96OI0IjZ8s3HLms1bi7dLtthdG7niuYP1v+zNp
INcXly/XMYLNTasae4J5rO/Ulaw0SKzTVb2PdSHDaFclup//deT8bTmhdD/o7HUL
q8c1GffZb6G1DXHW9fprkfAofzHZusk3gUD5ggWijII80UX0MAumfCzrVMOaMf+n
c90dSGwA1kY9glGhjwfBv0yqq+5Hoc0BYzGkbEi52HPdPdHZ2NkF4MjYSu17W+2v
OC6DgF7c50FEw3LC0c1V4ZShfiIYMVLHc/XK0FM88dAlD7CXadcYsi+jPzLxUfd1
wHqY8rENxY262kNh5s52BMtqGDMueyLVeM66ssboC3LIZEKYJrMikUysgQGCuUiT
v1jazKt2otnAABeyRUabIOe1Q01e2bxD9y2Je/PGnbtA3QbNrcZlsgKrztsDo9IT
MflLtlj6KYnG0xfY2k6HwSQUlB6DwLAncAasWQ4cDnNgfscElwA65XdrG52m71eW
oTvwI1W9UXXmx6J+bM0evha4EXrE2Obol5M/tQIKhA1tN00Uc0Q8a4T2a8zBEgZl
TKeMqF4z224H64kIX5BrE4EiVvd9K0Y3+I9UsmfJacBpn5HUAq210uud4GZuld09
qopmItrIYbEGYhcVFKxDp7nys/D9AvmTS8FXHS0MXpIqP0RglRi0QjEn0svA/7IG
BWEzMd9JzZYUT+tUc2eaKmtgul/C8f2869n6WDdwCK7fgkz6xyX8+5TzVfAP5Fb6
q/uJdYdxMFKFmJY+muJvj9bgbATSiv2qutQ9q5PapwlHDrPSMmpXX3VcaynNH6+P
morJtOaGRpxQ0FQz8i+By9BiR5d1lHKXc+RyOsdkKKu73k9ieT8ollk57s0rVum+
xeeDnqsLk/5gPlODylpz4cm1nXgfxZc4SrCEfhobHKNFQR5kf5bYGHPOwxK6NBTA
rPBLI9ZwxraoSfA3L45MKXeVqbUsZkQCoELdl5uXBoSHYWpUHm8kg3PBNvKF7LTq
8OXC5u4XmOycgs1/8sQLiNxj4iNazdczUrSuALhUu/aRpJflsF0NNlSKhZ3UQh1P
+Kmqqrv7p9zcO+s+2YUM0yNjFcGZyDcmFIgyBB2kD3x4LOYUNSGkB9HymIDGrkJI
xMJ6mBqqINfoLXMMuIWltL1kkTLj8TZhiThBSiHECks95PVznt6QGHcarmRdQBlp
ybl33amonHXHiYUlZtvHHJN2+wlbVgDv1MsrqX2rqNbxw8kLX2Ne5Btl0SsDtYxZ
1AWaVUUjK8UyO+RKOtpUn1w4kvouqY85oCI9I8MIcNCIO7MmzwHae+0qQaK70Kjl
v11XX1/g8Y8OdhTpmvm2gPRDfZ6pqdthcm0GRUXcxOjmH19VdprhtL5ztXwDC+su
UJdoO7Br9EU7fFWcJ4C8ld2MSNo+2fjiWg8pG9azDz+Z7ffwRJ5U/5sDlQMOFVGc
UnBW8QJ1Q7iQjT6tC4B0Ww8YmVIugoc0lzSqn5RuExXrQEwjNhoI6vRpH8syeN8K
UOnoPH9K8PCgubglqHH+dDXWYshB0Ml2yWYKxQOsyMiFROV57yrZiFa95ToxmS3F
B91aJWgsrBtA8485/eOZLpuKfnpXzR+CJAP9Q4ZCtunXhWC2fOGTEn20VMspAFKS
bCWuv6lQX8z4d32hcKZRID2viyaMZWOMQqrK3nrR+Zhei6hhNnCIr3+W7wniZLGf
xjG6tzBdDJGAEBlwSuj4wS+/rD1FFrA0In+1DUKxpL/PoU/PBlbXtsX1rhYe0JeA
fm04yrZGjB5PD68bxVnJ1zvtx0biyj7Vje5o8GQC6JFhEM51uSeUmJtMPZdrIHdv
RG7nrXcb/vYb/va6TeEiqANVk19zkR5/k0C9ei67e4uR/wU3cnZ1DV6plOXFnZAv
t3Zj/sq86XGTumin7f1qjDae+26aQNErtAFLqCM7k0YArILnZX7WfLYAAZd84R3w
F7uBw57QOGJ/Cih5MRpJWDUhbF/Z8JznOq/4h8lCNdDqgNjRRi8sF6kNDUsqvPlT
4VJxkcBiW90Mz0cbFYMVY+RkNZNMNashYOO/5khCv9yTClm+mYZD7ijFxW0G4OO2
/nXmhjNz2sluTdjZy9PIRlwJa045UY7fZ5WurEhEhM2mBjy/J41DQaMwsKOLUdDt
2z44TIiIJr7IWxegsGqezXKt7bPthxRxJwmZ+9ryX6DxHexahhzExmNSwTWS0iGc
sS1Zaq+sWzou7aanI3QFh6ub8aMmdzGSwQYUsiHL0kDV4uGJu6BDXaMo3runYM/M
5X5JH10VwbHV1c9JykpNTvcz4U5qCFY3y+DyFoGlwlQrbU0qIDoJ4Dt8fyAviit+
Py7ob6hqqdiTEpJU2IZsQGQiTe1KiNigJDV2cYnCvsq+XZDGJTc3U/pwEOpiO7/a
B1kyJM296T1sMsDYtwTbhmU8B5ov8lRtkAmhj7UrCLE6HZRRU5FAPFmZSZtqcgkG
O90btmjA0vRLgeg2rShdeRP7H1PmWyD5vkXnhTCsgniBohrlwnBDTBTPCBpCNTTX
FSZIwV3xptgd6+9SdDL7aTvVUChH+I9KTxILKwubm+8pJG62rxPOB3c1/ZM1SwRa
vm5NhgvogILdJtsuVTfl5HQ5vBw+tQZgPaO2wpFamSJReZ6wYgcGBLJPOVIIdqh+
YyLpFkLmOWcqz0ACeO2SiZQlilZFIoCz1Mjl1xKQ2nWm+9L46P7rRgPiMx+LxOh1
QafodUzCNSO/mH6KzELszMfkfeX5l3l9oSrT3A3kgcuByTG40jtCyFwKFXA3n4S/
SSfNsQ7zfV9zYQkVqYEcKny0LMIkns62NL8HtYuj5EwBf8vKwqpdEklgOZXSoX2Y
ReGtSHtw2s2DOB1z0xGcuOgfqGIbAenvpHzB7kpaIRLF3WVq+7AUyWvBpx0MR1Aa
GeN2TE+8DVmW+kZozN97g6t3cOMbSl8OWgtWEMd44swQM3Dl9du9EUtME9Zl43oi
YO4DeiwwCH53dacWBNs5ixmuY1mNAxptj9V/hXC/VhidugHMfUQmaTDLwNnd7sFW
92H9Lzu/G0DoRsSlZVSRsYCCEVo0BKfT8bz+ZfKxXiPzvPTyBPBwOw0mFlbaE66I
P8o5/d89hDhU0PFcDILg61i9uD6eY/BTmaMEYNfoppXyvrnt5bk+vV9iCTIWxSbC
0sV0rY5jmY+9h5SttuPBbOR2CDw15Fba1nCdeBAWpJIhT0+8VP8O97D2GVlw1cO8
seX774bpicf4GHp/CU0P2m74j/Dwacx8IOZHcrdHV95VYzgPh419aOdjNPe+pioy
27v9QeGMLpZB8tEpwTZq+27ni5ew0f/YOhojTJfMEqpBxyAnkN7s515YRPpL69k0
8E1Palo641KCIn45B8MrC34Rsn9tg8AbI/AzYtmMA/I5tEfb1Eel2rGZuBmk+kHZ
NvkcBmcNKyf8zJON2QmUXN+vjmuqL9Y0GgL/Xo5vn6dGWtgwl6O8UKgH4hnntAnx
UfSWdlwK/4s/vhFX+HG5tpTVVeHx1SRzDMyLQGbkRXe53NzQoIZP2GANOtYbn/kL
NPt1SN9sP11C0m1w6BVL42bcOlNKOW36xbMzbjzDJNEc9KMvqP+bq7KBAdbIMLsP
iGHBOK0ePPUhHmSUQz1jkKMGqVQ8hmqpcMIQTR7ePznHMh6r/bE8nTBMtKtYzZ41
Y4T08pK7zpcx6n8FWaQhKc5+Q2+mmdUdnGtsMwsVlnflQUoFK0AlWmgGAwjESitM
iTC8BD/hp+036o11b3/45G9/we5xHAPfAam9zCgG1fgcAT5rzVl27PDxwJfAMAlu
Y0L4t/b7RPOfd1dU8kEjAY18tUfEY3qyDIPsNMBMHF2DFIU9Gdpm0OoCX0739FFV
rq/+/erIKS6OlTeI5zwewboj4DlbaCisYnLBKAHB8BE0Dza/ZtO5o6hU+EfFbVpK
IkvX7lskWW3BFCd4pazoG7u57NSoyCys49toj35vX5hmT9ExwTDhjiGmCPJWLgBz
JpqjMDP6Qn6FcVnS+OjFXYsF+9GbMIFuAIXLyA+VcGuNFq22xhDPyvLsd9dwsvJo
4QnUYyhvZ5MnpwoY4S/SpWZw/zT8v7CM+Owib6n8LVsE777sJ2j8c4iw4c2mlJeu
ymXEFTQnZZoA4Um94Y612ExEmV6lv0ZSTu2Y/a+/D5Gw0hCkyTY/IvqCxSKERQ+y
N5FPCM2aHVVLipFlSXZYUp7aPxydfJoGv+4SEwRPgDh31xSH3WGqNLrTD/ubj5NG
JXiRl90WbGQSdUr//+eyexu1PkcGijQlYza0qceZRS6KDgl/nFQRsslqso+7F6oj
mvb3fvTxy9pDdf+furB+vIUIj3pRICvpluELms7E1QSvEGeBM0stpalTvrgpgTD/
YH9oPmh3IFqfCEyuNPTP80Xg4dG8kUyPXVx3ac/Tcm7Kd2KrseCR5Urv9/bYrUqH
VBHdRXx3X/DdC/HRJMGlqivy2HknoHUbQ8SvchBKCMCVf8VhDH+LawyC6D/lNB5q
1KM7M0HX8UZR7Oea3p+eTqvH5JmLe7CoeMPJjlP8w2+eVPJtgPrFz/g8flDZIGZj
XtQ2/4epFVGtaw68DX+3n1VMzc0lvxKuYBz13CreG89u6BHhQL9G2RMd9MjJNH3M
BrVpD1cWrOvP8CHnpBgwetLCTL2Qzlz1lZUrtK0imhcJjX/zrzJY0ekzPNuevC/w
Pd7UzOnQic2utAMmhYKwpMNtBnXr/82RRKG3l5FYGbQcfB95wpfckN3ov2dLWL7L
UMvZ7XFW1odCaxyRfi2F6EvWEto2y59+p6n0y+W04vq9YFp7vp+m6O+z6qlUolqI
2GdK4r0Kf6r5uqZZ2EcPIY9SQrHW4h0EW+h1vHkan/IiNA5DfRDdVqEYjxPqm6lM
+ZfLs1oAcxL+uSVEn9ftvufVXy0FJEDpS/yQOZoO5Zmi08+ulg9QAael2sLc7bc7
rv1ZogIdJV46/8R75HJ8E+ZJ0ceZWF8/bSlqWpzQgcCD6RkleQLmCyTwlry7cFRH
b6d9Mi0CpZQnq1NKc8kaaDxqeUjXsG5ab5O1BymcnD0R5w87LWvcD0EF/xpzssQv
Nowj21PXY95FPi2/vYL/jgVTPaCHLDC8Oo4DAP122abbyOOSoCTgjWYuaXjx7L9i
byPivA0EU9eYbihCqm90VHI6ErojrU/bQqzrksKiZvxVCFJ12MDnm8fAN0DLG7Je
qE7Z8c0mXqOItfz8fSN/pH5fUwKRO0Xwdm8km12pF0RXYwIJ8vWW8bAfi1MjybJA
TdvZb4TaBSesKE6qlL01DP6XgTCbNeMs4OT8k1UAPfpMEwNnQw5Fnh1B3lbJ/WTr
8WsRLTCy7zHA1DoIWloTbnvcu+9SEJZamt8O9iqudiB0ONDbQz9/8fcyRKqiyLNS
CAAbXZHoYztVAzZCfQ33x2ZveC8Z9RDlJvZ7vIF0D6Qt+vS8S6SOU5QlgAHp/LAO
mo70+IAaWZSVwzwVVbIWol4GTC9ScU97rlOwx+vAGxxfh3fTRdpzKMYy5EmoE5Vs
Si/yeXRnQ7JMM5WdekqwzQYQl4uj21ojFxwlOqDh5RZZqYZl/eIIrr9gPlNCWxcd
/5loecH4sfUtDWHEEb4xYM03x12cCEmUWdE8z1FaW4dY4s0FsZrYv4aTkHBWaQPE
eRRIs9ZQDIiSXG14UOsaRxaUu9og6fg+QE65NysQ6cTSPZ8UvKIT1pRO7x9mhzac
lKgTD+z34tSamojQKnx1cWBl85LZVzAbhss/Mz9+BuKzKTWphEO3QC6RmvlDPeb8
bGn7u5PunCla7CCIB85l6SZrgLQ2xMse09oKgnnuM6BVKbduBZZlgRss2KMCuyso
afdmkTm60WcepehJXihV5iaaA4BkA6xc8xllbhbfzMVSm3GVwR8cc8zw5gVRvJAP
L4z6BoT3U7yFkp3RWvGCvgkxc8ZXAsSTfPzfnpLQDHpdpM8eaZxNAxzusbbtWZbl
MdJtayKBF+lAQXlaW09m3yxmZU3RpmPuMSyWtcegWRJyIpXWmbp3xy9IM0mqDUaf
3NE/7xTcRPfLfWrr0B+6lZVY+u+/mA/e6ARwvzmj9GG3K0N0eqhzKZLEf+7AdyRk
1U4sQOfLUIdy7afQsb0P82cdYGKCPGfzw/nw99kKyzsZIvABpNLM5pYzePq8/E6d
2H7z9jDS/JqK38Q38XpNod3+CyEcB22ZZZsor5r117WQrTSh6YqMmEaLPVjn1lmI
aovBbUwuaMAahp6Pbi/s3wRSl/Ya/6YvWbUETWEm2wpQ7QFZ7yL01zqCh3w9SA3q
MeREjMdj8BCm9q0ZUD1TheLPv+akmy12x8k+hdLd7ij6X1Mv3Fz0pYrdREPBupB4
x3433ZDFxa7dVLh6YPZGB9468K/AkIWpK9B8DcAgDOIkzjc8m4c15uE8lu/U8Cnj
e5r5Ezw4qjoxVymG3aZZ16gGvuheTr0G0xKmr8p6+baHWqUb5XGWpZjl8l5Jw2M+
MCHbrF8VvYsyerArquHgxrd6xL0E1mNrIbTG2kW6yHyi6Z6xi2XhVr/tRgupJfOY
jAq6rkvAPZuGrMWCS+mY4G2be2y7WLI+eEE25e8u3GnFpNeLBrO1LeWIZlGDvCL3
8pNOaQzyV00/MFyY+xUhoAOPTy7v4Drym1om8DgkENVaLFL8BTMRoNASEx4/+zRZ
iPBvdBz3cgQAO2vdLWspLTdjtPBbPxjmFntpNoxIsr72amOKao11QbU7zsPNaINU
Vw6iT8AESebF3ZeeEOzXkeSegIKMbeUJECnssp+6XzCxO58hPfsGy1GQ3HoRWOES
AOmXvW5wFI6XNtEKZSx1/WCrV0eQLJOVRjzskcmLthj/Py7Pb0KjJB2pFpFT1vpG
lp1nKO6TUXtBu0EyuHDgM5sVYXR105XB0UE++YPZKIsrNAX0utKNuEtj8wcVxiqU
Tn131pNUFjNxCOOfSOHIF9k2j/s05Dl8uLdlGg1NoshV0FP8p46wx02kWUKTefPi
jUWwXr/5Lg/4U9pm18wiP3znORSckdY8b44pgmn6WjDrVyjS7d2BDoWbVsW2g9N/
Lc4HdGAT2PQ32jnPsDR8NbMwZx8CZwkH9IZeVy/nOfjDqbBl1Iy5GjalN0BDWB6l
152roIyOlYaAVip4bzg4Ajo613EpEwcHpa2c7z9fqyINchhVkSRASpjch4g/Yj70
BnT4axxOwEL1rt77lnUIcrXOcsdCqLNEUQBJBZ4jcygjjiVwCGLAvpeiKNOwf/5L
o/P5Z3himQR19xK3C35sDE/xi4VjEpMVKl5b8QOHpTa2rTRZYrva5jBaF7Bf0hoR
pBZcXeI7fuUijA3GUW1K+oV98GxempbIpxbP6BjcbISd4ZrPqkq5FbLSMjgIMewg
4pneQlwxsbmF78rH8bTVCeyAxfNxlIdNJ9Z+4rSUSh9VLFgplDoZ3cnjxy/dqQLi
O3bmR430wLhG10qmdk+640IDgcCpvwTXvi7Mkdvw3JK7MHJ795tp7kXQtm2r/E9C
zwJw/CSupj5XWIQm0g5v0+awLV4WPXqu2XclSxE2Fi+UWFXy19VtZnRa0X54oTYX
IOSmc26Jb7VcWD6jd8hKbd+sllQcojjhpNlBdCooS/i12fJl9FXE2JifYpdWySiN
G1wWrdlEoKJqKe7MPKHF1eSNE+hE5OVmX6PD65zCO3om5IqG0FfsEsTbU9bu/H8/
GyrPr+sLIWA00DsdW7pqGW+rPo47CXsNhwbGlgCNmUIqPVEUf6JnYdfX+IaV2hEl
a7CVqcHQgLl707opM6BQv0yhbOP5Oy3AfP8mt91Z3Xqu9+sf+QZ8rh8MtIZTx5b8
Ry0WRM/hCQfRVZF//POQwrXxoL2y3w145JNjAy7liV336p9LobQT2yEJYVIZdUEN
J19Ncao6H0RNRTpSPULa08xcMuSQ7NCr6oTPvg9dxclZIkLuiP/pxXunp1XRgUa6
ZxibkqumH3aGyHk3mUxk0IWocXzDFaII/73rXRyR4+FeP8PH13UQ11WVuhSkjRVf
jK/Yiqspaj0KLF6ivV8wcCI0j82GLyBtVysIWHtn2YdUGUdcjV4jxkMYb6/+o+TY
fOqwKp7A6IVb7qmBeYOadcd49xJnRK0lScZ0d5C0mDzuRrKs2DeJOjRaD/B702HQ
SyH6SuaHjHEcxeOjhpAr6tVPtGlM1eH3VdhDM+tHzqkfVmRODE7C/qdYlm9ClB7i
6tfkaUJzZDflsrIkft5YGb8bwH8m3eVHrZWSp5JgFkvgsTAPsp0/VmP+S7Bz+0aV
/54UNi5/5wdI8RvrExUmkYgW1YMMq+osR6xO6xuAnR+/BuyulddRcFtoavdYQnAc
yEQY/OYr6fBqGfXZBBZKPYTNJ4nZewvqUrLUbld+NnKC2/pSXucw8xQh3zfOCy6s
7pPvCPuaKM+54uNNhWUzJnvFywgMj0NhZpSceoISl7t4ra1Kocm1g0V+FW5uenH0
VhrPNimbyJS3/UydDAWMxZ+7nk/A5+/JOuK/JkPitYuqgAZ46NQIuh5w+xLUDsIe
jmYzrUT6agxPKjQtRRS7Ob7cFt5wPkLOHKWT5KMxqEqhTpKdEHoBuwyTmMA8+7BH
pxZEiq65sjhvJ7Ek0MLtifG+9xF9OJk/0+cSEm4BI7sSfGkO9QJkS07bflvfS84Z
pYdIf9Xtji+RxqQfOZTudflZP9yl3CwZbN07LAZErOKiCcSMA5UjjLIaYXq/4OQh
mFY1dlSXBH0r2gPzfyfWTCxuyHHPaQt4b78HBISSKwmmX07vG8pufgT5CXdhN3Ey
RaV/S5Kamdd1idZfPZPlS5dJETnykC4mK3oCS38Oxkna7CccvRWrUVgE+20An41t
HuksR8KypFa2z9qXWoPErVApQN5mzCnKC7DYLwaHwTbNwae8xgJwr3YfQyuTXXHI
BIPhJCWzfpS7Bm7h0rNEi2BYa0iA0M2GRPaqtZ1JByuwumjopLufkm37huW4HPhU
Ey/IM6NQtY1pqFCxncciT0pqBpF3xRU3vwYPPbI93DNK8Z8Ijwkbi4xlFclHeKe7
BrtEqM3uBX+xp+KG7l7Hl4RKmufAUE+qyes2PbHfN2tV0aXxN1ZnTV8fHNetio1S
0rajtBd2s0vUBS53AaV+aTn6wJOhk2//I3STdNFghN+WeSoiM5JMQyli5L1v//B9
48JR4XkKTiY7hKMELZfAvQQqtqVc5C4WprcofzXzmoxfMTAzEtW2t06Zx9dWY0+U
og6c6A0tmLxAcWJ9SBk9xjTFzQopL0jrwVtazKBlo8foJBmreNCF1bfGZXzuDsA7
1P+Sx5BoJR9XMM2MFZ4FcHblI9zP4A6dg5itYZpMl7FQSJnqdNp+tuSRfhgiJGB1
2GpeYzC13VTpbKIT2qmdu1B+JH855XM6/XqjzbZkTIszf/0uge2t+RviK68nCvmN
XZDsxdCGYV3uQ7NsSGfmtCOVqTS9d2NtSiqLs9KSdruuXfGFffoZtUX+nF1LTk4L
hULqTNKGw/6Vt/GRohbf7qZx0z4zMkqGdDBnowDRgtOgemrltcLw8A1d9+y4HLwz
DHiAxY/VZ6jHLrRXv0ZpjHcW9M6jqrzwn4kOdcd7amSeyOG+ZyHrz0woVg5Tzvf8
yAm7ojdQxMmC0i1TquzQEd0tNeaR/KhizHHMFxf28K1w1C53V1/euCkSmPMnh/wE
1EbxJNCF6vkaaWJAFBkv98vWnc6IpX1mGaBAdnP286/PxycTZi9YDMfySPs7SmLN
hik9kvpXoqcMvt4Fq5DdzFK1rVBQu5eN+lGA+lBIb/y8OGb2ICTrtdlPAlP0CnBq
fOswOHO6TxKfgvAaSdCVB8cYLcCjb+yi+jzTErH+QT9aezlVwy1Uctn1biAULBSo
GsID9rfpidtHMTebATphGWrT0H+OpIstiNdAWYqNh3KRph53fFnOkD60/2tbiTw5
ocC4zojwhpijaBHzpkDO34X8SxfifcZDFJnwsQpY3sZjjD01qMnjCqjLvwYw67Rz
0xy4UrryV2c5qzu2Bd6rRqDb+IIzwmizzhrjjFqWTn97qcday5wySfiNo3idrDlu
Gm4vPQ5v9rJBZrUMO+QOC/rg7X+dXzfbz/JNrosiRP2rOPP08TUCqW1sY6S0us02
wzRkv6SF8Sb2jcGvju6ctDA0SFxwA2ZWGslwBiZKqRGvuHg78YDV9a80omQRTnIT
U2aljAFHsQeXrxT14yqTUyeWg0SEcLac7jjztz197rHd0EMiblk7+5rxifh/aFdH
MvcmPsXLmkKEKoTUadN0PSrhOp5r5dhuzYe8zAT84Nb7O1/HHfGUO2yBqXD5mYv8
iezoaN3szLoZLO/C0IUTvA13yPJqg+t6qCiIw8P6HD8IVkV9ThGcJH04POzqwuXO
cLc1CVXcSsvKyW3QXl5rL8Mkxx1pdNPVxmYkurUvxTa9ZgpHgWI03NMvY9yPHSDm
N44jaKL/AwSbONoc7SblDfI2zsc9BFPvfpMzGVrWGWEfgUw7dkuCWUBsNJlsiS3w
+4yoX+qeBOk4LY2CY6kIBelnhZ+iXC1G6QuLcE65ejc8AmLwRFdtYomZamSro4xM
Y7MRRJlG7Yx+njwj1J+FWN2nKI1JxkchyW9jnp7B27ofz/IC/BHUgRfHaS1sLh/E
emCLPT/9ls2mVXpmE42mUu8vaaWuX/J/W3Fdky1Exugpdgs4j4IlTcvoHie7O6nV
n7ya+VLLin3RH4t2mHAkMV8y/2RVmt/KdPfU4Xn2h7j2VCUPQtKY3ktpfhKwwEJU
Qu52tZphRpJ2QJmcPsI9/vu++p9yeI0dIHLVgyw6qZjH//5jPZMmgNc/poD7rFlv
z/HWArY+4WQeeTU5pW2y4vAbwWV4aJM2yy8wNYr9evAFYcVYws1MQODJSMJkWAOe
nzQr8OGLBVnz8XBNs35CdlXAmfglR3RlstC6xVNbFT2E7PvHuYlhHOy7PZQEzL1G
iredv1007YxA9TWqNi3LFNWPaCn/tDiz49wbU5kFnw2nUCFTv6iCaU+7NdvKexzm
3zJw+T0IgsN0Bc6ZkWbDuuWt7LRJy9dY2xN9v/5aViN7EWne22i2gT/EOy4OBFQp
HF5Kc63xBzZ3Qe8ETUUW+S0OIujiMcVCVQtkh9WhpnfWfa1F8bpsf+MYlzJsElAZ
ct/3prIbQiQXbafKQRSp5/v6z94NX10g8myIi1Ddb2PJbgrcT09/xRlad22CWggt
sQsqqx4FHayBr2axTzk+89egoJHlr6gaMAKaQdmT9ELopdok83vVBuKVWGU+yvvj
eGWTyTsKsRFycwGlGux2YQYFxDmvtrcOeantqrJuwSZriXhtmCr+hBywqdln10ja
5Yawmb880r5bHin5GloYq3ChwhmKZsm8hGdauS9pUUKPKNwOiFEoXG9RKeBUw8ua
+1/JlEGANdH5IN1OIoHwBilcb4szbCLROnqDxCumhS4gi+kQOO5mA/gd4KGm4Iss
efXYR9LmuRid5PLnegL0dAc47ASufkO9mwtNKk7C6FgPuUjOrex+Vf4cVKFG2lOn
vb7wv33kMuGCyGuPRg0cHDp79Ea2R0uMeFUqLmU7QTpYRUhi4rCShUr4QaVxrYgC
U77E0u9lkzt8fn9WfvDhlWupuOx/Xh76jULitcgJ2NgFm9TAYn32qGl1B8W7rsjN
p4pT/2wtAt22lOpwrnDE8bEkYM9lXeUr6B8j0+rJnyC5yzSHKUKzUD9T7oPxWkHp
I/LJYWdC37a8w4iCR/ZZD6dUD7TXP6DM3ML94M8ERDb+OfRVSKlhedbZ3TZDPI7i
HYBnYuZOSyDKDyYlZhe30X9x6FyvZPB2NLQh6kqV7Hl9OIkPZck2MXa+UzgoIQIS
jidSZxQcAw1oQBnv4HGOaP7+sJPLSpowIF2hF7IJFNqhEGTEyaJS1B47tvcOWhfJ
8Q7lX+nVm0FAUSlAi0VWoj+aC8AJyyst+UhjYInuMT3q4gWM6AD6VAnCmSaPd/MV
TOwPOKzDqvx4h0gPMJmXLGEWuQztpq35OMEuMGEoaBF6UhKBOfAOwH4K8iw+HK8+
bJdPP+d184SjM29LxUfuEMnCv7znGUtpub+DofZXW2Fry10jRec4MgyXmOgNGkBA
1kOzE67heHLnVX7MttMsR4lQdG8YOkO4B16gvQBjfra2jpA1LJ7+KaymogEOSYhe
x/vBFd0cAT21TCmYbFAHTqDztjLDo2grmddP3WiI1spBUEvH/vIm2y7dUZ+63tbU
vBgB3RJRClXZ4VXTviraacv4NJTw6SVK4P1BEnP5culalpJ2XnqXfrm9Bj52+Vhh
7ass3KUpv+8GETUmf92ZT5gVXy/BM55NQG2D6ih1zOaBzBaDoDY6Jcaio1I/A+JN
tGTykMWNmaf8QLe9jHvgoUFc/UEUAM+TIVkCwCzn34XH6eYWlUstNxPL9ru4KQu6
a2qDr9Iz0Z3WX63P7V1OY9J1e4Jq+zcTyr9w09oh10GtGO37MnbNZ4RrIKUCKc3V
Vmr39wFhj6WWOu8XWqg2KDtnvGQ/FNLbnaWvL+LFYJAiox7D0tle9RyxlBRxU01R
Z8Ilb31+eDSxedWVNKphBvQF4kY7cIu/pLcP1Cy/NW3oM+qDJTdY9sYY34GSsrVL
FJj3kquuOwY5Tm9hqOLbtw4t9ZskZTYBxWfXX61w2Nc7iKerlxK7nFBtSZnJUBk8
Uc28Nb8XCk2u9v4u4sZNOSu6tka6UKmTrddKyhgL4/toOadG30EUhHp6CO7RPPVl
isvMJslJhe41cwc7HSR0CoNYQG8asKnfIuCGkbhnfu+vYL9RwdnzLb86hNNFr31R
lcMqVBVDMs2Jvl/5leWEkHyaQyXs/62B3nYD8vWfkD1sPvLcQbm5Z3LsrC+0fojd
OPKygEhXk659t8PVBYkUJ0cRpdhn5gsRqSOg2/jCu/QGmRjRUf/7yVOJPIE8x7NM
GWwgCZ0TTcQf0J2Mb+1AaTQYlvBytVxMP8ag1XABnh1BzG1UuLAiK2mKGucDLrzd
eghijtE35e1YOsK/Ch4wfX4Q7vtXHlxn8OHzS0dMmPVrWRNlodauXkAOcbgaNYTo
fET9+wRdj4xlnwsDzW7APW5qMS0sWYfbyzPWYmUGc/crRVK4ISKCMx5aWG24GbO3
IuaeioLB3R3eAGEElfbqjkt8KoXKKW5I810/UR8bG99gBCGs7EW+j7qIbwa0X/Sz
qnG4QLON0r/ULgWoznW7p50SHs8Bw/0CPFzXJtL4k2Q+d8taA0nFf+d653bja6KW
HMYEhRhqH3COwk3tijCmz8RrK5sq7Iv+TqjrJiv02IIP5kBTc3pcaonobUUmw0JK
vYY6wKoBw2qgE2LXMOa+IwRAZvgtENNb5/cF7cph+eN7Q+6rXkHKt2f1nkGlGYmK
AWfZYMpH+8X0u7wlmW1w5jMzeJz38Y2Cp395dQF4hhRDhQu8Jwbe3cky5TukzSbg
a49BzS91QN7hvke1iym1zmZklOg1iqwkDo6SkNa1pN/niXR8qVaeMXyUKoOrfCIp
wbIwqhiPUl5hdKPci4DYOURJtQdEKboY1xQNUM2Uwrfb7kLn8ZuCF3Lb+HYZjQU+
Qfh0Jb6CtdaSQzUR41DhqaFlxItEgyTH69JIYljXN2hD3KpEm4eoXpAnaY8O/hBp
xqUh7g7/vW57ZAzudUv4XhPdv/LvS1UHrCvEzfaSHWSyAxUkcpsUr4FFlxPPtT6R
bp/mU2FQp/xINkeYWjOfpEEKoobQTCjuzvoT7kcGuMtjlUxlRYE2EN7Ygpq3ZBwv
PNBiy9N35KUbibmLgLQAPHuhgac7u/y7xLq5RqCc8hCgu4Wh3Hj3o9B0ZhPoeRJa
7f5GQto21Hoxqd0cb8JRWcvNn58D07o1pjHBTuuSgTaxpz8+ZWibCXPjzxb9eH65
fhUNRXHvBay+z6xn9K1xbdy9rsSr1VL8GBiw3cGGTZBcDSWUP1mqlfBfMGsn5qmK
h+80uE4urYStZ8Kn1fvM9aWpggfiNdRPKaUBWYzwjQCh7F4KMRGKC0nX/w9kuuz0
Cp0pPSexjmG7nUXgKqkvSFOxlmyTzjDmvJHLFHWPEe+TRjHyXTPMYDYLqn1c7/Gh
nmiE5mVjDppuieia05CqWiwJlP/OzRyX5f5W2hJ/bm7CF8AXdnEnH4+ovPaFt/zZ
8K6HHphuG2PjFrDAT4eNg4EG1dq5aE3RjCXL/5itzG4Q6U1R7OnGHlf2Y601J1wd
MrLNqlBFuic6ATe6heBKzdFi6Fz5isZZJmalzmTahZtVMvGszc3Sh7mxYGEyzQTL
2OsCWJzncYAezDaLkVNBRjcJj9TZ/NGwtHfBgHJdqGINDtY+0ltKFMdHzKpre6kt
EWf2nfCLktGO5s4hGLBwL7xm6FaUSEkC/lN59+UzEaCx34Vp++DQWvoj4w4Vlhz8
wGVmGswR07X11shsnvJIpv1jD4YUuSoSOjs76G5VBjQTFB8+5MlcV7PgP7WN3anl
1wGMwwCmAiKh2GstaBazG4S5+Z5s8CMtOqwlTyoTVpEcAxHtZjvMDqpRwCfvRrVV
DMxk/NF5irDKY5uvh/8bQ2YDooLEDRRSiDXpGlibEzCVOamJXWBPp9s565NaMEhE
vxLWsSz3wf0ubwsm7eaqQopkFH5FGmcnlGHKispdHu0JSc4Ty8RDI80Cr/zr2O/N
vb1Ovxe+vYUWdMcr/arynqlh9c0YxcUFl3H1xYG9VtNYEOBBTKdptkkz5MQRGPf2
Has5r9SMCDWud74Ul9dsz9apdBXZuVMtyrVd0nGYgQDpD7Ajk9iCkLL4pRPvRANA
zY1qUzb8FJvPXCn91I6y35C0DSgOIxZ8JUQ1zDBAA/JwBvJs7vtopMIUuQg/fC3h
ioM5VBTW/h+fIFDvoZK9vX7gnXv4vXQX2IxY22kV5qcI4Q170hPLECpUlNCDdG45
OPA1mH94FD59JAo+xcWH2VFSYQkxk2CmqMyGcNQUcF8jpcHv2Y5UaZ/RDV9NCYkw
dIaSQgSCDhhdwO3ohwRQYujVBPHc58D0ozSoovfT0qBCOzbOT6AoppqWzlxesx7r
UF9FfY448Ji+ikibJh6FyKJ9lSg6pDBDeSgmEMH682y1/ZWor7dd+jKFfpdT/y1e
+NQpmippHmhjZDKyP6HExMDnuZ7+HPV9Shn9JN8RCsiZAWBcxvZRP8nukF9KgVqb
h9rq3aJM5IPrS0efsjducf1oUqVkuEd6SnO3sRhu9YAbuYK95xuxeUT/BGrSg1hJ
nq5+w4w2ZeVCORpsNFcP9g0RnoBuxgU7UZlVIQNBHYIDArlMEF/aHlEmLaY94T0Z
tDh6set/zybZ0Z8YsehZC19HAIeEu5TUsUiBXdiYg7H6LnyYRoB7FLtNCPjkEURs
bF/0oi4lYeX9tjP2Gie3A//m3JY+fo4X74J0MYtF5oDI7/gxW0eyudj+AQRm8POQ
TmvVDGe4dlKekeaXixcVhhiN4/E9/0L9rSGMuCzueyleJf0eOogQNpMscTI4io9s
O4DKEmaQZOwmgWuE5nZszu6/YCcoWXJE16lt2fHv9FI5hHAa7FSUUxLlJO6UhhSr
GiuVi7ozgphPXZWlqQ+CQkU/jf/cLt0IkHTASGU2b53j3hsfx8e57B7TM1dE98dB
Dt6RTkCoUw7xJ8onbc0yD8kX9Jzpf8KnE2wKKhg2TorFfMZcYjYEyUtid3/dQbCA
cv20Gdpv03RrdIS4sRyPi3VIFvB2f8mCpZOdNlP3cd2VqTCxJmXcIl7yqE0e8Q2P
WJu/pjcZDxgjM0L4HZ/krkUUtkkYjj9NsCfzTcRbJVypQaJz1FVyLAhPMcIyh9SL
BHTOTYYx9Ud0/pjsM1/1SElVE35qeXoCN+16ckmXbr4cfPE10JVMG9GRwvkpocgL
7PhtC5NCwBeRrpuwu3SRnZ//7WLfL5PunLonhdcrViIdugN4mksGVuG8NdEq7jW5
GJ+FLT55tfAnaVs3Y4m1bFBDD7p3Pzt2ijUeMkBFXRoRHkM6PsulfevSyFyLBO7H
jOdLy6cmVhyWLL2R6FprFdsZeNZhc4JBO1EOnzi3hrghZ3OSyqhJR/rQTd05RSpb
6OmXbXdhjgvDRFNtO60TxSHZmCKy6qzdTAKM1KLE19UNJPGZe4fbqMLQdZ+Et1Dk
QmxgRAR8PQtLSjHHiZ3giF1c2CMq2TYBqERcT09THpR8PG6Aq4TGhdHhEUp0T/2J
Ad7Hq+F1+rPXA/VJzRHq3BZLtjxQuPK0cgYSxSqb/Z9qiqeeTE4wV76BOeQVSdLr
kG7vdwPkX0ACGBiw3Hbx+4LaXhIZUKTMOjWiDmSdbrw15num0Kci2B1EH1MZmoMx
FyHdwLR10Wy8ogu7dr0UlpfYHy93KGn9LZZ3MmxB/U2cSfaf5gpILa6Rg0Era0Ot
ceu2r/ZbKUFBsepa0LgauCXTCfX5FXdNcHjAMF4I4DTNdpU1slkjGPL2NM71vKNH
Fn+YCdEjaNO8H7CmNkXiv4BNE/rsnSovVJ4IwvhMhBYnqEcgkJK4XJ52SUOak+Eb
Lx+8nQnFqmJJH/KGfACoXbkR7FSDXJio4GdOROYRFL2//sWrrzNa8dTLx5z3ti1s
13PdinvAPBQaOjYq0F/d/Uf1ih0PGbb3lucM9dQ2GuULwVIy1+puv68jxzcKVc6n
3/NF4Y9HAiUXwhRu8Vq7pUBufCxU+mKBEX2xC58bAxbvLW2bJ6rUM/1/U9ZKKlr8
2X3rnzlASXE/5vL/VI695l8eFeUlljM6ep1zfFoT962b8AKHhiwACGWffG5UcZJC
cPAj5RGh23XBaWVz+gf4OvYicGKjWciy0NZjNN9LFgCML8RroU7v4BwAgA0pxsxi
x6VjiAyvLywA7l6NQBLdayHExhoaEr9bTZTB/TbRhkKRaE+mghtWugacBAEsZUTv
IzAnsmrpZcaKfAeF22PfnlIy1iCl3A0MivymKQtif1LJou9zpEUca0rpA9dqJ52O
FE7IXaNUxXYTwk/Abs8EjWnds5+Y167YgB2aPsZjLFfbw2ST/B1+7Ah2g290EpTv
N4f5iGyh07lmCYd47uXtRWUVDXILoGA/D/te1PniZTvxyGk9fTPaJYo/mcMFhqZF
eX18wqQ5j3mn9akT3q94RApwH/xixAX50j1UOScyJrlaJpF+wzg+4wwooTz/VpgS
BlC6yd1SAHWRy0D4nrzmw1vwSTEAopFaZQVr9Q2lK9njSpvD2QJFSAj9J0ldEhWR
ujsAVmrHQ98aHUBD0RVfIjj4YS+eh/oGZnDwuQyZWvaecVh9iORUP1gcn8kdmxU+
T5ZB9Gc5DMkEHPqDarE6oi+c23ckux/0v2ZqAf4dXhpeGhBEeapHeThdkhzUmTim
WbtVuDxnNpBanaIyRMZYwlKONRs92VgG1FBTkaka/Yqka1GQ42clGmAcG8gzAEf4
iJyrT8090iAU8KBWG6Nh1Vdtmc0+iZwlMXGVZXTjj8BMO8GdMIbz2/mayPQt3Tdk
PP18MQbw5cz6S3LyqlveEM6hzkvsVq02qGAP6EwYUr0O3GpxwfEzjyauDd6/nq2h
2i321YMt69BrCx6jebxJ50CJyR/k5VbiDfzs0Kk3po0mKyDakQ9D/uCrcTWrhYpP
tw+WVuoriYnh6ZKQ0jt8f1cmcDFZ9XyhDdxnCK6k4/a5yTL1ufb+kgF2Q9ypUUNq
fzGKD4qNCIVudvVziXW2gRCMo8gxjDfydT94PHBPpU1sSPoQ5FmRj5yBVyAC+cw+
ONLzAeCe7mJqqBfVNnoh9udXUYCindhEG7ll3B2+fLYTPBw8DzSWOWKmO8K4eIYu
IFIUzsBLxHoLb9761ZsBJPeKOO7SCuO1I+gbrREtjNhQ7ZNrAxMKWvUghTSgUa9l
RPrMvlu8xBkJ0mR+fuk4uv1qPyqcZQUsIhVY75qFvmAWQQXUCG3b8I55sRy5f2mj
2NRoOu8T20x4WQzMzqfuQP3nl22gbMF9I2fFCOLEBwAHhoqktd5tGPJCZO2JbHW/
17jBj7oufr00AOkaNLNpxBFunP9ej5LR3fvw1VqJBig0pD+MmOSWrWxCoHmhIN7j
xckQ2CVV7tuzayJr99fQuvP4LUZ1vK/ZhQjIv/1aJxvaiihuzlL5tr9nrexNq+ak
ya2slDV6klG+KmktJDZnaz62i1kWl59zwgkOkqEjCVyQhzschwHolhigPZQcLq3T
ya1sG40nOXmSeAC08PE0Lot7OChEAwWdBnGAqiWpv+MHa30BMgv+Jp50ckklVBfq
IfM80nrV5aNA9GERnl1bAhqnp0wEF+l9pGjo4s7WPAErpArdUALsHunU8xUbe/L+
wSH4Ulf7nQidKBuap7b5sakvwzpiN0njPbCB6e0wC717xTFtBSL2EQ+gdNqY3w/9
jvEVm3wV5la/VTjkA1lzXuNtDOfob1lHqLeytNu1SAb/E5s0OW5ovmIbmhZuhTjP
INZWFmxwH4MuZQgtLo0NNjLZuSPTDIQCvuqLplT6vRb4+TBYgoHldzrgVdqkMTp+
1SlrFsme/lnxKF3Rht++oOi+g45PfG0f6PqAOEp1zPvKKP5WZ/kNjIx7tSzWOp+m
axBRhmRMNGveLIatThQHFS7VhcRDDQ2vr09KXoqCd0mnJ5CMpKW6n0v6iS6dErWs
1ps08RYTo+3QEbfh6zW2I1fsD98Jgng3lmtnYdfkETepcpamcDrSLkuYn+cjl/gv
jKlMK+8IaW72sMb5GEDScDP5iDdgLEFd4gmG9pOoKBT4GdUEgcNNW2cHzKF83oju
En+6MseVaWrIuDOvbTK2b/hjltCjmobHDLbMhzdk8SUVzkFjnqlQpMlnoiIGUulr
ZxomSrGsaoksJN8P7t4LeWJe9Rt/VbTxDvs6utD/PBNzguezc1o6QaVODOe/2qdR
mn5nvM0dQ+R66XhgYzOLyy7z4HIGz7oeiXU0Cfk8lsPYRNgUXmisU3oO2L8xyxn9
HTAAwHUMJEduJhNACbB2W3NOB+xQx9KmflXH81tAykN3ZEiYGUUGOC56oQL8uQm8
IfaS/QZehuaWGiTdQ1PTYk9pzckQtyy8u3BGS8vAy7kKP7mMJSFJGsoB4wOBiXDz
tQzrkOCLB2QuXdZp3ahEkDCWL9kdMq0uunt74LhZ4z4Zm8zQSYM8ovxZQ78g0Bvc
22vhOpfgG69ZtUxR8B+FvSoFx4saHmfSYdoOqdZQMNlwT8VOKnb9Wj70npRyywvf
PVOdy5dmjo6MONh/NNf99thZuy+INTAR9RF0ZR/JIE4GCvFWkNQ88FUs/4+hM2p5
ndAKAk7hQGVko1AziLI245hLNGOuBMM8eyJnnOMiQ8aAatOH7Nf2SUZOEMQJLhY1
zROmu/M0ciFz6QfLV7NwkChMXr93VSEfo61qxTeKUWNmSNuisgy0ZblPGVJWHGmz
CKwbdv4dwbrmjTZgJ/A+SAUMicJIMYe/dhkfW3sjc4Rj/L3d2aSs3/LtAqmN3cCZ
DMKy7s7M8zPcVC7I8ojCAMHM+7eclBOuV8Rsf+33AHpxmoJXdLsCkiH/cNYaWxP5
8n/t0lVE4Bc12yF87JGySLzKGYc0RTYobhJ5bwJTy1QI/E9r+uPyhRQRJjxpi1D6
ZwNqDrpfy1E9IfXiIQMYUq5pizvqptyuDvXGfAUIxEBrrZzFfQLQ/zzwkWY4W8hk
Kqsx9tjQ7K74X0DDNH3l4z0nJQDNWtrg0MNwQLuQVfM6zx/SD47+UNbnTFEbZjvz
HjCAUY04TtEhNRIXN7rn+IwGo95kvIWUS4MRJWiKBMQ2lHig13kPw1uh+RqXU4Oc
3okGlSW3PaIrEznqAZio08+v6G/Q+E5DcpNpOUltJdn3AVL+OEiVSAkIzcFE9GW4
2hugURENQnmN+3LSVFqR9K9eJIw90G5/sWA8hONsgf45xRT7t7jhvRHaIr2QfhDk
rMUxQLmlTBgx8aGPhpbpN5c/vxs1vfcmNcCISS0BCKn0auzV5RxosiojH7n+kQhp
8nFxskTbrldQb53UEAAXTqzYhkbQGu66qjlepGwULFYLTqjtsB3Fc8fXQPmNK20I
/Jh0ltx+mrgHpeO6LLRwJsqvV+3vn7jQIogGv43p5lSWZDinU3Ay9SSA7QEW3/Qm
Z0M88UpovoAWy4NaJFOMXeIVNCQFf9wxl6XmJfOg0jQbFvz5wFoillXaOmKUqGKH
XXyldSVs+MaCX9KjBCWoZiIoQKk3bkYTbYy4vMBWKLkV1bztpGyXJpVJQ3Oi2/u4
2gGPGaT6yrSRBQArQW7ShkwpAxhhz9bfNn+fwMbOkEaI/gTmw4FjECZwlo9iY6B3
t+cwrBJtoOgOWFfbnrPSkUKIPoYAZxxtje+duhcSgGFzcSuKX9Yyl2bBIsvrZzid
ouLAUOyQyDF8XInvoVVHVQegjxm7FHVatkAQ42JfFkP2unyIhgyvlHU0dr+sd290
ov3pQLfJHJIvMro2ee/RaMLCgvCUxgG3YYMk2PaBLww4m2iV7ZdsGsSa3Z5We9l+
SnpKMO4j8EHnC8GEQ/osrswSd0pzKh7gCrWILc/jMnjpOpcDgnEaQhmr3DQT6SZW
Gv4iXkaOBV26SDDB5K41owdCT22QJ2JfDaVLHUqOhW+uQSvZiHJ4s1C32UO5yMjk
J9kDKvlSx0SCpk5Q0BpqQ4rl8xpPJyOi7piT9xXCS3T3owHx2+QdE7hxBply2Hzm
STq/erBZU1S/piqn96h3LhV4WTcU/5lztrgdiyM2dPkzNv4UN1wqBlqrbM1nReci
g+A89FvVPpNr0Qyag+JCcza+Do5WrncKnjUOr33hYgrEypznr/7F/b3kQb6hcPES
6+HH4T8Oej7O0g60RfuRy97/QjUwcFjLJUAa0iDM3TawfC83VFA4KfGA3iJp4BbC
kN6gEds6sruV35BPKf05F2NVLyk63J3qPci9+DwWiXFR7gXOu0uxWH4SC4VM1QdM
CsvrQcb/ktghE3BAH20C3emxv5jMd7SIv10sFBEsy/suUWp9K4gAbfn8jVh78v4m
+UmUFW2033NfS8T87LozgyUA5bMT4TrKmm7dHJSyQ/y43GjngwmNIJgzSiDe9paL
0Y3N1A6zwr6bCXVVIfHkjv0jLqj0LSEHT9TsfvAxhQ0pxKmemldFYFjgrddqddVb
WfHc2GB22xWgKfL3vArSDhF9E3wZB3EbkIoj5I97MzAUbEiGJ5Akri9ZQLYPll8x
Hu0b+qTxdQPMT9ycnL9olL3j0O97GHstAV7QYsSM9KqEMCpN4mFctUCib9qgFyY+
rKBHGvnxAxjFeYQ1XZe8FjI4U2dTNt/5CqoBr95m0m0ldlotItllud5friosb+AE
/MYjuf3/rVVAfS4QUefMMNoPhm7ou685qPA+uS9T0z9aaJFj4tyDrdkGUnKXJmci
vA3yx0ciMRhKT43o5HV4WkQ8pldxuO8dlKgWYvKT19KYTFB/OqVsI1VPaYUhzNLG
czPBLRDNXhq8yfB2BRqiY45vcYOJfyxzHlT8hgupRbeWWNoASJ7+viZeCKhjWlcr
8b9URFyB6ThDKWf1wHPrqd8JQvkR6EfFpw5fGxmQ2t2roawtLnQRzDdEj00LS9Hj
44tzoIz2+YSgM+I64gYkPCWN9uWke6gmVRfOB6wZpxxpFC1MBiDxq3Wzws3KUk/l
n7wa9HlO1zJXshm14DrvUw0IRdqIEzW4ipKfDWRsEtOtgiqmFF3sfgmRoaxdn97N
sS0RuOCmk/cjfCgW8d2eA0BELyQYlQZOaBj5mQTtaaNdmOhZogJb2XCWaW0Z4CBi
HOMQZShKLm9JB0qfl7gxbq4/SFEFhJ9/fJseR9zFsfaD2BN/og0lxmyc/pQWzdjw
ohoFnLBYRvTmXQDec/2ZoFY7bcr4/0KKusLjnXfUFr2lfYfIN4ekzL7FinyP59JY
axpz1kLQo9R8/Nhewnvf69hcFG4kVmh2IQv+jl3S7XVslgqLnjHuvIsZ5/gAqAu5
bV023cI/c7CZDEnjoxOrz5meL8QB3LphRkCi0aS/5D4WwIE2TPMOZJXTS09gzizi
xeLf97JlavDliikmBRPTcLsArMieOZI7Kwp/DDXpbk/ViPqAuuYHt/maBIbcqYa1
LWaSTwxFy3meO8nMhBxuxWP7v1G7yYsTwepnvJsqafJEJMk0qjrUMDOtvf1Z1rMC
kCUZlFIrlD2MRzjgphLwEVt8fzfcwgxo/k58I5Hsz/b+Ndmg3RmwyUrQnMQz2HZS
MS+Lu0a7aF0wfQoqjYbrEA9Pzkx/gcQ1Jc28AnWbcbZWzHdw8lRbA5wDXiO6bAHS
PoRzmTdTzIHEmhD+FkEwjnoonHuXEsRbFW8Hh+6CSyGP25zLA/oHY6Z07FBmIGfY
GF45SABD77LPVTzq+2lu6jtPoWDqLz49VAu5ke0bagmGUVmNvZ3eypEAbRSYXrOV
dNo3As1/pa5jxbgBA84nMkEx+C4Mb8N6Uh5akWtAWVNS633G3wiGGg0dx1b9wwUX
t7wpVxhBBHT6/japCMLqFqkZd2dtZHn6BNvUHaH1uJV4jfjc6ERYl0KgEpsRrXik
IGCTM8wCuNILVv5L+O3v4KeMfKqNL/a5MGGg2hDd6Du+EQ0aeT2U5a3LC08uwEI/
Y9V/JwM3wUkgKGZxkY62NwIOdKkED6KU5mnc8XIkPUwslqsITeACciuKqI43RkJr
45dcUOinM8Y3Z/aGCr7tnhwkr1VAIzCAZg62UCATszi/UslAT07b9bxMJxOXit1n
T+SwhF5911Cg7HE4Ztwzz40my8hAZBuW9mvcnMfz8FVambMO1jgEVbBKVDzFiBfa
3BsphwYae2u45qgee/dS/M4cnIgj5sUohea8xX7YxDmqP1biou31MhfItQPDO9Yf
eRW7tYv3hMhI5csyys5bbclZajtIkIpxN4Oy9R7DP6WONwI1qfjpVnfnkLr0axnn
HhXgadUhduyXg+w2QS5RH1B7OYzbEDtxi8MQRcLb4Vmbi7llwW6EkMqdQg6G9N9Y
Oo4vOZDtUqbQp86+uZTlZxLpBhhhjM0SAdfKc5RaJS6x7YeMEXvOk/1FvDJoIcwV
0A8LDbYhjcY5Q3r2aa27JCXao6ACf9yq2n/meIOANaPR5mFPVZB/slOSXPGV5j+w
dw+Erv1V33NHfk0pFxnDr4njGcoipRXzAndR7ysSuN15EWpY5oisDcPHEWso+//b
P0YLuE+jvN9B/NoAN0nCWIv3tdEZdZy4GBGLaxkQcr0Q7Svd9phu4MNmGod3nzT+
xNbIaMd3hA4m4sdMASxzMF0M0/NgLfTeuCBqOKZyc0E+kPwBdLAmDE5Cd1E8JuL/
watyCpC6C//NF3mCmc/NHKSpAOhmBoG/SRFV7/yix7OlFi2ZS2/VwGWhgkETo0+9
+1aQp6RPdXA7pNJCyiLq2Jh52CJ7OcrvQvTHRPLjZYxUJO1Kh0K/BBAx5GgqSZXu
3pxrtJZu5R+M5eEn3OG3hyW6DqhkFCmYBbOr4mHkrYuGWjBjPsj8hY9YqJYBAduj
ZC0HGkOE2yVZRfuiJ0EmDGaW9l+72xenO7rpqWdDhE5oGMLSHs+HIuadqKGQ2YuI
H9Ktk0ck9Qu92iAECnFD9MtUOrjXpIi2ubpVhlE8WzitqmD3+m7aGYD0zo01Blyj
MN78hM3rOXDkaMTi+XxNkV2/6b6L7Rlgh6tVbLcsE21fwV5NQM/RB1O8i4RCoRak
DNlYavYebc6WtUC3C2mDnuPefD/ofXsoOV5MSr8B3/94BjXyIdCLCNaplH3A1mYD
IJyNMVIoDH1+b5julFjt4fXvKtADyagpgAXf2N//pqMQmeSPuqdze9ASBbFiVHv9
WZqWMTIm4eYfziLOCuHZf6DvF3+FNGo6XUp0qPBM5nhYno+rM78gUoY3lpbcERuH
lVmYHOJuDtIfqWTs5hMUv7/eJRPeOxXWcWFrEUeEuHNWQf8WngLSc3C1pzzXYteL
nft0r0sJfgBaQqlzfT/KLf3HJicvJKUm2QQA1NGaLt7ZWFCZKQQOZ9x4BeuuHYOq
w0sYNdXvDB7LEdoDxcdUkkBUFZMMx9DA1k/jXzio8nMrwCu6lWgJED45Onvkgy5+
VSe3SWGrl77vkaK9LZTtA6aCxdn4c6QbFuTllvx94dmAsYofxyo9L5YA1QzpBhPF
LKOJdhlWr8/FbmU8ZzYYJio7JkOeooGt9D8FuJINWOc915YYgzzIwIXhm2g8U83J
sbjl1ERNq7cQ5IaZUnFqGN1LG4Z1zFBXxNU2QjZXH6spGw2bz7G0PF5Xpw2A+t+h
7x8bbjd4CXyM/2gNl/6bHZhkTyMgtnbC8+j3vJNc1mdv7Z2HUzR7NUNQOHSEQ7Dk
hNj8BtgddZTHGvYIOeb9zGLrRBjXbY8estXTDUuuM9fMwXMh5F4RxjFUWImSZ3HI
+L+qQvKvE27uTcg2s0IfLpquh8qn+ES6KETuZ0DTXIkXpqUESO22YxijErHKXamx
5b3fv8OMrnIQMttRYLTYd/Uu09TwUHDdYKnectDeRMGizhIK5QLGtnkOGvdHwXjb
EQxBpTV51rnUU4VYPSzPf6LLV0xl9CCo0PVfbWrsOaKni9ShPXGUzjAUf9fppx+W
QDX7W+flqgzPq/vjxFICGDx7HcIWQpdz0pQ5bhg9gaCtiHNhlUESFAqQEAdEkBrA
lLt4NS0E9yAQ6ks0/mwRkpbuYUWecwqJECAjLt2lGXK1otMUoLa78RirQEMhOUNr
vkpjEW/jQmBg+JauLFuqxBuFexk4+dK53rJIC2atlzBiWAvFjJnGZ1DokDWA+YRn
Lnu73Q+onW2p0MAj6e5uNed8xwcz2c/2nbEqOdarqCdULbRQFzKYq7f3q8NEsr0y
ODULyTBpmqVW+tExwcE2UnuR57Egd8cJfa27s6z7UHBG/mxR25orWknHG1xfFti3
pbge8wYJJq0sPvZvgq/XZ2Zi99WcVFQnGulSz3IAd8HQxIef7voKKWW86yuW3uJV
wnrz5jgKKxvoUhjTwlkQ+qP324mx+4ZBl0GAPdyAxTw9fjXt8Bl6b2iXPKd8b/df
S+pG5/qyHPPzGLXWnRFlzPRG9tcZrwnUjet0bvLX3UsQwDukl8qZaceR1uYZLe4J
h6sVRa9lr4xQ+Mf0JAD4t82vks5WCyI3m4fN5v9jHi4+FHT6th6y3Rdl99Vj1TBo
+ucQCJL1nkKRHceOJ5oy99PgpB+/3SodoUO5ZBpTufzX81RajqV0933drq+r4SzY
zHpUlpVGigNq/MI7nHm1IFNn8/FFQ5rYJIb1n9lwZh74fkystwfJXjdH59IoOolm
UWT0PPg6wPgKETQEKLgapr1qjAyoMRLRCGua2tTIinRBQ4ftHHDfD2WI0MK5M6VN
5mXHZeDku7UbuHgkJz02BwfwXYnV9/a6SMysspRbJ7GC9T4t5JUXXLBlIsByYtMp
lufh6CjK56DagIA1EjbsSasRrr7S5eRg+VWDe0l3RtOBpJ4aDJyISy0L8T4Cs0nm
+x4VPv3TPhCg2lClqX6yYgss6aqvX6C0XDD5AhAk1DAGowKrcxcEHuZP0J5xcmCi
wsQRRUZUzhMnZuPpXAfwzkC+PJ1QTB7A+X6v3yDznWf67On4wbZBMBiFhxiovuQf
PPrG1kl0ql84t1FJu9IRZldWYxKlnhrWC0ekJb1gR+p8gfwAf4dY2CdKwxzf1kae
Pd95eFThh/e2kHglDfqlQd2jVb0XQXTioBBETSPnIoM1Z4d65qyz+cdO4l/VfYNt
NYIZtPyaMKxeMqbqZM/DMU0F323ND5RYam22S9C8tyBwykMCy2/nM+P0Eb5F8212
Y60XzNUe9GGwsUdvAkWYblAn6M99S1JEdbODoUMDv18D2tNIWKCDTJWhvZHqBwiV
mBfPryLUsgbsx3SFhqZ+m+DNH2r8rHbk0TPdILpARQbcIu5+h4uric9PKfs/ogra
PNZY6YvijprD/zHHuWjC+SWi94ihTN/ewFxy2P5YDEjDUCm04XOuTJABUUAae0QZ
E6HnHxxNVY5Do7++SN0ICwmYmwdoa2Br85shQqFoQyZ0/9G6LnzvZJFT8sNvxMwO
hrrPQ/xd0idFdX57zihluu6/1W3yXsLNukAWFwVmH0IwsJNtz8Q6fMxTdnPqggnL
3yyfRTe76vDN29x4070ZScUA+kWch4/xgAYNzCyHAflkzRhcBqwSaY+XxKz64lcs
JUEQFswveiwN8w3iBuT+06lrlCVPXgxMvp4UsfbiAk9FSRqDW/iAb8zAwCQ2lYaH
oERCODocdKPub7yPuT0Y3KwV4wqPNO4YDvDqKp0Y/G1h0/I64+tJLa1CP+yxS8pQ
fKpSUPAXDwCqi/aXGQpurnnWlg+42Y+2HTMGX3EO7Xcr5S6FDerYbXYiKaaxpeAA
pJAutDQ2EI4Nl21tD8i170ebQzF45NLFzmCXKn+wM9iyk7SY4A6ZTLJEk3VQrpq+
BM4p8Zw1LNKYklWXjYufBA2vxEvRgGXIIAiH+CdXXOWGNlFgnwkypgObh2g9XQ/t
gJfzEMI7KzA14Wtz6ppYuIuI/pDRvSoKGQ/P+XuFbycb5FWbFvaeYrSN7FdKr1pD
m0oQwypHiVjmFPf6y4ux16AbLaf0SbEnyyQSqhUxTZ0mj6hzJ6KIRPc6FQQFfFfx
9mRjAkQ4CIerxVorUEH8X+qhVwsrpi1yvHt+QHSVWKy6CcUkQlJyjWexQvumsL4B
EAoxxzPjLV9cVrhr0nN0N3VvtQRl/dzoneQNtOB11Nd2jr1A6EidjJqvMnwK7Eoy
YsXppJUDmXSWcKIJGAs54R0yeNiFmp8B31VVIW+XgmZd6Z30JxvBbd4xKHkFORm2
0Bigc6ST2NVxjpBwC3DlG7ou1BK/J7y2m69sFlhb+m1xezbPByQV2nmxJeKILwaa
is35gSbsmw8TQ/PwhjeIBnNvzw1B0J829r5gPy2zh0l8xXgGn1wSxZ/IgWKo3Avm
FIermkM5oMO+7Jb80Q3lKjFu/YcxLcJ9ULOyfL8uUab6ZNzY4hEtLHRscUSY6veT
IswTMWyPnOcgy5Cqb4G+KLBkAMazqYlQrgtlyfSYnVSHoKkPIotswZSBOP38gUQG
GSSbP8LpApa67Oioa+7n1C0u6+lVgFJ/Rw44NVavMNuPg9Evlf0ICMvE6tWupVXm
HaRr6DA2axG4C9sJzpjLK88AyipE2fgg0zL0MZmClueHN+Wj3gBVFXaRGPadmwH7
vIry7ke5o397aBl8rB97+TkpRdjw5mlcmxQQ3XNNYTOTCOF9sRWAJLNcuU/olHI8
u5ptzBU1maws2mS6UQxwjkK313VxDW7DOowPqfP78NIJiZ4yYMUGlRLklYBvmJNl
WWUXRROcnmrYAluORBPr643VlgYrtZz12vQ//M1kHfMixxeC6W9CQGAeizjC1sbw
rYXnwZUA/h3JDAF+eGt2yz9FcYPt7sjGkkg+VxSZklXOixW7bsLwxdHwtmEgv06c
YGHmll2/vSA+i3xBHPY6+LtBQ3Zjb6VnNruS6qv3E/WKkOCW61YfzWkxiErs8RH0
6AbD6v1pr+NU6i/UDgXf/4M3eXmJXQhmJ3VUltBvjjdjZPAy9vEtju50kzoKw4+p
5nKeQcgmtIgbCvQ3PttiISFPLP5wlV8crbroR3SE/IIxv0A1sdPqPPT0Pg0E/SlC
PEJ4KvGGcQ82Y8FTr8YkulFe0zLDGLyxNdANJ8ro3G6THnsGUazFM3+VB9qmVwQb
osl+JOOBwbAq/iO7EySFP9Jj2PrXfuQj6n9NbSnOYMRQ2KffBsmUBh4CG3xTMYd2
nCj+76NtjedcMDYlfcpIOxAFOLPIiQySRept4AfpzA0N53bLZIaZzSB6dj1y9C2Y
J9nZcqtxcCmykxmNKAFfvN3KVWArGitWbnI91C1u4LC5ZjFjt17ADHlkEPuTYrFV
JOJ07jR777Tb9QyHRDMa1mhz8HqZF7Ys/xIBbkzjaLvm2alS1WYc2ZWVjLU/xceQ
NdC0DC+SErKieMLMcMQbEM5nRpFgFFSK8jqeYHe04VvvRxkDBwAlXFWzEpP/eGoM
J1Ho9E595CEyfqi4m9f8KS1fgvk06J2n1f6U8C0AYUGW+/5e1Px/jW+91hFmbTXo
WlwCVAY2d/bgZnggeg753UQ8mjKlOK2VdyTcSqW4UtkhOEAScdn+hPkk+nQMJKBo
h+YPS0kWTBLCseNu5p7J8A9N0vXwXICXlAF7/c+hLF57+iPSLSMED5gpd9cVst0c
Mea42gQ0+JcElqG8lYCjpM3v/42WSyLWJTlFitQ/QMw+kUaM4cFt/xOxLNsHGouY
DB0ZQWOpnzHY8WxmSqQnsvXP6rMMqN5XnS4DtRlhOUAGtsir/9DyDl4RD0zvRUJz
vqjO0+/FT91kGLgNw4KgX8Gq6/YhJJeCXjAqXAjQtMt9bpW3mh3xHfSUxWll04cH
s+sCgqaTQScD3F7Ggi2vLTaLrDV4QZRRS6OW5kp+UQlNc0gsdfmelWdXV+VcyvP7
8vRm3Y/ctgFck1lL4JwliC9Ejhh1BvbF8zx6Zz5Dklo6uPtnY6Cyz0KaKydMlJQy
qEy1ptZ0ht+sgCEijwEu03Z3C35BppVsRgnRb3si4XEug7B8z4VDkPfLSNHvCcYg
m8UThmx7sDnmsrELQSj1+KI5DU6Cbc3C56XcqLjqraHGMS9up9OZcXKrby+SmxZx
98cw21Q/LVarea07zrMfVJFafcvd7kfmZjjp9BBwedbv7k2O1Rpd3BELtYf438Ek
HdVcU9rHsdE4ZKSKbXXvu6DcZnJV+XZcD6bgwc8XIIgAid7wRwfrF5KVzmR9oNex
BVdtZtJZbnt35/Ls3imLBBb52+zA/S8ff2Wy2p1LEu+gb0GdvDHlgUHFnSKldVhT
xaRRij7T+BGeczdCJheRcDY+xltwiLir7NOxbIhXEnrZgpK7nJegtU8kOk+50+Jm
7gyxo8mYrP+Kisj7EyhuXExWtkbMipmSYWQY95S7PFLSqHPa27vKwtVAW0IMxuNL
OuNcLj864R4hlOhz/DDrEKq7nc2yaCdILD9Ckvn5PFSAxtGpBe7ILTrsoVpQHhEL
wp5FjBTstai+23j9aKr/hviMZfJm+9dMRquXi8KN8ELBzK1wi6DenpAG2ulAhoF9
2hYD3J78RI/bxCYpE+4ekO13hyA7oQ6xQyBD3RciFbrWDFCj8ic46hbNz1ojbVee
2HltsrJ6M9s631XJGn8igm663dgZV1ddf6Ax72BMMD0sjKgf14RgHBjQT5YRKgUn
Qqn9+Nnq1+26L9zv9+1Sl7qzS7x2pvD+cjGw3e/b7IPrWyMucOnHVkPBtotL3WgU
D9HDdBqdPpFFJJyw2ZgWJWMPmV0/T8Q/PamrBCIZoLcZJSDshCqJ9eCGqIWiX5lw
GLKK0+c+lXXnFHfnumMsuWYsk+/R57SeV5+oyRbNlUtH67/JzasWE+5L1UdFm6j9
gKVg/520omJrn53GYgWfawh6JlW4FVRpUk0tMrnNI5N5Nh+CPJQDAb6LcXwbQLUc
/3/go5I9FpHzYtbuCONLRUE/2vQPhygtWLRyhtJ+4IBK1PCS+8z66t/KhTxEFHyk
EVZnf1Uno9Fd1SwMpLLtaN79xnuQEOLcUCfm88NGU+jJPrhrkyh7ccNLz7d3Vidd
lardKEQvz4X7mN3FhNlIyNhIC1WWilt+En19E/A41M/a/N3Nts9i5CRnEPIE+qOw
hRgbXrUTNlLqE1a/d+Ps7UQNevQ1ZkwUhADFcIk4Dwvgqxv5pzQ7ykKboDiYZCq5
IwKqgpDqQ1I98wSlwW//G8VOm3jEzNCEojL58z82J52sV9yycbGg9hMW1y07IFkw
pP2ywbKUli9Vl/gFCO2vol6PP5gjcXccjzJe/20E7BJETdCtma4gp/U1mZNLuLcu
gWgn9bF0qD46E7g74wOA6WP7pqp8ITHzZaXDChyL1MsYnybpd5A/2+eBUcjiKaoM
tmSIzDJiYlkM/Ctj7uObraRaar9xSpGkVM+2+xm0Z++2qXuTiAEPE1pyCowfnBjj
VWTQpjHudYMrZXG3ZK3mkAIo9dCAAG9LA+ED4tRakJzKsptUeol75SVmBAq3MZ5D
qfGNLdLGRKodLJZsCdM7VLQV6Scx2seSLi1zth1NiEBg21HB2j8RZyidA8ZKeV2Z
aY2RbDaYwDXEN5y4pcN1PSUPWZbZUvDVNDbpSnEnxC9TGz9+Vch9AjY668gyNr10
RPgQmtd5UKvhbiTJ5LcH4aM4q04TH+ASIVicfjgCg68iKU+YornwQcr6IXzhNgfi
GnnTJn4ip1IjvT/5oEAXER9Mn8gRukw65Q0gcUOTJNvnpffPqYBysTAhhwGTSZr/
JD2feC9x5AVGVxTqjmPWRbRd6kI1OUqMEf5hirvPv/dnQrpciRUE/EehBkPwCZqz
0dnAVc9jJG1yjWoBq2x4tJ7DEpe6FtX+tSfx+U2XhhFK6fdaITVhz3iKJzsNoI1g
RB9JqUsicOewjRx9a+W9LabxNKsB/CluEz69xsKfiborS6Lz9YXmjOY8rqqwiaQB
UORPP7vTF+HBq5NqElw6VSlHiwjqEgfeoReFI80NNyZ6uTR4e1miItR2UjAZt8H2
BQCggI/mni57FUBZnhIXEckS3kFLcVrGebXWdfUMFghoQA9RMH/NvRzSzbHM+JAD
aL9oJIGWYX72GpRMM4kIncpBA6L1oCaJ/MDvjZhVAz6I5PI7CoEluvhKuHSc+tSK
u6/vBsQ4Y0KHQooq+eJHzHZ3gPn6jVjcPH4MyAEDH3axKtKyn7+3ksBtxBBUktt+
wvTvgmpPs4bfJn0ipV4JojwX8Dx11q1WXVinuVKMaM9V9NP91BHZUkSLg3xLju8v
j4G0Ai+Ri+eXkTymgj1XLjsdu6lb56+aM5eN5h8anNQWXCfhNfg9AKbeAkcBkpHL
3j8cJ7NRa57CSk17SL+B/9F1S9xE0PnBGiGWPCVwTMpgr9XomQoXAu8ASeeVzK6U
uBkB/uiXMSGSd7wo3q4sZAodFZ+qeHa02BnLmYyNdapjgprWDS7O2r5iENc3KOQK
6hgK0K0K53EqDUaKobmtIatuT3xJI7yh+N/O/yq0aiDqfAzflkoyibjpvTFr1ysp
ewJGKWmYgAYPrU93SujyHFCqHs/dx4FNeed7hutY0LleD4B5B46I6a1MXOZ+UDMD
wY1RmK40QjndAGZQJsRLGtpW7yNwP5MnxGXMWCMOqBc7+Jbxr78cRCBrHD0VakCZ
8Sy+YMteFC4287pQ08PbKqB0RmWLx15eSHEsOGhiSSjPNrH866ruf+Lhkz7KdS4h
raEIEgTf47QIQURGBztL3/St6wqAp58TEExVIDQVJE9Ufrfa1qBIuAg7qY1nQYTY
qmo5GhvefKBIGCZR1F5zWU/y2PwDF0Gx0eYfh+BYIHiExaeWfd2Z9+sFjWEUN2jF
Z/Zux15pABtL+0pzRqgi6qeYLQek8CRucZIr4xY7Pao3ws3W1nVd0oTPzO00lmJO
79Wl8vjY9utza36ZvvM9JuCcWNvaHMf3HUg9GUzoIh+znpdmG8Ez3KcQbrRTKGXz
W12pgXsMsTcYEoKV7/ed0h0RQp9DP2Cz+F9ycr2iFa2YX8+BhnVpKEC9INFEMcG9
mMFeeurFKLJ6sK8MRG1PSIHtPpW3BvcuG9h52zJAQxmNLdAXYX+wTPQ0j92NzCkL
7gnVL8GVRVoEYQKw2OaIywiNmvaTUfGR572ZUfWeIJOSwUN1uICqAQQ24m2UOUS/
Uqzw5gAe/z/uMAsHMfldO8mLR/ys00hLq7wz0NH4+zuZnzGXB6L/saB6Rzg6gDz1
yqKJT4NHCAKSY25p2YWtlnkKzObpiR23V3smlkzgGV1wD/4aDDzkAgn52kn39Q2v
S4liJW/zznERys1isbh8kVRnIbKn75p9bRBL80GFq6kMHEdemB0mU6SNRhfaWaAe
EQ1KCndGYpjCT9BDvjYrRLUKC65wZG7c6qdoupCSZCM/fcFbWgoVF3NXzHu+Aa9c
J3B4Tri09dpLE4+j882wWcK9MmJK9sApVsfgN/rjYS9lrmhYErqNE5bcvsyoJkm3
iXjN5fp9T6xdDdupz+te3DiSFtbuFBrnPlk8jY0MRlC6YBCeteix8phDZUMHMdKu
Sn0pgtGnahvAJtfeg1Hk4pAFiduMYSCT1DzUyzbeCtNXryiM9gRXzXAHiGX2ohXB
MNJoLKXdqvx3DyK6D1G0bhGhmSmAC42e6SmrJLCDr4OJZByy0XrRGUJWRWZwZcTr
NmND6a+eV5keEP81n1pIw+N4/dBllhYrtsh6lxipIM3IsJjuP19a/AScIUYRX5l9
YXSkxAESXZ9p2KXzYeaIYVh7TogobB5dSGV6TPG0eRLHIcTgP313CvMuvFqLy2yI
miWoCqnFN2uesEi5wkbvAioWI6QKOVfnCX45E/laiOPAeJ17mIwns2RbEiEFrQPi
pI/ivZtGv3qA12y5Q0Zo2osF5M/lidyOYK+SI5Qs6uORnemzBwXZBjA/i9R5keLI
aBWWf2F2OnMwY8Ou6KK0CTxTCE1P8BUnihIS9clUT+6yPcXhyRtX8fWEpXiOH1Qs
tarny6lQuq4FrR2aY2KdCWsmW4HoHbMT2P5WOpTPfiTGQj/8UTr5OdclZbYuDGy+
pqETsy5vqDjjmCZeRa6yl9pVlzSd8qqy0gBGQJgd0MMVRZvr1JnkVJ4cGsXFIJtO
bksoLuNjC6vNnPQ0AUSCZv/rXWAfBjYmPcSj85lutQvBVnViX3Nav5VffCqJBVkc
MUm6mztC0WLo463ptKS2KdB/WXrYnIUu49WXzq/XN5vm9BffSyKXSdjlIvRF5hkR
t6k8+/eUOQFO0NoXE8yiB5vaHEy8hyVslQ3QRYTOkaGHN/N9GFeRmBNdYvw51LVr
GGST6R+cxgnco7jBov+eSEFFWfR78rW1Lf4w+qb3fGSAa+D5lRN0D2I1lgZMfzFi
O3BoC35DTpwGCVLPv/hByDzxHFmm02ROatPWVIulVRShyXbf/sq+vyfw8MgkmgR0
sVNCA/wiQC9jIPQPoQb5zWF5ebHWIpjwcv3p4WbMDQRXOQDtieu8wXh8B09oVh1Z
1v1CMfb6eDnMHINOw9cPdiPXlOkwLpU8YB5fWw5NyB9cVkADfcwfLdDCu+lvHOYW
+ntPF0LQ+Qa+AifJMqv7a+i/4wapn0p+syklMyfyqqjiSgd0HqSrBlKGwGN99UN0
DeUGzMgMNIsWCqznteTvexJttvL9d2FKZRjS8bFSrcOhwpgDdFi/bpgYm5bObDAH
GjT1aecjoVU60duXOL8FwZBMf/ZMj/pq46uVqlRHAypoz4r/w8f9sQybUAeNOjTQ
yJhS48Gp3ZiH6WnxDDEVOUqL0Ly76+AQ/Ggbsq0YCL3JHT2QAFQj6Z4zcGrmSkNB
rmkClWDac1GtEXl6NKglbJqhP2AKv+eW7dNdaLOxkbvv7A6sqniHRL3jHD8oEDz0
fc+X01kDx5rfTmV0tyCW23W4fGnlN1LM5pCcKdtXAvouJGD66MPFIxgGm5Qh78JZ
Ke4IJ2vLtd8JDidhPGbb9o7NXq2IdG5M5TeeVgUTQBppwLutvIJ29qy9sXntkSVC
YA/E3evAsumhEqUjgsMZkfvIT/kSb40aYD3wDLY8t3h6j9VPZj4jxmaikvUI0FZZ
GlF1nQtqLS5DGMiLsFN9TskPI0KqgAlbTJqoDXM+utO1G7RG06Hi/jVbjMM8vOFZ
o7AhpWyfKu9QB07PrmcY+MGizKyCJEsmjm5kzb9Mt5J5Jn7NyZSMmk334cleOD9u
EMel84zbVuNgPdspsCbgp7Q9f64RckRamZIbJ7EDczwvg05RPj5ZIBvBCZfQ4DKm
l4oBS1w9JNWqcl83d8DSs4qFpcbdXRvDhGR5Z+RZuQ1jXR153ItQfq/sRKs2ry7H
BSRop9AeAQfbBZeSIZKwa4t+v0QLYEzhjlF+q02aEDRu24tXr5Oo+KzzGl/mEMjR
yo6uRcfcV1kGtINbZgBD8AXglpONHLv+JaodFCMfSH2RYQ730Vge3+tzaxT+WWG4
miJ7PYWHKofUOqHvPqyVqnfo8KPy31r8/Got9DBzohJ9cdTMdplqEZw9K0uN8M+o
9cdKvcrVWO2Hry9s3XRFUj+xLRcyocQXy0fRBNCymllrLaQOnt8ux+RVU5HbQMdY
JS1MGm4aWxmggU0wd0tFRwsJioDUtPTOXpDmpK8H/ncrlT7qpiLsw99A/FJE6Gx4
DO/ELdzfSEURyJVcqXYTJenv8yaKEfVyMn6rHXuZW9O2vD/9nALLlPlYaSAOk6Y7
P6ZpDxWjmuBwS4sgBdY9tBd1+BtgeHO+hrPtkPWIAdAHMwuoW57wY7o8oisErpoK
hmcyftzwqrXqYtlXieKruuIEmopmyPOAkJKUkaDoxUC3iGCHyzeRDuobWQ07uZ8q
qC87qGSz6142TdYvvIfLlAk95nblxO/YJvSa5lraATBtc6dpLQCzRhj9h2vXn698
tM8HnEbBgBpehUcX7eGh1lbtnMM6LEyZtP5WXl3xTfpRPx84LD4i32JvUHezscLF
2J7UtUSETHDy96HXlKkyhZD1S9UxiWcJfVhByJzo4Mu7tc+fyHsDNXVswmXw8RKS
hEjHvsLQPr/IiBG+WoJpPtG2tcw403J/LTR4fCeAFFBsXTgoV9Jq69edmRZdfiTQ
zfQbmVBi1ff99WeXhlzLJ/rHJCgbeJmd4tLzWLN3P/My4f1DMpffBD4PyflNXoEe
JAdFL1lSCwMaGrA+RNm19yMbo7jr83qAMjHCtgs+8aoDM8+y4s67LX5TifDORhOy
bKy2mYbL1FMxX/p1+/eUgxxBGGkjYPewMU1IFi34A61nCYsR6jQxhvju6exPg1qc
Bzb9uWms59RMGLAdFxkigH0w/CGLLS01VCT6NW9/73MCMxgNIs/8sOXiEB55izxa
pj1//Rgrq4ahsOQsHZVSbM2N3Mc7oGutgEAVYlJDfOSMsOqbQG6NmktUvKEcoyYJ
W+I0rAr5F4YAECrk6xAQ7ye58ZHVCiV3QNMGbKJ75bBwKYmPI6TeBxh82YOQmaq+
0EvoGae94zMG4U/D4cn3+Ln9ud99VqolTZ9V+Wgo/COxNmqEx1nD03Run2Qazdvm
j24+/kSjzZj/inTfIItAYWsARwie5IdKjE3uhVfys0Tqo/CEVFFF4hyl47uVE/2l
KlfIZ0/aB9/3f9On6CV+TnCWaL6KEVxp60ad0/s4GW0wRJyAyG5CVZgJ4auHHv/O
UsWBfYEq53TpNPcDZ1l8sPFkvDQ9R88PwDRNGb+ONQU0r+pTuWWEJS29lYw4m+xt
v8OxkuLFfi0hs4ZWpeA/WJKawlviCSn+h1g5j40SNjpN8TtYO+4zY7KILUhwEiNT
FBMcb0jO6rDWc8Mwpg+oDPZzODumGH2yw5nFIH01e3OYC15gXnT/0kBVLNQlmdE6
fFIA4k+tnp0yKQ6k+6xXvHc+RU0Ur8TdHUYgrQzQhzbhbEXCPA0MObD8UsgzuyeI
QA4xTeL3uPaPQvsy+28UeelJ78cM1a6XRVu5eZvoV6Ih9fH0V8TyQtZO5lFo17EM
u5uuOqeyC/yGAeB/F6NWgLfKl2XiITbPYmY8q0ZVVreIuba4c9+GSHFSnZCu0Duu
yFptKhGjQKQFxaWSJ5oF9V9j0bQ9AJbuvIRDTCcijbd2n2vt0Dv9LyCvcFDG9Jkn
EkVWrCaLSC0bn2BzLfwoWNPeR7a/8cv33ZAiOHvKOtt8EGKtZMiOHraC6dCco3lr
7cg/a3kdJri/g4MQ/FQO4SQjuMVOvvnXW0D+6WBUiVEKpO5846h4tsQrcf3AYVth
lOTQu8+jVk9caMbINw75b8O94iS6ObjFOcevjQRqOcoMQk66QllCVCOXe9gyRh7M
xOq0nA81Vauh2OG/yghbdbJ0bTRatPfMAU/f+4kEmlMyt2ze3v0dFheX16HoMCOT
8iwJHPT3cyFyaFwVPm2KQJjop4yF3eORARAPd4vqSaplJ7c3E0CBy3S/yfT2bd4z
lH4i4M61d2Uhq7to0o5ams8zkL02wuYldd5+0jqqa2H9KEk/xttoafI3OcsUeAxQ
6rcVbybqfAUu0aHtWJJI60L9DMr5v151ZSiDVBZQsfj/Z2Q3zEfl3aKRcm0WPybX
uhuySYdlBY1F1GbPRultlzD9Yro95RmQW48SnlozpzgMBCapUuIkNqAMfLRzt4UE
IaOoH6P/Hj3jz4yE004qw4WsSivET0q/bLeFzIEsn+pLDJk4LbKfj1bqLZ4XNCoP
iG0M/fB6W2HEluQh1Dq8UOoR0S9SlSv+J5su5O8DKi5vUxj/yb0OpNnwg3wamAR4
1EJS1g+9jpgfjNY1WKzIiV69eQlMGKnz6gBOZmBNbEzLo4ODdABV5OvpGcAY1f4w
yMTGnFC76MRL6TQ09hftCVgwR1cL1EpDyOBHyZhMxWiwgIoQkO4d2aCIM3SN7IcY
Kt0iWbu60ZqM7b14IPUj5pC72oHyqTuUB8ai30A5iJGr4rugCnOqPzdiIuU3RrTP
a89/wqRQ2GBjIWR8UPWk0Prfipta1NxgFh+P6JHv8/edAGD6R9yOp4Y9tRUquR1H
+bYwoRBfCnwxM6qy2IMg8EaJdNiScyjSK8FxMcDG/P5husu/NqLb7+HCbq+V0MQ+
ea7xZ5H9ugwim+d3cWTc3++j9JoMQazJKp9+jB0NiI6w6ZpGPH6DD80e9Wwl9D/i
3olWj2bG2+1fSz11STWu2nJukfuFOTkDqLBNJAQdHequxt8++3KbpIbmKdlXgpAu
k8gtYXje/z2r4g/2aklsFGX3fGo8Z0rK53GTPk0qe2ZvO1OUU78q6SHuuX8agFeK
1b6mGqpsZQR+lmKPaKcLWG24C/4/n+FsCiHePzSIuAnb0/L07AVpTQtt6voX5VTn
hKH45Tzca2qVB0Vcc8/LRg9EqleIG+7dprmq3QiwoSw5uNwKSd5RFqUQ2Q4dWS8d
bpXXoult0xU2TfBqYiJB14Ya0CjslLrWR6qPlb2bO3Jy3OigQLR4A/x9kVFPlWf/
9jeykie2UbM4HqY7rtslwXzpWMeghUfuD3p+UOSbOnq0hDkOHO8mryeb6SmdMLT5
U3xoj2BN0jLc3C4qNq585U7NyQ12fDiFq/ppMfVu61NjvjqYFCKsJAPR4/tWbHl6
TekXjcjaN868XYngFfiRD8XgFu1za5w9YkzYlM7dHpVK3D+1+4LNDCWk8s0oEhDK
xkhZNt2GJZEQNnO641DFOvdBZUHbRptGk9z5vJbBMZJq9E8L3eWjb+jZY9AWNBPE
mtWMNDR5ZWwUpwPZ/ElcVFQwPMvHv3Rh7YPzU6i1aR9yERy8S5T/sJdARWVKtkh7
/bpsOojvGe8HXsJHZV8FCpxsfmJ/0jHHYfoevu+p2Vu3UPxSNV7GhMzO6km5lbsM
L32OHLWBsk4MRQgjcam85QtaPRfnJpoel/pkWJkwPHHEDBEfbMGVIX2SsuF0cyEX
D4rYDD5HbHZcpGgVOU2EtxTGaYG4stnkfdZMnmr31PH9UuA5xFkMgsu4N3CAF5r+
GHgB2fu5sJUQxYl9lpmgKiALuVnNhCJjO3XNZRxQlvFumFGUJIex7mY7dsoOQhpi
olQJVq7qcZ/aCs+7ypPFcM7VdiYSgT4ExgHtW79uqsjhXXaoYlJtJ+gNprkVHFjX
2BMc4icN0xtd7cib4hYutjBsPVxiNWywF22V4vlomOpKpaXcs9OnqGVug4ydxanj
DYsM+XPr1xVHMyDznmJNx+9Pi3sRfAcLUU9u8Scz4plMG/UdDtMzffPAZDDqPzf1
7Ef6x4QzeXq+oPVzsNajeL95jx3LTr5am9ZHtPbQcw5nfg4ifuoVH+1nA8oOo6M7
gXuR4G/j9C+oeLLly8ru+hEqL7/+NBFECRR2dFpTG6XAIuWBVnEgUyz0M4E3vTGv
UOfDCcNMkP7eMj6pSdnYQk70w3kHr0hn6pomaUhSF8n6FUsDFNj1Cr1GGd6PBJVE
nwPU3yl63EB5hhpQ2ksfLVj+IeogN73yAsqDRyhGxfMmDg78uzCK6l8YHTL8LcVZ
j9L0fKMCg49H4l//6+p+rD7o58D6bJbzVT0rR8eXznrm2B6SrZ395BWCrNDJihWH
oTkHdaCpIrjeOq2bj1lie/qcvygm4DQxR2QscbV+cKRDszB3vIsBLZBqi/poac/t
dPol9dBNThGnRily0jwm4P5yOtdpqsutTrPF7qPbWi2M492aQL3nImb2+L2K/tpN
UkmyyeSc4EjDwf3l9cqWDbEMqiF4sUJyB325M9ZqUDUIA14Po85ROBAD2nvt6G/4
Xf4nTXKIqGFeVakihoRjDcdDhu2PKUHUgrC0JWdPD6nOSQchCc/97YmuocD55W+X
1BM/lvIwWL+WIz5r5dSBtulEv26WXexdL3G463BBm7y4Lxv0WcLTtln/OF19DA9r
Ud86LlK6LuVNCnThPEJ4s/Km3GTVNZBVtdyGz1y63UO6At50D/VEbgcJKzyzryPy
B/IbqUDe1an5u0u3bf06LcPAuhOHVqXW9/bgTkwZgdvTBNfVjIpNnOkUR/SVBNUe
a3Ep8Cck2hiI0qVf5UR8ais6C6SjVrzhcNsoMYf9iXbgmHKnLcysN5xiGhR06jme
RyTHMIYSAojSziBuNM1ScVmBVKepm73050uh0KScLx1fegqw6uw6yYlmkG30OVFc
ITYoMHdZ5Rog3HcsJP77wNXLy0xO8Yo3IcgvCTArqtFKvMy37gUKjMXMjz0VxoYK
97AT0YcYt6PoXzE7aL5A3ulovtVh92oUbcvBS77mwF1eUIXo8Kr5GQZLphoxp4BH
fuCHu4bXakBQi/wiXIEXKLpi3zs0qfJCUvOCx59R9v09xo/tO7lQVBQ7Rk/Vn75H
W70cPc+1fXi33BsmnzM7btrngI6BREx/4cXN7+Me2cjXpjicETPTpaPYES1WAH1D
dHr8QI0SfQZYuEIVe1C8ZSFoIQkgYC4nuAxrlHvl178Qu0kCN8KUuu2qKJNuG12f
1FWBYFuEjj9wkvuaJRfvGx8hdogXLsgClk/Cgq7USS6Zpv60RtL/xOAONdh83eoK
5qacluBEAdc6VY/VVNq0RZoNPZYSlj5a9RzDe/glReUcSXqJ1R6LGBySr8YYoLSP
aXudyK1GyC+ClN2AptUV/rcKpc/DnM45yqUwQT+TbFfKg6s2xiQZtGVNkLfdjdU/
okSoarnMErQSJGJRPTLTcw4G8V2u16pxTUDV4BWUGqYTcQKlTFX3KYz/k3AFseAG
REVo2mIVXzMmjRzi0xE2hgu7tTKim5NyK0qq/uhHqYvri1bCZiasoga3vZTRxXdn
SYk9+3Xdg3yiL+md9hvWNPhZrkinVqE8wZJenQkvnJsfma2RQj0LvlHimfz4kGQq
ve7wSlxOHBtnO5JvzkI0yI1C02hOQFJL5SdFKO4rji7RGXKwrt1jJy5K2W8E74K2
Y5IOCeAINttHCyptx1ysxvhrHFjHhiAORvVJ+azXxDYYHM73y7mVfkkOuAS4vyJM
VyQ9QiD+bsQervL8WJaM1CthFglS+UO+cmb5XxQI+Scx2SUoK7st/FvYLUIyxXYN
CbumAnWD4xxK+FTtkoaY6RYS4JGuZSDoax6QjBpsObbOba3E/fsYc9r8bCPJwAnP
nVCFn9jMWW0VirT/AuwCaq2YXDR+hKEOBNO7Qm78Q+q/0xZmL4psRkYXCpNyHfjJ
hDzPJGoA2FPn1IlvNN1rbwy5eG/iXEUc9kolV28pIECXtsai2cPEAZ07uvIqDaLe
GUzUaJSDp0PNnIflxQceXcREVC1O3ervBgF7sqmg/X85+0fTy/ZF8Q4cTXIE4xS/
H07YAiZcu/qXYbuQHcFgCe8sRQ1vy4304ssMwc6ERCiTBpfk1ZSj0S6NjMvX8MeP
dbgnJAQOoHUq50XXOMcN6mMp35bZQaAfXv0hBNczEchPmuuEMjEP9xdIURoruaBA
/A1PmR7OpmnUp7ygjxrNYGYukES5YbOE3oYXi5RqYyZfj3bzTL+MgBZV/3Pc6AtE
Hhf8o7bqkc201nehy2DCSWqd7/BDGTeUgtwUmORE/wJVa83JjfyvundgPGOrJwdM
+2LwiIPR/3Vvq9OQZ6rM+KB21UV0ih2Y0Njs8v97e+W1BkHgngthtq4SGy3srr1O
/DYT5OYtbo99upqG4bUhCsY6RIM+DWSK/5BHk7bXMkTDeKaEk3QNhSqI/TrsHQ1C
q/1eltK9SKSA3t1b7k1z90spq5jPc0qJ4b9GAd9vKxeX9F4kNxcqYl78gA27MAUE
bsUskA6rJ5/1F3OZk2AA2EeZ+2aKR2SXuf00XEz95nY+Aqf5EjK+AuZKZoYTHXh5
Y63TB1eEoMX4h6yf46OubzdeCo7gH60LMRgZPnnWA/+dw21nrvYjYbyEvK0lmyRh
Jh+bzqgMHphWM0KRiiZIsgFOVzS1vnJ6SccgjVQYnWa1kaLmVBU4T2Gaox4OBlmA
z0CrdrSSq14gZoFDSY1spHMUF6UROyTsCTPJACyIwQJvNUi+9AKijAm6wNAvzVXu
MohNyBt3RLX+ikCTLlcX5OL2HclVzHy+GYOxaCACt9Wchd3GubFtP4EeatGsmNn3
92bWcbpelJ8iaAjb91mv6WK8gelxwcDT4M3qwjwGd8ZvASi0t4TefmRymSANR+L4
uHE5O5Jkmq+4FFANd0KRKBEYzNobF04EC9B8VI3F8UYsABtykW23GIEGEfhCfB3S
3C271T4S+yzQMZwfysOPqjOOx1N2iaHfmvyQfhPQjXUBQNWR7AakvXV0gJbKmuXa
8s+dSjjh9cx8HAQ9LJ+YrYm2aAFkJgBtFc7niCNfvpHVxsbLDD9o16k4t+6tVK3m
hKs4TqTir1V6uzzMoG/SLyeZk4DayTR+nPsoX5ib0qcOxOiJyrBpN8rEut6+SRKa
6T8X9vqjycmrx47C9G/ob5y0le4LGCp7s0/feXRS5gRG/lJIVAxnsgkWrBrfF/64
kNe/tAgVWfNZnGbl1fKWtBTqCwKNrBswi4DSEEBzjcxdh+8sT0DWp1RPkND+zQdp
0dtPD+Kh1n8FrWAYmYhkKYdxHAyx1HKRD/UzqEYYwE80+V8JkBXBt5wSVQNj8qfX
8N+mdcYS9t4gdkLmzE03+oISRAqVItTbUpWshi+1HMEuyp4J0CDL6MvvTbjkyG8i
hoICs5Yq8isW0e3+snG6PYlvw1rjRADrTH+azkDEPypiw9qlDyPFRjClCCwfQU0e
kJC3bM14t/SW7+imJ3bzoS+MltPzoUPdtQ7ZGZBvJT6n8eCMlOmyrGI1HZaB+zs5
4rQhF2B6j/CkS7Pk7FvKTRcxwrOudYpGVeiTG+QppniAEIbQJIZIDNY+s0to88MY
HPR2PbJnxtk/Pe7JXkQY+Z6G0j5jXdfh1s6OuszBxFoQEpZ+paAbJLsYme/hPRtr
O/9dKBTvpXWDjgPFcaE3lC2WaqAC8r3AlK1KqsAlXhAfMB98gzIt3XF85gyY3WQZ
W1L7McdbSrwBTSFu4GVinlsaKZRKWk1/xIBcILn3X9GCDIyNNVWp4RqZQbERZ0p4
ZAvZXERX/dzj/PAZrOVvGA8qtS7yv2JfA3/vViPz+Mi6S63ij9Trx2zY0tXs+0lW
bF/000NubAFl6XzShADdS4mU6yFJ/LRCytqpHY9CgVRithNutPA6Xg+Yb8j5rczM
ltigbR8Shi6BI9H6Ty2ne+0mf5ZV5r8/8Z8UaMTyNiQfdloSRVhIEqdPSStFf4Fx
vU7TjJzPV+0rp3x3hGY2vLzhrQQ1yWLs2tCIjeB4e53Wp9+Jblyaoxy0dpeuYy3L
i+GFgPu1MiGUPdh6mhz8FTHDI1fFyztQx5ncN7NPJ1nsLdCCxS6yB9QG+G3NzSva
FlX6fbYU26mUWWTn6gttnjWXhs8IvW/IRHvo90gDNv7W+L1x5LJS8+DjXB1xj4z/
DOyFnpZShz8F3VwWa0zt3g31TSDXFbuw0Gd8pqatD+V2PyddDhfQFiSasZxnbwfq
wB2fZ0CIq0U6goHZx7zxYm2EvKHfTZxQuvAXjKO3JrYUOAVowZkHC/Vn9ciM0275
ZEccY6e6tK009mg/oVo8DJAxncYxs1aewLmv9P+tdJjAsvZ/s64pNwqsJ5d/0/7w
GZRfRHaz/a0XsTfnLLGpkpfk6MTdtQ38g92V1nGcd2OahEOQDvLMAxS50VrJxyHy
C2npr3RUXYlSz0mW19RJG86OIUyS6RDfHyUoSP9LNM2CeEEcHwX+mHI5djZQEUvW
YgOA4BwFCl8Gr9/1PGW/ztxgcWpD+PLPMpCqpoWcbU+XE5vuiwnYLBKPLij6LKTQ
dSlUuPWmWtOJKEvxu+VBunx5J8lQ0J4hrCwQo+JU7cUUd15u1BMJRKcpiWdHxXWh
XSzuSj5QOSC5E15aE/4AaXdocIkQHc0tMhiMgPF49RVXyacBjVvhltWpYQ5/pltn
JICs9VwJS+AYbZCZ3KXxn89nd1nSsOC8EHItpLKii2AKmDWcGl0E+p/YydL71yZ4
j0jPVisZ79GhAVdgklZBFlqt5K5oPWt15GCNJw0GVp6/c9zAbwjXK1X2uZS5B6D9
CpIY7dQNzAeN+GhKp7di/7mhYouRwrPyzgqCvy4Mfx2EcdDLrcl59KWiPMtzxa0f
xowjKyQc8ockipdGK+mvChBhEReIPwJN4saiJ6ND+JCRuA5y3zRePvclsOFjsTyL
Dzb4X2gMa+7aiekgp3vhmpqyrpDHToPgMVMlXwqT4NgfM8xxPaLfxbxFRMCqi4SO
xS5YCbOspObC7cDdGxTvuOY7ZjR2qwQH25TCjmnosGyg1FoT1r7Tkrsjp1kNZY4y
4trxhTzGKuCIRfz4S2qLO4wD6TgmLmDSmofhzAP/iRBYaKuaxARVPgezLw6eyTvl
qcmZ7BoiAemknRxNdsoVz4B+GRNeTHPEHiGAH+RRT+ZtrtkuUa8oTpXJ/rbcgpWi
fwZKxvfYCztvLOyNyTen1MK3ybLwWlcVYF9pE3JpCM6u2CD9AzFL1964x0cC/pu2
XgUP7Ttjbyu5XNZTZ7b18Yqs9b4+xPnTGXQcK9hd1jTAqjzMc4uyPFjDTcUSmbZh
RjDk6ex+0HNivtQJQlnX/6Mh/H2hTyjBxQdCD0mIkxqbWbj+i50VFm8fW31LMmq0
PvyUR0h4pciPEiPpcXK9q4j4RUP78fS7HoRWN5gfGp448S3x3pJPWFltgn1X9cpV
yjICJvfucUyykUSxbeNgWe3IWJ5rLqdN8wsOlsyhPx+qjvnEM9Sm6kfaCabz8mnZ
9RCYe4BikW6FUkwXGrkMjaAkGPdCCLfEpsMQOe8XWZgwFUKBpwVm8GmX1WlMrYAA
450eRbrdEVNgxaQdS6MUWdgIcUsYF2cqJZKerstBjwEiLrPkSlXCMmjGk1Oify8l
W11tyrIqLXIwJ4m3jGZ57CdeG1tgMJYep5u6gCL8dCLhOE30cwuAsA3lz2M62gbD
ctdG+1Z8pgwEspG5Ql1tMPv3SfGfoEsO7KGRR6teLJQae944ZbMD4Z04gvIeXXl0
LDxHKji++RKFhTBQ9d4osLTbJeBfFP5yiiJ9b+7v3ifAIxoCswm1dfd70vLqCqRx
0pHX0bKtsKtDhwvt4nvvbHAfJGuEUkmI7I7U8srEPgcPkkT4ggxpfM6J5RxtU/Qt
ybbHiMUEAda/1s1LI4xNHfXyiaT2TCrtsL5zXw2FPVGtJC2o9lKcb+51nzQcNLrd
dSC7zWFMg5h7E5rDyqDC21TfjQJF8W9vtmxLedmCaviM7gkYg6coERIdoD7AcYO0
qdCcvAO9LvslD7NZXRq+LGQcvHWchFBPVXLTPhBfenTx6ZGyuwSDUIQATRrQRqI/
gx4AcWgBMBUtSSBjUuwxZEi4BripomAnQlSW/dM+hG6XHAGx/FGZYvy26TUt4PQW
NBlkcWcjU7QjuSrWwGEakSGTddNy76Msmen/RiQ6DsQS8SFZ0ClRZ1X7S0OqZj1m
gOZ77MDmPnYOhwSQP1VSt+Rf661z6sj7vpNdsK3icTEVNcXuLgRY8ib3kiFDa7qn
KKsnrer8PFh91nv+dGdCAafd5yk+gmHwhz670BbV0gu1LersvEW/HWJh8Jb+hKXG
14xBR54pAc9QJeI73kikj9M6LCHVFIdsayW93N04RT5ZnPggFeF3xvVbOapOiDOm
jQIZoQf73gIfiAIBg1hQzxFPKb6lyj12n4Vp+sjcBF1u14rVc0cYxF6e7SiVYTyt
1SvOJlA97dhAo1rlzdInyu4arqQjIzvxdmNCwVce8mKsQBGSFX/WPnOsN91za/dX
1YDqlgsiiwDgn/PTJKoIlkmmOMYX7Y7EFVU8xWoANSE5oj+5rUbSZSmMOV1/uG46
e55XNnZ5ow7IsRBdMDyNWsO+kesZLU2gZl9yi6ljO5Ym3VCsIQlzGMZJDNJ70H7X
0iPnT9UpKXriWN9/9gqJs9sVKDCTBKPASTbLZZlIsTGiKuxotT2jkwjl8yTLwNB2
9gHaPQx8VQmAaO1FAZBJUAsTyQ531mPad5icM/pT/8/WhpVDFEn9SgQAMNVyAC9+
pZx6Sq6u73QWRSp+UPKYCyYCpZCSh1on/7UTDlvuzhI=
`protect end_protected
