-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ypUSt7tB8C0ufYPtWUMWBiXptkhWXzjZwod6ooDFNtwm6329KwaTGRuFgrNzD5YsYYQj3CM8foR1
b6Sl/IGqZch2Mdvzx9H1W9B2Fl7K6FBGgkRJyxWzEeHyb8ruKbjg4KEDO6/GZRL9U6+BOUc/foZZ
8h/KjfV97HelB9P6TgwSo7ew741eQ+XlERHxnYZSNfKNSbkBKGtu02i/v/di5a7lMdvBST7Dp212
bJ9cU0b8jJouC3Xzu+qRy2FY0tUIlw5Hc8CumejGzK5ig78ZtDMt3KAz/gGAuLUVkZ9NywWUkaPC
RuDCoxUFA0BRM2qU3tJjSOly09/GXdTLWYMRlQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6096)
`protect data_block
/mbFN7mLqc9sXZHORa7HEYFjB8vZCGfceYmSJe9I/tg8aew+cZz7YHj4SV/JV1rCWTfBFLmTAZv9
gGLRoesqPwcNnTgUxLZtEGWGbYw/ssOx094joph2sTKPsC2xyM7gAaFN+9ypS5+s3DoB7l+SHxEp
vFBrKkgLqEHk7Q1sC/TEPYz/Z69txU4pA372/dRlM5Q5LKmW9rY7F+m5qZshfSZidHwq9epxGel7
XCT6kvPp9Taxf/cOV469z1a+n9WbfaN92Rg7OyVK1ln50nXgNmauAygVGuweZm9BW3sEV0+DNJfU
63KrZFC9B3dyrwXhXprqC2TlwP5mlrzW9COqerIsFC3BB6zBDJUNkLWcCHFi+8pmGAFs17wDiPlu
evMowpH4YoXrPaqQgIzBG0aUnfThYQ9Z7Ry2BI5t0ZhjPP/hre7bthEE4pR1AVUsddgqy6Jc22fe
YYpSjjVbSyVru0umWDOSH8Tiz3hSia7xRjAG9i1oMQImjYr6yTWG9s74G/S+sQn3/ck4OKDmwSnl
7+7ynQsTxVxz3ZQl8IwyE//1eaNSOTXZtnO41YDvQ9dJEvRClg18cPB/kiO+DPqDUsdkZEYWocqe
IKj3kXo54teebCzr+widLxt1ZVlZ8e4ztTV7SyiEAHNnlnJXafbvrBj22dB1ggiJwYas3nbRIsET
iGIPpBpJ/tfbHQ8e6+WXfcTPZhq4+cy+y1B/+iv2GD2DYT8qVX4DrXAb4WDBg8lq4yHaVnzMMjcZ
PvMUOzVGmHWGKbXZ1CBhy4n09Qcc4082HJrWf/M8sRpElVaIx4s3cNAGq+vUjxEDqTztz6VD8UK0
7R5iGTh8UID+aWnB2AwRMXfkLNkUO6SH5XsvK3DGABC2xO1Wq9Nvb9KjJmIcV7xL/2ksES5qy9Po
b5hyMxqiAjPK1wPbGGeYeCip4jMFpSEgmeYhNorQn179MNi77cBuXpzuEJXqmVG8ODjrZzZT37U9
1uKIJi609QmKl5HxtQoYUj4NfHfYV6g3KcYueFCcP1SW7NadtbsHBcetTmNYuPUUDtbio5kiItpe
jlGu6TUE3TXXsCggmNo5fxdqL8xHAKp7RciwAKxrv31YH5Y0PWSqFvmvPNubC25zGUhJfN9FJRCR
J5mKlx/lrbANlimJDn0Wb7WyIB1Fzh9KSIWJg1k7i3adZJJvge0kw9QoAUwnyVA9d1Z6QrcrNCiy
2oV13CcEgAtpGR7rG00XavoikFXkO6OWjrfNQPzNSJBwys3nXzyjeB7H79T37l7XO9R3rzIDNr5d
IPTE+e/Pe2f9yvDQhcYPvrq2o4ORthGLPm6HA1ym2dqeTQNvGMEHzrVft2Apc80oVCr66qvo7/d/
1Q/ZaxqjtLDsY0UVychxduph9x8bKEovPhWDG2nRfiOwiIeG8qgJ/6NBwitB8NTuHiNgz27rpsDi
hT7nvhjK0wHnm9hFpFe4p1vFzwDvC1UE4AeGwa8BzRV9MbFDuH3gvdq7v962vBFMua7CIXlN6zHc
CtFWwVRmDjR83Z4yuzxUCPvo9rF/tiqCoIgDSp+ADdN0WCiKGxL3QLJesereo8/yllxSyzM9tUPA
mG3tydcmzhD6Cy7kXd9g49RY7FKUDM86Hh5Y7crI4gtZGRq8H/ollDMrbJiYwQwLuFQLyQ2DWNS7
tbfmDChfUc8K4i0WfjErSJzHpSkBUADmuwm5lb/xvXLdn1zRI8pmkiECtHSKpVzE/mwdtPGlrbXf
I2ajNupAAQ9twFwcz8w+U2Wb2gMElrpmGxKWrMb3xhO/gbVVIJ7TRqC4JCcVkEVXHC+LcFk5YQtE
HvMuiCoVK9kqGkUya8RIlPsyiDx3Y6ZHiv1mMMXK+m3rCfflXGlIJUnUQAYOIfjX2bhGUyTvob+C
EyzPsRN9wqiPRc9wyO6Q37LNM1KYXc46jVls3RYHTN8IS/YJxolc8hsQcBgZYQIqx9EtVLrpiEMr
Is50DXvngCAeOP67jFjTE1qyeLNMAJuAJ/1z22dqMPb34T563VAlIpqyc3VZIFYbPIjGqwPqGAmV
oP4B4JkcRWH0eNoQW4nLQUwbBXL8SlUkxrUIXAYCeOPDTRqpIXM6rwNdjSgkSNUaHCKVq5656xon
Uhhdg52+FmmKhhEeIC1uFSyzcZmzxNkq8DhoZq8UIg6sr9186aa+X+/QIQc5qLYmJ2PC/6RkVcAg
hSMWFmvm7BV7VdbYGqdmOzSzM7L9bAm7YdvhuT2xLwCxE/f8oC5DxQHbKYSaO4JBiE4b79S6J+Bn
bT0fw0xaalOOWrchKDzKwP0eboXkt/juV9xUCaZMJXyyPKyGFmFY2sGwhGT6mRLLUCvpgl4pCc3f
OV3XVzQNchjYh72HeSTk5piV9lVGIpUHrx2EKI/9/tpVGqF5UJ3IhvZGCIFykc5qc9Efd4mXYtDh
RXdbx+QSzmxPv93Hxy2uVFbeGTIBVpdHabrHwQR6hbAOl2dyM7YdTyM2EMWCEglFGkRfLyDEUBg4
FfIuXdiToYmAgwX/9s8sq8eU7FsE9RcoqgAjUWKrBRUOnFy3Ej5VDt/nb66jcAaajqym6r9Dy0Wq
WzpbJO5s2jASjIVPRH7TY0iM6/Eh+Yb0MaMo9wVwKPMnQAPjwZAJpOmD9oRuPqGyk0Ntgdv+Q42m
QfV6iDykGRsTh8Kcl7Mn1DeWkhd1e3/BuTzhW8oX+BiGdyk9Yx3RsIaRs9vkgSAW+d3OWOosqesy
GU6OpSo1jYmV/BOnsm+kAg+DRZ6W5l/1UjrB56+rKw6d6yMSmzVaQmp6Ip7OSc2kSmWodfTKzmDj
L3nLYY+HERq5zot5nYa7mBMEr4QxaQkTUL3B/lVAlTsHDpA9W9tUohU3V9CEXaBZYWIis7/YsGBj
2UvK77yLSbDMJnxU13Q7GLlVQD/uTMydp9/iOpGV1ie+tbeWpSr0GpN3AchuBnZ3JdcIYyDknslP
VZeIt50rDpIVtWAJJDCzIGrbgPKR89il2knPFmd0w7tOQ5GsMteP+Vhzrjn76CkMkhCXpgPKklzZ
P8XMfdNzRvc1XCt6jW7ii0mdf8oC7KGC7Po7XxBcFuPtcdeC5L2tfeiCCbV04adhepDOblqAVTxb
0H1v1dOiirR7MKqszG6cPdTjCbZhrq9qGPABkAuxvEP1hWheKi3PyGIXNC50i5K5kzWb4uWeQ6LD
LaYa8vKFfko/R2UQEM/ul8DhOsVtOpwPGe8+Mp6ULqFdADBIHgGq/4zdlEYouGJ21MOAGoMVupax
RzFtJLGVmSI+2IDI7xE+eCMlHmsc2sPjJglo+MbgixOArDxfbR1UkoJnBMebnJjNAWw8MZbzq0SA
a7FQboVFLq+GuDLFe+gC73OHpDzsXEoCfRpxUBL2WFSFG8DIKW/X3iwX6RPkMB30XwqNWgYSpTQf
5tNFwh8l6hChUbT7+hlNUM6x+mpqFFwVJg1alTvG2cWrRWGZUeh+qWTR4YGCk6JnQ/ofDwJDchKo
nv6D/MGH5cxSSsyMme1s/J1VYayHoBBfeu9Vext+dqxtgJbO0sx2whbxOu7OvI3VH2bC0gEiav8N
mdZ+UWgq4sZDvMHUrPqZUdx7BauZXwW5bpq7zG1VXoxwhQv5FhA471N3FuL1YPeOkbKGv7vnhxLp
DdfInLmj70eo/3VfqGCrJjNN8CWGWx4RnTRi6L4SYwCt+p+8yiSNWRxljXQ1qrltJ81sFbpMoyhb
SnzpF57xHOtYK/3ZPOVkrJxN02WnYMR5FfJZ1TvakqFNKCWWYvDqXp9vROxXqvY0xW35wHXdU8xf
0SjUMk5GhW0kMd8s4B9yrntlV9pc0nToswBk9SjTWgLZrhfJUKyMFPkMluFkr3/OhUYAe8fCiRGZ
LaUEg3SsmGnvDWCJI+e3IwSzdLeiC6+fRBY+HR49cfWbds3JHXh8i7XsWouJk7Dn7gm/n9ZrfLMH
91gG0xHxumX0OeabOtRwYX8X/fTIt8rsY+6s9FCtQfrxgEy9HFu0x79tOR0Xo6BL+X0tgpugKRiG
vdhRa3/RPDfreIDiPLkn9XJh6jmGGh4C9FYtgI+ixCdz/b7qZbfFBTdlfsbCIfTSnQHAM/dqoDPB
TyBqvGVmKx7SvwA1BgO8HcUg6Hsj/GsoJErOYKThZi84GjbPI5Sfli/nGp6Kfjs07LCPpo/Jq8j+
9UYjheDkoPBXTsyS5iJCk60egS7gL1h9VIckWUvjV4uhKB42s1AkKhZ7dtYt7EEmq/2TdtXoguBp
1XTjXSXs1SFoDzXlg41kf5awTux7tabzzPY0Pbjun3CetUFbCxC8AbC06BlWPHVt95T8mS6KWnIF
9StOUdsjGDi246jwvRsok1x0/Ky1EL1ucPkspK611UPZQeNiQ5kaCNsEwnSDI9z5TxkcfF4Yd7Hh
JsKVHsw/ypUDKpvfgQ2kchNbtrTaNznI8QUqdIQFERW0B7wysGUbHiBkSbvd9TtrAg8Ea+Uti7S7
ONReGAeKNV4hJJutEoivHS+sbNmvOC292N0PyxZCYLnOsejifbeC0GFRZpHWb1Zxic9vL9m4iUdX
dQVObD8qBFX/4yWlCS1PEQdPXIys5AFt+2Ae99eDP/AqkTVerTzxepH8Q9huIRI81/lDka99wIHf
XHZMPWkuRnkgLZU4n0kiFBBPe7UNkfzIoD29ndiuritgrT99yiw2FMGjnci/jFhp1vKNkolfHKSr
GbcFvEVX4hgQ0mjiiBiN7mexOdgissjGXlU7QgYc/04qaK1SNkt6lExNACi6YhORj6SFBL0ZmxXC
VQjn26sD/sGIMCfLYiFeVluPpuhk2e2Z0jW3+KYfVlkhjXig0avkRvJRZWPsusMQYWTqfVBiH8cy
SiS0ekmLuR544ovP5ky/dYS2II6M3DGOYN9tYyPhdIfvFEpc72nokt83LPVXE1+DD9ZGHNzOI+o9
xvxfDO8cA6amUVtTiwT2DgMDvixESZGPHB2dk+ZJtEhAo2t0lnvqdywKhis4gQ/q+soEF3i/XtuK
Y5/X/byt3VWpeE/Qwpe5GjhOxISAUGW6kCbo1e9VSQym3rNNduhGiC5bs24g4Rux3OsQeCvR8huT
m7L/uuOR7MZ2wpoULHDmx4ioSO4TCP5Wc2Pz0aWu5yxiJlYksYD/CZxPaR6kCipOWpwKxqUwtYMh
hFhxg/dVrQiJfaDiX3cBdtYsgbRgkK+EJNZpgEo3n7Fv1cBOITAj7/qY66CyAAFnzoofZzYG735H
HdRcGV1vt0/rhdsweZK7CN6pNnGHlL3zfi3gMuJ1w0ZEkl4aV70Uvxk96B9a6OgIxpBI5EHaE+4y
up6qVo+BCuQxNqzX+ojYDqIWYsY4NFhqGQJpSqEY/piib8bsYI5J471m3CroJSYRjeiuRNoEYy5F
1WfC7yBth/6wHrfS+rH1PASRyKi2+/NnSJ4mRE2FgcR22Cca3yKq9OHedJhdQe9tSvohE20FV73p
6EOe43cdCxtzmSc70KTB3bbS6r8wEZx+i2ATRJIkuBNJPSVDGRderkZZFCOFPsInLanPusJDWdAI
fFCCwF3flD/IwX23yx7uneQIWtOi1QyMzq55ggJtNXLKhmMXPwVCIpqohb+V1E6LlxsmbcWJwFBu
J34vt5PY4C+Yh1iU9jpCIQfVE3G6ApCAkSOGzIDvcRx6yfmrk7AESMOaDqesaEhVszWuOQGIPzcQ
DlQTT/dhH+KZ3Zvalnn6kuA6jcvSXGPfFd0Pjc7M1atIosKYkQCtbViiOhVIRART5y64oiP8n9wz
hzAnRgDlcU9WEoITtj2WVYn2JqDR1aM6T85WF+apVul/mHPK5ZEyrde+moy+lk0IHz0Y0BTZfdDd
X8oT7dqTeF/buF5LZ93iTE3/obljr+/7GGzFBR0bRQJCwTCefFgpj21WBu3eC2oZoo1pFyFltsBy
SP1yPnjohd/V2ErysEz+0jnBD5D2QzysCNTek1cKNd9hV+ZZwct2zBTSPOmobCJk/JPf9zAs9EE3
QDw+yNpPzli3/g9+FWt8C4oo8er6QWRkdP4JznukBZU4mFu6Ti/pOVS48jV0Rn0/RCgH81Eo2Kal
LeboYJQ+2+NOFP65y2hTrOpECFU0QFiG6k1DHyIELgIPNNzgUugjvsAYvzpts+fcc+3212nkW6i7
j5I4Et47rUb+bGx4Yk8y7iUVs3JHVVbW13BPZJZG/yOCV4qVqZQuSiHtZlxqKGXhcHAYyGYNSZnj
enDtclhqvjEy/BkcCTqllnWdP8AdCS8ts9YN6xIP3RUzA1mqtb+8C3t+Vm0dGJW1kYKF/enc+Dys
mA5ZK5fmPAukCTD73Atj2UTnSf26xJOw2v4tB3x/hbejOAlU3SarWHOHB18/alYXRL0uKEeA8o5F
mykg3W+5OQn9uDYVrrNtZfw/8rj26l4C2rItjQR+9nyLwT/N2FKw2l2/C3gSEuP4eyxytISw0b5W
x2SwS/SA4AvcD1MgFI+MqFXzG6LPJVDgUsutZudUv6iz6lnGN56tu+9kavb2BsuFIo3VXNTIp9ub
h7jkYsyY03Yck8aU4CZo58MH8gy/h0ofWYWWcwPkfdwzRJK8K4kacEpgrak1++3mgu/nvMQZyxOq
bHXvQSlGPm4WyrujG5vgaFGBFIq5l49xJNOYcIj+DhJaocoD0g7mXd9ysmKxp3qKctCYtKcn3wO8
bwMn3JNRPYJEP+xiEwp6kYZXx0uX7gdvcaRxBdfbMm/XOm9AfqwEL26h35vk7JSNG1QW3f+0Mwy6
Il7urQ0YIDCjuvRd77AeB3hEMaPt64wClRHWGe95A+q0hye4K238PYby/Rh2hKaZQjblQqG2NC0k
J2c/fgj+aoh4tlAaMKj7zDp5mokMLkqB2a2ogL3EQfYnHddcQkgtfDy2NuFmKq1oRztkK68YD1TH
MmGhN5bAoVLnyE6ZLFzoGs3l5QHTxQ/6qXJS59QhT+I7nuJcoYCM2lHbQ0SEh5BTx3WPiUoGYs55
DI7bF/I6e5nrJlM+O3Us4hx6MRPNrAXJWFieTZAdFwzqZpNzGWWG+4KILiYODgxFuny4SWW/+VMn
fOHTfx0mOCvZdEMsxuPBo0hmAXoWSstF5d7IP1r15Z8h6KkEffADi0vxyMWkdjbOVtaSGsUnZiQd
grMm9CfpofoBwVFk7eTXhtniKSbS/kAxZ5qOJaxv8zv2s+BvOvbQ9FYn62imkTvZ9h/4aStR7ysA
oFu3lPSFshKzzIYRwGEBfc7cR/4g1o9AIRYwFY/m567QlMDpYmISszCECxpNn1nQ/rsrHhZpzIWH
F4GoBsAXmgJtpOAMQimLGaIJChOXs1tTgRLlf2aDtECw2zdeVDrn4gbsJ5j9oIOTJ8kBMYEZp9Dc
JMa2+3jT7c9aYC2hlVOlmxxNbA8hOzSwzvRrcy6ZIlZo3W4JQLbSJr4S50GQysYIxJCRPhR4L6s1
Ibpa4mU+Jkcaxk3o15KdiBL0vuFC5xOy29KZU402p2VmiIyJGOBqYDE8Z90j6FBNseOfb3hblVKq
L2j0hZL5td4xLH2ijLed8EA1Kxpq2Ne/CSrhZgo35IxhZuBhWOkwxNjMOeK5rT7kTXfILxXO30Ca
eP+NG3jLzOWZfH9eWXKVtGYGXKj0n/jNZw42gELyEG9HkS/fqYM5MZjLDgDTYG+LQlhUaiUJZgqc
hNvKiief7lnbk6nAC2uv7WRL9741rPhoiD8Zbc36cLP71svuOI08dWjMSE9qsu6t/ruZZmxDQV0X
d8XVwyRfXy4lPuZ1SRD4ljXB2dH3fOLykuDA1MZCO89aMi0rkIZOv4LBkR/pCSdhTJxe2LOvTG27
N/ZASvw2S5AXxH7efDW4K+4tIzxLZSKasuKY4bFY6+Yv4OtMRRXSpywqLvKt4Mz2etZHzlRocolZ
5lIGlk5YCp2fF1zh1+LJzUxbtzVqJHEKvwWvoIvzg+Kg8TZ5gy9tdE1P/1DdbOlS30QRk+TYYtzd
Um145jNcgn6101JcgDoKxU4JxHPzxcs6Kw949Ld73wl9f7ifU+3VTJOKGKzqWZ5Q6SRKmIIA+5ak
PmGiyKVPRpfB1B3NJQaF02iKp3FBB8K2OTdCPtaZ8wGnCexuyOTjhdgBJoi3S+OBFlGoF3V6
`protect end_protected
