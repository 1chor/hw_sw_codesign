-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ILXQ+TMv/07B1TUov1gXwxlQtgbCyG9UhxUa07ysIJeeKrnEkJjqyadJtNq7s/pr
j+J6apsxhKBRavk6LlWRTOpO+GIgcyKbQe+TEyxIDNnPKkr0wQqmo0AkjwStGtSE
o04FkPVJmwmNe43VXWitHQuf1ryuCz7HHQ4fIc6tri4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 2880)
`protect data_block
yAfgKspNJpCIChX3BaKWQAza2V0zRqyWnjQqYReH6WkQB0JK/MQzmkfTb1uNH8cF
bUPV4KeJIQFLOdNiYN2DytVGFYBsjYSDqQ2aJLyIxN1MeqI3rD/TsvJMUlREg1tQ
rdYZtftXHFA+nDmDWYls3Y+P2DQTxEDPeu18Lcycuh2fs3hMqhmVq8NCCdC4R3/X
ZDenIovMwgv1KxFrRcWPiTQ1j3X92GUODfh1MFXtl2Xx/jhIEWJN3HTxKxCYCegw
W2D/kUY4qaevkAPe8OjAkk38RL6/tjJy9WwicejUWk1WchYauQeJ4qXpvN6Z8sbc
1XMrBNmebHb2PiqZVjTGgWUzHFCRuVF7XNkikRFvUl3a74sr8PUAWa/5QIXm7sn/
gcp66odiwvEniBxyGS0QdoXZsRUX9FPbiSyz6kRL/w6ffyGzot6m7vIuvQByhGRH
boNzfUd5Dn/2hnCUliVwbXrWd0IrNrCNiriOPyIeHpCH5Fe5SSmCSQoFgoRe8Zvf
R5o2DjLQemR/i5G/DQb+GJNgATDORRNf1M4ostXUT7qirlucfOH6DjxGFlPkm/Cx
bkSIhJvCGfgnRLYEkMSHfbQuCGDf5nLNcxM+Hyoaop1ZEe2K3XOJ/Cz82/XVJxop
LVR+jeSkOpEwWbvjnZBlhge25x5DBhBcLNjap9x5UHqoxys+fIb3Q7gkMF17L7PS
dpNdLIh+fKN7qvIvRiKTsl4EGlJepQ8QyhUBPdOz3PG34EM2/5XqROwUz/6vCywn
viaX/9BDele2LrSb2H4PXFUoJVXVhjbytn2NoMwSXAVq1zB73HDVIH9BmIIK/Seq
7LRbMoFpADl7s3lokTx3x/OM0d8LNIBvc2/M1R92QUp5V2RXBbDdMPV5ARtofVOU
tiJPAsxh6gjNC8gidKdSHsuqlK+W/+ua3guQEqtn75FZRRm3aci/5+bR+oi5UTaP
mmD/DL8vz9eCviLE4Gjp7G2HXDBNKVfxijGFUNXsqDGx2tZ4+jmPFMcV53EHMRCv
/gq5TfkhCCpg5I98Xti3zAD/0dR/r++6FNln/8fLwBCMotvZ2HAbCbsNjYiJRpFZ
veGzikguf1lbYHuPEx1jVwEUxuf4nVK8RJvxBF/Hvc8yxOzA6ti2zIeLlwIQrA1t
fgnmdr8CA89BTbUM6MjqmS8wVUTHB8t9NYZ875kmb3kOMZ0p1PBcaTeukmw4rQdM
181pZuZn8G75FwKVb8BnYe56O6jugewJYXuq42iZENHZYsBlofMA39DEtl/tQq8F
VUu7PP6nbp1IIEQh7bPInRbXOxkkrcAulvBuouMgVzFJLpHLsTJEy5cBhQk4o/+k
ojfrDEJAcsgfmnaatyZERmxLG603TVVZx1SatUpLtbwGNrvKkKrccYVQLMQ1/jOY
0wlnOSqVOSCz+NZYAUf/12iv/atPWje8f0BscQjNznA/OzpXipjbUCLuysPzK0DA
IBfmKi5nTWJVpeeLpMiHFJ2Phup7nb0TREll2unhRs3pNC1k6BKw2TkqCbSX+LQq
dBMpDPpW4/iDyC11o9LgDLqRkNNNpfEfIjQKnd00FxLk1n6iA7Tr3hgvN6hnBgVM
4OqhkzncITfKGifkleeRZroMc2Kf6DapzirQYL91GflWDYKkzQrWhfRA3eznxb9U
TlF/iJAxj5niDTo2+DRtPhzogRAZtuSY1wHKdixm1SAlkX09uJ1lYO7vxcWGB7i/
EQMZpnSAJdUvrmfcKXfDa5l9nOhuA7iD2J/KGzNyTDyee1uB6XBqbgbVAdowhEJy
ljlCi64gYo6GR6DvlVB09PegiI6D6tfNBQSwY6UM7egG2TJa5EWDH6oogiwdPgwz
xwGIfI1dIT+Ir+wndT8+getfkIOGtafz0yF0U9O7gRgBvxs9Gy5o8I9oCHgejfg2
IiG99JUsDWL4LvBA/RJTeExC9hdZgU6lvm3Zoenb9JxqR1WDRxO+ywBC9gcem72R
ifW9MgiB8TWACcH/7eCZwKF8W6wvxq0jD0OCTaneB1jidY6BXssyRX5il5oaT+dl
5UFNT207AebHQbyAruqxmQiMz76X8jCrZU9mO8/AhH8P/NjfCtc0z30brBLdKcyR
HyV23/SUAyAaqDtvfVZ0XB/8g0brTPN39L21Bh3VUD8Q7UN3sK56GsY4eQK3YbjT
s21ZHWEupYtIsxedl3CKzDy+xK9uGWBUrmPoJe+t2fMYBYP/5abA5CxjkNLtAmRG
JT5ihe4YmDrs6+TAlcdjUJAcFc9NXvjXueMbfPAJPFTLDprBr/YmPIGRjxtl11rK
ki3mnqqbJ0ukZyKR72HrZ2D5Xg7N7ie6rDCMhNs4yaJl/sVsIjiPzjxiQcWslR0C
ONZn70Dt92WgfDFgluHJPYI0kl5QkZhylGcd2qSKDVbgjGEdDhL3EHFAcQ4o8bx/
JUfpw/aYaGhUQ4ALpzjADKzu2WXTdPn9FPh2uGF0UVew9j6XYPc/FrticLZQ8etw
H9VWFZhy7e5cRYHPKM2KcOgu2gaRFAR8W9NB27uD3mmNKP4vj3HGD6h6a1cJdJCm
qbuEUFmpvhyVC1PbLPe2Cwdt7ifMpEKSvIWNwb5W+ayNXjwNFCQRhCXNhSuz52Z9
pnqjqaDxw1RsJHTCLrM8ag9SiAzxriww9ohWJt+DKOX32EQcL8rMnXgCcmQAVmhs
uhX+QJTIcAKNO3hVhmzLlH5gZ+G3A9Iwe3fNMKYcWNk7yL289wecVv78iUWp/+F+
i6N319KY2DfYbdnPCqLb0IEyzaguh/L3HEdProHgnXhtdCjM9+GJ0s21YnSunvLE
iZAeCGsHUXWeVh2LfPQ8rQQlKoANblTE2GAxmjmVto9vMHX3aXDZuJ/pAvFa/U9x
1KHq/VCnm9UuPDAm8IkevIgce1PO1+rWlycC5xZ7ZbaEhJxZzx+m+HXKnqxUtfjY
c5Syf7lHyAV+LYPw3l1xo727uOdRU8yZfe89NLdFh6HHnBdilHUKBO37URIL51R8
iSSLrzg9EsZI8Yk5NWx4J7L6aNv2nFwBRRdh0T/XBVGOCeRrE6YNd6ydxWCW6Txj
aprOeQrADvtLV2Cy/qZXyFQq1hkPw/NtNjDQ1CDZh5KJJpY1nSd+Vi4vD9f7E+A8
cBW7uuGBI58eHJeHVRaxjC2KOsVvlmGomNvoU8glwydqsW8GnwgboAZPQXlqWIj/
BYeMMUc8awTCxw7xTvaFUoDznDT7TP8EXJZVrlLheamJkd0xkJqoXrvSvovg+uMq
y1RZhyFowWQIV7EV+8KUcDEgIz1dHB1nG9neAcPHMj3ycY0d07/db7sLUdo9vvFL
g0FES37n0/2JeCbSmBH8zFdmwlbtPWYM1z2mxPHyo6EzQppVpMVNZxu0wOHisoZY
ibZmd7cN4xPf0fyyVWV8aDBlVboShrvMn8dprqxzAqPdYi0jxKhoNKrZXaNCySL9
nET7XALR5xj9hWqMKcUpjIjCx1vDNrarqVBH29PJKim20J5YQFpXX1QpGIgiTuyt
IQETuObtOjepWh2V0IZDn+lot+KStW9TkoSGaM1byAwcM0a8oQzn56dl3act8pq0
6Z4vkKeTbbJxYQSlHKDqfKiLbs5OyCn4+xUqVkGIudzxp6s44zwF86Ab9XFvsUZG
aBpQnhChoJv626Cmte0ZSeRFEhhtaKFeFD63rBT7xUtQBbBmXzGtAFCEU8PDL5Lu
t5beKEvRBVGJOz219LVWh/sIsOVDHlNAK6fl3YXcsvdRpinD16Nr/XWUeLJlQA2Q
I/yrl5dYHp+wHobZln0/9oxQ92vIerMt6unxT7Rw4nN/iJ/uicbXFMfgoKzxhWie
`protect end_protected
