-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
oHkImMDeA9a0veDRBgudihtGheFK2+2MPmvONT2W/p5mOVU5CZxNNN3m0kTZNBNb
clRYGpfUJXb7EyqcQPnLaYJ4YyjylNLjg/8N/NQwHklzTOT+2wA+97Vp8PbmYLhC
gaOF5ZFCBi2ercJzxUXuKLD1o5VeMgWKj6YCvdSklgQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 2912)
`protect data_block
/uIdU22fsIHtCid1dTzcafC+09exiw36hsJ2ENCjLiHuDqKJSOw0366LJRJWfmyO
IUXKcWLiMu4lWsdcwWqNaqwt/5qkw+F+kZg47p9vtrQQRoI0EZaPVhm6Hv/DAK8c
9nvxbPzQKYt6qJPVnjNaFH4eimvyNWceM2oCP8p2EFEON+ys+GyCjM15GXQp/S2O
iqPagkw/cMDd7gS7JQhZpis/eyNK/vFEAFgcQXzXAJdmald9vsb1Y0hHgj5yKl1j
y5Aam0qs34Je4WlxxstVmQyIF553v7lQrnPfpeM+1lY4JCrjGL9j5f9hYzXvAei4
3tZLm4hLx8EKVEa9xvA/elOl7oHM8FEvAxf0bLsadw60o0Eij9OcY34ZXICBgj6E
NP6usi5Fi7fGnwrfTuDzMPKedB4TpQHlHfa5Pa6t0kVH6YATt+vpfXaep/N6Eoc+
/ZHZEqlOvFPL2qMgS2uv3egNl3nhz2Lqr91Qo0N8oyRQ3ScS2nFr57QDffLCsQRt
+c09yCpbiTF3MdcGHBfajXDl1GMO0cNQpswse6idiNwtQ4lRyxaOdBkqqabMym7Z
ndCs9A4raVoBE/cBE//KVWi/IIIbbgeM0E9p6ALKYvJN3APQunCIezdTwpQOWX6e
wxebmVySyfutn0hWITBcCr/hJO0a/afWKWAaFpOOKvDDxmZZOljpzMFxNzEz9pSf
A1bATDcLTfFz8CH2HwFMgHDBu8zLEz7Zd5Do9gmOR+W1RQJqcJTSTbxzVdi0CHdR
+ZY9PfziQ3nYE8oVqgFuh00eAHfd8nUG3i9fXJGS87zDIP5246rW3B+OvNQYVqgC
XEae5NgPLocqlv85ikskMyakzoDgvlKeQDzWBR9wbDtzQ3o2ommqzGdYmqXgtwvS
oIdKGsMzFNQtdOEe4E+lBp38m/ixjzTcLfLCT5U18Ijh8Wdwp8XR97Gjt3HYK9RQ
1zqz0iU9zlLMdV6pvaS537Pzent81xIWJwPZ/HlIgFUrZMsczd+t6I8+11KhxFDU
ytAWe3WuNc9Z3AFosRdNVWka4vsg7r2gr81ZZ6mhOlMpmt0cVobD6Np44DPIKD5S
4yOEwnzBZiBn5KCEJfAaGkiO8C+/V2nl2jiB01Y4mJ7KJPwSEn2QtSR/KW4Z4vCw
c7fROzpSd15LDTCxu3k32DWa89rBSn5HwUt9W+agp7X1NUoVqUF2+0Hvk7lxJ3Wn
z0AmsUS0VFR5D/97Bu5NuNtJNyV0euwviKplQDtUBMngqi5TG6uYlRH4aY1Er6Kb
2SRw/OpONT9r3eIqdCKVXF+ea1v5GQGwsS4yKEG3vjrPafImWqt3laFbeB1GIA7h
2xNdl1r63QChZEferVVNrHX02y/piVGnC+kVHTQ2LvZlgJ6oE22GVN7FH77PKQ3Z
AdX5rjCIjMIGxH6dHT9rRFtgeFjTucCc1DNrQblCc4uBLGL4a6Li4g7TdRpNDL3V
//p/xhhlB4CvnwTCyQUlvp0fKot4sew6uiS1RMjl8t4/Xl3EhVG2VBBqqOCcLBS2
16gARQoxgQGvFPyOOd2AlMj47fvVd9sMzRwMEtuRHfPpLaBceL20yg0cYR7ZodRD
edoVZkGf8Axn26Vb7X+FrQSbz4EQS5lAAt0l+UhAGyUDavNeoNHnOlHZbWCUqdw6
VjApxidYtzeBmvnC3rZ/KolSo0uRYYTTlAsD8NOB5tNXSVV9PaHAeu6bd0vVfiPr
gRFicywFQ16jiM2i0W1zZZZYnHuSxP+zEPy0bNwRb/JKp7m2hdsHjOZIAPi1He4u
HeKrEzQ185ETPvBhWQ4b3hkt8YNAAjuk5S0BKwT99DPHDXxt+J5tNGLjAgSWsE0r
QdzM73MlEn3LHcXsIyLxDBSp6OhbLzfd2Kxu3DrIb58R+RlepjR88CAfCWkzusEb
b1RS5qtD0CjEpE5kEfQEGKQ1ivfGDsAoBypjEl38cYEpb0lnxsTS7Q54hKuScKA2
Ov7TBz+cjbAbWFqwQ/F61ikf9wm+92CEkU5AWZOLDiCX9VP8N6hC0gFzjASc14KG
GWjK3C5+MTwAA/to2gAnRcOmafZMtFabfA+rXMXmv1xFdylxg7m0Nrg/FJN/OoB3
8FTD/GYZhfMy72zEb4lz4eLyPo3LjVXTQaVmL4KphZCbpE5/pbXf4HrpA3hDixJZ
kalGgmeklhivCLqzYtf6H5TaXMj5GP0KlgxSwtR9r2acx+TdvD3eDajsZl0PTvKE
MaieiUac4ZCOnC5IfbfajGw99st+JuFDTa7VubSM6XuwKJJIeXCn1emez2ueYdhu
rfKTVA8aQiPL9EhyxJZkyVcc+UVoPt0qpdVX2+01RRTeFuCNWSye73VQa8jFk+/D
xJjVJxbeLWBnuT5nZnnaeAmXDcgiiCYTPD+c++oUCpVl0fdJ37T8HWBgHgnEP0w2
FsCqdCsRc6evJUvXjOF31tRn9ykWzRIgbXVFCgN6V+hRDt8LIeWUjeCxCOLhWJB6
gbNvCFqjgzGthpCpsehs7xlJlzZAtB76sGrGFa9+tpGXi3ZoAR6idhsnV5H3xqD7
g4Xe5w9Wk8Pw1DTRqLVTuIhCO4R6U1jANQLHkmbAITu4pnQaE8nPSvHKZTEfB9dC
sFVxul4GLWwIUtmxtUIzvrVCRZvw2E8EZUluAD9N2jpXLFSocZ8Jkj1ZW14Cj9oy
WCWrla5uwhiekmpFxcrMmEL64yriAB3hOIGJVEz1UbPFP5YKZInFINxTSj/XFtyT
VuuqPH5Hs64pX1hiSMw61ae5CW80Oxs4RbyxTmdmOtFVxi4ESl3jdWIjonCaLbpb
31woO9zQYYae25rISnh79K0YB0kfvQY5IP3ThLh+pZOqlG1YtI+EoLykLJPVL0nF
s0EzYI2WleAdcRn7tqrTJE73wLl0SMopxeYp8ij+hTeA/9IkXhkUhFBzo1y8KoPk
tojcz+2XLhNlLMJ1qjqc2gTCzGNr6uZL+hFrhTMdq+OErfNyGpS0puhn1kKoj1VW
FgoLOYci5L+ncnVm9T7f0Rgp9yV04PayEbRCosoCeU/BppdLHfhHwP9Z9h7qf0XM
aiP5C+b2jxFv/D5++SX3Jv6ARE/vVdv2oIaLhnvOATkG3El2jctC5ZLkhUZ1YLW1
OrsSXlI7bzogfG4vcipVH4QupjZuCL87vdY5dwRpWYBp5i2CyutZ1IeomwgnDH4T
QLE1SQp+6Jvu6lS/Gg8YG4SsNrjdCbOMOVjIu80ciUx9/Arg4ztGnPNZJAp9KlKk
zR6ipqKrSzhoGgpEC5AvNbjp2oNiN/zeI8waJG/zRINyftmM5VG9IJJPr3g0ucJl
y56Sv2XDPXfJOIxAq+25GeV94mpW3UcN8U3S/GXmlVVupnZy8q8bOH61LahWbQpQ
7Z9i2ZJCw6PaQkJcezDYvPoDxX+hY2EspLfcuQLgufqIobl7H7IAxmVq98Wc+hgA
Cz2tP4WW4jrK1V0llk3VZUXT8HfpOs96Ev868YYt9MSW8g7XXV0+GpdKKyyeNq14
Ud+Axo7ARbkguj1RfrMRbhlKRm/RkC1PR8tkKt+mLAvoaXX99xQC5hN+r5OSrUcU
oTmVVTkQW4mzpTovEPZ/6mkPO3NrR5iUnchCvCqg8bsyZlubNPxFhkVNI+QUF3i+
gdmolJ7IWdSPiIiK+7xUHBWtQqmJ332paC2pkDGdsa4r5+ZtVU8JTIMcCLAzXppY
GdLldbP2Ugyges+9W+dauLuFJsvCeheLCxd4PYh6mzwhrrBfJxRqPMnY6yAFzaeN
80un1bFjec8A782shciqxkrn82UaKScY1O8b5nSshAPaS5Rfn6GL/kG6+Uoi8l1S
GDe8v8B1TMGhS57cCYz6W/+uB0TLW9SJ6Ve0siUfImc=
`protect end_protected
