-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
/CXLpRU3Isvn4BRGl9xDSGBG6eIv3k5tB5JLoZVOOt5VlengeQMPS+wkrY45SAVH
Xl/xj0MtLO9oTLyUj5hT+3i8pDnuNYPJqh5fzwA+ZriGsOmc8YB4bqbe0XmtWn1v
sQkIm4LuIj6hLUq9+YukexI+Dmx99ZsWzqdoOvBtgCVg78ONdekYTw==
--pragma protect end_key_block
--pragma protect digest_block
CQYEkpUbeUcZSxQBrUjAIhdAa+k=
--pragma protect end_digest_block
--pragma protect data_block
Qf9Ian+MG5kAYr3g372N8S+QbmtK37VphjN4umi5VR3zE09dGXf5egoi+GJ7GdKG
ILafL3J4UtuCPipc7Jx/vcFjKKErtwrwkUo8J8nrYLtyJZ+vdqO7qiiB+ckauB3w
GEFXQW/57xUdx2y9LLZXQzsz5lhNOJHJ4u50U99uuhWFJvSFOdsuemi9iB8KKhXJ
CquiZ9KGNX4KPuP6MVq7zKOlKE8Z7XZh43d03aypXi6/+BzuL5ySwA+skt/7j4kM
czku+HIvZkSVcUyfpCaRgS+HHU6yhX/I7TqV770hnPld2cFH+VhyqG/PWbsOkd38
O+KgbHb/cC8aXKsMAPKbj6szXg+T8C4Nvb5AuU75kd4RDXzm1k1u3ZDHp3wjpX6y
80mZjs2mps3namjoBpLkdQCKJBD5LZKslVtN+eoK+RsTfqbkmNn90PrX5HO1eo0Y
aW6/zEm9h28zm71/vR7vqj+HRzYC9ZeOw6vKAHUpfNnhTFh+9UR9erwYKnGILt//
DvRWUO4RDx9LTmxVOstWngeWSuD4Q8wNLH3A1TMzHiWqG88qRkGSbr5ltQMmbvMy
AUPHr9V4phraIQpUGYikn5qYD/gb5sRSMBgM07A/9gw3yIY3etypsf7rdi0kPTon
iP2zIGBgiDLvtlgkuCwU1Xe0KVdbXmXb18kGmkhZYZx4E5qTJ9gng8sTaPiPe+9m
mh1BmTjdZLULbP+/BBxWuwFOBoMNeOpJh1HCYcmhiufZdv7gSh6tekg4Lt5jijIq
qGUHNvJu0Ntin3W3doPvfEYUg+PZ5tDKxR5J7JuDTHiQ5fd/yDhNuUHiV2b2vMvA
OwDTGaxGUjvi0Etd9l+DZMHkKtHgbQyOIEROcvGC9OtyyiZ9ZPHpJgISwwIoIIdS
ToXu70m9dfXbWF40iY/FfFehGV/J8E1AMOaaA7DAG656XkBp0uKruz98LwkFpvaz
sTZ12m2qN69c+5AVijJFVm0Rcb9uvf7o5ksGes7ipPHRvR6ep+yo7n+65a7KWV3E
ghHcu6z9XA1NA7s3St+cr3+YeXTP86Ty+3ySo61UKXyl2H5YoFFHeH/1NRwkgj9Y
xOqhjxWTOjgh2VC5g/vCw8H2S6FFCOrJCwMeRLjwkN457T4exa4Sr4UPQ59UJ7vB
/OjlIfWKpRwxYHxmyT7NDimept6tdk8K6XRMWAz7sOAV+xZya3Czd0yRWg/NwSK+
dtdZ1iMqFKsUZepviIcNxSkOPu5CpUaV8v1JbGqigUMuVa5NxatAe1hr4Z2lRfhL
bMZHfLbxdztgWDD8OCUDNR17pp6Mvx1eHEbNr/DtVjw9iez1OadgieJ7tz4wG2r6
yEBNKUgzMyj9O0dsxMHgpoZ794o38XARc6icaZegfvFVgrWFBqtlD5qbiWCT/29Q
q+ZfY9V6UljAP2k+jrpAfNGbLfZjdO9TSJCvgCggCEJcBiTZ1nn3AZkye2swxmfn
DzYQbmLJwPX7I1PxFUbNQtUZXIFf3zenJ9uZGxFUpqzM+3C6YVDOmklSEPHkA1KH
qLRBumEyExvj8e4wJ0bu8+cynLrjFvlbi1HZXKyWn6zQJ39WpG4AAvACS2AkezUS
Ge+lhUaxZGYu+LSUP5AzSjCGXU4AKjNJH7v/rrtDqUld3vphuh89b03cf5E5qU+6
SOKxrbh/ouuYyNOUyce0RoM7eDybdLjHqYffz7KhZ87K5XNHTjLxDHIzDKvG+Xe9
lOmzWE7rgtqRssHMWYmDRT3LjQWBAHW6zOyRLnhuawM1yr9npSyPX1zblPXJZHfK
XU67XzGyHH37ZogZi8I7htjimQmaSdKYldcNW3etsXRoq/mcwTtwXD3HtEYUZSs2
4qGt0zbbcGtyxQFVde3qo6dtDeMfbswhIu4UqsW++gYwoYJMBfDya+62/0skYP4n
CCGptwhBRtGlpbtNKwlwUuUEjKvPhXjmvSoSdsPCoBl8kcGWUHGpff6SYHX2Yxy8
t1hYYV1n0GjZAie0WiCbrTu91wI7ks+bi1N76t0aCjSyStjxYYv0D+yOBb6ufRfj
XIxb9GZNEh06IJmoAhzn12BY2ROkxEfQyNopq+6d4XnUAkz2xy6jk76/VDD0ut41
jQr+ZJ+hQKaS28UZaXz6kM2K2AGx4WArWrH5TYo0DvaQTYgnGl1wwBnTxBAPOOBx
Ra3rNr90pJ9CRNq7B/xracor+oeuT0pTDyAHxigF+cRxghL0OwgthGoTHxJzR3oA
KQ4UQ0I3hz9dZwENchQF9YT9PX1J3eGcnqupMwRuojpW4nuIgrNOug0LUBOh0X9v
wFpZR6vpQqXs4gSorkorTypN/IwVcwsHDECCPOYqQyDb8dY+VGh/PXrxmR05z4rh
dPA07YtKiX0Qu/saDy1z1OOQIZjHmkCzePTN6PwKI0yWn2r/jLK/VqIbQICDNTF3
1pIswWhfYiMQD0dK3CxgAQyMnUwZ1z7trmN64R580ncpAMS3YGvcUenB3QVMolQJ
79N7/MhOwoymeSxpGEcgLrVFjv8HIcKwRtXHmi0vrtryipsZoQM2KnpusCqQzNDU
pV7NFodGPWJUlS2vRd4JIVoJu+RiUiHxeqiCXSDH/Hg9CKUMl5mPp+RDC53IqcbV
upDgZA9nT9KrBK1b0/RRJhwJtn5qKAQ1uQATtGVnOKkQvdWKTJ4+2LLYs4SwynwZ
l+E6Gn0Kn1vwjmtf78eUmADzw2Q7fTtgU6AHgGGLitnbalgXiFe1d8ZFgL5AAZSq
icgNMvOI69cRUmdyVDNSbAUQYt+lxypTGh/9cvvvvWkNye/c/PR58tHc5D1fm9zF
gERRQYMrhnEYwq25Gpu9U+xWjNyZlsi2fLfIUOtk1bOZJ0/QZ9ryRg1FzzctIwu2
GiyScPpGS7aDfwIh6NzK5/vJNHw1TUdPh+m7e83RsTiwHdH+4s/+mHFe09QuT0dn
MYKVK3MVNIfrZ9EZEgAxx3ydc3ikLjNQAUuCH+sm96yNHZK0rGyO0mrlEgLUwtCK
axNuivYe/bI6JHamSyh+NTedlS9U2q7thM/tEkS8QlnVAveeZ3YbhEUhnHlHocU1
H+AI21x8c1z6CwEbrVZdvzQ+OQEeva7BDN4sqRN+FaakGt9nLeP2IjaPj4aA8OFJ
fmo2yCT/8/KjyymSDyJCH5NVh4TfZSMy/Y6XdR0f4cjo2EKgYesxqphKRH9nYXgB
kfI+6rTXo1SM58HmzqW9lsGSGij3xUwaohRxXpwg5qfW7GZgGX8V/qDcFHc9AFZ8
IiPTIsD0Hk6bYMBRhA5/EqwB9c28UjREPvZoEdDjF3eST1EcPkrhE0jHvwiK0lI7
DZ1zjgi14OV6lh+XTMpYWAa3K1bhd2RgF4sXOhiKsvJrAa8c6KwRU1fKVkFCc4qV
rMXXoY91/6icyh001n4Sy4TosOyFHM3r2XwRzFfmTlJCtig/X7mA3hexvwl2KaMY
01ZLzXFgiy19NU0QJUCWj05j6eUlAOdUrIMTTRoSXnCW1Jz7fXAGa+53y2TwAmzb
EhO4W3f77I9V0lz2qhT/DRVAFE35kCPekwQGfaOBcjhoAciREY7vCslZ8nV7xitU
vcs8CXiPbPCHeBORJscpCkigvIXD7An7FkrVKa+Tlsh4r9otXWwapB2HVnCZnNGO
YjZDSis32EuqF6658JQJZKPbjTPuTjBSHbfOnI45WTXVLestEF+hxD/J3S9J1GK1
R6veqTVIwdu06iZuC6WEUuI2KipadJj+HBCRp3NLH3wcopW3h60M6MrO0duqTzPV
3WPR6Qk59Q1e1XewpUdBh+ulkgKa7fys4atl9qFNLW5KMPEu+1eg+/K8YQ1OkpSk
Od/BiFYfevAUy6NuK/rTp79PIQ5K9oFgkpbfR1eYlVcmvu9kp4YM6kk3NkcPN+yt
scvhbKelwccjDc78lDW2NqXRCUsrXpkxQcATiUWfFkxu8/wz3c0Fv49W/py/31NC
EGrrKPEfTTtrUEB4WKokoFvZxmz5vHUB9bMVsx7hPDZV17TbKWPx+wBYp/pUoUvp
lc4qVK8qfZAUhEd7XKKYZEHRKVs39gPJotNRBwtyykISZxjMJMq9h7c/ZmrQz+dI
RbwAS2lGO4Pvg98/81A5BS006PgXajSY8Afwa0i1rG2LYkdFkynymUnk+ea5bH8V
UoR1V/vAEyq2OXv+trG6edcQNkwdiIO5Ec49A6HPNYQy2fL2QZDBqR2hwBZ+FKzs
j2LL3Hqr9r4R0Ts4vnWCd2qs7EqmXxbYr4VeWmXz+WabwVW2UD4ubRYBzzANVDaa
N05e5jZP7WznImIUzY18G3+kpBocNg9qDckQufga3WHgOv73sSXGWM/JGnD4v4no
6VEgLISqDN5yzzzJFTdnodRFUBkWZVVIwD7F1/KdWh2cdIWIQDgCGOEPca+K6kSz
XbsQ9bVwRFBD8P5Pq8+UIegMZ8fI165+rEzUV5AW//oKFfNC9O2GwVM6rGceBHEI
wzRhTufLmS5Y0LQDKtH+/imXS0kBIJeSMk/0Wudu0uYb/rgWx+BN7m8nsm3UpVe2
A/1YxDnkFmJPQCpl2aqg9yZmbh12drf1TY7DMpzE0pwtpxg7P+lEqTzei8ajV9vf
ky6jReXNbezJa4TRpXKLkpmgzcZXevRswHRKWXeQMKqB+Ggty3RRWZPjeoWK+XB2
I0z1EvhPPr+gfJc4vkbUY+bQxo2JNNjFOZDHX1HjDkVAuTq87C5XZtWiPSSH/RvB
QSxjPVrt4vzU1R7PEiOha21/AV5jrM3/Dk+MN2/AEPADpao/6EngjnFbB8TX77Oc
Dwz52tJ149MnmJjtZGpQfIsCr8E4Hc0eqDWWkTLqEs+J75ZfgQO695F0KUTQqoTg
7J9CwULb69CIMyfdrE7CtZBSfgJg9JbahZ2H7s8OHaXSM6g0E65rQ6/L1T1SOZRc
dROnVzWScVrYjjIO37LQE4h07Fb5/A6kZC1OOVa95mqFH+++V1aPXiLf/xoDTSHE
qZQe/CD04IyXM3ttJVlOverx1ywnm/PlOg03uavqAR2loUCRXOZwPVjVm6If8jtH
JeChMIN5eu+tHIEnDZgQK6N2xKxra9pZ7JLaM90x+OEaz07TfibrMWZQToJGDIvD
j+BjNAVd4kEjg7yVUYfFR8AdIQvzQJYAhn3LPBmd57v2/CkhRxQkiAca/AtH4Pre
d+R/1L+Xq6JJkx3ICfqDmG+Lu3NHadmP+WbfFrtEGxgoPjue0Sbwh2VYJV1quEJ6
sJr65iRG90zSOlyqRATVEfh24QkTp0GJVkwgFBbZJ7lXl8cEwXpK2V9Ym16vRfU5
3/LOnGGSh/+arDNsLBmvIN4A37TbWa+LoAowr6M/TFL6dHEueY0nNzszDFzWVC9x
3xGcMoprO+/IsHmkwhjQUZIzpMsu5zoMmI8bm+G+/6qIJWZojEqnVa38v37pr3SM
TmnFXSxz03Xj2iW1X4gsSXaFOLFVqvIt6lLbEoDYKTtOjdmMRgHecrIpIVYxeI9E
E7/ScMshPvWp1htvFLv7LH8Fq7xN4BmCxLr0yJeRjrJKXnQS9ly31MJhAFpBOjHS
k8tfwy0DWVa4j4LU7+vAnGVt44UUPBovfdwZ/0ClPgVkh6iKbpXsApHqsVrw2VwC
sDF5M7FEFx7PF0a+6UDUWA044v6tkrNbPYyI4yV5yF1bCkgNTv5AU/RGKe95VZZb
LTiM334UUWdPgxaZVWUS5BycGHhQECJH6GV4ilk6A5Jl25hCxhsnVezATR6sKbT7
E2ai67Ahion8i8+1CsFuL0RoCc0Q7oOqT0vqziNtwGbnbUyztGAKFtoHdYZZx78T
r+5CTv6FdtALFXGiotkt4j7Vp+RjGv7iXXDakpqkJmReQYNXj7GNRUrarHSvdYdu
zEHb7pWXLys8fq8oRZOLJNaE/rrBMz67gFUFiYP6iLHKdgJdkPBqqX4Q0ca3uDNo
MReGPwQ+AR+EeCtzREmE1Uldum611sQi6zzFjDzasOZm/PDUkEkNHrz2vWBw/vv4
7pOL0CxDbsOjwJFEGMacx0Q+zVqQyRk+A6MA8xzQbdEbtwmb8TpX9U+hWmrbhA6u
TjnxoroROCBSxRVgDTnavMEYBrfRPLSSuKuxpezSjTsDr6GU0jpaOhNHTMaU7GXy
uC8Xc/s+Zdm4P9cfvw5Eqk+sAJfMXNNbgeL8qrVNj0UB/qoyvveJxO13QAFEIhjW
oaSikmdhw0QvCokCmbe2VYdRBVnz5YZHlfxkxDWa3ExySyV/Z2VPmBKGGWP++xcX
8DblibLCZMwiFCqKWOcWuSEljLxqEV1KlQrwgMsPmwMtEPvOxJlevq0vGCWdzsZW
BTV+c99tHMb7QvzlwzSWLsFkFghZVe8oH7Xuv+q8WCS7NF7KC11G1sP9syR8R1cG
rdU9PoRH0tPJyw1b6QgnzObM8dLv258YBzSdWKnVxCvBKhzS6ogFwUFFUCPbQSe4
Kp2/e6g5nezzsmxf7LfsAZeK0q9c3zh96lDtQshQNuq0XS7+6CZzbLwcjvk2A/+5
uVvGzINMnhB7GpbNe2U8bvC7GimKVMLunltbrGPom/ltWNCYDSEodVwN8VOQpSrL
7rkUEQevfQpgowDWTmqKem150DLMe5+HB9p0bRmzMzHymb331C16cYcHYWWtHo63
3Wr7KFwxWzfnB8XI2Sy/NcT5Wpn1V3oiIbWepOwZiKBLSP5Xe5Xn9JW7UPCyQP5l
lZB7A2fgZIL/ajQouhL7uXVEcMuiDA6AGgPbiJbn0YUFyxi93Ns+DmsypmWaT3E1
9IsO0u8B7f88tuVulsvJd/v+KNyd3t5f5vW377zau7MGSWhgXkKRVja0lSd//ifG
6SCGUXOsUmqwziywfjsfURZ8AuUWVJ8I6/EEVFqSsRCjYPxkuwZ3zC37acP48tY3
JM8Df13XRRSwBkG4fCJ4fwTJ92IPFtmEWZ7H9EaId91InzDoSawgKG+ZgD6hvYq1
YvmzS/6iD+QF5Z1EWtl35BYUf5TkYgAvG3FUm/qm2IfqfQ4P4kfALtws+XHXc5qQ
UXoxeHBflHzud3hldMUIZihn23UnUyqHDQEeLRIdZJ72mx3eHdDdEUYoIsA7vW6C
QSnChH5RZeYgICUkPUF6ZHD0YmmHsXKP0Gji6MSF00NNoUaRQ+CPdvpsvDLasBh+
nBxa/1G0S9XcX+jkgQApQF9UktsKUrjhfLHV9YnzBqa6HK0F44tR3OybVTbDBGuF
vCFNU0nlPFOTTVbXBNcRACIL2wYMxhi8t0M+Xphms/zYn/KPe+i5b0O9gB6VeA9g
dzYXZuTL4OyhiSfWkMdPkR0Dwn5mm1+Fdph+tdqiwkf4Qpfs1hCfQ9+erZ7PRs+W
CaC9NxjX1wUQgefgSA+T9VxrS/QEzeOuiIPOtPDYXOgk9+sp1K2KvvOxm23F8YLy
AfNohmETmpn8k98DPlD9ITlc33qUxhux9sHmI6xq0kR1ZDENA0yF8Gltz9jotsba
YvcLpr7ChZ+Fpidb0ByChExmtFTepecwfuUY1VVbUo8KrScTHg0bOut7NE6WvtG5
rqzR83zBsYi3X0Bfn4g4NUXdmC6Slns0faMXps9GsEHv9ZXdI8VkU6djXk8DAF9L
T5PLgDxqRC+0pb9RAx4QIiQD/JKjFZhjcW+gjkSiYLxjuY8HNpoqph3Q4hHynb4C
4qXbM9OT4Ff60UQH8/pN+LpMvJoF59gyEFBdhMurO+JZEULnEc19B806O4J/dzw6
ZgFi8SZb+V74FxGpmbXlUgDipAgXu9hCjPUKqW33TjCgecxIgbsKi/t2S20pQTwy
VImfI4a7/WFWXjHyZeKA/ZW9YN4fRByx6ldm0yLhcYDPAI1rNfCK0XwqhaMgxCnm
STloApsPykzmbHDRdATTPlPzlRqrfqRLoBG5MgfYHKV3BHgM1nTVWsdIwrBS1/D/
vfVGMPL/117A9vH+RqYQLzmEWSgqmRtSb0V8HHWtOyDppbq8HQkhHo0CwTF8nGbC
hUnCRQS3Ds3i8Btugk9VPqAgouJecV+lNTVzkwcWRClXn346LF14cP+7UWgaim94
ijtlo+4QBIMYkcTW7Y1jWWmSDtDfYW35avqxYt+LQ3sv7n/N3P/kGMYrNPHdotTL
7o4S8kUWp0L41PNiubpGGVyRa03UVksWYRc5HnTxpQ4ChaaHOH5QXrZ2kw0ogHsc
9/33vHalbDO8MBUZDmdPk8inrLWTa0xetA+dOcRxTnqw8HYsFhTTOzLRf6l+uK56
k77H/LlYfWgSUZHlbBsckm08Dg9KpO0yVABhRadx5qYdGUQm9eL3utPoeLVtd1re
NinCSbK2wHtybClgnWjrUcWWZ4JxDKBVFlJCZfxjUGPL7MAiC+a5XLX/e/v2ameu
emCRSOeljGdWJjeszq9+7jvP1DNiNFmkMX1GjRXC6cS+selKOygOm6DMuSiZz/jt
zsngrs8DYP3rPYJYiJJ5RiZ1y7GQkq3QsNxKua3YOix0PxFx5an/IScbRcx+KoEg
3XlMZtuyt3ja79gqAFsKS7jEoAtiEUmB2t9EQ+NkQBo0IkfGBF/92z1XWPeD48dm
zX3yz85NNgIz9OOjjm2E+dmYg/UB8lVhwuY6/bleuPvIuBFIPQHlwuLUoOGMIVj3
2q27VZn6hi3v9IKkc2A0NT26JJJFc2g0P+WSHCDJcv1bYYdx8Fpyw4Yy3ug50SeG
iIOFBTEs2R8BA31USdHpk4lVtuglZMV1YBFHBQqfo4KfGvSxIRnSurSzgTaVcQ/n
OEPJmDrsZvnbfT53lWU0WMa0tkoSyWtJPXXpItEdRrj/T2BFO7cyqsmqbIYsV2/k
B+K0L74yrHIJGpI4bRJR+ObxGPxH1l45OID2SexQIVgAh8rEgn6gDDjE1hlR3M+r
Stf+dH3zwcqhMSZd+3chItnm5Mk7ECdlqN2e0LD1/eXGMIYOLTdGvgCLtRq7zCc5
QgjT+V2MvoNJkO2Ahtk+JDncEK/dTck3JtnOnrgOcPUbDAdw+yWC0J7t+IbmQKzd
xs6nmyWGZG94O+A1oDVKdRyz5/a2694c+beMwjw+kkgAHPVbvx4Xxnh3G7pIRAia
afCkG8EX3EmcZapboQMlSyQqSK7YReyfuFBeFkeF+F1mlAa5gRxjxBO9pim8SMN/
R5uPPKZGvTG9xhBF9YOrMoax4djP3tgcSJP1Xs/qaSuoSN6tnabUQsom53vdefK2
Q7snVlaqEf+C+bQ7Xe83rCF0D9RFaemcSuSXu7odZzxFewHrIH78euwYNnx13Cfm
l1T0yaEPYO6CxXqbIAWmgTkN/q/X693IegF+uZyC/f+794s7Vrc8m+DnJVZ24961
U7Qt74gvlHyKRgw7xNpY2hmbO6DgILhXOke2rY04Uyx8r4ixsdCalF/6w5KDHOGx
b2xWNGw011oEb5buIcyi+hZ3L9D65wqiOhxI2xNu+z0++j1PQ4u+lE9M11hiL2Ol
0i3boajqVNvShmnDnLi/A70cuBYjOkFMm6+oPRSIKYI+bqjHrQwCdUc0MKe3vgry
JdLI9cvH+ub9Y/SA8iWjB3ZMAr188DB++K8QopWliVnVeVgEPntjZsHsINEe7vAX
ayhuhH7UICaO3qFdAKN+qI6eoxvtgC196a7dw50NuZaR7RDScNmcSg9qeKBMlU85
0MH4JBVKCtZCHfQ7azCGho9DVdbp6QPjHoBudizDQIXy7qetOZeuSoIZXLGYU44G
mk+A/SgL5oZb5Lu9He08t8bc1Qg+cTcv+UJlHr242Vfc2NZkF99/Ii9oRk/JkWP1
lIFOqTRquDRMdgBQ7Jgy3cmRwJnsNtHhgEVdUmIi+3xbGi27yn6v6HAwxJ3fNYp3
+iMJE9FQlbw89a+VIr/hVt+cjsG6MBiLwVJjj3gZ8Pkjir0rA4GkaSduf3ueVAJz
E9J6U6fOTQUyDqlzzyv1oiDJZaiE1uK/ByVS6enjMcDyjD5RK3zPz1YC1dpE4snb
z8kxG6mqbHkGNnSIt3tOnxQzcaY8Rhgjbh7ooOyaXc3pZZjP4S54EJSg/2JZoPKm
3pWZRBrl3pd6NynjdUIqkz7IVYOLjicHiTK/oWzQHZWl8YOdt2ybZuqARyR8CUUs
pEkkm6g3TFMJV3r0vC5LakP4szu/7LMu3LJJqJMRGGNZGPL1jdd17r1qx+OCYW+x
E5oThFS/zo+TTd50WCw5l6YG9IsBBWhwio+tnlt1VxjdKprDMnG0lvYA6iqWHKgC
onGCe1XhxDL7A8rbww1IVLyEBO5JpjVn4he6HgeRvkepydwwCVh2TXj5+fPIlN77
YtwHwhaOc8580UDsJ6TPuWn/4aekmWEIPELfs8AO5kGUUYPKze42+PXycrOJpJxR
TGaLuYlg1WmHbmRdC0vDuApMGZW6z1TvEkatawIzWrSl7vSvAVeluNl5lxS/tUrN
cS9AkJzNHwUwfkeH/VTvcXV+QPXBB+ht5vnyHQuPZk0ctI61VC5iVd1ZjWGL6Pzk
VbJA3XbqfIS5aUJTohZUyvue5UI1Gx5LI8bxlPZ9rf3FGJCVlHpTZ6v3IIPNXbXj
Ftc/JxJz3JpnPcxNgMlCoA83XQOdWdsw43V5IVIoygFK2cdechEtg1xPQFMiqqqv
uBKDeBFk0qgNcHLdpiduMxsywaCpbJm8ItrdNYDd3V/khMXRhGnNNH1ejvDSNmax
dDZK17zybVSo9kbnjkm7x+7VWOqE7Y6rca4Eu5oTm8tkQ6Zv5YIYNZyD8209ixNm
VUL/pIaPNFJpqGhZlMIOJZwfo9C2rutCT/ZeR7ajMhLP8Y7TX5pNFiSS1mAh75t8
UuBqbu6pak+u0P5bEhWrHzZ9u5Ttqlz6Im+EjQmAlpJJoY4NfU7quAnAo+1MsbKT
2O0ukboHVmJkadnYNv0QUqUCY2WKjS0kuT1TGtFytkNDrbEOd3LW6OElFMu8SJjk
VPph8QuOiNgtZ0BlvDsQGjgWmAx+pBLPZhmJtEBI6K8MdXzo0fVdxZu6lvDJT19m
Z55aLLtTxe4Pc4kEVpwIyyZyR4hsOYI79WH7n08D0EBH9b0ivh+U8wVr677x51Zk
PvTYfx8z3Pma97io90KfQUcoydu65BpzA+77+08vgyc3CYtZuHrcEGCbVIA6WOLE
j6YK3QoUmpfyL22IGefRXEH0ycZtdz68bWkagEwRRdtnURfWKYa3DNOQhQ+1sHFg
Hv9xiWBmK/qb3HPQgbRnsX9/VhmBxkswpMqGYuiFvBpiFmHzdMfe2zleLXHIEM4O
YJtxr+Ec/ES9oWB77gZVctBnHIwSpL1DP66nJXmf2fQTYEoTFadVLjCWtBwGmfpp
hFvcCgUdp2qstXWdeedIY1FSck9h2KrZvhrVNVq6+hhQYqZtLljgfgROYmUUGuZ1
MMjpfYjDZ1b31gZb9zX6OSs2jL18RN8KdI4HZcadr+Ol/d39FIeMi4KDjQ6SFMdf
kAvzB2dvyYcIxqpDguDhTCxILutSl2ctr14XzPRKmzQpNawDh7riXoJcOMCyCG55
r+d/NzFIpEzfeU7JfeZxx5BwHh1Sz+Djmhi5U1nVpgKceNM7Sen3UXCBoGbMMj6S
wGQy9fMkdSPOJz8RSKBpMm8fxyrAqKtC/z8ZR24cQneA3HEHMdk2Rzt9aUc1rmIy
9K7WpXLk0stSwI4K+hFYKvBVDxIMbEGAPEPsOUvVBp3W0ljGXp+UiEv6V+ZFWWpA
9qgLvJUSCNItk7ucI8wittcfTifK5VBDoD4/k2eokH0m61PPqwuT7SQqevzmM9pk
exNZWwHm0J5uvCcUFEDapWJC8BijznyrdUPw4Lg1YSrcc0vaST4tQaDX8wBxP/LU
qn8W/l4rqhN9YG6Mcnh30VxOriVVUp0CrwJZk4YJdTOwXpFwiqH+szrh/6mtQR0A
0fFzhjjiiCbySTmBzJVn/LagAXOESddDNN3ZB0GAn165ooWEXZHBNv8/bCT31noJ
cTuJvDNjbwRGcsVAOSOD8y8zf91zNK6Jo0T7kT9Uwjd6fMSUsWlsUX5nz66vjHbt
oksoQ1Sy7twXJCkV6QkI34Zh91PTIAmjhPn2nmX5UaMlr3I8cxV3FhNFzS06UA13
8t5J4qjDfq8n5VO7PiU7DQRJJi6icDq6sbnt2ueeQdVZ01tc+TOdwNwnzIWcoGiQ
VNlMtGdq7biCSI/QbMJNzPXBag8z1B0ivCSoV6bseVhIXxqkRy5TfCbpnFKS1CrG
k4KFlpXKSEyskBZGzDVHbii8PtyBT362h2Y6wa64c+68XWTHivoy2LRlYnbG1CU5
Ph1inkA3uCtmSBaEoWYovFUzWys9dU7cg5JaXiYyoy//opK8iyyt/DcdUXMGJ9h0
CGYzfFbDQVD+vuYgL6TJddU/vliPLVqj60jUAXNEhVMkOOBKrZV6ixyM+Zyql5Se
q149WaPYDp/nVMFnCaW5QsXjKEuP71PtUEEMwA5++Bj/x2sBx+oGu3Ck7lAcAugt
UVBcJYHzT/MRbD6XdYiYl1fNY9Xe/Dy9xcohxld4pbgnHMkSzWk6Khz1b6WHBcuQ
FGMxpyTgaklpSTMKbO4aIvYZlAy5GYVZCD3ByBk6rPo=
--pragma protect end_data_block
--pragma protect digest_block
MEwKDRlEk9t3CxFpp2V/e6Nj4gE=
--pragma protect end_digest_block
--pragma protect end_protected
