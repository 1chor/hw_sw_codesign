-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
lMFWmdweaJT+E23dtjTdMQ3be7BQIArZrVht09PVBv1fAdPX+FSFacDakhLHNJUF
WYaEM13u15AxrAmZ684rGv2tdtT7AM5XhbXO+r+JzUhnw+HtfsTH7qakgUyrhDjL
xyjin5RU8nmiY1DKx25aqhd4ONqCe35p85omUFT/rsM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9536)
`protect data_block
sqMm+jNVdnQX6z/qADkkGdjgDidAKtPKOlCGoqqAoXBKWCaoDTsUkP9v1+YmZ+iG
XtUAaVsOG2fW7mSx935NCfCn/gCGs79nEtypU9UyiPr26lRqq8JCLU+KhUW+kf+u
jIIK5nFkqmG4+E4xm2Q9cleI97AD0ZaEX1xFGrXX63+gDhNBA6KjqBezwrdtLnZ3
LmqhEJrltYquK0wJpELfvajfRpIu5Ik0cqRhEaaq1kOKEX4lJy8uPjFOA2U/Rh7y
Fx/TZ0ngmfDcrQ1ODeYEWoamxBdrMmh1pX1Km004qhnpSAEKPyBzsUYEws88Wc6j
d2UypokMPHXJktnsEAxeeQkPg1opiDwyk/47KBYYVHouJUzYiGO4qyrIpL5I/7Fr
IVdgZHgaLhq4y/cWSoflxx5uNCfwfKAO1CF/24WvBPo9t6VhL+IBUhDnwNKOz3pz
CJhy9+josuGRNRTpU9lk1fzzLwlMBg63N9pZXTCxsYJsBAbDC2/jKS36I4Rg9Jye
uEt5Z1bbqqf0UEM+d47ERBbQHl2W0cfDbTWpfbKd8oYGaP+IfW+hOLkCM89JCbcF
zffyv93R6wZGg4qP53nzE3VaegLYg7aFotlUAwWP84W3pS6G/5VtY1ZOmBqcYwd0
psXZLRGCbhnhC1m//ZJHrGrwELsrgLxCYBSyJVZjkrJnwfDwVnh/daIbBfm3kLuR
bp958YMAKehYcTdPItWuG9sfUXkM/jOA+nfpJhkOMXBYitNbYImXzVwvSfyyrAaH
/Cxnna21WS7qARPwLftxlw4eNLIMooyU+1lgLxgkhCf2NapTGc1bE1rp8FUMn+I+
g3OWQkCOdHqHK4Eoktc8uBqHvDXJZ7nfPbkYrXxhGG56SWOX8eteQs+kOvOWyzLD
ghrNDXBNtMSuxIfmnJFUxxQZamoBqwlNcy7CQe/LNO6QEhzE8o/4XHpQuCpy8MS3
D4d+GmphcgjDZCj0U6+wkYSk5kDT+HIi93idti1xZkvQq5mEPdMwrJKrUiXl2ncd
syF56BMsnHhZeGusOz3MurPgH1oUU2Ae3dzK+V2+npNn0hgrgin3HetpGQKu5Q0C
zOQpH1QGvjcmjje2U7NDGQR4kUbY14Qzy6HUCXTm2o/fa54J18rix8TphU92prEl
WKGSQR4OC3QzFpZ8wfgqtwI/4r0Gtm8eoAouZz669xaRIC5Q80wIo4+P7ZKw116X
7Y663FREp1CbmTW9D9spJkbMpGtIkEh9yy7gS7j9vdxnXQFxBAxO5S9poDV92W4v
D9JOXm1wUqVW1nBRw6YDn0rmZl5bJPOxa8wM2e0usoY5AwY23K+a0MjqYvk62fPk
tjwjPC7sVij9MFfpBTqsqpbOUK5wnZnZ+9/aC/WHNYWtuTOinPD2ome5636n2xpW
WaocWxfL3KgPr8x06mAzhhGJMfEwqWlqok/SoR6wlXWRO5nhxYFqqI3PwHCfdaZK
xDpk2t3hrqZTjdW/FdrDwY06DW3U1f5Jm9I4+PlnbNLRoJuuytUIDbRqUsisxBt3
yR5cb6g52OiE49EbSj5gdpMkQUJXgiIZojhNmDI8bp8hf5uOsBhYIo4dnkGom9Ao
c6VqjYf2KwTIwgludDb9csfLDcafmTA63kcOiQ7Pu+VX3gvulTlN/o80XlkcGnen
oW2R7h1DvlHG7UWSiixlWXdDxjOYAlFB1cTcG0fwMBt6Ztq5jcMBAcriaMJWtARX
EKpO+zTKC503opkJQjBKnW87wnbc50KGUwE9HgY/72h2tG/ds6t6yH4KWbBdqLCy
EaOgqTvlA3X1Z+cUARWa+kAk9DSYRXqILT0pGSgdSFegl/Pj8POb/OCKkaWZ/2cQ
CRvz72/xUB9otJV18DHczkSKye6Yt5mgxDK17bV0Q5ZldN0fYVpEJPn81qP42ARE
3T3G5HDhbZ2vq5fe+wtU80Y+ViSsHrA85n5iYsJbcKmHFCv8hDBwI+0u7bgdtRY8
s+6hAoGvUe9X8Va4PcV8o3aciMYaQ0j/4yxgF0PqGbwTnDZ0qO35s8ZRPuDaBCD2
gJf2HwMpuDfTaECM/p2n0hhk9h0q2t+IVJLsAy230+t4UPyyuKMOFpowdI22ua34
aYay9FVnTOMYlHoHZuY5C+Ao7rFrasZ6NjPt+0NJ9h1/t124vobld67ZQyyV4qrl
/qJ7Fac6Rk3VRB4F54X+q2gmEK49npDElmB4W1qRqXsHdw2Q+YngUCT6Q4oZxcET
/KVWTTIBfajWhGqfTfxTeNSoc5I1ZDm/O/LFdrEE/KUQwhmoxiHMimm/XK8ktxKo
4UmjTzRLXFE4kbiGvaeJbGxFH4TOt2aiGCHt06v1MtQm/AS5skLHFhdKsWpukXaR
3IDvOFT5OYyKXKzdc21CEHKpDGfGOmMYbdvC1ZMH3s9QKuHlneFBuNCYvTme3tVp
5eJ5HeabUQXFhbiAc9oj4fnfiOIYO0un9B96qCEE/XCOGSqeThM2AXUXB6/RrPl5
vo9Eyl28f8ZEEdyqyv6P827Yxzvau8VziUZML1nZzwfo9W7gkQpt8cZ2z8qStPVn
REDWOy4KsP5DfEUnP+zM8tMCYd2JGUCwcldVzdV58v0zrNUuS1IYB7QIZL+PsyzI
q3cYHQPWIUFHHOxETZm1wkR6zvC+ZSVUhrcjo0FGuMcM/8KJmrl8To/2uQyMVyUf
JVK2qOQdRF6MrE7DJwvttJfM9+yT7A1vII3v+uN9NtW+VyE1nLzIxAOYV8dhVQk4
m4S/dVjdnJ8iZsI3ggkYyd9+F664+4vDexZ7weFmyBeMZIaYWZ1oOeEwzWyYsFRV
0vm3KbKxQ9x1PeZaPtWUVEkRBmyqKHO5MQOrSuCSLkROXps+V3vGd+gg96Kqi2g7
MYjpDm8QJFXft5l5Vel7bSVnktddFeleGmg1FpTD8rZGTOgVJFa7v9y5vwSlE35c
DIy835wVfeNy/l2+nmVM8YOvKOjIYqa5zbL2Zy6LAYogQrWcReRz9vfBz4tu5r6w
tvuA1qbI92QGXPv6hbxjRMAsvc+7OlNAcGoeUj3X2WB2WFF9NnHyqZM1yJVH2xuq
MGfNYqrp4f16gko8lBy0HaQ4wAwPrgndXJloleZr4YTymtgZgAT1aSu5I8bciBhs
cXZl0msbeA35Lxr6YW3XCpZozstC4LBHognxDJQ5GzI7cPmrPWhZw8+YOoUrKynk
f2nPlCMte4BqRtt+g/5BAPp41ghn4wHh629/U3yfdKZgUsIdXJh1Zs4efcG8XxG3
qU1CVTh+8g8ZdFzPPuJVDa2b7dO9AxB0TkGfiBnunUOHrP5m+OYSivQAvXF+IKKN
y3kFKN1thL/pT90O06k877fnluSBSiCc0DI87YyES9MvA0y+zKGj+GReLLLjw/Vm
EvCOZ5G/qTnNlK7QwGQ4SvFPqpNVHC72htGoNQB+OmNjdQAARP82mRl2rN2vryEF
Ix+FxQdLeGYzCK6Rwrn/6sAIegNP12+HFrvL9jQu3qpEPE86gtFz20nddcP7Ckei
C4jKIBEs9dt4JG1pa+VQ+66pPX7sgIhdl+5juMOE2KPTlzfVS7Yn0Z4h+k2rUqBO
h+rOnuzxCPLSMqXvtBrYX9sNHcZ88MpRBhK6XQtNL7grXV0H9CsR0xfuLqDqVkV5
VVKagy1uwDmKSdFuwI/5XVb02GvZggokp3ZJZZAzwVeTSwI9kUgqIWTRPYXgo/U5
OJ+1oMIIE1rXaygj6uPW3nuR4m0wnCRSy1QU+2kVynGy8P1RdaBTK/dIJQymVxTS
TQeWYGx3iFL9+d3oCYEfZWnXCtXkTGPhq9IOpaezKGgDbfegqz7/ExLV4B/dKQqf
tYHxMEAgCs/z/d3Eo80AIuZMi/L5AipPGl5cwjYl4upSlsyWiFjG4G3VGJiRNsBw
G/Xe9WP38mMekgbfzvPctBh1ZA7wu7fBhB2i3ExY9cKqP8o7jDcTUZvJQRzj6XRy
f/m/GaNQrAfUQSoyYNQ6ftHJ5YS65oqZr6/WVgLxL28SVwsIv9JeXK6ppUvJbSiW
1Ul2gRZoX8h182TvsJzitt7x8hYT/nrFj87/EMYP9suoOhbuvMUeghKT5gHks7rP
MzjxnUBSOsdywYkaWr8z2pbKtXp/tEX7e39Dq6z9USzJTgXImRSooKzx/IyFLt0y
RAqSe3+9KgWAKiJz0q+3Vkc2GZGjULWkjUOfFMjm2ikgoyP8GqnGTVKLwoSygyl1
uaiUooEfKQpmB04sx0b0cdg/eURHsqYrXtG15gyG1L5l8cR6hX7t7Px1Lf+neBgu
bPns3bbSlg7hNFih85IZB8wttiQq76r8v5motX9XtFLlCFsYZBC0sYd36h/u49ff
CZbpMfVqkrMV68Uz4z3SdK/OGmesSnD9ZJYySq6NR8D8sI8IBdrl6VYfr0kA59gQ
YmWShlayq623x8Uqo4tGCH+BqyGiaFpj6nDpRborX8LICMhCYVRzFCAtU4i+Rqyz
FjP6pjg70tKLL2Pwa4vrafAsWgOQcRoUWKPEWL/LDhqDfAkWi6DiH2vC3KnnKl0i
/Q5C5AzIEtb/p0GuO+UvLWnPkkvOrKj7jp06b5VZKjEYPcijV2JhrAXMu6szyhAn
y3QUBb9GAWvCIaDsHvodGx5ebkNn3S3QzZdgDZKHAYlkR1yBCLSWeg91kbasScHP
mXDa9eV/UKzkDN3l+Rm1wpg4Xo+vnBUH8Q4R3VPHAKPdl4EcFAdpuzkXtEbAUGOv
KYz+nksFArU8BZFY1CNy+w2zVEcji9eK0Gq7S3E8/j6JSip9XY3x2El/T2puWBUM
5323vbWvXp7GQWRuYruGNxWWaAwIJsNZBweCNlj9c3eVanBS7VybWbavvmVxdPDe
5tEPs9k791y5ouD5l6CgpildJgPhhQ3wTo1wpEf+wpsa5szxyigNmpIwb7X5P8tJ
s1xhrd68Miwoqpqj9JLav1up9Z8kj4ICPQ6cFSRJwrfjBu06fZksnF3xYCebjSSH
tJvXyVWw6l67qxLAbBwoeYnqBElnc1D0rytShP8dtoiEWRPpsWkiGioEwArLO8My
Hywu7sCk1iMnCrX7481eSBJmd9qbO8iZJEWx4+ZX99GBxg/Kaw28krF9mTyVv06T
HmGmv6finpidGtrMh/YDvbQ1Q6pt6Q2XtE2b/AYdVjD4zveE+xDV0vI8KlRy0Co8
XcSXwK+neCaUU8rYhLgJxMSEhAHXWVkQV0Q17mZQtuIPzyN+jClPAPZgG2XcPjM2
Ew8zfVZn+KX9JTV/j79RWHBYLA5flqD4G6lM1aPj8jAV42Stef+E9PYQo0xFLO7l
sTcIUd7PlxEeSERGMLAXkQD8DNLm54JlT53/Ixl7pScvM3cJ0xrAYGIlNloiMYp7
FxeAgA0PadhNwvnDdFR3MZhj4G2VmUOHzkTRenYyVE9+NQZFc3SQaw1ofCEF52Gx
HhldTunzdnKsjpBEjBhicobrdmcdTn0xlCOEyOg0Rk1kZtdVXy9L3RvNozAuSFV5
GbZ7uEEL7pDMLX//vr4svbDbDG6crW3MG4gX64s/6GC8lJjDJhyodVBBLmbqX8E+
zK73YoHb2179iQufaldJIQ0G3rQpJaTtvnUiOFEwzXFkodUE4MPo6XhHL9KgFtaG
ym8SYvfBvvPqFzvc/siYIMoSSDa9V69aQIbyEj3bQ7tz2lwzQBIQ9HqydzTgzhy1
F0GCC3i5m91awJwo0gcrv7f6jK5XsWGcLztK+TZhWssZKSmPXwV26rXKK6ongg4a
hUIoSaS8G7ndeUNxNLU1oEkLiaBuYa675oCtIG7EAYUbPElnAzX8ZEx+Z+Nn6iov
an+oCU4x9aw/+fVGjy2vWXvpXP0KjOEKB0FOwQYfAbSeP+TKa+E6X/3/GklX8a4K
wlu9LCvxgnLc38qBiH75Jw/nZ+6krrIrBfLwlhQejlPHA9W2Zlg704l6koIqhIGz
jrP1emp+AE0NrYTHh7d7O9hi4QUnptqAiiy2pUwVv5nUfpo3z7/lqwJzCW3MQs8l
MUIIvCpmMjuDniWwc/5d2sf8LF9f7CsOoJmVyssw5iaOlH0oDJi+47f1mvHsM/nD
s57FRjol8NsDHSp8Lla46afMZ48bBwixz+ebGZAvFQHx5bsZmfyx4Ij+jao+xvzA
TGlE9rvvZNKHX8dMSAFK9QaZ/ak3StIKZ1U9G1WlDAHpZX6BqK/1x812RU8B5yKV
e7gj+/HjQWjL3uvlT3tJqERCrSm8IoPITaXFiv9LKwnU9p2NHrAinF2Dprd3V6Ry
7wTLAKm2oIE5+lht0elSKePW3mfwVY5dYX4yR+krkxC1q2iIQmhFOCmC5rqsUdK0
LSU7rKTCkKMLB0UFSou0jJqE796PN9kMNfC2nRNaEq/+CZ+djAonXyIDLh+aCoaw
Bdcja3rdSrYtTvrBBQ4ngdhL9Qdm4HWuH782sU6coZU30I2XF4OawblFI8tOu690
lRW3RdDKiBWBhCuY8ipVV2zemSNqp9xiNTd39bvpRYejIvpCrqACrrJL/SyHD7L3
pS9R7Z167zTAvOUkuTI/23tuOANDWbgVb36e+AB+z6Y0KevXZzrR1zLnb913+MsE
y7HlTHs2tQjr0wlL+MWSYsaBvY0dYRFDsTozF81pN8Ow+MgGBonRPk6+Ya1I1K7x
raXbcrEGhVJmJ8qvaCKsJkhEcy019YmacIMdPd5OuAfrEOgvgwj2C34ynNJdFLjo
9kN11X5qozOH/+Wmrjc4DAl3LFWlDcQZ6AlseZBHbIRJnjUtEgymjLzMjhJk2K5k
wA6iQVoDAgX+uAH8HvA99k8/AY3L4n5PTw8uibwrc1gxdIXaGWlVVTvgw18LN8Wn
YGw/z5CwtNub7SN5dnxG1v0cIqNtPlmy18RKEGO7jR7hacMVjP09VUdxsCsnQCN1
/OJUDSIbhkFNE+XLYv9AWnXHYZ6D4spsisnF5P+453L9wUqGWpESITkrAoqwayNH
+Ol2xFB70V/YTssZCc8lxeTUvZhnYzq1PAFSxWguHTQn5P/u6+GlA9SCQ4QiXAeD
xcQX9xioxSL551l3X1yDN6NwszbddOYTOV83zBnYEQmMo0etV59pmqt+ry66H9Jz
N21hwIoNGemV6Ydv03TdDmsc6+npnQI58KJ1SJPKD1c9YGq41orkGmvf5lGSflhU
NH8L2Xz7Q914tj1sV1RXsbUxoASmKHq10v9l7+3xj2TKYzSre85NXhFHgPg83+RP
8tjOP/XpGdUG1W2WoKEVQ/MDxPYJ1Dv8JLLcNjo4UR1hopsW5CPkIoE6BpXWxCLh
kCJDpZ0cKiz73I3fIJi2meRHPWQuvVAk7CNWCjfivvL/2zKS4j6bB37CdUbya+BF
zhe+uTFYszRTeRaG03/VJ7N7J8zIvTbHV/GHCOuNASj8hzW23N/f5gDMnGLcohAk
AJsMydqWaczICeYIV93g99v0Ebe6ON0nvNRWdF4gSNf7yhNmB4x96X8OEq+oCoLx
7haREvks0sgLUQidr8nfffXEB5Hr/61FcIPFX2NuMhCsgW2OiIC691aUZd5ZCuSn
XrBJvTEuq8E3UFaMQBbesuJiS4zYJ1f4IbYLmtmlr0lyma85AUs3qhGfm0FlHZ9n
ckFZv37bxvWFosQEV0ItrGYHUOSxHPGjRdBvz2g/gbie+ZoPhIbm8TYzMVcUYCxz
ermH5jiEG4GuE/fP9EXCtWBETKDTaw+rGD4TlQD6b2eAkDee4kvxckNYHFGq4YId
Jvk8vWufoGY2vNE+yaO0sy2zbLZDZFaslI9Kz8WVEg93+HkjiHdqCDHlJg9KsVUE
u/LJHpcUlAKxBQvGtYPb4Ux7mNVCu/6ScxIZ3mw9K9XbYxu5NcpXmaPPj6HNztwR
CVLpIkP0hXwcG50KNt0bJ4kLNlxu1pwr57t8L9iBLYfiOqevQRV1S3rWzQaAOmk8
mQjC+T16YEO1l24m5KmgJIwyz6P3BULtmAjm0sS/WB+2pNByNAGTO/3pJf4T0qbt
Wbugu4PRZi8/2KkUoMa3A/Fk0+kFbQ31m6Ahl1P9hp1m2Z/Pj4pMqrDmACCt32wl
j65otL7fosIXX5MaoOW/wLPx59pfmMc9/SwWlN9y++U9Pf4H/8ZEk6C8N+gyFRe5
yMvtE4VkDWw6L27+aM/ytfYwmX9XZlWaHONbDPvHathJRz896zJejfAbPRn0Z/23
L2Y/GtmAlfIL0FNMztxS9UuF9Vr6X7gzaRd7PzVOaqhGKftlOASdMW1RKPiQjgRM
xVgsez4oMgv+wjjfkMsnfS107cb0HH/rtIMvnVzajqqNyIkyntB0s8tdKA+O1HU6
RegDIgqpRhkpVTmp9LgLN66CmBbrow7dZ/i+xKU7z14pXsK9X8dDa3HYC7VVKA47
u2L5gSDoRnGHZjdvgV62lHr6TsoD67Qc5gv5iGrh1d8zpR/dhHnD7bqEtOdJ6fAY
fSdK55MtzFU/MZadNJP7kbJu0SP+CwKnzRqjJIGgrPhbD7SfqlBVKNaDHMP++h1l
ORKPD0FcqYudumOvEvQ7N+2ZcRn40WsNo3CPPPUaYltbenuJfZ+sDGGKHRjn65RR
vweh+YIUKM/Tft6pj8ev51XyHpFXuDtNv/iQW6qWsTsF6lWY4AeGUIwuJxe25RX4
GosD2ogZepjwXGY+32wbMEPP5oaCNMovi1kXhCgp2r2Zz71EA3JTU7YRp3M11rYx
01H3teIqgWfXmXjy77MFMPzDa0A++DPKk5j9yArJ+vnvFjWFXsURb1l8JlRWksnD
d5XaHJ7K1m2Ngb6ypKE4DeXNOO0saniCOSJdVHpjoYiofeTNCxLNLClN6iiwlJ+D
HUtVFYAZ3AULT7aDMAFA4GSKGBg9P7ko7uJbl2eSEGj+4k6PpUiMFhBI6pUwTfOS
wihE8BUinJVy2Ux9MPZJzoCWTT1ofMPO49G/RGd9aWyBEVsaXy+95IklKYqT+hcG
jNeF27GAkeFYoHUUJF5OgWW8zXEejbyq3JYaLE/3zanmueOBVVduHH8Rltz+/bRe
8v3HDEcf3wK2KeQpTjysZZfrxohSV66naOW9Zre3fTUVyexGhjd/P+4IJc1MeJx2
6db4JNoA60q8+k7a/jJuafl0D2fsOjZXS5JSxyiio1CEIlCLSOxDoioi/zqOTHCS
UnCsu6NCBFzP1W94j+E4zG6yrDPyZue6L6hMqvFiyRFx+FpLgOTdRj2u/PL1dFh/
6JfFyxHT/n1Kh+pSBRr5ZKZlCkr2qyansFSrZTLFx1Ap8dboBDL3yAUitn2vp66d
hDQwhhxm2Jv8ICUlzQmVga9skdfK2K3z9nv+fJcLdUJjVx7Hyy98LmKmleIerLHL
Cf0rRPGf99IdkmQXRfLtE7zsUTazwcbPsKoGTrzvHG/PwKPphbnmW9w6nQQpI/hS
CYZvnwNeo9PJuT2dB2smXiqB5D7AcQTqjletLDuLRHs0JYYBCiTkqhxpPDS9lzd9
CYzDlLJQBH3wye4dZ9WwAu/gyBEwCS1DBIQ65V5wfxvmjKAZEf/jza7ggjw85VZI
Trn6buO60kqgroI4fT02GWjE6xG6c6DqhcqmuSO6B7p7a4IXk6d87XMDwrl5XvmA
fDxJNeq5Ta9FFUUihknc142uBUNtj65RdzYjVYrw2OG8gGKPjAC5nyW8GWxeVq5r
K05HRmXa+aBSZjDcz7Fl0WvoeKiPpETDkelUPKy5e0u5tWYwoxWI9prtLkHkjwye
7+Ij7opUU9XTPcR5vd5SH5cnjiDb9wvc7GhDgVR4QODoDSkc1KJLaXW7+Kh5YHs1
9AzHUKz+1vqfDTnRR0qJq1sJgu+qMsm1dMztHj2O0/RDL4epGePCUo1btmACK0zQ
5Zdd+5M1BnXd8hb9XftlrVQgEq7qRwbCBqY2uFolfKHHHT3jkP3T7XPUkxR6gYn8
eyB7SxWUPD09dXjSnFVnr2jO+InHwp1SK0HJJfcX9gCUV+h0+qbn78hDWUPX5P4K
rN9QGUrx2GjTLK9LxQHEcS5P0GxMRrVSv8iRICgdSsM78nRipqS8vb+qmi0t7ZFj
8dJwIa9ixWZoVo8PYBHtPG+ja46VVtWRZ8hQL96/sF8yJAV4Uu1seh4mMMj9/frY
Cbg97yDMchENSnJ1xcnPHiqutC0/cSwsTXXhZO00hS6KxffTh2S2eL5fdANFMjNO
FNqlcZAfxZRny64zBvG3foo08cfM0zc+Fq1weFd1V52mfXjyRY+F5yosfHXr/GMz
521FM5IAZm32drtaeQp0MO3nqWYRZTME2NZG1NbqWJ1sotP8QFcZsbY537MzaQWr
2PiF70As2bFpreAx9NbIOuXRaPBdzTZOd2F+unWqLdl13sT6vis9IfCQtcYfkNIq
olgty29bYKHA8Z1qGYenh/uqJhO8+WBrj3kLr1qisQpBU8SYOLa6m/UvypMs5zbi
hzJzc5dMmWKMEM02dB/psgx3Qag8Zw7pryAeB1ZbeHQjfC0wUAoY3NMf31ysRVxH
ENx3lMRMz9e9I1cJxMdsrWAeJYO7UzEzZKxtWc6R90kJldxo9tx8hl5bBMjc1cvj
Ry5e+kOD4FiXOgnFzk/8cM/Kh+D3y5nL5Py3OFm657n1fQ3BLZsIJCiPktOh3xZV
+67NKQ3Surz5IBZ9wUN0CoTwvVy8zspjQNrvlx3XzyFAch7cG+snsnp2bV86NTqI
fZcy09x99p3LX6x8gV/FrOPCnqkzoQl8RONiBDxGtJpPUEYy84SBRwuMqw/NbJoo
h29ksCxr8cB/18zn8iYdi3AZaOT/DgrOoYD+RcsSw1twdw3iN1zOMaYuMcvcWjgA
bcn/Ird86DnwJbgXzELHTg2utV+rW5G0Jrj6DtiE9DWlpcqv5J126e5r9E6V4MzO
UWTXL7wY6fWuAdTrpGTKGIMl54rQAvsuebZItuNJDZDHKJMYZm/CWDxpKbd+BO+L
dnZd4w8kbRmN4/0z06hjOe3VgYQLVulbBI2CFW26sBk8rTJz6Ndg7ZzTEERKdbhc
b3Dp6ny4aeom+7OQfgXD2zy2a3QYT6fA+sejE6zJryn9cM1cckJcILzm+RX2ijn4
60Ych3d6b4IjhR+f+XG92fbsxdTSy5NrPApY5nrkidWay7bX1r3ZBKfeC7f9zL4u
3XaS1bwjDyr8p72JdAw4Dyik0WG5NEbenMd5e3JXJebAkLixxTS0cuLQn8wBn7lK
TsUoaLArmKfjE6YkM+IdpzuORE9ZeBQ7SUAnSoxumMOoqEmNHISOki2/Tp/WPaIy
iR+I1X90FzVMvTOYu1wV2EBdrYVgn6ZW+CYvGuxectQPNlF62PlpflixCuehs9b0
0VDwo593DejKK6Y5aI2mQ75fSmp3f5gGhoVyBtyTa3hZlVCbo+VCUw5t5IBP7kZq
Bw0a+ZTKosTpKl6CMdio092njzE7HwNlaS0lX+sc1JDWihilSLaVgKop28AnMO67
lUAukykZw6pZgulZjB+EqA7x6zRCjv5KDuo+SmjIDqxh4m8NTtypnlzP3tSfCB3r
+Rlz9EjViKGeqst2Ww47XNv7ngDbi7Xq5SUO+HYxnHEcUff/xXHv1eh9YFWJqelN
QnoMS0Rso3a5mEzsEHkUtLdwd9GoqfSEI8qGj5q4YsgsutObmrLJTt3hewzlVvdB
ezCGTQwYdDUXX+aVsVPmY3A3Rb4RVn6rfFA1dMEWE++4v91q7/9HJxtmoj5wMuTO
IbVuqVNgOwj/vlNBVE91fYvfmVzvSTmc0MWQZUlClp9Tmx5Qp7wK9LrXPgnLFLpy
Gdg2tYFoNl9JEtYS+OqUGyPWVsLGgggzoCRlOqbydQf/VX93pG0dm8UNdiy84gHN
YXM0sKIXIur3267DvsTUKgvZ9VacnYkfpmNdbI+uVoGTXu2/GV9979DVaFuj8VUd
IvQ5rVV04YqGYc1coI3cEcAoYKTV5NtCh3Fhrv9uyJJ9l5LNsqw7qn7FvuYAX76m
putl8IDVsIaOm732VM5B3bSwsD6jzu1fAYSJ9cCfyTfXMXhEYwmz1X7V76J48J8/
/bkPZeJcNbH5QsgoEGeWfEWrGKPQPRYM5a+W+7j18Gv4+DmDvfAStdC4F/dlZHbj
UWv5qOTEaUlgqrn5LTvrRg5SdGNBoz28m4OrfzTiA8C4+fXAwS+jGulwjiQHpw2/
r0wfONfO9MSYINblP65/OmxItOBtatMQH3G5YVMqs1tpkBqaH4wC+ALzbIS4oGKY
CfzkMv8mg1XYOEgPTjEbZgCfiScdD4xWZwMQczQu7slLJ9CTuUk7aJblA2lWg2EU
u1HrQjmWPkoWWGoXZ5fm1Ha+qnowDYHoBaeLCyzH/1X2GgY9vIcCNNfwL8g5TKRt
6ZA3HZ+nSSnDV8YX9I2yPXGq1VkSo3Pzw09qDFCqb8FbUa1qAw5phSvaP+8yYs8y
/7gj/RCJ/4CItHeHH8CbYeKBJYYJHMPqQmlYbEYnlp26plW0doiTvdhccd06BsWq
0i35S+JMKsX4hUXb2swnmdUiSPKkuWmMyMzuqmAzoHyMUb7M/8pJkATzoe/ozPoD
6YsyJXBy2Tjw+RBzfyW8v66qOH+QnnZf2CPt4iymyPuAV8LVm26/GgSP07Xq0gkt
warHp4sRX5TzWLQF9K8vsaFpIWztyZAiTLUdWG7I9ZV6V0abhm1ozUISoaNUmE13
MHbJIpubSiDxMFwJqLguvjKi6WHpzHO6tZ8aGn6xQKE=
`protect end_protected
