-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
usFT5e6ziBHxmeVita1pe6Q0D6wAmgiaGqo32v8X93wZE0yuO39BjTzHj0cHKdKtk4Ddyf93TVXl
QAO8dZwexwgQJHNNzYZKas3m9r6IvVHTmG8lSlCPwvydf5RN3hCsi+q89/C1EEz9l/Of5h0ShOeD
4nKEIk4Oq9jS0tb7U3gTy2ai7Zw7UFmYyZ/YiTAMyPggdIHajSLfyI3GUOQV+PvdwCnJTUrr2OPx
NTh/68ffbgdn6mwGwaxJWrzg6wPs/VXJBjHlJzjWWuZykDLiwfGJqdUeMIt8CLZD9NXj35PDm7vM
RSAXmRQmz4ZhJjttAfYnEtB9iqBpte/JNQulVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 111456)
`protect data_block
bSrEXXyvyEKa42AygkUNHe2hLSek0gDFapuuCd/aEJNKMSeK43eoEnFfUC8qhgBMWReohEszK60x
B6Y9Pe/hISquLT2zzYjdPbngbIdnC/Iz2h/2BezYorr1XdTkkdwrXqylSPDmFhtK8BIIp3K+vHvq
T30BD1FniVZOcLTUiTcPMFodOcPgGRoMSz8u32KtmhVeQqW6CrQn3JchFy5Nhr49dw1zwExoRvX7
gPXBIftb8NMDxs/B4ty2Thp6AFBSk7APZMXze2QkdshAXpb+DS4Fl+G36sltOWWydlTOV5+Dbh+u
eR3tvOucBHULoZnpn7QMyRWigTB6ep1OSpGCdHxcoGA7Fiud+KdWjh9hjzo4QJp+k6kG1XoMGTdt
LUbiyhG2BExTVhxNz3efwYCri5GUFQbZ9DBWclar4ueo6k0s55wnske1F0WM/lretr9jWyevcVXK
TUdFPK/RniJmhXVa4KVtu5Ypl7nSEM/wY528f1ZIewU2Dot1Ih1Zl7W0WwhGZfvLGkn5yft91sGR
ETUzuDpwTTNrFnNkAd3sgzH2IVMV9LvFHf7Nksxer3ajcYP2/SMjE6bbuDQk4H7hQlovmVRwv98p
th/+dG73MoNajsu3OlQruKYJsQd4IGQqDxAuedqM23+lUhphWwksgOS+/MyTgytANW/FOWxYGlwo
bdnEg5hSERrhqjDWlk649kwCGUmUexWEax/rOwXnWhEC4pB0uCi7FvLbAbMIObVTxuinAROTkqtD
bbS60NIc/9k0+L1KhRikoZtA9E5BIe6dozA6DzXhZTGK9ROmrTd8jI8sjRwr528Rd96gnmQeHMC3
CodMd+8sUrGewa4vBZOeHlyX6k3XuhwXOg+ki6zgqJjzsf1kowH6y59qENB07HFcEa7jpJqIasUP
+f5M9ZbJfGgt5o7r6T2JoULjzskuptjV7A7Rcb9rK52PHqv5V3i1iaOscqHUfsHNAEMrge9QyKSN
XxT87okTCfeKM/6xEzEDTxkruSKPj2zx6ImZozw+JHenxbZg66hmSJSyrSUbX7vfP3PKcjqJrCaC
sjGlXf4blz9smN/Ibbbt5iojGeO6ttX/+fs4EmNZbiHDe0dB9EOavCbV0OGha49vaUx4I/TDuGJL
z4ZeJ7mhs5knZX2G0pWrKfg4KgrIKmf4Q/aV1ASyzisFfAo2qexIBhfRbDY3J9zlvSnXlsaSR+qa
KIo6E68LIim09QeP+HLUuAWStb14xBxI1p6FM2PsW7H+5F8ZAv47SKrwCrZJFc0SmaDQaGy6trxy
DxdcAbrkx1tk0efwOwlHzcOD25185RxubvFnNkXUbg7LzI/jYwvl3ytBpaGGnbOlpqX3+ne6gQPx
26GuAq4bNjt42suzE/qz4rPMp5yW5temH/Xc5rVstgqdViJM9Ej93lA631ed5AJB4yJRF+W1DjWT
dQVXVTTD0gzU4FIUD64ntXPIO6RNq/Ay4a6HFltfx5Ae4ImkMBZ+vUKnaeFTghtZVxIhG8Wq8KPf
K7oKqvv3AX8bS8YQ2qNQV2lR7wK70EXS99I5IFQwGrZnQJ7auoprXvWSeUsRaZxXYZoaTC6qKX26
a2omnu+x/XoNCwFPtV2wI/Kdt44bVfHbOJXzvXPca8y19dv8qAGGGUJeLW2TErDTDyFQU6f1DLke
oAL9hcnNiFTUJqEREtt8GZXXXMnlwg/Bmbp+AMU74vYMpO+FFcJwX7b7PooxNt7tPu65Pc+nBSQt
bP1KS2/c91NFay5BS2KEV829EjZ/08ZlqWOHMvKdLTGsVbvI3x6aZQ3LoIx7HmGiG7zBHiWrJyVj
6nMsCEZPmub5YTULu00X0Y/ycph6+OyvUMmj1l3R82IQcaD82kRzW6Tcc3Uky+ynEgMFJ4pCoUOt
Et3TH2Qx9fhbH53PgRgHs5U3HucHm44KbxQE5xkxVwNHyuqrSiGldYBK0Bj8o07NIlhZ4JxnXles
+CEQL99cMqaXoCHwff7RfWShCoBKbjDXodjtEDwLPQ/x4hQjTlPSzg4St10G1qbLe06HBGevAs8Z
VkKWBGJ5OB6aMUOfegTs3+NnZR0WWM4FHu8kNP3qqvW2+F2NiKmviaI9MLQshDxdj/HRIIeIqn/J
0H9UrPj3sxVuUoGSfyQXOSFMZKS+9uSXVcRJEmja5+1shrF0dazTLCEKSAEqSKETV0Gqxisv6hiq
UgJbNRGZSRlIyP2HrEnSL4+pIZtyHdlFRBmUpoIt3MAnOr/ezKYk+Q51MPBsc0Fjg5zpEw7IB91C
PIcM8V51WvKKsUNl5tx5UQS41bhq9zg9M/iAP/X+u2eoXURY8b2JB/47HhSwIrquNvnrxog+mI4z
l2OZuU7P+uUlGjXVmyDLC8cYrcTT8oOT0y670hi6h8pnYrOb5RxmNe5E2/KTROPOdw4WB0sLNjAH
7QoE5NMB6EuRCUl66BNQW8MqIB9+SoZV7dMn5bp9/hj3MlO6L2I6VBSfTJDvl8S512zIzxyeu+oH
MI9AOsAH13ZyM2302qpeObSWj7xCGMmf4pP9d+ncuyhFFEM7MUObneGVtWM68tVYU8ugWXtMaNjp
Topfn1eupyZR/JNmFCTal6HzBuJTGM4kcJiiGrYFQOrl2aKoJN6bm245HgtszKvhiuehScMncYET
/8x84AVgUhSrSxt0I6Hu+cncgIcm8N2clHGLSN1unBUA/viVHgNPmrcwT0lSxlemppj+lEllOOvc
jxCTjJAWJjNTalyFeO/G/RQtfiKRCU48ppKJVscekweJPR5ageNVOSyHxo73ClzypvPKvfuTATXn
cRmccs2ENDuiAdPe/ASwZFbPsZhBrxfdKWTTFpnft4onTDi33fgocB1OcFdTVW5Wqh64NWy4BUsN
d1ZsnHwczsiX3wcdD6iGazr82AvfRh5zKu8UCLeOimyFAxjO3XDvpDkjFQHOsdvCHLCm+lJpNgum
rV5EtABjkqz6uxqTYBAiP8NmAlDXBPQW+KaqjeuvlGGrFX/IcPIFiSwvt2xcxcRLXPpHbZurk92E
Chy46dRY+TXmmpnFTbI89hjVLAKq4TwpoPOuv8SDfeHBkdDuIFhExHJxoZL/6XZkQXx8HvAeqiIL
kjVoFtoIGLcsjRH70UjLqIhGlxifNs6pmbqKhoyy4afqw+9M/Hn9ARu0MuSxUuvKmm3Sxy+GcSct
EWxAAzcFjc2HT9SfjNts8bWkTohLow7Wrwj7q6katojdUJ9H7PSnFFhX9BO61B+1VgJVx2Nq+3eq
0NSat7D8NBrgb+ZbASqFGpv3zdo94YcEfwEa1Kng0j/EgO6/xmshaoolkjTX3O4AMyxJI+52IyFf
O89SJy0j1XMpjJ7B131VJiowGgPVFYLC/GMhowy3vxZoTb9gG4vzTjV12ttHLSf7SkcJvmzRhAcx
igg8Xz7z6DhpnBZoCQKyqBsfF0jvvchiV8Hc5U0khiXFpBgRyZDCG+GyrC5CFn2nhVEbATWHPEvZ
+KPc8UCpUp2FGx2mBLNbz+uDqkobqV0zYrChlvk8C0kfIZCHoqUcNoezJE+JEFJRdLfZJ27tkeKg
Jgey0fjKEtPPc6tHF2Fp8kh43jnIMvyAtXQcTB0qxhmAgOpakLSSI/pewr8PWnJK5DBIw4pXV+eA
KVt3j+VBVUdEXV1PLPE/qZ7uUwEN/5gG+QPFs3WXvWR8Wd8ZwkeRBitF5tS8+Z7+JGjP0QqKDt9k
DpH18yoJU2cYfY6z0hj7j7g/ru39in41m6xnOpH8EG03S+wJYHj1LQsCshAiCK9noROzwroK1ZGy
hUktMqWbUhh1tqhwwE/j0rT+DyQ3x04mGMZ4ulWPYFN0sXTPED8vp56aknad5C7n7GUAf/ywllBf
+Pz5K4E+81VeRgAEqbRmFbluQZj3Mhp+PfYF76ptOJTraV3GuAj3xzzlz2O1ei/fVyixmJD2jqmM
lIvQg9bDLijivcQJGaXb7I7y6kFt/WQU8B8s0rFPmMivyCAjpEcSvcqRxv42HNB3DNONYorDwmw9
c/y5H4U/IIS2018J9IXO/org+zpH7rmaCyrgjXE7plwhRoz1DDkT10X9Op7+QMQzuUK3Iyrh6M/u
jKGh9/sGCgNpMmBegQ1AHJcDbxF/o6jwOBhroP6Uk4fraRsTGhG41N7O8BxMoO9ovlD3X4Bglnyi
gypbfx1cyyKx7iD/Sp46+5RBVuZW3bIo5mxMNabik4LlHbAYCn3dT9n3xQUNUqDQwo5Ie2c/loy3
qkCTTRszayLYV/INu28fiXBhjerLF1knDZBJSk6D63v5nqYblYBepEpIZJCvc16S3atvt/pFe7PE
MvWSTZ6eWdO3BXGBckLINsZDC8ABZrR1a8fKdqKPNoMjJDiQym7VmwcIwIv0EbLhUpzb0zNS+5LZ
nf6wwzwn2ly4jWzmXZEESIk0tzr0RNuXjHnylyD5EHUPppv6FbaLPsgtMPq8KdGN11ylzFz68kRS
GQERBktMDE+QVE0Or2k88E9iu18Ko2PSWWVjE/kicoTL6HPBNzLeTkUe/4uOJiw7hwqSps7G1UIG
T2pryUxcsp6vnphfuEYOy1kKNdHRcGguw2Z3T3s18jTo2CpVUNgskpcEY8OpAGk5YAr82hIg/rTk
3ErL+KE7hmYGZIPji0KWaBZyMcKSJg22Nrb5XsJ1VkJTPjkfovTYUpiVXYnkfY1yI5Ph9oohVZhi
/m3LSL/cpGbZ0i4AjJxQp1g0Gg9hXSTXKewMW8IQ9L/fa84Fxrcl3iSk5PKWUz0FP6W/rCWYNrOL
0HNhvp3/tavU+rZh+qWrxT80ioM41ls9D2H+geu7Lvc1tw1cUo2DlPCcCjnmDNeLhI3sRgGJG2xU
iM6Cgq5Pycy0C42lNI7hlgjVndIsmREr3nmJ/hOu0/XJ1z+IKk1BC+2laEJ7z27DVfvKKHhglxwO
GWNy8FNEhGna50hWfPcag/kKCOp7UvGXrI/DjD6WT1eS4b4Qr4/+m8X/nKcposIVXJO6mF2ZvY60
T8rBlgY0YwbPo551q5jLRd1U/VjfaPyR9rDx3x9YqE/3egTGFM8FKZgSxn9xRawPpNa30AhaT3RG
lRx2c47/ox1NeNX8LPenuZTgodDIIbJDS+xfhDbC11jqXUxW9vschaDqnPhZkqc3yAShZwdJT7dK
8YPMvy56Xe+NjDBWOBrkqW12azA3oge5EQ5Lnxu3tTGoWj0livbH1MZiDnaiEQAM45Xc7LF30ScF
KA10R+xU1qOhwLYoCyltiMmF6Xdc/CDrqoI8jlzfXW1xquXx1iDI1pbCmPBUrm0u15dVxVdTKjZ9
QaRqwlzbRcWxigp2FlWZ4omuvgD8cdtw915ux1P3KsrEjV8V4V4As0J83jycDXCo4hxQiz+4PXAW
JOiko0Oi8cwusuwpgCsxttnnTiLKcR2nU6ZMT0Mh3NM5QDhLPOuHRZk4rgFZCzd0OF0G9PPTbxfz
R78d7qklCX9/AGyIpePej35+/lrj/nfASuOijd0HWjCDO2W1AeFVeAJXYjnCLeMd+LtNcjjnbBw0
5Roxpu1+W4KRXU8XHZd28AsxuJoPzq1eknU4RdSL92199FwUTeNzoj7bFklQtYXCxPM6nthCJhg5
Dr8h4hsZLjK4qEcoJjGRUlS+mZlMxECzZVZ3IxE9Dfn3DquOEmXRj2S+8whYh0/9Erdb2B9sZHQH
J9YRDRcz0dTpzWS+BT92KtjIzRsTWlFFTejYz4x6VRDD7nkq+c3KOh+tVjjFcIWrcC/XjK+UnD7s
wNZM04Z17Vv23sW37MRTjjwCBQuOGnTVnpgrLtPbYARU/dDvnhubT9aMdsh3WP7VyquSYfo1o9kX
Z0xWLg7M/Pp703wcxcXOZ5qlFNI0Rpurj/zvcaYNmJmNQUe3XQ09BaDNsf2UIhfcEgbER1+1BFjo
L3WefxGDIFyeKJitVzTL04yIGeSftJ1R5TksChjQGnS1EA6+Zi1B5JJ0nLdBFjj9jaqfVKlO0pcn
ydmZZ1G8LHl1FBFPoy0+H8Icb9WH6pyZ0HFAC2zey979nbLILGV1Xy8hzRg5LJ97bzm7VCWvnzPB
N9xbMlmYEw94CUkswv2DrkgLefgrM5Vd8OI+3xnEiBfoQLOjxjNH3W8HJKglrKhbfro/OL9sFA6f
P4YMfOnkBugg0Gk2kTZBFk3fGShkBV0wHMNC6TB5jdXfqnnC26sOf5FIx9+TKlhRh/Tmz3jLcgUB
tkr0oZzLPYIvfGc5N2+XNhDIRyMzsajw/wjc0uQBaF+UR8IpE1Oz3fKAuFcZhYQfAC3mTUGv9nUS
ksPeH9f6A3R+GOhXwbvxpZBhhZv4Jt954ZTjMIZYTmJLTUMG7AHDnb3vu8n3955RECkWLXOfBrUw
YUaeyRzcRGmRTBoahbUYcXotOhQhwNBDlp2s9QknozfGQYqgTXJ12lsl6XnbOtaYLgYXM329acN+
3IYTwww/76te6Lm0K0PB+hsXQNM2yb6LI6EkD6Q66porvyuN6/GqeqwHMsbaseRh+Ae0V7KZjewW
HQo1s5EyXTu49+KfR8FCWr5BgpAXwjGQlN9ivKxYy7IIXUj2g6im25Pb4TIw+YToMzP4xHKdhPdi
82IterXiJqKFPcWasFM1XhPA3+s2d68oMB2S8Yp1bxFnf1iI4hbldUYVKjwXPV+Nd1a1XR6kjmvk
3xragbFeOPYbsJIkc/I7tyO9bsUrrsFaOms/cZ3OowXgZU1JveSm4Vw0PCefn09GEzm+4PWxXTr1
9xsSdW/xzFimKWzwu0+f7HjByHYIpWmlYapS01deCk0Wb3kLykf0n9FTGh+8Ghkf1Ih0U6JaWVYb
c0+Ul5Ac0zfqnifmMwPEyhGarSmPnMjnpWIwrNDGn6n7RDsVkJaESZc8FxmtS7KmznabD9sbv1rD
reA3oZPm0PpVHdrnr4Do1UUapT1imbTMye59Lxc9IE44pop8+4kIL0MEUlafwDOKucIABD1E2vth
kGVurPF3BXOQPiThvHXgNPrBFrtoJyD4gFtnzXTVwfrCow5jmy8T+R1v4GKNBbSaGGNzdiKZA1JS
siepegBDfT55v8XWO1/DWJvviZ0J4rfRXC8/tgdCzdJttiMfNvAG7rQq5K1yt0H4JhlGPLtcDHkK
5AcTGWwO9LKWDsNFTRDvNqAlOsTU4cFdc2lu/c6r9YVL26ljKRJN3Ax7J9wTUdX2tnq+z7jwtf9/
Bg1RpNEGccQf5Pbp3jBInaVdfenOr/1jC3dmfVQ8UFr2URWxci1nnvPdl2ugZvNZBxrE5b4IdccF
gRMUgzWjt/5JOsPKaAgzb8SipwWByKn/L5MeUSRI4/w1RzRn7sn8YL8tu6j1XV7VoNH9AnroqzGS
gcYf5+6n15tI3XIlC68MPh2cZ60kOzJmezThGJfryjwpJ2YoZghYkxceMtjG7QrHrzitIlMeU9HN
d6rhBHotyUNNPG2L8hTOmpZBZI3HEpzd7XXMxiJY6pmQFKJ8xcqy0bgDZ7Bbe/WcCXyLEjN99XuD
+I01e4TSuoTYmogJwH4+cHe8XkoRhgRDM5mnRr1hTKl6XLG7Dentg3Aor/38D74OBe98CcU9audc
2U9GIZswF9BIP0TYQ/PRMc0wWtHbX/v1EUsVVuT0kwaRyKybVwDSWjmA5ywnaRPUbufR+u4r4lGh
vi4+T19h5w9L0VEbJL54g71Y6YvknKOX+LFAeDZu036C+el8CESDnA4ebYDXY6Gc06Gyx+erHdwF
LJz6b4CdWoW/V7DsqiIO1uRU0y7MDPhDPfa7JNicnE63hnJ4cSxyxuPLm+ixgps1JDLJ97UkfzCN
ce5jmqVujZBVF6WQu1B3gP5xy9SC7EW2hUo0Q4pQrRsAxMGjjdquIeuAFb/4z4+w4CIT4QKKn7hT
adkIKAiFPZuTj7joTLCue+FbrkRx0yvhy7qixuoUC125uONIWv3DQHVuy863PAe+xk85Qa1WbXtH
OuqEjOaMohi7dW3L8A0mtKgzG9BSz3rthRkNsvhuUkNNDg6pESE8+Q/KJvsNzbtENjbx/BeqoC2B
nrhqX1DvUO5F6Z65Z0x71fOTzq0vz7oqeTHx2TMfV/feC7B/PozGaS4VIVkewMgtTBASyfpmHg2l
Db7AJcCBHcs33vNCQQ+C7kGBWZOXmWNE4EltYqI6hA0hx7AKLgjXj3xbzsjR3Rt5Enx2pj2s9bas
7b8XPIxBn5neptly0R+sI4A5ofLn8kt5BEv10XRN6Boi9RIFXO/6gV8WRY2g1QL895uqP2a8a/tI
OkzM0vuEFS1F66pLHN708na435OEmz+EVdEImQ6sS1r6uaQgm67UzFJYeF9rmUZhVeAQNzQZ+tPC
O8s++zkiAalDG+6f1YCTAbeFcxM0mYWLEhrxfQqdMtMPYYYftfiFRueSguuKWshWMIQ6Oatvq/EU
hgG1Quklc8Pbee73gJt3y+i1PmXtfIe6sMa5oIUNwZqi7yAJGb0+5Z4062C5S/Zws4q6m+lWRPMN
jxLe8p+WqXb2GVQYW2ewQKAXPXRxb/KoSfyfxQHiKKnUEXm+U99MDZWp5gVzabpZc6RF8xGFY0Ps
kL7fiOz7DAmeoTerYIjxRZiTRi00mUrxDLICyQrZ4c1q/XsNLTS4NJh9G2CHhHmNeJDsKz4se9iH
TX2jINSz9X/mmSsNcDKV7DeyhlBl549dNhW02SNWDqGA0jeR7bagIgngeD32j5Mwq4kFr3tmpq7F
fH6KAVAp688B4JmLSlB/y82fulUl6sPDRcEHHZ2tgcUsyU0t6sG74q0gbzzZqFpcGS+flZMDFduV
aG5gxpc4mJcd77/9pnPIyQTVNhHbiEwK+zXq4yhuiR0jPHPctjYvygS0b7kZbQAmc0Soh/eyMbbM
MuztRd629Cfi422sWzv3Ukbr4aolNPVAJJARrAIms1TlgC5gWmX3Xb8k5WilNi+let7qDmWGO1ox
GLqLYKo7S2OccmBPKNbrxZDjLuXu2EgGh9w6l+TDlW2pG/3ezOlt65RE+DMeWEeV0QBHVhrz6HKv
jMqAaEW37Cqrs2lQsaMrFpBR/Ty/LPmhiZ7xUyUl827QoCrUwxCfypUfoGrURxO7DrQQvztRLPgD
M67QxnoU98n0I+X4JaszkRn4Lpw+GOd2HZFPPN8smp5O8C0BzSpRonmU+hXEALMacTYHBpbmcARW
objW0SoahPHzdTR88i67g5iMGR8dA/TFUB2Art5dkulUbALJ4c4wh+aM+srO0A+H3sSNMPls4GMb
OrGHb0rSxrao5P3TlIT20vngIfJAK7S2B2aSaFIdhfLK8ehRmsUqiORgfrX4yPklrdxsVnZj9zqS
8Y8Vevs7BBhPEnsdczmZ2BlBFXSQ+j/ntYBZAyesVvg7CikXtdGfwhPZXuBjFM6HetZpA1W5hd77
Yx6dhtyNYScVEVLdyD1CfyeNnsCWxX9azwn0KjbJN300UHlwv1HFFi3TXz2/gGbUIn0C6DHjEVUT
8oxlBvMsSWozKx0NCMfLoQ5oN/237H7qVOL7cbfXHB9baCO7gU58WTgRLNUsbT+sXShwq1a87g+M
U1LWmkb2LCncxtGUwyaprSrVnJudqDxShqLfVYDKZM9aAIlm1bugbvGXXb+keWsgmunE2p1SfceE
wCdpqxuAqUWgYEU5niJkjuFx/9BDljrZXa8tcn2Ny+5RR1RWHgzochaOT68oa0T0oUhqy1dHAsz3
3bnH8dx+57YZYjYycJNgLKOk6BrEZNAGnlMk0EmNUX4PS5Z+neNbatVBJZxBKOnnb4dT8+26nJiP
z+V0yPRvWXbO4TLvAerfrpg+vtHWmRWju/UCqwwBfJ8IQ13wk6EqXBUaZlTdmUvKI3pT29f4Zels
Gb0XPb28AXo6WAEIJDx3IbdpG4t3iScVpMjUSUx1iew77ODGYM7P+qmscOI5LqkUBb+7W88h9lJw
g3SI240JhPkIxHDRSLgcmV2SniLXsC0gUTAtXn98HCusJ0Is5LdIjH40VcfuVO3uc/8XjsTzCA2p
HLqXhwyUbUEnrLxn1J0/16qOg0TF9z2ahonKaDW2e54Okb1MAjF5dtYeKqhdx4dyoJ9XmGWXH2Ov
UHiyuySgRbXLTq+k7b7S/505IRiIgPFoKx4qNZwHS/JlTfeEjwmsY7poSVAhI3oO4Fupcd54SeAJ
j4fsVnuYg1AqqpQoraOOs6BH+w8jWogpQDUuOPhr/yqV9/hSDYxU+EO575MvtFt+6bJQauU4bz7X
7afGl2bivIPHN/+n2UdYWjnEoiWrJGl4QFqDLw+6QaS5owWvik6i1p+Ol6x3SHZbwCcrQSByQrcV
5WIGA0G0pWllhYCPug/pmEYasYBBMEB3c0u8Z6XOFI+P4LJ/LYclrAyXHHmuorpKN4hmZ/+zBXb0
9Fa1FPOQhB26w9FM0aCgzqnCB0luBI7DeT3hCoMpCyS0RtJuSeQAYdK0bLb00qrjCKFfQ4kRKu8N
mdpIqQojwHr6v1D03GlzElWrHPTzjEz1SfuXOJekaoSBy7a4tJLmq21z6oQr8u/ERKWwj2sukE7g
uEO9M0WO1ywTLUEHwM2J2HmecP4QbPq3Tr3GnRKdo7ZIn1lrIqAt+twaBqaUG4w4XgvINU69nunP
ehNWqtZ27wsWNthP0kwWbLRLwb7DqHLZ4TgHqHqoeWCCkGpT9bkH2VmTBVggXNGKQDFY81Q4TbCm
okajKRnkMJlQ13rNzJd2YnCNXOJQdppxS7lxVIss0yOqZH9gqRUvII70DCMZU3SX/0bIGRzKGaAB
jeWhUKJq3FsI52sWpD1Wqkpm8/AQtricbJKLYGJdawXwkpnIdFnwQsGnxpHSLSvO9L/i7Rv1p2vY
5YpE8m50rTK+0mpzG0rl5FdR5nuH50sazQnX2t7OOqraSzHoB5sRr1RSHDQ+Gw/B6lCkLpDvlpY4
wp2tDvP+YlqrOs7X4OxVspKDS/HwzJc6FXvOsNWX7fg260trPmCVEGkasbi4bt2qiqhIoUVHk+6H
arxCkJo3hWqg/Nnjx547GTRmnzIaC5xBLW48QQ9W4HMCBrjQWBK0gD6Xy90Ze/a8srB9qEk/bv64
ehXNJLiA/fe3CIrFODAlPgry44vam6BxiA4HwIG0YVk9DXhlspdizjkl4ekipq2n5dkc3m1UANea
4zpfTFYiKLkLTMJIHYaCU9tNE4MqpP4mHpnA48U6AZwJTP7soLjSS4F/GAFbO65G6OyesLvO22FU
8wBQN+SSrsbrW994iHbC9qU4QEuIzO9RA473OCnVoik0PLV12Ml/U0PUImeYXTCvljEZzp7M7tDf
2qSl7pUL9VeDQXNcArlsV0I5i903Q1B+aOYni8eS/ZFHo7WgQ3kB26dwK1iIHB1KgKXwGy9mkbR7
0E9Mt7VRCFM7TsayAmJAyyuz8C/MntZfz6sfADvm2gpueI+NFuwtFDJU+yrJVDY2pWYdtBWywhNt
rWkX/BAlrMktkOrr4TP46rQda4NSBqT2bFuE8XZPHNq6lRyaXtBHeXZldFpZukZ06d5370wcc2HD
FouNwahWzvjxVJDYo6JLZgxDU9qXoJWVMPdOMrlGN289K916ed4SRlzU45en7KHUiNdvRZBjRXpr
z94YBt6AU9HIRpVegr3NHqK3JqUzAIq6x+UAiAHu8++N5YP0eVFCFUbPfYrerScRq3gxyAMJNVaL
UTGjAOoIBKbQnAMnGNCJUZENK7EqI1dui86Q0KDgCQMbGHJYGrkZLeXo15XIN4hXsb9s20MFwu+U
ArRutny3vv5kGordfnKD6pd2J+scL/X4dwDehXXvj5mUOaFEQUZ/oU5BiezNtc86sWKGfefeu2M4
7CUeY7AyaJNPoaEFgL6UC5sCYpMlGZs5UEIXWZ8WWjm7X/ImZvB1nMehOPyGU0GjhQ/y0T/yOBTO
+oR03e+9t6DYuidxqo7L5SoJkQZxHJGaeaMTioR/8ewfphp8jldB5F6/wT/g1UKT49VN0J/pEIg5
pYOLtPXAJgFbveW66i95pshjQgOH1sCVrEL6O0D9kndyeGP1RQrO9A1THuxIhNZIWgT7oOP7vklT
kvdkrsmhVT0z1GvHZwonoHt7QuclTliShvs8sYTd9uwZDHx6Bf4+lw83G2ibC5EXlaAO6QFzkXnC
PIQ0K7HaeCEz7k5/d+JZhm+Nj046m3zL9ZMRbaeNIS2QwO96ESw3IZOPXENi3dJyuS4gl+gF10S2
Q50tz2Kvl1Wb0TE9ByIpJLD+d/4VS5QS8hLz0eXJ1mE2klPDwu2mCDg3OQ3zuzdAViPxKmD/yvww
1oKFO/D7zKS20/4hnIvAsAvqKfn0/edvy1mu4xcJu/H9bZY8j1CzsPp9ABy00Ptunf5KFRwaUkvx
fcccS6Qbj0JZbG5+ARTlYKqKTDHP/sajyU6rtSHsYxFizEHqtxlrs8ug16G+66aknKYu31lRHbK0
22qHRNZ9dZ3RG0LzJQ1eRggvqodEKsZJz3psvOihBtHyfsANI1VSQu97IM3rZGjsYcM/hTHh3/og
QkVDs4WwlkXQ4pX2VCXWPtuyOeuZ5QXc7z99crBqMDV4EGAknCbK+ytgSyHlu6ylZnjLsmzsXpuc
IFF8IeWps9t8Gl7uOEF7XFWxvRDqrE5XiPNAgCb65yfRzkyE+fJhUSr/QukBEsDJgnWThdVRtNq7
PFB8X13HplL5af38Omov7KPH/rseSnoI36ps1bBK9VZKG7JD2uRHbn7qsXPYZ0QNh/rV6lrINTdf
+h1S/OTH5128gbtZZtSl3smAuNAjRn+KlZtnnZ8Ni60scI42tlOafD9ej7yg2fHN7D6GgvXsi0yv
Z+GSymvaTbEZlmMBG16owTpB7r0LFROB+uFf1T95xaSDQR/c8oC9jqtSVDdVtswzagPQutNeXRdu
6iOFeq/1ILyMgX1KVyiZK9jcIhL7KpbidV9ss+WNbu6oTUMNfnzIAvSgW3XXZTegYECLrLNKIHA/
cagDnbs5diKI+/cV5WIRPoRwEKGkqq2F/NMF6L/a6HSZY9bkMXSJAh+E9tD1TnEQVHwzKkuzGvNe
tuBsvluNB21P+pk4flG0lxhSIg2mb7murSOm3KHJuz0x8YDBZ3h33ziDhFHI1bckML0CAX0Ko7r0
IC4Ea5OpMGzs1xJFsR7z1WYNd1xtl8u/44jxJgS9M+erHR0bg1OrdYpPVQX2dzPIywD5z4wgPYF7
T08CYt4FRxfoaBBBQGKeSUp5WQ2bkWm2Uruk86kCu0tZjVhqjF/gsAYzp9xh2IgOhnCWVIXV7i2p
RKJBuRGIqVAv3TLKion10Ne8HrV1zxIj3Esb2QJgUojUp9fvYOpVvfmBqP3JdDsf1kMYBTVK+hrV
td+dOQy+U8CB5ZW3iGwmdzF0a1zgscsu3YTa2p/FTbAglV0Zync2jscmKnM6ZJ6N3a4sdGIoizy5
DIJWBUiJwmiY45p1SWH6NRoPtTbfYqoFKmNI9Pk+PnGiJfag5rcFRBbihHcMIlIb0ITVea/lSyT6
I/uob1y31FBDkN6flMW/NIFuJC141g4CjyfaVFcN8ZVdEwZIBa00N3T8O5E3Qva21pwNslLghFGu
zm8lN6WlhTqaqSB+zCVDhqVjcanGlZOzrpmN8hlt30b/gQHEYiyoCwlAG83HCU4cUQzq6MJIRGpI
jD+/y3gEk82I/XsPZmQVH/1m+Me36SHmoH/awXwNtbIWdfnnrOO1sUJaPvt9jSlvGvTwxu3HQcGx
oi++4ph5IN2MiqIQ6nfWFCp8API6GBNSON6saJ4AZbGx2jyKPTgyY769bO8e9cTGFnEklERusbU2
i60Ggb73n9IfmSHQIofn3rrUR4iVOLqye19xAHv6e4d+/9y5HocGAgUntqMHrAAnwRiOFT0DtEM0
E6NcI7qX8LJNu8YB9nL3/W6ecLtiIFxWuPv36CDZyIvblX2Md5CcnppAjSRfAvoR9XVA9OVqDx/K
5Mfp8yzAG1VXgH+7f5mVEF3E2Hm6cPngUSV4uoNncUf6QAMNgzIjteYOrM748hgj91SovT+DiluD
3zq/Lid0RFPpfmE1/hwQfjNkm9T8kMNqMXS9cb/XKZ2cMn3bRM32o1YG+9s7X+VnyD3LUsSLfTJ6
SvnpIU31bL/Fjq/QjNJzx01F6QIANWRcaYkkPBFO+J1iK4xmPZWMyIwGoNRVUj8OLsTOqlwTSFRv
IDTEZYVD7pARnBaDcBmwdV7oVujQ93/g0p3CR3IMYGLOwxa3Nd/0eAVxcVJX7jpAx6vdpCn44i2c
5rh2LgL3uBF0VNc5GhgLeZZq+nYRsskmYeArza3vdIC05zh8izq6AtxU+rbnhfwT3e9j0FHDX3lR
ersM+4wNuwBMpqxPrPXvMNT1voSMN6sUMKCQMZ/4a9wMIsAxuHOIrVQhhPiD6GPhQl3gnUkd7B6I
fKZqH/asWZBN9v4yYdczJp+dkPhNffMpyRDA5ow7g2O1tTvu0RRIVknuyq2HwDmVnZK/zL7N2YcQ
6V6f23jQoTnho34SSSl+Xf94xwfd0deGcRV6CFJuOqPUk0WbssKliv8JU7OaW64O4rXl4ObVYzOX
N4a/kQsK4U3kA+IhbLexX3VlvraV7nu6n9JCOxQjQQdV+gl/nPZMQRrLVRtKpCXou+fUvrc0nF4G
EAWe0i9cqQejbzPC83rcqwo+LXiymLjTz7pJGgGLB2MILJUGaw3K/of88AFYHSvvqbaLnvPriG6/
EvDcQIVL41ys8lClDm0QboDMJzjM3j2rj3detbFuyhmyMgAmiB3gKJVeWQ18rekQJe7yHCdaOOJo
7GfLoqltw5kgK8vJqwAV5bJGGZnyQ9w/6OtkD21Qei28F81NnIwEAMR5tJh0/a1x6Pml6AI0xQI/
tzvogNbwAMU0ReVZXW8fvmm1U8iwyACPn2114Sm3F2/Kn8yDvtsWaTb8ys4E4zSXQlquLlDojfZl
TM6UTLOb3j44IveZkwkiDqCqc0yatRXm5Uae3KWEAWd4QaaGcKb4Xxdozkae6wQEdOFPWQMi1GzV
zdlboKe9wBiMvzDZd4uXpb9kvPh/wPdVc85rlkRAPweG4UOgCoNNOokw0R7fzfSgQ2Dz3+GcH1w8
gDjT4lzSEbH4GwoZVFAX+AHb58XoS/5P/OFBbHbCjYqXqqxkA8de5z8yMMf3raK2HXNpnpH+73eE
8BtjmfCs3hrFIBNFgy2jF15VAmHsSmOXge5lt3VO7pKhEVHH9ds1Qc+MERH4sDDYyMkpocbPt84+
9+vKdXDgO/+OCAHF2qgMmzAbnL1HOoi+KpNw9fbG/X0AFgiTgKmVoRe7z9l/VjSBf/xRwG53cktJ
M9rY+62jkCzgrnu/mG2WaMDsGnTsPdxaHnTdy18xq7EGTKqcACSCORfDnUz+ljLiZdkGMYlBRVx9
AAcibyUV7in75JmaSE33dIsS/rLqYBLrgQ7V3d+Ja/DoJJz3KszDQyf01FlOx4wfice+EZRThDsC
gzRMurEAWK4XftmRvbKRSVxR6fzoHDRmDnp9055Gp18IXYCyCl+30T42VpEYNvnX5VWBazFaDWvC
WpdMIj6Sjw/krFd/YpBylxYP0A2uFiu1AFH3Ya0Cc2sDnS+KgGzvjzEqUKp1IbCeSvTP0yEuLjOH
LyvUoWmdFddrzGiknHeoxD6/84c75XAa0Euowl+vaarZzZTWroNGFf9tQVoGcqJV4Xq2MGP31PEE
/+f6hO1NDDwgu2zXTrwmB7aS85Kr6SAA+afVnA970Q6T+s+n6nXC0rL85fZBXZ0/B3XGJ4wueQNL
u2HxedPUoa7IYFpOi451B4A6aDxf/NbWDTBumi4iHOebzpWtcT+mDu4RUeKc7rzq4Lgj0mhCS+Ls
Uful9Jgx/rp5n5r6Hc7Dn+Hu6MIvGr4I2rAhHrF8iJ6Hc8XAZVckPO/uxI5ajOT2tjh3xw/tKhTe
DCUfSbArWd/Zzpbr2I5osqH8UWG9RGTdu0KYetOeAMrx7NNA5+Hx6F5n9CvLFJcWibNBaoiGG3Hk
GK/AmdaFd4FzG9SbPUJ4N0DjU2SmT9Ygib5R5i8f2ZdQVUKtoxwgYGThFKd0e+c0pBiK/wPY+Dzq
Hnd7hLkDbgzmn0QYYD7U3WgQLMm/F79tT64tzF+K1EacSAhcTfjuFdWDKrTDGozEX7Ldo38z8yVd
0SOnIiBFIqycMHW9RZVM1ZNErJ6oXx6pFCbWlIfUiKHkTKbR5/0b7AdEEcGhCE7Esd3Cv+UpTBoV
+ueftIND7VtVk9GBdgRFYn/14TYmK71RynnRA9s5cEVXB54k3pgskE7B6b2n0Hez5V74KZXBc+EN
yBRuB0XTplH8sUQ1B7VyqtJI3u5el0mvZ+Zwtzz5hJMSQBrDbgWNCXxgo/Hk0lRW6ScD+aF2o0BM
3NnZaOpRwYwW7k348dY6jZykYCM9sAK0G/1mJwH3YlYe0Im5K/F9nszrUaFJ6LeAj6/zSzJtwsOu
VvQ27b16p0RcpW+1dInRzjeN2TV3WVXnDgOqXqV2A4yELOEj0kV7gz47M+8yFMm/AEZxky621D++
bL58MqkOy4iXBehzSVMiL8gN2yM26p1SQqfF0OUsWs1aTQ+GZ+z7ibNQD6ktVKPzZ5DzhpCOIbkq
MYHYvB5QwGVJCou/T9403VCiduW+sPOmH3xVPIXn++yz1s+9lCib+Gnl5nyEkyuSJb53sIJTv/tg
k4YU8H0Kfi8rcHx38M2Iznh6AcvElodBTh/TLzOgzY4iI6eHr+kvS73CLYtSSGiv/EXjHoruELxM
mdG/2xKM6G/i8mQj+qMrKpuDewk83jBq4oVKa0FcHIaTSE1qaY/Ci7N9H3lB17xEZR9irrjkAc3v
SnI4kDj+yXpcMROwMy54OxXs6iH9X7/EzbeBDs+bsn+rUIPumf22pFpw9XRSlvePtBIiqv9xBZiq
O6o8V359QWmFmVLuR5RsAjqyq34qC2IUztS86VcCLezujBxVhPhD+B2on1i/wTVLkJPr0FUUDaG1
yzyoEJlxu6fRcLmFbFjEtTpmYv8eWcMSB+sHEGrpdoLGgNnNNfriaIaRkTSasO9UqsOwhSQ9EwsA
NmVepS5jjKCJTksbS5fMst3HfxLucOd7BUTF5jKVXthxTjrxfFfNy+0PPw8f/4G+FRa4ZMTdfGDw
boPx7Dfk5Dcz+xmSOaY6DKJFRfFNbpqygsXHS/na1ailx7+a43dULUFwO5ugYXwUGpTB/DoLW4Hl
4eTDRiJAO31HKymUOTxbiYKwPxIz9UsJSCDZ0aXcGbClRe/NL2p/KgmfwcFFTCAdistVyPT1MdUc
hd23FagZPBIga3x1zcXkoVicJ29684la+XpL0sb6H+ugp8vSQ01YX0bMkvspLbfJnF1ntdsBRZiu
6p4GiZMkCrSb6YwNBioQI056+y2J1iH3oedqE5EcrJJN+eBg7enNEr5s2dxp0rgb7wlZwMDUOtvo
57XyczrlERIpcAjzLvITlTMLII4gupgNTbCRlsHZU1iaQt7qF7VZD8IoKam1X74A5TRUZ8/ahNrJ
v2hPPIbKqP0AftI0XkkPsFPpg9a9bJWufXNQoXz3iVcdSzfz1gSynK+o5d4FPMzl6KtBdHvw9vv4
obK5lqIxyX2XFnIdXivX51yWGf0Bpwc5A7PrkRJkLY6/7wPk8IBvZ16ZpUfAOyRnMHEP22a+uukv
JOUziR65Hy1VbXm437OQZL8q0qBfUwFY5AmmRn4jLudxtOdspg2vMVtD8i8UMdMGiFDxzf1Jpgud
OUa7Ds7/NiXpV7I0L5TYx7/lZ/uGtcaLNpYQc0ThZnVzmqkyQFAIRswOrg8O/aITf7UoxLBU9vgO
HoxhtMDX2BHMkZeqB2E9euUuAJ8IVyQCorOhApUw1wShq+TArSboBWKxRMCE5Jx4cEkaFBjvkfmE
3lxre31J59XMmKoOPv1xVBrLb7g1HZLo8Em4P207zspc1DiKy2sOIsT+L43L9mzmW9DD9Kpa+Whv
/PNZg4TLnMTBelDwdE4+taCAzoGh5B9BcRn2qZtgipJ4eOcN2f5Jqyee0/gyIOCSoLZ2dR98xnhv
UCW2qyexRi/cAgsuVkUn+T2PCeR3lv//0gTORCnDElkS7F2DXksKqEXAwqE7D2nRG2wIApp/AtjB
p8DUOPNQNmcB6fC1Q7/UJlpEoSHj09n5uXZ6cHP3AaJx0x3ZLyOLY1AE4iJOj9wnSjyMyk3ZA42q
CzXpXieByu4VvRUIK5DUNZ1MFm1lucKL9+12kYx0w1CGHNDOzzhHKbwiYy6PP1WPu7C08F1OpeSS
ftgtH3Kpe2eLWSZ6DliPkmxf7Z18W2DQ/9E0O8S/d46lAtrmvLf/hL4MPoxjwnxBf5bF0EIy0VdU
QeOwwhB1I0f6mH8cPgz1thiquRsk8oWY5qOQAsQn1525KTSF8B8UGAZ1zQ8GFdin1Vu74cs2NIEn
Ij5aCAgwkvmvZvQhaGDdhqdQyJgQrrDvd0SFerxGtTd/b03mJbxmn7f+0VmdH8+DuvGdVyh3gkJo
9yO+bEDxXRkpA3xEfDfJG1AB6SStpQYEg89J6Lukblphfz94WHdZmm+jb7EURTllcSo9m0YfrxlC
RO+KMJiebv500fA0VTZhL7gJ15wQja+CGDIQ6dtoOZcfctU7RKP+avMe/UHxfxCN+RCBoe6/2p7u
UvpoOeou4vZzpqxHgwaCl8hNfFZG9N8iDXbSFc77shM7ywIVx8T9yC5nymSMHD9pmXaR0B8In2W5
1B/Jml+T21TFanisCtkJ7YPp614Hl0MmKBeZkgNC711rNmtBHxAGgjn3B5p7V9KZ8NVZbUsGgRyM
+r9TyZFE0SaezYw7Xrbg9VekfFbq3p4QRodTtW9oBsJGVBVaKIicIGPtRpCO95iSy4R6X9EMiAZA
EhIDoHj/9cuiRCJzy4pG+EOh8DFUqL9w2qgQ4gcwLupZVkm7bT+Iaf7IoxDcv2Lz/aWTbPedkZQW
U5AlNLv+K7qF4bId3n6I/GO+EglHhFTx6FgpuNO/LAl7ybn8klBDbMd/2mcgmuViVzX3eTh5jBPp
2TTJbfTSNPPSr6V9hPyzEfZbwNok+MQMRZZChuZJqw/08c1sAfebG4TkBq4Y/dEuGc9qw2oVVCY0
TOlTTzJQ77JtYXRsI3eUBYJ7QjR684izg3FLJgzPugGm/H1DVrsJkSvpMFxh6vfyzyZjHu7p6KKO
ibF7btjAWsaAfhC6iP6zX21j3wUrVNNujX9CjES/gLp9Vtlup4+8uOJ+OhJ8AjNPEk+xp+AT0uYa
zJ6VCOzkdRVMv3pjCrWk1cLQr2qjKvm90Ib2MbkkslV5dHReCqagk/3HZL6Qarjd2tozPAsC3nN3
+YBJl9ipBI/ud48RNvvtZvHacBgyME3v0AMfmfuCl5DAqKNXcMelvGgBhKt+SXHjdavWO/WxebhW
W99q8INRTF/E/09cKjp3QM2kE8nY8oXeFkOtAwPNisf1Mofo49awFBLEp61F/IRp0EkwOlXrT8VL
tHxGYD5grBFOJmOZceA2gvGVRjAY1jeruauiTEx4bJO5PbCz33jOPcLlD+8Hv9QoRlBP/o9Q5C52
C2/PQXfplZdg9Uay6lH8GG8+nqhiqYPf/y29/htNtV6EB5qo+qeZAzSObguD5cKTumFkSqKoYPjV
3Lzz6hkMB1hUoVf+KHPbHQT6XE2Md5d7qGtFP1L0XhbdWhS0Cp8vG1G4MyjJrCuZT313BEH91Zo0
dpJNKzNmvra/xUHf7iE6v+/efYpu5BxtelNo0QnINYlhO7sc9pGInJHXEfxBtIqyG8ES8NHbOXnW
p0t7XtB9XqhXjLDu8rPFbkSm5O4qGwBnmrnH/RWrvMgoKfqk4X0NJFbWtIjtfTLJbHchV79EKb5s
ru+mqwEDRmXUaxwq47bjhvfxxXjG1c/CJfoSYwedqyMAcLAGW5rJP8jrObY4EP2GmIob3mK6wK9U
iuoQMzo6qtqEk2W9c23sS1OQlpiRwaDhgvEh+JjeQG0bhrM4RHaYuBRLGst/5HyZ2yywVIj/Kpz3
KFSNMoyvXWv8dY6xg94jfYhOq1P+iLLY6pXjxYetP5PoSTrEAYVfmqghHXZhGGlGvj+KKtDYbaBP
q0eX9TFRGSGsToZLDZrk8OBDusfcMsn1t1JRa0w3pLT8CRXKAr4Lm1cxJCIGkOpYgM/ImKORoZ6g
81FH00083mU0fHSiGIlsNCAi6qyaEdbJwCWj5+1qjgQE/xCAGYoyhkLzuboky4A6LhPVX61SsPEJ
/v0omC+hXF7B6tRwNglCC/fVDomSo5zPvUNEl539p65a1U+yA5VgiPG4smFllGcVqNUu7pPo/DMp
c9n4JcbhczL6bgnINeF6oKVGET46hQ7za5tl+Vo/EGXn605XQ8WQWULIEdZFtI372iFTO/sXffUP
TLZX/5PWXotBNah13oDt3e0UCR7FGmAXQoabQ41iYwKcuKPhFEe82oWXg5MCo6JaS7aalMHdoOyh
51JmPiCHnlSy1hjteFWjeDATffdywcWr0eCis5n7hl5qAmnVcMFoVX0TUCJnaVAcgDuLVIjZQBOW
IQhYHuju03hKnDbcA/O8OulyedyLzwrnk41GH1f2RG5aJONaKGfpF75mXJnyfmCzbkn4hfXbYo7J
3cucu5BPka/0Q4PAAV7VfAKD0cmBmsRC4bRVS4WHID9QaBx6Q4mtSVcO/7JoTbmGWbGiTkXbRfvh
uCIzPvHkGaD26fDkyuRjZ4PTnsPX02NVY3gxKVxXG4Ewm2o40x4aRj+4GaDDlHASVw9j/dDYiGqJ
ujOouAGOmbye21WZhY/DX7/48RNOX1i3tUs9lCPX1qQs2rINNSA47eLMXXsON0mvNHvQYFr3gVtF
ia9HNaa3Ehiwfr4YWsHCC2WOYVUkPv76ArUAPed52wV6A3IfllbCKfmDRpIfA+Ikbpo9HTf8V3pf
c/eCZjSNVitr7UlFdN53G3hFiIDuTuxqyJXlVTYGh+Zn5OGIOacsWRULQEpZBNJWOei9HtFiB7wW
JyG3bi4o6Shw7k/uc2FTCxSYim2LRjkBOClZaCYHOuj4LQR6NSs4xy52V5zQokAJYs1/wALdPn8u
GgxfW3XaJvHX/IZ0g6yFrGIKba9NjrvAp8GZzvGpsMJUAX2EjWo5u5+/qnx5o08gqwejY36pQXZz
XP/cW/YlyDupRGlHxJ68uhYMG6xJL961aApWxvb1Pmd0oqE9DmIduG1GF80cXMDHQFkDN53j17us
WmOCTwPimfQ47HN1hcXYgq3mJGeP9MeRSWieXFOWCUbAEjJ2xbDo/QruV4B0RJrULmSxYWXyYCnD
zfv52glN4MQoNbyEtQdfsyK3sTT1UpsrxtS0UT+6nUwjbZkH5XbW+EATlfksI2pnExBnxDs0sEaV
FOu4MkBOi7OhP89TzCUkc73QEzBX1jXUM/vYRH+oprqzogM6u+yxU8eSaqrQmJ/Q3lmy87VZexdl
VNHGTCcWN4l6ukTdMCp4fs+FS44pI8Y5qYNVcWCQ7M0eww9ma5NR8IUkgNmO+XlW/xkFxfb+aV8E
JE4AxskNJHGioy80dywrPXHkG8ye6khGV1v1T7SRJZxjUAqQcPdEZTyUDYbpD5uQx0ouiLqe65u7
dVilJSrF/fxEOZzF/Hsq7c5nXYRg1R4DgO+VVTRzCrmgbpiUKTgQBQw2xtSQMx6xsKYDLnFYwzP0
tQJXzqUFTdA8Bi7IpfuP126/DJDvFtqbNoL+BGvxnzNw0cF+avLZBlf4LqaU4FyjqMSxqIrdqr7G
vS+1cgP6hsPrlE51qplHpbadMWWHP2E7NcJ5iA2k4A7UlKjDVRN/YJId2c0e5vXqC60PH4tWM1bz
77Cwn+mLQYJYMhKiy9UHMi6cpeR0DvEHfwIYfUz8hSGFKx8OCDB5NmzltAUMdGRY6Lra8QjEj21X
aw6fuMorIycrOLt5HLkZmQrQAUI4dFWJUAhmkeD1Eo4eQRxXxSLb+lkKHtukjA3H+rDFwzWzhE5D
QY0+FewXomr4otpp33ANffajwxaN6a8S3j50IrpJjrTOh7VyG2o/U8LjQr3odS1h+Kh6CMNc1Qtz
ht91DLcdwKBApTRQ74JAT84umD/dAMs8bifiVlj/rQxjFHcv+kdejpl+ds4awAEFZ0HuSWfbyMkz
ruOSmo+f1zvMgkwrvhPPrgD1kxM9Wbh3ISati9Docy+qHxZBGpRY0IXNCdczGtc+1zUK13A7J/Uu
xM+Z9F945NRJF929HIVDUIW77jIcq7QJD/b3yvX8GSHfbByhwNRxRdmSdsNUhah1iOW6IpXBpWRa
YYtrHyP4ypp3uBlkDyAa0bgiVSp14tOoLFYaLDxDrEGl3ROUPNBaoF5pR3zGUcyHK75V2DFvHqD2
T4ylsYx6lqPJFdmYXTBL96TNK16oQaYRM/m7PqRek7HEwSMhLeFJOXc2/d6GGew04FgAmLVwgbqL
w+0oeVHCTMuQfMAjqh1eYYqQTQOl+8w2UYzrT570VYaYEoqHBzkmvCrnPL34bKaO3Kby4as8pGNO
YPJpLYB9rdP4ryL7PY1t0EUhLcFZBodDdzxa8w7gm+NyyytELSbo7O5+F4kaxJeWWMlCU5LttcGY
17yLq0E14gVs5XQru3fmVtLRvfuuH1Um6c1BS7DceWAm4yZYn19uc6aeswC8GYgY24GYJj0Zt4LG
wFzPDjqi4HR/DuwXfSDic/j4xAIbHG3XRrsEg2Z3VpugmC1lk46xLNUfJj0Tgs8I0LiTeXFqMQXZ
hXG9GQKn0Zy1/Uv8V+fRIjE1m+Xui48sC+QEmK1dfSn2i/nZDLNChSHDw4+N/vLbyKAw6uhomwBJ
DH0Mfet9OL46AjFAFm9nZV4Mf32f714P+Ii+M+XZ3N8zjuGFtCRjdC2sfiZM48w2JYxcOun3jDxE
2D6rSia93kHrDqWGQAeiqD8BmNazRNibUYH3/+P3VLfc/mwKqSDPi//xa/dU/z4IvMUllzJG1YS2
96TirVu9J1swSDwX+Jyu1nBcBpHgBnx45HFJlCJ0V2OSNHPUjC9gELjxTapHyxxTYJnAORWd/hAa
x9snjmWwdRFkPQZ1DwpZ7y66wHVbYO+3lVpQ7jphCdeMfWN/qWtQzlB3DVXpvlkV6gZNQ5giJiJ+
khMu4uxAQ6/q2fjk7tK8POE17WbLlBiJsz0Sc5Lo8YSOtxYiGnBeSgc3D9KCftFOuffieuaItJvu
RM6Pu99P7wX6vK3fPj4zt1pMrwIchSjBci+8nW8JWbR2uII171tVsQWnlmZyDHqFBnwXtMxhuk4z
drN57jkOCsAmHT9wdQ1yl+/gobxD7CyHCmO06rH+BMRL67terc6ibFXnZ322E3aUnnCaAKM6RyuR
9Bir/WEQ2vM27+AMKFPp4qTVblUNEEviBNQvEkYvvpup6yo0suko4JCICQ2WB0s+IiU9hbZgg08N
lVtuMs9tZLi7CP0ea8PwA9BhbmYWdiHPKgbQrgHrDpF7+HRS52oaDUyqaGUCGD0xmjAo+Te/4KX4
T2xGYZvynuM3OFN/i433u8ZyxWAzXXfaoQLzzZsvynTivNT9xHz+d760KeodcvQcXxX8W/G0x1HQ
FLcdEAERYMk0a2IdYT1FUwNHP+lKn+tPfLgzsXbKafKBPs6TV1ftGT29VgTizREqJvob6lfnf3h+
N8ykwqC1FIUKR9ErNkf6fIKoOWN3pX6iro6FKi7KqvxNVE00kH3OCHB1QKaibEQNjld55K9JfaaD
wl6b+PAZYIjjD2a87uqOl+/dOjy5amQXtneQv4l2RSxbBg1cfC/PJW4pUxLAuPAc6avC351I2Fkj
6FSpgaoADLRmWbZBxBCcvQoF9xpzMNP3Tk121LoOtkTHZ2r0JNBQaB9jYwSr0VhMvg0ORVCZC5OI
kQl7uDaPQgtKxoXdJKW6VE3FT/0kPVpBNzp3BqRzUxYl78HTxuWVUGALCVAySW1jg3QHRodaE1bm
evUABgKn0AzcRriR4YEPRBzaXVnHl871DVcqbeQlDyf2eNFNbcdL+6NaFRWuGpYSJnC7Bvj3fruM
/DOu/W3Aaew8xPlJeSb1MBhm9Y6bcJTSNdi0pcoq0s+92Xjtyjn21uXC5Xp9v6f9NDqXDaqzuAK0
HtgdXg8N8CIemXcpMV7EKNXRb8U9Q2iwPJ2SVwvsUyk8GWrvAICEWoAq/aOSt1sE/ZqMMNnYRrDj
Vl91bThPQqR9wx4/glOabpDsLIwvwpb/glGABQM+Io6bRvePIsAP0skyQqvUlco+kOBb/hDKRJyY
b+hqAwH+9zAZcHdYREarJuGr6lEmfEGyM2r61UXiasUJCPtKr4SCsTA+hqfrGVE7S2OcwzMCFgZh
gF0aTNACpeIsGWd5jKL330I1c5U6/2ZUHTmcIMO+72Pm4SSkrliqsnN2LDOKIXPaYN1SvK3pqImL
akiYn6fU0TBtVckWMdXJipbsLo3ODUPVXF3B4oCOVgaojP4N0uMtsZ+PCKeIjYhSgjUDND0/5lck
nZ3v4gGk315KRDWF9E3534VD7kInpnngqpx4Mgtl2GDSRguW68a6HUIcc4IUtI76ZUTBbqdHr1Fm
wGPtl0u8rbUnyNgpSmMD/9Jdam7yunhyodL0Si9JzG4IU8zWlFzaVLsR3rFH+kbKC6vDZ5T+Tn/w
HslwypN2+0SLsX4Mdk0gjN0XAnjlgbY5MVQgRLz0BeqAyz0ey9zf6jOwHO5FHK2TcfScYF7z95CN
nIq8klQ95UImkkZ8skbCSC9CEHXVF+MNDt+0lj7HgEPSF5yOgshIZyz7ZVaBJvEvlECohKVCVvo5
IdV8PsreTdsi8TK4Ro9qpQkfAmY1aPIGth9q7SpxRN8ZgNmEq5j3tf1w8fEtsZj4JaPt34T5EoEP
MUIIlLmCJnXeKg7zZKvwwwpyfWW1hluNpch+0Hv4844A7qbwr1wDjLEfhsib9Johmv1WwBMnkzRn
Ii97wMhSwf9a7JRmooeZcf4iTpFAViWSX1kzHuEVQ7JvrIXP2phkqCbQ4GV4HEK/Oeoppfojf1eU
i/EpEAOS1MNQFzzJ5XCeeJXThCkrdMVSyCbsxN0Hac41oO66ezds6anZasYyIZYGqbMDJsx2+ZvK
yKlY/EjO+Ijk1tCUPby5qNanFWVi8rE7h0bxJ14fVM93bLmAjKNqE+d5Ea2DZ+Tl8QiUWwOhnZQs
MHP6foIienrfwAdtFxScKM5xt6iJZyLDG0oNUf6APj0FiGY2OXvOJVcULce9/YS0/CNcS818Uj63
pNlqeBLCOHMsTtwhieeHqWPHye2L0R9wLy/cOzxFR9oF0Glddp5yhkwAF5eVagAVvxSkaR46bAfY
O0t5AaGSo9IhIbwFgAcBdeVQmS8G2i6OBlPItG/OAmpcIFTzB7aV2ZeQzR5+et9qFA0reXKGBb8L
4LboLLPW+R0f07oIUMNZHQQSrfmMxJvGnuRXOruNiKo75P/BqUYnr9/iVdvMPCGRZm1RyxTJkhvX
y3L/0HfNf+4ZJIHf2e4AzxhQo8P++gmOYRXo/rbzJzRpWQUHWOZbZx2i5NnjDn9O/cLNlBUUYKgM
FUhQfv/ZMnpJvar1Lkq9f9pG07ZTRq0mLahb8mo5Hxcw8AHxS8xcjEObIwjGQH7Dnk38leINIK+m
WCz9/3sR1C913f/4m1u3bZGc/8jweFPiOgjaLGCQh9xQ6YDmIW5XL3IGWcct9J0MGDB52Dg3Affl
VpHsSHbiC5jALujru9IXRHidLy5KWzVM4DagOxegjVTTEt1v2HizoJNvx7emFEaRf7e1HW8JWY1q
Xc51RfBn8J9aULewa+Og0DhDvD4oLlx/Tka6R7/rYAcLgfETo6ux/3TZTfjuh2sy1eMdx1vr8Yzm
D63l0Fg7neD0XI5/uhBW4JN0vRumLRX4bStg1IEUHLkhAI47wXoNcfRnAj+BoYZ80YtAEZDoEWuX
KDU6VgtfCDUDydpnCu5b7y1/gZ+6N0eRnEBxAYYwTal73B1XlCC/uit4JwF/w/aWVX5mVuwUkTzE
tg2Ir6Qo10GFRn9bi6q/E7NOtqIRquPazuQMm4b2271LB9Y9a0lqmdiG0jTpY1R0VMkooczt1qn2
LcAfdYj4UNwDkfEIcwtkW1vnQBgqjIdH376V+7UJE/i8bZ/A6r82A37dg3cpDzTSeps6orXnewrD
h4lNjoCUqaj4Mfasoi3ENINvk9OrmPpQctLEd3lne1yKuMH80O6vF3vmJLrAn2oEfiZF63cKVBrD
XkpDxnYBE7WapcLH1BWwaEBdMvWLn0b+jFD//mBUupdmEPANYyvKKy32ZRsTdYa6DyW6oEIJZFMl
vGM0ycV1QJPQUrID6a7rsfRm/y6JbAYT41rBGRhmrstnCdUlq5qlewEnthtZIakY1vG4PL1jO+gS
eWfGYzx33P3EwvQS6NghU/GSb7RGY9108pGbGzkiN++J3zfKAD7KIATrxqIH0h9jJhz0hh6gs8hD
WJVuxSagTop/i6zENTyhn4ozWm6OnhNK4zS0f54A/P6Uacv56CXjx2TG2XWus/aruP5w8t1OkzQa
4yk5E/f4BAj3RTmZCwoV/xemvIBto8IRzSTc2s40MAWqHf/3ia8gcz5shpEPmicZ3AaBtJfK1m4q
Ksbpf9D8l/M5597WKZWDOYBTWm8T9SnFD9LfoN9fBkNmB8XlSNa3HtxDcMEARQ+Bru7PQe+6l/KP
ekgKkwO0jKz7x/kvw+4uTx8pdfv52tKF2DhfScehc9XZ68zD5siuvw+mklyoc0QBsJU5op7uOZCT
yJXmWH+7eRD74LW7O/YZLwvYMPLpaAr2uJTOsQgDQ7Qf7Q8P3/nFuF6OWqbtw4/aJDIc15kucTFh
cxg4WgJzw5klqx06eaLrH+OsR5Ti45Pjq7fidOZ74VptccDiu44n69LrQ5UpZqd2oX+c+AV0Um+M
bFugb9e8J+3Qm+yMigzL+KygXLSAaXKxWk4PxJrwSsxxFvEApGB5tmb0bruQp+5CnhqHvJqMs3qJ
ge8mxajcN7Z67aWe/FztYW25taIFFddEg0tJDEDW8bo319l1j++N1fo071EDRro6dT2j84pL2shV
RI3vcWoq4oH8ZXdZXgQ4K8ZJHo5bjXt2RCf+8pmoWIop9JLfOL6k2h8vQ2+crBZ7+Sl1403gWPgX
t3OXXToFiifWRW7pF8lu0IKDJkgWuzvE+88sfhxjSrUNa2ZphJu3RlPn++OKxTjJQ8hceRDf2mkO
s7xbRMX1PyqGkfF7D15xuJPAn8i/GGaahZC0Az6ZfW1uCd8xz+0/ssP7i4PQ1yglm+6zEXY2rRcX
LPrHrzIhHH2iUMJvmSPCKpYNirkt0ak7I70y9Dy3jAxlV7UsYGLfNaXCHH/RXx1Qw33FW9mI4oh0
BJRnbwZtk++ESdaEON8VXjfraqc4/RZcO2nXlYMNKp77AmjetTxf4YTEkfT81d39tfnfDb6r05hg
xAwiYqrLgz1t6CnWw+Jefsk3+wm05x76GMIA5DYLTOludleiFYKgflVn88Yty/CN6J5YNI5gdP91
FrpVdtvV/A+ju3Su3yUSqAsUfr0yVjX9QYdyo0J7kSHo0V5yO+cVg86k5X+kxxY1Pdm7v8iUCbMi
I84WmLFK603eFnIKcTC9et2rQV345wA/55DDIT1Ph4cA8nFIa00+3FPJEVb+buaWkrYyukvmelg6
l1EP/HkpzsAQqnnoAMBqOL82pjDU+hU0oWdY7N3uJblsWHtL6IvXmUObGjsQomupjskNwlTTIV33
zgmAYiqOtEEIb78RLdoaPTttvP6ai1B2OUwt836WW4BBDHGbbhjaiFyexV3WixcpYCFhwU/1wHYz
R9bz3cZHn4yhe+3s4Il2Rwegqvj2NV+y/dgat0ElAvManQm9FHdeyKFALKstoaidFCmS/UMZejKS
/siqLX72pU5y0kUnF3vh5kRPOiVWszjUD/N/pN9KflqHhj6gycuL2Dc+gaVRJ8IJdwy40lC2xEze
Ng39M9WaHIf3pM6Uu8ELqqSt0LNQloEpL6/ToGb+hnUQ8ypl/E38TR2VAHSj7fPadRoN3NPj9Q/m
HeDB7Jwn27OOMBqLO8sNiA5sd32c3a45SmCDVei058jgvfLh3ZgaqW3sdZS9mK/9l5OK2LFoISUK
TApQv0qCXqP1WEZ+6dcNoqJwE8JyoLGXwlwgb+0NzYNk1BpAqFhufo2Pq4cKmQq59jsGayYNV+yI
RbhtIM9Td4w0mQv+hRN4I4/AghCj1rZv3GVT1WEXKZo8MbpwATA/X+g70QQ6r0EkRbb9FLoKIAIu
FG9nEQXvheBDF9SOQk39BpcfGHjx3zT5babHaTntJURg9ljDkOgdd7Df9+pKOC6O1Tyt3WNDFI2p
g2OuXM0h7aB+On+Qj11hNU2Vp8eYDNIxmqjtgXgzgfLvS9Q5tfcuzF7RkAxZ/cq6LQILVFECBhmk
M/jyI7tAVGafGOG31M2MAhLkL+gj2+7SUViHgOKA3/863uoQMffjpSjQuFPuSHSsTJ21K8RWqKg3
TC0ZpOw4iQ326VCWBj+WP9jNq7hNelElcnRIh3L6K5cqdzcb0WjWuSNTofCCd3rD8VmfzAB7+N06
VXjGir75FSHPoc8eLPN/Xfu2FRNIrpb2D3FzXUG+UiU/dAK7W1JrghOIlt8OsYt42KCZqhb4zXSH
68+AXf6ZoPpFpLnTYLv9/+a8B2BL4clJQPr9ilZyEl9IuAYW1gqbGrJtxxTjsfzFx96r7RNVNhHY
Nn9G+z0KI6M9B19FFLf/mh0KSo7D0/QL7GeZ7pvhYfMpZPUzKuMHxtj1eM16hMrO0IiDNd05V/5n
rSvB6qBQR5iwcYBCOxtCkj2soN9GFkxPIub8gLYS5O+9PdYchNFFLMAHJO68nHNaCLZFp1F0lSmI
8pBjD/BKwCE2mnEWFP0SIAcumsSFod0juL8yJPogSJDTfPUcmLXIoAnK6m7eAtGc7zd8PimPXGYM
GKYI2pKwiK51l543IWX22WhmFpLtbQRkMsy69kfxOKVreOrLB3T7n22vwluKhh/AWbu+jWhhyUQD
EnTWG9x5kpqhfdQIUw7aoZQt7gYdYYo9yE5H3khwIR5xVL4wgbwlxurmVfcXeBc4j5IG86I0QRF7
5+ZKwtwU+zqJEds46M5+2ygT1/E8SsWayz9MsdqwlDUsXfK6GJyZhU07qWCut3SBxKPbt8us6/pj
/FNQK86YDf2bXUl3VtvEqxivaSRP8FaWjXuZtSO/5N9Pwo5r9gpvyRGlOBMJbBgRyctXCQn7qmzo
Kx9TUmltQY4RBvsc50C3Z4h3LLUqQnGDe2VhR83fGraDsfdHO4pUu0WbMYasGY4EPh7ZgfrrSs48
v1mwWHz1iLo8mLAW6kOOrTt/LzYXcnImCyxP2Yozs/himG2ltRaIyIJgTG8IZptv4E63Pebiso0v
qdbXJqjxe0tBKmvQ29XgU4hyWVrL5Ky4dX5Z5pENncIy7aoCoKNIuY7QWfxlkZuJf10gsQ4GR3Qr
CIQj2g051TK/PKXkNm7J+uAP0UNpxob41JW/IbordgE528fpk6slmhjRwlcAYk5BlXvTFr/6mS3q
woS8OKGJwwKiEtDoeqSmuK2UvVEEfv+cpB10byP3qa/oF8sfQZu82C85ZP8eqGqYjLvX8N+igVUn
qzIteRvJopNncImBMN85MZdhlulECBLh+M7pEEgI6On5vonjaYRXyEMXmxT5SLdIYQZiNKh1aQfh
xo8OFRmCRhaGkhlA3veDmOpqT9UXGITbh41IQXaVs4LlLqsr4eVA/HtntJVEu1Y+aWSS1b+yZ+dI
aQcEyqan92tgx4d96bB3RhrlXLJ+iiDH28khpkOhvJ6r2Fi7+NsqOyqeoUD6BGz56HtlQvM9Ylpx
sXwCbrzkdjjTiLKiqBx4bw5Ya/M3GXGT2COssBihN/dhKUFXwVs9besbE1LZKRsSy7Y57GQAmKtD
IFEYN7cCsbLWEQfzvEKOKpAspaQQ4+T7zw71QKFIRqpIv1msFY5OMVwrFZxjXPa3PeAvsdFkev+C
201XPNMWoys7nqoOUiYVBAEAW0Gwok3szNNpJ8DCS8wCozK3njZr+n4P52KnB3ttrrx15GB+ry27
K4eJ7buWagpCFjGXhOnKXJKBmCmt6PJ23TvB0cURFldj/BMRYzhyLxc/VryhI8zUJA0e+dUL/Wa2
gJHwS1vXyGY+I4htP7BLpyGeQtxU2rZZPMrMqiQQmXh3bHQBRTYnUql9oSosruuTS13jSsg3kl6M
VVx0raXvBvmE15/8uZXVYvlLHlVQNIMYM5FHCeMgA0/3A7C20RdMGngUQqgQjRnvfD24OsypdcyV
sGUOQ876hrko7wMiywc1hEjiyWNJxWpcUF/KfKbgmwlQev7TBh+37cj97UT3IJotMjnGQi66A1nx
Pxvsf1MxuDXgDLYOjkC4bPJ2krFBF4+XO3LnHZfCJqeR1OYu5zeVOyfIFddjox/FjAOirFEV978x
9LvYgk6zgn+8JNqaF2h0hGQ7kQah/zzbi7m+xpH6loQFWJhOBZAi8IoibcpERSCKKCC9qIBuxniJ
aGvp7oW5cLsfATwNvVRRPQLJ7WoPKP3oUIfqzJ5Tu5CH1gLvVYf4MNY0urYvKIme4vqW7pYf3+ln
N5g6hG+U91Iz6tLH9tQOjPzJ4fePBE72XuShaAVf3CGF0BtNLBG9L/MgF01umng3OEPLNepwsvlq
sKuNgNnOw57mPaR1GUrbYh5qsotnYKXJd2EmD8FY7QGIqLJPYNGgODlHm5HbCCUcF2bsVxyM4lXo
PHMXbvLhgPMZt12ZnJAO+C2RAmVI02eLBhyjmMcjgw84GjUDpN7n25GuCzyhpBVEknZsYVV/t8Ye
eGwvYT4gNgVVfUfbSXCHKetlgTZ62h9Lm/YBHlztgSGGvVG7032YBFhLNcwpE+xYdYlxiiQirUra
pSqtlzolcPzhiXgSnRVwKSzHzqWhRzHxy6TpndkLQ4VuKphuCMXaC87quy26eM0Np0H+qo6ev7px
eMC941Bi2YnT/tsC9t+CkzyDlT1A9UflgIF3s9i3jUUhxF77j17u3cz0Av655ZZGO294b5mcqG+X
7pe6VmlCv4YOg0fOz8+o3kTu8ghYgoX6Y/dFSwmqEWd659M9j7VnZ7wShla/UJpoExd/q3YbncJP
CRq5bvILSRyarPsXuZkyiM8K6+7iJd7xdrSIi4yBj/+389m9GZ2Nr5kLgCYY2Nd7vkQ5HkgttCSD
Ygfy8OhkDyppQ/ixWPwP4sU7EtNpUGklDmBydChFVGdLDKg9ZFSiwDsft2Wn9n4IrxHGbVBOJMbi
DGN9hov02XzRBDutQ+Uhrf/Bc3JRhngASPlLy8TJgZPqCUjggmK2ET8y1sIWfJK8iC0kQ7hsRomk
BxyCZYieb1PTqVEXNONQd9hGynDbKG954TgshIKagbO1Wakirv7qRocEORcg/LcHC0Itzvl80Qu2
kAPGVdIw3eQX5Sx3F72ULgasaz8Tk4biXAnKV/i68VqOHIm7CKSsXULKj5igN8LdpPrdXddyQeMF
55wYZu2WD2AO9nn7JPkfMuoIRXa28zJbj9YKhZmxI2mKWdVXKe/6taop/G3lnz8wjdXl5e5Uzlwt
YzbcPzhW2eg+Q0mbPnPHTbPVvRTscXtDGhHPG9yr/nqNqabnvEZp3lftm5r3msyv8QdNpOW6fA1I
9pqgA2ndMFh0hOjl+yTj/LOJ97xmh9Wll3fWV4+ReVOhTH5AkXiNYoK83VdCILHE4lW1xvD5CfYm
l0kctl/aXZdPgBvQPRvAJww7dnJfmoJE7aiKI0d4PSInXJw4nWnHgihc4//CKw/OrYJr8I91O4/N
9xgCITfGhB5yuDFKix2ytoMcgBmwLSXvuypoqksHtDzHc7rVp2lDiy99K91vGc6oASEZhprhAh/4
4hy2TlGMsIYvw7+42daefrHWg7XDd00+BAS2z0VrxkdGEq9ZBSLignAq8wY2iPZs84EJzROINx4C
GtL6oAiEXnNUlKQzY8mOxff0tzHyHmM7q6spRIYTe30CUVGqmn0deO9E6Muf18nqdKjvzwQsIrPA
IL7XQaSfCgKoAOyjwFlw8mGNSbCzWGKD23Ub/JQPJbQ1Bv7CVd0Q4SOKZVLGrTOR9eknq5jGtMJp
cPv16f2PQPzKIiRM3EPQXS/N34wgZvhvAImjVrw6mKCJoeGNQCXSAMqdwb32J+i0OpfpN79qXzYM
1VWyYCZztlLWhnfxYUw5G8d+5TzzhNHa1wihkgnVDojM1DXS8EXDYW10wmn+DWmJRe3Dk5qqAlFa
6+MWkXH1FyNbRC6FmWo6xPcBImGKL/SldI+0YusywyO4V3FerjMlnT9ETAFZ4AP/digk/WOjEtLL
DHQbpUxsO60avAkWqjc+6jdLW6VXx2iDO8m0YG1xNg/9ag6N+gngBWW0JYPd8e7vmEcgVR1qQMAu
GVsTaMslQl9ZEz9UpSJCDw0FpcTS46GGLK3jkZ3uJTMIpYfRKM4Ro/TjGzVHeatNr5J9y/TFa2+n
d/SDuq/Vh8y1O7Ywr8C6q+l/+lJOnemcPjDzMXexqp1MiXSaHabJ/famkfovdyuXfUFeTQ/iMbPo
tPCWAfjJUsBhCbdym9Y1q3UDj7bBpDDX5GaR9Wzb7tyVx8YQ1beIbXGwQAO2Q3ryS00g0iMvLaNa
NQ8HNpla853KjaaPPJUgLDHjFjV3+IMcQFrxjjMz0Lf2nuhZHbsYLg+cK2on9ApAWrtXbZisfcWt
upkqpJHNKaHIrJrWG2S4V8ijzbFHhjyJSc+YVe3TGTmGYQmCayF1bciDX3chY7AtVeYLsoGmLMr1
fskrP29Jr69suZb0td3NXl5vDLm0p134vfYkKSDqMsGafgN2GKLarhr9LXPnah7dBnDqvhTZT9d4
Nmfh2azyIDRamVmcNy3olcg5N/YTlnuhKNZWNb8tBIRKNQIqU0C8KgiBK1ebae00VxskfCjCf9ux
b9OjL083DrjywApGqCyNFXFMX6HjEHOg2Oeph+kC1LT3yXv3bTz02eU+SB5p2c4lsBq4k2D5yuky
8cR1+KWWVA0mw4wyNMCl8XRaErnXjtkHMBPuuu9ZridHU+U9g77YOGAzgrsOmKuNeXIvN++tB1G8
zfbBcpSbxEHf7eSRS/veaUNkCi3pBV1eF9C2lHpACdKvuVTMtRgBagGaLE9Iyf50zJdvdlBA4GMT
xuWrXGUY7L3oQOP9f6DJrorTBaje6DVe6oOvcFA+Mn+Pp2MNkmfVBLc/nw+SsfjkSJgCQL+Oqa2v
Ky3rCtrIN8gsGKiDG7Z4tbTC3B33WomrtiWrjEI9wTe1YFrINkrjstrHdSjILBKI4x98UZ6EOjPa
uBBDJHJ1UAdk2myjWOF8tzboNMSNa8B0qGvyiUNn+a4oPh9favkywZjwGUpIdbVtnvMdYANp3udB
K9oebJZBJ3MyNkl4cP7agpwEfar3RVedZHYHW6vPr93oea2ifW+XbX/b89jkA+TXZb4WMjN7UC8+
PAAFDbbuy5g9IdQpiA9W/Zx3lVthcwWXN1zRpLijfpweuJvLHbaUYIBbIkag42LBFj2CSvMIZnnM
xWXsi+U5wb2Y426opk5h6mGAlacKGXWF98maMm2+QucUtqnd0IY4W4wBJIqwjN7MXvgjiFxeIdqN
VrMsNn8e9pZZf25GyoVzMJeGwDKvAz5Ye1VB3/mRrQ0z/MQaNrkkVcDT9E7CNvSLIrDMHqdAPWDs
YPZCJfg+iUhutnN2x9CilBl6enVWooBJTd9/4k3y+hMPxzd03cVi3zLMs2KlV3h556qT+nugIjcm
akLl4lY2BDICN9VHXb2p67wSZR94+Iphro+ZTRgFpgs54LF2uAFwZTXRWlBYnO+uv2qM/9qQZ7Fr
UcFvUWrle+xn3w+ir91pj/CzLYTRuL2zNnUAB4U6P7hM5PdDXbveNoyqsFdNrBTuEt6pgzR+0ZTw
e/t9Cc8XuC0P8XLntNyGJ0UATQeh0/saaTk8wDiTlaeKLALT+MoXWrpzbWNpiIB77drymNmBhv+R
mBZqyN4z2hanDFez4TnSwo7U2UIdVROT2n5EUbA/ynOfpKiF/tTiTCRkexlZz5otfxS+V7D0M4gq
g8SGIgS7JFL4o+MsE9Yylm1BZwjE+t/A4/N2rcTQigDElkNqXxuapDYkBjp7NdysRqTs0JAoSUt7
7sNSc7bD4m2jdL4G9FfzuNy02ZvyKx8bC7vABRknLjwwi6ov2KuAJNMSp3nqJrrd3eSf5ti65Utt
ZChYo8qneD64NGYNtGGHSxu+uH9ZlRFhdrlIury5DiJuAwfj6Bppd9LkaMrYwn8CWpnCnn7k/sXm
QVqZ8J3Pci+JDfE2d8/tP8SR3soYjP0VB404NyzSZGSquxh/PWq3n2PjCdd8qOqCAUymSizIqemY
jbX0d9KKjBZ59lxJxCezt6rMsqjMmrp2k9iqCp7ET5keEUaBAuhSp/VcWkOenCE6E5Hi9cVEFOe+
OZVzY9Co0QaQq9v8e6HndzdCYZEzZivGyydfHZG+4z1hWbsOiEbyMZ6cza8e6w1gz38VXe24bvmk
C/B0lJU+tkreZBhpzOCv5hDTUHm6Utyct4RaohLQ+BKPLr/Xs9HjjE+BXDvXujsjh4XGINZ1tVda
FXvZDYeaOjmSKmKb17W35vz/IepSM5Fq2bZk41okGzUv3ET1IUlj83c2csIAQN+OwtsXC2UppYJ0
HIHRESMu+zHfudDlJOuex1CfJyfFGWs1CNs4ruiYfFUwIpdnQrfQQvmwxNaL0uhAFNOrrltksqqi
Dvh+bJXNJlXsONgE1C9JkogePfpYZ4sQ1Y56BqOha9Uk+71Af7/g8d5dvwTBDbX6ghY0Zm5jdViZ
e4xP2T9Veaohvv3rkHQFcNnoXHpFgLBYPOQkfZao6DMNSaHY3wOEKIfd7Ds8csJuNZUsJBgefo1r
Uv1RtuZyGX1P6EnF3uJTv0H8uNUczrsie763n32fOynua6IjJvyI/Lwfu1ILjEOEOTxwLfpz24Qn
k0DnQn1IIXOhgM6yFB8scbp19lnSrvTSCZbOdyUGVMxI6c0l6ZnZZIWwhSbiq/MoFCgKDfrZDfra
Exd+QOX2v37w6j4xrC5K8cNRxnWOmGFmQ7KlLhrUTwBfTeY5wi7cl172+RamkTOBFbQvD0rJnvHB
NGvBVIf2PeliYgZVKmnh0p8OavQmx5/qt+20fNmnvMnIKVbhxcH6OhvUPakmkfzGEF2JKwK/xAdx
DATIe2zxCEFxl+X88vDH61pH2Tk6y3fIhcayQMRiWbODVGSB8ZGQLpycczeRt80Q1HD2bJaQlJX+
4Nl62c6CoBMwiTvozPFPc2uqM1JsnIpSbbuHPsQpiXj5dUKBAtcpKkMBy1VGTgk+Xp4jZLQesJro
AF5/+KkBtjg4+nHM5f42XckBiU4QGAe1bnOlET/iJepL7Ul/Cky+SC/Bu3uqvgmWbQMHw4bKqW1P
naiddqmlJafUDwOdPL1RSk+AhJHlSnRGiFUtEN9JzEaEORrIwmBu9oBxYjLl7FgV9rCneG9I3y1J
BLWEzjiIgOZVO0NLZjlIw+yRnWZqDeSMCpM3QfVsRdbbxOua03p5zlV8BtXv0ynIov7BS1ARgZq0
2mklfJi3zaOO0gyEk5qc937ueEWtk1WtjsWjrurJoV0o3jkE0zmWNHCpiwLGzHvLhzOhB5ND5SvV
htW9Y1/6CjdOC07a/raFCA7QIZzdTYkuDZ/sJ6UMg15e4p8iWZvgcxlDIv8R3nLbeHQNw4ZodxFI
fDynOAj5LfVLkP9T0HbB0GkwVvcuVcigCfs+q3TGXpvSTK7vcjoEAcGxD2xhnrkc1lik03vHJSTZ
TbwWXVB0AFaSvBRY60gFXW6s1ctSKbHd6PxmZOUW7+wMsMyICtLBSwvCJJAsurjR5Qn9WF/fPzw6
75g2GGYfNktj+DqQFjYYpZcPm2WPk9gvY3f0v3u6/cQPWbZfM9FiV/fhwIuBh5f6cVctYLyBz/od
1XCyyISuM3BgtSX0a+yn/grVgvb4r9NenvMiqTETOglHFLyfPRcxm25XeNeIjc2iUEN4v1ZPssQf
mIE3VVF+C57OZ1HTvLi4072PUO7l3zARfUznUE43mQygm5dHthqxoK6OP6fmhOEBahEdDDUr8V27
YOnNZUXvkVrS0zUhy1LnM1t22ND5MZe5i6IunhnNTPuvNBf0Nmeo5BmhiBz0acmDhhpZa88eFkfF
8IMqQKiFEaa6eVa0jzExMgjdJTFyiia6P0iWCPIlqMHifJDYpyI+5rFuDvN5QYDGkVahZZFD961W
fXBZYXkd+v9IsSBSpV9Nx7T4s2tbmVYbVtHZgsIEL1agTia5WxCuHhjCME/DuPk6pmXEk7kh8Xzl
QLUZNdsqrWq0MsLEUWeYbbZQuIEdt4BAB+EOGiAs/f8DnLzPhAR/4cJaoLn2oR46kOVJxLtYsGWz
iU3EyH+b8yqVSBzPC5xOCbe+zplhw3o9aBvmJ/X95R+a7LCWHriiXaNRsLwvH72o0r0B3NicZHwD
wathZXle3PGwKPiVIaRDAPI2/wh4XjWjvVdmsqf2h4hh9kh5+MECL5Jq4KZsJYTdoDsqtCHUqtDk
shdlwRjJwpo8fRhjZV5xEa5siiTdnria4qENWaN+U/F4+Q1FMSso/tSrmw9GU3vGzNP1tZy+Npe2
YWRa0fM9dp7cyRXkHUt6sWSb9FzbyVvAriRhpdOT3+4tTIAbxA79CYR1yuRoGDotsd85OGhl84EY
dp6Z6dYoL9GIXf66Ncdv9z/rbDGk06Vi1wZH2uEtgSpeLB4kACyzi6moS783gQ3lfm75MxJUVHOC
ic27ofR+6AeAkdMa+CTZtY6A1CQFRiciJxL+Q/6HquA6uH7GynJa6kFcTCgWrA7V07tj7DrFGwRx
LnfN+HYT7HvltcE7PVLfylUWuubxsD/tH3HO4ETu40/oAOYwVw7oo1lLJqL/b2x0NESotfhyIgIb
+pM30/PERdP3a18aoxQSRnFzZksR2DXxRw1fThqerhEEsaekv4OQ8r9kqUDR0Th+0h1il2Csgrtl
wPIHcdLt9KXaM6Q6zGhX2iuZuoDr/8cVl7XzcwAASbR74kZXSn0Q6tp15IXyACdseHJrIhTgX37s
hx5Lbd6q2IJAfT3x1flLs1+L4T2e68TS3OdfdrEEQsm0LxBzDsK3jx3PYRA4A7ljiW5INE1jLSAK
OAhlIdc7TkCbCuXhBzIGLEf9iRPc0oEOOs2eCjDxhe1u/7bC1zBmhdLJjsHyUsMDAARd2uFP10mj
ZMy37EweUvxuoGPkUti/tToMn7RSXZSMZZQscSNIGypOvaQl63boLDn3qld6139XcseY4UejSvpr
3/ZPGXkbMUJYLhcmQjgKPeFtGgL+4G91N6rd+6bw+wib9w22WHRIjTMd4edkoipjl4XyPJAe51v7
0KyJizejpBClaQFJhwOBDOJNusIV/uyeeyTaL1+XMOCkcz8ZDur0jGOKbBS0x5A+ILBGD7Rz/qd4
8T+Sx95q0M46CaZrfPjrpuMFqS84Qj+Q7oBJthLmWq3L930KqmPseIz0+BajLQyVT1+KITL1PWUx
LrjwDK1xF/SIOkc3BkZf8mzW0CWlavjxBPX17cb8tXncD8MZCwqPe+0gSkK7AX9OUqY0DPBZTAWB
SB/vDziYYCoyiKwMn62RTUYZowU/l+w+AvTHSuQ5hmg3Lu9pM3pJK/qtxR1IJDVpfmYc+3bkhK/s
kD7d0X/gmgQ7JowL5e6KJgY4Y+5UBsmtb+c8Sd4NiNinksycWrs95qPUN1UyGXCmMwch+jac4A+I
KxUAHj1UP3N3U1iizhdiorbONp++aQT51IRM0YldAi2a61zHeYaClo3e1LRyuqUm/qAT4hEAOxp+
rD+vDSOchrQOunWCMiNQvki2BJm0bY2jBZzGcFeb+yU0RvjUpS0xzLCtiWhDaKf4KZ64t/KdhNa+
ip0VdZVWCRLDwu9fPr+lXUNS0CmK0r6VLukzN/a+0LBQooGY+8SCcmN1/TFenw/SVMb70Ex0fyqz
EUHXwC6yhra2GUTpbserbfg9IaaZS2H0KGrEjVfP2MwMwDcYdazTt6Yndko0gxdm6P4HnejFMMwA
f0hyJr2C03MsBVg/gBgsUKadXVhFtwzeAfiXc0Lytu7sUB5Yyoy0h7EvSWeA5bwZwhN0x/2y8xQ5
PxJKHLF21MyO1dFTq16XGve07aIDe+psghrTj61feMuwFfaOjTCkcqTGHUUCR70hqy4H4f36HRU7
+0zWgVvU+ZHp7NatwDM33OMocZqz9qlR9frz1tHyi+VumlsXlFwBU2MhslqfnC2FU6IzwEepj6kG
izVZBzJ7XPcKn+nQBDhcCShIBpnZ7Ry8oxl3CqMZv7eWLYnDk2xQcuK87vUqQ7xTUWQqEB0V7W2S
PP55ruN1LNC0XHYxHcDYD59+RGW7j1avTqWr2YbJoRR1qzllJwCX/kJzy6ykA0PNUz5e8FjPH/fs
+fVaRygkk42qub5/8soAshCSOHSR9kLCZXzCMO6t7b8U610dH3h1yHJYTIYROfN/GOZyetEsXqX3
oVUXoWrzWWl5bdN1Ykxg+bDwXRZUqjPk8J8e126UIrFJjGOnqJ5tbbHQadcDC03j9bydm7405QsI
HN02GWb4DRLkCgC1OI9p9KMz1U7HPGIKaBI9esslcyRUhzTNeQOaZ1XHl5jNj88X4ekOVkAuNe/6
4gvemFGD7pLDpOtCKes9SGwJlE5j0471blpC9tKeBQNiXyXETC1fxs+glvFCPsUIWHnwCqO65t/t
kEgrkzo9NYPxbQTzPd1u5BzyhMcTZVE54+Zrv7TwMqFyM1EoVACckwLSCcsqiIqmbgWUlqYsahJ7
Bdz+yL/DA6xOhfz8QI6slV/rxgoE5qGlGkzsnL0IVJmgAhnRzIeE9mI+EWO3NVIY36nqD35fhp5I
tLu/laUpoVn+FdRiyTzDcxug0mjfY48kH0RUJbsf0D4MdBOG32Wy6vPw/zsmV7nlRlGe0n2pcveC
/GXa+2/P+4KUKgP8LMhv6G2BWyk94pGIqYNtHfxgqO5bzdUKYdyamm2CzZ5jgqJlIVHcubVGoSjN
usEIi+HfppAXt84qiBNJmSlTcE8NYXNwhsLTeRj4bF3NyFFvBsZtZjdBJoo4mK9oeXY/nk1/PpbO
1ekfLuCrqVIdnWSYgItQsoq0b6l0s2evLALJYuwCYCgHMRvh6k0uNBNKFOdV+YcjfCsAeVezQt5d
fRiolacNPMLptx1hbp0uCAkWTr3Kzpw2yDphZJxzRo3XkZX7PJly5xUns9QY/5XPk8ks/XO98QZr
GF9rX25Hq8qfDcOBHtgQPbTK3BaLe+JrXMLb5XRFkcTGUhqK0mczxmrzahrZB33xb5DpU3Q+7VRQ
3fSRqh7XwLtHy5qvFa86gDB01YbpGCheSVcD9KO5AHYmOy5I5p9tKGXbBH58PVhGIOUE9dueNPpl
mihMH1tIr24ahnz4GSrp6arnfWasaU1TxwhD4DHImD7+xyL1Xr03kvRz+c/+ddZggE/seHF3WS0b
z8QOev5H6ZLOl52NKmEH2buklcTdVW1bqJQ05Enk1xKQwquWu9JWJtf44uPPTprcM+uqt2gdvNY+
ZK6WyOhU4I4ht6ajfbsKIcCckFix4h9ivPFWEmhWa7YzMgu/TI+icEvAxLyhEa27wI/hTHAL0xOA
swABUz4dEy7yILu/fbjzi1BaiOeTYBPRz5six4xKmZZxLpl2XBAWNopjkbhXE65QBsBobUnabZQM
y3GMQuxs72Geo0uq8VAmK+tCpx+fgYqB8gDE0arUcDKVCUeGjPcoNMWz6joiBnFYrntrDlqdxZf4
d3Fa9nNYdKNKn/4DalGi2p3TFnG9iISUrAjzqp0rcECUgshgFehHgJDy3NGs+U28WLvYFwEhV0OD
bvNz0H1MymNXu47DaP4GkXry71QDbaBu8Uv7ZB9JJrlMnmE610ki6kMewGP7H+soNMcafdp7HrwT
7bLKEseTUNo5BxPeNODrTnbJlL8MUL1GS6ZCeFvbG8b+m0BR63P/F6vG58kMPtIrg02tk8MjFxLU
w3x6Clc/yTjF4rL0Lo36AtqoFQbA7W574sD1lW7rOFbPl3teMEoB428IT4pSswfN7GlQJsaVzuaM
TTLnZ3kLsQ5VVkk1f76/wW33uYXcNsWtn23wiOkmcgNHa9tnLGRVvZ+STp9F5Ys17CqMjZL99v0Y
ba+BPV+/HP4GHSdLFnnAWgRe3bTPGl/hR0Kf4ABv4fNWKqIrxceRElMY7Hv6dTilEgqybwFj2zDD
ZtJDHzWJAi5nEpZ5laFrfhQbQNOkzYze8cSw5Xj4GygNDXRcpwzLnBKlld3/hhu7lS7j+tqLZtct
x7JiTahaZ8ngH7ntbUr9A3xhlN20JHlxUa/ewr5+p/n/ROYRrc2ZOLA4QI9qrk653KmKOTLTzkCv
69Aj2xF0z2wPvY1ZmLsU1oN2TL7E4g2sLGDQO0tqyTznMimKhdni5CP6GUxWGButmfEXfuSyQFNu
esFrf+PIagrrVZ2I3p8Wjof1IN651rTo19T945i5cGp7eJXaXcsax/tgrb7GBcsR70afRyf/+uxt
JJkbgYG6H251HqVOLwrzTyRR78ACH/TjoSKU383JA4QN7+zjS72f0AYdHNDtxYEKk7X5Wjg5ozFR
Xs5klYI7F4sQnRjxtSj0pAUJWx+uHeA3PHoQG0uJeYiyAmBpPxqZZ9sA5UVNH9ixBAe0ecZP0tx4
l9a89pX0PzX/l6Y+CTTDPplBSmpuFofBGnaaojCc8gvBSFlNpG8lX2SS9BNJJG87gtflphR6YMdr
PSTuVPCVID6t3qSylUDax6Mjp57fJOlP9pe9k2daDlHmgJvGJINAEsHF/+cMX4l5O0HLhHxffGqL
i88eeigtXdvrCCdrMtP0X8T78+7uYQHkye27APUr5VHzX3mpYAlFS+rIm0Y4fCE/75EcdpLzstxj
LrhiaBiNSaOBAgkbH3OFDVR4zgOBe0k+aQB+pRYKBRYENSHKi136Vo+5h2lXVHG7Wp2n6LjUIpeo
JCwFO70Lmagn2zEsJ7ndYMHYamGoXkYrjeUTYU0oO2C/rkdMwq1X6U/aKLJ7DNQ8N1hF9I6YxLUA
1Dca6KEaUdnp2KxlO6uJxCzMQgnz6361yQn/FR7v5ThyOPT6jEh9xT2SgsbhEEnttB48GnvgBa+9
dgk/QTW0XPOGt8Yu5gMCKYlVW/aTT1NYKLt5gZ2XSDLO2OybBvnemk9Nh5vejnqnGCevREGZyUvv
uzZvAXcALhY0dnzkqubaIXr9UjxdtuZYNUkp2qUKyZytPYrAuu0eaAqsqCfIMkvmLDKAWQB+g6xT
kGeSEtTtZAmvw2I6UIvRVKfH11ZmqgYOQx7RYh3EiZDaq+eethuMhJSaNmbYhjCo75AiGinDP2+d
eQPAJw4IofPR5dgnyS1lRJSmO//V4z8F4vjkcVO+BNlZrjm2q9xoL0sDu3qTmNf89e+HUYQoj5og
o8Zc6br6HdIvhk+WHVZJtXzlathyDPhueRHrmMsGsQtlVKQiYq+xZKLscFzQxN1nVmhO1mQTROcA
AKDn1mHH333c8xGeBoaHdrFw/0ez33VdmCAnNkf8w2LCqH5qsSsxs7L6ITKkK9SMhydsKI67Tfqy
Y0Sj4OEchpiwlEAr/PvLxG8X5yvNgQx/ImFtpHaSnRBb8NrlMLL5MN301wKDYpMVbRs5YqoPX58u
JIEfTdEWvVzl2W06VE8he+G/bbGI8VfNJU9mQ4uGLZBmOIyNU0vPHv/6TLr7As2bH+7vE+2c5Fmy
a3lpquqTCWCZLDzfF5GWwKaV18nOtqQpKNm6vghvSGEg/byYLbRK+FtpRv4huPZ2hmhXEnxtxeps
Q70xtlYLnqUf+09NhA+928xLHnKv+whiN9fbGsfQ6uxP+SpyDOhh4a55rOWOQi06leoZfqpqVm0d
5/aB8ahsRP0UJ1qRMp6BG5oyczCpctrd6LSXIUHuiEPpTxcDYjVlk/cWFflFMwY6PWxq5gQlpSgP
lBzcWYbVQ1edyMpN0RX5jkNq6eHmftuAfD2AoAvBcOVCbCS7RmNX/59DB5XelXf9iGe/ub34/LpD
ET6CwqfkTwIvFJNUo7yNj2XX9SOgGVR3H6fZ473/m27SN339E+17PKWfxzjtSJffHKwvKsts03BG
PSlpdQOc+ivxo0tg9Pr499ah/tb4LlaK+lbWJOHE539gh8sU5TKZUI2Oeca1iX3gYfqTCxBLzKjY
w7EMUOXkyJAFybGOxNkTHmgeyvIa/efcuiS/ZCR/aql2CDVtl6pa4oAqiZbisuhd+SI7Q5E+hzlT
wbOlQRo4jxE/+lrA2YM9IqSpQeELHn7ijo+8Wyd6bdCnGJNh0itMuLjDIjxLo0W8uPpKjN0+yVe9
sjysBjOtL75wK2V3kRbmYxmh62xXXOxJfJnhGuUbIPwCmwtVNT1by2kTZR3mOHUR7hWMgrWdM8GH
cJG3LQiqxS5mZ5QLu8Zgh6IO21TqaYxWsfZfq4BQnxB4AmCAF2Okg8BwY51XF/j4US+Uzl0wQajJ
M0YJaSgEZ/WoVwubP/RWPmFilpqlBiPiYfkRDmVNfyuwn95TwlkU51AgqYSjdHPFBrcl3jHk/tT+
yAy9it7pRS9ZL+CAtOa1xiPnH2cDmDahB0P7y6Vdl6GLhwQpV3hDukHNORiRM+6+KA9BdOlOhjLI
TeTFEaPewA44ytYsmh6YepyNin6Yn6iB1fO04n2qVRwTgB+CoOIMD7VLWzofPyl+6vYrk5L3e1o0
YNYZJpl8gf0RIWSY2QmzP0mytYlgCgawL4noKAmKQZQ8aYvNIm+rX3C6Iiz5JkymnuH+bWDnV5wC
vYPRXmX5Q/EmPZFT/NvnbeOsfaEcrVv9Ju6uT95VlWnIbtOSV4/+e8n1Eb1i5+e77wB7D6HkYBXY
dDofXjfAq5nRKq8unmDY2NuJaAI6KJeXp1PEfcqF52qKpf10sa5OfhohvPf89HD3t9e8lCyAFeQN
aBdlEAoncx/AD/LyUhQOZVPnwIT+Piv036Vn0oGW0sqJPbtmFILydGUETb/ajgojDVdVZ/OoIAFJ
vpnf55d1IfnBR1J5MU86C2NvflO5yA4BztKzL91mhigaQgwRaGJlNZIxry9MWC1FLKSrQjIuMw8r
mbu8etiFlF57DwkaYqhuctEHDayOOw4HVp3njapLmDlFHYFf8gs2y6oB3oqebThkM9QB6lOg6nzg
hVgzjZh/Et6BGpOx0NaKDPmOFhZtQsMw6Abdl9nryuIYY2Bp1HaCs6HygvqFXNOtk6I554yjYzUn
TyBiXaaBE8YsgQ5M8h1zrrVp8Eyc6nl8o5u+KJoADEJ365atVQYQc5VHrECWNfm4xKouagC234b2
miaEsy/YghT1kPP4hFrmPd//DJu2au6sy/czk0nAhMcHbCecd2C51wGB9/0e9I+fQCImeFhW5w/m
MS9dmorhfZZe37KrPZfTzMsVpqxprGr+10GGLC9OCzc94gP37w7NkQdo3ELy1Y/76u1J5eINC8AQ
0SJ3QVrbOPqGUF7oJSd/P322ISfkwMGWikKvGVk2QRuJAWS3tGJTPCD8LWbzR4o9811gjq+22WQl
4SKFT45C5Qh4ZiqcEghzyqHbcyoUqg0Ks/zIQhQjAr9IAfxYbbgAj3REwtjvsBAWaS+pFLHcE1Ip
+U5apcZ28sX+n7oZ5y+tYuRudCKPV9lxIU/2meKs293GrZyi7sZ8UFpD8XvJECzzlBeLwt/ZsUtO
kuJ4NWj+nVs1xOMMfZSLeieIZiEE1cRqJisHgNGsmzqfGuPIoCrcru1RKdZwW+HFiP9oL4mddDpO
bwR44yU+Pzb+2kxQc27IkdSiqzyfg+G7elraJyVX9xQeGK19KnwrhSNohCaZbSCOktGX0bA+AmOj
DHYPw3Ke0QZd7l3t8LSR5mpbuzIYXTaF6L1Uqd2YI6cQ0IiwnPa85JovfddQHgS2ecauCd9srKps
6YTfrc3qCgwi2Oua+niNMsdExkYN+AUESRu1AijklGSWgXTX6bCA8XnFCjbuW3esV6We+T4guU/u
N8SvhvPr1GE1o+kh/inNL/3V27eUdjro+N2dVkkhdZNWSNNbz2qHPEYiO3m/KsVJKnILI2CcQpBc
hjs4CJzrOZ7ChY0DUlXkSyx+w0cMe6D8fc+7f0KHPC/aX97QSnQcHWYKDBrNICwmMihLPvtUNnD5
a0FA2v7f1BBjBJ5BZA4l5ho6r1Q88xXoLZ9zYwC/327sLQ1eIzkCPy8qUFM4hbEvUkYLv7h46fsW
JaXLDq8dv8olThtRKatSleWPx4gJ760XFk2Bj3qfkI3OZ8W5PEgLjF9mSlcmMXURJH54kF9JfBiX
YYho41nvytXCQf++j34yR9Z05m6vsKT1EmTO2W7MUDAoaTjEB8pX0Mhc29jQqqRGKOk/7crxhp2m
WHnh+9UOmpwu4Jt7/HLBnw8yNPj5fBcppZU/pYpDs1N0MW6w2Afau0wPOxATXe/wN/Yt/akasBGV
/4AvQT/v4geTA0pw61dW/HBuDNthiuG2X14h56gJ86bfSvwX/GYhLfhRxYdlF/TU5vXrIcvJ57/V
SoP/oqvP2mjXM9Xqy4ijKI2+ng1lf4X1TEMhK6RY+5Sz0pSSKfXScfeDzbES//8uCQPaRf2m2aHY
qmDk0HyfWZ7bGGno33hIqdv6K1g0lpOabClFFJ2Of4DyQ8L5RaW5h9IAi61XE20uRvXIFzmbUjja
GwMlBsWqWA+TZ1+qxeqyaQ/afayCY4OGBUTBH53fuXEDTooO+Ekgpqjt9Dj4C4UmeNu4ejHNbbQK
lDsox+mFVYNMnYXYY6b/Fw8Vn7/SvmL/nA62mUFCBQnn5xz0cdJPXjvKLlLVAIuxph5aH5tYTGwG
5fLgtWLebt1DerEGD1TCN8vzEUC5jQW2P9YNcRtxzNWvHF/XBm6Ft30kq/8PrNUIY8Vyuy+VZBlY
cj1K1hSs5D0Cq6OLbyMwSwPjHcpff+jw9bqP79TTKlTvn4eiu2tkERN0a9QW9zyHFrfre058XMM0
yK0/77fR0Qn3IvximuqcZWlVcbRytdqlv+W0KMcIXDVMnHw05xONtyopqa+wV0S12tZ9adrXiWxQ
LgvaLOHJ3SXWR+ticui8xYefIsAdbDZgpCdX6zV404JV1ZRGN36oc5LqrOfw6sn6wHjH9qEvYCVf
3RNAlGgCMTZpAd9dQGbz3DqAWAZfgqT+jjDix3xsVNkg/Jj42p9Ql+aSNXwKMzVxirrgO+DURB9s
oojpduu/8Iq/4gjclQeQbCpyW9bNcOj5V4EaykAKLfPiNGJoXIJkfzh9wm7VkhPLR9IxLkmbOGu7
cosLYYKkxQ6lu+jgv6lsSBWtvFwqlV3b7PQtpVYF/Q//Ig3OehH8ZGnMMeCqJISFBn7aRq6GKKPF
OMqZc7j1S1Hdf1GFKhEvsjKtO/Vq3hhb2i6Lz3MTDbmJTj9kErpEfhhZyy/VqmCo95setc2Hl2eL
RXY4g+Am8BWkOT8OTUspdTCZ+x3D2LlvUIWNik0fP2DwLkVBh9Rk9kL2b36krubzzVPB2zITHvO5
uoO0Eu9+mJneVE49gd4DnrU2y7lBK9yNvsGN27J1qK0Wc2vSSNlv3jw7E7gI5CmK3BcYhbXJ/T6x
XtgBQ7L+3wEaZW6N9s1wsv0tuih9OYSomscLXRXtHL/2Pj+dc/Sd7NLTVWEm109iLQSRW/RLIpdN
Axc+Fsv9gh38j6sfoa+c8DPdYXkrFbbN54pzeFAIKJj/0hZP1OZNcBXGjtTWp4RzM+k2n8/mo88a
hu7D8ap4NFgO4xGCgeaGXoMW4V87AfdgrfR9+xbkEC/wE/iCtGx19e8peLyECwWQBSKymaFziHeR
UnW9Qr1eLNYBHXHGBPo+t6Qei3VOOXUbHJGE/uqC3Tvmd8KS+iHZXpS7G5nVFX77gjcEyMh2RUUm
j8EG0N8wcABFHni0dAKlfox7uOEkkW7rvC7Y6QW5LDPLWLs3u0N2w1uWIKI1Z9vvlQbSlUYl9AzY
un7REGE0jGXb6NvTAtZ8nkPN2XJq/K7ekTf3jqMP2NWmXggbsBCT+XKbkZmpNo/Q88mhn39WzWI7
lvS1W00KU3k6QjX6k/pSbbIt0fXZIj8om7TaZtsoLP9Et28UCMUSqe/DcC784ETF4QRzZBC71r62
y45FkAxyTLjLZalFd+MY+a5E/k4b+Qmsls493uFn4Q9U7n6IhTiv/Rte5l1qsci8IUf71IP3NBVg
QkOP+VazQqIMXifyBk0OwoBnZ4ilnGx0I38yKi5iXuPvjMpIXbvBLNSoK/CCl/V1X4bMsYL2avYq
vIVkWD//uEvrRdoMbnneJ9bnQqsbLlvryFpb26oCmjGqeWrmmpdktraDAnf/FUxOWkfFQmZQGwhZ
UiBv7sQxf7cOww5JP2Lj6sdgTbv6G9NnIXx2xMDT+fprgbA7/0OMKP5Tc78ap/urUrHWHLfc5lc8
hgaV6jKZ0aRIF0UvziV9JSvKLL9R+cql8XjuZ13aqGQiTF9h+K3jf8pIvDQhzDkt400JvxNC2hnl
e/ZEK9HiB4Oy63fIqSrs3cA7DCuiCH7IP/vunR/WL+GQuYNGIKU6Y9LALifrGF0CA6UhjsVjRUuq
u3uT81FMtArKXw7Ng+mIOMonltQanI0EtyhCBSExFKvJLXKuwiv2jz9I8oBNTqUtXD7RoLkuaNVy
Gz+9NyLKmZxQFc0AlYYvCBEI/dqmka5nKwpntwB0hVGipX4yOS+5BrJmhIe9bAsSFHd3mMs65gSU
2PSCfBk/UwbQGv7ZHI7ToVS2fX35fpoW5WsRiIkb5Vo/2OBPUVchLGfCb6VDK8b0/yOTzsoBq6ef
bpDhOApVqyRYNsGIkhW+Lvh4h3SZ89bhZXo/Mvh1fc4xFC66vDNyG86QAtMOlzUt+WDdF7Z8ZsC5
JVzQEG6Qu9UZCrDIo9XHdvsfxBI1Mz1q0oA9MvnrWO7q7ogXmWE/lRHSy4QyQ8nc3pG5fsT0f+0q
yLG9iS4M+3vEzQZiC7BrM0BJ6YoV03yHGZMlCLXabQVBoMV2sCVJ79cGd2932V5lPSQNYnZT/UAw
FtYOe/TmUSuM7DXvnNKPMP/rUprLHboEIp/opapHfO30iZF/7qTx1RX1BCuIUP0XoUpy0oAptYlb
u44sq0TPRhM+Y4VhBzDQ6DXbhjVpPZFiBbyd4rU0al4P5oaUumG3HrnSOO2MDieHDvlXvKLbPnsQ
ANi62rYpAWiJfvSmIGGuLNzFPwEMZZX45MfZgE3rc2k1nFO/xAD1Kc1vdJQpj1U7DofgCgJX2CAN
3i+C5AbTe8m/xK/1sTdkUhvRijlFStKQLb6OSlVI/jjKWHQwrahhWDeU/1hVDaA2L/CLdrfprzp7
WuOK0swpH1V3ThWvQwxyN4HTgw4BVEsANKrDMFKF6+iCIgRpzYFnM7i0+1I7ZvRLnCnRT0HjPof9
dDcU/zH4/9tubWQBkhaSp3UY/jrKO2dtFQcdghdCkYt0aFd4HD64YUY9LImtSy1XQLixekl5I7jg
qEGqyLMPEskfksopmOBS56Xu5zdSzaEcjmJNif0S9FMnHmivtK4fvn5ZbpeUBxutBrQktWIfMasl
G4NZxnXlmgi9n+2OeQr2jB6Sawyzg3JD+a4AEoZTOOBE46y7bL2tqYO4hd5iAMsl13bDJl+Y2t1Y
tckkH0UJHiCbHV8YqhJM73QCrXU+43MpAp7Cx4R5Uo/PW9LTYF2RdMuaXi6aF9ToWmX5EGAHxf1b
04h0lyi4zdzgEjtcw/5OurqKoQ0yxEKkXsXpSxJ9cAHbxWGCwrBy8voyEoq14GM8+TYGkP7NG87d
RXACuskjZga078M7oM6DBi5WX0ajQYcVffy9Sav98iRfQoXdEiRy0n6h4V9z1yyb9gwKZlWmx2ic
kxs/zpi6a9t/oXZ/A2dQDx0TSugj+mhwvTF/DlFVhU6ls6MlPrlcXNjiKcSZ/kVQbFXbvg3zEhMG
YfeQkBp9TL+cTQotuNFRXlqmu/7eeHROKoKvDm2k3D0soW6LRYsjvzBu4674AKJkkepnCcFC11IP
4/J1rbnc80KVJ6jxa6+CS86RSwVYkwJCXNa5ZN08mMMspd+AARFBVRKJ715ZF0EWGDCPFFhyB5iT
Owt7SlQ1gKvANpZ+ZIGIHt3vRT3q8Y3o9gqKRopIgh5zmZEW7oEXFoQx7eD0QxV2AgUVLez3yEFs
xNS3O9LHe7t5hZVJYpvlT1LDT5KOrKlhoJqY5KrPiPCM0v4uzLKj1x72dF3QEUtYI9zG1aDZcRmg
w8zn+8QijsJ78TjEG1bI7gKdu00yt00dp7VSPXL/999+SG2Efkmc8TKd7WzYL5fcnIJxslKkol6g
mufW+vh9cXEqJLxVHOunTUl48OiBYWh67xk1Xo/q76aSSGNsvXsLiKJ0dUyW8cz7ZlnkHb9JGpXI
VMy/g7amSVnySFWB0u2ObWb8kbjKk108jGjJXH9lxe9GiQAyiFelDdWFyTooC+oK6s8I/qydFOUH
3/4xuRpvgRJPsuVaGRNaa9uHKGSCs60Q1iG5OBc0B6pplN5nVuuFS5VAoOZEhn0IbKnvvdCzLHyi
HU2JYHzMzgZucImnLPJVBz980vhGIMwVSDbRonA8CgN3Z9hZkTVH8KtYhSGLATvdrKwDaCBHqkl0
59ONhNfKqcL/842cdxmgj94yOFnZ2fMKT/wTnokjwt+oa6oOmBX/TnO6eTjsPvKK3x/yDpihw5vy
t73LHCdP+W0aSMku1Arjd7eEtvsOA6gJZM+J0PcunSbGW5x0ruI6b7zhZVlwYpvMX5oG29LwTdRv
rlbMp05pQIENQiEcLwbxH+a5fVbF3rTWvCHEtEjdgLTxaLgUcaMtqENGXluScOeizBEc81nVd4rL
KBiy/6TLDSlOazsWA6KvNBdtfxXQMDEHPvSTRSizwhegSs4smytkruFfLYCKwM8Z0X/oQQb3kgm2
O2vWYVSP1J8DkYjCOESpoz6tOL3faulzmqa++LTtEF5lbYdxRNcnIwSDortrSgk1VllnE30DTuzV
vZZIoxbuysYlGGSscgMlSym24rfMxaKwQLRIMIqROVX8QcsgkTYmYlQrzUWrWH57dwbkL8lgtDov
9f+9DSKqp/gvLb2d7pThLtZJXJTEtroGmTVsBIdB32i7jyfLohXSYGqi4UxApQss9cpRvZA1pnRU
2gBYXHeMaHN/FIpoVUsQ4MyQInVG399hf4xeLwgQWazT1BDbXIt9qRIRLlzyG/vrfILGT65IwHr+
dSaryAa1jAEp23U5RHBGFJE4vd41IYoMCRkTyBZeKetCOh40eAbzJm9dtxEl1acg9oqKIrkLrqel
qdkcSp9aKMYv1jkw9DYKi0mmJWlDXMamm27sqD1cu1tR2FHjH8GQP4TmK3AGqkev4nDiTRc2HRDq
gkoLZC5Wg5Qic2rT+E4NfxEHzbJeSlgz+nAHoAdQMRKSqIldiV1fuR4YMEBx+0WIEJwYjb0HsgUd
zYB41UhnP4BiAwn7Zb6Hyw50ug4lrVjOe0QjXhUFlRq+hEwcULttLlwkfNtM2rWrkzJSJcE1SsOg
k2kaOhvgE7oaTe++x66pE9rzfyCMbjT+Lfam6wlIWe1IQqHJvm4Tj/BUWryNUqzhjI/JLixVI/r5
NYvVwaQNbSn/9ecc7OT+E6UVEs7yLd4hHVG5nAvrD60Z2BBpTZLFb6LbtwmCBubOLOfLfaozNijo
DTggbLKf5XsUPmdH62+Qjp6rw2agepJRkte5fTg81pMomrAjkH8K9X2Sk9BZtRVmpN+lF668biaz
UdV4vfcKwJkANLMImFnxEpFB7TGb019HKKTmOsgnLGoamCXAVE2kOM/GGNAkcyOfsEH+UP4+rYyX
DMqWlwLQJ053B9JfoprNYErCRXuepmdhPVSG3omYn+8CZUZrH+VAuWb20QFP6FSVIrLNkdxG/TBi
lYJ0IkHlaDFbTEDR4bHtCySqTi1/6GdrQDQ7VRQkct+17mSpjAjUTW2kQoF8k0vsApGgbHk3a0bB
p5Q/sHZ+GShC8kjwgSX7hNLwYS/JPnawkYYgoouZqLZ1uojfCLZjhHPqmOwv6PzWCK3RJaJEK/Hu
VnZMGoXQ474r/8dUNBaYAjkEnap60Eu6NmVyJwhI80+97adRusbOVWwrzAO5y3PKf8AZIDRf6dk9
G4xnx8HcVfJxSjJFMWNItZa1LXgJR63gTaPv7o3obOGwsjlPw4UCKxeB8rbM2TXy6oa+g+lCrEK2
scZrZZobOdYjYrEG9MuVbMQa5x0hauzkOzwO09f+nfKCrFwL1+61bNihgXOBAgS1O+p0A7yKwSCf
EAov4QCIbbsOV2cruGj0zSn5bfKyol+YTN+GhsVyWbaZ3GSe3rO41owywARDI+xvPUICvV4jopVO
9R6hzihycBPB5JCd+O1ar+OFdbEf/KDQQqR40kGSTFFUwWYZ9UPg/0GmV8HHhfaXp4A6TQjWSGpa
Ho6mp6nQpmwJ+9d28z+thnylHUcwFS0hrIgzSQwKNir4oE2FCgftN+dRuAf+yg0XfEyPuw6vrui1
4KOJCiwgBn7Bn9tFDduApVr4m1WKBPxBYTNzqrbsA0bdqr6DlUe5EeeicvDLt7L+M6Oan2h1+OcW
3YqusY87+kW2dI83E2wEmW64YVfkZyhp4a/JPozvue3k/87TdmNi75matyyBEgcKsus83fWmAmdU
NFnuIR140Zl7c3/s079QO2cNm6P2LPPv7FVEnCFEkCV8kQwyUuYA1t2CRDIBZgilbAUcmmyI6W9e
+peCx5kavVqZQEd96rzLiKPbgtCZzWaErY/dRuYaG4DEIDNapNS5nEYes06MOW8e2lvnLKWXlfXn
I5u0tolstwvb4g8kWnn2IcaNSvPmXWFQjNElJhOO5XWQqln5X6fCr+BV4KpD5IfQpdeo1EWN07ec
JBaWQMIM5O0wDppflREv/ATPfKf+GCu3bQiIXUY1csNXohbed+tx3abxi0VhrEASw4eI5vCi+uzF
NZfZijwggOMRk79JP2rjAldHxdkbHjYEGL2ptp6Mu8qFhuufE7OykNkHhrYCOPZGRuKogHnmv1o6
tJllkRmT3Anl9R3BjifU85gIpPSIFpnQ8Lnc3Wgh6K6ohgGC10LIWTvymxE84LpMnIBkP5+Kv9iK
bYArPHL9s40JZHAtI0mgbjDa5kguGyDTA1Z5invYhy0SIizu4ujCvmCeoIrdcJrMqXum8/xHBFf1
ruqjBenz7buNu4wlwtIt/kaSC2U5BLWc2W/74cwAJ4Ak6TlFzPPD8KtSZ/Ljpt/qJaUf5SVrK4o8
bvzVx2Yo5BxnkZA783wi67qC6zx0YxKrJFPwSqQWRgJfJ7IFWislh6gy+u1z5Xn3VV+zhnJoCRxh
mAO9LTtelvJA3aBeiBQhHkzLRYiK3pbdsN+DhWUYt9Ni3/pGuT5o0vEO7uAuSGkshbn8eSxFfnEs
NLdTrJxrJ9GzqBQBZHnI4FhRrBFf92JOi4KSbnMajExkDEsGYfCV5bEkE7Gn86NVwQsNYWQGTwFE
gvUUEd5kfur0S7P7ZDmMh/eNTrINMiWSTqttoMme+dNw8LtgKUFQmSc3DXeURet6EqR1ReFKUdml
Bp9k3+LZiUrrmj9AFf43Ov2dg8jPpqNeCR6XU4BGFGut/GmhedJ25Z+GBZ1tvltqsrg6oiSE1upA
YtJ11/sPfPoV/vwnUInNkfAPnocw8cAd9/ecG+R4pR4mqdiVNUaQdxD2fsjsTrxt9dMBPKOM3jAV
OaEunAWaMSHwoQpVR87PScG5I8Bd5gAytPLJnymg7RMqt1rwCtCMegBKK+VnqU4DBnbbaAh+iTg3
jKOFy+BTEsUqs/UCcxRvVVYV34t+CJYQ+Lessu/Xb4qOdr7gsmze7LUr9rom4mveTLxFJL+yTcfV
ReZIwXH2Qo1RPx8g6k8XyOKOdO1ZIQLeZkpGJ45DfFKeeA8vLGxH+LxitYCzwWMp8es+ywX4kb3A
BkL1SHQ3kpKUSEuEkqI2c1SVjuLtfo/PPB5Eap7eJ6bLnO97coh7aPqGxko56+oKdD40aUssnm/5
pQE5iJLo1DO/86vdjysBpuJvY/1Wbwk6UesX4AXy7sIRdKdytFSavOeh3+pbsS6OEMBr3O8UrpH2
DWc5Lv6OOMyqROc7gdtddX6iA3exEBpGR/tXFcpF7ReHbLw6DBV3j+1XM5mZcfVzjZcXaR7i57oX
yszoKmAY0Z/KL6z0Z36QlWRjDHPrgyy3khVFVuzdDXWpjc4mkJ6IHHruqS7Dy8QaITg7K8LvQKEP
gXXzTUz8ZRVqx7P6XBEgM5xq1+AIfheQo5FdKfEbqXsBeGEvNQ4zFjkJV90yuADVzkFeQGJMmrV6
FqEnbJHqtnJkX/tPbaC8LoC+2/yOw99UkjhXmBR2QSEJwZ5rQ45Nd4LlPji92Gix1odMQWRI+Z8W
nY49VNLfwBLQhS45UBB36ikDIKebz4QTUDgtdyXUD0AQxY3t/PZ23Os39tHSup7jHI/okvQWzJhV
AL9cRFOVq7FFDqUhK1iRNYojUPr+ORzlwOwz20tbxjkA8FRszruJHvJij3XyiIZFiUpey49cY39q
e0n2uoSdEIvEwvDIRZYO7iuZD4AVfV6WKGhZh3pbr6ub/EyenX4TdbPozjijEI9Rp1pdR1ND0f7B
gq95n6ORoyZ9HJBfRW1EnspmTifqc9ABEDkdqbHXYbPZkBua77udDzonj6X071dtFJNE4EUNbSjS
zbZcRuunwe6EeadBjm05ESzRjCDxFib1FPr/E+D8AkbvtZpsO7Wbvu7E2ZxhX3rqesE+BNMl6n8g
jCpeLVS7mHQoEJjRP68sJ9KpxyyHTg5QMvck3Fi61TUv0yu8n8vC5TNTycEtmGqT6pzaNdwkAiWp
K0DFAqJGMGmwzz0J5YR2bXeoDkXke+Qh7ixk6ZUBbVui/y3DVF2ur+o7brpT/yXcRReea0oOZbZz
lfydpdIpDuhMRGQGE6AMgMdcgQ3DWiiv5lT+7kVB/PElfut2rgKuq6vGDCdl70C61IQCwb09gM9Q
t4mwEsgprBIfrbt98vbRqIkoxdtDRL9HHAtDVmby7m3jNnmGYPOL7Ssm0cXen1hjpx9oJXaHDs0r
90qg1Py+Rgviz1SA88kHxHrkL8KuTZKh3+ypr7u62H7F/ZkUSM/Y4dZGx2FiWwhAO2URu6Gm4CM7
FSuhIqqJeggdonOn5yBJLdYvUeP0JgmajT9awmZ0t5v7SLKtm8zoH8rTHhMDppIngLYh/KRO3Hhu
oeZfiOKftkUEiS2+5qee47pwAblBpyU95Hlwmp6aXm1QHep+iFl1BD81rHy2lrlemNZp9TWpdlxu
7ZuVqfPRnb3NqcchfhlG2NCOcjb8TLQGA/jM5rfsyDG8sJfUoIZIo9plPuxq7joI/pmixm0PbK/H
M2vCOo+Ho9SdicjNl+DQ32Dc96/IZRjzudGaJBstpu/KY/tLnrAwsOjwnX70XNGerIolZjWcElU/
+X2eGrGF4HH3VajSq7Dq3wWFEUtwGSGxhNM/kI8NIQuT4UEU6uqvQYQqE8sA4tDMh0Im51d1vfUb
r8zsuJQX8HgREtqbXz41XarXePg9tn4djvyZzfAat6dSgc0372dUIeVVfgq6kK58oq6oXupDZZZw
799piIuo0UomNcR3AM+a+a1KCFJnBvPf9QZqUepJmszdmBcGbcPEJZeF/6dob4qrGujHOoYoI9ou
OE1dfvNRtAcW1dZ60GFRR5PmniKvIhwZffEUR9LR+T2bBu6KLgu2APvRGyOtrdA3Ha1FlylwilxD
LEYPrE2ds0VLQsqQY9lm2enUhZKXUCEhThyqUqEb7LHbfrb04EgOsbKlS7YNfV69JWCWbPNI9Mhp
ltSRvxDEdN2044MB6rNOOZFiPfMPFQcfh6pL6stfER9GwQZBAr8t5jq+P55o9TTbjCpJbn2EcbSd
3nLDUyjPFz5B7gVxTLG89K3QYyOnwiYPZ2AW6WfmaV7U8wVgBOS2gEUUMldwIvjfROtpZEubstsg
dcR6LrGzNGr6HeX3IP2jm7wvAlT2UvvxRo13rk9CfJl7Oz8rPq7W2IgyGxLnfki3NFaV6XFECCKv
ors+EM3ycUK8pDMEgXv7S9GW18edOo5eK3Tz48TiXNdhM71kGyT4yQ7GX4FsJo/4uZjGAGxUdUcN
6BZ0l7fLJyqB77TmaQu2MngRNs4p7eJNV0eCns8v2F+NibQ0ExpwX9KLSvtUEyLqTaVhc7WwRiup
0rWAcn7yIZADEYEJdkkiZDb+0a2bcFBYxuLSMkUx6E7yWnzN/jz5cEjMBQ2DndRHDiRw7zHZCi0l
/+UDnqzwjDf5XYtpalRLiLfiAebjWWRmuFui+VFuEKA7u2PKYRGHrnlpUdAq+QgnyDGN6opaugtJ
a+xdTpCy34JvRD0oq7v5UY0mheRwhvCzSfYV5NKV6W+c87Sm6En00J1oeHBckP7G5BSE39ZhhoRb
dFZHirFH7sEI1vhlcsTsEdAb2sgYrL+Xmupw0u14vfic9ugY8VMuysh5yd9/hp150eg1YQOSP946
VOxTTFHzz32P7KLnN/5EDIPyI6UeZDEJVPJHztVikJCqJHx2DiIM72v3E3Sk+PVSH72x8/oB83zr
nFItbDBetjEhBqns45Gfhn+9Q+IMOVjUMhI9LfBzhN9rgh+u2GA0vgtrxrRgw3b7HQCG0jcR74LW
GKr1vg32hkkempDJCRM12SgURbHEKxKC15R7L5vGtiGuhL9cxcgIlWoVnA8IogGySKGH3xr3Nb+G
42ZIN/feudZR6aYY/qE9y/E06bc6qoO8Qxpl9NpMYYN62DCgIt+D15VorYMVbEEHBCGlITKcVqac
V74YZ04SugOO6i3cW8sXfuub2m+JLoc9QvIc3xN1KTYSaQY3TIQhzKZ6NNHp2vumT4y/ugffamsr
1kHQh+cSp48h2a4y+l4D3zK/iwvT2/Hy+P50KFYnheO3X2k1x6t9Qs/OsHzKuIfx2jDkq2bXeljF
49J3FW1LekERSqrjtnHr4jsnE1nE6yFelaB/WE5r/y/NhOUXOqEbly2VK41GJP5ay/bA3dy1NEzB
K6T/ddx4atbeJvQ2AOs/E40bVWCOjh9XKuRlcNCQ4lSq/Aekt+JEroeE+nqyt9RC8kTO2fzBm68H
asr+6N1wDflwINSul+da+gVwrJhRLtzrr8pJB+IwOK7VX+bfWDRqGUHw64J/p6in0EX1vs4YabK0
2kZ/LJm5kmmLXa8JGJQofbMzY41uhDwC/sE3Tz6kRTjW149IR3eA2MWYo5eGp94M4w6lyZxh2Sdt
gqcgr3IozBzS+lyoDxpYqhjJRCaGO0ALNqsxan0n7K9aOGJ8zJqn03X2qa7rxZQK5bC4C8IPTVN2
llTVxyl7/nzM9aAVgahTq/SQ7DdwEd5xML6QOK0AsMKR/2iLxicbDhUtRNKaxf3sxZClzPr/SxyA
s/6kdnDS2Pu+Rdw8F/gH83YVKa6HN05XdUXHMW7nLaI6flKW5sDCYb8S5MWTFUQJEq88LKtSmPPl
22Xjd6R+usxN324Y15FsbahdtzFAkoMouZdAcCWBPj0kqUcS+3n11qDs8spwNdIp+mCNY3zURXis
HOKhaZYJMWkPKQT6oN+PsQdtVHJkNR82xJy8dg/2mgb+AxO0MqctgWN4VCpZxCjbUiXVNdT6rijY
1FOZ2ZwT+LePm0QVCXKK+AW2YtOZL+Ls+XqVPSB8GgIFE9CYIl5MDXb1e4sVtHpIIe8NOCQ453Ol
7fCNJvyNsH1kUxpepV6lGcf8CYQmgKNJe+B3zVi6/2brc4OUH3soj93+3G321u+8QTpL5btGJ0zq
nvFByxru751Gvnp4qXVsRsBiXB9UEwM9pjBz/6b51eJRsrUs8GTjAHCHDb6Q+NWynfq/Tz8R50mu
vMVhiga2MoIPy/B5IWfKyRHdq9ANC/Imp+22YV1+w3Mldwzc7GzB1nes4Tj3cjhUtiCASIivC9+W
AfywvBgm493MxtzDXBCbhwAHiMvDgWeu+BvhdJRClMcHmoLe/321J9AFG6Yxd8/Pudyce5PlHYGH
+H9PcL2EplcOeNkgKDs9fHU11goUCBiQhXWEhTqQru+qM80xzFuXiHlLyppMgFf/ftGWkFWYd6jk
D/sXhmzRsz+BQHNl1X9loMf4jgD9vkZkHPxPPsZ8niMSlrlsIjxIXSpZ7eQkO0Be74dClu4voESh
3CmNMzajJR2stpNwzzOvuYWrXMxIaxVvRL6JLE7AEjTend4Yf3awGCRC7r+zoFNKJJ98aSZCZvxp
LrXKy4p0vjf8shRZzeEYXyhNhhTMfnHeApwM9TTxmCLIPFqjwK+7eYNvpzExfVH1rX4ZBMN0jVMQ
bbmDACBZcxKvJSLZ5YW1A+lnG5wprX1i5b2WGRAsxAsFBChiuJ002f5VraD21AFT5KUqUfYZLILv
QCIoIQ2jVMJ/EvCmorB3Jo0kZ7I1py9lGBHQfyoJVdjDhiSF6WZy7KosiMBmrIBKJBxUFwf5XdGM
SD/22fwZBoOdrZvI5EqBlzJQXRaygvh9qOaCv93QmGY0wyk8Zzh2lcp20F8AOv+uSxRFlsTOICRX
VQA7lLnUsFgHKB7eQpiwD9adTojV3+871PTQqNdR1Md5ln+pgpSDaINircJAaBy9uIAcE4UsCr9h
pCpbFhQYuoo//lVymMuk72I8fH36oE3d3Qj5n/BPb+WUoTulT5Tie0Zom9DrfpS4WqY2F/cZJOvN
oE9mtDAeiu44XPV/VKf5VNmSTWpK2FWW06uOiYyZKnmVaAZXlzgiAS/9gFy0wJbarluf64aZqPQl
2io3Y0w1u0B/8v/HXWatEZVoVsAn3ZRmRY2tbsvFiyqdLzy7obw0CMpZMFpBFB8/bYmk/ZiRs+ts
ULQz+xYU3shoycOfD6vstye0RpPb8SFO5z5ja/TUp6sJixzbQWD3+bApawt/NH3YoLaTwCaMEzqN
+LH+mHKh7qX0raQNpObL3GXIKQzeUgfQYARRmKN/ZrMXH6DsN+O2GsmSx6yaZgwbnuMpFEK/tzUN
zTQCT5kA0LhMgij+HHuF2vgUjpLIkeDqFrrqxadRbOII7F0A+gmCRsoRht01OP4C711Y0MVpFBdJ
5WAampF9DJeSYscLnubM6Thh6uQr2id9ipVmFINxqSTGJMD7wVQbY1daUyFk4yPjVFEQ3yiVE5Tl
2n6gH2VLn1xQWCQmflo1kX8NkXGaNwXxaRtMLPjiDBHmLQal4KdYVDiAB/GPEpbZKN9dTdj3xg2z
v685rVGVtv28RR/jz/0DXmSlgdGd26xF359VECjKpZ31g1FVTHdMNmfyLMMLV2Wvof25IOUssHip
GjEn36negjGjMfgPyZw7LVtSn3+lJt+XXnEw5BuLIOg9oxEHLn5LzJ/Udwd9Ojzu2mCOgyUNgRsb
yshqa2NZJJHLfqnxo3tdxF29ytoVR6UhnpTYPY8xTGrdDb03Urt1uo5URrICvwWCvddlVieI15Wl
KHhuQO/fPuPXDNB+O9Yhf5pKyuz2RGQWYuySRx2LeW8MHkJf2XgXMJk3X8QkFGCHEtR5XMNfuHyd
DSRsp1VqL4P8OSbET/RL+RUmurqeQDN31W+NIcDn/CqxbxOmBSPIlQL/VQL9xIEm6X/HHOBIH9BI
3wYO0iHrozdOWSciUHrLnWoKjykVSaW+3oG/HnAXJAfi01PXEnPFejbeCYFFNCe3n70Ga9DkXN83
AJF0SCbNQ6gKg5u3rIyH6aWn6AjyiLVXIcqS+lK65c1hHGF4Yn47Zcj0+iHNddJ7EDAXRPJiHZpL
cBMsDqtd05x3IM8d18Oqz2qKJrngq6Ldl5MlSim2i8pBDlqfN+ntPm8GgGduF05c6Gbtv1U1gncM
XavHrKdNQqxDgMjhwtxZvc6235mucsqgSOmGV2YrZD6rPGcPeVL4k+spJZb9IgaG/yWdgz3niVUt
I9y1QsxaySUWm7IyvEy2S0D/7uEWjOE94zB79d13zRXWg2rJ5TT3EX8Pf9vaPcW8TaHpmuWnN+0S
y7PMdmWTe4rtLTzH9WmLjLySEeFUNh139zIQVYeiuSeGLm4+JEKPH67XIYCVcCAAqLoTNKXw2Y4L
x2snLpVOClIl25dWpIdg1CZ/JeCOkUJQ3Cj+ukAJdDGzHoACNEKKQ5Jk2Mo8js060Dp8zAFxPYfv
A2eyiTfWte+x4wPrS5bqwr8c4GN54GymK5qSNehYu4JJVASv/knESG2kH1tRQAAyUJ3lmXg/Nj9g
3qxU07FS16PGtVt7xPe8dQnNupIrFRs/axcLqbZY6/5K9uevUaoyvqrI4PsBhLB1d7mvNb71B+ei
eI8wm85MdVQHkdTcWWlJksubwE3zUrtvH5wzK2AaHV+1S8AAMRxPNhCXTScNIfTFCodZOoHjWTYm
NPsiGkG3yzHMM4rNzTnHdB7QFf8iDXapB4n54pPWIs5gWSyT8zeRdkEI3K9XKd0Wdl0YbnYHfQIo
CU453N8iZA+1+utcO53T3emYO52aY+LJR6xizPh13V2TI2I5pfVOYH449B8WHM8NGF9/XXYOltwh
S97IVZY/2RYmfHEYLpH3eB+BsMKsBLIjyNcq8dZQrdpdjWA8Jvg6UOfFqL2Cbd+pwF18jDrtQfz1
pkgM922JhRhvG0occXjht49VAYf3zajFKpExFkwPOJEIDIRilYiIC/aeFfLVTFY5njNWdUjkX9p0
C33CJUkNLQG8HL5OdQ8JRiSAefap9FC/MDZn4k0MB/xGTk45GRoeRpyrDsgNLvpOln2iCfGMp1s7
QS9JPzke69mlwWQrH8S90Py5biVxCjqK6jsrmsQv6F/EqvnfR5qLOT2dSQ77YDUFFYVTEhPUYPJF
i/hHWPtbmihbH//Tq+3OmWS+GlyXqOOj1pX1bGfPrd/KyblwfjS7QL2wykNPBwjcYoClsm+HVEHh
iotopI2xhajAXtr5IS6ZkGdry6N+obw6yEukTVpKyfWLX3rrKoDCrXmZl9ZUnZOzywLpCa0li0tg
AlWBNYxp7qsxd7pTmML7mf9sgg6aLBgDQ2qInB2QVKowa+No0CWRvw31BhOAlR7VC9+NfMWPV6T1
LnsuOX7mimP97ZCTQArYziotohJx4dArIfSSEdhieM+BUYMV4yJUnruZYIB8G3TasweZcdoDuNm1
k9rGLCUkFd2WEqvhrRbYoxbIj63v7ZwKG3xL/5/fwE3KtEIgE8nuDQ/ormueuyS6B5kByZGmesJB
44RWq+ylRUWgiC6R8tv/B+0vI/gRvRNVBSOT063iQW0XpkDY4DW25ZXjt3NyRVEn2h+ScgUa13V5
9rpxLXfvpl1I9QbwxPAvDRNL443AQSr0za+BLEKl371SITbFr7Uv/VMBCjuLq4W8icxJ8RJj1MDa
VneLAfvu5+WilykFZLyVwHgq3WnSledbEKAo2n8AxIMNI3SC2Ln+vYsWmkWK9X7iVJ6jX73XjS+d
vlc62X1/QEjEO1UnjWYgiuVqshyaiclYweSxftt8fgGiyyE+BZONF1a+BYnELaMRCiKaN9s4uRND
7lE7hgsX1f9BekSPP382UR6ykP/i5lcYTAyDG0RgnNSWfrehhaNmG/4zuTHkOJGXbMD8l04Pj5V0
mxKmxbcB4qLEKV+9MuOkSGTQ15jX3XVTn+pHD914YN4vkFecXO1T2XT6K4cdQhN8ftjiy1uVBvnX
jI+eD5igX40E4yx4l+h7WfchbkeMG7ClYUDyYZTmFpNqCHlz6OszzvWUJircWcA5FwbO8K/oVfJw
WFU1iZsN8cp5aO3Sk6udjYcbEpvy2w77Q0BLO1AM+gvAgLNWE1zim0IFJ5H2oeISAenzH1DMENRH
RTuKKtJCh8xMcY4ymYxMSHzEqn+PQ4kNWrn42SWQAnTlU7tF+dGVXk65H27iRs74xTDyzB5pvFE8
uESAtbdTfxykMk2ywwCF0m4pyALyatj/iWvoZHJV5PsPvNUCIOUTdNW9ermkaZHMyOeI/CopRAh9
U+76rtP+FMOV1fEP0JrNwjRamFZR4xJYmDYylKwDCyC5DCqfjIgahqLBiCAJrwybax5BCITGhpKK
3elCUFKH5HL2XgIIggp1i7x0t9WipOGoVHeGpH7TtZs/Wfi/JUuy4rZs/LXH/TNkmC3oAzCD+84J
J36pZK3qEnE7fKSFIkLfFINNLxJLwiQ5iR6Jhz1BabX6pgWDnTQlVE41ZRcM/Y+fKVU9ToeHh0mT
d3Zos1FQaDwPcixBoe5CvkuC3TZWCOFMJd/D4GMa4D/lKpzYGX/GkpLN+MDfaxaSeX1NUQdmwPTY
GomgCEHAKoMGf3qcYH60Q73qvg36HZdR0yLEbavyA5bI93B1PuNkz3GVYzCpvSTRNuKV8bRkMInz
OXl965IxzunFmcEXtll7g7t8TYdfz1EqfiIkAcDAJTWZySqWHogKX7NSNZheigpkvK+ftIMcMi/K
d+mUM3m1QQEOQXzXWwgY13NGzkFkkuzPBXslQ2TvcysGUfqyR49KFVeniUfkaXZMU9o/p3f9XDlN
JovIDSJ/aITwOnKEpqhiGKUdg/GT183YLs/hj0U/Lih88GocvwnVwX6zPaM5Io0SJFS8FxULTYjs
gWU78/Xt56rtaafrNgAQuodQgWF37DrfD+UojKXz0FNJAC6jHsdUL4lsH2Es3C1okFkIkTUj8Abe
PfaiuWf7AyyrNSGhiyah9TuWj6j2yIVLsr2korTN9rBjWjmDk3BSfTSj7UecRFjOJmcqVE5d47U/
iLofjbWNyIb1zFsAy1rqwH4RRarzmo3XCvbUjgVEBzVKImd5iJPjZcYUnrFpTpmSr6oA6d5EKkIS
E9KqH/Kbaw6uBP0Rb6nEKGTDxTpyHjsVN8shQL8XT9wiJMpHeP/GD6CNkjEjwn8m9mLIEnomSJo6
wNDSNP4fnOHYHBoyz+wxys5jnEFVMcPq420+ofih0KelXBzJV3fCblB4Bj4zOCwJv6YGzEgvS/mk
nxjho6uQda29g6Kwhz0qHfQk5nr6dRB0ygamWQZtsNFzR/eq0sLuWDm2T75rag9caUQY8rxieNqe
BoXEXPXriXYyVaTH/W13FefuD1nN+6f035gDd6YxOFjFfP6WUUtnKD+V4Etx699XqCeQh83lLO64
uv5k+uRIsqWDqyPlwB9OLum9IOo4QOVU1HUNC0WtcnNRSQziJYvPT3uicCJYqYwdwZxBZKvv6DNW
dCERNXIIZPQxao/U6WhTkEcwiFVn222tfMqUN555BrGU1hNZySscIEPiYJE3FP0rXNv3Mhr4Nzkx
etFt1nanA/Lz5+eI25LA92G97WBkzVHK30STrq5InMfz1vc0ecWaZRn1onVVcGtW6mtYoamhAiNs
KqV/UIbXYSgEhWPoiNsbL5NOo9ovmGVDGZJWcy4C84gaE6oT9n1qOw8idRLI6hVmobw775x2eZ6G
xtFEYYu+vF1gDWcWFBI3ulqbGogRSRoEuTAcklne82ofYl/NtRTUYV10vh4alHT29RhKTJIh0LBa
2K15LXyOL55ZqVAqa9tOh/cIB12/aUr7dWw7stLqzlAJQd5y5Spcuh+cODbXzsbaPM4P1ei/gc/X
qupewP3tpIhP5xktJybveu4G6hMxyR7URQcH1kHv3+XAA3YhnKcpxVvsRi8oJJQOc7l2a4EJrhyr
UIOa6zjtC1m/RdbxIxj94CvdLA/hqfJoNHsfS+pVvQtcCw8nwXQEWtHiEZs76DuYcKjTgRB6MVd+
OXKcERnGpHoDGzhXuMF/3S8s67lMeiXFO5lU/G4MmQKGyaQ9FvlTKXu8GIheobB5wXC71ZpOuYX8
HFpJGmx3zZQwhv3/4D9fjJzhS6zDtgi3jXTDo+Gy5vkh/pQqpqooa/jlD+FAPLgdsv8x5OatrLUk
kDr/kRNlDo7coMO8Hqa6iLSRt4eQos85ju3rEi9PwaPmRGSndnn5MUPZA3Qw2KjdUGfiOqdCPoWf
kD1CasYNSTjtT5uFqF4+4UwsncXZZ5TiReMdtYQFMONwtT1cLFnGjG6CzaKolkJL90EjMrN2kari
PrpfrOi/kzzdltsiAoO1kpXNMKXc3FxXQ8CO57+2J/6g7cFkQOmYuPyyCQ3DD4vRLSAaEzzzw1oM
AbOt+8gkyzpziE69z8ylKbj9lxxK7+gjUnIhOjbhUQEhtDcE0QYGSrBJ57iKMOBVbhfaD6pVzqT/
AsAN9XhbXnKcv1AXHqZPnhZlv/y40vlqozf71Oy+R0A2t0w1Siig8MH/Yv4Ank1Qpwyr9YmGc+Lu
gj7w43zuEJ3HgV7sp2e18o2qRfofB+6XmyuR3WnpzkzJCbiq9Yy90GL46XXc7JGkitIDlbk1rX03
e+zp8oX/jGhpZdqg4dxPMvt0BRL5G+SfkbkLlSNjiEmxwbOypl4lgSJ9YqI5a2CsD3xqt9iH/Rrw
nwm6OySrzj5yvv3tjsOwJujqA2pC4Ravf3g48FHpgaW3MOodml75NdnMxwsWxQJebpWNNzdC6HE4
nYDp6BuN/AvwqzUaPkX+cGu2/rI6hvT1tPc7o3ufcrNK1D3Ibclq4Z+dwTCKXxYQXz3kfATttkAL
B1Uq2t8R8qjaERh7+G5T2iMpdDndPCH4jnVgeXRzouj1ZFXsozGvRNCpHrNvLRCEqZ7GAhNj2SKr
K9RWyU2Kj3TkkgtL4KV6Ny9ufXgJeenRz2X1G1I9bb0jOPTn8ygeMsbtvalIs3mAN1dyxlXBJHBJ
7NYigxTCQj4jWhhU6IJvkGMhLsbWfQ+31kDI2zM2Qx8JnJDouhgMc2TpUpyFBe8uOkJS3jT6hL9e
ym59wjG+HJNvwQaW3CPtyYRO/j5jxG2OjDSnPczwNWuklpoFKJn+q87JqsC/94fXBUnZkW8jZQFy
54h2vI9WcsHcC5j543w2gDEWldLLu6LbY6WXY9m3zHpglWigj0N9LWZC6oVNjSX1OHAeuuq8HkbR
RVuFXkmuC2yTNjXPMBHO0LnZIXqtS4BCKw5vhy9+e9Qx9upyzCZYaafu8LcKHG/EIbP+XK6ZUTrr
gaY7cYFdYgEzyL7DUya0uqD+abWHO/V3RMlxVMXBJek/oxQohuvIo4K5zRwETGsZk1KnrFI4lsgz
lbiqb96UIpoa0ks/OleFTuM9GP8cUKjj0xTe8KMpK5XMgI5Mi9achYdpCIYYxHc0jhpe/48dcfr0
vAwYLgTJLbc+JLflSL4xCzYr2yTHRuHmYkodoB+0SpdYHhskB72SXZGcuMBJEYsrLqI0kenLVENN
wCBn48QJMNfoKqjzOmMgkt/oIDc5qYvV5m904kBWuJzheIbS6OtAaazBIFMp+5YtmXfCjgSpYphD
qH0I6h5ya6DmtPVvYmCrfYWqIL+5GrCWe9wYuOkUXOmpzeiQV7LVyp3NHzUkx/hJdzpls8JZrbPE
29/dujk7uZ8n8iyEBxP+hKPBR/dcQQ9h2I/bBGJ5ggEVCpkec/ZgUMAQBFUQ6v7nf9nd7/BzR53Z
UpqLAV033ciVn6CpsHE1M0wYq3hV2Z/iFgqZsRZvXVdMYD17VhKzDKIENW4Qj5j8aEH1uoFdQTaw
YcvkFtQuQbbX/V427ZMrdQo3Jr4wsCktkF3D4qDF3zqS90PmPd4T2UKHp56/TUutnJajHl4UFhHt
2qbiOna+0Y1lM/l9Ei5beEgVuiusaVEcFSksrAM4L9b5KTcDXuNU8imE2rsc0D5rFS3UZXYQTt//
DZBF4KMLFo4xQQJXTU6xAzFzWtivHcr5c8gJQaBt8zKDJDPzOv6gbPMUMGHVkiSxvbmEl2CliGWw
gWHZNCrGV67cG2fCEvm9GM74iP3C+d3LLQff76ukdyxeJVnr+BBwYE58Jyb0CgrdNqhLtrDXtiiX
67XZv4FsOGP9bIZTgBnhxmJf9h5GCLQ5Oy1Evir1i5NLil3eCNZGq4XH0cJLpMI4REbDyhq2c/1N
pEL4Co4wi9KAb11jDdGxVbH96DYWSTUaV9YVvtPJ99MgwEj0iz+xhLowccdQCeuCgYODcu5xnrkc
LtsF8V/uV7kXKoXqlsCdv++80iemV8cyycZTV+rLpt9UnmtjesJpTz2VjOzVD48ijBx3Tw+V3wDv
TVNV4Xy78f0YH5B5gk6/F7AO0hhlHfoq8pXKMlXUBxEhUCGhxX1AFF/Wy1H2Kqknh+Q1uOTho5RA
Md6kzDkFmlZ917wdxvoqfN5h8s9jR+2RhZOYdgICJ0UYwbhHhkOKqHO+l042lJCFxpT3tSF27izP
QbsaIwhYhI5MZLhOJtq22RTg7sF1bnOlM7wPtoS0z7gxoJfqILZsEVP+8pMV1wKRgBKpwF80rwAR
5Nif6rZGdonC6rse89CpAvrYe0n6hClgIounC9hL081JaX31/mhSINr6snaIUTwPs0tB5O8j0sdK
JgpIh45nr4voqS1vjGpwF8VtwCcoAVQ0EmlWu0QxNJCg0db+h27XW9Dfiu5GNAhFoKmyDxkw8Fcz
LMgW6uQ+YsTsXwcK0AWea/4lhq1AP0OCkBR0w2GzttEvRao6WjYSA1JUma6cTLP3st4HMZnWAS+k
Xy8zJEvO1tywlSnTWzlsuR4EnItw4dxj1phrrkzWsXCPhBdNx5Nz3l99KN6osasj6uDs/Zn4yPd7
fOAKlO9dok+ICqVXmf4UFrkbSLCuiEWNGD8+AN+3BotqTNhdDoW38tZb8Is7ERv6y/TWBYE4qx7n
AmQKpkhM01fRQUgImC9wv+LLpATmBIsiQcBrXzXYl3DgYpbGxby3m9oh5vTpdiaRCgwNCIppj47r
TwZ9VPFmQvOE+MGdzZ6yx1W3NskC8BD8YWhLxtY/bnCh5TjW6LtR6HL09qIKSctYGZWfNtc8bGXc
3AMmXGKsXqaNIDeOQqdEWeZcRtacJeG/8+OL37zNlywtZ/tY4tseUBwcrTUve4iLPKRdNHTkcMF2
ypi4oLB++OHUsH88RU4pvSu7Xpuf7TThe1RJY1piuVhGTHGm4vs47dEm81DEMoScFsy4rEE5bdjJ
1o+I1pUjYVCgRMIAjiX6sov5T2/rFR7iKDsmf9lReGEfdvbMGEOStHNdwui+OhswjSfbs8RruD43
FGb8iJLV8mD2Q796HPCM8SepioZZsP5MzBtmmlSJ0HGa2VZQDQIU3Sd9XQyUJ5iw4fjCEmI9LQeR
YsKTsD1luv5IFtN5PFhvUCCf2Nav7UNmiUZptaiHjUvqQ/seP7DC7zwAMGs/KInOmRj0q7UUx6ZN
Oz+CAI3pQrHFg6KjnMhX9XvSkKiiU4OTTH9qKYLryv6r5AAnmP8Wy8FpeXsBFnB/FoYpdwxLvjlD
1ZbbfwhzmKdBi0DO/qYcAJBl3hmfKgEV1UxucbToRZHOO6XRvoQnQ13WFp8ujeYTP5je1lshJqVX
9luHTDZaJZQ8LpSoJELRYLJwe+w3tuvYSgsmKmYJUlBzu9SLFK66S0h+Hgg9XLXirJZ/g5yHapqz
kmUDfUoSUhOQg91HjW+glZoTkXhy7jCuqxW64hPBQ79Heo+ygr4eLu2WY5F+STO57+5YkdzuSCeb
CZFvtwd9K1c0WPcYmC50BSQkxupdwZOAWu2r4OQvlkOTHEmp32f068cg5Txkm5wiHG2w8VpmOP7D
uGeDNzmXppbuUdzqh+H2I+BdxkWrFLhhYDeHtZbA7pZDw+j4hv3YDidzf0neRnmKn6k4V4i1ZLCh
w/8NnySJn6EFratamvbKwvzRv39m+CUarfX8ADxj1+Z31PFXJJF/XTs/4/RCYGRh/IqAg+mXVjIC
KE04/Vjgx4Qm6iCD4y2LyvaRy/Vm3hIxzGTKGgkkq4ymygZFFbtwr7OmMlgqsd/jJfUd6dbQgn7v
LUBy7LnMTzaJ/CBpY/Ec+RlaizfN/nbn0J2JGPjbjzNdcPL5V+esyjM0+w7PF6MxhClJA7a3ZHq9
mH6PkbkhGemffxMjdo6JH0S6BYrR03OlC0QEVc6AtykDI9UG11k2ztS+L/9Q7n2pzUbbIpc8mvr0
fehv2xc9MDeZl1BWjeVU6n43vjbeljSEyZPeW9CTNScKgxEPVM00j6opXUTIUDnJ9o3vPurKpOuE
Wpa4o8jxYjgK9w7eUxZYzX5rxreqf55Z12Qdlk0/NTMPQJfBVEA2kK/sQfyvnHegXMOANEUr0AeT
j5IPBV63olf1IeIwovPewKi5r5L29EokeE8lb0vKyJK77WqXR4sEwe46nLDxaLrP2ukL4JAZbuqQ
BWJu0D6CEoSFoMPVK07U5IE774dPEVDNIM3hte7lyhNA5jtEWMm6rfkcI042ln6GfcTxV6Oqp11G
C6LU+hk8nV8tMAMq5yAYl/8Vum8+b+Q8sqPQ2BdqX69N2wcawrjhKLy08aB7ySVBe2cdy3wxWxrX
34cZdU5wQ5xPDQyU2LqXfN1gzTp0ttuI57PkVCKGID/CXKfcvXjLhzl6YdnwtgZgmWoGZ+XA5EVL
PFQ5Ugn7Hf9/ov8WQ4eCf9pq3jSdb8u9y+5ci+TVaz49zOiU1IiLyHYdHa86tx+DnKoq6l9gKEnE
BtjY1Pm/KnZj7MnuMIkbHarLHIJBFtlh6F/j+frQZuHeZ+b6GPIdXZbFPqH2wod6hrCQM+bGDnUW
aY9PECpPaqBkbtY+7ydCRutde7ccQ1vqxMxk6PqioouLw117z2mwRb6swqB+l7sPe6hbTXWgfGS1
F1nW3oS+k9h2rzR15yOaD874nbUjsuDNTvws2lBOyq2bDvh9otJDrpzk04cEXZZTkDqXOHsChg5y
UAm73v2q29uD5+H0hc8rwq9B5K8Y7BzGG3fsboVxBz5LzQW6OiYmEj9+UT8epX7sM55diSRS5gUZ
ULY7eoBC2V1Nk1kD91C2aj9PpPDsKw4r9X/m5hqQ4DhYVSYeVdYJbo/8HvmcmEJWcK5EYv6F6FAt
yK3U0w4wft/UEDJzLcKXzEMFCcxCHdgnY8KENQ1IRxpdtiNuDSg23XJ5XKbYZPL3bW9Pbs/04y9S
DSfQQAfuQhuYnBFeBLIak61/tLsI5gseVAU/vD2FL/HhqCHGwXhAj7NSyNFq85N9Edj47urJi9+w
xR3B+8UlzPNkrzdf1DVDXEtrz1Ma6xml2SsMip1JUQpTo619beqMuCdb+SFQ5Ed3zF3NqrCV6bpu
aGO8aH5ElKWaKcT20SdGCgjpy1M/9aaRUmdCZ3lOTpQQzmgvUjKIFkcIxX32T7zj1f/OIj1c2/eT
4jH99mcIlmCK3cze0Q7UlSNIUzDeX4/TMehQBjN/509xD5WireKspmOhRpdw4Nc6UIsGW1JHoUAL
XhHx1rWu2Jc42JAgj65la6sTRHfhey8o8+/DSVnkB+EctsSgCshLiA0rcTxQqSBJD+dS7SA/nReR
kAeNBp/DcMLgqosrgGS7vGiNkK2SkYVWIUgoVlLYflEX702DqLgyNejSMrKmZiVsG+SVhtbGIIdz
yMtktT4HYBc1mM4aYij1LuwsdLuATNEd+8xzqVI/fh6nU9h26bb0x7oLtTsy1eCKUDrGzpp9D10O
3oucmZiPu9P8i7jN32WSm/RcwEbYorfNx5iqZvRKQQO2MBfKPs4mDVHFgF7iGcGyOn4CiFIqBTo6
EN6PoT5tNDftm0tVQkXGfZ6O8bLyNDKn/INjDA1E25uXYf3oNxb+whBk1L9mjzWUYaqFyKvLjMgE
6IlcChuAd7hk3atFBnhAYoFq8Z2GQKy0vjwG9qXf4CKdiGfWjHV5GAv5I7BLfiAqcafQlibgWzr7
CKA6Iwmw8rKMiFfathmAxREXCL8Vkl6/kt8EMNw88dbKs2aWzneht7Mzdy7nBEYjmiqVdOtbns+W
G2IlhuBtIzpAKxLAOxpoCmp4q/fH/dzxgKy8p4g0WyEAPh4hkuS900M7ba8XYlzKI0O54YstV22o
ofILJMTnfPM68N6c1JwH/hY5bWzErllcgtQkMrA9LBj65mKTCbv1PkAeAR9T6RX5hRPCvJxqS4he
b9ofQtCnFOFBzVGAf6eQ/gtDNuwAfz82YECuyQBi3+IPg+CKLSxaWLNNxHpLWh3jn0VKwnv6UDMQ
fb7mW393JJCSe5qN4oDLu/Rx0MmP7z7AT00gzdmKxqKcsz48OJxEPAK57gTwOZU9rMYQklSSR3wS
nGOgFHy2mbT14lOO5XvZtPwKP21RPC7srdzhiJV5XfeeoPA7bp3myWmFggqH71U2PcyrxfxFaxbl
MT2dj+Y7XMVcsGw2dP5YRvrK1cnl2jKunzeMROdtg7iFOogUUNBSn+58lxdt+qVnsWUnvB7ef1Xu
E5iCzg7epgBqs9csQQmbjWhbzozetVpO2ZL3+CEIXc8jhbzNvOfIKMzbCArtLXh68vnj76RGKWON
U7S2LzIaGCNAD2ZAKP7lgOEtZeyv3ODXb3Vv+X+MAl40SEDoJgNn+EFsgY/qGAbddmUzJQn3DY3a
6Se+z68MpoXIyjABCQM+40orv9j6nvaOM+gOFO15LZ2VFdTLTHhG5dYTA7CV/7rK9o8y6d/AZ685
TIyOt2O3t3gJdvopGuZKG83SAfh35uxPvWiUXD0v17D7JhCF39yZZEObnSt345hrqlzuTdtYSiQo
HBo73XNPPfM4yjgr9f+lJ+JyD7muDzU0mDyqt1qRrnGft65n7Qc4uUu4uPAwWNVNat7vM7iZfJFn
RNIj0m55ooFbwrAcl3pgo1V6bCW/IoOUWle3orE/qE8pz1Tj0ACPssZrANsck2ZmT051pWGlUGhP
mZpl91hJC7pEjFVj1j01zcPUXw+d4Jxpvritc6cm5nPRKpeMmOYL8I5G8fWepiBRe+KJz29PnM2W
X4yQeo6kVAn2cCXuzyZHpMFKQoaNXH8CiWZMRwMC+phZPBR2HFzI3ZF/f5v58U4OkOt2vLWERvjK
5CzdH5LwMZLZUwJbGfyBcNZ94xG1U2u19EF9QPy3ZT9SYSYcxRSS0iESkN0PLheipfrSzScb1fx/
mQ2hdD8zgQi/zKHzvAJjeFfFK83AiQqmDJ9E8x+Ti3EKaAMXU9bjO38t/3KsPHBTNIOeoGJku3EM
GAEjFnnSKxT3+g40VfVkPBBQ+gG2qY1+Mn7La2zBwIfKx14zu7shDHdrZ/0QB3cb3O8c6DiCQCq8
1tTFqSNudrOa40mFbZkpoJPRGVorb+dGqa6XfCAetB1t+HqtSedOhuR1TSDdf/889/u3EtyMdmX4
q+Z+SoTZiHxTgCeilzVfrJnsl0QIvfXerMtbM6H9G82szhoOfbGOK9UOoSe/Q1+3dMHLWflfqdly
SXP9BO4i/SXgHQOBZsXrGVNkmVHEr5mlW8RNS7rXlm1yu0sDOM33Dh1eoqagB/aylEcs8htJNhQ8
N9pPsTpzZhmxCxGn2phfLCxWaeIsLeplaLcJaCwReIRYmmDQaFhu8kQwSEMNAGAyBXTpC7e4fXnE
LnckLLDHq3rwyVH/b0nP5IO96Jm7G10h8eddQmuGTLg5WItSBSYoMoBrPEa+Ctup313QQt2eQMNG
1iU8+mOkvBtOlYQVioDw0D59mmsEgMqvZNe3+lQpnEsSoFq72Kq1fb1Oa382rM+9sghUVOE+N8c0
BUFuN4nr8LzIHtaVNqy41RB9uxwprlA5RYyC9g2unojPzBw4D7CWRmte7gaXDWL+GK6/2zfF6Sz+
qJhhkEYfCEBBS5ghS2B26bKgGMMwTT+dgw/Dho0W3Mz4rdMOiwolH/dKG5W4GHKdxgpRbNq6npQ2
it4p7rd0K0WEiqHgGbP9UwR7pW41IezYFCCiQwoISCC0JexAGGvWVZvJri31GJORRJTY9Qkgka3l
8/KBIgTvsfXbiLnSgqgmHrl7OtaJwBaX6px2Yj3Lj4mu0I+h1KJDFvwYag2ULDqKQAB3O7UOYQLJ
OYi1UqdILGupEPYzTZ9rUYmKwxgCbasNKK9/n0P/0PoJJfe0JnO3Ffchvn8TWg5E1FJy7MXdpF13
bokPF2HhuivsBu+1lLl/6rlBr288UmIa0zAqrv/tr6d10DWC5N5sbWh1dczerBZLTyBPEC+/yWU+
TOwWCzz1EIWJZkAb61Fk11jd++EQ7vTZE9S4CMXNJyeRe60uUZlV3504DPA7+Ef412MHseFknNcB
4TdaWcGs7ynrY6ZZE93aKvYYNmfrzBatVSLAdbmgD/Zw+3O5WIEowoE3ytDs4KXzcOFhuxiS4nNg
eWUNOo9JI+pZeZB/Xz0tX1WNJgJhT+0qlsb83kVn7jwNoVOaVUjpirP2NMgyURwQZUO6dbo9580B
X33WGbfoCNZNXYXyMLoapyK7jibEUEijQOFfxIp6epNgaXS/BaFEhKyOPO89tM3k78XV3tqDYmRz
kxFjeGXGLrFyDEParuLnvNW1iGy/PzyT1Dot3cKJRYSbjaQSxXWNBKYU7tUyknaw1c6CnGtHCAu7
D3QlDcxuqpTzOWObV6E7FVhACrvs0xlefaZF7Lgc/C0ZqEr25vfG8dlb+JOaP8m8fbu3nnIw1Nkd
tab6096w5xDxsRVS1NzbWitluhRQZc6UXbVyLzndfXcmLu0l4kmdUMMgZ6n2PKt6miRrecV1mozZ
gU96lxQIELpGSgZ7xY/Hisq3s3WwVYI3bxIHtVXu9b8adxajYzbXewN6rnqEdqJYjFM3fZPydTtK
VC+8hvIGCVC9w943zSeNlwFr3uzf8m7LaYRS2jMEnQECaqO+5Xqqj9yLa1S3WxZemBjvcM6SMTr6
Z2OKGR3WotTcZXQzbiJaFm2PUq54u+cZJiDuhVsy/QX5bUI0qNUTEFU/ESppJCUjsZYADuxEC384
3Af5zC19X6nXaUruo5dtrWuLkycRCnmfzjgZMyZ8JN4UxeMpxvOwHCa4y7ky1XVYcxJCkCYqFcFz
NDEBHkWZVdEoj5PSI4Z3YsuXJGKvGg+C6VPEw5kfI/eYkZpNUZliYm7sC904LiozPwRBT94F0Fd6
xcanl49vTHIqQut2Ieb7PxTEor8d1gBrOzGd4qpubR+sF9Glbqe7pMynnQZToClsHCiyP4swqOBi
Dkv1T9oUgjicmk7GCArwzJF+zrFSti2R7UVECLLus7GOLNnb1y/1e5njgaKAmLDiLejZhXfHjNPT
mv5FSq+bNXh28KyZJKOF4HyBJbnVI45iuNK2y/qlkg299M50tNrX33knizZ/8Ko2jG71RdB9w373
/1I5TtXNb4Hz7Q0VuoVM3SEjC39ZHQKR8pT8NJDfv2GSL3i9u43e2vBZTBSstxBosVhOspByUqV5
D/nLQ332NkE7kdPZcJp83Mu+xZ3wVrOXGTeXfelYtEmUrC4nCvd8WeisJ3Dt/A/AIhv0sVAsUFQt
uFo+Z8FASEck7ayLlXpGZX8WkmUyVbpQpEkSao2tIukV4v5jozlmikY6apFiHfFHzcFggasaV7ni
+sspP94wP0g52D2MPxfAIUC8WhliZrYSi0E5xvhTdvTwoNIJfYzxGQC4waZxj6Mh/cJBAT/ViqD5
SGrI3PMrSanAlMmIBTs1mxUinqr9whFDRPPOUIOF03H+QWWJMEgaBTzJur5R8HmQ9NHY/2YqIqrO
EsOCQMWfglbAv48aJ8t+N7puXb2Lmk/4S7CLt5E9hp681TBqbD7XjJ96GOQgigjb5ef4W5qZKJ3J
EVM4edGUYai30O336MrsGYSiprP3H+M1GpWWf88ytHFPPth4M/aUrwPFO1ZwoDt1xM5/ucQ/StlG
5RcKmsSm+LqAOQU50DKkt5TyX/AZArBpNTaVfsgX92PLUBuVGAZ4egs/yYLuBnlPOWMbNXi2iukk
ov9zD3/fkO0i0avFhX3pLANOihrz90idy+pZHRRK+/eS3Xn+Jrm4DpM+pl9gvSk4/gcLv9jNC/Tt
JoilCoFdCrPh4PjumblW04Kb/OyhGFofMXD/sOsqST6UQk86srtqsakqbR51UIOaLuAFavrj+tVw
8LxJQwHzuHNibCXXruAELFl82D5jRsRai77vRsgiFpRQLhe7sEnlpkZdClb1bGpppi9tZzaEk0Ge
UqVXpiHxswEoXnQZTe5HR24ds2Q1VGYsVmZyZjNW8GzNA+Vi50J2drNXwnBk5wWdCjn2iJMnEvku
Fm9/Oa00mHiPU4B6MFyMhqs5VNL8686nKjBkKmOIXsK6LfToo/OKDqLdDupnN26q06GLyD1l8U7q
/3+6zYFhg4qAhiefQfPtnMeKL7VA8rtQ6ailChTHmzWVMKnfSwmPSH9s+DDmMMTwnyjUDvcTqPlm
aqTreftsuSyf1jDmbh8A7+3Wl+BjedX5zF7+WmuOgXu2d7wA6ZjSgXpqMpz+aluf9PNR++iQjYp3
PL/aKy+n3FRRsAwr3Lm99YHgq1VqjJai16lb9m2rM33jRUwUIbnFgLK5g88AA25ECWYgQbXFgkvM
4gbTVMuCkrqIdhpK4XFraLQu84Ehz4ivUFZv0mZQq2Ct6zG2IfWT3aIH1rwJc55hyMilJU5geOeD
OVXGc9Y7XBNABhFFlIiUJiYlyBNOYtLPIghXuhTxmlFybX8ZIRt1JRBe1NP1/vs4SbBRQYdV0ljy
AaWsOQUr7vbor8oEez4JfmzX2TLjMTWoWwvYm9lVlA28yGXa26X1d7bPHlrIXqIdiNYOEl+ZzBTe
1QwyO3FCP99V3jfCSy0DVDMnXfvnspNSEm2TRwLOVQvU6QfQbiiTeHpI05bQDgQnUS/9y7EcYzAG
07vNsrzWIQFrZ1nCynd0Vlv11ad5XSbSgEWvDLVL+ThTDL/TMjnGJdI4ErR/GYaWfDduxsyfPQnO
l2BJ5BSODB4Cipo/kL6X3+A9mjpUVfIk5h31GpxXGfzL9tcu71U1M801SnwRZkt2r/5G6EHEsx5y
/RvstwAJPiA6yIVK5VNLad4LdXgFPvcxCSqkBx4u5KWRj+88l32GGzWbsM6KCBl6VqxietQgveZ/
yTGGLuOW+/OkkrruuXQZgt2WBZ8JSmnAf68BQ8TfjN7p9XH8C3nymsxxO68xNC2oAqHhgNCcicNO
K2QGumww0OFSIFd5fK0hYQSmPfzGS7rG9cKxckjDfLbcSJLCARRv6lkgqw/d4zVaQaKLlmbDLBJj
c5ZoNC8tJG16QRxRGnnijDNfogLOqUsCqS5o++yNItTBrcZGMu6tFdXvYxQfCGMqeuVJ6bU8wcQD
/h5oyTX/3iiN9pwAhOIuxeZQhAhWE7h3o0h2FolkElW/rEBl+fel6T8tVTu6NtTBkaK1qBl2VxoD
uFbIvNm5EUjn3rBYm8DcCYmsJPe43wbSj/dMlmnd46uhmOo/V+XV9KQGHirhADaMi11nhYOBwLma
06QRLyt5FIaRyoYgV4vNsToqc2JH2lH9Od6/F01BXweVuQS5aiVqhfqSdqGyzDrrQCZitlZ1Vu0Q
DqMli0k+BPTH8KlapzZcY9J4SFmf7GuWVrgcLNaEM8DG+sN55GDBtTQXFKWfa7TmELatkPfGoIhp
DoIamZxG1JH8CuXI61qXZvIXSoF58yTI4yRSLexPfIj9k+4bB1YzBKxH5b4Hu0Arh/+jqV13KYri
wvH15VtqNe4soJektRYwcFGKdiBn2fuoBjTKXBLu4RdNg5Lunpa9sFw711wChEsBk+vP58QdsqVQ
+NapoB2MEBkpRLvF780m27CZ8meZOQpRPXmWIczb4Qxk2SVPEe7flTzwJy4+kg/IBoSnFoBjdEEU
Qns2UoemOoqCEkeQPlbO4a6c4Tsad/bYnoVhyfbo80uhQA3a8E/9gPegbPYhOglWQUNOAdTyecuQ
YOcHCc2lCwNZuLzMamwtbR9JGfQzIHUezdo37/lqEEyVepEMu/LRfipmirEGjWr/AC6nw4kZsM2o
khMJSwvhYbTBJ2iY661uJAPIjU+SsnebKMypoFquHQXR4JLmzdhxbOqALghzBGDp18rkwTo+t5Lj
8jN1ns2Z6siQuxQuOoaP4Jsb7wiQgB73+pdUu9j/nrDE//sdNX0JCPZZ2fQ39elSpeIxP8MSpglw
9SKBlSST4HwQbNmqk6YPE2e9TruvjkWiuEbVPOUDwI90Dv16e8DkgZQH8lRRQDsDNeXcXt2vkt5l
sHqf1ZHhZ1lQtOgvr3LSwed/pxoSpFyISlOXxjCj/CuGiV2kfxk10qSL1AYZRP1YtM/OsUP2n43z
qxUsmQbekMY1XZEawM+r/BqEFZBr8+PpCZIdFbdKgLkGGYjaNSA3RJjjjJPIxnKrsJWd1Vp7vtep
gGDjax2I0iKuDQwcwk0Ty82sFAa7ykQ7gHQXCFeN2IVk/o295jcYrQDrvOPeZJOrdjLDTJE8gcTV
Dz4gBbnCDp/RhOW2IF2Mg2d//qCAoL1KZeyETuXYtCgxadXFbQeZDLLkAaHq/+IKzP0uF4E92mdR
fFLXZuXSWvuXtjfl/QIEpXEeUKviaI+7JmSP7R5ntXbHprZDJXL/uvvQdw3+GsFtt5IyCXa9fEno
UHlOdIal8HwXEO+Ucjlt2mUiotLxnUMovWfezAFsVPI7Rbgs0g9/Yz8fR4Zd4sIO/4THPlrPHrhP
0AiCP8RRTgQygVGSVMCLqhUYyTFdAbz+VDO+eC6Khs3DBupDUhH03urxok//QB/bbybetyAZa5uD
HcxWT3FKhk+FmbLXx2mjbAaE9jJbjNskIzWr3lAPdWhn6DVkVj4c0ZAS68WdtVs/fNlXtsPy1L0A
vnyTELQoWIbAGW007FFGBi2kbxHWoyRZBRwtfYLVdUfBrYQ0M97Z/NveHpqV2meXO/qh00BWia9Z
n/wXSVgEQLLTg5jx1byXKoJRCo4Nd/VSTIgfKG7zHFGz4VFRRaAt8voBn9IJJtc3b4txZDyVKYLU
wEUOkmFfcLiM/NSjY/zsUO7/Hjrhw0DvRYR6seX35ME8mgh+5BMcLmby4kNmvq6o05Dc5lWgY5jk
kUslgJiR9RUzkHGlgoKgmVOUpODCHp/RwfO6oDH1Gw6Dm34xjOYIVnJtXHlC50RNOHMhbnGZMUwp
Txwc+CZORQeJgV0NORpRzP6QEA/mdIfKtd9zNwWIPZfpWyztwWONIV1Knl82LurcT8ZHpW8dbFhB
l6oJD40L8ji9Zng3H5O+/OSD+6F7onhlLnCKGxeBrtvH3G22pG2NArK3IuXBUrj/MiQqLm9XHz+G
ACwvkhJF8jRM/rZjmfHOO8ZVgh4UnGtcLPrpKjEVnpdAn62Ok9qZFq+gNq3H+aX8PdKQ2S9fAuv6
lPhWq9eXA/oTwB4WPeLTWtqyLYKMEuq6v7SYQ69nw/adYeTE8Aszmzb6R7/tX3xwvR0/Mp1sG5uV
q4/zLX+xgnNHQkqktLDN+DYw6jJ4957BJKyhsPRU6/quuksokttTsvyn+TfDoao9dimPr0alY1Tc
LJnl5GOGARar8UcOMJgkDhiZPx5xkGdNxEC/gOwmhcQsq375rXlkF+BYWjSP5naJeEmqFJrBj4TO
5KFyBLgpt3gMkjyjqMnUyMc/sil+RzdIh7Vwo9E7iwpR19vVZnNSx+bAmoaK1m8GlBCOt3v2x4Jq
nSmzDEXJ0DNAioD8Vp4zDXxlP0xxS/0nAFvGybyUERo3F6BCwKI3v5ONIRXcLyFVau9hzDn4tL7H
FdS22uWFerW3EUFiGh9Yxbl7Nne7GvWh9ZA3Y/S+ccImVzsmXpuGWhfPKWkWDkvML2nIgwRja3bY
Amw8KYnIEEicDBx8bVwzGq8mgL7Z410dWBFqwvjhY6mzcgOTsotx/KmV0syHT8yEGPLQ4SWFkctY
1M6RGPBGXuGgfmLWh+8LYxKUvs3rUS6JS96XlO/j8AxAB00Lv4cNj9d9Cc7hENAfHlPvKKk84tFM
/MCeh0EptCS/AKgJ798N9HMGECenqQ5xZ8iZu3TMHU9ac+VNzPy5wBVwqZs7rm4LF0mmvvlaDtc5
pqQ9aw/UgtYL9HZAhF6l9iFiKdHFCvh7d5+kUYdGL5hHhGP+qh08B9DJSpyFaRHJIFHVwSI//9rx
0R5vfyvjl/hTnoUIzoIItQnwAd83cWei507ubZEsdhARdlHP9C/MIAFF2x69oSVRSr02Dt6rxYF1
TobAlIYY0RyCzMuQiNhMPf3KrEVGatJ/2VuPnocwgXqUTvuyhHJPJUc8a4FKoMyxuZkzuGHAeIhc
gp9WYuB5bmWfTNLwL6iqCQE2HE3cVqXAG5Tn2y3ytUu0/9vhUzh6yrfPdDfRoVFbSvwpnpeHaI3z
72bb6zG4FDeXxoFLaaby4F2LowjtWnyDeUD4VwQ6zIxPPYIgByb2Snxtz4oZ7oblHjskgBancjox
BQTIKKTZj5pc+nWxm7R5SqPp4WLqi3RDx/VXWURmhOhR1TB13/2NxlDHN3riK0BJX2ijoxP7a61r
rw0/XNNM3+XjFoN3I7ZwFROI5GVzzpjinv6LdTuiAFOU4hBkbIM2UX8GtlDpH3vwG0suTdA0ATiI
qHSg+JWAVE5opyZAKVYTeHRrKFHvotB1I0QHymfwTX4DTj3Ll4qjJZBFEocsRKXXrHpbsOp4nTYj
33DKkw6Z8WDzeivFYb0lGMkCNwRlfJm8fU2uao4oMGfznJwLbtajkDU7gg53NqyEWmKGIWBXic7n
MGdgv5Ut5HdbBhh6x0NABfboCZzL7KCVUFoXBCWAoyNUtWHQxOenJ08p8DGJTcoe3JdIRcBCDGDl
xQYzvIFjYdR1xfTmSPaXojJZesnLkwwYeHGxNGQpATNmbZjdWkBBqQmhnVX0nzbMjPaAYi0nVqKk
3Oi0KW//c6Z/JImzzdTBpTZAD/1Q44JelASHgt+n0uoKsDHSqfVV/o1JI+l2GEAkP3Yzj1A6d+z2
ZF9L40H/cReo+TR5LjoqMLWhT6/HBCJUgjYleDEn+Jpxe7ccQXoIqzdubfSQncOedZaw6o7natBs
sIuxULIv9DSjj3oZpG9BCmWwcdG7Ij3HWx+xQTIl1GmPuyNkQupmuN5uVVNjB6FidOoVnEfv6tNb
KKnI/KlloIvAO2mahuSw/8vhiOahpt9jQ46Ipz6yIV7/pyGzmesU9nTRhtf7PeQOI/joowZ7ocbk
rz5Mmymg55Nu7uFrEOmtr0ZofBpRFZdlJm14kpdEteEnHvOVEuEWRrLnSFGcmnP/2Y9YszqqyzJk
BXcTZvzq8/POiSR/OtEfYFxIoiAPwstQ0rt6QbIzdl4pTZf57e0Kje6Rps3RERziK9ltoCjmQFKc
hIzsG+p8z52q54UuJovar3pSFBezEV6lzhnyNmj+vAHzgfYf8zrmttShQEoOqN3PpHqLaDASIVQa
wgTwcPVrbzAJV/FRexmNg/HzBVL5nZe7YFVnHSFvJUIPV+dkUVhE7eOxwl1U+JqtyMtWO2Pm3mU1
EyHXG5rXiTVdLhLVCx26m/Kmm4V5OgKAdCMeJUNRfGdW9KkkZgEt6ibUrvAqnv1e8ve31uZvtDCP
zwiQYAXY05dd46j91w0EYS4rweUXmyLOGCPbCtRTA7XHjdirzRaOSPEkdtuF0khfCSsyAqYS3ACY
5OGk5afU3KZmZrPOhvARJFu1yG+JR7wgy2D3D4PVxfpNTDUsj3uL1y+6bQ/5ykAlgJXyqm9vHOxB
pMRnimhIfJa+he5i6AOxgtBnznirFNzjBErxZOK6FMELyWetvguF+WU0+MemapEQP73r315BpOho
E9HwQXbrNc5u54GtVG6b/0jBD71tDgYlZHUlc/8YwdbKM/Jgn+7zaF21oJTzXGz3F+qeyfNtC2KG
XHDjXWfKcf4BFHyjlikbG45j4WeeWjOtEeJ5e5P87fqg512LNkbwbYV4L2OzzeTbfwFezs/YayOD
IH0XN6JbE43Be7zcKP7MKaJz4HHxoyzH1iCz8nqEwNFs5Gbx9NS3nF8CAwkTlc4Nb8IF/ILQV2OY
RIKMCcvnmTPfrKmlx5cvjjUrFRIDNht33KBWoJYw69fCYoaI56O30flBVr8/PjaCnV/RPLrqUXZG
DA8H7F6LXV04KnBIuwwsZdduLoV/epmzOeBCvLzKAAhMAlrgJr2WFJi8cOUcEuqW+vl1tM9jkouk
sYEghPZq9lWYf70Wbce1qiiTEcDhCWyeDvv9CahLM/jGdnsTX/UjIsChedpfQIv3/ye4lcEYPHoQ
IWio6rJyuxzSVA9u0sfUvVtgkzAtWSuGPilZZXbPNXVQ468QVz+rHeTQOjN+0ZtggiS84AyGe2cJ
4WJytnJGfq9DopJ0VDtK08nzJl8CmPZUU815DVdXmEqItoiI1gNLOfRq+6mli1JVTffXbljV/rwj
BYe/mSaHpvl6xo4z3MizTBRoBnBi7UL311kAfIDiVGl1LX36KsiN+8QK0S9kdyZpr/NPHvzUT/1I
meNfv8SQdbOA7bKPHk5mRyhNsU8/OPpWRIoN3z4y+4saxMHX7YHFx0wj+Oz4CvZ/QbYyxu6Slv3o
7EOItUBnDDZmIwd/vfmlyTIfE8BW22qxFBeB7c8GyoGn1XPK428H7eSDi74H2Fuaqd3p8pbA9Z6Q
3vsOgJh3aK38Tj7Bg+4oYXatNkPFA6RvFBtI29PMV8XhgZhcBNA/N+N/EXQ3CU3YNx3uY4uBaK0P
BPouUnSXPF8G9K5BKpfNi7JYTjjFYuEsBjmdjMmOnaSyZHRDPpEnB7CXU2qCu4dmxmrUT/yJ/+aG
LHptDH2KjsCtVVR2QG3aROjg2WWi/Zg/z2IKrhbGuNE/JDqLW0YS+724hhMaMScZ0kyH/AN8EplA
3Fee2P0DBrb2oZ1u7Kbqr/yNN3SfcYC5MacS/QqfS1pwsjEDy51g2QsfCSUr6AubRfDStjxMdylu
YkSx7Cw6z5D6+7O3b50LaYiaDT/81XfJBDnKPXL0XOUiLYto+/okBv12Bw8HhUsu7lP3UxKOzBnM
o/+Pd/IRaC4wo3Kn1iWad4Le2NGScdJp6f7wpyP/UHOb7zL38uaZDODJaEMBLH0UAwqk2mXGNyDS
L6J9F6iVGsFVOH+900DYaoBewfaAlTuPtNAFXOWqbwc2ez7Xo3Zlv6pOHE6ZsPBhel7zgBWtczTb
QMI9OOE3U997jEpiNCF+ayZMWDHHOoSalPsrKrOBYHAbhoVDiw7eLMHACLGxNUWPYz3SyPoYBEjR
WWPQkAM+KitW8nnZU+dVNdRIImNVCpVIpoInDN6nZOEBQZVwAAA3sbhs/5uPHLEsYKrxv0BPHtHm
7UHXtXbPZhd8UoEQyfGYsT1gCpFdkFEuF/+2p510BtEjHpZmz+yaTpW9kzN/wJVJ8Iox3XIzSKys
D0aE7p26KUCF+9CyXzMyp9mn/OQkv5hsQYtFBR5T2YC5yyIyeR7NPtHu0Xe41zNYUNivF0SA5fBZ
ujyyk330Vu1496VozyhZCXEFTc2BMbG6kXXuGkqtBJT+xTxXH+Z1zgA/c+wF5pt8ZlHTg8cVP9PF
bViVPCeGoxflh9YZVsLxfjq3wBVtPEY2jWrgg0mIUe01nDszQyqtgMQHJGOyYl7688v6s3Vjwune
UsIh9KQ7uRmBZjHQFih3W4qLJn1DaChysKph000HWv294PZ5VGuoS1uuuXQFgxB8awbrbNSq1Hmf
kJRLbM+IIjB0gYMwJ2aQQx0IfvzFghVg1JLwNHSPG4Mb7EKq/gfOCJwwjRfaagaFl6wulNhC5JgO
+DfdabKDfrlaWn14igfCwVFvGSpPQIN51RyLlSos/T7pGSppy19KcYKtm0X5cFbPHbnxau14H05U
U09rUJDEddwRAMaWXjxVqiPoOAObifWrU1fcF1LSK9O/iJYsv/5KEnYIb+YBrOPsphwMhkoyUrIo
8UFwCWfY4D/34d2An2i+FBw55gciBP7q8fIhfN9IylNB+tvE6OB93N5DQaWEHSu0uNljiaYMUSbg
P1XDF7xH4PJ011RPZ6RyiCUGDKiH5JpHQRT5jlC1CPXl0nt2nIAO9e+MF2YzYECMB6jleAkPgUu+
ZbHoyhY3cD5qAPEQAoT0chYYIiH85FqaaAJZXbaKoWPyYbVBfFrFNFk6ZQqOELHr5NhsWA81oEzg
bLNrmXHXOFZ/A5v465BUd02ccRPJVuzfticPSf+x7KswVy7dOlcctPJRiWOy3fspOg45Sl44LBzd
KZMDXkKCrAYOiNmev4v0PdVz3QlV/ZBw7jN3gdtVNL4kRU+ea5JR1vuKDy/TVIoPeGPU8HB++IOp
915s4zrlqmx2bsNDkfe3/jzw6+4CGGYiE1Wn+2LbtE6KzHLNercIhyXaXQMzsZMUB6MgUS4T02q/
ePs//vL3JiV1pkBREoLvIUpXbyhUCR29dYdqVEi6Y572ivB6DnVZfp8L1bE1O1GjR1dzvMGLOKce
W0tslsDcEoLbjTaNmB7ch5XSb89D7Njcj/p3VgAIuqJiBmB4DPChsFDwGBkfy18VY+XBtKr5asUX
+cTRaNCAUTOecykCfZo8XzbJY4Z8TjCkT+ysO6CyBTOvItyKX51VNXFKQy+1UOHmRPbHXqcEe8W8
SXHugDWpfeNzes8PuJX6ZQqDObjNWgAfSzzY00EepcJ6KrAseVWkflAeZyAo8FefOb5Y1/ZjAW4m
SBmG+/VYwFKwEmuVtlz5+BJ6McWe2l61ODObLxYQc374H6HdtmL5pD0eYj24sLbz/Tej6Hr6/ep+
IrJMUO553g+3I6Hj79ogFzXwuoKMI+3py580ZsylWKCDRCMtDoo0jHn8aOJ1pCpu0yKl7tF9ojsp
55a9kPZJayNqkdbI6jNR6T6k1jCGZxL7gNDAt9eT+lMhCZ2iCH/FPv65O4uZWRYzfF2isM9N3Mak
drGPMz4UZAQ8J75VgI9MjKyF0/Mg3MYo2ln44jW8tdnwlFgoFAO7/wU7+aLsiRQCVINMmqfyMTNV
A40Rif3epmFRRt9DupR6xRLUtjERSb7qCyFwqTc14FU7cqvQX5T8YT5AvVHNp3q3EeAAtvPLT1yX
r9/Q/yM9cpw3zhK8ruEWcODw7n05vdo2JkESqzmSnSAglpz3SqwTjLeC75gfKazpe0Iat3rUEIL2
uxCCK3AfzlQ/MVd94l4d9nPdqg+AW4cZoCypyXL2aLydYHE1XUIrQmc533meVPWFqn4UaZ2Wg0Ov
curBk2rPSc/Ne6fgxlUngPyuwL/IMP+ITmXJ+eJSm0+Oveodbkzf/rmM4EWxo+pIPq24jM9zY/6T
taleYxPQiFn76doL5viP2OcHlyEH/q1+nRfsXuyHJBXpF2XJaNxQKx2cgfB/2Ubi0VNOGxLq+BT3
risgWwZzKCPDqwy0csNCLLYQZiwYNAThVsy6JEF4iFm+inbYzpw+pTs/9MLoVuzF5fODnGIBlxSX
FuvDM3kliMKaVeT8uzZJwnDrqiyGN0b15msGPECHmSPxJ7s8SV5G0hDDxOnQ1rRezstax3Z34Jx5
LxivNFXh+BaORkuRbDSJaysSFcohwezq8WkFe5X+zjUJUZB9vaFNJaq0il2lYihyAROsMCfjLH4P
8LLiJ4PjK+1R48NQjELMk8UYOOrKIRXjcAFvrqaqYepQe12z94XG7mR2XAdVSFA+Gz3Gay9wWcmb
zgNycqoPRZ7HqJAyoz9C7xO0gtlK0rxt/Z/iR7C6nX1eA01EzX+7DS3Wc53q4N4Mrgcj85lyUhWI
E2/oclMJcjCiTiCesaKInVCrqzz8NVq4yxcBYoj7I1tOBjM2Id/zSMesdJvkDHmDAl2slptIQnxn
evnuWNhfonbTqM4drzNYLwqZOEvzNBl2h7TH7vN3i9qwDOGC9OQ4WqOF+l8lINCapKSQwf5DAmb6
r1xcD+FBsAc/x4Tt7ue0ikI2JzR4PkspwRkhrWPrzKoLOF6gp1RHezMjiNBNu3QKLFJhmnWkj8Jo
7WxR1NNKCQG0ALJLZSWTMAigb7gmQTIZx0ykn2Bf6nhPT6d8cotA0J8jS9A14KEaQBFZUjMcxnya
CvLkrgTVAO7BIWG74bBIPXjlw/XuuewjJJ8OylI8KRxM2EQT13tRUeEF8pMaB2UEO9VQ0qvNKyqt
WOXTps8l+CqOhtBtlbXxZdCQNANneWCuN+DoobXpOEwgbSfuBHpoIwUyzC281uNHQpI6va7bFh0d
5JojpvbS0foUKqQ6/oRcuGJk8Gi5WAOwzpSbZ8zk4ellDS6NA438LWmYq07JFqagaxoW1vNtSGBo
rFysXzCJAAyg2eCIMRtkP7V4MefzdzYJti5dcWN7NvOo4Q1yEaOFe72o6p9O87++koWfG9FsOzP6
LYktU/O7EI2YT6HNv/UWS6CoPSO1kif0VlUJgVBLE1QxhAQpbdmuWjaVNE0S4/BI6ImmNmfrNoSD
L9+ehS718HkPUrqvANEv2Xyz1raQOKP+6ETknJWhRPhfF72c57fpzgHRARM+OJuG6bjmW504tXqc
+TA8X3oLF8tNSjAobUkevM0ALI2Dn9BXXQtIUYQ6lhZEgJpSHVcPhad3yeToVaIA9JvwYyiYBtDk
0JPFp8+AtAHzUGVv/Dn6FIruCLLRnlfoJptORhwo5frYFus8RmqaaxGajnaWpvBDY7U5vbas9gAp
HdgNGDrZ9BdSt6eXGZSlPBAC99M0DvZoh4XlW41McxEZJsBbIg3aUUPd3eqCq4ofpCM/m3xQ3PeQ
6H7CgfGiHSinsmKx5IRtxtyRut59rc1bOhYGTBMqMDt3QaKtt1k6t09ajpNCDm9phrQhd9xDNElF
SFXeYRz9NiQed+fkVYVqTkSbnLEYtS5T6pcI14n/1AceDFUFfEWb5POD34D7RAl/hmgnrY0svAf2
7jpe8LwFkUiDunRVYlu8l6ipohZSUZmNJUUypv9xso4Fu2rjfkIOPQgFAY98Sty2AXxRiYMenHih
HM8S/QAvbCvLSQkwXfI3q8Kfcj9ck+jznBU4C0M9hFb8PI3s7IyXEB/Qn5g/UJzFaSjxDz6mpAr0
LSRHYW2eNfAKG5cCWQMvVLvnuGpM+1XzIJmV7aRAqNAJl5AaTb628xziTau04mdZxSoIxbHxItV9
pJ9fXQ6JGjITRAL/BTuZogpiZiKeiPrJEr1jWLMGQjcTCfdXv18XJkEpFK1ILQX0mlggJYy3qLUP
Y1cqyBiVe1whCWAQaAAZjd1JkWtg+hA1VhaGFK/tHOyN+Dj3L/W+QiVOgwPjQEzDLIv2JzDiM1NK
deRzIV9bPRerRr5t6oTei3cBoQJVzlQ1rpavMO8LWCj8/5H5RTSEMcV1L8qnKOL1Tnd6j/kb0Hov
WriwqZfT2hXqxhc60aZrZbIzLc4Hy7U40GpI7se8/Aw0Nq7EgWaXCvs/gey7jFmTBie5byRgteOf
w3EJQyWScSIM6hofJL/AhyXnvXwZBKhOEYbLAFLLe4He4epHvW+UHNhvle0u6auq14WazpHwWOz6
GZ+vLlFNvakZebllhKORIm4x3AA8TZam4lLZaADZkmM5gbuS+fQXnHBjCpPG8768NZ2hqktKByCC
lL7lAPJ9EqMJykIGQSRIjitoqV8anWToaRhhrgZ7BCwhgCHYoi66LX6LO/NJazNGJnFFEk1acxIE
jNqwaIu9tgVRJMnHK2R1A3Hku0+oY6tXcOggrNlsV5AXKLbsowR6OVc2pYoZR0Sf9wWUgMrA151O
UysubRgCjuvGEk5ChBGauJsePDbKmJ2kseWB12nOvPS4S5StYdegsij0mGN1ODRrJF6Wh/tzv00v
o/MOlVTuu8X2M957YKSZ/c86pJu1GCJH2ndUkSSSuHfROQzdeZxwiG/xvcRNGFmeZAOx1pKp2Eo6
itt6yZabCM/YOHUQYmJcl3bg3EPaRFdygleoplONeMpa2929N2qAH5BGAaWSBCGHjkp6kx/SURdM
SJORNpxDpOZ+NyRF1FOjdbHe7E+HXUvoEaxly0PClsXz/WUK2p23jktDNelNGIiNaHVlAZaTiMd3
Kfosm1YBNMyr96fvxdlzV8jpIEaOrJMUnGrE1NPlKOFQknR/Ovo5KKh8bYOazRa7+uxLRJyfz7s5
Yru5Mng5CUUD97X9Wgbd/YszA2Q6ctzaEeizZs79zUNaHU7nhxG5pURN3hy5KmGIyz64W0fvROsg
bOYJOqoGIwZGYZZJZH7OaA7uvcNo4/sWN/q2OdPnpAGZLn5vtoNeiEpqdEud2SUuaF/2xt+FP2ea
sTX6OoYk8kyoYPizNWP5DPfb7EfZ5hPbp/kaiSHD54LXuWbsgzGCS+17yMEda343g5ZMkTxID2Sf
Esf/QNyEZ3NJf0i4qADh7EGDdb8MJ7WSuTYcEhNS4b3z37nXG2S+VcFlAd4FThzH9KfLeFM3nrbH
waVaUg/hxufrSDJ+EP/lKwkEKU6vOwhQopEynGfedc2Z6xRXPfFqkoGuHHd930fz24kOPGPrUN9L
niBdLnVjU0gHFo0YMu039/+S6+cT2u8n+c8Ep7+ZJEdoWQ954wjQ4Q6O/PtGQmLju61ZPjclLnF2
Ut4rOMpgboR/2nLZqt5JaMAv5GalunGzCy1rULXToQzDU9Gitm0t/CQ7BHQass+jJEiAoJC/UU78
V56K7woNbWpat48MMWjdElJuA2U7acOFDKohiwOOiI7Mg6npJRlwQCvxThzxa6eAbXuF/pHzCWY7
p3/eyM/z0/i+Rj+KvMhcz6QD2hqO7Ocvu5cb2MZfuD8yVGDsCjOXQrb3GGYnuYMppMP4h5BezBmY
XoLu/xG+EmSRP89lAzXx7FKxaD+0/C/oooyo+BHwsZqRIA0CCZiZJ6+ZcjhClm742p1exIafw4fz
+J6HYxITUeAN+5dlyX8/5Ia/nG+Wz3wieOuHP51e8RvQRqKoLfw3cHrm/OCKXvEOx6xap24O7eNI
9noZ5gZcJ9Y/hc/9t5Xbksw2aTnsEwYzdOwVCt3fXHt/uKHZTOQCAdn0+SMtpkgjTE7M4SUrQzzy
Q7uHgExVAwVgxK+pZvCbHc0IvHMP1bCtsULL+43sOOs95//Hh+i0rzXm1cyD2Tno8bW/UHhkxPyE
XLvrHt1N/q5ZmA9N7hyNHsB/zaV2giCoZvwpt7K/PUkzqSi28rnsXLo6qRjbWn2yQbZi+9nBvQR3
C7SWGuUXhmwZktJ3N42KvkUXLacwLV1jcaOGm1WbdyrezNdasjqBamRciETYCC9tLqkAsvHExH+1
34BLJULTrXTmKGGs9bmPlBdmUylY9Ou7ZOfAouISjpHPNHHHfTuErYaWHu2W6giHC4d5DjbRCCMX
XT7EH8NMYSwcUd4Tl1CPZtwotOw0bBt7fd+hv3zvJLsPQaSRFrS5fF53uCEtKLc3MdBcl/IvnQ1k
39A3QjZkTQtyxZsGfqFkulU55vl2YolnZKNBZQLKe2mhFmUMsWKlO2OGSXraYILaPp3qLD8BToy+
3RE5l6j5MJ7Ct+TNui3lT614GfgMPyDOzAxA2LmANrk8mgKsiZH/a2y6t2nnkBPjm1Sw/hwF73/J
IE7wvNVwilChpsm7gf/G+mnSx0MSjXHI+ymVZdSHB/+IWihCagJEcH9nrDL1NuGWeUxxP945DDNj
nMXWoXz8N3qhsDz0AC1HLxpaYnfFubp63193Ei561FooG2wKr/YCuz7WFeF0GWUkQ5/nVLdRxdcV
hDCYICvII8TDtEkqsdTTxaYTqrY5T92dtnu1OeNFBpevUBl4xYf39xH08HqZxepc0Et4i1dwVygA
WKPMxK1y+XfFt0WJqbp+CFYZDNwMZT/NJkgUeBQ9gqS8C1cPdfRCAx//mSehAA4eZucxAh4PNp6U
4zuwlkKzih3JzOvq4hBkAAzeMFrVKYVzkbtVd7dWolY4mDA9JSFYJ67/ZhjxSUDMFJn/LJWHHluz
BBc0Ohu+y9R7lMpCO2Zjsi5NL3hQjOpaM8EDYxRy3dBsyueQhahDeGZNOCdbro1X/Yyouh9q1Fw4
fcXW7niUXFX0ncA2LrjZKvJR0l7IN44te8YYF/MUQYjZatR2cYwdg76Xr3gVNMv7TG/cxKFhefqh
itvufnoyBPF34TJ6yzd90K6YHvp1rmY8RccAUKe8Cb2ib/ReQV38tSjXV7JGtaEMZRkWghvLs/Ox
ZK8j9aEyjB3Vu2qsVQUIjSzgtsD6dp+dofaqp1UJuafno3Zz7rrKtoMeG3rK4ru/JgebJLWaQmmj
bXD7FYrm9zKsTmy4ajMmfclA3qfhbRxgodBrYJrZw52priEiCb+6pd7IujnLPZlL73O1r00dHbbU
NA3KgGpzLDp1e2yD/a3E9F8+TdqLbJy97LB6r0ZMdVsbYx+gYhS0K9EPPf/eIPdgcXIeJA/dFXLL
LrGL/YzD9Xl3v7T4X2gbYSMczk62GSzicAz1blTTsgvlC8HittQGxsYE7NZWBieXKHyJsetD+Kv6
c8ydIyb6SeBtBeQ4cI7mRRzt2X314Ei9zlSu6i5JDDblEYssBo9hitKtvL9v55Y1Z9dcihi8VqnC
YIN/balEsIlsp9SIWi/GATFCROv9+dWYg08ZjNF/H4oOnq5kljn/XapuMZZ7wTZxCeyP2F3h2Qar
LjlFWKzMbebOe8MXA8sk2W+xqBt36GSfaOlH17PKVD8OgUxHzc5VvH7MIkEOkXaguqcNFLyL4mU7
/UE8hnXGZG2QYgDQfz7V3EZ6Mge4+VrCWFfcLYqnG+ZIAa5Mi8AEJfu+FPg4DEVSIQHo3xiNu46C
d9Ts0KyJoeDWbWjUX0kZCvoKVqFvVJSILyLwXajMRFQ4iJLmFX801oV7ji9joF5QfqJvAoxp/rVI
ojBD6QVJmhIS+idAiyOjMiT0sBiNQ1az8R0XASWbLhjlvVwibCK8zvJgkVt95PCPtp/NVO1aLCyB
x+AI1a10ZOQF5WsenccFtumhxzEy6zgn8eazdUO/loaSuigvhs50Pvh+VbDzJ+zeCfJPMoKwcHR5
+yw5GhbAmbbxcFmKZ5h5wT8I6kPsfRDUUwbf+fMB9Vc/VAIjdSHnBo9ZXhijbMzlOmE6FNKGkb4Y
g5Vo4RgOf2jQnTdmnFfJsaBn2RbxhqOjQc6lyXrKN6tYcIsp27hrDUMv46PZryaqYuJJZPlORgVH
Ydeo+Z0xC5IfJ+q9SXD8ZoIdElNQce1fgOL5Qbr2fo8sFdc/b2aAFS8Ajna+TEm2rOkh9SrPbKoS
hFfZOsAd7cogfvTaWOqU/7P7J8aPbIrlhJMRaay8VdTXslezZT5bPU88nqmPvI+FDA3Ic1KIgYuZ
ktul/f1cLA8Hvr9Z0M4wFmI21v/bYJpfvCOeFqck+fqF0+TL3krpsGbVp9pX8xiGTDJWpYtMYl9p
xTx0vaSOrixjnf7v+20cQ1StTjlXNqxpZELqlXgTCSBYx5kMLwbjRkHUl/Ofq8rOzpjUCS+a+v//
F5OLIEbVZ7w05ULzFeYQVc8neY7bLJ1uLivmJjyzqBr6cdPj+64rUfJxUuE4hnHh0x88AxdNg7E3
HI2Uv5jeeytVsXxkLbTSpOqeI2yAvFrgPZy3aUTGtkq3v+yVbecRApZGvXYoirkwh5fxsP+Rb+aY
BGL/87JCDtX67oQTPw23RLcXIYDULVZ1l2UcLfWgyyNI89BUarmD6ddFVncp7YphnCoRAZIzui/H
/3fkL9de+xABpaRXbExa9mLlqlLNwb53/M2ViKfcoDj97zgA1vQDZhYxugHOC7slrWzbbeRW3Kj4
ZzY532vfgtLxeZeKNJhxtjuoBBtBUreOhgFurkW8XVnRd7T/u0EE0iWP2YlCk2GSQRcelVc9DJYH
3UYytFGf1aBOevJKz/4u5pfLxujfoTW688iFOUEyY4wCGVdp0VbUSv44lwoGp38maRjo+Dr4v7iL
fbB5nyx7hq6+YdPqRsyiNOROu+xJDPRpmHCgoMMP3U1XQYJPzpujE/q1PvJZQr9/9taedo1aD/Mp
Pan1ner0Da4IwFY0veliugWMep2h5sBmfSQZcEXRLcu//Y+Gz/SVpZ4JU0B+XRitsrxRh0xGqb3h
OjCFwy4+7oL4IsGKSvmhqeuYbKYvnbwJA5N2l5H1PUop8cVPnWF+s3Tyf8wAhMwYoe5LXmHTyxRS
kACD3zApcP+9tFgmxhvDtSoeuju8bgsJRczdrO/7bT66U0hEZtlScIFPZanAnYjZhp0/7BHGAX+z
wrkNcQOYXCqFfpk6k/g1dbzvpeT8Wu4IHKyYUDp178vOGvJmHEy5llca+5s3q4MVlIaYWDtlE7Md
szvDLsOM9B5PPPnCnlUGRkSnM5J7y2IJcajxrYQ7VtS66tUG/tAx/4oC/ukSWrTMmczcrDNCp22K
7DjBCVuH5EGaRizIAJYlBJnpnjFPYeLPOli7yw78aOGRdvdlTGaeX34R/ePmWOZMbRvE8RUSoUsw
d6Pagnxo3wbnHWTwLpVAuIc8S2WHU6thK+HJdZJmVncpa5r1SFoW10S1jxWS5mesVh+L0Oyaj4pn
x5VmyXOF8YWPjPi7jc+2ZGa/Xr3CT5SRpjoN2a5nU6Ndw3A/F6UZjYoYTImas2vFFNYrek5xcx6n
AZuhA9zS2O9HveAv2tteLATo0IUoDUefn0zEdruwAmAtcP37MaoNldnCvXO2CHmVUr8Gi+87L+VC
uTCSMoH7DHnfrerh/nm4zjI18e8t2X6aICrXiG3R6y3MtH+mxRx6PI4uhqXw7NcFABx2SezMn2OA
94503js9fly0/8R6WgaVtxFtcqM55P/j/YNndWQSj4yjITWT5C97yGxSzODiD0MNd44mDsal0eXJ
qatK75qGjOCYZtYe1kF7j6O6VVv3XyqP7Z5GZ9/jMdgHI0jlROoPAdcKSsyv4raerhvokmmW3yxW
i9q1Afx4BmYONuE0a05p5YAfypgwmEMVcr7X/0wQL7kFwuRARORY48D1aSQiSUW+Y43ce20/PLzA
rYnukLSiXYS9djfzO80Gdrf7+8+/2MQ8DYrXcGDq8pSrhLQ9ko8AQ+3a/M97EskQ49jteljaG+St
BpX+7hDFFwhpI91iCrsMy97B2TSEoOGWgL2C2g75O/bKLUbG/RbZgskvkEarUCWBwiLqMEMuBIpj
G9AdtOLPoMKkgg1Cf6CSYS6sy5/976fksLpB+E9Q0Cq67+zAUq45mNHSyTDE/jJaKkkgGTV4A5wb
ColH0fjgBYBnRsn/zFo1mHQDGyKRs++r6tSxohBsDIT3Zgv3qid+/xYqzpbnXjruH7BKsNSBiNYY
GHq65jaPK0koU95gX1ruREgU+vslWlgvcjhj/dIbFqPoGNiQLKkuFXdIDY2DIgbRBiaNfClmVEYl
JEGiMVsEwMs9z+x4eGc0S6x+Ix6E3wJeMmH6YytdnGJkj2BywTPxApRiG/LB9yidyyRs/jKN9JaX
cwxnyLiP5Cl2Im73BdiYW73HoJh7Sh+z7AAb+Yu3OOr1ob7m2bRqynvRGGXjTr9AQW2kJsoujyNI
5uvw3YTfdpv3ITOUbzDVuFyG4gvSc4H178F41Oh24kXK6lhwjmKzD+4H0JYHaGSSMRMqpe5WIwdT
lXEvV5Zc5A+S2A/Fd4O1z7ezo+6Oes0WrudTqZ+e4kzQQdJIa9tTsG4vaMsLHlyUiLufHbpEvPc2
lc5V63ZvrF/5xlO5CiIayaIxAvLciqC3zk4mJUtlpAAyQp4lqwp6TszOPlHSbBfmUY2GNs2V+KbK
oNZ3w/VyhKTtOA4jIHeTQZSjNNw9lYRXtUpjviH/HmzFPfMetswhQE4fIXuu/Lzj/D957rmZs1VZ
AaMjyQrQfS7wGpOnOTngPRLK7S+S1rdOz/OBjUVZHwCTz7J1mrViKPDAycm1SZe/H8JYIooMkuLd
wqucN9vhgF4wHyw607R/sC6+iOhczYVZgsddW5wPYqdCuDOLxmuQE+eOQMJPmfqn8HCcB3iZTo7h
c0SJWybpU0m4jLb9zG75NYZfp0d3zCMCxtWESgWTXuRUK2aaqR+feV4XF4UioXi8I1wmbiNSe/N0
pR0HHDkWbUxYLQWrtp9gJVZATWLFqeUJOlW4+zML1Zt8c9kC1ohqXD4jtLIBvL8++jGf88Zyh5gC
G5U9DJBhFeshkWRkp0VpmxttApLFMyM0AgjmS8Wao0p73Zz3UDOdZlRuYtfcKHIzmwTtIT1KWS0X
Zo86ilAbRZKuXnZtvGgi4ObKIoQ9ybiap++ch63wR7cTDG8Mwdjr2bzlqn0hPK8XylCEauVkbaEu
tZ3nGUu5OZrr/0aCLoNhPj/t+JvHlAjKiXO/EiyPA8IxD4GElQH18I+H8y2yxN0Fy2uDc6Fs8m7w
sVlAlQ9CUNDajUw0jI3VMnHcCq0nus78gtUARKdtM8QsUocl2Tbk+yJ28/N9aENqYz3e1+6g9/6K
cQsY1mJr0JBawiRd9GX+InBv8P50VeZg6qGbPk1NW1dzh647vJoRdzMOQ4ghdy5N1IPzuHP6CLhv
fK2AYp8zkaEqLIQkWgvnMPBkRb4L8Qqfp5H/LNKTrKUKc5P2x84rA2Vm2Khvqe7sRqVaVDk85x+F
CPCxI5pRfsTIB5CZAzgNlpMo9nppbgOgJIEzwrC05AXhYE7UycWI9fmzYXr0Hirxq4mOxMMDGpo0
HOeytNlob2Cbbn2qCbp/gNSHXjxTq5h9sZofjrRv2xL6MhxmITM0WmZ9xUT/CDghFvsnJsegvwv/
cs+z8M1RwHuNDUyKSSeWea3drPD62Z+yXUUWlXV5JEzXzzRJ89OSulx5Vm5tgXcESbeHxIuTZSOC
GhaQbyhzsVcaPvQ/rSfUbiNCFujShfNXED5OBgHvKFl0m2qoz4BzPldXY6Sgj2WvmEWsD1SvMiTY
Gwb6yMuwAqE0VXFyxLQPNJVf8ZGLUztM/Ke/QxzV9E0zU/MT2AFRpThP4OC7j+SLmKc1cDwt5N+J
h9qSrpg+C8q0zPDzF3bNSYL5NvgJ4qh60ZN5GuF0q6hyZPqwbJvukz0R0PzZb27P/fiDM318KYxW
YWen2f++Dva8h1I6IsDM++o1cBRLWbuyngvAuX6t8YfSYqA9DWrAL5wp9R0RRXOOBgA2VTxVi3Nz
umco3tISETlCZV8AjsghqoGEKMiJhy7n+wve2yNhJ+0IHc2Jfla8GxjR1NvEAX21V0DoixeCJvOP
1au/tCrIzqVPKcJcwl1Mx3Lxbb6veCtGwzPQMtEsn4BoanedwBL8Ymif3e4z3fujTBdPEDtdJO6V
AVI5z/jak40sJyZFLIesUYvItH89Vr+kG94CyY9nN88DmX/fSwCl+gGcGQxyvwyiyc1QEHaS+hCE
m1JQXO7NpoGDnE8uTSKhLi11iCWJubYjvN1BpGKFbHtFxOPegg0wPONYYfKTfVY7XtqKAqV6Sfk0
f/ghYeS+5aYB0oPXekAp1JxerOeyhP6WeJjxeb0PazGkmwuRyCGAOMiaayfEU4it08VuONi9kZEI
9aVs/8rNZnC0+b3rN+a6BSGtTxMmvEsd111ZOJk2xknFJRRn4iNhCYYpvH4FnQlM+riwvWZ7VjAs
kOlhSeizsGKueg/NdF2wHV48UkSJB8gGBFk3FABsRc4LlLpaXOVkbmbQWI2IDNOQeuxGxmd5qJzI
whgH9cI2ICny3ItQoyrlq//kSLEVt8D1ManSfbQ4z9ygPMlHvca2GA+6UH+JI9XnwXYNs1H/pIny
+kJh8s6DmU1Lhey8NXUri2z6Y+D5idiVoO+mFRYxSiyqNaWtxriFZrdJlPxnpkzbTGfXkFxovA6S
3V85OYPMRQ7Wslfr8bR/XbfSk8rG48PSzVykPqxLvKCfHIz6eowem4gAL50uaUlAdPVXSAuAtjH4
JvUPVFL+cVwjORlAw1hA3U7kITD5oxwnSAKDbJ1E3kTeue1xT8ck6PdY3OoVi0411wfi5u/t9r6I
Lxhi20p9Rot3MsnLn3tv9tL5IM8Rqb7pyp2G3e6NvmnDVW1Io1PQHqQobaqcvLNgZTQ8XXcHW7ue
BlPe/A368bowL6US/BeTWQYj4Qi9ZyI/G/xFNlvJ8CaU+glrBMrzEsfr6e4xNA7scrDA/20lp9ei
zVRde7Hl+1PUyUrKVQFAT/xCiGU3DDgCNlOAye0jtKxquVEGsG4Uvm8U2lFN000pwEDdTjYJKqEx
qQbpeljznXvNpZa4iJDESr+L7eQqhU2xQPsjvSBsNESoyrutWBic9xc46qGC5C+pLK8t4eKYkSmM
27UxLPp0ok5eFIrImzeablyJKoH8hlCR7YEh1yqLUfLTSxv+in2eHrbt/mR2QeWDgw62Zoc8r+uk
SC8YLXSt32gFxy2P9yyN8OOUYFhbOUZmdEUexMK8eyG7NK0BAm43qEWlMwDiUOoULbdhZw4GHJk3
Qq1T9p0k1AWdgAAu75T2wQtv1NpBcEiYpI+y1hCDXTFjqUSSyyKg5fZh/QtKhI240ef+nMFzsovx
pQUMJIIMgXgDnCrTfVTIYPKxYqooxXrGO7m/x78d0Ad3kClO7hCBLJFKTIO1duEZhiiY7sGQbtD1
56eDfBsdDs2A1iuNg0aeXXlZsunCNRXbhEn06fO7HIDJri5bybfUmpbfiQMOEki3vXRj1QeufcQj
eUxpNc147b7aLApm9thNkpWzJZgzCWsTEP08KqPGsa3uu1ZVFaJL+9y6WVb8YwdRUea9Lc7uYpN0
bjGGWWTPuu4kYAhb33MLrn7v+/vwXT4tWHXUiiA5hFd4eH9u+vLNuqf4Qki7kFuSOF6k5xo+ZebR
DVKcSEsqzeYgUxgN7P5HvKyZyDzSO29wMD3/YjYBUgsGEkneWFpWDJFgE3y/VyQUE7l4AKEYaVem
KgzAwoC0jcja0FriEGxxGoRd+S+DrX7A7H6vTNch7XTU3RGiTICARkBmMvo99pDTti9LPWftAOqy
yEDJnkSGknosgEUiWkkoDxDZyfsCBZ8nwpGpGUOKQhVPsF1A1z/fecw2elh3bYoFNtYJLUMZ43Lx
yJX1WZ01/w16+dtCjLxvF98BL9vXW0EUW3NnoluOD5HB75JY3slhB8y0NDZwEBeWSxaTY+ICpzM2
1aXbVAvl9WikZmO3QNzwNSaixxNdFQmtjFzp4hVIoua5z2AunioUWbHTiI+QUicf093PJeNjBS71
OJj9STGyO8PLQT/RCJKJ/HL1exvCPTQOLM2wTXkz/vFCFKwvNpRyQusaftr/CuRBR4jZLiR6D6vL
yBD6CwMQY4b6I114CLuJJKkyp6vO23mbXf3j2VNiEAi8eVIaNxQVNMV8L/WtR18EWIuffBu+7Ss1
aCPAeNNok79YgaLa2iejF+6JFMW6hqufcghvxPFjPGo3hU5p+ivyJJLWnabWPlZ+8cGEBBAXWnec
ed73dyuNzVuUtZYeHsKu+nh7hvzwsBuPSIEds2u5tqCGFyvgal5pSnL6AJstn2a/LLSPl2i0QwC1
5xB2bH0pYPSX/1TAaYw6n9cmZ4Z4ivby6CzSoEU3YZTjxUbdRap4+ol/vPBbHYfEmzfKo6P5PVu7
ybrPW7RKTbNCDLiny/Hex4ggoaoRdeF+9heZ4T5BHZTvgfLuPMSvLmHhAEYeiHdfmEgsHLsOUWYi
ApMwi2NOkd9/vJhnpAu9ZY2WJv6ySe5CvbOPscwUVgRd8PWLGDFjKa21c0T2ZG5CKNXKTzTvZf80
TG4CIapxiP1Jh+yU/uc/pVAJqCncl56waFmFMQRzdFq0XCgHqsn0JigK4u3LO3pmfUAuRfNGk15V
327RvJ4IQTVBioTjuSvtk5CsYGMFrztc0DYAYRH597zdw1vlnUh2CVOpQad+wFYq2xymy8LvplEo
nodot+uOY3ub2EpdCkDYDueaZjFjNVtYrqEzX5n2M8c6Yw0LRM+FxC5SdvLWzgmiWxWB66aujrdg
jvarViDtdhWXYSeFlyGAHUBMEdguAqaoFgaMTtvaZFbmuHycyHl6SM5QmAqjV73Ots4UiBV0SuTn
mhWdgHd1W9g/JHgPXVUrNyc6jWgxKHv+Nv0CQ0PkGIZMV6BnmMiWqDEaZdv71SR9ck3iDm1E8w8e
4hjumkYotet4TARW72YovYc2i+GM6QWscZ9uzddjlx1sL5FRWg7I6/mY8/s3LcO6xkXpHpdX5Z69
xpnuAyILjAErWwOBkG6BSPhCs4oVUEZQCs96luoFUBYoMgq9HNMYMASpgIjVbTOsSFWT5BeNZe+p
j/Bk3w/hf03YY62fi5oRPerErMdwPNNB8goVMmw7q0/zh1ReYVkYcqvdsLWZiuLc8p3R3bAHumQ/
ANeOzuaAsPrYWV6eyMDfcLzpSsY0oDV1raO73L2D1pIeKLv50fXIsnPrBNCZUCFAbGysmL3tRBFQ
5rh+fsQdI3E4qz6c+rfsrt3xeNTnQ+8v/4vAQgBCMbOtUTiT9cPjwgzxRbfMVkIbRTHCING+cVGm
pCYwyglHNFet821nuR6Ac+CiCn60GBcDYNIin5NQi6YMxcWb4C3r2FNKu7cR+BCrcLBgjTnn+Ycr
ca9okR2NcHBovTI5GpYY4z5wBg29y1RxUOF/7flG38OP4vbN8N9uPcuMWyhmWxc3ZgQhvCiz8vne
daxiFkZIKZ4d1ROewu66+7uiEAhhuA1Ui233u6DzUnMN5UxIsyLwfRMrCVikopTALb+JAeUykCUQ
8bCVhSdIZTn4CKKADABhIpLELBffmwl5XtJNRGjJJVbaSV+aGOyd65HrSyiSP2IQI97L7NodyP6D
+vW6/qny7tmDQYFQIhqjwqxifbrmernJ6qhZv2gPGuAmg64uufKi4IUX4ncMNiZI4lilS2oNtC3Q
iaC9WvbeGYlfE//PgtOihrcOaZ+K0kbXAycPOX3jjUQC0FBRha4ZosfB7Sgurq0yjxklptv5/5dS
nxf1uECgaQGIy/sWDzSERp9TSevd9xxEd3lc3hRnqa4tlo6Yoh6wcy4pSVBqQuPSI8MhXyhqeQVg
mg/6qY3tK+PoAJejW2eYOUBLvyIZqOvgVBm+XzNIAy1eLH8HSUwMLwUaY1gyFFVCT8XtUvNgQC5g
825WJiCw7aayacA39CLzp7dpfs7lgoEh1uNKYUxkphqnescEjfuQAyvYA10WbzT/ke3yIxZFUn2m
2DPS2Zp+C4qc7uGEAXi+ZH1VAcMHMFjYxtw67rBpwNnkJgJfZESlgH7CYMzqBepPLB1ETFU2C50z
2xmijxzCWbbQuwZBCKmkZytog9FFF6wHgv8XGshOZ14pRaoBAoF50/awubgBM1w/txhVzB2bDehc
ZVRsFx2zFgv6dm2vHlCiaGxTht/mtA0598UNTFl01i6u5QVLI50Wv8HL7Srr1i3xyU2LDlpfgRCk
bUO+im1Rb/JeUi/xTxf+4333er1bz7GfozBF35f/QYrxx6fXJrU/405QmmH/owcLNjacUQWNcCAL
ho7t2xlp+fBvNk6Zp8ps+XnpN1BqFlUGOSRqcufDgBl1Rs8zLRjBSsBD32YsgUN1U0fYZm44KqKp
wQqn8ESLXwiwCaP21aXslCO8AQrPaghZ9o1APLuVkH5aubWmgJsZ8IZegrT0RN9SOiRQeVcTsua3
/RJdfuOWhqkaWIUkmEvR71a6hqsIQo0wKuGXyjjZ6h8qmkKbpr0pNCI00RgxZPGfO5AiTS76fFMk
xEKoLUOPKR6OzTwnfP2p8VMBWDVCTcR6bgyD0qSRLERiwkK8A6i3LjcRhMokZCm1wcAh4iW8yFQ0
otVVxqQjClDhbnJPtLOLa6Mf5Of1XvLbgHjgefKWkxH0g2lo0cYrI/NFKipzkfGzoAPmNEkiv561
uF4po3oFo0CPI5OhGNUCuLm6qLg8M8NglPUQIRBsUANU2w3JFEK2++tT6Bzape3FgBmSXCsVateN
HbK2ZO85iJxVZCBEHs8ly/oTT2DjT3wv1R1LNJiq4mRM8dh56mQMEymJjdXGKKsN2qeZb+0jFhZE
d8fmKlDbjWABUOVPncjRcRU1HoTbJEqHJEauT6EWH/I7PvsSnqpikhmw8qDS3sPd+CMjAB+xGGeO
XvEBMsnfHwouaMrqBIV6qHj+QsBcZLM1T9qX1/uQd8fkejDGTHJSh1KMYu8Yjcko6wq+I6J1V/mx
toX4oQ/DL1TFSGxvVUxJ9+7HRvABJjtcYtuazb69M319fulFNt6369sRu04zY0KXKV0HGH6KVoQ8
UUXCX6Qc/136C/MQQCeXoLJH9DfTHbkMFJw//NHrz43xOyLamduIZmoxN7nXSoeVppvzwN3qvxfQ
Ds7A5TFa5eaZCDM4fHDTkwQqL0OTb7VPYqZ4QZ2fjjZnRVoUuB+yIBxqinYrKN9IloP/fIHKJJ95
VNBeWSNOPRyaFia8cCJmIQnK+IifRSmll36fX7WPkV+YF2g7Shd+Bq3xFApC8AUoJrJuuraSxU6Z
azJVU0tvj/R8oKjLQ6HsQxNkbj5Vl6iFv5tyBLMmpL35e2lxUjCXmdNNs3PWWxZuZtjK6078RF8U
+OJuhzjOia+hALsYSSMFGe257hXDk6aAZIHgpxs+mzTpF2CTnnhu9+B8uV/vtGtgVsRq+6epzxj6
wKRh8K+H93waBL5Y8NCc4RLJJ/JcVBv/41lBwFdxchCtzEAS9+rvQOGzFe4/phq1gpvVlmFSMczp
nLxejLHPWrMU/1L22y8AmdHjI1r0T3RCw98mb4Cy9c4IyLMXn04evgTW++0h25QK2+pLB0h/6d84
bWuVpOKRJnJjB10yPwrTOn9Uf7an1xO7DUCYu1jFZD5P3k89pefhljP+mkZWvxAFPlzYOrR5BOPT
TgTrMBQopu3jqUjepZuGx2QD3BtonGL1kxZVax14fj33CWAyeP17Swtt8s0xZtcwErq+D+YhbC6S
TC8LpwokA9agfB542fimY3o0fY2w59AVL1wzEbhrD9fMnVw1XMFbxOlB9aG3GyvaKSh4KdISdqAw
FYBaN9GVt6XflBjo+tMsqeXutPL5l7KaaZLtX1qtnlc0Fh2tIwJjaVPiguOBXsRbUmlFi3WQvg50
W8XjzFJH1aGz7cVp6wz185aIEYfT6Q7J9zuwYnJZSq0P7ibSfJCR2IPK6Y/I0gInzhwrfKPTZZqa
g2UvIPy20XnDe3uP6nT0mug7znmF52gKpQfCNNnibD2ZsH2QigHeyKQEws0g0OFYXU7h4+yhLE41
yBHNQzDkK2yA5Z5Cl8NHvU8M72CuFS7IB64egZvmLswSxRRUh2r2YOQbJMNu1gwi236TaHgZTT/U
xbG1+7KNbWOyG2WVgIfFrU77B/+1C33zNTKkz7Bynfmm1jiMtukM+cgnUmRdjs4rwTDps6V1xEBD
O30L7FZmCh7rwLoAMd07d9jqBaizTBntMSb+OFnFu9q9NR1sIkT+fgd+0RzD6AqGsvx30FhiQIQT
Lsa45KyG0p7Zu1ZkeizuXfh/eTmH1NkW3NR00/xl5AB2hzzSSnMWG6qyKmOmWfGX9OcROuyg/DdU
dQImiV4wAjax/YubAB0wL9Exo3z7+R/WS5V7oAhtt+242NXKJ3qddY+kM+QTDK79JbaXALhnDALR
oX4g/t/Ix/7MTnoa0kErCMcmAnyc0xkro2AKokCmHtP30GaorQJttXdbvZONiRtLRM3YL39cLg1X
3dmUuQjTctxsZyF+11cuFfwPxpiBFfNi2YVZKQ5a7mAxwGDx/uMqTMcJj4DHFjLNqowuu55k3JDX
x3zkV/nRtPaFYHdYoE31cn8C1uuLWRBH6DrHUaJ5CLpQTR5ay81C47cs7p1XrIIoW8aCuZBYEPFh
O2HtabWO1oC0gu4sMM/+f59Bagv2n1mdVL2n1XEBepnKmr1qMfKdvna4nZ+G3AUKOAv0WWtFSXIG
6JaQOKZ0MXMOD6Rtib1SNmITibzl/CNad811zrh4v6SKS7XnN78fxd+xpC/vwWYMXR/4vHL6DeYs
SnE+OhPty+38ecvFO8cYwtT2YdB0H2cFgm6wzFC5ex1x6RDWpQ+scH4Zm0rn4KcKhleo/sYYnBFA
f63JBX59OB5pK7dThBR4R8937F9FvGH9Bz15M91dS1IG0td/brA1T2gL8FTT7ZKsY3b/5ZdwNda2
TAqHSGkNTHD0BciExncdrKqzTI42yQHZYIHIZFYrajuY3tRacT+V91BR2vG6SvHUw+izKaxUvjUX
ABdshJ9f2TdcfPvFRUtWqDk7Yny2AVhWhyevn0ZO5WRzEKZH3SFMuPvw5MKwXkeYEtOUJPXsb6an
LTxoC78rX14CX0Tbqli0ifSdC5y6Mw2cXOId4A1BjzefKbz9dcyAydy/bLDtlCOTlqj9zrv87uec
rGGTmdhDlhwn5uwELKkiMI5iuxXhrlPwppEkqI0i0N3123r6wbsjSRqddsDLjlkaNrRKmWycqR/F
/bqm6GMWSzPlZvTWlZFMGdgnje31NP7/pZ/reYcZvNe0gY7wCd87HeevaPLjAXVGHH93wmQGBN0E
mpzB7Z3Ak7/xr3bWDFCr07q2ZZiZ0zvmxHDuPRO+ZUtKqwhDF9335jfcF6jmyKjUeSvHbiIm7yp8
uraOzdAVGBCc+oAphbe0D4F5LRm9foWIC3luxEgkLBU6ZtiYiI0dOGGtagGtQ5qVyLNQy8VvvP+C
Jq1o9LZoRaYgcnABqdWBCwaG2FRsmWaKKzwnbiLltwHGombLIZdXe5aH0oqOBGGY7R5xZgwWQFQc
ghqY90q4acjMuZPFFvcBU69S0CIbRendN6ahHlkdr1nyXuV+Qt77mz3rZH4IacOnCV5c1wnHfrkA
+GX3QeF5Y9gpPTIBK7AunZTrWUfF2QcbYzQLGv7PVDeOiKXeqjBRrW7hj0ceFocKCbuixz67tZc9
ztzmq01xip4M2qBW2d+2I9j1itulM0ydfjsCyLXck1IPTkImSnLbKLaKEDUZDKFDQ9LAbqLI+UzK
x4vrjQBEk1/9HGZG5JIMsi1g2KSEWRRFuiZ9aKHDVfVmGXN3keIwYUInDxJhW5AsMEQFMrZH1zez
nPUng3fZB5GAx3m64Qwrozvf4pOxMBHtqHSeXektCVTUpPJygBoUfO5/mwlK7JVw04UqaUEruWV4
+fIOhRpBZcAMzoJ19xHZrxZSdET2XgHrfjL/A0t/lmGUZVIZm4fNiAqnnVnFa6fvFPkLSMEOVBkp
RMJfW6tGFYVqJLtMEDDihST/ghNW0g9ZEX+YvoWZ2veQajbp784msdKGpEb5LrHu9LQsGaZXqRpM
ckYp0IemelPcG2R/exQoBXDLSOfU5YMCJBjlwk0KHw91/XNXEexyuS+JPQ+b5w6+yOyiLcMoLbE1
GUXuzegEsFo60zidK36Ap4Z9S527geGwXNKNsvJ+1jrFqDWeyNYtkUTJBudMIzydVYey/Y9l0aeJ
3rJdfZDNJc/lZ2aeIlWSgLAiBEl0+WLNuEHAA5gqSg1zv3i9LuQM+4ZLOUGNM3qhOSybpDfKUp90
YKStexaEIcwJD0Pdobz3oRwJoQEyAlc1UrxqcKpSjqPXHbhg5bDB7skcrLmgVJy6Jf5yXobkRR98
UuYMAWbWNalOnx8JFWdoUCfFvIpAg+69diSLoj7IXhHH2KsRycVxAKOIN4YH3UciQdwZGs4qsz9i
5JOiPZ1N2f3OBOd7zVU1K8pmWLBkqSlejtt3GbP5ntSG0wI0jWfy4ZL6PO2R9qDX0bCHQ2kWF1Ir
BAuQhyZlIwCgOFlLAuPNdQWt+3VBAF+RpMlboWItJhicm3VAm57FBPcTEeU1PP5ppCzg6Or49Miv
Hf2bmR57K3Iakj4NQlOACGgcEwCSLIRXuqjxazrds8nciyw7fB/YSsrGOTjEaxk3yAnGZMRRgeJr
KEsyiQAkbOPyFi/pExqWIwTasWjyeb7spY34qfocrvf1J7yMqikKU+wXapTr6EUETQ7NTfhiSHXI
y6FysxjgN087+WYBaG9EdyBq14Zxyokk0gKVhEiqGS2roaICr2m/EwI+N5FtsKXDDm2rCzTauIu/
M9B7l7uZhNjzOhXP3qdwR1amvmbn/CZPD26azBj8HJNvU8ugFjjXsj1RNvrFvIOs0souERqmBBKr
KcLgl55xfJgzlI6rsRMHg9h84yPyvmYhjIiTOl8nxDgAKmW3W69KLG5kkCnB0SFNIQzVFYjgScMn
d1pHzHCjDHdjzdVmBNwMSoll7maUOg7NMi1wMebUFhpXq+Kmsv0ej43S+JhU1WKy3pHorQy1cnRa
hb4mo5OEao694y9w9kZ45GWp72Pk+HydIA2HttmociVdMyBUiQ1iqnKAMX3yaxZsfxwpss2xvul+
r+djlvxOoRwLrajhIhiGr586zwkmsSO9if5cZbMhHJFrnWgVGu/yKF/ndrIAEMnJElgyJqOtZTcd
pmbt6rSi7hIw2VfVX2eKBMrfln7JfAsEtgP6pRHS2+NwDkqdFCMQfC8U3Brx668QHsGZ2tc9r/jN
oE1LgqJ0aHLye2ZAOsZTqzK7TA5YrOzRMJaXShbHZGHvTmYI8267s3u2QgMwZA9lx81dpZDug+HS
w6m0Haa8/CnEO2/NlkOcY4uRRohJ9LkRHVplnet3TuZht2GBK853novG6ix1zXsmvsMPJdAmJCGp
uNqlRtfhH6c3T1bR0Gij56J4UM5JHURABqnJjISOsnjlrNcZl2c2MBVSITZh7c+WrKARTfcJc5TL
6xX7sa76c1T2Se528wE8ju5VoZwCFcqrFLv4f6mTjz22c1ddE8kdq0gmmiWVnQV0z9ML2FWeLNy2
8IwBXq6GtrwbvcrAaXZfab7HQt3I/d1Yop2EbbA4I8lsGG4W4DAV5W3OL7iNNkplzRii48zdmZGW
tU7OAQT09tlE1RHnUKX07nl7bI1cRXO9bb477HNO44Iw9ftOU51ANg5PCz6y2Rv2GWuFz8pRSBi+
VMKRp0hGbQPHya9PnnJkSRYzF+gK7vGMz2wFYgSxDMwqncbGeEZY2XUQ7DGoBpbRi14XpIb4j3jE
bZl2+hgQiVroMgJxlHRrMbZA+4BNalJRPBsYyGWXZUAKicjfLsBSdzeeQY5u6eT62wRik0ySMc8c
w88mDpGrrZmAiwAz221H95qm4oB1A3ztTWRlwDKOKoZ7prj6EpennIR/I19xqeEIyO+oUlrU7V7F
MH4jZnHAZXXH88anHSynhtOmwzK6cySFTIAVSURTtrD3OLT26pHHtt61/80tMdKAJFsUnE8pCq2E
Gb4V6RVsw7dA6/mdS3zosv5c6IaerTL2O0x3BxhFavYsBiEgSifcAcxvp+bBH+TpETZ4KpSByr7/
zOmavkXqGkbwMvr/R7P894wyM3tHSKZgcMfvglErIttgxHcPwau916/wwEHwuobA7dIeeqUgp43t
9EMLPfn6t38CPYT4dEIOcZ4DTofCEj49NL6/GjLXqWSUnOkDmxgxGKcaA+H6wp0W9LNQBc03vS0d
Uk05sfnErvsNkf69GiCpUHiL1z58dmSzzE+WMSWV6/wIcBXluLKj4X8FWzPwvK8n7vEjn1+fZ71r
7tS609uFUm9KKZE3JkFd2c7JTeq19Twq+cv7tXpUg5yJjkpN1U6azJNnDmvj2xpQurdFjk2uNb14
tuxuzpef005fw100lponzhXZtlPgyt8NtIaOnVktVyPy2ytYmKFnXMVhVPsz5sPDw8p59TnOu/BH
J0tcH9STgvliskeLjmN26gOqektP8jde1tlDLysY/2sQV4f2LsVvZk0D5kQs0O5okRdJxI8NHT4l
EqQOGNEguRo9U5GjmSQVy8JXvgCdaosE6WNclqjYpsZDJijEyRGW5Ppcmw1q9fYqd7tFUAUhLBt3
4ysbd8CK8KBO4e0WMTToqKWlmzUvCsYAeO8ak9huCw3zP/y6R3X9BdVzx/oznTzuZomb2DCqtkdV
t88nDJJHqyhSPreAEUqUeSptAFw6kWr3DFTU+a/tK3Af+TXgTKtUS9v3SYxbjyWgfPN7UH6DKzB6
naeT9/afwyjRWqyBNuV2B0+Yebb9FCh8dbLO9Zvrt4jUdERBud6eF2w8i1vDGaCXTxUW6iQKpYf0
8uxwy6cE8OiAVfT3O8B/MsIPx2soyS0hRdN2tS2gDviZmWK40P9N8uFx8H+1iks4ugPiGb9YScTM
Id7dLMu4tZamq3B1bcraiDX/0BB13Fp/feWbJFVqctK0kCHe9v4KOIiM7F4EcZXdZDsoIYE9q2/0
qy2gfyrBWFd04zNpu8AF28bUfC4VpsffhhILOYLj8QDxhDEY9ZgFc4Ce2N+aMSK6UEYJ+ieCn/KN
vFR56N1kOALfKuXF3oUyfMOpJO4cVHA+5+UDtJ9HI9GvCXRwFPSLXi3cV1QEjW8cdx/UErvCe8zo
bh5I8q+oc2O4dmzOzwl0WCg8qvozfyN1l4QnJ5AA/ghWVUqnwjIP8hSEd+IYVZ2JOqMH/edPSDoY
hwlJqPQ6dCW7IqrWkja6LAKZh94wWjWEKBFND3lYlNmqIbZL/e523Kxu1c/J4Sd06NVxnjNmGPtJ
c6sprMbUrUZ0LR6fNz3Nn6RRaS2uNh+A6n6CBn4mlQOH0I6rKmkjq5whxAqrr6QZgLiiMyTLhZjD
yr6WPbDPw+ARxmooqBpYZQsu+3d164qW//LrcC8Vxnqyk+F0giK7VMP6WlfKPAIoFMhOrBhw1vYd
WUxLr5ZIcdxyn4336O0SHmM8wUHPauHAkm7MNc+UoE5U3kcQb0lADomPAB2gLX3eWi7E3MaGsgv8
qTc7RbGhRraWjfX7kJEO0k5WZZ8f0YMDZkwaClX+AVOjEEGXBWaezxsyuqMsQpY/Jk9iUO/tB6SH
X1Noj2G1VL/GRyzUHhk6h5KALq0clkBrYN5n4ShVnn3OrLgkx1RjstCVw1fLPp0ThxvWfx1BHZTS
k83EQ8hIm5xsjufDYSQiOL1y1hTRj5MwmBcUJtoFB6rsf5qANkQssyh04ygowyq5eUFjZoibMj/m
hO7DMtPEP6p0ya9+WeiTGfh+DYfMYWa+G15GrBSk47gyRKiUwU353NVyCf3AjF34t/ii4k5WzsKm
IqU3JfsVE7bQa4IlwoM1hg8iieTd/4VNOUqx+oUTg2HC6TdWOyNDiHgVUg763uVnwYtbb/fvUEFp
GefPk4P3dlg9nzH8s7d5M2yMsBFzpczyLu0afsAP2cY2oEwpGC5UYKaliOKNEN1XlT0uDXpQNFar
LSyNrl6Ismsd6JTimHvBHodeDHCQYfD++i2IOy9lpaojGARzn5xUX4b5kMbeee96rHQz8W98/7Dt
hSlxrDmDFfnajvCVSRWXomw14td0hA90EbLthpw4cgQIQZ6IMQcqz5xwvEOJWlKgfdm7oayB/7pD
9H5piQJ3V80YNaOODkPGdSoQ1Y77gjydwODGtAfpLPk9OwGTA1FYbJ166oH0nCtLD2PQWf2Cva9z
mMcUfCVWi9V+NdbkY5G9mHJyvr/wpi6e7nSEsEkAZGbu+nnrLp+GSDBRyKvFphRdYAiKKttfRzd4
oWmtLsy+5KFuQVuOvEHaDg3ZiceQ95GOsuLFpRFes8jRaQYZTOB/MNyb354yz7r2jiSt8n0XN1An
OPZUvrDDQMwwSslO9axFqgSR0eC9uBrWxSV/IfVVPOehWTvvAmR5ktygtOG4Z22qwZnxTX38NZky
W25m4o3ZlVEE2plVlHhmHKfiASN+aaPeEZV/nUDg1rD1FEwwocDUAMkyue8xOUAmUX8tzOUV0KOC
NxOQT3PY/Yfqp+ir/pbWC4DaM6XhY5F42IbIfqWgvEN/snWPZlXGijbJmozVXcWnzLefY7l4PMTM
SAk4qCe6SG1x1W4gCv6Ml2Dtp+CICCGGLlZlWdZtXtsIt61acR54noWNSRO6DXy4Ets4P0mQAWQc
rXxcYX/5aMBYaJZU1lrQimC0LGn+2IyQrNOQkoc/2uI1wK3IMQkR6TILJvsuHE6lfW+3RGQo2nRk
v3KMRAdrXrG9GMb9njLKYfIgxWJC/MiTevYOu/gmPrWI0rV+UqHPRRV21s13AqKdd0Ub86d2U9zV
I0C0ylnDQc4P6VmJBrFAyo8IL5aN+ZCdootwcKI5vMEWRi0v1z/rjXUoziJg7qsbptqUCwluddZN
mhAUIRlHJZ5XtGlmuFxN/NXFiyxWGyrU3vQjkiKnLeh1CNq3JnFPkqwUVA+1+p8803O4//gzrGsH
ZBZ9nfmAQzuEa+kySUsqAhZpypV9j0+jVkwSgyhDVi3oecMJPv9/NndKJp9ubLIELJVKF7BC7s0F
5zitjpzyQpSmBKdaooE+7ihyf/BoY9KLizgdAX51mkcWtbnXIUU7EAqAc9u8if2WCNcxgw6ewFL1
NCefIvDBm26KJJ3HqXZbQbJsCl0SylAdKp0oB3jQ7p7VGonkdEQJiBfpmnycXZ0htixUAUDI1jHM
qS/y1S4mFS0Z1CUjOqL4Vl4a7T9+IhHn5azgzKpRd4GLsFlqy92Xig1SEqbfm/Lbv15s2Oo95CSo
lsWyF3oHxpXWdR0cRH19+23Px+NEdU8+u/HGVowDmxX3GRflWeD22ip1u1JIl8xMEYKpg0HU3gif
Ebkeqp6CyAE/rg/nTv5UlbfPKmO54h+9/98jWD7HPBqeyOdPptR7JQ/dEQYZs3hgKUyw1HYa0Sig
GveAG9YIX1mo3PUVlTRbcdReeZ8k3q6a0aChtyCZ5Oo3DgU77HU5ki4Rqgri1bVif7yh3YSRnkvl
NwOwMpOU4Jj2Sy3TjXajhwgM6pv3WqY117QDYK+Ja0/GzUyt6zVknkxhAT60U88UI+GZju1uQ+IC
VD4Pgj19+Lqph4/etnlZe0s/aRiLjTy+4fkX7zsAQpRWuaZ+CJf1dUfE73sEEbPea0eFNz4/U6Cq
BLZgbcOWHYaMcEveeb7T72yeZX5LXGBsw+2Snoj9aiPUnV+KBKldubSEhzfDbKzR/SYi0LiWodk8
LS3CCyOwwSp1tXWHqzvNNZ5I/M8dlbhT4FkfXqZyG4iWJOSAMN3TPF3agni7HzX1fqfIdYW6RctC
rsn6doKnNp9pJuNibQ/q9RT+wmCLLh0bYiZ9BSKOnQtT68pEii/LrBDIZVxUuLqu0gARbtj1Jz3x
e4QxRZQz+GUpaXBvxjpKmbEIN3NB/DKCP/dC7N6QWggKE30Mxh5E1GHjssBoOgHidg9IUyk7jQIM
oa2ado5I2VcorkU5TynjUSZxEtI6buZklyb8g34I7sKhzH6XaggMpLJeY1eZttjXwNcwbnalX1Du
CDdt3uUX6X/1wCbi4WGnZ9qOXKccWSiOXTMvQxAClzy8YCPgBkLMZOO+0PqAdpR1DVH6VDhtblvj
jemjbmuV8pB1i+GEp/iIEiQbWs2e9sfoZ1WNobYLD9+/j5RHS8Mdjo+XEdwRKAfZg7Z2n1NGJGS/
7C2dTO7W/DAONtzEwmj8U7XkmAuungv2FHXZBIIEw9cYmCAvDhTVKuBtyD+/jDr65C2+psMF154i
XERCh6egqB+gVVEYLt5DT2fAB3JFuoH8NMGb3E40Xk9cIBTnNIpp88mqjn7iQW5H1qdOcm0UPRYo
TaIT0GOEKzJKWqhGoqICNehASIISeXE7smt5VHGIV0Kzb/t4YDIp+k7eKn4jFnEfvk+nD29nmCFo
hyV9K0f5y5XsvzhRxe/WYPxrQ/CirY5V+fbR+MGSn5O2PrdRokNvbsvjEzeE3hJHz14u25yc9GzF
0R4uHa4rQR35K4XDgCrgag0tw6Sy7LIe4PN/ki1uS3zcQKPCb951KvwzR7zKkM3a30zOewDaO2rg
6CutxO3Eh7iohvzNCEWUEnL5AdS0QexKjiiuZcSBclK5F8HQX+/w+ubNX2UaB6l1NSfRUFtqSCNg
+dlBUMyaxkDH5qYM4b2mwXUUnO3S9r1PWOPuCX4QXTvnSnNFFWVVCZQuNZlA9f7NwBZLrPT8cx2E
nSR5v3A5I2+ozwEvLFWTHn74Rr673mg80xPQYv7nOEkN/QUcXlwzT2nrGbYfaPAPMFp4NyKOVkds
PjnqJjx/oa6DiT5FI3G4Q7GedyDPpEzoklbWGBFLm1PJaeaGsoSgav+hGMqmVw3jGoRcJv758Q2a
+KxM2dLrifMPig95vAFnn7boim0z70m+rEutMa38SCf2WHM22g301rkAa7nR1sIPy+4NZBxO/Hm7
40Q1L58DDPMPrxa6Ovmrn7ZxymHDmpMtTJlfWHkOsPT2vUEeEGbRRm2Rx+t1a7Kw/dw05n889wDo
6LdLuiP04YIAm3dXprt40ksSJQhrttmdEeu1O69vvqRUYkbivja2DLEdM0usRyWhtNJHU/3izdNB
4MULgR7RBkf4OCqhNlKIaQaW83X3V0SX+aFtdjR9VM7iKtJKHL+mfUOwjzUfmeOUQtp55TFFjh7o
9mirp/X8soKXB4lwmXwKk1CdxLYQ6cSZJJbXzAbbZVlEtkXwvZwxg/fCWAPPLJhhpIHbpDNqWSx0
QEvUlp7Xw+95TEielqVq6NRav0w4uEiudNxvbwTgaHmPnpsGJgmQAonOf1wijAdeDZ9mibE2xFA7
e/NBY8OjMEgKkvesE/wFpWq4kxElb1lf25AL+yZUA95yFTKz61NtrV3arlPO2HBjk2PBAkOlMu2m
xSF9hS4Xhz5ZzIunOGh6WkwoEem7keTS9MHJWcnkss+1Y9bqmUTSYjxWo04iyeko1EG5wLyilCe8
4OFhliufIxVuRyNo/1Fj99QGsSfzW/ZRdV05y5Q45cAuxmCbiQRMDWxZgkCq5gvTflQDQPL+0HcP
u082KbS1GbWu+IyOOdJYc4GHNl+lvyVPyA1Zc5ddPQkrhSPmitVolHopzMvnBE83L3tML2EZJj+i
Pi/f0mbzgNfhaXF5VJBNEhyV5tv5fgJxP7u7+AeBekz6MwAZCMR31CiT4EJucSB13Ma55QcUD/OZ
jwIHMaiTvsKfmP8Li0+g3ncwXUVXUe8k8gjf2cb8r58Stmk93e45uXetxh3yDIeajqu1T4prySDY
MyeIIniZtazidFSQhVLuH2I+wlLHWL06zAg6Cf5v9DHAYmX1JdTo3eT04j5K2fPQRGWlJA1WGOYg
zE3AUdFJ9/ffriGwL2RPCA/0Ppp5DCbrKXQGdruq2kbNdK0yT6dYwgYweswGPGljASrQ1EP0WvXK
DndqPLZKi867wbQ7JlvpqiCniYx6F8dMgsk/ATTRSx3WMfIzno1VvBkcwaKxJjwl2pj5LIRAcouZ
SsJMzEakHXpgZJF5bUT3AhDhDCwfkHi4ICGESpDzuADurrJZ85HLwHMvAppHUXezCnPhws7BvoGe
cDfZEsYuP7vCBw0YBZJpfud1/9e7XXBIBPTOYrMbsQqPp5e6fnoHTjpS9TQAeXdYv2Bs94wIaIBb
b1b67SCNnSVgAqlIv1rB5xZarI5buR7lf9xmZg6MEWnzioRzLYFN2dk2rotRU/FtFI+ffo3uVuGQ
aEHCNtrlTesHJ08j80dPE5jpFxJ3wK0P4z/eRKjvCv1R/fvP4ulBHLiOQgFo/kZ58uoCSt/UVckV
4ViaTqKhtByRpn82SwKvkeC9H2kncEJYVaBPT31TQFxWUcLFRnVeyGQVeNfSiBxIQSco4D3VBxj1
MWpwOmX81zw0VMPm3YJ/biYtoKnmuYSXfug7Xwvd7IsxT7U7zrJ3y/kQWd4o4YE/d9oI1EmWv9L/
y8FZDm8qiakpVjzbzFb86L5XEZLdrnjiC2lO9cXfB5cUuwr5TgCFrRpgF2ik6/2k3k7pfgwxZDXo
MlUaJEUMkDaB/KDjKcG1U1aLYFpPVm2T51Dis6QoSgvqjwa4tItx6ebMMjvnCVn2BzfVCES4cOgi
oiMQs6FeqgKUdo9WnwpYxHs/Jdff7vkXyoV4suMpy+Dtt+8TOZLThF6Cn/n+XaJVMoPi3mNAIY0r
wNBokXPb5MF5ELOZBaK6kWC9fPYzeedxBt4eLffJAed/vnH/RTnyUaF2oLdsJLy9Q9ATFRi+RXCT
mzKTJNvOwjjxVfuKltuxu/p07yTTwAxmBGwvo2ypIjfhxNph5BX/CEz3cH9PwNe2nHhIKWs+VW+Z
auTE+3quxFIMxHTA8lCoDQrT0uoNzAluY76TXdvzq8aM0z1ffFoTDvjkClx4FJTbMRwTfO6bvz73
Eq8OrbxeMmXbMwFpCXhTp+ExFjYsm1pJrLduqOzocynGG3XSrSxPlutUpABPleQDSWyDq5SwvUwe
g73E87S/u/AMlPj9+dm+cb8dxULnh5DbOl95tSD/bSE7E5rz0WRvNYkHz1szJ21vv1+ty/yeAW7X
l1bbFImu2hVg3tK2BAj5GeBs2fCyxDIJQzOq8qwp3LdnZNBhrLlPw47QtqbMGR8d/TgRjJ/3DWpe
omPJibcRsrhmgCzqWVbzV7pxbf7YHNvqR593jARPvZik3qAlzt7R0knWcLYjEgv601P6wpO8kEyK
S9zpiygsgqjWHX1lYjttSWtXm0ocz1t/n5APilnDnY1N82h5k3CQ9R0pIpK+exy8QWkgMUbDaHR1
vMcgCZtS4eugaWctHmPRfcByN+Tn/JGfskXYUdxgAS851iPs+kOqob1oBsoUYlpftSbbnJnhkte8
cFS96PZMyiLEYSm++AaJhZbNflWrgDV5+IzaA8qqHrKeW+gQdi/sgWZa2OkmwS+hgZPrQOXx8xqx
yyNvpUo8zkZxgb4z/jbUzHYMkwciAUu9ZuBRolc0UjjKXQ+4lq3hpYgjvlSyTXemIwTgXfWkBLLk
o0W/uF7qI6AJNuqxuict1jT4ow485yxZM2fnmeQ4/Rty32Gw+m0d2x/vfsWB6mwns6XNXAKNFcHi
dWBQqb/uFs4IdoJc7TCc7KmSoNr6C2kA0+/CpgBXhJte1vs6OOnqPJ5HntuqxctyOOlbPcPI2efj
sQtfrSNwbYXrtPZ7zlFK6Jg+YmIxMIn1b7vPupxpnKAEKpHAs0/iTaIx+eFIMdre2z8BfEGDpezf
G0zY6kwlwwl/kI5q8QpLGSezCA6tCShLtrYiW1LhT3NkFXJYXC6eXXMh77DvT13cXUMtSiqcIoB3
bo7Nj+++z21fKJwv0kcQilx7tBHDTtheBrTHLagCcH4pWQ6OI/3hX6jrefCAdUMNXsq8jQOKsOrj
bOeuuKrvSvA+tDwEK+MONTa2lheGb1yrQKRkqe/xHZhyp9Zd8l/1Qf/VsjWEcOZDgS2XcfxJHZ/7
5gdd+H4Ct58JaVZ8iHWQWBV0V4jTH//u7jUv0yS+n0sZFv73u0R3R2L7CeRsyNG4eyjmXMpZFfcr
oxWLdWySq9DokRZWpz5IijGDK/feEJItEVM3xVCiuC58WLO1ybzECkbzYTdOq0l6UmgPTB1P56+P
or6K22ZahiP4u5RcwEkOOnJ+5FY4C9Nr95U75VcQYOv9X5H1lwd2l8vhn0G3j5Pw0vhJb8UUsi2D
oflCnRh1lLfLM327W3tKZSx9ET4NNbX00385UhaSocExTlr6fA+wCp3kL5SdHM827btkM3bR5xtJ
c0M25EDaPysuHtkUP5wmQX4yHqp2fpwnohUGfeoM+mR6ILzP9eeUU09UeQdcGUI1kihUW1sgADyd
USro/YPap7S4FzJMTdwpDHICfNnAH9oIEEkGmetJurJ4M4ayv/zPEWERSPnNlS12e1gr+Rc4U5Dd
Qoi7JhDO/7t/aQoE7tbgNEzaaOrWJBEMIVdkYpUtS1MTGGbEB42eQONGXueF3rQ1wUZFAjiKaAFl
Mgzp3Ii9xXLfaTDnJavbvS82csG+HXUvbVNjsM5zMkq0PnEH/bdby1aczbY8EjfBFid1FWau+J6R
zv+j7NSwNn4dXQyEUAWg6gLu+aCvUh56hTMbmXL7cljb9fvLft52iJDUvQu9m5nodJodGUHp9g/x
eY63kQHmFtCq+eHBecmpDdVtD1eZvAzwcCbda0qIm4iQ8E3URhuPZMbFOPbUbOtANQEp6QET6ofv
nAsXlIk95blLzxN27zWJIeIShqnueBvsD8hK/wLSFX5c3IxSSkcMlbBQfbOTAYwrX+zFDv35d0fK
949VxtYWgGDVhG6tvHldI2KBsUtAcE8vI+QxWom0OL70kQtcve3EcFmXQbwYPnVJkB1m8tihWw2G
XsDK3G/a0uNuA2w8aQtfZAO1EAq/fbK1zzWmp6gUhetepN9dtU/Nde8sKJmGIuYZLCcItYeuOfia
UoRshuhbhAG60hFqdZPR1OafDgRDfOAQXA3pmysiM7ulI63ujOfFq4ns70B1c1CZfmKPIg00TJhe
URSlS+hXKLeLbD2b87d4qceI0mnxlshJJxF4aZ8r9vn3hEYKx8541QGvSEMrhAnvhCxk8IU8EQrr
r+jk62O1uBUZkxSd3N5zX8yWX+574SV3MYQLNR50czIoygOd5+V7FRMvL/+tyXmH2osz88jz8SYf
ljPkEmfrUfISGtGYHY8BGaxfo5HpTehniidaecq0hc3QD06qorAlOsuXIBk/yjLxxCDmEaOIPZCD
d6mb/1dfl18bumOHsL3ieg6Gq2v6l7aQVbGQ/1Ko8k1/pyvsGPc1UGCuR/HpdS1NaTkyG5sIjgxb
d0D6xkaO3Gn+pjSz6FM6WzeW0zg83+wV8AO0ROCqq9hkJ9lC/BgBLMahJL6r4Uyd2Kw9WT9rIB/B
KptU+KPKE3f4tdYirwTPypQ3DOMrBzt3T0PS7OEEA+wfbBywgWqtmT9HWB07pnFHPI2Titn/SaXB
R60JeUL8OrbVa28+EI23hS2o7xoNkSQsyBXsPVK13DDiC30QpYjkXjXbLYW0az7LNrn3p9RlM1Du
IDqF4bg7tHvlv/lmBntedRx4yCDtdrXuo0MThlZSPiMmtZHTeHEEhFhAFGhK20IaQFSxjvGdU5FG
UhW4wxDxTmArTWLNbe9hJqVt5dZxVRmg3735uY59m7Cvw5e99FeKzRAsynMngCy4cq2AmQzeZBNb
R0CCKy3bkk0B3WJY3Pz+Sibu3rWiyPS+hEH1pCgMRwQVfrjZQhH8CW8SywofkONGGJERA9XFkW7M
HlSeqIT02DEyXaSBher7oFfgl1OZp0nWJ4IaZaHqpijVtkTdnkS2vr6O5tQIwQuBNZhs3VeLcevv
uYFA3iNMGwLSICkoU24EO7gAgJxF5qmIUQY6w8OcwLVeLfojyUDfh+gZy+GY7zLI0heg/oxEMKWm
yGwthfy+YM68vwdUrVnsPosPFOs0qhCF2ReaAmlzDxbdRUWFZXy/V3SgeEtRaOQjgUq/roCFJgVC
pnotCT50LOHWlDEij2snSCqNoTflKRFPYoHt1++LhOXJ3anMzecsi8qh13D8xTbZsnfb+B5fznih
k688ZiFs5A4IDToKLHD9eoaP6dEYuP5gJDP38IZrNm/DRfidc+Ux/e9r62EmWehA6b3NTrK0PAR2
w/RyHjbrxMcmOpqTXufiqEzzkdAZTrPqE4aDl4k7MdlkCjM0FWB37HdYMm+OF5W4Ui6xCtg7J4Ek
5Dxg06Cu9VI64RjPMhvxvsdjYFuulL1euDOB3FoWlDvIDTgJkx8s7ev/GT55UFJXWy98zCpjkqis
2aYxqlUoVKEIHMot5ogVcLMIgdwDtpjP+VgFvBVIk53panIaYkEkT8UYfd1oLi/RcnsFBi0oCvXo
9NLGiRGY9hix7jcSowA+VUPDpW7qBrPyaxiROGR9U+fd98aPUW57bUi60b46nt+HaP+GNyZ+7t6t
6moWyddtm9hwdxdz8MS4DR2I/Yu84p5uRPtBvbQmqDBaUXWfvE4WJvjPsbOzDmds/fem7divctCY
caI2gkJ2GRXeIOROKgnC10zXl/g4h0Re4RgtRV6Zh70LPsD0wHthWgZ+KcSlxYYOnd4Tb7iLLWkv
nGNsTK7+CqeZv6RQ5WtQeq4UhIZcDx8IsI3AXpOR3VDqbwbb2gI5N3KU/Yaa2AA27KMMwf536IEO
YV1ehTFiyAk7s6zOn1AqHxAlVIiJ/UrtLS9uScSz/uamPgVSWnZ2zB79Iilfb6l8GaCuBXMHL7LW
RqQfO7rTwtoIkY+87OjBto4NW1MOayVw+Ntv0E3wprFD/gfl1pf1UUXRS8KKe92tuqIxmnkfd1RR
90Kn3D87NatVcf5BZl8iaoeGLoRRtS0bcb3jWiI/kixlGT1BJkf1VCTTjoOvAEZElLnUx9gWp8HV
iRmKcPTqqkUskFdwRmg6SApbhICmjJW4/LCjVIQeupe2MfWvN03V/7Y71ZHGYAg/7/5vjYDRbc5/
fArByyHwB2w+7qodE+mo8hHHzEaMoGhQeaGncpPuAp1jd4uwMpr6fPP30PGQAt8AEqBHaa9s22WL
9Xad2GcBP4I2hj4LbCqnLgroinVolPjgA3DUtlbHcG3k19EvezED2JX/pUhJXISG6D7tCij0xulv
jHYG+WDd+owmaWMwf8hZiaYuXO/3qnMffRnW+awZ3PAO56FyzjZ9CK6HZNeGYfEf6AR1ql0m/UNt
cnSGnVMxIrRsfYzSn7e1JeFgHRatJ0TdmBdind4MxyK6SAQbHIz95q6vSlGPu6NJi420QYOWINpQ
E9SxuECF6OZJT20DC8lvSumwEbI3XTDUK2/OL3av9GxOVoZ5MCar6G9vrAJJY8myQhWgdznb5lud
QG41Kaj2bc5iEtqq3cZAIYm6WuKwAWyxF0z8wsGHcGF2TrXpJi8VEqET+Tv0w8HEcRldMV/QSLvk
KDTdn2Mq09OTgMEu9vxzH6H+kTnoc02t2P+Z+QrkN3Xw1/I2Ht8L+UBlGcQ6ZCWnQJm+WxT+5/P/
KFZFJlVbgDQs5Imo3d9zt+ah4HTtXeKFTYncg11jAwHigw6+cCjuKTFv6WgnVvop1R2Olv3Dsb6W
4fR/0Q9rnNkT/OphnHpjNT5+8n9GRhJqzj7FkeA0M7yslb/ZajGT46PyCehMovhnyPibeRF8tA6X
A9MvP30mWPvq7hXaaMRjiVlvZE5bkUcR6fG+ZmC19FWS07cW1lZHjNT0FyWgGI2itkJPuBk0n0sF
iBwhe3crpmu8KTk8iSNqZOlbmtp4MYHJSGqIUp3aZXj3raP/FtZ0hoO4+NFagjK+qfcnunApmKfG
rurgt4TReWqtos+6ZxbguY0sYydcu026pvJsouvW4+lcw5mOlQE/LammkF1othrtsY7mWkWpSQTK
nFRqrzdgwwsa0ukYJjIVk+xoppnV9l6KcriB/mHHw71vrmXqNBw55ujPrOxiKaCZGNcx7Bmr/EOz
QRztwCdzCOdIsBznHK+W7Iaj5wnZQOjfbedETGD0Qmtt4vso34MMtSgJluOIYtNTTX6nIu+/EPOD
h51XkXSoFzcXvTYMYUiOWIKrMC+0mF/z/ZoYM/TlO3d0fnF1oNf+YwDAO92/ivIQCBwTIF5roKW+
5al6Rd65Vd9h1xu+Fui5J2kLYZm58buk6R46Fjep3+s7uuzwygLke7TAgLl56dPXOldpsWcF4rDO
1kRXiN9HJ+0A8goitxwlXheZjuICcakg3pdxJtVuUXXhutKVvE1bKerJwfTqs5wfsd7qmG3ckUZO
3BSSf/B9kowSnDVlpUlek9BUZ+ADPQKTerARoU5y+x8cgVlDXConCnIuwVkjfUTQZCMDXQFgPv2R
eE51rrXpTRd1KODzMKsOFd1xlZSm5oQbRnIBRf80yhR94Ah2gqxOvCPahMUd8nllAcoUoKDsIltk
bEDYwVCm/el36qErl1s00KBcMj6n6RXMGw3huRqknkxSszzGX6xF7LAGhHhYeagyCEhwsRlPRIH+
AwztB00xUUrYFnKFzBoqpTb4N7O+px0wtOaxS/wheUfVKHw6A5yj+eDMsGdvOyz9WOG0mfI/XNHB
K/riADfBCfkUgkATwd8uzhuZVkwwEsi2y8G/Pg9ZuXTsAAAS2aaA+PXXfGgL49Exn3FHIFG8Tb85
FjG2Xg1sD1Tf0jDVVfU33DglNOIAB43b6UjRFDqCp5UVrCZlGwhZdpYo3K8IkQwTSAMkry6JCOX6
C/Cm1AcNvLTc1V0809738PSkAwrg42WqjOPIM+v3Fs3e1nDrgrkpNcYyw3BjPdO0RukznFXQdoDU
q9cVV5yll336MBXIOGVdoFl/sTo1CYO38QoxfcVfkaUr5SdDN6ZAxOW58/0o9DpFGIEmIdD5BKGm
47a/pyaxFWZvzx2UBvAIXpvku9u4Xoj2Q1X/ugMkBfZVqLccZF44M5HZp7sG4oGuvzwVxfVCKCJO
yFCFNjEjtfQRNv4b2HPB/rHVXo1ImJ6pLkZ73dez3dad3yg5emrhafffcWdgUXcJJ/blunhalUMd
JLCRUB6n0vdPgSCQUN98EbnDMx/RaTjUBZK7nUuFyg14zD0Xq18Vcw49xxJ2fXSEL1s7NC+2Vhi8
rCv0xN+lNUYdFXgr+MwlM0nh6l/amcMDQ7N5hzwP28MOEnHVKCY1gd2J8qVtgoYZOXWlvsl3ZI+p
Ug+jwtBNHQu28DKtpsjElYCbjy4VMs2mO6WSLBe90kfhwFUcr9bEkF+XM75hi4CMh9NA2IwZMbub
WLmHdN7Xim8LbrM/Vbu568p8fYp0j6NhtBYsVsfrmsMemyK4C6EaoFnvR1JX+sQczIcO+DwhV1xI
Qrsek9bYdCSuI1nJ+dLZ/KroPbEoXXIqFsa80UeKXmmiFkC5EeydL9GzadD7fkoLOuliGpbv6XP3
ulDVC4ODMDXgsmdXoAgG+SejJVcGytVGtz3oMAGsOxlqSMwTH26bxf0djbLOv38nYxg/YxL/jhAD
ToaeYhFaC3ne7LoOe02Fxr/spahWiKAt1RREZkT4rdqgLRPE2RjxOtTtZYJqIY8dhWjDlm6hMU5g
DM2aGcUNpLAlXFiqQt/h3GEkt+TY242mYHeAUKK5IOnu3ws8b4kGRkVsP7HuG3WBFdzsJ34+JHjf
uv6jYkSsKe2nSucv36KHOR6zpE9Xyo1Jb7gdPNvyd0xTUOGQDPwmKmMI3emiyymml94/0yn/e/RG
Mo3sj7+Wl1dETE+x37r2Mkl5+IXXrRwkSUfMFu0+2vgrUnRttUUTBBVbIgC6uxOIEa9Gggm4B/+w
+kpSmLl4pr0kJZoBVC3PM+POzheeC8TTfOlGQvwYwxfDH20vVEZjHr2hALZSs6/YfwXtSSsTXZY4
XGNjrkqZcqEnT4fh5q7qMSuIkNV970WYiBQh5WRvaALpFivwzDsvBFywZyKie1uxsFLvRxpdZJ7y
LfWW5Z+dUJdFjrBiUe3ddyVYotcyOkOKvcT0kmMQLa5jm6GZx30brt26vRYsH9jSYKq7BPFfRWmm
wrpiepiqsX7TcUelBTKjs+FWdk7rLSAvEDphYixZYN5Auz0rYEdynkUn3d6Bay1G+a/vs4kcpckK
DBe900OcsyUOFSRUKqMfXh6sVnMfWT88q88cRpqkyJZYtxBQUR536PapOwe022sV2qUHICOg9fOk
ks4JTw04mhfFJRqvh2tlkhfBSf1owGLUrP8TzNlCyA3xr1pu9+PWGl+gTJ0LpK16mYOPDH53GKfc
o+/IZCo+2RvjFJuxShlliXwA4vXv9FHcvnxfxRB4JzboALDn65GhF+R0FAtnbGfNVmHUXDXl8UnJ
nkJIlWEuV6/adHg7uAoFosIk+JR4onhLP5NX3dHF7x73/H06NNEvk0Gq1zeZ1R8hFvIs3vhSfQSR
SgBUqhO9ZLaYB1MV5amRb38JRietSUzTKcgymdeptBz2ZunzzgqfjzY9wyg8tydB3PVdEwqxHEG5
BKrDDbacrm4aN/7GFJ7AaMsfwMdKn7FazWnUw4TyoUC8blC7tCycrlbg7vYy+QKUDsCZaHGlVhrt
I+MN22g6bd2ul0KnCbWxMm/uDCg1cP0QfPz24zjy9EJTAjoOlHYnJFiWyl7slm2Nw5FQr0KumWNB
AZzIwG0XaYsLZNjtnCC+e3PhsgXwNoDs9qBvhm4+W2TbTGXUrw5t5JGTH9vtZyy8IKjjuoCs4Ge+
S6NXzHd4sjW9wOypM8qCuuCgfSKfh0j0pDcYHFVj1vOt4fHXBQaZx0J8C6d59Y58DA9Ga2mRNVQM
qnQEsjNMoYrqnWVBVSU08HSxaeP9V6IQYm5GGvdVHCoQc6pSiI16wrX2z75eiX+rL9DQYa1IQZXh
Snvz1XpBzTzsyxsqWvuL0czHTshZXMxPTGfcT9NYKL6TXhSuoNleucw0bj1LioB0vqeGntMp5RGk
reG1FT1K/Y+U/wPTo3PfwmJofrq11ntHanWUFj7t2e/OnG4RrdyK3JtMRGZ7xzFULyvNbf/90+sy
w4UnVY5uJfsDH1TQmmTOIlzuj690krgRlq98CEUPlAWcXwcKkaZLBuzn7I1qdyohyna7bDcAkO35
9llUvPEcUKwcl01OUX+z7qVvfiBTn6aiAh2e7XF4mnGxjo6zrl5mwnD7SSfJwMZ7HUvRz4wZXC5R
vp005YrzBVlY+3XMhzhQH8njbcQfJMq5mDB4AQENqf5Z3Mg8ycc2+5/RE8r4c4S1pJ37CTZ3oys0
yA4TfBtiCHjsZ87K5xkwux8Q5xrvXf46trUKwXPxAlvvQBMfQkRBP3ZN4f8K2QQ8BWBtzCiGoIa3
dY89YxKRxHnSTlGb590BBLUXGmVl0p+Zblx6NS5TvlyN6HSW65wI029uUa1wpVyUp1dX6bUhabrR
fAkUuYgdcwr8v6m3pcUMknVx2BG9MzFDL2q2P+SO6rJKTzvLZ8PMl7kzpi4Fx7DGlY3Oda2hW179
yxF+zKqbCzQKKY9cjF8POB5p2DNVa9f9lk4qHrkMSymUV8p68xxXgQWwetI5pmG9Gr/lU+SjknKH
11+OhguMM/F8dc11CBgaYA40VhZ0Ik7t4Kzs7XYsj/drj+v4knBj6IHoRN9jDBYNcxV7LYj5EOcb
KlbDLrfwuyIIaYPiKcWeZZvVHZ8yLkbniqKefiaEj6n0RN3ik31rx6CiS6TAi/ic79DBk9xKSbLF
GGwd5FrB7RRNrZulx+QSj/n7IY5SRGiXc/ZhPhFWlqlCSnTj/4IttSSfrEYJWXBXhYX7htzZ/UGJ
cds+1bvILN1eJUzR5SI41zf87YVM0rv1wrLwOJIanqf/oDjN4pABOzt5TRm+NQI+ZsfQunHX4NhL
aa6WaXONnpumvsGo74epfOPr4va8ggRuiVAIi555+CvugglcxSSV8l1IUKhG4bek79jsk+zGVKCS
Pu5ulEUs5IRZRdQSr/OYeRTgZotEc7h19R3J/xD/LuWp0I3/ayKptDxVvs0IzsXRdZC/2VdosywL
ogwP9cp7FW7TZd0EXLK+dI5ltIr0nkePZgvmzBenEgJqdapuHM9YEYKn9X/q2KpvJagTbOniDi54
x180+L+dn7hwYzktsZ83U6kxVaAKjVQJRIMtOb8jY36PG3yyHMQye9myMQH3UY3cI/rgYbAy9nxS
ndqVU1BCyXqt33BolnieVQpEk3D5V1cupsQj7alytanodyG8vQ9rbVoSnu/1JcFOeSyokj+KhMHe
H5FkR8REpEYDaeL3lEv0UEhu5vsakwZe7/5LsAM20yR3sENB2ubTaDArkJm8s/7+eSo4chaiMCUr
q+Xjp5JNYamynSEE1bWGRtSMT2b5wOIACZUeNM9FkO8EOKTB5/FOREKIXAAS0L1V6ZfXkvpdm9h0
7R5jCyimlhApovJ9rzh9FUNNG45bdpTDB93LNJc1k1ky09nAQ5q8eb4xTFqwkAlCklVFgCAaKQAa
igJPhDRrYkNuSbFk0iQaczVIiaoRD4f8Cn7vSR2El8wIeL9X7FI5NsvBfo1kVXbg/Ve7dJi6lfzE
yByBve8Gi23J0CApA2H4C7yoJVonRMeJPXk4wrMsU2gRvI2e0GSjScrRxSPti2gIbtZUr/j4p5hD
YYSmq2nwA5YXiG5whtxoRC97HKA6WYdlQvP6HfZDGFIJltaMNrpLIwcVSKyC2L0tOnae82uyFzE7
xW5jsg/Aki4aNSJ6wXIIzbAzuMhZjxONj/k27V9y2khMUrThvSkInGcRl68RJbZe8DyiNlzcbxPu
0yeC8NmrbR5AbG5LDqWGlV2IWy4g404tZNvSTxbLO5wzy1+NtcLkKnv6n9L8S+lkfbsYJU/q55VD
7cJP/DxL/LI+Iqm3M52oAWoCp1YDcQtS3ZsIqaQ7OnyJuHENFw9rMNR4T4Pfgqnk2Z9dAuWqz8ap
90rayFekU7iU5qHAbQ6y2i5jmA11xlgCnbfpQxlvcpYBDd3zFT3qXSZjyPX8K34oySI9T58aGe9H
0WzySHBJLBJv+1UQqy3wkzc9CAAtsPyDOIJYGG7UacQ/a204VGLYFc0k9CbJ/3g/uUpg68BfdkL+
m+eDa8VmqKf0cEKIGKR99PsnEcIzq7QtQiCi1T33MHeIBXZFIttmuv+Ggsd3gRooKh45N1Kz3fSN
nP1WDfOUMjZ4snIvBTgn+xowJuXOuPQBxj/av8DqT648m0OEaE+tF31NpakWZvbuyduY7TvaG9eL
Ym2A0UH8WZ3qKQSr1l86WlHJcAtzDOZxH7UBDbAiVtKVZTAl0lOpNCfD/3lOuG6QPCyYN25hd97P
hxQkwmfWcmkYhsl2qcOle/NcG3h9gDl2U/prRJJTx9XjaXV0hp1Av/j+WaNCfOhWJKkW68UUK/2J
Cj/DZaXr/rtsMY31W+w/hzPCwgxMWgsgn8h/A3Mbgb8Gz5r2AnaPNPCUM5YOUuWG8vU3GFe2hD6y
jqsw4C1uQ2usBt5jYgZUU07FJkWXO0ehEJvt3N4vd4lx3l9DJWqdmf2llH9nseAQGVZdmHMBMNqX
AMzA1pRW95SIOR2iFLFKUTBzUoM6PCKV+Ev4cs/6KhaxZzBztZjP+nSDAAu0TD4vbcBDKx32ko3v
mSKkztJPxSwwnUL1LG97MjCV5575Gf8m7/9XePH/pVmoJWV/QjEiJ0lP9BTmZhP8xQT7J2hSdHfj
QiJcswuV3Inp/08bwYGyKjig0M6MP6Q+dAZWdHb5nds6JpBVyBG3ywkYt4L4y0FKhs/oUPQZkdG+
8UFDO5fFW7V7ptk/s3xHw3VjWXa1D1taBxcIBvFChnWnHW6xYpf4izFNIldzJardTNbonWUg+Fga
lRfs2zy5aSaKKFZfVj6QFr0oqS24KEGoOMURKL4VpbrESnNkDDgsZ4BNpE9q4/seFsyxiQF7BByP
9BCbQsLtMSIPNx9IJTvIPt5JBB6w2gYiEtMh9uuEIWOlYh43CjZ4iuQEEHufCMGxpMCK0wEf3wQt
t3nUH0nuh1Gewd757jCsD9R1GxaHqslEQZsCHozzyG9JK4L/GGO+JvdV2TkRhzGGVnAYSnBi60ZW
78VLGwx5wWffwV4wqZOBdJW5jgwExzK+w6QZ8ZmVp+sjZHOAeAM8zGCE4uzycxrmVkRtc5w4+ylT
xRvhcbz7hOPlc/8qDoA68BaYCpJGxga3u421ewvkDeZaI6txHQozO0j+A+FZUvyV3/McOGXbUyCI
1qAB4//eIXPKTXYL1g8wkwv+YOnnvt/R6Ibz8IZLzOaCptdlO6Dd8dtCIOgS54OKWSdSRDnI/QTb
fj0fQC7MKfhDpgxmF/WzBaFc6Jj/6QECVNTYcqk1+uwtJErOMd0ryLCRXdQmRGeXbINu/f87YNau
hrTFwR/jJdZE4cAnELvyNVv67U7pLGdXFdOFQa61w21sdOgA8iuYLOKDRDnIDioxcL/XcVIrmxE0
N+EPRSvZy7RIUzwhbnTGN5NUVDSuz1HqF6jDM87Mf02XEua+gTv+cvGwONr5ZRv/USqaJXgFtyrF
dg+6mGcArZNmaCYAXZDXOyH0k4OoEa6odW6UZKuWDncEGvwU+DI0kecnXUJ/vuFkutV3tKq9iyg/
fTjZ0TdIxnkQ+Hk5l84Q4JDK96KFCO1+khwCGGR2ERvP4vcuvRIi9KFRqKCh+jHPZPWq40Vd+fq2
rcvZ+0zr6A/NVwzTLOLlb/mzR3NR8zYwQL/7CSfw3D+b2iJBlmSFhEgc0H0e1OuFhL9CKCrEczdR
wwo2PxHGCafmV19spd+OBFpEPOuLme3s2DFKWY7xfDJUZk4X+uReJKaN+7xPWmlN7xbMDa74Ey+Q
Y/CvCEOfeiSRmHrGr65vNXZACV6nwSItPjJ6xYfDxWTtO7nNim7vFFa5YbqsVmjv+5WGDEjOMFVz
ETllMhfm2j7g4TSX+KNjyFRCLGfxTK4FN4TtnsA00pAbgpL7VNMVUa0wR3fTsqe/1ZEft8bhIt5g
yRXvAXDL26wqcSOx9oZZ6YCAUEgXx6FvdthVPnU76RTdZEJJonZXe5+X67MNqO2x4zjsJuwvqE3k
6L23yeVfPyyAYuw2mWuiDcTd+/9FV87PLKdCcoCy3Sm1823XVAv+Q2RSQL+n0t1VGww8wnd9sIat
JZFebyW+pPBb3S2Cih5S/1RrltOldMPhfFeR8D6rpRJS2pnz971JItpL3gydXD7AIay7idD/Ya6A
HgrGdf/fvFrucxoaK8OjvOTiLdv63S4BzKkvcUXSp2FwSXLdxhsa1zdyq7uN6HFH7zSKs3hibIVq
kyc+RCayG++sqNsqnN8UE1+FXA3dwCJ2bGIHazPmCABnp4DusSKBoq6dEHZXLDiwklj02ZigNmx8
88fmxDuYEtHp7UDXRKQvE5Ibb9wfiqJ3356JvayUujBDAhQQQF0iYz/eYba82MASEBZIDd5y5xtq
2IF8VGJHYt3q1NeM1CXU2OXQ6mB68NAz8/ccDzeFoo5GavyIW8gHX0XvrTrz6DYIVCIIst4Li8ln
EDYbBhGxawkikahEjaQSe6vaPT5YsnvuVDuUOIo0bE1EnhpZ7t+mrNfTA4avppcntzCa+30oJsNk
Qzu8MGe+aCNmijb5Vw6tCRW57Dpb0WVYPVX3Q70ZDiLnd2Q/wW87A4TCjS09S+E1e1cLnYLEI5IG
yv1CbqXpO0Vf1o4K3UIyF5OkX5X4P1KsMUQO5fcY5i18U0c/U/Z97iCXlpTC6Rs6D6q35Z/vaN9L
6pOhzPdt1ySfkKj0WMEJukxQYrO3nq9OIX19c9fZwxlVV6ouLhKskRteZxFzvo3uRNtqr4OmX4J9
JCEWFwg/JPd6ovyQC96ZhB9iPlmgj8L3JV/sHjYNhRwGSeuhY0SKECmjmFF4bW7pZOpFBYWPd30q
21tUdMsFXcXwsSseD3+5S3untFpM74yofvPurvwTytXtU09CbQ3Lewo81a0HUcoQ4Iwp4xfp9mxt
f1aR2+XYeHj1CfZZ6ccHgONsyFiu3Gc3Wa5lWXQmwP2H1CL94Pq19J/bb5SOGrTw9SY15iZNv1GG
rmGnLmgMJk30cyPpfkS/DnnyfhGt177iMKVRavh+DDasshDGzvoNRydfPwJAf3OKYX9SDCBXHIdT
1ZTHJxD6tokrwWUrZln2pdsIgujKjm8LWPGOOVT6W3wG7FJRNDp0bLPsEsM3vUR11c+fq/Gc0Mil
D5Kr9lGLy+a8mJPslh1//Co66Q/wENDwJLFM1tFsZE3vvnfMLtO/zptof+GrorGlRf2cbtgTc/1e
fDq3odokdZ2rPQYA/lGGFPo063QiLTSM65xgojFHu8OOxZ4J6R4P2KbCPSYbgfj128yomoEVKNnA
B0tnKmMYec3ED29BGx+HOTWgTFKo5CJwnzodHJsJxcMoNix8E5KqPIhh2GcMPQqOzq1b3MjviEq+
3lXpOBbOyMBiLQlba7mQwbDzc0tFzzq116SpKvsVo50u2YOK1bVKpMZGQvpkyp2IJ9m1G4OyLI1w
cANWgxX5RoOD+47jMGGH9LgcMJ563fXxA+BHSTyfAbDw/17W/jLDSQvQ0CFPJ62iogPVYpc7xfxR
1+NYKNzBgA/lRbG0Lv96z66R1FE7pRyrBfxrzyu8rmMzgYHS4/vfX8cfLboJ87qZaqhgHjzu40/U
4Z1FUxWQB80uVYCo/4XyEtoSfK5OQ8AChGiAhh2BGSZ0pUZTi1TNsJeOw9K+WyytBCwdhlTIcuiD
Jx/2f0mQafU46EzkDzY9DmMgmeCPbzhwEzP2pIBCsZpx4BpVbmDjQfVm0Wh/wAuFz/k40dS2GvMk
poFfR+r4yxsOgQAq/eSSjVMP6KHlZ4d3L6OPVWDNIunDrmBw9Y+8TeTdYn4tpwydMMzUnET29zrB
YmQTIDi67YXNjT7Zc/kAbRhJ/v+ciH42Shl670i8PZUHChV4cPF6e6yR6EyW+JW0vLgijVOt5xZ6
Zq+JzNDpa0RyrkAfpZiWqPzJlSagttuHtiWoo505gNz4F76PCahnvnMNcW0+GXcO1Bp2SGp317RW
ePMDsWz9tX5sCQbpiM4SZMfg4A5qCZ/9xlT7Yw0a9b1IHYq4RH+YIqSjaV7MP58J95eI7GrXcqtF
to7LxjMxoRHH+8Ago756z/5GLziNmR4sMfrzQGEO7abhdl5+XoND1nZlYaBVUNwsktoi5DeujVjF
iXoMHUCmObNmbcp/jIa4XpY5dq5n58dHL1rFvzD1+IixJ1RLKojjXflMDmg4npEPtoqLyUehDzVK
vrWAwilBBHTVAsu+fXlofPkXpEn32r9Jc+EWQpoA4C/q7Llr3RS4Ajccjs1LnjbuimJKaIH3WEEO
7/N8bvSEd56y70z7YXvXAyhJsF+amtJb5nKhx5qSH47KHFD8n1dOktbbupSVk9wWeBeCWHvv5WOE
4S+GOlVLnE8X8Y+iY4mQXhcunaec7W/0XLrLyaWo7cA6uUDqI1blkRUkL3T6/XFH9vu6bhLX/vym
ohEbw5Lur0NCuhAves7Nf5UPse5/ZxovAHBUhOLkF/ncmLFcY8AhqnSRXXSqa48mBkiaV5wWuU+C
g78vqt877sZyM7QOEB65pXjEsUJBapLOQSmEM5ZDNHREvv1q9c+nT9a4a5hA/3P4tzWgTh9gcL0c
mvjeNYDSxiAzj4UoQE8lG7m+BUupRVBEbtre7604+QIewbf6DMQ7j6r94AnOBjY6c1iGeE0lPDsf
Mvj5dPZNOIqS/67sS8Suu7rbeomsDf+UUsyh0sJgSlGdsmtWzYkwctjAGtwAOBZRCJPCfPk3mekM
kh7IsMnmKOiI1auO+kB/Dadp+ktbsl65hxulw3pndZ+f8R5oZV052kNqmjb7DLbLbYr83JeS1DMt
VWI93FBxKAX2qxqtbOoaSCrkcJfclEZ0tGgj3Sgivh76l0QXp167LdgHIbyo5hpTeuzlfEKrmznx
i+Z1S09cwkR/KtwS4CV8B/X3kTecUyFBgLslFdz5eXb8mBmdlshccdBVwsYy3i14/RUFqUI6IpjS
XnxCxR0BDJwNAIq6hhV3VnRhf0tO/aVxbMqcOWuQNU3LYXawmwE+obTXu/YS7QCdREmCXufZUAA1
t5PLtFB0WOKvk3q5bqGv89bmDnZarapPsW1RYVtjSJ7vemOsn0ihqYGZfjbXU0XSmelt6y54gqGG
7u+84e++0s64M9EEPjS2jVt7i4dxd37R+FT0n542g/WX86/4IRd3aDwuKkM3IGmDwfHCP06qu6dp
RbR7zv0cIYbCtmPZaICjSmugOQkyE1n/Npytb4mZwHJqhYORb5FUht+FkNgkEnFNLe57sXREJqj+
yPEi4BuW/4zt2+thGy9Z4E7jG76Mf5qYQRRfd1Bj4avom36dR3V1n3iVbeCx+ZqdrnmT7+Tzh19r
aZSrNOO+uF8SMIw/BZrqDQSM7/cHju9jYJaNK6qzbUpFkafFRItOwY4OrhpHx9Z3Gqp1Il8nUYSL
glIFf3EkNztCJ+XIkjmnNrsffhjyEn6qRTkSvFiEDy3ru0IHKU+fLsq3nHjNmxDWO6PPz8s1N9N8
WAvgDeteIXQ7EhEARE7cko6XEWECkWNbxA4tA0MEqq7P0vui/35f8phcefZvqKwo1yYOo7gKYGeT
+HxHzMmfBxq9UgyQAaMoxGQkExSnrlani9GjkuFn/gLg8gOraf6+SKHPP4u9vvWaTNFdJ3VlQMUS
TiO2aKXVMscSEWEikC6P8k0N+nfAbzWqTA0B1Q6a/CqGGHN8yJSytUjRBmy6un70NSoMz/LxCqVB
4Qm8OjVkSm5RmjH+ZHUrAXcabipe+aLcOa9ujPt3wikRuYJAUKnMMhuAfKZfNkNh89Sj7sgwYvFe
FO+KfCjW0wzML0alpAWzO1OY5f3pIXAE1Izq0AIxZVKFxvp5uq9AHpJDGNqH7ghQq/HDVY0rtOBI
1QFWKVjKXfVKa/HaNrsypRNsjFnxbMYC17awtvE3oZcIGPELFrDNx86D3VE9lopcBTmE4kZR/uVq
ujiWizm77Hwqs4qqq3fgl4USphmwNUzwQVIthQK1udxFjAYtemgryDNHfg/YqJdZiSrLqkA6nmBQ
kIeAPYM14aAPQdL0HsoJTds7GUezqkz6f0Znwz6WSLifLOaU54ujVWhGpXw97oCU8MZPs9dIYcCF
Z2u1sag6vsG/wKyYXmupwfsgtC9CRTCRPLtBkS3iCT1DsOUJ8AIyxFJtEkOlnDeb3fJnEcoe1CdJ
R1H+PVQewIyP3MYr9OsvJY+NATZsBxRaWNCinBk8iomkFyYw7Wi7dEQdOKTRCHWOl/Pf2KT2oWyQ
DbWmsQyQ0rOK2XP7jUcG74QYkQguY2zBr0TLH4ByGeCJQeB7rbD8KO0byfbY2kHVHWGcKxW2BoNb
7kHzj2GqU8G0qDsoYIUutzXTJV0w5FO+5yRi3cuDqnSe3bCNeYrsyKXxEJyp+fyDT97KJF/li1qp
M7TOPZAQNWixxjsIrCdeKzxn+w3/3QL9wlhAh3tzyYp32deeMMzcS+ADNM470lX72gbs+Z7dO+b7
AdlnpRTiONj891ja7CaWyAywGUUt81psg9VeH12Yq0G91sGycSqu/WOcwe4xVlxvfvXpAyJ5jOEe
XU4a0gJ5pi+JKFKx2I4fx9QkRynxuRlmmk+zKWDW9R6et9lM3ygPSZ2HiOXBNpi0AoKwEZNVQ6uL
6rma6GAsQoVrUBsaaDsCizt+GRpL5xKw7MJ95a951xv2Vrg4WXB5RBm6LNfRZhoK/vb4rvJa3Fxa
P7UBB0dqHLo0ESQF/eLrbUGWQAuIG1z/KqnADvfyp+3MPZsY92LeSkdhMBe1aFI1vgh9c2Ws0KYQ
KaPZZQF1IlHTCxI7TjtOAQGbjQjalZh7lOobFHPy+/dtBcwKi/n89FdKvsq8j+oITcfzzT7J2kWy
K6sECGlE2kYQ4H1Pp4CBfcZcX7dLgU2b2HvNyuA8cbA7Wyj8zaUDMv5x5B4JUayQFmTvKWC+v+DB
9xhtbmoMn7zX2Zzv3a0pMGWprfJWxytc7nyXizWnZn+6exNq6dOEYBp16Y+nd9dr37IHr+wktbpl
sVDQd5oy8HXM1toWcqz5dittVTtwcS1zUmUROk2SHFcsUkvxXui5vL+PgRNN+3jj/luK7dtCG4sV
zK+IDu2exd2AtiXCVbDAVuGPzPBjW2+beCroclkkph5lzi7xg6EsYKFgndDzmr30katOFF/kyLiq
MmEKDq8lBYuylvXwu9rCf1kKKCqsINSBIjIEpEqXdd17eP3N2HSnCD4jjwY9VOwWhOCFMR9C1mb6
2SRX8+yF4uwewY1bi6sSBFlkbgeoWbHjB0pT72UUzgWb6rPCyIYqjytwhiJegJnDv0IoHzQrhwqJ
UIJyT2N140Bgg3aYoKgQa5OpzqXZeP0qxT4v3k5PAochcxhgm/vv/rIn/kLpCxpID1mJMPgv8bXV
ZBOPSIq4lNY2UYzuujXLOUH0MPPvHefAl/Scn90u7GG5gCdxkHruADJ+MRG6GTcnEGq28DH9lstZ
SjKGxFxtNlg5c85xke586xkv0MeFhY/dvVZUU72ws3xWfWGMIz2hMyWyO2wv/I5M0/uG9ZStxmQ5
T62E2b6m5JtWJqCTQiepFvECwOxXNUxmiArYyIiG/PNxPdtkE+f49WosbpH8mHX3pq8Kkm47gEBZ
cKCNadbcnVPIUzqejxSIsjeQz61m1TSqimnqodHt9z3EWi0JbQFOcnXj/qaH1suLO245ng+9WQq4
YJh6bdTlaRkEEi9EiGS1w6UjpNt+MZnHPULPazaEPETS3ACn8F5kaw6roQUjjn2pgc3abJe+q9po
Bi+0N4SV+O3zE3LU8jT3YYtVVnIMvQn0AsXWYXGnEfo6P4Lz2LbOAjMAOozsuktU6fexd0yqGcpq
ErnDx65s/vF2GPom+YJbr1NXjpNh8/igDb0QAkkGoDWLzQ6MadNr4ilXQHX7Zfb6mSxh45wEV/AJ
Yu+unWGnJzgynGY1WYj314TYu0+AZEL/2N7ZHfqtqlOGXZkgO/FcbxdQMXP/pjLzlTGJbPqjofE4
f4jHVmcpG54LooMonE3K+Ukf20NzNVK3M4bmsz4mPzVWfW/HPW1IdpJ2jJL2F/nogOtwv+RSPm6g
3WQ+RXdUQ76sQBaPX73hXmGRiWKC7jRfkgP91ZmgLv/J9llCjZdWltD2S9dPOJ31+Ka4OgvaY8VP
7wYRbeObN9nJLx8wCw9RY0k25qHosjIV/6mEnpoqfmDodVhQzFaak1eKKxgiXAerBfPgt8FwNW9F
dYHPq4q/ltXbLh9YaX+m66LkQsyDMYd4u35f0LbBAgNp47WIpIzBUMKFOINR9DvE/ovHVZWKGkvw
w5kjBflNRQIEYhWPYEwSo4HYWewFA9CCZb+JbiTE2zt0E/8NMzjvjhqgGkBqJTbC7VTWYXddSjNy
cyMbaMzO95B+uVOsZfdVlaEmNDWy1UT/SqiyWfWveYfyp//TOcNR6k2ofdIU0RJVuXMlXUJx5wk5
XW0Ltyyr0wu2kSWocg9O8z+9ziKj7go3PiW0Wzpl/BSUvOophGKeenk0wJpRP85WJa+p8Vjwiile
kQi6gUDz3qzSp1nq5aLFj7kw6BzHvzpSI3FGjfDLH+nVbSOD/mh4ndcyWBQVaHGTxf4JAleuVtEg
Rc4nknt7GwZTNf/zDxKnSjfEmMfE4okGdi16+XY4+AsP1p6tXfsqP/rurKuz3d0ISM+oaeSmS5cV
0WBwZSQH9g/fL0NsiSLWAS9yz3HA4SW//YtgK8R3L+FOFZ2PQ5KBDve6M6pFCd28oRWv2X9dMIcB
GJgXk2PTxoej39nmVR7sJgyibM/rRhUX5i2/8AEYfAm0e+r/+NQ13f/5eR8kGS+N8eCoHvZNyeiI
fzJOa1EM4JuhcCAkMr9OlIQVIIeDTyvkxzgN2OmDnkbVVKT00U7tx/ZP8EyhqzUoMcFrvDlkycf7
3Msd6Tdl+QmIb1Mj6dq0ANkf098FGzBr5dDx8R3JJcD0SO1eA2rL+iDSLwNiFSlz9D0vw05AEBIm
vVtmEXQnqGoUTonHuc0Pw7gOsoBhaothhNaSYUHNz4huXD2ok4NM6HxCQ6HUImH/kZbnD4uiCNfJ
ba9TyrsLOj3cl/i7M/sYt1gXMSZJu2Hgth31rtSZBHvR2FRLByO87YgGVgLNa7Jcq5KKSr2Ite8a
ae8Gpof5kxLofXo95WXowgbPA1Uw6Jp8i/SqtL5Z0g0nl6T5ujT9qx6yThU1c2ht9yznx5D4iBUk
f4CligHddf+rxankc7A4RS9kQOWQ5akb/Rrtw0NVYqKw0BtuhrOjPxPMAqjHJijcOIlkHiYCHXmm
dlKpPoxlfH474cEPODRN5VvlB8h/7iCCeIIVgwzy9TtIi79X19cToci+Ntlao6I+mG1EGQeecmby
jtHnjHL5Zz5q3Dt42xoeDCQoKJH0/pvN1JsPjPweMfKLHsW9rkPNsiXEkvMp9XVFBrzWDi7rkxaa
PNy35Z0FB/luZ5OX6E3kpKDPYYcqfRRR2KvLgDKWOBVDdbxaIaqBS3h3vmq1IYBrVzsXUjiMvEZB
HEK+jbRquCSJo/WNss7FqIdTDVEShAmrZzyQy5zLvVZaN/uvCIZKzH/EVtiHVPsgN8CMXAaSn5qJ
iOPSuz0Pn/ssAhFXPkyQO6AUWGtBpOiamSLJeiyEQdQhweWSfxH+807jW78JsHiw5TYV0aB1gzMp
u01KbJiJaBXiaKuVPBvkTUoP981wECvFgWI3TAJmo0E99b8gHyTm+NvyEIe9AIJLchhEsgaA7/nP
JpW3RWY0kwmUj84iBY57EKEUvyz+B+qaNqNfzlkwT0YnYsIKDC0Psj4+v55ly4GHK8GY3DLNViDk
fcGuHAIjhjz/XOLW4O+J0UD81pS6L3c/GhJ7FFG+1CbtK9jKKpG3NhqZsz0wEoi2Drqv6DL36VQb
BzIZMGnAg7t1fIfZoRAjIgQIMM7OnEfz7j4SNPnBcb+gtRAJ3iXVuMhhjO2PwCsorZU7J8iSmlkG
qY1XXRdKGotXuQZy86VQrr/VXUlcifZAdDSJ9WJqHewC1Ws3GI+VMjGu0NQLRq2Xy6frfvSBJMb3
JDjFFhbvf5hjTM/vEOLSgwb3QssNog9x4T4u1TZ9chXKYprFwtt1SyBP392Zani6PiL6XJwiDc2k
3UxRMeWg6+5pFEgmfhpQs3pCWL+w+X7Oawe8mXggWqmDCWucsNLYnaMVaFTfkRH9iDMRpJCK6ImY
NNhoSOgUKMdmMWsONkWCxil23L4NhKiND7tzmm4fNLfpya1EbpQZQOdkYv0PC1H5xq5uabTgi3VU
FDilEmpf5W3ll4qj/oX9qfIXNdhpHuYa/ochqH8el4VmwUm3hPPR4Zzy7p/v2sDVlzXA7zcurUo+
cJcg2W2plgSDr1TxmSPQqWpBS/yIbxZWmnmxe1ittJ2Y6lT5liF/9nlCeSdUioKiCEpTKsAheQh+
eGjcqLuV78vYHBro+cqEP+huKHiy7Fm6VBN2kDznXRwR1LsGXMlzU8n/pRkQ5CA+pdHG6d/XvY+t
wqvRRwzCHze9XEVJYPRiiTZR/QKhkBEIwUbZ+m3j8qTR6Y2GBjJ/rEDwfiusI6b3u+tDR+5F3l/G
gchMRsKJ1r+WIyK6f/Il4THhHs6QonYcqzWbYbeuPRcDjDXpHN6G+kFvWt4Sdx208HKKkve8wowS
exVklgXTN9VlUUZTzyD7TsfKipEczGnpbrWUPYCga3KS8lhPgBR1pVY9p2wiwGE040BIX2r1WBn+
5h8c15i4QRPj6yqWVhteCDJBHKIK8VTPk2t85BANEuFJGEsfRdB4g/5E8ctMhzdAr1n/M1jGgx7u
M7a0rdFC7lDhWkWq7Ulv972BOL8Gl4RDxOZNarJ0rT50UHWnunb4mOmYwafynD+CgmyHYvttO2tM
uFdzhtupZTLX441zFX07H85Ucby9pZg2ut0xXnmCP0TeJY5jM5hK4uyubVHMFAeD4CrdCi2H4Plc
UGQ5PLIYsFnRD8vft6Oxp2LxSXZw04zM7Nh61qSiOZaOdSvOQr46xp+HhY+XnqQ4CVkCZKnhEPUo
DyjzNFdr87vH3MxMM69lX7Pi5KnzvaU5pgH3whbTlUMhTek/ADdkY4tKFVWJKvxBKNYbJId0JEFG
5TgiR+IhezsowM+0wMqyc7Tau8KEDAakCs5dMEZA7ieGUOyIMj4EVXAQF2OIjFYYox/iZ6vUbxTY
p5s6aiDUwLa/xsT9ph6MuYTDtnEogmUA18Jd4LGCBl/lKPIfJ+0mzxuKEObBjDQOunUxmwE6XNZS
tQHVb6shxs/mfar7JrFIlAHTdFryp23SLzZ0z4ExGVXQq6uj3jbPPslZCKMolMudASXN9hCJsiNR
JqxXvcHlAGYfbHEQVDmC7lka168j2iLfpIEdLrSJR6ap16IJA7nGHa8fHXn8NRtU6JpCtKbUI8en
b4rTYyGiHFAX9pHo6nZWO742OGU59XpNNdTaC39lCj+hertyJWfeOaaCLYPFfvF9bG+/eDf4N7Z8
DDhqEj8bnCmImARYY0iMyqX4kCLRjIzmcoLm5siCXazIfzsOrVWBpPzjdW+2zfHZ+3t9gFe5RVpH
AIQ1P2ApqqJDkEnDLMFxZRnnSeGPKHIPouYCHRFPzNot8JsIypcNyN2Hp9PnkmnoISv1dlgXLb5d
onzJ/DGVK3CcfY8ndft5VgByfUAPNUx3JgxFb53CpYCcQEb/U22znkMpRYv3uW+aXIt5zliudg3g
cXUQ4/cSjv3CzzwfUwW+7XLq4qNSHwwK4Br6BSGM/YzeV0kyO3nTOxNLl+wxcKkpAs1lOZ0H5ECU
DCweQNzsNshTFnpdjLAKT47b/x/yeLETviM+hcWC/tz8tjw9VxQNOFvWwoUQEUtk280gfu/yGN+C
pxjtnczTuGZNh4gqO13gm2WbxevEnG3WDlvs+K7/jV+w820GYOoaJgL9S5WVAuMI8yGN9T02fGSZ
Hz0NJd7LQU/5c9XNRt3thLA5UN9gDnkUZvgSs0lKpK8VXlFYLMhkczewq/XqZHV2B72YH7sRjcrH
JjT7jGLpi0KHO9svxmjDdrZ9MCNLpGs5X9InGsaYj8hnbeTbZ0NygN4lbIYANLUyAi5Gev6eRfxX
Y8QTfZPi867xCytlCG5VycAVecKG/VJQjlztbJAEqkICFsVPHZBCZskc2RFk7c6MpKIdikHPFhOo
m+SorSGu42pgStFhRCqEMPig7+XVUaQePhmRbvNUyOR9sF7vPhJEoR1GCgxf84wJeL/IqPX/tvbI
Qnp2GJM8loOXc+GnMySxbhmdYPXT0uQHpZJ35qm/6zkZ9Owg+H2suusBryBFPWtplOKTHR9n7gxN
3hSqI06nN8b2XRGs9JPmpjSURj+6sknKEPMp03i+3qmxXKGeUxtI0DdUuErJJyUoD13TfUgYUF5c
WnMvpS/UCUIt0HkGssJhGusfGT0lPSHEXkWB1tQowuM/iv/94ccdkU/x8SqgCFt5aX2MQOrvmna+
ROxYj+cGZ/QTRngmpXbw4gyGMxRdwNcOI2ndl4AxgmmgR/X4vyuVOS25mtd3SEfSYkxABB56yxhn
J9zzoY5EsLJ2mi7iKv7pSjF28Yq6CFrnpPBswT9VZ1uG6DwEssRTmi4ogMgKzgqlSicKz/aVCWl+
4LWhUNt0Pt5a32JopTZ7XGLI04ThFLDfyhVm96544pIRy/Mm3DMAe0j3GGPzd2M2w5S7HTaX89vy
b9Mkaq6ByZCe3Q2ZLZsC/MdWfVBhSqkJ82qufUn1iekh7+hWIoA4r7Q2UUfcAwyztXwqftmYLWhV
4Yw+pUOAm5i5ntHKta4VKIFctrDvz/230K6H1oinngH0b/OX40vmAzrqimx3NoQsJC2JR8851zgH
xh1CdjexbnJmSeAOreeRHNYDo/0J/T03J5dUAiIgUJQRcL1lfjpRmzoHS/CWQR+0n0Ae4UerqYgm
LpgTlfqs9Y4gkXroTgXMzm317NZrirQrvTkiKKs82yUGTvaenZG6POoDkV6/AAoYdZj7n+ePq6IF
0H52DcA+nFbpCW4rCRRr0KNQ7DkRTHJGX/fvxZ2nkWYowPtpZnZfpp8WFlUkci2y0RvsUk2K1nL2
2WWmXo4/e+2G+/tBn5f4vxMVVJ0P9PpmIV3zm+nYuMOQ7cPslsum6kbw5JFFYJTD1RmYNWcUbanp
CG3E6ft8sZ1XIWGArCIFMAeos68MduwCDMJ8Vw9Rn2NMS84hCEpJLOxOAvdhV6oxQQ+amUa4UW2P
sj6z56o/3wMuoY0Dasxbp6fx8/J5YJ9wUK4O8zazkxQOvo6GFvzVFMIufSSnjlREz+/E4pijWzKr
Mk8vnfXVgX24xHQdPujm64h918JOpxTZE7NRZ4yun1BgtXx1hEDjYxaGolqv78opaOoFC2SD3Lw6
WFvfUtxgt+g9EnSuYyA9agGHYb1TpZLCAck/t1LPrpXUWd3u8GNaD3QFemXZ5qPcZfqYg6BF16cT
InGRdA7ByyuiGpu4eyX9JAM86vCj7uq3TtiamRloLZL1wc8CGva81+ZxVoWB9JepgxhkURfgfkXC
ZLqCXVIHOGE+qMAopATqCzoLmuuPKHfM0120HwsjW+RMN3V4JXSAUyKCwLRFm731DBl34aD/tF4n
h2kSqxs76GanH6HoHVuDUekQtUnEGTEai9gDU1WU9ErgG1cY84q4uiYoKTr0oMV2HgIhwj1hGzWi
UfYP6NeQafuC0V9SbGwou0/9uHTQvo9wAsALaEd2zjp0YxWAe3Eh5q7vVnqo72bKfifQ5zANGnUk
OVTaH5glMV5QeWES0Wtvf5xiT7Bf4fJDtQIta9rk83KNKgBBtu0qLM6jPsxKRuK8e/oSZGEyt6cu
7/DNDS8GuMd0jHszzOIJ5sl35xLC13pVbACzZaQ65aaITBLIm1G9DVUl7g9DR6s/rPkVFWf1ujBd
BcFAn26jYcCYMfibxd4eolTvwcGTP1jesZvPM+R5oAqZSJW/+sHj35HlSxF8D7txG0zDSWhWVspn
SLN4+mWpjSsOZWXO/UtwO64cxDzii9XmOCpVzABhxUjxTKX8WFicAjcl0uNOWeDUdQhDixkQCUUg
JtTems0GPajzQ/KLrW3CMiYFXB+wpXihxVkrG863yDvYBJTSwDAUCz1x00w3aQnLsqtE2Tdlqzos
gp003Uukgyc5n4SWFCyWq68NLhBYQG75MqZkyayNy4kjL5AlSuWgWCd/lxU8l/YsJaZNimqztgAF
VOk12EIyQH1kSGnIfTwNePCDxb0PnXDqjBbSLWVixfxeqTYCcpWkrey18xdZK4CWPRTjuNL9IywV
3JrfPfMXw33tRg3bID0wg+ROpZb9Mee1MeBI04G2GBOIRotxl7y1LsNm14FreGV1mXod9f75SGAv
86lMtqPuBVwyq1H5bJlaB54WP2hqFeX6jeXTMD7a1NIIf8EeeN5P+UTy2GQ63tZq1xIgK/kSWq6E
SK79zQ6jURneErUEoE5gNYxmq/NTmCrsGi3ifVwVuVsys/uBgdmn2heY5ZSVYraiOIRwQBW+bIyl
tWAmXD69d0qTq06PXvfXyw+K42W5c7mSftVM1lasDtUBIXn9aVk1MoCZT2XQawHVLflDgXYyF+qx
5AZSe10V5sBpf/ndetOhEYdOwNZLjlU+KRGAwHtTL5xJFPHs8NL6+822sJdMmn8B5sfHRpfEeIy5
KPnYaewFGVwQHvg5UccUl9p+zsP3X2ZYF2UK7HuRKGqxy1GWAY37Swse2iE1j4MnYritYfTRUc7E
xHXsiGglKce2Bgqo7jXmSMgkcEEtgJDqF63q3+BwYwhP6jthkXLhaKNKFEUmz1SqNOX5FIW02gJQ
vc7eWiCKKJ9By7hv0aKZSPYbPqkAcwNJ1QtViYO/rcbR/layHGwLov4vyDACbxpng1L6XEz5AmRR
T4qA8NtrURQyWUNGV4s/4tqyrPOtaG9Jms6KrdQwGO8v2+DbbBub08ZGQqxMEMUIgf/M/qWd3ivj
Id1YWCSzjvKISw/uQZZfCw3IT3T9VTDvAmbkF68zMXzjumRC2AIPh8XrE/H/Vz6X3TwBKuQd4ON/
tZv9tmw/UptqaNDZpYtL4mb8hE864HFoGwXRYZHCQhu2DBUjdRpAhCkO5mfmMi+z6HJwLp6WrNcB
r0d51+Hq3FPUBt+gqXCBMxwtNLf8U4zy1C8ebfvlYYhShHu/wzNK6SVQKSJiQ9mdiRDmuIHHawyr
8M73x6/w7WwPlswNxu9pSbdyOzvKiOjonujLBM97sRvHXDyzehEyVnmQEwIeC3edaTeOyu2Mu4/p
P9MO9GLRS09SVoSW3zv1V62DOboypRyXXi1+OvmE9rjABUpXKlO4ZEv9A0fSaabT7vHcWOQa2Uo6
YVV/L4NiUzBnRIXhZjWkXH5BIYJVskU9qKThmu6XDc+BWzBtxHjuEwmAb8w4nMSI6VNMVVYhrXOb
5A2rSdhU9F0AY0EYHtwHEGg/75RjvOsI6XO2y66WF9FR+gmnrUDXw4R4D5zJTwfdnw1hdJJT8LEb
gWi2afRktjoJckNLi3/3myrJW3ycqdMgn37KoBA8tTer8e+p4hYc8m76L1kT+ZXdKHeCPrmVuYJI
3O2HcM/3O5ePxtXRnI/94SPSH/00jyXtPjkaKkN1RzAGZnbTZ2crbFxp7qiWTrX9S3m8vgA51c2R
Zv9loa6Lh/7QFSb2umzjMulhbA0+ohXvOxI5f/b45PUYeLXQfoeWJnkGl7AIiT++u0ppC7YUq3kX
0o+lO1E3GDVD/R1GA46i+Yzfa2wx+oagQzQNo2Z0y3falvIM9n1PtWOOyvzRAfdIn6GBmRnl+9vK
xErHEYvHQFvIzYu/E8QUa2RsVk1DntDd0K3eg6Fq3BA1cgWQt4XxzWnx2cmlot5Uqs1PolhRnuUO
pogFYDBoWnUEtP9wR8URhuB1SsIdRs4JbXA3MTAy/1ZO7k6tq/LLfMugv686teKLJ2yzurvTOt1p
emY5Dhv0KDyK8lDIto5v8ESzty3aKUTDzW2mzztK2YEu/NCCeZjs2srqiQgWSvSWnF9Ye5H6IlfT
imXHb9RGq9g5siQywrz9OkZhGiX9XtiFCdItg2LhTOYRfu7hVcaCFSIaigWX3SCgSlBM3kh0xQuf
dnwTRxZrbl01G8eB+FZuh9yT2rC6USLprA4wZzuQj/2I2Saa0Hi5PuyiWeFExwYcFvQW5pQRHDw8
br5wdroBVC8GO33KHA2jqTJhe9f0GUkbJwZ8RJkGnjwYi3+82Y6tWqYK4pbY0RpGW/fz6m5phAc4
2CQI57IakY1E/D1jR0EGWf8ffeJuE+FOVt3iqxFj9CLiXE9v4sfYrypO15X5tSumt3HWxBTG5xuv
SimFt1lRVpvMAwIIEMef3/gq8kzC788lif8M/34HRqh+Xk1qHN8P38bcHmhUUAypLWIQvcQzeMbS
0SiHE8aWPZcV6N3oSZ/5TcnACdacFPIjrtENUW2VFAcCmNN+QDS1sIgbGI1LO27ZUqUFq+HXsrpV
o+KOE08eFLoTzWXEwqJ4Snlp0Vd74lZn24jxKzXHUMIU4IYULtNpQktTNf7Wa3Cd/E6eX+TfwT0k
DhmHeohe80vjjf7/T0GnbZ2yh2JbheOzfyilmpbqODPeUFMrD53+AHQYR3cX/A4aqz9txVDBCZQR
2ExClot1C7U5HJLQ7YJeJ9rfee6SjVj65LXVrRSVl0VNkNkG0JbhTl/6BTl6AL0Mcj29h2ajPCAC
giDLUnDuwZWMTljQuOGewXj5X5gospRSMRLARQeFr0Prx0Pjfctdr1HgtU1vAIv6+d/gLE/U9wEW
NiYrTuxS8FYWXl7Lq22WCSCCbgP2+wea/7dRCxk/K7U1I0WL+jYsp+eJH9ljmPEdltTjacpgeDqj
7YqloqQWD8s2y6Wutp+Tfiba3tJTzQhSeqp8zwRmNWhdTMJGUR6S5NtJrCobI7MXVUBpIZHEn0pK
VeMtcyfwDsWx8WS9q8uf86ZzTpOHx2Jo2H8qFzbQuPyGvnBIo7Vgkm4C0wTBA/XP6yqH2inF5SWy
oJ4K2uFvr8MEy1ebTns/A6wwjJutnpOqXdPQUPdNvYPCyh9eMKpaN74ilmtJvaCNWm2EkePNhQI8
/VTARVSHRIYF3IVNdchFlrwAUVcDXIe3E8FkVPu92arZizUik40+16xXtAM0o9AmdCHTpkh5uGeZ
vc+3bX1MsF7vNQCfDgiM9jHRbDwqQ9L2uWKHZPOb9mmsKe0rntD2nAV+A0PWlU55YUFUufU67UXd
SIhdGz5ZbOu37kbNLhYFPRlAn5U1te8OmHq/ZWrnirNj6p/lxo0UducTymUOZeqoGP6/w+zNmWNm
kCUQ5SVgJ52Abr9ngFxwclVQ2ZfSoy/5dxb74mR+FpL40MV19Y1g637N0tq742JpGKIPgr7+9Mcl
my8bwJE1pbBfK3myiB+yu5JZb1rjdhHgUm4AlK+k+DbF1KuhY+G+qi0ewr6WlT9ifBvmY8QPk5m9
c3QWGkiM83SHFdnxGPUk8kQE7cAOKGlWU+l8Euls/6iffspWqQ8b7FTydp6kUnBDIj7WAfbm2hze
aZZrPa2fJ29/H4lP2z72YLgR+gqjLRrTvI9BwMKX9CUelueoXbcVxF9yvv3+q3wgNseoCr1wrTgs
lMEZr1s9z7HZO/jSIgPEZ3L+4c8em5/T8J8UElJ02IF/0i9cfN5RKkeEQjRfZYXzw13C5g+k2nAi
un+qGcYo1empSCwlZQfZ6h9/UZokh7vQpZhnIeENf3i6aW5qtwf9+hz4yYf4rxJMpv2ywu4YZ1Dl
IGpAn+OYafdPA4KLczlKA/AmyQwvbSAouVQGpd1P/bdCVOSRrqQtIeFWxPauGchnAEsmWz1oTzCv
G0GW9mretHMAFMwKjZBIKKg1vaNZCHleRYLob45X3CkEaatvigyKpEtF9AUpW+0IqJK/Auc5pwB1
mE0QtGIhTfByyN2LRzHA4OzJw5Bsrwfdg6FUuTEaHe/KEX3DVZnVk/qKmqUbcE/ivxit6oUjmzE2
ew3knL/YlD3QqUekC4+mJ1KGCJsiZhMymqeXNJDpSOngqfZSkM7CWFcsMM7N8bkLvZQt/MgaGZ4r
z93sZzoeECv2DlFZ+TPnC85TTGffKa1F5CDyPlraWtlu54qkm7dO4dwoxhxqp6yJIiWMBDzWdmkD
omd0ZS9cwv0Y5Qc6VC5HhVlZRTdwzKsYkDKVIveuoQRXNkspVsVRvrniv9cumBPFfL8u/0cKnN3P
JlRKo8LZ7x9yA9bfApzhb7AMd77B2ugQ3nVSJF1NU0d1GfQoL1aitw6cY9wxHoCwYRpb0j6oPKB2
r0M0Ka/IRzYB91Gjp5xRQk12kRgrpQWJvXbah5/4mHUkDrbCdyPuniaeNFmwebJAKEvLNweM2ypF
qHdMswSFYKBJ04ibaYi2IIZ4h5JkWperVlezV/wMIClAr7w5Q9tO7Yq2xdMFAHGI9RC3O0BAUAT9
qWbQunLhwFBTKEQIi2Bb2C5RXFR8iAgndP91VFcFYqTh7Urv2bGtCYjjQ6FSsp4SeBnW63EmzKx/
jZqmXZdKdIsqSdHqpXhcS453AeDRda4qaNDz0FBFY7VzG5ObTPdE5Pro7UOrUeWes1lWZSmz54Wr
f1msaMvz3Nn71G/xqro4uEGRT0We89dbg3ZhsIlvvy6I4JNPbr4CjZghnRT+C2hg6lvfDs+NuPRH
UbXB8QhRReCXWJnBHcCoFbpOmM2vUnb9XMWiIW6BJwcMAe+REZPO7DTQCsWKA3/FBAtbhlcXuYeV
Sr7RFfTdwIkUvDdXReVrsfy3AlifkJIzTPzToPh/KLTG4tqqI4ZMBIcbZQU6UfWnzsmo+/FPr1zJ
VnPcQU7+MMxMms+tOgTW+70aQsip4ZymTYy/oOVIJlXlfui7QK/f9/bQuBTI6W31hDahvAIDJ8VD
y4Te+HBZjZvkmFm9lHnvfWu+i3Vl51qZSRVp5WQYfnCxhiuXFYq2W2gGvIq+cno6tcWn6pFosfFh
Ofa4kClfGE31206cQ+CeGBiXGivgzqH2hpeXx4Rd/NVtwOnoAAYa9IvF+M5vM7bV0ZIc6E0pN+VC
A8dMxQwjcdQi4oka1sI1zciaoog/4x1ymK7VXsH/7Oot8Oa3HW5D0VqtRn874QlZWsp1MFl8El7M
FnEpQ+QkhnIGQ/hzxIHyoHgKps7ZMIzDqJEi66vZOlLtI/rRklMjakTzZy+Vg056jYte/WQfesuU
Pk/uxD/DUPWDdVjj2ahKs2a0tfJwbiXE42aQqd4s5+seK1SM7OLskurOR7kKz2I+3iiEb14Vc5II
HAgyA37+jcEt2QvyP6pOLb8BO2O5al7JBImu+IXiMhaAd3hyO/H2d6G8FbBAgNmXN0Xq6er4Th7g
zXjfzHzV8zhBeRVsf187xZyvkK1GaC9nk6ZQLZWZk808kGSViJuivhsxlXVVmYoooyqv5kTbgU+z
w6umGEXPKI1CQ5WFuNLcPK+n7EN5qDb1sDlFV9bJF8yNZjPY2cIVl8SjX/JZ25Cp/XhxY34F5ERT
dAKLWTMbGb1oSZF6eD8I8+u4PV2qGidiPsNYpnwTAcqmNa/8c0JyWD3MBEBVp+JHnjca33JJ5kMN
zTOzg4567dNi4N9bOqcjMGancvM16ioaR2xb8Kv5GnSAd9KLUPd1OK7tAHk5vJJfTAIbIiTQQzf1
OmnVwDQT0Jtg6JbrzrJ2PDMgIaHWZtCwYupXayvWpYt/IBP8/Zdp8IwxFKsRzkS5dfOnqIHIfQ0P
MVWyx4OskCnfBriNAx57p2sIgl05skijtR8a8WZQQyOwwwj2gYmqQ1Ie/lykDHs93B68MaKYUn86
1wIWwFQuo3QGXIeG+j+R3O6R8J+ZQv3H8kZ3pPEW4FB2j7O3WYOs+4X/IzSYe15kvrOWXiu+aDms
k2tyYAE6L+WKXobDTQKXDnveBgKoISDQ9s0fm6MctEUq9Ih1pixMpmQu3NfS8JbWZs9CZfIt9P8l
ojasqT+IY7FuvzWmYt8jAR/WgLs9R+234u8wR9tDHboAoey1nqXGVBuLhWYlL6cXYzaPNtqsgLxv
YIH+7Gyzc5Ldy8uEhcOoDHb+DM+cEKoqCpNKoqRqxqUGlgbU9K7A7DBTQgfY93z5o+ME9/18jbea
BQi6KIpUTZ8PftTG9NhidsWAoeTzzpJXDp7gPav82odp2O8OqCtK019BoPlM9mPFwDiXZr5q0GnN
VirhNY8aCyuA3AzBgue1IHRL9th6Niz5UN/m7SPkrsEClbvQ4c9nbAUv9tRJeWdsW6QtdXs6Hp3y
erLzalpZK6p/OxaeZaIuE7FzHGkbyOWbkwWiDJ1tdcRyB/45H8DYJD92ZhKQ2JFQ4Pj4kBoDjW21
/6je6AU71QKHF+D5E2IXG4M292FS94uqK/L+AT0lqIhTV3PaZ9XjJSTce3SqcZPo1g0jdgycPEp4
tdxM0c3v25VQpdQnE1LiPLpKaYP8qgX+sRfIze2c73IjjQmehAmd67miwWwwBtvJI4yAdQUKZAe/
LEttZNXZshfOy2Qvke/EYwSF0L4nFnzS0tK1STfL0WxYP8p+FsElhQXc90jH0tZMApIP+wmYN0wQ
cEBJE3dPD7+LHwlx6VY5zZEbTdPT0yJoeHWEUSdBwEfhWz59WT4mDfgLzsSz8B4vmr//vZarq70F
bzqEzrcjK3nZHjMed3VqXUFaNT+Iq+7dAWzAuOotL6kD07dOGr1bNo86wJpsK7FyYt7chGFFwZka
7ZwfVPs5huY+8v9gdRlg0vqGOKLSzjF3qpP3zUhXiCgmp8D33FxVqQhcvhtVhNk3/7ozMCq7i6qO
vQZ+Kii9mFREP5xNPSiy63TLBFvEPLqybJS/wzcSYSnz2Xez+/i2IILbAR9Yu2EOMB1MBiqh0Jtg
OqVSMGrRC04DQouepuCFdxb/mKLdQ0MVvzP8ibtFIff4/MqYsQo+XSGzct5hQMjs4leHWo1Dvom7
8f+tJrT8rvQ5wDxuCD897Q/SScrlWcHLmuEk00qlKdGfZjjzWxx5srRkygndWAM2upbMVcultzIL
LbhHkLs3HDjdTcw066D6P04Orr2knC2N6Xgjv6C/IYGoZYF/wI28ANgFNbpkd0lIZL55tI65BGyM
vLAl3VsX/XrpAmeqTWwSkqRNzAATJjOgb57x6q3JduxC9u/YZaP/ikkGSTvF7enL9goLn/nJrrPv
k1r0oeGibkt5kAncKn4TYBqNB1/TAsA30DIK+pedGP0/azMIFCYcK2FAOi2e7PpIeZ8U+uiD1roE
gm52Qm6h8Twte8mZ7m/4eS/KSfIdhGCHgs5H77NuKCNCdqIv3Mtj57xrZ8rHZQPUUKbR2iMxrFtZ
txzKHVuP0jLoRTx9F/ABDN2QsThcUuHwIwI+esp6Jzt47GTJYy8zCt6rCm+ZGD61MnQgMFDREVgu
JmNnpyaBzpN/iWEWGTO9cKRA0VSQ3KxOUKlyLZni9QOiNJyUuJHjK2hVoKbMyr0QeSMdK9CZ/1Qm
lQ0SZZpxFEwwb42ptqAnx1Apmm4EpFIkQMkNAy+RxTvFhQHmKY9yq601zaJtRICSGr7rGxiVQhOg
d4BTNv+zZYPi/0o0hVk2DwWuZWg7E0eIFK8DOPdUez770lDAcq63eEhTMboheApn/PioBh3qML6R
9uQs1ya4wxJKX8gDR+kVqhSkLLJBDucmgBsYSc3311AlMZy2FgDOHc0OHkR/GJFckp2DhEb5ZH2b
8jLPlOUIAWIHlyRRfbiH9F838MbcPejKWWwmarL8Wmq1+JSJ6IhacwaxrAFMCNTvrbuoPQ1oX9ra
z3lQr7omXdIdtfyB+J/AW204L2Z/S6X4Ax9bhIN2wrHOyycQwEdImorq/cUkyKuyiLhzC05AMVFJ
hocrWEYCG7dTTJxR2s8xLxGg41yrgzwHxR/qSENvIYuTD0kNN7vLcZrLxvkEebYVrdC0ga43cZB5
4bb5IEOyDTusu9ginBsBOMgCXHhmlIjr9rZx4Y8jFx+HqeH1Cfga7eaRIfFUGMnoG36QKbwTT1Ek
dOSfYNjLe0KcRJ1dqxFc/zX+yAtxdKDLSpit9tfutznIRMoRS5ExcgDHZl2eaxXBxasUuV+xAeD/
18KFrb/7j8ZC3FelKfebCf8/vEGO2R5n5m3qfbgs0bAGXhF6RkqvYEmxxvNUPklAR+2m13fIhuk7
IuLfy+7kFpXxVFEojziGhqmXdbWu027E2HbLRXxuwbVcbd6sSejAqrj32kOHAjjbjWYMulgNuNjk
pGuWbWWWNCuf7eJcr5iLIeyNOp0PgyrphXJGeg/FZ8cThs/m4tWsVeExtIBO2wv2O3AjChPbK3SR
9FYV14HiMiwMSR/AAYMHj/SCCByfe3ZgVHM1pfBAYTqFWv6BS7nq5i77arxMyzhQ8JZPQyJCB2Gc
22iqKt50YY5zgMNpIjgnyqG82Vok1kp9m7hVEzNP2mErdRYhTOYjtDqTZs+GDtH85yqvS+b7NSxp
hK8NDQvIXBUzYkTGxjldKclma7j21/7gKupB9owZogR6kACXL9pokkxoK9lPWy6WArQidRTwNXIO
ukrWWVhMeeY4xWsxkkoQpXTRgc0H+eummrEDM+oFP1XroeSLSIv4YYonv4xlNZnFY2q4r8Li5MbK
Q758HTmJcj9FMP24LfSC/kL9ApdicXvI1eVJPbFkVHJJzOTSvWkia845FAJc0xP37lP+4ALjTeFq
wyL8hyfO6ivie8dR3r/WBHj7tDfaEbmIr/5hx+2YkIFnPPsKgsMA+ih8sbKlfGDueRgEx71/suyO
c8eBgUbC99kEVxtGuGNKs9rv9dRO+j63p/8nINwjcJC+beGFPEraJNe5exUA5kht5ljciQTRJmdp
RhSGX7ZkADNsRcZx5Hf6KJXsIDe93TL2xrmgssfXfR7WNeYZm+0jm6hn3Gsbl0nh0dtlJGNMmMHi
5Na8S0Y87XSrqW/Why/3R891udJntJEWKbQV0cMp5sI/PvHe7QlvpEmiyG4Sf4/YmVZZr3LvAXb/
SeoCYwlcWQMW8S1axvbm5RtwpEBixoso5IsKGofJwrPVfNMmqH3Js2xR72yBtOophwzTEKofyURG
Z+T4/jUBm5mSbSumxbd4VtQPGbU3gaVBLypaprmPqOeOMMX+OlXXOGx/hG/SSY2EOs3+aDufSGf6
u5WAoqq9D2+F4Q70Ub/ddzXpJL3y6YZ9SNGswKzU14TLezTrkV/Qn+wWt2cG10QN7DfwUQvhOjHG
IVZa+Dj5fgMbLB3jscsnLlD7y4nwGCHxh6u425z/alQBpRjNgDO5GC1A6T+agLtsQi2d4qM86hX5
gIsMu205nzcIxNxcC0odpY5xV+74moDVcdt5YfL7aD0haKSvcNSqrpx5M94ndFE4S5rIHGzj4xkn
170tRG0vLz2aCaZU7TDP+5bqj3znxhCPO3HQesU50vhh6A/JZCrHgmjgZdhVAfbt8sxB0FUvXoPR
HcVoXYXVu/kUlgOwhRr/rbCBI4jXrqUw9whCyVglf8wN0kR2GTwf2Cca7W7aGrQIDQpL3WxYbTbn
gmWQCOrAdTavm5RTxwd9/v2PKpfWMo6m9kDxyrPiqFTaKD9eYYhFDN0QEx0BKp9JSIJLhSbGRiyi
VXUUuG9Ede1RiDSrGkOZZTj8awdzQSts4Kwhu01H8VHOkLSFzZQT14E2NnMcqfkCScRTuNS5ZEAn
fstcPXgwJsevEFo6nAVLUJ8Pg00Y9pZljkW8RAn24PS0JQ5o1zyuvd6XI5ZrNHhj8gxHOjltIPfk
rJNuoEJfQYurdAEmj9RgxhkA2LpFaNjJiC7fsI+thw4edPGivT4AZFBodXB6sB3VGxGINKe+DG6V
Qw6k8OCCUcJ1mIO7aKezXXdDgqrsupQlPiD+FpbsZX4kydfJKmOMcRAABcOseM7m9t7pyEnYsPis
r47nsupxOzMkMqtAT/dEhNrsaJQqJzGbVLqpeirNQIcR4msOCDt45apzQ6k6obL8Va5oFLTsY9O7
lsVFu6njngo7L4kLlyW6DMpPELVh2DS2J1/7UMs5mp4AFN2BtK9o6FH/Bnulj6+iuz+ITaeRlEKw
TTdMCaEDcHImYviWPcNvLAsIu63d1RmOHWmNCADChBp8ejTnwhSLGlfs+fiGP3dbBDBjRNwgYCvs
zGtIxJjkDDmWD8MLiPF6wHxC0RxtOSxT9D7FBH3imwX2Ma8DidT9OhcbP0ZDVgCZaWVkgCh+2o0r
0JH5rx95QOuTq/eGV9aZzc291e83G6wNmYds2lKJbvkbCKbkgeTU9phA92eFzPP6vtF1taEIH/MH
uu5kz1HJCKcQIyLvbOnZCEuyOTuqs3ratdg0/PD3VrOkYpo6Jbw3fFqpkKCadq8zN5W1Vt3qbOor
ew+ucP9dB6oqh/8TKDl9JYjZQuPz6rholYbDgRWBZ0yWKlZtQcUf7pJnRBVdPt4GRAjD7lPl3fJ9
no9fDWX8zd/sAbGReFXZzGQaQMh0sb+e8c2Jzj7SA6Wjn4rYpx4Be5eK83YRl5RcOQYkxjaOzZxT
kGjkOs1uoVAo3oJn51NPO7KsjnQA1n+N2m8EBjt+bwBfhjQCt0s3+WrJGe7QlInf6MKFkZ2czhFt
QIQUriMGnQxyzsMe+lgyxvNWF8l7+oRoRTIiamceaCPf1hZP0O1nefd/AItRRg4ASg+QtFgtZ7VP
m/wuMcN5zEs6cidFqU1Q5S5XUC7xFdfXne4wEfM6Pkbd2V2GvS6kFGOGEULWw/q71XKKsL62RXln
SSjGpFvlUMRo81uvgijncBkn36Baus4hPaErYKzrwZGOxfE9KgutcpMvgqzij/KJrosTzUdCajT1
4JscTbi9TZyZYIRVjepDyB6/uI9UArRizhQvn4FeE2Rr9NvJK8/gLl27lkKe+z8igOH1jksWBsVo
TGkSBAy2LVWhiGp6zitOV3kshnpMsoSFk5eFyB0P7AFPZpWFxOzQ1uyScp8KABW95+P+XPBppgot
QWiqPVjETTy1O5HmmxwTOC3CvuZiLOYB+sXzD0WGohYA5U4/eU/m43HkOmMpH5xgylnMb3jz3QfG
8QcGRgz7l1Kq12ZBYPWNBFS0UhrcoOyjzL0uK6DOG0AhMP4OGiYFPxOWYVcT1/gefyOoyr7a+TKI
Po7yqoaxyUDDmMq4SEj7yZtL+wg4mZiAzJeyba+4EAdn9BzHkUzlJMvYqsdMv15MxwJFuvHldVRO
meQIdkdfPfjo9ts2ay9hfArO2UECZvG51xw223fnCnoAZicCMzRKKKLv+kPW6Pr7DRB2ojNjJHmB
iMcT4kOGfPB+p6S/Ru1eN+xEDkKe0v26V/fDPAtemb8h8dLmf3fgb47RG6jqCIqE++etyNPreg6q
dCutETg9Q05G9LPFuA96xQvzRXJCiOwsJuj+KtSCnXGz+yjZ+PjHuBWqhBATqtzY7nNuziEDI1pi
eyAuGRHQHcRPRGsoLW+NLLV/CFSFrIIlO3pLk1KpEEVDSJmuHqlrsGc8/KUQkBWXancN798UP+zc
AW6VoJa4okxpYabOL76nj1FYSKyfYSfMkIlK1tq39GkyO5Qlr9XyVROPFspNWL0kkBLsIP1XZk39
YfNXw2aEdVBsdqt9xSpJBvW7vAjThr6prZFoH8kovyLkW48y9qTwinXa9/6HVGOkdKv+tMkAKeuv
KsiLPbhE22uI3CFu6720IWDHT9HOaHY1c7/m53xIDPqDQ1ec5G8KuQ1VyvjYz9lb8YF1Q7H/KeIq
PEvMwFNiiG7unBQApOOFVi0ROo06b7T5UyeOh6aAtYVQsju/GaWK14hBXJaqbR9JyT0J0tzPDeMb
ffHaimV95hDEDoFgYYhzzeACAYBN92kUIX6tDkFbspxjIDt3x5YXNwYNa9BHDg8AbViPibnQJ53j
uFR9GXTzNCLO8NPvHrzni8LnaX2Wh6oWQ+Bf4Xttg0P6/YZMcRY4gQU82w51iNUbAsJszlz66hcH
ipc4MyZyQM+BwzwyeCdwKRfxQ9ywOaZjeAkzqKqu4T3BkSAe9Pa0JnE5wUTHClg/oPHUtAzxYHD1
cahcCm69ACHIPU8AVO8hNxtgzftOz5MFiMr8Qa3fWG5pq7pNlqp6hseXT1qA3L5Wq/CCcLRzpsWU
a7Uyh4IlNxURy5V023OADC7Tm2DpszYbRf0IY6BWyZUg4c/9Sl5yTraSrTfmG3mFukZKli1t7HOU
djDX/MY+Cz8VKFFOdG9aqwR7DO4tR/pe0NKupEDV6a2l+3IIM7r+QXkncSt1OA1ZjMFFYZO9yW97
BTjVlepykHgo+GRLy0QXqzkVLX0pyZGIG1ewnVDRJ+6SbqUrSl2YMBlYmqZoPiDuoo4iaG+1V2us
wI9nGMGunv3IQjxSLpr6t+XhhCSk572QHsO6qxv5fzit9BkwnIBeVnglNy7xyy6rBwWgxsRMTiXw
05/O34aFqoiVxl3tHDQjdoGRSfpjNI30832aGC1pAHqThS9wbkNwN3Cx+UoGkjjde4JF6lH8vSdt
KRl7AEugfwny/qdn7GTnSAfB9zIV3oiju+R9UYkHkvU71+ns/vzBHfbiBcZSMFs7yKB2Bm5UnMjj
GcLG2Kket11gESI0ZbW+R0pDfGyrbO0YU4+tEBil/bDRLMYKAuenSTQu+Ubw0HvYoI8YaTWifhHK
5kjAKydcnZnWn4dX9vDP9xmRB3wgRQvw0Xax54j4k+UbHtGgqKZfjXXk7OW6pfngNLBN6c4cXRVi
hHRxYCfvLkOG6fWdtz6kcpR9EWNCpRk8g9NzQkaHrUIDYodrkNNTlHQmz+kDFJ7k8bgqQTlljLZI
YsApVj4weUOuVuQsx0V9hGqFaooWixhRCjdnJfNZo6O3RleUUrgmZXnkr1cOKK58chnXU0gKX/D5
1xzkMk2hYoobCGYAUevC2Kzs7HKTLsE4c0FqYq8HlaLzdoSzo90UDqZ/s2ujIRnuWEgrxKgSRhsC
U0qqf9kweTkiia0/2AV0WCB/zYKQisQibIcAxO7BxTybBXoInCcr0YlljDQOg7osG/Hsl7jBb9O8
5kMdCf6RBn+Hy0utVgSJysqzyG41XMUJA6/jgkI7UBm3blvFGEN2TP4wFolegwjuba4BgUputGJb
JCg1ajsYKcgUsOwOvgIcPkio0iBKBWTifYjkzdf0PjEcOwNeTr0Vq+ENqdmkPaOSizbyEYc4vFZW
YL8QP4MLCKUzMK8HpqL2XbnK5u7cVwPkSJ3E1PopsgvoMawLmXO4LRsh4kukHFHTQ3bQKyloshs9
DDngeNbVIe/KOs1c51z0uHmNBmLHTINs0pX+FjkMgC41x4cRBj2S9jutSi2NA2WvOknQLPyHyEMl
3GOgXeIwNkz5HdaSXymHLfPXkKVm6qnTPqRZXiHEUX7n0JMMiclzcA2Mq0nBn7d6ADuK3VmjuK6i
MTtYK/CZNtKl4Suz7S2NMCBUZYmIwoC34JYm1D5pWegMvcXT3SJU9co74jx2DVItD6Nm3DovioMX
IzNh6/sr7igw+1VNHD4GvNOXd3JRrWl8qQDEiE2ZUpK2x4WLyLdw8wLCiRiH0Ta7+wYYCdiAWLWU
plBqhAvWNnXC5lbvpC9zQxuOqYugRvOVe3+vnSrt9DowBABby3VlFXSy8uGR/yAowham0woLmR7q
O+gAIwwRcjIA4Irmn0m6kMR91CIiFWnl/K8+TVQI4wUNePHRHTxb/LuAW85o81PrbDQPfvr9iMO+
aXMLgl7AxCtXobddsjgPMd4d3fL29S1DWEvpwjIZpdZ4/EFg7MSQnhBu/2s1Uu6VGxA7sIO0hErq
q83xVW66n7f6pGElcEa/ySKo9Bu5AS3TzRGXKagd99VRpZfJelphzkdyxr2mI+uTmSW1EbR2AzG3
+mOdD8DWpWN6jLQ+QkWV4aPzsFps7s2c4JzWGaeJCDGqGm2wU7rQUjtYn+nvOCZcZXI9OvPniK3C
pY/uTWjYIdxOP2cAf7S2bB1OrWuSIPo8yUsFiHzK1tMJyJQOx5na2m02XgjVwYftqPmtzS55F7jg
e0rPkq8xTC0eHDYMeJSMPtmamwgrRJ6Ur2+GrDkWOI2p1T9LTz/XBKbsFo5aoUU4Ur7xsQscF9N+
cKzTRvExw7jEA5bW/dHSAXgU1MVJ/PVICa5McnNwf+1TiBShfaXSn7eGzVQ6A+FS5lH3LJJXVUTq
2Bp68xmHRzzFxxZxY5p7JghmruxxJxDHFN3LqQ3PtWrsEHKoBPeDpoAPQ6M+iFMV5F3z4S4YxhTO
hnSoo8U234psYJiFhbUv7we9GRlHSCCEAMfO/incFqMPmcHUBNzrk85WMoEc0r09KFqoh1ZSn1po
otVpPGzQ4pLjxIFVHZKget6WSDFNmE4jSbyB8xGY5VC8vCUNpPMgkhToVBum+HA49aTFnLuER5N+
fzmg5p85oO8STKKpY9mmIdbObzzlxYVnc6+eEVNHDfDe+qt+QJzHCLIZZdWSrmcb7mfbPa9SInc4
2fTC63BHYrZh/b7Ng3RUDPJU5U/xUiOD1cRZz0k/XZxzatoVrdDGjoxEcxhox8TNW7MxUh9ZAD26
5G16fzC0OpTLNQ+yQONVB+7u8b1m7I1/aTsf/L+MtQvoD+lzjZlY2DFMJot2mdmDjt7WpPaMngRE
lgUWy+ovuLdpX0xICdh/NVEATaSDRO6NAmimBWyj1un1dPkrV98WgxkCr7FS8+QkoMW5EJ2Vv/57
SwyKWnKMvQdbqT+Mn/SFn7gnxHZjXxHZGK5r1nIAvtWz+uH9vnNQK5GtceJLUuPNBmC3vtshfjx2
mHO65lLzjhzW/t1mLqHTYAJHom7ftB3P5yJK/+0biNzIh1mnibnWo57HOLJ9AzBr/mGQBHTJ6ZeQ
uc04z2N3k83suhGjVnSCubsIO4FtSy2AAk7sKenVKzJOkNMMRlxIcfOG10/svzkB5dOwVTrcgXGM
77oWUXKhmATsfowS3nNYUmsH9C6LSR8fGC3qB/2g3mma8wQl3S7HT4tRNx3JlDV3TtFN2obUkBih
kF8auMQ9pzK9+x9KFvngnNwRXbzSJ4F6AhwKxAOGbxBhd+9S0W+mNgwQbSQovzlvjbCdKRPLIL+B
LsFAJK2qNT6Z+Z0fOKQ4B3ZwyEdPl/s/gik3SqVa0zL5VuAbcP2ghmeuAyfdL/i+WPnw+UWfHmeZ
QauIlaMx3ZFkebuQNiEEwaXcHC/D2hh6XHQOtBuELGGGB5BooJNXT870LbfoBY0Vza9ED4E4BwWn
j56S6RT5lFCGoDy+LV78+k55YaSGkeW/EJL6Nl0Qjt4K9IoqyZX5DZyNX/SGgubpR2JqSbou26S+
LN+DEd7y0puPwieM5OBaAaJxprZZBrnS1kcIXp1HwBRYzfcmB6Q/CXppp0FGsf2iVAUdE2l7bqJb
uhnzlODjKfNEGEN7Eyt2ZTUOf46yNI6jMfWmpxmK/1t16zpNiQhamtFdPt8gdq0i2JxNlVLbDmLD
jJUvSb85ekLpqOmPrkcX6+fTEKVZCDYs9bu0TBDGiT9iKrdr5fPc3R1YY4k8iT4RuS2rxMFNp+mN
+iojqtbiTOWYJxYnJM3JAF42tBLPYry8EkS8Aqr9PpG2aySWvrun2g5LNB2TH++WOSHDp+FZX+Ym
C+gI4/bhUMoOAeKBDSRD//NNmTEVeYSXWh8pkhdoSl3UKQwMF1yaBh3Htv4Gtq2xHokRofJPnk57
sDOOBlFayQVs84on7w+ff1XnTO0/zzA9Cqm+hBjZ3QzLYq6l6ZrVMDl1EYLqdnujNdNwkuuCgh/0
Xn1PzJyXkmWog1tulVayZLhCox6oWQE09u4f9jkJBNOvTxqWJARWvfJV8e2Pn3tvIgOZqq2DItlo
OPqyq44V0qoY/uh2o3HN2M1QwFMhA30UkqvpMnirFJX2uvYpfrylzkdkD65mmPEd0xR6yqjuwQ31
V5VVqjQryj81IUy1Rq55bQoNs8JDCmgTpx9L9t+vXP+b8wvpS8ybko3sJqOX94gCrLI7mDSfuJYV
4LJhGeKntb2qZxLzrdpueiK7+abzOmFHRoCrmd9DLqwmzLTmT1vLhMdU88S8zjBl+Uf4Yei0Hapj
mCHgVI9c8N3BlfzQYx77OXNF7Te9CvbADBaYzSqVEYeFr1XWQrWiEr+9fnQZ/ZaeWWNUYXoYhiVT
y5Yg5sjQjGB/66hrUDZ7E7AjmuVa
`protect end_protected
