-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
mzQoLFWXvRhyVzOUmwPJ808dYcbMXHfYrPHxVl4Th53N55HJ5jlLeHEYHO+2GonS
4rFE3qw5wKp42hrImhgslU7FFnfVoBrdua6I4qLEzJK/pmUiXN6DHhcZ2UTwRGpm
fcjaFl8pRllVq04CDi4KTY1m78WA/3dKxeIJrm1CvLk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10336)
`protect data_block
5Hzaxbe4mvXSeEYZXAf3Y9KzyrYMEWzkToqI2XAMjaxknrVYVcPOC72ahc9dcRhF
1s9y9vJIQk1v45rhxI6LxyJ7OxKDyaSyhmcRp3uECWWxoSm9sBuaVxLAEo7gapff
tgNUUaZrzrlfb5PgY2tpyO1Aw9M+TTlfZAlcpumWWSonlBM6jtP/IhnlJmuL1G1q
UiamWzcPYJwyWE3Zg4T5XS5kzFECLkbikGHaTdtg8qGxXZhqvGvVyQ/89V3FBTqR
HdiTCqNJggtrLcYFCOA6hb5jnBNWRKizT0qMyuGkWHuO9IWE2EX3BPuqUf/NDEFy
2M7zqX0tIjioUQrVvTPHvA/LbpE2fAC5TfR9Dpl4zZKPb/UQdxuGrsoBg2niIV7P
xPcu6LxtiCLHy94EWB+2HK0wRNWKGHUAnKXC+qveuHW+DM+dpNHQFWY9+8WGGM4U
dhkLms8JS9oC4Mrgj1Y2w/2Fz/YjwLILYwyldmHfJwmPogULlfZqh8GIFfJ3r6Bc
C5uRucxoDk5qIKd6ac2XO/ur/hCWGyT1IPS61MnS3HI2H6Pgh2AmjXgPeXJY3vgr
oWxX+ZSJkDRqVN3y/8O+t4VzJwAalBi39uAsJY9FnpZFV38qZMk3mFbUhHQPSwqu
V/tCUbOBZpPrNawBk6BwIoR9KH9V04VjaJDyoK95NyMIK1Dncm8rBbZ/OQEhAcXC
Ri8PLTfSBd+k3qjLXaMYQg+5Z4e3mWO5FtjS4PB1iLzSaf79imQC23ElzpfqU2y6
/dVESj9jURbjrT6JSket9Nf/ydywFaUNjTtTbkkDESlruyOHtssdoY/tbqbKlZaS
Py3lXuOQ9MRQ6aWKB5wEDb2DLHlz6RaDZ5AWwCkcmZl5Qggc/BfCU6OWuf5QIj8r
dzscbE1G02y76SKz9bUV78UcOctnkAKN4Ryj2gS0sRzmK30BgxENwk3wOpRX4690
YVhtmeOtUAjKHiOJBlfYHLtJ7rFckJDKrLkbVQmtMQXVlmkraVV1ChT90poQ//VA
8E4aj3nYLZjDS9pVzjz+y2N63KewnqMuv4hi0BOzMJYuLzHCLEmB9v+SB7o7aS0j
i3FJYEdbR2Vu70eEMtmRQVUrPspX4lVMi1JoDBKc5kJ/2Ayx3vkENzljA9bG4NON
jTg12iy36tsI8Je2RIm363IMAnjf9a/OzvVu5ZCJTfPB5ryKJDHBwG+7mvDEW8oc
j+QpmPZSRr75aswCVDeLTVeBxX3xZC6W45+88E3GC1k75Mg8n5grBj9AswGgyYBk
H4iPxoVU2NWKMoM9AseeYXVJ7u9MutiYrZ9zQ4OlIEUM7SXb/Nb2YbauLzXwcx5j
YFqPK7ebxUzRMsITFJwWV84eM5nxetsIGoKDmSIgxAhlfIcJFP2+FGGF+PDWJeaR
XKbAwLLTz0L5Vmg4TNc3oov78/oSQazte6VlDeu0AajHDVgTa6upI7Dti0fTWAPI
3xuumlQi+Rb4M6U/QlEKbHCoN0i3UJR9ehXCHcxaegDCPgeTLtcbL+lzPOawDlg0
d+JvSzbguQMpX8w4Ph4FSoTFJfKN3Ynxq8yJo9J7jA0zffwf1rJ97Lt1Jd8nKDca
+4SVUk9xhrYVwZ8e8DKhIEK+8zZvBHdvPGp64ZSLjj3bcOzUXZaK2kJG7xJLNFH1
hmZCu7FG0NgV1REzZkjEMx8+cIazrRkkKkIjCuFOJHAvNrQ47fZ5jB6FPLS4vOnk
a8gm5hkeI8js7t8OxPi1hguGhwT+CmzNTyPwJ0sbNWr61+9D4ZwmZy8ZpbKcAE8X
ASOZWZS7Ojv5WlAwEU7+e/HUWGnmwLVHd4nHDgRNiCScTNQJgCqsOrsApkIwxVEh
gXjPrAY0A/DlEi5Mw3MXGt/9UuRp5KZZyYZgKO2bUoINuzRs3KrqyYLHnU0sjx6j
/7Z3yZpkHuEHEm+iYXl+00k/CcESZmm4JybV0ewk4gOQAzpB3yMFVhSg9f+gBRpI
U7GLDO85yB9W2wivw+AqkKjjutgILUxQLQyVNpb91VU1wNaTm3WP/toHQcjVd+7V
5gittvig4OBw5AnIirCZmSBf2P5HR+atUUp8hm7npHzQbzRbUW/Vd32J0/4mx07Z
k8BknCNCZ3dvvJfFUSwuj7OoLqSMe7wWZIqqrUDBJXLSEHkYWbBgCA8hPziFR/Pk
I5Q2jfCUL5j68sHjVvZtDik+/g+1lAHlD5y+QJYOGsv6E8rZNkYbohhbvWjrBWt8
rAMqY3tFW6yis7kPfCuyfzpIp/bnqU7k0m3hthHsK/8Sj25Jlm8PV/Fu5Vgfws/p
nPayhBcXPWOUumXx1+IkUIOnJ9/VWAwWXh0c5ue25aIe8UIn08sHmEn7npRb0p7J
ylNUC5nmIqj/M70Yec4viVLjwab+B5QYnp2R42MA4hIqVpmt0kgSm2N5kxISJwQQ
38NPFRmHPLX1JQPB1LJi/+vQovac19Nhldwof/BuoVjt9Rv3/wc/q4tiL/bzMBpt
sc6i036gfK4+7ma0+DiJe0sMpJJ1B4J2xFroEdeEiEHTdNqh0ZQ4Mp9DqRIQXyfg
8lIT5XjyVNEko/T8plCkvQSn2JMCC+/uJwu5gp0JRSCT1p/W6muUiH+LvE7LrVcF
uccITxe8BGPdbmcbHjVAPsWagwL//Kiq0yMC/yzEp+7cZC8ioaxmqbR+V9uDg/cC
pK+TY5LPk/oJqfBabM/MwO2YQFAQGi7TWOpydpMv3jaxtn5IJJlv07NHOj2liuML
1d4sz7A5u68EQGHfeAgk5JP5XvpsTE6TMWC6fstyCAcBaDl9G79d17gCHk3t7QY1
8s40y381qQfcIjOKHcpy2rKBv/7dfp/5jRw9zsNq3T2xtG08+TDXM6A/Kx3Rhi07
NnOFCOpRi+2NODRzeVez5hLrZ4VbKUXA3H7lbmctOs9RKPRGijOlB0kZuo5FFLSO
C6Wxst8noEm16B4lnMSTz2P3TcupxHE3pyVf7f/iSukH2TWp1y30IWuJ+doVWJFY
YdkdSOEMfzoQfzOf8u1nP99TQDYNK8SEfLZLWwZ00xkjORTN1Dr1mAt8f5FLYCmF
tV+p9w1/0gUY2p06j6UMlXkHjKV0dgYeziVHXk2ju+N/Yp3B4XipATQdMdCcpChY
7P+bHLVarBgl9I4p3IlzFDbf0po2LInePd3t2MYyrrqqtNsIkEbRfuCK6wki3y4a
9qKalYT8VoWyd5ScDueQ+IJ4octRrzw4aAQ4EfLF8a5bl0tnOaFka0WzyVAkePFu
+BjiXSOXDkLiI4gtJR/mdgC6cFvZyuTEi3SRgfmeQ5O053R8ePqORZuNnKXaO1kG
TtvzdrNeT8Li8CHF7V3qc3XwrGIffVGsO397hikpE7lUTE4Am9+yYDlJBlIAItIp
rOiy4JxkM3d79zbFEAjDmfBTulubwho4Gj7rRlGQod3vAzw5ffp1u3WhIQrxSGea
AAb+e9HPNuneBWJbZQd0Dp5hZ9CZ8lTpq4Enx5XhHF5Ie2a/3G0a05LE4wH/dBSB
5wwfHLF2bko5SVIkKxAh+hJzVXibAFx/Cdl2snBKtK3gd0hIOrJrVM4eK99+5z1L
FsXnnw4D8cYhYjv8XE+A93tzglQwCLeJ+7FQ39ojS8UdH7FyL92Pufi736qxjie1
4IvB/XOMf0fdLVQFk0NtJSWXQV9770LeBPcuuBicBzJRXJgKojT00wfFpIiqPhCw
auasPOGwjB90pptDgJS9baxzxHxRyzpaviyOeJGbu29GdA5qlKYz42hqTBSJpTVZ
Khq5rCPhlILRELk9r8adwHKSFHLpUJMoDTVykUrYYuy+LQ11Xb+3qXkmps66ioF0
l6lj0zXPynFsGmPbu3TFPqvf7G9E7SvsvFvr10Zq/CNxW06KhKUkiKNYEymzY5me
fLuM5LG4cf+WByOHbg28iTVn2tD12GB4KzNmDSq6rv2gL63rJUkjQnzwyihXz2lr
vIP8re2E7yjO+hBrOxHiHveGBoKex3jVk05Z+tD72IEUfnqpblS2quLuE+vQFzw9
MDBofeIpSZlO8hUvEpv4C7TGaquJ4x3THp7VsfRFwiOKloW7fUbiPhlBPbrGMn/q
487xKJvd0zlgDXO7ewBgs+RRhl9yFLTjJshc3D5sEPowEK4CnXiBO2o59KK6NwrP
5jBN6bbcvgTC4L4VL5aIPb9IqbuqU5b12+qyEnJouBjW9UdQbdWhnorRMA9GSTZA
Cg1epoSA2u+8tHKCQqde0/+zjyAzMrL+F6AjEBuNE/DaxOqOMZnybBKlbXG0v9z0
X324WF3Q83JDN0ijyHEGcW8dS8VLF3eNkFuSAfISYBwwkbjCeJRI7nqaGnWwpPPd
69qJc+I7K0Yqc6Yn1AVZvspvldH2wT/Nq1majud+lkV4OgaNkfHbZj+K1m00/47o
DEAIwWNl41jLVIw/won65CQK1Nx8ADPhLoekAzmNJBJ/SP/ch6bbS56L9yKRRj9r
hqLpMdTODLf3OlIjuXbzU6dJ6n9vYN7eAUDJtkyop1EXOIzkD7/SYJCKcOFTZgwk
FgFbklNL9syv21/uphPYQPn7FvkA5vXewg77jO+4sT+tMUmWORXBZ2SYu+eLtPQB
l/9o5DRYIp7UnYRoFiYYNSrNnIIMDaZOMKprVjPSB0EHEKQmBlSQAkjkvJgRjp4W
3vyTpd+R+PpKtDidYgeNMkWzlSuAr5vKWXow9sZ7fdrgbOmSgQ1vAWWEY5kjjEnR
0aF9P0zux9AZ8f57iftpGiIRjI0Vdnddat+O/wcWGVZwk1I5ygybhfGFebAzwIVt
P+oLOT5xu1PZM9ye8LBj3RVza2Q3ewHVLegVGg8WxrWZ8Zv69W1QCbnhUAUcqVvM
zJIgJ2zbidviz/rrBvaOY1JyMSPnkECfHojFtDY61rYy+WMxuJnSux3k6uurA53e
g9rmf5i+Fj0wDoS2MzAqJwFQF0MLzWG249ebRgaMi7Bu3GgTmtaTCDkz9WKz1KyV
GC0xnyghtO0QYYBXxq9byooKCA/HqgZFaxhlc07IOFZlXyfTb7b1+K5+qYYY2PTA
ODbzFOHVtiOt9uJ1ln1jL1PppnChQnxrjGUSc+HFqEpWrWkSFi+JMGVCWMbTYoNt
ZgLZrjPslxB9aFBTNf+HU6D/9rRkQq6/gDkjvjRSzfiK1Hki/Bo4EyWFY4jNuYFY
gnQ//48ddzo1bLkIYH9H+F9XX73PC55DVPS1Y0KYaawa4M3amTBRH/TUBHldDc1Z
9AWdbA2qUKoPrHDrVpR3Bmqd0FHl6CYgG1O9rcwrNRHF+yzkP+XOICg388COXZVT
QAtE13LrUZEav3N8Utt0YX+K60DhWbJN378kPgLun7Esu/svzz9O2iE/OEeji3bx
ZktgT4p3vj457jOWYsfKQwtFpjGgs+dEXkO8EtewypFPkIf/gScWZX9h4405CyKM
0KsmgEcsR9geBj/PkJU32rCbokjrvb6c5GkBRJM4LrBcdo2WVxQxVmg+iIpBao8Q
Mv9Qs1xjO46VyRa09naJVKuA+iDxTVdbKscGPUsGuaBiSYGUbAe80o0LYtVIRSj5
VIr4KOCVEglx7trvUx1AhJlAH6acLXb1PY7GvrPv7zlFH600vIWVXwVGQxSHvqWc
r6QGOilAdySjf/lBvytRubc2aStZEE8nnw1w6icUtaOFjmo8Uzd8w0fa7Ast9p6p
CoXxmhJVQH+oXYPSF8SKTRPZ0b0XFVuel01ZMxwYNzK3KDLW52Hc9Ycho8FMcKZI
w7ae22nnxICh8LwpDCWDjcTkXGWnFUQBWxhLrkXPI60cuyM4h2htZRQHnqIdck1T
db3cUt+HgUFJIQlIXQmUISlLmw8o1g9yplpZRDawqBYSwbxzglfcNx8G+cgKXZ1M
PiG/F2CxXtE0iHw0MU7qd7oQA2t6gQdvcarUzGK4YA/OK/EnYBKrREAmKws8NZdQ
HHj8Vvb0kJX9zovwBCw56d2ZdNHkKM4m/I/FsfH1NGB2pm5Bi3xOykOPs6rpJHtR
WYvi0LmoWhkyyy++G7+ABTHJ9V5OWpdDihZXiQua0xstAKqQCs3q136qzmceGRGi
SCNh2g+E9slBtEC4moyeKhgVYVRfkJFtdUled0sfc3wgSo3LjSiB9rsQMV9vpWIU
gLHq82xG8d5VHUvctUsyYhFNxs45P1pgZwsdYF2lh9n+rSLVIIRcpI1zNjcNxn3L
XtbPF6r3CGknVIsc/JQKn+ATytilLSRr2+AgDExqr4WY+y0JIeCeW4uKTu7uCiRi
VPOvq5gtCBGva1aTO3J9LmycfieEeW7PgMQiu2vGj+hmwd8YYtKlm7nmQfyoDuVp
fXNS3HruA2HQ9Zs0IFXMAocsZv059lN0jfjr9mrw0dqrKmcyDD5U83jqDoT/lvA7
AIS59fvvbyNRSlDdiwWIs78Q1SIBRlEee26T4tuSvNI4/54nWD9mx28yYPzcIPWa
jRPinYRWWA6RuiP0pXfsfPrIfuNLfjN7gqWGIgxpbBHzm49YXYQR1qEz42jtKcBm
dZBeiFRFbrYVUTxZ6gGWnNAdQ94nPwItNG6RcJFwhtRFoeN01aV6fhqA39GtdAsa
WfeBhIaHFU08myDS8Q7okE1HoEvghSL0kgHpaonviz2dXVlv+kavJbVZQ9Td4O2D
YxEmV47AWvX7JN0scCI3vOwWK+syiwhcrBt0fpAGZudFDl21lexXOOgEL8sGJH7U
U4o9COzHxM5xyyCyqti2qXs0qTg4CiD0mH5UO7gjswiK2v1MlCkdDZA43k/gaIT9
A6h3eW9PkjcWUeeMoXA0o7m0iBZRMq2dQBvui1hVWRGd8doTPxTtmWcMnFudpuMR
LDD7YjnPtakNxNEX20QLsPv79SMYPNDdFXuKnshantaYTVM212koiinJvIvQjf7s
ezPVbG4qAeNiM6S/gmdhMSx9dqPdyYHJipWgSzgQSrFobn6ww6x1UNuJi76pO+KU
ISRL0qH0Krp+xiMolmV4f/Sh9YbTewCRAjV7AHwfE9gMMvB0jn3IQVcuFdFJGTE9
eUox8LjSZe6kBBSAvz5BqyofiaAZMkVsgVuhD3nPbdi1omX2SUeIb1SM2Xz5AGkE
PtmsymptScwTNT1o5y77u+A1I3SfOtzU1wxO0Nh+JzyeoPJlJXD3sOxnmmIRnaiF
jD3rb+50ms6OJeFuX16WWh19qsuLkDHa8748smRHVKF5qThMYKtoJ1tayy2CQsBX
UZfK+Wl1DJqTaE38/FdhxgnlkTKJ8/QD+XPb4xLzFKfLh/5TEv9R28hXxocdUiwS
az+y7u6DiJCCGQUMEt+C+kRdF2ZDiwX3cXPiNNsaBtyTnVyHp8IS+KEh8KjeOxYr
/c4J2P7TGPGVdcbDZZToc9/MfR+b0DeWWf0Fj4z3E2zeUqwe72A9vkn/HDUNPNuj
CQc9Il0fx2oCuX4eY9lpzh1AUcEtevGNNTDlGWRbj3oCdPYTFzDiGu4EsQDywuWq
zJv5FgzTZuZV2t7WjQZwUyrrAdxwV+64t8lshxqBqL6jiWVUFLyotQCVwC1Vxs6n
mQmywgCszLqontL3q/VYQdDlmW+PAN1Aq1a3YHZZpgIOm9u5rTGMOC8ELJMRMJvV
Bsdaf80X+RuUV8OpAvEq12E03KJYBz1n9WcZgj/yhqKGIzlTU3z4JTaojrcFiJOT
G5JHeQ9ZIVbxLYLD1OGZ19iloD3RP6PlAzQp3S2My2W2N9paxQQSlcCu59LSLB8+
KZHK0C8YExZbF4T6Gtq9VP0mtOO57u9ABpQrPseKnN0SKW8CjbdV+WKNtzFqemaX
Zbzl3epMdCKURwX1WQnGZDG5ndbt8fE1cTXn6HbFrU1TaTyGklnTSmh6a5J8H44i
9xuhDB34DXGmKlVm2ohTQESMlsVd1yT+kQ8pN02LledAcKvwY6PV1DF8O9y83Bf+
R8SSdJKD+CGkQfU8w+JhdqO5BS+YNpZiEIIvZ10H2GZY8EoO3fZ57H4T8KbRr7m3
PiSxTgyN+5HMF6PCtbHFm/Ju09rU20HRsFqz1UyCBAShedy/iLSF4FQXFGLRMBDy
mEaabzddgdO/rhOYMIh9g2fLruiPGvpOgVyEeCR34EDoMuMQenRZ9A0gDkjNuC4i
qeAh08w7MspNcCUY2A7TSaU9LKptZqJ7iHKWJfbD57m/RDH4Onkr1tQebcdc+Czm
Q499QbHRLDFz0XCmPErl1Efv2sN/NnJLXV+A1wJIhXUgYujcw1Q4VsKfE9arkeuL
v5nrsiTJO0sQgjVGiLK+22pXLW3YEVptP695As/eiG7rVl9Jh4P7I/pbUSbiNa4J
LT0YagXE87FE3nB66zvQtHmU29yPsYppwzfX+urm5UDwNW3JcQNSvuOMnQVjfXMX
QLal/ZcStf/y1C/RbskfQD5Ert0aXrbDsKO4WA8E1UnlO7TCDaG2ci10BiNo8ZkP
ifYBKWMsSa7HbaBYgkTjCPo0+CJNpkKG5nS7qdYgGAUwpengzDwDFDpyjZEmiglg
2WRFwFShOdFK0MItKKh5oneAD8Kz0CIaZ5dqx7Y1jwosCRsQYmOgXp+9unQBIZyc
VlDNgQoMimmcLQ9gh+SnQMjKbffNyLNV0lO7W6olhUWmam5QyA9007uBSOxCJ7K7
BTXWqERJb3/1kc+rdfcTg4d5VnrMLKpLKZbe9NWUmT+1u8foPwaJfW3Bz7OAaCDS
9PCyEp9ix2sG4F51naKutl106WjAk56xhruyOM0OF0q2ak1+nGONTaBUwup5OhvX
P7Bj7T6u21DlRS5n8PV690fB5bAY7HcAZr/yRamYerf68XMDIGhDTN+x7i5X7avG
Hkl5cTZ97RTvE5Mo1nd91Fv1k71FBPi/TRiZmWMP9iQa26ctgMWvF9Lf/z7RGkKz
ra8sF6X1RV92IBSvRnw5APDQb7fDmA04fowKgD97HKG1oKpuyGTOuVMIlKOmE/ey
EX/0dL3BzUQliM4XczCOhkIvC3/9IhlC7rHXpJoQuQPqS4W9ynUXJzoPmFiZKnOF
jlF6bdNfzDDL6K7ErvwnZL7ac+idLvtjE9bdrcjaeOjFZysvyx4ncpEbqGpw17Iy
WLfkMbN3yg/cophqdjQY9k6vAE2cfAKkQd1uJFIZTf8ARdvZDblKXlbwlHFgMLmF
vAB6oF7DTHw0CYOZQubpUxBe0REdvRmE9GRtrsGQKrZbzxoYlY9mbWIzg0ZgcBWV
IDAlQjkILnbrfHqS1Q5H9FdxKtr0KG+KWYAptqoq4mG7aMPLb+C2VVuYoBRhWUFf
VuT3fiuon42nQaD0NXEjkH+1s4ISSbf8ASRI25BUAHN1lZhGCxyNs8elRTzyFroG
BZvgFbU8rMBYpf6Dzs9834smhJ75gIM7iGtIu7fOLGPISgdBQcyodMeAtxRl7MYs
q6KX7ACYd5BYJiu44MROXxN2Gv2gwKTEZEl5ntXDlBbzh+r1hGKkPUQbhdulTiwF
X46Jzq19H5zSYmSnrM3Emk92uDaCzHg2hUQ0JlCYUnzu6j2+LHGTbcbJp4JoBhaZ
hqmm514N44nFpzxq4n2koLaW2OgYnwfhLozqJrjp8I8NpGajAiwpHc2w4fzbJP8r
DhPutgT0wn7HCvlUAfKMEVy9KpK03BzpZ5vavOrA2bN0Y4I4i//IqQrNmemVk+9p
Qjiod7o0XAJZ0/hmm7lfIlTp/P5scvLolYZCfZKvx7l4WJrkXVNsOKlWhzjeV2/j
EPwNUkzVgkUV6KIN26/s6gbV0ykm+FGGCDnTpAu72yT8hXfLTMo/O0hU+VNaR3nx
DPFVART1Vt+iFD0SnVskO9Fv6Tfh3E8uqlT9Y6C+S5iD+K8HPSJxjxJPNLNeKh8a
FL3wNYAW7ly1FLmweTNY351V300iEoXJO1dVrh2tLYPhC2y+64JUhqMvCYXY66/c
OlzTPuNIV5M3M9pGIIzlAHD6mkMx2Ak/ujGVmUd5qSA1d10mRspg4EtyGBiY3oNi
xR1T1qd/msQxeZzBNhl/4Ky4RLuhzsqKIMYoeS2SIP6nks57eFguC9jNJmPGbSaY
ewpxm96kVkob7osIIEuEN7eo/ijvfcxWkEsxcEE2x36ogAUXcgmJrxEBxN2mnFLC
rfrGc50hfC/k16eDOo3NKqNfY5XxC2NvL95w4ERkDOtXQhVtK3zgGdcXOln6v2ow
sNWurFXIcTA3y8jR0I/TIRQr6gRpIoC5IV+/Eb+9n1O7dbIVy0iD5nL4D1Ca/0vM
ReN5X0jlt3FIz1dqld0A7JSGmifpmDR6+G210P8+3cZsEtkh242jhTLOWAYlyFns
NABHC3hqzmxMDrxtuNH2U3j/LvfZ6T3EXyiIhDXZLeOtse8jEd2ktC2JKPRW/l34
ruW+G51Ja2YK4fpx0xpZAaxsWY218LoBuJ0/LRoPfad99SU8a01JlyBkmdFU9Uvj
GYHdn0T8TJPq5Jy3G+/1ozz1SIiaBA2gIP836U/JqCxPtHoOUjv0BB4g4yUrdaot
+tk15dW6p6JCqVYqvCGKCzSxz9T8iZuLyg77HUkiBQHaY9dB0DtHWGwuNxI46IDG
8B8mSpwjfyuoHe0MvDVkXgzwWeecELKKb5aniN90tJ2jkP0A+J8kQ3hML9E60lV7
AYWvI1uq9TNyAS7l6sQq1TI7R0kywBZA3zIxr3m6LAuicZH/LvNct2zArbl0WYRi
E1YmzRGMHGEvAT5Qf4gXVCgF+XWUb7pYIjUSDt2gUuMiTNVg58+GRq0nr333iPxu
lWSQ7IQzpPrzbrj//qVJ56fCqVaZgoO9Yi1uoLPbeGzjx/EBdEAcnzdiH1Xr/jQ+
wjjN2wvY91nQdRMpVyEJ+POVnXTNEC0wF027d6C/82zNHLKQtZ+AgDySJR2Kg3yw
5td0c+Vh0hFJa6xMR8D0aQvEs2d8O3e2dAa+Y0I/6zOQQjfQEIrB1F9ZMBykLaIp
Z6ci3W/oy+1dd0BneT+kp8n1pdxMTXK+jjC2EVgCqsS0KCOpuQXTMMW9BbW07Okb
mlyvjzil/A96C4LWKwzm8FbrEvWqrQOw95YAl4zi3OpSLaGuvjPPKTTLiwvfKQ0B
fG2Vd7bb6XaFC1sWDZan3424xIcqLCZ52b+N9YrhGPaxuOK7hf3jG6GQRz8Lrqb4
BdgFUVX27wWo66a3zLglWYuLikdfrxfMFDtg1EUw+QKlCmCXfs+d0yQXEaoht47T
VkcOXuW5hq0e7W3UUUlZ70sl5temFLtCnjfpnsAipu4M8hOJOVPngXDVHd6M4Fng
cXqLp952bWUgPFMVCOasrSTLwZ0JkolUvqOFjttGjRaMg++ZOtAFaBrQgqmdJrDe
wgtAx0pe/OqLXqwVQ+Nm5y+pcqomlIdxx0nIFkCSLFcNrcsFfJ7msZcXNAYCK9P/
iXZK72vaL9xxubpqeUOqNejPIw7TZ+fCJcQ17iIH15qLBij721xkm8g6vrmpOiFx
cgi5mLvrmZyy7ZMEtE+cGT/0FV5/eHPf4IsdfeFNejqVJjG8rJoOQJmRZ2PhVGRL
MAZ37Rc8OFJneFi1s4uRT72WpiGLffKcyBT2+GGwn+pfEe8mwtqTDfxSoan2t3zJ
ld29O2z9wdv9liwR9PudijE0CmkfcjxtIyMw4jUAw+CUL5vPP8gf4P8Fcdjxm9d5
FyqQaAVf2o/w4vYL6h7JYnfFSh5wZfJ9lzSgmZ97C1H9vALJhqk6h2asPzOIbfcP
X2eldKGOVKZzdouBFqJVBkjYuNFvhrdLgB3QB6V+rdsDu/qakbeJ4M8I4n4ydpfF
JRoj4afdNHVN33m7L0HbSfe2iDJ1Txb0NkZW95NWzpf1vipuWWUb8BJB6h8YbYO0
rJy0AVFAf2TXqWePdpHkn7UDTqKFsGSZDxs0aE3NjDcphWxThvToWRQnYHZPCwHk
CcLcEEOvz+kcAnU1cyKVSwm0WEApiuCL1yFvu6z69sHiGkmzic6V58iqwFZmetO8
1A0+dKn76joNLbz7xh5qt5TVoFjOBrIJaFR5i8RE8uVIoWzNl2XYztg6GsIBUERK
FH/L998/G8zggrRxbIG3mbJ8l1HZ1I2oiOG34HX6FOhpbYX1TezUIqtSG4MekFX7
opAiksJvYUbm7YCcdzVwRfezhoiyZqGB+Pzfr1kNA8jn4sFPREB0Tbd6HKEHK4ua
XJ53CaH93lkSFcztITYYj/sFhpUZkVGCnHXedsnJnYNcSBjewOdTJW0eLeO67oZY
HYGDMXWXjqVwEoS345QuK8NHDvUAhpzLwUUJswhNLlpVVXCWkP1afNuTb2eTqGTs
1xAGJz6TMSwOKHZaDUVLh+U+pGNoybB1PeBQfEv5yCFPrwi72uEjTFqI3RrRTbtR
KKG/U2FLAPLgiYZ+/BXUdowKqwaOPmxRXySgtITuUX3EO4BnFxBf3pPXb2RlZ+Cs
eYgkjg00C/oSFubcHmcUjy3lVS4wyxvS1HPLpdn0WRr6Omke1TQN1vXBY0Ap9LXj
bBNETxt6c7kAxbb5+gVGMoRZqeqTVs7p6+G3dc0JRT3fhkXFGxGUzoZzk+ekIQHi
jpG8XO/4nfXVCSnVleEBwKES7sQFJRyw6elVbAFTvDyGjdcwWafesrGxOZdSryli
ccxVCmaAK90dBUcIr37T9+cnHBA50hubL1ezWjI96gg5jFOziG5PkwR+y1WdJ6iz
OYmWxT1MPP8a93wc5AT+UIePvPUIt7H5C5areskmgTywYROrljiszaMaVJ1B4FNg
n/hpZiQByzMLFq5+wpzGrOoYkDf1md2X8qUt8d+Iw7PLzsXlJpdchKNtYK3BDXkC
DZ3bwxi3dmZUQdAGWJZyUvmfxf0dlXCkXG5Kv9REFP1vawl60A6JJ4E6rSwc9ea3
48h8w1wiEyFAXJw7fJgTIDfcBrDhwdI+kD1R/6Oa6pYRdVhho95S9eJcLHXCyjsD
otcbOewOo6fRSlzYUggge090W+jLamIC03H733n+OtsCHAGyULR9HVmq6aGjK0Ps
DWNIVPYsHkJoc62ZTS37rDh4o0nLPEpkDRykCM6QuTrCVp0IEjRXHJvZyRJGSzHM
/offvmztOorU59nYWUN6svvBmWYh7FmXVJ4CUB02xH6sPznolySG4Lb/si8PzBtw
T7fm9b/AseDXFaqXU+Dj3IcKLLdQJyzTipdQ0NM9UDswPguaMqyyHRvs2mOxgZgw
9bCwt4EAUrjYH4zznjlXRWVHn7PuB+qa83jH/J/gtaPnCsbjfHEYT5XW9bcmdV5o
U6Jrm8Isdm8WQfhbbm4S/oKeHScFOPhHKACN+xq72pfCd/8x87u6pGZ27M4+VxjA
jxnw6Y2Ll/0LZIr6FRlvaRJOe+PJAFyjmOw06yoih7JFVhrZUzD2R8fVqrkUHHpM
ei089LSEEQ5FztlB4i+qvYP3KsgR0mYVljeRfxgAikK47mayZVA2IfM9HwJoIZNf
expvP25c8BwWyQ9PWwaoshgHxVoKvxgR/1zQQN9KhGNLYmXvjmkULQFWcuYCxBJl
ArQowtOersNumgBJ1PHcGtX0U1EUarz4ARmll2GbbQZ9lu3Fclhkye4DLdxvdAaY
HBya6bGcNxE8FUs2c6AIKpzIQNt2G5uaZc+VpZksoc1pEVCQZu5DuShapgeQQIya
xake7ihlWmM9Xk01XxLVTsWvnsjTgXcBNW90BiWY/pxl8oJEnFM+16TxsOG/DMsv
BBS2b82cWr6ZxEt6rL3+dqLflUOo9BCiiMoM9RGce8SJsL+ePa41CGSElzW96Vfd
xRhWfIgQErs+DZhEkXLAKA==
`protect end_protected
