-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
s1JoKxkAfRJGpunTKg+ImFHjY2wno9Mk25+FpZoT8T0w70li/VBJlBT8BsNRLcCY
aGLBghN9dfzw4gQK212mslOfOzbWMbba0DsSCaJqr/O+qHqDlgXYa1TLi0taTnbx
tPfFaJS0T6l9dZaDNdQLS48HR0Rz1irwbAZnb9OwPzw0g+7+llxwHA==
--pragma protect end_key_block
--pragma protect digest_block
zRP+Bj4+zK+wZWIiUKT26iJmSxw=
--pragma protect end_digest_block
--pragma protect data_block
xp92B8Dx966cXA9iCHPG/OuE1iWOzJ/p0GODedKC91BMioY0bzzwJOPvsKw/7Kvh
LAWP5pMTMkyfmXXvZGsVu8zWVCEdYDclyiU3KWhHN3fG4ZEoRFmxG6sDURd1z6pn
RrpZDMQW/NcoX+LTTVjLW55s2q38FHCbcEYU5Kn8q3FMRWaodY2UEZFE9qjqwAod
ERJOGbIM17NM8h0PDT9hNFgsmrSSPEfBtYsdZouhxD7HrIfsnfs4u/NrIPiNsx1I
IpWIegd0cv1G59P8C4ISdA5Tr4gfi9EwQuLPFrdWMbRLhfFLQ3WqpRY/u/yw7OZo
nGCPdpdQMHG+OQm1sEnvGYsX/vXLCb821gWxWW8RufsKaFLTCOybs+58YACEGaBA
Zyj7I/H8prkhxUxygfm7IzUWljCjjGlDbGRcHUnJRI6puMpaQuzlsUsuEIx91ML0
wd4H4YcWn7XhjzuAfq7Ct1NnmxOpqQLbw/m5aQ7CkH96dh0Rg7i/a98lvIBl2kjL
Vy2QKM7bF2NCQSjeXr55uBKL7uq00kJJUPvV4GSKzZ0JioxY1kWc74RA84fKgUfm
SfOZ4U3G0MgzUNqGrw1jKpts1g7VqK1wg9Uftw4QeBxeMJM0oiv41OhwzjowR/YE
FJ50MM4Xh1uoqSBwBIoQmDtN4CDmj9R4UVIYQjiZwR2EMIjIrKLT6WSoEUX5J6DG
ys9ID/f4OAAjDYYt926ebre19MEgngGpYStbPa4Sn26C4Mu6r/EB+aVdt1wcQ3ix
yLwfEPIqz0qfJKYzPQSKn5OGopGU1XdHK9tSM1u3D1brelYpQHDGqYzTah+HGfmX
hVukod5y1SOyOyE7rXc0mGzwsFTXBSFQNkiz+Fi3ZWVht5SzY7wP1prGF8oaQ6vs
KsIbRZmTwbNvttCI36kJAV5MlWjiMGQmUU2w+L4fYOZIyQ0/DXUAOaet4XPc2H8W
ujAxuefqOF0xUTHwd8ZT6wtpdyW4CvPM71+rk4Ul2cgXCW9Nfng7M+v6KsZ7YZNU
5X89QugUlsOckXS8zUFmxvzS2llH+SjCqEPHwRfz9cyAo4+a9oDgKvxl60co9Nu6
fOplPtS0kVGMOGngBdrqqvtw3ATfV8O1Br+5N/pyddNAJkCRdkXCvNThjGlEEXsk
Fhdj2T7biLj7uNqVOMc6jp0hGC7B2q6gHogDuJTvuSTaysYxlL7Uo5IYS9tQzNl2
aRjLfQSMTVoa6i8duUaEbDexNdZKiuCuFSvKa2486+i4j/xVrmm/AD/ilhMTN0cU
jIIqYUCoIYJ33hS6HZfZkEan3eyIUJjlugtshack9lMH3jYKoLFvd4hsy2C+8whI
YecXSzB0ywZ8ce+ziQtaFSBUkRjiEfvSs+4VXHzOWQ7EtIObtHq2+2pugAyaDRrf
y04XBSLE9sJqKfUWBUlu5wRmgNzCdkTcxVdjsW5z2xZPGDHyCv1cT5+XW8ZZ1u0q
Hjf6HH62CUDdclGudTzHstp5zApNvYFTRdPXgcCLIoKqN0I5jjJD3NQCTYBOe0y4
Qa4QY0tIJQCCejEnC+b4X0kjYcE+heAKJ6xkRVFTlsG1CiBWkjGlz3tcc3+WqZk+
wJqRavn/RI1tS/XJt5CBkR624CGgV12ptn9rwRP4jQjabcT1mHwwHb57sxHnce5Z
RqL9023EfAj+SR4ho2Uq++ZZH/AxOFcKew2ZkkGSYj5rhxOYZeuDq0NZ4mdtmgEK
MNfbSXVQHM2bxKbyo4P5jUPP8yNY3IKghVnRCrPTH2GW8HQIR+UEfy4sTRoFW7y0
25Wsvo15cqcEjNSzKUZ3hyrmHKqkcp4KLUIVy+TiqMV81d7aFZ19YZhyGHE1ZVOo
ru4hhtthHz6YtrHTqatNTmXqmAOmt8wzIUnT76EI//IFWufo33myt8GfKY/z/GFU
21RsPELmMk8Nfjo+FM0V5WGCa0TAnuPZuqZ4vEaKvPuzzc8MLeKFJR6+9qzINxel
dcVEtY/OZ53YVaKbrI6ArjIwKoNVvpytNMOdIToOQLp6874VdfDabFPT/rjY7dq2
Nln2b8OR5XB5GGwxKwow5buxUDZYgTVrauw0yMW5+yAvzZ7P6Gl9dOxRD6BscVfn
8W6twg8Vk0Ghv0RwrDR1Ht+C4rW2BLbGBXVurmvuCnSu0ayZ90TSzGVbFqhdiPOO
v+g6ZjoDFB7RfrFW+PqKOquXaGZJuJ2WYGOsg0epn8f0CkB5y6bT5Gub2CzVPtZZ
03+CD0sJEZ4Y407Vsl/89oLxx3BPsS+XsaIjX1YburzbEyQhVay5jdabpb3wLpcH
BIdshcyn+QPTEOVk9JdpuKktfE0yv5nEVJ46bTiDh216M1ekVP8wObdzTq/GV3V1
EH6+yjQZgRz7RIMmQV0NPiAUdWbwYuNrLEZIcOIILXwt0Yzjo9Tac5UECYx+Ktl7
UYcGz5rWfZzywjn0bHaOiPZEVNT4EGgg1XZKsj6HdLxHOt6lKg+cHAIaTub/iUGS
yPci+4Lu8CXXfeGGMlSsIqlVKcbf+oxPndJilHBaPTMZmO9EQOXeZYjEogFzgIKR
xmqg3LoGMc2cx5ue0SWCjCYF0/l0ohwf4hk7s2WbWWTI7qw2msIJho6Kq4eWJDol
/AMwqtPEzyAZ0Z4RHhGU2ekKo4MtCa9lE8jWRDxhuSmCipRI3dDxp1cwyOT8Kg04
dWKde0HWHzSyjrGUQjlDJ+FMh1fHzLkuJFuLDPhMMQ7FnPT+ceuPQAqNyhGaAxfq
8YDxHOpDoWnn4qQBVl2zhA/aA5VKJmLgbPG0hVYhe6qYUI70b2PtgHrx68DUjK7W
CwBDbaHOzQiU7P385dTlpL/zlglRnO4wZcy/IYg0qei79js4UxUyJE30iDeUOsel
hSjjsVgtxp0wCUQFf8+1KC6OiIu18i7X8G0T9qu4Co0qiZo9/EytytGFGvdDt1TW
Orx96hKrAXZCiwEFtfIVXcO2NE5CWDpPWEusMV3luduQWerI2Ugp/fQMFPi8BTxs
UpTYBrmlLimNviR8fXzajFRX8XBGcyvq3iceDufXHiNSk/PqyJm0Vi/VS79WCqvC
rGOsgDVO6VB9ljYKf0WYTqyNHmpfQh5tMiG4fK1HNgKlspBzOGHjKMWdRcjIwxnD
Th22ZQlfI42yT6+5LEe0uy3XwoqKcMjoo54P/zzRT3yU9n5XierQMKdS8jhGGFPR
L7Em0cvBzF6/Czyk2mXUuain5xhPm7Ys70wyCBMueurCk4qiH4yYBC/7aqX3G2tW
sFLvkkZdXZjoi9AnzMpTaimE1XuFRVggz8UYMwXNNudic1ko6k4XUySb2u+GMz8a
GTTZ+2iWjwy5smeqT9/vIPui+QTNEOs8wWlMBTAw9uXNThRydob4SE5QOE5/6yut
hzmjW/1XzIrkrOxvQnzrlrAhxT912amDRgDn7H/B2Y24UwjHBp+RP19W9ksXTbGo
htDSRG1z9XDYCnL7Zn/x+50ZvZdxdKSloy5pRzynvQPHhmOFOYVeu6FKGGejRHWd
SIXrDr1r3iUduBD/gXwDuo0P2abEZk9it7Hs7Fdezc9xbBWardkYFJ4oXEIu9lqm
4Tguy6B9yxIpKC4E3ycIXDpeSTOIS4dSzGEMDrJVYWStbh5Vb6KoDRFUnitS9+uN
jf0Lus8eevegKS7Z5owSQHS5RZFW90E6up23rFHRfX/dpKyExE3FpMtFLyzf7Qy8
z0Yty77j7/qWf2oAydUCOAlQ7Cll/W+zjSwd1Qm1iTCbBFUnlh5qXo779QcFWOKe
HCgh2DVolKLkZvSaP8CIJ0vJxSyz/VXf2QqSmm2LofRxWf7rGggDjShUyKBzcNFC
72IWSZFnmqvpi+dIIJgMSAVWNKkLRZugIMTY/V+rNRS1r2ouzRZroQi6aynZZ/AL
S9UKb4BMWeKCCLl354+p233ZcKC3c1BtJiEmqj+6hr/yndROuvA4DDV1X3LZzwzU
UyjJwGHDsKndxJtSERlKuCWOzr21m5M7n7/1MmSnLZwNrYBwbfAI1fv1ez4frxDO
PJEBe1WF6yFXIihwMbL6P8+VAGNMtMPzaohZR8kaK41C4UXvR4/brBo7kY9PtQPO
c4V4fG6mUGTH+FUltleNS230r4Z96Aao6iQmrBTD8aYDOCbSmGsiAQDKMdWxqQ0Z
CzGgHAUQAH23kiVefMzT1KEgdgedG89XcuZUWy6psllWZs3ykO+xZnAMFTaySn0X
qRJEajbmY+dtfmUUNKgBOp006wyMuE1yGqKaMkdABBts0O9K6WpJg6heiI++YnGN
ZTt76lfbJu3Xvak+KgsR7GgHQWXyqDBRIZqnQ4cSjp+vMz8gOygnvvAhEXmXvXnR
Th8hm6G8x3sswjgxxTC9RB6eQu+aNfK+Wj7dwcTdUnAe8pLfUSv9aAeC38YjTKA/
tpIoAGi+a9PzR1LoZ7cYnny9vZ/fungrU8PVne2wMf6qwA+lnEKl7socvYY5YDs8
k+LaGOLA8g8PfTo1HjDszBimgmNjL17itBlI21/p3Q7D5DU5RowhsF8WpAkTVue0
hg0XELuUCJoNNsb7aGIrytVgDhjdbv0WoH8Lp6V9wqLDcicRzzJqqyuzEheBpr92
yoqS2IY+UdQa1+l7Y2Xxg1o7M9r7Q3ON2x+I0zTOgd/8rzgKXrRDntE6a7rs4Lv1
1+cpGTrw7dy05UBOGx/PrZqwL7eB8/HGQ8drH+jj3+SKvNM0o+K2uxS1En6XdY89
5AT6i/ferDfFfpej7yRdWQkYeaMY/1mq4nIylETNRMYR0BTEJSCe9xhkFRCexcFE
UJACU8QGzXnwRwloMa09BojmoaIa+++QSo4G9B0fb8Z0UqCJ5C86SLwvLeirZuJT
OF8bO2ox1AuqlqusKcEU4i2y9MteIL9vDtHs3z9hyTtpAsZEgt6V6jyxR7POIPTl
O4uhjFFsPpADg7a4oSBkm5y/SgF9S1ugWxCFvPuvzu0MBVFBKl+diaSNAZtCavx8
gc++TCUew4R1aTjZ0E22yMU87NHjDU7ptgPCkv3UrdclqTmKMQ3mVGVaL4VkwDlP
yaqCgIfmOV7BM274LLflzYRpSDNjf215NVSMwpGHIAX+W59QJIcfIleMVcv6yxJ5
QDv41FA/yAAN+0L3JE89xsSIqsy+P0LbhrhOS3wgP5GrqtIGkdFGNZEYdCwJqyfz
/oJOYAdyw2nSWWiuIlH0ymGqpkb3GVv5seEq+jC0PXWv8TOYfLANfN0xRPkTOCeh
n4l+aRYxk02EhcdvRYEKD7Odpq6lGVkpzM/ckFl+EDo2203JfwqxDeNgzkh7SPBN
dp7oahioid7+jLu2aAgltMxivwl6KnTjiRmH3MqkWgkl4djMlPnPaCDUpfSRpTD6
SSysvuE7W34dD4Lq8/l9s9InOqrz32HqNEsSe7QWv89t6oAn8TRgCvMLifLrZWFV
PJQEBZ3G9i7RZ87FedxvIIhP2iiu4Lz1UaHcGN/G13jxoO0q5uDoJFR5ObwIShxu
G4dQe/T+TeI5ty1VvfgmAcp8XClgQXUJM1WVpe+dvKGd3G9puh4tIJU4WDK9WKDx
qkIrJTdLoRvCxenwblzpKeDnsxETEXOAX8SzOPx0U++pQP80B+o/wTYMDMvQHLBR
n962sZJ4d0BM1wftU9L88b8+zMOdvX6J3dGMCK1ASyXNygv9hhVKXWvdNsd8MXc/
Bxx9OSyvCNDmYltMjNyvI8wkGF1NprFzOJ+uPSztI8pJNfIw4CygoOV482EYEEG2
kNIqGp4HeLqNEOR+py/JFql2Gv/FFA+DHFKTCAaLM6dZlpD5TF/oe6bpZlIgOKte
GBFWXIUppkIn4sgyW6/27nBCNDh2V95/G5wpDNnE2m/2QnwwtKwteeCUiULrDmwu
3l0qCo+t33OUuW78zwzL8ej8r22JTd3qI6kNi72P198+eWz/YRcYYKiuLIhHyne+
BwQTtEdgAo+AzmutvmOFnfpcpM0QLcrDetJ6dxgcUAhIHVOS6rMh0alm05fXerOB
OifPyFT5lscVwrH37wraBAs38d6myvZRsymTZvOCmFyxnb1uKitD5J1GRP0Dt7Jo
BQlSqhFroKN6XlWkYUIKrqhBRNLQpnJm1Duo/pSf1MAAnKGAkX19v8hqGHD0Kn7T
o9RuXIz9lD4BDBr7pB0YdoZVW3ohMtDXzepbqwCWXVV2/oYkNvubZtjJPF8c7LLD
P/EQ7IfYuV9VT1nOuHYiwSQXkF5mybfLgNw2Yjcq5rC2pQtcAUap1p0GRoKkgyE/
OutnvGBcL1u5qG+GcAdzec8J9x5y4vGpGKyqPn9QfP4/sN7vz1G+UHM0m84rrCpQ
VINi4dczqT9jxlB16+1Tmt4gh+HqlARySgEH4PAcn4hzJKD5EFJcRZdDGYk5BB3z
Qh2vlLttuR9hWHiWh97NhuaRBv2vUVLJdW8yucv8Cja02MvuaIWO628/JFbwMt2Z
h4G0/PjVt0585XNO5QcjlmlXjiai1/NnM8Sv4e7/XoSLwHhd1/oECzCm3O5TQDb5
/h7mppSNuuML25MtNWAspQc3U2ZbbcDjJdXaZPCZnp8Eeg7LwIpm+sVpmsaiL97F
H/56fIEc4FjE6PXXVdqnzAXOBIuXVgosjZev9hGUQAH2zKED426VnaFCyPP99+wc
VMDpC0LsWaDQ0mMepEitm355d8Exc+DBsi+mTPhseKfGrF3elDhc7aVqzn5C/NLb
GFtRPnL06ZSRgZz0pEk7VBYjIJaqz3AhHiUi/qf9q7Q3S4H0CHikObLYXLICbdgA
ka/eEaBTZp+h37eA7d8wIKWdO9GcecFeV2HDkxtCl9PhxGWW5WULZ5Z7G0hF1sa7
UGJGdjo1VshdUBg6owH+6gQHcBtaKDZmi3/+rYhpTXazB9Znb7EBnwJ9PNDK2vcl
Y3PxEjFqdW/B1unWcBvmCntkMdxGVPoUdTVP3l5d14ZTeo/IS4Vv2BgzN1zrbTTK
noEET/xJHmvnJ+7KmEW6YrhbJAKidgiMhMMk2Xx6kL/SYCLYQh0M3m4dy1JHUWu+
9B5gDiOWjPoc2ugISedV26U4mQuekc5viymAULB80dVJsAXX7UZFCOb23DJa5Sj/
oY9UV1tE4buGzputdOPkJr5ErobGacpGhEsYragKENJJpcoGpc0tj5XuTg/MB2L2
3RFUG7veMh/025/hCjbaa1S9fZUX87QI32ydnC0Tl12SXSdQmKexnyVZzI5EHB3e
/3IIOabwf3+Rel8fPVL2xPrNCViS90zoe+8NSNvB6zDL3CFmKWEsK8WGvnUd/Z5p
HPXqtb5JVMGs1WrPEaGprWXHlp9jhvqGXZnSuoNZjCWhBqpvsyN2ecc6ov8Fa1+t
VGw51lvoxVsLb8R/7qead/xP6mDZo5/mJ+etR4zoegSnUSUvT5AyVSD1bGyMsW5J
2PX5eW9hVmcDgfFxYXdBTgSsFDBKxcIJI9eU9bcqalAVkBG/It81LOZ1lfTP3W1f
q7+E0i2bBcVMpBtj+qK0XYSLbjm0vms8rhgcLa3uGZ+JO3FrRZpcq1pH+kHlQyLv
9/wL3VIHbWCrUJEChZ+KAt69gRQekloafpfewS7bwlurZ9GMzLNv7XsZdOX7lfWD
ObR+Qc2GtjvpEViVuH+3unV4338C+GeBOVk7bInC77dI71KFvCCtZfIn4A1GlH0a
ENtn1LFx40GgBgCJUetESo49pU3oQn58k3MP7Y/N0M02rrLs0ReG4MJofN0IQHSS
9qMZ4FfOIA7ndur/GrtiEVO4Oi8I64gQxp0/XH+2HfpSwpvw3lyg9QqGyRH0jABI
ZSTytVVTDkHGa1U+Ya6xtEoGG945ScG8beZ+/ThFbDLLZGR56nqHmtP4mcXJ2hNH
3/sg1YA3lwpDtPCdQNLllbzRUyqoqUZ1tclK4sL9emlcUrW4nljf1RmigL/KYFza
N+UOW91ueg910H8J0bcQaJY2AyGBzhpXKEhBYWee7i5YvnVg/biuJq+sWXQkuYf3
nzyS7HJ31cc/MRwWIBRdtlf5DGj6Uu0UcsK2lca0CrmgpzauMZo48gJQbc3lc+nh
MCdPDT/UZaYfsHicD3X6at7BfGOLyi41qWxPd83H2/nNdXOXJuR1q+h/A9lWnGf9
0MraNivKcjV682wxvkmfusmNSPuh80634uIRce6fE6I005t9AxDSeMFJpJbHIS8V
9pymEBu5QJ/w7aHhKU07UehMWf/2dNKqOxsZUdAjRCCW2Wd6GGrsSFN5QAr070xm
EnzvkgTmsi831vYXbGPKqVPJGjI108349TMVhYuKxNRMbIEz1k4MlixGfwx9vTkb
gfx2ft3Xye21oJegOLrjjQJ02/BKI73Rf2tyAgTT7tHk62Y5HUgSwb5ux09yNrOX
uOMh+b40YQEqk21PTkqLQCWAT2NVYj3PWokTAYqRtxEfPyLTgUnArH6NLN30y70M
+DIcDS9KPhxjed3nOJujWTYiyX4/vI2jJzr6VV6JiLyYxB7WGNEZ040ARDp+lbLI
QVjDcmfIsaJJ6VbGyDCEMVJiG24u5jGvoMfoenSzmXRkesNDahLrUpV8gFVAmwOt
zHfelL47ei4/zu92XvIGEps+ASHGsNsXQgkdz7sZ4hSSNj6QSCC+GICcqkcqJtYo
x9etwBoC2lZU1WR7X04eN/q6qmgJB++czLYlSUcXtb8DAT8MCjYdyoPHYeee0bCt
mr10RNrVipOMXdVL/+kWOxNPLZiq0q9fE8zd/+oWk1zgFrOsZXmCzrA46NhtMjSP
1aFhi4uZ/Yb9qgf3FhpwKRkSnSgg3PM3RqcZDJbYS44mOM2hDI00ML/AONCS487D
ssh2cHNfh0WKLaTa1WJH7P4vPtVRIwDoEFm8c482pQIf8Z3oYD73mrltZM2y16jA
uxcwyXTbUAreFz4CT1j/xEfz3pPT/KZbM/+7WS6N0wvhpC9T8PHaOQvoiM6moRv0
CJgYHEU9+JJzlw9aZqVmJAMy7OOseH5GrazsRzq3h99/nvIofNOkoHHVCo/Vef6q
cei8DpQJbonxHy3G3xet28C4cVzjWC9cg04u4B+32maEPrBSrQKvkZEzzwA0fHK3
DXM4hL2joatXzB2a6iEnv4uPFOX4ExqPnrXuS9WJ+7VLDp/Incl1Gdd5WoF7i3ia
0dp4k/g48MBN0oEtDO5FDCtRpWtP9PTvX+m9vkHTu2koaO/peAEMmMdEmtMUlEKb
v5cTGYYV0b5gVl6YN6uOBz7Eyc75MBWJdfz2FJBqh4AkP2IgTpZZOx6LLGl7b3cW
4wHHVUphSqbiPq2S81lwov37bae47BBcjh9Zez6VW+qgIApfk6UTjqeSy6X3DCue
7c2Td49lce5q5Eu5bbDBNH7azHluxWw4nL8S8822NOCLL6rriyCA55xkUlVL0IrG
TAn6wU94PEOUI1fQAlMBIgmnHiB08tv9xGjZWBatJ/cFew+Pohh7UI9b7dAWZGWK
sg6/Me6BXDkC6fyn2Idq6mVxply1qqg/BzwPzz6hg6VLfHi5Ok2CSrOeiQRrUxcZ
UX5pK5ybUm7wdcQVJtbg0NEXngcBgWcHBum9GJu2+Ehnrl64lp80bIBXflQLGY2b
qOQy+cJ5YUQa0uxuSKznUGzfLa4CL09Y5vzUdJ1iYwYYGP7fBOXAOlBBvUm+Sa/x
1K+pQ6886EBzFXlMuJ2T/A0zk/X+ZxNO7xcG8QVB3/dZk5ipLIPKxIleu53unIiB
4eFyRDzbmPTVNEx9o0mzsirzM8Ftu1CNj5+3nRRhT/qdciKs0Wx0IlW0qIysAvBU
JnK2aEOW7SPelqd/rXeZdK20vFK/iufSdEW5Bhs0Pu/1u9MgS38cBCuGDzUvBY3L
lepc7KlQUkLDYycqFuiChkHF6s9wJCbrTxxD1FysVhCWnNVMLNmSHXv5LGYa1Lp1
vhi46fC/2/npPjZwu6G3yP91qYWmqg6BQHTW7UdIZL80rPrDKgD+OEB5GV72b7vY
Ppe2qaqRo+L5mlKp4xZfDZLnsJigN17symRsYWCa1NJGuT9G2s95aTCVuiInWfBr
KZ6+VhiQ4tKNxeaSnYF/9mlLKa028iUctw3DiGo8qkJIioPiCcVjsRjNa4U4N/4J
cSHKPoKDF/+Z07JxuzFARFSB96Mthm0nBJcy9WWPN423dX/1hRUZCoWwBDXlq7jS
JKa6zkt0Ym3T88kZeQzONOzHMXtKY0bx9fB/rpCspoNaNmlCGRPDPFno+hdriFB2
jHaN7SDH9MSCvabX4Gp0I2MB75rSz/V4h3D7GJcvMqTA1flltaHdYuwLKDAEXLBa
C7CoT42rlaPbibWFPVVD/CObMdFq91Un+NpXyjE2W+JfrNFsH8xHx66I+F3Ho00p
8HtxgY5CYqmO1ZdXFB64rSydxt1e6edoXwJSLuceNCDpU/Fg0WqslezqR5oIPQ6P
BTytOtSMIdcAw6pzog2afIb0EAI8Z/+K9w2yFOi4rPyjEp/gs109b3Ele5WDqchx
5V/xJIvZHtjBQGbAFALAc6mz+rgYQSLIdmsppRV9cPjB5aYLN5Ys/RDc/FfPtSqr
OGGDJHUsP4TXHCXc47YHKES9N7QF9I6wTH6ujaJpaQWyuWFfs32ckcu0mgBUgF5g
hblVMEMtpKUIKGNI8mQ/BI5136QMhg9Dgpa3KYg0XBtNKkd+y5rXgzytZRH0LKnF
rpkozWVoCCXm9Re1Rgy0Mrvy/mcBZUos1xQKuriRG92dT65DlolsWq25bNzjfQHM
5B7UdkSlGPVIVStOE016hn2Fl7BwuqKWO0pjnxxH9eIf6epsnZeklJk4WAYvM3X+
uGIHccW3/8kmvUCtSLkrrbVhHBmFO5i7uUmgkuNt5QHAv1Utj7DPg5nqZBksS3rD
OgQcFReX8OJa6ZoOEHJ783KD7ZRCVXXJwg9xywrkeeHoLHQ9MMQ/nn1Xt0eRQC8A
8FcS6MWU84DjQEuJZEHuJeQ8jz0bi3SfWSPGb84yzQe3MCkMR2sExTDC5nZg00IM
9xzQH3SAP0iClvvUw+yuGwJnME0ICTpvJBVK2nn0zlZXrL5Djxng217QESl6lF8O
I4QFyHpNsfi05AQAsO1ya24XRtzmFvcmUPJ27MWPtLG8d9kZ6oeZUC+xCfpYUYvE
s2zUfMdtTP+PDH57995sSy4B0dJ/H3mJNWsyybKU002tso6FsiPMZsfFPwu/iiKq
ukmjneJ6h0nAUnCoKaQYI9lpDN65La53S9XmCh2qs4vALF4rKNq0JHAuTy7/A8tb
Gnn+lm+JPErjjsvRYnyuGQlAVpF6vUm6XO6bICy+3j4ATynnpRY5mPDZQNox8gjG
aJHZGxO+c5yQRXd19hcJlYjLS8gkDvmSj9s8Lz1v9JOoY04ybkGfQQ6y6jVW24JR
pBgup02thqmJB4koTtEnHp5qjPcf3p7wlys0YYKk/2yzYVIaG5WXv/LyhsrfbxMA
VQSODxW3R/SE/f2hP/zUpNAzFBc/tuUK4UMem3e2la9aI13rgs4yr9Di2YOGBwxX
5PiPITqTNBihjIiiv0/VqfNjrdTfpHFsXzcSICVG4zuNzQv3YG1nDytQMHLsU/ND
QmcwoJScJi55JFWk0FmK6nvlRyhos+ykiNMLhzToPH5bysxE10cvg2gWrb7pf2Zw
qIiM0Zf88VZQKJPm3inar06DxWsuBX9+UMb1r93dhwIJ4D7XGncvNdvrzIgjM/6y
OAmr4DtKLAIOXMVVsa9Cvuq34vvsmlL4B28i0Nt8Pu6iYiWm8yH/hl/OV03WY9Fn
y6qXBEpNKkaKjoM5DMpyDJiIHkQeM32VSAA5clIxXo8HNF4/Ul9giVEVSlOLc7D8
/GDhkiSmhQ0fXFMATEyYOzSIyhZO2+sGRu45eCZpg6qLFZI3+Vg5CTok+EvttQqy
d7jrzznzMSNkRf9Pg0kCxQKmqmqAP3eiOsuj/eEn6R6c+YYXpzUd7himgEw9adWr
OXERozMPMwAt1/iZSk41TmIwZThQu/7/JAGtZGr+0nVBv2SK2KUMSeFaTvaHr6fE
THud5wKP+dH1OAp9zPMVZJm2K11exFsF+oTzYE5jRdl2ck9jh51OpoWfk0iO+XC3
IP5Dp64Qd+JcVGfrxOVtaMCyGEVFPglliAcLiGzwF9/2TWrLeB2+hTzF9FNx+4ls
fTKiBAFBOzFo9iM5xdN43vUI7p7kya/uI6dvG0/vkOC7GQ75SuIEALHTRn7JJ8vN
8o8KgIC2GJtMMQTTsPY+Fz4wMFZ1z19pV3+VTu4GHgbwqQj9gog6WUlkmhrnMYon
NWY67VwVU+4z0hNGn3L7QMH6PapuSYJ9shdyc1UB+x93gKQs7P3oIRFC+3MU59dd
ALm8xxg3wOrCps6Ho18CcwLZ7pi5oOw4FOd6OHY1YNiA3RHUhVpcis9zHVDrIEAj
I9wPjMW3SoTuVd06+T55Qf6glM2AMBpZws/+qQbMxFn3ORcEPZtDLp4sh6os/OiV
YbWeEYvv5PX8dvlghO+7b+zT0M7udw1I6EkpS46GBJpARebBwiYRmzGNJbbBVHxi
b8gPGfxCgQfQ0DOcmuWCI2rheTFHWc560/vvalRJZqezx+PgsQuRPysg1OU2PRtf
FqZr6a3dWHeasrDMclRQBHp1z/aaGUNDrH7Mk7fIjeDa0FepUcVf44x+MvjINyaE
MuzgTMHi5j4q4NiWXguXUDmZxgPaqWmAx/MaQZq3AOz/mTlXfOSbyM8Ke4mokwsS
HexlV3YOvvxmusacErlQAKQFfXl14wGcad/T2ExndyK8oj76FmRs5EM61TDqJOsc
l8WTzGmF5jYdRCfkuB4ryxo3KAN8LKA2yhCKjqYzm7eWuAYov3u50PtSEi1sU6q9
gvaLoD95AKWtnluMm6o9kEuChxW+tvAtWYBFxQ4IlAVg06uxf6tfvCxvOEjNemgy
geBtxkZvkQCeAfrg1tX6sPmVLrRBHZFH3rV0c4ctw6Ajeb/psBBw09OXMEm34y0Q
JGgAiMGQ7k0eG2SWuM/w2Qou4UrtjxKxamAGYVRgF7tLw1sgdKGlMK62ZAc7E0Ii
EkF3+NiJHMKlmX8fQfv90hqCLX6B7nkC6wRHJ/X1cTWZs/cHaUtyEg7wsY1fnB2O
sdOUi3ENl+tKAzOUaR09uayw8ancaJPnWSzG4ZHyhlx8yNwCVZ8vOu5d5e4n+usY
bvbz9LnhSfzbXy8qEK7KZ4HS4fGtV0zoPmZurRlp/3UqC04M6zPhrwD0j4CbFtJz
LSzod/O7BlqJ8kwsI52ZvkFx544SjlJJJQQLEowdaxbZijbCkSoGsXSG4czM+fB/
Fpx4oTeNEtQ9bG0Y86dtv1/5TAwKrbDWVbPNfnTGQzZbRfhGnIVTRMJy5KrmI5c/
YLjx94zPs/dFrFjJXDO7Y2Zm6Er8ybPAytg/EFiBNVA9lcRUG4NaGLPntXlMqq6h
8hsqUSo0LPHOwO4ZQjcN9+RbUk3gHYn66TcMv/w7wO9EudNgD3GYd0cvEzQdwmsF
3JRSZaTnS23EVOfahcFvxFjvghuaK1Mnpnb8+NjpVqQQGkC5iPloPk+6mHghEo1r
6U+q6pivu9rj2TOV3Hs/0ceuKDdG78Z4MyBSJLYMkcod4UthZUKc6O6HGGqdpWXF
+7ZumHvMF0Jf1sxYk1SuPWemcTUjFWkv4VdDL8S/Lw2qtWV/LoKocOAYbQFBrATN
NirOsg0qTr04PH3h3h5DDdWPSj4HzgwRx3uRWb0sct4kCd3ZWr0trX9mArmshxL7
qKyx0RV2lgEC3oiaA0A1GcnV05vJ5S8ZaapFVS6QdoM9wBX7ErLRU/8knL/5pAoj
kva6ftCKwxdQbSDCS6KrBz5uzCKM4Yj8hhikP0KSwuo370+SIVOAI0jjIX+/Nmfe
z8lZztHpmkvTh5O/mTTAaNoRIP906K6ysgC2ImlNzYEnLgSg4jiLT0MPwlIy9Rr3
+Zxd5KSEahr6HwKj20EUCxoUTI+RwMy3268QyHguptvci3pQD2wZMXsjQR7K7XMm
/9qNTfsdSqcU6H8nXDbbpNsShhSSwf8rroHRSco8GiiOoC/cQcB73N736PwcVg8f
0rEbkt763KHGVS/KhixiW5SSkpxIoJjcrXFUyYveCHeAd57Io0zj4LOGHTeHvOnX
LQF4T0Y0wonFxEu6aOTneGnoatHW34bOQ8hIb7CkoMhnyPh0rqqEwgPXUcYffDUi
tS5NGdjpAyexN/x92c4/tGylluy4NHh98f+vzsW6Oqwohjt2jXN/Vpg0NUPELLb8
u5ESKL2e+pi/0/bw3xF7+Q==
--pragma protect end_data_block
--pragma protect digest_block
l/BVLWHF3hkdNh4XCeXjkAfthPA=
--pragma protect end_digest_block
--pragma protect end_protected
