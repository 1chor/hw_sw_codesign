-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
YyKGKQbIl9m9Gug3VdvTPjnT68tGLHQYS5xSX/YXwgeMcLg69KEwz6rPlkmkGxWp
musgVW23FEhIYOqS64xrMun0KZrroAL5EEt5YDKhXO4E5nrZwBrAt8HhZ9Nz9nyt
kV/HfOLE3/74WDsU4rrAk/49+tR7rD/Y89QyXMvNFDRJQRs5bHvFBQ==
--pragma protect end_key_block
--pragma protect digest_block
aySqBR5TAOuHRxQNflgasjUxVbE=
--pragma protect end_digest_block
--pragma protect data_block
HxZCwSADFXQ0uTSFKevGbab44kYRmR/2LwACZRqfc4D5OG4ANa4ffUq3cznzYU7B
Z9sn4D/iOvo+WWZgk3wbS2TuPglL0LcktS6sDrOEIOj+uHrIe1AehhgQqVoSRaE6
2HLBUaM5bEhzP3K3qCiGCER16UiZIMAXeRfhOr+6cFsIc95fB/68Re8MxJBoEogw
n0LSgl36oSRJU6qoaPVrk7/NNbNvULrr9W8tN9nwI1UdSAIAU/qOeMANdS34WKPC
JjZRv7ktI7UITfkQek60oERE5SoZJc/NYSg5CxRSBXBE5yL2KEYT2gEgeBRbsJfB
3NcTfCPCb7npAxEKzCg06nQr2S91BGEeKkI2FInwzop9mMnA/FUxSdvYbLLnf/7m
9RgLGNLH0qHtEiHO3meGRgfLtngkb9mdUZmb+6GG+uFtcsnd23+CxJwfn65Q1yU+
yzZsHGfJxujsazRD9rypVA+1LXEgJWJMbfffew5Qs+4VYdjIq94iWd0IXFxh04tF
lM+52Gw0KyGr7yHmrnfPFMBDIQjjd5M081TeJmeOZzhyyKaFtGlOpvnlx6+gf0zP
ggnYy1A0RNGvawVFXl+7j0rtIFeakTyU51NmDgaMpH4JZesBASTBFMwpeODE3Zsv
1bxSiqGnU8hOgdlIyIVhiwM4dJMl53/wQcPBghJJuGL471QR6JSNq1ft/699sEwr
ttG7RyraqgU5xutsopxDeMQxdbG0RFP3wpMaxPK17jt1w3MYj0P9dDB/phcCRHGR
Zsu16bcKXDO+kTZ7Bk9RIRGf1PEXYelDnr3NCiNoqrD0Ua29iUNAqnEjoFfE1/hP
R06XzBOSckppiigGdoE5U8s9AyyPDh/x921G7/LIUefdeUQVDjYo0AAQ62vJu5tJ
q8gSZYl0eWLnC5oGDEmgXrEvMMyD5Sn9mk3pHOej6NBrQsC8d5BAMPs///Mtsz/j
L/M5nsjCC6L03T5JcVeTFgyLuNvtjWQRO1dxkErr5GvRVbURHe6raxZZ3XyqdNlP
QPMM0IouIELqybd0xleBiiUUS9ZgOJsoubwPboBDn2Q+OKDmF1SU94RGjzaPRd18
85DuuhGh6zVzmG4L+SIUrVfKQ8f1vjvZcsV3XGjTmeJvsglRLib69AMBPyBpIwNM
XvNr9g6QV+BGAFua7puXjt0FQXlv6HMHXxpDYdNRedj8iUuyDsjJmDvcuiKrcl2U
u9+9VevY7lfHM24LfQkQirdE9wJBusRieBm13Nkw91ghWMyTRffrea6haqOK+rP7
uyOreQ1vuTE4iby7ne7k7isYILMf7hmt0UvtRTubkyx2N7MOUEoSEF6ghzfYthjR
cj+oV1jnNKGPoSmS2f26oz29Wl1J9mEg+YznnIhsPRjANYyoYK+Y+YAaMKp7gM12
EhKrYBXtExelMDXPGvy/ZWw/FkGRJV4j/D6j0KG17LW4tWohsxN0459TRUM+Vbav
e+yi6+EoImbNOULBVm8/OmRWK+H+Bm9kx/HroslpjSNoeKPB4+HQOvjxq+LMDuJu
o0lrYajA5UF+gqyoKFZDtcl6uXBJIm5hkjDFnKmp8QByniJ1yNpxKrslFghJK0Ac
GgLFdf9N3g5bgCi32tI5PSGx1fn4ipWL4mBmoV0AihRm8Ze47WrakvHGrvy5OuZm
ODqb7qLIeMl6B+/wlWtuGOTwt8ndSaRvgK8x3lTbLiKC8Z/LOqPMuSuygPWNe+IH
7QHx1+eLinM1jZuyK8DFee+FYMIKfww0quMHPMQrere8JkVKenDUIt5AxdwWJE8E
hIV6n57GC5iUezMUi6iyA4QX5TBLrsrfjEXoD6dbJ8ds+R6P1aJuxv1dqWfF0EtO
f4FF1r+KbA1ho5leKixpR1b8ZSyWRzmHfgH7xJbPOASI9Tax4n+oQEUSNj6ZKR0N
Pl1eLhcvFKjZTe606DwS1VHX7lGDkJ+UZdRXMPUmBG1DCv9vyHNqCciyugqbzGu7
3hn7Yt+CgIa/zQ3Ne3tA4KrSXRVSeMLVQD6cc1pDhcWrT3ipAOsM3xeTHK/NWvMd
pR1zVVXp4hBRSXzRthGD9sYdjmQMruBlJTqJFwAYfTW4UXAvbpx9LDXcPJghlMHe
K9YdliK7VFiqSUEIyuuO+AMQaSIIT4i/WG4LjhqnzNF2Fbs2YaUBGXs2hGmFMgu9
cmdDzmsGGFqI4m/UV97vAL10Hz/CZGwqrSUlNwCZQu/93F+pE3Z2NZzgq6xUzfcN
jcxX3SGntwN/VdxKiWaea6qSCjZ+lNq6Zh729oXwfb9ZKNJYHgh4cbnJQSI+H1GA
oBcz3IRK5YkTcKnp75D5AMeKnQzCiVB0plhtYzMwyw0VrkpBj0j3VztoDZ+N44vM
JYEFJpKfV2bcPrbBo+Chmw30QXC0F7R+/nMahE3msL4IxUhni+Ju3d4kaeJhiu4R
Qzz63lVM5jZb5GFV+gi80RqC/mNm0T1kVmpyzDXZIGrTg5IrWKUN22BCebZpwMaI
UJz/de5Bs4Fu8+dTP2TItHxcNsnfkO0dz8bebOPGSoWmoc4sHpRoZJuNUQ3YBOYs
9HTtMJoiId9t3PEcaL78KzeH9avL1+/Zxrgd6lY6xJXe1r7TeGrKhsBnic6bdqwK
Q5PW+Bs+LC1/M1Slj/rSLV/jAqgHyqlZo3p1iigqOI4cBTsmm4hasBHOffgUEbES
68jSNV/FOgW/pm9Pu4gBOlGVU/GPn1Mqx7HAMXwsbFa2+BleaWhxJn/5imw8+p/y
RPYmtvnOcogZnUT+naa+r4ANhFpLRSI8nOYAGXkYbLdkintBMWGOT2oibvuIyDBB
7ghEk8Q7sZWj3Ffc57ffTJYZ20WpkMPdhAU+MJ1H/lCgDvGY+yo5+EX5Y7QiDY27
4scE5W/WWK+N2Bn7j0UjI8oJTwWihNEgNZcZ58rOlKlGi+t2v/yNqjVD6gjXEYUY
uH95H/E4zG1xSzlB681heBhM/HEMVWoDaSnr5ArgPK2D6hgDOznIkAg/C7CwsCfG
bHBwESk3oTaZhPtmbSi5uelFhN/jcWPzZxdThfnEt51lsqa+MoadtwB5oHJWAaJu
bmPyXMJ5B7eLHZceLuKnFsSBdFe+fiHuMVkkAFHxLwws5jctsJ2qt2vXFDNRG8RJ
QqwNZ0lxePDeE+LIRTAXgTU6yJDTPcSvauhm4BVsSVmUolo+IqWCTsd8Q4iCxoqs
0UghwYiJOzztaZqqc/4P4C9F7JukHIpi0dutaLGxR405eGHKyJDLq2UhKM+7BI6w
WdWLYdV+C7+Szwhg10i7ih2uft9EKVn9Rta8pf492OoKBB63bJUUBNQMzR8bjXVF
elfdoQaMf3/SCGYq9J4VjjayKHopotzDWGMeXBAkG5gbEMcvuMBHGt+ufvqvovFo
U0LvzdnyjbEyk/tNTnkONr8m5or+Xshy6V8+XkAZK5L2KRileV0OJyzTqFYoZ/Zh
VUWraqPHmsUd73MXgQP720SsIYKN08xwWT3aQypRa+nMO3OdI+AUInCFyVqGLIvL
1S3Lah/wKp+BzeU/CJCXG7aYvjIMWbpGdDANUdLxFN0sgj/mC+Jz3U1cMRV5ZNgB
udrBcJ4Vq3ftk0VITLCk+wy2vXwP934aWbWJAtWlgW+yJk+AxgLcyNc4eBePj19S
L8p3WqLU1oRWpwiQzh5qpggg0Zd84cka5+2ISK40v8GAfuJl6Xyofg/FaJ9LwXjJ
R3H7c+hVJ94NeQ2okzDaFvG4HivQokLBNJEInBcB8bCvaffgOsJEGUxSwVcMV5bt
1gvjSzij9uL92NCQxi4mfmyO1jRpRj5euORAnOiU9HbfGWVPKwXWmUp2V6q0nZwx
faxjqYE+w2PRlJhPS2PqyfV5c6TcJ+W6PRS74tEKMrdYfdymMLYiodpCGH7f6d9G
EVRLbmJvpw+3tfoyNGHANkhZo9/WJpWDiYpWCFHzzMe9K8RkUMOFisUFGO/+1U+Y
3JRXQ312DmzALFVCgEy1V8DMObJ2j9eUxyPFxSPSI8+EcfLb67kk4iU7vsKiUWkK
cny08cinK9vsCo4SYDYQfaPJqm3s1Tzz7Fd9A2rdzvxVEkzUNG3Ti8UsbIBo7ZrO
yOfu1q8h4oF4/IEUK3LGfb3K9j6NgnEVskGZVmEduziqlE/gkBOS58874vuaAXAX
tz7WXNUaZYQn/N0M7cvHQptECqF14w0plYTG9faELcfjkwvF4x7b6pu1t5b1BbAN
qcDEdR+94SFVHj9S6KNH9kwhEUcU/veELY5PQ4vbb33eJDfXkEXlhJzm+u8Via1Y
U8T7rMw1rwJtMak2OLlOQ3ikZjD/AqpdzZJ/0kAUMuiFPmwGRuvkpzOukAven5j1
eIruJxYnWsVDQ0s34t4xL3liG2O7vMA34F/uGXTRmlN42CC6ZqB7FYaOgn72CBb3
awURZvSedZ1OGROiJiiN6UNQAVVB3+0byzdv5iIMJQpGsIwNiQZ3BD2cNvWDaNtk
SoECMAVdyxt8XwpQnmmbSM/6rxTuDQ4ysg1Sd4qESaEIs3Jq3jZfk+y7ScHegsP9
0vFu/XiVCZ8cBb5b39LEQaOqzFIcEIw+sTML2k6gzYdAriLDdNQAx7VoJYTtnF0y
xmywO+M9S9HVALwuGYyKdAxKCFVaeuALJWgjZcz9FzN7FolaW6WXmcx+Rqy6Gb7a
DPNPtOMy5c4zmbfDymrNUk2FJuf4xZRSeqIBU1tR/D0bNAz+eJi4P8KpkilsxQQW
JYRvmVfZHwey2/PaVWb4Xi9+Im+BZf+epaJqrDHUV/WXR7Zi1Y16NykcuYJgbWJ+
7gem/QZd9dS99EK5wSnvuu9IWZmL4BOg4rpg234VhzBEOVdzwPMhvxzWP9vgTt4s
XQ7V3oz9aPGmhgpaPJOXRmK9/Xxoqs4B3NliGXQc2baf0RP6RFWW4J2xJE3+SNHU
TqOEWgfkDlES6U9MEfyE3PvE48X4IeL50m9G0wY8pv7NytIPPUsyYSonVptsIcvD
it0OUa2qle/DVBM8glknNwAlLtfx+0fCxqRYESUshYfsE16zh/O/o2mIMat9qkOL
S66N53nSDJHbR1G7H6tI6MInSJzYj4bX91KytqY4OIL/9AkiFd/Bdmwr9m7Zdt6v
68JQjaTlBVvDpN0qA06eayeVFkQk0OOtH9sG0GbprxTI9GBreKuYMbIIOIecynRd
7EAcBoj6pe+VSVp2fkrpH6CCKqMw3KHYD0aasYUHnxigWfd6ky+3/VggLF/zxjAR
ZxwXHMBan0bWh59Qp8kbR9PiUpFo/IUghkMWbNfcYRiRcO3nml49RKWvCSzOYh2Y
vYVrWuvAsHEmvcByuwHMVeihif6zi8d/WVOf81I45/XDz39lSOyOFCIrvEvmENsJ
IsOzwL/9BHhFMdmFV3Xiqmr5gaqjC1WHRu06IQ4w3Tqs9/6BhesWuIRCQYeb52nm
LlLfItHhRL7CQ8u36KDHXgvKHBUL4OV1/sLPv9GwdzCbDd5Kqo6cA5ykoaGT0D4h
1lkcz8VpPKR/banAGg8vdgxSsKUTWwwDRbuw0u2n9mZvY/f+MgBlTAW1AUtQJyVz
HURuGHv/4K/4B0YomIzViDn+tzHGR+//Q5s6YFZzJOpbKv04Kk96FaXtCzlbpr2O
uwFxgjF4dxrCYIalNdRLQsWDGibjlY3Y/CGDEmiWqIZFckJ9FHAlCkI/CGtwicpn
Jsg/8Ps3hX8ObNASwd3+iJtXEnwK2ZorpOjeQr95SrCryMY2OseS/TznYYFrpqDA
PvoQbIibS+CWUg7QynluldegcEicDGoClbHpPfzZBLoDeKuPkay+5wVAl4bQaHuF
GjhS+qtXzFgCraYxRTXGsjWxc7XVWYFp0qTmMdCNSfo0kH0P2Jft/ktIh5dcAj6J
hK6hOYKKu04yyyYpVBy0ecl6zotRmSJZFdzzHsqMGBjSUoKmoGitn6giTawFNrxh
hJWcSPtCPU+teHkkGRk9yVuAAS6a10C4QMrit90mZCUjTDBbjgNegU0+euCy43Pn
C3SwUCuambVZIGEBpR0Ug1FGjIovuEI64ofzk9ShbC3bHvYm/lU8EbBMMJtEk+z0
hZ0s9wloJCTjqKD28LBIDsfSgHTtZ96qaGrGa3tu95NOBMiHKcagdBDg8WsUkvBu
DZ1x+PfwBMAjgFiKAoaPfMIIgKctV2hR2VgKf+Ap/PhyV2/CQRBoGvgSz2fpOJEc
gZRPU2A0GRvzH87uwK0Vt6QP9S3Tu6atQ7FwHIInFPnKj6bpxCPAZahuZiiBY+IM
YlwlBcwqCPd5rn8h8fYdr8uaRfmZkoVQyr9us240uEUxiHJkgjhY6ivqUrxlKAla
aGmgay8fPtu5ufrXClo71R0sA14Y2dSDZefu6ISI0QVhaSyctAiJfl+JNeKe+sgr
iVxziC2r/Lw0a+Lkrf6mPEmEwpRYFs2oNc7jDaGmsE/6sWYLpJUckE3krlKAW95h
dhcU2tB/HeuFmVeIbPaITTLOs//WMyQ+UZXHDoLbDNgDGBQwUedu21z6zDtnvCmr
m8I0aL747se72Y1dOiNcaIZAN5i8OmHNzoaoOGYuqgstN9SQ+LC9kHu1ifh2mN5r
wpwhIw7OVMXDeHn1kyY9bOmfAUjMPu+aluTlU1wpKL/GfQY9pEZ9rdzLIG0XE4LY
phrrYzTxiN1T+HFcARiKzdSUvTm+znXEvUVR3Df+w5zgrGeJ0r0KLYOMgX2BUjk+
9BZp9O2ImY5OJvhzOM4/Zyj6LVB33GMIAmG1Q8B8f87p32qxDoh03amO5D6FR3zA
JPUXUQ66sbDKjV5FSWn+Oi+1S2k249dc0/O90JJPa/R2sNC0GMCcJIcEj86ssh9h
u9GKi0s+lmPhBQzes1xPdt+jyeehRpo05Ho8OHS3mNiYgO+dgVXK7r3D0Pljl8tu
oCgkY0W9VnsBp9OQw4XaiMVbpj9x8GRtC34/z1E7uN5sd0ztxTLpZHhPiD4RWXw/
yb/+8S/uwRevo3HEYDmefN886V/GXMIQk7BbiP9zwYPP6Fa+58ntVbT5RIjweNxS
DtiaE3ToLaPTPKbs0DRyhkEf7VEebz+oTP9/0TXflDAjtV5pj9KKmavCCo3Hknh4
/XrK5LlbwCVWlUwYDYnRvtLMz5NAdkwT6xrZVDQmqUrmTKO+S5ay5nR63Rxl1i8x
3unwm68k7VooRWRF8V/6SCY0sEjzPjnVdzaxzx8sCVhYCm3g9E76Ou7GZNKMqnwt
m3agrHYTF/yI1OXd4R3JI2O+CM9qJgqbuuSvQ5DbE8CpmeHzbNHkctJpit1Hdytf
N6ckYLEilu8V3MGWVCfIv2L4StsmDZg/cXqdAeXKwHCt+d6hY98lA9BcDKBMHtBI
zfuYk1JWjujeFyjQMo6ThhpbJyz8xDltlPOssRnhuXsb168pAdrLwgPCNS2mLkuN
szxDZqvufYMv51h6UZ4tsWmOXYXWvLjBmCwXdvlWSo0dufKmvAi4cqSmoI75sr3z
F1zUkcqHUdgzN6OdPiUF/z0xjcL8fVUj4h2XWX8YLjSa7pX4P33lcQ8iQ8AT604Q
4x/9iBp7mk89fCPU+ehTpQJ0ASQtrcTeAg9S9DztJD1U8EoCmR2Gism9G5tVG4dL
s7yzVmOzWkgONfwtCDgB2jyj7vuunC/HIx0Kk/5CKJJ4/zAH+U1NKdLLEfMrJ03G
QwJ8Qh6m0nPSwvIdXn79ObwjB3d0rFpY1+ti5D+QkRXOccn89+ORYVFYYFSDbcQK
m4jLpkPL9vTLqDfmB3a9+/Putxu6bxrfYFK+El0KHV+Pc5RmEK4fcq9Gi/XfgFOx
DoazIXFND/P2vPxLta6IcGWnvxoNAnSMJjz3zdNgzNOXaZo9fAGvIIEul38cdC2i
yKwDjuVJKVcBGNXN9/TdWO+JAN+Or0mnfYOq9UglOlsO5obH1s7VxU9ct/jEsK60
dTIsEJj3rZhI0ZY5NqRKz6wbeHGMzl2r0LRleHJuk8TRB67QbD3oRFXQZuVqqFgp
l1Rjc18Qx/vY7Bo4OJ1D/fdtHVY0Uwyd0vidaQSR626rs58vTX+PIXzHUW1XIRtb
U6fOo6BddyOxcOG1aFw7FiLqsqkNcxMhHJokzQErYflWa0zUUNPiED4el3LY7P1P
NPF1bNGl8Bt+7BK7eesy37EFttkSdmAzVJt9oDNw8HJNTaGu0x/p5rAGPFmj6gNS
DeC2yrWJ+QwHrxBRgTveTU4lHH8XDYBH+7B/d5AV9cFx7RzyhBkahQ3O0rbd64CK
UYyg0lJ4CH7WHr0otYvK9VeebtjFrkOs3XNB8TjjwfzeSG38hQpLezrrK43sE70L
K2pdNu1U/lZyOu1+YYNcQcqNFHeDhv2UXaKW6yjFzY/xOQ6mS27Qgi386t6DJfwC
iVQRM1IV4q9x2qr+/MEocg3jqnR6upSFBmz2Xu1dn2cRWgdvkDQN/4GOdmYfnUt7
icZdkpNJMmraftMWl1kYmWePejVSWAMcPJf4e7HPO0hDpDnMM+hw6j0fs6VMDL8+
EzzhIviKhIzmHcA2NlxGphlwVdrn1Q0z7lbhzLJQ5VMPx6MW91D1/EOJsiltD4+k
Wrblgn69tGIm4q/5CIwqdgeIgKUHEStt64Vv9YiItKrhXHiAoDUnOZzZMR4vBgCY
rfWEK784Z9+gU8puL9W6f0Qa6+3X6OeCL3+aGzhx/dNWHDICtvA1GwQxsjN5ohRk
oMk1VqFP7GBJ3NgIZBEY5JHFFQKSOPl/QEKPo403du4CoQ2/YKrhsFOPM7a/teYs
UAJNnTFpv+8vVE1B88jXOf70JAm7XwKTW8ES1jhSpqltS5K5x0vYRMxbq2onkelT
+YRyNedvQbfZHC4xQE7d6PtPF283TSFAwvdY1IHDaHb11PqFKn+pESFv/QtOg22J
JMXKzxF47R+siGk5kWuzstNYg4xWzcQfeytDZp5TuNoILthwKT4HbGxxnqxp5TBZ
0dfTtswlJI1Kqcr1Ye18CdWPT5s/EX6E57xnpnGafWUowVYfEw2l8T0bhUvplsIQ
o1YKwPne8o8TVuP54BumnPXwKiBVbWLZJpi8dqMCON6ib6NMyBZqMrIogqYrOyaC
dueD43f6rJxH7trlKbIa1QA1NNAjRQW2OW0W7cu2dOKviSEqBxQVAu6Kr1oFawag
HIdiSEQ2m9qOv3FedRQbeCX+evzrSmxmtD6VdfygOO6BbeIVkKMEhdom2r5+DcS5
VDUQ9osSoppPkEIcXl1Xk6tLnCgcBYkh+/JGrbeSWEDiZ9qh9B1VIqr66KSaUbya
3Wi2DVVPDWSatZ9tWdgehC9aV/kGeYHOvMUqePHvmyRugOe8C8OU/DcPkvKzYoP1
TJdCujKohain1+OC5p6QLS6j09VeDAMAzFdQdan0J6hS47ZL/Hows0CUnEVLbgHg
KzY7ZOxFNf9/JjCtXzeqUNHj1DzucA5d3rCDxgtTQC0PAlbp3kjo5VXFM4gbLF3q
fRcIk0SsRaDIX/57foQKizguOf5m/+m5jnRxU52WRtB4U34TQPTGSV7ZKiw8Rbxu
vlef5cDl1T4qqHNrimVq6gRtkxw9YwTCCojb4FaIcIpAwrxi5XlHfvCS5tPmyzjB
+9n+N7uggdxbBPZaTToJEmCaK21pi4sMVoV0Uy3rcQaPGtTo/kJvVtqeM8sLy31P
CFKvkrJklKgl2uoa1LblT77nL//pOcDiz/B0eOpyS8KxpLGY92YJ/PEhTsqhJosQ
4GoKKO3gSTsKvqFLbmJToY2EoHW2AoUBkdydtT76Y3fHFsgvIbbxzlHULjbrinIo
YYesZ/rCtpS9TfoVu1gBJrKCiGRg+eXVmZOaD6Fi6pooF0Jl6euTM2nedkQi6oR2
+5Yu9QkbVDXU68e/YO9Dj53qF6JxEigVjRD4MY9TxWzD1eXmQVMlNp2WBFwQgvGh
57nFv4Gm84B8HfS+wvUHXU8TJB8gVa3AeYxGyaglQHQ5OO5nN5DAH4YCUMlqiQmK
eXAuz4gCaEqVnggLjOt7Vl5x1hP0PwhVjvO6MET4UzHDmuRI59GqsgcNetNKE6Gc
dSXtzA5doD0t0tJrftYOn42pOsFypiW21QT55fRD47wPiTUU7D8iHfYhtS4PonQM
5nlnB5gFkA+I9VuaxoPYHbpV9a782drdsleRGMM5vCJzSKgX0aP/KeAJAvyug2+v
DFV1bvFZnjHgWpj+eN75esz2UtzyK9PUxnmxEBTFSsZ6VhNIUFjHagx6z1NvOcg3
t4YQ+P+++agTMscMjUIuGVpM1ZQVlKT+L0p2bvYphJ5anSLr3rhqxvB5D/kDWLC2
sEot4lC2myUwrpg7C0v+sHzrgyKpcIa5UUJEkvsy7tin6WaZ9jGWuuCnfSdZAW0l
TGRgVBKUNmy0iKHcHzGxWLVh/5NOa+HPvWcmNT5gStLydZ4qqatQK/vrkitl0ruA
PfF7ZLExpOOt5hdQOXL7/mBBQWR1N410vJba/m7O1m5H/XJnWQ0zfJqtL/GId4hx
ay0jS84bJnguanjAf6XM45s20VDB/h6ciR3FF+55ZvX4bUtppkKXFY0ysIDY7bV5
r/6e+7tLHLIp1W176rivlrDcM70X5r5C4/9eVEYFFG2cr0BBm+fAWa+pjmwk9+aQ
yqWhtFMhUC8koQlTYTcnlcC+HM9eXaCf7P1LBcO2+D/j2S1z9DvasE7J2xe5l/nv
Fn4S7hOG22tREAD2J1pGKjNwht1pMeqankPIQJRe6vVHn6u5C/o/a8P1viUdUzqj
NVdV9ZN+XOe9tgNjxA1py/s+uA3NI8VbWATJFWDfh1p55P0p7QrEFpAY24n4t1Nj
Ke9ZPXJ/EdZgUkqTbmYa/JbBxAMoIiDcdYBHxIk7i4hqzusXKiin9SEi8hpIjQDk
h6k4wkBxi7cASi2dql4h0kKu2sahIkuurhXZAvQOjXbvVdSUvE2eUK+tE/NQHyAa
7flzxEGoi90FdULXC7WRx/hxiHRYs+UGtgFzuQmzlt9SAzasE7vu2nr5jRUxlSWa
tyszLn2256FSlpuahad8JmV6KlBspzvj9RLKTvcQddSWqDLdfTn3B1mH/7OzxeeB
n7VUC3S60jGMv4xjTk9ihFjeoomJ45D/yYQJkDY4M+ijtDwgyycrO95PV4Cc9QEb
rKhRefWy2qmVLMkJUtGx8cdxrJ4RTq0IRTnwIAC/OfUUB+0nv1U9TYGwU3NwSbmX
f69ZhazakD0PJFdrVmdw+ZVSXfsWAuDOjD9iPFyvwQIZH5Q4clQ0MzdXn1zGe6v/
K5sRjtVnmkC5aapVHpaaEtLsmIxLRGvqb4aLlUj63dlavdCty6tfmcPC9OOvX7HC
Gatmsx54KjAnv5VUh8QmjHBa5TBmhcrLLU/7Ubw64js8Jt9nh+ViMyFZrS5SWv4O
w3/2T6sSdE+DU5JWC1b34iMZwAhvYF0Tv5UG6WLyJn540r7J3tV++0jgVKVGQn7C
tjpUFTXfQse+q32RfuAaTwUpDucHg4xI/glm7qVF2H/eFCbeXO7jf9XNCZIQEiRL
LCPa5rlvva4r+MKPPN5tM2FloD87rSSMEsSb4GOARlBjj+u8wHrlDLg5ARpCeMhK
J+D24yyE0i1257Qxep0nloj3/pkb+on9gj61NLAZASu+GC3ge52BJqHNiXFF32dC
fb/VTQOINHDW5tIqxBGUGod68lLC/FABU6eXJ/ebE5L2cA0Ig4XDNf1elEypx96x
hH0nAUnolNCw2dupYcC+85d1zFz8/1q/Rf58H64DcqcEcfe3HGVIUUVk/4JkrTJh
nuORuhqfudAQeYUGGtp7fSCY2odMb50PQKTM0GIFsc9b0FZRzYH/Zlq4gQMUsF74
+Ct7pl+mZscOhxFDSSC6YzzgrXMAvMz7SI0JXsdq7URtT/H6LB0tf3B0ZPii7Q5e
DwCkPo7Jt2izpZja3vtzHMFaQ69MQI5ftt+N0B4To/51mWpq2QmIP3+5FK0/YQMG
RUK6H3pUZHSg4acOtK0yP5U0pBo9mFRBT5VeLYb3trQNSdoXrKCtfdTdmfOlw9lE
mvb2ZawIqrABuqyWTNu579qmOa6NA6kY7KEq7OGdmZgbRjmKn9KuFyGHdfNAV3c3
YZQ+GSQhTyTJJa8CLmMPCTupI1h87VZP/syNWesR4lXMkyIKzv4lvUwrr4rISusk
YomxqscLdE5RmvGTTIY+TR6dXo/uYYakWak5L6D2qgAckxvB0MCO8HxHlIy0hZh3
zhqcP+FJ1etjID1Yrjjso3BqnvRFgwDkL2an7pcPIbw7O4PIUY04d2p/zlY7MWnG
WDCQD4LTkd7XXxSihgFz/Ccby9XKLCWd5a+Ft8gX1aLBxiQOI8q8FB96Dh9gV+b4
OgvAF1uaQjzF3XTX/ZEFL9+6Jo7k/iAhe8v5tr2S0ItDrIU/O3FVLRkPSCWNHPuf
C7WODm8ESflktqoZhyMgW6RvEgNawJsgX4aXVnHBvyXggEkkB47xB3kwBFt4SO/0
uCepzwPSML2XICUvOfB6lkSCLRhlijWvsiUfR/A16dZ4uEMSnLXYvh5arImt4I3L
19br2GUSwSxes810H3bIKz9RYTodxktS5EbVRBgJ7CwBeDVtwS3aA2jgcBIY6EkK
SbHWRpF5TGER3aHRwt595ZpDX1jzg0BXpN0wWIwVQl5+jxjZvR2LnaPalAuIfcYO
ehIPC9HP1Vl5DVn3E6L6FIOeytEFxgpsKsUxdtRHF41kVnriIcpbuR8erJqAtQvO
wIc5+JvTsZv/eBjH/GNUxdpWkdi81iD4dC+ETp836p/CYnuVQAi1SXTA019OQExl
8TNaQj2TG/HcwBdJwsGFJIbbaRuhqRexnyKpnc475Sp31XS0O5aiVtIOtAiWtdC7
PLcScmc4u1zSc35/bApgFcLlZZxht/BX8j0chvf61jYxnM2wLIq8y9N2yzJir0UI
5apknq39fpmCANK5Hj4t6gV7DIZXVQHpqn0i0AmGslg7Mjp7QgOgBXsKFBYaW39X
Mju2FoPAonb0m6q0TdHjHdYyp/rqtr/aN1Rp4ZUqClctnzYlE88vBO7x9jGN0GSu
1N4J0edQjqB9WxRKNXv6hib9NEmVnJMLSGcBuxMTMifs6pG9bDLm75QshuLx5kbr
ni3QPU5EWQxq9sMLUiZ/+yLAoTZZSnhXFOF70cx6Y/wbQH0d2ftMQlWAL+NBrcgX
RbNeJ0rpuoz3QdB8xO/vh+DtBfk5NPOVqqQijOoCleG2o1J4CNLkMdyQfkb3nELm
ZwQUrK5ONoXWjoIR0vnfv1mgHu6/JNOcoNMEiTOry+EB97t8fKHObE2e0GbbRxVs
Y/VAYNfDBXcryGD61wqIdnjD1y3bq1YNc1DpNsruBKLObjcw8DzHYWCQVaiC7TUt
iUWbN+z9yXpPEfo9TWjH6q9pYeZDhtAOTiOx7z9RSGpfKBGjukyYdd0VeSGsD0iw
PdsPoMYi9Kx7ScT+I2wNDrfJqF/FDv18WI6Mk7/cTUZDE8Z1QGJvuqoc8OBueoNH
tvndiccTEmw9m9/USnxokzpgnSzNndUUeDWPQYbdQkHO8y+AQNlBGyByq8bKovdq
fDrkEAZJhXO8E6U3EDxFG79SBYcf6ckqJf8zdDXlUM5dg/Ni3qJqgYtHzc4fcyv+
NDvtknGVCp0uPLUy4kG6u6KoVTeMSF1LoNwIhYg2Pggyuwlyno4N1mTo/14BODzu
L5e2rC+qycOelMPmsbMNWg==
--pragma protect end_data_block
--pragma protect digest_block
zT+4LK8YifO9vtkrawQwAOKq7eg=
--pragma protect end_digest_block
--pragma protect end_protected
