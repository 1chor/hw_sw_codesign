-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ezMcygi+KadXoB5/c73rwGkv6jPmGaq9GNaGGn8jauO9c/HXYNXSYfs6b8OTqdUB
atQtgBkeo5CPTPO+Arp6CmqJ6KufIzPkAj0muLOqVyN3raPmaIiyCm0jrWDO/wVr
xOg066pabBdyssBiwow7OzycdDfob+hR4uu1kyW9FlY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 89258)

`protect DATA_BLOCK
u2LvfRf/K045izobzXULjB45rgozWDb6YC2xdWGS5ormOjRkerVy5q1xodbOUA85
y4wPvZW+CDrgEoFgMJrsGGF2MFL30rDmP6QrtN/RXILDRVjWlh/lgIWFZxqPKzLt
g6bSH8hyqsBjF2rr6yrgPJKr2u741/r8xVznGb+npwbaSfY2EskZve/nawoEJ++5
1RiEc1peTQbjMu7kRuEkYHzzyU3xVnqw8ljCfpUttMTG/ymK1VM0eDI6TIJCSPaS
RJ7ZQP9NY2chdW+OQx3i7rQuoQkH6qUUXDA3XYezk+B6EiaWTRh43tssSPOkCr5G
ZVLffITxV/fy7+wiVGwGTsQrILVSXuK3+//+7xRFumcjXJaXLVBMmln8OngAeSXx
dM1KASYZ0bKVhMc4vURV0LIhGKHTppmiE3WuSFgYhy5owUfL3NrKy1ZdgkVaqQRA
58ex/BnJK+wGB7zKqU9ou9ngcR4+a3sDxJjWw0Vsgxy8xm/Bh/jtuSea1zSMZf1+
Dx9njtZTODiQOpTsTxGTgt1k7mZcU4ySgW6hYu4p7Ide2CpQu6klKMwtK5XyYn1L
iP5Ej1ggj1fKDt9a26nKTUE7NfHWVoqsxuTDPxB6SQMRQYvamV7QAZ83FQ4hPf58
K7XmRscw3cQAh5qVxWpWv7qmLjnn77PiT6xXhEE3fFwdd51qZNJoDVAlk1H4i74L
dhT0XOJaBNstKgohv11OlFjhSx8VfYnpOriwWe+upFlmZIY+GtaZW+SnHQomynCl
931644l74AYWwNNtqxnNiWQslg57kve5aK+SgY0Z6f3fvn+O5ZWNnq4wi/MF4/x4
ZB6UU9ctjFe4EaqXXgULWsd09qvsIhncFeHxMbHEe/WuvUm1PiLcRwf4UCTZkrj7
VN7ZpJkRnSKIvtEJ3iM9l9YvauDmle3Z+WCq//yda92rj+cC7w80fUe0BpiqdKlK
UDAkY/3lICzSNrWaVwSOpn6QEX2+05JdKi9KHluAZpJWwgjyZDGvbR6Vf5rJ3G73
8XOKmO2XSQqUYTUWBZnHTriVaTfy48Tqg6WVvwZmptTQV8TBfjKKrugq4Lw4G3RO
zlc5lksZLYEw3u7BwqT7xOMk4N3wOsuX6JxTipRLPg8K2HWN/khP3o5oMNWqifch
n4jn229bi8++M41OFcEUhJ4vikUfWtL4FHezGCF4O+DhcFCCTwX5gUHkfTzIrruT
CBHHF2jqa5rTi0JB6CRJ0DTjLhIGRTSyc5ScU4CYj7i0300Qn33NR/De6N5TAkRh
yIetrdjG188JWYU5oB/HdK6sb7HOJzceYrSIKoNdBKQAPSzUrn8LvXXo5p/sYhTY
xaD4F/JZUOcIsF6QqO1JBTYI6tdph2flhYw+mwpIqX8zQN8vW/Tzt6LCzFjYgVWH
bGgd0dwYwkTcqFJWtVruAhidtEhhZgL6zxHkR4errx4aOv6m76jbEclfktqFH9oj
3O9bKdlYs3vrETIn2eo7Af6saxmOK+gEtGdh8wwqD5a2I91fG1IY8bXfnkB9oQmD
iaFhrbba/IbyUGlDHVJh33dzwx5LY+FrnrBR7YExrcrfAJ16NOnThxZFZ2Kw/V1I
hVBUORWhVdi4DUsm/iA1bFOOt1zmZrJOelxUZ5gqdI1JE/k5urePzy6KOR0oZMov
Ur7RmygmDIYD80CpBH8RJnNWAdSiHB19/U658oLfWl+uP4bSAnyU4iHB+lXtOkc3
cbOhkwyInaDZiC35s5s5516u/Qh0r2Xx5JAbtX/wNA5ageCnlxtFKWykXOGFRQgX
UEEtDeo7eAdGCo7p0jWuhNHl0DFWy6AbJveX9uASgRbBIaUKtT8XNxK7vAiNKAwE
v4OBrjp+H07bHVwyZbgJ34p4PUuATUZ3HxAcdMStdB1EnTCee7T2JFVJfycd8Kk5
9MD0LBUeo860QMfCuhz9Kx40fKUxbsmHBEJJW9c7gMB+Ejy//5W26R0DNEt1ENkl
62UnV9XkRRLxX3dzQmX8ynWDgaTnh1x4JpgpTLlbaQFkS5iITAMpblYIhF4wAubY
23fpbj9UqW9H8IOmTga4q9R1HukWKl1M2cGdTKNwWEoO+geex61ciAhXhW57i7Fo
JxBW//F5HxQllMvj4pZoVRW8qe/s7YBvBL1l9/DYW1FxIXLX6gq8G4edDhKv35hv
HuWuZZtTz+Vop6QMQRESg+/7kmWl6i7O48SzmeDj2AarWOioKFqWFySN1fIYWIIv
OfKFri583FZOgtweEJNQxw6X9cSGejKK18ojMlo3zikre+Cs8cSzo4d9FkPCrJBu
ssjtYeFpMbWTe3CIGzAloFLFAm0OtxwD6mh5u3cbmCJtuIMWAH6M1ZsMGGG57gVy
RYaq/KkbjWR20YOQAhi8KTxntpjkwd+2q3FuJOed7lz5GPUhB86msFam1cS0/e/q
rR7XM+bWtHZFFA8VFloS4Cxw4nPY82Yf5hFILiJlkOsaGftI99CZzBIA/IN0uO/9
yOeFza+PAEnQOMJVxEFgDf/b1oZtyvVzxMiAa4hwjhF6H8AHutSUVjRW4RnZGb5R
SbmJi9cZsbMqMzgxGeq9qUBs6/7lULi/ITSxnHwjaieGabOyxNSAQAmQdlN30DQq
aAvKJ+0hseFJqg9LesH5A/+M1PV14oamfIfe2jfAQ5N+DhJsYPf7V/6kI4coc178
JhdeFfxgT6LO8ftzQajrljocAYPAkVUJbnYPe6dRgKOWc/Mf3YWSA8jVcJlDyO4p
VixzTBIg1Z5W6R+qGGYeDJCSMQGMkruGO0cGll6UAhNYmjrQ1ZV7xXhvFkUy477Y
Yn6oXHBHhic6xSER3nl2GW7tzdtBdmJYTe2UriMokJTqE+uVOfVVHRVe+wDBHfT9
Llkxr/XVSkTfF1mXnqgWgaPLPFkr/VVhlbbQCkKc7M37oLi+W1Puy2aouRUgnt/u
8ZoKe0oDnzuxCjRZBiJXNrvlQkWhAqrBNDDMP5SB7YBe2JPTT6dNcR7aU68Jbzyj
OMsqgbUEtH3GCN66+OWT4n+gUQXX5gqSW9j9KwjtARZocm9Vo+RfJb73npqSvAyi
487XFW0miHHFeSe8E1W4//Y+VAzFeTur9ozfljYoOt1DqyFqvb3AJ5UthvGkGTne
LlcnQnMCraTWw8zqrANDSbFdRcH72bfrVfwD1IX7JTM1Rt0AI+ZZPEUygS+Qz20q
YV1lxkCRrbtuHzqEr6Atwt8IgPq30Qx2eJwNlQyUAEDr9zjJjTu/Bxec9C+nGoUI
HYL3pxfLMqN4X+54WDDbOQxwrT5dVXPFCNixSRTzL/WKqP0wyokLKfh/xMAt6co1
Vc1WQWP9x9Z9hNAiVne+YUmLXDzwFAd+1RQnPkldPkIlhdcIlmqPFZ7X+wEP1F7g
QzZkKrb2adxR6JzcDjXkCkhe+eLLSiC0ocJYKcv5yLkwsfdAGDeQrjy57jsog7kl
6FVbUINUpwJ9uyJKRvSyCJSgNxG3Cp7WIjCY+7ovl2SaahncJs7hkBXZzj77kfPP
vAUjs9+Sq9gYQ1l2yxmbDVT5ZfcA5Uf+WHpW4omm9uFSM+PNpCxcnapOf4i39hHj
B8p7mXcHiTibGv/FN4bi1hhCqLkDVumL6PK8R6Kp3JtYoZq19doNJhIy7joTIk6f
xU8piRsLcoZv+cnlPQBkfMjNvkuxXbbpqKiAtGghHkFpF9uWwjuGr0LfF0Vy2P8x
IhjAWJYZOPzkSt5+0FCxYRf3JRP4kz2wEaQaKNTpXxSrLfNq4/TxB5mQKk5oH6x0
NrKUSznc2VTmhNgmW8NOWObtqdLyg99dc2RaLKDA1Y8xqD35L925f3t7G3FwQNLa
JYlcE8AS1AxN9HF2TSIe2eRz6SKvdnWahMc+CrNX11g55B6wiOIpRFiVOPeBSDpH
1flcMJWTmfTujbWzoQQ9z6Od0XxYLzFllg/BXMBApTv93ElausjnG9Fmzr0PuO9R
BY25xvkckzuI+Ym3VsIIP44bMDcVUUmM2TzmKwE3Z9TD5YiPPCcBp9kbtfA2e/bk
Yu6kanZ38DknSHvKwjQusuT/OZ5cpxt68ybWao0U/dpRNVDKhBc6+0h5MJD23C+y
ZZxDe+lwXaudESv1rLeQmwCK9hUWG/g3hNWr70flbBMSopMEFdNAJPHgXePFUF9j
Q6qjfp1XW4I/AM/8aMSA968gydBrqZjpF6Kt0nQmNnbVyQLyXjHEvmF5c4n0o57L
+om6Zsy/UmI1UMHSmNkSulRzxvgStkHhJRmRal7da+yMQcyeL1OGejxRz0MJ9n6O
lkbginTNDZoJkeI80XrWF/WsyHJU7YrgF/S6GVakKTFo1B/maUkG9tM4svZBysjv
UcHheJ0QajsXxm7OT4D89DO9d9+aQDLMZBRHVmnO3YI3uRQDHr6xsHl9Bv4oqsMd
IBdjWMldBM5oyrPPC1EHZ7qaOjVqlGFYdgsRLzDpSOz0+iT+Ez8ohkoHmK5nnI3C
y1rtzpm3fafcxqW01atvAWDnlLktzy5U1ADY+cOEdSP6zhxaQKlLcxqbH50/9rOR
HE0G61DwZsgrU2JqtpfIZCjkgqa0KeKFH3VtnGNct0HKej03pAfEimUXrB5gu+E9
8+N8Z1dcii8wPDGuiGHLjYBqZbiaJVOdSInp4+dMracS0aBDg2dYC0gILvNV24K6
q+NgeNuOXq4NTneIT2dYlSo/1FD6CdgLFBR0esIbZhW1fkH3y0ffodskKhsEDkUS
Te3glG/BfvDFBpiohyzYKfIdATSwvl+37U9HSyCGCu/Gv1z4EkBPi4IK92Lei4jk
Zapxp1dBST1IHtHPQmqvhvxf4xiNjL0uiLvMA0F7jMkJEFcLrL3a/tayT0IpaA7R
yfBaqvuH6U61jo/5Gnlfm1pugvEGFRKG3aIaluUg7o2zS6OfGnUck5gQBNQy9i11
BvCCuOAKdJ+qt4HxQG4OCXc1Z8S121QRxAsgt87xbQKfQK/FeOwQ2y4ND0nedHXW
2rY4e1IH4QMDMjMK6XACW/IYF78cjThLhFC9QBaI6yjZX+NSQnPWtMEQdoiKopM1
vGxTpLznGuAmH3RXGNUu/BS4HXMOra6IuzRgO5jpGnb42j6qTv8KVoEWjremofFb
zRNcf3UfBB8mLnhQyqi9HcNUP23sqfBKP9akl48FscUAzSuxTN+Xg9sPT0h1IMqy
yxkKUesfhpe46ThbXcZwjeXIsaBm+6EFkls+2Cm7Yl5arw7aereOG932Z0EFCq8I
yD8Hv9quDMImGHrtFa6Hev9WzXJGij9Z5tKinOq8dnTZX/+CNznxa9Ns8k7Uztn2
jkgjE6n7w7yiv8WelPEu7eY7wRgkLVsxorsc/Enwg9dvUYR29VK52dJWrKV0UbrY
ZZ6vl6EeGudCYGFMhryf4g+dcrB73Jl0vGOOvOl0S1VRd9jHAx5GhxGqA7KK7vIN
+olQm3BkusT7iX7euCE+EyJd9h1LM0pANiGjoVQvo62zOriqZ4qWhMAFsRSNAsn8
W2u3oHaGdEj+LZ6qEYSMdGXWfRJVromkOb2YOMAxZBiqh0ZIjs0mvwxbiYwzFoos
o0jtaBO9DhDHbairFoqZ8M8V/salcDh71/J5aD3NjQZL5ka85XyCi1aUmWDk1t9v
ST7QonaxCiQ08Gi8q6uN4j09eQzcqbQnbWPXF0/wBK9A1cAw+RSSx6j+fDyZFLVl
HP2E6dPRDddl/Yy4pzBS5CQg+IB1UXFn/eqeJbSA35MAcYtz5sfadOecJWs80iOq
z49xjziYwSrsVB2LUYAQpgXBwxrQWnI0X6+XaT9uNDa3eY8vTOFTxXUQ3auqstpf
dVIE/G4KGOsG7jbYE5L7nlt4gL+u3FWzsSBt25j5eA0Xxtmch6kVZfjRVvVLULxx
TZHDcEkyPxUi4GnO3K1f/7l6RssGk/tGodMang/0/ZAg4dlzMDzjcxR6JTUx34FX
UuNQqnhtLb6Hg9SyN1rNNC9h/s1Xz14/ZxsSE1AP4dkhPlvTvfnoEkTGYRFtdQtJ
QcZrWbDaeG7RsYgsa5GUiSdZr8/YUcJvcOk7l/zwwGALz8MmaFAlxSmLkhT9AzlE
AS5hQoybnPsg8ZbgSQMhxUNL9y27xxuSJpbw4j9K4h/sF921bQqX/VWWtD8REeY2
xxprznSsVdmh55TaEYck7ZIpQ+jEnjDp34dO9b5NpJg924XHWWzGnsIkpQSI/CUt
QqC4FkXX9RXdji5EBPLIHhqddNgMC00IVATXoytoJZpDfoZrReTTsXCRTMDkIGe2
gjpGg5lKJNbZMj23boSSHwr1rfAGJF9v1zKmGLLYFMfSnV0kDQhqDyNDrSQ+SniW
D/t6hu/eKqxjw1z5IXunJ6xHFHbEH1VEIjdzDzdMJ2dAkEF+3aiQYzpoMSDtDvPD
vPtrVLEIBVYhW5kXwzcihHZzNta0LYOcbp2w26JJiyPRCcYBAqeLvNnuxQi/SKuI
y3bUC9KFU4MXYu/gC4m5XDvz3RvVThGEwltJwd2YIFY8g0EIGmi+zBnLrs3n5cT/
ekOw/Y7O73JHXFywZQYagaP+ADso54GP13swB7w/cF1FkTphKbVJYc6b97eshMWy
KVj7eFqJmt4qY26pjwZ/FgBP4Ys3mSHU1aN56wta2Cm/8ff9tlUbQHoJ+4vwPunT
ke9AGyMvkVXfdhU05l4177c/fg4AmlT/DAtK6j9C2fUXEzSn2fVi8ZXz9z+tZTzA
gLZX5PGOlvxaL92F4vwuShJ+cCprpqzDYTUOMXTGgKwSHh5VhnARP+pL5sCIJ7/A
9eHZdbXgHWFyUAVhPXcoa/73zrmTr7W5rWY4u5NEb/slSyA6/U58zHYjzIeRzdk2
xN2Dip6dNt/RZVvAtlnYzKN+1x+dfFAc0BB4zPnbH8AoJqloBQ7tVaG7/mZEHadm
PZDkrby/ATTc+F6qs67X9Kt/S+cd6QnBrsp68bJRdHbnFxjX53nc1YgQsDnXhCgB
XMU+YY+uQ4d3wEa34NToyWGxevc+5bi7N+YD+qELt/VcjWlzluRC0wbS8JrmC09g
cTmYomYJQjQYfCBfwiy9OAosXXoy3t6fpWju8L53Oo0rWLIx3Hvb3pywtJ11k0tJ
XWb3q6o3++/SmYmLvifSoV0R8/ZEorDjCxu0InxWZQ33+gto3zmPQfNfmQHmJNFY
swzLV2f0G/jnBdblU8tjLa57wiVBzb6zz3rHQZu6o0VY5uWCOEM1gfTJ3iJVzFY9
UrbbZ1Fva+igVTMMa+2QHaydA7wT9KJ0ki/7kP/tTaeAZp2UFA0rbQdVTXEu+Tna
DH8knrVoBT5LKwmk2vQ5vtKQIZ8U/prJWvh62ibR/4L8SbjicrZThQeyfykklUMT
6iSBzf70EHU0fvcscmjBzUgMHByzXO1KXlctXwO6GHS6A9HhpjfYytLUxy4EivqS
PfOkKdTLh+ovZK8hIrSg/XJ9OxUS0LdSUG91gkEcpao+X1TUPt3a//jHNiu35701
nyJV8QU/DaGlQR8FnBHw26cDY2xS1uBQIluveJiQBRrKNUJ9+61yTDnvz4k6fLaK
G9MgQ0qzR889bZbOrfxW+ijGIUCnQOAZ4Lz7cAwRfRjdQmo2heUQhs7vdXhOMROQ
BS5Cn9NBQG2yofaklNk/+N1zCrRNcFJKMPrDEJIUFBoGacXZaccUVAlyiBu5hkGm
qev98/TCoP9nbQlHihoZ4kOHtaotSrbAG4BqQFkFFIzTUAr0V+nAn7ber7vmcRx8
xixPt3APSQA92XSOvZYwfC6StLypCoU3MxE7oS8xNdp8IF2KSaaCW97NIMiZVkQo
dyqJmxnCl/hCaV1pkMf8nDcsGrdAJwW3pUjzsNnMaRrgFJ42TafonbGjH4GxicAw
LastF/OHo3Dq68leLXn6GN3pEtloMLNVXWcaKNPv6+1K1x4Wns6zcoQ7OdrID5YE
20tYH6ufEXOoGmEJiav9W1ZtppBKppD+ZX7Rs14Hf5QKoGKz5E8HX855G6926aR7
R0ebV0+C9NgP2DyItqq/qf6soezcVG8oFYJ0Uti144VrGe18n5HB2sA1/te7dcEd
UHhdO++SUSvifXC30fdoFNFEDubqTB8d/+gD6ATvUOEi0CTwqLFrJlRY+k26OgHv
rgeF7aeY0ShlZZmVmpOveBB5u8hUUkalyEd3QZTV96ArTJO1PkDmKrLHr4Wxf4La
74brDXIpqTg1kfq7qd4tBXvBsiJZQSodS8awk+O4//K6rf0gSsWFuCJy+Mdw2AMu
Sk5nzjzZpoevIe4gRvnptmBcHEUs8cYPb3JykJt7FDwVWHnz06gaiIGvLWqqwR8U
yHsDVwn48zNMcFUKDhD+OaxSRrHpN/A3QAgNXx2RwvxbfFOEtzDdjXrVlFLhh3Rc
vKSLipucUDtsN+FTmo7u6cFa38ulgfoUoJftNv8YXo4pp9blJ/a+TFivhBwv4XO2
920V4zdPT/X7H9lq+7csJsDIgp1evA3Uchs8Jpbv6eyoxJ9Zb208AB7NREHyfLKC
rzLp7p09FponS//XHRAAfE6282qxjAd4T1rj0XduOW7VarKizv0SPyyqPf8JSavU
2TbPfy7kFv/stC8H+tuQbTYkdSki7BaE4R6KVo/xU4WrpbYHAmffq9gfdHP9fB0J
QY7jF79Tc8i0wqA5+DLZNovhQyzdhA/rrU49b8m8Tu4wnUw1pk8mZweg98GQUcRu
2bc/oJTBas8VptvuwayD0TKhGwYK4xcnxlHjTDKtZ9frxLzFw85B0ZCYC8dMlWRe
w6elz2Cuk4IAUOW7/9Orj4ijX0m7Wa17B65pc5xAllD/Iav+vCw8QPwyfIr4G2t2
xs1LForzmgOFGW1fHYN7FnzmKQIzvW+MmMaS25lfXbPNlI8Lg+S2xNN2yE3/lzR2
unm5TJ0dXSzwg87HtcmS7VrzHczwZBRIRzsyAKjlGish5AqMgKJGoOrCzwaWxLO+
4jQe07zH7ZtZmhToGt6Ge01doL4ZQ/DxOIDeU5J9yenVT4RX/vkf3nx2k3E36AmI
PEZFsMAAoLwABIoVOBh2m6lM8DHpmctr9Ehsp46Q7e8PNdEHC78RIdKyvwlths5h
o2XIddYiW9tTufC/4APoq1B3KSWY0Gl1tQvK28eA790t2z/M+gsnMNe7lCPi3JMU
hwUKplIflWGD9BE6XS+MgjNclsFLLrVf+ZFfTHJ6A/s/6WaLcZ0UxHtFfCmStca0
FqnVxqPkms2qhvqR1DGgJtA6qy6ljwBxC5hRkfEuzWg9xxUtS1cwxQBPKpCNuCrg
22rwfdTGgnh703aa9P8rzuBOrjG4gt5rNf126pWk4ydTdm7OhN7tAhBwWE69R1+x
2qF4iQPZcAt+ZfjAw3DMJDLXyA/M/kBuSPKrSPrNQw/3QCBYTAdY6TOIrMM1sa/5
ZSOcw3wQ1cQNOWdrAHJt3wA1FgS9BFNOld2EesPf/FSCBzNkHgag5vMUCX7/lDbI
6lSXoDQT7NLBcNfwybVs6/498xfk6DP0y4YiKQ5vonadXN6V0drjKEaJpUyqDXjx
fXjBzTDqhFIASm47ZQFaJu3x3c9ZR0WOPLJqXEpZ6BDZrLB28jN1EzTeTVp0wahj
3E3OgixF5mFrDV8hmxcAoKz1Lrq/UVUGgzafzGKutHE1Hwk6zyWwHXjPKLldVgdq
/baODESdVp9TGH+JHozCiO9unWIhPO5tgXCr/X7XUJM3gCM41kT7Cgzva9cE2Q1r
6q8H7a5mDVlIpsLOxAxibItAez4iJfCQg3Hk8loIR7jXCKptIOe7owd1FXzDi+2Q
B+8preTr3OZC4EVe4D41k0ff20+7lxDWugeuxCouOdmgKrUmX57nl50v7qC9B5Hk
6OwlKAzC/70KQLveabFp3lugWmxbMgZPSTdccYXY3oW7NlE5PahNdNl4xkZYgw2/
j79XC0Li9SAZNhDR0Gogk4M7NBSQntbFClhtyele/RJIzl4+iWGo2DA7zECHiqyB
L1ESCx+q5LxBGrGp+ESWhaFyHg4721AYEhwi4VwQBD8Tpr5vUeuUmNrV9iOnxb+T
QQMtiKvwyODkhgUo31TRV2u6AAuoDV9RNTqIAwYKpQpbNdKqkdNdNuvAH2NNXikg
D5ZaWQyalSCDbZZTIg6sXSdQ5YFSqxOX3rndFHCbr34uJ2T0PS24ZGkpgV/yBvMO
gPehNtAsZLgn8+FXeKLnlP14TCxwEkbSw/8uEQoHgI2SU3lroJrhEubzMAJfnSPM
JF4O3DCuGDvcCb0oUl4vMmBKd584MIuNJ2kmiu1ebfO7BJET6FH9RMNqixhpwwyk
xS3gCoO2/McKj+fMx6ePG1KyR7XvzW103uVUAzzYxT6U4aC7lDYJ/aFPUkZCbjb6
wKtzPTyMPHCJPeSnCX5aK0bQYmolbAN+lpUPs2QXiD+Qs0aEMqEWU941YS7IioxV
v1/cJXRQT8PCGXfVUMBaRR0YILl2EIqbGFdlEJBBoZogQK+/05x3HNfvJWIhUb1+
YdKbTIMwtiuQolKJv2FHhaCTJvqLITzCS9Msv5EwmWhbJ53QRfHq/r2osmmQWj/2
YXdma8hdEQDgKH4BG+c+4dZthqkPE/UfHHpOBgaj2L/ck6Efsg06d3itB5+k8jZ1
l/+mRj/SUA7rEkqbslgcaCNHM+s8/Fr9urPs5RnFQ9ONJDZNkveK8FYake7yVXkE
pMmh71B/AvZtelovxFFLGT68+NYHWeCvHlLqCQbfjpPVI7ZVZHXsTGy6c2LgkiYG
kCo2OSHO1btonJsyvTlwzUw16XZv793OIieiRTsDk8PikWCElUyAXD9oF4X+INUn
6GZWL6jAVJ43lmql9fOTcJ2ry9NxDG8RmGHWxP80pteYY6YtP3haP/Iar4K6gh66
JoHwni3HE7rcIODNBIEvsCFbGw+4A8v5zx/oSIgF+zNbf7fnaoyHlAWS6DcUCHe3
+YmzXlca/JiQfHbAZIBF09jkbLOXjnjx9GWj5xJEynKQHYk9dL5fsJitGuimuxZv
g5S8BWZ9qZl9wM6EgDTWmQTnZyRvhjN+cgVu/pb7AhuSbEZ1TT+R5dU7bQ4jsyvR
Wq2F60Qz75zfGMT2qMpu7UW5vc7USr8E1514b+ZTh1OkvqRLCv7BumGflnnCcewa
8htj3WSEKXGK0Oiy8V37/sjDiG9mzpnSniRnqNI1tV4Z4Na+tBuBlqrhx2uLsBEU
pHGfe+8rlSddHTueFps1WjmONGm8nhL/npII1ruMniVeP6oOdUSEJ2e+XzeNwmpL
l2YRaH5h74CJgeCu6iBi85LY5UPFRnGiBMUbWZ8KKWTtsi7bFukD85/JD52d5/81
uWsWMCGtir553XSrnvnJUw6Yvg0+JaiPtDqjNyUytGvvrOxg0UVJIxAcmq8u3zG2
FqPZ1AN6J0WLhrC3916uyTwNQesKF5Ds8FJA2hu3+dS30S+c0vSBjZHU3zpjzhcQ
Nge9W9Jy0+IqA/UBb8vjB0b99CY4/XMLi4ijKlonZyFVCmVVKCHrN9r087B/Qqm3
VpJ5ZzG1ItAXIdEVGYH2EWfQW1V1TNh0kq3IUbiYeOl6nNL9qttzyntDfFMgnjRs
ESPWhy00OsrHhDfypYuhgY34sF1XKONdFW7R7014d5k9jPN5KHrOIvkyxFsRQW9j
4WN5kYBKb8sUDre4OyCqdT590Qjs3OtQjHbJ4BlH1eW7cMThWSvv1ETE/gnR5K4P
YV1N+xsdX8rZLooEfWZk2JsfS9Cgv1vFMckJe9ySW/hjMPWOhsXqvayGLBqQ123s
dXI6H2hVI6hyBB1JOxY1BPuop+xBNJl2VRTABjXfkVHUxYKIUpGesbSYTmZxS+ak
aMWPqMFes3eLsnKmgE6ek7Zb5X5Ocw8j7lvGxlBaBWuHpJfFi3RBWxSc4gYKwoKx
wsVAUbHxfgBmFiv7Rw1HEiDEfpbf+xkdRsJFwQRDP475ot+Xz2jnAsGSvj0Q+egn
UNHbM2NeFSz7vOxF+p50XMSaSqo92s/oQGN7oM4TXKgVxRS9YP1QqWjEdjMRS1t4
4N1itvO19e9NDIy5PZr1SN0o33ilc8CniiT019lScPZ1OJ37FzPYLmzR95RPs7zw
FdLAxjl3RvKXPV4KkayuptqqltXRYU6KWP6reEjwtkAmFub4NLbEjDBcT+2NkaFX
2Wg8AatgoH+EQIrwxXBJrdJlzp6W3Y23FAprdNsDPXVndLripCoYx5aJMKYK8Sd5
/UBAE3w4rlMfk+2VZASRnygIR4FNA7+rB97+4E0mdgWVda8oMWJenPyAeo017DYF
vK99Mq+O/nSjgtJzO8LZJb/W8nY766ZwfAqKrUFNUasesgZDS+2gBEWc9YxovHNE
MgSfOnyhvAb/t/6EOmptGszdoDE1PddyKkmv11philRbHlT44hkgxgnfaFSHlpXV
9Nw0Ojv+U9pEww0PkejCLyIuXPGUr4AIshPktuTr3kTMRRxXhIBJGi+QHYxzY4Ux
qMPVZZSj3klxHpzhH310ad9dhwRp0QeSwd31b02MqfypOzqQXxM/Q6jk4EmPbs9q
TvomZxoF7Cvg5xIwVVPLG5s5ceRm560pNpS3hZOxsusQMcFYa3FM07Tk9zjFwkH5
2r/w5Fxpm/Ix7wRb8zLfD0HKyidpFPsUinsTupkCd9Gp2uvihKcyRGiWDALKIPo+
ExXgRDFYrhxl/eFZ5kayRlKV7Uwmv0F0uGSKP+xITgJkECFOga99y6C8TJk3Md0A
CkjQPkyqYJErb39yQXTisxat3UP9yBAv77VdXo9jfHPXns7AE/7No0IQqJIxcBaP
rz3yvILx3i+R7VqLvop5H+2mWfHu7rK0qhJCN04tg/4EJsqMmwjjugsPo4Qm6e1C
sH1hEJZcrIEhQkZLD2xLJfTutRwdtTMNvsPypr6xnWx3AEahso0pUuKTJRKGXgHU
O2qdvrvMF/GlbuWmh9O9gQ03h86GxriMVm5HybgXYRfHO+9JhaEBFbPYAI/hgMLN
d5k/CHk9LvY0EPfHn5jWnivwodc3gQAhgCan4nQ5b7vPQyucjd8Tl+vOZS0xKm9B
JDgOQEWaCwo2uNkJ+ra5xmAI6ES1+lt7SnDp1lR3iqUC0zIqrO8S6W0itty28gTc
IwYpVrlkyfisKQrcz2TaQJIb4B7P37CCrYFtYgiQf6TkQJyc9CICpfotpgA0aNia
+NFRG08EvmbNTP7EZ0X6uQu3iEeNkcbxrYlqBg7ABbCBF8RxURF3RcZeB282nGUj
dQ7+w50P1WGeiGwZ6TkD1sMtEhyeU+CA+d4aHViXYiOP9AQLXxz85PD02cS2FeJK
rUs/6MWkyMXYm9BF0bogG3+rO8amV70kinTI5RpJ/vr4wdrF/zsmNddtViQnqoEE
TOWUUap4REg3H6WkAYpK/DMzDmkglQeHeVYHxNPn8IgeCkaiXIK/ywjOF5EaKm5R
mO7w19TxPQmHsWKLwQRxiFc/QAA1Orz4Z2lNHDEBdwYPmuJjyudYL33aJc38INFg
WPDa5rIRw5Y7cxwY9DJN1NLMeBIV2eGXVDYyrNQOPbMoQlZtgkIsfBKMHe9CYlT6
6vZF1w97TVKWYicdkZ1tfluhiWxXYYD8x/OR/DMSHdAOh2/5oM5LqgwJCfCYPENR
8qcHy5pfI7FL7w/pVDnUxNZYieoijm6UMPI+KUTZ5nou9hKqBFiQQYuIowPQ9BML
94F9nyFH4/6ZNC465H/2Rj0/K6+QQH1vUGQjCyzZQQh3yd3qXXn6EnO68HFScnw7
cn6sjQ+Xn8gGDFs2iplZnKNQ3qaXCPLMlJ4hbEZ7eWxC4O5DQnuclRVvEAHznA3t
AJ+Oz6qzIuSGJvj5HojE7tAeGPQ7VKv92Pgr/gcd0q9qrOrIiZI1kxEEy0ssvYm9
CTi1maOdVKKNPMoJR8AUhGkphEqDaQn0IheLu1jkSLOHLJ8NLo5gFLjKRCd74M8F
okckTWx3B9hWdwxbCNaUoSZA/36eAzCG32eGV/kNABeaYbAvuswo9ZTDFb63m68y
r76QCdd2Anur3+rlaprktiIk+FGSS6AU3fbs3oFZjwhEufL7dtAca5HTugMQ8v0f
mwoeuWBKlJouimj2Tyz5p+jXXBs6z7OP32ua7f6GaHn6lGAkoo4LMFZT2nArrzmx
KTf3XOdZdLooedMI8F7apJJlud0UnikvlT01bnNdCAz4XbyC/pxBnqroE49dndxh
MlaYes1GS3SbXERQQRtewXLClIMR3miznuvZ9XTBtL3auCj+sOjvWDpwR3ACzsCp
2Zken53aHeY+FHwx4HZQyGJtiLLwFDq83RsR9IZTkqPz8exvIusPRjdk/VNql2Et
9hVFt4wNYMrGtJv6Xc87uWl83rLIXYB5+grINmg7AduJ/dCKJo5xKHS8oZ8ug8Dv
TL/mw2tAAbVFticgYaIEMYXKN+i6rJOhFkYT1TombPGI1PCaV/1RO7p9BdFqyolZ
/OGzl+YchR3hhY+bxlre86iUURR7Mo9ENsU5a9x/Z+oYcaPTQe/1FQjfW5DeFpVY
ZRaP9IyE9QkjDTB3R2YJyURFhwS7nGcB+YVpfzpOXJ/0Qj/753QbdcOGagrzH+Dr
khpNQoJPGt16GX7k9AK3fOGTIXJMeHq6Hpc55AzeMYE6ciIrB350KrVDBnX+nxvP
LCEymzjrrJi+LDVvvXXpumASLeIgeG9KmC8xgQCXHW1IKl1pMFCmtWdRLSLyuHm8
fdG02qzFx3bJhBaNv3tPu3G23ScAo4VpB5OOcj6ensNr5LbFgBfM4w1WTtyuRmKE
kPy2QYis61RAjE2hTRhSedNjruXdA5bu/Ch3hu8VZ3NVSjxPhYLxhh4JJmY/rNr/
VE/NLZX+Z/x7O2RPK91w2OZSsqe/bV2RNX2hniO2yPkI5LjfiG3uNoUZB5Dwf0Lt
y61ccw315L7gQWS6njFYvQfOua9j80tnCawhq//11GpaIp6mOJLedmxw3EiihWbe
UHUtqc67+oW/7kXzydCE1TJti7VzSj2wkgY6Wb5OxSR9BfR5Qqzbl1S7NnImvCKg
5g9QH41SnbQK2XUdpl7Kg8aBv0fR0nyLk1qBGPXsZ+hG0KYeKabKPxElx7xXYe96
ycHw7oP7WEJlqlxs3uu6FZL7CRJI8NlCrS+XCs4T8l3+fR+KKw1sDzU3ERmAwUTz
UF0Htn7Ltwc85sWsw7qKROkbKbTPtEbOWyN90whnYPOnxNJq8XGcCCu2SIWEJcKj
s6U7bC/cVc1DFTBpO1onQrSlFRxVj/8d6OhEFql+JVR2xpf7sajzshQVgySVHKDx
bAM4m2o5kY3BCRM2mfgCpQ6sLouVYc+9xr7lxWytHak5bQ3sCaHuk3n3QYwuvADQ
4xKm/miItK+V7mJUJkaSyfmAhQ/U6pPKxCXkdgpdNC1QiQIqO/2eR/7efqdTTTgP
o3rX+ofxT+vT3Vwko39AKGkhgicQSMo1I9qzqztgAl4ERZNGvxpZHGRCRqZC2j+x
ykZTqgCd0RP9W+SRxs/pjw1W7hXg0BQ/NESs2MJ1j9owCST/fd+Cwt43dDSb/SMV
XRzVbRpQA1fGZtQaxX4e4tX4boqE+ThykoKk1f/Gu4NPNN4GA39g3qo06UCdA1dm
uhBZxSoTdPNxylS45VXcYrR3bw0C+P1G3tlDtTfvAQReAbqM8p+jRPfrPw49csHs
3T9j/5HNJq/afU2RUaJRX6koRpKrNFE9drUX/UYYitPhHbDaEUxmAKsfR3EACNBx
/N/CeNsKmhNWxTnNH6Kd8FJlmMZINRNjnsbYkcfqR6UybJCyj/OxgtsclocOg6QT
Xg//IOX8PhYaK3nLiT/fgZHi14RBjCUT2xFykg/Kiw3kJcKLlpxNsnp6+QqLxpSj
SNbEbbZ9Gf997IgSe0D0aSGtYPHgGG1k5KfoMw/UnYKJ9fgpiQW1yXe3wZNTfg4z
PJpsH2kraAMOVR3uSNUDF5N1ld2aOe39AIZ5xLM+f/ebNP6Ji5h3dFuAXOp2ejy6
bpf2y8plW2SlHFqQdx+JOylUwspBMxciQPheswscGef1EN1aEuMiRQBVKOORQD48
ReytOnaZTq+92tmpRy6POBCtvD5JZdG5j0m/8+Y00d36iIro4X3rkMmfG7PWu1qn
UmyvqPJMMH0ZUoJXbVLUx5lPtj3F9PeY4wt+A+ft9+kbusy+3rvYtuZmmhXjBxEC
UADwa/KAXEB9scNw8VgD69iq6tnyGCpuDDZMwwCalMNKc0EZqRkKlVJ8+hpb/dk0
ro+CiNKnxTm7xHW8+tndFNO4lbC41p82R69razfBbPPPfwAaDNSyWuRSu21LPTBh
V1eZyu7ijmkc+8RASOKbfqyTatn3AYpXtFrlJatZH7tDtVz9Kjd2mohkvnaxQYQF
NqLzNe8Gxj99+2fh9xiDpRc2K7DoRhdFNQ5kjm8xarF3rm3pe8bc/WVma9d9rx2m
8qNJWlPTW01TxkkTMpwee7JjLDvppZcMKRvi32aFK/POHjojt+TavOb9QBnCJsvT
uGRV5p5O/GsVE7ujGO+jSol9CpdK5w66IVBEYIRygfL6yU1eCPg4mkB2UtV6pfIl
ITguivImfPpGPP4sVPpR1iqeqnSEG/vAlqfFcFEeEQSis1xOkim0iCqbRz/ibLyz
fRISfPeYt6DdFQIL6yZPprx0xyB2Mdp7iTDtcr8/WvufpW0SUTHJMpGkX+Q99YZp
ZcHPmWi9w/ZOA5Q6BQ35GqGz89I2QcjAio5a4EBMDEs29ulYzZTjNq71eaXC8tcb
1d13HdL8OWsWpKFWZb+yCyFCWF2idwvwGCmXAMEUnTexLhDHNFlBYCI+fHbJCpS/
g9ZmNNQoTRo6zMpgLz6NNM1/rrwwXOv/8x2np7v/k7ZTNr8fVz8uGK68XzeAFiYn
JTqO/p7JodtHbzk+f/DlJYwl93aEUgK9Zsa6JBsQTGngD38YbvsJuU/WqACT2ALn
d+We27yQwadmC5P2kWW0ZIR8N50FOyWVnpOWy4LOtF491wU7xcTePj0U1CF0/xPy
Udfr4DGa67Ll3B73K3ZWOXluvCF84iEsLRnEdH174rcPrWdfs3K29pPe2aaThz5f
6suzK7BitkyQNPM68qHNhl8or7EebBshwwrfh60JMS9szSsT3LiYhDtwVSZiEmLj
+LgY3yGN4T2j0wsoUns8Q280FivJjma/tg+nvwLRiLYBtK0xW6eAzC/8uZWQcbDC
GM3+HSfNDVxuOFYKtlBGCJdxhlL2rIR8ShHrGf5V0RmBcIN8K9XgnRB4MC2KJtM5
QIjLDbHAUj0JYaG7NlA50vey+JXigCxlsZj/DnciHZ27Csk0Aoz29SHxJJmaEBYY
a1m3CR3T3PF0j6qHduCNqfQGp3Zv3T67ey6TlcY/xjD/5HXOKOinQV9pviCwrZXK
h88W/SK2+V2Cvsf6phoA9r1tMSf0KV2jQJYhhZC1Gpfq7R+UIhYIUKnJHKhei5sj
nXfJ05mlk5EwbgMC9oOgz7JZWOl1HG21EyQvl0OqKX6v4qMkOdwTDJFeSSYYgGoR
dWJ4V3PUGnSZZ09UP7p9HIn51ukpRQtLYLmYw76PA+vHZmLKhj6ti8wbkFYn6DGV
pBLp5MtGnN5DZG3ADExfhC7VtRZi9RSYJHfzGSHxTwmbbRn4JVN1dSzBovi9LoS/
TYdj+NNjkXv+DC2EMQVFC7VUo2G8fSI6YvyZv+xPSavrOrG/+W7J3aI/PeGaBUop
XEttlq6Qu+NjkyVspIeQMvSfNMw1cks26TC0uHl/KOJAlPWj4stY+TCtxn421Ug+
/Hjy2lXNSb6NxO/+XBYyVFEw1dZ5wJSCwViao8239BOMuUy75sQbZRQ+mSb45lx8
W/trXRJuIjRKMUbHvE3Hb6U8BnAvsO/WuYweHQp1KRzlO9m9OskfGuIZNGoUmmJq
8b35D93KhpWivk05qsB5rXyFPk6Yvvbg2k2lFdCttsgqqlUS6s+BeLCtTLenngSz
zEh9lKmL4/j3o6Pu0OsVDgtTqlrtCJm7FTfgl8Iz5Xpu2CPjqVCa91rlhKp8QSxk
wI05qWqThI/cq0V6wTSGWRE+p+79T6dbMJjk0pdi0VWUnIn/kbtOcDIx4EsFLYkM
usC9ylrl9mHSV28g1zBb8MYqdCtYGorYYf4wsfLaXr7O6HIyI7yTLt5rQs/5Wd5K
iXhKIWRbo9hRAbkUrO/Or9BWz04dxl9YEzGZgVpvlSJb22pjW0OTixAP5jYL9mTb
MBAJ0uCNJ9C/JGg7ULe/erUdX8SfocCmLdHTP2USQDw2uoMdqEq5QURCmCx5zsf2
wbRYBwB2+3BQTHaO6DdZJwsBsEyK5I0uK9cSSuzI3VDg9NYAYngsX7SljdObOyhg
ztrqjZqnz2AP0Q5oovsMZzRQYMnqhA8BXzSRapAVNXMqyki14KuqyPCgBledQiMT
zvCYedvNZa0sbNbuRy6KEYYc2vFhRScMOtLgxObidaVMtENTu3oEycpwt/jLyx81
e/WA4hrxh5B75ggqFYnTg+q53Eq4pvzCGinbINhASmYmbk6AUNSrqWkUc6QD1FbI
ApQgftbUqAaMriu8MmU+j1fHhT2RHOiuk9eO6fsJUJnzYF8DCbPLjE8UhWVEN952
bL7u+NJARz85jodc2J7+hyzkICd31u0L6FkAFBQWHyrnrHY8RG3UwertVHwaNWuT
B+zbY38aYTzg8fWwScKw2Tff1bfgVw5y75apyxDP3R2uuKX8F2qlXJSZVzE4IyXm
YbahbvoUu/5o8m1EeFrumbKq1/ryUcI9NzFGArth3m2J4+CPJyP833FIOvQFgGwd
Zqs1K1xLDAVE2JUySoz0iDstU7HfhwJdpQwGFxVQOL3FS0LX5ldinmXx+eFdGK9U
u7BwR5Qfe05tg+I8+hQseLI2aiZzAZGbjfwD111+PZWc4bLkD1VVWMW+DQ+pR6f0
JeBq5FOyEFWNr5MdWSEmZ9q1L9IjcWwEPibe7PM1gO8xKi5TSz8lOoSDRmVO9c4F
9HMVtYyIQpbhaTakNeDApg+rIUi1rZtiHsxbxFW2KpqYExB5yqq86Yp3/vRUmdL6
+j32dNAu/AxbgoxDRAq5n2XPjBffiAbsoKUDHeICaKKiFhYMrGjvoo/ADuRVpa1D
6O+bbP4FYhK5MyNZozdFKFgJEjy95eXqsgVOpji1z8K64GdPSdvcYzILqk/luhZn
PPOdQ3EVCg3LeClpEH+q2BHpep/M8BxN+b8krcoyoVF0n9KXAMKs39v+VzTO9dc3
t2zMf0xsKw8YOD4KG/b6VJaNkg4ejxwTxW0u3HCj6d5Obv1ahSWLm+uq4xkwudgx
W7VgY65Z/MEwU9Kv/5Tt8NESGKXRsZ19alp7//u0lW4Y9G1j7l6Re2doJUdpf1qJ
mcJb3Vrbq9ZqOVLWkHzuqz0f6uN2oDnLOixx+kk4HiCje5YFqpcWLj5DPbVkGuIv
I5QS3EZetY6DVkqRkabpcxRLKUgi5wZI2cs9/+sHCAqgmSBSoepxzVvZoTMYwKFr
4N8XtyQg6SqrqueZmfhOlkWbP/MZjcOXGC50syNjCzkWqV4Qer3w3IepUOU4KvhT
6RbJkdeP5O/t0MxCjU1PwF9i5qlOClkr9yZI0jj5VcYawixZtMmgG/1AYNkb+kyq
Uh19/EylZNgKJsSm/qcda2m/D4eigiXhwNg2sacbcfk5GEPAVyfZAbmzbrIDHEHQ
u9UQb0G68+9JynIIO8uaK793elNo6Q+FhtlyDCk/LhUWvc5eZhWd3XYeZK/c+98c
Aov/K97lhpMDS7HRx/10jGFJ+4Snf9RPajUajdTunxJe0RMmpKUR9EL+62pny/LS
3oN9yoAHt5hXG2ePaDRrlh53RvhTnTvOkhovttqeREL7LjDV7pXUqlBuNrutUFiA
NH9AUFH5MorbW+bdfcZkC+7ss/dSvr9vh3impDnPQZM+bckOyytPj3LZNk3SPJlM
ht8fHCjGYDg6BimMh23wAFT1fSPRln6CBLLSyRFaIdOWJ0sQDk6WsNtOxQ1A7kLn
AmEgvUtloLi3OSR0WaW7rp+BN4NnYWM4HE1ToE3ULv3qLA874XAr3NJ52SUdMh2g
MxyuOOSNU6NvEejLjTafx7xbj2bueDlmDlJUWD0yWD1zJEglz6f8ywBomO0Mbwpl
xGMesdocfeXHtL+JwkXFSMP/3oDnZJaZWRZsT60wjcdeTehlnSaeo1le5/4CLKnQ
PtdEnB5GksVswk55mqTWB+B1h1YICf5tPd7iHk0IMPL56+y+MuxX4KMNvENaHHxq
wDMeYj2dUtDpYymvChqImEkRQUzHmWF2nMlXeT2iaRff6FDBtMCdgFg6eC55qirU
SyhOb2mUIz4W4VMJB+iV9skDwRNWGEutNUb3ow/woa/2WZ3VY1Us/6g3JfkdS/xB
9TAtFjgClgZgVvjj6MNFZFePl3I4pHGXZHSvebjRjCZ3vr2TWW0y3L+4yhdJuJ4f
N1gIuxzdQrX2dx7DbXdVGTpSyFFsMhSmc4AFXe7fESqg9eHGADlSSjNJgqipHWCR
TDxlKKs8ScsiPfPxnZM6iP/9+ZOw8zmrX+OigB7wW9Tp9BZUVe7/mNwm4RPM8CtO
6V4qrj/2bv06TtIbTQs2/ZZZrQiTcnamnRGiZr3f5PMvpfSSiWOGRLgEdrxrjUMF
VmYzBXuikGxlnJa+C1pRp1aFn0j1UCnelAjQVvT8Xmqdp9rtWRmq9FF2uP/nhlgS
cXA+CU9WxFJQqPgwf6gYCl8NmCsZIHEolepqKci/JKKhUhpL8RDFqBwXIms9jPjX
H3Hm6EGhkVJFLR2C3NpclqRQdclgUiPQHTc9x8NiNLZus9Ik3UJ9SyoZ/DXIPSYi
PSplw/8KAiP86nCA2rds+eMWLhIQsdhoWQl9s/r3r6jZdhvXmcGy+BKMNpbFNuXl
atcs/4HeiAZWbAQITFiKyRE2QE9o+yAYxlamALs28AIAcLPMxmJqNUKXCZAMzRl3
i0k17aZA3Iw0eQyEd8FB4y2HUWStoUFtC30EeoVLLpirKWALk51MnETEAyMZcshJ
yKTQjRiHEi9Po0MmyEPLhHbov8CBbIp28CNtl/aOE/ShH5zlbHyAfDGTB6qtQT5P
4BwUgITo+f2/EDRvisuG2AnFh7up/2JPp9Ys2j3CXpZ+ZkGY7YOZPO2NZ0vc1WPc
wjHuPTKP1Z10ctzRZ/aI37aCgeeZZ78WJL/rdNX+a7i47Wm4o1EJpNCOxl9pRSKA
da3m4EKJBGiVxiU4j582GZ3n3upr3jwDo1a0hlhmP1+xkY+C18SPFnD2U/7qpkbs
FKegbtbJ94B0Pt11LaP5t8qR8nIZ7tgL8ccVpCzy63uQnqVTXfKkMC8Y/l+/YruO
D/4uxlXw/eTfn6FhRycl8qNlwSwRRbjJulO0JhIIPJUQBpFoifJr+FvihrQO/7i5
tAWS8BzayGNnj21tnmQrb9tVfJCb160QU2NzK/vMRGG4YRFb9UlTln/iGZ8nUb0s
phN9T+AEJ/gHTxqxFRVoKzbdcAEfonMCGwSYawxhdfXOP33jOZGXXc8ifX5ALgzE
rCi7FPx7Tg8c2l3r/KQ0eplT4XtLa0ptuyvhdH9puvncVIHDu0OwNGn5OMgscWpR
zqD1AJpWDiQcZpXkujrHmhYaWXvPnGnoZ8Bf/BR0S0ocy1elLW4JJ57Qi772V5CZ
QEuDP6UVxVmT1RBRDxANB8Eb0wlRkuy6UHHoZksHXV/QL3U/X48nGKntCxo6WHVs
LYYmzQ8DRXBob99s2No2NEocFurGxptcF3p31D2zkNXqyObiuJhtuQZkCSyhjUWh
xsQSlpobMZ9UN5cJN2k6he+w5LDH+YX1lyKUilSbAs3Jyc/zR2+0KintLuVLKhpj
MI8WGmI9sokX2M2eusE3JQOvhXIdnj1KtmS+8VzV8mMj8QH/dVXt9lhSXyLqYEJb
2WoK0ms9FAOJPPtIJ7eyFyTUmbOIe4tYyo/17S1pqffYi6wow1XaU1jsyfW2Q11v
ALdK8Ql4K5UYmhfSShgMb5WJ7Kyz/Z7QuMPeDygl9LisG/tFFZR/kfB4xkv1SEfH
dZbc7KG2wAF2DG4lHHjHvX/FdEpXUQjrRsPAK+XAKfJykMxVCg2Lrn4CSLzoDOpl
o/zZpzm9lTtIj+NU6mYm3xZBcVxIEts0FjWEn9wfKm1w0hqZipdMnsnsI28f7IsI
8rHrHqtI+GMoJWmG9vGmfEi67Baf4OvhgZ9pqyjJ/8Gv3n3gqyu5CB3TNKij73dX
y2S3Y+DNpqeSPsko1zwDM2pR3vlNaLDx8vrpXfglRv7S1CzLxaDPO3gAS9wPO+LD
euttS3/U3agjtlGfLDFBUnF3/8PXmsNMSHTLhbMEZLvqGiWu0iGZjxfrqY9Ciu9g
0tX6gikyLVKw6XSJkbrvTwYyoM///dnByBQOP4slRaqdKslc49oW0WyCJED3NDnF
QALJQnSqi5b8JsXEV4jyHV4HhrZ/TMdCavsrrsxiB52SJ4trMPjH0Di8FEZsq3aJ
PyVhUWnx+6sTHCbvjeUmW/kH1PLLs9pD5AREdexGoxHA+P2+NVsNXXKPC7qR+n4I
D6xU2jN2S6brXeYDFMxFYU7Y5b5ChRnsrYhhaz5g6Ee54/8W47iqIEXMsk6NVbmg
+Stm5yVKtha5i1G/7KMy7NbA6jzQ2xJ93M4XZKr9JLAV1FdSw+kgEzzvmSrz58T8
gFDo6Cc04foNFXFQPWt3UcCKlY50gxQDNEJoPCKAzLK5WiOYzcHDF+Dj2ts7rtWv
QbJOAkuvK+odYkYP1M6F+RXiDX/6hRRG+8J0bkskdzXMdTOG/lfCYunHgNFhJPAy
ennM5YKG4ZWFx+hw6G3gKnXHysNmkH4MhYCBv3gPyvNa9bnJDCIQoZ/Ic8pUdgLa
8C92SEQF9lN+w+bQ1k3S77q5O4vkw6+XwGRlxOAY/vZTW7mwG13qoTdQb5gaUrFB
ULoCWR2XeExKUl5eSwHfTjoM8LXvq5ML6XD4v8uT6IzDFAcc0EDaEreyPe9J01K0
PP/3ee/uqP7cq64McTYQc3ytLojeZSMOEbr8KxTYQiEwCBGG+y4XLz4KensxMzF7
XaUO8r30LUiQiwQBHEua4p4eW7PUDaXil3nm8MVS9Px5GkxVsca42864GrnrGs3c
Chd9dcRCaJd+QVFGTTP19d0IbjASMPzXVcJIcxPMzzmwKZY3UOQpuNxAfkGrIK58
RY4M2mViiEK6ybtj7hKnWiJHvkA+eu1d8tu+4aNx0Akm15/tHC96LPSvYycP2YZe
nuGi7hyN9kbgJYcznnd5lqZ2Pbucx6Z4W3lcCEVZqgNs6Y8qjnGvfPfORXN7KXzf
hfd1T4W0LVlLUSa+rjigKFh020SaXkpoV8ob7elBT2ULxpchNWSOgvhV5BZHw147
Q+0ctpUwWXAx2iIfVj3zK4nBlSnR+gXBNn4Tlhua+xgH8JpKXZjrfkPgOKatpUDD
2t0eVsPpMVBUiT8/TZSS06uQWj2N0uA48kIaU/xPtpDv3mKYFnfMAL+Ge8ovMoUx
CXek1jIodWXrh5241KRrGiMUXQmjkCadzuHvYc9MtsssfVqegqDhBfSuLFpIbluy
XB1PN7PREx3D5dJe4jClCIs5T6KdpGMeqKUn1Q0L357RlE6F8u0YX7cHvEGPFbke
3uGJL9AJw8klZaN0POT6y+ukfEzRSh6wsF0psu41i8rvn+IclthtnmWiGyZOpmYa
kFbM+7MkhjGpbuq8uR/RVSoAcQnBj+BKN8gAcDIesvQXbXXZnYsVGhVBXHKCV595
QtbPEn60kawj52weChiTRc6ANZKiMI7WWCqEgc09MorF9RuT8q4YRfglam6UEdMx
j+KT2Y7viXekunA4VP4Y/LSIPc0iY5gCx7+mzgZi7oXFxKw+MdMfGEHJqMOd7A2i
tbkWSLZao3Mx+B0DuyVXrUbHkH1McIqvTKHYX8GJtiMxa0odKH393yrPnFn2xXHA
rS31Td1vnKjLIRZuKaisKFV94Trm+aIYcR6A9d1GNGGJuvwSe2yvtpdZY8SyIz82
Shk2mIaPpSQEV5Rfe62TiasmYglANAIBLrUP3v6QXJMqCKY8i7PdpUbaaSBMFX+M
NNDBAPmrYESiuVGiaIPNll+8z3MAG2/JK+UcW22aARtQS6YC/27PouM8bTZGQRiI
7HkHCoR1GJ4c9+5Ifpe8Rg1N6sXmHQVaFwW4go3fqvtFXrIu3tKvZI1jF/16iCFK
LEKTz+f53D0A15iSSD9nX4WdmQEaHPLXmBBUapGX7kzZ1eNBnKm37t3P+Ril3JyE
Bvu1K8Gjt4t4SwB4kif/04aqMFY/MMJ6tULcL8TEmXYOXNG+lIuBn0a+YnM0KQjY
Y16tmIdQ/o+qne5PQh59UxO3ScnW4PcHt9SAv6eblsIap1+ZGVazZ9l/N6q21gyc
aNYAG8I94V8vBwzx5x37v9lLa7pdj4toeHxxLOgWH+51WHakwJy7lPh9Pc8jDzZY
ZAc36H6ICHMR0QNJ+7Haej7sCOsVbmATIy4LACul9PXlrEAqsnUALk3gxvzSPRmy
msVL6bBHgZ/09Jxfl2I+ka7eCrj0sBW7d8nMVBrMNgDadCK5UntzWrNdzql2b1Gx
FipH72BssKUa4hNPwWEzbZeey+VuPtywtVnXL9tprcRg1/iVRAR0Tdw1YZ5P3THy
ZA1uwA24i27ZInT8/quLvjc0QohV2RWQ5NFCr4/+BDrB27Qpvz/3ZkgrEvVNFNy9
dWK7IHjctq2FpJBvZXriT1X8XmK8cpPeGv/IJw0mfLHT6GtUg6Qtpg+v0+8jLwCK
uxM09Vg06yX/KJjm1oI4zceWMsSmM/33XynNm/+dV2/a3vSOMDgLtBkTW89/n2MX
Ieb29pLE0gYmPGidj1QrfoZIh55UvtPbS8o2KQ/OdNyOFKXi18IJG5w7rBpdfL6c
LFZYnvOOzIkpfqS3Td93ON+U84iGT32Y6hq8tR1pl5TUidt16311iNxpXuQIBnQu
YwAAt68oAjstYIdFoiEXzcptTPAJ6Z+5WSPonhB7CGhksn/fkaIy+Cy+b2L22j2v
ca3fKbbgEt92iYsWrDAtoiOyoDpOOuEMjVBFq51nmFEYsQtc1g+jzca+1r2TOf8f
DJyLcKSbTVPunSVDQeeCdrPY2soWEGbKohtPu2UI+DivsubYkSQKtCKw6l3Y0442
wD8EdfkSNvWRjSZaEsXheY52CdqlhJdjiKlwEWoMQBbxvruwxchUtPyQ5L6OTQIz
8y8Zg7W94iHWKZ1BCwnaURT1O6/5SZy0ng08Kd5zT8nIWQhWANIIZLjQ4inmwKdq
C9k59I7wUTzlXjzkQ/rWSl1HOCkS0sU1xtTupefb6vkC+MOEE6/PFRvdiWz1rQi+
QWjgAycryOQp90MS6YlN5+5CXpcHZ8ISYjKm2nkrOdFsAOKOJ0d5u8KKKoJHzHPp
up5ASENikFzS1eOttDrakwjeDCYU+ACvtDq/mcup2YGDFIjfa5TPPRkJLu7W3iap
Djhj9zkMaFCgJYUehTgMNH8DNjcUbUE5OYVx0Hh1vSNRKQhDZJGn2Pj+tnYyNYVf
vCCz7Z3RCq5kikLoZUIbt2/r4t2Lftn0jiet4JWgf9HOPcpj2xxWHjoH0ng2Oid1
wfSDi9ymvI0UXht63kV1zd5XCtqT00PQFuDyGik1kPsIjnpNSiW9woTwRRsfvqCi
fV+CPdmBzvyJwHm+ZPTgYjkWPqH3hKLZyng0lm5jUBFH1I338IEStghY86bXIjzU
uhDbMGsa8dobTY9s1HsvpEarSNGYo7sU1j3McWek+Gxcku5X07U3Bebnujk0tmiV
2rSkVl80fZjVNev0EYKdjmgJGTlrT7qCvBVr5/jteHaoCzGRN23Xcql1sNKU+WdD
xG2B2U8TaLEkDv1rAI5UrSwOK+La6Jvx6KirTLsw6nO1W0hIBhDWRtdxTB7PUj0U
dZ+ZvfeLbiQe0xUK0wOZbHulOdxEpcXBSgy+hHdaplLfrsMAqPn3rCul/3DX2c8g
q/LnVlJNHDsHm4tYKMA4atEFLuYwMhr7uwQxU192qlFIRt43r5105zRv9eia0I/P
mgJBlxT58jmFwaD1sDzMtpV3hZqeOyKL70fmtfbS5Dc3HPrbFW8VQ0jIDZ1cdBg2
CzfETcb//4CiSWt0amRMbcBrtsr20cMs6uQg2Eihx9AxrVg7Aofem2ipna7qj05m
cDlRfITNJTHuLMFJQ9uzmK6GCpbkKBdaRsjwlBcYtDctJtA+2QY8UTLrffzCQ1p6
GpkjUbw75ptJ3sN6PW7+NVzqyX/p6TxLP8FP1hbIzfGFH5VjimkujcpcOd5ZsrJb
MXVg+kkr43W5UPUAG9IKv9y0R0b/4iS5A1QW/hAh1Xl9EH8yQkFlDEMCYnpVCLIs
VopM7WanvxbFBD59fa8rAdMaiuIWLurCGWYapXYpoZOFfnpWDFoFIWlwNBLliW1O
iO/UWoJpxhl0nWe141K1Y1FY3K8Tc35bVsezKos+yPBfKDA3ox9GmXWeNAd4/jHo
0hmK6YOs3WOTz2+O8V10Jmz0TVM1yePcL7SUBGH6PUAmv9mXqHOYKdi5ji2qN0mW
GbzuiHkRg1RQfOFilCxWfhhXyNzuPIWDzkxveqMxM0m971p0+Il+iW7SmzyW2t6i
91sHm2C1Ikc03oECpCSVgJod1U58HH2ODD50kTph+2JlzbuJbd3IVzevfjGPI56V
kC6INsrkoeQIJejMMOSrojn7lcbi5UXIqOy/wTdplm1IMMRsJbxlUwbkJvy1t2Al
GqC0ll8nc3a7kKhQ0rPobimfFRhJZBvUTe8ESxzTBcS7M6pwQ6wLWq0lEBDVdilL
PkUAhx7Y7gzBuI4x/zxQwXBkL/+LWgr2DVClyA2POpxaBHFi3jYo6hh0Tw/6QaGd
tqPT9BflBpPDJZjRq/pQAS4wAmJSD6bg3Vj9BC7yPk/3ERRTDWAyaE5FhrG02IXf
ezw744AIcKbGWhOEyfK4WLPcqqAOCo1Lvf/wzBpKugtXXVkUrJYOT0+sF3rRq4Lq
Ih7LrU3ieoqVOauqwOjHz4bnBMEUL0I0cmROlSM4QHYKha2r1Oc10I+9NVDYQ4Xj
mPBrFG3iCm60XgOdJCtgH+oSW+vaVJPiiky32M49Wz6PfjhwtjiCZ+ulqsUCMgph
P4QNyqxacgOLaujVyu7ER4rpfWF77d8WkDSEku+okgmyRYLsRtt4rG+ARPTy2bTW
ukCZjsDlKdBGWr+e0MH4Rf5c+2XMuoVxsrokZDfMnLE81Wi+9kR9hIiqsMgVspET
eHosDux/dS5cBqbrb1p06NcKNtMMFJNSlx9qUcNpQUwPF131MBXjvz1Ys4Dw8WOX
RW0meOZ/AE736SBQy6XBSO8XlUUXqpGShkDqD8HymYSsi0Ewuul7UIGeyn1p06OI
8qMQtlzUX8roo3PRL8rtDU1fh085OGuTk3IzGUZD+AUnb8N4qjy0VXKS23wy/xlA
+5LVTXBEgnZFz6vdk4QauQGksKWcucODbnMYk+43IFFDM9Wp1oyyyUQ7xSOe5iJm
F1Kpr6hvWEUVbh5SajD3vaYoBS4w25UKc7Lg9jxZHlRHer3apJwB+3HSb5dJp1Ek
elfN/zHdgV/wMpXg7zvAVR4HXE+lnBsBUO2U913cZN6bnQ5qGYKvp/kTqLBw6AW2
jWUcQDxKi0B9nJcYFWwhOKetHNnfmBHqfDepH+Bx52edIVeUUJMLmcKIzrP44T7d
TNReUORscS1cpBHi63uM3+RXuvI57+YQa4cQ6Kdn/g6iGQOoIbR0P+yGFacVbIsA
UdD4k0XG09S5MQ7h49pAYyCcj9cix4Ijss0h3CNRVFF04lagWeBiWp7QOU8dyypT
uYRIeAUt2FFJcCmboCJ0H82CQ9AVbtjocfmXT3E1K10mHsYOI6w2OaVEIUshE4GD
ldXzY+6+5ghekTfj5AoIn0NvU2l0DySOoRn1F7WfQHuB7aPgr5V7RYOvBcpDhq5U
PZvkr3hKocm5hYEH4X2xJLLTqL03O2PBEhSGtqTBGnhrUR9+Sv9HZRYBKerNFEhI
Hu+/0K26hDbrlbxl32pbD4KpHPXkPJsCf38z4z++z6MG5nNuiqDlNR2h250PqvMo
vf6nDadmpNRtdnP4nG1BTrSH79iyA4w+xtH/ivC8lk0iTQSwiz0+nJQFXPaG9Ppq
h+H1E1n/1NrBung8pqYpM7o277DkVMlJXuHcWk+S/5yt9kGa3zaO8Uu/ksbo2DqE
PzVtBlpxvy+MouDIY36dH7eKIbzdjlchyKEIUsLVFBsjRH5AH5z/DoQ1tSyB7JnS
NQMKu6vd8QTzOa7fObR5i9ZkGuku5uei56418kHgW3ZCQpMPbInxiCCvslxCaoJm
rVj4MoXn1WPqnbGgIlD7Pomr7qnGQ4vntRQumGIZy9vnPHb69uejdDK8qY6wRNbH
1uVnaC6J5T7eM3PWBECyrCLO6z6eVu0DqgsABtLVtpVgIwPY8wuKuoYr8EvonFo0
KjvGWQb4Y/B/exxw///TeMX2306z9VHtRg/joZ9j0e5GP3UzL7PLJcWse4JmA2I+
/VovdVa33H2dmMTNAreCF9za8Y9rc7AvRZbr6pvAb/AQYEUgQbW0YSt4whZfZrbs
c1RLj+gnKl4GQsMERf5hp15zxzwl9LqsWpCnUByRsIp7V66xRFWrVlM6+7qj1yfF
gE/gcFFV6NDbdp9aBOx+mIgJ8uvW9HdFw3ibQBWqQG1S8otuc/Pl4lbeeoxlZDD4
TBnHTTSQ01BJB3robTk4XIRdcGXCzRBF+fVdIADtDTNjqkNonInZAxMNVzPVJ9L7
PtD2Ko/1zJ/qcSn8fE+e+YmaLYbaBC9tXVZFCVpmOmn7iL8vjalYEZmXHRMZxA8y
y3/Mto6FL6MMP7d/fv/7FpAsEDIL/8EUy++xaD8xhdY2gvJJuoOSeildnOhlNTgm
74exjS1/998uvdmE3LXi6O+aebgua3blKcEv8sICRBjHxPB0FCgIrUX1oNoXLrfz
ZURlKARpE7iY8XvkZT1d6ZETS3uDBwW/BTCxYIP6qIb8lO6mrudFQXG7mU02iUUr
M0CC86r0kZQEM0TOLM4V7/W+JpvghZnom7eEUVTyi5vVEGCnMhfqtdMJhxAmpD7Z
5cjbog9Zf0r2mHIIdjzlFNFRHzM6Rxg8e5J2l1L+KxTSZuOuTLKtBcWIKL5mUviX
8ihDhm2bmHVxXogtfLQMT/Rxaeb2y0HH96rY6X4LEjLIjAaVuiaSSq4aJgQCHTd/
ydHQ34C+nq/5WBGzxE29UshTmtzPGheH2sLkhs3KiFnIjJtoE6dpgqGf8R2PH4mR
jhmESzFFlyaJd4+CEFxsL2xTmX4oNFx6+vg+fzC/EaWiSMQnD9zj9Q8w4iXXsxut
1klLyoVhDUp8ltWbVBA1oTwjppVbhQyAope7rEcQmGF48W+mmtTkpY0yKz5PdCe8
NOd918GDYDkQsPmfDAoAcu8O+fv9+BYjJ7wiK2aCZWgqnPAZH54BDt3v/yvDFSOX
L5mg2kPert2FyqwqKznlFFUAx7ZqfSJjL39mTlW/GDDGJoi65rNpct1UAexDr/ja
Yai8QtmoPwFge99HhGgIEKwPAnjlr+bpt9/UV8jUHqKdv2a06QqYSreu264IQOut
dTg9kNFqX/du9aCFybaDJMqFkFqsDvra6qjlWfIpxuN1qykKbp+0oI/5er8PgyEK
GeAOllBXNFkz5YMM83zZftLl+Jfg2wzVE1B2b2FzdzmmpOJt6V8RiRASD129YTOd
vhEC2+A6OMLxE2jNrsJJb7DJ90GTEEE7wCjUuKf5x5ovj/xWQNnZu71bWSF6vgFT
SfPrBHRoE/oLcUsjD1gSoeI+I+wfEUNGmhL9fkXc4jtWi4pwWHyX8iQ1KaV1YQMd
jBKvmPrnxi6Q8so+MaYNwFEZK2N6+3yUqqHf2O8ODU1KMo9jzF4Acvaimc0l2wpR
abpgflP1GnTv3OJA3g8SAJftYDTA8rJzRAyIdaRew2B+KrjkCIsHg9SZEyCRYMiy
6v5fXvgnxGHUFtQFOEMIPscadC9YMgTWYZXjSlxV5YCcJWsx3/pSDttTw9MsZ9ee
BPHwiS22MsBEYIEWopU0LSmc1oPl550GFRDXwa/gl1U3s1y5io5U8OObMShkkJIS
kJjVSTMEr7B+kaxp0lWE4XgZoE2BvYXpK9ebjY0cffY+jWISo5dEYBAFnb3t/0Q8
AyBXe2+jqJN2dorQTUKFbxJVPRuhmyuqQ2Q64Qyvx0GB3NXyYTkxeR30djmyY6/f
Gnkq/z0sZ9kr/HYQVd0q07grttCIDwuvQm18JVVlpMU9YXTQet/aLg2PSbNN/GZZ
AAtiRspeBlEIMsfop+IqzOOANkDrKMPOjRR5KoGFIs8o+gf2cUiU1R5tqzJJf7aX
4pjmtoDQAe/YcjTAXZCX9tau6dts2wSm2vKMeumqJVSRxY01wrJkhbLg2NYAosp5
JAD6zwxKoxdzfsK5xuvinBVwbPUTopacPBX8dAKmv/kqLnO76Ofzx0idjwvnt/vY
9HU0makuiRF8e3KRKdtry8DH5fuf2yEJiajjypZQBny/oDnk/1RICrLl+MwAvrHK
aAwoNOf2o8mZeuzji/BIDlZ3LTmIM17K2v6E2vlS0B/5nxOIpna4L7TX321hmFwK
TyDt+rSBYHgvBi18E0YMV1BjBSa8bU82Gt7U8sZ2bg9kVJCcHtIuc/Ki1+I5Kk4k
MBnM5XcDfOfYtPcW3wNBEErXj4GAParxJsLeZz85FPL8CL8XAe1GYQfvFadujkJu
K1soru44mLDJGhgHgNyES0JmoexO6/5vJzKBl/zXyDBOa2wjMSWlnVZtmWoZe1e8
LNRd0kM0mSrJ0JLUUwl+vCg6ec4ihVt48JbDc1x1MAFuz6OFaEyvMCn3kJPc7vUX
ir7onQ2qBX3wHFs80vRa5a+nkZEqDXq6KVLVmLfBqRShOJCz7WZhjFJmt1OvvqPk
v09zIny/upr8MJolbZgR/tR3jbQDcwSG66swEplH1wicXc08iABjAk2jurERyqng
NTYfg+gybL0pBThiZDjNrhIu55TSg9djzI5tgTqNqapJpAg5AkWp/aaVx6Fkoz/f
yt1SxtwBFCrPnwddpDAml6mEH116hhNhCayfIfO65FqcWbDhgS4pl2T8ngCm4qMC
8BWPxhkvV2RlKB3IUcRSIn2NGT7Mk1ffkpJfzQ/HHvYM2UJrnqUfh1k+USYR3WET
XTfPq8MPvONMKNT661Olbx6geKHcDAw9CDioPHpY8o8nUJHnU3ME+Db33UgCaZ6t
kuPunZ75/dXGPHZmw+Ab6Yr8tHli4aaUf3mPV3kZ7w+4WaTVvZuoyjr6fbj+twmL
HAD6xzkMNPL6Yq5ZLSbsNEJG3wslMbiBsgoHIeIgSuk6fR13yqzn6jdxFda+brj7
okMnNykLrEF15fHpqRH5CfNuxj0fD2nsj6QCWKT4vahhxin119iPXsnzk5jMAg4E
xCpJslHZE0cVaa9IHVCxy0SPHD5jf5S/gM9g8Vr1Qtpb4pKZQppsAfFwb/BJk/T2
Tc3MjoUXFVYY2+b60AQ2S+0SioVEa2bZHevcPU7VIYyZqINmKsPLz2kytGrQVH9Z
Y1k9AvL/XnmbAh3d1f1Hnn+xNR43I00OaZZUWCUDAVVpy+aPfwSHn43JCk4welWp
OKKoGjC6NiRWEMsAOY5OeHdA75JsN0RCSYm0ArLHjreHABu+u4Y7Bhi/yLznNv4Q
6S+7HdlL9sehNyQqX7Z13ZsOdX3gUolANLNXyZ+Hnu1EW6iEIFSem7V+eESapxcw
eOJA9DKacfT/ChCc4Nd+tr/hy9YGbRzzFu6NBXEGktuGnKZlyXgXQ0xxcwbADk2L
F7DUgyRjQne14ciTEzeIKR9lmFBkQF0N2U2nLmdgadzbe607bVv1AR9fmFjrfePC
QWrl7eF9/6XK+7VuJAbKdkYAR/YTo3s+VWQNHO0x5Pf3dwH+1AC+f+etCDj96hSx
Va/s50MqyZcr41+h7TeaSlfHIP1MOJlMcAhFzMoQSb9XZUG/W2Bpw8gwbDrOqB1L
JdGf+NtRjpu5lhuxVs8xGu0wXXs726ib7fdHb6KD6imgz9Hupl1sx8eC1DR3JOLV
haHTWft98c8gVAS5bLBB641IwqcDGxtktXe04JAExJxyxabymeT2aFokCVKAX/vv
UZIZMukQeE5avFyeu9R63nEzqnFKv4MZDqgewQpf6C7BLaInRU85bxvLS6S/jPDM
KPD0DGf71oJUUiIOJzRjCKuVkrrUG2YZU3L88tPEUZaSH5E1K8sJuNftsO3+jumV
il/RlK/Z7DcoclXz+yVdpQgcY9az854M6o925iowtdRsfRXVymkTY5HiKFh3yVuC
6qbnn7ZsQHhLUGoYJNinfiNiZONw//pWz+6yf4BCN2fcUPgXFmZANWc9BKetahUE
LtbIyzc9Ugp853orSb7yEDsrOVe1laDRz2/pHldaWPJyJvuLD11QpIo5L/OdFVCS
OfIYAXctwTr6C03tIikjPC891InxCm8xvEdvkO2k1MvfF9UbNllFrlhxQec1ZmYq
+NFQBrK8LZCPc5y7AHIwOZjDMKI040RD6pazt9f5WZbxHDUy8r6xjsVMliP8HbL0
m33tZcbJ1u+mnWsz7uwXQtyfTqV8+JmpTCQhYHccQfUiM9XOwSm7MRbxgO4y3Nd3
iyORFSGmjk/p49NItRpZqR0UDSgh3RPQBySybYFQxiwEWHtHDWJwHUYpkkbgI9v+
CpJ8Y8UqDVxq2+xmcggy846ADiRjPVj56YuIvxtqdOgsK1sf2lYXh7QJByWOt+wi
9Sc6Tnz4lb7pvHYwboMvSq5jh8hVOwQxqqLmul7btdZsUmVaNdcY+uavpQg7pm9E
ZNNaGk8SLoydcHLZvqZ/M6pHLq6aHS9zdyca5awn76mNcmkfM5m2qPBrdkHFZnJV
3q23zqQOjAYI+xXhgcbhYdDQtbUrd0Qnsn7eoJA9Z4s84F+HlxiNxt+ZBKrZZc8M
2nYr1UElnQyVQqGu0yi/psrbXZzVjo2wA26ClSVHTtOuH5jyLeaOIm3j7MBw7SQB
OG46kQxfTsuAHdbduck0GERf/2/Io9vjC8j6OlaYI0gNDwrpgQeTcHtuKwB5R3HN
JGm8XIpp7Ylp2RfUabAF9KZ5qagaQHN+thKI+G+PmMI1yqiq682Z5nkBA1VCXY++
xfoUodz3rt9cL0Vt5Ybzk0dWz5wfteZSoB2HzA8XgDF+Hw5/mbUNmJV8o9aHE3pd
Jz8O4h6XN3uq0toEiNKDEuKojcW7AUYbatX5dg6iJwMQkd/szK5Cwd4yvTpX782J
30xIMkRP5AEQmFhwG7OrG16TBdS5axF7tTPLqCSOaobFMQy9AACb7YBEWGxccYvV
lQ/pBR3wkqqQWVkG0YmQo6gNAyfqJbtl9NZqUOAREsNYyHTkT4D4B3a90dmdYPYP
iU0+TZmIuoKYust39lBs3N+pW9d0FKtuSxchcBVOae4S0aqzOD2QgMkh/USl1sNY
lB1JsPh0NlZ0h+vU0z5C2GmuqiQLfIIuora+9Lq7Mxf1JwD8H/y48c/w+97tIYDi
tKCUzBWCV4qejfa3quplSUJVm1pqHzBZvZI6sT2gKb2ba5DGUZHOKT6JRGKEVxWl
ISiXHMEq4zU6AdsLthjkhGfewHvtPbNu7fYuIEDkeZCg+hwyCBcUFLa81cX+zFtz
5spb99srbZA3SZqAX0UhbFq/Vqa6q0khk1K/JUBZCuLLhUCmEEzbenum1pXJqBDj
nbE4VjO43T1ASYyUyqNUX7Mw3qSudj11j0R87+OR+s/n7TGDN48ryA/TNe2mwUGX
l/6PPUMuCGlOk9LGFz91AoNJjhRaPtzLq9oo9mG86sN3NELOtLrJhppXIir67baC
xeL1jL+ZLGuLRwIS7Ms7ssOeGXfO0qYK6LP2GwqboRjMYID2x5VqsCqmB8hzAFoT
mcFGMeRj9Z1XrKXPip5dwY/ayY3aFZsaYoOJP4xOmiy0q/WrJG0YRzkH/KQcFkbO
MAGU00Et2GB3FVlo0oMcvSKziDfpmZoSXofgCqC3v73J9WiY2ClNzjzOlekAURPG
D7pfI0oq3tL8Vr9luJvvDPCgl2BPuZ9HdGwMvF2EVRNCjjlYGODjF8xh9lRag17c
2z4cd4e4uWvTZhJ52BLQG8MNLzLYTg7rEfcppbagRlHHaDE+Q+XSTvrdpJ8lYRig
V0es/lA+DgZdAasWbN2pM0LwoDNEXlrRR+Vd0aHmXmcbn1LYvhDzOaDOgMrQ61Rv
ahPvAl5tSr0v+JbiwOVNujIt+EK6bq6vhUWHcrFajySb4Lcd2zqFZ7MG4AbJba8v
HD6QI+D0KaUWcJMnXn6lClIThLrR3PwuFmxXg9xEYG9cIdyvyU+mFZGdd8FqfvHC
2+VgRUiGkoWFU3LPv3J0qbvVNmuPNt76+WF58v6xk8v6oMzWQddyhWLWb6MoflD3
KaY0gD9iVcUtO9R2qa6Z5AaK8zT5gzS0x4mRC1SQe3M/gA8ZrNItu2WejxWeP/UK
/BapzbEP9yWRhuAsMWC54wQLRJbT6IwP09xeOTOToLjVJXaBkKNcPiPXnkzNdzVt
LOr6Uk875kOXfk8IpGXQtgpfgwAhC9tV1PZMG0Ao89suc6BLuX4ph5nCf/wz6wVP
yGlIUjsh3vytVtHmEb4Q8K1PKMBQaVykLdzVxrxlj32qeEqU34PcG9Ipw9HmCA/b
M+PYg81VTAKxZ1qbhLtUvn265cCf8KYXQYkWY9ze2g5JINVWu8jvkMvVlQ8h/WBp
fN0PjYnubPGSEpWwrk2x8ic26P8cK1c8mRQvAtr42sEAln+v1wjJZG60TSoyyziW
RyfczlH8EKCS0qeOJelyRnIqo3vRYA9DE3iTdhHn0T83vRm6oUqvtzjmn/9e9oH3
3ckev3fKn1JpnXuo93yCZSktflC1XQo7sbdl2HaBUR6kCTewtTOTE88dZvw6wvBa
/bqSkISehw4UCwZAahc0uNFM14Tgenw/iptrRBIIVJmfC/umqdcl1BTHqa5bOYjX
6c96rjsn8o5L0x/aUV6TmFOFtkNGZPABR3tvv3ljyVihcA7PY6AGy4siTix/gjTj
djSv4/4Mxep15mqzt7xTY1cnG3MrlHLwTJABaqkO2PX8O40e+Jwe6hOapN7xBEln
zplGUXrWDluIXOxMjxB/+pvyUOnE/J3lTR+kvvHzWc0+u42lWLFaF1l7/D81+I/X
5unqHOOf9wv6vDadQu+KF2VUbpeyRZ19RnE71oyMOX/vJPTWIAQHpAc/5n2NBlqT
nPdH1iwUDMBay1LTKHv9HETMIioF3O5+hvdPPYC4MufcpdkNfsyOArqncSAbQv3Z
+bloObcXFgcWiPgBZ/eI0Sh9bbTIz4Ange+gs7gVQOspKVNbtmtzsiE47xHRkkB2
oUbe6eWBbWjmyBQZ8K/NNwpuFlW/Yp8AUfo8u+KHGSRTej0AvGdSVIBwMMOaSWor
gcFo2tCoxAtW1BGH1v3BhT4ogjv/I+dxoLBzMaEqP+Ld7SgBLD6NxFqohx7RuI4q
0hWkO9KHY80I9BDtYfr1ov4PZc64F3zbfvPrvIMDMfry3Y+OG6XNQG8Ng/gUVdP1
KaTxgB2GWknj6Vx/X6NsmoXI3xXc7UmyhSrHV3e/Alp2JoRpwcs9dMleWTKaMg5N
mEjyZ509lEB9EnBV/Kh5OeRLxqNup2J9OHf3UA7QcKxtc+SzYm1lzsHI9U19xxj3
O4xGox2nNmivZ1sttrth79kbQrZv8+33l584N6faRS1j7hjMCq9OfeGmHAab/MqG
hxW6TDKjmunOgxirZ7hwvDyhyd8PBApnnPVYeDo953AGzV5Lg5zV9TwbIFETaF2k
wzu5bs2SKb98s6uiz/at0SvcPS0LS/qxqwnUelOWlCkbPlAv42GgH9SH5tQswL3W
ODTOYm/QTsJM2XvBSJ1jLrjEYjaB8BaBHyWFaTTQovQj/TgCzfxqj0+z28XYGZvi
lu4zgctOxvEeKIc0+Is4E1Rww299NeBOASbkhUxA/H6UZxKx7/12XJamVFKEwWFM
l2M63EGzLWqO7o7nov6tnm1fG3a8vFZU5OIqCO3qkH7swDb2s4rhK75Y+viSKdJq
L5YWPQGKPNASTJinOiYLiQa+8jY+Z4saHTzZ0yLYqn7Sa+y/KBJjvyl1Q6f8/RyC
hUrFdDQ5PEL6IXzFAT4BOTSLO9doftCxyoHatTbXQFXyE6T6As9AFlFAk7R2Sqer
o6hspYBd/roduHpYXPKU8Fz09D4Lcx7MtWRdWQZ4F33oJ0pSOWxupyzbLUoRI/fp
snMQpE2K37PgOdeYJqso1GXcYp2rKfS2wgYzu7upksuLxC3ry/rvVfVlHwpVfyMZ
M7zZJ1bYo01vnd7SEAdp146BET+z9BUTnZI1r65ZHgIQyTG/Dehjbbu04hvCI5R5
UZd8K7tXWCd3JryoLTvET0/GMxAjDeNOL1AyvnkRb2AKSVs+SjGhEhztuiEaB3F2
hvA+m8Ts8UY84ByDUxWGdq58wu6ietxZ0NpfOt/7CL7vu6XOicQ+K3OtgYEPUT97
RW6jmJ/VhX0C774WKdeD7cfzNYrpDiG/gJScxTjqj1KcIE2i6CEEIStcFl/NS2Vn
BUquRJfgeP9m27zIJc4UZ7xqSsQt7dDftejw5ohRvAFtnv5F/jw3pgBF4GBOQ7xM
wx5gUmQWYG5X0ujlTnc4sIRTZWISVKOqBzPnJB75r5ltUpIrpoFYdPMoQ4mwUtvh
hSBoT1sItNpzOLWSrs6ndHoGOxedEqxHA/qx/hVto2QBS3UzVKSjrlQvlMfVgffv
8TWSY0bYOpwp4S0tnIbmaWjcOye4iuc4aSAYO42slHUsPQs2W4zOpkNEZky+IaCM
ZZUfS+ukXrcSFrkKvshVduh5eJfHhQLxbWc1AGiTA7bwyRrA72snwotFHgEdeAXP
06v/bU2UrHNjva4L73jwaduMLVFADG0loGnsR8PSTRWIUYwG4+kFDmg2RHVyhHmV
nNtlHVWmn89nrk50M35HMOTVMp6gm4e/zmggtlPiiWh9l/0gXF12z4G/XcreGXt6
nZe1hI2V2MsmTg66AJGdoJ9LBd+wpszcR0dBzZlV0mb33GtdwH9Fvs8izynnMIjP
gNAe4O9rGGbwzJUrrUGW2oyJGlPhN3SLbk5ipkj31pK2LM33C9u8HtSxjyO4gprU
T0GPqEYvf0kCw/TturnbixeWIyJjwxWc0DkA571o6AuOfM86Qr6vxxGelYq7A2ik
0nJMTkOMni2Ix+aEOoMbrLgiM4ai+vv/98e16t6QG6821gXVm517SiF27mdv7U+2
Na72OWWuFX1wGU1vnmmjJ7y3sCDoCs/IKWaod0kdYKg8Yll8cidx+lVLSILWa0BB
V3cyQBW0pE1+L/Sx3U5fKJa5ZriMKoxGgC6jLgfjDi+ZmBYtmL/ewyhPr94B+f/C
N+UgQWi8crs2BRGvDWZvA+DjasuqxFELk00JwhcKAXK/e8IbqBXZIrVyHNOK+RTP
8v52B6sJCig3Okx88jNw06CBgBdqieWkuyHq7rK77P4ROte1UAiPrcewCy5ytR6s
na2X75kR7I1LtUZM2Nakwokc8zjEV9rjdi95qeODZJ3wqzJvifBaNXFS3RGblVBe
AUcIdNnRDG4pASTxn0F5o/AwdiFB8DX608a3fcB5iImXBEbwVRIhQRkU5kp5P9NY
vmFS1sFiNb8/9orCAIQxN4gtzLwnhruVH3s7swDne112kyQBLXp7cQO7ll57EUq3
lIGO9+148o9FTDer/JGOh5lcev6lS+37CKyd+mua8r0f+64t4MhL26coSs37KdIX
85r8pd0uyZpXW0MNlvz46Be+ruJDjWJm8nnq4dWLXkwLDSF12nrJ7W8JMZtNp/ZF
eTybxF7af8L4BpksYN2YpAPO0lmNYoYKMOeOY6kpKheDJ/MgSQG2KSbufjgz83MA
3DWjFqN3VYcbMW3Yk7TiIhMeC0HvV98O/gzgDwcbKcapXlMHqs8I335CwSgWOGRb
FeG8YfRv68Bh4UTpeVgsvRzp9eC3IePg+xeQU2ZPltRlzjrmLompDBTuqz9qabK/
DQgkyLS5rQFzk3myba0sPqhLBo/ZqYNAbofWIZRni03LLDn6pzfjmUx9QTImfvnt
qI2xsZpMgWf58RFzLZuo7Zx5zsbPjjpuqMbmlQDRy5+fyhW1VNqSbSGZjnHj5uLu
xgeJ/tYfNVQQzJiAZeejymf0DDjzsduKuPfax1SvTNyyBY2j6ur9xR6wdUJM8gm6
xXdLWhu3dl7Z8QnikM98VnnUp14wVOx2SmlnQ2KB+TOaXWU0wZmfgYWqpCWiCjpf
m+CJsgWjASs6/UB9blFyFNI0zNkJfT2oT5v/Z/+HmSXwY4AWveZj2ZNVSPtKdWM+
60jMocB5/TFJ6cJDRjNwuKEMsnQCXUBYY3HAQba3My+kFH8Wd2mXejcxosFcuEUV
iuAB9ByNAaZhG45NsDKgSJ02qMuXoqjJ3XJVmOe7kmZ0TOvmugh5s+1yfzCt8LsG
Dv/s3bn5Ba3ukeSeVxLaT9u0rtK+8VY3U/DADVPSrsgUcuD3T/5DWxL+QgrdCRRx
DLJPsG016JXom+uy5VwsuAQUZbcTYnSMHQPu1exhwd0jalC2DMx8Ck/19U2nJwSw
m3DnSqoNk1ZiRh4zr+HiIo936CgxIlMcj63Jz9OsOY8Bix2s6jBDhdMYvxgkfI6B
mRShiwlQxiBJcjPempKBWeZCvu1bDKYiIQPNBr4qcoXIc9UyCoocNE7Y+E4P8Vad
X8TsK9lhJyRXDscyp1ibeX7LJK20ouHZMudNvyjJSNt4scXiNQCjwOzKVUxYpmam
nJsCH1k1rBJfCoYTd/cPC4dUBdxbgPkXh3oocr1lexBX7Es8JpWAH6w4sxDus+Ve
ztkmq9tBq2Wev+lq6weNMG7NuAtZmsAXJuxwCuEdY3xKsUVyeUIGq9p0NsJH4PIp
0KvjLnpmWbI71Fy+5VO0nMR0WStQ4GGY9nzzPwMKGnHMzz+A1lHrBNushfMDq5KN
xCZeEqxKsjEgF4TGZG7+DiiADq25LJiNZv2/G8/h5ErnQUqk0IsohCge6/X4WErH
/vsMGLpmXlT7Is4CzT9VLPqlQ9xuBjewD9cu9WGP+RqCeZb1qg5x3BhxqnukifGZ
d7DKN5JzNi6nmO1G3Zy29GuuKG+77XfDorx35IhixmgoQ09BbIdck+CX6uRZ4r5x
BMW/KsFJEEqqvyO7AF/GfUVTwUStI0cSoUcTHaUcTBlc8x3QEoeo07LzpK2pOz/v
y4x60LpMf3CEJiexSVnhZMiAbk1BFqt1nTGa/GY2tcwXxHu2QsQitUOk9aBV5gW8
FvqrvJ7NJXZ2piVki0uVMBzCNoIzUn3Lq5UI5Mjt4szM3AQ5oQiB0KRzc9UQNM3j
f8K4sijg3KXbciO2nh8jhSY2WwFSNgR/SdqGVd1HeHaxtJni7aeqZ+T8ljM0pQzY
tDdjQq4Xwh0vrP/yiSgg2x/2Ov3N6zuU4MKiOH9B0goBnhfZnHcOf7U8L2SufvQG
Hxrf9bg/e2PITab75s58bE2Qrm6JVxclChx2MLe93gTLtL1CICJD2bo/dC6OSVm1
+ZzJH81dqJsCqISQJpxlIykCrciyN+5/dUNBPB6a7wW7Ub9uvPLal1qZmytTvAyM
dV0sfdgldyy+p9E9v9ec660H3SP5S8i7dt0kyvRH4ZkdvfoGhTnYuNTHpobmlcWU
MlE8pazgijmSYVhsl6+0lcWoEPoqADt4ZQguYXextK5d2H/RUTJ7uFbgwjZGcFRD
+ajS5uQildYlLnFUeGzXizt8ygLq+kmrOcISiWsq3TwWZHmJSpnJI8F9ih/0md6a
wtcjyluuxn2T/1Dr6nFJhimcNGRIEXsN3LOVsO20aQLEKKG9ayDqdWUV+YSgFMan
ehjooFxID5LE1bJR8503sYJBbw/bdGibhajlLG/MkjW8HOJCfdCGTznwuVEw4L6F
1l/yziyIEjboeXuZFDOj57XP32B1hnLc3/SatBmmant24kvG/11z2fpSAWs/2OZg
sXz86Tfv/mJqjke9N14+Yhvhec4VvKfzPUiHqGSxkbkxZcyYiS8WnsPYJfPelb9c
jbd5UMn4iIFY76QxfcGMNd68f3pSINhUtqEUxgbdcbLtBI3P9QBSIxQyJ7PWoN0U
ayTL40bnyQO1k/0klic3bsl8Yls19D2RQXp7hHRtNVLtXapFxrQ+MhvAJ4az4dVp
YkSC1OkJKDBG1R2OfW1wg3KQl6B0HgXm1pzJm7jZKYFlygz1bz2G7MRh00A7aEVZ
cLSlqPYiFxRrtSVceecSr9Ui6Q0cqzIyvg37wgmWJxaaiQ6PnuQT8N6Rqw0CYDk5
Ao0lY06Vh2gXKrWgn4LzfUffVJbLlIqbqbg0/oWqSAwMczrzrvYOz/vDo26027E0
P0AbbhvqogkXRMKZhURJLzLBmaZOrrv/2LtrwWrpcviy/65tdy2oM+1M0uYaGx5I
R+ddjnrE7+ioqeBnA9viWXti6ddn9SXhVFXduVFRy2G5rlMjxruDxwy2pGWB5C2A
+S4fvpTs37VdyCxXGX71+sxOUtjlYGiYw6z94zo2xA3BWnqQveAwm5AOJYrVOnKI
T5wJKuhGVdJB6REk9Lvgq6vGPYLkhKeCWoOtpf8KXSD5OaEx2M9RPVm2Y2BRjipt
ONjLgGwxG9Kx2tDPi2VuASLtPynrJvuTXl4IL8MJ+PWnE+c6EefnzDRpp+TFKw26
Y/lKmDmCqXbkJJhxc2pRoHB66jzDx3pS+ZkrEnMmaj8lKNiH3+VBH4zZCZXwGa5B
cwbiBC9DAEUdLDoAVNXd7d+hzMLfkNPL20OD/4FqxuLALH7M7XAPVoI5Hq7FfrT3
QKLqcEWeFXLPA/GRTnApXiY2RjenDkq02c19CRrNFFOPk73ML18hIKKtNCRzFhQC
ZWsOWWNTc9gORt6SV14OXq5tFjBf5+1Kqj+9ZCgX+Qjc//tpBb/GJExRfRE03jsU
XHvub5crS8HuBexa7nG3o2RblF3shTxBt6W8Xc+ovFPi/ly38aoVPktKw8vnltdA
M7kXWh770Foo2uWfMoTq8Hz+YpmckxuaqBhXCH73T+oymLoBtXuPm4xoRz6TXPev
eDjIYTbvdZB5jDj659i+2y7dEvVn7t2ergJf/fmn3ag7kX4IBM5JZQ3uzMVaQ1ur
BM2mrKFfSgr5klr3ztSsR99iKwyCZmGla6z/CEzXpFB+JsRPnoHSZGAkziTPBHn7
HQF8X0G7+mxHuW4bfLEBsRMhUc+QzbUKsWKyOcB2dT9OppqmZyomducc7LLf67UP
TPAWZUiaaBsoUlETwQuUrqDZINP9drz8oWC9hL8iNZcJjqVjPKbgOocHMmzo8VEg
6P4IQEcCy3pVR0w8gwXo7i5wZtNxyV81TYZIeSkqoco85EcEP10jXSwj9BcFBSBP
018te3bF1rAACSa+pJg5Pti0qdZ5OZXlOUgkAFbIJt0xUinLIb7CIAKlaZ3ziXKK
7QrfufKME0wcGsVSMgTWZbR7/I02zmhrTk9cHsNU/HleOo72Nyk6I08xkzBurIzU
l7aqghqGl5HlIVDfAMxwrRR9aIwb6ffyD3MWxhVyqBJMnPhyJXG59fEtrZQx7dzt
rmTFdictuFL37ZItOFeVnjpWLDgdnenqMt8UJZbdoGQS2Jnu5vw/VMqn6rzyLyIQ
cW0TSPy3Wy9RqkdpYJB007b8ha5EGI0z8zRpV4fnwu9FwRm80sEj+dijmRZHRfJd
3S5WgC7QYs5CoWrURoV+GrwQTih5MoNtNcDdqIbrQe8C9XGmOR3bsXlKsN2t1uEF
uWB+GkXL5YSg0sP5x97q0X70ZPY9Y6kz4oGESkcFch8PA9UzVuc6Y64/NU3P/p3z
kSNJu2fdhGffsXa00J42Hu/AAjBzV0vmUNUpsToQvCJIk2hbOy+Cv+twlTUR5LCZ
lwcTZlvW6EucCGj48a3Ap1g4W2kRdHMdXY2BcfVktlZIpf1AXm9YdXZuFSwhbZUd
O2g2/Uaz6iKbjuVk2I8DO6eRpfS+UmetAgP9M6soJ4cskucPyFL40sHuoj34BRBj
f5VOGLAsR+xL0reknQxJRgwgCxnMrcS7LmWhX3744aO6Fr7upNT6/2ATLRHnHosS
3h2mbbxDrbov3sH67TPip7iZ/GOiX3V8yKSpw8yYhZQSPeA/HSJZqFE6WQXzVOwT
IPGTo7P+JQoAJzq9LHphuc4ZIFa3xyLxvxjtISZXMImqf+PJ+NXlmpIH6oYNxKjq
4Rlg+zJPj07BE4DT1gPtEz9i7igrOTht297koKNjtduJ+639XIVC2C7Gihg83i7W
9vIStuwI8K82zv1TFAa6sVTwiPRdb0AYkHxV2FNO9QmE5smvm8IKLsPNRCpHGAz1
yBAGtv6VWa3BqOey4Ge9UoanCZI+Fk2DKH8ooHHI+sMkb4pu8jQ/a4riGaY/21yR
QgzqZaDs8SBpdfnl2MfGd9ukLkZc2jOUUE60toNmPlrLJkgMPP2NKOOZ8iD2MCQ4
WBs2ZsWCFKfE152nha5s0MaHjWL65O5BuZ74i6xR0FIS4QHvMxpFy1EuDxI3K0q7
uBvnXpafXd+P/CDm/0Ru8Dth+AAYwD1FMyFLlnHlm/fJpALCHaQ8uvPheSO+vHRe
CRffAlDpk+/3PsXSn20B+AcR0SZ7dENwlrjKliU7ld2EFbU5KqWvavyljO6KDLbi
5odKcUHfMnNJ5BM/RggDe0kREy6BrMp7Jqb53YkX0kpORRdKQFhA2J/Nbdmotd0L
u6jK+kdfyoBHscCd7SLXSKClIYhvnUQ7LZtaYRYy75UoEPUT/aT691sPknFxDA9H
/X55iNFZk8C0ciT0pv2PnwE84GM+63iKNtTSLhlXuZ/UUc6eUbHUrJQ7Bw7QnRc8
/qGz9F0aO1nmH40cd9TExSZ/5nr3lugJkgUQTOgZQ7YnX6ew/wTarvWv1QcGTh5t
RVRF01oQYjZzbVkdcdWm/rqHeOxQKg/1X4Z2hLrwn0R9m/XALFYzpgCSpX91Bimg
PgvRe+zNetQKelHaEIBTBYK5X4d6xxK8ZNnkxYns6Bj6N0yeC9YOUllZ5YnnamRC
F4Kci7Baem1tO7X+NV7VZdAGJhQelsDyX6tK+Sx07rkSI0N8DmpiakDQjO0irMpv
pNVW9Z4E2W2bIduBEs7vc3TViTiK9XJ6SRgfBzQ+I2Gh5lZdWgMrJK+qWRwNvtdo
FKLmxprdwmMqQj4z1LPd9IZHdAS4snq8Vhe7RVz7DhZwEppXMfp1II3aGFY7Xymu
QbivkWwAIMTfWDuNj9FV4M1T8/UYDaKTlXtnJ2WtO0mGJc+fR37LsQnLhr/hm+DB
8vIXH87l9JvsYy5WOTUIaSGGjRvvJ56e7PYAK9ao575fjm9yv9kNzKkxzYLIgY/S
WfKtoEYit7l04TT8PXv0B/rTBUOpVP5CEBaCNLd+xgKU2xskZZ5zrP+6zr3BNYCz
p6fVhaBmvDDV2Lw0WzREGsiHq4BQ2ka7t877eqCpz9S0OHOmZm5VeKD02IO2MKep
/FAcqz0he0YEab6/IV7c8R7byXBvXHG/NSUvXVeb3UUb+rmk0vsLfPyHPw/nR58i
ZVqDtW560NGFQCa8qj8YWJc3ymDGDlu253NSNmzYMl+pkeb4CsUSS4E1mrz9XFTz
9UblAqq3p/jPjFqh+xm6/2aGnTFT7iiqSfBiDXM/sTZRsoQqKk+zpDePF9g+JTU7
1qck7crBibwyj/u7Obao1YQV+NyZDu8Ewk5E05l+Tpy1UZOZcfasi6ofcbq+50gM
HoqO6UXL/8GYzHSeSfLnXFHNB1/HXxFMcbBViGVqizPDM9U4MK10kPDM2VG5BYst
bcgQndOXvutGI8B+kOcPhYeQRVn0S1tsO7YIyVCpwRnTJUyEsAEuHNMqPYPcFOp9
iK9exIEbvOwgfqAwc2aigLYJdBJAuHXBzil3ghJvx/8gATkCbkEoz9p4c5rEefoQ
Nc+64yrfRBNKxjwx5tg/cqL5pq5OvEAct+GC6HgTFOqX06IqPBZiiOQ0/AB7tity
yAL2BHP+e6ar0W5bgFO1Bq2nGRj7TB8R+oNThm2uzUd2USvwsgL653YDmeStzkqB
tyS/AYWVsN/owxiTiCXoEot3tO4kvH+NVpKd63xW9R+rnEnuTdZOoVfoQq84h9Ou
6MON+vAupViXfa3Hil15CHZBpkHG6YTqLnzu8AADWSoE1WjfY7AW/O6P/BK6zvEk
5yFsu1AoJjsSd4vgWdJZ+7fFgZc2DvfzS0tL3oYnRbomsYzUB3nVaJzXAR2QG87y
fuzKhA6eqWmzaT61RrNUNaKzutynILj+U697gxNs7155R/MKjP3KGhsTZM0STS6O
8GZrWqGXIn/L3kQC0N9owt0wyil3gChCOaYpb6+6aIUq6Csaydy1i++6EkmLMhK/
qvCJgSkNC3gCbLBj9vTNmNUn81x5dZvJOBy8fynnPOPtRa9TgR1QUJmId/5LZv4q
k4pEAQIKlAMHw2oosjaIeUX6LTbvJy/DqN/ohmQGxPMvPS/3oA8VHmDb/IbDvDuE
zcwyefNxu2i96dS+Ndt8bkAiva0Rg3N8a+wXg0bj79pDfwD4NExztw/Nhs3BmtXe
E05Djy2TuBWEYMvckSLxvJlhepRKFe9ezrjKcYlxWwyDgmEmDo+cC0hdXqJU/UVm
elScck9BB1ISyq/WDF/o8gumcp2TrYTktBVF4jOixJV8B99XulD83MUPYvWmaKj1
8PA+fHzIeSKUbtMp6L7/UUgPUwpkCBczFZcSm7vlJtd5mxOYFEhIZS7LnuT/5sIY
TNh22npUBxcc2fF1mhW2bboBX6xn0V3sDuufhnR2K9zgggeR76OXx7BN5fTJCHVg
gVkTrqQS6G+udfa/+2Un8RdJj2LziqLvvANLDuHpDExz01IWlOX/CbGCJCNucYnh
atYX4lXWhv2QsnJ9Cx4d4m9e5aL5hVYSgbYxSKm9J0rB+j8xBgjXItJG5o2kbjvP
Hp4aE+rNqWKf1PDL/J/iN4v2GpWvL84V1oKRF1fQRhQYTERegA2W2cO+aILlJB70
E0vbiJcTElAU6Ek5ridCqXbZzetOw3Xc47ScTagMdFJAO+o9uCkQnGtAdKrAfziI
ZSjFzAABiIOa39Xc5QSPJZARtI+jcUhUnp/2m1SKii2F01mPEe4EWkfY4J3E3Og4
vtATWOTmCvIuirE+mw7r+FkuvbahNJNay5hYX+5Day9z8kOzMxCrwbGXhWTKyDWh
wtjpgEyIsLJjzyxf9oHewEf32vgPoQUVcR8Zm2SzM4vduc1b7ULnrbQkk1m0KcwG
pOrPt5K6toF4NWXpPwrhc/cNl2T9XhdN+MbXfv7RmJylloI+AFIsQCH9SAJD1OtX
4yGBl6ALhSSYmtjRn1opQHDIKvRFbZLzD1UZWl8dAs5h7ybMdL/cs5lTdM0xhWIS
mQtSnZ2TT1ksZtZPgEWT3MawZVIMkSN9hfiewkIPYSFLI5F1OYoYJBN4jYmLPryf
/8Hs9V/e/cswCrsipx14+y/vlIKyR6ksZL26ulDiYyoKhlTCrlSH82n3N40HP0Ns
0EOjS/cfGPP31k+z/TNlY4Wb2MR6PCVusXaDZRyYoya4nE1CjOTFOlyGaGFMQ7e2
U3g3uKVz1QjoEEntJkRotpVga532+HNKaFDAvIeB7irmlv+RvrYgIxZiTSko6/JX
ThHuiA/g9zxEXpvTg7Y0pO5T/xzj0PJlNqC2/+dOLKblDH5GKz0mtQklvh0S/bKK
xZzZ5SvIxDhZIRc0oT4W17QKwiX6AKboV3VX/N3bE88nV2w4tqqN06jlZcMp1G4y
r2uVoaIEtV9GEhbue2iK8rPkwl5RZ5yvXoW8eT9jf60iwjfCDe81YVUbYztiUV+E
MpQkYESYocRWnbmuGyf3ePPoYOwD7i+gIusnQWVaF+z6ztq9Qn2v533G6hW/5MgD
Mby1H/qyoBV2yUbpH6aEVoV0skMbB5ecy0FxskOYMMrU6KjQc5u0JMwIr40aLBld
ZepOOzpZ0TNaY+4q/xgA8VaS1bxuC7WLPiRyEoJNmVVehZOY5litMtTDDIYwICPp
I4wix3bRLjm4pZndIJQ0y+sTTP7Yt52RaSyCqcW76GklEdk9JlJ7CWjEDx+VSZ7U
AkJBNcdrLeYN0RYL9zcqC/EdARq+Ui8HvF6TbRPlUWa2pUjlHdoZWqN2XZBYo3LQ
0YHZ++3ODKFWrE2TNPluK6KeOs5hyyjtZK0t5cTxRcRW0MYS4tk7dm6hc0tnUdGi
S071XqxbMN07LCC0Va2Y8W/sSh8l4kxCmzR8irQfsSE2DUgzOPxmsBHi0gaH3m+t
tQE8ERFtRIkTXl/n/NLvu48/0Zp9R/NbHVLiYvb0vNchMxvOQLIyhP6+0mB3ccWl
PvgKjx24oef63S2XjGSmZXvNfjv+p/pP1c5MbMU6Q4TAuKOQTbapZYHkUBhgp8UI
s6Mf3UByAp+4YiI9i3Nq66F+tTs8KbfT50LjLS2fAbKL0VsL/+1uwk0Vkzo5jDnn
jjAIx1tU5ifwV3HXPwV5CwduBknaEUyf85RjnptLUNcXNCc0HBrD6b5FEmjOIsLv
p1/bKlazDyinQc5sMromFWbEDd5lc+sBW3UnKRXuRVACiOuNQ1CG0N+ZNz2zFJ21
1atdTz8bBXL4/sJdQ2ELL+rcF++DAAS1vjDLGbd1PbnG9eSwp9zXMF7ZPcVH2Hp2
XL4JXrclQMXqmbNKwD8KF4SnuDwWakaBbuT3VuMEgzS2jyLgyjinfFLbdwfB/6Xv
3spoXZeqmAe3fO2+Gg7kKsTN5guCrrOsAHiDgjwO13g65xGPZakA7Un9v5eL39PR
AoNcbLDdkSV4GQIdIWY5yK2kQYT2MS9AKtjN/py8ktq8CVa8mrpR7jTHh6RI/djM
/HZ/zn7blJvSQKYZAnWiewoF2QuB87h2FPJnGxwxrVekjyky2ugKk37rC/OOJoJO
uwRcAAoN1PFx50Gda/bjaF28lWGMZRhLHblYXaKI42Ifitk6Hae0LI529Syrx1mp
kX2ne+5Mu+geIBvO6CwlCQwq3GqNkhI5kjKvyjSZrmFQWeI+mOqmPk+Nu/HVYT6J
y9VyCA0XKdEVp8DM90TnfBrTJMFzfx3jxWUzAgPHcjTcNqPM5GU7pp1WGrTgd+zG
zdyTZuqyz0MaDB31BdK5iEDkm4gReIYF9dcUPmJp734z2mLXBXyWPUwWPO9IDSLU
70nMct+QYXImWCvGVU8Zo0DDxLt0aOQA45NgKUJEfHajv34foEl5Hi4LpjWS0vSI
uLC30bgF0kRnDL3oVFAT0dbK/rq4O1rLf2fWPJl9ZD7sSKgny1iJrbFFBaGSTrvq
m7HxdMKpUoW7Gw9M36y6Qv4z/pjLQ9iKFqYxzNkAl0eykK0nBPB6hSiBXQII7L5B
rovPpVoQ7Y/kXR51NCnKXQNEzezu931g0rFrfoWzlZcvbcAUi1rnd/iTUmKHLrqz
ztcE6QijdFa5nuV2gZMYRIF+E82rsLgojTqf8al1ShXCJ5IIqO3Y9SfNuNrpEBiJ
wFKSAfCsLE94p0akKxDEawfOx6+9SajBI9pee0iqDBGOKp0HZFfbhiNWGJgNnWe+
pww+V2XBCyzuyBx8JR1BMwlUhRzaGdevlpKa6vvrDk0MGSRFcRDNu+YOSFDKtTkB
yenJmKVGj2NnYyNHCDtfzwn7OGBIlif+t/zVzAOVBmAQL/Qa4+6dl9eiialx512M
44jJDLxT5BcG0xYhybXsc/qx+J04jPn+tBIEHtq73tfpZhRUOv9ZiBtGoGgBaGEg
ROwK61TqWeYYENoqZoq6KuLjz2D6aW32f5gzQV2ZyAd0QWFxuJjPaIAhZqT/5k0o
6WhSx/hHj661P/IN4K5eop9wyjl/tqCwkeKSGNU4SDSf48ZYMDxGX7RNbsfimM0A
g18bh0GJVyfAi9IYBelr4YzV2YB4gEge/YIqAl46t3AHk4WXbj2whHyQQKISILGE
1NCOkUM0zc5Nk1CLupmwP87nBVc0Zlzr/cviiSa5FUUII87gZT3WOJwt8AOLI2nZ
EP1dpPFUXO0t6TdBLjalEWBSz7a0hO6w22cPeaepSKBu4BY+B5uG+ps2gl9KOhtk
UT7SV2Xk2nNGYJ0ywoDMMAk9oFcLciY8ZQZVsTezudjfVERGuru5K6LJz/m3l2Q9
nerout/oUnqLyFreTFWyPg9gtIde3NSi1S9w7V5fFcUMpzrK2+072FTsPzRYhbLy
YxKUKNC/QA/logqdbITjLO8Z/ed9bL24hnbbCID44Sl496A9m/WDCRiHGYHqbo6N
wauMmPO5sYRqm89bdrbKJie22SHJTxX7UFShuqA5za/fhhsY1V+z+d4Iw1q8EnHQ
DqyUWlsCz/MDvrFLcVaWNfRIZAGUBl5UxS3R6TTNfKiX8eOq2dzOS5mwBmqtkwaR
JuvUiZUsmYVXkBf4S2aERwpAF/1h+7UWV5evlQ5Ng0y/ZJjejmlc0yj8OvbDeJNB
DA7m4XhlQP/r9wgnLjomxBSQyirVSbXNG/h4jQFnP8dCah89hf3/KnVNVo0COU7H
+RTYjePMhnpCqcKSTSNIsVPZLTmcsFCjoe8lR/E0UlgSy+w5KgeYHnPUYBSO5J2/
mou0zflQwKO0DrSCZC/2H9kiM8vRwsQIqYU0WhbZijqwzjRTriZ+UYErMwtbvhXV
aeZuhHx44ClePIuN50tRdWuCpzheWW6W7k65FrGii1tox/fzAQRMu1PS4xIhOjNY
11PdCkHV1KLvNTcryqzJ+ZhpW2/lr08D5YBcXY46vTKViclSmpiqz9AjYYEMfrW1
wRKfquDvfWA5/4BfpKG29dgW7DIMfOyzms1zQpMTyM42gPcy6PQJl1B+eQeRmhy4
0RCgCmNtPY2E3Fwlhl8n4vunGjXyYxgtOmyYBDfDqIp2gzgD84FF9jNoVKizlrHU
XPBwjWPmhcjbkBaTk37gJ79awP13Xe8ziLEWRVDjPW3zUIrlWRZhDsoSWqYs2C1p
2PI7HWhwE+BE73b/grG8ILAIoJka6Fha7JI/8NbJXxbX/LxySVMCBULvRNTX2GtK
QvDaxyxdw3GlJC+os9EsUnD64OFBlVOvtxM8pmMG3fYyAypOBMFLpWEsQB4dU3SW
Y+Fs+YnEYImsm92r28ShhhiljkT6hx+fo3TzZa619vuYniXC2skj3IJj9kP0m8ka
J0lcJs1r/Pt2HGPVhE+Jxu4T3mJFyvd42o9UoAwUuh9pfEwBr4F4unK+IjaH8v/0
wIvyqLc7UEBmEkH40QT1MS7lgM2zncystGHi1qiJeY1S/EJxFhvr1/raAKN58L0I
ovpNZMERSNutG+Dl3gqxP+FQvnSoi1Ih/46RS/2F+jcdLrq24p6WKgdHxG2/wKjb
/nS2LMXD2qXx27KyRwygCCvP95sE+1hdbioqtW1xb5dRs5Lv1V8vtL/KfVOqS4/v
jq7iFN7ay9+4l6wlorETpnJGO7T2cnT6AgK8EfFjrOLy2SXP/zfFsFWOd6ObQDOq
Z86QeiUsFE0ublH3sH9qEKAQo6utL0EV4F992kAnYK+kj9mhTDMmf7opkJtXJxQc
gXRSptRrS+NQW1VqL8Qj2wlw3Og/vZP3DJiZ0u048aNZmSqie8dKzerAfWd6u52R
w0WwLi0SlwTxYErLq5dBM1DO1ASSfcM7WyBhrlQJ9azlcIsfMgIkQdQIwXNSOl4N
gTRRnkPg7Yj0mWjuRvtX7taSpjOK4S4QnOxsMegQ5gTuWVS0HCoRYpIzcu/zxFM+
/KAOlrq862QuFHyK4vCSLzukbZAxSwYRk8i5FkMHDV13PoJ+vxZKlrqnKdSogSMI
qutMOd0oYrLHnqEnWCPSxzqccCQs6F2t2d4cbYW1FEzPUf2roMX7lsDE2jZKS+dy
b+dQZmoIvS1Kpkw+vD0UqcYmXQBmHxM0chSRI4VMKB41r05Htm/KdFRrAuTP5Qb2
Yi9zbpetV/ccay3HfJa+nz80M14iCU0BtmgBpTBJKs09ZXN4ZdADleLgJ6ceoLCn
iz6Z5qzuj4H7YmrK8DB/bElR+lu9sjytTK1Dqy09lmbdA3tHmhmEtJQLX84T/4Ew
8d171dsyMeTe0lAtFGDzcOhMDbcnJxFywetpTs+yYW5jx0lJc7o18Ev2B1bADX9N
YK2jgVQKgTt5SuA0wTYJ3wYG+MMNw/28Bmw73gwCiz2ntse/wSLK+kwrnFEG1evl
GU/o0ZUrJLkfZC//OuOrtmPipaHDrDOyYdd4v3HZMRJ18TdCILFOLwiafy9C2u79
b45JNxwKgmUpGEq4YvOt8fIEJcH48dAgqfvHVwc3+ffQN2QXoT+8UXtFWbZUZrcp
0dmZebiS+qIFo0DcL4g00C/8Kr+iQSp2bDbGGuQuULKxlUAJ1pP0ou1yUZ6QxMqe
P57bSyh4abtEHhq8KFtGUQ9FzLtCLWEQbwhthMWhdeSVDxY/qpgA/TeqCXjIbqYn
djeo1/0hO/Gnc0tChleuoB2D/lqgSMs21ILlBCpQzDGpHZmPQbIh8sL+I99emc8h
l+tfIGNw3Kp4Csbn1iyD11oATSuVDQ6BgFLykdZiW4Za9iVJc1ARdcctV5pIDWaL
qucZslXj8si2xLhI5dxM59IhFvmmyrfWPbU6DwsrDW97/m3OCgIexdiDaH22y9tN
/rI1cMysLao3c048MqSYp9KFqC2RsFiT2Bwl7Yjz5Wu0BNdVXismrJW+DSvK36jJ
pqr3UyqPAIZLeAykOSTEEWsWjE9IibcUgqEGt7IT51ajl++ZJzFYdazVhFQyfgfA
mVAIOx8REOpYAAq79Fri1VlR2O1jOeSr/hB219332HDfncDg4cAOTnUFiZyoqc/R
DLEPCyp3c12UMt2bmaDR+CEMJ203UYaWcivmCdri9qm6WATRv25I1K9Te6rot30C
XTyEXAM5cKnU/UgepZrB/kFN8IV/CuEP/EK9XGpl36nH5VMLB45AtsnQaWjn++to
io4nOp1Nv5a49bsJxvrYGfWVuJriq1y/02mhgiJURxP2MsvUgL0YsCqy9T59VnaQ
H3yE/tjknzQBdMdU+SRHNeARUmfSakCTBQnRChRZdeTz/8r7TZs4zR2DogXvf3do
XpLq7tFSIzI64cuau/pvqH/DaRK2SSM40Og5/Ev041rWARwzI5U4Q3ZQboFKBbXC
QOYew8CfbrQobWicY4amZpcGTHuki/C32h8dKCGFgU5nqMLQFKgTNZMp9BEzMEvb
MXQsEgaHQ4CQeV8naxX140mBVf8SZ47KE2OyTx9IJolE6two147vFKkCCQQHHkzs
lr8xSwvfazLmnh9nVZt3Nr8I1ytS7c2VjXqPqOEd757aHxv6fLd03XP1Y+1DBqZ7
OXqlIRdZ0laTtpBNypmcUtLecGC7x5la4NsstLaH+Me5vTIc5X9KobIYOt7AMPoK
sSeHfGFvDm5GjgJC6+Eu0c1+evutcQO1VzZJ0Rx1/jfE+ralog0JssbV9Dogkn9G
4VngI7Ayc6k0HOahUIT0ZfIRRR/Np8tzCPoJLdJxTJnlH/wGt4baN3sAeFhS+ghQ
ENgUE1stSoI+E2mZKrdySjRl2pLbuHUmXinqeb1ZgJ3767erQZCYh/vYuV2deZ3H
jpBJmlXzvZkX6Uq//VzQfYdqwkAozvdqbRSatcOY230yUTcjuiSE1+04BCe+AXYK
3zMz7wcyYFYLOwlgOi4pAde7hgTKA5yLLF7bkXEcSA1GXJgtrBuSKJMzwiANFydz
EgbiX4Q1hsgI5XuC1r1/I4XMFIFkZlpepCXwA1Pjyfre59da9YDy7zCyVxSaUkZi
hsmLM8tivf824pBTB14+yIxf9ZlTSEOYYscdkrPcPvULmFL5VG5pejrqLFze0E8G
IgwvMKYMtgC+HZcaMWxc7V9ZzAnHgCIph/AgmreIFUEqkx1qMiU/ZO0MT/uN437L
kVS1v+dxglyEiyOW+PqJew+dJQP87PKfPc1wxfbzrom2azStn4ydlyh7iURaee1j
NMM9Faam0751QAWYG8zfqKFpttR0zoGLkO6bL8330w/s1mjfuoa6rJvJ+/MsiPgJ
IX8DUH7ObD3J0qDmj3P7inGwIABz8Gfnr01hJkq8DnSNMiwb0Oshi2CKPFaeT/9c
pA8I+rxVEKcLkFpaz0fyECZLFICa3xPUUvofe3x2td0AhXTYOnX1Yorl9TkQZJie
xocihCW4cRqlUBV+gR/vyD1i93uURjkwsONCbLmXxEYEtLAO1b6teuW447bSkTwZ
/y2lziu0jTs+XgPAXTeWvV8CByBoy5Mx4g0kfoOQLLe/Pl+1a7vD6lgMVjhtAJD7
QLuQIfB0Vzu2aYeDN5LhgWs9kp6efIOJCvs1nv3srhPBlG5NGp5DIRCZ2Y1lwXph
Eyv9jhpr6146qCAKt2PbHGLPqzL2QcJ1E7jEBxb/+QQtTd6PtP5WB+0ZxXhmoptt
adXeJ/UzGAZWnlQEztxewUi6bwRknsacU5eUgfQIgG9FoxcrRz7Xd9hX13pBgjTF
9FEbJ79KhtXRGOXadzFnu63gh449MNhmeZAYTa4LwgVrOPoyj3UnzxSQx9/rn9Gn
C9Eus9+j4qFpT03lhdovdkklswh5fIloXqlt8x9NClxT67wzz4S68AeIdEV7X0Q6
6OViV8Ac4t5arSDlT7NXfB+QFd0Wh4XTfmivSZP3pHoeZM/D2PSMkBpjejbxAnar
Dpbk7Z/MCl2YIwuJEoaaX0sp7GlksvZ9++3rsX1QjkQBL4YLZcTRIXXWYNuuvRY0
TzIoYpUreh0+3rEUxQKKlIb8c31sCfP9ccZ9XU1MAp2d/BDk4RarAjtG+3IlaJd4
PLCenvrgZzeYFYcJ3GvRDhGYC9zWl2DrSI3JpQamuaLxxDZHTHPMjLcPh2Wq8MKY
g6m3uX0R9aTDWN7Go+x2Ao82NzmO+26dhl+h5CZQNuIuL1cTh0OG5pnOnhAyfz5+
CIvyjkkQ/GNRi76lpK0dkNpQ7iSpYxyhR4T0t+BzWQ0l0G9E6w0GuSerRYe9tp+P
JP8EaPNmMn5C4teegE5cIBmLbS9vK1NV40wvLjFeMNqXyMMmIdNzgncaeykSS6Xz
GIBXuDVXsaOgEZcZ/aotJ/o4p0A/4m4SvAaNmWMk//EFurthQs4AJOjVVleQOSfJ
k0acDTsPPLWl1GgcHs+hMI4srgtmcbaC7Yoeyz2nd8SqivHaNsuBchXBjGzdR3Hs
ocXdN6VT0rd/xBFb/1ICwzyckxAjUVNeGwhZYgAsF/reDm0Czc7pINqrKo+fiy/A
WOgWsMIU1RCx+FqzGxK96WgQTdx2au4XmNsNrmh9akAKIv019vsm2u0nMiDDpd/2
mFwaGpiTWJGVl2YDYO7PG88G1K/lF54DJo3EVuBmvVVpzq9na82LBixGPXCQqXyf
6pEn9M/Z8rr740DwGzBgznd9KuSuacXr5sEumjRqBKLwOOJfuNzJc7R8WCj93szJ
Vs8LBAPeXNKQQ6mB43H8fSkIg4xqwfvlMiMNteNIhhJN5lFCdhyIhy589p1BKHJ8
qnfOmxR2x4gmhdzLKpWLwO+Q3TzgViz/gRqbfyPZcI25uhgIc0B8//lRAFKPLAPQ
gFWiypz/KvsPa0ughMWqBIMVxCsVtqsvvNYS3B/uHBlFOFAX4hppzweyw/ky2wCu
4Jt3I24f+wfZo/xY0rn1VJNnTg1i2rsjqsmTaLYjim6O/60tZJxum3mbp+aFD8Ue
csTVkbPAulhuodyzUe9ndJhlRECgfWlW6Y/i+e9LQUpiFJUGwKjr7Ivka1a7kfKv
KMowkV8OiDee/sZE/NcWZVKKvODEdm/CrGGRfEVxEUd/c1zl8Y3qm8aU25KgAV+u
6Q5FxWjGZ6KijCvA/+glwPSSu1biwBEJxtnerJXQqwT7cXJPLkJFf5WjCtkl56lc
Fu6WBkNoY1XzscKIlqpjAdu/vJSl++SGA1zpY7c9Skyzzlqu+pzi67Zv1/8416lQ
SvOZxaCoFxwY1f+vte7fBztC1DyeELyISqbiM9ymEyF5jF2SRRgOgliRMi56ZEWp
AihK9pItGRLmZOuZwuPgXO4n7qst6oSzUbQZHzwousdQx/XEvGUNQ3wf7ifOiTDd
lVohXxU4BG0HY23X8kwOq0jaWPkJWFzEHl9hGTlC4qBWTZiQWsiBLNbQ+Zh8U3oB
n/s06Z48fvbaQCS+sl8TFhKRHoZPcl9qeAGzhNmysymZI8vc6JMEr9HYbsF7FZ3W
5SjtZxAw4J8zVFhWAuD4wUGDvOX5OYLnwXtycjnMtrXNEWuDnD06qj7IDUKRYwjB
0b3FMGmNxg+bAVUfXckoDaouRoHgnYM5G+h0e7t6HXPYNHQgKQ45d4eU7tO8XVeR
Z0cf5FhYS1Brhs9v1/gVNC21M1Zsr2FcI4avtEjt39OTxtfR1tFRIkBBxODHvyXZ
GBxX5gA8FavTfr6TC3GqEAmsAN8Bez8pu3WOkfdHTk16OOzmIccl/iYjzFLnJFNK
yx9H+1chGnfH7EiuQtC/1EfLJ0crYBy8ptDDWwx4xZh7dOLCiE2D2+3g6hTJW552
MsGia71z4zCof4GCa/ikmiPTWjZeQKF/55BZHjp3umRWBnB2X/kK4K+LnGq0ClVw
oz7yvKRbEPfs9pWPLIiP9JaAP+H/2Vf+Sybh3Q5qkh1DjPsl06mipe/WC5uQ/9w0
UskavsdYOzwKbnQnOsMWfQgzXWtV76BqWePkR4I5CL2NyBKPK6EmNR2fX9Et8I9u
Xgz0RzBt57LT9pFhcyoihNDE5zMIA1nFYZir7obPjazErpyEESh9G47OAZaTypqC
j5Q+7KHf2Qo16JL1IwcYWGbO4aWnTcuMqYXPPa6mWVlvZCYeaJTH/XHJFeZrxm7X
+JBi/GIuRyXYQZ9i20/tziwkFBKMW/o6m7sPMO1LypCJKo1oYl12oZn2wvOEk+Vq
gYNAqUOT3WBhua5OKKDg1X2NPOXCbJZcmEv1WJW09at1/Flf+Jd/V1JQ/qEW46V9
5b3ENcTRX5kHjyhSr1rD2dU/lcPe8RpwbIMYiLTzndtIlKgsNeBZySFKLx8JNs1r
22rGx75GtcbAs7gwCS7skZCYqgsBFBHSX8Qh3mck9BL6M48K7ySMgeXBwg7+2C3M
DZYdhlojvsSxdOWTBHcWUqY6STiUyiGQiMVr17ckMIAZ6phdB0fZ4M1D/evAM//d
gNL7yLhdHTkz7G91eQtxsdBQfJ01xKsOK1KWqpwenspi7MbEGJcNbxkpp5ujHcTu
9NJ4pYDO3AaAsvPhcauyxU7A6JD+QBZCaJX3vJP95YYk7rMkJ9jZrgUX82rqokx6
Tvr4OqhwGe8La5f4k13dAU8hAwEKA/T0VmfXW6wHMstsfKxRpwKn8PDmfNmhJYa6
qyPqCKSYvg47iMvT1uc9q3i8sKETy38WezMFiUX47EfCZKabNsFvoXVPJoQZQJ7r
H4XGg1wFqVwTU59R3XU/Rr2AWHyt5sGT9U7IrjQKGveryc+tAqYZcq5G0K0QGJlI
cxEYh3MFOdd6QXV66vV1hYV3666FOKf7AFMqL2fHVQOf/Czah9UuRYAMCCpHJ9Nu
0KXru2YcunGGXpMRY2kVjYHHh2CX9wbsXJb0a1h/RVMufBeKzOx2RanHb86FRh4N
Sz0TSL+2bhI/f8ETI4mNf6/ZPQAMnulzJ3pa9NNjj/5FCuz0LJxJuC7cAzyPPT50
WTtyyMFFRzwODZcuffEQf0Qwta1/W0muUGooB2wLEjGMqaew7vjZym/nOlMVTRKy
D0sVhnIJlUByQ8u7C+62LwRvSrzOVm4sNoCpl1eU1j/wW5pN1qntJAH2pMMxYx24
sdNVK2Z8SVH4ND4QvC6KGF//FBIAjoyjN2YdwB138Z+7l9qJlS4OK0xL3mpfjQws
sx6ECS+dG0kmSCv6eTLVeg4ubrgfA8GWNb2Dl+CShem103ZariCGujT3oCSFliS+
tP64s/Vq2JEHkFNhrQcanWTkDZAsqo/qEoz5EWpTnJ8GTG2QdOP9Dgvb0Dv9vJEE
3O5D+R5Oa4x1LNRuEZBAzjy/Aq8MRFX7bi5U89hqJRmLvzSJVABO+EhMcv71EhwW
jHQNFK80rzAumD53qrZ5wBsc51VRDVvhd0MV9dXx37JMh5RBAbXe5sQoV6cn0NUY
3GfMm20azp/tDgiTMTUrdZxO8dwaQBU0gDPP3VyzH0lFtdH4FzY0J+kYCZOpM3GK
2yh1MF9rM+HWeUmsXoQ/lbaOMz0zG4bmPycM12CfIMm9k+s1GZJKFVGQbM74WhRe
iHjconfdHHPkiWVYwW2h9LLhkJUTRWTgpXmb4shPdSBZs+wSWWSQnkqIR8U3w5pM
RQidg8TW92mAIePjryb/9K5Lcham71dy+VknceOGWVO6NtoW+unKv857+MQPcXPS
lWA/M6bmzS7JGXvZOSGnvjlwCxG1HS4yECSk10tp5fiWgaovsSE1gcBTyiqxMZ54
2cia53VYmZ6fA73mCYUP892qc+zqVEW2IIh/YQCWqer6Dp/d9Y4+0KLU4jXov3hX
u2TBimcL8qmbRtEbNrK1Y2JbYqoz2coYYlSJ95h3kMJgV1OgMlvBsOuD9gWrpBQI
4QRe1Dc8obDxQdRAbD5dANY08V3K3mvFSuGRDnYEu3/R2cqu1qnK8/0mdbSlfHak
oig4RTnB1SpJCgRbYefAv05e0HrRvUUEJQdXQN0LVsGzV40GusBRtlgpJFDanCXx
+rT8hTt3VwBNQXiT6eWdymX9YUELfsFg3zxxNANh/DIZXCKC+yXdYXRZ28szYlH0
Wv+eTsltnPVKYmnBBB0A5m2JppPInmYAYZ49XltPZl01a/LFsJrCQTkmwnqSVUct
/6GkwwQreknVLvBxQ6xMjPh9w/XL/DsH6KbPrcvgvVXlAJEAkLq7v3atbkWEueBL
L4zipW5kzP4XVF+lVwysQ6S9wKsWj6TwrOfVD8a7CDsBYkmaNxmxoFGmdpKNx03w
oixeF5vnhmc6M3N75jq8KFdwHbh4EAtE7uWkWZA2b/mb0cvKCMw6zjXYnJJRhRa0
wKUeUbN2vFnes4KksFSF4GBZxR/jmRKRC977mB/Kwz0g8RRKt7ToBZTBdNLhdces
ug6if4T4u+kevSFeq7Dcza8eZK9G9LvnKTqZWCEy/Cos1ayiNBf10+xWf1K101rX
1d+x3e8ShcpA+efGCkn3WtPs7B+WTJBClSnQhFcf8hXboYbrJkOv73Ancu8di9N6
avX9Xwmq3nbeO4gQ0FHYeTZSsc7jxw33vSubygC9dpeppLRQAGH4fYS6DJIW/ZoV
UfGTIP9KRAP6Qs6DJ+QGvrWV1XFQjRDi9t/eHgT+B7HHc8PLdIRaLVycDHwnOQn7
aX2M6VcusrPnFfCUPKeN+2FK7cFIyikeMb36+fId0A2320hV6vyU9lVxqAx+nyJ5
hNMyQxq1gmbZBUlMFVCntaBmPpZmvlaHhs9bjW/wK5RJXKdKNy8kXPgkYxlXCAIW
rSQONMfbrGuqc9+m4M0ebl+fZtZxzA4lFj/u9BSUm6d5rlwL6myJnlLm4GMiXa3c
GDjZ8zh646/XnylPRW4HUoHc3HYZ8nXLW/uXjdXWjBTw4jjYNujFsA5BWPvp9LLM
npicMp3ok3Zt60W6ngxemoVi2NIkkyMRaKqHZBXW7jCQ438NRSvHcfUtX0xW55pt
K6/mE1zZnVImX6UFV64cCkCEMLgoVLQwy4w+m/TcBs+6ahLALPXmkDa2oFzgfJXa
hFKKCrifqYp0ydfGYdySiSf+FzZf+5a4G0dEWcJGMKWB2vroILAUNAZ7xo4u10Sl
XHEhBT6cr4zOX3WKdU520HyvAQ8ET+EOOMjPI24BQ9O4GAyTIpBjinVHE+oR7QCS
/phyOZs/FY35fKJftum+yjlxuzsJCMyIacLYc4e4Od9C4sjaQHwhA+BCbGjFJcwe
aQzTUI3ydaW0VSABmvjFd7txqpnfhDeMoWI85EwOYSPB2QYIsps3XT0dQs17aQnL
0zqe/1jy7E2kg+HH3m/NFWomCi1yF9Ag55B0CDGwvdDf7yT7Vf+oke9ib0NR5Ndg
S6xFISvL+6mTamc0ql2SoKCMNoMeHCAguJL5GCpF/Gaa70jQIy1yBVxT3OzNHeV7
aRHoM22bVOxL1LjJ32YW2RZX0Zh08tRVeih74aX63bMKxHb0W6CwDWs5ictsVxFW
3ozyO/jkWwU5M9vvpCggvKgljB5iGSf3IePl9F3KsnpIRW3VBgamQSdJMBzJEExp
tgdFig7+1kbgIU/zZAgNBDeDPg/22L8660EZiqoOS+FtzdkR82HeewQlAChaQgMm
qmH0gEdlKrc3Sw2PLfOMWLCpDajgip5ZwM1oA4hei+UQnXetVGQPnajB2ynuseub
tBEDLtFL2ttVO5w9HL4Z/VHORYMrCDMemhFA9Ha9l8pMukx19xk5+ZBj9iQaHn1n
hj+GaCEVBzAgshd9eFUVtVJqlAYK29EW/WLHYyxHq1/XqDDAmsU+9aT0NOxRWrmf
E76F0frDyiJTSyplhckjyg/yilbaKd05YmiL93V5E8eRoirDqAkDrovcW1ulhuWp
/8//GUhxK8Pgq4K+x862F7ZfADdNcr6EAoEZ5VSTM3voR2t5hbUr8nM3hrhH9QXD
ZEaGUWqVugdaTHMkTrzgWKhLaUPwr9LsI2jCfHPx/i6Hg1ztecSYCl/2oDRBbeWC
6BfCSSuMHTLyr982kWENLuYVzwao81zk9Qf/Mnv2eFbnfIh1egZNPh8tU1q88ZKr
jgMXrQrMYg2JVQfATJIcg3jYBUEvqfaJgkw97vkMAMqr/9xrUaAWOcdeeNpeCBn1
Fxq9umsM+j8NvOvP9tCyPCn9se9NG8yJRSaOz5gGDdqt3im73GZDKbOELuSm6keM
MkMI0m9Rn8CJNACLMcj76M7T2ZTQQM8DPHhAdZu7yZVB0JLu35ffJxuQuYmJyFpY
EMR5DR71tvWKTqkl+hqPuUvsYdvOoPXchXhddvzXhBfQ/kvq1A8//LFy3dXmTQFF
vkYOU4pFIEZyvkG+6T17dWrFeAHvGzxpQ5D7UakOTy8i9vvfSmW2zDFHDWpA4l6P
BJh6Jq+2hmNpdgyY2zq8+DVwEZS7QyjDOHBJDQuT4pE5CnnhGmcj+bDQfkTAspfr
8lwWLlQ4n7XvwW4UI4MK8H2xw2Mfp46uoiTyTjHMNzs3R7CQ6gtR7+wXS5+JX1YY
ZV2FFTqgYyZF7cyaPQph+/kUCFTn5FBxr2oxl2keKZ3QaAGZ2p9nb/t4vm7tEp29
+52lcJ9/q3biU4IaLQE2UNVRRdibIPvf8YbYIetBcfws7aubNEWhtoZagTzOEFp6
n2w7OtQh3gqI3uZ4rZWm6O44gLIY/O8/rIapgcZVWKPPAVRXper+DoaiHLa0ulRn
O1vYeCH41S7y74xCbMkuBrQqnPz4e4oXetXbGEwoZn2G+W+gZ3A8NiS8hq0W3bhF
6qP9y3ZrYFjQIa87vQZvsPLHgaVHYpCuwso+o/qM2mdjZv1c72RZaUPsCrXjT/k4
lEpk4Lm37hKQp1zsNiCE8Kz7SYxOlQKKT33fQ8JU8oP2y6Kj4qdhrm4BfRJWc+3c
KtWpE41hVZHqYspKajRVBtazt2uFUKyzaqA1YDHvB25TFYNHZr9X+6Ds+FazhqRT
nTKfMLbEcQZhEy9jk9nLgHCw2Xe7hxEEz7M8Gsr2raUDHACGLfQWj3kWboTnG+yj
wSmG9EihW6qY5J5jkyG7cEe2U87mLdRFimSonLaOYD2R0Dn4cClmYyHaFTUEy5jq
Lhdki7HnacLn57nf7NMlP7vxwGB2TNCytd5g0CYoabSN6zo74gLjnrTqh4eYcji8
FGwMzCbej6X30WGLfA9tvPckRSDys+qAcBKVGwK+y2HOI8hhZGNfE56Rc3f0xSLn
GblXVGxthb/srV3JUiEo/gBq176WWIX8t3zR+1F7+eo4QuZvIwXiGoo5N42zEAy9
Eg4Idwk5B6k3nkFqSfGUBS+D1lWZaOnpIaHfU49eHtGRzbAUq38cJzx1LdnmnB2p
RXxZzASvaF84uNhit4FzLl+bNmWRC2+ppj3OhKgxAOcVpiMBPzxiiCe9j0D1kqSj
VDNUc0xWTyBUi7zUZh53nHunQkFs+p7lg4Fq/LGY+cmxSyItCG4RQZ9j/HtUaA0e
KJ9mBdTn0gQWHTxxKZ5Ql8bgUtEmMmXjVkfRc3iTnlyphEtApZEhSpBsi8RhvaoG
DFAP51cNy8vLlMVEcyPvUf8IFJ+vVtpWICNNQGHMsxY/xKgO5We/qFXhsvQXzswE
IoVYGeBsGVcSEklzTp4CefPlWO3J1VlN/nbX9QvICv+/Bu1Cl8YdBgChXT3hT6Hq
5GMUdmf/B8ygKRyOKJpbxPpA5hZZ9cqN80BUmWd/gq3uXO7lsRZMKkwiS3vXzwJr
3iH8xNP0PGROYXXuMncE4paRIzvX4E0Q6wtYhJC5yOBpxh3Gj2sb1mgBggPykMQy
Qu7V02jZ1dqoPsCQAFjG1PalOFxpqclEWCoNXkbyuvljTgqwE/dXSmU50n7loIXw
4iOEcDasOKMJNX3zh3hKk4VxWPoIMTQcXmU9V6TXpo7NaVzc9DvYRbArS5T/xcY7
JVHhB2tAsv819OrdWLI5LklF8nFazLnr1xyFrvEyB4aPsNKAH1lD9FhT8MRGi3Kb
bkeEIbPfds2zYxV+Cb+E/eyrYq9ASJhbh2Q+KB704CDu8iWbSmk5yOwyLSONUo/U
r7dCTB2/mqD8K748b6bP/CD1Otuf7J/xL1PkG1ll9GpADAREL+2OtyB55ry204AG
Rr3keTE6xXtl9cPEC3VyKxlHe3e3CchNLq++Apuf13rIIMZRfIxQ2c7EQnDljKbx
aDxhz3L8ealjqF7k96Qtr9bP7PVLLXu5CJEjVKBlshAne/vHJrxlaz1bfEgAYyGA
PKnrbZj+nYeYv72q/8lQDnFfT0A4ipziX6EddKodM+NAsHImfrFS2J/RqTR/TnKW
5ah2eSRvJqPe7DKUOy1u2mXpjqk7CWT1w6eyLJD3YoPg08160iUbg/zIjFpm4g1X
R+W0PAo2qMiHqcJuq0pquEMuwcTOctg5eeUgjGONC1lIreDkL9/ok7XltnTQrBqo
3D4E3S82UOhSqyH0hcOmIQct6Ecgcl1kKpzUm5xjlQnXkv0Nwaatnn+QdTbjWBZ9
/Q5tHJ1TYC+Jr7VBP8AdkNfXuhNuNkrgWUJcETI7c//IhAhdW2hUxh24txszwbuW
xQrD4MIGRLargrtxg8NDdWipWZ099TvFr6qZkmbhFcmyvUQjYkWhXXOEBk0rL4TU
47S2QYw/LYhfSj/VUty9p45ZlUw/Rzpj93/lA/hCMinTy7dVwtUOzPe9ZDHx1on/
xBHu3eruocZEjfcHKNfXGotYETV3vOoQybNXI7b6DbkQfVz/pAGMIy3wVCE8p84N
c7xOZ7OwkMIP9S0t6pgjOgp8fJpk7q7UQ8Nq0oMWDf6d3cohGZwvSq/78eCpx4X4
2hb2+22M30BSbQqGoUH1duNchpe9GIVQ+dyJOUnaESLmushL7YWJuaM/w0kgmury
8xBFO1DzT5TXd+IY3+Oahgwol7P0JyqISEpIQELyTpMTvst0FCQm/l/OABSaHdMo
BftVEOMDkbKXcTLFmYhUv0uRQqEVfwGAYUZW+mtQkflXoGKt4rhifpzDhQS10Bwm
he0xgJcUTH8Kfss3J1usCN1WKTE6QknNlAb61PQcm/QrK0gYem3dTCvhnQ/Pm2JY
shmcZ+8numJrxA7sK7RXacfXDPPzO1IY4LnJGyBFHREPQBGldm1J5slMa0tX6GW1
+IcY7AToD2OkbCxwXqXt8d/s+Q1qfRt6tMxfBvmePwknjRXckvt76SL33F/Smq6u
Jx+r07cT8thJwO9bQz1b1NpGQ6/Uod8hEh5DqWNJ9IX28rWuzKa4aSD2TQwaIupI
FhvSOCobGyUFpr61iHMdYKxcChDpJAz9ysRpTv6zB4a0yJEhkkwLNMc0u9Y6P5d6
/WUI+Z3hAmJ6cs3bI6bexZ/tgi49jUSSRAaLNvetc6zJJSVMhSgAToxyAgrPEubd
HBklm/5XTJP/cLagX7BjSfwu0j/J74FycBvUDloKOL7bxxcfXbOxZ5qLUPX+CqhQ
vk+Bu7cMhPXYduFCxPpafIeuLzSJ660suMhRzmJ1Cj4yqPWFyblhn9SF1S4mUCWC
anp1jdQPIOPz0GnVCPXJ3bzvjacWKk2z7bI2Q5QVnfsgbryzzoPWGtzx5A2V8j4p
usa1TPPLci/yYfbPTG6AGMJqJkIyhGnNw80NLr/iiVEXEP3RWPS2Cyw0iYpgF5zi
noOHHN019TJwWzEosKZz70JLSNZRt441hc1NqpggAfQ7KhpVbGkAyJVjkFRJh5Hk
D/Q7tgdwxM/zCSc93g3QxLjaKT7GJzzr/YRvx54YFvpb5DKssxSvj/fVK69i2WNL
gaBUx5LJAnGMJollj2+6RA6BZ2WpFDFJy5rPNiWWYZyKkGsitC8Lxx9E/s1rm0gM
a3V3fRlKIxCMUUUQW30+RAySh3ztyvjhc+8bk9lropvKxXEjPRk7TU2TMpA5qyre
vngDchyXTyCmQ5Bdn9mOKjXW4AhSSGzjSdgvUWKdVmBoCK2AX7RCdA6X7XCtZa61
Ud/033OEiUtYPiX8fwGdVsibIe+pL43CvMEFXv8w3ZpHl+RydPNEgxxyDX/cvhF/
u6NU330MW5jO6zQueL1il9dHDETw9CXHC5tyVY+PDwDtGX3I6H1p4JdUPyaG7uZ5
KMZDrgYQUpMtz3cGtOL5V7C+kILpUlXH/APejzQ4VzYDodTp3m650horp8mciz7o
/8i3bjxzusjYa+xIS8WV/uuX8JCJEVAgfMV3VbKLrTmaQp38o66HOVU18LcdCZEa
6crsZPGsNCkMqVpr1wYcQZoMYvhbWbF6DsBVybwiXKt2R2K8+F2TLFdFZhZKSycA
H+s/U4PtpatUe3EypL+MqjRsYUsMXNOHe0djoxYnp2TdLRYRSDy0gjNsH01VUS5X
rGo1QO9+pDXIv8zuYsVKveNBLREkzwdc+pEwfabI4akiWK6Ik1Ydq6WYCGLTATWi
zkLhzBVaqkws4ifCrnttBayQDadyCMaKtnRNDi2ooS875rnpeB7RE2loI0FO2iYF
Srn4dMUeKOC9z/TVgisddlaYVaYGt/0I3k/yYRFpsKNSdRDJtc6ByC6Wy/y9D36L
jwXV9oD1YolZBPyklvbwkyky05nsJqzXHkNoCCVOR8F9la75XZpWqp19k73q1pTR
Gdm2t9F+Raiit50Fj+X3MTE2nU0mMfdewsoIorvjmgwvgt/CdRjXjQn6eshEUqhe
a59bkw6cHRbXP7xyI000OGWHLZtYnSVNWKum5sVF99vgC+4hQhY7YVgyrFgFMXli
li+XIqxLrk7+EPv6TpLSHWMV/ZOltsSF88/i2Kd0qOzcmjU3Q4DsaQR2qKdbj3JE
95SPBgwnGJNietm/OattGfLZRgVQjkc4n22br40oY5OzrEPaL1cd1iDIGpDSB1PA
d/bWjIonocLq0K5UeJ8r/FpjcbSyiyZwDwc9kX9IobXNfA4oTF3PjcSbhTfl6pcc
tDjdpKmZUAican9t8ZsmyrGJlA+EbFC2q67AMLOdWrfbQtQcbXelvH7mfAFUAeYt
a7aIhpaawc+7iadT0NSCdiG8zLAkAc+s59GgUjND1/OdwVvSKJ8EcLLzFN+ZeB9e
sij6hNKwNXj9lB6eVLJ9bQh6pem+Vx4BDLX+zFRTF02RFa1mdpyRL5yzV6d7WrCz
6/fUiE5CPk9uKBHIn1xrYIK2Qg6XlIY3SMgMn3eez6yBLH8xwI8J2E8SBE3W3b5C
yEkVqbYpnCv4uvHC5xGY03qRwKnKWmc8sNyFZn7LibcKRBAj+kEB3qeCePLFVlFe
QiljSS4v1l9KGEj2XyYPjXhIeI8NtNW32Fv/Yzuh/0lUTDzJVkl9Gi9hjEvRNTQ3
jlfWlKrfuHCYqaRdodMewGZLSCkXCC4EY3LjX9tW7SWNGB+YBWeLMZ4MoBdBK4b+
nubcX+ehfN06vedSpGrqsYIbOaG8Er0Rvj0eBE8Zx9Bi56dcW5qN9aqc5n2Q8vKJ
H+sdqEA3QjkMJ1L+meM1utfXQKzgMXbRG8sQlaiJ/svNiAXcJpjPRLmcuFk9I89M
MHePT/gYte8AV55pxbePqH9NFzAlnSALFxD37ikbxN3sq7Ez2H1xzY49KKPlln1V
fFB/Wzo7bA+QkVAMSrol1wRs0JVkFyaHqicYD++fyb1x71E03zW/rv4K2ZbxGZBS
wUX2F6oeJcaVungfbNWAnVENeO4exk5HORena7w4GAtpk7Pkx+5U2mbNmdihHAe5
NUWPXGhj8KuDDlCCyt94G394M1j29pVnZziHjhAEJoRYhC/NaduQO136ybQMlgr8
PgIq8gB6TiqG0/o7ik3amB/hyQYtbs6x6KneXMo0z265flCYfJoKYyiXisX+ka23
Ia4aPXXkIZKIa3nted+ybZcjSotlpmVVy7evcBEubClv3zbTvtkZJg6XnivtqJB2
L5L+4j80PE4qwsEZuXUzkUW433Mcysv2JxwRgEtEabJ/95c3CXmI5zZ7aX7ttc4h
tD1qiKafGT6VfcaCG7H6OtiPCCV9RZ8szKd3NgLTx7PXyXvVplR367qR/PToHHce
HH8awabUsxiUL69sZXHrR6LUoSNgnxIQxi4KLtV1CHqEG1dVRTNsi0l1aZWS4+aM
oHJcRAda5zG01/aStMDTaCR5awZvLmKoFg2MUtS6acd20WRh3727/swCWWR1+ALZ
fEPlY2lFOVLrFxNbGUVJ/myYrQ3pbBKuRyQVVqjUin5GJwAAhNylU7m2Fqv29NGx
CbwjdMVj2TcQtMROd/wT8Wy+PLg6bzn5NKi14jCOdkx8u2QPPJtPF0KS0lxdjGp6
1Ndr43n34Rt9X2g/IyLUZAu6gu1qRqQCSBFteZbadlgCILS/V+rtbQel4aPZLl4z
wTGqcOGdivmxVsMj3t3mfybiirCKugONCkysc2CAWU3zYiSG98H5aBoVDKSmWld8
gGjkWJ79Jus3NksPVyfE1fu3ut5IlTshzDC9CUw6zuRdPTOxnTzgt+RLqEGI8zd8
bVE6PosPx36DC3PONs+LqgyP7Uu+JN++nwWE6mx6BnFxF6yVF6kyjKHOJrEA8BKr
HGYDxD5h1OW3I4o0uOp7dVfkxYWjvAHdAPSIwZLAdUDUEjZx3BYbkpS7AVxl+xYC
Tg+P8+enX18kHpKsYFEO7RNVF8zx8WOfPNy0sdMhFmaRzM2rEyFeOUxOTUBsdQFs
79tmY+htc0quNCTmcrt1LshcoTLSiIjTGtDUeW8srWZXXctzPZqjdwL4HnUp850R
ZNnDcp7PN5H4mCRhnR6O8vY67kWyTxjYG+Y+foPGBizTE+V4pa7SU9a3B5tKxCDR
SliORP23craxKddym9AgPQXR15brxfeFMtz3DcmXnKCd7b2CiaD4PwU+OTfZCYm1
nRffwk3OP8Q6Q5Hz2GzC80hwfy0Pgr5FhCMFjOFInF9OlSgXtT9SaMMGqrUUAofL
Iuwrl3Xo1Ol8FMr2s8n6/3dGg3K8rd6c0l3lvUSlHHtvsf/yXggsUz9zAsfSzxnp
+EcaSWzYPzCDNdm/T8J3M++PhbEAMSuxR3LWXja/fbM0QJnpgewfD5kU1JxQYt5a
WjdbwEtMfnpkL+PvzDdnVm4wxVjqXqMXDij+1OlDDHsNo2NXUoM2GuYiqshpqD2C
X5ZVY1S82/hADosxc/v5kHu2pbyFQ2yIok5RBBx2PCE2nfjH3X7i6vc7QOYUxWqP
xD8bpPUkpQ98XnfIQAalYyWhMegZccvCLczRsVaaOR6dVG5E8UTqO8hvLbcqtIxN
C50NhScHWx7jkRpTPOles6N36KO2UNC+e7m30DJrWhTM4/3xWs0GRiCff7ywPDCd
4vNA05m89gDHiDxOt5LjG1oaA/fDcWrWrg3zU1hSyfHMzVjPiyFQ2c3So5ay/eeQ
+OYEZOukH3UrQ+chvYCVGmkTZTSGmrLwDyu4g3L7xZE4Jgd0NvSeEFSY11Z08ObT
QBL7uaojpTRQj2L5TfoEWDF3JCHZp9D8r5bOyl6BIVm3nA/BmeoRr8zqWIemvvSM
23f+asVdVkGwnrPoBv2er/sBzga1zlAi0fHoO3cjl/RX0ps5B1P4EqDZvmT3mPTv
i0hRWkVLlCmxC5+AKcx7ZsEE5t06KgmKsR/7GkUwkm7ZFiOSKUueJsE1V8GywcV3
JouLlr8ozTHQPj73OBOHhHJu9Y2KXSWs0yR5nXVkn/XRcaQyY78KDajZH9AlMqWx
UbRrBKNITHdZjz1cpXoUkuqVCHA7GOieaQ0jhz8p7YP4sZ8y6WbLjlZ9d+O9gicV
odPAeZ1LGi7OWOwmKVcq1IA1iA41H4TYQmWOOYqQ9Xwo7ObfymFs/MQlHmiFM+M0
h331uWcYPTdAn7YLVDYGHeJdicBPDn1DkHzlGk1/6z8Mlo4rskjfozg0OiZqeplD
UrSOx3bpYhIjmhmv42jXPJh9yTobc2qh7RRpKAu/64P4Yz3BSEy2ENYIW2ffFCuc
7t9CoFhSPwUFDeEv0ZxstSsqksULHqhSVW7ka9PUbIr/geq2yMuKoZaTcCai49Xz
ObCjkKayb2cR9z/C1ERXwv/f52ZHBg2VKL1FqkLMOdtT2iKvxoR6eU9MoDsKfPVI
69f4EsI0HrYDrZUljnJhK6gBHkwdHas9kCUXsYatQMFKGYbxBPlPBwOi+y++lkMz
BmRjZnBtt+zW5MfxgwWFhtsVrVuxD+eAcpOqJED57kd/kg3p5RJDZvuqOPRI1IT4
Q5Zsv9K0WEP0nF2d1S2ZMa6vs9jlwzNR16dCnbbQYUh1YLD86UofiW69MWD1bvkD
ouig6jfuPFsbwwyFAHPUsu/UWa4h2QrB7+c2G6DKeUGfi0gGoTn/Q4CsJrs1npPL
IsQIBm7moxVBT1ESPx9E4ILcdOD/WvTyvh0Ci8KYbDHVC/om9E3BEBiuBaBdqmfu
+c6XRRKDK9QoplxQDAvU6urx9b5TwFb+OQS4X0zB9TFivO1w2uU0KuA8ntFDAZd9
BcLmq5L/zhHyqtwFyB+CsrBIoqYY7pat0v5S4sPhs1fbDgKQYwIusRIgEFJudRc6
yjKjED1edEhyqQy52QBktAPn+LRieWOUy0Y+UwQBWhCPOUesuoCWosAfifPVM86P
fmjml/YeSYx4TmaIKITXsNMBN4FFgbGGI0MZE7GpKlW3vRz81o+OzCRFlQWFrFMy
5R4BO51GlCSg+uOB3tOkvz0pkgdlC3wCdJmiWpSNRZ0gL/HFg5/Q9B3cVnEPRotg
OKOBipZHH+9vHfDllwAZnJiHh3gaoxdDTkoltIJAIJKylGNfQqFm6m+mx1y8hVE5
CiH3PdEkLz2dPARPoti9DgctZ5R800rlhqovqW30yEyMm3sG+lcBQ4y/03Da3K74
F3+BgtWFEAwEQ69SzaJa4Zbc4wgmSkyFvi0yIsRueCyamcQ0OenoS+Fjt3/Yx8kl
xzliljlYlljY3x1j5d3fIak0dgP/H/dfqcMR/HTtvFoVvM2jvHMXgU3oKiN0VSDk
sfgb1hJzqPo74Hu6MCpHXfUDSiP1AX5xI6OXCgKmtxEDH40l0PxfjxrCsfXjBpfT
QKNNZwIUGHE0CTkspvrw3Uo3bihCW8IiwM1vSG0ly59UnBfk+ONJEBUgAxkuzWGJ
dlw+pkgCkX6Hoav8FRhTb0GLDaQgWail97Rsmq6+B2019q9o2fQX68Omk6rNCmiP
DNx8gfytxYzqsiHE73D7qdD00BS/Bt2Nr+OTbHZ/rUTAciy2FsIwhFdbb/oNdW+w
DoVTqytBOhl6XEVWO0t2Em3BmfpCC40Vos5J8DGvLvHup1rS2dgCWF2pD+16Lvgd
wxdAeM8GhMvHy54htu1We8we9rdEWGNi3TvAgSaySXqEHxXzH3GWBuT0uzXQaxSJ
djZAFecPUntNdxXtYqLyhJZW9b8l7/wA8VvUwPBMT0ZS58p7UBscgVAhDiBgwBGW
FSgEf6cf/b6XiFz/IxcghCwz7Ch1kG+ra6xzqAHpbOf20z4PS+PQxnPdgSAsMBXi
eoHJJMNZyzgwrIRi6DlUglSXmo4tuixZXkFU/ZbONZ1qyBg0C2cTjPmUixNxjaOj
xAfuMqBiHRq7OdabAtF96+KOXWwJnZgp1BpokrlPOxfh0b/b2Zq2fLJcEQiNN1MW
7z7RnVPKvrZDU/V7i4s8UDW0ZFKYBK3DuwabedvxffI8Y9fymDi1R2ww9bUd+M02
BMH2hx23Fd1Igj07dZPxFcdqrOo+GWKutfPRjnkVqOenO1H90N2QEvn4rqYM7TsO
QzE6+D3UHP5N1CLDQFUDgVEm+QtRrKmhj67avEbg2OdFJeGSWVPFtiGxEzqqdhVq
1b3W297gpBvl5vcQJh9eRR57sQ5uZNf+X1IG3Ft9hVfGq5Keb12SJc9HvBj1fI/k
ZMNEsUye2mbM1NbOw/rwplNOt1jiciod+2gm+DA+X05WpPW3V3eMbEmNprtP69Qg
nEBDwj682q5HOePgKNExrI18auqqXZV3fRlko4ZSJnZGx7Ix0beZJNNoWqaQ2biL
qNBe3CoRGiJpjBgPiQ99oBgLyPalWG23cfey2BXHUSFmn8nK3GjKJlJnUca2I+iz
jpgkqDTOM7Yq2CO+4vAQzSDWTiZDsNDB2e47XF+KWXpJOorjJcw0Hd8N8jl8OU4I
a9/sg/Yt2hAJjAa6kps9jYIggwfKtG9hXwD6xy8YuIU9tSsnelmDLPmBTJsvtTRS
FDyscruNvIYoP6ozzCqGKPrnFJqLG7AYwoUZraJDwBt7WL6qTuTqIFfHVYuM4lJw
zvAISVzMxkfaQFoahhM2skzYZzaW7yOZuq+/C0JqIpeoVy9t0In/zWVav/l3fAtM
xqlXtAszu5J82Gx+z0AOutQx3dkbTTK4taXPBUmmP94/yYaS1o5Y8xzo48mA3HBM
RpMRFGol76xLVAFj4jFeK2bDnmsG1u3sTjLnB9AphW4PAXDTVn8TmuecXonTFG4x
hZu8EOugHBRep0IPxszC2Le1XcPmwHIQYOklIAda0C1AVQ6RK/o6Q0TB0oHqD+Mm
s8BbHpE58SgXTkFnuV4IuGvnBRXHOUyAxnjABZ+JQj+Hn/FgRHoxpvbfwGtecd2W
pCRQZiW5069iVaQyqAjEE7ZN76Szo+dkk45UPRlegEagH9WceDVkBbFlZP9pPgQ3
cQ4of5YZu1FD0vbUHeXEL1bkiLuc9XJaG74QNnKnje+u93V7/uX3YPYwlo22Yamp
vgSrhtf6VQm4JUNcKg67448ItZeaQ4WOL/I38vaoXrVV7NIMs4MUsCnmdvpMExzG
Z88G5QhfodHmHpYT20QwoZNPO1nj6CiTcrlNsar/+aWaPH9SBc9InIlcrfoO+nlA
4abaky1xjFt6wgGbKs5OyMJeAKc9UdfTpZwXX784PPC6uh+B8qy7ab0Rgg3XiBfs
6uRQCfy+wASePkQ4M/BoS8HAVg2VfhJgmxKTCVC8hdgzKMYrQXnTBNTGxYH9IfSP
TelYK1nPjbzM/PGAc7BQ4LTFCpJfCvOBRzXEyLJ8Lb0Qe+h2ZEeb2lmtGB5aLgzg
2Vw315laDg063lrQR6d2vwtDmNcIOetM7g2P+3K0/H3u3iHtCayu/oqAtGNEKS0h
AFvKPL5sdm7TnuV6GCdYA+RTGf0W2UZYOmRRALOVgQ8uhXMumv0KZNn/eL9tgo19
RHhyXtvyQjmSIr1FpLkBj1QWFhodSDAg/xVqvaObzbllunv2RltBnBVpImp8RmCA
sJjywHugnt3fp5rI1uDBKIMq0oYwHTFaQg+jllz++rLi0mfMllp3d3qDHB/6Blz7
u/DQU5nUB6MTyZ8m2kCsCXNx+QtF7IeZLJQ7TblGaCNs6Uhv2cpIzSkkHFSWnxLo
0oYYODokm3GhQBwh7qoZduObjxr/RWYX+LrAtT/VoqsS6Sc2IXsNH62Qbu40bmdp
sRGXzcvaiWazEGIPZPW4PJAwhrdNf5UdcXsMRSCEFRHZXDQUL5QU3+OZhZI00fmr
Zu9NK9BhlphQT3EDGxI9pYWkD8WRzSoeWAnu7mvU2Bg+vI1a8g1Bf39ey4oUMyI6
H9nUxV4O2Mv+woaMTGt8AU76C4TWBD0ySuVW1F8Go+dU6Nuk6Jfe2nS/R4eadSFa
GQpTHerAy+eg9OQMn9CIces30g8jXqbuNe0ZRLa8rpTPZEap/KHVix/rUnQyMh8V
2mW8qRUAXE3XEzieiEpAiegqJgtEr+4lWqfGHLRnCe9NxAXNqQRrPfzwpgitO+cr
SQ4FSz+T5hfZI5HdLm5f/6ITWUgMikV8gyW8i7uCU4H/7cpKos9rbFDXohPaA3rH
sYnFf+ORRUV4b6/HCrjcoAam5+WzRBcDGsr2b7FGVHrwxTok85Llvklf7GiXoAIo
aHDU3913rnGZ80+OoT2KIv1bmalPMKH6R//ubcJUV4BMr0+PJminri1YycMo9ELR
SjaVdx+9cf7tzLIHCCcXQYilc0sqf15jp8WK92PywsW91t2M8TMbYbLG2XVbcCwE
bUniQJH7jDKj217dXYXBg0cSPbZzjx1WJfzeheQc2xdtCRAGfPJwl2B1qVnubF+/
xQjjKIJcEtTntdzKVvYQUKWdW1XMXXM9cZ8T2E3ni/sfu8VOmixd9SUyJyoDr6lS
ZsOSR9uSNd3n2wUgGz+2GFqs58zZGoc/vACq07qirXaDy+ytM8yTH9VP59aZwjy1
Ksg2bc+KSBLKoyc5izwycveaZyCki+hWotPmY/NVWkuxG+0V6u62YwCs02VEwhdE
XJd+OdMgvfSKYy9NmvlXhWgiXIsM/4qX657+PRqM1zYz1tallHY1sENsZII+rHP0
Jj2Oe+/oAmu1wHQvQFUu2cPivk/bHiqXRyq5eNcCkFXa26kCe4Rsw7VCbSg5ilJT
s4Vd0gwYnjzKEv7h14EW1P2OtGnMU2IjZhikCIseiJGpRjH5vcs+Qq4jimmlzepo
skWFCsbH1gVIxKqLC96ixuXfEUBWlTYHflpvDUG0QfD5eotN1O+nRPk9W86YMl8c
uSmCHZVj14wqozcSe7xAA8tCNnf0jyM9gowZpMfl14ZBFwQY/qBECcCM4aPWX9kI
7UPlb/ZOcJXSgRkpe9+AVBFqgW7UjwwLwBgx4rqhmz8bmwOPu3jzIMB77Z4q4ziF
vLK5S9a0vqKvY+/qx2GkHf3lk2kXOFoqc4P/VbLxB/TJj0jckqfbzkad4PlbG+1d
WpKpWNZL2tVZ4MqN3sFnuH46Z5+UCfuSPeTl3dhJxFgkWrtxN7cgRepnov1hvDPX
zyT4tiNl6aJmycQ12dNo8Uk882E0i7SNwfuLiiRw168K6uKILOAAYk+Vyp5lcaRh
inBZjZTyzGwHyV3IyITcluZRMki4kckMZ2/HJZTdau9gSqBc7/d/2fAR+lx8l6FC
tO0wPgzNBR4TieEK2+awrP34V2QrHtTQ8ux1NPi1eCwaeu1Ki7Jf5y1izSR4WR23
IdCSKs2/SxkydhS9Lq3lmo5h9tpPwjZtDsu45Lmdc/NB+aN46FgtvLP6eibyrBLt
2XCa7lHwRyLMOgnPckRFzz45u6UdRoc+UvPZ7bNYq/Ufez1V4AOwgg5vWYwPAKxO
NMzEpHtMF0sTDEguWlJPqJr7ekmNA+l9iag69l7oWWd/j9HQMEJawRN+F4IeN//d
DWsGkvZPL1mWp0v6nthUbOrETYKPqyRVEW74Quh+J8C6Ieqfa4QQNtbU529KGKKK
OZrOTrxGnwyPIGqH12s/J7DlBRYvR4YeA8qbuONIgNamhByJfcvlhrN+RSRvwes6
abXcn6v96MuwihCJ+C2hS6CO4RQQ4pTExtDPegevSZW3CivyvrOO6YCBRaZtg5BC
F21Ylx4yfAE+xtNHeMcukuzdj3gKdy9xNJSF10pTT7428WDYKx8LsmLiGR3AY2F5
QeaxE1OtTNM1VEsWX1lfh3GyoWUSY7695T4BXVHsZRtxdISZ/o4pF4p+DcT/R+54
UOJhi45qYggfYJjX0sQqj0Q9BKyrhhsmBU72QQwgvMdxfKwGf7XoqURBNeMH8Cre
rW1byA40PO4mH4gDvGMQavX/0tMTcf97vJB2DzT7TxsmL5bJ7hg5eTfDp4xnbfwJ
e9DeLp2XpkRqwhu2TUFtU+9QPU7kqbzgG4U8d244Yqami2b36YJM5RbWEd5ATZ23
rG2cd8x93Pk/PqRATuZ7Q/aTFS6Xd6WbqTgdZbOxee4RAD6H49zWa4l44eY90EjV
XbScj9KN8Vg9c+yGhRDeYYeRGLKK7n4azkCyzj2iIwYx63Mj1hmlV6SFw7YDUUOs
PNLJy7UUfMu3fOa9PDDVUN+3VDVbIhqR6D5RxD37F8FmySiUIiR7rX2SnS5PPU8k
KnDo7BR37oPTxK0km30fAoZ7QdrajhdjtNdcOtTFs3nPFMlR0TVhr9nTp7d/U4JK
jNKjgM/sqPueHFRJuzcNZAdXNybJnuQUqKj6bvTEyrpJSBL2XMU3e4uBAdYLldDU
Nub0vEbGqVhzOOg+Y4VOwyfjPMxS8XcOZk6WP1mOl000skH1slSMboEy+EdKkFlM
WLxyC4ix/9UJnnWLhTWQIMF16khNg8Vredek1sJHf9iFhmJQ19YpuLEWo5hLdaMr
MhYGPbrzWSQekPtj+KpdZoEBmYX0azuVyxOSnL7A9EQD68tdSIy15vcYIMhiqoVi
vKg4lcAyWj3czfUQ/xYlX5/Ou60vlZQfTSIg7jm3WmqrcbGrlrpFVu2lRQ2uRxRZ
xm/BJ7YQAolyGlee3qRiAqn9WdyTaLFgEKGgW9toZ5/BRzBa00DJ8Lo0gVTW0MMY
+HBPQW0bYrD4q5nyXvkNclFEjX/oe5brNUfVj1kOh8ukh2SBi1xgH6Z1xtZStinU
Ppy3gsWxtGD0PoZZ0yuND0sgDIbc75Kn2bUfuZwwZuTysl9styGrk4aOE6CcMLq1
VcqxJFsqLiRcdDtkIo6DyoVi3m8o01obGHhbeKpnVangVE1+hq8ASpx2245k7hJ/
mYFZKlehXQ9nRWqmfKYzEijfUAXO8n0kMv13r1smzpgAY10BkXwlBd8jm9d49Z7i
Id5m+VRKyRkru4pAP1gV/J4aN5Zt99qb3rRhg1x7VQGqxHYMsgt+5WnNbcdhVPUo
gCcy/YmgZF5fZxEnU6zXOookmmUHB3yX162VsphbeeT+Qguk7dtgECpbAwtcJP9r
q5vdhSGjgWBQL2kPKIHl322ig6YpXCUX6+VsfzZcTURxtMPFPBqxLiXPs0KPSEi1
Uec2udwHafxvdNIchOVPkz2I3Ewq677kQ71MLVrww1WgIGI0ONN377Oi/k2qv4iN
SVOauATR6C/0C5riCGX9kEoUFaK8xZWzetk7/X0sSWopHjAO/rd+IxsLudjQvVcW
Gy6qIaxuIV9tM0g/p/O7sJjtsA/770hLP/Ug9lmAnLbYTVfFXDqSMUA6TNXgPoxw
OGDBcLkZ3CCsBqh54VxItgyV1dAM4WsqQghTAp37iowappbssBPTRQoJQH+Vbrkb
17I1fWNAcJ3zs4Y7yjqZAnyg4M+JIp+IqtvPmDwi3OFPSHORV2NTIQ35o0XmBQBW
2X/yV7LV/GblfJOfnza23AewJT9g3l+rBwhyC+dnjpNQOEZ8tZ+teKXo0jz+hIYD
bEAl+kN87a0denglY2CVNPKXPocrh79CXLMobPdS9i9FnmGuGWc1jwBJjFEyHUVM
/mOKHJQeWe/G+yT7zVGm8wAHi3df+kOXDz1yMIHGxKN0/kVpWD7XCI8LJNKjVPGm
iQB1z7XibeuDjgfeybVlEpMAkP66xlnR+P1gxEOyVE2Erxbiw8OifbXkQgu3H4bo
WFlEGNiL5+7nf9Z5Afb4jh9b3KQNmZMIQ1FxVC3gFsgE2kz7ejawZpkI/Bb/4v2W
f3ZP9VsMFc0mILPdOnVt2R5SHS+d2qZqlZ3exl1VQRZzhHR+Xgwc5Kzq7vVILUha
HAE244ctd8ROi/IUFTpwlF5JEEDMEHB4hAX7LMXblBxPX3xq47+EGMgV59V5H6Iu
tQRWio/tnHeqENr8Jl41mNcHg5Xe263ScFOIzm891UNEQU6yFJDAa146k1rW/YUv
TK0dz1mXrxGHtnnR8jfikOZ8Ov2XumbVRYSAJo/onJUY2jjrEGYp11PwH2PZqbFr
Ci7YQKmx2U2gx0qF2G/YiG6j0pKQGH1ieTdo7+NnRM0CRtkwb+taun0u89vT19/N
+xlz4bjRBXMftA6QKAOostRr7CFdpBe1nScmkA05L6ST1M0ByWfhFdVlnzJ969lY
qYKJRJAGB/f0rBmXsh38ZSdPSNPdLqX07Z/PQVjhy29K+b5nhC4PVci8Th1s1eWz
oGGS5qPwsJxXhG02psZj66C5Bo8B6kApS3DJRFfjWSwrCLVJOpfPwNJpgMc327qM
zvicN0+XFEOFfZf3cq8Jqg7zbb6egFbci3XSTfwCEKemP2wQ8ejk8uDtpJ6SSNg1
I4DuirA0yMDKHSdEqIx+yEB7KYgAmirUWHwvTVLKsSzv9jXYnuWAQfIaiqX8IdMi
BhGv1gDajhpfbMxxMy7wkUC3A+cP0EeAQvMBSYm8kQl83FiN70Yw7dRzDt2q8KTC
aGqmY0e66ADFYNLcV7KLBq1TXP3Mc97naxOhTu27nFGkzoEZg5ZmH8tNY50MgMfK
4iIvIddDrzY8n3r0Yx4mOJhneGxtFGz2SxkvnZsRiBQVvIOKK/D2OFlFb3rtLBoF
TA75m0gpSrDPSVjT0i7G2RTsdb6AmOvNLUjDSKfi8HIQ1KZaYviHRxi2N/cCziaf
ornX/3KZ6LT7VnbWwb8KxihYeH8LxYumJA+xskwd2SUvlYh99uhidJGM80+44fgC
d/al1Ff/gnY8uLIusYpq++ZbtTtzfjabz21R+ECsd55SRsgMEqaHZkhOeBtVQNrC
C88WXxgtpalA79Zb6eIFv0qB2Nti4eCQj7kf6CcTujvrn+0LBPuerOJ0xlHs/7HL
UAiAiGqHdQM/IHWn8mgBEnxDUFckVCdhOTXlsEu9iPIVoW4uaDzqkgN9+nPsNXcW
5MzcoSq1yOfO2SKUIkZqRRpfzlfqdH9q8c3I+ESQuLetYMKJp3y1tNf/LTjJ3Z5W
MWKO59+bkI6YtWHxO40tWiIzsx1Xynk0nLkOFFu1VADhRxpGXDbhEG5iKfRFOQd5
nj5NBwHiwrE0ms48n75abStGCcfr6ttfI+u9DFtipJq2Sfwe5mT0qXQLTL+ZYAmh
fuA3YeyHoZaMt98+z0dw5yEztnt1yNB5YuQgQbiAWPnpOy7MX+F4wUfL0hefUgbI
4Wt098LP27IwGpkO2GNxYFi0hI8IXJ5Go6/ln5YjBDc+/fCqrOFSHTV28WIhM25j
ufHnpTMRuGs00asttUuxNQUBComO75fbEAjlkBHb4NINBvrRB54Ko8UDI3dCIkC5
OiqHk5Sc5XXBaELI6qnqzdUsxEcBq62sV5iJfhRKNXRqSN1cQ5j8qejS7/UpL3Bo
NUQkfd7vrKaM+byGWk8LuQXOxgMnK4mwckwa+liizXElJwTBcQUf64T0SFrWot4I
FclUsc8qVpsemJbuuQh13pqS9ba08RBALj6LshVM9EkS0lrzLlLCR1ZXYmOIi45b
LK8j1XmI3O4Ufs2kpXMSfbuWVX0BhBojmuKdI7/j+vfqQP+2AVOxMb/qAlUjHjdz
zNanKQs49Iq4ABYGFMSDC3vvus9nvgck/NPqXD6NFNyVQRzLj17GDICyp3cOzO8L
B9VnmOqXTSDAq+7S+exslPjYDEZg4lcRCFuSrbINljF47ug7kFZ7VBYTtSqB8M+r
d6/tSvHoOmHPfOod15gsSH+C1XtSFfgGVsQrzpN+aHzgudXTcRgrShkPu9ccY4md
KqnzBOqgoUauMaFYTqrK+L95J8S/mdXX1FMlnrfvHcHeHtVqblI1SIAJ3e4+t9LY
u1IJV0mdr50Vw084aLLDO2oJTxLbDL6nM4LKz8N6q2I5qD8xP/Tda6XguicGIv7C
kiJ0zrXCWaUR2E3RNKBT9LT1vD0f0l7MjxBryP56kz9aoiAQXnQQMPOSUrjuIG4G
p/ktLfAxKR+zeMvVpA4jNLlDJbWZuLBknI32WCtfpRsgVnJnW0G3SOfBVELFW5s7
Q+1Wo3JaQoaorFSpFeq0H+QoLtxI7aqbHWIT6eVzdpwNc3QuI9v0GU/f9lw7MTVe
OhT5OPGgs9gGU5KegCxTeVRSsw2eZdgdTb/RrVd8iDkRNnLgxRJx10UxGP6RPJss
RuGOhJKhPZVr+mG8lxpeRRFJUALcLOAqSb8UhY9/Qg//bLgQXw73TdsmK2K1CrBZ
4RM5WO0K56+a5KZ1NipZWIUq8Tg7+9G6puAgMnKmW39fXq4qFYNl1mM3l6HoR3ij
+uDLRstPgLvWCZWBs0XG4wJMCEzNBJLD2vZHucboDHfcvk71m0xAcvZOPSanNvh8
rDmCQsFeT4uxmtuR1Q34eH0pL0U4smxd4CjU/BuVS+MqwVZ3su2GkqpbqpKHypEs
aE3FE1zlD1l7/uZH5IbRW918WPL4RyH7p3RagSQrkDcu91NvEd5+Ew56prcjnSW8
Sg1Iyv7FTHaW1EZ9bc5AX9aToA0ToOLCeVdwTPFyirgWGEmimv8xV5QcSE7eKNoH
2UM5pjYl66bcjvFCxvQhTwyGtosYo85tUapLKjWe/CBZPYS+I/Hi9rZoQFQSw35D
gHJS1zfpW51h7gkJdBQ+PSkssmYVkp6SZFiy7YyEtoGLFa7eXkk7nlcFJZfkA5zF
A17oqgNZ6fAGVbGTief83b7EHwliDbqjtvLef2pYyIyEs/YyhVgI4Ya4i12NBV6p
ODBi64ZZquzLVShyg9MoLw0McixJ7fRyGrKqkOMfhtFmawD4ytRfT0CIuAluCx5Z
tr2iZTyJbgCMXlxkWhYwwOzP5l6Y76XdDk76SwcAqcmsVXA6zGcIvcsr6IGvDHzQ
hvxrlgOEypc6a+2MMhwAHrYYcukFLZiNV1+LP4EFEaVF1UxObWxLxuos4PH2DsFw
VtcpVSMsEEb7XUFo7+crsalZvdb9+89q4euDLbwUAfVfTN7RR7UJMdGZYnUvfec0
5YjYDR4SKbcrouOUf/bXnrBYsB1MBCcVlgSDPtihvXFz2DQNX5RyQmF+V+G0r2XB
DeS184YV40PXjVybTY0kU1PWNgNc+XbzrsiJlGiHmpE+w3EYaJSo1SbdsCeJews1
zpUX5C6sbDJd0MO8PihOHMvrZBqaeetKHv3Dr4v3VWXE66FAJ3SWncqg7t+9dDDY
1STqJuyN6eD6Oe9tkMOhZWmClgXT+t2EZIkvQDFU34kOCfYpao7UlHrmv+fly77G
wpiiPAWm+DNDPjrboXyOxIBW9vSiGDzK4445fE9TAcn/XbOp9QE8Ms1MbfuqWuFg
cUE6NZ1SLXf2D4Q8yHYiD3BVhM0Zh5iH06fL48XnNkaqeCgY2QWhkUozM1UOxYWd
BBVQzeK10TlsyAmbLxCJiJGeDc3BMlA3Xn6zuewvaRjW73L0hXlHB1n12S4DQ4Gu
fBFWbrODNqJl5B5FX9VwDrgYvJYuEz6ff5IJ896YeFNjrC2sBKh4/Ifdy5OcyU8K
YumSs9QTw7JZn/lLcve2z5cEFTSnfNthG3hP2/vkLYIc5CdXLLTYSxflVQngQC1C
alk3MR5YubFiQhMLj4qe/4PH4KBy/qHu5Fc+qZsZ+Jrz6n7CScI0y/gFLsOYOZtt
5jcsWwnawAKO4oz1mxZgMxJViMTDMN30Q8JyUi0vALf3ePe/4uPIadBesVPbKz1+
CnCt8B85GRpViV/kp05SxGTvGEjZIwXVKu60jpstcBVCsxTE6s8rQNNF1+7Twjhl
kbzB5uWRZXjZSCJo4bPa3kqervn+EmR4xUBVHPKR5g9F7pVcoiqP/2f6h6GfABzN
jRXkDfm6hbM6/eNrD/gAy1n7cjCURdF9pBC6CQ0IjQEjXz0HVUSJemt0sBC9ddo+
4xOyW0QnbJUtAQu5zsFZr9szyZcICAv7ymw5F4e9M21oq4DVT4iT+Pn+TLlS0CgS
PGShrsqAxEx5ou4YoA7Wzn+TNaniQ1EOoaYBn3a8L68pyAJkp70dpRUm27W46gY7
CMAShD9f+dMNsxKijebhwqtpGxLICIGstVI3dmK4vP4yNSj8Itifny106jRLrXwo
28J7Gmq+ZMGoBmztP99Bkc/1NAKbAg9Tepjz5rrL6Ip6PqX6hBxmKZ9unAr9YNJW
C3fZuJuaoAQ6V+m65U34xyGj1Iwr69lC9DCp7QA1PEm4uTxCPG7krTEW9Gas6nqm
ODOTOHsp63gMfUw/qK88T66DFhS2+EAn8Pz3nghhhgLMgMq5GjYdRnxIHTevEN+0
PWMOBblXYxRO7qypfbFuD1d1Thla1/uLl5RZo7ruVETpKMYFn18eyBhB/R9at22e
YpSFZlr2Zht/CpEEhb7WK0+Eac3xCOluhGc15g5I0MnwLCdJ366syGpp9OUpFepF
K46MNRWGcW6K6AJfsGqDFuJUxHBfFm1OiRXJhiXM99GAs+vYjMTrx9cL7bt7/yoE
CFyAoS72DG6XWpnPYGkYXIDLkbB4RNtHlyrh6yI6uFMe+MpXYPfskXykwustOGQx
0/YDzZR9NIrmujDIex/G9ujuAzr/bnLGxeTWR4L+n1YHUDxbWZtAa1hXmwag3KFb
3mdN1ORl0PBAxeyV/ezgbVEQyEGPnt53Y0ow6UJz5niDTUN89+i/SzUcJxiO+tcU
Ih7VaQ5cEXCmozlUJJbRn0Q+RAQS7TloHGxhlWfS2Fz9mm8ZUDv17i/X01cTs3ft
Zyj9//m/NJIF6Y0gzj8qfamMhOvSLILoY1P1yEL/YC5go0m5vTN1gkWIivdW2srk
Cxm9abd9Th27I6SQC49tLaVyG/RP+gmZxnBIE9CwyLUdSCzqDk6zbDedD7BkxrlX
B4ra9wXnyRES3BKbdlTWKxe8PjU4dLGkQcg5tzIpswP2w6AHdKgUQQbwWuPdO39s
L3dN+TGs+/OS41Ryl11JsZkvuvbky5LzzUozDKNs084odyKXRYL+jV/6HmeE3Qlx
8bgT+eGoai5K6cwmjRLAM1PD0sp/ypUImeZe7M4hg3s2lp7YEBXY+yNK+zTzmaKW
iTb/IKOhqRZ0r3XkaFfDTQctDJzzKgjRmOrjju5VlgB0GXshOYHonGdka5pnVtqR
5dIeOOPgUAkPYxo9wY2gE1OS6jc9aGg/GIYL29hjxu44FHJZYS2qVbH4vZUGlpXU
MOjW5tvX7PiKmv95LgEYefMpSZd7zcXZAq72y1VoDPVX3TR/gkgUyMLfFx7Y8Hwt
XIj8PKSBP3s23D1G3cMunWfV+42iAJyKixYWY5eayGmMlNEfq7NM7wwD7hjijHA4
sP6aLm2wL2uxhsGaTZLBsODMZQ27Ugzjkbyto/6Rke6U0tijTmAmCR/SycvBVyrs
Bu/0LCOJqw1hvzRyf5ni/IPJ3nE83zivXQacfMz8fE5oVH2/TCMyNClDNhfkriJf
pwtuZa0Rn06FpYC9bL8+I2wabLKt9WZdHPyT7zuE7bYNNgssW+fD2Ht7D0VmRF2P
YGes6CBJgYArNv01zvrF4C3k6ZlfSxYaessqoNrF6gG1pda3tzuCUF8Rg4/W0aqi
ubascwnmFHMkuA75TLKfbHWtdOiRPfU/YAwBMQvJE9WNg0kTMUgIb+aog9p2EWmP
u59QYu39keo2bRB//NlYbmtdPjCYZxFKbj1NzHAOgyldaHZUY4+Va4U+kruoE1Jj
F4fYfZyHYmEiXXfLn9eIvPbM0CyI2rS7W8xCqWSrJNzPkKAoZtBFeiLC12rsHkZk
5t2aFzQpVen8Qn2paIVAjTRKPqkT4xSwMMijcCRnL01uBaC5U+LLk/iyOXXYY6pp
HumGJc+Mwd2jq2Sdr9jcNpiXmZ/Jr8dat+NwZdLjAADwspnr8fILThDvZXXGWDgY
TcrTo58y4n5o7n3xAV3Hmtg4ymo8eewUHWTueOEj9pfsLWVsrYpLh7C5KGB59s+f
4mOnwsoYSdnrV63qSgYW8yvIw+kZkbQGKtoG6eFF0xfKHYWF0fu7YRTTnbdDl7fr
2HMiIXdTATm/MRuYmh3vw2w8Qml+VydkoM8Mf8BgyPYdus/WG6x/sLn++QLC9y3i
aJOBkfQUFrfp2aXEXuukQgxr8bsQ8b9DVf7zq5T0ApsKNgjdifkUxJyQaxf2Q+Ld
KfwiGSywxI3xuVHMC9FSFloi6GToMRW+Qe6nXtg4/s5qAQzSbr+BfyMUpIGVfhfO
sHSc+60JkUqpQ4vjyuUOSkPjxFg6MlGscX97y2o3sZVwQVVJe0pZCraGKrc0lEiv
trNA4uVDEwbgeLSJELM4UT4ayR98QveiMJw5+YeW8/Rv/yInF9Nc4ntp4tZQZ5r+
/tFqDkcgOkCTm40oPnOHi0+PThB7eRENKxgXURt9fYjo/NPSfosxpFtVK6RrQv32
p0G45FwRHZbO0STZfS+a+m/NeI4w2EslKQ7RqBEfHpwuoJIZE7y8RgocIyryQsll
r5YmeeeQAHxuuC/6WgmfKOW7cWi0NpnBfl0inHGXJ3RJEM3eOiyYbWzHBFJ3q7U4
7me32D3R2d9up95zl3u71PdNuVG1d0zm2p7ccxp88KZKLTF67a0EmM6Gl3TpOv1u
+9Vnv0tsnI0Xho61Ym7D/aXqmIkfoRMVpMX6dshbQpNGyzzasMR4cKCAepC8Nl+C
4al+ZupZkB69PkPhU3fEz9jiZxpmFk30JqMF5GZyGCjGIvUiMvN5VgTxpMrEEQzi
V7GqmTKOdow9uz/CL25JLtVGpua4d6MO42ZM5HsYZ+QWkr65DHwNEIe4sYZVVrry
wqvGNvULDa8xPsZoGxUixKPSt0laCe0q4Z7Swda1P7MCDJZpTUFPNahfwHYrLgjv
1ZG/YCeoioHAaEo9wncDFncrfRsq0C+Q/1IBBjEWEdI7jjDpHkz+nSv8mebvLe+z
kZXfti9K/OjtP96emmZqzrwYIpbQPkKTOTl70n6W4QOwSRGs6+5NYluB1Yd2PCV/
h+txnYUCTIm9WOwC7dADhXOu/DlmcXFo4ZmG9AMCGlXWYF1U6viPR34i+vPTFnAq
/FiMgu31Lm1YOwR4FaStYuVKdGUUzYa61LX1lHGUqsUjFRaEcu133MY5jZU/vEnB
XB9WUBtjZxKqHGmhGmYEbMZXo+Ewy7FSV/7Oq2zTykBFAEukUJWT7UUKVOU2PTSl
EXH897ICnG1X+nyKUpddqqr+ZQKQfFfHwddUjOC0HGV2ibQcNqGRNfricYh07eo5
i3NtdQpkGJNnhJeB3GF3ZpG/wPtggpcH0K6IOph3QTHUtdhQ/IcNp5HA66F6VBYp
gVKwcLXtWJo+YU3UMWIbJl3DohDQFp8kqpYyYV5LqZb9jEFEASqa1dWSnpwTUwOt
r2nf7zV0oIYdBhMptuwgv8mCd0yJk+ox2gSgR8a38wHAXSWCiiD16BO9V69AuQp4
KvMHAaxkJ8mPff04rnxS0DgFRLMK8qQF4Goc+kvafnVS2akv5MoeOnXm1tGP49a2
R1gJULFxzXUpENoZzQ/7bD1q1Tt6JQtdYQpCa2tRuw8IXlam0NYtittdU3NwURGu
EcnPUketOTsLZPVbevQyoiaxMaV5ftKMHI+Io90axeXOXjO//Md7rdkE49DUzorF
FQcxM+OkWJzDwrnelHQM8Eiq5nBEVf+jCKfFU9ZkEAEJa10g7b0T+xhizcPW6pgq
kdqmdRlVlrknbPDo/s+OInpP3PLcBHMd9oBAmXIn+RZ+sRN3RD50N1ngOEIBfcHj
jjXAQfoWNlt1mN3sDLAnO2UdozscPP5TH9WRHzF653V/qBM5qBtIAwbP1gj64Nxc
8mDCvggdjuPr8zFeAXd14RS6futmALrevuhz1adJX/7zIxBOZ0Afq0gy+tmGgZgK
qc82eDMDrQjmrh8512YAJHAcdoknpLWcXdQkyldHzCkJ9wWglMos1ykNkOjitSp6
sjN/U7UdRaQhp+EJkwVi0PDfPh4PpkrGjq/mjNHfG9Ml1x0E/QcmoiSLocbuf+EA
M/9k1zb2rnQ2zefffSJgBNwWIOeY3TxmiCQs6UUImTaaL5PhNfrCTU967kgxhyZL
8kcN+TxrHhqGhV4H/4TJ/2ukUw21kmnvyNcWAYeryXwNT39kR1yOlgyNFyeMFi/X
1sgElCbdzTxxI1IWhphhJqvdPVj7EVgDrHsi+4Z6S/1dRSFHY9a7U/kO1jsC3vf+
hHwxuRUjsxcp25qO1L3yTaEvI7KtJ6Fyv/YgaCHlahphYzDHR62pS/65cjejbs2p
B8llGUvc9MHCYEOG23M1mFPjvVVHuY9PHAUGML7aiQPdvEPuNbH5qkxs2V2mlVH4
WBBJ68maNKGc2UpPsZVPh2NGvXsnIuuHJkHnClNnaV6sMuAsrnKKlG0An4tJtP8x
LSwHydlornva3rxSFHujb/07M3IjZM02T0Jl/Wj1fW2uhejnI0XPBP8pBzQzuuAi
d7d976ZkIFiCFNNPAgszHmkGIfxUw20t6ZMKfXKq7VMkGoMdUEqb0rrg60ooxtMP
hOkTviLiWsq2K80LErlzmdg99kLkNLejFqVvgOZo/5PamTtendycKnnTZO4BKQnn
/f0SdH92qGx3cbIei+9DoHr4Z+SSvgnN/Tf0hX0Pja3zyN6jEz6TxXElSjmg5J9m
DRembAUEvbMyOFNesZ66073StdTAs9VGm2hi2abcNAnF4cPVCVp24OSHwrtTw7jU
YhBbCnXdznKvJt3XU7HdN2zyWO2gsjs1h3yJk+J+vosSlCC4FMSBu4vW39qJKYw7
dlYnBAbKYuxg/3NpVjs0U1ctqIRMt/XrD3go3fjIGJR/YRTJqk9YmhjvBkg009TE
CEwho5QXss2vUeJJNMVUnc68wRJ0zwSx5C7CeEaZLtF/4FXRswpRjUy+w2cdSv25
Qp3CTLAWLtWw85s8mrKj33Qdtvyo50u22TSBTjVgMDuudBuOH2bHlIEPyq5PRuWj
+RqDeH6tEgyjtq8ddqv2QpiSvqyRCnkUnoDCYoKK0TmYemy7vctR9Fkwbe/q/K2c
1VQejf/+obp67UfUY9V5TTOrIxYBpbSga4/FaHN99gQ2Epqd5p93RUbMJq1XwxRo
AyZqGKTN5ABbIYAnyalgzJ6dKZGCAJWSZ5S99RE2y1ZPAkVVBWIqZpjnan71x4rS
udfogrMSERbVPqS8gEkg/w3jgOLiqfJfe1CFtNj2OLWqr+e5Lux8RZyUmiAk0/xe
2nJn98Wszeojhux2g0SryF5B2LuDDITMmA75yeK5Cvx3imJnrYXbd2v5BOXO9ja9
50QwsEPX8cemWtx8ROP4x99xo+unIJ4g3Tq1RmVdBrvyhlLbpWxoOEM0EGm14BEW
ugLFZi6AGB3U5KavKoVc5eCpdcNe52ssMNfk2eeBYxSkEQI38DM926Zri9ibD7SZ
rkh0IJEVrblxflqDC9AJQcZSaSreG6OvbOFmguQwjnyPE6K79aY0nQr8j7/D3CxY
Gb5IQ3X55Rg5EBBdrWZxY0eXF258AY6Q9dsUafxrznRifqvLvLeb8KhWU+gHY8OL
GkvcUCYITwKklRYQPW/ZO42w7xMktrKDK3t0yXwz45WDXgxjRtRsGKw/uibBp3Ic
iykBhN0doPU7i7RSt0fvhBurBzzbiNuyKpYy1K5SkcUhZZ1zL0DldN971YdrbU7O
rMnpxt0c1Tg0bW/kMksdYIEmTTqmCX5qFzzZdZ4+y4HXfV8c/gqJDJWjmdBZ5Qro
IczA0TflWlF+zFrDah5OwqQSgbCt8+i02KWkQKAgCbY7lV3JJJe/hVBGDuqUCMmy
V+m49Nf1+7r1k0xjyU5CEacIRZEU+v+tdLAotI2wNyseEdLBj835F3KW0npcrcek
CAc93VMLXBnzScz2hrVbElOprfF+WLlnGkow31ymAZmicDBl/t3s0gFTs/8Wmzgm
FFk9t4oNrGbXZqFFJ6n685b4uskmOIMz1GfyII7wuqfY/LR0ADZbBNLu9KGn8kBD
ZVLQsIaiCLsRRONACUN3+qP+rl2Ubpq+HhQtJhQdu0lJjSko542rw/4Z0/PwNe5p
Y/joguGsZqlQpN/dYtu4YFwJICnO+OfrO90AumUSQqyVM460hX1cML3p2isD+uzo
ZxfV/mL9GcBDQN63om0jz45MIZ9aMK0MD3JqwYa02wmMyr0ORXawlG+GvkidH1Sf
UIz28xGoNBLWf+/AaidjavFqbiEkEUyAo7ZuPd5DnO2hFp+y24Mx07laX+nSwKTC
mJlpSrx9fEV3/a5MVYf9CoNlLJZTGVpak4R1v3WMyfBNseetPINaZaG685s1gq9k
t+R2Nwe7QggZsz58RinE/+YZ7P/Nirf23n2LLaJ83bvhSzmJx8/3JneFRHjaYPLL
l2ru5jTRKg3BpmwAbbixXi2poRfRJT3pLZshjrKst/3hd3aSKttfU0wk1vwVYvEI
s89swqmU0eh1ypxHtP9ZhAZguI4EAiDSqFizFL+s1PHEK587vqqQZZPblCwH3S+T
bnmAnFMkPhmazwyfI3MVYCv0/DKM1aZ20iptN+JgLkRXGALhlisXFGybrQLDdar5
UUz4r504KQCxA7epHpI7XOfKkgM7RbUis85co/lR3NjaOXFfHuy7/j52SaR3Nih6
fgagluk23WdGY5VPV5Wl+ZhzUgSrLfnJhD0meYQaPrvoc+p14LCdz+Sthp2CZ3GN
aUbw25lkFpCJ2CSu2qkjLFMAiFPeMDqq/MLapVQxVfP+O3+jQ+qpkTTDlmoiO84b
iNdcZfZIHeSt5QS4YtEnAJNkV0TP12jnZaAPf+N6C+LYBTNU6Gfx1Aq7gIjNilAY
nWVPb9xFalveljpcUrGi5B+ma1YHt5PvFq4PnaEBQJwDmzI0Cs3iE4IDW3MZU/Zv
OVQtt5/I14xBZiORnId35RUSFhUWj2+KXSF3G4y9EbpaZ+MkSOZQUE7CKaZ1nhKb
qVpcV5UIXeMS4l9AELgfkyWjuQH9PzVjRSmINXXho41Hv+xwu/59r5dzoIl8ALtw
u2pBqKhiOPN7BKg4vORAKSZdxsMH4BN+ieYFwmocIspyQFBLmW6rLil3dDZwq+Dl
Y7BZw3UtmnYYEHRsNEqZLF0xqd9zYnWIvztiy/B7fBXmjp90jejWrC/jahcDpj36
2xfjVifz2oZTDMG05Yx9Wj6lPtic3SeH4pydw8CuueDTLUG7+1hlOZdkN5KRFtXC
wUJ4HXh6T+wYru89AYdc/vjoqSxSETqZ1er+ayXWHxOiYvbUtAkkc92aQyKY7fRo
X5kCtWvk9TrLD59NZldW0VKBQL23sRicZcwW6C8QYg4wU29erqfqf12cmp9eNeFk
BPwcdLh9x63jmBCgixZOl4pTEDKl+jU4HzAcMa1/uQov9fLeymMoNy942Wwfqgcx
kaKQaSAQ1jw4f2kme4k3PFB+TOQQ1IYisNXu7wVcR5Htz9rZL7TCdyUsN0L0cPoo
NpT5EHFRN2FUouQJW4/S8uuJjxV102wZM0pojKrVOfSkta07e7dcfNIbVvNfcAfZ
sA/mypSvBnJyJOX4LjnBeF1fe31EcuEHQEtoctb4N4gd1jyDlfcrYtrh/b8hF0Pb
j6MKQzfrvBoVi66scAH9S1jy++rkDnxeKeFRdHRIs331DMLhQqvYJLrB+0QQYkl5
OVhtKm7viP0HBZxpmhWaWCpLlfkhs0hyKCaaijxrWIuQC80kJOiP6gex7TYwvjwc
Bo8NU0McaEJNDTDr8LyEvbI42FQKYI6daP4GKYGIWEqs/NScKNKG6zYPWWe3xrx8
WifG1fXJ2N1GxKezB2GYqJTvatj3kYezARqWv9bq1Ws83rYGQ2Cm5333t2br37Yq
7XmTVFGoJffwP0DXnaiWJosu0lzjk3CpOJkQubSiWWU8dbSZNPxrj77ia+hPZegv
DUY1q0TCkfNVjxcEDGMzrDGqOcyJYHFGYXjTtefCDoYAjf6i5rC24Ngcr2pT3jZT
uGrt6Ie6o0VhnZjBcNkxO5pyaAD6etKMSiX/7n5rUkzZUEATjLG3bJe9gosFRmOL
P3b/ku1+VOIv42uxcjA1Msa37NOaS7Ko/bd8R4FF0Wq9KT3YgLvFbe8VvOAOHm9a
xOIeiybL9iF5bWGoFBNKJez1/+vqdpWu2x2BdANgxEnBYaAMA52vU9COMLeQJPp0
540OmqBkWITurr+1YHVLJw2v8h5A2NubvjUo6t0CdFmSxAMEdtfrbtolsMYgxsXd
XbqOdok791pY38JY94o8/SEdJ0XcE0e73XaVaGDiQ3Iuntqvw8sg83QPfHu1a18c
fhcK+DHFhq8JNPC4i2/oVupekqoMmbnURAy57DgNOr/qYEVMtkZPEwlrWNq7+8lk
IRtoZoO0X4jh4KqCg1ORK7P4fztluLdIZZfL0NeH6BRWt8ksVSIQwaV26n47VL1Y
NlpCQSyJVIHaybew8ZbYJFq7C/FGet+Ni56n0OtTf7YOEDIQFRzGbVyBmOfrd/N0
wI5gxkqFlGQw4OrXcKb200tfIHNyFURdvs17/DMPRY4RpSpK8g9rv7LnGyQU+qkN
QobgH87RwbmgFeAWSzkjAOxJ7RHma79R/IgjV8pjVpcvWf5kRlRS9kqB9uT+3hfw
0TAGL6YDURknrJ30NcUt263jBot8mM4WebaKVFVBGe3cUAwd9e41m4WEcWM6StrS
3uW0cYiJzxOUr7vUQEsCRHwekieyp237AdL/zy6C91u8S2B2S4j+L9hOifTfBNB9
CYT9YhmPQexEhgCAKZuoQRCRjOqCiltuozFsneKpkIhwbK9vY/ECnUw+xQoVUsBY
lobDxkqCS4hBb0PpMcQ7OhikNy80jlh7THXy3PoAb8yFAJIU0Z598APH68pbVdQI
d3PEYYPteoZLMHGrYBNNcRKhHHVQiEfZx6rBaJmyf8sr7rt3S+5IzaPftd8iQkGb
nP5B59e2wSm4o/do5iXw7FXYecjvaDcNFBkBmUkhw2GonhOWR6rri6QxEgbPevdS
TWAlhLR5Z1rtGXT+6LQsADYI0WBGk5ZJ2amKebK2gFALGey73fGx/69iap3tqHgs
ezndApuP+RSlmXW/TPVF9WZd202OeAsbUbMzs9jiF1Rw1hopdV4g/5aTDDkoJyu8
Y70AEc4uDdQNSexzh4wK7s/Gd7EObpHZk2L0l9jaleyI556FO/K7ZWlSzcsXfJI5
1KUpf4yqGTFxTfmrAnziY8/yZJ7wjy53K22uB+BbdhhtsKXzUzr5TIXS4Nb/hPLm
4/tln3p6FhvzvqdNmpxmE+7a3YDi33Z3qW6afXLpuUbmvWyuc/1pcWWXY+gtM0Fr
6ieNmFZ0DwurutL1R2CCGKceRUP6uJOEwUqsd7AiMEay1xxDFKdf4KUeJxuIF8/r
5/V1fXIvbWukiQAH/38F3KgLri948EbDpobVkBJknj6Vd1+4l0TllH2PkE+Y/js6
5e8ZvlJxVdp68ldhxva+BEnvLfaRbEGQEfQJvVcUTXyskM0uXOJWs0jxENkLXBzI
52tsvagqHrpkOvGhaRFfu5MuWyrwU5d60czYo4HX3ricWTgQagDDx0kxzjNLsTEo
0Du1zabrT0MXQcOq2XAvKGXhcRms+E1PDIwwON2d+++sE3tQmVtLz6WvWz1J6F3o
0xfRdmQZavCam0UWoMajVhdAEOFWTvh1dSN2kfJI737t3uim2mYzmcUj/ErglmA6
azUF6/Fj/+uiogDNiCYbaSprrT5ulPC3VIA6s8px2f9VDZzaP1Fuxia6lRQ7Iuuq
RcGKTIF3o2oKA3+cw1WhP8Fc534NtwNn5Pb4oRhoWNeQiK5vWE6KRkR/JR+D/zw9
r1hpxAwDSj9MpBju1i3nHx8wQNIFIByTCIbnQFxXviwE/Xzcc+1x9R/anhhw7ShO
WEmMl41BMnREK54fsy70AZLuV0WuM2FeFNoDSPB3aTO9KEXZAzMatwdqZhSMnwwe
WLi75PAwWgm1facsLu48cDD607VlAckMferc/3g52XtQENPHpdIrnPvPrlBrxaOn
qvBal8jZVFoaUhM6o+xLtMnR/iprCpfn1CML+3B0DpQXJ049/TtxR3t4SJHN09gu
Z540+JlOONuk3E2Bsys7VRXUiJGkC8e4sz+4UvjkEB8cIEZcZp6PsxUEsyvjszA2
6b2BucnsFQ2HS4Is5CL3Q1g/cqQ0jDeC6wXZqIrhpjWEbyaScWfLHhCm+GkGd6Kt
HZE/fSAThNoYaQmuDL2c1W7eBZtA9EPf4ixc0iIBSfG4NEGzcJdCLZBcS0ybxd6r
t4+DDD/2UBb5HJ4acCbkA/ZIcetZe4MTOBCidIUTzgeI+M2BKQ1VTa2OB44ENAFS
FUk/OFfuu95GqjbyfFSvcQKpftnB1FHDhywwTzTRtM8ayNMF/AMuPYP9Np1F4m3Z
17iY29dqk6DHyg5stuW+HZczqG36CFB0LiN6jfNO60Ci5uLYbG3IgbveTr6R8M7c
uISQySqwSAchvBk0t8ZrJO79PguG1w1hb/XYrPOu5jS9Vq9f4U0L4njIHs/v7SrB
EQtnpoj2CCaXkoa/S6sbA0ZDhJOsXw6Qte+5qXY9eoDiZuD6KyF0bIP8/8/FVPw2
+M3WD+cfTbiiOepNK4vFs9A54bIHWVNhDJX7fWnkx/HzSAgws6l2CdLkIAkBJHi/
kGhk2zZK9qX63WkU00uNTIHG/yWsOl0EamnL4wjuRV2hpvkY2evaIerqzSbpdqYv
Z9RdTKJ4kaNQ53ujU14aV2J28cTUbDrNwImQSBytuFlOqUOJHaITMm1sD1/u81ve
iAXF9Y6ej1WzWxGaFBI8zmbhz10YU7i4BSPnrYnpqa+l+E5aibdT/rH/WelahHod
NdvtmN85YJPXgf0yiCXUL29z+vm2Noqm935vhyx8dorVQhYWU4e6nhHPFTf+uA3u
2L9fx7Y7Y+JR6tVzJttiTerIF344eKyTWBROsqScfkRXHhvqEmuEG7JKBgYJuQIX
7b1Oa0X/6F2v22uBiFjUBeM7GTfNYaVaCudvXcizBD8H1M0L7yM0rRkw79XbdZkH
Z1WMbaTipL5+JIy7IACYlWt+Ea0OqQU9JI8uxl17Hwv5+dfvBKEu1Nl0hskZS4CW
FDl+46MX6w4QcwLi4n2kPvXpE41+IpxHxESiGcx3rYhaaN2avmoU227W6JFoLKdk
VFePD9+lfpqbO0y4bVZa+5/uCryKPHTBLpDHxnjrhWwxpfj1WKdypQbYwLruZzEK
SFs9uBlJNd5y3uF7Sn89uLJKLx3e2AdrbjWhbPMt+2MeAPEpuKm6QHMDxj6pUuEa
KecL9gTwXnjOJ0M/7yHsHOMod/4MTVliOZACjkbT03HPUrMW+sfPku8wcfGncU8X
CnMgr3Tgjtq9LMO9FeTQmV+9100fNsFWuWj6hWZ9pqoGE5WP34SQVPZmTjLedx/I
tYwgpV+2YrvGbVRyGSItCrN7dvctUC1Y4xlXWs41yHhDWzF0HR2qBGEaP9IROITp
+vT3ypftlzBynDqOSKvs5DyrTZiz2s1wefvcRKHRbv903DkzTnAVZcRSQ3IhwJ1h
QryRCFUi3/ryV7XPYKaVm188zlxuyUW8jLyf5YxuE09WWXAVjo67KnI+5xepA3pP
zpOq9h9IB/AW8xbg+x0X2brjpzFdu0TDss7yBULoeZVbJWhrCHoS0WCo9CjIh2xj
sS/JEBYvs5ylx+ehj9Bc1TV7/kvxJRnKAZANj+AYoPkFo5t5Pgce/xxo6PX+SDZ0
rWBvxRpSUr24aPZSfitIRTdKyCciJ7f3POsJDhRL8bUo6u3ZcZetbAbsqnbxE9K9
TEFQCldyxFcUUPbZkbpFiPWEiiPEdccmT+1NAdT6IwYg6q1dReJBL2ombHPoKHSN
7pnv1MTu+YKQAaKIJcadsWvM1KrUswjqQ+CdjViQToSEIlu0d78jylv065KVbG4W
NAkRkSsiigH7MN5NPKx2/4AE/drnlc2WeWsVxHz4FCrb4y9rQKIveZVtHt7TOUmv
gztscyXgGARVY6SRxSF2G81IfZ5FrGD/nmzkeSozTNoDJVrTKhzyMVmJz1kMVQ5+
qPGgBtVbLzMnM1xoDvOb9AbaNQSFXVZe4Lv7F4+uI/th4AUCVGFpOttZ9u/39oKd
DiFR6X/5y6N3ReooG+hMtERV+2zOnU6SCJwL6I9llY+q6Ps8xY8VSLIN6B4Pxf7o
dG+6V1dJGB1eoLO7E6p+qzy5IT8RR4/i0/7Z1vgfxyLcyZz3gu3jQGuzmVorNS+1
7gWJd32fBA1Z4kN9V99A7tKPkwX8uen+nH59sIiwsYnPHLwFCFqxabuWS8RIgQ11
cp3sEo6gtVUsbouTxyr8QY+3gK1bS4ul0MlaYyqKR1A/zb8mntUTOs7rcuh3s4Mv
eK4vzMGwVme3XJMlNUyXmkEc7dfQwTv8CiFBqIOz3aj3DJ+mH/aXdvDx7UlW91fn
OoHrX2u8Wp8qW2MDE14FUh3DX8rVL4UvPoqlyE+WL2sUmUJsknnudrErhibnC/J6
oVLXGCNa8hJkEQsFxk20oFosVmDQd6yGfHeKQAUABZKKYOWZTfZVsU5uP9UpEjgr
55g8aFZhchsGZq9IiaclWh0XG30UanPki+j7503/V5KC2NaobHBSjmIfFw+VN6dY
rthBaERWkkVt5OJ9DpeopHh4vy1OEvG6HvzsvS8tLy7hyukOLcICrgNTZjYQdr12
YZVLJC3oSv8uEZnc936i3BPQ3NuH5jVm+gDu+MIFK5HAwR3boDkhheAPcKp/RwkV
1lIF6cbBdKD9yxobjSHJEEmtG2o1xF6V5FlKhR4SHpE9k9X0PajMp+3N+HljVTD6
+v51BuYXmwtrydIuUHm37G0Y8iZ8xPmyAPM9dxETUsUat33L2oHBbp6/kkcdEyMy
CG/gahRFyKVIeBAVDuk27ZsTeO5ZAi580xiZaYpa7CXARXrMSqCOnUJ8daL8qBbA
NtOy77yVIHKF0nAjS+rCPI4qmotRr/PbRAOpp4uGcymwacSBY68KT35wH+XXTCbm
M/h9qOF6lL00IVZDFsGgBh1doHc6/2PjgUCnno609/75T4SmmmC/DhF2oFCK8JiF
c4kQXUy5ZrFHUSJw49fs9N2T7de65wcIEsltDC/Xc5XT4bndbq3buqVUjn/5leIj
ic/SOLt2daacTGE/RoCUcB1njAPhqSTu3HtkJ7v+4+tbDaj7klj6dUnYpa9oz2iV
4dgLOU0R/jz9UVa6l/V1WjEiovi2tiRYOZyE1AEqIpvqPWxoD/7YMf5cXAVatMck
3xMBdvLESALTXLUhUkL4J312kgx85eyf6Z91VtuaNs3iRoKnkCs70MQnPShzEwxB
TzUMs3NwoFf526eVxnaXHFs9kenhZ0p8emIOCEROiic5LFXKAa5omCinbBmxIcv8
NIgmcfUQZFJG3XXNyM0nSWKnsf8tKoQy1GQ0OpGdqQOdMeE3mikq+0/5GG9irQfc
Jk6aJDjmwHLz3dWrgWbpGXuLHAA8CqsiewZporc7nG36YdqoNMGVNnwLSv7dH1wI
C7rJThUFj7tsUaXvCQ9NxGRsbIortrjVDv6KjAjkWAZC+6Mey18fsSy0bzMci/Ic
Xuym/YlehD/k/XaqLJUcQPs+hvjua6o68gZ7CY5bjRmCwzksYqIykcMgXTB6aK1T
iubRcOnWz8gk4kmIoKijNh7fSpWdBGkdrgXv1PdgRP4X/Vt5Op8l4PrMUdxMQpIv
KJK/6TVIInt489wlSKEr1G187CHMyWTOa7xCJnKka+icYQHw82j0KreKe48fRPJD
sf7+PodigosgWki2Ooe0CgYUulbzm0L5Lfh7ItZhNPkrCPlEnKctlI6nOc1D1NNw
k6qL4WSDHYwOJbTDEpYU1wnEs/ta4wwkAWNeX4CGLkREmwenjeC8e6hTaJtgXgzG
eeyrwWJ6J3cHBWgVivqp6QecyUq5VKH3fXYwLYXkrcNF8d7embMNFdAlFxBQnoBB
4mC33+zv3yHJdkjCk/tZJshc3+BZAwqK1EcdVXD4bReQc3WYLVE6+Vi/e7rzj5/Q
P4CwAtzecBNeyDXFmcK+uAsZUIu5qwbCzOVq/OBTIeEOQ4TidWuoXA7Sl0OmOH7O
pCmF2M//jZnrIv0UH+ktIDNWy/w/Ftz5tjeU+ve0ZE/KdRxZehds4KKnPRaWjbgv
tBmbBEc/ifi7lWhUEQffY9u4xzv9zXmmvSJOcuK3wyMqmYaTUBFZs92GockofOz5
H7gmypULLlCOhX6a2l6Ly8khM9NZ3dCF1gbMJaL3tkSCTgASTfrHwOsoNC8pTO5E
CwHRXQ7WDgSZKV1m8dYmxJMrc5UVJvkKnrdTyxrTZd1SAAbVaQfprJ+B3xNNJF/j
/u+bZepSk64xoUCZKS1R3sCOIx+/Q5UQHpxiJBLWpGINoMgqwnZaAt7ofsS9HHfY
PQgE3uZoHVYZgqjRziSngcbaeL/wvge9NShzhbOQwQzAbTwcGjgB5D8+186XpcvF
HMWP1cNQd0Ao8X0vC6jfMiG6Ea5VT1jSC91qbcLijhcrai6d85z2+Ug8QlaTMHG3
6MhB9tZcmniM7PqttJjzZR9UP7nUFrOM1tKAFJn65FM5LKQma97TrXDlmTCcnu/7
NMAFRCyZgfEA9CbLlWCZSaTI5yxxIHKDbQ6QGU03Le8GNLKIT5k7/O05hbvj4eEq
vfKSZfdWrUQOXO5G2FB4V1L0VwylfVL1Hx60qLosewjBiVZ2YebvYsiNhDhoH5u3
9UuHVFKeuRgYoMpK3qhJdls4MwW/xddjNNuf2VWLYu3IMdZ5IEJUyKX2QJshTVxW
vmSBRi7y2TYCui02ebFCnidObUfjsASyGJWRSc8iVmie40okTcQGtni5xxpMm5Xd
++IsjhSL/HZPcnE4Pm3gTOHYlBSmYrkMlZnNUaLIQh67gtHRyts3sH7jbfgk7/i1
qawe/Y5RmrLHeCXSMBTaA/oMC9qkY9ayIDxERMlUiqt28+g/JOjgiJhn8ewi7vWK
/NHNv1wGi+16JFYU4Ke/06DnyKUaetku7VnSoOC7wQQtPmNBuCCGCOTqYiTpHtQg
8rWyDzywtJImBMNWs/hLaB51phW5Exbs3OsSHZDFl3skTktGhTd9pBeJm228cL70
RFOr3294p8uQUJEl/MqeobLKn7Al7wR646RLX1h9ZISkFAoizx4zjBn5XdR3PHyn
0+Dbo2fA199W2AhsC+aQ2YQni1o5Yg2VxMPQ2Ok8ddoXCbEoYyA7l2Yl7b6/GvAd
R6/rndiAalnroIXrrBoN0aFfIZt4cwPlB412hcs31Iwb1Fc24r3eSGEkag7TI9D1
PEFoC3t5cuhuzkDJn4IXAH6ZT9KITlElrmgkzBC/7azOyxaAtdlq1hm7JMmiNN1B
Nh1/CQ79ui0Bj9Jal8OcCe1eSSM586fTVRoWq0g9uKJkme9tOk2noa/cOdZrBS46
4IqIWD67f63SbPMvJIk9qbqpDJF8kyLVBgLMEIO++CZZPf5tcYWe/+UCBo5ejZx5
qdfbMXwxlGAr/lWzV4xp1J8ALKHMi4Y/XKD2na0rVsbS4YPp/NUSWEwqd1/jmrYc
EySpHc9hMVJZgU1Z0RrRzJ6h8y2u/rgcb5pL55t4CV88DX4r9TogjdSAvxCo1ptv
mrcCY3IGnwW+4UBkzoPLtBe9MCRArrsQ8auIf2a09/IAu0TE8A0HrVShH8MEuqFN
cHL5gC1lBs1T5BxspXoFuAKjnAm8Z5quKU5A11U/oP+pyFKaUfATVGuP6o1/D3AG
1xBJJX1SS0PLVkS3x+F0QAFIwxNRrRjRHIr47k8NjclLdP6J9OJkWtP/USYdgbh1
wcM8Mpru0dOiOewaGBNWNhUtWry7Y78BBUAhSdsaBDusjmhLA0k0tL37KHDQR53h
Qzd8Hz/RXmgIZ8o2rAGtPOGfe7NtO9B64p0TnPweOzHsq5zzyvQWcANXvgMdD6BY
TgG3/2eEF47ph45IR95/iE6d3fzVr8hift+wKqfzES6HNlhpyfTJzOdTum6fxXmL
G7jnfmV2V1NT1pZwJJuOYLRG8WuFNesBog2jDIxkbazTWhsVdxdJcmkLxWF41zLB
nlBhVEZi/UQE4hkCOFuaMG/MasdjcpdgVbXKH5XmxZRbt1Qd+BeuCLDoBcSFNJUs
cnaup1rYohhW0+qVZVUOQ0k+K/J+7DnXM2rw1kq9bfS2paCx/OHndrW9Q8Ep+sUj
CdDskTaTFp2MkpgOPT87nfElXmvFfGcqev1XqxfaorcF+nW2hERxkba8VG7iiriz
O0wmjx3XSpjCNc6PUh0QwWN1UKSkXx3JVjOelT2dW2H8GaPlBytzXj+x6TYeJrZN
GWvzdux40JtoImCeCozqExzggYZGIbxzzu/4BzFCIiMZibpYe/G0+NuUWQGmA0kG
vj9BJMVvl+1QwWknXWQVGofm/f0oe7MaZht+gYZsOU/s2mEtwbSw1nu6XLLiFOJn
jb+NkGMSmmO/QZWMb30RicU+2OPSBj55jQVhFjg5v3eYfQFouNnJXYWCyeS/VeRM
PetaxunLtmzihpHQwgBL4cjxUPKzCaf7HqYzBPbOzWKHslIDZdZKz2K8qM7q0E4S
VStE6mbmgZzuslWRTkgLw0UTjl8qLcAfWgxiT2c1PCsz9fXUe/Yu6oaXH1HeKl9N
jEOG6PNMC+NaMrBD4aTm7ZcN01C7IlxsBy2LjeEFb6ckUIT46sFPoYzm5FzmqS1E
+GxQCttE4W3wDPfBgva1Mhr8Ryfc67dhjoTNoEuInNr9jC7ucu0BPBxfJicCDUt0
5Gs5Ak6yT1mvBKHdr0FbB0la7AA2sJWYovambObH7qaP1+3qOQW/9abYmQQdqLDM
jwgwPktgklIvQPScYxVHQlvgJGl8oyjBSWiEGJ8qdMthuTvKx40ELvMq52Ox+uxx
R0mdoxkC/udVp7n9nSF+AORA8CYTiR34ntUox1h02FnQeIps4BSsCL9IQGi8X/KO
XbrSAf5spnq3ydt2AxXskrGkX0WocL76usqM7FI+IlRrc1etmQbc7heks9563tbj
TifS2DwYqtTF1iSugpZiPzpeh7lzKoDX2aBoODaMUu0bWBZoYf5w186C2tv0O3Zr
zQyx5MfGnCPJHafixn2OOrmes9v2RIJcX8aFIt/qIz1uu53BMibAKWHvTe7rjnVh
pPOZNvOarYX/+U+4BPIrXLJzLhQQH82pPLDSU4shAOspBfBHaXqREnbGVG95QthQ
qXhBkH8oHb8ZJ8ABFrfsryBdMhwdRPabGeL14YXe0+us8VJ2hz/hA2oi+65TBLX+
3GwxeL93BBxvM1+3pe8LfkU7g3itjBq/AQr86CSFhFn4Ko+JzyJTMCTivyb/KXMg
OOZtInVMEFsGuNXq5Qnj6+hot0x/OEqURizHiTZ+RtY5mbzyNvN4uPCngbNgzIHA
NXhL9vqjDpbyjRNreAeLBHDssKkihj+ng5077WxJDUh6RZeSLJO6qJhCoqGaEpho
h/Pj1NeQ90KsvnVE6y9BYhrFtNfYNEw5rscrKxKbqGJTm2AymWEyx6rOAO6HjZki
sUDzLQ5fkPjniRWyNCktL1bNvoG0KXJhWt7LZsDpJzUQcoHdhp8HrB2WymS+mYjB
lMXquqRKbfV2VUUMP79GLfjL6xfoAvTIEZ7YY9sRFpmG9YYD/FvcmX8ZLkKzBbd6
geKQJWHC+vvn5SiMhvFpaGNUv862qLfPJ2OzBJqutEsI1DrAWH7d5tMppzxS4d80
ObnLwQuf1NSkm4qG1Ff6ktd6IAE/iEGW502gr4QpR6ecWKNTOpxPomDAfKEr9vuD
HwBRsivBhNvNV5x853t8ksqGAjcdTkO8P/Ur166L18yUtdWo/X8Tm/UB6upsOaud
WPoihghuy1qnPpZnRSokGSgW4wFXorBtOdfZblR7l/0b2Dq8dsUS4UP/xTr7t2AP
pqTRqospvShV/J1O5ShLJRl1gz6MF+HVbjSS9mwu59MIol4qKa5GBnrT+6kYVgR5
2dhRtc6woei5xftEq7VQ2nUL+QeNcEdao6aXT37apkF2IbR4zLaCL+Agtj0/fvJ8
1jV9v23dSS6gRaUEl4thRZ0mKX4b/ZHY89KcTrHbZ7IybDmwPIIC0R93M9GSVt0P
r588uCFszMk9f+qg3iDwEPBhVoMpaSslhfVZ032cgAy189+9TmJ9dDjZ/RSYOPUb
X473rZG5RXI70G+fy/hCy+lQP9A2n0RAscn8OnO8IF5nTJx0uZva8WogRuY9L1rH
AGhcHJP0HxREVpwzykIAnQTWVe+vUTFDGQv7+c3cxmNIxyDLwdEeRtcObKjZvdNV
0EIeoV3jiIcRpkgSa5+ps3F02gSU6n6+l0gILVseckCt9BxkX12eHgQcB7QjsS0g
4jVOqMbBB54Hl433aNog3MKr8V/g7q0CoX+9tgVJcbofukZ7BijrOY444K1QZi9f
S1CXYeXdl/6jNc36Vve93+InQIk5LD9IyQ3vXXbKjxwEte45iGMIqcpP4zBXCNY4
7Va18KMnd6Hntkra28ZFStOr9Tw8egGy2AU32E+LU9ppTwIMdXiHDOhS6ev7YDgX
SNIMKe+gnyafz4G+dTmcz35HGDtwXmKAlAXLKKAopjbr8hOXYTIFolRqwd4/ZfxJ
E4JDkKgHvGVt1PBd0mJ1kcivfqB3t5gA0hEigNxDBtyhaiu33FjaNi7kxiXRHao4
deJ4w2AAQ+BxJLcplWamhamHj50+L5ovFCYIEUZnF7d++/mlepmI1wLtkrgQkI9I
yx0U3vb53NGqfC/9kVof+xiBPRmbTA9fYAea79SMDMXVaYEGd5h+mY1X89479bwf
NvXldvxeRICxgWUZwO3n6x7rOLddjK/8m9L0LyFQ6h1u8381Y9HWJjqvbMsU4njS
501PayLYCaAJDfXMh8pk4wuR7HnvSVE1ERUsPDkh4QPDruNtGD8n6ZtDiEVk9qFr
TK2gAiUkeq1HhrKOVfiEB+FpHEJ2pWKmraCfZqnbp1ifS1PAB/dckxHwU1cHX5cU
5ayGtBYFYzUUlZrM+w6kJyMt5ZD/2KbPdqHQkmtv44JuPcSDy2tzKpQ1XJWUZ820
lble3LXZsP4sg4MamLmUwE4HTCmPHUUgocP/fybEYIHq8F9nTrAAHv4Gx8MfvKt9
V7qxT8KUMk9SHqdwhTTdU6WAjnN9QUa9tCjPH8gG0QikgAG7XnHw4Per7rzMb+dD
9K8paQRu6+5ca8BhzXHbv+OMd6FBTNxI8kukOnZKMOj7kzbz0goFelZ6+XT/qCkH
Rs7HfkX+sFAV0iQljS6TbZMllQULsBJ6yyHj/sRNWEqXj7BM60cAgys55pxGRV7u
0n9DQDvzkm10hJUIUEHr0LX8g2G2zCjHX/Ncp7SpXcrZR4keeP9tPh462o+8aacp
NxLfkF31pRIUzBdPGM/SZs59FDpz+d2uQbGOTJMuu8hxTqPthCKVCjBW6KerqHgm
x4fd7ru6fQsY94JVND6geySQi/BipVKqrV8ZWqtH+q5mgzsUCFk+vPxjOr6j+bC1
i24AIYDx3y3/RCqc9N8CPiREvKpI1DAIP7StJUD4oV5gKtF6bh1HlRUNkHptvvLq
wfxo+LpBGx+j2rEB1mv+B6htBHqbylWWRjb7WDH1HAiIVLAQoE0jEQqDg9V3XohI
RKBq51tR8B0UsQnpOGe6d6w/YpoJcBbW3RgiWlkXgmfHc8iXiIztGWCznLPBzUWC
EXRZYipiAGu2BhL7zfOM2dy3GOVF4i9FbAO/ZIqqgI37mUXRZRtYFfRwYaKNZ2Vl
O/v/UVSovO1wAf3yoJKciHI7LneYCVSe7icCz6QXc8r/CNIM46r4EOxFtK1FnUz0
s+XiF53uttNvQC/K1vmpGTvC8Rr2EpWpqTuU5aIbGgIrggJvPGsdCHrwNkw3lQh6
7wLBnelicKt+oD8L49ym8LVjtcoiUrEL7ucTMQxBtm2L26V1oTPslgv6Kn3jm5YQ
lv5hzSoy1P9y7eQBHJAWxIoh+WFEhNJ0G3zAXOSQORI+Z/k2Zsj7OLDEu4JchP8B
co742uoktmmwc8xT1WickR/kEIBUwE3PCZYlYqnh0YuLTSvLpbpQ4KVRRoQiA6bt
NXUB0UHfkvLpIarMTY5X75XL2W8CeQyBzcLG4QWCzJKrkOBOgzHbMpptOlra37vo
Z/zFr+rOYQizOqV6qDRRPI+IS7nNcfWGJ4kxL2T/zafQQFXEcGju+4afw3siQrN8
QOytP6pN3VVYJ+SsYaFY4f1s10r938JF9A/ceqPFQK7ZVMFHmvtteRdH8hfkk2iD
H6k46dFo13fHTa0PgdzyyiXbTUBy4/Qiz9VjNE3xxLJYvCJJ9g8rPF3dVcQ7EuF6
J4JFL1z6LZT8X0zF9pR6kOQ8xH6Wg7sSl2FBjnyk97DfjEvbYodegrGZZD7igmmf
uHF7UYErYbdMoUvguRaNpbwK/EO7Jymz6QF77lgOSV1q55zKSk34Kw/MovhUTn3v
zQG7qDShXgTZ8isjodLvHXqKAeHOoJQZ6rHTpxOxnn03NcyvYmlnyVsQmhkMr0Rg
YgvmRDBaiVJw6pjP2jRVseJkVUsLafYThDPkhua0H/YB2brnhvIo7FviqiEu0ZdI
xyKUGkFtMdmLXEOZQolDyrwctoUdR5sRnEdK86K1dC98GfhBvn6dHN/ALZ726YQ9
QBHdH3PK1GTqZrrQdjp9G1TqL7Kl0PCC418ZlZu0SME4KTxd9HuFW71KDqv+sU0E
oxV+Q6q/WkidKRVtCnwDg7c8bb8e+z5BiQW3ruU62LCRoAsoGRQk1nJyg96yQFhb
Yy5RWlJ7UWCWEF2AK86OqIRVC1PqT8Isc1xBNGNocd6eCvXyQJ8DbnmPuBFLJ91c
W28eMoSgDrg4miPw0pZoJGmJ6VnSiebfLfc8GQ3mHQSuapzxWDHdjvkXGY/MrLUx
L6PjbYIbc78RQrjphmsemV47j0M0loH514PCfZw9KOYhLNwUTukip6MbW/QNqiWH
5M7nUk7sSUY1KgWDtqW4ta9Q1nqpUNH8VGEnIH9dZRPKYaVSotB2cK8SSLgfhXFf
35gfohb5TgmwRm8TIgl6/AAiqXrBbYpnh/NBMzQ4+KmcFVIREgeyYH8npyXto6vx
6ii2XWdRp7XaThZlhyqKYsTV7YftN6Icg+4LLQdi/AgQk9QgrX69wxigxeRPFo+M
qrIKQiawRAYZF1M0jf5dfa6rHgSP6OpazaRVVL7ZuNheo3+M+a88ZMixDiSLVrMV
kytjoPH6pr4B8/9ZcMFqaomDlLXF+WjgEs1uw8Py54L205R7CXztvR8HU2J1optm
ZkhCAYKgkt88RJd/84nkXlg7cPoac8tFSEp6WrskDQHr5WpPxhKxR5KrHOBmaV+o
4EiCVKfzFrl1+r1otQmeO/SITzrLooBzBU0jBBZ78pVFYf5nV4RzuiYNXObbVtRd
afMgPsEmuvqi4h6QwgEtOX+Xtg2KFhTobk1mncjn3cpFh07GMwG8MgjYHdPO97Z3
2A/elAfaKchUVzF7T578nz+qPMKT/EASNP+L3EeCdSYvuHFT6rIgY/1qG4yUPfx3
9mKhose1BI2CeVTS7c3daZp4pfhWAW0SVW8e6ZLiK005XannFzFmwiUQCQ8dTQbH
3rUUO4uq8t8JU0JAOGhw8mWtA5YpdEmOkEMoZ7bPQwCqYyVbDhaKTH4EqCHuGdl/
/2KqLVSgbqW1ZmjitAHtJKFAV8Kikel0wVaWiRhtp/G5ZeECak8o+DG7bl5TTidw
aX0wPu7RCggLTHoUW14nnHIuxU/oOwB4Ll+VmrD7IxqZK6T1ds2drAZizbAXeai1
fQcT7Xd0Sy4ruxzOdd1cow9VHHWcw3iVz2qsVkVQ4fg436gEcaLJxc2ouzCnFcDQ
bvPsNX+n00YOOEii98g+Y6MU39EfDzJFkmx48ru5VfNC4sg+q0PbhKFEGL97hpJp
CYZGolrnZu15+kuJdZK8FFgpg6Uc+CkAwo9r1SQ5PKfYsePONuUTSBbXlWv2w22N
kR0aNow5M4dgndf92hGN1p3DyUPPjt3pSzgTm926RMjtWNZpp2vsTxxMxHqHJcku
dmSzp5aWuhhTedIFvHVgtFqQ66vs7xcccJkw/djxyGdEVcNLfWggsqqQhJCJ2ibn
VyVOcYJB5V8UE3GNRnBAr1W55y7e3KERo+k/Q9ubHmtQC4U80D7v26Q70UdfNiG6
fddmnUI5yKp19JiTEBAhV6TipM4uOV8pSbW3ApkE9sbpLs2EYzalY0cleD7QY+lm
fUd7lWjdfzTUhAozcJPrXcyYHr9Fzw5oFCxALtKPzjuofJw6wbnWh2iReVinteej
4NFFRY/zLw7tm0DB3E4GqSvVY1jg2nPdwG5RtWWLY1q7qv3dCc122w1hqoHIRHmO
sWUd0FWMw1i4+WNNDUSojqMOmZAwtj627lsWrbe4GAG6vbljXUKyS4UdnANaPdni
J9SiH16zYpF72arXcWvt8IKSNWINGIx0/tAy9wn6RFLZcZek4aWDVYyx01EQ519q
/+MkHf9DeWKGxXU+JHxVJW5VrDjJ0PtvquWn8HUArLBazHa6IPBQdvdIwMczk0gP
Lr8kzNuLbWG7YGt9iS153uOxc7f72bjBWGHuUkUJ6qF6qf6a2SaJ60ldrIap4i2z
fjYLZhiJp5u/La/wQsoMcKKslxAxrS8yvsUFcCfQVCZvBk5Pyo2Qq9jpD/C7SBOn
APzP1Ybk+UoEEOFSxJsK0Wtk7EVtiDpO9pyOwONg1ksyQv0DzSd3I44xIb4kvFJ+
eK8txXJVk7iU1nE7I4j1H+YkdpzFEZMv1JBBLJBSJKOpzLjgf+N2ukbQKoNJzGhK
9k8siO0eZASTARs4mzrlyyTRlDTUOG6GIpc9KtppuvzFCqAx2WhWTXadO2hHnVXD
bvJOC7JglnNwzxV/SscBBdju2c7y+3661YqSDmIOCW/5YGBt+HPE600N13oDGXg7
zv7WRkMmk+aoDAqnn3WYRFY4Z9mETL/ZaQWIJ+iYOvbxWEJruwRBgfz5Aq+HuC6G
hUD36qbtUAvdiRJ+Vaio2HQBDo6xsS9qrWVlU0kZJBNsjQLp8XeN4u2VHj1cXnXW
D7LKJ+3qkMIHcbVLICfVuanYSv1X1pKbA+7/JEfHPQTp829zqG2mzqgGA1vG7jaA
8oxc0+29CM+duEr48ufGcC4j8gCqF0U/cD60duwI274NhOxVVzyb3fZQ0lcc5Kek
vUrOqjvX2zhj4JVJ5nxh8lLPsSzyR5h8Gq0HuksjH7W5FGtcaropJoBwuUQbFDhX
cWv4+mqhh6KDdnNyemJNGvDCWLV8t9WLl0xk9xP64xrk2WhCJHVR89DatPrYd7lT
rTT/NAaSjG49rb+O2LtcePzaOZxZQHai3fqNf7uDgNWxajHq3sQplecCPM5FNRxq
EVFgRN4hlf1elbcPiexTatIR50HxTeUQHwbQdSj5E8YuWdtJQmVDldjEwswdBIkh
qdhn2eneZVeReGPrSOoGdGj93dYcU0UpBFOkZ9sn3mgi8LHO4p/c5IcjokGn+IMs
lpSSmzUgA/7EGetuPk0odgz5ktdLJM7W7TTorCB5PBlXmLFj5JI9est6I4atlCxS
QcX+bwNpx2g5fywBwKGx1bbQRJ/wTeDCzbgJK09yHiURkNXv8dLaBJbO0lx5g7H6
ww5X6RWUJBpNppUb8mqi+IQ9e8zdUjZnQDpdsYeDm0jglZuboekFJF5UN48+em5I
11KdN+LdciOcAuANFQA6zQ7LStG/hM9ASevl4SeFt/flsCZlv8kEZjYfzA3vMwOC
LruJLAuLzrBJqL+9lI7M1FZQdvgN0WMAZ+/hT10CdUCUU8qgkM+6eu3yEH/pmMD1
5N2YGpTMjpGKBASJt2/iht277DIhyDOu4mIHtuqSN9RjxmCdyoUktk535AHkZwy9
JUVVskbJBZk2WjTcVJZfll9gM7qBJaDkJvq2eGTA4cnozUvJVZSADEDXT11X2Ll+
I5oXdbkmJtxeBMEnABOVvmagnprOEYM2X/onaqRk9LIkDKS2seU3p5btnC2l72kE
4laPXgx7m7F+QppWJQiH3pL9hsXJdO/4heAIJylYiWFMgCPS764oMgvs1W6xcZ4V
COq7+TBvIqdYfehm8z2XgiPo+bTchrVyhlgGqYa99Ra/83WkUVmhgHAZpTWIgj1C
tmr/lwVSqvkd3zva/GFUiNr3XTCk6gqXcWtCONEsnAf8G3QMA+MRU4QuW/l6RVuc
+6PSoCY8XG3Bs1Lx6uvTJOjTiiSo+Ps55ycXLCfpKsvNkjt8+nJrPdxPlhMbooC/
4Lpeq75gB1xp4FaU76UKtlFXIa1/xiOT7J5wCxsGd0G+WgRsR6kksX1kFO2fYMLw
9yxN1O6Oc475xofVC7eraAtoq3kX3mL/t5PtijHFApBnVbV0PNR1BLe/Arrlhc9s
IfaS/fOGITL92USI6j3oEGeHsPSKEKBq3+K7QDqmlMRIDeb7QlzqGuWV6K9BOTng
bP8PrLmxBLF7yMae+eDcUfW404kOVoGEzURHFo44gASogjREMeVBqQbYJfapsIeX
xLtSKGGlIp2FWcbZunQYbMjod03xTQ1G4vWl8EIWmqMJuFQRxUerO00496IgMjS5
QgpbgbPvXmVhsjDdgQYZvkeBRXY52axXFIbMPjJUqOQq65cEzlQx+PQw7lPmFJNM
eDcORlng2pFR9sXCgBl1OflxxT/MtVvHNlvmFsqKvhcChm5iJjxzirhkenpt0qpr
UNr3jes0jq3AxmSS7OWf0Z7iSgDBKB71uRqAl7J57JYZ2r6Hupi9cCETgCtt/HNL
Loayl3t+Tv7QihGCy2bv80kP6z2QA5BWtekFmEFoks4Hb3dwTWbewJyxroPHPLxC
XaR8MW2C28bSR3wjNKgZIRah1g79qz6HW7HpLZgrm0Y7ukda8GW6fCNtKHZ+Jj2D
MtGW6+vZNU2dZxwSESX0PBadyFknqjyLtlweeRBrBEA9isb47bIE6gmdN/4TEE5J
PiuuF7J3VQ4tJMId8xsgtUEJhsQExXcrfA54ysUwk8mbTkmOSLlDKJal2KD5oIhE
LMD2GAOcDBRKVhhNODbMy+rhYy5tqWZyGsO/I3xYc79/fHjx71yaX5KLG2ocSzCy
UEazYrHIcMmua0JeuIG8hYt0Ka0w6EV76f85BZ87lYQ3oGW/EsRBLeb5NyPZbgqC
HjLP1k2lsAnuK/wllfvqVF32f3X0tCAUDk2wMpRzKOJjuch2moPYgsEEwamTRW/f
07Z6FnDZz7q2sJ/K0JxYox/plb9upiwBk0lAo31rgIWvVwmaUlBhXcx25Mcqn6G6
ABbGLs4glVP9NgexAVB3SJkoFatQc8XQi+SpG+F9tNrmF1IZcCm1hgS2FP/mLIgv
9mSCnJ21PZ2A/9JoJctO11MNcjqoNf3XSO/IBhECTZ6YkXdkZI2aEtt5CS2aelii
HTmakL0vgha6F6bjy8GtO2oKbgjRF5vELzG1iF/m+Am8J2W/A1svJ97juCgKEzde
SD2EKq5kIclAp0vnm2UWrh9TBvGTWHyz+CQDeGb9ctfb4ZhT0nqlrw9zR7PSYABW
Ee1t6BCkMYDpGMUC2ekOyQqzYMwcro3DvKIAKXLrLI+lrY8B//BEPIPTIwoQRjen
HfbaE1LZx9sGnLRzgNt90DSkpCZwhEVfr/vCSsXB+OoSAxpTBCXHTjiRg2lRWvks
UVQ3AX/LmDU1g6coJvAO+yyLVsX9rl9Flsyg2ooH6HdvQvZP1c9NAwCginv3AtxS
WeZLaKy/Id4/1BiSGoBmZDJ7vYHfFDG4GdVds4GZbHrxiKbLQs09kmw0DeLF8l6p
jyJNRM+VklCEFA7OzxtvuCf18TltS/C+mB8KDQ/SY9xAdZVvyzWmJSGiLOfDA/U9
6wUQ9E2RLoNbUjfff3LIseDh5HzpvpYSySMctFeUZOPykhhl62I9gm8KnDzCETZN
y9j5TeX7ZWl66QeW1hnC3JEvJFrN3I4uwavHfvfCUiOFAs3Mli5KNUgQa9EFZtn5
5nfdmPAgPiOiaGsvylxDC860j/6Otuf2iweJOWLQqGEjF6iVAErTSOy2HIyTCTY0
f09/lglm2FZers6G1FCAQr8rqlbtM7+JldSZBmiJk5PX1KFg+cu/J3UW0f65a6yF
jx17VIWF3KGpVy8mJhpYGpxh5ozaL16PyNYDAHOsD9d8GxtPeohqZR4J1yzxp4Js
yAcxWL7JKhVFoiSSzUdHnUXOz9nzCrLwEqxXD64G2P5tYaykUaR6Ys8dTyRUJlcZ
7edoc/cktz7G2lsNNn6rSxMRQm0A8un8FaY1YCB018plrzdjW4DDlc7jabtrC3Io
fX577/Vy6r86K0JqPgvgNW1ogt6G2s7BRuB7bFfepwuXfW8M3O64Rl3+bJ8Z39rM
3dOvS+7iTBfNx0MhSmEVziCXqUr2eE9UHFWGNxwugZtsCf+BrtCd73tTEtlDGqat
pDawem3QDDoKfbVXlBJzGk4l61bJ+w0QjQugMBmWIeStBLGuJUTixzNS4sMRQmUn
ecaWdEZG1D5wQ82flZq1g8mDOpLwb43GS53/UcXfTUKkDTf5pxrFjVRs7P2wT6jI
ddkG+1IU6vREdDZ9xPbHxgHpLpF+qHWY9SWFhbWcu7xobGmEk4dw+dvSrsRLBk5C
tTCBqheKC9XUBpzlQWdTY4/iDxHk3qpcHKy+m/lZrF/z9R8lMXmN7KLTdbeJNdZM
fEbEkrnAenuaHqULfVXZq6S4kbO/cY+AgmGQIOOfQ/+3MabsswoPKU+59REpVrr/
bVsSKvQMQiJIIrJCkj9d6GkEiwikpSBFsh7JyhhqYtVsMJX4QuKS6LidARiCgB19
oTFp2f/6MGDmjrqVWIFdQPut6afCt4T4n4Zbnt8lT05w2GkhEUJCyJrway+jlXwu
WFnXfjKJkh6qd2IlWhdu4pnxFuKJrGo1/vSrdAF0XPeU/Ak2ug0RTXLfXa7Xb9jI
GaHO6e7P2R98uYvrNLhy2iyfHXvLTB665DBj9C6/G1IC8uVuEkkvPLoVAtTIuKuB
REEfmy4LO44kGrsbJpKF7vAjVUSMQ9yu0ugJ+8wOaQxwq6Sn+1UKaLkocBQE7pH7
8xdAC+AwZpGTwujq/HN00osd67WRIfworn6FhrAU1XAj3WDHViXEBr/hVMXdX/Kr
O/w3ni+2lZO9JtmRvlfI21voRk62qNpG/ymsCPcnNtvBIM5WQ3ZBPnILKZx6HdAX
VKY18SaWTslPYSHFhOgTJZ4MN3n7rviPU0vAsO7lau81LK6nvnHeGYlVD6AHUdg+
63yfhpFT212EYIoIPP5EDFDMW0sy1F0FZH5cDuM3knBtOywIwZfJi720yklHD5pN
oFHcycLblV5yQRxz6vdJxgXg8hJcLbfX9whYt80Xvf7m7oyJkvNU9fJVciy04m2+
couhuM/NupFl46TOecbY4JHUo6707/UYzBMJMyEF64pnWDcCqX2nAUKbSLgvrtN+
FJxG8dyFjwsRUvWx/gV4Yj4pgTaFmiBuLpy4giQOa+gTvhAgCrZy3rliMZiRKKRh
V76uds0+HISj0RxPz8GqZ/MzzGQNqEoWXLfmVDQLplE8al40rP3GRsm3FHmToiln
63OnsiQu+Ki3bYr6RoKhxnlqwUcxUPJVgAelVe6oJIO+yJfORp7S0FufguJNeFxt
WzP1VLvssx0eD8lqfvaZH/+g0AUe7lcQkvT6Hbs5nXPRSf/euSWI25MXM3dXtDy2
o0TL7ZEwr/KjjpwNsndKaMlJSaQyZt3j/M35n3uxYLy0GFWFbJYBkU77GcAOj/dB
h6BPsOWohkrPEd/iHEBau51GbpI8CJ1mdkllzYQWc5SdOPk4HLf8wYZCVefj3QMx
fiDjk4EMRYW2e2JAPsWQbdndSg+R5lM3PwOu10OIyoG/g1qeoqUBVIamHyCxu5al
B+971Da4n4hgzOLnQqE/11+wDM0Ty4+wQhO+P46yF6XLmED1hg6IKMEke4IwxzN9
A0FYuMxgcSQLS5bModIjtFEA823puuhKDqO7pXQJSEEvVASB+KgoEQFcqqg4E7ZL
7PbDgxNGL+9RIHke8lY/AuXO7heCszADZIKDNcESdtNz3TdYehPCImHMNS7fINsq
iBSpG/4pS2kDBmLasQmO1k+zdBs5IyrvOk9nLSisoZ7jQOWwCJgB371dHig3qLUX
dlHNFr+XYt5zMGMRXnHEvGNUe4vmRhCdPnRi3epjUw88/yE+e4cVKhQq3zFY5rbY
GwmbJfBwRebeO3t3elHxwx92m3HokzVhOve9vdQ2EXzH/JV/C6xyQTcqBRkA3sa5
eFQXDtm9Ow54WQhV1Evfa0LozyohygLgoZGEFKNQwq3/xWRGDwl2Pep/twUDzu31
N+CnofL0LQTp4Hefe29Bw2iGEYzr2yt3O5//45bJunwWi2CYy7Ku1Xm6NEJGSQDq
mp+zrsUVjUPnb01K2GztMpqAJVV8D7I/C7hprlvrNC0db+dGnSkilpHHivSkQg4D
y58pDN64rMo/nHGfMZUFRYYLKt0nclUDhjxLOZ0FBpZyC/heUanSJf6SDREK58J+
6DZgK9KyEX/ayT2UTkyAQVPDbEoxSZrGBTy4merKaeXHajEcBrrLq96q8F5iNVQb
HQSz/Bhm+NtE2aYhb6dcaNcZLR5IlJpDT8VV3GhZ9zgADayEvPTeVfERx8TTMPX1
uTHZ+Y/GMRG0p1VE2YgiWNAziDgTM8xNIYiLl/rgnrK7krHu9Vz7CcY6XGBBl3n2
odT4JNvEX1A3P6X1ausPlFF6er4J/JxxnwKTx5xHrpaQMuUVADabfe8bFbF8hnv3
p00B4Ihq+g5Cn7W+4moKXa4HemO+BbhRrr0sufzXJmGxD7WiDO7XAvdxGn738xp7
QZZgo+2jNRaig5w6MCO10pBqdpY/fp5syLzipcuotILl3qA8Gj9Dqql1Ihe3NO4N
2Dlk5pR3bNoc/2ZyvcRxq5hJgZPXVDCEBZTfLxaQBQxx7vDv0NBdIwte9yyKLLsF
RAhpCzIXHbA10ZcE9nxY3LovXdPvYdp6koi5NSNDMIJ/Ut6XJdoesLmuQiTEOLGv
VKhnbDqxCfAvh1mzFj/imiBC3E//2PwoFPAGfJnZ6Y0CiWRcUWNQbj6r8vdl3Ojz
7rmBmEQO7ARkyyHWHzYJNSg46C9/IFbespHL6BCY1dJSjJCD0S/rMxP5HK+5yCsW
ErRCFZd+X5xEaUzMFBB643P96l/Nf7iv3fH7C0yvxIAyw1oxlmaTiFb0gjo//AgK
9bRWorTtOJuRp5O7Xsw4jhDAhLaaOkktYNmnNdqwSWLAQqGIJD0/CiQpUQeYO8ob
+azeRT2rVxkO34bA5IUcm3Yiy6Pf6NpvTLvW/Tr7nnN+1mceKCmAN+OiHB4IhlR7
rkigrQyg4+mEl04TuP9wyGq1ixIBQzRL4khaSSOHdrwC/1YjncewcmKfAeOu76bG
lxR/Ak7E/aYwE6fl0PqX2uQ2/WSGFJw8D9g4a6ocPrSEoB1W+UDvMlroMPvoyFvW
lPDQnrhhYIIQcy9rYhD1Q1QhMBNj/bzR3mJROnrvFt7gLQiwAew5VB6jAgWzW8nc
zLKeiGTpIZoPWillvjHNNPDwR07o4Xe+pidwlFKmsL3XwR2u+pc0eqEpqyB1w47B
ybgNp6l2YR/Ed4cLxgaiRpmCLt9/edOQVWhMk49Yp5CEApvD4wQOqxMvVdwpERda
x+u5+oHxX4Gf9oTFRUDln+y+BnZw/hfJ0utm+A9NoqpZPiuOWVTFbTet18vXftdc
Q/wQodK+dlEhKO88CCZhI+61kh0yjtNhOK2yRdnBRygogNfGOPnRTC2x49yVVqUn
Cd6mpJ6hnWwYsbNJwc3m9F8fc7ojveOZcp/gtCrYlDVo+Jej0Blov/km5IlzXZ5o
2nztiiq+STeLyejAi+Z0lnP86Jpx2FbD0s3ClBczOh9mXyxIe6RndCZPWPggfBQo
4Hhq+2D2b4G86MqcXk3eyPm9+qdbcFsLyTS5oPE687nuNwju7RCO4tuEYlKW8WjD
JA3jyEdQcTNViV/qT9bR6Qpr/I51ccdGDKkyf3g7HD91pf5O0gJC9fS9IT6u8PcT
0NYbdi+1NPZSBFZ36w8Had/IaMnENLvit/LhocC7JD9ujfp8j8Lbd4j3evyL/BQp
gpd3O+TibiiPyUoiwiyTlhJx6lbQ/e2LMpjVZa3E0EUWQFK8zCX1w9XIk4QQJUrx
Dm9rCpXgujQJsC+IZdMrjxwIOArs1NLW3QTIjXAuRBb8Vn+2wgzeB0dZ2CaxZK/V
ORwktNIUUEoaNDmGISbHI3JZq/RMyIbWWKU7NrK8gDuIso2CswbhUuJgEIh+nMUQ
wsCOgpECRO4hLcbmaBxmTb455aiTup9MNf1KMD2F3Ft83dldyVaZjZRsK7cFCpl2
UOBrRfpADvkqf+nir4LsIyTlojaDtp2ktQjl/C21LtLMkpXX6w696hJc6/nUC+MJ
6Z8op9j75a+Fai/9dXrA4Pdz+y0vtVXeopYjQyx6KEfG4ap2ThwWUvrXg4xdRfW0
+diKXtpEcYLMRwal89+eZxTwkaeXeTM3tldx36tGGSxs14KCzjzzgb+aM9FRT5M5
4IbgjA9/rPNQiUjkUzd0bv5Z5gF8M25/z3m0R5yvH/DtPGocoV/BJbbzLxmtHxAa
Mry7NSXGYZEk59WUpE2K5RvG6nbPAAk+PSBlLvm6LqlqfbaV3g8DVN+fiehz2gW+
/cTIZGBbr1smfrWKtMmXuiX66YNg7mCs+9lk+PGFbd7gO3POXQ4VED1xYLCya7Bf
z3qcqyS08rwWvFbqub8fxLg2GMa7ILkIgwNzpB34hkQeinCdr91HtlOhIZaZG6Go
XZ2BqxnqVr7l+YG95ceTeL6OzCUH3CvorUPW5cElUO6MYpFjSdXx0kR0xauElnG0
8sSobfw1hX5y7A1uUzn1mgu5s/5S523vYX3ajASAWjgkcZzDxoug1naRL0Hf1HNb
KlQOilIchwtpuiXZzo1NLY97xrny8JrpdVTMMGdeGiFr+9hyYm35DcJ1sdhJcIOG
i8z1eyWJ+p2Tm+pBUA6HbNQnwtH5SGooWXLSDX5d7R+LUBjoQ/kiaST1XrwC7aqU
cZay77s5rgfRGR/7TDqM5zJwFgQzpTZrs6ow8UkshjNNj8pco8qBzaj/4SzzXPal
12V+3S0Ojem1OuCQQSvNCHXWnJ2oclDn9syN1XgXlcYMztfac1Xh6qEYbWtxv0WO
JkmLqaBB67ZqBOaP5SCxUDBgH5HmbPZE4ABDn4cOvWGbzRZg4LYo8i0QBFX0IeJe
9lvRyrRdbIrU2Otfj44Ku6wjg5FBYDwL1QvzWsPBIfrj9tbmsDGaKbMNwY/CmXgO
XodyOQYUmShGJEz2tvqKrBFcFJFEw11i+Hrnp5MJHHeqdpVjQ/RtHapdqwgSbvNQ
zwSKPN9eL/h1x+DTBSjiJIYeAy16qZ8GGqJp74lkxxG3dPrBTJ9FjhwNipvHsmD/
5fNXfyAUIxsGUCimDLo7heF8sl/4+1qv5INyQQxt8kCZ95fgToS7savMthDGwXDv
XM5UVmNkpHgOLZapg8RDJOKdcFw1FqnuJacppaW5nmBVhjnMuMsWbB7HaQqxvtrs
fYkJNtvfUDYqsDh2JQVcxhRKUz5nUW3o7CCzKJcxTMBKuJGoTYfB1xe7iyJyaNwB
41xYdU8fW1PMSbBKY9AOSHRxIDbJljO0iL59IwyMsK/0EWNnF7RHqs8/sfDVzhSC
ahZTvGwoJFrFKg322HX8LfSUlzOCBxVGcMzGrH1lzSENfzO9ozFlFtOZtxZ2ad++
W6Aw07peDQU6rYZ5ji1/7TPerCvqWxCuU5ZnLPAbfTeYdIRPmKXudLFPEFHtz7cq
C5K5L4Yq9my/mMmI5z3pDXqBRgxYJj+nlTinikAN8pW9HVL+xXwq4ypRJNYv6F22
VU2lHbVtpTXQXwwKxW4VllVlqdmXU/gTl1JOwcVcliR3y5cToUZM9h+DC1XKKqKT
TjKf22Gn6rJtE/4iPNFU0IBTIWzpw5p+V2hmKiGD2ByAEBb+BpavfW+yQLDJlRvT
Yd1Zwp4Ycj6qj7qXOs4+wGmUZHh2zlgKV2zDo1q6aNE4kWSDFfyvS82NJ7tbUIUq
GuqvfMuM5PZVjVrvrYUUIKmmgb2dn+3qRkDSgFAeDXbYDz3mJ5DQUnmacA5kdgJL
UTeclo0S5up0ogYCkhlss57J1bcPsp46yAqDc+vmIiexU4A+zOUUc3gbueOuRACm
piRpSrpBvkCtS61hVR2irwW1ml8w7ge4K9XsTyd1rX1JFdbNwuoAuC/ZWxQPB2H6
vhglrirB0RZynuydfwTzHlvyxo+o1bDp4p7bOykIehzM/AIh2N8qQaQDWwed7JSV
IqBODit6BiBIea6feiV+8aLt1Xf/p6BKTSZ4p9DO2YH5VSgODykht6394fNBVpPi
sfrjTYtwddcbjVXmSuop8oc2r78K34+5y+kB7srMf7tsmDB4eUfzidWAgdwcNtdm
lrtCZrgeYsymgIeiFvY4t3p3Jbg98Rgn6DNLGQUsi6rlhXV0Qxa3AQXN0RrLZkNP
fKs6xpFR6QKNgcKoqCDMwjp1PqI4E8VY53rKmyxJHYOl85u/ESoMLIRFdJDs982N
JxlUUncMx7o9Gj91C6das3AQRM23JJLqTulilVxsuAm+ZIIbQ6Pj2GqKQwZf59L4
3+uwAgcRCzKWaA8OORJ0rR/HlDQVBmqML7zVYBOQponO0eTBei53pKRV+b2L27m+
H+f/HO2QCk43nG4Ly4IyrSbHYorbRGiUGu+eCbGXi4NGF+Hj5ioW/JgVJvr9b/59
1m6TynLe0JaT8tt/SaBBtx8O/TAZdIdU1Z9+rKu1YWaMx4bxZoi06tPyzJWubvLW
cVXJuN9Bypj6iKeH2XUgPdOTY9r9n8pdgpiYEwLx3l6yMPE9cKhSFkAhXYcre9QT
SqewT7bnnClJzg5vNZmutUx/PcdT5ObFoOM3Y/H49HuMKlwSiM0nxdwxamoiLOR2
OJs4re6nRw+vpitESAsjUpn3ZJkl8HNonQxfTX3uJ9M0qN8PlzluSRi5utWOs/gi
RNo5RVIuxuhnVfqIPfGmyCIXn9f9QdDva+ZrTYc0lezI8NY87d5OBUXAgUMtcwTk
M5Dl9jD3BgJd+yPtl7NSEUIlVcTw9uwXAH4w8rhaVpRMb2rcvXaOxg2zLi+/27SG
CQg7NYgfN+pPPjY/OsemamaM7YmGY7k8fzYkOJRkJE2AzNlzbF6k6zki18GOgC82
UxLWqwvBBvojD6H45VNLRHlT2uzwu3ppQe4MUCauoqI+ffYzoCTpFoCyIGnEGfp8
2jZ7Zh7Ntc/H8OigVA19I3guTEmACJ9vS/VB297vVhDbIXLQZ4aeYB56fbAIEFIb
fZ6ijsayRhKRIQ1dCSEGaeN9M3NNZGiSM14Z4ieBDwXnAoAV5ZnbJRqpUTE/JaJ4
Pf3RZ6nUtog4YsOSZCV91Lo6RPbWk71bGeBK8tNU83WESjIj9HIVo/aCCgEsvhgy
PXZW5Nqw5Nm1WWUJp0exEVU+dtiOl8ZQ82drScWO+2lslsnV8oD4p4TJqQeOsn27
tnP3u3HJ31+NECYff6nnZjRAljOEAdyve4JUOBFqL6HWzuLvNH02gXBcZq3BYz6J
mLTJ/kJT79UyG60WMyARS3ly5edPfkdII2juAytRwZsAgYCggN0t4fz2q6Lw4rVJ
m4OJMeN3VHTtLuz0cdJNL1RMGzIjad/l982F2I4PAcMap3mV2srKCfQrlhwJv+sH
Lkn32d5qAkNWFsRzNGFNDtdn+SgtVG0kz5uVj3GiqX3dyZ1UZFo/5MPlQpxLsBKZ
65f9Eb2fCb3HQBJd3KrJqnNQeSIfxPW3M9pGPI6LVpAtopcFu89Nz4B1XsoLTcJa
QtwUp3gFRfDIkho2WiA9IXvJ/i8z6H8pbyYIo36idb0BXLDPVUzEPp9SFGg+t7RZ
Ll3ax/wn9VC3klCscueD2yfcpnFhRj4zY/0geGD7uFj3a4ylGpF7+eVv+FDXFzUJ
adYuYT8LXnyxGdw0hVjZ24cSpjCVnWeSbcoSUSmNlqgU6m8y3eDYi+2OIpq4Lg+4
aYqU8drybh3tz/ib50dBRYCnyrXCnF3BC3Qkl7+yfoJJM97wqTXlNtgWx69Sa24W
UcTuazQfYVvLTGsEmHwgUdC87qJvaztEgxN3BA30xc1DBqMynWFzJcyGtDpwE1AC
O1tptE7IAgRXGtAvuCI8d108TxKEfj9KK2BWAslckHqQc0B0GiKuJAm0Qru0B4o1
PsS3owj10KF4nVbKpVtsH6WxdWuV1Zrc44A1kTUGdmiJrkaLPLEWJnHQW9xZTdz4
86N4e6VqQxYXEzyqmD03UiQUSQpp6HeSlXvc764Wc0Ey9h6yfxE4wcm32oM5EHXZ
GoX6+2txl9gDKVTYicz3taIWyOsUtbCQ8cWQY9/45mzdqlddvKrTvVz5yVc7OD4u
by5fLAxvsvRIKaOuKI67uhK/gjxL8vTA0JK2lZ4SSzTlXqncjFS1oh7DGr0uwZ7V
qFcLqvB55XLyt/Vw10ULEozQvdP7B46KYl60H9eZwm9q87soqum/rmNOsrmvgL/x
7beDbg+ZvfLuUCXZC9Ye81gvHgBajZJHx6s5DV4CwiJPCIBGnZ5C5CuBIn7ELY/m
GHIgfmAd2mV7FbuU4FcCHGKcrJGE+S8wf5bPuX69c+OdZQY8R5zpUqGsbKRJdD8z
J5mxbRYKccRlRXY+oN9yzZ0UrLOXw9lK3F8p1ZczWW9vjHFw+sOz2DVNwR5dL93D
Xy75iQbdxBPTa44KZW2cZLOkE3W7ol4a6vb11+YUylGt8cDZX2BWEqUryzrb5JxN
3+7pdVZ1XSKE5pnbhJEkmFadnXsXVVrSwTAMFxGwybnlyvljF5Mtj5NI7KM+u9ns
PKjINNcHq+L7kPZDQu8fZOwXs7GvR5Y237YWj8JkmcSLAheMd4cm3g60yhIjOSgT
0lELNar1HqLq1f9TGl5HB7vY/bw8sqx70Ungjese0pr2Xh+CbDaQ54tgnzE6goI0
jMfrw66KiuvS4tS17YXlZJoe/Bi67U3hPIBivoml5YDIMqJsqTvFxtctraeKt9OV
6xvOBGaK5r/DcAIqPV67ytheY/AhufjB2OofHPxw2+KwhOaE5oykyPR7buEGMMc0
DOTHFqFsnTXN5kRIpCjA+fQMmJd9pJHpHKMpCz/LvL6zFpg5MckiiSa87+UjHGHc
sDCLiZYHnOdyRvUcPHJPCEcjLvIm0iV6xJHFLtBXQHlbsug02RS5RlFSydcxuenJ
+RlxlzIewVHNr+iJyWneTb6Xbn5flS1785ezGyT1ZH83SUGdr8htTLqg4I2B/tp2
8ElQwBOItQknvCCc8/7VU78Qo0W37PAcpBZJQFddcYrRrSrgcv2RkTbWiqdp52L7
1jyAksSYFbdY62eyqJuSwXMfuXZ2qlu4VqFG64oVdolCojFQPm+DwUWEmELzgBEI
i8x+VQWyETvO+G+kj2VcoD3tQX/d4UwrjvhWrvVILvy7069HNwiSREUujOjIaqav
44K5+jcFHZnWiPCrvYGjEyHKc0NF/Bf+oZhKkf4RSpXz+iiYsnw2gXGXbb9b0SmU
wdrMqGymc0RahocQ7nkAdeuZ7nZNahjSL/mmgtNuWoqnW62X27YGumgHEPnIkcZp
n0MvRTIUSzjLr8+REzMbdCyiR2mAPeMrSHoZHGwLWU24rS42ne9gGZ561o3vtOqx
9Pv62dFP+lwdhPwyv8jgQXCDRanX2JLLIAh8VihoS2NNFlb/Kh9DDe3evIlV9JSj
RXU6w+kXt5I33EUJCyMTPUFW3hyIh1FrUaO5539u1jezXru+kV40JSHrqNnTbTes
ImkhLObt4yvN42nujIjVnFp7EodAgIQC+s8CHfqsnm6EmD81aPpdjGKEHliBJ0fm
/WX6kKzclYCjza4bSGXBk7P81mA50pBoD/LFaS2RP5sPBh4Kt3yvq/OtgzLGZiYY
Z7zob7rMZdl1yIYAyvhMG32Vcoh3nNKKxSMihIR/A28XviX8Eg2ay/TMfa+JVjf5
rSJtFRDJ2qVatHi6KG1Vc3XiEAtxpBHItYs2rBTFDi6wugPVmbbymPT9wFQZkr35
csi9eAh333FHGf2i3a08WMEYT7pdHxe6OjZMpfJm7I1v0vOLoGWc9Eomczz1HhbS
Rj9+gQwHEMbBs/qw1NMseGZcnSp4HfFoYkLLoOoWPQ5riam7blb0hgZWDeLyEuob
7OvSBQyx2vcxwA4g1cBqQi4W+s4iXt0/2kcErA9Ohvz0ym3WUP6v7dvQzoGitVKP
EvtEsOeP4vSYzqdJ/MkbU5syVwqH0690bfsw1835ipn5B0XEQd6om24jEvAl7XjF
RHTdtxO+gnFzUKICYEBuuE+mxpHOzwIT/XgZVn8tCCkR0+USZ9EcDziYW0tEarmj
zadyGff3W2sxigetR6mgpcgp/9TXwXtGrW0Puhb0aEbV8etBERuIEzLYxqZj1rWG
W9DWQx9MWnD4jIwYK6OSOoigxo3RhFnI2KDIxgdJLnaTFbrIcLCW5NLDDO7P0OOO
K/25lNjPtvhNpgrtyhNG3urcf3bjYuNjR7Dh1EJTJqzNArAJduFy2xqOTMAhO98r
NyAvEimpJ91/pSgDZgbL/XzPOgkjfWz01Idub1Zv4bFIuEGbRK+NnqcJNObR6d4/
qQEhuX1hCsFm5QWb9sGdCoII0SZ4BVHCt+k6gwgPw8jPmQpReNYSqmyGgEqoOYhZ
veHh3JxsFQNAN3br8qAHdqCH/fsU0W4XX7u6oQSeVwVyEn51bdOVNZLX1/5JfNJV
TLk6jHJqezsA4GztJBi3UD6vug7AdzvCm73iygbsrGlTb9JyJUdURmRBUuHBfpaY
QwwYMCan1YS9IrDg2xcdWD4Fb0gHY06VfDEmFWZPRhfx7dwNjrKuDjXBEYVMQ5ta
pY1x/l55pdJwkSqlVXnBx0v+AFUhq9YLCzGR4eSfeUxxGr4y7qjhY2/1RrA/9IAl
Oxxuz2ra4OGWGDTJt5zRKnmcD1Qvhq069xd2VD8SgPcxjuPQPwcXEucllHi+78Wl
Krz3xj6LPLjb+/URX1ETr2iYdls7aavdmBwXol4qh3xqkmY4okwcYHS87vaz6JAl
gOZVPYk55rVWg49XtCgXYG4N1U0oJ6AWih3LXDy5X4HUY3ZhrkrqTi+m4i/R1OSF
wrpTNy26M3I3wcPaEgsleUTWUMq/zPrgXeTuS/A04GCNg7MQn1OCGrSKr96jEReK
/szVtuWUvyGS8Tx2a9ndYrsRrDCCbBnunJS0cywVBWbSZGowOcWRhfLsK4zanPtA
aSjVyzk9Gj2y/nhGKhxsgmhm9reLvpyXUrnsWNak7dRn9mnVeZTtaItLaKRCzFtz
XzwWX7O76NFgU4yl8u7wqq78z0VmwaaQNrn1+yoUxzkzmrGisxTZykgQroZYIgtg
dtNRDETcUXJHk2LFRQlagW6DWwaW9SHLjcgCLL4rd2XIhFGRyjuzQ10dafEgDwE0
GhPI/KROa3Lf+0R747F4PVuQmbLU3F0tvQBMVz6xsYf7mO3Gp0NxG4MBkpGVakDn
lMKpmQRyPonscOjia8lii4bU7FDC5YnTK4An2KJyySLosmGpp6r7KZSS9yx2FFd1
gRfc4c+ndUkUqADEdHjPEF9JIWwiUbM0GUM1p8XeZib+bXaaVpOEnjY+XsB4jib9
wp604x9iLl/BFq1JQd0MO3HBn67vU7Ca3LbHV9sfxnSBaRQ6X9H6AjVeQ8nvps82
FcmK8aDZVbsmdbONrbhksaKXSHXqJ1MAkslus1jHWE/sH9Bs/+vgF2Dg7MWEm5Fj
L/kggrKEqtmwjr36kU6PZ8RVce3VRe0h0fC9INzrxHDXiGFFVi4WAk09a/1qa2BS
lkfgs7A+FyJ6PuZILP3UdhdlgmCeegczUizmjJT6tKyNo6V17G0rf3p9t6sA1v2g
FpLgTHIYjgTfGQu+PHQxkC92jdgl4LhDrPJeidRN2fAG8TJI49SOMya6U0ZXapFT
Vrmudjc7g/vVwefLIhXC/HBjtaEdE3GY0GtDUQIUUI2P11SvRbZ51FgDcva6egT+
N4NB2qrj74t8W8zkE7jGIvjwkJPwI25vQY95VTJQzuc2ZRM0/DYunpg78m7cFW1F
/n8s+geKXaWGrYvs1tKtIbZC8mjEkQnJSSvSXT68SrcMU9ab+XtQZMPQrUnw3VnO
+wCpIFuav4nkgDPLBqJHF+t5kaVM74c82bs/GaKnqJNxjefMBqZxoF9KeCJ4+Afw
fMT4cz/BEZZMHV8QMByhcZtxWwldTSuj1lhtzySWildzI41sSVCus9+TgaovLAOr
X+AnSL0iQv6Sk4Hay9uvtf7d4xKV7/wPvLRAPHs1cgGQtb3w0umxc9DfTpTEsv+L
X0FaPakiIiknxmzYshcEI3vFUqfFhSIHA34kllhHYB2rPuS07UcHgJv6x801Qv05
lOWUgt1Kc4yOh3ZCnY5Fzt92PFE9rIBORjr0njE8ZT4lEpFbIbhBryYCwwnCQnDs
/dqRN903wpbLRD6gWObUGzB6sVqwdclQWtyI/T7CAiB/g1Aq6Y0yLWkMwEeItXRq
TjHuiTAJ/vOwWQjD+O9Lp5Pn1/6r6Wm1n+hWTyn4cvkbmBiANBeUd4NxypYy533r
niQH3ma4EoYSxfBsofO/c374TUS7HN+ZQkFJvusQUkIUGRLxR1OW5Zp87MldW+3k
hMk7DYnZEqhYUL+WYUkze6r6FHzjMW3IRnqwfSIvDI84wrG9YKR/vaBVwtyAYn2e
a//jseBFZ31TaSqVFKp4ceKdoHt2bzF5WRU/TzlNoSpZS1zyGBBU+VlVgNZof0CC
Sn61oM6yxJVRiGxtHlzp3CvS8EelGRX02rjc9ABty1uG9KSAMJm14bOyU28xU8Oj
KcjsHp0L35rn0MNNE9dYRNqwM8s9m+va8VWq5TwxY+55IsIDXCY2GZ79hBLF2YMX
9hlQa2FqZtwRI49A+QmlQs4r5kaijWEDzqzwfeYaiF07fLoOMbG48LCJ+IdI7whX
uKplbWsh/fjmvZAKv0Pn5wmjLzPhvHwR1Q+o/J8G3svKO+ELtnn4lrU08nRMM8kr
Ts4ny3s9/g5Rv/6hnAyBvb5DGYm1U3Knhba3r4KdB2v8ECSaZ7z984Ft4bq4eZv2
F+rxnIs33/aTfd7QxjUv8D/JfbtB0oA6z/jnZc9iLQuXolnAERm2ln1yXnoWgOPo
LugOX1e3+n5ieHvYX8ZNeOqzYbw8PCvI9+61KQ5LPIXhOSM89FpcsuM6zDkNvfPX
lnA38SXv7Q8ZgyOTAPF+KjbyFiN9vB7uACLetG2pMci9ktVY8F0AmYEdLHeyMLFe
BuWdOBCN1MNtQgmBB+jfDd8RpQ5gxEh8p5DT/z43FveBOlxk8RAgNHLHcX6aBnwK
rDJxgx6UH6JldDApzN35Hvz/sGeprhP02XmPfzrIZkVRsCkbu0cxdvkzozpbz/JN
mHLOlrYrhawK3x9FPn01Srd4/SnvthysRtHaJCNRVuEsUKG83dHYVHphqwv3p2/c
JTOVolBK7hTDOUgfpyxB0y49mafCJv98SkL82faNU6kkrIhlShQmwyhuWRd1M088
N2UdX3hcwUQ+avbOgrvlFKdLQJmZf87DBAZsOHdHxPbvXa1hwtGRUR+sI4jJTrTS
ZMs9as1Wm/NOC9K16ai3YvnWR37BYQWW5cpkVkjSkM5Mqgc8py1dfkjLFk1IOQtA
oBoUxb9pVpXhWtm2mFSFNHGujA5N0136c62ITl02mGZoldfgkjGXEkxK2eefbhPE
Ka+jOXvfJITkbyR1kXQc0eMQ+M/VNQ2UowItzjG4MaUcfCXv7XHdHR/zbIKQ4TDU
PpHgOZF6RRV5AeZQD1O1BjVaTai7Id7UaSivuQgMhAinF90dW/pjKtXGrAwomARC
m7m9ZlhwJ/zMSozh/FxAxUX7d7BAHH1qNRI5f+BhwMLi484nV/6UYLHaa4jctURt
k3FLe6fpiA5ZMlVXgWYc0NQlAvEi8Hh6EogCbsYIcAXs0E3ReJ6u3qWh7gW6FYeu
x97TkVXg1xNHbrhVTS6oi+PbIf7ie6kIj89yYKC/6cPMP0UvQ+mhKQHMr/wkr46c
MbClLu8eFbTeanYXBFe42tisUNNDb5CE4W6c65iG8J7vbEoF2Xsx6iQfqQXPpcEI
dTbJfdobfGu6xX+Q/znirenxksRGyA7wYavBC63SyNbJHSOcuoETCZtgbVZFx/+1
YFzuPVArd1bW9Isd0s28KUAKwYNLdNGp2k/PX4TbQ45MpZ9PrfU+Gcgyl8+UOY/Y
vh3mTxGQIsZNCJobUcqrvLG42uV58JMh08lLmU4GPBWtETVHx0Aadeic3VrpdGgz
`protect END_PROTECTED