-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
4RG+f48Puq5RcbX20VP7aqDsF29iBCEN0zqGe2rKvyqshZEVNN+EHfXrJtYpRb3U
UlylIeay9C/jM9pDa9BZJIL4PlPMb8tALzgWdSC70FsIIZn1GUU0S3Vjs24jJX7Z
HtUwe5FzgUxrCxjKsECp+czTlLFPatfO9sjC+08SO8lg9EyKGOjO+w==
--pragma protect end_key_block
--pragma protect digest_block
zAq4wBzZPx8QzkDBMkf8mrdUVW4=
--pragma protect end_digest_block
--pragma protect data_block
lRjrnnF8fYLV8+hpqt6J7S4mg2Q5wBBfV67HHwrHthVyZ7HvQC6wlxyKEVPV42ga
GdNUN3itH8RcMPRwX4/Wzje329/pKHJsrWv05GndnUX4y+w36c3JKlx5+68tgZ7m
NvQt3A0nCMWpTkFwGdWk758gxQns4qvMsqp0LZBO0r4/45tqza2n9/mrBDGU7FDn
xsuQw8vPwZ7PU2ZOv/o8W7bP1Q9BRVtyc4bjhEZiytyyLPoO3dX5UmOBo2uo+PFd
oaHcr2zlvzUlkvGa5pXLhCmpYXf1z0T12Zp5shmRA9k/QKRTy7OY5SQBpykXy1wh
1DdnpNs6tDyD7diRXeWNWtavYbgfV102Rctoj/qbMeMoPus87AznVOK4v2qo1enN
cbuMf9TLjULsu9pdtdXWKsVPl8DRsDmWnA+mbjpReypTxZJY2NmX1PHLcRy/01uq
oGVTxQ9hvDF/sGEheZzFMQ8x9UqtgHinXkq8eks982ToAQVTsc76g9HMmTb7DjmU
EmGNFwgaTmXSxd26TdKO4tW3OHzDDWMJQOmZ+rADz6TPAV4efKb+ZUbvnIq3S71u
q/90OVBFthaJwM+zW2iy+/Bobs/uzYlufh4y55onUJOVGXBBP3VFU4S8H43wVsKj
GsBB4w1efBjMF9QYycCfZVrmjQF2OJcPB2lPDWIVE7S8Xg57imseQNVxGqpUSok5
8QEZWId47qKb3jubV2jwg3hg6qcQqtmrJKiXj+AMm2Hv9mYRqQHJyv0e9MTWhPzW
1aCF0WzjPO+dPVf85grgevQhfotwTSBvM17K3XDoaJW7WAjJAGCU5pgbz+8ESSKU
pX469r/u2V1YZt+3D5RCbCzLpUXi5MCmpmVOXo+aSLJWeetQqKi9NFUa/q12zsXG
0TDTpLVQmgR3+LeUu2kEkvw0bAGBXEunc+mq83RQf7GvrVHB7OyJSlOW1mM2pxJp
+w0FO/ErTmBvsl4IKcUYK/QUB6w/Torpy70fjZQpYj+uN48DEl5/UaeUg0+qJnsM
ivh/Q2jpW8AH00zYHULOa++66ZArt+x7FV4c+Izj2GM+dLz91/uekez+q1Lptvgs
QCyK6i8Kx1M0rkHqJOgIYAJ/MYCX/cYh+5jXK/MAdsFixzjTBZjsG6EQ71xGwDsH
WE1mh53WWrtcJ4nsvp5A8+qafCPOgdg+ndov/+heXHYmaJVViXHoAyu6qakl3GHa
c/rTiKDt22OwkpXGyY53LgTQqAZvZJQSFNTnsRIK57VTalJlV1+cUvTZADMw10QG
hYlemXVSFA0qOJ/sOaOnkKR+Srb7hVSEMDeDuj9RoCWHk9Lna1KaAE11VcGRYXoO
Q5aWUXxFG3GvKistTIDxsPFxdWyVQTdkGgJWctcltofbjIkgndyeGn8kvPtbFHm9
vOgWglQOWcy5Yu5lYRMycPu3bYIKPJRY5tZfVi6XKvjY653PcWJ2ppfuSGPBXG0i
WOsYHaQvyIl68c9NOcaaRtjCHx5aDoC9WNcSSF/eVYoOrf4nNXONNPlIBDVFKUGR
5y338zi8u7ZEFgtqq7I4+ChqehEyeUs4+HfrDfNdHbbmvOivE3PpjqyVmfi91bRv
lAubJpxH08mnCTr2owRLVz899ql/vhdKg1Tnhpe3c3KMJJ3jinJdS3Y34FBHuu5S
exiiO3QFbF3HrruHBtVnI0UGIuPeV91qHonC2WpyofQASVAeFRDiOXhNukNElwGg
uGwc2Se9nCV0U5ivjBUhV96Sj0JHHT+8Ovd7akojf3DmCHYnjOIQDFLSEy3XrMkj
zqiJQqckhhMK/t+PSyya/mwTAyqHqcgb1wFfSBAQzLEKPiWiIygflc9TbP+Cmzdj
hLtqeRs+3aHZXScydwYYuuBVshZYG4s2A+KkexI/+CdavZAvyEu+zfBXbspkG70i
NA4hlZSj8gZZiEcaYJ+uUxXf6MekNun+ANx0wqtk8glMIMasTTLekrnqzRrki153
y0AEUjY7tBZ+FAZggtwXQyTOl/gsGy9ZUA/btElGjxFTEzYgMM17H5V/QAQEds9o
lJg3PGMzVzLCBu0oImBM759l/s56//H1+q0NH4+LXaePTAbsW4xO7rRHjX7g+Z0H
SC8YRROkcW8KjtP7zvK38yVS3Hv5QqQgp1jTgrjHAi37DL3/o63YTtT9wLGkS2Lr
Q/gfLPrMK6s+GTElydOIM4Lq8tm9uPtrXQSsTQtVGu8N592+aFPB0tR1bOpxihf7
di5LQbQjwmf+BZF8S39ATKHab5av3SwKPIlsnO6gweTds7ibvSn6oAW4i/Hm1Tm/
GHxVFl5RUupAGA7JmAa8A7R17CxpR9TmrE+Q88ykHJNmqKwUDLSOUf7qEpThENsp
LaV0t1T0cDJ9PrOMntU14/v9ordgWTXj0KFYXxHSYhFnIhFxDRpoJo24PIguuIuD
1lnOtRUmlshWVtnf/2pic2glEpiR0fWaIjISlYNTfE+PW65QB6fLKqzqbHDY5Pib
zRqBkrcmhkfUkMY5A7m50WAZM7YykYueM2ZQyoSrh4FRawEdsL1BJ/UR+DOJmhj+
xBabKPkUveT8I0AoY1fXbKIGsaD5FRtG2zHpC60igzqsq1Wl2LceaIjYdIGJdzO1
FJtX9cZlgtYFEYc7hwc2R92k1ufshsQusSTj2zMdXHZzBg+xLsDWFChHDxnV7/Sv
XFHvaK7zZFwQKSuTt+8om+FU/mRnhK1kXdMd5BR9v5RYvGqTt9kYdDhw/WVyQm0A
LIUW+bhImU6PpZzA98roq9nKFAAqPc9b0aKN9DV2ri1Hq0zjOmJXY2IjmrfD6h7x
QWzSpKAJMH1ic8B8uNFQTsA7xT/JAP3HWKzKpd/EoPzn99sb5NgqNaABMJYiX7Zh
lwaOhOz/61AsRcd+StsbGW1rOXCiU4GuzpD8XmjVcXs0zst25l0MveYEdguhYvp8
pun80KI9j2SMdsaCA7HsJTYDMIt7g/CPjLQUCbw3R0Bq2dHVSsYpG7D4bESGhc7a
bTLCG8W/qnKogF/77QUVUxDRqf8+GgG3TcZTEdGniYakXxzMJZ3mLZOkAGF7qHGY
3AoLyCXK2D/uXqa+DPwPYCj2Td+eYHp8FP0ejKECgaMgLvF+UigQcJ4LyfklonYm
qDpANBnS0XChRQu6nkL772dufh9sOg7vbp7cwZ2ml1KzCBXNSOKZ2GLnlsq2TkTV
p5Csq7vSuzMwTmuN8dLQTRgys+eEnm/uQ2p6drSN721Uprls2hce+3eeaOtcHTTg
34ZNPHw73WHfYJlTD3i5dkAQB9K30cl/B79HaooLrWGibWaLolYRREj5s71u3vSC
5sJaENBkcyA5CEMlam3dH2sOr6p1maMKL0p2nY3aaQRl0do/0D3vEf2h1f2dDEY/
U6GayGxpTN7lNfnzPsD/sqIy4GitlUH+T+Llwxurxtv7cxmJ3HOOlb+QwmqrIrDx
6bk4TVugJlulsz4V9Poi5TJxzWJ3LrNB9N6Bg3NF4WrOV2/2ZZ/gEP5kRLS/e0bx
j5raF0SvQfq1zuMSLdMmorMClfFf43gJIrStX/UDbNGAIuiQtSfLxI+SKZHXusDE
TEdPMvMkxb8juipy6E0ewi24i4+L6XXQtyuJWBH9wa8+S6a8f5+xS9YWR7V9yKHY
bNcx/Oa8t0WQQoLa6Fh33oLmMTW1c+2aefZAeusCkZQ62/hMdJEIC370sQfOIjWL
AJwfU/T6B1g+rZaYbde+/KiGNc7h65Ag81vJf5FE/GmgXEVCJ512EqYBDwXOosyN
N1GFTD8pFu71U5By5rPlfBurWQsLf2ZBNKCAbsLtIHqqZBQbAQC9ekmMXnKFOOC8
fzY8WEgAQxX50gYfi9Zdvdkpm8Sg4nKPer5BdP2+/PzkM5HWIYQsD/sCWgUh1Wjw
ML69AScYCbkuyLdQdh673Wn2XjZ3vHUVZm4z/3PlW8jkCERoMrA4e3CslgykbrW3
pZTDKaou2ixqzVKKJZL7JEN5MQVN0fzb0jJwnok/Mtj8XoGzW1cLj1w8TbtOLAzz
O63XPmcMp8tHltrG6hivxaGIOYay5lBFmKkjDWYeWV7gWqLGKvM2j9Hv+Zk0qqa9
3Y4aRrSDtyeivSpPt981pI1Au33peNFnnTl+euzNunu+dyXxZW0e7rePuyX8viZW
JCfdKSwoj0dhMexdq1ils0vLp5VEpF/xZLEBsJ400GScOaK1r8YDc07DcIwpseM5
gYgFDzKOevPb/y6gkyx6RNaYNsSrQ8w0xcKXX3SZZzfhiboP4q6Ajrb0c0XBJ/24
HohkJi2oYsOqTHF+PKf3V/wFLjOqWu9S5g6n395BTq8BKhgd6eYr6gwtIX1ap8+t
8F94ZrcWhao8OmBRrNFwiKKxgARmD7W6liGUfc8OFelmL9Ds8LNEKPaOFuSJ9N5M
FfhveETXbYsEjx8z/ISvfVYpOczy5BrWjn+zSqRalIU03kB+pRUJtYgnIhYfjOBG
4aGVYh781S47HZc1T4NaCTf/9ahXCLHYspJ+WFv69CMBNn+K7aNEjinXbyghc1Uq
0meSEUqa9BBzewlSq62EyXyVzlQRJTH3gyhB5utRZESjl1rmowFPB5ofcX66J57q
UPytxtdXODyzo/RqlMxLg6UUYWOhxNKnjVMwxDIZ+H0BHBNUFDXyCcBZ3ToP11x/
v2D4CHWB6pl/rJjSvsu2HhU/CUh2VtTtIN4CW8oP2raCUuUhpV+7nNVt0shmCwlY
QJkfCMlq42zjiJgyjGxaY8O1ljUdS6q5/3flFbkqhZQabSUhJrTUc/slESechbfi
zDawv5B0npXGOrajGF6cKaosRzyLP3jzoIobJGD+b/VHRBBCQdZKghjzzVoWcLrn
Bywvg74rcQgIUaIh/W47cPbDLH3kIFdm063WyB1oThK9RCEgDF7x4mKl2FI0VFKa
Nd/KBQHcG36SrliFqBqBT3ViaVGJA5zvD94XthTh5iL1YTk4cV3N32LbZSZ8MgsO
/WV3Uvl/muePdQvxTDkXRi7W6v6X+YfC20QpTP59T7xiNQILynBa8zRnanb42ndi
CI4jD+n0g3/f9DfR0I1U5XI36uRlxNHjMXVj7GSOsa9Ti5fZ3G7iIZlk6s9b78qb
FlM2jhoOlGsp60i3+kk4iDuLMRCFY1QrnvFizzO5rcSvGp3Uu+xkhyNeg2li3ERd
/uqTCbiBUhdkW5L4RFcPzvUNpGmLP0xpKUV6sBoTf7xTCg8H2Uy/ZQ84hw+ouZwW
Z3DGJSMCToYk4b21Q3/RWMpDfzCI70F0V9QkzL84xJJKJ27Pt9mlmaUIFtgDcEHQ
XeiyGFpUJb4quwneqWsGkDeOIQN6AmzdPxxT7gVPy4tS+O9yT30cOdhT4isoo9AL
CVxmxJzIG/3loJOH+rUxz5e02ASjcwWn+xGNPxjRzPxRBPpmRvofi5+byyfU+K6P
llLtBd3HZt21ZKnJVFaB0SKavgJ7o5kjcr1S+ighRobN2OGn0xlR3Wat6jntD9GF
hhrq5iAzA+hT0ZiQFcUDNJGL8S27oK4F4qLN7ibzasi0AzSnvmUlXfYy/7Ro7503
RusK9eSlnuid/RGP6UGLSnt8vSOtYyU3ePkZcAYfRpuWtc8zYollBM7P2z+h5X06
pO/2NP1NSj5nPYohZhKaD2I647yCrExvRFS3qmi5PSM3vtXHAXZW0ISJuubNS+Z4
1HN+XSp9s5wDw/esrMO2X0RiDPhIo11XqlhN/xoW2n0c7kcyGVDqjqEmsnP4lHGW
GZsfHcqlL1QTQcw7ruqk5ohYqh0r9nbfwEx+Zi2dq/+LZXGyhr9j5BUtNEitv5Eq
GnfNfFsOzo0kKGyqbSGf5B4yc/rjByMC13tUN1L5tEduDCFwmuTngNdlPSSy+48z
Gzt6XhYdXHbl8btTyvsI3FL15POF5X+44SvYwxx6JwZoXZ8fgcXUUuuyLSVkM1Qs
Ep/OZztXmHaCbmWZExqqgUIk19QprI1sEf2tvUBuRfVWMiMXca4l/UR4EQykPuQl
xhqyFZIXd+CrOPIQUGK8V2H3RrDd5D3IwGWYUo6zcKJEQoOKXjFHyI+JyCAJD3E7
z5YodeZrRSeDLw4CIXhRAN7dujC+n3/Ejkx3OdHEvLoicjlOZqtJY+YQ+NNaPntR
lMb20R6kGrbYNKMMGWu10vGDb5o+FS03ce0IHKUJ79TFBjjbk5Ia+eO5m/sycnS+
TvkN/qwfDCXBxmCq0gBtn1i3dSi0et6XiPb4sS54RPOWd/+iYoiUQiSp1vErJMb3
V48W+9iyCooqgtJ1+rL4fYLKnZe/V6TeVSefq0KJP5rE3pPybw4kN2raAAlfeodz
lXpDnaQXgObGs2OzE0sml2gKSgTqd7lsqtYC1iBFxD6Fgb10gnbTniFGcysQwga5
x0M8rMAL4a1lA2XtSq5ydp5MXcqWzrKkJftrczGPhgfUFZdtgX+MPVhbGbdGwpUt
m/WXd3kxQ9mCAI9KOGh8HiXI51WOlZQBH1AlOmwkoZKQXvFq2vzQFbfBbnG6QpTk
XhkRKIFp1QADdzryh4qJ10voVb3+1i1lwKLkSdMGa1feQKD9udrF6dUoKIAsP6O5
TvwzrTtuTWdLOR4WK/cTLFVCmvjiekpG2Jkjxjf7mUxSCWDwyIswEqntOTOgrM+L
b72PHvjiLjMuBHxXX2ucdrPtmV2RovXv8Rwk3jwNh1oH7k5tBC9Cdq+5V9Iep4Qz
XqQlTrFZr6tSdUQGNWfgD8+aBwkdH6aQdSY+EsjJM/snKsiz98ZcqZ7ibyBR7+yx
OxwGFszRI8erJvbKgTFXSYt45PaF5kACgMeaGkGtw0n0krm1hi9/TPKWoeB4lgjI
Qvxx9HkhFfRsW87SyuoTAXjRqz6Zx3CL/ccp7+kXXaVBcMgpWN4NTG427hb4jZcI
w3/4xxksUEeCfQXZd64zDI81WQdPQlJcJsUfmLzrTjEtTSN/yAajDtRVslHZ9tHR
6zIWjx7Yx/Lt2/erlPgqa9ZSG0dYN1SFK5NABvIg7ucFrXB8RYJ+cs2pGMqjylvC
g+aUgYX5j44dgtqAMnFBwK2MmStq+itDfXWWKgFHMZga74G2SLcaQXmIvU/3RXBY
bbSMuPYwIl5g2uzWlooes63ReMcpYtBwNimaze0YW6w6YX0wMxO8lhUY5M/byZcZ
qtQeqH1PZkCsiHMkM4BvFEOVfYCm9t4YCXEw4+No2r34anSqT0hFl4HDQrjPwzmd
ffeeY09C5pROELhEAhd3TXv1rzOol465ZOEStXA3PHoZGVkoIB7OuNMjojf5+RUm
kQXgcjUYT8LtdRePPaB86nIB9ONZvNEgxEaflM+dYhrz3FUfQwXd5E42kRTT2gRh
nHu53AIEwJlI2L7QXs1AyOK6bm4T96sSnW/YR9/iL7PjU9GbBgJ6NdBGZL5yrbks
/RSrBlCP4VhGlZXCaKxtZ1dKseYLysjQcsbHM7GhNeePkfFSOZuLNjMUJrQmpSOi
0abSSf9ujId/30qcF72zh9m6VlCW9ksRZb0/Mkh4X2pqzsSUxLYrRw/bN2XjdbnP
k79lu6B0rUG/ogF/PXbaNYHgQPp6x0y3PFM9c2U3se7ObO8QCpk25sUEoSvb490v
N3CwJC2ONUI3uzL1gbUoO7umc7NtqNhv6Uiylg7gmBpIRxuKKGg4i6lgzID0Vpb7
JCLKqraJGIoUY8Ygk28K2/Fo0VcqZNTH1CKGu18V5ixwEB2M6Vr/w/yxt6IyW/pn
gQS82AYbD9wLPGv+EqVkJtj5FUKZtim84K5+HpjIZXREHp1BdfeT6PuXTyO3wN/f
DV+cV9/ZGtdKxO8irYHwoSoavssB0X0Th0Q+1npKOlMVPIjrqVgpc8j5LGYCuTxt
oElRKBwGc2Y8RaRaoGP/GVtT26ahUoFCGWQVWvTijQtJY4YzdQPrD2sGZkZuArMZ
1z71e39a/gLbuJ6MjrUUFAp/ROmEwM3C/fdmD3kc+vMm74OfO/BebBcA5nvlHOUp
/vDlHCVZHG3T4CtiDQ1sZ6v7Fi1NTsSu68kP/B1esKkHS1UhwvNAN265vDRS8tA8
qH9gSF1ZCXcfEqmXQNqTnxYS7E7cNHv5XM7yLPpBu50gF9FuXcg7tigx/P67xhNf
aK8pO5IGI2X5Q2R2B7eGuegYQdBvxQqaEd4XffJn9XWBb0dThBUxrP5AVZDKqclp
c/u2rD6ht/PnXq+Br7lm9xhZM1oIzI7GQ3SeoaEPlwIqph/eaj1ouY6ttBI+rSB0
lqukjCUKmhM1ToeuJw7Aq7qfhgb9L4hfIQnaWb7e5Q2RgrwahttAoQOtrvEX9vGY
+6p0kukq5U/xtE/Lid1FCdMdFNVyJm4oHBUE1E2uYGjLhcZzY/4Fl5rVW4bfHtn0
jrBQjVRdS1975COIlv0f+p2dkWRPzSMDdglHNRujsYw9di387930WqJLhkuli6UC
pW5jXXJILFlGL0jUXIwS9r7zZ3aLvsvqJ1NY4+Farm2ipMqy5o3golIzqNJHq2Iu
cKC51cFEZ0iKInOnz582gDS9Hal/VhCGC6De+jqCZccDx+8/Jp706VVLALF9kJaD
FgpW+gQT+5pUVFYuzK7qcRtfq7AnlqoBURECjMaoZgcUb/m4bP9x3raMeigajICR
M2P6TNqw68CZX06/XUml+Z4AZLVw99Fh4BLYDnAvj+1Bif6oZcAYX+8tEZLvyKYX
SWUQN7xeYvJbDGfoU1tO/AWSfo53R4EDETZhT9/M+d0ReQrHotO3WlUY5XvLBPI8
JP+zQhhVzrZOdQ8rSZMA2XoEZ/B+RvXkU5S7FGk8MJ+l9dQGFi+SmXo5n3FRCdPt
16Gz/OntX7YD84Mkt+Tiu5SMnwCT1yULPLUOO3/6Sas9RJk4xg1A1GykN5gouR0k
WacMDVUVlNxxyPnG9mjCcMhb9hQ9Ym3Q00GwbOyw5e/NtqDKVgW+eOTijDQwIUbm
uu03pTyzm1i5+DlVDWKTbooQ3SEHKduTq5yqMu4zEgjAJJw7RkLEybV4PkDcg/i0
Gl384nfFuxyZ6hhAtALzxot0Iw7XW9N5kU2MefIpgkazkHtYfi/uO9ZvYmm3n+jH
JFFdL5OIEC7DXVnh8QdNXPsLLIVs8KAxm6xnmhtqyOhAfYGKwhrxKm4NRyQsbqlq
t42YD5Er9I/LPcdcHwN7BAaChw/IDhrbN5AGTGmR/+GlT3C+sBkEJ7d+cAvWnaKV
BbjEmRY3wz+RLk4XRUP++9Gre8DvFDYSwPzX98sdtZMOvs3h0qTRrKgSsqlE84TL
boFkddDxJFuqHve3vy8sPUbIR/lTCnUQMZEAbZhcAGrKDh3VsocM7MH0QMoBQC0i
ezGoVrwUyoGdCi+aGW4WmdJ2YnOqmKQGyYlRR+4iMKPBMsU8Nc7KYj5H4aJ4Qlf3
6jjILGkeUHyN6Pkp9b3uSVSy4uiRg5Zd3cyqUDdCaE2Z2GzOHKtYttjNtdth/qsf
LWYmy2YEjYE8vaOQIg2OZ8ZKvU7U1XOcasIdvtMsGu3ZihAPiFGFIf/2u7+5tI6S
tSzDrHbi1HCbTFpNM4dSeiQpVgkdaearFXx8KInAA317cZPv2Is4dYYtbENpCNh/
MTOM3woZOrly/RFdjSsdjQGrdSEnwj+/uVQoIeyTSYVWxNkWkoefN4TqSASjddlj
rUij+UOoOUaYnQOLp04IKUNZ+fl9yGj+eGzejQS92zYz5vAhWBlCHW4bejiI0H9s
QdQMwNT5k3+DM2NZZIGgT3RYDZ32dST+POSiW9+7sjVOw0xXxmtbptvOROOIdQA8
/ePU7NMJbHEgY1CY/leS4HEdV1cvjOjQC47SHdpXVpMq5gOiGzQSiO07UgkxyvLK
fV5kDA6M6Y6bAHMFZZDfZfOmUfJmMJ2M0DtuL6/yIbOPLj3GZhyfgZv7RbiV/MFO
dHt/uNv+5j+kAnx8fDMgjle8KPQQ5A3Vebi/At+kdafsCeWz58DNMcACR9qp0VHj
mAdDMJrAzhyDxsO+HQBBQU2IXZ/GhvlijTwt3HeTzbqiJ84VWCmvEFemYI1qzz48
RArHzAN+N3q01LOGKpRYUvy0UaYKeAM+2+8VJa9yNJBronhm3WAltrTCw0/koa08
sLxnzLlPfVySPyjf2EFUKF0i0swgWF5Weuv4YKHf8l0PYADhA6te4h/fPt9saH42
t4zaw+NZbgIUHFx6Bdo8IanV8wisvpML+4eKqeiPgjDFPokspBkMLi8nU2F5gmO9
0KfCSDR4gJK7iCNgqCqpkC3dDt0WeHjC38TyYjuEFCusKIvThGVceZkhwUYTjDtP
ahw84vFkXq1Zzzfx+DZa0TCbvw23hZW/u34x9M9GKbabr6Wi4eOhE+V4C6J2WNED
yS8zz7a3ybCAJB506tMFzHVgNC+1biGW4GBvlbpx/N5SFNkFYbrE1llNVFA2W8C5
ZtLELpfK0dgnZvgxyLxpDLyIxZrsUA9ethpuRbMqtsEAF97ydD6TPzUeRuwLGTFp
uG3e5u4b6JMnZztKjtcjKgYySIPBtl1RU5MvB7/l7FNEOud4gBQD7RH3hDioo2eg
4hkmluCj/sH3+9ba4oZuRbcmbCVlM5dvgzk+qJD0PvMUJ2fz/O61Q88TuR/Eup8w
HJoMOoqMjV2vt2agVBe7OY2YUkoDdpGhlCTtqoz/7+QezaVv1RgaHhSYUswAFX9V
T3lNV62gAgJIArAx+jnlLsIdzipiY7S2uSsYwl2OOL6NKPdBusW5nH3QG7sqxImu
WoUNGgrHVIw/fvWupUA6HLNk/gDItC9z1vaAYhbRzqdLl8BplBse9MehTd6XmdNq
6dh/Eef6gckeLDfZeQXUoyr1TQsNRmWzl8KIapTcaTcqlsvmhiTlwYBJGl2PXSIr
Azi/yEY9IbGUgTXXCYjQ0Ym8+eXHyH4io0rh5WYEKho1clGacLvHYFAKWWWAvQU7
cMnBsLPgl5/1g/XSF9xdkwHtIB2oDklXX2yohR+APIMuSRGqcqPmU6LB4E9G9dZ/
zJ07+Hjc0S0Bm69XIdZDUxwSTLI74CqWht2qTG9u9NP86rp/O8C8/ck+t/nrriiA
wlZbokB1o1nftnEvdC4kCQshrKwpAydNfkOBa7N9mWI1t0LKQt2ayM5Ldm3tZnrb
WK71sGyTy5PMpB3YAuX7J1rupndIF7+wj5f9ylL4gCWTitS1rx8JyC4/teuiUWOj
AU0oKQ63ijgyLDNNLCzL4K/sxH+6O9MjhANclYauMpJH8JGOv78bOM69FOzB8x2g
UhFXweU/IS8unoAbeM5IEDSCr6T4gi+FnHVG2hq2Nb5K1EvCOnKvh+W8h+itOeqe
7SVmtQtHsGl17WerjCv+TYlFGJWUnt/kmrORg9rWFTXHJ8R3+1XtN7YH3zBgf72h
xjnxh5IwLu55iloCEZGGQqJSndnzC/BapF+OcT4ZBAblYAmFymrbQgX2Oznd2tAH
JdH3T3IMeeYLZbCeb0cR5nngEuGoyhwc44eRaIqnzcPmTqV6vmwH9ePPsT+nENrt
MckGNMSWYZx2rP8EWe3PAXbfEsv/lu3Kc8Ic3qeRuW2x7W0kO9GqDMLj6Pots2Pc
v2Z0/oKqSnMAOo0poNdbd3nH15DR2Majt7+5ETo0UIaTP/+F2fLr8W0Lm62N5zCY
clNmV6lHkogj4UYoJn7qG/ZQqMnRE1RdVZhqzYC5YCzVveESyDphl9Gqr9z3w6CT
P4kk589vurPWoT7tncT3SJzu62hSx6AjqNZWNvEHVfXkNH6IvByg6kRq4vYW2ojF
5qCahHATRjDIHO2w4LxwSCbgQKStzzj3SdEEs8/qoUqkpuJ7MwzqVXebKv2WxDiN
K5T1UGr2qYBXO6wLj0kc9xbMgfymbeLb0tFRu5nt1JHw12oUsYvnSSsv5/6Scd/a
u/3Y3+MTWluCrS1Gfwo4H2bKRetJlwKD5stLCtflgprib/BWAUyuRQP7KD5bC34G
lKajvcAhs7gZq42QMawl57gy4ZFlmPb1rrwH+cZdKAViQN/mY0W+MbxcxX4IbT5+
FCtfCZ4LgSEqxzgwrRXJdAWaVn0uLYo6bio2E/UOS16UXpiGRaw2m8id8pp2C3N0
gHJvWz04aQ+m12ntYRG58Nb2rpMOzv3OP9XgzAyuauWImXaQYrIXb7GjpfTajt11
yPDIbJrH4jdfAynYDbr5hjbq9ppjbgtIBm6InoN/Boh7km7cgLP+iKNH+u+kzhRY
nggMyKOn6imQbfisWGgVsuSnGeZgW3MKhMZBpLD67wf+iHSj3WSLrL9rF5YNSEzG
fQYPrhYRq+F62ypAYt4Q3S3XtSYEoGjNJcR5Uy4n0IrbsYQnMSo+2Ys03Tm2xGEN
HwuMtb1yGJF17VxeYwdElaZZ1XKJOoIDIflpLmZgqQ4DuRGwWvgMiEbhqUarMRUg
kAgm8gA+pDWAxufuDMAVnwBtvnjruHNnwnkS5l3VKehx8a9Kl4gisOij51NN5Tc4
47SlBYRqwCy5eUWOmUF7Sk+gPYyRpSHjFpsOEIYq39Z/W4rBkQHGmokZ0IH1OfEE
YH9Q1HnllV7vX4UeriN5tATUIW+J5LMKi1qEvbQXSh9BKb9NSAbgFFLdWVNk9/YY
xVPyfQIDPARYannGZZVIZeuzKR8T+S1xja5izz7QHM9T0EE1rYtnN+y3wDHC0VBH
kGqGt/UCAmfPcKcFiLtSwUlZOfQWkZb2gNa1vrdLjUQSNr+9u7U4jX2ft3ZOjoXT
fDxv6dEjuwqYYDvfjVIK1NikqFbpIUP9qjnSw8UFUduCjpwXt152av+e7NHscRu9
ru4MsDDD4WrnLKRUbyGuEDZ6hDaearqsGK2sX4xLMCHIq1mnyt44b8cOGlL+b/6f
16xrVLcbVqIoB6GiFAsHGK7LSVXkmS//CMwxByMytovsgNXZsOPmVE/XKpkPIkvX
JpGayavk5s5MztuM2CQmgM50yEUhqSegPkd7j2iaT7jkf3Aoty5yix9FqkisY0/i
RuZWmbKUy2rK7g0IzgRmS4aavXJCTVicSO0AGimfS7OGuXuMk7dmqusZ0MrTwbyd
MCtuCm60ylMex8VVj7eVo+wP5c29UzZMtIZ6poexSOCIFpU6JcRsQ4NpaMjK5Kfw
J8TIvKCISn/r3fbM7LTKViGuHGQn1ZJQ1derqaZQ8/rXQkRe5dnRB8DvWAVJ3wre
r8Sa4gw9Pe5AEVEEpgN7Ubf135Ex+txX2LOKtSvs04fQqA9Qb1y/2zAnvlw4xQKz
R0Pb28BwR6GUY6XPTFe2cqLJfE+T+9660BV/lzvvW4xCoM8z1wZ0CcfYSvMvPNfn
3ZW8On1d8H0syfeWEvQg73DYK/5kgsLU5E+9B8KGLFTr9bihozOOchA85YRNNH7j
Kc3XGRkJvmcAST1Ymua82GtY0aJM9VRbOjn18DBPrezG/O/uh3ocf5AL2f/qkK6Q
+1BNCcK16aydZcCPH3kMn2ocWWwhjxSMgfLRhFfOyF4VVvVaoHgBsjXdiDY3Eo5G
ytIJpp8kJhJ9Ot/PoMpO8LQKFXkODkZvDfLiJmV71xOms9cMz8xFP/PZ9tS/cV6T
GMcAN+iNEGZlfa3Qe3WQNq0LtAWQarzX66q35DzmVEHYE+jjVrWsB8JTvcwVtCcl
yUMC7fOZ7VDED9HLebucxRY4KfgQnx0P4zZ9IEYkS9CWn64VVL8s1Hn0kvUiey4a
yWZTD8xBCnvU9XbH17/aEhOhuaxqCPeemOeGWUNuaEOuZELbQb9CXZcNiNE5egVm
ZfsHgUVPnD4hDOwL3SsmL9N8iGT7ZCvAumHWclC7cs3w+2zusZIOWiX5mHnG89iu
LbRCEb8v7hDiHqE1AKe0Q+1PlgMBMkg82qSFeQM3N/AsOO53198iiTGVngXsD5ha
xbVBFQH8UBi3Ievcy9/Uzp3jc5ZAZ2qaKvhZeywexglYPmQCabHgfNWG2qMGxwqc
F8gzFRti5GlwAdeQ1R21bTWl/rAvzTyLQj6bSPoHqADH7S4GyGF6TImvCmZvumJg
mh4XuLnymfcoVhPAerRmVULf9qxy2e9b5gMIjN0IilkSbr+uHMuaYFlmwxDlVuGl
Ee9hae+DIlpZDHn7vppt+1wzUZ+0gcRVylmdf73HnVu0bhDKJtaqX7Rg0UKDMaA6
22OUjCR06U04HE3MX0MPjGJW+3ENhxgXMBymMRGSa4VSrs8MHc2RbC3jpOYGCXJ8
0R7CD4JJCMsIPSE+aZ2XNmyhmUx6VWTBy7PrpjFKRM1lpKpFfd1zh29mY02tPIYt
71fwarZg4Itz+JnHK/d+KsrXFHi4kdThVO8Dj55ebF26JZtJCfOVpDaxxcN7wAZ0
TxD/TUSJYZmC2FvDiRimtIlI8gvnN7Rau8toSC6GQHvADyStU7HyvLrAwQZkAnf0
rE3sTZRHiXMKThiiuMsCbLOXIBjBhppmVTL3666vy2BI6Z1a8T0g+jS91q9kAhCL
vDhWtXLQezJzl3HIT6ThShwl7KW6sPr212zAqXimXUiRCJcMNnnLTVwmbFWpyCVJ
9yCNeK5qBbwFZXpNKBPFlRhFO/Nju8dSkrxvNK20XoqRFOIm0huKX0R8eqWqGZ8t
5UhhZBoNodQs00NEQwHE0JxInl6oY9TGWyq+uixdJ1ETDRKygtep0uhQJzxXNaoq
WnVko8RWQ3+iYjiagHh+a7n3nNsn2tNT7dtw8wWXBAZHtCM3jx1b007Ib0i2X3We
sYEA+BSWyhXhXR9mmZQWMpYpi0cF5Pc2Autgr1J5EGgo4QAS0r3grV3EQSHOfOgQ
Jm0+pVwzgAe0eQu+0r2kXRldZXPydfuJkmh4zlCgK7KX7cRFj6cxakiT2tosb50R
eD4+US9xMDMZxAM5WujyTLwWRkUqkuysbVVhGtdXbL2Ly/JasA4n8dDqGzH9hRpF
YSDzVxo9syLtR/SN8DSGZvcsbpWysbQuJZxD9yCsX+ZWo+G7pYBvQ8IGmWYNbu+J
Z0oYNA2CpCqxHIFrDpFpjyFSfkAD6F9sA8y5re7hTLOfABX41d5gFrb4BlsHJCSa
IqOcWod/L4BcusUDPVqUzaivHcHVRDfbX/RVDd+e8Kb+9HVfdZTP4xh8X2C4t42n
PlcFD+9aPMNsRhysBm6/1FwQ1O/VV7Bq/Jc3OwG7QL6A8pr2zub1PVgvmyWP02My
Zf8herCIr8dnoZFi17J/VVYcS9iOqE2fWn/TKB62YsVius6GY+rWnUUo4igX44qR
QBplZCTWSP3yAfKAlt9tKZb8/Bv9Amse37qWXahcjmebX62wFmCk2Fe+Uk07u2mo
8rkBexg2XfPbI80zWxScBbC1p2dsIzcHTHXcJejezVgCIDcYapqVWq7H1NtdG2zc
zMoBuyKDmIVvw84TW/SCnUgG/Rzw1NKmd3cizhTRXbuHl+Wy4LkhdsNnKHAOe206
TseqsfoFD3ikWmqhhxF/INOreKDN9pGrKIWM9NWhXv4CVi3YicdEomVOH1qeiTot
1ia1LataX+l1XnRQbguOwWeBY9y/lpcbPFie5Jyo/CoOrAAkixesIQcZOiHUlY1Y
+1QL4t/JvFImgg6WekBaTLnY1U8oGnKrPcQKi2BSxTebemKKXK6pnAuVWujeJsh2
GZSOJcyXfkwOMBD4t9omm1TlR+ajXG9RkqkyKSgm/liJW8o91Lryv5xsEIPJoOu8
CiUHDwbs8jeQfyvBgfMoP2vKptArNC7k7Qi0sU3XYCI1rDDoHUWdOlQ8Tt8X/4sB
e4n3Xw4VuMdcaItQlVcHXxKK6PPusGVcMLEeqMd+9el+mWTg4Cw2OZnyxIMoN3KB
oS5BUaXBEQyuWPIY+vmsGO4T4u1zv8GfhWyaMvEgKDz7gKBlPuH/7g/TcEmwPgUY
UCmqfpnSebukfOvztNDcK5UBRXwvwAkGWLHTn84ds3/vijryQmD8bAVEddy/B3AT
Qf2YVuZV7JaBl1fZEdFyvuNbMDw/UhQLX2dMpV8B8UEzoQQHZ5YCd6SjkllTcg6G
RUvWTXYlMV5GB509516n7Zb+UOYRWJIlmnfMwD7G2J5E+lHQUPTKPreW31vl5jC4
pzn725E07OoshS9UVQjg22YmqTWIs2kUJf9Z5h7Rqr6WGdwNDeHHU7RUDlkDsKz+
NHkoIgqxXIDzLCm6XYLcX6T9Sr6XSUuSFTe2Eh4cd+inl33a+RxtSLT9JW+5hsPV
SyMpkaoPlIevDfsTWai+l032N7GWmFHdP7bsjql8TG5a9DXgGw1foPKtxo7zkWjf
ZOyVW7lshaYWXHxua2WmzuI5GQQG1nJftGpp/1qiZ23uSDq8WU//CJYySdZlCdmv
FwZLDINR75Z07u6yXiKKoDjtCF9w2nzkHi5LAqGIywISLUGv6vKqKmrwR+atx0IX
X4I3v6jkXxaUeVJbgLGWsVhOfSd/yvG2dqB937lEtms7edBB9oBJZheTVwf3rhBW
t6orSimuTUNGWN5h2ipA+xPm1tdZ0FORJAlzAQ7WOckOYYBfS/atkom03gQ+BJEQ
UsV6dAY5m0x2KSz4N/lyaTJ1Eizch48DXRkggZPdy+pDpicC/DyRdPToxCoLdp8a
ixIvxXxjV2N6MpYWxerxupw/sisbcjKoEUpucEJR/TaYCIxCItPXBE0VqKLjdRT9
9VRL6/RJuoQHMDhSVu11WG5g2oZQ36f4Zo/4Iol9lZDirt0TNwxLQrk5buU9eGTJ
aGeXKGWH4R78A20jW+XdrcqKeSTjeM0YEXKcNZsz6dQ7MCq5vExfku2jNr4dIkIB
z+QkgnEgdSc7fI/Jtsj81/rPFl9298s9IFEJTIjFkfTEAfrcQ22cs1959plDRZM/
Inmvvxa3c8khjU1DSGzt6UuoNam4AdYjeie6raIGd1EUbvblaA/yuh4kqmsEy1Pe
pMY83TVne3HuXvsAcIw72zGzwZ8xUoJ0LAwsHYNypiTyP7PH55nzK1JBGbg+8PQy
Jfy8iC8vT/M5xpEJ6tzqTroEBfDwP430Wbn0+rpIAIIv9d78hgW4O/7Pm6R8KKtN
+dObsuI2ExqmH4CFFKhWB+MbtDBUO/D4ornwTMQIfi0iYg8VLjMop4i/eQwk5X93
cy1obD5+UromiWzirzH93785WQl9YRiqc9yf+F/AmFkOhID9gRBd7kR+NM0CFxBA
GeH+FPjv2VvbW72MQOHvpAaPE6pn4FN3LkCejMGWtIo8IcmvJMdu6ijBhoy4NinW
n/PdfK1p+CzGOFWpOayYvslkB+vPCi7zLcxmnu46R4g84jpZX5BKim5rOUOSj0ro
Yk/1Z5HT8swjyDtRdg8qbf8AGV9arTaN4BpIYQRiGnBnM6NbJsq95uXaXX/GY0QE
JBI0Gyb3nPcRJ4ckeVEY3QrHEmiV+qKsjYi5viQqHh2CmjK8Hb5tNZGJqAusCm4h
U66K/yeGMey8zbQbpqEV8ay2zkL1qwsBjPqDT9YLhdRDYiYfsDe4pgHPOsubUJDL
YNmbQrl2SwlNJIP2TnHQDbcJzIVh+9j6CycpXd0C40J36Rh/NLmOLgQNeGBoai/4
M+auLCw7v/k7hLVJHAb3Lqbk3g5vhwzYJ35soPeUO87BGUIm+ID6/JmvVJ4DGE4R
eu+633VoqncvUgfBeBVtIl3MMJHmQi1yUZT0C+dNPdoyTltkmWdcD4gfizjE+Jqe
qJrsqxK0Fpbtozp1n5gZnAGnHEy7sOgNfqXyeQB8xSoj4lPGXgsA9o4M8v19x3yv
RusxSNEMH12pEys1JGuCqTME7V8cdGW+G96uNMKA6jB/QHOJ9QxJnyHwSA0H8j0v
Ha3s2sJoFkuviqvcutn9TkNSpG4fa/cKaxlX6LZx5zpOWxHByTaUbfMieYrGhvKU
Pl89MFkaMof70uJW/aMdoZjvTpq7xIG9frkNepJMm5xf/MaIcLTBpxgZkSN6iXaY
7lYC5F/qtrG78AVSjDT3N1lwGpwZvmxh4w7KEgODhpN1ItjIJ9+mhywwYUhcs4Qy
LXXZUgcwDjIwSsKBiCbmVQeT78J0aLpx1PiQP86PZJYDH5uu+1nZCrkDQWclXvtF
NpqeCSB9mPuJH4UcyO5Zs+ex52AHONGsXVgPwZQkH1k8i39eu9uYpsC56/CPX2jF
JpWtlFHpLD9zvHTlLpUuNKHn7qI+mKi2Xuvv0SLRoa8vzdoI47mS6AX/AqixlyVr
ort/e6YP2TpGT8mHWqYPGr6kWGMiUyIVptI3KCvYbq9TcL7Um77lCVYNtjdtf5aj
ko650ilAink2U04d1QEd2YKJ7YWWXjH7eltK1jtRUje3UhBFrdcZ9obHhPI81egD
f8cjedZ6Bn6cEh1104ZnCF42/VyaxbeVXXsAM/sdTtIVhbADWkQBZyptsIl1Oriq
2M79Am0gfEeGuZnCkqpkjURLBZtWVv4nzETFvoT626+kGqvnV/iNf+ZMb5VKcpdD
5toc0kZgUhP1GI+LhlSD8Wne0JqAfoy9xKm77lr8Vyw4sat5j0I47UfcAW9F1c9l
7o2P3GgIWaHfj0BWc5VwjOt2jLP1dLg8L2siBcljAtchaKi/aLIZJzeKqiN7kt1A
CCb4QMCLWuGcyeMsE+BT7QiRPOIrBxGbCyTMomCFopns8MIeY+HHWu1hLalxpi7G
c3QaFlFkwY/xTpYFMtCY0Z6qL3l1DkRTQZShV835KeHk/Rr8s1Jhu4vo5ojmzJIB
FgyKZ72e9k6+2heT6IP2jbS2Hd3be2N7zC56psZbpuIY1oyh8ZLf1BKhmOjktvSw
gquBSwCgH/9A/K7mBJBjw5vHN+ZHVbF1kra1sR7MDxSBTQiGNDjKd4K7z9yy1NK8
DFtO96erMUlSffsvIG6DKRvAWutcYy7Pt18SINawhxYzNDBAMHuUO/rZENTDL8iO
Am6jBSeq5BKGfRauOeJOs85JqcUsd/HrxHCxFgHqWGLGweGe7dgAyMvBpGYIVeY4
LfFh/Yp5ZtaW7UG1UF4oF/hA/c9h4h/Qj7eX3o94FQp5xWHTFMltz6Gbihxp/dwx
4ApGSDJ6pT9VxhKfh6cVmO2dPbCXKSzVSOmfqrqYwORnwTiuXCGwCRabXox/bnkZ
atlvPptM7eSdcDfFhHPqfFTvd1DSXlPlSwE4/MxemqxzfTK3qRIJDQXrrguqNQlb
f+NvOM1my22zIH7h8Vrb+GYcdwax+MoCZNqdRV2owSNLLG/ZuV4smwfvTVghism9
/H+pYHRJjfUAa673fppt5srdAjGdvWdBUEGZSa5UoGkuR7nRRRm3GQGrrqtROnx2
xaQ7YRHpcX6GHqHtIgYpI5Q5vRIqDicgnnYE9UJqy50CMC0cMYM7xicwtM/Vi+w5
kYStNzrT8oItp00nujwEv9P7D9Ch+wdvjhGC2hhTB15dxLQ4ZZfojVw2BcqbP8+W
sW4sL40YPnXqCwUwkwUOD1CI6FxoWCe0MHo7yqULXPK988U7XlqfJKN2jkqIiC4N
BVi/OWg1SmkC8QitREkMBc0flgI2XNhiyL9mB9hODabCBArZTERiBKhAxBa9guqN
MBvXuqFjanG5o35toZcz6rztGLT1NX0CrPHnWXRKPe04eJh1IIPpHJXn2OAR98q9
+f+51Vg0djHO9GdACkVliAlWZjBTRz0yV4YcbqieQaWIWtNc/Rg4Bh5V4dQPvXtE
WeDFYgemrUhSXij2B34lLrRKtldrxu8waOFW2f5Hf26JFiqM/2feum+ftUdlf7Iw
LYK7EOESy7MvqkSx7TDUaAKWc4thNMcpLPbSN4oBwx6UoySoBHovWnRAMnZBQgU3
tiz6q6saeAU01JoKeCQYcHFayYB/uU5mixO56GYazrSeqops/WG/TNm9zo6dKiFH
i35LMZ6Nms8TyvfAfqRhyoKdN1/+8nRULXtKfXrZg/uTfQYqrI4AmCQAafnSd4b3
0xMbUMzRbySzeRqN2tkZSQdBNz8IDq8FmAqPIqxkPl4e/wzrhG0dwJ1+sv6x3q3U
TPP2Pq44nuVqbFwOrgd/WHy8soC2ncU4ry0PmNiye4CmfXO9bZX8FveyGILOOU8U
7ilHt2mjZjOHXnGhS068WybGEV8KByyAEYTJLkTj1DLuk+YMxbsIrQvZhMeqmrGm
7dOPiAWs5jauQjHwxd5v76AAFCd8bigNp+7z5x177+8quOCCaSHt6Mqo1uC6gRLj
mE1p8Fqt8QtlQgikA4Ti0gQEC0Q7VGaeEaOG2YZmuPZD0Z6lxPETlaZ6D1aIfmLW
VelwIg/MY3ji7aaWGZnKh/wUeHN2QKqu10zVNXrJIHue6WMZM6rQBtVlhmGz9Kwi
TcRi0uCxp5jZCMhq2YkHdsIy92tLHlleK/mifSz2VoDycSDP7vj5klZ3Mftn2Wtg
5kRYOycwzZt/iORt+dJpiGvmDwRZLJBhwfCwY6YUR1YzCGn6l0jDjp7D1bcGk8kh
Y+yRLMCkMCmfHMza5K1ZT3Vlpjik6BfMMsYB/S2PN/YolPKmPHLzzh9TMqbXltJC
hgtCBqr/lJCcbVfz1s0E3InF+w6mNO0UTupUHwFWABWdEKCSgKbwrPkDkmji0goB
pJnNh7ZA5vQFKenNgGia50sLeovLl4TG8oaUg7RMmOE940rPlFzwsliw3eI9w1M8
xqsYvzcoBiurn7HLUlsBBG3tfEF1nlgC2NA0nakG3QIDYr66DMIQWMdojFCl4pml
TEljTB8xrztkkvQXWJW5UXMiHyqGns1Ts989raI0LP94py75eey2GVLdaWevqSBp
MoFXmu+UIy+zIqF/jT+DsuMtZTIJ47hX7JUtQ/oE7tiBEK3vwMuu4U1tRvtDUzau
S3H6b/cE5aEYg/YHtESHfO59vscLt3INuo23rc6wG6G5a1J61Uhr9HhmZTx+OvCn
GjxP9qRvDlZqkDbwx8i+f+YgtGFg9/E8Vgg4toDXdTqWpd44R98F1CPdIuR0toSJ
OkjpCy23WHkzMBmGIIPISkDMcnoGKuJPuEQPkrg0rswQQcbkvp3mtIqDZiMUcr0F
65JY3z2UR53gbE+XGXGHOecQtTNtJNY4dUOFVBHP7tjAjTKn7DnjwbR0yB7gU3hQ
ecsBKPFIkgKd2bqX7d8ZOJbIV2PSdLSo1ZgnE7YrQh2G+6koZ0V11MRHxU2P4vfo
hQ+YetaARH9DPB7IF5fOPiwDQCNwP2tQG6dZjs6jZ+y884c3dAZqGJJ22ECMNrqI
cqYdIg2yBtNKkIj2AllM6+Adk/d/NiIlSNYLS4A5GYqFCXWoSmVwIit9EwO7E2A2
tKmEjNKG27C7Vpe5uKrSaXpA1D3u9Y9KZT5IYbLHWE9ZpAZ8UktXzkCiOg7A1YUJ
Yz5K7eTahEzxAvk4aKwNRbAL8vFYg3hsEvntPiqt1d/oxps4UwOFfbsKO02uQZKp
8RAuXI7E9ZtbAFSdvstTnaHiSSw3tufsu8MVGwxnz4Mi0o45imOhrbSLZMQ9FnBd
mmjoA+AJdiUs54OwkXZH3cfPr6uiAEbwiJQzibRonJqGaDy3JUAhPkF5lmmHmYua
nYMGh4qepYwOi/E3wzsZ4ukA3w3f9HKcie7cMy5svpPjWqdUpG6awskKu/aZnzqs
dlNF6uiZXMmeZ0POtqObi9o+8rZauJyFgNQfIpJ5VsdiB/f1LRA+Zfee5uoN/L/7
PaHa29NAE2a39TzFtN5uuP+Wsdzpx8JKhmLjhG2vCJ6jjSXDfXroAkjA9ncDT1md
Ej0BEqo0PDZeocC471ViEKB81ls/aZZENmttfjBI5QIeOBeREuXME10LDAV4SCrk
NOk+veTDEJLB8Q+mSwLVTjmTYqhqkQsp22qiNhaq+lIoiz1goSOYHdSdvn6OOKOD
4OloY2MA2nbB68Ro7ir0CJ14ugMPywVSYn52s2MYHk/TFOHEiIWDBTsxgRt5dA72
iY6G7eMbHpDbHJHsEGSoQ5RDDdVGyLwbXL/8SM09J0OsPAeL0Otj7FnfeooqSai2
fCEPmjiYm0urf9shE8sBUgvmm+aH7dvCIuNJBusVlgk7L7z1TKMenTeWAgu1bp9h
+pyL083fPdEdekZE6En+TssDM5ioR1T7VHFo1GdwKNT5s/9JY4mXeY07IkROvtbW
rY85V5wDAbdrDEeboPiRNcBXXTeXfdTODH3A+iWPi1JZO3tq5lI0lrd7Mn9vu2n+
vZ2XOn8nhfcoNmV2PpSOw/vD1os4x2hUv0VDIrV9fY6RZiAIeJlRcHrQMjZD2CD1
T6OO4KQGYUdI5OUjQfnwG+gV53pD/c2K6EMNrX5V0US8p5LGLu0NQmbI80sYH+X1
jEd41Xyoj0aqerXzXmv8bs5MV2VxPlA+jolYeQdtGss6VChiqF0WrzQ9h/XNMFVl
MLkeG2gtPO5ScyAH0nbMgRyz5rdBH5gcNDhH117K4qlKhhRgkQKAzLb58GiUE2wn
2klHWIJqlvuUjW+i0Amfm0a6T03AxDD+3NrIdRUSYf4Z2k1iOYAj7nAlJYnXzXeL
fO1jxpzV+hF8SI8FAK0bwLH6d2nwmZ08FUpK4xcEedlqge9IOWbOtVozIJEE1+R2
aouf7FXxChTP3lDfWt7ML2RLWvcNl/OhrOHM5BFm24s6K1JjL5BhvS69+7JgmRKQ
8qIRdSLP7GmTYfIEUnzaUF0UVOEYeth93UQdP6glsuq2+8TGnPqdwbKOrJ+pIn8t
s4jJaAI1HIkacIw4ELgptKunMOcLVzdAdPQhqgkRgjHj4TOJI8lHCPtqSa12giKJ
xkmJCvjCLHk68bobfHjNBzw+3Idxn0Y207u2YxzOyKI6Qyj2a9onBGkMY44JbX84
e2ppkHBtB98A4/mixj308wZ/rPE5IDn7+YFvKqJzOwKotTfUEeHBybM+shuu4Qns
KuVqlZEMmZRMZQYRC2OMldGIUlkQcv5maSG+5F7xyO97dRYfTmMFc0x2sirnR+Sh
AI+OlIiP7VNRwcC1wefq0mSdKvhk4AuzQIVFlmYueSNSenl8aspDUHAA3voa/A5P
P7io1EsMGhBCUSxYA3IxAifU/bPI5zH5pvTUy598bvaYriSa25PH3OSjyxkx3Zvc
Zz+VJyod8+91Yk20IXQWGf6QwQE7b1nrKQvrfbtTN2avFgWR9vNXFUnXtH9sp4mR
F5K3vKNkUFkkCCTgBMtnxdcEBUfX+TRGUeeiZLdXh0GREJOATZ0mO8ihfcue+w3F
PUIA7Ih/d2N90VFdVWyL1V+81WC53+2JpMl8rQ9A9zZjpJUozjAzM2iVW62t7xuL
nfZaBP0PcVKqCdsDNJ0Jp9wBeENHpvoAFbaLxMzhdy2yFgv78d53AKRCfHDg8SwS
DvFpNx16j4UPCd1Nknflym/GKtpK5VRYDUiMUocfA6KVZenHlgSzJuX13RNEKBuM
0UF/vTMH0q194902FkT+CFpWR1ZWLktDI/eRRBk7wrk/VkolkB7S79ma2r4ZVgA/
Hr6NMa1ixHrLojfyCMU8vekWLjkX/YkLzHhcOlAU+VFJwNStmHWpCGH9P0ykQ5Jj
v2akUrsjzN+fmokf24ro2/LyPKN0O5tr+f4mTIGhGuHOcNSuE3X9nVaz/9pb4RUM
EwbFhQTulhWtmxZ3hundIpkk7nupsyBl6U56MaKo3YwkVwOM/XipO1EWmMSMKsoM
kNKpfMFSAu2HUbdcvha2XLxllVbg7pW/FJeIYBTrddjKM62uCzIB8jsBuBlafa5u
ckCzCwJqDhVZzixYeObcLhyw57cdU612l8OliaO2FBZgAkz65Tzw8cqkHHeWbrO2
2H2RilkRdnU+wiLD63vhxEPn2bmNpXXLXbqdPxTzj82a3Qx0FsnMUxZzKOi6LXM4
2B6bgvYnV7AKvdlEdgw6wJEYGuHGew0cJV55XkxH+7WZtqITeKVIbNKykbO5j/mQ
0KieuyMbXs6XhWrEVp9QbzIGlfXb1kDnB2SnZXWhTPfFUpZdSwpj0nrzgklgpH/P
m5wz9knrAGdA/PUfOc53UMEy26L+kOWKFP9HCeZbf+e+GIXKnFw7eRvSjdMwmsLI
7svmyTL1cixUO32M4HxgBdrWuCq9BBbA44jWO/bXQp9055J17GCQTGamhT6wX2W2
+qtXHZvrm7olR0gby2HZVotVSDbnfr9FABbnjp5u5I3XszqqYnqdhGg5GwROzXNQ
x5CUDqzsFM68AxhSpmojyFq5hsZw65VYZ3Eu1vp4NsBVbY7EtWSyUjrKvPDYH73P
aqgYQGBQNZMNHPKKcvTBywOV9/s5H17C02a2kBToe0ZoOQQKPAWrcb8Jz90FKnBf
3AgMXhrI7/AVEhpPTZc/YeS6ozlVwrgzwK2BG6wwhiF77LCa8Uvz6Mv6Qm0HAzjZ
9mY25TA902r2N2BKNthP9/chu3gstMOZIOPq3Lp6BJuExBKCKfw/w4KoEMAQrmDY
Dnen0G9FYGHpDWFYVCbhqhI56c0oe/XcMC+NXIfn2gAGK/8MOdAnt67znOXIEHkl
m/4C2JyStM6XFjGkVRK0MP9WLpNChPHP5oedWAsM5OU9tjvP0leYcZvT7J2h8CSA
sp7zSVxBuKo9Z9dRKpQx7YIAY2K1UP4x5M0Am++A6Xw/z4uf4WXEe8Y/lZeMBEz6
m6sw+8NymhkyL8Y0kiUECmc3FrUYhISu+JbmjTaybK4PIfrkIrW9kRRo2VFFtruc
zWlxzKjOuK6SxUpxPi3YAxQxOXm3+q3G+RHq23wAzjouoofrfDANNtTkqHy++Jd4
cf4OWS8Orum318KpzQ0TDZC1f/OI388H68YQKeYFuuc5Xev4dtwy7TzYx9U4CpK0
hBg89MLHRTT661p1slt4rMRA/m9zPiARY+4+ziC7ct7fCq4Id+XomKM8QNgBVRjm
3oWm/aEdbNiO/R3NTDWpyfewFpDqXZfoVRtUd/kRFS/CNyIsKRdi1qmMm+p2d+wi
VRzupxPK+NO0kePGbPlOErTJ1OGwLqxrlCGsoJU4dN92OwbADsb5A0QHz2zzs+9l
rXw33SWYk9sWzVWdmzpvzXGSg0R02UjuQtKN2QLH92DK5u6vfhRSULm0Lh2LuYIZ
vK0/RMLbbl1LredSEYlXJf5ib1YngRgNAgc8E7lWZEC/P/NnQWPeVK8AJZ7hu9yh
U2kQMDesfH+SthtEqe0IPUOd2HuXv0W2WDok7SOu9HDcVt5Tuo7XQyV+tpTRTHBX
3Bj2yMH1LeiTeMqxF0WEkZfimZTaSCMMHMF+pZIbgVzZGYSswlPmbfv/LevNCdnE
hr5t6Y3Wgh9Y9eDc0RE2h/8ZCMWcySstyL3h3rs/exZ0hNvdKADwWWdyPYSWmGTN
ldv8rIw3yNrYfQ5w0Rk7KehoPFZxiaZu64iWsBPg45PzXGskgHJSeObTcc680gcJ
Q/mWh6C7bTIDm5UUAjXnKYtSqVHEqJ20ve2rZYY8FnhPlN9UK4wONRE4wQ9ESC6r
nZpzet8g+m6EBKkf45qXwE0wMIAQYsh7IRRZVQbnWOiW+WKFcJLZTOS2eOTeAA75
KZsLv+xWh11wESM63HS9GNYSQblHT1vVRsIl/nY+tGoLjR3fj9oGpryd8I/kv0Cs
wOEbFM9gvHc/Vul22qZlqZFIITPXcAhGAxtrku454HgwX52pKbrCa8AJmlrg8y+H
cUEecjC2Gc4wnQqoCdF4uVrWGPbPqnTcXlWXucCtMX6FVcFf0yHEMHSp/8Cw0PB4
YzjqlsA82LQ/64cNclXQWP6Gfth96HSLX9i1mPy209DjSvwgfWXPbjvKpgoKSsql
A+FSHPuCtbtYhzyxohTLrdY+L8jr+vR+2xbV2LEw1aiWpXOsf5kUgjeBnCt6BCn6
SGQzqaudkyb3FnW2iRlSpjYBrbk/TZI5rxC6IsE4qeME+vIUBItjQn1y1phH+Y+E
NG3QhC+7Vn+uwFcnDfNKTryHU7C0lsVdStfFGYO+RJj1J1rCgWA30L5EYmG9Klqp
9EpdyVRnBDaLCD9FGivfCJomaXII/Rt7VNu3qN0BYgWrxvjYW1ai3Z7uTRkGkwud
lWzaFGozgRFkUJfcACfgkdShP+y9fg8dwMvg1skq7i6/E/NgDVLt4NfJbStHNl2j
G5gL3fAHsx2KJhcs8Pyuh8whp1jVvvzPkUTxfVc2bkGa5QSN0mLQwEpBmfmdPiJU
xWBtzl+ypYwxUmpMl7FRousGqGIKgde2o1PKHJuf31etqj5op3BSRvmdeIf7fnwG
2QpZ7lcJPlnD1CJOP9cuXKW3J1cP7DUar+jAQqQS5jjbunn28tTk43iFcSvaqS3m
Csp43U8G1w0E6XVaz15cw5bbGKIhqx4s4DN1to9Ml0ZUx/HzHGF2ouxWgQUbNpvc
l/7FQzifMWUZJx6pjX5N17woI5/zsoss20EJdowNJKxsK571xxWxN1Ejn6mlMDUt
/Yjz9obkI00vjxVCt+5CcTbNJFcTPcK4jc68zP/cwAm62bnuUALeZYC1q6BydhJp
PiR+NL+W6/WSd5F9yhbOWAW3r0mkrjnawyw9hKGpalco2ieG1TGnEGSjv82ow6PT
VVXezso8yk+EoeVm5QN0qT7TMl5ry2B9BnFy2lUxg9MQFwRRhmz39/aTG6wZ6nsG
Tdgm7/LvquMIKy7kGlIQCWyAIekh55QeyBJlHrapa4IiCq5nKiFkVKlgx7LaBpJm
0X/E7mee9oOFV2z52+uQxhDSHKZLs8Gh36aOtPPSTUSOj31EYkfXVAAVSnGFg7AV
6KeOB+rUnRrEJkedaKWdYb1boZ5hjP/jehLOVPi46EQKX7dWLmzBrt2uFUY2vUIe
r0GA4yEehiehnTkqtnLa5U8BofEm8GBGJd8cZs3h7Uusn1Zo6wmcSB5xqV04gdn9
Am7y0kNqLucILbo5VmxzeNRi5uBsFZP3ikhHYvIniCr60CZs2UAHzIbsWQD+HSpG
9MTmMJSvDUOx53jFSkJlKjBnU//+juhQkjvCE8rtFFXasmQB1OIm/knRCJAswJsc
7CZHDx+qwOTzCtMRVN6n+flOAAFzdUaG/MF3OMglIJgD8HUkSYGWCReiATfiKCr1
7Zb0eIyCdYYjGxaDa8Ea1lgXXITmjJkp5jkloGkoCEYTAOShdrmqwF7WlKUJpxpl
t2YmeAWL8ydstJ/1qcGnSz4szbNyURXhCF72tUZeAqsQK+MKwQUjsX/K565GAgw+
29zVYYWz5A1TvU8VmibqDc98ttmHsFJZqGGWUVuvHSi77DmH95E5zg72esbWDjxB
v1s1KLA4TyU2UydN2G5+oKf3+lKqoBe1Eop2y6FhRUA0wNjO/fa5khRLYkuVa5Y4
Fg4uyOlXXOX1cXpNs2pwM+F85C7x1aCMcr5yyC5mRyUVD8YG9BmDZZIuchTudukl
KDffTZMXyrC5He4z6/dOTZe1+Ze2K3IDmfXGywd+QbhqNMSjvMqxpPZG2ETBCsWu
h4cW9MtK8fePKRGowb8L92G3pVICZda8fHODTFxGVsTRLqVX/vR7+EcG1ZZ1+1sM
0yPIa/ccSry0TnhzHslhAMx0T9D6iqfVoY4zs9KPnOZUKVHyb0IqK4JrX+3WVmP4
c61OosHTV0RD2Z4gsXw5q7c5OC8Me9bN/AfW8V/WsVtwaPNqT7r7dpDCQsYDS3j+
IAo4Wb6eICEjuY9tbAdVZWfznr2squn4h3Zvw1x+N8jHgqIdZpsqyKlkiJStStKI
8YKHwOPpBYipzwQN1Uw6GDi4SzWIsioMW8HFcNwhubPxqEUErXvJDzX6p96Pp/bT
52Ns3gPy1Ads0AM+yckmXD5jc8Q9EFJ3aldgKQA//yPvO3wXMgC1gzyKOuvRvyh+
KX7becyg4QT2/336w9h7OpLJKrarpqtRP2fXNhBNUPE9yjGbMIb/SgTKD6mKvmC3
RXe8k7OwOf1zufII/bdJzXhHLzC9kUvD0sO9np0hE9G2etnV9kNDiCwWDKUZo1y2
TBDLsWmwGde+VG2YqdD68oPBlEwScPD9BueWtst19QqOfTgBfd+37Eo67x7/aKQS
7mQ5kSodxMNgxm4WnrJFZx3etePaRKEQx3NK6W5wIJ30XAFExnplqfhKf0CN5NXK
/GN8+dGfetglsmHq8gAEhfuLFE75w7ZhMUvqNkKzuYSSR6DDWcKk4QJxlfnXN9oJ
1jwevE9bVSwW1dbdy/XIhzEsNmX9ZRJnnJ/ctY6ygROvuEYrq+LCnhrI2/PZAMMb
Nn+dgcO706W7ri0uR2p2Z+aCBRzi1VpLOMqwFjT1eNnr2rRkVFaJ0kXEFVEVV5/4
hS5kXgb+RATBtPmQYpAuUWWTPDIDC6YXhIgGI8NEGHBB9jwnBWX1cbqHFIGxkE4M
YRieKNmTau9ti6WspNsIyuvbz7EMqYf7laiYK5liIZCgTGE7zOG38KvwVq4Hs159
mr9NXd6UYEQknCJ/Pqd6uvSG3su/PttSP51/tifKcZRkpt+OY7Q9wcEm3+GLssnO
CntPLY/KqpstZKykw/sxdNPCTDllsSPXKs4XjwL+Dll6N/gI2LV/N5Wqm4i63KSg
jUOwo8E9Bo4wISjAOs3QtE/sdMUxYMtmwLGD00NlAJRh7gPnFpB7AS4iwztn//ty
EPgJAsHjoiKDxlVfEdTWgT/pqqDJ/nPk99cyDpDzcvPTHBgpqFOf6eCnzrWYq51T
tCgRY6gc/MvMSnP/eJws1VLnDqzR3+H/xbWr+JNJINLY5/pZILIFHrHvsltmMigd
0qHi0qw3TW3yuzJujrzvwJHRtd12RMquRpJM5LddvaZTzWf4fOsYYuOtz0hZsCoG
6g6Bo/VciPFIjTGLt+i83Ezs7GjXb9lw5NHuwwoO7GcCVQsz5Zq/K3/vCcEW9ALf
c+Dv8rP+CVO0NBVRgz7wYr7ebH8KHVJvlaRrpbDIuVkN/ryCy1EQL+nKJJHhLibL
/gmMmQwLQvNAjZZb4mNSHKxUGsVfiIdoG5f+vzyurPBUECzy9R5FIpDUk75KusQd
1hFic/f2NZyaQA/xox1+0aGn38IFQGgZg8c3vLA3nuHlK/Zs1j4L1sJegcLzlmgT
LV7dA3LZKRt8RxXWxhW2mxZmXSg+dXT68sS+Rd/o1U87xIJ1ZbL/w3fGAKI9mhbt
vftVSWAyQ2vb2EX08N0NvfjR8PkPmzWV1lmM7pjx1B1aJa7xH2mzQeXzI66GY34/
xRLdwwvc6Jwky12OK74nJBywPXGDtCMYVnAjYZA8dKR9jm/wlV6PVNy2LBYOuKc1
hF2JBkqjbxwlSOsAkpP6lljR96i8ymjbTPdb5ObrsazIUdthLq5fjTte7s8/LZL+
IvkIc6OWSvF2PkQkNV+2QlTy0dwcOXMXHxQ5B8IMhCDf8d9DNBvD/Qmwg8PDPLWK
hxxHD8cbrxkJOjo+uiUmL/DkZ9E2cGAdXJg21jWlSyPYItRk40skj0tSwauKtxPz
mK0c+QDSDA8IRaIMBd5yJEI7ShpCyxvipxPgP9chPYkEhulfzFfm4SqJ7Ku6rlig
hvcttyOGXm+Mb3EY55vpraOwxaSkvl7fUSg3c58tC6Gy/KLfi99UMGerzz11TOao
QUqkj0zcwCHzqr+tDE1+BINaH83nROY/DZPs9AG9ByKCYiKJeeYH1gGsMtsUGHrd
zIfzoTtCA6PRZ3wgsIAfJpnqTa+USTTZ2csQ+tS/gYEzgFUoMBb0LlYYoehj43b5
++yuDOtkthzOgLVMfBPirtYU20uZArwZ5fFsr83TLwgSSmLnczHxYa5b5/aILD3x
BO94GQc70hJ3e7+WDzFN+IrRT5ywc2xy++k3Bgcgz2Kjuz7G/Ql8TKXqOK4pzzO/
ccEC9Sy01jWLHx+//ngdFbpBUzmMuOpyMPYHQgGXo6Z9LlQfSo+D75V4hc3ZDha4
daAJAROmkx171AfVXtu4F5g/j7iw795nFvmrXfoKT6jJ7ZN+aumxgkqZg2tbD6JQ
fzsT7IFyFnbk7pUOZ6tnrlhYxfZzVjyZJ46rSg3y0AVi3RCtaTGNCebrV+qdc/lV
Cm/UEyAavXJDw1nES1Yuick6HZsZSQdGWPMf7lUI2cZ9XVzEP1z3eSHrlZUmarl6
NqTX1MIU3oB9DRcJXNV5wXjpAaXmtYm1yhQmcfYeIY/85Q8zo0SeroB9Avo9Srzn
dhYir+Fjc5Sowk1jzPwtgNn4JMeaJecGRiEBzhaUq/5sjv6x4WjssSD+pKsRTVN+
rOWjvUxgVg+omQaX+Tpf/8HJLb1N26O65xhN9py0rl3lhAWFMjl80wCEOHYjE+f5
p/MIvUv4inaDusr8lP1qRMr2eGbMLb2VZCQKhZ6ncWB39aRFCrtvmHBrPd40eoVq
/Ab3EKyBQr7N0NxlOEbEtqplbISfujeSlxXphb/PvBbwndR9uW4Ycit0lvZ7ZWED
j4WDphjYZvHMxTg1IUkvlstQnXOHuzQylZrHHo1MHpCv3y4hbDk6xqEPN84riLXG
gOr0nT8aSM6p4x79NglVMMPyI4H5crnTB5ksIu+2eqRUhsP95i3dmi5z9N8X1tuc
DFTyH6huzojsIdP33yKItZp7Oc6nynFvciEhkSTRvpYX4gIo9ExLPjAGDranVJHS
9Uk6PKOR+8Te+g2/RPoRBJCcjSnDJa1/YCNe5rqTFK7aBUl7/34Kly7A1YzJsVHY
bFEGdKZeuNI5futNZIdSS8fBrEDiTZKRNOXi95TJMIieUpsAjqIrkALKy9eerHoW
ZjQpsQeSQjeI5d8O8s20VpieN3Vd8rECCCTyTxfAmHz2gd1KeH5SBL2mXRykewDY
w6MuNv3mxvDudVWTv7e4V1WgGdkk11/L/4uwPGsr179rEFFNOCoayJUonJvfxyvg
tv74pcsvVoDp7SK3SKKyd9uYH+j7EcnyDigNMQule4iB1Fy7EhCTjEj1o35IWbKa
d10mx3NYDGkdhY542Tv3Dhm6w96EAK8hXeVoaNQjTAFd5F/rk3fodY3NWLiseSjz
n0eAdHwwtL739oEFAjk9i0qqDiE4zpB1l6vCHbnTtW0FLWr0gl7bhjgFuk8imCSN
L5lXrQfF8l1DtJEhAO8EQLjrtUcA6Ech1X5sOupHhEdykj9Y1yARrY03bibp3C4U
KEHVjRPht9pMmjtSG3K3r4/zfKYu2W4tFoTXoXkzZ+m5/8NlAVPNYA49EHgwL+e/
wDp0y3vOBD0bB5+k5GwhzXhAZuX6Daq9lYqVqt29clDCs4IcqYrudQzUtTw74Gu0
K0TsFpY2ldQMXXHE2DNBdytYXrRXc5/EK5K6ZcuyTXaWF7xZ8OpebARaPa3/hwj1
JeSf3FSz/xKx465YiunxcekMzzGyRsblCW3ynBPC/DbVkqRu8g0YDjy9Dvj89Mnl
A3cXdDWKf83vUr8JwFV8R0pIaEzPDtOLjGvET8BotDAR/NeBKt0ILQOAGpuO0qED
LT5MpA/+JrjePJvB15xdYx4SqduGLHtezgPhwg6QmLcUBx5mv3MfPd7K1ih4MR7O
Zrux92Rk5KJhW8EWdcxVn3RZzkNj35Dz1Sz/Y2aXPIcsO+7T7zeWpCsr5JhAeopE
x/ruxd41ZwCMcB/4bOQBcvr5hLw6AVgiVB23WdvrRYwc2hPGGAUv2pTrukSEQF8c
8RZCRbc5gg7yjM5VdC/NShPqRs5R3Qyg+VwgN6JTxMXO+sMlgeEWg+OXGxvg2nJA
LFsTF/Ij/fBkTCwNTCyaiwV9VUYMJn6tWVf2KJu6T8mzQOxs+USm6l5KMz0Zk5Uj
Fq530Df+1QqasT/eqw2kMEgCdWML3W+o4zRBs1u15LGX2VeUlMz4FaAyzGYm2aGh
IwxQDLTaJuiuRzqrQzVmyLiPeHNWETkmdl35EFhpZ4J/YDCi5W8Mb8+/3hZPP0wQ
CEVkda8m90Ae9pY8k2haEgaahWILnh2XtUT6Xlh/imPFl66zbESEjX5jGeGBO+xu
XkL3irmqiC0nuh1F7pYKyeK/nxhk74hiEwApqz/9po7I/VNyJT4kf+npkzGdoons
ZWkDrYM0iW0QAyXYGNHX4UKPiHWc40CziwlS/3MlIaP4PMhZnrPypfGu8eByriXZ
HX/d2OIg17w7HZiSjk5PFc63KjxQh2uKoUH1QPFwE97OwwfLh4vq0U1zAKD/XVs1
Wk1KF3wmfa8EHvOvzNekfHg7pDY32nx+5LrzX355jp+u7OiQsMCLQi/eiJ5D6rc8
M1zuf15jNlCYdUixNy8mX95EiIWd79CNu+QUmgiwjpbxcRIwzZeqhVHRAVEDto29
SysOwly/bkBINe6zGIzdfTQGtlfZO4n3kQgFdP/TFvoR99xdZy88S9Bms6zemuWk
qW/yh67tYTYBRE9440ogw2zO9m/vBjctZBqsb9YhBy14k4n2NZ4ncfSl69x7FVhL
HatZ8Iigr4QzYISvpy/ntW2BIpUnCwcYFPwRr7INSvLfoPxM1ROMy0eyrmGsL3mD
anP39ughrOjUYwXUYLeNtLOu8Q/d2BNMNy7z9BEFIvMEWaNNyRpWivj1S4PfvVdh
hKu5OJVE+vSO+gvIA1o1nMqTr7sorSFzvr3we0bBPZS7vABQr/ZbOx/Xn7EJIk+h
rIw+yH+0n7g0DmLoDr6P5ZRGJfegl14SONaETRVp+My2aRIu6fJFZa8m4d7si7Qx
4ECceax+3+XKSQUeaV+2cNKU5yRqb9VnsBM9W9XDvnpLqsm2SZxlEZcyheTxIN3/
xWzLeEVJLfoeoNQu9VQm6006SkKLzhz64D+XE1zQI+BixAgyr9jd/z9Bp0yjQ/xF
la11YWCuvpvDTIcXRK+2T0RoITvQ5UJxIOLZ2PfpAzTZbH6yLY8s0pzZlseCiPBA
GRVvd3VIwPsEuhbw1pmpPV5E6t6XxpMe/XP1GEPyicw3v8MVjVX8Ms9226Sx8N0V
XoHp7FqDeC8AZzv+uYt7MYTKdEYC0NLXXX3ES6sQA8ZNv65WmCXit5azBF1R6k7s
+wLi4eA356/DE9sC9ud3Vhw3XNgwS54lwujEG7oaQ9L75Km1Ih2MXOLW9GXw6u0g
Z6EO4KGBMnvNocpU1PVYYoA6r7XQkJ4vYqfA/NjDVq90po2ruLH6g6w2pQsUGOtU
oi3LNcMxz8lA32upuvYG13YMnU7VBfGfMtFUJYjhIsxFVSo+8FJsOwpKt4VVsX7j
gDBRhGk8HVn9zuJJ8/RRi3vxRIfhET+NGHuEga6JGq086pMn16PaiStlb/ZwrYO7
FQRuGyuBDx4jtxn4l3O7is2cxWzidN+9NubN8WJeUn+09I2khHWNioV4SIImB8jz
7OUfE3PiAA/B/VFCVXMwTE0oBehaEOK2MgZlA3AIqtnuY+dlXlX6j/i60MncMNBg
1bpwvGzlf4kOv58Rhh1qOrsp0BffCdggDnsef1W1dv5aknSrsrq3Uvmw1diFQQlA
LBffBTEyV5AxZJkPCyRjSuq3t2EOCPtSzZuyREAIpiu7g0W5e+wvlV3F8x88YvfF
hUkyj+Awf2m+oxVrix8o56L/mpUu9B2GIqxyAuKIqhyJIovdGzB0goUHPin7/xUW
xDZOHLIxm1p4D7R9MSzqqLzyp+8qlpllrhFB4Q9lVmOkYixvumDGBzS3DXogNhIi
XvHqkc5tjFwXPJ4c76nQOO6obCggTjTDWJB/g0ASAbQlgzSSZM6OwIheC7lzsxPD
Dt/oBBiXCeqai3/gYWYyWnVjm9QXPnE6wkS2BR4rq9j7I8Ei+CgXbnIxfbql2R0+
xQNf7862Hv+/dBALg94s4+FeyXUiDQZX6xZgQcH0y69GF6uxXphxw5JrYGAnWosU
SnnECuhOoaxh+Y84APGlFmxK1GBs7G1+tAG6OE+opzKX+2zSX4903A3WIA642iQb
zmpGW+eMiQimOZUH4Mmmiyd8lHUgP6iekuIL7gt4j5pYkllLcGRQcE4vALdfyGSa
LNaACEWoMgUe42efUQp5ENG0Dv9ZhIpZvXPDXHMqgZWoY42CEUsjcDOIKtjT6z+H
cbR7OBGXRbZ4H8cS1Z2nQO3WhR2RF/flC4h09gjulNFRRNVxpq9Dk6I7e+2KwUfF
T8MNe8BNu7dwLqIXqQwi/JdVE1CzRqefh9KbwPsqJrIAqvNNa9UfFNTLg38Bm2lG
SE3r2gf2WM3ztopnHJufmDqWwuNU/uaDk3DJtJqgdpyWKzW8u6C2YqPruaZLt1rD
AIcvxZDu6oFgOZ28LgY2W9jdiaskc8TbjzBz227MwUxaGdWsGgFjkKrDzrgu73Y3
zqTVf5fm7eY9v8TjItSOPA5QUs4WKzjnlvVEnPqKXcyY2wSyfWfPAljoTQg9ZX8O
MBAn8L7nFmJDYwEoSFEO2iUmOkkCfWKXD7Ghbkpbo2eQNZu7XPaQLDGUMyLIA9Gz
0M3rB+C2MVuGe1abmDHlSFG7cYaqJyknLmqbXIqYpjBGpGhANXac7wPl7VLwC7RL
3i9h6wq+TJDlYp2xKbLdzS1gmJfQSt+Lv6hAbHh+XSsxQzqb5+lVSNKyN57LYBvP
+yEOocnZIC0a8XEBMEwnzgCOGqOrTmJwsm0lPTMI8v1WqeHqwZWMnBC1Y9PAVi0j
lzBS5r3tE6kHuCVM/wKd38IHInaHW7zmIFfpEHwlbv+VB3cVax/l5tna6tThq6Nt
c0yW7Zyi2Dhzs/byuRY5llMdK3LAn6hHgtleL79FjmymMlmrZU5altpYhQxAtAzr
SKnafC4IIth5NgPCEiD+9X6mBDuWA/iyYgCt/7eDWqE/GnH64LqLzGnxrlTCl9mR
GVAHQFLSJEGKkvA8UH8Fuli0eJKcnbhfMV47w+thYq8/x3I6nuu0s6m5aieZ4ufC
eWgPNvV4NqjS6dsM7OlXauDoPXkjyuWCCHCByu11Ejrp7obIYgOAktaRMi/182a5
V5pzk1gKxE902Ok+pCH+RWAGpkhMagQtjPejKSUWoHSV8pNobz6sFOF46/C99kuX
loVNri4UejMB7QW5Ue9UmTBAfDcPI54+uc73uDQo3yWRyyr2dtnctrhERwQEcTk0
cEOoHg/qE9bR45M3m+Ty3kn/QpJ/sDEaQbcj/EHCqpf0IkiL66A5nKlXq44djuXJ
Ft+ll5zn7dXp5tB6HFjLZGTCMdQHio4DvKrSrSLJAkZaFAyIoWNwnlGbcDbJ6eCH
wXqIT0/2KdLaTxYbR3oRg/S7H1S72EqUu0LQ3qZm8w/9SrzOpJv3Z2L0En8LBfNj
yWOB8iaF6Kpa9K9LBcWC8v0TVuT5EuK7fUapUEYqN4j6ipU0IApV8dKC+5l3M8kj
GEoLGEYwx9o2wKprFps22D7YIpDGdzqnliF3ULOClTkiXelJADTe2Ch1gBJWQm1D
rd/7qs4tfJmQEzTu4il/B3vBlYvhQx2b4I5cpMYRIfnS6qehkHS/3KEypzoMCE1a
XOUzv+SPFbVwHFaTfywu4p64Z6qz9ZMFEQKkM8/k3yjgz7BxGvGRl+4fSRZobQ6E
3kkIaRsqhvIcH2DrB7UecZ9qVVqf289FOr3KLPImtYkPLgE/vr98fKjWTgr0xWqW
F76SVbeJYR47tsXUs01lc7tuKIrpF8MslpaKmWaY/XzwAy7DuqQbF1+68v2UIUXh
a48cckXE/91qB6JDB9h3m+gagiDZSeLdnCH/VD7FhvqtIPNQj62/8MOvgC0wOYPw
Q0KozmHqg7w2i3/axr/WBX5gmF/dqJUIs5kMYBBYL9AjExMLGnjTPl+vREk6tIgO
aY9iijg6/IXO77+U1rRSLGZgiIQ7OVdMs9gcXvr4GA1rUT7VJL4x7aK9lj9fOrvX
M/H+dJKRii9EeGjCVgOX7UDV27rN5RvtPER/J18TU62ftJCkwJrNweXsmq3R56la
EHIX2u1dKHmP990QxPV/Hfw8CEhT09wLIA0r05eTvNN9dSDTR0e4tJcJFWo8gIRS
BHW6P5J2yJ28OVeeWAIFDWM6cq46aYFKxo7QBT2DdA87fO576xHMb+Jnzh1g9rPz
49iAiyahkc87AgEpYYXnZpfujzCLazDUEHkhH3DARVpQklmmpU65Ezjlz/I3ys2o
aJKSjQ7gxUJXltpLrMMo3mRm80fZp7lQzb7GdLoJ2cNAlc4YhUexVE0HEvvy5cjB
c9sipYkDcW0eNx0EkgLWS66FYm5UYgLwq+Ljf5AYhtrrQS8F6zSJoa0nuZ2oGfDz
Xvr1uZz4P9CceiZQ70naSVXi/qD91d/r7fEqmP7YSj43Vk20D4pLLcBYXeYjW7aF
5P/j4q+Cp+vqKLJNkK7VfeEFaxdpkiQAeU/yaLuua/t+VmFlsLyPlsLFszPuEE5b
IsocOBxsyXbjoVaFMOjjr2ZJSpxaNiWEDhItzax9EGDy8X3nxh2sz4WIxhriuzOa
fvhEjg1dWdsxZ2q+sQz20lxMAapmnSTl1PP0/3G+xVno1HOLF349+Lm6b3JoeTnr
m0rNQoWHSG+o8KUMjSR/vr/RvstP/6TDi7tK2AGhEfyFV68341TV8fFKdEjRKUaL
5smgI5JMuBNH+hqqSMKIvqW9ez/zlTiwXy/434xh3n6XXG3zFR5AbCfNqU6owvlz
Zzvq1bcwj8oiIJEx3jd5Th7dpxYg/jxUXN+/XR0tM3iC67NUCcZlVX43rRq+vDn0
E7bHr4kkwHyekXuaOPT1N3ir9ca6yktFQLAh68wgb03uxuFWX7C2eZ8ltGhFx63E
cqs5FrZKHXyZZ+3YeTwcMIWjcdOpvVxjFBqUG4kN9Q1JMWhcCbf5LipGhLZKfb/u
KhJRiO1hGP4ltoqMg/tI+yJZVIuk/+9Mn9vgciUJO/AJ2eQsaD1Je7E2D0gEXXog
VqOfEHtvIFZazVjar0mkSoDsZJYDrJS27SuCC7Gh3UVDN7M5FUzsjdAUspWqo6Jl
uxBZZFYguS9sdab3ctNzKRQKvq/cnQTdZ6+oFrHU3uwKXjWNC4T97UbNMUm0cPjx
SoDo9Be9vZ/qtpHp4Bn9rYTfeY132+rKJqlKMmhvDy0Ylg24vNb0Bfy7EzCJu3qE
NBUDXkFzbfdxBkJSwZgIPNsSfgpzrT67rdzsPi8oiMjRs+KguwYr6ockhVFwd4Ms
bWNn2KWJoBdHPTGIssq2rojjviP+mr/FJURUWDXV/o/8qyGHSP9BS7kJ41G2gvwu
Y8hlICM6T0Yfeag+coVo41VXosJTqSw5EqJWKGJIfJDSvzidOO4mJLrRfyGJ7TnF
aQmqD/dTpbpsD0YZImgPVAbC5WeUAcWkAzFyeaqbKkspxkNyatxNXYqgp93PfX9x
UGD4/90DRSZBD3uOQ9IojgDE3et1Jol6nWd49+Ou0BLM6ho+8FwCwDUKRoVaO+P1
M+hLDh6b773gsHgL8pOjBCRqdy6XTESeT5cibtNCNFYvl9smdvc3oR2aRojd229U
h3O4RtZ4pFi5o8xSs+NhrIjEwCL8Vi57k7dho5weIn7vPr/zHd+mOpRD0/4HSzRA
P+8Z5Gqq8LfGLBTpIYYz8vfK9FCutxiyjZPUHuAMmJOoseRw8BaxF7a9pQG5cz6t
PGx7T9YtEusY/ImbyhpoNJg/CdDLhJp1mQpBhhk/0lgYzZb8XgFc+88MJ2r7jdNj
5HAEjv2h7NAX7LPz38kxz5WmqiqiTO2ldIr/i5UcyLo6x8rpjnCXAxVptd71XSaw
1+nrmq5FplUrp5cqpMWU6HfXI5Wk3Dxp44JtAV6bL7sFxifcCmwGNmbjp6V6+yUG
rhiFmcjiuK4kb57Oy3rgPIA82m0TW+s4igUtumKRrcY3iFf/qd5vyG0Qa784f6Ij
RG0b8v3voasz7jz05PFowTsvsuszYINOG0seicZXe7/Qig9wfSCgUzAH4tsGD8HZ
gGtnaPpjGd9Jk6tbTgBntzUvL1ba4urCk5FRWGoILJR9TZNCGJMGagMIRku0IqlG
cfjafYYbikvnWb9eiQd8aeEA9YVPUhnfY0Cdb8lNa/Yv8gzGkyyx+LeHDEJ/Qm+s
Pr9UKjRR+QG8qwuhim22QreA/kQt1+Lk+IsEJFp9t7sEqlQLX1HRr35hTmMFP1NA
ImuSnewL56pYySNAvd/grFBJ3HmyJ6fqt7QTd/BoMunWEpRrLG7nNoNUHhrpcCne
Eb3EGJaoUTa5dqvBYZ0xdFo1/FmRz5cEKGI9fJTaOLHJ0TsWIll/NBeQ5SUY/oM6
PSXJsghM6lZ5GXpEu/VrOTXvFlVh30mdt6vj3TUJ+QI7IKReIDT3PvmK3Q1ZWFPs
Xl53GzB5pzpo/n0bFLhiGOHrn6P5F8HrMtHloBSPXYSUczY2wBhqOVDp/dN7kfRH
yBP7wTSZLXIdcLfE/a0ns1CJK0YHJVm3oQ5OVlYNlLuS0H6RzY6ka1rOYv6Iykri
woLxGxBeC+7koN8yHRXwVcdniMpc9Pi6Byv9YUCCu7KJWqgqKSTDIR+aeh4HJaDW
PnCDTmivOUW0mldCP868Q4GrUXT4+kk1hvK628upde877ZtNxFUxKFnLZrYLdI0L
LraMaSW9czfmcekHKYYDIVJGRlQhzuwVCKbQjayjfM5X34fQJIxvTPtt1Fgoiw5n
T5vMgGVl841t19+5sdnMLvo6OHpwfMbkwDn2nEjSS2NN8QX/HDvWCte8gcGHVjax
3kyug3BCUkNQ+gyznZmzpRLMS9yXG+gqqm8aauOyriUiTDGVj6niAxIxbCERMknl
czO9xD/5F5bLeOGCaDmCkVnMfSISmqmr/FY0ZykvI16zIfjRGzpb3YcU7zySznOg
j2cmQr1Mh1CIkEaejKY42Ji+zDrGsZQ9gsKdGuwb77D9I1ZWm/t0IFvVPYAzspBy
LQ3xaRdp/SjtjKbSF6fWcLdKT1JxTq9fY09cSUclzocbjHWprRg+duPo+PdjNQX6
qluG6naW3Zw5Xas78h9ptA/R4m4PSCOnI2OlcT/rA2lMrf0hAoBZmav2+6BnLZ8S
5REA4Q003YRvSTZipRIDbo9uSaicRHf8ltEpyV8Qm800kxddOjznQibFJ0rJgJCu
20cJs5ADdYk71hoPrVIFR4VOiBY0ObvxyaFFZw6Pn+99yYRX5hbDMY7fwNKm9rW4
9HyLpffOynu6CxzhIKyi1lgkAkbGdUC4JBZ/d8IQ+ab5SNW4RH7w0HrGPdPCDpPt
BQIvR0tTUch5E4FxmO0mv2t/cDfxXfZRsdxWFnt8lq/vXMzmxgI58zpsEnySEpjN
MhZEkZFG2k/8rvZFYZDUeqM1OekvusgElwOweuuZYqeLds/IDUJ5UJteuTSK+saD
FNnUGFrp3m4MjzqOBQHEjTXI5c+IxmNudY5E98tKfT4PmnDXY8WuO+1SUb7vw3ez
fqAi0qhK9ZH3lwhXi8KYznrQNbKnk/MCIGEEycd/sc4BNMJ8ot7wRrsFy774oWAs
H6eqFXAzNnDVzmlktCvNqtEZgMz8BduIW0G1mR/1YUR5gwPEDVbtsgMHLUJSMuvX
pky2vFia8lFedTNCEMKjrczgL8BxBnmuZqmZMZ+uz/JRHUsnBfmLWLuQv9vTum2s
pWkixlNha4CjWOYzuAHdiTs0EUtT6vvK9HehYWH5mWE+mcx+FnDsdacl7nL6cxM2
j4sYDB9qviiQ1hZtPr47VEgEd0kCZ1MwoNjDHhCAEASyMcyHeTPMKt1c0BWM4F1u
VE8fGzk9u8yzT2Qkd3iqypjA1XDzvDvf8FATHUgEla4ioUrMhG+yA6eqIaz3kmV5
GNCk2kJlg1MdKXt4/lXO66UrOLDU7rEM70YQ4Oztie1eoDW/ZlRlMbyezyK5XrjR
OX/cM3efjaiMpWPJDBJ6s5pmqKl+Qc+Ax6VlEvWr0xWFV5G9oPtSY3OFCL3kJsHk
VA4nPJTR/TktZPC/wIDhLLyiVtsy3cK2tDxTV1wFKt4zMie2zq9Qfto99keGJoEV
UIby860nXlxO9385oE4CyJ6PljQKawq/ZPR6eh5qZksGjpt4qWYlAK6h3kr2xJW/
BTOY1C9+GfE4FbYg3zPEdtd+4ROww/yTj/sGRcn5MJqe+cX2BCEMLwanGK6xhahF
d7Rvk3o0SQCVhaNyLzS7HCfvLTGZPdfzY4r3yyaCw+8U1+aAYgBaIXj4Ytj5qMp6
mzBwX04uytKuSzO62jAXEku87TF3aY4U5a6tty5S1DhAP1DpBWwgyH99sa7tx1DQ
7A2a4fnWG0IL4y13fgPHRp25ocxDkWEWroRvXxP26ae7HQeJ75NY/zahRf0mfzgU
O0gmwAuhl23NeD0kWVmtn36tVRjYsW0Nvr1XaJ3/1Owv4k2sXje0P6zotS5vV++M
uB/z0xgDwnXwQ1SabKB/5YUdRmM9BMWFAWpj9hjUeF8leyQ+9+16jGAUb7UaC1dE
k0B2PIBzJfUBPyFrX1U8a/jPRTIEvjDH/OSUR7Sm4qFNrGFazngFYkoE0guByIPA
8ZjDBndxhsJadbo0A3qXvBl6v8n6/vdPXFCU8JIHNNJ0etuwPSapSzCNPTMqRoow
7Q0hZULBkuOZEAmZGTZw4teJ1W0fXssb7E7ABgu+Idal920g35TCG0FToVW6QyHP
1zc/WtJLYp3DuFmkHnqy2wM56x1ST6oUakW68pcpo53ASdj3y2cS29gMxL7jtceb
V11W70/V2iOqro6cxqkZiubmGNxiZzw7QIZyQoHZLSn4W3V+4oE/zwclBsoZHWel
YzTaeDMSwWBNSiC4jxWPF2pFDPKJlainET35SgyjANemFr+fMKjpuLz9myzGf5da
umpEiXQNojjpI03oIbtjMkOIS5fyx7fwTSFuj0MUqmJUz8OvNIX0a1tlwmbB913p
fM6ucwOOqXIRLkQEBsZ31Lud4i+xxdBBg71FsJFDFUWraXe5tpXFTCpYCI9lTCIg
Lkca+EwGFgxisN5DSF54gtnrN1XpIacGZhmpY6f/d9sFXTps6A4EcMFM3EBt1aIR
8cqxt5Dgbuy1sV7ykquGozexRzS8ccLUtY42kjixzFy6gWsef5NsqfNKQaYGNsEM
ESToX2a8SYaf0Lba900O6Q55fUYgQVPy+1TkU8YzVy5XKg6FLoYIc16c+5QJfUjj
m/B8n7D5eK++DsZoQRMndgM0fIWLPTD5jGLHKBfLykpjaKAlG3hzx8OH+sNMDiIf
8uZue//LcoRspBgJp1ErIImzzrfnJCbvwWbaJr5ruG6WWtFHnGEJXRBFoDzFUuBy
l4n0nO/3FxNarzrUXJMuudButzmT+akGaajdeVnVlB1X8TSHzhTC8YvztEm19os6
JW0M5qxcZvPgk4UrLxtZ+8dFed/mbHLnhcjM6II/sItUKXOKgouyjURk7licnite
RoREUsoKdR3ZZxAxBS9lbUszJ7rRkb8TNxUVbjMbjs4XTLaT+TSvs5Hf6QkPaupm
/uH3d8MXndeQfQ2aYFCDl3kZ0Qc1GPtnT4na8q9zTSqU4yyE9RLv5B3wc1zwsCgb
kGIZzXWGk9QsHcr6gQbOhRO/I7KWKkXFznyhbz2mdXK0CTFbmDbE8lyI0ozVmIqY
Xat5/kGWxl6LJwS7jmzOLyZ80UDhtCVEQ2d4eEnH1vnZN676omO+3fBcDTMch8RR
Za2nMwJqVNoJ7ijLjY5I/DWFOoB8y676+fSrQG8wksEaRSQF5iuesl6ILKA08/Gf
RgEIwIosJ4hf4O3DxQt/E6y+p00GHY8EllA+mBKWitO6xMTVk67M/Izl+xdEpvx2
NzYxbVuJpR06hVpBQ15WH74ofJRCYi4hs/ruSq7oLHiFGSxzoC355qw9IY/+zED1
Ro9Zk7uO7Xri9ybIfJcwZVjMInPTA8LeRM7SKhEhL/2kGcS7K5M5/+xA9khocyFf
nATPIaY0jo2SRLqe4XFv/rti33ZANBwCP/EPW5xUpYPrVBS/6qcM+aUtJnaAW2kI
F2/pT8S1omv8uDAHnPV37BhVoZVFndkpECvV3/3+NfBmT7BB7H4Geqoy9ZGKhssZ
UfY38EEEls2ZuZPg4ItgDhmIrCEz8U3aNI7dPz2MEcKoRJTffcAurj0y5Y+2LLjS
qiWQDN3hfyNOo/bl23kQxZ+N2f2spxUXF9qo1+ZeS458u0kIBPnmxSVGSlw4qKb7
hruFDjU5FD/xwiIgJvnYh0+zX9I942hBr7spnKt7m/Mtde6vu+/6CF8H2gWq2PPA
+IG9Q4UKF2qhYKJfP0IDFwgCl2nQjKQaCql4pA8TUAppEYe101JjrEQXONEOeQIC
PL4r+XYdYpFqJXhJ2GQf/8FIwmZpe9F7laUm5TrzKqFuXR4EIuxlk6SMPPB1tmbY
HmG93y/UTYRsFYrd0gbSkV5kNWChxZNkiBaPOZWA2Jb/oMSJR2p0njHJYFkQZAfJ
Oqnri4DQmcQmFmAn5pKYCKgPgFyMBO6t0oZXWPuXnpDEHLq1h1mGKzlezeH/3Ql2
57yLr2wKt5cFiHFFsyqkjB1QrwKDJE/66O28i8NGKnI9cLNb7H9K2fIx9CDRYIwD
OESWHUAUYtaz4lyAIaS2dIcd/G6YCtGXcfeYud4DMDtnjqjjnAriCxZujlyqhHoN
/1jgT/7PV5Is+WVh6aCV72wxk7B0sbQJ8BIb7u+jctMS+hN5HcBMJsJ2aqBTGg88
2AVyGw6D/LzAiP/42grXSgDIGzoOjKuas9N5Pq85T/ZWJ6PiWPpfBHylKH9xcHnn
X0HEKKKTCD7oFEAKKawDOg4sCWOPUtRAYYo+FgF4H5+Hgv32BDG2K5DJt34P5S2f
JEQWBn5qgMMP3ceFywBun3G5R23wPQ4otM9B3rykSQx0mco0DnjgXl58TBwWIhdZ
XeUl22qCIURINKXJnLlCh+92jJQNc/wKkwOrr8BKMtVv1uDxOyNtO6WoBZbFacSV
Y+2rlJwH16QvR/FTDtSVZv9UTT/xHHyrMthFcmqB0RN4kTzMhkabZTYiUklIPDk1
xNPIfJZBsrVemB+538SKxH8N3xlIigydSWi7VHchrFH2kaLIJ7/qDdtD5v75579Q
x6WuyPZ+VbELGhk7wMhxiSEogmZOTuwIlrf4idP3Rll0tjyFO1nLRi16/TD4Srl2
GnRHnVy5iB4W34TtyCB/fQwpVbDKzA+S3TmoMAtWc5LZo40+X4zIu3nNgddGSEOz
H7+zP1+s9OPloIVQ6W+Ti3X0dCu/xTC3xxbH1KVSW3gxxAI4qN64cNwxkvCG3mBp
Q8J7m/zKi6gwwh3/Fw4hSM4n3+xo1hHFQyk5B1Sck9cIdGrGX0qiyVgngrbSehzl
8HfaUeXjmT8c3YxqOa/WVh3CIVW0Fi5SFZVuVNW2fJqY7VQWmQ8p7DkczJ/edME/
YLBja6AiorcXor30TjKN38mUDlZ9qC0uzN7Uvo0VBGmDPNQzu3up+ZTiarf2Bahd
3A9SLLx62cRM9IdvbZyUo+EFHfb9nwK8Ll9GHq7Qs2pGtOI0OH9A4qEgGX85Efzo
0W8FPs8gQkhUcAW2zwTcxKGz2Jlp9MdujaDaF/abNX0sPM4Xg2MubMSDK+i8hZoj
ocZk6QMUsAZWh4bMoIQHaLDIxjkQEeOoRa0rj2ijHu3GUoms1TLXkZINSXFkTO26
PEPSOQAhxqTig/136IfWf6MqZK6L0RHbn0CoH9GC2wwA6HhiXBVQmRgtekbW7nN/
IL1Clj7pStE5kQSmZEQuRA3REAn+VkyihHWbNk4AslWTpXCzpae+wKPrn+aaJwx2
daY1/XmAL7Dlk38ShYX9cRG1BSqUwDFDxZWmx1ltp5PlAw0BUDCHzNVHSl30swL6
XYF3bokvCCOmO5XHETD6JC70iPXu5Rg4CwU9xl9+7aEGZUmbvbBbuaRnkju3i3YP
H+DtQnG4uCBvyQtL14hL3h0keoEgN8zgMNeyqZbrcDpbKU5EZvHHTHhDS/XUmTq5
2HLAj0jOzbafDI0QReg/+x/N9nxIWrIJNISHwNB6XgY/a4HjhwtEk5Rjf6gPmRdF
hM2AOGRBm5sLkLYB/iFL1CAoffEAuFv0qbfoDW1IA5Em/A6+WROKqb03vB8C5qTG
1doSvYND4Zx70wFduw4wEs5OoIgVSPiVmCtnQb1dGBcnIcATZFa9XEhbiUKzdeoG
hFALENRKv+0xdygqKvr4qL1fbHenzoIYIx5eiAW5K2QKvQnEpmjaNPQw0GdupoJY
9lY6HLOJ+FpxWKzy5D1uG6dBI98SMwPQIL09XZfLC0A6u2DK9M+U/h4HdjCDMppU
2G9I3HvDKpJXAWsEAPep7ZHT+QPqqivgkg7q09rrHo1SNmSOj5QDywxk1a6UFNkS
2j9A8bS4yr+yXgBnK4UmQglHG2EU1uRJHna41BDSvqVS8LMOHJnh6yiyijgcjIOM
xB17Q+hiGOdmjBPKz8lCTjSgj5p4E2xB0IB7MrLqFSCT4jgjmOwAfk3ngqV+hBww
tU7UX+ZSFGMYVuyqdY1wDQ0UK/ZPH+VtleDAQHsu5dDkVy26sy0d2nGZuoeEPEQt
MAQ5VrTIDbI1r1oTLLe5e414AdUxZuLY8LDCoVf7suMi/FFLEyaIQL/N8P3cKPUp
RNnl7jhPSGLorX63mIc5J2xdnRkDoAOKt/+Tzb48+bkBQBdVV59r5tFUOP1mrvIn
CJPoVW0zWhzkThAl5ZeLKc6xc2yr6LrJ8tIMAjyTDo3I+B99leSHjCU53TPLmFZR
Off2fRbxWiM5/MdfvjYn25BfhSDkL0nxhChT2v5Hp2+B+JOIIeuRPi7KfWJ598yF
Q262icW2AndL7J+WhoSYAQzQw9Oh2IkG+LeAnlvoVnrg4GUyKiLPGGuey3y8VhCQ
jPOQE32emiodIYN9O/vXXTAPmYtkbi63bkk1DxxN9PJLJIZSaS9B5HgdGT7g7oqK
vcI0aEThAit1tuzGwgpGtehYVweCH2hsN1X53sbMxAkfXGPFSIKD6IN+yAprwpl6
6EcFm3crhCIVSYsxsJZhPIAL0IuHaRS5YS+dG14CcRKOXZ10qylsEo64J0vcAwek
reA9Iv40LPMMPfeq/y1njGJbsHMZmWhV9GaQ+Dahg/lzgHcsi6trMNJNzJ6sSTK5
Zk7gOQvceGCvzceriMXUWBAUPFNUTEEcyrhAafjD704ZKsyDOQd3AFBboGPRu8LM
7mHvkOwx4RiMWUWLIVynn7v3eP3xw8OMCv9PA0z2Bj/wkKBEWsEW+F4Fs5nNXKXN
VADO4Pzf03W4y89FTRG+5TDV4TJ8CIAk72FPyLCgLpP/UCw5liBVbw6UjhZNT4ST
ANRbuUXVQgGeqP9+Q79cnnRWRKkR3RrYx+D83YmJcBkRQSWs9FH05cKVatHOD4Mz
EXUAIR2UZ0d4Q5C8GPLtFCAb0Y4i7cTJeppsUG67v13OD6Xid/FzF0SpDeNmwU2J
xGhOKzT5tMd5tID1Kd390tRLfx3DEs5/64XjI6lrN62V6XEogJqi4iOWJs8mZxA9
/htR+I8GosEP+ekXjw/om2arzNghfx+ZQuBRx6wwy1MA2TeT+8DmpMMwNTN1ctGu
UoY9bJ/dj7gb7i83Dt5ka5RXi72/Xbpl4XYMOWdws8xvnmZlgp5zKckJTDigoRF6
vKntWYNiTUa+oOPrD3GKRi1M9P6lGbHV32Xp7B7k/rLi+94nr3MsN/Gi/heXka5W
p5brLny+Yn/xEXALMxBDzoqImRE/BrCYZ3HaU87nuGTiz6MQln9wMI25ROawlYic
dNnShW/VyrCWOOQqoHlBS7cmfBDbMrQCukaIxvoQygPo50v8Vm5KqBVaMOXhKlXB
CZiWV1XLMFIDBqE4b7vT1bBUx90D6zyKjvcMpeXZJxqDoJoJxNLOF2kWIprwS9Tb
ruF43Km5enDC3e7g+qws+oEEN8N1D8fBUqsCVZ8nLV6BncK2/hO7Px3r6bZBy0kh
HhJNwOlLiZG/B/yboZRuP8KwBlsK/EpIcdUHDsqIfp86iMnlnM/+m4krAVVQ/jTJ
mSmjhyC1S0fsOXY85V2+PJ1m6efCYuzMopOQ1OgBEDHhxvllirVLMutMNv0/5Sgt
CfOxnWhYHNihiGXrUkKWV8DvvlaBrHUEVRmeGkYw6W5aapLgaYlt5SWxyB8bNlAq
4MxdlLCBMD8vl/H6wbnTu9yqecOPFolGURumHeHUp5QcqbUX1AzaL+59eZHJFO9N
5A6DvpneShkk/RnWmky9sQBBRUBzdJccXAAZS750ht5nUrP0X2YsrE+GBNrmIZnj
oC1SXmC6zJj73kN7LqnZbq9DxpI0JKsC0oUfdSoSm3kKXukYa6/7UsMiJBVF6mIA
hlmthJT2JrVbvHfMxofL/OfdCuM+yiFBGw0eUmjIkFoIc5fWq/XXqwgmlouJ2GLy
RUD0jVIHrQf/YjN9TL7Fpxl8o1oV5AWAq5f40ZpSDeqIB46w8eUcyIr03dolSY2G
7ZVjHtqN31EByqRmvNgza10cHk8B8BUnJJ9q8kHNH7bEkV6EsB6rmyNZIdSowUOy
/S7riA4Ta1suaqcwZYuJXRpQiwIbfwEt3MKj3JnGIbXxo3OAIphNGedvDJf6yDjW
gyDLe6N3eQqUcmEuzkos+Z2I33wC86UMNG/d1cTJpwqpc8NmvVUa0/UAPp+3Upbl
w9Ek3py++5TBBR4KWnnQIvFwNogTjaRxHdhOKEYbDdC0v6Qy/OsYG5fQieqKE2+5
NImq53NZ2GSTPXQojvw32T/SB0YaE0Yc6ZrvLlWtLd7ofhLw/2JM3FAggfFg2NBU
8QmipmNFtj+Z+u7GO/n2RADHqCmlH9C/SeLMZMbKBTfzbwZCB60Wtp2q1iAuezPD
XkMJk2uLelWPylQgTeH457cabH/Cx2FogSZ6Z1oEBJePNEi9bGSiyxfk7oZ5zsDv
tTURekQNiGP5wJttKYnpynwP6+f9sWudlqfPfV+B1jo41fIuIylmDEtgVCA4B4Vw
nRqSWmT8p6uSE01w8jGP3OhVwlO5Dgi/8b5t5jaf+PPXGkTzk5kNiorAJ2G0fTJh
O0Q4fl4TAKZ5UKN7DX2uLHqmppEGSsRgXuOpQdjmBzR0C/8gal/gdoxnifBIhZt7
MNpg+4piaRLo7xPbSoOiKzWU/Z18KySBMW7pplAIYL8oYBThO8Tj76U0a1mZIuno
VtdKPf3Ki+QWSTKNooZ2PLYHNR9WY8M3UPpxnvBl7PgwEC56IReatZIBwR3sdUlj
OVp+QKv7YPoFTAZlbMRD8iWUfDOtf8wb6W/GrlLF0QJBUtKSUsltfPy3WYHsbzeL
n1pyDG79T3jOpTswLc8+paoDvwRP1edsjsLxj0SerEk/j+ufmduRdJ04+Epq7epe
S4P+rA1/Z47ProxT6xWei349xg3BPIyGlt0YDU8WY2v1ohlm64qNcr7f4JlPgUtW
nqQx4yZua7jaK0+veu/nttXGYKwA2PYNOjQjHh/RW7HQQUW3djC7Te8WepOi+SLx
HgSw1Ld7giJuACkqZMS6OLpJL+EL2dtFtSv0g+sGddkh1hPEqwf0Cer8VUyiMgrR
vxJdRBKLpgxjod2xoJdqLBApbcc/MZniY0Bapuj4ey6TYqd6wlBl4XMm409oGzSZ
Tdl6ggF/6k+9Vxc0/f5YNTssc/SBbq82xbvAjo1s6gh7hWm2KkV5tz/nQzJ/VTgG
zqYYRS41B5a+mVGAw5paNrQVhqp3GxZwKQKVa24469KCaEdORVvq1s1wFJoKzUnU
rXb98YpxraEiU0Z/i9/6aEXcA3A4R/vpKfqvre+SOtxhRRO+WG3HmaQfuogBpRbH
IF/LkciOA35vl+lVvUA3PszXqMrbx93o9D07gK+qlUV19hj97T8EBAM/cHgnPaug
7ze4gvtuMPqVLDLIIMnZcFZfMBg5Lc3f6UTmipK8ejPJ4okAmH3ENniDr38oKVkg
KwB6f9Pf1WQ4oB1Weapi4dk3Ln2wyEWbbhZiWUED2RzGP/bT9cE6Gsl78wGLF3eo
4CpjY5v8VGfaH5I7dCQ6GM1wHHDMkQOllGFPsGrJQRVMPOeZ4FgMJHZRyOR5MYVn
AuHQ2rnEx6m4/DfMeKqVBO3q/5O+bC9uibx5dtu3fs2Hwv36OVRNjpLaehMJ4Jv8
mp6NIgsc/QvwKd3uDTa8eJeKbNxWlE3iUurD8Th8st2sUNawLsU9ebaZfymITMpx
6StGwdD3R8JCPii1g81ML8rejJn0oHsbTu5zxOH+Kwyg4JfU7XqzkmYXmkSq0plz
MHCPr4duI5KO244n0IKS8AcpmpBaR9FxD3YnDhJKX0soN9VFkdLRmr4Cey2vmkPi
KdBE7fVlFGJuDez/lCBqWleFOZyhNuGHUh/rIfUgYrI/SWaUfai/ttBlJg1HlbGb
vlnpFJR99BIf70fiRZs4wSBzL1sJc7JdeNwX6ChZZkFi7628fkvHpus+zvx0MTww
S0+7zATT06s4jIWQCIY+njgjp7lmGsSJulK/fT+LNvgtnHRmORe8a+CjNbLNPAHY
zdBcK1mSPHaokIQtwgsf0YF3EI2LhfueZ5BtpCc2wAQZoCD3ZKfN3t5gPklsOBt5
T8rsRyS8KAfb6NIa9csLsN3YZicbaxciqoctMJHMck8yxsRmIl+7jjDQ3Eim95mw
vPJAyICyCvJq/tbeeKaWzuIuUZQd+P/eS9ZskYPJthUOdFx/uC4RqeBkfbNJyb3z
Bv7BjPgV45kR2LSYQMAlbW/S/+iCRRI5ZtB/uqEa0fiw1GgWU7wfU9oxMYCSkp4D
3NMQFsVi720xH4fC/zJoOfYfgxMQYkl9JqTX33nluIFNsO5zDOvMDeHpAYepja9q
1MH71qSLttSSi/z6jOEQMK6brxNvvSeKzIx0YcZxaG2XXltpO3e18Xdi73+p52h/
AbSHTKcafQt1s5yFvwIGHo8qm0Efx7KN2uhqG84dVr67KFcOWUWvR+FAUuJ5LSyT
M3dAC0DTBJU4GuEF9JCj9UMpm+AtCxCdF4TLRqnDENfBlqvwxK8jlSyhRRLgXoaC
BBHOTSc/OMOLg5pfQzbagq9Pyky5NK9qltgf0e7fMDv0ihSL7NfjpZc4vVg+zbbH
T742fGLu/xZYpfrNjq8hsHlNJB9hIGtXoC3DkqFtOOo/bF9uIqQuRE/lBTbjl65P
fxd3FliM+RZ5X/k8MU4wcyfUv0NIF1Xti6VSAByL1wc=
--pragma protect end_data_block
--pragma protect digest_block
pjU4FWBqsmRF43GJGoQdspsvq2o=
--pragma protect end_digest_block
--pragma protect end_protected
