-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ugDc2MYfdce2gjzawvnQEZ5dfXjb0AELF4B9q1kDtnGGgAxbiWcq8Iote0cpSJd4ib9vUavXQE71
2AZ5sjdm08nFFBREpaPXvXcC+oDKmzYc6Xxcb+9+5G9R4EsH4KxbQhO9YDN2ztMHt7tKqAzPM1Em
NxW/CZa3YGGiHZMwQ95HkVfsWkeCWZPUUSj095s3xkvtg2yrfv+PWN8rbmm4opD3V3rq9PADs1cg
Vlcb6yIOi44p5NsWnrBgqo+69VD0q6h8oeqbE8v/Z+KF03htX1fvhYCp7nkVJFTmC5M0KKj6NwCh
IQ0WRE9n1k7+HMmZjvhemqWdRzp2vGeFv1jscA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 84752)
`protect data_block
ZDxCYAMwNo46XzGHzejKftBokvSUfvfANUO2fhd9IKryUzOkHrscHezYbF5VHpyh8RC+o+9FXL+n
9tFlzvNmyfQXVb2hi7RLcNUQQVF6FCWRq8/CqsdXXHwGQ33EszKPxtTTp6PZ6knAWqzspGPBCrop
ZdrzYn0GwM0l1VUDqX83GxgqB2+jFg4lKuqK6gAVRMSu3qwsckj6WdwEmn//o75nbN1bchHB7yIG
RXO0rWmHVYh5x2EXmYFbicb0xoSxlv/46VXj5mKrlKRWrhYbcPTGg+h/VMJ6g+MG/OdiSj3k4swd
b8EAjPgEoSvR2NmQNb9x3tTOrxftUBz55BW2itATXj2naQCXSHdiJm+Z5lgcNlCeuJs9Rg6H2BZh
ffD8Zwqi87FyyfkhxGUMXH0EOHqHfc1fwvyqY0cO+j85n4x3DNrza3P2H2tati1l9oFnEiR/T26f
CuAmc1P+TaarfWSiaADM1hLmqXnpMxoWMLWZAm0ND3OQulSf40fyLPvq0JfzFDBV1OOW2Ik2KmmW
nySZr3VG7JCsHTLJl7oOvzTBTYey+p87g1DolwhzA+UP83xz7pnfpR/0UovWkX4pPgb3x8cUZ3Vn
RAXlqhhNvMj/Dst0DyKBasquK2C/t4FWkwogIEhzE7BpKJJhTQvyIVKm0aM7/NtSBrTw64hG4g7M
xkPSbgQv0p88hfT/t37qG7Q7AC08LQZLmmXBgblv16leR9JLxhiSpXjwjB53W9utnzfrYheVYYNk
P+//jEyMLVQVIQMUdZeaOs5MLk3p1g5mmfRjUHupxHan2o+K56QoTBasPqPpxeaiqtg3Y9HM9zws
qHbZ3PDRecliHiRfnUMSN2G0u6lcPA3BujDAohsap71K8aSL/8qRpeOdfluBaru51LBmbMoU+E8l
eh3IGSeaIWhOov7yIN3c+ixIKFAvKkzqESH7uDrGxOCRu5E+g/Zxhafc4nzbTR/JugBykCHwGJsO
YVX0iJ63YlD6ojy2DAK6czkZdWN4y+uajeQOJjxaaJQmlwoyIQwXp9mIIyomI9iV9K+T+48rPgBm
z1w1ZXwx44czrIxcE9PCTn+IJajHTCoL8ZmYKMk/30epwLItITltDLZvTPOpy996X2eD19cRdkSn
DmXAnO98+UkCd1xtIo2fwsUxucoTPhBG5NPXk2OEl84mgpCf76aqVWpAgSZ/hG1bE19Sh3sLWHw5
TUaNRvTCxYiJpM51gkuvUqsEkEjolSEkkvxxxpo8rV1i+uK0MUSW7r5VTLnqGJfHADHytGtDIe6s
N6+AYOeBxFXlZXCYx3Dx57RZ8QYQphjUd2o7Kixl6xwfwFy9Zpy1uHXcOj4y/nodHl9CtRdfczgA
OSa+ldDYXj86TdZBDQ6U1X1J69GePOq+pePMAIebszt+q6C88rvwM9PXEJc7I2MzUCqortW3ev8K
wGmZDP03oOsfFo/X1eXOQzSNi6oyo/AntCTwAIgCJ5cni9X3kK2KsDBRdtA5T/+CRRiqM/P2eWUJ
osv2Bs/6q68Ix7AfQURGdbGhWIy5sXRxJgTQGLlO5r+k5qYUzyJGC4j7aoqHzj1Loyvdprdegizk
UxkjvuFtEyDVA/mLJq8XbPSOj4soNzQASh2pA+1hMlmQBHLS5XPE/6y++/0ma+8eM+WoY5286VFi
hrU2N1uKRzDiMXuCk8Mk2oiHU7jyN5esIsI+TbzTyuSdTtRBDf92dSL7batRW6GDjb87NApgnLfP
9eQAklg7zXgnrEUNtTJWuyvGw2EqnTp288Wnd0G9duH5xHZ0xeVcSBorlhBkUW4+u7sDVPT1Zzfj
Ne/g5PmpeYbgAqUFFLnPubQK9GpdsVpV2Em9phgxyfoMtmZAucWVo0tEmTiFrfx8Yg7vcFB4NpJ6
pGMbAEsDCaqv++vq1d6znFTxY1M6RcHGSra7ZFR/kM+odZSshsmdHu5/PLHajoXpr0fI84fNAW7T
O/rYXiIrRuBORMumwkpPPm1Y106quIL7dacc/UaUBZYfIZmSlvoxzYYSd2ytPgUs/P5etFiEuZaQ
nJbcEPof9nOyC3pbU+ydpdbZgTrYRbUSeb4L+zVSBSNTCcdQGvX6otm2Qb9a9DUe8Ncc8ohFZIUf
e64g5Br4PEQ2cXxazlPiHNHCWlOlOf4r2auYeAHauzTnPBPLDBpZzKo8f51VyI3JXAlirs6fHXQg
3roqwe1cO1oH6HO9x9JOCsmsLax9nRrzL7p4pUTFadPaZr6gWCBc0ozPhyB+gpzZsWlsaw1QVvVJ
3sPyqcK1MnIMHctKl3SMmQF/UIJ9gPCnfnJ2s3aiCTI/7tVB16/IS2o+XLC0WBeg7/h++Jllt0Te
kN6rF9Dl6gTRRfSVSayf4fr2E2c55ilD139LtCiv0NH027usb+Z7p7adHkOgRvsbbpsLTDpZ7AxR
ow0HszfcHpN1dZjXRC+MjzR1aeLWlbY9yBfKQ0yGpaPXL+YCFipNl79wz9kP+hYCI//C7XVofeKT
LqkQGvMAwpAqYET3feB7RAvbsyusPaaDWbTkpTKwvazcWL8L8e3aW2QtkGK4L85YM1N51yOU2+l1
Ppdrq2jEpsT4LuinycNMu2QaE5h8jTJ7+9VeEyOrC2VDeN99h7OIZDxHOVg4Yst9S8yz8u5uZMNS
PE6C9nAgufaYLk2f7GPpsKk9eiso3mTUyqVj/JhT/LWV1xrdTOAMtq20NdlPkYiDs/aAEUhNsp5Z
U+SVdFX2nyYsZHJvqNIn0H/DAGDXuZJRBlNG6r++LEySuOYNuoFee9gr/zBg0wYy1CAePMIXnX5M
XiSftvIX/BGiwu6Oik3YryfaODdv03LhyQ9dPwEbSIa7+SVNWLBdoIJwq04fohr4SdIXJnvuS/Ud
i8rqqjSx6loLggNSVZXavmHsftOojGgoU0boOt1tg7AbWy/3ptfDgwq5ghMsrInmYwfhRMJTeGiu
LBIW6/ZYqwLwdebfgpPn9vF6kXbEFXutyGglFVSLyz/Lt11csxy4MzzWhX2SeIK96STmtl+Y+YIq
FDlHvRNHjPQtKcKKczxo93JX7OnzV39BAdH/hmOl4cIMgX9lAv1Ac9C0PNeMg5SWLzyPuzP1IqVB
iYjHLVinFDUAnhpQki4qk/jQydcxWrn5iO3kJbl2Zm/pi1/CvLK2XKRSbsysWsBGfiGrJPLAvE+x
izlMWMCZe/CwXPLBzJld6+Z/vf0tRKTZ07JBnv+8W7b/1OV1Em+zw5B5VoKu7M4DPNunfgHnCVkv
DHrUdkVvfP0t4jrrmyu4i3ybWnOMVSa45u8SIesNPkjRjKjJJzcik10ozVpW7QyQ0NM/rpKqIZ//
RMBvMdVxM6fRst90bZKksOG14HyYVpI4kLhMkTEimkooH9Ecsx3wFqPv7NlOUjAc9Xh1XuZeMfZe
M9lPvT05U1PXhAZlQlrj6OQH+7BMueENw7qk0SUjRBHbV4QffrJXIiFqXkyqbk58nwbv9CtPeguU
YjY3eccaFBDMqu0CkLNkpKsZI3dGJ3yZ05lsZRJ83dgZgxVwxXaVdRydxfBgxz6NwUO1o2cjhskQ
9+J9F9t5T5q81aulAL1Ec3/58VQiwZGBG/OyR+18rI3u745m+HXmMcAiSQO1fFT4LoCNpoPMAUh7
jir2GQgXGdga9+FLhHHa6moEGjORHxfy0qVYG4ouyZVGwMvRUMUybYJiSzoiMB04ZdB9osIxRi9B
FMEQ0VQaTqoWj83eBqj88sbxpHqIjhA8yfdPHxIFFMAWU019pdygr6nmUhIw/TVZQwZJhtgO7s0u
sSyDfv2XjafyNdvij27Ueo6YEgfwToUdFQDJzyTCsxXw9CUgHpleFmROTXL5NTOtrL09ZIQfnobb
af74L8sIjgwNXzyI4xd5rtRdR3J7XWbed4ipB898DVvsK8WwQDM8ZOfzZnDzXn6rlzsyy/8OrC0G
nWW+IRzag7apK5OkIkwW8vjmRXqrgJA1AihNQlbQcLK+e/Zz4+ReOHPkyM8Aaq4fmP3KU+60RZr+
xslHX063fxNHCIGuBfqqvGa9ea18226ek92gwT2639dn7F9uOUxwCU9VzB8IT1/tMl6BjRAX/XG2
MiEnf9r83uIZP1UEkF0jctS1kZth6IDavh1nC5S2JbH+6vT8oovVXY1of4Rp76wSHz1bfbqBAufn
j4D4M5NZUcUoDWQe5yPvi+mmA3Zp73lZc7uirR2058t7Fx1wsP9GYUE1Ou+AdDSMwwgkFKR3RDk1
+2tmlzZtcq4oeaIKq7p8yQZ2CmqOtQo7ns9xpOQlkR2062BLUK7zoQLsUMqGvPwzlxwEF5j4Gszw
OO6jsPIhLl2w4BNUmYJ0yelQXLAWRxI3TWUXCTAcXfzyAqb8fbco+yIpLYfQ2x/NE2SEAJfF0MuM
kiOMb2M+oBbSquIsfOnFDhHXFmW2i9qUmT+RJ593YmAP46GkR8924tmsZjZn6Ru3imhCPuGtqG4v
p0s8wSgowg49TTY6wfzt/tD8TH6Ja3udJXcyB8d5t0BbVKa6Vs2cNfGkehNDiqlhYQ6BveDKsAuv
WwJB73Bwjn9N/b58npITzoNcXDbegA1SdSEA0n625KEt7gk3RL5/JfBGDl4I/q61YsTdVY5Cad36
A7BgmxM7MNXfDBhoy7JBqEVIcUf+eUlCkF2jbVkgwsT9Ln05idrf39Cr+uJLC3/lrPOVa4abMkNJ
dbmJV3Fju4YPqztWJ+MBOe12yZydiW3BsqcpHz7nhXAwEqStvYbnQn8i3/jdYrABRCeJQ+RVnhnJ
hHyn+oiySmXwfl3gwD92siMlU8XyRDumifT4dsvWDmAnuPZ0DO2qOwUUw+XUElBcCAnfM9rTxNf/
NHHi0MW3Gqq3wuwdQd6+xi2V7nBs5UlcBWw+G5duTqUzkj7g+c/5eVms/qBGE62ugCOwbh9iuiWD
UCKcGwUpKCaLhD9zTSNQKM0Ed4yQ9OvO64M/mdfhSyVQLZtj4Z8ciYl8Up0oe8TMU5MCfGP62T2C
BKWyyJpOB/wcU8TDe/Wzu/PlXr5IAv0KZC66QM6sh6EIo7hN+g0DmF8uazBr6XC/jsC6Najg5i3e
kQj9l8hZtJU0sadtEeiTuvFtBkxGGdls9bfyKvqMA2fiiQ1MHWsSjxl9ZCogIkFarv6X9bKmCmvl
PSTb8ZbBVfMrUusKtIOuuzlphka6MUiMRFtQ6/DZLDk6xBcTx+5mTcdaHq1Sl9NHM8RolGDMyXEx
Cy79VefCLem34JIRDa6M8JpWKJIK5ZSMmuOHb8viA/BxdK/CJhs/6093AAFoX2D3b84G3qafxwHB
T+UDNQ/RATg82jf7XY3Uz5VYc529TBoE3y/eJkv5/LzGFdK0p6Ze+cj/DNtPpAUlYaJvj0fZStHv
wNOvH1E0xUEbBENR5/HBWClFgsCa63WDnSAyoOKZGlsTyzhNlbadUSUTksPqMOLtr+cfdCwrwsv5
SnVoBUaCN2r/jPYQfH3w0+hSQ12tW/GTxFskDQX7OTxOGhlko1T0QSCS6SUDg+pypJxGl8QG1aaA
U/2b7r0xyWhuuFjCC+9MoDgIlns5OVNwIjJiyGCq2UkoehokC09ph9TzLjldDcanVrEjG9eiLXRm
kBW6aJUqQFmgA01GHQY3vHJn3Xn/hCT8wB7h32Vp7xG1RnUmsrHAvkm5R2naiOzOMB48SBLxxFI/
S+UuETnS2h97z6ov/M6xwHjXkwvTgIuwm8lV/kSOSPOGE1sEmV11EpjROvqetbRo0oiklbJ7zndB
/F6T7ndEM5YWVlm/u8YM8mPRop+oQ6muFReWVeMAH0qDtkp+d0GDgHarF8jrsg9vF66JbCd5slHI
lHMZZeyI8QAmWt1PucUB6nYFcCzqDsERQDh7drCq2fQPcqk6UoHP5daYYqTTKZVN2JVATkb6jwgl
t8qDYqYvMlpnzCV3JGNjN62jB4yJMpT4HksKKv9CoBdu1glR07TDjuq+MWKU7nIBgKPpguJOk95Y
tvyp2c/aZ0M4wrlpV19bgkNNkVSJq7AljwyvEUXj2b8em2nxnaJG7T/kOG0ITmkcsHIsrsUwshfk
ovFzDqoDPsQG/uKBhj16I7QVgd2WHWyWon9+WC35fRERrzXDlzTFXjDvQHIiT+gEmf2H71sxy93f
S35+60EiMp7e1bjUioOGOCnj8d8+YkxqJFmsL2SW7jq/xksP9vkoCmhbNSlxAB62IeK4zgVSXtxv
HiJ5mrCa24I2NlMVOT01xkKo0N1EA0UC1gK4+IU/60BhU2aCaZQPtqrHSaD4MV5L8h5eqkHN9YZc
COV5uxP3+ulSgl4cFRnS6PvsBWeXbX1upP0tUpkf2h3+75NJkr12S0RMh/iiHmx53Ehh9DtsrNWQ
HeTbjDPZXUECbfSHncP6MRKrBvptLmFyN2/qeueFqaNWUqQ2K/biWAz+JYuiqjxK05KhUP2NHFeN
6X5iH6k9P+hhU9gpsHNrnj+kXaBtYrtjrZ2CHxVcx1+zKT8qUgIXyCD6sXRRBWDHvW4DoIwmCBHP
EmwZBRN1sWS4Iga+aZYH5uLfk1dTKnxwNff2JnjXWCJLUeUJOmHxH0PZrVHhIGCMlIO6Sc/si3ot
o2bNH7WS55/yzfR9cAOHhXLdGS4iV28GHoVUqo/WY1Ra2BN5FhPz/BlA+5RlJotLRQha2kwkTQB5
CuQWkNcUD+UGD6VuEwcj9wfw6TpJTEOvKlaSCj7usHPADfGI1VuZP7jiCrSmrJSaxr7RkVJN0COI
wXC1uMmyW0RkApO3aq0pq/VJkUH2nlHklNJhPN0HU8QOfrrhVJKeAiYq3+HgKmelgmv859LxHZFz
OkrDJ1op3BUpagEJfPDVP29j29pYxq/AXEoedlE4wevK01L9HTJNw3jzh/3FCZ8AU0TcONT76MMG
VeAlQlo0+qQIK0XhjV8c2xKjheymCilizQc31+Mw9l89J7/ZcbAxNddhM+COXxs1pCd2jhz9AuI6
+y3lQyXP9kKnDVI86V4LMGwec97ZM4UIERxmOY4rE62FRz2T3Uzu8OOZLRqD30kAFC9NYM1rs5wh
8J4QHvD9aBZK4sFpuT0OHxWetv0uU0EfzmpTbQfnJouECYEz86+Bo2gD16nMWqm93GdTCKf+e3HT
Q5VhvVYAJofhXL7Fd0fL6qkXvjviVU/gZ1DBuPkaGW5ESNCoeI5OTqfuKWdU7mnxp9jXvGPDFCoD
kIyGiLv95aQZoQeWEa7nzIXpx+oDxs/kJ1KDl3z56ipdLCVxySDZ2imgvfAy8mSwfsQACKoonCLA
HpccPZKqAtLYAg3/c9IpJQOQw/7jfBJ3V58mrmyIMgJwRqD8eJw7cK+lXvtW1aFyxptRqvwkg0Zg
BoKzWlUcwbd3pqvvgB8PtQFO8uDwRzKR3KqCqxb+D8rAA7iEmTzT2F40tORKXY7C3vljBJuVgcLp
6+n3NubNlOAOlYfhMqs5ZGMRFavxj0n4jR63uaKfUaIb8L/zeLWELX7xVbB5LM2A/cvH5nPgW87C
6GmanBEI8zd7oIaUe6nRAiH3WDqaZz0O979tkxVAYUk8l0Yq/bGmfKgY1SLy6YHZlH7eQhPvTntM
HFVIjaNwXfGiMpQxws+P44Vy5s4dDVM0/6K+MI3B3ireXoOddvPMPxKRYWMwNhNP4XX9Wls8r+et
yCtb5h7L/EysCWQnyFXNGb19tk3+f5bBWE4kwtVzAac9gJHEWmu0U3To3j/cfniGm58igXClvmhT
iNb81bQOvSOC1ncAiLaH/qw6ucSvBjiNjCQ0R491/WVHs/CfDIjA0+bhVe/Uy6zLgVXJYsFF4qtj
fXb1I90Jlz3xLqc5RE8NbSdtV0c4jKBVahkAkbx25D/5CqgOOO0dx4MRx1h1Myh3Tn7AjQ0nZzyD
cjugWCJY0IvVvlyoDIy6+N2lavwy1D25rJBpc+sVy0hmwMdyNFIv3MyWz6EFSyymYqoxRR9XCbWW
uBz/W3/vS7hXJ2RQQvtQWEb2OAi5TqzQ6E67kIGniL0TI3y7tDjT/8VwWjJK0SJRKQiz6EjbDVxF
nzfDTHgQAafRYThCmPRTAnSWXxCZ/wF5q6A1T3yjKhjYMOdNVsx3ngEdUCCL0IsuQSKmGWqOY0GD
9kSh6FqDf5BXPXd0dlT3xotf3zrm23Zj2JgkOHGtQC48ZjguT3KNt+F6BNqTodIbQSy9YlD8kkJG
M2mPzgqtzn2rn2KjlUzoSYCi5nNCem0VNm8W4N4yO5VyJDurFFmvoK5K1NV7z9Zgx0XAmmThQxla
LTxX3xshExG3IBOmmGXH8V/4dNlfXI4cP4yq7zKYGAPvl1z76LOuu8pOn/uq2Xd9AvprcrTevm/z
S01OhEiYgN5PEbBqEx5KbkhyQgB1k9H7Wig3323qY9gjSXLFRT1/PT3cxMyGhs4rKmORt/UKEUGU
Sm5i3wEGjxuZ6WzxRLNVlJch4iIKa/cu4ng5g+tf5nmFZ+o6j8kPt9Cum2W102MPtjB2o1rRzPL1
S+1OijSIswd8NVe+alhLSAuDYI0xcPeq9VaCI+jGHFgY1gnDl6SAFIvWxBNFUIFdNeu3SwWvtpDI
ux/OithLUwj6JuP7En4qY6XiJKDthr1aooF5/9mlvPDz5Bmo9JHLs3sZMVSKO7ywfhpXi5kU86iP
3tRj2KnA3OP9YKoDT9sWdCSquMa/TCD62J9YV8EQN79zjOnuadeOlBVyCNqvLez6/aSTH6YNjXDH
xpQwIuGwwzNyYQ2zpkWTELSBNX6xY9gTt8WnL5a8JA93AGla3d/bLX/OigDkAVj/mqMTlN+eOmEu
oVB15YUVy0Zi8i8Cb5thaqRefbeR63Gox1ESPR278lOMpAGlWjtFMDO2aLcmKaEOiszHfnXNsM2G
xe5WPfpH3Ywc/whbR2u+KhLtMJnpmECtWCJUtsgSAbtjzS8WepjhLWroZMLXjZaWxNwgglk5/7tU
uBMgAPmHIA2nfGfLeXlYjkNrnQUvRQ5BlF76H0WZXNELYd3vzu7R+BZL4vEMmsokX1LARRqrtn7X
cgGStRIGwOilP+JyfU0H8IN6MeZ8VCQoIzM0IEGDRsBTXlHm/YY3736f9r6e0YHgxigNb4Yq+KII
blpnhWl+dr9gQ9xXOmdYt+nIIat/HPoTeLUxx60gbvQcCqhlaH1jjmusoZYzxdV7/cM1HU1qxq4E
YH2SM1JO0lv3+R3VfSzrovCSNQnKUIh6HAPbqtOLmDcw2tYIVGEAn5KuyX6nZSqc5TK1Cp9G/8Er
UBRALxBKL8DES71QlVCrT1UIOOokohVtIsd/3k7+rGN945kVE66bwqG2YtezaNKbBG+9MDeTKp4F
xpGgp2+fiQKGXSWjldLi2Jq9j57bXSvhd1S03MCB1VFUj+EXfw7hjxifFi1sa+Pu1qtAcZX/RgjE
rAh9OeVkRnPxH5qj5ChUN1XyqOmuQnLtuy9ZR/alP+4W2zf5tmbCPfW9rFNQO2gHi53iCczJhkcF
O48wy81IIXZ5q0R+OG0rlsqoPrMsZjQeCOJnE0VKNwPTo+y5M1HTsWipFJgut9DzAe6DjdjP34hl
UUIUohLSg6r4YGR49XwXHmlXVBXrEigUH8d/34tRMn8fpf8M3DTa7bLEPVgF0ADnlFMFcpxW3f5P
SdJIp04t7V7GLg5DV6TjHrLxFr/XjNBsVjUm/075ETEVnATdAq02cMhb6N+CxlI/sM6+wA9okYwU
5jGTAPm/shpT9sz+xC+B1vaGx9/OLxCW7rD0DpvZOQEwEYlut74s6V5lhIEVHbFv4cnqJ+NuGzdF
U9XFpts9pcvvhPiD83odutLXjRtIWJOfhgJ4doUMAbv16iuwEndLJhfn5/75W/wTxKkn4qPeBjD9
DaXRIW5jVUoI1eFdmBGfeJd3PYOvIJNrvBt6ieptR7rMIpJBvDBwqPwnbn/zIB+C0aWOE0Vj0Kex
7uZeV6WUGNsN9ToE4D9kVca7GZod3oKMTKEqv8Me3fgdRs+aKAHHC6iV3GkqT4BAn3tM+o4RVn+g
vBu/tfcwC0q67P3i1SN/fkMcy4HaYuqrxPAEnfhkfrPGge5w5UsAu6sByEW++074R76QD9MdT6T+
phGhHDdgNM41zQSf68RUBEAASOvdxRfYi3nQAUDziHqryaQqVn5ooI7mbbRbogmvVtstWpuGMcLe
UAraR8gnMeMHfc88zU1mrccEzhHxeqGCSNEUzNpKSurhhLVRDghzmcBmdJ0gyg68N20lxGkPcFIg
2ttMHfsycK96NB4nW3DaJyk+eNJ5WpfOJJdoJ29swF4Dv8UQv0xd/MwdGJ+q7f9blD1uHSPoHwpH
YArL7WXjKSOAfjynyM9sVn+Aa9/ylXn+H2/F/DVhBK7vqIs8x0Al1o2rb8Ea3P/Xdwtu3+RyPpTp
u657fdfic+tcjadt/rGqfntBc7Vr/HnDNjM1FrDE3KFisU6mZXF2TmpFe6+XQugf3uTxUN02F6ke
tDqBsjoK2iDjaCIwUazznShV62Toi3UsuBhDXPAdJr1wuDMN1asWRIHO2yqGcr10rk0SW0S7hJy8
VuhZP1EUr+Q6MwDVOj0/cH1lu81/Wia6j9P5ke2th/qg4CXK7xa8DShttjMyr9YcsYr4ggvUB8SN
OFfy+NJES0p8+9KM4SRKk4Fkwm0xMZGEku+Q2f77QDmkfDvq/fKVbZOQb3aO87lJINn/538VR7sO
u5GHla+/EMd8yYFKX+QJ096bpqkLZjUHRC0y0MIEl/aLV4qTg2C24VqSaO96Bjm9A6XzpPNUJTZE
IcwaUV686beDKJ8FpzAJ6QXo0mvmfYTNyoQjrrinFfEbAZ2POyMHYiU/j5AOt3agPAJO3YDmrDXi
9fIpalMXlJWjWXNEV4PjFThFwIsSG1tD4pClPcjkyX/sZmCbEVtBowoa6bqDAHk1UnubJU0jf7HE
j/tvDga+vdAaJqMwZvK7gC6YJJU1fAK8btT8QxXfP04hzZppUOP5vYObiJ/HKDjFSxHeGl2YAtjj
dWSPRM5aJRQeqi1NXRiTRQTNCWCTRJVxe2bSUlyPxyYJEv1hUVuX1nfAc0BXfvsjvKyajgVtbIZl
QT1W0EvS2d2jylgj1sohTUgako6vdKVuPaqcJCRa6M1dARjb+J0+Qpmn8mODBMGliifjw20YY4ls
c5lz169CnKOhOB4ZS3gjI4XmhfF0tn/V0xcSDwwSlCZ2KTsZe+sIpUtXwwocm40bo2Hd4wqtut1x
PWALQ5nAxjaL/MtHlXgCKsw1uuxmz+h/1Zv4vB9ZbV8MbiFzTbAMBTdSbiqfwi34YnU6/ips8Hkb
jUSU2nX5xsHRyrv8+gAAULHW15O/9H6B5kJfQ3V+I+K7h+cBl0KSP8IJpxzseaEailEvKfz6NJn4
+b5HWWhEuMMPfxiMMmzR4/Zxmvi6OcKj6YGW/WxvTHt48IXNq4pwLo+U2nj859YfuZmAUNUznPla
ThSUuqiMeXs8OlPqoH2sCVo+rGv1RMHISGH3+kux6CuZMDgqceys3/vr3KfG7Vre/d7kHQurWQKL
5sxYhvM9Y7vh5FYXprSuajfNX5lvJjgheqLqjHKKIM6GNP3Rg98nFYMlgIhkPQUFEQRNCbvOpeeV
heuPm8RIToGeAFo4zk+3jMePadDySeptNL9pMDbh1T1iHSA/VG6IMN1O6fn6BO/q014is9PgSGEP
8jHrgofsntFlKP4G7Ri6FvzFL1ME+4aF4Gnck7uWVQa3bUbb07cDsUr95UDoV/jhczoGjxL2rwhy
C10Up6JJ5WdGjbJfGayDqpEc2KDnDqSsC+BwynW9DwaSHQH3ptSiQTItS9FJG4D5wVwxbeyf1FX3
aSQ/f+GGxS1+nhhLrkqe/F+Eiy2QIRQiJMiGtPC9Y7HBBYGD8/efq8aqGKvkVZx2cyYL/7DZDRMd
UUqpviBXcvuZS/4t5wPkFd6KS+7hs54YtfWPFGzD2AM/xQGalfmqf4ypqe0na1se6TC/mQsAqOJ/
mnQMEtyNxUQCrPjeMZy5nPM7qs3VH/VTf1LkiN/64aJPF8VoijM66EaPTIRJqIRMio9AypAmUbP1
hVoRB/mJ3j7evIyyl3IuBnZUeL6kjfi1GRrNMTb+W4PRcsDRmX6468Q01DnceY22aynuwXhFPR34
7mcFK95nGW47oJtsxII5G9xYNRRJIa03Gxjs45LltxaOYkGTQjIPE/pI+GI36WvOzjFqJJJYx2me
msQayWH6sb87pHn6wpck8WMhayjCoosb9r5BQ1qIeAUCyJ7LpK839PyKCQt6Z+O6WvYop2YVqRi9
EvfXfd5zM2Hcps3XtmhBhWDMkfSILd88bT6DeeAtB+76UtvHyy4EZM+Ez3BXXnJlVe/cdZ242XZn
KlkEj/4Yug6b3cXLHrEsoFWAxGMn1xJDx5vcIozEm29LnkrtgoaZjXDVA+/ed5C+1tqB2GVL7219
DbX9yhmvfQ9Py9K4i4T3hrX8e1AIcgSF4fNCu3lbvLGIsD1d+0A6hcpy0d41UmMl/+KROXBBlsTh
VwAk3ZA6XA9gYxeF255M5iZIfpATDPqdVBcoCtEKWweVPDl9KQvN4+JrRMBqVuYfEbZfnl1LEuBa
qhSK8x07G2qcDvCZJxRxGL1cFoFSs2RDxWjiDduM9FJuQXbzwhNfA1ilcwMkXsGtSJCZehliSwUB
T3iDP9JxfWunuhOR2/tG9Mc846zrxinLNNc0z4wMJQynD4zRs0qIpUEFie29bqNNr1AhuHNGEqeH
QYqeUUYZpDqm+XncLWp7nXplY7MwSBOa7dkQnoqM1KXvq4xYSKUTCk+De+q2z9K73WdXkcQz97vK
BAevq+zplvgp8TFOURzTgTbjrw0b4jAQg1b/2NEDE9McMOQ0cSYRwI0kBNwqhdFlWGm79IDU8Oag
9zMyYQELf/C9icWn7nWh2nZvZff6eUwnF6gTb/BAw8Zmw0IARue3X/zNn+d+YTBP81rp/ZsAJUEa
9Obf4G+v9uKW7rmgXoyD3rlCC6IlGG9DqPas+Yd6ObhUoIXEgjCpJs9ghvY0lWn1gIjHssOjIEFq
PEAPY02NAwhSBxRgP73uoomItTh5tpr7eorNy/uDYHEOrxarBUSq+BWq6cmpShF+/chjKGwt16kc
0D2R7RDd/dTX4NIgiIb/TUuyOZTTYrTHWc79DFh6M3Hlz/Xfq4jfWbg50saQWG+n1ms4uBLO9qTz
Hs61kk7x/33O7M2nJhd4U/Xd1L3boSzVmyFBPJdt7tmJYYiESlQNZhsBqKMofgs6pg2jVeMaYWxr
0EtVYroGqnW+7WZLT7Pnzm6FX4yRsCK7yZa7INxP0Euzf63YAEWaP2yrVzOJ8Q+XncGRiipnZ92A
njts3J/Sw4Cd+kBTt4sTzKFjzmhP8+dk3CNQ2zuPY6ExMK861HI2EnzH7Jl1FaHFC/DKN9wBokry
C5rLSnhrfb+kgSReqDMZ2MQ+T7mCIN/heJIZNn4IlsdJBQ+XUYybSkrUa9mXDR2aXfxCqUCTLZlc
dXRgdoCvK0nPKmzdZFDZWNUfD4dz98p1U7NQwG6QUKB9syT/VVEL9MOFgrkw0AU9A+HaJgcj7Cyr
URMRHgSTGTavuW9nHfrDmDu6LnoqO9s4rgPnOFYZRw5Z5q+dmqa+ZsJcpgY9466KF7ng4aVrdSPy
o/4FGOCUkN82PX4UW2Udlif/5lcWgeGP5PBe5vUA1o25O4OUDnpIIwiFSIrR2Rh9A553X/0+GsdM
BL4CR2xMzb5IIjeQxZyfzI9YrAfnpb0zHf941Iz1DhKGGpdES7xBJv6vVBW3M3cVjrkf8OmpoKQh
Fmm5BoYN9f3B5ogEqNeoMJNq9IKvt52USWHmFdk7VzqLAcvSks8+vYFP3Y/IKBNVdQXNGbIR7yRU
aLYmfZtvWTkgs+44AZ5Ppv7rzQxMucP7iRfBDilO3v7K2V0JcHfQVr7KWAh4kGSe9PX5BZ3d/qG3
Ofpzy1qLGLJTC8FtwWOO9mgSEf2v9F+EcEo/FXfYObeRwLejYgN8FqbsPRkoT0OUuINuyUQf6vHT
c5wYZzCpYDMbb7Ehewjx4czEupMrQCBk3T8cVZf2UL+9xCQT7+EXuSg1ZQHE9RyHBdZIpONTNdnW
Oq1HWOdO9+7Mlyp2DOFGF7XSpG+bdqHdoLgc7YpuWMKvgfl0fDLyAsqd17+e5zvyppClMLYT5GSP
PnlG8Oh1OPO0p/7LYX3M5nsTEukwHbeIxOgftqHg/cB5kzb7kj5kF9zvYCmPZozTWWkV/OHv+yln
CraltWpKlV64AL1av8RxpIDxdnDv9gDbvHE5Og2YBZAi5rz4jyHfJOSX8LEiZW8KILkwCYQyq1gD
rzLbY5Mey81u9e+ADiOZmRZobZJ/o6CvaEVTjR9UvNGQj/xsAswixEmIClbaSpls8DVXb4NkiNeb
FC5//SMM7Uw/XqXV+OG+FY2rzxu8qzenI7hsFSB2IWn9zlDfNO8UhbO9U5ATIGKHrM2CPTqjzWOP
PXsZf4QyEyxYOnthvlkaXlK3iLVMbCzkW+d9Td867Ptt+k7ioxs393GKoJOFF73CT0e5oRAhvpYf
Ze7qf5I3ZRL54J4Pkf77YZ2QTJmWnKXJ0HbqcHGWBaY+KbrNAaU+dpxk5AuM4SGYcqWFDY0kEip5
Ilhjjg5NOdAN8yEShCFAE095exWJa8gNJyOWsURpgDWlu2gOHtNMw3nU342PESgUjbP227lcFXXK
DxlLV+pzkjDz2lqYjt+iRF5LFz3Ms5I0kGgJInx1KCahy+TBlJPOe7z2EyN4gumcvm6Me5pG/+tw
2ez2iwYKaz1fpQ1W+83UPEt8tGv/oYgyo5jIG5b/QQ4YH/4IjqW4o1BShtwvGT7SrQMhfGrlD0Ho
VnxsTcsAaDXLM+ijrEC5uhSEuA2xsOyBU6MtEigTpWDCn5uedOscPHQiMzbiQyyzYspz9zdJyCwA
z6cWq1P+slPXWkXZXnKEcY0glY1sPK+pTiawhGsSS233Lycu5VxYFOugrLjEExAvhy32WP6+t6SD
8tZiLHmwYXA7Ex9J1g0DOlI7WMu1gg2OgVVClnc8f1Yja5jjVumT2l7LnQt8VX+XBoBDT/jL2uOr
iBvew3I3ieNXr8xFMNa8bP+JyS2GVm22R0YtAox1dKgYelz0mcQaPA25oRXgXhu7YsprDloTCQYH
tCfQiZ7hRIYN7jHl2RjfAuLRpJsRnlxEpfxZx2tUn6SyxCVZZTj6iahgQu3HEBLRrcW/sx57+EPu
IoGpS/1y0smeTQE/Ooti8uGgOFfOOsg77QQ9vE9mvgdi5PBHpaQWHUBV7LAuNY697hARGUiuvNO4
4wEMwqMpCiXQH0qRP3BZiYKIMAUFJtZ768zrD+t3iJQhvrB8ZKoASQoIiV7m8CgGU1ORpLpEeiBA
ySwdeK7wI3Mcb8UrvhielDM27WCj4KXuZa8o/vCb5Lqw8nza6qBxLtyy++BZTnwnE6c8BsyxQV9s
uRQjxURPqzuPKIUydeZU9N+zjw8x9sweW8MBAoYAh+nUMC6Z3l3hvUmkKn+VFqNg06ZE1pzEqdVM
Ul66bjPxHP8Rqdi7Ucn9VgRy+91Hngl8TZbnKHmCmSJhlHorNeTc/JJ74OXrK+hOcW3HUd5yLMmf
wbFuplAPt1hddEhdutr8vtX7oiDQgwRvH/xaLxnnEcGfjeUFK1SF3G+vQ5LWzReCuFtlZf+sGnEb
6Q2sF8qxTBDz6lhgZd/MTO39TPH9azj7KLuamupwViK3UpNKoZyfuqORj3oOvOrIMxKj2j2Rv/DH
GLW4UgfoUAdFGBDssUaH/tXrxtEqnCR5v1Nu/5MbuC5oYzpCGTacnGtyqazuhfKeY1CVptNWGmV/
cmdbUEMV8AUnI8MEIFNSQvVge3Ueb8zabmBTpS3lg+jY1LioyyVNORknoV97+DQJvnQjvDcN3s02
y9gKvczl4aJHbgdGf9oJqLtS4QxmSYn8TYR/16jsvUd4n/jETZo7iakqqxn5X3T6WXj+5LBILk1x
NMrd2MX4HGUBzOw4fioLBTNMXrRNntMTTdy/vlb9X0vNVJfv/d2erT+8AhARKe6wgBYSyt1Ca8e6
QK0ekVFbuoWn91e1t1dYMs1YnuG9/BIqtzNRHXszug1ILI+9gmqywWr30vxVEYr1rYOO2O0b7cN2
Xzb4vsVTLX8P+hxgVfUQxFSW1nOuLoCClJAas3LpA7RfuyRKtO27g32mEEOgApxIlHrlZjnEl7ri
Vg1v2SYc4Ztm9opFfYE/s/xqUv33zze0qywbduWF6rPufCNeGFHLFfdACk5GxKI5UFlT88iD+Kjd
nMS7bcHTpAOKdH3Sbrj511Jla2z4ew+VSlo1crI5JO0KfrkUQ1OZTRsgUG7IKJO/ces2ODiXqwEG
w1dQAnaOlzMrLcuGVvv/HR0REq8kNrW7pEmFO3mlLaqfwS+xIJxv6HUNoSt3lNj5HtuCEGWJxjF+
E8xAed0kdPd0MOEXtMnxY/rFxcMm6EkmH3qotlSOmZ64NqaPBd7HWUkXRSgVOH0E1GTCufff/RGN
bgWZspcEoQ3olFNi9Pa/0b4JM98NET8KldRmmBdqPoS4d3vJ9Ak2avXFmsx1lowA133CwGLXACpG
5vkw3BL+RNq3flB31MTwdrS9i3qy5Sr18WxF1u6uG0s+UHQLeA5QsaXBj36ZYXBead+jdIzNib3u
plombBqH/o95+ERkKU39Mt/0NQIAkW6Rtc2SzmmUbBS6YNIaAlFBfY1qTnlKQEDOaDgVHVQAgR7g
phdz8LLHh9CkEDkNAffQaq54jLb2we/8KXtxBwiz+RlfE/xjRgLwW7hxYaI4s0Ik2Fv4f3IDoSvs
kTYstgmmiJUcR6PI0CmCfG1tn5l5H4N56YPccwY59Jj7tL38HcbD5LQQcdlFSKPxdz+QS//YeHiA
ha2zKZow+gV98IJ3Cu282T+Ox9JQUBLxVpzbj3OMrt5P55SEleoMAc82Q4VLFVGTvgUEp4Yi8vDF
5UXhOMJVq8DpdDvHCuLiQX84mtZC92lFM9LTFxZEF53o6Ian/xdPjCuTClkbOwQ1hOkGRHhTNehe
6CFT5RDFbmnquQ4mkcA6RgMUmbAm6t6NQA4sOYbMHsCDu+1emG3C1GPZWJ2OszYTJg8wpw6pQIT5
rKvrWGzz4MxfOm8uqH3k60trdr0zB8JXV5xp+iiOSN89kEPb9Sg08hUseucSRMUN8JVf9aztamfA
66k5y1I2eXImTSKxYXwKTqMLWgtNRjqIS+J9n/6YIt5vWGH7COIngyFOQkxW2KG3jbMQ3ILQl5eB
0Yfa5J9sU8aa+rNVezOm5cCRqqngTjL7la2Y04GH/YnnCF3DaLbvoWbMtqKkd1hugmuraFhqS4BB
kSoXmXSqmeRYki+vF43tfOhOfPNAtRLhaG+KVdQueNZW98gMR4QgixxGpLNZLoALWlxtdHMa2oUm
Fx5mJDKGjymiJo7haPd+aE3Se9+Ew6oVgi/HRxxVTC1uHV9vXpo7eHn01PKub1tgsqPN155bK9zX
8Qi1sxjTo/ykAVmx9cMJyGI2EN5fGLT8UtygPXzpby54hSeBMxlZQMdP2QysBfsh2YOHgOIga6Jq
3pFQ+/9hNRM2233HLcjbUcWHjXbkLg88GOS9f4bttO0mP+O0TbVprQBscnvfa+1XhdfaMy58Ui01
X2nsWdQ/LW0jSfNaLwVdSwjpUnyVFNDXsYLIeNHLJIVLeDmSFqNVdvy/h9N7txL7BazWYWuG8pnO
AtcUGY3MEymQYlrPevNLf66XeUXgoB/SBjh2AH4UmSMdgN6ngZ2gTHB3SybZx51WtDq8P8S7hrzx
ixe7iYp+CFxWV/L5vBtn0j2e6Dv4LwPbFMhJ75fNiCqNCXrlzudf8y+rrEliOjekuP5mEZ9xrjCR
7JXgbqLTfbDtLl4efK2/MILK+i/VrpFp2rU9BNSy6eZqoWygcq6pMgk9pCjI377qz54Hf7VHLVFq
ylDhTG/MshmgaGFsUIP5dVLjL47ENIj8/tVLQgW72o5I+Pjn4/zK3wKMi91mZIsAuAvrXRzBMm3S
q32reeaGokgY71ceVtcVW6dQhDHASy6E09oKmKeFSLq5gxdjLUVfWKXBhnvYXhFmtLpfW6kRkAL4
dFB2RbTqC5T6uX2LSsm3/u0B0+EwvhMtjR98VFZKMO6zOAEGuDmAv2KyNL4vE1tYpwVNP5/D8d1L
+xUk4SBpthuLpEi+49KIBEHLkVPIkqdtZDTPke+spYdOc7I9VWJxe5U4Y4K51wzSiX+dY6pfiewX
/mQPV4x6bTAu/cbFZI6teGkFn/mOspWPbqzsYM6wDBdjL5mInqkgWLZJ0Y+RJM4ODkH6S4xO7AuQ
hE10HKiFGtQpV2fVIgpHcbMKQ7GbgtwzlIX0j0GTAn9tex+f/55D3K/weB18OTOkgMUGTqyjPz65
C9Y1bS2FiMM8IxEUhc9LfqFSktqrqCc8SL023gJlVKVJfbj+pJi4djc9x6Z5K50WkmuU4djEgYqk
DFAw8UH/GEDS6yC1maq67y8DRAkJwX/NLb7Dd6NFwp4fyiBsVastGjp5N2Pft91VcI/e0d+anBhE
D+VGCPeC9d653WOHBJUUZ/D9Xot2bSHMrsczPDL/JBhEnYiEPIsJasPvdT7waj3ZLPyjZ7m0jTcL
IifSbTA0GwyR5BpM23k6EBU/i9nhZn9D6b4cIbLBaUvQn7GeHKYaKv9pfQDRQv7xWwVPwm+y1zpu
ziCIlDTAP+EMhrOznBBWA86ngLI1xpYCjF4K77R9V6nL7qXKq7EUsh3SBiVyoL1ppBHcuZxq0rM8
n3DMibshAiKQDUhan5XVSxZ0j5L90byvrIw2lD6Qus/W3n+gYZbgPUQK2v0cFQ2BnLUOa/ZCPBk2
0atLFWMaAWZzj94tCGykb6CMzMGLDcRovaZfYYmtI/AH6Bpcc317rOwQ2+C0YibkU7rvPjW3piat
fZSWXrvg/1YyQqLHvfRcJuRm9pBMtFQzobsqXCzPZeV4fJbhSomtvbdvAVO2EWSTBrSBIiC3vRJE
B9oyOw4fW8d8mtRXScZRX2C20BqjC8op0nccwjpLhDOBG+3ba5/kAvHyMr9B8ORKk6fST/knGTkK
fJjOmAUB/biqz495447hm2gRb+TAxRsQWmteLsiOT/y66+ITCvhBd0JhQqu0dkVDcm7LSCEgubcL
8AmWlhzPPd9BclaDoV+fYIM+EQ1bs38fo3kcHIvu4ulGQsxHmxzpifXlclPGhjHDPLoyaRDAzfqV
bKdRgpXKD1nBJv9x9QQR3Ck7GCUVTR/me7Pu6jbawt7LZP7lXHgUQpG+KM3EBSko935KH25vYdpp
0EWSNVl9axf0oZtLQo/WGYi0OVPCDfoSGiZhH3+7ma/ANeNo6pEZ7jwW8cDSLO4qnRGkylDWhjiE
Tw6ydG5hu7QazRF0/FOgNEFsm6Pz2LSnpHxaQEuIR+Ulh2beLlbLkty/DaFBisIMaCjbCeG3YssF
fIu21PYY/lXy2KntJ8PSIfBjzHpJsoctE3JZOYd+2DOUYxnqLTy5r1VoXZR+Q0v/lJCjc+Rj+NyN
aTzIWLxAmCsbaUbdQdqTKriHbpk4gMi8QyjLIcZfgd88W5CVYaf7KulBEniZjXSbz9M5h+Ss259A
z8Ctc8Y/VUMs775a4IXLUOK3p5tlGE8oCHaK0IwrCcgtGqx8Fz1SF9vnzKpfvoWq/HcxshB9dmFd
LySj4OhIiBkkDTROFQMf3mIZsXWCYBkJc/wRjcI1iDXM2PLIdWeERTPerDim11NOSLdL91cGJCk5
eru3L0r7hEWBs20hnH25X4YfXhAOfNQ5k0K46Lvl8sLOJoZ8dJOdCsOlEFsaXp2aVJZ+mKKWRxmp
Um/tsoMz1DJRa5vF9zGOTH48PSEjXKPtQab7shF/fqCoAdfaidhyYfy4omAspc5C17AECVozQxqi
PJAuGWGR+Gm/Ka/h1Y+fo+PHALYiz+KOG/inOjpA7VMY80uqJdahVZVr5TqHSRGkeuqvPPkP9RG6
0e6L2TQ6+gvxD9OvHEoJ8YA850UZ+GWXJDtL4wo4JRXMV/we1b/EUFrftENRp1HoQ4blY5Y/+gaF
jdCQxha1o+k9qc60IbE/iL+ogPxmxX2yIebO9ohZZcK1NrfLGxgO4QeaxAcZpxHnLoh7orBY5cMe
p2822MXetPlxFPhpYUe7LbMfoOJ+Fy5XqQUSFSxO6ZNSDYzdPRj00WpUWU78FbCksI+CJ4m58Vb/
nTVZacHZSJJL7O9RyZHdkic2Mr4K8fcC2eluvuF6iuQRk+STxL/xHt+WGm1pGatC0UsSTXU0AbtO
L5wSGmGVrIdTXPFBvTmCyicEb/FrrpKbQbV3hLZUQzC+uVoBOUKzc4FJRA3zWDA9vDP3zSU16YYG
5MpSViCuXban6J3kVpE0oWticsD7mpwXjFPN2sbD7NQB1iVZRA/7JJ5y6BQRZ+gmbD1LK5yDRWcK
0Wn9VFGjOCcuwyAEmoHo5IQe6gWyL0l7u6Zjs7cvE+q15+ftVC3AkfAcOWWMHp+a/UTvRNQVsdDC
Ih16hVDMWPtPG7gByc+Ts3S7g/1N+FmQFQDM/aTGz7UlQSGWM7g+SyKKeFF9vEnz63W+hhO3+1zO
sMggTnc/xhbLq68eGFShWRgfp/99nn4lLMrHgdZcZ0rOMWyCJqaPylh/SYFuViKQ7bQKwQfRXbu0
2j7pNqGlJEQdx9YY8yfFasOrmriTNDu6JngZpZ3QUVeno8h7W5ihUpjqeugEoVvgTWAWxR7lrU3u
+wjrh1wP6OGDanEHCFySV05WXQfiAuoByXmtBQDOXt7RntBcH4fvCw7r53CWJbYF7N95v7n4YZLJ
GwFxhukwJZYghOK7+xQ+ar3vxbGLr/USCi4o+3KqugBgvW9/ZlVyy1nkruRLXgooPk+9ihzjtYyF
/yrras2LHIj6UQQkin4dlDZjC4gN6dpI2j57A/t0+gRvWIMSVPBK/JVHgtyj65grC43C2iF4nxPd
+29WUly19Y2yaMxsQt27g5pgXETFudTiWtlIh8qtkqmkY+Xje6/6cPd35LF2XQs1Ty2bJ3QfUpYf
mnNiAVwNOB6Nu/lMmXMwNkc3/omLxEK7cCGp0rciqpCmVRm8ysI7xqZ372I5SRm8s+9i/Lq/Cf4z
Z52yYVGrnxMkWcYB+1wLZErzcYL/vXW34lPNquh7D7VrMKTWid5CIQxFPTZA1ckTBQs6cMCyVYc4
aBRW06z7rvWl3eam5R7I6XjckqvCZlOP3ijKAYTYIw7kEbL8iVaFHBK9W05sHlnl8zz7NdMOXUIf
wcpRZaifRPwsyoAA2c2H5sM9GxF0jJVnjOvEP6fZt6d1dgNDXPXQpA26n2k1jLR2pI3WwyYHv/Mi
7a5IRcqEZQIu/4hXOWcVIx1ycEQJqJ1UhOicUxMfMjmzT/5xqPTUrHfHI34evQ/B9L3pWidkkvAy
DXbhf6kOUqLxppNSFLU81CCzx1ufUlZU0JYWLA8StaFREfXN8aqtz0wq0gewQKtv3tTEMZUcbgMM
Q7ofBvxKvTdMW5l6JbtyTQYC1FsS7TJKDBaYuGbXGgFaUT804lHIn68vjL3x2t/izFXYmDJVuL7p
/UG7L3jS3tz9sf6EuzidR5YvWX0Uk3kF5qvkyrWnpK6Q9S6RqB0P4y0DJ1FJIc9jK50msFxK2pBd
2Tbx4x2fe+uI22ZHy8h3uF0NyD+W9I80G9IaopcqMqoGHKQOoQGWtoXQjT3aJlTrU6P86uUFmVAt
6m+i9Wv67KWHZ4LG5kRNzrZVEaEZt3ZlC5fB/yCHPudvSjDvwXj24RATu+B1Y74aZMs6fH6cOPAm
nVxGrkzxz8tqslB2aquKPIWvisO/lvIE62ww1Stp1lybNMfl8MbFQEw/xAIxgvMiEESb/utyb6LW
NjlQIGC9OIhilpSeWefk1OgnyEiPv5sxeHQn4h5OTd+FXg5lzCNMtPxd5j2uBERhiHGTkJWDIoTm
RQtbqwegkP1/bSF2jWOzQB9Mx5EnJW4YKvWPFH36Mee9PmFD8Sc+5VxGo6do6L5Fx/V1NL7oFzGD
TEfY/Msj0Cr8Mv0tUsSRt81Pt7h1PcJu2E9RYc+sEz9A31g7D1nPf/fPvOOFjDZI8KTe9JhwE+R6
q5VlARuEaiCHxxqp5R1cwbAAJvSz6MaRNGEOUlbbBNoRhCkOaDVwcfHP8YHftKE2++uJSZhCebLS
uM8R3CnbUcf1AleFFx3YohoRBJAQZKkJcT9/7d6PPLXgpwTqLdReJa0w76BpkH949T4NFRY1n5te
ZtxctPBCO7cR50F+nFnDuH6EVWkIwjqzrlKlkVcw6y9UdXBZqLfF592rgAyPuk+ovyjT0oJ7wF+D
0rYo0sqc+6w9crcVVMZ04JeiAfIbz+cy0NXgVS2UrOzL5Z8GoU0sBmSo7uk9mlOhc7hBYe6Qw7nt
Y7r8N//c6gXcJU5FbInYpXDmDP+h+QGeMnV1X6iaTBVB+FKESrfbMIo3Qp0mTUaBnUSX+lIp95uO
/P75ocSYujudu/JoovoYpn5z2lQ3f/yAfmPD738B/PorJkhlXdlkFfSe7DYhPqTX8udwhjYj4LxX
GDkE6gDvZNol0tXompNC3r5WlmfBQK2BC4GmnyohCIuY8bfOot3E6riZZrcF/PF6W/KpW5EdnJjS
ABO2+kjuXWv4Km8cZubjrPTdpB9qtQG1VqJ9uPQ8GwJV6VQ9xpsmsJ7QiPwWSNVm02AmJ2p2y6F7
9PZbRYIP8fF0LHvqzDBEX+Fyf0D8Au9pH/8GTVxhSyVosFVgJZEyuuewLhplB7iJ2osEgQTauYaS
ydrRAI7cPZ38avS8+sp6hEVeLoeLOeLepwUibXTHejuIrvgvVyNzYTnDPgedyhLKCj0VMZO5cZnL
m9GETz+ZIJio9rJQnjmUh96bX4V0Uq8Z1NShPnvu1lRDFse2Cw5w2yK6SAnTYjc9YiIT+XM6/cqi
u4B+AlOdc04VUIpdkztHpcpciljtXDSZvGwzWsazukSNR6RqdRolotbCpcQ7gZz5ei0aw5dbPWSO
rr3va9IXP+1ZDuT55aj8opNtYKMszsJSL8U2m/LUxPGubnhJFEOTXY+exl/hw40B4P3EEq0jlI9R
MxbfGBrWrWD0swK+DPkjUnfLI9qiqJBBdHNHXtcgoBMLYaVYNMnHAvXUOxAPWvCLdr3EveayhBJ/
cP5iXNgLJ+pi0b6utyQ3atCRD/S2g+tDI9Wjhe/5NnfLj6lo57HdjeVY1zXBLPqNi9qmEAqXGmJk
qpnXwpHRpAXbu/4kHq49AzybdZKk5rpfmTIU4/N3i5o3fUdMPFXaM0h5rwZUAihgQtVBir8n0oqk
omoR/tBqgVFKGdHCQIeRPQNoy6BIKPTb0NfNTIOV+kJDTwW6YSpJ9IaHFcwo8iRMPKqQ/GQQmyTD
oauV0/2q6OjeiVm8dfov39S/FgEZeb3GEXgU6e7WJWQVFQJThevsmd0HDCGYl2kxP9z31KqxbZrb
Sa4Bh1KIQ0Gd7vSkUJJS/HziAxcptKS23R5BiyeRY5awU54YijQtEm28QkAPHWtOMZ+f+LC0eGg6
Rm65rXh9IjdcVM0RhhWX43zzUH2qL4Gz6GlVbngM1ePLokzie4xst4bd9XFLUkQyBZhkwAMx5kC5
wGNvIRq8FvfmtMxO85t65h+Xug8sy75t0VCRWuqRKka6Rpw0OeWNbHUR+pC4qiKYeFkctiV7AupV
nn2JXh7ZZal4LiuqAJjnuxhcdlBoqKWngI6tnvKYQ/1D1FnaPn1VfZTDCpSZ25ma79uNycI7DQOQ
0d2ynHq2tm+SefFRmR7Q3zOapWtMB/DAekIR5IAyMXZ1DrF2nkbCALf7iY2bNafSjDAiWOTKcPpz
icwuo3kHDdOCQTn90woLZaVS9763zyeQI8P2zWbweYyCUalpSHO8Gqf3Klm0CLkTrl7gUwEiaseN
gTprZE2N/IWP0lAOJBHd+B+pJAyjrWcjDZB2Y5j/THGNfXXdgncV7ZwaRy+6qBwSITnF221mbHih
meUt4tnFB0VXcnr7fu7FWmHvszNitmPHlMTr4xIPEyXJdYFsGNjBInYb8kmcxlisZnKLi232dgPy
EqldcXA8yp+nPNGkOOIlaWBgciEzRMOvyXc4RK7ofmT5TFo0pWeOQA+slHp+oDTkDxS9mQlXrMTI
OvIQS0VphyEiByfdGZVLpVAXiXE6yjEPc+JQgsvqU2tzLtmFc3SUpVOD0CrqIG7LNgKzDMHsehxS
7mzp8UTNXcBrpaKOR/SW04qsEvonFZCW/ioaATQG9khWryssC+hNuOi02eDuG1+08B6ullU5y6SV
r7/aqoPisiwMglGKJEavNlZCveuRdhx8m+B8VL8Kp2vRBIkT7vNMTMrg0iXiglF0DupDFHUhDpL2
7Q77vRdqv5CsK7TxVuAR1zlCoJTtfp/wtvhA5JrhR4WCbZPr+UeKLxGE8Ql+0YGTVjHE0ZOyIBGm
ad2kP4cHbuL9yq+ABmxkcYwCeVDisnAMqtkneUep3WFs/XmquJilx0/1b3Unu8NT2jqf2fdfm+Qp
QX1dwdNqK0UXjq1GzkTIde6EJO4QbjTEZrYxDjBw0HJCm8DZYeuURZKGuWZ/j0h+skanaxhjAw2w
kfghBtsMrnAcXDq7hhzlgEK8GAHZLfXppi5SEVr1ZhE810/VrKVw1ePQM7hyxZwqQIxrjQqg8Y64
B+zdsyT0IsNKabVwDcIjBQa8rB9WMos6LDH6V98MHQO2pZzK4/Lfl98Y29J+pCTgAH0ZXEpv4hJn
ebypW7a9Ogrl2j52djoCqM38+jefZJK1jfW1H/pePSKdDsaXB83rpKw1KLisFSlob1yaqMVRWrVF
vgLl3rX8zUwZhUQYBis62P69hg1LSbVFNGYOmCOV331avOwfsuJZfkHhnXf3YoRIrPhwlipifWif
aykGmiudujwUOBJhp7O8Fbt5ZyvF48/eorZaJ1Uj8Xq5bUbhfWidDeBK+IgAyrHeZ0AFiuOQOD2A
ud777XUMoDCe2ZJoe69EhXV/txpScEbzcDt+syGhCw6jJXHko05YcOERjxd6CXiLPS3fkA33PNGl
fyATq2W6s7cM2mowVTDADHf5X+fWFKVnOOIH9OKC2COCfAMAr6Dn5TEp2XOgAcMKAD0l0ISHb++v
K6ClmMr31ytubVKSMRYIOYGTPC+FldUNRv2Co4CwYMddrlFAh64ICpc643f/ZeJF9R2fqNRlUvPn
DCM0OBgQPCcmi7BylwH+IAGl9DcG26qF/zuElFz8p00ngljqSIx5TcwbcjpTTbkSw/X+2bDJnTL3
bNUnyaWbNux9F9cLXN8LG6mPj7biNvzSuEHCBstz1WuhljBzKv2zVkQtYqqM6arvdgBhxLhnOqp7
VSgKqEuXgQg2dPcUTMesx4GCK7pbLl+SsokcQkFDBKF464WelMBdq3QH7PXOT5UIkROIg0PnZaDH
TJIJAoNC0vngd2ozLIdlygJJdJi/PYx3xxJIGgvxxXL1DtmN+nyBPkxKolyF6Dq2kRzGbcAIU+Wj
cjKheqLM6MWyJZ9xRg6nh4AJ4bs8tI7ABgYNm5cZBvwwKicH1v6cO6N34N5S6nrixkg2AvytlQL4
9+ihdrZZQ2O5FyvBpX/0SU3/4x1XuoIft8bZc8pX08XJEHSrPVej0Vvym7BA40mxIWN1U6kuY+ud
KOUh6/F4gDG07zfxA+gBMDb+lxw41ZZQ9slJO/pShBhdydQ5yiLgaRZS5pigNLgSPRE143WfxoJi
pdj5RFm/0Os8ou25Gq9GLQ8sUxOa2KV2pfLDcSHuGLW7Ske4SOuiaM4JivM8b75Ih71X7hmW+dFg
KocY/Of9a8Bf7G9adUFybo/aeREj0mUhdNnVhh1fnkLb4vvpLBmC/JjoiUCGMSiOaN7Ihqma6+Af
tNAoNBy3uCtfHaKXcpqyEO3rQrCNwiB+dL+gfRNgROy7TT0tNnc++2qmXk93JrYs82LBK+uGT3fu
R9CM0EvmUuYfG6B4P1N4++1aAiQIxvl5UGOZdxhkfDK8GDariY5pTmXtW+fh/kXCTFLS2GI7Irbt
VwETcdfNDtSUOlGkEdswrsuTwn289t+IuOStB5+bQCZgvvsSm5B3+MZJ2lX96KA59WpsJ+5ZmWmJ
40skPONNeBMt6SqKSS5NBV9/Tgh7JRhhZlfd5xaM7I8X/pUmB/ZuuuBgXFIz3LITxyUqQsqpQ9cX
TjpFF5cZ62oKtLYnZZZ4+giKBE9VMKz7CP7ojeNsj26QVerrY3ueHHBiHkd8JmN1JGL01hD485pW
ptO35lfMvgSyx4ynF6GDniaz1h3iBPn2tcor1fOsPd5AjlOdilEAIfLStop8vGamdQd8Jgr5Hqb0
79lYIGRoodtdBVPrNeP6YiPX7rPdAreG0mPl2Hg4+6wMfLx+nSi8G6mxpRN8bSJZXUhx1LuhSv4u
Gd1sbegBduFHI7NBuhcZilQBqO3cHPRjVDuDm4EV0f3D+JAgf/HOFejHcnvoj+5C3pqNSYLYmGNu
XpfVTvmXyUESm2LvFhLC7KHDkoixbkRCECiYuGXc/kfOgTB8dLinYQoL9AHg2cTNjR/Cmse6eE25
kJgnmADhTVD7cmDte3S6AoohndkwNWen3d9Iy5njpZ5peLTqrpmxAbeoBkKQLPAsepc8fBNZ5/h1
+w+qBJi/zndmGDBdQIyCJQbPYssVsKLKgeM0TTYN/5P4RM1bOamYb1NytWB1wEve9CBj185MeXOI
u4vHPrnqDG57dml430rG17u57yjRHUWpl8ky9wgm9TqhguIqYRKyGq/zhZS0gN43H5Aw2YiMivtx
uYKbuVJrEqBi67/cXDWmWeXS1d+knt7knDABw7TJmOqvAMOFOnf173Dk0WKZwwL/q2HX6oWod2Kw
KusvQvzB2qn91n7HhQjbybUwU1/HQEzVIL9VH8GbCECt2IWe7+QCoMNriFeOcKxjCUHZXkeJUDZF
wLtvKb7amDFJheFns05LqpSs34VAh9Prctrf54B6bg59PCJ5JW/ms26lnpwmV3Xk4d0rDnmCot9f
C0OSTaMaES6++UGq9SE1AK4+kb28y1OqqQIZaFE/MJFVzGZQ36L+HOsAW+YF3PFHo29V1sgO4ZAi
xZNO9rzjSSiSqXyHljsZtwwCOfxuUX4DZQb+DljqdvdrBalmOcYJrJC90zoOzRlsZ83rYWAFN5qT
tqBbwwZ3/JaEexuj/X/Xd+/7pAlv/ZXOsIcPsmUB95eBf/4UKviw052t9faRjZdvcsjgL8gVs5/c
+ZOk4Aj9UlbVUUuhcMU1XWvtaLq+MiapUGbUoWI0bmtjHgP64rceeVgCLFn4/UgcrGAyLXQ0RUw0
kQ5zN6ppQqsxsrije87LIf/p1KecVnsjFHutSn66JfsIp8R5irVfp2reQvJA+dgSmAu7m7JmX7ME
NieqOHJc4n5iid3QzBawhGVgEwC8eeOxkLb8zKX5K2XzAhutkoKSRDbceFRvo3hF1VOpc3Wm+zFA
z6u1286j8gCiOLVvc7WLjOx/k1bAGNKEhJ07rzFYXt70aJURWpOkrAUVgi7aIKZM3ACUqo6OQkLS
FZmARl9YkyCytEkMortL0asRhHNSko8GUZ9jsB7j9oCTuRXV8mx2BOPhb+URiJ037GPJqJu5EDm5
ows1f5PEVt3RpZU/A8q2qQH01jNs2RwuVWnwt8EAJVePbt8w5A3qiAY+F1M63g43ABF7pkQ46RZ1
Qj9in9MIbatVzzwHwfye1lTXkgWkosqqGEj0kWBzRQymB0hCwS5SbM4lHUD2O9bte3uxcTenr9Tf
S6FWUMgV9xnQwv92V7mFiEzqy0KtG8E2Vc+zhx8dkr+pXCwkbeO/hBXGfJC/Ki63IMGodUbXnZC/
mBOlMRi3pJfZFtAfsVc8UKHB8Eu5cK+8W+r3lf9YKssdZXB3FQ2ilTKNEqEaIw1lDB0bkvafFN+d
O2gN43rsxnfUt3rLFHVibT1qGkUoVKV7GWISkej22OWm0kNZzSy/M65eiR1Q88o191eTshfUCAaS
qGGhz9b+qILl/+XyMWpmShNza3YPXFPwcjVbPqrxs9HYkTxvbBakU0gaMBbI/1eabeuxQkbO3roY
AFqRCZYhasj5LLGXrzit3a8B/3KpqdQmPeygeJPGjkrYyAKXZpHoQ0oapryp/HII+Ez5K022+1qc
/Jz9F7xMkgRcBDxA+6dPe7mfnviyhr4pZJwHz5EbwPzMQ0kg7GO9V2cCk7daM/BYC5hK8yRnQJ+0
pdnx5c9tlJ6gMnTeUWZZAN7VENgABNdrMbTe5tzv1JeKh+hadb03I/LOPC6myfffF1GX31m/IvRw
Adcuxz5jUlMjsZ2h7qaHSJtlIWoTEKC1U4m+QleWarkiYaO8apbLtWxEfeXO+44n32uyhTlkY/Ju
++HUHlDJm7burW6UAWdY5ASyB3CTTsVabsIcGFceNyMS/s0XQquG1MKIZn9Zd5GmwW2CO6OKbxBA
C6HglWqyiuQg5KEMlXl5neLXVX9M08TFq8viwKb24V6468sfkyDO7uzOjk3KmeC6B4Uv2zX240b3
gSkOotYN5kSOWRl0x63V0Vj1KfREB5BhLVvxdBnywCWeYL7utxK07Nl9xJ5XLobbXuhdhK5CfwtP
AfZPvzBm3KlBVM3jjxEyubmXrAylTenvuyyy0xSvm+vcajAtu1bZSz9QMuLRjpuJU2JwjxjEi5uJ
2PnnjZRmecx03WN2rPTAP7J43Gqbk6eE+IeWKj7np+Wvb9+uTcD9scFz9yd90i7Y/NlqtnslnT7I
4JYiLYKxRMWgJXk20vvvej9LJrkzI4I4Po+xH9FIGfNrTV8Rx+DlsDRXSYbf9tkuOY8ETk5+hkcP
cnjFw64CGG1thdXqSxhSCBUtDkPuaLu4Nev8JTSkorLO1nZIvibYUhUx0w3frgpo0V+LOTAkJeuE
P8DfdENlNs+oCb3QNPIpNBSbHHWYw57UE5I00+QwEKr6RDnLNpCGdaoeSAYkEt6Q0LNjnVEcOLKU
4jQplydr4mXRRBvnaUA8Dd7utvAOYo8+HWX8ZIzSmuZanYc03cDilH6KILKc9xjAzlt+eDV8R0ol
5KqCKUrnIkbaAKqpKXuUHAoFCCK1tC3PPRFZJtUrWPQoQTkSrXCw4j6hGzNyx4F6rx3kBCYDiQ/I
5BF/iO6JJvWgr8aqe9QotSVk2VhDCujC/uNB2dPPk0sEYGwxm7T7Kwc8hg8O3TGZbw1O+PtEeXMJ
sDElp7vBx2tzPBH4c4FRrDmhL8AJkfI6AuD06VXV4chpfwdAGug+oRyF+iavpGLEdou2jNF0h2T5
N5cGSjsauhNwtGSI4mfK3zxKeI7LduDY8uA69UWcmSBR8upu4su/Vf0zdLFKVoOb8u4IMz+N3472
KeJ0I3gf1vAtRCucPgiy1lI0Wzx1clZXTHdLhqIZHDOiPd7KXovux2xit7bvTOrr+teVYdfZllZB
FuvlBs6FNZDZe6qaeSOg+CzUQFgkrCoJhxpjk4TN09wIfMFKNTitQmaqdRypzRnXWNbvm6cKuuQ+
qSpytfyEzoNITLtryqx5ywEpz4deSSvpix+ajIyzzwoiPi6xE/PjxNmB2bIgb2jgmvCaU6rMoPc+
0kp+dpEQHcQJenH0ZeVjxwoEw4x/Gn7H7bOGllPHpe515D1DAnPy+C9kMibJO9NdEndjCbdjcemA
KV05XOYz2qG7cflifVzyBLLjilnJc6ewI+KUlOpKYFfoY6DXQ0vobZedrHv5neKvSq/gOA497nTm
NHLWZ+BgQXd/fd6uSY0xSIA/PiqqA8SsYFIjZ3cMqA6H9jgX5qdYLSdmxXoRWW6qP77zn4jtLHzX
ij0fYmcZQ3o53dMrZ9O+sr6OPt2g089lJlNMZbAGaQ16JpYmwqpYWKzpv2Px7ofJlLbk7RSLNpjT
LORcuLOLX1VmV5tQABUN1X2O4PmvwoeVam+fnJlIdgj0I4brCeNO82LZxHekXOcGNgYvglCEINHO
kJ70cNRY9vsG0WgsDI0IZr5twoQMVaACpM88SeH/hobg0Xpupo6u9bUg7+A1hgnEJgKl0cInHIPp
+oDsMaEgr4UsFuZsza+2/9Wh/fdJG2xj+q/WX7GoZnEMlGC3eEeAFk0Y3ZnMLKMtXTgKSkyqv4Bq
T/VsIJINEsmMCy13+1TnMacsUMaFOtNjZ1SHraQ6UVWgDpEUXhSHXZ9Ro1avwy6rNf0QcBj9a5Lh
UyFrVqBDSvpZCtOdd4bo4kYVa1L6fG46iAdUwJzXCDpr5H8IbGLAESCSwVLtuNo0gzuNHarIbdTF
XALBWOuH/SmwbYZnmZAe71G5hEeQSck065pSJpeuHR+6fuUiCcr+qyJGZXvwpY79MZ2YuQuF/uOS
oCwt2wKXnGTKc+NvivtdPjbUkBto9QN6XJ30RMlh39uD9d/fdXH/NRe248oav8xeaXW1uImtg3oW
xhyB6ktNu2IALTC8eLW4nDhrb4V743nbxi47Aj2CnuNVJUwF/hWBE5k+tWKnPXWi6lmpaZTRqIfo
WtRNdD1tiwHKu2CBF0u+1wbAxFUNxbt15IFOiUhdBp6H462XkljD1wXslFRVlP/+n5BcTEl2nBpf
hrix2ByJqBT7782HPJGPkzW0gTfUTjajHBfg9HomVzI2caaqumq47NK+XJAfYw3EL3Xe1SfuFkIY
IeQ0PhZRABSTdPhqSHwJyMGnOs32k/H/L2bviw1HnaejTLq1BATX2RiLKhaleKyzP0bL/IaLGrC5
Gtvv2Q9ovWzwKSdjnGefG0LcKC5V1PsYDCWoN/WRdtj2iHw3VnaeBYdqwhBCDZdD4YTv2fhWBwWM
iwJCW1Uxtyx60n8SOgtYSf0YkNCcPIaZgPfavQXSBPOxqDj0ESOxB2I59b1Dec2GsaB4KgMmZLSG
Lhsw/IE96pgbyW9qdAbzZs+dgF1nousr/vY7sluFrs8P5nlFpHDh0vJTuRJbuZ4sAY2qcS730sqI
Ce/b/zcedco+P23n/SRfxIbB1oBvet/Czgl4Mt8Lzjsj6D0VxusHFuKR3FJoi9SbbaKag/Wxftpi
VXvkPK5LpQrZCsK/4GZhJ/kg9Dfua/eWaTTs4bQjTThiuGHc+hOe16wGoSgCRsEUYxvkePjgxlXh
Xbv57Qgny4glLZlDzERDZ1+S8UbksxaXE3SzDcSY6sWEf9uwrfDmeNUwgcAMHVnYSFvnEgLECKLL
Fh2bChUfpNpfDwm5lOU/4+0eidR6pfQbSjjf0NL07MDWretvtk9uNvwTc2PqqBaVHgV+A5Dc1Q1D
FKzuqNcVnIb/j2FiGzuvgtjGaMNEOtKNe7tgGeG9h/gZ0ibe8JtFtwtWSghUV7lN+alNbeLZ5UN/
XxDqMOA2O00qKKl72zwisJqDg5R1dQNRO3z6OUU/PNHtQCDYkzBBntTsV4tA9T11ppTV4dQNSEhX
G6WOOtm+FhXiZXNHrG3q4WNtXqWFxyRZQLRwINJ4uJM2NTo8CGSDGQ63A78Ku2037CW47SWvwCP9
obtRhM8Y2mdXtOzAd2/5ZTam/tKRMf87p4stTzAyyUe3pEkkQfXsr+Eq9nUrUzDD8cG955a29sf8
W2YpE9f2qKKcmy/RSUhc/1Mi5eeykug2c3JBSBOUkZ3bf4aXT6Yo2lYtdB+wUwMHZlrjennphm5r
YG/wPp0Zs1U3dwxNBACoBgacbEM5VEmFN1Pq4r6Tk9smNdP+9S9IvWN+J/lnV8/hF8OnTooHVGdQ
TfL7jLQxjp7Zp8YR+jxd6YJ4Hj7XiX2ZjOr87yE65hnmPZkzswxqwb1IwK55UPej5HeP8573C7F9
PgSrRDPr/MrbO+iyUUEEgPl8A1gkh7BtJEIaJdEBAf5dxQJ9/HC1mkesvio1xqPeZwLsm71pJurR
B2GRIxmfqumyMxKNjfKdmCPmBOPSMdc7FitIkNZVrNxODSFLrwqNY3EvTwGLuNTCAcJGXoDV296a
oq8PxDM/EkvbTFr69Ybwa/7c8geO6jgMwhp0E21zs6YhcCFa8AAsVxtI8l4x8r1IwBigJUG8lZP/
Hiy8f8OJvoBbWPoxHyu4L+m6ZWAmITXcHlKeB2ohFzS0MpPdf++91AejI5s/PxRqDHJLrBO0JOQG
Jj5KXCCye+lwtKKlPBWWyy8cuFme97kMKNK/djGkppN0vR4KAQ24Xqh5LkjWx4kvTmK7abrou/wP
2QmT8Y20fwAvr+vWuy8mpHKzVqqCbzS76j06aNhsOiOuWH/9y7k5JvhtJ/16RO362lM7WN91ccFa
HTIaaD9WR1x8aF7uq4CelH5s6sn0tpTl6hWeQA9d+ei0G3TtE3K7B91sAjTx9S2+Zta5bqUKbwWX
W8Gjf2jRUJdN1oClB/EsPSeKiyW+crpwx3Lcd0NLb0HmshGjfiwYnACpCNc8suUnYLRcIuNqG23R
mHPjOEK2DsJmnDL7EiG9QZlUIFlEgCXD40AwvZNNkp/rhtR63FK+HANjLmpRV9lb3OyrvEnpQGHB
p5jSyGAwWFGp6q/ZQSUJmxSslLr+i9RU8kDZpDXRsYYIpZiWaUL/TBK5Wg8hufq6T16F6QmSHLXv
2PkCOCE1t9sGZHMYb/N/LBAqa3wdjN1MtgUufC/xIM9ARb/h1Kf7TjIWkqjQ//N2LCpfblLeidMq
0Xo+wWjP/pBKHvptGHxKAh2GQ3w/g1UYEFZ9BQL70TuPezFF2YSTdxzZtUExOZ3088ou1ctxWsGT
CazdlFYfHoni1joFQBUatdXipZTfHbWFQBe5TBDdXHbG25NBmlTsAJ1V1SuqVzc7ztIRAtoGQA6Q
k8kgeqcv6dAcF6Wb+Ap/cRUUmtmMp1/nNrNnt0jCcJQQ171QWYXNRZgLC6U1Duzij8n2lUS+P4Jb
pRgvqocJ8gC5J+KtQxteJ6UvRzJ9SDG1CKbmbiQpaFxMoiqU4+GMK0endHZhhvceFMslWBvCtipt
kxga4ReqEYa3siic7352Qw1mHPSjPPd40NH378xQNTM19B/ifq1qbA8thPLNMkWqFwodDSgix8J8
7pCNLjIF/nbjULEKBFnuVfKlku5ESqtjVNwNV95vnvAe+bZNUWGbn5VaT6wmJklP4sxLzrFCRfk1
HoRHOHjcf1UPxdZj3nYQDr07RxlUEoqTARlCewkRj631xl1LpenzyqpqURQhvTMSxKkM73Rgv9Z/
+RYWdV6kIQfEkhGYoD0suTxtUB6nBP8qlsr1jnzFrjccI2ZWiA4r1Nd90MRNF1HqSHlPtcCMKwkm
LnJjc4NspHPVQ6txIw5CbYd7+P4b17+wp/QBJQ4fwzTpqfFipnPePwjZMRdNe/fLjNFEpnXIOiCi
VDEnftzrYAUKjzrGmDGChR0+YIZ1fgYlW0lhLRBVfeNcCH8RcEYG+xg192h1xwu2D3JMVfZbGXEg
Rh9BY4olSzeyhKcCpsgczLe0MXXuLCt78Li9/lGP4ajzAWKfAQPqZk0Z5H4Qu6BTDGbPLz/mxtQO
5lSgfj4CxcPmMljzcTcC0YM98nzuVrT0i0LGsSq42kEiu1RKz0q/p7qcaGVxKBne/5fKRfC9ek49
OD+fu/2ZMEepQ/utR94Mn+wfWD3TLOKu4VFyYU/fpuJC5L1OQmBr5bOW0H7lsWg9rlQb7tcPYnTz
h/blWiAI6/Exi32RmvbKjPXXfD4ucl67S25xbsix0vTMuoXglcwj7Hz9giZ7YkmUXiQKm9rPgEw5
4AqVuAT8LPwIPLlwmGhui/atJDOCSM2VpVjh647jfdoZPCpOBn2ueMbiYjxbKc2l4jHN0Yzx8FiF
IRz9eOPSmPoOlWv60YkxGSzKHBSbxwCinlKgr3WHNDPBN4S+xXH6rQM2GAiVAEgWi7rajScn7fpE
9WIJxutVBv+Vkx9wCZELM2zF419FJxjYBfD7f2JLXScDuMG6OYslKpYPAYGSZ7Jmx1IHw69qQTKD
R5Tvb+b5HtBkTJTwNxb2Be7qBO2tkgZ9a9+kH/5HzUi2gG9JPoqQtk9dCqBivsq61PXawNCFIy7L
Pkq4bgm5E9EWRi05t2s+1F+vIB7sFaoBrjWR6H7leZqPqf5HXYJdU0Zhy6aQr/4PvnrnU7Oc7JGS
xPVsKOSeOlQlrCAJ2rdYj6hVTPllVfhKX9hKwWdKAFuC3GvgskKsViCQck8RTPshdg+9CRKLz0pH
58ELKMwL1U0x6T9N+CIT1GJitReRvPz5YvBStXQyQFHiT1YiAaWpQaUfBPvtlkvC556/Y4V40VVP
20bsfaPbUTK4oe2i37jzTUGSpQ1v4NxRHZyqZMf8mPpzuacKfrDc70tPVlG2C4A1qi2j5adMmrAp
aKHjOQXwInJRg1B10xGomaHQCc02OZPNasfatXb573rPBlMiGk11WGu0BUBYKQHSMO3clTlREHKN
2T246jStsslBclA7rByavM54eZF+vB3IK7iWlQOfxkglEoIpJHnKcdqN/KkGj79hdRc1AevM/Efx
mEam8lJ2cOhwQOznOqrYqHnK7moTYLNKPCZqmBAncaffQyI1vVOCrMG38xqIJ5s19HNBO0GuVDdM
iDzWth8T0IgB2C5ixoN2OfIz362nbOvF5k/+3+F1FAAjmFfcOEIJmjzI7IgJC3mFvnLMdLOTO1zk
hCEe3RAl87mJHhG7uSPnsuPGvyDbxBRqte94hP4Y++dxabhJihx7zE/XKaKXagKpy9rK80/ym+s5
j4za245aQtLzlLVyXwmazLMX8nMM0GBH4Lb0Zpslg9CSOD4GYN6ZcRMnoc1ba3fTuc0DbFftsS2z
/GWB+GP3Q8xe4LPqMx/s5E38EaK4F7ffRuOQVBdOeNs3VB1BvJ60bf7j9uGurtiiY2OB9i5DrSnI
vfMiPQEMqMpYekhx4q3VxV/6nMXHVRgJRvTIdJX1eSgU1GI+krs1DurPs5wga+3TeooRTj0iI1gI
zUJWEArimCb4+/Rq0jIobj4pbWX1V1n2TpimiW6Kx+XnjDnVkkJo0YKo0On9LzkCxJTtbyX5YZ3l
0TtuIAjGq6Lx7sM30anbqJwHthen4obHNKEARifJf7SNApcPyH16/AAMZh3cWPejIh3uGohZgjJ+
ArCKEMnVIcaaNOPV9xgp1KDNkoQE9CnifUGBbZMkKt6yScvaZUVjIG16dh6GDwKRjNhCRpEIg8u4
XA624Wzev/40wcnS4iRud6J32yVJ6zM1MJeoZTjz0VIWt9M/F+gqNuLp78ADKyuXON9ggke/h2yZ
mpEydEdr7clXtuZr5hW0YhSxmfOpWlh83EfO62dqlBlQ2pWtunPNk2lDkzbgpm+avcpygjt+LwoU
ftLk+iVXoE6UGfYRxVXEFYZ3Yk9/3RYAEJgnP37ZNXAPMRZ9zRFFWD/8j/fyRLmm2GM6J3LkkFkh
fhUrW/6JhGYU8hKL39J+9CPlitR0AARD+OfXLHNGyQuqmjFUEyikii50uamyi1Gm0Yw74yxYmw0b
OGBdfrOXlIj+0vfqNKANZTBIiih3DPcT/1dErbasHqDOHQC/L7xh9pFbppJWc9PjsUoth9VBG4B8
XRyCUW8FgaBQuPReWtgI/ci79X0O1EqvV3/Nse7H4wH9snctX2KTKReeKHRGFsxe68kIP+LcEYF7
yWmynrszomnonyUjsl0/SVPMus9NgiFIBaYl1M2T4uLJFIcY+I8tf+SR5X5xtVhcueQeZOKQqLuA
J1Nu82WYbfxdvSWs1gA3rXgeGB7iXI6ieU545iHj43c1YujUbetq+MTBTHvQ84aMnerfa81vt8W2
jzAgHiTFDBwyE5TMUliHlajdsEqpCsrxGrp44bq1q0/IO+C0MtxKY6EV9eCrwFQghEoMow8pUGaW
r8NfaPOLRMejo9b2Du6uTCtkilVz2hhWvvoxWcDUgmxnFD0aYtGCTe0z81yLtCsC9mYp0LIP2Xwb
PZhSlAnzt4R1sPXntGWxXeiI1GYckbv+ypo7Ps8PnswsjX/TJjuvA32JlOBfYWcQgyMdB3jomepZ
R1bFakGrdyp/j/J4m9k5fDVzcjT8a/kdkQmJLOVFHjkdJ3o526qSIJBdYrMfNnL9c9P/0s3Pm41D
89Ra5JU7VQkUfm9xiTPdMsEoEUDmtQP2HhL4a7xde5mGn4+/XfYWmklKdkXw/3z0akMNTfsYRJNc
JrVntv+48Hk4VHKK0Cyb/WVU+EjZ6+YpeDbbVYCk/6/3hLMPRoOb+FDj1zkabQu2+T6QqkVlhLF4
RukbCugW06iciLd7f/rnfzBJsGiA52A/GuHcFQieJTxiF7E08Wl7tlN8UHGHwrCiBr2M1Wyz2I3j
Cqg1aABkjK2D9se+Pw16gigOmwk4dZP/Kd/wqldcKGyqkI9Z31jDg2R6cOW56tOx4SYzQISIApi6
HqKEUx6KJuD0rrvaYGQ1or29UuSpXvDq3yY3SOpk/cdpkc+eojMp3iXjNiOSLmxhBxMWmyjh6A4B
h4kFN+fD8VQu+YEWYEcmhWG6XP1qcG4qDLS6DqA40HWOOVYNN3L2augGl04Mxr4ibTVe1ZuDLen0
+53ZWR84Ox5C3B5O01czU+N0SmbSePP/BJ3y8dupXEv+X9sSRiPK5tpWDqfVJX41/apMftdFdMxx
w/gL9s310rOj9vNmyXnvt2HMqwJpGAtxPp1Tk0AwiDNvoHb+DFCv3b8FmI0rRiY/s27N+Sj1+Iwd
JL7l75CJwHumtS2g55uSlQ0QWJmL8xybxMSsthwPLLkMRnGgnbIA2rEkXxy4lbmM7AZAG+ihTuZd
AB1HeRNrZZxhR92GwkKz9Y9yqkAD8yceclumXpjEF3m0DQAS54GKas0d6T+BI0347vqnEi3lQskO
bFOClTt9O/F5tB/CcokATe/onZm2Jc89Omaxh6BvxqHyl6AC3nhtq7pZiy4GTWBFotBdxe50E35R
OdfoTwXD+w+3cGSGCkUQgST2nUHbIOgg66IUiCdkQtnk9UchpM2xgIqPwoAmuzfRO27aI353Yixl
L/uswovekBwzxVaNZz3F/CGGhYVt/Zk3DODQfYX0hWap5vLO69fSSJMW0ndZC7jSOBBidHGXGjQe
tPkcXIilJ606qasFxJwhHsgJl7mVXySe1ZExrbhh0gm7ea2jv3oUo6n70eFysBZq7j42Ceh2xGUG
5WQIF7c6Q2Kc249QO5UBDEf6IjEJ5lYBx8O0LiB/eGEonLL4/PmDX0z2/n7a0OVL/2HvF+iJ9LaL
km3udutE1pZHCoxa+Qn1Gu3IG4tqwO+asrXy8DLslfp1gakyzHrygiCL/2oivIdmSdFIpCojW8pm
kGgxnAcUS0lYwcKKy+TkNPc+3XASc/gEVfFEvpSWaG0LtndkSxrx31g0rDkZjchZV5YZJFV/x0q8
wnxD3UwRaLdUftMUCH4r5HvHtwcZhSwYbm9mCWOPt8GJF4LwCsiyKgXpA2Cwl3PQ5afqULfxDAK8
uK9Yi2hj1t/axMn2h85wfq6U4dF9upq7zyD6Pdr3zMbRmSwBVZlxm1qUqnn6OrIyrIPZG1oe6CkE
DNsWaKFEFQJlwAawUOzkXEsxHw7LDHDTA8/Ym2rVN0tVraezEvu5dVlUfKdcBDhHFNitpmOVanYf
oepa+7wnw0WiXNDkkArV2rrkguFvvoFSrAmtFR7UYhouaMTWQ0c+p1Fn1RdVXhz2QPeLLWPvnfUE
IxAd5FgdLiu9WZIoRYMDd/1YKQJW+LcOdZtQMct0ifuK2a9KBAMn1cA0h7xLnJ0mtClsIFrt1Qz7
T3oUC4B6mB/p6zWeTPDoXg0/hdpejBFxAdQDJuktqu6R/2Fq5LK07r/1o+EGKz4XV8yu/T9HjAjk
ygFglr/MXsyrnw4Kp4AmQy7Z/FQqlu59k+aijN1kAQu9Dxj1ZQrf0NOBG642pFupBdO77DuJqxOr
TDJ4vp+qN2MsImeqP5mTdN9zjrYKPYLuB4x2Kw224Cz/BNw2AjAds0tPwg/K/B54FjaKRMqhGGcp
0itagk5Aqc5AKaoPXFBwk3DOdkjOlTmX4FRqnm+PuslXi5XntiDdFhA9F6WaIJT+vn3p1r6KOS/i
lkPtENpc29E7vkBUMcRbcnblXkWGF8EAaw4uf3cn4rD0nkytusVBVmMKT9oMCC6s62UMeWxD7zxG
FBUNHgPloSOsSmgEjweICKltMPCsER0uLJZXEWqRgCc27jvA0D0NnzyI89nqsCGwBRd505ij/bJ0
9+c79juI8F9IlO7Njdq5lrOqKWXiL4ixppQp18u5Z2rFCTx6xalk+4yN1bs4u/WGXTH4MMlY3eNY
uzgcRACdGRCmCGcU2UBz7JXjs282F2O1yujpwlU34HPxmvaMNrkhVqsuJ/yjeCAS2qgdYWZUp5mX
P1q7LES4R34DCvPuVw/lPCoB5DL6p1km/nzOVBiy5zrj5Ox1KoLQ6/AGcIo9FFh03eyyi+nzLRSA
sBeIwqz3QbIpjL35upeXvtC04kUCm8ghKXV5SeEJG2VOy97BIC68jIAn5mg82ZyqNKOT1IYKv1Oc
KwnyFOIhRdmyVZ/tH0G2Or24MNWsR67G1xwLqr7YYehMHkeRCd5MSDfP4dQ1l4nYXUYKeTVf7uWP
KUVvk2tiuZQPGlgRaHxI+nduiy+lFGXmwN157TFt2QuW5QrROZvell8z+3zUueJ2/8JsxvRa5LXn
0gsi0vABqqLShWFhpF72mzGxO0OR6RFZXLWcRCwkGog7uwJi5X82vVmSYNijt9x7oaTBfpByBA6v
/jPrvKmMQjisjvKTSvZj/8RWTJehp/zSR+GL607OoDiLOspuaXTVKatkMkMAXIn9xSCYQVbr++lM
oDkf0IE7riPv97pLytuQBjinLfdrDaiPZ2pGrMIuydn2WnTZ/yIKAAkIcsLUOnoW5slQZ17UEQr4
u2CScSsQbUCfDfPmHhJ/X2n7+iS+GVAtmKTbwYHN0tmJQ6ZPDvH/9Gxeh01EeIG4s9s9lbd0lYrF
bJBcfqDkwPH7N6TzBUweLCZyeP/Rdi8qIxZe4X8kJtqGgV1ZqgRNHo1UL+9Unpe50wC1UHTtf0UZ
WajFM59KwnG4lZoP1mU0SZSwk6yTbv6Gl5q3/4E9XoEO+xlxNQAapDE8Ao6WFG2jnZM0YsAB3mtF
/LKiO/4oefkOK2xl2IXFjvnSVR4VHnyXXizpuJhppF+oKYAYn93SIf17gWfX9Trjrr+cEmtalLUv
QhjC7VJpZawFrXowl/MzUXDsNI3oOfo9kx5tt/cnV4xpBKLl70LM+GlZHJFbXoz3cVQbLpCrDqzc
wyra7KkYfZ41gmt4Y4lv0GZeLVKA5v8Lf2n/rLbJblykPvLpxfQ0P0AtJMkepbzgoMxoQVyKejc1
cgzCFkp7WDSwqjjakT+yasllrnznFvrG1phQqWj2dGV+KOPQbf3yuq9O2BziRqNY2MwmBd2yKn4p
ke/cwkMnysm/T+3af134fSokwGL6X/rSVbABXweNyja+PM4ARnYcX5WtGaRAegMUGJFRTmLINrqN
7rZHh/rGJeVt2/4n0zuAft42hkNrmYrnVNGkQVv/TRB4cfLXvAWQAf2DiHenqFlKX43+TSarq4j2
JZCFxq2KK8mZiwkoF33h0wB5OOXrmgwNdF12w1vO9kVIJwDXB8Gj6aLVB8biaqcR/Kp3dAurXVte
j4kCNp1PjVUyfQ1IG3Ba436VRQvabhaBYoin5qU/7UPlfGL+/ohn4Bs7wP7CPcr7vfhu2FWVXoSA
m4xsERizr9WEv97jsTBpq7vc61NfnIE8RsiBm1rp0pblfaGQ8npUhK1dgeHYmuCVGuFDP4pHQlcX
kXOkx7kd0ME/F6jPj+b5HEsC5Q0hhaKkQa/jN1QV1dwUQGyC7jTMJejPP0zDtXPNWW5yq13EmCYK
GzJvXF6ymPnnz3yQPRtf8ZNc4Y+mA0PthhkXhg/lruh+5KItBcam6vlzHJhtRrRCX2eVr/5YFj/4
6XnkED5UWiONyhCfDFhlJ9Zrewtsaf6pA426zfECZRkRf5JqbSZVsABbdqkMXf4gges4+/IC51IK
Y20UakWrpso27JHvZPSCUXK7oag7OdbrxC1pkSu5xVsirVz/pqiAuiwmGGWGqQk7Mrgp1TEiBzmC
9fqx+DX/O/XO0qH0P5aCXs4LmQmfxvZkNfbko5USJeknKpoAWEYT12VV6WemCPmAPjuZW8khVWe/
ujRg0JDB7Q2TLSfFxZKi2U07w/3XqPWsbIYrFeXwrVKujofnpOQv85PkWHDgcR/0o+Jqscc9/5xl
Uuyu6RzrsFN2f3EcDK04s90rFdZVSGmitEdCdhB5u6o/jfou07qPR1Xg3WDJKOE3fWLiREyAamlU
LlVRFdgt2taij7XfHmneSZAQ95xpc81on2GgMZuEmKB9LDMkprce34ofigFlZGv9hLG4CPRhphpe
6Ua29GWQJwA0qb9OKq8o6PPPBGrTirIvtzc4B73CAxkDg9enxXjINVsK0ccO+JF28dpDJhqeEUKR
Tihh2EOMuiCPdZozvuCQKorGZRHxDjCuRqp8Bt0vZX5KuLEQoxmuBMQQIFjlYoY/Y+wXb6MMiJ1L
d5jKiCCZ+YkZ0GAVlBjbaIRjX+WXzdhWw53fKv7P1t0p7vlZOVUTNVPY+7nEnS+yn8yuUOdK/wvl
7jdbsznef9V7AdJqaQ3Xg8CmuFo9g1hdSQhdbtLU4/m94qSZ6lH/xoH/d+P9RBhH5VZB56/R63VI
lOJbMw3CcK+/fk8kfMz4ibtla74LOkeXF/BaYv8fpT8lV86PdGmFesThA+WXSO81aYZpSP7Y7XgT
GQSdeMaNmJTqLS7B85yC63TbgQV4E7GunQ4El2JI8afRiRqaOYE4GH4nvMb8P0SH/IqJenZ77rFl
Dt4PDnZRdaWehNritbVAHQDwHffxtyHlvNPr80asxdNIFBN//h/pmOmMhGzP6fFTsTHbPsbYT8ZV
Py56h7zOrT1gf+ZyUiYep239B6xDwFddm0Pmobf0+6Lw+nO/aJqWNSF4EZCJRmKhWDZbRFpzdh6x
XIffgj31DxUiI3+anw0KSdYono5cqFVqhsZvyr0k7zMdMjqUOOEbwdugZpD+Nq7oRZeAUuxQH0w8
nhpz6QYbNruhKMFXKMHa7CcL2Zhtf/IkHeF0gqMuLxfqi0E8Z8F2AHQ2w3iBVWJedI4bol572j+l
loQG/cf0bJ0Tn72g5fDoN0Waz69BRSFPnIZ1f2q0OCPZ3lfgWTOWaCYTXaX/3+oi+Nw60dx2gNR1
6BKsbUHo3Zu9KNSCUFccTS07+txx9FGYF1oqlffN4vp4V7OopHquD2brNUMB9O5XISIIHxRJNRuj
cPOtVejwP9tzSptGdi1//iFmnNvvmCzKxdr5eVzBG0bnpMxCpq6ftIbTK5m63FyHVL4S505Oje7O
RT6B6yE+eldX9jphFuevlq1r8WL6SuCrdL01+SougpSx7CIah8Isr27bTp41yqPgvfZvGZX6G2rn
moWVidp3Tvn9N87ltVkeCJua3Vtg8YhL8IUHLsPxarlJSccm0D5zJE9L5AqcamSKls7ZWx61+7kv
uvwViMOKbaTAEiTg1eY7zS6MZXxTQMrA7i1yn2L7Yv5dPYOMjzAIrIxKT29NNB9l3xsmziDtj4mF
DzIgvLL7eF57TajqaXm9jH0WoSBrarue3UFILS48u7t2I3/kdT/A8mhd6L7lxzJzmsXtIaq/D/56
DYFlpYzsMNILhkmhk+kaeDt4CLMTD/d7xOpx3ArJXvPxE6fjnkT+8auOGzYxLcKN+dz8Ss0J4EUC
LeswunJrx8j/pE0tndUXqEs1CJqtomfIRExR25nYNXX6bVTumY9FlP7K0YFsV/Ppe5OoTwmcVDEL
JxMt/QxrL6pzPKvbtPDMsmZmh6n3F786UmB5KJIfTU8MmUfrhszQtpehGYhfqL7/ah+Tw0n15bxS
O0DxETOztTK+mVgNQQ9ocouLtoxVkjo5nE6TkyMP0f1dJyZgT0ajW+gMypukL0xksAjwOqDoDC9Y
p+mv3gzIHKLuzV0naLis7z2xwbSW4YaP9h5m33bB7r1dHqOSqXBl2RB3UTFo6ulwtQ1jNqPCui5N
nG9a7gBZYlyofhGPWdbo5rinAXDxu2YJImuswQzQVAjABkr8n+02Fk1QAXBgqf+aAwqqhgolMJg7
eEY9ZgcO6khM3KNGjj9DRgjp3e2QRz+areOkWx3wsrxE8oHjVB29PC8grQ7RRbSqtV/jtap5oWwP
YdTTuqC/hiMW5MeP8FUQ9JrvFg2BvMM3EGltHFyPwxOISPX65vceb8Bdj+IngiIkA67G9/5cRKVS
at3LG5pmedJ19elAzu4lLCG/wQYoAN6/vhHCAqP456hvPEai+R3OsBrwqXr1qhFlXXtsM4nrHZy/
5T6uAH0VSNK82ipVtfS5ssMlP+vigE4DXkfiYgoGVM/tMV14QIVKfljzMz0RMXd2rUkONp4MQ5QH
wU3zufFMOAHxKlDKnFvD5BoWjhG0FX6fyr9WU0y3Ewxoa7sUOsmXAHnUft0tK89oQid6BrJ5eUIS
cf2beLEx2dQJ9Gq+QulEAc8F2fFDzS35nOY1dqI6B9nQsQvDfOZB5lZrHttaXc9I/P/ZA/OoXD9n
4X/FSHVcHJHQKgBXk1QVVoOJ4EGQD2kjUtyu72YmPwdggzUWQjV/4v07FDceSMxT9SlRbtyPMXiN
KDG8Ufdab+vvFmhqS9Q/pJX2qIOIpOuJlaj/zt4YGHzcejVQPfHY4NT8aBYTiMB7eqSjyhPaV6yV
9231FnwqPbky6D7k/27xY5hPIre6Rdr7VYe5lRcvD5GEuXjJZjV6EB0HSGupjCeXn3ldRhMWoI0b
aO+ve330tD5XwiOOtaV1sgJQ2CXV6hcN431VblZK1uQMMfsZ3AmLgV8/bZgDeanUZPBFsV9wSm+Q
oV1+aDPsPcWN1aQusUFqW9QqTJQlyKB28BtyD+G+i/V54F28zg8sRtG96rk7491xUNMJNOuIiHVM
xiBeVCXX703c90dbqqqdr4XXVUQhk9zmL6eQdP/SghQWpnueSa1vE39ZHZ0dLB+iaCokUoCKLzWn
uoFjKZ2eBowbzd/XSzbFU6ZzNyBrasF+lUhL4LPG7jtCe8/LfUOIhfKd5CKCgJSDuEZ86TByQHgw
7AILfRSf8q3am4ptoDH/kksw/Nx1/B6TZwlDdsKmfNNk+YPnYxE4hum25matrtrNu5RFRKg/lpwJ
Aa9UNYBKh23Mt/vY21Q0wOO4cOrhZnkpKX7OQwutbhSKOcEVFlevE5ZcNVsFRPCgJ+RlP0MoUod+
rYS2vE0wE4UnqOAt1pa3znC8SN8DwFvAkGGBfs/fVLfiyEFeHL8T3UuPM7bslxCXoWenSxoDm+3q
TmD8L6KD22hA1YpX4+Jrtz0hWXOfZJfdX6wyqJwTq6kc1NQcTQBCAP/yHjTw5npqWaHbXAlJ7Zpk
wt8Nc9lZm1nFSChNj3iXtldXUI0pdEetg1leZANLac6OvLQBAYuFjSexJSqhOsnN/O4yMpSQt+i0
q+ryxIAPj4udLGEX+EYVLBvw/6aV/xdd+uhaqlro8nqkbH14Xwuvl0hTC3WDDZIF/FTm/Br3/6Jc
/cPmEhqXpajGZdFhVRMAZqFjR3BMjifKEdn+fg7MeIqZYGhuSveKfzTd3aQ+3f+/qxUAXwc1zXkt
gTvVpznyu3skytxZj/P1FLQs9jFQg6Qjdjn8uPPpw81f49OG5qKrh7QyXoMkPRdllPgLJ13+JjY8
XL8LCcHd7o4YP5EzafzKIEe/SeA7+NPhm8zloHfl1UU83MpyBv7HxFkWdplMH5dZ8M/ObphdZ8Hh
BVbMCxeZecpFaNbz2ZkzGQPvatM/osAKE4uieTFy60M/nGlgdJEoZFLvuyDOlKhoRnxbmGJfvjN7
geFOHFFrFimTOzY2ywTbC6TDd1x1Sx1hR0UrK4eC1pxTeYcDzQ41tTSKucfbI2ii7hm61UD5gy7B
ddRYYtDCFKkYwZzIT6K8tvt8G+0PXCnNLQQPljh91ixgxevq/M5hsTp5voUhyYWS2veqMklOXtyo
WUvDjOAN+cFNTK2xkq1BOafS2Zntm0tXYd28klRpyWd6EtyiRAD8B7DCkGxGGpzreXgqPlHEP5Y0
LoVz0CGN7Jm9XCvkyMBTYARWLlF6SUcRK/97L8GZ70/6PpJs4WM8CLvGxzv8wpEhg0YHTVUy0j00
R17HaKuOBOovtumuBre+beD5WuvslFkmRqeqtGppq8y8k+kY8amldm2C5BIag7K7zUFdD1ZnevLS
RGpP8EmR6QyhreUfleJX15f1heYDjxMphcsb02zo+18cAZ510DHNC6kZSle/wbeQfEpKjB3Pd4iP
akARypeAaWWcb2RIXPIMIYV9TBJ71gT5+Gb84x+wAOKFV88Xt9qH7WfO7eg66r7CDcdBqpEUxyqy
5ZrpmdtPRIFDUAh9nelwMp30ERFy6RXRCA8LQuE0EIHl5Nb46KMZ5lyZpaAg95rSDBpuWYAhQC7+
X67y42pbxy4ttYooj8TuSzlyv+8GO4bTpx/+Ye7SNwgJOOSidn48t2qA8uhm2wQIo0tGQbBhDKuh
F/ciIT6AEhllciKzfWeFA6dgu8xYRY6dQcJcZJH/EPpNHCXmZlthdB0itVJEYXxgHYpq1mvH3s/s
RaypOWJy8xc+72dVbhdIMWFrgada3hxNYzSE/+FoQGL9WjGm3LYICa8szzCmxRHiR37CCNMsfcJX
ix5wFs9d7Ds9UojSw5xRf/wLBHkaHJQJeQEPf/0VK+KeaoaWkiSgLmK0sF882k5E8n4ozhT2s2he
ABOlIEo+kiAfKOt4UbGi2KQhslmLEdqtZ2XYsxN1lVKSzssht0/PKQUHXZdttev09gQyFwfUc2bG
7b2reLAL0GFNjFCm9W7S77VsLdDC7AwSgBXkkhSY1nu7UPe8IwMls7IUgAOVYnxEXR4H/ccKpeoF
21RRhkt/iX0DAE6xjFFms4Gb5kDyuLGPzhq4aFhPK4ir4SZAO1jFOYBrl1evUX4zUaM572nRarBy
n11roFU7muBg3apvK/AADnh5uTVsS0gCW2QXQHQPIsyI0maTNNmNv8Q3EssrIMfF3Mb5ek3tgUVw
bOSGqyon3uSOm5Mxa8zu0NZtRgH5hTRrqWrhpqNnmSBDSG88lDoglERce+Jzaxdj+K5wABV0+I01
/qol+QwwkDESDv6UTDggsXi5YjHkReVVFWUG5dOu/zy7t/Y6h/BGdkLk1oYDtDsJd0FpsZ7fQoQ3
e+tcrN+QIlQ4RFNaDEW4bBQ/v5+v50bgBF3A1JJFUl7fHw1x9k27VcV7GWzFD8fQkO+5uh9Nb7p1
4U9lFU4sLbbPfAFehrxpWKclprUmrTK0EIC6Pi4i2J58Woqo056hyTo5+5kqwQ+AcZAvgBQXT9ld
G6AIB+Y+gb5UIRpPkFk1iDjlHLp2VzjqdaXhaWKAx6rAHJXh07PNGRJCLsosxdhvBZmu5caoLedB
pvl5UXQKtbQm2muCzc1mkaKlvraPQwNgDReSXYAcLoWWljtKLpVyQiiqBEufsecO/wmkunPn/KCd
twORJWdY3m7gwM0mRfZtBZFiSnSr8Pm02gYIdG0Q+PFZr7ZTafDgvBovTsPTS6FD9otHNfMQXgaB
d83oaDHNWhDDP6nEUrmdcMV+/lV/geiiAZoekP1P4lYCk0PJm0wzMTAX4fF5Dce7KNzxeCe/Sub4
+OjowHsJUAhvQyv/iJgwlamrIAPmC+hcgtqtdCxGu+k1GwQViHKyI9zY4dOcw3ovotSOBoklRx7R
i2drPkvCTKbyQnJ+w/8Ix7U6YFcRNLaXDNnpflMbsslaoSv4cgRSvzWRzq8Twt5byqxmXytPU332
A2dFIJcD6318Dd32P40+qU5azo+MRK/AAPeygB2LYKDTehpG8GBhBaLAxSRoFkMF9VEyzPsXWK3q
IQ31V0qfsF1e/UNA2Gx6QCAuBT/cI4a+GZpa6jS4glPnrYFqRqgM86hJwN7nnt6EuMs48wLTcwto
NYWx/4CVBQtY5w1YCscoAwyX+WD3G3pbxD7EjsHgZKce7M6n/plDKSvIRyzKl3QGLOj5jMPmAuDT
vqEj78FXGna71RJw+qRvezEZMK2wTruN0dbmp91lbtEzHjWgRhU5IIJluij79w1CeX6RAUbmrq4H
G4aSKplkYDdFvatHjPBZ3A9GfhqoN1GebBun56zJXA5v2r6EHbGBSi4jwx/35CfzOhVi2F9N06F5
DLeoz0R2tBHORdfXiAiPc2pxdGDbo0k3W583B1D+/jDGc1tyBbUtvA2fPR0N8P5Bnc2HHjKi1FuU
BW/pWZqz7Lg6hrvDOKgK3B+/aNebzl0ZEjOWoBkA6LyeMTkXsuSZ+h9h9ADnq2teHtoP1f4y30FO
rrUbXXIOLGB4V4Io2kj3rFzmw5wgCAB9nbbl23Wqdo0SlAoHcLKmQTqg5XDtWh18G9IeqqXYYC0e
DUBKeIr7V4uLvicqHvYVh8yuu8tARLXzNGpH3D32mLSKZ8JON/xN5mUxPODmI2FT4IYPCMdIXXVY
FLyifQ+B+hQ3ilhksPnPYpYeGOQYy+dagDfeqkhgvMD7Lr9kjyv0wBT2E+GbG+h3Wn9LHcufU5bX
qiN/w+RQcScoDQ1eodQyQ19WU2L9nfppUgFfSgPeNMl7zIt4AOocAZoRyRmNOoXO52COGc4FEeon
dZlk6c58urGZikEtpDZjpPSV4O5AuiePD5wFGoF5HTX6IS07FJP6l1LH4alf02O71425vkTbcYWu
noXxz5NLxFtDg3m+Yq2VGI7xjOTooK0/MNQeDveawRaUskMc38/mbBAah7FG618IV0YhbxNY/rLy
F4F37fgyQok5VvR2DUZ1mt6cp6vxXUSosFFXxhJmJAu5nBk+yOAtnaawgcrV3gNoUKXrqYm5MwL6
tn8xrOfQCPaMSpJ7viLow3K/ALkt2dKSu4dI6fCk+atS7aaA8ezSJzRaM7CFupbF/RFx7JFI4E41
E2CQzSHFm4noGmhnLGHa00+9GDaeLsRsaLu4WrEnaumJ3vMLWKIsEpBnRiJCgj5DtvlwvU/mYen8
xqq7XIbxSywb9/yfNTb8bNdPm0dhLT/IfD95yiEL/6uHq+CLdq7+CAk1SpfK6O1GcqWljaGkd5G1
RwibIyXCy/QiwNbUjGtiskdqIEOtENH4H70Ms66TzkCPbGU+Lyi9Y+mmg3a83Ztl4atFKYqzLDzt
RGR325Bh4avP+I0qIWNj6QEOndYDY+5oVk9Raax8D1UilZkNXzNC5lRU3bz9s7KvlvTrN9S6v6fE
MYNF9r20YCQdhs2ebJbZ/wdS+LQwOABCyJE0FxA6uMYDsHUPXjjze8UmMQYUYw7Q8YwPbui4TODN
nZdF/pmqd8MQ6o0ngPvEyu75Lq81EfaR15HfkL4a1ptiLAsZQzDlBwjP9gbXJEAI3mhnoXIh5ViF
YmqlXwU8yWR8TAfHRhn0EVi3ajP9RB8I3zY+quGZUR07tgJAr+kPiUx/wERWn66cjU5X683gXETS
EPTZ0oTlq2RJZeoNQbJJhmeC61QcJMkhgBkjG4hzgxdFPs61d5q/5mLlwOv02xM9n7RVORW7gnxV
4DDMfTYAMYCEyZBqB2cC5w3OeFZrLEZIRX7glWk29BHx+zNMz5O2/hHR5438qSHkqjs7xWNsRfKb
iNOeTXoqL+DMcKqp7UzWPPHB/fEPT6KYh1z06xf7w7ixgGKpjeqIAQdrnTsQH9ljCY4bHJZfy52g
5/wq7543mM6zRVEySQvBQSFMvJe+BrQbRGt8gu8DcIsJ7QvZ7z/eG9A4iS741DSpuGg+uv/6ewnZ
EGfvwLB5NCo3KoQorulgxgyA7SOesrAKbhwIUCQRuCqbStG9dtG0V8qgBC904JFkwORY7KIir+E8
cezVJS1xyiZEl39gkKkYj3oe/FFZOtvYwIhlkBkwVM5a3YarT7NDl0v03uVjAwQBkRV+8EUS5n7Q
lIhAfPqxqZZVL8sXcslh8iX8TZNZFrI3WnbBpb8HbtGnVuruVY6qxVJd4uJ6qUKeNdI5mLdbFLyr
IQlK22I5JyzzQh6oM+H6z+zmIzciAOD4XA+x/likGPxCVIPH6e6T0BLkfnyGU4Fcu1EntE+af0hC
ho7Av4/nXFKMbiZbHBWkXwdZxUvfEaeUNAo+M2PhRUrkyrXYjoM/ozdAHZOWduWlP7rWHEMhVbZU
N7SV52K2SsfDkpqY9LmoYHe2ofOvjuMwdnNgoOTxuHlJye8B7EMYk4h8yS8Q7nnjvR8YnER/WP5e
4IG8wOzphBDEwpQjihnn+3XUCNCzDE4sxDu7PvFeJsuRGrKybU805tmeZttaQDhHfrDMRXKaJfru
NGXnetwgt5cah9rZ5/GC44HglwPW3E7QtAk01Uf2nWL+xY1F5nf7mTgqE+bqo87lnGqS40BGjaV+
U4BtE7fPQmQgBhACRiNH1M3W1WUNKFhtptTTc3VDZ+tPUiZam7nVMOnLfEi+bdJVfNw9P8nXbeU/
2WxlsTriMXvxw6faWN901vfrNmn23AXbI9rM5XHKBfyUsGfQoCJ/I+5w8LSTGTsVa4ekeNieFdE8
VMj1qc+fMdJ0qZOdSho6snrN5EYhJ+xxMiWrSYhO70B5t/51U6dE3XwrV/Yy1pfHeDc21r37OIxY
kKOs/VX5W7tHwyaHyC/Ub7RBlDhjtfRg4SOZjDGJAhJRe2DpyxNS2DH6YymYim2LnNkq0JKuD4XO
MpXoMQ7l+/JLju9glJtHA5qyhDWdd//4zABBZvBKGcbXfbgte5di3JOoPsLcaQdpf+riBwwettER
lveJO3xw91MzREaCM75ZzRYLxShg77rLujbn7bnOFJNSvyCR6Dz4tuS9egzk7sqs1x4M+Ptfu8ky
UK4jXtxCTvBFWqkOUKqF7jw/tjqlmAQK3nzC0KZA3yM1DoXJtr4UtXpamKHgAD+1Gl8smkQRyfP/
duBvVgMas6O5scc58uE2t0bjXhPmKoh/2Cr40zRH0p5Lje4wokRkYOOyZ1u8DLO9fAs5W0T7vtJ4
zVjIzwuVhKMEzXaEcEEYcLeNmqMkkFgWGXd+s6hAokL3GEGR/gcGjsyIMU/2/HceCySH3A+QMlUv
lcCkoETxNs4whI6ejWSYrddfwRK+bzJMPjUWlwFnwh3EmQb78rRmcRPQrj5KpMSpNUWk522IPr3G
snK6kXtKfBKZumjD8Zelu71SXL77UTxOOsNGFgQbZ4iwJn+JCxkN1sxrJrswJ3N8Guuohnn/bFr1
9pvXopK4EuWHkZVz1+nGqofzf6PRsfA/2cvdaMfYPF/uNJmMKloFtlzm2TKex0RhkW/luikUCtlG
E++3g3bPsQJG9+DbJZiRP93RZdvaAyGwoqzliJcwaNueK0PgN6VENA9K8QY9UkysSSd+8QvEvkp7
p+omSWJqu2UyvlbYOHJU99yG2pGR2wi6Z7RiBTFFMVpZmXakU+xyzkRvUkbIzawJYl+NEusbFhSs
az60AIMoDFBjE6zQoSzgJ+YVYTuvrkmtcMartcN40L3brXa0yt55+tgMc/7+lmOS+2kspkQ3xqCN
7JePCFoqefvZ1TuV3rz5jpvNgSEv1hXaV10/nKfSdT40CewGs3C+tz1rQ5wpIuZxM2/ZcsWDmAL6
sy89nut/28V3XL9cGABiPRFllt5L0HS3XenhuovI/+y5oE67/q2/2DsFf1h9DRY7oPfUUbJvGUHc
+cyDymu2wTaZxZoROpIndUsKWmRE8QcpLTpOqo1lO2x1BWV76K5S78ofi+5XipZkC19w7R566bGP
PmboyBYha88wG+2l+HG4zFGx3kahKzvHfKrEgxZyfep9YMRxy+RQ8KVq44ooaj3nkrzZTslXC8S5
KcIN+IXRdkOm5x9E1J6R642c6BkT5kMQi931lEyFFKjN01i49JrnSSdLOcmyTMCirHBy+bcaCSgd
Kpn+q/AaM8CXIHGr8E35X7P9IwimdcCwbGCAncA0SS/SXuyfcMiTsOOU5asIZRtDx+RftCQmdoMK
C2of1eYdC2YJ71ZI0Of5LisEgaQGQXknTUH0lY63YTBoRMEpYwpqPpS5VE6pePpo8TPB7APM6ilX
zKkweZyh+TXkswUs45QgeMSnLpbglNQUXGKLWhW+8lCZ9GRKp1Qj4pKH1hM2Q/8zRmViFMJU/dRm
yNg+WytUc+a0QDaSPNeT7bM6WpR5SPwUPtsji98Z0ndpqUVHjhaRGZ1LVe+kEPwqfN4loLDgHAoT
A1WMNSc13jhrUOOHSPG7xSanoZLedqHvfC7upEwhNAxZrKpL8vVh70mX4AGzpVXxWHqm5MrwIZH2
s4vMdgVytIQ1FXumOWw5a7QcvyIci8hL+6IYwncMRpaRnnHVH4skUzABflsy/rI8dAcs4qC+XxiM
NWUE2HTGl6WNqMyrdrB3/DSDgNaieJFOgpGBeFbdG53r8l/vt67yxPyWPiroieZgbzN9lW3AvGyf
OYZklcBwkB7+nx0Sl5QrnDbT2B8duZtNz7ppVbQQt1eaop5ljl7PZJAv7B1/4trL4C6hZQViGEd+
ZZlrWOSXJ5EGMVY6LgAWSH8qehFo9uz71IEkB0qDNQf/UcWvU6zxJsSUOp5V89Ccr5bj0pVBDRUN
Uk2gkmtea8D7TIKsgjet6fpugR8i9U6/SfObmItMhdL92Ulo1UPzKe25g/Pqz9rfGTAy/JPVl3hv
fX/1kzk8PnhK+bOnWFDji41i2FzmMaO3Xrvoejk8a7iGbD+3I0mq/7eqyrI23hkdwTHZXWWzDdXS
T7V0f2vKac865sdBf5lTxcywYtzarvLIPMsqmf/25gnfBMhlJ+qarxNbc3cA/WnhxVIOMWTDdVTG
WjycxW1Ce/0dO1IYagLu9kLw9gX3sDS/BkIHOzep84G5b6Ykvgj70+5veaOfPh1WP/mlPRQ3bogE
Wm1mNfTIq4wdepESz69i+adrwjCSPnNcu9yJT3TNNpaLOCa7DJKxXOX7/LYsrsOIPCVnNMW63CFa
3fosFhRsik70kElfgezUqPSvCs9r/ZmLFLSgt+r9MWFrXgomTq+UwXsAwSmnmIf2VlWS6jmONly1
mdBFZ1hM4dbJbxajI9jeEGHyNcM7OERKVO1I577yB9daGNu8q6h3NFh5TxqqDaS7Vm7cJy1+6bNx
xvXhI9goca0V3BmNDP0fWxxukiPAzx//T0m63w80u1GBJoKzL+466kKwbmeQnrecaSbXqSaC7+A+
9MrTCsvt4l37PMDAMdK5FkSR4aa06FcCs2ghu3EyU8Ax3dl2qLQhqnQmzKDiqxNb++xZipmCej2L
pw5+jcGZ/gb9vAnI8giKKwZ8sa2nw2sSRIDiq/cNznVZy8AzC6FwalJRhRHhbM5rWs3EqBs9li3R
u536M9MNMH+9l8z4s24r1SdjAjwD9QG5fmyFaNflMD6Kk00SKTdbi7wz/NuCmmmSWrRv4KX+P3e7
guZE5ZSWAeBeA63dxp8BBx61UQxjE3EtsjTxDlhG12b3AjTq8NuohC6GJjNOzG8YcnWDNYh11TGF
FeQftEjaoszElLbVxbPinxijJnWxC/BL5ZszoS/Bunu9imOEm3HuF3yTGysT/cZAwgCdFkuaGh29
YB8anEnRx9Wmah50j/x2fu3WqXDPdDCwtr8RZ0UeQnV3nFPofk1dtA/C3y2X9jHuMt0o8dZpFQks
eBywXwUHC5+E0IsT8/+sGDPBSS0o5CnsH1bsXxKTwueytH3GuOHdkBGrTV8E06/h9c8gbBlvRct3
Cm4zMMYnjGc4IAhiW7AKhBEfl8Levz8dbWJC0k3+8q9/RDIJDgsxCR4yLruMyENK8r9vLU9WcuGP
s57XGjBUUYJTq14YjmteDAuYiJ6UbmMQdzUDO9AqlLMLM6jkuAoY0t0M/IuLqu/uDHyf/gjUxr0Z
yEzvLHW7pnZPcaK8s2WgMeZ8SHNj8HGWWS5qJWebw2IDkUBBbJjDTBclWQu3qTOYhQa9oGDvI9wv
9vTI04qI7QTc+pyqdV4YHUZ7FjQAXXrbBiaJuFysraYa8Z1We6EhT/00Lj8gUcN73bB+6HQlF6gZ
ecJkAHjh6/jWH6ss2ZUDbA2e7NVS7Y73j0hHDqzo08rI968byNVCzxU3K69IKDEykGyNzPkG1Xch
ibFKWW8GUAoTbxPD9h5RPCGnHVEEQszDpTloVexVo3igNfKNaFZV7KzGldcl9eV6jxk76hjd5Ogr
H3cY1rGWX4bpRv5l78bcsVqz62khAm2rtIeH3Kd+HnviZYQ3BTIrtAX5q4B8CJQEPb+24C6xyqi6
z2G88qUMLx8UD16eUUM3CbwGEEAgD3EgaqN2gBabFOz8Z6S6rR/QOnv/T6UoxmcZ3QX+4zz+9fH8
NbBwH87Le3ZqYY2iFptvoJSPKGkp0BWR7cvnHdRtDAaZVN5RB/Mzh6599pd8PQcspJRk023KiTpF
PMO/jHOf8BDY2oFe9625KrP4xei5PgW9hHLjM+bQKb0D61nFWV2vm4EIhxt8WNE3e+bMj98ccTZV
pP+y8DqmkuRNxh6Gw2liqebhFFtVlxCsKqndx4Le1YkkM30llo+gqr2PBdP2ET/6vqeVhThecoqI
SK1vzrIqMZRJo4dck+mQ8iUoQ3FGFL+CP75JQ+DX3huK7jFoMi8MRUyQWz/wyhhN+hD8EserTOUZ
lFDZOUIiYO497FPddsdvacXkdXZycUuMsk7UZXyTmXq9G94sq32p6wxyfAKbqy4+BT+456T8T4Ua
9FNno2N7+gH2D+JCnAjZhwSRSd18myLGFciNUarRr96TlFkekOHr/TrfoUIlaQmrxXUwuVwK9HHw
0wrTaClYGIReVEiEZatwY2lMScWgRr6ALo/M4oepgrc0FiY36KXTfSsPBbLNWQu+RDtzNczxO6+T
+ucGxQbj5zXEqdWeQI6LhYi7mRSLLB1s7KTaPiFfz5lIg0dtMB4NQzKc2a/oD/mf/eWUo61lI1xI
usWlcrB4Hzm90tAqo/Ua4Bg2up93FO4lY1L8KH783VMocj3u4FdhxYePdiTNOrkGZHGKFW8raLmr
51vl/1QPS7RIM/yHdbLVRWTOjCoS21z88kfAtlsw2oWQZzNZicu9zLLUPAMMOx/z/I5Cx1q5AWUb
Qo/tNz36jYA9EapYBeeQn1k/3Hl42DEZdHOleA7ul6GanNtFLqjA3j8HzC8gqzVL/F94s6cZkJmn
WU2hAL2VwodkqfstXaxEqF+8i8DYILnSuSvuelI337L8pZoW00rvU5T8rD2ik8xsV2npJVYkJAUi
9UzSWFnHMSdJnu6qaMh0HJgaKfqgKklW7L/LzbnAFEqt7qsF6Nyxq2R/mwi1rJpycGO80L3xbGvI
iQ6KzJWI3unqpOrZWhrJxml45PrYxCFWZeu3h9qAZuFmxQ7cn5BNMlKj/InJaxMBJAXZvk/7ByfO
dBPnLO+mPbeFVrWPyM4hTzlEoybRiPJ0ZZTjp1pFF2aRUCoyPvcVZ8TeBWpio+MguAzEXITGtF0P
ISrpV2Zm541wRwoBqZOtCD7PFIOSG/mWLC4O/m5bcYa0QxOsAI1D4zBaa/oEKAGbpijLeQEZHinT
XKhRPC+6xpQ9Jf6RKDcMHY1vGAtZ8KPmrTNclcY5Cnt5UX1ZfX//xLNgoK2DCx3eRgZjJQa0efev
yj/X5whLd1GX8jGDqLoP0ohCcWBFu7+3nEi2soAjvlPQlsEkiI+hM/uTlZuglloARzKmXFgZX8V6
bC1//iklddnr0sjlgk35TLolt3/kDEe1NBNKKIKr4opFIzn6wR/z9riWcaSoGUfVmGft881KFYyZ
yhuuKjGUK5ajilrXaWiTAOqYsqDVpMUMzCST7ShyHH2OrLha0VXkRsduEg2fmm/2DunfaUlW+qaK
YncOK5W9v8HneaA2PjS/p2daGCSaLSlmU8gekRk0Ncy/l8mUeVRrcZ/ydc8FE2ncJofoJoop4S9N
dWiwnp5Zp1553ExrDyQqOE/59YS/ohND7lfebps5OmL3p8nv+8xUJMBuODO3qnhoh8LPY9bZN8mB
c4L0EY5+ov49FWqh5YmfLhBYQFaWE3MVkvXp0U48U/P8IBpldmGfPd/3rKGcJaLREi1GwTSa5eZD
s6pIRN8ANvOMGzZZgyLf3a2YUO6iL2ngpC2yzLVyeIRBrRB7bdz5B9KN9UFYqgoCa0x2cvbOMH+u
v8tO1dcL4mNh22yBDvcMiiG6APv0gEpD7jrQzKAu5sXrAiufCHQvsItUvHjIN7/XceXBuJLy8KSE
AvRatNQO3VeHIhPGN/sABm/Ygr6wjFDwg7qUhK4Gn5zzk+bzh2dZx4fOJrcobaMyEWN61uWZV5Uy
R1HcdpBDWq7NY856Eui4JrkAiWvjeN1aDTXPSX3V2HMgHiKEJCx/zBUF1p46lxvGTImnjdtqKC0J
9EwXfZZQ47SHAhz7m8dEQ5Len+5DWyOkwFQQZkXfYyWjWaSbz+GwVUtYdyUuMIUtob3q7MBrYyJT
vzoWwp02YKfYLr/GCwCPLkOtUbfbMj+k0K06D4C1pvd/1fDhy/lazdE42Ne/T1UhdF3hH4v7yy5M
NawQq+uAM/wQMTcspgnKWWh5999TDvIvb/1ndzCAXC7yZbM+N3SNtCc5RGk4Cv2TXG5q59qvfCdK
WD5SLZCle4t/nEbmDUe4hbxKmNIgvqqDEG9XW1FdjyY0QrdsGYnW773ArUQ8fAbTkM9Qc0RIOcXq
mdgVH9oBqGpPYBYXggsLoEEinDinC6zihdbaGUcHGP3l/i+QRdU2pKvrlqahxfEeN3n7a7kqs/Hu
+mgOT4JGuFOqsPP/zyGB9/0aPHXr00ZEuwNaj+nSnSe8510m/GLyi9K1Uaizvb67WClDHOMCJfXI
q5oW2XwfT+U1eTIx3b1Si2bEag3EDzdVFADqv7TtTjtG6IjiQA4Kfncn7kUY2aipXKLuXgDzcgN5
4YoRkCE9w1qO2fWOMGIySzs7g6X8KBKc+2mh8YSm6MbAbvP6+FDb4LkRSC6ahQ6ncXnXkKcLRK4B
xp4dEed/8z/wBXWeHdxlW043Vh7PuxfiJEYPH38E0sRrsfGPBG5nntuNGJoqcDouGSKJBuHjYlUC
jDAvoJmr+R4yf7LKf+IGZ9jfenylgr78zV2E5ne7GD8jJdmRCQy8YxfLeWGUdbwd02tMTcLJokxZ
j2bfusC0jzMBwnen5ahZ9AgQipaEhASlkR8kPHbQ6eCd8E6tBzzPTJTxPilFBn9Ge8eLWqisdUph
XlZ24qM8yvRoz7h8SrvmjsZMnu0XrXG4WA7k96OCCYuHr79e/Wchl/+pa4YaGfL+J7qhcaQtFUly
GHRFcaGL1Da3qgvfIJf36AIFjby3fR4pb9Lxm1j01DswFPYwpvNKAmPlZ8Z92h4jN0gU6njOKXQx
Gk6TdyNdYGbbd7FXU3ZpXI+gPlZQqO3cu1eM2+1eWXUc86/V+cW5tH0+vKgThaMo+pJNJWNgpHcb
io5ZUwMKQlcuPPtIWYohfDPke1MuNuNMBQ9KI88LWjN0VhNV7+RkUHNQTluuX5Yolsu1gVIf66ta
KvOCLyrqGU58xlQX6T/X0h7ARPls5H1dXRRzy7unBv7iD++Evr3ZJ1/nfr+yoAk8mANsGKfydS7D
fkgx0epFze22AFCmo8Eu5uIhCfBOSke+Ya2oZNY9pdurEL+O6OKnYywln+tofbrU06IWCmLcq3cn
bD/uhQ0+htkW7HRnSQa4iSivNm23tWm8JGBE4oq7gmnsjsy+QbAl7E9hEpT8U8tmcwxyRmoPgHv/
hwzvAtnczVewYSrHQhM+trx6bBugYchudQtkEnGAsqyQppyEOC8HsgnjV3MY4JY82GF77Qq6Y9+G
tHV/Ue0ePONEva9CwqyThwZUr5McIHecLz+rX64z4SIuMZ7osKEr5tIV7J3U/hfR9G4INhQpthRh
MG481ZEIrALkBczX8X40IWyoufFa1lCeqFiOVl5rdvT6Lc2AfQwTs302CSDEBfpCCZcSIBMXVSGD
0ysreWKQvzjUysTIurI2HXZLCfHNvhXhFKnXbC7MJFkEac1Hp4VJgsufjgN3JxSKakHJ2/G2kgJq
uyYA+EIZ7Z/5i3URFgdAPmt4dAk9KsiY9fMf4GuUtRyUZOBcvcy6JQRY5di34sa8JEVzLRJ6WChv
0cuenY0LB1NJBuwbIGIwluCl4u99JNZIZNyNx7Z4foPQfXv5r0m069z11TzGXknusZJd49mobF3k
2bdhdNxdhaIcPjVEZENUCretiJhPlJeMR/r6ZkqKwTJXHE08kP9nDYLn36c5HFZEYnTU3J8c9WT4
qnpx7sdE/TMbpl9ZiQihfW9eZngc6myh09bdMM6FEkUW4kFHPY3BT0d5wvD7sQ50Eix3dIZ9ydTb
1glmY/K9eBhz+s7JkowcGXgDqRoJt2hZQZ0KK+FGdOWdgaH9re6PebJm6lzzTB/BWn7ZAO2aggvB
WDfMq5BaZUm7347aly3jdo4pYcalyeuaZH6L8EZNp6yYbhSI0QtqzKTadp2/ujIv1ol+DskCKOvj
33WwEJ4TprZpApnbHpw95xr8wYGkKwOYwnxEJlb4gkAH2+/fjw5zYQi1yGzE7t6o7v69tPNTMbMN
mfT+2pYdU01eV8rxn7aKV0QwtraY0/XXJyjP2msSwl7Y+sT5VJUYsL0BJETLIZfIv8jauSjHYIsJ
FGSCcMnGsRkUGtIhscbYBKimrpYHQ2NRIL/R6JdzfDu1x1+9aVlqWSgbcOVjkz7IJfpcStRu7Qub
E+tLcAwy6yFImZ/QXWLtkL93BNeUYMOlgsreEkKTDeF3VHLQYBRmAJHRnjNia10PCSCMQW05sU9f
2OpnRStnof5dXeldlEbm25AhcwfkOxJLP/LIdFOvUeHb2XUwCGujZ3Xh0Fc2nrGhMzCuG+QlyhLs
P9bqWOuqRmn8hk19XdJqZ8k2hb5b/Joe9WVySoSPwQBrKrLI6rVZPgcreLRzM8Nl1YQ/DqjdGMSW
BALAGeaYR/j1goCGf3y+bQtHVp7X7XjJoiVTC83iZll+buav2jACswgXXDTA/ktHhnpbdoMc2nTT
YprmYBkaNOySC1gqp+l9ijdolIHXeN1VhQnVip9TyYqoxuTyNvRw+IceHybmlFZgD560FLGYSevY
wRIbikCgiTHv4dzEpiIzQ31TrbquyR1SbrT9hH7G1v/fFNwV8rWiKKYP16sHoF1QUsf+eOV8Jh+0
UjDs3JMBf6o3VD/wlXhf8bZ2+TtUcI5oMM/8XBQhuXpnL1WFyXuOIYHx1MEhfMFNFFAzO4gR4LlZ
hV1xpCeV1YMbMkF9BEgDnGnsynEQa83idu7+kv5zRTLYk3GSFx1IS8KePb1KlIZFi8X+A3oxCA1+
u9lgYDBMmxIDFPDry0QdRCJaS/p/F3e5ZFtzdYqFLA1zT4JNynF50Bab+kI43UmXq2m5awHMTunl
20KvhQU2EWG1068ev3wx2lxBD+L9VvNhZ33o9uwUiNWfnnfsqFMR12CiZb0KTKn6XfDF36Zb4Z1H
y26wyKy1+qD+x9FszWeL1SqPcq9f2XWpu4RZxL19eYkGbtSAMgDyA5Tin0MVUHhImBnTpccLLWoG
7wJ0W6MC0uDaMxxYFjAaFW/KlWdqTh1sl71lv7npB6GhbBWx514lrYcV4a281UNPBZAUNlgPwn9s
ZYwwLXDlolB9OV9b/gb71UI4v5r/dChTRBUntvXSbPnHm81Iu17k4EvNuv9SGB+8wZ8w+uzgYpSm
8emQMdY5AjDoVJMOX/qENDGGgXvsF0cVPCE+a7yB57wmNLNW2XPca6oMGKxhaKguYHIbJfB94XEW
QdaiLQEDJc6q2lMQWR0hIs70+RhPWMEVELuNsM71e94IECx79FWgV5ZZLN0LrM/SzHJGNi6WHbEi
bG+4R0NOlBxOrreeKNkS8XdswBtwmKtynSlz4rw8XQh9dX8yp1sGCaqseVYdMHYasUQqe7Mb67c0
V0zZFjA65mjrb1M8w10/EAxJSsM+ydwTnxG+49nBW1vQ7BiNydzxeYSO4DKm0nlx/YZhcdBT4vt/
4WdIc+ng8gKai7dZiT40plp3QGNVribMsEvtA31gsvcV5xMy1Z2yvzv9mqmj7AiFwxposrR3NmZE
Iba5Lz3DxuA6BFxm0/tS5Ge+sEJwwnnjSTXrZihlWQ0UVy1iE8GNM8DoqU+P54If459y4vE/6ir6
SdyTPY8DPBsOr2AUrYa1A5Itz79UyRMje6hVlr9sxvGnx0QU8BNNrgjY91Mou8Gn3MYZapjFjqEO
uUtuB65BdbRrL8rgnEsJz22V5733w685d1CsM7Dyxy7mAPUXCpsbhrTojvJ9XTkH3PxNJ+2Z0aLK
QIV8+TmXSKzZmiZXM/pTo8SQcwx6Int9Jhf8cI39WNH6rJL5VV9LBKA0BYNpJ7JRxrkHaZeOLelC
ZUJZWM0ln7c62+6v+AjjPSL0VhtNFZ/n9KobFvYbOQuND9vHdekAuZ7nMv2ciV7I/MI/ya5hxAuG
AmDd/xbo0fitc7IXK4BQMnCtGc7uYEiDpuaPTuVMw2PZRy90k6PHczelKWMeG7lNgetKWzSJYB2+
WGZRKAHanESTVrtPYOk7inBXH2xmqte7fsD9rNRNSatH4O9tDxV5mYa//Jw0uHvkAebrn8f9QvYS
rJLeKbfj5aBunhwtJZFMD8EAWXzhKMbsMCuPC2LSbfHn3MoaNqKvHrX+zNf9+Td8bjs1abMeeGU5
3DKdTeYWWkXZLPqtv4HRyx3jBtj8ViVAZS+2lHzP1eFTp2gmvmQsd3eyW20zhUky/TTEeidV0ba4
n+Kk6k0gcAeDVn12HGYPyvH6KhkZcuhqM0y5ETKua83a1w/rtOqgiqH9/BEx+Y7wQBBYIKF4x8oJ
4BQZ3K1poeoJ2ePEdut7tZo2dP9dLf9rD4NZxc0CXu2GBqOC8pcx2vqha0z83xUv3X8ypvj2zG3S
C7lK9T8OKON5yzpW2/4V27nFl2bjF+LUmGfkQpZldq8WK4gf6otKuNVyjemOp+bJIIRGL4TB/FHr
mDaw0sGyN91pY7wEVsjzPMq5ogsglA4D39SrYGpcESRdgjSB2XRz8ISfKscpWl6lqO0Njvl0o9CV
yigByD7Es4L2oQarl3ZlV4cdjnJFe4R3eu1IQHVJlD6euzRLajSG0strw5K1/qby1aNuczROxhNJ
sSU6nNc8E0IkCSo/L5ed7Zh8cTKoCewp35129HgvCYh+AB1iH8i3If4QH1vgbbszFzh82m7JAJZM
wuWy9n+8aloA6EFgu7E6nv9bPkP7+3VYOl3S6MQF/0swfTy5lJrRBee578QH73z2awnyGQN8vAG7
kFEtHw2Tyi3WfVNe/dYrMe6Bu25+T2yu/M36IWoyMx/0knGuslKzAN1bjwfH9bT++IY8DDLgH17o
VAtHvehvFEixAVD76bsFv688U2Fe4lgdU+iiDAlNAxbvmLbrBo3gDZ8PEQpvMORusY90MfE55M03
8OEd0xOIZWUC8Giw6p7U920KNwYYooc69IM0pmwQXUQT0TFmHmbxhYEkzHq6dA7DeM/3OEPA5BgZ
KMWz0IxVWlCK/YVHKClec9DejsuCzczLmrT9SVwo2rg6wId0LVipaJcxDCutVNFiQZ15lMjRXJfO
xpdbLK8/BA++a0IggP1u/BfczG1V3KChrYs82nfez3r9pYujwXQB0mB9G9dNpDHkqJy1H4syo6Qq
UAaebtucWkO7KvfTq1Q4/NPE3CZlBP3Tl0/Cvc19+7W0lCGnu+1cP9shHJE74aoJaEu42DYgVdHf
quP/E5EL5ozmaPyM2Q50bSJRe2943NzArIO3KuCv4KZWq4bWtR/EN1C9He0FsXy6/q2F04h4k1S0
NnzmPZhmIajS7W+F63uTiUuBymT45NIiJbyJvIgjMSY6yaUhnNNBFNd3wV91gu7FnYNeRfmJzFhP
gT9yXg6yY6XS3Nqh5Z4tLrmAcqfPxr2BGszDX68tYHE3wVmo70y7M4hvAqhkcFUQh0bqVK2iTszO
CBXuaCIopYjBvn+SgZk6uyy82vzcaFrgzeKFVQO+dHJhU0Ozv3auV0qD8dcIF8Y4uBWWCndgLcjp
0ngLnHFBVrDD7EPgH9SRx/eUMVaxzhounGiR0ukVd2HiTsi2kz1VFbeMzUAyUD3IT+jXb9/a7PSI
04Bl0Ap8PF1hvOXoaWEtaswfXCZNONyCOmbYijsgtjStBPA9v7eh1TRazAGn6IcFnH3r0UJ4TwOQ
DO6ZApHw6jw/859rvs1IaGVz+lIQIouMb+Q3eCGDfe/oqdqU9J8T9ovfDqGVgnLZUz+ksww/B2xd
I6iT4u5uLSJgrY9B8XamTg8WkoFebPOMqeS868qAbZ1cDokqKd+hdb5Iu8MIE9Om9UUw2VUgEN89
wut8priglVf2+nRwbwkS5kkzM4GeimnhomwFiEMhjGv+bT8xoyR4brQxv1BFhxcYzI8Un2N3Q0qu
6w3PdBZN5E/mZtrknMX2fiNXuK8vPvAHIefwluyoZGaTCFX9N80JtRA6/aSkcvJkOvCKE7cAm4bs
of62owHJnJ3suinWYPULvenKE1uNJchu7uVkiObXr7Ezilw6trs1faUaOnklLhhVuzxolE0cgQ7+
95EU/VfyGrC7QTdpW5t0nvZabVqIG30RSPg5BS5B/HjUMcIhImrdGefjebKAEnYpyYDOp8ujBe+u
2OECZPLiMbn0ot31J8mUeJyStQiExFrZPQgvzSj0dBIsAkZNgU3mY5oC/6/ILq3WnrK+sBmrJymV
btuyv22XSPCeormxtAp4Ia/T6HRpTX8z9YWY1xNoeJG4dZXg0NLSz0tloEPDKmFPOgq7jmJyXBW3
PS+cAzubXxGa5SXUHKosn+ua8JAeWK+hybVUU6tfYRm7wbvxiczIXgYzyroYtiijptiKgRkUpwLZ
HUDpyjSEXKzoydMHeybL4mNbqs1uFs3xtXhyH+RO85kjiaNTemnnZP0nM1nGVAE1oNd8jkddgL5r
KM7OaPX+wJm9nZjIqiIW6041QU8nsoC+lXpFsZG4sfxUvAacALozAZtMkMqJd7smmClXrYco7hee
xfEkPPRUwWdQ3SiP/MqFBhEmyiYu5Tk5d32PruOhPrQH4AtocH4avjdrZXt2WsTZ3KHoGz+0Mv7T
rDhTCPMVqazfdBc+bizm/4aZFybtDByTMyGLM6WPXuEjizQY/TUjNd7QbzHe3p27WHcOWeyaznkj
GiSUgIei8ED66Mon4a5xyuYzR9mCSHXI/3HL4EGbSxuv0BnqyahoJesRwhtkXqJd0JBeGuDRBY/M
RfOZ286VmPlPfxJfRt/CDA+R3gNeQpQPZAILDSbo0ylJtAScW3TMnjTzhFiXzt6JIMKzPz6NRkoa
Vebz1/sf4bPE69aAZCoPmLP6S+Uccv/+RDWg9lc6prCQgBGRCHBf9+Hn01lCpPDL8eKQuWIW7NYD
DqQcWeQaXmyF5JBWgGIeEqvm6zmM/lf9FbX3jdpqaZ7ppZQJPyx2Xh7RNvWxr/t3pw7gpEAD5zPK
MUdwQDUfV9D9uL86dnAWhLenx/8kS726v6xHiN0Dlc8ugD2qrXaOF0HkVEBx5cbzKGkmxu8fSZk2
nEBUjQAbkwpuBit0IHpAe6verLta+QPrybrEBiufAYPRXvmZYxaq5YSSURsUn/l5pbaBRBSxuK57
Z+31+HubIyXqckJ2qdVlL/lk2dhRlg5D+N5qXAqU8ZLtKyQwAP9VQ9UO/Dc+gJ28EnC5ORxi3f1H
CaCPEux96++VHt53DU8fD7WGx0e/QDyzVpu4fKcvgBA7zhxinHcbGjIdDOKYWXlzvv6RRs23zha/
pO0SJmvhKgwtR1jEmGi96gCTz+vRY3GqKS25rfkPGMc9rEQosO+WR1wVVpa0Z1AV/1+hst2Jj1Pa
qOW26oZOO6iTFPx0uFMf0pRYHQRb22tpIgbLnrZ0E7Uk2lo0UmTgyRoZht9Qyam+QBT50FiYOAYS
tw8FkOxhQChjWrf20o+4YXDKow2ZmWomS5Zez+PbfaggWCUWDKSHPHtBy+5GfzSMKfrpzeJ0rN2M
QzUX1bryaS3kGdnxQYcnk6BHhD8oLuZ3dS2fEORvrBuGct/lGRG4YPJgWK/B5grGaDpAIPTLFAit
RkfxfdwLCLGuXtBnjHnMCYM851/LWMEwETBnNlqFszYBEmtCb7GDMSryWHQgnyy5aRfNOmtT43qO
E0H0tSoQVD+ARVwzvbAPqj48q83OKJ/co+qr++LvXig6HavrL/Sp64SZOMNWFFJK9ZyTM01C53pq
5n+7WynCJ9IPC75m0mwgB7i4ZSSf2gGhokM4nAE1Z4apS4TwtMa1ukDleeG3SNO4yEFVafyMUQTB
TXPGfcJlRd5gxgPB+sNPSBCNh0E+G1dJq4XREgVxndPcZi1BFWmy4UjrN5iADks1z09oHbyr9fgg
qzZn3qxTQ2tLHKz2b5nhoebhvHcnPHrvQjYHfoLZPPgn6DkE7M7fTvd41EauoX3npWOLoYBUz4BL
mUHazHh7a3VG0MbH7aWEKIsDT5at5QM1/Ih1HP3czso3sun47k17OuJEIXVuLw/iHirA/nqnnVec
uQxJ3g1ewQQW8sZyugTXaPkEdBUS5AvyS1LXGakrTNHP+qSOZOnYmqfXMjKrZJmpaLcTw79AEj1H
q4OnN8GYd659pN7HZ1PoRtQ5G9cCWEIxu0Z9e536ORLNM46yifo0y+pWtmUu1rPhTaxsKGqBRu90
e8izTvJE51D+2tYst3vmj8N2A7PtB1wVjDwapT6kb4IyQNMivBdBxWGd8FnXoAU9wO0A4Rcr+EcJ
3qK79vBvH+2+DdZ8Fwo9/6E+8G9j4Akf0daCnC+P/yXYQZ0q3kFo9qElqH/M5GyVv5I8RYmxSnhG
XX2R4m4ZW3TUJWM98CokbybOEMVqiTi06gK+KhpteQJxy2ecWH2qWjS4RBHgWmmcuf0L3TILlMdA
GmruHBUsFtqgmVfU+WJNxLpUoJTIi3OMcBq+YTOFZ7x6PlEsqn5OY5RWXeUy/XWLrYP+wPYTkH6e
kw46R14me9t5tzukz/Hq8QTzbQlKn6B2G2J5zpBB4kEImrPafdmAeTIBvSJqFt3aU+76kf/A/Nox
1ESLUbgMV5NZJl9kpqKQSLGQS9g4NSvCN9NNbpdc3Dn2fX/4D0/Gxbdc+bcNzOR1xQtdJhmj67tS
mc2/bY3/ZSSQKv/N3AAcSW3qITCpE55eKPFtpXnH86L7DHlba2rTItt2ONXW/UPdoPR5tBvTFqUu
H6Aqip/C8kOywRjMOyslkRekDmdGZyKTLD8/yMHySVrP/gz74xch6WI8hOCrO84eRam1nnLTs9r1
U0PioDh+r4Wi7KeotFxsGmEcshyYp08G5m7xoMZa1+YqFz2GGcigsYgz3jlkt8tyjXT8sEAQae9L
3ZGgICBQ0pCj5IVjdPCfG711eajGXuWLmAn2qz8Q4hyWz/S/mdwUHR9bwkieMc5fZE10MYCNjTYl
iIUQxd7Ms7p7WJdp6ctksxggyuAqjRYeykl45Li2bEM8hT0T3oLk/If3jY9fyMlKh3A/ejJmS+N9
AwKRItKLV5O8ghHS7tf8BrvWE9cSKmJUGm9jftjibmiOR8nitNRXhni2GQKnFhKcF1EnV5rVKCnF
ZscNXwgbAbVRHRcrT8jd4wrxAsncfNZRz9+H26q1mVkxfCsHGtJbWPhqIidTVGXqQUslqPesGbnA
dTHna+ZrX5sbBuZW3y1DGu2/TlhiT6+zxlr/i7U27pVWYmM9tkoYf6cYyxHxoHZS7F53MNQgDWDW
H3T9AooJbHzXQOJZpcm4aMtjqnOkBWpD+8GZOnz3+sGagS8qt1DfC0qcQGThQm825P9Cink9xHXW
nJskat6pCJEZL4hnx7hRTTuJlSb3tuy/Hgk2Ctw4lybpe59T6/WLnzUS2MuBdv2z+TutIIulwGdg
X2T/24gyWkYkmgc6wnSdl9kcj/OzkrvMp70ZhbGRb/GoE5ljwuPwd6CLdssTitkoismAWmBvG+1w
MjKIsnB3bhUZtfRGGnjfmCHaOGX6zAWH54GAEZafAeHF1dQonvpF8HiKv8FxhgDLBeed2hujYo6e
+r93dcBG/z6nNXzGn3Wetl8JVvcutl+zXT9BQQqNjnFlZZsrAi4/kNPZeLg/PmNKEkDljBVcn5dF
CcMUl8U64xEySWpHOp7RTwSXebGEal3siw0mN+VNpxC77f3Gj3EPh2npz7XL8yP+ESrlsAmQpBhn
fyCb1gfxaBnDGgchKag8wtMXDyAxEqT5KbPaUNdEc9dff6PFMisDRtjtxdIJ4txj+wrIfLbLNFZF
bOBMTRLzBvrT5NdHwDfvPyMybzT8Oc+on76TZe7ZnVooFTpI3RTi4biY2SaeEq0tMXiRsJabxSRk
42VhuOZKms/T3PT2Tn1SNnCzwj/Ya5dKfPGaXIWChQ09BJxie9BTfj7PpVEC39WRKMtFT+USlLeg
Drl0op/6A7QE6nEmKopK3mrG2oHU3Ax107IVdDftDYnfX/GEPNMDXPQJKtL4WqBs2GsjmIcVXcF/
HycFjx0PUof2//tcv2bTh8N/wl1OxmVKqA8ZZR0rLwBxabWJ8EapFko8FSt9tA7vE/K4cVzdaCEn
p+IL6vyyy534PLgQfxZUw9Mqf/H3HpB/0wOWeJjjRi1Sj3nceWmDw/vEP+jNBoVy/FBDX+7XN16s
CqsF3Zd04Mo5+qf+Y73mYy5upPyF5k0QdOwsOvWKIHasIPg3Sb5LAjIdqJsjxAJ15I4wlhXP/bhb
wLbej922RI7ibKygiPeylAfhnZc6+9imbdt7MpTXTkv/Q2VGSAg9djFUHLfF4IKjJ/Jm7tEVfWf3
f0yABzlv7sV7RValdtryTgHdy8NVZ9FgI2CFRHw4P+1GUA7ID24JRWTRz9V8EXlNnL0XQTkqa15b
QKOS6wWIJy+lHJa5hvobMNayN29tcNI1cdRrAA3vBSXOgmgZ8Z53/EIzy7kNYSH2SVrvXWDeo2DB
qusC2koQgizMvFsWFEyz7iyEHG0cg01lAAUha20eU1odYosZYkypLN37RvT/a1NxGTkJ5bq1fQnX
7/KzuS8V3m2pDLBr1GvIvTss3mSPTPZHxUHcs2GyZ2vRXXLSlrGqP3i5lzVHle+kLHzGGXkobK3x
JCDVmgEIdLnGNh2w1/UNegY9f0uzmNIb4bHk+/xzgiHVBeQleTlpQICREOoSQLgBjZ+0S1SgLcRi
ykwCwvExE8zaF9sp8YMz2Zd0OQccIIRFBq4rSpqKGOuwQSw7zocsmKS4kE8xosXJ1FlPxKRcHkoX
l+ZPODyu3zw0OhHsQD+siOl0IboG0+vmkWwcnXKDkpsSUXxwJHQa1kn17ZSBRoX+wu0V9WSrsTgs
p8MdRPGBy0Z9+4z6gJ/6YTFxciVRr+sCdVIetwanlLjL8L9ftsvARS3uELUXoydWatMFrkPnOlfY
yjCsxAIv4HVH+fWxSnSBBSiq2JiKBaGlufX3rpEzTVqbNOwygNmX/tg1Zd9GzF6Odch/rnTXFwIX
mwSrmOaTsG2IVJPPeZSg+jlvkfEp9I9x8A3Wdas14RT+O8VtmjlWD2ewdfSihZ62IM8hmpXuT5+G
eBM3uNfQA88vdrOFNfTTbdXNPJb6Un1YDFRM3vDTyiW3D1ABm66wd1xGogH6ig2iS1fdosFxnXl1
BNlXMmoi4LHmO7Sueh42AWGj8bX2JpcpKDiy4ZlhcLQmWHec/ZtD8NpcwKLQse0W+xRYjL1whmbC
yJnuzdJ7c2ZrWnkCmJusVjSi/l8O+NciUDhC6vfdnFffr86b0wHaJjtVmezL22osaPC/7CPgLYDA
KsgD5xoTajxBBZVj/rDmu3UaK7yJLv4qWNrusOH2lMtgjru8cp1hWt24s3UcCLMhUwc7haLo1dOL
TlloC40A+PyJqDT46qIDI2FWeHnUGwZqqnOW/RwtkNJon9Chb69G0maNOJ4ciQbVr+LEZ6zghC8H
AonL1cNy0P6gYhpQ3QnOk0HbaZyKIlc5LsZorBs2eg/Sfpn79flbFQeCfxJBHDKd7d2qKSezV8BD
fMvRPTFHDGB64mTQXFVK4OY5u4yGrZPdUapk8ajAdk+pB9QBs5Gi66gACDRd1kBnxUecgikRWUE/
mptDjBEecA5jIw2mvI2IX8XZP2BqP3YV55gBZijYCQXoX5DgslHe/I1OiFSMfW4B8CGipogs4Z53
B3RFdKNsRQHIsnYsN02uF1Q1CcQb5wAGLftwlySu8Q0dLZOCK4jRAVkQtQdLtw3XkVUucIWKga1V
F+b50wljiJhAix0+x5g8uXT7H2lLBhjHMiBg5NbSW+Xb1JH6vUfrrcamPzUGonWUgfqh7OpIGznr
DI+2uEZHXgKXeLlx8mDqLJ4m3JbbY4Gj0xQWec2JCe6Y36PzVNFq4O2DgcLqnPFNxyZHVHxt9ltJ
x9Wtcms0OLtSWA/1IVFAF0o895waSGj0gDRdw7Uujmk2D9Xe68kd+PfmCkv6ygY3/UKIX0SwynFn
FM9Grc8zH/826yTVl4Dx0It2ZCGtSJ9GmjN5Vhmqx9cH8WRPhIrhSb1JdGz/su44QKwKn6JA+oTh
g8cZrFRlbxNghoCG6e7GzYHOpFg2o7OLC+oKBCWfcNnE8bJw9sV1a9avD8/aBTb626pBR3cEvgMQ
ALrKVUHnlX8d+Pv1CxupUMGkIMeCuUSfPBKz9yeWv1T5Nk0n+6n9HhbWJIFrDq45BowhaR4jD8MS
zw26dllbI5PbzdsTm0orsTjict3nV5JikA9H8n4XslSXq3Tqg5+QQHJpdpc65HuAcZ9AivGrePrt
CmoAmBMAvFfjv6lHlrCIsYnaLaw1SegVM6XvoRvLu3CdZDCi+IwW//wKwc/39cDYR4F9jceSYzKF
HPd2fddsrMX4mCBft1PY5MAMZJHi5/rDC7QnrUBfSQcWkkSh0R8X+doPh5Qp+G80IxDeQjYHNI3I
9BM8LxPdjDaoCvi0vl1jsnHSj7qB60bqlm3XQ4cw0efCNZHujO9VTJGecKkrQUcsiZpUU3XFGrY9
QN/ZEwUzbpxtGsdhpjkP4sAToffFfXfu/VMxXGBb9DLoWAemX2O6v/V0CCOncZyFZrIEQHESm/9r
3sh1jZ44OodTWlEgJyIi79XaA+2YvAbduAki4ovxt4STHytne6t9iUnc6h9HfPtC85BTQ3zgBScP
mO6mMb4RjkfY9FwEqXaR7+/G+2AvHukkRgSVdNKlvsEQ57Aon+yR0uMLQEQiJohJsolbgXtZr1me
btsTpEAtiTMOwaKVZeVKdbzs5liwuWqZHqXgZ4GkqEO045yoeFkMRaROuVK8k61q4dX2d5Thc3MW
KT7+ayha3S/WapD9biu7gMsXTttCfOcvesYOM0DYcPWVxGWKqh44nDnbQTicY00MLzeRVqsTLMuc
kzaQnkhjvD6fAlWWUtkua2pgrOpnasDn+jWaLXWuLK1mF1PJMIr25YPh8FmD4E1hU751/9XR8MBW
zUZT0f73bU9AIAKFfITM7ZAOmPh7gM9F7C2GpQ53KZ1q4zsCkujXEbBFBcfPnMSZrsL9K8N+oHlR
xV5y0xE3USqG4qXi2E+XrrPLanUqs0iGY1FQWRHeZ3MX+j/rPDUQU+ruiBCRjuCjVdXIExZIgNuT
k40ahLflAACSl4+A157pVz6ol5A7EmQxSEiz79CwORMfUtWhN8gdIliErchGLGHQcY0f/XCpmRrt
XyXjv+rJ/go5m4qFG0BW5KB2A6LNeX4EHPBLRg6L7rRxBrC8bEibXvSCm54sL05tENHbKXPvdWn1
xANrUKPuWOqrQI90Fvf8yxWi2/j1NZCK6KU2YYPAihBgt9Ij+z51iVoIMCKcXrUnDm3rN4mxK4DS
/Eb+CNU/p4F+oZFr/lwj4NlkKliDhSqHo46XEe6k8/3PDwKfutv3Cfu2Y1V7gNU2WyOmumygPNI0
P7IylZPYyNIP6CgzTh+ZXyc2oF2sHy+3DqkjU307OeMe5gjOBdSuPfeYEtRC4va0nVhU+Guef9Gw
PRsihf5T6HZUzcMvaS19dvbsoJ6qtWtz+DxQvHzvJrzHRrP0GnKWlf+axAjcW/uxS5p5bhWKAS6r
oKmEGAyN/c25Cmgr/XhOyiXTRbqhRSIZuqNKSlzuilf24XoqVTDtKyrX7+h88cpGDCeSmNBY3IVN
9XvCx3S7UQG7YqT1QPBNpF/JVAi19jQn9uClIT4/uyxDayKZgn6Zoxf5QjKDS9QQ6ZpWL/n4+jl6
pBi5lqV7gEX2lOUp2mw8isqkzQy1TQRe7GAB1hPR1398/4IktgAVDnDAVImrL3V6i0AR4x2LlAhR
1NHZTRmsLgAkT9yjmD2ThDKuJcOjv7/C+/fr0riE9InQsJXTeiUwRzBmKYlCLjfLGgDT/oVkjBR2
RRhSMwjdbBmlVR+EuJZxoESqjxP0cUcXaLsTvxH+3luuabSps2EXYgjtnoY01TzL8+gbivZsV5e+
8k4KLB3gMfB25d/FpF0avNn25K1Su6CLHXXqrC5emaokt8AJshJbr/T6aU5LebwNbOx5DPl5VQMn
m4uaijbEsn+PovhjDKC6rPrpPf9zE6WbnDHnv+FVHtzrj/gf+3GslgnVM/k3YbLrk4dHTE+L2C3y
wEVZwUEx6fUFdTvfqBE2GIKb3poRbp2a0N1smumbfwB7GXT5hMrcJg1tuZaMEoFBc7jhLAihqUMR
ssPaj7HUmlTUmEzhc7PHXfEaE5yNZ7ZvXkqxBQgSbIaobFu/vJ6g7CeNJHl6KbqFSIQ9bO0mCLK1
4nN/PxaxuNFqExT1tO1soyeO4OoGnvbFccqDUikCZNnyD7D50T7ijYTvMjSI/HE0ho+HwfVyZjPG
x4+8xP8y2mKy4swhlhnkulnLxlR99nQ+rl2oqnQPxrK6xa1kyW8jEOYwmabMeTYSuuICWQSpCN6W
slC58AToaDmnA54NnTUcQPUIWu51nn5ZdZsCPZBPng3LMaZFwl95UDtEjK8yXkoxNCfaTuWtNQxP
k56t5LPhPyGs3ISJGTIL8I9NyFr1hsKZLpPjqGgnrDKrTxFn0omj5bRjKb0Tpk6n1as5S1NK+iId
aWIh/w8A4PreFXuf0j9bshAOrqKzvdESLZhLMPEqhwgHyx32O+4xWb545ti6NA//X9upapPjvpOY
8h/OTnsoL/R0jmC8YAtpOPSAcNqQhUSaLbh4ZfC5uoXqJUi2kqr9C4SZJfkZd59O1sdeIM7r+U+v
RDDvGJX0wIB0xPFyprQp9NDWivQZJw/6vRApawAk8D/iudaLrXnIlbkwXwj2+hHw0zUVrS7CKl+U
NhJO4aXAchk6opKNG0u5N5+af7fOU4BguRM9xp1wXZY92L+inKvqKXweoF0q7nSvxLD/hq3DXFG9
P2RAvE/5zjnzbptwUxnNdYIwiiQzlyMmoSDjqrMJKz8H02AL+O1pYS/6dbpYdhkDCo9YVJRza8u0
AQ9qk2+wLl4jnL0JQOnl8Vs74zd2L0mC+vZsx0e+05ppxAVLGZxelgVCkIdeQ+aQ0BwDOijkL/nl
XW2nvjag0qKio2kORlJTA/jCdDFSj9M/5ta8219ys3CZtRD7VUUylqoYQJw5nUYweyzxHCa67kre
aNGSC1t4l7VVBCXfKeqnLOm2UvDnnklUZoD9R77T6Lqi/k3/J43uw07/e7a8Lhc7oUOT/x1rDPy4
GsSAFykssUN0nqe3oRQU3Se7rf3Dfh4gRgcvkM0XLSqA9j5cSDihNZz8XwU4CNgtIBRIDQlxwIwe
I0z42pReTPUC1UfkTWZgXTqRTU5eLRcWhsAqXNZ+TmqpyofCWrQWnRZkXKmf5bD1f6G22GX6/+Vx
Se9iM4Oqs2ofcZi+vRGS/CiBXdGjIvW2EpDO+Cqz7o6V88MEfmGXCMJFpyomoubs/GkBlxwMfylJ
a2I5nnxgWOnujdp/pVokGbZaLUuVOFvgW3lurzGAsVLEk6autChQ7DYd4vxXFHc6z/X9jJwlQtSJ
jd33gL8HkfJ1YGJhzKySU9Haz/vdz50bvSDUxFcbfTJf07ZUylKHACssWDHeL5TGM5t+fRaD2LyC
EdWTcvCzgCDb2tANZKf2muGyoj6N5F0WPDrefwdF70detbXivdO4o/Gv7yRwGIMlePNaZqWWKOs8
GgsUKnPwriNpDGxad/pVqvgZ76RkYel9vfk7cn8xgJiviKw9OEQRB6mvaCiJAJos6w1So2jAawU9
leXZcR+74X+i9uO/lEDtKme9fttx6eIBBTOd7JiBouL+apPesis1dsquWbWzV7AIdneV/ibHV4+B
rtPaHxaZ/tZhsW2LEoGqi17AWZvp/PrYCfSk/xziK6L0cvm6OfqeVe1AgPsN746IkmCIsx1Td6qU
NpfqY7R3PV9oF3Yy2w7ZZeJFNCypEdV7Rh/wMjqoUPWxqpEY/e6hQgMXZkpsk+TiHg82WqGsl10K
t4v//qqgP58l1k2eZ+IZOyEQ5bFwx9+BAiQ4QFMZa9sF70zzuYDLoNbcWS4b4V/rd1co267VQK8U
UZar+QsYAEj13cbFaxfEe1ehdGFvLbqFA5EOtnQ8jF4cSdRJ7PxmvR/tg5J56bsuN5k8tidOaEtc
MuC3FIM0soXI5Wj4B6WT51leoivuww/gB7HTwVZXkbiXOPxfkxobkhmyQbWiyLhpxjG5E+Bc+th/
abWtyFUrhTeWBBXHftgX6N4/vTUNmtjj0cB/q+nB7nQ6f254jfG5J9LzU608l+XyzcYdiEFFzTvD
DjxuOS6lpfc98Gz7uGv3ye/iN8iGoV2++MpwYmVmxSCHS2z3bxm9mGjROM3HI/RlZKNfuL4VQqMc
rjOcZ8SUWwvql/bPZL5pGqqEGX7dN33uFMfa9oagKsgT367c8fUfytzXGlMeqfxT4EAjCbAi79to
ULYk3C0tgc9AoYnV18d5tSSm1vm0xA1yeIGnjF5+2ve5y3NHpjVQCvQ9Yg76wc6YriHY/avhKQrJ
TGM+IzljXOI8JHef516wXeAmd8h5PT/g+HUG8L3xB4fSY5MTD0XYrf1YUdv1YBCSdtbiuAQvPgHJ
V4lFb5L6FpZJlL9kLEzfxBSdEdI4TH1mqgoGFbwPCMOYop6JurzucO8FHf+RE1NcjV6lPNOcsI5X
ii6njWs5KAJ87pz6LuNmYj5daPbwYGx8wTjsI/vJwSLw8+KvHPepiJLgKZG83Vp8CHTNMFYVEeOF
n/HyvA7TYYFkogxc4fHHZcd2F/2mVxLQbClOi8bMux+8u7fs51X7NTomMtDpmFFBAhYOlgI+kcmX
nLu+Q8vDSWVJVAgGGTeeW6wa6pE6fAdMFECgThHGUQQxpKkBDAErlvA5jF388UWwXGuAc2QgkEYr
hvoC5ipdvupT/MBi6OMXekrt1c7jD/TJYnM5n0jRhlaAxcbhIad3nswmjvfCDB89Lbr5hNTWmmXB
DlX2+PWk9hK0mB9IAP7QJecCx2KlW7T+Z1Xm1SOFtDqHWwhpfro02AvF6CE+4gzb1FhVjSvUxSWW
GBvvUwe48hC/nvF6cV4eV8Pz7ZjVmSSfVE/PzHrx0vh7QI7h+ckTCO9NnKNQH30CPp+C850LK1gZ
+R0A47GzpY5hWzktboIsmPNMZy9lPLn6D7stXBLD5Ce32eSiMS04KWkf2YukdOV3zd8G/NPO5VTH
ux5T1CsDWv+neyK1EzMmsmGbIzvWeBWQNceBCDRN8U18p2jvNKflZvYJpeTIIUN8VaYYko0/bCmn
vj2yNs7h3z1GNqQSalpm6ooCiZcKIxsDC6lzCjQbxgF13iwVyAoHPOJLzjF+Xm/unnXs0OHjMjSX
jxsqcZ63796Uqv2BoBeKheCrOSybTKJe7uMKjE+n8ldqByVqXxtRXH9dNCQpbwoCa0wCqPOmK6ev
NOxsbc3YLIxsz2gxPO5RdEvv4fGauXGTZ3dnNo4fe7RObbJnZULXjobs6RLCFaQmdZ/EfQv+ldo9
d652xYZb1K+se/hlaR/qC5lz9BX5Xfxe1GMSTVNXaKOQ2gerulQAZHjzm/3QAjysz2LlQrOtDV6K
XzJCXeY2Yzi54XNY3D8u0jiJKwyh2mp/KL2ayV04wPgFs81YqazVe2Lt+7e2J/ytE5abDIh6r94F
EthnOeF3HRJtSM23xYxooGlE+rxFeblb7g3OMnKneIwz1KciFhjS67joacazqNGnnkIhExEzTobR
iKE5jY7319IjjDci3ZZbzl69LZvkwfwqcYfWEMa6mEoxQ7qUrG+idVk6qw5SN7vVECB7ZKd4EKNp
tHKLL4GK8DvLyowjsMNpgovRogitGZvxjvE6XDs2WJhBGcx5IbRiQwN8UHRklO+6DI/nLfiLmw19
qP9E9uOZ9dgSm262vcHvsGngifeva5Dbg0nUm0faYGs0uwPvWcpRr9l+Pr/1HktiziELPIi+TDnc
o0htFawF4qCIGVfjeXsaaaXMpUosCUroeV/LeoMfqJN/nY3iFQD8v9ZKUqcMRhjDnHAs3LDVIAqH
7aER2ybSDvdRRSpDakZ5F8YhfYJe0InvzPx9qqdtjj2a7M7PQ3HaeUFjUIlNruYeluxcG/laL+6k
ORk6Mqf3LMrx+KJj2NxvIqx/FyEzOxIWkZHoBbBI76Wm5ry/2IMwe99IAGapupWcLBbUctK3mYNH
tZVSG2Y53kVO5rq1iT+b6BB9XPUDLEaEns6nJjHpxdfIzR+QMiX+AoOZ6IKDqNAG7GaacEQEo7LS
E/iHzwBLxj/kD717rYS9JFSswQ5Mxbh6VRtYNgms8/MG4AQ/0s4wu6r/d2hIdz3IvHMLsvuwfZF+
dDYgXeZl+y1O2chIYbhpUUptYFV5cv+JAtFHomSXzvo07lGvMSQAkEmdy6hBFOpufIC5xrvt6GI1
u/0AOldwf9ooOPwD6voE4E7aom2D9M5xUa+zgKEjUm5ukkT5cHPl04C3HNi/pZZ3zVszWR+J/qLE
9QmIOKh2a7gntP1DTAG+jIAUcV6fmM95WrVKDh2RlPddwL+Te5g3I+vTQ8ZNjK9wbpab0To7z1a8
YPCTgb0JBOwZyzsn7v28VtEQq/J4RRg6x2y6DijZyZ/K6K3VhTeatH1s558F/8Kbleoj0NNmQy8f
3q092lHvpd4OwFPHmF2Y/9Gj8UNm0Sc40A81SsZwteWO+eAv5+im29I6ZfFEbtQ5zh1vx2abc8D5
5+F1k3N0e433VIDO+CYl3jTHNJKBbOXyckR9AtYurVa6C0cybLa51iRhjmOKWhBy+NgZlNGeFmE7
YIXD4Pa4yT3c/4f/tjhYWHLF5sPBnG00YcjsL5foWUTBUEk58DaoiZm6MC6HZIM0hMPotG7//lQi
vPLRf/xlu6dWnyGbfDFgJ148a2J7EMq/KWNHIfiI3KU/m4IvO/Nc6InmyFjGqMi6X0BrsfN/7U1K
0YpEtW3siQRXg01eyQbIkXAmUFpM5gbCn2v34vX+v1AVv/MipnVmPthIJ7MQdmp986v40Qu1VB5P
cmYMoynkcSqqS4riJJ4wxD18E7bj6UlzikZ5bxSrboca/PfVxwT3ZO0T4tr7oZRPztFkOFwrKOqM
rc5B5lmt37hPkoDZWe3/xTqOGnoGs9NWNztYC+iM1cWdTHnOJFp0fxYBuqqUbd+mIu/W2dnacgBa
5Cp8CXWO2ht/fJbtFCqdDbzQIh5hMYd1955g6vFfiJJ0Wi9iZEmRz8qKGvuIs2EZlcUnQQQb5qML
iRH9zV/kIKLWV4Isim11EuERgXtw253celyRRTYY/C820zNvGl+BkBM/O74kp7SwtuPeiNgAruKw
piftT+9dTAjucDlFbq7AC6XkPyP4j52HVQuFK5SDx0esVc6VH/qSTwDFu4qsC38SUSxZtPTwTyMI
yCyxdQRLX7BAp8Vpie/QpBVa5nx5ZnXAtkF/K1Wu2PTKO1NV/FgoUCxgc3QPbmno4TH1zCcfIwbi
vXU0ZyUuz8m60HN3d8+gH49Yr/DGs55sYEvktilL43fHVkskuiC+EnSoZp+S+86KGzC7CLEgsFSC
ipY5GqdWg9J6rJ7FZWghbkeT04pLd+7lzTyTWMA9izX81TOn8LrrK1jrF56vQCi7u88fMm9S7gnF
jM4Gae9qFKBBJCei8llF2bMbYyXCaTW/RSHV6mEJIQf/g4TbHmnZz50Az9J4L8Raag5W+c5FWLUg
6b8A3s33LgzCyZErX1bx2OtYU7I89er3jM6VGfCy7hFwU1685klj2nY5oUb9sNh+gknkIhJmVMId
m8DbKY13MDaPuHeHZVF3WDPm3o/DxOHtJ+6MFHb+4J7Et9AECStEMZTWcfiS/B3OlQlp2bkYHUrs
rru5GasEph+QjpmSLH6jNRtiVsq+FBw21fki+r9r1ZDlq6kBqrnRZpSAhcAwNDWWHu2TsZOPdp6m
PMo0hKQ1K1wxBvS3N5rXVUzKBmuVePCjUfBYRR6T3Nf8OJH+KXT5tJaeJ3bsl1Aa3TSSD8g84omN
ijodNR0qz09CqR8NjS7ERDhuYTzCz2Kn0J21tIbMdvN1RJFbQXBoeLL/PVDK78PEFR1C0CPx2Cl4
cS1BBxxrYX4LXZCpye12VxCKXgfdOEUmEg3jY3Q5WAc5sZ7Ld90FLv9C1yOs9FHX1RN6HfUT6/Sc
0w/+8By06q6Y1XGP5dwJHWf9xn80jX0Nx+fNzqrwb0Xz7YueIEXjVguo4WICeIELbtZADPl0EcrU
XBKva5jEAbq7KSg9/aarzU1jDFdj0htCV59SuueJeUj6RwZOQu+ejHSM5duflvT2iVyM1FjZ/ONm
TTjw4138kluXseVC2jiOQ9R2R64UutAtOt/tD9YldN+wJAZ7xVJsEHlL3iljbiuTYtOlHk0X+KPI
cc9JU2O9NLZj/JscK3ZNKa4pakalDTyhKzYMnQpxnfWcCt8v1Y8Gmzbw6lcENFQj3HcB2Wy5CI2g
Kya5HBo2cAb6t/PzV4aCP/wZuNCXLu0vlCMh295Pd2uCw9841I3V3FCtJofHl5eG9bywl+pKftn3
nUNBGbDd8DY7AkaK5hpDuC38J3B1XrCNpl9SzRuZw1ksHUcvdn5f2zUZRagC9mCVeY5FN4qA3xRO
D1EtL6/tJ5UV3O36NWaTLNW+yrt2UBd0RpgvGHtu5byzhUKbtAs/95+kcXmGTpdiG0IBO+nNdJoW
2fxAKoZCySFlUHJdNzMtLuvmHHeNpTBaIOvEkIm7FSDtXg8WjrCUx7NttcyXNa7z8jfWj7BaCU0u
qIXlrr7Dc49XAJPcuePG2kTaXbVTpFr3P52H+dEA4lJxuV+M94DwZ4FmGLv+wSWqk/QQ7Vt8pEtG
VLKGcuXIZ27bsqyYib+yB4xvWqEH/JzSjsDMwtIX+6uJ8SanIPJpvGGN6W91RDFbnS5HGhSP6STR
ZyJSizAiaHnJHcjrf2z1iBmDdwERl6+fQDgFlitrdKYg/ibVdQ8aaPMLEDCdY8Mc//G0Di59uXHb
kJBa+VHyCKtc/amAXt/KaPdeLuUmYgSrLApa9JY7tG3hYU0ztHnt2DW93dNUB3ZN26xXAeSo1f7I
HjWCPrpy5ogsbP+s0E69qe0RIhclBdXYtmZaEU6nQ/g+AbWpk2K3BPMgFyJ3uocQqet4BRH7G7Gc
JahqQ5tGUumqh3q35K+8JQ7jiKui781DwQbFrKqQzc6giKYSpidyWAFTV2BajG+De1t4YNE7YPNN
lfBVA2XfyugfCRTIHV3i7ATLyJq1ghcpzs5Ce6y2JuDfGdBvzjTBsUD29/7dCONI+hYP1JOFF8GY
qO1fskHgxiDriDFbc2HGUisi3JunkruDIXceWql6bRfoBGBmOuVy61QL1hz2x6CdmnJxSgz4jPtA
MGNEwZqiWDWY/ynoEn530HqA4yCWWICY7X/PoNXBVXI8mqtIaE+bnRVHg/ATtApSv1rUzqPyEpdC
nezuvf7070QQwVT3PdYNaS0ZI76loIBUE037FYgbiCZer90KVQqWFWBferggy+RlM5wztK5IV+KS
Og2dAlRBhsMhbqjQjw5L19CEkUAFaW+N/D/g57uCNsF1yGNn77JfVGiLM8+3NOu7SCjE1/NQFLyo
zRT5iLMr+xttgOT9Gl069s6t7dak3ADbxOKAq2MPwtKwv4RWLbGx+npj224d4QBqwmj0zXwcH0dX
AjYWVU21Ph+UXUi1po3Xx6L3E9rEGxIiZGK1a00t2G993j1dZvAIG9qEyj6J4UsqRPH1e0qs7Sen
vW4jTH7v/FgO7NXTWgbMQNgqSLaTThInqLteKrDSCR63eQm8p2b6U9jEnAlBR9X/u5DMWTIgxLbC
zthBjH3PD6BnQ8OgN0AYolv3lxLWW77SEPYrRJVnnVii87UnaYsJTfdy9Uaayse1XZAW/bk8sEDu
lk73eKNsxGkIdVUDFtkmdO4w9W5J/44rZT5JT4aZHukpYZhrXCPJxZE8bOJ65zR8itTVsQUYla+E
UcybCay1mK9R3fz5gl34+w3jEg6hwBbo9RbvqC5mhIxRgk7/wNawCz/jn/kWNJFFdCiNr8TnIpk+
QFCC+1UYna5KURz+6rf/FOYFgRRcAbmxZkuvfExx2hKJcgGqiO4OQA0EDYGVJ6bu/HgMpuUwBvz2
9pPJVQrvXb8IfQ29hMMx3iDpCtvU+tQduqNXoxT4FZacvQbxhr6oj+e4P+8kikJfWTlQRsxEEITy
wF7RGtyQW1CYO4JEcHxbJgJg9nrQ+APZ3AzODnHvnxmzZgf4jSBj9Wd7rcxeOxabTmNiMWRTHdL9
CfZ6mSGvMSEL2kJQ/O8Lbx778W0WNqZyVMkFxE6FbiEPadIkwTyqZZByCFHneg9pfyvw+DDVsKLG
q7wCDhPU/BbzQIALhvHDXE1gYf8JsMXAXdN0vV59T5khxFS/GLDpJy7TQunHtRe8Y72bRHXQXAvM
JzkeoezPcdQbyvkXMKvh8iU7MK9jFCp/UlQbjl96UbH2JpJby2CvoDM9sohhHg8YKwJVxG5e8pLT
ore5UPW95FAG/cLgw1DaK4XGD1X39NQv48LpcEjDuxSqDh+W1EHd7R4JH8OeJc/SLA+QueCjVvsd
4Wm5rM/pv4cTWkMhhyBqXDbrQMx35Xmzro1EB0A7QNg7rL5sIgfJgF+qitzg8DN/ecF2lVzlfYJM
7eFQ3BxGUDtRvlXArbnEzsNrpTWnqIq6Fq0XptinO/4FNlRdS55qXydEiprzwJDCDKf/PjcAjWXx
cQKUB6Pu6PA2ix/Ad2audm3hKClf4m7hZByShBdOYq231mpn1k0oUlW+3ovD3UwRYzNbVDFEgjm+
MneUhSmXSkDwMz3ekgJYwR2BDM2mqyPgraviZ0YvGawv7qCRuOHpMkKYd9kUISpsgaGBZLcgP0OW
Uboq5QIcTff3mmH8DokOoyhcVqSlpUrZ7h/j3reXPYaPgsb4Y82jN55ocxxT+Y5qZZ4d/y3agbcG
rkYHJyWXrziJW5kYCE+2RKJVe/GBN81OrPalTOorVRRgvctEcvcIKX9HyuEnEISi/71soBtwg9Wf
oODWKjlcim6g02k6eDTcvi1uyzzVcYiEksPgQF/yJTK2QAqCJ5CXdO9xr9RAe22nEyg57Mri/xcv
3A71EeMbKeI9M53NWWYgOjPjUI6OOQDwCGMHfF+TbwltzvEYSY35J00olAJfuqTLEkbObn/Qg4La
kpvB4uGlU/vfJoZ89bZc2l3pFfy/t4cNjbITtslqdMVlEKCjODvyWhH7M0bbo9aBHKgp+vHRsNP2
XsR70KaxXZ+MFad0/hKhjhhTQR/mR+yOlF/cvKX3rU4snA4CZ7x0uacj+yT1/ZdXrx+oMTTTEyHF
r/cCxA3QWk1W7TQFLcQsBoy4Fa/Obo1RAktPqRYJfhhU0LCm+HS5PQQi0EMNQaiytGNZLTYQEUXJ
kRY/eNKUaLE2eKytVLPB9gm0maiXM2xRScX3NcCFTvwFWaBFmP8/ifx+XFOu7Q3o/y6jhYN3y3vy
wezWPcSia9+/zsRYtx0ARvgOvqoCazi7UJlRN2Y0X+CF4OTOJeM0hWxRLMyBE+ghh9mtljTWo0mW
YKruxaFUJUeHc8gndC4SeBYbUg1y3XOhk0tlRBJcw4VH+dK7124qS+h2OQ01ya8ApxdmMXYpf+e1
vK7E/U5YOv2atQq7+MJiWOBjeu3rlJ04Lp1LVBG3UQrFZ0+skHZO8rZ4Hn3K5VckeUH9ULsd7Bad
fO0rxZhL79+fjas5lf7WjtgVvxRWJDHXlzYnt6C4zlMbTOUaRWxjAAm+Ylx7JSXmZnBT2xk4LKI/
LsI+e0x/HM5sWtgoCVmLOyMFSP1s7T9dkZdhB9/M7JxYDYdWf2NbjO9E8td3IymU5tKSmpAs3G7E
8uSpgGb7R4809ZbPG8NmT0ygIddCO7h4oIvWC8xm3qNBvohCqI+zp9J36LSMp9rkodz/q7lCHtQe
up4ZwmEHqMdXG/L3sn/rHJgMCWohz4gdKLBAQkOGIhNXiN9u5F6EN7DKzVxdVRC3aP8RM3Uaza2K
q+8ikJC1XVoORx+XS5VpPbw99ULewvPQ44A/8QAMGU26fcsagP1blsN1x+k4NLbL8JWgvo37K4ps
GTyDbYsZ6fU8yoToND0vIMsVVH850QT3I4gx77izb/P+Wjv9jsQmRMmOtxkkZH26t1F4Ze6kkMpS
0h/O6VZnZy+FJiNgeOQWG6R4bCz04uaEGuuyBvT3eDY22+Any6SKV7J9v5hXAyq5PRYow4By/1uJ
y0o1tIm/TiMaspbHayAv7Oi91sv6zxusbQcZ0XXrEoqh/GMPtPZlixR4uOAlN9vyGuGxiwzf/Ou/
R11NaYVo3+KS4ikXcPH59UCyc0VbMULMX35qGYExodPjR0FdyykCsikxLgmsGwrJ9r5FHC68aDii
b2p+a4+9KAvplo1RmhApyWpHTM6LFVE904JolqLOMb7mH5CYQrFVCpn/tY9a7MsRAA3ZyKO9abYk
wi7WnlncGk81eeHLiKo5046Ig5CUhOI0f3+ZB3NjtBHpILvPYSLfwhdcbl7ImCEwaiauSrGFmzFP
3XE2+ifSlVpy66xPgQWYH26JlDSclxsTfTqJUdpnKRInv/3yKrD+97g2QhKxI6sGL+eqFUHXrHl1
DLgzsSw966JGiJKXL88JPH9RmSGYY5zye2gaJGVy86QSOjtLw//4EkoqH6XK4kd35it3FiP9y5fC
WByOqiNRi9m2xf1LskOOAzgpjw12hFwlFdzSSrmssl1iAWkQA9qSyPUwIqq9yXHOqBTgNk334+7X
T24q+VSBE9xUowURxn1vSGiFLSpTWsG1c5KVzILl8SBIxvi7Ii0Y5Kzc+SzMCrlrJEosIesB0zOn
LATH3QBoNEVpixWU0EH9ZS4IWKTdAyeP+12XYjsPc2uw8uumved0GjTg7uox6TQxhpMdILfTTvXU
+hcVtqO4OeHRZgmE4RPYVExI4rwbwBbr2X+b4v0+SEjVHauJc+K/v0/CcFf4oNddRPaE3XJeiWwM
+mtKrmLtF+vBv8u7YAGL5LxhLA5a2Gk/LViHXyNhNvInMN/TalBntvkle0nMDzPjvsh4b1eOSkSW
jmVcunvWK4c1RQMe5orU/QmMeo4qygU0H9tIegL4qvFP/bVujHtv65oOfwk8LCKaCN29zEzxkW/v
yiQOqQ+Y33aGu7vctxSRxpvhrbo7+ZPn8r6JZYR0j+X6dZf46aCj+SOrqSI+tL1TTkQ9KGpbC3oi
h/wOMngHBiohZn8fZYrcYNid9j6Xy7Z7NIx7ytGmTS+9rA6Yu+slGgQNv4jIOgudoblEEVH3AE9y
z6Lw2/4SeTSViBeA/I8aDjThMH47vp6ZQYMPRXeclr3tQ0/a+uXimUDdx0QLfJqeHCnAO+0f2yZH
iz2Ajf0+ha8BxVQcuLh1bIn7XztRMODX2GLqZeyn+Ra+hjWINPkoF4/m0LM8Zrq4I9s7fn2xnRmN
lZORI2quhMh0di9Z86Am43D/Z28ldrESZdB39Cksa4076+n2RWpa4EOvAYoqakMTwlGCAZbNuH2r
D5CY9TAnbmxPnAgv82kOfCISunEsMDunT1MceSaTn86CoUdPzca0iEfuqiiApQ2RfeOwWr8ZXPfV
WrL5aW4gmYrbA+fMvd9euXw38tYcSK4R5hMxcqWnvgp3m13SRycCA4q9kETZ/x778uiEMlmPt7NV
Ois/WCOirPS1UnQcGvVZNFK/eWzuERzB7MYcWyqiZXxTZbjPA93EdTCwdK60bxLIQEFz8HbdpRjw
/ibLHCfV92HI/2CYxa2OWHS2iTyU1LQtwsFTAZzoJCROXZcmJdMCSZnYXJT6h65S14hYCc1E9kFC
fqYJM7iWCm2i3Ti7LaZphTA/W8WSYyUbZGqtfT4e3t0+ENwoWT0cfN/4rqde1jNCpO+dN8ZA47nL
7ogivm655zU/VmjFtWnl9UDIJoiwOQ+IVxbJOdNo4g8hw9oUDCX/YsoLJuwYkYvr43YSC5PyYBOb
3ShNLdGenjxH3C1zQZIE38z3PuBSqKNb2K8ZqEYV+C8KT75Z2NcjJUnZ53xhuTcuD9buh8KTMO0c
IL5cRNTM5AhY6YbEAOrEJTCo6alaOZMAdpLdEv7M5OaxhQH63a5A+lk7ss78yMOc7y7yO1c3fzLI
ch9BC12fx16aNlwzpdGLnIJHmTiS/FrfKqNfDnCplUr/iguiUETbATpdohWxfRJUJHhzU45iIni4
xQx6WAI+mNIoV9Fycz1ullteVPVN3Ugx9qJoh+mq3C8vSdbot0og6OLnT36vQ00hL9w970/WHFwC
bppjHrcVhbZ6G7Tm9F/jPWHQfofjfNsFp42Sg86qk2DlVglxbp6Pimp/ZJN4zjLkH6vKD1z31ZAu
X/nhIfQ+u77jaoCmKpZ3ecvVnV1Znz2BeGH5GmLkJ1l82vJ5dD9KtFIq2YoczqCFNDWO4q+3VWrg
0VOSWVdZNmwovDestwxkFhHNJEEyRy1UqxAamxdSxaVnDvjADAvBCfBpa5DzXJ7TZmJW6Tip9Cls
DbSvkCt/Epz1Bbc67vZMRstT1AIYyt3s+BonmJGKdNJy++SvWIXPHqpoQ6gAWoFkItof+EWzvFyO
bQ0/ySSBmZUCkPsqDZxSen1TgiaoASvWNhUdLOcsjv4tz+8zrXF1pu5P7FLOjjanOBkBR5Uvu2x6
VrKzSo7BhLwTDYV4up4LzLK2+kj0iajhkFZyo4FHiP5YpnxPXT99RH2QgL3s1dFV14BwyLldVLKm
obUmYmZ0FxZkVCk3cSsdiO4nR8G9RFvyXMQGk4rEv0fd6oR/SD5bmpoQOBC0n07ST+DbhvYmI0ew
gfBpdnesPNfj5HH1PaI4gA32i/NV0fYTo4AP8x58pfudGNr5iGvC5XFhUtGWUrfFEX5UErN4SCa0
s9pa1k7by58pSMZkBptkji7+O4V+RHFL+b0cQDD7u39UEI0rb1rc3Caw0B7zQ8pZgdltUBDP60le
uo2qxNjPRvEbBNpEDlKnglcdamLNsP0fwa68Tzwf2sDfdi3FrDnSFnNZVZBWeLFCIlZIK+Jf09EX
DCgdjGvUR+PXCZ7cRcVW6OnUA3V5lT5v/uHcsNYjbkjUozttHRsHuB3ZsiIfCbrqUFDYyFzXjvH7
L4PpoRppn9k72seHtqbaNEafAzpvwqX4vOeVriLkaHDgGhd5CK6msIJ9/UBAuoVhkncKBJHh0Giu
Z64ptDC4P9kD846quJp3vnVufp6ySuun0KWS8DLcj3rIei8nREC5OVYIXdv4I0Sipf/XAEWsIVzk
s8zGwNBYG97v61K8homHfZHJbSXcIdHCRXr1N/yV5Rri1wzyTzHEE+NPUzUqp+5KCtjJYiG7ZGPT
TjxiWj+DD+NivYA61XxfMwFR0f2UxGvVEE2DLYxjt6Ui6BUgY9NkxnMNpVWbo/eucnaKu0fo6WXx
b+ejMY8hS4AdBuNh0tVQZ2lggcdrhq8Z8S109Dk22RYFdyfRNvkFJ/2OkAeuXoN08iU4Ep81+T5K
9nVcs4G27GJ9wU8h8KHvua0OmY3pGRuiseCfwKrswsvQugvnVli5hN1kWqUhh0Mej3PaCVdD+QOC
3Nk/yQeSLtobxPbdlpa+yIP03BcLC/ENjk6iO81nS2eHXAlvsD5xtHwHR/K8fu4Vsgd8gGzvJrqX
rX5li7MXuGzqSMn2j3rZ+LYj7Dqavtobvi+2gSRoGStHvhUfAIVT2ZKgNQNOhx3Zs265EKWnQhXG
K3C6oaWkl1r/GC83M0mR3N3IUTlhjLrrCBVzvPnM8cwMsQrtm0NYrjaagrk2GRhEjIKprlfld+iF
FIOx49qVLAQDCraDafaV4VjtApc8Dr8KSPcEVdxZgdQ8CEdfnFFSYPKm2ox0a1FHX0rOMsTF0CkL
pqkdJvymrYEWBaG/pnjweL8MiUoaIsgxUdEiTdg78u5bRdiC+KJFtLlz4ALit1BFaZRye/lHvjwi
CP01XRdZNWyOBKHvVhcPsa/poyUCa18sKAXlPeDhSiL+s/l/0o02Goq0Pjhzm+6mPPi1eJyF33KA
Nu7NSJbF+X7jgBElk/KDUI1PekqvoYjRADZtkZivPSK6sgwcjn7s4TD4Zq5+xN44KJDrmFLsChmJ
cTTIV1eloPYx+pIsV5O3X+q9+jtzzNIPE9H/IhCKewEDZOyYOFivHbVuWrk0tMGGFw9Emzj2jTzL
bRecQp515lOYsVMRTAMnv9xs5eYMaVu28OAsuzXlDSoy7DuCmKD+esQ/VyKfEdckyngJNU+cudvs
3UHap1Y5yh+W9Dqls2WvvFd/UKoVWmVYaw0N1iNnlJJqrcRwUYxQqV7rDl7mpXFEHRMF3o4yIqiu
8nNHcwxCaBNX2zQBbCRK5FDmP1sZI9ZY2ws4q8tOeILpRZt+n67lj725A+DUkAWldElBUaNWinBj
deG8NA7OUjgX7coCP8HYIcey8VPQBL9DyJu7BpDVq5AzLeaTGYzUPZ7gGxgdAak93ifXyemMlXmE
sOUa7kLPD9KqBROnojR2KIC2H9T5gbbX8hgF5EXIS6u6bx5bk8aYw+9SjXLWPj9yEJ/dntGTgCDH
IKtmv2HCRPRWRddOHffdPyaX+g0QvEaFFoi6BNM2nxoAsTrT98+4O4KQ9A0ertR8ew5ANTsyWXWN
GVbUqlPQ+EFVKQQSNp4lLLDhlwHdIihpWnbdYmmqEDDs6B7Nwwl4IEY+7TucjYqwJ7rWH/6jE63y
S51L8ypV6YHCN/N+S+96XFrWsDNU6rPbbL14+nDU8Sc+JME4pyLwNI99KLhiTAFtmiCrmsQKMylz
KCXsxZyXqgmmxsg389i6hsPdWMryRN52jyWElZ4eg3tM5u7+mUOuAbVf74+PH7Xqmrrph26a9scb
S8SbxOlgwfWCE7Ht1N7cBUm03H1aTK0wjyNlJHHpdK56FPBbET6nkesllKMgimj+0wXsgGsk/B0d
wxVcrdeE7T9oui+R0AuizcMJDfNTNcx4eNpou+xK/J6D/Dp+uMlJs9qvdQoqTZgdDcBiqaxgeagj
hPmxtcbx8AbVaPixTQmrkIRwzFOMPqwNz5Iwa7a2Vo3SWSBWYfbZXsYl3FAsWR8NVs2sLzTR8/zF
s4vo5s46PUcl4bbahhSsDDxUCdqLsfViC1eADlNqlqc2xefeKbugLVscV7WyZUJ5ar0Jefy1wcSF
Hd/pfrFG/YBBz6mw/7cZIX629z/U3vc6jjSmUgOZXl2NnUoKUuWtdmL+X0/4p0iXWIv+XBg4dTsB
gL5Im/WqBwBHulAFL35GOASp/wS4IKzNImWdgqghOBB4ddbIZJaX4UVQZFVznKrnC4mL8eL8R7pm
UaWXw8nCPuPsQ/SU79SLWo6HOOk8uKt/dUOhqWyXPXo3aWSVJHVBG89urzK35A0eE+yBfHNWE3U4
qcUnEGMxu9QobBBb+bj/scRa+IyePj0lOV59+3w1Iog9JIWC7CxYflgVshIHxZ48MIH7CR4PThMe
WCSAjQH1Vn9W4UMWN6ljZUysk/NDKR4fcYWYiHLN4nsim5LaIkFhPDr7/sYsO8RRFOy/sCEB2avN
rLrOV27iHJ2pcooDy8GVqLOyTNzMozXcFXK/X8NSEijaJ4ZXTMFKl2yzx422NEBoy6RV414Y/SE7
VF/OWLe5/XG3Q6yUx9Rp9bN8CZ9yqv+H8yKbxr+mj+wHxAT5RmnqnFTVFyjILU+1rV61janHdNrA
2caFozsdDDVGhWvAn/tJfeTk3pqU0Kg9CR0O0MVTk+zei6rCrNFVSqRJyIqrFqxr8DcZJGMGBUEz
kibvWvqFR+ZxtMXqKbsQliX+XQ0EksrQM/m/tZr+glQ1lcXrOZn0Lm3JhH9wBMZHM9OBksLPNSr8
Vudo8KnrMDjxflchwSJCQK2WcA2+RseXnfG2/cY8mUYxTxGgpuGDhUi/lnMg0PMa5RXWqREluD5v
QG/aoFOXhdJCwUcp7bl3axcA/VQLTZQ+ZqSUkm3uSNjT60d7EepotOtGRPAKS+J6SslpXZULBzNm
AsErsTfYIElHXSwRJAvskUQCFdHLlHD0l8tr0Ma5OrfgnvuYPlwlOuZOLxs7e/4f6nltF64u8uA+
RMLWp4isChZ9mXMcqUPR+/XTI56Yj9HP2yu1erAhJQwzuWVIIN2OWaEFH63Pilg2kEVGxQ3bO5Cn
OAxmOvdZcCh1pZ2/o7S3JzQnDL8fYNuf3Vh59+MjFF88WHE3qHIuYRS0yvC6A2FP/Wr9y4HAo+DJ
HHx/hD3rnA1JUoMj6jJ65L80kcfLTA/5qTOpdvogOrgV04sPeDIft2NyohKeN9WIkeGHuGUinc+H
QsS7si2Md1brVjNCuaCjcLu7Pt2ekpqok9/FyZp5vB7mkQ6CMFsrosm6gZNNutQnMzrjZweP0UbT
MoO2TmhFHnW3InS/b0gRhDkLZsh/zKiRY+KrygNY7+10cCa0h4Gjku+cWSCACHfYfXVD+MsOLygL
Wx6VRFMz5vYsWM35QsiFeAygXgWMm0bDPdxT1MLitYLFZeDdAPnkhjVXRfKR5w5v1sNDGj32h9vi
Lr7uWiA/6bjPCgWuX8/WEMEqNh+c//DkNYCO/+I1vKqjIwJTjwVOIbSGNvhbFJVBWQKFRV0mvBzj
M37MX4jbov68MK7bQQ/8EfiQ+ClZ3pydTAgHYw0OZt8caQCyALgCM5SMoz3SyMiItWgH5fgghZF5
aaCCvK8B+toYwMvAEViXKolWvpezbDVuoLD/WjwYA27oTcDBdoXdoEi3/dx7KuPEc+qZPe1TemiF
160vcbd/DDL59CpzIdfnzH29kBW45YlSE87EBv4eLFnSjSzuA2Wq3q6k9aoU716uJ1UR4rEur143
UZKlPPir8VgRUGnY0K06wLxoiGFhbIg5JurRLnWPghvqtxe6ihrgLgdz9kkQ38Y2c7e84WL5levM
BO87n30Ua3r3cupmw9j3Rd5rKNbLc9BT8BGalq0xUgnW5yNy8DcC0X8TU3L/+V7gHHaM9ee3uLdp
+LfcXJL5R8qb1zeuqaIsa7WHlo90EoaBQvDmeNjP4Ro/muuVA63q1JjiOKRndjixNDQkiTAIB09m
Jy/lcXIJDRR0z6YdLEIjC74EqmF9cXeirp/6j+YHc7DBJELDB62DcD82d2SSSXScKw4is3AcjyBY
cYA1CUDOco8AkKOk5itz+u04uyiBPFoDmiskoz+SJLfREBAM+twvHy+mruAhIrZh0tPZyMUlzp4e
JsEq0US5CfV1tW7kdNs/I1Z35kl63SQJZHvN5y9svGRXH2RdlQBq91WS+M47FYmyWyny5y+0tCDi
5Ma0mVOHeG7RTQjUbpWJpA7WoJ5+UOrbr1JMyBtSF8WisJfCS5ptleu4TMTKnYZ78JGFBB6eO4y8
Gb86x5FiOK9i5oN2m5dn5DhhVYE3msMJyD+pkyKrDyzsdKjVMMQRaRR+eT2CX2jd11v6O9k4r+8E
xmA3AuGyU0N3QttML9q6MUCf0KzDm0tA1dqSRirbVV1z77nhrk0sMc8kWikc9aZWAWycX/DVaucA
x25hFD+/MJIzIUJWCZNkVSdq57QwLm6/ZuFdqk2tBzLCkoVouTQAB9UsZHxGe/3YurIU/WkL/WUm
nbovQ31pB6FZok3D33PWi96Or2OqD5uMBCgj/ZoQJk/QiKSwk/zlRWZXaaaliRgvQZDWn43QuS3D
2icDuEhxXtYw4G6E5s7H1KqF4gm8fQ1Z7Lu8mKot9IM9yOQB01yiKd6diBR2wCxbRJu2+b3u9CPB
0vZc+34iGgkEVFeuzZSM3JqkDjOqNBgRF4YHywcCrIXTd4t9ajVFbSzWelncNF77e5J4o1BCRHXW
GBsAOlZH8IxBpTzUZJSmBh5tNq6ISai1JZweHrMa3sMYSsX+eFuR7m5mo3zBaOlmpsxVfHwy1C0D
N+YgemUYTEHA5f3HtJEqm7EBKPlRGSj2t5oPviNTLy6lWMWt/yHlAwXZ9rlTSSCrbtCXlwbsouJz
E5rTEn7mQ0TIe/eolY8wda041JaEVqJAYguZT50LYAiXKkJc4Lk2+gfrGG+dJ7w8WjvyO8LHZX70
y0Naa6jzbDY9GiVnaYNOkwiSq0PoZX7U9F/7w02enjInhAM3O0jNCOMkqJgPubARNW8jGKj/Gseu
VZ77rGFuSSyplc3rqiz2wyZqhHxsCoRHf0LdoXgF1DK2VAtmYu1jtJGxlZUy/f6lqe2he6OawWjh
96vYA18EuZpHLSVkoefqKxeFxL6CClO5pdyLikecR2TmzyUs13mwHRrFEST3Msi26UxGBLBW2JsQ
PF9YpfOV33LzPsc1psIC50zdwSD5ZxA9yF9zoCjSLIrVbU6eZHc+Jtd/v6vAMmvA3dM7ISL6gY/W
sNMw4BA4H5/VPV4Hx6XQFLFaZvLuR22X9EXOi+JxbnAWG2D+E5p/C8wB6vgQFMH4/VSA170qA0sF
Yy3jNHzeNoLjVqB1hM5kRCmdO4knYah0rxyc6swK+4jbsHPGyUze0GraqG82lcQCO1z7q/+qMtBV
/4fCvXPv3KhNXQGlsTS1a+oQr0Xd3VoCJmrOvBGj+BMpVNWN6qTDOM/uVTpUuseC2uhpMx2PidMl
1tnSrEc4KOq6kN2I21p+IWVZUiYPnu9NZDMbURuJ8yfbifMbJnt/CURFCIHvGrFMEosrFL6mNfqU
pqfVYJIc/lY3s453xDhJfKt2gmHrDi1ml3TVw9qYFzpmZK3R5zbHug1bZJUECp3+GkN/p/Kif3uY
XeuDuM8ZigGbmACVtsfw01kHRUXGU99QXSYjlCyhjoowYur40A+5YpuZKryAd7M3HIIxCdfu18Ws
84OGjtS55vUmu7GzCKSaW7xCMBEEjQUM3Lvy6/nW/QroGpWiu6Vl3zXt+qfTWs/LovNv3fTsSl33
icERVK7Az/RAgQ0o0SB41YPKKEsuWzXsxxe4OGSqyslwevRrRNe1A6jcJHqJ1fVg6aIpWGkvfQhV
sqSYJgbmXDm41gDeRM65xidPusUl7t1+I6VZ6Znuo0TMwqte8GFpsAlaVmhKT72STyMY3o0kf3np
+mL7P5vmlGQKFDTB5YG93NCDTJbhXclC+jmI4i3P+kbK+QTysTW6HYJ/ew63Qc3Jsh1DvcY3+HuY
/aPsjxMsXNswj51sAkjI9ThotenXVbq5OGU9plRJARJpBu9YU6sd9wJ7RAdPLeUwRWjiMvssjfQk
Ym1u48xROODU1QQbfkbE7x43pdx73pCTOctfxtmgMUntJtfkFg0V3+9ZPu82eJPEQ32WhEoI9AWK
Jn+PM1EyShU7zhIfl+TTKzHagDNHXts6nHX3//vhtcE6E2F/DVKq+brv/VGRb0uG8Zqhl/toLW+a
ue4HnD8dnhtRv5v+WAlmykldjorROZeYUdlmtrdn+l9J0zL5/2D2C9nKTeZjTyo11n5MSGpfGsz7
Hsi3b1WTV/5MdcpBAca/Lp27bDxFlYbvvlK5Gr1DQKRmHK91YrtQmtx1R9jozVpDdxCVuiyXBWiq
0/6m52iBMW57hL03Y2KQhKeFwongJQgrDw4ARaFNbkFJHICptPsGEiDWowW+fhjjVKdXNg3sPn4c
Rbdz50KhnUkl2edUptf2sSE0TdqRkSos1NaAsLtIMXqDaPUyjjKn1i/avRCu7KNE9UD94wnSq2TA
IgZCO/5zIye3HjjD9LQrY6bNE8T0vv7zNoXde9z0pGpBfRwjHg4dmlIh1bVsVXjdqGANCGzkwTfI
KZtsCotTtJQ/ZrH5CCvhp7WGYcWwXdFLKhOb07u0tQf38yoHBcaDrk+cpnsu+sjCdTs9TwqDhoLm
IYZrIwe9tlg8lPoyipQtMiycN2iWW3U+37OSpSWez4Fi4dWt4HFjnDgXz9VVFyylyOTP5NEfmfiu
sDjktceZEYSgCp/66Slc8U8XYz93Ie13jEDVc0W+coGlgDvwvM7nu9d0cEf0LTsmQB+RPCJXlip1
pCDqJlLoIy65sHqeToaqTyyTy1djrtAksQDvrQq3kmFaHUppwQECWD4LNzQMyWcRfyyIJHbGRRXm
Oz7Bbj7B81jkEqm/bMYZaB9oseZIav3V5rVf8/COlXKqgIawFpiIp0nljtjFmDuzLRIHII+tvaLs
l6skNuLwidrNxLMq/elcFzf480gBksFdOOJRGZkWB0zp8AmUKsRf6n+OIOHY6T/8pfiEEjyVEWHB
1ZocyFokiY/qPqogRfS4bBvQcO9e/cHVTIsQInpGj+R3X+sr9zb4x658qMFQXTw5xeQYA7anNoat
REKksaHsKQtlL9Re3uCArVbLuOAopYn7hFvMesFUbpoLnL/zGfAfEaci9TIqSIdDS/P5X3zjN3bE
jSO22x7qvGJ5XgN0yVUgRDxbdgcTDlQfDmoHQf4zimCIUYFXIdlSQmEWaocHtf+vBUSSaa594Udv
QN0NPqfiG8BfJ+ocgkLHsK/W2zsBcYahAUqVMX3P6EI0Ln5ko48CR8lxzfJu1wLPibetwVvwqQBa
spqpyO1G2MJxolodVbtWV3Ah8CPbIfHY9HnQ7l++TaQq5W7V5VPPQbYZZE2x6xlGI/TSVMKw7ZWM
dtSTnp1r1j1Iap1CfehjQDdfmecXx6PR53HB7gLlWyDF1ghq1SN/+MYaPTsUbif+4JlofWJCPX5O
ZBke/NdPvwni7pZtnOiwdvRKkLEyWWUMq2Nl0UL8JBVrbXRgmbQTZHZCEjUptAIOOUyUdlwMvgiq
PqXtsvd1ZCi72bdMUNgK3EosJuzCVuFGRsGsG6qaVGqKCBkwkLyrn3EwYKSQKq/lx5TYuO9C3Hlq
ZC8X67BP8mTbRLlwkKLbslYB4tzQ59TZG2vsYh0jVC6sCpgHyukAVxKO11aqgTNBA19yHjR9LcTX
KsHT986P2E4pOPq6gn5y/8fsIWc37lM3cUNjFt1kbv4hGcH6kizN4w5gTLrmSGRmbnY2c23yo7u7
P9dlM7awz4Z0A8CAVxvPEaN4OxAb74CxErFxPa9j31kZc//o2oZUFd3R48SLHbFD48f/bS4J35ub
wId3z2ZAyrsb5/KDNge9F47yoSfK5/GXbk2IqiQkA/no7WS6XtRxVVZeQNmTDjg2tIUV5zty8T9M
W2fsDmn7PiA4uF9CRc24Tcg8eKSpC+lu66lBpuAIWUTbzNyFC4Mkr7J1aASlmU3bA2DDd6kDzjHz
UGHnFFNFF9P4c+tFvALfRRkm5oSDihTsFtQqnBgO3TV2vQEucy6aya+vBWWZFc1Lxnfq0uIHfclS
rTUs7KuHHHcLllt7VdfdOPuCteWUsYephUSUsG9Os/DYT8BdW/ccnkOeo7EO7SslVq4jg+KWcz5M
tGPDYQxqBjxr2JtFUlQ2faSDS+JkQnBdYfdf8+VJRUZivEvGXdCc2Ljv0bB6urx7b8004WOBe+Od
FGgDQCfxISWdBTUEJO1KJvXVV5W9PVESx8EpdnvHRI+7r6UYh3Od9dv+gsFTGulRSeXYh6WOp5jK
0xrjPZZ2fFC/4gsSDwFQrEToC8E1g2rZbyUfLwr84GY9omwjtt5SaQ2uglhb3czgXzk3WhuqJvuu
9LpzRIG41VmqLd/yIJHRDxWtBTYvPvvDAZ42UwQymBTJC802mm6QVlWhk6XWi1amAp2aEAvIAHfy
D0AQSPLvwMg2X5UnRirUMXgeJ7Inadpvp0oFZbFZYWI+9J+B/GwGCANBy3sWMmbem8qxC+YaXvrM
hV5OpwxXNjPcD2AHP9X/lsrbjgCO6a/SFcr+wjMe+5kTtQxayAsPMEmCcS/EvBlDe3oQ9bj8B+N5
+SRR9Xd4LhvpUNVjLfstzB9o8KddYpkdct1yWba4HlmSyf/OYX9HMDNb5kYqjeb31ja3lmplp+XN
Ld2tYPT/dAYzh5kBH6X3E3565k3gWuho/QxKuHag8ykHWgJItEwqUjtVzdtfdiKOqj0ywAw9jwZD
9rCzEpQ6hK9wcG7/B6GlEjTWz2x0RI4mgXIylzpnwyU9SsZMVT2RoMoD5fwwquOUJkx7dzoZyMA3
dS1/ALn+FKnrfx70P8fVLbV6xmFnZ21tOT5zOLgN5LhQVWUnbiXw6qp+LXvb7jdnw/F115pkhuvb
HtEaAedd73iJNHoU2NDIZN7sINrdduAOhDo5Lqwwd1I5tqrSiE2CJJBKUgxvyZN3EqZnNtMQeSuW
uL8RnsTEj5CAJ2wkZJinea8bMlN4PDYA1o11s35RNDg/Jnlygf+Lz4wq77eE/ntvi0xrOh8t72iM
36oVXWjrk+kct6B/lUhetO3ToRGl9CZlGRlCqzbVzFX8vwQJKIaWm7OEXEd/jTGjbB0zRvezL+dK
2bxwZAHtjJ1rsLC5FaZRjIc7SOLNAVgrY9/XsyAAoYtIflsgV9OwPymdV8dFMDc/QCotJLTnEKZ2
zl/Jv3gO1NBNa+eiqoY+Lrf1R8R2xmKD8KPTINyHrUFYR+eH1AuCqtBN/x7H+laVEKz/kzM6vDig
ajPEOTQkcSCeeVIVsMEKjkCG1p4Jjboq3G5fKENbPRauAT8YYCbWNKdFvccQEXsqXK5r/LbCXe9L
vRzTSi2njkc9R5Rmwd9R9Vjg+SiknVf+yWs+YPMVq0y2ih2lQpi7ZAXgXtF/LluOCK9kKzmEJmop
S3sMaXzxd2z17lyejezYXueQK8sXYfPUwYaKpUuEX5Lqc1xY1Hz4BiC4HX6HFn6ec+FOX8rMtmup
cK1QYHa8HEDdkSNsjqkMZdX/QpdV+nai3Bj0LGdxZXCLjoLuZNYT/Reu4BMrAUOj15uspLN3UzHm
LItMXm/VkxEfjgPJiuB7Tdygpx18nM+k7DkIOnWi8Oc3z8J/xiAqxcG11O5Pwja/oQUu9hNTv3xh
iWggM/wXC0dOYymGATRnkBvRMdggcgrdzm/9hyZBF61Q1lEEAfPPCZcqAt9TSfu9iIEJ72yy+Rsd
8xAY4Wjc931ESUQPXHxIL78huVLWRmT6S5nEtQh+vR9Q0HQbFPPhA69r694zykPILYxJmzq8fI/l
jR/lyiAj2vrPbmVyT9OEcxxVIzZpeOnq9+EOQRZCkr4GWh62YtWAWyyIcQb5DIe2FgbwI5WZPryE
1QJoevWLetbh41y/piPAOXFs4ILvny85UuJG+WU7YXD8wG1yBLO6zXOvRNYZj84DgkFkiiWqhRrj
Iq3hIe+uPgpKeeogyE9iZFIbYukX4rUSsIfOpafRvRJ3Kk5ym+s/sGjjHJe4sDeRrE5zusWGQ6ph
NYDjVS6Sk9P2nMF+2FRMI2r/dedODtCt8aJYNzIXKRYM6mfYX9RGLMDUhDRwZ3vE8qT298wJdOXd
YgGlPhURR3jCsDK6XFRV6xizOc4K7UHzbc8rxUc0yUP73qfVyQMdJmRVB6zX4RMbLDA3tqKXDm7X
Pc3C3oDzjqII4VG7+nU1EonX4V15bZK2dettniPlEnGDF7666fGeec2zhUhiTkweY7+MDO32WZnN
DkjzntAdW7gg6ssFT+goCKSW+IkNm1xR+jrNnuGMhL7pAQboGWLfiMF/w+0SIOTLSJeM30NUMfoi
xHwueE+k7C9XLYymlpjqYYL6GJlmyCJHZkVzJcriZ9AWfu9hU8K3HzkGRxJTs2Hho9+eogaDkG53
CUBwbtvBSblndKZFyw8pqjT1SQgeDW17uHSHudrYA1tXCAKEdRwbl+j7sEb5Z+f9onaw7N4Jfks8
CFuvxmmYczwPfdm9ytR2Ya7jigkWqCBQN100u+vxGWBaL/BN6rbDzs9xoEURW+MyFApDpdkTnS7+
e21pq8J5x3pHLTIqgFOLnIvAWT73veWO0u+IO47r9P0ex7wSyS3uiiOcdU0SDoZXhQ4M4pNKwEav
s721GTySbeRgDd2dq/TgRQsWbfI35RwmDaCMJfG0CucrCSlXkdJWLET1mhYY4qQGUF0AAwtnwO7e
ZretmNDR2UU8u8vnsys8qLhviFhhjZMvHuIJuuNElN+x7HBu7yS38Avovw+SDHQBnwCM7Mqrke52
SGEFwjsZJWZgm/7495R4oNqg0vE8lzw0isDlRpv388rRW7cNs/1xwCnCKJwKf3dDKi/dJYDXVXOd
hqFAbgxn1YFoaMoqkLLz+W9ipxb74WVjj52Z6U81ugesP/mVzxBpi9tXh6kCTGNtZj8TVSrUGjJr
WPjOiP72PnLEFxsz+3Ylsgmnm7oC2u9VsaeSXi90fAPta+3sO4xbpvdmoqaZfKmzpR7gy7VQayR3
Tf8fIRMCPKmlMLNIdJce9NHSTCjF9pvzMhIqJNztAcJPjzlUR6kxkn/qNdnDWhbfHdvlhkgg1p9F
cxigatIP60fzLG98RN5nvQy7PoWm4r/pHOETHh2WuTSMyUBw3l2oGYr9I59YyrngNn+BiPQsYF/2
yEp9oYZ8+5GX04r+eeWyV91Sy/z3Yj7rUpPTAm8peEejW5qOnFhU/GMKbYWIyi4esU1UGPmWRn25
Go+Qu2UmrOX9tVSfMOLEEKHqW6BnsFNBV+Buu2gvR98GEdTEBHYztGzG+KLUCKYHDPEyxe65UZ7T
T69QN6e+dw2oremqTtKLXHmoCMn5oajD004ilXdXZYgsfr2eMyxYhW4sBuRPcVmxYj5xmbuv5zQ3
Igs+KxNK8+XrHGKF4+snm0DW175XpZgqQxIx7TPj+imowT0JUVrRO05Zi66zPosnR+JvVcxC4NeY
LcowRNAdlmVa9/eOhFsVc18TS1FXWm3Q8JHBwbYRda6Ah/qnkv8Iw5D8cWaOXaOHZK2VTipfbrDQ
+VmVVqXpofcStdZHhypOi44d5pV4Dw4/VXA1rupphzt58I601R0uc7aL21a9lV1SpeJVXx0CGgTi
gPHyYReFZt8dHjN+7GChm4AlI983QYj36N/mJyJWMfx+3gl7nplBJ3vBaMVov82IMpLRVTH2p7DP
T7iN3rvUZcp3I90+ODv2/l8myCj6YeDj7XnJCFZWHCuSdEUstf+UBpm2Z8uPrNq9PetzGImTMlNW
IQezJnyiXzY8BI2yMSq1wDYSYU8FB5bFW3xTSpfsoS8+sihJzOs8b2kS+87Gh2n6bU7K75dcBSkc
7jYgAlhEUbmgjoMD+vQXeidUhLg+iOKsdtVK84EdoO/C1BCzG3aKOkG5oY5sx9Lxd9hIPal9dKOY
/l9yYW9ZM/4eeDlFemsdWHMsTLrb9G6WMHvT7AMbQ/xO7+dB4s969v0n29t23cTXU3uHhkKQICRH
Se3+nVOoZ181yFx4FJyG/uLkEQiu3ZpYqn9MlJyxv7yyOtwX+KBtGY8LEZ3mJZ1RsRas7mSjHwW0
/1uu1ScMTzYQxTtuRTuu6XHSPlCW11FFjNwI7SGt5zD+GNMBqWWtGACfYAPc5IXbUIyN5NC6cy1N
au1soqKIJ0YpMN4yp4wDZvo3z9rLKz1SQeoohbP93OqObtXYCSUMF21cL84IUsA2ZFMxLDJK0Jyd
SMOr1T8HzSySrwP/zuajE+RCJATqoOG7ltbpR9cfAEc6wtUBTOtZZruOFSd5dbMqiUh/ysfBTH9Q
7r3oLqbduS5V9SsMNp2pKgN/vqFBqAjVql6NdGQeXhUthPIhvKTLA/vf8PbTymAFJixEypWCmTj7
jji/+jl7HoObt18Ee9CS8He3eBZcnsL6kbnSLG/IDdJ1IIiwHFo4xi/+WkT027RuoSH/4lYWoQax
bTc0DIqnsgrI2SheE7ow3+bNqp9ygaxEqgtCcWtXeh5JhgurZJ7/HeXdI6vNIXYlepCNzGMt4yfg
7kIxVt10u/4qLNif+gAwtvAPanUTIliPsC9/5L7UV01mITNExJsZ78dZ2ngscXK1nwIpM21/Z2XU
5DdKvXr1nsPDwYh+6Dgip4aV4TAFEGzYRXAe2OutnoaDf+tbuebMvGkkhQRpnyrcgJSrRLX//YPX
w448r7cfBt4EZ0+AVyqfESn3kw7juvZmv/e7IsAmX9xpHHzQ52kStTNI+bxcpxX5oEG8l10N+SWD
XzyAJBMI3gjLxuPPq8mxHQVRrLOwxLi5zTAzFtjy8Wj6XuUfWqZf5oQ4qQzmt6wL8E7h9w23ZLWP
AOivb3ohOOG2Z7I+5xO8p9QF51MLgjMBlh0qNJSgeFhLTjz1Z2olF5T96SzpHwScJ32xiim41A4q
Azpuy4LcXnJK9qLgtlp9YlzkHZHXIHSTAweP81mCAYKOJSAsest2HDApfDRRkIgaWDJUq3LcJKIb
u8WHsXr3EaKtWg7wIeDeMZu5FQeR1Uog6sj5wZVReEBMSGf0G9dJAAFBMgq2CuLJxyJYBAf4rgNx
PSsttksikZ47POXWQ7p4a2NQPIqqMWBfLKi3Jfxsyak0snLAm6vDlrg6zvVAssgpKU439qJEfN1i
HRD6vks/8a4DjAiZe5ETQpfQ1JPRI1wl8GQLx1qtPoVBgDo6ofvqZmMTPSoNhcfq58w1TDKDMGeh
e9l7mMgIW65hIG8+Bsx1rT5AMuoP65WDAOsVuCWN/6Yu9Sf7NhV8TBZeHhl53UY7mB1yP8MJiI7F
bw8uI6wRlmP/jvOddp8wAZwZcr9onUjNqPMfF3dArmh6OXD2HHJFQMh4H+/Intk3VsfkXbTQ7Kri
6AuFPPwr3FKt2DOqCuAn34DPR6J0OSf8xBK8jqjE8joMqrp/VN8F3K9ZgiE6b4Lnkc5sHSim4U1l
U5SfdnDcWyDsyhaNo4OsMxeONYcW5KEoZyO8H7RRY5WZ93bB+Fz33hV+2f1D5BxhcEhtBqRom5o5
7R8LQ7MehMiJ1lDjg/p3m7HIZfT7Hbi6f4EDrVypgRyC6n7QXE0LGgzBRm7qJuPgNERZeTrJt3/1
BpRm2NEBBzdiUsI0KFc5+GxSG4EDnTqMoM404Zylp02mUSxhqU73SJPWKm1yQ8KRWUCHoqmdQKhH
z7WFobecoURgCCV698uw8BAZ6xIO15vyQ480LYrvZ8QvgBK1tcxl3cpgqQqAWDXpy75wHaQt5yUF
+Vam9yeK1xmTmeXyHILhXgKhBWU1hTow9lU9q5PG2ko3nzSRa0vc5bhvIj6VbVouwrTTLZTs8xNy
hNLUGgWxfDb0wIG/EKNldpSDIIzqftPQjyv8kUPdtVEPK8aU/FlcsLwnh6qkXjhIy73cOgxTYNGb
XG+XAd0jOBDuNi+v6JuWIGX2GEX8WkynGW94m0k3cnHSdJbvf+k1BUXkxGf4qdsOtdGG3xhbwDJ7
IxDoAzoISZ6WAts3iz51JJfvuy1DGkp1hvcTEByIPO8RxGRFyYC01HfALy+FaZo86KH5d+dehT2j
/akaGLl32gDVLzkA5a8LCGD2rDjcWSdBwEF6g+bW4nG1TAp2d9ZSTsMLTUN4wynCccUJUf+BXdNv
c0RhWv5pO7AUkNlYbCofwZUhD0zpGTwqn/bXCDq0LICPgxUPXZBeaUPvyigxcCxU92s+qxFGBUS1
9LNtve+wWfcSnMITdkeDKRzzeBuYUJR00OU8Sm0rUyOrxvnxHgGD2To70He/0ftzbfwEzUNiCd9c
AcWQJsIKHjkjOUvODSQiBE6s4Rr1q2WTbjYz0heV0Uxm4YOFHY6dPM/dUVWzgXIBkGJcML4NXnw+
26orSWja4bOdseNVVnie1Jfon6ZJr/9TQIclpUpnfEiH7IIslNq8EwLfA5cCIKfY9vh3G/b92T1u
x/+YmYVuMNeXThuMH6JCwxZOc8HtBHD29rDsRnfBX2tHj5vujwMVlx7G2zHdDJrOZboNOxxBUejG
X4yuP6siQ11fm/PKl16HGZ/5qpXWDjIeouWTHKWyxryfJ1smA2iiwPvHNzqvW2F/ax3eA4wVJQ8d
emEqJqXnZaHC2XwCzij7Y/nzNvZ6WveA/BwbDe5S97J+uqO8n6fhmXf2GLbplJRxVPjVLNRSQikB
a13BKQoa01kQtHo/byIZfWUM++Z54ecqdcrw123SEEm0CA7Amw345MFrrPxbry/6Y5Cd/HSuAcSn
2l49a6i1XfE/KmZS8A+7zvk3AalNckEuQEIMrYkH5caRlAHNrV8RjEhNpV7ufnvs7dnStxb4y4lG
j1unKA9LZuLGe9oqXUzvLJtZ3JgRTpEVUFhXBtJFuDEs1pZC8aUmC+PzftvjaS5T3lcvHLDeR9qV
7EMT5NMlLZ/fJLe5wuL2DH3/S5Fij65UGSgEv9ZzMm9d/8afPkdPsW8iZHF2H/mmFrMQrAYB9QIF
I/f63u+pf1G/hp6BZysQf5O+xSficUKQTrXd38t74KJ3zR0zyVdNkaBtIZlDUUHc0IifoKxZw3Er
KtzsoKNDxiU4VSDZQwJMdE7tfHk7YvEe8ny9dBKbqCW5EoqJLLbQRnw/1Nlrvbo2Elv5NoU/2xKl
QYL306gVRKC2lv4OKx5+NluOk4/NOoVwr1Icqpa55NEM+f6XjCNhcnSDQGZIk7o9tsMaK2LLYNmT
wzeNIvO4AbfuHVcxYwfU5gfLLFM5CSSuHejjXNwyCgBe/sELTM4hUyIF/3jRy1la1MwWBG+DiMu8
Tyd18LU4XssyZNsDQLgPDazN7mdBPipUOFIr0/scEg5wJ0VNv/rsmmyOlvFWy6ohtDmHUUTBvJa1
IFLtHdzyfgrSyTKKFV4TSuzTe6qUJHHVgNM012fDA4nBERWSsP8Chk9ElwQ8HZob+jGOmFG8SWGt
4W9qKX6D2pwpIYwoT2+Cj8YWFCmHae+SDN1a+Z8GWNDOgsbQ6Tos2IXA0Jc/wdDCbENJaSCy1L1/
cOGyH8VGlTor80Nv81ZignvrxKMfU9COsmowP08EjydEox0+1i77+u5NFD/lMZg6k0F+evS+ZJ5b
5I6rrd34Uz74/RCn6ucVfW2w8hUTE0/sZXLUUptR1xXX7ws7LjWpppu/jp5g+rv3MMpyeKdlXi7f
36lAWflAqoocJ7vak2jTbfT1yspniLg02fV99f9AiBwjnJqATG2/j7w/ibyty8TLQaRHfMVKUzB7
85+Z6KmOMywCbkQgm4Pfd9Od6cmCRUID0oC54XOFPogqCGoWdlPT3uMxgr6Vt30LD2NTaf23XWi5
UXk6dATwTrsvDUqHBpb1qBuB/FYcYhHac9pSnUz+zMx+QDgImx8yMc8KeWIBZjVqVZXxfrLqG17O
XS074iBqvd8hL009zesU5/2bVUTIuF9smhZyTo04xnhLrBi5Y2ZMMHGH7We7/oDoEA6V6MPGFVFT
jCArBaU4rnriMGfiDrvZiniUtuzEqXZujqiM6PIcmK0q/E2WcXQ3KQHCECCUCBtdc8nWzfgQY2xf
/h36ltaWiJ5nQNfOezzhlwPl7aOeOIeVUm70Z8JQe5xTIpiw0CPVhHipQ4O5Em8Khhf/vDWpQB5l
9Rj//91EQNp2Bi+8AuENqvp1gLoejCe46ytTNhnOGeV0catOVVfHB/BwHytle1Wcr3b2Z0XAMtjk
/Gklb6OFsyXtIT1HBh32nQ3RjCv0WfPtxH00n4w9vgEgCrbrJlV9vCGQuFjmv1utblbxBLMeJqfU
AMF1DY4uwtS3pspqPIyht8t+YX9wmjx72WgdYV0klMVev09HOtOjEGj4IYJHHHILn+NKrXa3JqPn
RIVBLgA1YFJNdyJemK5IysuUnkbefREj+60hBXBIih+sw8P1EWziaFDlJw1EQcKURDY2fAwENKi0
2lJ8C+RcS/+yCC91UbOnTmlunO3TYFUHoXm9Xd3XrbS5HjAEATte4XiAbk5oas+1Qgc0r2TQV2Is
/ID7voWkf08EKBZZOZb9vlI1Wk8210myHJ4c7Gjxrh+ZBAz4shG3WSK+Rh3ZVPnyLFv4bwtvfHol
6IpsAE8YSApA8k5E/ieTN43ZQ5ggs1NG6BVN6Vx80scyZ5efqhsOMpvIHay8Ca7q74kA8GKNxKdl
9YbFh8FbtiPpU1SDf/QeuWOF3wQjMKB898OmgvwsfgCx0q7/mDgYKrZuO7mxwzHytX+tzvFaVHXG
Xyj0cXVhHfrFlI+KRvc1zTaNH+4WY3Nxln209QRJVhOZa9nzPTgzcZE+95YxR069m08t+WlwuxNf
duiZGMzZA2OE4jwpn61UM++LGLzeOGIckdU+IWWrUflACRAQ+UJ0336pKYrc0rKlMWjArSNWQDPs
iT1M7bj48ghNKRNxJSWKKrfL7rBMkQDg7x6yU2Ho+j5VEWdn2m+U/KBMmn+f98qScPvGBs6OG8Mt
NsrjS3YpEdtGRdfshv7CcT6XkEs2l0C+6f2tISyBwxAlMGrjT5bBZ/yHK6Ng33Jxz5uCMzApt6IA
YVhsnKh9NVn3szCN1aK7dhI4OfLARihnlD3wwhuMerU0P/b0dOlTgQiIv1jXaazUkJRjH3g/5GPo
Xk+bOxkozqtBUC4QYv7dbAD33XFcT4pupeu18h0twesqVZglXAOVqehorTB5K9kHLEi348/TdJbv
laL8OIRjGgwUdOk6GEceChbGroFJDQ0FI/QSxX1vb5k29AgddXC+Ivd7AmNRx80UmxQruZTXQdtu
tV+7QF47H50yMNvSck9qUpRXQK7KeexTqtfPcyyXfmmoXQCxi8XM3WhcL6PKEHeQkwNqcBHOB6Bc
q7UIgEkO9U6CiJwJhZO8qf0GYM8Na8bkMk7fvmDcoI9CZXyvdU5q3cT+K7dRtDiDoShM29ZcJ9Ci
+IoOQpuYrlHYZsI89ZD2VwJt7cOFxt5Zg+jGc06AA5VrzBFMtoktCIvjxXa2gCNbcJKG2SKrXTyH
TsYCtDwXxOZdH3tI8GBBAQcQEfGiJ+fYHhuGaQU1A042EWkwenX7BzWZ7Qrg1dpynUvhjJPhbP72
EUM27y2565IOi2PvnkE6wYIRYMzVRan3AOUAO1R0ucz2OLmGxEIqREoAIHqK/hWL4CpVP3xqfd/M
HmVB08G4BOVN2eBBGnAyCnVZPg38fanHym4ffGru00i5mqbTCOFP2XBSSufj1flPPriX/YnDWPIF
ANfiM9x1W4oVtVkMX2lDbMPGRQWJVEcdOHxNuDIJxpqAJ+61Nuwvz6WVSRxJuMWWzoqovRZ9xLc0
cyz1frS3cSTXINQKaOZCM5SlUvK8XlyEIAJyTmwIrwvxMDaeWmzOPdM335XOK+xeDZ+izAjLREf+
iw2aU6X6sTryQ6Nt7RW4p9HIuc6Qa3BbF2h6qPSZQKRi5zX03djRC85wIbqiJR3ACgs6HJE81ifV
Z4yZRVRQSmKmcjpYmwKmIgYUEG9Q+iaFQKYMgoTdkqksaVqMVqTGg1uRsstZ2IwoENXo3EZUlmtq
7MXzPDH7XqBe0gonYDHZ0tnsnc4/q1jWI8lTZB9ybvnx8Rej/MQbwgZBuzIJ6EXMMBG+ox+jLbH1
oLvWkRDqFuMFlJ6oFTcH7SwPj71du3r5KRsQH0FhHJFyLx3Y0hA8VewwnaLqk36oGyl+h4k5kfun
IO7CPA4gn+HJkWVtKr7frsmP6yt+rebTgypsBNl08ZFQhTCOuCk8hdS1B4J9zTuZzuDTZ9+Sl2/V
7z63mrF5+cbmnJWPMwbCpVwzH4/VFxQhGImJpRJKzXtkuDDuNRIbtlO//nj6SM/n4S2yVpglar/n
j/GaBZU75MF2cxupjH4gMu+1hLh8PjFDyzgxSvsQgymtocq48NPhA9bYahu1faSs1A2huFpp/cpt
ZClbe1J7/RpGczDHbK25f3DX4s05571tQAxVCAzbobRBbECBGSNlosQs7oCZn1uvmiC4PvPxqhEy
umGv4blmCVRTW11mD/IfuQtPpJluvApC5gfn4PortZ/yGDJplBY9SIMvr6/wdL6ruLhZhmqy5/hJ
v40ilAoV5bMH+tpVHchzXEw1G9BUia2eBxHDqOT3tFwpNHFjnNQfIpj1gcCG1GKV6NDxqeo91tPs
1wP3QNR74skayvGv4uhhvN5ZL8//1QkvG6WWJMvkGl7nWr0t7Rf4N9g4zQ9XhnC2pk0qr5b89tLe
OzjPh21p8kjMinYpcOCKNWimYQY20Qxlnkrt/+dVxQ/s+8P+aMX3Q60LsRIRk/JMYWq/eEz67H3j
goiK6M8ESfsKO2DAarHFu9VkyoFqo7hLhBKAVYsIeE4wzTrz74uVbNgDl+7P/nDqQ1gYrJFGOAiT
mHmAynUSHOuof7mWochEXx4duxAfqjw7ac5Q1xZCGBGwwVYYxABkH4ruqzVymDmf3S3U5/UoZUWu
xH62Pkout3vKL1d6LOUNaZ2ibzRT6RKiJ608PwVFS5Rc4CwaH5Q8TflF4dEr+HN0tuhtvFEIWtC4
pWEMu8AyfZ4t5dsUVI0TOdUaReDr3e8wV8AE1/YBznl+brzz90kiah97pr8eAL5ufwThzHxNiov6
bdbMSVoG1Aam9YA/QbDLiHuVkdorvVLHI0APwEpB+xR0vwykjEXAEw+pXT5lWSPv8EXff/42rl3H
5upfSNVW228oiHCb+KkzWsdqlTDNh43RfjqpNk7W6aw5B/oGvfvF/GDz3RH25B47T5wkjoCZhr0G
4dIjVu6UVFAWmg2X0k5lS8sfrKrV74cK+KfkQxj+dsD94GJDI4GRjYrmBWv390CW35dDGt3EZ1NL
7yHWjiHbz36V3vNCWhSUnpQMN/OJPel9NFUqNKI64R3LJk8q5OERGv9PKnmi5taFwdD/CHPvQZ3U
8l+mnMnktC+ZY27nLcVa3J+PYKztPWzJIPC6nSs7ksBrgWmwiwvIe0gsXzoS6G47+UK97Neqvytk
z5JpELOdX2nzv+B4n2WX8+BzH6mMImmW7Ral7XUq4BdPmRx87sRJO/QTZWWf67tOCK/HREghEAyP
UrXho+1w6xGavsLQBFSYN8IQ7VRuNwJcqIoWqS4x6lK1SxWgvhqxWV8o1tMnHFHtZHl6ZOcOYmms
rMVNLLNroB+x0v+LlsnhLmJFW2YvfMlQwr6Nb5FXW/zuoxuipMTr5I1WfU51JiUK3JpViAyIe/rR
8DVHEqHvwndB2ToJYJQODa+i24JkihA27DH1LJmveFT1ZUWZjXtfGiiV2/TiNLv67hzsk5iUyEXy
zHfYxgn1KXWw7U/hBzVqJRXvHvF6bjwj23GQ3VSjdqHGENlObxm0crTPzfTIediOvlzYRDv/2X2a
fOnrCR9vG12cZRLCAtG07nn0RFxXXauUcld8Smpx0yys3EJvZsZh5poD1tQO3DuykP9Sp7pzKwSg
46J2IwovaB+eeEPgEV5kuXfdaOWZ97OFpSvblARZyUj0/OOdandcuLJIteNvj2eAf6QPksHS3C/r
hVMIUG1IfyZgRkUPpk9TY4N6VryyP02jemMRJKWnhwKyXgAAVXAA6ZWaYiVHmmD5tHgweReCocCN
1jW5g2sbHyqgQKvpeg/kadi9TpeW087IlbAIfwypYNSKPFvzOeDvuRHT08OSVdcUmxfdubKscFA6
s5vJm8Im5FIEN33cCfG+eM0vosCYChZQnL35Heeh4VvQlrZfymS8QrPtJvhaqiKSwBKpgf0s08xs
ryZd5bQ3qM/pGAQQGrM/S2+UKiOvm2XhJrPmt522z5Um8lfs1a3ZPidXHWM1hBKjX8FSpwUDy1sx
Yx0VRVR3qUrhmS+3Q6VWwTbHMGVlPo3zIBqjFSHrlci/yL+axTTDOPQGp50A3OBbKFgzsUH3uP8O
8Rmv3ySRJA7Q7tP065wTW9LplgMCn8/s8bfm+TSMcDuha+ryG1ywlvGisXgtkDNgn1cpxwYnV0sj
W2iZIMaoB8UcwVPbJgVpyhoQGPL11YlX2AhSepmqevkdkFcKpNVAQ3hE2tyo9OrF2nxRC/843ckX
rwjmLZoEePIr713bfopEMvAMRSTp/t7PUAYo2o3p/6GumTZMPbskl29SfANrwuL2KpqqyfWsDmJX
hL7bU13wMsGHJZ8oNYoc+u1PLIdaVQ25F88z3lgdOirmBeZTN7KGRiLSihMyccnNzyhftIC9T4fv
qTteQJo2HCQyk6J/V2eCQaijCYxtZ5sFtNxjUzbsa/J2BMd8YRwavpLu3W/hLq/NFUcvwDgXp5YN
zwYttZXjeVw98jJAOVpnO++AE0uFPNG83Z8ejhjGya6htBQr8Gv7I/+Xqi/xDZ3NYV7ssfhRwAHA
zWusvRR1YScNA9FmtdL4tPFS3nEl4g1+SV0CUkvNwtF+/X9WTM0NVfcNj/qOdodu9mj74gwSCO5s
6xqT51y6FT7qw9XwE5CZa3H1K8wtCcZxKwPcO1bCV61fzz/njWPTGHZ3KdpbvXgowL0u0ucgzHRQ
SpF6ag9Z1NFaSUYQg5bO+pSyjKkKY8LbtNHUMmpHy35uzGSQqWVMT+ofIsExORm1uBGpR5SRA1ZQ
i018j/e7CwGu3WMe475zaq6XThduaa4Zon7AHj5YTkARdS88NNMH3iTzD7BdpSRl+5c5/MTQgICQ
3AyXSJpNk1rnq7bDcWhwA5F11iX8byFlZkSYQbcRbOXwGJ1AanmW8pAsGxhELwyuJ+dVjF6zbCB3
2YuDpEuxg/aCyTz5YafpfROiJ+EBIBsM0CbIoXrHmKC1FFjgcUUUwzi2r1WthjOmMQm2kG3JI1YG
9FFKO1SrpTvPb//mfRDCr+HI9YA9uH63f0ljFEbi8Ju3wPNdRZSK/+4HaXKdAaGRD5JO3fESb7oU
Xpk4fYCsvbOks3jCaexWCeHfw14oBgGU009XD2F4e8idr271I5v6E9xLVTpt1xOie8ff8B2kvwfD
Dpf7XLEfvdIIc49lFc3DzLdRo7+tV8tRuC/vJFxQuOce3ESYV4rXLPbAmXeHjlwoTv/iZtev/1Wu
0vCj961YvdLrIJBO+tXAbEGzuv0g6dpEqWBxI9yV1nxBLecpFl+AaZrPPmKYD/oN8CkHRL2Dm4+W
STWBRFqzxmzDNpfvODgAn4B2XTOUnkwm00HBLNpzJpPQctKd0d2Mn0BaFLz6zgc8LAzCWWR43HBX
R4y/4yYtgZz3jz8pZsushHvkxtmdpFJIdEk3DBoMf3SSI3ro86xmBdKukLNzAmigUfpQScgzAf80
7G7RFjI7PS82TewjCuSqU2FcEstjjmRRlTevMvY+yAVZEEI27NgbRxI0d3KhzSoQAHPPdglr52hN
E7+1Dj/coO7/L8cqUZ63vzSJmRfnWtdKM6mW5Fm5+AMa2Tu9e4LVU6+RKmTdzlySZQc4UcIfW1Ps
pwhHz8Pd2xs6jG7UthnitIb8P89uXu4B/1+b5+iHY9YCqOU0VQ8jwferPlpNHIAeEnsPqA4vaL6V
EBgJhh76TOCJ7EjjPXw0GsTlXK8mUCId1TvMSmbcQGU68aDFXoXlCp9PxmiygaFGlbKxZQuz+697
zCSvBUDx6BBN0OtxUbztaWd3DZMq9FzjQaIfKe7N+05Rgk0xHqyf1XvwP/M+Ciuc1Jn4iuuz+HJj
aHFy9PQ+NiTMBr1Fgj9wAldJwg03onZhQhszBCAMnLk8qh8IH9wQTPGPOrGORLKJIQ568a+GQNUi
PNeM3gR9GyfcbUHYMgMNqhOrEzj+zvucKaYdORjptYvTJo+7m2es9gNs2vGU3obkk5u0Os6G8nm9
mdLghRn0t6YI+5n6UqfiuSZVBk3Ub9lKqkBHHm2LJxhdp+5CI6y9+AxabfmuL4/TFNs/0NpZ5VXy
mc36cqFD7ajmmU4CEaTeUotPcUdvUhJN7WK+6BbVyLwfhz875elzgDTOsiiK6UySE5VhH434JVvj
OO6QxnYRaLQ6hnFhBQS2RVkYTvvyRAD1nRoQJ3EXsqPlUDp2xi6LIGuMnOdWVaWoCUqU4KYWbwPn
n2ecDdOzqSLtijQnjamHhkB6YA+Xk1vcQnBp6uog0Fe5TWBHs6M/lGACFK6dtSBz3MVtiZ8CSJEP
qTCNgScBRkgFs9YQBlqd7Scpo0m3BB5O8s0n8gIzVkrEHLwAUwWihvHq34XGWW3HHPodf6bweKw1
8r+yj4wYpQdpfsAykmgWFrDYW1eQkjuY0/546jP0usSE+c9jZ/2WDMrwGPW1DxFvEBjgEinqspSG
esfvCtMYpm7JbD4SuHsM5qYbrb2yJFeGtiP2dHm4Snc+EmcxOVuDqTeeZXf8KRYOQD/LmGq443cD
SGsz9ta2vTSgSRTbpCuTvic7s8EY3bsNThUB1nw3YZOZe4PqyjaF7WYI+vn/YkmphoGM4pYzkbhN
gg8Ej3bqRl/qjWIyjS/06TDXZkakw5G4qyrqk4/Sln8KudFYYOEO4d1VWYWjUo9EBwD4AWK/iPhY
h36C9FGpy23WD7x748CsqO9zjWL52AbF9+PES15eteO/n5wZDFEYjwqgpG2DDoZtv5GsSZ5zZNNO
J9+tep/W3SG+Q0QWtHNSW00x0ZSjyqgFZKFve4N9R9Rxqnjd901AVc56FporZQzNYCvQAn3pQ0H3
cywgjfcUhrxtEVOPMNdDVA2Whe4VI35E0JBfulwgZNcahOpCFAN7EJBQVE3Wfks6OrnnVb2PLKK7
4jSjlnVANRnmiEHXLYQZ8fC6x59ool2erFHRAiIjC8OWnecji9U4Kj2rs1yLngZTDeKCapa1+5pF
2jVH1gUhXAvt0WpmO6P9zNrhE2bNY6e6vjsp+TJQ9AFhrYaKMqyTKcTl+I0LBBzS4JmiUb3XiwIO
wniwHNwe1fd8CcPTW5xHloKQZbQJCKXH+GHPPRhjddqEV4B/rGyGHNPnMZRgWDtcV2liYGGM1qLs
IyDbI/yX4mi2aFhGl5hHK4/scFjXgiFY1OERbu8VRc4cinUHU5NdMAJ5t0BGssCNqh36iK9a/InD
5PMup9YVacaCRsEcfxiMdZnJx71nckD7YQZjOX1HZsY0ofS9WBdvS81nUZZ6Jw2voQ7lf2QeRsbG
6u2llBuHIUqZJVspr/OQ7nnEdyIC+v1Lt4x9KmOHY4kprTEKNBnUrDuqz4b7j+Cp1Dako3HsyIqH
RXFP0UdkEnMGh+Bcu7E7PU/cZl1jMCyzRKy6znQUtoaEJa9WHQSvNr3PJVCuPmsGJ/YXu8KHj90R
Sh0Pm1g0NSuHl8XO57OHjPeG8PjqOeQJt+jf9ZLBSkZUNTYh+9jTUqJczcZNE0Vke7ypxYuJoosV
FDM9qm/A2K3UoSaMP4Z48a2CijbjlUEH1LCNznXf5OfGi4foYL7ImQAAyM/wJ0wUz38c2r9Z/khV
yUkwT+LuQnIAV7mfqxtsOBuhzptvF3oIcFIi4xHvWQXRGWX9H+i2E7qwbFiTGFaiiLoSjmkKKsOW
0Mu5Li/019XIkZJttONyIX4VUvy6ttjqB5LDXH3/909tqyMwZU1CcolbSzU5Rn2NAglwD0CAm6wP
uRmLc8UlSAQr6EDxdd28NejfetqeTQ+PQ9LvISJ7BITwNL0hP5gNmpHbDImnd80GyoFZ4I7Ji1JH
5bJSThUOq6PPPRfS34Wc/03yJLCstUgx2rdeeGec2TcjmvTGBZDnGlPvnc3dTHYs87l6LPtoxIIG
1RHqHsFpIPSDFigadfXNty4Gf9oujcWjVCszjLqozqu0Ai0H51rStgS+zavWZUl8oKLuZiBLnu+V
cN93qbnFi7jWeJj5WZalohuNL8wVpWRW0l3aJ6mOgv3Nb/5ztcOj2o2IGO/nu3Adb2+t3fdW8OS6
SL8Yw96LFNf+KXtboMJSCckbGZPf7ehuGqMrVao94JKbdxNcuXUfwXZU1k7Rq4jKTVO5BeSLIII9
BghUv+1qkt5wj5p3Ehfi3iRjNHDBRmA7kaurC6+QJ5Rf5Y1I+HcpesHW7rqQhPpCrjXADaRw7lxN
LeAUX79cYl7D49Z0yd8hIBgO/jLYZl7GP6mH4dOc8M5NY1vkUa9vw5PDWpG9k/01JTZ+zJdQDI3S
v5xuzEUYZqRz+z9hV4Ubn5ibO4X8AtT0CWO1tSlSYgjE/Ib5mxpLgUXjwnjVLf+pumlufqracXiO
jjKgZG0QCHeNpHB/d38EelpzHekCxD+aka4ARB0UOTwU4hAubT4pN87ac/5OMinMx5VHkdUq2oc9
V3N+UAuWqoYXH9s+9vPha2UZ+i0U6/2dgYqzHXCM5/qm84Uk4byX19CSJgSyR9uCXjfNmdKEpzOh
5KnXMvxFtunEzzV1Q4axpaB3OGJkse9xVvNbOo6vb+3inTmDLx3YxujDJNChlVoIa8/bHWZ4rvCI
hQ0RnE7aHPpCzySh2ucZYcG9clTmGETRutFZQ/sC8x1i9iA8CUUj2K3cabud6tGLv2axy3w2wVp3
Yglmd/es7MDz90UvuFfKfGOKMqx6ivWl53/RmeifHxgqCQ6EVaVQV3Q49wutanrRXRLAJQ7jSH+s
ByWnE5lMQpBKeQL8fK3wBTQrJ5bm7x6NsaqML4Wt8w637+s+hCYdBtDE492K5ziimi+cBQ2ArzZi
UdQKz8OAIbf9/R0KtTzvV8uzCm6CcKv6RWI/xk9E3WCqnlLs9yFsIPBr8hL527QBdPIkixegOY8f
f5GZ8Gq10tq3If+usyHZ3AUBggTkAxUZj4PUdIj3Kvc7kpKs/71zm3oYXpjJIDAbdCG29KtAspqU
sqEO6MPH3tjIRkdetFn2JEID5CTQGI29lr75odeC+moXVVbOZHdS8bHwSN7Ywgx6T+6G7G3qLrvs
+4nIg1n0cATdBJqo/qaqS4Y/hcgeGGnre2wJ2ECD8h4F2nd7TS94Elfz6UbZ7sIX0On9MHlffHiV
NqKxID7I7oHgth2mEV91hMlgZSM98yGmsoaTcGRt3ioI7fawBX8g4FQVt9xUq9SrbKN7fN6MTMDE
g8AZTZel0M/yzJjthVv9ElN/y1DDm9Xi6XgEw0L9YGS+q/96VuTFrfmvLJdzzh/Wos8mvNS42FsL
4KgZGZ1645UdyGgxcVUHNIvyGK9I8pMaz4Y6QkkOnsxCbSgu2q6NZ6BmNLMmGgzDrQnasIFl2CKO
GeVPXjBOpDNpU7ajhGdzWVEpfn1OPwl3uTO2l1cM93GwHkDesiq5SI0au7a/VZ1MEwFFDuT2Jiht
hk9WF7hpaEMQIaMuH9lPIPOYetIygZpWaWSfbJ26BbfIDEsH9JmPjhqwMibJfMhlk8pCkVI1DINa
MccCPGMD8J/G6XJDalZAL9qC//06BbwmF32Nu+kakl0bogBzC+wo9TaWacXEbEJBtX2TRjqWfNgB
UJ7zMb2Mh6WM3mXrmMcb1/hyCYrp5sgmdUjIjEWZUjGK25KnEs19NwSMugLISxhomkjDIACA742W
yHmRsRYuFhLT200UnowjwdsFki0JJM8nbtFZt2TlURxTM3zob2goTKkkVhVeiW4YM21Bkt//J97E
4nhjiuL3YyJVodVpX+VG0j35557nH2KxmGQCO0iBA72iCsDbhWMlrvrMXGXll+Tje3Ahz8CKKctE
lMyNEhK7WLvt/pZX5SqG5oM9n4rPD0bM5bT3n0O10Jis6hJ2GN0zXQH7UHtrlPDyBvoBRyz51a1+
RF/ahTixRLLfs/UJsDhPvrHOA1jTazaWgpFYSN2C4wV6+c9oEAiMdo6+uhVZwsE3eODwjAb9z0GM
8+FW5ep5oN0Vm/CK8WrhNRvMTQB7QzrKpEPehOcSw6ydshmRFj9B7rAtP1huyGK5zVZ1gHfNJNmb
vG2K9r6Utq5SSDQvauKAIKmBMp6LVofQbxLBrpDJgaw3ZqTVG2Oq/mxiWdIhSdmenpE3Sn9NECcT
o4C4PD99qsGBgkICZysGilGojcuYBL1un0kVds5Hr1D5dz4kPH9uNiaLbgI4uEjVFEPoCzLlEDE+
uIxfqlFdicw1K1V2NCySUMbq9ShA+q9Y8wqWc0yJIY33qB/jBlUkmSK22mO5xGZXRL/4iDhZcnxs
w8LhhMwBZw1Hq/Uoz5uulVzxQWY6dHbzvS1CQ8BEs6AeNsiilnndPM42Dj0xfhAPqytFqm/Y1EAj
nHpL/M7US5OohpsoOJ+k+0hmcONvyVbX1f4CoygLLxww7XTv/dgYIVFs4uiVzm/vG1rLOtOTOBaS
D6u6nZBwixrY3NWC9dVY4Wxe7NKVvbq6D0gcMGMQARIDEMw7vx85Qr9kRGTQPAvBAbfskA7LTo6l
E7DR2qbToQiQLQGmXJwakata3gzqQh0Krz1t73kUmVB1KojPcVRh0CkrmNx1ABK4DqQKmkEsHTSz
eLvVwR0w+WRfvroJzrEamGzBTBFaKeqdTToHUD3zHszoELtjKhVClH6jKeDuhKP4VDXhIRs8dJV+
rbmTmoAdlZWOwMEDPM/XlIvgi5MwyOVPH83dgTKmY31D14rCOB0OZGhKuAPthVUMLeqy9Px4BgSl
nNt+tykN5vq4XtXqv/m97+9S9CsURkkIfiH3SNM4qbncAjjwikUI27btLEu5SlhKubwO6WVsZhRK
ctnkWVEMLCheCQ7/wWeHVXSGTgedANGwD4xQD0DgX/v56HC1tUzbmBsdHhlgYoECpyClH+wXmvH9
wKET1It4cMZWI9jZayjniurp6WGy2SUyA8YLEEt3fsDesZHsuDiBevd3GNbjwY5kDvw5d7hCXHes
qtkfWdttgiN6RwfiZtGRkUSISaiicwngZX5WKvCc8OLwcaBIL+j6d6aJaZePRL0vvOekMBDzXs3j
IVq9rdIrhXQH8qq2+HhnCaElLe/5TZJwFf/Uh5FeNBX9YpCX2enlZ/QPSqXZQ6pZPqpV1sS0GukI
Psz4tFerniMQVVs7s8D9eM82+hFJo+yrqLUlTh8C2sj5/6N1siO+6bp6UDhCdxSbaFhHaLIHXQi6
2+drlXZ8HLEVvv/x5Kg1tCo7nHutYUjuc2mO8RWhTfrWsC9r95NtiRqfQZskLQ9tgtS9pa5PU+OX
TzxyN7knLnqrCYqBf2Ei9RuVod5BMCL+afvh0TKddm4bPBHQ/vp22Dj7K7R5PeVAB3oSYmgvVhrS
fx1Dq1OCpOvYWN63U0RewmtvRnrWYisb/sM3wHGCYd9F1fWmcJSbT/Dx0g29KtnP//zvY2x8zksi
8XUBIT1hrwkMs/ebuOWP5EFwOqmeTyW57yN/eqE/0TiOW9W4q5M5TAz3dv4IIN5uh9tvpAHGdDff
AXv7cjdjDF6o7uyxn1uEnN4BeADqCoMt7WHUOcEpNMZmDg4pp4e0bcpvNKKJd1sIUxIYo+rPumRg
Z221ElUefQSCLmmmJs3eeEoVaD5WBWGbzI+mcAAuZEgqoeKvHSiSYlFRw9lkh3937KRenb5hD6HF
HSmuz2jsyXje4stoxRElcaNlq5kNxY8Yczj0qB29ZXbps4njfT3e9khn8h4u/S/dF5iwVnkLXJBi
TUV4q7PiJYwUDEi2K0dFKUJkEV6gdjFNP8xVBIzl389pXxMyeVU2MPESrl7prYOC99RkKTZcwu+j
0Vq0MGOZtVDUdqqOan14UxNAFvvNZa5QdWfQC0GTq+WuUXRxeuPrt5pAdDUUzbP0i5tqT8R3Mizq
Q9g2r+tQT0FKkk429+FCaAMRhOi5wKP+pII8mBUrjhvYQDJIq1QQ01e6ggG40E5cVA3q/ESAJN9a
JQBUH7UYJ/A+IqdEWgO+AByIypeJX8EHGxhZ0llGFiU8LOsidZhIO06pxOXWCULzXpgkkQFrctQk
qYwnEQovfiWlwFy2Cwuzgc8q45xMU3boZD6BVbJSAsrFxwlJQybeBaqlZ/WPRTSV55/hERZO/NiG
Em8lMCViQWtgLgOX9/orxJHgXA3s0+OYJOLv93R5Stl/FzzGLpL7dVi3iNnyz39LbHPrzZtyRVBU
g92U3ZFMGSEnsxV+XKglEZiJ4ea9lVgDg5saLTXt3z1fzyXYSrT0oJEtttb8TGpUgWL5eEam5bYl
zjsHEAkvKrBlqGOnh6bZU5mcAkdb27GI8blvyrGnuGE/4kXcCzq/9Q0cLkhwFgmTCpFxV1Ji79kj
CyrTNp0FYiGQq0elaHtVlHdQb8AE9xL8SrDOG5BXEGQ8ETNHGCvZdu9aeannHUQl88KWA+8+g62v
YzXS9J3KEuPDzej65aJROcMXe2y8jKobmekh6sb8CH3tAf7dLINRAOdoBq1HJ9hcWhK6Z8B2c2kl
8Xk4gdBpcsGh6buY5n/NvZ7yz4AIsoW2O5nYETBBK9NhPh2v7CGcKyyxzlJloWlkfhJOlJFx60KH
JBWrVevvl6/JE1aPi5ofNEGDdxrCbceibE8VG6PESAr/oAVz+mXuPAafE80z5Mf6lGOfLlHlcLcm
1vtRpb0Qa0ByTUniE+8DcuuUrexxRddGtK4KDCBqU2YmrRjII2GpfTuKqT6sw5pMi7yMMR5I1smn
FbFhCJDoO1qk299/p/uOjQiDR2uY5qy7uqk9vkNSoBNcUuaxMIbde+CYJeouQsBuDeG90T04vNLz
u0WcbWz+oB8cNk+v8Xjnz6tRz7Y4A3ZpJ5hy/6OdN9dOJxOy6845A6pRsseQFa/ELavbewlY4fKb
nL97W8jmBxs1LPg0vtX6HZqBOwpIer5fQxUKNuhxZW529IU+L1gTwer4ZmaXvQB18cblRf+dIExj
1IBn4SApmKs3MN4WDtxjmBfMitggrWZ6Ng4JwMvfVP1T0tFxPDw16ZfUMReGPXooiKASwN5YXz6o
0b+1GyXcATBSsL7QOpP9kWCY2K2ecjLSgSgyPNIhTmEVxMNuXf69+I/X1/KeuLbkk8lxc+H9nCQf
UGY5qbiYKdBeebftjv5nWNpBSYN+r0gSHyfqB6R3rQwCQWe83MVqg/ZBevTFYyQybS7VFbEq9g9Q
jDM5/dAZB3eSeM1Le+mWdf0JssOMSoR5gGwKQ6sdDklFcFCUZNOv1xHY2KKReqEn7OTtpO4YNfK3
ySCZOCQ2c9IOX/hvw14rVc40JPkU+zHTmXz4jRbFOEKb1cnHFanMRQM6bmPlZwJ6NhNDk5y2aWdE
vaQqb0W0KVZKJ3+CtvMqFTNaEAs0sQm9s0GKEJD+3ViENiIQmj4gwmQmRRjIeuqyXkxRQ3b7jnFN
65VSB20hB2cMWhRjHUGLA4MrBa9fWtRQ8ig5vMn/888rVm9bzKmN2PTBjT3UZDzTKFKok0p4Z0IT
gseccdy8e0vlyTHEYJ77Ltnp9jBNYCCRtEiXaztEqwfiMBnNKoBvGDiKdcnSUeFZUeYx2KWcty2D
aODifqzFCpdP/SlaHK9HP9lKuw5Vs1E5V9EYyz5er+o6eIsWqEnFLgJg65fkb4vpPw6cGoM8/QHs
R5O5vI3EuvBrw/BEsMMWXmKc1j4L3TAKlBc/KFZ8rte5M9C/x3vmfZcTuvYAqu7/KnUOnm5feuaz
oywH22ayPjy93d1h/O26nEn7tkTX+T9cvGuNEcp+hPoyqeu4T5dru5/QJpPtriolZjBmMsp9pBiD
e361fNv1nMIo5UuZYuyfAE+qwNLWJPrxf49r0wpESq0E77URiLceIBWfOQQkiWo77frdjH8uqlaL
Pre4oMf3LuxelazKPlKQ83w9a6A2jwZZ1bkOcH/Rr91ImqNesHtO9x8Znw1SjQAqLWX8aS/NJR6M
SWEcEddVfZAXKBFnvhjjufXH0PxqLqQtEwk9nuCJhtuhLF/8PEkTn3XaV29E3W30psBI04RI4iuC
zEwyndCTe4O+PBdbUGKP15yu56xQNKkWWjRh5sbEu1cac9jnqx3/gbtMEvAdnUTR89sBXIuBilEg
yWDBSaZGrZ9b+O/JZBnqJqajkepoTCWeA9WljR14L2h9X/NLvAXbV6CScY7O/6RwXbqR/1TYYRL+
Nprw2pk1HrLKJUc+wsrqP4LIcdrbVZEWlEWQu6P2LEXgVrBTa7vb58sX2l34i1BigP2LadNXHBmB
6LnTqc1htSSIFRPzgBd1dk1xu3FLZ+C5YE6vIG+AHa5RBvMIGZy+pSTQjBwTbVos/C5LvIFO0xp4
AXukDdY9gtJ0fHSAKLSR5T3/3aZ2KAszbBOHeBlYQ2GgsVTNOYUr4xVhVWaRGocmnCR30lbyJX52
wAOYEXVp6s4tpYzcm9OdqaP4liGmdftK41mrq5nmAUQPbUe28WIqWpoQBEq05oLBymVjlJRLRPds
yqvhsxzjqkp9Cw1QVP+08tCTKIJ1MWJGiNcJeWMFB5gFnz3NPcwQ9HFXKQ5r5F+j9bErRJdBebxB
WvoecCv5QQC/AfQo+doCHCFDoW0F8MiymMahi0D7dTFO9tRD6xjxZCzIeJoWSqYjkyaayp+OcjRp
9gS3u4hpiKcxbYtSkh1c1jdMtH6ObGuUkChpxFcjlnanQAVazpIxeGPODyyk+uAn3GL0ei5rDYXR
TJ4bOYDt0IHY7is0VIjmoclorzFmW1z2ZTa7L68+EhML0n76Yx4koEhNDsUaA2gNBVgHVujJ4bBC
AUZOohIzBtS5OJ3zaT+5Li4N2UGeCfXgBbzOfkpyp85wtgl+zHmIl8ruqaNueihzG0M=
`protect end_protected
