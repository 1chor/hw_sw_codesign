-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gLGHdsV180athhFyQt/ZzQ4QT5Lu8bPE3YSdyN2/oRNIFQ83zs1AkkQSaN1nXuQx
nk/VRnr1HonjTEmDdyxxRf137gLYTnrmURD8+t07i7kC2xSFkvwapdmlsltS+Yfb
6TPpauxFkX7hngrv1vcqjlgd7Wk7F19WS3g3sZLX4/I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 3563)

`protect DATA_BLOCK
JEHrklFWeI0fgFD9GEJeekd13qMyEAne7sRfdQHn+y9NCZF6hDaq/jCpogActJB+
pypkocxdl/9SW1pby476A68PwBxQhZLxsPsKHQABRVp+ILe7N1lkmMtFqLJ7ZKVn
eEsd8vmw1LCjGZevuj1Au4jr/NxGHo5JuDj6O0PIK3wG0vffNOdxvchkjpgFcc05
7sd5BPtO+CV7Qr+n7V6LgqyY1/pPD6qddAvUEvCOJzZjWbGom7QyxwhcZ16kiqxs
XMAIEMAkJ4pr17gjyk29akQ7+LKz1DAXtI5CxN5+YUD8bjh5zgOEIhGKSVQ+Tt5T
uMJYElO+uYXvyDQgF0RbEDR2Iqb3hhUTaS8OLA7IDwq3Wj+afeorfcWx04A9cl+C
pJkx9gOdSH0n8W+pi8W5Z4mKmJth/hYyMiYcwqqwQgIYh4Lv/kCKFlyS7IkI/AVk
gs8SHR7E6PIYO+BfGIQ1+j+OSwf8tmWZza5jqwIdBfrSRTY3vRtroijt4gD0ZL2y
eVtZ233Fb6sDRXG95nSkCP/qvX0VK8BO4x4faqUdBa+zFP8HXdBintIBqnLMIBVo
BHBqBn3WTHvWNRBVxEOzzxqtcBgd6aB+qSKl+21rb0AjoHe7a+uk/KGo75w0IBQA
L0hG2TQ08ISx3aHaZMFwnj1gneYNWEPIh674tcZgfVwxfwjdeDaT2u/pZQu+LLm7
FUY0VeZ8aXJoBeSJ7qmjejl7nJehP86ZxCUtiRU+uJmw83YKV1z3ao/gk0/hn7IG
MhbMLwPyWMiwbRAcXdJYyzctVkYXHpFSskct3qprcJmrhB3XUkPcaQiTYyNl3jc7
idhIayVNnJ9waS0WYG87tcAxlGV9SZL+ZRKgeZW8iW1oBM2xz3Ipz4AopvDR9yKN
7EF2oQUnwvz0YzttADO0weCzRXdqVagf5ZisHcvebjE/c5nbXvy+rr2OMa6lcPRs
llV7ENZ30h+K3tVogNz2I9lSpFUfbRaKNcPPyfMK0DXq3ZMbWmZ+ky5skRZmStc6
er+HQBi61gHSIq9m8fiEfXIjT2tCgQaett5vBoX/wIqfE/ZWebDByaaKMDdE8dSa
zpe8iRxZ2hMJv1nhszbJ5sa982aXhhGGyOBd31e6BeYpR/ZPmi+lLvZ+IyLfT0xO
X2trYRvS2eATsVxRwmBVuuDEMSStBHUM3+jl3jKjeLIMgl0BUVBfhdRu8XcrMumX
JwKBnI9garc6zg9QOSRDk8LkyvIWz36TmEOxkaHMoOjXdnIfSbJKLiwmZ+3uFDjH
Zby0cXQEtKGhq5B8dnX+ZX4ez2tfSttiWzVcN4EcwTEHYLIvQ/66Yv1Q79wp8miK
ytZGrnLxJPeivXY/tsWZvRK4CWn+tVVzU8zsKxShQ610w+Fu3ExHd9k9QchmIHIL
U6Q/RZrjBkdq+dLVYlcgx0fW6XAxbkoQl9V5yj8po8/T7dnrf+C5hjiSt6qDm1/w
B631whPwaRekXCoDCvFfCnv2q6fqTo9vZn43+mmPuZJjj9MKv3tEEGeZM4hmlAeI
cGvAQ4a/BN7Z2Izux0VJ+RfDjzKBrudwD8qf4l2gqCwqhFGzsukRvpw7qTYTCdqg
BLpUO0hBeKhARgfu987mSmU35KaFFsatcaJLoKdmh0BoItWOR3QFKD/yoEBMduS8
8M+gbec8vVkxNlg6Nq6rps5Sm1PwUOOok6D71ObnyMJgLOpCPry1pz5frHJH6coc
VqEbjFkcNlv0eErcYQIydYZhmOCaZWNkh0obk3f8GRYmYmNPsKT2kZInYPpL8RHj
pKJuBNWsX55guPwwbwTaUMWaal0eL6wK+fN/vcj8bwIHKb7q7GLZevoxVrorSZMs
7Pe94n81AiCwmA76+IbeGbfGtPx9Gc8WhaA1a5Vbv8r8mJY+P3vPCXzpDNKPnm+a
gjUk+sZsH7+HzReDeQMP9u4a7C/4+xjcgfVA5WossTFu0VU2Bk/DhTnVZfoKRHHE
TuR/CJHnZJSz4w+P01poDIDsuyAUojGj7NOzzsQKa2DGPBIi8FKBRmh279u1ks7S
cwisU6tHe1JKxtYECtlNq/FNTFpeyxD8Bd57sWWrnj/O3DLujXPR/ID8nOhCkZWx
FEM9fVb3ClwG8kBvkVEy70i2pHd0ZOiDGrGYP86/IDOanUrMDDjsNzYkmhh/ZpHe
1pepwCiRYqxb+auHymW/7x7qJ/YI8DE9gqozrC+p2U/et7gvJQ7RRdkNJ8ZR1vJC
3KzxtMDlmNoPtzqCGXYh5UNFjglJ2dEhDeElI0o6LVLcfQxDoD/8gkrfezN7ia/V
Xbv8xwwXCh6/UKgxqS85rnJpIKk0Mkk1Hrl9fzVzHfhLXh7S1/8n8GHoxWTg1g5X
C8IzpvsaARn1/a4YQ6Cqp+byH8Hiesw7IpuO/wVQEz5pDk2yq4IlpA+bQ/BOniia
4AQ49sZnI6H5P/Vtekhblz7oigc3HKoHKPKGMNJmMUm32rYUVfydZpHfMX/HZhtD
BP51us0CYNQDNNGXAvDuU3FyMT4ik6aJX5ytfZUULCZoTUFxnTk4nS+zSorsCBeS
2xGhJkhGX7AEiYCvlG1a7qNRpNuZOSlIhEsKEzv5Zm6OIYKPm9OHb3vmQ7HJqG0i
GM0D5Ntba+QS7KxI/QmRQHSIZcljKzTWfXumicgJOvRfAGoQXg1/Cdp/ue5gqKb0
WQuD+rjIRgIzb3RBrTgFAIv1YKl8yg5ruqkAvjYn1x7MeCKssTpv8+QFvPqSwYxx
P5SNBR10yDCyhTjuiRayUL0qZR0x4j2u+ALEqNWzB3/R/M6axAcHGTQ/dkGSwW9T
6ZG4j5Z0rFeimzmqQ8/PREIH+d04MKdnFd7W4xbZM3dMsjfJ4I0vOzkcB1PSfynd
tFXWYyNIXJ+X5vFNlKPteLsVWIn2fnXBvkVxPah0z2m1LevXdYRSidgTa0E1Pjjo
L+o1hBxVKQah4Dz1hw0pPFRq97mACJatYkZJd7jBBP0/yvQyOFFnZqJAJmainy26
Obx7SBl6nyEcttYyW6hFpOtjrkRPav50wa0C1zKWazmUKFqmfAcrQPbshb/IQPvv
nMC2lRh9EGloFJ6b87KAbBB8XDi5PQNCv8SrN0+C2SjC9jm0QtO7Z72w+Vgi/SHx
/y3jqv2Z+w3vm0ltEB23f0GusnETnW1WPRfw8EDipNLphCMHTYGOtRO3mMp7p9NT
krBgT1aKwwg2acBJ6Dy9PPRzm2eFNORn9LZQmvInz319LFA+3OG42DWeliOdxwRL
EeNs4/miouJjhyT0INg1QwkJyitR4kwt2sx/IAP8M8BHZ4+O0CQGU/3Bl+E0Ptk2
FRhjK/ttJ/RZ5tgW5MKJr67cA/7AwlMkol93gUf6Bltnt2oFlyV7lvA4FIH6PwDt
DgWlVkbK9Ty2+dY5A1Hfmy5Dg7zYNRv9a96ndO29hZ9CYhxD5zREZmsiwW4l/r0H
EKJ24npLAu/CEfmGUPI9xGJxO5M3gqNFc3f76+rBEmj4G3s54GxRiJE43zCpAZpH
zj33CZJC8RzNF1zdmSTs/F4Y0Pt6GSMprPNS2AkrdfMTXkEgs6TuqW7ib02LjKCl
ajPK9sUIsodrCvmmzaejFzq512Vz0CiBXJwD9NdmXp9vNWO0tm/Y45/CbqNHA3Ld
pglKOBvsjb/tmXCC7DiwIWose8qlEYK8AyCNp98CYc5Gft770S2N/7hXTjXmOeo3
ewvqheL9R2FBY6oZVfbohb7QyYs3nnMDHzgx/C0uLhhK8b4YiSWz7h3R0CdVFKOt
dJW2VE6PYRRL+9uSPR9XqkNMMZ+NlFR30y6RVrPVkrRnv65AzmfZ6Y3oQExIu/Nv
V5v41uqegpGtm3CpJmsIIfv0AF4azsU+UC8D3fhtbA9a6M7z3/NcGCqV3vgLmYvk
i+qx3WDS8PTDvb/FpqBOjgPS2odc2ONfJ16xqFoIv/GiLLN4GdjkXNgQCD0A+m7o
5ooPocusZFxddjs+MI3Sr8rtJv7O0z3+vTS+U9lCwrDmPB+WKoLQEN8q8RaV1LnO
THUHiLSEGMl3pnX/02gDe9SbepX/APyiWlJ9IGEMgIc24Iw46zB2+/XRDZ97PsFi
r/RDvC/cCmCFyuI3AkHqUOcpaaA4U7OMDX2vLF//KOiO+FYYXgOWxmYAkWTQiFQ4
7ggwGnSvT8EbsgHB91M6lz5a6Je4wx3axYmYM74NMPgYv8XKDcjCXqO8BQDkuVAV
vqoUswVxlCZZhBgezUNTQjDLdPYXgJaGE5D8EI+nJAJc7obs9XOOgExuK1uEsYzP
3fNMW0Gr98RQZw9cnngDTtULKnKypvdVf//yC9GjHpt+b3cVP1EcMYXZB3o5IARP
3ZNbXTWz8QSTq65HUUsNodnpn00z+AvERDoZ7N/h6K8w6gtGmJmH28Yf0urvJZLH
PZHB4NM16Qh4FZHfU5DNB0gZtaXwy/5wesyzeoOdGtXojCvqIc5LCNw91o7l9VOn
Bop3fFcj3NALETsbFuc5nWRzbzXeFxZNqddIRE9eFbcEqG4Llzy9nnFT4WSRbUjv
mbYwANYY/WIdB6GzbN03kmCF9F5XI2epaFCq/2hAwgbyQX8Dv4QhV4Fu+Yk8snun
m9b5cerLi/RqWYghK/k+0EwT1jBN4PVhAz8YrYIzIRTo1tiDxIASINf8a+s0j0k6
1C+LL+nxQdAUDJ4r0RpIJofBCJe+gsevFGBuV7j5d/b2zVJvaKvfdU34Rt3SO33r
/7zhlW8ZAGngIgIZB+TDGXiEoLItlBaFgp5BwwRUZvg=
`protect END_PROTECTED