-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LcpTy20wTbZqmJWZocX6ogcMvgmSjJy8PIXQ2quC90V8ULoJ32O4sBMFrttXFIctliLDzDD8McEJ
Xncp4DE+CDkQ4G9RHmO8z4C1jdPSwBoBGWPL1RmyWQzAObsYaHIddiISqArMSZBDfjdt5hFUdKFF
KdZ6zdSirvL91YaB2BEkzO5gEWRVGz81Q7n6trsXyAPURMsQpjzCuI4KXNJ1aotuE2CTIZAtPCAP
LuNsIf1XhpQzqxQ4DxRdfR395r1v7IyNGtfyLoVfsGVCH1prs2+iyEOMAcxUzbVfEIg7587cnyH6
VPHxBqf9AKyZNJr2uL65N1lC/hwyLbL7Q1z7lg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14336)
`protect data_block
Wxtc14z7370hTvGTMzrqrkryBn94hDW8Nxz1L2FGCPMhJyBShtAOAPW+n3BqyZxnhFzTTYy4Yz01
7a3Vci39hori/g3k0ZHxLaYlHaP6dutt5iiIvIcxkc2L1knURMAljeSFc+F+r93/0PehXwFr+krL
07A7sJ5DzRbxlUCJdi9X1hkijZOr43cSFZRf/EEy0ofchngimAW86sZmaJoPyMBe58S8mvo+KTe6
MtVtvrpt0OmdnNBqg/lignh8uskAGlfM8Scrr7EDV0Q1gjCNwVgxHNkZqm/OTAhZx8hMGDD+RhWx
s8dtqPYoGmTC63p6NBWG6SzoYSTUfanevqtbblPm9I7888GheWejBB5T32fSx8l5nl0o5mmGLLo0
mRkDBeY/Q4HtkfH2IqpUtb85E18aBZZ6JSH11n7Fog3gmdpebMm+fKNQLkO6RSS1R2XW8DfPKlPJ
symtR9iAxXJd8PrnTxU0yX/JQ8r2Xu2vv+S37Fvh0gKMJX3Uhf5JaDE52QgOl1eszy/WZ7hyRisD
8nXWDi+ElHKXsb4EzH316zjVFkDE8O7CWMtpr2cLgDKQYlve/0fGCes1fT+p0P5j2T7/rXvbAkxU
dALZNMKotMaX+CXdxy6nVagQ92uBgrnOGZQPJzNhCVWyFBOIg86v2Sg/MlFAIr/4Js1RY4CToe1P
8fKikSGLTI/le4+CDzuD2cfjem3BmWTphnUpMmlEDQbqBw7OCOVG2VWNUPCEGgmYn7U+U6j14OFq
T+4v35gG9aSsXa6qdai8GR4NgSROG1U5dPsK6M4lSGknQDbbJJ2aftQfFyd3RZY6rJ+Z0oZilhUM
0ur7a1G9Ng0D2i13mBcB4IzAkQ7PZdALHx4bn09YSz/zASTjFr62Ax7C5VRoFiJd18o0gmwhaCXY
frvTQvio7kRERomNBQ+k9dyMrDbEdzNEq7jrjY8z9Mo59ODqZqejc01fHxZHgPEbcTuEtfvEvuhE
7I2KZ/zPYZbKzWEjLLVI5bnR0Y+rnLaNuI6sd0DvwPGOTqH+Gy/rSLDqHCRFNrCc/P+zkB0keS7g
4mNXir/q7cbVahNyfyBOpbi3n4ujnN+w21h73/dw3it7f/OefZgtztvOX/3wtwcEqpXJz4VZIpp+
zJjRiKwP58vvPSnEqNZ4lfzJbgjmEUG5c86DnzcRIgkekgjpkHEy8g14Dt1Bag+o+FF9Z1bNeQO/
SE6ipj9MDNLnac+Bf0uHrwwIZFKfJUIRVgJ54UBEVTsXj2l4u9sok6U0T6HtbXogS3FOgA3/W5a/
hQea6d1wmlessahL9pg4M0e5n4EnKlRX5ugxE7ya+8UPyvGtqsQKyOzfhfSQvRENiMSDH0zqUzOH
sIpjM94iHP+luJNwrRQsOAlih9jM/54cniJAUuo27vCvD1zkudT5F6Nd8i2Z+KoF6jdOsh306p/q
0a6/rVdkAqlj3Ie1uXvZ2GxYjGF7Dxlrh1qAXmIpmOia4aaB88ifYxhucwFwFLdtX1qOP1Xl4ci7
tjfYp/1ECnLjMHT350IBrytIpp4GWZpKsw7L01frkAKmCijB01FEskAzni6683HMPfVoI11oxemI
g7qLbjRGhNOC83u0V+F0m130mGWuKGAnfosDjIKv6OtvR6K/fYE952DkipfBb6ytRC4MGICyRKnr
O//3EXv4NIqL6cypm12ON3NmP+sL/wgLJstCM2xhuDUD44vji4G2gFYsiPOVk8iGvGpUBGvXyc2m
9iYEUmc8+Jxs+ouvY2vkJ6KlfS/b44FZFQZTM2WahbTv2RpajXl7x9ULmmk+gJf1Of2SVinbYstm
V9971zrKIEKwOurnaOS2IIC8p5eGwoa3vsEKOgBJeVXxH+HxPVgVASpieQFu8RTCKIk0NIWR0Z+U
5DbHZmAIOc6wTo31azqTuID0YIXSPGXxrxthMq0hq1PXfCDEG7jmyBEdft8VDjd+d2nx1DfUWN3r
OqWTdKOZNDujeAEjraA+KDOm2OlP0VYtWrYUV6yjzHlg6pLcLcajIhUxSApS25vGU0sWB5Trb5xm
QrXoVRVduyRu3UF/OU9XTs8RieN22vx3wzhYMjfQwQ5BACK6PySz17n3y4e6UCKsYAmvqo8gubyf
7XnILFNutBJojTbUIKiMjlMbElPy9D4wXOVfU4uzmNGQuBR7FGTFosP0xiKZ2Zlrf2HOrFsCEn2B
dRzelK5nqDPQVhPcFvV0ANYXFalrfUwBHJCeCJPlzXptRktyhsYH+T4PIUQJcX8xsIuCIv4VgEsH
ozXFqllGvyYsfWvbPMcFDAYrCLoeG3DTmSs+kdCy3E8JFs0LelyfURe1FRak0rIoEfSsUV0ja9oc
1FDFGt8+ZzdeZxVgiHBFu+p9DxYJQUbeWax1SsXhZ4640zMgg5qaj88Y+3ykTFzkEek5BBq5q3cO
gb83w5BeIHXenS21Y8VSvV5hVDln16eXE1X4myXDPUyJWf6V4/lE9AZJeW5YbwknNJgaVKcfUdcM
rgKnAC+it0ngKDC6P4bcxrMAP8P0OD8twRrwJjOIIvOyHRppDsZwSC1Z/7LhNjZ4mQXiOMFxRcMP
dhdN3CG4p8vxTtGFV+pvPus34lSUyD+hX2BuvG+T6OcDdtwwOK1dWrUH01inFSdE+zgF+CniNJnX
pAr8rcWYQglrxNd1JSFuk0a4gHoF4m4ARVtKmo2uKQ4TbsXruoTPxilVJ2eFm7/m6A/0TuUx/Ch7
N/3q60wJCNT5M+wXGdFxNYUyx5eE17Ex4MNZwIcEgMEpLTWOPp+glrLB6/4KT0/7m/M/n9xyu7GG
AVtX86IuB0w/UI+Y1mVJgp29yChnDZmBnOec6f8SB2Y26KND1fK3vZ1Vhkj/SqCikbPd0s+o1w33
5r6aDtBCvN/1ietDpYbkVDzH4qdiCfHrgHyrTjOYcmIx9uRxpo7JDu3WVbPx5QjwmDLIDKWIVCfn
Xja7oaOSN9Muoyw76SadBjVo7Tqag1ZeDq61hxB+Y0ld+wUn4tROQ8J4vg5ulrr3EE+iVOfr8jvM
urGBwUdF9V78FKzJp5PKdxVYzy3BbBRmXUXOwxRjWM1hf4vcZ9ROYYnGsEBRYPX+EPpExYUbufZJ
T3HmfikjI/l3q6pDUz80qj+C7UkAu9OhWUggXmm3UwF6V7R4RM8xGGvwxrXiKDvRdKpwovnNgD2L
Dz54vrSDydFwNnrgy7iNJ8b+lRa36+sz1dtR/D4DC5BGQVh/ptI7xnpnEMaWEqN5YcwAe2vh0tF3
Vhd0zQp8BGLUTEM3AE4DRu2HiadC52wwxM7lHpENJ7K/1IPzwjRe+MFvPk/ggE0WyHWtjUVwe0TI
C/XSxG5MzRtQvrkrzhj0B8UNF2ePPEu32nTzLgxg2qolhmAxLmfQV/CjELbu2N11ut/zVxd+3fvG
dqfhuqSfEDRi9G4CdUNzVLFb+pQi7s/fzlmwX+d+fvLqCCjIf+HQjBBHYRWJEO2/uqSIuE1v08Mc
WTsc6o0VEtKYRqn4vuC0ZKQTnmzsIhpSdNUSo6SP7xHCzPXwo99JbV2mJQgHXKNtzgrGWwqsY338
slpBKTiqSkOlDD8PviYKaHB191e86uoubvi5Y2WHEQ9VwkmJGP2psoc/ltucY4guspilvSbA2W3F
oGMVWdrO7WyL8LNJvqnN3KHscY7EIS4IT2P4xXLbb+qTKVR6qA3jkjxMxhBQ/GZMVDi+pROlR1IY
Bwh4BoAtrRv46CsXNfinpwsa+eT1lSFWAuhUhkmudkSWeUptGBiY4RalntYmeJPzOOyMWOS1AYSw
Wzch2S1oETQBMSKqCtZOth0VVb/wu1AgA9GnBTsYsOvc2us/6vqpgQInHDmbUFyrPmDZzNniT7Mv
9Ia83YZWTsUOpG6eBAA7htMFgbKZ4YvK/wwUCk+zgI7AV5GrGlkCGwR+jKs1fG87yaCBApDNdkX0
fo6DVoNhW8DTyZN8HtzrIcrIaApr1iz6OGVcwppUhFw+phLxSAHYyxGNULgq+Bn7djQ2GTHvypbq
UPKNYdB0khAy+KDbo9YJ96hpRPE/0iv4zAd1TcFlUuKXU3MnmI/n1q8QyCI4dCsyl1cyOKc9DlJd
rpz0eTMupvcTjSr+Sh0oa1NjBw0xodDcMywVN/C5HwD83SZRkR6iEJSJg+oSqdjpPYDelxy9KKwQ
bvJ53hnkoNey/UNPRQ8aI1qFYcKBf3mIYI5ValQgjsh4/cAhk5Eck/L7MHw43+bepRu+5kXhrLIl
ZTgN+9sokbuHX/aCanRTUpfJLXvIV66v+UGtTA8eszk2+JUrEkEli02fR6OeaT1Qa4HIPFH8XBnJ
75yy0HPKSbV7Gjug3y/zpTouHCaXMlbbTxgTh82yghGWuyjUgk/fle1wezihNfJR9wSkG8KTP1CF
FhLxleG0CbnqTZtV8/CJaFmB2+t5ukG+FnqZNTD9UrgLjqQkeVmle+cLqJbQ1vK1VsRE/qrBwI4L
SIZcQo1h91Hho+tBDjwLDx3oSXP8hKWjrwo0t2IcmoYMYREWzQqOj1v46jPyeQqgkoE6F2c6nBwy
9U3iY6RVayH2M/zY+V9NtZOKDIU3RrwIo9fnGyyamwmUjE7semQgYFwLXMw/n0vIH3xiGTNsaMtb
M4R/pNX2JyDDUcoC7uB4uvmLvlKTZCOtHMp2lb2pu8s1wy4mQ4oKHPUTQnCFyKyBXN+uosx20tgh
xbg0pAeuszWcfJJfduug4s6cDCBimqehQHDyaZcNoJBvZ3Gb4a/OY2+jYTDVVOoelgZM9ZRspuBg
9TFlH/BqFO7DIPDvXFXC4Yym5LEssW2i9LCvEhBojiH9NjpaRKrzRIBbZIMexvWw1SUll5x3rpj6
UjrgEuhXRyKH8ikzZoKY9IKtqyMphe0cvxFyX489cM20RQqF4g3aPgXbx91fTGVGkm2kOnS9qicn
jo2ZCKcDa2vLEMBL6EhTNj95MkOyFGj7polSc5CtZyN8tVqg0rG2rUEMwUIiuPtsC8TZUgOblTRE
ekHPDQZ+8Me+obRthkR2t7BnsisUlrFcBVURP9guvoyw/A8BKYIVYUPCwLGilcn4ztfeE2h71ZBI
5QnzZbm9YeKqdHoG1+hDkk1fX/Qk/Yqzo1/SSYkdptWogi1CQWRz24CfkmzP/ycguVg8ORNgra4V
B3xB+/iIoLvnhfYoQxu8po5EwzLBU13eXuJOrAABJRDgwZFFxQ3ED8ouzZgH8nsKJtk+862Apxp2
si2cvO8ndbgevrF5zdKkB2Bl+1edlKNaxjQkqJ4vhhYTKiR3SCtqEWYOPSEchxKML/nXtTutwOYg
WYa09ls/xVI5outjbxUnAqkvUr3oTDKEoU/PTTuNO3uU8Lb9zTSw1I2ST2tiEKKRC8agLkaYR8tL
F5w7C8EvFrY7SSe2YfIluBFNQ5lpbzeIjB9rIZoOTxPUVwKbPUInXU+mb6nIVf2MjCF3d5UyTRuU
LmZuVRffZnYP6mXqMZg/UPatyfvmWNBkfztN8Axf3sjZOcKdQxcmTtCeiOM/7vJh3el/k8JaLx+E
ok/uuhtTk4VIgcG0uEVpf9GwR8q8gxQmBCcXl47SzEXwiwjbl2g+XuOQfU+ykZ3CUVpFkWdv6mtI
r56FinTO1iBWnbOE7Jtd85gOi9JLGAfuambTsUxi6mDP///hEHNHpE8PORWdhlroxUc0N2r6hp7M
Z7cVdBWAjktoUx60WSN2hhr0O7Ps8kaSlpu9ODT3MvSP6NtnnzlA5ozCtW5+ZcBLsBrSKbRMGDZ4
+ePvFtTCRaj8ETPASLUlBg3BNisKgegVY1Gq8vhDR4VF+w65AdfGiU90iT4dJY/ZmAG515Jgu2ur
o3pHY4YvsS6SHIzu8TXo8phU6SaXnw0dFteN74E7NvwJLucs/GTgL2mcDef0a0oDL19kNLN6ol8V
P6B7I8Mr/Ym2io1jlayBwD76WlOO7dsNEKCXpPh41baF/3hX0PUW9Tju0or5vcMfA27hBJErCbm0
q/dJtBLGvfmmajEAeoKbxaDpFb5HiLE6+drD430EpVfklztMb0PWWE23ExthV7yZPqtRGhMnfwyi
yXLK6i9OZbX/idvMernLzcYIgp1Wz8YN/cvhsy28fnvLlJSn6v5yO9xXoJjRTPVqjeCRICQha0Ap
StmgAeNTi/JIkA/3vZzK219reRp2U6HJawDBVLn/UiMblY9jJ+pr9+WRKTm3YqakYqYsFw37+hSs
wjzPwm27hh5AR87rPlP4BNSDCtHts7dCCT8KpBoBx27jbkAVamvAN+sk2CqBVFk7JVyIEYn8A3j/
pphUcJJHWXRyrGZgV2/NXj5BcJJ4fRY8RS8WpkSLGd6gH3W+6j2kVGBOrxp51A0wTqB5xND/17Yb
zc7UvQh8eXTaBkUB+FWIP/aaLx1JyDw0c17tfQdcBJLDyhwGBaFcHWovQEiom4v7NSPM+F+BtNye
qkJDlXJIrecVK1AJ9IviY5vqlGzLDpklhz1RL9Fl08wHVYHn959H5Qd64RLAuFKF0txzTKUSjiki
btbZwV1546K20MBy4B82yLTslpy1+ESh1pe/tQ1O2f8MNTfi3ZU1DcbwzwzCUHm0kDm/H4y/WOVL
DY2ska+OClZGg0OODMdPiPjmc4VIIesF7ydXwVyu4HzBOTNeD5xI6BlAcmNK/dxXIPRTjS3qPXzg
owOk+/bowlyavZ+OroOdLpHJh/TYDLz7Eu4jrpKEPCgdKqnsjc+IWjj1D0CNE2nJA5GHt8IzNTLX
fBiRn00VIzCn4pkri27ZEgT/t7vuW2KbHKdpWWw3506Wx31qAMzoM2C4plMzs4DAHP3c+ZTIbG9j
DLFMaymKk1oE90N25m3M9c/nyWE6xLcGrvE4eB2M4csEvrrUJZp3x1B4ZAzSWcnY73L2GiU8YdDU
zcTFZy3FRbjiRgZ1PzlfrnGh+v1sDKoWGZ3Iov7h5Rd5gfSLi4+xSefxN0Bxe6+hjg5AK7/ZUvWq
8FsIrMWEEE5LfTk8sjZpdz7TS/9S3qolR7poo4vwBO53EkzdjV5OglGp7zsXjCvuZts9T/U8kIS8
5QNPdBNkQLcNI2CDS4LTohhrZ21uuudVeKxk/tOgkKoZboGlxaxD/IC+Vmp7W2SrgVSpVEEp7q5j
zaC00rBKSDvK9VUm2AlCvTbrY/Cu5XcmdEIPVGCyfoQZSvMaODcHuuv8K9uDcztPuOgzRi2h4bwl
GtfvfiPEd7iCxT4r0k8qMdiLFl4M0QluJOEtq1pkzIHpHYeh9i+g5QkgDSXUAYEM+Y/GAdfbNyyD
u3JmWfKJylwSxDwhnDEVnQuWHnSYVpv33sBbg7ZWccfMujeAMf4uf8Lry4joYSPwmql9blZJBtd3
YZeKAsEC7tELoOflagDXPWxmx+wm+fZ7B//7dz9FX6eGF5efD3eZEk7VmDmOYEX0ZYzYbC0BPO4s
kSSieiQDHSDhi13dfO6nOzBP20G6jzGEVySLF5fFgfDnNlXrS1wkGLk9TYV13sxZNShQPfK2Ly4P
PAUXArWdtUSuEOhK5rgCG/7kamgjWn9eKzCKYf1tfLMQLFrIc8k9Nb/tSBlI5OLA4cSSUYVu6fj5
mvAsAawN8ry484j3AzTPa22Pt3P7v4AEvBPiIqqdIgjhs/QM8jPIy+J9T289cBTYKKtaz/A1zvCV
7hhUtxfyArqAwNmHCX0AU5+6T34LMc3LK9kNMaeTPIu0ihtKV5kFo9CIzfyXrGjfrZKwmbhP5X9m
S/ZjaYY2N/RLsxJY6yFofdMnFGyCmeXrpXjpgDEb7IfyCp1tnkv8JxqSD6/3JQ6NJQAFPci9LWb4
rwIO0a3fH5MX4GyiAysoCoxyu+0iba0MYgMoy5HKdsd4Oi92UqW0yZKh6Ua5oy9ewdH/U5pR0Fes
f/3FKtEqP8WIOjbeauq08EiZz1d7GFnQFZxknMV1sJN1RQVncdFakjLpPYTATEGbFCkNmyUeDfgR
a3K9Zmrt4tafKIepgvEsgIHEqeocgXJombypt/dtnP3+kyN8C/lWtSmuUGKONpaERk8zYWd06rG/
56/YZ68zewmotk9s1bw/bZ9b/VvmtHZmBp33x/1MUrmGUNEI8WPBunrq3AFssOcWMwibu4VNnsiZ
dLnl9ABDP4bkTNvMPJm8xAKKtHMnOLkOtH7dajfJ8XQOXH2/GSu5dKcAMDxVjyhOVvcRUkdoR5Pi
XsOFiUpDE8Nqk6d1Q41gNrIilZwlPlVy9bhMRYmtUkjjBR+znZdUI2TgTe+aSSstPhlEEcAvSeRI
hMrrgjgX5XdpMJgosKSw0hQZiXzwXqHWT9dUFuWhbBgvTcfJcF6zn10JPleFsXLFZEnaHyq4RfII
SPzbBsRb0UC/IPlSAvl8B8mrjN9zJ5BTb3kM8pe71JRvBR6+J6xHznrOTCYNSEFEucSyQqYH4ZF1
LfogdbhYpR1Ps7wuNxs0xwTgxU+J6kHCeexgORMjSit/t13jtTSNhQsV627gnc7Lr0/FN5+yySu+
ina4uEhcaA+uBaIdG4VD9MMFNI6AhFV9SY/IhVsVAY0/ynmzdpetjzW1cjHbBUbTzTRHsDXD/7aM
kk3FUyhCMtBh3XcjCarA84litKJqc+lGf/Ki3LvLwYzlM80NIofCeFctzF7HdFm4xEal06Bar3Ps
b2qApoDDklAJQDvs1W/7qiUcK1czp7TJg0vCKsBQW+yEYuGIBQzHqb/ZhhFnQqW5eaFwB5t9XNJ8
n+rFiqJOYF6FHwveFcuuH7SzB8h8TF1RnzodmK9Yz9TNYV4g/hPhTAb0p21l5q0XoulwLjR6uV3N
5UEOj9Mvo9zTuoQm7oYI/ldDn6xjeH0zKJlWDB/yJ/EcJ5DhKe5GzUzqlPYRG/yMl+SYxANW96S6
BIXoGt4zL+L5fn6kSfTjdfePaVnIpCO4gjF1g/yHUg763dExy23/4c5kN6NUx2ZU0HdEAIpgKrru
2mlWs9TcbChJH96kGFegCi4R1OLncl2QC+uAo8wN9xO1oa1XlWD6FNYd4wW9n7OfbrPJisyilXX3
8ubO2JSe6mFFVQKQy7CSV3YDcZ0cyZ49onqTJ5iVLSbL8bDllw4m4NGYXby2UyUT0p+fC3g8Qd00
RfO4lTbf9mYWQR6GiRed7MPJYeYuOYkhtPN/CM7+WBDGvadaP8Kuj/+aSZS2AfC/Q8SXywRBd4vr
TCSyY4vbunTdiHghuqEdEpKxoFfxuaBg5nK4uPwqCgj2ASSqhytiSwKKr9TUMScfTpywZ3vhauQR
mA6gYOGZnoz/tJa/Fh/B69VwZ0dRIyo2P2ai+QEvFEKgW3Ak/kooj7qHnBZl3/6JjmsT6T+LAmzW
dQ/VIDGKoWm8u/My2LC5bt9JYcXF8NSlEaB+oheznkcgwc5WcSugOpvzSU1ejBmB7Bn0qIwCKaAA
VG5I9okoo5wBKNl0EcE9uOiGTiFXAenPD+q2GH5Yt7TnJaMC3sbqDYyg4vNdXQ0F89u2UOO4UEEt
SXa+D6vB9okpGMxrglit0ZB1BLRGTK2eX1MH3W+q6oWr1xjxg31yaHZPv2FEOy8+VIFIyywaHfeC
uKTVNT6T0E1Ss09zNRctX4RTrP6FrayqLdDdFYjThLz7Hwg67sQTlK9TOc9O2pg7/FG9jFE8nx2k
GiPrK9gCvfMKzc3PAZAkjVIs3JsbjldQ5kBkFoamyMQwItrq4cP4Ex2fQiv9GfhinIJT2dvndHWv
iLNUeZ2R/EwwCnQcXCL6oWdHmr+NtgsocbBvEzKIfG3SkHz3nxW7JGgNxqJ+YZf8f8yCwT0Y4gd9
NHFmO7ZDwmkBtcKr9I6dvRqnXnr+d7W45Tjczxe/tsPedBOc5diPlWkKnJRpTTOfV0szw9TLSTDh
aFdJFoUERbd8FyWUMqcPEq4ra9RAdonsNWNk6dSiItOcyPITm+Qcrab6kB9jKwisLY+AlDJKLdFO
Jp9900G8MsIo8NKCPCrclw5N+y0dXjvaEKWwLuzI5GIh03xwqo8OQ/h6XxgjGlFkVB6iLJ2cxs9Q
obv9KhowX0MjyFHWq/EfjQsbtUfnPZRRU3xjT6zs+mUu5hmPIQ4m4AF4b2JupkGbfL3s7bBpnwCt
pd17gwbOcIk7su/k7VJMYCWTlAMJTex0v41TBSK2YdcfujZ7KZlO4/mZ00hlJPFzE83eJi0le5yd
ZMNO2oJZ+Gn6AzKMGgch8O0Z77fS9zFlu99ZC5qREPDcepfIzDp4k3TTWryRMUyaNoj4tTYxf3II
uh4Os0C/7RJTwwn4LqxCyytpMNPOgJlQKETQ3178GkNAiULrBCCOfGSrJQMJVHtLIyiqrWZGNZFi
nMJ5V2zn7/IX5E/llc3KV/G+XeAPK4XFFsyiIFoRJM2z7PgHTuRKtdEPVBWBfa8m84P/LU/8oMzh
YvOFZ50FClZ70Q1zmHITQwMPBLZpSxVkuiLN648S7weJy0sGHgsn4SsUf3W8AY7lPqYc0diNJxsH
HQmkfSZXztpBqlbgfQ/tKboLV1yucmBC+k/bEe1Cp4mlrBd0FHofYQsm6XeKuPFWu+LhB/YA6fp9
N3+Jo+/gTtQXI1UZKh1Oti9j5lFtQFT8y1kM28uyg5J65whxfkecF9tjO1rZwKyXQ8bP/8oFwNZa
ujAh4rPVBBH4+xuPgnfJ10vxgqbJ4Vo1lsi78cilQejzxdNMs8nFZ5f43469eFrrjtyW3BIda+1w
l8Xv+7meT+Lyxh0xz4YRSXw121UvmVaCKNU17jnMJvY634QcBQ3d7e3k3WWAOz2pOh2KOHBk+FZz
SeR5gMug+3yiOcV9GCx717X1D2uTBh5Qz6GzpoERVSvQMqTmrxQT9ae1NET4fcykPUkI2XP6ZymO
EgB2hp4/POi7hVXixMEygz9d6OFfAELmEgOatSM24TAIRMcJ5902V/Z5SUoX+q3bDkavWVs3DTR2
3EPLnjFjLeZdYCvpuzfFvcnprToQcZG/05seQXBNigHE9s99Kq8GoQh3MciTCuyY4vFmJ5o65g3P
YgkWYwckGa9+zbdy6+iA8dZs0E6w3cqAKB29HymyYSIeirc4prAKp9q4p3H3/RHVGYI+wB5Ct3IR
P+8lc9pNDzhgmJQHORMzWyknZTeCSSdhA/oGUqtmsIFNCJgQVPNt3a3LIrG3+0XKI1IeZowvFV0j
/c/sdkYZ5B1H2asX7GobPOV0Ti/UPLQBNMLtvA91DeWLKzE+UuQCbe9yc7Blbp7EHdERjZfhoyev
ihsgnTDmHtUjVB9HP+VBf52EM06/UVVp7SmE3A5Xwbs09+R2PKe8AT5UHrnrRMUSCNzH/955aGy+
pmUYy52SU+rckK94cn6ytl0udvOCubw/u6cUgrnAJBKKy9JR++mSXkmdJZZm456wi8f7dFydrTH4
zHR9f8Wr7UqFJYMGhcYHX82fErgGBp/cjHn8kLQQgBukpCDAUGbll3ADK+iuFy832o53LZk8e5fq
51dVEuWRd3pyMBL40pAyCfZt29jTE6SqkXaOdht7T/lPw/qPebwnswM3O++orvXJvXAijGXDbqKs
SJFGDgZ3E5okCo06PEPeJeCvw7aBj8U7JiVmFHi++TTWuUoeE9hxJl4UKHw9XIW8bDcjAs7L873N
QuH87O3XBg62B38v5s3pnZGDMaZDTnCD/DhKEy8BJ235c4KdlZ4eU996PmRRzqHM+GjqdDWOhPBp
tRGrXappEGAOsObTuWeMnwtg7FN/u1znFrSWu9KvfzoUdGF19E98o8SeYFobkOUDpOpaEEE4cYge
EzjVc8JaNyJAdxH1ZatjwO7fm+pq+0RxS4NMg8jOCvAuJSEzZLTrBHSc9EdClbvWBhPdblZz3XqW
WdpfktQqDcB5AAiN+xxDAGJQrnwbWwJWOxvPtyjH4y+tHJ6LCzelrvVncvavK0xqB9D22hljWQY1
XgIeZ75Lr6zsvQN34wPaDG3YrLAmyWhF+dEjOzrEB8iymCZNidQtfY4ef67pwQKM+dzFYPF80EeX
eUadhJLWrEIR2E26tk3aLhLgsXvokR2iCRzA5/ljknw2XrhOW/TMwAPB7YBSrSvLP19SFCpq6TBk
e38zCyeA2bFadElV7Ts1P11ZosQ0KMjbZrBqOWfGCd0YDyb4Ws/V6C8C6UjUPQVj72E1cgj9dNqV
JCAPluc9wir2OPGBZwgZ9DFoK2sZu2xSDb/ztAAaHh3rkrfzhayf4Fu0AO0fT0YjdFSL6xyi+7WE
qCeDyptbic9skUTk+lsN3uMaaBVM304iNARxJRDCAthBv3ixHfldpUGw55PuHfBh+82AsD/LYLfX
GRA6lDJLKcq+4kZlz5TJPM+1hhm3Dk6dhBVEi3MQon3IBVfPs9q67RPgUqgSPX1YBDUwOp1W/J9O
+yVqzUQWhQj6tfRNaxhhjbbxAZNj/b6AKtbgr3/8UgjFBf0+m9LzMUjsYSv3SwLmFbDUHBUfkziI
s3UVLXDRuXXj7IdsXVnvaZC+2e4SEtLDloA++kf2H2qklOMYAudDXRJBjbn1U0cB7wA/g2N/Hg0g
OeJTZZbU7D1vq1lArYlCy/kZ/Cq8hN0HmqgPX9LSumZQm3e3/txsFQyxfsPdHW6t2M6NFLf4eGnL
Fg4e6bogjgfLEqdZV0dLgXAO9WBf+6ldfgsfo80HnLRa99O60s/YaiM0UBvawG3QRBw4/vhrr+PD
J1PBWiqFy1PgDa+85gFLqR/pMjmijgm7XnwYtoS6xtvRaGeoIdiEHeme5e5mM14tp020qQokKkKv
Z+ISr6J1qWdp5T8j2fXyVaDku97/jK8uIIvk3U/cI4zCkjr909RsaXVliyQZ45kg4yXsqMj6s7tD
WWnA7Zl2W3cBLtdSlbe/8ArdH2ogz9Ugvqcj5GmHY7Aet/i0wx7EbRZQ3ed/mHJp2U9U6fNt+f+/
rNpH8gyawxfqfJnOlimK0oVMLdzK+hmnluq7PcaX1o4n7oH7s44cAcM+6ajQd+01pclGBY4y73CN
15czBSlKRmUwS3I+3PwT7VAUSFBigDXsBLlZbl1fPrAvYkvmCBhA4RCbR4O3HZZj1/i+cY/TBxSk
AUCE8SQrUZBF7g/nS7UGMOze36v1gaGbzLA4Hqs1cvdtSuPX+08KZOub18Hln/Qi+R09GoUQbcs+
/WFqacX2GCzaWKO+IRpDkmb7X6KBo7+hlEfOzMFa4v+YcHDCMH8ym4/mT3I3AvcSzo/48TsuIU5B
msj9ZyeLIt307yc8N26XOQqJZ9cTWg+srcR7m0kkPfILzn9mkD6IlA5oTfUZ8xFQXQLxmO/GNcOs
Ky7rqqEpx0SrEg9rcXF7nSTKQM5eTCHbAD0822dlVZ7K+mZwYwQC4teDKtvC9g2d4KVE7Lyv1eDb
pw1XM/N7wxtboZu3N0co0avbEsClWUPbIaiGoM5/AaFBycJPOGaoUdRwOKWG7retKemxfBzWEPyW
oINoj82gI9EUUFkC0M2sTpr1zs2tFKZabzJl9zWvJBsbdSE/ttjO0iQc62gN0iPdmDnR5kCqSPd2
YVgG8DpBveAlWf7Lqcf14wSj8M6SfBCanDY7k9Gq1Vzxu3vvh7c6lphevgKxrgKxWsKS1STlNvYU
DwogwEdyzsrqLCjo0zveGzcO1pfqg+XpccOxWE+aE1BwLQZR4Bq7WNITIAnPjg/zDkfM0b9mMtZO
cZZix+QYtZ/3xPvGnr3JtQbe+qOdbhIAw9vJpeBAD9OxLpWu+oztH72ioI+c+CsbMC4V4nzIL0UM
Zv0gRJO+7MnfL0rn70v0d6jQe0EFkXr6ZmcwULPg3CykaEe4wG+R5tcK0YA7Ng4NnoJd/StrV5/j
HdVbZke1EwJfaLIQyFL7YEGH8CnIoKeJm2KNSUzxbEXrMgDXuaqb2LxJ83KoaJ2paCihst0oDsSo
a7iu4rk/O0+J7omqPUoZPlG5OgHLG35lx7hJMBh9vfVudL/I3xfSSE2nFphdcMgYHnPMUWkZlfI0
TCTrMH7QMt17yir68hPGN2WaqFwxK4q9CkTbuBnmAyt3XXoJuNMcYP9NLd8dz1OXEK/4W+HhjCdA
y5ApnX8yC6Yq4s5TJNLFx7LCwqIzzVZbDRgZ5nCS088heG0FIsN/7i/f1kMr5Xl9r+1ZgmpEXnQm
KNgXCRN/PQmIcl8Gdia1bcxmKPhRDnKExp3fospuYZAjNnU5PsIukZK17/JBf+Wa5e5YqSOlhMxY
oy7gSQe1wOXKW7Wxut0keSnqk4y3GDSw6kIjTYrA3FS5ooC3LGC2RSaZK6Dg8vZR0JiX9YtDk+29
EGYBk1SpRLyQivH42SJQYqlHD95s6SfHnwdvPnhumAWTYpEkC0BYkvmmWu1aLz4fkJ0+q0crjZiz
GSR1M1OOwPi+VpxXMKmLhwWnOXC4YcNn/4YiyczPnIee73yecvlmBsn3IGL6TGRqZG65GcmnMLUR
CPDHOBT4Z+NCe/YgOdt+9G6GFihx2wsPGjef03TcySgm/sgnmB/FdYEJU3McjjUYSbtqePduLL95
QyIdb0BEdBaa/PffgMLbVpK3LLXUrjpsO+bTzzEygcG8WMMhe6R2P8vHIFwQDW8CFDMutzZi3VXB
21yWtlM/gWvwbiSwTqnnbYV0pbEk3dmLxgNu1YbYB7Su5c1U0wKCPup5Sr3mYKnY1z6ylOMfwiIM
EB5snrqKCCG2+XXIjiRduIHUDCKI/jGCzgNXxZjY4Pgrjb7buctFgPasjJd8QaZA8E5ylQKAZJHF
H67+15ArwBZJ6r4FH59YD9XPixBSs2uwdXFjZge0SbzcZfAJFx1xh1gesgCOy9zaT7J2JdlrfwlP
he5103+a4tuJYHdbR2izy78et6ZPoeIv/65RlPPcHqCnFLlRGb6vhtklCs9w/sdxajQoMNgi89/G
/RZXtQvTPYYXBIO9V7c/UU9QSZWz9qbYRVs+ZLl6iiXY1Ro8G5nJCz9Yo2pdW5W7UKGu8dMtZJHn
ZMGE4G8dvpZZHX1bpglb3UWhKMd7zVp9I2r38VK2BXbLGjubGRunpypF0AYiBh4B4dTB4g1924XN
4PlCNOKcR70kbBCVoHum9osc7v/NvGYmBquqtkPLrN6oMTMVkgtB+8cNMJY2ndjufhK8dUHvQBWM
VjSKni+PgRGmFRnZGq/cmtfURBeSE/o4QNJfuyCH1EnvW2mHagL8WNmPurANojnH+mSMjBXn8Hs4
lJQqlH5ykx+oeuXQQR7y37H9s2yZ3hJnJSLyPBFQY783Wu1gu7RekFYul3DvBwKBlR6/Q3EZ9Zyu
nMeOul3DBCKZEU1KUaIte+GXgSPbI7G7TOgyuWItOma/IJM20qVSJCqUgBmEGAMu91Abg1+c9Id9
mm9Bd+LdW6oiGy+uTSH/+c1DCYxAloGrbJS80FMgBz8Jp38NcU8dk8kFOXcItdlR3xKryoug14Y5
8RBIu1u3Q9L5cydQt/mWbEz8z5exMy+td/gwBMPkCpf7h88990cZx9KVuALbhV/X/eyLJyEY4ic9
wg+QgF478aQXZ4eKk+F2IvZ5fcEN6KjhNF3dJy4dSVpnf74M+xCzjUWAE+g4nm35HbJtmxOSUJwy
FhcT7INly0WT+1XiWAqcClnwwil/yV5qoLbk7kdm/G50jjZFRKimnYddruTwHt6tcQYG5q3B0TZU
52ioKtGgdV3LMmam7UwIqQD0F0F3FCaSzLHCghbKMieM1x7UpZL83t4oSUaf1vkJSsjEY8VcQehq
Dxs2H/QvLXNBye7NE+Po1hkZ5K+1P1gaksrxBNIVeSj1cVccHN6jlCSzpnBeqXRdqO708VrF/mjg
VZVd0Xxo08PI6zn+2GoJrDK3qnWv7DfW4VJjndIsv1Z8afamItOuunfbn7ww5rCkd76a0FjXfmwx
Jj4DO0vlTc4wwhWSiK58zAzhBCf3SWRZPIzf67l6kN8R3smeoKE0lbfW26UqHEvgdtXdno/Vh2Nx
L3vNPKgDV8mT2G4juta6CQlzJ/cQj0E+fOLPvzTbnMJakgs46DDjOByMaeLCPV8+wBq+lUIDALeb
+s7e4d1HWD3/XTACR6KHOlODVwINbFVheyIhTLFmpE9dTNWBSjur9Qz+ii+ZEtlPlJbWvPBsnVnd
v5amCMAFejOyxciZL/o+943oRGNxbqB8n/PAbYkSMZwGHwrOtlzx53LrP/jyUUCMS+ddMJe35bCH
4SIgeGzQnXZBnhygDLvpE9xDo8ozV4ATnzU7lDidlpd5p4l9lnSUc/HjCQdZEVVXYdMMs0MUei+A
EidFzZfz+XaM15MMORRdJgpvB5OTsgJKbUq/poG+5Lv8cSfnI90f6/yiZBU4fXVCwVl6lZbzoUty
28yt8qRH8zJ5Ma+ZAnKJcjNVPQwBo/Mww82M62n1uM3O4TF2ZGmG4mlg3jAqAj9Zhw+AOA1KE137
YLE6Sms+qqpW5k/8dJO1McjlhfVxEDkosfeZg/KxrKnaEwgWFFn3GZCFpJ7BCKIrfFUJ+sssA/Nd
We7hPjaASzW0l7gJiqOHb2DAB3zEyYwooachTTB2eKnOT4VoUVA9cry0qYbJmY8RvEzWFA1x+t9v
BaB1all3gE7CCRHYyzALTPM5q9aGDVKJ0UQNlzFyhjJZFAhr8pItZ+XfuFCfY+eywoFsGxT7l6vK
vgThqZyZTpCHDUfQpe1L867yM4F0+Rix4xskGiyG99BDY9UkBK3qwrJPrWvf4cc3MqMXgz03midj
1tYnltrsnvpfBZIya5oFneuDVCBL1CM0fW/kxeWNOPhuBoEgBdVSHDLF8yy88s5A+VkAeJq54gQp
BbVjSHFwxUM67w7Y0wrNIq5oCD3X/n0LU7mb2WMy5ndxCyqh6rpdjChTMAvxybmExZa6E8szeu2C
mlQYytZ/+2C64cChpit+C8PdHT+iz3Sm97MSSytNX4FyNyVt6fxDMv4Uv2WnBdUa8dRpWfBAr8wb
hrytKYWyJFEYmLFrYtC6nsP2/LK2A53fDYJN38Z4gDPCGbF8qwwZEkVbtsCpmYzG5EUijGJL2Gya
yY8cGZRkgcDo9jEOEZZdMtA1o/1l+h+YkmKZ4OGZ5/8pqpFANFQo27shcZTt7xQG+rrX2KUk4UUm
CX3sVCOTldGtLPR/ER22O12P+2iZBQmxWYIlE8cWg2VQkSPWlK5y5UdUDi918I45rz1HnncejmVZ
w5HgLzcuH7a12YM6qm1O5h9E03IUMc6btGhqwdv/X+zlT8X6wZay6FZQM/BqW+zJqPTo7/pRyL26
4f61Eqv0YqRdjmAEsof3wAzluhFhhdy1iUhzhro9vRvhUa4lcw6JVThXkMVI0z3I4v/HUVKL2luV
jIzcG0eGK0ag/ffhw1a2mOemrOr2PyyOFnIqIExDVDhu7zfLUlROBxoZ67NoWdnyvYPPPMw4b/eM
efCosgMMBHP+FR3VdxfFUH6Ett7Ax+HoGB3bqpIw1Id+9m9x8bxYLXWh8kmGRd2ce02XLvUIt+aP
dSFW16WNR/K8tR55Uf2RowQfs6DL9twya8aOZV4shn0zo/8Zx5sAH2DQ3Eum6hgt6f3jZMm/WYVp
kGY2EDt1GIa2TJVbL3u9TSkbCVw6/jHZzu1gv+/aRuf60YOiy8lAydC+3Cjx/bSENm6x8w8xzLN3
ln8tck4uYeGa5KPPoYZFcHZF1U15rlgTsKxn4zd2IPxtqG++HeU7dn7TLp8Y3F0z3KFgPbjhOwkp
XEmolZa2sxYeLOy4N+3Sg3sGPU6nHhpbdXd7+JwrZzVUSZ/p7ejKpSoQbxAhYPRCzPUgyYNFr+Hm
wYxGRX1meSU+BFfO+jOGfsqMFHHRFygsbbAbYKPYq+uMsr2b1hDdExhPwtnxD6bhZyVPs5Z1FFXi
BV/y7mBsgzuG67OH0gq4xBHXsmhhx3MK94jCLnUNdrDwgrVVZfcl9mMB0iXXzI+jBsWHdlfnbALX
EEqEkOaFnABQ6SL0a2bi+7MGm6E/ZhLzouXgP8z8SdN5xQK1Xdh1N9BAzcsghwBCKVgobMjMNc2J
NpJMf0DE4vsfBpG9o46jyNSJptOYHmeD7iOnuat6e8ljxltdhgED3j+NDgQNiKNXmrJBancdFYgP
SIb46/imvpY5EoG6f6KkLvOURC+WUKYdkeRu1cJshPVm00pmYSc66mBS2EggAqHjxO2HPa51fwr9
pU849GaR8aNZFF8UJrAYjm05TYaJU3iIQqKHV6OlGS3VQ1W2tE/Aeltd0czC8BiIJPor5PRXe3Cp
u7HXFlEleo3ttyzhPkn1uV/bB+aoYg+oS0nJxucOFdfaDNdyE/nYr1olP9T5MuSsskcKiVNQNLoR
74Do4xkhmVXVsAsya5vvKmNe+EslfRohU8AaiJoka4ks2s+FXAorUjx3i0cqzE3zhkXx8uSpSv8h
hFlqyuMWU9Wg3MsWBuQq1H3wAG7SzSJ84J4qbdd++RYLlsN9upTwATyEejV7qYyUuvq6TK5w4c2v
RjdqxyYG/SJSRG3ID1fK18+FEPSwZNRiFaoxEEIn+NLvvJxpexMGtwXsUYZ8ERF7TWk4Jb/dYnta
sADTHCJq5P+F9GBoBFxLRiu8FeYdHgIVJ0GGGLeS0HtYuaLPclIbZLRdL5TTu60nNBdS/Zsr9qQs
NNIh/Ap7tKX/2Lb8hLmrSA/ojb1aeA2uzJWexzIIZwAsXTlALHTywtoxlYPJIbL5tvjJpZGppolz
Il4Ut7UeO1TnwUyY9Gx40zYazq3CcsrK6LG5UbcTF5jjz27Fk3mnMbY3pY1O2MVpqPvvV7hiKNHu
zkpWGnNR0qB+WFeaOXeWEb7tCS+Yk1X68XoGDyY47aX1haYjFzEn4Zd1CJCJEnRkrFFyAgnILOcw
lfaQFEYXEiNNWXT/a6fADbuJzQxSs/X53DMELFXMlv0Pja3WzIstX8yDvfdDbEK1AOujP1enViwY
YoDrg96W8M3eNzpY5c2GBT5wxcojzgDvnEBhl6N7E+A+wqVOSSaF83gmt/0kKK4QlgFXKsc/G0on
z3V8eHwn+r6pyAOCguNBVjtUH2cI44gQgBggvj/K3QOVziC+jpFn5jOPXqIAMisVRzJ+1o32UsGX
nWG05nnfN8qZJeEAHAXT3F52ytKFyxXNJh6qPh4=
`protect end_protected
