-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
OnKLAoAXFMGfFR11OEARw5ajVHidgDfEq8V6g5kl8Bs3Z94zK24IGXewo+gIEDcT
f86E9R8CswnqNxU7MrH2S0YGg0M+exkh1bHKQNxsf0aKpeNvsuarECpSNmmWTepD
+K3af5pJkZS7U4dIpCTZ34tY9u8v/fea5lFXd5cuxyE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 121943)

`protect DATA_BLOCK
jCIX+BCJ1GCNs+XHlYMisO03UCSyNjwK1Tj2AF3mo5/hfldHfGIyVcfVDheuOzwH
mPj9J3fFVeIo9CdE46YAbkWM/nEbwsSsSBY9Nsw/XiIxV5OAfX9dRzVawTRmluyh
KFpxkuAf6O+wgdiYR8AMYD3tbcvf9u9jMFcoOe4EpXk/aUNS4hhW27L5WNR4a3hy
9NEWy1BjyKFQwrjQXmANWgjrZF3/EpRfWAFjd1PeO8O2l+B08xOENYuvlkuCv8R5
GCyKxgDoPMJgJ9JAkvRQSok3FbgtNtz75Y36jEsuf7Sirao1TH3CEBpUHaeEBHVK
TXlpwQ0gfjRTCpAxRmUjh0VAFbrSELwBtrHfkysRfNliRP9ZvdB/rJ769RI+CDAL
AVd66UDl2Y6qFD6ssEEH0Cc3CD2Q17z5ucuhnfyAgdd0bIv+cqe+oeRMZWJenHbX
aGtrh9buWGpbUkDbxb4kzWo1QKw4PsIrlMApEgMzpkKvsrAYkqyi/8MJiNkCS3JK
LEqcQl0xda8xyjwB1baLsjWAsL+SXSUzQ4/WciyyVjgEF1NKMC5JifeaRRIst4EQ
bFh0VzxTajGc5+LRXgCbJFozRGlcqA+prfl4ubCqQMFIQoGMMcn5Pvnb6oNgQPhJ
fsXb8XI6SYecOH8KfM9lQX5B8ZxjwEl0IpSJvt+1KwWbjtCyjmnJKilxNrrn4kL6
QkxS2ByY+2q3hcToXFLHfROgRPkzNRCvzB5KZPx+Dzl2SlAgo+chn0frnoO3Bj++
Av8ASAMrBQYzAVPrTcyytCQEuwPvd429mv1coBzBel2uyrgL7ZXCNMmweSN45U6f
Lul3dnl2VJHzJmuA/WX4NZO1FS+Tel9J9w1d1Q2tCJVJ5KajVRYfo8xw8mjdldqA
3NmV0y6yV/yoHbP/dLuExt0Fq5oPL2+FfMR4cJr1P87slAvtMZbOoYLavpadauWs
Nsslg+gXH/iPmyZAOOuFSRx4Z5qUb0M9j60IsAh5yDVWb8FTCXxqmRrZ9Oq4TR/8
o5PAxnSeCzSlF+Moa+5TUdhH0MRRBeulvppCa83DagKMvvIkbiOBWgkegxw+Qsu0
GiL1j2Q0SyrtpcDPiA2rzlg/Vv9nCmD0QV9+gkllSj5yj4HF2aGcIpB72pC1N20h
mgcX+As4RGRZ7KCiQZd6WhOxH6gpMrTZ93OhqD8/QWezRibKDR9NOsiqNEQso+KJ
gilGEWVQdfInUJ7xRLszl6FeA/vRFGSC6jbbqm4o21pB2KYfYbZi+IrSTeTxzh3E
vPJHZ2X3lMsuopINcfwJHr1YdmmI6jm1e4awH8O7nSwX4KssjMiV1gJfXnv1KxTm
vwHicOeDVlKKzJ5beRrmMA2JQwjGMQ9/kBOt7hReeDyuDBhVTEvHncunezcPf1cj
M4cHL3kDcla7lVeq2cYC3qyAzVJxLH6U1Mle0B9EalNxt5EE97+4BObD3EpGWj9Z
kLBE6bQziEE0ZCbEytPGD2t0T8D70WqgNaGzjf0XYEFrXyMCge47iRK5FFY4crnc
kna3MIrBjV5GCTujLdv/WXSXjbQRUWFdTnI6HuwjUeum5SIGa3guiYC9R/DRaD1r
5hxxPGRoViFJJ4G109d/UBJq7wS7Wn0NSs7HDhcWLXYfKruCHY/wZ+BGMk5dkoFt
zqWeXzS/httQ2R7viOON/5M/uODgZX08wgWr+LYbjiy2Z9Nm8ZTU9FQwHiD0CIw3
fuQibDhjuOxCUSUzyfyoixz/tuvVEl+CnmJl06GYpFrJorE73LbpUAA7Z9mOBEUa
tHYyx5qJsYC3LNNTr0CZt21yxJIbdyT5coaseHJD89F0mES75DR3+fH7T6pZkhPQ
6EJv7ZhGBDoaaJN74zhIhGQ6cabIKt9bsfy8DmdNT+XOM8/p7LkBTTO6uohkrbm7
eJ+MN7tcwUJQhxw/A5nPRO5s9pO3DYU2IEs8zvjPstFgO9E8+wxayyWPUrbix76y
iU1RySIXCl+sWc4Uah04B73YvEqQ2dV6W1ES6r7ISgAkxoc3DGnzcxd61AU+eddb
818XYgLO4WDT71gHIr20KNK5JX3NdxVosGeNICSHy2SiMbqHUlEBn2hwqmgUalzO
xpFspu7w23Ukl5l75FZqQ7wqGA2ux24FDsE+ki8vGDxeM0ZpBylwp2ThBbvGhOuD
WqCeVe4hGXLbr1ccvc6RZw5BET39zU5iSjbA8nxEc3ZXOgKpy4EkWpRyhW8rUuKv
4SjJmqPmpWZRR8/eLkP8TLLuo6dxB7ASQmYpbRS6YwFKqdVU10JkVoIDO2b8T+dx
i44gTVuehSggnyyr3naeq+hehUlti4CO67nYTfFDM/5AkHa6dBl0cTs0c//VKq42
yz/0q4XR+CvryEu3gDLWLU4XuQHnvkEqB5/ZDpHUk1/zjdTXtQUVXo1vXOhnw2q+
zSMZd3At3qXiGhjm9kPs65BC7Z1aN+PnF4DwdtNu/b0h5s/eYPxsZ5GItaf3tIop
J4nvSXnVwtFX7NMTtSTXJTtcH3IPqWovZTq7KB2dFfRlLcWB2f9VVPScBnMoPzer
LUoeLCY8mqI+iDNFyDsqSb0kaDpfQ1QJWuUfMWHkSy4eeQ0+mbqGAMoTheC80S3L
4KpHZYI5qyL6qFigrqk7w/gdvmht/4eHnCNc0jMIwfIj/LiDgCpESdySBTpX+Kqx
zEboJOByf/V8Sh5QieyIOmfFJDcxVs1GaO+vGHfAkIqkpOZKu7UL5DSC9lPZFfCr
2KPBwQuV8F2B9SwUOQ+mZD0ilOsuA/sndcbi9v1ws9YLyRf6NWf4xwmjxQqTi4GW
gH86+rvAG8VJeQoHWExXPiizu+Y3adSQAyrTOv8xoBC7DJJabqZXvhfq5HJmHPL1
tORC2lruPULaGg2XK9/hMXi3WZhfkasSkDzAFUAqqgd3Xs43VxNSD8/yu2AuMInp
H46R0bpRCshWGLuWYKCrnb43mV5OYXklEFWUYviCTvJ6UkY3Aay8IEh7QCQbLT4l
/+nc7vkDkJdiatf0wZ0hM1tSaYWvsRuUK4mJ7IeG6ZH4vX3n1TyEH0Ob5AKnY/tn
L61ZG6b5vXJLSZEfSD2Z9Q96ainXNEv8XfX37KtNOnzLsPEIZDKQZzkTr6AoV+zq
ufbADAesEcgJYSLGdP2AQXod632PjIIDe8FQMIp+RhQ2fvYmAz2FHyMuxZfIyihX
F/xiV0oUvD4mTHsjQOOWSPBVU8wyxLU3JAdiWz0ulrLfsCvod7lY4SEoGL+UGMip
IJd3qz+kPdThj81sq9nqN/WBq3RGL5LxvaGJc4wHiQSV8Hw8mR/PEveuKOLk4+qv
jFQpcTcQyHjlN8HxDzPskpxgQh9Soo5C8h2Ib1vJzGS6At4i0SeewGaH9/9IdWEQ
8Y77NnXjrNNQdGwyqYGSlmwFnL2JRIwbkzSazQvg6pf+PFZziPzwLCDOwsgwR9vf
zNOolHzaAVzclCLvf9JPzb00CZbqw8kFfUkT6lx7DpXlmnM6vPcBfbXtrfX95NYO
2eajSwRopGGyDSAsEa6YKWh5AlkknDVVPej1tS7My03IWyY67b9krtoJuR8OYeVk
mLKtrF28IJyD+zqCFMYtVQIr3ACqVqEOHhECbdlTFDX00ZcbJu3NlUiTsUz8uJzg
ydPI+54EuTg2AF2aMxpztvtkQ/4kRqIvzfs1ZtpZYEmO8cxH4hwZApCjFhdH8TFT
edqRJ2T15Bt+QMZYSEdbtzr/KV86fX8ZyNjxAerly5jqeK/vKrM7/ukVym/BuhJU
pLI9H8Xuvj1zywCtkUXk06FwFBKhV4PFnEFh3ySlkHaZbVW7yaU1DuUR/zNAqRKd
IupVziGTq+cXARHOHvy7vDasGvQqaDd5boeKumBDPk0ya0DZOnG3TRPQZ8WJOIsj
atqY/EyZhBqe/iFsiNHvHvjDuH+gwRIrMz8AGf4aEbFdmQqvGC90Zi6fLIW/aqEM
fugU+07oJ8Q/snivdYuDPvLF/1y18CNIAkwaYz0NR02gxOQUs4Nvn+ULo1Z4QZjJ
JZZbRX3dmUF6zybDGYUJH1evJufc7oqxrguAmUCuv6/N/ahozTk9rCbrlFLzESHt
WjzP8YO0TNDv6sfaHh7xz213hP46zIjz4riL0mXWvN/sx171BjjzAxPFpQV+/Dfa
Rhi954bygh2KhwrMbSZMTlZpSPref2sygo3Iak1djjMcERiYIAHVJ6xQEH9uxHM8
CT7wOaNo+X6WviEKomBzyQDGxGiNVUshH7+uwZu6HstW7r8h9Fq1a72w7mWj7Hkn
/LRHqmjiK+d/T8G7FI0DHdB8NIh7N6Gr7sDektPhNJPWSDXXQb3/vEoOAxfW2LsT
EKGCLQe43zmVKKtEfGzM5f/p2x3SwFvE0HY9m/A3q2MjbwjikKOyNndVky0Qjaqk
H8rwOLwpCCn/9XPumyQ2xRsYIiWnYvgJLltl84POJyj+A+cznHLBQU09a7ACjqCh
TEKKCMd5913dhOPy8nTsN5IBZYxylA5pmlp4V2rxZmxuZvo2TElFB5W5WYdcWQA1
zTz1DOEyS6h9hjquyJ7RfxeB+DfMExB9K1g5lpJ6qV74rKIePVgfKUsC0S4b9fCD
rYig4laKeoCuf6JQLEDLCctNt7Z5yo2nKxoU+bz+IjMX/f7m+yHxC1hZcKQkm4Lp
Am9Zt1ZIfziYD1acF6N3Dx8jeiLMMK5Z96xLSdE+MZlJe2pZ5n/7PXghlxcr9E9A
2BOmLBwyk9RKHr7L3ulpdh0zi1uIrf9O5XLxQdtp7jJDkIhlxWIQ2IS3h6BFNais
ukUR5KovLN8g1ydUG4U4xGmJeDCMpB1QV8L2GAh9flq1wXKanQSVcC8ASySbABKs
/+E2QSrpYmoADY+4U0v2n41cL7Ti1faeU/jHj/bKJdVIckKfG5ZFj7JDq/FX7jpB
vq+sm1GfUo7E+It+lhIO/PRUmeigX931qfxXmrvYR4wRyI1yNEff8OLfpWKV/H2l
+YaVsllZP10+HgSAbfqWHmUsz5MjG4IbFT0MgOS3pC0FFG1aMm5iiEjp63f+f0HC
f2Ao4F0sOkHnnumsZVNGizvBkeqkNrq+6JjUFq7wdWWJt1+p0ot7OxG2kBvK7JQQ
C3Ql46Ce1L8KDfJO8EJeY17hoKIHhpGb2qzjDlGtUXWDxTJVV7IZO58RDsq+zdmr
AwjsemvJb8kIG9cWwbGeUbK5WslNUzeauGq8rLU4hPOYH6F2HIzbYUCZleukXN27
tHCLDuwPSCoxYiQAdu9yabiEY7F4srgiou/fDpgDz2tT1oUFfznYAUHJhhOOiqEe
W3rh9S+mJJQbuQ8f1kQs7uIzLHEi8bOBaWyGIf2iEdHMM5fTtF+xJzg0nGDH0IMN
/dLO94MwLoi+zVCfjO8k04OI6N1HCQ4775Zbig1ltRXiv0iP8NXbEKwcXhyjwNVi
akM33xr9ocakn2bwU9pRLqwrteWq52w43MKsNpEm6oNQFoUzidVEBJWWqeq8t86i
uxRuhEjpbQVL5Wyr6kKySJh+6F7nGOnYPTvrg7IZqzeNfiM703ODtmjpGWKa+GYK
c7DonSxTVWzOrWmauDXWrYEUuGwaewEkQh+KeH74nlufmIHOKC9jAktkCNf1JJxj
ZsRQF6J88HUkNb3JnzrE2sslxvNvr6MmsMY+Mo3bnJxRcYgz6Ex4YSGZ403IHfwn
gFlHEi/RO1GB62dD8FuaIRPD1L7zQUjXpYmvVEI9AXFGLWSB+wiJw3TbD0AF728x
CoZwI4BntZrACoy7MQ8eTakEPVwljm+k4DpCXkXBkhupKdA+qaRIx0lt24bhPUc/
GufVA6d49KRaRbmMIubuhF0ejLmStBNRnViumlgKcTfAMHPUsdWsaUnZe4BUBYrN
Y+aXzg0lYmP1ZqPi+vCuN2KhfZJN0j5Bw0TEEGc+Bv0qZMFD+4wNsy+DJd0EmQyH
86jzD8SyVEJzWhEX98524C1gotA+2R3eIN7E8r0X3cxaybbgSJZu/cOfMilZ0zs0
GQ6PTLv6LghLbfdiQyPHtS5EXhyrnPlHPuEOZKeqtPsN00DPfwfMC7BAGY3CHo0D
NEk8UyTXO0VlPXpfgISa7D8dobdlEtKx3twOeYavd+Qc5Hgd27PDAyszkyvJIfjd
L2kl2RDDrcdUfHVadTLJPtKfBfGAfmYsMZgVB3D6deUefJOGeVkiBCOHstFx+WJ+
Zni2xrA9dExKsOGrOF+qqyjiu/fowbi0zUpKJ9Qh3G2XM81qvk9P9ULBQUWDdg/x
s4mEcQ9V+7taXaPo7PHAq17jeCCibedFHmXAkeqY3FGPNZqwqQInltf91UjUr4v/
C8sshWYn/hosbvNcprDOrpzUGbDTSBGOupN0L2S/u/KSf6rtYdUHvhc/+4kifYVf
1zL05eG7Lk4wn3hEpcSH2B0PjH+yZN/FowZiNoBUrcRwz8f8uQtOQW64Y4JGcXad
iAsDV5QjbSIVK6mUJjwqX1scxGlPIBBreuFvlc68/nDgNc1O1/62mdsuR4+mEEcM
pWpw+j+D8attGk/GsmjceUgt+qD+AmWeNiru4InuJGTZAqs0Tean1yNLLXScatrr
TCOXEo4IDUQHULz1hbrojidjf8F3vAdC87xpRSAfbmu/1rXWdTOEd9AmqWGY/OXp
DL/GIwWwy7xrOmTkU7JtckJ6Ekp9ONlAn5OhHhG9OCF+n0sLO2pQthaW21NMpCV8
1zaudeRT7vyTH+PfLR1dugGAsNBgSSnLzbn6WA5uAEFtRu0/FUcIux0ySgzpZPKT
qRlPVkgit8vGVKiVhki//8xUymxPunYhscRVA+wJHmLcZmG70NcuB6suyzE/v7Fy
oEuNwI4h1k0pn9QUqQBt29dpd9oJVPaiK1jM1kwut7m6L937Lcnd7eltfUr7aMKS
g78X0oPS7/0gAx7UC4+Q5b+44+50NPPj8R5xG73pVd4/ONkfI1tPGyHaGIC3fgKh
ktuxDraYszPmH4yh8Jg5XGIKpnGFhr8eSwWkEW7nHxpgUpqbNkn7hEJY3NYtVJ06
moxSY2ZoxHvXbKh3eOBdMy5gaJvj/L/nHTfSXyIhcetIONhiuHDh0pSny/IpDNUo
ME/q02J6R8PJLG3fQptiAN8ErmTJ6BSBvEIVHl9t6QnNyfcVucKNGZ7ilvV8JnpI
hW9oLmcQfEfqziOelBaHZOzn3T/4Tmunz1wdKX0/x8jpNshfGUgwBaY/a5Bvywpr
DIR7K97NufFH1BF2hXRYCoTqnWzdBlZ7blnME6IO6jdCkN9SwRXE7BwP5gyedpj4
kMpa/tQOlvdf1NSkVdV6P2M5DS4i3W+viUj9qUIWDXwAA6qwC+V8n+vhzSHOk6FV
73ErLI/lA7aBTB0BgJNlMvfC8NOlQ2dyTfT3jgsC4M2Y7RqaGJxCsqWlS/+jrYGB
aq3iQxPq0iIIBkTkALkadtSM9GUPGz0CiXGzEhkcHOkk0yK323rcYv3dO8f4/9IH
UGUon777d5nhua6PZF/eLHqEF/NAcGmD5SBL5BPjMIHaRuXclgvg9W2wHupqAsNP
lNKfizCTAmZWX/kPbJkuVjSnI2tPuh84MxghBipBwaUbtRdK+rqycYquSeGuIAQ1
nN/Jj4zloj+eJdOx+i4ge7nNwa5NZ8h7xwV2AYMVr6QYcvO+NZKx+b9ILYskNoUe
fKZ8QIqfkuTGuICbIwtnXX2TwIGkw1rShTohroNwsJL2L1h1PUd+hiHHogd/WTCQ
tunCemeD7N9+JQjaInxb0ROusswYlEjgsOYvY/oGLMerjbYBGfEwOPKNwpty1NiC
2pBqDWEgUwTqmENfdJn2gcw4pdYLrEZvNOiqhEygqp+2TZ58cpMCKLGuZyvgMDit
KqFyIo3PrcKPWHmlv4J8oN0rauLl5I743uA2EtG2LAY83RoCk5OHzW7oZM2nYv3s
ocJfmz9xf/HHFTH+O7HxD5e6VKu1xN62JOIfh/gNrErjIff8c0ZTDAojinQhj1Tm
/uJQpstYn/6R2X63MTet6uDe6RfT02s9nL8HwEqqrYnpOqUMmpDqiSzAaZQUpVhS
catqwVCOeD4IqIh+Od1J0ULnZJRcMY+tQ1jm+kHlvgJ0x7CG/3W73cmjHGaOdmhU
/xpaKnGRL1Z3MeZVkeLFbcbUPgJVAQLZ9NBgOvUjh93ma4Iv5oqm3M/Vz9E57Jkj
htV49uNCSa5m3hf1ry3I655scMnz5Xl7wOZTXsMNwZnEbK/nEdv9b/ZMs+16W/MQ
9fBXbik2ehW4bK/wnCw/4i8JFLZeTMDRRzIHDFzUq5wTuyBLXtLmB1glvOZ2NIKe
ZMQ6BFC0oeYRPg8p7Xf7QvOKgVklGA9LiedJCDXreFF+ghacTz/ZmXbQL3YEHpPy
LRn3ODZWefkmMbxPKfCYaewHNcHkUU9eO0X7sWoWbLhV/xjyG6TDbkHsPTZknkKx
4E4MR1RtR5rkOnALKg7aKYsM8BwvBd8ebthH0phOwysHU1LxDpXqSHh/SHujT+CY
njoTCkdwAeWqKYLAF8ZNqDQQkBIeLo+Pyh0aHxe5u5P4XyjGOfwpan+yGxhG7jE3
J6jhLIGIoWql3aVDOW50HDeAdkkL9uRF50W9+3cKx6paA2vM4pY4TIaonJLjP1tv
KVZqWpprgHduk4JDqsoktoaKA0VIYA8MXK39z2mzCAZlxfDjz8t4dM969HTM0Eia
g+Eo95mbaH7ruPGZPto29yZPC9OrHXWUwxE6ds7sAtHysFjIKI/ojOjaIOzuLa9/
ZnzjbwNM/Kddb6h6q4uMNCqfF2MCL4UUmYIV1YSli+UcUziP+28+u0nYVQRYGj9b
d1+4YdDX3COFpF2o9C2d8wvSrCj66JeIjyj2UmhHQ2lOSePtTieOmxDGX0PKlW84
7wH1Cm4tMPDtFb+QVb1QM9YU9LI3GHHd4AjjUGh62N29a6enszHNECThQw/o4Jd/
DBmuIZ6PJy7KV62DU6FTARr6xCIK5O44aWH8pD9vt2Fg/0UiNsjOo/F2SQOPFFcz
9viUItOTUvxAfqFQhpHJdSwMIkrxe0BAdwUuDdTIqGVEJE+y0uLTqz840U9ds0va
P6/X8dellF8yRf54Evu5D2f/H8k22feEE8DaAci37wPij5+7x5gJpMVfrW96Bdcn
SBxu0NMDMvF/oGoHelzK73APTvFsDRH1WBT2xF/I/iwyox6hQU1OjJlxObqh646r
jUvlnMxf3DUvz08lRio+hp4mKzg47nKmj730UpZm2c0cLDPzovFNYySroaVMH8iV
EFcndf0ZM26PthR+9BSm4HizEcm4wRDOwrXt9Pk/kUlQfo1tmkduS+Gy9NNAUMqi
9GICiQaCIMBlTnbEQ37mSCbN/THfuFpY0SygkRMSnK9T5BkyLbwJEJy8S7jcfZV+
JV5Rcq3dKihrmH/2sFWG8F+JqRdwwm+X3cUr+TdnuegiVf9jQdm/djTtV79VJdql
uZjSAisuRk0WrNDJ2fZ14CL/kh0bJUsAvycD641/erSBu1FllfNu0pnrG6zTSXnN
JUWetAh+Z1bQP1RGcW953fqe9M8NJEVUV7r32ehTHOBte+QwthZ4KKA2WQ9JNNBg
obQoSdjbefX12n5CEkbDSAXeYSYTNegqSE4CywfHBajascI62/760dneBgxemphj
XxpzmLJ4KI7qsF/dgfx7W6+NTL/Tz/IXH9FVids4utFmsOAJus2jN81ls5c0gdeK
VASeRTIIR6TJtd0hZFGGf9ptyzNJlYrNsqMU2Z7Kt3w+pSUVZTJza+FIXcBjoyGs
4fvQulXqEOvmTKqI+vhLw10NRrIo6Thvu986ZnRV93V2ZoJ+PgQlBpDaXLryMyHO
eg2ErKG93n9L4l0A7eBVcVt6+TUmn7kw05SDfBfwMK5DBu9uCBac/vAL+P+PP8M8
6o7UE52V64Y3iT51CEE66ZA++6LAv0sNDYTtCqNecJ1RKikGZUQRl7LVcOCzPV1J
RIGNPFP7ihP6H8LV7ptQL5GKmjuUoCa9geyL7NbwdO/zvcsqwAKFL/ttxzyO7dW2
ZaPDIrEeZ+mRXnqGEI0yH7kleZuQqAaOD0qvfs7H1CGOVEh9498meoupgnjhP8gY
aw61FxyUgAA/nbrNVgdiINJTlebMN3j0RUkptujYiRYiayeELGIdUEt/M5kYxP6+
RQuUsjch3QEWNyBRD1cVqXqc1Io9vionWuUnZBaQ90Q99Nf1EaNnqYRnzZgAEObB
+jSEbbSiNoa1NQfMbl/+0FfsQuDHS0AU/lMSia2oCqp0InchewufXPaqkTM40J+P
nDYhSFhXGck6useRLLMfAlUK+DKkgnhtL6LWClVbGo2gXuSLAso3WlLRYDIoqn/Z
7vpUpMRDQvTvwqDxVffYwhBXcoquFI9020RHUBvgsx6tkjdhmy466mGtb0OmKfD5
6JnreyxkPckrVKrmFl5ekiFqCC0RZWIBSSICHyB0JeRuhm6dtFxZDZu/WWKvGxyx
dltL9oZIfpLlLZbfz7dKYStzWy5N14gGJI4PKCVpA4ES//yJ8vxmPGx9KxUtOEdu
ebD7lvvCw5AmJJrf3RslyHo/SqRyHJAnd8YXWKYyHWLRDAyH490vAOgfLSaxtX/P
wpW5p+b1rYj0vW4FJoiRomlZJSnbO8IzB5+1hAzY3SMoWjUvKnLID06BSqclEB5J
GFfrY9WdaYALHk/qyQS9jNMLUzBN+ExHse3tGJ9iexLn8iX91MBn3AL0Lxnb67Q6
zERY6MvKL5utSd3la/y4ImmAJSrelxl2DWMD6P6HTtIQgsiQF0Svz++aTvITC8Th
Gz3WDjcb9jEcqwg7jB9g0jpA+Jz+GTtEWPx/pFOra7VUTv2+Cg7PJK9xg5F7gjtW
pFzEvDtAzbUOTtGBoLaLDJQK3X9mkwtQ7fQ0o1GVGN1aaIZoKcYAxMpr29JIBpxg
TDsSkhy2kFj0rol8HrKFBnlk8oibF0or5/LZQtKTFOlF3WDoUpn7J56H9GslS682
5Tzjbhzk6BtlzdclAtzUQeYJV7zyadXQjaWJf4rLo0Wo7H3htq3vJEpYzDm4EKK0
nr/JeoY2aM8NKVnht9/efrGE5Lgz6GHFMXmRkofWxtrpBHluNC1bjZRoFiRqHGnj
MTNPCFQFV8f/s19RivS/7xc+67/cbUdctMtTBgGMLMzu7M1LaNeEjxHvdU9CoQLm
TYH3grqv6sKCgczBkXyg9ihEZtmvFmYjxjnE10jn77z3A+AgEXFeMzmhYLg7AK0J
nKqTMwbBQcpyyyGULQvR9VOCfF89loeDAHIxA7avjbGlwqrbwDU2CuyUWFgFN1D5
0ysTJciNZniu8Yvu1ZUWBEpCUKf1q7n1Soe7tsurJAtLWcqSQZB01QnHd0QP/o6A
KE9eauOys8wPbdU6E/tNX6SO1hBTAt24dRfxzoivIYbUAAHLk8azD4zl4HS6s2Pc
21pcvfBY3P12NmoghexSouYwPZ7RhvenJ3TisFHhqRS/LDeME0DYd91UThqfGdKc
snOu34Fcbc6vWmyrBcbJZP6xr6iVqV0V2kikVXTD2E+iFdswH64KjhjQBf5K5/qq
7luneQeNqyFnTZPiqYR94ov72bF/FzRPwj207Tesy6+gGFhx13asiqStf7oPZmqg
kFW3iN4FqPMta4mfvlDHSEZ3k1t89n1W7SuznqSG3s+JPWK3MuA2v0IHU8n/E4cB
WGKJZDu4XOwMVwM15DMcBsFvE+31de6u3AH4UluM/0GWIuNBJfJ3rzMuePCcE+J3
VCpNQe26dmWgBpLJozUP7lFY16pIY0yWEjed3c6/XGeP6CG0c7mx2VIMq84h71eq
PedOU7gbiDlJikWiVTE0gwuY1D0JTnQxzxhj7UeIkWrBAu8rrVxebWw9hMcmZ7at
wReqNYW8dWGlZDJSMrZPjwI7Pt3oE2vTvSoQgKOsctqMfwzuq/Hx0WDVzUCp/SPa
WTPZk2SiKk1qRrz0bKr/vFe02jFplHjktoh0L1iqCum+fy3rGxo/1+cpoU00Jsib
eDNL6MyWTdx8a0VIKXHUQmSgWK0Yo5KsNOnicpOkhW+CeNmYiJ9JfQgyfdmiV1Nd
1SMKfF4w0xKrU9Z473zl1CB5IqNNzuk469GVMkF4h/xtQlpUPOSQdEgRfdPpFCIX
KkngpW8ndaeTg/VN2qOdE6AJzilOQ4KyNkpW87pxv9eGKdQWUI1X3ThRxdAEEYuq
D1MJjUDMOP8WBXiFVw9ZMoqrvKA+c6WTyPP8T0bSf4GxBUH5ZGwUUwgeHToX944h
dn6aqsVPCJRdpt75IdHQb8ctubPL8EjRea4iupL8igz0Mw9Cmq3zDVIqw0lH+Sx0
aPF3zVSW00aYnVg+OHJEO9Pl8kZDT5/HcIhVDbX6t3grSDgmvgveeJhQbGY3fijV
zCyAEbHCujMiYHviOuk3T/P+nn0VdMKeWb+BTJ5gW1rpQG93B3+JT+qbG9tkt72M
OIBlC5rka2eEEOeWcZLbs4EUPfNiTnPikcN2MRHXSq6D3JOjOFNgGZe8cxhunF1p
GHtMpeJgkl6dkFT2drd8mMxY2/blEAHrscaQnBWXtCVaK2pSNUOhZkroZknfloNB
i0CPD0ZhRmfkebJJOaUR7ImSnJzc4Gd5DtqefraYqDh50HxroMUgR2KIYWOecGiU
yapSrvVkFrld6XmjuVs3e+Pj6DbggQTsDDXVTHaJ4HH1nZnJ+D5tosRKYtLVdpx2
HTM7fN7SIpWlYZSFxxzXDPRImWxlIhctFK26JlJiIKSvTusa4d9yuk6BEMR4+vN/
qk2EZeQBJLSmcv9dENYSRZBOy6kjxgubiiGNwOCRoHMRgNZA4W2aiCegoPDOC+TC
YxOGsCtqTUXroQE6x5hPqjZGT4AGzIgx3zxE2rP84yCmYdg5NVUEoj1QTPHm/XCb
XH0EHJqq0OD5DV9Mc6t6p7Gr42r5wlvjzMfVPpTm4S+dqmhneZYsWcXBuZSS1no6
GPGSTFpdcQmHWrpBnpE4iaiKHfJnCijTAX/+IHhbCToiBB+bbu58ZHEHc/2Xy6Wi
Y7mL6J1Rw0daXmqSAvGMZ5PnVOizOmsWQ8mGkVmEhWUliC7z0qq+PZmqwXP7pYMS
2W1lUrRUGOgPE5esSGznMjxZM1FfMNLC3SYQxpDE5M32kYgjSvAXVgXUm0oCmhnq
xWAHY+kS2BW9hvAgYHWxxh9tMf29ytmgryylD4u861AF+kYUm24dft/7Iob/RYZ6
LrXnZ9f+xW4yKOgn2P92lwqtmxGFYwYH8fFDZyL0AJYo5w/gxFya0Vc640o/lHV2
NOuhYsHtFjWVIw/s6M1EOw0P9cimlATryEdmiOm2aBchJK5Fd0p9rbVdS8gVNmQw
7BFGLAhQ/XdOt1L7vWzYAaeHm2Oy01s/OSaPXrdk3KAZLyvORChOuJ0VfU560hKj
r5Sr5yja8/hOPq1BcNWsG62fNa+AQ3aWX4M+RQXn15V3JUQ4JqSyvuN5s8oKXpmm
V33AJmUVVbJ3SL2nt2s2z58kpYWFKG+yfvSMQDCntJkJg/utHz56Sb2MIMuvv9/v
3pfvaWhg7S5BqX/s3/orgZKfge8FsY7TDGEYKPFyYuQetialmZw4IDUxhe2ew+iD
kQpjEr27PNRF0f1Fbzv/nI6pfK2Q3+3WOgZm0xhSUH9Aiyp5PubyMjn/D0c0kLjQ
yYgvY/WBvgXfmfvppai29ILbRXYKnBPKu2Xr8AkmGoj6+BOku8Qb7kKW3gIpfGKj
zJowJdEpc81KlcR75IqHvaSgjcXKkQOus/MyfKpXB0cNUe2zbZExbrq18M2ZIHfL
R1zjIJXQEOHAXBu/P4kXbECnD2djy/UQ7/3wyewzcj9hD6d9jdx4y9nWPfaCsBqq
mYtgyGPQOqHS5K9A1ZICX5APN8BmFCsKlAHv4dbao0S+Alu2XRUIAeYYObeEuMPE
B1WdBRxNY3Xy4Tv4LVwijlDHo3EEobpER7UabadGizsce07JsOKdZ9VHa2CCx4Mq
0rIHZh9s1jt/vaTs9E8UCPTfEapVYOY4OMqTI/BmRW8xpsaD7/vDby5XbjBU8cbo
cxIzyfqj2QGrqIgAPZi2hKlkR3PYv6hiKOf0icq04V7rK87b1Ec1u2UBXczFxZ3P
VgaSQS0jYhNWa0gQkjcJJbzzCKDosM5E+pN7Lvc21F5XFibUT4oUgBnIip6aJtAl
ANpxPJXdERmQXj1G422mtnxmOz2oOZZktSjwuYYRSM+/MY+GWK9xfiwWJFo6VfTC
wYnanSwiECMkcDc6ossvL988hMxeW5Jtu8j2MoC1OOWM5MGqoXS6ghn3wtrcexJp
EdpL6OScRNJ4T+IdAtRYDmWunPfXpv3YREaZrDaJ4cvM/Rz9q9ILXRnG6xqT/AmM
br7Ta6pwEfMhXguHYEyUVGME1b4fE8ytb4nkdzJmKQnICD9yLZPGygdTzI50W4N0
V+YLdJpK7hb3e+Qoxz+7lafkmJeYbGYrWTEQrCZvJln5JKqqgz6kfIpIfXtze5yd
uZRL+zdSLS41orumOiAl4jhTBdGLeb9H1jzMDlHVxbhhWUOu/P8KzcO1pl/SGK7F
odEk/F61xuGmZxgO/T1kw73EszbxH9HCned3CUfZazh90kuCJgZyst3HLQdSz0E6
xA4oWM2Edlzgp5r19iiwP3c1L2sM55yV0ngdsNmMyvyLQG5VE3vvFbKVcOjQvAq1
WJZEj7qoY3v+BrGbBZqhWCVaaUAr8WJwoqYbXgouN/nQIT+2TUnQtek1ms5ZGh5J
4c0H+y6NpaEnkTx5iG0/aizjpsrobslS9Mjz3QA6sGzhTndtdGiHJnl6q5qXLQC3
xGirBDuVwkRRu9W64WMZqSs1eOtRe9B42YDfwp58S2HEJzSprZVCG/Vo3sMTQ6e7
4wbCfii24+QAb6JxEaFDrdtfbTgM8+ZifmNoCPhyl2gw+cjJhmPdPSawfkhrricP
ZK5j7gjuYoSbRRq4tSclH8m5k1672GXc9fn2ajufnFVYkzwhQDO3c3/C9y5zk8AE
LVyeRyXt8seBw7PyIA0H4cJpBx2xQCVcipjRVippJeKb/Nx4oVkIJrqSJ60jcKLM
nmDrftjGj7QYZvrUU/sgLH4eKo4hYV//5eDB4T7PkKhsfeGpn7cjCA+vef2dL1hX
JqHmxK881Gm51osQ+Mmtu3RKO1Yr6+2e9H1UA/+R8aTjnCA/ekTCW/LLxXV31R+3
B0i9vZc3xyMbVehveYjuRMl/nZTDomB7f28k+f+er1GDzr1G0O506FOKZNCal0fB
lBmdtC+13aK6RGy+P9uE0ofxcKbROZvfH0hDh0DN4/Gn1uXkBpTAnhFL6ebae0i+
x7lmFEQrp1pq0TMVDHk4GNZLfpIoUNlrGPra6oXT1gErhPH4GI3CY0PzDm+d8ALr
RPFjDsG/lSf0CcmN17DLmH+aNx/4X1AonVxpXSH/guQ07lMITHs+/4KaNROaVLiF
nUD5lHQRZcrv9FOwX17dS7Yn+1LILmnP2qY8jw4gch3C7vSjV17S1kgyba1GDGnz
qSwtDMB7RPNGWSCk9sND3uRnsMt00bHEqCfRKmdzzB2O2hq14UxtNLusNx1s3xT+
zJjgS3XPbGcE7ejvLebcZSE3C7YHJJn2iiExhtCqWjyr4OkI9ji4ScvtxxohyQ1N
KhX8f9+4YSrfzrzHeIS7e2NJQVExvSYnRlkUmQCo0xQz+ijCvQsMCGC9M+2n9e/I
qzPrJUbU8U33adI/AX6dmFgbidGzYmLFWHXPcU6CyVG1kZXjs3bNZyDgySHhqv2t
A9qQ8BoCh6Rc4WpNILMOiiuAcy6wG7XvgMfN8gFsVuNy2icOLIO5PZi2C0TmwIU8
lzyGWZXUzQSq6uHAQjHEw9/2Gcb3+7i/R7EbclKl/GoSVHBfVDb1kilWGAZdnfqz
MDLjH1O5Fg/Ly/HCemjbZFeEDtEUOYP6FSZCpASldBFHUCCxWMHXzElAaljxigUw
lRJvUsN9eDmF4iqW/vy5dlewc6sAwDYs4yMoZuP831m1inRHoSUVzzPKg6TNyism
/ZgAa/LhtEq6YzY/0CQxhEOax2pfwgKtq1ArX/7m0b6PGjw2mYJ0zCQnEnlb8GR/
9MQu/Y4EpAsYyzEA/IDADpip1789OunkHbG2CQytWgnzdGtP4QMJF33wPuJ7se23
m62BzZ9MIfYVq8BSFa6xDL/MelrQASNOGaN6YET3OAPJaECKzIVOExK/ti4EpNEw
wf0t5sLGtWzxUJNi8LqbVmG0ggDhS6Q/wxzjWko9w+WMuW/bLFPZ/8e+3FhJMUyC
EmSxIWTdjIMesKtSGHRhpYtGnj4Adeveb+r9Q7QgHNX65wSntk5VH/4b8oJL1GMf
FY7zWoeu9n4KX2ZC+IA76a1c6WhNZ20tNu5Wf7nvwj3P5Z1Vw7f56rYBOO0jNNI3
PUJnoX9OQr7lOR+f7StK8nf+Z3NjoiCeNFf4tjvW0iAaOL7Zn8QlqBqC3wRd28yD
ldMH5mtkH8E7JOd+VTpk49e9o6SnZYH3MaftZ3IyWMEJQI95z5vxahZjN1Ugurcp
fYOd0Jx/2D6fH3Gn1JXZYC69Z8kTN4kPXtu06MLfVg4yC3+i+WXuwuwiBxKAe+d8
XTEFYId/x+Ndw3b19ZvW9HKRtzhLIqVwQr7JGFb+OugB8B6kiD1NtmT3lvU2j9GF
UewbLeJpN3okrZ0fHNPCKzW7aR3oEUsZMyapexd/kmN9l7y8t6BpSSPluzH9HuhO
9LEpmYjET01R0feX/szzL9WjKPiKOwS+DyScbSailo5W84xWommmSXQVU7OjYI/G
pc73PgOI54LOzdq1hKzo5RraKUbNmP/JH1ET7458/Q3rNIvSGq4i2tfrJgMszSxX
uph/frOtThBFiR5rgJiMZDfsKfr2nwz2PH9Bc3r+nsh/DVyHSZ1qe+BUoN7cPRUt
w1kk5xTvYsrWsWv/6C6xIBA22Wo7KvxPZHnGwr1Ey1DyQioEZly9Vt9nOuOhrAmU
IOfBUQKl/BtK4kwso2JzZI67HvPs2bt3/1a5v+iY77siYXdR8Huo7tVQahH+zvw2
s8CocL7ykslsHuhbJuyK0qARHg8EqlF59VZ+Dl0AJEGh3zQFo1T/hGO/TVHnMgWg
PH9koGbsB+ygBI462g+lZ9N0Jc3MO5OUsoJO5i0aI+J6yWc+hmBZWGSz+HhS9AUZ
obQx4ahmUqvUEU4D2RxxMMFAxyVhTIQowmbNKpZ1wz8cKupwLWQbjjic/J3Le+sW
OyL9KYNfozHMw2TSeu6nU+VZy2wKF/rnHZJPXdJcLdjP4unbdWSFziee1zooG0eM
Yh05UIEFUv6jqqt1C8V5ZtbWpisR4wJQrnhYpbSR84fHvo6lV4G2dZx2MNc7W5+x
Yl+nbvfh1wtDWZkbUsygIjAYgDv3XCjQCnsjOKnmUmNdU/ZVWNCj8cSX3aqGCO0o
9zop4/XqywPnhd0LlsogcS1nCPrJmMBDeQTAqWOBg+48DPjM5nnF+PJpTrR377TX
r/ltwy0f4vbKEB+/0Wza4AIA72NWmudwLF8O00ALoYiHKwoEA4F5V5Y97PgBvTFs
kk2oacRhRmzxKythEWrK62zs6/YpCMTtO3PyDolFKZnMtw3fJHrtVUUmcLS5QUVX
YQhjsS41JBE1Jn6DfXGP6eghUhOXLWJDDgJ3P3Mw947hs4O1Wai9BU8y07KEECaQ
loHUbktgzoh1fkUiklwo0pWdrzznGhoVW05pt48Gax/Gt+QAHmJsoAo54bXs0eTA
52/qj1md7p/C2jGfYhd7txzdLLYjIeJVycWLS4yPzg7bSCkSrmfilgYJvTpmXH5w
1wlq+UdpgXbQYX1+JCdk/ay4SWzoR8aFuhPjRrEbSp+QW2MCk5bH64QFsKoxdERq
HOxxH0VBLhHMFsYlQpRtPfyUG4xZb//d71BNBScXfqqcCWPiL9UPk+bj5ecpMpo1
uc5xx64DUNSWeBZD3z2s/VgDJUoMgG+ffMW2zpBkRxeMcsqPbxsLTN7AvePZys6A
oDhmJywLktpRtcFZ2xSTxRTkEuZ+YeDvg17TYwT1y/MVArDv8nwN5NQsngG3nBvQ
uZpGea7iJRTUE/b9xhMNyBTn7ffKXQkSt1zob9agY/SxL5EWMXC67c06nDPm3wDM
Vk/AZhCWUgUvSmvpsYJTE1ZvWbOZssSjzBgxdmm53YL4c0LZIIo0jEWJ3jbKeqZ4
EhqgffmIn6CF4/Gyn3NuxSFECoZvCCv2Nnp+9AxrTnm/wePZRiEijmiC2pgR7GyT
LAGcYDHHcAudE9kvJoY6netqVoL34B6snvtdTmWQWST73AWlo3qRw1jqmjA6p64b
tz7cK4eWHOrIePRTTCjo/OnoGHaL/HpJaV1fuTkYrfr1GeNwoK5LTEQxEddKy0hO
CnZem5J8JVONDu9XtqE/OzYyRuEb0ke4eZRLs/THszFgZ1MrIcB5sffu8D1UFFdS
pOlPZns29ZaOMhbSbasxs7flEXYIBMu2K1gSK/ym7Etih6k2mj+g4maKhic2jPH1
aOJrcHDC/8SKabmeTgi/ZJBdj97HGXeoBZysZJqDhLmL/5/Sd2yb+A6QPP2nkbwW
ko7CCxIkXtkgxQ1h1s73F+fWbIB5ZZ2mLxZ8J/hAziIznOVSEGOCU/mpPIgDS/0s
Dgw8uK1fiXUiO57HE/I1DN1xB8vOjFaPbfQpqqRXF9vTsTErYGBikTwMvDshjs1f
uXpiPF036EBaInpI/i7xpd3VjHxR5ldgBF+uABTDBGw+h0RBDht3qPkGqZGPSCcA
tQNmufQQ42vgniPxKAwKzCIycws1TPlsWDVtl4M4ehlAxx3t4bU7fF30nuCERuTX
DOVegfXxXFKYpUmP6Eai2+c5EmAJv4P69mfejG6xaQxZ4B7VeDQazGO2UHwhPY4u
TEwCqZ9u7FUxZfo7oAYx+a8JrAXfV/EPwcqwmgU0J/g/Rv/P8wwk57FwgPpKWD55
R588trDcnnGk2I/U8nCm2D2iUDA/9nAcO/52yv1gmwMo3HHgYElIK3Lh6wnmu1N8
rCRIhRdy0R0EVDVeE9h0hiM7ex/lc0O5KB90GLlcVucQvOhnEkEWzEMUbmeQPH5B
qj7rA4VmoojsQ3mzBnqtUGZmm4jgPwl5CKXyxp+6GaNDFVfc5C9126KP7XbkSgFK
2jpjaSQU/zrDEqeOIhzgfv3K6l0gWX59iOiSVCc3M7J59UE5QtjG0k4uU5r7sXpM
Z5Kroo2FJ+8m/zbtvxazaLaDIK0Y+VB2U0q0vbcWUviLlkhNaqkS2DCjSxTimCmu
PCoSCpwxPrk9JEOk/L8IRqbDUbjcUIx8rhCt3AY+7nIr7nepox58UxRqM/YhbC+H
8fY2SyAeF/ONAjAEeVstVDYoE8cVBe9EXBY5O5FZ0fNFQudMqV4okB0peF9X91Nx
qeKUXiOpw7mW2ViweYD1J+/V1KSnFDWwIAS0VwIkZaLZfKbd8SUAA441oYar8Je+
IFVBVW8wOaERx84/VMALoD6oNkFryykPKvIHstocCx8kofYxBJECpFquAT7fiV26
JVFJPCxSUWrc1p8EuOhDgGA5cHIFaBqjts29TgzSu3Bp54Pwig2L2H2XYejfPkVS
wlgN85ucwGU7Xt3DyRvAw3H7ieLZY7dPJLIDX+syKCBML5R+kz5gtDo71XkEUnSj
YeZYJNG35jQRJ5s9ut+USOVBKgrB3YJmsx1EyXfaMF5FL1fo9pcADizYUJSeZYRG
h9SebRhi0U9QsF/UyPgcAItDFZhSqQwBk3NutkbzHF8sHIYmm07jkqIFkB48C22R
6sr7TO5KC4dqazaRdjTZmKybflgwE2NSXfrbgQqmNoILFvDU9+qE0UfJjKmneb+1
JHFZjCNKBwAJrFiPvQkHDOC5IyHzcHCJD+ntr+/d/uUqbccFTdZw+z+XqDiwcJNm
2cGmqypBSu+dQhW09ujleXv5/v1GS0en4b6lvwgCddAixymyC0VtbtXPY8WaP9Wm
XTcSk+/Dy+yRDMafUKuE6O9TAJEhoGB9EvuJDVyCd77KomOiXnCfyDu/r+E69KtB
bIgBSjb1sNSKaE8TQQEE6F1Ya5PQZT9+DZmQq/d72qIXnXMdCaQigpnuEPcslO11
xJTBCyMBvaYnoWBJFmgGNRil61/Tni4ls/lvRUJ1MzidunTLtohjLsQWDg4gY1j9
kMDVjhl7kD7iBO6XfSveaoM2YYsX6biZLDnFm3uXceYQ3WssDl+rOLtyG5ALXKll
T8IgEf1/Tgkcy3YKGSIy1QClJ9WF98oZe8c079LR5Sx0oi+rBxb33uS7b1ezSYfW
WYIRQvNqgTZnQ3n4xFvouWjYmaURY2ZuHroEKBoxY8RdXtDkk+ZuhsWtI/4kO15J
QYMMs0caBLxebUII0ydfNRZ1Lvjy7kyJnGX9gWOaIJ0rTt4AvaOOANCkbQD++vH6
W9n/j5joQ0XcbwTCsgF29Ep/3Y+WCXwNNYo7/UbbGWRnQuUFOLXT7e5DD0k14UKX
5nHOOMsR1qHVcXJL9+0FSPYgw+osmKTOpFwwvGIyz6/0Vh9tbOZlLY8TyzEseBZI
70d+H/D6x7ORWFhzvjJajrhwhl00sRXEXZq2V0YRePU9Y40u9DnDuVKwrq8DjUuu
OoeXDX/m66jK51+mDhP0td3Zz+2xB9HAQ0blbwsqn7R8wOI2ERZmfqfh9jFH1Pbe
4Vsar3hUCKjaTsaJ3RVydXMF9ENDFqw8hlg7RWIO9WsXCj/v8zgQbiI4Se6+4JVH
qjLE3k42/IT7O/VTtpFAtvfF+DG9bVdZzbz9/PFhnwpdVmz4XzuNaEbM8uWfN7uR
ongddnkzt2AjxF9t0QO/11lJxSedsXq/Iu7tQCl3EHqlSV6vhlrPn6NHEwOXwZOH
eUV6HimhH8iPzxioDLdIfrKJhcw07GG2MeAoEyZGi6I+h0jn94EUlSxJYBCiyb3+
1UdHRO5tTb8JCrUVtbj3NpsugQi6cuPJI8/0tpi52CK233izBt79hiCrNdaigJVi
ZVxLEakDVQWkw8qLahEA6VZTkr4Cd0MpsFl8+syZiGhL1BBSxHvUVSBm9/LFAIh/
4e2FjD6BoFRVFWojMoCs81jZRHlnAp3mPC5HrO7dO/gITPRo//kIbKG37J6UvO39
LAxu60IksTDd3wsyldBIylB3SwLjqjnvPVd65lFNmjBy8UE4pzsedW+hpuNq380m
fgd5Geh6POF+JkLDLzGWSiOw0Ippt+YdfcKzHrxKAN6SvU7pCIDfD7diNIjBn5Wg
crrFKBa5bBX0Z3woiH7tZlEw+kTx4mfXLui4oSfC5UyZizUeEhulJFX7R9z+4HX1
bHFMqy8pm4yh1So568EylMvmvNZqCkFK/KkPYhvnXOZSXMO3KhgSFRz8xAGe958T
f8JuRIAZ9D99XN2CCUrQzv+Au65R7ZoSz80csO2/cmsvHCkD8Kxr5Qp7W7LKy/EZ
DQqG7p99bycYBQFYp+t9F9iHDxtqnqxd4P2YNLhkTogR9Yn9c+vPRee5418roxLE
QfzgHDmX2zY8EEHWY2bwHD3QcsviueMWq9nWCrOWjp4ma0BDFoH8+cVGRFf7B9e8
N1hIk1yJA+mciivzghAY5QvqnlUq/cF6hW4RNK+5OiWle4Nha2GQOrnLXlurO6Ki
xnkZTEeDJyEKRgD6VXdoWvJWtH2fcVBCLgNT/I04c9SnWllrSGXY++eGryLkiny5
4oAJIUdPN7ewfCgGNP8938Geccd136do6ZEx2PmgmucBuVlE1n8Z+/1UoadUhg+u
rOepYnEyiSB812WdTBMm05mOBc7XKIwNf5nLfWAjiPiEfuyaSoXwZ5vzA2+bVtp0
VJS34xaqET0reIW3zEaznjY9GMxizQ+TDLYCbu7hLvsnZPQzdMvvVdFRHWVHpW3k
hOVjbRmLMlxeetsS6l/T2naud/oabknSfN3C26Fdw4Y5s9FocHDGnlRkoMfYTxpN
Z8ZabUSIMk7sBP40fHCJDtOySO7sAZapxJ+AYFzsbW6t0gVdySo79BVjtwOXB7kE
oituLh8I5URGcBScpqz0EwAwd5NKISBGL/SYonnf7pspky5fnJ9Jkd447MxT0d7X
6epRDuAeHw2OrEtNZac346MhrQXPQQ00dZU6l2M9YnDJr6eiHTM8Y8PAZHGGlkSb
ymfACkIU/jvP0AiGpisl7/5iG5dk20+BtRiHrXuxWwA7yPp8Hr56BdWpNi7POQMa
XftQ/05TrPLyAZVtm1wWsW3EGAjo8CnTrhzyK8P0irLuwnLOWYyGZkFrK2+N1wc+
+S5mnvezmd9dHVSIKuClaNLgQo3Dva8Qbqf2My6yvv1syB9t84Qjxap6B8/o5l2A
5kC4NqyPNkIKkakUKSzwYWdrZg+gOIaN2BCfcU6WpiP5wrAQh0rFnjYaPhwBgJAQ
boC4BQT4SP3ItbK5q/qLzhOzVM8j3AOP/5fUrKWY5swjDl53HKLqucHxYT1ezgzi
0ZB2R4jot5+1dR9e+QnVr3PVsBjfuU2Cup49MF1nbADR9J3naE/fZS/cMGqsTnyn
JY6Ui7bu03qt3m24n9rTL97MN4LUCu6aJRLGw5L+OaeIonXzjmd+0rxlmCgMuA9l
EVn4DlKFGOPdGcsIbY+ibAKgbKDhugj1TUBBCJL396So7P3x4iM0sIr721OFjh/D
JYqCy/K6disFE/c0QWtAALYGgd5oBNULF4DMjYeqPSzpYubznqOkGDLSKRnpC6Dx
HeO7HXQYWkrMgftDDj0/uVn2YWwfqhO4ts/qGwidF0QHXdZ80IiSLrr2HD+va1Db
YuQ7VIy3UhcSiQ8jf29LCAS0sMT443dfh1cROCTwerFrR4I9/EyFcA2/tRoX72Zp
Ff0fvA+bWm9hjL8QU29M1NllbCUMLUnvjFgLsHAtxqIunpAjneT+xf9V96NgS713
CzNfFA28OwrOTTCm7TKOdMQENmXVxu38cNsLT7YxZdZi32PvIAkga5usmwf/9sze
4Ad1PJ3QJqO5lQ+Xa+2q2KXMaFNv1YF7mmjGOqVGRSMNagDx/NdytMR9McZ2S9K6
Ke6L5LKed/vLDfYFZPkxKWPVsqzTOWWB/ea6v5OXTAczSpLHbYsG+6LXCMpJcvu/
qQcbpYx0pMMoF3ue/RVvj+L8zyocsYdM++bpQvJOFI+J4yxaw62/gBLGpmKrbJZU
lXmKIVfZ9UM1RCPuW33klDNG6d1Gf1EG8aT8CF3MWm008F8rYN+QI7jzVhvgNFBZ
RWRPiTRjNNySHLTTZu1QIX3xUIxGW0ssimytrzHohZoY4jWMoGWsFFqYCCjFsPe9
GChFry1IwQwRk0qoZ5vzyEKqJia34uK3vXyPcBC327OSOQqbq32JUGHErZrt7ZYS
mhdDzY6ga+EIe2PklBmR0VpdZ34sxHtJbZzBPwBIvX1t0bsmMxuLDGGVYcCeGi8w
mbrhubSLxYJxuMbkysahl/Cf0SDGmzNYUb3X1uF7GOyAD5aqafb792FLsJ2EZZi2
VJT3R44dcG6j3162ORRXL7wlN11YS+URpmXvuWECr75wCw/QF4npSgpG9QpZUXx6
GecXVDRghTNwcW4IoksizvO/C3yBE/TLH9AKX8JpP3DvnIBp92vLC75QCFem+b/P
YQb3GdNHKSWCL3Xu1PxTpy2QfnbqaA//BUkIAS22s5Y6XQrjfkHeasYqisxWvOZA
/310cqxyGuWa0d1qBuj6qajQ9aTElrazgy6Tj/U5OU7/iWhjQpiA8niM4p4u83Sa
3VOzJgCXOO4QfAf1D8hhs3wp4nP1H+fE700AECFsKB268J/wNUXHQ/OemAn1d4fA
ChsPWXGO1Bd3VXjC8ACKWNGlmN5N62z4y2rz4GaeV3h+C8idAeYPhTbWdXORSR7D
Clg3rvR+OjVMsLj5zWhw1iOdvpTzjm9lwGCly9sQfL/Bz8w/rq/VqaKj64Jfg9MO
laQ+C0atggevS6Wq2vh/8aRf5RL4PhzoI9SOx35W29VQkW5erSkxg9Q0tLEx7eSP
1u/CWU8EOBkZG3TeC9MGUks4vIqG48JYHw5RvyxTd1ULu6X7wDj+ZC+qk60hzI15
hZMjoku+lh5+RDqvm+iAaxhQmV7tClANKKoDAXhB3B1oaO7LPqQkdq9ej/xi3Sps
/HPtMGDpWgr+B0CDHuckV1PQ1RMLdoKN0Dxz5jDn7QFQbaYL6hDpNaIdRAe4Hv+d
NoRSevhSWaaMUNC0LfLxqYAB0tE5SGrNBcPVqPkJOv+3emkzUNWT687kaSuwLZWj
pncxyZLREzgBsceSgA4hw1f/Dw90XVKZUT7Po1cO9ARUH4VpD/Lxs9ir2+JF3OOQ
4CkP0CmIYiIM+g+XeeB/7tfyA/OZeMGgSl4r4/FVxp9wC5JalQa9JoaA7t1aSSoZ
V5gGb6iCuOPu+D8VObUjv4iE3rxbhoUH2r0phj7tjHuL4IRFGxv0RUTtmkXypq5l
CloyAO4fAdP8X3Na4ylfYk7ZLbzbqFhB+VWLhDbXkeqwQmVojyY54CTClEeRpD2N
N3KoCQrgjRtIom093ylJzBkE6feTev7kK7dNNk5dwnBpBASpXtXruPf/Hw45YXQx
GC+f/l/5EKKNAVXS1hJmxMUjgI0bWkf6RSXGyshb2wblZ/Pzarx/RQnt6DdhIKzG
/gtX104ZoMNW3g51WTngHXCZIjqoY5VU076x0pzZxnRzUPCsVCiHBml4kqOXTVp5
vd07XdCOaijfSVb+yEZ/FLa+hFtl6cp1cradRBCxFU+Ph4SUx89xpnRBril5t4cs
Ja7EgGRMhTW/ivCYbWRt+vSa1CnkAwRu5lBIVQZPK9sYAqoA/oMC1olz5Hu1pBGq
VxPP90QI7NRxbaskF/d53FS6C+PtDZB0JM3JxHsnRwU00XOM8Se8JuoSRIe2PEvs
sFla2sMkMzXEjjgsSxfag+nuj6xB45X0LNxk02/pHAotTbOkVqzh1SzIlvQZe+Bu
wc8iLoVj/BQEO0RPNqhDpoqUrELlbTmzQfnBgW/h7y+slQTJfXzKQZCDv3YH7ZFt
UzC+h5pzSrYhDMR8ZC06reFO3SV/AU9rSL45aks8HMxXZ8Mv5PRagHiQRhDTrz3X
7wxQo6SyxTG2ESG68KQUIRgL8ikBrDulmUDT8dhj4YPpESjA0z3oyvyp7pe4FmHI
qYhOm+Xb5fEC0/w539eHyov7irsZ0WeoLT1MkKSYLrBFszkx2NCLAmNyEH5bfErB
A4I0YWtX9TaW8W74mE73c0dhl5O18HPs7ap/2HKwX+AoetFUzHbx10MXRnd/WXBF
AAVDAFlC6K4eWH5Ao7R657duZtwtprseMQ+Qu4PUvHWiv7Q2DvExestZpoNPi+h0
InCJqTqyQCpS8eUluaXFExlLc8O1TuFkPcTDWMLOZGOwoYvOn2QafllINkx1xFs8
SrxJkl044lKEU6109n79kmX77owndAFY73xuutZT32mrqNzULRUBnbe/ijQ/rIa2
GMZeXhztxYGgOEVICoPmz48m7Sfyh5MSfbXRzH3HdztDYAxhekw5J1E3l1WFSvaD
BJSUxIQ5GuGFOCVykC0LZ2ENdtASmQ0F2Hd/9lw2D1sLIxYeo+6bCllOd2cikI4m
QKOC2eHhxPYK6ouISGtcC7WsSYMlFZ2cFne0jkyL4U4Q/IxBuNZUJUlrRZYep+ED
Sgqvq3R6Z+Scm9UoX7R2mzaIUvjoXUzyj2ttnQL0PBl9YEE+6jyy2CzzTbRuGIIE
40NwHGiOc8+PwpdetXBnu8m2OzAGDLGrMhEHbcZY+XoyxtESS1u+GnothYepfjOz
czMhZdwAIGsSFF4KhWDuCO43Ebez7hJXhZP7pybFywgVyrGlHFzgQdqQfYpJyf7b
+1hPb2TRJux3xmQmUk/AojE8OY/p26xtjXvZlbXK7sXybDkVD8TZavOmSMTcIjBe
pa4QHkKe4nYd/gPopRcfmNqYIZagTHCBli6DybvmyMWNeum2eH8av7Yy4ZyYfwQf
cY0temwQRyjJwRP5nJGIesnymSmZU2uYe21qDk0o+xjKXa2H2fvx8s66VJe6/awu
csDGUmSL/t6uv2vvObUuHY/OggT9FbjgYhWVVQFQSr/VcBpqFxlcmF9GizxEKnqd
bXw0BK5F8qiRICjGnVXZV7BLyVd3qAzbN9Q1SuAsWqVl8Y58ro8NcQXFNzWvyPph
U1jQ6gf9JsyhdaEgRba5Vxju+SaNcyUvNeVr5qFuA31cAGxHXIDm9c/639FQzan4
hy9Krlwp6BGw762kzeaS6biuZC9h3kU9zduCkGWXASGiffDPFhKylMgclYP9Yr8H
a8aQ0+8QiCN5y/w8mzwdW7UQH0o9wewXxPJ1UAxI8mRYz2v4upcSi4pjTcOZa9xu
++xY1s6vQVznjx9YQBzi2+HIw6x8J3BRF2UWkV3JDxT89JiHbCx6ESAaV+VJ5CRv
7YyDEMm5F21/INTtlRIoVKNxZ/0hAT1mqF+LZ+JW9MWwo0Dg0TRdw6XLxPwm5zRQ
KRIJLV7TIqqv06WEYZbqlwCje2MLINecZDKT8QGH5rs+/mRMDNSbPnX1IOqjK+jS
2z+yHSSdVyGTOSiZ7WUvMIFKhMjuBYVdvpiCynzVf1LgYABX0wy8xVAlTjNuC5SS
QeYJdeJ2cqNzdRExO8sNw48hdm0LVWYGh6uNPmWSubUMR+G/uUI3hH6lWdD1jQqJ
92m6p8jBeNSnLomeDGQJHV87t+F+jbLGM/Y5k1Y2J8S5ddSwG2sbigJxvlQZbXOD
JlBg8rc1aqrKFbwJFoAGNNseltc9HednoubF201ZMJ7AFGBaqfOKcErF4QsqJy+G
HQ9fl5RHGM2LsxfG4XDgLCwQp1wy1vRyjpsKUjP4xLBTf0T4/ikLyEAVmZREy9if
43Qodp2XhCjK3XKmjVxYheSrlwyoC2oF3TyVC7HDfuK8pwz+8FC2mUy00jZ/Rh8f
Tk/eS3qDlR1zv4tbaa/fomrV5CuNVqYPANhzSuyVm1oz3YcbqiLXg6wVpfaleFpg
gSWxPo3tTkddfm3tbpQjLA0XXy3XVTk47tgJxxdmstsbIt5c0HOe5rgGxnhGleSv
PIJmxhp9z7DMPP4ezQGUP4Z+KzOHx2StFLj4bXvBOOv2ExD+lWvHphbKyAjWeMVL
RDzKZQ5706a0Ej1i+Z/4A/Wm315tCP1/bP79wJ1rRGrq7oRlxfQwLdjIcNy/cf2b
0Jhsw1h9C7VumaYkkC23yd5M6TRtnT7oA3bBIgg9194CVT4/dCDOTV+F1L0j+KCb
hZQDFBXQ7jH1nkujR/GgycwaO4bbOkkRA7ah/aPYnEMZpo2KBR665OERdZtQ2fOk
L2/NRC9LSOgAuR+UpafXFFkcuUwnMSCwttOWOK6/hvnWB21cCiGaCN723dd59HE2
Kh2xvOraeyS2p9Dh9xofvLw5Hn/D0eSRN5Q0wNzqAKnWLD38W9L+cc5fSI+pDdtM
lkdxxOP9yesKxYH60s9Xe9AKeoWVCRAaYveiw22qQfAgbynKIV6Ks1Vsgt4TmFa9
U9ka5v7aJgnap2LI2JUPtVedQcLs87/XagTpQZr+ZrZt7aKwnj1OHTSNDjobFt6c
B6b87HV5LiXUhIWH0tFnalIzC5kiYiBKShc2ANqOCsYl3ByQcOqbndIHFRQrdi3U
r+vJOnZ/65ZCEqEG0tVYjzwOPUtGxeOw4JzOqYZFLGoi1hd6JxoZ+JdkZJjxK7Kd
2jWHcjMCpt/0K7Yjys9c5YfcBg2nNR6NzevFABpHXtb6FpDhOgpN78j2ydg8njWk
2dg6/UJRJac9Us/XVFeQJYUBDYfCLsLf/43IqlQU2yGW1xaUn4VaWxFQ971fINW2
zlZMpIrLdDDpA5gKb7cjEVyMopLc/Hko6NFRUGhqMXcVZgf8+qFsgM3qA0ZNa5SB
sTo/CSqfTZFrrQNj8fIkY5LfS+iZf141GJl8H1xBJYysb4QMiZjW1FGH7aIOL0H1
CZ6rdjmdNtN4seKiJggyz//RY7rs/vwTGAPx1WJLJykpZVJIcjNULzPUlBWqHUdW
zGACW0FghMLb3fRikUqFU4Q3My9Q4DeUwX134P12GgYiKxvMNE+NiTYbrZ1r8hP+
jAxwV3ZYuivsFnb6fUwt7Ufmx5lidN4Akp3wt2ftSnXTmu881MRYJpshsRJfotzS
5225RWSb2k9KKbu5xrQvz5o7InAIsbM173uV8Uolv2faFkjnuwibx9sln94BFJkb
Y0aa71dVqvRMnnARyaFW8vbMNnZDhhK0E2J4VZ5O4N3J/mx6ufoWw9lU9ws/+l7c
hotHxjBgsdLgum7C6uUVcdtZTPR/znqvp0r0PvNhLNhG9bBZnHesoiS+nV0/N8Ck
J2XLaa59p28I1D0vGqHqh2WkA6HXAkWlt4R4W2epX9OGo9/IJvMQxd8JgBKmOQvZ
k/TKbit/JOmVPycwRgm67B72+iN8H54WGRzv0twibVQBo3oqkt2e2Iid0EdBFZEV
VosqwnXkENRHvG71gGyaE84vlcyzZHVT/t3mxkCxASkUFncF1JgKr9vUx/OmQePe
aWPbiPYZWjR7Jydqn3r4QDo+A5Ueh9nyeGRWHGJk9w1ngMvMIubuYYR89Kli8NRa
Jpq4gop/+rLU3rtvDnfXZMsbZBLit80a3Ro+6qdHCyh6AwMsee/LzRs1eLhW9+MN
RFYDsSPN2q3Q3N1mjXnZMzZPRqr71+O4uCSF3NoE7CJpx3QxZH594DkxT1e7NjJW
VcqaKGdT/xhMohDw5Mh7z8Ztxv8vHmx5gvWsNSIHdW2GTb508O+emqAgPWZHhyVk
q2xn40GbrsRZyPAsA6UhboPhcLio17U+LR40tFU59n0XHh0/7x5TasiWpGbeq7QD
zY+pdovNhAEVRjbPqMPNJ1OEe89LwkGCMXFjE2jYztLTHIVZxc3rFH7EWr5htAqG
JdcR5Szgl1eL5HD7KeeEacDyh2yW+I2Zff4T0xudOu76Dm8rF3LZiOJSi6Rc7/OB
IavLfgHW6iihbk2b7dqDClggMYs3wAkHFjp/6EfViV+h4pWv5wLyxfUu2yU9lueY
FWkbVjRFPWCTs9oIj0Qv6SaapOU1wXP9nyXJ0cWnajUmf7fR7+L3ElW3ZHWiWa2v
UJ96lDCh3gTw2KeJ3rx+4t45gq7CJZLknIyM1H3LOyjdgF0U5R9w67WKkCwuiBP9
VcIsA+9TVjUnfWYOrtxlUKfs4mwSLoHCLO1/+yua7bKjJpnQSj/WiQA8Rqde9YpC
hZD73pGeqUeb3qhUiOqKk2rlXbwZG5K8z8sYa8bxe65vug2Io4sa/bVLBokOWGDl
x//qwC6oFo0j2ZgY8A0bxaY7ZAnKkQe9/UDMj+GBOF6kk50qqqVUXL+6kvN0G+T6
6ze+CsFdec1hgVF9a1FG4ivNYBSb5IYie/d4143rnjjH7Mw3rN8aXtFSYuWxBmYI
wK3xhIM2t3fAN1ADDv23oJYlQjf4FxVbhwFluaj2jmHEo70hMtxDtEuNBOycqlK3
tuEOE9sJt8PdOcfcp5Sd2Im4u+thVbAWNCOue7OCV9muB5JeRNrCsNAEPgi2ifUq
Q3tElfwRxNblgNTIfph4twxNdi3kPEgn0xbCqPLVzzTFGEsUdgn5D+c4VI9h0u/B
0fXV9HbxCiqSehjWV2+I1OKRLLZV96+FBVbUe4qTI4q/KBzUfHNKEmtPQ4GQB/7E
QOh8wmpKXN5RnGYRiRAi44oPJctvXBmUGoqzo9adgPhRVRoFSIzQb5nya2IBVAvk
ppRyW02082B73yTE1XEp+zVLHvEYB7JL9f0/Qcrzdgx+GN7vc+hTVNUez+dv8ZTQ
kL9yYIKolm/6CubRzUgfKn1J2KEmipGxLpNITXQysoGiOBwVVq/vFKN2RuMnM+Pt
k/K3a1Ot6h4ZG8pI5j23SetrpB6TSEY+v0+COjRxQxPp28//xI0mJe30PHIsrv7n
geRFzeed2qdL/sAhkYmLE78Rv8q7MMGJ1uBazXuJ9XTqJj1u2ajkzzB19j9wHyd8
yxhR+fHF+rPGUEXC1AY2Bb4pQTdsLvhf1HjyXMZf7CM3XOwfCqlLHnhdR4xNeTi9
nIbgXeAqRy/rEsebGXCskKWX7dDr1Rk5QXefgzd8vo8TJi7LXz3y6zPM0cLrMA9K
OKJ9YP0MOO+aYecJPvR/BvZUmnhuy6dYzCG7gcTH/p9ICYT3GVEnUqNJb1jUTjVD
s7Q6Yu2VebXlAsAuKfeGj77vW2waFFJHVdYlgLvViolRPYDa4b1ViuVKdzr6GTjO
iQX8Vf4QBk3sI57KcwuVlP9yeTm4KNb89eVCTTL5KdHTR4wD6parpwH8AiCxdNKw
6B72UXsl00RAKPONyUEdQYGu7EizOpXF4NXRtfgNRRMQVs0Xg0mR7IPxfwHX5n3o
zzM2VR71tJlAuGu28i8JjHpMAEz9U+h51nKKHDs/7FNtd0/of7l7muO9yYPq9h3y
TQpo9U1n4gS3csZCTVnkWQJog7/x75ozHQZtgZzByA9w5rl1HfiEdjxthsTSOlfC
n507Z6qgbVqjZedacI9NR96j1AqNIirCFI06R/0h1GH7v4m2xAYxkbULi7362Wkt
f7TwHymiYTreHmM9Sx6RhdQ96pxkVxcPBnOeIT2KEcmEU2z29QMuBVqgWibX9VMD
T+mtvevKw8gPG1A/SMMJyp3LTcuBzvuwICfO7rOMllpJhKh0ptP27RvHlJSyDSgR
keKrlSjpWGO5Vxe/maNGZdZE4rTD94IosBoReff4YCCy89kPJxwcU5A43PbC7W3o
jz0SmtAZCil+TazY6wV7rmz5nlKSDUoZUM31mrGlSvdZOEO8+N2tMN4AJzYNsjxK
9UZ+eF5kW5IV565YBcWcD87bjsJsUQmK7UtiTqmabTUGUNi5bq8GBHrppC+R9YXn
6lDD+HguOcAOjOfW49hXeXNM88WHVZYRbI1fez0e9dSiNh/sm+Mxu3EvlPJDfLw4
mT3crMLa79d+ztTlE+zvgZ2TqJgxpz0BfO45hMnxQctsHGnH6/Nd+iLzoIQdy/fp
hoVq7bsReD5jXksT+sCsU8qn8/Q1LJPTTStY82uSESfI8wP3K0+QKWA4dddo4Iaj
VTEFbMc0XqD11BnK5GNe++Vb4yjBndIi1Jlu2MDx/cvKnCCaBEHIlJQdeQavTGIc
czMqUXE4zTEJ0f1ThTEB4Nf4qvkGfGQG4YJy6jIMvLo9FTtlFtZ7+dLJUt354mfv
1gUz3Ep07kBphDMsjtIjVy/ZF5CY9FbsFSe85I3o0uiDHIyFITWTt4JbD4LNGLAx
BxKv4etxrXH6U4mzWcUDibQaHMpjLMdOT0B5zR8w4Z47yBx3cZzCy5dDDb8yzl9c
gn3tXe/Uy+ym1GvpuFhb/76bPBo6VZLcpcEyvDcys9sIhlHWLW6h2y0EOc2D4nmp
Mci2NTJG3wGuPPLI0nKpEAw6jC8bNeEmHyhCWEYDSHGVXV7nI6w6fXFPIqqDhg4k
ZLkLyQBJ0zROPBTqq+1aqBhXh9rblnp5z9u+P7yTQoWoBYC/xBOiZexUVinS3X2j
9j3aJcFT+k3nWjEdczAhaRFDKqYZmuQVnPzk8HVgFLavJoUEOb4H0HeS95xiV9o4
JI/vmMqVYIax/8WZmVOkJSSFIH4DRm4Cm8GlLiYeDQeCdh+JF9DtuymTcHhFsKXL
dwxty35bwYHtqXcotXNwJGBVsY/kzIPP814KJx239dW21DMqIyDwmd7WAgch/nTt
P+JH8io2PWFohgottVRESZthnQL2F7/b/BlnT53jg4uNayHYMJ6alvRLrfL8sK1K
EM95dgEdniHJorKy7cIp3qbnuLce0mPHM5Fd8JNw5g7o2cApaKg9jc7ADxehKq6c
Z3DBs7lWuaXsVQtO3qZtQ7XTeuqeqmnKQU3kyhedcK5l5GmC9upsQlJddVcwFVTZ
o2vH7CqQBebc9Ml4N6ULhHGPdKXxLKzMQALZSdUrPSfz9i+o1T26tbadnPFyEnXl
JtCeZwajnusRtsN+o0pB7nm6YVfCYsLDBSz1CZ8rLS7or5xBsUD4Spt44tMpya+A
AcrSNoN5XsRML7iD4dv95a5gBJs9BRzMO1wm+8Ybda/xzYW09B8jmr+rDlNloTsK
p4E9d8rNgaWA09k61RwU2S/+spQcVoTqykHbPC6ROMc4YhAp8JIE5BQbxAumhIze
LsD3CpxoNBN0CTMP1m8VerKmSeIFOHwJATsyEfiCpiPL4HnKcSQkIQSIY5+n8Jfh
Lk8jyPhf8GWY5smk3iAE0138bMv37JMSohH5M4JNmDwNlkUWjWOTudZSGa+VX7VF
zgyyU8MMm6p4i4SCbypQxZNx6bE9el4QcRS48P7xwHst2YiPnBCBRg8rdkwJqIdu
SWJggG0fUnCAZYOX5od3u846KwcEpVnvUl4A/h1aHPrLbNlTpudm32bDYQAaa9WW
BRXPcjF1+srWEIStCwEXOZ6yUdttzcu0bkoJmIIOxsX8+rkYW54+PJciT1GwpXsG
4pJkqP9bmxyVFqSUFyvMQ1xl2SRYGN8Sfl2wLnT14NXaNEHt7Ux3Wtexc0dA616y
j7NL1Fy7FSZgRurd+YSzYB5J70ce39ek/qhZaZWWUIkh1we9L4gLtxyMeMq9a1Rw
QFCCRwVaU6GFnynZhRG02XlpkJqYRYwE6JLiNisIOFicl1FoBOA1uJtNV2UJ/RXf
ukmJxfnU0OEvM5ccLmNmY8wPzecJWGrhbv/8gDILTWuEAb1Uho0Am9+xDClez5Z3
gkgF6fdatcBejP62lDAajau+4SSsP/pgE4WOw+5fFNtZWI5s6Zj68ONMkQWatQ4d
tl66DlTHZd0AIuOiRFklvAe834btf9eftCjPORRm88zIYaBeyYMQRF+5cSG+6Ts9
ZHckowk8ZtDpPi7k4YHVDEIHTAf8SRSKI7b0EjwaYrmmmaYxiEWVcETxevpm45eV
gr3HKCdEBkOlrZ2osUEN+tK9b379EHdCVK4fIPIFVkIPU+kpNAMCuHP+lXK0+CM4
AfAQ19bc5SI6lcwm08r9S4SR9l5BvyGFO3K+zocmsXquuhQ8DhyCFhn36CWHWr8E
7jqOdXJX71WXDgjYcnsL0ZRibrEwNXVX8nHONaJAWomOgDBlTLFxhDTEPcS6h9uH
6mvXIJ2yMafm49EsahXI0ZCp3kUCCD41ia0u/QvNHU0N2Z2lPEm+pIsi1mzO+ZNt
Ww3veqqyZQ5lMQcTcbcl18GGK200OmwAMN/OK393oJV8DHom7T9SBCynFeC33VsA
B9jug0brx9IFwpC7YdPphphZjsIxS3bqdTrp2H/Ja1DMtc+4ZDG6VGwJhX3ksZHp
JXTe9TpHQ/HNo+Ly+0MWsJ0BaW3ZwVwBJ0whxlxsNvpjHbMFZkC9Ojo9kuVn+7st
ypCA9Qu5q71bNZi1PC3mOIfkW4ozVsF48Wsp2UFSRyRhaBqH4SsqzuVUdtdmAyaD
yyhC5/tP5p0TDKlWjtZSpm6q/Kzuv17DL+/OYBsRWtqzLh/ajdthSPMbXMYoydM8
sx6brHkgzDUEQyGQZTL5uKQYB1SWMCzA2DikrrYVK91TWxcBJNAR2QfQbSafpDKk
WWp2Bl80gsCq04B9F8LSNhtfaTMBgpVLjCyTErRBBQJdOd+lBejPtzR32LSOz9mv
8TL391qUASzYSr7rZ5RnLNcM0U7AAOBldoDbx18uZ9wNYIHA9P+RHU+70Y9lK9kR
NM4R1H3c5iSeGRWsjc8DYaEzopCORAThH+330q18ApXyl9cc+VXU0fmVMd5s487G
euIEzGFFRXudC/h70G1YK7uwLDOzcBdj4IFjMSpZn5oxyNpRulpylPH4+kSX0AZR
jlsYebv08gaewcXpHTLy2NA6EBNb0UoyiiILIaNDMKTzqd6t4WpsrJZtCPllKYWR
8C/P/MZ65x1ec1Hic7zEtCMNpupXRmE3pvc/tduOxBlnQvIEjr3HqPlztJiPtGyf
JdTUzJ5dzKHSYRGQTh/CXeiw2vbFqAqS9rsaa4Y++qocIzTE8mG34uEpZW4Hvjm3
hQLeCVmAwnYXzdeET0G0+WRx8YG4NTWTLozpylTjGfnanii05lByEJ6C8/24XDJa
Wom2JpeOU94s6UvK7CcpzOW8hHzatZDwOcr8jF76wJOJHbePEJ2hJfiAS61HmftH
Rsge8lLBSMxEfmmNYxFn0saOynrhbbQeyvB6KekV8g4ErL43ant8aLeUQJCZFEXS
ENwVYj2FnMCFf1Oq/1TEdsf0O+4ehJ1SLD82ioSzxiWuJcjAvurNK92AJLrRdSB2
KbSS2KwQwmtSN8iNsuAg5bsyFHVkHbdMXoxUu8i8R+K53o4lDJhR8/Na2rBU2xhn
8VsOhOl5kxwhI0j+rSxYF32BDgQogafmdfmcctNvXM4neTYnQjs40XWKQB9/WJQW
hcVtEthVzILY1AQ5OCXfJOMEEqQ9i0ZwRvMM2tSlzfFnAce1EeCd5OMgBB+sgQqa
aYoQ0rk11VH5M/ax+b+nxdnhGVRAsdRx71T7YUCe2G70l9TD7o01UgYVDUkXpFcv
vjOPR97tdOadXcAKXqBX2kIE9wQIIn2FNzkPRxcLi2+V2oNVc/uTtVy9nMtWFpUe
I/84+ugi6iF/Ujct8bQG6JKyY00L3Fo5Gh/u5GRSCB2HDUcgjp3n2V5znYHeL5xE
9qedpDUM6q5L6g9mozPCF9tzr/qZlhDE7zWOlfxSFaAvdT73mvs6WcPwEXJ5hUFz
gsyqDLzLeOG8j/WY2mCcCeHhTsLxW4XciIYnTmVCs8HPLKLKFDqhoKBilNT0TOPY
7WI9HGihtYCgw4s+T87pomLkeo5bLjs9usmrUrs23ek8YSo4CblIU09m9Eh6F6So
6LWj92slRVyNOVI/byapFxdHsxCHkRtX8nBYjHBPz2oY6sp7J7//DmZUpKkGBZ0M
N/Q45b8UaF4TG3ZMP7Q7jLCD50rQ0Cs5TJxEd5Nsbo0y2toM71FQhACzhHRGIlYN
vLoUMExTocJu2t870JmLKJGTFdq9/MbQ9C3RawJJqY99ebkr3qXkMf08WyUD0K12
b1UBGcA90UeiyeDQNnXYziB/EsQtvW0R8zuGIxNjXnVOwiX+so15uPce2n5L/Msy
prSnewIxiAgWaJQSK7Q2JGyOLTWGtgnJYWB+Io8ZPH6HZ8+erJFB0iMKhItsPubk
8EuK1ZXXbEa4YzRbQtsE4oVDFd06snswj/0yHZe749U10f2nepyaHBASr/R6u2WY
xs7SAVH+odAe8VIVTybkZvnIpQZDXucTsrkfoagElNWSiH2jAPTC5pVT4ewMCQkO
V3glq0/ffHeLxfFInvGysAHu49TF/jtl644BFjhXIm26gOtMMgpbBb/aSq6mfjQd
wPXmOEhP/kf7krZOnjcvDvyJWQaOd1vtF63VCTjmP6hikOa3FHikP6lrJtXeWUSZ
PNsbXirqkphCAlHWIPW6LmcZKyLVWeX066xW2Brg2bfSusooxRPNVkjeIV9wXfbA
NEXM6oerAra3nMCHPrtfgm7yiB6Nn882JfsBYAw2oTYWVOLPZoE+66VmJ+BcyxSa
LyfBWhRwPpjhoGR7LIjx0shxNlAJODGC3z/h7lMwET3O4/8M4evTg2zOPPNwvY/9
Ce6MFunmRqTY3U4tE5Mkv8pAVnyyDd0NWNof9RmdB1X+TOKZpYMghEqN+bsahIRM
zKDC+0LNEafITtL/A5nyX6PsYRw93g9n8CjQRrB1iP7fZrSW4mxQyw8sv1IvtEmP
dOjHFOrd4xYVuPkVJGOpf3U6EZ+IYwrADaGXT5dGnG9k9Y5gMtSpMXV8ttk2qDAm
yoD7edaFQOaI6/DQBjxv3L0agimHsDTsVax4O/Gckh7YNv2ogILGDl2ClmbBLC9H
78jjxOj2CfWJEjdtIsTjEfsexRHf2ZbBfuvO97HxIcF4G4Sd84Zc+hoRKEZ4PWvP
CU7GnDd3p2Lpc+hYBzBNeKBLisxx8o0x5qwIrq2PDZ/wA+eqIQOXRdpUot4aH4Kx
8IJC28rIxrVcdLbQY3cNA28NWrSPw+kL/dOE+qc43ulv9GOOSB1nU/Uiu7fP7a9n
iTcMFj7asJoABR7BmcYlTzi24RcOJQsfUprMFDw/RYlYhbssNC+fmNR1MYVeStKR
zMn1m7PQKmuwcRjwaCpCmSh8Xo6I0VtLkzTe7sHPKMnOTopSBha/Gp+iONGFe+gF
/dTluBfrXTs2EPS/r1Vi1YBxZgRFWZKW7LGJjcortBQAMY999Nh20R2gzmwK/4Us
vW98G/qXLNENelJE5fgSlCqWBPS6DLsmWzYxG92sJFh/ontdrbpmJSwkKnIerTp9
Js/8uc4sDTfeHyKiO3eouJN59A8rh7BPc7AK5nc59Bgx4RK1osOxWGbm6+7ZfAOM
WZsz1Rxtl1AWZ2sm5xRqTIipytVNZkKNI17mm3SBMkyIStRbk2RaKymiP3wR6/9t
wXnOJ0ypCbfPgQb4hnlMFkdvpU506ZLz4/9a1zbPjFrou0SFaQIg4dBVTThWMQwG
BsWnGxEsvgmh72nTR3qEUkwBGEibybYEfQ/mzS/c/lbuDBLqBZpAAWvN0S8yAg1t
UgIeuU8YqxVfI5WNPi97LQZybmN37MtKomSDPnLigmhpVNZfTF9Esgd8cR/OzFt3
vbq+VcL+N/PkraiG+/4oy878n8tTE/GDMUXDD8Q4L0WlcFBhMAhXIslHjbDicscl
UGSHF0WZVhVqTkaRWGoAZkradEASoOhmWDAIRxz+2sGRfQ6L/tRXLVe/QkFQp/N9
zzYulmBBqm1P/cw8eW1JIHvMz1dnFWqIPIMbwM2ce+QJrK52NuiK4c0NT41/iPMZ
j18zA/G+gCeB6R80yPIer33+waxGX1odcEmMyassPfmyo2iNSy713TQYM/lm4X/S
I8/vyzxLlfHAWn+s54V2dMTptTfeyE8DmGF+Vxjp1aN2HrgPwi6c+OWAGYzeB6IY
ydaj4RQriViPFx9RB57EheJuTSPokNC5pdCoRwsBLz6X9OF5h0cLAL8JkN4CT3Fn
gf+xeo/tqy0kcSoPzKDaSfUz6zZY677lUy2/qbRGxzEsCKw/2ARQ1kYgOLfA7i+y
ArbF1HddiE0rDce17AlZM43AgSX8LJk6CoCu8YIKGU/nWdtavBfmEVB9/YKwpuuQ
8PcneF9t1gE0tk7EZ9Bxdel4CsQO/6NEf0AviCBtQ1YXIYk8vpfVu8PN5a8vr3oX
y2CZRSLdf51TzRDR3lwfRsnsLFaeP4bTrMuDyIEzTJOSxdJTYi90BlaGlVnJK+IW
aVniDJdEVnhmYVx2yY4OqKFlY+sC0kbTOffxsy9W1+ILUSwzyuWs1U23dNUlGYbE
UPNWdZyX5tSrxx/I2ShW/PQ4XxAkENLfX2Chwgj4tKETXOfych2xoQfiF2+jaT+O
rS0OXOBysVW6hdD3FpMqFN5FzpuYNRITrNjQMkcEjs8uXGSyAYjbLbA5djJmFJSU
tAJFwdiCXi/o9wj36cJWAJHILbJKmalKahg20YFSUT9hH+TSdJGtAtchO/xIDREx
7+me9d7gNQNC5clntfQ85w6oLZWmzgNb2yHGUsTdENtBDUhHzLrOCL+JT6h6LJeS
TY/Fje4Y045uWnhSoF1E4a985QtX2DwOvVQge3qGXTOwCYCn+k46IL/1EMtX6TJo
FdO5oCwlpANh9ec60gcyz1m5aQQkMAHJyZSPTix6Q7zPctBaj7jHjUq3negjWVcO
+DPABttFf2R76Atk72CmwQIkOkDYAEzog+VRcT4HcwzIZBwmObUSulsFOMoVEtV5
oz2VunioXhEH3CSa0xrgiblAIzpWt5DxlVsyVoDTC3RuwuHFXuIo2MIzWUeNOpG+
6T3prdZeigdWaVsQfJUJl+3Q6HuhgLWZVNBznMuP/HNQLcI2Sd3gV1KP9Iyml30n
pXtMRMFt17dGypjTSSjbvy7atw6ctuR3/4xHlVO4ymRluNm7dz4bKDOx9iEhy8dB
tgEViDi08O1WAiWeFjjGm9wRHGL4UhK1Q+PkOc9KPpD0AuXV7XvhXGtrsrJ5fsCU
P9EW6lY8KeynkLDdbg42WffNIvS7oqwoeFWXSv5IWexZBvSWtSfaXmo3AHwpSbyr
vX59jxoPIRJbCgmCt5gKAbaODCQo521ia1yl/qK+JfIplP9afMh6tmjpFX/UEojs
a7W3Xcy5nfzAwotn57Ur8/oe1qf7vcGGCrOixtN7EB4EbBEIYsrPDJvv2G3KpfcW
WKxwBUlux54GzovZs6kC8UDHUhCt9T7cd0xUNySLz7D0LrAf0l8dZj8GtSusdq9s
jNkCNkXyNpi5ZtXNel0sGT8f4vvCUMrdaLtKnFg3L0QQCNqVe7bvMJPdSBx/d+Sz
omwD4JuTsBcxg51mKa3U2cZv8sSnWSjiwbPG/GospPC5uW15HkZIoClPSaDNOKay
8XwCSOjmU1FIkvlidIHKSsCHfX2pBJxmARBAAV1M0Fn9XbqhzeNs5QARVMoci1yo
KyHJHTDMeNKTSKznPBZSEXKQZt0ChfsV9M7Cu6g9MFT+S1PAeUICENWq4Pw0F4fa
JcFYovF/9arqueksAhsgeHnnCXjzmdTM4SLZH+PE0tHGCbW6KpAbOaf80R67ZiEr
TkH5plMMXmw5r6RyEvsQTE+ql15FZS/HK83O0DLQdx5DM8ojs27VVQEdZ3IfmbR8
BXW5ra6SwQw54n7vzSzH+eorAaN2GyttAYfipJ/oyfiSSR8mSKKDK3SzpfUS8DtF
wLOHA7Y6VI9Zifp+0PgDUXqUOIn1Stgul7/UmPmVYXJKwFYAiUromIpz4kHakMlc
nw5Hey+ynMsxmpC1fFp3wUzJRo/uGdZ2u2v3VyIaoHzoVR6lDkxevBSUK8rwUhfE
Jx0CpQAUIYOsf9QoduOpQmh7k0hPP9lxzxt+9VqRiyF0Q0vCjMZiNiszUIfSI8v6
ZvMhYflehtTQVe4R2hTAwdCdOtDT378+s066+gFN4p6ACRu5S+qiGujorKWAI66/
xFy+yARsqC0qd9PHeRQmDZhUFSuaNJkczufHaJTryxBFDz8ETuuIcEy5Bq/hIvyW
U6oJaafIFClvaxkXB8aCRnjIH/QgOG2XI54m0vrNfQSu1w8DOaZFEdWaI6XIqhIW
YqJRnbOo4nD8VZ7fuk/ulPUrosTcr3Tdq+pGrVNNvn5KZvLFR9o75jI8sq6GLzyh
Fz1/ZX8PJhCbY55AJiE105z1txq3cdEol1IsGfcw2wViMntxFJdjoHstvZyksJOC
8tN1HVtNyi1PGQ/4lMgeOdSAnQ0kmKYM5KL8Kw/Rie26OWpvdJf5NSKow3eov0Q4
2GTHKGeqKf0k26dCVbLz96jHOjLpRwFXUZl5C0MXp0OJT2dXezImR187xO9inkNg
URWdyD+gmVCX6GmFDBsM/AXAuCr3o5wC4EzUI8NbCimiVJs3iGC4AB47ayoMKAj7
bnhundFnVAn0cfphsgB97GCj9Z/IpOVobOjZzO+vN9q0Rw2BMNo7Fd/NQGNMxf4B
FOuGhDeyD/SXcQWA81Wrk7rJx7pzW2zmBde33OjY6KcommJiuj2qtdp+4Uq/AEkD
M8GwtYp8mdMG+HzrC+0SXALVrhuIwyHi/b0PX+JOitbIH7/oszUBvXuJnaOM2CuN
43rZu6CeXe3jhdEBLThe5VQi5OMGGFGaheqY7Ie/jSfoRNJkQFDu3dDC/OMMxqpp
Y7wgssJaz8M4T7UVnjbyLyADQN2DKJnepiJE6LNQo/bIVXuHXN9b8qjNsq8o70qw
/7zfuh12HDOIRr/royxI4+AU/dm4bL+zwprDXLBz26LQj8lffS/wxA11h4lETXO8
8ZP/qASZAugwrRCY4g4luzYGGlbjab6b6kHuCzRisJWY6WPu1AKRyNR/6nihWkck
xji3YrHfU+f22HzKl5c/OgcdwVqYmDtt7XL+3Z2O78pWL1yTJnr1p8gfPJG3RIKz
V/JD5SLa3RvKJMZ7Ot0iVO+RW82WOyfJbfsmgYhroBxvYwHGrimtZXNLSFt6ZlGc
QfwVo2kLlwpIEwqXM4HOKb+9t4B8/HH91j7NchiS8Ukki1DskbYhBHjL7Og/tHq9
5jKNChYHd/aWxRUxTOHuD0W2M/SHTqS7bwXvVNdiVZSuLpELeLZZIDRHckD1NzMd
aF00TdyjDUFf0Hw0juFBIFXGTKi5VqONlDKTuBEKUOupc0Wm2ooR8mQQOlXcR7o2
7wy8aO+mt2xVJq4lFXLOynHSi6LB3wU3AOnIM8EUZzRQrY4hejlEv6GgoznXFqDg
XKsYNhtEkMURJTS3rgf5TtDHejOaymcmjNH7OYrTGH/YOg5DK24fRZywk7E8mFOn
yWkGu4vhOpJETm+WcUkiz6/nH7oNHyK2BxSbuIXmGCLilPX4HyxTv2ETFT04hmuH
lTF8um32BER2uENMGwB5NDbRYJe5OhtgcRr4YpLNzxXrZFGaz329J/Xo5u0/L0yx
AZmRACFp4xMIo6iwjP5c1fPkkuWpc6heU4c5/NDYq9k84DImtVEZ+ZqLPkGK0noV
2KDYF0PbDEgSSc+0naI+NXRxbWuXVNB2grcYWCKMP3ZZ8sinTpQYXD9Y7azLGwE1
NcdrBnDqlXDt8U70ssBLHm4SxLxpGTOugnsr4Pl5vSgDHOTiyQhN95JUUBjvE5Q6
3V+FD38D6bhnD9LACtf9cdu0nI7uaGaue/w7XQrKG8aePxH15rWawJp7DRm4DFuR
5So3kKpzC37ctcW9CYP4Og+ZhOmK1yU5Xm5059gpRK/qbMsj08AGZXKJeQPSfIKD
dxwxTPuyGQFKyktEtmZpsfB5+e7Z5+7ncu5D96vttvDGFM9R0N2KR++rJVrGt5yN
uy0ECBypYYmPgtVWCLfyRlEK1DO12WZ+O6VtpzlL/w0/BkNqAVbrOTrKpL6X3UCR
CYZdzgcqa1RRsolzGGllQlz0I8iEBeTWjk8D0F+LMXqp8ippAshP66yXEXTMSx0w
ZLgxGomh0iJoRgScNLyXCMu/Y+2mV4123DE8qovBQ94Ms7uhrzfr7VkpTgIVTjdw
z3MWX6Cocl35A+T7+/FYE2JhpwIqA+sNeQSPm8jKA+J1OaC1+24l6fErOFh+PcKI
UcHBdx+S0WBXjBiW7K0Te76F0lL31Kgcp3o5yaw19+HeauLHi5xlxEuoYsOtCnGM
FRc/ONXch4qB2GvFNqb5KjxS5sRh6dZM50mO0ATEKegq0WfduVm4mX97tvggm+VS
GxnjmACBzu2ilg4/hvPzfZbdE3P5Na+v9vlqcFVTB99NvgaZMcHm63+ZSZ5K/QkF
Zc4pRH49HBK/ZgzKNELaDypynHyweyD39mApXeof+h6ilZkHxbGuL5XpdroEc37A
BRKMh7YhL56lykl9Ab+2P62RWv3wJGogPe95+XXlnracOVXdTeAuSMrBbxW3ZQh8
u5Jw4YxnBbsqGO4gejAZU7+XvA8ioFFJAVc8DUWaQbHyTYVbc9ThcSFEACQTtNuu
xxT6N4d65y8+PpZJk3bV1jELVWMLJtI/yJjr8ajP3kwP3HQzfMIYxAriEutKhYBE
My7acTF60eePTGzeiUuqwDKsfoNlUMBuCyuT2Q+vQnNCxs4N5yXneF6q/ZLYjv3q
NArjbssVy1YUsxycFjtmwjCIZ9lB8LiUF1+Fhgg6hwGIhOmHdjpxExP4iOlmQlD8
AgVo3ivfYBR4LfBWpfAV7CkqVxDiu9/uU8195CwYU8tQ/AuA88+Myaeve1zf7URv
3rjU5eFiCRWyYj+GkSoHeocU908dXU/0Mdj9N0fwBfIHHEzfYlfiXhon6hTZdt6u
WUGuUVd5mgE8yVkMKN5wQVpGc/eMjVmZiym78HjBRskfcfOrE13VVgZai3QtKBxT
CExPdA2Cick4cEniCTn1FvC5n4GWVv52yK6WUyyAWX+N2zOnLlBgwSsCbl0O+xe2
neduLGmsAGLLVC3VapWJFNycWGS8rHhaiIgI27xJuiGEXEsT47em5CF5RcwuWjU8
bIeJmG8zEuApyiabZ/9l0mu6m/pW/UOwNnfqP0zLqMyesEoIOp3fAnK0Q0Ika7NC
L5gbF6qqO9d5WCQy/J61DYmrizsUaJaGLdwCrSXvX8Bs1q+C6EBtX4cPMCjcuBvq
htwAgYpvWzKffTpBZDLMkyQKMJHYFezs3sduGzB60eRLnvNEKoyW6ogihlOLcHPN
OPL688OoE+aGgETgBJ3GEOXJW6Y1lpqRevo5WdoEBvDILOqJPrVuutsm/xu3JNY1
ZkCd0s7p1hv4rRSjLxr4MrUakaJFmVS6ibFTycsDB8zhPYTfDxceXhJ2qHvprBzk
BKYxyAbXSkgqXP0Uscr8G3STqzx4aVZc0khHrSDiOV+4owHfJShPs9zSxTvaapWV
rLdzugWBBDB6LuGw1f4FQDdLD6km1YymYbwQ1JuGkpQdJYmkStemNYxu23ZgrjRC
+5J7zkceCtIn0y66rmMj8nFuY9mv87NpNrNN3ElJ8mU6C1al523kaIDYRVoAPJos
9U+V6wpUBxTMN4P6OSG4L54eHeAji8JqbnURZ9am9kdGx9TAYClbVU9FD1u/5agC
JrHu5hnc4uLGyhqeaOak5dnYwA7cvNjdI55n3CsBMNw5IRZ5Hc/VSbXFOzNQz650
rgWNZFsSgWHlZ2D/BBwFmeRT/cKZiYu9qd1JHEdCmqTjfjU+fJnWVcG5P3Kqii/C
1kn3mrOVLzgKEJ9mpX3vGy6adlEDBh4dQ1nmxvC+mmBBfAB+ntlRhWlq0YhGbsgs
McJ8TMMA6Cb4rDjvsmgALGdpcJ2CzQ4ti/PGPiQWJuZYB3iniiQ32Lq+gjBo57ch
yHScE2On7ZUXEyNrZlX0/7PMZDI/A7/+SNJrdsR+1Ug1CvVs0lk2oXrO5/9AUktP
OFnwtAp9WcqdEV7EnzpUppi5+0dGEX0l+pKEDuYKbSNEfJ3rHvHX2zFN/wDcV+xP
vtYyckN3x6kkcj2Dj3ubP00EPAGM1XT/3p5cZUrZz49bwkBWiF7BKq4LPRdyzTT7
OWujjL1SmX8ZQQLWgwol/uWWgA4JTviPUYLjRe5/fVZv0OHe4MNT9FqRHnYTru5R
PVrRuvEtxmmFawAj7MGYw2tKETjn7p3B8j2RyVsl9Zy1gB/Ez25jZTp/w1lU6XP+
AE8ovtsi1UYDJUu9Z5eH6Gqep4IqYPJIJtcZNw3QhDQvJ4L3amvL0L/W50YzxL8h
6p09tsqat2BT5RgDm49Qy8kubQYn8TAojjiFlovukevC5OmtLTfzu4DdDY6x0iW7
LwxVkmGYjDkYDYmGBhUHbtp6WY8yKw62Ad5rxs/YaSQpXr8nSBfcBSI/+D0gUXVK
mVJINp48s6pBTR5+MsqmjSG7Aivce7VGFHEmYfoWzsOTzduVAgG3WOz/T+qJW35k
KOvDFzlQr/fQwo6caX/pRd2ZCKhe+3ZsNGEKl8ZPXnBV8FYZ4hJ3NRu8fYxbG4t0
NCF2TDIP3NUOCL/lafCJ+fFAcpIyN71Qo320jD3jsPgyFXVzIdo4kUd8ihit/GJx
7UfVrsMUGV1Dk+Ha/SvtZzPCC9Rsroq+7d18CtsXg6xad09+TD58EQIZt3bVhU5J
qnKmoGSmcaimUyr3tS/GJmI36GvfC+RyOA/o0kG/crzcooMjd/xIT2E8k+jyVlmc
9lcCL9JgesGlKgqbZw9VSJAZg75b1UUZx7L4EOqSlz++sJpEj+cz5/Oso8kr71Mn
D1dqKJpWOewGZfIkk6atLjZEcKkfrEVnqci4ZuONvcYewUEkhezoZP3zwdiAR0gZ
Hx+6TBZeeuRHma+elWZgIfylOkSyjR0UAm2zVgxDmRb4eww/P+FJgn++8PGbB2oc
/ugM9X+vM/xVFXKXUGZ+6yAYbFaCL7JJ1c5UVrpzuy8aBq5Jkip9HcSdIwq/QlsT
C7eOU80I6GdP3Y+e2AECSRZmwTutV+jqzQd/Fvs8THcwZkuzmPpI4FTyHm8G4dG5
vFIFWVGZra4L9Dn7usQ0+NT/gQil2QLnBsdYbeOg2RDwkwReC4NqkA6gQ4P27Jwc
wgPON+Q5de0TskYZu56HkRGYXiUBspSncW9+5tAmre7TT5Aj471VOWioZZbNtJGI
N+HAnWmaJqJ6CSVL9+pmXoUF/4VXdvqYAcAXomR2RgQi2eqtcZET3w7JYs5zBZ9l
na4sYo8JVVRrnspR659vOWyCB2R449nDGofGiafK1B4ar/F8JuYg+jDLKXuDuqFT
HBQR2aDpSSUGOPuYX/+ypB2LEizbzwTULCsWTVx0KtuWXHNUx02sv8afJi/VoBuA
5Y1OZ1NXx9g1tdlCUDo4LWwz8og5/cS3bdDXTOYXGVaKmeX45ovTndJ/7/DY+Tlx
cgeD8UOKMRyPVKJ+yza+kHzYgFAqPvMG4KSdobQEpq3DOgz7IO36zEbEOFS5KtuF
JGttqEK5Ujb3qlqmgRSTHyYoHSCd08DrDNiGpj0wVJETGA9IoA1B7eYdhEWL4LhM
LpLw0IjjcroqZwXR/vaiAEqRF9P7Ajaw60HhNGtLcg3advh5kfHvAiHYZAvGxS2u
rRZBA/aa+u9rg1rG36slWGGEEqINgdBELKglZBM7auZRc0dhLSkqz7kBA8Z7FHNg
9aadbcyVf6mLZvRIzzks55KJknneWiuNK5T7ZHGEvFON2XQDW2lgD807ftzip/+c
TrJonFputIWzQoSQhirqO20yq3LjxxHMdOyEE/0+GuTfUYLXvglmd7ZHyjEXVSpC
KPEKtkYo6LSmb14AsNF8BdEOQe85hRU1D8bzbQYZK2goW23nN2aIJOHzV1ApCeLz
IWI1ukJ/BJEf6QrKUSZn4fG0hof0L0XCXdYpX0zChIiDYtDCrP+r5PmH9E1Zx6st
R3LBWrizYD8UbI6TY6ihge3HYw2v4ScV1YT9RKQ3vQV599pLHDSUdZQqAlKVhx3o
eH8gjLF3H7Q52xKf1cSmj4OtbkTLYgxBOM+ngVK8eABZC1fi/fKvnX7JAKsV9pbx
HXPxuhVB+4Be6S0HZV/0CmdpDW1YfoM+w8eyE5pjjuGK2T79EThwv8pVJkjZK39/
Fl7lrrtV33EohsPrVc31LHfYh61UyhIeTf7nZRD0lFw+/evk3H4bgLlPtMwBijoM
JAxuXRpuEZXqFYa/2ceiALKDBoXf1C/6RMFgrG6yPatztUM5PuCkrWiDGfA2cri2
mMXmj5I7Acfn648hecg997NSXzWIKRpSX+5DiXnKepb+lFbLk+dkBNd9Bj7PNyLP
xrUhhTO7Xi6kuuTZz+H4wP4nu3wDCLwz6+/EBE9BvS8vFzhMP9e0keAZ4Mg5zbnx
OVlZJjot4ErLlpNarQe7WccQN1TbTfUWz8ButHKg2m5wbj2r9bPGCfhp8wvIlM5S
J/tXxT4HJz5Kb6eqj9zG3KUAfWpulVQU9L5HPIFuFNXU+L28yRad2CV04631aMDP
fckVDVM0miYKRN+3hTMXt50b17kgvZ7iyGbZPbpPyDp0fPtFQEoEAkzh2yVyU1pE
BjB5EXxpR1V+HD0kQ31gZ4xcFbQNPC9okanGk3jmc0LPCdWGjHew5rS9YSuBrREf
XDJQwzXc2jQ6iuh/oTybqYkRKe/hK5HmmqRtHOCypg+/wywubzZZSQO2Q54jHYys
enVx/uoUM7xezkSKotx08xVrFGW+RiSU5l36hWRz2lJeYM7gTC0CPssJRor6sWXW
WiDYnxZoI4tHiamvzbFoMZUYYZxRZVpxQKnsi+21hb3Y4TDIEqazEDQwx4BGK6od
TBO4B9jEmLIY0O4PFLQmaZy9hdeH96bKc8xCK5m1bqdHqoO30u1MkmsaWDZXLnwh
DrmZ9tvAyCQr4yD12tJjwHC5Sh6zfYsh41U4N4QcWKp30Nlt942qdqaO0v1MWFBp
brHHiWgTLtceB4FdLiQrftnVs6Yj6ujGNSU9BL8lIcispSCeLLWUTrHM53XEO9qW
zwkSQIc4cqEqiBm63F9EBxaiiZ5MRFe1vXJv3og9fabcex8Dp39nDpZdHYUgsv0I
qHgSRD3dPKqJHFjtdfzHCH5OLlOB52dKdVgUiOT97k0Mtz7NBKQLSylzUvf3bWHs
390bfl0IyoJr31xGGt9B0FvTQpKe/ePU6vEz5zwUrJiTUnqQX0kKcQGvJRcRywGL
KCo63y5HoUffufkvjiUEF7re7X+Ruf6AfXrbmVohjh8KgzA5lk8GX8bbSsUodShx
APBJxw0yD0UT6pXEiXbVeN1530ylo5tbDf9wrrcwK7qQWSPiEx7raCjZIc6nqazP
Ux6gDei9cmV1zsFtiCaazHv+EWWgOAw0S84csXt5qTtsTixdtj1ZHbGS+/fryqtV
HiBYpepCdpZpQ63dHJyO5D3EsTTUXEk5mA/I3uTEJQSg+HlvOQ4wGgT/mWb0gfIt
4EZi4CNhx4bx/AeshHlnQIUNPSgnUJEoFHSZwnpS4z+GYk+wau3Glqa/mrO3WliH
+BqHsLV0LcWC7eQgg0YrhT2HrqwzbX6XFfsBa4gKrARMuIUc2xgFq3l4jGYbX0Ht
euH188WoaRc+bOzt9Kn2mEEBsqG8Qu71/U5Tf6ro+Qs9QyRcjcmyvYOPKY+sOeKW
zz99DGTIn15Rd2Mq1NVslP7aswptKvjn+J8omCb7QQHiSnnYN1rygNKRcDw8bG3K
bMr3muVdt6yd7ogMIOis7SKUSFq/PwK2SGeYBF4zftYqpiLIbOOc3TyxU6bqG7Ns
cJ5Bdtm48L808N5Eguxg7gy2TpaSna/xkr/bDyu+RsRGhqZVNrMlTi8/pjWxEzh8
uFVbmyOiXuDuGSV0S/KzLPgjoSbQLJ5EQ4loe/e0zrbFZRdu76u+VCFNO2wen+DD
hOeMc1K7+U6UIMqZJ3dan3bz3IDvkNpSx426uLXRjkYvDqJK5WtnzAD3lQkWPp85
7oJ1DYC8g8a0nCQPwZKmMY1DTY+aUOSNBrIBuGsg8ew68vcJkTSFjvTJ0p+4PZn6
GId3USYp4L00mdgW+revkpuZguBa98Ev3Xl0eiLQmS+hOuqqg/qB5xqadF4cj/f0
dkb/OHkPwtPzg56nXix2M+ql/OnIsNfR2xlKdlcCig76WkRwAFeBrz2kQf16mgqd
UCRXD7IKEihLKoK+7svB7UMSbbSwOQP0RVga5frx5hzZ8B6N6dP4bQ9DdXauULYh
PZRiiZnTniePHVUVpIraKgZ3ARR1YsBr9AKOAh53J8LZssBFRddoq+p2l6HGmI9k
OzgpuDm+VjoTx9mHpej+KW9fp0suAqk2P1aiS8jUnpuQXB7LKo1+mc52w9GhdhUO
/YMwzu8TnC6Ok9fM5og9B5wp7l9LmWr3e8gfKT9ObkrxU+XP3OSghb4BcChm/n+a
eBfOZWRv3Jg3UqLw3Ls4MYzKbRFT8DVZwP+oz9CvCTnqMvfExi5gwfnnf7lrxpgD
ahijEsRVnixGcBWyrglChMkAQ+Mn8TTXgCco2pFBbVqNhdAMAmu2GtPkMQ64b6ln
jIfXoxhqk9Vw/arXShtzrGNqWNCLOZID9PULG/e1VB1VRWdTYlrQCrKTcTtszOEG
tphYfx54P9el6kGdRCocPTXwlvT3YkJ3facsUxxu1beCnzicDc8MNRWjSrvdgI1+
/On7HUlNacNUKUjQi6bEJ15qLPWAD+CSCzBSqPdXCotuQhH/Gw+o6u/ad/3xt9En
jnsnu2l1ZXH+5qqTSngl/tjUTKcbSGVCqFHxUqqMlG8QA/q7o3ONext/Y+N6mNFe
jKZN0+sZsHas1LQSGd0nveiHxYbsAoWBZ6n4GVIXiHjdgrzyDgCLZsbGZf52Z1z6
16wzjZgo9fODDaoPttzZwG87zNtFB+TZSH1Ry3xQ0Pp8H9yvUHZD/Dp7U41awQi+
yg4KW2zrxjio+PaR9DG7myA99e8u7X/fCPjTkojFwpP/I4CM1A/5Fzmrh3pDTIR8
MFhjWbRiq9YjDKKyZuaMOX+paPibHzSOW6BzGMceLIzLcpqnMcj4eIK2HkcBD/Ri
eK1pP9o9/0iSft5TY9hbGo65DpE29BdCmc0xZnJ/byxpqcgu7fvrvyoc4uVmOVeM
GHrvSW+6LCNTxkz5QpYNM5gQxzgWOuAWLrm198To4YWUTp8RGNYwWARUBK8cDNi8
NYMyhNVaR5ghVfXG2vqYKf8WgHOxwv36j4WYHYdrN5BmaXHXJbw8HovqrJhPgSIZ
FxWEm5E2jAAq5XMdznCmHX4b4LVb4JqTPjcPfIKdclDo53DJKgDgjRpZFRr4fZcM
O1O5VXpFq7kmeoRR8lGUBuAYCodRliuvgG8l3c85QZ0H8q5/WhTk2rZ2lKsg1Y18
R95+y2V+clAS7o09B9KSz4Pb3yKX8TIpwaiCXUYq+Mp280Fb3pDr2aWRdphJMitx
tIg25el+UX7FuSvdRuSueqoNS/m/6CG22g/Vv2GpYG8OdA4wn4b3neBUY07oDZI8
tBgEsmFK3rfdRlMIYrxOMVvUoDvW6riJYMC6pi/AKqH5SkMLg8AyMvGnK7+eJtKo
c0HHjemKeAbGwzzAvwBl7P1fT3O/1sZVCuiJEPQfflql+8s8+m/odhJtA7UpmLhY
daL7hWQdtl0g2B/zqOpffbVmJNbPoE40j/pEYcIgZ58AxL+oNt1sEGiWTola1ERn
oZTuGd1Pvtu895G4zwiGLYRktwPeReRjmVU7aTml02NOWu6Vpx87o31mfqCU033Q
lRalxk8h/1RSH0I6yrmhotD47aidyGC5/Y0w9nkj4pswtkkmLa92iu7cVQN34mg3
NrVkip0/wgtDjjI1Whij/gg7vT9i1gje/F8CaRUYz/HINSd42lPS4XkSsIzctlBo
811OvkLy3RoycHNHU/zb4KL5tzs5vJb6vCQ51MAXOV/MbcKJKGc9NoKBHQQ7cBTW
ru+Lm7GuVco3b7JUPPF5KIKOWpwQzM87UnVBMphA8mh6TL5vb3SbEaLJZwhadu/B
v1L1/29OlGAE1xJcirv6tNujJ4tpft5QxUmu8SaS2c2eX3C7HYwHDIACy8tUnI34
WqlxgK8+uLoUnwPoo4YNy7fSSaj1Vtusq2UEyrlgdKq5oUmhLruCL2ivw130ebWw
0YVBo7Kn8OBxkgV3MErkr8tjM9TER4Nox3EXE6Hy9FjomYXf8DKnDP2tk3HU8tNk
ZvpcNez8GkrNLH1KADW4VHEfh8DSxQMOIP5ea4fsXG27rg2eF+qsISVngewciX4b
ZLtwIjRGDDMao7ljtepeiXVr17pLkc2r2loPcRM8tGpbnKBd8quRcOzbx5jsgNeE
U/CrGu3udvgTb4F9cOolCQbObgLCMYOpL3SyfxuCsMCEAMtQ8Qko1mArunAmEtF0
0s/G+3W6VaX6vjyl7r5DiJf0hz19nUccWKCmottQCs/AktaQefQk9DsXYWHvHb8J
P6yD4vj+47kvVhiobry45SpZbgbejxfpqSoxG53GVgmGnURS3a02xjaYOvKJZHgr
qZ/oYSpp4ZPiMm64TK796PQkJCnYoHV5y3zq9bGyCmiydMmQZbI3jwsQs2aYTQE7
uf8rA6n5pHY6ERXYSfwlQRYXoCkhXjdkddnwnAoKsrEGQB9wOLn8OETGnJHtiItT
3ZjkCCCam2N1V3iZhVGcejoBumUMMTDzO+Duu2LXad5im2mYjjqd5wFDI1+AsS93
KAj50IMgGgS510i83W8qDHdeWdu5mZNB74oh1zjobblDOlyc2orMDYsAprkK3Lbw
VhsfF7o3sZLrCGFAvf/Wgcu4dAjn1R0VBGCWFjEOmqwpBybz1g6ay/iwqk6Qg+N/
x16VPvRc2eEhWY1A6h1wQ4Gho71hei4Da3KxjI+hp6UpQ9WHEAp5cXlr0KbIY6gC
nERVJkgYpnSDjw5qbrDj9m+NQ84rJYK2weGa5C6Cyx/hXX81AFOMOp8BIBVzSz9P
dgebxYs28nz8Wch6hc+1yVtkvDKXsoiQgyjJ1XdrL4Ko8RKM8addswrisFHuZxvz
v/pBGWxE9c8ZWpo22VlHuGGz9tQXC/28qV6ijOoSMiBZOVR3ivhZJQ43u2lF5GVq
mh2bOYRDJyGzaMWzgMA4shruIvLFLC8v0kKMjXQ2p1VIvlv54R2ptnxb5XJCoJsE
ll9qyXlr5JsEqX+dLo14Wczic8Rj5agiORF5siqO8M52Xq1C7DN4FZrGpivGrVyN
GtLfHxdBlCUCXTDG5BAuwHy5XoqGjIUrvTmtjTrk0PJ/OfP3Fpt/UbZRINQgL1VX
dj1A3o/R31E9zNAn+4SmYcjtiMBPQupOpjhBg9gpfqXkZpuc66e6NqpTz2WsPVsZ
eZ7FJjI/DLuPG5SsSOYhGLwZN9RjZu76hpsB4i5EaLay60xIS5PlTbnu6bl2M1EL
Cvig0qAYMAvgqawQmFrOAewdS92x1auqHaMYT4vux+cPl3tbyfQv9ijQGdEqiO7c
XgFzugt62ygS3VKBt0qK/fRsVyNlTk64DYe0rD2Wdl+xqzDc923zsVl6QozD4oXz
57hgzN8cEbuV4bmqTepr1hfBBweq9KNvwqJpTQIg9Xiw2MHZ5fJs+z64haGyEbV7
spUhlah5cOup+i6bwxzffcnaho2fCRr+r3tfny6tGEZUMoJqlmZ//4r6Aw1L4659
0GwLvqltqtZ1rtYDZ03wx4+C3GGi29DdK5o1hYNfaD2lZWAkttQsO3ZhEYiDWoyn
37LrIpyOZy0P3ge73u1wDTzrO3DjhtBY12iwr9rEy0u2IT2vR9XMIOW9Cf9TT8zf
r+ivGbY7Acm4rYMgTMBRtK1OLOr++0gusW0qZPwcGmJsyFuEbBc/ZPc0bBI6kLLc
Dt985MWDvXxJG16Twkn1kQc+YVPC2vk9MZOqhOzFGyOFZdtjajEJNTOov9/QNsJF
TMP+IAKzFjGGU4HgcabxUS3DMVtwk0QEx5ZSpwyHbyVkUjvTiUa9gNzYZHtfGV1E
pFmrDBbW7Qh+GFuTiK2HVxTKGGfZ1mXiT5g9tSS0i5Ru6tZHkQ/2J1FzaBtUHItp
/v172pJZWPc/PC7vMIorB0I+gWu6CgrCeou5RL8847SemR72ze0BA83CnjxAsvhT
dPnNnnSdz6pv1RJWC+XmV9jxvmGX+97EeXaEsX1fqfRMqWFDPuWf5in49pE0iS/S
A+DzPvOHpif+PBMVuwYAMT11oKy/esq30ojb/kigX8Chq1QzuvJzqEp+0dkxXxY2
WkRMdYCLnrtSOUsJzYPJFbYkyKqF059aR9ue5ct/Kj7KsWplDBNfjSlVSYLfxe52
CJpuzjZpqUgs6dV7xNt8VuHP9B95n1V6e/B12WS/SvgNQiYxHBO7WyKzvHfB9r+e
m+efmFam7hZZqQ8SW0Y5rvsl2/zPBCAQT6MY5gsyuote5JVnUfjGHjxNPhqrGIUa
pbYqpT6z5zXkxRveDp2sUJhYBxxqLSQ51uA2n0jfxZ61cml/YCBJzSNQi0Jcou6V
UxP5OL7ra7BcCJcZcwu+iGUOnKQ5iuDK4N06A94KyVdgrEtd0DtSJi1zzqH636am
iNyH8nqZig4VlJhxbfPADBiKZzaCNqhChq1+fpBWJUDoqyFtTOkBpN7+udPh8DjW
gqmv5s0R7cjmrZzGiYl2Qh3eXO72+3bboqa8WlNmPA/iGJUUuN7xft3weLnrIc9m
mqWITCwT5hRCxLqPx4A0MG3Bbe1u9aUyIKzepelkAKS0f2fBsMdEnlDq+vzoFh/X
014IdCSGGn4cAkiLOPPHmvYhod43JkEw+VKR45l9Lo9ileeKoVRj57CQqyDyj1Ax
BXpDv9nhBiGAanfgyUb6+8Nu55AX44ptLL2VgWTLTXxpfd6WKq/Ld9BFRoXkeIjg
j30J4+E4es8Zae5xG2rOXdjEovmp6uBBmOdqTDIXhEz7cXrocG3tbZNrAaRAXq5d
04JFzkdPY69FhTlSI11w4JjeHm1OXPmzs3jNWla9oNGJT1YApmxHqXdxgft1WaB9
xVJjjCdKmHMfa6DXYdv+wtE+yyGtTGcNdVKlUbS2UPAovNwlaSD7lsDk/hlp69q8
zUG3qAqZgqDF9b4QoOUbDapkN7pN73LlYyVRRekNnjrorz0B6sfZ92IUfQNNxhyn
+1+Ae7K4g5HbUQGSMKbHgA7XMXaqYmi3e/DTUOwVA3aH261AsmC3QFZLxnap07G9
uMX0YMG7BYWsNNCD/BAKExwFAL9JWFXzG0YXkuFdzIRuhXXMWgPLDV6kj0aIzr28
QkOLD5iDPH5GIr7dYn+ZZu3xVWhClsfPZ0zpBlh4z6njgqx/KLU9nt5puDzof/4M
mnTPDu9+JR2uf9RMM1Ae0wLe/QWauCOUkwWLrZgcP9FvVjoFJWuarmMQeu2u9G0r
xzR5CntBEszrzCi357gM18ljtwb0virKtIL/LNDMStIVO5qS24MeEX5rPUKeP4Sk
5YlbvHuutMX0Jqcg2hKuV0osbth2AAOhIsW5NqZL5FW8ZTXPogXoHUde4iJrS/do
aMrcLYQldiYPjnh+vhi4MeQHOaPwz/LiOOMGsY/4XDx5SocACnMXrgMjR8xnfsXB
UvIEGs0Xjgk8U85QX3sBNotsnx3KY9wDDlr/n1D8niVv/LVjTqdVV1h/ithRSZOY
uU6Eqh2M5uqg5tMMI1XO0vBPGgecyE8qLPsTBI7zL1LQs7B1ysw8rBJkie3Iuq9q
Kru8rKVlG1P3kaup5rQZ6TIuDKiFOcp/q/sewK5jfIiiQ0oujtfj1OI1QCB6FX46
Byzj6NYYqjVU+PCg+wPs41sJ9Nq3ZyxzGkU/ljtAXr15VJhftC4u/JoCUr+8hPVB
SLkYNsjdZb9UOnixum7ilH9jibp488yco6AMGppBHhxBJMtZheb+kCjAC6gotN0F
YQqxXLov4aPP2n5p/kPCM6u9qo2mQFWYvTNdj3UtHz4gHY/cs6jYn7m75Nat8L+q
iduTdgIAD8sO82KhHOOJWHOnhRU9zKMHJOYhvn1bJjVKi4ZILd7ZcuTol3tDLa5F
iPlOJTxDpbhwFrqQauUf9h7sYY/+BiXx5gF1PEBdKeCGEHs8bCL3YcJ3sQvN1OLK
5BBn3bhrr8yHNOViHZL3IP1ud0WZooEgJnv4w7kt8HcYAXMepFWK6s7iUDb3q5B9
Qdx05Xw3hPfq9NMtWYbZnEpMqYA3RWsTqEqIXFB/TiMQJEw7XEraP+NIiQ4ut+1C
EB1/lC1Wq5ZgwjxbQgjP+raoSgABzqL+6L2qhNs2BUI05R+YfLbhEFIRxD0O8KUm
vozIoRH4MI9Qbwx9J3MAe8B7tuZLjv6rIxnmvChbsEsuhCIKllXbZ8NXiOttC1un
tRqmQ8nmzlmX5DTnbdY1+CSooA+mhKZ/z8BoWQigmfsWQIT7qqqmHk897KhyaP1k
l7fC/O25i2GFqbk5TlMFDxc9Oy+stpClGkMbH1OJdOOr9Dq11ngeZ+Az8wCEcLHn
tuMOd1ypLB9OfCKcBQIo6xuLEJWL/VGwhLLDUMrpoV/a2P5OaxPDAd4OnGBGULL0
kqmIdxys51dpXEZlZb413g+t4m/SWgSkoRA2rIFYDAZ4Q5aVTPqkrjCrSbePA4gw
z/FLxRsyeNd/f+UWPNUj+e2+Z3cMoyWZFvCNT8jqTkeSzfSeBkRa2pXXxMji9LaL
3DOdjoP23T4YJMAJsVAvhLPfO+PFGVjQBFCVQU3/dXvowcUI/UfqVYO7Zu/HZeI2
VN2MyT9KlFHEiYbTlRj94Js5v9qQ7HpBugOSXz+P4pPMydO3VJrG5h87ILmB+wk9
W0RAJGjTpBfrUF0n2RiQWHXowalzGQeBt20AVhx/zXhUDprnRS9f4IcuAoOm0Vfn
c42HFXlpzDqjMOYDBfOzq6jXz20W7KLvggc/BUfgpo0drmO5drDhBbUKE3tGazmF
pJU75YKXKQCyMDsjyn8CUakSRnI125JpDwYZnMyuHU8lL5m3uTf4HcQdTsrjCvFR
Dnut5ZVCvhFnNB0hlYqRkjlVGk5xQzxIYJk714rZw/C6Zk0Y+ds6uGaYiC6cSdqb
q6uyYATZlpzqhXP8kOzesMG3YZ5+8lgrBI1ENdUECllQKUyDH7xLl1+s5tsGhh+M
mzceFO4RfUmGF18OtqmJXZXCLUHPK8NnG3u8ITVZfAIkFJ55NI/aE/OEYRMvclu+
bBV3GinNNY1JnguKLt1I8SYfXTIn47TNUXr2mcFOWsjZ9ZAP7EIufbSQYYB30HTj
jVrtmrx5co51I2UCHwEeEnhPnnsYe3ao980rTrIjSQZTZmtRXrWiBNcKuBBO7YOr
sGIcQqUGLOp/0mSQ9GMhkebxVHOhbsNoHb5Dm8wZwNJ+0Rwoufh/x9MA8qyOLpXG
+5hfPX7crHtNFomzh7lOJ9xxMi2yHDvcceiHAvEy3ktU4cDMq5viH8CUkhREcLrB
SYsYeCFIxQsOlXLgT87DJ3OWDIe9LyT/JEmJKvT3x10uZhJEN0u+X6rJDihDLlkt
0BG3rHqjmFYMklsPuNa+jpeIOOtJRiBnOVKiq5p8exiCk4lo10kX4Ey2wEL24PZK
B9ENPGcUOguc5SlfgspxWQi371b/xt0/LolifklIx30+ku8VYlAttErTSJV1Ghnr
9nZ+h3+/7/xJsZcx6uIEhcshHr8M1wMOS6oyxoJlL2jCzDmxw6Ka68w+HHtqd30g
Jz5kyPUSb9KiT/q+CZJFuwMDjs09CVUOt95KUa3bEzxTOrcyBepZk3s0z1ORQGGf
PnMrhDG5LTqQRIRSwqacrFScXMw4PSDjg7SpYwagwN13+LxkNbU7Gt36at0P+vyN
NZWtruu8shBkeZdtX6YT1E7o3FGrPXMAXK41DXB2mhCBrdR96LF9sFpLpP3nPOFn
Jm/pWmWFa7a3FQH3GFFBSV9p8G6ee/b/QxFm9GbeHk/pYEyYKW7VvYeqThQtA8rf
r3djE4Ff+tO5VjHLyf1UEZrPaTlwpy08C6EaVKbGrOcqzi6sd3DDrocYYWtDB7vA
3uDgrsfipgNDijbMPz8kcGhRQZ1mDRBGZVO14y5NBLrfDfNOmKcmxFVd0NsOaqxj
EuMqV0sbxvE893uOShpbOz7pWsGAoh1UI6j8qhQB7gK5ySuB96D1+B7gL0z2YMLq
qbdYjv09xen4XKIVLkj6twXMv2F+jqHqTVkOWi0yFkK5/GSCy/zKckWDWpZnO982
7nxvzIr6LZXAUoOG+EPKg6F5Q3RDSFUJDPNhYX7scsJBpDc/CNQ/DnGCn7uRnYQT
qFpQoGXjgnj7YCZBIY0egdLr25GXS1KYWXgzj6F2x8iCI1+0VJqsSZEqg/D8wq2z
jzQnAJnVQeNnocqW3QDWDM2pFmAGRk1CskY4Hh1L46VlIBRYGgH1ZqONSTQnaza4
qXTAeRftDQWgl4WWVnstJbEv1yXxwdYUGjZBTf7vRQCloayxTN0lvnfPq6YX0gIT
UnmVx1jt6jPQa5HBpKyJ7tqpCyHX/+B/GKQ2DazBre+54uW815cRAwMP3GhzV9+M
xjAQkFPXq0fkFD1t9UqJC+JXtIzeIiojifQvh+F8c7xeq4AnQm9DKvp+CMr2w6LF
76x8x3OEB315gZiglCf5jWBsLdeX74gmhO3+OustKMr0F1jCxQOBFjjqm/QoKK2n
W6aiaL6+y4JcjpWZgaiGIon6nBbbJ3vbJL5BKtzIOAa0+C8Wg4/TsI9/L+T9Nfsr
9Xj8bPYNjekTwvCnHlVjNgOFZBILeYyOI1nhbtqW3Ysq6Z/obhLwKX2Q8HJDbuc/
8gD3/Y3yd6WQwNf56rU6/ZAJFgYFaYqqFslBTnEI3xWDGkrgesHU571SqadJXBRX
IyMN90cIP49zokTG+K+aLVjZurM6dTRmnJOTqPf+WVqnPg8rBzAbXLtkIYXjrC0H
/pGYlQLjC5Ipvccbf3rsSVBglD87SQ6Z5x4dIzS8i0dA+xJSG4iSWQENPQZqp9uX
Bzf40Kpu7YtbRvK4d11gpp0/ue6bSvBPp5fiBWJ4Ooa8iH7somk1inK0bhSw2nOL
luufII0mcA0d0vtehqPY9QuqccBbrXoFfnijBeo5p6zdBC+vLrZRDLGavFmJJJma
RN1hmdjc9bAd2uKGRxPQjIh4K2SU3FcHdBAROnN5c+7Iby5AXABYI5t4khYZ82sJ
LSYILacrOYt+wd5No5wRry5rpMxF17VUAqjd7Zd4QMGEFPj2olLYVO3iLCQ9IDrB
MNsxTC5VshSzxTB0BgmagiVC8vIRvBIk/ZH+keM7Z36SP4Hu9t2FJZgnW2yCwlX1
koh3LMM9xUyKeb0QNLKKueLZwuIMUIo2DONeh+FLqV8v4t5m/YQDA3Md18RBw283
vGYmoiOqHS0fzITQcDQk7H1UTgnHmkm4g77+jKyOcmyBsMIbphU1rpJndU3bnG8p
81oQzFmHVEAe49jEjIQqPbdVsWMge+3hTtJsgMbDdlERuQy6RkHa8vDQVCesH3ng
XIjefX12LHLITN/2wFVM6OFP0KpQTRqi0fzMV+dd6IJ/ODHdSbnTZ2zHNxHy9qO+
cmo3DCRWUN5HEclRBTOrU+5L9RWqahmS07Xx/Zr8QYAD5yng+IbfkSHr38h09PCG
nKORli2CWdsbuHRYBJPkZTEGgqLa8LYAA6XQG+jK3YX4h8BFFqV/4C0NqpdkeaS+
OwMxt2f2Xs78l7Xl2XxyzWWCal9EVRHn871byQJubZkEHQt1Z+yBiz5GZfaOczx6
a+Sr5T5GDEKVWC3uo+Vi4nL161KcLSi3Q+kEjNfOPFWC+AZVKLRuG9xmSDGA3s9Q
TdrACo/YMn3eiRoSzUcLyBZqnTqyk8ruM0J/s6bJLTDao4qLnkaGHB6i4FhM0364
/jtfPfCtG3Zx5U5eM4ikXGaaLEz8H7SDPfudtzPAmI8TFHyJvtuq4kyaGcx/sidf
JX4Q6xx2HWMa6o2GAx2RCd+s/58jOuJgFUVS9QJguSj8v7ggIWRwkcx5dPCx3zxZ
QkwDOyhbJtpKltjFm5/27NR27QEG+0ATzeUlXOSimemzz6UdOb2sdVFIPfvPstoH
VTqUsIApTnlOLpGjq2x7cSdp2xA0yTrGEW6YIUGimRUSVeuOyizmgJEuKUi8yp1n
ZRdV1NA/EFtkNET+3ANu3tCKSFcEFUmh9D4cbmvbK3ErLTD+vpXTrVQX4VKwTQmg
LCRXi8om7hItgzD9qAISa6TD82zQ4mERLjcZHRJchWuPE7XdxOZsa7vk5fF9GoiI
SS4DPz5einlJUPLm4cf0oSXsGwj0vCX5l0bUgHW/QdE5eANy70cCfP6tpok99rAx
bWTY1WgqOJOYWAZ81/heAIqApaciYnVLIcKiUln+crEyvVS+mrSoAZQtjPv6D0lE
87DlSx93XYAQ1mwu49BqPypgW3GT2GD8UmSGL74bt70z9lv5xOLRGA1jAUO7wBox
I3HiIqkgKN8F3IcDgbwAGgIURFBX0AzyABL1qjEA/Nz3nLLyeHsryQmAIf/R0b02
vUPXMYenw8g3nftdeU+gWrjdrgwVL+V+fBBFQjoLNIE+QPTwP+sFEwwRLEjr3EMn
jdK7ncXD3Y87nQdMyslTJdrmW88lH6xH4XRaihIaY1cmLvAu6n1MpggMywiibXvg
bWh+m+7mU7jC31WZ39QKwx5zztGYlxkGXSjx0TW7uqOmjU9CaKQ1MZp1nCPtn6qU
xd6XIpHvR2c64cs5M3Ld2CnsJnP3eoVzeWq3CzSrci8Y6cdPl6G+k0EniurTw/Og
8OWrS1iZ3x69DusLUtdPLJXm0SmMcvC7kghLzNfn6z3SrQjHPlM/SJJh89tqYS6Q
Z5N+A/H+jo1Uu3YacfoRQpIZM2sVbGe8EFNHbSgp9lKqfENS/VdJ89YazyjZ4x5R
Y8WYfNRKzTFb9o4rhPEsBiQEEmBJP8EJ9wPVWqrAIbqAbhwj0offuTpeLP1Wz3lC
A7jt+CWcEWcvu+SxkuQfxwBehLWsU3NW17IQG//K3syWffmy+m+/laFfR4lBGuvR
pShG9gdJ3HZTrLdknpVRu6Bk+JISXGoJS7sC2/zpAmDFoWeZXhE1GGuBEJ6cR1nX
L9k24hMvN/Pc1W1s7z8h5bFnh4PfF7zmL7YrBf54dyPeX8nNzASlPliByjGtpanU
48d2irG2jd7tm0ueXninFGbgfheTB/LEc3VAotXqCXDB1SpHDKttEW6C15KSxIDq
9lpYIdmON6fGoqQ/8pkKrUUnydaKP0aIZRFrb7qRIGuA9K0PuaKuaExDx2zt7g0U
YCl/oJnAYJWO6l+U+cah8XVlLak0UoptL6/Klmi6z7qG5Z6V7Pp0yrFiH2xk2hP/
+ar4a901oKaVB3QwSu8KwCRW+fhfrFu0C9h75KZM8gUGLn3aDKdA0aeoasubgKvu
FULkMScLzbNaz0w4wL4+DFNZ0AdAn8a8Bh2Z5ojJea66pyxdrBSVjW9AYdrUhGgC
dfdy55H9hAMbKam/p9iZ4pX6N1aj9EW2KkluH7xwNDsCizAzLsdzvwkaGcJIySsW
WCrSCOQB6YTrm7UPamoXKH/JFQQ8zVrlLzym61k5el6eYqdsaOEpVQ12Fd32z6S8
v0WqwLALWJDlCYHR6nJ0VBIIA9hbsGgAuXkstCzY8y2cDYhFlovquwdGegDsMcw6
5C5nACTI9d8pf/JRejWVw0WO4rkTSSC1sgefBDmxqmQUovB1LQrwxlpLDi378U8u
Fp1pUdFE+xwUHaQtZ7dG0lMkGtU/D/N4mpCdTHXt+edcyXIlo9T8gsxVJ4h6dHST
wiLmhIuTc6X5TgbddNapWc34D0ynNUP9s/0uBhyY5rgEbJy4yEhFqY5ROSnLtnXy
VzSya2QeCgKmfa02lTxRfyejBUMQPCdsFgsbg/9c82C4D/D/7HRfs7lgi6qAsBuj
+Zo+VicwiqDGaofvtZPbGUa+jqQ3Ua0+BRb7sSlHTEVnev2fMOnchExK+/KZy8FK
FLDnRcwNkWJ3V2JlrAyrsDxwcMxMbwU8vIFByXo1CmcsfbgWXe0Bzj/kZMDUhLuP
Be6gX2jqqFc1QipFm89KueqlLMyDXMT2sMS75SfmdF0qCUfqu+fTGjkmt1dnL9jf
kHi44NiRWWiKGm42agKrJDjbUa0drw46Qj0S3MtGmymTcAs1ZM2mMct325d1Q6H/
IcqN1+lKCeM4w1Yk9d2mGpFzWwSFjsznxZB4jgRuTYYBSGTqbG4UAAIc5kmV7mAc
zb7UNL8k9NyVULluZTgzt663rY3ty7qPOiXdyHzQw87njOJhZh5YjT1B8jO8iL3c
XyBI9E6MCkJ4Ria6edrvQXxwwhBjjKFLWs/VtQfjJMJBDWsHKiNYSjk8DOb/pgy2
YAEwQXo63RvFodtC+n1EEjkH5YKJS9YxQM5SskN5iq71uC4DaB/f1PKoeqAnW5aU
P4C/kf90KiMFumZh+x/0mEH370V8wJR/F3qu9PhPB8X4AhdT+/6k9za8eer2F0W3
KvT9Th0jGa0PzcHjUc8fl48cTafOMCmWc9jcCjrrdgqHWhJGtr6x84AYunxpyB14
JAlnf2zxG327GXPvCLp4NpeGQX+3Uj77VbFzsY0suOijswB6BaeJa2eTXjKV1vxv
Lvao/xZV60losaKN8w8z+zz0AfHPozQ3eu5XvkVvEn5nKH6Lrx8hs77ZKoy2XEbp
oVc7yqyUWHfUfMj/ZuVoShAkHheOWpjpIEZTqilhGio2MBV1GNcwspqH2ru+NrO8
Leh3xm+I/6lUQYLyRo/jbMRxQOeMyx/igNXvuANkFKn6l9z/ozY82R3MZ5wmOS+p
4uxuRmlUnGxN9D0yGHH7/JTymn9m3xZ7Hm/bAxav3iiSEihgIfNzwV4OAXtlF97d
y57IB6sPHW7rEfQuX8KUVJlcDohbVW8X1IpTZvyJn0LyULzbNGnttYw1axV/62eD
6lHarGCr/0egyhETN3WpmxUAnRWijTa08a3i8Yv22Xxdw/ILujbqgTiH9XhOYItg
TfwK/+QxRbhglMJ9epwgZaHHKxuek3NjtRpgGg+g2UAX4sW+bGOzh1+KQ3NtnRQw
cXVgFAHzsCS7H+OGg52AnbAYCGNgDxlqWdUBZIoodQMSIx8neTHmYmtESblwFoj6
JDzDZu9C6L7JGM1jU9IZ0r7iwvQmr5xDVpnJ0AA7X47oUbBZ9kNDY39ONLYSULhe
XSGpZ8PHZ4aeWMzC4U1xQJ8shQTiT4ov5p87nwe/09pRLaGnUvYShYF6/YdcdZ3K
vjc6OERJ2Cf152onxQPXE81PE42VBwdPGer5XO1yksh3QUdWHCvYToWpFhooyg5d
t2/JLWA6x8V/kiiLI8fxLQhrpSrf/mI0V+AJHmtT2bQRQ1F/uImq9qp7VSLNtepI
S466YPrZAyAohrHbrGAz9ujNHqfSfaV2k6PGAzijw65VjCX6OMarH6kVdb4AYpp9
pNA6ovWBVBa82FEC2aWrr77sq229l/1Y+wo5ie+s2WzNHewC97bd8fQv86MRVYmk
6UH2igriD1kqS+lbqsk6bY5/C13TVeAeMnUHPkubscSDtzpdsoULMTwNLY3t2/+B
2yk8ps5S5M0BAONzjPT+VoW2/i3K27OdDwrGwtRObjaykLH7mkN76airpj0QAhrp
fKQj6yKPLhTrAzSG1169dUAfhiD+YuBRXjdOw4DWCxyeiJq6t5Jghd+VdpjE3bsU
hm+8DIbEu8Pa9RE6gTb2Bto1o6cFHb35ApYUm3j6ujd/095zRryPXGXCz73lrwTi
DIVf/yCbcKjcvqCwFzwNY1jcdGT79auNYvWYURiUFiAW1APdT40Sdm8Xu+/PVOXF
G6XaxlWz4ejuNx93F+BYQmgYt/SXnPrH5YLEBBQWHEstFrHcR6kz0eqCitDYwLoV
F2PxzV5Mvio1NyMM7RAh7lhTapNizGbtGEDpamHNt2+hMpd3FaezTnINZQsCvmQw
eCFqYTNpMxmjqlWm40UaFv9rli1B5Vog5cWWxWxnEWhnTf9knbWcCNbqOYCeoiCx
sVhrLa6g5kamaW69p68bX8LHE6063Fn/RFxLdSbKKbdNBQo083zTLd8DJkX5ESTJ
CkXavxr8k0fL4Xkktn9uW59FY1TzlIPH/L2RcjseaImM9UD4n3AfNImjjxDG7gTd
/X6rzpvLlk1Jjh5LKD1KXNyw/6wqZUByjbswzWGna0ITInHAj6NEc9GLtV9LzcVA
uQFfFdpMpnN+JPcrSTDx1EVJ4kPTEUtGV3QgQ2cTliXRl8nQwL91sY3xj3HpGIjS
QVolSLFbimYDLteDrkZv0wH6Kr+LlZRgZOGt4h+fo4fEKcQpGCM1OYSYjeYjmubt
ICwsWxHYNIlGYJ0Il8PMKhgrUNcQ7yyQiDHil9mrxTSwrViZ6fq/haxvvwC3ulCA
P2MoR7feZsMWcoFB+geWPEW42Ns2Efb/iMA+l0+ViMkhGV17tsjgdzH2Xx+UYU7Y
UAgAeHwuF8qD4uada2sK65mmireRsWG89ItcgZEZ0dCOJuyZP/VUxTjXNyUptCHk
XQlVCLXa8mrB4quGGFIs0YlvMKKkwylpJJWnf9c5QdMBsDNqegxsaB54nbhsgo9+
ApKtFGS+jaMnOel85XQRpX7VQL008kOLQnO9AKzjJNrJQxdbJPa2Sy7QkGdECZNj
Kh0djmF6xp/a6Hb4p47sVj1gRpdZ4V11ecs/y/KS+lE0C1vx+xSBKm6PZ/X92cMF
Iv0LwL7VIgnuPmCyYMr3wA6i/W0HwLqzYMQ4qdzP+omSJV9Y3ZIxiqvhSgF+go2C
dwsJdpt1x56rDhE3+ji/O/bUHYyi1Kl+Vb0TFWvS8rKGJnPBpR1yoJaR4H0mkXyR
Hyy0gQForsd79wGvmq+En/oh2usDCt593ENsDiRf6X6gs/3aXAgEWzn+VOBlBHId
11UU+C+ssuF5T6FNwwXpGnzfpZh7ysDKUAhL9hrdzv/ZaNa5PPPDgGl/7wFuvn/s
O53KVCAsLr/JrImy6rBebYarRgwSJbp3gCCOm73d000SeOCsOkJHWTsy6p0YVPYy
2fOe//Dyr/ion8HvUCkyz9FAxTVFxPGIKY6cyynEz2fZs7SnJxpfHESOWOIo/SxK
p52iEQKrW9MJ2dClXsIghPEBj5dx+AljzogXdVTvs9fY8/o5qc/nqOUcIpDs1cJi
ZnrlMxdhlv5MGA1d//E4oRtN9WJOIK5mH5aZo4hfKaBQ92WFd+IvoWzOthYSdQk6
V9NlH0Y8+N+C3cGTuj3XLOfMJ5VE2agwMQBolC1RU0Yw8cMGCJiD4dLiHASBlfb7
tIXZ+mjJIZTuERlzpK7G2j5xAwkkv87wk0HolZgr+MSChD/E+fAsPXKzyqDvzmlw
DrTmRzZU39kLJgmmtVjkjnwiP9B2Bm45UuEVSFePwiaBa/0IUKsYMTbzsmJI/oyT
nYn1J6jHNEkBpxLwB0PlKokd9JSOPMp+u+CdnpyABEAUVmUZWJ7CZ/Oq0Mwk+leQ
ZqZAFNzRw9ELtkcvQ/+NFptCrbSB1rYlgvL0NKUOs3M19eGtPZ9eOtP3MwNR/4GJ
NkbcUsdu5ahWOQb6ynJy24qW92NWb87Juh3MXAiuoGa3Wtk4WdjXrDStqAEb4isO
K/qaNpBXF/kNKZbmkTx+6rKHE0TXediS4fXaEwu11QLlOVQ8JdNzQubW1USwowrw
95GrfH0qU6vfvEOEBSjA3Ps+AlAdSWrL3NG6Tyylxgofas57BKpBYQPFnPd8Kcu5
K0ACb7qokM/2u9uFizzzILNZ80vAinvPyfgzVd80KiTstFoFEU7pPVuUAX6H89N1
JfYU0Me7OafQvaHVQPdWCit5LTGZdiPSJLkQ4pKwUYEJawYDsAStEwJvTr63csKK
RkrVYn9Ek+3A1xcBdlzFahdsWXDGyaKmvmlTjHEraTABjqC04+QDaYy917R7KBFc
lXNylK1Y2mIKvNmWy9hsQXY48cCtotUU5URsS61r7+w3Fx+RuGaQUuI+02V7NHxj
FQzXyWlOuSXPrUHwZjNf+QkEQYG7qfoO+JtX/uZCJ5hBZtQTrX3oQ9emVWPgCHXw
u+dK47qerPChbuS+vghdDNviOx44qtwZcqvSgS3q/7AZ1BMG+jYBdD4IAcJUAYRw
E3cngLYN/QzjqUdnw9lI6QHjPY+j/7cbaWcw85hpVQIGEKBanGOE7sSGltkgVd5y
MSk2M4fFg0F1dJg5aaDO432RR710h6lmni+FMwU04jFtoJAQgbJy+p80gGIk7Lb2
srVwRCmOPvbmYgNua+y/BU5GDSiOeGoSoFPsz0XdCgKrCUn6KrcYRwNuI9sZHdhV
jj9uOhBQfb9cw90C2bfUJHDPHdVyTmvs3TF1JXMCJKWqWygOekGgg/XVPt6jIRsk
5fuoZBdbUHrSsugHUGQQ3mY7M0qnL40mzn9hnlCRureMb+HcCQ16xeFlJl2rian9
KTtT/kEnf/wKcUhDgpB9V+BgMLkpWPQZepAdcmjDuhmZgnb5bozmxFL88KgqFe8j
wNIBoqGTXmygTn45xeysBkcZHywZnsvN/eUNt8cRI3j1Sny7JDX+GfzI+Jz4gC/B
528K9kfEg58C6/QU6KeOKLYoED7D/bRAWPwzDMN+nM4T+OWdOPOmlWLm4ycT4j2u
NaA1OiktgiiU0+c+vou9g+BhqQP3YmJ3XDbRFB+mMVqakkUNB79fQslWXRjl2Ee9
KDKPMsBeUGFtz0TmvBtxeli+JkSY0BcMM5qsebdaSgx5mHEkRmQx1CC/PvjM1XDR
nZayzt496+68893h68hezcU4GItU9eBRo/WgPW/Z0ItOl/KN45LdSh3o4fxVrbEK
fCQdWC7G/0pJSIOKUaBErVmC3aUIFxRiJB/Bq1KsE5r0S/DKBHc0+QdbvA3CAFgZ
ijn/MvqghIAmm2jb2qDNmve/MFChFTOVtAOyiP29WvnbsH45pSXSiK0PIC+2FWnH
JeBulCUo7MQogCBHGIAdinNezSnBUmnofS/ktenuqmw4fafciPrQJ/o9W9vOS0c8
+3+F7bplicE/HjEL7EqZEmYQzkQ1Z8mAYse3agjou2RlfCDuK2maCEYTfbgZPoOo
nGGeOqIahoGpK+V1OYi/hF5Vona9PjRWd9C+BogaVaNumwPBjHh3/vqKc2z25kyY
NXIm+3Um9NXam7B352SORnQh/FZu/j+otbuz3d+iqHd+HJxuhAOjtEOVLpLX6C8R
gUNaFrMPFvE8T0ldmWC9P1Q4sGGCfrPmM4ugMJ1n7RsvL4zusFFajoiyx1HcBXBr
P7ozjXhC+hz+Rl+iyCjphKnEMa2aDU2GUtfOXQY4dDDsl5pscZ3xJoK7xbdKAyO+
I1PvW1xnd7CXQ9hHUY43K+FKfCFYgJRhMmZ5CBpE0wVkGxo6mlrBlbB1jHvBb889
9n3KKdo4MjlU7USaZhj31WP0J1QZM/GImMifkVZmJB0UY9YHlvIbM8w51BhGckzk
ztGNr2RITdlwLVKkI4MhW/V+ei7OCn3CXewD6JhShsYhEzNeLasUxf7J85aUvJ/M
2RNBh1YEpj9fFsmnBRwCaDiqkeAoKsUnMUSgQvfpzpu7PdBamm86BJDZKnZwlK4A
C1KlrfcSQl+v4mCJGqR3790OSjpk98ge6DhzJeDAfu4sP+Hm2OzaRIOGNR0zY59T
/MoFRFdVRBCyoyl9PsPZGhtatA9+tmrwNRLhP/G21N09pTebkF86BHA3WcVeCSU/
l9lhr5YsEaoX4tEcL+ffvqSefINN/UB3J/BLwc+wRad1zpv/Wam7y8Vuh6qLVLH1
UkMs1MWbcl5a8N3/PThFrXDIZoiSsSNd6fjrxP5cqarzjw3wmN7cZv2xYNtyiG8t
BtojVi9V85+cT4mi3ucBPmezlECCHNPZHBewxPUOGvBgn5J13fYcsWbqMhM0ZA3X
b+NM5nCGqd7DnhwtJaaxoSdUfcv62VDSvhX+TR0nVQQc6FJuCqhcvOT/juv46I40
dtDUZ9Bm7/G301ynFOKkBt4P+M2zcIRHGwuYyBp9IJd+BfD7HVjCKQONUUsv1sbx
Vxuct0s1WcvxO8vO7JQm6gyRsTkkdpQ4klhlZyWtx64YxXN8c7wOCNjNmyzL5cBA
Jfy0aUe23OM3wd36N8znYdsyvyOWO/OrBzzPf0j9D678VnvGgxBB2bx7aquuenVv
toEPxpDWXg+bRY4KkRpUBP+xcRDEc6JP3T1i1Pb3B71MxCPMEa1BwasBtBHv5462
EPF+ZTlTEPNYL8u47DgHqjhsgPKUdDBKB0HFnCtGKe82pxpDxileVmVoFNjoOR50
GYiazAWoh1QvOWT+9ZCsL9g/fbi2EjwTUYhSvP+j8uJadsKKhVJ5oXysbJREPzZM
f5Kf+nl4fsp3traUqGZtk0055ep9ot1pkIVpDp5uTJ8UgRWpliqibx+Cc69QnRmF
Ks9N4LHDYXkzMQN80fi6Q0N+jw7EQ1EJEJmHI6yu2KIzxkU5wPP3HgQ3DrLMkR3i
VxBfAMQ6hwDHBFOax3u0o8rMYaRv6z0lmwo7tITO8BaRaT40iTlifDSvqQI+z9lx
ts7svmA4/IOf9tuZARpzmUSlvHwMBTxHGdky8gkOTL7rmEaokqBeAASTKntYsDhz
1QqyF/nI9Z9qUiRrnwt2HonarOGW4fz2bqrkMI80t/itwjU0h1UfXMPZVlxOuEqf
OyWzpKLY7v3okB5VcQZnAOLO6u+ydiD2u7eX+yVHBCCTgEOv9DnVOBihgi5xXNGy
l7Ghn4+tuqKcVhqAzGozUfkGqI28gxXCwHPpULnjrbDt0ZSU+dYXSXjAekGCk9vn
BrM0860Hu0uDG2S4BIDv+a11sr1hNmklGNRCn0tqAUUdtEGuHKwCQnVeDZDJM6iq
Ksx37q7iXY4R0TgbzYrnwS8utLgbrlsfHZCaP3FWbm+JLiwf0W9xrIhpQGcTfELF
Z7RBVuVSVTV83v08binnu8/GRkrQbkcXe4DewpYv3fX4dM/BW2IvBHzo+yS2uoyo
43pXIIkNpeJMM2fII9r4+Pwn91/MzGdcMDmTGi6IQn1PYW1Dh2LkWZD7NC1sylq1
1fSUmyCKRw5qH/WrZTUY3KR6zL7xcNnGR0/pzYH1khNHo37/5A1VE6SbNFW3kHe9
OWuSVqJCIB/3pewedUz1uges2P5Fx9hXfTnHPTGxEWBsmIhZObE5Z7XtP7DvIgyE
wSBxp3fA5dp7YZRKVU5Y2uYKdX4yi98WWQ/D/bKT31p0Yn+1R7coTb+B+Qm+3TPM
xuuhAEzOFixUEnk72MqFVzWKDlcq1ip02YeJuT4me/eDRW8TQMdb1brXHkb9yhOB
fYEM0nsBVlvR14gAWFwhB9MixptS9KQQ762W3T0bcy0JlHbaqg0hhYKp9jQ7l9d5
dcQMeZlLj/XpG33+yy9yhPcO8ozr9Wi/Y5qexTfNj9JfDchD7RlB1sKfhXd0sRsJ
oIGIWur0V0I4rqjOS3PuI2J2ltarPzzpNnMGUF81NGkn96L5rhjYYkfOM9N4wFmA
vLHunnq2spC8sMIYDX5FUFzfypAjm/RglkRREBeq8pQN/nxBy0DNRIUyprK0OCYd
fR5v6WuJoyWu4lOmaMpKiACSKn1O//vv52MUb+hcjcwb16LC/z/UAkrPX8fCGvGY
HBEBicwBF0QvhPtFwsJfWzFUTzyeQRmMqiXXSxDDIcqQlF1+oqttbh8oGfOKAQCp
n1hnHYM1a+5m6NrYKyQikaLpCHGhoIJAyyAMK04gaTdPnKRyf0lhXBY14XaGh/kQ
oR2PVVaj42iXKyeE9VTDuAf8qQc2ftN3pRS0I2kET+X3NR0MDRak5npXWo05GycL
HI19hNWfF2X2rQwr14x3mozFCBXxQGvT4u85RanFLBpZXyWkDkQ7tDlEZRZn3aV+
SfWFnW+S7dAsT+rKajM4mPxsepSyPCiNUfrjw3jlrQY0HTOpBUDqDz1kO8Dm1hPw
xtts6fRO/E6G+K9R09775NbZVVr3ZNGfTHp03FcW8Lh7q5qNJj1Lsfi+gDheRQMi
ydiK+PrcQPY57q/QJZxmlTPjXl7WJFTfLyZ7WcOMlgrR+RZcAIeXC7UGFlnYsEVj
3AFPYCtiXs7mSfKW8nFHC34VTVivS4h53/fNwCrfJL1zWjNehdEKWE0VbikuhvMr
zCCHJ4BYOwVgZOa2AlmW9JCyaXILK2kV1Ri5H3fwqkkke2MQ/8ZEp8unNKlvfh/b
gFXVvSexQvDnX46Fokp4OLEzd30kNVOmmRwgHWB4uzGRDbrlO0qaOtVD0pzVFeNf
RYwtW8vlC9nDR6pBt0aNzB18ZTbWQlv1lJ3vOeEzVxC/ZB01f79QWqqXcRmBqDjR
h/3WSDFnuR1IKptIrQPYuw5JzLZhGMM4bS862YZ7oOzRx7hwcyj6aM6D+dq0kErF
uliQnQuj34Wp6NICnAxxV2WcMim8Ex4cxVBS99Gzz+2I8I06fMC7AIFNKNVoZY6F
yZ/S5b6LdFGXv3eig05bXb4IJNM/p1IDjTaoK8WnTcHqQvrd3jd7nHnyVxmfJ0YH
LZEXJCpJZFnRbMnlDkz5eSEFPfqry/MHZIQA8jYiBJK3NRiybmlHYEYWhV2IfGU8
U7AdR43RoQBI70v7Eu2w+NjUwicNPetbjLlWadrkEG/bIcX/CgiNWZb95WfHZqeC
PEn9i0ecb3gbX7lI/ooaIP+npEebejaq/XU+YZtx0/oGjmP8RYrlUkgOiSgzdVis
IvmWU7KYCOmuowTDyvmVcF9tt38n3J4NanGO4CISglEfdiyWXVNof/BIaYSzL3o3
97maMClaK2ZgzYrBuhm7Uw7weY+EL4F5wRTHwW4JDSguLsASOTwGY1pArN/8R3gU
/w9PEC/99OwFlh1noCO7aIIIfRWw6h8BugTtptFu6lyY24PTfVRF/S9+SSkJlnOS
SrQQOuXLSmDyBz4e+AvbTxpl0mAPGM3L0xZ0g3ty5gezn0yqByQBV+twgjed0eai
8Cf7i+T+mxTi1+YrkCmdI2XXWxDqeLrydv2V3xDyKpfh2oLeirnVbYIRdwSvQVTO
YVDY4dpFSUz7K1Rd6753Am0jr+I4KjGDerOP65XNcZDa7lZiYQtGymnGmz/jTtjM
LryPUN67raOGIQ+PbTbvxmKH2E0jjKMKAqcE16Y/KnkBqbrEB9PYWVjybGFzryIz
+gXJPRN4OG8Bnz4XxdXZaS0GysRSQiLd3Xahm7O2ZJC6zYjlcftk6DPu8xDs0r5m
Tq2zLqlPOW7ZZoFFlGZ22xWGTpMHpAC51a5xQeXNw/NEfIvSSRtlfQM/i1sDqcWk
BRxdm802pEYGB3n7//dPsC1WEKb+t2IEjr+srJCuvJfLYA6QfaNskFMS0w7DKoUP
6EnCvS0qGZWLzYZmgn4m6uzAK0Cais8gfwM0DkBo97ErPho8wI1NHX6taqt3yoQh
aydNhSOWE/JzBAOyW0Wx8gJtheTh47A9nDPCr8MfHSF6xfOyOh9R9/InZVKktsUa
rJgNaa5hl9C2n7i82WWvKMk9UDTftHxj54Q/iiYjhWe1T/UzX7ZF0cFSlfdDgpQq
Yz/z2N6RR7yKfAn2mHKPHwTARL3ksPKtCeS3z8LAjXKHiJtPphcapCza0e8NVan2
HZBuaeIWP2vzZ85M/jw5yu++irVwzSk7tjEBNm+RXZZkkLD0Scm0UhgCEyhzLbMY
8CcZYtvOWeB+xShWgFMq2FNF6fD17Ky9pBvdTUNFwOjZLeoF1eL8QhYvhz8KQE20
vAo2fTOXh9g6RI/5rJuwkyI4QHvy7VTe8g2JrKQ9ZyWByZMQVHD9bZXKSgWMDS3k
Cgb5kL2KXMOZ6hXSxXQsTzzFWjHdbq+mF2tMzeXwBJ/FZIrQtfJOQRhJeN1e5pMr
9941JOs0MJfuzAz2OIcqRonJmA1Z2036S6VeB49AMr2SR5W9uAxE+57DdtljB/jX
L885UTFIgSfksg5MHh6vrmdMsYGZ08vhJ3nstl1xZ10+gjO45ijW8Sgh1s16c4fL
h54y1BAbnbCieHnnFoJTKLQTGPNFHTfUQMzeP7SisT9iRzj/b4+ha8SnvLrJTNV9
OjlLNUZV1UKRDEh7v/o10Cdj+kaiiGgF8KuE7/mK2yGKiWiLe4VW7IZiX7yoVjML
wrHkOZ744UOi5hez/H1PW8e4AVKbTTJ3ZlOx71sH4AdrZ3FEYudnh6gUyv7aa/8S
TrG1Yc68Td4Bb0SXINRWVHZ6GG2mvDRgP0wN/j3ZkzpmpmYg1Wmzb7lAez5qcNku
wdsuxh+AaYTmQnojN/eJYlq68Oo8JBsOohuZcCM7NAks+lCltTSU7XkGEcvgaQFl
Gh5jmtvur4gUDhgTD6nouM889efzzANEjNUwPrFb/I1e66cr/L/OFNc3DGjWFR0p
+ph2lz+vHLXNTzE+Xc1Ok5xa51EiPphNmepUphEvMszq2I3+c9fwhliZIAAmzTbq
NM6/FG+OKiQKxdkGn7TP3iHARr7xw77ySiZNMZlENw44EUihXPmrwtMYYksTVjI/
nBbQ6IHoLPTDLkyqRCQjvwpuGSc/wcQTc+1rji8zC5qSPyBYjCIehtY2OR6a85ht
5zgLm4ZAifhQgvbIuQJ+sxoI5KY2lzE/Mj2ioWSqFczJONSlU+lZiu8NAd9sxFZ1
tc8GDo5foviyOxr0I4mNv4ZngosK2QaLa6pB8t+tCzmvEcCb+esKElMn4VEN987F
CfEcF0Qkkh6vt2goBoX6C/sRWDHabimYdJa6uG4oGMSKO95iSgLove71j2LtLAoG
55dwJBhy19i4Tkg71XfExUkcouym8nTEx7Ll4RnbTpwqUcfqqcYvLei9GPQ4yP7o
bRf/vGPwuqF71pgs5Y8anWztZV3XszDbg6ExBT3v9e2ekYeqJXgzPaFO50lfvZ8k
QAwiNRmtD/BCEPnFgtEQfy7w4HXyhTLlOIcszxHboVvatNq1T1U404eHrKwBXlCK
0oOX06N3uSB7+DVW1hbK/ES94gU+we/hQh8i7GCQKfW8jAI7ZHNYGjj9+Ri+CV+l
CLdFxEVonk7pmxqucvBIXhMTlarZfrrAFcv3AR0navNfIiPedyaewAWwnas1AJpH
QWYsmRSx0bPRU7mfqzr9Zl0YYJMZi/9PIlcXY7C2ptKSJmVQKL/5IJEshKH2mcn0
AhEg1vhc6vuWMyzps+IbQBFo9Mv/lTbVgWuMiqNAbzaepFpqgU1IoqBu+LAgptq3
1u3ALOf550m7YYImYXqbjH9iycXkESxgrzqz1ycs7Y7ze8N7xGUR52r5obFdigtL
zA1VA9c87+yg015NozmdTeKBueL5nap53JpHs0zoPHmsywVzTnNtBm4j9otBNE9U
yvv9CWgby3/4tLuoLI/68uK4h33j7J0PiykwWhjFIvcikxGHW7X2qhkBZozHzLZq
hL+wZTyDhUXG7u3w44laa+O8s1PqaCUuwe+o9p+9oiiXaXxnapbifUd6BY9iJfsF
0Cutms4yWTx70mm1TGyggYI+Tm/dhjDbDFadBNK2Kh5LVnSlktdytMhkwnJtLnHv
+abuMWmpfkc48J12xw3P1dlRcj4Gomzu4ZUNN/Ogglqhog1+7MxASKsXHzhJOQgC
XHadb5Hf1yY4se7T9w5vM6XCV9pNBl/pfTU/sX7J1RlTQ1VepdJ4wAlYCDEOMxjb
STwev7z6yupx+FF0hBB9xpwUb4R2p2ap74zKNlQYSsjjq9b4JupR+hFfOEghRDJL
K9KjLJP8oozdCEA/hU8yKtTEGC7VwKT7w39uia5quPIUIMuH7ZEvfa1FiIiF0A3F
HXf3wL5l5QFDsbP8yBv5FKI6cA3ilNtOhtv7ofj7x+F4UiBq6ZnCsGif6CUBtNgG
Or65ajbqaJXjvlTTVd675Al8UB2+Z9B/cDNVgLL+kD3YAM2nnp5Mls+SbHwMxVfk
Go9EWy1ARdwne7IQ0jKrJu3aMBvz94mYlf7diGE43WmRSSZ3qPQJmNxgbWb3yWFo
DPS9XWyWv6xecDPepxJoCqpqn4S5Ca+LtFk8fPyxLmRnorXH09uioBdsGUdAwnkd
t3oOp/PWW0zSa1j0hQmveTCjsHLk85Du9bG7QTSQ81EIypddrERRtlrddE3B5a8a
FpjNzfIlqU//jHXoCifEmeYoWQUW7zRj3d57cCkcHekwqR+gESa6pue/JyDG8ODl
nZAgxaOLepDOxPDamsPLqXMIYQGjZUKPjiF9BynH/BbHaowUzXfpV+0oL1BgRSQW
qUdDCU0gYtZBsYKLxXsW//EaKPCvSLvrPBAXQIbXBX2KyiWY7HnoeC1xlBGLgA0y
uwfwREOKPvV9/EqT+Vo1na9UcalO3TQXjcBi/ctqdEVK8f2JubTY/ek+Bc+zjWfV
I/d0Wzc0zk/l8SqGQvIvsHI19hHcJI69k4enJlVv2cXVZgRR6k+Mh+MJmqb5PnXP
RRkT4/9tsUeqp2iZxZ803ZiVOMMruBC1SHwIT3J9ZlzaMmIXRquYfoYk4XBgIlWn
1dPnMzjsCCoK2veZdJ3FYxCMqd/gchluf6/Pgi194jjps78Rl2n9j9vdqFaq9WUM
F7iDjInFrdEPhAxOJYIoTM1FC5TWxndMFOUDaaJ4/r/pRxTLdeM1mjUnRwRSDv24
5poFn8N9Ifwtol6TXzZlexv1gDub5FbrycH6DlsmztXaEQTnRJ9Hcmb/2nPSSF6L
B0jlWbqXgL1qIQiddWtq9YKa4AcbsxcHYvkj4NstJzq0iUs2pagfUx4evHgftYU/
l041xz2JRVltmiv097gGxDlxlIEW3bqor/1efTMNvndwgH6AW82AJ7y7DCVHYaS4
hD3uEnR1BqlFFZPc6ZDdfBTP9xVXoiKJKOY+8Y0hgpRkm/0w1Dj3fM0cvsgQ7AZm
abf83E/XGOde97IL/q6bT7B2ha7vdHRvJOkeKizbyFIc7joNEC3bbnFTb4ZYbL7n
5m1MqVTcpprm1/evvyhv6U9p8+Wv0fsucB01jfsr86z3eWlVwbOQvfyNujfn+gd5
Y8SIier9+5RM0i3efrRpzpbSly/2lRtdyV9vIABH80Hk0+Wnpwt5/hFnzJ/AONm7
QsOdSkbjE6JE2M0Cv3FqZY0f8UJ7R23Am3Z1a55vUfl5eFsydf5PyqQN9dV2cBb9
h2jPW4bkeLv1AWT1AfbYTrmEOippcd/OmmBdbPfbRjzwVWhOwYyykXqldd6p7qNu
H6N7TJoLF8t94I0ShZ4k2uCFReL3YZAv00Vksk4VPGPsyd9w38bUMIc+4tU4JeUr
Fdd2ZyWJiG9QRfEG9o90r2tGV5m4HbSbAYVjZhAD6CRGtmSMnONw2N+PbZ+FLjQF
i3fRnHwVjbRiP0DqvMq8/2rjKpXpEoyNL7bnDqo7iZ6y9GvpQzkAvSL+efmax7rI
/7mgID1/+rH1OmM3jdf971cIRJTJ3X/jliVIbouQcwaCoxv6zkcvjNiGPUTBYMv/
Tmf07tAFvBVzE8bHcozKLTAKVurM7nPpxSfl5u5A6fWdHbZgtapKUacAlZ7vS6Xk
egkBMILBExEXV9nHIrDHztHZ0Q/velXtehEWgp84yyIwJEvJsJ/MNxtezpTH9JYu
zQKANdkTHcEgvc8nagAWqjdy1Nfwbx60AON13lZhPlMzA6+qzvivCDg26xCRTsHl
rgUvSpYnpHanAupQlUsRvWl3tyyKHImiKW4S45WZX6+zWJeoy5Er6hRtJ4edB0cn
zE3DWR3vOK2T4Lo7BQOigvJ0eI6qS+CfWZ6G2QY1Z7oZwVEKbYclNUJXG012YbL5
ZjgCVWqujlx4J/yKvrcNNbg1UA9eGrDICiEHZmbLIEXs2Sjsjn3lTVFCIHc+G7OC
BdeFuPEUGUiEuHXHSAnZwiJGDJ8TR8CFfAfRmJO3uuEdTHbajCjUcBEVGo1VpdT1
WetaFycgpcYU+coNmJBwXNmZUsimJlItJUYbtx1vCMS7OvBimXqYceY8t/a2Nyos
yVaa8CROJCL9iI6v+rKhaa5ST9mLu+lUB+Rjl46ckC5pdF2ULcunqXq2lPTX5C8M
ahS06KcMOE7ODD4eDD4rAXUI0z8OlX6yn/yF2236CoICEVR3BvsNWs6QcU6IQ/Kx
KUlpe1hgScRRU2/5x0iiy7sRj6UNT8I4JAHgwkpTIYYiYRxYE/vFV20Pfr+IKmtm
ziPnpUnaL0wNnsRw/g7jSqkhXOsRKZ5AkYbn3xO++AP+t42SqQqM5MiNzt94tFH0
WBMLuxovJbTc3k8MV1gHpP1QEOBr09zsrhIvGDmUCrwzbSiOjdzcNfQLRbKi7xpH
NfGj7aH4+kIufPm7/zE2adrhx1IgUxHfhElnGkd0dX/t+awTiAz718DvSbAEAPi0
Ba0UDJtrroQS3ZGVJXXH8jCGIxl/qmlbzKnt30iTMpBBiDN6eOvRmHtEuf+VDwJI
wofOiISVPQUZmwwXH4lXzOZuuLVQtCpzQj6JYhIrsLqf5J3HeMSr78k7XafnDqsz
DWevwn2UepcXM7Uq4eYGqgw7lbgHYA1BHj5xZ0SzWuoIoE/Oxm+vmYPJ6je3RJKT
BTvSDwlHbYI6nhgt9TuBPI263/rIKHYlnhK5v7UJmOfH59sQl+nTo6dRbM0ogNZK
664ukoVojGjtyglOFLR9hiTm3Fewy8GhyR2PReUSoXTr8c8TKXDXN3hwOuT8jqHq
FBCbVTy6kYNCai4Fp+Jr2SUViNJyvs2fQorYdoZXNiNa3HHNlTc0V2Bd1Mc8rBAE
vm6HlncWNnfa7kcWWPUF2NE6dDnXXIqWR1F8h5ftLsYYt1bzrYbiHPNkbXq0KFLV
W6pTl+tAQ4VDVS+1x3iNjMoa3isDOpnqLGZYSJR6iKC4P2ec70B90w4n2o/6Y8hn
dNqllVcQnPOthLafwnUUlkbXPX8W8Jwq48ps4YsSaUk9/8k8oGDUshvaq7UxlyNp
OD09xUc8dP5vaWRnr6qMMUV5pHup4oGWw0GYuqs4FwVWo+GfuHo5tdBZkmswlWVC
b4U46JRxLDNNfxL0wj9mufWyIuknpQ3191Ef1RYgt1M4Kbrag0uf3//ne0dAPPhp
A91SXA7KIHwOzkw7HW5nroShcYrqKXPYyi3OdXuvGj6+V96eBe3WuVuOZqWSmD9S
cN2Yx59bp8PgfrOfgu8ClfYpvEII5GWsLw6mz21hd7x4e8twnwkndmXPPJ/qIZf/
eJfv9JE62GV3ObzJlVDePVeT7N9LGQiBcrV5tRFkc/eCb3EIci563hAnfY4smjqc
zw7G3uLdDfw4ts1s9wKADIFGvfT7BGjGsJd0O/ZS4GnFl52qBIPsLMElyE5JtKkq
mKQOwltWd+8UiyYdqh7f9WCbksGpCvyW8Yyv+VOzincxs9oER53+Rv2G6bomrCct
nvlkVkqfCYbRSooBy67pfn2qGJ+eAcYGnYXDKhh1+t+PYkQa9QDkBZyIBmcp6uAG
YnW72Q+hf7sVBAvuKS2WuXzMjcFiZkWiBpnQy5hR3pfJUJ6K3jpsV9/uJdk31mXI
p5lGcsX0RkyBVAXF87sJ9g+GfglV4zY/p2V8us3rHP9RQtM0AOqR1K19BQMS1Yvp
qIyQePc6KlkievxdgMrGdHCvTfyyd/+RPDs4qSuTlj9HrIbJ/IFoOwbUyVclq53c
jTpOzL0qtbbnlwhiGI1HabNNAcw/PwWoCLMDQ85hxwPY5Kt68jSqRm5tetN8gBNg
/RTa8LRwzxqeoGtJE00jylUTnyGz7WpFKYTomJ0UqYfSdSFegppvnVO0LXiOxvDG
J8QrveXEfPFxHKygkA49kCZDQUYCiOisKYXP2PklSYq4y2Oz1MtD4G9mTaTlJpmj
ZJfIUFZvyvbCZbJb0s01Ri0ab7GT8uF1a23mUmWSRbM3RtnlilRERajQHM4iHD76
dJAs/oje0E60JlMFgv2d8syBAWEiGYk8aa/HOH+kqjy9skoZuJwXxqL7xUy9NqTk
sqz9cAyGvz+n/QAGkFzRaJ8bqBMYAodTEMRye4hFPh3bzL+BYtAuUKTU1Aan/TpH
pjR2yY8570Z7K1RuAgu/oognzaRTmi49/o7x1AGkHD2tnzKq3PIAwmUJuqV2hT3X
0XY9etgM6Xb/yMklruJq8od5CAP2INNm2cTgzilC6zJ+G5l2WU9amNAemdz570e+
chGkIKd4oQohI4uzFNa1JX0+B/veSpyCGRgFfDVXrU9UNQD4ThlX++RUA+5BPAVz
OacIh0XgttRJKLX3eg+MvSjPtU9LLWRA8WmRHHs16TLGFEMAXBnn33PslxExmkO6
mlMitLYsL76ECYLHKfRsPqcr9pC5hI05Q6At1tEkidFZumoYYze68bm0CbFIhirA
TRD9lYINbO74vqDe9YmBjudRomXg+S+edGrehai2XxSYAa42hT3gcX5xuuO4HqgS
7+f/YadAsfsLBH9ILDSr2uU4ToTc7uK/zgGP6SiREoZxqeNkhybLaSWTKWo63Vs5
Lez+0AaSkT4mjfCbe13M5F50PxBP79lB3y6X2vHllbmDrzOTzQpO/ag76L6VBDL+
Q9lljOrCawec7BXcHCRyJ92CAy5K3I00zT7y9ri/4gYav5TRAGbRup8jvuoFeUST
xR+uklzzTL93KAWart3ocHenCzMqvkjQocEt9AyhQFc6is2TKvnFJMy6RZoTL7yk
+GoG/dKChRZwn7VIMC/zK6Zuv8f9ugNAXujn9kAMHjoTqnEb7cehfoaLW9TAopi2
Vk1bmHFtnaiVqnnTqDXvqWwz2opdNBkiRGc8j7f/MHKezT1/NoTeIoVPeBBdb8WD
5tRYquQRjRMMKPJ8vhwIeGGZcow4XyXVMGL5SMditBxPQGs6fEiOgDG1+37mD4FR
PGsLeuZPJ2dob4tP9mIfO6omayLcg2iuBeg34mTWuRB9B05X64Eh32I5FbeZ4U6/
C9yXNnAYQrJd03sLFuxrmB7P0xiif1zJVEbIvnpOA2X0TVawTeHe8wPqLKDzdkh4
ukaMUgHkRzXXHYkKKHsYY+JiPujX/lRU454g+oKQfbzMzhuRfdTwD6gBCraLLQWc
9vGWPCSi1vG50rZRQjamOdjO/eFhFqERTwiNHNBH9Xo22NX3Qtc0iYP5IikTUuP3
mT/ZfAX3ZrBbp4tbxiATgKJ8SUu59ZohO120HKqlLHEGXSeOaw0dmYHX6p/m3Gkv
+ChZd+zVUYA1c2va1OKZX80a+lktfTMRAszu76uwrm9PlC++MSp01tCnYyh5LjDS
mnFntK3Pa+LXtE4rfhNEd+0mz6bO8rY7V5qP/mKe4h3hgCyAdJEFf7dz1BmTbsPk
TzkrDJPzL1CJ6S9cqx3nURXpkieLBm9OVOIlOE5U+OqDeVkHOt5fWbB7IKVwHzvF
sjVX3PoY6JguOApkI3ru73wIiWXJUlohVqZhHEQ7Cmj5djE377sa090/UuhT6wUS
yPmie1wZZRBAXldNhRMM8PH7Kvv+vf+2mzG5RHBpk2+3a7G1hapK1ale/vJozCra
a+8KoGdP93ZUsF8n4Tf6z0SjCTf+VwYsnxKMPLV6TwP9GA4uJ9nclzc3YrDpl0Wh
6a0DP1CF/g6+IpjJT1YfbHSWnyAtxLpq/ASTw4to6agLvxXOS5uPF30P5OS6pgaS
Dh240qkxfoVxevU+WXv9KW20CR2hz26lPPZ1eLZgEQGk8aXiNV21EiUjRNOULtlC
i9oIJekdWNXQL9nKmG5s4krmVSGW/Y0n3g0Ufbo98U1Zljjf6wpOKSTFu4uAvTPA
D8Qr03CZ8h0q4Ly2KtegiWltZAqG/O03ggUecX6677vHepPHghs8KBsrl/TgFxpF
gGXaNGwOUz/I0GJkwkyUPtBgU080DQtpFdC453YuSg8LxHIOby5XSC5AS1h10fNU
6XS6DXuVOMRr/jTknRcHk+j2acgqGaFwgvAey3FyjQsb6HN9o/JdOhHRKtxoS0K/
XVg1HNDa0QyUYFpq/fTe1vsGa1at0kmpEFt8ATgC+6U2dkoGm6PvNfkENpt60DAo
9Pr9edTGo0p5OU1iLEaXZPVl6fAtyyhPIWgNO7yRdQq7QsuqrwAdF+juh5hdE+QR
9dDPDS2dwKV4HDjLx+eh3kVaei9SB10Slhg+8HUPHzIdJqk4ZwGEOuVPdDuoZq6H
Yn9iS+cXRf6uLuqKd98RzCnAqlG6toWQPSPS8IMnvRgj1hT61rSY/ueP3MkUR7rh
w7OA+p8ao9L9s0LKyakTE55yY246jh4Ym0giTzRgast7oeTnwsw9OuPlgRQ4XgvE
KI9qYHlPLUewYFuiqd19vMCUR8aIF6aqvL9C6flWJhcyrT/6ascJKQm+Af44Yetu
Iednd1qT15qm5d2KZap3X1Pd2zEhql0LF+vUiyPmYVceMqZ7948zGcaHPr40A3E2
HR0yU/2kh5arH6s4uBTglD4BmvHVFYLa7s2i+zQ7DmiS1TwiaZZU/2a0xIW56wxk
hZN75Zf5vC/MCuEJOX0xLeGlOPJpMxx1j6T8rwsuBGB/ugoD9ybXXLgdh+D/wdLv
7gUImC+N9AUMKtHR2q3iZP1ySQtOrc+SWVWDgNsYM6yFrsK3SyU+9OZgvwmU/dXE
gEuaprujbm5WTheqwzH+UL5nSm018inkn+UJmtzQTIrVPga/F4KgiZj+BZlDLSKq
NdpY+XvJIoClhTgsL3/WvwdECrNbRJLkBikTPeHssg9ipzjsp592F5Ovsu0G2A6N
/SQLRjwBSpNXE+mU+IgXHSvoeQ61xHta4UOGHK3C5qdCTLSqlqe2ObQO7M712Kng
MMS01yEt3IgVTELSM/BP0SuLxj1dPOSiEr+qcg3kNwftEpfab2DtTKyZIgYXGuQU
qZwS4p+pMzCR1e11pHei2d5pF0slNWRur3q8rMlLhbNCC50NkvUyf4GW5HasPlJX
Pt8lwBEmThblYu4KX8ptjejJadikhyFgzKmnKSGIe7H/hDt7ZDsSyL0Uww+QYqsA
3qNG8aNEbPcoeaF2tJ6I9AW/NvqWZZx+YDTbYnHKlArv2rjE3UEkKaZva0RpEdw6
SstBU1/5PzLSmvlOA168qd3WN1IAT1vjKuWiOENPWcJ+TlfbTiAyAWomuebxH1It
rtB3LaQNyHwOSapv1rAc8sQjHL4tSVTnshz3Xtr797ZyRwyVbrPVKn2u4wVsHaJo
JttgCWrWAtE/PFtCMGrhDiH4zkn7R38XVkq3saZhqU9SuXGMqLDDrsdftFTd5ywL
ctXeHb6s13UU+QJOU+KktMTF4ncA6QxUbLpnKK/U2qQmXsM5teQ1t0yI5Qhbt8Me
TWetsRt7yFDPkKZZXZthqBR+Ize5IRcilCnBiEaySpac7hYm5SgfDcHkDsP+oRxX
kbkhIv3SekE1+oX2t1lTQcYTX9/OG2NnQBePPVIx815EgOmlfvyqCyNQ2s8yYtF4
ihYaqKm7vyag/V2nvSgGzHQlkRfWisR5vDGWsA29jHG5SVOv+CSAAar3ToVIiDiO
YuIj7QPBP82zyzHeABjKsRdS4kVzuPWCPcqSVXMwheBq3AHKtgQcH4J1x6KqwJvA
qdQeovgDeQRSuL+FaTXAY4BRWJSwUNdn1og4pasESlBG+n2q+11CIIyjJRlYNpKg
xHt0N/O8JcEQTBgfaDGpCVPDC4Zz677ZLNJkjy3f+N6/CY/s17pKbWWdIna+r0FR
PSpSf3id/xUGz77itfEN0CC8jN7iEqKGdPLKtL4WOOCQRqap6VC/23RXzp1MR3hK
rzqqAMqtCMsHWNghfycW15UZgNTUjHINpwZp27CKBWv3ahu3SCmAbJDAf9WybTUk
jgf/3c8RRCEeDKZB6aUn47gXfT+C5NZiUSQgCPqAL90RTeHk5Q+IAtQyHrOHOoQX
8CRtsVCqoS7EEqM5kuOJSHJqeXGlflmri8GWy81mYOxnf+A0dhARe0A8Scwab5fA
sJKVdE79z3/Sz2/UZYVPvJWSqX5mIcRMUej0nlf8iyQtC44e40dPmylR1Cq6jRSf
pkqX2cKgIfcPM9p39x7wJSMKtCv7sOQkU+3yxSXE4D5UrpdCU+J/HxtA0KLDa6x9
82uDGnZSyYPcJOUv3X6iSqC9xVE5WYRxMAc/yZnUAbx/7TAF8d5QXAa52VlHcP49
lxSBGI3RtoUFfaV+i2egeOV1GrigWuomGuFM8x8e0YJUkMb/IDzuXoFiXCOEYOF+
cSjVHtreeuboXcelW7s5LFD9hA6a22rcrrrY77X6s7foo43VRD6I2J4C61rUxloj
yxv9FZS4sSaIRSxQZIoNqh0J0FOztsgNDTOYp512j0NkZZUp+LpBx8U3xIWZvUAX
dY2TI4OwkKWIIKzx3CN9ldG+sDftMEysSrYd+aznZHVDpjLFopvFX4MiXxiDbqdV
Nipb1OhxpcBhNb8TGHAc173SpzU6qRyP2y5lpwTkrbNK/+hPwTPKgbHyWCHGpU2Y
ssB3H7JabRtskPnKWp/LYBvXOwy7genoUsQq1lgyPyVSqkUpMebEwjfBTMB1wwxK
xGJx4VNCf/mJdoBADGEkgGcw+3RMsDjD5sewC548MKjGPgvTJmQgNRZ1IOfrrt4r
+gGEeT6WM96q9UHJ3nKFl46XCpSaaxUMSQMgrTkqLbKko5WZx0+mECALxu9VjILp
hSQbl4a8KkhYzcYDRp1wne8NgOy5mtcOyuLx0F997xzl7mk/jG44WabtMJI1uTPN
cnZlzVIpZ6eAmuzr7tAROfXEU4ImkMz6eYThbnbxQ1n4FlhLtqYj8ZRMj5w/ePWD
XyVMFHSMGkfW4vkyq3mvBQfd0M6+r75C6z9b+5wxwx3/nY1mLLmu95QrQRK8DWxk
54wGqeSdNROQDJyfZzjlPta69WBd2DerSs3RC3VrQGahO6XsnJeDqU4AZjsLC8az
Co5JoQ540g/D4X0YjE+W9ERZCWHTWHB30LU5UiMTiuo6SocSRy+hsmZbeMvtVslq
5ACaW+GKDefw+t495+vn2r+aAU5WwMxyLz2hD3SFQ9WzwVmDE6NJjqy4l+czqV77
zcCdRPd7TJREhMb+RFAQsS+Pbpn+FxWGwPdEcJZLJHvDygwo5awFQxnkm6Gl5r37
7LwKSdBoNwnUsfoK+SsuI+GpJJOo7YDXHzwOJdSB5h6TIvaBR3v0+vZ4rU+uCk+7
ewD0zIxuvQ7lqgLO1ltcxpriOCmHWHH4ZiPEO2Y1oazXcL2mQJ5EQLoEpwrB5Fst
p6wooAAhYsbWj8DTQvTDgBXaT3t2cmnIk24py53qZHm6xYZGrelcn5s1gnkTGTij
lzvORjnvxS8Eghd/COc3gdYvwIhTv32QhD38sLN2CvSOIgNgHn3QVz247MyGxp3f
Jqabb/vZTrCNJM3H7Uk+2gHdKZmvxInwZODqFELMVbzkDPFsQKI4BqLIihTUwzAn
dmMUXBvyrqRpNDCHoGeIsoVbNYl0WJ1NZrpUch8Ry2GSSDO7tJP+/OlSR4kVcpAO
HRIbeuHEMIQMsojdRKnODUz8sgyC+8JjcNWPuD/n4uzfJuWgCHiqb0u9QNKRfsbK
hPXDtp2fG0jzKjm+MZX7PPwO/bZX5xsDyh3ycaxiZtfSpu/U5ssmmtjW/O0o2IVd
W9Y3VwG71gF/ZGr6HbyQuPvhtbBL9OVLwmYuES3k9ghfM3YAwHujnBIkhjkEzdjn
l7nTMbN7DgGrEQtO4ZjVLSa0spPLiDcaQwwJVkmgQkevOUoV5c9cV3WbIXkF04t/
KcYwukJwMR/hkUQSMu7rdQIoBybKb/eY4/dS69b37As8yd7jwoR9UwEbI7IgLF1K
1F7yYUMZN0L+jm/A2Or96sbsOeTDQp/i6V4z5tU4fqDfOEWIXwfEp/ZVVthdulhq
6ExrCA/QyfwOBcYq1UwwiQ9JSaC97sAoV71ZaPCJY5AiV6DqYgJDPX+MPdFHE0yl
aCsBxj8dnSBvO/q/Um2FcRcC5RQTCONNX8J1PME31xNM/83D0uKbVaOMUnElQEIM
Pnr4Jzhwyrjm8iaTdChy6TEpv4mz6xryU4tZ9lVOVNdyCy5j24gYa8rnzsOFKZ2o
jhAHA+KOUwRjyaMUDQBZklWId3k57q9FgNP67HKck2I8C+A8nzq0KGx7hKogchpa
8dnzI6EqzGuJbiG/qrJ3zYwbo+tRttkNB6OlmmqrhMflaoX+1aCWi5hqbSL7sNJ3
5j/SWPQbvwrKqWPSuQDjQCoSeHQ1Beyf071WFHYEs7Iw6wLDpWRimRH2Y8iBSmmD
aZu9e/Yv2ZrrfgE/ehLup1rbl6ggSs3bYx4u7BDBy9WqiNlp7fCpgLJjUP7B4ILr
SAke19rCzS/AeP+XB6L8uPiGUJU37g4mvpZoulDvtDqQLIozSAszY/fLJ6T2a2Gr
652eygqriOpvohXmckn9kqcNL7Dw4z6XcjVsTyrilKaNl+o4q2crSZxuD7mVao9R
VTgPZ/mjTecAtJUkBXvmjLFle8woCKbL0HtF04fzujyegGdfJ8RfIyOsrN3vEaAj
KzmWkDH4wfIAmzEuVyXCd13Cz7222VVsfRzO1V7nfWahxykgG2HSd3g8Smf54au9
+oMes01h9RELMmAu5DJ4by9pbetkPtrYSrGzHNw4zH1+OAKr6Pp3NSGPnsDlCP8W
kcbb3d2bGBJvR52kN/d+nKSfWQP7El9FVl/TNqeq1aekzOu0255scOYKGEWrX0em
xyBezlUaHrNYPREoVWUrJ3lAvruzpjPXQn8ktLSTDSCR4jMm78dyN/DswAvlxepL
TXEoWlmTBxbL82VgkF+nYdak3dgmaUeW394cNw/Um+30Yoq4UOwhcpDldbS7s71u
e/RPA8ngX/dBpjP+ykNlxNHDTF+zVXA/qhoIxn8YFmmAdIZXEBHsEj2zEObwZmnT
CIJbC6JEwD42icm7PUxKbFKUzyKWwCxjAWneIN5HdquGtjVYERjpQIckVc8jUJ4V
oZBWc67D1r8g0Y31Cax1rhMJoE0Lj3PAtpxroaMPtq75y5pPznUA628d5U/t7DTj
OiZ1INZNPiHMV+GdddJCcGxjvXhtQiZ4JIntsmGrhsvwS/xVQ0SFCUSXeNbOE02g
OWnpNChQhLllfi+IglGsxp7P/39y8nN+vXMdqDonyQE/3JBxEEY6DgeAzZPVf+AZ
ZW20XHgUNCd3CgePvFMpTealrKSAVHa8DgipHLH7Fhc1tjAQl6vuyWZW2wgTiz4l
VLP26Z8hN0+ILlPsbWrdzBh52Q7yU6VbtPExrt9awOEfOuXzONErl+7rJHrb3niV
4G8uGeWaFFhG0dLRh+VzSGoyhZAmnRrvLr01D2swwZ3mrbupHSe3Fi3Qq2wAlHZ8
K+lzN9ZBPPYuPsAUrqt2VzzSrGFnN6DqpBl0pU0x1eDtRNFxSaQR7vZnsPVM/9wg
TV1Z6NmeuZNMPIZGFq8M1dLomnjKaw4GepkDkhyqVkx2GZsdLCKZ8MOYVC2v6olC
tQ1qSzHlT4+U73rRQ5obCVepZ7axKSYO46ARgR5g8a9Dam+5CJ+Bo5f1oroaFZHX
EvTJHEX3Fzc67aeSsegI//QkvuppsnLgOYxKdsrGWlcbIpTXYbX0hZFZZnKKl0+6
iyllR2KhcXXD+Jke6kPHo3W7gltvPGaGLIQPi/EM4mRoQQs5sso64v3aF7ya217U
7ynXWnG36BdtqCQcDW6Zryy5V0208xbr+PnS0eEI0WoxJiOpAZrCbGnmOLABHe/Z
b6z0lsbDb/c1WeO/L+SLtNpmj4Vb1pc0NRF4FiLpXrXAaHt/TrjBkQpP4z0Yhkyf
qVO7JKkKthiIZpmX00p0jxQ9tIjTe9ki2NdtQrK4yOZPXHZ3tIBqLk95bqoc44PS
Na7zKmS9JjVEcN2BR+8VAehUoNglEngcmilSytcK4vI581yu4FgOljRQ+ODkl2g3
x3oi3lBWHA4AUb6P5HtWzQEef2aPiAh8g2au6k3YINr4H7XcCkJDG7kJlq1G3PKX
Acr/YSjcI7eOk2JmACetk3uNOjCSOJ6yiLRHGaRxq0eGDK5UeUp1kKEBrwNzEwHV
siquFwY2xxbIBJln8MGSw5hdD8uXRD7NQ7CKFmiKliEpf6jH23ni9XMS2eUGF/LW
hkb/LgWdj6jhdDwvJV/8IXUwh8XDxIb2CdEOtU4YVVsXPs0gZs9oPRPq28hjD6LC
FGN4sJIVq/ytrTwe1VBvSaJdceEwxJLrVR6ti6fRbHQBmlhyR9KH+45ccgWCK70u
RYOOEu39zUEDG/Ya7FcCvAfpiK5s4fNoaC6fh1PQiYkLmmNV6IgT3YLNtcq3RhHy
rLH6HnGbQN/QHgIsWPy+83l4/vpo9lLym2hH+ckiCaiJ2w1UoX8NG/gGdNot6hsA
vw+DdSOhL1+t0EXkjM/q2N30ZWk+oXdUyJu5n54Uv5VKrouxjKnmUwhu35nJ5EOQ
Q3AJFIj6e1P9lEQAP6XUuV8thzPy5TS8oB4+uLdG3EYn9Lch0uycNxV0aSoCuxWQ
2B99+wD0LCwDvjw1XgTm/AiLKTzQDtam/kgLIW1+naBzeCeM/Fo89MIsuclC0E8O
63NBHUydjGr5lGws4JDjLLnqCZLjOeOmRkaE3xT8CNydI862/17vqGXYzsaNI32h
eDBjqmH5myReNjfpitYlEYYRowx9JmUrpA5utle2hHgLl9edmJVz6YElNZ/GkC5i
5eRyXz9ICMycZ6IF43BX2Te8v6vbdqlXKBeKbwfNJ+TW4ooRCxIHorkHF3I40d/J
ESqQ2ytHdjcXtTpYqGZyxFh1osBdjf16u8lPwIFbCy5YV2tJZEuW6tbiMBmwby4Y
McNkhHVptdMKDCGW91MrtkMmW1CZ4XnWBrpbzuAL31V0h4fAnggvavuFpAz8ClCg
mJpnLLjIMEualtm/MFxg9725EktUXMxUYxrjnzc7EosmECZzKUC6Wx1g8AreZhQ9
5qdYjOfJuQNCap0pWEo3CDhczsQ9PBn3a0se0YLn9s8ZRZ+HuzXJcHISdokVW2jV
mM5OK1Tq6lFI/7ZyauDMhyTt/6ti7fBG0WaZBJ8OQgT5DODfK98UsS6hoQ/zKN/e
RbKfeA1fYFZt2mi8qLByU+tqAOt7B1nIL/yLjgWmix1VBLZyJ74N6Ix4wjAqrVkg
EXKsO9eKsm6sUZN5dOCVt86OcpenAggDh6dBXT0Gy8V14ZmL44ZJSBYORT46tA8y
B0ZpTMfVW9ozb536kBzLhopQ4uSsy+rA8thsvJSKfyuPOfEsgx75yGRiCuOLh332
J0Bb781Po0d0VAUtVQUgRyt6kviRBSsy/31/KRUm4Kh2hK2pE0eZcTSqL0D1qNS5
RDqm6pq3vkVpB2pnI74OX3q0A4JpZzn7eJJw+YXdorIanYsCZU9OZVRjFVdeYMfu
zwXYJFcB/E1LO1M1i28LEaPVZpgizU/6uyjgNKwxNQFdkR2jTyX/aPg0NRZ0NZPG
JmggbIN+tue8wZiWzHPPWt5BWOiGippOSF1bqTbaOtl/5H59f4gff/guTRIsrgPM
22KkOet2laDwOp81EIJnuJI6cwQtcTYN5rgrjQekpd/Dh/hsMdHJUgp9hUk/mzIl
jjQNOYtFBdRi094CiQRxfnJRAlVMD3gVngvoiR6vUO7+c6L5A2o4fpf3ndMv0cV4
uJrGuKBwag7vNlnfuve9/MUrJaOcRwyfwJW8+zeUzEppDkJ8xeUEnFY+IzqdF7eH
ED4b0FmgZGb6cyaowAu6M8qI6b2vEmIzha2eqg70Kb6ZrzmDCljeczbnAiHq3k8g
lfemXMAY2PAEd2itYVIASgFJArDL0zrS8dOS9iaW+B/dOVO5oU2cK3ulFX/4qqe5
F92tIhdlVdIm0cN/TrcLhxYQ92NV+J7oclehxYkuMztEzBevsS0m6lXSr1JL0mer
icNFaU4qoXfWitQAULH8CEJ3BOPVEEvUIIIEYfxxLtRYsYDDDSYyME01+HI6z1Be
JK9SQRms4F8yYKA4HpWR/+a2bJwmyqDk55lQ5+jULiQpB9Lynq3guX3pUFPOzqnI
0Zuj5OHsHr5UnDU/KzJ+BERz2ZByRQWwWw55mg36/BIHWaQGlKBVHHwxbxELiKhF
SlHjp53kC92cOMFmEPqDHcjqth5Kg3k5vFX/B0ASaGQTmNDJh2TQ7qY0x8RyAWR8
qGsUQhLPVRhBy89ATguvna/Q/ekJmMCcG9ncjWDDJGvvH6VPIpIx+2ovj3ff4fOM
pWDWZvaUNqcyvJg0dzUzY4s3NZ4RwD30fokbfq7RYzxFdDbj3dDhn8lE0OfT4fJH
em/J+2kWLYiHKxjokuKhpiUdZzVuVF1WzPkOt3GtZysMD/WoXJqHh8xtp72hv7Hq
xIQgF/Fi3ymeKIYN79UWPeAH9yzKjz2YAiKZuCd4c94yOxHPniWDO4pn1TUbND2C
uJ8I8Kj8fgMI+l05KCNiq7jLx+Oh9H5vvth6LadXy0GCByNXVIEsfa4U3XCeumF6
GJXpBTT9QO8g/u4QSUE2T1wzaQvBf6adcuOOeTGvv+fTtsBdC8oRIVnI3oIJGzVx
2VhgAxqay9Otnkr2ElyjPczLFORmbuFcA0oSGKEDZ8nOn7iA7YbasXi8LFIAPwXr
3tg9YZrM91CWd+nCg5oSDvQd9ECJfkVzTGltd3ZK/Gelwums7OJBWhnjY0FrpmXI
OnA/pHCzWTDJr5xadDT8OOe3YAU6te38v2sEsfZDhfXdisepJJ83UdVO8B6k7yCu
5GORtyA3+f3KEcQJOnDHO+wAUGKTGffcsKwXpyUjjnvefhknx1jzf1gpZCGv/JNh
VouEic5zvQqG3EvW9gnYJaG97FZLsH3WgWk5wn3yC+Lmm8NZ3PC3foTBHALS3u1A
LmX2UWOB+9nwLD0wTCKUwzuUAHQX0ZLVI2+7uHDTC4e+Vv+jgS03E0Ah/24EiwSk
1FP2iINY759eij6DU4+LXrK6rQ7HkShD7dRAgiCcPVQ8Bwptr2NVVMb2pMgjJjoN
Thc7pig06CoPq3bE1X1jZV+vaNGvtkwixe6zusUm/isfO6e1DzqAmhTfeAuDkbN0
2QswORk/v7ALa0Dt+Cql4o7b2ZFbKfatAlVGZ2WwfA/2qj+kNdRfOa7qYPGrI+r5
gyOxK/UgFrjN+brITXkhp77KNOtt9DP7oUif1PC+XzdJe363rrdC3eQvQp63CMht
papUhVgr+D0z7xe0LEMU/PoP+f5esFrXx6ViTWbTh7HvyA5Q2brLF6yWsCGYwQmO
xvB/1es/Uhh8z1/aDAeCsWf+h2IdjwhC164Tm85Aq5u+AT9PsLrCXLM7sosMAIwa
nMDVhFZ0y9QgSZ5Mcpqy2IFMZhiKlz6qvdjQxg6pYYw6FmYev5DmKl49cT7Xb1oS
jyjrS+NLw4INnnOXLhPhg8dpcgRLgrm0T1jZw4eUZYFgdbMTmj3YCnJCm3PX9tSs
kvfgdyy2JM1rl0cC7Ku0BZ5AKzQ0c+sU/KoK+/2JolV5nM5Wj2yfI0u6FxCIs5TH
7t+S3dcAi2RsUAxZS4MT7LMkHDs/CJq1/SYM+S/CX5D0WffNiCLYf2e62M/vzhNz
3ulAFvncEWt1X4EGgsleFHO5yROc1oZWiWY73oF/sTY/r5N+XBVmmzpYYEUatMVw
5q+HAgeZTh/HfrWJasPyFirsFtKIUGZBFRYUyU9NvSY4ZXOeY4gsaCtO7haa3Ot9
kslAbpFuCpP8dVa8TiZP40UDePB+0Iloxl9/j19FzjHJ6+S+SI9ciQ8e/0EQkNuo
KvnQrnXlUOtL14X+lBX0ac9bX8sUb65T7VaS+qDmlA/Eg8VL1LHsTIFtZPqWSnx5
v+t6Ynkoryr0NMcvobkMR1utn2HmXRmE0VfzFjnYV9mBdPCY0zaK09bezcgv+js4
bXNVGtknkYV0R0ul58I283BGC333BMBImBirMUcabuDl2aspVtYzx21JB5vbOz76
+3YVfoSoTXy84lvMaIzE6A42+vdxgo8tDBBdt9mLLJKeMQ02Qi4Yj8Xxh0c1df6o
NhCW7edf47SxUsSc8Qeugy7eGEW1mB9hAjTmEwFgq/v4emXdEDPYVh/tHoBQss2C
IyGuHZ+luEpLeTihUX3ykalop6ntgjbi8w5E9O7rq/3O50vYfafvVRjkP7v0Btes
5PaonETrt1xj6BHs+aEi2USwRSW3Q/2s4SoO4v7Xufcjo6U6zf8CicjcjO+W+aXm
3PySGOF92akuYuZBDwMs5lXLisj+Mjjxypsmo8SLFKVNfVNHuCoam09MiUOLFnyb
M/Vu6VvKYHRZsu8b7dnyA20wFz3GjtTdZV/9NNt8gwOjxYbFOwbTmAEY6U16e5JX
fjmFxxHHeYaj9k7oY9vUFTbPJ7/9JyxO+zLzxUMkvSXHz0TZ58eVyMNWfLJ7SM2y
luJMsdg4AW4DqclzLMUaBx7v7LLTyVOXv40tyCIAbXUdWUwdpHK46xbAcXlhcr9f
qFKlUnG77F4rRV8JpKfA5j6HxiWwCQ16M+JtfxMBy57L3gLGk7a1XPEiJCV9uVfM
buzpZ2AHiqJJ5Baz0U5YUL/SQCs11orKOZd9JuzwST5xqCidZLq4mgCoattRGKBm
3XaomnPmBwmIce4LV5wP1NSFRx92GyLmRLG3oq7OPMzPqRHjcZU7gA6HigK70vf6
fKzw6rnTDmCi0BAfgYGOBjKl1bX2wYlYwjRYDxssHu6szig8A4Tb6trdRp0+DKh9
o1NkFcdydpXAQNIOZ76GBIu0r2o0oYxaph27KjjQrdBezy1xGf2TsjWAQjfzxlMG
YFgAQ1wdWIT5sHe3jNYnDbuZ4ZWdtwP+Tus1QdRPZNsR1jECMgJmgdPMXiTF9e/M
RZVQbC1fT5v80cWJjSrof4T72TVFzX1yw0m4EvU7LBGWQjWWX8ZH+M5V37O7X8Pe
nbixrna7fQgdPi+nyHlOUg7CCD12j8C7cMqNhmDPz4iTdyjpviyQXiyAq0eFuq9V
vx+hHAJ6bzKzyke/JlG160hI454hSE1qZzX8XxnPaC0dFMyURn8ejBVSGSOpm9Xx
YaLSzI5OpQhRBVeNuHvJBC49csCnT34rA9+oNanf1uSK8yTScJxfBE52vzefO8sw
JkBkbL4gJZBRmqj3wq/fiQ3PVqztxTG6PqCyyptlk/0U/TV1/hNfqtiZDylXIADp
42cODDkVjnfLaqQCmsOmBtmVhli/4l4uzDgYt0NZXT5H2KENsDKEIDNJ7OGca8fu
y2wex+h1AsDkJy16C4TKHymtQ886eDyCR3vfuvFJcHkG/u+rHGSre6Vj2RKh2ree
IrrVPI6Rmi5yqINrHJuNcageVcL99lAhl6axD/J2pWVL3nbPXK5wc98xoR1qDDUw
6N+8rdl8A/XNgMl3b2gxeDUE100WDgFF6b9mQb0qI643eXiTrKV+K/I1g9BXw6EX
On4MCXK0f9jEczbACnydbQ9vJZSEVvbyqQVn+FdUNWfZ1uec9tSn0TTa1tP+rXYQ
HDX6qEmM3yz/4HcjI3MvpcKEL0cMeWJ36+g6K7qx9F5nPdqp+MZKjT0Y9D5nyGYs
EQm5xn3xxm/GMsg6Ut0hYekB96ygcvoKQveWeBG1cmCx+2RotL+qpYYBSPodK3iI
4eSpj9kuRXH7uWiLqqghVe1ACATDuqT9jYrbzbGEdfgOBCYKsknjyrJ1g9Yd1YnA
om7jHRq2dWazm5QVNhwdxAOzGQsh4+3Cx78cWrUg1fcFuRMKfyEvfNm+MYwRG1cx
7frPZMM2maYzfNO1jWhHzmRqM1YfTVTp+4TbgQc1wQ/KRqiw0ps51YJ6Mxn9o9Lv
DU0ninXTUQpRun/DYQxtlZM+xpDNHWPXDG2LB+yDdvMhm5rkp3tckyDRx3Srctgj
Yqaoh3hdsNlM8ag9jqWFs2IrPQyujG6r+fPoIvOWdER2OCP0zZ3irtuusMK8TOxx
i+ME+ygoX4+xs8Ev2Cnci2FEb4Huln/lyt4LbsNM9uAIRko607JwCoQE+XuW+jZ2
gB46/SZ4MNqPsq+AF4eXG/WmiLGoxybf96QKRUQbbqW1PrLjRL4g26CyckJNX0J8
s0Ojj2xiqm29W/IggVxz8ChhWZcb3qcqQt7nlqyzlBaChx8B/FanMYG0NqQbetPs
v1UI1CLjkzVfgjciWHQXqD1SJg8ftwRLvdWUikkgI9pakMhgaNrI1V6DX4YXXqTY
DXIfkAOhUdzEi+Voj5T8Snyk0wy9tVTYG3pqcG2PiFDiXfSH4TYrhcyVC+2NTtiA
y4jXzgViYjCF4OD5gO/+5P+/E93cQSHP106OjLKeyNTUr3EBpvHFj1LQ/aRrjFLp
WbpZHc6Y5tEc58l+io7W1i7gXVOnY101jT3yZlHmky2bmEyMwoDzNNIhBELSlbEC
cp37SDSlcy8UStcGKPfW/I0bD5z2PHe9Ywjgz8ZdPIYYPNCX8gRhAb6Qrp7Q4uHP
lZ96SaDX9kkO93ZWhUTJf4E+wl+lZt3Y5ZgOkZxQOrhcII8Xg205tZRzCDcqgiQF
4qcWFqUnx01hSCpbqqJEE2KFyE8ZvMSYXzZ2bfxZDFa+trCxCoX6pqRBj9KlDyfr
jAqX5HjqDiVeIh10SDEzhQH3a2FxjPF1POYr7O1CvPGCL1T+RvzbICevPsQvQdMz
7QTkNShUydBEO/D1VOpaUDkONFsr06qGxVhxj75IP4RGv9821CmnTFkYZwFXGGSG
v+D4AwSe5YObU+CNkQrv+YVJBPk+o5B4WghiO90KboP2votA4D6HJa3oGjvXsHCK
Lc6DjxlvlvbNALRolYhz4kzwP32cQ8Uar2992Y65ngC41GH6AVRW9JveNacQhert
0sN8uBOYZuAn6vgSUD2jsBt4a/zxEmvoKnGYHLLw9jL6r9kE1WB4vrfJkJ8XQKqi
qj8PE2SPlsxZ5dF5IxPHJiYnQvlCT3zupA1DrMuci1V61UFP5pxh/PgDHuEdbzps
8PKdeJrGKXWkQD34W78PDW1lgMjQiOPFDc+BXNFjOO/R8QDMh6qGKofyhyc3erXn
RryrzHQmq1PZWKKYzqBKYBXtRAv6r2bQCeIP3fAzEltcGeKFix5XcsESxYCJCEKE
Jx0pZGeUfvnj+TKc4nBu4MXy8SkPXyQsBzxHP3gZOAM07+hiOyJBt3Y+71kAZYuQ
u4Vi4ZB3wDQhMvW6moRMb5CNzsRXQffIgufJEsNcvcppEKAjhiV6ufPIp+1FML+x
Yca9wcA4MGJdv1dDBPzNqV7oQecYVOKliXe/3qdf4hVOAPlZdp0OsJHimcrrT6YD
6qrbpaOrY4urTcuQbfFnS969VquNZ17Xf5V2kHxq5AEQk7K8yM5qNkFuYFeLz0WZ
0pUbM4oYEEpufeqlmyjvHwYYPkQvzWVpZoKQn5vTwuUScyHjGK74dp5M26w7a3cN
RCqDUxLMQ2RqY+WwvhsbAxEIgiPpjkVkHoYVuUyFxqd3jLnSM9Wfjux5eQAp/r0Y
sbHOaA3mUqJOvEp3weNDpVTjaapb3Jm0u5z2Ns9yPBACgSSyJNp11+z7MJ2wHPAy
NO02zQrxLaloPMbZeXCk+KJTnymmwOaAzyzZlaDyHrTlbNQ7Uj92wjDc9hXstie4
T3n8SJGv8yevm7/B1XsoT9TOSuDusLFH0B0RRZR7Wgz/xJOqZdio2prJbI3oWoKj
Xb1Ua+zIlA9fHOw5C2SjvpRWVZmOT1YSQli1tkXlB/e1sloBXR11sdChZGVqlt/v
yBQlXv8kVeZA0fg3DFClWg65VYmEWcf7taNAeQs3kBX7k/IM6gqVAWQW1Myvk9Uy
C+AQWrcLY05rgpB5/BOWJ+RRlXSeOeJQEPrT7Zg5K9mk/dtTYKDt7LDXyGYQDg3o
VMitcLdU0/+xhU6fKVCSQl60buu1Eiq/udI2qg+2d1AJPdpMdqEjrKXJdBWUkKN+
BeMkAPoPXaLJMkln7g03KhIO5eB+W+/NX00UtdHFb8a8H6z0moNPm4oRPdarpo7p
NyHTj41LtrevHGMFRI+aZ/A6cZAKfe3aUi1Uvs5WvIdnqOFievms7TzUf3PwR3ZC
ep3ev1W3gXJspAu8WQ82X7OyrXh5ch4E42mBZ8qqhXYMQ0RAOdlVj/jrvsY/XI+v
sZCYyCUhsmYhCNlIGq49KXBABfg+UOLiS32Pleqt/jk1eI9nzKGmjVaqxq0ER8qI
0oTJ5mqSvxbnOJ73oenx3rEKI7d5GDH+3/aUpWKZUNC99pe1vrZftXQzFLJOaV2X
zlWiFMzfbjoHumql1Pc1buMna9DEpMsx1OAOdFSMQ83Z7ZWcCHM1IhocAD+2TOlo
Xy3rGL3aSz45728aoZdQmA5BIN2+CejO3ez5AmYEuzIwR1FBInY09Vdzkombn2Ac
1B+jbGoagNEcgRy9YbQfZtA3HlY+6UbtEeS0TYlSwIlTzb51S6McQaqygxvXSQOQ
w1KepL3TwyuG7fXvOJ1u9cjTWS1aS94jo/0Kk9N+HL+0k5/zgORq8uHagz+htS1j
gXBKvkrhdUmdXSvRhApqzitTneoGtS+Te8bwdEtTE83OpeRqzZ1YIRV7naLabsq+
PEESvu3heAyrtYjflJshjqh1SIvoSlNqvvXmoALHKTWu4ewPvqnWOonmA8hxiG0Z
gi5rRNLf7p4pWduEUMB3cg2i39OhTtTAi3Rnqwol41u1PDmvIjR/kGd+4wa0bRO+
bmhE9ZFP8rN+NeZEFCBwOK0vMQenuHqqwf1vk9xZHNZU8c+503rLvsa2ko8EPVi3
hx9N7hVGqCDT41cjtqSNJQDPhwH+MwmIzlSRdVdUWAydwgagf8PNle0ya3+W5ac6
/GYEVOrgpTVgWJFJ/bkLj+YZiH7nZn88Wn1zwuD8ZK4W9E4NQYbhNHcXesxLo7o5
VirawB9IgRsAVYVwOIk1otNpOuV4iDuoO+eUeIA1fr7Vv1IKvhrTEjODTY8ZVR8Y
SmbTMYHPtpjgdmVmuk/lbY+gsrFteDPOfVR6qXsSre18djbFQXe9FPhsQWlRskcm
P6t63TD/MrAgu91OcsfnkSo7GEBvWRJ5NyOW4B+zU5hZPZ6Ux0F/qCpgBcL9LOpo
VBPio8J0jEmlr5oLuR76PpuYu2l3O5Xha8DhPctwZ5fx/GDzSdWU7HxWZqVzf2GM
iNj1fOz27o9DgtL2PxCSmn9ECZKbkdKJtfmCB8Ngm8tNz6ivSH00nC+tlUH9wCeY
68PChCcIvuJTX+mtHdsGhp4jiRkAtSa8b9kjlbezT/3Ksj8gy+HSnwsI1MRd+olE
RuPXSqCnvdj4pJ92u342hDERumIxmqV4GyZshDXC7oma5yqsaqr2Cg7we9kCcKdY
MeoT/3wQw5pZPySIRz/qDp3aUHgakOLaPJjIREInQULeOlIiDKSSupwndxhz7qaD
MKUCfA+45kytyTZyVK6KiX9QIAZpskPEqw7E7JbcLDduQ8xmwPX6ifimIN6pVLE0
OyBUzXHCQ/42BWIMcEA0jOunY1jADduEcBDLAcDbXs5jJ1OGvpkLfLp7FV1pQ/B+
z2CX/Lq67atyhxNAfh+QOgDqJCwmST3kagHytqqRW/hgZS9dxNDo/r75yzA4orjQ
vrWtxVX8Vp7HPIX2TObGi8B8JcMFcVOvLArMIQytEy8Bs8fl2mta9zv6gD4nd6nE
D8KFXSxSnSUpADd2YENDBac+KvO1lk0qGtpmlYf9wWA2zPChThlRK+bmASS8uKHf
tTAcjZkgjTQ0hdbaTiXIfA5/xZDc2tRjy1T2EmoLr9xQVqL5dTWWCqMltTlhjnVo
2DQZ1WtgDdGJcsI7sj4gfd1pEJkCHRb7Jsm5Z2zGEYmfCM2LV1NzsZX8TqrX1b0F
Slcuvi8RteCJtaW3UFpAsaK0JyyVZXizZphn0FSrnpkXekayYSJ9kM7n51389rF8
qk5SaLq/196GRBZ64posqDtOpsQwrxgI7sZv03W3w9WHHWubjRMiecTTPj2lAM6+
ZGSiQymXbXxSVhrrM5WDrf/jdHQptQHUKG/lB/JSj/ouOA1CF3OGLN4qeeS4ZXSS
7jyE8d0KKrauVMxZAmg5wRlh03hFQmnX1TFbia9WQSPFZB/3t3eaPufZoj8SPWvy
k2PRDi2m825R/fLjUtvDBYzSSTxDequC0t2XWtqAirEgeOBVaxiCYUpnuGd/qzZ+
ZiNP3GCEI18yUgjjAnCX6w5sEDrKjF3A+kYYl5321FpQmbTGZMa9UdPyxdGlkad9
+hQLQLkyb095vgc3PCU8OVhbMn1GU4pa6NjleC9IippEeq5JEvcSygpnU0jWvgBy
fULij6GspIdy17TNn1tarLiJ7qehDtMPf5dMrAMexCPFefKes5O4sgsTZQpuQyGD
2p1IDt+5p1oDJXR6GUYiOL5VlomNBqY+jca8kZsTHaoWGmjC5BEPO86+nRjW2mrd
+FUoBrT0ognYsUHfRlhbv5sKsLwDa/tlBVIJf35QPZww89ntdD0TuWwi8X6ufPzY
ECl/FXr/IoukofLwB23z/0kd7LLI5yBvZKh2N87+eGblHU8j1SkdnqYbdYzCNl3k
2SsNtzCcHC5EfEMfd+bLIL/OIlq54UrOVacfoeRBDso4hgTrbTKkvqQXrZkuqiCB
lpsZGXlI0IHzUyEtxro0WAf2pf+mLCzRJ4tgRjfZFda929WCJitiGFP24cbAeTs1
a+svI42A8tX4WSMfe+BXHMRnt6ETx+Arw9mLL8dIDYmOJAOt1kKkzCy0toisxAvo
mrQwrqD7UUfCN/vfrLhS9ZWGWpdJmhFV2hJ43ZPiRgpgLmgbRjt8MMpfhsr9P4tb
eqAOboCBJKvJTPcmAvDpfthWOkCfXvdrWztjXwU35OgaX/vknyv1SUjK+i+EwQfA
Vi6u6aws00tqO7gLrxMhnCjsnL94FanEeEs24+wlMKPGwZR6ZGe0h6kAagTuB0/Z
9qK+bb6GmntSMJSexMPgJcwVYQKBgMTon8U0zOqHJ/iHu/i+SSLnaLKpcUwFdxqn
4Bes5HiZu369vVxpEDL4MgUFZZk/EjJ3PdmASVlCwiROPpO5cTBtITW9foBZ5Jnm
tor7c0dtnJOmsKchPREj8x2z3uBnb0jT8WOIFyua3yT8ENcjP4OQBssFVnfZBVcF
IYQ2jGHr+2RyMR3mwcCPeVB1JZbkfH/NcWGXIEf6Eu7kSnS+5nDGSY4lA/I6mdyA
vk9DFPcnoULuXfIPnH+9U7+QDdYPaUbYWL9mAiHPDxXS3SdhiCmvatsEvn7id+Rb
vp2aO6SwYPkrHVGOUbhAqbdPSVaRzIs79afo07F0TCln26N7RVCEz1x9AepMSYmF
Dl/QfJtfqujwfEbceVTnnLzjQ3HpeinYyU7du1XxjokuLrmQI/5HSV1g0Amsxe1O
6REjIrxPi6OQ3+GP//F9c7bZMJynXKrS09+9DEOG4hRvi+FMP86TdnXDiQ3mGCaz
q3YdtPyKlcsCM2Nog/o1WomnhJgM6yg1kPnFZbL4RNUH/xd4u6z//A66Sx1V8OEL
ecoVUQOK5YR8YaHWipPbVfg5mpffhjmNePFqt2KqwMaY38z/OAs1Bw3uhD7tu1yw
YB8hvBoit/eZq2MC86pdjCxj/7Ux9M71FWosWPB0w4hdxX9s+NkYOoKnguQP0pmF
pLe7X0v0T5xkk2U5ZqYwDIAxhiBWtSax6hwF0ZUk11W3DSo2s/ZSQAQUzegEenTL
bWu8iFrA5AIuZQYzJ1ZooGD/olX4G3R83DYXqYh/Xa6He2wbzMRSFK+oazXY4W0C
7LVoK4N1ZJ7JEXZEXr1tV7xCcBBoJqaQqvs8/f5Awpw/elLihn3WBWCzOHpxI0yi
95fownFCogPXIcubTVqr8NZm0oPMhv83NY/DUB0yJSSd9Hw+Sf9gjCuF2Hi7MIYN
sSPiwyxV0G8X050y+JlQCNA2ghecf5S0FMFckx7aefl+UGIKj53kfWyE7AZxsmqH
Bzp4zL0sDMMM159UVXk4hBgsOr/XV8mQk6SM3FhNWk+mSI8mnDnivkQY0WHQSCjx
x8FV41Q07bVNk+/xfLFeksrflAxXhxPWMMo2lI8Q23E5qMe9USO4acs/FkBf/ovO
GP9XhM7CSbs8UJqoCVYXjqNkRestTKBWNw1KUcH0kpxm8NVGfE/5DqcnFYMcvPnp
AqZHD6qhVz7l5KGz9J2m+U4IuI+Gd20yBrsleLxajufOyutqBnuPucOFSoWlzYmn
QTggWWkg/CtGsEEkTJ1mschVymeE84D4y88PVK9mH2ZQ3HKiq7kZ6NfU+LdJm7/j
plr4BsjzLjhKCaZej3Q6yBRd5sDsXt/pY29FqmFVxCIwBzoX/AZ5FlyVjdDI4Ojx
jhH4pbYuGv4XhSZNpfh4WjcaWwVRmiaNrYpOPqoBOHA6e9pDgkjPTzJRLY/zPauV
zYtpm0svZkNeIIexSZwELBQjLMK/XdhjmaKbruTmHsYwZ3uj9IZbnmChNQgakFsc
0Imp2jfRr2QXlffWvfzvO4ef4W3YSnLTCxWL/fJRLBAbZRR9UaCqnI4LTcKB0vLT
ZAXNSZ41CytjfG3CMrjC2CiLzE0sdLMJGKXt4xaI1QPV72+F2fp1zgTE6PMqUBR8
Xy1UYPAbnI21WySFHhdKK7+V1CfK5lm3uaNkMHMHnF0ie+xdo7mo1a7UEkvy2jWz
H45He+VY0jXjDUwA0kbOro+Hja28IubOSszN8mcC8GAt+6q1KDwUIJVu6KqPJUXi
N51pDCcZfN8irFcXMQY83NM0h6G3bqyuRjtXssKhSFFX1SIuVyx3fdZ7BcXZS9dB
0VwTDNvHS4QgXBEixCtqk3eiPjCoaBJOlWRsM/+SfOKQMjZGV1pmZdHJVWVOhsKm
gLLUzyMwin53iQNmoYhukZK74g3Sj4yG4yqhxonozGvEbxx2adM1wkxhd7c3iefm
0yx2YRL4cqdVTv9tEw/pZ4WIOMQEwcnP1Mwp/ssL2uzl16Bm0oPLQVHZ1cxKrtp9
LtYIxeC399/aiXUfpNaT3B3VQUHQ9+IgVodffXudoyL3u7SzzhkhHNVoCJSghfd7
lmOzGwdKf6vEj/FgI9EGponL6JViyCN1rP+wVUwL48bRBbnsPUHXqVZ8173LUt1z
FmQyLw+JBKMhgXLGzQuP/5EiCrCuyHYhnoz8+sduARPGeyEB1BWizezEOCJc2N6Y
ZBi0OwEB2DBAk1I3HhuGKPXU9KRR4/+gmj+iwBPDddtRpVfnqDQ1r6uawOqAbsNS
c0QeY7K/1WpRKfbSCRESIfHwRDGS1YTOYLgLRbxOK/i5rnCpg+5mrfm6madq57Bx
sTnXI8stHcfosJTZYtSnb4m2fXrPR/dFCKy+fVwZKLvhgUrWpWfUz/a4+nsmn4lM
z3UM9FOZtvbCEO5mT7f551lAEJCyx3G4Mhkb14ErIFjUJaQUykCl3nvG/7Xt23Ab
SCuLSr+VgWDG11KsXYB+sv+dxLUGaD+cHKg1odqfOQcZKZOBufxDSZbhN06nimmm
2Rk4J+5Y0RsiKlSpYRE/BZrL3ual8vSHtj4EOqrWLHcNf0ypJBMv0iQA2huvVILL
lYewofjduFUYlubkRMgic6+oTC2JxRi7ev2sIkqdBHXB6nwTIfmFRbZhlx1YjLVf
uQL5sPc8wIY8+Bi9R2mhP/faHTQwB8MXkIZv6rYBmJnia3vewF8o31nUC6O26rXo
F16+9B+S+4ztaQFUtbfEJ6RA/9L46FT2Jnkmx2LHAA9BfwX6NA4ENpbeovbK5vPe
+YB+pQ0OvDQVXopYBFuDG6ey16VGqL2uzv8+fN5o8zZDeQ8OAsY508F2N8f1NsGN
6FRMTg8AFnqpNvfLet74ULRzlXsoKmfml2V69ZaJ5vZEvBlcIMlnAwuHI8Sh1A0I
aSiBM8XuLYXNT/IGZuAUQeq5bj5sBduLb1qDQ6cbflJgLeYe608yAFveQmDRM9B5
ROrIGvGWqOUXMCAkQT7lHyzhGPU6B7QLj66Rmim8IQKyyg2S2QB1V17D/zuXSaRX
vI+A3NoBkzlTynhbVu4xQeOLXgdqBXCeNUp/QnjTs/Wj1VEm0mDSkfV+yB+0cFUY
bR2GeOms9H3I1fkJavsRFFRj2PWqRPHvhp4H4ACBlQ3uZcT4OPlFjtgIb/GXpjMj
EAsnlZSSxo2qechwPCECJFsSp7tQj0lrhgqKAzHGAnZjJDYxHIJsm1dJU32GL89D
/oCUyYWTeIiJi/JFLq8FELlU5WZqRMjcKeHSk3mIvJNiEtKAgrHLiOVYb6vtK5bY
fFVm/SouYFzjIomuIlGT+y9dXAHRldUZ06cHQFYYBFjXFqtGyt8ABwCdGNFsMLX2
R8ny+RORDyEkUlndWZRqUuU4tBw8UHB6bRG01c6NZynTbU+D+ia/60kw3655r6qc
A321m784SMvh0FdMGhS3m0Nq4GyChE18EQw2AtgXbTq7kCvNVFSm1a4vy+Q2JqS2
H6uFjcTUMrGGSo6otk2JD9vpIXHnk3FqGipNRPuy1MJTZKeH+/FJhTIdRwGU/heg
5I58W91eQvGU53nWGccfwD4sFYG79Z8sWV169zNBNCWghtCPlvBA+hrzVfwxY4Sx
eNKFcGC0tJNvUYwd4zAkCfgMgZMci51Hc6Nc/QWvjw/l1kfKYGI06KfkfpWF9GwZ
hAZHQxeEMK+aKd157KcnQyDLD19UxArDprJJ1VD1CXCDLfuIko/jhbZ3qgE/YHeZ
DO3Jbgmcfk7l9hLsZV/xBoS6EXNyVYgy/0ym9+UjEZhICEcnZ33sdVsHy4i5y3+K
K8oW3L52cmboPyNn9xHen7ZXE1PdwrY0P//BhnbzuaXuHgn0hOptHVAczjZwLCnR
6gdj82jyJLKU+4O8NG3UIaEabo/fDWdxYDLI4rVnef1kKAYJnf3g67G9cLZyRBbn
d6PmjNThcLzQEpv81Le0PSUXYukHVHZxAoEMxpIfV8pHPaLcR3UmVOnv/6bsGRPa
lAigPv7Mx55/iRp9BM9EVuz5OGyN16wg/SjYkkfWpf2pl3UBzIfFsUbWRUBG8ESD
CQDCDsnc2Cg/Bc+BX5n74ttC6Hd4X8Y5BH7XnPhkYKWYqnc0VcxbSHmugoYQaaRJ
JQM2ahhZk73/zbYMiDcShyDVxbQXu8etpVb0ZNa0HNJxqZbvHtEAi9mCbEwDLrU6
ZUy+ZVySRnWyN/Pj5kOtimjqnt1OrWFxHpOdSz+heKOwabQBtfkubh9xV4F+kbVi
pJIgG09qoW8qZmeRJq877SZSLx1OriHtHHtNlOl1nSzoScttOihEMo2L2Pj/4EBT
m9URilotrAdm8k+npIqy8lR+bnMlDVVtmO9E/tLHPPPbjoGWP/6cF7C4ox2thMCF
nBC+ZmLGBFUVjeJ90WG8xpI8ApONUPaAAATN9+mwQicgo/0t/2DvaYuI/UAxnVlu
5pXo45qi1ecw9K9GSD77beHpInj1FfB8+S/xcQ4vopWBf26tW7Yv6xmbBcUH6AGf
Qdb5YcRFoIObIDWwp3dXeZfTx/YzFbMX3IsObqUWfByTXaDnVEWnc6MbivUGVwnv
copl+MdA6aI4a/VVwT0uJNV899CfMxtf/O6qx3zyEzFlALMVZD2iHCJDhsYE4CUN
B7aqsapVkp3uliCBGLEKWkqJDKPo2nrQTF85HAUxxagZVVQ/evaRY6PhVF1Q46Ob
Ds/RisjaWQOkro92DvOlw5UeHw3aPvw8KUKlHO+tnFDJTC5a4eo/Meak1W0HaxY3
Zu2RM9CfLV1rYy5OW1rwy867unh1JyABcbKXsBXlSNKnoUGUNFoGv3WKwT20ZGMF
L4I4Vgbv10ZknA55k2tFMwSn+55lasySIQGB61r4ZwlhgYH642v+C/IP+Tfl+jFX
dYRJRvZSjrtCklGARQzwqaYwHesWmBHpohIoOyUGJ3zza0km8JBVwTVmMpgeit9o
u2EUs32Xi8GPfKAcet+wC1uB75pMZ59KEeDl+OBMgal1GMu72e0lq4CtWJiI6dxu
gf+Pxovt+xRtJSAe344vc7WiHlSyyx1R4QljscxiiF1Y+xJNoQ7lbuKE9GsnTvly
9cv/pohn8DDeiM1rDhVy1JAYxvNjVIF8Qd6CbqYDGfCFSXtKszPi34zskVst4s/o
hKJCBFjhvI4NGfKT4/wv0wsV9yoiKrFxjwPPmS3LCuZu7o8+MkJsm8Hl9oPwZSQP
t8pHxhtt9klGVLC0Dt5hH3P9F+0eynRf+qktWiavgl35QjcAQqVYNLYIoFxYZP2E
C09YnPys0RzisZh6C64rENHKw6qakyI9h/2Fyi73ijukPiPEF/C9QW2fVw/GeWet
H65CgQf88T9U32dON/PizMPmwK7zheV9wnLvVvf1ARmFflHGr0zrnd/rLAyXeSnG
d7E84GvQYIjhkKk/9CfLtID+txjLnKSPlEmRsPA6uSXHagM457xThA+Me6dFctEr
rzbbVBNshknO7gONsu9c1ullOD2GYizPZ39fMVQdpEdWX/iQSbWOwrZQzwt+vsK5
Y0RO251WY/jA8IbX2yShPpCJ1A16MbWqq4MJGXSwQElAhEdVY2mOVE1wBpPhLwZA
zeGxmLi2ZFdoEW0xfLTDBkZvkYol11dpCtDl6B2eSzq3UAKkLwdIm4cYzL/O26bb
fIKaXUor2Hl+c76hpPYqvssdVZoQP4eGWiUjllGW42DpFNg/dvPpipUb75ioG/e0
EXwODKBCFN/8DKLXBQeHHVLBIuagNxTiSrVUtEkd4PXPxpsgx5Sp3q6tUVKrFsk8
FqueCoTL5gLcPksnIESonj1dXjGRfsxnOazT08LnUWnrjFxM/ftC+ArfB65LIvpD
u1bE1gfvqaPc4Blx1UBBxM5+0JHAdoezztyR7v1Ys4gbVTKCf14cmCTcqdJZ77ru
J2yqvconx3Bmbq9+LM6JeSbzYxf4beiNCEvIakuq68zLykkKBN7as0skX4IeAXpj
wD6er5buZxlg7WUxqsNg5zE4kvGUcjypvQvsSOMP1K0+/6dbm5UlLgfoGhUVsVZt
xGdWDkGOrnRgxVsK+qF+WMsNRwycWi7Y0wmCV81p68wcYF6xEONTa2YwfvK8VJ2x
cGIfw47BHvSqx3WM8WqdDgNpkXDut9CnMKhBKccIFBJvwewdVsYGBdH1sFDNjBBW
ykIrCnyneBO4cd8DBVVwHysDc1lkpG67tFSlH6K+ZXAGTk3IAAwPkp5icvtiy18H
ZTY0YD7sVg5rv9zbJAx7/y9CfXYPDuWKTHWa6XS/qzYond61I6M3cgmcHj1iXYSa
BdSPSclajQQ/5CieOa5PEpM6bU5TriprN/Kw2Wvs84OafYN28WIFS1OuJlpymvlb
bNS8cvtokwWFo455BeCHu668brY2wNK5b3IK5pZr3H+7lUVYrXDACN9Di0kPCea0
jwAPvk6ovvDeR67Jj80YngQhpQfmNwYoLzQBw8Z1TIhq7i1L4zMjDV+L3wQ5j6bY
Q+d3yyVaM5f9ksczHwH/BquA3Nda6zHqIbSWysPo+7sS//vWiv7Yl+DL71obIbcw
3gC3vtESZ3x9RLseEAJdXzzPHSqhe9u6mem+Qb21sghfut2/em9eF5GEn+MvPAuG
/Ip9dhyYhtBeWKANzmtJKU+YcjxD0RzoS/MgKFSqeUQEgduJwoYiC4/oFC4yBCbY
CLFBEEe6ZfyN1hDClVz++EKn3kpGO95K1ph2Ypdzz6I62cPVKwBuiWerzL4krcXF
Px7221+xd1WYe07qh+i7RhUEYqypCHRuq7izfTUsRzBat8dKDBEHE04mj16KkGdQ
MOH5TFzgVi4wk+BL4LxVcnu6oxDCSo4+mtdwaq0/FMRF9Le8KYQ7iHrVt/ublKHa
k9x1PF4rL+xn5yHxwGlr3OPjn9nMWcfyR2GZeizxGywDCwivx/FqqOJYHUMpoClc
EezWsPfq1LnCKPk3l/TiZzG6ilZMXazKYGBLLJTa3sFVFCMrfpVtVpGf3cCES1CC
ibKCnDBvrdNLZDYT6KlMzv4QfQmgwrK5ohhphgTiQP6IenU74g2qrbuh9uYp5wcy
Xwg0mM7edvtzToCJH78j8S1BuztsNp+46sDuX4/VfXg2jELd7RCT5XZBA/wwXbqj
q2p0VFy4578a7OuT3GtrYi1eLSOuqUenJ9fGBIS1BFibArXPPn9jMeF539KKpQaU
VoMvYaUDRMezMpkvfnTRM1YomN0t7oKF8E5nq7s+EYprlNl2tS6FXHcuOHRyTud4
wrvJO0rk94SLD0Tr8nnn2dDv9EQmAz5QU8h3G0npzG0Y4dULrBoYaN4Qn4tS7eTy
rnH3yrY2KxFI6F+XoKAVGhkQOdKNMgr29L07DFpJJQxMF9wRyOziVi1eJyak4oew
/PsVk/nq+RqIWciZ/wtJ3kiIM7cFML2tY4o+lfbE4H4U+CUnZxgz+pcQFa4bywpB
oDoot3thBLgIq6Z5usPWKcvC6ubskgp6ofQPr4BefaaC/RGhmd8CjsRtCyFjh4sq
cdDxtIczKwoKXRwSm9+usZ4PsFXLex2GiFnqXmIeHvXXSGGVCS+r8cDiqGLTzD78
Ynh/BSeKPihb2tZAIbvkexYYfh5vjTqG+2e0OzLDWUZnonJVGnjS8CKay/lgASd3
EyOEZWiTkWpHGwTTrCYObhcShEw3rsHQ+0gkn5BwtlOrxXQ6sj7SN1sSmoCshpZa
u/+LNN0POaykwDBThYcg0CNf9GGWn5mSiWV9Xpcme/x32W6Tthq57xWEMNUdR1Q2
Nz4r+yjm7U7o1ToKyUUq+jzR2HlZP7QJ+Qf9oZ29tW2YUR8IKa5LokmdcWvAsgdI
6my+H2IuYjCEcyxrd8VJstn6dFaX86/bQaLGGgHpNAX+WQCAGlZ/CnNTmMUYmOkh
vijCaAMj6G1hwa93Rbyy4r9Jq5xDr6XNNyqz+/2/6Mj9Op1sFlBh7SgUpNnXvJWZ
NlUScM7B20a1IDypbdJMddWHG5lExijCGCezo6qnjROOaRmpXOStKgDV7mFUIsvd
jSg4+dLGcxlp3VJ7YLDqW+E6it7t0svvrckJ9xuDeJSf5eBGHFAf9hyTtVyBmrTS
4ksNOP+Zam+Y3xt032EXuiVZ9hw89IFrbsJwv3xGrZwAPyucyo/C2s4hpmfRQ4hk
HDemj1eILit2FGyZvHJP4chBddWou6FpRZx2NB5/ZZDgUZ6w4KFrjlbK2OlMBpy5
pBbSh2yG58XG2YwZGWH6GUti1al+05+Od3MddHcSQqYC4slMpVLA2rwHZFK2w67Z
1AZR6DPEnHdOWB/uQiD4MR85SqPrYJOI9Udg4kVYJjVMzbJfVLejGYNWyhFDVdfi
hk9ewcnKqvQMvmxQSotldXtKyyehI62taQTkH/vDc23qYasIgplSjVqKtfmBA/pT
dtxm95qErwXN4/6rmn3YNmRjfHAl8ZzgpfdOtLhjgdT0V/Vns9YF8Gj7qdfro9cF
FS29N8F01wHxwkkGxt2Ug7nW862u//3OvgeHQ/J1jOYyndhmvzxV6vqmyTEF6M5q
/VPp8TqfTCTCiYhtOwy0gi+tfB0h5JpZQgQb3ufxC/VQ4894YChBl+nRxxkCT/Kk
NEILnQMDpfDA/bJdWjsQnYKuQwkRwvXVPqOFV8sU43xd6cnCTbIjwOGZsG1OH8MN
G0JleZZZ2tb3r5Q36JaGEj2Q3XxooGcAqDCfkltZ9F8T2o783TeY9NmbxHZSGSmw
f8B5SYdizPmZq7xAJzv4CmL9ZuQVkXAciuYgpny28b79QeXm6kIhhy5zmiBfBpmR
yXDvgwAmSxAD6LPm4hx+cXXFzgQquRrqmo1o8HP/3UcJRNXIqWYh6lgz/QjuMipH
OJJwoEqg9fjH3ir/EirQt8JB1uchnuFNPcmcwJc5l6C+gsG23B1Nuy56yPIIQkq7
xqyuhOG+4rQio+t823Nyrn6J20hm43JAWvZKmxDCNrsSpIoR/mBJwVORhnyC0fs+
f4q4A1pofxqMKP0D8yO9eO+MlEx9Lzj472+VqUP3sFepJX7FUqeHMsdU5gKpmGr9
5ZGzxBFAgPnnX/NnDqUu1u5gKLaodXJatY5sgEhqTTfLdmJ+ZkPY84V0dhoU657x
NK7awUIqtWX+iowK5qlFXCfJgncEPDx9K16kvmA4Z0+0rW6Fzc8rPBu0ETxGkZR3
D4qyvRP5FFYOyIm9pepnrMO+z7Nuz0nzrOhYByKHF/nVtKnUUznixl9OgIt+vTj8
DBpD9r+7Y2VCWjS+pjMkwmlQtrnj9kxegt4M/t9178suHrtpPkDH+ha2d0UJKG1M
qYSCtjQRbrvNRQOLyfJQYw9LADhRDeRrMcMtE7/PR+HOtvjGE8fPTbJPyG60zALn
SKgkLA2pl3NvYd4HteyMH+Dy7ZibAuverhVbUflVRaJ8gbHs29wzsSS2bAF678XX
LEgIPd2V/TgzcXKCVpgdut+Q7j+pcfau/4upZ2/t/4Vjflta5OTaIaSQKf/YQ/UM
jmcna0XZdopInT2d1ZUBp6aLg5SrNc8xQu1BVVyZ16rcnBtFewUV+YR1wuReAfhh
emJj6BSc4EYS34qYHBnb0Jhj2vZmCIufCe4uVwibt6CkZijNk//9lR1OyYGPuC2X
ZZIDv2N8zO/aLGdiB8uASCFoARCX8qdmC5ym524mGjvIWS9xKJ+6XJrCtq1AieFg
MxSVCAH4njBxdPi4bUTbbB8In9LrasAOyd17ITWSLOtL4J5JNHxOB4uDqpzvWqdR
JEdpu7cr9rbMLjOTi5+WHuV1vqD0TFkDDxGInfzPVaI0hS89nsSj9kf5ifSneDDU
wsRqY7J7ZHK89FauL/PmFjN7xpIg30mwsrJkDaJpd/i0aP+V720+9jPTh9MTzPte
SOh3Uy2Veq5QAEEFUthAJOOC97MWKZlYwzHkTSjOEI4ywZwWiiLZsNvAP24fU3DC
mKqGzAHvG1X9gHjyReAtdk8BxtCCNtDAP2puwua79MIdtWonPSPCBCSazOM7vaXd
E/zOcS7gsVkGdyhR682q6TfkmlHUbeZBth4dPjFZ/TLOlGWzFlDtYlGfq8EZr7QQ
s0asiWWpLgVQtkzI8lQfUxaHU2jFE9n3l6yZBdS4M5TsASJh362vOupEQb+Ch0ig
TxsXrR89bAD7g3T18mJ5Ly9cyCNQdoH6ZZuOvSL9mZ/O713whQw0YbtUb5GGMbEF
riRHJ1oxynjLbJVdVoWPYg4TfB7xl/7a15SMCldnJwgi5wF6zzq9HMDIFrGrnt7B
oflctoub9tjzDUzfHMLq2Zm6pQ2gGtOXcavz5DKsy7nNXo/MkTCLSD85uBRY86ex
N2Ds4RhzwCzKqyJuQGZMlkM1Rv9e4TPZAEcwjZAMettT2HKPhZiSe4jt6kvsyAzX
sMTvLcFoPxvU0sxazn3y4hMwMm4dZnZpEwzUAbex35GCl4rZoSZ94vdpQZWCxMo7
bK/GNJvf5SOmNudhFoG+2CYYDU0Wh50WhqRUQvy8UOSh8MOLst/8CqlmD5M4+mzV
sCWfFt5SCebt17A9+jwk+tEhZVb6HiLfl1l5vpvX9QelJt1I5mYr1nuPRrl4AFXS
dlqvD3o29UalCzSG9nP+xWp2j724zcmhY6JQX7jy4lKOjJH0+P2TebaPfFGml9AL
xcZ6u+rO9p9RuyglVsZGRruJDC7V4+x9NbTpdutTPELqEzuDbBpPOhq/tI1tFaxY
zZxm2N0UNYoW0E3JJB7s/J3nOpOfxE/B06zid0Sesp6UzNroTWiTwUPb6sc4nx6Z
w2nYa++BbtnsmkRKghlk1AuiNtASkAeDSETDB9vSAFcjYloYb3TiUzOfO2vmbryQ
hbP0BqN+t3/BjgEarQ2jSlN/etdKtzICxs0JWbxodNgpPU84GoVtoJyJFFgncrcn
Yoy8HxKsN/1kKfFaLVJ/Pmp9NjA9qLlns08s6bS0wA6YaRhyTyP2sejeTQpz/trO
OGhhQpC4ZScdbJuL/8fSNiXCME8D4IwJkhlzGFHL351tYTFlnJh67arucyZsGmJI
F9EAgePCXAuJFxJXnfNzCKHAHTLtE9ZvxxqiDoUZIe/II7vRKAFrXoyrKmMR+6AG
vh9xAHwM0eVXhgQQaxzL62wfrf8jRCrVGnXg5JYdqcWtdJTWBzT4G+V+l/J714ze
9Xm/0+rZNqt+AYCpbZChLrV54VHMuv9lj/HkaCT+CbrasSdisz9cvZ4hnDort9Zl
JysV3Fm4rvVY6g1fD0zJDfoMKSe+rqq/7fYOqbDkkKGZ0lzowfWZRJnW+P2B0ddD
56uvbPFa19WGGNFsPv9hOuVHOzOpqxsg/uTouiUPTl2gJBUDd0GkDtF946uIZ/Nj
kdJKzvTgfgVwd+u8guJ5aOr5pAU+s2rxydDWT6Z5LW9sN6lRXoHyb2SbX7bEL/15
m7LxFPww57+uBOPRCDMe37XBoJVUBolr0xvPnvU3Czh/13DgDNk9U+4Dj895njrb
wTrzB19Z02naESPg+3mdumdK/9e5D04DmLa6VdundZ9bXQgjc94IkEuX8ppoQO2N
Js7OQnrwGFaTZRpFtVhOCBdArUSDUi/GPySSj6d5d38RUgZcpIBEd3jjouI8J9ot
IEWO03OznT/0Rc8s1tHphY076IXVsfkIZ7q//Qos9DJQtehH4juQuekxH1J5thdi
zGU750PEJnZXqe3EsYz5p2E3lb8pIvEQo99p46nuAJ8+ggFguqZEIU37X4id8Y15
FIAtvfPOsyGVq60TuczhE0l22QT1yfRba03PXm53jcx5Oc2p/KtdwxW50Op5uG1C
IT1lkvSggrYsyMgLUZKmZXfpNjjc9FOP1xLca7PF+sDSFrFzgQqW4rKmzkM+YwYs
Xg0rmlPcCiLmNWiZ+tVZr1dTnNH8QaDsFHOFWfWaAfsRp1wGZofw4ezRKuh3rh+W
bI1FrduNklZchWLqUxc4r7FedFqLHmN11vLgjR8JKyWtkEzUyRtQYbxdjoj9KRmh
xLhng0vQ61lTt/0Il8Ky6kPClnFiJipZs9X9Ukl/HcxIbysGyTCz8MnUhfV4db2M
urpzLuM4VHOcJP2bfTLSC4B1KV2B7aT5yTGHheRFS1usHPkuiFkFxV2e630OcOyW
LjRDopah9XcGj5/YqBIXfs4WNStsdCo2lPzlIJiNrIinOcrbkKtppAZxHqxXBoOn
N8bvrqfrgzDBUBkADlmmemnvhUR6yi94ZkY5fQwaApeEmPrJUMAiGhTPjYmRuQYV
HP9pb+qoNCMiSmtmU95ItvYt91ZxS5G6rfFUQJkbR0xQEYDzyQZWYVvb+jjal8zP
J6IvxtvTnl/yr8LamOsW9yufZviQqhsMHqCMZF2E6RnU5eIsrO0TdBWjksWHWjxf
ilwFJJwpyb5sWB8GC51MxUXDPQay+RStFMQl1CcugGMtXOMq9KKd0cA3Xs6KEsRu
PbsSp3qEMCj2i7tR8oudmrcOdRpvVmSakVMe54Ij+QaoQ+sGh9UT28BijLHqlckX
uGkVS0tCoCqZlJnX/JgQ+xjbTIgWhJo+brj//YVzSukW3O+iJx69W2TtgYC2rmft
IxllCbGdWcJs+kVZDKLG1Gw2lBM9OyaZXiiSdi6KxolqqosUOLgR+1tRT9t4V7sB
C4ImjNHkdxeY9au1HaKX9jN/1isKNpe48BXli+ug36jtDZ09YLATD/NvwBohXScG
pnemmn398kHDQ776r+TCKAYus7LYno/dvy4Y+VfCpz3rgLkMMJcKDtMf1UwJ8Pd4
Yj5Pm3guhAZib4k59Hvf/AkTN5CKKZN9bP2rKVU/vt9ZqfDmkhnNn6HytKD7U/yf
FBd2QZwYvXy9VEz/tQ2WAixLb9wr7X+GZoCB3LPnCd2WL9tY2Ju5Zyn+dmwQirN/
+naVOB5HKIIcXRq74QR/9Dt99Si0LzLnbFcE4o915/seO8hwUc25e8gpA6bzmuRo
VmopbkYEAYv5FCdsNE47vPpJV0eOiqlNToJeOH4oppDrl79SXZTs47qTxqaCus/o
3QXjjLANOCyh0+rMGXPnCO9QRxVm2UWteBKztfEb57iE8Nyr/2nwxPI+iVLp3A7a
dXNtZ6Ui745/HlUqLtGQvzra0qZImKTaS7KewB+wH1OZDxEKaUOWgZ51Ct/abuOG
kpzPIKtowoCLJ6/FHU73S7IAO05h6reD9EiqhQgoYywBnnyrfSUnTm5p0hN7p1h2
UgFWu9K+VIAelf8DmVNQWsL2VfL9QDUVoqWP06Qhq1MGTPx8SBqUX+bKNS3RdjLM
6bXkQMvunI+jmy6fE47rENF9joGho8ui381X9aBhdwHTlsD2V4DR1bQ6gMAa86FX
pt4jncep+Dv+aVUuzSJObXFjpglgLg026rK9IXJnptBP9OMPQwJ2+1UXlmEa7DoI
dGT0smXZmOifmeRQ+0pRUzOEAFuaj9t56lg2h0P4E6cg4eDdsgN0dHLMKObA8T3p
NPdVgaXkwHmhcFvnCkpxYaU6v+szI9rinihpKUsFzw3nDjT1ov3VPjsAIAW0f447
lmLYuMF488UQIJp0msJsP2DjGMEl6neWeXc7yT9L2M8PcoR7mECi3m6LfYI+UOJe
2B/QXpvUka5BTdQVE5S+hrf0fLrCWT9H0k+WdhdKvPQQOrmUNDVTFjvhHXw8DW1Z
lhplf975NFjuoNuvx/wqFOGAD/6DuQmUBZ1RFruOBP3t+G5MOYa4JeesyD4zzHZw
SvuZVdoR6d2I9CbWa1pZUIcUWJBgVOr7MAkWWX/+kbaqB/MjPS0mA4bOhIBEKYw7
QdwMVovdZufcRglbiER2mddk9FSz9+FJ01ESXSAu9Bjb4AqZ/6rkcpO02LYEbbdu
8nxrIdsZmLZckeYlLTIipkIDQ5cl8qjaDb3tzr3HpAcMsBiJhpzRV6prGaI4rTPo
kdiRhVxnJJuR0A/XHBuL84q2aCfR05ihpv8l9YFCnoKoZemzVZsFo7UwS0acR5i8
iwKw4ckk02NWZvnRMAsoeaZ0J7TQvpgrweyqQyr4cxSym3u5WnJn9utbheRz/jRv
u08Xz5xFAKaMsCtTNwcXW/F7awHKT8C/MybP2j+NE8ZLyr6kKyHcUuYk6bEODuyd
/IpdWPMN2DMyUlFo4ivCdIwPByJwUMacBsCh26nmx91fpzugT0q7YR/nIHUPEyf9
Lqq1ACFQAkur2D0XPoF2cHQHnF4hul785f9pfI5Qf/EnZDNseqG5OOTtEA5NQ+AZ
N9V+ZX52KoCIHE+lvwYmUcJESYt67MYaoI+n3QJMgFeOXv/1TxBmnfzNtbjCrsH0
nMQ0++xX8Dp9ebwir1K+q7t0+G/oNzGSFlVUi7nAP0Z5SdfyJYS+UpUjAT1DVdqp
XdBtquPjGgwehc8YyCYjPotpkMsyPf9bCc2zAHhG5LaTKuTPu95WB4EBQu4MHpPR
1BAoWzjCsRj3+CQNbxDyXIjALuvYFcDeSOzYi3xGKszMxwX66dcbA7/20TTjMmzD
CaCbChwGAl6OS8qbM9JijEfR367D8NXr1RepOVDSL0Y9eslyBIi+HM/1OZTydOJ5
eN3kvDvp9r/DYlCO6MKH94tZhwUSP8i9YbQg3OxyTa4RnJAfBvHyfTSsWtr9bjy7
UYD881jN20YruxXgacCUlHVmO1AubUCDetMpnE0G2w651l1qgbXkq1un+JAdC9Mr
wi2SxTE6mnTjoYAxBd+OZm5TbNeoNQ9aZ1Yb4yH2qVrb9Xqixu29DRwtImpyTKED
myackonw2T+JARUksHsdGxIQPImdhb03esvLsIlI4E6QJu/lXet0jUcjqFiyqShY
k/GikNJ27HImF202JDIoEq3FolWiz5e6gVuX7pRRsSsz85J/hZF1veQkRbJQimxK
DK6CvcKlnRdd7D6K3cTlTSd6fESTpCRn5ip03i6IUS/aNZJDTeSbY2cfGnLG1GE0
9ziphsINNO5sjVYxORWvdPNsIcVQGf6F/yaO3zIO3Yez7sMsgeNmPsgqp/5ZFmI2
EQkL/hDb4vOA/5w8CWpqWxuQmd5ML9kHfA/eG/upD75nEw2jM03uVRYEvNRRkP4C
rwoEGhj7TOeJ6KRUYCYsBHB74BheB8lc9ZBuAoOalGv4zsLKK1KGn3aG0vp/IQrd
blOBqhpQUE8NlriQqRSprXmoj/EV6gnxP4A17k241VdIOW1frz8IEerIrk0sRS0c
CFHIYReOg9paIP0El28xD8ePw5m8DMQNCV2axP70SV+8Yo8Ez9LCjqyVWTx6pZoh
QEz3duZTOifrWJx2sVtgQYx9c7sRvLhawgo//KC3p5pqEtxHHYAEO5vSnpwsoEaq
Kpov6nEMo6L9EN4zYuDqw0p73udM1WPOFrLxXMwNbpAvXR89Gb1e7qYJETMlaFHa
b7YcthKqnh153cMZmjxonXb5UUQhxJqvzD3cOL1kH6sKEqENzcx6Z7AnVsIyhGeJ
aSzkSg5K6TPu6m46kVj6AiA/rrjdsWw+EvfXcpKpzkxcnLGrO9GoVsoMABqD5/Av
aYWRJfCwUqOZb5gHUyft3vxu6XAIqUp3wqt2HHxCmbK+WWhDkxYp+GOc2SGf4mnc
6WsY27u6vPdHd5Jp6na1sNowbyEd++9a0zPF1I9cpCVXqgagelesOVXb+idckKbz
Abw+lPyCmjcDM6b0Fai6u+dqxhmAjQlq93tK+1eX2oIzTxhZePnPDvBy/yRETmuy
viLL6WvSLHEm3C6uZilJuFQalMY/NY9VuhQg6/5cQ3wQtl2AkEzZ+u1oLwIYIJs3
AcJujQxJ9q9rhZXQ4wlVuoklmAZpeC1RvxnJWunpIKq3okQKkbjBRQQS9VKbnZ5v
VLIqhKXgX+HYEJ662JdHxOT2mAa9KMH8o6nRLgNVYmGrc5pqmK6C2qN0kC5a/3fS
C3RrCWNDh4mIvVEq7NXAgDECx4KTx/Q0WqOE9p5D987KEIfHGMwsAByyZJ+/xC3c
eLfD9AuCDTEYwgM5j9yz6UTpktsh5OidZ/Y+fokBQrGWVbPGUeDf/yZka/QW+ldd
lsrC1U87BKK8HJliajg7F1V528n7hwyieKWpnwCm0rsBkqOsqg/2La9dkPYv9JtW
Cb9aO/+IVGIaAdJSoEUH0rnL+EqDOsmJn6x+kFuAg9Ljja/ky5BEZO5xB4bzjRRn
m9jEld1n8Xl1CjbU21SmU0nOx53L29ABVo5IGEGclzsWAc8emVXE9COnEV43rftM
A3WJ8H7hKfQdNN2knf1A4/M5SwZRE2b4m/2/j6q6e+T6zoebf6NS37BbXTXfs1Oi
PFL3Cw8Wl8qj+o7L1AZwHQF897brFthZKt6v1wp8HC0D0uaQMzDa9ax3rALhBtYA
rEOYyDtTwaBs+i3cE0PMwPXS7aoS1sF7/LL2AC/1512zq3GFORxwHq8SpFmAEJeW
RZ3oe6yYFM7xpCQMvZS0y+zFaM2BuqLY8jK0uppHis5PF7xvZbjC9YNzC6MMfRxU
x5nY5HNvL7Jsqm2qaK2tHbuJil/RcXyCJqmD5ug5du63wlSA+Ny7JV1qYYpxfoZw
jcUbo7EUz+eDHZyIAavhilW4dSr/350IVCtmHI8IBc9vACHAMeJoJFtu7xefkQ6u
SlZrtPVwKCpEXUvEfI83c6RxcT7JLF5Ylvlbm9TCRYZm486QN2IyGUWCWlE8uTwP
DOZkooPS1eYhc36vZEYgDi8l4e2zndLuk3KzwBqSsBk11qYhhUBhWeBmKn3BW6ym
ZqGIl4pSlLbQn5KIdL2u9wnJayCLcn4N/8jTLUGfF2GxYJ8BuD2dxIzMpPzxW9bu
yyfttrJX/dpIyy69ct+Aw/EZGAk0WdmQg21Rin68Bdw8qEW6gB7/V0I8bXRsEkMK
+h/rCllXB4z+9duGNP7t7/zoFLSfnOS/33tdoPDbCCT/NV7J45RcmDpMPY7bexQU
Xyquzr/J2lfS2E3Mjs4DGFHH+XjuWZrgbXwfGe0sA94Tg1EPutjU+5J0oh8ZgtAw
nllUua7PV460cF054bpb3m851unU3id7ew652iwS4aVF/wBuncobR3DZS07zCaTx
KcCQBN+tMy9QIcTvykw9m0DmsCp89A4QxYccyDLeQyp939ginnc21eHI8vjqPw2d
VI2Jgz4b5ucWv4KKemgfjJHVtelH/eYwY8RroIgyo/5XiOtYiX1j5SniYrY45JWn
SWXI2dQiHEAGlPre7yKm2EVXWGYH0ldtJvODsWCLLB2YaE4+Xwg+ASeCEjup8k55
pemCYsGs3BjbByVamxTEHsDTAq55qleu/swKewMvzn98WXP3n8MEtzqWTC4SzyDI
Xgriz3HkaA5ZSBPFLGamasorCcB8kDw0fpEj6GkSj6udfnj5V5tSIfxSuq4/rZP3
/DX9NrbVuGmeFO9MQIFoeMi4Cbk6TzvSnZwPuOttuuCgGYKSeFk4XRd28ZTtF/dh
3KQrJR/l4So+YHUm0FaZf0jC+NKaBwhlQgmmEGGBWgvJFBEorxUJaHbEjXUXY0iV
MlHZdbPWHWESnDX/JGxcCbb690BIb2BjJsUai9zM1BMKlFUr3i86+r8FVO9eZrsw
4Y/El0/5XzFr7jcYz0B1rW7jwsMt2DH4nbL3S+0eRF6W2yTanTxqpqhb65376obo
ryF+HhBMP7at80z6JHwtBoyPyEM00ZLbROqfNWz55lOoILAK+DYKyPEf8wK2mnTW
LMXxCUyH0p1ZbStSiXvYU5ySonBbCIAVLutEcP553NUDOpxXpErEyeOYshmBO+mM
A+g3DO5NLCLbfGPBkzaQ7WSLgO5GamQ7QuSp1O5L67ojY1KkmUkU6h1F3fF9E/Yu
6g226qGThN3hr7g8/aBhx1rv+VCaBAQ2zx5hRA5KP4dbggdd1CZ2mNz7GZgvfz33
bxn7FRVXjVW9x/IIZBIgaKOe1IyKGnGRQnB3mKX3ahHpstfSghghhdFRQsrXq4D7
mSX2mAjFtmaSfuCC1fH2/Qjdtxq/FZ8eTkM3/sByjXJB5kNTdukRYrZXNUnaIAMU
NqmChwESRsa3QR5SdG2UXcsbPVG08N4Kjk81bTj2Z9Y/lto1zT9MRBgcOefeM1CS
xwh94w32SIrd3y9UOmmmmjkKNinCiVLK5UlitOFwowN9kCqVid14fPnN93tVN/xa
GWDXFtP8LWq6JRkrRoX+Rpp5j2OjUxGYma5M9vMK3f2nzl1mHe0DSZZJDQDZ0pu/
0EvvUZIUhOZQ8/jsj8XRHtLLnwK5PByPqLerMAEdqEyYdXG4gYbiEG64H5BElu+/
HEQ7XS07KkR8r0t4ROQGOeXKXEx0ctBodgnEbBw46d93zbOKD6gclITFWpzOLXKL
Gvt3qk5IdNaOq+lD9MwsTtHWGxKBU9+rXQ1S9/5fWTBEHWrtIa1K0y1JC9oaHe8Y
1nJbC4I6nL+ZPyc1tNGlCVyE3tLBt2jMrgfUUE4OYAurKtF2dP1v9BIQ5GG9+xc/
bvgjSON6rL/sHra11WN8ULJkavPUriHrZTLagVkoQD9XNLNb4fTIqPx+x2jPwSuK
h7faXZaDf4nC+N3cE1/Bp/pJRoABuOK9y5aPwLN8cb056W7K+elVYyk6KeSj5paY
iAOZclmVBEDaq3bY+9rUBW2RA6+a+6nMyU72gmXr4Nt9gCXMFZGY55PjCu1LAxyc
rGj+oKh9ytlfoZobZ2UGe6+xUpgQgTDc8nDAtPoiaN3gRqT9wp6W1PA+35VYhfZb
Av5nzr13WL7NWDv5MQY5BNmO4k0wvaRwhVKMvyZ+8jZVqwd9/fljaONSywPFE9W7
l6Ke2oM9s20KFRYVeQ98OuRpYBspQPS19Z+RLZTQUeqzi9ZQ3G0GM3YJwn5tVCLe
LtaIDxHyxk5e62D7mWqpyIQmgwfOYe37IbP5d7fuFnWNlAgcPatlZpHdvoz9tp64
deacxsmgDf6RABk+bh79GfwqFl28W51zPmI6PGaL1JygmDtM3gvAgZ9mS+b1V4/u
+jKrHyLv3jCBy39lBKeqdqFnId7Jw3aKGR+WBNN3ugYwzy/r8VoUttOWz3cc1NzR
+HsMTgYPGWFDMTvaMY4H6FzKtNtUU+kUFG8zT/7w1YNzkf1zIvhBpt6GtLcX5xuB
hpyJ7B0yXwy9A7sSC8G+i8KfLnRqXeLMnPxF0L6cs0yZRU3pgQ6uiCfT9cMBAzSL
Qf9ZEuX18TxeQLrpmczK8DSHPmcRr9potW2RLnBMZmHuEUoUAwvemUhTMBASU0ak
ykLeJiS3RistGJFpyvAQh9gMTTM1kfev6VOeUmIXOaIKJmYZ7r3Q7TJ7oYOpBP7h
OYkB/raqusTKyFK9D7CTTZ3GwBDYYX9SWN9nlgJLtGlA2BfMikFo1fShZipPwI2d
zuY7+Dj9j81XBrwZEdej0n32JTz657LKpsfhFWhct0c2wUaal+GMw0aIxABf9+Yf
tH8k6w74q52xaWIgdbHhtUiu+2VhxAOlAPZYUnERhSQ5SFAPN2c6Ri6ODPuldF19
QQ8KyeJUMLziQ/Ko5EKkMEQNuOgUIVkr3ruao69iSqRGftM2IBME374EKetRkkrw
1PCxwifJzZ/K5+CryNVBmAC1EcjYQWm2dacfywjn+D6dv0VuV1iEq7Fdseu0Ombx
j6CllIzM62R/WPQGFEz3DKqZm6N+mKL0B2q0eKAGo8PH3Pt10ijb1Td0sO+Kbz8y
7vYVlcZswtuJUwuRRwrWL8NxT0T9jFPLTR7Ou1BtcUeoSxtB0Mry3OuSUeo5nTuV
jJc8VncuftdaDOcqttRA23BSe4EJ12r5dKyIpQ3lb5b8WnSGpSQ1JXem14xyUCve
/elXTyJLKbyQAzJ0iFy/1b3hHF1JV+aOMr+7OPvtgiBh6akidPgE7ivgytq4Mc5s
1DIG3OqUb3bsx82Wkpm33V7iML/OhnDKpoJIRZwJKe8HPUWKxZraNIw3pAmPOrC8
w0rMf7si99JnzmbgQ/ak58AMYhWFFNYM0AkTrNg2F7geMU/jjAykRR2mVzTciN/8
7QOVCd08AyEv07JsCpiq0Ewqi7RazB7Vu+/XCfaX1v/hGjnIWVv3KEKddZNRocq3
wp0XF4ksyJJOA5+vZHDyFrYx5KYcnsuDZaOSGNXNOAPgpq/PYUsus9n/KfKJxuCy
oCHSHKXw2tIm0+zwPzZem0jxKNooKO6s1x4dm9K82jGqNjmyYDnRu2Kz7p7s5NWy
8ILwvFRmDF5i3w4uCI9iA3CyfeW5Qs79sfyTmSDU3llcw0VI1z68O0h7e2bRNq7Y
HkZ8OrThu920lH6jRLUFfg7doetnnILaDaWyfN0F+FeLb05xRkCB+QgGAfaVqsi5
x+YMFESnd+t82iT1+TDG0krLBJU20OWtSYaaDmda0chuVJ1axvBoUg5hu/YwZzkz
0kOTUWM//puAjptb4Exm9Vtgt3vBhG8UPibFIN+Ofkujmmptbka1mvFiO6GF1bkn
0KNmb7fTMFI5BgtSRDG1vthpGCnToUUN0bmO1Bl8cN3lCTZOYhuv+jqs0ON/whES
yFx/SAoZJ048zH5F0dKnuluMVH0rbpipZpAfJko1WjP7DalA/PsSkIda62Ue7ktA
V9x4xJGH8ERoXYGji025oWKixdtnQYR8hJQgKtv4z8w9AvKqV7Bk6IhwxAxqEytR
PToZi6pDuLZ4QToalkIIBtF6Ue1k7klBrWWdnW8TzHL6wIVKjRzVRhJoq70SlOy0
arWxt9eQZr9lrvBuf19ZVwnFbBtChLBI4cGm6m1bCnl80lYVAgoKFenelWFeIiMa
1OgnPuhMU8xn6csyLYRMN4FxizTG1sq0Gj1WzmteoyHnDdBB2QMVnYDgACTBZQek
JFfGqAxeyFJl7Aaq/96bAHfMDMYhWEO70AgLl4s46/scZIP1qpuiHcUaRh2k/beE
vtTIGcJ+CY5m1CCuVlWuNUwDsZB7/1yMdZOps/LV565lxEQ4TfDrYySMgA/jJF3p
8c/HlH8H3ZIhB+3B/njteJmUVj6Cmi0WjP1lx0QT5uQaqUSzK2rrSCKOT2bOgCRl
NxpzqkLTdWxnJq+lmMjwzEwDzguFE0NCsqCzptCrryjXBqpYR9Oo30hI62d7t9/7
FkBNlW4/hJa1ofkovlSxEhxciXOcZzfJKKh2Wy8rOCjmAHn2XfxAxtdxCqL2+/wB
Pmez36AkEgrRWbmT8/6HdIlkR9aYQPxcjTDwPlu+kJdd08cGCWWim1ZBhQd/802p
8YJGunp46g1idY5NFEcPzNXycMFmy4crqWUieBaxrgGwrh4Hbem69/VeAShREU/x
BreaqkJuL+LhVJhFBY72o8kiZ5+Q/8u8az2FAxykPwDu2x4kD0VhfEBxAYOdjRWe
haPn7b054f06ZJXeH+ncLOA1UD4NGxMM9d4Q0QHjWBEq1Zb38JqEBs8zsYn/BWAe
+QMH1ZOUzEMNdTuyFnp2UwvF2Igjm/ZoDMJzXADJgzBog3tjciFbDI5Mxe4GVuwQ
zaw40FzrDkH7px4quEPo03G5crUBaEekaJnQhYNDt9gLoV75BBALsmYDqWfAPKxE
/qN7zTf3Ok1uoSDAxcJYcXjGIH73OroQKaT8kzHEIsE04qGKtUkQWcFNKH7N5cJ7
PSx4yfRD2kEpXUCPkPmjafGiM+V8C/+FGPgGZcm4lVKTR9OjQ3yJSdcSjgB+HDcw
ivmk8bbhX9CTJsRuBBoPRO2+PZG/PfUaMOyqupqZDo6mgnUaTUkztiaOZ5IVxVWr
xnYyXCFDymKBsbkSQ49Tcix959mjKLPw5aizcBeW9PvudYZ1487hCORUI0p5F76O
TBbd77EOOufUST9gr30v1ORqtzmPRcfP9l3K7KisyhwDE1gaj/R1Lz9RDfwFP99F
cG9pai+2JeIp34O3vejogrqzJ41DOVdvUroAdt9EHWjzhkxX5ZNDw0e5nrqR8aJh
O0kVdxdYYE+w8CRSk8iO1bAlR+7lmE/khs7rZRrZrKsvDXb7Wv+8+j40dORfm5Mb
rf0dU6PmkW9tJ9Px0ycFp0nFSt9qzJSOk4ZndmPTonQpq29nf52Tw5LMUjnX3sO0
vLp/GbalLrNSPIsaJyOt484Bf8np7KYoDq9wsVb7sBng0ckHvm4eiji5oNGmIFSL
6O8NX0rywKkbEap9FRmhd6Czdfs4Gbkuw7N2HWpB/UGeDpDe2a2Wm6eJJT8n7Cir
ZtEpbM/pxzIwhPEJBmaxmIq2qOcjns4hFo7CR2v2wpwu1Ur38ncxg+hdSSdtLd/H
+xVrqHhra5ga6E0bwYeTOZqSV1Y3C/8JALcnWCpYfda2rMUOcwQ2OVE1XR6H1aSD
ZnNncB+CPVmAs0jHvaBBrAsGsFUtEQ/kRJSkMop7MFLUCZkqpjGShFAAFJs08O0q
xihyokq4U4ghOC1+5kMFZJQnwBF+LK2GQWPimlF/7Q42plREH/iXhkfrryFc9jeZ
ZNZMtI7ffzrtkfsqwqIL0xgRWCeoRm5qLLxUVUW6MdyeRiPw3sHcp5235THeH6i8
EQjOiE4JYXXpRqvBPf80nThykvtueqyhMAgHWgFD+ieb0qdtznDg2vq4amRcHhPI
141DS3dHlaAfKQ6yXRB3mUdFfaIk67uPpEmc6OUCDWjplTdD0sM2T4HpBtj0a7K7
nmkq3by04jZ9Qr8ouQOnG2wfus7x40QvFFoU2i3AJmwZShq0kDHqjIMjcp5OIgdk
/pKKKmtgZiDUgd1xXf1uvLW7OoT0/af9On7tPJiHSbguAzV9KK0HSzOzlV6DcIuv
16OOFRa/Wukj1si+WXwIUVZQJMFpBwpa3uy/YC2rbY/0sck1Lepv7HDtGFtL0h03
Neem3bcqnUrPYo7pmFK0ej/8yYG4rv0DgleRc5dq3NFFmAzBN0LvMxQhvkS0RD2i
0K9IMx0o7RfflkKxFoKll7os4xEuAQoSrnkWO52qszuYtgvFh8hxV8fjOvie7z0n
ru3xWA1IjMQOplcCXZRqBWpSNZsSYB4zHk5Kwdl8/l7qvxZ9CvWeZxPIV9dI5MEn
RAn94yLY3uWeKkCGeSQdNXhd0NcyygSUdph66GQ4Ufq2Xnr02qBwIj6RyAQ2sAkZ
8rAdqCYVAszPlhagQg+8E68Q36ciZnKE8Hz2poBgT+yeCpJpIQ/NSBhSuX6e66g8
y6ljBTKZ1f9b8ipEHL12OkM7KmsnQ4gH+C+5sqXpVrvKZAzP5pNGF4TvXw8S/X+e
7DpNEUMgN+1etlk4/M8+bWk2ccVIr8HTzLEsx4qLuLgeK//pw2IZIZpTFwZ+/qnX
4bplf0XWgp4rbcZdrZ6WLLvyytpMpHaSxsqiRpMoW8K3rBxFjHr7KH5RfXqOpweX
rnrT45/iXsXwY7OlvysYnMuThGkp2l3+HPhzdYD78+yphCW6Vb5JBPy4HPRwyiic
cSioTvfYRHpbT/AEUWvA2u1XGCqIz00XM4rbPXcIpCo1RhUvCVgYHYFQTkbigoAs
ZK+ghsBCHbHV2lpo5Qlu+XyWLh+YQl7IrDVuFbqFarBN6hnWBOUu30i5vjnPRbqw
1RsePgo/6uCYjFma0r38v2uREgoFr+1DrQwTcNy8q4ch5Ei9CHstbSrUI2Im6laT
62JZuETk+N8TEP2O2imt+gMozz03PD2CMTMhYQV9Eu0TRsj3oEAuKLbCkCvfeTNi
I9F9YfLb1pydi+rQUfdvk7ZOIf7OK7r/PnqAD79vhrSWgj7zdFaIWFcjnP5QEMI2
KJH9IhgoABedGBdI3p13/IaOG8raLgJSm84gWeawirXocKIzY5VLf78DPeLn1FKA
qSaN0GVJEuv75csW8KFszmaY5bxQ9C4SS7utf+T4RcYTTCj14ZgOjxxCyy8yecI6
kI6T8N5z0FQCph/CLNUCv3Te5fsjuwgmXIRkp5taGrmhhz8v3jORClrUtCfmkLYi
kzUdrXWFVoeOWPzec3goRVR8J2fTbGoOR0GBAaWmWAJzxe2DhGSGly3JbtBurmVv
VWQy6xad51dtezdkmfwnJXVswMH3ytAeA16w7CJUwEtrJhrDQWhgPWIVqiASRwPw
E/BWU6F3xfzBrJZdP7CBtB/ok7yDxl6MALcmkXz0GsLfCOdQbD01U1Kia6+GvTBC
u8buhE8ZCn5sxKYgUgTrvgl5Xjezn8PDSjUdoq0lUIEuIj9v616yDRRvXhaM4dsu
MyUZbv+mVDPlqIdNIJKcycZplZ4mmT4tEUBMiCHftoDQ9OQhhzhquLCO4s7CM4zZ
OqnYjnrhVlNr25ftCyEsyPeEwN2RkwZZxBWoYLeppO1TA9iiHtGrqdoXEodZ7uVB
4y3M/nKXFiXpuiMaCuobkhyn5Gc5xXfIYrtyCt6zODprfBsjagrF8ItwDCwPnGqq
NIZbkH2DxO7Dd7VHkix59R5GjbN2CrpJCZb7hmwC/ubC/xeOoPuSxGEnChAxegaS
FqaPWEaV5fNM7QjQfikbAyUMfK70lBhRr2tjJs8EHs6r2gImE3TG0MiAD3bYfW09
QXR81Ft0/qqNUpuEO5jBWanmfKKsdQ+37Ioco39yUNE8Bh71q0u9vw1FDwn15fr7
+P29EeW/3P4/qlMlUFy/+N2pCmDsv7Hs2/Fj5SAXQgQg+2vYQoru6dS9W06ttVkf
gBAZUMjqTbJCzWPOt7qm5iwYfMzNIHINYWo6ABiqf2GvgBddF2oOt3T+6kBDVaKT
jBZ+DGfqsFTwYOS/0dNyZ/T505y7HGWacrFOsUsPeyBFQkrPUY23PQGfz1resgIA
wfNUL60PCrWn1WmHgxH2dxKaelnz6uO+1jqKhWRU0En95od4XXCHUcu8PfWwG89a
216dd9p6yVt/IP78MbChL/DQCImfvVaNKmsKzNUOrb9YpXb/RUFKeRaGbIcmAk+k
hi7RIKq3oAxAHb3oAZEZw2cGi42owZGAx4jbNfYUbWoVWIPfi9nXl5YIXirIWP6a
ctV/mRldZP8gzLvzM972R9/5XEgJAQLBAbzwdeWxwGWmMgnalLaio5KuyzW5s10D
AsSjsgRyJdbJNTtsa9ROVswDf/E9HIWA7+rWB60gCHk9JTYvfwER+6BWTh9UckuI
zSsCU0XtYqHQPlUjwc1h6yRi/o8uUunOGmHGLk/UKCRPH6lrlK1A8m/u72J+6Tz5
AuiOI9n94yT5/oB/MKY0h3zskhu/MvSKhY2UAuEaEG3qg4r8MKRsWYYWroruNwbC
GK9T6GBqAw2sEGUKtumrXqrd2abWmc6vKGI+hNg/7+kRYcK3xbE2uAWqdhoCThM4
q7IR0iS130ggu12ulZO8n3BfB7m0gDs9jcjT3C/HUU/3zdsjmHIdxNKGqfgjsxVd
10XH/56NaL2Sc+1csxW/Pn99YlsH/QH2JWRuXPrbufwZ+GPnAX5P+frNXDFVn06o
zSakKq0aLF2aoL8qXBXh1XQhODO/KzuA34NJovIby3atv3NEMPvde0z4UNEGXA1B
2e3M19yGgatxsuOM/iboispZKNgMCJt+RiTPOmmaaPRhfv/wKS10YUvTPKaZ0A6T
HduCLd0urnItfh0k2LmBB1cqbfDiASoALdWoNXL1y4kUONnoseMn8OoYAF4MKLW6
FmsD+UhZ/KjkIVsRwDLfstFKpqN388VTT6sgGlYY2v83Ej66OuGhFUj4neWwBac9
Xi/ai5QcE7Zj3kGEC1yNCzWvaLph8GABBtBSk0WqyP/7+wGlWtSH++8rciCHcCUP
eu09KpYrT/mxTAZQpYZIB503Hwn/NsINXtdUQkvpamLKD0yAV1r99SPler7Sms7X
FiyDdSYS+fwGY+bzVEkBkZcTFlgLMJ1QDaVF4ItUhtYRP8Uz8rSamYJbEpyFFMa7
5mJFvq6YDY/xXl7qibGoEMETpkdM6+6awkj3VoAZZkdbjL8timj9YuS7vRC8KoE3
5kQlNiPXSdNQePW/HuEc1TR8+vKsFNYkBXcD0srBVCbiv6xOjxLXonbjSgtBjXwy
kUd1cdW0EdLx/+h6N+rcxah3AppVl+0EUmqhj1eA8yljw2QpOBpM/wqy91Vd0yGl
rjvBE9T8QnouWOOXlpBdNDDmFUHVTm0CSjLBWcy7sY/SnH+7fWAGS2A+keAruJxl
6r5b3yKaucSRPajNqP/yUah7CiTcyEBWWzylLAX8ft+vvc9KVsKPdQJh7+r3+Sw6
3ZyNEh3DJ0YWEpFZhQSiI/gGlJ9QBRI/M6OeO+s548eIAXhQTQB5eX3jvLMVOqmt
lwyZFZihkgF548wci0d9FUGYhZFzVAZCkPSpANGV8q809pAEx2jqiwcezyqWkRR3
KO+7W5tBGainf5mbf8FWCe7VfyhR8QmDwOrNoLsfLh/2ZEAiN+L3vgkCgIJPoeCd
uWIDjttNU/tYrRSTs0byK1pBjaO2iAPRltR0wS85UlXLx0puiM69+mAgzVxPD5qE
iHyJIMM96tL4I41F1oftwka7gjIoFMe5xrRTKDaznF5KIDsAHattSrTNI8433UrW
XJPpOlPd/Kh0h+FrixSoW/gRY2TmWZg0RMORYT7mVTni+dQ3mCw/lROwK5NXCmSK
2YdXJpM2x24ibjrYQHpeiMOzxAwDYkTNwoTa9nxnZoPodxdSmjhrhhgtpOEhnpS4
plAWqlSLiBj/LLRKw6uLs97ggOhzstoswiDPuc/NF2smeaDhyfQglJEshVRWJ3zK
jGWTo9LVdqnZwWnluhzKOq7Tck9eK3WiPJaDikLGC1OJTKp9FJwQw+SAB97glP22
XMYomT74WEwprABgsf4xt1EP1PeamL7W6IrZLp5GCghXmZnjMeBRsXvjW6nXp4vP
7vuTtZc2LVIc/9a6cwQyo9Iz4FmeK9QHvenrKeS1NHn5SZYmQu8CWoFZMqHXFvIz
SCVUIkKBLm/psnmG2INYJx9C/pk/MlhEDht3SMlhs+ut1ANv9hKTC67dLNpmflgJ
Rt1DrJVZy7T53L6p5FR6tww6OuGyTN0EzVl67sf+7N1SFZe6wPwK264rJ4rEBUET
OpuyO7SzDm30AyAHBrE07JN5rmo5h0j/ARIM9byLSaSkoqpIZK0GNzZbfDeoQzu3
37Y25/OB/GlYisOEqrM3MFsQKWXXF5x3FlRkqtfPngruCJEIKeg2WeOGr/iW6huM
toANddUgPjeoKVyu2FqK+z4uAPD+JWhwsEQC64NzodcSmmgMtq2RN8Bflw0Yuoxq
YMNERiatz9kwUyEMurqM3rOJN0ywcm4Nmm0ps+2S1T26acx16aKhHSgqFZ8bXgWm
ScoDp7ndHwHiQOt+FTCnJ/nlo2lmyXQDCoa/D0NAn+nG1AhzdHJHm+ti3NMlz3Rk
pIyuFDFYfwt8q7evvSKpsdxGcUhvcae/qmX1xGL9r9KNWTOcxmNhtKmQd3soQUFx
ZPvozrFu/V5zwYR+NgJ4yDOPphweOCl/PpkWWvuhryq4DPzrWkQ15ATTW9DXSB0t
ZUCuKrMVAE77HSbd/OkiL17eZj/Ow/wEU4TEG4/zNAbOIgnIUf/qVLdXBKl8RgKb
yKPJlA/wJa2zP9HA+vuHH2BD/1WWC6xeoIRktwkyyWY5JKaUtyh8+8T8NSIrPNtm
3iyelT6mJmGqw0t4mHl09g/rLAxXyixH+oXCEOpJ9BZCCfBOi4ISVCgwSQrFAxLN
2AGjN569GWWpefhk3e19PPpQ7RvmojfiRP7APspYRYrEMaSXtLYdBSFgGswh4XJQ
PvCJYi/aQCrSUl3UwxhsDKh5ihw1OIoLBDWYL48fPccxxnJIb22jrIJ42R4ESD1L
kUmQTLzXJmsnu4NsVTm1fJRujGH0jYz5nbDJuuDBwO06AxRHf5vH3wOv/nY2W6OT
MLBdt2+dAWLEEfBg9yvlqldSHcHZu5XHQL69TICsb/kAL3bhQor5Sc8BP3kjzBSi
zbKnJJFuCWK+D9ZMxDhTmE12rC+SnBAZhlwH5h1tpkfIikEQahJlt1BYU5KdzVvp
iiDL247jPiIVMvlKrp1chnaSk4WkBfEeBMP5NX7iLIJbTNEXvUsg4JisBc4DaWWp
F5Z4DIDBhwweT5KIo73Hxso/Sm8Gibyebd9hJGrvfrDnC0nRXa8OlLM4vhAuVJVc
NYo74heoVaCfucii+PdzyL5eSTY55RebzGG1zD5w6IPKhNu/WtqRDQli4xyTx3F6
9hZ3/A0FWaoFKLiHTn8/1jopxFiqYB0nu7t8uLv/B/PpGtyNGpErhFNvqz2kAhZK
1H+3TxAT1p/CSKAn+6x2+H8JNIi+iun4EjPm6Wh9rn4iPxaNneIYwDRRbRp6JjFt
+QPfDA4cbJPySRBhL77VR2VJ1W1LvbmT4y+lB1L7CORFyWtnnRVNpJsReBh5tE8o
GMvJM/lxzt3l5faR71MprleEqzwCZEewXx966f+ZnPoraXzJ6qEGe3bMw/W9Y7N6
frc72ufWy1bamGGsPtVdJTGP67K3QX0+pQuGyV1jER+sJKFBpmv93YFTZJIM7uev
VmfmmxaUspTh2aFUfUCN6EJDLQJqlll8xAKSoSJqijiDVYw0tX8iWrO9eQMBGFaE
DxR5eo4BENIoV1Vkoo6Takqhof1T8DoEhz4v5w6CyBY81+OqD26JrlL0n6fduBbG
6EQTi6G4SIml8zXDT0Bp7UQzKfJFSISQROKNGeJOaWoQWOSC1bfJbYGu8+JHjcVl
UjMAy99Ggc4ZlyCAsQ4UzwGY7rLtR03fdsqiZdgZwLlk5JFu/Fe7Iesrfb4X5k8D
0LTs7Vqx8jJNu5oLaVJI56mmlJEV4xI5oYpe5Etkksgp9yAMo4GPXJi4V1TLReB2
hkZMN2KxJHlX4htoZolJv3k8B4FHkZDQeSLBtRn7s3XIZJXLxs5yy/T2e1LlOiAN
IG9JUYHShSyqMMU7AsrkXY6OAhDhvFOrQiONhTokaQN4QvuoY2TQRUmfh/1kH9Jk
QC0uD2F2fMfkJcmNqt1AuFrfF0j4SCCNQemGY9NbM0snxgCcpp6CbkOMfBtm6Fgh
LM70k6Ovy6eFeIqMzMYsHcQ/HMzhOjt5zBPhvwOCQ83m5J/xgq3l4PjvTnH9SzZ0
ckauxZHG63CAolcEwXnC5rpL6EnfTkcG8EYQp5Nor4wRPsQ9oe+lW4EaiHRdB6J4
Qq2CGH2T2Wu2iB4VDAgyhr0F+c3U+dXFrUSC6/j3RBgNdkzp0hp2X2h9YvaJPmbE
lb6fRDb5tzmbmjkKIGQrr3HErgDy80USG2w/GdW4xgqbNXqh+QxZn55nqpOcU4iV
iIUbC1ihdZThMhnNzJNO+kph81tIoFZ78BlMVFu5EOvwLhOzigpbWcb4dEH74zEG
ekDda3XarU7YetddbjhZxE9qMTddFlJZ7qk3Oy2K6ZoB5uY7OaFIVgQiLXIsueGu
X2ScI4LSfhAwpWxCKBZFKuONF5TEy9qV/EWR+eQkuCz3nTqXRC94ZuckN6zZb6Pi
nb6yN00cgmiwROimdGw4/OVCxfVk1gIa0nWovrt0D5I3pBkn/dnsTsC/27X0HymF
IdEfIhNO3bmSC9nJgL3mcMmDyEJTsbmrCkhb0eRQ9FReWjMplzHCBYEoVp5hYX5q
to6QMroW3yFXEs83e58G3Kfu5VKSxkCCzefhGJ++HMg12coPFBEVY8FBnKR1eawO
hvzgxqs+8ftQ4Djb1ccpQSSayE37r7QqLAuce7e7aNZmQNQY/WNC1AO1S3RQM/l+
qRozOeLo+re/XBSpq0GGPv5GG4g3VEmRPk/BbWVsjMXKWA19vxzPFcojxdRg9UVT
2ObPe5taB5N7y7nTpAvHG5S2Xk8puDNQHTZfprUHCEazTQEwAMuQc6CutLCgoNKn
mxZgSNTzhEqRavGDfARA9WKafiGEOsTLoFiQa/zPCWMRdrns+Vvf99JzNE7D4dKU
kThr8G7Gu6zEfZaGyryVOJeiya+Pg9eWQqNDmV3j82aDVWBfEhXhWCTJSBVF+HsL
ETgdrFBZF16m2B49wy8XCrCjrr0l1IkV50RpRugK3mRXGVwf9JPj1/QNdystVfmR
fm1LYbrzZDHeE298Ok41wZmJ8bprCroo1bBpsH0GGlwomsNZ9ATGXUsJVqJw84nj
GMWqstWM5UpYW+9Ye1/DEwxkI1ybypQ4RFVTyg6yCn6a9UVcZ4jDff3OfbgwThOO
rwItnRz/1VIVP53ZQlkcdJYT1m2eB6lWT4KY1qZ94rtc/ZZIaMy3gNDK7Cv6Llmg
byU6ybLgGb9aftd90wqbwgJUf99Fy6USLomCsu9T+ZP070qhLo8b4gJnIu5vAdIo
/jKINpl2f9DGQMYh3B1Whx9eycetO3CLVYco05jKwRjF+PN8fByUYU9Nns1gTKGv
utvrTg6NN6MvKZPeQmjuNtlgXvzwATT+vzXkwkbLz22OIXVW3P3X3Vgz3WKvBYp1
DSPEY+g2uiPLr2OggWtcuLoL8BTVN4c2TYDC+NYKayaNXsbcRV2QleSupg7oTUr+
i15FUxvJozjUvmVIVzGq0YEk27v6e45uTKcrnVCAIw8t7xcTBIbcvrpY0iou5mFd
AdBF2gepNBhz9XneriKhILwaOQuymiIImo+w52xt+JmQnCgPwjQroQkP+zOvA7E3
bmnKIdZY20UKyP4K2nJr31feglZLxEBFpjudj5gdcjU1Rk+RDVD0FV27XK5DDiqw
hfgau0ZwyD9Euy7sR0CpJBT6N/UefyiiBvDIMm4/0h8TE6fmMOf6s7EfWJGjsILN
Yh0LeBor0rXosW5pbCV/4rr7f7ZYvCV19hrg4PvJ/iucB6WJRBS/Qn1xfGyclWva
AHdODUedk20VRn2qvwA7iZJLBPzVsRSw8Gk0TvHp/Rmzjv2OCfc1OA7syxUxOLZd
I2fSuZjR9KfaxJCFys1IGFTdILDNS9lKct/PFiK32muYN1UYCTmJS2ukBH9FQKLM
1AXnEkjIOTStMtcw+mycQAG31OVEHNusnDDGhGkAivU4Y1pLKhZXr0Qu9g2/2A/Z
jQgdNt5Lp3rIwWi5p9M/GRAxDxk/U1jVIUqpKACtk4qfudstcP+CjPCGHTIw2D0r
KrYZoyB1ITNAqyVSCKME2qGyIUs334AeS90UqIdjx0SqfcuHpWcXiRfSjH1drfPb
/uJLiusAWJXAgd0AvNCvJeWov67a35zfOj1F5hbhKA8VUwDRAkE+s7IxCH4Hbgm1
latnELT3eqy12/IFkZrvBBDBj7C6RSBqt5r7yuqSV/5c4C/Af5YW9Vqff7dHC8BH
S89dD6G9UOCCTlO9faThoZknlRtXv7CZd5pAuiCKI3p0nafgSrLlY2udwbwOVgVt
GuH5i+KeAercktUf+2oO1x76j8MSg//B1ik4TJymhP9f+8W8x1ukgwSW46fbxgLd
yQqH9KylLAVRUOOVpP11PvTq7Q6Bw2BRWzpCBcGM0I1eB53TP/+Kbm9CKaUdEFg9
MZ9h2zskBDyX3wvqueRh6o/QWdOdJ93BQ96xEaYOV8NWgUFVMID9KXIRIfbxU0Va
B1oIBp3JcSP9nhc7DATgvMlj4MReFLUBk8F82dRtpyiLwvoQJJeCrDwi8kWwqjFy
q0wDpU5noAA9T62pkKzAo8m6BVj4Wc9bjhrosghB13o9+C3wi1dk+lPshoumIA4A
IqRrkIjTFbx7ub/j5JwoUHwIvvmtzzslh1RCqOdKE5rb8Q74NJHccwi9fYI7Cvgh
5FyK+xk/+RBCTscGmJne2GhIRr/zgkPlpfulfw7dRhebvrFSSfa5iTYyBsy+Vav6
tdPHSgmfO2QIQfaLj5ashM9XSpfXCQoFwcaAF2W/1GiT/iLfIuwL9p/p7AkIX8Km
RFairZ4udSaJRMp/vZ6BB0MbCF7kuU8i44CdQzMit9zsE9Hqd8SZgCabbFjYTucL
UIfHv4NUCHgfEnBrk9QxhC1iktNKttoUv4nUD9/aizwypSSeF8lif/QkEUfFusiL
MKf1YzDwdC/Je9rNjABJuvbbVySpxy0HNmR6c+w2iBke+qm4U/ephm6dNK3wCu+l
kfLa7Ika5k9COf2tOtrkR4UMIYrQq9s/k+LVdwmMTP4pUPJXvGjwlbgUgPXHEqKQ
SgfRsK4XVGD3y8rO2pw2yxomo1dt07Zd7AdZbzk1zugCrrTWZw5zhZ4Y11CqKUUm
5GE9aKBYxYjuyh7w4ZaM86myspM8pA+sq1JdbDgQCTcKyVpF4Vdm3TUNOMjA+PXM
IQit2KjEZi1habHkxW3YXZSgXfOrDGMVdwQBtIKHcEMd8r5X5Fgg0KeGcbRfIEoZ
yTzRIQ657OWETasgMdAb2XbFPo6o3bGEMAtiqJOpFL9YRjmRbuvlDYuLS9j/D7U2
1TM7I5Bs2k/7lvHjQb8a9qXRIPXFVe2emdcnqlVRj6GTkoHJQ9SInsiZmg6hVkBL
oeu+QD2I37FLzkOj3mh3+HaGQy0Cw1nZXOMhZiyn1xuGh3zGG9CT+SYfKAl39UQ9
uHmDXOExt3pPF3cQIvCQETAq0BqI/HYoj0HxzsD3qhmBB+jaJKWNGK8l46HumTwp
KCe8u3DnwUgn2PBnlPQ/UkpQu5r7p3HjDCLaPDW2Vijz225ukYUlb8yCs8OHkA58
Wgk5gC8cCQ+pFybpVNv8oDO7E516nCe7dUmhhqAkJjBlHMrBS0zapw/8mpysfsa+
C3fPEvSriYZNRa51ddxGFFlxvkmxjryRl8PdJTaTQv8R8/sCk0IXBG+h3J3iiO9A
P2tG95+XNNnzglCjJTAXXxWy4GWLss7p9hv5qpzeCkwXtB0HTM/+8eCB0xYKGEH/
QSbNBZY9c4BipkTzrV8PmGVPKuRqigmZ02Ha7JBC7vcDgrUoOjrSs9OPXXzDKvxR
XmNCphnQx2o4T9fd2ICM/PVyNnxxwPqwVUKFvKBnSpo6IdBaJiXUCBpZpWQi4tq0
MkB3pQbVEwnExelmiqIevZ55t84EkAOOpChFDZfz40GfPhuY0N+qTZ6D5oYHhxzk
Xf0FcJZG5Js3DanshwRy/vV8oIl0YmUkj8pab4GveoE5hU8+abl7RL9E+3wUM8pS
ZP3awzQflXt81hdnIdb3EH9uNbR8wGOLQz8UpWQiTjsyclK649B1c6tdV6eEgo4d
cetrhnv3JlDyux1rxgPYjEhK3wZj9kcpvtCLdXBDDH4ZIh3vnd8xyzqtg0maU6wU
1PB5xXnmiVkRH8o5Zk1SAlHGANu7ugRqUJHIAdC6I4I5ccRQF+sfuHxhR6ay0nkp
2Et5grU6+A+amd5l/ylWZLvvp4RxNi2bVc4IAogHL5E60OOjRYejamUK2bs00qky
WgBoCKyoyrp7cmGT0UqMoC9N0R+yerFP1UHAD+Rd8S1IVZGArAXAbRpk6aFKyzg/
Fh3zS6nky9cNFkLzi2oGn5UiET1jEdOqu6WIj1eWL59kmZi5QrznD3KRujgNZCNq
ymHeFswt5aoTlIFos0YfyDX4o37VzKxWvih8KGuxCFhiw4hdAmN+ToUmdpitDawj
Oadcuri8nFrvjYgQzbWKdwlDqqORWij5hJ1U9gqDjpMjmcyJf8mqzvyeB5d5EgUg
KhWflgNcHbUsSMU6G68rUeKqzMepYQoRmEzXR23fvqy7Sf1ywAdUbKEQH8KLdPew
Lri3B7PPHl6F+aV1KzcUXK/uONEy2E4SbZ2BnSOUjVUlDbNsAQu10lcym0VlOmz8
N/PYPbmPj/ECJhPuRZpTuJ9SgYnCr5tupg0xRAKdWn1SyFjirt21hx5C/AEWP1V5
SPQzbL1SKIxdRfMWcOzdJGWP1B5zlwvqD9Bqrlku6o+CuGuCL6T7GK3RBJSpzg0x
vcjEQQBXqeWXs+OYxYnMefpkxc27rvXNorlKxmwonjded+6ZvrC0LyrlrHR73mWi
cOT0epvA4Lv73u0dLlJHpfIOQQ7YT7PuwWx1JwoiQ0Z4+0qmRsY1mTMWuW5HYTLP
xrOTvqORGdnw47f57I6TV03Xa1KIoKerXy4Ynsz8K807yy67EXLVd5ssPxdppiBx
j7xsMSq8RZfqPe9qLbrXxnooQPQSvcOxNyC8Mf/hiXxRpuQdvg6q2jzc2sjVpcEK
6qetyYPMzCXIPYIPXck8GjWzbexXI1AegC4PrNvI5YxeAUoN8j8Vgd66lTi+wO0V
6MR5rdvL7170G+wWtNz0SwBZpxxBlI/G4+kXQP8k68xM7to1TRIO7eJrMGfPGvJ2
vh4djdWqx5rsiO0cFTK24HssaTb2r005dQCIZ3TIIPUWq9ADRzO/PDwd7mklzK3f
ovmfQ0UoHuNL2I4wwTCdZVeAA0JMWEA+aQQANiF2zRa+QqouqVsroBQbo5XGR1cA
FYy1yLQvY+6cbiHUFUoRerLY9hJH1J1ADXsyA7szMuEoPgYtNmQ0QPW2JHxBk/zB
bNS4cPeqfvG+3S45bkj7HiIEyFJVdRwLzS4pXH7SWZ2nldEWIWEH1KIQjl+A4JcJ
6cK6BGHFvmVm35sgY79x//2SWC0KF6Kdr8x+OpQpGcIg2GAcwaR7dHOOWcNsOdze
Ks1P+NnkQxOL8/jCUTnxogMZNRrteRvr7KiC1e+v7vMHhI8QK4FMN5OYyIuG+kfI
x05xAJKLyCBDKHBgeEfCRKmfGrFI++uAv9XAYgnlA+PhHHwz5+JKa+maVBotyYNt
Z+8xZWfZ+d32LqRWHdSSqhdq7VVLdwl5hn/CTL8y68ro3rGUtT2J0qq25lB0Pzhr
Dj15y3gGJVkoYIUTC2aSkbPujep/Dg944I2fhqgEFvrO7/kW6flN6PuBbhpAQA93
iL07PJZ/jDnwozTG6ycVw/NNaXMkFhIoJdDcfbthrj2ls2fsVdd2924wTUBr76wp
ECp8hccM/I8g3N3xVgQ8FwmFdKoAeAPRrnOegZeLNdZAgBFWHSbeWiKFYC+XqjgC
eKReG7lgLyp2O9ndWRB6N1Qg8362nvlxeipBFKrVqeJWLoVsEZuIJsS1XyIdeU2M
Ue7c8Y8rVTMXPDz4TJAO+KFwPLOKY6g2+Tn5879lAF5Q8v5oDIKv8G7Lo2XvizH4
badJ6C7vefYTLfzjcpU/GuzaszurVXDNlZnY9IkWp8uQdebdBUguwH47l+OwwOlg
TPReOdgdyIUE5rtIWj22t9RmNdn52VxX6sfiJPIuFK0HIDAjcJzIAyu2pSZLKopU
4zItj342Tca1dgRm6RokNbI4sWVtY38JOPsbKirAF7YAGLhIiBC+BIBPWMLkd1wo
UJf9J6nY0C4Cifq3bReawYavRiQYKSQtpKyFxB9FkXRXwEyOsClHMw8oc6ORT3P+
eAnhUScthrUC1ThIi5FLiA7BXmxczm9eCtOrW9U9nvLbdn+z4dowMY8ibHssmixY
qg++IOmistlADWTdvhxG3gbZLXerqoYyTfxaLbEZGqviNwJmNFG+Ge2HJtOvuyU/
Skb30q7b0hH8jCws9wpvkGGk5oCBrMEXvO8tErP95A5koKpeF5lgA730lahPGJ6n
LyIEzLg+kpKSnbpQMABfvavFDVL5qqy0CQHDZFEx/tgwdxKK/DF5qaX81XM4AhYV
t9AiOGJss9UdREVQO4ukKCoJWrsdnHIUMWttbZCneFpzO5Pwxs4xogjgnoI8RyGr
+ssqC7S6JiNtl4cE0xj8TU0qaMbZZ9uELzGD9YHazL+TSzowtKq54qrpkpJ5tQri
xI7NHeYrpp8v8x/rBLD3umFkwBmW/LLbRvBy3rJaYKe0KHtk3kCWw/b/6eeEcE/H
Jg3CxqIrs4LnHd3PZgd3K7WKCbPuoxHykH5AfTo/xCyLNJdiGHdZce7om/riWg8U
iMbStgR+0Iry34htIODoS+gKlirflI4qVpndzx+hBGIa5CU7wmnGT2hwhsKX7cLa
Nn3GMkm0aNb1BQSA2+7PCm2HbF39rqLp5Rn04g8ZG7JRMu+MJdCc1DNduYQI+KwN
6AeeDR6xIt3p7MasB3cg/G1P9gdskjcPq33jezPiLdlrlQUrMH80tRwjmLbahadY
wvdW4swhqQ9Pm5SLJbeu3Gal6VYMrXrpJyoCB89ADQUmHr6SgNPD3ZIaAo/vWYBN
8tsaW8XJZcPuHPn8gH+YQA1KnmQnw9075hRZolxp1RTOQwExm0cFIm6ujmXBv0cF
rCjeNIP7NT2QRylgdmg7hv/Sf9y1uNgL35veMeLGEccIEdF59kwENODJ1F+X5dqi
Of+Wk2VkHNCAwP/0HmM//AaDsbpQR6AmsjBuq0FxeVtM1G5aIYJp2lNZnbPmcOjM
mxZdQWPFDr2LAZnfAEsulCRptCKGy07H6Dl2o8HSfGAXc0eckVU6XLUTzJ0pKvDl
XfE02l82oUo48zplYMBHE07UOFzN3WGbG3MNtLgXKoXgP3tCEz3KaJT8ohvtGN5u
Mf+f73iwR1IX7m/0WXaj47GSRAqShFzIqXO9L8/lbOr1aXfwO9xiHL4zxFBGb3hI
osf0lXhm872x5KPV/hfo4wUu2m+q8eH+BOfcn1vc2a7JQ45mwsf0AXiVsIxNWXQF
vKyh373L6sEgjwhNTd++KcdQyxpBvAwttYXSGExluOc5mGoezK5cg9TUkX9+hRai
XwXY6yrUEv0ZW3VPNvynJB/kLsNt0OfUjaQHT6cqUc3H8nofF4HQiumPwcfkruG2
temVxCgIsVuiwE4m2a7jeD99rsbET+10hIa44+Au1u6J5klT5M5nO+62PF1/+s+0
oOOEEtdYemu3SXDiUge1pZ+HzIkP7/Xj8qgw8ZBpGA2eEvDQG+NZkZRFNaOAgyV7
Un3Ax9KW8dUfp2FXW6e1V87lFYAy3GBuuYVMzXraa38vTO7RzU5CSenDXU/62zIl
MvVdoqVA/YzFdoe+0YpOADepCBAgD81vsLP4yZa03/rXc1VQKa9yQtPYXg3evAnr
kL6CWWPujPK5Z9e1b1YLX4LHpns8RxCGU4aqHFpKJGBlhv3CqxV90HiA3GcbEPme
5SKJN4DefARDY+JkTCKbl35vie2XEIZgeORT0RG017lgfFHvXHphokRwVLbiZ4te
p9KXkRsyeqmNG/fBWPy/g/3OwDOSJNP02p7xEQ6Zs4YRj59aJ4Aio3F7S5SZ8pEY
JuvsTIysaBoOtjxm8m82S2qIxnaMjGMcqTjxLfUsmCGjOzdTenYaOJrsrTtkLmtW
5lFf1lrARv++MKqEmIhV9jj6hAnQsp6hp68Mpv7wWNp2nrESYOZj9Bc+Dw/l0C6R
+fFvlFIvpwekPuuudUDwMV7lFAxok+29RFsG1usu5k5c+/9pYmXQvwLU/VcCMP6L
JJJU041djRkb2Y2q0yjZIgyq64RpcorqAXyHUtE7KWjlqTrh37Gz3pnIwG6x+wNs
FUP9f6jgMypcLGawJj9mARpLppToOZG3RbHv/0V/gbrYs9jwfSRmlQF0lpvvo4Ui
2q7g9vqoYXcmYcnxuED5H7Pm5FMuw7O8leBBeSoxlu5Ls19Tc1Xzdfr+SFw7WSSv
0oP9wFZXbVvF4AfUJ28xTugh9+xbt9gU2CmMygrqQMaRnpNv+uBRDYOdx3rDa+Ft
yiVbLS4p//t1TS4zQAFqFm8RAsQ2QdxBpJ2UPb6sz5kB9w8RK8wJkEsCHokHVcgJ
QhlKT4i3C5KRh0wuTToV9kNI3bL+C+1Q2OT5W4WmDuLUz8psig5wU9PKQ5BzaWFH
CGMamjNFPOJiQw/GpIhLpB5dQp2K0dbABg45dE8KjuHzLuN/qu4lfZ0je4fNV5np
Aue4FScgztre7eJ9+1N83wXdDikX/YBOncHLgqALyJ3GqXCWHg7tVyPo0fmduo+5
pm1wo6qHgmKUHKk+zKKIefo1bjmGN8gmBjqax6k6ZM0bQ59NIpGN/59t0M0oT6Lj
FZfL8IAA5R84267/P5m6E5NQ1leHz3NIfXkmwNJaQYeXlFBgmHVjEAZ2M2urSdC9
VFp7Lv7U6z4UF4OJ1A2ghj8uHzx0uck/XPWZjfSQXP1D84KMRPJFM/Ctbe2hDYZq
me7m/pEkjgmK0/ndDmdLjyfWK3auSLirhbUSTb0ge2gb9+CwD1yTjNNqrrVtPTrM
vH3byAuwby3futNgYhZgcdf580X6r8OFFWJg8LWdAxCxVJSQQSm4XBh4jA4sOgdN
oQJpbxxNmnyEzIzfGFys+/67py19Hn7CW72ig1Vd441seLTjZVE9nVFVpSd7I9iM
Vd+qWkNK/rvFtaYR9tnIGu8yqgMaQ1K23V/7UHNXyfnivy2tVg76bafEVuCBbki5
2qpY++jCMc1O7JYyaUEmM2oBja6kPoJvJPmy0zAMSfPtU+RSJTJn/EA4MPQJFuV+
F/WobuZvLIZV5NQC+/jEWzyknmWfpq5/hu51ER+nHOlJiNXOGK233uVUonJvfQEG
HpBhjUyaUYpI4yuKuYfH9RwvQv1ZQr1ysdpUn5g97F03rR5cuC1D164Vjna6rgN3
4YyO62jqnxP81sBhetK4SrupoVV2a7U3lmAUiIn4FIr4noTEhV8qgtbKmLQjBVNm
uZu8IytOBLuXTQMv80TRzadVwG+YwER2gX4BKl8AoBthc7CameUIWYXXfw/Yl4dp
u6DV9LRo6DdRg6LOsnkImKpumhbYw4bigqHVVKrsM8+pL+Kke+2Jw8Cqe3iBTwC5
XZq4Bob7TxYxOMis8nyfuCFJllzZqQUyIrhoiqHsoFXAR6CCY97nw0Ulbi3KdaZx
o72EOAOO6VDMm0PkMlTiCAI9E7MnMIIu4imV1ns8POpjHzs/K+6i83aElnaktLam
9ZnStROmVAXvSz26KXhog2m8rv7WxVtoIftnnvGWY0elsweE8A9WHCI+A4mPdeBp
9Dog51R4JhVOYA4NIuyBAQF+TmD6nX54BGkDzkBAlWJoa6+qVkdSoQ7Z9s5c/m6V
XUB5tVrTcU7l51renXnq+FAkwlxXGmUZ7JfTuSnm8/2SM+yiWeIKWX3ZrMblGPwm
hO4R/48HQHOeMecPTbY5/3D+TqNzI+L3H+/S00RsbWG4aS/fUfoEpkxgu4eHc+YR
PGiEr51m/xtHOII3VxUocc+6HKOhWZq0WRqGggj6sr5p9XYqade8i8Q9VteR5xPK
1mwZVSMdEbZohLiPH0X9IsQjHvV5dMFd9FcVSa31wsDy1jU1cZa2aYHt6KOgSXkl
g3f0a0JXwGDkM/BOf0jy/+FCSevA2n/sIllockGo5g8zxRzfjUsNUJSDxTIiMWM+
ESyhbvH43QTCr14134OEizNBCM0ZEv2f32UFUocZa8oQOfdUdvD8UAD43j3x+H/s
NLiAWBFhdEhAWTu4gZMYmkZseTlBNmbq1NeC1KQSlyksvGt91ppx2FWcGlcxGIUp
kshamk8SRnQDOpVcx7tfkNfS7fdBkXiHJnKGkBhWhGONDZV1qHSaN0Z6+eRMwC2O
2ZUNYSG10toH8T/742noxUPsljKdhQHTVH/eai/31mlmZvQ4dWWjsraK2nugg9ik
0nEhEzgQuiTBM8WAvIWLYxPUYTh/eDfskrrpZ00pqsEIQ2RqiIdWBLzmEW4yQF60
IG92CMVVWTrDtor3DAdJ/Ke2zSsQPmSjy52z1qnt7dQ8ByOuzgjauiZUlMm8lADX
SzDU+DbN4uVPm2Jbm1vc7wBe2os/NP16PAOgk6Jdn0Cez6O6NgSn6ZCzlP96c8p0
kLHKjfDiPUmxrY8svdQ4wcqmo8SdJiXbKfmwVFy7HJ+2MbJSsppuW4lI5m2JZhmW
+J+LE82AQ78t9t0aRerXU6kseSGWf7+PwXEsLfy5lKv/BtvdJkOleoboojWfYdnR
197V2EyB88StUTHFTnLjIHxB5q1OrmEClmM+rs+C6LPHMaNvUFqPi8vwGzARSFkx
fu6AITbthvnS9pFE5TSoPlv2v+S4wh7pdVyC8MLv+4Qs9sRZtDNb7WKzqw5TN8Mk
xkhYnBswtaMa9k++DumgHOoE96fgtB13Yy+kwcgxQ3FPHkyzr+/ndvYpMtZuhnV2
RIIvz2sprmFUvbdRC0/d401vcZY/38jXd9TtCC4Kv42gcAfj99/S1527hv5qlegA
rA9NQu6CkWW4+5i3kiIMsR0J/OGkw2NVzsrnLXQC1msZKa7DOiaWzLgMMDje568E
c9QA+iniDEBQgtpj4TyIM3LbdqJwXjvt2XTb5CpqKpE+qZlmGpSi8G/nepbt1hSj
oSRmXINDzkbyBFyy1Zs9Ft0RY80kIo8m1j14AXi45K1K7t1Ec6gmMEUMw3MnYZ9M
cAVD5Q6muomsThUzLijJ1cPIlfzV6KCwLXtOi4WwYh3z/+1+sFekdLM8sV3tclk2
fjt3eKt9Pu9wpxp64d5kWr4J8UrQTnScCWdDgMv1LgH8tDbXme8D28DLea5xaDSH
C1o+OaMAp+TThw56xDm0AjP0yrueQ2UpS7TKd34ORgmRwlgWmJegvxUsy4V9g6iS
x0FsVYgSgkmJ0/Jy9rRYbs40rhMwIvHrxl8J7cmqeXhyCVoGEMZqNY1cvrWKMLnS
yfjO8eB4XcNf6GiljGJCFOBSnka7VRlLXml3V/QUV7SDcd4duwlRfVvpFM4pBjdh
TlsAR7jM11PCvxVBWZ1dJnL1RIKkwjfyKxWgeqnRmBzHGJmUAqSfYKSs3c+S9MMm
1pXd3CSQrJ16Bd/XK9AiPzmTushiHt5nk5zyR6HwainUWF++MG76sQLq2/bAwOIG
2AlZzOXNzJWP652sB0Ddt2m2i153iW6F/YPmMhFNBPn7W1GzpA6iyLZ8WIfl3aAK
z+6vwpvmxZn+Pgwl0AdTpeGIOOxK7kDges6qfyQ2ewvWMp4tloiDoknimJTTsN3T
neDNP4iIzoqVdAAjv9EAOS9tfczK8v1KlMSkHhFYp7SRK0VmqpOMMhTgAD/qdAz5
CxXfQ+l/vKC4hrV/GEGd55B8e5LC4TbwFWDeguxQ47pdHhtcoYBsDT2SnQnRcGtW
szStHkXlIq4iFA1fOPU1lNhj2idg8B+pJeLNHLl0p5mB/DTEJVeE/w53ZTrPQvCP
wy63RvbbBHDsmclE5H1ssl6fBbt32OlEWjlXINKfN/CJADU8MgU2MaFjhxmSp+6v
4FsFwv+IK7Jus1XrZu0SSRJPRt8O8YIpY0uIgr9+oBSSoe9aIvJslTThKqRt4R/H
/1PN4I4ZLQOzxavCvpQtwuVOAHoCKTzEmm2qL01H5VBs6JrZU5qL9bGSV8QovjIA
V1csqJ8pFxCOW4s+WTDNT4Y5pST+lWxUQcY/4uKyheGm22jd68t7RJddQLaOmxet
6W6ii8Oq8ff7CYNsHIxHuqYy7eXjYh3/eaSG7kQ5xRDQdI6yipNvHv4XvOsaC8cP
d+AAZUkg/n1o4EUCIZnynqMM/xMXSuHM4lchRgKZ3msiamv0f5ksL0HFBxO8+d99
PXqjfYBcb1FudJofdjz4+BbrBS4UNQ2Xc8EIVywvOIAKNf07NeRu1D/gOBatHtnF
D+OjVlvLJk9BqBa4pZZPRs1brrUiFHF900EmfsrV+MGAQbjCbfQcY3Tw3uBbyRnz
J0/Vw7CKuY8ibSWfhJD+nzOaHjloys7Jmw035sYCjUm3Yk0WY/MNyakPQbNynJiV
MmQqReBCi/s/kgxKcCCn0Al14h4u3lejqBBRcvmBKzmN7s6A34xGjar+1D01hka8
CYaGy1Rgh9PBteZlrfeyh93WtZ0FygUNE3d75vYN/luwumJrxZkTEaSBzwbsoTvT
KLhoCVjTiyNV9itcnZ0DKt5bonEBrJ+jKPlfq3TLZ5UGdTmSy3miGgTlt+MTT+KT
+nZ+txDubFgXR71Q+aAYFr97sRz/hoLc8L1El/f2rwcgRlaDycAug3VHGVwgMI2H
hH9Vwj7wZ4onTv2g2CWCxV7Rxa41+uyKIrmRcMunAvNxJqT6nYbPmWjtHq6bAxd4
easiLG+vnDfMxAjg7Xf9FYEuHVLN3ZoMUUYmZ3H1xGinpvv4JDyWnyps3s86bcVT
H8oFFZThEPCHp/08MX9MuwwS0qYEWN1f0zIYW5HCUeKMqyYs7Jz3jauCRRPDU1oN
hK3nzj9pTzoJWvqynniIOm6cuzHb1Puch3QLkbAQ1BefxIXgNFyPFCApMDsMJvt5
yy+0kJ4F7cRmFVQI0LsAwvBIgummtPHGDCCvywx/R6IBZMM3+trjMNQYaWRaHLos
LigAaS3NlYDunWAcLXdMJWirvdVtC4f+ZyC1WnLcHhepa4S8NWY6G4N9mXGkzWkp
aMZ2KsR75n7028VzGNxsRBkvbhxBW2doV8sbpd/w64vGix8tj80Pix8g/IJ6YGyW
FbD7iedoigm0tEj5nsPiUCtMh4ttPlVGei1qpXrqWvB2tPDIFkiIWcINPUuP3POg
nYPolhznPmNXCTt9NTZGpp8+V3pO5RSg7B6LCbJ1skWNY0m1j6CYdUHWRO7xA54t
5B9WaN25rBbkU4QIfq23vs+Yg9nHDeYhVm6zOtXKE9efiEtm3wV4Xcu4VFYLTgtG
wLJpVUblDguUackEh8Ncy2XaLDLjTeXeFda329lKFi8oPASI2alO5cZSp88FSB/c
sEKa2sXDw1OE5eJw8oY6kfSEqcC0W/Ez1Xfft55twRvn3WMMm9Oa5OKBlfULRCUd
YN1jxni9KNx0TK1TiLd+QZyQB+CBcPkuoMYoZWRs+LG5Ylp611yxrad0tU+NBwtk
ALPpLRu1YgRBp2uidm3GXuJGm00vD6kXgDleVHcMMcBXyETZbcj4e9slEohRMTPX
oLu5KV3mWBDL7/e47m5UBYEIevvEoeMWCxXNLhM68Iu6tJ1eG6uTLUeDaUpwRUTf
Ad+2BXR/nAfPIQsIiGusoUj64cwdrxaATgT0TxeJEIcXHktxzgY7WiWnMGg3LxAc
vk0RacIj31xvAtZ0GpgFfeSRvt3mKsap7AQXesrDreDiP7C9gzM+ZSp5UOFqW/aq
uoI2QnvCRt2sneu6l0SDHawrrEDcYMiYG8aC6N+Tqm98c9gzlb1e1rGGJiqBTgfv
MjY2w1ObZVuvqxJvqIbUWz3N0KrgwAF5D6wghQyWmNZP/oX9/Uqfqquxb14SmAn0
AE5BT/n7yT2lBhi0JalnDssk0IwpOaeTU75dRIKcgmczz2GKDbTpnuBTqbzG3tQe
Db+2A378QCITFm3xoCVvKk1N8vWVbYVWRGxEkURDBaD7aSfyi8LvOL0SMFWAzW+k
E5rehgPH6Gb/x0cjZ6YBqUGdQMgEQv64CDL6LemBonaMvpFP9732C/OuVhAiQwii
VN1TT+KZYcu37vV/Os8XyypiEPPmhp+2wITkvq+7vYN7WKlicHHg8Q5dLI4Fn8r9
zJX2L4yg92VnQydDNqnJJP5TIezleDTb5AnNimOP576EgvNHzsbQZDQRgW2Z/IVS
Ofpz93qh43DUiNhVEHQETUZDU4uUBY9fg6KZ9axbJEaXYgqpfgmMA0mOzPrSzNR+
6Umn1jxV6tns6W22l4LPcKqJ/eEkw9Lb3V7tkLMJ3dG9aCBtAvCYb0PJoBwwTLt+
+22lJbPotB71CEroTueguZouIoRYglvjejyDGYUkZYRWynQVLCuonDLmMNPCLm79
phLHXB7yFTJnm42hSlZTf3UcnLLjHapIn6q1bDjcPctgPSptSPBSMh+4DVgWunWH
j+0SDTnH63X+yYhvwkr5D/5w+RzVOBcmULsr6jFA/8lDvQonqiWcBlh4+TSBYfU8
QdGyukYOHVxf5q7vsBRSqNJLRDcD0eOchtb0Xz8qFlJgY3Bi4a3sVolohPt0GNLd
fjYwrCnyopMU31TIqSDDb9Ia+9kbSkrD0eRgQfH5xfEsc1WNgR788+fvuPPfxROn
cFwp1l11F+FRZPGfDfEE0aFDIEQYQTgwcyY4jmBe0C95IjKgo1Gw3eVNJxPgd/0R
PPaVSMv++S6TI0s72K/OXSJftnOf8oRTpR2HbYraZJ2CXhhOMZincFi412IaUF1L
bQtNzGLnZ4dWjIUzIm4VvQppuE10+s26UclgMSKsR5gS3vKA0D9W943CwFGX1NR1
iy3A9Xij0Blk3JFo5khUDmzyLnh83XZxaCpkj1wPjg1FEg0sDX/rr16pEr8ZPiI0
tkVnVEGV7Lt40oZzI5T+uZBuwFzRPVgQ3IyMKmRVXcXUtju0fx0DaHCnzht/YmBM
p4mDIs13JXWg04RotX0nOInOKkQ96qPkuYyCQcmFulkSCAvjhJf4Dd7FKarztTB6
nj5sg9HsJAWamK3+wNAuLUqvI7nWsZ71FydLLxi4hCv8sqmwYQh5bCSZzXc2gTWg
2sm8v/rWPyPAvsd6Y6wk0oVIY2z3UqKdCfE0DdAQ4CzpFqk89jbt7kBBLw/I8lvL
UhFSyYM0tb68IAsJ8qM6sM2imM/kkUqGIOudCvYqBEhgf5nQetpE5DnjduWLbYJx
19R7Dkcy9oft1ynP0LKktOidKhJCqn8ZzBBG361+4UDb9//OTNe2EgE9Sv5NJV43
kk34+JGHqviibDaIKZ0yeiuvzEebN0VWhhWiRo2CNv930pYblfnXVFGTmSGqQuhO
1sOmBCi7GoUEo1ekP/77oAPCfdHus8Oicowa5SabXG/71ecOBgwU8ICCCoIuyDam
T2LoP55+aTScI2OMCqLHPDHvxQ1/oLVlL6R1uh/+6+n4EKiQRQSLRNSU+wJ66Gs7
7UsalT2ek9a4Migc6oDnlUDX0CZbWVPli9pnsO4jLOsqxMVqBU5tW0gx/Ab2qxi0
bi+2HG8L8TswMFjOBs8IAX+0mevJoVQS02d2Tf+Sp9G2SVjp7CA7pHlBCttvjJ29
zbNV2egNfM2y8bqrgdiqwn/WGYXO6Ad7sHI0fXgBY/E50E40UHB+rFw6Kk6/RBCd
2yrp1zm21CPHeMktnIiL/piFJmaG9yEH2gu/iKN/HbvmZ7fUA/eYlrqYW1V6po9k
Z91z3wOIifOsULE9D/LJ2BSELILHdQRQC8tGpMpmj0hvkK9YlLbMNAaW8OVaLdO7
/iKe7SGWGk7VkI3hO0GvC8/eChTuwgqHanVjalmHjKwN2qFsyN3nTJBSmTucrP99
TvfDKZMuqpUm0KGasdmZ5N3iK6RaIB09GsQ1O5zcNJOlqMRd0X1XBhuIupT4ZdXJ
lyiK5CWe+DTqGmN3kM1hCktsG92Ioj9ZE0+QttaacmxJ423Y3LWROKGKoxOcvvbW
YNgO20yPuFp4VJML1Z+GUfGlNuRF6bQCei1DUVjpipbWlZtos9lZNicummuVCTbJ
dg1IvHNHR8yaKC49IZufeAezEChtu1Qx2xhE2qCLbWPc+T8SDKXE7L+HL1bO6Dpk
RbtS24XoHeaL+h/kUX53GeDq+5+WZiCCubvA6a7+WT6nzGrUjBN3oq1SevhiWqIa
es2iLa/v1JRZgDSm7Qbr1ZN4+jeHYgsO6saGY+L1Hlsj6/YdPIR5zLy9sZQLpqpD
bZ3lWiGdUiqHJlhkbSbulqOQYRajRS1ZRmgiB3cxbl5RXfZhzUz5D0AQVgzHBv+h
cgkr+1Xnla7xPRd1Ht/OAbjA95wD2XcsNZXcX6OKFjy4IJRj9UmRrVIANH3BORgc
wp8hJQGVdXc9K0ncLmePdjS2BeRgkiDAW/HXJ7Nh1Il4OwbJPSa8eqaeI3G1p8Oe
OiG8sieVKEoKvkUEi810GZXxIh4hzC3bXA8R8sfRlotHYpgJGN2cDMQsbjx+8O2n
DFvi8yTOxJOxLa6A+iewPB31Et4p2L4QLADMH/wTqe6QLhTSuRY761/rb5iQgv3N
egcy1ZePW4wV9qH1UMb/4KEllgNpCfT6V7ES8eIKXNmS4e1TUXDVSmfaqXdsI5MC
rBWhdG+u1P5map/HQqDzBpqYsqeQd3QGEQirfBwHYvbogPVkxD7szHX4AeV+vY9k
TRwBy0R54zxTZTfKdmFFFM+cXGeTdi6GEDFcwTwIqzi1zVbmpvFSkYSqrS8sZd5k
1LBTc5JHEa97eR9uRE5HWtbFj3Ii4z6RzvQObime/8enfj5q38feGkeCNIPfjA7I
oUAVJfMvjioWhstXYI8hl8uhGL3Ls6tUtL9MGUNoG9R6Ha8jEjyo5z4/qsQC6JGC
9fcXNR1p6k4sR+IkFau0Oz4aY9wGoMFSZrurs8UTUofv+Ht8ttlW79xM4Y4hjyhU
4zhCjj10kzgtDcxmq7GGJ4cyuW+dRvKbXXujHNvg2ybNikaVdemnIBUT7zlKOUPi
rj/ujNta1DUqgSKzJwxblFiwCKB3erMXp7sVAoTsKUy6aOeEteb/HqANJzPOGAv4
TJphLu3oYsR+QuPEXytfqJJ01W101VlQ5gTbIszmKZE1uxAICgDfxkASoY9t16g8
+DUnv8EP6Db3OzvWhcrVmaezYSw5SLXLsDXqOvM6UEHnDeiHI9TQDyaRcGwT8xP2
LncYzgFtffDCW+IhaTWVIBNcCm98by8z87hL619FmoxrfLh6v+0TtukVnL2g9Jjo
aQP6MK9zy3AfXQTGT39YDvif9WJPUesp5KaEUxEgJrPdFAEuUqsYXzJ6ZJ9e4oBA
NbXT2fM4f3PNvjbB7hWs6pdbCKS8Mka72nmdnhgMVNl+D/H4WGYwEbby+57hCzaB
MUNTd5XEymUy1TH75OAi5paU6sNXD6sf2t89BVF4ru7RPapPCzPOr0s+H5SOhcO6
uj+4GeTrW23dbMaSBqFWad4b6TYaB8FBQKGJO7xSgQMO8KdvYPV65/HGwz/P4Z4M
ten32C8vMIj05PLiBs9TYCw1+XGwUtXZI+ArR2IS4SmXkZfvgTGlJ5L0tIt/K/St
ax+Y0abvw+KwEjEPj1t2ZGIfQPcAb693Yc9xYkjAeAmyWyXBDmV84KYC3YMVhgV4
SBw7r7OCQzqQKpIXOhhRr4NdOzNnapFrvRdmUAX+oXTZkQgngEvf9hDXUJOxJ6rQ
CU+djvAP/jdPUKKJI2F1/pd+1z2i9Rre1jEmw/BLCamjwnBnMAfz4TdZmDOxEiB3
wsWQBeNvGSRPboFr7oCWEl+31lUKGk/9Ikt7A5N2Z5GNc+Z6hEZUhEA0DR0GubnY
F3GRw2fjn3JMjZXpqghluK9hmWjTKm04lCPBf8xGb0wWlQ5uTOwf9hFv4IaiQrHZ
RnZfclAjICpLjCAnrl2kusEZc7Nvzwiv6PuMHoDf2AmT725Quo0sv51dz1unhcUi
DIK09xS0AjmXUKmayr3+MhO7iUqrSqKj8dODeFRvd9j62k642qEjEVY3kdOJR7wa
x8TrKBnzWKyBYO6hLZzLurycSksHcwpJnPkqg/cFndT7ZAh56Qajr/xBsoWk36PS
Q5+oUtNCzTNm1oSa5GgeYYIAvU4foBForHY0OryVp1qqADKMh/p/nDTsQoSvLtOL
VX61dgmnVFze6Yk3SHYwyi2aVT4oh3hImYCngdizh7p88We+bths+DkCJyKSMIRe
gBr5HlJevEdybQBf+hFLIa1siVJqzb7uPGgmTBpPSCthvtSfAJqqcl252mcTZnFY
T4U52dpz/AmnQqbYPDn6Q995Ihd14xywNfc2m46VFcpYO3ceB2I6S3239RmIk820
YQaf4+4K+OuUzPIz6TQSIEvUXTd5Eo/W51aYW2380FfqdLmmtZjZGosHTZ+ggIRt
QortwW1nNSKsPmyc1wjQ800cxp+bujq6XKF3KY+KJwfyHnUdN6w85JRDJ/jWriKU
5go2L599OoQ8LtzCJeJRZkz2BvtGMaV3L5mywuwBawHsIe9+BXXJI3xzLzkQxkQD
uvqwhjiWg+99122Y7mbyCgyFDyNnNrDaJUVSiyBDo657LH6Zx8GdJo7KvhBek9BZ
bA9ny5YRnRDzaGxDFyso6JSPSd5saaUoACPnnnc8394luUNRzC+50d2EjGXOAW60
zfdYAj2rlobXWVOio8FT5/GPPk0ujQSkrtEQEV/GL07Gx6xMDPcyDnfUyzQBfD7O
Fnc/y9YR9GfoDp0n8BuxmDVDukG2a02Es1DQUTw+cYzwHd8/A6pSEeMYMZpyik9E
H/EEEhoz10h4qOEVwA1lPTvj5A9jvtdNxCguZzDG/AOjdW9iUPgBmZI2oXFRrISx
/XNz/UE1NCyvhK7FTx1kU3fxS7JN1vREYqUk7vcIF6iYKj/N9gnED5Zt9Spv5blR
ujGPiqlX2buA8EZsgQMVOvhIsWqq+W5yqI807K3m9jClOrnLaMOMPJpeHkj81RN8
YgITNNlL6i2frvXqJse/RlTf6yMszASXXYINu3DkTmYrjvxCvJgUqpo6RNMbijE+
r3MOtlI7Vabeu7QBXK6+xWntFSZ79dKLXroPngoir2U+jb2usaBv/1dYh8pAMIkA
QM2wvG9ddq1dFJEnYDy5VIhfUavcx0DAjs9+EnMisQ0QjlrEOjNDqvYLE+MwsxYU
LU+oRthlKcqHHwmthe+E0KY68AqWT2cjo0snQODGX3qIibLEel+ray1U2j0acJFp
65cpiK9Wu2oFpo/Sb2z17SVlW5m8I/2mI0MTP/4O2wFH7W14glcCH4t6is0y+Zuy
m0MwAP95RgHSlkjWB7f4I1Wh6uJ93Tb585bvDkn9BNn6cWK3hoO9ndJj3PhPjoj0
39BxsZWiUFAfUU0lt/cQzxjznYqFUSLstW7yxFlc8ZYwZB6FPzfDBji3NjzZuhqR
Na3qxfq5eB6UM87WPaCmdSHJTLqfGWoECqiD9s+rkiMirAHLCRSnQUAQOiTHq2zg
4NtTN1KvRA7pfBNKtiTVHxVHxM4N7B/lWlAn023FeiI/Hp5VH8JzYrWDBhy3l2d5
wWv4224wkXWpqqX2MVj+jsQjEPXICqQZPB60G8qp6wriOQogIOn10kQDesg5Lx5g
HHPcZsxochAZbWV5rDKo4Kd3N/zDuAwXeQkaCUwaPhJJBVfD3AXllT1794KSvYmV
Cnc86It2KQ7eMxzmmrXfWgsuqffE35yDRA+gheQu1KvUNilesUOKFJsP1kKI5yzL
Z9pFd8UwzmUexFW3hD2WGL8kbTFjehnc+YmTXTrR+N/qK7OEWJiWGVXLAEB3uIYv
Iu0rG5aw2iu1ZJjly/fTjQTcY0TfDWRJe3JnRk2bKFyoWoLVDeOthP8gbFiD4GC7
UvnYJlPP+1JU2j7H7g7bqsrTrXUtYsdIjp5WQeEvpOWpN3dgKIJ7bwuT+DBrYZTB
MjsF3AgeXPDDMpqs65oyJGl28IPMS1nUPDViBSJpXJfJ1DvKBe6+Amo7hU3eDO8g
Vcvu4TXtulEgm8QsazqS6Dc6UvAK778F33E6gfktHEen8CbMDj+T4TL+dBUhJkgJ
IPIw2JEkmX14Ppf4igBpn7lw9Sx0jXIIRcbIpZPOxiw26fLp2uHTCGdOjm5aoFFS
6BKmWSNH1sCcOroeHWL6iKfKXuOQNPWBROGtdF/OZcwBxrAxwYuqCS97U2sBLY5g
mF98G8o/1Ij7dqkZIW1dALG20PjH9ZX16HQaQNTWSYglL/+CjFNR0j9lkY7OOwqo
JoEcCUaQlGrGmiiy1UKB0Q1TJQkA8ytb8dUODoGN7MSgOeihwCOIk2jRtbrdKPZZ
g+cEXBtFIcJ9J69IyXr+EzfsA73YDjpvLxAkoVbhjrKKKC+ZeINSmaZk3t6YsHyE
zUCIpiF/VsnCQPhI9STZIV1/EGPDBOAPgUOhqreq94TLCZyodE5FTlXmyBvb+HAI
kxJROhYGAxfMK1IcG+57WRkA6FqZQuGS6wz5Y7ACi2eglExl5cNpgKjW+SUscmes
kNe2MDm2Xl+/mNHW3uMyydmdqE2IukqkI/7FDZAhe3k7JSO5xBYsouPkzoE8sZ8n
EQlClYYPftUCSvPEeUG5EEMH+4tcXZMKcSdfqATDS87At7YLrFuc0Eo/w5HPQnUH
pMmGfRa0EC7XOpMvSy+/odXuFlHYYNttLUMnJCMZ78Iu8y9Xm1PgGbz2Wwevi8Ej
lLx/Z5A92MX+tLno0oiDzYSz4u2Wtn4tTSP6Rb61CiKanz0S3qhA5bbfufB00zGF
GHE3aehBUl+SPx45jmpWmev1AauZzNRbhT5tizp9IBaXwUJ/roI9w87MnidYU8Dl
ePiF7i5VIYNSM+FYAVgHzQNi0H4PHhpdDa85pmFx2UAAt1WhCyRRGzp+LoygAEQj
1HF1QWIuec7Mqk3nNSluQE7H07MSZGXsqQDi3kp0bn/r5L95oYVgyah/05AB0qw4
dqXU4V4VbRp6qqBnHuPob2qTN1gVKwtUTGPAKWQdB7mHcz7d/2qX1Yazmy6t6vq4
DdWHdPYaVnLJYaIPGlChXV4SrTHF95GodU3NqFVFBrwVHY5KKbgrgb49a4IXgTmy
dQrP5SdEcUOiHcGsvhgAiiQGUG4aaSnwF+LbbBoEYobQ7E56ig7JKSvtjwohPPZw
s/lPlzWrndjSRUipT/3VVw5MGOmYMoniCSAmRrTWGWjMpoDoXwar+9JDvaKQCoAK
CMMRs8gmkgSwh1GbGm8EetnAA0JLU/tYGKDP21QbVpkeVn0Cq2ForweLOWQa39eG
u5ESP880jRp7+AZWjAhbT4egI7OC5C+Y+52Bu3audQN3qA9IbvAeJ3ISroAqtFiP
fy6CuHDaQMFdwGxSNCaLPg31io/bN4+V9vwXXNE6VeKzh8g7elwePTkABjYxQV9T
D/6aqEINWjY8m6/7HF8SLMBwg1dlqVNytV+Ys6UdyjejcOwpO8SU7vnME6V83vCK
eOzfTDDkIgp/9GX8CJWXG06KW+KbU7elcONx06RwrmNcAbK8utxtvmTZm8lTBb1R
GzwU1o9V/04AikWgvq+Hnu0eUzu4mjpnDDWV16fv65MmDAsCr2a4J0DOhjXwgOBd
EvVhNABLhzo94sdEtiL9yHtfgfSxhXnrRGDVKT0UTNpXvTmc3SSEd/bTnwp8jKgR
ujy4M81B0KnmPwnECBZuMyVExM7e+DY3udmhERM4BnkujDkHil+zRFd+xKTulXGP
MFQ1G1B0NyPwBP5dtZxGe31257aJE3NJhWr5CJl6E1516ybm/Bg8uwJlURBaA64Y
r0gnPC5GNM+rzNzxnwBULRetCaaEr3fkyzz/qfZZIKdLaLLN2OCFe9WsVcdncYjD
HMtRqtv4e4IqaSjE86ypjVhq8a/N4lIeZ9eEq8bmvic3whrDl0y3/ocQgDDuy+25
ItYZtMoUCTaKmldBAdihfOALk12OJSjCpPQIF7VJ+GNmV69tac/oBgt9BnEG2Z2h
i/iLuXS+ssjxfBjVwQI7Chmn1payZV4V84w5nhfLZQpjB23kj1zzvtk084v4r9Cn
utf3vcmrUy0wzrLbExB7XTZtmHW3b5rSIuZNmeEyF0HF1SCY+uGoyy0AAD0wK14c
1Kx9AoidXE/oHZMLI02dHLqeiPkLeJPBSNuLVblh9CmgEZV+t01tq1J0o6aSkU0l
b2LE9Br89bv4FbbOGGyF6ttLS5YfV66fl3eH5DUrNerkhtdvFXeOekGR2tHBgW2U
4bCnMDAN9AU5/ARLeM4xoiHSB9+1hCfREYF9xYb8ot51W9eUD0coiVtRWqDm4B51
2Wm3aLghOc6Li3+5LR/vv70Srg+tRW0pGu2zXSgKbPnY2LniZ3QF3p+NRmiPiONV
qp35o01xuei3aj8coJ0JOHHpIwqoFI9pS6H7zcajAOWEYv6qVhwilxzz0p3xV0N+
xRbMMjGdyeXRdpmsvcVEbTi1/n89426f2P58tHwKmGsGwvrNnhikxQP2B3dQYIXx
uMJoqW3NT48SweZRAHXn01egbnYznulW8ex4tFA85W+zUzG9OsTT8PNj2YHu45Oi
VNqJjZ3rW4+SqCAL+EhTs1taKAXcKNZ6hAzLFWMVff0hLa/EoE82zorpl9FajPZS
5mNc0QCTd594nDYTC/2EdZwRPUCtDWSZSZGNB3Drs83+q68SvL2Gs0S5DWXA3sCK
xVBaCQgXjbPiJlGyzcW6VTR3JB43AfvIF58aayFI+0sfDsSnyLQB5q7I/jDH82AO
ZgH42Bj++o2oqaMhtxzgvS2FkbdBHDzTPFVw+wqN19AAua7TfoY/ErxlvUXw6qBl
1KreweaCLUZPnV1M3LGxn7ttw3TIc4dl4obR6oGR6TmUdyantUvs4Fc8Lva+qEWV
ywSmFpMC8Y5cnREMV2JIVQJeYb7kOBZf3DSS6lyoKAuIuumzs6WGQ/ipDAoVptFZ
19tVZlYv8J+CmJCwaREQTtosAfVmhil6qK2NMg1fvE/PZ6x18O7is/icLKBne5gj
pJlRfFcnecxTJwe25o+5GmCET6fapC5sF1M4b65MMyjcLPvCM4ezYXraa7PSt6XM
UvkymFznz42HBmhHa82zYbla59qFK8m9jGtOFL6pE3D9s3xsxD+buIt366t32tGW
uD10dCbEgMvw4MepPtKlWId04jBWBYn3EHVNAYeh8vKRi+Q+imppRkVJ0dPsP2Ba
rA41t9I14zFvAYgSDRwKPM2dlzUyFnCpRvsCVuN7tN+Fisgangck/yP8BMUjhusz
8jEDOsx3bf6KDbpFJC7hUWQqAbuEyaLHUMBzMYiUAl93eOcL5lB22Ss3z4NuFZgy
taHBDIf+4a0af/HXAi5F1GXGC1HMLgOOrIgYX71stRdLmRHulUzLOhQDypQOBkGa
vKJ1pjOzF7/NCwywwNWTmQIZbsuLBdJxgkkzHcXZZPHZdTE8VoVRdKBxi0FjcyYg
KR1IQv0qUmFTfp7GCDJamGFa+sizWU1ebTYCgVLiCXqTjsp8KGuWfcpqd8ypJR6B
awaOY39XHW+IILysyE3SlOG2oyhn5mipXd2/dxaZmibvOLuEgk+umX63eaOKxhBZ
J9wV+nrfxlJSOY5kUZ8sM2wzFjKIL0Y9hf7IxLW+eQwdurrL2AdTfIuPkACeW5GW
NGG2F/MGk3nssT+efDI2KgxmjLH/yTXZbGVdcb3wrssuv39cFdCHey6S8h4aTPV8
6JVMJhooQMV+C+SpySdF+36pVbR3hoc7Lb3FziodQVZgBUtd+kwHlNiaC/QkUPxK
F3mcHBAxh0mAFn+Cd01/yYyYmdunUV8QK6dVU0wCYq3q1F6AqUHLSKR9H4ImzZez
BTDQ0BVk+g8SYBZcbiSyvad1ntCAFQX6XplvBg4sKyJIpHwL73AqVsrZ7O3nfsYU
Z0Yp8tDr8CLFMgQpAyQYGaLvzXMPuLzFy4O6LCL9uTG5pZrRYpkwX97zP5A3KtPe
00GGMJSOwDAxIbUScuepIsfDQqq8x5S8vJccp1HErsIETQOAg9LweTvmDrKTvWvt
0gGgPlYqryBqxvEBlkuq0NLOGcJ6xCXUFzs03kYclpV7BqRJHapAhypARyMiirEU
OcoJiFCJ1JYw7OC43jFyrqLwrT2idF++mkC4WbKF5R3c3qmWTA0II28y641lDPxK
auxy+9ZXu/RGR6+koeZiH2OBB33u99q4LPOgu3uuA4cPo0tVXcmqInnJd9Ap8k9s
cS0e4bx9twdaOUTxy3WhgORD+EiDKFbgD6wzrq2B5zkO2oDsLXpi16gpBxw5C7si
QI47eLpsy5Se6oDa90YqJB07Lvnia1MjSWiGmzwPOxGDzndn79x1vMUiVvJ701Wb
T2ZXGv/g4d17zmz5PcKy4wsDhuZ4PH4mmYgIo1QLzGmwRoCxpxASjAP5j1y+knnC
g1auoGc9z9C5w7xMEDaBK4WGHzZC4NN52wTdenrTJsGSAf0LXisCJ6u2WLkJYtk+
CfFFJxV5bv5tWJTsqPY60p+2f5bPMfUbEYXiB1xm9IX9dT9+h+yT1KYDWrt5+tAM
+knL5HWfg9awl56E0gsHPa+hnXSQen85rp+2b/uBjUaEPg/9oFO8iJX57Ij5DvHj
rwnpGSwYnRANF90Ep0KpqWr+lq7d7cu9bEkDYN3OwtSZfaeaSso1Gfza9VM2saxD
asceRv7ss6zequOR5jK77l/YCd6uqawI65Hc/Q/E23XTq+YrEHauKJnXZk7TeFk8
l50FLsPzIcXuwaoJggDVRTftTR1l1lM9f18mSGoMeaMcsWyJMtGHTFgluWJsJ2u2
uqksjMOSHCpzd+5FIMbHK+XouUEiMkXMQYGbcIrFZRXjS1XDV37y5U2+ACwNTD72
Rk/ge2lB7/rQWjZL7rqFEPZgo0KU5Rp40uKIi3l3EtLNRM8mcLPTDNTmyI9xHrzO
12SjS1wKqzgB8mU1kppIf9R8NKvn27KePzGBryT0rUD8vaorYs+H4UkQIhJWm9Bc
L0Smzm4L2un4zj8dT8iG45nbWV+Fe++Lzw6c+juYk8zXJtVXsFOgjZ8OgA9hC6cj
bl10FdEXteIHlGL6i7zDGx9dVVlDtSBhXqyqiOrR6A+gM2wTtVFa4TeF9IVNLpnw
n7q3XxOOOzxZ01bnzHa1kV/i8RLjqD+dP53dvdGcDRGs42dFKU7phwE7aW0r12rE
4w7+xR+ipBqCkdjmfUJrO3605o7jx3MrthkIl11GVuLl3dCLFYsOFcc8LFUZf9oC
25A0fZ5pP1Ec+u9z1rzta6fxgdh/8iOWb0euaPZuISF9+6RqDBuC5MHu8SMB6fSV
o/ezaL65SgwcZNjCjPBw7XOOg/2VoDk90m/uL+HAdAP5O8IN9Xiw93fTVSW3u7cC
YG4ZpHo/lk8vT5qeMOXEcU3pv8+KIeJY1OC16nAJ1JUfk+u61MvGaJLAU5rV+wXp
CZW+MAZb+MTF36F/dHg9fgURiRG/KPgHfoDzxAlxxYASSkO5ypHG6TjjVYpe5MwH
opVkcvxza17BsDXayKrO/T7NvH3wo54kAHiKtGA9EsjZJbbKoW5wVOQuP07UaShJ
2S0cz0zh4i5OXXEbSdyifKPBvnqUMnDTh4IcCMDMR6yPET0PxW9anP44XDeSlPqC
NXbfgoNMevK5BJhisIpb97G5M9w3E6rdJez1pLYTlypfjlxX6R9B2q8Nxj1SicsV
gpxcy2EdaPGqNMjvN4oH4Jeis6Nfz9AGbxBQsx2XBOV6n9EwKOnUF+HSg0N70NYp
RSK9ryvaFReaU7T11YCDjTiYrS7QRv84HrDQbjJtsMs7cFgUB3+ojPFLgcmIefIE
JF96bWFmLvbLsvOf3PI+pK7uOUkMmJAYgz22Gn3ZyGDmV962umm4Az7irDkvTRVm
0dMcttvMeIJ4SAut9+ZhBfe/NzrDtITJB0AsCP1cjFrOgsi7zsjUOcBxrTJ2Hvjl
X3WkNZcnMLTcHXiyn6X2Sp3pWmRTSl0mul9TJZiGogLN59svWHRuw0MQqoFnZ5Hi
bIYSguZiIh0ox5YnInsUXzElbR9rcOq0skIlP5i1nbpjjnVHeMziDXpRe846+iGL
kkAgcd8xh7EuTdT6f6oOlBhJk6Tpo7W3jTGUXxrykRJX+59fOLg2hTsoam+t+IT5
XfpCpDFq0cuuvoapyIRCSw61AVa0tQXcf/PbY/B/3o8QMjx2nd2T0yOSTtYxRse5
NAeNXa+/sSUidlJnlk9oXYui/QztIqXJcstWAWd/a7XLsRyoN6XzdAK+tXhBSQwM
LBhGk+y/eZSeY13A9g/hOEDCeujYDP2yjd1bUzdDWtTJTde3dlpegpU7F3hng4BT
rrzBpZ2eKPS4Jkg/QQaqQUYFUYvFXrct0axrJNLkGMwPQw30D0C8/33bqDg3+1PO
DXbIpc38cbUCfreFJVzURTswHFzQtyh0+Cwptn7q6ivCApPncf1HjwCabF+nCXYk
BzSWXWcJPUfqrMMFfd6m2AVbyflTvh45vrNLu6Tvf5pIMGv1LcPxWqYMX7o1aUAD
Vk941ZgolsDoN/KkmJh3gGGx0AKKVEMo1kgQQau2r8HptjBUdXVigRQgMFmeCLmz
72ExYf3B7D5VMFdBvwGYgdvC10VA9VOnKTo0pkaKcOlt0P6sUFoyVL7ACLqxel90
n0Q98pQG6ZToXqdvKJ84HlD+Q6tW1G0YFwa+TDvFSENJBLPdEhsg8XEWeBehcTwe
SdFmZQ7c8cvsU6FbpTd+ZZlZcZ+fx56Y3crd8IE8KRWexcVh3AHs3N6EUjqFiUMR
IjkbCc0jM9PJUI/cMG7JhMZ+AGEf+Ij+LLuxcKAKBa8OvcL+SS8jCACP1bM25Zum
jKbjPia5q+58sbFJg5ZnYZVCkp9AsJFUhKg1i/DSw/3la/kgqKpo/+XPD5l5BOSD
hKNoUF+qXQuatBKAzS4mt6wewDouNqDQxVQgTEeqvNx2zoRZBZ49oVIrGviHXTa8
Cm9/fI3yq5X+QgAzSrLH+j1ecgYlIYb897c1dwhXMGJMsEsCN56F9Z7HAjPS+3OO
lHg8PdrkUt2p+XPXM1phr+1x+1GcbGbtKRmB12oku96H3wkGiyq6vcOoZe7uSfj6
iaO1Mxo0Q/KS0KjoAwrFjAd9TVCb+woemBsWXjyAhhWYIwbJzruJXvFLIXMjGR3n
cl8PtU/msjuNrVSECc4jxIJtf+uoExgAg6Su+sq/1WmTymBoDUen+dx5MGBwJ+fd
BwCp/KpdIIEDmJmbN79y3imIFAXCo710aoycjB/5NF5XpVfxw+qP36lnl3Le+7e7
yXAKN0MSoyW+7EYrc1ieDYDFFdK03IHlT3y/PGFNERlanVsIg2IDD65Ux+xJDBlq
0fMb8mFd+NPhFRSo1Cpr/iNAFJxx4Q4RMp1tu6D2oHe0+uTq8miBAj2AQciNpvr6
WI9okRK+uiKXXwQsL6agVYPgFr5DUUWKhfWrD+lS9sfdhiHRJaL4KJRB9RmZKn2x
fO5q+d/gVIjYc3Ll5OLAKTpvYV/cDwXnqjhT7cXhmhQ3BCCyzB05zeYnsNgfpDOz
u1tLOkHEvNTUT1BrO3kruGemTNzXCBwveKKXHb1m8MUPqNAo90T0PWK/ho2rLLZy
85Ls2m/54uIfhMLKpW1yXhsgL10AqFfGk4xX54XQiPch1vmlMeXDlJDJFCcfcrYd
4KLn2sbGpyiMizFh9fWDVumsgeZjEhQJ37T++ze948UnvzewMyH3ADdn7/lGEFnD
cLsyVcB2H6HTsNoWUfGOQGZ99jBIMeKCP03pp33kzSKEHD0MMVx2nMa/RnhpjORm
cIhxsGiio4e6QQcHtHxHOg82GQXtc+/fIhRVRn6GBUhhGhkhQzKdLxtpZdFJwdVk
TJtp2gmqyAnViA0lA++r1b+H35hpKIRvB+c6/mjbRI33/dWuZoGkF+iAHQHsEfRr
SQJAKhU+JJmmnbm38fk7raKFmJEULnWGZha+Loo4eYYmItkCf4VL+5cu1+Sn3anY
8MoCaXfwRqUjxMpw/RZSUcyJjWzYn0skjckgiETusU38xZBQTnesEFmFLrjzwQEy
IhjVlumBOsRwP3Uo1b7tYUpovyR4EmYymWW+43bTHoncLgFkerkkRN/bxeoW7Zrs
kJY9s/Ix0EJOU8RL3v8P/GOIADy5M+qxd7kaY/QjvvsNa2J3MHelgr0yLP1e7nE+
75aTPnw/9BexWcrCLwx3mFbK/dLFFgHuQA++BFv3pyPqDyQViOS7+0gcViO/go/C
YRnQEsIs73TKVYOiF9HygAiUUqUIITzJgCvrwQ8SdLt8qwi6enBnpccZ7RvU6wNv
YCAKxpopJtBxsNN857tILIVQ4g5fnSNerhaw+g/hdmT97uJ3lYXiJ0ujqq/BG8H1
ZduFU1jxxKbU/R+FFiMbOrYm70zb8Wdt//9z1zvidoW4WA747S1no0p+IcX+By8L
TYz6uFKho/0AUYDLZVOfGQiEFBFr7W0nIQ0boNhn2zGtIV296m+NXVslNyh6c8J2
sv4X1z4E552WfcRT7wmO/zr2ABIJUBiB9v9H30n/Kr9hr8zzLE3Oae97xn75VRpY
0q9ObmOuOvgFBj5OuPOxoB3SjO+yGCXLa53+XJi+07DJJYBpuJiWvsIiOP/hEzJ5
IBUslKGYQl0fjblL6oKXv9I+nr9b3UlxLnooc2NWAytC+/sIV0SnB1EBm7zNSba8
OeaKj4A+PR6N4IEgnXDfrMEYEKAKBJFfED4zpwOgw9t//ZhC5/4nUmLJv7IPGpt5
jVXD3X02X/kK/pvBNrYrKBh7XotJ0tIFbDpUTUDsz6efatuFe/yMYvQt575ppBsF
EdahMlczpslVvS0cfE0GVj9sXLwGfkLTRRTqMC2KV7rcTAhn3qpETc86/e8VHt9V
VRUCV61UriVFexeNhzQrZ7mOE/Zjpz73CHPWEgXBT/uvga9jfM0ojpTLOgjPYFLs
s3Ynz32f/jsm33NfyPExgNoc5tD1ZYtEv/jWJqZTHNknBPtNJcf5kEpbnxpHXd46
+GC++N+kQlH2lhq/R2O8HTvGZj2urY2ARYxaBk4NYOHZ1NDhWBYGjju8V4zZPM5s
GK66Yxyk+YCY30fX2MCIiXgvem3FbcbSM4F/KHtilK7bt5HBOOd04TxKx8KLnZRJ
7AM+MAFf5N3l5iFwUPuxhC2lish7WiYRJToGK4/J8v1G5BNBgdDsH7yiVhGIYtOc
op6+DLoZWGDN7NaGPj7TmbUexbHTcmtj6D2O/exyOnL9h+UbLZBcoT31Rtf1oLZg
RBHHlSx+GE6hAbph89Q4cix+rfL9snOAOydwEMPs2h1RTgl1Mtzm8uHhuZ4jW5nQ
47f/IFIB/RnjVagH7ZS6+wpzKSNSLc4JYO4GtfJmoDtekjlV8aSB+wukb6M0BaI4
cKhRCwCf9Mmhf59Vl8qyqiuYhWAWZT2MfHwRbFTeKwYOFZ8u1LOm6csDnSokRVoY
3a6AQn8KcMPulQXXeA+rq4LaSyqK9GhBZKnKnqZKDphS+9GvbSL91Be3eRjwDyIM
viP6eiP7WuzpvkPAHhZUw6CnVU3LIelCnfRoskemBT0ZqZWO44H19JaKWDLeFzDA
p/5d8rWDuvxKuksG7LA+LO/WvObuG0iKo9kfiRfqCdpkw/w/gcxH67HTdCR5vSZT
kSRHfVfT+fYgIeQGZEMSIJx+jK/QOHQ3CL2qdTsJDBAiFyreWxZXNNpR7A3zGbC2
8do9qjxFBnwDRmSTaNT95Nt7FpE6SqPiQmddfaPr2fttINZbyFFdzUlkz0NhuiA/
8z8iqSdZ3XF7HGTWfCcGQLTW0tue+zpAjMvz8N2gupmfJTfx1/yfmBM+NvwgLbyB
pYszvO2j2h8wbJcSA7Iu8uk/rldR0Mz/53Upd+OZJ8wRAMR4JeIW/R1WB0xAWjI3
Yt1N7Ng8GsZupqiMfrXE5I86pWlWh9O/XAbIMVIo7FRT54/3bZeGUTkh9thFUxtl
937g9NiZ3fqvy6O1YvrvOPEVfvzd6RALch3ONX2d4N6M4G91Xy9/C7w7Uk7p723X
3SBLaJ4TTre+iptVY6IGv7TgRhfkZe4Y+53Hjm3fl3cYh1OyidyffG2rg1/eIQZT
O6eVyy7vXgLHpn4KrJ0/elU+ye+GMOAz7D059TxWbfH8yKXvv07O1wGuwqBRnFAa
ATt3btKrhVPD7NPY+TW5mBnPo9Ry3a2bdGiaM+qoCa+nmT+lw8eGkG42VFtMAN5/
J0N2pPOLq8Qddb06xx0+Ox+QNxrID9meQ5GQ/ZaVnu//uyt8Fb/8ocoG5tUIQzkc
mVWOjWAaRwZ5Ux8rouV8fdQCQ3+L9Qy+KvhJGxxiGgh6FEPSC5Po2n3ILQ3YAiNM
XTIM469bgAIvPVtLZY0REnEYyPe1xgmLDvy9/KKsl0qd+ooMDKUJvGTcmILPMqut
Xvy3TkFcuzdzThyX9EkO2YNerOy+kgiipc7yms8UylhZCzuY9ezLeideQzmBhp/l
6VsT7Gt8UY30Ofa4oYeEDgMBEz6912MOY7pg01lU6dOMf3WzEcPlmkU3zr4w2IaN
jtopN143eauTgSPuhizlWSIbwVtKmXrxIfGP1UnKzOKBVr07aHVecSsbZBncjPp8
WHFnx3IQ0Rb65DPIf/x372sSAP2kN6P8qit3UklHoKpaTY+vp68HPW4ag56RN7j4
h8jj60vxhFeLoRL8KSUfOU8nstYF1Jbvy+FpIXepprVGRJaTvhPmr7G2c1sOArdO
GVwKknjZXTexFtOY/TVdKEkSrk2BRgLmhhqE3EpH+OTQEZeBvnkTugcDx92iX41m
qReiVFt8k9iAS0Sa60yAhOVU8JeYEP3NiBoT++SG5Eq9zQqK4qJspmqkMz7sPDQ7
rVOp0PrhzfWK/tVRtjEA3tYFZYvRCT7P/xM/f95r3pS6XMI6PzSbD8qN2MR5r7JN
T0YevrDAMF/Ku4MgbyCaoCvIuCgN4P0uHE/ZzrtJX0+G9ksHxkGFwfb1G6Iiykid
PkVdzJiRt8/xfc+7wTdR7JSUtnXK/nzoXOmVEN9p9uQ5IxekZExH8O4weP2rgwlY
q74hGwl5DJxH9pJTPSpVfRsWPJn7li3AUfKOTSj/RKSfwFSD/ciC4z8OEmUYVYXC
yUIRTlvM+XRK14ddS02vEsMUCA8f0t9gwwz+RXSNyAoGES0PMplRCgSZZYxFkxs1
GaXzzLy/A5PUbNLv3s4X9OELOfxXTLTO8WJsXbvpGsJTLs1VuXDrw9D7TRUlHtsw
dFXF2x5HCCDW0c51gga6VmiE2Rmc5JVk0xfnifl+to9eVF3X+YsC3nezoWFBLSBb
tFcz732NbKg+k3KvT3fdXVkYDFRJ8aqby4RjxbA2kRz20hX5jvvG2zoUF8loBQY9
cTSsgx+87tQjYG7xBIiyASUXqtq8lEdG5oigJxLbBQUP5EghdyvCSF8BQEt2hdib
P+TwS5bzCic8iPFPBcBGN4NWFD77Hi/NEG+pggeDOz1fUadr+s5GVTa+RrxwPJ9+
Oq2+MrTOyuE/7Fe2Jia3ajZZPUYBWFhhLiPv5qfb5V4KsJVIsgBu+YfMcWxGsmN1
89wo/MphYAcWhL83SK89cSR6BcyXXTYeAuaXEqnkPkhcYS1UxukVdzEwvvwywPOe
7Lcesz6FscMkUUeCWX0a5zSi3bBqWgZwmQ36idFRgFc+p/0sWgHPO8QVN//EbSwR
EN8H37LNm5YeBODES+t8EBKKMwshpRb4H1xUVHq4753OQmWC6yzuB62Sfrn0Ffz9
O+j70r/UIr94RJNbUE/q009sOFWc+2xBUYbsAfW60IhoPB8ft9xNTUPsAliIANda
fl/BEY7wdxvUkr989wT4O93ZUw1jHYoWi+N2o1LWrby+DcrbOmMSPequ0CF/wS55
jExoDSNzEimJ4Q+eNdMusrJNkaJ9r94BMTtvoQ+44lTHskeoTDB54QaD1pb9F6oS
psMWdZy+FkqkInU4f75T9hAcfbZ72obbnv2q4jX5lyBBAr9z0nV4UHyRL8gGeADN
h40jVADAUDJcw3M24netpydBHKkfaeJfyg2vlElw2vjiXLxZi461T0bSVf9GMGtV
srDSD2wN8OA3r0u2U6uUaLX9+PPKxw86rPstvcNRLEZWiPVukesAoICm7kOjFwlk
/O+GYOJ41B5vwRzSFeFAzGXqGdYsZLPooi557gFjXv3a+EZO0L31pXR4e8wIhrR4
7F+dJ9z4oc0gpCf5BwpMXPR2NxPJ/y/fCEPNWGpZGq9GXgWEJwiPj0CHMTS6IOsO
5MrpeX7NOb3ncpWlNbIy4gr0SHny+Do1ol6SLtg2j5ogC2fZKB0VilRZ28z2e4E0
q/gFJJkUSVcQnF+Y2VxfZw1xpbSHEOvEBkGZHiQUzWr6f2eUCf2TW5STrl2FJQ8r
QkmK9D6V89u+Rq5Prk5iPwRMtfidWet7hg66mE7Yz1rRaiAFKxf6PpHQWg8tmmve
clDnbpi8nViwfVLoaNSKGiQRz8Gg49nueq7DefqxFgWo0JqNWRqXGUQiRqWq33gq
OkrA9yN/Qu/wm20XjgQvo8o6NCOa+Rc2MoLRINikTHow8t2orgg1BYmljIDH00gD
ddiU0gE6/YfWJqBjkYpqJg5v+c2YpALgDClKS2FoFnTgYTyz46sotHEGow/ETHf1
wQOsVhdiCEXHWX1Nfc4Mrqz6SGCo1oHrdgnMbI8fzL2cR7wEzmgNyzhYxzSHjyJr
ppfrObtsrcFNKyQF+FbySuqzT7CnDfcn0kb4RIo1eBBdiZ2l7DIq/TD1vZC+6t3H
0ZJmP0NJpJfGhxyX8n9PM3lx6K+W7s2UQoHzhODqwn6bbvYQ3ACtOLmvR8TVRR9y
0USJR2CT5a4p/dClOwSARP2PeorJCGuV95zyV7d2wND5vZlc+mcmCP7k9ZZGRKCw
KOcs/Yce5HcojxUfaBRRtNh/jslrdu+D24B5fkO785Xbtzru/XOCQsPtq65J3/YO
/XwaJWAD4spqmlnBcUGY4ofUgXTHyXS11b/FDYwr0H4NZ37uM4fH6quZ58kTBczn
y1smp7AhdLpjY6H8s6ri6Vbi0cTiXc5/VnvVs3kGcXPRWEAb/MCPXuQ0rnoZvnMS
9j+o3tR5W0YE+NNxeEh4gXjd3HPswr0Xi9dk2qlGSjeFEoTYRaX313PK8+eZPQzI
gOHDD6zYaHpoyCAl2+H1kxfw/wV4zXoFBzqZaOwfkaDJBm74kdfcSPzVoEr06QGJ
qCUOA6yc5u3Vt9RNfTxu/QDV4D4jNoxF2TigPMwzeRyZlXTUsMVBV08RLw3xCyZm
9uDYlmbArxNH6W680DvDx7zEvgClYdukL0gGVDQqG+sJdoqvjrIvbllBKPa0W2r/
qx3QCzxU6D6FLHbUBN6ZG++BEos2rYUuC4v3itoTmR4217MvdHLhWUQ9Yadl8z3b
2ak3AZdddhj9Mc+Z4AA1HDlfJbEEp7tTnsz26w/vxoM5NOr7cj1H3FUuMlgq0d7M
bwY5bxm0+JJCT4jnfK/7cOYSxtz3CN0+RRD5TqZ1NPXS4+OGYu6BsHuhjYYRReRI
gHITD2WnbYWzk6df4wH5daid140sUK1GbHVvn1IBJHIfITL140felUI5p9n6QdmG
3fTpP6td7Gg7duileHIACJCqhD00KviQXIPt/3Pk456NRhDD5FLlQt7JIg7RQl1w
i8TjiWp7KtDhuOfwHOIelela7sPwfuTseHyfI1UDB9GoJWxSDcn2fU99f2YRqsfS
lV2ScnZvaYlCiZv4CA0SLjxl1SkgGWyoTezJEsy97xYcNxzdxp3TEhDPT1dZKdCr
A6vJKVpMkjbx/XW2+3veJBf1QuqT8KSaIaIyEhw5n/t0UOHPssZeU+Ta7b9Fbrm9
/EX8Y2GA7Rd62DcEkzs7vOFWiDSkpbFraHpNkGIrQZbzkfSNAL7qSVKHW4aIk6tl
04tGZXl+6MfvJl5WMeTKa0pj/x0hukodyGFzfVfaRS8W7+lYpjrRK7uL3I97eS8V
tbOtNGWT+DsdTe3MTJ+fNnxswQ/N+u9HzH5MAmfHiYTIeAIWkKRMIVof9xLivq7J
iOmtRygsgKZ9xbPFKb2MW+UoM/dH7kys4oTs9JUOsICqK5Pbm58qzSF0nDjVb+hh
gLAuvPv9IA4XUKk6mhDBxVuXeAtdFaCGzw/N0sTW4EhXzJ4lHRmvYiw4WJpwWUig
B4+Iz+kf0cmal1vsEfXzQM5J7VzNiS2YgvP80hDSWlMtL6cU30fDdHPNYZldH0qZ
Yw8HMXgASRH1N0p/M3Yazo7aOrSfd7Kht0DuGo7rBw+JvV0gCt0+OilAiG5vXwrM
PgsZ7cvYi9QDDyJq1tMnDpLi+s6OgLDPmntIaDaT9oH5YVkekWI21xU50oBK3Fc+
fYozxfVw6uFZ0o/4vPVjTUUPUP4bCKljl1gIul48q/YuBzmUpo0F45w3RXMJsymH
VM+UUTKaaNzMDYLQd7iLAYpzu5Y8IV+Y3AfwHGC5GjvN9HVR7j7+Umd9TOqg0a+a
hbKp6NmXKSmfwHtw1QVXjh0J/f5gWlgsL+MYt4qcAUR96j1K6N04Eh3RIhnmHAi3
LmX9P3caBVrt52V+I3gfctuIU/4ZlsZ+oBPjrMtptRzqmMUCly8Wdjk9j31ai2mc
QSvnRiIbwA0aB2MJk1a3QxeZLcooilejIEKtwZI099Ip6DmA0WDoVH7Dy+g3nTZw
IO/x51dAvT+EkFoOnZkx+XqgKQujyz+dEFAFaMqquzd6MCJis23X48j6G0VowYL8
yMust2CPVVYbT3nRp6EY0wJHXEcy/V2IfRI4D2kvVSTs0QFLqVFQSUmo596bxzwr
qA8cdrpHsW2koerpVR5ncPr5Gh+SblGSY5/Hd1yQr9aa9tOszU75+TMsVEcyW//e
S3KHlBVJLVwIc1hHn3fZGhXtib6/n4cmyQyjnkhpZ5/Ju0MhoG72FBhDLvEQHPpF
CjcIOaz5SrO3RHXnBeKBvZmJHdZIq0if7+6MsSaiG1LNWuBwAC02qJ2I3S1godEx
7IBiN17fIdNsNsJIGGNx/Omcx3xGiWVEIFSCUyRRWVOtaB8zcmgSnaNbphkhC5sk
7izIHFva3TwWIrOe1f+Rmc5Ej08LJZAebBzSNB+XRzhpmgHFLwvTQcRcIoDj+R4a
/7Av0s1UGGCTsxn3c//Mccu160Vu1moVrlYpL8+Q/L6vH15Sasj7IswvXJnZKd2j
ORMFOvIEEpIEw0/TJTRKJbw69a1wms3tD0BityrpdOnjWtE5HMkzKGAHKAaaJZVp
Rg6Qxd9G0C3+RJCWNDJ8Wv4XHPo/MYEl3sCtRshi3QS9d7ylTbYMAp6llv/KNTd4
mbp2owjh5KqaABHGsiT9OU6re1INeAJOUKz4WVM9LlnnFrAIgASxy9MWCFY/67PD
r9+hDznlnIge2KB/yg4DSB9uiGFNMp6iH5RyITpfD4blcj6TAJous3XRKBDm31pp
l74Yv0VcyicmsSe+gAJ9D/IhUe8SaoXN1/5f11Pz7TWqr8zfOdSspZ0wwcPL5Y3G
Rzn8Nfy4VY3L13UGxX2xH/sDJnHnsJohI/KQ79LlilnpzLwM0scndUVs5upNwBnQ
jh8Synn7ekeiH5rue/xZDcaGHmHcQCSquzsiYI/hkMbKc6ZbnEi6+EF2xAbvA5yD
YB9jSp7Z0wOfD1WYfWw6xz9DYGt+IsjkqnMFDBkcbq2deZH+pdyqj5FuNkNICobP
D8CCwCo0KVyD0Bs5co8cPkxhZl+vROAcNOdj61mpmuYReQOEOVlQWfOT9fpwgh8B
mN6YdMVxEO0oGJafKcnSXZ9VVWRj20Dfm814k2nD3BfsQ7xyBF4M6oIBiLdvOQfd
PR4bfSNTOkBlOinr9QqCjYSL+rUZilvz0Ct+DFS/M/2LA7c40R87N/h/n47GmR/e
iR1bS75rrlPJABJx2mX9vtBmvKGQAns8GTDBbota8VejYP4sdDiEPKAMkiVVXvs2
zx0oFA9bCc8Rz/I4rRgjgRtaGJta414VSh1LPaRcNsu+Hv/Z538rIqrA66ZK7fDC
6X0NIjGLcyJnIB158ALYRlXT7NpkgS2Vt2r4wOuyHLZNkPQxikKvDbK4xjZUA/S0
xg8JwxeWGQIm0ds0t3sxE/htPJIqx07zYL9kdooLtaC3sowmKsWC3tQ3e0Of4CXn
tgXMRpavNk1zbM5JC+C5blYEDvKpxfdf1H0M77cPGFl+zfbQyFm1Rkdsa/ovz8tz
KHDUA4V6Wf8/JspZxF8Mp8omZ/dDBXWn5+nVYn4EQhnDwdNYRTH3C7OGjpn/TLCf
TKFDVxMRh1XFVEn9DadRt/alEMSwR7EsWigv3NzAMdrqkOS8ZYtSHgzEvP4aPPKW
BaqyOry5ppi0/b/q4WC8iz73TX2D3sI9LTQY0hVuoigQHpGb3l1Oe7f2jNQ5KIK6
5gPWkzi2plt1d0zyOjibC+K1EMQfQjTQgbWN5RiU2b0bZA8AzlLONJS+Mqqs+/23
xSqTx08ziRVdUGO7K9eURZL8nbkmn+IUmBUYDL9Qy/7qvn0sfpW2oAPsQyWFvsAt
VxMuyROVVpMQncS0xxXlBLOGAZooJ/+anBkm3kRPnyIXFBsR8cvt96elsNNQvMoe
d+kaTKLPCAtgQWDMiGzKT2YuhLL8YtdYaO+ZA+yFOQC/tAMaWZ56xrfKWIaEs7at
h/OMwfwKQM5z5+RDOqpR4jRqenK4QxEVQFEJF46eblM0I3QMqrzgtnslj3xU3qgK
N9ZOzKtEOs+JV63JAVNs4/DKd2r5x+rt6Tbuas1JqlnDXAQlZZE3vlBK1BOMrGEj
Tbakkl3EdtzuOHeJJ6XXCnPII4C5J4cLk3AK2tVOubroxCbtS397M7WmUM7//yA3
O0jOEYwpGX6ILIgXFNbRI6jzflLIHCdxNbwgKoGPS4QnsmVkU6WAuaZlcz5W2LKV
VjJymTiwmcn0Rm5lSfHcnuAp5HBavMQc4DiYUohCp1cmN4T+GO37tgXEhQRydjce
FE5Xow1jlADKDlpVu8xO7f9XWdGvGl1p5cIs1I12aYvlWxRG1a+EPA/7AAjRFjnv
tzfWPugsQTwZnOzyYAo0WSp9s3PHkObdv9msSNT/ksZamP0pU1pmU3sD/JhncpFK
GJ4yvlOw/aD01cQri2QeRE63H/B3hItLgOHGORJl/lvI0PfziRYEng3pnNXasQ7Z
OtKGdQHo6zPILEjIuPQFbYH7olx8nH4FewPb1Xn++QBWB1wWNkjXrDAY62Gqm/rk
s/NX0Trp1HZRj2AjOddQIXCSsMWKLOEXmE2pqsFbqb+WsGXzlTlElHPNnjskRpgU
P3jkdtMcIL2YxT2lJ33onslu8Xsdxp9YKOmPZmipQti3raThsbTYd4bPkwBXAqBV
/KJBleodpNelEUO3x4vJyyJ80VibnCdZcUJ/KZQaFobrLatM68gyvw3aFJR85Cie
3Oppagw2fo708oKOAarp+ErPDmnxI8aPOdPBG4X0dtz1GUJENyS8kvNbDOcoBlEr
TvjJ76m/bJ93EJfqOBqMAKqKsAT96/4Yi4Q3egk1NagJPDcL/nYOy9EuVxL0Um0q
ASKwwXZgCWK/NrGeSmnm0ZGAY6X8x09OBfiMdT89mRST6IhUIUDM1g6WgUpyzmFI
XFQdgNsS4BH7rEqM3j9GvwzAs28Tw4616Twylb7XEnttWcd/ZIIlP0iF0mqR9Zib
yLSlXsaZPBgJSQ6hFDejDj5KeiRnteaTAQL/ZN5SqE09JHv3VKVIc0DgfM/HqkJc
GEm9vKCTw/D+jU+oDemvCmA3PqW/YEW07cyqp1zr2MHcgzBx20rTGKs2cYmpJoYA
qCGxZDTWY8Mr/xaJn5Ao9uuRE0W+NhVSBv3Ewvqc/X33cE3H/AJNZoqTg17WwtpE
VXqPsI/bGdSYNq9lXPP/FAY7coU4UCaUrRi4A6uyHg8WNc4YtKcpcKa+2onVeSSR
tqIlvCd/PGJEu0+lnZEpVb7LSILiwTz0RogSOkmKZIH7eYx/+8Go15Jp1A5IXReM
M0ocG/5wUkFcqAapYeL4wGLfi5j+g1lYu1MmBpcj6ye7AYXN65niotjCEgl323++
APcgtNQAoKy3TOKMlSd8kG/j5QKlRzuYsq6x2a6GEnYN8uyOC53J7SYEJLaisiOG
2Cj3lZH10bvJnLaxouV5LdKn8Li/yW1lD8DpCddI1/QGW0nIAb7T1OGvRRJghECU
dqUO4yQ/V+dhRhit4euu+OXeNPMWAxs4v7Rb6/X3/84Q9NGIZUhycZtA8d9VW9xK
V/ADqBI7cG5a0Mb2jvZMD2cqXJMMS/hobflFbH6w3asQQCUwhTvmpZwpTOTDhigu
xmHKa2YIGt/SHG18QN/OrGmFdL0QIBoq6qpkN8Rr0r/49f+3vGIdDtdSSR8jiIW9
lqG3fXs/I+2feb4dj6IcT87RnVQ0XQP9bzvXr2COquzmpikRmFMGzFIEOd5ZwT1T
xWhN0pooSuXeLs0BOx/UHQUYM4hTs1SdWsh/VqsPd/U9m1dy8MwHx/Xw2JFU0Prq
96esFFlwFjWQ0UWId0Clih2/HA2nbZAOsa0REY4SVoXObJJFvn1vaO5puxxfN6CH
myVMNHHaVxzi1I9hhsHr+CH7j4cbLoOCP/8qxh+RO9skicbd46d5BFUaskWKYA1K
e4p5sTw4KRa9rCu0PlctH/SUsYmcJe1Ho/+hZnMT5gZdSsRCYEjfGZpDH2VyWaLq
d2iAVA/C1lSJiT1mHOQSD+VAhOR2D7VCBipG2TqRjdcJ7uY9QZO3SGPm7W8twU25
ryzmz2CY1QFyhOng16y0H/qy1EimFPbrnaX/P5tOHR7a/WHAWdFDypQfEy4CUDZ6
iHjiCtJPSiQPcTJqfQ+Qur3iNYEMaMMdlKRbCIHvqVvEdHRoMle3eoHANoNaz+SP
s/NP6HL5NVZbprrZTbk2HxjmDRtwnIam7QtIBhMhCJ7GgDPO60QzHPGJlWEuRQP1
VbFOqBFkEPK08yr63W2/uHku+3xp0B4NULraPrgpjOmfOWZBkSCl/fY1EvSEIQ0F
NLSzbtWdago+BUJoRAK8k6BcoFdHcS/1fdGl535UMgPtS+h7ygI7FBjP+vQ7L9XK
oYmDtfITgchP3t8fRojc16Ic1+RlpVTfSBcPLH00wiSnGdaXUtLhANrWQP+AHGY0
/7Hdh9AasKHARmGrrU71QK2b7ZeQHQJFXypmdcFc3xcku88ud/qaqc1AzPynhtJt
16PJwH70efwAZVl75E07I324wqeHR0OHGdTRCDm2+p0r6oP6ngcHaiYT0v+J6ekw
CaVCUjXIjRndYrKciubSkc68qtsuo1levzwnAalJN8vwwUiRj5bdbz04/ka3AQjT
J5hwhJwg37u2E3BTh/Ude6u4TL5CC2GdykJFXSkVkxwq9nY7nJeGHA2gxmDO3xUr
`protect END_PROTECTED