-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
c3PD6fPFl/mQIPtJouenG+hNfpGaI3utkzhqvC37jHl57FD+JH5ee3i8f22GGKqu
5OKQ3qSkaq15JZ5RwqBfb1lYOxm/UVEVnNNUz9bUIiYoG3kFIpjElW/DLrsKo42+
1hZoCEEnOFXwYU9+OdEp7XRlkwzV/sBt9nt5Kx3QKwjKPgZSbF977A==
--pragma protect end_key_block
--pragma protect digest_block
E8N5Tofo9OjwVtb+JSHgNJM1mhU=
--pragma protect end_digest_block
--pragma protect data_block
NlhFLNWL0oTAJ7G9sZi/eiDa2GFXAPIvCAK1KTuQud7zL59aVo45w71HVfOhlfs2
FRs25jKuQQcmgSsbxU5E9Kw6k8ZA1R9uDARc/tdHDMMJea/fI0AesX2yCca0Ai0T
86guoisO9w0ulfP4jl0t69eyCDmbXEzBGVnrBxb9U8wdo0VcermvhaNfPa2kSfeS
tDbBBMQYKJzkSN3RPqOBnJ5VZXYUNsj55dFAQR1An5yr2IjJQ8qloMXQ32hvsxDs
AyJfe4kOkpR7evC/0H3RRa6yYpxNAfkqMphfs5Zd+6wiML9vYVukveOSKA1H0pSE
e1EpdqcrtusBnc3g7qmaDuUDYaZvRW6Ky3e5SprSEYuLxPeuLgbs1RSfoSw3uE1p
1zAVYJirhZBAIagDuWluXEHbhqPT6IktADaKXzaLRTeQJdLTI2VZaKqV3y1JUEHw
9yQDQVjpf4VgZBtzrCT7ldQlvNWh5uJpclAdvGDSuxGULgt7QExdRO3koeSvGqVE
VQRo088pv/5mv13sRFZLyOTOgL5VVHxPYAIqehAU46mEmO0iTBkxgK6ljAEgNRs4
hx6EqcQAfFyuDzRbamlkzEPLjQkge7EFnkrRDXm20Revn3Z31JP/AaVjAe5ZJrWF
ywEH98rODQDPAqdsA2FGGaYPD/Z9/CLxXkSDTaWjA9rdqYBzemy7a/rU1ydojLNh
Z6srdIU9QBnXdy6LHZTxH/ZbpOuDmG+KUfdac8102CDd5JT2HE2zl10EI1mT2KGS
l2gYgIejJYbwhnh/r8+FO9M8tmiHH0Ig+5/KHECd/3BvwdtiU0OTLoAaOZLRDKP5
r52StdAht4FvbEHgSjSRmypGRoUmn1OVi4U9tkCB/Azg+XBpcebLP9V2oNqkvEEA
8QNVfmYVNfYludsfJcj9WA5iMTBd+e1O0zkxtP3RxTedrugoJVp6Jd+yJyznF+qN
rVnLyxLCgTgjmPb6pTdFvI4zzkP7Wnf1BfTg8ycYUm2P/ir8+HqcpmXeqI/oPMR7
ynQvZm4fsJ1nuOcIods22r1nDddcPGVcGkLM7f9unn1GbufaZYOvU2IBv3H78EAy
uU7pyXJl+E2CPjVRxZqAl/TPr/789AILzZeJjG6HsEesdaXtrZlcw6G3rwTca7qZ
AyKYEZbxnMJUzVDAOkNWy+iNuESPd0qZHVKIAiFCmGTk8PHe0PQI+n0aFHE8ejav
sQXtyvr6FSr01kGFV9cJEQg3dHyZ2lbqNH6KEC6a87Gm29Z877Pgy6uodVFx71G0
LlmdP8yoKAIV+nnHGVgPV2UTwH3ZaBtNwlJZxl0Yu5mcXVS9IBEnwaPn9ivWa3gG
ZGFFVpBShyFO0NoKGU69FcGNO/Phg1DmEUeBcOQF4JKHsCD9916CxCVsnsEus0gH
6I8Daggh9Ol+zhG6KO/KHs9GpDnJHPahlrqjN2/137/KPqjr2LBmh0DdVvDeUWSF
Bz71BUNbI/P5x7AzDQspfvpB3XVS4hgqoPb5P8RPKn/KmpHGyvFzIUcV2eBDW+0l
QUbSAiu03lhYD0pqwJglbi+4EuJMMKr2POg+EvkYAVongtqPuIqrI8qSgoTNV8FR
vrxCtLQygAStmNMtUD3B5GwGU+et33M75mVY/NvXb2uv94q9cqIBtz5osjy5mTnT
hUniRCG0KJNRBLQMn5g8/ot2tJHArTqUpzpXUWP8cxfV593RJci8ybJAh+3s1JHE
Okb9SHENQEnNPj4sNN4Xn+yeKFlaFiGJTcPXXWIdEx0UVaPRmwORUDbaeCKYX9xU
f89A6kKmK1hArCDEkB+IpAoKBTppdi1+55vFasqnfYEAA5qls8te3Wnjm0FrxfU5
AVSr+DN9naXbx5Zmldy5IVUA4HZ67TQ7mi/2NGOSEbM/UO0ag2SaZSeLnYAzuR7V
SNw2RQ+z0JYZGdk6JJSD+Su+k/VcuW3s87BBZptiAYaB0zqLubO08Zb6VCz0z4MR
N1NNsJE+6ehVaQ4k04ldD5SeUYD4kHNhXWtKWpcBPIklu0OqyRmr4R25UVqzsIs9
Pk/OfOn4MMyW548+OkGqQcOBfd19t97LHJwWJH8ey5Rnw2fnFv0cVm5KS0I3WD0O
xCXB9nRdUiuM3gDR7oNjFH6fvOCMlM3JxoICmd6XjeW72btU/mMr3ZMjAS5olisO
71vztlY9iMN3Io72N4vN0+WJ0fDT0J1wvo2031N60fyvDg4TpFdH27M+2GkDtcc/
1GmpwBoVAEC35xHuvTpzrSW16/h49lRpNhEd2YZClZvXC9zd4EsUFML+7c37hnBY
4POely8KILgezQCZCMbplqNprWEa8eFCLFfnDMc8sEdiHvD3JWAtaPKwKnvxIxNL
a6Pez2GroSrLRBpjcc8KJ++suT+ZrlXbaZRBZGt7GrwT5GrNHQt3XSi3JUREb7L7
58v285N8Ixu/KDvJhwLcMdvdzcexb32tyr3Yeh+NSVkCitnWIyVvul0RAIGZV+E1
gglaDhar3teIv3DSpy5vy656d4qNtkk0z3n5QRa2xWsgg6mHy9YJ5aRy7utEiYmG
FISR37WAmljxtVUXfn+3yOLSIRxhS1FoGtv21HMHn/UODBWgxMmgcFS9EBL5znK0
tDGO/DaQgKOHDJ5JnnAMAK1pE4M4DXFpHUzwAKEDfrhv9shwZ9EnXlWygp0T8Y5s
zM0Q2kuMA+/qEGzpBUEF3ljuSZARtgv/oXYqFA0Fzvt9xT2lUuTd+RzZ08V9AwW8
J4Ddjct0BfHkWN0JSSkL2z/zr1cracq4Epsyr0p3mhORh3UHOOcnR5eQ6XolKry7
uqlGraX2De4pq7acofSI/iIJB2fT2JQLAdsAB3/9QPZex7um6RaT5jbcV88B2WDA
hntEFsREHpluNXRUBZ/PQfTWP8Yvq5/WbwpoFCtVidxdaDDbgYv6kQehN9E4J0hU
uExokKi4sYMp++uAIXa/cC9t3452cEWGBTZH87lmexQpWBWTafoK1k8+qrQGL4o6
mnEoSSx5AVJP9v4gmt4KZhdXrD3wovryzSQyJGSV+FXtSG/zJS4Ls8lz7E1SXrMS
2DvfGnphA7aAfF555EOVmLHR8rn45TvhW62w/M98YIMVXnmd5DeZaJCncNvIuQjF
9l4dnJpJIYo1A3w+Ta4EYrm1MtAJamvhX+6esWYqneDdrpNwWDbUt69tj5yixx2U
1wHljLTboK824pNM1ljZY89bK3ApWnMMd2vr3EKvu7wHyX6vlL8smlDjMcbLVK4E
7nNNYf6clqz1gIiaLmLI29jCES8J9C57vawHTBYxGJezG9xCtmN6OofVg3wJnnCR
NGBLwMQnx+OKNe1K0v4pCamvN9rN6prLfP6G67cjNFjtw9GEqKmo9Q9XqEWXqMmO
HTfZuLFU0DWAkDy6cqmHENBV/9Xn6Afo2FMfY6pxR8P1hD8vQ8R4fWGPv6Rg3wPr
IQsQWsrL90up3hbuaWd2mRC5ohaqE2WtxWRP06e/Kwh3rWUpuD7fKlC3F9EuNt59
H4NnH8pOxIxS/cVtOGhO7XTg91bHNaSPNggfX5nzdY+j0vbtVVpqxEY8+lZYDBxu
aZnxC7emtYY0gzsWPsfPTgVOgCvYe9cbUWIHDOQn+5jfHS32p9ltCRrEza5KHFcn
T3UZgk+mtM2A2nWsfcowAgpcz7nHA0iTIJqj7HifEfABfXKzM84itlcv0lrfeLf7
v+8fcG3FQXVUb3Ok+Tgz1Iu4k4zGnCfR4gLd89mknoqnmW+I1oQVr/TJEm6YuJ+x
oAtgSzRHQvbwg74uT5JOd7Lhk58fcG+IDMNB6aQeXfUWKKZhfqLtaIFl8f1G1AXi
iWJ8eZ7rIncug4GsMiwu24eir1D848V25j6Z0e0cumlce62nyQ8b7CJoOBoZLjbg
Br1Nx+Lc3RBExNd8NhtOT9hlBUylxdF4WRpi7Q16UdHP0UnNF7ZyYFncJxDbUqOq
BwS/Lt124/b2vbi1qcJtBJYQMILrzgs8r5puv7F5FZNa6bEVcxzCJogbzmz0sC2/
860MJYLXN50huEOk0tkpVM+rycipPU2nFYWN6utqd7vCwABM/DLDpNgTpzFM81Qy
Dd0VdNN5X6K5wchu8UK3Tqu9p0CcTEWpxEBQzezBfbkZVtz0v+cBTmzzIXKruzxl
BVhAwX1Cp55791rKKlkBEUoVNkcpkXRcaa2ZLmVz0L5dnKP+Ve/t/KB17AZAQQvE
lu+yOygLdcxNjBa7dvyXOMAslcAQu/ILw+ul89m7fqEU2R2qPLHumDIQoY9PLuL8
Ya6rFAUwADqxWREgF2o7NWhZA+Iz6r5596ywxqVZYHjI2gIHt+8KN++2DR+yckPH
0dlED2vulMueq9tck0Gthyd9FKd+OVDr0T/IFkowNPDmhtmEcL19Uxdrdj4FzoCk
QB+nMEW2ERudCvgTkdDE/xyRJTXhMey40rzSRAxlcl6XesPYwSynMyjZ8d0TJ7Lx
0myhlgdHEtAzCE4Vmd5/YxrFz8tY/jxZ82ebRKQUsWGhidJaw0z7CxtS1kJFb0Kr
7qGbtdb04K1bxv7t4hdElS4OaGImQNfivTzZH/RNl8MXwxxSn4/6i3MapkkNUYMx
Z2sFn92O6cwmC4tj/8Rbp3FiNEF94zyvVfqZGGsILaPpLc05dhen0YEsrVqD9YpQ
MWXvXDMRrLOAV6C51qdMcfoXt59Gbj6c1YLJ7IkszkizP1dflcj9Ep1W/nrChsPO
7DVb8pZzml/sBUKjE8yZhUcavMMaZIWdPWfCXJmBxsB3xZQc7pv/SxT/60a7aXbS
NF5R7MM87mVVTahXJYMud6nfG2Pbplhzugo6nxtObtyJXbdMj4cZFjPKc0vLeLJx
bd/ZjiYRD+84oLZLVP62OpmFgJxrJCjukk5v7sKFB/ckLubWK5DCKluctdFERJ7q
IDIPf0hubgvRudcvO7WpJEOiHMdrOiYK10rhWIWeM2uHZlRSHT4EoNcPTRE1O3yx
/SxR+1VDD9fFliLz1OLKqnxM+sS49VhKFVEm+tPYHsc2EizZ5KIWlE/j2B/jWMsA
qKGpLAuVCmXzGIhnOvseUN6Aw7MY7BS5tfu1BYQb1umvvXoJPEWe4xWccgIx15Z/
E+u2fXbIhdVmxeiVIsW1rwdz+Y+hcPydmYIsuYxzwdXeFUXQAqMlkwUjQLwolAEM
T8N0JS3Esncvf5E7gwbiYyLybsUw4flSBGtx1A9fxXm77R1+sn+pPosoumc3OHmq
vlEo6Ak2Bdoq9Mq23PEl639QyVlC2ezViRIKt1nfZPMvg0CjoT7UwUTtziHnNAtQ
cHfv+HbCFRqzUhage0nntn9WwTWwP2Ze1rG/4RsDpkh3ZLdDFo51eKzCFgv5l/Cs
+cnGsdf319C6lEaRvTQnoMHsevGfZJo8jONeGFXxDTE8Aw3OEJS805P58sERMuEK
sqzn3ZgKTdL92p7rlTaCe+QU5ctwGagnyRxheGl012BnNg+eAMxCmdA0D0PyB8XW
Pu77DxcrJ9pi1x3swnMQPiSZmhLdxNpGjd1XUG0IwlVBUoGicQvjDxHKzPtbg66O
qQEbRsKMjkhfY8pIxeTLVkSKtqEwiEVEDE4I7h1dZDzZiAH098TumILzNtu5GWI5
bhYQ7bd3YbavqAE1ICCg+1tBpgvM29u/4iI8D0j0LHaf/Lz/D69h3UxzrCUoLtOl
+5wqZ2FhGVRz3oemdIo68z5jiDe0fC44jCj0JLGWsyY3ksHJm0OPMY+7xuLf0dlt
Q9yK+7nMy0vJM6NQDY+OEYGqld2itTvKAlkaFnwmGU56Hx633WTmvE7mR72A22KM
M3KXzpQR/FtPEIBu4NAWnT1zLH8Agz+rS5iupNm5J3xoe4FsndUd5FYVBdBbR7RR
WjlGOXcDit5+cIK6AtKBLJ8lOyyOTYGQG6LCJUiVfO5ZO9vAvR+h4Jw0ghLFhrfB
QE98YNJfSjrAofzQ43ZU4TeRO7uL05kFvsw14RdRpPk29wWRz3rYpncdEuUdA9qw
VwwgJsFD9i4Wa5aF99JeT5ieKKHQIix6oHsYI7hDgIUtGIGjP+puGOoc8lwk/7Ye
0htmxNPon/90nDZejpUubJtUQDs2ON7UWO2kkXN97YgkDsbywQBdIeaKBu1VEqh6
XM+14q6UJtJB38XYVRS0uGJxOpRQY0CvRZWQbTx5PCNV83523fkMCzUg78rR2bt+
yA+3m/hEI5cAGvO4VN1FF2X4XosJo9Pll+PHmCWXrIn30D7LK4cW34STcTk4MJJr
1SuIF0huO7FT6r0C0ZPKuei1jkiFPdJSW7l81ap+ThbbMJxspOpwLoXNZoIHojxo
M0O0JCY9EqbdSsrmh8T7sTOk6a3YXmNKSb5MSu9DU5rPYrkpOcfwQ5jcyodDsJ5K
IYz+JHW2ZZxWEpn2OhOo4xNQoHk+1O8EJHDkUkX476mHVXe+2kAZNbp/2dDXOL7B
KsywQrs/EDoGMA3W0t8x79yTNXGrxbLEaO8j/iQMqSZi+Gthi//h39FM0lZB83mm
sKzXfR1GiY+6MOZIRBjP83MZkMNwnGgJgPNhRsc6TR/bN2b+ZQzm+DhOg6FAYASR
IpuwE2V0A0c7uK7js3mADvmeTMgFmzBl9tMzjEUyp1wCiP0ScKK5VD9bggoBycsU
RnG01iTWhpT+EUAcPtc4Nuf4Txqk5oosKzI5xbLDuwrZZwSm5bAlbmZrWBEb/Rqv
nnHwqW1/SQh8pUvn+qb+F6x+YJnd7p+xcWbB8v8X3u03av++xArjdgKdvnz9Uq2s
6x9CtnO7G0uKTuWbfH8YckKHHTQrIlNJW3GSUYI7I2GozTMTvGzKg9xCo6oZCopM
8eT8S74I1I5OvBb/m0e8CKp4xshiMnE0q3ek4d5fC+BTgKPiCxyxOuKBYN93sGPj
BtqkpKfqAB7v+ti4RgIa7iJrSWaCLPvSEYE4a7Pl6uQ0ICTSMurCLal5XFyIIh20
KcbY+JcDsWawnLL8IttWXfXpSU9MzvUxIBj5emIJwuNfN7gynGXC6sDa7F9/YWY2
At+GtYfrnR2Q3L4IR7NB3VgEXPdNX25+KDtnMaUK3M69GKYdn0GitIu1yEmcsktu
YLiAjtnR+bQadZhNOmnZpb2V52CpLbfbz87/ZCQTXv18YdaY9qfKZzabYTZCbppf
oHevOwTMMXYxLcJ7JbaVYShs6muK13WTeM4Hn9jFO+syeSneNLuvNLBRZX2FkEQH
VVj7P/ZkS8xln7tqG5V18v/cvIcRcdjQbWTPthxJ8QwRReOWbf4/PeN5AXolnjay
yQRyndM5mkgz4g43a9oIz6k1O6ppUxEhcnT/dqKvFn0MyuYGcFsXMWzan7Eh0pKk
QIpzZwvFSkeEq5g7LPG2UinDwhEiaum/G+fKB7Qob2REGD2ljd+lYZivEiRJ0BSZ
B9MEWz7pejhUWPH1zsgoAhTgENcGoEwhJAqpTrtW5F71dsauLsYgS0qzFRsh8s6l
0j58sMzQTNXt7m4E8sUGAfckceoR8PYjiAMXnKce2zUeztdEKXWxYsr+ZB/24zbH
kRenHHO10UPMXf6uXGG7ZU6NYYN7b9lPQAzFeeVx0vRzElEf873/qxFmUQGVz8Br
hJxYBTpyq2zgj49lurdQ/d20umzytVV2yXEd5JVeQ7HmKOkRJcaO8wnz/48kUQES
G3gVQCNIkqgrjTkNTY7h9TvBJL1/NgEwesZ4rOx+6aDnhAIKndenJI0tixG4LQ/u
1HP9yNHR0KEMBjUAapqYukjOEtysFmnezmNnrEdq1vZ/41xee/apdTJE6Kr2swWE
GKuBWCVrTtTTBDYKDLxj3adoeSkJ/fPzVpZGxSNmWor63ON0J4NKytctmdcTOn33
GkwIqt4nbr/dULiFBeeablHw3R5RKUXRb5n1dFqcSvj+rcQB1UapOSv0ebNZxZvk
lSbgMBF2vI87/fGInaUvT9xsD4c53rKyKdgln/ZMJ6ytwfAIo6R/Phlmi/UEZ7j2
njaNiTD4VYOYP4bQe7QYbkAryFbrmOW0sb/aQsmpuAUPbxwwScOb8XDG6aH5ekS0
DhFzKjYD2r0S8famHxx30uLtI3exlZPn8hWK168hKaRJ+21v96jkE097dlYHqk83
E/LCfa660+Z1KUVQaONeKHDRlbOl/bPL2WeIAauZZ+4J5459UMu9kmrQugX5+XZ5
pCJtEcUayvjz1IzZt5ptgnGKXYl7m3UPx12h+gENilsAcstKIva4tTMaGGCCjCWi
lrPLM3ixa+iqPUQRNpq30YPPEZvtmcahCjMyU3S22gDhb1RUaMY9uF+HPgyLtMSc
kxAajk+kOhaTJzFWNurVATkVPw/IMQ08dCtdX6z2BKYkrqkZxgdMxwVZvofP1FtJ
gY9gMb54XxAjpm1kg0Y+vmjtIuGXNyvEp5Z/9pb59+DnU+abR4GzdzZGWn1ABJ1s
LG4WCxW1PIgoYKJgEXqwVGx6mbg8XuFFzmH4LoTI8CrMuPVC2VlLRAV/a+c0XUaB
GrkG240vV4pAj5yN+JgCS0ScPhtzbzir58DfmarFICYbG4SzuwY9g0ISFJRw9ys5
dzXtS9NjlY/8tGhSC8IvjT1/MrY3cNA6n/avq0MgS3EDU+H76drsczpUDOE80IBy
6ZCh9Ho+YwqklU9Qzfcd1J6i/GvfoTS60383vCRlUApncRPw9/efiTqcpQ9PsCXX
uDQIkGNC1gYoERwUaVP66NNeeXazHDa/TNDS3BSWS4oBPDGOjy4Xq4Uj1LJQcdmW
8kud9036XKqKRsy+a0d925xHxjk8K/+a39mW2ZrhAujkj3O7Yy8O694gKZThc2gK
nIsXtJvMWK2YdEkvRRqxEnGwQ/38vX7DeU/m7vvfw3K7D/tJ5MQz/v/8H7jMponj
UHccqleh8PjqsTQkCSmfRqQyEXPT9KCFkOKfSdhRN0oN2tlucXjfHhYDp3+z2qVk
vHAWou4/vpDlppuejKcOypKVKC2UgqUBdbJtrH1pIwitWHmnBOiiukscpU4a7w4T
acr+UNTMyCzGGg0/p9SEnbDRketl/K91OoDlIuA3Fkd+ngzQNL1jr7Qd5FrnDWNg
0FQZsJDoVqIKOq+lHclxso0ICwi0cr7Uge1AoseTEzUucg0+iEtJXGdoz6NDn4D/
viNhITWCS0P+wmM1Q/6n6EEV7dhHNfKISsE39IKkuup+NwARMbmaq8xPqDPNxuko
YTcyYmNMUT55Rt+AR2BvYXeOcqx0DzeIHRT8xCCy3JfAfDLOxOaKlBMbJwWI1pVw
L/2dwjv9HHXfKVWP8vzvHWvDREhgj+CENwFdow4xc0wXCZvE6UF9yQVbfUPfSWf/
yCH6tmg0snKnxrGhC7SlGycoLGEE2xZ8BUDamrC/dv6xEIj7nIw2etHoStkV3jl+
faroflFqBDyaxXttjQJ4uEQWhBzNaqDLal6/81xdfl5ZfIxkGFQC6gYAnKTQ6WM4
7Ycg2JjpBuSrl3wEapkaTlyhsrfYXovBP9dw9CfXm4b7XGpSM3gN1Z3PITQnyQe3
q0f5AFuGdxrsEKXK9YlthjMJ656RibDnUjytT+lniRCAvsjNIbg2V5eOXNqkBFRy
Ydwi4QzW79pr/4KTQqU6fpR6i6b9luA78xgC79IGt/g5L2KkLo4DnOkWSwZEcaSt
DP26MkGdJbo/FcVDpPzbg8d7DrPl6eNfW3jASLtROJd1VR/7BMW8l2B61ZWK2Y+Z
54eHa9ZRftV7jUkLbflAcVezhOiAuZvNXb1okFMakymTunWb9wuSHx22HHX4jFkc
q1zKEtnm7AR51dmbn6VU3M748G0vidtS0Od9gXjjwNtqgQONdoBEE8o5yIYUQUpx
E6Vj9h96kI63o7zqJQuLsvKT7YclI+h+a9Db59e3JagOAKN38F0MVtsSBMNjakgW
vkhGuBjLEASYxzzSVi9iNPSq+/DDvu5c6ZeYa3ZmQzqcyX6CP2sun8FNLlgu/ISs
uq8Ic52NDmNLj4+XP3/aLUOjzW8qkY1n/r91Apcec1Epd4b1tDHXsJzCcqliBX9D
sZcVJH93/KKmUifhwGdXMj5o0R9CKs+JASeYnKN6qDl2WEL5XMxEeA74dE4ukcVR
o0/rjhm63K9uVE+Lw2NJ2onZlOxlTUGHbPzJOXvQzoWzpIw3pxwzjZp7AK4UAwxV
ovYDyMzS3UsbjQUtj5aCeKN3YVZOHs9qeub9H3Utinh0OjTPnOfJzgFm8NkfipNg
GC/33MVeYtjDCz8wVIMZ90YjjGtq3vTqEx+iKt1RsuxmDmuVovuwgA8De7KdM4TB
XGCUO9CuTnmHOajIsFkzwj/ufwyF2OfGKQZ/NKDcJfYGtj1qEGU4BWOFbPovuqtu
xBgDAujNdIpC1re4+Obc6AV6RSNYuJZduZ9hDPvAc/i1qt0BF2QuUJS2RJ620BjZ
KKwq0sXNhohPPOO6o5hnTaX/O4Ux5RWL5jk6L80USFAlI6Jp5ygckcEfBDa3/dsC
c7lNK6JifCAfBISk/5OcgbnDPeNgj8EGRHo+eJqHUvcPxUGXHntOr4oLKbQeZ3e7
QD/QUkVekuX5lg1jJxMyBOAmPXDmogxlZJzC1pbdOYvWcusty9u+GYBok2zaVhei
40J0wTgxN100YZ1VZHeD9SHMkHhqpWDp287uLZqSN423BzmgJhSCDFtTP1kzwknT
euHLD+ooJpGQJj1WDGkzUA5i3JIOBdwUOC6SbYikDCVKFb/kOW7/lSpKaJCqrauv
Cu57cbjP3Lt6yx/z0jJEgFQRP4x6WaXqK2GGW/ragoHQTxNPu5TD/jQTYt8p6447
XTRiJMUDZENpRuFUU4XPmJ++6F9HUASzPWHDekY6QftD2TmbQHHB6VxGz9QJSjpI
VuglNFh9nwNPMpkQjYgBbXmB/yFBg9T/mXyf8ahzK5vN2hIC7GNHARS9xCWgobB2
f8X9KAouBlp3Q+EhsBzjBC7/cGZ1e2BcAoTQAPjaQ1XS4EqYRx6MESl5yWb/RdOz
dV38z333GTOp+iayRJdFvs5If7Wd6LmkYOUqTI6scLp5J+k99diBGCMV8EI2AL5M
BaRGHSmCG8JHXtI25oZHfkWujTVw6pQyGuvpBAqZUBGfswxGgGTAJbaw8xQzmuD1
Z6AFGQeG4q/oAqYjLVBJ9yE6MkM5ZorqJ2lFRwqsJ9Zxu6WLZS6sC1DSx1JJw4O1
3EDq7Ig+vqf3MYM8yL1nX2YkYs7s75kAxbPERxsg3kyLhdjNwEjTrBF6HkvGHcAS
8mV1IDGB0gUKx72d/5Qotnl4s80NtvpjXsf9FRNUs+vZqluxr3rNrhmlr9tkUPlt
qpWqz3rFy7k4XXIaiHAQvwjsKo8ZqaaCWL3qdjP5Vb9s7XCelNJ5eoXwL9cHGWd8
Dz6bqQF2LLqQPtrjbbwMxd4EpnguH3G38o2q++AoRp1c1hdBPjeaRFI95SQAMfWz
1Kw5qRcIOh+lEDg94ExL2qQoE8npst1ZyPpVxIRv6CIjPafEQGuI1G9W7+yhrJZ2
eu2Oir6rUJmPhVt2QtrOMjVIUX+6djrmz1pP21whbWXKM/6NOOf2Q2qTabJB0/AA
Ff4HOcsbUhE8iX/NvZg3hAZIqbk/5fpSFyqM3CCAuwaEAEqRwE1V2foXExByVIaP
oj5GRsSZB0uS+nDPbxzz2YlkI5++1G9of6/aVMwk4m5RWvFEHZNp9B+G+5nVOjFF
zniR+DoGuKmZzn0wzrZSKL4IXSjZ9pYcwqp9PULmJOh7QnssE33snHzhshmHO0ux
BuWUFzlNaPajFGdsazRWinFyFAyy//WanMU+v3Yft6aiXgAAGa1cHX+XMzKbLQbf
7SYB7wuPwH4lWReqagC04AO1j/wryx6n03ehjQWQZ7JdhzvzaRYPaft39d6YpCTD
P6ANOQHi3CA4zqB4wCW89KDLnQGD8eacyutkIgtE3ZI0GY9Z2cskoPnkeqwfwM2I
e+TOGWzTpG1GgimOr/Mp6PE2g8S5S6728i7y3poNaDQuqY/xXKFPnT7bmvz7+dAq
pJfgkQS7Ns55630oivvAwzS0Odx2pXJLCNCUhIwoUVb2Lpxyn0gVFYVQX9Qt0dNt
3XuFRHCAbD+oxeRUxREElza+LThX47nRJV7QBj5qjqSJcF7U03oXg6Q7sYIeVJYA
NT+A1/wfZYCT2YOHvmm3zL6U4wzPnCuduSg8AP3rfDq/71VRkpmumAHiHuO+efhB
o6U9tHXAYzo2WZ0ani01lK745rDjYSwxhzzLSp54SvSBLAo2aLzuS4h2ZPwNIuwR
Dr4E5xLz84RItvJi7Pt1Se2FQFwfXN6Z5P+xqycIG5RAJ9W7GiZyi+410d96NdRr
vDnhnu6k2R+8fMh6F08faIQOBILOUQyLwKOgusIPg18emarorWwnHTDjxF151528
vNYgF/5GEdEivmjxmoTQ8r8HPpCL23wxBePPoGE3pjWjShlb0nbGmE0GOarWh2Ga
h+l9fzureIJyZbPeZh8jWMO7HLmSaDTBHqmOiNQd5/hFDf5FE4xUVb66bJrnRcNV
fPTo2cDOwLUn7Bz8PEosgBtWZ116rhntyAVp2c0GvHFqSTWHcjFcwC+8yllKv0Lp
yB2f80VnhfQ8HsncT0XDc5DQj7lBMQgKhry3EjYtTnPP7Q5PK97o3LCwR5syWoit
c2Gv+E48tDb6blH036a1dqWV9gwcYWGrLjhqM1lRUaPcpakE5BHzJ26v8mrEc73x
70xndCOFmSoe4YfGGgDpc0L2yge/H97UGqvg6fjdtAuJQMlK7ATenxi6Hx8gFiF0
cH2lWzcLOwi/N3R/B03Nu/sUXUrHIrlWZrSXB392f/GMU9OvrCy6WnzW2qicdA5p
nDLLtF6n1fUEc0ugEl8gBd1fOMV1vxAsegkL/gy1haQXUGVzthHq6H0ksjuwDnuT
n/JCHoBA9hwZMoChYNJiSwwVn5m0ISpALbLmdtw0rqKyskcEoRPG8Zngxw5Ihq00
L0KUvWAekLabAcCJovEPHw==
--pragma protect end_data_block
--pragma protect digest_block
67cEY6+H5xAkqjJ4ZclPPpNn0gs=
--pragma protect end_digest_block
--pragma protect end_protected
