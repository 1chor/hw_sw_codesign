-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
3Tv5qEQPmA+Mf00MUBWvrHByt5otxVJULbHGcBgC/itnA0NhqBQSjZHnJtOIEapZ
tgM8wEtMOVdN8KXYiQHBi4ZR697+BohogwiWEIIx4qczzgZ5F6iS7k5Nd0myVRFB
dMlYYlHNU8AlV9zvJODLUEgC2I+HDeJ5dwcdp86s63spq4RsoszBmQ==
--pragma protect end_key_block
--pragma protect digest_block
iojn/REikJIPHUxImn2IWQGwMGQ=
--pragma protect end_digest_block
--pragma protect data_block
EbbzFUoimmnuFUIb5K+bCoFxJM3Cb5bKtSh367S9K0nr7gBV/W/2tWZrUgnSEZZ+
Cqq3bkpHV1zHWAR7Vj4/xMfkwJ3OGt6Sewmo7kZBkSdnYUoHiqymPrq1bFBQfsd/
IDVope+dDzeRfzEZOcAgbuqTatlduK6kLIghpWWd93rsfB6Oyw3EHNw27wi9pi+F
I/AnYXd09T9EHhwVhOA87rMgZJLpW7cAsC2R7zDvVrwqD9F6lmvFBLJJDqjrkKVW
/YHmZrM72+YT4TbHhBw1TwhpZbd79kOiJoAO09yDOgC09cCnFemiJwpDQXU4/ZgG
fzT/ziCPoJ6BjHz/20kDO1kyapADfR3gfhM+96PEGTPueFEGiyDwEKDPU9XvsBwe
gFRk0vLWD5ljDSz+I0soWHFtml4tVgtLnEdHtMwciGGUsuWZX6I45NJVRfyauEeu
7it53z9sHagh/krVXr3yh1i+6EK4unahL2cXRwm94bkr9B1bXliZgp6AXy2ErJuX
p1Mcx0bEAc/dht9DZVKbMZsTGtpplezmEy84K7KOAb3+Nrb1gIqerkHr7DgtRTx1
TKBY1DGahmoKTjNAIgTrWkDg1QHBL7vgd+ucLz5uRTiIJUEGjsHQ1b29XAH9rPEV
kHSrxuAgmZKl9PqbS7O+qFEgndjK34xcqZR/49HMJMPmsCYs50lxHDA8Qo+zCGKj
sa+bcZvKI6ub1dlIf7HE5Ar+SrWc8zT1xoxEA9tfuJKrwaui23k5RVCYa+Xi+mBu
LmwJwIffRKAlnkRdeCUYIm689cxXwLVEXdbzFXkaNp6Zfcr81X9SMTSG8KJuCBbc
+Z59OwMH1SJq/QC422Mh3PE5iP8Kr3frB/GdzcCzxnSMjo1RoXhdaZZTQrznB995
EVNooWZeu7zxjPVsUN8npNK0Tb9VWuY6jB2q98iaxy1/uRNTspVOKtpwH0oLAgNR
uWwKPE1MJlJNLXk6thdPFfGPsVaBl/ZdCV4SuzXNHN5TaJTy/07QW0xDiZKHfXbn
zbPNSwMhz+tH0xVsxLbY6Nz1txPeGhH3he9B20HSsMVmo9qWPblFYWqZmEOZRuS/
aSKPZZ0VMwiM9RwzrvFR6OW7fEUY9h9TI/PnSbE8ZNdDgapzhDv+96KF1u11HxA9
33084GR1vPfQH6c6htIM6F2MtJtBrJl/SWRZ9NpH9zNh22mDXauPMtZcRLlpVhMn
82MjpSLd8uxCY4BWHmrDtqcP4h3NyECQqPfme0S6gWLZp5qrp0oPYlp4eQ3uerLE
NLvjdi50YgoAQETp4lBzPNrUhOnXyZNb5ykxIl8I1cTUzwxYzoyEid9QVcHeq9uL
ieeNClNM/MOuj4HqbEivPVvy/VpTlUBGL9oL15FYs39st0DiL3BZfBERj65mrmsP
kEpOzPd3cMhyq6GwNu8qJ4bhqw1yq8OLSIO3go5Q02J+zAbp4gpUH2DcbapFEMh9
G/vsUfnSRkJKF2KyUj/1j+j09JcVHKZO2jk+mc9XSdDN+mFbS2k7ZN4Q0POKEnO3
J3N3JfGTpAD9pxBYZzf9vXdIwQrH/G5aqc/KDi28MIYwUR8DElShd66YPN107yNG
84cK+coCBZjBFn24VJFsKsLzSIAFPktoiAIC3eCldJbDrbCUOuGPcPk54tuS2oY2
xsDmqxYagdbqwlCLiQ1C9Pyoylqa1yEytw1d7N8zv8lbKaPsLQ/eLwfvYFoOiBI9
f9iOfvfsCYW134eLBTb1oqfThQJGKpofNYKeUPi2gsi4wodkVp8YhKB7NLpCmlLK
a8aXgQj7XbMOl2BHFt9C49ls2JQQh7R2knUJLAKxtxH2BHvaEzF7E1cpqG/fo6k2
eDM8YCXhndZml4/C/X5Arsyl47oN0FIzI8qVBCqBSZSoHmRv6QHshX79qB4G12Er
pr2S5eG+2HFpqBfhGx3xhPVmM6hfVH80BGzWymJLHnyxKHi0g+1Lz9HgUvVh0wlC
SuyWCkGh+hDkwZYCxpuVMfIt4lurv7RPYJSJ+ThVtEFZZqlqYUg/bO0wqwDA0LIw
6Gs8Qdlgss//X2y5vL7Eu5L7UjOjxy4Yyyaq5jBslneyU7vRuDNOZFdz1lrGShWy
YoOJGN3/Qd7n6qdTEVx7tul/zk3y9b5nE4h9PnkDpLyxcZM9QPsavQkiAMgoceHK
5talPyXDHjgQL3LVJTtk++/8w4Hsu1TC0kKJSqiwfAgOAuoZuWl4k2zMcTEaRIsW
eaxzS2yxoE3pZTyQdtuKfDUkoceKnFTHrx9R7emMSmoCBcZ45wuMG2/zd5ljbtPh
AwLnkNx38Czo4W3lJA1WRuSI80LQwoo79I7rs9ngX74UX0JPSi4Jih4lk4BwZSX8
j1KjrRUD5eTk+AWZcw4qRoucH47b03M/v9Wmmzc93Hh/99Vuzouy57gQ+th4Ov0M
B6lpEIZkdW8WLu21rTmL3C1KzM6xstiDlS3x6wOiQMS0HuK5/dcweFZKuPjMAb/5
2hYDmmdaVwJPfXDFGgCuxWXA5/RFScdlah9jT8P3MOVGsk43DQIqrTghj7+3do7V
5/+mqEhd+9x5VZDP5XOlwsXKznkzXwX6hKMaMtp5nIPMOLGTX8J01vrAlQ4AVaXz
uGGbx+YDbPK64pnzPKInLLPDPgPTujKQjcVSAFFbjrUkhIlsB9RT96FALfiUCyMv
tSA8TIMKJWrsFI6vAvAAnBWi3SGIfS3ApGXEiwk+oy6HTLWL3Am3lwgsCvtfjLal
+baV8lS3Lxy61ubn6hHnq+zUOtrcL7AmS4bMhaFlpWJbfZJsXXn9k5PxJCtGPxne
ZXtX5sEI57Y1SeFOhFwJF9xIQ9YsmD4+0bTD8ifX72uloLskRyPoIdDX2jdlCBfm
ovRGQLV/aan1rAm/rmLQasvR683j3vSrU0nwE5qHlzrBvEEytxzkhvi3Va25jxYC
6HCZIZlT03tFxCojppqi5UtpmoJZ5yqswZPY5nzfkQrmZU6sQbvwae5CGqj+9r1m
SW7ImitPfEBbG5Jp3DGDgE0s+4IjfJrIsDBqMqSiVcK7ticLP9ezWKV7RPD49kYz
GyALu5h9TLbAtGUPCU2K1cuAM+Nt4BuiXf0ULB22IMDL9p1iwz6sn33s6zKoMgcG
DoOjeHHSHbyoA/Fjr9zZI5VoUquLNcx4WgDlDGJyxI61Fcs8ikYfLZQPjmsXASD6
NLZjQImbZmO6b6Q4HjYCUr1sRGKvR50UPBXihSLyOcOmRqmgf7DHIEX1iLnlk4qm
9dElvXoMMUAYeO7YklgvQlkH5CfXU6eAUouBpvWz4dvvwmkYmTWzEPpJj9+nkyz8
X9T/acIxVCXIgmP+Rhym+7f2kBQ58rpMCVxKvEmsMfFAkucXZarX0HtBx5uT1xi2
mj8ag2xnnBnKyTZ4y9olRc7bqBCsvSGFgLV3+e1xUqud14YOtJwIFMIwhscxO5OL
pW/Pt91S6a+5zNN2s4QwHLW1efHYQv/M3rEqpcxYaraLMZU1WKmUCfo1ymRJ0ymi
fYC51VxvcXEDLHxDUVR+RS7IiNffVpkyoFfy3c7/mCagTaxLyc5CyESSekxnFkZm
uNAtIxts6GldpjxZMRHqz77G+hjcAnd9y4Uz23jNRNdflcTRBGHZ6ENlGWZDYUpa
sMEZDxstcGFCzJYCSfPT317e8EEng6t2K3UBUaz0zRuXs8Ju9VeR//Yw6dfARVxx
jV+wGRvXzLbOBZ69zMdUsjN+1d7TylCLuopmd74jHmasE4uzA2bFErNZEaK9eF1E
GmPu68h3mrSRcfVPJ0VvUcJg8zFo4kqnrsQx61n8T2X3XUwH5CPeo5ANw2/b1eaO
DYNUzvSD4qHYT7PNAKz7kEa7AU/rJUvmYK9Pr5qPF5qYKpDt3luIKapjl2SwKbNh
PVx0EoBKIAtby9JrGnoCyzXIplc1Gg4NHAfo+KG/43xrp0vw1n6synp2Fxj1wEVP
WUFMk3clT+h2XybBoHLM79BmutfU/obvA/Yw5aHVAym32ZUC/WF4OrmnkoyXGsNe
T4cl931mZjW9IRTqUxkn9lU5m8SCQ4omuq30lh5zJEsVhK0V4WX5X+hhjR+wUsHY
6c7NX6egLXGA7kUEaee7vrhAMtyq1r/aC9G3j1SLEH4rZpWwflcujhcXcs8cb3um
jaedvAnH//5RLf8IeQFLR7VH9wuivPFnFSE3YHxfenZ8t3yLsLWZNH9J/Szs/Rm2
qwe4clA7ahYt1zNRyERIc/LGUudFhDf3MZI0Kp5DBnZZ2eRHe9OKLzo07QbrG9x2
2k6z3o22ipgjDPcoq8wB1JSOBFMg0EOo+byo+v77coPp7GLrYNuq8XdawMj6/xZj
u+A52cz2IuwFRxha4v2rsqqRIBSwUaWR3oZoY0W2tUypoJDVSIPIBsedq7jZtzEq
zAnE1hyXiz7ljy2GV2fQKqs2XBLGbt3MA+yTNj6K1hu9vMG7aBPf9E5Sm8U6/fC0
poqL6NTSSD9iMfK604y1XbrVKAQIJjvFNGNegkCxqUeZ1B2cLookbtG/33ix+zQ8
1+tfTY46wMvtZd22KyPhjYofGaRrkaEfr44zzeAeNTZXFZCHO/mXZPLJlAqGSUcQ
SLTvOZ/Z1pkbtSiJUa86M7vy+gx0ftV31x9a36HIEePVUW220RNCyqEfyrv7eT59
wUebusLbI+KSXevyTUFYHohUWIQK8X1YhLEF14VPiORoPITv/akjmTDRf6G4uXcA
OB0gU2Xyd14NU2Oo2gIwlcyyKTGnia4QWc94JkMFmgoelnr2iLUUGXeJnSDvNcBa
NXbFyO9ez5wo5fYMUL7zEw27HCBS/UXFxvfKJckTLj+rr9mNbEFU7N6RC15DOEck
n8Wr6iddSTYjRmkW0UjClZoG9qdO0xTxEGzaGsbSRSpWAKqVbFyaoV+COMINZzHN
4WuD+k0dNFIrKA5aO7KaV/bBBgtIFYQ3daMWai18nw9EhE6bqkqfI23UzOoJp1hC
xdHe+L4RhDp/3pyyZ/eL/X9HDkQThwOXhvlfwz3QvTVqXHHUce3f9pHjKzRnxGJm
MDwaawZlRcSPfwWQnAXRpvI2nQtEGzx1gUH6swj+JepwcDE8UQeo9KPsJJJqTWsg
bx1TGX1BRZuP/r4M4gvpoJkcdrj8LTzPuuPyKOkdBuP0QpPelOQsdl0e0QcqM6Sx
KYr7HqiIcUedifSWZb8qnXNwjMVxXZccWNuMJhSK35C57olfQd0WKzO3A0N2wPqY
SP4iw81AkqzG6Si0dAE13ywkUkrDlblkjn7Y9lq8ngymL0Jq1N/wdY8rBl42khZG
PxhzAHbGV1jvYN4V14DgG0QEsNT9dsIsoOwjiwHzIdkKQhTEKbBCkNggIHM0gilb
9KoxRihHZfdrm6EcAsmlLlp+58Fbw6NuvRcdszN7hzoJhf4yZgcKrIGj9B4CcGhi
UEiamD6i+96ZOzigbdMK5V7s42ET1QgIPAKidP44u4lWTUa9y34jFtD4/LKDTKw8
M01/Oh2YzLq4kOwxr0prlCVrkfy0zKujG7ogbbWOZfJMUAHzYfuvotQdZYiu+qRO
hIwKbCZgGuHEbaEv/hYeM/KB3ditBXZ+zwHXLzGZtxxgyegZBz+krUcV5B7RpCJU
lfCcEtPGO3ExBpV/aj+D1LilvEaQfSQ66AysUt6Bi01KpLsYSa8/cS0pIi9a6woM
bJf8ruBkqKHxpsHsAmk/Qp5MxiAuRGtWZ+cIp7lhvSPz0bI0i8I5yUxXJRHvDqa2
HjNP/XgVicfwC9nWexYmpF2mxOQJ7YEJo2vxxE6j2yHbUfqzXXFBzNCmZDnTfyHd
o/S2fVZrAcZ2KpSi5uowTNGMCXYJXzCBwc1BC0FmRPBjqm/KQgbnR2uOD35DkYv5
Iw97rVoSv0HW2g1yLgnkXH5X/w/25tgL0hoGfqdM1yjoqCS3TlpFySzkn0rJb0Yt
2Sm097HiJks+3ttAr0sW2JkvpDHMDKo1cWn94UOKt42SODZXda6LtdbCztJtneM1
aSIATWyYxapZSYEgLwgyWbOw8ishaBn/WBeMgw5KKlvzkMKbYUSQS+dHkgMC9UG8
gdQHnB2t6ToCAB+5EUslImOPofCJC/f7i5Gmufoo6gmx1DGkS/EhFmKnrXLrWiVt
5TStr5+V/3MJQgvR9z2Xhsgun0XWq6EdLooMMxZ+nfsb64vVh7TBT0fBTFLv7nAJ
jyzf0vPFPhEVwU9yyAlQ18cNmYIiccP/AwLOV/7yDDaAvhKuwXsfm1t0TnWECosv
k3j/JxhkrEJ35+p8u4BnIDISCXTR2fUFboAZbeKXNLxxujcdXBPPiowG4plXFlvS
tO9MAaA/WAggppdvEasnGubTSRNWVf6Bysx0rCYeGHW6+0mBRVtcRvSdmnRjWL7Z
stMzp17yZiCd8HFv1vKS8kmCEZCLsEuXRwyi7anj9vgC+tAQldcON2MfNHRjV+Xk
p/NBZJTlaseL+eqBQC0v39YbIpz3iDdWi8lydm4KAFt5OYFfecmfafF68WMT/Yjc
SDECCuS/9Jgq3QbYcpysVwVod7XNwYaqNBplH72nGCO6lxhCXO23EOxyDbEDy+jp
Pz4cY6tYeGOEhfkS+Ia2GjBiOg9DVFLb70n3bBZDR3mC3/H1ZbL7Ybdw0DZ6X5mK
R4ckSzl0eRtgRAbjBT/+nJ0WvkEzhs3DA5/3ZbFMBS6/zscYej5A0jEYAuO95ivS
tIRWbISo7lNqR8kz0L0JursIABwqH2lRoawXc8nZJV1ru5xQ8TocYTVKTDg9qgFn
PtSO9a7OfkuwZQiJJDlr8mFsGm9NUg3HwpQGjJOVdc277OzYPk7YYY46BbZOtGb4
xkpRlAtudcsQxMZE6ZOw4KzmVZyKGgXLpeEz8up3+kmwjKT7UqwXBntkRLvBvQPM
IUCE/Koz3iKaeMC3hahsZRJ3CrLl+D7A1tH246P9XfFpyQPOBvFKKxbiOdHwc610
ODcJ1lPPPfFytTJo3NSt1lmNdfpyTL1CIaaK9Fr5yJxX0IM92VejuB8g9u4AioML
22aI4oEu4IOLpqVtfWqW+m8Sxv2Z+XT7hCnlJJzBpK80vwz8EJRxGn26u5eq60gt
eu7xiT3qLIR6G52y2SlJEekcUs1YOvVBuDKmq8dtWml8L5JzJZX18xRMPVuP0ySE
+4cvpCjVlN8Xjhv+lznRiRvfVDjZPN/juEfR3sjxOv36eqrOFHciCh+BOOyMn2qR
cb+q2ZjLLrnOB/8glpjU3uyLyJr0NFatiPyhyEzWjOO2FPwvExzV6eQ3n9auJZW+
IP1u5O/8eNqUbpSkVIJ1OfHMh+HRCoNlW3G02rE+MuYHqtKSNQRqxGW+MPrS4rTC
QlCZKPX6H0m9kZGaV+trKS7LDGBFy2CPPL3CxaN5ho0S1fmikI2iOWyNpaeEUJSM
0N4A49PHFGSMUPNZKwjHxDMeWlxH2rlfdb5zcwc4IjnAfv9veTiSEOeP5f25/wu4
EPeRXwSku8GJCMbsJhCGkA9PH5iUrcfG3gEhqKfMQM9RMUWrDg78jLBhzCt6v2ln
cQnIA3CNDIKMmejBlfMZn5GvgdL9LbgHkMXuCk1JahdMAryvEGIcxN8nWdU6uRJ9
wJTer7uoPLYaxw2LDjvqVkewN4GBfFX1BRzUzKey6n2FWJpSr/SNgCy+2OVqEYAo
nTxniRPEGQ3fhitPpO3LrpMVg6mVWxIykA9r5Y8XxMI96oL7dqvluA3qq8bQhOn0
pAzJpuQoVYMndrrLtq7JzjXAN5qVvEuwguPEuwwwSWUAsMj97ZNco7SwoC3FlTZs
5pXzEccMCue1WqWljydJFPeeR37cX/Am2V1xuLSd3HPFU1Xp0tXX5nT7Zs5nf11b
fr7u8xVBWukX9mfJaPluWucyipCVCoV6U+eHazDm+SzfBvuJiQeTFmBPSqPk/L5q
sOuZSYi1sCIbiWn4lHnOrmHPUgM7lzPTaMOr3QRF3R0oU2+IFT+Khaf/V3nsr3Ud
d7aWnQ7HvBtiuZ9SWFm/D8gw7BSpKDfalRRoI/PrZZ8gk7bhhMMK9Mu8WjyGKxoT
R2gvHnBHh8e/8XVH4OPZKCOWEyrX4PfvZrNwvrz0c7u8z5L7Yuav0EcZAYVRj+f0
/aOvO/vVFyOu2AVgGSF/YlVvRUS7m88BFzkTlU2OBN3lwSRt8TMWMMqShD04xN4X
sWp+SkUym+5WokUOQaWzDnw3Aif8tVjE6oWG1GhYlKzTdVEqyYOIm/RWzy+XKFZL
HaPNCiCn/JUeC3YWm9hLgBng+XGE6r5n2s1wRhb4nP53EtEO2HX/19hOE55wXe6Q
i32VD09wyFO3Egtd8sIS3ckRV48U3OkJ5Z9rdVlfOx400FjlfzciVDfp8plHforf
j/4PEuuxzHSeDqgyO7LjwXEVMiyUKNCyvJB3qr3JoW6qiCKxbJbasBG95xp9U6Ap
mlPJ7e0YHwjFB/R2zJTbTwKml8cQolPbrYYjh17uhDTCQrWWttNeYvsGq8J1vpTi
8r592Qr+H1IOCaEEbLVGEW2N3uvRxh7HRD224hScYlnh6Vq4msTlnEF8OlK3VD2Z
giO+iqbZaGuCLEC+dRHPH4HNmnzpz9YnMAjG5UgHnopRDhcOVzL0wWDt2GA5N7h+
or5yRz8RnHUXXMsmPt2r1vWYubhGTwIMmlapLeoz6wCSdNs8UsAbOzrYkJZTIWAx
aRUvOemsUtDLWCYbsFdcczImiVz9S141F4vqe4x+ZqmpqBELvN5WK9TiAaDArB9h
fwFnILAyxL0KX1CnBsnN+Qdmpe8/dmanZp7oklV9lbI2xdyhIWvObrhL3BpCP/5f
X0UyK/HXryidleoGNpQQHyJV5uomSIGGBp4iOxsoh4de3zw8iFH+3oQ7cpSzKqMh
9WOUxSkb4sHCS6gw/nQR4e/zAypvfaJSr2vpWzMG+7NUvPpSd3tXOs+Eb2w5xwmE
4vRbuQFWrYN2pDh6cyOFOraMBl5rJHMGrBeg8PNDND/8l7kGEZSGb/0EUVju2bbw
Ka7p6TcvSY5HkqjkWHXKubCbAF+WD2kNsV1GOOf3VKBG2k8uraz/KPqUE/1X4Wcb
VAqOl6ZmnUK8XOx+f2yrDVh2Ho0XVolOwgBuMrWwwb+jydHacMa94gi0WkiO3W47
0WH78Wix2Y97MHhX9F22DfMqVoaZO6J7b6FykHCEQ1ozUo6UI+2znttJL6+k2RRq
UV6/PRdXLyJ1FpTN/UvNLSjxzf/AFt3WheHWpkMpulghnl/c44sj21neXv9sMg0Y
/36ArSD+A9QQ7V7IDE8A9bRdoB7/syv7LnC1TNcTbou5ZkCe2sYZzCIZqKA9BPeh
KHmbX7Xa7YPhZXW1cj5bONT5I8YhdxvUBw9iQrbfdLH7hzkYGe7sFKzxNNAYJp70
8ON6+R1wEEUUK7dBQsIw6wKlrd6wXFIwuqvtam3KFF38MTYHA1ND1NKUrDNvOFWW
PZWyrx8mcOpRrHjedjTVUyKaLlmIuNTj6/6Pw50vEEiZmL9ilq0K/SG9tNfXuhAB
7/OGt7fvvEPp204lhe0bb3POrvYFtl0DhzJ6EBqaZGxP/+/8H2e0EnOJZSUrIv1j
BrElIy3utISQzKDlVgR8PQLvnr4ZoBgosCeNGysUkW6mP0TeTWhB6iTw0z+me4/q
9P7q0vOcBaUao9x4wH53CTjhj+AR9DiPVKVf6Pk8RZbD/8OpmWnoYN55K9QkGULe
quMiUh/pP9YIH6aC7JZmHkmy9N6amld+P/Y9adcBmZ6bZmfEJBMLzBw8IgNG5Zh6
offaS/ei4otdgCBH7yU14GT40HMDOa1qaiw3/rgOgRG6Y9cgstVENmrhAYEe/9E3
c8wGfwYb9g2LForav54kOCBikIwEtPVpixe65D5fBoDR0abmlMMep29UAjbtZGov
05l559b2sb1UaRrcOc88abbgyfT9WJ4vTucmMR6Qk1CjIHu5blMpDpSPPPaKjYKE
Z5XPu9EBBZVRbv1kdB+Zsr3zuVLqAI+t7fJh1OcZnwm9s+4veIvAvNLj6A0WI1Ar
Oxn5ZiCWsnD5c8If85EvAtemfQlk2VBtFQIanmH1iLEJE8Dm5vKYPHLW7V+pjR41
e2vjj/ud6iVK5FFuKC0y6ES/aRx8eU/AD9j3MOxpg3tEdL01j+NX7kB6Gh7kUtvV
mG2BRb4HcEn7jkdipO0ZLkYGR6Mgth+puZ7HCXLgp/djtx+cbxbssgutWoTJ0fIT
T2/Kore9TRhgoS9zLfS++cJUCbQFwjq4Zq5rTZkSS2Khk3HTpoIc8huDKykTHG2G
yzJJNs9bDxrjkn9v38aALfcy4japlixJ8fgMFTvrDOgNmL5Am+326BmEMQqb3jPN
vP8sTCkVgxjFNkLMIyh2uz/nxhz8F+ZZK9MFyFYSe0QE9h589GUfAplbC4uiVI6W
/LDMxn4JqwGhZdmfKEQPRz3oa5E19GsSRvz8ghclPTFd8gJjJ9kqv6dTHxCJybJs
1grjKA20+VvjXA9M3RSHBULBhWzrPf0mc3SwkDmlH1xylPo6WqAaBb/o4flT4pfi
KnSz1FFVG65q6akcAB29fSae+fAYgCt5FnvEJBuWl3ZG5rfHpOeVt0Vd8Qi2/eLp
4Ic6CiUb5xybZarBSt6kRHs1qQ0P40PM0igsMqmWC9CxYs152PMhS7bcCywaqRRl
NGyq3959B/AsbeY7HAGdBuNK1Hb/RR973r8dABjZfQWov2pe3WqmEDXmgbQ6cxsb
tOARn/ak8XYjOK5Px4bsWF+7LWD6hZUghE+t3uHEWBlU0cK+9paePtjd84t+ru2M
YQMEe9LsLo0SBWENzxek4pxwQk9cjKSAlVVVz+6dC3O3Ax716IWHUsnxtlP+qVT2
laQFJhIAohnF7PRQmv/bJs1+E1r3xYAv1LlXieeSoN2kcZPo5YhS+pSjMvJ6Jmck
eaOS/IbkP8xFH+BwOWbxpp35IUYJCbEg77FbvaFFXHx4Wx2zfWq8rfu2/k/XHdCq
uDrQV2R/NBpBKprLiUz54yCXyAyrniFN4lGg7ENhyebFbBHsGoBgPwLKCCNMfCs+
GEwptoVhU8h8DJCU1Oz8uRGP+vgE8cHQu56N8HDVCfh0fFa7bafm+ACg6YRN7d2w
FvWeRCoYIbivCvOXBG9zsbSu+r+6w5GsHXEE+0CKs92Uzh+4ev+T6fLRv/qdl/VB
m1P2CdGZXo3tTxs53m8NzfZyoxH+yCrbB9wwbfnYktzziLCTYWT5jPplXbaZcWAl
vU7Chm9P2nxttDS4L2aFuvmhMN0M1ETisjPauyjHFqrEA1nLFwcPDzB03tpAJoWg
0sjz+Rm8nfx6zHqf1gCCE62EOlcuPkT5M9Osc9kLYcAyMw1AAyPtk7TkkaIp4pA1
UUMW8ydJUjmJUbjFBp9ZVrcSupGnKlcn5WMFaerX8v+tLveFhoQtuyIPUq0hN7ln
eGcTG6MUymdkoGcCeNXWmceGFXrAIIw6n9lnE1PR8bw4kdb5hxrTLdoY4z4GjR8E
/R1CDGpZq1yRWBXpMqbuQ/UG3i43irCH0crBwPBwmPoVW6pyOMLZPlF9BKywRQpf
8pvNBekByo1DctXJomEoxiBBQvENOqtlaWT5lsrihq5mPZuWrVm5W18lHHH9tV3N
aHBaqyQhb2LaeOMAANOfSYahqXhaipwMvMImlSiK/vHnneRkRh9SvcGAC7cKJFpN
jWMRm5HnFdV1UWFUKXxWl2MKgx+Xp/AguaD0At9IzgB/eWGrXC5xAOczIK4toY79
AYc4tVetkSh50D/0DyDrmIbXyjhyRtY2nD5rh2bODQWDuxj3BXV9Exbqv6jJv/uO
Ty4rF87ae1N0OIY+HT1MuQn6Ko97FH3G7TBFtipQgMyA82BzZ8iMBi2GDK4B+ylk
QNqbxYBgTNQ2/uWpTqOewwhwu20xkzpOWvv6r2lDZ0cci4vCmWVKbDho5TQSrba8
MdeyT93UB20L+33nY0LD/HulnFL2e1I6mteoRXe4vrUBShlJJv1vtrhnGXtP2QT2
Dlf0wanQL91CHwNE0MgtAmZGE9cXhRlIJ/PxNRurKFSDJqheT3ldaTIxCDj0Wulv
vAPLrhgI1YNprHfS2hXi0k9nK5LI1KG/ugdg9Ll23Q0vwwwzbIvM8bzn/43P3/2F
TWeCNM8zuPUWbuBxh4kncXjeShrCb/LBfQcEH1WcyqUmnYJplPRJfAOXRc7D5Aq9
sLN+rW+IxGAykNQuhOt43k/W1JLQXQs+jBv11P7ThyC+ohU5fre9+5bhYDXin68M
SHYSrSEkpiy9UWhgjlVGGgEagLPk04JelxTrHFsUX3NMw9DpKjHZuNeQW6WoqQI/
mCChMGTiSzESzhGWvDqebLaEtki3mLu1CzGg4A3+HlHfydh/9Vfixi7zOsLqCCQ4
GUPzkjW2G4KWooqrdJiNXp//FDkzb54bmSqIC+sNT4g3BfIN3tkrUHZ9mcD/nijU
gGLGR+T5ilm/5jJR2dLtqAMZ9ZMfJgWalM39PGab25lYRADFgwqvHol3mzC9i/aK
VnqJMts6QIdugqYrtvBSWrCiiwmwt4l38VJ7QN18ubxWg5YY+xr5tsX06xzBAV0y
BvpooKfJbSDHqOularA9Vv2EeiNGgg6qE7O5ZME2ZDuBQB1HLS15492qXz5Ly/sw
kX4cmRsfVZB10ZveqJHkdyh3w4NBKyIU8SE93FbUcuDzTWzOmPyrzKwR6Z1Tr+Q2
fBmPSZuzpw5PPE66QR+6X0ZniRrDQ0dk9uGePCj9HfKxihshy730I/UEX5srk0bc
WBx+07xiMxisZNfFLkcL46urqsBJqHMRjkR1st3cXtKK7fpdlkZh/VZ5ELfipq3f
huJU+bdEv04iE+pR5Gh9dUjpyaKgaxo/MpSkctPbWIB0RA/p/VuL0NGeI8Wgh3VB
bKAdfI950872QOClc70mUH05jMsKhU5lNb4bHdnf2k/kU7upKGF1GWzMq3fWtJtt
YhANAkXVvHhbKX2o7CzDDmY38Lzs/tJIJrsfLo8heFYHWeZ7wqFudn4ZATRhERDg
jXIQ1r9hwdLc8m7K+B8wEeRTvfffOESfZnQcavVRv4AAtymjFIMHcfN1hkRakZCP
ZRvToOPIWRzn+ERmif9/3JGYdWMXiqIPNhoeRxjbcoVHG8vKf1HY/WJaPB1QL43c
IhjmiS+Up/JEFHwykLx6ETr6g8pap+D795O2JTgHkAm8j1TiWSS1NrTh2QO2lxi1
ZqRA5XbrmgEWTeeQ+kWu1LvcJVtFRBErblCxpZTS1NSJw/TylPgQYP3A8CpedvDA
V6MBnQXNOljTXUQ3k6438hmIqVJ3HneTVI6HBxxTvBsdXw1MjhQNC/H5Y77uNEMN
EeYoQPe+dNv8hTH0O9JGU9zJuf//+g3wK2sfVk4GvY9Dc94FQmqdG9KcOqSHHkDd
9Idx/x5U2EDzoxZuw3whc+EGNZ8uv617dXvrES6sh7C5wCCJMSQ8uNkPMk0wfK2n
gwSurQ0rYS+sP1JibEOEh38pqN3jYC5E3lACkPA/6jTqWpDmi2S2wLvceAr3qoAB
dui0PcdJukVy5SwP2oxMZfatliAs2ftS1BkjpuPQx/TQDZTB9Vh3GtQJ3NaD6KzN
PrKU0EVwRclfACXu4dRLbMNHfMVOEFrmCpWqe76EeHRQ9X9py2U10tr2D+rsJWXk
1MhxgaZ2PWPFkVtZdTyaUi9At+y+LcTosCR3RUE23suwTsPj51zbxOdzo5bNOh67
PxK2NXumgQ0prslPPQoVrQ6cH4SCoubwjOKbM1ovZNecMQLUfcsoz9TCFa7KRmc7
AogwLGfS6p0/bQaa2v+bdaW31WFiBQI8f+l9MWT1grki+y/tSU7/qTDdnZ4xIu1h
Xl0ipTxQD/IZSyqCpM77ooZEUqFtwYbqGvVkULsQQW2/ChRrniqekBeobZP3jEhz
nAOTxqllmdvorbR438THMQf6HbG25Ez4MxUBQBaMSJcXYVIKoGv9AxMwmsZJaEiG
k8gZEYospm4ShrqXm31sn+2BJhGNfm0O6jQZ+/AWPE9sAtYMKteAXCy8iI73sQxd
G5asqzob+zGfhhJRb6q4TrxvdvEMlSigr4p3C4fOoGroxaU7xKq88Mzry38olreY
/sNFmGqu2o9ue4uz8aaDpJGzLxhEx3cq/7f9W4bX7oiIynQ/amxAhP7RT78f0bud
kkerPFReQXUNPtSqNwYOcxrgUi6l6VuNKsZcgNE+321YGkwWUPHpoQmiGDY2TuzQ
zgZHIaGeVrRxCjH8pGaSUp+8tUQfguMucm47Mce6IwrJSMymEhrKgsp2GgttiyPC
7rGufNfIlCWB3Nx20wk39CYFVx4QxMna0XKwJM9KMzM7nQGl7F9pTL2lLnbgY2g3
gt2gS9UldNj+qej+wTwJ5bk0OcALsKcfmDwA2RLIfA6huihgJMkhOt4/uiA2Ihmv
gBMdUnHjwA/n2cxJslqBh2WRbWh6XBUlfs+RrIFIewgNXL7Ie+p9Lmw5k93V1s+9
VMEJ+kt1zX+yD1ku3SEeupJ+SWi/7KIX1q/ir0JKF061gQId1Pu9n8YohL+tG2ED
TshymezREB5U3qOwJSHWl6Razkxvo8QU4M1/qH38IQkcIYtd2nhs4AiwGBQuXYRB
CbtkziTsD3tws2mCbeARyNbp8NpN29qlHE1s14WrkrBNKNib5bP4LofdMtMopUcN
UzEb1D5XQW86ewHhkcaI+KMOBKK6Hgu9xN7p+5iL7R4U8W2qpSDfdgZTTYthhhYM
CZlh9nwJ4+Fv+j02UQVrndk0tq/GRydiP257QU3lnCsqW46pkvLiDeBAHJ3YaH1/
OQQiADR6/Gy9D0w94euUDirzXwyYKRC7+bYMT1HzhVa6qNRF2iXBiRI+cJA145z3
h/JKBBqnvNlTzyWqaRHYxa+eJU2Md1wV9LkaRh7/i34yaSvow3NJXVqviSAg3T8y
TSL/f3kjY41IU2LrmNarqm/sZ19fsC8R9mceimRxZmHl1w97R+z/i0ObsCGT0r0w
jxZ3e1qdPPgD65m3kYZEBpgVcCcGd36E7nbuJISZpJ1DES5J6MozzvBekhKBeM+Q
0APx/u8cpUDrUYFv9qdf9H1jqflkM1cjkWNpWPvgT1rzscYNWHTyDkIFX2qFFl9X
Jc+a0FTB9Uup2hgVwkuKd8pj2Il6LKyrlEm3xloxKj7DJKD8cIlFjXnKozVcxd4W
SuitW96zT7FdFP2peK//uVXkZXQ26m5IzJnLHz74xK4Ccj0cy2kznxtY+X1QZbr5
Wdo393NGd3WKXQfKYI+Y4Cq6j/bWPu6wiJNRszQ9uOlPXrt9LcV5de9Mr6BlArNd
h0AdcFa8TvrponVfJoC1qwE7sjO9lBkXrgVPw3ermgBF5Y6PJmbjumPRsPpKuKEo
xCbmr+/LJaJi8P6YhiCz46G2yxvEy+BF12eE3XCTIRvKV/jMMOfPPU3rNieOntb8
AXqTatfvdccktmTj/f5Bu2TaglSB1IvjvrETDja7V3wmjjlt10WKulb0zNsiBG9+
EWYQYViss81vn2kWKGRMkYvxUPgOaN3VWPHlXWtGz1XCCmf6/cFjZVpOl4JFgIHy
4wNPFsmnAVsx1l2/ygtrkbMw+tsYd/I6cZQD9ZZqh0yO7jwcqzUwjpDjNixiB0hc
JlFDFaVqw6fUXk0Lx3UHOZHsgzUjHEBIxwRl2wVg/cSI6EudgrPqUTjn2/In6GdY
5Dlr7FBkoKQRIYSbDkRRsm9BQJ8Q8XbvYm3cnfoNYk0e5d1rD115OUJcfBFsWFKw
DKnixrVLeoRAEOQ3U+wo4qLO1uj00LEwd6OJKrbshcFhNralli2pAkSwWguv68Ks
EzJAeXZQpyogTQXsofx7RjBy1Np9QoWOlYa7QXMrHWdQl++/vGUZvnxRomheawKX
zNuwBOhGKEs63kCVi5Do13nAm+kRzFpW+WBP3JVzpmPB+LB1sUj7ketm/EkEbY9J
2C2hRrUcd4I3y9FS5dVNoRxT5tQgljbSQaQ6WrgTVGuU9KUuDa895l1ntASVSj/R
g4WHpXg/VU6ZybMHA2nIDuyEc2GYVrSzx55A9tDg2eJM45661BqylBj3mnZLPJ6r
uKmL4chBww6ZGriiO6QgyolzTSXl11ypW7h7Okjg2dP5q/iEPJVv/JuBVTUlF8jS
4PR84R2KlhhUeAeDOS8C3chkv+OA3B8HKKkwCr1ONnbsLHSxx2/QVWtIwlnqcq4A
BEhjpuwk74WNR8U8EL+JrzItfE8Ozkn7pgq0fP2V6bZfUzLww02wbt2nLqDcyLp8
fY0M3lxUspXMN/r7YIYAFWLPNQotKKjuJQ/miiF6ndTxo9HiO5hkdq4MMzO5CInk
LQj3BG0RRUW436Rtqv6k3Zl0oJDhxH8Oe51WGzqkXC8HR1nVQKdFxO+GaRbBbghb
QOFPHdZSLy2HhxOPDYLtloG6i5MvmaqByE5qS9ONGGlGxc2DAOjqvU+hKrlzK0ia
1x1/ehZ7NEf8aACejTGdF4yigMAyHv/yZGbUPYwpR1zDvFzpj+oijh/kOu71Ag4+
b7+sPKaPuzPZp61IALKhlOYIs7nHPtjIc9YtSTtGNo3jOQrLImFFGreV/aDTuHYt
Apl9EUKGHDEbxNPin7a2txc9tON4Z8YFPpzzSi//NVwjT9DJoLctLb4zanyMYGVW
Ic00jN9tzqwPIOHkpOy3TivXO10J965zOtlzPvORnJ9tUfPGtRKcWM3bIxR0g54L
kuRajmp+qYeMa5XEheouW8fcINKTMVAf6jOSw2MWB3Ix1M1ZUCFNpRuowQfiRob8
HeEZYJdb5+5JOhx0qy+fgQ5KKH+lzbqxsKuHQ7MvxJyPYWPB32psMJGjkWa0QUjK
t062juzek2bfZJySCFJ/070IfQgZTe5egK+Dhliyd4G2pWHrL7oTCImjvzJfBmS9
IQsYtGpqKBLiKuvnUvYe18I54u3U5b7z1hSdAs9bm5YxR99s6Cj9KH/0/QB6GNTB
k/O7dOyhN3e2cOWqIJfXlomDfgHxQjR/1z5Eg10XcoAbQWyrmektOqZcln9/QlCi
Xcc4Np1gHB6h6W4Qj4+BAGeUz5UpZwU16m/xQSdkfm5dOFiz15i8zlvdauviOqY3
nU4QDLMSoErhsTkpq010CmL41RLMMnzV45CG7LjK8OavAdG8BBKhP9Nw6cm0sMOq
HgsNdbr7LYM1lIpWDd8ks6OraDw8lu6hMFgcWHs9mrffXV5/XV3ndK9xfAsx6Nup
9qUuUKNb2lRFyhWQcrNOR4TWHNTKoOXjygmAoZrKzgXyh2Ef3oPdLD4r86+Y7IZK
rAY1F0ANyEGaNR7rAcwXJzlI1hgXIu9mnDBgY5pVKIB+eA0t3w6GlOuzDVEw1cFA
5W/kXAw1ab/gRnz953P5vIki5IsBDz7dKTV2GJM12M7EA7Uf7PFfONfzbNypy6N8
APlQoM7Lg7WuOYuEpqBt8kR2L8Ep99K87ThX174Ej+EO0S13FVhR53dIhDKbIs80
ELsnW+596eTpE2R9rWw8ZPkCcjOIzDm6jgMvof3C+n+HyWEEnE+LI+rerhEJ6pmO
XGPobkEp47dQENjWtSk5Tu/D15XexRiLDGjA3TJzryKSWid/4iH+s+lTxgCPEF38
FCzD1kiLpOOBI8Y0a7kllQ==
--pragma protect end_data_block
--pragma protect digest_block
LkD5vNOiV6q5ukF6/Cox4kC7vzU=
--pragma protect end_digest_block
--pragma protect end_protected
