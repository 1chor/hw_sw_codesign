-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
C0KkwffzjNku72TrKwLpJQgc0chm1WJG8VxVFooYEtF3RoTDNmwmW0eoWY66qrVt
csyRZ+ErM7+ywoViBavOxvsPqCwepmjCa/vGxSvt4xZML9Kg9In73M5+w9y2BJVG
Ht24Ra9+/zmYqHiJxWRTOBMCIYLW7TB0kWgDSCpqXdE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 34496)
`protect data_block
sS51X0IXyiy/B4Vv3bDDVnzoRAW7cs62MBSRu5s/Qysrrk6t/6Ur+Wa8KyAcg9T4
3DMTVg/hLOdHShgMTH9t3egF17SrfPY2bdDXl3FrycbXLB4Au7IoUN9LIQd3uy8p
sLpJvH2iLngMqNu/I6GFYBpWLGFbK2S3sFQYMGb00b7qru0AC3NT76AA6BtaAq6j
yC59i5UdT2c2QuxWmdz7y9ZFYHtLd1BQdS1Fxzc7P3dHBSk7VVbBs1AGWVSnCwbF
zzn0wHtC1BAyx0oo+upmCri+v7S7PIcxDM5ZjTk+BXKHAWfV3V8EPWKdQaF32BeC
DpTkwasdNG0dzb7IwwMi/OwE+f1H7ybumC9DW3Q65Kkl5QSLLS8Kz0F7fkvRcELu
WK8CeR9lFNElAMNlIZ0MFBEqN91fGKHCrAU69KRH0sqzkw9jh9zsL4nR5LLibciD
U0wG0xSTSvRgt28Z4CWLdyNlg+EmTc9q2MPNVZfgqf3/Ir4Lv0Bzts8Q9oDpRUR7
kOgZaNHbqOtsSeYjKouWH21o0KtR+GIUoCvCRAvtrBmK0sRVuWHRUzdwhPb17rkp
/ERiF2gOTkInFJ32ubK2NveQEg6VPyMukauYjOQYogbxXQbuDFoA6IvkkzYRJFQg
9lre38BROazuMU3qbOBYdVbpb7AHxa2Iws1f+I3AP8pijiJ9d28cp1hMHb4WoaQI
N5M2dLiAWSRPHVo0oXd2nzBALhA/06P15+gaSRNXSctgkDd0mDIM+5P11yMI1KSu
+3sWZkqHXYPmqpyFn3Hc5l/Zzy/nRXW5XuGnZP5m0o5gUpEHJW89qKmBnDZdHGi5
IUnM+ItfP/ilo11Ki/R0ikbH5JJfcUqyAS5G9LgD+qUF0ITPcALFX3WIuCSTESx4
Ph2E/1Uk0KVQVJ9tLfgm4deRRwUq12IErNvpgI9ha7TwC9iRkWj4f+EkfhjI8NP1
c5x77kCKmcrpU0uE3l7xfh26TF9u4SFWFEFLMiFBGY+umoVbz3DEtUNyKdafvcoV
FX5P5srXJd+X6PvBAI6rf7yMOK6QaY040CpYPNcGVEU0IbG17menEfxtm59aC4gz
kQfdychYAzO+2p915IARKEhjz80AgZp8cUirsJ82ZMTg/r5BSC6/v6Th0BQzfyKv
RIFXw0AgbZGAJyLX3NVQPLpV52ZWYTlMXE4IDFmG+HhXoJZiC0tJs4ZNzgFsEVJd
fb5hTPsJYGvvM5Psx5l/OtpDM/OnepGTabeypIHvG5GSDw6a3GMm35T274VhckH2
EyI5uOFjjiV/sVPn5zBFJn4nE6XtelGPo1lSCwFdRysNNwWQkrvkTR4bzaqVxWTS
9RKPfMTx4t+wgK66eFxYJwjMdLsZF8PNsau/+luSHap8BnubQefe5b4r00vUKFsJ
NiRLgFeaWGrhWD258bM/KepN15XBqAeyys0LE93iD+s98TkxulFjrGM0Gr/OYKth
a3jsMsULAzzLEd3fkgPHXFpmUs72LFXlOp+60qjttJGUYeJFjBRb4AJ0TLfhiw35
e2XWRZWVox9u+1aDy7wEqsHv/xfSdHKPSyVX611uOUqnqMeEJjTSpAtXTsRBYsVr
cdkxfWZ6+yk8eUGeyNFai5B5z0CwGpA2s6zseYVs2nmnhcKJmSC1UAE+zok7JSCM
Y9KV31B/SvkEairXpVVnN7e0ExRLq9PgAgMYw+lUDWzDJ/OGozdqd1w7Xc61W9to
TM3831oWFA0DrV74ifU/az4xsotsDgVEZBXbzyvBOcEv85o87WuEIY4K15cBfCM2
Fq8NLSlwWrb23u5NO5MKnDGkMN7LpSQy5ABfEj4gO+cjdKd3yyFMtQEEp7CBa0PK
wyzimTtulV6vk685uYvf7p9YbZI77TXOy8QmWV7LOaNpc91AEU2jCe6+VYU4//qX
IKveYtTKnEHijvgvbZScVRl3L0y82CLGlN5dp/KOBanAchqNQYHtdMHn3FuUfbe/
uh4PC/VKE8/sKWnAb5UWV9WcDWhd+ceFDT4mCLXIWWpVuqevaqAlEKrI9Unylx7V
R6lvYs+2FYGW4/HIBC3Fu+0ZjLoi0dw2kp/iXM6nyHJZktnYuHPh7RQVAZd9IHE3
pWuMk22EsPVliKzsKJa/UAl2BswBPyKJnG+8QF1jfqr15xqHdjI0z1vLNOYTwy0g
do9Okw+/EI/xlt/xUKNqaKgLsEbz7YFNQjlZn+UE+revWRBr1RAtyeal4mme2dW3
8WHMTv7sr2NysTpiAkJyDLnpnBN4ILjTDEJOffR5OIEjgp99aPryuT1fPVmsZLqZ
pINWM5Z7fmaLy0CUxbyXgULpTmnFKWllgh51Q3ouevmFYqQx7562b9x8QHVIYlB1
oAgaI1maHNGECNB4z/W31WxHw9FUTl1gfI1fRtKwYJlHzOjYDG5gkiFDzZ0Y5hn5
GRwjwsBQXoas1nrGf75z2DV0fqJJ2hbBPVh79h88fZmyGHLZ5WIE/2M32GKJpuLr
Y7ZQoeLKcPxmW2dxGoWsAGnn66P4qUoARRTIxjCYudj8mRacQaWTbDhsj5OEj4zc
E0xophPlcp1zG2g9kJrCWab3zh5ZuiKC/ilhD7tCHnTuVljvKsDTzyQx1+j3Nb5y
dQZ0g9SWXwIqqTaLa9cm5hZ+bqjcuzBZT+Q19l/HylQycKW9jrWBq0u9+v1csWRk
x+T+Syipg0UKAYLLy6arRG1QZj3HQBYe0QeS3+VX3p6MM80d3cnifQOfZvTqtrFA
qOfvEzpNbsbDDFtEbvMibAo5SFTkZH/UvoWteNJj4mlIuknt1KnWWYmlJhDFrk0r
93+bYJVFhhCc7fCTgJ1/gNPbKt/RujW4RSGBrl0Kks1kMIkJbi3PPqF9/hWmS6jO
71LG4jsownbx9PdBSREK30SKkdozRJ/2FWECf0pv1Ge/yEoYO7PDlTZdUJ0enJJ9
E9PCTk8l4lOXeT86Gsgj/kRXsqT8v4XUvhoikdKHRnjnavGaOlFCRq1kj7G1JaDN
iZW3PS8XgY95ea9qoYlRn44UeN587Nf5Z8Occ5XjN1A9P909WXzjuhu1m4PjAayG
uYwrrANsbLXSXoWlECtXhaLV/1uuMcV1Ve/oGuTsTib/L9gs+JU66fW6TR8fU2/3
6xaDa0u7KkhvpfzutlSSvKhllWmZKJrzfksvMnGGWO7A7P+iB7QZDebvyy9XOA74
wP/umOFNbS/Z/LMpMw2lkCxrAAEnfB7svLEi9YWP+2ApTL5JvBRwkf/1YXaIb8oY
Vkbxgi1fWS/SksFhbeGgXp5dmoaWjnegMu7XM7R/KJhzQ9NL5zz6KQWx9kd1cx00
Ukkd+97pkWz/YQl5jo1D7eKh6YBlPLLVfDO/fVBGys7phFGPZ5WnjGQzpuuXZeSj
lg+lbm3Xm6e2KAhT+KMMyCrJqla7zb3vTycTaxZo2/5MBDcjkRt3T0awNKXSxylv
RtSNzLaRkr9SEsRIkpLO6Y7hWC0fM5YRZWVKijHWW4yaw7CSmhw1F06fkq1Q5S1w
+iCwtIUFjxas8nFMLzUtCkjW+IOZ45ItFVRq9UsWl9tW8OPJKajuI/oK0U6iiLuA
OxLF9DXyqWQOx/jn+ptDF/WJKrKSzmBmeSI3ZPdFykXsHRSPvldAGn4SJjg/IwnK
ItILMLHNbx8Ya9jxfFkzFnlWM0e2NMi4MsXFQ4isPIuDmmmKK0VtOVeVsJzibH+3
XavwkbW8JaicdhpyAiZsLJB3hCakLHXE5av9a4GkB76XR5TJtGhUPJf5uYNNbqVS
R54iHXQ9fPAT1UpQ3AoH5Oni+e7V4lGsxPLQ/gMvfEiTs+60zdvI2ln+82DWq7Uu
Q91z0LAGh3a5hu9CUUvi5qTijm9luLQYwpU4liQp2jRWpmu6b9+sy8c67l/A6pc1
7MnvWvyVLMWvQywia+U0PCA8rUZ6qwKGGP14XkkfRwrHH5x3OwM8zDchKl38VVZT
GUy2vB8VsozKcFlLbuZZlcXJ3cczHPGXNtUInAJu9CPlX6RVV2lM2xUCJYcoqCr9
D2/HXFGtDrIuX9+DR/PkfqxvhqCOCFN5u03WAscuGmTLXfHMH7ZSRJDRtFum4wkI
N4hh4gauIdowUgOTgivR2+HlMf98LW8ZjaTETs2DiMakinAM2atmAV2v5SbumW3w
W5FVoiEgqbSHhdDmlih34O57hJiDV1flbcsbZb5rFNkgqBa/hYNNsXdkPe+wtFYO
fsmj3GxBxMEO/L7EgK4JOFsO+6n6znQpI42FNvB91NDLM6KhHyDU051Y2h/oaU5f
g2vzspvDMiZPukHN7gNWhDmAfKnb0i1B8WjPW/ve2MvccCE8ojY/1icJrRsf+ux+
hDbp+/ErjwoPLY7f53BzUQsL1pgtTUoXjqK9nSxlIH6YrWu0aDBgd/lPuHarnt8U
dS5HHWTW+iN82yV3xHPoZbwP1wWlEQrmkYfs5k+SM2YsLLOcAb66ToPw2fo2yLfY
xVa7n0wxzWAXtoSZPBVjWpFyg+JzY1xfgNZDrtR7fq9dGk1LnTPVTJO1VBkLcEYa
p9eOiLUocUj0ht+kza79TbpQZz0glO9FjEMW0CweqHd0TDYBN4EBp0xKj9AflQqg
Xy8OmGEyLOvMN+SVUjAiG2JUZ67ClqxV1aSxXgcV57Jrtd/LyCEmlq+fS1tVCpXC
QjgGzzoXzFcvzD3gj//Q8p0dQpv1F+/Rx6l6fureQsZfToQ/6S3I3jTnV1m+w8VJ
c+Gb9qCPQK6CF7sQjtzpPza4VJKRuD9IRapNiLyV8hc7s+1tO8iDJBdqru2KQ1n1
RKjupw0PxYI/ZHdC47npRpTzYAmGY5AKrfgxq0xTeQdpOq4KTrlnWdl6GkZy3WnB
2BW/jfXVkFNgBZZ7oboKMKpUqPfSLwM5OHrB0HWFtdbQnLvMdwQ4DoIqH+dNJlY4
IXNuW5obPAb5JQYSXA9MYdOFnMKiweZPPMQU3JUwJJ8NvqotARZuoHBXoNHRPO94
Z23t/q9YXTB3PsjM1Enqe8a0quiyLfUGyskSqfqkpDAvW3ZRYyVOqfKp/JpJeyhN
FA2CB9Ae50g4RA2U3OZUA4y9YDVL+JIWQikhzlQ5/aRX+/2L9nxdQyS2pmXL3duv
KgJ8rlrnx47gFAL0I7BeZNJdV1d2K70JS6E4aDa+stQnUGFjHTFkWF9OMvs7I1sd
nBqNDeYZGWq7fsuc51WwrISJVxUDnfqQEdE/jQEAcs78GFIZtmD32Cr+CKuN0rqg
Fv67EG6Z+jyQ50cOVxXFzzBVZZUcjoDqiogCahAKk84qu28NIvCn+EDrPyCtSxK5
1c/k220aELOd1unren4UtBZaqz8oqJKZ92CdWdvLN0QVmLAobAv+qlC29phqXnzG
HIihKXTdk5JSn2nLYqUkZbNxp4MEkU2v20W0gypUAKwZeGvvi/8mmXq7Cy9CVB4/
KzVWFGldFOcyLiRZnWBwsg3LuDGe5+Y9+IJK1yYJ5ebgFOzIWAELdmoQmr1/TS7F
lFaQyQbvJNYXfCdS+RLi5CoTG19cjbo8uU1sNVkgYBE047ZxFg8sUv8aV0giVD3U
D8upzU81Wv/Nq/hBaFVtS6aUipAy58V7SaBCRVi3525MYCGPEvGEQbPQci3GtbbV
qPPTtDD5mCEdRNW7lZyC6CXTkv7RitBKTgkUWFOsG+yZzfsuRXS/8R57OeYfUBYB
NKvCzbL0QmeJXXnV+ofOmO5I++vdkrFFHnl4BeMU7ZHds+n4japrwJMroU6eLLuA
J2fIG7XkmyGWVMfWC57HF2yjfNjhy4kYubZGwa+KLfF1f7ttLI4aw4O8gEAVR0/u
5ji4/+tXGvzVPedEM2D9G6wvY7UAZSZ+0wiGSy5hpu+ZPaJSzQRUi7eY98GhfM3F
1YYrRv2e98O9iDOlsucwFHEHIHkJblGMfyqi1ewAfy4V0E3n9VQM1/uYTgHPmfVo
yRFGr2KjbtprfTOUwUO5Ag/gc9EnhVW08HuFV4z8yCWvLpo0VOxAD12yuM9C//Zl
Sxj3IdU0hQOfAOlFjjGntnQQeU0Rk02gmnWkPEEp9dzWClppXOvtnXkSZpRgL1e0
h9j31Ao6dR2hO8nISEelstQiDr/lfGQ1JiZEqRjzATGep4gzp+LZIAneCk50LchC
ceAKHHsORI/C5AE688xAsI7XaAVSA2ZzgOBcPMc2l+D/9ojTOIOYw8rAyO/oNydP
InAzbzxmoAAzHxuL0GVkOnEgpiqXdDh7qBXhe6mQww4XonmDlqxgmR+P3Tpo9EGw
vTPuU+kpEGKqvo5y2fozKzAy8/HkQkCXJ8m6VKu3gSc5npv/e4wsAXKzTTWScUtL
Y8ds67K6WPJ24329+XF3R/P2NMrd9OXKgy4qa612ZXwdlyTIVPHP0fLH+FjNadVE
twmf+qNg2AG/9ni2j+QDSg2LnbMOVsbFzqk8aB5bWmSTxM5VusQzaOWdRBldxgVD
j2U30dKf1Qb0uGZHdc36RlzwMuXxnusGNl+SRHtluYVDA7BVTlqg/n/0lXkhqDHs
ILwJQEXHsrO0qQy4mtp7rf5TEdLpUM/KwO6TsyQgCQp1GfFatunKmqtVOEnKeKIc
GkiA4mzZl7ja1R8iuca1tfasUYt8JuhdjuxDtUVbhcs0KJnJmivswAydgHZPqs8i
yGnX3fF6o3WXYHjNrhsGzH3wydSgabUfuOpwAM7Djx1u6QgkRoAMopFioupndQlW
BsS59SwP3w1ahisiR6xzH8cwLgVgBaawW+nbzybVOMlQpE+Zy6oKD4Lwm0r7ipIm
+VXFgxpfRwIHeVf1UmDLKfpMDCTHitFZDMAg1uks956uINF6ezxNZ4jHxm2Fon3E
LGUU/x7R+43VHGXO++pVaBVcGkNC9ucO/KIpTGw8JBjX8Es7c2/pIrylH1y2SBbH
ba7U71qJbpLLRGRpI5NsyfhWO6/WsPGwIwQLBIMtDCNNEkeo3s9FSEy2XHEEhWes
3rX2o31BhVu9C6PPvGTvy8JmXuV5P2nFA9al8wkyKmehiaACyVTQ3dcGgzAMvIfa
h7w9rYOnZq8zaK0B7+WTNhqR/ZZpiC8REnLmcex7d6rmTgWjlwrs+IHlFxfTzA3H
bqSxqf6vb1RU7Xf6pStDgAS65QOn4DV3rtn2kwTD9iuPi7w1qlGltyjgBdB0XiFy
eEu0yTVDmIOXwYjL/NwjgdlbpYnqNczonFDuWB7bs8j18u+J5Lksg9Kb04IfFuM3
1K/iucEyiBM/B9Bc6IJmvW4yTwCSGkJosB1yy3b5NiEGDhYAmXb/0nnIACs1CXKA
bSMwLXpSQbW8X3b/afgHPU4rsnzoeMPA9xJ75X/sxZpCF6qHDXUCoCOsDMp8gpwq
qcx79dtVcoyizxSanrfHSTSlDyDpHPCcGyaCtcun0Xl50oHQpWqwRhvu1EMzVIdM
RtgQjR6+z+UX2cIGMYROz466fBZdGyddnrvE+tJlzG2IVtoioCyN3To40Fw6c+aT
bU9/MY02sPa93KkQLL7YPVMUmzHlNJMecABCjzWQo+nIZDT1RsLFP4sFuMXx+c01
1vJ/uWBbflCub9gBghqoGfrPuMsx/jGtcAV3oBD/2RTxt1q5brlqh75tEo4I9juU
+LNB9JZte3Wfz3rKVCFRFjnTZ0F/THJNo9/fVGRvdBIxbqiJn/IuxyhGraxqcS5r
IfiYF7YjJ/qy+pfv3Wz5WKu2LnJeLFDit0d3vjCdkG6IO7r3y9LKTr5K3cjKBIf+
L89P7BMGiA0OZuETdDz1XDl6gz+ayhnGn0nXEOSOUT/xP/1z91nY+/HdIw40BCsW
uoBSXisQ466cxRnqEmT+uFa1wZGPBORNTiG9f9gTp7M6Mwp1CT/JvmsZ3L8+MAO2
GMHhN01gtQY6R0+tzCMpSRkKQMywhsTDkcN4ZgGa9a1kuMO/+65XZu40IiUFu81Z
WBustuIC1bXyWGKDnGMPE3O9kLj4OFY5TXCBSSpvNDDGgOcUXLGnOxxGpK5owKgt
0mQsWd90fUVVGOavV7a6UzDML7qQs1pFsYrr2kPdIc/OufyW8mW1rOllRYrp5HJ4
HHZfw+JQ3tc347w9QmQmMtPkeHxvKOsYNc2pz2Tk5Ysq//SAng6BzNn+ohqXNlKi
KceaaLAQxqgaXM/S7/axZsoYdrXWmBbyQN/KkdVlZdmXMzHQ8rDWe24TPGrHyrIb
uM0CnvfqbmB8KON0g4+uOev8VP0mgGGUWU9PDfkXWtyAEnKGoyHtNs/Zj+nQvblt
zCG0PAtz7G+7wYwlq5//up6h5QdESkqcg3FLy6wW+adAh9qsCCElNVkdx/BlZsEC
f9IWM2JR/uEiQ0Ke9SLZuZUz8oeZZNlmv84bRAChdWQeZkXipsl/ZTCC7jaMzamI
0tTQ+4JLb6AX6EEuKet1Htx9/lbCgG6X+eNRJL/GF5CePZpisD6leqjrLJ6lkhf3
yAM95uNdtKfn+v+3w4cxRC7ttkgvTtnc/+ZNQjaoBcs+bC8aU/MO1R9VkCqk7XLy
sU6qM0tQThDIx2UTYU+xZNpoZtfGJRbW1df0Wlw8SwE+cmepcWqttftZjoPOqmLn
UryH4bN9W7MlFIe6jgoDEjFW7yLnxU/sz6sISYq5ileXAgXXtrU7q/1zRXri29cP
FzL7XMrhYDf1Hq85tJfSovLFpYPnBjcF6L4/RuG1WtE/MzEryQIV6SqfHU5MXioD
aONCBB07aoTziAsjuGoLvrRxejG/9uEaAWrXR+0l0wUubdFbRUS1kI1Mc5W3YfZX
QnfWXTEVY+8DhMLwFZco3Va88augIHnU1jGDTGBps+2+KK+zjHwMpHq27+awohtY
oiYrWQSmhjthif/4c///ErgnRxIOkDEJxdj3fxzrdhmniVkHoh+M4McQteEiFPYb
C/wA460P/dbjbd9uSMeqmxwd10bskniiS4X9DL7bNBo8BMBYsa/4+IjqkXlqeZ4J
Zf+cHxTAdmLX3sRzpj0nax3CDZW+p+H5+ZIS2WVKShycJhXex5vLpkOXL+CE/j7G
4IIC6mAjzksLPjvA98YXViwYGS+/J5H08ulRyR0RX2bb762kVeYcYUDA81kroBpB
ifNRJZn79zjCfDj3FpCVihuVqbTeYiLfh7nJ8iD/YCyyQuHabf/BOAYsG5MGertD
uFltoHOZCu2DQzCCT9xIyqmFiTX4DrW/QYIjhp/f4RygoiWDUSepLc4mfUr7ns/2
whr+Jbg7FG/gVZhxGMVAjAIx4keOIbsz8z1zEf+BGGsxsMh6D93K0u9B/N1on4AV
jMO+TO2CmxYz4/rXR1PciWaLqgk0ahSICD9FFFNBND8tViCy0ju0fY9yKopyzpSo
FtZVRPDxzvBhbO4N2DeTvhqmlaVwSKvSygLyAzQDVIIOT0wf+dLqBxMTA6x8zYTU
fGH9m4Ot1JbBUkEys/GhuHmXK2BSNvJwF6+yKWdmUUvu504hDJniGonB43UE7qY+
HfszzhJ9nCO4f9gEQ+cJ65xmkWB7cqpvsl2I1Xo88hpnyhu7Iii0XUc2XQUel1D/
van95jnuufqE9l+ZzqWlmL5UCptcJ9fBW32+p8lsw3e+hLV6c2Ap32NxNgtC4XOZ
VHSzg/RygPT79TTWb9v00d+Lg+jvSod94xF4XTVAfM0SWEK71imy2zJs7rWW4jC2
j156R75LqOcCKqvrhWlRRlFheMh+pX1RzGvneOJOLN1jwofOUs2XN9/6P/ragrPm
QzjCPv+hgFpmBVrZdz516zZyT6FEytqzBg2i2xWZYsRaXWYU58s+og9Y78QKT8rx
Aft6aPyhigfDnEM6LKyV4uzyv7i0zhKgLBpH/w+wFhK7R0Z/k/4xbt5W4YGYw7x1
3l8xkKrG+FvzFZwgW63TIjsR8UEMlSujhbaEWsNFYjD/JamjIrPgLXrYOHpy7uV1
f+0KJQmuRPZRrXxGT8temv3OJ/U/OIRsPFuyGjyDyykOFqKymM42jdBNVuRmQcf2
Ggqihjvu14mt2wvGD7yKvD75ChqpKMXUn1YIZEf2uE+BUl6ZULwcKzqzJ4TQcji2
5g48AlhmrWPiPu8yqK39HpkMNJeRaz67skEj0otf07fym1wwHns/M82HWzljgHhe
9CBoD1uZfL0qx6ASfifCOd6fTMgqhr5SgwIUf062CSynRlUJOds3oCVIgYQ9ODyH
QucDJbpUOjHt3/c0pfC5y/aweG8xBgsDx+qJLIVTIBGYzRFnP2rVBJ3ajCyauNwh
ZsB573Dr++liGdxmDtxATF9OJYVNFf53mnsrlA9lmkfh0TSiJhp31i4TtyTKnBVc
d7wOt32XZzvsnhexT+Rl+8hJiSN4hg/ll5UADYQRdBj3H4sJA+AUjvfFQ5G/RTbt
7SlPEIawFlWtLVgL2+KkC2xJqBQdPZv9xHyJ/gjrIXkCsbHTeAd032sJ/tF/nN9P
LLLJEQ5e3VPheliGaPb2hHOxltwJAxa518JGBbebiwJcTlWlNW/X3MePBE+sYu26
GcpcYU+/5h+Ewu1OM54b/H9z1/csklNzWaiBNhXV2Hinw1eYZqlrvvbAzFDL3daC
wgiE69sxlmkh2ih20DUatoZTQvfyPkxV4FtCK1+WzcFkx+Uh0fMwMSbFz6nGZIp0
IHwddDBnZF3+Kp4Nz0rZ/gkJDvizUXEcVffe2/ouSZDRTpPpMh8YnvCaj95GM3qV
/xXPtr6lmP6IFWkK0WLf0U1wkiQ3YCF/rtrG9jayJDPHU/m4espnvArPlLKNCzfk
TgIQ1Hn26jXcxBRyPhQGjdX5jzfj3Ah9JqlBe/raU+UgRu1MVUF9peeR44ySWIgJ
NRxq84+5unpCnNbPDV55xMxFAs6t0gmEPrTEjNT4StawdDKjDfO0X66Ol81O3G+T
ySBMIh7ilpncYg9RtFq3oCvMcMlaIVXfClqluYKM4ufF/Lao3SRLMg6gRf87Cqhi
MlnlfqVvyWPPaTRUTuCOfZaS5ttyO8+qK1TeATR2NIA6d2ZQKlc8NKDRi2g3pDT1
HkEnU7hM30TWTMuAA5P+v657srJnC23c8ntpoVUYwI4at4ixzT7T4gK6Fh5S7ql9
qBXX8lZUInY/af70vGaGdMQEHNDPhRMJXVI9lLtn3Th8GtaRB6gB8bc1oED5kswk
Zzpfzggbc1IW8dB5cW1Alhvs2qHks+9yzeFwtuknNa8QMQ07PGEpyvpqAV+H2qCN
q+lsIyODDH7BDiMd97htFTW1WPo/kPrCRgWqYrYi538BTqjF8QmPXemD7jJI3vUT
7i0c4Eywtb464IFB3aG8i8Q8Ox1dJMw3JKKSvqZtTxgsNNiCnVgUJR/aRv9BXmKj
EqKJO0xmWZp6VLhW1bC7+CeEV0JWX8UMlPgdgH4pE9su5obO4sM8polH4mnm0JyJ
JcZ28Utb0vtJHauxTYvqv/PpkrISYnuBxOfJ3UnXkogIrGWnkRCAmTLES+3mW5e7
/6cM6gVBMlll4f/Hsmrt7/aQzev4kKhe41PO4SbtiQ3VpPpuS7G6vW4O7+8ts9dq
QK0xXSiDCSFUApxyrDxY1zqE5W5y2WmK9TjpREaZQf9a7MsApuYK3eBQPZqQvwpQ
Kd98PNtVt7za22xZPUPN/56s6pa4Xe/aNnldoUNFMPfUKcBwkgQHjn3MYk3kdHly
pWXlf6wGJFqK+vw6wD10IdJQKgJy8UYNMtShc7GJX1rlfn+i6T9Lr7sLkNqiP2gV
zXuHT+he0mWbED863PE9CxuKPyTj18bjtfb5QBT6uWveUmE6mEe4AJuagvXHkwLH
E7VzKt4mBvkHAJI08vHARFQ59kMjxCOEktD1n2mhxRMmZOr/+VnJmoyOU2ERRnKI
t1FPZDjaGrrIIgHxv1icNzFSrxTgI1kqtHccJ7J/pzAdp7NWw8uF+4nlbbjdRPG5
r+/oy3X2uBTI6awJ0eO3OkQ0d72+GZdMBa4ZETausiMy9ybArjpSK1UnpBu2FD9F
PVLKaqStoQpcSbmmoFtGHNVognR/Xif7F0V1ZUcPm1PJ0eu2KloZfNTwhyZmY0lC
FGRAuGr7RqN2Z1gN/xRCKrFgvjxCWm6TrjZV4bHZVY+/Qt9IGINZUzGgEN9lA1KS
HcorLWpea75ozQC28x0hUs80hDqOvI0T85VNOVxKIU+VO9oHgtkYVioF7HsblxC8
Zk1hXTpTxFXBLbQ2szsyK4bmMBPHE6ygy/ZdspvPf7oJOWchvd6jzjT8pzr3QH4A
z4lwmrGcCKrt48nayojdGDTZSa4g1ydIAxRT8KYGcUAbiuuBVlMtm4FG/P78DM89
AKyoheh1kb7nkKsBKSQRJLuwQow/jiWkN9QFIeauuG8oYL9YlJHUTtHmpUdMfsr4
zjc4+i6NcPZNgBx2e+SuF8ifgRDSh3AP2nYbPTE+xD1UcN4IX7TpnIwilnA93p1D
KLAuIhhAB7DdkA53PlBZl3GHsXOp7JSzkArr/O/LlGYlAbel+T7d4rKTSk90muIf
X0wxDVzfN/DY62GeEcsgHi2V7w4P/JudFCoqJDiM8WX8DaYHpRisdbufnd9zsq08
/BrCOa2i/FH6ZVQriiby4atMqy1zycXcLLZxdzBwu3Zp+cxdWr6VIizOsg64i9x+
KYk3c96rvtbYn7wU1byJ19ePKbk9ZMUyf+YxaRuqUlnlFxRl8Qka01lEmcXSsAcI
pQ2+YVGnlAc0VZ99AYddfeULvfBfGboZB70RcIdYd7NqBEvB6otjaZKPCMIqkjUl
fc1PaWzwwGsaqtHJGh5Ddpk5gzFyPt/o1vMzTQrGEhH3FVklYAIB5u1p2uproVdJ
9uwBnmmpBOok1yIWzqY9r6etpsgZEdjzT+NpR7oGlcKkY/3/pjIMwQfYQxFFXSu/
fNEd3il6720/Wk6tc5IRMdMQKwMJg/iP2SwuPuZS5CHdmBjtbBcdtUheZFqoAtsA
+GD2/vNxM7mvZm+nsXcyzFxk1770mzWoh/Pk0T+OvpUck3XX+hbzQkBWWP/owxie
5n2WTDCabqgdphJFaecPXTYBy3MXftKLuyOAw4PM4c0fOBOT0fgLZSGwtp42h3b5
jOrakT81BYMCEzve8qU0y+xSoZ+QNVkfXdIgxElqswZc1ymwKzRQQsdgVzsSFoRh
hZqOKPLz02h1xNhuo7xsIyRTwQuhJBioFPA0ygtkDTp8qTJ+9MSjlsDJATC+trmo
1VdZn5w5ThxEasfy5PpXA5bLSrLV3G3EHFHOWfK2Gf3aXVhaulvRu75ibSs9RvJ3
4KO3efvuy7iriiSluFDV5Td2FFk3XOp5YA5UNnLwA3sIQOapH1C1uUZpt5CAUVFw
JmAU2ntCW7DRYU4S5Lex6bJ3vPZ+Ya0KMIyBc9sLH3irnTHWDBCR0twaFWBTngtv
0KZy4XZhWoik3DuR6Ip+njk5+ZNpkXHN9FLmGExN43jGr8XEXWmv5UREyR/nb1Bh
UlF18AMQZHNv13Rd9qYd9xd1sNzSZ7hKPNQmbmkltpHyIgzsb/9BpkHFUia1hTUC
6N6tTXozWD4A2fmnk4/H4cEGz4pxidH7/0z7C3ZzcmeVdMR3APF/epMsiLVm9sZW
l5RtXaK0HA+cdfg4HU8PuoNlttrU7J9nHOmf6tKd0mb+Ma4Mb/xu/8Kf1MS2K+cx
psmcWJNO2vFHYVyQO6K/GG4HedwWnUJzGaanx3WZQCZwh3Xv0qW4Li8fde4We3FF
UouYG/u81sNUJxSBywIIAVtn+aJSNgNv8AMR0VuMlMihfiANpq7llvax1mHaVik2
ALecvuelTsEkMAc9HiPxWalUvwDfcKDQtCvtXWLkIQslvtyvqCMMHYUSj8DeaFNL
b6Lr1GPxTOaaP/+B/CiZ2Y9V3qVpWui00pQnqGR0bLyXi4ZUfr6V68rPsT6a3cqG
i2wJ7396xi+gNcgfv1NRwOy3eywo8HlPq5mLk5gLryh0hiZs5mk4zGS4nWJhftCD
QAp6VnKci7tJcywCeDGx4dQ5ty5YJZDddQJugJlMwU/qPxOoIwoMYGsHhzVwTrYD
Gc6k7224zvUamd/cRXOGAEO9uj8o7Usnw7+0hTvBZwNg5ikBZ7F4iPrMSypCn4Tu
VTB4I1j3FN9kHgxEFMnTAlNJATuEcathvVXtZmF0jb9/QnxJdGfH3OeUL8/DDKyd
0gtY+47P76bDjvuGid9pouVtIRjkin5ieeV3Wo2rEo+tt9PnFptba6zvyJa7Xl3i
10WeX9biTQ0Yphs+nGfN4M/dUpJeTPEEuwB0Uw0o4vWitbWKtyb2i/DCvanz7FYr
Gkptv6miVEyIZcBT+t5W5XhO6hXU+tOK0WoSG6FW9q4sn8TwV3qRQppXU/KYIDsv
3eZByJdtV8oP1EpIyR4HyLNdlUUK3kDUE9YtbGpGRxE4Q+ZNWdUbTiZ4M6qQVWrE
eJp7I4FsDY8r2I4M1/Xjd4zH5QjEFPpX/SanxY93/yeGE6xjXjuq3PZWZkLL+IMF
Ojji9ahknYpvyD2vg9UiW4c8EaOqKv5qyLRUSjscB27KNpXAlK/HNyriohWSJGwH
t30lkvziqK1+01WwDzQnZgOp1uda6A5IBYsd3iNGR84WG/nKFtOrk/wE0Zov0NgS
3FVCnSFXNa+gf1RpKyfiPjgCshZqQwMO0DV8LvLJPDrLTuKoyT6uhYvAgu9jotRL
gCUUzZ+QViqj2y7xzxmNCOqXvJj0GyxnvDhb0VrRSix0TTcdPlrdMAaSIzNj3TgZ
JGB21q4AlNeGLzIF1iZVmRn+xTBuqzpGe+B6BxQ2spSYlXyA+ugsaC9CC9ut4r4Y
2uvyLLJi3ra7NT79W1Q16gV2FtL6RrURLLs/3SjIJZ4XGA5kNoEXTIgrfTMtBm11
BKx1OJkMn+t/XvvCJk296iFPTiaZQvXjzZWCJijDSIseWMU4JNGk4hsHpJZZ8J5z
cKy0fHmhuAEn6DwsR3uUnWj5pBvvu6qXstpic0557EgopX9lx6GvyQlmBO6Bfoh8
9Iy83/QGsgBKFarDDPiv6T962i5Z69gCP2cRvZ1HzuAwNH56GIS16LhOjyUCfeWf
izCx/2P7KO/bKCcyDiBisgOrXQEg/oT57gsXfyIyLvZRWdm+co0HsN1YVwDwZU2/
Y6lY9BRK5rWNbloZSmagsj8ERkB9TRDE6qnZ15IbhpPLCzmMjVky1GJz/BwcKejR
/M5F4XjEdJPVRKxW8xyY6fKTnLtdGlScuBzEkmj4dJR4O6Gd1wOyaQ2dn04oa1dQ
LpbArQD44Lz6eY3Ml4BUU4kFTCDXb5e74va+h7eEtYs08lKscM7S9chgHkdipVmc
+SHXRMiQHgGr6VpL/2RIKoHIKu5GDQuAVhjK90anVyLQEMa9DvOmZ6nmr0tDGGDW
NfeQg3LV6uLFdN3fRQ7rhCnVQhwbrCgpN7DPoCmmvmLOrw28Cmv4rm4FPq/Mo+gL
q7JQEiAihyq5+JO2how4KXJwSgO8BbUznPh9wt6xqIgADNuyFHRcvYIkX8aLOGqF
yLqkMAXu1m0FRbyVywNwNvN2DdvKg9ppDD+PQIXs9S3TlRdOY1YDqS/WvtGJYzp1
3ybJbo/k8xuBvqxmEspKJcxdguaEoI/acdpMg0KzOWZZu2OnqVKik0MoUZj80sMj
pDJZ4q1RSoxkrbdlpRLyo903lJUVOBTqu07Zq5ehhjL8x21v7pysIKBt0h5K4c8k
bYBjtsqFMjg32C0MPD7rUtF/63ldpLcuPhjjP/E/R5Wep830Q68Ecd2KuEumWVv1
KGBkOTdV6Nxx4lxzY7P9ukHYozYYD0jj4EpPMK77yRBHXnDcmHDJE73BV5FqQrEI
z3pCC5V24zfqsC6Crn+XiJqEQYcjrg3ZYdIjIv2j1zQrCLv2M10axdb/xoR22PNq
4zKvKML9UPwW/8QUSASDOUb/o3HGRc0pCHKag/O7JqclFya4bV25e4Y4NuIPFOxz
c01WhCjHvhgLTXdpfgR6lihtN9790bdpqP+c1UonPAHElwMvnLzExmBzOueP90ia
jmBy8uT4wkmdfSZQOE+5i1LU3x81sws/VCklqpq7NE4iNs0IbndW3+p0sVpw6IUJ
Kg0TOwKiGmQV1cYxmyOuAhjkOSA6F/v2eQUfUuJaSX1f5Pf7IKE+NiPIWX6CYqa5
+HTJSZq66d+MWfQlw9RXfPLQ96GogHy7HjFq3mOwFolRws6yqHDtf0Y00jrnsTGD
bH8wSJ8MBfk0zSZknJpq86cG4ybq1WIPLgUK6mVF8E/MAcRP6b6vz0jRlTI4D1rH
YCBDSwasBuW+DzgoCyZ0bEQHQNsEXAtPN3d0Ek2qngf8X4XoGMXQmdsD0PvDn3cq
xBKuhM1BD0r2yAJrbsA5spaZK+YBOOKerrolBLB8Wy6EMind2qXaCWx+U36Se6a1
csI8BKMGKpaZYUl6XZOQvI2ocnJGg2qzc+0saSEk06JfuBc/EwTMkzcKZrkPLOd3
CxiRFSLEGBgbnnJRIufYCJGf+9VscpoNAIoNtFcap1b1764PbxEcLIr1Xmx4DHyF
W34vFTrj0BlGHFls8cm9GE0apg+kLQKS15GBSmKmIsSEENtgtIpPBvSk8IqMv/qB
tDzkQseE+rM9TVgOECKIB7tL8nDF7zpb5hcjcCq66EZne1QpA929zL2Fn8PlsHks
1FND+FCVzb8ljjC7RoCJ68vvFTTLIQoVBOJp+46ft7dxlIKEp3EaOuklnSaVFNl5
t01yIjG7xwNoD7aD+Hiessy7F1QwdzJ5S/tAOkRC3/0Nkc2/I7RvwsH2ILckPmYO
Ic5NWiZjHEy+KGFoZW3qqiVtqWqIoABYzdxV+Y/9bLda7bGRDVaVZQa0YHN8QDI+
JP+PCtdVLPfSB6wTHWv9ilBgEK0Bm20Zd/ae9GQTLlvkpYHQhSNYs4rmEIlantnk
HCwLqS6HrJd7z6jXn3XGreK6p1BUttbxUqD8Ehtm+yqDKNuhJD1hCrC/VI2kbMWA
1agwm/mMLUeyM1k30bZ13dWOWOyBATSXen30zk6Eq+oxZz4mG4t9G9GwJ3VKm3fD
6xfAO/P6kHMCJDkYwuiOUo2DkxQr9gNGiamg9NDQm+K349VIwB6sOTM6OnyY1rd9
AY4Wn/GncYQa+dY18oGurfuGU3zDA0dwBcNeFtmjeSJoTSY2ZiPbnvnD0CaMwJop
wqX5MB9gtWxe8NIX+YS1XoXf9Xi1jbgH6KCqINyMy4Aa3mClPjjL/OKC4bGjbg3c
w7vNUuWnOIIznaJhlxMXmiGbQVtwV3TFTAGso05k/DahCabKIk30bmtuSlybKUm8
Sd+fKI5ykqRWinmKTq3WwrM6mQo0XJeTGTvuIJ8QO5tCHMa9Hz31MbXTOuRiSi9V
UIiEFdc1XdeTvNcn47Gb5yPMG7Sjc+bxezZhkvSNjvwjRi25scjKAtNkUUEZ3D8u
Ss804Z0kZhTmgUyxPJbw54UafXU1XqK+AHFFVgIIO+nISycr34oMyUqHPx6ovHUh
sNLjss2c01v1CIso7+i+83NDJyEUClHm3Gde1V07Xwuq/auTXr9DNs1khN7JAQYG
ifiu40vqTCevIQisUqN9fXmqC6Bkshew/eoB3sn8wKBfsPVEBVLmSWa6RV/YgKZr
TT6wUSCxVdhLloxl+0GuvRGpX6nNOl0bvqtTSn8fsYyL8FUW2rCWmfElpOUdn1u0
5Fg+P0Y7/Mqm2hLQm4hUCQy0AQh4+85kSL8oiiBwahy6UbyeZP9C7pHg0XN1Pz+X
ofOe9KX/A9chT7mKow6xVybrolLTbYKxDV86DjBzeNxU4doOd/rubGH0nGNiqSw6
6BenWM+VLsQFY6By1XnmUaKhkfLzzH0YT6tqltrfTPenvqgvlMH4WVyTCw9p6hgo
ZiP4S+1HiR9mkUUaGFKElPvAMOXgSMUxzzrwABAOF95Gl790bdXs45AssQ1JiuWo
SzZbx2RPqUzJQOOkqk9MUeNlwBHo5nVtMVmd4ZZfw7EpPBN/DLUXBXYnVSNyWIms
wjkB15nOgRA+c7C+VfbNcjdNy8yp4lbm+dmQV2GLVgAC0458RFsmKMcmp6RiSn/t
2IBMz2/PPGoT1WBUO5f3jeZ2MZd4t/uziqxKMPn43rkSWISF2j4wfdDKvepDWh4N
ysUfrR2YKD+29kJrEY8TvGkBnk/IsjC2h6ShwfnQhmbc65jYcY6ibR3RWxID3mcZ
Pf5SULDU94k/IOU8rvCY1DJI2ZHGI0+CoUQ1+4RrTQ0UmNLc38jaYs5S70icyueC
k98uPb9/SsBJsd6ADspzf5ONCZV3gOeftLEVBsZ6UCb/DYTitQw3omszuyxk3YGE
qyYN0xS8xuctG5ARGp5KFmxUrl4AmCCWaZENCVmh3/f23eyjOXcIPrrSJi1FSaVs
XHz8p0aBDQamO8yUAN841NVJ/wH/ILEfj4zOajiONpA8bEydM3CxGNKaBCcy41lS
hPdN3XkWRM5c7MWB25dBLCswk1YDcZBW8scPveRKsLmq/+g968wUI+gXkamYsM61
e3oytJI76ZnFMdHVRCrap/ePv+UlPXBTN/dSLI328wJURP7TbeV/a98fnVJCZjd0
lHHHESxOogrQP4oGsupwCgR6bsZXddLX5KXQS6kwDNOBUObyUKLxh8XVUoNRJsJv
UuAdZOMOekJtz2yxDmLluGR5eJJ0b732kJw9xvf0KntX7/yuV63tyEs6n+Gm7mPR
cqKC829wI2jtitlakBLROPUQeJ6KqdhJShKPfLY2N55YaelolBzfENh0gk9KLcfu
9uwLqwD+0MgfeiRSguNUNSum7mbFpM41LgKrgN9TVZz16b6HA0Dtkw9bbimjmTiq
A1Rw7WUzGYVUprsfX3sL5BYookuLeXcj++JLrLBuJvdqlXBJlfTQSuj2ytn6sjaO
dzM2lAOmiCUASN+FGsVEVYfbdsErxCc1vzOvlS3atLFT64L4ctJsSkc8HcA3VZaP
OEH/hNtLo08Lx2KFEvyJpam875nouneLu6podBF+6cD03u4/YVVaapN1XVtFoaIp
SE3HLYEwWIwQGiysBKR/87DKC6bMk5rIlJAVdufJZl2zixWvDZr6dfZyNimBaDKb
/ZhkFmH9n0hyhxwxZvRR6Vs3k93RHwZbaXQU9h+3u7/wacZAS1SohrhtfvIwj2Lp
a4Uv7kCy1WzABzZYZyT5LmWtNMSZBIOe6N0pWhpufRfeSQontAtGAFhugEMedVEG
LoQpx5fTELMxk0HDp2ywI5AqYN24x3M8J3nJZYy6rrqJUkL21Wz/k9TUalCerAkb
4PSliKq0ObSmB4W0SUfDHY1khnd0JpEDU7YR2nY9uv2u22Dz9XnMzO629PRqhBqe
HzJNyNTxdG7s4+/zgwJmcnsg5UuCp6tDrE05s7coie8Urq4cN3OPgsWwko8SiVim
YnMza92g2ng7UYa8A5eN5SasHrjirZwDNjiMrQmmIFO9bfjKFjLSXYbKO4Gf02Ku
KDO1iGgDgtPEAxiB+sB1b18JIPZFKYyEiHEwzDurdxwQETC/72VEIDzJp3culiA4
SrclakFJCjZPd6af3vj2mQiy5ArWxDcElzjzHoZMZd90Iml6lmBU+9yZh/05ShJ8
1pwGTWJHcRsoHt1KIMa4CpvmBQ545DNUcGgWIlQ7sp62jZfXZwBSaTTL5Li593cp
5UvW4kRo9jAh1TbK3ZI8vexFtbf8QS/i8GbTdAjFsJCfswEIJxWQgkkBq33cZ20N
rmaY39ZjK/UsOxR8Xb9sUO7Ls/c2FBT8pGiCurAuQCceuygUCy9oOt1e20huk5sX
2b4cjV7/gpbVcEAdXlDlmBSYaV+b3vjhmPN0yutpSpiGTUItk+DkiNNkVpmb7A2r
Yel4LC/9PUfQ8C/dXccKnMJQgAZGvO6bFWYSmjtBwSowaERP/BGj6/RMcMTtkIH+
rU2HANh647MxdkI8Z9mq45hbCB23HfTh2jdkE/1OhkioyuB/eaZ76pHQcbbMmLQL
hPZjcMGMbPKwBofl5goGtseuH9CoARfPpmUtmEP9q2l2vADhZ4ZM0uAWSNX3b82X
/Uo1yt2XXnVwaO9SBrRqGZU7KdzKrTiCIFLEH/Ld+Y5ldOBCeB2u6dXqf5ymvuSA
zp2BokVZ3vvGKlW6n7FKd6kuFMuFAPhjObB5aOqtVpf0pnbqVUSlCpSmqWPLVkyt
mvp+Ho4YEnd6Ser+jwXZv/u1k3JIfhUceJ3yZla7dJn16Qx+DvmYAktO8YECYJHJ
tVNwYFjBH0TtBk4c15es4u1dnyl3Sq70o7vitOyZqUbcoQ4gb3LEwN1Mon3nJKk3
UgB9BoFCxbRNabpV0z5YzPYRwX7EHG2fT/nDSLCedniFjriozp/6aevQlz7VGJjy
a27eHWsIfQn/lQxiEYUb2vvRi7AEklPfs+8bXVovDNFjhkbdrl5Ex46piWQjmsu2
VMxi8Hol5rjXD5EHDDZPDxqVsMwc4vq8GACgQWuuh7W2f4IPtszgQa85+d5OBllY
69j6+6U+xiVu81C56cCDZo9HIMLC4urWS7t0lJBD/rol6dYbLFtoqhc5Musieejd
F1YEP3MXYONq5rSMBF4eHdOzvMHht10eNOStycm7P00624bx/OXA5slqA6QaAfhP
HtcEw0DajjdZGA5cWIjHxeHizkwWMLGl+3Fc+bxrXGhAhunvvjBK8AlhoqASEa4M
U2buoGlTuorJpO9bpC8tUk9ajXolY8VELBhH4Fnms6+jrLl4Uehjz4ZUrmuPDevl
ro3GpLfb7gVmp95bZ0XjPXLYmxMFN8C39ZxTM01wAj3qlGybXRA/8EG7AVEQr2KU
YuOFWIYAToroSAQg97SICubHY0i/2WszLkkfCOOCyfRg6zmbtlu3527DNZ3LSz3M
Q/l1VUU2E8Szpu2A2//c44S8rXsgzgpZ+wl6ltAOMsbobEsjcmwAQYUxUE3PUUPf
5rNc/XOIkqsZNYy4WgTOFAWlT0J1G9/i9uKFzXteoMwMKnKrsGX5/IyONnHgKeXD
cw92j9Qta8HT/IaObXUiXfHxeW4BPyTDLKFV14yiWjnTBo3rnyLQ6w4CsrCHBQEG
OdE/xSvvf8LjC2R0E/JN1yYPZ1KwHhks0In7J4q/Xh0wE8yz10CJ8ccQ1p3aaR1w
r1l17K2te70fAWE4lmXVa0+XPt0YJ0zZGZejN9TI+0ETjtVVJRyyLtx0qfOSAKok
fbK02Qb1odUdMjOyJqmmCeSL2UbrPr5skjygffC6ssg9+6U5xX9EXTakd2/UxHeP
PM7RKV5Cx3txKkQiBdpiVqgeJVasedNePKp278mQlnkEVCywGabrD+LowFDF3wE1
vF5+XdByk0vna2A96aAWTfIhhSSz8euqipSYKnYmQJ2/8M1kM5U4JYn42GvMI+33
pTo5Qgfv0hQsJhp6psMII5iQiP/fMkgHV1SfBg4kY0VsLiTXpJ6ZDyIiVY7nGvex
B5w6NK5wn3JL/LNLUUrvZKwurFPbJIK1wo9ReaJonJ7aIcMl2J0VWUiAfyzVkIpI
q2jXdH11y8XfUpklG3j7FZRudZQjyIW4PmsEuY6uYYmppcHk3uZzhLnqsEcILXM7
e2Y8fzkUeuN1g+HjqLzBs5ue8baz7c9manz9k2/7CcH7SoMTPzEz9vv0os6V0wH9
rMw6+GnKd9xXcmvrhQiV4SPruWIykO3v2FI948eugUZxC9xTBHqp7/qJE2AuC4G8
+xoFW9RMbpvF2BWQiP/fV8F8rh76y3iAiOMeAP+sO6wQrb5Mm2xlE26aGFrzAV0K
A6Fm2OechAsS1qKnabenNo10SetFEaBjBNxl3hbz4741L1mcV8SN3jlDplZKCaoD
qsEIZSSbr8Ej464dIZL9mtGpXz1QWGgwQQSb9XlyqWT5VIwC3jh7cTHRRiI/duy9
tw/CMiOos4okHKopEIMb4DnFa1daEILdlWmntDniWYuaofBS1aZImac64v5X8n3q
fGhxNmxaY4adVqhrXKbdtlXZWeven15ZSClf0rEa6fVaeZUQXgWF2SQHa77d+fF3
6CWqohuc6fApU1cQKXjgQ0mlBvsHKhiJDYmSwDm+mIifrrW4TUbcA/5Z9sGkhCHp
V1+OtRITO9F5EuzfwopZPhzu3wtpJqBZBOWz9g5+sKQw999e3OMDJCIEwKkOD7zX
8kVSI6RuE//Xw27ukJkD57jbV6NHfiA6t7rcoVC3wfNi+O85A1b4i4SPWXD5jCdH
0ps4VC2lqDjma5JjvDzEhJWcIQxLaF5vWp8Bugnf6Qot3iHm7y5enncGqQs3due+
ac+E2yWo8ZT0ycYsCi1mlry4Ya3Vr03zxM67Dxnlo8Qun792osDwHV8PVbll//Zh
PbLDzxq4O2SRSL99QN1ZrbrzP0NfcN+/o2jq8nH9mWEiBXnZnbK2c1+eR1mtjcLq
6VbqiM94zLtsw5Po7CgeJnKMogqOQbZZVRpPXr7roogZHlwjDePzXBRC1AC2VOP4
MDlFeRIWtRINI0bogLPO1tkUWyi4S+ZO+O+EjFMTKEK3gmB5l+nu/MuHHaYSuwNS
IYLEzNYMIWI6j3PXuuPsH3St5Ly4ThhMbKsvCOPmvvqfK/ssy3yCotWPpeZzlKTA
K/c1h509JwlRNGfzvMjKAPkceYI9JnSNcT7iJNaXm4oHewKvZL5ep/AYW0ocp4hu
UE3D+nLC+jGsirqvdaojsompF+yZJ6YpDcGMqrp6C0ZFHkMMKs0JZ2qrHrA1oa9o
f4hI797t1GdyNqlLpNjOJmlolQyYYnMMK0KYm9pHMzm5E1SZR+xyX4V3dJwOonTt
AJwMjNGLapyjYGiulDFdVzt4dQnTYZo1DovQz1pnFf3ZbR62gV+WpXhW0GGrKilY
Bm4Hd6mOm+xE8IjwpeC1EwrE66nAQqIk0QxrUXkyY5uW7UiuxodO2vNakOxhtG6m
LiNzPXy43UTw2Y+286vcEaR5DkrpbIIZGPLuxg8cInlZWyB/VpoZSCGIH0eOSKVC
rNj/rEFYQAKHJb6tUGWD4LiLvs1C16Ky7XYe+J9ZgGSANQZTahn8a/WCW2c6f8C0
E+szeINdNdK82TX1K0RN78fHZ+7uzTTEuUlCA3ItYQ2iEkLP492LWD4mBT4XozB4
nAAkr0Qbx5Tt3xV3QuWlXMzC8CR1hZeALBp3kneAPlondsWIKZAc8C4e4E8mRt73
IUX5ySB8AThiZ9isWgaD+oDfMqIQSfT4r1AN9MlzYz2YO1OLgiDSWEnW4SaFDCgu
ydfhb3Y/rLiyDXFF7aV3luNA1wKN4gMYSMoOx9M7l1cItp3nFLoJDPPZrT7VE271
RCim2aIfPAoVm0NSWNEu1GgopL+RKpF303+jvDwEDPIKLjpnFtJv2Aphnqm0YFb3
9rU9I6uCSTNMn2Kp3wv7cl80OXjewWH7EB5Kj69q3VFnO09dwJL9FAznS+cpdYXu
Gsiqi+6LKwr9bB1gFOG/Jx2Xg+tobezMTnDqkQB+TlRmJlN8sG5kIqVo8UvG7lDf
i00BFIs40NPGAYrJid7ZoCszqqpcpMDSCtBago3QnEDjeZRW0T2Gc2G7tNnUxNY1
wOKTbwj8FNlOd8x9/b20wXf8xEvUn8ziuBAwS2hSHRv3J+7fwwxvzQn1OzwZ7TiU
tF6m5PljAtNi3SruU6VZnOhvZnBn6BFdyU8Pu+WmLqKMRScq7ap0PX2T/wnb48yD
Sj5nRcKoORw1E5k9Nnn5MguixyR1BC20du5BcTP8NfofUfTWpXyVBPV2oEuTwd9e
ZwTT0DqSODnIMa1nS1Cc+HT9GmuNXaI/vkp2DR9lcvTbphha+cf03BBpQp4C8uKn
6JRqUXzsyA5egrgeeCgxODGbpto53csjWbBoPz4Qsk2STIj8+ATQhiKqBGO5x0Jb
l3NbpaMjzujUeLoyQ461kBT2sMt4bb/GU5m1isXdHXzvadbAFKsVBn0mxdJHJKZ+
eB3BIHFi/an6BUcpxl6HifRNtOnjFVYtBboBvL8DxoS81uZcLdLFQSGhETIP45ct
cJzUq9XRLyGY6mrYZWgiN/TnJs+WQRMJMN9wQTaRSuwaUGe0ws/QJoix6z9IHZXu
O7VHKODV6G7E4IEcwBclL9Xrc3kJ3MF6UCjXFTkug6S36SuD4mZHUvlEaybl3cWf
n8C3bbjB6X8YxVSd1kwKBN2TKrtV969VA28pWI76/CI+HQlhoUjmuKHM0fK+hA3k
DWY5u3rzhst7oaimizoRgUozQawBsZvrLAGZCdl1/zbc6E1odW4DOdm3lAOU83Ci
/YMAjUZONsefz3/wlQ/3dn1NjbCRVzSyNqvFpGtxl02Mn/2zov7SGfn5VuyLuuVz
99jVkeSowAJUkJy5H++tY2aee3m5/zkwvWFveeQvYQNvGbXqrrK0SLT1lTCi/j6A
VtMlSl/KAfdBRP+Cr8VzSV+ySh6C7cZYKrmnGl9WHAnp/+UQ879ytMshyM6+VRDF
RImK+41Uer35gc7xqWGNxx4+qGVS7Fjq8EzsLScMipUhKTYQjYE+CMJkMiIla1YA
QCAmb6LATcDW80UWYLBnX2sFMyjF3DlPRxo91qJtTFMhNk1mqe7TbJFZg1de/9hJ
8qRetg8s4HiumO3SEwlOSMYDmy6B8KM/vVc9l6Ua9vPjai76bd1uPRneTDRnIJDQ
YgNRLx1+4UrlfJjCPGj7JbuujtXt4X2EeV+k2qMebX6PJ3VA86iaBYiXljrp6rDo
DPQFMlNDSToj2KSIZwvRgNx2lBZ3b9zkdzhoz8lupBuY7l1CVUxpOF6bbLVGlqfc
U2C5PD/HcQSl3zKtPsStmWQVM1uFWs8I6l8yl4vnEHdcU9DkTECJvnbXsPTCkVOC
nWPHrY1j0/U42gyRLwEL1KtGmMxmxaWkm25QTaaazcXuEm26JYczcnSSPNQ+BiV7
bqFSm+a4X5di2So5IS/KWDBy2tCkjkH+i2BT6CuUha1emnR8ori+QHT9HvQGrbXn
hvM5UbNqdisI2h6nTavVb2kGrPiw4M6Ufm2tEqcO+NzlY5sjFQOEz5MQH3DVmzhV
OXukz0h1VFUprHKEGiXkwoYkjbf7MHTq5XKirI20e90hKNKdm1ezHsHyav/h5UCn
eJcvhXcJDmuU7wJLFGqEA37Vq6ChKLWmbENUpfBMlVdpXuNEIpwJCQxduZ6C3pJR
D5Gm8+3E8Fq11otarFpU1/fSDUF4X00854PCVsN7r2bO2kKloXt99dv861h16gqJ
VkP6kqjzT26T6hl7ijQiC0hPGFbmceUDHLdRGBWI5muk9i5NKGILa3GVuu65KSdh
iThMmryO47M3mWicgqx+osydJJb0uF7MsF0iylnY53yq5lFrlaBL2YcHIIxgPFmD
EIaQRKjarH8CoBeYVDoO+lVbrcrBD21nZSJxpcGdsLdi2ZURG5DpVXLkdcGsdert
8DGbPuLjKpiN0FUR83f4hQBZqRuXu9GLfF0t+Qgs5GhSYI8MY+9YK7uuFHRAxr3C
KYG0OjIZ4+Wss91AygzFwWM6dYx9PlHm2v69KXeTjf4t62m5MIJ9Op9/THIkJmpY
7YGkoieI7NFJaLiRem9rb65F8Rgwo7GUxSOQrjiSQdBrJCKIkm0NzeuIYDht9DOU
Yf1uznoVeSEy2/mIZfTGIHMOsHzPaB5Cfy+b7wbwgCwJIFKdt8a5Iyw9Db7XYv2A
vp1Pt5jNnedeC786SzrijpANohpZrIcJYQcgpxNUe0xbs1Aq3zY1lrkFfqtTaNuq
9f/AT+nqq42vku7XQfeAFyngaZsudz008cSldI8hE2hAKMMMg/QLkdEh5ut/xIYt
Ns2ebNqZwy5ydjNUYwLDWr2XsWJ1ytNxLpfF/rnllaZ/7w30LZbHPDJGnPd7XoKg
as7TgVGgKkkckEgPZhcon0CJ7LGjDe+1PY6+4+KuW9+0D39HQ7tnUUDVbJmusWke
1LNBR2zxvvQgMayls62rvTz5s45398BXooVC/v5rtjlQJ6XC4LzmsGucPUBjDzOa
pj69UIEyUmSN2MeuLjXihCh496LbVb/ecr50+zdxUOw6MYYV+9S44/1YhMDsz+gJ
Pi4R+ytndbVgTDWoYrAaFsyV2Wi72N9bMYyvMFo5Hppf++VR/dZK5VUZapqdH1hw
F1OL2pekajmFt8CAxMmsyRrhulvZzhxC0LkZmKV+eqIrfEyMqW8IUmLlFJdxSW9n
YTf4abVc5nv9vAhZ+llAC2Uw0NP392CoqlK79N3qPFZcpAqjxLpEFhl4+JVP4kMe
5gfUYug9xv/qqxgWQ9u82tyToN9FEW8HXtwKLTSCXnY7T6nSV5R2zi+7WSeeOdYu
q6ibhGLBDjHGtBDTop9MMCA8ZMO79IRBhbClKh3MZLmuM9WHrTMctEw3FKNeHA8r
5ONwHdsgPsl44kwE7xzneGvuK6YfyTjszHfeOCeA7kgJklBCh+C2S63aaFcD/xUn
38sP9zpp8azYg5tckahjFsx+nsnYsHygKEA7AwcoXn5O6UPmND9M9ptZLAWuBtsk
HakmoVGJBymB29bHpzPdMANSlbPrUv9o927gVbtitYRnZ6a+MF5xkhfmqvJh3qjy
q3V3LbEeQYcEHhPRHuijNmMnAfIERhidvNuNcfHJjTYlz/XM3U2bShF1oWVY+y2I
D3UZF3lVyGjVEDyGU+BPZJ8EgMTLKJQ0sUgoYU/NZ6U9pBR16/kKwVk0t78Wui/T
XQ9WeMB0/5jktxpqy3GaKumQY0JPZ55PiPnYoiJU/WCTYlmg1tlU4ST8ZP6G6COp
5z7WZQZKnRHG9O0cu+fBi48DJjcOJYiZZlNmh+dvVG29BhT7y6L/SxbIz+PmqvlY
8Gka6HaCPQHnS46oVkSFhD2Q4td7YeSr8wrHA3bQvUo4sS/SakDmsF7G2G9Zjlfz
lhyusd3QfVQQIbPV6zUZL24A9TfdVQ6rWOsiXNnU1ubAf91hI8tj9lG3lpzhvgim
2HpxwFyLRRoTLMrokiVPUYal07Cl3U+MFoJzFfqZP/l/K5EAp3H4w+EYxz7JAsas
JukHvZGmk3skq2IdT6UBQPXKiWKOYD8lcy7Tzy5FYC4RGo/ty/n3hcVx8I/wyb90
sRw0mywunkxnGULd5xJthvTUARa7knnPvEJ+twr5PtdOJ72ip90smmtZTFhQt9T9
RHxbqEdky4YW6XHK094Bn2yPP1AY7MyY/kmMShpwEb7/PZ+9It7bpUETjywVfNKX
y/otFjGpaGJJ1xOSQ3g6D8oA5QDJaSxBUuqt+JA/GKx91Fmb0fEcVvFd9l8FA08f
nIKN8fbS2l4bgNKD2mqp740hH2/t9te/XfhtTWrq6QXNcxrWeqZTIZUtAQgB88FY
HgUDxHnh8acF/RfnlJP4sbqBW6mdke49uCcNlQUQMCYIFMcAVBNVokWbJ0jKjQqn
joYhkVkOeY4o3G8OVfMCltBQn6hA49XUayPMDiP92pf/Z2Rgg2ADeC2TFF5HE8J3
RiBMizxDv7xWkCf2MldErSLr6PcPmYFju0KfIgPsgbVcuH3TnM4lkYp8+r6QTael
RRKwMsyP1oXuTvxCfqbM15czEvDH0El/if8YGUdJBjfUJabuLr8qKhm2bnx8r3ze
wfBnX7f/B/ge4GCZv5UQPAbeDnLzf0E6JVAL8fC8Pg/ZdpsasKCbcZgqyrocAUEX
IDBRZj89zF/bCGODRHse6kNNhmZ4paR8WX4Pi06jpgUDegyd4j7YrskD69vkEgPp
SdlHZns66TB60t8hRLX4aEM3D7GVbJJfrnVYD47H9pxg0HQFpkKCzUHtJtImq/4+
q5PaZhqIqSC3/WGCumX3suU053FRpXEGsp1gn9YcI3tBoyWq+xWOcNcTP+0LSmOP
ECf2LDpGWjUjoxgTcdn6Qe/lIkZowbOxiseQFwieFUDs1a1bxVU2aon0Aox+Z4XU
A9Fg+O5C5/ikaWRZUc0EAhJhuN1yIo0Eb9S7RE9bYcnobM90kG5jNuDlKZncwjP3
mmz7NPekY632pU3azriPD224Ny7n4y8nD+NM3GZWlgEqCtwl+Vh1QQ+oNLVySrzL
g/tQAYshJjTYiBUfAvlqT3Xv4nRIVv4GPiBD3WkSFO1bc5Q15vRIaBIHDCowz2oa
UEVhR+DZWHZg60JwtSljlvjYPbuPWU8rMHFhsQhMiZj2iSXcueN/u2Ns7kW3WKFw
Va5mltNWYhzjbReLzyCTCBJVGct99h3kHUKk3yjG0EEgR+Y9oPzefjqZboNk+Dow
lUrCX8c5nX0i8YbCUFVzpj39XB3/k/W52rWqfjm8TJKAjls3VAGV0Dna67J4IhLh
9YW1n8i5eoDWYnLzh3awHblZJsjdtq9XRZB00419kav34ZoR6b/PjPrMlX3oCLNy
vpPaN+8YGEC7ew0cTy8+3wQYESEeVAot/telRXX0jkQiOEIAc+8h5K4+hJyYnP31
9PatG/nJf1TxWcSdY/Ck1Vwzz0kGt7seKs40CSwgeyEqQPekuT3jkpLoqIlkUx4B
QvmrtsBoTr/qQGbo876/ftangcEPpyJ21TlLus5oNnPDu5Gmc0/KKlrGhFoGXGWh
DlIaU2XjYQS/rRYgP1VWNt1h8XG3tEX3gh3WAv8fccHnPJ+amUJwcXfoQ+WLU+ro
38HcJzC3a/RdeoyNUNvqKece8V1N3D6YyCegd7rq3t4VSu7pwY3hDDw57nWod4cx
EBXAjSnU+bcrpvhAC9QUuH27HkznEE+mkrjXMQE9P2+teUP//mRIn4XUVu3K3dKZ
G8hBRFLA78iYpgymZJBdzeSP51bxcNd70gqj9Gzg5xPnybi+ULHlHDDdWp8ePc9M
IXvdtf3hswzkzt9wnsy0m2xGWwyW2pL77UPNrjuCJUJSmj+MozTTkRiz1iw9H1f+
d30hZQQ74fEYjsTM2W2j8wvM94F+snxoKZuKkEraBo0zygG9ovcr22yval7AEsNS
6oL22dgovEtrjlvg0kF6+pOoHxe6/15cLWWTOd2aktinf0qH8V4Ga6lQTXI+25Ng
hRxLiGb//wLNfR2T63WrYQWQx0DNQhY2Aq2RRAcW/BbE4yJ68iTfL6hWPpUCwlvI
n72KVkhqFrlG0yOWZklf2KRH/K928evWdTSRG13wPl84m4ElpX0OoKVUgmaGRrk3
7DjiQhbuEQbD9eUktYCVWm+zXVke2/YFKR7+9BrFUlB+NOHzq3sFQn6XUXDMzEn1
RAM/tOrAuZXxfo/h+kr3CzF3nEiHNel8CKoueK5izALg5hpQBCaeIdjUCVX9KPaM
QNEiqTfHqEI/yLXXaVyMmey6PJO1R8Zlv6vg98R4UHOn/oNJvV+H2MExTCXyFgFK
7ZlMv1VmMwoiJDuU/UHTJytqpqNXDnXsNg+AalNRPNxO3oWs8C17bzpnTKxYZBbe
TowP45y52djzTuVUn1xnrOhKABT6KMDAMjag/JtdduS3dYZeHS6EfSl1KjKaO670
q9W+OGZUyWOk/9RdEbFbqLUWnXxMSra24/gOtqoCijZ9dSJwXqEL3gKltHbayU0M
SfQaXm/SrIc2lnjaSp0oFBVoXzRb/qMuUsK4/HN43wKtWf8FhtG+nj4eI6jWmi91
haPFbx+vo/zVLsjhxVAxytIiahNZOqOYPbAC0oqdqkjh0K5lu5gmgwZjTnctd58S
WCUCbTWJVVSghKl7cOANU8Lqyq/knzfYeWN7WjN82RQpneXRFFrNtQsLVZFie6bE
TBc0KN9mcRrtkSxqCaYXHFT+5L4At6bWhjt9VlWpNGyNs1dnWIfpgGHlnUVdtr7B
VZlhPFsvWp5xmox4aRMuEECtekDKmGj8vQvuxgDbKC31XooqGB3rI+xXvlOufGFo
l6pY4iBJhwlGv8WuUSqrgps10+WBo6NmMbJXmiPemXqDEnXW0Wm04BrwGTmTWz7g
1GUFSbyOSREVEt1E5nwanoqOlkRZmgF6FO5aFuOurVRipyfw40p0jsARjx4PAPCM
b5BFc9iGOj1oisreYyBKESjP1Lulz2cAw8nEkVzve1hkdScDxCQZY68dZ5LyeuNa
h5NQ1D2BOAcS6XEkKamk+5DgFScP96hBwEQ21yN4J0itIfY42iM1xa0zNSgnFUFe
e74zUGSxKrJtrVMZUiup4lI3mMMtTibiCfTYg6Kwdhmz4x11v///EzGDHvbTsmTA
dzVat/UrMZtqcXKqpNk2ic77QY6xzufnEReEYGGoMxBqiu7LDZ0rILwhpMWgNezH
cjOWzTHsHKuvgoBXIMoX/BhiqR9m96MT2N7Bkdr6EIhxBG0KuRtEHG1vqUTYfhsU
JtZk/u2TMQTMabYIK47AhlLlmkhbztKIxwFQCtynFeQqLCxUN9yVHZKK6WSJKZFj
ra2j+PZ6vnIs7n2vlqIZiU+g4Chlg6kZhfwCeYTzpeFzdJghhlO1IzggdxJSn5GS
UphmTk/FV5U8kTyQ1uBQK6Wm6jyONtwYkfbBSfLhnkt7fh0oMH5VkppOFsk/JtUH
cqEAKp8sNfibw5NT0wYiYixZx/1H7xVc8M8FESSNdapnT34+OUSiindUc2+zXHn5
kUem+W6EX6VEJhI/47nUYVf0eiZaYBoHbZG7wHGfPflkccvoinzM5BTrCYdFQJxd
o+w0kQR5LXoaazWn2R5fCMwI+3tqPIeOzFl73HGDnVTpr+vOu+6otAPpXLbUkcqt
5S49Y82tP0urVten9hJeWiAnBGC265m9FvID1NE9broXHmuNHjvEFEk4QtwQ563c
zXbx2V63goUCUBE1XKyWWBQz/JQki+rFE6+xg8OI8cNY3qfiU/zFa6eyh2RFVB4j
YJzlmYnWLRn0+tnCEzzfZpK2Beq8qVGjeMILKElKDuZFg5UbmRqkytuujQ0HEalq
VXZgMFmMl3NkJfm2UxQp9ZtE8Xg6Xy2dpdWkxE7oQgxIebWi+MjCkQ79LiVdyte+
TZbiZ9uAJHO5BMbuvEh0womRrv5k3wmf3dnQ9Y7RvpyQHUXJClOp6ARjG9m5IWdR
BJ1RxGGwkbT1ai+CG/cLYvxQrLkcRX7wkTGjWrc+AUnHhnlXcdqi3YR2oZlWrRTr
3CpOFI8mwkTGR4oBE3qZz2TgyzbNxk4+O0LymySOMPcq5BKPCZXYEzziJu6XWE2C
bbvYihTAioCT3Jc/d5oGYSdnqyPDNI8zyo1+9GMZtcyfambeYa14ox+0l3ORxxfL
YmUUeTabFsQ0L7BfXC8rxnmjkpoTIy9la9GLB8+/idvN2AfSPI3TmLdLqH5v9a6W
Z35Yvqk+P5/elGK2EH1ArghV30U1skRA4AWj8zccSUZeMNRjyw4OdhWm8MwbdsMO
wga0xPDHYbyLISCdV3TRojsHqqX2H16BDMeaEQNp+8QFTDFmkADrbwyZ60/S2Aow
HOxIhOB4V+UEcwO42yApzwR7MNo39Lrom2NmyJhDtnY8p6Db6aHwB9RhjEWPBhyB
Dg/smG+aeIFXfjmZsehObOyvJtW3nPdcWtaXLjJQu8Luzg/pjQGha2PuDheD9hte
P1lUfmodBS/r0Qq6CntvsL+w/xa4zk6FC3tMo805gxL2Ng1qv+G0m6+Pbfa2ntdY
+nMqjcVy+Uv/2GmqzFsuC6c5yyVcHa7lZLOuZDAKPR5wTKnRmuf52jROzr69Izy6
QNOmYGRqX/T2qxeSuSvjTttGxeFZAJOvQSnAe1g8UM2NunqysOOuzIcxdkGx9AXQ
yorijfAFvYTvE5FNm8wsiCmLysNzHFyDVWBAos/CgxHyO6U1i2MWAvjCP3T+UW2v
g8l1BgS4Xy/ldX40jC6DleKRd41WWEnM6xPodJvr++wdh5FUuURH419pjLNjzvbM
1bAmHukN/MYWm3PDIYChpm4w8IU8IAf4/+kb2ivesQmoTe/VWDu1ba5l0DTJX3hf
xl/UpVt5917XhpsEiiv30FPHXpoCO3BbTG67h/yIshLNIusr836BFgLkFKbPiU1h
mvmcXMKhjivL/IxW22DIVTGmrLxHgv6SjrClt3sQ7kqniFsY6Q9YCZiuWgahKsUq
5u3EsZj3TVKJNm9sB4iS3LGU1b2qxqMgQerJMo9eGGzl/M4K0ostsASMnPBv8C97
O39NZV0KYbnhhweVyBwFVyx+xTCklA+upF9cYxYX5hb9Ayvf64zem68kCqy/Be0s
NyVIcpFwCQXI5Xb/IEiHjOQFQjuhTEQ0xGQYGfmINrUBpyl3r1PYaZKM95ZQslqN
30lIihKeVFzgeNV4tiRgy7VNzhP5WsLBmAO0sr71VcFgqj7VSWNJFer7uhZc3pi7
COXe/a4Zw8iHBIA4m1wqUzpzdUbhR8tBrMYrw/gsOpxxuNwNwqF0O5LfMgA5VPF2
D8z+R0i/dWLbETI8ee7n+zN8okbxzq2NQA4b7Qn8WRYMmmhr0n6CPsQyxYbfmkIb
uMIXCAqyCh5gSDyvPcLZ+Zo39LPmlaQ3MG9XkC+eGOTMHNcdXrk2zxdbB1E1JtSW
czUahI6anHdhB+MKHnpHvzRaArYqcKEvQ2Zp3hYSuM/pWxK6yYlSPj9VSLw3iiSl
8q08BB86noxKhD2zEvtjR1HyX8yKlJOyOWamyuEl3wBjrBxi+rOPnjFJSg0JMfhA
1kRvsthLnb6DdoS2uPHbTribkm3q19skCGFWR/s6y6YuOvz8BL8GAVvgImWaZ0Gw
E0Rqkc6ARljIf6LnZYiX7/28edsC6mSro03gJm2iRzyKgt4BajGmSHtVM3enwp92
ybHIdr6JzD4Eo2OlNkoXi6s2pSHnNV1azeh+K2xWFQcGw/w61NSvauvf5weLZj++
XHax87si9WSCy/WK97NSnyvLW08mR0HIutV6/OxhU0edpbGor6YIuDKjaMIxJGWd
c5JVCJ7810BEYb8iboRTTJWasuArpkaQOQcFDCD+ObDJQM3205JkCPNqlvPFyB9k
O1jc8LoXkfg5TlkeaUu9kU9U7UmuLm4BW1lTzhmMbhmKNN4gIncEuqyWCzmjf3Ky
EQiXV9cdvOS/5VBfVmZfaeVGVdb9qPPpaxVquYzxbdN9fuYoLjrl3o3cCzNcb2+p
51ofoQFqxKyLVxNkHitDWzMsrjXE3JhleB7pZ44k+rNiKxqcOCAVymvOSpuBHQlO
pYsQ+bmBAiVHQqips5QTeJWpf/L4KANx+7Ae8edLkHmvF4P79+iWY6SB2oyXF6z3
JX7OAq199t7g7p2WQC+2SXwXv01Z3+Bklu37a1ApQvTJxtW7XMy8wCNqSwTqUycC
G0jxbRsq/MemlqO9skCuqo4lV61jrfSAnpSfkLm2Gwn2F9bAXeXbuZY5ykNHez2D
CUNcTyaRlX/RvLOnQSrrxNnc574ducdtS/XMe8By8onFdzJGpa9EoDC/otH81yv/
FxfddeirVU43UquvOWoXlc+VXMjnE94GUfLNo+ZQ1+SUOuA+EeoQAvKV4hsnIgzZ
SMMfEi3SbmEoZF1VnhXxPzs87En0GAPdWTsZe5UQZGBQmOsez2E9RsCabDn6/5vb
n6JDVDnfJoSGWhch47NNA3U5ezCMU/en1NzwLCJfItHgoyKDF4L2braEpgQ2sG1q
qxOkonD2WryuEU1ox1lNBm9z4lNjrNoWL6/tFgoPw5ztXRyGZ7qNHc6Vfr20AN5j
b1IdVeOdnxaybXn71LQtJcGAUzf/OVS4RfTM53lInC+mEMI+oqjEo5yci17OPehO
AxJ8keRfHuuRu01DcnMWsY+c92ckV0MgAtx0y1fRqWanGKBhaj/dUoQQa9sAWxlo
CjFs3NZQZFQSuuNOsgTDjuK0o+aJxbOH4uO2C/n+l5lWrA37Ix1Nr8ZIcjEtBdaa
AeH7yXjUiHtiVhGy2iO5Ae7KlabRgLZTNIhX+TEQKkYgTQ5Zc69J4Q9me2TCiDTs
+b9QHflKeRcTP0LY/7z+YiEg/+KpFAEdFMLwKR107esUdZui1YGNp+nfrSoh8TPb
xh1Ik1ns8h/Q95SkU7dZ0UReZGfkWc3sNMp5OMlD5p0oD7XDmFV7ePjcKiqttniB
WvB32PNw7D5kVTvM/nosSHeQOnEnEXYlkj3Lv5eJLGdPtXsDv6POQOFRpq1JMO48
ZrDKORIndW97WfxJf8GsA72B7qc1TiuHS2+qesQ/YuKR95kIQ+wmHs42z2Ony7OU
4fGqYamxMykKmejKsjtMVgz6CKjC/wEwZ5ECOyUC+P5wLDrhVbY8e4UzE56MzI5l
kzv946KXKl2CUVhRKqEDdj0LQHc6PSe+vnjCp/cYFTPZ1gywTUO1+8wHPq/W+nad
0TARZwHQMhVGWqe8ylCqH0d1ke5kMuteKnEEgbMuUCyoNyG8vqRK2+yc9bStOeNj
HyP0zKCKX7blfGTJIiHAwW16uRly7WJ4gRUeiF6L9b7IW5zQrWyKgqCSndjFlvFR
wdWVbZY845pg1YY00dLPib2gz9bls1y8D8rZWBV89S1TxQ9DHb14zBBx68QyieQj
HCIkaYS3eOuz+v4H/xCIBxEvOoEVedlr5w08wCB3632Vh5bucnvcZL5u4TBViPGJ
S4jRQAQuBWeZ1Vb3HUHuB0JqJDi5MvWDzmzsOdcMuyRy4HzbPZo9TdnbFBNa5S46
fpZwVlvJZTBITZjdO7QQv+36WlfXUEtUGO6x8/icdVcn1wTmGwesgD4Sm7Q/YJ+4
c7eVxEYFQj4P9+h1OtrEWdLztM/mF/dQ4w7i/8+OfyjQmy/pC/6jlNwKbVjXwE+2
UPaPBpJ3KT2Kl72OgPiXufdG0ksx1PUsgd8Mtyu1LcSliwSaWZmm1ZnkrLFH3g6S
B/2LKyAepbkgTjt5KC97A5jQ7vBE2wf44a0BD8QepynuDGoi4HM72RZJEEc32IGz
mdKvb6NSb0NNgPEkn1fd3szUiZgwAPKXGDcNH2mKzQ4tvd0hbQgZR82FtX+u359d
qniqCSo+joT+2CzRgNV1otIgl6BAf8E118dZiDX+2vmKUiNIsSGzc/ugc5xgiOh2
FpRWcrlRwL9bgtII0n0ICcKiW2ptogh0BLPlfsPSXNwyFIfvDcrtiTZEDyJquDBB
5rT8tlLhcYHpiLgRAHgkb/dZY1FnQ4sy4Y/ASBwatAFCKjv01tFPS7Kz9z/yTkJH
YkQd0nk1CK38bCQRBWXUrezQ/yvj+cQIuT9NQwDF8kRoC/CNnsz8+Mnc+Wp7Sd1G
c3+bo91Cfoi2ij9eWiraAXPGAQB08WpCi3cv8pb9Hwt50q4pL0cJCZMe7HLfMIxd
NcjQ9wl17S3xvm26l+M19s4mH/jNZ7/Fpy+HO0rIGQ7mJxdcTC/4q85eCgN3VjXw
6zGt3zLn2lqIeyqnce580hrhO+If+IhPZYwPo2rdvI7NUfB3803feionlp+mKcpM
9tRgBE/HNOwP2l6E6AcOuyaoVqrnAsq9i3YRs0hbt6hTpLQfxKeTYe8Fb1QobPQ4
A+v14fjDZPb4G7pSzWRhAsdPbpXELuXJeLSizOSd9aZ/pxM1TDNfNrcRnH6TkcN4
VKdLXq6/Kb+Mvo66u0vhWLkXSqMD+AVvpPAgXSod2Bk88Zhhftso5XLWO2/InwCJ
ArOIkKK0HokZhlI+ecKKu+U8ifpOOSqvRALXnWULrdaZCZZkmpV7xllTFVS27883
PtFz1+pnZvBLQduqsY7ShdEUdaB4OLGEFPc/xHLp29GKJK/MC8RiTJL9TUDkAs/9
cbV0FDedVM5a0AzulqRSDjrCpHB82VdsOx0GZcYUFHg0ILw1OxRdy6UmDhHOA7nc
JrJGzTJoq3vGx4N5sDP59AUhFJh7E3uD2ZJoE/uoIVJPBYcA0as9Qmc3nqqhA04Y
BxczCfermzZhtEHHEbH5eM9phsRCbxIJuhpfmVlr5xrpavhyj+0p7BPVfouQkUyA
wi/gG2suTzs22UXzitG8ciRYNK4R4Dgv8bJIt1XwSZPBMU8dOPNSmyvLyWGcg4VQ
88qFlQCX9HWBGhCO7rfn5r1J0Vm1TQ2h6cazEwQCjwkxKq/kAHC6pfCW4NSoCXE+
8zXOi4b5Qjr6RQugSvkHqV/FyFc5Mmjc6BWmZZTmzOJ2mdh+M0+f/1M2pfE36sOn
Xywl2GhY40+4tXycZRBUCh7maP2poGaOgtNVunOg3AcUQLmGjqnmP6UAZyH7LuzT
BD5aQ4/Jx4uC1YkL4hS3mYXRS+8xRbpnVKdQNTfeS7H8v2tButrwlhZsMRevuidm
6k5cH2LEaJjKTtnr5Ci+G8JWUmWxttHC5sdgziQbo6qa39yKfCb3hPCfj4i5ptkt
d0McXBO8NGc9Zk6jNNm6QMdFtbGZa0NCOUc+j88/bMgV+stJA+u2tfOzns+DNRvb
bpoA8iCTzBd67hsUxUbqhXfK4pwe8qjKDzdPyjfUZHbIWqarTlIIo6X+e/44fABr
tgx1ylYWQFYkb0Uqk+3isxTe2YhJRORkKvNxrXvAH3C9UucM6VAkroBscF+NwzUl
qvkfVjIY0dzFsui8XEfWxURGaX6Sy5eYXGBMlnIiVg9aPbRyPGs8Gzy09ueER2tn
/5Cv+DmA/KamETTUtRvLHlGREMtVV1LcZEYWvIPte40fzm5n2vKbMarAFmAHQB6T
vfo0K2/vF3UHf0H+UWt89z0A2lR1E0XRyOtwFHdCT8RKtCPHSbwL2KDZWxgzM3bD
KT3Be9+zvDKbN6ktXl0Yw/1VQgS8D6F/Bm+ddQlocVopVkc7sa58nnLoZY70FEdj
QPQOMIEfRw+sPL1jA+QKM7WiDRs8yCNV1u79i3Pv7aVE3XdjE2xVGJA6/AeUB1dC
qfCBVEBgeVNv3jIeoI4aoUB9bfT7bWhNjSlhl/Xe1lbbeM16FqUqq3OHwN77JsOX
3euoYZjdXdtcClZ76FkBqfhYjd1b3DRdd5NRz/hmWX1y2m7LkjkkVsqmbo6rU4Pn
SQbx4kUdsxPnenasV6msB39keq7phsqzekxG0UkrzL3sltLq1ybs65vp5qQshdtJ
SqCMm3csRCUXS1Be2itfGt6Ttzx2Kj5A3oTZCgKAAJcWpEnubj4AT9jcWKnGQXLB
xun4i+0oFOtsh/0cXwPVbIjtQ7J59+G9B3G86UFFFIjEv8UGw6Tu2gPTiWPcl4NI
CKFE6msY5fhSDQZRNJzcjErmnD4wZnCDJtvx5YOrjq2YMGYtwtTi/cjMOuAqQiGH
lKYRYhT/5qNL/0PPyOU4KhdfoS+TbaOlqJX9+QgToNQpH5c6pf5bk1jkOXM0g4fz
8mc9WHyqToHTl/1y4Pu/6e5nSuvIx0VNMGccmaqZb03QfAveoT1iQQmwzQqMPMhR
pFYL3kHEMhiALIqkWSUswYph7tXomjSzjsy0wxsmh7Stfd6Ju4oo6yYYlfABp+Aw
dacI6yfGDgVksc5S+jxONyg7ofpRnmbfDRwSm2bTH4nG653n50AGndHGU1VhB6+Y
KrHMb26RE3o5Ugfn1X7wQr+Y+HqmcpdN38aPL5wcbrULOsY6533uupzpU6EcaNzL
whbfnRoH9yfksdxBHrAYMRPpyLy2+A5QBK/T2aEeFTQa+/fhGt3zxowGvQD5Mtv4
NdYE+bwDhO/FckLJ7yN1MiU+kQ+rgiImI0jQNPfPJpt0rBSips6KRyBUAB0W9o06
EoZIPfLJYZwpfcklNjEhFfzGleGrM4mUvO0IsW5NbIe5qVcDS8QHv7ZR7YEjDYBi
Ye1/f4YWOldaoR2Qrh+9B+oVSYWtS2o8w2rA+nCZaf4wgyzq6BJExPZ0tw2vjap5
JaQD82IhWOGOVh+vZS76L5H8q/quFUGe3fYSperz9KnMtRLD0vK8832PzR/zsNcM
/Bjwm8EzBA9auGwzOiVmsnlgiErKz+y5DafHytAt9cEYpZSalzyL2jkMcNCdqZt+
bhy4mr02auCuUTq/Aw55DfphswA/OTp+CD1H3/w7YIl7L3jX9zy1N+4BExdME2GP
SExGsiy7STg8/36Ue7CCIzC8ofrfVq9nDwp2y4Z6wMfLXVhYDYTrLNV6rfOkTZXa
U75OPgScndZLg0jIVhfWDq2d9l7BW0A01zMbEpM+MJ5hoObcqMMWZWOG+1Q9JT1/
yn7iggvDrs0IFLhbWkieA9XvDQIoO8zGk6qCbnTv7g93nthuEJjG/BNTZ6xcJ3ZV
V6D7UW0EHJyBAEbPaoapUcnu4cwjxkhzsNZrU7Z11WXDs3KZjVEdDs1owH57cmcW
4w4+n2w6v0M0Rs89gGqjnPvUqcrgKch/AxicUbdNz4Hdle5XKSyR1Fi83EsNgTqt
RDZx8FwhaGES1J2IOdYQiGqXN2UKGPqZCCjg170QvNVn8i6ivLRT2SGMreAIt28Z
0mXhOSGdZOSsDvFSakAFwoqyPqDTiU/dvH/P2via/5jKANRBHmIaullL32m7FaIh
0/iSLR1VuFAqwnoj1H2BP04YLKvo6HjgGy5+vxrxd7BAx2SWC25oqEcqrn8rQy1C
82feE/MSBWOjna1PIgVbJ9GnisXK3sKDQvEafTCZzlSMdR0N5YO+xtBW7xa/nNda
eF/ujUHAf89Wf3+jOX2PwQASIfSDOEYUBGb6L66RxRaqaz7UeuJKZfO+Yv6cfm7m
qDMmKH5CQptNbaM2LmoNKJuXfEtb6uPBEaDcKoJgirXJfSY81l9Ww9QUPL5e4XpD
DfkV5gXgYxtbTsgWbhwEYVKA/czxo1FVHrhWE+sjRUQZPlFTD4TdpIu63NUghSXn
1VZ1F7C6rJBxZs53392dEUZxfy8q3KmdF6I/nIj0Oequr98/ZxAath1L8WcTwttd
pYCGBCq+9+2BzFtboRXY6owwxMkXrgAreMmDxs6iJa82BbZPqaFjfw9Lk78mC9tZ
MTs34GNihMFsoZ7elku41bVacgJVLN/11OkhtSj3UJUthlhHgNm3JPJ+Nwon7hYr
FISB//bHNBHeMAaY1IfXxLvKUgDrbUfvOKNjvG4bW/pHex8u6X0aLp474Pluh98D
owHCLvTiecL3I7Nzf/WDB0WU5UqWfrak+0dM9VdkXX+EtvajIWQbSrMAvF97bjWV
YauaJ+GbjtRYkl+fdfJhcrT04yx2fMZZfvQsjwq66Op5r6VmXsSH6PjzhkM9Fydi
ldYHIqd4+oduf3dalL2ZhzmiKzMevpNXe2IsWVPYx1V0BeNZO2Vq43RPsKdqp8Lk
MbwrIy7nZFcqQSVG1HBnL6ObwvL/CL7MkgyzbAwsgfoCFa9m//LdGMDo8yWCJTk3
rLMHt6QXWo9MpYtm7jLioJufMQ8rJO+9PKGbX1KN7Ro5Lz0ZBKjX/5O99wo3o8g9
j3ws3IhqMF9A4dMdSGrceNpSQ+htQInlRcZ78QgxNQvwinegbEaXdwFEwikykFOY
IgeKMHmJxoKuNxiEWs23HBV9/gpYphzFdpKeeVlaKxyUkw27t9tisVuV++3iCWgx
JO+xF7YnVXQnOQ5p2XbYYFvfGuJWurTL3htgxZaumXvnMqt9PzEU+80uaNEb09aw
liW5chsQPPDLLKzStuawav/YmUwzQVjLndIDeIzquCtdZ9p2NJUDbdHrP20kad/y
b4bOsndPfKxvCOyMK2LvfHpgVDjLku0ls2xHNxgXJqI4elgILjxP44YmUgxrt+Ba
JIW5T+YEendyaihs+8PEYqFV9ikC5IxjKuNeVP6xJhBrN/SUtNffZszxtVKaRrp7
40ZY0Rbx9e48KWM4nc0U9g/uwrFGUnF/hK4e6AQ3UDYrBbX+kdaMsyBPGzHVzqE2
9sQc4eNZvO+Haozn71BYKLO2tQ2Vxic+/CR5dLgNpFt42c1Aix54sH6SjmaQgMt3
PocrGVRpCE/I6CWS2sguqDBrZdm9lflSMA8fRTIhH+8HX0LT9+cAkufHa3lCTJbk
zzVepW2tV0LHEWotvdrZ19Ay6FBSSlyZWBL9ZR1FjxXiK+rM2qje6D54Z2jxmwS2
FOOsC0yzgHxAZ+QOVEimtCa7KLOAVfG70/vVWi/7wIpWQZkdI8l7T4STht1vHzjC
0jylK9Ni6/I8xguPaRzoOW3Ob9twmko6v9J/dwPNIM1fCGQBDyiiehTkLzC4LF+Y
sKRz0XNQbC4PMG4l/pGixqcP2t8awuuWKUfPOXDKZ8nKuqmujObz/0WeNw5W5fqk
1FrkJS+sa9xjrra/Up9ncGs0CJ7xfBA76t+Jp+MmB32wZukoba4NsiBeaXIHd1a6
HWcuCR7wtLxejWC2c2SGSsLA5vu+/NZgAuQ52FHRPSx8kJu6suUGltw6TT1OB3zf
TeflOtvRS0oYOxwx0/xpE+munxxIBLpSUpEEwUpdTzIVjX2Y5ZEtm+JsMp2IuX7Q
KV7kJQHwho6u910UvA8JEFxkrJEs3iw0OJXciI5dRgN4tQe3rC4wPWfnTsqvr/xX
WdWaGv/eZjXKCQtxmoervOGUAi8N5GKESUBUKyFb8/hX/gA/LKPrTxsumT4vSnEk
Um249LTI1wjrffPi7e9csK1jxThMr+7Togw+3rXuwTxD6qvN1m41ufcOFC4XWU8/
eIo4lVZ4sD/a8PZtXAiiCVBBhyIv6wosDEoDguzcHqo+bFoWxIDLv0twFqprTwAq
ul6bviSRSa147D/rv0kuF/yCFvfV+mY7lOz7U5okozWJVFcjcqfQm2Xrw3kDuoQO
UGa6T8IaEZ+HgpZUy2ObZC79VRfrXcHHVNx6jgeUyhAOQtM+V5NzQiNDKK56zXng
hG3/YP8UhdAg68oTtRhyUC7ED3FoRzDNEHzNjrqNcNv0mIoLsO6bzl+FJIjH5YmG
61CeQyn6AmbHtBjW0uapoObCzH9uZX2lQV6Im6yHJlePS1ro4U+D+zDiYjPxxk8x
U+vUCRiKgML95KwQaZPO6s5xPMlHtyXHKXks26Etf+sYbh1a2ge41nZRO4WWErZ0
g/k52Zd+j9kdqHDVanFThtZ9M9UKo0ppxdKSnw4tNztb/tB0+64zVW20RJxCoaEB
uWBzn0g8TjEObl6fe6EKhdzosBRYkM+mds9YyXKMxPvlVwKDqGyfkbuaIKpmZKLn
qFdJO+9OS12nG67jM0E2q4uUEJSrYZUoa/XDwftfKoK6CVeQzBQgk5W7so/uuMLj
dXNRw5Q/kEGU2StwfvFePfbKprzoy8SaUDU8lZ2fEThSExup3a5IhZCmWMz6JQJU
4GX0/z/RXYbyTBnnOd8QOfhM/TlJ56vYvlF2tN2EGkpxenScMdQDZylPnASZ7Xe6
MVX+/3sRZFk/4gIeb375VEAVYaMwiuwGyvnvd3WAevxpwZTwWFRWAffTzxY986gO
pMgWYQCTVXLGEsgMp5Vb8rggUYRodUiyypygQ974F82ijvMq3Xg55ckbCCGI0z+3
82sxLt3ws2Mm6BHvxtNdl77nNYpuBQqy5spV62Z/KAAiUChOhGaRMQe3TXdXF2+E
FawMui9YDywLuPGE3oJfIegQ/Qg7HcYGzHQENcQBcIo1fQeMB3PgDtSh9rIxLCeb
/IG+nkzOngXlwHXlF6SbpAfCdTeZr1ZkGVwGB+CO75en7u0yCcweuj1p8hRbtkpb
42oU8qRosQKXLherz9HdhU9RiFizCjgn29jg+Klk1Z5AfrXohgoZuXYjjwvcal5N
rkIP7MepgV+j4oTpm2S+p9ole8+6s+dJ0L9Ce1zCIxD2QPq6M11cWv25BQ1WStRL
NrPheWXLBh83g+bVP1yd2HaaVyhK+19Np7dHLojIDXZrIAtiZJusc5Ayje1Rxh0o
ml4zUAMxQXAiN5cXJTYRYKC5IhX7NVaxxKrn0htLL41G3UztR6hC0+joVZ4yBO6r
aXfCt5cU0LPWacIfcUH65aSsFLYL4whFL4ZGPumfVXWAiMDLgeEvwEnrUOmMPED4
/8bwl096O6cmkB3x6KFsbVIYUrHvK4tTtNmgkfuyYMnIjULF4SWYngoDT+1X61j0
XkwgrKDmtYCZkgADhkmAVLorbzGeiEs34sVn93Azcoc1uNQLSl9dLFcr2eFWbNFy
4f34IueGq4APAX11+Xgr6njhpuzFJe4WdEiP4cMlVhbHttptJ0LgETz6EWsfhQSS
rvSN861HvTWQoCMigYyHRPCYYTkugYpo2793sYRMnhsYG4SFdaT+c2yHSlSrHWfl
QsWgGzRB0cgZxmkf65fUq5Gh7gWZzHNSW5VryE6PCFNCVDNCR3C+fu/MoruenYi+
sMQIAp7H5VGk4hMjFxHHV7PKBv2bxObAc5vREt7jzkW6iH8d4V5mCAPKf/y2/RHT
5ku34J79fTL8wlUwaA0/+dtZmEXEG2DDjzl9WMuYjL561R5Q4isSTC1uW+g79bhO
l5xcZylhBpUanKRHIHptojxPexUvcUwitxh5zkIAsI48f9qop0P1Wby1eH7Pg3e3
ODRiOJ15QKDrda8adgdsHoF4FBasWZU8dmAUXRplwxq25n/RwpQp1Azvo6Rhnlec
+TkFrEEdmhTJIBPI4501Ua8UrEVYAUSflx6CXyMhAYsZT+KdkjPf4o0lGbzztLGF
YsE6Vonte13dbSWm+XOhsRK+1f686jsopXi5WarO9jYk85WVqn2y2jrRrC+1SGOy
mssir9QTeAh5SfFrr7pHLCWayPRkVtmEqZ8+E7XGf8LVUjC3lOzoVSjXFboVheHE
8H7ZM3oCywJzj3iznt/Bkh5wQdAbWQMb+1iK1eF5T5MeDBkrzdqMolv3fO86DCyE
Kskc8N75jLYaCpph1/fY0VQDXPTxy8XgFfFFZD3+D1LxXZDcg6+EjQ698WPiFnGe
di4Z7OYK5/dsDPD1HnEWd5eXZO/TwB3q42MQUYQc+8rPNdeVqgerozAb4WvyXX15
SKmZP4ZYoxe3VHdre8JdPDQS8Vwa+elCN6xBlcNtP+rM9w4UTpjj37Ha8zkDSefz
mHY1h8Fjg+yKtPcqB3aQPdGLjXQtj+n6p4eMf5rCFzXhgBF/xXEs2My3DX5GIWqz
YXUQA+CIvfWbrADs/BkggaDAdZZQowgzz+DJAh24oX9z3pluQ6NhAhZSrYdNfeVq
aUeGJkk2+wPMpOdByYGZM8Fsnf4b6qkkoZ94EbS4iJTchfsu3CM4aCUYqt5kgNXD
1GAx3awUl/WO7uyKPp7aRvOMv/+KUAqar6q0NQxE4k/Us0W0QPxvs+G4E7ORQjq2
/AIq8Bt28K3Azrp2hR+u25r3BRHXvStB+AmKaQ8TINkCyTx+QuR+/EltYJIADzmH
oqIqarRtZQPcA7Javl66YXxJcaldjJEYacHMySWn1QNQjKb0RIPmVd98YSfHRcG/
v4+PkDVez36yQXsop4Qwh0SnLR709rpHfUdK3D8QooAHO8f3d5JiV5540Y2GWUE4
IwE+6ar4AiKTQTf8mrcWCy5vJ4mB78wLA7QztpYblgz+LpI5sjsPZnoc4+wBYwC0
FgWtzleeAXlxVrenPnU04MnmmG5wXippxck3KhJ9kwNuzDvP4GkokXOC1Z/q0rgd
IwbJfF+1WSxhc0doda9efG3PRFiKO2jyRP4EQpSzvhwWf5gS414z4NGnihl5R/fO
dEKwjlzY2VPbgnpqROHaclHj9x1UqKhP9X2p8HDKJqFOVDB5+Ns2B6uZ5IqM4BWA
zY0tuutUSZVAEl12xQYFfn+q7/IVPoY8fNCyAH8Csviwf1lv6dE2tHNPwnVZtwRh
Pyfqhs7zrlZyAMlm5P4Um3DCYe2VnCVbN28XBlH7xhWRkftS/WTZlp8dYVl9jVvC
0RBUJ1mJQ6imr+6HTyOrMOlvDiA5XYniBUHVLcuf0xqrqZmQ0QfL8zLVDL7yGIZd
cQCNnn6QfJ2Bym8kjQTqIrXozRAECsCAU6VRwLbGPvQ+674ajLiFz5WQpTlhXQmI
VZDcW4M5eAt6E+BsZ7ux2No0JEVXs+zz96eYU2/Ye1VkXN6/2hcwPiyHtnnHQULp
vAXuKsA62XYVafzlWZyax+ZwSupJY234YjEesyjbqbwBUklBshj6KTc7oTHSXygk
TQ5bvR/lu+If2zgwhj2KuzRk9XXHnrHSIQBN7JZ9/n8XjKk5pf/bBtg0+hwrv2Ai
E+/sxRzp8fO92pYuFwG9V6WJnCsM+mtLLMdP3AM6eKATvtx1huyDwfXJ9vtQ7H3e
j0rt2x5wfBe/hyw5bw7TAwOHc83z096LSjgsckHhVj9tncKIge0vDlo8yRxOH0kf
e1+ARBdiOzYjhDghmzv7t7i3NomNtpbdsEu1dQk8yDO3K3fx8sWkK9yAI/ppeSIA
AF6NkmkaEC+Q4D7ceq7ybsZ9MQy5CI2xkJ2FsF87NTn7XTbOBira7QfvrdM7F+k2
54FUJrF5jXmgAKhVwF7Sff7kjM4dBvpeDU+p5r8eQbd2b8g8lHwqD+wC1vY8fglz
OpfCwfPRuwMIMymhS0blGuit85hbGiWl1pDmUDax6giZQ5Ani1/fBqkJXgnFCoVR
mx3QfiYCqu8aGusoIatpoi4ZmrYCixqYN/wUR/HAVMmC7dgXrcBz7ZTkNotYc37P
i6dMwwreevMVsMt3h8YIzfc/HLtnbNrFzPh3TtMreRyhlxJUXL+O41v9RnKuYodi
6yoOjdmWmkNIsQoG/e2oj0JY1/IlwgWTvFzt1Bch89kfUtSkxbKs7eGvTs+SjryA
4FIEQsi5rLHJ7Qqxbf4ftbUySsDsvUXWcsnHStNP48/dGeNR5k3ubyi4DHpVTzDi
uUqoS2zPWRYkc6N01HBiFI5NX2YH3WYfEKbImqBT8bQ1F9enToL3drBzTeHa82Ju
rL7pSd+N6Nj3ZCeXuMEOkDoPyxTSSwBRL92UfO6caBB4a8pPOOteS/Uhj90vnP10
XHNSh3tKtV16SmXR2v+rZCmWoVMbwHyo8PZq3YtXKoXiEo4zfkp+9YXk2TCaT4AD
JwcOcGMEqu9sXkUP6uPMMmW2Ai1TP7ZDNQQQWyEVZD5f4SerOnKwLsb+joqMphEp
SlzQfc04w+4TyNejYHjdTYoTEwcEjKvZCCWENVq+Ky9l86O9ErlAhQm1o0wVP4lJ
1w98Zm0q8jnyCQ6D0Iqdv8DBvnnaNMzKnxj9YdwikFAP/derDqIOJR+xcDaF+YCi
faJKR52ccwxZepjUj6pDJ9R3bz2tyzzWUBGpuuoo/EhAaMnjIqXN7FpSyHA+53qn
YlRfMqOCMY4/aYGQRJ7jgZ8D1Umu/v0fpJTPHt94wW32YgHEGihfgMicTihDuEYP
r5agzvhlOX/f+pGyncwOGuef83JsrnZpS/iZoljx408c0yg6LMxl51NbBp7OmR+U
9aqeOLDbqnd6MKizYmEv302irWMpejWIyvvo1kzTayu2/t+YySUTfszYoatieilA
T7Q0RbBbJVY7qxnZ4Co1eKKONWc2o3amGHx97WT6gVlGeX9o43PGnxeLKuZiIthg
nfPxs2/8G902YtZL/YOTwRBHNVGbtH7ydJST5uqyBIF+5AxS7Dbv/aR0lph9OsW+
2FKMzkwKJ4QqwJwjkVni38V/O3KISHMkXY1x0KaTDhHq5UXEi6bYDS3mS5N6RiDS
bPpIrAVbqcn7X9rvU+YDAwK9El5dFgrh2Y4i/bfif7L/WPs5oAlwfznlkzQmTEFb
WkQyfttTmitaL5TqVVAXKVlwn1cPGEohs0koA1DXqZ/riMKPVsqbBMbZHuuKKgF0
gUeI3PDlOtiMIYolIHN95AchqHAt4jX1WMLNUk81sr06Hq9ymGxO+wFZuovJIWAu
umY3L1sjFIONsG7HWZWIaYHAim5HcZp4DdWn4r220J2LjQXoUkMiHR77D474mMSX
imiXWmIkhHnp02/fqlCG+fKmol9MCOP8BhR89AB4LWJyQdAQdH3mZKuvkl/84s1B
SvdW8+PhtjztfjJ/7cHIVB2vKTeyoHU74yxcfK5iDUzM/2Q5mZ9ZyIzu4FodBBk0
n+tC25TqMoETC/IpBVQP/hohEegipM6SjGd8znuFtrICrgrMIi/+MZDisPGSHLJe
meZUZNGc5fkTHlJ2igm7tJw/gm0hKiZ9xa7wjXrPsOJ3NhtifjQf8jw/5fOBJBCZ
oF72J0j+fmnzrAQHhPMsV3lFP16s1FibCxGW6/b2ofU=
`protect end_protected
