-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
A+jXZ/E+5hN1Qq7JhykPwHSVyO8L9aL3ZuRrsuHg5iKsTqor8LaTvI0G9xmT2iEl
Qb58oVGbyeXHR88qDpXhST0pmaz8r6i66kp3aq9Dgs2DuKw4CzMywfOl31h1MXAs
R8XPJ0z1RAN+sSnalWsFzLK4OHrAKF7OsDHncAGZcK4SNLAPaJIaOA==
--pragma protect end_key_block
--pragma protect digest_block
oU/Cfa71++bTpJAsBbVqHHaGzEk=
--pragma protect end_digest_block
--pragma protect data_block
yrvciGPX8uXBDraOkLO6uvCVk63htG9+9xxfghtlzhQjAwtNJHfnjpWjwtZF83Ic
NfMs7rSChIbx+/pVFWHwzoiJnv+sD9Z0XaWYFVvIngqsPLU33D8sdOge9u8SlsKM
oFsVX65hjB4tLLZ2zlAr4l7FWv+zbqjxxNbiYKzFGib4OGDohMXkI54SIVxSGzJC
e3y5vY0t4vxy24yPSi8rR4bNw/dgQQRRLp9x2TFLWHh2UUBt+YpYNDxOlfaEfsbe
2keYnrNjqqN6HUO2B917o0QUW1H4yI5dGZM1mMsk8np37pibqadoJ3njJm+lpBQM
eDSlKYjcq94FyP6ihHc+qjZh1NIwquua2cCYk9HHzkvbKNc6hQuk+sdZgg6oEdc/
D+mztKrL7NSyhTlruMP7WPaVfxrlI1EFjKJp1SX4GoxQ2SkPePvHxedZmRW0xnd7
r0Tyqvt3f3ceZeKW5tOiZIykTXtiIHCahzKpL4kXGJ/y+CczkrkBqLguyQPeoumx
W7RlrtfwvZ/IsIKW+s+C1LEHeDwn1bRKnO9RgtzcyeCqZhs8fjFxnKm1VEpfJg8w
wLA7UBlHwIQVZyurPShAY1IetvN/Oez1Zs9JOeC8KIWIT1AumpN5tj1esgPtC0r5
ifpU+MLMV752wD1pyXpZOiakdq0hRtTUI93lO4dfzisWUGhPNkwqnR8BVXue1N5r
7aWPZg+U9jazXsx0RvHAwMYVjten7EPOurzMV6a0hUMzm4E9JSM9/PO5dutTv47b
dMDrHu96jF77pVjHVmi/j+xV9WCeHKmqiHz1ed1UMvM3MKftF1Ug55/MCRKI9ibG
VLGkokY/1HP/HRnXHFuuMpr4rqK7RS5TodzfWO/CLaJoKREqc/GoHiM9Nr92D8VZ
KbepKSlGtiJDcKjhm5MUNjj47N+ukFlFTgjcjHXoukE9ia+eQiAIgWuhtXCP8L3u
u/dvCT+DHf88Gor6mG+wqOGK1y0sJ/varYZtWb4+MwPyHPvbHfwU2gJW/gFFXrps
YCZtSSoO8JPGuxk10JYeubx7SHy4OkbzcR+DR5UwMMybOadfoJ6+C4jHv0/ZopF8
BeTk8IHjSkZS0D81Z+3SzmJq+66vQ3gy5e2U5RhqF+xAxu/uiqaBXtMPZmuURGq5
h0LkkBa5+NppUbMXhGfUDQcxYejnsuolnwyZstCPWiz/93oEDsMrobz5Tr7Mc2rv
6eyQtdBCLntNtZ8YOT8AbB4vCYtDscx0WzwHWfGRD7DsNGCq77VD3lIJW8PEcr2k
b9PMhar0JSSDY4QylVdZgrZkk29Ov20YM5hKK5N5sfoHQ5GkhuvWq+riKLFaemqP
rarJFVr+7IFpgGJE6qa4CLLy4xebA/2fodMlH0sXYCFAfT2+65/Ea5+ddwFgs/L6
6KKQn3qHNYosR/ey3fu43HJqqNfQlKup4vNj77Xx+DfyXkg+4HcJz9DP/OvW84dy
Q6fJKIa276cUTngPdTh5am0DPEoTm1e8YXbV1yAWJ8oeGnWln1dBaIJe9pkMwMAK
a+Y6q/24y5wIyE6baM2pB3OsXVwf/JlhNM90IjuD9imS7/BnStjQMhU9+QdDh+Yv
tYmDR089UtudP6hBYmbEpPJ34Pa+t0VO3lkuSKYS8vVKsNN8KOFdXHap4ey82W+O
fvRz1A/HfvDPQ78T8tLLQHqiTK2CWfjX5SgKsM4EiPFIFxwBzI4RsqgtZVyB4wIG
oVk/QXZu+JSRMUCnCzhYY643YYn70D39IeG8d032ME0f/bDw6QhCUmLv4+Fpee38
uxicHsLKlbxaWhlwQH5QSPYW7QKmKR0mXkmSTgIgiRAz7F4Lczk6uLV5PnkIBT3U
BikdqXoHpuR2CivBWwOyrkQdaEy0aDN08syulcLebiNh24pTcDAudju1oYRUHpvK
ikiHQ+XsFSbR2fKrMvstUCV3nj3lHefGzZ54/CuqpfQBS01kCewjv5tkgEffOoeA
AMx/OFrZDBHW0uouTxqleEg6JqPnQXfa96wr9VbypTdf/1gucmEeGh1gCh5P7BDc
0ZH+zYxp7t0Uwbgtf9LX24rNxyNQZp73tkT5746rf80fnzbFlDhKNjOSZMkGYRBq
Mp9L9WwqDrZqHye8CQiKecL3guB5lDo7QSfmUsQUDXgFzz8YMVx/0CK/0ZoSrV/k
YgP1jRTDcj84MxFYJb3FiLFx+ZD8/Mct6Xbs0KeTOW3jHtjWzsMEzjk8IChkC18Q
kqqmkrXRJobGHuBP4uZ/5lyvtx+LFxRlsQKJ2A0p2zCWW6oBRSp2V1ESPo5Ii1gU
cca8Mb8DgrNLRC2jwrAz2pAmOS0KuX484RJ3zkm6ahdm3W75TK59a7uMvzi2xLlO
Fk3W0u2aHTeVtiwyjpyQZLeJnW9vP/PRXaRZlNVpHH6hBIELDwsT4qJB/qhm22cP
QlKB2zBrVC0S8FeGG+wggsYX8HjmEhBO7sJHy4UoEamXLSxcDkwm3GcBW1RS2DJv
E5qGT3AX+Cem8Zyl2BbHlp8MDEXna1lY5gWPscNcQ7ATQYofMj9NNFn59Tb1I2OH
M96by7GKtNjWe8jNQmxvhXkV3LkcRnUAPP7Gfi6K9j61EG+KAGEWsTmTaUmqdkIJ
OZwfbDeY0MMY0ZvBzZmPldSxVjsHzsqm2HLkQZNqi/m5pRiA9i9rWlSrTtGFA8jZ
YTrjhk+rqJfC6MGl3gb2H0WftBhduDP9xB8ghrbAnzyGzjkJwuOQu73qKJkftclO
WRuqD/A7E86ZDfYVERf7l85A0Dmdj+YOU6hJHvY7N6B4LStosjIWAGUrSZkA6vrj
Nq1XVmHY37fZNflAe2+f1nkOr1+rSNVsGaQ5ee7Z9ICxY+NmJiuYqNJ1Dabld+vv
m1SrreIm/d3oEkirKMXZxxH3Ot8TXGFId3ZZ3s/hNRQ3myjzs1tSaWZxNcpUIKua
cFb744393B1r73/LAscUKLPSAlzb/wFUH31agELhlvqhTEEjiEitbL2MRcXEm6Rj
xAMCQz5ceWHN4Xi2WFs714aHvUBNS897yOTgJ5nvuZYLtIG92YLpwMU9erE362cp
8J0WfX4ksE/IDP3PEIMS5UmVRMhrxIE5NdL9jVFihAz1TQu0D39P3aDBkCmt9hEK
ssVjQYxcqvVdfLFMx6V29X86T1Ghzp+S5fSk8/jL/KMtQBLwVdcAEwmNUHT1Txor
Mz837a3fUPLGvcIzbOBUhTxkbq002kDGxD9aH4SRPuBKIrBKHIo1X7+ATzVPMq/R
uExoWJU7oRtAoNZlzgQF1WY7qfwizc/w7LncXeRzc5zRaNCaZZb+vtfN4fsCCKZJ
bGw6J0kowCYGrSuVWsASli3BOlvdSA67bCS9h23RvoS2zTCJGYA5i1qN9V/U3XnF
Mhmu1r4+vLysl4JxnVzsldHZUVlaXLPaIBQCS0prUDtFfd/kqtC5I8GOji8Tu57h
24x94KMYPyH4Trr9Ez17CKPp38VT1DRuKvs4evDcLcclY28J7xB+QJUGCeXQduvO
i8b/OhUQjwoPYdj/zxfF67SmUX2ufCNVoxjnRNePlf/YIXfYtwest17mlh/z0LiD
81KqvijKy02jolGZSzRK6DMxyGXGPpdTV+Lq8icT8M6KZJT4K8Ev/2N31iMYIlHZ
FuLjhxAJwr3vrIW5umLEjXCK/+O69fyaSFmu1E46QWe/i/2tVbqqW3j21BUWLHx3
7P6Kma/8KbDMUliv8zo1+coy32Z/5Y/wKvTJYlU0RfPpa1aGrwI1CajbieZBDObY
PHt1/TcUzpTCTcJKNZ/yXmq9wEqoElZ3WwCq5OQcKJFCaCGtESFqcb5b9GZgROdQ
GhenyJDQJ7sgzmXZTv/GaSkhX/XJxCYeH7aPlNjb4PGKNWUE5iy3ndWVhppSzgaE
xEH5jIVFoyO+lJ3Ae3Ebcfj0tl+tEvKDcMBKMnlwdsu5jCCyc+Mt979eBXwR3HXu
0HCXFOOTwCP/arheyLrLs0dWzCuj+IvFqPx+AkBEbaZDULvCCNj+mdJUlNtcl/9R
zsXUGM6dhygQHCk6mJB8QxdofcbvtPjGAKLkXdtOMPhFoIh/kyVUUXl0ZUqeLg1A
mMplmAEK/Zlvl22aMXSFvnQEKOFVgu3Are9Cm/snAkgZFtA+snHQnVH/c3WfGH1R
nV/G1JX7iUMdd75ql0Vx7Ws3xKxJUobdR6SHCUiPuGFhcN22FpqJkSxLfBJ3jsNg
/9hGOLSGypI30Ap23Ip9/Y7ODZmMPR/1uFJBEFqgITiz9gfqHDTAw9I3vcMz8ePB
b4b5GHd5ShNqiueoFQoT/MarqqmAfKogvo/+wfHRGnNRBdE61U5zqFgLAfA9VBcn
PP6xyGwe79l6ECR0XOKP04iGkjT2nStjAgqb7Oyj0g5G7TY2jZlMa+T4V0sbbOes
g2PoUbIu46a3diVjawf2W1zSwwxtvhHszCJ+HVWIp5tya1JaErAaRF5ME0alm53d
tW1jLgYI1lc3n63UbdaPjflXqvGVWD4NG77iTANbCCQpE7zB+QM549bip4FgrWR+
FMF2ut73uMWx9K2+6ALGMA59Zta4/5UVN9X5w8i546xz30NdUCk6keYAofPHH8ey
RtXleffah3yAMK7EiC1cdxQ0bTPJgx87n1wVkbxqJS+4nOl367XlBPd5HxdhGuxA
z6GKTex6PIWHp0SvShK/VPfCIJDLisB5C/4fjFXNAg0QJoBgchSbLMr6BWG/BuzK
kz2X53cQW2VXhN0JiDuEOLSofkUWL6R7cZlb1KF/IPOuyR2AP2RVBR9nS8n91oJe
X0+dWu77AVrU3uko7DoNerSSHyI6lq7C3jrmXbmCpODPTaxBnhb14xqjiSMm81oe
X5Z01n8Mch93EpgFIKzeuUYa1sSem8XXRLjwacl8YnBQqFHTV646AT7F244Pm44l
clm74fhaa+xvAvIREP9bskXPclQpiBDfWLQmkRbJ7W83TfLkeSbRI3v2n5xw5SuV
9BzMquRkchMqgk376jahy8p+uwQ+7Td+ERn4fkN0Zpg3HG0Orcii/MHF/o/QEj2m
5szUAigOOGOmaUOKSAZtgeDVkZAeyrGwdGiAdMNYIKE+63/hmv8MkGqgv+50a4tY
kr0tF/hH8JR1xErU5fRcszIQYm+6j1YDJcoO/RVAEclyqT3VewoC2J9tjLlalag7
3wPwn6PcosKelLD/x4KzEi8dOXMBOhIssdsCLuBmBdHxxxef/H/OYrVTJ9RG+Nav
nfnEuxE6JsEj1DXntoYOuYPTDNdwaHk7Ieg1VrvfrFEpTefcnDj4NnO6dosemuJD
s9kCepOjOqpEbV4X2DgrUzdtHv/CwS8kB9FOg7+s29eb/erehay/Yd+As3DbLH7m
Ny09p8o9lYXGFgDPO/j1DsO6ly/h++Eoa00Jf1kpQQQl2yy4Aq53B0/lu0JupkW6
2s6RlTK67rx/wfdrKWQ/8XHd9Jbn8HzRJqkwxTnKQWfZxMdUlmERpG1jkKm/h//o
YgSgjf7fUQmCWii2fZgpsZsPEXz40S9cryAFmJciBmlz9BGs9oCQUSjrgc6fMPw6
5jxZLJO9lKL6Q3r1j8fzBquJBdfXWW2ODNTh/vD5LKfd0Aq85+FuiCUcR/3GAywl
bbdMZ0kru5M1wfixIjbJmSkEFxfQcumHMMPz+NQt9XzrlG/oXrfwCkvOpXTRMT61
mrZJ9SrgyAxxTDt9tH+VDMLppXTf7mWi1O06GgF0m1Rp9LB09+GAHcCDRp5VDQLc
bDnwyr21jcTF3neCUhu7yofzxH0xKdPGkXWUwHOsAszYSRs4oB3LbpcO4Tg167le
WKcsk74UBiz3QKLIyCH5fm/Yh97ecKGIaCpfn/5wDIG3N3zHaot1G+1zJH9fmAkh
Qq8bjtNAksKleEJkp6ph3cPF8lut2k6FhjaTNJQJ9NEwv2PZUp/l8z/DKd03of+/
SUcTsMaxdgkTjy6iEvBxZbHJA3Q1k4wW/UH+00Ft9SOG5yd1539AV0MZtBWtJk+Q
LjMfGhjnhupLf+i+qMHg/wTQtRWptxWaHkSyUW8K8cnr9lfK2XJGi7AQMlUvQwJU
4BCj6Rie+NpEJo1OF5FGnpv6hGBdjItMIsFIhg6meC706yNkweJvneWnuE7/djQr
zte4zNB1dF+XDFV/9WCiEXVP7zZzhBvDRqrBnk7/krcR7Lf++QfB4mvuuyH4R2jO
1e5bhw/CP16xtMfB916S5n19PMuNPv28E451esHNo5Cuh1OahqgIIQ/6PG+0tF6D
xkbHVVtVIJJIJjp2IQJ+QG481lV5CRD7JHK4MFcMhdxF9pensYXa11lyiTnv6MYP
xLX2eM6UyzteOtfYuFw8yOIdmC9rvPlI7eAKTcvH0028cnZuz7KmNpLvZpzyO3u9
4NVfBz3d1fI7VsTh5XOTNiX9qqj1ubmK74DH6igiwtt80to3+nXQv1xl+pG2kMw/
b6GuymUjdXuDErk4N/paU+0VonFKpOmF6aWauHdlh2DlgGVfZxLHONi/6+0vTTCQ
nRlWBI7grNb5ibHM4V+VTrOHNAXYwDI4rwpj6ZowM7OixFLKEODr+nRYGan/y+MX
Dyfmz0dQ9YTZw6FgWetVcy3nId4KdQrkuJydASCMwLqrmWNcLi1/KAAEpOsSmgyn
2b0BcUbTBGLkaA+6LMBMU0BA9N8LE5pEVsxgPPrzaa4dg36eHZ4b3HC7XH2qG1o0
R1dzGfsvEzJw5GWynzR/v6WcnMroDpyVZeQqXPYGicIqTGMPQcTLYop4X2AtplES
GE+BfPJQ/CHe5KwwKLd6LkMYfs2DyR0BfCaIEcan08E7+XlGAODdwXc4Fbbt+y2x
gqE5pp7Goy1qQRqdJn7rUHh24RyLXPtQZJpXsW6m8N1wW4/xU9XaSx4o6QeQq2TB
R/PYkrMLdf1kcjIYEAJXTR7IJi84/FpaMnu/NbNy4k350nHaFjl64P3w6NO6aace
uAJrwtDfS/m7jFxr2qq8dCpGFDBTlTjVUl1wFjhIJPnz33OOFtgXQdz4kn/k2eHY
FXHDhIsKgApIWNzoKfhHasiqLIxZGF4Ay5woKs9q/jDi8QcfR0PwEtf/Kj7poiqH
fcAg1fbhzVVshqiz9XhnrvKAfjVQCFXu2oBKAuq/dcF97ZHP1U/wPJ9sTyJ+nxh/
nhW4bwr5rfSjCJCBAzQrl9UMHMVxI8Bk1h2m3O+j1Sg2TelxuD+sb0Us9q/ka/b1
419ZIrnLxQX+oyAt2C7pVxcNL+jed6EHiEE+LSmxfMItUI1Cxxae6by/dU06FqRH
xW2079adsIEKobbzYJR0j5eqFtA0ekQCmNu9Um6dQIOT7QMkjmM6IJ9YFZN3qyRO
m4V+BKUrJdreAyaKzEmXJ1/oUjlDxIsbfjEoUDCf0J4QycNSYhqTMIOjAOdsjnuW
UL13zzVQicd1l+iCFb2sfn4o7h0vxUoTvxMuz/3rUpIyDJxyYfBgK0pEjrvKIDZW
5FuZhCWPegELsDGS3EpGvO+n+K0tjsgQwQdTJEsU1qTSUlVvpVZ6RDFsYHBUJqdS
OjDFf01sitr58w1jaOkNflQDexTJ+M5veho6YevhdSir5dGQuArf1C7iIAq7BQk8
FLBZJ4bUV5CvVlHfzYTb9grYr/kfxQv89Z9f18p2O3BJeJYxOa/Tr/2M8IWF7WUd
73fh2GmRqRuYHB7CX6fNCi/qRDsLSAnJzIFMTQJ1APjl+R+KNJAXj/gtp5WMhBJm
Q7dl2HTxzP0ziTodfZYn/VqFbzS1TuA6x/Cyy2ay2V+zBgZYzDvriVjHgvdoidX7
Cqw0R56pLFKeJb0PaNmOvYM9atoA7SERdNXBAlaXxCLx+MvetTKpm/O+IErkUlE3
SkG8mKYDd0pbEdzamP1/Bs2xzWTHbCZMB5+F0rJiGYf8kpO9iUH18UXXjonQ/Gyv
dP6LH9onRTCIi0NOdnNGBmmOKa5IPm4SVDsdI/HFCNQGQoxND45uPeXNkKMptZip
ICPXft0OrbPiNZe3+hDzIL/w9NPPdALGOTcgv+E/32TwMBo7847J+ohFeXIWpd/M
cU9XSowDmY5os2JSTfryYP22geUGHSg/sJKhqjXLj9LsywqbnG0dcgTGj9oODsE6
NugPf6ZaoYOOnGomZHIzwvzBGkZb2G/qSW1a7z8+KoGvlIX3POUgK1TfvKIb2Poy
kgIbxfItV9B1f9BMZEDJkgo6yNyQJJ7kLelPOTtJy76x7fo3KyHHiaWXiUVZ7/GS
/4oat4xcYJiPWtkaGFDx01boPwv7uunn3EM3Iwz39+H+k7jqk6Yn5kFam4TpqA6c
S+oE5+xsh/hO5kOV0WqUBzkAVurFeSC1KaXgqcmGxcj8AZloCJfvDnla7HK+wQGK
kZMSaJK2NF8UuflxmsmlKNlkFdyXEgVzCLzCkRDKdRtK17M7qCOaqlhPFos1wRwV
6xQqj0pvashJcX0K8DmfcA02i6QC1Dz+eNY+XqzdEuWD+7mEegpvgEVK7GQAiIM8
OSyI4ugmoM0+d054dX1DWn1vhs7HYxJhaiDryVEG1q5Iq0wTsvYM2zWZTeWtgKJd
cKpKxdjhAHkIkq8mxhrzZHWvMv4kmgUovzybpwPXeiY9bQRZQ1D7iMFbdu/X4fLe
BieDjZx3CRBc/OCIQXQyFhtrM+BXCG1PCXwO8gqbvkUTVkN/fVseT8tsHpqke55N
0/AZtWTyRcc7f028k9LG/QYfGwvRKslAGCEFa1I2yYJKEtlzYPTywoNbKUVzMq5R
wn6bSF4vVRC6wcmq7zKtOLnAwh/sEhZMCcUwu3IMBcpr6nYbTMFB4EUQXw7TtnBr
sFJ5tNTir/5iIVJg/JnHXngEg/XX/pDJUSb1ZaKNRbFVrtet1Co/RkesF46L/11F
WxMWqUj5KidENSkn2cDd34JTwK1kB4KmGrixs+Kge9x2AlxP/vkDd6U0R0IypNbr
RAOPXubk7ZRAFblZlyyO4/nsR8WylVyUQLTcPwn4vPHNMVI7Pe+Q7jWKSgYE609G
ZcQ7gdYaWZwk+nFDnt7njgGMsES1IRlrMZO9G25No6us/v8tihQ7o4o8ur16WcJK
iWWRKESuin9D+XV2YywlZPT+CaQJlfrFujla6B781c9mayhF4ISMBX/jSB9Fjq6B

--pragma protect end_data_block
--pragma protect digest_block
M0u2YBemBaU5HXS9rk+x05gpJyw=
--pragma protect end_digest_block
--pragma protect end_protected
