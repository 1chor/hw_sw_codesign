-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YXf5x7Kqw2xsNIvzpKiWlQv6CMclBqvInYfWweEWn2euGbEuTMymaZLBAt4wrr5OsnaSlAVUFFSH
M/JyZaoaDN3hGXluSwnI7sX1R3N/rJChJYk6GKj8WcEHe3wIGZCmlATPbFR46nhRF83/Z8HjWURe
SaGldOCmtS/cqExBGHrqcbpfqoeslmwU4G9caBNcNR+IN6cEu7NAH3RZyt2wZEFTPaBCHAtHZ+ee
X4svEBW49seey9M1VxWUYOTdKFMRYX5gureNSm5JCeM6N3VxJMIJBy7lgyo7rA2MTY7Erd/WMKI/
1lPDBv+5X2n0WAdao9gwbquwwEmCosctb22hpw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3584)
`protect data_block
Qag4QV2ql/hbrEWvZ/drTlD6nDVub6G/qkE/cAWWuyyr/afRzX45+N3kLRh+HWQCTUoQ1swTbXTY
fbkBZ7NGCw0Gyey99d7TMacdLbSRoyH3vZINfLppvKjkqarMAav6g2sNMPtm5nhOP2VZsCuejgRr
rps2S0hOpX+9CdWlgQkqeDPFmEZtqQYbI3P8kOnvwt9PjsHk28iCY/jHy7f3On1ripVIYqOJ8ea/
7lTiRYXhn8R+FB/hJcgrAgmXVWNVTYX0qB+M6/U62k/aSxl1RrIrGLcATpAeih6j9iHZESS9eLiV
CjmWBL+HFJFp5v+HyJBIMZGeEkQRGL7LyzZSIR/dFxl4wOI0UZuZijhBaEbD2wCjYTXBO6AzNQXs
VNIq2vCpe89/uLydIT0o3SYTaimk3+vSh9v6UyncvF4vBwpxxzGw7vwUHVoKIgvNyh3VmVvpALmq
5ugzMYHcwqzW5JqdtV5zRqjRcBlaLlcqHIpQp9XgNrXW5UZcR9fJAqhljC+9Tal2wOc1AipOBDC3
SoLVoVLJ/0A3hJEY/zY0+1KnWj7AApBPL5e9RQk4pZQmdUKD8PgOoWGKj5uqpBzOE962/NQHspkI
JqxDY2TOTax7TcFuJlkkOc08CyFiKPN5X3BWnFb+l7R+/5OZ/00R0Z6rtMNfySUERe0/GXNFaLCK
TwFlxk6k7fBVs75sKaw9qn8uVSeZUpsUbCyKeQ+nXcTGtaWCe7ujTrZrDvyyq0gFKoNciFYxtWwU
y1UYJ/SKXi2ahM9d6fM+pFVT3Ke/5siJb97jXCeAElRptu15Vy77Mfu2ql4p61Xh8i9yWimtWWYz
+VdOW//rOs2RdATr16moKdlXxanhwrjtVlJlKQABPFvKLPCLYL6WFRVuySko1ASfHXcQNBxwnqZw
/V2koj1wSoqPycYh+mSQEab7c03xvw51lyqQzEUGPr0NqKyqv+2RCGTMLpKj2azcqrUKUSNG8KEE
6BYSCIfoDCYDYSmPbzUj3k+6PnBFLKCJaxiMwi+CPhLiLztolPXgkRAHqxTRLA0w+0nr8muB9qGb
NM2z5DLvE+c78U2hDu2Yxt9U0xbdEPT1E+3/j+Z/ILS4JxyDAYrxKp+TwbN3xjNsLPD7r0ewD55l
5oNo9AU3wW4R+yPOO8CXzkyGUELd+EvZ/ZPAvGCdJg71cgrub72p4kVSuzBh5pjVxlLuVzFrGuRF
h6k5HcZ5e1Lv+evfuI8NvwPvZsQ+Bl65IDDlZMErwHf+yRBxyxp0FZ1BM7kEEIzjlLYkCzqymxAX
fS9LwWb0NbfYDA9paiscO3INIT54e02PkbwUvDIPpELOi/a1maTvABbxRqQp/vaOw0h65NGFY/4F
Shy0t1DDVQ+RhSOuTzkXtdwjCCGuSQApayehMlm75Xnqsqwfr3b+FxOq2pHVu/7IDExrV4sqFnq0
doR5/JG58M+Pyg+K72m0cVIUNfsXR+HaLpL+4Eb8szSgkKgemZuDHYIc+vfpIf/YslFtBq25YZFR
Ho2rnNzZRW+51MdP3bL8ExAPJXcnuqLKmhh2Vma+YSYzWkfXesGay4CuZxu9yfT7NUwK54C085qu
phpUVFfKgsWKmx/KE3S9eb5n79lrSjRGdXi3y7kNiHm0yHR4VknqCKiWP5O2evEjBg9M7NM/juJK
YWrZi3rz6JlF3Vmo86mjX8QJ86L3LmE0hj8TAdulxuMKayECHMEF4hj9P+HEBZ63HReR1asOWhpg
bivnY1qj01S+jTSA8bQIsyxIk1aJsTO6d96peJJy8cDt6ARYnBvFIDZzMm4e709kbKs0/xP2Tah2
ub2n8xbDK40IHFsPKX7vkry9qOqxyj9B6P/Wlu2KmPplGifROW4BiJt2yYmnuruz+guPtOkDQ3o9
fUJUc8IfVZGXeZ3KCyjjSWbovhjhDkTTZPuA4rgfCxzfiTnmrGEgkwlc4+4rlcgMZTzeBkdXrffo
h4suPF5HGNz52nOjGQmL7M3qmSFVucMyu2ayBws6HhhiWu30Wo9FCKonEy8zOnAH76z0LYeHaHHN
dq1BpdFZIp+ufu1X5scbgwHcPYp77XZxlW+xv6I3VGKcLsHrzsNcue4v7n2dWbRO9GpftBfZSLeK
1rViYO1PtDGoxDvB426ALig60QUPOC4TqInWcP+xUqr4aLX6GSXjJWQNQplvmAMTzi28AGbMi0Hi
a0mWZUP33A8IVCi5xKuEcfVFIpfzTY6yGvcT1eURfwJ8K5tI3xjdPmsbAKgbBntju5AFlGvLU6tQ
cSG4Mpn7/+cr+n69puvn5pt2TBdkDqLG6xQfZ3zOmJPm5ak7DJs24zkGIVki60FKtcZ38P074pjT
l+6fnN4N+yY0o+ajfopll0yT4pZCSYW0NH0hgcwVyyMBfaE7WV/i9WjC5LUqymcBqscPjtT8GoiZ
be4xw/iB1vMLvjjmL8h71v3huonMLLbDwmhqUDLbqEs9ktwBr4v6BYZ8I95/ZihcCCQGLlrs+xUe
nRgl2nM6FJC418+r69tGa8vThol0WhTjboL8NM78QRmccieC3sn8qGlt2AQwWygumRY9eyWwBKoM
Eg8a/Ll+wgGsvDDSpkrbBfY6lDfc0Y+VLOG3o1VDqp8mPdj/7UWmS++V7ZXdLehzdaHoPpD38DMF
jcft3YlU4pDI8tss0V0RYzDM5jMKe3a2JbgteDqcxa0L6O2aTRD2XJnunIdIphepr3htmbUbLJOB
9bnS17UHiUTlizrE3bcT0i3zZxz00QeycNF+WNWqKrE+jfd1rdZwK4wfNkUngWku58WpeLDSaVTh
ICCuPfpHrlxbXyXQQKcp8QJynEhmLRaaM7BrBF5QvN/6IlPTn3krMDY8Y6g4zvrvcoB+jS9vWvwi
m9dpy8rsNppC3D1kM+N9BFKwC7+D8DI0HZr/GL1b3NeK+T/BBHn1ayagc0nUhA/icfPZKi1q3Mxd
SN1NMCyE3M7yKCAn/CYQOUfhSf9B2Q+t7OrdFwZPnmdAry+ESDOxMMmGqzV4ajd+RB0SCU0DOdAL
dbfp1O4TZOs4YbbmMm4sEPbZzCWprFUIDRAFN4fYjR40KZHrx5EvNiVTT8626NkgpN0f40Xcmlr2
Pi+pSkq5Z3XYhDYiz9ULtne0B7q9atP/0Ui67lKITJX1bwIZiRQ0Hfyqab9mdtmuJZDO9cgU6WGn
hNVKp609ok5B4XW8nh/7NkXfod4/3E5C6+9eOMF387Degn7ATg5n9pWQEUSXoKWStcNIT0Zm21Qc
D9W0eQ7NXzb3YnlQg73GQA2r4ZR2jY6+I7cYvNB99S4Ke/jvCqeTWySAV4Hru8xx6C6A17Ic2M4f
hYY3aztujm5jYOvjYjir90xf5priTC3ikTqpq3vGU4ZJ+0WcAur25L7aymy+VrfQ3S93Vb27KegP
uM+F+x/hRuiLqm316BaQltjdJ7yTzPf00f8t4fGFiFcsMQx6YaOF57jpFPaWcuF69/KiYI+PvN7t
czRRO6ps/f5R6Xo+KnMRiMugnJbIHpU70oKYPrVuD45pS6Bj/n24f/0ltOi2CQKAPNH1IOdD/NYT
hl28coYJBRY0F+ljHhq9NeH3YMykFSNH6eoC0v+sT4AtUmWGyrTQnFSaUnDLC3fuwofU+oL3PjKX
XIRMQnzlJZ7P0tyVBCtWNsLLLCdRUZZ1Ydus9/8vKaIf4A4/2dv87PhVr2K30meBbMnSub7i8wmc
ayoM8rZWxwtyOhPrz9rWwXqGVoqnrnvDZWLYc4tMoKuRUtx3pgn1F3dJZPX57zkomeXynaYdq/0b
3x+a0xVtrxLVfzfuAvmOaK2B/OnZ3+RwUJDvubgwD0E3uB37esuOMR50TbeCk15YpXEpfaxatKPJ
/akiyI87mqjjKpukUKBhxpMefvIx1Rt8VtBYC0UB9QVKax9Tx3lb68xQSRrLy1/PGi3ZJ1bPE5t+
6fNf9sg0OUmSLuFz6DBmznPwpi+THb2XJzVSPB+aJIKTz8O7jkyFdzgWyCw67StjM30VkKtU6DDS
66GEy4SKebOjDzyphdqKsiThNiCyWaAakxkbyOjCrs7DOuDBtyGee43na+B32qtAXL0zPCeB3YLa
ghqyceeQY2K9wp3f+UI6JTxQm4aRiWY/uWEcmakcHk6iT7P97ofW3z+PCmvVBaWd9Sy80Vmhu4IE
V5OyE6NIQVJZT4rlCcyxWGcq866r/1Jse9PGIX0lMRSQGKqo0Vl7cE/SMSZtFMQiL8QG/1njeHsu
nLL6I+MbNRPxICB9aEVthh/se56ujs831OTcC0QDPvElYXt4464AGBeB/yYam7/v4vWgSEtQX5eD
sy/FihMaN/YUVNG2sGD/fruf539XoLDOEYcErsO2YDCH87wxRP3pJBi9vdTdyX5rQfSuJN+BKLIW
q3mSFQLZyDtxb6qTwc5yA7jorNSYFX7UmQ7QYajK/VUdv6JhtiFH50D9JNRzcpLCIPr8bvJXI3Ti
kcE1xxZk0vDBajtIiHN19o8Pl8YRFxJjqf3sHdyNcqJPcQC4UhAXEYo2LYTRD4vfdRTNZiMPiQDv
MGtuWL1TW2wxnRKx/fJwJhSGxKMzUWG08p3hZiDveE96F7ssXBc99TqaI7/gSC6WrkzTp9LvHKV/
79iu3ox31d5dRUW6ZmGtYUFgX4Xn4Yv89h7NFARcY7suQxB6nAsRFfqmSxFoT4qlxyZ8xpPIGhLR
0WzuA2t9fBspMByVFz/YYXP1Mg7sKyRJp3XCW6FUjCZoCep83zOmVM+RMdWYCDVBdoQ=
`protect end_protected
