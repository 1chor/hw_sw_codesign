-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
do9ics6FvsZi5wo0ydykHT2br1Fsh9gfzZ9m/PZTO4E43If/VzHVPy/YNVqZgrRW5w4eazQ9imm9
Oq6gwTNeEp9jEg93zxFML3CWDJ8TyflcbijFyGQQVzbi2FmAA/J9HqK8Sp+PMHne0iV+ZAeigG6X
k5JR0xomlMD5AVVa4fjZM/WJP6KSQXMmLfHmxiXvVX1pK6rgYpDdDh5739N1Xs3BSjBf70Q3x8/l
53gOi7bQe68Z81p1dvDjqavkOFDdcRhWLDTEww3IG1wSi/S/aqWEYMsl47EiFQuZM8+Gw69XSk60
tKHPJgZ+rQUdUTKkEhrf0jtSzgioiJnd65MnUw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9200)
`protect data_block
RxuVmNpfQ8qNU97yEo1E2qZAl6e0n5bSrZYdiOHXYMElfIoWYojCyPyyGbmVPzHNo+PLPftzGcfy
Y6Yl9ixnAQcIfj5a31zRkgQIdQA2sDuok58CpINBOCfSnuuBXO26b5jawNSdU+5Ax2hf2ztRJyiG
7vn2ShUMeeHB0V0OF+XR3h+DCEPjAjJSRqPRPk7warJhPqZwGn4+dggSg0XcP00SYBbKId8PgKvA
ia/aqNCweLGlUJb6gR44oyOKWj42QCLuVFNoTuEMJhlBBcye4yCCEmTOFujWDlfKSN01ynUzVgVj
fy8yLdFFpxHV3zc1B/YNdqqJnc3bZc6YLeERczWpL2uYy2lX+V73WmzDYyo4j8mzovgC+x2PXbLp
EERoKY7vOqmKN9xdDObS5HGklZZzNd6WkIyhtQpZoxWVLEd0W3uyO0O0KqZgFQX98o+3Ro0I6xcV
vMfgucwrK7KHLxhG/n2UQL8ICL6rqnlEslss53UTn5r/YOL1/VCSFmEoVLDT5qv3QTUAwkiJcd1V
qJ6n/XqUHyyghOZ6FH1rS2nq6QmYtl9assUlxylYOFPMIwtss18T3/ADdC4+Ur9Cet+ddxGdTQ8y
KGl3ANXmgmpQQykb9Hdr4WKTQ/UgkzxwWqUc0B6IvR+dJ7be0tmN0yByquUJ2t46wlpuouRvqBX+
3oZr7HVlkSx2WluGEH4YnvG+0io+K2kVQ1C+SIuM/6198Qqz4HZASMC0f9b2Y/GUg2mhVvVoCftT
7b6OnAfvKWxEdst8Uuj/y90v9rVwQ4KD+V4F68rfm18feYhjCgh+bG7N5d3sBjJxc5SEp0s4AZAJ
Ye+YOhvFH4V8Acebi+AqOLKlF1fiQgUlw1ENFWl+u4CPuBfn18D33NH/YmZ4VumeExloibfhcaC7
LIfbnOQdaJgwn03fB/tfgMvsngrIyRl+rmAvAE3FG5SJlKFuji3x8DOcNgkEkN9Vct7hL0XFNJPm
P2AXKtBkRQyfiBBZLBzWVEzkG3bZ/BDT0FlDUhlVPdKZG8AQ1dYhwMKK5GfvnWJ8aisCsEcX8PF6
KuhkUeQnkB76wohKcBnWMz2ayPIR76gWQguqRZ7ATSvMePLsV/xGplfPcWVYofwyOgDgRKTylsPC
pJK+l2zZNLSTOVm9e/dL+2zd5APKyPHBAMxjfX0PgYXKQBEulMaS0n/gNN0ZphigcBEtssLKLNjd
R2d0ZljO3ygyjDDIInzG/9iPibs9yendXQBhDu4O7e6fdzL51wxNfYxmNS37QN7L8ZW+WL4jlthZ
0/Un3X+WGxVerLBSLUKEJ+L0gmmeTWnu7CZzahbA/LRSinAp5bS0yg9quayYPXGmwp9u12ogLLw+
++m467g9YwiA6TWDIeVxfzJxGGE0aPXr94cfFf8bzwUkTfZ8xjR/gIgAX5paXAn30WDOBgCX2kbL
ZIe6MWsd0Jd9qXAVlZ0ZTcz1z/TbQptaX8mrnAY+hwNvwggeqKPma14La54tkfIOKvyOxaLQHeUL
pv7+dZodszTwUEKj9dYliouMRRlRBWrWsXYauifv4hYRbVUCRDj0fo7+J9lBZfkjI3a210RINCHt
0FUKWRjm4/4pGPoJ7upOodAG//naHD+azUEYyAP/A/gfBRdDQZUY+/NAwj+6FbeAW60aXAFU+FL7
ATQwBDgiB9aAYl2IEuvWUNj5noHDp69P3U1CvIviJa+EpVD2pv/tBES6OIlhe2mqkqB7Paul8MpF
CnoGA2mTOFxZ5qvhAVWdgjFrYpmBF35wl9hzD/jsyzbn0kNaAZePB4Sqn5y7123SS++lNySWmXCK
0DkXIAOcbAx0Izo8xxpc7kEWDG2v+fxoSMarjBvyjBJ7pZJtY9AbC8L/KIGtx/Oz4Gm0fLKlUfhS
srmM6GDFBq0a75GkM4Obkj5x8nmbaF4NZYyCMPiXIOL6waMrBbWNSa+KbNK5OByxDVIZw82rY0N2
6vghNyGXxHA00eDehX7+iasMCp4aIvkuMhPpIckiYMO3oi2F4L738+dX3a/CcCHxwibgUx/D23Du
K9FaavA/s37t5/qwJ0RjTfYKKDH4Q7MxydBIAIRzFk/mxZBSJCoeNhCDegNQ6ZrrfNGojiCXh5kx
iy6OMhd7xxs/rL1QuxQUXxr9845J9K+2un071xGo0h7V5Nnyplis+ms7TuBIwVxXSE1bdOH8HvWN
A/s+VFrAkaWGPH/eRUe68nmAcxMQjTkM4mGmSVOYGRc8Y9vz4aySA6jSCceGhwdvMqxlVh167F0i
IYfQbdO890gFMXw7nRN7r1DEWf8mHnZboiE9x6tj+coxoheGpF/pCtP51ns7EtpH8X5vPOfwrj9m
qQix9DUnMYtp2DiMpKf2SR3IAd48Cw0K5SFcL3IqeQftgU7g663WdtVDQXTQQPMyYt0FScq5Q47D
ICguX0YFCUiyLkC2SnSrt0IPDFrtKZDZ28OYDVsx0MNNmk+8dBbo9wsE+mMYzTvz/XP0od6LDJEf
XHt5UvQs03pGS8hr2KFH2UKXc1Q+tHGgWoHY27WhzKNnzingO3ApTb/G9Jwv53N74WoCYaSOIC14
STmDOMaRWDSuExewYg2YszB3TKxbkdfCw/e3TXTA3TUWOdEY8tyE3ZOxDvlUqAP351O4tXbXXcOV
DOj9oCunjL9OOJjeGwCDUtM7HNp09cYYh/ZxoVC2pbHgS7lNAFZqcGXXMP7sC12wC2LvSDfWseWo
6c29NL/P/++bqFF1O3c+hdEvjz62prldlqrPYMygIGUYo7woCGmLCzEJbR7DJFJ6efJx/kzcPvS7
t5cwXop5Tv7XDw274yRmw4zqR7512lYDq3wnDPaoRcVmVTJ1ZFGTBcMR7Wo92V6jPicfDxoim+vx
r3aTdoVHeq9WR8bffgAqoFEqYSA/6VZQ0cGrA0lisAJcnFOLO9LXdQKslxWsjb09B/kDBFwOZUMu
ZSFJTLGz03Ge+FhVWhJlqk46Kr1KR3h6vGFUruMx0TjHk3cQsAhJtIgFnsHn4yPBWOCqMLyTmcBo
fpehzEmJANRLPTOpGBmP9yZCth5RfrOdizIx10CDxJ7GUYa0JK15eyCFB2QiAK3QbBJcieMnq1n4
rKzYx5HWTD+WMhby7JL9x+fueO0Bdy9s0jlDQMRApu/Cm2a5yuSOMiOPLuJmSLm/dy1DC93lJ0db
sHehd4TpG2HDx6Sw1yUxSfJPw/2aATvuC4xJO4UfjZZewA9/Zruonc9gSwoL7N3hiQR4FFwKhXJq
3UXQidInBjnmPlOX1riu04UDR5pE/CiPXH3rmZ39prEFPaxBscvHZ51lFWK72Xc0ezJ3JirbDeG1
r6VduVmdJCMM80U5MZ+y1g0snfbPoUf8YPIpLm6yY1m6vTpOkuNY8BBeXcKZGMwGNoEOWsz9Za3k
TYG+2ut/b0cZ3DWYC7YWjssqMabEkZ5FSjKt52eRaPo/3wgY4aie3/TqL5R25MtlXQ4p+g+nEvzv
iUnrMoxgOqg0oENLDgolvhXpOwvVxVgyXCO4e7n06v/5sX8x2MfPKAmpPGeXmoNp/IF6Y1fsn78+
/LN2aKQiUINC8BEtwk0CMs8lhUmJVETNtN9d8fb8rWAZ4U51bcG8YWOfMXjWMwsB46lZHZbY3zBy
2U+TPj/abZhoWge3RN7S5QR9UgAEEcM56VfEXA3n+KpIjmSTdvb4FRBMY3Yv+lagmeiCQJ9RqV/6
oPLRyz1YQEfc53GwhjOxiojYlJItRDPRvJfG7SxyKPy2szCLc7y6toIrCAFKHfy9StIiYDMfGLo6
1S84B/EQTFS5GirxI0jnD8HFvcPMWAcLpcTYM0+Vj/Hc9YtX9K/YMzBFZrfcE5n1h0pFNAfYQBsd
0GprB8N0Dk81SAuvoZwhLwVcbqzkdiAgwa8Hr4vIkGGv1DESYTSk7XCxhvfkDu7qHvQ9VNrVquJ6
Efuy8/ETEN/hDuXohVkRFk6Fh4U4QXt/zcNukaZ5U4q3lUVrWZ9IDfOG7EQ0NC4nofJccVpCj/Yf
23WajIMofppRqtdK8u0xNdfc4TrDI6a6kE/1oSTiY4MBLU24h96jQy95gqVtLu9J0siw2QvcNu4C
LFfRoyViDoIyAbiqXVY7D75eI+VxxdS+ifCX/LnZYkD2R4ysFWh9vPQE1n7baU0YLtHqMTKmutI0
mhSVWFFI+Qif4bbA1Lp5nCemW4PHB5Z3d982Me5FRv5xVkwRqdlmW44l4PCY3A2Ga0STR3IB2SIL
R/3RZeJdLRke5DEaMftvcBgGm37EW2801KHvyh8QjbWB3XJb38KB/m3ea2sgVUYUlB0Vu/aOcq3m
AoXrrN3oSWTQ095ey14I5Wwl0Jjp+GP2iGMYsNgpkGYIFaWeojmUNiA4qLu4v3foV4m1tkgWvNeY
TBvA67fh8l9CPfkbzI+W93LLUXKM+WdAtXUC1pPoepav7BIX1ZMrIjiWhOKW3OC+tGMg/xEblvUq
AnBChtYW7OlMVL/DzNTzO9Fjirob2nMmsj9pNiXdmnK7mTwxb+fWnbq4vCcFvH/52sCtchtoYvxt
W1730TayYg5euYcYG7ma8GlLAyHvsqrZwwNewbKdhshGKKMlkRGQE/tr/P3ijY42J1tXY4fygK2i
kEhV8zRMpPwFnpYep//vl/7A2srhBgL/XihNcRw/3/aN5IR0PKk1u9mQX1R8ZufoPqPsiR4h2yuC
lKwxoRSP+DN5yPuAd/i6+M+suLYJGyoKhrtUmnXjniQfg+6reNu7b+6e6JOCuKBCZy14C9kXuG2k
mpLkBh/vu34/rvAsDjbRrzBmulHCALxuavEeaMC0dbWuiwL8cmCPxvMxaVlJPIT54Xd0PzdFEgCT
Ndi5BBuY37pgliEFdsNaYy/aeL660DDJT3XMV36Fg5AcZI34xZo5Bch/OOjy/OEeRWRmk56/on03
ckH4NxHe3GVc9csQfR8z8n7fQ0AUTGSIIMIZ1caAbQpFt5KQxin5gN1Rf4y9LFoF7u5SDXfIcYJh
VjWwWwgkrFJ758/oPKbGiyMOSV2yDPK0Jalw+cV79ywbGnx9jbQOpapiZc66LiXn+JuOvVlfMjr1
TKocOOWyoAcQ/la2gnpUgbs//2A8b/8sKUP0Ss1lY/afviOffCh3GSt6vIfNA9nCZ8jant3uYJD4
uPM6EBfYWAVSf1ZlvyK4c46OWOvcG1tzPzcIYNPwXTWX48PcaD0dqoRUIqFnDwIwILkkaz9DyTmJ
PhrhEURAyrzpicWySgGk81ZKTo1FODHdbgprF4tIwFeYXvw9UrYHskY76gluAPr51GUWoOME5z9P
//J4yYiG4LqJLUfvDULoTjNghkD+ordmrKduk25o5Jd/raHAhaUfnnEiILQKypXT2KcortsEE6k8
RSQrVIaxQeElMMf7XXOCjh0Qm4qo29BA0+ZrIo1Uiksj2xsFrRl1kQx4ba1iICDlLPWXyAlDb57j
oMDgQXKWbSViuyZalK46lyxaBwhBV+PR/xeUHNchGxrBiTJ4F4kb2OKwPHajOuASx0DJmc14n/Df
9C588HvVbk9UbspKU8Ah575XCr7ehpSD6YQZBKt/RW6Q61tpiSjdo5vIuB2z04RtFOazO47bXuuo
naf2Q6kKm7D9J4hSLHAWJg5jmSPDvDhVa17sm3i0Y8SiPP9FAmMbL4iDS9DiIWhR3/FWg4RlkXjy
k6E3wpznqxkxHi0lPjK2OBiNRrez04W/h1+0ZFcvHfdJ/n1OnPpJ2FDFC0oA5BRctlqSVb/VsDPA
qjwPfVfS7qcL+DYGH8bC2vG83ytCGsqk/fAsfYtqVkAsWnAnHXBypPhFkhah4bSqlaONZN7DbqEM
nDhkrLD1eDhUd9r7mQMepAMJy0kZ8mrE0aGz+0xzKFo76nmagIXESZDXhRbw30c89Bz/Cyod98VN
78cl2OlhjwO+RPWZrxI1IwNl2nrZSyJ4nMVVEZaCxSb6ZWdU0pJ8Ngf9ioibeUhNZkO58ms2Os9Z
+GtumPTTSbKIOGulNH/dbjFIQfXsfh4pti8Gp26fyDQR//kJco6jyvMRsHKx/CA8jgJ7umA5eTdv
SdFC9ywYrF1kBia/rysNjfCvT1RxYwZSthACvIEq7rqoFBRymz1Qv+4Dxywvv+0J3tqyrPcNe6ra
L36RZVWDtOfygcAeEF/O1mqdSjaMVoRnTUQMYZN8l5fNylwOpBNLK6aTxHVw8vYcAcOlpuOVF7sp
p8TohjFZoPmv2dtbp/uvO61wKb9iyr45kjtyAjWGlP9/otTzUBmHPMmqlUPGCYJlwDqoEH1Uq8tm
l661KxPoBOb3Sn7dHCqMaj6Y2u7Mv8DbSdndWVeRkD8fvMwlBQslu6Ff8SvX5FnkTKJi41M8Pg5y
1T7Qg0F2tYdAoWrJawBb+sM5mkAeB5uQcQcEYCEi6W7tHM8/WmU07IUAe1mCo99kbk66s/K9TY/U
7R4QLATMGY8gARtUuVEzVxd3pL2pyfB8XmOvHranB9jJYVHjGGAG5lCMex/KOQ3ViLcLX7sfqhi3
kewGtpYfsygwPfcgDZj0UKUaLl/NZgUH7+2G/p2qf0+x1nx+dF5DGUdKYSFNVY6N3WOL5dnXzmlt
N4Jf7I0N+Aw7n1e+0ezoTu5T9zEeK3B9nIq9twDEKmKElYOJdNUUxMHQLXbffwPPGnOKmierh+B4
BDjJPi/dm/m9LDh5KJ1GyHtQNBXgQcAh4tHjL1TeDattF0la+AJJrEPdKPmcTChbZ9WY8tDPVsZQ
gOKiae20eNgUz709i//toUu0eKClkWdPXAFi98XPuKTqgNVxx9nGiR7r6vccrLIQi785vjpgj3UV
OF7X8vAj5WwRx6zVRBCgZYaNp6+CwQ4eNldSbyOvdzwsNQbRNSCbqzg4oplu3sVE1xv5dywRZmi7
iTYMYCuw2aPObIucRjY/O7aUBWD2cli8Mj/J+f0j3IN4L6ZgQHoy7edVhjGY7a8y5tvu8DRJKZDe
SdlhiLbTr9ImIeBBE2b6xTnYmp5YzLZlmAYl8NiGdPY2BvRyeTUnxHyax1r8ivTdNpErGDNtNLhD
dWdUb7HU4u8HBxCPjZw4eqB6edYVZoHXTwqM0dIbxToG966x/pWV/gV3xgbHXMadnGc655O+MiK7
RYqBKXP07kJmHLvNVbvD0DyQRgFCD2uLXyZrSGCFXMv/Bq6FGUVrUYxSYsNKi8KeFXidwdfG+MPt
ERDwQAhhyINb0suncizms+CATuMxw86YlcKYr2df2VLITtlW7izcwlmeV1Qh1TSXsoID5T7CAvlR
6vQfIfmW+6eJKlBN96ElhwgjrLYO7wVu9z3DRyAstBoJZbT2TldBcNLFSvwqaqaVRbFgMc7v2x0E
WoudQXLjPf9Ai+X+XS7bgWB6WDjFdLHJcud7E635JTvvaWwEWFYmxrFAPHeRrX099bse97fPm1M4
B30+bF054cYe0k/kkoC+kBfW0A41JTwgary/99LHQu01Da0js4eDXyLjfnE34vJ335/h1XZFSAz7
ynDOBWgBssAL6juhW2nOOJK/OhfGQp1IrPd+WhABhobuPl3xFCJTBfnKQpDp1k6BdEmpVlrX5Goj
BU9fSPClVmWxj1DSpQizbsYRbjemvevTnHNRgHRaRGB+c+3IN2pduuxGH2rbrZepmIf2Fr2V0ljc
9Ki//PICloQqczWZl5c21SObvcUPSojZnZLUISsw3Ri6zQ1l9P3G7dTWB5SQgpHGDZtFI8GosNEl
7TJ6pHrDe2b0dPtQpyDS9D5qYFv11Dc2ZJN5xyYTziYQhzrHeYBRUbNa8ZjUCAa36CIfO2fVIge8
SK71I9JOV37ye16kZ9Gfq115H5w8MNs3vjHzKoRVkQZghSiraGgd5JP0LYLR7poO0OhOQDblmt3M
CN+6sjOJf/ZjbK+uMwbwgET/SgovyyFImQfgPfuKkb+9WbRZRWJIC73s7yN3CgsxtwQ0jiO9Zj/u
zUBFpKUPhLf+JbfqlrnIeaUKdS7TXP7mDYmslO6Py40sgbok6nTn/3TaVuYrfn2r6oGjtTQRyGSs
vv7vpnuanTHZJWGBLZTFEyg6GcP53RLbFvvuMi91XEN14OwWHSIQwHGMHlKeDKveWHQb1gQwhf7G
p8A4ceivrcKf44QfLHAqfUrjm9EcaASBngtBDf4fqUWG06g0sk/KfZUZlw9cT5G3KCuiiJt+2lz2
jWzb3OLw3g24e0D42UqJnTcQ7a43erV/MQYGVQst+Cl9TY8trrIWJg6pDEsXMCJ1QAvP0RVDwRdt
kBL/HLocvyPimnIjHk52I3BcLKvXC31+HAGNXcrr+BDqNvvGfnMqkInxhpQlamCgS42ynLtjRZaw
3pXJQSZ1IvEh+Q+qLL2VHEU29vskhyrrvc2aoXa97T7Fs1zpPIBLWTbcimpKNSH76SuPj8b+ihZs
TbpmJRSfYdsLavUmkzfDjLnG/76LBEGosz4J0u0ogs3PFGt0Nik7T8eBiNXlgBpWGf3CUsPGlt8c
P0pw+FX06kCA32+6pj7e/w8qfQaBBct8ZXic6T1Qm1Nm0ntiU3DWQ3JpLrtFjMVb6kGKZbMvM+yY
1MLhprL8slvbOmI/cWw5i4fkEtRn+N7nkHK7dzZnpjV4UVv7YFrp6G8I2g+3f0EaewSnqUCtQfve
HgjGMprpOEFAAFy0q15BrTTK82xgH1pfb1SnXkSHm36qNLInVgq4PYDfh7EVKr+kWFF0eWkPk2XK
zZzXwye0pWGstjs6pg6rT5hMX8j/wMzUe129TILrncWHDMQ1UohyJ0gW6nGoDd1NjPZtr6NBqx+J
Jl1W8yLNVZRegxtgLAC+//z9YSZQbHfbY8oQaWQcgBs8g7cxL3i8XqFZYz9CLlsmYbulePLWDeXl
z9t2ZUSugi4+a1whD3X0fLqL7HudkzlFbJBdgKRbso9ViyOzyVOCk93fMNL89Sug7kVLA9JbbWSS
KbgUTgvjN42PM26qLPL4xHerKpD13nduZcqHaZOQUVsYEvMkaHaR3vrnblZZCyCzWYlfAsfFoD15
G0Y0RPE+K+p2J/xaOWhc4U8bTfwikNuVs/0m0oljgAuDs0Sqt7sWbj7yAzTjvSBEV65iwhN7n9CM
Zp0by3COjLuJfBBsZJQiHnPqTi4eZwz19mOEPL1RQqxAoGRH26w2CesIylADOYOZJpja1vRj6b+X
JhYUJYc6KQjqFUXQfVaz82GpwzMeGObXrI6YVNQhMSundeWfj3fDVbigavHE9QhpRUbWu0KOTXcd
4xLZ7kLl1I5qBINOc04jxpngW6QkkE/5X6oy4VzWxBdOqoL9AYPwpRooenETSmDaLwcalp42DnUC
MhhP/9Db2YqsUPZe+jquuDhEhC3WyZKBdjHTJSQrhWQLp0sqMIr5H+iuWdWuNM5hCsw2mBBMnkie
9HjB/azairSMq6OThz0WhSIwZI1qqnZwaDh2hbLh/XpQcrk7DzUa1OE/C36JI0f1yYDQkNASsbSj
f+RIM0LTHkWPt7rdDKK3vHj0baAD38gI7FdOsoueRI5bcOXejESmv97SfAob22T0OAaWOHt1nCL8
wD1nu+arVIBfzXCcTEXbN1VVp1fopEuCvHMoYly6s6KubGc65CNkRwKKG2JnLhSx/I00vTle3d1k
ztsjbogAWfC6H0dp5n31+LbttsCaGK6HAxSYzaX2NWWiz81bOZZzjsQP4ecXQnzqkxA/oVxhothm
2ElcdARjtkVbIXYuf+RdrMYMpxIi3HlzCHD/tbQ4VtXNGDuMlmK22/H9DmMXckTabFQq2H+BJSKb
FR9y6Xb7YafbNcf3G5dTsluWq8zNUOEmZtdf4YUuDvBOyMQgYc/D/RfZZN6sEaCIdw5visXlCJSO
+kU/qMmiQnrgsE8i1+e3GT/8sFp8feHYhkc90pVKPMdaZF6rRQKWpG+usANB3vgO8hijCIWc4Kx6
H9A/EryuShZbXOK+sYIvXtuQnWnxehWJk+PYbWS26bqcjtQoLZGZSgmPe5HBFx3rGtWYPH2Ntqwj
uDRmRgKqWjSV6M80/IXbvyCgG+vmQ2X9uPOG/E+oU6ehhbABhUc1N9cHUrCdl2puphBkWLRlmNgC
nveSxAUyqKcvWGbSyM4omDld/TsEY9kChH4lX2tLjaGk4q4LQ+c24HTu4Iwm9/OCrVolJOmM8zWE
8l4rJlgIomlcDz6LIrwYcEUdDWGdPJzwGBaw0EHr4hwGnbKH1WbNUo6X88q7BaJaV2HESXkc7dWC
9wRP2vjfj+5rxM6UZk2e2h2jd8iSDGQ/80fLV6wnwU+4ak/2btOMPo9IdJcV18ISNaDGWQyQlELw
1XN6DN4NaNoJrf9070qPadNahcRmyZA5tZp2vCFH+/k0MOx8mpYZOm1v1y+1A4JYJWgbmnPiObG7
h4dfSm1gAAWE+eF7v67F2FIPrk7Igj7Fronn8fLc5KG07GxoSyzFJ5UIsycKLhD9LzglhIRCxi9i
KaxhhJzOxJ0IgztQP6bFUzyfmd4sexfCA1eWk2ZOlFDm6EpZojlP48BMsU5mIOn3bEJieMI7JJRg
6pBBe/bdXeGWVOuxUlog974QiZ/vbyhHGr0X3O3mBeeljJjnKRMFeTv2WV3YFyoff5uyUc/vCYyM
GEc99q/lofvJGbcjxpGanIOSHk56MLU0GVdWFdJFhchuBBM4xzGMkqAr0P1A0QDx3mTpSMyVwpjR
OV5NBCtwOPmT2bpnDIDh7jdPbZm/3XTLhGPSrikorGtx368Di9MyjMhGBDwhDg6BZtxdutwTCcs0
8BBwCl6swD3fcwDfJ3LfYACyiMtGG59Ss74qC2JvENcaP0VENGDNjPQufc7eep/RKd6zVd6eRAhg
JjeBQyi22xvKQfeZLY1gbRet0jikx6VIN/gxEj1IC7qk6hc4l09oAuWmBetj/6gE/Hc6y2AURB3n
nUi+S7tjU8Oc8b7e/dUp3SyVNlATI4vn6DnmflFukSTPb/a78lwE4R2eBn8SG4FbfdwC4ILbu5I1
AnrIyK62V2X7WkqkeOqgb4mGmYsfwFObfvqFBEJOE2CDSKmfBLbw/Qw3uQCErWh6YkVU1awQ5Ebc
BTdGgxzrsOh5GolbeyKXnIh7YG0Cib2xPsUWXHWSI2aMsXD1WsdcA+3cOvogGGWY5pP2bsYzSCCo
/juQpKp2kJ/10fhrUL34ejtDQzIly/eO2bgrVugjjMZwN6DK+0ZL8fDUYsk9II+GgyCFV9Y4KxDw
T0eBq4peLFjVqimd9O9RpT8oE3GMLsxtfJvq3NgNmS8KMG0qHhUMkduVNZLvKsS4zmKAmHsiZvAD
LKsk5Ue4FyxmA8KTIVny3DByCORLDe2jG7lbz1bTZpj0rXeusbUafYk1sJUCXS5JfRieUERyuKI7
9i18IZohg2gse/HJAXo6/61GMK9z1YAqU6exozAcxDMlHPPjSlqg2ALFouZl0E7EczCGfYvDYfc5
d32BWlfBpQwehhX9H5nHjGrN/tTGyKEvYeZQ7ILxWvWcxpR5enc+gXI0XT9/vFFy8793qXwSv2c/
ToEPWjmJU5687b4hinmAfDz2uAQTW1jOALw2THgrsfakX6KML2qva6rI3NEY/8X4SyWPBu62Tb32
NH+an1fA40GNtf8COUXnek8cGgIJlyZCr2TQgP3ltOxJDR6+X2xvGkwLNeYNg+g6fVHxBpf46aLh
qwTE+ihkLNGKdUWaWUA0mahU8uKLtrhqe9Jf3IrWTtA9N/lArwGjvKK2sy2MJSikRwuK5FSlGhU7
UNAm29CTqF1YGIIU8H1mkul5awVbWN/Xv9248S7fkmUszj2C5CGY8fVxKNkiipB64fk8WKfxL3IE
MYm2L6zBi/7Y326agAISYUJwKcrIQ4MX4vfGu+2paKvq5GYcnjBYK8i39doq55s9lIRlxb9QWpFA
nsx8siiZ5sRvosGD/gwGYIhIXw+M/XHbhE51ernSXaD3Ru45YLSG02CGdK7ylZDU3xHmK4PT7eca
G2IQcLQQSugnWTjeCXyl2npiweGqSbQxrc4ePg4rE9gGB5UpRHeu8pfW5LRlvz2i/yNI3txjx46F
PalcRZ2I1B3jnTdI3DiF6oC7l4U41vCg/8Au642+lX8PtLED+w2SrzB7kT/3kgVrqwYq4sahqGsG
ZefaRsd60KEN54r9rDx3BFVvwz2xao9TAxmgiTKTdQyiKvje+MM8YZJtICYnMnPtTslJ26NlNqQ6
IPSA0/gxg/h2LRu9SAqFjPziLqzNrYM=
`protect end_protected
