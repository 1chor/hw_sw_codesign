-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Y83RR2smnoohquKoDnDAMvDbV8JiKnJHZ19EMvBiWLtSQS3MZyxsjMRTdRsJQQmv
E5skA9c1PnctTu8/E+DgMIsGmJK/Ui8nEoq0cNgnxhhsj1XciCfna0xyns8PhSbu
1QMHe4zFWcg27dvCxVHrug7r3iuDbICVHfRvNNhTl3s=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9200)
`protect data_block
UF5EgOA6e1P1Vct9fbfcRcEIiwFxeZiOp38rVliX9UVVFCpsy89XGhX+4zkB5L6C
a3BvSTuJoc2PBpRzhKdiRjoCiC9kQUvWrmMosRuD/0yrJWjmVKQELSb7MpvIfNEv
SAyKg4QcxEHYDxSZiCFvUunKsHgwtk6ERUbToosIZ1SKQEj8p3L0dme5unf5O44b
ph3B3bEMDTj3q3nGlPbeGn5AUkNfxk/f3qaEPqssSZHMPOukCHvULl+GJ9mmS/HR
HJtbatXawVmfC1hjXfbV4J0Bg2q28DgApa/WgCcyAnCsCJ2HF1vnglhvAnqkGA9N
dF5nQu8Qu+MAJ6eGIlvVdVMqXDadiI9PmblBKkEsO7qRAAuhSnMib1QeMWIVzP/R
e0EtKmIO9tEWZp6WeDg7OzcStdrcTCWT/vf4pNs6e8CUw/xLjV4HU+PoyFT50Icl
LoaY9JhTCqq7RftWbGZUvmjYOgBFPxHhZk1BX7sOaS3xSJnfwSfxe1bVZXJlTiGk
4qD+wkMo4U9Za3vjumaVlTVrYJo9UAAxkwN9LJ9VEUx3ZGlIBMy0+oR/62z4V55Q
OFbM225+ApfXbOs3j+JdoLijxQPzPQATCfj/VQ+/sv81ekKsWDu+jWy7fdVoGlOI
spti1P+V83WFH+NmeHB6f14DLGwvJNbVia58RyJxkkIetWv64bMN51vj16Hxei+N
b1vK2dthNQNQTjrU5KQonPbl46X0ShkwhGM5+OYWc3guIGs4OhRrzjkfYjRvSZWS
GyFWoJOSwcbOkdmbodVx+czIxYhpljsB9O1DBUz2QrRuurnY57GM0JK9qZSBmLCC
PdWAHyOgAKA5R/TFRUAle9mPk5PUYjeMpIlSmvZ//8yN/8mvPNJlpXZ5FUl6gEE/
ZAmytHNauBC0nVBef7ZvoyYGMi/JjtV2Pl6xDndG2Ae3lo3Op3wdWkvW2W9tgEJN
OrxRR4SkPghfKn+H6jlvTjtl83WiFFMWv1upGaRVQ1iHBhASdXOUB4Q0e4YxKicY
E0obXKK9XdYKgIWfztaEWUTBWzZDKX+aV0typYGEZ2VHnuEIfSdmg88/yR/u7O9l
grNyJyEZLwinMIZ0fSVgLhQS1at7F+gIki+PgNprZNuZ4K/OeCx+7N06oRi88xlA
fMPCTtreLsKMEoBVrPnMrs7K1adLAybtrnPg7RWJSMIRLMaKNpZscNKqYJXf+q8a
uAUPd5ehhq7teeFCXNFvPK4AhMD6uKw9QcoNYc+0rvpCNjDQmNiEfBKYPuZKuaeZ
YjbDjhhNXfSUzWMGnSnn+/IjvAditvQqJ5EreHSpMeI+CKSoGBdxsig3Gdrz2pGC
nIEP1JWKQOZxClF4iE6eDBS1tLizkNLa2K5p08Wf+J4VUrmZM8nptpOxaiZ0mnMl
Tog8lE7Sj7cp5qk5KFNz2W1NU1O4BrA9vrpU9pB2acG9+G9AoBMbUOl9wmm/Y6pm
e0qzu3CPELsJB75CB/diS7vUjfHteRPm5aFAqkMVlLry5AGs+kLxONdiotuVGQyT
NN2+a3zXZdR6NG4Sgci1AUGb2i4xY8D1l/D7XvJR3pCTNznR0Z4jx6AT4NnMp8GI
kuTD+rsRPS62vIfbRBjymABMC251bmSC39GAYHJexIyANOYNLPI7ptRf+pUz0z62
NUUl/NqgvzCxAfMzkAxlEvbwD3vka89C4SNUNAy1+qEU+Y97yKd16TdFvi9DqzFh
n9B3DA7K5FUhzRX6wGw2OVzVX6zs/URebsT9BswDLTBwHxKJIRnhanSx9sj/Vt/3
TW2ylZzqCXhMCw/GArWNmoDAbCWy+ZPbo7LNI4j0SBOxZvd+g+f8kBp4KNIXfukf
+rhQNUYuvDbh7RR80t8mvVmVEs+cokpO28z5e5SacOS9jeoYIwFi9qNA81I3FweA
5BGR5zqOqvlyvRbCDWyzkgPbU4/gumeC19fZs0lHQ3SIxV7m3tnWW0ry/rtnf8xV
WijWS5sbnHqDZch5RCyGwM2d4Rkgc0XtfODps8m1/7Mnu0C0LUaKvLCmhLl0chR4
4f9Ab550IVsy/blox3XZJs9ZRs2zI301V8YY89MZa31SWK8saoXG1RWiQ9lAup8W
SeraPBaM7xvG9zF+qjY1wiC1sw6kjHH7ZI338dWiSsJW6TFKWOqaqkg08Np/QfoB
BkxG11YuDl6GUxbPqzUUo7it6mWpyDTBXNRySZdYqQkffPCQV0yDSp0S6WPkVzi5
RARjjq3oKOOYs9R/99wRdnm3TYE268fzQWTRoijR4IMaS/ykNGzNvsywP3va8eMG
4EljNmhsboPZyu0rVCt6jeTcMBrdWnmoEngAQ6zbU0kws5bK9G0w/0qfnJ7iDXOY
9ePGzRj52bjoHNfDY+6mUV9AV/wVOP0noWTdVm8a4X+HVlqgY8qSQknlKI8MMu7u
2PkQe/67C9jCDX6zu+M+o+ch85fRP+/WvWhAywpM76j1rLRTeJfGC23nnrIq9m6I
PUGqXUap/8v/rs+Rf9TF6zqfCkhotZQdKrwseY8hlMDOY8nKlj793gR2EtKiwH/o
diGXpC6YJpxdbd0Tsjf0UqUqnP1sNkHzYsXtrEST4qRhNESyFpBVY4jIM4JqOa5Y
cuydi52LqBjLeQsNn8mndsLWBBQQyXCL7PQTCI7Z/YyErS0W4U367bOov9jyqFbd
pFIBpFybHsOE2xO+XV2txO+2j9noi4o8zw02n+GPSsU5XSsk/AU9DKBOWFuI4nHF
gz6GJEmjhPywkhG3fOLcdNNe8yHWEHc4nxDY2HVPTLct8UwLk4tJ3mlukXmED2vU
SbJ4VPI8cWtYzbWZVm0yLq2YQuw6IN7m5uVfIJIDLeNSt6mlJ7VrnpVIITLsfM01
2gnyn+1wG9tXLvpo1ROkQ4jEIo6FSQZ8Vt4Vz8I2of2UBTPQ2NB3Rhqx9ziwgtIr
QZDNsEeNLBhofwICxSCybm6FjsC6G7gsg2Sn2uPNadaoQEKKq2xwOhBKHrH+3pon
Mwdwma9UzMRTBFiD0mdN8y0/JVlfxSfjUDNfxokNL00K0PzKAu3oUg8KmWZ+Gnme
8kxIgf4/V+HQ5cP8oCWPLdY+mWBwOyLhJnJQHggPZNv7bwARKijkQFyjHNKlvZSO
YISDPFc1RnNpE2WF4AFQhh9mpMXOWkYTdGOm/uGfoVQ1Yid8IupHElAstCYgn5qg
CbmHPiyQYmpOQspePtphhREI05cSeM/P/NHWzak7/tPSL4D31XKOqNfPPpcMpL7w
yHfHwpD3fCgzCy1lJwL20zMLbYXsTOkRXv+iM4uMtKNf8g0RsaJ7Moxr8fTdg03d
0doWxwPNEqwv3T5L2SeTwC9zy03Oi8Ds+g1/7UfEX4ric7CHwWgY1Px8f9V87j2W
t8GGGthuBVYUca/1nQ6N3FYVHF2b+ucr+M+WJJ6aYmvlp+1fTs3OhYMJLF5WBd3P
WORw5xmweCg9x/dUmH6zHvqitqd+VnwOX/T1spoLmlWcM39HLSU5a6w34pDz61my
PecIt5wwxxWcTLIibZ/6jlKPX9aP326QVeaZyEJkT3VsvucU7E/Hmw8VJDCH9JJb
2KpddxqUOzvQMmYN2hDjkHXTyjWZszh6IjU7cXxFIwzdjJgKPSODCG329RtUGajG
EvDLZ+A+n2RdB4J4taT8bZm2inlO57SdjdIvmcOT33OsnHYwJm84Zxbm9dPEixoq
9eNwJCvNn+/HDNziaM5W/lZauWxmk0yTSi828aEGjNw5N46DLuKB9Fb+BPuAb2Zg
NGT2AE23wEHocwLp835E8NIIZizSmuCceqEA5nnipFDf/2tq996qWQjYSVTLA7XL
s07A6amk7bJ183h6UMN/NJ+WCP9R15PFNwHBZ68PsoaYLZXDbxbh75avTFxDQaE3
fLDtt0ARveQLSaXlsAkXwQ01YU0PynY0Z2djzM/T1aZWPgv+U2WxNamnQqBA6UZz
dMXbGBgTqU2JHlqKFBUKcGxceN+MK48vVhY+MaDxWBI+Uy6v2L9JQfDeWXDlMluL
So4u1qXb8XFSioIA9Jz7MG1bUePsKGdudlDHWks1/AuCsI6hfs56sxob9OcqiQiW
JnSlJr+E2hMJM2VTO2F/a0TEc4a5MiNiCmAS7cp6HYbnVHqCuDU5EIEYy4Os+80D
dOf9Q1cABbdXn+NOfipJeCKpWOaOjWr0XZbEQo5nqDDznNIXDrheqNM1/j4MS15F
TwOMJG89IAek5RLi+KbULyeCA5ekQ9SvY/0Ajoa40eKHNtnc7c5tAw4eawyj+RFZ
eYrLk6hVella8emIGdprdnpaGP4rTUZNtWIlb7sOWUHKOfcXhfwLaT8wl4R29plc
OdLFUUrYsXqRroogWGKR139p3d7k1aowCJ7iRBqCRMr5tuoXDmPVjYusIg6990hh
Vr4NHuyKfJz61RXUdDIlmjKD3ErNfBHj4wCbiG55kFZM/clHDXkrmE4soQX6NFgi
7ofnacH0n5jsbBiSTTiSxSMJ79nqlU//3saG6Kp7E+23KRNOTHNqgp8ij+eBFjVe
gXCv7CZnY25ATOLW9IoCSwDOnqtlrTZY0TGZPmHYSdQ8+aMdiwOHwe4RYzFdOXbk
bLA3VwFThd0VfCtkcLf2mWekxM20ki3CJgFCpw1FDpLP+AvAOikMUQOpVn0/hRXv
8QHuN+q9VtZ/qp/tqUJH5u529x7ps+06g6Goi1IMwm/4HgU51VjQKJjs+F7drOAp
nUZL/6WICACVi8o5a8APdzV+WmbaQhxjLcv1CS8V1Re/G+9NhDVAq8lZ+05eCqUy
C2mVTr13gM4naod7a5W/5jW+u1szSfp8vl0fl1HMGqb9rWgNzsDbj+5R4+hb63X2
7TPhh8VRt+p3KyQ5uTnevsDXuuZLVXxZTNLbWtIk4ZuRDiu9UJhycJ2bZXw4grcG
i8Krbp1cITNEMeYK3GfQ0x8SkQdKjdst02UoIFN04ooEYS687gRYyzn2QuJCYjud
KHJmO6pRn50/u4sK+nUNj0FEx7UJGFJiRFCgYezJTvN3d948D9UwMnSU9kgk/tsk
/PyWrf25/RrZ/kHd3maUQeynlmgPtuKjfgy3LTs299Ma1Q143nqHkStWTY1TNqHc
4URf4uDu6nqqyXzThjcbTiWjMHIRZ1Gz+HvrVFwyb8fIC7A22jANozbt9SGSRs2w
3EwECMS8GadY+kbKFPl1yCKj/AmVzvAquDyq3mXT7ssa/IYfzZVF4B5j1YlCrly4
QFqGaMiSba/nh/XoQEZN81kwOGBnJfiJ3JiBqPXsqFN84CBcXsFER+mD31+FS7Mn
pZf5OAGnnrTLbUEuKMiXVELhESgwGiYgwVtkvC4DFM6HH77IUhkMjek0DwwQTBry
EPJA+xnEkgjMyovLln1cI3k917vKDu0sHlHLq0gh3tikwc2gFLdEZx5LufWO3ApT
PWQE1Lq4pXE1bCRTJS8QAFRnOvBoRCXLmIBSfOK5bmx+u9VVxAgbos+GBH2pDHUL
XHohGwtpgrn/3Y+liE7Ecep5e2F1nKuvs0Hwvso5yt6miZOtJ9YvSxUefpa2YeZC
pDxGj4E4gCmG68oRSk8ormwibys63wHeFxHtiIN2MZ/9liQGqkHceuprvB+WmW2Z
8wzVsFZIAXYow3D7FxCn0vQ4GyZslqxWdbFrIxjBwZy9P7o1NX6YPY/FHGOSao16
bieaNsguSCfYzqCcotAnsW9knJc9AS3hXAHywVt9yentoM3uY3X0BCvMiJ+fb2K1
fjtkvbHARXyniEWGKFTtKl6Or1Rr49sMqhzmcha2opCfQmKRY8ThLz6mN1p8kx7b
ODFragcYeQ0UfxKnan8fELIRQO317y+OjLGIYNoDg8kYVIxp5MMwnb9qz/ho2n4r
Smr2Hu+ecAaueHfQUlR20iKUY3cUuzXUE9oKaBUt4r6Uw1ZGxvpSAGcWw6vwqeVX
5+O1Y1p4WHHRBQLipDNA2NsZMqFewAb6r7c6G/r8e4ABLCAh6Jn8n1JgUUbl2COE
WSZAOQ3YlucqIDdMpZRjRvTqoFggi6fxKvtAyU49XL5ed32CL5Jwr3dkqBIH51bF
R/t1b8frxNGCrXCh8ZK99o8hKFxRVohyxJdQ0IvP31+WMZgTl3g3RgBPlo4V3/DX
a/hlx0qLY6ov+l2Zkku758ZBR2WMQgZplT9klaztdptCT4IzS4nWI3TAHnYoCxC+
/YlkkunNxX/pMQGMng4JV27JF3XrAQkEx8XzkqzpLKE+stNHwYx8EYYcRTymcJ2j
J6emr+mkhOO5LaeEXYLo/OKEF7NdZT6YX+13iSqtAi1Ae1mr5esAXwNp1rSruEKj
odCe0N+gZ2GT1YOYoFZ8IlT7jLwETBYInflVosI9G95Nl7urXrIJK1gwLWRwLEbI
DuTz9kN0HtvRzX82lYiTdBlBnX/uhbvPEzPAG5E2+yGMeVhsR/7g2p6IwfBI1tWd
Px+4RWNAIEk/7J26kl7N6gF29qDzAUNs6uUjhI9k66P7xdG1vc+35J/flzKbMTby
5P/blWL5XR8d+hYRr6vQ/06DfMIsafKIeQN6dohR6GDxmenZqlPGFIXGR+O7H9YO
iqBkzc7p4kueq0ZecAz13V/CgcxY2bDFaW2Som9GKLY3ML9bdsnS5S6pwerzhFhY
lrm0CWGSc+3R0ZOyl1I0Qj5T6xfpMBs25iLd6//FEt4q6Tw8zRL7+COljBoHIfvx
N055f/Yr75CaxyL4CgDLf9JUGT7B3nT/ihLni6rIo8U8qB38BSN5N9ZrJyk91ZDF
SmE1yfkhXqw1VaQpPH3QeB4IbCiiP4NNUTXtTn8TqG6pfNSJ0CP15PVJhM3LTXDD
mYtbyMTRa7sxH//2Fv+XkNs2aBq+wamO5MJgj3hHGOADE1DYqk5XnPRHgv+dAgrB
P/ce9ftqqZxt5CwlMumKucxBTen7tamJmOL9lMAg0sWgPFm3ex3tQyjgymg980MF
G6biPHBEclpdptfQpkFdW+84pzIz+93bfqLRUlEKK08Tw2nhaTBrRG9vLd7AMqTR
6qkybQnPMdx4Egn1Ztnd3YNnvyoW9Kly0USRkHdE7gUoIrs7db3Vmao+PgxY0dhF
KxLhe0iTrTsAzi1Gju7pO8KxlEQledk1DCKFQN9Cte7OYKtoLZI7YtA+pajaCkEe
QFBqiR+4uKrWggDUKsripn2JXdpfjS2rNxHe6GUTxm4mIMv+ZrUg1AWSDxq9WpJz
AGth2ea/MXDZqKId7okL+3WhGygWDLXLhQpiiPioAEsCLfSZtK0hmpFNjKdSxm7Y
U7rShuCLEbNQXRYknFcLe/wwKnCDHfeQFD4opqSZIgZC5gCNq4XBf60zZWP5jEkY
+u+MMBKPaL5xDPQzUClIXYh6KN7t9p/qwke7zYx7HN6JWnNxKUziOmAqk+qqnpzM
c4j+iNO/lmr8F5xuhZLE11uwMK3gQ9IYZONfQCOGLqN16C50PrmiCkDIsm7JQu3z
xohCnOrGpN83GeWFe/4/FtjpmhKPi7z7oWZ2RF4i5xzd27ewrhmBMSNIl2R3Dp1N
r9F+IQErzueAVjsMUgyp7yBDva9RUB6lNfOpJH0gldlFm7a9HJEFaqWfCjn3F2Q7
EG/eUcRvlbJl4Ri4nxbD1NipD0VrQK02UevyY6OKtBUciNVhvY5hp5NGFQjeaXH0
q6v8jsDjZzO1NNc9i1xZj32qevBSVfadimg2KDRoiY1WOu6Rnv257DCIPqZJijpp
EjFTG7j57tmwXzB16TXfhoFadPvHCxHVkzrgsT7RuyfmclC9Tr05OoCiM5BqZ8QJ
4Ffku9Tc/GLTaoCPJrr2CYRWGDwRmNRiCYz90CJh0k2Mm3gwX3uNbUp3qurqF06O
8tSNPed5cccNodcMPorFEsdcKVDgZrv/OaV4d/EHBfN6/Zw/j/oeTeHa2+oy3Afc
tI1gSPy/s/qk+p1I0K4EK2JyqQY1no4dcwpECp/WnBCoazMZBaEfRMLF/DhK+Cmm
XkLFk0u0tzQzCIHy1r84ma8A+GPArzHUKq8QwxFCx5UlnaVhgNGL8JeS6NPtUL2q
dvzSBjTBmWM5NEDB3e9lRceANKZ3+pFmpCzgh9kC+KdnTnN3YZD5MAsK1iLAJRKE
QCldIIk4xz8H1Jv0MeTtVJT9bo4dv6vfY3FRivSzzB4U1mX8RALaN3aVNzAoP1fA
dBUhw+pEhI66KQ5qoli+Us6zVoe1bNmlv954jqRdonZnOxRlP0pr5caDpf+d7gj/
/P+sog+IsKxSUt2fbnMdqWTSUL1iCBsJH9v3gHFO4bA9TCQzykEYY9HvxjB1y6A5
AZrjV5YYI4oN/mL5YRHiUbZqr9dMGD15tS9CtcB782vexdG+YvedknVRqR+W3y+L
pvqag/jp64EL5BYfi2jdMZTLHLpEiPF0v/2PL20NYrVSCcDsqQhTWZ9gPxiwR2V9
sJl/GV4PriKgfDBwcbz5ag0Ih3nuvVmzfHRWA0i/FPROU8TKMQiv9fzcto9BoEIC
2aXvAaZT78kKsxpRCp8WIdDFvPQJRzSgnxbWV7zfh9gaX2HveZyUrae10PIVXhut
g/Zu0ICRiQ/D0JYZE8223xTPZB+9ixngPt1sQXq6ywpev4hOF27c/IKOWgkE5qoa
QzmaA8TA24rFEGg1xdssWp0Kt6drwhfrdZpwMTaCqLN/1VHwgaBsrT2jPgWO3Cja
GmDzL157DO7EmEJhU1YdmH3le8QnV0I+r4hpQ0gWuMhsprO+/HMlHXhpDZgDtosX
5ruPa1LxRz9yXHfUu/9ONwkPHF8UewXVoavZcP4U2hFv/1NsqPGIHdOsmOQBEXNj
+WV6EUP1IcsQOM75PjaeiqxENYD6V3CKyMBeJ9/e5Hj1wDcXb7AZgYIZWnMbFtKl
1TKMTBrYEL8L3TXMRI+BvqlbjPEq0djFMIcZ/lhkGRXc8DWWjkO1FV/kaMGObCV0
zD4+5c0V64/GR9kpc2oEzYAsnCe3mOPAT4bsStGx7j74PBeSr7xs8sBk5c4nBEyx
TURLopSe96gdOFeTmWLClVc6C8TO/55257kMGUVVcgU0Btv5VCwVFDsfzAkRIsP9
olVpGZFqU+OlbFDFqzjOSiH+Nl9s8ccRcqmmRN3BYUPkfB8EDaZKrQZ3gtaPAw98
u77Q/UpCRk61T4jRVzwOl0XXlCtfwfdKeohMLYBZaqplpV6F8+BclemUptuf984x
p8JfPIOaBGNSwLcdMf6jm+xxTm2yoygOLSR2Qy5BdSvEYJ5yUaS2/j6t4ymy48md
cEqvyF5xMW3GK8mAeA5iLFkBfRSCsptCzZsngYYRiDThbB3k5Z8QacqmGcBsdLC7
PopluaSR5JPJ0bZDqJFthv7J4laV7mKESaXwjP5clO8NfTs76XV24uG+s0cyMvrz
VU3LpnXbG8iTeCjhOD1nR7acYYiSB3dM1cMMgHPGrDHuk7fr7H6JI46d+jLmL9jh
z4cQtOz8FOKruir9TCoVenvLlR2Nil4u8wOVSeRFZkx5oz8HVkEW1khaGdx9l2h5
i7LsFB57acbIMuADiRkZu728ahLVCe19ADC7nvCxXJnY0DQzHoLKA5tS/u3LSVb2
lIYW0+/EVWTWXVh+qER9lJaQ1E9f7bl8DmzJPCgV++HlrY9ANfxuZdHvAvA3Taqh
vr0be+THMCkhM9nwBmdZ3PgAqAjayDcmbN3HILLiNSYk4prkGAgwZZGK/UGIWqW+
t18Ad/8HBlVBDH51tjT6p7AiRcCKKQq5DtkNgeqyNuqgXqNQSqvwWtjFBqikjS4B
rhkz9dImKABCe6q2du/vkDF6d+O9bqfPN7MABeoC9NRjzbBkUoyPT8RSN1t322sN
usXKWUGsz4tOBaLSyu/Y/m0N1CVtYfv0wedVWFrAk6GB11CfoZ3Por+zKman0V6i
ofDhkDBYSeo0fJsTnR79JBkYQjvgMozEtDOjmsvfnGbQ14kDSAN8TsuoiI3FUL3F
cCnsX8teHjmNa+EaqEqA+jdhEdy7b+d2cdQAnbAmc9rBBQOdhOvKkTk/CUChL7iw
qtux6+zY3mPiW38wIerN4iJM0bztq2tDzEFRslrxdobvQ8LedR98mKRKaS8mmfD6
Ai2zfQCvKUuJ0AVMDI6zlHgRao4KFyV2qoECEUB9hc+uFZa1uvPIUjYqgjzXBs//
CfffJY9CLu5AZhDBhByNwKqEPdPOk0k/zGZ3CPAJHbduwt/4SFB2J59kk/1ey1nu
doPY1PqJh1xUwX7qK6K7jJvHTXyRzUedtV1Sd0/O1A5q9Owd9UfeN3dqLVRVtx7l
Uwofn9tHbjDNKaP3VkZRDG4HDW6A7gdInu2MqkZehQe9oT2VU3ifZYM/jLFuX0oD
MR/LRk6NO3ZyBC6S1VWEJC9bBlfY2z4E7lWVf+NuTgI09Ez5AYLcrbMpcXg73egm
EGsMBdCwKqd68oeHIeOUgSboKsnlHkaVAj509p5Ykh0nZQkJED7crDlkueyPZY6H
XhQX6KVwnAR3tKWMcblYDUpR1eCOWogLKO9V1Glu4snQTXOVhNRB4Iwlj9R4CPRb
CwUrWzZ0o7qMTbphs4jlHUsoSlGue2WX40oFmp/LEX3wnNMwVvJrugkRdyVkfz9C
/mwunWTLKXkqGEucTOTK3jdK223MGk8joLmIx0Jj1/p3mHUSmqFPonpn8d4KoWEh
bmpgzwcZtrAA1OsZCJ/dfbOomFN3R2EzgYWBc0fgJoGNaGxI2diBBGdnoOXwxoEj
eRT4dYYv6bR23s5SaxMVtRwaiQvVikGsJ/cwI59DQiVYEn+Z8+6w3zetWWUHT6S1
HKRzNgcoFQ/7SGA+vsvWlRh8kGUW8S6XTphvt8RI8bpucRGBwVIa0PW/wjNAhvsF
hZhKywL5JwPepDaT6jn5cbwZLej+9tzkqoEyZ+AO+LVY91e2qHTSiXCx/ycr9E/z
xhXI02/SrZF2RNS/nb8wN/VJjxlceqUAqIXM4PwxemF5hjcGLzXer4AsJVQvwMsU
Rnbtwxw0Q4n9HktZCxF076NPJwSDf/aZCIw86HBF9+BG1buvbrsuh/mHjxlTlnxZ
YznvWJLuv7TJer+pQnAy4QTItBSBcz5GES3j5yhCPMmUvzjx97yXjA6jQSss/0WB
wkiHZSkGUaZkjlSn8G0sksXQMxiAyThNbKoduOMo2R5xRIt+AdD6H4m7wA5teTsK
sZS4eUcsWPsLCbp7Oq6MiReM2/Uj2f9WtoUil/81EDwLk3iDO+8Igb9Ha3J9RP30
nFyXgyKJ2/QlqiQZGMQxkus6gUIM5mH94N1X0SGCgqJJzDhHelLHXRhg6vcbWLIm
jYkS4z2LgzfIr0xQoHUXaZNiTvPb/FYfAYHQ/Cd36KBFLlwC3RKN6RvHwUWr9QAI
bKZgceqzxvss0dNVPzt2BfLVto273cbKoCo3Tu1SS/7HCmgdBZC5aR04F8yVaoBK
xPesA74u2PJq2YDuYAErIydRI7kVKKe3MIs33ACjJkHHY0Ts+i5N8A9v9UnQAVrS
MP/Pp9+eBFFTNwrGm1Vcl8etuWgY4Xocfp+sCI2IXz3vEvqBp7YbydRIFca8oXe7
016yuO3r1CUmwJo5qflGkNMgWiSSJ9756CQntkWft68hwLMW1SKyEng40ID2Jl1+
4DtbL/+YBqZY3ol7BfWMqYjulgEngk231lRF2WhulQAMgpabpc06mDEf/98Q3RAz
4uAMITRc7RtFbUnvf1jUWBam0p6xPyznXEKTnAGA/vvPyKtkAk3qNQV9PZou/Ld9
OfpDIFKwFituWhjE5UYNe/5ybCNZVT8LzIQmE/MjBsj/1MyCDKX1MokEbNriMpZ8
PRLralrjN0TWcPFuasv440zF0E71HD07IDbYZPq1MQmFspCUKDQuZqwK2IqmjGOD
j4MU7yIzVbz5zZ8zZwl/DMQWp9TjAkU3Cs6gBBsRlIh8m3OS0o6/C98RYj++vJww
gOKX4b48z4bG0qLBds9f5mbFv+0kdgxLijJ6gosHtefjziUJgAfDoAKUErqKK1kM
/ggDb5+oTxSGI40vaQLQLLyhj4rUgJvo3vrwbsUjTbrzs7XyRQns8DtXoq8Bu6V8
9PSeokTS8gFMmAjZFbUi4Hnn5DobRYVa4Yt1IASCRXs/9F9hqBZ/6Ly/H0oSRGYC
FcBbIBw3TfjYT3mJ2NQEGbCEiZ23HfrzP0o5ah6p62iNT3GRoJZuTDlfGKlQNBuU
hnULtu8IeOsAqTuyIEbKc83dHQYkeZluSGRSiAdiCps=
`protect end_protected
