-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kowC5cTTiEpSxqCDeRLzJgnMcrMxlwld6SXwaGgZ95UkwG/gnAldJzdj5DWQ42dJ4Dq32mrRirzd
PXGyY16t3ffugTa7gMynMfKa4E1/YVMYDHLZMpEm8tgXxJbNMSQSNXVx/ey4SO/nlGca20j3H3SC
SUO/YS/E78ArW0OMcXsHr0AnGLQGABAid9FDCKfJeTQMmq6NaZoDgMn2N2Sm0lopommIZ3uGISQp
YTwvkkEpsi/kVaqJZMR1bYmVwkRg5M207zvExvAR0ID7Gd9LdK1cBx64gXKMtybjsyBQdQNNJl4Q
0MHN5k+djUlyVn4T/qKo9gLuRXL6Keze2BOyEQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10064)
`protect data_block
6SYEIPG67cm256Y2bNl0fCpmqIK5n3cz8TZq+RsECta3CNEGGf6xwzeoK9lWdQw0Y0G8DdBNLBJD
wzPWTRQuoj6MuuiELScrg6/cVZRJ7kDCKgfLhqKOfGm760G7FcWUoDSeRfZVcPhJErXJ97yQbUow
JZYBfck8QiDbbsZEKp1gsFsbTnkNpj6HZKl/SKAT4ZQ6tZEdbqAISuKM1X6EJgFaZ2wWrsZXS/7C
snzu5g5UHhqs1w0eQI8m07FcqSnJ9PNAbUp+7zPJ9yt1iU7ayfK4ywrBQH5jnhqNWLQgYyIEXkHZ
jjl63TEytNU5QcPdl/IbwEDhKkNTzzNSAHTaWkIAYpKMQ613AZfOLnHNu0yKOnzuRXZugfvQMWro
b83kuWs0SSBnAnuxGCjA/wV8MaaX/KDVvib9ekzrf252OpgePrGsTz5V8mEGmJC2cpWRq+se7HFg
P0uU2MbhrZOzqJ1N/o7wloAEQ2efjVGXHFQ2QY2U4FehUY9igXYWOaAsL6UOrHs/qBwDeit51ppS
+h77WwbwzT2STLJ/YipvJTUyPCqzu5sYfdlGNsDbn7FQkzMn5C9XpxeCbX3tMxWus+HnRPrHL0YE
Z4al98bminJ2zPi5KVB7GytsNDXlz1EK36pntdsbMX6jpUUV8fR6CGmcoxBQ3QU7pExoczvGlRcy
6Zi5z9dyw2FPFXjMCrJ1MH8eNP0pLM1VkiWqZVbhrO/VbgXK/IHxUxap0oO+TpVfjM+W5xwZLr7r
GMVqO+lLpHRsNNs9AATXiz10Q7thZbvLwHz29NwLxiTlJY48i1SPQDMa5ACgbNnap7WeKXP0xW3b
rUJdShtmZ49ohTfpDNnsRjO7UV/dTq7jLsO/n8gz2OIoHIxRQl6vwSxpbHZt6wdZpEBRwvBq9Cg0
XiqsirOe1KRjnX5tj3JM2ZIxbfHhXCeNR7Dv+WORONxpJO7YPpEujLjm6g3SC4CUv1CbAPZanhbx
ptaFHOXz7Z+fGLH8B0mC5rG67MtDAuSTLjbUdUyBlmwD+hLjvq97if/5F7cUAH6gBZmK1chQUjft
1GZ7Fxt3ncnq5hphZ6aUwK4d02l99i5NfekCX7oBjimQaJ1lQplKoP/1doOIbz3q27quY0IN42jY
nHXwJkLc4TPROnvjaBFCFCPj4G2y5ERjsHwiO0bgvX8xwDQaeU9UnK8xGz6odpA5R17PnFw+B9M1
GQsmFWO6EVYI8g2UoAaNJMYKqpiHARy2hlnBXwMvQ6yVylkVPflcNC/dLvVt1Ma5vbGHLfdPZFU1
tw7MMcs2QNG7FWU/l+LssfBilqPjxB3Bo6MfnZW02nqp+m8nTIAPj3BlWqtydvIi35UkgH/cjiD6
aDlkQYdEUmAC+btvnQit0B4/JBuzZ9y/nXG5JH2lVG343lIlw7XEojOzP3vIVEaN5DC38M5KdJyX
8nZbg7aOymjsiYjdmSEidgLYrqCFaQ6EDI+/pfoQI3vocwk0fNdn4vJ6VXy+eSUL60X2P1+r/uTK
EKuwgn4XlhrsfrQh5KkRNKuScBjtmx1lKhq8pEe8M/iCbDvcWqPl6prwkPTWuAgPmzvbhEYwmaeD
2eoasxSVD06QMYXI9C7sJo3H8ofBgsE91ux9Mhant8qxu0s1dUUSgAJnQxVECEzYWeS1sUb55thS
9zHDuWHwjphKxmb1iDIKVk/IwLCMzLLf/H3UWj0oGu4d570podSjSuRZaoPNNBxdxPwwB6LVcEu+
Ehpt2QqvIok3L3D+WbgZbzpA8PE8cmqpwRlnkfpcqzVjajCfTHwAOw8mbcHe1cCdfk1AQEP+Lyid
VSSF9yEPGgbJCpoZnBg0PuDXTY+R4tSrOGSVL08hztjvoN75JfkxiioHAw6EgLmsjv+L5kcRiSKV
FANQWhTGiK0Gyyz7Okd7/n/9gozHgLEMeLAE/3AbzxAEXJtgZrH/2SkVBnVIUlncuOFuA7VchKyI
G6wU4NuNXxhPr+Fk5cGWLpM8/p9vKKfYGHb+t/loo8l4wKJcZ1B4l0EOmsdsye4fXBoR/gh/wuXp
16Jp0ArCxLyQ0M3fm5JyAcw28kRGOCI+khTR5L0+2QRo+qNGnyXGRMwAKK0AG4/DdZllwVBla60u
9Z1QllgSjoIK5GCJXggLynJhFh+eSMVdxxwOKYbyJ8DiIT1Qqnllfrb2KWvvYzH6YItu3OODdiDR
dvkLfKZZtZDjUh/cTVBF4ZOr+U4F+Wo0C6lsp1eEtAhx+nWpnkzpDkGZFLpZPqqfKJ7bSVMdpszX
rSPTwvyEMQQSAlp9VfREhj5ANWF/w8YEtr1c7/BIlS+hKhp6xi1P5W6WTFCmgkG579D9QVqkeBvv
o75V8wCGH1APBds6PdFHDh2nRQKhN6A6cZBLqY3QpvOfv9jGLnqJxSAnSz6Eyj583u9ear0GpmfS
nnUpwJQfy9W1SKkdSvpydKmRSa8Io0Q1TSoO7TlRrtEZh3pxz8rw4fBq1v26mYoHrr9V7JC84hqV
FT8rGnAuqITLdi69pSoEyx7P3Nu1eS2ajRgEa+TtAu2jKqX+YhYn/8FJx5bBBQ+4VZSEDv/EqBzE
ddfbJF5vKBi8H8AKa1tTc87vvBXVty+CMSEGsPl5iyHgsj114XEeVzky5bsIuOh6SJ3tLw9FKIYS
TEfwolkZ1SarB8kV/AmK4g4DZR9Q/bCVZxwxjtomjEKB3/v1PF7E4gSNFyBghr8YI++RBZjFKPbC
JbMHc8HrLANftnFdBMzyjr3sNcTtpNCYgwMVgRmbH5WBB9ErCpIQI7oYTWTipBJyXJx6HWQDvpNX
HkxqAwvN4YXV8tVSRXZktwgIV339IfpL8EFdIlTibqx3FS/UFWjXDY/BpGXLIW5Jmzl4Araqbb8O
2r0x9j50CKxKetPMsan+1eI1GOYn/iZ5BjfhuFVQT6HSw4xorJ4kit/+fFdbDFqcWR7u3WChaiOm
HmKmzmc0kVbWih7B6GT0W2cBP+s+qyEwNWcmtioX/Ohns2UVhLh9c0sRnnpW1vvKNh5Xh7JcCi99
2D9Y7PnblS7JdTNl2ySOXy07kXPi+d9z84EkXoOYd/AgJI8obWRrP+2aJ4YmYnANfBOMMILGvMlZ
it8X76acPEQuq1ZwlcHlarbp4yju9CPHtPfpDOml4Ic+TgcbixNqD0q9EROgFrScnvMeLDDME7DH
JP8iPeFFJdTZ4llN9hkgIXufOA7UTSvFZ+FiTIdFrTuwgsewxyL+OwMwFEGJmLXFicKVoVc8Yd2/
RAy63w2Lvy7BCieRwNbqk2rqngaJATPTara9RHKLUCVa55Sf0BhBEb4bJJmTKKUS59TVPaHHm179
rhpxuyvolJGtp+dikUw9LP3DcTP6CMalf2Ktg69dEgLtF5CMyYKyO2DShmTrSIQ8EQ4tOzLjvoIj
GxHpz2NwcNoaeI5FULQa4CDqG5CXHZ3fpMbAF9TEAeDw7pIqOy9OVUY+HDqxmgxoHegKOcMTm95m
QHAMmfyZ9KLTme2ubEMLpJjvcTqmKbpHhhvHDQ7mwXgXT2DuNTuB40moS9jDyqCUdUZG26qgbopc
aIUcq0U3xWXdtz+zzPGCAok35Cx/gWIha+5p92jtSQCWHyyWE5lFvL+5QQg3n1M2hKbvjrAIuR8m
0j0ZJGbQH7xVtNVpqm6XhebIjBMSxMiAXLa3QtPxvrzhgBwgudx5lU4AzpzjDMVkV7wtF6AcFO9+
X+ogQkFPTqlGCK7TN0h7lZONK5SDL4gDBtl8hJDGbbDY2//3tHrkn9nfB94UrydTEwU1mQvHQ0oB
rH+To0JDs9wGYoe12wZ+DBNDp5t2PiYPvEvNldaDbFokcoxob0fAH1+amDw6zaHVCe4cJGMBSO2C
kkXGJCm0I7TbawH8tCVPm0ukSzD9UjZ2un11VCto8B+30zi1hCz2mZdF+ebnhCo/X1WS60r2aqeg
sIdfk9Kd6bryWwgrHrwmdZBEEKXmoULl72BhoqDVYwdKJCjrUzLFbU/BgJAQpsixo3ShHn8/E5ms
Iic9DeNtL05Q98pH2JwGFRfH8Nn+kUt+eNIq/Jg/NulOtH/evp/PYLUyAhIHSJrfrzuRSvUSW+MG
zCtqaq5E2DBgQ536H/lnnsdyf/YELHi2GAi3b1SNhwf5LqTYhYZsUBbMnTM8zQ7N3ttrRfiuhcBh
LkauT3YXRH8ww40VGmzVC3nfpAxeNfmj5BYB5YfWittyJZX+LgMpM6/dpGF4FLg2mub6QcBoPnFQ
zK3YeKT8bBLBCfC1shJ5NlRW7GmH//CQ+wR3WVq9j4nB05gxHx1RlZB6DdiE62qWH0pmrqWPZkKK
WEYktmjIp6IhZJA2TWzkU4/2kbexgaY1q+K2RocY5DaqK4jS0afqv5BeKJLSSrK//LxBboTTo7Vl
dRcqdXmt+Uevm+nw0ouVLHhiFEZXw3ebq7MqOvcavg0p9WzxI1UnPIyzqBCaWKLuhqBiBUyLm5QK
h7cZyrIHxNC+8jRLX9zV2JTI5cnGxto/ds26iXqSXznfAnzmLZrCswf2MI9NStfIGeU2gLYkQCuc
AGgytTGGGaO/D1DMo+w8xOroRGSMIHjWJu4GYFeJJdksiYj49wCrv78JNiKoWWO7StCNZr0I34hl
eadrdVy2W1nDKPTMzRwp33DNYHvT2Btb3F+yHRFz2sdPo+QyW1z0L9FsG3UswI67gYq2LwfAKfh9
CJG+yR/fj+ElLk8gR0oqQbfiY1HdW3BU5qOjJeO0XhmEUXNcjvkeZC/y+dYFG9lUZONSty0bTTwL
iH6ybrSZDtgpz9v9iEKiCpNsWCvaOOsb0on78o/wwisHchgp3IcsWou2kRYIvkg33nRFzB2YS17f
uJ4WnWCvfBCFeBucLY1VtV2chdEvtIKTspr2gfsBIrqQLJPoviOK17dNyU3Zi+TZqvraYJr6DcJ5
V+qESCjs3lXFdSgGMksUyxH0TNQEUO/ngEShp7FZOPa0/BaT0tGH1IcmU878zML74P8kwo1T2QpC
Twlxpbj0XxsBRkuL5xZUtpdzcZQY3VFpfZyMiwCWoBX856102jjwy+wZ3RS4s+D1iin8DNxRvIPZ
NcQy/iZSMGr1qx/xAh1Y3FF6Q02pkYisxVaGqTBk1uwXTlxc7fP1rYR9lTzihddv3LLnsuJnP/4f
0vkmToPfumRwsQd4gjMQipn1GY4wVid2erqRJ1Xg6i2qSzy0nuQ97rHcuQj2mPrYVZq+wk5GsHgV
9zkYFTb7K7IprR10rgtm1gdk0gRFjzt8YjNKmruSGWIyL9AZKg5wmsreX+sl1o8DEII/hKF536Ly
n6F5QSX4vNSrEfU9g2CSCs/cGriqtqPdUNpEKFYGBiLHUwgFb27r6YiZgsKC7/+/1m1ftaP8/sVR
WH+YuCAT6z2Iou9G9cgE3JJnw1WmrQ4aNCU1jurcwLxOcuTRroEIE2EoMfllVJChbQcgrycYMtQi
FbY9t/HzMa2Q25oIS8d9JYbJHZEGx5jqqlb36V6XLaGjUIVPHLgf2Nz5eLENAWJVPCeFyei8povM
aKaw8D8IQmynBcx218PdrpAk2cFldQ7aE5qWrmipyhRACndvSKryqzcs6/6PlDIsw1OBqRGjLN4w
+o6aqJaAm5sKpRa4Fbo1MaoL1orKvuM4AI1vMRqs6oReXsCL6tJWZH9/lp0PzIDW4ZXcPzZBt9sQ
J/8I5AgidyFNM7JV2yaiX4QKPbMjoZndSAGJzZctZxVLT2Ce6uwm4zMoQdElHujM8VVJKRSopqOR
b+64ie2E5wIpXE45SftlQeISeak2BXjJLQ3fAPpYgHmOe6C1frtgC03MFqffiZcsTGWXQ87BSemF
LTma2tvhPa1+7FlpynPlepZ/nrIIVbLXrZxTz6IZHW/btEwcjSPuQgLNfHVyAZUhfa0fZAwup+2R
groLtpfjlZIdU8wH3reiu9Iz4xzJR3w8JTeHd6+9hqzaPM0Y7ocJ0gusSXQTmKvw9Z9xOAqqnp8X
a417NFpQqEaGavcHQ0HcPyPYylTVEvOTlE5jOK1sd1ldgAD44NQ2lHg/Gc/ZTqGpUm+duKgW8jGO
JJmcSx5cgXtEEUPB/dqk0nqJNAK9k+mOlMqZMXdyrgwIjY+pzbBPTOT+dFN/9A2/vEopYj7dejgx
liO9wEdzHmra01Fa8C0DnlceK6n7hVLEqhwOxwuFs7FexQPyMQLt+PgOGKU1RtpZRX3l9gxOWvqL
fPeKsDq2y9Ie8WfL27KPtNKfxmWqycA6bgEjalGft/6XHnJkPZ/0trpTQMk31Ar7DXA/Xf54yobt
jAgTTfZeL3zx6CvohoG0zL2pU5Bvf6ZTf/QbIRDueIR7vaMwj0ZKSCsBhfWlh3si49pklA12WVdm
M0p/qgKXKn3ZDd7RerNmUyQC6Pb5QUl2jJ6Ls8jHTVjRB9kctizbNcdgZXZ/21x57VkTiharVB/w
7H7Ptkn7sArLesUgLR1t+8VgyO35aYhOKJLTduu4OCUPYAqMRQYwFSi/q5f9izwhUIQwX2CuEC8X
re3B4skN63l1BaqMzsyxpeUvsY40G7N9LoVgzZkstyrG5PUIUS9A1yYDsVUn5U5A6+YoJDLfQiFb
dkZ1m5DZyfj0fIFI2GCUdDYh4hqi/7Ava/WsIMObtF1ZK7eug8X1xFkPsyNyNf+QP9QEPbOy/ztI
FqQYiqxqiSWG5Xh6XM7I3LWbAyRpPkStXfX0DqVKyc3kiKdRrhUKiJuciKEd9RTLNqTzU+Xl10Xs
/ue0zR9srAw1cUs/U/RRP3X5ZOtsHU0sBAN24fsUKMWgkTAGWdtZQ5l2bPOEqAmwIdMu9CISRXLa
R/KwZs4pDDSfdwm5nTYsqdiGilmsCRckL/eVD71uCXqBERaIXmH2wNIUpHFbRZhnrH+uI/Xe5TWi
ufRxJ7SJirG8ChAOg+w2KHP3mQM0fjvrsgLMifaEdox8WcpamaVjJY3GWG1odpH8i9T/o+Z07HGq
lKWzZjoM8kV6Ev1qsr1b79YCG5m77ZEIEneHPedi0nJBv3nJk/O45TZ8LSp6IHQARa7bHHG/gRdD
31rZsjYLNgU+GdpqqzWQ2w/z6SNW20kU+5wKfvVBapwInDaD7U22dZiHpdgv81ZJkrsQcAC+QXvw
ZUG7aOd1HrgczbrybbMV1P+KjJ9fEhqb6ppIP+qG6fqUkyruZa/l+ElVesBJsAn2IYCh/J2cS1ZT
H58yGuv5dIO3jRdPIBUp7FGmWcRSbI4Y73N+kZUpTCDP4xiX08QGXFPhnwotEnCupVwmZYzgZ9Rq
rU8wsAOA3u7nUvtlUHC+2mhAx9c1qObxrsvjV2l7N92qOKDMVk2Iln4BoZrtJAaOf5c6wA0L9N/1
MR29Y7B6P5R87Q5uC6n7sAtHBtArAa4aF0RvMkaS3a1DBdVS8T0BPBkmEHeyhroaVLQTtTdWmq1D
eS+FhqoVibiR21z74X2bOeWnLFjCyTUAKhJVnmKE8qaIXyGITxeS2PeDj5JsklWWJBySHVtlzr99
YrJKTR2kRzkX9euGNtuocW4bni/pCN7NUfpYeRcYBRGl6PjjVNkV6kRMMHMKrA7javp3uxgvcmjl
i93bk82KeuvZSJUuUBp4zDsA6KXCSHEsfKwsK9AvM6O3qIGOMnRY6ieANh/PBt8QhM/3abYgrnPK
zUJhU5LC0PJ9Q1J2OWRLcpVJWxL9UjW9S1ceixNaXHaUtzpHWAguK+SHncg2ZwcKGa3Qy1osZikW
EBILiX6RFTzLnqAqq5lu6vVqBuHDKQgogmENNRr5pemwrPKMeAfbDlghBgGJRt+KNVfYjPwaruOi
O48LDtnQs92+L34KSqoMSwXROIk86am5P5RCwmdi821FRdulqXM+z2A83kk0KG3sFTvHtO5BCmXu
WppaaRAudLCRrfx//X+rHEDocokqT2Brjh9Y1J7ITxbOQGPCleAUoMU0BU+OySNmYLamyNgbzz7z
azguXZCJNOLHhM4ORLyiAfzBaBu6Hn3E/IGzZ4i5qRZ8AtgqIXjUinJY05/NnxZ5mcuACH8Jt7sj
xlqxvCrJMmQUMSjudOvw/W3pwKWutmotXevk7kOLAzKCekbllOQXHCcEEi0WBTeHIyyGPmcYA6Yl
RryrJwIMXVlv7Y76ltGf49+lx5TjUiBbOR3+Uvg0hUhExECDMzQI2WdbYtfqGIfBk/AlRsgViPfI
W+irZ1yWlYhkTK8IIv2bAZ0xcoNB2QGNbYqQlf634IzzX2v/Hy3K/3Tuufh66zTc3HzZMrTGCVn2
d5vRIqqRCLom9+jEtrT2u3VXok+4wcaTYhky++qaHuhakKMnt1KxHuEaOF5TXsxOfPd7Gf5M3GAE
TPEW3JvOpJX8yi13PRdtU60GFz13uLS8rY0vkIJ1JUyXE28vhR+IWxzkVaQ9jHGA7Bs0Av+URv/s
zUKa+rrmf3n2Md4vhq/0OK8IhEjF56mYBo3Ev/ABDSQPyW2j8SOQ8woQ0QGlfWs7qVbsYAcVE8kg
QqOEk+R3wVX3LlyU5ntXCluhUx+ADEnHAW6+Yj0Bv/EVaK/5iJVqXRhY8eA+BEN0ZKeoh34xXGM/
YbA9HCmad8zu/U4KLllLTr+nUU902F/FAzWeuEcIYLDPQ31Bn0w/PFf1I4UqOX446XZsp6vAanA8
MRrhBzmVuXPJZ8a0wVMy/NSexSw663+8O4S1vcxXh+/MRepNCQw3d7ioAdVpWKq0U/9jVWxtagWs
d+6+L9BDWTzENl2dxL6dUUlMIP06fFYsiyXhkHtDtoUch6TJL5A2qnuL+QewHnKU9rqgW32uzTZV
1MKBJ9ufWBNMIw7jhMsjtQRLFUVnpdyhxEhG0UDh2PRxDDc29PzXyP/RbOK9UTBgQVjAcPlXQw9Y
mzTdVPqPw3o4SwhqkOR8jpxysZ0nN4DeVNmoDfbq52IdLf4DZW9A3mL5uvToI2FnXRHe3oi6cS6Z
UFKvM3draVTiObchsGk0C277Q+KE/mI+wfl4Gp8nwGaKROogihm0ZcF7EXGYCq4BH2Mwt3tsJMxb
x/nMteEs2InLiggrVgE47kcmJleCdo1CfpF1qCkIPH3mtzVeuI1oNoDM91xWx50woZDC7n+xuTHz
TtKrY6p6Q2Pc46NNg9Z+d2tHwCZFI8ZMsRUFrQ9mtUMudk535JCiblyrkjQn0DLD0EMx7fGExBNn
dRiaUyUd6s0rGauvMMmCZ18hUHEHffRch8lxFBDTyrAmwD7vZWOxqE2THmwkgX8/2CZuJPH+eGVo
FedrWE5R5i0AeSw8SFPIkNFmKJRzIQmwtMtdI17zy1MsDXp8277CvCFStUjmQIHPQBjgdz3giWkl
o6xSVLkJJrd4oDUpeXWjGzwBjcQb2korr+Zp4kW6TZjqFNcs1DfAZ4AkOmnhEumcw3SDyQz/mTeA
tGSBhScy19XdaYjw0Jmmq7Ckqdv/y8XhpmepWEHrxiuawgdJpgOSJJE2unDH8q6Ns8zyR2tKzEzt
7IyQWnAcZN1tsZvuoCsvqFf87C0Mj560vIz8p/AOSEOGTf7KRGRfyJd8zv7LMjikF3QHejWheIVl
jzPDD+D8m/Mhvr+9a/w0QlRhJn8jkn+oJ9t1auNnX3wJmDsUMomdHdI5fv3TxE1ulaeLHV6p1Wzo
W91RjoqrJNBrnf1MURIZiFuvYubDVEJDN4lLcyaMvsj2uwbrETdF4tgQvSd5UGlVcEHHi2WHtb5v
yRu2jjSaU+2k8d9tEPN/RFyLHoXrRiQr9cVkhAIpeMM+TBhxJSF5gtUVjQBfkyhcFRoK4H+PdY4R
K6fSxjBPM+IFt3tTjFUtyDj6j7K9F6AcCGGxCo031rF2yj5nojYvsWga/bM+0mL9fYGQM+lkZLvM
ZQDDGJMbDKmeyCtO7LUSC4wI7jxXVsrK7wfcITV+EPo1Pc4ybKsy17YRejNlXriB/XPresWrCdZG
S9SpM4Qnu5ucaeIkkxe/adOV/pcjK1BlLc94r4Mb1rNQHU1q6PM0ncUU/dHKvyPXUBCSWC8xNnZy
aMCFDEs+Y059zHJ26T95s99XlT5hNI5SH+ZRA/iBdr76pwwAhWD475xCU/gppx5N1g5uIz6EEnE2
ijMaYGUC6TWAhTWoNok3jjU8pFIKC7KymCsDIJXMvRyFP/LjsRTHh9hZ3/DTyGymdk7Qve5S2Bgm
ywqPT/FzhFrwGSEPHcExNT7EeJB+j+ITcBwMY4/8bte9lVHBIKJjTcca5LdLqCqNIkL6JXR5l/wj
N7WxEVRW+twqr1BinXv+zKXjL4XQgoGKFrxnCkF2T/C2MmveOhYnMRXpJTtZpmbpmOWmaZGms5z1
BOPF7v8T0UCRKKB9KIlUZIPIgJTkMCLmaBusYEy+kYhWkAcGed3qEVsT77xS8plU4KBonXFYajUM
DNf/s0TgQcReW75LABou9PmgKKa0VU0PFqfbEXnK42nkPFdUN/5vKGHIpoobyRngDlGFNR4faRFm
0SpChyzHcSKYT5RpEwfqiOremIx/txtSZNtDw8raKn0RxasbdrGZtRDTlowvyvDZHkuzrKzTo1LE
wKTcDtKqDNIhGpaWbnLyzEelUCxUh2O/hXwKDep1yHJ7Jj3WRG8vGLHf3P13R3bvaBbOy67hjYmE
lhOc3dunJI/T3Xykg02N1SoPC7748z5gpP5Zeph05YeSGhxvcyVrG29PKkza4oi0UT9bmRNo3CGE
Ub0w2i6+l3EJjMEyZ0AEL6XM/yod4JrmsCaHlqjCnc/ooEQW0IFKHhrTmExxGJWLUNiYLdqlc2GD
DxH9hB/Mc5a2lG9MNvLkjIzNku1SKBXOjSDqWmIuOZl+0D34EfHOhZ3dgdlryopxGvFCz7pvAMUX
wOELIE438UYCODLlrMbTEzMU6xUp/lNulIwh5WqQ+g1W1GKxHAjZ/lf6qEFKWHT2q7Z4+iQ3d8XN
DdFzmfMTxseqmxf4a3olPSOnJ0gaGwmc5M4A56vsZDLbWLpTyqYTG14X4nboAqZTOPvblitxmOAW
48tmVCCyi7qb7wgCRmkp8onUQBINoALjYmWNxXMBaSOPg0j94OuR2a8R1jVD6fyNQdBaF9mO8YRv
EB5HIOs2yJkL1EVPukB8CKw+7+IAX5ceEB3eiooCfteY8HNiHJpRfJ87/ofwf4vnavRUI6XldeDo
aJekfstWb8EpKyuBwxl/jDI5nnz81/nlyobHX6UurkOo2/fzV/hMfInXspaf1hg+SIQUR5AftLVX
E15VbaO3TeGzYi1Ypl7WuilyeYM7NSkR8ag6f58/pGw4pb9UvUf5Zh6P2zCj/Ro3i8jYTc/HmEYu
pvWPuqbqnTspNFzdp2SIEiSyN2Y/hIfmXREv1nEqHFtmmLcIDqrAwc/6S0pCUHgRHUZiNPu1vF5k
t+aZJzLCRSuAC9qmgOfG15dD6a2h6mG4AlxKwaXZS4OqFCWJ7c4IRv3pgR2IsY3juQyZGq7R/o8a
iDs3h3WTJcrYthLrgymOgX08WzxY/jCDH1Uhm0yMFBGtDpedNtRQLFvQd4F82+h2wT2dR0I0h8By
Y+K54uflJRtjtW3oQw4EcOZqf9Iynqqjx5Utm/u0+3t1KT/UYnvYEzLizniX8pg5UqLEgDdlsSNd
uSkz4bfgOnAzITLQLsUtg3V9W390PfYuISpep+PjDbqXOmKqXWAgFjU1DyEbeWXczWLHr2XJHTKS
L2oJZxANcE88sLPlSgYsNGqlyXrC0AuN9KGttGvk0pBy48F9tr5dXrh7LBnFTy4htK6UC/1KPh3i
qJA61YtVbXLyEpm070VHVJwVClzf6OOFMUPwu3xYLGgbbBxC2f7H4p3qwOzwb0XleoXHiWHbHhVr
A7xiIhH54zdyElQhqLZVGVuHGMjlb6gaQ/YWcpNW6AuI3Ab77UiV3H5XvAe6sqgEDoyLFRp9tWWT
XicL/hV2wNSwCkwfiO+zAxKejsQ4KBo28TU3C9NZC7I3H2lkAZ7Exnh+kp/sHFkve9pBO1A5oIg9
RzVMmTyRvpOq3eSjTUKgLH1c+LA22EEp3XyOWVWyMC1qwmNgp8SP4zYuZe7URUaEHH+w8CTVPQYz
dltzNG1IiMQACJFcB7B7Abzfn6t10VOmQwdOHp7UZYKPr4UrWAjpADVl9/i2DpWPSyz2syqgPvwB
uHbP3PrHKRVMt3ZfOy5Xq2/HccOwsmrbAKITy0UhPlnVpewKI1FrBW4yXiZkJ5pcU0rdEOv775Lj
fiy46RSg4UQzDcNb4ox0Alj7zELv/pSXVNXOwx540pH4zZQ1nylzmXPDEOf17ebHo4ZI9I9gnCjf
KfWO2ZgG8r2aNiO+eRxPyu+O98levkCkys8jLwqBVorQONQ7hItFYG0JcYS/2g/279V7qYH1X3ET
Ba+0AHSzxMXCublHUzPI72+VtvHGLjJ7UMKYW1OPoF8h5VZ/dleScE7u181+KTgahtTatRXnX5ac
FMRJT1+xYJ2Z4qRONEQzdafFawS8mq21LjFDEezv/J5vm67ZP3Ve7p4vc1244e/BLCeYdJZ+FSUY
9bktnPbVsWrKYlATGhYWFWV03BIm24O0u7UiMILusJmlqIGgvVQQcnJotxMxjDwOfZjlNUPz4hXI
L3HJD9m3U1kCtuFcI0hpxNC1uMrYeW7yeJdjaOkHOSfxO28+x7x45QFTpWmXaRzc0/qEbhZpIZ94
hJHVbZJu9/jB0zMItgHSodKGvKMNAebVaIfeQPZcdTLFvrR0TD0axc8PVZFiDZKGt3k5X4yKYoBd
idTyrCeCMNwyMcYqTGkJFuCTnNhmQx0Nvt3NxyauhMzPhyAnF0FEqOZZ1rSzwPDbwm7trnUkpTde
STS/k0i/ii9HMLIBZ48pMPvs0ksCCJ019CNmS/lYeMVXPiufhEpUojQpPytwdzrXJXIsA4VpjYRc
Dy2ENKL7GvbpeivuQuLtuqt7N25N0ZU7YF5Thqbj84OYAUuH6aWJFD0kxzlvS27q1cErrx2Twehd
A9XXXhvC8Iy6zrSllt1EiwZ/xXK6CL2is2jJXiCQiE/qfSKwBzEbn+ivQ9NX8GSXL1JQlL51Xo0M
jrJwuS+TujeVB0o3LQydRqCgLAhGU/zGTrlyUvX7XX7duA/89fDTrcMOvrVb/vdcVLU+r8QH0ZbB
r2oIWcUhNAUJlAdGFOhn7uPsssI9ImLTw6ilHmtLbjUJE+n8n68pK18CQYYJDw8K9aeLi8w/MSeV
v4Hv3w4jnbCCkfIOSUNTIRkQ2uhPhOVEFUOcG+9Q2z9Ai2jmnQ6z9vjuvu0/zMx8yIcLaLJ+zqJc
emxc7H+1av7Wi5orqqdhNX2a+zuOSUvMhehHpHRE+WYNDfAKxQ5xr4/6f9+fPfGefKM/zK19+RFF
doxJphM4b7bhpRCNbzUHm8/3IXk0eX6W7XYsDKdD0+c=
`protect end_protected
