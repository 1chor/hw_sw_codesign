-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
uk1DFx8FC7mDCJ4szhyYUuuMocuF+JWuGAOVCto208lajf57cegZJXLKPFvUt0zc
nI8+rpgQ77GywxwZJ4pi6SxzbYwi2hvXgO8G6LtyeAw7RDncncxS8E2z7hEe/Yaj
SynKn4+3LQvoWdypTQAObw7hEwXbAR9ZCRsURYbgOa0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 14336)
`protect data_block
HViqR5M9K/bHEYOfjcTnPDh+0IZa2jCkF4cUcU1fNfz9PvN06ZOQvC0ilccV7zUJ
F5sKxYr9KCYU+bKHBXlpPzokl4xALoI83cKDDoPOI9a2pKNVD4vGLxMkXhLR7VCJ
dQT6nidTxXaVHMKws/gPChiau3UUS1X+hkaFlUJlVALqFmgohxY43f9ETcMtzin3
JuOZxnOUOD6Fye7PURTnumlkno/IS94xztKgDtCPutnNY1IIRRMRneGCw5KNrr+d
p0TOaIPoySgBAgI22tvJjozr8Ommoa+h7+R3JLJlIkdFE/fMPinHw8Z2siurZhD1
2p3ZijPrRH8z5Nk7ZsOw+W5N9ctUJEyAXXJe4uH+VbWX3pPHaZe7W5zuss1rc6en
AhGS3eRobWHLtImu9xL3HUQ2e7nKWqHh38Dxh9hGKjRydy2bWCCSnJiHa2SlOSrY
Zwv+rL3ybX3JEaRM94GRSFoUr8xOLgorwqTGdyNqthbMLLk893ILK1/OcomPuHOi
1QRsgaWZfn7ZpIWwRtG4HJaxIThBB7UK7IEUPYsd7goiA2Cv8PJaOsqoCjSRVYWf
h9G2c3LqrFe0WbSodJkj02gapwIrwkcBeQ1p91oseSg7ginRqFYeZGxtliRF/IOW
Xe80DZtrAR/FYPKAWxskJp28W6B9cVtQwg/j+tyQ29vR+SOpUnIw8JhSAXWPDNUD
UXqm/sBwRBxv2OzaF2+5Yv7ZsV8+zA51TcVbCwW2hTEJe3LWikyTqiDhq6E8Tb8Q
bsBd7NjsM/ET2CupewNJpiOcwW3KWtS5o3wSaOz1I3qOLk3bH49vRQfx/BfnjSsi
Fk4Xmd/Gs+Xpb/iVgD1z/qUBKoEXIi+hQOMUN14FndoWvojvdgO3ryu9JW3oY8XU
E/2WISNBM74wgjm4E6taWm188nzA6gg5EmwJYGYMykGaxPlOj2PMc3TDfyAfWeWL
Yp0NOU5U4ze0UR/RVcGqkH+Vbt8Y9Q+6p/JPqrUbEu4Uy9RPrK8dxqyT+oj8EhM0
HOGXgx0bfJhVyhEdbGsY4qSbZep0/zp/2+oRr3PgC2b3vUEUlerFC3o8jhGT8y0Z
o65iZD20kVIF49q+VlPUJHTHv8Gy5/kU5vfaPmQGd13SwtC3yKsVyRAAwG1LMbea
A8awNlVwJC6twq5IPVfzVlmJFWIESGtNLAj383XNekQB7QIkZK9zRpHLM2tHmbs3
P3h3u2FhdBRn4mkeLNs0UyVpF5BGWgqBKYdZ9e+MFt5sy+rsTRz92ajlTOO60SuF
2bhe5H4E3I4IiHTR+yAzQ/LhDIPapl4VqWLqVdJZa/Qj+eDsWrPm3ZuX3MY2ecui
u1qA7nIUgfaulwXmrAVt4oLKekFE/bziMPSbBeRHMjI7xmmk7yCdWW8oVTSZE7H6
Q2x4gZ3ATROjenjR4vqM8S5l5JvBr5fRjy1lPtZbDlW9+b3FuncEBRxXP1xJrmyl
es9dzZDfemq3YXXGdbNwZiCG5JHnnBzy9pQrZvAR7QVZX831G6/LnHb+qlyZmgCC
0tI27qHicHh0gi5yWFe+vn9yE8V5MgIwlS69+vUQlNROP4bnJceAPOG5V/nC+IZl
9DSdepL8+SGBOYgCK0Exbz+HtbcwFKlkp3S2drQckaqYhM0i9ceWpd40PK8jSVfo
oG8dnLHMUWqlxQ55HYgm+RqIXTfYZnpGvU3ByrcU+xSD4wHFTFOLdXlA02gGGQ5D
5nTO9BJYCOGu2f/ueCAy4kvwDp0wAJHlF2nK7FkwO+18k6J38g9cP9EdR+2T6Lkj
CPQIFdMpD3q2ASlIzl8uhVFJhd9dDbfj1IUG8v+QJNtrCG9gwf/KvwE0ll9O2Dtt
8tBmtx+2nvtfQyT578rSXjtpywBXw3FokMV0aGprfk9Od3JNcz8iKxlqU8ajU4sf
JDZjTXH90KiUw+AUIqRekvg0C+dLvzyblpWr+oqoHSk7d3Xd8LrdCnnFUwXcGo/6
a4VfznTPsAoQ22rjXQHftM67/HZl+VjVCUzzuh9EMnYfgoEK1sBRxvDGJf8t6F2+
QRjVNOcNoMdkdqTAFnbMsODp8HQRGcJNZuXHYiRaOjwuvTdNIcRKtzXS3OcvLC7q
8Lel10GCtPzIlk2S4ibfilkiBnuaYRjieZxVVtnXGwy4Z1AN8T4A87EulUtoU2rc
j97ZWp3o6pb3GTZKjiUhyN/zV8TcZQ0Og/80OfVStsv02PL2RFYt6NBlgw0CqthC
X2hJZ6l1APPE8d8O1NJpRCmbad2wlvfsQfB+QEPMx/cB+I/BtyrPBmdFS3Xi1iu9
lJu/vyp4aYyw44xJvsK++oyYIbmD7/p33fiDX9VflqfmYroTxrjkG3B+amUOSCvI
ld9Vg7I/Uy9nhBi35V97Sd3r9xUq+HJUJ9fLtxXNVDhsStc2lgU4thJIq4urL3Oq
XmrH0WFFscHX8DhUlK6UYok1e1jy/WwryQvwwG/YDXLZWzkIwuEW5mQRw55enGwt
2neuwIu8VfpdiT9wAv+8ok7rp4Kfm/fQNiasDXGf3mG78QC1Z683xQUYofjEafk2
gyUMe39O8/cTzGUtK9rEMhY1L/ykhBmZO5Tv2Rugg4W99HUGSAsEq/SkgAseWU73
BkE3V+jKy4eM3qUI7+eZbZoPTPoKiN+RZrfd9ORMDcZsVs2mxCels9j7hoNwaMaY
ATjEuSk3F9HFjkO0awZ6qbO0keJij0DyIshSbR8uhhzuo2stBLPx3tHTYMPwviDh
ZzIXtYjxeW6bPugr87zsR4Cw0SLVqO/8tlYt7DD7XG69niTxHU0c7Qo1Uoq0miZu
u8VoyUKj2sVfxgU5lOHv3KIcxSK1rI/kAb0NfQFC85JOIw3rbPZtfnTpSSeXPvyW
frgcQjRhgvdvFegJENfeGuMgPmxSQxQb+Qbnx8deAWj0kIRlaqr/ZqxLrSeQKJ5D
/XBiz+heNI1nUrul24sEIADpxlJ+ZKEwx3SmdF0tIKH307U3xBEYDNboPsFpClqq
sL30/BisWOBcvb4jzH0NE1Z59rhFw/qlSoUUqd7BBje0cwv7yTnjusLCOJszXmpP
nQju+JNlok1NnzLuJDdZa3hb+mJ0GUUymtDrKPSnRsL9wACmpJS419BkVCs94qlv
i4lhPR997gzsUYZQqv3EvjQHDmKZPHahXIZWT0JI6bVsD0AhLubyE/yhpHoh2S7/
bTeuk5kZ2HpqpOPhL1RzjMM5iVXq99iw53UManOP68PT6rROkLGNp6Fa2pcIMhwB
5GdgSnAPiBI/Ho1bD7NhVs5Xht5nSugudShqkzb6xl2cXPKYIxSx5qL3u51EgvWh
tYNFjVAryjgeqgPFAUKbjkwK6PZCQD6i2j3I31yVnXjAf+6UFYYAPI7HIe85Zqvt
K/lFZJe8j+BydRc/eeUvJDvGgJJ4eVvYmssh4GHKTRSM/CsLruyfFIy+GVM0XuJF
FlK1ljua6SSGpgKQO/Fetfeetdgc1Rq0PRmRMzbMdlCwhS2EBDpI6R2RKSnt2Nfo
MAgb80CCGxEi6TwkKNGXikG2A6ctj2lCKZcnIpihKyi1RJMoqiKM4tXvYBwcLTp1
3d3VBs4QZ8ZOS8k5d1rz8snovlM+zFC566ITVc8+DwE5ghuAL7zGYEwUc8rm3aL7
CpE11s4M5yj7D6ZqLAs+ybKKPrzilm0nrT+XsK2768XIPE6QQJD6ZG8JtW56txNU
JLpq4zIxeKJ3t30wNt5iiBMeRuuctOFSwHYoedLGEWkCeMCwzn/HPIL4+KQ18So1
SoihnMU08ykg+hETbmg+iYWqgAqTiSl6qwVwDAzJ3MDDr2EtkmnIL6ckRPOimydO
LdndBU1TMFJKp50jRqlPdxG66zu+hePI54Ag4FHgrm9+onb3XDxMMtbG7PDXaqtY
1/dxL4aAUedatco40DT2WpIyjftbLUaNj4KhMtAGAHCExO/0tiGMtIcHS1VPohtA
5Rj7F/KSEnx8Cg8607WicQUMKh4OIrJIPPVERSNoMe4fsB5p2tsAO7wHqn4iRQjS
XiawBoqg5bBeBm+TVU9BzVuRUk4K5ytsZ1HF9K5MznreOocBI0oIdrkv4d2v46ks
NkFzWIiMITkILrV/AFa2jJlrDHlIwp1K1IXjT+z669J7EyAAJtpQPP0TJ6RJlAsq
TG38DJ4ets61aKmxmUb03MuOGrUz3xCqhOt/lE5YD+A+eS2Prg8GmurEaVzpVbAs
LY4+UI+ku2NYfdcPRXUoEp0/Mv2yKZ7anSkcr44E3B6ny4a77M/DEPs6JK2MiNDk
gBtWp5jQyBza4Ui9Qx/RHQE7f4rGOjMGvs9lBQe3EHEeD2QOtf/yFIopvvB8Bbah
A2Rk/sqNOv0nIqp3ccW/mVkGnvXjRUEPJRl+5MkzmsBevzU7hrZ6sqIQzcxeQ+yg
fC6uuVCYOdrWQZlNLFwci7OlrRPfGBkKT1Uveryoz0HNM6BdpiDwKhH/Petg2RCS
sfoZgoKyz3pJGWMj7ACEI5pny3xPQYnvPfcj58fkckDininzJn1DShQB7gsqKfup
Lbxky+pqUWuAl5Gvn4/0RX+2ax6dDSAZbKDC9G05mtn6H8qzxxtKy+FdkKrzbR+1
3pxHF94muQIUx/f1WEUkWlE91j7aNYz2qra4sd4Sde4cu4DYVhkHqycKeNy1PkYw
/HuDfY4vx+YFjCZu2vFEbcOGe1uaAv3/Dd+kG0lhsFDEHMM8WRIgD+bngCmwWapc
4vT8SbNWWOSNHMUYKYm0pZnwu4mQLcEpMl6Lw9A2KqSFl517XPgpB0GoG/svhMbp
ON3/+/BC9BtiocwghuYKK+lXy1ZJltcMuJe3tPAHfDZpH4h+u7A3Qy9Geefg32ZW
2uh9NVFPKI9DXbnXsR0ikn+uvQXuwHRBRfbxuHaPiD/jg4G9kVC/eCTQT3fYeDfg
K47A6BkWaeUewjUeJQZxlJ1/yHNH6Ivz4cilNj5wvjc8ECNpVb0YVWfVfFMn3BUT
F8ZeESvxwD2vRhMjaDBUq55dSWzdqVoWGPcOJFtw/1RwS37YlhZtp+np4xLYNn/L
72tHXV90KD3uW989jlpMWoMww/n9ZG6QBSQ2OsoX3uLiHobCPCmfd8cLkvyS1uwN
IAdjo25wRM/t5uDIJ8jIthwYZSbJtOOqc53j67BJ2UKOpWWWX49Q8dlphLcAHSD3
a0SgAU/Mu9sDiP4Ii308Bn9Vjv/TurstA2lPqJDVYCFqcJfiLocfuh6Bsmuef4MN
E466xZpTlZ4Oo595npVsceTFk5XNxkWsZxrX16rYT0+Tn8HWZIo/7vSax0cunC9R
/tFJl2ZsoTwrom4hTfuKJ3UHvOMmoB7OtRF3E6H5qzn+W+5fSL4PItAutulE+DgB
RgM2cl3JMoHh6UUvDI28T5R6/FtAKJnaInHi7vVl+fl392BfJn0g839FqcVF0ndF
geyg2jvP7gXEw4zxgcfSGPT7OnsY1dWfrq1ICmyLMzYnf/B/EuNkU4LDhXdn6Hi7
AgSwA7No+u3KXDLmGntH9HoHZWre3v7uP7n81CEYLUayhAUTtFQyZxhe6wfHf28K
yj304mIcrT9cFvDUU85y0pIxp0JK25egOKJRe4ksjXi3EfcD4nZyzZT2FXrvfgQ3
r9CU7HDoO4ePHfmwJQ1OFhTyehh6U/bFd5xk5FFXXKlj1mw3gZaLw3thrszlId3G
w97N91+fdPOpmj298fUIGaAEOIT3eOP4W6s+GzR/y8zTwif7K2m62vKPUvelpM9k
14ByIysfD1/3rwn4HlWBvchdcDjhAquqcAvVp7TMLUJDxYN/qbDpkhLZqfCQBWFi
qDMNYJrX89/v+8CyMa9VQa8T8wHj8M927ju3Knsx4tZ8/p2Sz0i7d6zBx5asBOxX
kKxg42D5A41nLcgtN6i8QVhYfM7qlpT6L7T7VgFo+J0vV0aAxJB9nj47o/rx4bv6
Gumu2rViKzYY9YwUAPZp07tmxJvkKdXfn0w2gt+cQIMMjSpzSGXLPqF+lolqx2fa
Rga1f9z3UDLlXcSgXEJuWrmwYJotnz+23HdZ/lk5NCS+d/ugMjX4J2lwRfab1GNg
DIKTqO15rbER7ODQ0W0zYJl4weEA0hi+Z4mTdjt768oUafa7eIJvCHA25Jqal4MY
Br95Ky8MptCbz4TvJQetxunM89Aw2So6Y83ooECDSr1yEoFjyY+ANthKMihR92Aa
IrgraX85o2mU7WFbg4uB7Cc9gf2X1fpJVFQURuZQzTxbX2iinUKUg9oIe12o7vTN
CW7AKK0EETOtmkmuHfcRgp5R2X/tLoBz0pkJ9e9/kB6FOIaY0mdTDNOlfeGkfVT+
qJruYghueC1bq+lvah7FF/rd+f9oY4llu5lbKNYZ+dVoyJNFyTjYpZWGlBcmf3+g
SGhB1KXF7fr0gfT57OqPmRUMRoir0CJ5WLqGu9TAGtkVROr602HvenJHioaGgBvg
TgQz3W/csFWnVBqI2sHIR1vC7PyEYWmWGxybI4i4YP6PlL654+KdNR7+klBwIxu3
OyWLW0e8EN649P/9Lv6kPNkD2nmSm9qfhCeakFstqP4elLO/2aK3AvSfR4eWgKpf
LnCQn1ExqcbhdvnMQ4M70SQhfalwwWq/f3NpYUZrOIAqciwYxHVEmEvaVmP8ddDQ
/SwneRWU7UqHD+dmSYfODmSxJWOMHyprNpZ76IMokvSqPWp3Dygrv8hGf9sZEzPf
HRGnhhw626JjpXdHOq1gGhinFlvXFcbV2sOm7GwZol7fkIa/rpS99EiWx7OUKF4S
p3g6ZV9XN5Rn5Op/bePTdyuJ3iPi7WOaHLnzwaDjLdc50sYvtrzjBHEY6v5z+Rpv
pcmjy7fQxfjV5ai84FFC6/YasuylX6SX5SOJWm4uyS47FzB2MmYPe18rcxJZoNcu
xSIMHJwM723HCRGk5zSP9Ljx86ClkzLX9OI5QFAWYPgP9hLpR1CXbxNwjeXRNaIZ
NNQDh+fBiiFNt6c1GMhkPHGO+/Y3Jvl4Xi77eqs3KcO/A/Z8tkmyCk4j9vYo4GRw
4QFNE2JP+4uyjqgydDv+KtH4krNygI4uVEt3YlrnPIQqiIh7RPftiQs3ZMid9aTB
6PrzhlQUrkQ1tR0qUz/XdAY9OBtNQBtPvAtXmUC7979xlxMIq7+rlvPUtfx+VFoG
1Vcx7PrECSS06j/RTjugo6pjZbZw2uO++z5FhO57mcLLfyZvePTo8v8N0eE1R4Zr
VMhEq6gmtIyNXaoL4qklgcja1cX4q/PtAdQK+dvaG5f0n+uHdOlvmezusfiVp+hk
QVyrTlgt3ThqqQ3bkb52NoAdw8p+ald3CvDn/VrEJrNHkrRDimaZbT+QcaKBCe78
KvZ9d2cYV/QB+8v1yCkoVyCS+Ml5Sj2+bHvwSTkgFAbD4pp2Z+aUYq1QBm9Nwecv
Eg9YG1Dg1t9N92fZTqQjqCtwBw5yyOqTk8k1RA/JoIzAujj7A+fk++sApEN5rVp7
3uvcraHHRQ4MctHLCrcLXbZrEBa+JEmbfZ7Amt6dXUsxKxBnQQKZzI+viCrzlEb1
4lIVoNGNbIB6S/Y9wwxt7kL8+a5x1C9WMssFSqaWSJCwgP67gJz+i/s8sbu8mhBr
QWgxxutEYPv804UApw12meT3DAFvZGDYCMY8rZsKmQtq+ysxCWwiI905pQmbC8j0
DF+TXJWP5oHAUHW+0OWSNnmoILsTYdXVt67TFNRwJ95M0ucNSvUbfLaMPQH7+XbK
PS+JiwWMRpkrVGDN1Atx9UnVJ3La9zZW36Nu93WkRvDXN4w+TmuxYsGUzSPVhuEm
S6y1ZFbV9TQQIxcLl2Vp6c0pev0mbwqdY3BQ1ZtoUQecdvei0gRAIOOFrnakISFY
a9AKIVXXWXKP7frSKuZ5N+n3gQy0xE998Uri88rvSV9UbhO7lyLIBPcewWjtktXt
DbAXil4feMu+4oK0FpaXzU0XEsTTh4yvQWVc/K4LWFctSJR3CC1IrqY/twX1JgcU
GzqIZKmQOYsumWYF8DCqSXITh6b7M8+SWQPrkhqyq23PPeN2q1prJZR4HVZhZURP
KmQUN6l70Lj2tO+Ziqq/aonq0AjcYG6vjtQk22pSoBRA/QmOC/UsJfoBi4E1qs5l
0115L3PW6HtpVXUSDkli+tyYRHoDIvFTypHjSjDCzjMCJUX4BFKQbrtgCjUdaKEg
TlGBScWP5Utn/rXyd1HCVRJXxVXLGIVCEBaLIra7d5OuKvbEGI0Ce5ORQDxCcdiN
9A8twtHETHMGFOKbthMxikeuXejvx9MXp6qOMm8f202Sq3H+zr5T3ViXhwbqRCbI
RaUA37/KXcR6FDtqfXTqJAZJeJbTrIalFWKSb1o6vY635162jccRS6IcupyiCIIr
DGq0a/uv85/huC3LERevMP14NGMJPeGUSEnudJHbY3zFhyvhiKLmf3f0t0OnBdjh
l92pwOB95c9EPmEYf+xYM2YjSN5euHOR/XRAQYIi0K06rBprcqXiwHl/TwxmLTLo
FEFR0xis+ypYDqSsJ2FexAfE1iWyzaMAboSkgX7j61h20a9AM8dVhGOTU10+9JDM
0idu18If/bFgG/Oa9HvIZhp2hN8UwBWecYAQvEI3idNQ7X0I7GnfvXI0qLIkkLIr
3r8FVRratgvdkfvkeeGb9UR3kuhH8ohnM07Qaiz/0v9jfWdYsyUPVl/7/2YgLNUJ
gL8nvYOAv9u0sDZGr0V506HFBTi9EZD7+JmGkd4fO2WX2jS6Y80OyZy4bBOepm/m
sK5951qiVPig8Q/CnNh76gRHnlN4aUd4FGXQ+rDKsHkNwceAcHYVp8FIjDB8WMzM
r7EW64WXkL8Ufiu1O843UwV2JEUv0YtS3g3aJcpL6q65GkvD5DjNUsOXJViJZ97t
yGsX2WAyjv/nisU3Oj9cDsKs9fJV5ciFXwcna3y3IJLB33+/2clSVJlcYJSJT9zr
cqGVJqQUlbLO4barDfE/ARXkfWGWlUFQW2YJbpFnqykX+8byyEwpYnX1EwzHhIAj
RE08bO1j6qgFZuoV5slf7o4jAs5iOx0d4mKWxsP0vN03ATe5ork3jBawDuP/Kyhc
qBgsn9XdSIi90GQBjFsFkV8r5pib4T2mfKEL0ypJJplgWZUTiMFMMlgp/cpbfA8d
sFoJ55A4t+P55mxyu+GGeLDjx2XBUgZGCrMHklksIgdbHsJsTe8NOuqmimtWSRAo
Qt6KYIoSVeBuW4pkpSAFeC1lDkMjVsUwTH++2nPH7YW+4H5JJrLl8d2J8qu1pPty
F5PQnBaXTiBmlBsYvQYRkaysItPaWKUVeamuPp+E40MF3J4QNjau3lUv9CjeufwS
bFPkxdMwdTp5ZO+cH5t6j1yWXzecEU3MmBDrPeayQ9boCbZjv13h2sEtSZVQsE+1
sbBe9IQF0f0EQRQIrO26nuXYkvhtcp4pTtkhFmRiKR6Ia7QVMIn0fqhRgXq67fEX
xhAHExT7ZIHC/V7e/IghTxN+B41KTNpx5kcmGVhLDeVOOWE/zclaIXDQ6kTCOnU5
If1Th2lEVE24QPz9N+SjXJypWaKJk5cG1cc/LmL1tnoTPMU2mAgcPH7m7BpEvgOV
lGRVd2UtFw5pQTinMgTChaM/J60FTZx8JdeX6yi/GrDIvs+axKQrGvIkipG2By8/
bSRN4tFfyEpeuKDZ3IvvCV0TuiW30XAV9GRX2bU81mOIIj7+evVA1tYzEn12YMJ/
jLGxnQgR9HY2On4+Sn6TmkV7KKg1qM1ReLP0FJAxudFtaq6Mof5V/pr25jymcqo1
xDm2ppWvI8M4KAisNiClvpWYDErZ3Q6zUR9YABhy5uZV56B/rgexvuLUGCx8SCyB
FoE/n/nzg8gGqzK/0iHKLPR3GIXznq+H/ycL8rX0b82g/8rG7MtV2BJ06jNu/9dy
WSIaypDiG+MPuQ0NFfSEwA5T0zfLtLlIVyQYH9PPd+/0aIEQBMORUlUt8Jxrne8z
SFNB52Kwb2jvJ2aZ7D0cCZij4R2qotbb2Rvcvb7OIVUl/iZ4cI2tOwa/yX8AYPCV
7ph1i/btfNXPukki6Ynh0GqNZU1YWCbkpwDH51g7QRokT1/Rwxhy7nnp3Fp/TDYs
DzgrjG1QTIhxpIUgGQlKX25gIrPKw6CWpPpyQoHSUAg+DHRiY11Gskr+Tny+gAOk
S8cRPb6PXwZwAMgf2O0RP3HXpJVTh5+WJ/I0KBv60fpOO9ywvbRYh3Sa+eiXja4C
eVGpUWmGJGeNsX2rma9Sp5CxLOnv7daH6PNp3EGJWDZCb+jG58CYsgagImVHbA9C
JLwvNo+Y0orB0L8Pt/3gcjmLs+WBMViNH2e9u0e+6su+viUzCOVX4GNevZRKZQhw
q7BstOlEIWmD+gdAkQNGrPmuPV1Idwwm3gyuTVsoZvomAczGzhSREmQrmk6se69Y
TPy/5fme7xG58Gmh0zRxdV1h9jaWomPY5GmUQIQm0vXua532XPlJBzf3SuPjxc/q
eXjx3quq0kj8WWU+uku8Pzvj1asR++NBgKyzGXFOIS7f327e2tw7vKid9JLIqMv8
pjbzlIb3qamEjkOpINqAFOsXja9+Yi4wKXGzP1tfFQbzdVTehREsAPpF2BZR5LGX
Y7tHr4puvyE5yyg+v8YarcYe4K9VgtrQWVxPQpFtX5B832cQYmrdu9ButVuoIRxB
6RWHkiPGFyiXNSutu7YO52/qPESOAnOnrAn6S7BwJW0HdFRBN7cZx10bE77dmDta
Yjlia/NFjW+LWHfUnvSJ04q9S2pWtAAVi7tzvH3kQieXWVxPFaXvF9GZEMgGNMBy
7hdpwPJFRz1eFScJoHfsfdPkx2kauoyVQeevOT5tZQxOpM4T2cHKZ3tEwjMiDA6H
VV+0GOKQuDFQgVLLUX+f6ZWOTNuAFSuXg5sDjU2HyYTs5Gg779f2+KeaoWkEeZA5
8FKVH9j8ZoYPbcK6Ce/TiM0i45y1xIJfouDTIkfVQlqSPL5f3hNn6cGzr8zBRqTo
nPrkx6CFb9MsCqSxmVBBJsdB7UDkT+5YdeN2GgOM+yVrpFdMr9zqDrauOZpzkgAU
sM6QP9Y1VTXu5e3y2E4O/hLZ+UF2RR2fihJKX0yW5fx+lclUCsSUC0GYqtptDc5O
tRUFjV/PiPnBhVmmlZoiTEY31QY13/9XrNszHkDinF7IYhuOBf+kWYWNcCvSXqSm
YFn0MM7Xcht3MefxsofG3vKgAysRM4a3vhEdApwkauO3Kr+dEW+QvLnYTii+R+vj
kEJBpJb9WVTSufYHzqWBjzSThrQcejOq4DUXhznNSdOeNLSYIY3wVAYe1AvUgJH0
dkmnCa8w6fGiq77nUJdrvHxmC+fQnK99EsNG0qtjM7LvFkYm8tu+1sPhLkrBmfEG
KgDPsVlDNa9/ABaNl5RbhYIg6Z7ZAJCFF2C7LUEQMPQQcrF2YJjZixUUegn8iwyT
8dDxl8H24Zvt52TnuYiisDQc6US58eS6DH3m7M5yD8SEs1RJrjRZs/xTalmD8Trs
DXBHPuum74Mfnlm+unAjxbBgJiZazYpW/1aBVCQKQUi69IudpcT+MuIHA88ZEeFf
sYj9OjsbdidApye3GgcgniOUwFz/RqeIlwHMzMyxfJmIO7DCDEL+C8hrhFv1fzot
EdeELX5+hjsmBh04FpelMA/b62tH1PJ+4gJXw8W4vhBeROwqgX506DcsV2G13XM4
BWwT+Lx8tVfREr+85X1nf6+/X16144HwdKzul6WKqNFxXmoUsH2eWjSXVIff8D+3
HdN3vBUyZtZ2Gnka3yNCc4wjUeL3E4g7/xhKjPd4v/WcUHFhdRFNsooCSSEccMck
OxrU1Uu0UtLrsVBnIy/EFuQLQ3h/4iJ2OzUd+9mUdmpEke7YHnmMU1HXhxMshs7I
+QoCA1bawifGzZrtKpwXQq4a61D6BlRokN/PLui3coxasQOKxVuDmhI+ZyShtVGF
QXcYzxTsgKjTXxT6GOP2Uphjseve9mn5JlQ1Q0PneK++6NjJVPSGXQ3aW4I7n5ra
qxF4kGoOjG3zrTlnRTddY1xs9spT8BG/xmlaMFWsMe3R7s4dTxJMhHkJdSaBAGpp
yzxNQzez+jmbX3Zsd4rwUx8c0mGzNS77dBnx+m9+PoDN75O0H0a/op7/x9t7WI1h
ItSVS1mzabyqzbaFX+4EDIHaVVSGjEI3lf3sRtUGkZa7b+LZisPPabxH5w5A4L0s
XdkOk3zjEyxEJLFzsecg6L6+aHCSTfC7yzAQDswWWDkkdNM0XRBqZopFVmezDKxj
7tp2OgTlz3Lvm6aaoQNL4ZC2iuEmjVu3j20N1erPD2wOnEjr240rV7FXKT5clnth
RJLkO/VKEM/DCI/k8NChljsJ6edDF1SFElcyQPP3gCQIL7D4ddgMP91zg+bU0cmY
3clqXDXtM2WTFNo8Zih7lhXCveCF8Hr1lrCFq1K7Fm/YjOY6LfFjZmqMPETFRv5O
U66oodASznIt2D/1JInlydnUGuSqidyihCx83WF4/lQehWTAwZ8DhnvFpTRs/3FA
lbvRzVmj5n9L61r5P2p7Jw3hLUIcr7TGNVoGgeD6wbQ0ZmfZfeOMjuSD4aZoFcc9
poQ9FKTIdlVGdfY23kC2n2ZuEKpj3f44vuwFo/KkMxynYXfYadsE6U2yvULBFjON
pWP28nYsJxPO5FconFu2AjQ8XywlUxBkOVOjToDyJkL0DgNApZO3aMY1jmsgcdWt
u3SyyWWZ2HR3ieU89RgVhp8j9fR5zw5tDd2TsWfSKx2tn0bQFSTqEkw5ttG0A7qq
cMqkAK0GBWyJVOmtyHastkeqCfwi4MvZ5B88lYDu7nf6RA4GVHzwWoEINn6Gurkz
eTYxwA7rzfby+JcSqq2zIfFzDUzl6d/u6d7wJkWpUOQFKiJb/w/HrbkS7Ng5Yg1v
nrc5jMhpLoJRobgPDDJQX9GMPunR7mFdmz5Im5qJkOyEKgGC9WCUaN1B0aQLbYe7
itLU2rT/vGplomnU2j0LptIytaTOgd6gfjC48Bovia+kj4YkEEm2z6tSq1MVt9xp
NLLXCT1+jxQ7kuN+7s+8/RNsUZ8K8QNt7gnevavHPr3ugpo00J/Hehf94iXBLPGV
Kqdr6o4804OVfRcHFw1kYjWvIKzoqnY9fXdWePv2QQoYWYsn/MQ0fR2dSqBtzS7H
TkS3RJpD/8OOQPln6UPv/lLEjbNnXz5pyq8dBeIcy6Fa8ly6G8cAY9LYQnzk1Q9b
y8OxXd+DlcjmvT0PfdFOk3g3mu9374z8I5zQQE+7dRYFWipsb6FRRC5baQlrXGH3
+t58+qM1W0Hf+cHLTpCUehsGpI/7raB2lp2aLNpYVYVj+zHLNvbay0194GIAW22s
TyH6UxoKKPiLZj7hbaQylv2gv84kQEq0sahsCWOvDrRp4+M7/FvZ51+Z03vKCKIz
BwZ7tcjxcLRik8IMSx6QNmDoo3Fueip2uI84geaVDdIajuGVJd1OkEahndChlPZT
Zn4rlJkrN236vajc6Md6ZQKyg37F0gvlMUvwNTT8Duns9G0Cy0xQlnRz9HLRv+y6
5PzOrFDF8dcwCJekQmAYJKN4B5JyabQhsFHbdC9RUapGlIMb6Xk+9tjK9BxDle3T
d8hOkMwrSd8v7V5a7D5QbMV5FYblMhqdCi7dEuqvrK9m1PuJwPZPLkBL8U8wtN1X
/pNjhPr3C8SJJ/rYeknL8R+MT58/xlEVqBEwJGt3qlcRz5q+YcGtEk+AJo9J5V5p
IYk8aJO9IR8b8CpbJU/W/BXPOiPeQH34ILABWHQfe6ep+HvyXYJiikgD59TqBGFc
Nzo+WnzB4qtAT3mMLvxSeMfYD9wYhTmgR4axZ3iWuMzwLxf0w9oB8NzVz2AGfz5e
ysKaiaVUXci/VWG6T00N2Wb3lp24VeHZabc5K+2YIODRL+tFMb50louHPV6/gFPY
beJdax5HjG8M4+49fpr7t5rObfnXvUq7IknZt8oezkr7iIbOwgjnuwsgrlavegfl
DXO4jE+F7OgE+36xtGI3McF5SnMD2kAjHbu7FfgsD/hqxNqQikdXYt8k1R+sz49+
5UYAEGiNgn/qZavkSHhIRIh4vJ7VoQvjvP8pDky6kHtYt/2FRh5QlXofiDfh9BWz
rzaRGel3Bp6UIJxJjzd6dNtzEEdIZBLzUXdwgYu3MRXM1MvAL14Uk0RJPXU8O3n1
ytNPILCZb/5JzemRq+RW2rvlhikiClW8/IdFe8J0By2CTDeartReSBmAmRcwbOZF
6eqqFG818cKQRhVUEEb80uyuj6pEFgq5A+xcE2Z3AVJ5NP+YbAn0y1sc2XBUNj1S
NfW48LJ8hmuBEYMgjSa+gmY147zy0GJNpfXWb1vKvHONheHQ04gReu44VukXPxmh
M85enpW/3TaN0fpLY8YnGS8lIv7Wps9b68GaZqeqMYNI0ifGjUu08TF1uNww5mn2
ZROJXfwFlXHNfeBebcm+OQEFl/EZWjg4piuVV3/WgJ4DR9citz3gqogbyb2wMFJ2
hfZ8CkO9vg4T0bCM8b/wCwjSD7wnVzl4i5BtpWRxXx5AcujfHd2X0wMAcd1qhMN/
kfVTFipEcc9Oq7Xt2lwjE4N+AXJTN0BsFazFQ4SN6QW38cLv6WAF0/zz3TPKXMdB
OkIniZOThlRcawJDXRP2Xp9Uju1QLNtqaWtoN4vkig5mAkTtfyIo/nZFmoFIjqf9
br5apqev7P/057KpUsOH8OT3sILFbFg3HKjR6PvNXmBxWubjw1ILHJIDvJwiaaKR
mHKoumkuvs3AGDv0mvkUucQpPjKcDkQ3dpdaclJWvS2anS/ShrdT9hmoxlgNf4nu
TBvifoaBD/au8fsgKyZPAxWmPXPkZwAG8vF/GJ1B3tNSvmr5vX4H9NU+vJvVZ7wS
HxAqIxRHdwSWJ4ToeYnS/C4ERAvQy0coiQfpUBnHGFZ3hkg8AEG5OMbG+z5fK5CC
lhWaMYmE8et2RSG4TQItjan2mNp4UzbCIno959jh/DcXblb5Hit8hdFF5WLH12Zc
g2xsSLZfcVSoPiOaeJ7qs5aI3eLYRwu72CC4Q8p944fpyr3eHv8bV91EJ7qQo7GI
txdMfSNP+GsqHaSUGkXFaBw15wwIPrpRsu9hTagXfUwiyzgJK5dNrDFWGaDS13Ne
CY2WGKl0TD7cosh/Hq4jDJEe8kRxFj+tJjckgamY8BX4nQUsPwiPv1XFykMVWhhs
/ybXW69vhxgJVti0N/NaQi4RCfdZv4dsEZved3Ffs7jkxGGzEAjRh0q0Rw8BNNlu
gIR+M2TbYbKImbp40/hIvTXC/r2WhR2BKRWh8CxSNWyzPZML8tg63fk7wi4A9mKg
Y8xy25A5X0quDBefDutbvAaxVhKJdmE2FhCMn7IjtkHwhNvfKKHzpkihcajPfbo5
ipKz8xSYkcNnfpymGgW8Wi+gTEHTNeWnE/O/lTK+qzH4vcjwByWFNxRTcr7b0osR
pP6YDROxsS4+yPysyFMDmwGvp2J0UOfi3Ltk2Z2szKd32pClOf0z70gjJPUN49hu
quf7Sv5FNfU3cFUq/vweyDoOubA7pLF81LNCWR0UQvTa1QArca+djyYL0Jxx/acA
2Nfmos8s/IK4cricWEKtxvfW1cd8rCRA9opfbgvC8AH83sSAWeEge4tlZfjtcyxP
05kgrf42LjUxv8qlmlEXm++NH+H7i8nbQdsrykw6aaYVNtnFe2utaR8v7T15PsL3
/88+9l+z1yC0DmUJXejgART0w4nGNFg6dZRUA8qEuC0DezJeLeXbWgIhMdSJM0im
xjc+wI7RVZREb8k9he4AQh/Ll6JP4QrAMgjw3WBMgG2i/RFsBm2g9E2IYRPmSKeI
wuci690dWPl+D3vNiDyX7ePZIs3YUOvdJ5YfUthB2swkU09spP+EGWO1I0CuFiWe
MI6Qv7rcHg/utOcNAz4oYc7KYzD7YupkOAaPiMbBhibIbL1AcmY6YXwrblhudHGj
FGLOFITxGhzDGejIp5dDUlIFM4QACCyluh++yX6ngd9NWVhbQKDJs8oVxCAnwbCy
CSJN1KNLyVoJ7Pdp7CUZhhhKY3kriAjGy+Ft/EyjrjTj/EEIaf/p9pMyroTgOC1D
9G3YAB4yxi1DdnERClEzJOgTyvZkB8wV5jiAqfXTSFppzkvykKEt1LH4UTlEDJit
6KKdmZ2JqoLkfhcRnzHB5zv+bU18DnQcELEMtRFwsVcTq6t3rVrSAS9RGPReUaIU
sys+YgtUBOssX6uyvSUu/mxv1NXRlNTc7Xe+HNk0cEeU0D9f5BWx3V7hF68WPdAn
J/pwPRjmG9wQ0s9oeIGAVxDFBC0JAF6ft6RVwcPgVFt1nUmYJYNnR+nrtT9MSIy8
mzHq/nKDZcbeulUzV6L10ri8ypIAf1ScoxEb7p0lmGjf7lIfDLSYDdV6gcNN84K6
e1krOqizKPnPLpBK8e6wYFSvFIUVZEFRVm8kvJRN0rHgFyTuKYt4BA3sZVUKP/Uw
WuxHwWUnhoU0Xg47y9Bn3DRoMuqG/AUc0gg47VeHmWpFsOgS10X8itgA7NbXdYu7
4aByg0ZYG+/wIY4L5596hdTJSi6m+L+iJDuH2hzqvZGeC97HN8/pWzsfGi0792Q2
s7kGUGfpjr4KTxTgLtjeZZfT8ijVhkYF9N/qv/gjskRCtriJDYflK5M9osefpCWo
7lluFZA91LUcLxhse8B/U7ZF5H4K5wsp3XKoc12XIlX6o1y7QOuA6WtwtJesUasw
F/Cn8fCIcZ5SQrn+j5n6xz3SRBRWnQXTSfy9ALVaWRnPnM5lUHgmT2E7Ph3nvDsc
UB2tjG1IXoUL7us0cjkNP2S2FWkx79sjY04FWeoiBFk17CvucsnwHJ1y8pnjRAID
X2EEIO3ZqPx+mku7wb/6PruO6DMo2Xf2MbQMrJQW8OSHKVCzRBuCX2tZVVdKJuvv
4SDNc32hWAiP7sDAbKcSToDMe1DvUglY2mUTugxhZiP3odG+Puez0i9X3k150lxR
nxBTDsdjKLHqr/GDYuxyYuZzn/+gMiUTUHA/bvSeWWeAEO6FfxYDuzWU93JGW+hG
TNA7PMwXjDQ2A2DiDgueVUZyvdprGIwO4lpydq3kqBCWAh6f4ZDKmlU7FrYO8+oQ
xYc2Y+lHbdcOFQiflf/87URs5eO+HkO+w0eXuGp13xb+DEZxTPM2wYC4Y2+Vi1xM
CMKecuSwz/wZIOlshA5J1J5fnCBJVnq7Bfr3J/R0FOO2yP7wAG/fnaAOvM0ZDsYh
Fa4zdBoQz3k4Rhe+bU1JWrRVcmV42bC+sTowhiRRzCKjTqocGjc0+605cWdMQj7G
3jHPu6uilEzyQLlsD7R4rrkZ+DwR9c86AlS0b7ljHsZB32Xov0hVxfP+cd7ulYao
nfHl/pMT/vaSdbVA5a0l/JbTAzHtThZi2NetLq9L4dvHQSwiDXkfQmz0Zj5TMaPv
GeLim4VrlhJ626KYnbzecF13DaVvDDgnVxXCYPqYU/1c20l36f+aI+CHGTqoUd+A
CIHL4oI/D2NPAlMybHXmIxtmPEfGf4MhtEE3pvAf2uJ3SnEpubPGFIW4FqBjvGqV
MNQXJh5JGldcopPY2K2OQK19sz3T+Nlqd0XG62b3JamwByX/FncLOg58auNYI+Bj
BgxEzGoBYq3kqPja+00wC9XX+JNSuSNt28i8R2EGV3wvJCmUahbSZAKQH+jUbpQv
GsSdtG8VNiMjFmbHqPyQvmVnglOU1twOD7YLCjHOv0G/B0p6dkkWe+sCqr38F6Jk
VAUzJ7YXSQkCyaGNVHgvNJj+yYikZJop0Drka6MxY2Q6b2TsBQ6Tvo7mGmhirxlC
/lm/FaS0kQi6NghTX4w2prjSF/5t/p8224yBHh+5h1/jB2r9CXr0/nbA7BbyDgDz
9JDf+mOaIOp3g19foy/PUDWMvx70G3M9kfBgajT75DXs0jJ5sxgfaZ+qln9sR9iv
eC5UvLHCW73fa4UF5nqNeDDoBJuTCD9fhWpHmYLCZKwozI9xtkwS5vQPfZ8IrRCf
1IFe4UrMnnxNlNXXdvjy26c8laJYRMuZKIpTDadlSC7HEhNgnIJSPgmkCpx9wxe5
2yybFbmIl3hHS2itYtUiCM6k/xiXjgHztweOxcqOA45sVNByqB0uuIaNPSa8+8zN
lUjwLPnDxeF+WNGLaoQ4fN1Aq66WrT47mpxwdYYkXR7p8UtHP1dTC2U0tmtbViGV
GXu5gbf/bErgVnHj+YGl1tz+HYC9GcFy+nt4vmtdr4gkMIYG99onmUfxAvOp+GnX
yf+YHs5/HhauUwRbI9w99eyWHRj+95gMsRSO9XBhR3ymhtNkP9+jhZzUXCv0wibM
UWFUUq2abBucOKZsrr1kfEgOBO8g6mBbpmcutf8Plt3SynWInHjPMZIwO8OsBnT9
nNem44vPLrO7dnUrY6g62Xy73oIOwD8sL2e4TF790OmcCP5G4htoU7flmvJt/uHy
K7FTkXklrjvXjVzD4ZLQDA0/JsZ7zn9J0Bbruk4sksmgd7nPG3Q9TPitf8/xZ7Br
fqvGe/6fd+y24cR6xyEg3n6HihxMjTneWTqL1D4OABrPZ+WkdglcLfPkEjkjxb/i
c+DrgCG0mmRW3qk/T3RiTm4YJzD+VFloH0ON1qGJlRoWtnrS+owHdyYCbgLfxUBG
iNx/JoUSe49ey2xez7SxIkRPuS53sBH7Cdsd0Ng8KYB9k/nKidVhnljoM+/2EqzT
l9RCB8TTVgqXsscuKvj0NV452fjC3NOGtwmuim2bUU+BpwJa6fl2RFWHYG/HKQCi
6zV/feZu1bEtYoK6Gu7+fAUU5M+LNKEQUmYyU+j9kTyX/dVnAGdvoE+opFeJP9x9
EDv4cHdq8fiVGCOR0jaY3D1ulHa5IxswuA0NM77noMN9rCiVhpXadXyKvHH/s2bO
v1O1AK0yvpE0G8OKwWxebugFVxC3Pfh9JOxiCs0b6ewU2p/Rs5rR4GmOA5yD2+j9
1JX+fTEEqJELmKzOg5Uag0X3C2xqEV5detJDV6YI5zLSmp93n13UVagDsNX2mTnR
0EA4t/84oWevzXtuRnjcPI4KuyEsaiy/nSNVNaKLXbU=
`protect end_protected
