-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
U9HFfm46M8Gkl7zSeQFOs5nIwBtW/Qhvdu3Cv6RwrupPqIDxwHRaJ/aM/z/DFxd0
Q6D2fDdC+V4AODopyojr1LM5k4vfTNJp+Oo3cboHtXT7z1L8w0DCq84Dmv5a9FeJ
nrwgOZQtdn2ajLRN1HVDagEh3TwOaM30zwfHLwz2hhXuVUBCp/75xg==
--pragma protect end_key_block
--pragma protect digest_block
yo+ilPjqzsx2GG6CbIDkN/yqwJk=
--pragma protect end_digest_block
--pragma protect data_block
b/VFWhYTtpUKr2vPyWUU8L2MivYRUYDvS5FkIyCqnQkT5uQI+Sh7nQkJT7KZdRj7
eTJMGhv6+psfvvJ5xLDs3rR65PBpXx7JIYDe7fl6aRtNdWbDpNXsmzOPJBGz3r0T
ufnH5+aPfimenfhV7/VXoWHYBrIXmhz2qUnErThoU1aw+jfPHdVnGkzyDH2ANh45
OzMhJnm71vKCDACq5qMBTq+l4xHGYSgWQSqW6o688YrC7C9HiOg/CSL8u22FHwRe
KooRJtRb1iKt+c375FPWQYvBVuSPPxlnFivbie6zKTnUITzw1HONAaHMtW1d86Pb
hquCt/VSiu9nch80Pf9J3rMMCIBCaYkAo3q7arSRD5j2/sxXLnNj0MBoy7K4HBLw
5QOB7wCvgDskmJ8nX3m61atUZ6/1qKqtHMVgZ0zzU1orH0lkibZtIustepWNP/Ah
HfCQj7IoE89kqdfTXZZqTmv2no1Vdb+ghTGr1wD3CAHTUzgIXOgGhJ8rmdu4kLao
whdZVGqFhPHdHLbUj841Q8VBtVsKEOXIgjZBVrLyykJFUveGU9RLhoC5k46ybW9V
ZFiyfF758uR3abOPqdPRnC1xY9o2TbsuKwFSjl54mToDpdRnL6QPkr0JAz6sB8H6
hXP/jLJ7D4xz7g8H4kaV6CTSSW00wpiJhCNsx0DxQzfZpEr9ikNndiM/TLD56pBz
cabZ309B1X0m6dG/jUwKHz1k6jitdJCh12U7I/4uE87Gn0ME8ZolruvDdHx9NzW8
EUckPWFObbSnt/ik96WElz+MO1HlVWIk77Vdo40ozl895eCHsDL0XWiluTU4tuoC
SUA5vFsoC5VmaAqJXSO/pwKfBT/P6qCg8k41JkGUdH0CG7rWZ8H5X05rfPXz4WCF
p+QX4U7GZ14N/IzOjnVfIJNfutCUdlW9abK5kFnjn7iNDPwYLkegRxnoYXIq0TFt
jP7YiokPBcCh+CBmOvTzyhJyC2zGDbl6Qp9wD5QY/y7Z+ePLak6IYjBzPAt3yYWH
hBH/uLXJQBYt7MFaRpn221lFhBn5rDxXkFXnLnmxP99goXzXzWnUWbTTqTCIMFw0
f1ob9sWTs300TcvbiApk+9GF8fxgNAlN1lsKt1bihd3hH+cuD+7l7zljuaPSp9T6
40LW3mXbjRK3xnafSa2nH0Dz6ETnfOrp8gBOB/cXZJd5uI/4meYtXqXQlMafsFie
7XbAblh85w8mmOr/yW7RJJRikG4U9ayq1FhQag//D3EzEucZFwdUKhr9echSlFAr
kCuGmfUw/uB+xEMydKW2WmUQwi4PGWHosTDoMkxm6VeS7TV48bF96dKsixwa7a3/
a8uVMD64XfcrUYOVWk7pWksWZIk/STJQvtJufPdt6oad6pmNypqJ2AUAHF6vJUgO
d6X9GDvKao+eq9z3ccHmiZI9uNI+aTukHF2nG25OOfNqNIH1t3PDAx8ziWYUTRR/
zev6F+YIiinqCoHiMe5LKHGEDSBmGTD6VAi5IyN6mOBQ+ksEofrxV5SDFqFPC2rp
Gl5kS8dLzEXRaMwT4WLvFBb3Bzj5DefyiObv9kddcb5mOzFE4Yjjzzmo+1bdMVZ5
AHFd975RqUz2gBfikfvn1gjsz+PY7soIO2p3c3bFvom7Rd7mQAEl9Ya9FutmPUYu
qMHjJ3VcPLZ63+auibUHevX+xvJQcH6lGDfXglKJyll/IvGRv0gKfiQicytmf2tt
JcyIuIfqSA8Rg57AxMngpiACYginObXdcsPhzKfD5hGF0nRMsbxGo6lYikkyK9ii
QO96NeygKU6GzvdMUmw3W3s7DvM6TmtoHA6P9SKzwOOCPTxDcfGK/TtrkV+vURhf
W+YmNQnHqBxQLhlG5WWmxRj5Ybc3SRMcI7DLBR1kOEv6W2oU6m1LPD2J5t5uhuJY
X1/LUqGl2qUuDrTz8ZbklrwpEQS96Ct0pwoLBGZLYnHZ6Aufb2I6moOPQnDgrE2h
ZtBRMi9ODepVKSx0oBd162KOnJX4U5ywt/iwbNtW7ybqcgJHBIEUDJVyYx6uehJY
Yfe/64cwfteVkjTNTNgLj8FldVcxtXpU1QE/NBiqJ0UtwaHLWeuMv8oK16sefKYi
NQfxTelc6WtqA4Bb+7GpJ+d4/NbplW8qSZkrtOrt+kMDl0zCgagTuEA5kBpMVT1t
XGR0R6ZHVsx+Z+zLCV6XWoAyE6WNpuRiukGVCHOh9iy/w6p2xpQc9nsRhXVceGMg
xu3SBl5OoHhn7J/WhEp9lyinHaXBqGHHRGq2ijYlI2ZFBPizZ6pCZQAjKA5tXEWm
NnOEqE+/7gog3NLBMmbqiRC8eZpwze7K8hMlAsO6xwmwvBu6SKcAklrUiEotohUR
BrBc6Iyk+xj02yyJ+MOT7EH2AvuTdS+BN2CDeXjcynFfZsf1dA3arnNeFf1etKuR
kr3D89zL1jnwiPO+8bebUvtK3zrF+VKHW3VUMvIwdEq/p5AZCXGlJFrJ1gOq9rY6
+5hG8ld+PYURt7fc9qa9jmT2zrMZV8R8qN3A7pV45/npRX4hAUmbTug7/QjUrNHV
FswXhYsZe7tzqO7LPQq/idZq8Asfq310FSoI2lYRDz8BVm0IphviHNjhZoeDN0H2
ZnlOPdchEsNmSCN1d0nOS6DWn+SLIKfmgCWqwK10fqMX5m3XUmgDy5CHfSj86UVO
fMwdljjaQPCCkFLGdA6kUvRkUbpiTWXIlu6RjdiZWwoaNNtUbyzNXJ8Y/zKYaynJ
Jr2MDvM9MD1VsEZu8WCrn85cQ5yoxa3H+lyOpV2gaFNra3dTkPnob8NQHrV8OqlZ
G8wkgRWY0c6HdRey6iEI2T68rOI6fdqrqRXcp9BpZsHHHo8GQGPE4ujFq827D+kE
10y6p5ovBQhnQXGRf1GbO5rQ7Liue1D1E3XgOQzcDntoA+e7yJd6dehgmQGH3I45
TM1+V6e0+8Y/DdSmfbKW7z9VlIMqgGzEuDBIWRSEa3Lcv0cTFbfGknjhG4KyNxIq
cNDTBM9LO1J5nWXjh/aXHF0HDha5mIAm2jEG2BarH1DIdhdj8U6Mdaj80ij/2F9y
dzq2eJVCsh4UE0EbI6cvLuE7UH0RMmcyG1kKvysN/P6AgD8MLqvepA0saSWBotpL
kqeUNTrUCxn9+BpVLHvSfc6htgJQKvkg6m5w+W1vZpogs7b8UN29QvXpYxsmt8uw
oG751K2GPzyEaMg1YI5mzmaZaRpfP19t0y3GrMYDah+JjXXHTqWLRY3evbMLNWn4
eE1gweeuVEzZsuhHIApFZUD/9OI2Rw1uvSGWp62sQhrg0RSwSOwKWmgze9p31HOz
kDu2QRN1oAm+p3+7PFSW5bZDf70s4kVe2VAeEz7LveA1uNn5xA6TIbzRHdqp8PH8
MALcWLUQlDeX8s+PELBPqGcVUN1PMEaivszmSgkAWp1zlxVuCn48ieAfs+fAHJV6
PO/2kxMXcQRJG/YhIdIBdgswiR175W5c4ojB9NzQyYS4y668HmhXJhJigjiE/uxP
JR4KMaJQh/JoQlhRPaRAbTQnX2kOj53rKAsvPnjRgXVHZ8L87aRslVtzPuCJwxtw
3FfJf8o0Z/yAO05jN9cP2lLEhbXX+ZaONbsYY6JHTq9/GaMcAY/EIyZOz6ZOYTmG
Whkf8kH9ByH+KUXnqIKoEZArkFSrEjwO0TOsB8ejHOCR4rCEDJ/vnLZHGBazJDAz
oOKvdL9Au8q482VCOy/XnGPpnbJ13/nnk2XxSB/SYx8YX6SgCUQGRqzgpCNUX9Oq
ihMhc/FJ0yT1NPl19U0PhoSTpSx5zUuo5G6XfKalie/yh+7MlWPu822UT5s7pJM3
XeQ9W0mEZwmlesCj3LdvqAn3KHJtTfw4ih5aZRhWeg14tghopdKbVh7AbjPslyGW
OpdQ2nIVR5r9En1yOT/4KuZk9Vuekbq8ewrkMExaOftPkNvtZ42SnC7bRpV2aiLz
4IAWnvqxfkFskj3dz3KHgzr3W8w8TR4+rNaFldbUdXeFpkVtY52/1tm9grZwmTWx
sL7HLKzTviiGcdzmY9PcveuDhTSoP3Q/HQick+9z6eauTlcVDBBWMkmuu6J6czgR
lhyFIZtRcgNq0JpMqOfKkDtiAaWgOYBgqtgX5BAkuf/rGrIAoGrjIkMSDIek2Y0n
xVSQx4/XFLH/8A5cJPQAig==
--pragma protect end_data_block
--pragma protect digest_block
okyv3W0JYOKA2nw6R5xk2vjktCc=
--pragma protect end_digest_block
--pragma protect end_protected
