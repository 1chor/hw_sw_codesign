-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
q99/5YiibixJvke4E0UfX6WZXYi6BgHQGg48w9Dk9l1hCvt07Iqp1ZTyF+xGcXJxZPqFWkvXgt3u
RLAw0e4oTnZp9/XH8WyTmf7HK9yvQwgB9krgJ6LxT+SiSNWJSa5WBV7UtXFvQtwyBN7+Hr50XaX8
HJ2wxrDWf+MiTN3PPC1ZZYFP/leeLo7Ho5rIrmSAUT5lZIzGysLWkt8EO58nXn75AGOWm+tUBECF
WBGSiLjt2utWond/C+GeXKGuAmo5ua7WpN6Ds8bqeNMYApcYHjS/026aB+xuCAb8VLrqjd3B9c23
bXdJfbZ1hnN0lkgDT5huK9svPSTPu/9IJ6PYHw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45984)
`protect data_block
hXFTtO240FWCXgoD78ydnhvkOwezH/vwjC/wDEyuf2giYUwvcltmMnIkfCK1nZvmLRFk7h2RYkJE
gOa3sd1j4aH2T0WZCEYycW05/NhbR+wbVVPA1CBPakLPYZ++CIbGiLAYsLPcw+MjQxaW0GIr2J8Z
tm+QU6M2Upvkyim8SrGjImm2xiqNMUsYkKrHfphdshoZQwlaqY4Fi+Yxb4WZh3xGjOZZmGzTWerh
I1BjY8p/ZxzdOmCF9mK2CYkZM87Dc9WvvPqSgxZVQASq/eHRFk9PRICr2smFOUvCivNOK/K+5qXU
KqDkdzvJCqr97u8KNwW4VOfd/98lz3RXEh4XNQxXdI7oIqiXNCtbkwnAP9Kkh6MNwAdQCYNqPzyw
KXjfyRG5qf+x8oDUi1Dhrq6ysXT6rjXbXxDebvhylawytusqkrVMKs3k2HEBa7UXSiJWseCD7CQV
p2mOurh6gTbE+FERmIRKQUPbYtgbjhpad+pdML4oksgY6/s53QpbX6+sKUj6ddW4OO3BTLmdja8A
DEck/MiSxx62pckjEoGheYePRTD2/i2DujBYgLESDH69rlO0TilJvX6K2jSkIGdLBczeca9wYELv
KjSczCu03vob2tUHQ5KvaixMAHH/qYs7glMX1y7/DbTWtA+otbBm0pYJm9IitZZSyU2FmLxrb6lP
I+EXLXiI2mFRfEfhmuwC7eDUDy0Ij/faDHzSiokJ5PngWl/EYbJ4iS4FFDAXGndGb9PvZI66oEeD
vm1cOoy6NKIdrhwJ7sD6BBgJuwjmV00Um0JcP2QZUFlJw28j+6lOKOq4d3KeiVEcCZrITeAUQFUf
VvM1TyF84eV3URUOFa/WTU3Kt+einn+/FEpykEoKIz+PI5n7RsExQFuH6krjP/1HXe2RY3wgPgJT
s940YfeN9qB4J70vaKX6VSIMMozPN0SHCvFG8/6pyG0cHOaSGgHPOtrD6k9AlpxGuw6EKgoF2ZP4
92Ctp5KvFXz4/X4BlgYgVOf7NiZci0CbQgXLNbDUEXs7Jo0kvJl7Thi4SQOjgdWd+GPWWX7EaPdt
zcidWC2ZCxS4rfeE6MZ7nh0EFUHJLDQ+DG6ciNM+0I1J0+qjD6Qyggu5y7l3/YnePdJ8RrB6asFb
bd/7m3+lv4RM2H/zfyKhx+wnG4QJhu9/gUqFWHJHhLYBpebZr0xVZC5OSnvGaNQciEOdLOKrlaOq
e6SwljteAtztHgS4F6A+PbFGXQYJKiWpNDom54waQzUVo/Hytc7CJfHgKrzFjX+37k3ZV+Uujr0d
egCZ87VP+23f5bWtB631U7k6/eDToyNMSAYIe/iMJBcknMPGkjnC35aW61LfEwql0HGq789XY3pW
4RswiQ5Tv7BWX+QesFL3xkOobkHtvrGW8i1aJ0ubEvABpd6p915ew/cNo9E8QgXenUC5U15muQCE
L+Xe5z0qlZr91JVLekoz6g/BsMnjD+9QG8h0oEja1e69ijPvTygZPVQrbD6mErDUb+LBTAYREkKS
aXKs8sQiNKV6BGNt96BvP+Tf24uFzhrLUcdUHwChBAjHKVfmyWNZz/5PyHxFbUsNi02e1QNHvvEO
tn5fy/72eqGnrvuw29wRNwOybE7LJMlzQigJWFK55UE6Q+rzYHmIg13gmUdEgEXGpW6uzQXzP4PA
rx/rPQm2QWbJLUHz1tAI3ex2lnRzWZAODRo3K4rYSXPmCnyeqHZXA0ERtz/ULiqQIzsQfIZOi/Jq
eGk0z1Z55Ul5/XYDFUGcK//0bcZcaKIOu+1PoUTNBpImJ34R1pMQS4hkmQGRbZtoMzzZQjAlrEWC
XJdY8sNVYwptGkq6XrJi2/RJHGDf1CrPjRmlBq61GFD1Dy5t+4FlaZiFyUlBTOd+VkZaudDqXR3o
wWgTHbtMjN0sNRuhuTrxfF8EWeToDssUVeDlZib7M2M3ORYstnB0UGpl5XHKuCg2Ad7RV63aaRDJ
wL/jzEHpcKIuQI7tjk5wx5ajBWWumHd/REy6cirruSL20OIunSeOIwRryeGvz8ixmIbvAq6IirUX
VYNkkjtaxbXION4YZ4k53vxHL9aj5mViF18ZRKwdCkD968raCPwLEIe+pgJl+wd7nop06Pn6olUi
sWwoXPQBPSQ3mGz24VmdNG8p5mWZpIV7IkUWPFSYWyY1xnwvijbaXImhafrVOAeFYGgsTt1B40xD
WJ1PnzqtiN/SejWJjEGIR3gG94g/PSz6tGcjUk4TZ885kUxlkzMIKrhtu6uwl2LI9u70J+m2I98U
4FACTfGky6DLkOxWjMwGofh6ZKcFh2KOBNkbkXj6F9I5QSjo7bBKJdBfv4TxSYpAK33vwP3HeiYU
AaiI/0ShCSyiHj7DO1qR7XuaNeGnMMDs+h8BqmD/SgQEvKZHwIz8G/zIhWz/e08lfn2oIfyrBdm1
gx3tMXRWef4rOv2IzwekiEoBY/M4A08hjDMV+ggjJ9DiLpMPaz13WfimbI/P2+5sdb5k5Zzp29hI
LCA64BCLPec4aMOmy9xIQM2y8bSESI1VDEFWrlGABLw6A043mS8fBb7yvuHJnQM+76xzMzmaLPgc
mfjiwNKobk56hqxV1jhm/3lK/7jm7QBcBPNY1ZQ9+qzs168zWjKcoNZdEEeF0/jpAcMo0naCyeRl
QKsiEqK2MQm2vJ52WBXoHWS5m6datE6B3O4Y8El09OWX4Ob8VYgTKpJfGxvd2veK8DidSMlxz8nt
27wGcFr7YlUMkLcQiw1pGHMBT8UkmecXeET1e5MY3XIUUYUVbtp8QvRhpPe+p4x0EuYL0H1r4vcM
XgGBb7VazkQ/A3yovJ5gxcTgFQx6poalZQRtSukjOtxgGQbf8I2EyPJJy2nDSkp9vPPHhRYdmWxn
hMGcbrNROQrgTQf7Ub8SYoRb6a9MN3w7Ru0EtvAj42HaOFItG5qcaJw1nKPgoMUtBtdGsu+6WslR
mvqMmUSUUNtvgu1UIo+cKDQTmRWgPBeU7eEQ6VBNvl9WTgLdOJtHcr4oPDfHVCoTjrSPUydYP6Vj
DW1tLQcQo5U79qc67rvc/6TtM/tXboTkWQQ4G6eEb9C7L+YuUdJmOJ9C69GO2NmIPZYFWRdIpOxh
CnPCvP9xDGE8W5sySJxImpbghsFsAARdxV1NmdxtmOKEJYr4rdcqW0Pr+6KZqJqMur+3V2Vn0u5X
FSfwym1tKr3Spk+IDmm0wxo6pVRFGuV3DmipoeWIQVlPW9NG0TJ+S+qFJSVyf80nFPxWgnEZ7eAm
jBVMA1yy1kLptjI/yrcrFkmLnumh74j1SS/lnlr/ef2DWu5AUJNmQT7x8JhyCrrjrBcTcCZAmHOD
vFIKrgR0vVhi18QGNsWRX2TQbx8XXGJVJBI14wHjvyCk/TaO4yJfdheumuJargP7CbmiEPFRPHt5
KuvJhJdjlvMlfkb6upZZLT0FPeAemGSeoo/DkIGNT8mE09e9dpA8QNygGzWhK5WT5RvVkRTvU36h
SPcEZWQxFWKKNe01QbKozebdaJ9EPvCQk0I62H+uO8agMEpno8T6TMqSI71ldzr56SQKNgDUg7r/
Bu1lU5+Y3PxcKxlAM36xUgWEZcqF9hfIQv5FvpMEGheqhvEcWbxqWCOBHMRWdVjhKyG8qkgADHOM
z/9HlucxjBqAX61R6QP1RBph+NR0/cFXKw6ZVjGkXRdIScBa9MULycr4bT/91oSad/tOdh42I/BL
kqTkGx4tyt4/mC7SbdO476sTsnZnVRuCqq1zCIZR/rzDPS1kmOGHHQBbX4BhUevcrQ8YmZjxnDzK
3T3zFfeqLEkrs1b19icYhgy6hyKEg8bSi0YxaD9bGOw7ItG24hDMPtRu1FWEJkg7RqK9KMXSgSoX
DXIeyzFiCrlll8keO+/Ok0I7k3Mx1c0HAvvocEB3XA20VFctlJ+tWI/piAEDEtU64qH5HUSN8BSE
3+424oAzspGSh52szJC75nqYzJLgynmnZVzl+9+HToTlK1yw1It0w++d9GeFoIHu1Oz9BByWhTyj
pi8m5j8DV5mlniCQSKjc+5c9/ujmcTspBwF+aOAo0m4eljR0nSWKDqagUQ4YdI+xOmP+4kR2rXnH
6u+nx12HGVPDVgNhG8II4P9+kMnqkuK7cMIXrF3aDZeT7YFIk2hALZWG9QqCa2IBtyXnm7MNFRff
2ybsUwhqex9DyEKrW6KWN4q0X6BeBZJapvfG/l/8cS7GIWVVEsEzdcU6fN/IoIDRykjbXVUSzyZF
1tWPCJVXFo02om80J7cRI+RZyIXUBOR2m2uZSzlYAwy78k1pcUfXf+46JHIbGmLk3ds9ZgboNM9d
zfamiUEoI+p+p+ABdyjPIGRmmsYPaGFazktYfyhO2bUCxMlBqbKOjs/Dx6hOV5jgQu2WDUPYVh6a
EZWIyvZY8NQ/tuAeqapDljSr27Pwrz9NagbpRTXw2H256+ru0F6JjOr8uv63Cj9m7PR5MzImMcli
ge06+u43tTBK5idp5tSYgt/xYGcM5Sfy+C6TYEccl7cKABMRckfZFAYug4c8mqeGHwrcupOVrKkh
+XZP1QJMHRqM+8GW5tgMgjaOv/kU293Q2RDdbBbjwuypvf/OXzSlBLVN6YofMm4sWr8RBtcoTIY0
wLN5GtmcMxLbXivIVl0A4OYX7gJ0+24SKpj9O71xNcPQudr6xakYrSCe9Yu933zbTvWrHD9RvOsi
ms1UpfzYldN3BuVK6L/W0ofx+YQc+Af7UJaNGMGX8hBPLC0K3qi3RQU6vuNdBhGKCHv+N8JYbsSb
Ibn+m5rg9dW01Qq6LQgW+i2xYAYTbUey1oFf5vZgzL0yANzwkiiW2GXnPni6mzUAoNb77YWBuBMn
uOvSqNX5igdlCDxNywoaFTVoqKHWBhi8nRgVJh/Dh3i96igLNvhn1FELBRrezqIM0I8M/0Ilx5TJ
oWHqiIeZjENnPJ1biQEkz5/FeKySC8652beoDiHSRYXXzVfqqMOzXRN2dldfpOSf2VzFFXFbH+o8
s7Kf3pMs6vsDaRZGi1i10OnVKXhO0Vcjxr1e6wjBNs1MXMAy8UjhKgII5o/WJyDtytNp6fsa/zAi
c7qJjYiXO8D32pSxSWFxEuOWEQTaRqPYusk5GIOrnex1l764U8jlUiMZCwzIBOn2YtV88zecIGJv
8fxpe7Cvk/hJ7o/XSRuAgKhue1vZ6v+W2gGr4y4O5uPlZObPsse3egriYZmMi1f43DbB7SwleikV
Nei4h6f4CnU3xqbaHEjXmufvlLh5du96f33BCSsxWF810OzJYCxDoMjET/Opq2ma+7DB/wOyj69L
bh090FCUQsh/+GZZxbKsr/aprMyYPJ6GMN5gfVlsrpBwE8RlSB/FhCnwTbpg5ijDvlflpUAkpv+w
80QW3VQl0WVaC4aru51u9kvuPaBHu4RLWEwZOxq8T6PhPgYQY3MqTMDcf52HnVWidPIiMrfVVpY/
dDWqR5Z6J82sNsPheIw8cxjzsCi7DEzwLL0NjucTUkEPjGE1ZW4S0SXeW7Y+cf35WXBbdC+LFJH1
xWbBe0R8Ow2KjSJW9Knd1Z86vUVDjgGHkCOOLY945FXSZprv1rVU30uxl+4RWM9d6j3jOUEh5S4z
ZKmeaG1zThkr9gcHbPSQ3MgnUYBFrCRh4J8JFtoHuswoN+Ak1pJwCj5u6mx4CIHsbRFFAVFA7Nc7
ArgxrXUOD0TlHAhotr1QqP2IUttXSwVxwTY1RSpaXn/3rF2EAEwipLDTej2lD32Avzl1YG4kJHly
EQkrRFap9TdavS4oDFy64DVQynlmF01pi+cXEB5olG2jucgL1V/BxCjIBT4g81mXW/YVVBZcop15
UYR9PXSQQHn+2c0kyqAGFapVLqVf41noqc1Wn8p0ms6FqJxyQUaoAWhJIsdKln0uUAdzqetpTr6N
1U0756zOz5D2EJgoQDWliOmO4Zp7HmMwo81OwHMjFcH3EgZK2h1BJnAIhKWuccTMg92vK8uuHNaT
1SUDug/LZWi4kDCowUwWmoeP8g+LV/Y2BzMTqUHgyHnOXLwE/9ZvqkB55Wfnxh/4pRtT9XvbnkJ8
I0agrNm847UG4iHCaFCJs3+PIPucBS3TYPTlNWWPeII42owXI7jdI5E9C3JkfYXA+06SlMz/1Zsv
rWUbTo2daJuGJUviK9b1HkL1T+tmyedWkSC465VXLENm0LgQih013Y8YbcRQdO4pMO0zGIbtSs6X
FadvGdB6yvYgAsxxkSYFB6UfUalnQ3x7H+d5W7y2hXOFMlhxrWdd2PlaOCCkBibjxxxpEvm73y0m
80iB4GI4qjDHzc84zvk7D7vJNhePwRC98o6DY4CvMTXeuupR6XtYij1wjZKMlAInoWmF3LuzfzQS
T6ysS3unQxyf2bW9TxLHyayzmJXVVAHj9nJ9OW2ImDC4S+PCD/mrlN/XBafvL+ha+It2DBy8iJKE
n3N4b5+GTgcW0tr0knroyA0njueRzO/rc5CVOqVDXvNlcMdw8gT0N9fBnFIkwFBg159S+r/1rXE8
St0+/33q983pcTH+tHpzRCwLMmGVr++bqvRuzTeCPw+yN5oNqmuQE7kmf1tSRdDr+e6L5y5XRT5+
0LrOqFVX2RRZxsfvj1OD47j66RPlAk4P3uPx2LArHTpqxBXVkD3aBqC+mUurnzYxGlsZvjRb7qNP
p7yabJtS5saxvxtu71WlJBqZslJiqjLBOV2xPhTnrzhp2EFyBYjP4za/l6He+Wv1ZP+NRPn//ki9
RzwkTxY8SU8vd4pGzffbEW6iudFmrRZEJMlvY8RbesPqkGKC7bo/to3jBdSmuLty2gCM4FIMpzjR
l871lMT5ZEB09NTwbskJmQfxm6pTv4yW8bO97kClVazx+z1xP9aeR3LuTk3c6MVTjp90ESJA/amU
1xsxsEwxBN56njTwlCGnLM7SXwTSUPuVkSrngAYM+QL6RtAZg5TJ6Zr3+FtzRZyWAmrK34WzRQVz
LPiRONVtoh80usDp03ifPID5A1/e2LjW/I6BnAmXadvcGeieIRyA27xyJY9uQDZORGP/yO96pp/c
VulqWce0XZvfeDwZK8CpPR01yVO96jwiSWDHN1n3P8oo5Gt+URa6st0xZmrk2MOai/UlpYtqwgsj
YHxqbCTecT/EcjiuNrSM6rxD5U0M7ShTErVh+0p9B2SYKZhJ0wVwtOYsb6ZVO8gnMfiwgk8h8bbu
4KDnlS+U4IIlHwdniFvpH5vHNYimhYFZbii0g5whH+UIgJKd8GCKoVZyujD4n33TVXdN+X0kbyaI
VTfm3cxAbOJYLyXPEEOx+LFg+Gp5IWdb0TIagycMYtvsC6Vk74/AExX+OyzbvxZBZ82+G7eBPU6y
ePQwhR2M/lxnHhzYdYn5/y4y4NnXr2BRa+PxvTUHlkffwDwI3IoAeaR+DP/c55ufGNGqw/bgIn7W
H5AykH9qFjZeqxz/D/SkRw3NitvfdxnQG4+rC448nFRyZKHUb8RjdPWGwh6gZaO/YhimSshTQOrv
jD/B4vqCR4iENvimykCytH5Sc10b9/O4eTSQhoJkXkyy4+pHe7cRqRhlTHAKf2xU1eFeXRHODi/F
afVSTtd7zcti7XirXzi/9vjy2/fQ7/tx/tWmQPDhBDLqwrQkagAgEaM7VPXEinDfLTHXmSM/r5DQ
vLgywLjZSDgEbCKmTcYzU/wrVkRCr8lUNc7HzEh6A5/Rz4buFvsnDMcWunu/aRh5LlwRUte3hoTO
HviWh89qfQVP0VX+y5F7H4AMdm4QloAXuFrxXX5mrEvFQtQasztl/LUlQ3w3pW86v3QAEvaG6O/X
q5Xaq9RUIO/sYvp4AQqNsfnSTOy2TkJFNxVFL1ee4PLNay/u20AdV19UPcjnryWj93HVyzO0IZdV
keJoZD6OZlMUdVAHKDGgZUqqihqPdG/VjI6Fab2hkrTEqf7pPGYXRqDKIiFQ3wt2mPsCUn9BRQJe
dZ1mBs5aWmKLCc0yRrgECqzQXahh8XHKkAZ5yzYZupdwkggERc72W9iVqbZHuYt4XNtdKUn/e1tf
SmlHxEcYdGZRmv3YnVfQ1+o7ZUfn80TJQOYIxu++GuEiVprRkA4htdMcc0UytPNc8Ztccymy4Wx7
rYs6QuI0BmjdV5gfUnkbRuCW3tin7l1VVFnRgTWyFddsZ7AvoVKW9/Bog0yqp2YO9RNo7cjNgh7v
7rB9YNkKllyWoG/LNDXgbPSU01BPkL5N6DUZEBI0FqdsTOywvL6fF3jiaW968j5oAyH63Bs6O75l
RKwbVENmlkZ0OeTZhCVj2B0mBiNfeqEfsVVIxQsUaPbao41INrL+riP3utJuKVcJupqKLv2Vd7+E
nfu4C04YRWTDBkGD+r9kh/CmPWUaibpNfHTo6N6FC/5LXwgPxzreIgQPGxcmFgZkgRedyXygGZVp
gqJvJHeecKRNMcGqNaKxqh3yOLLOJn1l8y/AAgM7OLoUQDIM7W/f1zggkufSYP3W7C0/0FKwxcB+
4rr1hxKvofej8Xt449xwpZQVBtJL/dl2N7ReBCqFPx7f+kOpEwVRArd0icsMg2wradzs81KzFRVN
snNY7NuIlDmBU5r3tBYSM0QOFVIAh/X/avU1xzHUfD3Mc/7Y4ajRh/OQTbn0QzUCt8/6QSXvdWHB
tJUx6RddceAFcybvVt4BMJKA6MwWiIGFSrMbC+annXwDTFvj2QtWpH8BRWE7uD1raU+jplAY9X7Q
p2eJpGjp3SANBb3to4NFSeqZyDEyILe3+qY9eUkCWA2FgheAzyIlb6DsYuZlb63l/KOp71k27Tz8
FCWngq86FK5mWO3/cKMh55pY9xxeJFE029uBrUtZZzesDBlDz3wY8lhnpGXznyQAu6n5CS5xkzSl
/7N8tH5tpoDFoE0Sve0CBGQ33P7H27GacjUqn5wSMRskL4ifIjLPQTP9EDmCSvNLdgiQUSdKh42i
0eLDbxsNW09t3Ni7LUozv7glaYTNED1Cd7nnZOj4j2J5kmiFON6cUEDffHrOEZyrsUv1UdtZbUvu
CpaIEAvcN2d2qQliEOVGSsfJY9P2tIlywVCEkT/iSJxao+OpKHqrkfsjNKHUazrXZhxgp593gSpx
rI3USHXaqMF2fDfb1oC5NHuPXd5LiDADCJ9ktQG4Jqp82p6iYjaj2AYfbxOvRUzBCBKnVknkoKzx
iOTsDBPZxND2xI0MNAg4UGqPLIWlHxcnu60bpSPdcr8YHGgFaeVeF5m9p7swR9Qq43kwWa/nXWN/
qXTL9t+lufLvbmKWflr4yAEVfDkXM9rqr3291Sp82VzxB1C5QZWzlRf73YiqOXbI0QNG7HACyOtx
NYx+J0Z1PD97ROEmcq3BANqw/G5LiWPI8yVS1zMhYt+VUUS6d/qQnZnuZn+CXdPzlo+iVSbGiSW/
TQnAheOr4h/1fvg/MzLcyWppkDWZAKEV8pLkJAlvpWMvYR7cTHl6VQIojDjjN851gQC+lHT9+cex
1c5V9YZ4nuGQ61enrh50ck8H8agUDHBCIiL9NTaoLm4DMOjGFihvkjScBmtEQiI2Oxrn12BgT9TH
o4TUpuGbtNR02nocOyB+AiXg5sCnsas4twu5gtukE2wlkvoO7wV+DXFIcmI4BhQaZltKT5snXFIv
e5fJR3Oil8mJB3exTbzFtmWKuZOuxj6C0TQ+iTdCrO+zDVm2MGfCAc7DxBAjz1troYs4YYlV6SVa
ONquod0JPLUiZ6KxL+7ywCk+o7uE9kdDPJqFuNGa7Drdh0pLAm5YnGGoaFPZANr3jp5cTCIJv6H9
IIPDU6000K8zWb5ym5/Vcz0Pfm6vpLOhT1SLbnWZGLd9N503wcqaUSy4vQ8ypecNUBHFfhwJDhKA
exA6dsPb1ueAvaW2ArIZg80IdhP/eQb2JHXgnEyHQWKyRYm5iYx1beMsL5Q8U9fup+CnXXjAdllm
xU0uGpuvO09pNEKJd/8AAUeLq5uYpzh/XtyVDX2AYcC40bdqKruZ3OlSCl1JGPCex4q6vSbU6ZnN
6ImiEdLaqmLERGo5jBKFQGIzKAs+4CeBLgeY9bOnitkLKWqUlJJTgw7spt06FjApsEJWR+teiQxk
2BnMlvMP808rvP207vLrwFh1g+0M9+mMsMGGVnHGUPvDGOaAYZdana4CG7MU3AFR69tYvwkKsfs4
wvvDTkX1TkoLaLVOZsdsdSvwAJccTXA0JONfPd5u6RR2aa3Z0wHpWP9T7JBvYqGY7SXVX+IIkII1
vJQ6gZxJZVry7hbXZ24WLqnZfy9hdrbQe8ssl6dwo9+5uAquXDqpDRI/8zfRno3eHaoXlr7eGldu
El6pg6kcHtnNsSuSqLdGgnPsUJ9xRfUkOYMd8oo1qk+FPaLF6czf5zuQQ6pvJBAZSPbC4CjUfBWV
HwZATKy62clXdOs8tLOWKTAtvb9slYxkqYBT+vaDkLU/KgwYAyLPR0OhvoNxyAgdtWI0TKK2cM1b
Kf2iQqU9CYeAUw4ADIbI3vYdMzKPbl65DtEcqWRbdLmT05xlI5JObeEobHbUOqX0POUiIf4dRgJW
+Bm7kTidRyJ1ZGy+OfyLCTwpc837vTcsTduNEV+lLPqpXizfJlVmc1FKIKaa4oDOCkWahPq/yoyD
LH8CdsIhhZAIjko/aqyk3c+KnWvi7DoH/DpqfONN/dL5Wkksh8WuPiz3zb+AaIbWmbnQk2d2rdjI
9VupCBKjm5fEJb/sZ898YABAh2mbrLXvkb007knquMoK6aSid/V6DUNftEZ6Rs1fyjykbcRgkRQV
F3FEdc498PPo7CdyBRroq+sOlVQ1mJsTi1nKhin4ew47iVnctuPBbL265kzVw1CPU0Kiqyee+LT3
n7mc2A5BeA47lm61rqy9DfHgZyLZCNNTVkL02BNu+fXteNBTIJ/LxBYja9BdDdpTB8wpY74PpHhW
22df9a3Wq6EPps8VyLFXXMTc1TlKzuP7dqMW47S9gTPCJ9ojVpGtnWE8N0WjGlFaf8Bq0jHMQ4e/
/9GJqbog2x6Vmfno1iViXgr1mzXmHFC++Bb534X9e1dN266TQsizAtdLN5qru9D5D2NpKGiZudcz
yZMW7IUHgHXoH/Caq7vg8/UH9hUBg/SZjyyH/Lo5GecO3KmwVrJgB9R1biqCubvjIw5ztmi2/k+l
UQmNUGDk6nbJCzZ81cPzoKXICBno91uxiYXgPRCfqWDjQ2J9m47KhKQtkBYVvLjhDiWgDc3o5dwT
4UHUOC869jY+yz63XLLjeHibBIIX3V8ag3XPkUnDdGppV0m/tvUwLfz6QBTZWYiKwGSEMrOZx9q+
gnsQ0LPkWfOND0RFuFbqczFJsUmnRSu7BfddMEwvKnxCKjlN9JoQnXoxqDvdY3Q/w9gssxJwCpzU
tMMaqpkv+XWduzQb2d2MLCrgAT7dbr7tuO+7sqhSkTSkScNV69vvqjEyBKgm1gxbCAhJbazci6AW
1JZAcJ3fgla7yEHc4OgmzVoVAW7tD+3NKEpXsPbT60WGZZH/jZNn3KFuQHFpqfEmorR3B0Six3bh
RCu4k/AAg2PTvPyLj3N2cKLc+QBbC6QJS97q2JqQVkGeyNktRkfXy71qMTFVEHo0DjIr4i5e+Sje
MyMWjZLgXi/EhMwmbbu1zMreZXw2L7ElCFNfsf1QvsKuY6jcMp5tsr84f9Xb3m7B9wKhWBF/IEYe
H73k68f0zUPGyls+GfFFbekV4RJwDYB4PP+eRa4Tlt/8Iyn3cHMjaFq9CfuvjLrOTMPxuHWaTx8H
rTSUhkolNJ5dRkoohoX99PxjOy+i7hRCtNgincE8v5asUzELQg62IIY5cCtffdBWVU0OEAWtV5Y0
pHugumhVnVvlbmi0SUYlFoXoreUM5xhpIEjjLrxH5lBo81BJmzKMLtwjkTw9X6Q+gPoyNuiSIekt
QBmRkzb2Ia5SJ1I1XxdWQch1EI/9xHJAaJcgTnO8TbnVDIfUNoRb7pe3dN2tegYlba0Mo5Z+/mcE
Rtc012eCZsEzQQbFnPRDIGwf6hMVG85JkKA1HLd2JbptSlOpQEKpfGq6sDxs/B2gus0Ko9AgvGuM
0459gyIaAdyFgZYi7ViylR1e1dQOyTDFF9eYEV63Ba22LJZxlw7guR33ken4yWA/Tvj90CxBzid+
8jqKAxOEt/TPmyE2uZrjCnWt7IkPMsGg2zzmybezl4gMKeCrZyDh/4ZJXNVLV3FFMQys083KcUQC
Dufti2P+/paCwbjPDJtQRbmCFn9U/8tHwV6qyzCnnd5ATI2k6TePFi0Za4sO5JgWvUY3wlZuSbj6
o0BXvZCCCCHne2UsfypYcAjQejtRw09QEuvFE2iteH0r59C1IWxzzwLaJPw/ZTmB1yYnmcOhova8
NpidewUoOCPlSBwwhNm3rOVpYkAg+36Fzw/dezVgdyABvR8MsIv8QIqAqLg0yYp6xyvqkucPxEhV
fcrInWFnYY3pVSuhS8i7rO4/eL2pVt4JRmQqjQvJDrHOR0qbhFUyFZTzddTMleZGXnaW6CkGEzj3
cVb//UrmK5OEpqrlfogFSP7rKUgcnkfHTeB/rZ+XU2EfxPtvA7PdrF7OmPc7QfuIOTZe1CedN25D
0E3Rr/rMx27KXla44CjVvgooAYtm81otL1QLKAfwB//txsnudaiCgQCnDoFDp899bo8JiySD17Y/
abLgBvRMO+QWkUZnSK5KidSNN4eXLvZyorLqRxu5Wzbfo4InC4IsITr9vuyuJAvhJ+TYn5r6t01X
ew/w/uSJIKXdrLpsEotxS1AnhJ0QwA/7xxZpQmUpUZwsy2vh5dWHtUhPyXJBB3yJHiTWFd/dkz6b
XDqsN2ftGo/AgbcaDpgLqs4t1gTGI3TLkjtrWBqNHhVjh/3PsiN/QgPfZZcR7AlwSMsOQ0qOnX+X
OfhlKeMRA3BWBPNmFYbHUHaUvLCu7gAOVx39wdU8VNPL5r4TJ24LGtRojixNQsDnMnPiz+XF7rHA
2ZDH7zWOHoY5fyV6935BL8gIBRD+H4t0OD0oj83bn8XK7d3jcRcfQv8hb4sTSY7dVjyBZjbAPmBy
et4GHRjlJOTZiUilwwOBI2jsu6GaY5FTWBDHw2u8OC0iiRk++0qq61RsZu/EmAMRrHSM+hKcK+eE
tOjhk0MJatjfh1o7Y5l0FIQZiVgAk47CGWQnixy1wm+HwybVo7B+xPUmNILYcvStTK8NFxPDPcby
4s7IiwMj0bLzwgYdNpl2MpZskbyeLo3yzG24AvTYfvC7HB5/1WFZK6q2lIUU/31xknXtjp4Pm2lS
bGYPdr1tdyqq/RAFSVlBzqWvd/4qNIrgH8rQx8oYr/nvQNh8E8c7sPN3+b1F5W33yyicGNngt7/L
kMqvMHquGUa+YjYl20vGUQvX6mPMFfQTu3awnlu8E0qpND0sFoBXdAkK/pqmIcjisRB8GeeXuc7/
/6UfgiX3xUbGl5vFTmCs9S/bl2oGVA3cGz8FxvPbjbdkx1cAmDl7sI+V8iVTwFcZE/GrNlI97wtY
07XrpcHMEArEo9kz07XRUiQt9cDnAYr4e9CUuLiu2tXsBPtfwWtt3znWkcICaVCQb+SnAt05kTg9
xJ+DTN7YvKYIzHxi1MD5S+ZXqt4a1ZfL5b4GZg0xdQKB5kEMSo/OADJa/QTEL3a74bQZmNE2FgWj
SIylZMFn5L0gIuuLrdlYJUSSPEsJH9gmd1kS+0qAZWkmeKb8yQkU6bpuPhG5v+VvnMJj6O8UCDqW
yFmIBlQrN6Yf1fPOI3sEVCyL2/zEgX3iSIMfvrZcq8X+ZAslBkCI7j1l4EqITGttig/sj8MAcq2b
ST9yh40WvDLtURgwhBhyuVTbipASTgeKHfu6u+X6xnV//bdcVJYRz5J5QIGnqgkgeS3IXXjk24/Q
mNF0cT2gaEFE3EPylZukP4ZislfzP1KXJqVweonte4JS7eAbMo140NSt16i5h+dzp8oyZggvkcb/
cF9qtBa2uBt7ruHa4004CHR28gZHrpNyKbmMi5H7xu8gm8WvCgDc/L1Cl4EEC4PiOLHjtvd/K6hm
j4M/4LKFrAIGgaKDNjdqc0uhNPyoDd4XHEvvdE9oPUmGIERAEXkriClb7GbjgZBpMWyYo2sDY1IS
uaOl6mpCq/20wpRWt/U11ECx1DKuTkf1bs5XFRMQYRX6cnwUhbPU/CswgB84p9Gp6uDgLS+EtPwD
lRBP+KiW1Lm/MCKmvidkagehdJCqTEPfB+8Y5mt+xRkHbWZAbsTi9USR+KvEyKosRb8vIxS/xuX+
cZeJSiDFbmqFWk1suZQGIVWVW8lWD9cOPStD0p7nLAWk+gVsuNVHJUQb9iet4K8myYwxmKJvOoJQ
bHOqTES2pr5rzrcUqfEbdubO5tdULeWfMuFaSnFxqMLRnPxLGgoyEdYSOZMEPANGRUkDuXF+8XPa
37QguTAyQP1ypERaHijsp5v4Q/nctFD9TE8lnhjd1az1MxcQLguoGBey9s5UlTkS7te1fux1F4jw
nifZrGdsPps+jIzG8wzJEEsMV6lvY5yxsP2NeXfDNXp4D4qQOHJ045CWj7b3X4Lm7775DkOUh9yB
bcL/oh8pwV3izYoKBxmUtHHSf31iNH89peydG84e+qDIpXv1N2Csxf4HCkCUrM0uAzPVreoNYFBW
D8SRXRHZCwo8DXfXs4fKvSXT3wQIjlz0lIzB0DsJMPOgFJXdJcFnQFULb0vss8HGpwD0an3p+TF8
GXWU4J//W1mvQOqVSIToq3FFyVwbXkPWHphtFB5S2U6lAG0gw6uFAr8ycEV0HxIaTjOB6v8Ye5p4
ccxdZLZ3mxcUTxytvI+g7d/MeZMDYSU0N7SMWrOyf8m5Y0Ck/sj4CgOSCS4PV8GmtdlahPSuL9p7
bSWsWkovUDYj7+ZzdXB/wwDV13eM1WfDvsm6u31W7aT/0m4M1+EjXbS3i1CILGgEnwxs6jeHg2GU
avC7XOD77o0lpylQKR4wcI5dCedTcWFoA3JXoHGx3Q0K+Gry8JjoVX7/jkNaIDRp9ipopRMEP3m8
orn1J2tfB4IxNUJzHjyf0W95B942kyVlosF/M3fE8TMdHj2sCyco2adjYPM1FUKxJ/CTsGRL+bnt
+wIw8HIwk7AITvs/UEAi74yzT9Nf15OsjkNU5Q69D2qmltYVJLJMk7wNgW3EKDxVqjP9yAqAvAzV
4ahZzNRmBdcQ2Vt/DAL5FnmsqtSIEtucD5Msth6WDTJ5HZQobTq/darRITMF6oW1QxmWHiWXXcn6
UxLvwuP5RI2UqDupRI2UPb/Gb/KH3LYNrlvVwGUBdMZNaOhRg3dLVwPZ0Vd5yUDt12BLen0j6TNn
jSubfTyWyX0ZQKY8SvhysoSWwJs3Xa+UqsE+N7e/LK5DGJpq4Vj9FnWAu24UeU1rJ5+YvM2Wdk1L
6qzRX0/1ASox9cOQsYjTwycnAkrQFIsf2Kcz+H6oz3j2iwlhCzOxyf4u6d9sBx8Zq0tnWp/NzAy4
DyY7VIsTCGTGqyyc+VZxIUSn0+8c4C+9c3mwbiflXWahGwzmp8jH74HP1vAZeIfBv4MkgN7VVu3X
iyKdG+F0zodJRxTXQtjD8hLdu56CcXu7Ii8gTD8kUABL1fojzfKvdDVEhMp4h1PPZx++zxaNCdtJ
f+LbruAMstVc6NJWnhvP2nEQZEwars34Ko5ESqwvWJNVYk2iTN+mBTyO8oSasiz+0jLPg4fFcHFn
fH2cMHg8tLOQIhN1gBNzua0MEikPA1qvyxUBQPWF+BGVdFPQPT8zC3DSMJZZ5e9KBPGQzle5Q+Vj
RSHeHyDRhOVt85dybJ/whVITelHMgx0dblNqBoZPbXUYUdKdVnkG3Knw0g7YQdAbqJtMz0BZkf19
ASQkKjd2Fx2btI0EZQje3mtEurz2pbGHpkVgW99FHqpN2vchGCBn6ayQTPcPzB6n9pQtB+ZFXWgY
CqGccSqygBgRbM3ji9RLLuRPAy5sZdJdRdT2sAcktvsbjNadGTxYetJy44NROiYXA6WAVOV4bhDh
UF+w+pO6p6UXamaTHHQH7yiU/knveTMmRxdJQuVxVxMzboctsODBgWual4V1qVGJfMWrmojEDI+H
Ha9mdKvFdM5wlty/ra0+EmffWukpVTMbjPAkrJ7O0OwTOPH4Wl6GfAH5/9VGeRG20yuVYN2BmBrD
pTIo5jpjdUSwjBnBMaQBIHeK6MaVM7IdzRcx+xwtoWQhPcORJMMWOHGk331shkR8bMqPExfivZ5h
SXs1uvkJNlm2/JucrFsZh79pE+BSB3XGe24M3ZUwxkSEcJ/3S9qEec4+8/W+Orerc7EOeqMuS3Kv
lfQs6ffBlqO+gBMBff6rd4VJ8lS2/4JDmCjB0TXhi0v6JcEW+tBHwj7v6c0Nk9oc4tfOPZTCDK5g
BE/CCnuS0yozUv/8xs6VDnOcg8zJJIAZNzhovwWmy6YqS+qUlpdifS6vWGxVqrF8lEwVZ6YGRAfa
2BIhqVRVY79augRYT9Jhvgaj2YLM6JMJmyauH8WNhI/Cr/9Qj6B3ZwGlYoV1ErM9g1xPpIIMpaMW
+DeghaoJueQPqldAJ1WDBp4D/woyf9gX7Kn4MJckZJA/UQKEp840uxBygPrUwPkH4PJw3Sco/HWA
hPJl95nFYk7hltl7uoFvrBPJOMdP4Yd58AYz5pPrw6l9i7oRJXUpEuJ0m3GtK6CKXpm4fMstyiPn
DUdWATvMobBxfZtarn8jbFl6FGx1Waorep5Rk2pIpdXlvt4phJG2YEF1bB1Y/Gv1H3tL/cGFC9eh
TzG0q9+5nKHcz0Mbzb4GeXiDvYhN6JF9sXGqUOVR7W8Kv4H0Dw680PKNNu/L4yvu/MP/NpPkAECM
CpYtu9O9ebAcnqyezrXpYc5fzNrf9wHFi64nZ0eeQTvgIzPZ5426+8yhvw+Z+WpVzNbYRHV19elI
npckQ1vVA/Ktlayf7xB0nj0IfjpeKE5gW/U/ojbhRHGYnhr6/I0DMlcLiefnD3snDZ8/MNW8OSS0
gAPlgvfztGAMd5MUZBfCq+5dEJxJ+LcDw/Qsc8cfMILTDU3v73PP0x8BB8BOJ6s/ERU9UgyYkP6B
qa+nwg6YiCl8CuwCvtIXfNoU9Djm/pBZkGyze3VWflZ6ywTlk3t2iLVP+PVuNRBNW3/aqlOEv/2g
FWhNww8exUIUjImeLwCul8CBaZ54H1qzbAxLQJUkgwEI2W2jfyvhqbDBwTlA62I2lUddONP8Zt80
CVLR2rKTI5dlAoISku/K3KyKrM3+kM21ghv1+yrjUUQ9NimkvPJhTog/Af0BWauKVi9/ORv4IHYn
TQiGoXaNboJN3DLm7g/ci/kz0w/MLGxE1rFrY9yAFLRBCCb9Hmd0JLOMN8SFBiCaPgsd6xCGxqtu
NIkk7NrI8EaPujkmo++E5AVaFAIJ/o2eQTh/aWCKR01LlNFQYCedGTi6omSge+rnmA/bl0+UpALM
Np7srwWDJa9Iy2uaKX9dnQT5rsZp1QLV1/wpY3EZTey9boUzv+cHzzhEaVq4FBJOudFyXxdkN2ld
bBV1zi9POAk2N8UTMW1FMxE+bAWsQgycuazn2cXmLVaSvtQiEsHCNVK1/08dNvGvUMrFzbCIPBY+
P8sTR14WgcK6IyCZqcm2Ikops+jJSQEjMolp33kFYYpQadoZEs7+w6U8iH9/12hdCfUpkoGQ1o7/
pP/gCiRP+kYuje2aHsAviYLdhbr+LVf1mcnqRjvFSUWEqmWXHg1nwn5eY6Cr+U8/fdE1uRRWLfgC
YdjEEh2fA7Xrt3qpvHomk4vruZRp/zf/qfp6wYU/45KFJP6zSZ5EJjZWmfrD3kEz7fA47KIKL9hC
QWpHkOgMQNCa1u/QnmlDz/SDZ4rzAcDlkCIQ/xxMQ8sd82Vle1VLdnzoQmoln7PvrVTzs8CUcRfw
9WvhSwOdA2RlJrF6NthxlBZtyi4W0pBBRKgOClBbddHRW23R3MySf8BT6tbCSiKFvj2THI5tUP4f
9+5R7UGHq1vdLrE4Lyx7CRamLvi8V3OqQ+nQmPOLoWBgkyeklZXSZGCePZSUyM8V++5h2z23bZzt
MDgLFJFJHHhWkM+6NIV2Uy8JEmMAVcGaW8q2haIEV9WLqXU+nKz11ZXpZon2djmfcC3jtTj2is0D
V2sLT3iwoEt6FsnYRRSdBHvrAE2vI3I2uql12+DaLXI9ZhqCxECSaZ23gV300F7jmdm+JifYzdSP
UybPwNepUXlUlRrV+gbVbtFOdzHQ27cuIFDL5zCgywrbEN6rv5yq7gbzKLbovd2wfnBOQKWMajoy
Rmr7Dz5Fu3MiooedkOP8dKGzpBNKfIc+Qh4+K8gD+mi1h7a5jY4pLiU5kktaMq4jkt7emNphXsel
4YVTZgvK1XFD+Lj0TbBcaH39O8NqsmwjRSy3UV1fm0+/yUyjGy7WkqcwytaBdQ5iOra8yv/HgK1q
OkGZVKt3jduSgoTXBHu0lV85kOr5Tb5CkgbvPAVMzoAWz+XSk5kgxoKBoDOX6C8lPMQ7cAvM9/4O
t4EZLN/b/jijUMMUKpB85BcxA/6fttaFiAPogvkPx2SCy3jCEL2j4FlXr99pLebC/O+DcVoo6NZH
UVcepfAPZPQyEX8whC56T1z78UGuzL5iezSJtkTzjOBq+3AY6P9z+zT4SwRpw/AhO3RPT24RXjcg
cbHbqMsqQHNkfRv61m9BBm+9mgWFo28YaW0nRCKK0g9W4wzGpCIMGQlqmJ+jYt/XfJLn5R1aH7q0
UlaR2gK9lmVD7MXQDZvcHeA/xqqIpyXILIBzGCikfinAkS5xChifj/U2B83mHr0kMeMATQ94eSay
bwgs+Qn7R3IkGt4bgWahnHSYOsjRqHRtvgaueHC8dA/HKIxcNgpr9y9/DF9GU/ORfpDRqaCYZ1Z1
pBmO2dVnsKWdSyTnCqLl3UdY8w38U+/h0sJzIge3sx7UQHQ6B6pclfeFgd47X0BGGeZvaoyMlQbe
+WgN07PM80HVcfz5UsLCsRa1tjtuaTWMue88srgjNp7YIvpR1Cgm/SwjLlGA6ac/qULbms58Q09g
FiYTRqeJsceFPtXSoEF6r8e++SrLxIGKurGyt2ujTe1c7PqRhTzUwsL1ZUJ91HdOgQhdvcV8pbY8
mlCqjiDJES9fi3X8ymfNYdHS5ouj5DWgMw8rw3HOKRK43eTi4zyAVqy0XuukkPYPjusJ3a3YvDqi
KJtlVKKuFCMnfAcATE808DNC6ukuTZAFmBtsW9dGT2L4aMETO0rfcitsGqwlEP4PV/aR99Xm+cXp
G6rvosfLqawQhifhIPSr5SGx3foftcsj4ARFoauh5q3TC5Xb0GaXIrCbOd7eigfqsJVPUKh62n2B
hHxvQzHiduzAOTqkInpc0d4ZR146O8jw1s3TtFaBrOWh1ClfY1CgDawVivBpM18iZMFEIn79oRsZ
/C6Sfp7zOZsnSYqAwLtJHq3ZlkQGDQ2CGbE7P3NvgmtAjr9Iw7O/pI7FrpG7vo09j2Q2eqUdg9HI
M9CO7dMK3SiNT/1PybV5EXGF2Zn4tNd9XXU5XKA8HDAsnn5fAmfrrf2bbKnoL2sfOEwqCHC1joCz
MdPc9PzflOkRNG2yYxEQxqzW2mSMTsVzqfS6ScmEfrzqVRSCfpj2MAk98WjsCPGcGxH4YKcB2R2s
p0XFVn1Z3qt1z/xKRk4iYHhTTNYG7jVVh6ZILmvGI8Cbn/9T/Ih1qBfbe4eebE2GqUnSGUdpc5PM
y/A/GIUNG9PngTyKdRkg3IrIjhunqK5FBQUbTTTqFHC+W5O4iNJXCOIrq86Sg4IK4qtEypHgVW+n
S/mhjSesogQQP3Hej+l+85YHQLmT2uXgsQc7BRGflaBd82Hwqr94Fdzujyn4GzOZxXYKBD8WM4EH
cem97VI6apUlYhv4Ct6f50McmL8WGNVvGOXXii5iArXm5BFSCMRRnkLXW/TDAvZZsUJdKxg1D0ul
LkDkQcGS+HplyJQWADcKUSf3cnTQy5Bm4YgZwVEGPDGnsWnm7jicj/hiLmkb8tD01S7CbX9mVEqd
PXWx/Z/ztApMXi6cRIsT6msw0+R+9Nr1/y2gwNFSzgD/D9mzqDWBkT/+nXWiAbqA0K/yNkwCXWiI
jYyTRr3erxmGsLMNvwQQnhDqJvEgySWek5J5yOhqO30B82peLIfHht+EAcPrRUtwErXd6P6U3SP/
vGy38eKa7Gye4oVXEVzzBnX4EHvdiXUxQkdbGdS27cSMy8kNVc3tAnt5hXNL44p3fxtm/dTfoEzA
hvmLDojX5GdTQrTTcC6mktYmkkiEgjgaovOwDhn7zuw3gD6VTjuNziiSjYhpqLpnAkedcentFmWz
Ee0koHMHs1Oa5zr16sqPh2d/hBcDjCOOjmHinfLg51U4NBVZkbZcYJDlKFPqZaqVlwdh6IJ7KkzR
b/TsMEU/WqVdLiJdvIBJ8vr7yjjhv/6/VQ6O6AZd9ayWsk3mqkB3zL0ddiYnu3Lg0O28RwhWnebm
PrNOLs0fesp1aId0KGg52q99Z0l5MI5fmGYgbDS5NOgjFHaFys+Di/RekutB6yGLwr5kAtnbCJRA
bMq2Ql8Zf6q2TH0q4xEWu3UOQI4x3dgVJptla3MnLF9WXZcPzyghmnAyv5vaNlcFnfJ2oYAc13qN
ZKlAgxaDCVoLbZ0wbDe4D8zrHCWLFzFYHbFuJele3OJ4ydiy/Mqlrx896oN5hAHRDgFRVkhV9Djy
i8PziVpGIfK4zWK9IWXx8sQ9G0Q/tyHpW3b/a0yp/AnaBkQphYj2iDoTdTKMrZVJfvwAIZw5LB7P
Mdu+qaYPvZsDr+LHwTTS4/V32JT7sc5HRJe7c0t7FG2PMOOKX4ZCK0+vzunSGLA4QVhPjSk7R5p2
kQ2VgdNJgSDb5oKLXeZfgzoGhkIgHJXtc5TcazjPbywxXTeRNb7K1nWBATkkh87rebOL/Ydh3rRA
+ByI6Acenrai46dh13EI+z3TtEDBLN1TceUdGAKp98ZIcqyedu93N0IlaO5Haf/VRrv3pQ/QqZqR
QjFAwlMYRRMqUJmQtuOvIa/3v4ys/9JXph/dO1nMH8W/d5o5RyQxBeBe2THMrOPV8JcEOP9j5YGz
empwc2JbXLmqz5cdmYbptcvy7ndsSaw+ErxbFnrgiLCjy0bhiQ0PHnUcWZ2IxhhPNhzXhmBxHPur
W194ca2zuiyvnhHLcro2Yv2W3vxpnHFVUHIuX0n7sNm1p1OmB/DxKGLGOia1TT58IEQMDeqK9JIG
p9GYRrBvqqEcHdm4h0xzyrN9ncNXhftyqq/vufrXoU2ZF7MYkM7O5U82nSvt00cmmR7rfFPMehpC
5QgxoyiA7BlFxQnkiU3yLZJAzUbSrmDTK8/czRkgKI0tO50tAvVR6LHCKs0dg8mhlNk6K9Zbkbwf
IOnh9GljsEO883OSx3wNFPA7juHEHKGZHPkPLv22uuarbFIgjnss4RY81y38JhK5Lr70LTVrbN/U
BDno7cGe0wTuRzByNClht0nlbdQs0mkrphoEVPqhoJg7142lpn6PQACesaF2hpH4f47oyXQ/WpsA
AIr4MPXQbO+C+ozq+Wvqi/Ri3FXHi8ieE3v4h94T/EsWL48To4+nMjYrKHxBmlg9sAfd/TIqZxvQ
pXIddaUiaTreFP9wyOCDhqTASurV+cHK540nm2DtQ1+VP5ifIHpIUmi0sS6BgBZYDU3Zm7Fv8WBd
sM+UinwOBWjJlVFSqj1jFXZuh9WdcGzVTKPVhX/x1PEdwiXF7bJb+RbKkeBloxIh3xz4+uDTcu7C
cp7I0l0paph6cWhUyALakrM8ek6gaEOsxywhdh//rGHxZCfHmilSYXxHPhgIa6lpaFkgAnuEGEUz
oPI/WGDpqFYIKA5AONSaA3RFDiC3vDdWiEcGc0QBP8wb9uI4JwAfShyFh4oXNtc12ijhPjpEa8EE
6M+4sGZcVkh21HSdDuPGpv8I41RAqdJkLOLvlDlciTjijFRKWB6fCwT+l0IpUecBAUPhpXX6WAXf
LepClUbz+KhWNG4vBGAiLPXKzH+eYd4j9fyoDo6Wk/oQ0OmNlmFeccma+69tkVJDJXZKYxNFK/29
W5gq9Y23OERdjmH1LbFzAS8+Q+oDA/dj7Ut9CP/2rVP8KnppgFpbDwAAS4PLhyqnEI+qET+6rsd3
qRjU0Kw4hvxXTTUC7fAIlKgW17W6yil+HlsMvebEOu8pPvoU/fSfDvrz6voLEbwQQ4zNbA7wNgYy
kvLn4Z/ucRIRzYkiB8udCfrVy+Lm2IeZqcjwegHqpbLKgyJVbOUmw9+cvZVrZBBWCr8SHanxIL/7
fiQdPEw4J/hGnPiKKgJR/08Me8YkdVb+sAETDdmRkqiYO1C3rb2keGT7cytkxm1kfcO47+0M59r5
gngxy/G5KjqO9AMb8vpEMWLVllbLn8OyoOZycTiBKB69/8dwFQiNBeVFYjCZ/tV2b+qLn9WgpFl/
co4BNDedmxUhdo9+J0PYTND5qjHoMgaycGpkHiGqVLhDn8da7Z9Bwg8Lo4NlF8ZrhhqIkE6woLB6
1NkZM24lxAROG8f+QC7gVspAkdi6lWkOA/bz382trArPNlIljk3DCOGQy11Kd04IPfUNQFlhnBLp
oDKUKNW0uIYF0EMocfwLvnGHHm6h4NudFKcsB9fk/jLEvFHce9GQdFzGf48WnWSvvz/JqXqImUYe
yFIa0KDErlRlaLjKSXrmTDsDo0tIartQAhG2OKG1UJRWNl/eB06zfxt07zEt+X31hMOsW31SYjIv
gsA1zmz5+gRzNEs4XXC14heK2apSJ1xNaeGJBvhGY6WiPYGxDbkB+JJo1gAn95hyEnbigzCeB6WH
y9VN/CAic/ZtBQUvOIUaqsnPeQUfFPsl9UQe5PlgvW8zAba78E7F/CZBIzKXAy0igH5Ek3HGwI1e
j6iIpFgAjDfxOmlXkhEiYb6Bf4TIK813Bt4iBej6qG/M/WyL6Mja6oAOFjrh71h0603vBBlXD45m
ZZfL4tFNeiqqGM//d5N1/e+I7gOiJ+lMe0d5lFmq5HKcfRsxCmNl0NpDjxSn1WQ7TTgO7mq1n+yJ
E9Epcam8QoWELZseVk0b60h+Axe3Iksvh1s4Cw20OdvIfGiNr84rZDDjH4bZmCZtcJbGP8Ahju+n
YJZ3Vuz4RTd7+xb6uKUIVCy6dnPCXyXncWgcLtaHF23PB0DP3IK9k03EyySvenfy/e6s6z3nj8q2
p6AD0r6+V0sUlRXLu5VaM/1WkJS5Ex7o9P34hqvf2rjCXcKlAVEaCqNVzK7CkW5/AQ03MofwOlq+
pJpAHlZ1Lc9YultmcLaTIjojCdE8qMvKEVtYCmzio7bBsqBmJxE9awr/O0i59Lweg6qo1AaspN+c
TGIuFZOMsDT4wnVqOkyS6h99WMapfhzSbZW3GK6hl55qLUoN4+IJkuUzlolZ59m5cXFtNfqu3Ahk
sKs7rzN5sGXYuhnG4Sh8Q5Z4hFNOrZaKRrfbfIljLyhNOQUSGMmybb+xlJ+hiTsEZ1t2Ff9CsQbb
OAQT780WKmIygFmROr4Qx2CGk2K8XUdD7XA+Rhs9nqt5bFJ+82lJN+9q2BySPJrWF5loa9MUhurd
izPtve7pKYEZuKDYDAYIvfH5+YJ41E77tbFQEbIt7Z8MBSZxHUjml5t8WPlYDn8ckzuOn/i+XDUO
83HtnLBiZMJHnWbtBhu1IaP/Cpo8YLwoyMGQymgTmCclmRwgRPi52SBNvp/iHYqmYhIztTQgOdIo
HHBGGZvdV9HzfYd/R8R96fsUiKiV98nBWqALlFo7ccOOBncnmH04R1BLcvofEQIqJbH+l8+0uU8z
5VBC52WpCMatzwojkxF0AAOYxEYvVOd072qYeW47QbhcDyTK9fuE0l0VYmpd9aK/3fPISYsM/SvF
rus5uj7wbKE6+nZYf/gv8+YgnFik7S6D21evP5ISTVn64SU5fNK5hHKZMRxbb67Q2lojhcIvwSUd
BQnRAz7drl1GDmE+4dSwagJIdVFTIczlLtGb0QTojK7fU6u9gnz/Pw3Sia2BK0lu05OLvUib7AM4
uAO3RmDaTfGgTOtYtLH+BH7IjVkgGEbtS/6Vilr/5kmmXM0Nhu9bU2R6jklc4EZE9qlQXJ9kDvpq
IwOeRWngl9rKhzw/t/jecXiBg8oIsuexEQMzTI9SRx5JpOzuObfZqNyfCLzNjcMc4YZGODQeWKel
ggZMD1WRlyp6PMdid6GcjDyvUCmoKQp93pK+rkiFimPGCr9uLzZ0zlmST9khgv6MEQspQ6yYFVt5
+62bFtW0o2y5fQK67SoAwSr0nGdeTQD12HhlYrBHYQWCCS10FbEWJDk6vwniyaNsDTUBaQQRDVEG
3BfVYRPQoXIS42GBF+9wCWL8XwLrZ291Na4r2E99SSdwqjwuem8d90jvcK1lkIADFNX+GM0CPQvh
pxuj7mtRzW5cpgPiUVlrZEH2hlOVMah5t68k/r7BxbdtxQ+89ebCwCRcIZRD5AuyUDDgej9Ho1Xi
lZiRNrjNhCWlDlpH8m2+0UY/p7N6PUaKBd9FkiySKiDX9q+T9/hm79+pBKiDxd4DkVS1tdn8tfe3
WiaRnuVbU/a7mAH5R3hXxFwe0Do4P6wXUil3yOQtkpHI+U9cGF6IUSfSJmdI8zjiyz0tSxcasGcC
GnJYZ6q5kBt51VWTZ1cv8aepHFhB9mhzamsIlnkzPwYkiQVaINODQhCfuypBRew68UsFbmXc7XnO
K6ihsoF/D/03jDoXxZaC6sE7bESHmntMR2iok9/YQ8Bz7M3m4Pz4ik3kcxl9X/09O05ciqWdnyA5
lGqjpwwzR4E6sjN3S28GNIF5uPcpPJFm7TXxTmzJ6ducVpUkwek7BSUHSO5ENYNJsEIH0Kn1Q7S2
FfdLctkt0Z/VpXhfnrdi6DQmsOgeln2CoiGcYDwqU5cssj0gLp7mj/cdT2dnpUugzpKCLy+1IHXj
3qzEfHwL00bHFRiQkB3pNF5l34zpAGao/nyxu/qaQZ9QPHbGOAmg3uN+UMPaYLhEEJelHhsNAK2I
hDdBHsXTtteV8GyeA2JnPY80ixZdDosQtlrYZ1ACIXoLapSsWeYdNKTK667eWg9wZQkZa4QX90Bj
1+mmWfeMgebc/khZwKBcjTnvwG2H/53bhBIa49h9/p3ifIXzJX2nKkUTZpsHZg5x3CPSJJ+WaC/w
9ICy5qZ7VY8JfuO0hQaFLPWBm1rFYuO8pZwwKd0odHciAlVDkJRKcUmcDqiHuJ0TnF0kyx3wrOfm
5gcr/JUWvZC6LzvFW2CpZErR1+BgfGQKcgas+28gx/v+lPjUTS6y9SXYDlv3BjPxSF7Zf4nEFDLh
+O3rmHw8yn+IBGHpj5SzOg3ouVo10fwbcqbDvg1is9sy5nsmwbANPtjGDRK9+mXfOHxEZV0gX8vn
iTt5AdenKjmEXn/HMRBx1nvLZbFMTkmwNzzPz0LNCYoEXEfB44/zTJcN4tZqIppDgkYNkeoR1Bpp
sFk5pw/j5cgGeIZzAw/6eoh+HN1ekfid96jz75tt9M+lo20ISIr6LvVRht8sIdHfhQPEYbsJ6U20
biq7RtM47OZ1sXOXx/S11p36qelWgWJCmK3Sna01IDzcEUadxiojkziRa5MyvIIR5CPB7sbfwhnd
BGMbiy2hSkeJCceXWCUPGop08BsBHcQe4hkng9TvjEaW9/FtxlVqpcVqmOxfMUKNwU9mZTav10jW
//8DIJs2uojSqVwrZE+w7Rb2d02Ku6qBpf7qUiS1xoOqk2M7/aA0rIpbXo15PQrFfFzpJCklScHm
Ds/zF3geldWgVknkuPSQOuAgpOokZklKkw3cfPGykqVOQK8rYUzDS+WGGPw/4FMtMbPrQc1hdbNr
aTIhzNR7zgUQjkYdoeetj03NNu2vsQmGH/dypTw3+A6iHUtXbnIn/0wsOWgMyw/q24RMBSSgnSP8
dbgZV/7EWie2UK12FpD5V8afpCavS7Lhe1+D+ecZghRw6sehOYelGhzc7q4Z1NTSin0PqBg+mqhw
ePB8/yhIj/auKSwxAQpJLG/nqUwMPBjEvionv03pC9JhPhSGN6IsyuqMS8w1Ozp34fU0slWxZCVb
93CwbUNXcOh0h9f4NyDzGmH4Dk2noHJDeAX139V9o0JGtj0nRfDZy/i6iExaZ1PDsghNyCkprKx2
UCSJWNuGI/LZVJnqCJoamSfDwI1vSuQbVFpMB/z28X/BNd3gUskTD5wynUuzUWuM+tznWom8CmqY
qyb4lCAjuGAvDgLRKVXHlAAFM1KMjWrUDYf9XUQuN3+UBNx8yzHeNQMkCt+ujeqV6H4+pdgOFK1P
f9V/j+87HAGPu87K5epEeu3ZjLCgzQOZym31hoT4Ygrm2AOkwtOqyCCsmKoqZaDFKZJI2CVp3HJB
PsR2vLKvVbokCO2KGy3uUYbJS+DaehehiAdN9frR1PHNB0Kmp7vF+HWzJukOY1+aXYnmOzL8VyI5
g/GWZL3QfdYNCutVfR4/CUkx44p1lt9tOkIT/O6wmjFKmBCfEYAAQfnuBn3Cyr4LSnIT8KY6y1lt
dmtW2byJnCKjeKJGXwzN7gVczpciRSkDSECIXqhqkBNQRRy72qMseeW9JdPmWfX3itdhZoNt7rFX
M4nlrFg8RLqAVv+wkon+OHtKJlCsyBqy1D+bvOVMCrdBFKV7ND9zYv2HQfz8L202H1/OksNeuyKB
heK18UuROv3upiLHePFGXzFmszCDNyYOQcQCVmqjUd0elOQAI5vkpKhJcDWJsga2eXJCyl/rppzm
ryEi7W6aPXzTh5GLN76oA+xHxoH39QBlDqa6GAAETc6ZGSvm9rle/NE950cq+78UR8hpqpBcn7iG
DFVdRCtp5ihoyYTFCR23Z9/QZmdUVXrVMIFrdfuf+ePQvl6wPBc8R3HxAiY/he5TfSgJCH431YZG
XKCb6w0XEDp1VBDgDZHnOrNNt6C9o9g7vsGQh0LfoiywaymldnxFNSXsMs5/R+wuaq06gxu/tV1z
F2FmF5BEosEhCbEPvweR5ZZ4vgBo2EbmtRBszmrAO9f5JoMvYUdUBib5zwDfdTD2bWv2gh/AHp9d
u2dz+sXWNxhYHso+s3CW8aXTKpADlmVnPx8LFCn2m00MmIsi+6F5Yxfhi3MxpfdvpAi47T9nYGEo
u090lEE5zE7bxDemySTfup9/LmaW6wDaFdgUDJMGT9NKczgYnB0poGKNYcB4wNODC6t6oVK2kFcd
Zm8EbFqIg74p/lh5WRyfcdNlbOkSZCM6dZVACua1ICjzPaNI2JGDz/nF2FOUZAlzYIQiu95PuY4x
3oOoXVZMIkWgl+GvtDJcCl95htp07q97Vyj2NkpYbwiVRwnkm5gSRsvRw3pF+IeXcpYuwqYFAVtx
W0nJGbS6t1DXF0+vWT64jooh7a+lCri+xEYCB3L6WVEHFSBhg1QMvQf/te7dV105QNSuWXhBbPZ+
s/YiBcWCA41ofasP1VTgr75vLkiFX7ZB7BdnHoebhxWV2MBXbhEaqcbgoBThs0oDi2dPpltIv3Pq
e9LlGmEK16yMXeEDD3s1fgtxUf2zB1/SKK6maPDUSLGsav8BlmQB+ojlo6lhVeyLdl3K8YQRD/fx
ERM/RZXbfrCmJypyFUUpARBHq0ICoQ6DZcY5yvXPpo9ab2FU8NUxWyRf4V/kOOG/yWhu+CtaiN66
JxhtNllf8o6NywAXx56QIkvVEJV9oKKRaGQ7vhw2MOUWVPWiidHfrXk+35njPA4aqQd0L6o6ASMT
OCrJzbAWZoma0zyzT0fTv/Ro8RJUpwfpPMEAC0n/jMpROR6Ap0ZT/Tksw/Ys0zuQ02mYAUlei5p5
/nVkUslIBNf/uOtBs3Qvkn89sybiAi4ZPTBGwwDC+AmKeQk83CENkgm8Sku9LcNsd6qi01G0C2nT
PWETalLytk9Ir9KifjBgzZ1pqD3fxE34BumJ4MLvRjWLlKIKBnybC+Brf+YsAdqvSdX9R87Dx0L3
5l67EF+KrTLA+P+R22Zewkm0GOdcmotZF/v1HjHawbs3Sg+LT/yxOFNgZZpGD+JXMQ8WvCg6MQob
5fUeRasjEIo7T+qV9DMKPW3DZVGxf/4CoTJjTQ+EMjucsJqzEM2mZhFkkCJ8dHVqDQhl2T3gEbuS
lySemXNFtRg9K8QLexq1NEvG+QCIfCZUUMOHbkW49c0TusUIRXTW8Gm13aYQsI2LBqhhaGNGf2eR
YOVAtDW7KgBQusmtKWoRtAmUOQLJNjCT9F6Noezx5TEj/4HTC1DvvgzyKSZhjVBdWc8mFNq12gkR
leYRevq9r/fp2/x+peV7uqOaQYpFqr6OM4dPAb2iUqGwNU1Y1ZYemWjzllSprkYlQo0Rm5oOTuBj
Z4GWQn1N+KsJzN2VO4J+DMksFWZL0AZZtJOG0N1Zw42DCpGyR9Gxb4ABNKAfWtedDbL6Vc2kJ5Xo
VNgm5yejdJ7BL78uwYuMjhH2G+bPk9aRYOrTTlSZtprfAp+CX0lGM+DmLYkPGcYW+dyZSx4tsuE+
KF2Tcy0Yy6a9Nd2xtSTEQUmsk6ZVrBFb0DG75yZMLrcvB5pugVc3Q/GvZyvsVbmGXkczEod+HLVN
ZaTGpd1OC5Dc9fXimNF+8gEegB5MPQMxI33+XmQ7Hf91xtwOnTRxl9CKVM1NaozzCQOHPokcSscQ
aXLIGbzRj6LE1JCg1EnfyyCOX8CSdEXV3CVn4sKyfAmLqtFRG9yj136QANeLe5I7du20sEDJCDCl
o0AthzNliZ6r3iodNJVlH5G3iOSwTyMR4rREMN7fO8gppgIVzWsSf7mVoZcPsuqrPjTl24qo7cBO
03KyFhv4lmUQFKRN33gtq9G/hf4SXJsiietBD0tVtlnwvaX05j2tqvlj8kHKzsHLkmwu+F0tWV2u
Idq2ryZF3oKR17WgF/jMc9zkQGsEGkrxpAbLSeWG/l1W4aSGsvlZ+wYFglRs9ICBsYTnMGyPnSPZ
aY/zNACSLBb3tsP4xjqlAu9ywDQ+9eI9gzqXyfjPrbjB5Gr8JhkQ5yO7FPuKLB2iZ8YH1g7i4pg+
Q7nwxTARUMFSh13wFAsSaATEEZF/L45vBZTI6zlr/d6L7rOBzhHCht1y+32U4b03M1yFCYe4KI6g
oP4F7lmkyFEBbsyLYAGQ87pt3qlplqPd7hVVpSJsxv4cSC0/wWAFHK9xFvp9ziF1u+w6q2OcG4MJ
T9DKrdCf7Q2hYzBIV1MOQf0HfQZt9vl+D6j8ApnGRT4hzM0IIA+x2x8LGTXZDOREGF+PECOP6FpN
AeeIAMZMXsYSpTlebCHVra6hjQKgn3TbLj3ioqQujUJm7+39LYORiEe7DXB0FfbuXKfGmalSeSX/
AeGm+ve4RZRQ1DKTLfdbp2ZiRIPJuUgFxMpIUV4h+/ZJChgHQfzj40VyqaZadpSlP3jcogIGGdmh
OeWEGguLj3T1cFW0LL/qEO2esAHGwtD4SlhW1rb7KLtBBkWcbSk9If0nG7abZpSFprtr3eIyMcN8
5qSYnNOcL/pzbkJRzXJHW8zzFJGKZqfo1R6lppo3fS/XUYOlGV0leQC8sAkA/5CXEhscqDMwUeOL
o2lyrGCdDd4ZGnONu6IoN65ncn8rkk2e2fVhPIjVK9lU26i1puO6c1d1zFQF5Qktct+dXmU3q/su
yTvRXjtFEIQ/JlqkmuEanIOqmY3lynqLREb9nZ3AYVB2b6FSVw4qOvYFimPE9lEbU92yDQB2NTBl
GfkSHCkyV1Fu94UjvSF4ldCQyVgM60Q67G49molaf8prLw4S/oGJokpLfL0jbG/cV224cKsjUyA9
xH62kPuGPIE3JXmdGrP/XISqvHp4wbb99zjVZ8vN3sJGjW+M1HYqzkQEXkKoxVQ+XrnG12p3CN3M
zBX+NmOy+uqEjzJqd0rVFzq+2u0XFq7uae3Xz0wJTVncPmEpWqIKxHgRybboxOcDrLVr3ETpVCwA
zK/HH7FLUa6ZklQCmVItdobbA/OM6kwo5W+Lo2xzvUxvqWnFSlZtJiNUgiSavbS6YnSbo36M+Ya7
K83lYqEfZH2QNTeEm5+FacR433ca8X6tN8xO2a50KiIclnbPb04BeS+S4RrUnMtIMii0Eun+PQfW
UkqXJgNhP7FXUXUpW8zCiocYvj8ZaUp9TMHWgE5ZgXWaiwBEBz/rSSLrQ7ccXUFT1SFVNExBPq/o
HncYBj3xmun2FzrRJZnpLKVl2NywDAVwkDv409ajwq+5LjyRaM+LSvFdb/gKJYyPvG20Jc49lO5r
HUe+f+JkAVLmRki3Oo6oru9PQx/xfkC0d2HRHMS7AiKOyySsv7D4DFjlsMG6mq9uhgENgYc/IxoP
h0BCXvRzeyTVPqpq1K54tf+eviDZjQT9PFBCU3pUKG/QoqXBtubAm1YJWZAErAwf9HyHVxy7Z459
qS27BmNsT3NnuRCN2qizGC9Ktmih4OsTUcixxPTG0Q/f9NXymCgvBhG5kJuBLmcWkRmHItHn8myK
WAlDoaWjIM0pwmZ+s7Rs4t7sB363momnLctlzpC0ObMyxgWkKm9AOqfUkSD8AkBISGsTeOv9e3nG
+zDgBK8LYMhhtVG4M1kySrcA7EwdbG6l20FA8alVAXQskVLZNVjWIY6WHCn9Uq9/LcY7Tk86wzP0
dR35Z1wRJ9Ldp4FyzQ6mwigSUZUsGEkF0CYhtHT4g9Y070ApXFzMdklSq4XW4w4djF/kMB1IELFe
jSYIDQ9sPCOJ+3qQ+8qkBOGYm6iZ56wr1Gv8COz+J5wiU8frhU/vwG6q3kdJ7WEjOU2RgqetuP3C
4TcP+r9wW6il2LEQQo3ZxJkWn86+BKA+UaFdMCnu4lZRWx0bIlB9GLMadQ/1DYyoyQf5VV5kh4ml
guC3WHVW6zIqr1uusX0u3dHt5YGnLqlPBHO71xtoQk1bjQ/f9bo+5mIdlquN+1I+t5HpUZ3aazfM
rQbz/AUjyZ865o+LW2g9uFRv4xc3LdzZEamEY38MWsGzQ5xc7+xM7BBe6FTSu9wsjeWVM0SOgwXm
haYjFKrq4W4U8dhaOVIIzsB2Lot2QTTvrOflGkFvxtuIP4i9EC3676Wo6YHu1PC6HaJy9P3/X05+
sfv1r5UR+xkui9IFPK/lGHFFij+Zmf3YiTQoqss2obdUDfOCPu1a7uL7WHjFTUQKVEjyC4wS/qnL
ERuCFd8fRX0uhRI3orba98HajBOgvmKO6fBawpdt/nHeMRyXHnN5P991MdbyOrOiZ8FOyASrmOVZ
8UIT35VzPdKh10u8IXU9k+C4Hkr0w1sbdoBqzDSTGaQjpmUATJrK7+FoyZiDcfXTLZsVgpAwXhUr
GLs0TSkl1XRVp2GvT0ESH4uOElo3JO6e8TJRQ8FsQyN7bS7AHDK9a+9yMXNMGfQLdGZ2bABcRy4z
jlDyv+v4Q85iEDtujXSM91fZYPH/JkOnzIkc2WAjWDpjl4YEHxWB/obDU09axhYvAY80Jl50dnW5
KeD1NsOUlv9+ZoUy3aFwl+TOkIWV+Blq/gAMy6RZZ4PK2bg6a2TBLo8fkps7VLYZbKX+uZnT3q1f
1Nm+cfxiBFp4oMVrfrF2vEB04LUuhVQcwocA+1zr137Bv7PO8UAB+ai/xztZwycOrlIXzqUZOrOl
LJvtKCLc7C8/3AM5B3ZlpIpAo0HgcT4/IsWBtZatE7G7GzbGG/wsXaZ/J2VSkvLY1rL/v88AF6/1
Px7dc3H+7eFzGinCgqJPlaEUEfqC/lag3f5h1obAyhixLGKD6t4PNGvp7YBUgSbGI0+TNMhvZ38/
6cvb+XFNQ4Y66931cm4OqfTmIBrR6WFO8UoB0zSUXT8q05bG9mTC9szif0XBmkXIVVAXDmvtQGQf
egXfi0MZ2BVv3Fa5YerzTk2vgr9FFufXLwxt5+GHwVMApuH/ROM/zk4RZT5ZPWFs8Hpfoy7qA9Tj
SPzzryNVgCfoh3f0lJpRpgxIreHFJjBJZG1Srop4iF0drrbwpa2fZ2odXCIgIacLPYTUBEiyXU2x
ErEWEvNMu+Me87qSHMMlc4jGtsJRGDLyD7PtuRFO9akYHgS7qCkcsFDn3riVZ1m5+C9c8bACXcyH
gKLL3WknxD5fahMb69vw0OiY1VDx8drKzDwtgdJOPKFtREbH1rfK5fKX51PacW6nvN03C2vZ0O90
+wS5CyEU0dB5rZeVaFCgyqBzvTMQLdeTeQ8DY2y1ruaItnDG8YaVmbM55cEPB0dDOsxTkJ+bMcb/
g3MHqOTxi4iAMVhF0AcCEa1SWri9QCVrmJvVZ0fr8d5EAtS36XO5n9nfePiBTkQKnbkwHR2faiTN
QL2j9yP1pJuJhNP6QLjUni5Yz9w/FW9X/bpdD+g5xbHmuK/THXNN0okoJ88AEK4m5g5J3VZaptdD
qvdyDdpZCiKvftFZNUR7LeOlwnUxIbsR6n5fQ7kAkLhbCPm6TSPAtQQnHRTIwVfZZFL/mGKvGwkP
I689uuIHaeQbfZlMO6r3nhRcjWA763JIsUHV/xRZ2/6fqzO8udf/uOV1wFN/ATQgWbQ9EAwg6zfn
hhzXnkQ/18rTHZ2LWdA4urFM/7AKrzgkvPyR9Z9vTwJsRf/kDfGGOxJ7Ffm1mbm2HwWxEZXYpMsn
+HJmCPqMST8r00/5SwvwSJIZJ7ETREEvMyAGAbq+sB645tp0A4yz66dj3Eh6UuN9trwShSnWlD2Z
t1L1wu2LuIEEn5L98sTKwWaDEMiEAl1L3tPythkoe+MlkuteZKO84+w22QQUpb+OAtwMadqlY6Lg
clX3jObJjBS1mrrHtiEPXxT9Q4TZiqqd7SBiox4f73iJRL26QMPIW1k3dFl+j8fYIFdsNlyevg35
BWGM9E44Bfs6tNUaxAP6NGVtKTbh8JKVkb6VbYl7TdlPXeLjbIoLlaq1WMlBSQ6iVDmm7xVsKGtO
NgSfbwIQiuw+ffRETCPbBLeG3fLl0GJOZYaglOY8Fjf/Afq4vv6KZry2zi4N5oERl28+HRLCVqOu
yhUp/S4AZG6g1H28mIXptZrEKSksJ+Vh5vLXMyLEzolpkMZCPbluLsHfMSh9wYF3Ea/6tbXpjDIO
NK+9+gUchNd027lamyTBIT48NfcW62tjI/kQJl+quEkDBqAO3yMplPqui10hsM2fYFOxNqHlRTqh
7pJOwXOu4ls9wn1PwwHHcruq2pq0umZ0sbczoV9croNdid7dIXnWImCb4yTM9IREmIszmbsjJz5n
n/5sAmgS34hkeuRHi3V7/lNC+gE5KVi4a+KNN2zAja6L/HaI6uJtuSiOyQfnsJTYp5bkMfIijc4q
g4GnduoGsGkiu3pmAxo0aU3389bWFr0OySTTyzbjirTbCQDDOGAlfqaJ1bXxRg7s2F6KS4mo0bdo
8p46rMXM2PCnb2dE2N51H1e1ms4olCM0ojZjQ+dxzfg3c3v4dDK6qDMmVk5mwRmVQzdEdHvavKcS
7N8KhrqnWV3bQgQrqwc9NgqeIw1GCKQFXLLgOI+pDqYd2Kq4uowHQkL/taRAmkIv3l/XRXUC8bYA
Uglh8rWCnyVR2FjlKgR58nWuAcPUodz0HFfcNyhtjihpJ0SxbAw+tRDmb5g2rKTpTcQzOjOkCvA9
OT5NB54ixduvOo71YRVSMTtsJjG870ew2/sla3S8mN/N/KxFk8HYbUu+2yfVVNwTT39weLS+Jj3+
F+ny1YMu3O+McqrEB9FLhQTA6Ne0KTmQkRY+DCDil3FlvsbbyRa6nFThMXgi690HYglVvqD6IU9K
tKE0pPa1MNX/LpjIkXcJlJHUz8VnrjhF2Z7gFt6G1YhIpykKCjpE9dxbHNxJGRg+F9XROHpb040J
5NwiPoVM/W3SxN6Dhz90OUiJJpuPP41lncqIGoDT+TJAaeALUJy54uEpF/1lgJtuSGU82YBoc2ET
TlteBhWXuTrQp9ek/4hket4HN92DiQjMn12WxjcUovaD5jBY7dbpuPT4pxqgVy5jcMJYuySN2K3k
xo3I0Z5zu/eHrbSOesKWT9AeBd3FqYI+6kAaUZn6rWkcOO1+f1ID/M6Corc7zSA/4c1s2WywwNj2
ucf7LgJ+oXpCwJHQ2ul1Xi33ivtC+OzPUmcpibHBguh5g++N5u1ZYONuw9Xq8p5K/iRG+iq46vDk
CULsC0y/0LZCIdqD9BIUGHRfmohgCtJH64jOjFiA537cvCIg5s9t2WT1f5pSoVKwO6+1vi/4hX0h
RxBThdW6+Lbm/W/YP/f2JcWNKAFlHcy2UCUxJWG8WAqzD9dmpc6hsXCV4fdO1O7QtKCs0qOzh4XL
yzK5YwYUXENi7JmOlk4Da9agUwVh9ef12+6zBt/OqVnT0jNjSzVOPDywXtrVIGF57IzfUjaoP/T2
iaTdN3xgUkMmCg3kpz9OQ0hTsb9GDkg/csrkCkAmR+GriEKKNNCyiyH15uKZxgNpCgzkVir6p7wR
xmRBbvLRep8gh23FnqFdjwmCcZF1lxC/fgBJLBNz2bQhPm+p5CH35+oDLURulScKjiYmv7Ho6HuR
mL3NCI5I11+1N2jMng0dOLR46SzcBgD+b4/bwKurBfPfZT/VDgOrDtmG1SbeJu21fW728g6GZP5s
t/DY3JH3hO12V7wP0Jqf0ilNHeDN8G/NywBhZZ+Eh655VkNG0kNAL3wK6BaPco4plzFxYEVuNRgC
jEO7Q3RIEJC/wtHQ4rV90Y1TRxqE2dCJ8UzAc/6Ozjd9k/3QMuVxUgo/px0tgc8dJ/+XQS1qAlLA
BfaJ6khyNauDdm6Kmw+fbPMbTpEJb5b9f1njWZ8oLQyrQ9jfmqZFuS06YvEsBwa1U3+SOP/yAlDE
BUWzXRUereTVbfkZNECSHx0Q6Tg2L6/ZF/ANpQ1IlCCHR2aFoypsXPD5BhaE22enDYP5QLKC9o+q
d8JVbMk9M7c6ORzUAUGfs3ZanmFB1knmHOXpHLCc9lqWdLndmjAj3IEqBCdVzkElueEaB5xCdtpI
nODFP1U0r/Xk5MoYotBn82raRdkTiycczrNFYwx4iR9uyw1tF8n+gps4jwsfVmdDv6ojeiveUUJX
wbF6Rn4eBnUSHkRddOu85Hw5kPYMnZaiqhAbUvHVLm/uVOvmkarXMOaaiDMZC84wqcPHjKqeoOlL
mIqL4qe38tFDuYwmqnhfswnYRX5stJ15dTW8wEy2xMHku1HupgLv0++y6kEZBhgGg9Zorr07tuEi
TPTn3hEFMKBF9wj0ZX2x0jtz5NVvbbLMStEmOUHERCm+4QB+2ljsda+oAPiczJfYcAlrc69h4Om/
02oMQWOOjrSqnKgt5jp8dfPJcremEAHYG+NXeVGkQMJ/URaOsBaco8R5Bcy4zQdb2dkisqLc5Wcp
xUvNptGBR1mZF7Kjwsux69UujgYgdBA/Q7FKas0RxDpcQTGsnZH9gblLG9B3KYG/rgdSBoOrY8fu
d4BcfgkS2NR3MTc4h35O0D/+OM6x5aRmi8A+Nm0h2DOv36A5Q56bnH69tWe8T/qTyh2PkCfd5bCg
ZMKXxFSCoSQtkjPqNdJK2aPFwflyxKUpJkekR4sWip1yDH0XvFKgHaOtlvZ4nysCxAMw4l52/Jae
m+VS7WVDuG/YILNxQ/LhWm1ewdic6d8ILcdpSA23L6OFJpkXibavKmCL07u6gh1DSjzwqff2/DGT
PsguTo3NSHVMMSfBxLzNyxJ8Sq/weu2nER/BOrJ8eP6EjsF/bWHqjFg5VB9qD5DgZ/mlJQYzuNMW
Ukpc3pm4NUq4dLPiBaQSr1sEal/qT3kBDwOvJjuTI9OuQMzN4KvHknZ76JwzzPg5dpoLkpZvq/Ka
GVNmCO1NZm/iEn7HeHprfmu00UR6x+FPBFYT3l9zh3NBgCIeZa9h9G/4efHWlIIjCkShgRKOo5Ty
yhwMUIQYuvwbVyjpgEC1CN/tUkc2ox7aa7jvfOgdXLl/PXfnT1lGOCOSjC6U7bFagrNlQphqMlah
xbPlrVsof24r+FqIhhXhd/TMpWox506tdKq+zNb8clTTopXzODq6GEJ/hK8qqSHlhE2FkKKfXDZa
PUZXqVlg3OxTn/9GKLSsAcuBpKolZZKdfWO5ztoYGlTQp+zTh3nzPg8crDQTrgvdsjOjBbwRCNXb
yS2aBqtoWHnsxHBlAuoz/ifZIOFyEiWRY+N9oQaEOFDuZ7Ykv6WtZWVTxDx2lE0fWnVvLYgcn9LS
zg/cAHITXMBR5Ofp0QfrJLMUYZrLtAZ0IruXaEP8HevPwhEnU7VojBXlh5LPa26Qcobuk0Su+PCN
9hGsMX9mhZ6Q1tdd4G73dfJTrsU2w49qx52Lc3SGJvx8nLF4jenZXLvavYc96ySSU1rvxQRg4Q0W
aCDTCotoItnNW+qTDWycR1iJescKY7JcvnggOhsngWp3B50Q1M1KOlQIOu+Un4cCPyAADcZ7KxAz
H4hsvQtqXAD+xHfXZzu/M75c9JRn5TGvJ1ToeCmXtYLvBuSL/R3Fi09L4A3UvsnaAOGisP7a8EBH
LUedRGj34KZBLDxRUqqlckkP6d9cRpExvM9/xAHolSX7nGNwTIGKW18QmL+NoW3wpW7OAF8UGKGv
9wvRhGCo/A8WCqI8AokO9cxZ9WFSl17FfHwbFK8n24XCtEccenspDh9W+36louLd4USXSFnf9hnq
SOD5uu0Q3liYNKeDMRL/rUCS5Zs0nlwcCZ/qroMkYp/PABrkBhI2s+M6Y2ubC+0s2CTdVIRWCNML
dLF11jtGY4NLWiBuNUHk+0Q5cx9gVAJlsi2CAGgUDtEcArWyO182qzK66RXNTiZIAowJoIWLtjcl
PUp+vu+Kn1ssSuqBp6GfQ/3k1lwSjkBATQ0PYp02mjH0FvFb4s9o1NEfwQtfiWYNvSU5Fx6BYMSj
w+YeBb3tnbbDjB/15fKWZkCfmzcsyMIqp6339FM9xxjW/g5HE92kCOVuQPVszuGN2qvkFZxx1uxH
gU2QS4uywHpiKJMpnSxJApp6zTAcgQyRCNChKNxgKVwjNhVdGyDpeaaTBRzSxcgokjY9aKkrI4TL
Jp5Rhm48E39hYAVSUgFdZsv0Gkmj3R2ibofTEJrBWBmXOE8b4q+zzTUKgCfDaa/4CcJPgGvbqBPa
sKMy4JJQUG4j/BaOrKgengn8j1Jic+Jj98MKY3EY4iisOYxcp0zAJnXGcI4pizlFPxlwgwVKQIuW
iRBT49bQcnSn/UQ5TomS/fhYyK6qIIHk+0hjTIWkY9twrzHJJ8AW5ApwMqmv5XHiyUOk2xyS0ib5
jrRo9cy3wKvonMOyXUsncI+X2rQ8XgToBKebfBs6g20B0CM4bSXzxCR1rmlBc5hveEYbEfQf79J4
T02CwmPutJwx42x4s/OdeVv5hM/KKzJzacNzYNRGm9YkKTFO1bN5KhrT4cwZAx62LVtNG+yCLNDT
mwbKSAFL1btIxpcmOCCPzRU4mT9v/oInlaNfPvD++iVJfvA/Q5YAqOdWX5EDjs4wgO2zWdogX0R3
vCCWnIGfOE2teFHV/cAZziH+glWCS557K6IZEQDTn31q0fYyBsLQO1OCVW03ybfXpDfr8urk/sbV
fH4973SDyooLZXd6eNiXIcRtZri8m8i24mKKF7Z9yBLrXmAgTzUagmTW/NO6CCpgnSNIJwxosods
NztUfQtpeDIxu/OfQEhqnCtrhJ/OkwNiCQ1sJ/KYOSkubv91qIRXJCMgZSqFNNEzNzXgWVRpUH1A
P1E8pp0by0vKmouvL4HBBIBlpDPO2Jg/fiHucqpv2tebP+JRl5EUS1KdrDKQH0eseyd4MRSRXQ4e
BOZoxE8Oghgdn+nQ5PpcjNkUEW6aoy92B0oM/lnIZ7TEvneXsxeLEjEM5YzSoExx3DXwCuWc0dVF
PnivHkKkdbH2HzgpOLWBWRXE/F0qLdj7QF7GDRnoB9cjMC41cOljjNZ4ySa1+MgyFAhiQ/o/MRjw
e7lqQcCWGY8wJdS5G3JDdaJnSMc3HCzUJjtOr/a6X3rO7hBjjBJFs8L+7XS+ltvz4QofHDrWzQvj
/6n2p0tj4xumRYyiMEWzIZLcjr2YL5DS+Dm2J8yOo0gHabPO/qXOvveUrJr6ZCMVfgXEG1YkT4jd
Hy728iaesRn64ti4QZwHCpKmhkoVXwEf/VYYuiNgCjslJ7o0VrYQxQncqtDdxnDBIwv9FEfiuXNW
lCIrl83zkh+C7RW7n2qLSpFQZS5JDgD0qeEpZELxIqc/zErbob4j1AVCTVf9Vn54MZ00uNvPcKmu
hq/oAvbFEJ8NJlYjGQoDYkwW1xanQdmj3IKBV+U/HnGFWcI+G8eAQcLdDnc8B0ALEcRv3UGdXoA9
XZWMTTUrTKFgom+RFhQaBxX9ttU0sqvfeGvNAxaEDbeXycpf3fL+39iaElvcUARRVhprJLcYPiBy
GI16dhaHFr0S6KyUHYeLObEJPAnOmpOn9YbNgFb09QJMGxtJSgZBVCozl1m122i3r4E8h4ioMIIw
GVIYz4Jw0Yfq86fg/92mdTnHbUJVeX5+WBz3prNC89tqSN53EOsa3rnwVyrNFPkfOtrLKkEDwxRu
UaAX+zSi+cLbsKloB+ZpuVRt3DmUz1MlbMaqsUCsxbED65Ra3ucPpp67dwsfZ/Jp6wuHfbEE/yC8
A2yGxBISnrJb3CuRLY8B32XYtxto2jcWwFdvY9olH4CXXaItA3cH93wbeag+ujStf/E+p+Kyomxh
GpHMt62wfWdN5tLoRA7jtuiiaoBZ+xVFW1e73CYigYFqFKV2qxtEKdhdLkQxS1XKP7x+HFtxh4yU
Ky2W80Ei8/WItbziE/ZFCf4T+mylHWKPTWhFvRRhBn4fkCW0KXm9NVT8VdNeMkDPNyo8g+/oFljc
RhCwGK5G83t0Y6aTprKHRlklnsz8KrqTqx7qCeECdEAURLE0jrevF3ON+WGTaGV3hUAWnzr8RW0V
8sjZ/WvHjkCwiJ5MjFGAt1ANFRPinRJ9E4ZFjSfzpnaUhfh3Wr3op/5SWm1fpTZ6+AHw6dD/SfTJ
hcxbq8dAxTfhtiQSXnGwQwIVblvN+PyjeaX+/Lq71VjxDB6VwjWXtuvmdlVEbdPhk0mwqr13u/xq
ntu3n9UKCLHhPVfShPqlE7D/IBaAdukJXD9jnk28uXcv33yzU+s1hFuS9alFYwhKEaWiPghS+CN8
rHsFz0lS0bVviFXbyeN+czQP7D8+OmEiqyGhfvyZYbrh529+xx5a7yKqGTPTE+vWUIhudg88OI7u
wIw0Fuj8zzIpkrpRZdQk4hlq0cwWBkjUS6wWzI7BNnrpLErBxypFAnA1QZaeyXvLEpLYSzrG3iRO
TqBp8YY/zTMKikMLnXyhzuN7CGiUo2V04rabRAfjWKKBiRQzqivycorfnl14OiGLQxR4uIO9m0nH
eaSrOz1LCx17CWbZBn7L+8kMRa6prTvNK35vR3lznDbdve9oARSgOt7CUKaDqXRbsW7js2v702Of
H4KrWkQ1Gx7QP4/Z7VvY7mwHPxVJWXVW1SlrTW5Y145lX3ECwzbu4lwO9cBj4E8hg+bjCZKwhc/K
GPjQ7wdYqdScYv3srAm5NEIh0zK02DBedqEnS+d42ARlaw9xrNBqe9n4xxgTLxVKexAPeryaxhyf
MgC9vT8JwAsM5ug4t4LkQgekNhveUEn2wsK89Za30Llk0d80IrFhH3eM+J1bMOqFY6qdy2fxoprh
e2F2HkhM1G75lIxxIzMmklTJwODhCnLeXCzNa+DoF/ts3hI9YBbfhC8yk9+IvGTVJanrO+FJLxCd
IpoV/RddRAHczkx9vxFslejqGQ6wChoArNetDUvb1wqMPY4nXN6mu2etoMnQnybLlkTHSJP9V1mi
CAvACWZiYT2C+Zo8sPYxATtIrsXp3Spcz+keUI6HNySHm5jvUKk2peBeEcE7BGI+yHoOb3GY/XkB
ktQvz9oJ+msl6ywzukr0IC0QHhvN/zdFHfq3NER/+yvXCwACCbtG7wr7K8I8qlld0ggjE1NC2xfb
WjIm1Hht+GnzJbLPDXQZfWkMimI6SIz3Tu45dttcFwpyRNq1Fc5adksDS3vsTK9khBBOC4gUdBTI
KS8PnsThAPsp2exE4YhY/xIS2Bn4x4XLz6LDNMHjHOh8Ibg+npp5eURKRB7ugdqwfXq8DywBXqnk
xvXXi8JELlUdlqJ5roQpt0RxU2546icmLdGX20S1NVcc8PVQy2X25RFxHp8EvmEXDLMI5Z4YTtIb
DLa7DdJE88srKggsxLYusBf9m3WNoIksSbrXyz8YQb6QdntYyknZQarVYXoG2RloFv8k3bnwfycn
3TWvItmfpmwfPUO7sTOrSGRTIDxjExbFrbiB6rNy+EOAC2veokYW8CQ/zjaDiwUnXTQw4+707hbl
GTc721by0phtvsij4Gp3R+Y8zlv9dzlmwVLi8Xt/FzawjJsSNZWiBED7fSmYyhkgGccYR21unDDQ
l9Ojq7al1PK4QED6f3IQhEY7sJuyT9MUI0IqzzE7thbuhD0VYpcrdGx32oQ7QD2hCFesM4GdyWrD
+68Ncgs0TUZvnvT60d/I7mfuPohS9YYnOMirqHq4pX+Aa6vfc5QencjRLAMbDo9Sh1K0Vym7l4EW
xbwWgj8pOl8VE5fvNEERsL2os/dW0bdU5nnlwBbgyU7Y5OIGCL9HWg70eFtkFUhHmHf3dT87R/xC
KfzwJnusAcA/DKu/W83Z8S2dVYP6EvIw2f4RXnqnV9C4yznqRzQwrG0xdUSLFylNOliGAXbBmF6l
7MdmUk+wmiAfyhnYqgmd5Q5m3YepZCuUECD7NjkIkpzqBIpA/XcNifQlShNlbExJvR7VEGEDdsce
Vc+fsncQcs0GIS41HmYrR4Fw504L25n+MLq372RNxA1PmUSbZCioAdAldml0WQGL7cJIyLjRvd4O
2Liu8ohOol22DFbKlHeFTInr7u/e8zrVd7Yc7JN4cj5OlZcdgrv5UYXHAYHoUsKORRFFq3unhduR
xbXQH/fSIFLKYnM8PzQUhYpCHVX4+JLFZZLvPyfpdA9hAtm/i2Y5lpjLdg3RFA8FfQcZbV0mA+x5
QqlkDGTqUT2lJXKrSYNuiT2WAE+lBUO3bBud8LBCMpdsJfi36uiWSvVF0VznonQtOpgJuCwy2e/P
aNqVD1IOtiRv+6u+Rqw3iU1ecA6QwO2Em9k0seqmfWMNlCiaOlh1wYHdT3BLvhXYBJkYAtV+GzjZ
dRNN8hhKRQHpyJDarzZVdR7V1hJSqOxPCcnAb+3tU0kcAJdjjsG8iSbDslwp9fg63Tugs8GgGCFe
aTkrhY8xqRBf128+ufSn3XOEuJn3WKYdB/Ggw/weuzlaJ+x7/FMAXvKh18VaORmQlw4dKBjn35A8
PE0UvHUZguRAL+8SPlFt6PeH8foIfsetXraqDqQchTvFC3Qk71aSx1yfUSwJTJ+R08e7H+sCEhmQ
Kqh5RtfrVueEw4yyHP69nj/6JhEISblBHXnhvYYAvgg63fO2OsjE9dWvECCxV/FcxbGK73Ctwl4U
gMrshDg9DF+biZJXPCCVTY239O6xhmSIsxUaO31nkAQfsycE6Kw9ehUpahF+YmVKFDJKB9waZn+u
14AU/dlxVeM9Em14AULQMQHjBIZ48Wm0bPd+MkJac1VqkYCdFFk9tlObw2FWtDwWqSZi+Iu2awot
AkkuNgdELpxOfIkCwK6+YDijyEiIxTyAjIbxvYRzjOJfeQNXoH1+6AQ1ajgd0SAEe0dJZaTC2W3H
gOWbc5slMou2sMdIi2NYFNEgrO3y1LE7XSl8WuzUOh18Pizg3nEoyKXqpjxm99rOwAyGqVHh4JwR
GjjS6qOMDaCuK2ZmOZOoAQowKZ4opnC6ELUsVFWYeTHTL8eW9q4vTSLRd0CPAu90EkOLGJg7lTRF
F/VBJmnWJix9eOssYFRzOK4q5GRfmfKb6P6aGtekiVr3eZhCcai0ExYgoFIA+5p9q7cvidmkUMfe
hcoUfAJiSJNjCjcrlGEr2ZPc+Ru3/uWvo8V0iGp7MQRpUsYTwdIE7QAZWCMEPvSwi09smlvD16Cm
M8tzRxEDah4k4wEpTv6eu3xoTkI8QSILG2pM29fSyxGVQ040UfAHES/cNlKnJIAsnVPIh0Z/kJXD
3kuyjmoATfOrIAdBobCNnoKxPPX3w3ixug33jyYhFGjBn+D9r5V4wI/eUUoq0XzqKXPJ/n27xLpa
o1+HxBJX3Jpjm9FO9K+OBMafYSaob6HXfMKp29lcrk96jIbx5sGyyHKett3rOpoglt32yBqLz4vP
AAfvr1RsNNRm9W4V+hg7vl+qtVr78w3ZPZDloo8D8cUC0FBSCEyOHYfUyYVYPKAGCTkYtjZlBOHo
49mPpajyqujeX5zzsHJzP9TOJiywUE01jMsk5Eiu2v14Hq23UHhm4dGbAVRwMIGUcucneaaQgz38
cTDmSoQFpSS4X95smz7wvls+eNwp5BIkFtaYb1INLc01iyGOM9uoq65OSAjluYjImvNS4Wi4feL2
RbMyqRQaP9KjRE2FE5cfCgsGVTwhkZ85fITdZvxkLZ4gFZdNHElO52Rn/MFhKWp/IDVglv2ivhuB
0yNmVRGaAFCOk6sAnPk1Ll0WLdiC3UFovGVnkpQlUX9XBIC2Ty7OQ0ofV2m18F411EebHb3dYPTR
P9EJ1vMw5DBQ77i5ZuwcPWIiTUUCAhZhMGSaE2oTTL+fhVWj/2Qnwl46Bf1QLyEnzeA+DN0vuNNC
LDtvUT+Ot/92rOmO+6fdlfDh+NgTkqgWWS1NQQQjKr1Y9uM1jFNtnAaww1OC8HRw/u4x4NMQuJUD
xTKdIXCNYLxuUYFSUlevu2VwS31pNqzkOSOAioJiXHGqYPEPSJHjOeApKvIm+ikIGejOrRBrXOd2
kRPYqN1Dmu5qBmPh3zlMFynXNFaifuJxkQtsEXGZAnFmsGCtCwPE65hIQXS1Wqk1IIGBN4J+q2S5
kypq89YdejbRpyJKKf/p3XyRwrJdY8v09a4+tKat4s0V52e4a8oBmubj9VFilO/d1kqZabaNaaCD
cAtEh0DLEzMWJYcars5/8AtM/A59Ed1jDHYokEpiV6EPeA53vX2XJl4Z4lRMKObFus4D6NvIgqQI
rMnRuN/qTBP3Y/6JaBw4Jkm7Y96itegW5VZ2rzcou8ZI4S90zruuv7qZSEqpqo5IhGzmYpL74w0G
im5UNQ173dGi0/BmohbwqvOyJXThkeN+fk80FuLzkfU7bUjanAGKGCnXJ9w9kr6qF9cFGaEHmyTQ
O0HcNUM3dip+a0b41WoHPwwqs+NWuk6ExLF0hHvpqGzZpXpdsJtDJ8fuZRQWPgM+UcJzmqtk0mBR
iCr896gKrFQqLgzCoaiXhmsiYJF//kQjqj9X3GXD7nfTQyub8M/E5xs4hwAygdlZC+DZdn4XCXZU
SvpYmxUbRgfMBoJDtCo4Y9JC8yWYg2OS00iMsEXWpJWLsvAnRuVLkjUbMyr9oAgYZkvRmRemAJua
WovF2ITXo3rhsA1Vej53Mg2EJqowTIURY2tvJu9IxybdvkcXUJIsYTzagxoWANB9RuMpKeSz31Fd
JuJtttU4ME/1oveLtfvhB0I5OssB3EGMkrDnzNzjs66g9MMsa49pU5nPA4qqATzFTmR0oN/rkm90
8Kvqy9A+85qTYI1zSvo7B3TCeCjwX7gHbA416Aur3NjAUJPuVOF+W14qGSi2R26Rqdq+W33rof19
+8fQaI4URYkb7OPimG1ACMcMIzzYdljdkwaUDLwIk66LmYOS/CLbGC1pjLc60A15FMl51zi2tW7R
RJSvycCjebq1kDu4bk/zostjSBseiGyImLiIiIxbD21sYir619+VliSWgXyPr4rOYoPL991Qg9+p
e/I4KWfjERlWMav6/aCpATh86j8Y57puRrF0mc70TlluZYYRdu5ji8lC9avWBALAjBPVi1bTXxQi
vpW3zeUidM+oyonv/UYCxIlnERnh2RhnmdXQGo0nYlVldBox96wmd0UzkNdQFuJJpeGPi2+J/wRu
9Q+oimt2k9tmNfxNzfniYf4/Cnv/p7vLoVvt/CZCnNScMIMIeCWAZnb2jN+2TRUBDJwCp2ewnxdZ
scK68odBGf7gXdApLjFeFvutK6aK7gaoDvq4mpmffFrZauLkl6tQVXAiKW8Gunu1QvpB93dEUP1T
kqXUAL14bTBT8y2Ixt37t5VQeUS1zzWK0JnRI8BO3UbtWtomnZuxp3QhTZGB0znzRSHwH0QgH3bm
pNhszbCx9FytttCZuXRb9avFtgRDV6AsIFiAdZnSInN4Jv5UlZ7vlZ5OK37C3ffWC3pxXhvOUTNR
OvmSQpfa+v2i5x4VdpOP33KcN/sF8ZHHdUYB9axRTjX2GWf3RaOQrLIqBg0w6cK4V9Ugx73059g/
jb05nNeMx7richVn/2CrPhjjV8SI+1CHjoVjT72uAuSEimkJTwPuh8hMq26ikDw8nx7kvXUxRj66
myMnCEbfA08KfgNSqHgHDV85ML05OZMFqfD1xUHuRpNz4azWpLrJoq8QUqo/WwDzJVHbRpscUFFh
TitXv46/B6OL9PzVMafhLb/R4QbNThYEDBkyTwRpTHKLOmkZ7YFRWfFfffUL5s/5LI62lwC0OvjP
GwgohUcomgxkfh1SrboYP3Q2TmJoD3VHeVziAQWuKUySye//2sugttrqW8ma/MaD6gvRwLyouPN6
qRaOgkTuxTngrtMcu4GkTra40/sCdLnQvpNYFmIcbnLWUjuTDpN6yfyxfvH4sZZH/9aGjCg/+G+j
RmuLKYZ0QSRKEopj8swZjzgrvsyRIB76QJDVW4huWrWzJ+C4R9a1hwU/tLTKLYraO982JK0m5+Pi
J+XXMbf2y4A3Cc6cLImrtEA8INyVqviZaxVPU8HP/6YIc2JSlKznUMUnyiat+5yVWOAPsterDUAH
+4jW2L79oswWh7g0tuZZgxByi6Nhh/Xlaliy1ULn/jyZuJNAHAaQ1NVMlIRrIWYXXGWwnwN2Geca
dPfS8Ulb32UPOEatmW4xzV/JjwZ7FOxJsTBZ9dLGY0ga5wS++xazpP4EApFJfvuLS1JG6TjpEhhe
BYJ84mz+VwoylX9iy3FXJ/GOmBAdGXkudna2J1hVg2tW0HT7X8NYJTK6H2vzLQQsILdBccy57oas
luH2cTjTT9jKgLA1pqxL6DAxoUAsxQvfHBPxp2hfC1MesAMwE3waBJTLIwt1/mFz7sLDero1fcFb
8F7tZCfc29od+hTTRvvAxBDtRD/JVZoGd2MFWrjFS7fpF2hXiMAN0iKpzeTwFwXiwzUJF4V5FN3U
fCzqMCZoyri2t2VhOXT4WYxXjzegFtDuxesUi9cOMegzkNWU4vb3YdNzeG4mLKMO6y2CK47jytH5
wwAFirIeRJx0VNgdc+fhFjb6rfJHWYRAisIC2HCUzs23HcJ/HQAbMxZEKq6GzRZdpMMdvxCya4aQ
baM3KfgOzgjIBD+RVrmSa5lotZn1x5R+EvDwsBi5ji22yod6yBLsoa4PaO6V1XD0iZHR12P2suSM
cF0Ks2uJAdbH3wOL38pwIrat8Yh3WiFTQO8uDoZIeAhRctRPgkgZLHJFQsRF/W12Kx2/K/ecxF/J
+aZ48ur3PE6NCWm2/pkmL9zOVx2hbpiSyipEIEZ7D0LRyeluRHImyDbdEX2W0WYRUb8DLcwooQXF
ke1oJkm1ArcyJI1bNl/BEaAmYkT5+5+KnqZrsmxUpJwIdMhQfO/2sWO20GHaa52JfruhO0d9a3aa
llvB2YBa7cyhbpRT8NvEtKbafiz2ANzXGb6ZYMQq9eoGIWYh56CQ//e4RH7Lwkb8g+NY6mQI3rP9
E8KQbgUlLDHiTzLCwY92B1ltRBD64cr0NhCtBI+ojQbTbEs8M2j/mnytUGOivEZuc585la+gd0wE
p9Y/pUzWgGP3Sim/mi73iwiTFDPXklkpn27+TSh2eLegx+1ZsGL1/l8me3eU8o6dMQUptDJTGxYj
RGdsCNfsmNiRPgz2/BO3INqejJ4Psc+YHIIG1SBt7i5iAYnbyBzjYZRTs6JmRn8RzOtS/DziNmZy
TrfBrZny2qujfvQqt0PmUaGCH6G6RX+1zM7xh5dfn6Z8eNVHXgODde992oep9/s2qrKL1jNVU++s
q5eVGXmjfvajvKF0fEF014OY9Y1mup06CXnyRt/I7QH3/gIZsheb1zIMNmHXMNAp003yB2NzQbM8
XqMSllIG42KICMVyeB2bi9zb+j/lum+meFrvjt5LDt8d0TyvnAY78JTM/Zv1OTqNY57MO5GplgK1
Z8dQx91DROoV6ReKwTbBkG5Xugui9O90bA74bFCTociYWUZyv+at9cIx8o62M0W16XfMP68QVH3s
To8Ac1GtO87oRQ2Xiei3TYAjuqEW90EQjeyRYYPaRdSxkTdJENOg0LdD+vOQj8t22ffMmgvJIkYx
Um8vPxcEUuGlTOfv5njZHaQlOzqc2QF0pnsodVbezM5B4MPFW1/pT9FKUp4tho4JQ3aSpLkZg+hs
p5UMGmtWWmn0cCiaawhKlv6MVdeq4LUq11UuxwPDWyMIJvAxCdcDGqI04Rzz+suyiwL5g36Ca/u1
6+CR4vzjyvydd3HYuq7NuHjeE7Xp1OtNFZkzRddGyW5iH/qQVTi8aQlX5GkNN8dm/enHw1tEYdjD
gTc5h4ArbWDiD1piXW3x1E3R0DacsGhrC46fP3FGvxWS1p7f8SmmPSYwzxhYng8wPwVK43YRxwtG
Ct92m7/sWvLhP/ppO3OXkk7bBswMKeEG+4RG9a9hxur08loI5M3HyKmgROYCfoA3mxHJeBWp5z7F
XOXGJOs49paVKVtm75uVLHUuDESimdrit/t/Q37nJjjdzZtyTZn5sW6Sw81qPMf1UTBRGMJ2siG2
4K7gz0wz8kGz4Hb1uY4HxktUCx11j3lU7NYs2FTjs7TSNcR3BB9iOsczA+U7M6I9QdaXqaXWvM98
K+R1vR2TSmYPlOgWL/MbCzAzRofGDG9eBAxlO3fg24St8CV+DiazCOQngGbmeKqIJilhVX2wRSXt
nVVRVLx1Y0mX6GHKdu1TSRD+UH9XQYqrolNkvAWkTETtfkHOG+3tVb8pP5GSU7kUDrQwpYkbdzRS
YXF1R3Xrt8pzDvYUmh0XOskfRtXQLI90oxw5Y6fqiNi6GzySRbLsP/eN4ILMUr48BiHRpX8pJ5Cu
ViBpTvbSRjRlzmmMCGzPnA3veNCPKZs1qHAOBHdNhI2DksnJbcrtJ0YROnHJwtIWQaBxZXn88xvf
EsvH5HOoMvoZrsCFhdTUfR0pYjqcIu3/yTilZB2GYg87ue5LucGHD9mZgGxgyP8mYu+3qSojgfEk
ehlx0AT9KP/LKpXRNR2lOZqLJXAMGI3WzIJXc29jxVGdMK6CK04h/hXMxM+PgCKSAetUtw+lkrAt
akdVRQZ7Vs3iBCvp8S6WGvJzrEOlZyoHc5WEAnwFLX2BQVYZLTnfR5GIv757MRiCGLsX3lwKTDhB
BMCwApJvuLvxFjn93MP4bqwMgCdAH0vZonr4JjoaItYRlcybq9a8bjCs1MqJ1rYOzYuqi71fAgLW
/HEqWYTZgTKbYhFEXeNHM5dZRwEuhOJIoJpWDDmCv8LVdw5G8H8lmVLIDR/MVsgJIucxM6Tsvu4N
EBMCIVv44QB+e0I9jlNloFVHtmN9tUoAjhFCs6hhKbR/5J2WHKw6x6HXP8r1AanwTd41FQe/Amgt
J2pNKalJBfdHNUwI1ctB4r5g/BvSWmon27QtXPSxmoRLpYBIqizIxQiMKMTFbruL1q/t33oX4qyx
/zjB/y6be0C6uawpjssz7JgUK44BoVWj0nrbES6lvC+ytINehFvB9O+E/E1OAtwO7i7svp3JK8vi
uarIbDtpGQRrODgmC5tXce14DXFPM+gk2nOGz5qi17a42CKwLBavmU8LoredHNJUuuaSocvTwSlr
V8xg2PDguzRhuokVntigc5wM4R/hF1teW1XsU+kqgRCGQ9R0Gb3wo9MEMjNcRZbfeNIq6vLqe1KM
7uth6z7XIB4+IMjfmr3BOdc4GZfWSdebdf+fAF+S9c+hSqy50Z/l/ABBgcd+qGgcOjb4vHx9RfxF
KzeriNqRYeEMwbhXsldWeFP3g1DrZtS2BYOxSKdVm55FLd3RDC0BFSieyZtbkXU68K3b64pd+ZPk
EYRm8e8MAylKUMdC4TSmeIzUN2BxxX1h2bMtsBMxxrT0twoIQSz+OyrVEOp6LGEHAteb79cYg+Az
WXXZoXlcng6OpmP44ynXNV3r9+2qDAvksMxN0Vjjl8jAjkfEpAEGCNxj6M7rMG4BFz7JAUch/Lju
q12Ux1H6nRhHNdmTG1+W6lyONXcYiMk2nGONFhIEX3EWW2z4eHRCaX2p0h9707vG1utR87pQXHHR
eIUtevFlOlZ+ZE3fJez5jkLFD5mN3wvUxGG8x/yRU1X7Cc3Sve0NM3EQRaxXinHZ2NN8wgOyhX3k
uQ+K9sCotv/yQVgNDw/Y4A02HpCuLr7dDXTTgKD7vt0yPzepwjtH7Nmz6doL8SuA4z3wmbbWMoWc
S8pICM90tK23cCfTktv3pA0u0nYVgXK5Ln42FU+TOyiC99DR3PHg2CKjWJdmBJqG4/aZZo462rzy
ldaP6Dwt69qkhM8wNd/wqrV2hSAzQv1hdwPPwH6UEBtMPOOzS1HwuEu5ESqSZQjTpGjF4/g+4yU8
uSZwUpjkQnfJU1HXszEmxwJWeSzu6S5xzQwgVXTeJ6dRnLUGa8SMRHKcqsh1yGrqxL0p092enm40
luwEiXwryTcvRTF09PjgvHFshMs7kpYgAa7vFMjjz+sACo9PndHIJRq1q6ZFMksfmYoS0paAitMY
0DaRPC3JVW0WEOFHkZAtct11kNFEQ+MLvQaLqFKchdQUPFcJeeNjm4+TnuxSmm00Yit9ujDom5nm
gxtXaw7LPo/2bZs4jrU7L5zlPn0FhXLGoyjsKq+jrPA7VJoxHtba35WvNdHNYOd+YRhzoUHevv0b
rn/DYFgfj3/dgBsMuFvsCZe1yV54XwhXNQt6kKFp60uvcoHLm+8LTcEAKd+VnztK9CjGptnSON9C
64J/u13st9+DQ+q3U9jkO78NZltrSb4gatY2CLL8YSajf/Pqw80fwj0Oj2pIDiFN2GHkS89K48K6
yxv4/Gc071/UGUQHr/nycubNHr6fzOs1t8sKgpHg8ZSr++Cdsu2o/HRL7q4IJ8q7X41Zug8WUXHI
yxepjNgVoXGtmYSYi4cFpawDV6bbmRmbEGI3QlYpMSx2CY+ztV9HcTI199kA4Wl+K0q4bPT2gwgt
ky5RBAtwPZgDTNaD2DO5Tm3ShHw2hIzCanVumGzeDwd/5DMGVnvv5sSA0AM7JhirLhQe5oV1w7Vw
dP5hz4/YWlth2BrDIxuu+zCVyJofV6BbybzHKj96cUMfQhghh0O9kMr47fVEax7mmKsLld9zVxCj
iBodGRWVXML0Eip51zSrzsobq2W5XyYlzz1DfNqSdY9PennnxkKXdLXWL1vTlQyfHKxOHzemrgkG
tNT1lPcYcBYs1JVMixRSzkX/YY6tYANjMJ/MA9F9C3W4dHtbN3OArDIRu4drjpdzb/5kTchaXgXe
1h4vW6ld0AzTrdxphzSIzAWp0NKp55IUveQp4uz+hiGp5+3sm/Jmi8kr+nsRJlmmYPfjLnMaQtFP
fE63zl5AfwW+8L5kUJAc2k1srr4oi6UEoiu9j+YQj8HIyhG20qurQoW+upb9gbTfK/p1H2HGQdbE
8jbY5iGvi/jVGh9LFo9fTod0LbqduDu9WD7F2dyiv4veQmYpxaoTFeRNwKrQxAWib3ghfMsSwLPH
9DuSbQkLUaMRPwUxyNS3aNV2BAKX0Z+awkyOo2oY7SPjIFIHRFvuxrW5dROI34S1xm+uyHJDBuVp
GoetmQe7e6xC1L945VDeMWYcVdye45S3b97eVZyFA1I7K0HJ0F5dpPZ+Dv1lKs+TqMjtIfg1ZtAi
Dvp2p47RpnyDwucXr5tgpeUxF98k6y2FGtVfsc9+F/sXozfkeltiCfpcz++bvzNJ764+T73ikhJR
ry8OKDNEnvpPpJ0mQJc0C+KXCrX9kErTvXHUYZOjcKD5zYFQdgvG5iQsv+H8qAwWMbVtS3YrbiFO
tDzfWtI6+o8yqnbyAIKs2Xcy1vS4YSWfbS2A4HmgmRJ+BfQKSK2EW5FXWa0MtT0oCSA9EsWg4fiJ
PFZfTH8wZ+q/PwN2KH/lVZw7gtU5sgFd01cpbzCxTUpRJB+L795ARWH2pDyv8+nD5EnEYbFwQnNY
NYgTjB3wivkbbVxany2QL2AnZPASXBlyR8Qytc8dOmJgkub0vcYhSiG72CyxK0JFcT8lC7T4rDpN
u2J1YKKTTdP21a6EUdKPJUA6LDOm+7tdSn+LS57eLl7uzsAMAouZQHrSZIBZR/mA09EwR33dM0Un
rCZrrnnrJ0FS4+rKrm+TvVwAWKo6W2hb1B/xmAs0vMZw8xMHHMlo18fJw2l7KQeKjcyrK0XxBnz/
O6cQlPwysP58bPb2gklzFRFnivjtJdjcIwOvY/LLc3lwgJaKJknA0vGJAqzMWgIwG8sI+GKklkH/
UpJuY1hjLgijI8buMgJKgNRbCEURLKoUTuSva24yzKsDvPdn25DJHOlJr5D49jwgjBsmZJWx3u4e
tBnR+w9fX+pEmcYfyLHbKw31KFF1Z7cXa9pTE0faBiNM6EXbxJKc9GMJdFBeqikxPNAFg9zrwC0Y
DFrTTI0gVn9GVhGLcv8iePQNoAY4XZ+yLJ55tJdKGbZj92qpb/jCHY2AZOpMdJiE/32H6AEsyfVi
B7hVYucBjWqacafueWeyCbiN0ZRQKKzwr83LGRjaAV1QiAVCv8l9UM8ooW0K0Hg4j8XXxjFL44gm
XwsW/QQrCoLTrP4lEM6KoEuSqClEGHnDvfBBRZnNmpcaZXAP3lkc4xi1f/yObyAp8w3+uaHs66nx
gc+ZUGZEHH7gYNtu1mLjL96bo9e4l7WRDSVVeXGXOBL0XFkFRBg0/SASQ2B7GzekYGsJCGmkXuaB
8oNY1kkS9skdkBMY7m8Mcz6xi80giHDg86X5iac6uvr79XAOy6uxFWa5nFPjknkQ8mr+MqpvXWxz
60nw5hbEmhkjnpyIK7v5bG1DKde66pABXSPoB5ef9VKczTQLglUq8R1taRqvOqK0kLWm92PvWTpt
uF0ViFcOLNRKAac4uBPTFch1r9uboQqeUfE2pfbtHruHfKqyLB5KKhzEUd+Y6jF2Aju49fu7NW/w
/sV+nq4k3cPRLR2DKHD6xJ/XaT2myr2YVbHYWT9Ykapq3v3aMwNdlZQ5JhT24/vUj4FCgPIZ91Oa
MxDWJykk0L3oKlqFeCFo/McBOZEWZsrGcvjLBF/OsrMVAZFt/tIr3aeIAH01I1lzmw1FtaIuZlt1
Omg0MQRl83q6QZa4JCMQUeMQ4UxjjtuFFuIdRDxwHsWw1iksLAagjm3HkUHoyD2J5HqilulJo1Nb
EqISetVQ0SvAxqzpKe2xOdEk+bR/Uxd+n9oK2XOrxHsBGfcExJ1AkXdX6+oGSwo2mnCroLhg/Rmc
trXNPWdnBss8AxBGPuBVbXyHDIM4q0s53uezqJ5MprRIeSNG2cAe5JXKMY4qGa7GbDd9we5ti5VD
Q2cwIfD3aT/2QrL2JaNgBtO+XXBwGOomc4vu8WTjsA93Qr3op+NsNh+UrziU7Klbozqqd41J1H15
Kx58+BKPVnXcYZnxWdAZ1l+9sSmKM6XawVyYFS2YCDhg9LJRSGS/pm4Is2iZk7OMlUg+hx49DwtL
8Pm3yM4nAGCnJuc5UDB8kN+v8YSgM37/Cg9mW6uLAKqv1mJ8evN/LDoEv8LyX9D+Az1XWDRvpYe8
eCIcF+3COo1nnefdg52as3/h34HeNQIKitdSb/fTkaA5gky2ste/JYz76KtAOhQlvbV+XdfLzgZP
y7cR7jjxNArR4hxN920GY71nbPIoLmADq9McU9Sg2AkNDXY4sd0yeUSdC1frMLTA7yfJ4XZotkO5
p+OyN6czt8IWtTKaEod3FjrHGTvDyZqgFbNh6DUDW94uRgiy4qInTug0GR3cZKlbIrz49Q8V5Nxi
Sh+C7oRmbs+RzFpiXP5mGTijVBls6hfAEvNS+AVgpYqeT6LndNptAFyIZkIsUM1isQdtHFnhS4mF
jmxxKmTYRDKlA2w1mna0MZ/dGtJuSt9zyP8fMOyd2WTLUmE2XQ49ochzSLIrXFoG5SZMV3J5GNtt
QkGTrkb/x0Rq6H3AhJJTQbxJYVcyHYaEUENURWdBzbu9Xp3pevWd6k5oKy+rhLoKLMLTbq35TWSG
oCcQRfRsn1P0aFIehjeRXNsiGtw53omoEjW3IgqqW0NJud4ljTLcgXfWPy7J6uqjDae/5z295A2M
J9e7jr+MtCEW6oFaYF23qHnbsGyPoKsmo9ujPFqtyhlXP8NS5WTQD+yICvZM9Rw2U3eQ+F5Av4SW
P3K+3gYUhHyse3A8y/93Ps144+4MfsUywG7/MQW8QS2ZPJPfQ5Zh85vqYKJipbQAnJtacDWRR+UO
tHw2ChCf8IJ/UaviMj6Sm6ewxPlTq3gZUrC6EwHoP6KTtF1zH7XdwxqHWZ20aknW6TwQyrMx018D
CDFc1//ooKRLhYs0pibyef9bfeBiEp1lYDBMIAOU/B9Se0Gzxz6o/vTSl/hPVE9nzFYIS6n43XsM
A54R9BV/Xi0lT2LM+NwR7gHevnOA2zzUtCPkt89h82ePrxpBOGghQszl8dEtDbaP7v7FlPnyl6nR
MuqNBdHXdYWLjHEIHpXZNZIDP1pf+EjHs4WnMux7nGnAQEVFtjT4dMUGxVOFy/YqSqzspNuFr4HT
avF52TuxJSsMMDh/uKmNOL/pV2JJ5vXPodQAZ+aBJb4bcAhhwrXTXnSS8Q/nrXSaFiLTeicZVoEB
x0m8aotDTBJiE6Or31jdWPhLW3jyzyStAhQz/vbc/BnPzJ6d8kFCMKTVAPVTAZHMFH8xrm/hPIUc
5005l56sS24F2W0R0H7SXrLaDO9qCwvlzmz5Vg5I9Cw9QPd8g6UlFPVGW5LcaMhHnoOC/G6rp7y3
KaVrd2G/XLqxVJUMDm3F76dAbbnzZKL0b8zLfi2uZudsC7GIn7HmeYjqVjNq1Zja7XHNIVVzrQYR
G6Ynr6MqT/LN6vIqL8kVWyf7FJ9ovW9h2DjrKdqT8NjpKf2EpZ6hvoI5LSTbfhPRQcMWRYs1NiFm
S4QMo+SOB/PZnrBpQbErs48gBQkzovZZij3jPWUalHIUHaJSXuTAPSvpC+BItXz3QlgE1O0Mzs2N
u9T42f4XO+zv3PHmbXVAc2ydjvWY39QI/Ol51VSGQvPMdF5VPQi5p4blhlZg0Y5AxFgvZFn9BBtX
ysN5mI2VTrMwDGQCytyp219FZSPWG3u1tzm44vuOa7ed71Na+ZpYYVyRy+RXUE4Ou1TlyAkzBKrF
dkB6nrZXCq8x1dTfaOgp07JKk4ygT0UkFS/7RIXN1aVditoK6n90p3iWCqxT6m12yNELATj0+LL+
1MkV+WPedlaAkwsvkYlLEiVJnl7uQahPyG2bkj5Q3Ti3QU26XjZ078QGcJyv0DaOBnFB5GTsZC+B
+E8CqMvfzHm5iyoP0SpzeTBixpOuRzhWfLRW51xuLiBV3OyDcONRvNKq+SMN1Z1ccF/o8q3MPbVp
NUmKNr059j9yf9sJA9kc0dOsnWTpp5FrI68d+YJzY1jHN4ZBZ6SmNoyBH8Q5PO1pnr5JkTbKZ3lA
6kM8/KpL/cZY3+wVhMoiXXKdrOppPvbMWWJauP3nYJQ016R4ovhlEjbzaJGpOVPUn6n1SSDbT13a
vIL35xEmvAvEclh5k/DY2Hq0ZmN3tglwA8Hg7VgQzfNZcjhAEReJMuMldJyvINIQCnwijh/332Mr
DaiQ+nSnHlVs1HT7cq8FczV1sGPUmP5pj37hwzAFwP4lCt287Q7VCLVsh1lCLFw310qJKL5Jxu3e
8XU/kCksJJfCPdX6Ck8xz93AQiWSfaxV6bxuXGPP7TF2bjzpd50VN2JKkaH2FM82RPSzgEbERquT
C6FimI1gVCl7v/RWQfosuFy6Ow1Uv4qokMnaqLJVy8cdP+TUxRtLl89+GNL1QwHY75JDX2P1JZcG
4p29afVdpynNo3pRZdG1XZqV94jlojlsqleXnuQ07CGsES1uMCp3uYbHSkXykMWx2xZebfaNT9cR
4gX8FvnIP4LljLIeBYwvbc3i6IRYfTNy3udtCOG4XQsWJbnEnz22+z5Q5ZxtKV4f6TnPQQiN+snF
a8EAVe9W4sDDRs660OqBWf0rpqtcXYje+918eLx+flKD6I0wj6P02FFbjQ5jDwXPJwfO0AE2E9y/
qikP5igOc+kPzkS9UgF3oD6sfCasSfwc9Judr6goOwVFlHA+1g8otzkdAXLTzrC8DiR/XuHQSfM3
/1pRQ3KncBlLvrDFZE6vyKs4MjDYOZpboEKxxh5ytrEQspPNd44fwjx0I/BZNAHWfjrzB8wNsL7J
RTcwJgLkGhF/GWpu05X3vGIizZfJZog07lqZV2X7XaJtsJ97WVH6xWoy+EyOD9hnkS1Wxr9rx9AA
jLQh57yWWl3XioeIkJXZ2vy/8R1/At3FZGF4KNRAWMio5QaQs2HDLaj9JT5JnljjqiK4Z/6zIWdO
YYLyJjcl7HfLLdhVkfE8Af00QdB75Oabi87MPQgT8y5ciu6jTMMhRA+Muwa6tROmFY2LT9Zg7skb
sB4bdkZhv3xGrWOq6GBYwraTxHztRKxVfYtVTFoBdR0dCeLCwym/MFzX+plYqFugLtaQwaLF2Obp
RHHKjs3CyjSYuDm94rqxSI5VnsKBX1RLXsGbgOy6Aw1WJVd/Tl5MIsKYXH5hlgJyLVEsOo/SRlcN
04UVoTsK/+eRF+XJPIMyG8PJ8C05ZXB1gfV5xIQ7aebPsQEfUPPkjFyFR0uMcH3zMmI8iS889KI6
bx7maAe/O9BAGZNAyDmITX7BYTmhm/kHCyh3zpVcKlIm+K1LCgYKZS4+aonscE6V0raY+umoGuxe
gIHxkdCgC5Ios3ZlcAW/f00AJTEVLxmaO+Vu15dAWZRncFvPxZoz+EK12MMRyuE4gwVk8yKwZ3Ne
ys+G3UmEWtjScPa4msrePmV4GC2gsCKUgaG+GajdwXDl5mLHAn+7OfJ7lp1+iE9bYarSErY8pbmo
G0MzDlYD63Kb8EmN0lTkr3RoklI5jU0SanJD9v/EMGApWD+bHy38LULYgxJsLC93iY3GlkM9ftdA
vvd6d7TtOytCG/YIQcThOfZ6OgJ1pvXtNVwMPVkRmin7n5Mm0no6WboVpG6bjisL0gcTxLJQad8q
MJfOITNxhsnytiEurbRqAOiNqQjmqPppFL1p5ipRWsFTEVX1DJ3INUNb3bE2gxdFtlBM8SM6q7wB
nDAchm1fJmXw4Drv4svtDlJor5jsgfDC95wB1TcMMkIvRUBUFoZQCJCPzA2z0sQgFWe7rqzlePsI
LbJKLtqaYXn3JI9W/lrYNz7ZwAevGemwPkBg2lGduJfykR984suB4hqUbGY++O+OEp3NQ/sFMf84
Ya+c+YyqEYYHjCsXFMFQsCvEMBXVb34IpeuL4Nc2irxuzbCfA/Dh+QrhqynoKpCDx05fiN4pSv9Z
UHXvHMnxgq0GZd+taslEeFbn5xt8Ywf7meYnsTLsfitINL22LFgnWVacUloXrPGm1orLB2gUJeUv
Kgbu4XdvIoiGcST+GoCEqMbU3LSEYTxFP0tRuDKadfpKZm4yKZ+hpYgwzsXvSDJw8aA8zg7ME0i+
kI37iVT3KjA9woq0FRu+c1UJAz+9F56bbDTy0kh7A6IICOE3ga2NZxvjhoiG+e5pAh9obw5mkK1O
fhiV55+TutPzghwSVNbmCcXknaVFLHwxfb2RDSzy+X0vTCoWMvxIYiEzH6pNQg9Q0hoN226pKaGi
dWwOX/f1YK1BEYn6SHXNgLZ1fZgZ26LAGmQxyM7ceY2A0lyqVYWp4saSbbpINv7V34OC+P07gxO/
TT2Hd8lIH7TnTU9MWC1x/889YhXnqHlGeRzKCGfBltcmuSc27ZbNhQVH7sBETFgqzbM7/iSx85Pj
zFjmwBb66kKW3TA9Lopu1WyZM5K7VHTMxrlu5NKd106doWz4QpNL5j2yphoY58+45baXTUuQYxxI
lyPUfe3p5qu59vMX8qC3caXEmWpOMW3/h1u1HMnDlEtXNKKMJdgA27HF1XrMLC8K5k64LGlfp0Mp
yzUZTVGPKnePVgpNKBEObKCI4BrsMvKsfBQJW1bnvYrLp2azVrrflYwfNYo5WgG2NqfbgUvtYycG
mKfHpWYouvASdYf4wnJEbNFuZgvJBo847f92k2YfgxmteL48zIG9poEwj68wVjd9syPmxFrbbAmb
q6Ak7YcoTjdnueX8LbmHIPcFc49pdu+52cKu+6P7JndNWYqsoV3qFGuIpqK2fY0ikqoQ1Vbx/VSN
1EZ/FmskmVlmr3OlI8h2hwQhf/T8eqaJbJSSR67sb7TewrGpGb3so1ZhThrlA5qBTodO2ZlRwvvi
gCWFPKHaA+mtbLSJxFpVqna4gQs5KfWlVdZZErfaTAJL5cGG2kqd6QqfdXynIQFwMnnp26/YjPlt
syXXi+op5+wdopTHvE0ZeiB69XWYZCtyfbig2eg7Iyag0Tyv7mcFIRFGhvSTdJz+mgJZW2Y1cuR1
wfuir8Qt5ScMYFnIQiVUPpyveefzmAtZQLnwoenRuU4XQfrTsUuVvsqm/59HeS63AT9ur44meqb2
k3aGsEITurupTt+qk/bPd9NbgPmWZTEkCeVX4tT5zTy7b4GEN2Czc3ZGLmo/CKlgOU5oic6+MSfo
L4wFLIY0adsc2Cxsz/EJ6R9gXX9tYvSyjXv5QYIZdzlRzt55TPqYwqUqyBYKrd6if/d6f8bQWo6F
lvsfRUKhoUZHeMl4kVVYdu8QzEnKJiz4Swj71hNFPP5oj9wSLNpDJaorAH17YMDMGYYdzYmJ+eVg
+cU1pOUFPh4kQLZwJiAnBR1G9+8lNO++IpXhKLIBi8gJ54yfTuFRandAQ2inT+185pCIiSjbl12E
f0Ltcki0qReoxsKZ5ES22I06MBp2JhRjCyv2/lFnEKadvT4xAG13MBhkWBV8Iu95sl8+85AG2A5Z
d/l7vnJ8Cb0SmAhjpKH+WxXE3ARJpli1NQWGRx0EDLhfaonGVlu9AVLWBP6irdqrVhu4zZOitP0d
jANClXyPqcFqx3D1uyxeCK6A+7RRfqlbf85qvWvQ1uDN2Ac1fE80XI6r2wZSmopXV3NUzHF3gHpy
8fCI1iqi8hj+g0tGiaoG046BG1umw/JAFMpeNxPoyvzARVGGkfG1gDY8sYTz0LDrjLjRAxGyzygB
68hyJ8hu3iCrRMROTrFyXB7BzoEhkO6XmpVuumkTBuT4M7YRS3sg2gX5Jur3XPlbmJkCLR3Ja8BH
iqJDMMU5vzseTwsfzsSDGhu2hQlOnKmkLgyQvJV+Ic6tTrh+/zpb9660EeabyLd5X57NbPtKCHRN
PMkb565Af0Te38vR0Mm1PqLeziqJMyxz+r7OHGS36vRG8W6Vl7RFvFSS4e+mIbVlhLwWLN2eiPO6
3AsPjDLjFAkV+QYxMiNVBBlmQXO321OwIcKfAZeMq8egNk/S2CSk26VI2gER/7FaNzn82wp2DkWP
evR3LOvQdYtilTqcpF513OkCjPXYKepVelYlWSm48D0NVuAG2rCp7yDKEPMceDEfAUIq2jfPr70T
3/lkumjCWI1lS7GjItKwPDABjPQ1QrTshgAFYD8/POh3nC7LqH6zysKpqg+QoyBtCla8iueew4u9
EGXvCRed1W5CCru4yJv5Ke6onAeF0g2ZswaAyr+5PeqT/mVQ5i4sXvPewlj6hhXSMrqTrGw66XmB
RLrrbsIwRCMRGJw1RQBguLMUIfgNHI+yn56B39yVPtAgXbXm2UqqUvN5w6YyVaoxb0L5HCHYfcm5
fkOEdSZfUsSxURDOyNoMNwn+qnjj9JUqQdMFzwZJZKa14U8yiuIoDu5CLBngtJ4yD4PZiD+ABGHC
yjh4JoQ0VJHpWgdroTf+CJGc0Y9q7UajZKMiFLhlvVKCEl73S2joatbDXuoLZ7aXxX8i35gKXYjW
1c8R43BFnIx+91q5VVrz9Hq3W9oKdwqNgE0bjT1J27kCRuuWFxcehEc+xk7iOtXIjev+MMiqpxOB
WH7mLe1GDKvyZi7Dmp5wI/odhMvF5/gsfCtQEobcIIe4N8OXGD7rEOWTzg4DEFz4UQj1HN6BeSpj
NGTp0bJkv7fyYOdcP/rZ9I+xah/KV19vw5wM3YfI7TZfAJ86FuUPnVq89jJDFnbIBV3EN+GqwUZ2
Rmv9jYP8iZ4bjhznawQpd+ZGMYdRguACBTOXByN2zMXP4BFHAxykcuErdT63HbT7N1mJfsnLSPDn
LOMVhyqzabXTZj9oF64MIHB2gztbOEsqJBLwOqG0KJT9NsXGqxzRpLoClZTfgiEutHgU+8xOxyPe
dCunM63ISfgpe1sORSuPEJdr6AxTtjQk1Y9AY1/TAuThsQAm4FuhE/AyeOZ3Ctx5di8yIZnulCFT
lwVlKj4QpF/j8qjIe0qJ9L3BRA7bPcURErXQNzmeJSAFZKMEoi0cVcb3tLvnNIpjbw9y5Zczi4gt
i9lKn1a0PuvOjwn9imGUkoPWyCMXXKuLna8/Itd+cs5hIXYPOyqX7FkivLDt4XtuK0eD9ekmK+Pw
TO5gpcym4QDNWsqS+a+05ePLnUJ3OmZCX1iWp7XC1GgygOGMUvyqFB5yw+in5W9KA/Rebe3S02CY
8ECWd3HI1ACtFmF+HHP7MpFSNzAI3WmarJooYel0L6IjfPB1zA1cmkoJ70OwjrwL23WR93Axeto8
ydnwc0WLFJD5PQln8gcwCCg2GTR1a901rkFSU42BlGIAURR2DaCj8Hb0AaSwAhWumNnULpPsOgVK
xsDt3qzc99gUqZUblCWQBFcNnrLMReOrS6OGqq/uO/wqAqSt+hB6dSjaJwn7GU7GR6ZWH6IXdIXA
nPpH29LFDq1kqcWyFzjNol8xcVbM2XoOVP/lHvIoCnLcreILqqZZE0QrBINSitaC6zwUTqJm7A7f
9uouQIcAB08x4vZh+gPFVK9SpdpfByncJCZALZgbL5VP7SVXVB7yeuA5wqgs2HKDLpDLm96NatTL
emLQN2xzj5fhK4xfIGDY2zV6dTRgOrbaLh5X7uUVVggkMAa4dHi5d3GJAiwkJWPDkaoT5KGEEBWI
u4ac4PbzLA5GQPtc/AmUbGrD0l+6kY5KKSNOYJJ5ruP2+k8ySo7P/ZQ3ZL+NxuAff38ct3qDtBwQ
qfWzzBnd4ld+DU51iWt58u1vmcnQhZlvVJfGfSaMuMv/4sqZmFfWrSQY/5m5tECEczW6Qz21ZA6a
O9Eiz4Jg14jDc0H4VbAEU7aRWsCYgwCRZEQlQgBK56Y4Ft7l2HnpKzrgLYxS1spEoQQ4A9dSt7lT
7mqkq+EK5PMtHrRLxePeYbxIkdIjiZHdBcQ1/TB9LjorqwJ8OT4se08HQwGS5dVieOQpcI18El+8
PYSI7IVtCAXcfpBN/GwIinnHbIRkIowKJErdfG73uPMGQQMP5uQKePxe0coi0rzFIrQLYXPiND0C
c+wcfKdzlxHUtyLzfgSKMip2h/ughnSyT4Ylaspz04jIj3TfnMDl0lRXmw10QGBVcCHHOyy8aXRl
I3Uf+s+EOyGmc/0q9cJ9ELlKDic6gW9eAPTFJqnMJ3mmlgVlsPFzcAR7xpanLcegBYLK/4nvlvDc
hDsYkTWFinlO3dsgQ6uVzPWv3TGfDSaCvwyFwy1pHFRxUikx9P/qtw3rLjjHWGyJ50Ih6sbO+cPg
WN7VsmWBYZlqZZUrCAnJBX50UMvFmzpVTKaWzMr80TyC13dC4rqaZvk0T8ESBqK6NUrlzFKSAeCn
MobEo0SvLPMY626Yo9geIyVznrSam4j3u/zxGsrI7WQu1YDk1jI8fFgKnAu3HzCgfdSO0n/59r27
ie81nGOSkTqC4AzZsyf/fICIBWXla+kGD3VL5RBYns0eS0+RIfRFvPSzDBYCcI+scmHjsLbCRHk5
hs4ohJOgEiJLK6kAC9+X4Ko3/tqkFTNQrjaMXsfhx4N6LEXuBAmrT+dcEqN7LrBwE3h0OKFc93Ox
dHhuR4vdJCMctBnoTDyxjRykrE6QKHBr0erS9E+OmkcqLKHCbFBg+ZBs9TaCaJKhX5SJqeOV03V9
SjHBROKN4OBWjE4pqB/rsXZMbaN8mCEfb8DPwe8PauIQ9T2O6VoN2nUu6EhEoPAPlDhrY9tAiXQ3
+g4aTixVpMeNLvxWhAS6rK2kghSgYnuLZSihUL7gLm/tR/t5y5eTXf57sqronS0hptZBRm6WLnns
La2FuKZOorgCZkl9iMXPysRZEP/9kyXdHbbQjaXYKxVYRIqAAYit5VH/xOrVEpy3Te2nPyDY5XZd
+jwUmUVcDj7n5jLqzKJFjULkjB9A2RKOcNduR3MCqmb4+0W3FvgVNj3Qa8hCQheN+XEPHCRBFTVT
IZ8JY06eH+9+a2GsehQwkGCAhNUmIUQULVxYEMk8z/BxFgcnFuyUfRnryMPlEu3yZaLYiDzP5AWK
CrQ1CApIVRdf7nqBH+oL/UsaCDQ0bpf/pyab5hoyuE8dbCw5GZMrgO5gN/alDgQXfxxL/vnUkxWV
H/NRM7YcirNC9iRqLbnp2pXa36WbJV7dTyWnvJav1KKYh7z1wQxmzjEZ521RrDUOkBXgGpg7sPMR
nOp6c5GLfzbZuGCj1oBlfTbucj6OrKWoDbxqFGjdADvKfFC7C1fW9EDBGxr2XExgtYY2EWN02A6F
3kH9jW0zbfnJk/IrX+RTRGzzTQZQaeRWPwR+9NOYsNGyLWYf8iKLpoZHoiwKrDLFf66aIlP2ZeoU
JGZu1A3Giygtr2T2SHT/ruWLPi/iMkb6xvIUoaK5FzgRWkJCeVOMVFiajjkv+CtrIGLAvnNMi45K
38jJEVnAVwu4K1pQPXP1qQ36H4tt7C2JiiA90eUS7b+1RgwRAYbgNzc3cvQTXmGHO/GZXouvwQMf
uAh2pxpHWW9PXuRdBzSMrSAxhv6FuOkM9rKsv3VMPHWP0S6he7nu2QNf
`protect end_protected
