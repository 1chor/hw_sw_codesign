-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
XbKxEVnRj04qdXUQuqVmo6Ujpkb14Oht/sCUKLuNACRXBHn/c3PQ3VfUzWDjuioR
OK7T6F1O8hV6xRwCPsFAWjEJQ8ASeYaoTVz1i7lLuXzHmD29leNiSXDQjK6izI2k
MzpfIZ0vzkqCtrwzJ0xu/Lume1qR0RxJZwxXpioneb2Kt5wBDooUrg==
--pragma protect end_key_block
--pragma protect digest_block
zyRmsS04e7Uk4c4mZ2RL1QUMlL8=
--pragma protect end_digest_block
--pragma protect data_block
MlAeX3KA7FVc8ijOAuwfdS+tmvnu7JaDF5RWcXdS+J1ZXr7OUhElbkEjjpjKQGfz
11FO9aVTA01aMh0ZKvoS5TnjJ8DlijBjAIPPkimUI3L2sRyWyi8CywbiR44R2sdd
LQ1SMEQEmuELnPuDigVqJ7NxdZUHaFadL9EkxK5oIvM4zLBnQQYL4If5mTbpdUnW
5uRiCOVJ1wOZMJ+HEAg614lf9YdZcZw09nyDkyiWWzzXlsaEGp/FsSYt8HlOOHA8
7ZQxO4fTst197lANbubq0zu8NSCVAFwgCjR8SBj1a8WTo0Me8pYlmbuMeSq9QqVZ
6r+4VqdfeR0M4iabIhj8Af7YrFhhOW19a36ImbXoHiToj0w/N2cxRt6zQWHqlmIz
hKodXPIIzW4ITiutX3XIpd5+1p0qC08vpQO6mAlu4fZf5FPGuLh7cjzOotXqlnHq
WyTIBb1D/DP8meaua8ImLKm/qKRD+IeQVSBQ6pyk10NP8IyXE0fVmQ5fPotSNUMh
BdxYq3+BHUKff7AmhPm7NsxzTtYL/Tl5oAU63aZ/43kBlu8miJvtEtBE9in/X3q3
4q8yKVaHffo+kBmM68oaenWhZTrJi7XIDoAFKltoSkwR0zfnXK+Ak10vXjGuAQJS
Vrns1nUJsd0kWulnQ1cVWUALk6OsbtmcZVKQmFd9Y20Kvejvmo+6xxmkEQr5AriZ
ruKmLAIKiK1ia+tCCUNtP1TCQxWZ8EBv4cV0GXrwvuNMoBpxsLc+SdykV292zdp+
XmSB1XrPc/e7KTq1sCQETwyrIDfPPQ99Zy2CrxTp/FrcoN4wP1oFefcmmtXBL0WS
3hnhH8fObFfn5v6Zs7vTyZlUiPB/o86Nmv8wmp3MnZpIr1rEjrO7lKwcwTJKvI0Y
+l6SpobMVka3uBfUA7qXpoQcGD4A/RTt3XKoSsyTIVXESjWsQh1aMO9ofVWEqq7D
cq+1Q9HXK2Eb/L1VYr8vHUvZOWqEhqFFQDau2tIrZAtOiQ1rYDHAmTZUAV5LWoEs
5+WXmSHoKxpvD46e9HuR/UBY4d3srJm0XFLyJns1nEBYbJawsQFHHzj0fKGm5qFd
fanqFVLEnl8Tl86j+7xUhkr77M6e0WmhGmCBOsxT9ysLozmzrZDCvwkhkFJ1vEbp
rYFH9w7ItaMOS4y1GMKvI8p4f9Hh2gZa7wVaIALNWheBAVn8T5YXuXyprVNJHV/q
AeByv2SlKu+RUrMPE+DDlXN6xPzl/3Jycxh2RfQ8ybPMMUdZPNtXj4lJDK86gOmj
pq1MuQ3pZ28aDivU4ZcFI2g0Gdz3S6dCegthiBrA5JLr2mSlLwLLfIyrPjx4NS4y
/XzviWGtEmqnmuq1NP+wA4Z1yh55GBDY2paTvNru3PVIf+4K5BJYIF8P2Zp/uEs1
mLkmIgPhsHbsHPkRMXbQoPMKY/7e+4tm84ETOwZVocA8h1yrq38/Umxq0zPJBu0f
1tZ9+fy4oIhGNycguiwuwldDP9MQjZJuZIYhCCCWFJyuXksN8VyReIATMWUbnHGm
BYgj0Yck+UIETTKuLeiAKVJGoEFPqNvKnV/gGNLjQ0Qz4dTJYHsmVDM9r26N/4Vx
g2Cweyv+cYbq+2abfxdYEkc0pz+FjXGf7yOvbPMAF0RmSMpSSJnkn4FrZUsqbGer
SiQPgwrxlrGFDvemjQSikx6ZM68A9LdYkHMkPxebkLIXmyvnxnPgZS2CW4JlvayC
liUQpJTuvqtFSxNbfj3TwvsqjZgz8byLeSrJCn7hJy26WiWsUhkGxw8+S1tJvU5N
JQDnrBclOAXy0TE3XCE0vQqW6RiPfpSONDDc3DrjFGJ3cyOibmV2YIQdxbJLnB5i
pSPSD10DMYvjbrL0XToO2nRyIjIzj1AAoFC95iXMo6C4CYNBPwftoyo+yYZQkChY
6ZcI4dRcP16HWX7IJsf8Ynq/uY7g2QnQRnUDQB6lnQ0CpmUuQK08ZeaoeQxuQCrl
ODpbgnvAy0l18361FjhQXjlSa1Fr1ufMrl3KOHJoEPWFrt/zYdHmRzspVvysYdGx
NIu55lisb0vyBhF7yXuLW/FyTEgkxBsaf63AEQXAsSB1sbvBqe4oGpTrWUEGCgOT
i3bY0502jqZXULvZ/3uArREK+FDJ+ppIInL/iUnrqQI0Wyr5Vje6Pn4DqXL1dhNV
sIi+VfvZvHMJbhmFu5x4JxI7jwjwjs8alGtZg5E8aLZ30ta7W39Cf9eRJoe1CQEo
sjtA15RfdDJZW5M8EWEoGJFwFKf3rZH/SSQeGm+G62yFPFq56wJovqlpzG45WFJ0
YPMnN4FezHUv9by5BRtIEnjDd2K+5xIT4vZ3wJ06uG7Y7hQtKN7UJpPAVJ+UICPE
UMZV/YXySJowmjESCigeDYmwXtwnA2gZOXYE129I9BP6Myiwh4lWJNH1TrwsABaf
uCs0zfvea+LuSYGM+YegbQMn+WaKZD0z49TmSFwmljWqDGSWbpVKaLEX9UAn3pKe
yGGO4PE1mKFxV/5BilTo9wRey1P7mRbNuhcDnmVbHGldn3RRJBBwmBbE4M6ZW/HI
WEymVN3Q4V8vyg++z056YGZrjmuEzeEPZDPJ3YS4gD918U4/eEexOYmt9eh9BnXo
M5VD5Kva6GWHH3lErgPaPwwxU+WAfMufkp7hcLUFuc0WUsCw0bbaMgJXRl1aV6Ks
i9nF//NRQjJGg33RIbYGmBwa/Y+7T4H21K//eIjeD/ovIwYTemjwCQW6CUpkrvOd
PTbTOfSvuEPuH/OqhBedkxBVv6Jes28DFEeCT/jDscH+IOrjhjm9fGnwCSHZSzdh
QokFI8YNSpLcEkz2NzhQOeTnY3mrGUfqtstn4nzKLfnaRS67yQ7CCKMhvRGXS34P
M61YWUjcFWhgB73ptrozIy+VgZ45tqRsHGuuUNRf1Bsfa3LLXx0ZB7BntmBOoKXe
yTfX7pNAEgSoFOYxX2CNWU8jQoNwUVvv9V2WVnCJSz2/VsPH2ZkU/gXr7WL1PAs4
azAqcDAHnd563eQVEym8bo/bs4Ck/ZrCLQd0U/2fumWsv3vSVmzErXASVcKfcPWh
ieMlc56yM/WXAr0+3ffMrqRnDDPJaYi9KlU5fyer19OShU7Hf77EmU9Qz+MWPxSJ
qrrxg0JgavmMR0++p1vGP13RaD78yES3Rfd0hWOfq5EEBjFOhCw3K5x8YXlJMAAq
yUV3SibFSJppF5jzhrQcK0930YlCD/NeSmkGJO+5KZvR1EBGHN0jPAzmMFFYnSy9
9DBRVhIKyLBrFCiu9qNcmJluGLEAko9ruqMqe5ltK/rSCCtIGbWtcYiHLsFwEIQM
WGwZqM0Wt4Go301UN/nwr++hw20XbZ4BHOirbFHYiEPAAR8ylRGyeaDpP0wBIpyM
tlqlfBkcTpMYkIgbyLGC/BPebAVZCv5e7xT3UTDZxEia/u5jJvXZh5cIozeTdJIC
3DQtGJ6aD5+TZ5FhtfMDT1N1nkggPEHACIlSpLHbydWNsJFYevCEMUvBfVih2+Xz
0twChpGPyPIffzIGrzttp6zRtN0tsm1K1ODJn22RbKIhTAhkqEwdmKhTMODR3gi6
AKhhnUgfm8QWw6Hu8GVzxpvasd6ndVZWT64EO9UD1WcUWKXU5zmgpmniTBEEn5T5
bpyRRhtZePghw/ohI387q9GCelIyqVrU+17h0+emIf6SYQnejSjFzi9zQ/8XsKJO
Pf46mdLe6st/h1xq/m3npwroc5GMmeskVB9XTOOpAE+0VrWuTQSrHHc5EBHdsIsc
7t+gRjUJFDgkPrPSR+MSEK5VyS3jRioiMWN40J8O2yOtoWJkJ/xY44B/ZGjYgjR8
+WmMNQPeZDRULm52qZu5I4eQV0ALxq8tZe5xN1YT+R44pG8URQniuQ1L+gFDyzWD
o9y/OojRGSdVmMI5N50kJ/7AsO0F5iZ+q7S2dmueE8n9Npyb9mVxU/RsyYsQMyBI
3f24OMwLMTUPYKZWI1BfFwG4/CwhCixZy2ZbImBkSmQexPMOxRGBkHrivsggrz8y
9UFYPrvmM/oWy5rp7Moz+CrMnD7qCr73t6hRh4eDtCR+ANLXwgUpLvic1NFj1CsJ
hZCS1xungCoQE+HB3Mj5Gm4AnDTvqWYpgVxnPuIh8/6MWccrWchzoZUwDHeZp55d
eXeF2xc+nBy141Yav9W5zEJSWHYGjFAHSmYJ0938sEjwlSK3FrT3dcTiYL3ElYsF
3ju3/eb90n8g1ETHuVd1Qg9j77KZ4JBkHfF/b6H1oKiscO/vJdbBrhHxdOf13Fy5
/MsKpu5jqhTVrFLxFKsfzU6ktaLrtuC0yRDmYcDndS4jjimM+gA5ULThY5R/wIKo
A5Q5wgGw5RjHrqDlaT0/Kmc05Wc0FmQjXWpYd5c7he8jqSGormJzsihLCW9868Nc
gjRhjJneEwdQ+c8/eUnSzLxPeb3BuZpX6IJrpYNERN+TSy0ab61VEMtKnumn0A40
iVt+kFIlB3DiXCJ+QvrtFA6K9h0EQ9yZ+yiWP6KxjahDz5E7x74FyBGur4cAFndY
KnGuDhKGIErwdTHz0/jinCYkhAEo78PtnJKZf3Laz2VnQdkOEHyT8LUWRsSyyiEE
GdZnf039hdT2RsrSUAnuNZbFGFRbOGjaZDhLJAMyv0PUcejm57gqorfMj0qzVkim
gPuiTMhrPj8YnRTsWsIwPgA+GWdqViJ3Bk+GiW9TeZryD0icn3BFUDFaZabgW62A
YevDqvwL0wrAFLLV26nXh6gX3y8lXWZbwhQLQU6DjJzMC6BLWYJoTuCzWagaPaQJ
PeWdBhRyWh27BtxErREuSLfxhrTioz2d0tmlXkxSWbpIIWAdnOG+kiKqf0qOXC7x
QB0ig+K1ahvNIbtUNPbed4nHrZkoNl5K4SCi5VvizYb4qe0C91g3FyZ3ZvUjQyOk
w3mZWYHFDC++HvmCpypB/R2GvsMhug4GvvIDbB0E5Ds7Q5fvaLCILbxMNwjsOaDo
/5KpMvuVRKGuUzebRVEFybKMXLXovRTTaDs84jwkxgcbZshwi+PnctrB7rq+jyQB
BbDcgUWAh1GfPGIvCL8nD3qLy42QjjPeGSAg44mMsqBtG259OS5Gi5X8cbwNsKFl
oHvvL9n1PrictCAojY4KNmoCx/yewt5HSxG+5XEInyxAQ2EKMEuO33mDAYxgKQP/
0eS0lQClzgKiF3CEhkCAKzBH7KiSYzgufRTONHKgKpGel42BVECWIWsza4T7ZkD8
4RFE/Nq92DbIIFCFAmA9VB52C8s10y5ktFE5QzqYGURwxOEt0izvglCL/6U03fSW
3uCSPi5E5DkydfVRzY1VNhhNrP3/C2CE0uP20d31cER87vcLQvNtWpf94UotqvRj
lT/1g1AiipaaRKwnNIJsVQqLMH1YAMszD1OHvStB7rxVGf0ml2MqCG8yeneiAJc1
NeJmzZS2x534UkjAyeydIce+EQHVT5n21lseRgI+tA1HLdDZT5GgAjL2TLjHa90b
bRAHzGYvnehYqjuizHnBbd0jbiy3C7MhTOfO7fRscPb+rQr5THcLib0B57lU2wL8
s/ZltKo44onxiH/3GTJClYl7/RJ74zFi/ql2/nExsL/SjUbKPH9LM6Ffnd2M5Gf3
VMc9Jh9BubxTTeh06zRaajjnzm5Z9lirHQCmCaqdBv0LwwuYsyggida5qjKoW+vd
T0uol4lqDxNK5hbKJSM8fB8jSXqZF0SCGpIYTrDc06uhJKwz95YjPsbsqe0Txi8T
DPLKaA+G/ftD7G6ajQQyUvT1VEG0GZtPL9gbra1LMd+8fuUPkwt+l42s8MpwP7fU
K9mbDPOsqMaO2379K4GJlHpkK3IPQylZ0M1G8GwRF/ySN/y1BMKWsWC+nssoPWdf
bgu9qPAaYfQPi2BlfNR0fQla5TVWKpzCuJbh2m//Rw+r9clvwdJBIZHWFcvuOoNQ
FhSsEEgDMI6o7aAwZN3R1sX1peKxoYsIpS7GVV+Wp2MuzhJbnXxXTnVnjXjNFXLa
ZGigkvglR2hZDlLnapd2WzULct4zUzRB+r8Dj3jnr4FKUXH9DCTaSKCEieSV4HTw
aT4O+VAByMIhNKAZWPJkpb2ZpjfWfEq1NdnSGalETsDoN82WX9nWvZLRZdDPEJLD
BFWLdhDLwnSOOP1tS9SEwCDljjHevH1y26729/szTr2KBtcfRTYLIwvFGyUnZi83
AACgnOYazPpJkjSAclo/RWO3MU2JH5xXWLMpeq8jqrf4FXJGyfFgRcjaavtj569a
FdvUWiwUuxCehkEdWFa8jrs5dKNftvGp+gEa/Fov0LuGd6hItUdpah2iOBRaABb6
UTT2m8GhxXhY3Ems0+ZiPTBKpjpy6jLzK3ZrGDYKBRk4IKM5q2YWHN9ffvvZsV0i
QJSVSaEDmHKb18fZ+qOUZJinfTkxIPNi57xBAw+NchSNo/WUzcTU3C62flSw8ShH
sLjk/kM8namNIip6Ks5zsyeNQJNPQ7rYOsM91LElLeFi9XMgVAmsB0gJ+44sm2gD
bVCbVSRwm9Gpi87WE3Cv411WiyRlVw251kXUGb0F96QvRVNjrxthYTuksDwGUr1x
kQ8g9v5FDeMFhLVvotwfRSBIuDmGwBwS+ChBNFKKQ5MQYmcZ2MERIJrnh2X6Rm27
OZHUBsILYkmE3sXHuIlSzR9J9hR8MOAWMknvAvHpDmfCgjYaNFXKjXMolJaF3THd
FfLONuj93Er9p05CT5WcXIwvKeUl5aKZYCy5qdM1kikH16EoaqFB8zaiB+vtZ1dE
XA/qCV5fr8xncMnGBvSFIEiya+KXCw9LGnMOfiwjBCDBUIVvucIcU2N3SJZX0zWE
laanpt8qBGXt0jqopsjj4FwQ/O2vBvx4e4HoQ2rd0jl164ZIlAWuxBurx7fHic21
Vg7VRnLKWI0HLMMU8Xm/LhCGlJpLcOWfZEBu9+jTut/9mbRb/kFYOXbVP5zn+lA5
DqPufdf7GMgT6Kn9idGXfuklRRshkOOVmDyqgUCiP02GlwRHpIGoIwfnZTvcAUCk
a2ER7mqK6bM8CA1ryC/8rncsnS4UP9yrzSUmc8mGYnmgiP5wnP/y6WlQxPpObMFg
FBR0b5QgZVVc9IXZd1UAwtxnXR8DRvbB2u5RlORqVPbK9UMyRFKEfecI57Yti+bM
6dEdpaEjWGf9W1xH+p+uR22XW7Cr3wYAu/XGzb42cHeEyjTtzTijRjx4CO5qtwQB
k4mGZYNsLMy110B5CVCQKTwSjXuYjHdGQCW9b+7hvX5/eW6KpL/nBnAVfBYpoCd1
3eTlE2BtkIasJlR4FrQepfD4Pb88Qtk6Ze/UVPkaHGfX30YXVPcRuEEjPmrxdUgD
plUOuOcPdOgxdQn2JhOQLBkJyjk6KpBFCVLfkQmdXlHypmDI3XPeFuYJKNbploLE
ehmCwsNKdwfZgmNKNzVbXfR6soek7IreqPH2XOMN7ExJEv4u1sM7Dbep+mL2Cv1T
gqH+AKIxMdYTXb2XdLoKUbl9RkDAJA7fSjX8YRkf/juZWXkuVF1h/JEa+XRYAfaC
8aLRxa+PbpwU5WL2R82cUoOfIgxKX/l+znBP7yFlryWc4hiVroAsKZIDn2/dTvK6
unMvXpao/R9tn02tfIOWGsyYWqeIfJ6GIhwbk92WPL9KwFZVXaMxQAJNXx9DOyPk
2UYk4z18xYKsq0RReFUYGHKDg3XyeGRjKhwZO28yQLekc9AahXh6lr3855X80MJc
2kowyRQSVQyLXc3tbkUWoRCV4rRi1Wl+XjFIdiaXsXP1gpILWHQYY2s2Ib/ZX+jy
varlw8BhultqAU9Au4WZkrySOetpezhetItbaqmaQDITEzKsMjpA35TUZlIfeIlb
iH0vDvSGM4xAMsxczUAX1XXDDoh4vcHJRbFWGxvRdWImOWGhzA7u/jIbGs7t8meq
/bjDuF1rcQO21vvrca0Z/5aKpX1VyS0x7Cdbz2kIeCsyDWdgJ0NtXRhSm5YJC3YF
3dxRsAZPYhsD5UxCEhnKWVge9PA6AKjkqKAP3WVj2d/d4+3CGN/j3r+aNmgC84X/
NyKtIGZRHn1uYnL8CKw4MclB5RDSUSyxYV0gM3QE6WZZuiXWUAHDo1FOToLH5eXq
A5MbzY7HArZuhblmkUIUda4jj6LdudF5evm7uPIomNpNVx3InhD8qDCGD9PvR6b0
hSw2KPFxgwo7Z2oKl8RPCaYyOnAYpylV/N2U7qBW6D8D3qVYIl3qNKrp8yG56q+8
wgxPq3fXgDMQhBH2eGwubqv/Z/n7b6V/nf9DaEfuZhK676wquOZ5qAQjw5nQslZe
QUa9T61uLJpEC3Xpw0/pBs3EiT+d2lQRmNUBa8a8IzZy57n0/LOnp7b2rAM/2CfT
si+LWMbN27hoYGYLZcVgn+N9ul5ut270tqc5r4e8TPF6K4pdc2j5LbWTyaem7GZK
7r90EKLgaYBRaAlwrUCpa8paCaNT6Ukl4cycyNRE8fTKVBQ8NK/UiY9yVH7ysBLr
MHOj7LXPUzqU6rTjRaYvvVDacXZClzp5xLR7emrp4H5kiL8A8SaF7dtUMZUaenwU
q/wXIQBk/6MMTBgsNP5XgXHUOOcRoTM+5R1zK1LC1hC7457ZB1bJNfeqEtM8JaYA
Z+ZKmZx6zuunNtds3nIHQK6TOHESvfNsJFqKY1hsMbwYWwOrwn2+QOHsGO/Vo9sj
KgXurn84gWVGeUeMAghYDvRom4gy091eiaRwxl4NR+pSyDdnp+eC2wbkR4DkEOKY
rEnSMeqluJQTIBN0EytTSOQCx89o6rt4KqeJMYsl6MJyTSo9N7uVoONsyLOL2jLt
2fCDO13Uj+CrpJExRgJiaTAuCpDnGZq+ft9ugZr9ufP1tKcrmmh/VnEOKgcWXU17
0f/noDDOIyIex6af0YO1RGfccqxTMmxCchR/bLd4nI1RoAmz8JK8htb2/H6GNFfd
0IaMz1zYiQxocMyScroIL05RNm/u4xR9oKKp9WDvV53uSDV7ctyaDb6JqX+A5kiA
tIJ7Obb8Z9XkH/LvvQmQ0h0B8lv7wkkc1oNtgUczV/fT7fJpXKFbvR9/PSFSzygN
VUwzGpcN9/bsCKk4xi7PLTMhmNrjo+4IZCp2Ka8dCyWP4vh+qm1sKNxcObAmVgjq
Lxqwf9HvGp94A2FJiNY4d3phAZmwzq6eby2GyT8bn/1J/eUeQLCtEIxdF2TrZEdu
rauNX9hz2ND4vJAM1AZKemZEewotz0IERC//f/8RAfN43ONlA1jEcgyMdndhwWVp
WJXnQ0Nfjohig5GiFTAEWA8zXY2CqjIsWuc5AB+PcJwTWG1BPeDL3IkZEtWZDlZx
w6KkKODveQ4gpV+JksvOUtKmzo9Y70t4rH+Qu3kNCUHZtSr8VGgA4R6HOzqyudng
/mvcudwarw6UBcbE7XZi2dJUGk7QyhUCNGbtIQdQkXjw4SIpynQ6e1l+Qh3CW2z6
M8dKyYVitMqLhMyTEeKhe58ydC4kmTUCep+0uYaAl5uM69LtBVZK6VIUnxdMMRUX
9lEnmpWnxRXqbM8b0XwSiw8FBjoMS6vq185gv72TYzrwkEFgLBmPZRavQnq6mkFm
iq6zCrqmAijWHbWv2LbNQ+IeWkVOaCgB0zHeX5PmPbboZaHG1AsMG3QukUK7stAN
6ZQzMPYFHbIYZlvnnNPFqeKtJjTXCYStLD6omZQIhzt7W+wV55In4X0rV6w3wjgv
1eRgCrGkUFtd7WXyGsgBpOkThs5NlBZ+BXaEhtPCS6yT4X7fPnTm8YeO6Oe+pR7S
JweG0XW5NEltM9OEXNgD3bXj+pPoYUb/Wx1fd/H4lCGcX3HH3pdsS6JkN1NYHSnj
9IOyrtrrvV/CeoiKo3koMJZI3gZ3lk0oYQZX6NxL7Yys3Aw8yZ6K0WxjJgkfToKC
jraikJ0DuawJ2z0XLj+3OxO/VKsozFRz2ryLDtSx8/+wIPQoepfJjXp7U5eV6do/
V4EbC7MRFdHWOBbhn5Gbnvqqt220y02prRSZUIfWFqVQw74I7lCaCuBRbmm1yPbT
WsEC6BE3H0AsBHyrQMjdfY7EuyaFJMjkMGGRgi2kqkCtYDJ5AtH77QQGYld9OjKZ
lETQLaQBeDeCvfDdchLhw2cOl1EDHBLcoqb8Y51B9AL2mkKjpKjF/cSWje+AZWUB
lW9DFeGhhRjKwzw1Y3BrQjV+4RJPcAe8oR3JbuvILQam3pir4Xq9kpPsVAVHnhad
07AnL01fBQ5QHCTeY/49veymXUACC/I4eWDcBEjU6bA+ql/UMLtVhA/XSWAQxZvH
K7splXugTt2UPyyzck09P4MRZHsZulr5LBxd7TKxjOL1obez3GmqmrZRmAnHKqqP
7W4z0eD+HEg6CSUUCyxbj2zLQx91jUFmm/I3GHO20dXFM8i5o0BX0Ijt63sbHGGP
h0L3beVvcSr2LTJ5cExN4aum237usy6hDihT43RoFxgEWtgoBCdHQSl/Nxlf8lYe
uakFRWu1wUIi0ufanewjPi6+U3IBEBbv37bUSPM4Xm61kkBx3ntQWJHEKDctnohD
obYFAhNWN8f4uJC0AJYLDfwJaUwL83vlBthuw1t5gtHgl8p2ysqqRVX7bvDxPKqY
7UEskYhJ42Cl1ZzeBFD5AmmkPCW+Symu/HEsjCSxJTQCoWtGOgTfuksfgGx/FtPN
JFx+MTQvLhRBTAwW7tL22elcjLiBjLJ4jkd3eUEKVt47HyVQGG9OGPXFn0D8ktR5
xznq+Sdhfsmsq3j6AOJkIJLp8Au9d1TKGlmMlrrBNayVRE7WJpis2K+LLtzyVhaR
80hJ0UHK3IQlbpMeduNqFZRLsRhZU92RE72FI0eOhmauV+EYo0V1IyGczcmc3aK2
K9Bhf8x2lLe3cmPJzE8xGVRtlrJ3gWGQeq9WFVLkA1xB2sRa8F/dYzqwI8Leu5vk
UgggAiarplAzRiE8vl2lP2eMuMVDOzwweg5m9DBZaE6tTAZMkb00cXBKF7GBat1w
6tbi6j2lOz+/yMZr6VItxoxxXMno/sNhKzXVAMEY67ajpST+QNYg8+x1YIOW3Fix
roGfgbdaHkaj+mkiclIh8aTcSCLgPB4uLIZ6n1e9tuschpxd5d2th3tY1TEAiMec
XswNs0hiHzmyOu6aXexZrAR5m5ZAxDFazVY1+jqfUdhcQe7RY6WYPIJ27h6jvrvu
z1uZBb7gzsZTBnlOqEBUuOz4YT5vMYpNlABdyegOO8MRUPKVissqhWodHUedRX+A
CeDZTBUOGBY3cGtZIX+ouMQc8gWYH5T20S1Ay9FjidH4OcFaNNAkS09GhUUGhcm4
h75KWEa6MUDKpsyM35H+SichwNmPH1PmeZZgbY9E2DlC6JHDORTJeXBH5aK6fyXW
7T8Txw272tTTXfG335JlotK5m1U+UCfeHb1mFJjDUqCfc1pzHBhzARS17gBE0xgN
yV6Rj0Vom9/41mUMW0yuPzesC3VI79CVVZClF5itBPFTQl1G8vtRCsuoN1GvjCDd
l3oDRYciyGbqhweIuzUZeE2ZCjIniWy4fn0VQCMXcmhEdeCWnjRGwVCHIMT3ihk6
X0Og6ePM2qLp2Wdw7kTybDulnZcYm6a9Uu4kC0bHSjTTVs78ACpBCm+ZsglAtlfN
rntWEu2KDEb60FoPXZSXVjfCF6CTB1Qslb5nyIKyetYpOE0vYOMQhYc3YMH7+g+H
yjdisgVLZrgrxmZkZyWNm3DEF5NSgBv123TlONjtqH2cQPiEZPOEpBM2qnsHboMq
yD2cOHS0KVnnHsZRANhhsgzh1YFegy/xXdYkdOsejBozzGT2YgyRm9tO92bahbU7
VvcjmRY7GV10ECMIkuL2Bu7jleLnxLMzycMhQQxqQmDS8Dl6kR6lJlXR/HwyoIVN
nXYluz0+OV6nXV4ENdCjr7GRMHPMo5tH3fBsY3kX8hBjbOQXy4u6LOEqKew+FWC7
cfAuFxerso77WnjLqOHfLw8KVSO6xJyaSOCAAiqEQpQebXBHxgEkuMJYjCu0gU7e
qMDtkGNKKA/ub7D2pZgefV06fHAe2T7mbG+pkaDrSE4pB6B/DxMJgMD2QjoQ7Y1t
G5ZWmJpkapkxrxALGrIS+/AscHS0UOwlvS5J+ojI3UdwcqY96AYL/BpNc1gEifLY
PpdwoWYQLeKaI+WngU/JcFIK2T4StIO9sb7BpnnoZvHtVEE67J6spx+8LhDWFBEb
vKr5qpKYj+i1J3rtLwuI2uN4doTCfJ6CU7p+9dJZLNwBdVFucPWdzD2iz0jVTJRH
bJRQ/Z9g9lqvAoGKc3+8p6vIF7/rVuroPlxnVLfjORyezJVcR2WEFA/UQ5iOAMdY
DEJGv8whDUlhx+RtoxLkPd9Q+KlyclspbJEnNxXoyqqPzmZlolEZnV2gByiKyv9x
4Wu4VYlCk+O/GIx0xobGQvnHc02ayPIUpidpytpnnrGCIGK1bSSIkt1dtd0B3DOz
B9tjjCs+S58OmBt3TBjzWyoXOB1Ie+zhYGSV18USUfz91uE4YjzyHu9FuqwCnnvN
cfa8Z8Hfzojc6Xv/K+jfoAkwdSQ9U0SssFGTVKix7JXRae2x4fEBHdH7M1JS+f3t
B8iYZqeBOgiyp2LiqN/zwZ5etY67/AyF3e67O2zdzQ6bwIBbSEf4wtVKLWiftwVd
GY6HWuD5WaKOM+Ir0fPL0dCDuOhl+Ma5cN4Dqh6dRWWXQP/MRS7Fs2njhReH9YlZ
VjkixyPKplXnn1Dum4xhxPgru9eo3IVpNQLg21Yy+MNC1BdqaRQXwWA+bgz9Ia2E
bhovG48KO0NNVpJO8lKFh/CSeq2At5y9ARxB16TGi/BmNxQui4nRDI54rnkw8YAm
rQgPt3eulKo/n1W1/G6XpTeMj5FNIh8+uaxA8HjcpBCAPDqJ//q35sXAwarVXtPt
3VLxbqmPVidIJk+2l+q6LYRvUrzF6St8GiJsdcXTbCgloU/r6oAvi12AfvbFMD2j
X1+celt9ATzGL35wa4lCVMm8fyrQtJk3vpy5S3gpIlx1dAnsVmcY7nYztQXoH2Y4
6Dun1yc2ed1NTmALq6G5RCwLwvJPRr30yf/AgFEob2edGFiX+kL9/1gOAbTeRhjH
is9o59zU5nOeZKrTslpb0dK3zo7q/dI/ZpkbyWV6fZkjSX+3vv2mw3Ubwx5ORRWj

--pragma protect end_data_block
--pragma protect digest_block
pUC30EPGb/cy1Ms7X8iY4cgLkIQ=
--pragma protect end_digest_block
--pragma protect end_protected
