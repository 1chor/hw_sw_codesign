-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gRF/PnrRY2Itu0YwkKuLWiPvvhs/zOu2eh3EHy8EBTL1MxgmoM/CjTaEKd8uhF/Y
b4GIbybdEKyeDyg2EpECEW68xppoP4DCJXtgIkYws4Gjf9T91I8YJaggG6iH1WoO
Qg6GLmAiWAePTFEjXrJ3dAxNyRANK/05dDmfDDN5Jz4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 17442)

`protect DATA_BLOCK
xmOM8uo2L2oSdptsiFSVMyC4tzcFrO4G1ArX71aE8lmrXHMAZlSIT7gGMjzrlEk6
y2Mc4mkSkwiTueJm48b5prEWxdBaOxvCDfW/IByBuQnmEGnincTcuKcf2uVQ67C0
5bDz8YS+MmiOd3IyFZcOP0KPvo7B/untG1VPyrv3J0sSMsYIAdhKomrSI3VZrNm7
YbIoy/6QV+G+E8Xhv+GiV11N0Tk9oaDTInigxW5odC6p4MnrlD7/4OO3Ub18w+pe
Bq94t7A0671OezAsVBtJLT/ev6FitJl4Rt0n8XSa+5XzAk1GJzlFfKKrLykhzU/b
P82km02lvEzvVI5skQjxZ4QPsx9KJHtizOnO7wU/XB/BzHS7Eu+wyC+1n1Z5Fchm
K1/1xZiOiyPOg5twj+fcVUE6vumS3E8XoY6MSETK0go+zPQF0n69JcRs5R4B26cv
chFOJNZyecpHNDGKXPlxPUqtvlXeTl8clnrNhcILyrqaOV2t0QVOXw2B5+hc4upg
HbSMwefreTk+KHwdaCpGZ4RosUFgMp2MNHEOzUX9H0JbNsl+9cbXBDQmW2/C4Jdm
QhXWODDu9pYOxGSzCdPGD9EB8gw772LEaYtyv4GHdbw8GYKJtYP1673QYrFdrn22
OFeEgqRFhKn5tExtphH/lVV0gwrsFDxnIge8f1LGmrfrpZCST00X7pKTebc9oart
u/3VyovbvrI+zwYiCsOTl9rD14GZf1CO/i8TXVmaa6bY7TvPb2m89Q7mrw6p/gSd
JRyQhIINHu28ULuBsKVV1YhWlffd/K2sfKubILzleR48xK+/dwlVrZggEj3YgSmM
AoohIVtFwkvazxAGCRkfVmhRYnzGlZ+aiyfqosulzx6VB9bKY1nY8Hi5wdrD9Uz5
kEjEoLJEN2Mt7D1Oi7dV1qBCnCl/1pw2cEJ3QuoQ9EuxVd7giHp+vX42r/hR81QM
RnFckfzPIJDcImlnk5k6w/oHk6HVdf3sCR4qslFwpeZwVCQq3ygFEVrG1aJwrEhf
mASQsO7COtdHbtQ72lc8bcZqihgC7jM9rJ144GmNvSJVu4TMWd976+v4946W+CzB
RXctSzjnyGVwMDl8h3ijpSkT5h0qewldnyZbJz9z+t0RBuFNu63DWN9o+TxqRtdP
7kT/N3VshuWjizvfUZlAYKhiEs3+UkhGaVeHYTcbrUW/feC+ahPE98k2riGMNy1U
vm6Xr2lIoWUbnyezHO06Z8CLhjEqYt0Gu275UPrGbWDFcs9vr74b9qsRObynMtQ6
t+GNyx029mUfhm3wxarCmu5Jxo6+E+ElZkyYGC4X4f7MO/MOstEaFYUTzxDPiP8z
hiJB2fMKpuYLFWsDENwskGjluh2UUINdEXmG7G7Hn8GeiHDJ5cDIp8vJBF2UXRsz
e4gFHwbDQ7J5bKMWj2LHsDske8yFwIxbSEG/eAX+JfCCTa029uRBJwRgLACbNa+o
OP/a7SyTzk3vAKVdRRatbO6COS97BXIbcEwrzW2KylcfFc8LwQ02yQ4VQGev54Do
wFFr/pvwN8gJs7au622VNRO0FaVCqxp/T32lLJCsE/HmZn8OjvSS57+6FIzlK59L
IgMyM4qrRQ50AihwdPCMNyfG5dtkQ9S8D4TOWYpAgIfvDNLUBFJlMGnOuJOzjHyx
FXBWRqxm0uzEEar3Q712WCFQIdkG2oQsVr/iMUahiwSwDd+dDlknOMe0VrezxXEP
C1vF3SzZRWJwFYje6bksz/eMpa9QVlj75PZr4ZrcUbsDWiP3xHKcqpqOqOoXCc+k
BqPtGMMzqLgffS4uBOsL+N3KIUSZhrwePywPHffsQeH1Iu6lAqy16hVit4z1UvDZ
wja+zuMdhE89p4UPoQfJusYX15OhoJJmP8hOUm5Q2Hty0kXukNbhCGcXRE2VSkrO
iEe6MNSoIh/iIS4L/28zBtcT2EfBI0J36f2r78bCRGAtqh3zW/hUlcsfsJaegKoY
Zx7g0oXHV+O8bHhUthEswogae8lj5kGWK6/Lt7I6VVy3C9NTMdnox+42d4opECS7
tRvttTUHSEONtsADDaCDsA1eEaz8h9OMBII8cDyjNtGUmadHKTunanJHe7dMO3Fi
MPJUua7P4jePnqnw1zKsHc2HiZl0NAZw4jYc2V8ATWTJWUY9cQPGQjI4sGFaAYl4
Nlf1QECPBjg3XxzP02drh0Kt6iH4/sIva1vCXFqvX1YzPyQ624OLBZEkqoSy1JNa
v9iVZgsoP/dlo7jn5ckQasPakm1xN9gD66iBrW81eDmBHa/TrFPmKz08NConYjQM
BhzBZUsgcobFJXcBgaXIZdCXC6t59mQ8JK8bj5ZQJVVmRv0ahwjUvz5J4QVAVVW5
vqzEPCyqtCtL65rHNnuQ01mL+Rz6dPb+S6njHNSBPm7PoHI2pUmNgE+wHtNjAbbs
PFQA0J7bYW/wTZBl4S6UDX0bzoriDKe8K7RH2J6ENo/WIxJmZwPnA7ld/czn4BJc
HSazybpvNENA74qL6cldWkINhyqTghuG2PN5AH6e7U0mTshqFfN55jwnecqJNnk9
OZObwrAq4ADj+6z/SV05PwUA2Qp4idIfh/n/nW4AY9iLvsX9K+q8XI3xa+joUVFo
GgZf12jY7vdt2nWj/lD7FR2uh2vHlaDXCVfpJPoE2N5aTkDIxwgN3P7lDU2VoVrD
sByHnI3aEnue8TYAbpVBUd3yh05Xbo46BagKJTiSxCYHQWKqmo/O1UmGuplZaSbD
7T4pf+pGoCG2L/q3YM1HkMNRtv04XfR3g/vABHVZQxR1YFoSs/wl+58BoY02aMou
xGezqvXb0HaofN8OLszlSOxXYzCf5nnczeHFaMZOmRfRK3kBrREtCnDMuZPZZ8P3
et28J0k+7BlgLsDFFPyksbgEv92KL2f7Mfhe7ThZRRdmnkTlBwVgZDmyOzAHpzGd
CE7/difNlxAVmMwtWvTCBdWXmgao4dc7yB+tSqq91WAbtZFNfcmtztA4ZdE6GLs6
GOgG1g1V2vsDhRKS1XF7V/JyvzFrdePZK1ifesK685V6uVplBjd3LVUTNs4686ca
ZVkSuNBhcDu/bSczqxmFFUVHUMcLMkU2oeuJGdGct20iMFdZK+zeYz7lbqM+XitH
tIGY41T2pQADbibkF4BA4yfj/CD6I29uSpRMmJ6jQDRJYi70aoy7yGFONO27clKk
huASrONbHlrtK6wWx5xQTI6/Lx+/CB1pCdzJ7q1/ssU5ieOSJdxYUZNOxB7zGh9n
kumQf0INmKPkn0m0RXt+OQUvCjXkBIllM7eZqHCTB0HiWBOyiBQXKs1jxm+FhEL5
tTdWBwIoE6gioUqHEwnipqRvpxe/rBINL7ZTD8yQV7j7piW1QkQbJ0vgmqD2LOQe
gva9WzVaaGoplU5/xxRozQ4V88lU3tbndUwjGN4DwbY8TPM0PcrQbWebsHsCRdIE
xNf2gH/D2A7HvNoGen6/F+Sw3nXNxXHkDEnkUTqg+s1RidFchOtqVkwcm+cDih4p
ZnpGO7oyg4cDs7lbKBLMAaO2YU1AmiAPtRaKQ/IGCcMm1hkihrQ+lzLfF4KzBYMN
RMAEKyDOCrjIXpQ+vxDqj2IoTz2YIq4kcDGAe67K8OeIzouxVdPfB5TT8zzR3GK1
ZTZgzaqebeCJtYGcRyFYX2qfDvZV3/NhH2fnwNtKtWAIpiIBuYB6bm7wDQbVJdNm
T5mDqb8DW4hbZsALcKUpTQPqS7o2ZS5GO0K786Bb5awNyOMx0Al7dxt/mYCSQRsG
1qqlev/ZOve+D2swfiIwjq0aTdHFKSViT37+H8JeuVmnzTIh9y0Z5yEK0qE4Svv+
E9uNUeOi2hTX9S0QLuRuN3OjYuq1LSBPMju+UY1W8GJunEaYBa9CyTXIDPuq95BY
q4wVPtrKXX37z3DHDqFz0654fYWpya0vZ3dL1J5fOdrrro/vBguqCIAtSRyi2WCr
k6qkTiQ+TmP7l4Gg1nq6a3zQEc7f/U1SffoG4NCrEb4w0ZI0A6Uvcue0k6nfQ1bf
dTBzWbFGGmc6wibJc/j5a+WRpq2YQaF5OLksndtDrvLMdJ0cT3U/vjzPKMHoPAlt
ooVDtAIp27a2Ifpq/bz3exj2B2rb3cPpDo+/5EQnNNRDU5cPDVrlvfiGpv3AccZm
TN6I+gnVFA4cpOlDtx3jZX2XMSpE3zYKLezxFmfp9GdXRYSahZC/7ZCq3zhJiZmY
8N9uR8h6SXSXWjzcp2yKGavpmXb0NRcyiDMoh9GmciZyypzsqDyictARGIcJEiyp
qjoeSfominYgWixrql5d0zgOAbRieYn/wuuzoKE7BlJRM+O73vucMBqmRvdD8vFe
rDPNQ+fBdiZAPWYEm29wd89VRoNonV5TzTtO2jDvzBK1itXB5R6rTiszIx4Ccv/q
dx1b4Y2q611uTXEDZU5yvnZ1HDqyFBJh7HHUv6OjfaWvRSsWg8AtixuqrkJthgiI
gtzoQ9w59GlYUWMAM4ttNnGUU+mMfmmDidJOLNanUPYl8+XShpN37IGh+Jw4a3dc
dbVY1fZUyfGQneaPFCTSA5DWw6GyiqeJnIEFuovtTmH55TbHQYlWp4oWsFECwZk2
Mh9u73q0jQbx6lh8LNtQmAbrkZ2fQiCCeKzru8QiXSG5srNrM5Cf59hbMjLfXog/
sg3YApw3JM7s06fVLrInUq25oPaVvEFcWGS9sraCkGTWW30y8S7JOdzc4XYGGGNQ
TkgM5hnGkDa5bEp6qqcucEUoU1pI598vHIUac/6g+aVghUGPO1DHRsNvL+mfkEy3
l8aRs0luXlznv0zFYFTGTgNTTs+riksv04Dkh039UqV097ZZCOzSEuPuCJDMj7N0
qMsi2lxX3U2sW4iuxBw6vC5Gf7aF6iamJFasysoJOSjckANWaUee6SxOBjhUjcO3
Jxib5D24lTIeLE2CvbbWnR6WV2sr1SBuBiybsC1HFZVNBVzsqskXTAbq1CJ6+YDn
O3TaD3mkJy3NjpXP5DBKV98qk2QXLzwO110G7US3hQ+mVFENlI1yAMxbK+3hzyx8
unooX3XY9b2wJI5uChOWUs37LARkCUMTY7gf6BOi5P+9VMkurMXYcZ9axm7Mm7cn
g984GGmRf0FVsGUW3mO9bSKvsEkkbEik9921Di0QoKyn2DJ9iSag+Eq2SFEIM4MK
DsrpoAUA/yfwqY/+PssMg4eRMQwQD47J5WIjcFCDnVamiPcLhUqdeheDGDT+whyx
4t3HJSIJ2eJxZTZGZP18jjsz3+9ZFxyt+iD0t6035/P1EII1Mw1FNGzADAjKE9zC
DvSECrPjSQT+lUfjSBZMwcifSzydazilWCzkp21CRLOZa6WGZoJ9/X9QuSbxapg5
kePmoAeoDmNeo5KYN0X3sYPoqv6vC7Qvohejhbc/ZfWQC19SJZEJN/i+gexbXWk9
L1XMqLChlfgCycxO2iAcf8XN8TivwcWDvwnffAzGO8V9TbaBog0tnRexD9ohgsqS
ZSPE6MA6qhNwESXK7viYVbgWY0g1l01xuRTHbhQhpfq035yzojQEBiXOh1HdwZHb
T4NjToqXW21p93zaysaGFUEUlNa0iS2v0zheUq9zcARjsqClyqeUedqBtQP5shN2
eXGnByM70ybhM/i9lr82uvMESog8ckzf1zJghV8PU3DmrH8xrGgoxcC1zWnkpA2+
hrMK8tdLmCnZTsiSC72Fe5HA4WUJeoI0g9MlYmPsrgQoj2T9ZYgbBsSk7A7IPytG
1Cy286Xc2zH4zgOQWKPSGLD1nyfEsO4uyQUUGBcDP3GL9Q844xkw/SvKYvQnayod
s1d7iprYMurcGqXSnvDvhBYhgY/m7o31q5jpKZZExL9VxXEZ8Ki6FbqZSh8G69fQ
dHNPwChLSobJqmmjtC/uItVI+zsRZpvOvBDIvZTusL8Qd1zxVC/yUrh0JGskJwjm
XDvKXbNxs3wdSHgAjj31TqCVbfl74qefFUO9hbv6AZ/3x8FL8A/aQGH/7Rpo0NoA
5Ea1MMfTdF0psm+ynxbDiN0vdncgH6sROMFTAUts3Ucr8P3u+OOfUGyW0s13uZ1d
uF6NY7w/YG0zgrBE8Cxc4phNP+8gz6itm37Wc245w4wieHKUfPnc6et0WW+jqIlQ
KAlEDB8lOQPUHLenEJgpAtK7EXaXpjNQVbClEdJReVYLHXTL0VD6kwCsvQ/tT7OZ
AvEg7PmgRoXAsKtsAtDF1GsNId2N+ScITw755USBoClCC5Jd1q0lwmx5T4oZBlOr
wsFTNOILtaEcxXgmElPjNHtqz6QqqE3Nny59RKveKcx+3tN66t29krOsxEMCuW5Q
n0Mr5Ew1oiTkKRni/m36pCayXSRQnBh3NkVrtBKLoSjtE8PIOb6K3LxTMeGfZ8+/
KfOzZ5m3r2uPz9DgjLD77xdlh0SS0AMxgS/puJZTxOtnTYhLR0z4lW6jpnUaMyID
1y+sAwqD2lMXOl/ijr2t8G+WQ3cEU9WEd0x9enUeCg8YX/+e31bAfU/v7f/DUv3k
FwyVETalvThCsERcfXuu13a6ND4kJjaxEEj5ttbUxqM6AWLs/gw4R8ztuz7qNu3y
hQMuFtXD01udfaKpRSsdV/eMYWV8eEm8Z0Zae4AcnH/DvVgdDKGGWsgP4zf+LP6W
0ZbNm3VjJAKbF063MeOA+ufiXMI6OsJ/AtgQ/6JFwhY069M3u/tflgx/NMhfOq83
9eNsAiseEt7erVTbH9yaPHqNvSTgrjnZ5bLFWhiMrstDFxnn/FzdFKZJQFEYoyWI
gCh189Yl+lmAwpQpHMK+oz/pNSoi6ZljM/1Bnf7vkxxlv9FGTDrKeX4+cD3IjVUn
249Rh9p2IUw8JQQ3/Xd7bT6HfWhhOuqv/iG6pAw5SNaNbAGyucDxIQLT4hWZtqeZ
DXlaHnKBs8t1HyAlriNeEuraflfOSMuMtRMu2lIGdptsr2yfKK3DFnMNOQOYhLaP
ajseigiV4AjBGYLmerJqX7zSY0FaoU13tG2JxEMjgA32grvHlqkmScT7hEF7pcR5
XE4L1KvK+1Pqa+VR14ueL/eeK+9bwP8B1SURLbK7Wx4vPXjkYkwuNDb2mvfzCN0e
6EZ0WYaGuB2s2AwmWzZpWzpmOKHpSQ5svl7rJ8pmfLUI+ln1gt4w/Ek9/6dyoSma
pXscFOI5w3hyk2JmJi+AKgG91FH5wZE8B6mnlakEaMwBu1Tp8lCgPVEw48C1n2FX
cZ+1JsBDEy3wb7j+1Ns6etTRlnuAdldeY9+9sXTUuePt6RmZDJfDOob+1Tq3lQNj
uIwNBtu7XmWtwar3N00sH5tunVArShGaFvk5TvqE2VUOrlAoU0GpIZTKJux1TJ0u
VR8Ww4bz+dBrHE3oxxfmg7QD/MOjZ+4pDoB7bTKfTwmQZ6Eoeh2llivMtL+eCd/B
5Kf64570l3vhqL+rIpKRzjvfcN4Nd4mfQ15qOojQNnyHDzK3LOd/EyDryM/+6HZs
4vTM6twvkP2dozkFpUA4OomX7Ao3Wt6+MjGpsSV1v2cP8JVQjZ6XALpYo/pzxc6u
CRecvw0Lr6n/LsggwvKp8FcvMS/4HcIGuIgwu3zshTvQNsFOej7/+vUN/v44TxWb
r4DZxL+WIvJLyHGuvtNwJT90CnVB7mh1Oze3c+2MfmAv6hkYr/0cQlnoYQQz5SFK
oU7UR6px3KXcztV79d4vaUjXhwXgov9RSVdCoVRBcJ+VRmRQkH4raSjP/hFUqZnc
f0qkHDsBTrQETxAkbERCrQ7K67cVkYv/wknVab61onFgewyOwQzI9KXOK3omU6fD
X8O1KmZK1hJCT6AIDiPsBy4YC2ittdq+0wFQjSR72/LjYburravWOoabWMx0b3q9
0YTkQI2FUPkUvf8sINuLOYgv6Xo9SSFbSTIoayDEyA3LWNrtdXu4vVOmIGwECB1G
mGoBpuhzhKZ0hvSm3l7zzkf2ms5Ztd3xXJTj4s+kQXq7qrjzbg9RBfVzZoIahj9f
TrZeTQupKk0eAcE+8o46NMNBTiyh5IsvPgEyBQVL/jcd/JxH8pKyQ+jUTa/Sy0+c
gqVs4r21+vX/oEJnRTIByvuQ0w8vwlQLCxYQeza1DRoZojFVKPAo6azcuAE2Y/BK
wE0BjOmrz6pc/hjyua5vFcd9FzbjpNtHTYDqs5Nko2X2vqutWYEHfIVPEfvXaFpo
UbZ8Rns2xQvC1cH65A3PeC0PZyXJ0j5sHS/gRBaTFrequwaUVglPfJWiWam9+Tsm
lBfGFRa9DOCg9nQg5LGzLJKaJllXcKoN02cvuE8kQD+Ugz3ddVbTcBBTLtRItsL1
O4m2YUpeNEeseaVXj8T6zkhGYvSKcgUKOp8fCkcc3xeQBZr4g85Ej/XHPlI3m9Iq
WckG46Pght56a+BblJEyTb0TRBY5QDWbj3JoUnpqhrsu6J1Tm5Xl5udnvPFAYiYf
Cv43U3JMYzlFPBRr3tL3qWalb4bh3ArC/E9TMMqAeJtVAJ/yjoCjlsUPcmzork1O
EhadxP+VVSKeMkBxs9G7aH3xunJjTFpEkbiZ23Ag7LLWKvM0A4IORYVkOhdmYAxb
zLh9RFHeK+Mvj1cyA/veAwaB5FIGFHze/MQ111KTZAV39sNP+2gft0FRFMh6onmt
bQfYJbWhJ0z43RUC4liX20HI1DQNK1doIoqPyvDlZQG5LDy+QDJ882pCWtF1dU/I
ED+zDif8tEMd9eOjIa65S7rhEXcjl1xoAcEUra29WdEgFIoEUEYBL5KXYDVXyEpC
V1/4tsZeSeiGX3SYoUqGiY70mHfE07embYiuMHDAxGwm2zZQOtrixccNlNjhKavP
8KEV/RV4wfxh+MlhVEfVvtstsB8T5sacVp636JQmWLBOB54aMb1UKCYPnAH262bq
tMSdLSKf/e2iQ/FXUDP+iJuWTLTYC3oBu3gVKqW44T5I97DnThHj0ukvL6vy6qu1
fhE2X2J0kOv7SVYadCkMMaAQsdr38DUVtFASzOeszVovkOqHeqVNm10LJ22SxNVS
+vTOlQbEnWx0t3XsFd53A+s/LqRkzS8AlsRrEAIyi0gp0G4qXmfWWVBbLROuMXT0
qakjP6DDo5d3IGwoYmhUhQG246hOWCUVIF5B3yZLClBSKKaCPMuM0BRtAEOr9X0V
thOHb6g6fSuIdrTwmN/qiJS+xabbTSnXMqQ0lOgzpt1G32a5hvzjIdWLEJlTn6IQ
rzg52ueMRcwOQxcHpFnAw2TeguTzr3C093o7EAmb5Q9i4VKAhQqPZD7Vd42eos3Y
ClneB39L5FyTTnmr+beR0WiutAljoyYhZIHo6K2fweeNg2yGaVraIdTjHaRFpfRX
HL7epC8XhGjX9T5yP2S20i5pCtheb5xu8G5m6SpsiaAFOxDwAZxr28nCgpOYOguc
2UiIc5kvS3o9ixD1jAtAWM/qBQPr5U2dJ7yrE1P3YCc/m0HRyz4zWMUyKq4EjTBX
ed2D8MDbTun8ENEIHcsfw6U9JqPhN6cqyR+TFgnfGbdQthsOYVnNm6TLFRD3knyw
/fh+Z1hVrqHjyl/i/si9Y7E+zOHzv3/2pVN+0PxDMJqbDfI+EWFRcAEO2K76hwji
NZjgn7IBxrKxYcROxlcLe8DyAHXHAR5xjSi7lH5Uql+k4EYwAf8KV+F9SSSsqaWj
c1NeXCNOvYkUP02bDScvUN77NwXy5nFP/wkOE3z2nIEhjAQXFVgS5WS93VzxqT7g
ZWN/4dPPgQZQ8FQWNykGh0S6BJEhD7ZjpkV3BNiF+F/VSUAEA3jk9AIEZnKz/cfF
HWkQWPOwjPQT9YGDL9811ZjABWHQESICEfBE/mtcnui2bf9mKdLlOOx6jd2H2Zdn
bXzvNvPFZfUGDXMbpeSHW1b+PBJgHHwzdSyZhNmXLhDP0tlCBlRq7KrzyH3SDO/p
QyLJ5kiA8V7rmuk41kiTKGY9IKl9mZFjNxHwt1kK9P/eTi05Oz+JecTxSIxW0Wii
h/kZi7jMS04Hi7E9lKLtaOTJyWIHCdBE1qFdRIW34gKkAAr2UCwxx5T6LiIiQch9
tV3BmpCjJOpfAGGw/QawalGBlZg88nwaAkjVNR+O3lLgYBHAQZM9+TPPCJPdLPLW
k9NYZ4yhhJec1yMIwjHTvuYWg40lEPlA89u5R6tEVlJ8bKavf7pabxEFVYtHCnmO
suWDpMnLM0/YWk7N3c4iDXGAQXjPseYUy4hDgnb4hjC0yrF838+YM0RB/GNcGbM8
Hpsr3nCD4kJEn5+k7d6u9EK/930OMMvEpyPyL5ccpRBAs22el4i/u/3nLOEHeASg
djtOyPzrXBBsj7Nch6sqBPfVsIfWhKuc5iv1EiKt38AHCWnNfyKhI0FTGfGeChwx
KtcKWcchXf16h2xQT3oozUuSwGcROH2ZtKdaJ607TynaiyzSZwqwepgKrG7RazQO
6d0LU0X9W+sNmkprJOKdwbA770kpdCHLgbg34UD8+ywt3/ZSAAJhsQEThx/z9rTT
cedywJP0fDIg7vGqj+JDFVvbBdEwlQqPQr0/cmQUsjbKd0tKkzZnSQGfkvqSSLyV
Pj3XDAPhYTfsqKWT/EDKMVN57buGULR7tYvbXNflnTmohU7hpENu2niI7dtjf3y9
Uf16rhYMyOULFVS1UVSZo97C+H9QqRnq1kinI1P/PTGcsQkR6GdFckG2YN+5okKp
BRil1Q0wKrJxttWTl4WvJJ6S/vR1R9L4UtbeGfh/5/r4vzVaqcxRdBJkX8ulI3ZN
5/I81MrPUbKfzRSRE5TDyve3MvWN/5QQejeQmXzrK+W2rANdWYVydLsOhtRwLgIB
hGNqvCz4MqE6dTXzE+fYSuAjtm7igw8Cfr9zv5j9g1uPdnrgsWS5JdERFvJJsFyu
Z8hEcBCsJL6vNUbGsYBvWs1d5wr6bpHOt7PHrJgj0QtYfaSlqrC6zIsQxTCOY78H
oFcd6fPwrG8LcfR6mrLHlLly4SpmtSEQn9L3u830rLBlZ5bClgYfRGIHEtgGh6FI
ceU5WtdMQ/r1fJL5cdw9HWmwqDjmKsyXvud/xQ6nEaEjVyV24LKJT240wnUrbvxW
eHnka0kdFY3LkeiNXotdZgh1a2gmQsFFnT4KFhHitaNZXxlY+J+Xt4iAcZa9BUX9
KnymQPuw31izMnp5SSI23eQK1bf6tvDtlWbxTb5MjrXe8h11qNlFj4HhUR+l4bjg
xk82HNOmwp7DNOd3jmt39YkE9vUzEbPY55I/l04ofcqUOngMjlUOxWVdTRQIxb7+
WGaecICygO/yD7gA+Z4v1sUq/A9i0ManvevVGOzdXjX8P/MDkNrNBJFAoNv+FkJs
8kR83kjFCMkrc98Gao+xo4qqPj1iChh10WJwPpjOGg7Ob+9A8Uo44Q8JoL77dDil
PzTbjq3yV39wuFBsTEy6vuxhsWguA7rA2bn8W5c5L2/7F4SpcVm7Xm5lS8uQsvTE
4gjwmv1VRtZ/QYFwMeZ+At3W7FsyPJEJQ/85ylcuw6FL9N6gSTQXSworyGbLatVh
nTcMDUj9vrA48dFi1Sp1QgbKEMrOKo3I1J0Cmbev3mKbnuoBmGKj2JPy1oNvvmzb
UEcHCgsnUeoMK6oE6pmeZSLtljmmsRxgCr6eQ/gUhaWqYzMYqngNrWwuf1sJLTQf
oMBdDT4sMm7FxLL7vHOS3PBGWuQTN71/bP0iuJ1I3lbWgxuOx7VkLL5Ex8BUWqN+
oVhTOwivdB0L0B2K4RRsmjGVaXvj6tD4A5XsskVwxls+PfmhzR04iXzs97dpZ6xP
xRYgd06BuswIRvKpaRNclRN/e1iZ22lJ/INkufz/5W/RDn75WC1q9QpsY2HvdXFb
ihpVgdcGZxTkkN+5YUsrOuJ9kFt9vvhxeOfuWzSkGPQhrsqfi51rF+vDQpMBpJmU
X92yWwKfNxOWRMFxkTUAQ5O8gIps/IeUUSnM469sGcBeki01Ni79ftuUB4x4c4hK
TdrpRoN2sFbRRqJipTqsow6mM2tdNZ3eDfsf5k/UPP731JRB5ddANqtUlhOiCiH3
05Bf+qmiPlL1o+JhSBF4C06jPrAK6gjDxif0OMBBVQ5XZZabVmT45GJqq3U7lf8N
Zspkdj5SWoFQnPH8ezZAOKRzmkkjEyJG2OcIa/FtAcYWa4N/tV/gHYgt5s622wO0
yMFBACY+R3ujnyqgRYsgyXBzjmUe/a9exAb09CachLBaRdYIEF2+nY0mAoKmsuVa
of1GJH4ieDWmOVvL6tWbCJZQ0c0An99161A3mUk/eLVyQOTM5JwRQ/t3mJdqc1kn
LqyqS34/xsaP0NZzZJ/29r0ffHI+02P93eSF/gDkr4dorJLU3vmgWWe+nCHVDO81
DKo4cHOra1oJveB02FemEapAoiKeFXymIRiB6EVSplN1J43GqTY2Tu7OeOOaJc0B
TwRp2LlnDPf5jWG18OjdLhepa05YYHMrS4n2gRkuDivKGPiwfCaI1zMwSi/wV7G/
sXZrIvt+3gEMdwfKTx5ayCJF6WstCkpfsOnLegKYtXAax5mFkfMTNPrZ4T4AbsIW
RgGccYeXhoj5NcUSEc/ntcfzP2rtThchX+O8SCmQu+pFtQVzwgd11JK/hwpYJXXu
Nlka0FU5QpoXu5k++8BLmPVC1wUGlkfpeEqSS9bHZEBngzvu7A3VJp41/6t6Ivgh
AYpa9XY5Y0jHHkDo7Y2IUYynNCbh9pzRxkYSShDMVZLk+xAPyFJcG+MH3Xn3GfjJ
QabtorsNCM5R4aAFhow3pAenaFLyWdt2/uGJSFjIV0B8CeIxVgODNH3QpSjMH+W9
HHEyK+h8NMCBZQIrXai+uaRmo7xCkbkIasEGP+kvFoe2Csqrhdyj4UwjJ/XIKk4Q
Z30sK5wK8nrFDrENBP6+7y3k5HNoCWK4KoWoEsoSvMehSs7Ze449P7HAXCoDjr4x
ITmM7YJLvP8YZZCOS1bczduyfIwTkJTqv0KBigoua6svob94TfIhF/tNdngg+qBW
BO4A5TughXxVQP+GaC2OnqmkX20rO24Bf2iVlvRR9jy2M5H+5Pe1WHhpDZrHM2ZX
bRumtGnZEaGjw8VljJZTG7ukUTq7Tq4SGVC40YuU3rgrFhhEAFtpv8chGL2E1TlB
4p0UpWwx0sh2emHpymlw+q1LkuLiux4Hw1mlUiV+zefiFLuyyNjv9MuIkHrFokg6
38/GCvkiyfNmQLAADK5La4wD84UVdEMPD5LTyJK3mWm9ggHB2OHp/5qMS1ZZB0Yn
C/1c+FBJOVlOktwMJN8gsTd0fhLsP95WPKvBsQ4JQJuXgICCGJ5zicYKdSgShakP
Gz8icAOYeHXx5Ih9dnud2dvN6cVXe8AmQXpdPscQ0yRkJo/pVM7La1WuZ5pBzBuw
fF/gwkNUWNN3mEnVyAwOSyQJAmj8hU2+zd2GbbmdtTibIiU95mBqeHWqyaQjRh78
F62Imgc/Hi1wlq/NzhClQqsfjoCODdaBt73oPMUIcGMdr4THVElezSdu8R4LBfug
bLM7gcefY/VURW2AH86ItE+v2DegOSuy+0YXuhojAuLFXxZ7xYZlVFjERbe1I77G
6AhZ0DE7WeKvadczC+M7dRnsdjOLKpL5a9KNfniSdnKAOSuBBkZN81tATAQRXBPG
NKbIGvOjoSQ4n6a08vXWjy+bgsKZpIrqItrI6VcEAIXDAfi++LGvHx38tb4LUa3J
x9nJ7NDEqFn05fXVXZBN0wkipw2xi/G2J+5knCM9mWDDBqqdWjU87t3D9Rb09RAG
qZ4mLVhHB8NDYtsgc1gmvsoAH2PY/Vygcu/j7j7bmyFvBPjxuYAZLlbGwvszfy87
1pdF1bCrudPlCWCTyrE4nTi8BYcXZlDvZYIBynqvw5OUPOnCH1K5swahGq5ltZsU
6d2WM0j2OY32XF/fkc5LtslvkjQht3vXf5MUTH/2fUtVWsjD856d4iqo+Krm/ZIa
sJeIwpu4t/E3oONrhItL8rZx393fDW1sQvZMM0cA2yw5RHzT0H4fU7p2XBcejt/d
wmvOoIolCOoZWnGDQdJSYRCS4bC893wARs0kVjj0h9lk5tSH1ob8HA+AjkMTA+eM
3B/Y+0QEznD3ZcmWbosv4IwVVsjdrWvUTbkMLypvxaeuOALn/XROs7wpb6tbNJiX
Vwf2746w5Oen0TdymkrQuvRCQM1FLcG/dxxJMUMn0qN3b6lzdgMrLQ617lz0CrFB
PCxLMSFcXwEJu1LE2It/dMMB5BNfTApJ8W9BsjRTH8Wdw242SQHcDZhbuCWHWnzi
/kDydOivfL8anJiHZv5nkfmtHuEuQyfbenYr/EzU38LfHkRFhouCOMBP6PLPnMDy
2Ktu3OOJaplcNj92r13mMZHxUVfsyIhfzdI/kTOlt/AxTn7t7KVPS7MRlM+5TpmA
JVxWCyvi5+liWIo0WnL+9mJwybuDa6sor/fk+9/CQybAXeGdw86Mh35skV7digzy
gBdGhLzIiS1QHUr448n92Mz2p1jPoV+jMCz5+UMkckeozrZ/DvrOvuZ5fPDgRZ/U
WwYAEHrsrA2NjrgRnf9sCgFBC/MGQeIyOytktQ8poCZ7ZKZrHul8mz9jhiDbvMGr
OhC1t9s3BFmssS5AKcIRz75Bay58Emlwc9y6ZNEeXGlPe0M/GV/hHPrB3OekwmSt
1x6GB90i5vJI8u/HgxKdfGR4+ZldpiYTiCuf6Lx5wIdF9AlRPQczPWuIsxnrpZtL
7vrHRIpji/V53nVA5TDdxZ4GuJruwcmdyL5Z8mhgHJyAAVbbdcVB1RAXFsj8Ed2b
2EROq70NHXxDM5qIyTtcmw01NiK5aQbLcgVHQ8KcWEz4RofXJv5zm8n57eQ718Zy
WrnHC4FkQQunipMT1s1wAnSrr/1rrVotd1hKVl15//RdkiNT398BDkwsGg2FaFhw
GRLHeiXaJE9qd9OQMzSS4XSk1/bS0cM3yiDNzWc2WubCbz7HRwdkcLXkcHIwKsRC
NiOQonuyOmxee6+7B9VjbMrWE0JVou5sNq7fu+/yAD2KMPDoJtlVnHfc6LzFbgWg
4CkkRHnPxQt9XVOkedzB/UrqfUXyY02kzyLTV1D6TrWmwXTc5ZXzsPglLKcKzT00
z9fUCj5EDoEQP1FN+3//rzdsgsljzykVBXSQcMesd4yvUC8xewbbkzxi8iK1sZ5u
EvyQ5djwvJNfKiDkIEVl8iZddV5MyLs5jBAHGL1FWXtQy5cFtZoo+4yEkBn6wSjv
JZk0nBDoMf210nEo56qJ7c7mhuwhFcugAva4WM20gwvMmAXpM4i67FIUZVz/6c6T
vhApX5QEhpAtwmSE3ZcCpf7XpE8z80FcYzc2cRIRwJn+F2prZ5wN1Y6AHrzOsJ0r
LYIRR+JIGcFyRC16QbpPKN/cBJDZbcjcbI4JqOm61hSx+VCzEEwvonOQddsg/Qvk
/FdfebNLq3hQQxyfgdI+A8uWqK5Yase+EV0vmddNKGeGGdZD577sDOLcyhpfdoJ9
tO1YYgmiMgSk5mlnKhC2TXejJ3tunmGbmv3cMhlsnXBEvLNLY2mGLR9+6rKYjmvU
70E3FECHEaCJixqZsKthv2zNz2+Ehx8wiRUhXmnOLEhcztEWsLF31HyI40uKl9ZG
Qg2sgWntF7dQG51QxwTJ2q+nFT8L2i5dejGoZK/UhgEO2Bg5eebE6l9cpkS09Irt
0ceumsLLORzRwV3F7wbubpQj6V/NfJNcIIACz73mMHXdC4X0Z2gaAzZv+Bir/i2E
swJsGzuJ3Jhz5K71iKD4HsSQe+G6m1fD9g3egygsKaFYg+L1lR1SYyDs+cTZnFUw
PZCmwRlFyyqr7bj55spt8AdpVaYBt2FPgI6xnIdsnjd0x90muuVszlzVbkIk87y4
bJlhCGZZS16PRm03bAGypew9JjtAq0ZAD/JUFHLrpv9anbWwqHd4mh9GtQtngu75
CTHQoaSHx7Jc9QY11DFeGcRg3+ZMRvFmKc6gL6rAGF7pFx1iEJbQ/HNA1oReJVCb
Syff2LiEgz3sY5Ru+SHILlt8PRcRjCx7fVqOZ9k1xjbC3DlCMTYUfz/YXjJ8EaL/
65xeeqoiEATy1ZwVjvRKXAfS6HahVGqbf+t2UbgJ43I9gYRBHClAJOC6du7pLA0A
zxP47MjZrcUYoRCDSexCA/8s7Ez+gKnrgTipJjMlrxs4Vah25e5H6uJdZI0M0nSi
bkeke3ZL34A8i150nne5ObcmzpTRJ69Y/swT55DOdPoSNE8Keib0EnLdbfxJK3Sm
Oase1d9znE5LXZr/RdonvNf6LNZf6JU7aKxIIpPFJ4QFKrf+SrkovC/QqjjaOrKP
W83oiKqQ19rYYLTcOjHLokRNO4Fn7d6pVLcl9XVzlYm+nH+Td5tOT/oMJuRyy8zX
SbusVKrCW9FJzF3hL+nIFxVnb9aOsrFgUsWF9ZFqIv8Gt6tA8cB6GKFwR5aGRuLo
OxjlCx6bJ+yAF0EJ6W7aHK4d3nXYwU19180DIrUQSVeSJCM4KlTsAUhweEkc+Vzq
3feLPpWzFLqYctpUNlHxB4r8fUIRAZttrwR4DAL24+hxV+M93cr8LFnfvQDXJTsA
joUvtDNaM0LAVCy+/im16bl/1q7M6KYd/tBhjBsWVeL7+KwwsHVWy8kt2wPdPnTZ
Hwz4WqBvIqYAJxpQJYjBZV40aRNdUk/7NQcn93Ej6r625cJYEuzTgAijiA1VLHpj
F15VhQ9JDfQqriFcuGUv8luaCdXrmi8iUvc2YrQFvdn4CtGZn6TsARaK7zxzT+wP
ePAEQzQov+GhxTWSHcsAi1XFf8HkByQVPCpogEAXqxEeKxotMZYNQljdq6HqgGuC
b4TA1QyTeUyj9Lmnwz3r5W0j0ZYno+y2s5NQXznUEsvmVrxK2Bu5RV5dSxULilbl
cDhPquY7K+3DOWKiWdsaWGiuNNh2wyKueczUA2xbBsWj1OPNCo5H/tiESRPL2TpH
ylYiJK7c7iwcruWU92pFSgYg2N8s5KMlHh1kMEDgTlirYPZT6u2l8Z3oQrRp3sJI
hekHT2Lcx5AS0TR7arSTIFQYlfY84xrWQDH7DJ9J2TWZGGcQOja8KDz5c7CnUJG8
qq/O2MwLJEgTHdd2C++deiulbIzk+gnAqZvPn5WwiqIzSpeeABAjOtka6XUs08mC
OYqgdTqtuq/eyJ8ai+OleuXuCjdW9mT37ja2Szdp4GVTwzGAJsvB+GSBH5coGZAb
frWvo/IXVTenNk8/cB/oCgERW4oT6Dk6pgfyfVNsnnQDZz6A+NwOlzL/eFNHUq5U
USKwmdEi7GS/fuXJuU3OdWVpOG+/kFgbe7B8c8Hrabg0XXRkKKdku1n8PEpsVkeZ
H5YZ5YBaho7t+854GqymXQaP8/H+xltRQImlYNrZKqo6CeQkY6SFnx5IoH7z4PsL
X+nhExVD+IRoa4XJk/2iHUvRb1uhmioYxiHDMehSeaJdIv2dplNDHKfvzRbUEXgm
qTPuq4t2dhaA4mtOyjpUxsOGsGTj2yyU9PjK/IXN7Tvd20U4tmL7tAhjUKvJ+qhB
A1w3BfxLwJPvM4+8QrEWXKTmyx0Mh4gPbeu8B0Oll2I6wbCXHW6Q6ZjFhwEcLadp
KYnKXg1hfu9204KtHjV8J/MgSKqvc88Km7yRarJLATUVswnTMmYVlMwaBGoqDJno
4ZyKae/0BBvaLj8hgcAdetQqf8rgBgKl8KrS0YoSlAUlVEt471mJ+ynavVB306Rt
jj9298DulMUlvB3VHhHhELL3xcgK/uW0PBg8Y2DfJwEJYxx8+P2kAyTNcrMtMwQI
4TdncugdARq9THmHFNcMSPmTZcZfe2c27P8E3TUTpY3XyILSfQCvTTCiQLTMJwNY
KRI1R+15A6560CdPThfZvh16pVr3oeIkbJLQLx9bVdyMYJctBOw8Rqug9VE1iWur
DpsSYUxjU+3jC7oamAfwWPrD8IBSaVIeFERUPedCOIG1LaiBgILASzpz5nivT2hs
rGlE2/WiaS/CtlkCHNId3/d1pVApbWMsw+2AzjZb67VWFvaFjS0DyIhm0QcFb0rW
z9hUsq702Nty6+3RJ/M+bKaDCwL3cYWVoYnW70zTMdTxt3r0ASXOm3R+4HPqDCgN
EuBZaZEnhgyUf/+v6SVGOMxziLnSM3qobWsoq/FvLrCt6M+OJdX6XKukrVCLtiHu
ANLWueRkOghgTjVnNBRPVhCoS1e/JI/ZQgvp6xPd0Z59wr4pxghfHeNxeqppp+Rc
QPa1Zrrk+NuPNbmsTvZDJ8GyfMTQcCp8URGgvdUkl5p5AbF4XDURkoC2Uqbw7PKo
FNtZ+ERjFn9Jb0UNhceuh5vNImvQSfdl1shRPtM2qFXpG+OqKpqHtGsFx4MD2I71
32I1wqp6bf+YQDbGUTK+hncWpfXrorbVoD+lAFCX8/ey0dH9lAak59RRkCqsKB47
kANXH04t+mGCrULXapKe7RCagn1Z2AWMdkY8c7K0I6e6oK0wy/K3Nk9NTnaNCUaD
cLeOn4FDFcyKY2tW51ZO3Ha8BJo3InjGD6N5o8CeDisVVeIDYHRtXm1n8WP9kKVQ
j8ixebUONmhp/mBxWXtoEyEiP2OsIpWo8Nb29nNTOriWpmF98FS5s/TzJaABIZyW
iGJEu0T6kf2Ml6R0UmNcaDZ4BNCn1sotWzX8tPpJ3j2UKTOe2c6ffzBX6AbzTA2I
VIjbr1i8QYOs6Pskxhb/TPtlW6aDlJKmq8gKbjlyaFTEkuUEkeE5Egnfpl1fNG8Q
GIVTUXITVplh99rmu9zLcUGzI0l2ZN1UrJtcw8+KNqBYW7eZjDX0TOAxTyY2sCmt
IKvQVsYpasG+cxxgsn5y2Y7LKNIbWNLZivBj585qneUHH+J47UHThJyrTp7bxcDJ
qhdOa4Qw8ZE+Ue6beUWxnOE0YWuXLbrQhHa2nliZPOYN4JSf0eZ/hH6g5W1/Nobr
RS14dQtoJt+Zi0GzJZaoNwMc7vrjxq8nqST3zi1692a1lWNFhJqp0Pg2eAJtH7wC
9hKJmtu5UI1qmaFn7qbKC4VlCQsHro3UlgcrwlyOxllTyUaIu4wX677E/hDqYPpG
hMj6v6BL/nBQWZ54kHB7EkmCB8j+5CF11tAJFf6kPr0LFt1IbaqXLpWcixHAYxGT
iEVjqJhNHXbFxhOy0Dhk5wATRIi1yhaDvWmeriS5/8ceykC2NQbOiNfQ7yYU16oh
jO/ZLntHMa4ny8tarXHvkxLuH57acSFboQ8LLXHm77vRgeW4ruoWQxuhOGARS4vW
uS2irLdzkZkjJqm1YUZGKJd8XQBght590eOyn69fTY8UKmqZV+Opoyvsoiey16z7
62L9WYBPR06RbrKirucgSqTkvldb4DGZ1YPQQ/y1YOtxBPdzH4NN9Jzixi4PpEGA
SWRWRENZJzzBJmtMUgido/dJ6dEpI9sMTKjP2U1c7GJVy+as3BYcuM04NTv5DbSm
hH8hoSvA1LvCV+pt7J72EHu43wbYBFrF+KJJT2eSz7lSXku842A33fqIAVPYYbxw
NGjzgwg++FLrletD+xc3QJZyhve+M0QGA3vyP0iqrK4CKnwfyF0lWPqT1P9gp/vM
huRy9sgCBj+tsjoQoqREjQcHJ53dy60WeL9N8zziO0UGwzhMVVEBNBuTMSa28gkx
rVQcO++U6rnxUfmQDQ4dX2DJFZ+ZyvNPa0FrvXGegRyZl0p1Al6KCg9U0l67mwzY
++MUU3RIfmz57yv8WSpsQQQTANTNwAkP1S+gBvclR6Nm+onpVnOibKxZ2JJ+c2PI
Cr+nfjDzchlIkSFiMKO5gJUVdgEfc4qfmWW4wRX4XhsctIDteLCviSLpYJ2OkkP5
hESugm4G42ZxHEED5AjdP6WKa9ylBKHnJ0ZsTK2wtHHpk40A0QYZHSSTR2jbIkmy
aXMVZeiu1tahOy8/AiR1no+fj5rf9trp7g/zyNGv5BBacM8A8IRtpmpu5BBmuC/7
9dJ+mZxssdZqnl066mMiV9VidDEdCTDP3/E4zh2tMB+/v76qbUH3ZcnZYCwKYofz
v3PzuugiGfOoMFoI1J7qzhIRjBsftQr+ZYcRBELx1B5B2XAD53b1idRtvBButORw
lO9yDJiAh+vrb6UHJBpBl2f1flndN2i+aovNC0GSflTng8ThTDcZ1gVMSKzCHNW6
WoDjhvlM0Itdi1SMSLln8eq/OnLq/HM23Q+BnDYC77il6qEQNc4eNRNobwCAaPUz
ZFdMuUGD18eSR7Scpg4rLDlwiMWe+1ML6nNBUKkF4Gg8GIEp87lsqofMqaXNSJcY
zD3MaQ0tS/XQEPimgggYfAjftFTTTH2G5/5nvzK33hS2pH+L8bGvuj5/PCX3EdFP
rHFGQ4A46HM6h8zMsk3VxJ47bQag2sgDLNUK4C+AKKzxupXn9TEQKUHcRz9ARKqk
ndVJTIHILeuTCug7tueKxLiy+0WUhQqxxtsqiOXxWZOe3+1Cqex7QmKgN5Nbpc4O
KOv33aLfCrJzJ/XP4Zd5NOfJTL7A3QzRFtCUV/b0T3VlZMFOgz62Q+OUkDTfMVvl
A7o4LD+DE24eSnaeVm5nv2UgMXZu0QboM6vjyA2HbE4BOF71kw6JsLy6k2vg4c7P
DRm8cXiH4NIHkAfLLI97LdKfx1zFVvTdSRMlnroBgXln85A530WOgDVWzKNVk/09
r7CbY7wjH/D/KPB1oK0lsQPOM0IZbIU5LSSPQDUqUP+zyFfWqEU/egVgyZpzZP0d
WeBjwvd46Aa3M9zyRKq6LXFAAaQ8e0f/86LYIzlCPoZ3mZ+rRVFe4w6yxVykwThT
Ys8FYdBexS5iPKvim45DzMtxVGtDy7Z4Yj3rPBFKh4TItg2bgqd4xhXcuIrdx9nM
0Jq8s4SoOi4oD0286pkumFUx2AiUnvcMas7dPeJfjp/ZAimq3oDnemEHUbe0pjUP
H3QH+/XUILPyPFIAu8UJoV9Ft3OPFx2RziOqClGiI+yhDYWEOudaXEEYDl/v0Sea
4ayXxDx4ZrAfLXzX6s1eDLUO7oB6PLifd9KZYRwcSdVoqZvNVHEp5DSNwVgPkUAi
4xvBsMFoGKxYigmnZvm8hEI+QdAezSbedApUAednO+RFLkKJNwsKOXOo6Y2/h3uN
De/gw1DdzSKf2F3n4ozlvGY8AHMzJBf9YDsOZ36cuom6FC9FLVqeH0JIcfeNj9EO
iSnYUx2YS1xoIfoqgZ1a3wHLgSUI9+C7SSCZ8VdIOZ19fwJ0XL27fuZFPzA1dFYT
PzaVLo48L/HbXS+nwqpMxIpUkFRdqs/0t6v5lbhrLl6M8+5ZpMpkHRPfcRvejt3+
j+kUKPwpj+//I5cFR7jNP9yOk58uNZIrUgXRRxGx11VBvCbGX6EfVxIFY/48eqay
TuV5b4YYnINZYsGnrZZxgaiJgebagIRh8+WkaCXu43nAmV8Qc1EsjdyXREtDlKs4
xGwwxg/tUrdQmmizRikAA+iyKKjiODCTUHr1Si+he6gGXm4Xhc3qVPAA33tqSH4q
NQVdmrtS4ccmwbB4PbRJuNqv4zfPayP8skZXZlumGRvYcTILJxLaP5kit/22FYhS
yxUuo21gdr+ukS9oIp8n/47xtHBiCQlIuaSVAOlaLd9358ABiNsxr+9b1TAOkQin
Rjb8DnFTYQhFpB4tBMBa0K3Fr+EMnbEwGGY3wfwtzG++Ab11G6V9+DP/Pv6Fi4bt
yLFqzFvgKw8jGq63JG79SX+OT7OKrGxzaLWuTcT19nELD6yeJE79DPV4XMtOCAXV
vpFCISM8yfJaDul0YLmK/+LAbaT823j2ognp+ex+4yS3J0yNi79jm9LdZHS3il1B
B7Nj7Nje2qIWXCPI+Z/pm+tJYbhgjT7nhAJ6Di9Kck/OpMJfhrGEkO1Sowb7m/p+
coxfK6n2W7rGl8SrVdcz+iUehGJ5mBHPxErw24AOe7Ch8Z+oaIwo/N9K4DJENi1+
fjCKOb11ahWWKlSlYhccMzRZVmlQSvQdTKLywX0aGvWYQ1DXmsnC4fCJ2/tmqPvl
Zs+6I0IkfKng74zM9eOpLknQz4NTDmliSEZevx9bQoEjnKCsi+ij5XPOcuvij2Nd
VC7PWXYHr6XSgamiVmPRMSS+eMhpzlm0SH2J/ZkJEjRKdNOBzCeqTIENXNVayohH
GrKFkUERe+RgMBw332g61R+fMtuHLv7ZGW798t1tkfNyaUfg6JAdpWCrfDdInOi0
HUiHdhQ+C5cP/11bbRlwjDTknIrnwljVx9FvyUL7QQ3/0JH+S8WygonHedlsOptl
DP8HinrVq79dz5wZofljcMqWTO4agm6Fd9LWhz3xl/K43d1bapOjjM0mkMFOm1xv
ODdG49+2M7VTU2KlbP24jtTDkZQyRoZ2Mp8JcxGfrD+b0ZhGOOKR/awqjE8jOSAm
wyxb68nMn9UoY98NZlJO4DLNF/qaxDPzLwjE7IgA3NWu1jZu9QcNFxaAT8rskGJL
hG5iokouSW/cHnnKLc/UDgI5/Dtgnp6W5TsvM1zt5JhJNvpUo5B8OPIsIFNOe+Dg
in2xzNXLTJGzeT1f+5ve/Sm4wqZ4aRJIS8XvBMVpuZ3zRMgcckxcvdeUO+iz9cYm
bIOEoBtuc6c64Yf7lpxraglPZvWxRd9tHzK+mP8S6eXFoACPsfl/U4lG6YzLQijU
nK3kV8hb5J0J1J1HyZ6bJgyCOlDVFj+c3GOhdDcH940WdMthbjPUb6LnhANLKPYw
kbw70aG6XRLBjscTwyuMja6AEybZOPE2UIRb6JNLYjIPKv6P7Y0kg1jwS5OqxXwg
N+pct6ZGFzLgiE7jZ5oREHfm7T8pazK1SZbozae+vHq7T2Aj/kWw8BICqXhHzQxV
jSTI0ESvl8quEU7IeCozOPy0MnMsHiHq36pfQg7N4XAuZXd1ipe+j3Cwt0WO8qHY
ECbg62fr4VK7K4WqhTXRxj7Gckq/G/J/WI/RsavqeR+RuaOz9CZ22SSQoRJL41uq
TblGt2TcWkXBM5fCQ47qGoUjsIZNQqHHWcNlW20MlXxcJz9164MijgB/8WOpl878
F7gcfxqI94z2Zoba/Qda8tfqNsofP3RFXG9v6HbNUq+W4ot7Mu1x/BiY+0uNAqhY
ryqkFRd8zFqoiIh4MGVA2aSczaYW9UTUVt5tJsWIXiId/YxJ5ufM9ibKdm05fkxL
ACv/daIraNDrSitc1B5wNCDgceHSdRynNDp8yVuDsz8NY38L5LHt2vz5mOANQDiw
6u6fKw0tYanidBtob1sykzplXDUn4Zzoi1MXG6mwCAeYGdUrYEO8VqFTiXgW5DYq
`protect END_PROTECTED