-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
SadRbdsVk83SWJqVXpzo66WTmEDfZ9N+LtFKOz1SwUwKJWAumRYK8QLEHF3nKF/J
aMkgE7rjwgAAZI4hEtUFJmrgPgzVty0RnJnDmgUzJawTZBX/tZSDQDemsNgQx2oM
ZHGemGxX5bDPxpNPRuLzkWti4a4uviqVQuVZsLgNpPVztrlcvtPCfw==
--pragma protect end_key_block
--pragma protect digest_block
9q996sf33O5BkmDW7y1U7TsF2pQ=
--pragma protect end_digest_block
--pragma protect data_block
1ZRT06UEjxVzOPUa0iOdpN1NIXxFfkEsn7onQLMt+y2q2+bd9+WxtmAfsXc7rJDt
CMTQIXaxXi5HbMf4Zo3WvWA3XrXqNkfrLDLwrOiJTfaZ8q/KDDsxtZPxk/0N7RWb
HLjuP427yIAoJnQzSLo8Pps/o5dvgA7izDod2LOOXugKUvzDL8YhFvF06ZgYzaIt
A8yRbKStD0dpD5aQVWNw1o4xcQ3YKDCzpfaqJ0IjMwVuHyo7S0E6IjrdORi89D79
gtF6YAztJXadZyU92O0GSck7BYF7kmxW7qNgEQflGAbjlVrdtm8D/wGEUPbGwrSL
P8glDmjhWK0dqjx7JRX03QuluJieFNnkhtClLq8D5iSYlCAslMWICHrJAACxtnGX
x8d0Ex+1bVaLicOmBQvwrT2N74PUBHDrSHMxlM0+aBQX9iEExEloBWyhSn/NLJ72
wueqJboGSq4BqveTGHnfjCml9yNhiirnX2Il/a3h/QxfpfxBqAJ4hyoTwzQiLpKz
bCq25VMzG6PTJSObpEeSutwJ8cwrfd61oqmpE/+hrnUO3vYV8xzdUTCe5pXxUNND
ze5o/219qcyWQ0r4rvh8AJ+hCuSjn7Kt0uhCA1PADTgxIvvcg7wd5OZSdqfFQ3Lv
3snYPsKDbhpMQlHzn5bbVFr7JyUq5QBNvOBXibKrtvCnMIsu9a++vdq+E38GaSgD
aJO5iMRjL1x8ZlS9a9LHlg/Je3omqUybyD/3i1xoOdRSWWJ5M+u7LsypVSdgfVUl
I+X3+Jz7mtFrcjUhKOqFbmDDug6X01r9CNNEJgQpPXJVK6/G+9mV4vI1ThCsLmnx
+kZHRzQw/aTO+5m4px4wUAvNgpg704g3jYvIGVTzPKiySSof5RDemqbL9mNpYgAk
pOuAb29Tue9dm9ywDNF6eGgJeCGGskDf5PqOGVITa+u65ImB5umxH6Sm6ZjW+ONy
LJcABQMB42a2c748Vft+/DA+0NBqcO+J7D4lQvznObgkSlqM9+buVrSPBIeGRW9n
2Sv43yp1dmiKvP7pIHmoxed4tSuhVr8n6BQi3fQkEfAQqFIv/3S6W/IklW2OtrMT
+2fWp3mVk/P/3f8y7Qzf/8aCLLE5TVLL3naF19kqOTHDqxJYe9z79Bkl6xf+USDN
nYt4+WgW3ShwizLxPN7js7qrSUeKpouvP3yHNz2Pvqo3YezwLF1wwCEYBbttGxe7
fzThVP37P7ZPoi8drjX0LgTQBNhE4QNvQFA25ONlrTH0Rb8VJ49RIUvtqh9/CnAX
YtBWF7QGOWXemZhZ9JCt8iq5YLduVv2b7WEfnKckkz55SRlXLm0B2JjPIWVHhvpl
bg5BlDMY+LSyAnDsNjdaXlYoJsrODbk2bSdJ8CsEKitXW/lIhi/GdQGZalhE2nmd
PrHMfkSBrKvc6ttBEBjXhYbG/1Ca0hY1RYVHQS975jN0x9WUe4tg/i106n25vuYF
zkrROoQ98eSf2RjdQekAMvcpra485gegXkqGdWE2CglugxSY1GTmREDm40lFoFOf
LC1OjpXYrCWSqxSHS6TS2g7UUOmApgm+kfCZ/2ZBtXYzXNR+gVn9fVfEblRhoiII
ntNXwSfaN8wX/bqv5Ju5+x4hJYCM6L62RdjhjHRTQm3CWQO3Il4M/pXM1QPgJgQ9
oiYMdliFS/xmg5MYUIx192tewc8DLpGsLQhhrz29SVA1B1uWEOIK4BI5CPNzYpJ1
9p3RyHlJLV2sy/wdiwqXN93exkoSzG0TySX5wA7o24J4+aK2g79cDDmal8cM2gL/
wWbKdZrZ4nk4iNTqvLfTyHyVJ+oTnrGONs+zESMDFuoR+s2mqiBKBOw4jIBPRe1G
MtcjQnqN73T8GLFjl3Rdj4KG1eUoiL0GHSZu45xBFw9WeF8n14pUcWoJaQUty9DC
Boo6PIZVNk2VcqNE+7arX16A0Uf54lFPbRsL2cfni42ezZT5ZXXSP+BfJ4zFnOxB
3O0vK4sB44rqjrb8kD3yYAnk27wrEJqdyCNEM4WZ/3U2cbMUZoMbDuGaGWXZ7pbI
W1KDztnrAuVZoNLSBwKun0iUMFfeYTqLss++VuN8FGTYI9hOAmmiutTCtVwLYP9Y
zSbNLOaPz8nAN0wpttbppwN5bGWSNm6I2Poc1JMalewoPek4OF71QP7FALOHML7l
wc0rlnLjOO1O4ofHmFUmxD8wUppuoG1CGJxnFDKRcIiKGDj7ubK25fkcAy42M48X
0CJGcVwCJyXSSBVBE4Bl9U0l1Co2RH8MR/p66qgchP7pRoAR6bZYfYRAJZaVpl7I
2jBnHNH3nzRHOx7yAwmaHe1aKhjgysYAEQ2PiPNoJFad6a1PW2EeawOMj1O9LGto
q+3Nz44FTGLY4yB4utZhEJnRz0InqoVkvCzLvSKwi7iJyJz46bM7e+zebJqxOn8+
NjxNSsEd5wzmx4irSOqElAaQatkFXrJWM2PmiiezFxdaHVZXJ0U9Z1VC8iU8ZhJj
b2EHV1sajH/mFSBm7pNT7VYSBGd615MnkHpBkK2hE0Zk6BDICC7+fGwYro1M3x94
mGvtgV6dwDC/lxeAPNJSts2QqfDmPwMNwTd+0WtLxN4jqK+8aqoDQbl758oPVMen
Y0cyNLexoLvLcWU2Rl/or6HO6n3/jYtSeiE1sfWxO5IhAponcDC9Qq6QRIZTapql
U//Vg2dUX01a748t3bqtx51L9WORi4xEPkr4ojeNM1QxlAbPhkAW3QmTnwKnLB7t
2IRQqJIZzwjN34sndMt8M+6zf5tok4T6h+AjuwQIidXgOXEheXpmikrymdlpDCFG
q+C1tq9swIFE9B4hfQsshan6yll/GhCUJd96ZswhTlyrDysharsBwxUdJMSMEYM1
lT0IBgvKlrKiFaV/d0dX0YkncG736JPu65Bkq8fgE+FI0rhWI2pnrlEXrzYeIFeC
UXS2sfIqq6/1kLDdetUG9B+HcZnTOG3FkYFV0QW/9euPe423C7aZEm0NVVpD6M29
XUpiEUvGSiMOxKShGBsJVrlf0YOVUVto9t4f3d5crJN99tOPnX0LatuAKk/bXVuZ
uo6/gv8SKcjDiin48T6vZSBLW7cwtePFXFC1ZI45BCOQS+wFPeUKEsAN5OXHMsz0
Dwphj67dFX08CuaA2rg/g91trwo02LaqvTP8mmLefZsSaJPdJVKCIZs7WCo2RlO+
Rokx00mjuMT+BionL0bJ97KqLkGmHU4hUws29jFhIODLF8fv6hHiMYkNurSobOp2
U69aMFBR+ejcKjQzozHqT6oWpqWPov3dW8HWApGnoIDavoB5v/0wuWhqoLn2w/fY
kRK0PnwTyuSYz6TF2CtUn/7Va2JN5UkUR2sd24qTb71Jj+u1mY3zVufZBW5Gm6fy
Kw475fbZmg36g+IHOqP69EZjeaziLKaZxHW5FRXEma01lWvF1WEOr05JMZnLlFQo
mz+Bm1y+c6O1rKn9f35o1MUr2Tc4yvtMIht5ySMDxZVPAfiZuE34WG07Trp4diQx
XH8ezAkYJnyZUWC+9Ld8VmTX54l0MRjh/ACXXhr8KzGR6+9kICOWSRXNDKX8q76y
oktG1T1yUyT/spJYLOyh+SI2TfGab8u1+tE9rkeleNMogdWI2J2L2Iffzf9bus7F
eHmgW5ScAk6Pw1cRWudh8VsrmgAAzE2ODAHPppHIHR/00LQpNKLfcoIpYXvBJgFC
bV3f6eseP9BOqGE113LVgAJFaOlQ0CHW6oG3GsmNZ0uvc52sMfLiK6G2fRGQjVta
bQC4qAx8Syh7cjCFBEkxzVQRX6Di4IW9CF5K0OEXpRd4+7SfcF54Sno5Do5/gYKV
yzhCSR/jvI0C2HWkfVHa8srQHMU+QiRL1b3hqE/ZUOPLrFONtlVWGVYNfj28yOnI
JIiKedwChZJJf0IBaBCTSAcuyjaJGZEZTrUjCpYhvGKYxmEOwkJkKNjWO++U6DRg
9JNajgfELOWQ18oyoydx1D3F5KAEhIWYtdlsf7jq9DjZSZ+03WWkHHL7X0TAV1KI
UQi/Dz6ol5as535eVd5exC78UdAKAZAMmHcMTgG9Fvoj2vCMy23iQF8MSGSKR91b
r/tkHbJaPKnqo4hGLUkW2zQdy/RRpq4w56dETmxWIKvylooiNL3EyVTb9DU49WCS
B2gKs+elcl59PQHLrRTlTlEwXz8zD77elCZqnVbMZM71PlUgbbPe/phfqBqJylRd
6gZpAhp/QkPVQxCBImdxSOzio2FHnH5pz4g6SuOtdZjNyeJsw/Q1xRX+oWSHr8eE
d77LU8txjcZmgeIML5yVgyFRaJre63Zr51AHWKPYJ0Q6RXyP3//tSIyJxmrjfIOR
yibgcos3SZRl7FbNkhYqVpl8Qf/afxxe9q4egh0H4XAITl+0FeiES93rObehac3c
Daz8UaspXyywKhkg5e13eE3C5uvaD6NTgJK7nBW9WZso2r4N2hf266aD3hvlLGiH
RiauQ6FNqOPML+P9fVW90iuoyEKnAi6RsGyxG19FFDbBffa3/SmTwwAl2pUyGA1y
BDdKaUWg4LW/a7q6h+pUJ3XI2IE9RbxsH3CqVFCn7GJzgRD0XGe0LDnr/K2PGKHi
PdTWUIoztpIoGxcDmySCreYMMjnCCweh+QSC0xgRvzlPRm5Cqo9s+2P7Zp/v7Khg
Jw5rIbKuxtlL3xwqExeU+NUv+nTQlT8puY8tZGXq5U10N5C9z/FZ462Hz2O76bdk
/KyTcwr4LgS66+OVW7o1GBQCLnwBKJzPB8/ClJsb8YEn1nEFlE5TS44KPqmgYsqU
RcFyNjkxA8jAqHhHC/dJEiWvlApAvv0mDjX5howqdVhkn846QbwDNO2eMAXfDVx+
X+ZmnGhf94L+ii76h3aSqBUs/H4PXTIPO+4RviJZUyZWuW13E5LfCjfPWx1QQjdj
aeOSQLzLC8cfmv6HMoWLdZhwNTtu+ipFlUFE8SdEfivuf1453uLilBxAwVZIWJOp
WTl3BFD2vVIYZkEedZN5NTuJu5vUDK/m2Vg9ZIgIcDciMj3seHXMctJdytwX04/o
AAUSxSJHQQ7i1kz+k/CT7RhYD+/oeB8yc5TQBhBP38OsQbMHCNgEKd8kGSs37xyk
8cPbcnp5X1dlsuk4+0jBjphcjYJ1Vo8cEtQ+ZfndBcjY2WYd4tB5+2hpBacCmwXA
BuYwefLAG+1+4jKhFk1wJ5ya3z4xH40zDHDZPapVcV2OFWpokhU6Qv/BCXbSXnIk
/IZ32319F9hTge36gHxe8RP7Mbxktfkvnie65GGtf08PcZvvmFn1DUFDicaHL/8M
JiNeBWH7bjYr9xf5eCP1PFxK/jadqRyh4+3RxvFe8zMgeb9ovnnx0Gx2huoO7KG0
VBkBtpgVxpXwPyWIvTU1CPpRKpnVcEClR2JDkeq0G1qnCA2z/6xe2EsBQKHenQib
WKKyE97brmu1u25DxY5MW46tngVEyD7BDhXy7G2hxbYKi08PUJHbLF0K4TuZDtMo
Jt/iUVmv84gZAgOtYk36Yy/nxNe4wnEkCXa9/dSRR6qa+oFcORln4XiThojvLZUr
re/2ApPMCuhT72RaK5ouL09Nr8qw7Mcqf+zRw2pbv0Bfyl/msHVy6kJoofA9QMcX
TR/xEbZYL8+vElmLjGHy70Q6UjBto33BkrEwnqu1pr+EhPuymYjrXoK+aYM2QE1N
CCecTd72T4gQYuUJdJs5uBUX5WW+U1x7M7LD2uIC1yifgjqim2+SYUhDq2m9rmyF
M3ph9+hHmuIP+uigh5TmymLSiW4YShithBfVgH24I0YbLMIsmG+iBoOTk6PEyovu
nuDH7J1+lmLx32gNqvAV5dzvxahb6WLPhP+cntGU1r5FBYAZ7ZYHyTccrhM9tqAO
A6C4WKpmn7a/usBiXuV3DS8OhWo/xyBe/In974EF8109iRh+zEd7WWi8798j/LOL
8nytfWa2IuEG5/y3VlbSLyDDfsv0mGH1MS7fkZTTG8vgldUwPn6YUZqfjrRTi/Gh
hKjzsqCdV1EZgTlPPXMGZBuADXxKbabrgpETy5IwrHnVk6plfGwdhoOt/H92HRqt
03tNG553N1fJ28/Zu488Gzib/sfkTvqE9SYvfz051mT+0McGKJG5ZTgfSaoJgxHY
Q/OQMLJsSr2oJzn4vKbTO7srBcsY1zODBAKX22LsuUcKLWmXsJSfm3HNjkgelhjJ
epVNqHx08iRlpXgONYxb6hKbONPjWazenWyMLw7luMrVwQ5E6jaJMPgYcy6WY3gd
hQOwqZLnQmIfZPyyVAn2i3WefWO50SHYzjTkRbwPLkjXjNU85a1hsJVgil5mDNAj
Bw9/62jjHY1WnPCagp5yivExMKEQ2FxgpEUb+yea5FUbehf//XckP3iTSQ1NHAyL
wcOVhC7v0iFzI0ygs0cSbgzVaevLMhzSwCArk94PELIt/N+xxHaLil4rlsEZmquD
m0sztGuRojEqtaf8V5YsyqKS76R3YHAWDBPnkwqOXa8EdAxJhJpjffRH/QffX764
nnQi/kmPu91pi6iAg97in/5dh8c9MDnpwhbvrT0GC2slojpmNRvnZw9S9mbomHcL
iYQMpRbMswY2Lr/PKAwgxFP+fWiizFpZAvuXezS70oDd2Qhg01LiIqUq7TOUSuuK
H3O/OkxIOroOdF5TSJfCX6OwnbwLOPJFv+YxmTYJCzGxaZOlZXxIMfU7fH0qfsqT
9sG2Dk3Ok8jX//SSGQ4SnIatZIeWKfCzqKyGYomDqhiU54R8s+NWOp7cWeBvvUrj
3XxMsWNIHfJ0RsVDHppTWQRWRamzYLdiFwpc5IVf4SpBQZ1wWdB54hNJxvI8SBm/
7e/dq0zcjYqZXAqKhmxKsnou4PW+bSakAx9WIU6PTZwrP3iZq0wXCxIr9+qzcuhI
T3Ry+16a65LGz4HMTovnvONgvQd0ImXrLHe3nsCUhiiwYa4h5o2eGzMn22XEJD4q
h1CYFp3HQSpp7laPxU0+0I0LBdwhrBIfr/EXutMb/kadMsLb/0VFA14ArkIuk06F
Q/tSnFVOGNKv45YXi2Xsp8R2NTB2qYBkwtr2k0phr5oifKK2zt19eh3HlFR6EvU0
GGG4tdxiUoGu2ZOGjs41IMQFP5jR+txqI5x8njb07UQPAmZYUJD4Cs4n/o39Pp1v
7PfPeGloAWlmPTGkqtNEep9NG412v1m0A89dz1Y25FF9o+X1dT5h0kUp0Ek6zXhX
srfrP+biejmvPQuzHlU3eWQqI66llUGJ5Coggw/E02TpsvgQ5Gb1lDqf418gGOTG
zFHSsneMzoT7VOoHClR9kIpxYhT3GfHFp0ZTg3iCU35ZMCFCRZhWJw0WtW9C7GOI
hBCcq0/+MFXOiPtTbh+Z1VdGzAVci6+jr7cV2BjpzJY8Nj3mH+NMnSjEZr7wa4EU
KQHs/v0Xu0uyPgJP1at8qF4aebqcQ0fylqBhqjbpsrAI8OwRjdvgVRP42+gWVSgx
FUNIftIgWeh2Mc7sKLeJsBcFLULhFnc97H9GqaXxaj8oCW/HWnpBh3lGrTVUqQbS
I9x6SXyOt43OgK4cd24V2BLGl1lKzsLckhKgKmwvCJk4TVAOcq4neEq96+HxHFQj
EqnCnKfTIHP5lvCjjggkEiAUA3iA5A25JCTiH4Z4FSzpqp35tAkKhrP/McwCUZKX
Ka5jyp1f6OiLQt8PA/ujMWQxGix65euT+Xb19pt96uUzV5hKXBabnuLJEWJMDmx6
GWW5+pss72Iaw+74ITfMhu6+Yz8XMfjm0G0naWnRzPe/6Nlwl/XRcsMCODRS7Fgz
70taY74Weje61bTqNhGMBKjHGPDlXJQYE7EwHdeUpxXtfaolBRvIhCBaV5GpivI9
jVom9VoSVhYhF/X29xQp7kSgVp7wGMB4K3VZT6UiHW7lDicYcEJrseAC5QJbJCZl
JXfacY7xQR6TvbMPZwv66bk5Yr0T/dmVSQ0GuL1HjZF8WZR/fB2mRHmXZNKbSXON
r37ZEu4H7Lue8fS/T4zll2j0+YQ2fma/o5NwVNU9TpiMyMGedUayBaLqRSY62+oX
veGx09zYSwy68DJjm+G0NKDwYvJvgf5y0b0UPTMBcnuCAmQDeqhiF8WOrUdwHc8M
9X4uTt6SuNXqbmLrVwh0odDrN6Qu6u+GE4pIa1FvUuBwtjCVz+5ydpP5Dve7KtWe
/t2aut4El16ZWI6JVE6dtkXFhWICIMlzRxtbkHlw/vn2Xa0GzCDyL59dwjSEnpYF
9f4SSPMZ0Ykgezo+3MbcHdD6bQIcQu/qLd58J7aC9RqkGSP+AlOD7KGkJZx+LY/x
bXNtsNgJ5X+3dBs6WktloBX1C6eTKXG4Y/1zawr6Va6PincdvWCLHkOx7iwb9rtz
Oj9VOJIMQkB9KmdWWO8pifz945qR1yh5jKQAXidR+c+PccSFr/JjVQ7imX7nmwqE
sqVjKQwtC5STk8aZAy99NKe0uksh/qOBx7cglnRbuMypkAJSNKdfhOmHeU8ElcOE
j7oBDqC8jbD/E5wJ1FmqmghdQFsAl2YJ5/N9XbrXy7BbHQdYHBSxksZL5wKRX+Jo
O6L6P8+yDtsHfbaEywSOu/T8feo3jfBOwH/CGQYyZpXOTZs/WSgsflZX7InQ/slN
FUGlkV2bM9kRBQMcrXW4bAEwBKdWva5p2hdRLtegUof3jhTbbuiyKCUcEoideG8b
mll6SqQzz41paJyzL7KpYNFiiBmH2HvQE/Fnp5LdSheW/ssN76WMea/3GnfxaTmn
JXisR+QYxGsTbCl0qBa13IOC1Br6aQjLlrStl5XNdbJbXZkRevynFVZZRIjdHcSw
/M/8zR5hHWC1WqmGkr0MZ0GS0gq/zL+67jrRb/IKF+30ZZfTmOhSiIQ7TLltr7V3
/l+l09B+D7170YKD7HptFLOZe6lCrNPQ0kX/VO7rTrtCHpTmTeiOr7OqxZFH+zWm
6F60AhY2a+MJJIQhwrPPC+oQPghxshcLSyUFEEykNLp+I4lY3okL+hYInv/bl/6o
YF9lFToaiGDXR4OXrrDuz43bnPVuuAdrSMeA9FSu9jeawgKdykm0tWFb74oh4GXZ
2ndXwJVmNyoXh/FshLobqBd2QUZ8yQzlZYDEOaaJ7Ed28+3ghIxuKruigVUlk7rz
fWLJOnI+n/2Vg/IMjaR+M86JdfBa4zSmbIHYfurD+OZ5SX5T8UzqaW/yu9VuWn18
+LsgZXX1HjQJDlVilidpOENZXW6ldrjpG6dsH21IEH0mXxVmF+WpmhWWsvGaJD6o
cw5KujR2qQ53F94JlpFe373qu74lG20uT1DcEDPu18rtLGpvLq0r0nQfFDVnCc+w
6/mGVy6Pbdt3EAMnWlA/GiiAdTZr+2BzOFlBUutxTnk8OaYebTfcWxkdI2dbFxEG
/o5lKg8n+40EPOq95llJY6zoAqGN91/zbp4w9yYGj1ENcTRdpSX84x5e4WLiCMhT
7UWKcafkOb+xDwR3Xvgo46qElyJBugDli+JcpojVLKIc2AXktlv07qu0fjqybsMw
YWu7ANiwuSPk13PZcrIkL24UP1dmmoAKW9JN+EHxzCBgTirZY4jGzQtWb3BITWGM
LlhuCSbwem0ikm49lSHFsOYiBY7mFH/RQS1C7Ki2IF7LFVzIITWMEDaj7tJmg1oX
3FNn5oFl899LFH77nC+8/Y1EvYfOY5NmqffdRx4GmjIotMHOS5g4w8FToUJS/NnU
pOcXPVUN6lxat2LOTQqaGOtZSF7BirdJi6zURNrbqc4qaTlhydqW+C8ivd2n16ST
gYnjkLIhFIhbxSbiUEe7qF1a0YQDTOy4Jn/mlPgAGzobfsQ6RdIakDCu226vjJeO
3RBsphFW6agYxbQa5btmKvnfTaJVwDwC6W+sB4ptnauwxgJUJ6Por9xGEb1eD0c0
vzFZfVRSMNmnGFlOM8kXk6c3EDoeX5wNEeBsm4T+ZGBlO7NfgQecVCpE+X5sZX2+
tnc0ZHx1AzzjD1GonXhiFL/HIeUPiXEsc2oB7CzFJ0YQc5pSbbK6BYqaB2UMGjdR
/zf7++Dlsrbr1NlDdmUvuIKhpbct+e1G4U9R3XVophiX4G4iQIi3rsLgrvqZzeKv
YfApGzavGGlYqrWG4ZZ76KSoV/hQY6rcY6b2YaLFPa/NYMWPhJkKhfqOtUAitvZ/
1KVL4aeNGXzQzvJqAr5x5vzMB53dcDaVwjmycJyNjw98bmY2EVTjNwoS5K9aL2Lp
dWj/eb3YTXZTPRNjSENQhXrR1VjGGLEbsmG2NBjVugs4Xa8Znjy/iJytRZOMHDsn
qXEpIsU7QiQPqoprlSYKscPeeDI6NeGKcHyfrs2eIefjVzxpfqt0ncjF3r7hvEz+
mFqrqsTLS9S9yZxBEJXoRZ60bjSpKE77QBo0ehXs9tIU6RGWS2psNs7tX/lvAX6Y
M0Md1aTR3XPRFzybCNwubMMYChK4VJgjPWfigZLNtjqhVFikXzDKmJz4lrBuNUYk
DpEHMMNP74pxzhG+s3me6IxrQGMKFw9P5iQAOvQlvXM6zKF1GpLFqxqD55iOqz5p
XLRZ0zJ+yBeSYh8gTRMnTnp5F9RArjjt1nrNy3wDwghVoOCAH8TtkM0fk8jJ4LLZ
AO/3Y+xt5K5lCAXYSxCVxElx/snGjs2NoogPFZ/yWWWGeFVYcDabDNIQPjf0ek1f
LvNG57qO9Px8YUvYtU6NaibbFS4koriCmwd3Gc5w58KjniSmb4lTwK3Jy9TSyBp8
Sh8fCr2Vht+KOEWkSLWIXPnldEFCYUMLq0vazGk0DE7qg1wbX+9yi7EFA3c5wPIj
prwuYTl1WTIygzPCjThKgJ7LgV8awZk06l0M0tFVipa063NoP5/LRmXKxEr/FYy9
WyNMTuKNCcJ75RxAb7xizrDJDEGke1ULhwoxLZSfHE30mLE3FtyMjzytKWlNivpg
DgL2j3GSJXiu1Z6JKyTfslNV/Kbxb1tobl+5+nyjy8UTev69ip54FyDZ54a6KXbB
ytE31u/84hOSgdpTTg/HEJkuo8pqj8b6TXr8vlujAynpmJ6Q+a1RTe1aZT8fcZRp
7LjFBMVp50dJAP0HqoRCebqo5mtNNo89MVV0q1oab/SWiNIlaqj2r8lQeWEzCft0
aMODEzWDzeGBiQA7jSA8bozAtoyV/4Jfl0Qh5byV3kBjseTSriD4WxWWSRYkbxKm
Lf9yHOL8ywfTUSAXHJmr8tAB8uz5tU12zEXKarixRrEXeq+Y0S2ptjT/P1XTx5A/
YOBKnoiwMKPf1Au49/lqOT/HKnqcFMpwKXWxrpwI2iH8VKHQ1ATS4Rt2HqujRLb2
dHGveLw8jX+jCPEJ+dpRDgCKU4MTn0jo62lP5skZuanTqPRzYWYfNpCxlZE8YUf7
ULqzVk7ctlRAywaiODENEK/FyNuMbga+ty2aSAldTcEPq79HlVLfsQRoiI0zs6zo
Yk6CK2g0FykBDgR7zayxU8cheh/2iiCAnOwkfT6nSwrAQxWHfddTuYvd7u3Rc5Ln
wW61AkVqGvwDeOwzsfA39/zGpb4rsJbWVHGE5bkG+8aJOGYvJPX9iJ/SweM5PeKx
+OnBA8PkcPfj5V714IexAvLuAGNSaZHjMzCzCZgXdo6FCAn8kLdxpNsDQ64uiqpq
WUKmYyr4hEHdxToJ0Dd76A9DX1RXzvd5jKUDMqrjJ9l2r31CEegskGP1jEi6JIJ8
bN10devc84yBzbMJcASJTk4OTbVsWt3ZJyn5df13orJxHQ74HNsEF90637hjdpmZ
uIhNLvJGA3kKnUnZCZWh8ZBDXiL7vyY1SF/oRx+ybUw8cCSaFg4tb0LwGpqawTpL
uhnAWRe6ck9rnW5DrN8HB9KHc0JU3ZpxaoyO1MAlXRS4sRolFOZ62HsYv3m8PLx5
SDLMDMTlf2omLObvoN9dAAi4ym7R1Qb81NVCsE2FdHm6aJUydT6HHibVfkHrbi7+
iRrklAMA6QwrZ+nlzLTMMhqeEGeZBi4oqFzY9qG720NMqz0BvFsWeFdL9lWWCP66
abp3Z3ULmDHoT95iz2UpB1UAygOcONY0sKeAsR38mp8XQsGZwA0x3mRQK/ICG7i4
vH3txl0hUcZI2nKoW7LDpaXPMHpfdFb2PEOGlRK8Kv7AkvN7b+kV9ss//bSH6jx2
mCzjY5jLnrvFrFCGPWCdMaCITLwAoTpT/S5lnHMA39B+idVzc77+J55YFFBVJr+0
wL7gnpM3iaQXpDHRT8LPuMzv8qjNrPDGgmMgAaI20M8nv2T7RPl+9xRahvAS34iI
MzFWXRlGfh2KOdNW9Lb9wBd4kSyRS72RHe7tQ9mmqxtt/yh2BF6EBq7lOQIgJhLR
JtCbCgbl2yTh6APiLX81YPtTijy/vWhSRweQqYANOTillLaTvpZbNL1p4PH5wgtu
7jKE7UKLDWyJmk0VuxUCjBG/YBPI30HptCuxFP6CX6r7H40oV67//Hko8EFR+84y
yy1WVSiX3UE+pOY/oDe83yY+TZywzWKyrLQ+N1uEu2GhBDE1TWeczJKP3x7KNsiv
2mKg7gjkB0AO3CzZ8KtmwzuKppNWg0E520bOU9b22v75FbWEI6DN5ixt7gTfX0gE
IUlX2+cFpnTJw2nmrjBthU1ICkFt6JlbrwjSfV2QOF8p9xpmxLciHW40wjDmXWRR
l4JLIn+VOubaeYPvXJClFYazCAsUAhH1zhFs5gmONUCOnLhFwkoipkUV3cPmISlx
9MLull+Qr1OrAxpoWYgKNdxVVlOHV40IbDzWSi9PsdzZ56D4fp+G7cZOzb93PphN
GwjnlzLsV4tT7e5xWbM/zja9HvSPH9tPk3g0FPKSYwjLAZwf5uFJ5c+EtrICH3vF
ueYwF/LUk1uyr/I1mWU2QaQ4kf+vGHIG8CHGVsv5D7L/oK4NG+gVWcQQa1G0m6TV
/sR1UcMKK8l/w3UVZk/NdVRG5tN1fsegmCMFF2Z2GRCb4tRZQYQ1wVJpoDlI6Y37
UFHLx4JMV23kiPkbwX9x7gFkScFwt0TM58u1ZgHcQ4SyaBUd9ertVUKK53KoREX3
A5OJYRAU+yQZ7VEcNpz+1JuwO0OH2SbAFKNl+Ci61pnkdbjH+g+SxMhxaw10FazC
6aVPLgGG1s2fZRJBWILdZRUIocbgX2QTJZLYNte9fu9smBTUUk2i/PIJ36l2SDn2
0mS93sq065zdUDYzcYx8vuMeGg6eqd/3PouZ5YXFFtNVP2ew5/Be1m+jcAN7FTRp
EpzyS+4ApzsOyV8nVePBjt/JApy2gFxR4F9/0nPxEL/gdtyGQRAemav10FoOkDL/
Y5D6cTJLqda/gVoPh6oTNfJoEvOCM+5dXeCp1fj/rf1legFSRRAblKzRgvozYBZr
tOI5EbWx60TquQ4FzB6iNzw2fwVDl2KnZ+w+oLYVSJkO30tubF/CfkDcyby5fSoE
wNhnjM0F443LbYgC15VeOJIzhM5D1gd35+6dxLewZHu9kLC7bnTC1VDCBhFtDrFS
cqXToWE8mEqdQ1QfUm/uNIMjwb8g61UnQMEMfpPZW1C81mrcHY6vU9x7ymcxwKeV
+csPE9a8IUISm4eIyvs/A4ThEJ5J5/X343LJeyPBJ0oYMO4s9mWSUuEDisnad6Op
0cDrKUnkGbx1QzxdmxjgIhQb5Feiy5PPcSBXMbBBzSOU8Gq3p9Ua+Jr2IpX09W9b
4pxhj1UmgLtgDs/AXSXd8evukiYdUylrlSBON/OnOnuX99JDTupSiP7PoaaCfQcJ
ybCGBACo9AynGtcLihfxZQVENtqdFJx8WcGtfFCXCHwTcrWYmcHhbWP/9J38mAfF
kHYs0BTmDyBDHcL+KR4YZ9GgZME885K6oolym2OF9b2T71ssJ/ivUbCKYaOFHryx
AlzttsFOjGfNpirWpNF643Z1X7HroQckwp3snx1WXtBzC6S0i3PprFSmDbH6aDOb
petJVl4RgiYpa25TkXLO2Yrn1kG7eFat7IGwROHP8vn/uPLRgxuWKa1k3XnH7Rea
8o7BdE+SQD06vXieqJiurezwI/QMIdJEBZt2cBah+bXQxUr97edAYB5Ujh5ZHVDe
fMgbLptaiPU5szuMXhmZvrYldCzz0BL76V+6b13BcN/QjIJL0aGWKvHUoGF2cwXC
Ml+hmcQ6pM8hJ3KOUNN+BQHkXCkw6FUg/g2EJY1I/xpo+cr9mUuVf/eda0qQGUeM
KFaBf0+qS7Cwoezo+T508lXfVXxqau4Ie0Dl8s2SMMdpeX3Fq+fzcZK54apgGj5p
JtriEZ60QqOWII9qCX7s4JaKCMjojrT4WMpvzRRyubXlhSMI4a9f2AToqzZQhvOJ
Ok+U/4821zNZeYNN08hNBVctSC9sHmfOfKkG4MWFhCmk4o+TiM+nEMlK/HgK8Uao
i7lHdsnAs3GcYmiImV70gf4sBCWNlIEOJ0GxEOS70SwZPef7UqAM9VUdg0mlK6D1
rEsZyoZb07VEC0c2HdixwMF9lszs6wcbKkaJ5t7RS0BSXaR7N11B4P/4Xy6I5H0l
5HxTyJNQbFVlU19PVdmRyjim0mOFRC6BjKW8c6ZuHrbZemIWnOj7ctRHBYl6LwNB
3QmSQ1vxADy3Jms/98YzsdROcYAfpngzA+WKk0X3w+/YpJakD7odkaJjVg5kKcds
zBQfgqWFrUH9o0uZcwftr2fKy24bCF3sK/Owg5rWUqjkLKqn++A7Nj0W/OHH7ZUW
9Os7ZZ9oxacSce4f3PQuTaOu5+MhpTDJ6oJD8aNi/pyM5Owz7P1tlAFx2y9g8vWf
Rhf4GDlFsESE7CJJUacVbo3gUxYa76rip0UHMS6VaBXBpMv4yIufKN/7zGx5maF/
vXVk/7m1cunlaDS7EdiHyqD8wylmGDd4lubedD5bPkwLnnDJtWQYmJGpEVpJWBkD
4cEccwEoYs46By6/6Fe+TdXYhztEBOXfYXa/jnJ4Hww8FXurA+8KarQ1IqXQJLsc
+DhvpE3iEaDcHLXd69vb8zcRhPiUoTkfPirIcak6BaFuqt10Yq7rjPCdOucLlBqW
p5/1c9e1gcnbFHOcJz1ul4I2TOYcdpob1y6M8uWZkxda7RpCFB33s3PSzPYljZG/
48HhqNABL9mflg1/d5W2+66nNoAy7xSG4WJ8m0fP3znYHKYXQ7500CgCVvOQbmAf
8g8/9RK9bfNB0hkqSLRVZIF4MrTJC4Vzz5vi9nRXEDKWDhy+1dgGFr0hbqicQYl8
IBj5fl6HVYzRqi2GvIpNkZMssrdy4E/BZ32jOBGXwd0TWEHnp1VI7RYqP9+NdVgl
BmLgdggvfU/4pSaAIbRI8PYqWovHXOb/jplnvg0KtxV3GD841qjKMV0V27X/BD9X
fUM1doSbl87/PbLilti2jyd2wC66yZatZGBj9LiB2int06/1g848fOipQoice5Mv
i0uf8GaAKr23u8f+oFvZV+3YpqG1FIZ331UTo5MRkbF/xPMnRDeGuCa5/1MzPcnj
TAwBU9TgSxB9WvRKZUt8K3LCKwTH01DpC/ar+56F0lp0DAompZ4XtAcaXDBxeQ9P
dCIfnuK3vrDuQYQCTBn7gSDwwmMKuMsS4HBeABfjzz0/ujCokBKEuvo3gZOs6EqM
Ybbt4JOzCccM/vrnB+IKqCIieYN7WstvwBjUJB4pjBPODyVpB/z58WCIN6FTiTbY
2Q17IYwLfEeWFlCHeVTQuWJC6i3zZzXxfuSNFxqo/p9m2EGsuJ4yZ/GVsq/Y3fIH
SFIl5xAWJL9gf0vy0ZNBTtv4aNJMeeTDFtW0TNFHSVu9utCk73ETs8UwtJNh1mET
+ERXwGyiU4V66QKFWGT+9hFd01Q+gdfOgeUw8wditEatAm459LOKnlWpa17fxnSf
ezuSe9lJwjNqAdkKgTSz8/45m7LknlSG7G3TFRhc159bolesmlSHd3HK8OR1fnK8
+zof4FGqA14WiD0WkujQxPNLPW1/j7qYZ428rcQ2rAhX6Ki0RjNxrYlTHNwaaS2y
PvCMbRpAwJ6mLHlSX/LKJ1SAP4trvYly0/iJDbLkLVzgb4DmX3QaLB/DsEgk4Jl1
Dqp+c9JeHWBLJuq+PPqTQ8miBrRl3WOqhR/JJHwBfDUdtOjxKe8xoWNeJRj+CqcC
whfZXhc+OfOUqa9ZtbAKTk4jdy/n7qczY8ziurh7mgby0bwBvTWI1Mm+Q6iBkv0u
NQgOOM/sr7yO+HN01Nb7S/xY4/pD+A3tId/jDq+Bdizf+FSLhz28uOBZEbnXA9yz
dwe0AnyyEc+WTuKnRXXwaZ7IyxuBEkWUpopGbnzj6uAIhcUTBxo3tBVNi2uLK+3Q
XfaY72fUShkUMhLjOwnaTfVPHQlrLywI3y84Zut4fDnS9wNAoEUHORUDmoltNndj
1HHG+8suNol+H/g1IvBUJR+QhSTfZdoREl1NIP+sT9OqZjRvLp/aa3wedt4lvu3M
JBHo3qcxo1MHP7T675stcOoQdM8h8QzQcMUr+XU9Yi4/Et9ArrW1o/B22Tsouiu8
hIpX8Ktc5M3flMPACA+GuV7QH7bf/NMBZdNI2DmZUveViUuVnyfUIGiu/94P4F6I
TSTymq29+TOM/Xe4Yol3cw3rjTjUrlRQYL8kU4pcVa4orb8AS8N7mi/ubSgIL3Yb
hjJGr7dzRfxlKgeOvq2BaBqs04Xv4+Md5rhm7Ms3scr/Fqv4TGaKCB8M2e0OGUIZ
3mWoRrzmff/QlcTQT/6x4h+jRL3RXIGlJLgKorz7dNoSnBThAHZAeJr7cc8XLk03
ZkfdCM5utD9uOlPdXT2SmihF27FcY/NnLAK3YSaqLyTJMJIMkiOhwXvdF0Ww4BqT
rWRy7GYKzKHnOeuGPjAfJgrXvAixwPe1jlT9CxhD2ucIYV2RMCXQRxg4ONzv3MVv
zoVzWFYG2TGKZRxEKIokGM/7jzaIRzZfxPZSbdo1sVU2SzahPAkSYG4IRXN0j3GM
BCGM0FJ0o9OqydS0bsgsDn085s7hluxwHtShxmjJ7pcMjkh5xfV5EBqz9yE0sRIl
fXfyXtAvhhXRC6uIJnWEDkzzRAX3mpn+Re1KUghqKrJPFu56PITwIurEgwkWAjDp
g7+4UTfPHFfo1Q+AFI2Y0SlzNy9Ybp4an8XGcsSQjh6FoT8uQO4rj4OXDkJCHKE7
Xogyv5MmtN7Zp0GO8yzZdU9w21xWD0jVgtBav2dGPtbxLpLAK2YV5tPmlMwIiTTu
MmuGeK5Ccjmg/PVtZPwEX9vD5l6kSGc8naLe+WD1ZETsG2nykj+M9TbSZSTzqzpB
5E8Z4Gp6Q33bwIKqbOR2o8lt2pyBa0nu8d2RHYQDZkcpEs4eMuMKVbds9NUy6aLM
isWuiHS2XHIFewutxQDmWRWupQ8lNlC//6saLZBJ32H8O7t8Zt576znfS0jJ0cnx
A6K96zSyENW2r89Ip80t5rfyxQR7jTg6Z66a6bfiog8zjXmclhEaNLJYJvQrdB/z
vNNsN/e71BjrwiGKuvcZldRu1EtwGFsOpmVDbcxkMo4L9Tzi0gWS1Asz7k2aG7uT
c32Acdqi+867+o6Z+2LkF+hHI66hJ2ifWeBUpNx1zbcyqEY1tjMhdEZ4QfSqdTd2
bDwXMwk0s2dxnztnvkoTn470+oQdU6vcPrCakWMwj7NsztaFvtnkXiyJT1sqXjK/
XSGAkNlwE31qRoS+AU09fYeAaWdAh9mspdCVPv54Xt0shclsA6UEvGxnA47BQCjW
fvT2Ftca3sQRkfkwrgyilb4BlgdcGasFPnX+I51pfF03kgInH6vsAKhiU25FopuZ
oGMtY5x3W/Z7XG1Zxu5aTyXZ3xf5PE9yKvowjf4btHthS97ZVy38HolgtSq6B+ui
9UJfWzDuoMIpSTTiVXvvWvfcwtvQQhqRRIG6QPFSmkNaTYLQ6PtZkdZ8fKG4VjvT
B8/6VOSUdP849eFGVR5g7SjeJ9M2W1X9xTETzU6mL28GuFPSER+jWaXjWq81Q1mA
ksm8DWRyATGarLYXDVfu6XogwL6K3PT3FDtMzXaIrpXM9uMKw8h4CPK1N93WX1ks
kOKjhXBvTo+pDwEK4ocGb/seQVWZG++FAZfGJzwvxSQCUfHhhpOPxwvZ2q3dJrN9
QCEjivIJSJL7tMHXZ18JamQYtGR4Zmr9EA8rJ8V+GZc8G6HmbufWIubbcnLuId9e
CmahC2f72xdFJH3HdiXdirN3tLoB1z69TkbOR2ezNTmTWkcjE7A3VQEaeVNRTC9X
bGfPoyiqAEDlMmagOi6kx5b9f5LmYpDGLRshj/TVK9khnDQucfWEFt6uBFeyWgYh
4L4S5f9FLz4hT/1Te0LCOYigNN3KmkTU2HXj/AL4erSUcik6gKkCk0WVjBaVug96
3rH2W32aohPwe4hxYzPfF/pISENLdDbBnZjLH+Ms8/NBATG/aMFNXiIFXn7DzPNA
fpAFxTArxIri1ij67PC6t/01qDbAM0VD+FZqkDPe/JuVKfsncGZ3+19OyXZgKJBt
VyWZ7Dj0zjLAyTLH8PJQ40nHRfEJS4iDajMVNd+Nqe4l99cj4VSJsVfEe+XUxESx
NnE0KWmj3rZ2q9UcLWj3jpmZFza2QuUaM8KCmAbYo6ddaKOnHIJb/E4ED9UOVoqT
z2tuO+Ix/CguOZxg4NylK0ZfMSBgtZCQLnUKrfvz8wQ323S2aAnYThhJ2opnhNmU
XC3PPX7WTKM4Qz+9RaShnZMlvhxv5EeUmryP87ODaaMT2ay/DJKzZ1JNFPL1mVce
/aZUpyIVGMhULlgxOVrPF4W3unDyGV/SZ6ZeSgV6iN/93sQyUEzQ1LZ614D42sFc
5qy9sQBc+iRNWrBu4kR4ks6HCxfOM75UQJb/ICHmP3qSLN6VqdkgPPw1Y7HVFbkv
+SuFFaLYllwVp00Zz/BYSXsX6z4/5t3Mu8buw5zNDx9nLVLRRYneEITTkkY+NzFF
BOBb1QnUFi2cEc4tysuqiDIH2R5m3Ux2q/eB+189023ALHwuy5AZUzYufL5VhvHT
z9ch6q8Zi00WZyR3kqUxxlUH4/HwZfDeJ84CbO1hSzVgcPLtK0Q9zrvs3fdEn5rY
etfE6s45CfbPgeT29ZB14V6QG+YQ+kpE8d806aq9s5oLpuomddiHf6PbhnenTDCU
I50xLqWW9VTzngZYNYz54lT+gwtbQXIEDJaxc74uLK0NRVEaYYoCU45QZrcrUTZL
Sl5/ioAu7307egn6vHSGHr2O4mFXt0U2GwDvCXHpByqWgAoZb2Pa+SKDJgIV0Dqn
YaYL5Plj4PAhzSggqDf4w5YzizbajKVWu8sc8657MiagagJKuLveO/XdTV6j7LHE
2OtD75+uo90abF9eOqhU42oFZRCdJqlf3a7/+cQiIy6vZzfq1l5bxFcLy+Muzele
dItCskA16daxaktLXKnX+3mWXoAZS4TMIhIWe1kSq249ySF7TpxL7zPCq7jT4f3A
wRhqWmDjDMWfzQGzfHkJMnl7WOG9mQNKfTl5CmGH5htNa8aMaxfh2VdCurJ8SsPO
LEGMrlGyOJGn3hrFeyF65pAf/4OsYduMvVzIW2YUODSJgGse80T2X+89YEi87TCt
HKBNjENAGtPOHPfnq0BhjimU5KCOmJVbyjH1zi8sroTKuFl+SRAIBpNyvtrOF1O4
xhfVmOFUNTM2c15TZDXNZebsq08DiKunysE5iPJBq7YJpnxWWmKaWe3ZC/Y6J+//
hVl2sO1npQt4ET58kc+agZwEMCFEXxn7Jt090UVO+LKZxqii+FE2P01UI1jA1Nuf
zjk9HgtbqdMKNIsWZBszmrKVg5KKNYxR+BGk1QOjf6uF6nPv4R62mVWn9dutQJEG
f/PuLGiLbZHJleoAaTn+a58EehJavKEGOCNqO3jn1veJsz86Ctwlzzc12IsU+oKB
tc9+QvsIm+LdP0jy8Ct73L7VQQ56PfPyq2jiWRAcxkzKwsiXHaej1GYzNWpPHiAt
9mHt8Jgz5oa2gpBs77Ko2G8xqZ44nmLn/BqNxF8RgbbnJ+eqjb2oWFYdK0Y8YFwj
7NEy3G00Yx8WIEvwscphFTZD3/R9kBLn/FcPE6pKBKPVJ59P7OoV5Hg+TjaMgSMD
y+ZuiQspWvcrwh1GN42v6/5rmb4z0PiZ/NiESuE++Qm86iokdGJQaplbjAOJbwIA
QsRAk1BFNKEZ2/B+M2NedskJ1BRSmAYOf7swlGzZ2Q05G9heouNTstngNRxf25gx
fzCGs6+Rl3F4bgj/J5SioxeylhAvYgkSaHlNyo/mkVYawps2yvTGAiyZNOM99OAa
OOrEJmbnjwyJjC5HmchrainZE2DQdBte5/KvAAHKZO4BVCj1W0DUET1vHhqsdXK6
/bEJS1ZiwL7A6s1J6J/KPnBlvuF5aDU7IbZ5Z9wzRnIP0TsINLU5zCfOyv86BNSL
IQr65p4VdBaDqSxP1wF4gKoYgRs0lffGSnKMumydU7dxLEVMWTii11xSeX7Ov7ky
UrL+571uJF1Ny3nkP+sZHv8otiaJJBSrc037yKUKle9QQRj40BTWormMDD4JPWfd
a9DONLJDq7KUhF/T21vSNG1mKRink4gVZqj3y/zaqkFPItv0V02JzsYEKAy4irOc
lKFmFWPCVGb3s+0IILZkoZ9P2S/9btMOz2Wx811MyIbiOzqTrkUfd9i5TJ3kuB5c
d3kA8rg+ij1xs0pz6TJkQx7CX5HW/SwTHqVvrZYsDCuHTAxdQCNaDUeknL4VoqyV
LtOrCKsfbYYpkNkya0qZb9pgndlFp9J5bh+fNsOUEXiZKwYPvXs1ebbBg6FcGlzD
fbTj9RE9CSimNJgBhFdWtCROPQgsTXMqdeiyQc/was1Xo0FbhRRKF4qyrrjG7DCO
f5KJhGHAblpWOoWAeQFF13lGDEHXw7/pAN0D7aCTyXP6nlhp6qyk5PLt1E9NgG0S
1CYiO4j4ua8ZxGq5VwWIvK/9jz0dZwzhdyuuOfPBvUt6RGizWLTQj5Et+dsCrzQJ
SkV1F4ivpkeNiWqzfFaAdWTQ2YQEkOawrD0kt0Tk+skBzT83Xl3Wx7K/s60r1qow
YGcrBbIY9244MnZME8Lnw8EYqeZO8+SC2mHRKyWGi0903uraHqlWeFkJpC8F33Hd
blyfmDnHBgNhQM0UEsK3x4cJgCdwO1gnyjYg6NNnaRBhQ/L7iYNxORIQmBUEdAXY
gEb4sF5pUhMvqiHnSNyRZhca1ofX/dW7Xinc49CqWeoHtRgC5VWUEVD9pFpqJm0u
mOh3UDmkut7+Kf9R8jXMTYg1j19vLzqf2kqg9Cgae86TkMhPuI8KrCaJ0aX3z6Q6
Amjc92Z22GQ1cy2hz5gnL/XYORhbBVxtY+cirtdUwDWQLcuPSO7RD5mwpTHo0TPn
VHMkO8DhLAffwH75zIzCTTpvBWa3KPQYsyZyQU3N2rhMbITznAab6MxWzqxOR2+R
ijhX+7XV4Ot1OEA+8KDlwTPLR6GuXIs36iUx1rXV/itOrQZGsJ+V7YkWdBrm40YT
107Er9WapDbM2lTZYKGZrBeNeAZBJqLkIQtJD83qtR2Ob0BTaCy30sz3PSnX1yqe
pdf+MM7AQ6m/fk/4YfvD16sIjXbOYVF34uKbWyhTYeQpceVke4J6YFldJh4dYs/J
kOv0HzRPgxJiKSpHSvBzfM7MO6QixxHEVtGLzwLja3GKyl26HkFthMCe6saB88vu
pPYGgB9bK9vCKhvFJdJA1rO/F9o21U7N8J4UcYTOuj0TOzhfgMCIatDbeKmAxNhe
OLtSm2S08DpitSBJ6gDN1V+Gx1hfQXhf7CkNwaXfsD1S45Y74Ttp8qyCSVdav+IH
uWT8JQ9SFp0UHkuRP1CPnAfO69+Fj7IapB6VAQCwZgRfQdN2apqRpetHjjF2YaGW
qMsqhQNJVn5HD/rhOlpJf7Fltkf4g9j5Q1KwLVHQkbpbGYX69ySymFPvWEXg/wDX
QTDrzaHLbxKxTN0fVfjHXKFbgauioG13uTRtoqb8CIUPS4HIHMdfWxqj+OiebKBL
hOZXILaOOwKchHGFpaD2i0D3P746qxxecKS+vaZPn9rxFQWYzyvcPP5OOnpnUwHP
lzk+luESjWOts+t/7sSeU3hcEiS4rETDmLyIP4eIKXin2z6CbbqiBYllHCD9l3Sq
ufq6EGY1q/dm6V6HHC75utIrOtYcovoUAk23ZZkbcsCBF+yw3Ixy7xX70ZihJCOK
2hjVO5b9YUh57zNKbez00LuDriiwCkmDqh7x3vH3DxPWxherqNBlgARoCJ/gUpzj
gYCt6g8MwR++QpxOhHUeJ5FunO9TD0kxfOd1XxUU2Kk620C4Xvuo0QcHbNZJ6sFR
3PYNTbZTt5lHXW6dW9oogO0WWOnpnbBRrxjKXJVBSBu1d05iD4bLkrM3JfcSgdJG
gLTtgizaT97r8l9+TAY/iWzDUIpcyGYO8agEgaBOLflvgl6Cv5KNGbFwYumAhmCU
g5WBRoRN4fS4iYHIOKIjSbixL6+xQll71pFRyEclDoUF7XP3DLg+NBLBpNBOswFN
8YPsUtIwWe7O5A9TrQ60O7mZYpK1mwYXAgiNCtKd6/Ax3kfNHs/b2swH5cBowLcj
Fj5fh+PijrVjv2YOAcosJHOyLsqTCUGb1qGfm84+MpMbneeBPcGImnx6RxNXULgN
3h5A6GCXNpsoboGC8G+N6lUd9YN/sChFddoZvdfooFU8BOTzKGTry+Iitz2j5FCD
W/coY5lbdpOsgc7m6mQW+Vp33VZvRRe2kVP9GrNSnoA+ud9FAhxVFOqS/eZWg5yN
8TLCBRjh+41jP1IJB1B/rRj6tmriYuDjDIUVF2gFwqzmuujd9Cqer6XsvJocM5HB
uXoRHtxTG14oXRM8oS8YuIzkAq/VtxVmlWLwcDk9ryZMb2kt+ZfjwqHuLNmItMe7
J31cSiODtrQLdfOwf9GAFx5CknPW/To3fDUKpGeSEauai24G/N0EoUyq1Dz1mZLK
57jOII/UmgHY2hojxgFqpuJLCyF7OkY56sc/AiAgmimAVVmF2yI6Pw7JGkKu62dz
bOt+iSXCPWthpqFdupuLr9bLJAPGn92QXhSOoXN9Ya0I8Q6/H7DTC8FI5H1Yf5l9
/nxFzt91/B2VAQvWFLZLxMZhCIYOgvnNhL6xbTs7g2y9UIL9NZO/8E3Es56ShGLc
tPSTd1sO5g6cjDoApV1OOjYN6ghqA/YAYH6b4s5hb4OvOR9OjnaeT4QUP8tBJc5x
6tdOpxt617eG3DjLCBra0ICQ9jwQrxnbZdJkcJpnXWJDdtL1PD8mIHaezwQrjxY4
r3rOcGqQPpNignLO1LTKzytT2M6UE9ZJF7yzM/tCJmZcAxRNLdPTeRxNuJ5+ubjT
H5NIoohHVev7V1XSpmktjJ6kIIOXJMgMIrkAMQMCKFi3cnChrszcn4CvWXHfxEFx
Xg3ndbXGVNVOVrum74/xgx6C3+m6ngR6L45ptryc9Nk+9kkl1DOaUkS7HhB+tJr3
ZtgGNL65bMWZ5QCJ0ITEVwhZoAil0NtZRdiSnqV8ept9FRMddwuaOyjESOQG6FZc
wxE6az79JUp6ahWkxFIseJJiRfdn01+4rpW4MaveOhFjmGOH35gKY2sji5BAnvDG
R+kR7d2od0XCRJN/0DmIIfUI85u68e4unxmd/sLPieHkWkpCK5FGBWLv+rv5re/Q
eGlPahjvOu8HIHUOwL9WxP5tVOmf8XM2zMZyLoxH9JdPapuwvlxO42yYv1s3GAf3
n3MoLuqPzV0WRbpBWYTXvjDgodnpOJXN/FyXed8230c0XXxZ2BvnDBZ66WnxpiUG
3KXXdSfJN512UjIibXzSLZvAn5Wl0NjxkllW95wZOEmLLq9OEZCY2zMRE3zC6Zoj
Cfcrr54c2CCI5CBOuACsr6JzciT+utoU3+BC6GXQqTZvPcXq1bk//QsDI0I76SB8
3CmHlNbany5E6wkpVhge6VKbWKWuj2qQ24lz8F1ioNKM9UdZOTsa+Z/e87qh/w4h
fvR4NJnAY8FZIT+7I6yv535uk1FnTv7UX3OR6wkRX89XJnERHF0IJmmEd4//PdfG
h8xLZOEv+MMdLtD4lQaYW/cH+Ezv3ARNggbxSHtLuAMRpiJ7U55Yl7sv6cZtJKAZ
sFO3VS5ZS9BitI5rcDQZOLSUJcpINMlnv4wl9vpLwN8sZZ7Cs2VTfoY5IhELfRI6
8PN0IGkk7Yb9YrvOrDnIRlHu7dEUZdO6sRotkyenExuBQWcG/Vsqw1ukgyoXUtQl
yNuSCh0e9UlI9XRTTTgQHZGXGknqZBv7zXEDBkAM3n0sHGiLNOGYzTYTT4zuExUK
mVGP8pSUob9NisfpxfAMHlX94P/RopY50O8SQyo1Paw1VFMDaU+KRVzPQeO9DvJO
sQrdXVdTsIXbPuUhmYd9cIdphP6w5FqO+5uQohByI2N8YZyqm71JdBdZ97HPT3Cb
XobFYxOtTYN/34O4tlDlCdcFRHlYB5/FchpDnWXFq1AqLBEmLHyZTDrgHGcrq4fE
wB7aYkGskrC8M/dF9RWZKo8Yw+AEm1GIkjTchFsDTTn3zGD3X2LTFyUkkwRLl0xC
N5lS47/p4yHXml3eAovMzi6pk8/CJH6bVybJ5zKSemH1+d23P3E1Vx4c+kQdo3FO
N6shxA8mLwu1q/oSvD0dtQZb1uQwGKAQeJGEufWr+UAoualfHtyNW8cZCs+JLvjf
waCpZKZ/9RtIVLx2z1oqksPF2NXrR+BDv9LpCoAycdCNWWH28mMrQmn6rdnCfe77
myDbhGjDiR0f4vTSonnD3SxUiIbntsrp+ZhCmwVZ2DmgoUpWwTP+2LtfY8UbXzBm
p1CAPFYW76jgisT/B6YUnU4mf5zL6JuBEddSTRn3jIKQkrjZvEG08P87adEmbXfR
bWdJwO44q+yz1Qm/xRksolGNVvvrAo3XmDDVsQ7+s99F3e3giwija+0Io4WG19p2
EzHTjwpv6kxKBNXdPjA76hv3+NTWRMEpMT7lsAORL/WklkTeHQgSRZ1rj4WNVPKJ
e9ce1fvaWUJCrfKCQmk/7D8wxbTdm0lBjjl0A/qq6ewmrQYUwpjUufVDtkRzK/Zc
Ykd18wBV9XiflaWNxwBlXT/KBqAsQ7m1PchumGqor5b4jdxBPTUwRAMeExbZG7p/
qYlCiu6gvvPxwivekBwHqA2NOhqHWCLoyO0V7acICBEP4iyLA/YqJnbZKsSUMiI2
uRWtHorMydZTFgLPpePJ6Euxa83xMN05Pw2KSpzc3q8mGSf876xyKfLiF9qXjlel
pSdFsZknhhkqUdVStJgHnajj0GxUaPT0T319byWPfDuTU2QU6TDolevh4CONaP6E
9yC8tF/fjMsLhc7/UyA0U+gA/i3m+GO4pzN6N4mYpBRmB6Ix/FgMuakCe+ZO0G+o
3pVmb6y6jgEKIvgdw+Ziiq4X7pX7ICrD9zE59T/mVJSA5LleYWnARYWHc1qeaigb
odi3E40ukAM7JogqiUpKMm874LGqdrblwpZLq22FnM9b1mmm5QU2MnjSpOlfYwmV
yA3knQ0BWjiMtXDe/b7WRaTaIeg8FgblbeufBMCQIYDmuGXciwbr3zGI3VBy6fA+
2l+tosJhtKnh8UtdsnzLnp7bBAxdtzPpLZC0gS/Nkyd3TuxP3m7Z1WQAOVdLaWFC
/Zs8s8qOXQBwS7eR7gwduOuKSon6GXSt15pEtm78HwUuvroEabjs4GDzMpGaaTGN
IceMKxZhkazl2o5uQyYC4b8I6XJTpBgS/X1NJwVTco99kwZvvADEnnXkVUwtuAEE
7kphI79pbQLeSAvnmHqQMBj/tyWHWDz+90akaZKpMlv6TphahkfDkNGeyNe06WVl
X5tbnGuNa9G4iDC5CAN2/7ED8aYZWElbTgct4hwYd4jJ+qTrlL2d+sG5JxWRG2cV
KgcF1QYXimx71eaIPkkG6nAE5JMiV+TP7nXiaqgs3d/rAVT42gVGgOByAUBaV+rK
/q0K74rA3RV4eV9aN2kxcpO72frL5Z/Y5HRJPsSHJtvTzpNk8x0ySrp6S1p4HVv4
UnKO3LzMg+KBw4AKx4cY3xebEHJXyzxTkvTMF1XIkTFu5b11fy72DF+CgRGj4dBU
XJXAj4bD7MDMIQGdLWlxYuNNBV2zZebozMjoWLd2zQ4s+g6AIFxzx2AFipvL8PMR
sexW3TI0XOnlsEewpFNBeJCtdBzeAQPLci13L0CNy+yKmXq4noQaRutIHAYVZWvz
F6ZUVBdcMtjurEgE55snL34R5L/Y7oRM+Lgo+k7CgGzRjlW8CRDdgek+BvF5b15P
F9Wr2JSX5xf1PeyQ93rZSQ2uli/RSFc9ZAfyCW38xXxi3ErUtgdU11/I059KWhiD
KSk64UP4GWDRJmMF08jJVDYCE2u6wAJfMiLEFBLHzFMJsU49IR5oNc8vDV+E6a4k
3MnSFAujBQhj9G7ZDKyUXK2aPVbBEG31fKxUK5SBhMaSlCN5cI5KhCGmnxsyn/ZE
J4hPxXckmGA968LUYhyjvSyr8rSppDn8o+DGVHlRuwA/g/PbosGt+vrBUkx6IWml
S/TSwjZWKYg/nPZ6cBIEHpo/yCEwD9t3flo0CbGMdi59+xfnOkRYcJx6eCnVTsOm
sJIEAPsr8rPKcrXP5QJHginNNg1RpjZItaJqbffs7ihAM058q2zaG14KWTfPJlKz
TdEfc/FRLkYBmiLxlMJQDZsDah/WIm/Id8U349QAhU7BdexnFyL2A40SP/AfazUV
BlY/US1KnkB0iULcQ/43d0YBjRbNozsxZB24tn6sBWQpdCkzUM18mzyZBZgjnClp
r7QBeCE6ANJ63Ud8FoF/dj8wFYpLvI7QQDbxoP28/O2W8CBJ9ZkcbQi4Oxg1OkoP
9+HTGg2vKk+stHCJdsIceg6fMGM6h7mTDoKq/FAQTc+mBdYabYFC7xPiMGSrZkwR
uQg/ymyXtQUZ/VdwSBQSUz0EJxJKHj15bw4HTiye3y8PeQGm/t2hCKH30FvkTfiU
QZPaTnrGowHHcvnGuQu+stMwqgtOY0IV4O305qpsFjY9uMtTbqtNrDYdiMLFOuFO
xx7HHD95Qu/mEyxzwvCYIEca3BPKxKRQ/aOznWtet29eCzYIgfySaqBAUprpICS+
cj5a7CmkMo7k0GlO3npE1zbMsUrlJ3uzz7P3AJCbdur1EXXWsPAQmE8pFKloz4t3
6VUPl8/oMiT+/bhg7jWtnWgwSEAf+7YM5xOqwRvRWkVR1SpyLgeq4zC4+mZn8sR+
ZJ2rQui/gbAQ1A6L1bGLgt58ZwaUKbHOAnQbVN8tlsIJ2IEFeEARPXdY+cJ1C5XR
u5ZE7K4AguJW0QDYr8yKg7cc3kDnv9CfPrSQHrCQ4pj4AHwIRT7ATzWct92WtHFn
6v6pkwCd6TL5z8SPSap7LM8xbJiGQ7ei4NmE4vexqTzCIbihKLdaqUFC58zAKp1f
THNoNeMrUIuSw5fyQAFvHE2UvQzpjKLIuW2Oy4SgQboKaptTvjXiPzfjvTh/OH7a
fWNHqf/rKFWQboHbdP/lHy1YcAI6NYkJhLUbc0uGj9mNGi7UQDX2L7QyEMtszc//
EFBXfAB5++twlnZjB2a/ZzNV9Peds1Pvzw7Tlsz2Zlz0XrMUq4tPfkixyYgcUFLu
2ZT2yNrR18REnbuyLP7dNFZXt1yVx6KXQXib97G+yHtyBgJ7bqFmguubA7EDFCOp
0pLeXwXWFG6N1w/h7tVJG1uzU8e7amvuVNlb2sStze0dYkbCpoN0IeOAoGhzg8iR
sgDu1NVRJQTWxYArd0d9zRivDB6Jtgfos1IpWkvH0a/pkggMqTtWv3A+fMlY6B8p
dzUTx5fAp9l97iHehBnE9/6B976464xf9x0UQAkgBVT/R5G1PkglHyJBuJCFRJiy
7HNuwGtiZtpsIgfBYlI7+SK2jxja/vnPU1+92fedvsEyqt0tXZmAdn/kDDbhYtkP
DLrsFQoC6mIKagBm8yLRetGcAOWWeUR7V3iAJ9DMT/1GXcYt21Hc4lzxcSwhjPUE
RvZgo8akW57R1GdbiyoAj8HQ7Mkzi5LcvnWKEXTjPtYNtoVQ7s1V+5AN2OCcuTi3
Ycos9jd5qthY2z7zg32kYtV/mJ+LwPo1NxHIjC70a7JeHkFZTJiW4wpZQz7QcrAQ
VeW7L5iiFinEkGFHlSn/HlcajgEzFqUhPDlAy+K6Vdin5lM1iJBySHOTGPMmCpH5
VNcFatVz8X6XPT7RTsnX7Ffk65ikSKhKwZxsb+giC9buwmyYbCXhWf1HDCj35OTx
ENIdyOkH1Qjrf0SAc8rAhoJpow5XZnEYCR+nRP+5jUFM5gGuU0yJtK28z1yuHwBh
+SqgyJuBRy3AJ7ucmtwnJPzgqkzS46eOipBvh1jOeImdX7o4Hrwom+47uetNNNqe
8SVJjvCGSfzt3p6s54P38ZWg3m0GMf/kMSMl6RQ+BvoGdO+fGio8W6ux6TR4/3qO
0vM0r0VLti08AnnM20/IOubHGbFpqv8yj5CPXI8G4k7QmOU7E4i0rS1+71mTzZsy
tojfC3hfjz1/q2GFC/qaVtthGXCivGweO/LFhH9MjKtHW5e08ziW7dU0OMvaDXzI
+bg9m2IepYcB8trxk2cDBuUpAApOHrT2IvixA9fOB0BaIcojLAVz0v6h+VHIWBxR
xt41ZWe1WPi1d+ve5zZ/2mdBLdwYPcvrDTwODB0PcexcUffeq9MOWvQGAiHs8Xv4
NNRwqESGOHO9ziWJ9HquTMmnXQ+WyKXz1LTk3hXXVemYHoizZEfjtrOEvKC0GK8B
LhN7Lrq917BwbcooBJ7ftjldKHG3JcKZ/yW9457eBTGAauMzNmc/gjzO7YnPMtL6
qHDnbThozFR/2WArq3UioFPeTYvB0cLCGwpTYPri9SBgXyQDqtxeX3q8Hw1BqmlF
1EDUqWs3A/sR2MDGbalUod8Di8SFrNcK1bv05D1nnsiu+9sluBxZGzpPONKhlQmy
MHphRNyU6uzkBWj1Zdkx85ZtLloPbeUMFgntK3Wi+khihMtzzlbDdl7mmxa4wpMH
wXSXEVSvVzIR4fXEw0Jb4jDYAtSnC72aAFTVGV0KZO4faZLgeaSwVkQHRcM8QDSB
QGyQWWDL7XLnuNnsw9PiTzW8psknj4mVQnLZdljlyBXfnGnfkYSO2WglLt1wXRT0
rUSaox+1Ybr80GT/mkTavnIogmrxEIZT2RsA4MzyZ4bbkHujZ7/ukgcH7R1Tkpgb
0jEqOMk32ssCF40FzM8WrMl87Z/5IQ5Gw2Gpe2suvSRT/WpOm1bUWvaw+9vwmM63
eOX/SWUQFc4N9iTvgYzUgYRmJmdKId6SIgZxsRBCXzLwEjG24RZKA/Ut2gxV/lbO
Qa7CS+hMFGg1iiT9pZytBFjToj7oeWJ2Ys3u+lUhu3enEp9g2S4ZA1zgoeUdFCqb
vk1h0fHtn/IMP5kKIL9MXZWNgNfk0TzKfl43014jz41mMIOGUbx44X6M9G7EkcVB
Cn3j19+2SSfebWyCZlRA5Ocqjz6bgZ5v9xbQ8BppC9+0i3zly9tsCKuSIfigcthr
Y06k8zrF+6wvilOaCqC1I1dDZEFiaw8/pDzQ8S/MbWlUM09WWhRrVjMmU1vMwsUv
I5qz6imIl+ovlgc/s7USpXCjWv5ms8WEFUukaVt0gJTpjs+2A79ZEpRv8Dm3UqCB
fZSAM6ay6z9HiLkvSkqoTYNhqJGhCGd8nc9rXvJmnm6wcPcU5IqCWntf/RUXX+V+
wr98fIKDII0MoZsPI+axkbUUYCGKUP/CXIdGf1wjXNzWBl3YD4z0ZatExaCVAuQo
+Gp7jk0KffS5pwN6l/NCj8I7y46/zoA5E29iba6xq7VgXQn4hLhOR/87TE9pVKOx
X0pxr9FHoYcYNOC0LwHpMY9IIRTNb76fhnFHJQPQJBRStrvIhls9Q5RPn4plX3gm
zGKkgOdcLjo2QnxwBVOdXoNAJq2IzqgxQm2+dmINgKIgCCqprLlaYhHb8woBUJR/
Nck65ajrse4Px7taqVPVOBIAu8QhhR6ZNBzt1iOygNBoNmgBiLa72mJa4ZtLrCb3
7goMqBK+cmC6vEv0N53qwqDt/LWUjr0Gij3AJiGc0jyIIJIIB16hzxh+Os2KyCI9
Xjxikju3tTkHIjnfpzssyjJLV4jjJr1k8GaXJvJ3G2LVUzdiRdGhIgb5Dx3VH8yG
EE+PYOdQDUYOMkH/n5L0Uj9KdhB4odTdJ2xXv4hJNmnX+AZChdNosGZPYRecCl1F
XlJQk/TVYbznHlIW8TTGWR5AutQEaVs7XEHmicQ6ev1E+2Pppbl2OQNgO+FBW33C
z9cJ56y0FzT2g7gUIUv+OZW8y4uEEI+pkf/kxoVJS4sj1iiPzs/S7zbHKxHtFdZj
XTIMHc1hc7zTwPOjaoNaT0kEBW53ARvdulbDTSzvQCjKgSJfIjzbwhectMFWRXjx
p2jbUIfchObYusUHpWOG9D7xZSpv9/YhTMiD/icVVBTwSu75riWHBb3COGccifBb
dXJ8o04w4U6yXUEBB17nHKkafal1BkPMcuEx/ElJpWEaQbp+iEAPvdq5d/L3rrYs
nLWjPEib1LTMyc0+93YyJsocEbPygKVxiGMPXPIkm/1mC3f0T84YTbvvDB3PbPmh
mDM+w7kXmOU3EU5G/x48D8zCFERN+yTLNVVKv8qChr4xeEx6KZzqe88HPpdP4vtG
yZXPxKQOSIW2XVaRDFTGZlgzMwGvT7ybFSAgM7JZAj0RR2gRyG20WIhqbpI8oSeD
cnJY3k0hEUxA9E6+Ban3I/02fUCE+sS4a+/7M+lWFWOUloijkZcT6TCJBbyvBaxf
0bP7NF6dhbD5s3Lpq6KtRx8jPcu02IMltwp2syfbmRCpsoZW71mps9Fudy9WOoGy
yEythJtySfKMlKkfD/qh5UcTyZrVeAXMNFpufo6jKBPEe+3Z0uaS5ehAo2cMZXXs
5MspPHUy+ITq11prpr+NBr5lkF1YoAWRIAlVIXONJSRCL4VuiQaM5LHNuP9hofg2
ZFjC7G2hYf/wgPYkehRar321WIqQtY0BUS4/D8NJbYT0jIDOnd1moxNJQZe6cuJS
hnvA/CUbxwG020Sltdbyh5Ao/Zkvhm9iGEx0hDdLXv8r7sdgNp1RpmxzJsi7gPga
LJpmYy1G684wJAjpEpjZmrNeSd1W4QfhGxVr2hnaz3a69yHZsyIwzlIxNiNxWiz3
7ZIrAnc/9k73Snn5RAknKLwIxk2kx0ZKxdYsA/0gVM8ew/Vsc8h/PeeDZUhw3lro
DVH7PZtkiobux/b63sxYahlE9cZf7o5CHJupZiHuvXjF9mWKtcCLdC+emNkV3Csd
LOe63D3hVo6E+XxTe5hB8ab0XZoI0qCovCW856m95HD0fkOWIgb1ESt752e9ns7Z
pasHkOS5Fy4oJsqyz8hhFmnZCOdgf9Hz6GCgZauXEw9weytwhiATO5bdX2L4WVBy
1tCJpqkxQKRtE4EReyPr07ajDHpeMrNm+eO/Z6Is65U5wiPtulv4pCoBCAV/R2e2
GMdKSGaggCTtIOSR97DQDQOlQnV5ohA60YtBSv5Pa+90kJi2Nb5TcEHXYJC62dCm
QYcBjyfkFwHTV0wWfdj1nWHqlCoLwktb4XPQvyg0+MUNDmp9ZkXvNh4uMehaVBbe
HBwjOXV/GkuNBymb2FSJQE4hS99JrQcIEgRS97wi6vNyd1DBXsGsoihppNeBYO1u
rVI5ctK730V/nXp9zcnfeN2CG19Id7YLss7km8KEQuS3IvD4Sc6/t5dy6ytLCWiF
LNdEaQ+GH/dARKI3+UZz+ErkxDObU4N6Enj+UG1n13pg1AEgAUR3q17LPLJ91QDh
tMYZxTvoaQelgXbnjLI7fwUHUoOjl4fOU/P9MpMw7jDS/WottiR8rt9zbiGCEDL1
7i9ck5Ri4TwcCNfVVW4TMMsLanZwhU4xENPc5PMm1yFnsf6KRYZWSgO8zIt2tyZp
Yf6ailUElbphEvM4dfZ/qoIP63TtAM8OB2eIoxRkqJXomvGcnX7E5Nm0wd8j9TKl
n0ANsltPxO4jCmX+d95JX11OX7ugRlcEXGjL5BAPXF1ebAAmeqacynlvBnWtFUZt
7R6LZc8pvekpL90GHvOvqfka6uNZiH+DRgK0tX+QJDw+PO5GzGx91kGlpn+2cJMC
4PB0oYwDcRF3/hVF9h4bcZv1UFXYvUdKHw1IEsHGFDoNbHKxN393j73REJcSw1No
w3s+MsXhiZFFFljudBH8sjaufV7LRPI0zstGVY/hFoQ6Q6GdsabDaUltfKRJA3U3
Mxpaa8tKVWbMM9WqXcfKHgownHVblfKTESgifN+zPc3R4Ja1MvJhWjF7pF3x6jsS
HFCh/99tboHf0Q0laf4Y4B/u6YEoGljgw8eAuMPAIi4cMOUDtrL5iYsfYATcq/As
CGr5a2pCrT0hcBGnrZpKWFFFM4rFt6mypd507ZLe2pQHZCxf72OR3qB3kYgGh14h
I2TQtN8yg0h1TkoTNmduAC0JadIZtbiw7gLYRFzN5veLYFJAa875WdUfN6sdSaOg
LC0mdp3Ii8QKxPeHg4qy6U10bkz9W2jzlx++oiputbhPE9zv5O2sEKlAyitKII/c
3TXjdzG32kAzS5lKZ5bdZCLYlboAP98sOm+vc3IAI6c1PApFviC/IrFTMxRYAJX5
5JD8GzyvmDc2B1FBwVNj5yq1d2cVr1yXneSpUuv4RDsZdt/C/ar85VAjkzky9AbY
RAchl/zkUzaJrGTy7Ktv48Qc1+IDC2mJw37HvaS60KwphidZ+I9Aq18ixDiyz0Vg
9hJmiDDji6dtyvmIib4vz09UxEZck24Y58Dl/sFbmTgmhsKTAJTVRvyTXkmFA0yw
d7hsSvzpHO7s08/3MgydjHKUoRTNVqNqBucWA6e4pl44w/C7qGVCqS8r3s8Q5fsP
SEIEeLDbPXMNtUKi2U2AAg155QqfHs7suW/Rd/geTWI+90TuB9HthSsFKXvZSsfe
SAmeAkq97EhJzH4cfhbAJvT4HzUomE80ZMU5utMJxSGL9a3xOrgPdqYI+W+yyYqx
DS5x70BRwK1q2YHg9FNTHagY1q4xopKeZSbO13kUN6cxqY0BJEgZn0NY4UFrHOnE
FPtlbhacskEq6amnIz7bgZNWUsGWcSQgwjSq40Iek7rVCtbgcNVynEY8rHXiNcwO
7EcLOJzhWyS3VkkynJZ+dd5+S3UiG3XrQiXd4RCSxBptDblGM4/FOMKAYVZsfb+d
45TyCe4o7HZQ17WXdwaCy/4f/1lGlK2radFDkAGdqPwvJ8IbjmwjnobMW2XL+Im3
ZpHoGwwaL4qcEtZ+4A3fqARsD2z6uP8xGtbBUPhMWM/nROJ/vKIaPMwYiMYYjgud
RQNiRlApVNOANUBwfwniezgE4v6FH3tNItbxnrp/EnWpVWNbBxAzIj6BiEzjYyZY
NFbPfmcXk99o6k0UScB2uAFd7AiMXBxd7X/5C1E+w/3xAT861QuM53ghBiVYS8dw
fisuhCSmm3NY2NAKE0BUb8SWgdMNR45cI4Zp5wN+01F/U3UjuRzywdjPYwCURz+B
11IdXveRm5ROlkMgAUxn7EDQlS2fChkrOQQcJDg2TWJDHkUjZIxQK+TopqIOULfr
C8ZEu7EfBRk8rAzqpbWtASIRZKyLg6MdxdXLc4qsqSFF/JgiF3B53j8FfidDD1YJ
x1naQITt6zxKZJ1CAIu9beg8VBnFzyK2ePb5Ry4/aYH1fF6v2cnpYu8R0Cw64L/U
ek9NeCpUY5ukJ3Uo2/m+TEoGjt/RMRb62Ye17BnCnIxqojlScoxHopk0xgTFvS8R
f+2Z4NX85rf4pCXlWA+7Poj2RMCgS3+nvQN0Zr+jRpDwBV+3YtOpgLwsFD2NLtBd
zGg9aYKFmhfWGIM5wxHNzVpS+aXtzaWNpQAmolZBISwxwNH1z9EdkWL1jk4qWwty
/Ph4AE3sg8SuiRlVhrSzx555kRCo6XL0HjIeZg8SMCIay8b9keG+kNPGdvJ7DeaY
X2pJwTUFMGwCg03W1AhwF7gBUE+r+9xuIOilTNzS81rCOw3OnnW8xw7OviUgBiq4
yjFIiLxPShqrVGa1/Fksom3mUB+Pc2cwmosHopO27irKeaRTtL6D2COXIYHwtwaf
gLIbea9/GUqkFPW/pUvlSQtMktpgLR7C645mU+IPamD5SU4vEN6/7d0lW6PP65TX
T7y3GSPCy5woEO+YR3c08Qkzlh4adbcBBESsS9bWaIuM2h29t5J6IIBt7u/dvjRy
SmxAz7AoAxwyuOs3ZyJiY9KBXYRGqIaWqQi/IOnkqK+WoL+hONg6HVpu+1vCJNqb
PlqaaqtNFNtCSxA7FEQoSAjnC8q04KUFaexjaUx5T3N1nO+x65D3tARam4Q8kFLS
PC+AA4AVvk6kPDpBth4KV5gQ+hjJz9eXlopIz/rka5pFaJfkiVs7Wh2+VqAbHpgV
7eo9e90/v4zW8S9Eqdb5o8dh6ZI4HPekYz+8irXvXfwVMjQxZsB5voOzNt83nb+5
Wk3iQO0FIap7Tr6gc+HS+mTnt3IYgXiTccEIUNh4K69qRuYvUuuLoJaMg0mpDrkk
/xWq+SEN9t/4j4uy9KBFP8AkulSxypxfGWxKue4YIkKsISS0q4brlPyvmw1sTPnn
RD6fxyc454DIN/4ICzc9ZvDBQBeoPDYoHNK0MIzRwh7Gn+cxfS3YGEAU+W364yKr
CXQO4BEPKSXO0tPyKFjHheQwHQKUr8pyMg6lNWw1PHsX6fm/zBKbR3tIVYtxD9+K
24b8CjQP8vLeG0Z7wOvmlOz/Nd2OXnNVqIaYa0vaRMmSh60qpxQYuC74ZU/7h6lw
9liGrUlMPqQDrnKWufV4LglqkGrl/ea6bq3eLGwfOMXcnGkcdWfcy/pcNBdOhvQT
PUVuWB6W21LXsn95gOEzM2Zlp/M+FgoX8wAcZPDSvL/EMJUKWIRnynf1GjlY3jaa
tzMpBS+Iki+xXB3b3g3etfmEn+GhEIjPMVQZ+KrEsAaO4iLM9YwfNqPX0JhyYq9u
Hy7c6231CCgHjUmpeFEMyZctla/CuzIPYpbmq/LPh9GOuUNRC9bgqZUkYWFH8p0F
QZ5BuMxEprXcT+wcQ0ZYuxJ0YSZoaUM8Ypi9N+WRYoRatrvQekqubGetHniKOWqd
xU3kweiVgfqorw5rX6GtFHOSCjkFw7gahmGHKDTPrNnmcq1WgqlysunZhF1HvnDS
B4f9JfEcY9mwb6XzeB4/BQBYj6oioUQ+7r3C0nIvB4Bkb6kJGKFgBvDdUfUPrSos
TYsePBpWAP7EKS8bmdtiFxvuqXYYAivL8speQcFtohZBhvuNWJJWKjHMSuupsz74
fB3R8aheSAyeAetwbbg6Hw9/qc+HC48wamsp4ENm4EVWMydzmAf2X5YG0ZE7HGBY
C6I7UEx4CIO/tDimkHcFe2RrG2FMhlw91sWsvuxiqTfCwuAH3Iwgwnja1UUd9aBj
uQYhtBNUuQFdT/4GeMPVQJ7AYWeQ3dVKGUq/7oaOxY6vB6GUwPs98k2DNIbRzpCN
hnU+fABvdi3BYvdgsLmh+WiF+OB2yKlguaXB8l63+sn/KaAJUrpbjqmTuGeRpczn
btiE6WA9zAsf3cPBYc3ti1IUXQQ5C4J35uXkI1bxNtUflSUYr5icrss5QXfhgjej
b8mJ3UwT/B2yYvrbMOBs+o0QmuVii5FyIb0pr34ltitUXlen0ocRDpA7CtkQJjVT
8OseHGCFYVG4vt28JKz+CFOCGO23nnNQorZV7s5DOqjiF8tEhQsd+f8fmnG2dKuG
XniqIyo7RiteWjYWniQJoz46QB7wZcPcJPaEOUWQAZ0Vkjff+BJsezNr+LiD34AW
p3/a6arJTeXzjk6ttZFrWnO8J8kjmsYDVRs5G6l2ozWfi1uwXwEDU3XogGqXwofG
gx8tSBijVVwThJVgM8Z7RyHrhzei+Y5rnWTaxMFA3evDUZT13g2kHLxdaNSU9IMz
S/ofCqGinDUOVZ5i9QpOl6UVFisfJQio2EOB7vXvg3dDaWvvx/vPxn7rWHeQXvj6
dJf6775uHpYEuzPtjns8cpVyjw4iGLHrY1qigzS4JYI8dKjY5zgsfkbi6QGlVFC3
WBt0fKxuUyfueyDGh6Qb/tpr1xw9KVJNR/TqT+fTi0BHS3nzQCtwgzfU1U5gIQet
me9m4ZNBwBbSxql+jjA20rTxKUa3RksjfsR7pvft1a6nFfV2N76ZZiJv5nGAcNT5
KOe+vUyHBtlT1JmfaBg/Eo3ugr/vbUT/cweHJ49fUo/UO6c2d/6SgTH4TE2D4kIe
2qyw9clQVf7dBcT7wSFVaN8vC/b+vhUhGAZpVoWAqMhOID5fuBDuIRtQuSxlCw1q
TAi37PjR/RA6vC5+jbZRTgEjUz/HxkdEa536PwsndN+sgEhsA76OIwMAxJR/66MS
cSB4bXI6Zdia4kehibcVFlvk7g0bHiWRbGTMBThUvcrIK4H7UeQkgrkBYShuundC
hkWT4qIeshq4R6vaJZJdKgArtJc281a+/RuGwGnK1ZMmYwNPi4Y4XVQsAfbwQEi3
mkhL5WKEVg8v9CuDZMQOABwlj5oIMFNmfd2F4tZo18uQaHviemyIKdxzKF4//E78
yPAv1QaAgOdZkHEwige9daqr/+bv6zu74VIqE2L/5YDei6f0g2+eVDb0Ilk6GOgr
p+kP2t+B8bi77CVP7tkSftRDItHqqNFqu/LBVzeqSXQcGybXXcXYkrW/X+6Nx+8f
rBvpQQC+fHELdXUARcNd92FNFfnyrTZeoOjMiLM0UkndB+BDT5+cDcdjIvi23x9W
fLM3ulSW2PkzkQrYE8je58g/ahfu/4Gt6JQ0J12UquPwokHBsrD7aSO1hw8qWDZn
V7guIaf3orCEwlIY8eJfpmsUT6+Abnv56INfGrnqdAd+7nNZ4f9bOYN9fArbR9s/
d9pfB6o/KKg6WTBxbHaO5Z+l4wh0DVzalc7Kuh5bAMgmf9UEBKWPC3MbiWBDuM1X
o5rWjNQGv+AhHc7adKiQRkNaSZk7JeO1abWubB0Mgl7T+cafi02Ub/VNb6owgROJ
FybKuMLExb9U6UD+Zz/DLtJUJigk/fYDONPwhtAqdf/tKj4D2yvpWar4e/75i758
MRJ3QA2GqMYkf7NFdIVkJj7RfgMIT6cSHPBVzr9N1VMEN3Q1vvDlvXFKOGhrROzl
JCOnrYsIpDHCtLtVhPjSbzQ+iIzyYcDOqf9MQegjWnvB7X4BA2uGxB1+gAUg+r9E
GHoLeIq7xwhgDMymG7n4g7o1XJGy5s29pULGTgMOOfqZqFYhiB8MnpnEJUT8g8g7
dmp75uZKI0SjnvmaxHN0Hl4ZzWIyZShEUqcp7BZXqRnD0Nqxs43kbTvIoZSD5+5v
Rzo+vK3BPdK35hm8JzzIcQWjXRVrAWfwtDb42DepqXeff6vVDPYIlZP51bNyNrJO
BGFK+PxGs8dkCcF0djZCSxjF4LolI6ML4fhst46iXmD/wpcgt0Csy+4t/bnLptli
W/fYRDSSw9Ki2pc1kBhzmOK2wF/O5QBsDTgJguP249NuFnD5erHh5ZjfauIi2/zi
94xrExHwATpPt7AwgDjEH7nQtkeH9gchbpgvV6CzqLd+C/93H4uJER2Ts5QquGMY
iTko3VxlLhSJxcjJP4qnBWk8yJo33D1HUWuYgRxKNrIRWnx5H3IZYYSvA7zFunrG
+Pbr96Xeuch90E0uXUSzHC+uZ6AiGYfBAM8CjCpvgDxVM2brpxg9JLYbzDQ7sCj0
vzdw9OdgYQc5NJ8dyABkqE+PUOeIQbVrz7zTkGMoEvmTatftGlDlF7/kC/BkXa50
c16gQcQqpwGoQ+iIXDpfxDPv+AiCyNjrwV3qnATlV6d5ibH4wL80cUovRA4t8vpO
CanDibHY3qgdTOoScjdA6OJK3snmhrmasyHH0dKNsu2EMTEtwwuVgxb+xsTrR+k+
NBetqaUVpte/S8eMaUe7BeGybADLzNnz4mATHMcND3n9mdctvUMgYalSzQJbRHMz
EIVRbhIVZke6g699J98pHXPIH4ajayb4HTeRM6Y/2qU1EalqLvKmsJFmtM0Ouu6f
atyTW54/kOOE487uIjoA8LuiVg2K1ZaSknmiwq4vJv/m5cxqO7UTD/c0fCDxWfkJ
osmv/QyzweEESZKD7t3C0jrQz/sL7G+LRikE70d7mQxgOXgXEExqIo0Pcdtop9iD
kIwQ9HKA9+GxSG9hzhmdHdc//BTQGFdnZLkcvwQ0dODoSYgJPCc7W3oB0C9NLrEB
Lybke858LwadAyZirLgDD3Q0CeqfqpQKOvbdnEuTnuHgL2Oe44q1t3ho4j87kgbu
p8GUUKS1IYj7TgIMeJg1de5mCojR7lUQJZxiwmNk/eTxS37+PIJThJsAmAexDq0p
HCKOEda6qov6VlUcqFXdB1V+5QYdoQYow0afebQjkNhRX+dM0O59Zn+pr9paoGZ1
i5mNT4QE0TS//c5INXwKl0ZKOwtWb2f3yAqh5v0E2MOhQj+oZMZaTJatANL3ISnI
YeKx/yy+XcpFSiwYOR3sbFRlDmEQvW4mBfs37abPmUWlqENM7rVwcS2AmJR2Q26p
pVxDgUYCREz+vFgfYyrdsgOD7iVg/0btXUfqMbKRd2l+oP/qfI8oEmjJY4FohMNh
zEKINetOEVldSdPX6WlOf19tuAjkw3zBWynkuT2+s8hwvS24Wdb5CqRYvR55jS4j
H9lu2B3xPr4VSbapSbD4FivFwYYdGrzwfV8OViQM3YXwILLLihlodWbqPuoH+Lxq
DOMOtDot9cnRuFZgXjmz9zZets09nVk9M/fjI4v/wZ7T/sBFTcmGFym2M8FTqbCH
QwDZ0gAha9IFStNUyOVH3wJAyLVN7RixH+z+9cLQh0sI64aTBeIGDg9lNtg/Etw6
AA9fxSQc5ffWLteh72zXKI+EzK+nt0/XgtiaJuzEZW4tSwKBgMdDxgaJT9v6arKF
aEmG5CQg4aW/L8UMPyVQQiS4uKC02cx4+CzFtr43aja3cPdAkEOQCZxzDmIl03ru
PCQ21VjjFWBGOaokCAW+yKrBdv6ZzDyffAWxnN7BvA0OvRzbIyZuGkX92HTvrCmp
bXJw2KuoqkNYCkwVuZkn3wS3hcUhR5z7qduTh0NR98UHhjRiePRuHDpmt1eJADjZ
WycjCbPsphjdXSHugiv/gkqWt/MRXQEDqMFNzRjoCrWpz4OY6d0Nu3iRPyuuIG1G
rSCxfLllKsFk45mrADU9JzmHr5xeaPBKK9O9q/EO2eyVfrAO9rTAz6sbcM7PysOF
ffPNZZqbVIiPtGC8pM3e6h1wCigdh/oI8TaEvHgjSNHmM/8uQokfsNVgdAxF5DJl
Z3+zpni8CylVEhLPfMvJ3xsxIzMX0OIV4RonyVE5fjD24OgE3OFLQ/loQAeNlUFy
OCQ2M/oX7sU8HNZ73TrB6U1hiE1G1A6gL6YE1iNin5DWURZlOughOY79LnYeukpk
2lBAbA0ejqKCh2R6FthrUNURXpmna9tjmSNfpR+qEo15zzzdEIBufE9UrOcwLOoO
Dqe1NGllJJ2wHl2N7ZAsjZpa/hRBPvBrtdlMAk5pIkKTTq7KmQEe59Bnj08wNv4Z
QaoeWwQYQ2PRHw7AKWdmSF3DOds9RTPagU+Y2vnI/lhwnTdx/v43i0hbhUev49qW
qUzo0PVKxbDVEPPkTOd1a4ZApxeSlmrUlQSdHwlF3C2ynjbL/UslNwtL6jTJ4mTG
mF7XBrjet9cE0L3LnnTFTwncdmElWyvJvaK+udNBaZjc2EHVwxjBdJu1BpNzukR9
nY0LEGuNsCiFn4MkUbG+tHVwc8v5DN27FU/+LOoU3k9d3b0y9GeOepm3NQGf40LL
k6RmSsd6jHHUD5KwgfppnRhmMgM06sjtCKejAQHd1eprKSNxU1rr/eC23gk6GP6V
UYPteZe8TAr/TVxitfX4R0cDjqXt24tqj70tUsFj8GSbjj2OEdvxL37CnWEywVOZ
NKzyUm18sEVeeJQyeeP/UuwZzWDanJBJ6SzmX6BuxZYr6EikifSvu7ClMyvJCSzZ
gjiJHNJE9rzoPDDDSgzHYfMmLbuHmqldAb9oJCkoudW9YaGRUDw+abrwU9syhE1a
32aqfn+FLpi1qln8szNvmrJvV9HTuPn0QkcQv10qs4DAfA4R9cnRZwVJB+DH6JJ4
FS1SJM5TBLEfjPWoi1ruO2a20hv1IP61HczKAFw38CAvtmbmqIRGJP5fy5nMDYrJ
N9xQFEh7Dzd5kUksPR6LP6tl1RPoT+SuoLHbY6WFmAuBcFSv/0bwB4eih4bYhHMS
SHH1mwIkr2I0nYsJEFAe3IwCJ2y88nQ8I9I5CQ3W+yt5+t5kz+F/0G+XyDrlXXSn
Ikm/s4ef/KCj6wC7lNjbS2cRIg1MMrD40NVH33yludR2+54PredNdv9yKFbWXYPw
SCd4ljvvcc3oeEkZJXeib2PKiDfWuBccPyLmcbiaxgKalpO68xuYiTOb0amZOaJM
wPO/TtXKgVMGC4cxYJTfDYz51+wz1Yldb2/yBmHcCVzKAIXuoQUcvTzbwL8R/xln
qE2iZGl9BB5p7przFEPyUkXKwv+RMODfpu7tqvZ3KxzPK6HwZgbtM2syL+I4d2H+
ajLDwY+ckz6qjpaCZqg9WmlSkvjnVZqzugsu8beIM6PSkj2ByWP+MLTxch6ldZRg
v9B6grMHDovhw+pF8zFVqTYV0Hg4SKVF0G+zTuQ+bLfGG9QSsNQn2GEVQ1O+j3/I
CP42lM0Yp5qTR/bLtyP1SDqcz7wYUjnAH/yM0tEn3S5NJuKoJ7Vq93XXGJe5+KzM
+wyC3xEWXAuuN1LUX/B/XsJwZVPowlNWv8UDPo8d7xmIqmfL1n/umxG6ZMZeKgsP
0a7y+ZyiA+VH2kCXU91EGZlaCmgdfL50UvqU18jvrNFEK7mOsZFVCqnjT3DbklrA
8pgPUb3Q0ZMABzoTJjuTayB9RL9FXxO0cfpTKmwW4SNVqdNKhPb8ijpOafeSWHA1
zAkpwKIS5Qhcq/coMbVYqHFjxbCW8SnvQn5Im0HMUutS+yWMiZk3PqjtXn+TjY6S
/P45Zq+zNz5Z6Stmw0fZO256NTBtXcALdVsBob3akhYKeKPR3joZScU25hjOAHg3
Ev2RF/oyPA83CB++dE6YZa+nHhUUGG1XNLDpM/xsH+MXo50az0eZmvesjAT54oth
GHZTkGh5lavig+nZtMzVHwWQI78IS/LRg9X519R5dSlO4QhreAi4Totr+r1XcEbw
gm8copbfkp6toIpdKI5W4D0og9pwAGnKooyvN+rZaFYOPR75MyLdCGUv7sFvkt+4
qZMj2p3qcZHMXHkdRs/CLBFbqSqmYNST5AIUNwE9CBB7KCGcDD2/3hYjJqcgXl3/
96NraPUfMx2O3TtSR4R7qCK/6IFJwkxaAJJAqqWIK5BGdNwB/c78lWJZajRtLTS+
2DvEvBCUoOjsmK12lEi4e1Nvo/pFZMi3z5ZtZ3Qw27iYagU76ae5n2AEmnlterBR
AJyydKMr5S0KD9VBBbs0SMGDDQ6Fci6P3aeZsX/9/u7zVUU4Tqkof5w7NBQFpL2P
EBGJi8PNv5p3v5lKUh1GyFJBhHjHYOky7rNjvABbzQuC7C0hyUekVucaMJHW+ZhV
4vgLIuoJKOiMlehxRei5QduVM4flpEiJlCAJwMA90d4gVO62Qpc3xNzQRDa+5BIx
2pJB/jtgKSEs3QJAbJBcSX4rP7i9w4rq/lf20shMYjShBNfmiG24IPAVMJhh+4mn
zCvYWL876tYWVEAjIW4/P4OPX73bxoOvLRCQ8f4ikBJaUrjxZuCycBbM2AG/1ekC
3bSni8SbV1ruhuAZ6Wyyo17rXnk/WS0KDRswqTzzRt3rbZ/iHNcm6Zk4/yEieVlZ
TkvwZz9FQoxivl0tihwgmr3JNQBoZlC2xOGUK5wac1POjagDrRpqFYUf3ixEM7Ac
q42kAAIAG6gdFuFloBbZ4TkZW8kar/IVxEqHqPR3LC/MVbd1wDpypG3uKuaIkThx
YtTiz6UM0NTZxfNB85K3pk8fR2zd+YixzoX2WebZdcXS0KCeQeM8lb6boPsDQlrf
XwzrA7C42iKI+X3VNcsvgkY3QXBgds1qxbxYLzCAfY6zgxLJTW9baTHsl76g5p0N
1muAaVXLY3L0QTOQQoPpuAd8makhlestb1LT/HD4zkQKbCPBx5MVYYWU/c8t+QK8
IfNbJPtTYUTIitMlTz3Pfpgx7K/JyWQW0W+7aWbxIKly76vw7UehAvwpuSPJL7ZY
7EOc9105t4Y97Ow3fh/CSf4eWIMjkYjlC7Wu0HHj/5ymUxQd4I3zaXpK71276cSO
2UHRzGOr2SkLh/gn4zNXzlZx4ks3DUQ/YGAMkU3QZIq0LMHhs4d2H/zVIiFyJqPg
l3B5s3jOa/xCb3Nq6XGAzwAqQUimOvd972RepqjS9jLzqJpOtQTgl11if0flkAct
UGXxLP3lj1RpPWkvnqtilrOJo971UA2nsMrnskzNds6qUeGDwh5BExq8guUHLtW/
6Cn4PLerM9nuSza8JqfTVAJkvSrNTm9u+aIl1ORilbwQFR8v/17tdelczs5zMARQ
PmsmDW7HjHfLxYzFv5TClLgriCiP81nCVNneE7x+bN75IRg65HLvtJZQbcC8p4Hw
wdN9N5ziPUUIqd1il+ilP785eiLC/epYona0bfxWXwpmA7oFjj9Z64g2ohbc3FjO
2uHxiRwO2Ioq8XUq6UElWK/ODgc3NFyd1I4HN9j9yQjNdsOcIdnjJMij1OiAU529
cZrUBCqRnicuPr+DXyEsJrdxQS6Ja0yf9cnVkkicXF81zjc1QOi2Ba6Cj+tXyPuq
j7oJ9zsEFQeO+/GlEJ2aHxobxUsKMC9cXyFXwEreNBaIA3J3Wwdst82Bh0Rx6ds7
Ib8rFottXbgQsU2aChzVAPO0dPcnpgMAyrodeXCRV9eEOIY+YrYtZQ7if8vRrxCl
RHOMh+GEsvx4m9cHbTkGa597V4DpB5u4uOGD+3Xq5QH4+OakxWZUJxV2Flp+nZIa
lfVus6RA/C4hvISqNSnYuo5yJVyYbN3NydeUcL+PmDcuWJUtJFTCp0D7qlBAnJMg
nFVJk8D4wZRYLVCTaAn8lnDD8rx0Jr9GDpxXvFMhTHrExugOg6GwJ0HoI3ujE2+S
HEyTR4SnkfPTJxkQjQQtmm6LQulTItLKdE7hpD/S6E5kr+Cb1vajSAndryo7lxqK
+IYUKzO/a/VxFwgNeAg9aVJ8/a8WJi09mqMhJ7cpOAVcKp+6RZuQIbW4tlCYLgrG
/yChadoAw9pCy0ZteEle/SChBWXo4bgzJyxLPPeWZwPzEVF+me/UA7NbYmrHL5v5
qh40tkcc2rLpREBGVY5XVk6o+MJnpVwv1lKxFTyVDXVMAulaR95+WyeuSTfxVtki
id0JFZc96RIUMo2/Wy5Q6jLOTfo5pPfmj49pfkmuHLbyRV0thPZLlcSo3ivEVWSe
9pmCkXBu9kDaySB04c2rPMn2uU3ZnMg4srQgryKKOGXaJtwQP/PUTrn/TCc0eWq2
e5yLn8ApYS8fSqUfestbwc8EiD+komablFMVf6VsO74SoFjWfOWaPuAhBxNNJ9F3
iHkP+NY0i15T6IJjPj+zewNBpn6Yy1q/uQgKoAfLGtrfQRDGxXowJ+ri9+nIruOh
U0VPk5AkSJKYAo7+mHcQAmWBz55sYJl7TB/NeBiBA2ACxBeZsQ3yoX/xupAcXQmn
rlv6QXk8fXgpwgVzkWMD3G+4E3/s88cTCBYJvV/kofB70FNsQTZtFXY4cCwazFKw
OsmzEOUs9SsPgyZTzjHd+6Rvb8AMrqci1dXf0gFj9PL4IsY2SdUqQ6tsdqW4uIA6
uXV954dfXLLm4r2eNrnXbbTThK38SiWIFtHda0kMgjKEh8N8D06mS8aIF1tdBb2m
DtJmm6hb9LttsKmZMzTfakDF6cHPV+Dt251k6YuIhcZAkvEjdvFVgHEjh670mmCL
VWdu9u1iTKrMJ2odmj1PJUHiWZCR3L7UNvfht8jPxP2AaSmxn7mBtoN2DBUe1nMK
fI3oZQb9SggK4wQUWfrDEW+rf0RWFojNpZsXw5mEyY+sAE0gaEgCvUVkAV+ElWFe
Wb1TKHRHX5pLvh6d/+SyBkGjNDRDCFaBq4XWICDy5tyCC05XlXDtmRZv9Fd52HdB
XGsDETY84+nccalUIC4cwULvlZGNIjtWreA9An87k5LDFUFJ8uamoq4GRp56/PrP
qDcZO5bzYwKZ1l6V8jmjLHuT77tf21xcAJioISAGFo9C1jk9KthPuzbk1UJqX+3d
VxcvxDF8buG9AXVBupPUECfh7CBRhHGxjifduIw5UioGwRUXu356+HLgwvKWs0om
mGkI1JNzK0EzQEOiYxKn8B6LvtKDZdh4ZTfDm13wgbhxWica6dAN4IaL5zXd7087
Gc1BHNra/Fdu98qgeOEv2UpKSpmZlKrIpBdf9KUh2kl2SIRzY3638k0nj5/eVF73
7f1CUUl/8jXc7XKLgGmJ/8asR/+j+4gHs/lfelOj9MDcLzCqx1RLpwmZaD+TNVhX
Eb5jKImxLr/dy9bJYnNHQyt1gwzsK1OeYAR1nQcEL/rfBs7iauEUcFPNLFJEJxIh
X1NUH61FCf4c3O48fQkDqKCMVFNMEl8deykCyYS4dFTqI6NioqHXGJnpLwrwOyzV
Qxsxxe2YxOQpwnqPNXn+uEz2jkNBNVDCunal40gbX0fZUZoHPeOkoMQWmC+9Jbg3
5vE2zc1vRXBLAWUsJuuY3Ylecjp+lyNz+vl/JnZ4wJx1UmuirJH5WlDuFt6Sf+ra
OjEHhGLFBvNfdBDp2uvWzefu9CvOAv+XiE3qHWD6il4pqNlMf8xLYAGUT8z5CcAA
/8Q+F+sj6wOYJEv2Uyt/wg03R8bN9lxNXhaHA3aMrsaDaFi9Sx9v2inoBWKWR4X2
OXQh4K+PXAGsq+qbmRD5abRul7zNDkU8YEYPC5+J9mOhjMfEdHZIqYzf+xJ1N6rQ
xPhXpr1DsFZ95q0vBNp3bGIlA8XozaDZLynS0UDPPHTmM2PPTOh3VfR3EeCDsUZr
oLJH01K2ir8Ho4PMx93b4OxR8v9mfVmQwJJulKkitFO7WY8NqJy44LSR5CeuXWp3
Awch9m9DT7cTk4pxeOo/srfjfhTEv9hjDLR8/qcJQXAPivSEDpFlZKX+7KgSrq9j
UhnKvTVpcTKAYuRgaLGBBf60fgbmqUVeheA6raTYyKswHx48Lwz79ztmtkJ3n+K8
+0CccPEA+KPH14IY2sc9ujE6VyC6Dn7crMKkkuS7Ye19kX3aBqiVDotZtQKGDcNZ
R4cTA1liTTEQ0VVF2Bysxuq2p+DoM4r1OegBhveOUSSlX6qVqUy2SJ/6ulyu1YXX
GUU9Cfam9QWi7zwA7eWYTPvXVPBrohbmaazryiX+bIc0l/EmnXe091YwPtYlHsPk
fzlJ9O+1KoVy3PHtt6P2gDBewchLzlrHGxFGeam2f4HM9fSPHzK21E7kvTRyxCt8
N3Y6W/JwKanm0YruiPvdLajXyflj6QHVePPB0YBNRJZfLWRdAUAKGPxkdK9RIZM9
plPxMy6SW9p4CUjVkIE3aEVNpD+gGY9hy7pmsYOcDU4TIXz/WUYxT7owRAZQoFif
TA28oTFggUfDzNQ2KACNSmreNex01bV6yOMA2Q4/538cr3u+xdsVPXHD1A+ZDTmB
sSj83mpRAAjvnQIG3F1jVAXU2DSOBVFAF8dEbjTVnHtDBLG0D20/wuwgT71wp9oO
bKdG0plF1y9+AtiO9RVnxNfiOUhwyLzwlag8x4ttGS78rfQFa/9zWS9RE/Ow9dDz
zZfAGZF0hrB3L4dIM0VUsubLnw2yeB5CUOMIt/IZ05MRYyfMiFu3MqcGMaVni3VQ
BkMqIxGaXhOzrKmUT2UuAIzgfk48ljEcSvEiM47BcXPH+r4ckxT+5dZIS2Q/6kWw
OHdAfbAlpx1n09GPd9yst88cp/UAyVsNWiZZzSsnutXrAZaRTvb8b5f6NoFUZCt4
iOkAJ8R6WRFXTM6Aq3hSq0U++vNNnJVa7tfjru0XJmmEs5bW2zyvTCu++3EP+jfe
CAlw0mKSvpSU8R/V+CjsXWHXuENhMaI6PflvM2tEvojbyI0dLYYUvdVuifcIzuHQ
7a7F4SKlapCZTV6t/1JTLmUE1f/xGOfP5Fwd8GjkvSHocXn3NnWeihvLy5argy7i
w6XCTGfmKI5dhyRIiGXHvsUOpTw0/Hg7MDOuBvOja1XY2nEvZuIIb/RZJDUosmaF
8G7ghV69I/+dfUjQxIvhwShs/Qe5LnC7oNJujC7lg3pcmVXkj4WKZgESAaXkHYIQ
WcqIvUoG4MEUh/Qw0RR6hkomN2Pax81T343iNfzWLNX9ZMrb4zl9Xq2oBKqJ3PM8
HMn2nPUVs+HgLlt2PYwstT/EgAQopSnhuGYMZqU4MlN8fCFjzuU7w3lCrTsmubtM
XZoLUvTGp9Pe2Ful6ex+5iF/6HGZQ78yHCW3r+1tkNpt36Av/v8SshieeiqMifzM
cqn00SH8peRu48dnSTEHAWCQnphhn/6dkcz+8gxXVROz+q+vOIjAl/SZtluzZDOG
8tzMNtBfbeljPreolJGmdjZssnW0dQjaC2S5DIjQ2tR0snwaUT7QB9v/jJJFO8bv
w7O07i7kAWK++aYinv2bGPiEIkbn7+7NpZpeoVpKwV8qQ71uc0zFQpnS5rsFXW+u
4Wi+TTEfJI6PpDLtjskaZwOAD/r/cgYbd3XDI9K+NFxXbvwoYXyQr/AvNsRvTizJ
thmOIa6ReR3OCtDTZkvR9VGvXngjGe98fyFCvjnW4hm+wNVXRTBXRCGDg0xRfIgV
cqyGiBKiqy0RDKVpIaK4IeQX5kry8+esg6weQYqQoKqXq1EX/z0/kbJ0n4pRJc54
Tpf1YfRogE6frYtkj44nxO93IVWJZZyDxoWEzYtdyDCXhNxC5Oyv6xm9SD+tF1Aj
hQ+lSJEkIEr5BL334hTu9x9jinza5Y8sMNKsGxIgMk+H19ELQF8P0gazdldJHgA0
zKDbKJ8n+ldkZ3VrY+lfSzLVu5F8kDg48XFCSRAFvS+hplLBVjac5die/ypGNg7E
PDIIzw0/u76v+o+r8e0HGkVpURNsXBWTxJUVcKmJv+b2RLt2TgM6Fb/n91xWdOQN
ujFT0xERnxd+4M1IXPDz/hOiZeNB/tuken6aD3G+HyDQo/UpF5173MnMuyWYBUOK
cNdHJ/dT1/cJ0Q1shiclNUU1brfHIyo7yOvp8K/xzjY7YGJXlMpuwTANuw85p9ta
Ct2sE9gVJrlck82fCYzcxwoyLmmYOrIsCzVs0J4Nl9WmI3aB88A9/nOplePjANNK
QQWDIAMfktdDzITgq/R4KAxkYdATJLDt5VDTkRgzBXRu6ZDOUiit0dGSH59u5Rw6
bEPv9hbP1RgYHgmptqK0Zc8lUmkjJyPl3hYHwsoA5MZA+6veQLw6ZX1mzbOBozzN
ddYWKEyB6HS5QW4x4P/bDJqEcBqfW/bB1lxvsRuFGKRkuLeaFamO9uRtqY7iunFV
bUiDL61BjLgmUwuxYo6Yjlk0NLJDAxoLTyTPHA1rwpUMxMupvDa+S4Kak1UOhQ/m
Maibg7Iw8T7eS3pWDpRC2DhSFjS01NuXjuRgEkOzGCIexUWRC1sBi518LUimqzhS
sm4usNHy6jk1OpTI12qxM3RY08jjn3zEAvyC/g/WmLMMg+E8dAgRFeIwvafpz9FK
6XIJOi5+FCCwhgv1JLCDgVyErNxd/8vVJlx/FdksxfQksjV2G7GyErpx44IpxaeT
e97Dl24sWJk5+GDXvfdvomPP+gaVOP7YQsKKZnm/NyvKgjeDTQBvWLf8+yGcM9n5
WtftFiSYK3/iB1Yvjk+eBE3sHxk/Iljf2S/gU18M4JWHhQuArC5QWO70aBcOEvTP
KNAP2IbwulaWqt9LRftq59Qd0Cy4U+AOOODK1PxwSvfByy+CuNhepiKihnsuriSo
xsbjLPs1oIaYpCtYjh5eiuDnBc+KYvmMRNGzoTMm1SYRk5KDJbBJUqaNAwCJvU1V
xnyhb4k81MA922Q+erWSCdqR+9Jw0eku3BzsfsbcCRXdEcC7GI5qOHGRrX75omhH
t55tmldUuF3EO7lhHTzw9djybKR3xe0956Ol8JZAooIDntBvI+S34o0s8rZumHnh
mGoHJMTlM+LzaRxRwWMeTgIeEp4KvygsrspHlR2i3IMUyCMDGI20C4gyWNQZYbuI
oQ7KXoMqHyeTrpMIToJP+XUB8IlRRLYDnLousFVwpSR9Y2dVgnt75cHc5lVDVZSx
VG5lg/7dYS+2ywvssO5/9Hqlev/h+MXlMPbatTmRWE/SBSLFMqOCFzgSw85KAUJO
bbYT6ALPI0XZfzeIokNqFPeaR+ldYXYuIPPACED98Aef56o1W7/RSwlsb0e1tlOH
zeKKjixujTsOd1WG1BisJn2S/f5e2mUPDxmuhwp3q5uO+MbScL7So6jtNwztVItj
VRNsJ3TExXm6dO54J3LzsIL3CTjtH8jnSe1dwXMntKn9W/oowN2TBLTkAYOClEC6
8Liibavyu2Ye7yr+McovZ+B82REo2KA2UbURmRJKkNEARQLUSICezRdTnwWwR8qi
hOxxD49yk/l6x9tiJhY7Ce3cZtG6dVhGmZq0zoYGOG/7c3Y4iS0jvvOS+NoMv7JZ
DNJIeye4YokeTRl2VI09xP1Jbx0JzcXm+dVVSkeD4M7PEqWDR+vaXdvtNVLJ6FrB
ZB9E4uzdfuTHB0NuX9nad3XVf+WqUJIlkyHqodvcJm5UdTrOdQQx5QAAxw7IAfbc
gU3F2h80+hV6O2SMABtyFIIYiRegFLdwStt+/L5cmlz/n2O4fem0xN5Ta5TYR6Ln
pd6Z4w271VSZt341jqO03+gcT0JwBNjiDWZGpzVwsIGXU3H0xRKnrUW5ByxJEjNt
qfIIgbBrjBOQB/UiDaebSI2r1AWWJQ1iSlf797fZfJB6vRqZtoEpMnG+E2tOLDRU
oB1p6H+BCOQIy47nQTKYzLKkW3TjHmSbprA6l1Ve0Bi1X7+iEL6sXsbp/CpMa2F7
bChl9T7WgP5tw5/ez4qxS3YHa+GxaCRAyxgSEznJO9Qki/hzAcrI5CMn5AL/iSnZ
V35TzoUkFE0we0lpQ7Jf75ypWsGeb5Fu/K95dNpxUVbgo59k4V/ZO5iDoJNIFbaz
G1t3fVq29tYoDdYFYKL/S/Z6bK4jCG/y9eEw+BeDKP993pxld4vCwi7PCeGz3Fl2
7kI2DW4bs01qUpvhov15VbpvqLHa9DV4HyF6pJL95qF/7rZ9t/Jmi6oglWSwJOcx
nbCWzUV6hS0pk9NrdF5iNEStZ7RnWgxbRgX07TWI9r7VKO0dEqyULp3JjtYmFPJe
0GcE7xMJ9LiQiNwliozqK1q+usbPFJyJc3U2gsd+nG6XIlHYqRUiWJMf2DeoIs/v
/4jF9lmqfnelU9eWRawv6kEs0z+cYZFoANwnvgAvzlLYEQOQs46YddRnke6YLgUU
hV0RXZbvml9nqlfRoldh1BiuLSRwBjpy+ixwjwTjnUqeziN3OHfzcYjGiU5xzT/S
0/CXDZB7iKrl/QwccbEFTQ+zjlrrUMOpUJYf5fX+sXcQuI7r5v+tUp9+JtaNkVSq
5l6PqlN+Ko1YZSQT7Rv4oCe+7hU6oOkC35/8OiI4tmW8R9VIvEg8umg/RsefQi32
JeHmDkLl2NLlJnFIBGraUzGtMZnQSxgj9bBUqPIw637D8XI5L1r0hqpe61D0KahY
dOWF7Lsf9uRpG4+lRRLn+JjEJPuj8OafO8mpvjyaUufwugR/W8LqIFEeuWDAcsu1
yFlih4ILw8Bss5PnBCNB/KPx22u6hOexN4N0JjR9G6RQaqDdV5BrZ6Lah33UnRek
gnJanNjreUov2vG7nYMsR1N88DOyroRyf4fm1Io7LQNRam8POWTBjlzZ+vkYPFo3
NCIkrVOKgnjcmSS/cj9s3CCdr29NoOeeYBKebFqGg9eH30J4sodVOsqcWVX359KG
6iDagUm2qtBUCG3mIIoJQ+cpAAnlRMZckVG2MR0DTFAsI5USL430Dw+kTtV9PHFw
D358nv9jhm5srnKOYe0H+B25iOOgBqq1VxHCsoF1TnE+nX8f+5RwZG4NczZUeSVj
qi4CaVHeyebXqE5BIkOPHT+YbairxK1AwIcVF3G81cFKHU0OTbMF0Qnrs7Q00QFK
08aiynpyQmV+P/GfHP2GMvAgkfFtX2X3uv6X3bKabBML+fpUqMC68wnUpbjLLoGW
7Gm+kdhyhoU6Xl6e4iCQSoBSxx7qhTLwFXVdr7/jKgRPG+ppYCX4hptZ3N2pA9jn
Xxm2apBA/3OXXHMhLz1yJJqy4tZvxJMDruJJ7eQBSs0phv6yoFrAQIcWVPaz0jX3
M/eZ5GM2PJprz6+0hSwcG18GKcPn1klpTN881HfY7btTlEnzsOeTmnBwTcjMWsqd
w+//vTBj1Fltwb4KjRFghfy4sO8hhZRlgMQJf+w26oTF7WSSqhYxMf+GTFI2K5x4
iCRM93z066cHUn0C/zpXV3G8cgssRlM6oqL11SdLv+Z5SsmoPpq5iic2BM+6kaig
DEPO8c/bZf9J+0+mamG3WJrPggwvLzv87va4+FmSMo6n9+wMZyFCJIqLiGAttYhH
BfMR52ED5JCFzGXuGCjHkVJHPFVK6u5V1eSu2GondizIiZ/DtFXWhcrx/Z6/9wkm
HbzzcK8UEyx8bcEQ+gfJbz6wvDzyNTJfVENWhLDYhBC6Rg6RvM7SgGkPf8tF2kND
tvvUVdQzFIYITrQIxlSjpLH1SxZQiY36XHuLIAFcBO0tl/sPodQoqSRbqA7u7FVU
9ckoTtZKPWA4hB9JLdVx8NNbG6cB20znLIt9EtqEIUHkUPQ0FUhti42WTUG58aUp
OGAXI+RdMShhtYXPQLRjWCYzxu/uZGGbmchUnDVCDTkrsGkf06HIm9YAR8b3bIVm
fHeagbiifaADJ+ZRukHG2ZEpPZB0SGwvfTqld/LK0Ig7jWVdMJ9GRf1jTkkHn1Ft
3ndfwZWnaDoGRy4hl8FpEGS6pruz6r2rXggrXGPJrXJGNhxsC/Mck52pUDLTLhqe
VALZRlNc207z4Hl5036dEgQmbX96YY8nUIlYLOzTQ7ejcgidb7TPbF8LV5Na1JSY
6zZjdcJi+UWlMFlwkxr0ospAYYJwLLvkD7Qbci7aDVALiaIFZd/pyyWMdGgIHZAS
B3Kas9hfm9dspRX/3zC8O+iSSnPSE84JDiyZZ7QjIxH3i95EQ83QTKmPQdxyC+jI
a+9n/5lDGiEmJ+sZ7uTC67LLDRfs7o1mw8O0cVD7WMDoUffWYwl8hzzMiP7VKYW9
UsuROAdRqnw31ZPsHGbfkn4FS2NOEhTCHuHzYb3v6+rR+EQzbtroP+nsFSDPKy2U
nj6UroFQrnB9TJfUClHE1QNWIEdifcUoAadZYFMBJACR/J2kvupDPsLEI+scIQKG
CigSP22XWzpemxdoEzDUEURs+7iiN0mzD4fYBDTVRpr9dxL5jKC2NFUjnUblc4Z+
gO+SoXMO5253mR+0GCarpKID94ZszLrFZ0tQXqOq7rRgqlqAoFIWRVhlo38636pn
McrhTo4evtr6HE8ACh+/G84RhT3vh9ZBpKT/rrRlSv3YqbxZYPCp/ZspUnrwTPXT
n0gIZ4f6sGtyhEGco1ygTDxzHB7rnXXQKMJBrlYh8nrdkF4cD4lPsfeJlR2bVfeF
NTrWYgJeLJmzTQ0okf01RvO3d/O4tHCDzYl5yykiC/sLXFU+kLpvTVNPdKgY+g8d
sANZxNwPqclTsB4AdoIRXiCqseYfGhBawK+3t7/W47Dr8BVirpdWYRyY07Hg4wbH
1oqORkwHeIuJzXK9NXFRg3W/G6P39NzFIjzssRcYiD+QnmPO6v7j8irJyOOXl5D0
1SgTFGO2VrLfzmHvxB7UHS6cSAdXe4ITqeTlT38yJG5edzYR2NAJ1VkXcG6Kw9jd
SE3JPhIDPi6K1UrEQdtUOHdSyr8K+T1MPSiS4f8o4Rd3sWRGJ4++olUrzWVef2q2
CZ62cmhITAv3pyxdkHXVZhDnK9ykuddmTAlEwafkLYjTfznosvKt12f+Bp+h7HDZ
gJVxREgHZgdR9H5Tsg5E5AUakNIiZvD4Hlvj15gqwbDyhtHTj315dlEXv+EF/4Cy
iGBQU241R5OHUWXwiAU+UAa1kdeuiUY2tZQH9BIpglptvjZfZz0VEm93b+zOXJ4F
vwHYNEpGlqdv0Fyxby4wcc5e7sewoNpgid86OGlHeVDt14rj4/wUFoknVjfKttTo
beglK20zPXqLaPASzlb1plpG8B/+1s1gtjqiHwwLp8Pvt2hF0KWUTCi11t0LvGhF
/z98Zgr/VBMCO1k5NMFZh9t56uzImv/q0pDyVnfM261jhhBp73NXXfAg06aZG7vZ
rkric7NXUWpxjxN6R3IHSZ2Aua66aflOwzm2r6PmBgZb7pJ/Dl3/0iv1ma+A8ZSL
Nrb1XoWbkl+q3B3r8Z1xrii6u80bSNT1+NUNeFRWlMX5lgYfcJPRwWizK25nyQFV
pt/lhovgtfSuH4H77sEVOSr+0uij8/VqWAW1+DyLcq52Qbz13YiEcYHm0oJ0NlGx
7GFKfQjMQx2JzMRJDrmtJODIWWH/EmZz2e5UbOY0N946KnsDxuldPwLrsOlclrOO
YLBmx5XNiz3HWJRWrEtbbZ7TJSTdMpmQCUohdtAd7gngF//S904JOqleUGZDi0ic
D6U+XvcPaaM8CcFC1mKN4JwhcDgrD16MN9kydJaAR+qA1xwjZxsm8Y64o6rFPMhK
HvznalJGAi/vo4OWEZcdbvf4O1PG2499ckkRh9JucUffoIhlZtgcKLnSwMn1Jnpz
5sbLrDR3gCkZvIelgyvxl0AfO2oBjVLXhfh1xPGGJa/I7g5In4okaBNmSp8/Fkdz
g6OAjxrmYtTAZXjinHoB3EpW9ROFaCnFyN3w9vgEpsunGuZnbc3TTyyzRes2dNix
zLznzdYd4aCNRMNoi48gc2/R4RI6Zb7bdsuT79Cv9/6e/GVTilx8gBDN7DV5soFs
bg/W+hceITMtkdswnmfDHZP6PuCcoZmhzOoDZeJWrD6YcLjWPOKT0Noh85uU6h/y
h3YxuaAoHNXNTh+nLhsDeKgwfO76GleNcZly2XQBwMpeo4nFNJjOqoDcbwPkouY1
e4hVG1fblpesJROWUIbmpnGnD7JVpglEZxTNjxv1ADYUO7ZJj5SlHUJmTJ8CuyV7
lFcMba6kDriQp/XG64P9U4CyyNOtKC6KHl1QRyj6AJ5+K3B3skD5z7EnBFrxlOUm
OqJ/LXtqp0syQrNNOyLL/QcSa1TNbeFfoE53GoAkmD+oRPRIQWr1VBLdT5eAdTSa
gUUBqCqgMJbyeE4HK6wVdBF/z82eVbJmJ/NdBrhQtUmcw0qOObvJPV6LCIertQac
qM4JyGXFKqSC/UFp25YNlDLm7FBWI5F+NpywwQ0WOhNem4zuCUCN51YKBbblvpy2
CTUkXQ5gAA0zvtw5GwE52knkbFub/J0DruqSs0uf/0RFktnSwShWhp7NCAUMd4Oe
4kPszBYF69M8gb7tI1oX/Ypq2DNPCGMU3cP8ws9UC+df+2nre1g/UrdWMYiDiDwZ
E8z58CyWsKTHKY0lByvN88rUwFUdf30RtqO21ptOgu8l/7soooH2Bf3uDLJGZgeD
7yym/ljRj8hN928RAgeroQy4mqvBAJ2fAxhdGI9XXMFT/Fbez3B8SJhfweFh1EyQ
z9/l812RXYiiO7zlXpvSwo/Ok1YtQb2DEcZrgI6yWDiJT4D7WsCRH/iQle8kkgF/
U3bbWfLubezEgA1LG073l17ADQN4/tCl95j3jm9e6DfhTvTO2LBRe5/4fhrW5Z2y
xsmxrWz4c6bU+HXYIJhF33VVyYyhpa5HFsDW+Qv15UkwtsYRSeXvhMagJsxqQhIJ
CrrvSTS93h+oCW2o7rXCs92PMqm7T9ocPCMX78NBw6Y7fgmkEfcvgDIRyZxrtBfv
LESGRVF9T04a9Y8dWQoEOB9KiJ7GqZwdpS3sAbt9pt+Fnteej0HSPO80PVR8SzJM
nA/3TznTSeS3BtyRKWhTXqUice5XBZYT1yv9UgxgA0mPeqJsbZC2WL4zQCj7X0ac
hKneNZXUhxJpw72/ujaFwNiLHstymaEVFtqMdIaGIgVTfyjFL5w5wJhMl4+h2bdN
kW4xcQhJuGfvQKf0PEKn1LtGh1i7VrC8GmG9olYfbUsuLdvE2SEr97g4wCyAFc86
mZ08C2K+1CXT5lUPOuoWqDuq3F0Ty7VsEVir3F165ESSDz/zGyYF0D2tQ/XrxTLf
ryL2KBCmDdBAJsxD8cxp0pLvA9FtZLZL0InTAEGTw5DU3aI1Cq2ISOnRtJjXTRiZ
4pc3bUaMzcsQglJP6nNBX7lFaTpKHWDrMz/sKnqLTrzSU3PXBK3xGXYP3G4IuPj7
DW09ahF4ut3okvbKSZjjB5YlfoxRItxYRzkIVSgyEkhTunMZXRX65BhWd15CSpp4
QJC/v3roiMVKGVk1i1ChW0q1Z7VFHlrfXUaNjNWJ2/+K5jp18Z/Biaqnl3QX/Jas
YCn7wdwxuIyhiQkEF9n4JcgNI4akmATOYfIPy7cUaCscyuJj7YlJq0txOufUUShi
xf+pUeOr9aUWjLvlzpMZVelv9uS+iyfUDbz9TTBsFX3uU5Ee8whMTg1oPQWUx6b5
ocukcUcpJSfI7hB0+ViRROLWfQF67InkK+6whoJRdYhwSCxXfmQYqsdM3zQr6RGM
Fesfj5ZT68ZOqtYUo+1ih7kKhg8IY4NB6VVzAWUKzySl3qmMPl8eSYDSzSWX4edq
S2dFJE3c38PuqQQA8ft89HCwOuG57LZK5CGadacixNaux4Kh+Xik9ZQ02jCpZJ/x
3OyhWjGLWEbsNlZt/lxN2GlGl0RDjc+BuE23JVlXsmoIUszfN94hqZT8cS7VeAMR
LI+O4uF8WZgJffTHWSuTo3+znbulp10AHQufuziUOIe1DKzT3ZOH8QAcy1V4Dnwz
ACguEQ1FzGs+1dWuWrlX0QQGV/3+3RJDS48BnLaRsqqaJZVNSfJWzh1V9KYP4g5A
UCAsvVNPnGSaX6fd6CrJyMRKCvLrwJxifJpKeEv7+o2/8UjkZ5iyhvLsV0N76lYP
Vz7BbLlSmL0tXuPqUZRMM0bdIoTj2ONggRS3QF15OmPcsutnlpQGfIA6l7KQ/nq5
6LpVgjNX5/yYkdBosJW5xEu/WLty9V41P1gXo6gr4n2+lIBH2DY/Hs4ZD0hSFxAW
6jmyRFbSANC4TLxwixOco8p3zhucHs3O97tIvRTWCIHYcrD+6PVkVXtU7iVulGNt
gBByuYqp41K7Gteya3uichJaFCUUP2V5XlAp17+vudUTclwmG56Xz+vsozR5Fqxx
zFI6g4z7TYjF8AnvPcDDFlyx3Nrqdv/fRGt3clZ5BQ/rF2PZpS1EjEbKlZ7iwy3i
ESfeybnCBGwoC/GyNfsT5upCNYQvDbQe2uOmHHai+VcP4m8fbG9tqDE8grxrfRYW
mpDiUxlUyhkzv6b3I4d2eqTUxMcfUeHPTslWZwCn4wEBTtajFGeWZX0FlqhT354O
6BFjYr9GLOnfgn4in9rJNxQiRtaiCJ3LLt5TaUGEhHzhqmzp1nc3IcmZHwnOXw0f
/eM34lSj03uTXd77KhIbv4Kc0SkkcW3+Fd/Rvl3R5wkSRp0DXbA1ZhkLGIPTzDTC
Yx3p6+L+DGY7RDOwJTW4tIBVGzIVs0G9n5ekIPxWX/dchgzePZqni4fZE3wt6XTE
zz7rnfrbQThO5oQQ1Eay3JOqsNU31sj+HG9Xw11w9hrQ/7+XmOKkiffXPTfvggAw
KIEQpy2zNI3QOnJoYvsPZ9UAhJDXr9hNHPkXcK3/Y1oF+Rn0LbAj/X1zQlHA90tb
1XTBwGLWnIXitVbaNnMt6cz3MFhn9EGU9N6sb+NxYkZHsSgZQv9cLxdXTvi7C35T
6ZoSEPnVRZYP2QBM8hgivBvTU1xd2AdHyrKcOqKiKbFdyYxhHziHA/fxpdEAzyz9
ZpJV1LlOwJyJIsxtct8Tce9qJEmY6BskFgeqaZNpogTnFDYRAyeMuJ06F9NHTeQ2
CcxwpVXPTOHz71M7668t853ywF7ydHcTBm1B8GpvjtZvmU62bKXol6A1saryp8Zn
rMj3ev8ELLhUUx8bvRgF90ZZfanPInYdQYK/QNSOFhZiFm0l4wO0jmPbu8CRbvfo
R3LV8nK3A9n+I6ZLmC3WL4ZtQokHfrdIzU5Vaw0GCwYUBOSl9JqCMs2dGBJK+iUU
2CsalTsTVcrn6+zwU+qoTOAcQWibJHXs80InBxYLKEyS0rZ8vObqsFS2GiYngVaj
YCS13Dhshoiah/nt4HxCuOhIHK+d8xETGoKHEa3KxRyYL53n/yc50CPi6lYgoRgT
ucyHko9i/qwLO/HMWprZX1gjY7yI0ogLDJ1Jg+iqxSkCWLobgkWNgU9Ch5muqEZq
FM8XmngZlYD1AQwkA9Ek4BJUSkO4X6JSAbo6OkXYeX28Ck83pK+EF0tVlAXgiwu/
v+HYZQC+OL7X8sojmaug0ZPjweJ1UALO5MeeaR6p8Jn+IrhAjgog+L9lPDwSxKSp
LZfkkIuKRtkZ82b4kM2OuldFa9RZyN0OzlnHwT4ejLn85PjHb1HWWmieKrbXzRm7
OT4mZL9IuQb8qLKmynTcviWzPqW58UAKg0VmSt2VM1Km6sAFoGpS9tl8OP/ma9yJ
tM/EJjEK6shB/QDHgOmUsqFG6zXQuBTOV4sVvV0CCJu+TnUtv9XCTLURcQwfJw2P
MjnoaGLifoNmbt6cpTOqk/MJS8kC2RLD2M3fHctY06q9eoX18A9Dhq0QLMaSGZ94
mFdULKpTaAoggeDC631sZb2RG7ECPbEeTy9j+b9fhauARiU6Y0bWjEk1mCkvKToj
NJUlGlVohFkx3ORd1g536VTriG4RflCa5bD0h/p59Y4lkninAFoDrKFBv3eA6Evg
YGgPhMF/XRgCSm8msYZ9nb2/hU82grR9r1Yl7fkK47E8RxfceRA6nMxO+gjzM7wc
a9+4jf0hwzQZ6k2xKrS1R98r+xedZiEvyBMnj04swI9RxBZ3SaQHQc40N9FPbNlr
+wdBt0NMCG+gxN+os3Dh9FB8+9SELbnxwmZlJcOrdsNYsviyhfYYfC+mPPVw3fXu
z++NxAfjI0tnLjJAGB/e7ZIDtAdUiLC6XCnSVe3arJCXrEky+RuJOp26RTHGtUTl
HgS9S7WDyGoh+M7AZ5Z1Urdt4+WEAzG1nVuMoGENH/LE6IFu0OYfdM9b76Hswris
S03CIZfzds1YEhYW0h2FKRuLu4KXzewTXs6V7+xRqbil9uiCsb3/d69jbLUOloLS
mPjLCib1fiq179yic1BnV2XutO7WeCKM3ONmknanE/GUuc4pQUPu81IP90nSP8Sh
0F4VpALN8z2iAsF/9PDlCs0oeXwhjsVkIDpDeN04I4y07ey0UNIdCroUIXd23lN+
oTx9SbS+AUBXgsrKZcNBV2foE3j+4xkmoRlS+aCFXOVS8ZEcYEpx4eJUNd1gQlD4
228JWtHIjV7pprlRO9A5bvRdzI5yclJjCJ0UAWqKqkipIU4FXRMkOhoMCgzESK3x
2ITFABTIBdz8FhaxQ1D+2SOn7CX/q0AKtd+fFgSmNxQol15N/OYRqkhn5XZeYZaM
w1cm5hhCi0JUt6+iEMqk+JqCDsJUB7qN/71GFbwhCFayoHSYE+8/beajzfrWXis8
4P19v+RWwFCV1mPGAKq7oTjQbcV6B9S3nYSY3LiycQfku4BkiWz5i6hg7Upu3sRj
+qTBx3wY/nKX6ZaKKdyLiax7m67ghpp1LlrNAAq5UpqHRj4YmFD6pKebLy613MHS
jSPgh1vaKGnWICnAg0h8C0jOVE9ucnP28S+FNdDKhmmOU1LIChon6fLGbZT4iTjE
Ihcw118hifTpvHhCEs7FxNtxORwZ1arQeIRnFLHikkEmzrQwUJhjSmHuW/dstBJX
1vs7FL3rYgUDF5PtxUHuPZQMsg0IiLiM74M5XLtxLEvWc34NwDhq7Rg1l3UAkrnq
iO3J3xQHMbYjEOErTM/Js5ulW0F54EYFagRa2RAlV9XSxyEFWEE6tjDvpDca7/1F
7uYRBOShaTFKaSNKm/RcHGBjggS6RfJH+LqIaTfMK5J0JpSSJb05kAGCokJMAXDS
fVjZPNvBVCwSM4DaiVQjM4R9qzCQ3TQpquN+6HzpXm1I1FZNwVsOchUpSFDNtVUG
8cVASQ0NEpLz8NpQUvadvkGFg433r4MzZ21qsKgDEgOlJhIlk0gdJMVSZqj9VkX0
7prhQQdB0O0XZDkiSu6TSIAkabmXloXqipfsGhufqJL1jrkVxg94iTpszFQfUdGh
HCxyzOv2dS7in9Paoi4MJ8JER4ZTMkP2rg7fSVY4bTFtn8WgYTDWCBWiaXTYoYVp
zz3h6CsjF56wLfmhCnH1AZFOBZzl4iMU+RL11m1m2u+Fwhx8r1TIHQCySGZJcCZQ
qha0lkpcGte3N/HRiSPp6QYu/mL6fZ4rXeCwLznLZwWQauvMPlZJT2rkCz6pZFYJ
W2+82b+6HnNLyrOVkTrhrhfLapxYiCupbX8wch6iD2UBm9SzUKWJg0FDUlmqAXRQ
6ZKqfOQMmO9J1TPnzrH2u/6hoOFHzvXw+5Qww+IjeeWvDZuDi6CPpH+0IhFDkqtw
n+xPEy/DUMQ5FVlDDoQNlEJpE8HU1rKxts6TZud60JIY79J5RE3vtcFZ5qsJbBdl
meaWOKjxv7vQ/mqTcV/V+XjC9cLvexWZaO95+rBlPlQ5s4xjpTDxB/hCzt+W+119
VZr+Zp9dUjz3MxTWM+4ixkNugJhoaLbe6L6VBwqnz2QzREMdlST4wIeEECFokOqQ
WRdxOQYKOCyajEjCVr18dLZQysdZnkR+eVAUKltyBRFSssSoLmrkhHl1B6DD0Mmq
nTa/FrHdAWBrIf4Wr9LTOrxgp/XH9XqpsElnvs0WdwjgUNkOJxwy0r6mrpuLzJgP
2r44lbhanGFxtNUAp2PqlbPq//LPymSRusV0RTu1cpbE3yoQSMCvKmIBFrENfbpj
myixDxwUxdUMMjFzlV1lNmeuf0WVUiQRKblBCrikjOKc3qXTkQurUGhwUEB1Wf4c
CoZ4YH5cuYHA0OMNkkwNjgxAjQIK46LBul8ZKnhKqW6ZE0EINeN2fU5Z2Nmlj6Ki
vUW0tNM7fQ4eVFiz9R+fInDMp50JWE1a/JiAqGwE63qpCDHUOWKKMjtoItA0m9bT
fKtn+rpaVOwNj8Oe70YwnN7+BrksXSDrt5KlKmXT7FizQj2i67iRPrRzz5i71sqd
w3vZfEfityFIzrbKd8MvGCXXQR3t7t+Ugl0kbLh+xJrNOJ4555QLwmNHx6Uaay8o
VKKF8O5y5qyayEC9T8hV+rzI1lyk6Rgk76tLQi2ALH5I/Wzpen2Yo7wV/JMxn+JP
jPhxRLy+Sc2uTLclCP3hH32tDx282eBpueHjN+s81FFf/n7MbJGgk6MY65R416rF
2OcIG5G1IU+0QUJY8rQ5m0DMhza9naPrAyDw7m3N+2HLTzHMvKti/5ezuUJ2OB4q
hHFevctZdEkEU3ioTxLIIBLDdLQ0uNlSeklic68Teu/b6hpvGYHtZko3ge48WWRY
x9tFU9A2zuq8c5BbYfGEDGzisZxMwvgKyHcZvHM6S0tpilzNsKGncX+Mz6yleWVp
5O2H/EzFjVGb/lI1kmuhh1Jx29hf0kTTosezUY/eyIHkxy+A+0R7qeswblGgOUN9
PHIwDjkY9KlAjRCr19rwa5yCuSBZcSKJfo2Wn5aZT01rjAQgzcHnFZTjYPaID0KX
Oe9RoF/uJCxtTd825aGph/f9gtXb+cihgJfrUw+bKph6udQbFWZNHFNFcPwT+W72
Fk1kRpAdQkAIbokdeS7uU7evvuGFvZg2PyRIgxUT9aLjLKcH3kUJYGJ0dTqpj13a
UaWAwK/KRAxWkuYhLNugxGigcxJrFmTAZZkri7ksHr9KMXD7j4t8GNBhlloIIphO
Mm59cIICpJVZqCKWD8urKpDeJ2TpSEqz2JDxWeurij/wkYhbZ1whltypDZUIjsrC
mtasUurIUARECbV9D6JkrF252+8AKhorxQEOtjMHIVPWAgCPgGmIVmWV51/HmJHX
qFOZ3xMsVNG56YAmyqy7j/MOpUsDGonLbwqCvhmkSk5At8bfyjJgMs03W9U8MkKS
McBZwJuo3hQZ9zaPDpdfXOoMy40dfyzD+OGoO3BCqWpc0EoReYKkrPvHyJcMXLN7
rdnugRWdwaF8l7hdrOjkvaiFuWn+mb9gQRCEom7EH7Zxc/BYqennur/9w/BKkgFn
zLNaz1FVriHarTsEXMrkzDG8m1Q7lNfvvste4Pt/n55OsL+uqLfC3Dj5HIQgBqHz
F/O1819H4YQQi+kmA+jRhrNLxOQBMkyJauk7ohDLKvEJzRDttXPuSg9jdly3tQUX
AGK3davPg5dvVjfd3UhFIYye3UGzx4gJs8DrF7yw0IPyVTxRcrYf2AGQXC9K/QZW
JjCpTbYCeN6k9kvgGSsQN/FD+7K+s4/Sv7Pqpi/GPdEb+SCbQzII4O/WVh4FQGO8
dHF3F9OIAOfbLhL4KzsuwnfCMNHPSkKQPDS8DfNH4D5TQxat9seg/da1B3CDndOW
Qv57/hb3Ti+idKBlyUrQnzjjuBdu55JrqfS/h2kO7rj6OqMF8v9N0/zaqNncMdFs
mWCTbpWG+kLqQgXe4+lLKgX0HiTFWgYHdSOnWbLi+A6+04y5tSc7cV2JGw8gwLaK
xndOXeu3x8mjLSWRDOVjMSPyGIev9ZcwtABQwdIKtRYCnMgqG/8DSJc9MFJbMEpN
ijRzlelTUKrKQygCte0U22ql1R7NwqxR+oKZuyFH7A+1jxuoUlNw5XBD0RlPt1u1
AKhXmYWmloddaOApPajG4OYm085VYDIq4MTfzMuP/vGGQxD06aVLq+UW7APVkp9d
TdkyGXMMzfoevlJ0v5WlDQFVLW8tfebUORtpLVdMHvVd/aISqBR/qz4n5em1Ow69
mzbfhGwITPD6nqOJNbWNsYpwzHkHtSgGP8pcl5FtRIy4zSuCFUuevBWaK3/iCYBj
ew0uC4I6F42CNx8PYHmQYxpbbPkHQW9hUYxymaaKfzNhn2d57bKMEcaOgWzSAeR5
fI5kDgcSrQHCQdgJLNL9rQbrScRk4nAQb1HRM8Zr0N49+hTFBiZ6M+tXsBXmBhwF
lJqLYj1C/XIiKQLhheEmOiH5kIBVqJw3AFcSOerliWavpCFFVvFMdSAHeqXAhh8w
8Ob6j7gxocZeKTB+LsaaZFn2MrUfQYRowMcW9LQ08yTjx9XqCVGcFY21R1vo/1OQ
dCgDWQVDxx9tNXVMYP82CPUTm6FQGGALW4Hqmh12XYNj/Nbq7763wRfviSkfHdXG
KNVZsedLUO5kIzPhnEdH+tA/Vadb/7tnhqe5VY/AevipmGsskx3YVGc0BW8dJ1tB
P28ClixKnRRwvCSznqAh+GohLKOie7MtFkGBzi3XNmxH+rv9JipPQnbVkEaBaBTp
VE4iU+wksC+cpiFuKjoRv6CjXTwID4JVF2KESbhKV/5VjR56HZAf3LRNx/9H3PU0
H2KmWpWHBmGl0tffyUv1a6S/mbyP30/7b6geRYhcPctBECotROOGQ9I/EphJ4Aqv
LMHlLtf1JPxNskKEP6NQNj9F1mmqHU/jmSBA5HsqnSK5+nPF7Ka3l+UrT7BetAPr
GWKOY0WEj6XCIAXXV7regba2OcviZsewLKVvz1uOl4O6HeXLqSBodX0MLttPlomi
Sbz1/OXpnHjgwyOkQN8mM5+uJ/v+3yrV6ZaXeab6HmG+Ngngz5w3HzkotdqxAf/t
Zh6QsjZX/0NZ37unMQfe/Vp4ZGkG+opqxrhvGOvVUlPPf0m9XJeYm0dxfiHcft9J
OwUV9EB2Zs2Xi/q58nOz2UasyrJNidHyPzt6I5mHud6TutdooalyM5r+A6cSs7xe
ZtY0DA5i8QJEDGUpbsQxtg7zRXSbX3hTAq+rBpkKkVnJDa62gGo7HLUHXZG2/at5
udIPppIJkhUilyeQnMeI/kFisSipS+6OtumPSUwjltUh74j390n5YdMEU7lNZASu
DFhK+jyJNcF5BwbYuBwMRxN/99SUhOa66nkaFIm+oqjDNDA2+oShYggLVamFBHvz
aTYgZlssI7S9hmmVC9evojwDbgMxQDQTxtNLyeK9972qMxiRVJbwrBWTGsZBUOuM
OXCUQt+vipIQ/Qw1dsdj5240JiI2Ey9uqcflV+67bbpbsHUxOK1BOrBnFP7cUxra
qCpPctHjT8LH20GJVsbFS7WjuGCJeQkHzLYNIhZMVP7eYZ5CQFYwJy28dYvlafT5
zvCSkOERZ0OihZLBMvKxTEdvsC282QHIaKMx/rzE720EUauQ2oOJTfHLhgtXQ9IC
yyYYKVjYP7sQs1RQR8QUlRi3h/zs1MKuoY4MvF6dAJcnlyGaX0zvre5fPVAuLu2U
aBWBkwdRRhlvhte9yk4mYemvGVNXiUFgg9qFCkXAhMr1t7T/c41BgP5u0Mc9JduZ
088GLMPk8QKMtsyAg+Y3GNiDg+bae3jMo7QceuFku29+NFmQU/I18F3zqfB/pW8g
e3sfC2sRCCChP/B6m5r/LOYRjf+ko6o8LKAP5X7eTS0LJFzKFJiHyawGmLLbHDeR
QFSym/WccqpRnpIpV8PR/evtCMrRgzLRNA+GYc8xzW8CrPYGYshqQ0plEoDznvgF
zDxgNEW9RpPjXvQ2TCPpaVpeoCRlniZz/kdI5/ZI2kv3Bdv+z0M3nDI1i1wELj0I
qA9PWZ0XXUuQsfvDmwTGldCPVhsQqeTCLv+gVl/rBvU2ciyvfEIy0ahjiATGwoFh
ejal5Eq58CK+xqVjmCERJf++KFyFKs+KOVwrhAsHbN0Qw/MqHXHCMdgwZ/tg/JDo
APlIOma+Qsi56DEUoq3q3JU0aG7BPPDoETmfvFEZFRRY6hRHLKRJ9VyQwMv+8ZHl
nIxLrDJ8E4RSD54Bim453jIlE+KhTDdJUJsZQGP3cXWkm6186v9nFVkaivPaytWt
LCi8XTN8IpktwfFQgE9qlhCfliaUjK1yAUUn6jM3o6/nBITKLKMjeeOa0CAaz7QI
vY90ALn4dtlUGf8WYZKZHfcWdvc3OeAe8DPyI/X/+RrixdDsFo4EwoF8xrP51puo
ZNovMR4blYRCl3G9GhOmLSPRx2DJNbfRSmh7U/jXXNwI8ulahwBRj4hBvWVwdMMe
TZe1n7pygzCVjd9zWoYU+SkfV+23DyU44s/uKhgL0JMZEPWwE7pWvsIC2ksFp8Lo
0nIGVjQNT8tZce2LgEPVW5+NTP6NsvJMRv5nPq8QOnjaut7L448rw5B9r/j/axgS
kr2FyUH6KmF3QHQlpZthvJ1VnaCGpGp4/2WbTZmUa1qZHdqu721orwI71JRwAclq
bicjnUO/5rLw35jYZd+gzGzrT0lB+DKhJ2oPVq4XCo5k3+9pUF0dnF211rNHpw23
JX3iuI3t/czGx7WYVl3W9rYRqe23Srv3FomLN2+FZ1irSa1aV1aTqqsl6lP6XYW4
7ckA3PpguHh6ybPhwAVU4TQVEmrMJAKrv9Hgmfb496ZrC+ndlbpa6EK0f+ercz/F
yqjayv9uaUCU0Wz9ywgGetOQYI4O4t6XRdiBvh3VCTboqrWMQf3yoGb5xj+kYFWh
X+8Zhq8OLgpqIroyqG2nROy32GfTiCekdSVDEDc2Kgcle9PgCdPyHiS0yJmiAiZf
hrDQ5HvX0b9wzNQcq2dZJKfHtEJNViMd6KWXOodTiwJk7JcBFRWIKO3AdkdwJzn+
yDLODIO//mNzNY9Q7iWTYNwBAgy3tPz/Lswxpey75rvtPvE8o5LGSSXPZ1Rzd/Hb
l58MzUEjl7/h27W31UNGm3HIoxlfaLEDmtHQaxvLp26EZYtQ5pCDm+3C+TKaR492
GBLzr7vgKS7M9iXHbpYU80rn51aaH9xm7IclbW5B+riOjbYW5Oy/WMOR9ou5chXf
MCDODV/kqfOQPJ8NoH65aZoUWqD8nKCR30q75WglVPoJjOUZu6BNkdb3COetDZgl
6w7Zmy9zvuvE+pQvq9zYKoGhKf+8IXT1PXFDe7F765aimEBQuLxrTBEbayCEfTGb
7UkLDM58w28SUHVEZqQeAFl9uDKHHtwyFLOfHyVx3pefYvGDdH8CLT9a4+0U62Lg
VNTKjwAnKTSLb2KEAbWizmq1hXAl96z6j28hmmrZBOL4jmFcrxsWqApTdGTkXkIT
fvjtpX7h6gGap87yrYgI+yb7+plJ3bMWHObaTgh1D0Tb/qqi8HgYF8ulSBfQ9SYs
u+tHw2IDGXRGIj74GDwAJwZanpokAr+NlSDFLeNxAYrIQoGssFF+dOGLdlrmxlMr
xo+meRA3AlxwTBta5D7ih6wmxzexyar1M7nBbLtT2GjaZEt5c4VOSl4K2NukrFgg
oVSjlVusbiqHQsHYXkJONWEcJITeF7jcaoLIRHMoi2M6Zs+Jmn1U3IRxrL3Ot4lv
bM98SND6oyCz5/9AKVqJvXVFrUsuoWcyWfH6QD2Jk7Y6Nj99mOGdSCP6dMtcapCG
EjLntm6HIW3/Y0EKQ61v2oK6ev4/ViVQgvO4saasWccoOHgeC6rqjthIl2RCeWS0
9bc1i8gJWKtMh3342BwlSkAsBtvjeDzRn9jBXiOVFq53f++igPUPgs0yb5MG8HFD
pABI1Drtu77aNmUXZ/6I5rzAFUsesgxZA7vrL8ww/dQNyjz65N8H4xIeaJppu3Mc
aO98dWlBabwFStwRn8IWyh/LYBSIcN3u75I/eBXHjRjdde0zXpS5tdl4wTMYwmi5
EpMeSDW34PuGZ31mxpDzOV4pi0Fd/3ZXaKP7Ol9OwYXOVqQRaACP2dhQpiExU3tz
kN/tX4DiGEQtrZbYgOiQeQljBIp8/hPPcxwnhcZHRqTc5bOxazIh/ENycrUmMJo6
nueMv9bFV2p/6wupUg4e1HjXyatfAS3DryQJ+JJ+dSkwj/Bbzf9N4p+HDoJuo4P/
TzpxE+x3JKMB9JcVNyn4dMThDR/WdgbcPt9rlxpmXUtjV3ncC/yip7PxrrqR25CS
Qn0wU71kxYVm1tGtD9Uz4HGXuvlX0WYPN7mGPqxNeinhASMSFkXOBqOF7IgvpI3W
BXgzDOYDWt1AnURD6B09YnU0GI4yzmid/vKVyDtwvsRI/G4/Z6AU1WKDy9tZVfTv
pcH8d9MlXgotE+qBYK3+V5EdyF2tdtOk6WzQbwLyFvIo2fDFylw4zCvmuxINaW17
nh73o/ouevRtiyXY124GBcbGL9XsB5D9ph6rNvmCgsgkJ0sLb60lDgYfC6OgjPrE
9oQVs9GVwqNM5QyzzIH0QfzJiFyKCEXH8YDBzIM6W7gsAYyW3S29BesD0phf57i/
J8/iNLgOSIbg2IsxAbLxyvqxtCJWNkb0C++HlnqJy0ZeC6891N+8ZYOIbONVmD8E
QWBROJjwd2cc3wdzcntn9ilTAaI0X82IAL+C9OsfDdpBPHPeaRB/e88locAWUBpe
N5i3dw7A256NpoHK22Zf1gFXlotO+i69JgsqNUWNB/1tMwOUN6mfoyPtTVSpZycy
c1fsHH4rUGpSEX086ODQME1VRFoVR5LXqKU/Ox2RX064EDrWutfzcCmbq4nwTd1E
XZH3KY26XLkEKuQZ0BRsirD4fpxZwH2h8H7wD9eF24ydm5UXLiwUhZg6y/Np74kl
OF0UjoSfIMzg8NfZfAlqW53wPAgK6iefcslqCamqLSvmeY33EyqvtPQrNRA8MR40
UlES8R5czzCPMNo8Ajc3Qp7VSFilvOMwCGtwpdswmLnBwUIDEhcOZQBTmkRr7pbv
LZklpi6pM4h1bm8Z94GxPSy5bLPe8fh1j4rEANsgkbrTF2YGzQTrbKlaebGTaMyr
CMo1byQVzHZzSwnY8TtY4rtaMym9TiKLOCyz+q6thO47MsKqwcM7FNELntklU/IQ
BTtdbehi9KgZ36mpDHJHhV/1fmZCz929QGVll4Lg3ozzicTFxMy7CWgfHW3zeqcR
CCr/yFdljjE5fEy6i1fZTuWVdTXIdAex4CwSuB3PSaSCz+uG7dHoSoRxXiUxs3DQ
pYt1UgK5OyIK7J7Ku92zhpo0U0h6IuMTJ2UNdEAq9ni/u2FkvUc165M0X9pRSIa/
H+UobP9nJ7SGKGAWB2HMytvwmhgsn4nQsn4SyUXEaMePg04GPBN2Cxl7bTT0v50f
L8Q5PzlXdeoi6WzFsbph2jOh9kPUf13GYDuh1gkIwvLKI3eKyoZC0WL2GF905XyY
RNzAcpVk3S4dqae8ZdHUY7FcOA1cwWQ+MkMCIBErtzgMfsdhANXEkLj92dy/ECwv
VzfNbskSWqIU1cpJdMRnPA==
--pragma protect end_data_block
--pragma protect digest_block
t5AdjzcCaZdSBIC5dZxTKe3t7JU=
--pragma protect end_digest_block
--pragma protect end_protected
