-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
XnEYBKyKfAxTiV8nZpZZT960ZaYXGkPr7k887dgqdlMFf1vRyqhLLuMrvvrtvcYy
VRJxgn6pxECSdRs0EwKsaP5QZoyZg5etp6AHu4QTw69gekaSrm0ipoa2DJYwTfz5
FPJJoZ9pIwS8gq2Zp3o2J+mb9bACSwMK22qv3tf9jPI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4530)

`protect DATA_BLOCK
7ps920Fe9SldgniZaUV70LCEmJjYD8irmOKaCPeF3U376bf16sVx47Q5DKa2LYPR
82pJGWAhocthyytf8wS/Yut6/SBP01A3Vy5J3Uuwvb+qTAAF/kvBuamicuwp5HJp
+yyobl1boNP7DJIyIXYQhW6L+tEbTlDmhfHZHk84x5vV97uYP6WctUmCmD21GqhO
SFdPNi52hC3lbzIwkwnDqxw50rNvkYwHr7OvsK8+oW4uUdjOvuyGBk15+/u9Efqn
T/SF5Q1id7ENPQiSrobVc870EFfLJPVeice0DQ6BxK0sXbD4O2X7D/4evfWqZIRe
beMmPx0NmlR3VMmmaG2+N0knZf6wKd9I+dV7eUzDAI2n3hLEhwGaH3lEaXO+LXq3
uIh27vTYRTDZ6210KknxoKHfdxIPSLAX9Ux00lHURFMt+coqaERpdbIg8IqSui7B
38q4/ufwp9RS9+uMshokKre0m0IEsCTodMsntx/zRlBqArcemrb8ExTKOqISKOXk
9o71gS6ZQ5a+CGsshX/SauSmiW85VEkVocwPzaxT/mpnmjlj3AlZdYtL/kEDNHsu
U1Kpp4pVY0zMw/oJFMp13vqn46oFTzNrI0zGZ8sVEjyNuTp8whKpO8eutJgp6jyS
saDybqSdNDD4NbUNe8EUmG84uFULHkw5w944rc6dkttkYU9yHuRItrI+kOcW6/rK
an0MncUx6QIrgyC0Ym/FdOeXaRQeTL/aA89cX/a3d3X/+oD58hKMM5fsz0jwTAIf
9gOvqGOc7D9qkfY02ZRcWm5sPE1r4grElGOzjHeFbqXlOEpxPNcWuYMHeVbMnmGV
qRPzlB3+Gry9Ii6hP+8nurpq/LhF8YDHWvtwTdAooCnzSL6NI3IS4uzbvbuMzSY1
EVKYojvSN5e2RX3qN70xKwh/8TVGmh3mcSL02tR7NmDkV3BevPKUrXjmvTjCQ8yQ
CxfWVyGXELbg+GU2AbRVzccp7sbkO0y6imWCUlhS2kHA7xJ6+pl2isAdBSoyLetm
g1tnBAg/EzyZ7PwlFiU9cXTBAjf8yOzrhj92D6JBdsL2NnNZT3+2RXdQjHH5D/W4
CDMZCcqDCYPtV6a4dMoafOTy3YbBpl+n0dLm/rFJxknnV/HHYt3WnpqQCXkEziRG
TEs0kinRNGfHtz0dHAJrlnf3sSe2csPc1FDVhpxzYOlG6q52skxU/czD8jhsHkMy
oSc+qKeqG8gYLAYqVwti0G6urYr4FFJgloXyi1066ZjNI5w+Wu4lsF8M43zKMMdt
kT8VCdIaYSTUGpJ9mUxKxTVcvu/+AYoyEHzHvGso98AHJp2lgASqfwB0PEP2Sizm
hfG125kts3Yr5Ys7BORlFPqbJj35e1sdXvctifNEGHN0vXH4sPY2bf2UTY44zgOl
T2EQ0YbSLHyiukcV8zpmownMksCpNtgiJtR5B9uuPNUcZr8JVAypkcCa4nasHrUq
n0k7gdlG612lZWt3XImwmoZr5MI3fqR53rcCFl1J5MTURdzhoNIQl60JtK9T+1I9
csu6gWMAbWCdurUjDy2tEfnOfY/VT1f+fEtt1Note8tes7KKzqC2Z2fzHjQc1IV+
39AdoTNHMySEL7bMAIVepzEJAv4QA83isuSwxv/Rh/iu1XjyVe5mJXf7FzS4aVE1
CWaYvp8S+gEnkCat8WAvVnb1pytiFLFh2NyvVJGBg3XbvypzpuCLPFZzOQX1Dnvk
+VmSedSMi5UDrmbwwoNHm4DhefQugSQLCQxABtv5idOwFP+Meo3uW/G5KBUtQSAm
GhHlqCY2VVUF68+0LZQ5Ayu3CQt9iDjBc66iTkdriCxsgJWCuuSmz0l2cyS9DkHW
RqgSETbHmE87uQSV4KTC7L+xEdaKNsLMTBSa9XRamRvgv5GNZJGLvXXkST05msmI
oU+QP2FibsbClfsqbXFw0B2wzmnzgnC+uZJpuqe7f371Sl7Bpe8+37YaIypXEw12
JNu9orBHidc6nTMUbgTbeHkuR3JGokm13zANZq8mQN2upnR733zd93y9fiw/Ernl
/ilOeNGzl7YuDxtoMzMuhxj92NJ+MRTi/Bdy/U/FPmKX4kYzB7pw3Z+9Y3Bk90y0
9v2Kh0DsxjU9mAKfeLzDgbam+1wYUMT/QmUZpRbjPsDpCw1cSdz0vF7f5AxBjcsi
qBeN1FZ9xmFLENXGGPy2PE9l3GVaovuw83CnYvz3zdjNUn2hVNOlg4KvNEUaHjEn
HO+Qwc/3oC8e8fL0ML9kKGfbNZiUCCL2q86YZOjSENjFo6QOueyWk0mjL0FCTB24
aX2sk30z+oCFVoof4HgubMYsKzmKEKMFJkRUjDDJC7TxpwBsaUB7uf2N+jZUwkC7
yiVrxUUCPragjccsPSIK+VzLkEFA2Sem7U49Zl/LrIJGcEtWEKma0IAPG2307bZH
39C1lgJLHNE0zV8kwWYghyF0vSN8it8/rH23dtcRYflWIxYrLHPUBJQtOI30z5e/
SG/u3cRdEeU8w24rRQuQ7wVEOodcVeZO76TMRk4krLTLSL5zP2hxyU2i2tssucxU
/OzbTaugn+ZUHDDMItt8vzRKO2Dk8OGlJECryDuGTsUmv/y5lt896kleD+GGjXOI
Qsz1WYvuY5o/V6g5s02x8eNdZ1Ha9V3EG7+SFSgGihwZmcemRCtnO4a6M2AYldUM
aUgq7Zg6fuCqBxGBSMeYyo3nfLarKbWu8elB/m8G0flWSBDFuPBEYZ7eAFGU2Sd3
OpY0E6vbBsSkQXxbgVOUiwlb7lqfGWLjed5UlZY+B061x2DCC+uvFWlX4j6P529N
mIEpvoSv4cn1bbPFWnZRrf70UpC/8ucbR/kGrycUYWOe53TuDWCMKN+ZdtavzAGP
tseISnG/PTUiRKv0rlzBwb/xWkQQhU/yE94ESrYEQRlTSF2Z77BfSwmN9Uq/HbKC
1ZZHjm1HOGibWi2WQg92okHOzI/9u2hS5AzZJCn6gX0/YVoAGsluC+xbbxz1oKUe
vm0eY0favLGRqtvORz61PPnw3NXm6WoAYDrL6bd2ku0rLCVpjSx6+kBfWeDGS4EE
rLHzHnoPh7L3g8qrL93mUFXFvsHDs2PX3STC4yloYMq6n+Ka6djSHmFFjmoLNGWy
JensJ9mg6DnGhDmfHp3T/3oLMGfJrhsKuDnXrb5HekGvv3QeEUDUdGCHDZQ3hSJY
HecRYN6t0xN9ikAmh+a7e+1Ef7aaM5k+Rlp7dmwvIFZlrcDxdhAm4PpEJxeMgUZg
YQnwWhubdB+89okaSgzP8CSx+kF4tBSNwxLYvyUu0isLvqljk6hPDa49G5YAnu3/
9bt/T8ArffzW//VRHg4taqTA0OrbBvAVlz4G1qmqiUWo/hR1wMHfJZho9UNGT8AJ
uHlvz1z2RluaS5dDxcKpX0oWDccTRzeQ1DlFhwxYLtDqDdsTrtiMYnqhn8vWBZU7
GJVBCqRqXYJ3F7xD624QIdXAipRYKS29Hd1/5kMsoNeunBbYoLxAN0aG0mQUmLAT
r7NJOg++iEmIXNOiMQS3qb2aT1JwtRPALUnbB4AFOlhDgJorke/C0z2wCwbRT4dL
GWX0r6iUhsX7xi7tzUgMVNI/39UsdjzWAkVnRS1R9dL+Sca58gE+SydSmCMGO4Kf
I4hixTGE/iAFdsa+WgQZFjzynGXItJWnxwHKW5ms0UO3fxU3Txv9zGnrtoHggs7P
lSssHdBPibsJCq6XzTWevgjFHGbasX7i/sNIN9SmFEF4nD4x+/ULqVLESe/D+5BN
8YL72TajLa6vHqG9kdouUMl4MlvE6Bm6R2LTrH/DbyvV0JX9VB5A6cvj5ovLoJsu
x9dupgbJQ8XeY/SjTqNOsxUQDdJdaIR/W8zh+NGU4lF4QGAK8POTYVg1Dz3UzILn
Q1qqBtcrN5MjW0ww++R0+BSz0wHY3gdGkpNIHY9rrS8zfd8xAZmCqngjfNej5IMP
82C2/6BJA+fsSN1hPK7nVJQPCxA22tpwAoeuqsjMhHIGtXV+0CV2WtS5FFDKwVm2
zbUayNrH7fOc5VgAViAyppJky8dy8NnVqIrAgjarrix9GOJvRWxOEABkve7DjGQq
UO5pqBYTXVDUlBpiJFaCyHfgZfxdQbgStWwOLap8c7LS1hH7u4VoL0c+grMR8aK6
wyjZ1EeJWCS+5of/TNNdrGmxPc4K8PF6pPX+Gb/nvhsyppT1KTyanPEOvVPW1Z8X
CDn8PeE5qb5r4jQmWxZZ2fFgm76SmpQN4FqgzMUxWCH9vJgmFdHwUC0XAefJGuQn
c8bbgHZQq/Q/iahmUX1dGjLzT1luR+m9ILrPaJF6zfZCjwJemkf/b+GbC2W7yojY
UhbUVmEEZ+WzA7hBdqsw7fx1qHt7dblr0SxPPyISULIbK9QDQCfSRAUnOLfebDPG
Bw6UlSt4WJNuxzwDBXdbryzxZYkh/6XWGBs/2NDqxo67BvA0F3SIjIkIk6yscEcu
yxN4NjiJ0/pClEbmrWbUZMYSB8IIg1sS1av/fPqRGkb9KXZezozIyTpO9URWBzhf
N9dH5s0SgPPcHbuUvEx2Srp02sVJqwPFdCtByfa0bf0xkL0RQ2LacX9+U9tiKhnJ
XR6AUKG4frFTD4B0877CC3Or4wRWzJdJEEz7D23FEvm8Z1PqaU64cVFh7LwUSbAY
SmpNs2onHlWuJRsmy0j5m0kBClhihfIl/8eTGcK1p9lB+fz1lOX65vmqnG3kqrzM
HIACnYloP/kNvtdWQkXgfGNskBfOWH+sP8R681n+TU7sbU6qorjWYeatRfWJt8m0
Uifuwyts5qlEPZq3jTT4WT2vSI6RU2VwcAsNJAJXMz/DwxIuShxbYPb9prNgGpEE
B1LUV8gR5jkankaV4vmFXJpDqvN2d7pL3VL9QQ/wDR+/e9OQ69hgl6aG+Elo96j3
BFzjcWlnuqKU3EydhukZgfKK+25fxH0/+Xnuox3xs49IdMnKlx8XukaCa9wg3tBI
nW1XhVMirItlBQnyW/gSuR3vM0zRxmfAVrnlo86+p1XowOofKcVborJlA7yOJZyw
pdIKEEce8L1lgMou25qvBAzxFEbsETZu46GpIPJN8Uc1XG+86CMJuBnGcFO2SzJj
hLzZAF/5BthiXSlSpsaG5di8cCbs06jx0lg2ck1VcZtHdryrZrc/W/LH3ojY6vwe
6zgR8imdpZcORKasL+usIiisVoWVPb0+XIkyhGxMCiZURWOoZt/GA2tVroQFfpyz
SyYL5f6660hDeTJVZrXVYGRGivgYwKXLdLP3OH/Vhpmow+yLnbrLE1xpoYJqrb2z
UtSs0HKan9ljTXVsAIW04RHTCMJwy917W2gQosghqT6U52jdbyWjg+WBogehJKlo
P1AYk/IhVbyanDhxNKkPKCkPnJSpOQl0hgY/I6n0hVQdzm/+m9tvTCEIyZaiD49Y
4eBv2/AtbU0HgtiXvyZ6+gcpNQ9Sy0GOhQ5KebYqmfm2mJvaWiMtpElw3TGLACln
BdbLPWHAXAW8a6c5AFp32k45q5lyB0P3lPvTCMOk5alFeWq29K1gz19ahDQiELAy
uwiKe4XAcE0D48AvKYuo2pjfIRy+yEq9fD9+CC3C0wm0sE57jwpDDkuvBKf1QZIr
64JUSkgCDNzR81hF6GJdZ81WtOlGQgduZNd4aIebzGRKO88ShfuQXjM2aSAb7JSa
k7ebAviieq/X2fOUhtdebNmL7izypXDFJA3Xq8msvZ5dmQ54QGqoYgXQVEYf9SjF
fFvdbO3HjjdsGMAvlnpV4Xd4Ao4+FtfR+8o+1L+6ZAIotRt/kYADqQOPQ5lY2GQo
/aAefEQVCBAcOERWbmEHctZMY2fhcDntKtnxbzhEDFiE7PVk3s76/9AmWCFby2V2
u6g+bMlekDn3jiFT0GwDRd+cklDEmFC/pgi36ff3H0/ucIh3HK8isRZV3sGLAksu
Px0reQYqNXLwpntYFtkIAbX0fPjrcOCSEPf4T/qPHf8dufd620ush12/qHVkErnh
pnI5ufDT0Cc2KVNLDbSwdCbMfG9KDNrFjzaHjYjJf1/lFI9R5yjloprt46EohLcc
`protect END_PROTECTED