-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fiRqZP8wInXZYhGs9vkSQZS9LHhA4myx9DWcmh6uIsBN93RO4cxWox4MP4O8L0bn
LFYNyILZPq8rbwAK0n563YrSDdKtTMir6G9CDLQiq+hs00Ezc3DX9lrYvC3kbDrI
OcJoeYnxPQCGY6Eoc2a4J0kynzqZwcdhlo3dhioft0Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24365)

`protect DATA_BLOCK
Hv6mLmeVxGm11zCoIKJbU2ndjSH4QchEi3qy+/ELHr92FJema4VwB7emOphtDj8J
7SGN5YIUvXgOGWIwxxad8DtAJ9CCNcjrlLZ+hpcoR8UbPJZV1ewallh36y7K/3uc
HPuuRg9Li7mjMe1GqOMGoF2SEBQrm4cFqlu9SePesI4OncW38uKimiTUpkF9VvZL
8qeSIaPNNK5CH6qjNzoRPdBjabmsp+ERHi+HUJV0uKtLokT3JocMIxYAeWbs2P/+
ie5JDOpS3F0kh8ZLiESy4vMDx4BCayblFWxOMKMau0avBP7BEsVJhUnWVnktwZCH
FXB/FX0l18lMgRys96a3t1KB2nHNlzKu+qXjNoho3d+u/Ni8OoTEP8T7YYkBXHQR
KesHaaTy8SXSOtl39G9CxosIvFVGu2nLmfo26ngCNzDHEwC7MEFDb1HFpPadIYCY
IVIZDkBAgEwxV1+DSGUHGwSDCgm2VlGwBPKKqAZlHrzsHUBXXcVg1lR6c8sUocsC
7R72C3yC6/iFmQtSeJ1kfXQkZ/f5IvEjz4Dop/KFqq4sLRz6z5fj9aS4IwhoDu3m
F/Pyf2IdlQGKoWF1PBRMHW1wJki1d9huKIjUUFXLgOKVAo2JYpeKIvAuf5jrHkF7
UV7yAj8x1QoTs9x5m9tLj3TsONG7LE+DG3udy5FOZfUERuQC+FglQ9/0/xwivS+T
IKVoUk+8l2zrK1Z4I/SJnmljeNBqSxfGru8LLyP8ej0u7uWCd9DqMb+lAl8/ajzj
bSIIV+EYLE8eckIo3f5wz4kDQkDidpTGy1g78n8cweu4CRuQKPHbxVH9IBUXd2hb
HCJjMx0fAjYv/iRgj44Y3qCnIkkvD7wwCkaY4oYuIx+gCtH+JY5VZPL9pafmnk6Q
9/uYrIKB9mPCpep7jxiRHMafHUvrxlO1L1pgpOU+6T70EviKGTman72Ee3HE7jFQ
/f6Q1WPlGdGIreEjbb2XA7lyTlx1y0hxNYa1TZh802QG8jVzYKWlIB1jWI8EOeUu
t+kB9Y5JxtinRE6KhF37xIP6O5/EoSwSIYhFNOhWkky7o3RJCHvVt1BGZL4wMs7I
FzmPwsUcJoF3cAS3hr4Mlaf7kkRz28UpibV8RwTeZtFXq1S7POlOV5/ZWc4hufX/
kE7W3t+BvzKgK4zsnBxaadhOT+ILoIw03VRJfKiJcY9JVzMFyHLvIcZs3Uiaj9Pe
rAnYUnGe5iAJpnnZ38viVgoaZUccc4+ue1M3SItK2T2nBxg0qzRDRjTua13K0xPY
BHU2epkmUAAbrNgDBSELfgd8qK/FF6npv6zaotatWr4wakNSJp0X9+YULgMvl8aA
hczgaw7NxagaPrvvKTdhA8lswB0WGvb1ATypO7gYd8P6hUrnqB3tOHYJBgBhWlRY
pAt7mxoY8VYoGKDYhLUnOMZNdz9vq6OutzjeQKrP7YGkFxugK5tXoWCJB739Fa3x
kdHaIif9/ZcPeE6A6lwON6Du2iy51rBEmzBZoP1zWswVBDE6DFyqPo6AR1octQ7y
Q+/BjBgpu2qY10Tsy7KVCGkIDzt7ISahovB/IG8S3t8RajntAGQIgScS6Xs76W2/
STJUG7nnEfb5Zlr12sj+nuCifpJDTL8T7LdU3D3W6dXcc/td37Yl33q94O4DLzWK
NjzsZmmkUYZU0eVKL2Wk87Q9beZsYhYb3EAS2jMKK86K29oeAFPToeQusfYxtdDI
p+w3PNeRDVxdXN65VXneRtAzvbVZv0l3iANwV2n4mQ3rkeq/xHByUswwo02s+eLJ
HKflB04TEbCDWVj8AgcVd7qdSllP628ZRxANJNW0xBwJX/adtXlXs3bfrTNul/Ax
1wZu86eYGH3q4m4ntO4z1x0DV1sMZtY15o1UeoA3z4fWo4ASb6feODUwFC/ziONe
PSLq4T6FT8Th+5IVKUp0E9l7DFmrdcT3AgUzmu67E2LX4ZCIcuXWunoMru79XlWc
LwVK4pnUApHSfif0PiM9OvAb+J76LA0KdUh+BiQ/zSNft2PvltRykawZc+F8ytXy
BkEX8WxGeszTOUUuU1/YgCp/Xd7rY0NXBtiMrldxEktcqImTe6sVcmZrim8QEwcU
hutYQq5KcpAHrWZyilcHlZZ2zP7sJU8hLfwgJsT5+e1E/QeYKq0P64SbqoQQ/B/K
cKcwQcPQoxdkyf4djD/lhPXHIaezR4xQV/VqNDY56qlnAA6fa/nOtcMq7ebZnqkw
XoUz9YLpak6D2hKi4xA4H50QQq1c/6KVa45//seFKwgZVoafdR8/JmgJ6WHyCcHr
hXiOt0VYQbldgxvdJ4XMF51fbzFrrzNJ9bnqbFoqujRPJDqd8uP1EgZqFsbkqYR4
QUEoCJNvmTm7qdXKc3fB4NfIVqOEXBOyNfZh/qEFEkX3Iul49ZbRtdSPhJzgZzOg
qMYE99li266ppfDiwzPlJS50ZAaMTe63pGCyRc/ayEygSx3w9rsqAoisoECji+dn
kQMxMsP1BpwedasrOzcNPE9KDyv5E0HbNrX0+hjkgKZK+jSlNuk+jml+1aOC+H1w
N62NZIXM21tRC8sQQRH6LaD5NFR80dhfE3i6eEdISiCGqNSWqzqLa702urzKXz+I
ivvVy/GS+Vn6Y5HSzmPvxh9F/IpBNXoCWvtijwgRimCM4egHH1JdnxfLwx5pDTNg
OlhvcjmQzJKdn+QatN5HkSf7ujennn6nXbSjSKK5kJ/1Iz8Ow/NYGORGWfKsG8ie
UJkMRdcwtEixS+502zVbNECrFiMqWBHx6l+qm4mx/mdcsg2AIM/VGzgmoft1aX6Z
roGiFOPPgw9SgPUsHOQTCEesuv6EvRAD+wyom0Imark9UoBu25SM9VOPbEX3MxoG
E5atVFqhUlPbuNpRb6pq8lyO3LkDNuqjx2L19v0GFHcE0vYrO5z2SEyggG44oaDc
TspGgyOgdNz6KzXF2V4CbQhG65FTYySrs/GsFiqm/TcH0ozoNQ3MA6zkhiKSKjeg
CsAL71FzXZ+jK2969XXn4bf0Esk+InXq9cEIw3m2OS5dT9fiVMRny3W1yWUme8fg
MlL9gqLw3pMtwmFkwx8Vhi0n3iJo57NwsNURqr5n2npnhT+41NB74Wreo6o11N4f
dXGONnrWS85FEl0Pz+E1urv7kXEuzyZM73MJXrV+nDViJe5EaR6SEcIKZhtBr7CE
dZoP/271U7pbQhKBaTbxW90S6UCp1kLRbBG2zwPQctINgHXMWsIK0Yk0CCxfVh86
s4YFjK6Xv84Y+Q24DzGpsY0eA9RAbhFldxhZIU38UEUEqqCACRcIIx5GhyRXX1ow
s8vDHMrkoxmZV+uRATj5Fi1wVFGCNPjhdFcYH3paetgiEa0KJkmTtwsRpRHP0h9+
AiUON61cOGWFLwx8UixfASKbUDB4gEw/6PR1FN4MnIwf8ydcAbRzAbcdnI+ep52I
LahkQDVgjmWExUIne0gL9NOxgGe/9+CCoQCoTZLe38jfDcsJHZe72D21lIuZRGwW
qXqdz3d/q3FG3ZiYVayIsML822MZ9stW04U+EiHy9bsI6o17r3MUhKqqcwuiH1Fl
+nVIZzRfZhl5VcP/0QRbTvIwqYC1i46qT7mZUn/TbxifDgaEjHErVrn7HdlSPW51
llp/uf/Klm7fxd3zKmUWcy3bhox4cDxJaIc3sLEtRrOgLwduvkrPBKgOfdiZuRQC
qWuhIREe/BX5drhxwsKEYj4aU7XvAZMYkfkswYUxptdZUV7+aNywgeMoOCKri0p9
stqOd1KlWjmIvMOrhUlvR5YI7fE7vGrwZ3ugNYS5x7eg5ocQnJb/shQ2cqGKUtxR
wVudC0YpLnlx3DtJP1KUWcOa0Qp6nWEhumoyk/aAqadgtgLG09pVvg200Kk7YFZ2
Xdz3g7gCeDIwZuwq9jRQhnsKPu9KTwvWBpsuL81ulHK+NyhuE80T8qAwAa+grUS5
nt22CPz1bmMq1D+cYWFlcUUCapxLRv/Ea2lOI2wko7Q0LmPELDWv86R5YOhhZtuH
IHlUVvAQW34oghQfCh9oBDKp6ie3VHJfaDS5xPuAltQr0MSj7zSC/LVZM1iEaWYu
lj6nvkX6KUCl6y6vsCGg2NRlvk+E73jkJ+ZPMiOxxqmg/E4A5+BzO8eWULHd5Q+3
+VXsUQ10wEV0+S0CP3fKL8oiGCtDUM+A2gWw9WVi7RSJwv71J3IM0scXgza0cYAr
kfyMTwqbIgAKe6TUfWrj+TjNHdB1LZQvhc33KsY51+fgiDk/H/02ZSRn7GAY2Yra
D4ZDvT2thCvwRRTInqjUcUp6+KYdn12sfax5dyohXk7AqFi3AiI84k2K1O/zltPz
sV2/8/x6RabQ5zc6RHwgvcFZDwc41ziXqIqKj+90uzQv78l5q/FAEsSjCZt5Mk1E
7dabSd/NpB+qyMedbp3SFHdCz2aK/NrQyitnm0+I8STIAGymH9hFX7j2ndTwRq+a
XQh0Wxja6hq/NlFvsceR4cxZk3TUrnFBSkU27M5U5AC9J72h0/FuYW6ZBOtJlkH+
S6tavvW9k+NuJjPSEUC5sy889vh/jHRmVdtLYU8r52DzzJzSTg8+bp2WvKeWwKPB
h5dZ7rF4LFBVSj8ZLx5TIQqg4E1Nk95r4sZKhJMqrqu8m/LX7FNqBA/uelCBYp8r
3gQlub3uId2mYhXivJurtcuYy9OLZGGnBl4Qt0AozKPMBskOH9pcBB3r2qm+MjIF
CNvz4/uRVrvZlwX6KOOvTL6JXMBrOsGon7xXYHGydYhK9iFE7J5ubjOQ7Ip7leoc
y8Hi7Kpq4wwJCaoMYogYUJEyiR/v9T4CzBKxVcuzlvFWm3OdhWVjbtIYhURYGeKy
wpcxmREU14rytNEL0YLxsMNfraAnVHPkKIY4bp1AgBZI37ujy9btPZlT5mknjMQv
guPJtaNUPYJotYchqpXcCoO3IR9p1KfFzNuJkLh0Tnr1yh/GQFDNOT7Ff/RmnUG2
xrvlo3tP+dTlG8vxD0mGpu/8qs9gP7NuFUUsOaAciaHhVpKkbFauaO6Lv7NpZlZC
LJUR8xZHTV0/AXsCCgPvTSKWpm1WFMHympTdVPs7zV53sTOznw/nZoFaCliCtLeC
Otkk6ivBjoXPyxcnqKURgf/5MdPHX2r99Ek00tJ1zsv6bQjZC5yAoVqxr2nq4GMv
gKNh6uICxTVyQ5BigH58zc97PS5NX1nr1sMIOewrcIKYZClN4fvTweIpKKjp5+Lq
1ukS4JZExn6mZfiI8eX8CXwVKRwDhZaU3L+I3nYFilDXQcR401Z7KpU5kbEy4DMH
YatjP/G7WG5jPt+pzFLm/xbxKCMCOEzUWTJkupG2It7l9WYuo4g8j4IW2nZY54Ry
DzpufhnJtBpmGq3lXbbMIHl5FsfsXNiKgQQG5m8l7gVYhz3JG/E5g+V8qIeFoACK
92rt6BXgoX0sL9lG9isbzHF5gJohBryytopXl/H+EQzCrZmQViUxTTNytChE6OmP
CefLwV7axQuC1yTXvvkHMq8z84d1Sm8Umr2R7qXcYlw/rwQX08EjAQK+MuHBqm9s
O8wK3qZ06DMwuBMYBJyseENQy5say0SJIlpJ3bGh+7xZChWzoKBO92q4oAKJUC6C
7fCmBS+VY3mODshRtEpWmQaO1UihiuSKtAGEwcrvVvVZG7q5TV7meqPTGkflFqxb
NhT5AdgOq55sE0cbAs5fpE6U6ZpiwXZKlZ0snKCHB2EeNDnX1WvqPTWzxhH4xW3V
gbIp4wgGpys/9LwgaG48otp/7cTaqsrYI6E8hmE7mGSXuiqDW04shGgDnuFU+T9Y
Ptis0SNeEQyQk+KQCG55s727alablqTuPL2+nWrh0O1ijqEgyuI0die/UQPpLLj/
QSaqVix32uMQZsDmk6UXGLIXj5BjjzkY5JdMD8jfhoZEZ0zHUWF4ER250Vg48/UH
icClza1Aw7QJ9s7ww8AG+L26Ikktu3pc3a4ox6urZtO071N1EOIzAfZTMcjCvB9K
AYxmlyNgdhMb4r1zjD7DyF+kQ4YqM4GSY5FGdzA5m2HpuumtgK0VJ0PcCtDIRnrW
K2X3dh+en+sQNgfmadscPD9fP36gNbOnn1akzpV7AmUVXQFK81ABEEzvwZR35iA/
Zo++Xnx4F9CDUiefkKC9m7OaWb9ZjO7LNIWm35sq65uNpHhw5cFhsK95nw1zbww4
yHovPqFTJz1+tXs+fIgw4LcgTFr9B4E45CIEA/BK07bymel1EK1VWdf+JiiX2oiK
/gccY8cxMiw1MpreQJkKeKefqwuct5VXXlw80X66eQzjK0Dx+5Vw6vMVTWYkSl6/
KFjBj9jSQDa81KmqOQtIbcF4we5gSt0WQpwRWqdplAFE2YLLnWQYv6TkhUPKeigR
vgGd6B2qg83CaxsMfkaa+U8MB7BbUt5QU3OK4vyiwojitTYD7YNSk1tSK2UX0UIv
hDRntfsVWOkOOrl6KCmxw7nwye0A35bOCxfuhxhFHlBRjf3WnQ2QDZ57IGVhSKY0
07JFZiGDNQ97xYp1ILm0kSYyyH3l1NMuuun+hCm3zQkl8A0rrQ/iSG9LHDh4eili
jMvk8jlmz9p1cmjyQjmvzL8mLj1epEnHY6UrjVfgwMXZ1NBHvPzvpr9vLJrsu69P
ahV4QHTB+gUTLiNfc10aZjTu1FmcOHcVMuNNlNgnfpgd6AMLmt98IuN6i7ctzH+A
5r6Fgc5ZEsXm1d3O5wLmI7u/YojOjz1iTyclcm3aSj0WoQ7lrJppMdTcRzZJLxxa
cxC30AwC14B4jGYDxc37AGZP0Hj4RQb0udhVbqd4GB9eF29QYwOuNV7UCBmcnVbs
A2fR3EdRZUi3uCx/vHwi/eIIMkZv/12pTVJFGpmDTrzeezbvb4jqrQqQHIP5RLsT
uIQCPet6sAQ2duXQBuv6/4oStpDYIVSM8QJiCiL4jpyyL54oS5GEX4QZDbnoWqho
TMrCnf2ryF9NssKyeuAKVqt5nwU5QiyyUvwy0MyziiIYdjSSdBR851Cfqd4dsw9X
Umhfcqe5gkDhSRVV8M4FslF2gabwvkqzCv9ZMQ46UnlZYPuj5gZM0bVrEvbqE+32
LzWpM/EgPR25bThhi9tFWLb1DV/OkShFW0Sjlnu3uix4u27NHA4MM3pMJ8lA7Dg1
EwDj+nX5nppzCbSOML0ih3sWVRpJN4vQKtLdLJc3zLO+UnjdBQyjQUaOASYxyZ3n
mFJtDC9ryJ3wOkNZmPK9+71NCS2SnWARho6jJbgI1xsGNrh+9ZLsoKYO18rP208U
UB0N9m6/V+RM7klZImQ+72QLqRCBXPrc2FRM5ZIWuhw4fpMg3/cElR38SFndLf6R
0AvYTDU7eVRtWvYeTLST0uirqgN6GmUgQfDWKQl85390VfA8PEtYecN5J9QBIfWu
Nmj/PDkhtobVFS7rVgIIxcvBYV8qSRhX1RyYJXr48zjAiUKpkqwYPcFoc/WKebtT
H/mQ8t9kmurDp9R9VdB0DPznKJ/pXk8nbjH0Enqp4+h3Y2sl3BsWZGFSiiyN8kjn
0Rqd/8EQi2hMbRs4o+igdtPFQD5XHiDY+pAZjhPJdFlyBJjc4ikTOnA3cbF7T77p
4Nb+nywOgvfuOeIm3Z9HHrxxGRtIqCUOa5f4npYvsKlJDKPIWH71Ul2ltuEHDoNx
FZDFnw8DF1EmPx8xbVY6QTOKXFZFeHzWWCBNXD1Nx4DMTauGFpMLOxv1c9AAwUrY
LPlAYvSSkp8m4Hucqtpm3AtlCHYsWw5s59hW00r/olzcQE25IbDgx5bit6RT4xAW
ZCPZYb3T3JTFHb6t2TtBIARvbVkOAm3/qEQhm26QwVNxE7xytzkDEB2lw1FQA52q
qywj5yGbFZwoT+pqJE8FEUWPhfJjIdWg6ZTKCRJj0uIb2AyQV9R6o0uHUs6oNrBD
9rmimzmXj7uaMIIWmD0HDz8iVIzImv6or4rYIbH2KZDowR0u5zQ2tfLaW6HX4Gg7
pHK9FmbwURhllKz7vMRJ0q8rVkwg8bMaHEb4l16aOtweBOk4lgZVo5IjUIr5XrmG
L94q4eZDJooE/95tKe6qiNjKXFO0mUmlTM1FbjTNHYSMd89f84bzmL1DgA3/KmST
UCEX/eDpTLL6rC5J66/FSiMKs4p5oylGyywDLN6Qe+6GUbIDXy4J7UMnJ/E+Hn5c
QkjQ9S6SMOLmn74AQVjCmTHP25Ivvq7teyh6AcmnQlbnBg7RxIMLkIjA4+1zYqXT
z6L0SyKdaUwdGAVgLq1QVPMYLcsBAQhMlhMw8Oy+oHX0sezoO5s0wpI6UMI6wVHU
QC8EbXQeYbBncRBxlydvEUyVg49uOrDYe/Y6SaC5J7qa+QsX0SOwBSt3klzzxdqF
yb5wOtmI4EMuIRQnKKB5XnEmQGLN7UFVzF2gHYG70OJqS7JAjVOlruTUSzQAW0nA
jtmtrwIKGfUOBrKL9sPMXTBfSWAyn0390CvoNQhm63mFqYmTkzpb5NjmEfiftydv
heRrRg8UQ561Nh9yAW2dcjAhQyvLgpLbzY0K1uwCPK8wu3WpTHrXpiFYsbFyXujC
Ir7m4Pn7DxAzc/I3IgxsXAQStIUXr2oFQ3+7arkErsz1uD+dcH8cm9jTBhQiVBhY
cCADWSNF6XRjuJczGq6VMEznTNpG3tMH75Jjn+xDgzPFK8RNCsYWI4576h8VAsGf
7+UEXflPARBKavqoIhQWRvH6BrmP2juAW+BW088eCRgyQ+RihG4dswI54I0uVWV8
EGPoJUid28SkFy1nW4zra6ditND8JGKYzdt3T21Q2QLf1V25A7rDy7UOwxhdIQnC
/bctt1BrxID+3+lgfvNcz7YPMxRM6oUgw2EYEaImQONFg4537ep45Vm/yWSouThc
4g6wn9riiS1M2FkLcAKJp0c+Rx9CDYlDwllfD9fs+Lpz6aFdeGV+8vOvpZuqDUxJ
d4WqJpn/Um9S7ktn6qiNLy+IXngdLVL9SpcjOLjkk9sSutmGv3rXWovmK2iXlzrx
UnK3mlXXQnICqiqRQMmW+uDdzYiLNp6fx9e93whqMmXZ3R1ynNyz6yZt/ELmRrzL
t7EdUNqV13Oe5xTDMOApte7PuMlR6SFV1oJn77PVwoYzE/inF+N5VPEl1+u2hyd2
5ZH1e/W/HxZ9b2GOQU/XJjF6CNuH0cB3sMUEdXYt/Ucc5Do/jYjMA8haE29G5ymf
s3+xuUMOX2URxuZFxe4kj6BfKt9DmynKrkdQrKbqsAKLYR6ODRR0DQaZSXsDEqMi
gppj78E8+ZA8VtNxJIibqKqByqekHq/YW4PcVU6EYRl7GAvkdsoebimzrF8o4+1L
3T5k1TYrcro+yTFuiPVB7AS2icsr29XCTEjMMCafpmpYq3MdmBq0fdEJGg4rhBH0
Mdexap2fyZiPkggKx47cnt1q+MuFVe3/zMRAomAQG0t+GTMwCUblQYj9kld2rgq/
1Kq44jU7DJS58olRN/gikF8ZGvsCvPTZcLAHeiBxUbEBrD/L2bdhuRDZfomc5KzF
R/cQKJmH0yuUTZ17mYVJT+YlApqWfQtaeq0w2hfsI6Ti+T/O1EHfJfIK9BOnBLWl
N8cpEL2tHUxXu/7PkPHhtpQT9bcUGdZSVlpagTvIwhSlXth4lD1wFb02yPJnNGVe
8eXMYGUdYzJHkeM1M79OhknXK9aRmIj8OYdP4otkvMYRzFa2xWjPvLfcE3VA7/2N
+vGA7w2I4XbMpj7pFCJ1VQ7CCJl3uoP4CZoTEVUZpD8D8LcpblyGnELNN134kiNJ
Y9ffYmCmOnAoR8f3dj13jGMqXo1/kHid6y1C4jk+km8L3G4/4ukTLa3Do1xf4M5E
lxkYTq2ERBUTzaHvP5DIdWO3r73DQAMwJw4OlijluABmrrEmwLlqBk/UmCTEMSuO
5NRV/c3m+cr5pEcVIQDEPwubTKvd3o0lU6BBOg97hLhxZknTB89T+qM1oiOyMxVP
7+mbqDJXQ9K5jNojw2weAW9b0oDHC+qM8Yeck3otRgpusdJeUiIexbzyUmLpx4HR
l9C0y2EwIwLJKoIAJnNokBHTIwghNk+FhsERmyQT8Wohat7d6Pl0noexo4tjdK8K
+YZUBB5Sv9emA3CmDEcV1tp2eMPHRaEiY8xrZRRwaIvFWJmziFuKmuJwCJHKDuiB
S0LPF7xRRK7lMoV4yjBVSXKKGPMnNng1LAbkxM17EkIqog0iuqGrlLQG8fHLZrX/
TGjXJ7qCuYrrDGMytlRbBb7zrFdp48LfcTJYI2Pgsio4kStIa1SjIeehf00WOUtV
8VNnKZM3w+d9mKMDTOu1fxKcd6Q/T1iQK7uUUsQ7Plr9zHMnuSKj9KjS4r0WUrWT
Uqw9S8j+GrXcnLmUctHdRLWha+MkFSqE1vL+6I1RcXZjKmpAx0ONvQjKCGJHTKM9
TppZH9qUlpDt4aDZDhDhoBtEJc3CcYrm7YIU7sgg/TinZ12tBzPELt7M2cI26Kl1
ThIDxU8r1wYUdZUC6uCMUJ73uAD/hT7knq5fY84qdO67rXUIIYuxLJUflNF8H15L
WgCizlQJ7w4QfaRd8FsGwBRdQRNyptVpM7Z9zAxCCAyY6cq+Wq9hGNQWJa07b3rq
6Kr88s9isB5GIO4VLTJybcjDNaNgaZwIorTcd7qXLdV0GNlQ+qOnwNRuCshKxJfK
TmwghZGLu299BTYpC8nqaG3YzZZf7bOdx4owXxIOzYZd7TVJ62WIvsjX1JPHSV3+
W8XUrEWcDhzLsAYby1T5ncUGvVtUfiv4KLe2UmaEq6pfX3OREqO2QHx80xYg9BiU
4wOkUQYnX24jXAnxVzonFjf3zZ9hG5yMWYMH6WF9Ir4EB8ODulA8zYU9EXU7XHY1
fI6DSiP1UKoKe7brORb//qqWD+Kqg7lR9693oE6Qd1d74TtmKyWEw9gwSjTgHjJ7
NqvjKoBic3dKt5TLYFwZb2wUW7/jJqVTijMTNofJumTSpSHeSV+8Qo8sCa1TEDf1
E4EplwI2B+inYXuTYa5ogdlWSq5Xz6nizCVgim4qV0Quy6E8wFbpySAjX9xrGS3R
zGIK2OqW40WHOr+j/b0d8slZNXXPcyMSjGhDu9tdF73cQ6184mOJG0HZKyOrZ6tr
LAMnqCl+k9EUq2TlVaWvfc+nPwesx2rHi+mffhlUkflGAqnHRY7I8Jtm3rjf9/S+
YsLrZUSU9Ta44CMqm5h6NBA7dyQnCPp8eaw3OYLpfjmsasikGOgMlycSLkSIRQHb
H4QWqv66DF2BughwXaKpN7Zhv1y4ZZMs/LBQ6R1ASGKgwdhoiFLIXplYqVomCIWY
bbdnoMtqi9i4SMB7Bb1PuhkzLPa0x7U8KxfliYGoUjnLAIuJKQy8yKjrBChNKQMC
mLRsBobF1cMFenc3xVh0r9iXxrRLdo1kGQrmegnAWxo2XjTpIHIsMcdde5ooH+33
Nuznps64nK8/3DstX5TFDQaFTmArjlVc0X2PHAeYzJT/jybqhGzQC8S1TT2xf8hd
mUr9NK8j00uoEYQSXACxWhkNpOhkGhAJOPUumuRu5uR4afsEdxAdrb+KL1adxAbA
XdtvN+MoDsZ8LdB2FjUBy62zookdPxbLAGiCcXNNq1PGVs8NzbxAaIC3oeLWobvM
Jl4JNMQno9pP9TNEv5BWgDGCvGN7eXAHohDCH0WVfIfrN9RbUv7H2WlFwHFZx3Et
JG2JlBVaI/HmmAikKnujT7q4r/mlbhBkkY7U550tCHJBcFhiQGBnptfWbaaEKE8u
9UjcSOKErGGTt+lvUI44/QKam6QKi9rd0ZlTUpM45em4uOOlRWY+h9UzA1XlvtUv
Ik5xKIT16ukMdSMplQfCfn1WqJWdk4YDvERrnpvJSmgFa2BccaDWI0NbScxQT+bd
7saF1fil/zJnkZS3ElkphQsB4TOny5aYqfQjcYhRnYQ8kDNZAPm7jXE+Du33LYs6
BealcYJuN/OmHVrYiWPjXmVIIcEtkOT7xNYvCugs0r7BuR9P1yMhibSyCLiKvoa8
IFZqpQaOQKtLTlU64zted2BPYnfK+fjg46Ww+NJdsj5VWBV0uqYuLtpujjs1u5E0
BQag9f6JBYkshzTbGF8MEC/xycFLvOwCfKaKq1SlCOn5fcfd4TzawajeEfcu91En
CikLy5PZ5cBo6/z4lZRT5JT72edb3pZJYItVz5u84OFDp8oPlkPipgcTg99kG2h4
R5U9/VFq8EjiqNLNB5qandeROE79EYsiDOYYTRjjcHA5oL+ESuBHK9//t/nRvYnh
/8xBhwoWOc/gKkFsiap7oF7LOP3m+nf/M9kp8OxFv2NhqiuwbLurtrYKVYf8JBdB
s0bTXKzpQiyyk6DMdQTu3RScO1i5ROJ2tvpTF6STtXTG7Xs/WxERImwLC7sB4pHx
B3ZUryHW/Ewyhmw7QKpdybtnliZRN80Ag9J6v07H63hK2nKKvICsAw/kC8HUtsHL
B3GNjTTgVVeoPF10ZXng3k8HepDGMTjLgdFMGfRTDYwQNAaCNoTryw3OX76ZHoJi
0ROtZtu9TSZnQLbYmKeZ1NehC+BaFj3LQQ1JOQqLrmRn5EVtVgNeB5FgUNxPUWyk
pMtAbShnHiW1d2NiWryReB9rgeaP/TUbu+dL2ajAu/Tw9bPY6uYN4u1sSFNJGdej
FuV+fjnxRKNxUsy3YlVwKMx7AvERII3qLPcn5LXYCTmr33wTvX733HG0XKO72D8e
xtIs8y6OsfeEjoZ2bXdWvmBz9gS77/MujKLXMHJ4acNRhEWxj5sjX18liLWrpMgW
OUwtXwY6eI3Ek1cAWqA+s2XVoU4Wd/Py7LnOCYleoWhGLeQFMMhbrx/lB6Xt+K3D
zWfWi10QsBsAWxJ3H3KcR1WD9Ufw9HM48CO5U7fZjNaYNtsQ3rnAxBmHIgh3JFk0
k+YSgM0bM6HK6Ul3me8DLXqrOxrOA4K7ya4NlPI3E0EkLOE1nOCis0FznVgDrTjT
MwzwQ7LgvQR0TExpvLQ/g3XYSM8fOr9zXxu6rSdTNXOiLz4siHxVvIBU7Pq1TXyu
9gCKXWCP8D+XdXWBEWnqN7kePR6NcQaIurPifiXAe6fG4nMbRDTuajON9AxggPcB
xPRphFeDlmQBZAS7gMQqDQxz1AcmwNixoHKtJM7TR4/JCPbxNW0ixZu3xIpMtsu7
dKluDxKHxdaLLWaqAcx2jr0COdROfRoBilaZjcmVClG+w7OYuWySO4BcKlDHdOGi
ck3K9CNGn1UoZ/5iYb6inYiejCFAyqip/09KaGjSveNSmMeMu/FgiEUAU5h8427Z
1mpKgKF8dhpkJsYHk7F3sud+bG6NCDNQtO7sOwUQRRMMT8EV9nueNxUjah1nYzJC
GFICUsidzZnZ5XyeU0J5XmJozqssrdw7H63AsrWWu1ruD3AEFex3H07zvTwsLcTb
i8H3zbIfsBriIBULJDVtUhUEug3FgGNdgyC8OWYl1qGxSVlXt1wyB+QIYhudPzRp
cZjtYTfLC+M8h/B2BPIRThhNYh7rv7u8YYeDVjXochOeWgyTR7t5z/trgicZKkcl
4jwWfTCitUhTpEAxa8+SCJP86+whHdCtpjSZOVJj9r5rqFaUSB/7AwoeuzBIU4fl
aSQC0K1nVsOY0qBWqZhsiDtR8Ayx4qNO97gLomCs3WoVvdNu9syRjIAZLMm+yMEy
SANwvK6Ai7Wqa+IA6l9h3FsneKkGy4ZZbQxPzpvB6pJvUsA9ii1f8BZyioFjFJGy
ioGDnWpMCxuif16+Cw+TfIKoJa2MBeEXV6P1JetwnyJTfvleQfqnWitMjL4bPZRs
Y2Jhd8hlf1F9g5xzlyIh6LJ/bUE514QrglSsWn4nko1iWrRC2VG/YdcXqK/ptgWm
6QhypQIyoYnlkzrS1gkFJtkDZdo+C/m8kN/Anyi71sSaU2yh6yDlJJz5pKRicKzC
+u6iWbwImxbs5Shuy8xRwxsADfMCii70/UA/aOOuDxrzd91HpbZqJip+JOzYLFF0
idN7qS0kXSO4uYUcD6qHgvtxvoWlLbv5AJamn7awSaOUbKbwCkiMa8AIhfQW7E0D
3DjCbBVnyP5eAxPVpA864lY/wxYRTN76Cnobpdqg3cCixz7MPLr79Fg7T9VzcfcB
zdFgu2uLNiQty/+f88+W2PLgj4s+SkMKVeET4NYllnM9I5enTo7DZBzz9cO961QI
yoAtYPfdkfCBdghnjyM8pWoOVlTl9XB6HXr70aAtBWxrhagMAlhqB529EhNKpo4Y
euwMlpCkyQritTe0R+ZaktYUMqnmKaBx32SicdvTfFKRKlr2TjPp/wk7Uw9Fg84G
s9Z8Hg/kAZolB/XJm0fdvlul79B8R4dPOVJpfQxjCUuhv4hjpUlsqM79H2ZskPpr
jXqIEnCVHDdNMjnFUGu4hL66KYkiHJXghLpefYDJgVVrTPHOarXG299uTwOH8OKq
yV17QMxckMKTo+8Crne2aBXwsyCRZgaxqyKAYi7gxLBkbKOj6cij3Tsg+XxGoKZt
px0rUVOvJvYlGUJ9CMohUH0q7Vjp0Hw3+Erzj0hf6xVNAZZ3rrnRkfZ+5clp26eP
z1chkAHajZAAso5y879q+EakEFEfhtD2iBid46igqxj5D9Oe2RMsP7CQfces7RNy
YrM1r5KNXGv5ONUkW0fqBEoLw+sYgETuARHbGkyIRbSV880PEQtMO96WA5vLs2vl
MAknEaH1rmZEqz4H0zXcuaSIgbfuAHiX5q2QAQwUt0zD3WOBCl84IYiAMNpDUwE8
1B4lPy8pUb7uJmWY2BhcavHQVmIEtE8eINq6TveqtWznIwp/nqTa/I7SdTeMlFxz
XCdE7W5jUCyAjAfzj0Htq3usxCghymdjUKfnnCscfV0Qb5aRFfHxki1n/avRbKpR
6fK3scGU2iuPFn+wjyXjeFQFbzkt+rbWOvBCDOQdMz4wjnIFq5KGS8YKZuNhSBEn
/rzVEpIVew/YYd+yKR6xB7FKR8BtQcxNg7n3d6tANQfdGUuJWWIg01OI63yc7oOa
BwBP5AMR+IhwBPVvVcT95xkmJTBWvqTyZac/K97+LjoX29p6No+5zCE45Ihh+069
pRQZVuveSgs3C3A4ap6/4pWRNLH1qPdiCa3o+CO64sgL9TfVlpb+aCFradAczxpG
O+BqE3VtW84CBpo5YqFihciQu3C8+qM9zFDymy4ZD4ECbGyGybTNf1azyz04ZQUn
vooAHz3S+PVk6uq+xZU7/aOwB3aoGbcX+rT1XoavaRhAX/Ez4Pi/W5fYHNf1SRZw
8dbi+Q1cDy8sWlKfClIaohbFrnmaAdRqhdjHBz1jMvHPORQ+45ga4ZRtp7GVtZxG
YG32nmqHjxdfLc0D70BiF6vdl8lIOkOHGF1hpZW4oJWCNqY7ZFe4kf1uBlNnizkE
5qN4+6EQt9fPuAl//+iHuEdBQqh+ORCMRoAZelnFH0yy90S7S6bcPqJRbXeU460J
25UlhQtqWsY5XIGWxbhc9zPpOUD3gIbWtdxaTISiwvGoq25LpZWhVfF1UVmtEpE3
YWu05mLURnfMyHjz4BgNKU/6RttrCOmg9NJAGO0r751SGa5Pn99WtU5la1y11OjW
hudHgXa2Jh1hR0lUM1RYwV2y/fn4qK/WAiUJAcsvuo6XFbKN+ND9LkpWZ2Q57EFQ
vy5vHg6urbe8HbxWKD35glnjQzb/cITMZb1f9t6rXVoT8qR80sgqRSsQqnPpGxd/
zzv6wD5yTt6xRmN/OGOsOaSOLX2T3pNm1QDVUGQkPJRa4aalpEtNJ+o1sqpTb8Yu
Ks2arU8l8jFg0tKdQaKYKcPjGcGw9EznxtVqk6t2TZUW0p4bEphJ/rJQnPIaXo61
fcJZaqdJ3tvr6PpQGUw3yFGh69pEx8XfzvYo9az0bEbfo1mt52b3YcbKYyEgaazM
q08jrGtdtHyqtT1FGaSd3DW2ObjdsmiwHoDx3bMZs/qu6xjuq0gnGXWC/wRBBOf4
2ptHqrFrMep2ZuhlZ1CJp0/NYrxGMBocRKJpmDsV99FBYDko5V3AyVOlWciqs4KI
ejCy5gQg82YCj2Uv0W6zHBFnD0unHYR99RCoPdtpEjE/wqLFmyEZWSdx98mkclj3
KBZOl9aU6Nfa9FITrWeOpbT+eS+9gQqj7jNcz576iphoC8uSzv4f9jgUWGwaBmGl
oGhbFrT0H+Etc4sM6Lwr8fwWXFhHc0Ei1ZWrcxEqneWsho5nWNHKsgu/V50OPEWI
pxtYJ9TEYwpj26xdC45kKvc4xnlliyO9D+DmNssmydb62nm+/a+Luh45n0bbRhim
JY6MIX63ja4vywcr6hgaOM4YSkTRQ10MR28QMhg9SsCv5P4JSF8sTsyCBQXZZitq
fyUGqR4FpfucfDJvGlmtCsZC/zUtlwo4KbB6hUdRKzxqQSxSjrhQbpzo9FcxhAos
AAWb6eDe3vqCfbGURt1TY0S1QO91xOZmt/l94//ecjTcdSfiiVONx+gZhKBptwaA
zi65ZGDkDhe18x5hLCj2u/6XF6eHNy7aiHX1UGkJn5XXWmdj1KPc8R7jlb8xQJUt
JjtXMrD/BREft0Ci6eNl83xuW1E+GnZF63MkC86Kg9Rfbl3Ns1xoLDJkXSmlKzNs
/pv0JgpWAe7nEhmwBMfaEjNeARJH2KEdp3wgboOsZBKj/fb9mbyB/AeKKRgaArhb
qGjI8CvGy9SENXCCB2Hg1XM6FrKv4HdiPQxXdpxAR6A3HFpnr6c/O14G9lNQ7BWe
FxZSmH16sxLJTyQLjKtF/2GiGRx/AQdn2J8qWhRtNrOFpdA0QPk67sCWGVwv96fA
1Q6DJ4vzm89bVPp1BghQDbpfZUi7L68VoWR+mj/wFiwDYaEQUD8ZRZagkrNXFHnO
M/AkXXfODQTuPBwY3cUeBV49h42HibvwpFXRfYQHLcF3FI8Z0HjDKQVxt1Dmd7DZ
z7q1na+Vka1iiLny2bs3TQhHTfOC1aEBp/u0aVdum35v4bDXYiabiwP1MU77TZpB
nq3NsHNpMGdJP3tjqpnQWEwj+L+AAXVc5VqhHBbNXuqQjJ3X/Md1pvPaWnVayrYk
KClB1tvm9hl5XqOmk4B2CF06XeJSHf8VTmP5vLkKa6CW9gEHWLqwFKjZh23m4tu9
bpIdqz7VfoTp3ku6tOtJ+LRCUmQDoj3FEOXmbqjbLFaiuKQ0+NaTR2uTnGNBPRN1
v20QO1Iv4OVY4/caD5nBhCtrtzsny/viwkOvoYANzFfCG9wb011lJrHrX/b1RCCe
EiYamWJ6pdW1bu9jp/0Gtas0L34kK13CtBf0EcqXyAP8+krhdNH+3ZO95bopKfeT
8ZXsF9ts9+g6ebGHrNOXoNlq58mW7cOGQTr6OTXRQ6AJ/3Ey55Las/dG2R+8l0Cx
rQ8j6KbjP9MVnjWhwP+s+L+tm7LHbFlGcpcnR7nCDIg7F5vcHxW8epGgxijf5sA4
U3Aiq5KH9uSKxKM3OO7y2dd5iHSNAGT4+o4f5HwUq+naRdSy4WvxmAGugVoB95RT
e2v/Qthezvs3BIZofpex/CrGWH8bO6tiBndgckLi0dFeS9K+1ogUAqCSaohgkeZI
xbM5Dz6v3dJDONehpZ5zrc9b4xXFKdqA/S0pHK4WJQDCOP5fYtaAXYmvbO3yZ1oA
4PivMDmL1njN/n96iQjC3BqjbC55/oUsGLiCsQhN9n/GzPZGiX28JnTtoQBDa5Lo
OMgmX9lh75P/J5u3lPZgGDhhcQbT50xkRHkE4diIf+IKFm+nr6C1RHK0W7UuJmu7
UvO8XIhvXL3VFvvXjdpI+9x+VPtbmoZIIYI5LFGZW1K9PDh5+FqnvJ+Nd9mo39r9
vSPMEn8fO+6MbjJhVpuC9XsBcqo1dTbr9YbSLVPUmpTzqc1lX5+xEJ6XcZ99vMsq
r7svJquuBYg7ckk9qgfuBMIDsep5RK/BnQySH0a4sEhncUgqMtpLDne+PC1D6iwT
WwedARatNHsZJLmFyWOkicRLvGI2QXQ61krQKNSL5S4HdMWkLacxjYi9A/0v4G9w
ALsSvyLrscFQmaOtfXmOTwzT71bvGFwqccmL1Gy73LbzFhHV4MtMlSdFwi2Kp3DI
pXXGnJ786TXZzrbCEnJGQbd0yYFRINWXizu2o5J8ZqgY/ddICyrh91JaSl/3CapG
WCT+x3JM+N9OOPpXpwhXtbeYtiRrq3yf4uHd8p22wmscFR0p4UjtSy2vvjJmCFWy
anOvEXi5jmx3SMq4JgBC/4t4iH+OwIUCHjUj3iMTj8G7Id2YCQE7FlZkni+KxyIP
ZwBi0jdu9vPCeZ+RNxL2gikOU6A/tf7UfRg8dKhZUArqVF5tKSWjq2MnohAz7wC7
6Wh7JS30AzLzFMQnVh6MpOUxfMrMoiUvqq4fOXwSWPGi8xjNAIq6/IP6zKBthVeq
dRmTwABzwuPln1rlOqcr/Fjuw1GY+0CrSTU7nPFs87tE+VbFJ/ED7dOh485OsUt3
mWUgsCRoRCI1yyGrIS88TOEWTCQPWeuQ1pcZMc+5CeisNbV3jakrx2VTvZHcXsmh
uWjmi1tt3Uz47fGVKhq1higBNj7jAJ/rnD4dZupX+9/u90YnzXrHSgEUgLVHarG5
mVyzN9UosMQhZRczJNRyhuiHO9aYJk5d39wqdLIFUSNTpMaV1AWt7Fc7BAUEbcom
URKo445EooeMlVl5olnjugpDZqtRROEwR0jTkR2ZkKHAmrAFyKXJ9SLGeyLvxLSS
tUFt1K2+JnLej4ndk+nMPNMT8Un0v/icMElSka46ehMRmroV2fkz7hB1SUopaFbT
AbTUcmq5KEXeGe+Jv+DCoPWYA8suBCbLuHsvUKcn+b8NpEpz3JCpqG0Dyh2nuCbP
NZaBZV8grEoCpsI26PdDUkHBoZJE68TR2ygTCsg8Ti/1vx/+dPzdbGcfVj5zWK0K
RE1Nzq9Wd+Ov0YyJ6aZYX6d3w61k0J5LIVa/33QdHa7LNgE80zJlAEHa78+tjK80
TDp3xV9GWian9itdf7h6AiULWi1TrzHpS4xbSBmnfLO1J6EUbDRtma/A0t0gy2JZ
ETz+LMrdBYG4i1SxWNz41H7N1pm/hP7Ma+doxAlW1zFfuajZOqtskL9sYaYZtgOA
XIdw/ab9FY3+qqZcd6WtU2oc90cNJ+dRMa/VPPkTblSiZMVuwWEdLUHlzJSjHTsy
dgTVlPy37kCN1jJwxxQvJEdWXAOI64Fk7FCoWQsKWy1SnNiDSqW1lKGwAuIdwgPb
HBtG2px78Veh2V3jM8KglWnPfWda0Rm8KyjyKFEVSY4+XqQDJE6zp7Bu/ml1aLRo
aBKK+WcH5cjhBMHdJTS9S8JwDD1JR0PN9WZBARY5bfufr9jJOSa0gn6cYRnrJvSo
O2Khl/ILU9sU4u+Pk+bE9VN4Pi70QpZ9UQIc8dzYr6A73rTrRutKebGzonuPZ0dy
75R2xJevmymsqWClaVIr9jXZ0GmC3cKwXqk1p5WyZHSiuPvCp1J8MjW/Qt25ZzWg
Hu6D+krnvdJFBuASYp92XRb8NlhNgohGgrA1ZKCDYJEkvAi1QYCo5fZ2zA5O+o6K
4RGMRS+tvP8mnZaKEbpD35TTYe68Ka5fnD/qECviOrScnrtvVGInP5jVUXLUZPgF
JrkP15LCVg/udwpgWOHCMVLHuiarcIONo45lK7X/GyFpZfEHflIDF5DcNUGOkV6K
jPZE73FQ48JSY5SbB+2kHyffqkWvHXtF9sQopkA3e2Z/Ip7CZ8B75vqpPzbBchmX
oFzuDpOYqUfT1UlHjr7YYJM8li7WtHJg5+UZdXVkTXOsVBNcq+5G3p8NWyqOL7OS
NbRhQIOjC98+JWxx7pZOXTEnyAkihKuv65g3Fim/a8FaMsMWmxqd6iSveWVwcKeG
ThUlUMj9zsIOgPrPpt9f3MX8yZ1/0YujgYdrvqPBZ23+OQjflp42M53CUPx8EcXR
lFPSk01KFdrJJbyVdRZUt1B+grmncg7oXKP2P+6w7CaUZD/ZvU3kqCY8DN9SFL8D
QYAdxVHgJ6hkoRuBFy+BAegHwJEzLywKWR4Qf/gRsjefxVFe4eQHkbnlriJXwZ5d
dkQ4Ihh96FvJksmrE2WHt3Uo/nIipaw4FCwxgEZekZespHp8eVwv/7F9SkgUSfY9
9TILG59UL5/p9noHxGJjqmRUzquJCIvIwycOqlHMIoIAXTicEz3B7CW2Vy+PxqIg
LNaMUbMoMb8kOsbhkid/kmzBqoQ7U2P+okUBInZQH9fRHEN6yv2/EDhkWA0eeqp4
BKbAqzYSvoJ8nf00M3yUrLs0mUXHGi7Spm0H2EGjm5/buQYYcN0ZrgxqSUS1tZ1u
nsJcCE4oXg8Tve+uznS1LfxLS9RoI/5Muf60YEvn2Mwtbmwdnanv2s8/NNkKaamR
6Xr+6zQ8RAq1BaE73EiKozN2LocJY37GEfKsoVsYg4tQwc2F/s31zOKNEKZ1Etae
NM4x067WGfZoB672OJnI5m/EN0N9v8xJA3pBXw+z7rLMinUp7wv7XalQHuVOal7u
3+rbaJNW7z5ruxLI9IyL2BSysgvBNlxWnOUQwnGjdO7i0JDr6rBLKNczguFHbc/v
edIKgVdsroeISN4q0n2ar4XOI0Rks/7vmNTV/KCiYvo2CtOEUZhrLH9pzOVg/LCr
rMp94EAq7AOIRXwiyN4/PisdBP8Sr/0WCMrpV08Waq+jDSA3uCoNkhm+DrLtHMGt
0+t916QT6scnD+zjWauNqIZEMioLBlR61usgiKb8bNX1jTTvoGSiuhHVliz7v1tY
mSat3IjdQXK7ytpY1uCx/V/G3BXWa3i0OomenA+D9/u8hPkYI5SE9xNoLNVvBl1P
9WzI0ZCh+RcrmfnDh4i3pn5GbS8a+hYUp9M1uSN9wfQ6NIUpsdcpDih/RESHgEy/
ABhqRWrseK6Meutf7PAI2VxQYVmXHlGNseLnMHG8pwAx2ss0i3WNApf6yknzB3si
7Lybc+6en665tbNKUqYxqQafrV568nQLqH/BlZnNrXsCJFOIUsUWd0L4o66qNIzn
g07TWa8OMgXZtGljvm2o5BBudLyWncLKbu4BdpX+CxdYeG9H5IKU6LUylBqbpZWe
nThgwhn1yMysEh8b7pbQDDPG8W4IzSRVbcynVa5hS8c7CuumWjHDr5A0mSmLkWlZ
oeoSHIB4zP0vL5aPd7hGaKEldCrHKWil1lVAQCp2LBiYcJ/RIpX7C1CD+xNPqaOA
Bh5UO7Grr8vEsP3Sh0jolIpKN3OMZV4SdoxK95Y0cFrwWCe8ojUc07sr2nD4koG2
R+jVzWEQA6M9U1PvOF8AeTIfOPiR2WAhuO6R7/fROIGigsD5kQtgLCKGhT/2UJgF
HhJVlJXWmJ/s3Pqbqsaaj6GDrHjKeMgv/c9ozKn3uvhA8L/u6oyrfLuC8zJ8n5l+
rOq3WV7u4gsHjaBQkXFP7dIfc84JRSt1jNWipX7PUNdqxO1rvitHwBNKjg0l5Qk1
rNcB0a+gBUfpIg/Al99gmhKibTs1R1ziQTYSCNAwaWV/xLUafIp++zBvJO3wTZ+H
UDaKBF1X5YNxunCylPcaq6NYKCK3YmO+RzlYzqJCDIJaCqDCvRqGp4Ejb/YVvogf
TogAZPXlZWwJXhM2ZSsahYHNvtmO9g3ZhJQaphe9Gq+r31mMua/AUM4V045KcPO6
KIxioPUQhazTT7ThqTXs9MdzaWAoGLy+meEXb3QL7EGAoOOVo6szAspyxrLUYznk
JP5rd3rlPFyyMMvH0vJHHIy/BaqaiSiSSw2QoL9I1mvMY0SJ0sAMox7mQBDv4PO7
joKtL7pIhYNbpdNepEmjZ2XX4lIG5navhi1lELumAYlooWw48Tqk0C4npJSxP1wB
7DyehdIGdkck2dMKh9bUfmZH7AiRM+IHoQGCJRlXPxFJygNAZuZjFNk7/nDc7r8E
eZZfNEaJyrE5/ZUBPxWeT+5Tatuzhk2cK+1aRaW+X++yBWmPzs6k+y3bUubrgU9v
piP0nDyyCyxYnzge2x3zTh2CN+H7pNa7vD0f7bDdpbz+gH5HHEndULhIeZG9UQqW
fsu72RWKFSaYzGPQwBusortXsDJqgOcEk86FVbGFriDP+mAFeUuwQ++CybmMotRx
noL+Szo/ryecPz5F2vWb0MNW2c9jmHoNEYhoNxVBZM1UmbAd/O5hkY5ZSB7HLvUU
685WKa+YHu4moTJ6vqhGtyc0JlqGEp4Qhh/MngUdkwd7N3buBO3fQb3r7f3WB0/I
VwXIFku+ASRwUKE2GbxtYvCPIb+i/Abva46PIOtQcv013IaS4vBgchl6cDc7iXBj
wIs/m/Z5J6yIkTk46PItZOxV1NtigeUa0B0s4fytjTQm/dp3/yKS2rPBXMpFAfu3
3EIIgEcKELbWoDcT5YjezxXgTlVhvMvPPLLX0lIHGYZaJTM+/gmA8q2Zn+uHK2fD
P1t+Q1hxpOrevFZVwyxsrqPvsJihXwr+rGSHyw/242VSY4FivNQ1Zvmg5yZxAR1I
DRoUX6G1G+m9UNGy4Pp+RZI+fqw2uX+da/smijNqcowzsvxCVOJ8leB5YQt+oec8
QdFWo4IhniD+JoSU0A1NBpWnNt6kaLgri0Y+E4ueYgYFsnMLip1hvrD9E1e5h52n
//EyTyFYjSW+u+79snBbLVmXVDy9xH2Agr18xkiNtmEQwJ9lOG+pL+U/SS0We7dV
72M85mcvUc6M86BUKfXkfd72skqrs1pBbAqR1wWhlwE1Zb2ukcNzLNQ0C2Xs8sI3
XFMv6b7oHuYoZBDLJfp1ZBp1U6NHJP/zv3TEK+ghroO1gTPm3pkDiUZpAiGyud80
XS8dPag0sZsgRdnGXuWJYzmJGLvgfpardushbN5VL1Kw0iLiCd/JHIPA0zVovBqJ
3uziaDBBUHsVlfMHAsIgZwcmxWhGCtCq9LjtlCwAs0++TcTm1pbAnqnPMLN7ZRYX
c5+VFIMMMcAcYj+pQaUmssjEkB+INBuuxCQLNTRWj97g7QvnxHD8gAPuSAbTST7d
NL6LiImkGyWuxrlDAOEOaCl19tr6ZH3PwLR/2vl1VxujOfx0ZzUU4HXqaKZ4l8A6
94RihA17EtHs+Xq6Ir917mWPWri/OaYulE4OYuXaaisJwvzBGUrRSDXuJkmPUIEs
vfnKRQ6JRCXA/DQ/JHUE5EAnXC/DGwlMuV78mr5gqX2nZmpmCwE4KIHbcVtRnjuG
LCiyMlFN0NMR5dbwLl0kJyki6LNNq7E8flm2ipFRvhlMDAa6QnhGQuAMYqdWGcv0
dR8fWqkM6Nz4zOhZDKRj9rsloTQwOX4JDoUms2O8mh8JBgqiGG1XghwhK07708Jp
NGF0GDDjocveKjcpAH0C1tNy8Pzn63RmhF3RpOi967oNC0LN3BjSPfHwcilb/nBK
LB5GIu+4lWjj+9dMoNOadG8Nxji+QdabEQ7iTHXyiL8FGNo2vsgXdxbmFSCKf5Yn
IKAB6UM2v+xEzPmoNyg6KHa8bKqlCwV2Ld4Ky5FQg6VVU95WsVz32EFcCamvhOQe
YNWX+HWk2ou4HRUzm04rlh/BgBqAAlweNtXVEEtLgA/2GrwmDs/riIbnacXeK3Ye
QSPq45JLGrkhIJ6SQxntM75wPgeb2mAP2nCSIweD5kLjYKQaw0M56X5+X1CKtgkK
TuQgUw8cNhgx4FfGxpSNxxZARHSlKni+YvfSeLRi3jj7s+z2zWYudNFDa3WYaX45
QvR+fYVGZmTI+uTqwCfUK9Y7Vwi2jBdjvHT3bVN+o7YCk+/0ZPAQsSEV5KfEAED6
8YztGYiIOsYYKamL93jhhjtu/XSLIeazk6jaJeNAc8RncIZLI3bnwxKLGOEs3dJq
j9UvwnEvw2+eLtpOXKarIQXR5d573/8gL+iBsB0O/OUwXq3/N1BbVCYJw1APZZdD
mtb504532oVaF362c0Ik8FACMdGBtde4EZIl2FC0mvRp1ea7ZeSUUb1ZB516Qayg
CbrQy7MUH2xIfwOK2SHMa2mwvmy6wx+ySTzUKOJFWT3KnIAqIbO1nk6tqBnLE8Oz
djFhsErsJNhxi83un3QT4XAJhljkzz2n+Y8gvF8ie9j0M1T2HbdhlwX2leX5j8wk
tze4vcwB9V1HuQ82j+w4zUdPa3aTIpEP4WimH3fr7/MJfhRXh9ygI/7N7YW+OtyC
hUKSW7SC0wChnHsXIlNVgTRs/OcUWmvU4k+OXYsiGX/QFk/chynrNI+2/A9UI/Ui
bnBiKssTR+yHOr9hm+Q9e5GlpkvxQvIRS5rUMbCdqV++08UbqRt8NcNldupmA6Gg
RqUY4dOQ7IfQuOqN+czXxiwhY7JgJys+auA66gn+aVLO628xEE9J2ur44f6qmlyt
deYU6yzkk1sA7DQhUmINDbbaNOVE6SBl9hqvEnw4bdp+p/OCxjCjHt4c5hZjY98/
nCDpZ7sObstig1pgVwmlTXwSnvAQ3TjvDZRgEzhAQPN9u6i8IKMwYMoKO3OXAbgl
PgY4ijGnGGbAUfEDoVqtDqZtRYC66Gd2mc1B8Zujm2/KAUxofI5ThUOUxZK473hZ
vLjJE1d9eWfQeRi4Xymlibid90Xy5qHLz4R6qYH85vT3kcyXHNLaxQepzkrgfJsJ
gDiXmLvvh5fmgFGxTkEOVUviGlI7ovbLLervPwN4Pg0FIBx8sIz960kXqWyN8Yst
fP8gxfodpHUqPO2LGFEc3Qx2ogch0CjKHx5PsyAz2LU5nwjQ6umdi/TjtuguPcAZ
LnKzddTnzfvqYgGONb8t64kc5YKoaI08BMhR5QVogjAlWBaIygeMki8jzDdUm+hE
dXjL5fWMqe0gmjDOW+9LsA9QVOPnRO7rkOdNMhy650BAgzy32PmSDlwQeZ5TJuv0
UAGxazYswAD141R61JAgLpeCbaXQI8/mFxM3TB7p5PPKRlUxfBa+GhDuy/RoS7JD
DF6XQsqN1kgVszy1yUJ+n41D72UN29CzoHKFmiHxFZZsOrx3PGR2+FsGAFJNAD0j
Xrry/Yk95YTD+1Sio9nt3BCdvQpPWsCbr3F9VmQOA43fehA01vvgJZ1BGLOeO6Zi
IRjZBIx/glk8339SKb8Rj7cLyj5G/l60OPrCQ77s3sb/JIA1nkR/gFlPVcnB9O8k
qCSsFdFMScHWJZKcy9B9heetTVq9r1gOUfwgx3pwWi+/h0A1xh9wKvW8ysBUYdm8
rx1pDEfwdnIiPh9ow2mDRKWUn8dFi6a9305WnSwZGJkAE9ZTPd8/Ztb8KkYqtEvb
J6wFA0/wRjn21YR8RDoqEeM/xHzP7ht8zXjkOM2Zc53dfZGBAU8T1rpcLhxmY+Wu
neRlKbiSfGw2OiWcxtIFZrWGXjducu/6mjwxprs4rJLMqOCEwpTvfWCaFAGu1dkW
TYUfY0WK8auz34nNNxxnA4XA3zlQCB9Pn+LQJ7+EtUopqegovx34Aa4zQ+jir/50
DYP+AclL8zKB9frDqJTJtyncHix06zdmiozMdaVI/DH10yvBjMC0xrUodL1s17FQ
MQbu91Qos3ZKWNPy509ZfU6wkpF/W/D3EEf/L1uGTnQ8UPtwAywlQyYZcO1IscLx
Dm/riy6HE8AawoHn+jjo6HWii4BZ4c/H7Z+gH7Cbx2hYbRp1CIVNdBDbJUzjswOC
E1PdJGaPdQR6/1H+jgbPFR0gx18Q/AtcjFDmQgbUZASFAxCs+56yPTD4JnpY151x
p7MWY8NGYubX/b4nS1H2VNgNevjI5+2qxp0xtA18NfzUOI8qt4xoGweNJsyc+hvt
vDNsf22N+t+uAh0pFSqCLMlx9HTyV8o873iMy8iKHFiMEIrFpZs7wXIUEposl2uW
oF9SgXAnFGPPObLH0Xo8HeOZhfX5PFbQSF1D5sBK67GMGk+0lanA2Ui5jCnXETL2
FnrO2nTzxpC7RYd/FlwNHOWRwiLicBLBCn7CTm1KSotW+cmjjSqmQB4w8nX6ARaX
bHb+rc3b93NwQcRrcuPxISq5fT/kBYPU8a6u7v9SdUNQoV5H8via8mSO3yjahe2M
A8e2M+6fogXFDkAtP5pXDaTHmm2zBgp64JgfuaOVXhoJ5EhG2WDnW+koCzQV2AQQ
BEQqth8qeXwUnHtoMEKIKGoLCAH6qefG2o7YJY78xbQ4BGuApaT+s4Ju98FweASv
9/J/+Aaq9pSnl7wARP+IZYtCMX5w5LyqQ3KlDXQUp8o4pTlWq2zmkcfOl2eST8qe
v0TeQCggFm8dGeKLYN9c0cjXmrKNehWy4eV7fgciDlgV3WZwjItHVP2Hu8w38LfD
9rgxNe3XnAkAqH+aaxB4GB6dyUMRA/m8Ipz54EuHvzgRs8SOsrAaPCwSocTsPIKf
rDPVrU+O07jXk+JpZfN22IPnPCQ0SQU97zs3kYDrrTDQMobKl11LVhX4nUwV6T8c
tPGxfnTMIOrH42qx1Wx8hx+W51WmnULqr7LPFCnxhj6gnUm2OY2/taBm95OM+auG
to5TPm4VvxqF6dQm/hNu33eTKx9SR8ERsMRexc40VMH/65pe4sRMkp1sZED4rhQ8
CNbJrzRNyn12STyoC49zJze1rxohIYfkWQl3XGiyGySCXDhD+mKAukyXekv7j3eX
rU4X+gYnaJ2Lb/xrZihzkUzxqDmWA5+9dH3buS14D/SZ+7aJwfcxgjIaidpFFd7H
W29PN8KPC7YAOCyeZ8KYbt0mOw6RCA4lrQEPyNMFKl3OhmT8MAPS/NeKEXBmHX9g
meth44D+8f9YSMJdj22yk5NueEECkdgk9dYWLrbhqsxSlSdlPWwLMooX30+9kOOK
iJJObIJmQ5yoxgsSksKZiv7D9iwNS2K0zqSRpibJ0vjc8MRiqXpIQWfh54PpPOff
WUNKqLBjoDHw1U0pR/8LcKRQa5/BkSZ2aBtihh/dvAAjQP1TzAVY52CE3MUgFUtA
u4yyosMzeyhcG+EWQXTqqycWkOG1HxjozbzNCQmo/yqRWDcSsQihLCdmGGMqNOdY
KY8p5/NDx+99qBDKfCuHtbacUaItsAMjQQb4DVgsvGZFDul1tF801Ytr5UDDsGn6
OAU2efDZZYlKDXmFtJoJ3IIkanmCGEknNgjNGAXQR/UEZS7SASfts1cl/1BNMxw1
cjvLTrILMOCSiNKOJnUHyKVoSqkmyBC0YE2DyaViH6hL7X4LE8mYs8qlYMIZr9kg
dk7BaCvGa7Ff0hgm8B6bibGflaJxIISe8JYY9K+GrZuIoiw74srNiqJb1Zhr+Ntt
vANtibKCIPEB0cMViSqjpZ+oJza7zli7gtz0jQ8uIG9Q594IF8nnmUFwAZI7du2L
ChugjeQO2xkcl5P0/zOtDS+tPros7n7eJL2Y/+fXDOAWIBqsOxr5qxvaDkiaLVY3
+bwCx92Bn7J34TpqQu3TWRjJgz+T3nMeEGyqa5dOmHE/FDBD2gJJ9e2pg6IonncQ
E1jsLHN3COOo0xhFEdGdWIk16mIkKuyPIbiAf10qy22zS1tfyTszx9qSyhRPaKXl
q/dum4k7ZQNCMY1DNIU74jeEXkOmG4GyWuk2d4VlP0bxFcYBVFh7fNskmjiqSRle
cihLjRLVvT0m1RjQBAzKYViA9U9dZW+CTaeAYef6R+nIsPT9D2EwVkiH7ispMzJl
sYhGmTcqdF7IDJUtFSYK+OTWGib2oV7KlLWiRffhh/PGcSb7EVSlbeaiSQnVBYud
3N2JROnrIeZ/JXF5V4GlkXxjdUS/hpUlSoDkv7hOiz+qg9uuGdbjKk7TS3mECW1/
2xSovzHfRc4UVg7k7HYChHEEsRKZziogkjdHLh2K2/YoptVPEAFfd3mdxJZHuRj1
6mUH5gLIYPpSb0XqKbxH1azHy/1cSuBlLS6W1sz4uq/aqr7LV3yymhl1EkWMl/fx
nKhPhU9CcB/j2mcuQd1Z00iDv8aXSvulSVw3Fsq3Ju8dk3i8sU/QpQQ2tf1WE+/W
ncHwjOmkdtRcXqnY3Hl7Fy4a3enoPFY3iMkBzoDmMz4ji6zKULe1CcacEaPJoqna
zsa0ap3+mV4EVx7Q225hst2Njsb7Yw40Q8eoo2D8FRl0zlkeEkW5i3bSyCL4ctMG
kXCg07yluP89CsbqmO8s3nhgbEWgGcgEOgy9N/HYLN0l3aI+9TKZzJXG2nQaYpp1
CCZiK2omQtlFRf3+dqp8IVQqJ4iPQBqhko7P0Lxu0ypjTJYnfULI344irS1SRzNM
992JT1FpBJL/fdLnm+OpOz8yVo4m4QTGyokcnsY+mzpYU5NJyIx9ImZNMMLml7+g
juvwAWsGoqpZT02M55dtSxEA9HJhow212ECvZgPAIa+gRlUF5lNWmEthND4NGbKM
EP3a/8lkop53bFRBln/qlJWNXmIneF5gTww9et3V47H+4l/jumK4fkIq27AQvXrv
auxWs8pNHvnAqlD36e8xQckRDd7BijxjwAwNa6lH/6wAsbnZHhSeDe8NtV44Dnvk
EicuvGmXZ/w4PVMC3G69NdqKMUN4m+sQGLPlybt4UnRPPHTzeNn6nm1Dq4LwWJS2
8UVebHxC7hD6zAqi7SF8H1ZgEpByrE6gVxlaa1dvpSVFyO2XtfFfp3FTmSUHQaUU
pVPPCefguGuSMF27OW1K0X4AMZRM7rsgfW/CYydFXziAtdaZtyyiezFSw3c8j3Ca
eDwV55NxoTChMYR9RNEb9gncFuPr4NWfWBBCxTulVZlson2ZyfSy0BTgqc3R/OZ9
5LCTEQb0wkhkbnmgurVYOx/OiEBhWv6YW8WSmsSxBDkt9J2g5yI35pIfwKvbKwwv
XxTGOXMHf/4UxFBSoMy7r5dc/Yj0NB4TNbKoub4x85RMxgghTd4vLBc2U0FLum3C
2p8jCixobMlik83BML4uH/eFFBTB+xdNmgG4nlDb/+Rgd3Tj//VSDSu+aMuiGFb6
hXEUBnA1JhmJ1w+oQJ6IGLisKp7iuGAEFJ56YDElarYQoM1ZYRcWD275axRtIkPu
pZRivrB2S78r46l88FP/qsxnSJ+nW8ZIyILUbodGZynAa6BgE/GK7MP+hTGaqLUD
j6EZrsAh2b3v60WbciM9nExI5zGBignOMGDTRv2vn+V+P8xWAQvpEE7FnBI33vJ9
lQv3t0SNdJ+iMF99WWTaet602d8lR4sRVPQ7hw3VQxXnWWCaXMztQmaT82GZWksy
/wnN0wkycX0uzaDnM2J08EsUf1184SldBFnpMhntxswfNTq9ko7p4s+wSHobVJ7p
9mGwiKjyxWITfHH/9Z5wyGXJ8s87y/Qx2ZQAvW3JZaPBsDeOZCcaiCp9cuhX9y1U
2i9w5xI6bM30JsYmSkvpAzF2oZXTbylrzWI2W5PK+UnzmkFrAGr95AFbwIMt9TEN
gih3xM+qFtFX6wN3kmbrVhW6yGCw2zasq2cKY1itXsMxs11nTcI3bSu+uonm7/AR
eD2oFgb65Vm7t/oVrnzgWWh94N5nydBgkcVqilmf2yucUXz63oQoqIL81MMNcr/I
4vMBYve9zBRxftdloBYO52EPsH/Htk3kLT8rqH2Oi587ZSbTjmii4WwWQxdAL3On
NusZHRQQDQ5EQW/sMh+0sLYN4RSTDUY/BIcBEQxF++XYScU74n77yAwMae6G+KMb
6PvJFOrPe0LMyNOO1uX5/4/j1gC+23Fd2hDGAi/kA7FgChmEicDE7p4gIqAsU4XP
10YHLCa+vstJPLSA/86aUno+06ZnCXzWpYAgVJmRQlKjDEFf7OUyd53ZzQwIC71x
IBO7NQ/IYDbCcKZ1qSjaBuTYST1ddPIghAr2hKr5o5woF982tfh19iwFbitkItVQ
mxC2IDBeQH3zQb0htSWgVtTK27XMLnvWKyllQIpTI0mn/Kmzvt/LlUDqUPPV2MUl
f7xrMhmPDiqTZhBlFq0eaiQ52+gdQBFSuz82i3xo7diPBTdWPGB8HABSrrP+mYFv
29m0malNDNlN2vfomxwE2ZujWtPiP9kkEe98oEtmax+EqPJaT40uvG+m/Dh4yL4G
9nH00DYJpdWunSNYNhRgXiXe3Qg1SeWBQL8MArN+nEdRXUPKr2Ajw77nVHGS1Bm/
aFls4XIqh7h2mnM6GPBENFeSDLwp8Av99m6h37fXmEL5WpHk4+/8BWSXm7zI26up
n3LnDQedFNqPFQdOLXwNwj2zkuZCJmHuAt4IrkSxUvQP2varlFAvyS/rAJjYShpM
F871pQVquqwylps0L8MUuOsInORlQ+WI8nwM6maUj4XF2qD5Ohx4YPk504XrfP4g
b57xt1aWL6WPxePC1AgQKU3QvRsM63o0fbis3SUgowt4zgarLZj17yQ04pw+Jq0T
nAipYCCjDr8gixW2aI6j9VshSX/RZnf1zaYMpf/HnUIfKpNpBL1Q0E/v/rdPBGsQ
cuiI5P/oKqVIMmt/7HlCZ8V7jHG9IzD82kdxcKcePaZfQ2yL01BIhp29i0lvC+NU
H7Ibr7NI/nlpk7sXTuQZg/K5JMG/mxFVVTH7BGhy5wGRNnDLNZNj2OAifwLxIGSm
Xys4OQe1NjTcXco3ZJmzJAjRbDt9ny/TpoyrJXTto7LMPOpJq6J+BeOSiRGqBzmh
RZoPqy0M20UINJeP00A1uFuwau2eXoxIhhERCohLFydmOBQenezWlhDgiNDKevKt
7u53apysLebrLzCMinkLuSUNpT9X0NUaHWcCAKa8uf02A3BetIDBXiDBdvtUnOJp
yZ4ln4sp1jtG3+Ev0NcARGbcaroUOomMIn2RxNu91DgxHiNRJrvUoKPTD9w8FVwR
N80Pqd6RCwFj6l3th88MJC6SET75ANsoIW2EnJ4p2OjEZyfLgbVt6CGc9FFJo3Vm
BDbOzcW4EVDRK5Q0ogmnK1PUj37C+ONBiDMVKO9HyKP7AKMZjlwPmIS8OL443qty
QKqp4HMsu13ZDC8s42BknnmT78ksH+p5imZh85GvdApZ2gJwMO2Y3lcCrgbNwqqH
EnomMybc5b9ELO1JvoDGuaQI24hzW3vP8f+Jy7HV7w2dhW9Y0McHr3PstPmh/cRT
lJxGYh1RQEXn1QVoEgmR1h+5fs7Y1eLcAJfkUjtzX1Ouga/c5zh+r/01q3BpEpdp
Y2CtuT2f9RrvSkk264qwKfxYD0xommG6I700V2Jo2+tIkn+CXIrTPTes9ZeylJMW
lKUX0SqYWjTFqQgmaAVIElqCkhzoINyNlQsg6tSGkNR70oef4lWCDgyU3y73yTpI
lA47ODVFsqfNSyKPgeor6JzuOyMEXyzm1dqAgdunPbocIR540zmGbdiFJZm5KlKQ
ZbkoMKYXlE3afWH8bzd22pel4SWZMpJCJodMqeMbu4+LkO8tkJ6E7gds4xoVh8p+
jBiFJIKRBwErCxDY0n6hRM5++S8updP2Nuf01/nAka2b30fC9QXqyAg4sReE2X+e
+CzCKiOa8sgpGppAIAiPBd8jGZEQ4px45umUZKAC2e7RvQ331ygmAqqccoxxQyn2
C13ByPexN1y3ZKPDMTe/pPcZ6iaXDa7zo7lwh4hWQbTTHI8SRcZkNzBX8VzMnilh
C5PEtGcZ+su3I3d7vXjmFnNpLvb+HGHl30CeJ5XAX08m+ySDjK3FlyRSbU3QhEG7
WCJSlHRuGAYMgnsrneN0+UlRRxzZ0eZSAAOCBzWIFnZ08ShV1f1O91T2ZGxRudZ+
5nJXAiRaBAUFvfP9hz7DxFepBJSO8TyvNqSf74egLPgdkGvdoawwsmXfyOnOG3i1
NkvW5KygSUVvM9FLFoDU/VLb2FFdUGXVIhGXJW/M8lhbiQJUwjz24cNyzDBBWhSb
hw0LpSxl8MRZj9DPZDQ7aFSTE5rtuUq+emXUXfd7j453x5uGMDmuWYNnvP9q6Fqi
HtNXr547frKOuR3Rq8/GTztAdvRCc+uTUh47OaCh3FCq3lH09BakaAObDQqtHbo2
ji8coC89R3uQVqY+vj/ae+eFvx+fIe+G0Q3MNRDpzch3jxcRyLptTqXrPGpk34GW
OsDgVjejXBa4qsmgT9uB0Nhp8nNU/IcHkx4XwJEnIHidHVNmrgQCsKky/ebdIakn
KSUWONdMwV7A1LOpy7Q4D150J1t2RAuTWVTMV11QIhk3ZMHuJI6vGlMTYvLcNcvs
FaWTQbIcZHcOrNIM5gT8MOTpam0d6+3vSQhV8hwDlhXkTf+5FY93apkKNrQU1AjG
OIPtj6Xh5eaiUzm+bIuDs0tUG36WoIu/BNJluUd57rK7z0Pw9W2voxHUBjRy9+wZ
O3BsPw3yKdkWvWbRMrl4o/ZQGZBnAHOxhGQiznnWzWqoVKr4/M6GLtFCVyxn9psW
Yf13UrWxzlsLSyF0nehEpK71D/ee+Dn8U2yhVSvxJIbT2WnPgBfDP0dHejM/0dvW
wyyeB6tUEd2ALxbiNquq2CgVuDmdawvrJxdSALX5fCLxbWJ4sjWS2CkFEpz5Mdlz
wnkum5B8LUaOEsaG1adQb62KskVAyFFq7gES/8U8bNDix6YljgK0WrpobvwG9GXL
`protect END_PROTECTED