-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Emdrqgpu8QjGa0jYrqZlwUdnegQGB0aAP08MRqW6YqcQBqskd3wMTQWgBh5h/mix
w91GYzfXNs6yhe3eJjMwwt7ogbzq09hBGxHqI9b2RCmn3QVUUbZZY9b4eyB3W8Vz
YzQwsje8iIgJ3jdsxlM49NcVRA4lGdJVKqljaa+MJ2k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 111456)
`protect data_block
a4x8Tt06dzT8cq7g9tT0BmOfDTYjC5/G9jaIMqdWvZX739CiF2H07O7wNhrWtZvt
gmbBwVjdiry8qKscedzBczP8YeBJFx7SX1ToKohaAa4vSLULyeSajFM4sM5CXFD8
+t63cUe7b2yAhExu5LbrYr7NLPUTKsNT7lLYoJXC0C3C0pDm5OJ20gRUXRGTR2hd
WIP4kGrtTQIzfjTZ7ciYJ+Rk6K0PlpEYlWG1sXWtM6lbRrMsiFPpkRq4rKHVxhHB
zRREgyBvFnJUe660NlllaXygmfP0cDcvlgiBK9NIMmrwCByxFZNIavgqYdJOL5qj
Em74oFgkdLmZnzyj/IIh3le2ChrmNE+ggT6r4bvRhw6ZmqW/qJch9/mhcRzV4Byl
wxlEwma1YQLHM7NcGdobBPRljphGMr5+diiiVLZbNMqiEZY8R7lwwi/0G0SgGjS5
lU69EfeoRX6/EpBNqmcjByOt1FDpJ7OJ3zZLcE9iCrqj38BV3rolzvgZKPpNdFhg
3jpCSzpsv73fu71V0HNqZ4/Om6AOf1pmT/UyAi1M0qJLztC7PXnTi1hc4syYPEvU
3sC5SSKhNo592yaSnovPSYBXRayGkZcdRbeZK1z6R8pt9p1FqsyRvjkwUvP6Su27
7sDcMLxk83CTYTHdzlZBRkdfaoANpeuyQBSJRqb+3I6oeJVMjqjEEDZgyN/bbxLi
t/UlrgK05DXsvLTwpIUmH6K4N2kDWHm7TYZGvfwgu4b0KAGYf8MQS0pwc2oSeqAl
MIcH98YNHuAW4XD9MvzOAmC2zUddLGiVPnpWBAK/7Tyt0/LM4X8T6tz9AjeGAe2g
mdQ4QC29os4nvCQQ+E7pMwG4XBYpmnYGY/cN4eFhsr5RFGCTBJAApVqazp3wj4bL
tyd+dbsV+rIwRutjSCehbVncHm+H8noAoFtY5QnSgXI21GhjzJZDhMGkLqAqNcod
u+aQWPcFM6nlHz9p03luNEhenmnQHv6wS0p06VK635h3GgT6L+8FekTJjMXypwZv
eZOJqSZEQ5PC9W6u2Wu6NgZ0g09tBlePnmCUA4d03v+xyY5/gVJFbyGWnS7tYyDv
luWUy8GvjWFkjKNrImfUZ4WhtwK8z7yVKVFaFv+jfuLF8jNJk992mZkfGryB0yFN
66wCSbphkuiZBZ6rWpjEb9uyc5/6A7TWOxJNHYDj851uzyUztPrK5/+9jIKNvcny
68FBJlBJ7ZvGKEfRbzTqGwRJB2egUyxJFgyenuOfwu6OilLQ3MTT+Ag14sMRMHJN
tUip6fIOdbfdZE1W196zMljp3IRQLnHlfs5fTcZMDXoz4R0m8oxoGafP6cLD59Fc
Pj6Ack386D+Osyozf0zSFIe6jxbd37D5G2e5+Ii4+QTjEq0L5L1KBjVGNA8O9qtB
sZkhY+kOGt14lQ7QFefdSpBAwKGwSxk+dbqdLNrbfA8zbQZuiKkaAOKgtg8fdH3l
a1rJeuXT5WN4L7fIt2SYXR57vB4NLvCYVx5T2xdZUy9NpSUOzzLleetPvQPPmQMt
Q+dDLfXmday/9CjkuMMmo6ch5hOlVzxPGBtcFGQ4UCYyocYnLq1X3TVc/rsxUP7c
fMBnmwO5oQbzXmVdn9VfHksYGWCAuA4adI+28jlc4jz+eiR9w2V8BTO6I6DrxPar
Rdp/7I3dEDyw1DbWbgtJugeby7z5tR4Rwb3iLBrCppm6w0B+yn72sJuOG4iE17WQ
8r08dW5rgiR3HBIXzL/4nt+3I52c45FxtXyjxezO+77FZE1+UPAfuWbT6VZrfhmj
g6D2KkOSzbLUPfjWnbnROAGkACa6aXP/ClLNiWrhRCzPDb3u3h0K5XWKKfJtVSoV
UdhdJMGu4RapW1CqwVGKtkaJ1i6w7nMc7srZ1FkwuGmZFz4ba3lmHJ6YlITBFiBg
Ey99DTm95I3J0J15rZJnw5enHTosUrKP4DxLj0uub6PvgaJHy8pxmx8Y1uaGyhig
kDlZzyEDKOI7z9u42j+s9bnQfw2h1Z1Xcom10Z1WbNzxoyl2r2GRcwhSWtTPHU9/
WQXY/e4y+w36iyDKGJdfV3BQgUlIC4Ye15DkGiFDpi//c5QNRt5eg53c1reNoya0
cj9inamCUkuckarjC4ZSLkPufLHyGWAqPJYoK5QGpsic+RVdcj81/fRKIAJP+t90
LWSNYXAjpI2TjCEvukPuM0R0BDm8n0GYVhcEVMR9R6DcWbU2ukHdM3S5VzmdFmJm
NKVbfWq8dHTw1kooKkxTaGKKa3XXYQAYluXOQZovkP23UNOuB3gb15hU5gwggaec
Er68cB6CgdO68bEYGVyLL9ZfssaGu0qTGmR7lqaIGJ110624Pweo2UjXr06SJK5I
oRB3lIAUYyQe8QQHMk38jE8rLKsO8zETWjK3JrkeWU/q/zq9ibQZ0MwyWFkmUG0a
gGEaa5jey+0jcag9/jiBU5LOj3qyCxPzNJy41sra+xLN3Fcb56kNchVG4uIAlLHe
EOAm+s6fyzZrJdMlq+BZQhlvOkXofawO3IeWJSXlIWBMhgjU6fbCrO7+sJG/KbBp
FH4eVYOfP96yUOd4UShMXLYoVIirO104PWFXOUTkuY8KVfT837fkbvAFoawjEyxP
KVCaGJg3gZ03X2WRfgFTj0+uZKBP9TBIfbbqJBhWUp7Qd+fasVQYLox26l9vvoT8
1I4YymGoxRXaz6/kZ13JrKtoH9zwQbaaomLbm43iPRO6SO7Z1ReMkmEM0xr7Uz/o
U0sy27BTAQs4W9I492Rn7Uz9JDSwquIT5oZT2HjMjY9ARCKQH6FqjFYO01v2tVke
4iq8/MEMCmJ/04TP8HZAAyLxUgVdHwvMJB1uZTgA77j9231lAT4jVsxsk8qWubBc
wXkPDL/MbvkNqJAfAdCl79EVS5HwPIsnO6TY1AmMnll8GT3/jkjDNj0ilxI+A7zq
t7Oj4blONhy0T9SWYOxneBBjfE80ogwaAqvhw7+UAVDataSp9oUMQ4P1bjaR/l0I
jWaYrTK8iBUuo9tuZSPk+CYNyxfj3JHOim5uNCxtjYAeLmB0fWZhFf67TQDlDTVo
viBKOqfxjNLm8kt7pTw5LP4UYpREfOFmhsoCswLB9gbjMtjgU1sXqMxu2MVE1Ix4
5qAWUo9OA2uoeJvqefOy6b/jUSuyfWuIdEQKwchsNnEgSBEQRqaVFzizBYnWJ0Hd
seYRVsxAWJFpfzOhDLxO9sdPCQ+t4//ixDzkx4eK7RekwAHYq4XYudDZn4bOIiPG
EP9uETUR2UYBdJqWmvRbRJImdfZgOeL6jy/DiNM+Wt+PUEJa3YI2ZwY9HLCRwFxD
b4UxVcDVNqKBd7wo5kElo9hu4knwhQQwpxQP2xXSIxRMxMNqoSS8FVwnIxsLGCcy
BM0F6FSHSpQuqpZ/DhJfsAelS44SY581o++V6OPDFRw3RtfOeNSA/HeVEb01Wtz2
Jp+m0wIBcoCwi85CjMsUc6M3XymDr6yrnd7bhfTfCWlA7O6I3tnIkbGOXOvfmcNN
EIlgubzuA87dVnEonZYm4vfi7MF3SN8XgEX0GoBY4Md+AnWUwYo2UnEq/JXDffGl
K6hITjknU//qbfK6A/L9j63EolEMmyVaF2eECEtLvca8daLxSCZkXcH8SOWBJIxv
UrVe1bEBcofT7APe3Dobs59B8RhyK+7RWfO4Hxpl5eMuPcSunzyzddk/uI1KWP2Y
TI28uNdSYouM2tBJsbcRzCPG25QRa+yv+TwhJ6Kcv+726LaBo4JpWg7dGXN/++fs
Zj7qIHSemZ1yThIwAG+TMBeIMvNC/Wbi3chzxn8ivx+/8u2XzvdhABwTuezdwuGD
pxlOgpK/1yADKKX+OOv6Vfs6rK2HRCeZzgbJ+qSoICIlFrcRXiurs0ntYGFlECFl
Egfgs9SDdalWhbCiHp1fWUMeYQyXk+nY78s8d4rZZXgTvcRTgMKEkcbiC+DMxNn0
EF15/cU6hhK1eWA6FBJofwivEX7FHAwvSeGUCFF7mOSE8OuEM1+ETot0uup4QfrK
ihEQdZh193j8nzI6XK1/Cb2ZbnR2vBLTlGr5kK9kRI4qj1Hq7e7fzb9LEx7jnPLU
3d1fWiACe7QdeAgMsg/7WwMCrNuu0Xo/C+CcxkR3lDUSz8Lue2qVySpJYk0EbTOO
v81ks5C60SxdaE90sruh6pfMmHq48cXYJugDAol4HON5KF6tljgojxi1NM1cHr3U
8msTRbSJHyRucdH5C6/0yjW1KAk7aiaAHsXrsBbBlbkL3CDDqbHfreYwoDC2lmZZ
wGOdNiaKv5U2HAF9mevTLrTiTkDCVbHsDZVccfgX2iXyNwJNUSHW3oJIwaqmShZD
BZkrwzc7lNYDeoH3XZ8/ugp19jm1uVWKg1/7pUPqIuh8lXln1odE9r+4jMXcHjL2
rInnJFTA7B0ABiRV4NP4vry2L+ySUC220X4DdxTMbDFPr4CXjFf8INx7YZbHsUWR
d5Q7Fu+w2o41aAE6t0nxPCzE5EOU3KeTygwuiyed8x3/6sRUjmFjmcGXUXZfCNHI
wDSQSHbhJ+xWCyQ+yXrbp85yoI4HCj3mJOYFTsJQhO49pF26GhwHMo/A42OwT4H/
7awpVuECmigBFNyiSDPuyKBRIGGMNFwpZRa/8XI+I/s+NWV47/IXwzlZ9kl6mEK5
PEWVCGVyO0PYN8705pFrsREPLNEOYJOLHnZL5HxLGJdc6I30UcwLF0uEsdrVgVIL
lSOzv6jnM04gyZoa6k/zSF54EAmcb6hCIsm/0BvOnfAF8VhgVG/SLlHYJ1aiRHV1
rnt/Gd8HkKgJ6/Ljat1OV10ARQi29r0Q2Cle2wwIHMJZp4xRVkCE+VK3SJCachMr
hRoVpUPfL2N5f/hmtn+wuYDFYirxYE0h3MlTPzRqfCWBAytAZWfcmwN98/EdrCKb
tLBC2Heo3vaZEYCKvNTkMb81hTgosOVAad1Ha/lGgkShwkd9EhM7iW9yyGyQT9Wr
+VVGy5JCLwBbXP/+xFkC2N7qcx2iU+SkWmPmxL4wMiGsxUF+DKsGXmCzA2dtgQSR
v25LG4qIXf779v/dQAmekEqoaG/Ui0MbGNhHMjm7UwXNzkY6s/CUV6XDEpOHYF8f
VQwxD5gzKTZXaXcmhmEd59arkJbWREx2m0IB216hu5ciYdxOGFzgBshIlzxmi0CS
m6uAK+XcMt2Mqv2/qCWiSK66q7US61/BK/D3oXNaggvi9/hKiYNEJw6G2OuKHshr
1EN+9Aa16/Tvi0XUK/OAIfOHQ/Q4P2XPXCMs5j/jQwPFD+U+sSYKGkN7YfM+Y4Pm
fmoLhr2XsQnIddCj+XSzvU3QiEtmSXEVWlsVtuVrvMqywruagfXRUfa5Wzzd6kAk
gHLVsfew5wOzDaQ2wwvEVT3ql8XUPlQOHoRbRL4DXZz0QGJGlqu1WwcCeDrDn9ew
Xd70lCbxPOEIL1Xy/zDEw3We1i+YvhL6BXY+kihpRynU5YjRwPa0Do15ZJGraASi
lCS9/BkMLY3jIZpR4BzjSu22rgHRXsAqLhgZVi9fYSZoXYEyO1F4iaXOBgJptk/Q
eOYNlKA2LTGMTppL8OySYpRyA3Uyyqc07H9V+d5PEcuzsgbBiojTQIIylUjQzqq6
nOnnOyEeVx0s59fElyFnv6m+4piIql312QwJPVE14UwEX+MQR/z79G/XcO/AWurZ
PwpYHvcAfrCcRnlxedicqrk2rDNvrR9j61t18Vpd0Nms+ty5CjWua2sDyosQEYjb
AG6OQrEcjcfbMyAzaO0p7z4v61OfrYq66/vIXb2UCHbSsMA4iOpq4UEo00+jzCiU
qr+nq+Yu86U94XK8r+iUOI1dqwaVoNu+h6rTnqAzOUeCbdJgcAUGHso0ULE3cuSa
M+VgRGXFx17h0xBUzKoYSt+0/UtmmGkgmc0aLQWoYPmUJ3ejyYMnu4b2tnT9l7pC
ziqcsOi5JxfFuOp4TB7noQrSPLpVp9zQ1TsZw8hcLc8hFl9Zypgochxq9YtKcEMs
b7TlD9JjnL6R9+A3q6QzJaKuLhZ1JYGcyjnxrroCPyDre3fKUEAN1SFOWmmf2lOs
029ruOwi/O6h6pvX7tNYuxM1uwQS/wvcSZiraNvX5KpYbCq3THDQy2ICTY+4x9e7
TkWcM8I4dQ8ED7RAhptYuJuJnyQsMPD8RfWZl1omKUx7hPChDsUQhB6L60pfVboB
NEZ6Wh/xGZhhUqTRJ+nivP6eLoiz78AgMjIllTV5LajZNna6A/wmTAocjFT76W/t
XpB3hmbH5cWkkC5UPwc3gRwpPK8Tc3xtY/KLCrM1rX56u0LZzNqaqqJQxLJ9pF65
IP5KgKzy5O/MgWU2zn5we5L3d3mJlpUClY4WjA4fBG6FE0W2cni1kavceTPC+DgX
UrQKnCBARaNoP6rZme5SHoJTwlDqzeUJpyZ4tKXlP8eCDRWlCfs71iAQR63KK8zC
AAmmke2k6Qx5PZXWJ/Nd3QMXa6iX2UfeC1c333nRbIaTErsvfR5r+HiOInMJmd+E
qPHRASLOFaS21HCIcsVu3n9V3ZGrArEMStX34CbuiktT9EBZj7fRMsoglhLa/+if
BIv11gWOeZGTZe8uilb43TdmYrQRYF03J4pcZjHD0Looi6qvuduAR5aFnQWK5X+9
1wjJRGmyb8zJc8L6M1oLCejg0uUxF2Ys1Z9YqInlBUwpSwjca/Z+UK4Tl0AAxTOd
aDqSdvERGAFGW4vkJHelEsMnDjQjTG9dvAxVoMiX8waJuguC8B87osNf0vqc3RtF
73knSg2BOIl3Q5bOxKsP2ZxJjw6Sgyop812b5E70BJRIEkugD6PEuOmbSoLTGlJk
4V4oUGdAIjhEieEo5godtBAwndro1PTfND5GKatyz5M4oyE5yeO4Pb35eIjXWEX3
/UFV23BSSvddFQ579FvDr9+5mORN8M/xcO71hwpP9iis+qzEm6GMxDoQjLifTCXJ
Ow+cG5ujd/e++Qx7ZJUSG3GU2Ylu23nxah6ay3w0xzbwEU/RJ7NxRNWFfjk0n6YE
5gVhSM6cy/ltYLqAHx+uetohqCQyBAF+AKzrEnDUuo2ZBgFJqpnEA2TKDE+KMRBm
dLt6IeVbOn8SbS+f1+GcITy3YVMnK0rfa9XvmxrYy4WIu/jPOAf5Ou6SIZMMF1zX
iJq32SbWKZ/vfxBjVWLtcAd20exJPGRh5czO2XKtH1IKHm70+vIpMsrDCMYBE3Ea
TwogIZ+DqLROhoEh0p8TipRhLjAJ379YRuSD5uPPL4A70u1quuVqkW8F6mZvv8gN
xn03ZJWYaGWVxSfIdov2w92kMIde0rM25rjuTCtYQ9cKJhmYnzud2FKtZ/psjgxy
Z80ymiSezstSZjxRnH9Hxhpq1haz6TD4jumBGZMro6J5i/YQbfc1dOo7XIrl4Rhy
M7FEWv9bk3nisiJb5mvyXZBjDKUmVIwrOYRqAqMh6vS1EF9hKK+O8wBFLF3rDsqj
BXOpM/i1T6ea41Tho8V/IAnmbtqojbLmypWXZXMJPUzSILjpx9ang3WfayFn6nli
9KE41Ay4wUWmNBsrTvQzQU4gesQtHxlGDrafXpEGJvejqaHyGh38fBIvDmiyi78L
8GTvy70ffGc6DTw7QhcT9jgf1ZsM5DcCjA4uL/hpeHS70HPispQ9SGvNCUWMmxY7
wuwYeArx+qBMRATAojwibvrp+ezeXqGcbvm6JA0BweSdfchPwt5wl7gET9GguWOo
M7sWdIiIWXdzijebw7vikuViuYTCN15J7OVJmHbB5jHMuCGoP7Zf1doi5UWhSxiw
gIyFa5Hib/pyKlKmEyBacPBw7I/8kPRYz7OM3Zp9qa3MWevlUkN1sVr74NjyO5tF
i4a7nZsYnPIl45OLvSJmslQuBgKcnBrZFE3UyNBI0kJKgmklZikaWnO3IljsMKek
9gaCrYFIM2xxbHoJ4kxfO44S/gm34NWC9ETvpe11osrepOIAmU4cr+t8YdmwobrP
H6KqIK8uNPY2SIDGGVWrmbCJgmiCPB4dJ4I3m6HghdvovJtfgESlaKlAcNEfMeCt
WMpcn6XoR1FpEIXYnyMOeR7oS4nPKnyGSkWqXQATi+MYjgu9z9RZHMKeo3hDHeX5
3Dk3Fe5W8An1nUlWg6pPnFT8cYs42nUDUh1YLAKLaGndFbgsuCz9S2NP1cCqAOoe
LNZ1OMc2qXRVr6euDgOQnCCRBRuzEu2Vg/aIBMuNBxctwyOVm3IoBkcvWl4mOe0c
U/GCtaHY8kc88yL5rsFZxTCQ/fWt/JtUSp4Gb80kY0/RZykofcgS6MDTrpYtyLtJ
jqKhQhouV6fveH8hkV26WnG22Ee5SuBRC2GvkX30++tafi223IOA2JT0xBD0byKW
OtR9UgSrtwPbNQImGSrsM45fLojsQkCNssaVFqFIOoS+gEOdzpD5syN6CXD5jETq
Pi6Ra23zotWSUkVQ81fEUzZC24ftDu9E/yAwKEvkvab98t/7mtucm63gm0KoEu5y
q7JwNCZumaXWJnVvt8t/hi2xIrxNtdLHBZToQR+bMJEjz6Nk3ut/8fWzt0qcPYqi
00ZIlYkHQfLWQcrSFoGMFbEzub4QCyv8CSKfXUwk7zqH2PikooYfgA3Df9Wr3zex
X4yzGOOIeAK2vDtI5Ps8+FEqlkKlDs1A22VdFV4H/c63+eqWXqQHiIgBxov0Yybm
AbyqiLYFrOqHtWp5yz98hNs2OvLk/JvVTAIek96mb05e6vrFPisKgaofBJHiVHPc
EzO1SpTiJ9cvv1Iy3SfCSmmq1YiktpnKJ2bwwkR5lOJWmlcFokNuxSRkV9M37ols
ZLRbmZzk9/Wm/UzpKjQTV+QwsBNFHS0fXaVaweyQ+XXMWKIQq4566QNxg8iyfrGo
0Q4Fo0TO8T54521jAriPUNXUovnkAFyqnC0Y7gGymH1GeaNru41PQ+oHo/6kVeu2
QWyNWXX29WmxwQi6z+jUAzZFc4lOnZSXVoNaD2rfkOm5ZxJnjN30buD19G5QD3NM
XiA2eavf6WMm7MGx/xzAIJpcMvK6fBGlZMYYwzTjFPNoT/a76yiylPkSQNQxR8jl
O9wwu0wJpISl9x6axPb+yoGWRpPnP6APAX5QEazeKr35A+G57pQ6DNRjaOmo7jIv
6Llzyw0dWD8cRW/4vXn/UlLdr1AMak+catR61UtSFhuTASgmMvA69gt7HZA2cG6S
iH5+HX/jdO1iQvgkWDUuN4CDqSxnFn5byHc8MJ3S+6HlxcMFeYdzKPJVJcOnQNAJ
OpR/Td4hobx4odHdyyED8n5ptDexUSJi6o7EPQX/LjPlzgnpBmAfLL4bKtMMD5SF
gciyjohGM0JXIaRwTyO03Bxq4qziP6fV/0bq2xZ7KqdK8SAuFobbRCq/376tWpYo
VLck+qDKeON58tUeWOG4DlM/8GGTNgWr5MYTbxK2Px9yubE0AnKz3/jHhNu3rEs4
fCazt4CvZGiVH8PtoPRBFixypX9aZkth3E6JdjvGK8+5ehaACdOQ+Lns3YFftXxJ
CykrvRzCQ759crLLCui0+Pmrs5QrIWkxpLDnUdRbHAkOwJ8oadJGk8tXWld7QjLP
lsQLIqQ6zVUrzOtINp9WwpR8BbjjLr4unZNxtyIAMzCwPKIoDog0NhGhzeRDXB5O
WTE3yu3TIoMOn/nz5BdT5lIQFLHcuMn8q9OOAxQIF3ajuvNjVjhb3d8nL7sngB0z
uUkSBNioXttaFhjDdAB+n/UQFlbASlIbHnHAjXX3t4bRt9043GB0nxORu3BPtvir
PTHHxbE7b5aOHm55oJrDEB9JzFLokWDtlY60XegxLJ+TAOGu7fjd5bT3Paid+HE+
hKeGxhh03S73MPsYrh2PNL/FubPGPQnk+ee7W5gSj3T4pqM4Tk0S99yjCR7DPwgN
NyeSuHnh2T+kAwu2M/LRaQcIpj280Bswg+WSAfZDYFHS+sZ4EjE5tm8LeaAqSjgt
JSnxuGSBAs6GTYxOTvM4Yr3XxWVlqIJuv1mfGdDztD8ZqMO5c8H3OooqwZygt6Ph
NSrb3jFmjxvP84d6BnYyn79uKfc3sB6l+pz2xunFJuPs/HASQUX0rG5QgFKaLCmm
ME7gVNEM6T+fqRUcvoLKTqsh9yF3bsn1fj3H6gxZAXXttArZGbQ2e17Lg3cAjsv1
/xs3oX95rp5hgSb7OTVLCAdyl0H/ckUvmt4AqkWG1ZTzgRdEeEV6Lem4CUCFfA6G
9SXseJ8bixvDwIFLsmWr4ojirCJwEMyC4S6sJ4TV8UF9eDD6OBbwUSenEG/lZj+d
efav3zeDdEC3TwxHBGyTzX3uBUZ0QpTxH/IiEk0dkXzLTGDoRPTrUjFSlhOJyEfi
0HXghFUN0JFGqr8GhmhRTT8v7xduohYELd+GJN6TCTkFBnvGpfltYPa7Z0FKlFhp
YWNdUlv13puCZ526Bs5lnyv7bADQxuXIEjWuih+OCnnDoChiEk7ftBhDnw38x3x9
JX2hS8LKZbPttES4woW0hXNsuR9Pyg8hz79cxAfehZ2Jd2oNOjNy+UzpQ/vCK+zd
0Y8P79ql6X2QPPWwVIzH7QUHU5H0F09txwkNwPtqFGqh/Px6Q5KIKZOlU7GYw30c
pz3V9gzHpZjVN8Mk99bIeEN39kea1Ao2Z7P1SfiDPGx3m1qm5sMN1O8rGMicY/B5
dodQIzzUL9CCj2YIYtYhfcz0sRwhWDwC9zyUNyvcrAHaarVKn02tY5ztH63dRYdz
YHtBmzPzXtxtcpv5oGGmiXxZ/wGjv/qXVzIylkt8VXcHrgtgvnTBXEkCPa+QBv/G
OOdbOwj1PmtR/xFE+Ao+ih6BoMA7e/KeFBxzXEtRWIAes0u00dOH62sQM6D5Fl8y
3NuHOhomAY8FJLT/WbYrkThoLKlVPdbLVxadAXwrNVvTkIvdsgYSx8BfMuGFTAt3
bB9aXVFlY5ZswdDFlZ+JpSiroKBP9v2mTHss9uYAv632srKxlO2Jnk8O39UoOTY7
Z9aN/sUBqdTqFj/tq+RmdKXHBvyMj4jf+zUEuM1x1xXbRE/r1vIYx6hrFD/Wf6ny
uYKpif3e70HzzdJ5nRgj7siVuQix3y+3RMZkb0owYA4/sTCSRc2n0KCioCVnaZ/m
lGdjjuNAY06OM72RveZd65qFFx4PfFLCNMAHeph2YUFAROXARFdbWdKYlo1xnC4s
hlHeSniBtVZpNgmFkPqTUKgD25ej8kTrFLJaNzbNhzWjQxvOupWY2TsEIBKLaK0F
JaOIVUZfE7w9bnV/gIVpeYzgi/bPSQxE+sjxz//a7t/JFL5lyNH+mLyy5GOwkzhE
R7H8CvdvqioWle6hwWafYQ+cs+ASyAgbLjyq7K51jVWfbbPe23/xYx1ed9stITjw
dCyC3VXfsiloDY0LJAAvhuazsi+FdHsZoWrcQWO/libx/1qvXaoTP3OXVF601QZt
AQM+wfIheaqDa6hzH95T0bTn/r1eO/1+32Fek9urV78Sn1ahZixeFCeWcxfaYxli
KCova9lv0aHIAM633o2HL+O2jiV4dfyA+X2pvdgMJVbFMfaON8CiMROS+Yjb5dsp
qU5c2yIhX+7fgrbPHUp3Br1/nUFzMrqcxCNF+rV0u7x/gsSuw2cRwnwkEUm1YC93
Lf6UsFr3KU+8P3gogG8/1NtgedjAmXZg4N+CXoKpslHV50f2QqJ+U96q3uVOjMGN
JX56Mw+iuGPLG2ZzXRTYvPOMwr2plWjRlkaSu72nk+wRA9WvGI0pTDoYmK0YwV/u
YTNcs8MODgx+Q/LTZu+hHTOyjOuOYt56Xp3aIFaVekur0HpUEB5pHlQ3LHfPqdn0
MmboIaPnJROjb2fI15kCMxA2PZ1VEfNHVNLMM4qXPbdCskqGeGmUWJFf6P1I2j8v
ErtHbqUVeA156Z+ddY94AcQTea9IUebj3qzaXhc7MWbAS7B3SX8+2+O9inZ7hdKq
WLO0Uc7340YGAfdKGYJDsul9mEqEn8qIWW+OJAXxn3jlQMrYVaVaPHm7Ox9z2oDV
VLPuqQy4OZ3ECWWQoyLnTsFPb0XTVTDfo6st/7T359sE+fhZGwpjDuD5lPRJmohl
LXXibXtC+hUBT8dutK/syrAUa/5U3W35P0N+Fm9NUpKdIQDRlmVKvDFIzcHS6fuY
Jb5vmu52pSNXzpHZMbBQNtLdqupWIvmEg2fImOiyRYvPvNIef6sJD0ih9hoL0FEC
59Q9gpOGgNKVLI4eu2DkVBIVSz5ydQjUjOPTElGqHxy4m1ZKGzN8g2AmjY37ZtR4
Q8i0vddG53PBMFVSjuAQDSYE9Bc5RRegTT9vdhdzL9ZacQO+pvu6/Eh8RRkeiXyE
j1QudPl5F0B+4mDiQs0vHHvknm0Wz0lr+1j4HKqWND5yPDv9Tcw6A2bAgZhg6pbb
/6XGqW9UJ0FVKsPOya5Rw7lOtaXsr0bkF0MbO0HyGh3rGen0nbkBhdNaKePzDuPm
nqLecIE2RMVEOilJqg59+eh9r3cf+NBtzQhlzhPaOcJ8osqPioDSLzeQkHDWYA7m
pu0osU1R+ESrB0kNzA019Ngz3V4WryrEDlEgcMBoHlzuaqX2HUGIOZB5eCLc9kp/
KwmbXBV9ykjKty+mW9/kPt/366Cd/o1jsHePOMNSkwI1M/uzLJkHc468eDiIRepE
9/RvzNjWmm4QtbYoO8OdMc/ABJMdp3dav6uuDkEK3AUrj8dwfk8S14rlaoUclZQs
SSyiFOsDZRm9hHijyS7nxrqC6b23YNvvzV0mfpvjM6ECQ2Eed4MLJX31cFZ68Hez
3WvPIEbo0u+FRCc7TcUohg0F6419GrgdGZA2KUnGVPgyRtOzE3xzbqgTPys69Tt9
yOVqTdmH7AUuNaIN4ir5IPvsZwAAUSrpzIfglRYfCWTC1XRg8czz0BAZrdhWZqrm
mSiX0oW5s/8sN3bF1kEh+QmzBf9N/H0/A7ViFBzJ34f46ywTIFZQqvb/HnUtWpxb
wIwl9gPwwKRQQPUqsECiUqEO5D3VR9IwJTAUay0pxTVv6OFKH5pDsnxkS0P7furj
sSMI+AM6NidXxc7PdJ0HsBSkvYFGfuXyJiB7SYYojOlQpLL+IS88b9pCim8Bx+0V
lDos7X2EQ69PVyqXlYuWc5FWwZ1ODDeYPGyv+3RjUT23VIdcb6oSczufok7XHRpW
wCRoznQVVM6yTCv4YUTxDthPGpT+XksscC0C3HT9XemjaOaw5HrhooDXhdDeFjYr
ZroQzmKbe5LsXqgXsE5ayUzFtuLXfXwIsrfUTYt9jWocL9H2DxHJbd0t5bmURh1F
ahz1FHIFehtJ+BJEhqpTtuzfkMYQkRF0rmDgLraWjDeVR/UEGsmmPG2JKDT+NUjw
VXequuMZDhAmxN8hwyyDWJJq2h1ULcfQqhzlM73B7D+PhqSyijk95GOswIpO+lQX
YYUcAr4Fab7ue5EFfzBohH3te1GH9aju0plOz2Ep+0bm/5pTCcx8hIwyG4lEoFxs
RgDE45f3BWKdphOpT7go9obfYYkJL3rH8jXhr9MN7cCi1U1YYIpQGVyz9z+toSE6
GrSrFSvJz0eOPQ8UQL4DXO7juPYb3m//nm9nQGSNvyvGQagF7qa8XAYVawJdxsyz
Yc4g+lsDoQgN3MB6TOxh7qYObnOWei/cc+UivHdP834XDc2hUI7td4SONi3GL7GS
BUq+mXJF8VlQ7uPV90QZTF6BdzfdwZ0ppttOJdpZtIYrGBgU9/rOgdM3K7bNeHeq
pDCs0YFtQmNcn0Ouuo3Q9wr9Jkg0ovK+Cg6FeDytKqU5RcCRzK99T2JnpoY7utwg
6kLjOnKVsysSvEwjp+XJzZ2PM3HHfT3SV0H6IGcmKSyZOTKnXK4ZVl6pkk6sb8fw
G584icp15S4+8CN8nUMPrQFc9+qsF4L3oHvIFIsR0DYoVsZUTd7tsPlp1KENmcFp
+O+CiuYlD2l0QzeYPVff9EbrKy070eenhJltSEOyFHw2FRZsowgtJlSweKjmbAwh
AtuWq0Law2+s0qXtmji9VetIccgxojuPOvzCDAlqG1kIy8ilVOqL2RraI61Q5jpL
X1aWJwHMUVVQSwTKL11ju/yVbUf8cYr761L0M1oS/Fz8sP+A8zfse0BaV6dRXmzu
WUSv0nYXn+SL+0pPA/9d8hkOoRJl24bauCePCrRUh2ipxJzkIt2CFsu6d+jn3zD0
OJ1VYCsHJbFfcCpIPvZsdrSSpOTw7qzRyy84s6jzjeycL0ES//rG2Z3cLEyx/Gdm
01BVrRd8wR9r0LV+BcEY4Ai2O0OHimAeyQZn7P+E0/6ueSTtiavFqv8GCg8H7sMl
A/BD2AgyRnm1eyEmtMz1z3Qmo4TLpdlP0ruT/5CEQlX9q4mYK3BorD9vz0Qdxf0f
O9a7sIQGkoE5QiQFx29LpxOU6PhYpqr9Cj/BE6UCFkuetcIG7J9k/87pBpIBghV+
OYcWP/RI7c9DXomIJgyc0e7t3TX1xaIYfuRjvjil5ZGs5Yj6zlkf3pnV2Jcr3xeF
btKkYBJXu63q9ser2NvfecRIl16lGcoFRZyV3Efh4hRLojHby88jzLVcmXswXda9
YIYoAjhyWzM1CgLRfqCqmxYXP9hW98oRR22/SOxoGDYcm8NV0U/qCc8XQG2LpRW8
eOWzJEY0tXhXSzl5B7lSqTZFCjIohBbZClZ5iUZqyuS7LzIb358Y9zX8fbuF0Zut
SFYdQXq6MDYMJIpiREfiVJ+geUBRcybtolM3pNweyQcDEC1hmEweC2YLvFaie0Mn
rz1Pr8EAPTNxCHypYdfax6sBjbSHBHZK+ZqQ5rZgLfEL1yLQsFHxwuENwohzxs0C
PabDjnF0cA5FUTIMYmxeb7Aly5wPXeaO9XBYQXBSZWZI/RJpA/+J/B5/tGWUO47S
Z3NvHbL8i4ziV5/fzVlPQMGnJxJ45eTDmh1AexiR1Vo1LfdVMGELB59yiR3kC+yA
36j1nAV2UOllihGGH4BegOYKoaaeIznO4smltrCEiU4WZFQ0giiuz9cVYzsByvmh
ll9sHwLIeX3Gvg4A9MYS4ltPPhu3ZNEbXfm4F9xqIlSsgw9ssEYXZx2ZR6WeKZxo
XwsIjnV5W+jrqNC22PQAoCfAk76/+cUqjwNpWUcepMeE1524K7F/nYCUXNX2Jt3S
1WKBr3jIutsEuNs0QCixxEeGvqzMcd8sLMkxGasxujSW29+0HJupuQ3u9KKkF24l
NwKVivqWD7PK35yW8OrNHWkoNmdTkyPvhC9JfgbSxE6N4QtC6J0fO3ss8jJ2IIPF
3dczK5o3fAMhxp9R3TXnEbMQda4BMv7q73Y19xtRCyJhWSUaW6s0aCEkpbamr/oI
zh2yr0kQQrkOtpwgAdWhUbELiNQAEZOaeYvhc104XFq/N9LQNBuwxXhdWkrf9x7R
OR07X7ALIn5dF3pH0R1UxfroSldmpleWBK5R+l24oFY2Js2pNrkhdD2MthyyRQMg
K1DztwZ3TdDaPWMoHFgwCOrRzBHnl7NmMYu/G0YcxSilds4osJsPGiUFxE8e6Im0
1ZjNfLWTavrtJOFEcUujTB5p09pzRy9UCiqsHaLRQwycbZ9XFnMbmtgs4jCpAVl+
Qaws6nsosD3tYI7PDR/Uut1imMq5wJJlOmIXXFB/bJK/HsKnXYVbNuZ4lrWKD4LP
u7wbkI+/tNjF0+rLaP+erKhH4PBrJ60j2uWskGUF1Ie2N35GXBt9rkAz1VnyO2yE
+17NjGAxKty8Y4S4LgtLF3cm9aySVyCPF2g/AelGbGUuIYkV2RP6z7nfbqkR3GAv
zUM3AO0u9paeID8jPgNAg9hoP7P6qSx+ANbJFlDejJ/UEU3aehN9E62oon8eSdCJ
UwhWkDZ0/vR8SZFeOEy3ukycfyr3sCzj/Sk+rSQo83QcWFjc9Nh5OMXMVq4XWrOJ
zvuEIgPyZiiU2obAKByVx7fWzzAs63w13cOD3kirjlzuu42XFwbArbp3ZPQguXp9
eQhPwjwEI65L6vAMTwpJfPxBDqFF0WdsvAU0Xkw3r0BomYzSmhYI9phRgq7rGyh9
lsCzHE4glXekUElsG9+8vA4JwuWo48ix9C5ShF0QZs02hghN7rpztpfbqCk429P6
Jt1pV0ObIxWRG69t35T3Q4ZQjqK/rGn/dlfDk1KAFFldIK2RJGAQzZyGMvHlfHND
V7m1rSjP0sWrOgXW9Mqi4xijELeZ/B9jgvF2ux1ZXwNgXS/HI0uoEfGYpqsOgzo7
513ep/MGkQAvt6fBRRG95s4bcWdv/8uj2GxGEmI8ram2U8bMHzFdbdkqopnJiGKV
hht574o9lXv67lhUIQCy9LsRXouLQloxsCw0g+pCJBX7a6UX5uce2ea9Y/R7FZ9a
PCwjUGXQ1FkafaCkcoXb1CsQdpDBuWJaLBR1REiLu3YqUfxppwVmWIJlXx/UUBFc
q/WompUHUX5DOE8NHLvBt8lIMhL6aUoS6X99mqxIu+m1aUB8vV1mJ5BqYP/vy7zq
SojDYij+dC83bVEWwsMY355vrZVaVBWSE5Glyfek/Pnrq9zzn5lehOszIvTUhL1R
4+HwkP/PwKbkKWSkhFwdeJRujbtDEQPZZmCaVAZ7GHD2RGazNl6sF+Dixj+73XKu
bWH0z34FLfqmXskw1bHj+B4gSrQrEwbhk9zrdrOpVOHABYYLuTSegyqcJP/oAs0z
YWtDHO29mV9wQAX87+wRIVH3tt/GLeC9uC9QSqivIY5+NfHy3asY2rhGflLtdMgb
PPz2lQOvlhv2TxzxxL/BiYNF1lIxugt76LHW2B57DV1oCILH4M0G67+q/Gtst/tr
qwJ6oQinwZXbDK5MFGfhRFoy/JYGA1K8hnfwm3t1Wqh470FTg+qGSNsmz1xB9QPi
9iOacltRgXN0jslKdmGJtWNYMhL60i7CjbP3wVoudIBtzDAzuCkKPuMvEZYcOMys
hLHrd2XOS8i37ibn9/TasCGZYcCIcNVe14VIgdPUC39FBNYcYQvbyb0Lkm+/zLmx
PXSCmv11FBXRKI+y6ZPx29zA3s/3m+fXr7Q10UdS0LtsSt+z8ey4IVMsoix4qwra
Aomw4xV4yS9/Bb4X9NATd+7IOezQsjPvqA2Ofg+bL6HX7X0AI9l6jlUnO4k2/3iW
hzzzj6g0pw5XG7RPRNvcZ3BP2q61q0PWrTUOBFs4KaarI1475NS948/NelqzhDhU
vu3fwD49dX3bEWhhZeuYnmhW7zNCgf9ggeRB3ch+BRPxytl/RVTS3b920OcRR7k/
N4Y3TmNsOOYYxXMT0kcuWaBwhk5B3MjlE8rA654MeEWi+tRq1JaVVD8LcvpGGRmD
4Q+B+TU5riiyUVeaecmeWE3EZxwebOZ3Q5d7pMBpQXN29k/HAtlgm8B/M56NDiLD
nKi/tKXd2q7ftRAiaghNfaYRtjy+oUgpF+F/BjbzMoBAiUZqMajoOY7uBJCi7eNa
yZj6p2vrJuxBks65VlBJH4QrYTxhjLoLbQtqbV/CiW6L2T4JZ/ks9nkAVrV3FPir
0ldLubDBCJaUtioDvv2t1a9hWTyGUhbZZsgrDQXuUlb672hNs4fU3uPenwL+0cAV
cAkYXDrlnW0FOhRw/60LG+F2QTZuvRKHQyms0lu4x6gQKAC6bVgnxpzuK/tT2CN9
uFoVibzfzo/oXX3WDoB2Ex6UL8RhnwXvojclfRHtR/PUZXOAIh8aDW6q/qv+Apxt
JtRW/4pF8N/0bTjK6FzH2mIPFSUlj4Pn5nzQG4GvMfmGiG5eg9DuLdnNK84jfJnu
GUG9Spa7kQxJeArH23ku8cIxCt1AQcvrIzSn30yoa42XUg72zbfGrHrthiZd2ODN
O5lQYC2ISxfJBlJ6Gn4/V6S61OL8q9SDEOAHLYH7fe8ZdwyIJYnTjw+7zswoDsbm
gDIXwjG2HDnl5amELVasAaLtZEupSFXvWYN8hG0kceG0/2eO/8nWkjyroD4uKLKD
ttsGOxEct3WXt01+M2wu19303nsc8f4yjTZjdDHeDw2+8w6XJTf7S0N5H7iaxyEs
reiYbRoxHTJX/W2NEc/HmAwRxmsH5IQgkyroHO85oGsNaO6v/TRSDHZQWg8uRaPH
Tp9kW5Tt4fPZZa6H5oh58dWF2Fg/8CtIJbetmEwEo56t1x+GTsNaeyVk2S7BdRJd
yw+Awpoq69jaC27YdwXpR6cmtcLOZ1M5EghQPRjjEewQr8saqY9BT2gjvEpq4kn0
YUNKtla6GykMLFVJCHjGZlS3o7XP2C2oMt0KPdHnpgnxWMVzkgyEiy4W0aiCVrvt
R533gd3eprE/7YZ5CEiLXT3SQv3FCKGKrfnbewwqXj3IHX+CBmPnWgyyZLLyh+XQ
u7lK0M77AFlLKrpPloX8Z7e6lUvnGSxAQ4yeTj8L9OcmrCQUuv6+Zru3iGott4LI
UwH7Ea9voVz0XKWGKqzUcSAlPulGyN2kB7lMX/cRKOMMwdlLd+lfjE9ODrqCie+R
lnxymDe3QXChaugkXfc9PUvUuDo10/RaObI+sBfhqJEpLCXK5eA6lWDEnssPI7Gi
C/QWObtT+nrPPgrom+0vG6HA8QXqiSxw7HbqoTCeHnM77xOrqwadp0ecw2WOgeJD
3CLA/MM1kUXaK+QEdjsrIZyCTIW4gwLGzdTfC8cGwwl1k1rBSv03oZYNkf/nZ0lU
82tyo4Nchmk1hoKl+MWQ+AQwgOSa2AHQ/MM31jj2pprJ5K5t43EIZhyZa4G3vQiO
j2OlSmQyYiW0kCrIl7u/v3TgHWmApZp7zciGfZb4iSKWn/Uo5XWUho97jrr88d7m
6C9Mz3VF59i92Qi8vRAzclcHHOzlmnkMuKDSbUTaifn5/eulgVlSWmnrPGsp9SbZ
IWvES2zh8zfD5sbAmrOGUaDRQmANsRn5CYFJ4LDdqIV483SxARogGR2R3aztd/JG
SXzr9ol7tpWFZf8GTnM+CRlIK2EAYwRFTlDpAVKf4u5GnxqIdcxoH+gntvgMpUb0
O6DPDXRmbPysQRskETnX6smhxy5IofnQGUMCPFLKJ1dY+IlxMSA2ajsludO6vMEL
4EhnAuxEtYbfQplCufNDWYTXPvRycjLCqBDAKwm2IF7VlA+Q65vwvfIgxnwKzkIU
7+7VnltXxRfdgyTI8RQ3BNReeKB2g5KfGASeqgqWIwewdasLo9lR8Yl4SxgHI9w6
vFWbhwFX+26BJMAKFtum9sWlJRoTAsDb1WCjgTN3cjvKqeyWrHGh4bdUVFnwHKKj
R3Y+83lZvANuO+GFDiIbCYbAN5wEZIQSoRoNxsVSJN2L3Pr9OM7beFO0sSIz45S9
rltrsF9rLlqTH5xjBBw8xyYDTYjPC4u1t/AlJYPLzkoXVk2gLaui9TrBL1ZwiybK
bY+6q3Zg7pG1T+cx8wjkmi+PNVZRIJktl0zKMJ9/VPVbdi+lHpKMuST2+u3C8qVd
oE4ypDGvkcLFgNjh/JenQg8QOv7CzCp3xy3AW8gjjq7TgZDPGkxQDBhotJqGubQr
95QgfmGK2cJL1wVQ1KJjqV7zZW1bjbUaIArOsV8gX85sIz2oKWSbecezwhEIC6SL
uz5eC4hmoG21nYj9uaco6UZ1/vL/k5nxzExhxZZyE76unrzaZfvrlKmD6vbUXubU
orSyBea2CI7q45Y9N/VYmY6R2Nunuw0Z5wf44xIB+cJoyOWMngBI70Zf9hG2i9xk
ivbgeZMQHI8oajZdFoF9GePYae8+U+ViMKYYpkuMukOk9VQ1a2YsulgCc9jn21hf
st+tAHBG5p0F8e5UxMBgt9uyATflEkNcpzlsNOXbHKhxaNLDAnq/mhwAgvaJt08d
dKX89Hg6bs1Cf4xjH9VueX96VI1oczyvf85TALRB+AbDOfdKTQQUnNLva9M5sMsE
X3oAoZbJuHvsUItsswTodcaa7KzsOE9Wj+u3PaTiT6dblYqbwtLR+H2Guops7++6
JIFIKfaib7323CKgL+524saLo/owmYuXnumxovNCmnxpnKeUfU6Aqhsjo8BM3ci5
uTYHUQPSviTEdzWDs/rwBELefEzhd2jWbSFhHE/qC+03AP2oB89KNSZcPKnbmyuR
g94HTxvkLuscaKuSDSIU+f8xCctBZDjA1u85a38Hna8ek00N/Gfv86eN0tumo/pZ
PJifNv9HX2lgd+ASMo7UWmCyXhqjR1aLyoUNC3reZGFJC14Dc+AsFed2xlE3/ejZ
2FV7bf0ZNdHUer4Ho8oUtFiTDVAKPf3KBbcPXKMRypYVbEZsr+nEsJYGbf84og0A
wEorGhhwbmTheX0XHjbOXvj/76oLAmUn9fBl25bDdPDdJ6IXB3wwqTb1gCjAgTQT
u0uoxK4hSJTm3tiHr3DwH7HdCXHvCmUehwgkHcQVWHTBvMqufMl2W1+lNWIjp/j/
3o/h6kIrWrvIXzdtAEunK5xd6K5YV0mq9KO5Nrzu18D+TZfaaHU1ugyxehuD8eq4
hqDltwYQ2OQbtO7hGBMv4pco+v4KlBzeTLEO7VS/X3pEHT8PwpGgb4QNt0CcBAcW
bTG1RkPc1GX4b2eSoAZbLhZAZsmARAb5n6tbPfqeatXYfkvdojVPVJBsZJ2MatkF
uaItt3vEZbN89WkitERvNeCgkXRq1dXVkDGsfuJw9FcOj3a2swg+CgZvCQzb+lNl
JJTTXiKCIUe+M/qnUjgqSFtUinIKzzhNL1ry72KmiNNkCk+njbeiP0HKxPkiCK6m
YiZyaH8G6Ox94SK45u/t/RN3hAFC/HkoNjkAV5MN7h3i28NIzz+FzLj6OiZwAKwJ
1YRebMGDQUN8FVYrIIK+A5JN1q90qP20rxWimJF0z1j3Ex1P5nASmcdztZz9nQBf
UaFD76xeJRf821Ax9wcL6IqGCpecAF0JniqReswI3N0Dw5zE5tN4ge32CYjYkbUx
DZxnnJ4t9Kcg1cxxaHo4ppCA+g4zBMlk2D2ICZv8CfGDlrSoVoYDM2jNxdo6466T
cmbNcL1j62nyzV0aMoif/FafoENDDQoxyX9Rmds4v38K8wef05VK42t04VBvOhTi
W2rWqOG9zYabSDMop7433Qv5GH1Ca7vo7vDCQeIRBSV4POMroulWn8peyej5l5+t
K06podaUtvpBKjvdYQLLUfv6yL0Ad1pCbNbJoos+h8ntSvtYDlwLRVRk88gLuB4U
3mTbg/T+ZA0hPL2P8Aj/cLeltTzKpRXyQeu4dPHtvNO5VfNF6/1AEiXRawSyjYiF
+WR9XNqNl4siB8AtPO9tYj8cpOtKPAVMBVyEohmhqFmPjZfy33HFBWVRnWWbrBk4
I8voT23MJ8xhatr9+PPwf4M2jidM77Xebwarhylw/E9bwpiP9OB5b/a10wa19OYG
vxEpbgaPaOUoax+bgUM0lIPEvKaCk04uKCkB+ac52I3AZGyx2+qcDIZJUzLi+IFi
4ZcESSWiHB2TqMZmgoavSDUO2CkI7avK5pfbkFjOwouO0jXMJTWzsrJHVIRnnahL
jEDf9reWfg7Qh3ePvMT9Y0AUSTx3dbETUp8uOF4yuqauk8VDk6v4UE+Qk+B3/lTI
sneFEBrZTRyIb8IRvHEXMuHU4xbl6oEEq2hmIroZWv35KxqJK+iS5swoDG/wALmj
CIX1MDXgJMplLQjY5emKNPBaUTNdODsxgs+vzQn++gcB4YrCopV7BvrUUsRnOugl
mjXuZU/1D991mRTblI97Qp4Hrtb/eXd9JcVJ4M0y9ZCVqcZKXZ1+LeC3Pwb+hPEU
L1IulX0ag/3sprrx9nook8eZN0t87z/Ahyegq4aNhvehvfmFHKF0Ka9yaCQ5o/qz
or2g0jtmjVO+6rOjGoslXzssoIj0K4vPkZfWsccfOpMEml0x1+H8Eb3U+F3O3UvF
JLe1xc90YqHYBIgqIvUceZSfrCrL9m4tObDzhKu2vgjB6Q+lC7Zdera6h4jcEyj+
OWU0BQjn69UfENDXcfg0yj8By1dueQf1pdJ+hH2/c5oi6yRUt+xTQhy04WUuehlm
oEotMpWbPlYnbSVMhAoyQYcq+g0Iic19NpBnqNW8h7vhcY+MHoUJysOU8+x4HP6Q
9IHnwuWb0MwCu7v2x3AGl6uRevMV5JNA8JeTlyxM7ThuaBXVmKs4mCYDBuYWNHMb
eSF0SQ2p9xtXArf+lQkhkhDiAon291A+e+10ybD5ZnhGBKAHrFtI9WH5dJ5wcP4c
NveARSbwuLTO0cHTPAK1DWZoh6LaasjP46Xfq9SEKxUeqpFtd0SsTwjVGSxc2d8M
7QFHM2J/3ItPqDR6qPw1FcOlGQC8qEUNQ7qMqqw9eM59Rx8bSA4+wk0RVV472pmX
W6rxLAF7/oXyplLnsG/vhvcyq2pbuu3expuYI5+/n5ltbQ+aODjwLi9aQc0l+nGk
n7O+hD3NxHQcFg350aREdKTjzbpaCG6vTkcYl3pgsBLgjes9VjQw1pNxnwj/Jblf
mddFsmyZLW8NOiaZjgrW6wcdlPs4SlwwdeCMuHqaIS5SNLtLnqQS46c1yEL1iXJq
q13wHDOTzmYDbbwWNeBpj2qRPV5rlCXU2fGNJqqZKAzQ4ZFMTfVIVFiBO5c/i3GD
UG2oRkaPyWe1SmYJ+273u4b4eTCr3lzR2oGenyjaVI7CBOttFyo7AfS2a0w13COM
L7kRzHGv0PqEV5E3DAO5qiIRdofTyW8RFq/QGMOnOuQhNPuk3Kr5IsiXZdqwXT3+
lj3gQuikl6suKH8wvws+Wu++EcAJzE09q/NPvB6NKQbsG+Q2POxTwEewkxYP/syd
rBrokHAsOt1dTeLSX6HI8Y3zn1gN/Vgu0kUAc3PcTK79Jf63NIjA7XXx/r47oIZc
mnRyWXgo+yljkm4nRkeyPgGooOd5021iU2HQ/gpjhd/vQqOG2saynBgv9bbIxD5z
+ug22Cal39HnKGcxKsw5fHS/AGTAGRJC8rBvfzRZvpMDNYIT166aSk4s1ykTBN4V
PtdvxZLrgkQ6hBkWfOOD3nds+doLSXGwmTJrlhiPP5L1u49tfP3ut4QuT6+NsNSB
Nwqy3kXHul1IZGP1bV8I/p8E/luEonc1JgeuQxQWOltnrpKvJG+Qs2rChfUFwx4R
jXWOYBHGVK8A+itGDXOOTCuLuUDvoXXdHIM7c8vOOKH26eq/3Ez9VJFGLQhWB9q7
eciJOtLts5gxaYcrpOr20I1BcoRoxyiYdOJDEzAOfDTrrMus6Az21m8FKhhIpcp2
lNYLgQXGALzOYmS9cpZCDvqriEkIrjb52tnpxVc8csMQIbsSVOPiP8lGYZxzx6kv
P8rrW/iXvdbWCftg9Ko/Fj7v1fcgOZiE4LM+xlLJ2Mp/9qIJD9W9K4d7jbia8sPW
w6+62CsExl6WG2RGvI/MkNdCSpN1gyKZhU9SUGUv1LAIEp5jvgUpNV16gfvVsOUT
jfDyjjkhyl0xWmHFpuBbAJkUYCViJn/FjujgwqNFnc8kVQN5u6R/v50hGiRpK/hF
z5nqZmLeCVRNaQiWYcdOqk8eoPHDnNwRzm2QMHAsQBqdHFnyPaL15euANJ+x8xQR
DAMeL3nwHv6srsf1NRRmUSyqUZSDmxkFMFQCQWylQPvqvoh2OioWfsoknp3UFRxW
YFpu1mYwe+exyniS69Zbufmqv56GWRUSi2n48u3fMaYQGwCQfFKpurLCVz65G5pM
BoEjSL2+OH171AwH5vCieIjt4vZXZyhNNwfKYGKWwsawaC/FHXSvg/6AHXZNpjme
UYt+qfM6S04hZ61XZabJGhnN95ic3ESkvjTDoDgxbJfdT2smBV8oyj1oSM5UR7RL
2wWqeEQlD722nCWlp7CwA6znJaDkyZwGYRCthx4yiYUNc2phfFq2EoRZfGKn/BzE
mIT84pHtFoYHxlfl10sV22Bb3XHAmvyjRYQQfoZv2qfH4xupAm7WcACxfy7RYdZW
H+Ikn27HsBTPGhCdFNOnUvpqAF12Rt2QM9BoDUz1lJPk8MHwTULRbDMtqRv0D02o
oKXlbNzUahmcbnnDTz32HnQ69hhUZXCuoqBh3W08k02nO8wyaZf3C0D4pZ5NpaYo
Rb8sT/g13vJd3ouI10E+KTbmBkcQBoJsHJGF4ZzVrIzzugvlonpGKBxZlS2ClhPk
pP0fwVCBm79GNcuRfTw7rYKafzu3jy7C1eJVS+i5/EXBuMfNa1LhWYEKKjWeTkVG
49Vtga5juxElpYrMw26j8Zy6adaAALDtUz2WcnbGlm0olGauzJQKDfGnlIqXrzIi
YIhmpl3R4ZrUc3GK+Q1rzLC+mTxUBetkWcTP3lJ1RdMOOz9h3SsBSE7wivDIvBTH
w27+K7J88zo3RAROBxdwfQMnV+fZmDw6dzrLwd535Cn08D7ewv+0Obrb9kwL0LNP
Q3TUZdAQW8FghuUInwQ54Zvxy4ntJYNtSFJ81a5B8F9jC4S2LEr2XVpzbyO/tDe1
laqw4nTqrIH/i4oHFvgMDp379PS/sjR8k+nnTIPsj7giAE5dtLa1gS6Yw2mwI235
jRLxq0pEq9xBGjoeU/gDg7wGGOfrRYxfdgQZFGhU83y0O+nP9qRtjobvM/a6Lrvw
PEUIxfY98E1eCtrjl7Ua7qw/RMD3JmqRjrhBdvZhatY5mE8p/8rty4GkqgMsvhxh
lGjdAGM5LJbNV5Hlb3Jzrn4+vMrET/4muT6srm7o6+SnEyLr0L9ZakcBoqJVAqoa
jo+4qhYKlsQ4bClEw4q3xOkIyrstML/ZcbPwmW27jOow34ioBuyGEw7m5ITzf9uu
ZkTjwT3uaREJULGwQysi6JEUoV0dNjaJ3x135MJCy3utIcfsc+GyURDaBVmqJcD4
CjLv4SDDgIiQq+MoSIoBr9Ccn/gBWs2YLWewl6SCY+wqmIaZmIPNGfxfmSiXIFcb
LuO0LMla5jKAtYHqKmSPQ5yyojpu1KRqjDeRMSGyIZ1SyQGCMfv16i5ithAEAHsT
nsr0i3cA7SxTxYXwBOf+bjNTJxEl4G8yqhgLU8nQggR20QO68Chu0sTVlNSmE49p
1hisrlcH7wQRKqLsGMMfJFvCQgc39yxdSe/b1hE0GOtgkShjYtM5WrcE4Rf7ST+y
+dTkhqsJVgJ33taEmaHhl7qE+FMKY8P3hT2aCJK4ymOf+z/CH8PgJ/gVUkxGpZWS
qhkkjbcRiSa5JyD/tam7UXT5AU336hiXF0AA5e8K+7IsYmFt6bPYY/72zA/CUC7+
MGg5VPXFElziOmbtOZOjTIvE7XeAYwwU/VBg5tex/IC0502p4AIOti5ztZuJHlyC
bS4EuYul6skVv0+9Q6hlkqg8MvKlYG0+Jr3cJqB32OW6WvaM0erOH+t1lv1PQAzn
jkmEj1vHqpb4GFcg1AeWg9/fPnUCZgapoFsnQ+xMbv6BIrvWPW0w7MJZiXESMHhr
kcDkyGgT31s7lq49JtgTmxroSjKCag5oGTplWYx1IRsG4c4QKrQH66TPVSjhwaO4
MsC5HekPdGLXWfOHmf9qAYWLlWfpz9MIgPFRlmabHqnlG+eZa51WpstFAuJ+5bjN
SyA2OEhCDD6qXgel2BNGVxH2atMM+enrQynhfAAsw2m+r3iWq+p7iTTIYEAWBgJC
YNjwYKbA6Toby7neaB6kPcdW/YAotfzY01WObk5A4SLWUoYldhM4v26YO/ZEByzC
HaxjujbDkJDQ1XhFNBZ8jYeBsTZb+m4K9qdrioQnU2eELmfpCkkILoU6mQUgXCqa
BaOg9k7NFr25MDVzAP9InSw175pg5Vc1jZYD007b3zeTSod/EG6aXMt3ukkBDLAr
O/Tp9XSezcbyDzHeSEWT1haq+05zODwa7Ggq5K+YZAkhmr938iheDeUQJwQtueDM
ayYQhqn1rXi1vpi6EOzsHKQZPCFEP7qfleTCpXp8IR5z4FaLbvpLJ1PD7/aV8Mbh
IrG9JFVz+c4Tj3K7/cNdPNtCNkivcM2z0aUtD0Ur2ZuV8AQT+QLoWcm31JMhcW0/
+MG1181RiOYjNG+6BgeXa1CSExjkBjE8KCEwjxNvnhJgYFZ1D/KHwKwHGUm23Gfq
u1FVvXw9wjyBZ+wHhy5SByM/Nf22C4DLL/Y5NsXWjacbLbqqJa7W+m1TIuLAqW0a
gw8fR60BRpJkuYSEzCBeEIG4Sb0/8If7yNaZYeR9eKLqD4kxgEhqBnjx2xNBFdjr
jWeCUe12sr+quXJ1J2/ScMKb3tq3nBBJbRLzbw0CFlhH2oDub+dHSxL7pLKNOb7M
2xWwnIj9LqRWuhxd8NQS+i2ktE/URg8V6g8vfQ9ydCcF5YfUczn/j8l6aJxoqOi9
3qS8URlD8vN6oJzn4WvmxnixLmofm6q31n+9Iu+kz5IAUrbpJOnn338aZcAnoiKE
0ElpWs4dokCcyiwfYnm71gpqZVe9CI62ZXFjh9moXYuJIxqiUujN9I2dWd3B7CAs
/ILhqie+68SNIcNIQ4+DTYtrnYBOJcR7EBrVwxVq5AhRprOJTDgvgVd6O0T60g71
UvxgE7Unl8yBpCk8eqNipnzbxRGWRpX8zONW2i6ZvE8UWIx6PdJHhFGfcuKbbnS8
EwNPCwEmkK980ANs1ONzsUEOz6lPattLuaTNG8cIMAeqBuQ7G1WpBFoIBhdvEy+v
suqtLVrOIdpq8Ibi7qCPplYrdE/oiCAleBolwKu/T67FEQrPb39lFAThg7jwdIQS
bwkgIzdreGhQrsOmvc+9xCEtrytZh47T5Cbh8ueniQuQbw011VUtTG52mibFIlSl
PcW7NG0p7V4aghcN+Q06whzll+aB9UmEnQxGv22hu4NtnCV8+fxWQaq1edjVrDsD
uXum4OltTdNBmsCk41y/PvlFxy+lzB/RTqu60bgzhgqIXzkjAAY9vR3guKzcYj3j
Y30bV2MWn5eOv6e9tpQO2B7u0DD37Eima3nN0NofDPbjQ0n8GzgpNrt1W5rr6Fdi
axJNR++Kv3GsKaoYwoAFCBY1bY4lOFuQXCmZctapKXpE+zzTPXW17zFKpI9W4FyR
7f30Y2dDeHJBKyvqJUu06FzZRHfHvlk3CFCLdmxedFZbEJ1Rfkls/l7MeM1aKiRE
0hMDghvQZY1dWA0A2VIRFLSoJkPeADDlJP/w+RQRdi0d+45IskgCvTTY4Lu+QOVk
okgSjSWl2Ldh9sMBNGWL1lt+LDTbgEKP5R9U9VgijZ68Aty2m+p1vnn/hJqZBH4P
DCOQ10Ww8o5XEuZ1T/jx5RqmmWlUnO2wTjDI3+0QJLHJZSb+M+6vrcAJY04MnnW2
wGeuC+DauwUSeqbFkUgVi4myUalJferqeCv/toJOMQZ6JzsrPlKXBsM/SQofU05M
NCiZ9pnhdxif3g1/iyQ1vREcdEtgfYoYa4s2VM30eSCO/IArww0lpCzaOpOvtuYT
8RJqJGJiNgP0fJ61agMWQiywLV3qM3jD5prdCXKgTbevTNKXtAMJCuPZrnTD/RWD
sVUaJULDXQ0E4rxDAxVRZfR5L6iPgyUwO/OwKFJ7c+E+bYaPs3vGzvTFW+bjbuyx
ak+0y0QrHmUQQ7V7wuN02fvXhDpxFVquuRWnQ6rp/1Ep1atf2RsqvGqbBjrPqxni
d0YLmrXQJTpRiEeAMkX7HiX2NYqTPQuXMFkUzwO0500nysJ+rwobXhqe6u+vEP1q
rFzyph7CVCHp/RV/3zAjRHUSSF5cAprkNMuv2t+m1qh7nltW9EYRCJVUosrCJYX5
26MUY9JZ1ahko2Je2JGqizcc1eerP2O1kT/UPTICEBWNuwjE7CDsDOm0tleLjcFB
5VSK9E2VDZ0h6yAPu8ZzuY+MYfPJdlb3NQWG5swmW+/VcYBGQhRwx+CStq7kkc0X
DvhLcNJ3LrtXLMeIYeSOilvb2Xm1GztEx6cma0M5j1ZSf3oa1jtc3dtFHrhHY9YE
miJZ/wNUAo3fiazObabFwiFJqVZFng+Mj3R7VBYULhkxX2Oe0wzdul8Pniipbyov
UtgBQIYYrZufPRUvnYvJlPKFq81LspCQD31qTb37T1zn44tWweaz/2raX9g4GgEt
8hYk/H6xIxPROVuz/9npzImMCrXTW/QvSrIvbiWm6Jzp9zLEo7BTmAQTCAnk30Tb
3dePdWttZZyRjoBsisBTDSuTwLBRDhnbKtat6uN/vPQa7N/zxmDYqRtvatmnLEM4
9AKhUFteJelWovwabDxjwDVbSJUBeKUQddXjEkElU2C/O9Gq1OuOvcE4vA9KMDyW
YLcaYli3QlSkfGlTM15WJ49BxM83fnjte6WzLuoKMa6BZlxm0huAmks7usd9dSph
qQhq/BcaeGdOYMjPQrdeXqX/KlSrdOU5WMB25TqYp7MZZGr8TNCXxAUe8b/z7SD8
lDjIMXxSLI1dYVbioGhTuZegtzZRYSvpet+UPi+o29JoU1VoOKIlyMo3PvS3I71P
D103WKFWE5sOKZcnYJRKxLry4gIiWSmDSsmpGST+aeZQhkjPYZNCyyRJYK3pkPJv
VGrCio6uXb4AxG4wZPGToJT/ePAC47fSNNptzdCrS8s1MZ12BYREtXxfyBT6lsfU
ndEgOx8ro7w5E8ccCP6symKZV4sHFjdPFSR13Mk/uWbMeUaoa9I0aly7lcx+E1bu
PlCOjWM+zDW/lPF7w1sGLaaHDdJr44RGRN/FXdDD6g28bLlLxSKuCb+yq669XWh4
mEf1pnjsCSOTniquI+TQuwfHue9sliSq+pSW/a8/o35LKhkDkAi6ssxDfa7mloZU
NmzewceqrOEpm21izF9ued0sNUhUFKlY79IFyLnlypLRPkjUtynlMnJRPkRlTsio
o9w4Lxe2Qn+4Rxh04QY+Uqj0Jj/CFJuQlbSZcXiR2U8lFOAqQfDm1+nUQQ95A8DT
D7eWO4mer4WRcEpyvk1eSx+tMwZbL1xlxEB0kqWWwy81tANaY/JWXnUnWTUB3ue5
XwFrak95vd51GAGYBGP3YItFKq3heJMjKRDcJGh+JKQEF6oFGXvZCOcTqz2HupaO
1htfA+E9p7LWL3dNXayfRNacYcKyA/2kysAmpStFZ9rGEkc4BINJqC3rSARE4riT
pC0otM9RX+gMEJhXAYr5Vrc5N6fxQ4HWHhbGC7yvC4uVImjUsMmKTGqhcpJsE7Fp
qICFZbYJUnl1G20IQqVyvG3zS+zNl8Z8LKIUByV8gRBbL+BXgO8V8z2VIxVBvw6p
n8OEIp/D00PvFwXywp/Iz92CZaReZ3TLMYvQUecfWW5U8G/l4C2w8EG9MkujHmG+
ArjjBIAO5jESJrDilyo3gRufGGHlOz2vjRfdugMPFMZZH6SFBKfqsBdOfRwVdk28
P6VL4pNCtwC2nW11zvwvAoc4EegEM5yuKTvMYLyLuIFoKXL5goECBHXXfj6MDEmb
BBlegKXGYtk923f+mcOpdz3SdM5U9gAzGLlwJGZvXXMp3KiGqKuMbW8t19OIMqNs
gg6ut/mMoTVXAJpo64XeK9PIctYwqBNfbGBy27yxlWiOjTz0JmymSn6OXs1EV6R/
EGSM1KCQ9gjxoYt1h+D3zlRym+Dh86OQUNB2P3m29+Y/RHdDCf+Vj9Sty54uezOi
NVm3yXbzzPtLLzqfQZYG9g+3BnJtHng5qxVnSpVTto4ENZR7n909Xdfs8QcgE0Ez
nIBg2+DXpi66Lq2rc+JAfZjkl6wzQqc0BaOwY0QXrn9M2uQP8eLD2K9C5rBH/hIs
73WlMBgEcBeP/cRqCvpzGKcs59dsyOacmXeOrOkviqSx0M/wtPwZ7U5mTxsNYbUN
YkV/qnsJGLVBlddf33Dx0bdTUJ8xCem6/iq0UpII81/RLRKrOmRjFo53i9lftSIY
qxwUsVMbK2f7Yqv01FIx3LFJuMLZ9yHqQedGLAmvmp4FltwkCsVcT3+n8oJfcboa
+4KT7ONpitm7OdK3mqsu2DNjQamCOBgr3vTzTxx70/4+JqFu3Vs1FK7Em6O4i+rY
TXCQGiNcUBFYAZnx/jKxhsCJ7ivJV1en/uTryT5E4yHersoLDrwzNqiZFbPod2Pn
PTi7n7WOjKWkMoGTnoEBIp8zp37zxMPoT8daIjv828x7Al1Gz73feCGDiYzoG4YJ
3Ol9lkIpyfFpmu43FeszTfGgaIYk5pfxVuAe3dNLAykqsO5ju7gHr5SDRbi7ROxq
7kZPomdJkBMZKqpvcu+10oYSP+XiJtFOncWhh7LdZZSZ2Y1vAcAX2lFp2sME7Kn5
7AZFby/GFH98paHy488wGrbSIY6GR2tDxylr5h8nygkBtuTihR3/gVw4SSdY7vDQ
wT8PrsmSj/BglMbFruHJsQ/44IDsCx0hPtLpxDmerg4mhszJ1U4czdEUhmsjgKbd
8wBN+hVZL3NBvbVErBcUHXHaf7euLOW9CnqqsN/SKkFAXkLGQ1MXTvEj05R9Q8n2
zTwWtAQjlOu/lOHvQEi28212wwnDf7etPhei14iJzaSZmnjah80QJteAOewLfUms
PhtG6BsDKo/poaxIpPcoUpKd1Pp8Klk1Ijl/b/2Yxbr6zG5ci29IXcReqRDbzSz9
2oJUZbDIP2mg2LPyRyJ+xDEkuWcHElr8cBo1utAITM9AdUwFnM2nhUuCyXCAVyXL
CjGkUvReExVGaET22tPpAfdyV0mHvZoNgI2HYh7ASclD83eDhO56UgY5tpr0K7wl
wtekx5ArGH68lXvBNEcl/R6HWu/izxoxXtDs/UU5A9eQHpSUnWl5VnXvKk1tRR14
yESouepCTTp6GDokWXLlJ/xMZI57bEmt9yODBNxhGfYkpouTCUHnL4dx/qj4fRoH
JdU8AF1MCPT2aHSF9O6L0fC4X9u5T5tQMkNeUX4SnWYeVSNhzsgYKiCsJ504ib+E
cgTzma003DEufVD9XyICH6nVO0M9JkRIwAIaz4sw9ddBn3UAPpLpYbB5CauDF801
pA4X3wYqDThuNoyLX3OmQk6kLEjLOfrvloOe/+5yAUt+LFu2eLIYo04RaEsyPkqf
aMWfAU6Y4/nIJB7Bz7FQnn2qz6ycZPnkYzn+rk1uq0sZzS5yb7KgSrOCXe/JnqGk
VC1tNTbdVrpuxW+i35AgmjBx694KPYzED3NL5CYhQ1iZbbBs3XdsXZ47QkBCnNg/
FMlhuKtrDetlOArH1+xupuCSI8s2QlJL0c25UpZBqEze8SeVY8QvzET8WenJz6oz
1+bsQIFyjGRNN0k6frXPWfY8cypRJMeOleMj8RoL5/6bzXWis5T24WXAQxxoCF9s
ve0JP2ThpeR1GjMAo0odEHCW4S3nCtzRYA2aaWqC9Bgt1Nn1ycAKltNkbfLywKAw
d/BFbE6XGLoPkbaYZ0ECbjZbyRGOEkfls9Niyxs4ALPrjuG9pfIKc++kgIYjUzXY
Fu5031lHQmhY2qgfwmIaBUHMnN4CkghuywpFtjGP/8uRlfVvRYgOv197Dab55lWS
hnx0iKcSBcNkCNh0YdCgHLnTN0hbVe7IAIXpeKCn340BstuGRKmsoYFbgKlFnZFQ
9q5De3MpsvXanrnR3DcFkpta5XFZkDl8GS3HTKnZbz75E0QrBbUfa+2P+tVBSh8O
YkVRm6tv+Ly5xv0pQtP8irL75D8Tmyg2Pe1zPsC5xpqEuL3zsTi+XPhV35oUGY95
lwoPJGmR9q4qdc2/p5BXKSTWtg+QP1vQktiKt0DbmSMXAtGVK/ShtDbQQJqeU7zM
pQ3l2lW6OFwkuXuc+mpKrdZX1OgzoYby/qi2a/866RiBPC3Uy0hwsQS4/5WApLVX
4W2MSUBWILeTKQCJjGUF11lCFEHMbNaqrTGJqJvK0RNpUgBI0yG64MHaZEkUyu6c
Dqy321ijiNWGKo6O5ZmvyW4avrNN/KCLhMJERekmiwH+0qXjETrdyeJsos21gZwa
1od3dAtxrdNhIpy55MluArJ5/6e6WDSRjmTeZNwKYQdjsbVr5cBGdMZWijVWiWr9
oHTpEz/eYam9hC1Jhpg6wmPjMJYQqgmWzshfCWMF8VTQda4uEZWl4QHrV8Ir0m9M
ieUvD1WA82xYkNe0SjkVSmYqsuZ7R8enVFuaJtoLV0WSdPNicm9sgKDLQTYppTSD
G8/ZFnIqb/ds+R2vm37pRGMPc+19Trtggr4BZ0nl+YTNHnbQlynE9T9HPS7dlDdk
q5+cp+YIXiV9AhyfTukTwqpQpNp9G4538pu1SpaHEc5q2QJgF9GG9Gavs68CTNl4
NrrHy+YRMYh+d+s3Y9Ext0VYKrTri7l+8nG+x6lx6csz40yE5Lr4H1jtI3msJrhS
IItuhRjjkEh+OCFnbmmxfQ/CCxLmCENuVM6L92zSyINKKZJbY4KvBS1l0bCSFX5A
3y4rOSG3XMOHTBSGe0BHh595DlphZoYxLpZTDtnDfKL5m0b355uLH6XRf8JKwxsq
6Ey2Ef8dHNvbW91zYay3c6hYkPyWLiGhp3uRJo59aAkpJuA/Zh1cWntRrTnqnojg
8vc6GY5ecZGwD0aaLILxUGaIZfIOCfWi8+l1MMA4vZiZ689MJsAcRxeQlW/GC9it
jQdztXFmrCq2jmeeAzZxDB8yzCEz0D51f/7pVY//9E/MTY1RWzBoiacyFvXmElvl
8FfTe8NHOqX/9sqBitZTYCGcE1csSctirtMvi/uS6JTinx8Bdtjj5knDYxTMgnsW
1tQ1F5JOWl9c93rNOrnmnP3lbI0kZLh7mbGSx1btBjKLoGDz6QlBtnh/ytu565ou
2Nze1HLJQWXnqiAkK5Opfug6u3y54YsMKZ2OLylAGzCf0Y+ZssAR8tSrw3EYRN6n
G/Hye0gbsgFhXoa/0twYMkDYKbYYCBfTKEuyQ7zYO4lIVMfPz2ObnfY5y3MQUJth
g5Xq5ruJWZ+Lgv7DlQUJDqx0kO20SwqW6phvfA+azyHIJ/1kX3eCKja0AKsdrJQi
NS5t93NnJjs7UHZLkKdW8j2BjAffvhrXeUDzbSy7KmsnJO9zkaoRGwdMC9qi/AM+
tSQWdH4pZky5EutJeiQyoE2vVKbQOs8sx9a7qO/Bz9E+GZNIun++sJXfLOEza4QM
lIZGk+K416jLeQW7gJDkJ1qps1RWntIDXo9XxXnsrfLfunwyU2TNj68J/xBO0X5h
AyaQAELWSMfmvVmhgUaRz2wafTbklmEiNnPnFfCAflBaRKgrTFTrDn6n5Xpzg8On
XouQ09+sbdsg4u53gyZJfDaCJMWFhwC/SrHuOVevno5CQoyj/B/BJr1j/fv6HjfL
mxsfBjqJ6i55Y9wwcIJdPymR4CoZXf6W6WRufMrSsiCK/5Yy504loLTOInmUEJbP
GeYvazjWCAKgaSVpPfacv944E1G+6IAs6EW4mXfsydzhl2wIUKQKIf4CXXS5dz7v
ejIqJR0pSlUFPF4r0Eyy/dFArnvmCPDCjsfYxx+y5MpZxEXh4k6tVKW+zeEwP+/u
hmgid6hKhgKbsvmocdcZ8oUHnaKIjveorn3XRkjBsMk379Rk+faOClcmEeyTpKDm
Yj/CqFUwW5vatWu0uAITDUMKdFAHYrO37+elQt3efKxqaek3VeWKwIzG37+az4VC
AtZuMc7w4ca8u55jtRpGy+m8b4Q4D1JKzGPSfLSBXwOdG603syFgDX02nK48YUcs
Vyjh2oHF2gyN1d4iZM6GkzawOD002T82onB/YaW5vqjqncXJcw7SU8k330DA5cv+
XBY6U4YX7+Wd+WgWogWZxt23OTxP1D4/gk5bdY8X+GsjyrimVTiq7SbIkZvX0c+A
XoqDZ4gNks5o5rlta7sJjSi1N+d4MBvRmihPCKiSf8ppPzbZ6YGdQnRDtMxJ+zpG
gxk5LCkrUqqcdcSuPYfgSVLpah5s618PueJ8228yZLd46Z0ID9y2MQ2MLRA5naXw
gMpFjtjU6CAcoR/DxDFNX4hn5TVxn7MKHmH5P8Oqm2gv8y5iKFxisEQIxWBcW4OD
gn/vPCYdv1Dyn2K1kSNqy6wqSqqG2OCY3wMOtoUi1GpdU9ZIrXvIZK4hYq03oVbX
hkNxHJXy1IjF7JBf9Zz8LScG69c6pD70Z/p0RA3sbpG83XG6OMnEjszGlxjVAY1r
UaC4qfAlBg2MV5hUXXXBZ9JhoFgKfYQ49pFNyOk1WO5srqSdOXQG/qUQSEP+O8y6
j5+IBkfXEKAUG7YK6dlWduimz+Q15NOGZDM9CYAtq81VLC5Gto6eU6HLFECNkAMP
rN911ZwO+zjYpEqXCLSIj7l5vtFrvi2uovYHTdFpMzYVCfMdlkazCjyRzzHsEZKg
6d1BWtebsxjNgHeldyk4RV39A6pOYE/vGWGY3czzRDZ5rgejNkZ1okYVG5dGEf//
ttk8tlnoRy58DAjeJnRo/2OxBABDFvzbt5HTAwrM3wnYUnsM4dmkSK0rWO0PhJR5
OMpRmIFaELDywTBpoU4CYtU6d2f28B8UTapq3r9btSdHM6sL2AizGfywCxvvfaxx
VVlJLshgPUPBgIAmF0o1mGrHdSjIjmWb9aobvvebqlZ5FKE0195BH7eYEGDer1rx
iaS7M+8oXFudqdwHmdh0p4jqcA/WXL/cABHKs92aTycq8PTo6Uk+UQLxeZs7Dw5I
AT2CEVYSyniDDN5+LO/KprSkeNeG42FQW+YvtpJFmXz2PtGppduOJhNcFJuYZ1pW
aHybZeBAWknUTMjwWSW4LVhBsQfrE7taFjW7QmtAlpDZaHBv9XKt4zTeT73/QmTF
p2rOGOuRe4lgeHG+Dlnmuc9PUWEGIS0IYxQvTHQaGzaaDK23nSqEee+SeOHHzjb6
Qn0Z2sdvlmdiAf5B0Szhvc5n7ECjKKTbQFkTSUxqsDkn/scW8+ZBFu83lYtmbpPW
MD/YCR/WbmtM8twYlXtzeDnOsKQmzzl2wLyZb44e9mANuk8HXhL62mvDli51lAJu
2s1m7HSZAOyJ2vGkuPqy1XVQXv4fvWfc+fIxDLnuWQeiEHwtyrC1IbyWOz2DNhZG
3oi28UgsMo5p42CGkvdDfS93dcmhcMqaT+RmJIFjYzgj6iwTsNgm5WFwuxvOdMMH
QyosjikSSzfY5h4QVVFk7HNZya264VsGmuJyu3a5cMFthJzuXjkOrujywsFY92qg
ku3mqNeuXDxhzM7S7Q9HlNk6mO+RFiqejQw7/nbdM/aXvIxBY9lxy7NA3N7NMoGv
gLSLVFytMESdsX6rLvQWxdGXP9BmVC/ETcqn2ZtqfylQVzveybEST5u72tIBmhNZ
Pm0kZnh9u0PYMRVAJuyZGAjetbuwHGYkfOOqAB+BhrjiF6EloAM6C295dFhfWpDC
alVVCMfBUCPooFFobZ0KBG031vaNik/CQfE4b9SREMkeqUts0zKzmBx1avGieGi4
9lvq42syQFZzP7RVfp9sCs79w7uTzBJGuSpm0UzrfvCtiH4TbCFx9bKwVt1dlxv7
fEnh3Ebe+nC03+5+OMTzVtrjT5IDdWXpwoJwZDsU0uM+tUzoUbY8p8hmlMcjiT/W
czz5c4BZDtbpu8PBbbnkplCfQnGZx9jVuR/OrgrkEs7RNf3MNJX94LlPjZat24R3
OKgTE02J4y533CPTrkLpQDzNu9FnGdmBdyUdV+g/CHK4tgTCqtTBmv0VNVh3cySP
6IN0ZfgwzJyXDl8zT1p+G5JWPD99I2oOfwpdHTe4N4gTYEqEFPpeBZStUcLahINo
60geIAQaFtyABZiJNath1Q4D8wm7n9VY4EJx6Hzq3MX8oWoKxkti4NHWrmO6mwBZ
yCS84cN5Ky/6b3Lj2UyDJya8EZWLUCIGJ61LhALtVjM8zHFwsyvb1j1n5dNvdQ5T
5S7aGNPxpiE9EPoqtPeJjhzKfLrBzcZonl51kaqKRK+wYE7aktMllvPT1gDE5Oia
SpWt9pnfW8vGoe7XKRWPGqqs7PGaEMjEPS0SvDWV46jWqvoNIdc3VragRNIRaqCn
GWzWFs6n6FcZjmfZtDatNQxZjWy9hy+/72q1ov5OhdkoD4UXBelcwiv/tIQqyph/
co7U3Mmdk1F9LDJILIr2TWm45Lx8MX7xn5N+QkejnvV6i1vlVehxC0/0l+KZi7e1
/DFKmbRqEYi9GV3d+hCP6ewOJJ822bNu7sxFGGoOyAXma6XXTu/0tH/S/OyvBi9G
3/kV0GuCklQbsvJSLs6b23fnU2tZyjmpxe0AYEImpbAHgOCDIPGLrCwkE6M+OYkw
gLu+Sh2tX1L3hHwsX2/EUVtcMl4/aJW7e0YFEQytw0JMZKyO+xZAn9ZPayIGUV30
3rEESALjYsW3H2eQP+snwV3I/q288akzIh8cFjhOP6drYhAzVB918GEPusxMdj4J
J9mf20olTqtlACx7PQPJ+QAFxsOzqfzeE1SyOoYIftoeu22TxBit2qmcPuWk6KLR
SUsLa9ylav45VnFU62F7dtMFK2sRUFIea5J15EaZqkp1JcSipRuFRkAVTFHaVDSB
JJKDdEBPe8iMn0i0EaD2Uf2MqqYwsBGX8cqRipujT3cd+hyvhAqkD4Z40SqhvKDd
CwgRMYTDQ/wbJVpaLyG+Xu6wBu2RK1aIOJtj3EqJhQZ4P4AviNG+vpijtb3WIqP+
PCFkAYaA/CfiBcg/khGRKK4zT/qb1YVctmHYskD1yDqFrcCt/yYQvGQRAc6l8DHB
HeUw7oGiL/iZS4YLaJ/JiwR7foeOUYa9Affi5kgn7OKraMFYxH9P2O3BACytE43d
A4HSmj3s+zAWSPX/FcDleVUCsLRcMAuIvLSGftL5LoopKVHWAmGhfsxVWQv3HDVD
tyDGZDDnv9XrgP6dVOauqRDOaUlMXeMjDtliuSn1IFAcDDabylk8SrIi4ZmbxY31
y8a2SywBKAoeiEZPtgwoNnhnxt4/hucH7D/XrwiBimzp+AwNwARNt979kD7X1idP
mW5E9zDOBXkOrQ9jwCa/STxMWA9vMV3+w52xRcm1b4cuvhvFxUvqF1Y7bOAQxESl
eDQZ+hDgbTTCbFUmadVnqHc+gWYHyc7cd1oQC0TYmHs7plm5+GpKesWSPo7uDx9W
8nsdSh1ZTiOyA7T0uJXQerrj4uHSg66Z7wMwDjhRoxHiVQIsEj/TMhRUyr7VIOpz
KycaOWyWEjGFG10Xt2GpnA6t/lL71hxZmXwm6OA6/F5g8Vj0oiy1RXD6QLjnTgAY
Yzy9IBDgFouqC+x6Dsvysr4QeIe4dsXz6WKKhelcbdNydAPrGWKndMc+Oyt3oJeJ
C/GtfxoCXXkJtnlf1d/ZcCFbJ5ujmLjDNA8urhRsqCr/6VfJ2ZlBCzhHDPynvOiT
qAUrqZSaOw9aPvLXjIJxmQ+bLGhqxMQsrzEHjM4apz4stoFt+QlwDCnoqoKUyej+
B2WTgo37m3Buo4KptaZ2eora2LRTMUUBVePRtJWU5UrHvpj+pQU98OJqsVeyP40V
KchPhJDB6QoEVfveH43BDXboRvLUNED++YJw0VUtx4o2ISsC7SJkek3idoBlV+6i
GOwBi9RNqjFlnkelZ93DC/PLwejHw+bkJqn7DXwoq+YV2Y3aJeyg5xibZZi290eB
X3YR1wzJECoVCvKvnUQ3u59+no2ZI4UVRFHSJAPuD+x1080nOyq2UaPd37NSxeDC
f/JZkbVYy87iK4vj8ESDXpUuqkFkJc9ctOYLEIJHpylPKUoJtCToGids4yDtGDzc
w/QIYF1cTwZB2U8vfpF/T+f7o7sz1WPK45o6cDZK79cVEFXyptZipHt466Z2gyWP
38x8BwTvuikjtyncyMCZ3OumtDRoCcQHMMVOp6KZbQpgHnfHCD7HIWp0FymnCxGz
MzzR2kB8RuT+aKTcQIugOoPOaif+SEOmiigGrMfv45/g2H0DkguC+aV0o5XoR1wO
BrXMJO2mYRd+txBoJjf7rUPgPGRaMNWYFhGm++M0PWQXxboqXJKoRXD1uX/E00VA
upHd6nsth0Roqz4/hsOmpTHx+hh8l9Avv1oiiaA1//C5yBlZqQK+Fj4q5csq9gvO
dHyO8t5AMhdCLLByvgoh3ElQt/SVrDLnTIMkRcMS0bGMN32MvbK+LV5CJ8W3LQXb
jRRVZTuqVljHxoxQjYbmfgiBTneBzso1rpr3LsHWoDnKJJR/DZH3XHS03U/09wbs
D+U2rJED1Je5rTe5+8tydpq9ZLQd16nJKEJ48H2oJi4ZL+N8/JI1WDQVNjv2uV2T
aOLh7d52jK0CwAXG+GeeXj5eg/AXd+Q97QFrgVXoQYal7VqFIU0GFaFP0svcOfU0
hIU8Qlf0m6a8UMQ3ZC4WEtdgCcmCaXFzn1Z5JQb1nmStZu/ISmaeEE2PwfZTyB4s
vZWSmyTP9vtMx8iX38MyNbQqyI4SzmjRY/Ocew8y7/pglg/gl+niweCvGJWsUi59
iDQAtiZ8VJGdQJOo3pGUeRq0BjLcDOuccrVGtdrNWKOY2GYUSTSwrJoGs4MWPaDI
c03OAsb5jiQgqd7t+79cC1dZTGSM+mURwVx2c/oPhnjd35raO+rH0Wn6N2TH0sFE
a2isXIy0rXUFbtS+fUST448zp3QZdYhc9nO1d0diyEVxeJpVmWaty/8x1M+A3O8U
mPeYWmUr+ELe4oJRn3aU4+EBDiPcLFCe/xtUCVdOlY/7V/AGqTy0py1GdN48m+HY
CD4rItY3PV4mmV0S1465TcNi5/CL2KasB4GMx03l1Y3hVHEICBfZL/I8oeFRbPxI
vtkN+TryUaV3jbtcSGkRlaBH2Lp1BMkhYNT4pFfQtwOW5R6ymgfme7min77DW2Zi
Ty4yruFStyIUBhFUYbao/f8R28vhg539s8R4TwdgRUAFTLwxid2ZQdZMe57G1AN6
PHX7E2S/ksfKXPt22k6hUl7HPodgUWJQRoMdRx7VNCRjoow0GDS5nWnixqO4h5m2
jgQBzzsCuzp0aP/8611/IL4MkkvksiyetOjDG77Rh6JL4e2MJzJnR1UQ+6MXFNFE
5nnUkE0NQlNXkjBElsbKg7mmw+SrAgKF3H8VJ1xZo1TIUovyI5CwDmtZdgV6yUl3
KNaATXodh37E1WYI2H0wKR6eCSiJ+eFe6LGYhTmgCP1fJzIAd6zdq72ntU9oPVCx
igmBYT3nGFiMZVutZERysWGQ8KqCJS6HMQdCS4ZwpWj7rPrBa0RnrM1pUYAJIvWF
blc6asPepVsyhj2i28J7b8CALhDpNfjN1XYzlbPACqyIj4nVPqqGVLTPbVYTXYiF
fYtxPN3Pw9Q10Q2LvkNBJClcHsnsSLFhL+p3WBOhvetUSVCSIC0l3T1v91YXqARR
EbYQ51tsP5es/id4XV4vH03lg4C00PMR36cXai4bN4ybur7GsbolKms39qy+LE9B
OXmVgUsQixdgrob8FAed6frysTIcw1FZyC5PoGXblZSfyRoUmbEFOPYX5Nx4hebS
bHOGBfkLuDAmp1h+CKTV+qxfyBtkmZfXWNQ8j9lSQSoEmPoa4uFM1loo8jtAyJog
sIyQB6QaBcxGxN5gB6wW9E7eL5qvE3t8WTxMQOyIGBFEX7NF7BwWr0CRDi2DtegN
X7aZH6NVysLBJbpj1ANhC+ox6/V9wO2Nnm9kIwHtnp42jrGUiGaorFguFxWYwGSg
cOsnP8X6+2JqnNsZqa0HAmiAolk9+LnmiGIJeQCaxlULB2BxbeL+qoDBDZoVtEl8
8Acc93IdR4udOgS/6TwZmC1TKX1sUbli+1BcrN+tX2lgVTqA1JEfjdbtQVWMuHjz
Fg1RttF7vQCP9BtHzfZg8XTxVoq7i2qDb8TP6sJtTUa7NoUQN81A25ZBWn4to5iD
3OUHpCT2SteuGE3sIX863QJuPk6mDVpS8lAu9DmSaD1zUVMHVNmo9XkJAEVFoTxS
umDsFBmy7iinGsCuAY9ej9w074+Jw/NS0UUjsy+8SOWENpibb7lHVXJsslSC740d
BKE8QJjnCjPBAQ9d3/kTo+wpa2xAcSH10A21b5mo2epE81ZPy+AipHxqZWcVM6ut
3MgeSvELsbXwX9tN2F2kgQjN21bloM8shwvd/B37aM6jk8HINh8eMI6Hpmu2LkmW
rgQ07Cf3QX2d6R557QVNnDEkgpcQ/xEYKN14gwwKFafKaHcXMMf0NJ6FMnOgw8cj
SQF1eL+Nzm/w33yeonCFvwmO5PgJUDlZD4X5y0viyUNTF0Uo/QBzyGK0hWBkGmP/
QwFFTEUlALPH55mcim3fEhAhe7HGlzWioEOIjm0IOsGfUn2A+2zeqwRYR23FoJbZ
h4NfHK/TekBZJ0VaUrWyejj1vuXdfx5WrpE5xlHjB7nK22pekbHFwStk0O5+yZEc
ihwoB9F+QhLe+DB3XyzpXq1J4/8EpwmVC40xvGDlY+zCt5ddbGCS0zTAJLLtv9g6
PxqRopQKCSxD+GeoX3jiJDbwgtgZ9F1qiQksR0osU3tdkKW4R89d6l4cAVSD4Cv9
jpXN5C/RWPe9bj9q24lXIxeAngQD+CAjN2eW9wIjYX0txLiWwk9hxII2ZIA8id/V
yvuq258lMvQmAHeEnB7RYraq3IJO+9VS3qWxrEJ9iQBPqoSfmq+U58beAql/4xSS
WjYgeQSDyjFCTYb0/BPjabYr9IiHp55SFkGiMkZ5SIpEeBz8MApIrsKhTsaHatB8
VerWFFt3k7uyW5KntBPyhNQ4yQt9y/eMoV89Ud/OrjmmyoRAJRCylKu86UEcuO8d
tYJxfmImgyV0x/Mq/6wcd9PLNAlc1xvU8SPbYthWCGLXjfIVaujNBOnixawC/emv
DVLzag+DH1lu8GyXz84K7lahlUvEnWy6dkrYbABPu+KS0kp3v9gwjEJddLTKuauD
atmZ2zfdocP9epDvtmGwepaCiM4g8BTULgn9Lc+l3nWwHjHfL1aZ61edOkyJqpnD
8AoVVfeyMC8VIIrybE/yGVtiKYRcuXGCDLKj9OFMcLXEE4rVv3M9/edhl0Q/JEE7
3mEcXODBQVzOMc/Fx4krcSOLju8cXDGwgprYZ5Wo7AKgfw43aoATaAv7cPPiFUt+
+iZ8E0b7BmAULefV3PjKpa819oFXjwaM5aP9M9WmqDmAKrQkmzPI3iFkEms0+390
PaPXmU/muXOz/T4hy29/Y0IAnWqhfss9Snu1R91qh+R+dbmwllbcz1esB+XhPPpc
3XgNVlOiPbnYtJZzZ7+eoSwCCoS7hU9SdBKPB3af2JQvzUFlFZkrx2NwHo6hLP5O
j3372oI9BFDR3arcEan67QiHHf5hqiNiFphOrJtlpBOlhSDdY9aGtrxgFtdjwHVL
P1iFBKhys5dchGkwa4d5IEBHtg1DpVgrNf2xxZ0XAmsWCPgn2bvM4P3mW9H7HM3H
05XYSqNfSXP1/0Ko2jRQTa8yga9lty9Lz1QYvyXTKII1QdK4pn5iQlDDi5dgdc10
qBpSHz1aog/3GFQ4KI7Mk0NJA5pC92zOvSmDx+mIncPgVG5J4Aa+IUR+PBLKjfLG
5RR8bvvBp+dSG2SKuUvce+hXnd9PYr9GUTnTd1nc7/Oxy5a3FSLl/mGKDiBc4CiH
r5zlkw8pHbGF9HteJGsWJxpUwHA2huqIJ82SV2W306o5iQ1QW5t+4uvNhZd9vMhL
Ntdq4nhZGHrDHXNxhVKqGQmzwT62bg9DfjT3h30LjchVZNiD14ZCYUfanV1kVuYp
cGYlBLg+D9aGaAWm3wTrypAvtJCOtRJutJbuIOLtnhy5Gao8qIFsDcI2MSqQg1rP
881cTgYJ3g8SZFMbVCB8+qVK3T6bHTRVSh0NzAXGb2fIhTSyR4G2WYIfhDyfPFlC
qL8PJfDKzWK/7UXmypBUnv6pfV65tlAMZUW6SrmtNBZAc45uqGPotUnoFEQuhkga
ESMaTGN87OaYDxC/7b/1MmcKboYkuOJktMiHWAQKyNMJQzUcNSAjVE9aXh89zFxS
8I54ZcfSlDyUMnAsUrFdGi1KIhSPUfzBtRHvCi46SHu19VPdHYz4gUQ+PV8NMqAc
UiUrGvndAbGRV+67vf1Z0az4pGvSiOP4YHX2YsKC20+1t3SzgwWrKLinUYH/lEgQ
lqt84KP9pLWLR+ODpdxDbDcfQrUHgRohPNUvRkPoxtM/WZte1vlpfI4Eq2WXHsy5
05PVtojqqYZ2bABO7tFyv6Hv/Do+Dpye+H2oWkKlVcGr7SMS92AaKeJB7P6sJcNf
HJYUtjFHsaf/VD+Izc6AgZuM+7ddF25ZbFNkhZymWZxmRuEvDlg22h+bXavDB4g2
9twxhOy1PL2TuGk851cbEzso5lSZuByEYsfRDFSamxVxYfWAmFshhTVK/s1BI+xj
BR7KozPS5Eky/GwFdqJfB5FaSRjHbO7oagE9BjSY60f1gg16IwJNrP6xp2f6k5bt
w5UD0WxgI9Uy//xKQ7hA8IC/SVkgyrF3xQ8v3rolRmIRJGLYkzWYlPE55q6chEZM
GP/uEB6c908jyZiiaN1EH+n5TGKRUp4tcEWqduGyKfzXBJvfanhWjEqg+XQXdIOe
HP9j0qE69nyXtHyAhOPHOIBwgG5k8DwW9BTgOCwMeO+MiZYDvOz+NV8HySHIsEN6
Gm0BDkg5IXIv6+mZdUQZZCkAYnpYneQlFzLCF28+H+W01cBSVaDpC7G6L6otS1YB
9mpW153HTF2mhygty+blFrt8HJ/8K3PJ5buBO5KJOK8BMx09i4wB5coDa4jCUgJ+
1y41xu5EUV0i/4ICAb7Ylaa4rIJdy4UQ7XM73YZObne+H2GNljAygfg01GL3UN9T
WeQvQ8z/Sgp0QordEchSe7sMawR2k0JyQG8FT7QPvUvvcm4hzCC47I8TAHXKbBuE
uyAIOqdH/0vPwTDSIEKhi7k/kEOu1F38h0wXJ65dX93xzKs6hzfnUshU0KOlhXNX
P2fpSPVnsn8qcZAgz2RNESTd67D+Pven1oCWKOm2sNiqznsbwF4/XlAmrLYn1put
v19YB61hu/tPBAtrv9FRl8oFICAh3AE1W287AtMbLQhcvuatSOYdaY5kckt3M3sa
cbaGhhj9hFbCijUIotomGSqvWnLoEs2E8cyVkNgCrG3caggTt47Xq95eMf/ypxe1
KF1zpiakep3k+dKljbD4okayz6hKjbtAa3RFu6QVeLwNb9Mi3NQvC7WSYLyIRIf6
2EkoQKCqKbIpQ4T8rC9/uvRT1AKwhz3aTql52l1pFvvEPx2+yCbw08qWoY5ZnKUk
46/2DTjmxoO3th1mIIQj8ikTTEZ8AnjrNIkN4rVV5KsZD7NpDoY/BUcUgXhKaBOl
ukxMVpcfpcg00+sL3m4IxrILMjgZoTgFgcVtvMMOmhbFgOucgxJDsyMkIjk1tgcl
kKNdsP9rC1GpmAWyJ7nWVOMW/+mQkQYtl3xHAd1VVGnd9D2EsDzO+QffwPIUu+CR
MW0+0sklMxfNiWBM+EJ5SkFWd/AdHH4G/tNTAxz/xmgZTdjHOas5sNrKRReTq6oE
5xFHUwKc2p80Z/p1AnkSPGEqawJPZIPr0QcXn3CV1gPUOvx6/ZfOoDh56dj/AZiA
KY+Y6mRXCtwIAmmX6USdJuWr3uuk0mZCDmV8MzWDcZ3zU6hL64B5avrmRCTuTMPq
iO8qq7CvolAZeqJxdT2xlTtU1OIpvXAReb/UndRnuYFO2LVcyx533rGMM7DSwaYd
OnWwjT7PGWBCvvXO/ObmsqVXGMTgvnFqvIK/fZKAqTFNP3Ghjl3TqOoHqkFLcEFI
tmT3ecp6nZOcbTxaWpuT9w8Cy82Qmoc6s4G1QhXmXuNE44+ViXt14HQKUGxA2ORK
BLtFyqpy9OqVVIKam/RfHfYDQ3l0XX7tnW1lt1kdIckeVE9QEEhDMCX/ZSy/Z3Pv
J6N8uD7c5YBtUiWfwlpxhDsB4LPiZoI/l6m9WLSW8YVGENjEocE1ZGYBiCPy8fTP
YZSvLrFA8d0LEVyP651Iwo2YEvntdvnRjZkhaJAzueWlsRLhgha+qyRw4s8Vyv8e
ejVZa78uskcRQPx2NJpPLoiV2v0NnaG5TMt9tPuuySHS4cUv0+GS3fcHAw/lyZIm
sBllqmcio8y12UcKbhJ1Kod2Nbr6ZT4fGN8F9unvufAEul4A8hGEy3jrih8I05Bv
WRc1pxrdclM5nAjlw89vU3n97RErSIuxnh8k7JXxAthrWSOoCC3OLeuBEIJj0tAX
mOqixg9rjs33bX4JdlgA59orTTuGTZ29P3w7jWm74sCPZUzPOFRe2QQR0qN4swnF
Hc3V3FY4nYkRArxMs6DjHo7/+I9heZ/SJeyQVy76SJPml0bk5Gnzd4pe8Nn7OJxd
GloSYF1zxur7VZGnIss4V9Q7KyUDNFdzPgFr8wu3wy9i2j5zwgIJw4NfLCAHkAl6
FtPWgTgJTgvzTxLPXykWpY1r1D9ojifCObCOdv37yyki38gN2UYnj1xUzK8WJEmN
eVHSlhCm3qtWXji/dUshOwoZ4hdqTd2JLZgToEIBu1SprbmL2/utcsomnPuTk7TE
AOkK/ijX8hcy71a8cJuGDj42sJSWOfk8PSw1euenKkdFKuas87mJ2P3RKKWJ3R1D
lRceVlVx4hRl0LChpcJ94ALQy/lOe4Dg7sPoImvQF+u39rV6DwGBi9i0p4LmoZSN
fC1d1fO8m0q8d326o+GEezgf8K9WkwHiEAtGrggIIIRbURYJ2KOgnDQ1jzvI/hbu
YpTwXyL3lUKNV/MT1ar+82MFs9dKL4E82VnqpYNYOBDY4oTtLLIs+PeigUKGSpMh
EAMO5ZjO48QDVe5V57uJI4SlFcNp44yVdA4aE//mFFcty5n66LGH4VzWlvifDcnr
lzLu3/xXPHaq1yhiitkJNlUIy+aohPaKFfCe/p5S/Q8bHPPgcS54+iEXimUTtOt8
uRTm2R1IVC8Di7uOntr6vcEV8IXY8NLnYEXBI1T68gFhF4P+ehZWzoel2KUYh0B5
sq+5RPAElELqBB9J2HUv/bTm3Ek1JjCLl2wuNVlTVSWJNIT82JupKjmm70e7PT1+
eid6k8+er8g/fZp7zyDoAD/Fqr7/Z4inUOC2Jc46uOu0xd1CsrbnSbCwbVVsCm0n
vzNU8S9GbHXju4iE60wPKZDiY4PdyTEbJCt/lpNKKXxMEgISGsKnZqa6kK1aI2/g
V4RvfIJvrXFW6X7F5znyuOGeGjiqw0tRsEY0zLSDNZYxnwqSKLuql71ZGyRNnSfG
X862flW1bRKkMj4cekeknK8OLL963DyQ0GfLnpQ7t5E88PsKzFmQq1YVK0MYWUTC
p6TMGJbdUuHxUxFo8zI4rKbsVAavA+GUStKDjejjaLKdFBtl4g1IPv7trrM8tAcV
Di4OpgBd6N1u8q+376krAAsGIb6IY/jvAbI8bX2NfYVhWjOxQWK16/E19YR4c0RF
ZjVDn+syDWQWWh3OKGe+gUAH3gung5pR7E7DKGElR6Z7euuPbzx6soKxZBGXAmX2
6IcZ6EUW9EfpZHpS3dRTbu4QasrVjtXKnymh1R2JO+SmDg2f5v1GmhrORqbVWMih
oT9g/W26E46Y3iDQXE5QJem+Trfwvcj6UPdtvxuBUN8H2KLqgXNsfmXMm471I08M
2Pby1pzT51sB/FjYx9HAQe9ij2QgWvAeiOn1KYAzHhkkD0ocvULwMv2jRR2wFK05
PePY/fvyi5JZldwkPQRyAo7gg8gbCmMo8hbUKkHKAIug7Rsqx0yNMojuy0+xq+ME
Ob7Fkb4y3YPoKs/ndTm2oxmq7QzkBDgshpw9dUW8rFh60vmgPlB4ZjJguQGstRyP
pFoH4mqRNiM9WU+O9+OfxA7YieGY2xsQTKjbzgp3oAUk9UD0o1cdDhSERa0IMMLz
OjqOuPkHSTOCCjiU/+Ig1R9JVpY7pqfk84bIVb6aZ8j55dLLSNSSnUcO9jI/7DAh
giI3J0ONVKmDj5AwbEh+27SqQ0jriac5pIBAEMbciR48xmfBhUCgP+yTijJsSlaY
xJov5KVqi0UVzevbIPDhbgPEGpKWhLDfxgahCDBNwJQoYjRlWK7ddheFiUWS1NFs
b/8TDj2zH+k/fOTl65a6nyfFCl1mqYno/owozf3Vfv0zrTXj2vxmbMRwnNJn2qwk
wlUHO+0+eEINzi+XBrPHfs6LDg3ekmquCXlF7yh0hcwBWY1uaw2F7TsZbn3ZW2WL
YtvBn53gnCTCvFWSczRxXipZUiGthSWuQpMGgH577M7A3N06T71PKm7bvgmzzbte
jorISBUJA+1tmRSl3Jw/C9P0UrPoj2OS2UDZJEcBeFnL8wur0zbCGgwGpHzv5Z8Q
qIL+hoxOt+raAXw61HUGIV5VOZR5xum903J00UEavlsUhSTdSwbg+EH/opuFcM2K
/Pen6JPEVXTDBXAzQotdoyrlr0WQ+VVK0nIWqI71aqad4LmdJJb0XnMTQEGrBtfT
hR67XqGJ6AnQ155b2niNt8A3sfu0seXQYACUUJanfWLsZNrk/8MhmOPEyxIbmITr
85Zwdr+I8nP0zMQyaNVXduiVjVc1a9NCRx00hu4tp+FDIROaXOE+dLskrR4JAqHE
rrPqRgvzRHjIiw/E57b1eBHDTyDaxfRRdkdz04b30e4RlNfdAYr3AxSknqzUSe4C
YzLnLbbTIryCNGVdxUScIGd1/sI+CXCu8U2zzUw5a6cO9Ra5mBr96gbpuZvtiqv1
Gzpfb8hf+pwpPIQ8PikJ5HkktTCPVIcIsVJ7H4VbA2Tb7euxGZ9pJyQQ2jTZdxJj
2d9zFtfArE1e+pxuf5Q03VcxGVyGtzahmnt2WCSryEuh93/CTxDnqcVRLXXbU6aQ
umQL/EjfzeQFTC3Tm12X2pnabnwC7oCsatFfLW8KzKzZ/D/414oPrAKdibGhSf5l
GJRDgC8xicPiWU1RWRlgUZtWZAPIWe2dMxIfzg/hKw20WlS4KPXjYvikuZaCGQHo
YwjFv5mqV+fN3HaaSkv6UkGpL2Yurg5VGqHKQ2hihxKw6oNXJE0RUiTFlZxkNtJz
YOIdfOXsivkrgjUNRsfrYeDtMjT3VPjlGR9CKluPFfgIToKVh1aS1edE/K5phBBD
MM6eK1fRTjbgu2YSK5I2R5azmgiXTX+4FrMDlm388JQ9KmFdlWldweCJkYB8v53y
DbByxWy/utuRr2OvI1+1Jee99xeCkXi1VRujLHAcN73WLYjjIm2Y6ZzUhoF150cD
zvwbB9gUGdyRX1HNivmosxDYkHgPXXQFqD6RC3spXREuEPwumKf5RWD68guLE828
GQ39nTfp6w5kGwTmh42+AoNS9+J0A9aCtO7/WXCWdKnxaOHlGSRn7s/z/Yaio4Kr
GFpHQlQzNYO61ycOVE/Mnqb/3ya0tzqDhm1gih6gOTw3Du5zHIMK3LODFqICJNcZ
2OSV4bMiggqC7X9KMITgGPiY4nBMZ2pS+Bppbjqo9kTFri5XKV89FwfY6jot3TXI
nx+W4Mcq1oY0ObF+0apHIv3S0WdSv0TMbNsPbXwVnoeVLw94CMGZeNncDcK7KVrL
Bd3p4/O/yfcaUTt3kEuaW59j/5Cnf4BJBetAiu0gBZrrRsE837lTglpS+qqQvoJx
Z739WRhY8zRqIasY2uyDJU4S0Mj7OihIeZd3NpUzK/dkujrz4iaGbToNbt/hJLE8
fGL4GOnCtrZ6cs/F6KvtGwTVL97GDHB5nZD8QdYUH9xjJcWJ/z5KOXdIoIzuMaXk
sU/O7tv+cDXsRl0uBuEz1yfqYmKI56yShoIfq1UpVhyPbUsYugZvHxtdwtDWZTlj
zYcDxtJlTyN4R0Ap5mRO1C+d9bBZa8ow24JwEdqotscVJZcJcspe5KMhoTk+6K6n
X/bHjCDSlXWUxI2ZjphUmnQTxR1D0dd17b+LmA5IMddkQiHtPhLrLeZVjxk5G6DF
1ez+4r/DoCbpzEkRYsPhXYqHrj5zdXu/so7dw0rMLQhYcEo5Y82ce1zJSYrDHEU3
Ar4S2v8mpkZ/rhxlHwL29SU6cM+i58FOcZ7in6jyV4L1VmHj0W/2ruy1eFwYYDEd
tqgN4iC2BKZA+pqLHtN2WpWQ9RvTWGMhNTqzytgAXimPy0iSbqKhDRSuckQnJ/Zd
vwvGuUQD2ICy46dvonJprYMRKtcL3nowEPtEskQ85KlOaHYRpJwHzoyqSJtkM8mg
qE50pslD+smPmyFCTDzPWpBvu4KSvqVSV21eCOB/BQjnDaj0w17IvkvzEzliMLw7
06H4DQzYpIZhRJcFz4ecD3dypoTtC2SAJ4LOXhqw8V2ykgG5AOEtlenhzE/RPOhC
mHHcRlKGAvIbaa9YKy8VUzR43jaL1zE98AhEA4dh3Tjm8KGidBvRaKYS6WS/H5Kz
z78hxdatcUQtqc0v5zNp9wHF/7E0838u1oOmxxruEE3CPTkBFf7QBf5EcNPF+eyT
nTu4BF0fzcKcS+QGDH1kzGws8SN4Zt81FftuM+3Gpjganl4J7O3hNIvd0INLTQEQ
LJivwnHeFuWUF/bxPfYH+G7dIIY0icOPHghTW76X47+2+lVp/RX4oT8SWc+uAacz
ed7jSiGkSbu49MMcn1njkIoywzDUlhM9LrNOifj2rWzfq7Iex885uZFuukRK+6E0
+yWo8zh3s51MAkJ0up1q+vl0wRCAHeykL2bXjrsXfvaKDsrM8qGWY4MuFfEJm7U3
n7Js2R4Dd14jqJyCNVS/aAQytmfaEHQtQ5474MLuX3nBQ7xLWVQkh7EoivAxuRbd
Y5QnyC7T9fpxh8zVo3H1g3KaA5DBJ8dbw7mvU5XATn/w21B4YYTi9BqUDqyFXbQt
YYg2GGqMB7L166rasnHqjY2vyTeyXVYFs1kQZdbZEyArhEsOU66JpktIavEY3rZL
i3ctuk3QKTyny5USW6QqgZjl4/wnb6J2gNfA22RVZ3XlNESxkpboQ4xPCpuCevbB
jcwOGrmUX7lVsKHTz4Wyhuz8JDdoVqxENYxchmzyUfC3j5mwO9hFiTQazN4K5yQE
H9xvllUSHkMRMdypb5xHCM1NOVigHy4l6hggJKC84SS8dKnSDgFrOGQZhTwK+BXi
tBra8gkpMMRmo0DYtPZzzLNZY1AJKYTd8fGAr9uEA8FZ6D8seBMX0GbDXKSyl+PY
trPO90Q3NsrMuCMdR7j0mvB32wXWGPRmaCWwLA0q2ICBS4B3RhQzpmcDlsa+zjyn
yzHImhHzIx33mC5U5pnqi2DozTBtEYfxgoGtAbK8Nah7OH3I3aVMNvV8Lk3+KpEA
giYoWe+UREazjCAeXRL6OIOlIQCpIii1THVGgTCI0P0E0jPKregTqLshGJ7rD7yK
Gii/EO1an6+U3Tapow5IYfkt7CP/KoEWIV1uKTB+OkhqQyICiYImEg24nxqoRjPI
s3TTiW+h1Fbl8VcJ5Or1m+III63jLoE6VTETR8sWTP8g1SIdzfSBHztFe7/ShjsA
icclM4GMew0hkvcs3zk7xFW2+p2Qh9dgvdSRrmm6wjyxdYOiXM53V4lkS7eApD1z
IJ9cM4gU+dmWoOAkM4TfA9gGT8pmVSe3LrNwvhXMrWd8Wr+xW8ZTFj/h2gw5A9C8
KlVElOc6E5xQP/MIO3e/PtJp4AK4ABLppEULeLv4a8lQsoLDNIdwbEytOP+LqzLd
iKJ+9UZWsaWoNcD8/NmtHAAi7Yhfie9lP1ZhURuAY7wSj/pAALgvHUwcN54y25+H
yeLTC+fg+GUVBtVdP6LJgNN5pKz+7G09UfR4vCggKh/CpEvmxWgVZ5gqvjjHjEcD
7dVlTCZy3yeu2krXxdHvueHE75WdoSRGaW9LwaatvXi+vSw9pSEuEHuMuUMYCKLK
TR0Bzl06/d/iLowPS7/kQNBVF22P1VPgcJRA+Xo8+N3rtRIVQ0wnhop5qVo+vyKE
K30ijHjLMEfdMQDfryyY5dBUBWPoIbsLfSJQh0Ul7/A7qFVrNNZnFzWjswglYhZi
noSRVk2qq50tXityne12DeM/3hHlbkQlfrw0tiW7PF9rYfEmmU06Y0g3bAReIhbt
gakfY78LoYI7IkoKy3YoK0OZkaUMAH+y5joysOV1YdV+AtgdR2X2FavmFnNxzRPo
FP8D0dND2U6/zh02AKObPYy2TU9JV4fxHpi9hRtN3y1FjErxJMmdoIbzoU5ah7OE
yAMNjWaAoSdu9HOsEVijRKOeRhHzmBmgb9H9s+42ldfg/KgIFel/BqCm+a5sbezu
xm60EEe8c6V4oBZeI6xkOBraLm6y/352JXK575tsUzh8Vnno43W2t5vdpR4S/41l
lAy5pTYGRmptqeoGgCNYeWkY/ckvPK+XkGZKaH68DTngtPOM4olSxA1NW+8FVCmW
Uub3izl/bhEDJQat99w+IAOqih4eao01/nlSTXV9k7z3MBh/UdyALlZV3yTv7URp
FHWswFBn2+5PtWp+6sj4msMvkD0MP5SkGn9fypL924HQQEIDDVxvRo8N6/YjjxC/
KiWPPFP0VZ5FvgDY4K1CUDyZVV4oh/NNuRwdF4YPzRi/BvZ5BLeItlzc08F4u29T
L+l2GHo0TjInm6vYKBuDr3YCTsAuJ/Gx5emTLbjz7F6KqH3nIwaZB/oR5ThOY5em
Gn7clmhYL7QBhe0bQCCRh0I666QNLteDtsJSEB8DGJ1YlWr4SQg/MPwbI11qYuBa
MbhRV1JY5WVhtjLtM1PbO4itjwglMC54jDpG8HQIgyO9VXBf3LjgN2aOO+FtDHr3
ojB4+d167QmGWGCfhiyZofFCmlawzzDUKSEEy/SAzJAaYkDGMveBqjKCM1uR/WLq
iuXrUlIjnD03ABLIT4jiTPxYnOmWfbAF2UXqQ7WIT/ch1uCczfB44heqK/PO4zKN
jwav9t6yrkS6KAnAbUE97uGHpHhXoiDXeJMqcWgz/OgM9NqoyxFK9qPaMJcsrMcS
aRnsxEf99yLoI1ctqTDZSs6Mu6eLNAi6iXTNLeCpPW8T4xE30wVujWz/+YjjwxKg
F80+SAp546rha/nayrTGyfYjSYPDdzN82VtMCtUxk1BUN3VOQHyYsR1GeidopRbl
PgM7XRgyhpdUxTLdO78MSVgyOmt2L2CAWb/bKOnPAcqaphkrUpim2PcFp2VoJRHX
k8awLQaf/v6mGhqbprfNyLe1NGSyKQDGAPGoCeqr0HkgqZ4c+lFdZjsSyUqWbM53
+WDfruid31Ij9n8E8H3iFE6o8YS5MAWLALNMOkYAJwwjhsc7k3udEPQxifGbLPKr
ZmMOcfjGFjKK2Rso/mTO9NMXEycB2+JBFuzZFxnyLvytL1ZWGvwzoMIFYE7U9agf
rJHPqsr5LSs/wJ2SCOdfyxbydZqqkR1HEk+2WiZl8AXJ4ye7oQmmFIDkDAeDy8zg
IJgDdOBFbcUcoYV6PUEd7W/dPCNRlsNreaO9xF9Be7hHlDfo0Wwoeo3aEKsgGxrx
+eVeHLeuLHu2beisYx6dmMzxBm0QbcTmQVKyYDAxQIYUQP5rf4l9MY23fiX3Y2K+
gXhbJQyZrmx8aYG17AmTL5YWwQ/DpWnXXhjo1EpPkaUYJE+Od8xc0M9hXh+WAbpi
AQ8Csw5d6/qpaKnAQ/ARUlaVjsPbB/YljkT7cOBfJxE0DKBK0YGhmf5QAft9v3ut
RmMSDFdG3/pQNzZYPeJoWsEGD+/6MV/SmxznkgdrZE19iaTsBLFhGHSoDPQquxS9
P9znlnHRhkDndCy+javlA6Tc7dj/ySDlQz+RxzcRFQavRVvh5ICt3DbwaeJbevBA
c/d5p8spfwIah+m5u7sPPMkYOz/Hm6kxclbeG+VzPr42ClQJDWqo8PeZiIT+/AUH
0mRESCH01pT3j6yMAp2Gqe69NlgL2DmC6DgudhZYOkK/YKdQ/faOVLSMyC6XMPzf
cCTH1iYI8WrP1qyMd1MY43EjSK6EkC9Y/dM4RVF0QTkNcc019Tm5W17/zentuQBO
x69YsWy5GIv3hB8XX3XjkQuLP6RO/miMZzznTdBLFLIbS4QqWIZrS308gqZME/8L
QcGab4Owega7QAQQnMSs4pd+vXz8NKrxwMPDCeXvr1kAwYbZNYvE8yR9jJs5IyLO
DBsfQ+n84EygKb5zxTpC3xtrzmKUSuOY2TcKh6urj+okL/xWh7FKxJjzqLYdZsF4
nlb9vVUmFlh8lWJd0ZihJvJd5MtfILuLky8+eZuqkZtDn16gXgSesF3Q9XKzWGx3
7q+Nk/MrHs1o+1tBNC7jicbGMwppv/mltn5IgQZAT5OudMDHav1VqojVGoZ3ppyS
qij55x1xyW1L9FfYJgc8Mc244CfiKB2UFxxGC7nQ0M05oYdM8ERItds0oY46f+oo
CaaZWa6iVm8gL/qcfXkmuxMMiPeEmo6M780abYETJfulITvDouZtNbwVfPhpy6aV
WivrUZ8huGE0KwiSCDQCUR+DVpfIn9ncAtWCxSFfQ1G15FE1WWCza7taCngeEaGy
ETZpbb4ewkGseHKiBiwxlhWCyJdP20G5BcZ3a6QpBLH/UNyOovQ+fkAQiTKeS+u7
1kmuieyezNq9ajYiwzX4KscutQEByNxCjN6wLwv9JeFy8SWWxsJsUi6vYutCsaxT
hvb/3lBokof/wtMibvV5kcu6pKwRzzDgKqOlrY83nd1e+QystJDpgxg6+SHo52VB
NIc7yWnK+ExJHNYXAZbnjsN8V6Nn7l2eJsCIlXS0LC+Wcik+9u+ifkdM6vLgzmxS
etWEJ+Ev0/edrn8BQxzu08G9I/vH7nkdq0T3VL9g88s1mYtKAkb7n8KATl2Bhd4M
HrDQssd2ySGfIHgwhy9iQEAckWZL/+rnYuIs2uZqu70e1vAnNaU48nE4BJZSanqf
EQaLBhGcX4CuMaNWrf4kJ+z6LpNZBuRqlRA77kPIQ1iJOOZfhhTkpHmXDvFbWn9k
Th21yo8+sSmMW+kHVin6Fgjmarlc1sfF4k7FaLMCQvLU6WoF5eogsslHMxmZL1mz
6VwxkQBwdpggZIC9pJr5MX+W3gkhXCpAZxe4AIEmLF5YC8AyGTSLK1xi8RdtirLT
7li/Z3UWeRKo1fxAPux14njw9MKKaA9mwRJJvkXjstaAONjkEvXVHSjIbTJuzzpo
O6PFJfSuD7fAHkbpy6WQBZgsjoxDVDC7QzbUCUKNXfTgQ1WkeEuF/V/UeOg/fruI
t3hSNcN96DQsU+2VfzyiPLry7Zw9hh4GOQLN8rpnI9n9Znxku7spcYUTLv6231hH
/Tbx92BtJ877RYhdvVHCMwVJwxGcYaMwHFkOkn9B7x7MEpdzxBUtYHA/Sfc7k7Sm
COuC/wedf2pTUu4K+pHpw1ESRSVDWxbPtraxXU9Gfoe1U3D3EQNb/WgAfpCkhXo2
corXUskGskVyxuwyWxbfs3qYLaTcJ/QB/455sHXXY12kXDlpghOkuvORPeFacHfE
ePj1GsxzlW/vKbblTWOLw4hiOk6mqddZFmoghedPkTI1Ann0R76grR7hE4e3qoPR
VrMNUs9QdaYOWbvHatlc+wG6t0L5r8P3mdK15FyX5OPsTiWdq47g0rqurXrImvb2
n/Hih4KhdRqcBSqTwc2NpJvMhPUQilx+fMvBmYbtWbfEb6jdlCX10ah4gFqE8R8x
dUlLx7BykCzaLTIvu9gMGrWCv4B9Ayov54sdpRcG6kt6Mv9HtlSh6GXYxa/Fgp+E
iccCWyDnRmm6e4EU5/gu5U0M/Dx9UdXaqbahXqJ47jk7HSGDfvMtZckboOD3zw6D
Ws2Ffd2qbmOXiWj9501B2U71B1b7lCiXOnSd3Xgs1kMTT7rs2aYHlFWrG4bU9qud
ZgE99ni2jVQ7AoqTe5MT3fPXTZeYUe2OEtoStkDqckqKXQ8XQMqjvSN1QLzLDQoV
L7kZcQx/0KarTAbO/TeSMfay7RX3kXZ+/j1YjxN29xOP4B24iZM35c6R1y10kTFy
/I75qi2tTeqAGWgLTDiHfL8bVZtHFI5ucQ50kYFejUCR724ZnWhNVCwUyOYmggGI
+YJXOzsZR8x0u2uQJpIv1vEF1fRz8SSB76oF5kcP6cCnnMc+9rUtl4AqabFpI8fM
3q6jHnBIOuZtW3LzgEcV86SI0aNxzOP45mEHzlfqv9mIfAKiHvIQUW7aG2OyYY3r
VUN7u5dfZ4g/eN/VF9/FbhPav35k+t39nrNCDKjBZ3XASV8qG6WTWLW/CWW7JGWB
hMftrmMd2e0xCHrmpjYGdtXJzn+4wv0ZPPqosMyhNzhwzY30PTxZqYK31bS8CROJ
Dyoh/uUWm6ATwoTc2eSJtILU44AjlGvPSJVb2a1YfRzSXSE5splq9BYQ3oHVA4pV
W9Wc42FR95UYgsRMl1TaP2XTo4IRn1ihkOU+SSNk45fdsKKkOY6hsxH/dy77ZtKe
e6UdkfwY+tKA1Vwwls2QJjx5hM0hIe3Xun29qxAib3mLbVoC4r8Kf0grAyMdhQfr
T6fRCoh12qLTvJLqv5n0YDfSB8rxjxIqRqC0ZyDTyH0Zjw6hyteKmB5jyJvQasUv
DCSRxm+TnISdKJF8uMv0wqVqh+ZAfv3GwDaAYsrP7noW4O92TPBjlrEZJXln9AFr
QUzX4G+mdGTaRXReuMTtfDDHDaZkIAHRo2xrXcfl5zZ7z1gRQ6KX8xj196YT7hKH
fY2N81r0nVyr0Vu2AU9s2TqXxFQNJfz5dAbftejtExXceUCDBrixLX2lzAyAwtOp
5nVxOOWB22hUmNlXBoKJYyR0IXxPoJkeGZs7LXzJR0B6ojQLcMqHtGwFnWkzWdhQ
AZwuYC4XbUXb+BuFewPe6848YgExvCgqJVQVVjNmPPN6cc4ZcqXNguSPIIwNvVMq
7DbdnDyU+z2jT3pGCH8e2vKsxkKuJzsJK08iakbvYHm3UwhwNoUpGSnWrwskN05o
IkUOCqVE7jpJYkligw8t97wQPQnKPNT4oR6+RUqaed9FB+eaYhmUzDQnNUFqf3/Q
Njzvh2aWulepqSWhpQsz4U7lOkKBoOQHYHGTB0uLPqHBu2iqOvzH4FNwahseDztb
1UgzMIyl8ZRhkvsqIre0Qcz+8U8kCGPRvkUkQQszwRAF2ckjJfRoNtvDK0twnSg+
roVRgVj3G0jfGnthdWO0wiqdUiplZlUV92EmqOcZLrkCd4jL3vE6weIGNh/d4Fmw
mHw+oBlRFGN0osLDAIbbKGbXSPREu1onpceaKfpX4O17csLdFlwnyEttwNCwYQRq
Qe1C+Q4MCtBULFvt53AAfUCtDpye/EIVdaOO8NI65nJZCwBwTt9EQAWlJhPlfyn6
QyeVPCGWL51S29Y/dKsNNu6rVl44QWLnAzKjH84rpQw/W8tNB3O+ghvOZ9/bXyDW
lf4ck+CLRNXpTZYPWcMVJUw6sY/9eGen3d4P8lVNcEqeUjLQS8gfJIYtG9CjTEz4
pupk/WD72A+P9i+G9RFtAxp8X4VCoY+x7N1ZI1f5wU4cd26CKDn0lOFksIi+IRzk
xLhFBkWjft0HMClW9c+YCXe1JvptCTFCCEKgOgm0KP7xQn7sQMbosXEBffZjEoce
euEcyRhqxFBUkvUVSEzStrqK+iwejDZAIUSUjDmbFKw7LnWSCR14fujAG/S5RUR6
gWgWv95O6uaw6uSUR8axim8SjzCZGnQh0fO2cr0Eqxtv8La2sZGBGb8i0QfXqVCY
Cjn2vn1unloA7IqIz5VOb50F7lutK7z6Tj4KiyIIOnr6LIVwCWfx62F+63lQdjWM
zphOuV4hWEMvxlNiSq6yPjop24qStKBbbXRl+bCk7DfLk/gX1Tb/XtZzzBgWgSlf
WwQKbsr0IxgQrWbRFhyEGXFKDih1NQP2cTzx/k25P7FahHMwzjeO/m//lWlb9Y/X
5lEbLYrDoe8HnkWwpdrpxCPiaDIy6kNraGi/AcQfRsqMC5sXQb/G5HG4tBJ9EWp0
8aSZvl2QCtw5MEHMOqs/aq/UcScd63wj1OOltMJWp/6lssQNgFfjWgr9kfBbnMs0
Z70t40p2OA6ZuZqkd0vBgUlzffcyai1SZOYRGr+BB+IeXI6sMTVFaTngQ86VC3hL
X9XPsvdNitkdjsTlGL+k6Oq/BMhb2TBwldimG97POoBQK9WHLJCx7+qshMHpwc/9
oPTWkU/TmWsWtAiS/qDRe69xRLmRu13c1L5MuBlHUtx2QWdNV6MkkZQnHoMYcTsc
4RMEDn8ayFXGndMbMsN0Y8j1Kwn7W42pGY9HMuJD0QsBpX1eKCgNFR5C7HI2pejk
/v+db6qHj+N0sNOuxaZeX8buf1PPPVhRF79XYWecocvy9GCek+0TUdBl/MI2AaX3
yzVesq6x0GfoZHHUoVTtRUVvhwVxkIjwAwjqsX3+XnMgZKXWn5gWLVz8ZsI+B0sr
M/LuSmfUZU/Zpysk0wkebzrQlAZJkifO1KO8PsFAECIf+gu0KLbbgI6bg32IjsXm
9ESZ/1ZtyLJucQooTFVJYz3vd5Y8go7g3UYZ9ZSUxrl0gV8JCR43Ep2AhMsruytt
QAi4NtZbJz5syiw6QwqK2/TzyPGlF7pZpT76RhyNDLRnpvr5D6HfJx78Ua80+CDd
jiOQ83DyEuC247EJYtre0zIBcFe5Jj7H0xdtLOkM1CODv0OEX0CMS3Fu0iLyNfSc
ppcdyZiGweyNlt2A/U9Od3TgTId4H0u6eNTj7XfUI+JX2BOtqxgfMbSKvhvGoaP2
A1xdC2KnO/eaPUNYPFSq42R6Ta6qDg2xuaXtTxTlxe77mqLmfEURPJ6dWibd9Ols
k+rXrkhv75UGhrWBptRNEQ5HVVn25KV5ESS1jAf6CJlZjMMHyVyjRKe6QiQ6UlTl
qAjvtfl5TtjytEQ4V76xSvbsT0GkUfS6ppQ1Fu7SYw2eUjWEQ0KtpEQ6u+Je5cfu
0Bv4muYF4Z3BO+VMd4GwWESBIj4TUw5zbZCV155cUlAUx3cFUa/Adjn3aCxskXPx
3RmGDXTA6PKNHywccKCTXAWJSXjEg58xMUGsGpToB/jGNBt8ksyXJcbfOMCDop+u
Rp4UBQC4+IC4sE7w8gmISWXiSWWGx/Rw22qXe0/ic1lkVIxuzTekBkqLeiXGoyyS
5ge7L+FOKznmYaNilpCErB2hn2G1YaUQ+pBKC27tb1jvbiP7ixC3f5e/bu3wQQDx
fb86lpNN/x642/eDsa2K5HoCdhpWzK0aN6Rd+QREEAUb3Gv8/ZpKMGssmfPKFHTY
CHypVGnf5fBgmBTHZbfXwSfTxlReQBMeV23wKFqiFwDM+Z1uTxUTm2eZIg19yr+R
frLluLl0zG3ge+8ofyrYDQtR9KTgPbAP+d9L3aJ+GXTeOp1HPc3BAQ1ldgM3yXJr
aZjIcSEnbP/tFj1qRsqpTt9J5laBfHsw6TcKWa/Xq3eJOy3hueTIMiguxDLz8J9l
rSUqENYBPADOchGVVWZ2+JuwGPZ8y2FikpU0OzfEhnOBzZVdBf/XDM5ctqjX1gC3
TrnCJasNMyE36VygGsDc9P/gp/4rVIfesWPkTstCD2TLnbyTsuV0TiJWC4NsJJXz
bj/9l5j13b2zCxSEfTUQaopqAbtXXjo3QVTgJuXR/fwfL+rzUqubXCgKB18kxtEx
drWObaehtgmLzpv0qd4J5m1HNKQdCRF6IALFING9IHtAUtHORXj5RCVksNg9e04G
uOywJyeGE43apPksqdQLYXsHWPCJk8GaTH5WaT0R2j3OHbCwlsAIm9hKqHAAHv/3
w1sk1sqjkLnic23NunlyBITu+GVRr68wlDepaH69NbFj0lZCdMlq9XW60ppgx4Bk
RLoP1yC5jpwCKZ7C7x1bN5yMBL/BLCCkP22brhbHRhAULn1sqtPND0W9mhUgawwk
f7Z3bhqsHTRqRSGQ5RV0ZMysmP3HWwNesjfgFhBXbGXiSretvj3dw8QC6p35JOoQ
t5ykvsB3ei1qgQ7SheygG9fA6F+cqF2CBn5UgL2HmRCb1TTMIl9cpBzHZAGN4F6m
4kaliQR2DTi1YERiyY76ph/vKNHczLCkIjaUOaVlFkFW+0UKIQ7/KUbOiNzOGnii
Rxpzi9IkJiPrjafo2+Scz2Kw1c9z9E/4JVwmt4SFkuShePhOHThaiP95KBzY6Ae4
pkbnZxTbeGyk5myhzjyLMuJY3vRAkxHIxbvssu579KnvbZevLqMF3tVwvlRkQjwD
eMTcwR3s7UqKGsSEs71WOkSLIbqytoTyoASu7VjAwFJtUgMNYRsF++1gm3cwKISp
DIEmk07U4n4fTupUyLrxZiUa4kpm2CobxKWDuBq8PIFKsc9dme8kM5rQyeUUfNyG
Tgk6+Yk8f6YuUxTNAisQ5F+UES/lnT4VagRb8SVzmpdo9zgnubaWpm90HVW1LIm0
TCCwpRd7JkQLM8mUrIj4KCe+6vEs7XajQXMepb1StqiVnprdl50ntpLZN9RD7Nxn
oDrfxDA/uvueUyshBih3+uI8drpN22YWQUm7vPPydF/v4ZrxSbDN8z9zBSu42IQ4
BA4g16AIIyYFp37T0woKK/VNyJTO7uN2+B0IKHod8/M1SkvroThypxm0Lq6qG2kw
d8rTQRIwJhFsbH304iT77Cqs3cr0ptqFpuCvNmNkhPrNK+Czx9MuKLl78d0sF7j6
qKHx6VNC6m/dRdTQ/KgOHwd39NtOidu7QkK8/UT1sgxyUn+lshcXipxhpT6SgNlU
3v7XEZIQuVypcf2jSIv1okRa/dUc/rRqtqmNHNvaipHBnedQ7f4E+5I9UP/Lw9Lq
pt718ZbA9/3LrumbUF4CycRE5iEN5T5XoSRJzBG7M+Vo82pmCRUPTW7rdQhK4LFY
mFQVCK3V4wZJ1F1ugFsGot+5GpHZmQw9+7EKkg9q+CFCUonQhoaorFBPmmJaXM3v
TkZ38AoTDY24xaoVWQAZvfTHJj4F7rcyPkWa4tL6h9MHzv/a12kyAobWTSZLjK7E
crOBrwADx8Ka1KTQupxmPZQ95QfrIgy9w880PAoexz/qu41o/1Z5EGJE2U/MDGcs
HfmYTUHeDTUbOUX9GJ7rVWpHkwCh+vEAuQmfVJ+Lu0Gutu2FnXwhEVYYHWY1CZ8E
gDIOmINyQHzTy2HsGGP5n24gfeZ/qA7uCgXrmrJCtKzrPhznXYxPRwd+Lhog32sB
g+eaX1MGI6pjPP5c8FOoirLQv4y3NOGeyNdwCYG2S39Cb86aN5+YArvkrO7CTmFr
sRdXaebog8P2KxEmPJQmXAlx217HpjxDR9gEGd3dQ3lxmq1UV7xZRBDTX/DjEBwF
nDeoslyK7CmWjeg4X7a6yna7pSJILTlCth5tSvK0Q10qp88jhelt+7ig4Gui09en
USdh9CeAC/CUrXZDV0Eci8MxsmDT1q6VA+j8xL4LYccupFPE6muMwaO3fVHZBXSC
Qej4vsOV+ehUyondixBs6357r/1kqVZly6QcySXGpGlmc2ogihYvWBDOl2xj/s1V
nGtr0cHBTryhqluoG6KXmtZPNasnzh5CaQbWKeorlHYvC0G/2Hp7KXWWFXLCEnQF
AimCuepBmxJTWd3qnV5n+h1E6yRjHcZf9yJthxWvOKq3/z9Mdfx0NjkybItzK4tJ
QU6s6W/YqYBiPBw8cCqllmpJXa0vhEEB8Rc7IFQ9fCv7c9X27ZINAX9Rl9zNusBM
uwGYvtJPNBBYu+k4ORZeoYoAOIVODF4LvXbpBr5slzJcjh7oobvGqX5DBrn0fQCp
+NTrNUtIQB+lRffgTdK3ro9G3v0pq+CqNOYpjkNnAeJK4Mhf4TX0a2XFvOpVuy0b
vRvw0OLDytdQkQ7p7ad5XtxY5qXDOgJErNHW2y3iNstXiNFIMIl8ezYMgRf2Ez93
vAzOGP0+eT5wS9gadPc7yURonmTUG4NULW299iuOB1DjumnfFky/Y/w5txoKQrIx
hbLpWNr7KNAG42qOc5ySWBQm/XJnRdNgKx5w3tq79Usvcp0kzoJuhSHTHdm2BfVC
MzYjo2FRulZKYG5OIhzx6ONQiLmYxvSEUwpNdjY7FMOoYTEHGOZDHuVD011wmT7w
qjUXgWb4gCvJZzX2swkYF0rAjCeLT1Dk4/h8g6KnIEEDwJBShuIusTUqUWzxCIz4
uXh+rZUTJI0vS1cjEUkjcIvC0as9ctvQKOFZby9Anc8XQ58ggq7LSs8C+PgPchcB
C3PUUx3o1VsMm+7Zu2Wze7/bzGfB9sl1w0p7hZwjKcvHCF+gxCVB5vmWiFp3HMyO
pAAIyb7hkmPysVjazQcWIiDo8tf9a5R56bW/p9bhmclIl01VZFJzt1IvN3Lnj4uN
2Lc+jTRBWQ7XW3Plup2fI0K892X62Lr8fTvAJg47gJ4FGocRFuh3fYSf/PgpuFdl
hVbjOG3zKRqYpXGhS4poL35+tGiOguI1zZkzEaYokSIrvZBscwRSKFxkkLriix/b
8BYBcavBi7n1wmNDDuMMB9RitPRrpls2MqQw2nxn9ZhKLgxREc74Gv7bv+53VrcX
qZnQOKP6qYkAbYdCqi//GtOm+rRyInWcKMbJgMh6TmaQXtXuXhepFuX3giV8svbI
1c4K4fhePNHS90hz946mlGdVV83yLkPsz3wBcR4SQhNtlqf/mvkJ85YlLo6PRmQD
Zq/g8wThj4tvEdUg3zGCtLZ7B2D0yTF2jQP/pz5eiRYoeW/qXL/DJp/0F7QEj8lO
y/mmJAqSeBP1zEdY2exeNprJyo2LGbJP+d40rob/ziTzj6LG64fvw3dGeOuCJh6V
V9rHogMNHpDr6YT8VJaJg6ulV6K8TqavqU6Ja0PKQMbRu67B7PDX4EO1/nmjDaxG
cMv5AHYAqpokhFitFeY8q1wYwVmWI7cp5+XU5YKnfSNYsHmB0mQY6o02VZnF9rDU
npaJRm9u1TjMuKMH53Ot1h9wpIg8fR8XYbk/eMKWgSJd8x6qzZ7X0kUh+S3qa/io
G4GZAXLkw0aQwHih8P0fDLkm8CwYChVRaHHHdXqTgvoPiiddDp2DtK38bemrPiWp
l6/RPRObmFM03+79wVE2FaQx+S+SjeZOJLQe4zFEOdTGnTJXJW9H3qGsENyFeR+X
lagBm76UJZEw36mAba1DGK6m9FyCXjpd+qG3UCbtrr+NLQoRX7EHwCmoh5A/5s68
lzXobjtyppyTvtCGRVuHF4A3B2BO0D18WEpUu5aBVXMQNGhLZyMkk/gBuvyxjmEK
kq5NoExJm9MakG3nU9/bKzgyhTi1xzfMCxEUTLW5kNJZLtxFb+VsA7qJ07zU0Fq0
wTN+DOkFYRkx4cCmPAW3GgmElUQ7rYRCT+GWCj4ZbgK+bk4HnyEOZxRZDadhz/ds
s9zAOXv82ofrVI++QojLewuOxRKGlbRu9QZ7MTdhNb77oq0c59YRUdlemlgnRCBP
XqB5APZgiFttc+mRK+hd7OYBUloA+gO83rHftMRgcvWvYGPsyQrKuXMneKvVimSP
px578Gk97WPjyXyRpIDkcbJd5zLKKCwaYRmJrXV/FFrw3Ykm4B26ieAqD0s/xYrw
HOdLYF+jeFQuFFfeRYaQRQPPAIYAqNiYxT9F/gTQfN/EXoWqdCuoWZkECcR5acz5
frB9Z/lmx+5nBvULZsl0q1OJjOyuHHA0R4SABBijNIlcy96tGhXntASCy4aMwtDt
VlEk+uDqLEawBwU6fG5WrL6iDvte7nnweHOXGuz7g+PCR/jqkN5jiQ2ERu90Aw4I
ETS5+dba3Ojr2KJAvKrCvZE/lEYBr/oBbJ/19aF0qwIfA65SsOonllX8U64H9pD5
tB1STVK8f4tVzC/MP2BUC8i/e4Tg5qN+9RC0swsHP3s99HeRQ67DuJFJjdbW8kHM
rF81w5zK5fR1QR/9P4Ug1QS7k58OzV8mWdbRBEQVcRKEkhxrK32Y2tEk7iGSfG7+
hXHQGs72F3Kc5kG9qjwrDVSXq947m/ALkxWHmai9H/eWHVx13pED3eSON8HJlLtq
0Ce9fgkHaOLyH9RmJhAyL87ICSulQnTCmp6XZGsOgvPCReK2aU70eO9LLzxIYvZz
62JSdrdu8E1Yz2sYQ3x4zFuSYgxmExCLWSToml2R9hy97iXXBGsrcDx/76h1cEae
RmoKjd67vfYsXFtaf7fmU+oYlW0PWZI0KK6eZZghFa/FE+oXjQ3jqQzqmjOg8eSS
LTA6TJ9uZCDG6eYO5h+PVnXVDOHiw6HnSp8mrOCk100O+ssBR0tYQ11g8SYvl/J8
47CH+HgC/nyQcnNwz1HlRO6PXQ8Btf191a0T8APuEdnHUCmvUCX43d5IKtQ+Cu8J
92raJrKxmX3rCzT+SVpebhu8X2eS3mTMBTLbiyQeE/MPwPtpG5aidnFuTsfaZZBt
kUeBlyOcLOVQNOp5FMOYvTjCDvfYpQ58MRR2SN2kjMrnFxMkUcCZHygsx/VVkMlp
+gNB9kPDniLkI1+pTwAX8uvQdgpevVJL5WVv0DjHMxCBIFK6IZ8n/bsu3DZ4C70l
BKOmcTtHkIQV2q4Ildzbz+CZwhFvrby4/nOViAS43XDVyw/j6xGMoDCGHujbeCdK
4ULBA5pEJfjnamyPRFV41Xj5Fh64VzHOAz5LDGflyBWJGFIpRGtEZcjH9baC/+qB
yeKCLwHdXqfGfe+FcaYVLYgL88Aqd20BHbOujraJhZKTUVaPq6SdqWAakF5nkgKh
FuiDWw4HHRoBcum819eWLFMYZZTLHMncyJPsToNqa4OApQQWei6jyB1a+8FKQ/Lc
1h5ATv2haZVewmMx7cXoFZrc/POEU980mdYWnlKtHgJEXMv0bUiU8gZipXz/oXaX
w8JKaXhv6xzaaaYy39vSSAKdk/c8SQ+HkeHA3MlUAhIQ9q1d1OL7lPyDC7Zpe8VR
thzV1BziyrInNgpCAreIR3eDbl3GQ6j1l2OhAXAbXJlbW46CK6glwKOgtkW5hczs
wlL+9dZYnNTcSbWUxFJGrlAhO+WIS9G4N6p2sSdwQgj/rkN4mZdECB5b5WgK3a6a
Yh7zb5FchiGfjtXFTj5g0OzMCm6YrIA0A6bqKxEGubVWsVDzfTUSWOrBpV7wBNZp
+syy3yli7seYGLCUGAwjcn9E85zsKWtoxiuSxpGJjXdbW284mQSYZRrczJqeaImv
9oV5FJecQgKmvC5524hOoj3lxj+m8HPtwiY2QNc/4NbtEpB9DwxOgUGEyIatd8NI
z6Vu6bDRdtpoeJPJM8NVRvcza5U46cRgmX2o/QQPQJuOE3WzqGSOY/8v+9WPA1ry
+njWtQ7RxTCA1l/Uuk1GI9/2/3fIsMZ26uR3U3iY7BHMDNGywmIdgsrmMFaDz3X+
b1sw0X76nBTifVwaSo1nfPzKYlshNrJKfWu45XKe7/TqQh7PvSihKpav3v/3c1bV
LcJs4KVQErrLSpimguAuuPXo8RpGDgANVNCqkej4w3VAUSh6JngSGovlka6e08rJ
t+OQHxg3HNmXW3MXcGSFFFELedNvfkH00iuGIhJop32XWhW13rZc9aMGQWyq/p+9
C7kjrfagDHAgcDumLlKWXi39XjOgtRmySSNLzqf+8M/iIGloLUoWKhXgiaViGUgH
1POTtwwWGH3F5oifFvzknWN/rL1G3Si27O2h24Ao0ueO3ZjnWClwQfeJ2BRX5HkY
B6jbc74oQMmmwEXR/zIWQwTdPgJpXjyCYGiNip+nZ9ApJFooPkIPuIVQXuyGH7Go
KBGr4PSmWrlBszqDE/uHyXg9VPHIJnA+BjIdVLzLa8VGt8B6KNNG/SPbFTgkD8VX
YurFdQoM/oDjk4HN4fKUhUcu4IjWpuH7r78Z142ZV0KZDZhGkNpXUVdJtu+5Zw2d
YuPCuHNwkL/L5hnS0CAiOu64G2xwQb60ZwcRwhh6t7Zb5bpdQyGylmuJhmH7/hsh
EmU+MJIuMVE9aNrAeIE2MCDVB1QrBXDqFrMSYKoPQG5Q7JHTPwtaZJEPvgTwNgFv
vFyMxcZq5+TpUq02/p5kNhimnfGoIRdKMSwtGFwolQEufz8o2T/Cd14e2CRY9b4a
X5aOiBhRDZufsIukbQFYuHHslu/HaJQbTseHOmyLJQCtyA9M/Awa6MiqST+8NLXN
RkVHpNnEDDrdiM/jWNwke5Pc82u43fX8sj+LJZm34BiZGFO9dO7pA85imEW/vBCV
g1ZaZo14rH9j2S/PV3Z96CUaUjfKuZSvDdPISbDTC77Ajw+6Ah0F15mIELssqifs
vPi2BySUYSAGf+WceAEjuyoQDRkzHREAUUIQaVvSvyX26niUAtWlHLlW0KZOiCqw
wQFnQ3rbk4ipVZDJ9I2zQq0efMM+4uw0CQlyobdeR4Mwn5HU7T72FelQyASZbUoH
J9m8Tc30fvsKfK/de+G9Ced1NvmKnrNTDx26eqyrpqoCYNCMoaDvtdcfP4BZgAB5
JU3Ip69JTpJ8bmSdo/gqTnlfx/laPpVEGT/rKBfmoDfX9MXn0SRZfRTb17GlZLmW
EqVfRD53N8jWzxeAGompTVRYXCKe7NmYZCdjoCLSojODA7cprMb3y3/GbYC+AJ2m
tx66bnu/54pZ8gJoy9AsPyEdUkiEk1nmRmGgQFHp50xzMuI/tY1uV+gQNGkL+wRM
aTqU7hbjobWHrX6X/HBdg1KtVUTMT6WDkBLaE2GhCvbNr9wQ8DFJ5JaGfHt4Ufrs
I++r3ZXjN5XMEGWTlEb20R43pn/RanENs3g8jOLsuOBt+di82clOo0ESk/9Qfg6o
yb0vw1kn7Vl9/tLmpKuUc+sQxX9WYNdCH07zoGuR3vwT4F9CA7iPWLZ0AX8mHlXS
RXgJ3Eivhi6PmBz9xRfwfENQUSEeMqTQdTqppLJvYfrCg1kCfwREUnmZdcXTKGZ8
yeeP4sKQxs63rqjvzY74wB1OhmFBmt5JeHIGrgNzbm4K+JxIQWkhWBQ5jx8AKJ01
APU5dVSxQWsAMEmV5Ka9Yyy3grimn39iRNtjyp+vluuoltbt+jcNxpeDXEP77NlR
HXmvrtIwOoouEfgwUZbtNkCTQg7xs4WQTaoY0cEO0Z2ceEYJUIgm+ihdUTTIVpRi
svp8RSUEYmJoh01+04e/SfVGLYPyNiquQoS33k5I2tx0AdcPtqhsfzvN8/vIchIW
D4zxo1fvKQzxqyoqxR9sTuS291DiCcqt15ZDY/DIG5MJClufkZabg3IvmV2kOdfv
D9grWxdjwhdpSvtufkDejDzHA7YlbCQIe+yK4/zAGMuFY6RJG7l3OxvH5KvRkEJN
9qvDCa0Faq67ot2Edh3/6kouB9ZTw94eKF3kBvdwiVuwpRgHqQo/nzXHfe7VT3ML
s0F2cXcrBqMbKILfKA6soibx79O4it9P9+wb60CJCcneqV/m/DBxTBkpLIGYIo9V
L/RtJ70n+fQbiGtE5jBWoMcM8kQzueki6YYzyGkue02GO3tQ4ese1mmDgyVr0vYW
rh7XZLbUsX3bwOK3C9l2PbTyqG3CynNqGsb7vRsz6tB2bWtm8Bdg00CqionRkYER
uRJh9WGGQc1KoCi9FjkcYR/Dgfl7wvaa342YiFmau5pbRpCKbmGt9EjjryZ38Kiu
qPKW0KjK1Gx1KR/aEVJaTrGorw4kN8+Jo8JINhSXUnlyVsSNlX9Cq+E+M8oTngWB
cXtoervSvPIuwqlXafDamLcPBFKyy9Jst/rqye3GoBbxUHTG5ZKV3bo/v3h+AZLB
f32KfHrXO9G9K1c9tCWHJd3oDZ4tGH6uL4Fouu/xlED/TRnv/BVImQhZjVXBgbjL
l90aG+bcyUrePuRZ709mbvwxfKk6LQn5MwNSQ46eBffrHezAl6VHE/Ne9hYFVftO
uLqFFuGSczMOCcDIPoZv9/Qo4gPVmpdVt8/ywlOfoXVcgsboviaiw6rfS1lWxUwz
TVM/dPPlzZhhgbbI2QHHreg2w7hNApcTthqFeWNSBGYEVzXCFQXLiuC5sQpF3K6A
xrbfCLD0qx3AbfCu8pJ6UMElSpj4PwU0gpmQxPYvqhybCdkbJsEB9x+AxzsU0dv5
t7vlXS4Hsxd001Df8ZHbGCGGMG1PUokGKLORh2jr5MISiuPP+QGCuPW/et2UyV4H
/B4xOf2vuU20bH06OLnN4LIJ9ZkcUPd15y5iZlh4nSH15b/B2ETtz+vbAFYu/W2s
qFaLNVBozc8bo0MV91GOI58jaz6pw1vtft2FXm9kHQBp/f92TUDU6iTK6o8/FDM+
UHjtDkF14cELW0XHyzs3KDoNlQScWx1BygKFeVY7MYIKAv/gapOK1nDikT1HQ2wL
Djd2d1bwZb5XL64t0bLK6/+IMXXIqs6BHHh0Zke2TGSha/zUtfReN9CWoPO/lg98
Zj8SWC1kHEH3aJzxX3Yl8REOw/MiP1n31rZ2o7VnUfp4uSfEXwb6yEbqww2WabCj
XNKgBVdNy1Z1K0Pb2GM/sEKzlci72zQNexMnqwTp4t1xEmO8RtTCodbWASPe9Ne8
dxeijKgLH6pgeTxQdF9Kr3MX3NK8UkWU4m+ArgIgwr4P8XQc7xRbQ8qw7cmFAtCb
pfdgW8LqsLTzLS2OBwZpoA1uU6qlYkpPi7FD8j0GI7rb+meHYsctmDbnpI25zeuW
5d/02UgNePdRwFPHG8pqYK8GOFGS3pgO3CGfIELVrsT4gB3Hgh/a0oCzABKrrkTG
4NwcBsbmD20g3VMDaHalmHNT70SCkVJls8ztiErKr3Qs6EObGHPUjya5IlBKEVBz
MT2d+HAqmTbgUFavOOryZBLS2SauK4vkJLynW9HlS2vaRRu3FUcv+/z3spH02NJH
DkccmSLufOk7wRNZRvW7Je0ISOVRtBb7Qkqc07gBqgkntdMUivIVXZdnZQYeD7KF
oXksSrcyYJNAux6DgiYLft+nmjdR6mg2hwBhQPtbJHyR+oKyaCnhsPMz9Msodykj
YxiEMkqQd69m75D2eYa0zDhih8I2kKwlWIMUpiE/lBBAO9nJdB9g1cZyh8oZ9apK
MM6iNrUNwIBscmjDum7nx5QWynhyn9Cvt5WgT4jPq+h27F+CHfTRvj8LY55/p00h
1lXu0Pwj7s2OIYyDFv15hI3h4sGAJLDVuVWHj7ZOaviE4N03siyXRvVYiZFaXX6W
8I7/3MUDYufj34WyTfh11Fm68/XYz3oR1kFv/39OyF7SxGxe8DdMdl6ihQvRr+Id
G5YoJyYUTqk5x+VmU3RTIsNb3XpOQLa8e+TaAw4MXYw8OSW/VMiU1Mm/YLd0ZK0v
SOYrJo5/l+ea4sF3thmwq/opo8HkSeKijoerlxd3cAGUIZOBxtcAuhtTCIDS37pc
bFP4JEEVkVESHuzZdwHUVdhOBo8VLUjHWbhDpNlnfnO3as+HupejA/KNTeCI4t6B
83zK2ZnadWTOm3R+ACiP81fwh8P+HmCuBG4gQVeUEnfg5bRNZb8tPnIkRhb0tG2L
xOwTLw0seXCb24iF6Lxa37WmvQAHbibXKAzPC4DWNxFiGMZD1dsXcpLtE8xX3DLq
s/4VQ0pWgJyMmO8INha/6NSwNUBrOBQB32w7dSKPk/wwcCQH8Nv5E7s1uyPCZg8h
h3CBFV9epTdUWPzlSSWgpbPoLzbu/slHckAZCOwz11ng0zljjyXsYlZhGyuY03iK
3o8xl4el6FuM4vLgQF7QqtFB4mMfES1K/ZdGuzf/j6k3DvjxMT8trNgQFhgwHPWF
aX6Wen08D+z49uVOfEQC52BMTjuSp5WIksIKuesANtTwDVewv2McC3L5vVx2Wvjd
wKXl3rdi0AIqUpMWMMaaNXYdRRkXW+NsOovVp5Wg0c2mAhPLLHrUA1B1ruLxz7dV
81r5qx/VWKaj86CbT60wflNYgdABpnWphEa6m2eCkz684qd7Aw66Tg9Sj/UQF6WF
LqdWORW+n9WepSqlksZWMmnTMZ80Gcmu6Hm8ITdv59KdystXdPDkT3wOIpSUhFDY
ztu9xBY0iB64RoOeT4aYGTD57Vu8xh0h73h/JOvuXM3toDRFsxGmMuoTH2UL1Aic
mu30ZTjxgcsA4jojhTAXZHitrO6pufQ5opaAEXA2+6wwCdrUbZzUUho8ZeG2rVXd
aA5wEhsA/QQOtF3lnPltkLEiyqtfI1lmtPqri4wuiuBB4gnVwH5YF+VfLY/hF1em
XYJpPoZoUg80OKnAClMfAGLqDQiVMh2WHv9vWDuhUyiw1X6hwNNHm4Thm6w8BZ7d
1zzSsTWayK5aGZcDCqoanpXrkUeXGMbXL/TiNB9U/Bhy+RCmkYw2NgLm22hflisi
2DkVAFsUpbA9ax83kh7677UGa7hzjlQwZzHxrzu6PtcZ2WJSR7ZBO/z5RK9Y1sKk
aeG1vSR93UesULg5ukJs6hdIrni0haPOH4tuTvhwrSKcuVuHghnd0qJ5F75doBWR
WwSwgTr4ihA3GGqPoPglPdKCyDrRzQDECkQDTUBmQ9GyWyTfrfIM3nndt6wFDPMr
gNy5JxTvgoC4CSknq6bSQQR79vgBcclh3Mf64XRsT+F7Ej4zEIf5VJ6LXTUB37cU
fYzvWv/9YUXTe5I861nO0P7oVMwYKYH3eiq9BcCfTYvqRFpp7sqwkS5lGxFvU+3q
obAijmifK/nSfycNWPSdGJL3fvZ07KDKU4g2IRTRdshwJSkMS4LFm+KuVxo7YG+P
7tmatBhyFLRfybWu9RkaZOCzzUQ2If80gbFUDS+Z9mcaX1gK+exW5OKR6sUUJaTv
lppjuli5DeuP1nb1zWAloacgoZPzSM3IFcKpvCibyn5q/ycXVP4IY6Az1Ant9/Ii
btRJ7c+QZ4d6GTVNXxDwGjbwWYa+T/lusT2LWj3Ldc64Myv9Uh/bCxv+5QcBChBZ
COR0OeOkwQ9pAlZlTLjL4MyXYm6fs/dkk/qfkDupaNf0R32gvIk2RRQAKwJvKEJJ
hzAtO00rqw8hzgmSJht5+SvretgRJwd6YPjSpLMnrzp6nPMtqEbHWnCuQs9CPNly
9sJeo1VAakQLSdznXlwrP1A5oS1JJLlX45V+sy5uNwH84oFGcbiM7LB7DbVbT2Yq
nLoPProOCsf7P9pRGZTzP22hYd+6woqaU/O1dq9WGXv7wBAWcDksp7ULqiwQo9cS
hkD9zaaD0FHYwLTWSif5dqX2nwsoNZGJYpS3NXmDLsbKKhGIVagVYV4YSEZa+jGh
xYWTtZushOTePbpibPsR35g0QC90pNZHDMnzSpIRZDlcvbhXwkcX4bO4mMVHveQ6
6OlaE60jbDHwerRQPr5YhRm8zdWAR6Xz0aW0fD9jq/w9cWeJrASjhO8Q/tti3DIp
oZ6ramkoDuR5SFfRFAPxpU43lAoFvCq7hhVDCfWFj/L9q6nNtEhxAEdoZyJtTsA3
iRuDaODB4HjmjgLc/vh59rQ+qbTLgQurilZRWD5zj6nrHXzzsDGVhDYnlTuZAqEb
8gcO2+hs5sgkv+HlNfi4Fuv3wLc5+Id6ZtLkWabkBW5eL9XHN4USTsdQNPNC6Bhe
UQrGKMsEhNv9EOm6C+0Y3NGYWrLT8CDbU5ldA4gWXJpEQQ8zxWvUPMaNxUGvEVzH
giI0/AWseDqj9Gyr79jHWdtIvLvvTRIPX5ao3Dva9QBz+okCaHMzGBOw0j4a1WkN
D2tit3MtaJyDso5Y46SpuVPM8hy4j3ZxOwxWRefKDEYE6vetCDA4pjltENqAgcPU
HX4OkfgvO7vEwlsiNXQH2CH4Zg42RZh2ypNuBKxl+IWC0nKm2rgfmMuM1TA/lp/t
Rak6XSVQ5R2pvWHPvuu1vP+2mSKB5zpkJNjrJPXX+4S54RD2TA58ruRPA3AzW3O7
neB9GhPQYNWHiqgAJ2W+iX6Z6tSitodf1Uv5//uFZX8vRGw2nlIeDvST1ZhzF+pk
+FSHrgPSf2/GtOUQdFIvFzoY9LFPZqEzhRjVQqlHJYAAt2PmVS7e/v8X2K4wxQA4
hRH72l6AJrOPWI9RFmcEb27dZhLVLbP0E5NDNdY2wTFW4nUoCYf3t7B9VAtpYrp+
fYDhI734SctDu6Km28/Frdfc/rptXmxWew7j+4KLuaIOlJMBUqpiy8kiBrT7f7Q5
AlcN/KrnccqI6Jzp4ZRnlh8KfOoXMGMHSeg71BWTXIbGY56WiWJC8zTse/mepJ7g
pPFnEBmwbp5T0g3DpFAkqIiaZExwlM3yy48QdgsoJU09Rn8LjdhTlCpmeAH9fMsY
hAVjleliLeT85VrSWi+RYSco+6JpOGI9mTeEpJU6Dprw6WGHYPBeg5mumailxx7G
LB971MKVQsx5iZMw4nmhhiiTL7Hbom/Y4hs80Fr3LUZjJg1nin+q+cJQYWGUb0da
6e48DAD7Zj2xyIz84ipfLczjWSh7/bvD0tG5cxc1siPTJmTAJqYw608zrJnVLNRs
YryFODNF8h9J6wmAYYKTnC3iDLbQo6DTHQcpvphYNg4lxTWiqmXg1ilhEIO5ijzI
Zwp9mzzd0hw2Qx8t8EXLXhP+CoF308nOwN8gb5ON9eN8Dj3YEkuSOwS/mdn95Inx
Yg5PbREqpE/HiVyIH/mMg/mfVeIsqmuxP/DSqtAvZ0fCTVsJvHBQC5aTOkQ86YsE
oCdLILH3al+zCIsGto5275q1SnTtVwGMfcnCOkrsg2W3wPDdpvtZe17cj5beK4Rd
G1DMppSaLlKfqbNlvUHMi/h9OPhjkL1Jfl5qQp7X+2Byn8hDx8Yqx5JSX5bg2VMW
MBHIR9u6fjme9g0Bpc3EEA7c1XCkhiP5j43/aAewLcCVX6hPxDcV0QfPp1m6T1yD
IvxpRM91nz+WXualvYI74kiVkNOpSlLWwFvJ3Up59Y9DpWZpmOV0Z6PsOmgUDNfC
Bol3NhCqF64PsC3Q3TxAuRBBx5XSrgkoE0QDe0oUm95XnmPImV4ntdSjwJ07kDcF
2tGrWL6/sUZZjzWEALhdhkmFzWbFsLptkv2Z7A7WsokxXhPMzbw1VR42yovyOPPA
jQvFwpUXw+aN+PZvcn5gHET3qfkTqAvmEApQowCZQ9AvWDp6kmMmy7RQ/R6LBEyk
3VbObEGgTpY0VZOit+S2u+0NS36kG35Y4gMW3RqhNXTednzFYAK9ocSt2czKTE6x
kYQQJDDotJzlgBm3GOhZhKu/5wyTfw1NMJmM4djTQ6+qiuPG+02GV9LyhkiqngcU
zwujltyIFy5FT7d+R3BfIbZyB4s9yhXTWv49wBDa4x3LUFx2d8hYKtLXrqQQr50M
EY0vMM2ositnEZvUdmMuijYtScqhI+v60+7xDvUz/hc+6EVRuSu4pSooAErnYgLy
5eAANAyIsZp/wobD4+EXq42A9KG4Z2AqUru0ExYf0Sd/40m0NIVaEYV4eRLDT6Pe
6ft+kcKvHXXXfZO+VYG4QBaBGxKQHm6BzzGR7sG6SLBnfJDoRk6CWd2TFPbLbk1h
3517ZA4MvoowxhwoQejzh+VKFzVoJOWLR25cz7cpzTepeszbmoQY4hvnBCFHowDz
5YIZeXG9CZ44QcQ5lDgHbsdQwxhDQgYjO8FAdY6v935wPxSwegVylPswhV8rkzYm
j2WiPJCZqmMOp/BRDeSHuzyt4aICPWKA1tZCFAwgVhxEyTcsqQcYiHCBHAVnOcd+
Rippi2ExocrxE5RSNXnaDMtQ8h4ycpqSBc2Hll/6RVGbqhx0Cd2YFOPTsZkzP0Ln
bzsVIGm78tN/WTfBoGN1CaEDwjs/bblyztKA9Zg2m5dAGFxMQV/E7PLYxLl2tWp8
33RvCyEq3YTULL9ujwtoO9nBo/Zi6hCfGmbdrVgc3/wghgm3p5JPxXhrr9PO0JTs
kjirR9FhIfJ4sBbUZ294Jr+gdQSfJsHQ5+YnikAjxc7gaCBmQiaCFHnuqlqe8fF8
Os6W/otDMzh0fBc82wsSy+TZk8/I/H55UTzJ7d6apJTYXza89aLPigdJrqVQRBOv
mky8rtln3UCTyEjWWVV0m+nl3itFcQ9YcxOYEfjfaRXUYa4FGbkQ5JifNRfFy+GW
n3TKb/Xc6xLzQ23aa7OEGW9iuB74LYh2c8AEwLKY3TERxMWeFUqmIx4uoN4BL6IE
5Hwj+BhhtVeuZ9T4SChtzzkh9Csb6/VAEQuwNBXeTSUAiN7yePfSnvR2x0B+BnTl
6SSEnF8W0NfOVJZNYUC6YdzZTeI+acJNUL5vNAuY7K8t5zjO6syyese/8ekduSoC
gJmvGTiO4eCrHX1q8tnT+EtP8+QwrV3A8uiuyH81cuqHA1uJ6giTKuwrR1EbiEFM
GCL0cuMOaHgEipCjvr7EL6UyX/6U1kWFQqpib5jVhWt9VYtlzmfK2eF1WeVvG5vR
AUb1iR3pzrMW7ecN79Ou5x2mjNVaBWU8tNoBxXLelL+KvRcWhPA6g4PuywYEyggU
wAetfHT4JCqvzwAeX7rzyIILYN1htX0IiCN1lyJ2UweuNrupg7dTw3ZqI4IB4Teu
KTAPgNciM+qeuTj4xueJCeEhVBM5Y0wm6ToSlW/vy/3ZW97h+5v5i/tjIOtFTdPN
UcshrwljbaDDBHRu7wHyfdUG2Mcow9txna3Kv8hHx2ShG4/D0EXYtWE21G64jAIn
cENfeKCLVyXaZ7G0YBhf/B5a7kaTe2QdFicTOuNWQ2K+PPWixsabY5rN0yFA3sCM
L5/J0SeOE9XMN7IprDN5iNimFD2wer9+7DOPxivmQOpM71cD4vHWXG3H2zwKR5e/
pv7K5Ngw47UTx/BIja9lberzQ7ExlbbcbvnS2tvl/I+BfmWjNZpnS3GmlICOHhfe
tZUVM8AGuSUL8ifA+8D141TisLIamcAubtrZjF0F0K7hUORGCVAY9WhjQmC4/N/D
dULpPNzMlUGTCWebNA0Ht+aNPUiGcgwHQsJS5KoKG1IQm6JbUZqYgq5qgiEKhPMI
TMxFnnezPY6Bj2HKhIBEhKuhh4wafPSInJY0l8CnssuaVwQfW+g8eatT7LGl8R9U
vUAIVpSLDh2nxe00mUMUxFlgzmIz/2hjvxj9dX39e+OWCq7BSaN75OaxLKV8ZXab
YhwU1wM2riK3dluOQsgF/XOTafQZq4TxaFsAKw/sVFn500PKdm0yW4fN6nWvGl+Y
kEVgex1C5GypWemDHWCkLKnni5bvRrX6MS3vXk2M+q771m7Ux69fUoe1I4DRdVbW
GnF7kUMpRVoou+Ct4LTyzDxZEp4qdObT1Z2TdDvr9xxgJmlNpaONCM3jxo5VEScl
cxrP4KXqC4kBt/eMnF9mpBxgZEm5StBhS7HcVd4kIKLMf3rVzJ/kiNn4XWMVgY+s
7EWJfeKwEjLWeswMRjoPINHh9bgzyhfPLTusPByFurVjdV20VgcCBlczkFGkPOP9
itV/jsyXIdaC21kho9DjKsdNy576oXeXl3MC7sfNe3gE7ZhG7/tITjwUo7LSsWJh
m3HpyGuRRN7NW0qfxDpzhMY+l+D7vE2qDabwTazESajz3XkuoDzAjYAJdyU1+TPS
qvYzj6+5pa9yY8ladXH2MEkGke127/lsmzLPxTHKF7qjT/Ji0WU950LLf6w9LMAN
WQrHXTwswFxnDxavTwKm2n2F7SsR1lqkS2igJql9rR8qwOGg2hE4im4smYFjMeiI
a3oUrZBYnrGo5LKwC9dhknVytJkraIH/hhdCm6nhVLfKgOvR95hS4QKRvS/4YAmW
Quu5jttBCUu+HjdkWha1j+kegx0PoVg6Yru69QCJYES1zVF6Xzcv+bBMg2CNjj/9
h7RPu4H0op5aJ5SGAeSheLeryeHy6eTP3pqfFEze4S52KSrLAm7L/eBcC4tkjdA2
QkAjHJMAkefVf36MT4HdY/MK11KvJoF7N4DmVTdVNqk9BSk84UI6uXoimT15eeu9
pApdnZeuXrSpGXOf2C5tNzT2AgXUPdl/wzCrNwLcwtRQcMIaI1zdVdhJYXq040EU
y53C6Hp1D7E+R6XdzJwwqpKdjhrSPFie6WQdHeXfmzT7dVW4VQfMcN2TlfdXJzZK
u6FybATvhj33sCUvNKaH6s93yCOGogLNdfZKcLVSaCczK+6JcLLOQjQMRC46ndf5
oYnVKd3+2+9AKJWibwyztuwScOfN2SGjeKT/vlxwe0iz2W0++0GvaIMDghiRuG34
3OkFyrn/TeB2+ZAmi+60Pa1a2Tgv9HcM8w4Y9lO6aqrVMuGNnLUHnbgqyTKbP9iJ
gg8sYyxF5KENKjsfOURWUmrIuNK6XHHjDSkHOF0vte/xskSl6GRrHIhkPvr1684h
X+tscg3vtowUKwb1S/fuGqoJ5m4GsCvhOKArRJAFLqLWXf3iFB2OR3o5T14HmSBY
gxeoHTuZgOE8Qw6VXOY0+TolS8VItiy+HVbvvDt/2OL4x/+kPgVnwZtlRn83FZEa
Wu3qrUj39PSQjo3AF1ruUSohbmJRbMyn6TYnSQPdoMEDeShAsTQZ0FtDymy7eQsC
Es4mWcSYKc3RLkMQ7raN1F8iG0DKeUwfqpsVEBOhnHL8miVwgggNxz9NV8ToO32e
jtHQW/u+GGTTRbq0MAPPBySNWe3EXbcvHHEYKkGAarh6MY1bGeLha36zxqRYb5H4
ApT7yu/QPsluAmXu3/f0JE0Q1z5t1nbiOx1n0AXAM4MPvws4pqbmRb5NnnBSnBG4
iEilfX9xPvXems8kPQEM+i0ggpkt8rh1wiC5JSt2UgN4jfAiRIp5n9akS3Yy8coI
GY/PNRs94A4N59OkUwi0i/E3epjl2BmfKSt0Njjhb4KhFoGWcWHNgoAQK5YYDylb
XlBxOLGUmzWg8j9k9smSoEXCvOpp6WA9OgM6aQ5zJX7qZWyGFp327K+pBdMU7i3B
xTi4Ns60+kL0j2CujztSoXoN6j66Hps22U5a7uS3ShcvWcBoNOQZdYVuyN7Dg7xT
vbsZXpU6pL/+hSF3/CxCFbyduRh4y1MegtEKJFvYuGWCjbdmWC+PFkoIXFgXspMJ
1bdvM2bBtu9ueg8ei7OmlYDKgKe8UejoUvjv6etv+3BNrLVgawEUZDmkjQ4FwBI9
FM3hIzbieLIgZXfSRb6/h3yo/KRc0kodITNI298wN73LkRerFpBG+CpuO7m6tKZj
pAnNYUai44Rhe6OBWsHp2nxfHhcxlkdU2KzkyRoqtoeKn9s1LcR2guTYe8X0uTs2
kzcHaicZ9dk6EaREY5MIvG+IwCMugVuu7VLRTcG/h563q5G2I0mDyzQrF/gMycG2
HGVOjt5gtVCrwpFyP756F80Lv775UGBpN+qRSxWV312vtRe8kRq4C4pMGhRyTvIf
TFw552mM0wWlqmM3NqKVmRzJVTtg64vcsrC90aKJYx2/BRbmOgGa7TkQ5pJ4Yp4r
dqFnNimYKjk+zauXaCFlUM6fdpmdbBULuU8xfIaVPH7SqE+qraWxQCHVUbl9d2mN
MXDwThek/oIXbFT8l683HTcy+/ShUbJOCHJvhM4Z+ep1teysTAtgFGcl/X2iXN9y
z2HZlE8BtC9yA6hkLrPwJzqhHHvHvKhKWo3j5fbajf/fknkqutCQDxKCJkZQ/NkI
5uaplpZSgxSN3Oy7Npw8dviJrwLLAz1htMF00IKdAiN6b4GzGr4qFxhX1sVKG27m
79sXzMY8ErWMZs48Kym+/aIqwXD7I6zf0fCH3zwq9NFNyOFBmBpB1E4fX4DTJ2k7
Pu+iH0apI+IuuidYwAenKhtpljMtUWR8jK8WFr4qCpxhQCSX0EmuXSpoOWRyxkaT
gQXjwSmYsbVxWmgwBdP3riUsd3bXe1YDhVYGFRjUX6wMFlPJfmkqVzkjJ2O5un0K
pHX7Tm7k4iaBeIA5sGkmVaoEnMSlGA1qCawgAECI9jgQdydwWCKbreaQ2H2aAmtf
8ZQlYJsCCY6YIoIOOjMKsi9vvDf2iFII28jE6M8GACpz2mFPd5o22uzglJ1Wftvw
lnbfJfdUKxlTC6MeLVkDPqZ7lUuB6Q4l4SZNV4Ny9j5KsqTNcHSCpC3Mw70FZSHM
ISnu9zzKqE0t/FGI/BLGa/4AB1b+1cQHB0OSQ2/KaRTzTK5tLMDyQLOFW4mRKAKk
QwhX7e0X1xMJxgqbSkvhvZOf6yLqAGHMwdcv9uvJxF8FG2jWMlVIootFKwo8uiwW
Ds6CaYCIgyVLSNvMko+baI4Qg4Mvr6HY0DmGw4KhD7hZvhhQK7qHCrfE1DBKdMce
dcChOVoI0Gha50uLZgy3TG4XLGzs0G6/ctrxveACS2FsO3SKax+y0yj5UEoz5J6T
qzffAR3IkQrV4NlVHiMGYsDGm5PV2FSKDuS4UDQRiB/sBWxMHEJfSUHr0aEi8qeS
th/v6GNy5YAueh8gHw4w7y+GtqFuISSlfz5MMjX/A0GzUalxhUjfjx3JSFRr0+RO
1rDFEykKUnezBmyjtgcYRRcM9pevOecnGgNXoGiNLTWu871xobPjXvA0c41Ar2TA
GZvxqxRregE4rpf/GC5dO5a2f/MoU97yBC9Ab/Mi2JLkFcfifHuWmvZF5gEUGx3b
I7yekV/nXgAPxIFnl+6I8YVEvhfWDCNCfpMofsegL30ptwXS1SqTwiNvZ3+wdOyz
oIE2jaxTxF1cYz16wo48QDgIs1B/F7yu8SYcaZ+QQ5z6pR/SRw9T3ijwAQ1RWsuR
XFvhbZSHJmcayOjhxRC4NF2eSOD+RFWlwP0FLiKfbH+lpGlxUfHJEBn+eaINnQ7u
m6uZlj42trkUG4F+Z2H3cNwXYn9WYgqaNyPWOUKa2BwxIeIyFuYfcwjYgnUq6j/6
AB+uUngaPnanb4DRMhDZtQ01FWbQvnxcpXw4tF2yyOYK6Lole/6c+QuTe84mm6Bg
6647GVNHF5lGDRN0/UxK3eOm/9jPS/R2H4NzHKbepzHaJNvw/i8eLRmPARfV+Yks
D7VE6xvKuoxcdywBL+RGjF7be9k+WI+uFwcKPZoF0QoIwy/vNMGf9Y5z7RfB08hs
Bjmx8X34seqosTxGfr/FaOFLYFTk2h28YlxTCmqh30Fnh+JYml20LojD9bY43YAj
mBhucD5SmaKdN5C0YXkA9AvbDKMOc+OHzLlSYjImkgdBTDO3RV+XAv7QjUsfcczm
CgJOPVZiLbhmFKplztF4jnyj1KVNxAFqrxNdswx+JUad4hxqLmKirLWGhAmRgusK
ipwRCbKCFd8H1qSkPhd+tkYCiUZUZHOOWXdT4/BMm8eQff8Vyc8R8r/1qiG1nDXN
h/m3FFn8o+PoInWEHuUBbo65SkPqyxWbghI/aihEdLs6v/JSrqqsI9+7pnCORR7W
MaqQzc3Efvn81dIKffur5bgrAth5k8pX/GMjiZwpEXgNe5JyzrfFeSbzUyQwh8Ah
MzDxtc7vondkizeLxseIefkfPa8ztsyoqGRVQusGnOc03D+YuN6RbGWVB0hmhh3q
CJz+TSHqJmLm1BuyxTcgB/6jzuoEAKxfUWz7LW0TbCAfxDAmi/T1fXeKUpophg+L
1viMxUIw3L2h/z+rCFWMj/twL5XaPUou2nbudlTqIIsjiWjOGdoE4eWHJP5Yox2v
mEagJp7sA5a3KkHK0GCEGGGyRcaukSS/mOMTiUq2QipcBNLDODZfrmebT8OrRJYX
4kz9SIQ+DypfcCg6q5VgMNqPD8V98sNqMsNwCSn6MKtxrX7iKR7eJcb+5DWLJrYk
DNLzVMtW23VTDD/WIEQ9u2NGlIxeCo4VzD7otxhTRGRQB3XTVmh/8UbPXx06XD/G
2H8Gczu/73xPSSyuaWPsiJdzQcEZdkq9rziSopv/vZ4kEuYyBOgeblzI+CLrOp8v
ykER1ENmlU1KDBX5NGcfkXY3K0MewgMCNshvoAvQOC+IbS6nfTMS39yklMVTvsnm
ZIvIktCIh0wYw9JvMqKbUaO0ji2OLfBE9fKwvjAunFd++Y+SPVCwUvhXm9IugdKh
kWC8KGCOUQN4FkIGi38baA60XE5leCw7Pg20GPqU0s6bKo3TqPmVzk11KhwY3owm
nPOO3XI1Ji74vnWDhOcvUoeKYbe4IpIL2RN6mZR3WHLkotYvTrKleFJpVqR/g8Ls
7TGI9HyU8Urskpg1i+qLpU21Ii69X9OMSrMKXqtll1oHdwS8ntA2WH+S6zrPyTvv
jX7J6nodj5chH0Qrsibv8KxwSM/k2wWUVIqiXvegtKK1S6jEjG04U3fWAc3Rs9q0
0bKL/jYGjD9Fahdcle06lS1/EX/hUq1o5ibevY12G9jo47OPbtWLJMjz0sydtqON
8Nfp0u9c+vPR/movM7kWvWZ1nH5PlVvIghm+PagaYveVP4kkQKLDBeaWixPYr4BT
ufaeeLBKZD8Xjw4u/j1bLi4MYSCtIDQCUG3Ddv3CTTvnXR2tx5nz/qPrnnSSai5c
SxSUvte2s49m2wDjpQiQgleDEk1udRs+r1coGHZV1zJ1cdKrwy0TYQjdK5xqS5qD
+TYRasJUFuH72E0TVtp/Jzu2KnlOXJNXkFVXfewmp4gvnlDan5Fkiy+nFAB5vHcj
G63Y1U8uPVKStdqlZmJaR+CF4D3fT5jH5dwt0Q8KX5KvMQ89u5w0uQqvSGEkkRgo
QR7GiYdGhfWc847FVhAUMtvzhQzCDgk3dHlGColSpLiLGns+kI+l49Qfy1+HfkP1
3I0JkDdQ99ClsbpwRZDW0/EEDLg+NgRDxKtCh/iwiArUpDeAeHXVk7AKzI+5n+Vc
5CgxLirie+IDrLzny9IoJrpWdtZmFlk3nLKNWP1GGcmWbwlv6J2T0OWfsspaghTd
gNvioGNp8vs47hC1vX9bgVHjMFiNSoFLRKhuRxIoFuy9S/ez3MhBL0Lcw0EBd+Hr
nGEobT8SlGDjOkjRhWm6KULmpht8APRZLmkQgQ+wrUVDeaaBCZutHmGcUh4MdHbp
ABe9BjJ8i6dwdhoiIl/8aeoVH8F5xSbwKMvU1toJ/BA0/Aoa8aSmICBowrbC0nak
x/CMi4xCta0FTgsnmH03Hr+S4KlMOLbCrd/yxX+qkZNJYRRUqoz2wY1y6yRF22AR
kOr3LeHV0TOdo2Huk2a+Z75IbGsiIVhotrPUniDg+88Kl+wH6pe9Gz9WjWDDzgE3
oDuORBMBZzh2Bb/C3V7+cIeNHd7qx97Fozxj5HZpFY8mhlHvrRN+LLPfFLIbnsDX
p7I1CNRbJFNRDbYYDotXJLzliLmyPmbSIHPJDIa0JbUaOZkZEr7nyB1l/PpT5sA+
ixfZIxNKCuwW3J/M7fvAx1KBp/+K6FOym+H3qz2+Q1EIz5nJIFoTDAIn4sqpitd4
ikR2o/d77a7cQQazy9Jr5qB9hxZW8/nMm5DZPxZtR4op1tq3/7YehYZ13PEYll8c
pt8V4Blw18Vyb1XB6ytyJx1LQnL361CE+h+hPrltPbS3zk7gwQ8yc1/QNMkYupJk
jRHmcLGiDfqx43K5OCswSFQVEgAzEitVirnOEz3y2tfxkSAnohQqPX+4eHpmQ2rc
1NLtDGlKCyanNZLic0sDnOWZLujZE32vmnhJEv8aPuxCgm3KlU0RL8OULZtRqRzA
FU8QpJ43LgxjVnLRsjdb9DPCAklgYUwFtYhrWlwhS3WxhJudF6VYvHAZLi9YPg/O
dGpLRFzLwpr5N4XPhALjD55EEwdUiD1w7CXocF7b9kUWaO8wT6l2K/oDzgicFFW/
aHGa2o0ylUpK+0xjLUlYHG75xAl47TodVJnI+pHkFA3rDZ7N9v+uFgKrtAI6IJ1e
7TilvbeIG8s2Gh2KALpaytuUVMh0tZdm9hsPCbCkTrbRfUTHFNH5eX/3dyZXt1iv
e06xJtlVbijeEwTttt4SaebF0jVN20WKcNBq8NIpCwOSnh67AVN90E3amxSKJN10
UclCXm/Gr42HbTwp0suVc2VxmaYLWRuoUdU8c7OuAVkSCfWLCQHrhRTDat5AuBFt
52q7o9H7sB9+O+XZUlrVYi1VREDmFHaHr+jK1CXGwJ6IKi2xHKmRjSqaFwWOpTBC
rY8ft6gRcAAJ+lmf0fRsKmlcKR96waexgPV+QD6tpNnOGLmKkEHB7u6MnQnk+0+1
qAUyXUAjEL4xmn2VYVdGpaD2ODi57rxVz0ji1qa7P4Q93d6IX8yGT5mZC7RueUZa
cLfcvcIEJQ8yABgDa4puy2U1K/T0HVUkC8/C0HxynAszAjqUmc20G3B+Iwv4ZXRR
+VlzBF1macKXmniaL24Xk1c3WtmWoW//3x+fp2D9/3aMy+eUMNYiWBzuW03ilSZ4
Ae76lEsgSjpAkzhljgflKkgP5y2PIFsBy0oNrThSTF+LleKxWfmjD7HAp1MYT1yI
BQZT9aQcVMOPVe/iAu9zJ7dRTxx1mdLqAeWQgqlJ9XV/jnykEnC0yG9s8kQWCIsA
6zgqojdR9+RqN0z4SzHTWRW7ni+5GVOdTGL9PFpY0Dd6fo+G5s2EZmII3bJl+MUo
CqgkZVoy3Ev83K0k8p4Q0WZbPvff32Yji4LR4pO7bkPnSqiiets2KVrueiGjboEW
y4osm5il6YoWtAmXR6QgrFIaXFGba7BQHlAiyM8QV5VOJXT2yjvA6h2S8fkNhH3X
tIaniRPNA+VD+Fopv3mLCL3XXXLHIwfBkTb73dZBvBBZWuI24bXG7NFltmvHm+RF
J6PgYfPxFWk69F5P/n+DOje+m3stTiZPXrpOJHHvjJSz/D0ZA8IeCPBHBlgbFMDh
dIZsBgWoRJL8Hj/8EUkc0jVTxtGezZJLDcEd/dLWfUkvPDsiv2m1G6tvxIYHeX5e
F6MHvIiouXYl23vm81WvaMb6uZWGtnqPYyLYm5wSAdY1C2PhPE6OUSRyUist0VnY
KOBI3I6R39sfLO+lLRcCwZmKqWFnPVUNKspN6sCChGucqsVPgeIKPdjnCgDvacdN
uwy6sxW2GJTu8Sv0HMB9mgFFP0kGYU6YGCVoVxJ4vWqCbLHTlcdFtprWD/XXdMN7
ct0Qz9tED/Z3XkmmlKLQ7q3IezB24BRFtxVaSVJp4VFsogCtvG7FHFP3v9AGT94y
EwJ89aP0A9ppgssUaF3PodoG76KRh8dFFrccskTIUqowGMFJJnhMtACHhi00B11r
c0w8FICvr5z2LOdP69XY9Z0AzGQXlxZs8ILBZFKN6Pvf7krNRAPndP8rIWYOZzbt
PVvacYWaXGiWcabLV0XpTUy9L+GU6hWpPT6ANpt7sACzIinRGhyi/OJMcQOpNKe4
rXrsa9h3SJpkGCu54gmBERhdS+RIjovfLgNSqj4Lq27goAeFOwFuqceB8mhohEQA
ME27MWJzIatzbl9WzRxBJlRcYQKMlv1q35m1IuATAjxrmDa+4YMR2p3SMTTJaWYA
2jHieeHInquML5cZtE0KmCWUfv4Oymli018CoD3fkrAMbuMSOcegrdW8QuMA4eER
ajjqFowMKVbf/K9eCUi/gwImCEoEIRhBzJJ9UZt6qIdc5Hfws2mDIjYeU5JuXwQz
PkXID3oQWI0I3n8FKf3ZPQbL40+phjdfCQ7vZQBMxrabzrWXna7SUlitxNzzMfqj
8s56Ej7dpz8viqTOqwdoWBP1Ypc+11XG5Az34lQ8Hwi8wy0vRa/BF1CDWJgHjfV+
Com8TaQFARl53b9gkOJAedyf6r29Drzj28avdXTUNsecOWykK9hktrtKqRIZwHgN
XxuOzSSv2fMrvHLlyaGUwGFEE6/Fv6z8DLCedCynk950MOBqfYfwl4bkNzyNtgJq
YtrlZ5m66N4KWJZOYI9nWqidFr8Tm1yHoy6k63dgUpahLWfALHrm7d2yfKhLtMGf
GVpD7L2BzB0rhSQFj9kI9uGCLsmacC6PHa3od5CVf/vyixZImUFEugQLuC6XDFOf
zB2QGa4VvQJDQ7lPUhZeYNI+0qxpdL+Nv1iUilHAUPYSOkLBpNBfYloeSL7+NZ/m
MRkqnlMMY7bj8P1FCgMrV4RY9ZpEbe1ya6pd/lBXN+DwrmfWIZFW+DKoFbcthNJV
GMeHD5O/BHxJm2Sd4dMRWb1k6QbReh+sji2hnqmgu6b9iksE4MSIdwtIoBs4yFYu
4uCL0O6/0kap8iUzWzPqHwxbxNH+VaYx/H9CrBac5h15qUzeSrME61kAg5C148Xi
jAo32SAg8/hsBwzMwglZH3C6xE5EBsGiHm4yQ6v+cs5XVCMqBm1YDVf9NrkVvw1W
lIfk944fZ6dInMpRk9z/o+VL6dKYfe1w6MuPWVHNiFSmDLoyK+05LyDCdH30+eDO
hamOXnNgARgxPAorw0cIqNjSap2VTr0VUmhaoLhz51i0sCeBuRHMJnZPMUMEvwV3
9kSHQUllcQVoDgQh7J9HQT7QqZ89etCcboxgowPcLeM8nhlMPfXghRauKF3k2zVv
4FuO5FTNNPGLjcS921jeBvIrYDAFT0vob/8u3mEIwYoFqb+qVqS2KghqaRmoRYUG
hD9JDagZp88DQfxef0UmGdih/CGNpvMAkAh20vZ4JiuGUqpOORtQBl8hoIAatSJc
3t9tRZ5dJlt1VvorA5opFg9aWrUZ/sEplX+bZS9ln7FLRBhbCrZs0qMPiThyP4JY
apVoWxqBMJpa2pfDKs4F9J1GjQgvKZmqT4ll157Y7ypuk8hFZ63K4eWQDwoaLjJw
MLsLwL1SJxjPWkCY4Wipbha2CiGDEW1iGYvWuMV1Bjcz9ZdcCgMRUI7s1VpcxtK2
NlgCjXWd+jDNdyS8RtD+CAc0/Ea1dARJkJNOaHd4krMM8pVqmpazQ52+6aHKWoKI
i4B6gbpG21nfF0CccVqgh46apEZ2pKrgIyTG5yAAFcW00FuflwK1MkulT0C0YkoZ
wAxWcRKUtvkb3I80ECP1EPz6pffYW4k1VOBDzZ7M38wWZl2DX4va/2EIwzeC8EgK
fEWcsMcfWyQtYIOvVaboY/faj6vey8acmPxpsaEO4YCU2ZfBMMfIUS4tDidSWVei
UrQg8IVJc3LLYtm0xqRv+pIn+Ari3AD/WkPrBVifUJQ4qOgv09L/r9sXqU+UT1PY
GEAXtXCWBW2KbRzZ2hMz7nK9hxFl7VVmsYur+vQPPG1yvBfiiRTh1QiRiDD5+X2w
715vnDZYRxbKKJFF8/yzN4D08bRDbhj4JylsxiEo0Js7KFxwaXPK4dKXj6Iygund
Za6CNFb9vRoRd+zFTeQmQy6Gi3C91Y/T06DWQ2MjwVDofK2D4UpeKDUpQBP9gedr
eQsvzHR3NI3Xa60wKjsR5tpE89sur7k9bqUhJdeJmSQGJfzWVbPpp3Zl4cOhmYUd
ECvycDxUqvSYYZm2SbrdV/IKz0WRdCwUBW64Ymy5Wls3RmCKE6tFxdYuc4TIN01L
fXHfSnt9TcGIWxl17VQ9cH/eCYBe8b6590s19q3yReyglcQh0XzbYZuTyJ7GicyS
B3rgh93m1xAci2Ew52XBXIPDzCl5t7o4ld5aPwbQ5B6PZ2mPHd1cooqjlZf4awkG
JkR11F2t5H63+yd3Woxa3JkqIUiwmj5fqWK7y3onR54BAg0hXh2dKA3ZoNUPconG
sLnsmmibZZcMe0sZNnGUyu53C3zua9koJDC/N/uu6l0nqSFKVBP7wNOC6JL3JUFi
74ZYx0l5b80zO8o69zIjhGEEmhZE7Edp1uIjuXjfwgkV2ZlSym3SSZWRuonMtUVC
wvYE8PBkz4VaUGJvK39BspTuo83BV6889j4s8Q3Tcro75rfwS2sUQrhjUBfTpo1w
nM4YO6OMW4wjVHfDndyWs/bAcbaTmWzFrD5vy2WauNRpYa1nlXJtiLAKvWf03vcx
+DalY9jcW5UpgPNUGyUnDEHgnmQ+nsWn50toHuhg/Z5KbQTtJKM5piHIF9C6DKE/
64ytdeAyizkFdfPvaVj+5d1A/HoarSnAKpKLyf0UBQlVA2tVSUvBeEX78HYVM4SK
Jg5vBvxOPbIXbRedJ8g0vyQSJlFY10pKT2ZHP0iN/WqcoHicTTMGxq91OpMUNze/
xGf8rVhED8A9O6x4miHYNTIGscOU9uzNI9pDkLoZ3UxYGLxaPwppH+ziS4Nx2cdC
FqdU0CdarrZRtA72cH8psDtGYpQzkDvlf7dEAOkK5GAFn+658Du/uslHf0Qnuui5
iyWnmZpp/tG0cgvE6URyXWcTWh9SovGVj48lwskO6Mjm03GNr9OYjoOxkUot8/ZH
m6lrIPh77uRJgMh4q749Sxk6gxIP581B+9ZrWfStd5N9XsYFDgEb/EcsCb67KjA5
guqQJUFJGX996j6cQSw8tWacEfRbRUjTDd+N9KxuGMg2+ChAAvaJiirJK5t7YZ50
UzIXyaIkB8arQtOjjdlC5BhRDw7GhgmzwbyBHY9iVjVFleFUbf0cZf+03ymdckWh
epRVL44M6BSUImx//qwFV6rfF/xEgf/AMSJwiOmSIS2tUeNVcbzIEAdu/AsTQJpk
sAyUHBoUmoV92deulI1Sh2yBmx/a4tx0tj3pfTnzWxVdpqtKNe2k6RYoLiY+Yedr
YcmszFrYrxVf+xltqaaI9vd8XoWH1QimQoN1Lx2VFfdNnB7LvVJ3BHzERRZnr9r8
lsXeVL7SEDcDWBYETznPD/9Bio0UvlpCqvCsBj5rqCxn5Els51TSM7LoI6mxRj8i
oagJVYPs4ccF+oL92fWabs6mZIIwCAT5klru3ctq4bKlJ8kN5LDfLqcn5atiLxN+
WMQyD/wNXrmJYFwoIkSE1dRLPOGElUSB728kIqb2/LBWvv7tH+0BUCxsy9ZpFIS9
Dx2aa8aMn/40mQ7IPpl3QyRcb0+Ud+QHo9XqUZM8WarFaTUP2BPN6Tsqnn0xxIS1
Ae0absLe5yI5TQqtW0l+vgNd0VVHd3eUh4NtDF5eQIv4q6fYVjihVb6iAD2qjmkw
2/uJYmBQU1WKtx9e6dVa1DJhqfOU3kgZ77vs8mqIrV5XHQoYm8RqWUwILSxo+6SP
IpFRADgFK/peB3QWftslxkTFlsL7JXYheC1Ge1JKAom3iL0BVb7ed+xLtMWfblEM
r8nHLpZUuXtjGSRhL/ZuCYDrUMgERBmHLZaWTWeKFXFr7mg8W8rUgNKsOHpQygDN
qp1oa/nlBeETIkXQvkjcSLBNQ/sxDkT5iOiwo7j3kw1j4biyYu49EzFiB5KVleBa
HYL4MhfBmw1AizTf+BPdjs5aqkdlRlUBQJk1EVO+X1I4vBeDWF+NhEZ5DF5vpfvY
y/RB92P3Hi6gf18w+LAUu7LO5oS0kAEeS+zUTv6nlhBhp4EkeiByAgRXhr5k4Klg
bCO2dCqd3VqAFcKYurEbd62BXt2hONdsbEQORx+Va3GetK1par5rWRqvlrPEz/ji
9tHbcHvG48/G4gRPoKh8xxtCUEGarjvKfONcToSbfwMjlccmQiXbug0Lukc7GyR1
ZgU/gNiRZTMBfcbT98NlPcRUUj6tScfJm7MenmcukSk8EMNDYN7ib3FTtigXokIs
gntF9P4OFxckWFSJUQYtpGbP/1VsusCQLNLgj6I6pGsoZBolCCCjFmT2F3k/29Ef
LxA22nmy26msgdALxuYjdVIRAqHNbO8FWYHV86EZ9rrhVgplD1BVFLh52AM4gFcg
kReIUbOnS77mGhjMDBhiVdpsmi8HabSq1kAuZL0Xr9E2ewjge2R8eEkqrqr+Bigd
EjeM/hKKrYd7QoVqLRN8+n4MYmVBKV4p0G7z6RUy96ajn4mZDUzcR/oazdUgNiTI
U//iPBNxmRC/DeEzHUR6VPpx2Hb3lHCNPSS4UzoUTsar2UwGuDF7yXxhqjbV0FYo
DUErnXGh5u1KsHdu2vaUHLu4xegvz/bqTkYo0TFPV5Unu7iFIgPEKRtUqA6XNabi
8kUQKs5mbBN+YDo9ad+vXrTG+aoS7O39c4L95ydmkvpYhwBIkSuygQYZBMhgC1cz
3aeka4EtSXtDKHcGKzzrMC+ExR7wX62wNPV10Wmn/X9jLMhM/r4OQjuQMIxIfR8x
1nvbKdret6OprQNV2Zx9p2kUCKsdYygSC1hH82H76ztvUcSfYBkAJzypoE8/vBBS
3E76CHpcgH3DJlC2HTW9SScdKT8rjNlUYBX90T6896D6piOLODLMG4I+rerIJG4L
pjPmU/OHuPwdnq65wM9eW0/7UZB8NntBfv5h5O95+4t0Do379E8be0Q9QssIN9Oo
ocZRpWMFndoNkyAjNUJPePaIr78rzxv3sbQ6bLhF34OQk1J1OQDhG6Y7Q9k5OQI0
Bn0gdnY68bymG6Zt1Tolxi7wlXidrqoSH5yn0N5yTkysqd56LG0z+4W0M8a8XFJx
9nalzmyUMzto8lh7LpcrBcnwdhJR/GKB6fmLXsBXQHWSdoJB+rvjChOVJ5qjXZYY
3Tj/dDQB2rxqsWdhgXqHSAiU5BZL0zKzvXj5pARxtHlRmTDigmOAapBNI77LHzjD
uiKKvRQ4X8utctPqSaQki9xGoImgFG3Y26/1wiZRvZBzOzkXKUZqdPCsv/urrsqW
qL9/bHt/V2SIaiYXEbjnks47lj7SMeay+3sP19HAdtAPQcLoTkwPMyigixgMH3YD
QGq+XPiTDCGsiOTSgfqRLY2xAtF3unXxYh8ZzUtQVb72RNs85K8TBNgOkn2QZ3R/
ZDpb6i+hIpY5iRMmyOcJR5Kv2DrG0w3mwWePvugxd4uVt7TpXPPdRYBMXUcKyzVH
6VUF8NrUp0UkJOfiQSboNIkJXQHpM0L6CxCxF/jaoo1qyAoVzSEVtS0Nhn6CWq1l
57tiwAMOCwfik1waLLg1jJQT1sc1vO3WKHc9lmstsGPxwu1bEfcZBf/bBw/nSGVj
8rl9mHK5gSSYcnYBSR5fC/+Y1jIVnJq2bbvzE81sH+jyOOVsmZ7aHegZH1dU0NUZ
zPXVf4kaUzLMD+ei+hxjfW1e4sWwi8d1PNsnr/i8LB9l8XoY4Ll+c4ThM9TBxdDa
9ZHPZHpvyV93thGSWjYtvOiiN82s2b7PXFEgB44DFJosmm6TD0/ObcT8dNlv3GPi
MdgaQm+S+PQ86zvPZVAamFoQpEVqMyCi71QKYYl9n17DsOHzpNyHct+OI0NptqWy
Nlqe78bFjcwHNJaQDjiSRL9g2UxvCTGkGfyMS15Y7PnxdgFVrGKouyY6XCPwk4Ht
lEVnPM/ZhOKk9lQab1K6dg0RCiejGO63a5f7pQzn/D1KHoD8vNMCAjtExWFszDNL
1QyONCy+VmxURohPDWEvC9Z0nyIBcVRN3cufcrHoTnAJ4zqc7G9JGHOFMnDdV4qw
5+4+RDvedkrmvDgWcHk9I7Ws3KK8roUxYhUQ7541aEbN7O9g7ZmUXUGCyZrrD/rE
EGjPCOoquWMyppnZKLdIcR7ANW7fqKI35yp0ftIPzz8OJonjcwqXjJ21t5Tz39vt
k+T7M51xjHxGOgSfyuAOp/M/0ywMxCGUrhwyx5dvCEeB4ks9FlOexIeA3OgEKT4Z
AKVwldllqA4dyF6kfYq1XovAczNq9Kguk7hIFjLNPLXZ67YF/IId+bsTGaWjoLiR
yJbPoo3O1S+8VSfQpwq9v8InDZUIM22659Dy/G7+DhtGLXbVgqwcJOM1M4U/nT/p
RwQnO2FfKqSDtOqaA2aVBhPsnPosxqS7F/dSU73hIhxcmDYjdTfz3TC8oUbfQAeh
eEXyIqL3j1zK51y/FQtmpB49SFIfremdhXNAnS8aRu0rZHmTztfoXTUX+9Wx5MIS
+/yql0vjuAqOQPI9wlMtMaJnoCiaG+JsajxWhlRwvxOUQETYEMZxHcnW1B9HsSxq
q5xiLyV3YZhpH+0iwu7WZwF8RFhKs8k2QYfYMpLVaCKVSc2UBsFFOuGn+cQ5PVyE
aRQT+Isywymu6ko+VCNkMyTfUucCUdvoR12HXBblcET/sWZ1ghBuX30L7brU50YO
d7GHMYnkRGFo+RWcpZi1twWIj0HnVeFfN3TX1R6vwBf9txegr8F9VP385sNFgtRX
LaRoFiUCg7oEaH2k4BzFdDIkgAdosdeSvDLiq52pfhqu37W/2mg7SEjucexBVfaF
p3shVZqvqclO1JOCTX+/AAvI9pzQs96SMMmfJ3PlGvIpROGlEyhjLxQSQE2AR2R0
v0Qk8aZkySyv2vn7C6GjPbYXtuXPZYnFrd3GX1BitzPpcK8zzMHotvUZDA9NXzBx
qPhJBMkvvUcGzXc/BFZRulE4QGqE8rfyt6pmt9purYyKHJC0Dv491R2203LcbDhr
ifL5bywiDqaI4X4/xUbTOore+xjFc82lvFbxs7zty9TFI2eU5yiktlgXJCcD1+rM
LyRfgaLVkvEl82O0ZqjLzGQtU2cfkLPVWRlQedTmxv5fPUJWU8TyL7rZXeRnc3Pu
LyyRSLktFgL900DdRhGrLgHp9xCB7Vf6gTVdAOME+qTYq5MGuajg0n3fCgg3Oqhg
mNCOO9uHtaqonkRAP98l1x9BbJb2ZzM3fBcnHQD/fw46z3UJ7iYCvI4D0FeOFikZ
2kimsvKnbllGQRjla/3RNigEmIrkEuc9+MfQdHZ6dpSDzM9JiYgpJu2UkQ2A4Up+
U66OWf2BbcY65YBQCMcPtoB0uNesM7bLjhzlxvA5s+AK6NC4mJ+PVUDRMOy5Ymjm
ZNLUnOOShkl7jF9lxtglwOzBmwQwB/Hh4/nh4hGZfAJJj8J2ECZc5x4/pIdudYOX
BGWBEtlgEBh798i5glmksHGZBssZjvxW8Ii7/FMK3TbuzhBGZMB35ywi7iDDchEb
yIIgzGNIwZGinZDs8xPw8jXw16WJJVhjhxIZjTAMBg4CiwuXL6UYbEAqVR9MC4h2
aDv1xohbBcAZAsA59y7Dm81778N7g2YpOeJYsjQrAdrfDcKrDncDzdsnguVwQKKA
Y30hoOnoGRBaRoVQR9wI6FOW7RGhSrJi2F3sI9n7BbYeY8S554Hnpq5sAKkZrT+K
hoXCanaOFLY890WsuiEKy2xZkaqcjT+/E43FXIVyP0b3kNiK4g8dGostIoRPhOcN
W8zRVEcJz/HK3hKsqDeq+HRA7QGs369LuVvehxw3e7FViBtnSG2CEm1PpLeZ15zO
TycKaPVShTItPfc3l8N2/6yX6b/gqQD1e3ZgKaGiVesQDKifUBDerJCuBBWj7Dy0
24AGndd+IeCSr+ytm1ujrPJxWeYQ6ghUMwGMxOSF+P6iizt3Cwoe9dUCtR6T62Af
CdcKv9fMfMqpjP2gtyoCWBcehTtgK2iD1hBuWLjtG+As5LygrcUiwONNcMmSZU9p
qMhHInY/3siquC09Ty2gFFoLyaQkgU357a8uGEwgRuUQE8xASqev1oTtedpgQXb/
vPmxoPyF1GAf8xfOG4LQqQybyMIBL/RAHOQTASioEPc1elNNETKR9dfmMyHP/6eM
pSXXx0viGrFnt6BAaRrYYZis6I4MPFhn+emW7TLXLPG5zCl3ksuUs1cdJTLvp2j8
pusBTeLWxlU5Tt0RXyrxeL6vMgObT/VqnA5D6HMEImk8WEw3lnoLPOV5FWa5gXcz
aEGIgBpXrK9noSHLVAkrEPO+k7vhIIjYN1nYcQl9eFNTKcK6gAlZbsWMWrw7Lla6
6vlFofeEARxHiVEXQ/i+6/v2gRozs/WnHwNTJ4FaEtj5wMf9MhQF383htBq7z+PU
n4QYZLjKaM9fKpHcIOv4Ujwynx6HeHfEpjQpm830WbjZ5do6MKvQNovqcSrCsFp/
+UAYoBr6Y8GRuA6+Fm3NaRc9whC6ai9o8f6wHAmfjznhyRZEXbOXxbkCHd8qIDRu
HeG2DMBJkHFiu8c26A8/8a91ba2Hlfr7QCktP9yNSgHHrHt7ppA0bY/pvR52d0iR
REBvT0qO7EqzaKc5Sc07vBGxcjkzdAiEWE7cuuXRg86AMvMLejf9pr954iU3+ojI
nNgq2UDH0VMFkHzWs+nAM6KBvPmdYvqo6Jatd1ZWBL2TL4tNHcp8FtGio7iL4dsm
wkzmZIYyJWR3ftcCQRw2AvcVRXfRXS6QbwCPqRK7K+xdjaF8LxIM5PlX0O1/XdzP
Qd/lvJUYtAWoLiBHYzH7WEYlubpoLEg7qtRf51FHSjjWSSx4e1kODNYDXAMl9niQ
VTDtgEdxEJ8NKUu+nD6x1CSeEmhJx1H6i+U44gjp+efyM+5oQ1wEtny1gUi9g3fx
5BVdS0mhqqZSOAUmDeIe0ZpNl/dIrOwbf4P9oQae1pPhCmwG6GiOmi/Q+mEaS2Je
WkJbsZ/N9JiL5skdWRG+ehOtMXI/vfs76PpOF3u/PNp1EhDWeX/iXimhLAoYhhkK
G3zV17oCHxkMIQiKLgrESBUGEpPjxwjVf7+IQgUBmumrgyOXEWPSWDKDNv6umBPQ
gNY+SF64h9aEgsXBFRFzKnRPb4eILFbInY0/cyzl3ZShc32nmM2647+WRFiAJL9B
BBq1dwPWXHGoFvIaH3HhQ9aWKCU5kP9YWoLLLnsluavNo5UuoV91JmH01AyPM+HI
BiqQjSaBNSxJTspWGXe8CGsWxlaYLM4RRaR4DWYARFaUX1T0Lw+IAajEPCZgOvcV
Ls8lWTs2V1fwusWyBIp507CyymPT2JvRdv12MjJdTBfcnBsbIzjambGYXAfynP/5
5Hhz/vHlb4AQxDSELGyyjehlj3BoTFetNFSQT1Or5wsvMAUyNbA0Lxy0dcxUXK0A
ODRZMZbKzx7ZsdUTlfJvmOVJ1ciQQCNlacWUwbQIdKC6Ox4jbYEi9on6DkUE7WBY
yOPplmcXjZCuAhQrSOOWbbvFUQvidqAxaO12N/wdA8FTS0YzkmShdYGucD97aK+y
kDb2irD9i/rQ3VUed8rVry9qI6kOwCzxFsM/DcmGBJUdd9oGSCeVCd3cmd4o5olB
eeSYBDC3R3o6iUe9cgwm1J/ahMV/wBmwnBUu3ykywt8A2iSy9KzK+qRVTABL+lvo
56H9ML+dpPhnm4OVHMBcPJ+2HaLFWsvHCIxIe0NJLVy+D47d0pjaEMIxYiuT/tA3
m8si34Z1mIVKKj43sOyNPsIEYiq5HZz/IgAI/qei7VlOEWJcNJKbT1LBUst0tNlD
VkWjOMoEROdFwCCHsKhFYwYzEkAyhzI2rAn+JB8XrDNjcLaY+iT61uYJtZ9E22Hu
hkyOlyS+nrwi2zo7R8A2k/MY0TvkfIZuZSDwFwIjGeEKHzAHh1IXdVFb7cbZrdyY
m1V2+wEABSKsu0h1UlSvksyBVoDuC0i3Gt7QxoYJKyXvxE4MiguaFNkMznzI1f9g
JBmP12sG8JxQBoGaeFWrDfLA1020ynQ2Mbs0cSXSHyRBkqOPLE9nooeOvBSWbS7I
XIzQCEyy8ldTZoC0WdPXS6ROpJM2NPLGSKvLilwwA3F+4jxeW76YyP2Z9ekC7WYw
iBh57ckvZbt3RWVqmJ7fNSC7g2xkcNGoGO0iTlRfyeFVpeuFnxUB2oX9Y1F7VOik
VRSfVHvr+QFr0NSV0m7iw36PKZ4KsCcSeIZiVEi9LFhXpKzK73m7LzCG41Nntzii
YZ7uAr6ExgEV0S9RWvrW9cQLMwsHaHUq9MiD8f9nfWyClI2RpPm/LzOUCa4pG16g
9clmdEH3GNFrHFt/K/BLHgiHRJSed75XZihmGsGmqXhuRyoID38wViQJ9MUfeaME
SjLw91kRTJACQKvMY/Bm8YeFRjCZY2KgsaynZ2Jk6Iabb6oHUK2s5NbTH6yay9oB
oqu0qe2IrGUA4MckNeANXKoFQE7R8AOyjz7qJqnUXm3UsbM4DDkli7SdI4ZJGL+B
i+ec4SPo4w4+OFTjR36I6VE/hckU+NquBXG0Y45HQ967Y6ug24j5JrWb2gOgJ8Mj
fXyQljXXjfAl0vWjL3BKZ1YGFdhaph12qI+KTXwFmjRR9QNk/ca4dVf0s0KR7mZl
pXl+XYI9w25jTwQvuZ8OB7d7lLPDosTHBrGrDeOF+mHwQNAeshZ34v5jE3Ug/+8E
0SeW1YHikUDi1qrzI0R6ZwlcvRY6FQATZisMRM5f7dJFoJDDQ/2e05Wv44YqfFSY
Z43ql1VnX1Pp9kJvDETK9VBX9OjnmMMEeJu2aTkVLL65wH1l9V30avfYH+FcI4X/
ED0dGgLiItrHytGIYEYBS12+D8tQsyYAO4qga6PRF4yix9uOP8+XEx5R6gW/ErJk
qZnSFXTeyNwiekhD4rpnWLZMG4+ohtCxGU2Qr2eifLRxc3KjoIyAssqUSDb82yln
Y9NNTZUx4/6ImTDGeciz8OcaQYt1Ulsaaq7Kp3CaIGzSLwPbp703a83y9FcU2QbX
r1GOixMsl9wOSNH/bSNNWkCgzPm1NpfJH3Gru0wVwzzBgPKp5n6sAqtqWrVmWC+2
EfMedirDXqSO12uof+wyLa6gsl7b4yeNDybMt8ST4hem2wiPNtSjW8HqnLEKNKeb
sawxM88CHCtLd19f/W/wFbi1oyje5JJk1IsQ5zIaNS8RAeaMaZELhJJ7ffxm3IEI
d+GLMvxQAg76hlrbgSV9EK2G31L936dEbbHrNn1WFeqZLh/0wS16K48ieiCrRSUx
1lPZI2srvyo2iZdaPlhiELj3/IL32cQx7DDeLacnw5U1wPOyPQ6NkWv1mD6nhRFe
rGQHCuHJy61nzfK0EEB1SInyAnS3b0BQjZmMCBfDgu4ufyT89Xf5alDqpC8Oq4bx
W/slH3gUYToyNC3Mx7Q+9IsS9tf5ks2dgi46CeYvaqjXy0yAHGhdImf3IW64GPoz
m42hefHy1dacnQ0N5MSt72CvP5cU2n66AIyfuMX6VIaJjMUqz1fjaY5Y4+2jF1UY
SMmdigVZPR+t2rl6yxscmatyu9YbiWbPowyvnGRkjVUcuKVR/0rp+V4RFIIBWkTr
L7FaFpDF+gurGbJCDZbnqu1i53c3ISX8QpiUtnZt2tpFIA9Gpz2fLoc/QpqTm/4r
yy0I2NxU14TbXs+en/YcOkgZGtEwJ5MXI/WlxKj6sPiEQbsJMzMgRMObLCgwDwuj
P4ls8SJwQ2jJIDXOHlwk6IASXz+HNz49x4FOYXZgNFLubLB4JgeahoQeYp52W7Ta
a2HOE2ZQrS3ezOSQaS74EhhTkZPzArBR7PYcUDrd0FFIYVLppezZ66tpMnsLMh6f
AVsnzNtBbbCw8sANiv2RwZekdmt7y1e9Vk57EvTwVBFSojJI4gwQ/XI1ZCd4TL/k
gpJaNRg/qRMd2nv2asmSI2xkR45YZ6ow8cpNfU80oI7S+aU7b5te+R4IAHvye7nw
P3JJuNock6BogNEoe0kEhu8VnvqAVv1eF3gZUBjrhbKMMKpFpNhPVOV2E9UGbv/1
xCizcBRifZVbp5DF6gZ/U3NuDODZfchuC4VZu40rIr1hlP5p9PuWLR93Wanvic8f
IMf7LMgIr9GTS/fBc85TaFmYhusEe42yUNuAlhNYYUKX0w9GQMl5w+Sw96sX3OYe
CRNCkBub9iUCbLYTHkww0eLRwvMkFzhj5wRCDKphPGPbnFDbISc7k7Q0hNvCH6lD
qcI1KonHmo72K+u/XllaVUdAf5yofhqxYgcbeNmqxJNe44kOld4/z1sfuEY248cK
+EehmIH+rEhvxuNjuT+/bANrv/efWXH2dED6i5IRh4dWmR0mtnfr6KszaIsV1zlW
ozAZyLbwTOLFFI+RNmb8qynC6NfPWELuxWM9UKHZdmA6M17aTm1wUlLpEXcsdH1c
frDKMTRyRqmUWApi7cKhKb9StR3efNAK24ZJVxp+jG9+NztQmK0IvCplAeRmExRR
eWIM5iqI/IQpNfmlSMyhKO8M48VkNlGIyJUPkJWGzhIX96BzP6UK6/DCbW82lW/R
Zg88cY4v7qPHSo4fdnfkGoIIanqb1+bKyZTkGy2tGELwP5pvkWT4tyDjkRTPxbcJ
L/CERtsnN32Hy3f2lT8jX8aBdDCwguaUvvPLcUqgMUFkbzzUwxjdd6V8bUhtpRTS
r7vrWba62OgblAeu5+7jUxlrmGajICz5pH+B+ZMX9aOVjKZkySlBfJgoPt4D5DdY
GuCx8F/8XEVRJzAC0SqUmWPYsYV8uh8E9hitDVkGt3HSMigiKMnGX9rAQHgCrSEr
b/bJuSWifa6u8ZgB8uH17oiQ2tKE25blcQ3eH3pbrwKxfdynXkoxOoHF6KeGpaPe
OyuUpwhbkPoiBUrA/38MmUG9jcQwCCOUTjSY8mhN1zQ+2znrg+l/UB8AOD2r3WUj
XMSJm0ENi0H34yaFAdKKAqqibf5dqMr/l8GKrUInCqOGFVCUEBya4vsG/0A6rDZn
w9eJi7PkdGtzDfSK+w/BikQP2pojaxm53dvM9+BE/gmbGch1yGnOAfZbcn13bbZW
bIt38MG7qUiW+sMv7tXrtK41d2sg4uDMcuhy/x8S21a+YCOUKzfXYgHC5WDSwX3+
CiEcnjWAaxuOlkORQK6GQVgHhjdUPzue9uKh3JW26W18/KtGPFospBhsnwWl2pzT
H1UZyFtv0Ha37NnG15zlAr3Ie5flogLqq++Cg4W3E5BKunZpoQxDN1myMcNejoEY
uPGkfRfofneNeJufF9my2XkLINOLIK6p3Px4ST7ueB8qgAgDXbJTVxe/n+4LInaJ
EuOVWFHLc3Yh0w40gD5+3s3QGzbIhXrBzEz1oq1UAW53ajQMGrmfX7IvvCL/Gsjq
EO+3am/vHZKKWhXfMidz6vJNyUKqVW0AN8zwvfuSNOGLBenXIU3jFADle0FvdQwm
3IVEbgKGZNSDXYxlSTifELD7Fh/eeAsHTTSnkByrbQvfZ3TYR6QLy200cjOTCvS/
XgpWoE3dUNYXTx58Rt6E914dxdF0OhqQAeisk42O2B18Vb96qXt3qxfNG0fFv1PG
AWskAdG2fYaB7YME4k/EMbvh9hdHDJ+S80gK4/WzBvjnBQ+/pBt4BK0PuFGV1NFw
KXqLZMIsq4K6dkhbuhv9eXzpsOFP6P7Ecg6vMbP3vLJa+FTidt3H/gKj+4osMvy3
RCczyfsJuiGzrEPYSjaQTDkgrBQv8xQadsncfHfe5IVmepfGOt3TuGK0EYLSwgm1
zoSacuPEJK2P9RLhYJ3DA/4KwkpGTkwRYaWuc+QE+tr6xPxkmW6Pgc23XjxvkHKu
QayOirWi77Gpu+vXVYDFp/gBaNz0TmZNyx/fuHAnrzZ8XVC+DD3uSVM4520amPLJ
aHsmPrnNODgcgZWVE+NLcsYYd+8E69oq37ABKKx8ZtwapMrZXedXueEX9nLXeVfU
g9chMSVnB8WkFzfr23YyrF/gInpRRWBpRm9vheegX9FqQgpgFKQD93qZ79UF9Atk
DAcfAnyyRSlLk41ulYmIjMKv1yj5RaFC9XuS4oK+hssyEBT4qj+5+SC5/TUMPKq0
nCrXPFRUClL2FLTHmgGl5FI7SjWIaKLDQ1uIEgtLxLgTmysNguXBIUu7KNCTUgi4
HD5yOZC8EecpsuiijiwOuh0UQUs75uxOY+M3ldl66wZBHlt+uTq4G0ETOLa4C6dC
SSsWPDTwHu3X97XMIap2HG9QiN2omz2vylEXYDiAhwLTHXIf4ZHliMpWzkaW4x4E
5My90p24H5+ty7/eW4ultBe9T1kXaOpyjv60xN5L+52ltk/PsyHULYhWCu31Yta0
3N4y+iXhvA5+OU+e5ECm5aQluWHoSLuVcwgmtFTkFKC5S9zQAL/GAgZDi0iqgWar
XDmtP+ZMYTvdhd5LcrmMks5bdHZoT6PtA5rS25GTIzhhu+94XcFTu51B+hT1os6D
3mbaO/MAiDP9fZFgBdvdrL5ZlcuLiieAvjbAaImnZTPR1VekhD0/snGwpJu1+dTX
/NTPJveIJA58roE+Js4+3JyDMTsSw9M/89adINhA5a6lg10ujcXA5Ss9Pap/Y8kg
t07+YHwm3O8GCSXk4vZXyCRflQ8OiRTllp9rBCRgZHEYoDCJdSCzJfhVDRD9mhbT
yNBq3aHcv0HqOeEAkNFL5E6tIEptRz2MUYmdDjMn9hsZumOivIW/Soz2a75eLZga
HM3nG52/asbDjEdr5R/lGGkWaOvALixAS7syUfgWk7DyxpQYV7aJ8HZ0+HPXYC1c
ulnitmzRmN98/w8RYtyXj54uStvGs9Aor9xQ3D850cyhxTAKdBTqbm+yD7L51EUI
QByGN3HshY24cklAc9go6r36lq07gWX25SVqEQt9FF6Ty1PNhnq2hlYLDVz8Mdda
6/dsqh9A2TVh7vV7Hz5XvIAlGOgLTuRQVZDwjzFLc7BuYDvMDWa7dLEcjITbz3SP
z60SPpgA3W8lyY7VjOCVGlMx2sc7zPLdS3vznAYUSBD7RYvIEnGD2nj3pm4fG5Gc
bimeXfw9iW06aDICj4ZOGcGOJOfjC6YsFonAcmZhDXjQRYUsEWMQG4fqK0By1apg
0YekF4Mf6Jke4kCj5Kl1SdTLfBDngNVP87ek9xt3njkpIPwDPDG4LBy3dXponXLp
TVsVHJVztOiouOEhiT2efMbN519oetVVqFtiFvaK+vx1mJkaeW6Ql6bGXqRCowd2
6YBW77lL9ipm5XBiEp5/vPx+8PmH8yFo5fWn2Lbvyo8p5M46n/lbW6oNCEUPL+Ta
A58HKMdXKiWoNuT6xpAhQxTjQjAbHuuoFIjl+wCayQn+cCgWj5SNRgCqYGk3bBQS
p0kckl8kqZkpUiUWQ2W4PINzVKgYUx596jIxoiqBIhJbEZ1JN9fP1pVX1RaJw3Mt
sulok0aRC5t5hMRozNsDBAsgGj1hj8JBaLmzqFRhwNBfKTJb+DZcgSvaz/QSghJd
R402n0f68D4dfdVzyvUyXlQ7KYA/bRsWS68AqMH1AUdsffiLoxNkQLmQrWbhp43R
Hhq7cePfh6vQxSYhrKFk/4fk40eK2f2mFCsomvGdOgAvKEM4UdozNckawaAtPMG/
AW5UcDGsdX0KATvJM/DmBevXx6Dd8k4Gb01jViAxjF1Oll4jg0Z5RdHBvI4E1c9o
1vqhKgC2K7wA4V/kaXL7uYfAZ8DOYKFHlv9T11g3VxEQqLrt30kTnKTaGL24RRHM
sHuBXfc8Oe6QOr5hr3gGyJsC57ZKw1flM8a/e/nlZhWjKwgvkBa++rri58TNFoT+
ZHWZZMGFSeIuTOixLxvfFl/gucfHwuOoEmff80On9xm1QVYTHKFmic+Ic8CgFenL
tWrcNcL62J2vHEfExVNtjsaYsmJmRD1iW2UiaETjvWWHQUvzGXJJ+eLq9NyNT+sF
qQ009En+p5FZCSM+diUtK/Q+gydiL9j4h/CuGunlSdqNC6lxzjRLETQn2Z7JbqiZ
PqzKtHLoCMpgl4Hh1XsEvjVkmhV2aDNeiQXvY7a+BAQ8n9uAFgIqJvmdFY7sLtUQ
k01GrV0+T9zI7Z9bvBADbSuxiO+x5jwafxnXgqT4J1RaDZnyHqkfRXd60v8y45mO
c5bE7y30LQFB/cV+IAvo+hiI4FjKguPU1eDunMm+D45mAyeBb5F+h3Kz1Qa4VwM+
6D5BW7kDCOUS2tcMyCza8prDz3cAI6qytRCzoEj2XC/nL9w8+V2mX6rdOh+RBXlF
EuWSB3BN+TyNBa90mJNy12Hbeoap+aSOykDinsRH0UJgtXu5ALVwDrasoo0v9IvE
hA1dpp377QBmNfJyoax2Ak/tuiffPzFuzeZQZ3/1HkPuJQnaqBqw8GOPbNWkNjRc
7IUDku2oSAzsh0rU045jSEDsELwGLgV5bJLjjdSmnwldPZjj77ogsnMWpGm90uYb
aK7SA5pbbLfW6p1XR6oAoJ1B67RiFz7uqf84mOeur4V2tna43ngkhOjw8z3z87zV
i7Rm0sPLV/1HvwVKz5tAaMKGgbGhjdwH9QKL6MAREkepi/F586jzmeok244qPc1V
9gfwzVL6tSTP7zUiepoH3ooCVTV8cEKvV3iE6Wnc0V6vQ+REQwRtqyrhoOPrIh82
MeYcWWZsFvsmDtwf4hODFOB4+yukCLJvEsPlhDNKm7+5Ysr3lpPHJo4lhsjuckkA
23k7UJlprja4qkUpFTT9vB9TzGguPpB3JbJ4BzRUxGE39UcinurSIdLeHow+oL3p
SDMbCoBc6TpvUYsChUmrcXNSikmVNqvoCn1Rhbp0lCzAGGNO6mkPnFBfbL/7znLj
S1jLn0w6vFzYvxIGyGBigx/SX3cvQ3HBiIf3hdxXbqX9tk/jw9o9qW+lbgpYOAkM
j4ggl8iWWpxvriSubshRpkGwS18xpzPlzsIv8/Tn+wD6AcsNmTJLp6/jj4unwDzT
zUy7b8F5iyt+BxGdNpHwsajdoUJ3f/rioMMFKzzEB2cuYBZ6GIA2YSOHL0SOga2k
5GbBNPqPVBhMpoSMlswjtdZ1HhvSwyceHZe90/6L1GOXxEqUOxbNkuxez30g/tS0
/buXBAJrtNiwPVggESQ5FrabaSJ7Ut0G4jbed0LE/V6G3mrEA7le0fY7Xf4yR2yI
Uav87sh3oUfwIQtDDig6wioXVb7W4+r1rr7mOpDBwZsUtrZPmSPWUVO55uKDob0a
uY5h5sGt9MmKuq8NQ8qyeI9ztHLabdPrZG+Hkzp3pJF2ra+HUcC8XtDusyyBtcKt
kF+fdtFcLMCn8boA6rJlACN1MgYomQ0oT0a9NhFN8NZiDWB3Q1ZxWM7n0C/2JzdW
fLbNyPO62bq5ZmG8M2KMjG/okPW4NDqUZvKR0YISYJjmd5iFcBladlepuUFRnWhc
qrjTLIUbmHwYXGbVViGU+pknoPpgGrStwL4+2sGlbvIMpKMan5kWxtbs5Lj/EJou
WUxYn9Xq1uj7Gb9ItKS9IG1/UvayTSFYpXOdSk1aFoxNmB7ogpdmuyDPcHLpkuq0
gwUZCx3GuidsVcHnRV6KzrDu1ANgvwCRk2WeC9XHV3zdwxHB98IfqoCjm6o0JUkS
wHSW5/FSVHbMvlMWV4BTSS2FxgBEVEqMmklxEQuhJxplt8XDXAzjFhViYVi4Razo
goSf4wXXRXGwrlJwvkhA+qiOGDqTE3FZDEHtIn0jjDNflch7eFS6QxTSNz92DneM
0LS81KQN1XMl8/CZ+x9eXnoSp5PKLKjrmY6+mRfNczILKcSn3pFR/w0AJfRMMAK0
N0F0dls0/erp73KCgS7sgbcXaGu4pUcY4oF8XK3GiJqVLi/09sSJ5UXWY7a502Lr
K/z4BMjBDNtKsq+WYlOrioSKxfTJ38semNlPfcxSMRTYGk8dpQNb8bJ8Lwjj4wmQ
EkX4y1FjettAm23uF8DYMi3tLxvGJtG7YwXjxsd/1Bm99kj2HKJs/3fEs4HkNzmy
4Re1iJypiMErFGfB1qCjQQKyug3+K6j5HlCNPh2uxSMA1WppZLZoi4sfiz8De2xF
ichygkOeEVdipWUlVheKueCkhB9+fhL8D02h1PlKRysnjexRLp6X0jWYknz3ExGg
UhUP4f+zIWtlDMu1CIpJ8sJSvgMhouHVeTM9ifS54j3929ZZS6VpH9dBiDIxlc6C
2o7jB4B+Y5isi/8/jEYYAZNqMQRinXFMP7jkUsxHB5dN/+9CErG9yPGZloSmpfjp
Mt2XAZ64pb60U9IfwRJFTP1DL9Vq0HMhwQ78T2VzfFPGNxJbDXzkSU7ZG1dtd8Zr
0sbm22K2IxlSjewiO8yQzevQSlMr77GnTJQF/K2ScpDiBwwGIaN/Qbml1fpg4O/b
lAla9m7ilA6ZfjbJ0FX4ROI8/Y54GI1HOzpFYBN+cLyNxoQE50Ke3oCuNryIHeVv
uIG8GFPFCtjCZSDHvj10UBqXtNZe/zVmzHmOuBdZcI3iZBdkDU5jlDwxyXfZ1bdN
ZGEYs8RVHcQv+CRLzLuHnumiEO6b4O4am/413wDjjzQXB8QWZLxLOg8VRzoNIQvh
M2aPx7iKCzyWSD8/vsMzAv4oGxt9hqOZOuoebIlKSKKpkXqyPkxHZ3povtdTyEvQ
h9mRXLoPrW8ln4OWSvZE+xx1aimeaZ2NbqH0Rt9J5ZavLVsiOZJPrqBQey16paSw
6UGigJiIqg8uGe+Eqbv5Z9FaY0oDvav9A8dWAP4QtHRhwetEkcOFADLKSL2sBGtS
IL8lukm72rMLz2MgMSgPszNMS5DXa5GY1HrCtNUxxzvWLC4S8nQSbtYjU2trRGmq
FoCjeOgOD/CrnuVp8iNjXe9GdqT8t9rSXbie5yjnbGyylxuDTcUuctn/S/Ab8Gyu
Q5paxsAhvhZKDfBO1vJk8ENCqu1dI7l5DxNH2BGbROrqM5G1Ma9IOa+zJAWNuuDK
T1L+2XKqhM5LX3ubYPdpMQwOhMVGQ+9/TnIRWFM+vuCWvunIJMDtGtXHDoiEBOq6
S9CThdSvnpwH02t7eFSYf+FId7X9bmMFZKp/A8fo7399Db/jeKBsxPLTclGnKRiY
yijqQpA3CLWUTYtpUrQJM3C/INrmYi9euoFK5grGlIhk9gARd7go1ue69/bwiPdz
+xpO6xwG2n1Sh9/RIjH6AjeDCixzucWzN3L8WfoPg9Yaq86S0XLYDQavpZofXGnK
pwmomrloAj12kYSUhxhBnarkCvEvBVBhjFo+lzgazZ9mgedNv9myUH6r2DV1MJU+
nw8rM4EPsfPUX64kn+quidYxTZOXqp6PslFBrxuQLKSC8v8C9YZ0+Co+opcygUfI
3wIZtY2fm5A0JZ2hILCQl4jjNohu13lLBnlxWvppdm9I0cAWmx6rL2GlxPEjw7cI
OywCgiU6G8lEBjYSnTKxPg1EnT4gsVmkmQ4s6HW6YW/GNU/PHOzaaL9ZTlduRpVw
273ZXpN2hTW/Yh71QbR2nGxFhviaVTpwcxdk7PpM5YhS6xJ4WGSC+oKs4O39Jzvk
CsRfUE2j0SbFVQqYi6qxjklqquetQ7uWHyotr2riCqoLJ+IW5d6vWfepMiBEF/ro
6m29j3m73xPz8FPddarxq59Jv96kDpSIbvKy9l6/rNh5imqudrkmeMGXVE8q7CKG
AYe4kukobVZPa711D/laeFu9SxrBx7HFzO+DOHNBqGA9FjDgTYDCtKD1BJ8NguLG
8/SX7k1I8XVg1quDPDeX0yidvndDzfG3JhC0cBpbz0yVGfdPwIkVUWk523e6TnMH
GpveyKDI/3R5OxiX28H+4oemU0ff0JCng2xQHpx5+UPI0Ttry6zdeS/CU60ZCJcM
HTd6SM8r8OlHbNW4B3m3wdIMMBx/6Wo221vHNJ/3kT3YF9hmiffcKtDvIC7a0jRs
4XzQHQwXPqZ0q9/Fbd5fzImIjuQbr031mUEJDUrYhTKODnIDTiy1o/iVlZ9wvMj9
YYZcw/tiuvHi71eY1jPP96/HbDsY9hxtClP/HGy6AEUkI2P+exBxW5iPJ0HqYxVN
eScw6DmwylIOWaB5SH2V6nG0xpZJ3skTUrAT6edi8/KPkDvNkjo//d3oYqWdFZyM
pzWzf7OqMSkNC5OcTnrxDUurGPs2pOrkfCIY+/wwm7kkorx1ZOgyLkN2Cf+/LuVF
+FJ3/MuAOj+R93IS7KC+sPEv9C7Hl9CPW+thtbos1YHcgl6FTKcRSJLGDfwZ46L5
g2qYJ9t6JAQVteWArTaNwOZuCuJZjqHAllinVQaZ9UlbNT4FFwUOLDYFYBWiqnjz
rWwzscFUAU4WsC6BWtYdRnb4nMxFgItsc/0qcFD8yrBuZDwyLNO+/5D+EsuQvyhd
vLFb7mvH5pi98kGftR2wA9GCYxneonpe2TbgjQbwjuF90p7LNPMg0zdg8m/GKT+3
rz6w5K9Dvy/UT5zEpmJnsxlUiJv2KKgdmNcqw/NcJoEEIEk4RREQvZqeztrXnO/7
50E89I/uvfhsvjjixM0wq76rQxhPi4a9zJAKZC9G8j9yfkcGzMCfWC0hoGG4t25E
SpBimjm8IFUXFkLGsufOU/NnR+IdYc6EtoVtlly+dKIxx9HXd1JcE+9CYje55kAc
SVXSnulIDl7iD//FQ/ISKcNUdH0eeQB/jYjfaQpYmZBXu8BH65lFnZPmR209ojNJ
9GOzcI+pQswJJZmxdZgXLCHPYV26udrv34HqfK6rXxpt8ZbRyn1Z6G2w3I4in2mV
tJy6MvnKveHD+h8f2RwKBKrQ3q63KYx5/svWB5m6TT76Wh6oe2FX7hjh2ogzc+am
obG3te4DrdcZ0G0opy4sUFjbSbw8MEpI/L7U+/AD3E4P8YzFjL+VhldTNykmujWg
YfWrMY2WOKoYHPxi63bR0vMOJXKcecFrLfzNe68HglUwl6SAMEIHIyNe9XyN61Sq
/aRtFOTR6OnAP9LwRdJZ9+HE4Q+ZkP7HbUtAPGtTWa65ct/vTd9HAGZBZk1TkZQS
ZzisfilV/kNKa1+STlLXCx5wpW8Y6OofNkCGEFktCn7ggvDU6ubkLRHqoIKNY5Eh
7ZsvARai20t7vmwFlvxHVnKQVN2YrPc2iZzcQkmmxKFBEbLi2BV6GB40/qvsecKD
HiObuYUltg63dP0JlVmGX3oz7dITuV5CJoKSLPOSVkqzI+JgAvEF1+Yv9oSxbtug
pikV+AhihQJ+/ObtUWxNByAKGjMR8gjRKItVS5g5gJT0Mv84yul7P9A7CHnjyuNx
dzDjICqJi/vILclOBWriZ1m30P7+j1Ep0NlrFpGD6a9xLHW7nCwGXSIYudz27uVU
EksFoXypQFuRcaKB/XFycBv7Jd3bxbntAst1KoWTHlCXW4fiHD1VE7T/vrQTGRtF
K2Ts4T7SajO24CYxUMNLzp/ViGERwx9vkeTSjOAXvnXUplPD7bzeOFEmStsigbQC
cxHl4UWOmjrFnYX1Hwfx4Q0VUlHIt66ZhuxAtQfOcpIFrmN/a9HAjdxVmf71DVdH
HwJmMoUlzF/LQd6kN+dI0HxMr60SMGbt2Qb7pCFfEBBOjhFhBnYB7vRTMQtVZKyX
LGyLvWMrLXsh4KhI6ShwqNej2zCE9f9AMk+02O4D74o0JFu75jzPH2UIoQNtsdoS
q8kbYNOrpxkojqINlHTzIZ99RxFwy9hm6MPQHDxveaz28mdYq1fqCoBC83aeUkdi
eR8nee8sdcMwhz1KXJOWPA5RG2dihY11wEUJP2QBPx96+f/QD2pzq8+DfloM+h7m
qTFW7ri3EcvZhDuBitNIeG3a4yWukg12C549+f2nhd2E4UmSr2SwvylOacyFqghg
xfG3OANGtyxEmYGklDLkeEFmFo9KuTKQEE2O9HgP8GJzCpr4pKoHpc3eOMFI9B4T
t/TyCQ3xNT7rnhNDAa+Yy6DvRQhWlEy0GXjXVrWKFbjE8bM0aVLBAnNDxTgqOhHA
SJEmwuwHC4DjQrKDhbTdgw654c4V/H1I0krtB80X8BGZp2ge3bRa+zH5/OKyB/lX
lAvtyTnPQ7xspQG1FTA6hrUxK/cngSZGdQ8OTXSjwqkrxc1WJVDpQ4OQIoqcUl4Y
MBZp3tsaUP6MCCF8nw/xX2208DWXpaxQES2wqDS5OIAnsIpdUpsovqSte1N2dZCr
1GtMWWAdCsWqVJrMGMnTuB0uCRh+iU0F4AWKh3B8+4Jp0u5YIObI+72XbNQsR1+h
2tNXYv5AqKvogMA/dmXHTz0b0BOfi12eM6de71TVirjosqv87+ONrdTbtmwP+AXX
BEMOyFaALipBxDIh/mqQUHUMR2Xfav2OQE4CC5MBkW72lQ8NUQk5mzy8vs6uEpXL
j9xqPgfVqq3ekADBeZkWSAG/fZMVH4vBURw6g6fc7ecYddUZkuSiZq2PmIUpMx6b
j9cO6mj5QozH1g7UBvrq92rpKekBvWEhazErfeBEsrA0m1t23Kh62fZpzMe2YUNk
cXwfXgfTayCaer3Z4duSw153v21IJLY+mCxl2s7a3IjamsvOaIhshmN84rb/6riL
L5cFcsl4sSQH/sPlBqOfagOtFIUFT+MYuz6geLPeumG0IHgwpxi4yLSheII8R/sa
hHAq/gVi+1c4sou+1/dHVroUADUO7PTNNTVVJdoyCNdt/TBfLwj91wSCkUzHK3H+
DBH/TU18UVqeUhuYq0m6VaKmn6icUwbQuV7eUO1HFJ9+FHJA42v9OMZ5jDB6uj1r
+mhzGnZO1laK46rGcAb1WOAIaUy/F8D/3D2WBfQ/BAQaN0Zjv5/pOcv6ZTS1F27u
MC4awmthaZYVk5eJlTSjfpPrG3ZCttS6/LJKI1Xj0eR05RkZh8yJkjDXJeB2Kh9S
Z9vgIy9bi9badjqh50N4mz5cArMJNarJGYNR370ysoDiGc6N3oa80tWfIuYAMp6i
/CYK13nkCtfTKk0rYg4Ng6Cj/0FmOdtPtyCJG8tWv8WsBVENNEiO1tXBCzWozZhv
08Jd9GC3h7rk9RiD70UrEbrx2b5zwxEakmyp7bnS5cVkL3NbXlS/L9/GDIhk5x5R
U23APMgaFx58RCN+AeLB0uFji7BRuOxzcXVn/jeaAoxJF22WK0I3sScqF2dtxBmJ
mz5+JoBTjctP/5CAVqegGKDFKuxb88POu33eRV8pOFXjoV2MyoTj+ulDhj5qF45q
nixrMSja2xk4shkRw5lNzoXaUAJHdfEifIYVgzVyrttEsJXfSZURD/A6ljnUQ4Gl
3EijesH9eNsgA3N9mrxvHRG5yllE/Dq1I4lejhR05dKuqMxfqtEE2ZrnZHJzMnuf
XuSsVqP1bZeFkwFqSjwdOEPvjkAGBBbta49atY4/SD7p0cJWOaq6kMChwW/0jaAy
BGoL5+9xuhpI3frM60+Xhi7ovP3Ghd2207di0lxBC494y+OXDDg761BJXh/hAbsr
4U9noJ1559v2POxvDk2/suNy9WuO2HWQOG0rPFlpYrw/mRYN+86buFerogZAlsEM
3TVXcyfoN2T8HO6HhO6Lx8D3JZUJp4ve6b05ResXRvdFLG/UvVQw97hlvkpnX6W1
3TU1U5zniXg7n02nouqLgI3VK4lnIQiPlY6d0Jx6lrgnbUT8miJGf01mFICcYt18
iTWxhf+JMZ6BInnGtrdXmryf6HYyVYBUyyJkIilr3zniFW93hbbRpS0m3gz0m+Yi
d9CkNnyV2ham6rKFfOt0h+uESS9jHJ0W1EdmMHiIKgQAqTlR9P5ttnJYo6nEjOFZ
NHjlEwoi5Xx3ENv+x4a/DJLr7Ju3taNqUIBjYSvGW0/edtDSQL2gzRXVePD7B/Zz
G75W0jOH0RrmIOhSgYi6B8bmhv/maJzedDEhnKCasYmsR2QLadnjLrV/f5korWO5
WQE/noeLB9dKNDzkfRQoUM7wQzQYO49SxPIPW93iaYymmu7V9gW/g7ZB+slsQdmz
XnuovGCISYmrqf+ljMoZPBvAdi9nzML4CNfW4TpcOY92MS4k+x6DzBnPM0PpXVoI
PRPBIx/axyKIiqS0mrlQ8cg2+nscM5pFy1a+8+1na3BTjVAWLovzpiS5qUwngTK7
Dmt042L+vpDCurk+BZUV9IstnJdGiaf1Mmq4zlKHsVI+hgG085L/b8VVLuyzHknP
H1YNYOZvaj4o19o1zRAuL6Uo/mMBVHKibGkcx8XMxcbC5MRoa9fsMu8XDjnizFiZ
rIjORkrXoEevJJE1S3Mxy8vvs4Ej16wSxshs7CPxSDi7QfB3b3OJQ2D9CD1gshoe
pp6vplo9rYlo7+woV86oQQ1QCvJwL5TwTxnrAnEj+V4TVYwGl3/stpceqA6JjEun
FUACtdunkc4h7us0cUGcunaZ46CIBRazAIXKEKlUkBYmgohnvsw6SpJiOO/jMGvH
0A8spikpmeB9uF6wBxaY5a+u+gR3z6PTaVsy1PxoNbJSQ5XriD43T/WZn9Trt/dy
y1/nN0R+p6nq5GhC4AUkXb1L1KAVhcf7GCCBBeHebuaSAQdC/OS+4bADrIU6mmPW
1rI/YcTP3ty9FRWd9Ck6WBVwOs1KI75artOonv2SXT0LdbIzzXPxSEC30GNR+7pM
d58e3BCd+y4GS4iS3+xWg2z7tXGYfqLgSyXODiCve+rOC5svrA55gPbA3m9I21TN
HbZShY3gcC4pbnL2fuBqp2cmS3L1iWR//wdQ5Cv0uWqovGLpY8aRhTxTq2HqwB6M
ulFeBnM0cKYkkjoRMXvu5gwwjXTfoIHklLuCwoEjRGgkUf50qR/85iiLJwPoUNBB
nvgrrIkfOxXkKDEck3yA/WFeX/Of3WKm2QpIVr0AqeGnONiBNVU4gSYiKuVMP2PH
SQaKa3b+au+bVhIVeg3x+x37Jee5Dk7gyFoW3uwSPKlWjGaorZPEkq/j5jhS+j2D
/lXANdLzEnfAS0prRUBZxXir1sMSMvSOxBmFrs3pN5+ofMd/TNo2wjC/7E8dru1d
zJX/ZvhTPelwUil+MHRcM3V6oBjMYq1VeuJTKdcGwAdlZu5RdOhbP6vKYB7jd3k+
qV/OgVx9/+N70cQMen7714QHCat7OGC7eevntlntuloewSgV0N1PNLigv41a3w0s
vXUYwHkgs5BefVk7npSaI3WUc75Zd3QuIdb+Bx6jxSw+U/014zrCf8ENQ+nfxV3r
eQZNZHPKbwXOspNrDw9jOYjDLHFceJr+a04yvSy8PcoZ4ZsvDyng1rL3eyAvBqzJ
l/N5O8gpjGJJ4IXl4Fb9zz8tETU+sOigyfmCLjxxjvVPFCULyqY5izdqdaAgrrPs
PTgXhdhac4aa9YkIvZj31+eX97rGfAywrQtl+goGkCqCq3rh2k90ha/bihznhLGg
DPPu34thaY7uwxTsBEKUF48D6QZG2zauA8vCOQBz8op/Kvd1HmZQKbU1uwFTVAAh
etJXSaAiF5LMz9lgfT+9TyHsBfEWuH9zp2stxzx7rvSiXHEpOOfgQncq6Kr/y3Ww
RPG6ja1Fk5VyqpchjZdXcp9axyPyrYNCI6mHijcmFYFyZMALJBwWdWjghKavEjgm
tNQ7CsdK1+aXR1/U+aJwUaL1bPlQcJLKvpGK6FtyZlnPlXOMAwdTjmZIp2L7NmIg
3ZnloYYXSTWXGO1V2nMLXjqyPwVNtLm6nnL+6TiykrmtX+8jabOPG6ZzX3lfd6Ea
K3ytIBwUS0cHj9IRmK1yLIvBf29C/TFEOXZHe7H7s19Wlh8pLrkRlVZw+OUTnVFq
lYDoyn9UXU5BLrcBpuxF9slzViu+fU+Nhh4MwQal0V2ee3nNyJ1v6Zln2sii5anz
YugriLoFXQs8ZcxqZbO8kXt+Uz/OMs6UxoafB8ljEiMpijDoiVD5PKfOuku21Y12
2c7hStVKvS1bFjoH0+jAztITgJk9+Oji8iRVl32Sp4U2J/gpvxgtqoQJyfgEiPxg
Ii1lU25bhNvUCOvCZe97b2puwP6Kl8qf/H2MPZ7jW7y0xFqmsk1YLlGUUPYBWceR
rdOm9B72agEzH1BDXuzebjwuuF3cSgDTAyj3yHZxqwL9ENvGvgni8EotmwPr7jZ6
y6UW6IIRCEmDLGsO/qT4BEy4UYvEdrlLjChfuATeVBFgZHIz+WffORPTOt3ClCRM
7CSCetTggQssAvJ9wY9C5xNSt1UZasMNMTD81SUpd9a641R3zODrcfRyQfDdK9+s
na2GE8p2bpOvsu5i+Yrbd7q1CfG0aZGyM8hwFp+SWo0/68rnDO+3Ms5vqD4SJRo+
coe5CwGHMqn3Up1cGKh0cmCBsj6zm/IPkL5KaxqYOdrIkVCtpGKBnAWjFs2ASSzJ
La6Bqo5dKKwIGjYc167TPqYfZgt2MxkyeONxnFvG53WcJuPVU/ajWxkCjU6gAAf6
sPMbNBrQT2gt5101DIUdOsuc6OmVIYLsTC7EJLMF1COCT8PFOp8hbIiQgHRmdxY7
Wkby0JlUVCvcwqygao4gNZoT8aNd3OYknd7BUvTSQN9A3+R0IcTHC7ctkNIauRHZ
c0sQpd1Kht5kW483Yqme81RHiRecJ/Ynu0IxhjoIyZYSyFjVm9ha0Fg8z8G+l0vN
+5lUbzZkZydtWUIczeuYhSNiCnKQTlSu1VVuZmRq4/Ctxp1unV8rs+uw+x90VvnX
00TYEGt6jP3sWjT4oukxFwyxQlcx34LZc4DfnKtm1Yi3qC/MLOuXC6ABuBeFNBdi
cKPL58hEmCYT5G3/yozHXPIIhlsrwAUJW+k5+cIpYrT8/Os+VRnblX6MeppIJYfT
kKZ2M5cuwqjOxAHZsaF+ZiEZ6bQ7Z+zmnsfToq5ALhd6h8syK0Fwqur8leYUqysP
LgvSt1SYGpeKbQB5PPOuC6pVZTFLaUKVkNgfMeCB14KvnvuHSzJ2Hu5aV9rrElVg
tsVpeM3KDYlDznEJYBUYEVwtC/sBFU8ko4D/f3AgM0aQPUZdDOVPNP4AwQBvAb/x
wofETdwvCy20Zlh/eXIvzSoGJtAfw25QeL3eRuJlkrsk9O2dhivZJlhCPQCbgzmG
CRFUA3ki6JJAdNV84upTnEYtOQWsWdBul7blSqiEnPmx+A8odKlUvybLVyoP7Fbc
XFxhF31JhewKg+Svr/OfjnHg+aAhGF3BnO9p3gQsUI7dLXv5R98PmMaafD1pMTPP
Ui5dNIYLiLX+RGH/yAMqK0zkIJskQF0wlWtn8vsK3w0lN9emjFLA9Qtk05BknudN
oFOdwZ8uvJFFJqn0tQw0/QoaLBRkJ04JyWCfNk+XvNPniIiqt6m8r8sleg46c+AR
mSebSIqErSzkl3IoHiT27AESnsouYemHz+u+TvUYdAc3UfM5AvXnUuOO9VPsz31J
YW9NXNcETkBYom2Zh7YYbh0Fv884Y4XxNOwQeB7BFJYYLe/evtmIotuWmDmfBB/v
zkjdxtRuUClzyScgPAqhCFZDWt4GytGQeoshcGhcuK88rGKzSP3GyrLsJGTyWX8F
UvKnyZSBcAZMjkz2Hvo1V4xZN2/h20mlMsh4ZR48QKszgKW6rco5vfvey6HRMEqq
9Wg9ENi4cB8iXQ5x6WK8hDAY9av6Nqwnr1qOlMIQOH2SjMkKDixnViADGP8l7GwC
Vhba8gwaTNaTVGnhKEPjvlD4xQx9O15l76fCVeogpjNMunhmhm2WsAeLhBfx0Gl+
sjHQFNhv9/O5Ka38k454I0x/vKnWv0HrT15kjT2kILZkPil4se9uN5tjfZqIx6QM
YX4gdYt117X0uu+AAO2TatBdoedG0x9h8jeSv75knKd4nXgtbYrMTStlJA2q88lk
8c0H8s3C5iTQDFUNnAyW1Jc81F4ku6SGHiEG3R+6eM8q4AyDj7IdtJoL4yL2Gzu/
ian67u3aJa84YM8OoDy91FK/qNgmWtagQkzTEeggpMKzlRIUzIUxwlAQX8GLAEY1
5Q7jE6vZJOmDxqM1ZNWNYWSt/Zrm2cTbfujpwxd1syDqrsm+l88PfRybtY2Ux9lh
6rQE/eYH5xciSgT7LTC+dKDSdLBZzF27p/2TMx+WJPs3iDAPF27418craAv60SaO
gyxJAU+iOFKFAQTjqe/2MRNLrGyPHywQTGC8BUhRgWCiEkNaLCeNga7KOFJ498Y4
nUFKwxum3v45Nl9cl/d+zHd7DhTUNwj0NxsfjFClOpaMJW//aEBhHyCijBDYi4TU
UJAsu13Z8q4oLNNJGnJk/tijTb0P4t3QZIS2qxV1rHk4uUdOUXVHkve4cgHB6nc6
ZRRuSLag/bh72rKHfKm8CTt/5KUUjnNH7rhDj7jO62j5i11jUnoRW/qzUNKM+w39
yn5Lgp9l8RBWJ8Ie6I5eD/+l+LDRsCmsgRbu26kWEYrXVg0iKQkU2LYWnqta5IF8
R6FxeopfSRuiqyG0SsQB8zxjNcnLuqbfT52A9hX/8RBFBxXfqswtTDi9cwk8rCCM
C7MLTERP6GZZK0iUdXWgNv4pFl2H5yqNg43QDcriYDRW8p7drQem3PdSUm8QcXbI
Y4j7a+3X6JpFUXSWvFUDUA2p53L7lKL6DowZs5nsuOggvx6Pf8r9bIJsrxaqbj6P
jQclgfmx+wE4hU4MN2vkv9OMjuEC4GGE+uCV26/s9L4h8LwnFeKA5AZ8D7fJOlHR
SqxAdNTEI5+UFiASa8BN8P5Dck6kdigvMHG7sd2dMs1OfS/O6wnGFZVc56JJzXmD
g+Ew03EhcXpEvqsuCEHlpo7tHqFKlzMehJj/veEIvnidSvrE4adOXvxO4gV6skMo
1YQCx4APG2VCp4vPzyeOZvePQXoTLnajz7OfosFzPcNQfMNEiBp9PLK4PJlXQLe2
iHQumxrpvS2dUytYz55jrbp/ygKXcWTpcs09q9mM2FVLvL7P0ny1HwdrBEYj3yl1
zpsPMg7//O8gVcabeVvjZPaCu3QWeXkjQj9zVsC867u2VY4mXD4+fkGAzw7fYOJb
k1S0JcNObgZt22SCSChd7R5JBXVoW1JuWshCw5ad+sgHCOvl4AKFczKhVneZznqt
CIY6ZVzz2FCZwd0+UjTt9oDlo403xzKM5h4JcfhHoTil6asHTetG9tkFEAUTZXTd
3qaUz4pOLPw6Qt8vXVfbAwaZblfobR02t42jjai6P+fwC6C1x1AvAxiQA10S+yjx
/rXQBoKtIimteDvW9OtPqWiRkEJpEUl8TcYXqITGVXUlBfTj7ofez1c0kf0ytWqa
NWsP3l928E21D2BYZ0bK+pNrHpdKYZJw9rV6J+So5Bd0ZIPZkAk1t9vamiJ9suBx
i9W7n7HbBd+VTZboMy7iGZa7rcFTOJLSM3GYO6PbZBhdKaZekajrqiWGlDe28f9o
dnClFEdDbHMVcHqbdhPdc8sxpKSv7CHXFhcxi880hX9d4nL/W5sC8376KEIi5PQP
/lq3t7cQZbZtlJzv6B5FjJUIHsggNRayzwFCoG6uZrL9tu81DxNirvGW/0K06sQC
7F1lmq0cn+BXCoTYBKkdJO4O6CluaOlFMHsopl+K+CDvtSqr6JNqPkNHyhbfhWNP
TXrM9KC6YPu3Z6HZG1HI3YW47ECEGz725wlKhe1PN2tZuUQQp/Om2x+g28Gyv58M
L0Fg36q4Qrtjkv5eLHd3ucj7EgmXK92Oraba7xQCMwolDGxX9/qdDXeFwJvEU7b1
Q3OJepjVAVuXwwGbyp+pa9NS9wvaTO+8v2XznsCjQ/YIeV3JsOGVN85o99avaDZz
CxJtakHgjmgm73CNDSdq/2NKbBzahXb0BS3JGXRLO32p1jM1RaKhQAlXpVOMaWmn
VjSJ3z4XJyBB4F1h/zdQy5o44J415XbJl8ZV0Q5V7qHzZlFMD3x+5jRCSS3MVlN6
s1beYAD6ujdGaUtL/U3M8lmcXqDx8WQCWmI59ctuC/gNLuKliCxklggHVZqPScnc
o4Xr149Ott5tdrMhglwi2jU+Zg1oHstW8273b3jxbsqpfsbfUzivRzKuSUGekHCD
VHg3T+fCNRYEmwdqMphflWYIM0ih8gTX6w34BlvYfhhcerpWMvewFBBhUVcyEJNQ
tG0g7RcOaBNDtke8xuIWv5QJKuPtG4U5zKlrRTQejgNe/9x1z8qy2F/5fgoADNNy
Q2fdmiWDSfK7DEpXp5IsTAHqo/hoLHXvdmvlVPeXzWtjTmcTvXaB752pUz40zScb
iedvDP3ly0vwZY7vZDMOXccjTrU9OHE/LBl143edptmQei/Y/65NzSJGJ/1MSjKv
DhauQyiDR+A7ihDStt115dhIb+fChQb9KAEmpnfKdZQupqPUhgReg53tph0+0MtH
7vwarf3nxFCniGIqxVNaW9XRsNphbK3tt+R/G6ekYw6MbkyZYI2dFGAM+MKqOSIR
YJ7B3rG+AbLzaDfFbTJSEUWx0w7HbqhpngUEBo6deuzIly0ijtkuEh2R7FBYwNP5
n++tLqvCqTa/P/s4D1qeGN+/9Z0EHBDad/ZhXRczCkP8ipk+RjobtSJc9fQAJeKl
Mpru1NCf+HVb4hx1XCLJ/cd1YGAvISSypS5s8jtPp2gGhCuEBLcpu/gbvtGadPR3
CdEf23sasLMh3IoYMQ50PjZdnUf7VeIn+N/0bNktFRd57Jak2vNtvCNw3Nq12tSP
t7/UwihK6EEMu2mhco5wGAA7QHZ9XIvd1Ae9W+4szmfLIosVj7R/bR+FOTOASgJO
qli6M/V5DoptBaLkoq87gRCqS1wokI4T5b0KFz2pRXC9gzTRQ3MjIAwdicnEx/T6
/+qsD5VBBV+qma+Msre5nRaN+dzPLAPBR6mjQErHr/qlNDV9JEaPxQnRSrJOrkn4
ijjVCnnyWfYsvFyxXYtRYQJj3yRGqJFgICb4UIShL6P7z55clhGIljd3pZkO9DOr
+ftrJqLV6G1GaKou0qmhhP2P8m7tokVWkr3h3eOoT+X72s4o+tZY5TdrofSU9aPD
VagRD18R2ggAhiQS9suHkvmZm5ILKgjudgeIQUAN+Oba1w1rLrxuL0Z1FVIuAuxz
4zxrPTo4eG+LKs8QJQpkTxaoTAH8H9E1J66Oq4Jj+/hbdA6JkS/roYbt4D0KHEn+
ddywvqMC7QlM3KU3Asa/KyUFwahfI9o02k6HrilNcRGlQZS6NscSk7MvI3VZZYuA
e/0t1BxacYzysV2K9RjfZHX9wKUx+mFoGDL9Dj0MQbwQMB2p59HwTHjzzHzmeAdV
HFsIqhh30IEoFowdfJlfvaHUWutDmi7OWMAqR8NwbtL1vLCDGYkj6WwnH7OnR3x8
YK8JAkDRwDlNos40DsutgDKBwTHnWmxQayPMnkfpWAYI/3b/7jb4irjcFE0g21sA
USFjzToWCD3dlzQX+hXPtWUezyo0fBWbv+xJjVLYMzkZYpbDFs9chdk9a1LLIHhi
kjq3NanCcOvXQWw8WFwnj5A+vp4cKEVbazqw89ht+JxavqhfFx1xFFsoloWkenKg
SGIfIWp77WpDJX1rez0GdO8h52M4kQDsapO5Wv3ZBaaFsTSYH7YFb5oxe4BqPrgo
ZZYpHUvIT1D5k9Q5W7KweZccnxo0F4pc8aweEGgsmlDAE+hxk+UcWnJCHziIs+Z0
hrqjB8QeA2Czz4V/Uzj5ZpM488pwMr6vll8KfLOsH50sNTgRdSeFKYPW+db7RSyR
KhCkaH0eBwqqCUS+Yi4gklBr8v8JrWEs/kw51cdVdQ4lJv0q8eNvyYR79q8kCfCi
YlJ1gWFYCHDVrU1c6Ty3poxLMjWw1vNdKA297d9qWpf3Wb9a3A90iZBC1CA4V1NV
Uee4MAD07qIaQ0bUm+jb0SMn1hj9RVS2Y8COjjimKZuban1HMyhr0ETl2j99H93i
5AxyKI5atVyQGnECY7jgrsiU4RVMRYHeif3TXeC1YhWIGfyYCbhFkUzeXXdp9/FT
e1l2AUMX2FWNzBpMw3AHrHAZH6Mwj7dWVr6JKV18racXWqjsyerwgSFDNaOxIM6B
ph3X6gAqxP5aRaCg0jNATBxhNBFKZWabVN3cGPjzczeegZoxUz82PrszT//nypWq
DJwDdg/RwS11wbV9gB8EzGEHzl/p1rWDqfgYbO9BTVMo0XI6SqqZJoXsftradH2k
UJ58Ae4iA56a++50IWu0nGjLcI5rVX5NSXgukJHiXG/RLyENQzJZ9/OGe3gwvIEE
zrJ7P3zLHJNYAmQoG0dUnj6SjlPx0OmMQn5vSnYpDjHC5SuTdF/N6aupWYRYzExd
IUMuFOm+nw41Nq4CtkGG32zIVMUCoppS1kmrZ4n8T7XK9h380MmSUThGnK2LG5vK
KPwRKEPdA8ZQm6IsFSeBx5YKuVUU41ssSm92TllUkMPQcK5/lIhf6eRlgLlkHE5C
pTCbg2bKdDTiGy3OjyvtFO55gzW3cyCMzfhFffk6QIzQvgZBg2atfKff15w2RfhP
q72ky9SN7OzFzKYeC/ptSDgbUFkxjUKogrtB8Btn8jLllUJdpCH7mtXPcsGvPUNQ
eETHKhaQ/MdzagNy+nUsn5DwgKRUvF7QyxPG87CAwze8QkJHU2twDWlSUjbY6LA0
TzPtRATNRCpTuORYW1Taz3/5uh2jWJcfzL8iiVu6zsFyGvU3ffoHReX3M/45MovJ
fReBY1aTX20WwV+VbaGKczYI0l9yYhW31oinbrlrVTAZnfKTptMFJlIq119aBXcV
16Izmr+8UOe+JkxNZ8VbIsdvEdnyVka2XgMNEjSQ4oFqiTqRPskVf5NmQAA/0pFM
vVsk174D7YnoCkydppRfgOQ0mHqXSyrkMlTRbqbH+j41id45ijdlOQ/QAsPC4rBj
3+V5qsH+Sarry3rol1hpOLqoluXNn/IxVrdnkbYArus8E2+ZM8WJbcSpdBg1P8eM
Sx5VbQNs0gBst8fevRBv9m1425VB5pSlgof8GwiPGrGT0PzAR2xvvuaNWBtboFIJ
yxRm+P1dkYIV95jShODMcnGd7q73sgwMOQYCJqreBnA92qOfxQwuxPQCoKzWlsEn
Ie2KeHXOovOonZjThkPkKf574hKxsYXwIfZ8bO4O6pPUnWbRuywVbKZ12hQTfkrJ
DXDbg7kGm1r4xLMJCkbvLVx00wyTG8AJ6zrIZEjpMdzQ2QMCfvcTNUHQ4DhbgH3T
7aw1C/VntQeFjGuFnZt3lD30TPnadSjSikRy+7hPilZRpJIzW5CRBZ6jPB2zoqtt
inPcqmwScsroVXATnxrxYGxOntfuwJ0ZHHNnIjzeFTc/rb3HoTEKUhH6MJQxpuzV
b1Z4aVlcEaVBb0nZoZvJHaUVjpNRdRrItUL/Z887H07C1rzG0kDKM3t4Wm2VKmAR
F6ouJAw9d4n8WLY8HU/a9oq9yxqtpI3rlPcpWYtiIJjl8V1NqcJ8EpRODI64WK3V
godTpqBwjVX4Om158wC95n2ew6Ils+yvb6PFLl08Cf+BmFTLj//pDjH8K4VyZ/Wz
zlKzb9tzxjtMwmxGrKohjcwDkOz+VixPHx+ny8zwpHh5aLv0BO/bN9lBsHgXXB3r
SHBwmw+yiUA0UqeoIBYLMoo8tFK+WUNaqhDIFwnhs4OGpA818S1WkMYzBqU9RqdT
Nl8tWTfL52JU1LRrzVL3Kd5fnKynxkRjDdgwB+2bdNtb2Co51k/yiLMDZ7oq7VBT
p5GZi9F24lrGEBoBl/w1Ohoe3/jZgwCGctsC3uDJnqtPaFcHLTpO5QChka53+3mE
YlBDE/X3hub+odPV5a7DGNZz1uNj+P0F1SpHaSKs3cs1Q9x8XpmpOa2XU9RXRymz
4pXFEUlMbKEIT2OZ4iJnpNRDYn5tqwdaYyX/7rN3wmaJx4wCvTDRVWTuGPGIi6SJ
ChBkqPxamw2TIRU/Q9LgDCe/g2t6GZbW3UFHN++Bx9Y/JUCDV9wnEXCPDtxtYyE0
wAXLEjfA3YkvKr6CSJajrqMvs5PSTTDvDNc/117tdAgpiFPuOuCx4/D9JBZDlHuu
5+IqZnebY2DPIzqMsRVRYajqBDjeLIO4AImyeHzwyvAq58/ueLP19/TteqRmoHh0
zRjN0vI7PdqixtneGOMCL5xxO5LDVANElCbRwEFZLE8vXXMu0XrVe/fLAAwfyxsh
YKAF34s5JsSxxk+0W8bhdh3eYtP0Oxu56SxYpe4uZTUNMzhb4yxbyYjFhQKy9jXf
L4lHd5x6kDq2mu5+mhPINyAAbyh3lCUpUwB79d93qpFepqtIlC5NghR/EKoV4jTK
Fs6Nky9fkQvJUipYVU0JVDZvnk6NaENyFEVXibMiMkTrdAvzx4MvmOBqiRWfNL6P
XeMl4l4VVWiWemUbacCi8e1TrtrT3AEe0/4UbXSVV7IQ1Nj/Xy6pj5h0kCFDV/Es
+9kgsmamEXLAmxO3J0qWGCo1e0GiRE/ayaUlo8jeTVdE3xhN9wdIJDQ7vHJPQ5GV
87Whe3eFlSEvuT4lubC2dWanWlMkEs39n9FS/J0bE2miIVla/UoqDnS2ThBHN6R3
FGHD096rfIjHGWlUontiEtkZL/Bgu0Et7hufrwUhr27OAhqx9YL2b94evPo6uTml
A6iZ+jpXnngDmnlkVJAFsGzAOKgmITkEArZlKlMRmswS+vu0Dfg1NgaOiPz+QBGU
65gpKQQ6MI4l/WdfoeIqhq6AmnHlCjo7UdRQF1Maqkh+h0XHJ4JejqbuaR7SDt42
nh2h5hNIxXiGxOdUAyGFeytWH1Z3EHTcBDUZCfIHqtZ39jlAGv5wHX6zmPcqaEfI
KNbvpIPz01pnYZ4PciIHJsCOpGz7mwtO2OlO3Ftv+ZrHuEKuRqgItdvR3Juir2Hu
mnpwjCceiTQ+f97sSETXIHFGKSOBOF/+dCCi85QGHKuM7/putA+Ab8psbHb8YXmv
uaeQ1Pbwzw0g0h9Ej0XK7vdR8fD0uddvBHU2MFClrIZypqZazKJ27l5PhKQEhbwC
Kkocjp4f4tZHU+/Vi0wAmswlW781/jGcH6AdRTunQZm1shk5qPGhRPmY9rms6Ue7
eEoCub3HdRtQvPEy/dx3YyR2xgh8gMKlIR2m81n0+mOugLRaJDDtb1Wq8Kc6LDaT
5CNjWaj+9JeZnHhjuoyrjch0MHYBJX4pNuxtUieJCv717lMA8LXweJBNbO4obLXP
aeOvCDKutxJBdImHP8bWfgV+UKw8KWcE7vYo3mKtWj/NJEBkyc47VUsOitsSsoM7
jUcpi6AhiOCrO3p+TP5b0PpkPLpl6iMUqcr0wXuLh5CQnYENXe560f79wTv4xcJR
7D4x53RgyV6287HcoRU2CfiNOsnr4rGm+0kBwczU9XDV/QwRqrqTEpNtXKnmJKtT
Vh20jR5zw8ItC2aLKvNRs/DhCFm5oCTekanmiOCVX31RPGdN+z/6KzkqhrCO4mAe
sb7QpJfvto4tdhjLsN6/uz4ZRydgj9caE5cMaVYtY1D7GzDPBr+0OHZXOEDfvPdv
8nrPNIwBmGEHA4hY8ik6HSWktauSHpENHvgjbA0r9STIcQ0WN2UyMFVfWEAD/TeP
fDmkyMSiwOWSlr99yOJ7MTDERr/XWMBb+KxijC0viDWyOqu4pSTZxpX7x/2T7Rx2
nHnRXnJeiIpgl1zYPttLZbXtt5PuNlQBkZPnCwkLkZCcE0yo+8i4AyWslQXyfq3+
141y6e/rQAiUe+/E+vhO4CcKoJkLkhT5z9mJeioRmSvMNh7GpsvPU7xuqGEqjsmo
Gsmen7KPEYB67DAB8ISttOPjtEWegsitMLtXQyuOp771b5J4iOawv4rcyKECV/iM
1GtpzS7xdpeR0LEFk7c6x6LR5RM3x1MvgcPUaPshqENEEGb9oZ4Wt4+9mf9QCQiL
HBVArVk39CUVOJ5ixR3QJyHRNAWkc1pLVec4sMtcZdWY7nWdTBPrHLCGR3JWGmIN
jNFsz45DKJ+N1nARCnU98iqn0kzf+kUnvXwRF/iUrAf2Fq620Jyz06jZpu+guLmi
bYdJktKMB+rYAlNAMhANKFls76qQ1q370/9hiBaG7i6Smd+EYetqEzYUO0qBcQpr
0fFBvz8jtLjOgmGT46rEd2HKi/viCThAogercK1k7Cfz/ciaxIPv5Gd/ivxLnA2h
1NzTxITtAzLsA22/F/L9NFSGD4OIyH/BEuOIOi5OouNEqMU/6k6I04xrezwI/Brq
91NGpl9KUvktHNhyu8Jp/ZnFiL4BfuE31JleT4FQu9OSMGlw5V8Jt8oZJd53T3K8
0GCQBQBZgfLMMVKApbxDeeGtjHIGoMxDX/imerYrHtq+AdkOwbbc2VChvXaeugsb
ZRkrOW5vgf35A7vwwrDfXAMqfcCGhg4eqsw2T7PyZ/SCbB2so/UyN5kd0v5DUYOF
X6M5JeRZGQ4QWfL3htpsnl37qC0ygDmV7UMfDtCyLq4EQkJs2afjRoBkGz/eunzb
AlodbKDauJmfeNKgU5cK1GgdflDg86DI76s7uHptjKp0J+IQ2sbaT2J3L+qjVHbN
rqTwC4YeIafRXhY0rcAYMZksHNpnl3NNfTwUZYFlPZHreLuabDcuwls8n7gi2Apt
P7XxYEZ0wu/t6R8HWtmRdjOtqT3zQxaepLdf+q99P8Y+CS5LqLpwXk10WTlEb+rc
6bFcMkglHSSgEMg30kw84RL1btn2yaWXO3WZBP2KpDFGNiw/o07trYYst40sRx/c
vai6/vJfzduBXgZQ+LOc2cVOKu4up9oShBSnbxPGZnn8Y65R9UjVmogrdtLTzWRE
JnZn+FPTf6qs/LG8aaZzQxZTdjkaBSBVH3yd+VY/248X9QpLddUBf4tJdm5MrYRt
xifRUmqEYFUdDUaAuSOFePzhd/rILNCYIO4jcr5s4yVb+R6a+7CVCHhmcyyh4bit
XeSjx4zWi622SfWfcn2bMHcsAcZr/Olto0Bu0WuZ3itLb+fuFch5EsP7EL8YJ/n/
o8IZ8r3Xgi8zesMhHlFXvpHEgDaO9lR5c714sy3Iab7fnJkNlu6GkZ9XWMa7Xn2i
GZ2jVdwruT1BhRXfFdwkIUuQD28gjjoohTEQhhUjOye7dNcMYRASBQQavX9ElzX/
z27frkEKECBRYdmxpj2CI0ji2vPFFTm9CHnmCOS82TsjeDlyWTxPvpCJrspWPdGZ
I8INv37/liaTDmyvOVOeleeuNytoU38A7btloUi0QBjBd5wTWfcYb8xIPREaaNM+
4NwfCOR6/bldX+/gwHC0+iwcc1b783h4Ua4YvxmszYXxZBk4TErIDzFsQjuZwuKs
n0vpFWSprpnnbT8bU8qaPkg5hqGW9rVhcR6Ajx8rvSPUnrk5P1qDZCtpFKy9gRDd
JK0sSKIKLk9N/yhFHrHMcv0ty5k1wbO6Oxma1ZUo2Xgy6ONTZuogDOGSa/m56yo+
g9WlYewAxqN/++CfM4EZseWWHlzEYp46d7HxIsSIiZbIafBKU0VgrkB5r9NltTez
Z1BM7DQPrIcVHjzgsH6p3uWV2vpNeTv6aV7LiFuy+kyPgFR3TM3yUIdnjwvQsj+w
rXdD2Kr4Iaxtkn4L4lyOYQRfiNXGXGXiCoQaCx4a6pVvLcbhg5yCVTKnd+NX4w9U
OtTMnULykudmOkosSFvvfkVjiJdc6uRUrpONm8Ih7PCw1h4N0r0oz4L9ykMlrxYH
3D9iJN2LhylywIjYISAU/8yOCy3rgnn5R4aRDtNFw0UwrEFEOnPE+a+QXQTEArHW
b38EnOVV9JDFwZ+lz8/Le0fg3e4/0hcQXGsOnp4UKDdetPiVxTBCJxdK0bPK4hd5
UmjwxF8gRqykWjWpSKnKtcZ2cTph7qaPKfCYcwUgSsEdqd8y3BGFQicdxgwJZ5z2
sIb4FNn5NuB68HGKsncuRf6mP2RALLDbpFrtqoMwDrBAQ8dAvNoUHTltiKeJt7/5
dEeCHQmT18TKPxhUEIlC8PUKL2LszBBJyPIbv1HJXmoyB91HyX28n6sEnRaXR9zG
uZtmVB1pRKUNEfrB+8MarF1m1f/mdDhiWeN5MWNhlE6TT4DLUd3th+jIRCtS5St7
kq5eMu48THyAH2t3kXTe4h0LePVNnZ1s/1tMgH0Xg1L/3IMJNJWxB8+gam6Aofta
K80E5efxt0QJYXEZ2bpVcuGp2pSy6KiN+e+9ObaM7J8t/uyhf+Z+ZmttGccQKSig
6ohVGkFUBbnlqDeboZYyXxR9Dtjm+IXCGGTBywTfXpvqb+lVOrmJE+MXlOf+0+8Q
937YIHMCZ/auFDOZWN+KyzYjiQh+NKtwbZhkldNqi2RY0mJ0TlO/KnZ/iUR38gcg
ESafwsxEIUYmyv8XZ9s0Lnf8xzTiOla7gKxytOSKcC6o6uGih0Vuj8iKGiNbO7ci
U2NPuzGdfxN0NoAW0f5VamNcrGI9WLiKQac5HhIGV4tsYG88P/wI7hEO9fxd+kE1
VbT6nmqB/x0Q9LskbgqZW69tZbPGPEKlUe8BsWZP5udnr4GVE+ZTvhCXMiaLcgQo
aW/6ZS1xxr7Ar/3N75G13F2A0JfhJfEVr9dsI0ycMVoW+I/kEYSkY/y4ycrNXRgL
q4NZhZfJ/+xaJaywGgHAcKPDb0r2D41Mzuxi1J5FdUwqFdqiy+wXioAjY8/rUH0D
wiPDwpf64AqH6In9C4QfhFvIc8fAdrcyPKnlf/byhNlQPAX3R6R0nL3AHd3oYIVQ
mNN/0Q5RcPB7msqXfzZnd1hpTd1w79AuOOhDpT5FPkDZd7EZMwx++XzuYU7nmFql
WtQuSWN9yIOSWVOi/sHkCO2JVkJXFYAczJkTzlNsoqI0YmgOPNp3VM99Yoyb1KuE
1yQzYK+z+UEsNBUiaqKWAO5GSEamJolsy/2LUN3nR0Rzk5KrXmh07n5W7HKsfKCU
f5R8RnkOyB1ALrKKaIoqp4Dl+wAz76sP/rjrvOXyn/V9lH2GDX/994SjbFAay4T5
m4wtVFrdUolpAw4fzgorCfgD06Au+3LmOwrV+QBdrFJ9UkHnMVud32wPrkFe7It+
rVZHSYrTg4ILWEsGcRoJD943fu4yy++PbR9G9wlzQ3DbEBvwsYa5UXNT/ols0/di
wcunmGFRtUHRANVLUKtqimM5KT6E2aXnQLc8FzgYYKMMVw+/BmXH/qCe8ZezwzLn
FFD1Bbt2QF7fS/XgbYApTCU+v3oKxqxZt/oq9T8AToPe+SkLCGnscyDfh5IaATza
0rSVNFmHg3L3evpSCjw3/zARXNsqxsb3u47bOJh2viTp80thfqH6KN3UuWY/h4dR
YpvWu+Jy3MN8vq6wbEsnqSZcFxOFVDPsaX2jkDgg+XbGorzep9MdMHUkFbcn4RXV
vSSPyuVCxmDHhbmwnyGLP2v21mPAaRByarJDlnTYvbWwesB4xW6sXhZoDD5o8/VE
f9/pZSVdN6XX/ixz317nz9tL5q1I8OPNBCsXBnLYffKGGhkc/t+tWTmTqvjtZGPH
7DM5ioCyjbw2hGsxsVmPjupyjxnfLum+DV9qK1d0b88iZp7vhLt8sqs+LYF3vmXT
IRt9Ztm6ZZaeSUOkZWPK3S96A4WBRVNXD78EWmD6TCkLoS4w/HQ/GkjrTwWZjow3
7mCV5CjesQlAAiMtp0utWu1ZrDY6CWClBB16XjUIx3HGA//51QBzRsfsJQho91Yv
BNXp9o5001mnr+K7HUfl4nBqaauyoKR2O0vvnhB79EyH3JnqAE+GiX/Z1p+jcVF1
DHu8o4Xc5njDbKKVwrBlrD+WilJZONsq3KSBmqXvARybAQO2pXhpGQQzaEixX1RK
l62GLbThCqF/yEcHFKPyAH2vhyN7Xl5T0Hjq78rexqnUi/Z4oyZn3Ekc3ON453Dw
LSkF1kJvE9A4YW033IcTJpcVSOlkJ4JhVzzf2B51O20/KRY2hCNf/sFKS2cWuMSk
pmUbKId+ao3as5cQv9NMeE4RBLVGKXKzPL3e38Y91y2J5bk27i+NGL7EDsSOwDv3
dZNuSYbDr9bkpMQ3rei0w7c2WcjwshnuK4R3T6R4Y8cE1Z4iTzfy8+HThf/rsKOr
pbOzkqiJetFyn5uDkOu1CbOzVTwTD72eR1DBmC4TANkoY3wIEVJ8sohcrUrRyCzZ
pB/e6viHW4FiR+p1J4mD5IOcFreGbNcFwBzKs2rjevbjWEHaHBxg31dva47O3i+P
Z/QTxstf/lwj9AiqGwMW/Q4X73DOZfEWHxYLAyRs9n5uVZYAZpTxwpQ1s2Ogc9Vd
I48pefbMal6c4GCuH/EeoNuSgaS8LINCkq5/mbot5El3lE6WyTUohOitH2CEJgy+
Y5Hh9r2ZfdF31Wug6LlHvmhd7SrsvwFE48kJY9T5xqgBk/uRizjy5hpRTQnhnUUi
EGWCu4A9No8gZln2Vlo/ndrGHbpaQdQzw2dovcXb1bpRAcS0U8Ndmzd0yPFoZsrp
xn8Lhh26C9WfdaBiqBUGn6tYN9VS2XhYjFDsMsvlm5igK0sYCF0NgQuwCw8uvOvY
lJnZd5mVIM6Bd49nTS30m9m1bW5sY5uKY7ZX0/5TGEmjFqmMkvyvVCNX2rPSdczL
sVtp0BT4LJnDDi62LCwUAzt12CNvAjXhW4lsJtpEq+G5rol4EZVKFWR3gy3kjMA/
A4vvSnRmX70Sbu/LF2Uaj6/thP5CaGQWJfRcIfM3A1HzOpkA40rmjaxzyLIGujeG
c4ILQ+6a3T+PnXhmSNpn9s7tNbIH9A0JpnfRiL22F/mHyyKFmL61Yvq/GFe+nxap
otiHlBoWGFAwUObwrd8OG0zY3JUBMJ55E/IlnRfzwxW/V2Vv9sPc7qh6RQd7vMsc
qCxk5wCON/PiUYvawMMbyCxBbfa5GPUM6eSQ0ApnVFId/qU+efN5iRi0FWKPn4E5
Zp6CwlUifHE/UaOQhoO2M89omviGkA3FVcX60mJ3KIIAZWkz3borJ66w9QbBkJwo
ZnyxhfxZJOhPTdPl00H63s4T+9XIYcaJSHP3SR/eC+DhJ4ygSwZnZJ6hh30dta9e
mrKE0WWf1w5tx6bnTm0taA+IOAX9mi7aQanPGP76ErHY6jUaqTMSi3j6bgBf4/6j
GTOudvEVN01Mq4aG9XXHZ0wLChj74+Kaa1M9i7J14fIVRhEaZ5QlZKbnXNMn2YfI
6qcP8TGpziVNMoMVLzmOa8YJCcpWg3oI/pk/IdZqAFBaegprxxkpjL1hj7JFkSe+
pBfdqRR5H8vnB8gLdfVPbpuv3VT+MFqTOgDVX0k85I66KJFVyiDv98DbEI3wnY6O
5EpScXyZZaaz6PjrpMU6YTEGPpSVsGRmYWo0aZ1L7axruKptsNjr226nTIERKMRR
L93sx20rUQnl54vdZAm4UQ/0cNxHbu0AMNzrq/i2XiOvXs61VpiSA+cKzprON/ru
PQeo7JNpTpRNOqPQbLLs0GS+j4hI/suVGmQ6Xtsomfjy1lIs7YpAEelPUJd5peyn
IepfJ91mCA+eF/r3u8o65/TKvdJ14XBMujDjIChe2UCse4uF7UOVxrJD3Kkfh102
e8be1kjqviS1l22ev+9d5jSi3Nzk90ivzP23UXEmsyabkhI/bRuwJY13VBKLVXSs
oOLgYYLnCRYBCYlFoEhwe4xmZuVhq/J81//UJkW1/Y1ZGMxsfA4Ijw1zwCnGQJZt
GXPjVACnSqEYYyOf5KlGfwHZVB0eWsrGAgN2OPUR4OhSTuqUdwLCXA92NPSysoCR
bjvrpIxvgKWIiaUdmcD4DyolT5ij0cHIMERlHQgB698J+QhN13M41fyp+11OHxib
5rIYJNlmR4WQXSSm/V7HhxsoMwmMD/kZOPVmZFKkrNNMrN5Wh3uPnHSX9wUbNsX6
QnUx0gn3thPf+7Hv0nn2UTrWmfgHpmKlkpzr3VJr+4l18bCGZk1c2/CTd/ec3VYW
o9GCzJIOotER/mRX8UN2EgEVr35QHOezzs0L1/4mDWzIPDwgW+kLremW42KKE0mo
/kFoKXXVr4n4OgpSsJReMBHDtVZDAAEBI/sQ60KKoj1FDO5joWiV8I0SchoI0u3G
G1hnvsejhYmDIATxbxeC6cmkjU0NDWROvujDAu7p6MOg7zNtQ2zkAQGYjA+D9YJh
9Nq3ceEBvPJjtsYDOwbA0tkqSS9I7fCG0Sib5oGOK8JxdWCfOJE1xhwObsKMN4Xx
AgwmQID7ZeJEtNWCGBY850v6NRMY6kOWb/FUHc2mAKFsN3G6R999kqU/TqizS92o
bmLD5FHGfHVS9jtJCdEZCHmOPsJXcrhfCAMfKquol6foVPpXjDfV3ZorjufmCb8h
t+So/zbyo+K4LOkbfj8IlP8QppUk83BfJZOrO6QAA3bIHmFdV+1VSAx0hXQvehSr
GufIFXNSecdb83/AjxtX9DQ6YBg28SxXxPFbqLg16jXs/XmGHo2ZIc/AGsY66rFc
tSnhsFqc9pANx6eZ3rkoUCdywyJivcMRGucXrV93NkzIVxvRPfYvOE2vYe2ARcBF
WHAnLul04Htv8Z/dUd1Ovtexa1sBX4C/WA9EDCszNszywM0GCkyUWx/UNAkd01ku
sbaVoVyu3qUe2a7wglegk7fueLW9X77TV7KFV+eN4D+oYNBI3dwx9UFqftrbpvkK
CKyMNz9D2+TaRqd2WjZTnlaNmzUVaEp/UX3FC+EPatJzMsCr95eOQ3CD8YgdGsUs
mIs8EfvGZHOREFaRBGp6w2JuggGFxXd/7YotlAhUsAlNE8FQuM/kb+hYKgeb1mzb
/w8DmxS6S2SMHwV4kRDvbzeMr4r3hl/xKU6vGeyPxJejfxCsT/BckZYosrfYIx25
t9Q6Y7xDvahwCfrhmpX9FVQ/4zyjbcCvlq53BCIuzJkdwnwwUQR67QAjDMmCXfu1
v12Rl2t6UYr/9jxpYjnon5JtOBIe3bYekgj8xhxNHWhc+NnD4hnODKNyV724+AJZ
xwnby1Y73+ZIZJhNtG9BXtC7kmG7UoT6pue02t4/OwSgH5vqAAxWhnb2wkCx4vS/
Q0HdLcQWI5Xbxhq4moJRPz3ImUntOcLFoUAhMO1cZBXN7DrHZ/gE44Le8clk/otC
1Iqa4mwE94CQ79Ds+JQsoWBMBeYRmw7byvV+RHtBX74sMrKxjvYEGgocPilmEzLD
CYbu1SqQh/69+jGamI/Tz6Su5cm56oRmf4rxA+OyBohz8FNW0uqFNLZkW6kerD4q
PLixDfOO3ULh/DkPD2RJgdo1AHRFImXGlgXEG9Dg/bs6kaUJdm30y+pYcxhuv7j6
nfEy0PX4UMwK/KGkFMoBcF2MEbgfARtxR5qRqcU9BTbYlAxZU+lWkNh+e0rec2T8
0YZDT02WKdwZrCBy8fbQl0kCcqsKfzxK9vevKBpocpHDQsI/WrffA2bSLIa8Fen3
QgUl0VNXws/G5qFSKfmxJE7caRLmY/kxkO/zOOM8tKyuwokafkJ4WUegIDyCXx07
WHJd0Cwr96LlBEbpWfKQzNi4QL4vo7E55035l8QphAILlC4RixSPuL3mtrUqC5Qk
WDW7KOWJ73nj2H5VlyJqDmQoVPIwfMHvYXJDTMADOD95EMSuCTZV0tULTw/p21n3
eYNGnmhX6jSvmW7IrRUquoMDbG0qLPU6A4IQMHCL+8eUUkoMSCksJEsX/gREM1ou
blhE4rqcQKee9hH0oIs73UFvA1fEIW2NkGa3gablzMkdZZWzjdCKCCI4BK5X4YfD
dxGXtkkhrMEja/lt0UVZoI+4tNppITyGYhA3H9HmKb2jXsBwkltyWTj9xcCG8KfJ
mRhaYmqjVxv4JfZfVA2jKmPrJwGiWn6L4aOyygKjqjxKEiPPPROs46JvAuvYHx/A
FDPL179F5ATy8ZSdQ+L04hpd1+fKDxbGZ5s6lF7bEhf0gYmZ+lMw67VCnuld+Ual
6ytAwynAWeULDOpE6A7DZHyUTDZb74SxMncbjhYs2POwmXztFhqe3Sfk3SxRbewA
zR2DSSZl6ci20XAhHDZDWHuY4pmgiScKsAuuLRnh5uJJmh6p3joeI3tDvQZXYwUn
9SyF0GwT5if2RzBPPzdlH2nGEQBGAuOUqtNUWviS/UIUY/lMtDp6mUF1qNOEZ08T
GMj7mg1FwMqbkrOQsQOhGwmguBpAyj68XOJflRp5Kg+ihjGvMHrngSkU8bVB8qBv
JhDrmvAerusu/AHRoK6RkSaDBHRtfNut9xF7lPgi2pCGIUWP5f9aQeG7dJRFb70y
GbZA9O9Lsxz5WLtS9a+NmeGKzh4lJ0zeEffW3AaxRZGnDC1iJywgtO2XDoiqpFgg
LqsomG0Nb4Ki1HgYoIGjOMaINZptak0rMy9YX7OHNsv7IAw2pawHLV7LqGBobq0v
CH1enaKhk4OxeL4X/qgwbnA5tEjuCHSG+NFR5Y/t7X1m2kdhGDgDqwKJeej0wI+H
pw0ohg0/eLFfhhe0g8IR94xa801nI0atgjiXRZ5z4r/ye9GAq+eCqX4j3ZCyPBYP
3jxC0E3Byb6noUMSvINhoiDmI234kpOpMKX30LlmpttjdWjSlu+UOw4rREQ4oRLH
HvfwKKgie6/8twMZKItmty1NDKFdspg7nmP4Vp5bhi1c2Ovv9qsvy2J4srK46Go7
Vkmxgbdtj2c411FWa3P2I+QxD+O3YLXj35sjGArVxLSrUHhFuMflryBS3sRoZ6jK
Km7xMukiw1Hg/MLS84L/g9o3gUShCsj0TTYdmLO2tqEd6yOxlz3tCi6Cc+hgyaaB
/SzMDWj9KmviMIm2ld9M++bqFMy/KosZqDovX5Yhena/38iE6Y+XWaH5RcXxy2zC
OpGtUQGw27IIQqr+0FcJ3HGD6x9xso/UOrZ3n8Z5SNCYJ7pzr/1q+9ij7sBvB+NC
ZSO4/8mNwDdzeBsOBQMVbQKVe0KCi2yb9PqFE9ZuzU1wNI+EUZmC43z64TtqR48p
3Ol1CYmWH9H0huj1TSKIwM2KgXA9QXspW7FZAzQxLEbNv7Ozq3BUnl6dFkvmhjiJ
KwYH3vkfj0UPDzzZVRUjdNbGIRieUFuR91+6l0vLSLC4gGVqa3KpO+xGsc9fjkvn
BQuDKAn0mwclx0tio8ilGAj5Ae91jJ19EZf3gnYZkRG/XFDztSIJkoWtT4Tfgj6A
CHyBqVHJhT+YRVSwQnpK15K+Lrus/j9IIFBshzWVWq+l9/oYeDCY3BLB0Jx9FFZx
kfJq+WVSjKH2LSX2qNhLP1swqNTwocxcv7UGmwJayXJdGP5RJJzHbs3idk15IV0G
yev+dEA5QFgsSnMUR31vqIQxHRv5d2dcgeIXwkd18MysIEvgodsoL+bQUuw2IWj/
ma6Sapzov78sU3x97hluk0oepbxBWB5wsdMnRwaiM6rnz2GKjjnk01/Fm3NiCYmr
7BbuP4ZM/mqRLQUZE0hFXHgHLDl+jF/n0ifsnztHEJOa27onBF8SgPcURXgeOu/E
7FHUJhH/eT7tTK0ZxciEcBTXbQ4Qz0C4c8qYhd61MNg4/iVs/88sdBM8XNFHeZXy
0+INP3ARNaeSLzA1jv3cj9xZot6EBKIVlFbC4Yq0Q+wIEpOS2TafOczLTtSGsAP0
8e8e3Z687gxSYLsq3bl0iBMZ1ppPep8LaOxIBiOi8VtqkpV1PrlsO/pL0nqnGC2H
ypUAFaTcGDlPjwlbjL5/fwQJtEo60G+hKG7ndgdUamQtC4vaRmxhv9Zk6dEWeb3S
AhhY1o1s1a7C3aDdQalK4CpKPJqHzoX/Zl1wz0S54E0JxQrYBqrld2tsjxbDUvo/
SgJek5Rn5nX1EjXHFDT6FdqnfyfKPW36My6Yllr3yK8L6nQjaeqvkWVlcrXtFKo2
9aktu1NOuMkcJSwt/4euaAtBr6g9GfJGT1P6zqeCOR8yXVb4XsJW8hmVchWpISFn
nlqvWgH7Drns3ChVP2uBipWc+JiVx40DSHNKPUTq/ZCq74+6vqvvk+ufwlMD2Mlx
+nW0aYkLL5VyOqeG8gYed5bE2fmVU+S/oejJYiGEcYya8gUaxLd7cbzI0C7fvoN0
7V9smy8oO4Zym5R8PCQn9N6I2+fpOKnPormFfzxJhfXZ5+2cmgt78siYlK3Hpsbz
0NzShzfirurp5cvodXbeFqt2zuYqRoPJdEjN+9tTnVF/X6Fh23mFoi7WUjLeAbYH
vX1KGug7qN/hnrLNHNepGYGn6jv/qZ0GGYnZ3nP5mMNTvOFArmAEKGeOMfB3hXRW
LzZjgmOJEio+hZx0JGOkV9dHHAmyH1PjafUD5KMsRscq0nT8xeeJj8rXxnKfGv38
J1b5DeW+5pXMk3FezaaWQ47uqh7SXtNYnQ/DjKy6nFDFKoljXGRlkal49ZMktR8h
UpT9gywJ+qqSx+eflryTOmcEKooFrQIND5xaiulH2+g0E7vn3MqH2Zcudi/DuMe6
cJqmISW0lmJSLdyeXTtKMSxCuw2a5w6lKtNvf06ISYEC9iAMHBop8nCvqnWJtZQM
NaYuVqm8Qd1rjBE8Xp9eeK8rjU31gGpucmN6qMFLU8wBMk60X94RJlujhCttdaLH
Vl5NjC+naSkOZ0lECXEqt/wueea+uJGEnEyt5aLgv1+5d1u5pDsvxkk5lFfXrZyf
zT3nfvaEno6NuoYOhIvB1jd01z0A1F2ALkQ1OTu4EJtSIzILxNxSsNeHnJ64PlWN
mL+WFdWqfiktfrjADukSqMgXn+prgIjckEy65+pwNTRRGmopeZuCSNXOle9rjWeN
loq2PNbdtpSwYaS2tQ5imhLbItGqVVwjanqbzcyMMWEJMcYHGtyakDKCqsca1dDm
2uUWoKkNBFBpYzS2nr0ewe0k2dnnL5hSG/Nbu9fxnK+eSr3LvroP999jEphsM+i8
NZqXgqM1me5Dz/LFQHdmo0GIH+xpvGVmuZjlxnU/9ybvpj4Zn0toy9EQSMFV34I+
bkvXssJop9rt9X0MkFRasCAOwVmrx/SFjUzryKzKlYG368ucsMASzBxLaR24sOdE
WLlrX189avjaNkCttdfFyM5IlQVbw51J+3nmlN9MZu17Tn1XBR49VEbIbZSAQ7/A
POy7xHjUy4/wWGxTz+2KyxIAT6DXHoi4YujrWFdu4ys63ZlErs9wd+pe63vObZQZ
cc5nY/RPQhKNuzp73IEH4htKcVqcl89IMOQXw513Gi7vz+ed2SfW+/4uAIsHyQid
FJHssOkd8kW4atBmCDVjio0hnoqdXEPHM4hL00hqriOpwb26exSqecxDr+pri2Ww
IU9+TeXoBiNenAZ3aOBXF2d6rOixkZmDceK6wp/e/cysstXE+CeakpmQIcZlY86q
Qx2v4CTPicHvAnGSFnLc5uqvyZRK/cXm5m94KT4dmwlAa/ZFa89hPG6omZkdLUbb
4I2DDxs7sAPT/IvAxFftoedGLO7p6Y9uk7QIS/V0K2siUhFgpUQVTfZqZ5Ur3jxC
1HFAU4qsJZ9F874EBMleiseU8udqjtse3BTAakxWX759B7O5EJkNPXjJyfzL5S6+
iAtYYlPZy0DO0Rh3g2WC9GcE3gb9kjyXVioR9XgEftXI9n0YUPqDFQFVc/or6Aqt
yL2lqEOISIrlf28akDJdJR2o5ClRbjKsLA+flMRbRg4uYXDHHz+leEl0VdRD8Qho
U0yGgAXjDWSfG0dl61Sn5TJ0GbYT2Z04d1BUV5LdXe+uosUngnkqWfDQKHbOVWkB
LsMr6I6i974YB1j4zLgXqY0H1x649QQvA8YSwHqRVV9VM9fS2BNJABub4Iih5UsQ
2RiT4CxjVf5JtYgUSFzCLsXLJH3v5XRilx6J4iMPuDLjt0/m+a/msWWJrDaRk4S0
iDh/LL06e1iQloLvzeYWj6OrP502R+c+F60jV70nQm7vIB1Z9IebSn7Ncaat4kgA
npg0+Ltr3S+H3wgUD/jefklRYpNHfuddaOtAQ4XNgo/boqvvlHTsK8DnHLWE85Sh
okVycy8cOTXLCTInaA8FubaLi9Imd9TlQTYxL44KKDPPvLBB6wpLlulSKw1ZDo32
H2CSFziv1ygIHTEEOcSO8irbqq7PbbauXLEL9Ey0u76PQzxaSQ3u+58lFhNwlJAV
kd2DlVhJXDci/uN6QsWtbkreQUN2oCJ+C03MZImzKKkwivaZWLYUVnd85JVyETZl
YHSfDB8uAG/chBpSjqun63Mz93ysTL0/I+AlRMdyB4fKnPeI1f/GoEAKJ8fb5amO
Ml4sHmxMLyG/WdltRB3fBxs8k5+xbaXLsnIN2FqyPkDj5Y6ed1VFDau0ombE19JG
XELwSIMHFR5RKLQsqC16ygK1eXmd3uvSuw8XSyMNanuXPQvnjh0gtwdhXXfkNbud
kiUmi04JHLdPnLYclFiQEOAbFNAxkDfooivWjxJSGBsaZdla0ZBRcpLW4sLG85c4
yemU4nx+MXV4QT2XB06+T/2s5EdMSHy9fEnm7Yl8xBv+eGt63dDkfkfb5GOJ+UVk
OEHmK0G2G1UPVtXj93qqxQC/ogf9pdpRvVqMlJI9tIYN1DTgzb2h6m8+dXs9fHdy
J1dNN7Rt4OjITZeTFgc09QKOrHpIadhKobjYtdcRN12FxjX6dOyfoFghvO9thxFF
WbOgqg1DNXAfCkJs/LghLs8/bI2ftpDsNiaCpoXRGtvr6mV0r8zYGaDwuzlUmCi6
+Xeq19KGp6OoaDJMaXv+DEetFyiYPwt9lxXeJy0kwSRGkcvdbeKAPojY2uxQQhaG
mqOPjZgGB+PP/2jM7V0bB8bvGIDRHzokvw466ZAZ6qmLu8xPAbnm5ADq2+MJef74
4lqLO+Skp6f9Q3DLNhkte3zqgLkps3RP9+yIpSj6KbqAIR8MGN4XW6achnhir1Tp
ENTLEIuSIbWpV7LH7Js3ZdZ69uWnAkME1bO3xpwhvOXwPDOju6ys3Jsasl6VL/8a
kds4Eed2tYFWpeUKU36A8Sr1Wy3tNlDKVETOU6yggQHJoMoCT9ICrJESW6rjWgBQ
rHpkJd5ATOlWQ2eyxXCi+QztTmwOpGSHLwGR2UDKzFtFWPHCKxzDpr4esWhE7+yq
97OWpbREFCKk5S4tt1WuJvFVZ+ohneKqc0MtPgVoENqBSMrRDj5L6KRiMzyloYUe
nmr3lTgae8BvNFls4vEjGLINpyFWGlAqpTnZIuOoKN/5zVt+uwlu0FaKJH8Fd1vD
VjDEps3ahq5Ch9R6vGrrV1fZwfBRrFKtpcylpQ6eXbvICwj+3HkhdW6MQ5UjLB4X
wageeJYWY+HQzoLAmPyXjVY9wNJ5FmgzKeHhDET8LHOHpvhClIjcPUdlNNdUoSCJ
mXjrfvGCQozFEo3EbX5HbBGxjLFEp75jrlvC5oiZrZEjvHm0Qx7OQv39Mn42+kKA
tvqk2a5FDwhtLvb9zcK8sz8sWIjyr+Y4JRLGOX3qlpwhSWsiKCcru1pI4j19vhMy
bBzy0QmSfhodqNPIBX5K7m00Z4yOCed+ZqMKx+Y5Zsw1TDC++GoEOgLEOnK4ve51
8eQek3BKhiXTkQ9ridAUoQuZF49eWDt9f2qQu36PlZj3IU4dciV0F8RkYMp1WYBa
Ur+a+i7Zuu38hgS/7GpOG4ULvC3tQT3BnsT00tO7G5cDe4QVw6bTkGQCbyv4xG2B
eoW+eGAVrhhVlSfC6GbMB6TseFS8Drdnk2ybskhGS5y5br1Uyj0GTb5+lOF+h3S4
l9cmpaAIV2G4Sg///VlHyzPtFrbDEppaHrlIsuYlKN92MrZ0gegkn+oRN+kw6QrJ
QeEAeh3K5PCx8ce3Mq72J8V6ctha6g7voGx1wG/Sep1UefLeoNflnoiSoyqZNUhp
kqmNrTGQGP1Fvf7qF5nvwlGBeRMr2zUwqQWndUnIdxVBA0dqTk3Da9VKFDLjPFwI
mzgd7evK3iLD10BHoz0/SWHeTYyq/1syq/jAqmjBR/XCnftINJ+jXN68WvOBvCjw
c3D55cczKcurQ345XZwDZGxClICx/Tw7ziYnQ0LzyoPSYWDUzADWL2EaKWUogsL7
iIRYAvnh6rgQDjwbB7T28//Hz1Y88tkAo1sgJ7ay3RJ/Ok4dKp/mopnn0dmVtG4K
7SXPpaEdSshcShsdrrROQLlPvftM1X44EzmuTg9Mmeg3Qej5xu18wqp4vzpOO3pI
wuWB/CuTAqfArIgCfdupPC6hzuzC5jJ+m2d+tFeJHaMhm6esGrhFsz7fbSGfN/Bk
cgO0Lc0qJIY/gCQgkdQuXj90REC2DlanUp76SVRQiFuTr0iO8ZQr0ts1O0NleGO5
aimoMIKDn2oH9xPa26ewplQpUhDI6MYBE63sAXn46sC9/90XQq2WCV225py/+9Aw
EGi0KVszxDhClzQi7KjRK9NBAxkc3OKZFTB9EjkCtnBvsfXcq2Ikigh3p195Buwk
fUj3oNhIBl/y2APiPnqMM9y7ccedeSGgMQ7WbqNOvUGxH1I+gyk/vWI+5kaicQai
b3annl5vhY26X8Ya6Tb5lYP+FntD03FATtcCycdfLpeUuQP39e9BdW73mi6R+4DB
ygs7Le8tGUvJZNuWfJebSDl7nYkoqnBonMhco2/hhNjcf2Bd/8+YYmddtClcJsps
MfAjVHYYErxd1bD8gWeiLavAKCwmWC3vi7yn1XzNQExjOWLKsbRrbggxjT35/C8J
yXpLC+wSuxOjz5nlH5/Es3jZfqLpK5Gsn0M08rAfqPwe/kpg5mQE1igsvI1lv0CO
I/QYfUU03NbY5VcMRSzWMmfLwYRkoHxC8l/HwyOpHDVcp70hxevZQDh/3rLk9rUI
R9Tb4kWLRVI0mqAVgNQlLRLIxVhMAaxMJMMBz6Wp60eDKuQPbQBQBgFR20+6UHRQ
ZLhOpJ9LUDym1scc6Ht2twvIyy2bplRi4vvXAvcV9CBMLcl+qRhhdmYFTUlSLe3i
eADpryWRGs9QZ8amSpEN2lXPeRsCtyQfZIGfturezHqXqMXNJdC5/uGGG8FS4wWS
0OVTsTyV63OOC0elMJAyNeEiXTnxCZKd8B8TOTuPWBtWi/BPRDPdNPqm1dmcmAIe
kvjnwUJfPaOktY3Lh5rXxPPDKFyUKboPNeZk6UzkoWqpOwslobVO/zYWUA3MIrFR
lqsxrv66EasUEyJpp+Iv7i6Pxt1Qa6EaQ68rnciDpl2SmwVZ+wIlKZ8+DKfGWbZ4
MoQ7f0jo7xF5i2mE/pBqurG9xoEoKpXT6vD5eYvLIcbBg9xgByGOf5H6jIu8hSOX
uoiJd0G+0QCtNOasIWMf/Nv6tPmQcoiCLVtJYYI168rysMjmWSrYpoVreFesfSbk
Qh9fLO/0EMCLQVzSnuioGF1E5mVzz2OnKpNCcYR7kFS7FTj1r1jx6/Jf2GEc5MMT
mfKK+UderIwr+WZeNV8NzY+cfxQjZwMbONrz0UgH57Cawd3OGsOmNfTeMMZfnpKz
miO5NeHEDV2Aptd4pFjmQsrMB9hKg8Tvf7eiZol5RHFWg0Hpq6xC68samUcO0zlq
yFOuijT7WDbmKGNJJDvunYDkXayDWXv0ypK11el74OBslTAKAVXzUfSJgQBgnaAv
WvjM3E5iPLhPJNH8p1LbPXIqNf8ZKAwLS+8cMupXxUKDBj39QuNOCVqjmR2KywFp
1rvmfDE3pW7Aqm7Z5xaJ6wbh6AOLA04/2g7WEQmT9IIRhgJV+OEsT6m7NiRGM9/0
LIwIZAXHj2a18JXQtrzuB4tZheMYp6OmW3clVeEdocH1Rc9pgRJlKj9xc2uzwByF
XDAby07EjLC0R3gaw+acU4TsoW3ZIDz9StHLyPdXvwg5ERpVi8t1Q5BGK8SmEPGP
AvdxcEKoBGcynQWGayIZx40GY9nHKIDNTlyaZIPjOcPkd2sU3zLTP5pWOS6wTWbG
G2rkKPpp0Kv9XWjGivnMHUd134XxbwcQGR/Uz25GTSVenY/wjchOSds2Uz6K5cyC
tTqCB4LfPGhrtKsstTX75/M/No1UuB9ghSjQ1/5Pna+k62wJmxrfNU5IntlPcv8I
4s35DMl6cVEy/ZgERYpO7cbjbi7M0I7yLU96r6viT6TIRNilsbJ20ztTTv31jZ9a
EtKyauPlZGQrrpONeYvrdY2yZr1kNkMMH8Mwg60bxLZvPx6K1Zwm7m4UB7RhaHhK
42cu8p12c4hh1Zr6MN20/Kp/5a0IE7FMq2a22d9rLjYy0EF+SjBBl8OQ/kznc2bW
revFBh1lE5vDH5tG0SdFfoMOz4+Us4Aai7mOYNPSS9DEw+VXZiYJma6WDQb9Bs+e
csDAz39dwn0yTO5Sq4hqcgDVatWSR1afBU3Zps0x9McZzD7x+2WAsFd/ufhRjnxY
nJgJubQxnBOh9/j1JBEmxy/usXWM3xW7T/jX23j9kPPUASH9DN+VpVs5NORjuETT
jREdvxC3Nbxd49gB1BuGDxZZzqEKEPX3sq9GwhF8NpOz/L8sN3JWcv02w+xg2OsC
2iRzbUugPX9Ag0cAuztq698u7FrlvKHedhbizWpmbfQoiB15ZdsTdGxY4zoI/nZs
gjYH0K7jbQA17shGNWMrXyzH3gDK4d52eNTEZKpNymEJJvpLTi7JKf0PzdCjG5Yw
L2inrO5ULu2YuLwrSt7PWA/pakRDuYu6k/iYC+/t0i1WkrQugCBLtoLdfofSRceE
k1H/Qmb6fB0sTp97efE9FXeI5fUVM2Lnx3mFlwFVm/7zL5nGIanT8KKS999QUGfx
C/3G5uuEFHZmthFFnnqchG/aNZLqhbyTS9elS4SNO/pvX1wj5kxhRZEgDAzrNHw5
/YD407vCWV+WNlDGsswadDUGiB0T7qA7dk4uNxEb4TnXK9PUS9CUDqqyPpdtiVQc
GzM2MCfNZ6gnFC8pKSN4msf91uJl2Axiu5n9fo2L9pbF2C7Id+QpNQgLBHc+2lAt
c0VLtDL54gQdeJK5BZoz7GZwXO3sKaT3w7a32z59Z0D//adMb2cnDLcUqqR9GMQg
jmyQly6RwYTFJzecFqRU26alw47RTbHNUBivo7vAPiCd54l0hGATmei9s/1fcANo
xNlfQCC2vF1IYmlphKm8WP9vP5FCHX/zRpSeYsIpzFgSyeqqZZLRV1EHsCz9Yuze
QcvxFdEZmpI9JDIft61GSq/LkwxF9tO5sjLBSwYoEUKZwCVmjf/2xGc/pvN6BXW+
yjPm1tyb8TxZ5rAmQwFuZ26Ype4CRdih9GrBd0/XZBxfyC3cDrPxEO+/lJdgnj4g
3qVxMwK8TKXLuSh4ULmf4BDWrF57JCAootD+7gzhdQ0vN7xv64rXQpdiSYZGZLYu
cqj54RlmWzgF7CqshdAVzUzRnIMv2o6/56H6peiL4drZDlY6RtqLw4iPAXKUCebV
M60Q623n5NCYAARB2murRixxjPKqazqdExHpvWyHgcp1MtXiBCjZmRZvsmDgfCZ+
IUYWuKwtVmkYa+rU6u+/BAKQpErBkK7XqrG1m7NkVBa4R/DaBPYb4hhCSJuokdBv
bbr7zeDy/Txazrf1JfZrdm5X5adjdABSsmrHaRb5b60xNsJbhupbgBHR1sfY7LWs
W22vP2TSi62a50+3+g82uWya+psU8ZSrmpWScRsb0nQiQJ+KsfCoQA0oAslLVG/T
mr+sBGNCIzTgRnACFtQ8kFsr9p9HChtpTSd5+3kyqThht2mLwLPrfwWaXNSwtJ1j
uyppX6SQnDb5UUcdrmtT5cYxOP7BYs2fWZfddkMB+t0ttPp5fFpnQrlUwHgdJay2
y3x/BPlDsk1DZNvUiGRZDlojgqrAw/AeMYoKAefmVbALAXchTbuxaxU2oTBI9aAu
K6PAwFUZcZauJBTwDOxGenF/8A53fkJwqgiLBiDJ49ZmU6hdUaZwKhpv0ACE/OPw
1T08OhNo3ilRRy63X7eJQGwGotYTHCkm1Z+YqYcbcj/DW3qiJ/88wE3BgYsU0tax
kseK4fOrenw0/WzmzlYdThOnUjMyaoej5oX958/Htynuht/XeljyrxMWixxFpNoz
M3vueVFQzHo6pV5RhRkb1u2GvwBCVYSj0bHmXH05p28dW0v6UwMQ5MtqnwiTuvRl
VnR39PIae7pndi/V7Pv6crZc5M9g/wpmrMlWtR5u85bTQp0HDF5/FFFOe8bTXB5z
IHYaZ7EydWJLZNb4ut86HRjGqu4LRJBC4L+EdCON3HybsX/WZe9RzcL7o8EQsqiQ
e7zQhv4qYshRNa10QkoyXCvrR0dkzOVP3QEZgvu07I0pT0NHeuwM60gX+TuvW5Ni
ApBXWSaeTmdi5rOfnuinhDXhxZB2H9x9ZC0Zay24i3kbwf6A04pQj9E8bFZtWZOl
8P0jGJawbK3c+rTmU6UgXYDkdC6giQoDJnpNGa2Plpp6CVE4tXaoinGiSoZW8x6Z
8BUPfTa3eiTMgRYG40jfNHJPYEydTVuxmFlcfIxZaRgX5e1zF5H8RRuIfWMc2SFf
QwTXIBM48ZZlOcr4S3TWzJo9wLCcKyCaB23XzHqAYGBLPAJXcRRd07vOxUXah58G
WU9130/ZT5RiZ7FtIOst5CL4OpSd7LPJPojCFmTQZmsZmrNE9XxZG31iASHkek+Q
EySf63LIY1H+1ltU3V1MH53ARemCMwcxYmtqtF/TnDdduGD30NjWbK8ZqdlVAys1
2Mh4YKfEx5cr+XnWS5UqHNmXPZ2GZIrtzWXi7Xo7FtZfXcfKJD1WQsgJbuBTKnUg
ZiDZT/q/lGS/FnDxb1jXA1Mb+cNVu9/3IoJt3urjd2oxLR9nzF0MLuPvMSzJqfkX
bZ30FT2+TQaSCz9z2Dsfr2KF36wfSfoU7qwEUkJLj5t+0nFbnNewUyj04LbIDxdL
3fUrKpPOBSgnOWOr9zBSECkaO7fpdrZy1QfM6+GDOTwsO0ez1vDNZT0uQpJ0TGjF
T181Hqen4GIPhdEUGg5I/DvHgkNijMK160XJ9wO/2Lhbt9RmVu05kwdVBAA2kF4G
jfjluw3R2NvMSdQsduLP1xAFg5qzNju9nfFjIbaTyoZpyytfWte00y8ygFnUsMbS
GrTLIW3w3ceIi6grZfhQOjvP1iJtDeQoER24+jF73IwLLChsyVyB7XHe1IhfTQTj
CmcDJw+24LjQQCOxkViEBr79UHZizDbvuJ2At5NbgDirTUGNkn+zWoJU3R1mkMXy
309tD4m7ViD4qJTosqYO7cpSDvHPw8YtN5SkaEODsMEsd7RE9Br19EqqSxa1ErXw
oeBYJ1QLu+2QTOATysAWtv6UGTOoMHB43LLKupsr3oQiqgfds0QhZpacnTFbYWoB
pp3FJD+SXt/9G5RwotOzLxqTwbjIWw+cA95Z/m6VMEseB9vACWr0aG/YzY1wewjr
hj20sQwk0Q3OpTXr2XkCo4AnSOFxaWgnjVnsZ/qLvFLJSFA9GF17dEXqqaGS6TR4
Eojxl6qc8TDloMZrSdgLgg+HGUvFvcRH1b2VmVPi7ndNViHYqv56LmnKFbPH1yEu
hRS2t8vdURs/77QkRN/A2hTsxC4UUBiH4Z5jxAfkTPWBFyfCd6x6cqkMrxtDr5Dw
qYYH+6c6xWgyz5twRyahPTNTIUcpNy1FK6iiCBqYBxlr+EUE1P1DKvNfFPQcrjfU
mmILdgzfIHLuRFnVWzTbEIAXl2nsCcy+w60XmYz8Oy85dxFuv7FOVp/hzke02Ij9
bIRcbcGGtCVgR6ZPYHHDgmpeSE/luDoR2tZd0de2Z64ils6I3bvIsBOfjvIghPH5
pnFfqT3tuiLnf5iNb6WqjH8F/OuUrYLSxVbN7DjPplm9UwOvXHVnNjhsiZmpGuog
+BorXs6Flldv/b2EVa1uT8Od5e6YmvTCHhO+PlcN4N9hHqDucWdlVXHVk9BXuQmX
ucYW4+NTBJlF2FWRq/ZjqmyLHcWqFfjSHpZvJ510S1BPLODuJcGWHO5Gq80eM7fI
QYG1aa531iA/R9fTCazEIjuX2ygs+7asRs5ziPqsDW1sG6uH88P1O2IJpssH4+Xc
J2Xk8eItx1ZzT4OepNzMSIywaEqmbvh9Kdih/couUt4AY27pkDWykEQGPq8OF7/N
dI2CNlLbNLoHRPUi9EZ2F49HCVIsvm2hFzLgE4nrAR/3/oVhLCQi3abFnpDTKnHB
HtXuxaWzVQSqiyziG5ePbquSY9huxCs/lJ2R6Ixl8tQWMfMXs+dmAQLBnK951UG5
qPDXkFdBKwKCdXHQUVxZjE4MJugO8A99Xvz2+Hk+V5UsQdt5Wh9rDGWI1YJRtYKP
voblG8Kq3/tzJsKuw/1bT2ymEPn2/ywplP6Af9bR7ycw5fnMlNkge+chnPUaN/cn
OU+zdE4y/OmokmhDOhF90V7fCMEQeFjy1NIx+AhnZjEDmcnaa6bYLPE3z/lxyYr2
pqLHHMc6nwHtUaW6Xz44CvuhEgYuUySP4NWGPCFPGI11S1hQ+vqiaP4whUhPeDoZ
+y1iBPdtdafbkcnhOnrRgE6ouTKkzO1HvIzldOACp5v/0/HHqmd1i4l1fszWM5KZ
i3aCMmGmb31y4clhXCQaDw4uXAnwMARtvndkfRUnNeJsRJ9Uddk69gZJ2+erKRoV
BSZ81ruqUrAskmFwF5Pln8HeCpk2F/vr847FR+VK0qxLpuByAgUXw/Z8YZf+xTaL
ZKcg1WEgM7OAoXhhUQ8nAEVxgk3VCYODqg2yqmujwJPr69WW7aYWBBlFi5QzkNbT
ldBf3TtdSiZFfIVNqDOuxn/dSiyQUZwZzNHRRiP58+7vapUyk9fKKRNH/BDncXmf
7h6wss3+V8oy2TFsqzi5dpbBKR35Sv86Yglo8AtgDrAFqk8ljmPs83YD4MrDS1X+
Cqtj5DpGSvaLp+YtwuWUgYL+zSdB5KH4GY3ztl0G16n7IPhywZxblf4w6S6xl59Z
81I64uzzCDxft39v7DJ0nOXfTEoAxf+4pCLf35vHKk4y1lmoIWCNgV60eFh0lh0Z
3X8r8SHzZfhPXnPJLqYQ9+dfl+dufPf1xVkN7JV01EEC9ey6hMMIRig5AzsvJoHf
vY0ful/1mMJlV7tPYiNeV2pJGyLTyehVDAzv9rj6ZcO13J/SbxIXhIqKm0Sj3dta
peasxiUGUJ+6JAG5d1EBi2Gix4Yz5gecYE73jLlMA8logjVI92q+xNLFY6/zNu21
ym0K2u6ueHC1hzRdRDpa5UWoDeRpjdCNSsktf0ARxaEIncmwmM9YX72rzBTc6LWQ
2b2HqMqLMpyL628Sn5yi6Z2kUED/RpaLry4N9YPn6MzpD0EjlgXq0f/O+V41bcYb
Q1+QSQjPmoL2kVdCm5anQH7LCeMJfFfMB7Tij8TJTCnT6BtjsKbZ9D2v7AAHpGGy
en7b7/YjKC27GBTsJzDHSUuLRDMKzttItFfsYy56b1kJJlTWvbEIeZv+IZ85v+Y2
ra0vrgvDdDAojKQq339IO67nQoEN5X4+YrRu3aV7Wg9fq1SZcHe65TIqJsi4b8ai
sBrPYmNAzTUpTd0oqqTzpay2GQnqdGuUv/9GqKkBTEmHcDJALrWyE8PUAZDkj90l
J6QZNshb47UuLBI9Vbil6MJOrwje4iZvi5eb9ALHDkKV2d1KedFQVqPIYS24kEwL
fMaDgCFgbSVZ1+ARQg/kiShVIOI6diuqpghMRKRCrAn19APB3E6deDnz3nErVHog
tErkvh0mkekBaSUNILd1ctoVrGg+lugJh1oVp3uJyVtyI6J4cznoDB9uZzxrkpW5
An77Ujaayreauduz9IwYn1qaa9BkI1LvKghAR7zwx+6JbzC91sPHO2sEcyvfSa4o
sde+gemwnRQr233Jyoz16R91XZFzE6tFFxS7HiYXwTiG24njvpcC3K91sLi7W4/I
6zx81vIwRLMg5z/xvHP6DI9Of0f6GSO2K5rRaQgM+Vhcdllf+k+sGYegB/Bw5Lyj
fKaj5qC5oF2H5+Te1qZLJ5cnv4CEgRJFqzaqYBUr1llLyYqWrNMxMdUgtkeMppcn
KxObhSL7k0klFy4BuAfgAlsOpkPN+U/Qn4WYvq/0m3Lx4aT/syNC0qhauJu52wjr
rsDNxWYH7fdsGefmjrZlDVgQHeaJ0+k29XKlbz2he5YfrBwLEsiI3Xh0gu3Ul4Q7
vRooWE0ldEQBkW40UDOThW/UvbDqDT7JIpzZoXmkOe3W5xZKoGfxZFoXtJ4c68G+
EMBVkIomNV0THIjkT1cSAlRs7rVehUgB/91NFFgPcSXEAjgHJoQWVClX23FR7x6N
Ehn1mzfLpJ92VyDdk7bnRjgZ9lq0j9tGdtniug/WThF7LF5CEReSVesSnsUc/BOy
d/7FXgRj1mI0/Qriq/iCR1wJHQ0tZHZUBYfr/oT+2X0aTEZllQtAdAAL+Jr0xNG3
c0YzMB9s97WHfTaYq2xdInxLFedqEulNoInvRM9WvPoNdu4YpSnhuZsOw5RLMwDU
GmTUsAeT/6czMVVJFxZaheO0ogJPlcck8c1Wj7iwv5w80Wvs31KK3rH2BG+sdrDl
so7itGez/i09dWvLSAimGm7empA/4FLaeKFetH9zM/3XMn1LgBdbNLw3VboSnCV9
BPhemVz4/m61+KsnibGZ2gDUedBkkhwJHXrX/VqOZ5jNqOU9cjVybdy9dJzYn7jL
cACqG7Y6DISQuWSgn0QSkG1WGWBc5w2Ul/oy2SW6ZsANsxZm2eKCWs41k0nF0O3U
b8irQCrpKUtibHDyPWbS4tUtFHggWLdhg0SoLkfPCwwXhWDeQOXKnN/QGaAYOkoP
Z8T3vq1BjARJwzQJKq6Qtfny34Hr54e20SZoOrBzgFaZH5ObWGQKoSbFoL9tzFTu
qka6b2JJuN/b0l8JJSBXjERsGhA71+WgVRP+CHYhxwDYEH+qw+MnXC0/Z8679uKK
jik//F3eFsqkmDkJJPhWQuwSsbf31wXWX/MFHYQAo+zHLUob+zJXSd+q1MGWbktb
SbGO34tNMkkK9Fb8msM87RwresSulIFZZ68oVyZQfu1ljmFm15n7wsWHKDAcpnq6
J18cd43HNm3+b+PyjnUgj1y0P5ma5WUYvKhBSUXPOsJodiBlB0C85504GhdZGT37
H79NeDZqbKpeBHRxfgTY5mE13ANsveEz1qzU4ffbPM4pQTVaKUk4Pwo7P/sgQycu
dzzlhCZjYyVZckYJJMPAtEsOMSxVe7jzL8Ataw0gRNwlTATI3Dl53c83qHHreu5W
GERFYYOzkjE0+eKDsbxQ8hYNQ33V0Z8Ah9CV6vmUUbHDFc8U1Aoh1Y9GSkQVBTIj
Kvip+04EzfDC2Av/lVMsvpwYkwi+GLAc2CaisCeq3D7bAshKpzAKeL0X7bEIxlcU
ejAF/YbgY04sSsbCb7Vn7X/xzS1KISGPAtz0W2qUm9BfCg+Ksoox0equUrS49jS6
waEq7OutCB7ozJm1zL1Hey8+MdAy4AeNEA2LJGqu7IrXUbHJge+5xB9TESniboTo
8ZZEwnGFnLgUmtH+/WgccefA9NY3/ebIA4MDrw5lUt+EDQkFkT6Kjm/nin8euvJN
UC11iDiwqkADq5I+3xcX6bYggAXP3cGGcWe+wzO3+rHs/scCQCwMPSt5/Pa9mj/X
m3J4TW9pjKABNzomBEKl42jky8oMoIUOvrdKqOGCf4v06NpK4KyTGeqccccdUODb
vJmi3Mqt3PiuJflSgYacdsVRMzWOSQGg2sGc3sDTkxfAaMg7S//G4gvHmYza12ca
woDxpseO/p22gtVMXdyiqESl/w3E0GcjyW+wAwrefFISP+pLurXal59pOtZz76o5
m0PIOU+T8mE7kbTakkW+V2wMncdz808658uebabSMCq5hEcl6KaNhXOs+zD1FbmD
H84cOMW+n/+24EyiPFOAs//xyR7iVxt7q3Du1UerIW5bDPBI9nuu7zE6f8sNXyiU
c6ck0eWiK9ZRDl/YD7f02nRo1U86DxTm+3xBKdWqUBPw3iuWlCE+urW5w/ufxz+H
uSPHnirT/HsUSKMhXaaddBBTu25kLueB32GULaECLob5yp4CoiLMN+WxS0qe3alA
YI6tJoS7YzEoAmlYE/kqmx94iTr4NEGfqNEdWIZtZVqR7EYtHRPd6fxrndcfij+Q
FTi9jKK03rN+UcwU71gKx3ITHVbMO7GTIvvAoJnR3g7G59PX7pF0yp3IcGj00igw
b945Lp+KnEKlitALicoVABQIIsvOKWiA0yNtazIJKw6DTgCaII08rYohn438H9iN
eKL88pRO23Xk4BtSfvAbJ6c6/dS7FswQb9CYWpvzOjgUjgMS1dwfVx7suzteUVTa
E53BSa7fVhDEH1kHl/2rXmSMTEQl++W5bX0AiqdLFLnFaQu79VJGmQcNymsbBJx4
RKMN2TpATLsrQ1efcpbsFiwlCpFoZtrd+yKcbW62d5LT8VcRt5NLYBCQoBjTjByH
Ki+9FE5nUZ3ErfrJBoIJqujDo46YXqnUj8p/eA1k3sMm/679X6asqLXE0I7Gjp07
MvJ4QdM7Cm8YjpGdWZVhbGjbm43hDlt4fwzCN8tOMdF4djV7HYPrN2JelYZOfZfK
mzBLtbj093azHruNEYmpuz2hK2Hwzb02bqxZJgBeQ+Xj3/6E60w1Y7ckCOKl0P30
ZqaRntZcEPB++0Y/bNKIVC/vY99ne5A4jXVkvsyPFnP1kTEuozTyt9uJSAQyP4t0
v57uFaurOgxn0hyDT/lFpgqXjVLkIfMKDLMnU/D7NTfmw68y2+c0q4cHJxmFS5G5
dpm9Tm9rjg5G644Kj/Tx81sOHDCgbGoTtZkbQ49dTehOfoNDX0i72OYLDEwOinqI
bkzVA1a9GosD9xJzwoTfLAZp/DcsAGZO7kMjeRTTL3g2SdYFY24vd+rYZNlZWAHU
4MrQvGGcfje0+rqYaRhQCpoTK6RtRAGtDHVLIxQETJ5tRTTZArRFxKtYTOYoIgl/
n6PUdw4oc0+suS83eYrTTjioZZJO7bEtHIZtl8X235+S18LVC14tunf36+agu2mb
OUHLRb+pHRn1ZaQcsp36fG6HXCN/fD1/yEjzRpcG4rf9HTjILevGMkTUPnDXHL4x
5GRrxrw2b/OuLHkmMtJSO7SWJwTvP6W2tNWoevg6ccwXR73/FIqfwlfCK7WUlahZ
Do3XpNr7sg8jlHrS/b5wpIvTZseUwoi4E68SEIk8pdeZqsRNEETWWOzpkCAaWtb9
jMdl8gqkVu77AYCbtafJHBU3GtKO+wXMVO2J5i7jLp4AmAJOpJVOQ9gs3brWLc3n
p2+u6Q/2MKy7oc/ViG1MBSBxPUVBMsU30znQTiCn5V2GjzWYlsE7LF92NLgg1sFN
bwL30FbsctLe+ejaH4s9wVEZrZh3cR4xs7KofLZwsimj0WaeB07B0W/JObHdsdHC
qIzxRH1hHHfeUPB2Xbm/hO4J9uJq5MmPcIDXtrcrXEh0SFST7rOnPkNK/mxyNX8m
spqmMJN4ZWJwUQh0sQ81gTVSmOzufYCpQqX5ERJYdILlRtMokELE7VPQo5bw8AHC
CLWJveiA2EA3aEiwCo2T/TJUT7B/yUq2jm2yLzxLF1Qh7/234tD6WRSN+tq0ggOz
BwY6O3phq5AtWbj2Asmcqywnb/r/mihyqYoZQtz0FLahI3D2ZJvILRiGFu8nlGBr
uv0lZt16HaGrtfiXxOc13lmc6Ecz9w5xUrmmOj8ccIFUM5EEg7W6vvBFE7izdHZK
jb1p0oj1RVCNsJ9rGMP2Ga5ZfgPJst/fPGXKhrewab8i2e5Mdpf/or6QtXQ2t/Dh
swVGlXcOoW63yX5oWF+Yb/g+hUfZ8mMTx6dHUWpR/wQ64F0Xsf5VaB0ex1eVaI2k
9P7sVgFPdlEk0xhmetlJjxnmTqfToNN+HeqZpUm/CB/cjRyxpepwtRcVBIGBa4D5
N9VITa1/4pUhQ3E8ZBP5rnyLcWfROcaHVruWlWelgfl46MiUM5ScvnDrcrZHE6Nw
VVNOH9+Nk1bOYhHnLnBLPdteWrfTfUBXdeP5hz0b0aU7TEuzxXdYZtnM3h/tEqYE
tNixco6vJjXG/xyOeGHtgp3GJnuO+kfHfZnKkEJwIiJEbjvFkBnqoSBydzo84G3Y
5ngHG+yj2qUU/lqfB3O5eHcRJxZx2uw550ikwcSKrrSyBg8exXJTk+sC5OQRWxUX
q5ClTyswYhYRM1ng/biOxvZkicvZqlEZksUfGsU51nMF4qLWJfWz0jV0D/Uv1MMY
hajFcFKTKCJtLjKWIW8Kk9+UxybBtVF3SzM0zX5LoI4K8Zoe/MeTvt28ABloVkyX
NIpR7EAK831qWl3KSaiIntHaR9xP9JAs30BnbUS16GHDfC3W8DvYI59l1I3yHP5m
eubqG8/ayBtGkR+HkcoDeR8hqt5KynKglSWnofLYJSXISN2+dVeXXix8TDx2Sumg
oo/1k9Jgb+gUVYUv6yEj9XrCQ4Zm3MZ6i0N7zlCN0DGrTvl/ODZYndE52jOBQ/49
HVQyadCztN4FW2SWmGPad0x6CleTD1mL5m208vsymxfP+T+dwNbiEOe6ejK/4Nak
lEz3PJosLjEdV2gMFKoKe/J808z7GgpQzUWcOAID5TM8kPrhwaik1N2RbWdJftTJ
SgGYJ4P4d6DE5ahQ80+SqaH7eliC9XHcdQSJTqD8CQCH+Isk7T8DnT75mcmlfqQW
jkt3SIOcj9URYWUutdBf+SOkhP50EJZYMBEnB5bMeEFioLlrKjBDWeVnpJfOkCG2
9JKIkoN0QaNCch+IA0YuToGFNNe1knmhn0wz3TxV2yyu4lB4AzUWZG0wreOok3vT
4bOoztV+gUD0i+X3OTiWJQGyyQpA7/kCdFelsd4zvR7oVx+04nrWjzB4XJJ2D3GU
/3Wn7rgGZhOgbAKSWhZNeN8zleSW439tBQVH0DeZOziY7cbSyrnAdkMPIFMZ23x0
lKf7RUxFibb8L7dL4sZhBsURcpNXOfcS7+bp/wPNmbOWjwsEybXrrsHEzoI1Vtc0
unNFfoCv9k/D0RKRIbHq1BZfmLxmKojW4y25rQAV0UbN7YAypXAyewsmKXxAqkkq
XzgfIt7+q6VWTwHBDRc5KP5lDdNoVc2oU0NnPYPkb/W22GG8z+m7Aft2Ajx5CQ3/
7KbGOepbadqsC3bHkSW+K5c0kVy0PupYRMr8wf40jCQc86TtDRexkX16NlDt7ejX
oJ1CsS+tKDpUnIKV+Vq1Zq2eB5bFiBskfeCjLreMBSpeQ08HBWjE8ieVT7Oi5Jdm
PSrXopEo+D406g5or0r5kLIZ2gDfs3YfVYoEFm643qOVJz2BuJqtIiuoSjQYeewE
pgcaaFj1Xh38CsiWK99U0RYb/96bRib6GIdCPFcL8CiiDHoszlksVCWG45vusGon
JalfwjjR99OnqtCC90vY2611/iaBypQkEjtmzGpwFmQPVif05QWqiKaHL+Ftcbz5
wSw1DYszjC/OUnziE38Yu/blT3NN8nxPKPqNGKz1HuD1r9uxbkRCDHpkVlYMt0MQ
2yuTYG+pRW/DqNbPp5wJkvT6TpIdDQUj3LKP1FF4moliUlKhLHz8LDqnmQpB1ZRZ
YE0Y1dOLqUXkxYhzNqVviCgsc6We0BQwHrD9vnvOrRun3w9NCaIwrS6uHYzG6T6c
NShNpaKN47mn7mnLp4BVzEottRILNLzPArR0TAax/1oG8ptfn27KjtDJNM4OTqvR
TUh6H/PUVujeWXds+rFGaw+hN+7xB228K6vPtLYmKxGNXCRZ5/9L++9M2AD2eaMG
duGjZ+CuSe7lvM0Kk7tBCpu28mIGyOHrB2vfFEljH8twz5RAgMbAWPLIhf4zgmHU
1HV1Q6PuLkei28pTcLg/7wWk2QOft1BBKqh1rAfp4qyMzNPDlRYJXAIvCG0WO3bG
ZaYh9xSDJyA499gJFgLR1iwI6nKEbxeaqkxm18kQpSDTQeUtziFDfTtirrANzvRS
aMVNYAF8YvoC1myvb9TtDT7M381nur1Htzt+yZspj3+DOakq51Wsd2wo/18rPRXy
xzLd62gBcR+bVIy2eb2ndjUN6rSwckhtGxEJKWp6omVqiTW5g77gL13dpH1cZPe5
YH3lTDmP2nANc+VevstVqStnO0exvWOppOEr04Pn9eKIvgyUoThmBj0iLMgoHk/3
84o5l9D3Jg68a9BiJEG9fepYlmiM4rV39k+SIulrs1uUbZxIyES4rkpB1c+Q1NDD
GY97kuG13fkXqeaAiJuQaZ1hSa8+Yj7uMTXrqzJ1H7aljriYWf2MK02iBG811OKq
lmvHskHcK2D5heAlIx9zH08ebBvAdwV57yFcR0Gza0rTT7076xbOvYxSP/YEmqkn
OO1ts3UOHjrQYcPVQ0TFcHYkMWfEP2kIe7dy7gA1IF3ZlUqGOHUzRkfYJ8I4vNeZ
2mgT1qLP6/i4Gy2CinIThtb+OeXD7jx//9NUiG6cNfohAc92km+27MqtFg+HdNvP
hEa7XiFTFcWnH4HeojXyH86WLNgYbbASlH+8feoS+aJEtuTlgWymJB+MB+azxWMe
zPg33l03aWOXLBa4i/FJI1KD3EQ6i44C6MdFH4LschwbZUXJYLDgpkHoKgGFJH2q
LvZyiwjGR6wW3QKPuTfSa1gVcpuZi00eq5o7JhMSR1IhVzScAFd6IzOx+u607QSk
ETq9aLKFd8Bq+bDwNSnb7qJtkDGKjhV0m70BlmuRIaKMuaOh5BhLfHUND8NQclzQ
QhRLneJa2ru8XHiaUjtLCpkYEXpY1VAfpBsUeGdZrFqWapePoutbTGcQqpriqbDa
b94F2890pVAcFbuzQalDv0SCPW5QvotYT9y66WmZMXXkt4alIGJB9l4wwuFkrakE
ro6za4T1fNpDUcSRpQBkKqV1U4riHk0caDGblSi8p7dEHSrcCBOG5zWPechg7ASf
9NWb3DEGXwvlNK87x2MHm/R7ZnWI7sk0ni+EamozXDhHScFkbm2Jyps2KvRmTkbJ
ouynIZKc45dE9LHlmCnC/wZgusKNQ0gVVEnqX/KgWcDWCF64e4d4UsLcRkWzTsjV
zPaU1u3mD5U+kINgPAf8kQna5jCQdFhDtIQb2V+RUN9q3PkCCHZ0xZn6QEhuI/2V
173ugxR/htZnNMlwNlgbv1vilgKYADQoyQ5Rko5xu/tvx+JKBJ8T+KAfHvWcQCyd
l5aj+pLEvQuE8XiNG4+1vsP94GnJfcmIjTnSOIaF1PiNSj/vPG+9b3zpXijWFAqf
adkSRRXhcrOEorX9leWVItL2g6oabgwtT3W9BE2A1t6mMHnXrfqaIiZf0adSe6h7
spgE/nolmEXa35OOG4mDqD7FSsley3m/spg6/vAg02VL53F/+9wdpD/z8S0sd7fp
xf4mPoaE0giOStFBENzGYx2hEEhIKE+UpUivl5Hxo5rtBB3TciivtZ4MUmcoPdRU
/4dZi7AzLlUF9dulfY37UayboxCtvsihqS0pCMMpEI0SowUFrcdT8F61WMto6GqK
SCmjoevj+VNdPSKyF+Y6Rdspl+3MjQWBuQCHVcg6UxhVyK2F6YW2MbI8qQmF+kE6
ILHtabGcHFgIKtNZgf5dVu7k+9p8BdiAEcX40F/9yj4eCJ0n+Q42+H88l6lCO/EM
rwKeRsNBzGwLAnVohBORxajvTrSoJCjfsYLVbQr1v+Mm0xAC0GVSc7yx9rLbp/lx
bmT7qmdgDHuPLvmPVzMSGFgJ27H5FadJuAHaj/dylBK7lJzpbOlyssUbblTY8KoI
p2KwfUZxLUvFsvS6MehNA0l8XXRUotj00cy6ow4a+T50THF7YGbIfyW2MNVgNI+1
cQJKOqemIOILn15TEggPmr/2e2DUMrD6Un/CwPoEY89FQ+6kzhdfvAk/S8GAIChm
fpRdi3Y2V7VZEZpOg9imro0fig5koKhMCwASJkAufcZEgPMhOvuZmszZ1Gwu7RI7
rAua/oenRQYFGVNqHGkkGgfE7D4JA8zxovACZ4nHPAM7V3K5l6+FD2zhpJ2biPZF
g0LaiN631+by4L4y+iY13xxjwyuTdO54PKJs3FmkZeRHWQtdS0vQhQ61yg+v2Z/9
GPCDpKTBF8MVHTX7SZUwl4i8Q8DggZ9PZOdUwtrY1IIphR2qmzx0uMD0t4Bu1J6y
ahVosyscwV02loLkwoyy+mUdObq5BWjLRNU6BF4PSvDr9nrtlX4RCyj/VtMRH784
zBPmPPJ3GvPnFdSM5Evku7HYDl+n0Muj+FWHni6VV50fUCwYaqr+mkKXzKiKxfFF
wu1mnAUWqDLr50+Qv2fGAFpw0ZFxvELuyoz4EvkH+RZXHjSPxaOoBNjheA8MimTz
PXODTTRQEOoRFGWUpFK3B4VfB6tCFj3lZnHUv7qfRz15cuVXb2x/LRKeIbGtLsc+
qZnBDu0altdY6Cv9MMl+zxtv+W2uMvnHl9t7FBEIw8kNLJe+Km3YXf0RsCn9+8i6
5c/EeYizYFwtjMwS78m3kDaWjODp48g/pwUmga1NZmrqX78/09HQal8cdNhsSLwB
ymeEmTdY0I6jwFeNYrFo2MzM+/yq6qEIroAJCf70F0vVJNHtnnNBSRZhuLWBG01a
jnNulJ1vzMdwntCGOyrQCHel9ryV1WIAk3KIrk2QUlOZQQX2O3ch6XIJ4jdGUSHu
nM24TVwZMeJFqEWYMiYgRU8XYUL9ROBCLc6AuMDKIdLhbN2TpI/5yW6Rs5O94YFZ
WaaPKDnTYztwh55MLPieoYmr9AOTcvjEeKsKivArrudpRzYp/XbMT0JlmgblY1go
YWFEdmsq10msja6JsBqPkW0yflrratYWolSmTfPlYwwgHoYuj4wUZ8LcqalDhTYj
ch/FcVjbZ/BScfU528+rx1Qs/XZN6zKcG/32V1C1FY/IszlqMSCfYRDOROVzVrZ3
L1PEiS28N5Cs7mxxGdN9+9TAfvSWdOrRG3GGHd6gOdllYneUuQkGQ4uiIZkeL9tL
1a3ZoCALrIlV274XoDTbBfBnh8ghs0WbayqXamn2MA1yydCoT+2YtVUKNs6FUy9D
TLX7mIo79iArPRxuIWCKIKbgErr1FUlrfMYlmxanYREAG3m9ZVyVLqddRrFhQvbv
fQekpSDAiuPHycx76scn0CcGlpF1Ur9XvhAWYcai+Zrhw89PVcCT+ogEbw5C6L0K
ljMFHSILMhJVWCnch9QL84wz8H+7di0H9v6H3pNG9cJqKlEnxZWChfo8diiH3IbQ
XdIC4p/Fr+u51IgNJEYQ40n3La8aKodBoMCT5Jex4FfZgHDzZql/4ZpPY1yucR/q
e1BT8ndVWEQgCw5E8HZKqGf+7FCH21fN6rwSZZtBqd4mM71fUhrfWMi2cr0Za7Cj
3W1f1LWZf9VuizQH+k+kfw2VIKcsBeLrNpYpn/MFMuolWlwH0KMj3xjeYcnItLra
gitKYOj+GjqHeCPPAoSvJz6PmnNfUjdbM8INbenQjd5ma/RDDuUy6uoAzIf/XBKC
oSezXORay1f+TJ5ubH0jlrPKdyuA8xWXyevsTtcjy2l6DUnzi/XnQIpzcotOQAki
uL43EViGahU592DJ/uQ+STyXtGoduL+uChhr9hV9N5e4Dsva2Nju2xaOucCMXkcH
fN1xvLqt7i7RySLDdBr5nng41afh7SgDr4ruY9VXdo3QofCMyrzXivSq0z7hp+ql
5dint7YMekrBuvPO9vrm9qtv26ZNhXy7SlqVk7ensKGHGAxfzen9x8cvgvAYNRsQ
JWB4HhdfZnL4HtNGf1nTMrhxUk2bF0pvcTiymDxF0pyz7eYpRFXUTyPCi8tHmL4w
yf4x0qWulFrh9i/WA4S5je1rl0HyMOYHszXFB5QtIsHa/ovZp6Q+P6YK+/kriKYF
`protect end_protected
