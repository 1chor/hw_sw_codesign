-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
hQSOMHN/yGDI5yMPkpV1PCYIOOeoyZL3dZc0BccgBK9/WIpqmNNy8LDEA9lkIA5F
GYt4XeuAGXI/vyv5z2mJwzxTS1i30h/qUCbgoev5VtC/cfkrW3djX768bP+MI6Z+
o2OntN9mdRTk+5lU8G5e/ou4mb/iGq6wJk7cfXH56gg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12496)
`protect data_block
EWOFX6gJfH6Y9EGWXO7kB9R8bJlN5aWnLTFu6Q7fRCAXIXazVJTK1QimB3wrzgkh
L0zZn8z0RRJvUu9j3g4IUkeTnO9ikFSLTODrRRJBdaB5YZstLAo9/R1nVbyy9qMt
QY3eCt88xW3Ny6CiQXrxcgtv0VTDP6HEXFHV5/aNfQR29h8qHtzUIJtDSTC5aBVt
HPN+SeZ+j4qp/chS9uPrp/13tJmW1noxnbCzItE3LBss8tpLDhjGQJpfmiVwscWg
ZtYgXnzWOK+KfxIC3bJEgjwgTHKlM5FAR9mYJXD23cpenGN7rghPEw4dILPu5GTY
KV4cgZgTXGJikTd6M5Xn0RIkHhpewCQkAMYflfUuxdhcvC4texC4tdIzlRb1J2jN
EEriNTxRIPQkZy/DW+xE7wS7NowCiG4A21aN4I6Snv9Os735fJR49BoEbSr42s10
vM2FftnDPESby/82zknYw2Ub94hPHNl3iTwLWzd1l7CZUEmB0t4ispl+VPsZXGPX
CffsEPVNa7/AbekqxG8/qVhSvjWXjBR8JdyPLxhAKy6nRIPtzE9OsqTy/cRVn48x
v5WEp/36Ni68uMg3tIhS23e0hnntMWMufauKMjsN5++4An7rlxetw+3xWqm/8dhm
wQLazsYAH1X4B7/5njKsNhTaER41Z6XF1yikVtaexZ02yLlPRsyJ/3JnLkGt/bCb
osRAwswxDYefD5zf5d6Wqt/t863M6nBj+GExa2zPlP2zrtZP6NTP9K7fSOSH6WRT
sxsrj7tCP5JDj5Wp9XB1772flAoLr2CkPqiqUEGD+mtmaPH/BNVqSUkppY4BWt2J
UIr7/FNmdiiZZxggQYEeekSllkPbKLeiyV/i5h2oSSkxVNVpPIQwFCqdzI3da2rT
UOQa4nXEwqToP8CJ/Pwx5H98T6pJTs9tpjLTCB59SXt2VfIbo3kxsdL3+xnJjSfQ
ayrJ9r3aApCXXwS1V61OaxaWCP3uOJkidjse1p0xOTNBgorRGo6zqNS0xkQuYDUO
ozh/E4H6UoMr+R55dIrInTQbvpTF1SofvyS7y9QYzXKv2N+OE2YUgg/DGgjY1C+v
b29nui18sPhZP4EpLsw1eKxJ/bIV2UB6JacqySLoYO3zF2KGtERT1iuVdIKT2AlS
P8HeXyYHQ1NyxwqgKFvUV3G3D8UBgPgtHGJiBZn2L4EGqaqhaIR5gy/pghx9E4sv
E+QsUsmGHNF4RjxFuIH+JjPqiCavd6Pcm0vNkAKTZhBsOMc2E7jgIWAu/lbrxTl9
6J/3Xpb+cQjce+hxYzaDzcWmHo8Xsf7I3GtwiXZe2T2OP5d2AfPEd+2TVI6h9mSI
T0fkuYFkOzEGifXFyMMKtL4ht0duMnU+ee/GZR7mIH0Nfbrod6N4Y5CuNN2HTEUN
5rVUMAWId3AgmbMLx4+N/ryfb0xWgRIc+tov2GAB40siq/2kekJkNDtRB1lp6+iz
G39PZv+O+PeE3ljYFe/yI6Z9c+n3Z4Pm5ViZUmxp9N8miYc2Cz/POPRc7g25wHnz
rionnGNaVlrjqlfr450GbVVFDPHaV5G9laijXgCWm9cGJUO3FJ4YwfBELSHyc4Nd
PNUtRjpynt2U9iL4jGUjwBTLn9G/n3NWU6htICi+tWYJCo1TBqCAcRSAloYXfE3k
CLE+eOHgfFqFvp6rx3LDOZcSOBjlkE8M5XrRZHrQFlKcFvpbml8tF1AhreriC8HJ
d4aksw0gBCngoHf6htx16dluti1fzSR++roiv77f5e5/T9wPR9eW9GssRkDDdZKG
DiKgbIgs/mireU02NKKU7cj9X4aJ3LZJuOnM1bjE5IWMhH4VGA7mszEkIuuJlc7i
0D2N7MpnqooHvCY6ft9P7paG3GkNDYrGS120ctKRLdl0okvLpsqIE6zA4kV3u3Io
D1+SC44WoIKFZ0az6rjL+fbkFNom70mgm8ACGU7YXTZoDqVG4sd33z5fACP/Dmr9
Gek+4dhmigPUieKqDDlsjUbpphyHuXkX5El/qZvkGqG2VmrkJYSTEw1+Ha3kUBD9
2QHlc/24OWa07Pqw4VAyZNjcpcK1NenZAQPMSrbMed93sRnhHpcuxv1MA0/+82HH
fCEN+aalSFz8KxrCgRrpMO8reJ0igsW9urN00tkAd3nypiYdP3balq48hYzTLK5/
QevNjCRtGlUo7hsZyAu5svmtJDq2mkdBLrizC0TRbY5wa4hUR0WHlIY/spcyE0GT
HYzG5k0wkhCU3c5fYw7GvgXF27TV+yEk6Q97EGfaY22DHdNiFrzuvhPjvHEppFpM
eaxOCyu8Zg05RJYhypTZVdZjVrbVz5zI0enjZlNw5//xMRcGDckg0NqCFL5obucG
7XFnlRsGnsmp1A9TnQDH7d5I2dNBxqbPKYvcmaHcA338OljtxYwSALl3z4d/wRqu
6yjbpymtv1rnztH+gvKMPMaPIqvdk9iUJl9uhLIviRzEwQ6/p75TxGy2fcpgieF9
MGrneoHsESatEhD4kk1bBgFaEXtQzFwMMrc3Wiaf+aB0CEHXIgrnosu0WNIE7Bni
xLyk7UL52xoRn98u0plIxIrYQ6pLURViFydtfevI7bzJMR9J447fCavK04E8mA3N
sF4ds8U595p6J25gaXGTHzfuh7ehBF4enSbFAHQ4BkwJMAhewh4l3iyrtbUBapON
E37AgQUH49wTJd1DgtlDwXNcLdeZTMd27tU3pYeMbyGSRhnZNfSzFk+OWzXC2LuP
3GEHnaE4AIyJSjlHjXzLufGVgNIH0NW+hV3QIU879wAAeRcNB2E4/1mQ8zx1UTLB
QP21VZ6n0GmzYdjr3nedtCdSRD+qKCjGaZNjM3ozoTlntqReb4fOtEy489Ot0Wr0
P3EcYC/MOTtx9BM6uPoc1uaRLhrnCJK8ihZdlf2Mmukko5tGDE4b9YJL2jB6lVdO
oP7r2eOSq1ChqxMS78aHc/c3XI7ciXJG76kcc6z2Nr4aMIWrYBUDB22mOjvAPbQm
e6v3YOoA2I+LfiIrBw2uoFUcHCZS+hI8DLRxTmg52ZHs83pomOP+0EiP9474dCrS
2Te/4lg3REE1x2Y3Uq/DMtOakiPZA/E1TeetmNb8tq+SxevCEFNq0j3GEy9Of+ms
SiX6+xwhI7fPynlMKeSkvo1nIrYOWBfrUbzQO8neBt1R9Au9yS4aSkzgXNXlRVqs
pzUKQ75NnmFHJZvSwvirV/p533C2KrWadO0WfFraizr5sLvNQHrCMPnpgwSo3C1C
EwzqMNOTnOWrW2tJO/J4Hnr7grwOzFuYL2qW8ifzOwLO8XqXCihjaEvRZYFr4taD
9TPwNq0HMQNnvTwmZ+NZwXI00TJljReBhq+wkRpA8oHruWXHMjHmETcfyCvMcXKZ
TySVbkkW0Cc9CXoWs+yydqugIk4virTvIc4VgsSuI5EWlnlnoW4mC0YJJyjsz0sP
tT3bxQs+hFEbD5YfyWJeyD1pI++tzbAGgf38vZlUZVHDC53PmdbajGXc0/dxDcl+
GneFo/E28ECowDn5XJLYfbreROM5YEUW5mSheE/mtonNHVBMFTqOBR2iFY8/Xkmn
i2M7EoNp6YnLzowUyyypIH8mW0h9EroDoq+i+K/d11Oi8hB8Rj7vh6Spaf8ps8hO
4KbrUDNKnrtRp92Oa8utmiASxxfRE0QhsTFPsqwyT7Uqy9K4RW5QGdsreYT75H2Z
4yZhJAdCb12mfS2QREYIKjvKuqhtZsSLFXHiyetWAWBvNifJOeUCnAoKehBVN7k6
FfvqnOdpTqWMOSkPLtyCOYA2EyNwb8ec63ZAYdBubToH0rpdc3sQzzFHSWS3qTlu
gHwJ6MXp6Mc7UK8crXU2adB9UGxTqTu7SYltPjJEJmZ5XquxZ6aeAZzYBSCguKHR
7huUQY/AtPGibMuk7mq+a/vjJeu3YIpLRqcbsxmjpOaylRQrhEWXuCGN3bKDe6FN
ycV+MBVSHqe+NWryZppGayGHSPFNphLPMHQCs+T+eC0pyBettKX+dqBLfQDwLz89
Pr7A4OY1YZX99d1zm97Z9JFiuo5XvEiYeKuE2P/C3sCQoZjXzO3eYSU3vp0d5tIz
l0564OM2BqTkSZtMst7gFZdjna+Pm+K/HeitWDZv6i2EckI9mOszrioG9UNtnVX5
YMwRnAggTAOvUUHgKCypZ30yjgnlUGY9vUXoQ2iYSviuBxiQm2tD1XvncIiiQEvV
Ta6WPSr1so6421xXOM16kc9FYT8sOLut9SLzIyKAJFwMzFxzzMIP7sIlIrQVmb+/
4Cwu47hElmtX0li4KU+ALC8q0YUjnA2NQqCmDpsCwt1p15fnUGBSG0qUjd03obM8
E5dLefBr/3hln3MwrAOTgcEQlO6Ljko43gWy92PJQ32tu3D/Yv1FT3HQOLWUgcCj
FBHCyB/uNarKEVgQz0MFA2GLoQZW7jjCo0yhmpn4+jeafmc+xEa1AuafFGvYpZQy
8kBkX3T5ctnmNTMrfIosQgybysbIuyybNjsLNRNhTv+G8qsbcNkVI0tQ+wzknfMn
W3lhNXz6HqWZMntKbC5PKzxQLU9MGcOcaVUf/OacK0YzQALthjCKlBIXhass3z8b
IhqNo/MFVs2lBWzQrMOUlrD+UntthfipmdF01OSs+5hMVIgtvLcvkvM4JYiGHxxo
SCFDrXMaCbd+5OoOpUwwz9xiphwCeeW1dpNT3bexwnmpCMNHwzDgJLsK8yuH0zx0
t2hAyraEEZ8RnxGXTRRLVmdgTfI/6ZgY8cQPSwsQXJI9sU5SRKs9g1HHcL/S4WH8
sGKqEbsq+k4dtl3FDY70iteg8hDQVGWsU3rPeW++nkwWaLkXBzr5n5axxfMdmW9l
IkTtZRTiZ/CSFvk36WS6rgPdghpocI5BoJxoMwglX/lr6UIdS4rhdwpMOBnePlOT
u/n3FQGVNCEAvxZ7p9R3FHxbDMSUzns//mhWpvQVC71QSzzV8pYBTY3zpU3j9U7h
IhulSj2WiGUTpwB64Pm2QVaAVdsVL+XkdMUDVP4c57t4sfrr+JvtmHp0abuPe0Iq
kurICABmRUwauyKBNeYqITINUt8mvZEPdydSc2yOJEUKbuUhVNHRV1IX8MjbETkP
Dn8N6NKTPrar8ZurntWq/199C/lUN4hcflSylmMWFnt6OSZQAm1oBHmp41az2i1H
XGXpk5JpsA96X7Nk9ofQWaLZmrYOz116Ais+vHnD2Gu4XleEGatAteUVMpH86z1j
eaHzCHPXAsx7YHY196J/+QhZiLmZqWJc3KsOexGlA799IGkoubis9rqXdfaxU/6b
Im40FF9gIakHb58ryv0wqq97YdKTzy8VdSRm1dgatD9/5Ab/uLyHIt2gbchkI+7f
wltbBHaidNiwl5ZZO+3SlBUmn1dGgmbIBUShX/U57PZLcEFSDUL8XgPhouLFt07v
wMCGsnZ5KkAZZasWiN9Eu2SsSLNJUrepkn+/mkvm/Rop1NwnkuNbFdAZGO9DkVsK
Q1+I8ZtfAMx2CVrSNeUp6QVThbbwgSl8xkBZQTrhcgAjoyPWjMFmhFLP4RdzqHQD
Yl/w+Kza/gLLdug15uIq+w6agHWTiagzgYkbUN+aEwW4BaM1YtGVTgjH4MC/JByq
M1mz0CZLlpqDvM/B2NFlUI2LcNOkRbXQEpIdAmw7jxjREl0b6aLnDbHBMQD7hb/I
DKAsMxd+GT4uEa1y3WGkPs4jIGQ8gse1JNa74cCvwVtSu3M5Febzaz45tHnkzvZc
aX2uaJTr7BZlXZ7nxFdbDrwEDOkAqceYlINyBpWPdZcS0CvPmBYlpi7dCx/qsM/U
IUfH+msvk8XeXxYGddyk+mVSYeoxWvmTy2ZXGsYqR172VislyoopAPvU9P3LIdtK
004Z84NC5CYKXtkSnICdF170TAIVbTKiD3URe8+694G/lkZPYv0dDiABAzL1cMe3
uxJQ2LqbIruspSQ/IhEH1bMgeYHnJf0jBQGfchOVWESbaf/ONNAqWQpMN+197pxE
njm9zLUmVMzT/H4kHmEG7smzq4cCkjjej629udngfFgsZ4fXiZUW2tKjInJgjYe3
l+ByRqq0sjox8AlBPSXDcitLqpcO3mdLP60JQWu0uoUWNy6+JKqd6jgTOa0L7Geb
+iVDaUSAi4iCnBlQey9W0YURrcG7P1aS9iBxKhsqjem4igx2TAMigpPrwH+itnL2
/IX/Px3O1LS1qxBiJdbKcXN7MXyPjuRgyvyhQ25mQHEDGb1atmABvgfjVB49Qspp
6FKSu7fONsx1cgYhgAMVNb193X1O3Npni9Qfzqbz3yW1uAeiVNpXe9thUU7as37K
ER3Itxrv07pSCcJfln5jILz3Etqi0AzL7vRzhvhmUFuPgNs1CbHyzc6V892CrDu1
eY1PpYZlsyS66yQiaVzD2r91IvjJCgzED+8iT5rkf5iM7gBnjL/AVP3W08/aEmq2
tc2/1AmWcXsH66zBksaPvRRWv9EhsCKPSv+Nnu/ZeDWB4d58KdYz+nB7NkiNM5Q+
27litC1XY53MP7x/s3jPcvQGtV9Xdih+K2w15pjZcgU2YfC8BCzI0fBq4sP/cXYQ
+bzxD76BJNKGA1HIBTsLti9/zU414EC1SLLsNglrqCcVC4yM/DVQVTOanzCSXtyF
9a1bhkc/cMpW/9fay9OEW6HTe3C9ogt4yo49ZGo0xFIy9zg7F1NZBwg57O2swMud
qKvxNOxt8IUmAFpUvRiHRXlxrG7j0XwGBI09THlpuF4uJuaEbHngq6DfgslZDCcm
iDli8uDHtgtE7rXOogLyCbqjh4aCN6uZVIWuPA+ziIZCd1UcS4hCnFIrlJDrnviT
ZA0WrvmANLxRcJzqoMKmFNB0jOF6oSk5mUwkh6fh+nOa5FpAalfWjmWNlwSjGP7f
iFLsAGFMbKENvVqZUbwb9QSItEkfDfb83tJgoDvikk3o/Wppt+JIAUd3APCt8Kog
XXWN0LafGvd0uH9XzNQdY6H3KYDibtE5EcyoG7NvH5Krt7LFLti9J6LjR058NpwG
74wXuoG47Z3gZtIC25z8tWdRdzQbqyt1yZV/a72m6WBIpRilmUvzlgqeUJsX2uXJ
YHzoalS03KzUI0UZKKpDynLIzqJphUPiia0Lu7AgfpGKiXBeRYq62NquK9oKYVl8
BkEl0RO/lrjcHMbIQahCaiZM0bVgko47ACbK2U4PvsYkvX8MLhtvvGU7g3T6WkRO
N8bv3NIuZMBemRUQr3sMu6r4WeoRp1qQtDJk0YLApIC7v5TDerktW6QddhF5KISq
1LS+HanBewSmb09p9EVooTephegyDKkj+V+OUJgnQr1MX4gLilkrwUimMt32BBmT
JgAeUP98SSfXAhS2bLZ1Q5vV3Mpx17DvCixjhmEp36d/7PWnwtapCK6caar7J8a1
o4plHfdf992kOsWE/LNDzrQK/WEjWXQkdK1S8jB4knI5YxdShQI9MqHD34V2SE6F
PDC7qg3S9ifcuBOj08HFFWyeLtBAvzPUqg0B021+zweIq+QR2llJeu3bwExWPDfT
9tX6Vs6RdIXVGqgtR3CoMmSfWKXr4hRp3DEmzXzfPppw7WVvUs8eA0jsOoBXLmCz
bbf98+rkyXI5L9yCBkiJlnn9HM7VvoZ5seMTXIEPrLZrxhZ+gFQSsvhQJlIXFjcb
bxZuPfvVyhniTqrNqQLSRGzo59sy6FV2533OuawKpd+qSx+JfXrv8dLKDFyXVY5b
TA3Bks3inzw7aPvjWmrPirxl6xv2RrBCtB3O3c6+hXxbl+OE8MGg1VUYGlI/EZhD
clYCesCxrtwEr/zymLgAstKfCFvKClQFe8bLDeN8UYpt9UNMO3CM2U0hKxfZ5BbU
/TOfm4rJCD/fYxfsUCMCd+nlL1IIWALNLVw2k/emDu9kFsdoOb3y1voofgnQ8DSg
n3gwF7hgo+tciX1swEvR0sd8cAps53GaQmI62rvYj6mYQU0d9juePqHE2+vtMKzS
ffhp/IvsKRXjz5iZE4nIc3tTqtfCOsmvnLeMNk/zElZ5h/lxK857FAoQVjrxkENk
a7k7B5b81Uy0w/z6Dga55MSaPnPin+7ydUI/4PdLmLcKffxyH9fyaZ6fl+ACGAn6
UmQPbH7gFO+xnHgCHt5h5uVYemJpfNUX3WdkoGFvnCti1T1ZmVe4PAsKfEvRy6+j
+2AtV/qca5tzbmrCWe6OjT4yYQ0/toi2pumq6g/A0MnHIEMFq2Ctq/maNJtcMwg3
mS3TZdvVftlYLiixxnwJ9hjoNnXVMctNk61Tiua/+U4KjdjUwcaJJCA+InmXqjUB
NXkshecP1fmI00RyuaY1Iryj4ruRGywu9LEG0wqlY3wS2EgktcVmE3KitAYB7eLu
mcgpVXD6ui7T6qvUU3fznKe3AMwVJKE7EYu5paoxm7vVMHLOKJZD1I2+lfsFG43I
6L63oqRRGAvlPCOZkan/FdI3K2ZlbrhSKJqTFMtLN22mSESVMwQrMoik5VNG6cdC
aMPvK+ZH48ssBBYt9TEOnAn+Vjg3vv379GJNmbduafoX9/DvoF/0luG6WeQa9lSb
fD5DMqOO3EtzeXG9VjpsxaK1S99DWm5XHIcV3qJDPI4zHnVyWwBXBl82EuUGqoLF
F12n+T6HnOTEz1HC6sBrukbjWWsG3oL6z7pHqcbSE0G3UVjoTSuj+CZJJF6SAhC1
HeGMR1Kr/npR4hpWcQgidQoXU1R5tXHIPrgEGwk+7WRU5e9isIdGHiNyiYfLSbTq
/6NMGbbd4QRNx56jIT9P3fsSbAChW+NIGPJT8Hf+ZO12p4t9e8e2bOSyJqU2s+k4
9vUf+PZyAX+R6dp2fumBwLJX/MxjZY3aIQbkkysljnt4lmQWwID1YyweElwbUNUo
xfVDmu99G+C+aoCzKr+/AlvkQaymXQgDOl0j5eGOy8dOUPX6xDLa5WZ28oKTDjSr
wMhn2JSazLcBUwO76ss1ICl49HVoRVsd3xYLllYhHvaBgw+I9DsHK53h6ibwhsLU
EARLMh2sr1CK8YrxZtvE4USugU63blbdnq1OYMnKTWepM26xLuui69rlc5sqSNZf
k2H3Ph8K8FLMJiHVG+H9XadfXR2rF0FodPncfMP7AvyOYNehNOalX/Xge2le/7Vz
SWfYkmduSaw7eOO3PUTowbfrYURe0vreyZCPT0Ly3NydBRYGBhP6eY5VZEH3ZE4n
0vczaP7OdeEcV6EZi+OqbTRw753yb40iAmxzYkvX0VvvyDP0CpZhmq96H/5vSOOQ
olQFFoHTERHvqLCZlOOeRVmKiPTJ8Cdv2fVnBQ9wmRfU4WWc6EpuLgRWuLZ7/vRY
/nS8cxl0Jka6vCYFSBg9tN+L0UVIRcC7QKbmt2Ap03iTMmygrSvYodo3wV42k34i
Tuw7SsclIHjRK30oQNZwAMvwEj4e+FIOXod8Sr+tXVuE0dhD1UTRwInKkUHuaGbk
05GRNoCTfjHXJqBAQw3PWLHWuRCdPgVTl7jPO+mzlO7QWEblNOSCcazUX75L1/3D
XPuDBk7ifpwqsLVilgWicu+JNOWdIc1UtsolCN0xeV2ohkRHedauYo2m+FR3mhAy
LckG0pS4plC46o4s+EMTOUoOU9YJDD3QV1IUBweBg4LD3zrvehS+Ff1h/tltu+PR
lqWYDpXIHDfH2DZWHxzuquZgvpI0QaG9dSO2Pkx45Gbw/oNyB6jUNo6qSj6Jk8wU
3c+bzK0twaVRQvt7L0m88kQQjZBTs2QNsmqw9Uc/bQxvsVGLCEgOfeltBF6juP3F
BX0lDgBD9qGyPhQDKZJvPAZdggfryRZNVX3a7eqtp3j8hMxCp8FzDORXvF7iRu/H
dymvF1gfwdKPsnGKkbXYxbcfDZsYZlV7lcCwWfjGUr0qxCspXVsix7A/afQo7OYe
ZAfMNJlQ+XWQHzuQTScNMX7dQRSWDtJplBycEc7sMDzUB90na77Lrjc8Jm0m54LX
whbZBFG+YwA38gUNzT64NUH4dyGAryNE+BsTNkdwPgYJA0Vz0Semrq6kvsVCZFJp
Y7daNtrvTGbLBz1EmWjag6E1JhaKoUiGmentvO68hIuZUkdxd4DXIGNz0R6p/8Uz
vV4wZCeEH7dLaIfcy0x5mMtovoscNxrm0FLeMTh276CC7Xgu9pUTqQKwMPbVCzz2
kYyLtboCkXsYklTFyfpHs2gkL2BEwwuaX3kM9Hb2v0OKPOKZL4gyY0Re137+rypW
gnUPOL/FnhghBTrxcMh5looNeZxzuCBaL4fK9yjcMWubOD9OI8oOlNLk+QDwouvj
3KFW3wEMyd0kX0QS2tE6gUKYi/Nr2dErhB9XaAg1rnaG96tdwadK/QN3bFbaOfFM
7+k07MnZ0QcOR6cJ3D2uZTnWVtCHGUOWxtpQHK5gcP1za8Cp2IazP3F40l+e61p5
5Kd2bn07qsLCs4A07V+K3Ta9JEN4uPh56obQxEEVZxP1VATciRhVojscdwkgqVQB
8guyMw3WcCUVlp/CTKnOrUBfXsA7xgZhD2DFT7kMAU3CuK+txBEVUZepbxvilg19
Fr3NWG+cyczCjnQO8gmUAIvhQC5jAfr0tAtJ1LnAr7V6qDeofDJwjUStVRKfQH99
pcFheBErEasyuj7Y3GISQjq91A7CbWpSkUwvDGz+ixOY5y5undxF0ETA0dM9YN8h
M0WcKp5KpycgIoPGaoGLdLCTfOyIdyGXYh7huWgEXVweW1sy9dZ60ihh0skpSbk+
ASZPHCM3sPSDctuwobVyD7xFDcHrvk+aYEQS3b9pjTW1ZOpNZJ7hmgXqcI1jdh2h
A8DhVYhsG7KQmQWyw3VC4+R0sqOWxl/Wj3heVzitgv7WrXeubGSFrhablZ5K0XnS
LFfjiPef02OXDm5dDch9CS/jwly+p9P4vrCABnrPg46XTWnVU2imu3SdXsPWNKCO
7egD0txkwoFqpqVhCEtWoPkDC6CHuHsGZXsX4LfH5m1FNugb14lutroYscgDEznI
t9rBRqb6NzgH8jbQWgt7VGR8NG81SF6WbY8kKPTg7QdR1TECR1QFsr4bGCRWDSIM
DrI7dafx9YfNpXdMOLdq8dzzyT/3TuMMeJSCdUkFv7pFljJBRu4zD+6Uz0hAH4+F
MK62FWXAcEnZ0gTxG7YqypPK8Enyj1nhvSvJNDTC2zHMOqw+//R/3IZIz88evC1b
YEnAKgKTa8wgOmVZ9zJyOMoXUE0a17Yt/fufC0auB9HwiKCg6LUuUKX50K54KFQB
IuO4JOvqMherVm46blyf6++ANt0Ku3oI9/yTZ2UZ9/xbXeQ2qxMsyNMc4ira+4qo
hylzLjnIW6mw82w//25N3TAtU+76t2v+HJSvD3lTAgO4zqp7tRpI1fwn1mnhfnpM
IdbSVIkLMdZChekXs3OS1mn/IcLCma7LxEfL8RG6K6dGAPRBmnazIo4tl/MjJZyI
NXZDiiXjxHkjdb2mHXxoEnpkW4P+14eQmD0DC+2j/N58fGlY9+HeNyoj9oKzDl8y
LIgDsAUfbZpMr0qWL1Y12nWS/gsKuHsSPxvZ+2hF1ZvPwzriv3JB2Hxr3SHC0yAR
3WZ7Se5KfsR7/rOdGh/780YMUzTxF4tx5f95QLyd5m5aiKOsBAc9oew9y4YyGnlD
BtyfZJeFeBO49fXpIrsNjzIwi7NWPU6iccI0sJOWoTgMrVuGyg0PsA7usE9ptje+
CUZn90QYCqoRruiLqJO/A7MPhXfJzrSFxl0a2fklPi6XoqWxblbkGGKoZWRRIsqZ
PHv1+7+KiWRPOC7pKCCU7O4bI7aQBCC08wM9jKywdKQaFFBjw+cT8vFe78PrxQBR
htEX88/WuoADAA5R13uutDpHcRsbzAs11loMpkDJAaBE1253qNm2ksfVvzyCiNCL
9choviJVTQm+5i4xipdXhkMrmpr1cnPyoxsUN3IJfhLqcMYhvrjNRTiGt9Hhcm6T
NOhmCDvLWPmpYAx298gQPW2rKMDR2K4Ip9wY8k5EJvVplP9XdBHmoW0ETKNRAH5E
Z6Z4xI3jlS0oaGK+ePf3FtEXjjasOTfGU05wZJQOB96tDgXbFHBFczrrOCYmtFGQ
99JfMLnVxNUROU0KHG6fGZQ5GNnQXotO2JVoXVCjsZ8ZWSL8a1qdgeW1a+SCWWb9
/91U3p4LDyKixopKBiFdO/7/d0gUeZAB7MlwZ3skLjhpZGjTGdYkMR/ZG1akKZYz
W6Uo+SJwsRmw8JygLK5cpIAavrcFOCNpgrz9/MPkaKscSt+fDisWGi37sWQVIey4
zqjQ/LPemzOP3oeYJJ5AVDpK7142+MmkrmeOyraLWVRJX+vXsTukBh44OjexVnct
s3xlit4cxIxqBstSS/1Irnb5UbzWoEIkNiEY5U4vN6f8SB2ijA2l6bSzEgeN62SH
2YPAVPtRopunWiuvLLuYvdivgggbRS43v1N6ept587ZN8RQlFB65PTHoXiJxnhQS
PbuvgRocpF3CaELN/UyNprzu8rBjG+DUOOgnviJt2BfZc/qRMhB//xd5xIbISoIA
CJJh9TMdLpRxQzy+N9iBAO0CV2tmKfLUNOaorP1GtSk6UOGk1CvnatcHM3pVFStW
3vnazZKXYcvW2vvzlLidbOThe4xe5wwtEfXv6vrcEin7jcjEhMS8sIiqY5o5d7GM
6vLC3G8durYsnZD8NPl7m0YP6b22MjxykOXmBM3QtJHyG4JU4pXThwlmVPoymtuS
ODHa8f6ln/dfB6B7t0xYDUu1FOXxWgRkeNUH6gDI2yuZ+Z26tReswaK0wo0t9086
su1R+TdoytRBm+8F70q+CY3PGaJ9aU2bm3xgcblGRZnEw1VBm0/GWOVX4inOq83n
6IGSFxGleWCuyXkMwxXpezlXmfuYHx/mn/VECKHGISkqL/jE5/BL0Tt9nnMpIWqB
B9INe/imuPIHdZhUNn+8MTQmbmTAMe2nGdA8f9JoeIH3LJSCS+t6J/7aeuan+5G4
jxz7TNKEo6vMM7bX5P2lKi5FA4UfvVax4Us2AH36EthhcxBZpVPagUB4Ays385Ap
1G2abnYN2EBmy45sb7CwnuvDxloRS27y5+EMA+Rl55KBZqRYeLjqGC92W7O49XqS
iaVMrZLAibNQyBUE6xKGAh17MqJNEjJ5D3iXCuUGQpw939dunpXODdZzhhU89Qin
3gBx1Rs8AaFZrRjkQXtA5HwGwrwNu7rJkYfyu7xT6RQ8xo1t/D18u6MhduwfHn3f
EF4mRL1vqGdjz9vPUpXX6e1h37J3Bo8eRhMAP21Vf4ceIklVHYoQnrAflT/d2ijr
csa7copmN41VbsK0HIjBaIns9y3OE1TJDlnuatxOpdPZ0vqN6ti47yn2AbYalgtz
4c+mQpZ6FYqPqKPFoWrtOqpL8da31iEJ85fcWWBHa7Q7E+SCGrmWdh+FWWU0AxG9
DrJ6b1vTlgMWqSPyCCRpPW6LuXOgmotHOeS7DOJIkQJwz/9ye3wy8jnfNTfkBVU+
lRCc/W+F+bkgKYZgWtXuxarn99mWgA2vGb0uWAKYuSukwTNRM+wgxtUuxIQ6RYps
+hMfHbehOcD2FKv0bHyDAJ+4YP0R6i7z/JzVl9K0aZzIVEPW9yO2qU0VfniU3tRX
0Nzf2aRdjB0AF8ZyQKZ7jayn5KjVgc94Jl+9SiBDdeCc2ylLnvstdVV6zI41HCPX
Oa173icYM5r6B1IMuFshivckJN4uQv84uQ83g0VuP7ZRTM7fbpEVgLWV0eId2CzD
BQqVr95xrGz4gbWsZdtI6PVJ3VfhonmWt9d3+IAOJyW8JSGf9nB4g8Ha0HGHIiii
pQQsEw+xgBR3DalzOpV/DtNXqh0fpLQGJ2ZAUMlezZ05lS7ms5pPqlkyEDqm1fs7
GIYzJ2mOZP/LiubmXll1UNQu3RiNCkGPw0CJbA2vV4ILstu6Hljw7cIXa8QRXX2q
yidYSGh2W7+5C5+dwhRWRX2vZ1dV/kgojKABgce40S68SgTz0ri7qrHAKPO+UmC+
CQtxYGiPqpzpzU74VVlyOSpPIacOg/He10ehzJ3jpod49FaiqPdj07Cqkwkjljh5
lyuTdJq4k5uitxg0EulPxtTdxkNy0F2FTI4CGGYJrEPf1eQfXSVsrIL3Rsj9kXlQ
+GSUjw6Z20bX6Gjz2ny4bDNVRE4A9qCn/5Bv7kdS/KTOfhOfGOhDv0s7ZYIOh+9F
Z6q8BA90mAYt8Q3+ei4PJJI2RfOdgzwIpRnTVN6YlDy4DGJ5wePxtPL3fvqLfi3N
lBXgQAET22+jklV9qeXXUN5/ukW7XlaDse/1CstAtF+z+rda8DkkE2WaY/7Uo36a
JT4f5+1vBxX3HWnjfVmyNDIXr/gRRbndVyMKtoyR5+fZvoFzTrEEsxducSFjqJu5
d3tUUjdUO2VYXoXZrCof1Shvn1y6JlsBn47zUOegLtJG8gFs6BgGlRFoahpCJxjK
z0CuxSkLS5+6lwZqPVkbNgFsks7yfNaKw5nd0Oyi1yiDM03YMHAv/iUk2/Uw4EeA
TVwjVgHU5y43yhLzoNk8E9IN1yxtEiz+2SpKLuC2nDqca8buG0wi6l2DftE09kNF
s7RLDHxabKmck/7HOmHC80+u/HTGt9FuV6p6Oc4sdSrj2nyRWQiR0KOippKJvt/y
3ghosbiZHzKcFqCoi1WuR9LrgmM71z4HhXIsZb8gMuDe5VYTOlEt1w+qFanj/r7M
apxa10Cir3xwEs2Ci0uo3iyP0KCVLuTbCTCRLt2WuJJDF17thcblFhReWQia5uyx
fGVUIyi/AJyKuO/J4LpfyWxS5OK4KUzIWwzfQiZqv6rgrZtZJJoou8WIcQ2bSmzR
njLROtAiYqKuB/VUbD/DmaMm4kY9IIREgGVkKF+59XnIT3yGjm7Ao8ZUM2gVR07k
+LM+2kTRRHg8eL4mFzVOijq1LHSW/YSUldSVdW7uKsYnN/VUTwb4l00NpMFB3mnM
TVQ+NzcezN0WGs+qP3X2POhUdxY22gFqYuKyHO41cvJL9XGjGFEY7D6F+s8v6PCb
MkWOcCKOjJUrQypPa5SjdfH/XaWntcUBYjN9RWdP2nkPdxp4OcxWhfKYMpZuYJzV
hnXyvC3MZFm3siX1GhOHi+EfzOzUPuTBEPAjidosOs9KPNvTciWbM/QPGXePFmUg
8hrIje//Bvjt4t3IYaSqMN0338sMtU6+mZUnw0ScxB3EE017jZNljeiFv5GKqofX
p6r/OGXb3usKkQzYC9QwDp3yo/985e1WkoAS98yl+JZtMU4RsKebg0o5ih3+d/Ss
I9k+ABYjRsIdigdQuUpaU+Ax0NERZ8HsQAspdfUDhxhbcqaGFAQrJUH8CZHcNhFl
kNuK+zRBIeDDSGo1zFr3Bh7mzvSv3cVkQZnim7RYZW16xPzEpUuMx1PWCxrgnyQN
WTT0RVsGlB6vVVyGhheIaEvHae/ZAdB7HzWJacYY/5dgRtY4mQAua9nQ4ZHzN83h
cqGVImEciY+szBqgRgDnrY4W9D4eZ5z+kyw8N8DaNVBc+ZOdISAXedCbT/l1aYo9
6BLCCnEHvrasw0kLwtTKn5lv3R2kaPxu2IaWd8QGaIdm4OMGUy/8xf7nnDzNYO+0
TF0NhhSj3qPJQ6UInjIH4o2+HmlMOu7qCrTYilL0fEIlI8Db2nyqTXtW/bx40Mie
mK01vMKM9ho9guGXQzPN4JaKjRZcxTjzm1rOxfvJEeSQGBdzPTUmSBYhAObz0hn8
kYbpboCI7uwvvBVjIBsWM5LFvUI9b49U2ZnqFSlNez+X5BMoei88w6txCWC16aDh
Gfrtl7mR5FvQ3l/68NCFMPrm4h1sb8GoLMJxNpi9C6Uusu2Xq3K2qgXR5BHd8LVw
78zFo0bCgSBqo3ZzZAGDudJRWcaztjdiivZIVjCAG5xF/N2ZqeFU9f5QbqyoIabd
CUhMoLaohS4cCk2R5YfSnVBPyPWNqzv5V4pIVBLT0yYSKphwThwDWB3ePnHYwdXw
qxaYDYWXH9GHe2TpoMWLWoLDC2WMzPewgd5gJ3vzVaBqNnmp9j06Z/y8Wv/rEgKA
fkKdQyerQCm45nHUPnj0M1pzbeXhMGAhIB+Z7Tv+nnj6A0Q0wjew0aJoUx8Dunkb
O/izVWBGpSSmKpANjiJpHSsbzq/uOexvJfQiAsay10iHuWCFb+DiYLA8mRpSuCou
xt3SFU4NbM59YsffY4z+lCkzQqXASMsDzqJCatiiYjCWCpUZmTb+STTRLju57usb
xWZj/HUwXrkxhDyWGpXqjzfRPtAM4Cptxnr1dnZqb0YTk7yi4nIREkRzaxl48Fvm
Dzuc6R5joNCVxM51ME/OXXRH00f7IumPhGD4kyLD3/Do9kF3Z5pBwxc+4s+5Tc7F
Vkh1jHLo/PS4E+jOUhUnlaT6BXwJArr/9/fyCTn+zKpJ41wbThTn0iJNSO83Czez
xl0MeUictsbyq5rkjg4mjJyOmWRxqbzj02qR+ZsV2LP/G7661way4jG1nVclQlyn
DyHjFuOcx+QU63Zsgj9v5hOeHae+I+aOfgeeqkPJxhcPcGyisl9vJhNfLK0BcJ2V
YbNrmrQUkfdc8FA9sNFNNwphD8WImfCRJw4QHnGQSKBOlllhwvdg/TPdbecX4Chl
5kxNjoOpjIzQi9XqHQ2lRQ==
`protect end_protected
