-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
N01auONliTIIKXY8UexMuzrLygrWTL4t2I1a5RC6ZxBlJlTT4Mfh40qogZKCr2gN
VWn0buxgNXkJ9m2nuqX0bCEzTn6AOyf5RVnx0IBpfBw+9IV0bRWEVbp4yPLBCNML
zJ/OJxWz9adfe4c4xqBTpC7c1aMfcJzwuMh+nyiw5HA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5100)

`protect DATA_BLOCK
NAo0eF6ZQ7RartRVtvbDf226J0kiMgbnZdarH4xS7atg0Ddo5vbmwKAdjTNIJVLm
7BglKcpFJQo3PhVdCkAtOsGHRHfo7nzgedNKHcuuslWEefrTQb5ruwFdTJoiZdNM
84+LPU+HniYBz0Xl7sWUnGX75FifOIFc1+hf3TiGzQxRSuosEQNvqig0FesmTVk/
i9L/oSGh9YmrRq3Ki4TcqAMZ2gBDdG3pY0aSYBXhCP5G6RYIGgFpe6LWBq15c866
pTLNfKiDKHRF6Hm907cpIkOli63wOh6R2KNBjvryohglRS+Wd+X3lfFUm2kS6v1o
lVN50GeLOKHlzp7iFirrDMFo78rzvJdZ8hOU/jgDGF2tJDexzE0fVkfn5ddwlz9K
sEwY84D/EbpPpdkkKLm0Z+8TCbbEJVB7/4aNM+Vrdh/tHBairnq+VEQr2fh9u+eu
FlYoLJ4DjHAFQh3cAdjLbx9tIZoHmU+8GSjpateSYfPtKN/fN+bRrQfXtUGW2qBq
rGyI6uwoRQwACYfm6oIQe8a9frrtxizQWqWloEOzivEqW2mftSQ0AxwIIgUfHfBp
939h+u5U2JH7WIJQuH5zaNGf4ZuMPZraU6+Xt6STQl+gMd5d0LO3mZdC8hMpjb69
d9caQ5yA3nEzGtWFEEliLOhlEv+8RskEVwLxSYv4i/pYsl1QN5x7o2a82VpMfMq9
boEszJ5/a0OfuelcRODyZ3ys8HmYFiROiscC5aJeawmig2s77O0b1b1OrZA408Ae
ZbQmDl3JKM06C5Z9lY9SbeM8v+ciNDlNcywg33pykJPdbGToLhhKRvbvR+DDYJ0t
fhLgYIn+5/1JnkPAjIP72reaR7YWVl9+NWdM9EKvmeBcGCXBhnIyJM5Z7OErZYwJ
wcg+v4PFVrGalsYaAdGZYs/8WppX/ciHBfX7BInM92R2AyZW9rsbHqRYJGsMXA6T
87wjo+UAeiB7RdmjSqVf5mND+QPoK3inGJmTowad+PIETNB+OSiFv1OOgwWbDFGd
FvoO9B5Q4OzT5cW9LEEBLradEk8ObP742IN0CMzMM/ii9HAW1Mwvc//0tsQJYElv
k/heNxALP6zfvrNAZPRc7Q81Dkgr/rPY3NDK0nE6mkFe8L8UvRkSFdkTVtDh4kfh
VacnAaAQQiYD/2PdQF+/nUJct2SM6f6wX7lzGMp8Oo3JVR74pjYdUvXuT94Z5sll
ISULS1xqkiM2iMcBaGWr45QphI5HjFwkmAEz3GGdngEM2bFkL9vJlPKjcFgXein7
Yh+fwikFS+ICwStrknbpSWgYcxJCpFbkTMu8Uu7nA4SjyYTLOhP2dEyNbb+CBlEh
2fb+AP58GW/uQ4baXw3Vom2X8FUtJdiK6pu0n8rFuWknKapq08D4I1vJc/yVo+ov
iWkPY03Blq36cPFopaD8Z9XuxKU6pTPBaUsKMOKxirPCI7pn7AoW6vW0adJ0ZSDj
i9po010tpZ8y0eOuTlvCwBRle3xCjpNFt9XxNQQCoVroyQVhaBhuPA/NJjUkIqu2
t1DG136GrDiwRY5gfPwaZY/QuBIAuuwvxoZCHglXlJMFaTd8H3cIfBg38ny1TGFc
n2pboGMVXFGaMXKwaQOLup181JqQk428bBXlUWYPstp01YJkcAT3fmJmjP8bQUbT
3nKwC1ewOXvCkreM0GxAhlqO6vYi5AZG+pkiOxVvo6/WZvETqyu1J/U1zCo+IA7h
R+3nVOtgBbn1b3C2WUPyiBTJOcxA8eXgogKtzRAT7mqOZEgFkPJyUDvp8D+zfjfN
ffFisD7Hfol7Fo//vug6gp42xLarU2wxZ5UanG2ylTXji5DEbZi51GVuI9y8uDRw
lmtxXzThYqFBoFk5XPnJmmKVxxm5QN/WUnhnPFlt6b9BLPGVoVP/g6VsBroyjXDG
Si54ciOcDcF/lQ4ikhu9yj4B1z2it8zSjlwM37epOy9WVl3toSId2bxzBTW/IQWa
8dFX1XyO9G5APnrPcsFb7Y7TEakd00JPI/gqTi0aCU3PAJ6iYnaGNVTvKF53NE4X
goTNORx2QliXQ+natNDcDr2yYeEkByQRoaIxq305dSGM7ANYW9hOC5G8eZdHzptk
qvBt/GeWQaeM+etGmDN5i2QoQ9n/4TcfzfEVv1y6jPVWW0kHlXnfNlffSbm9O76P
fJefSiiIvYzwlKsX3gt2MWTxZwCNEkZ1Ld2K6XcaLE5p/6267sk9ObYKv17c+WNl
tLROPrIIyF7Qn5euQ5Q4jLUNTuY45H1+LRJICvKOp1XDfkwWoKhobqhjCWAtU2dg
6eFDSVhybRlAFqByB8hw74vq4onwBvn5U9BmBbcmDDCDyItF/ozGLrRbXump3BKP
5ZotY2Cu+ZPGG/o5Iw4m3RCn9cLswkLLZPfDNWxyK0VHm9++rxguwoF+gICJHSAa
/2PIvT46JQT80Nmg0QTKVJgQC8DGmg/89nmD2lQV4GEhEoG541l6CH9cbIKAn9Ba
HSLZInwypX259sdwrAGGU25dCvPl6/NSOHhaTT0wFf8ykCPFR/rugKv2JGoBeBKd
HODTL8CLNGqhGvXzGKr7hh0zEee1BKiNRG02wI/ZsDqtpVmOU63uRSpsVig8PAW1
SyimEcZZKZBoirGrxIfw5Qx5ohSb4v0bqoIqTNlkj10sSG5QDc3Upwjx3UFcsN8y
3G5nlY7mQT+GONbwOyh8BAcvcY32HHsB+pe7//dMS/2uFYeEIsMqND56mC43S+qd
/Imh8Y3ikYEK8/BlF5FqGhAIZlBTz9f6IB9jT+iNf1IofNNnucgryACSQJrNLpxH
D2Y1oK2/DQouVD5x0wAjnOTi9Ud9Y4A0c/ONztYod8tjH8Q8xsj5I9LUXNHpVpmM
8+C8G3doMLIxOYnpwKq3pIhQMK2gSwLQnbTw23Gd0wf3W2UViuR08AxlgBe8oZhm
1WPJIpbVXzPN2FmwuUmqxsRCi6F3W5mZCags2EWoyAMo0xx5CwwyqXlGXSPyshXX
i0IZc9FS220drYpxBUxNmoc1CLZ0hnHRLllE9rGjhh+H3VKZuE+Yx/17FbQBGDUq
X6fEzsARX1okbhY5DPg6nFuucSy9vj5AtY31OwWAiR0lAgwJApdws1uLnVHwsvRs
CkpusLEGns+tlX0+2xoeEKxc+yqYXcIrt6+SlnKVkGsuRMA4iZ5QJGhywMZ9obL6
TaNWeeXVkUkMpBBZKoj6FrsI8YS4oA0LrJ5c1bfA6C6tjuj7tlCHEfUkaroG2UEh
TNkbKvfD1PBkbpGOf8rqiUSoYLFLNVh2OcxMMCCSfmFvBzVSsyL4ha9A75qV0TxQ
80QbtXJnQubYsTxIniEhtxkawI4tZKs6tQwALh4SaEaFaebafArBb4h3y9UfO8De
ARkZLArwgQ8awJ8e4lFnQ1LYXex/tVyMrs9m9mhF453AMimMFf4y8+rYsUjfrvNp
r0D0vtINChrBBZ3Qrv8omg2cf4Bz8Kq0zkPnjEPSoIGMyLI+F9MpU4u0qbIVx78I
zyAL4dhR+6W0uWioGmkpe025GDmJ8GkI135G9GzZ2sFfwbNPxfXVdvSOHv5ZVi7o
Rg+BpgXLENm1qX63iYoONPeGAHaTiO69YgE4g2FTY5YSJTWIDpqODYaJ6Sv85e5c
j36McczU51u8wyEsoBeUVLb4bM+vXFmGQpprJ0PHuAfFIsMW3oU5+16FnXBqUvRx
9YTJJnL8oVbg0vn76BTtJ65iUiG6E7GHLJ7Q+tKbxpDuWi0sUVMzYQzFt/2QAweF
xZrxPvyeTmevCzJQFyacjv0AKllYN92kw7dcAjyWGzh2dwDgprjm6JCFGAmNF8e8
jhz4Si2gKdRCQbOu4OmO2R/zg6JiQTD72dIOqNNGWne31hwbt9GQaXJHYFh3iwaA
VDKgl5u3Kbw9EsFQYPZczH/WhQbkPwH1B2dge8CXG3RYwLUhh9Dgx8MpjCoLWlH2
Wzu7rbelMQy/bJGycBPkMHFCUay6tNVJfmOp0pF1jXWCIBsNLOdE2rC6muuAhYkL
4MQRWRCGX5jlN9Croi+8Ays8FqfElIBq2pkbZJVoNo/ak7RFDcGasEAf5VUHMvx1
vJKpZYi4R2yexGsBLgySJtv2DAh4JwU7XEetLEq4OxfCEaQcH8ptkjI6yKZ5Sho1
v9o/4kvLN8ZfxUhWw9yJ10Zj+is0MYJ9FU9jh9nr5eGzU1m+T45KOzvAC8FhYZWR
Qzu+6Ki5YIcaROM40kRxjMRd48rwj8yL2DfaM3LaRIkUld8FdxwowZOJG4edTGJ7
YvcCVTssOhsBmdLd1E8/gxMVc2lgHjVWmSdejEGdUJtmDNkQhlRteOafkcTtYusw
cigxM1b2mnnmn09rwJIDAbHQkI01K6nyE8pI/O9+Y69hzxrytywxGHKOjpmt+Ko2
JY/Nq5KQY0wvi/5g5eeRQoMpPsJqtYX+DqzYut8vHRFQs+q9byk0eHCNJv2lPPgL
mPVOd/OpvmI/HVe+WH9P4WpxFnyb9qONCSTNa8kEFHQPHtRAth60KtyW84v2l+K8
l1Pi9B61VcdMyFZm/ohehuXNUjt6q0MAB1/aDbp9LM7P2inyVZiNjngTQH4qw+gj
Ajo8b2Hg8pRDP+fp8piYEF8AZO5+b7/3GM4YoGPAU00asfHelSv8eKoQiCs9KHKR
fsVlqt9DNDgFbKKFmttcNTVF/5/3iR+MZEwlbei8lWZmo+AGd8pUJPEV6OgXR68h
HitX+bGmAxDdx3Q8PecCaGi6jRaYHbAQLnaSXWe+rtsC5J1vtQsltkieaYcGy/4C
X+bvET2QabYWDVO6Tv576jECSsU91eJB3iB0zuW+Q2iCtMwNeFFgghnALR+Rtktn
sdBqlQi1r0/CmSKViKrhw3cfvqmc3II9Lw/5XIMlt8sFxBzZQVV+82GGK7pjrBT/
oArWg/gHhj1awej+GgxqV5adFcOtWpvNHLnRDHIs9j6AGEz+SmqAv6d2A11PBTU3
AVZjlFPNbTPOIKcRsyRX5xU7FB/o56k5hXQkwrsD73WULe8czuUHDjAt3DTj5W9B
qdllUVIMzT1BpWetgnFUZZjH209yxPf4t+9gZNBkvF9D/R1bG103QxQPaH/y8jvD
3zXnSbpw6j4+apdVgsKC/0Wkvlok9oNSBnkuYt+Pu1s2gbjjA+uHbV16HG1zKYiI
mTKH8VZJVZbBlSxQQU3Ky16Q23i9mehMi4WVTd8ZR1ignUNFcLU+tqx8G7zE9P8j
st1FB1H96XXynzRYl2bfL0TTCxSKMfEn9j0wwtYRX2gjUSo138Vr4YUU+/+1YZzI
VIjXmy/+z3Om8V/vgDKqmdi0XuviVoCvOdyhWbufiGUTGm4LMB1+Jo7WXQvUDpvi
Q+pvrRPRek+AF9zSiV4fTwT1EaAsIwKVRoji/xBw0Ltv0bCA/ckoAp9cF2UR4p+A
XRfXyHl6oY4xykeG7cRDLJUdtbzSrK72+s9U9VX61R/bUsdIuk5eNrZnHt1bJHOg
2XyfxUnDryd4gQTupytMyDpXEnhHEAq3N7KIY1lgcTSF88tXKUWy2efqVMtgF5Ly
udnh34qYoVn5NEkKhCfBN70kpt9uBQ9GoSUuqlzuM9hznqz71ysM39nq02vnW+YR
pTGK+lbG3Yx41aQgJnrw1vs0m1y3Cp5GOhHde/6H+PRdzHTZvxnRv0rDWb2QyCmI
y2Qe+YQKI3Z3hsg+YwBpPFmT8GDgxxU3pzWdRo2WW6Q9YuzYneA8aWujI5nVeGao
mvVNAzTkKrsssEaj4RIHn4cFJfNk5Xj8nE6pdyyf/2lRoDK6FrOaj5Og/OG28YGe
FB2OYCwxKbmTJianEbX0t0gP+fR27ujaychG0Mh63Ofm1SFY3tzhTkhGwrZwh450
brYKcTsdiTPAL78t8+p2FpEGNdU8JZcLIC7Ug+dvREM1lRSEqCqFCW7lsMkXoVdh
5UEq3MWXZQMufmJEqh+d30KLFTIds7IvjccZwkXXBzVuDLGvXR0pIgQtlgp7ue3C
Arg7cwp2he7/868GHEXkPtahFdUPkQfiYR53o8MJY/jAO3vF85DWpODJhYbP/DZq
JsyHVcHSbqRGDXy9b6TeciPeGP4kVEKOeQEzBvztsSkebtcU2gA3a80MBdX5543P
J4PbORx9M3VbyIVqT3DMcKp9gufLOh9HGbh8B/0di1KFjsjSHyVfcJO7VjpVFsyK
78AHQvJV5imJAThQYq5Ofd2EUD5dUp5diSTLQmGSc/lgwm1SXXk7dH+PqCt/ToHI
ym9nktScFhn/33YJNrpnWJmRXe91o1X+hRNcO4/FMQaBrRSjvTblluM80FQ6ZEUC
d3leVw85jA3WdoYVbQ0kVzkIiUL/BWITnJMr8r4wDdTGP+Vm4ZDYR9+nRWp2y7MC
MXPvDVpO3XvuDJZIXlTc3qMgpr7uIO4fLLQ8ON3/pjusn6jGO6Hkd02qTCmAPYoZ
AkuL2zMUXlfhxgvspZSJCjGOw7w36Th0yLwh1d/Iv083DM/jG+8yCbsx/9qGXa2j
Mo1oEG9sYyErW2Iry4qQOqvQOt0tqNoaxT7mV/cFZdJIhbcZNVJHL8siHQAEcfuc
ppOG//msfcO2INQkGmI6le2jTPXITXGruEDswkblmkCRo0J1Vgs9ou5g/EDl5n5S
zLY0oDxEWHPg3jRLqRIB0gxuk2H9giMd+ESD70UprSkc8W9zP0fw7UzZehYtwJLI
EHGEoV24SKNrYW4vwldvfx7O3+57QrxmmyBQY26KQQXzuAbKyG9g2kyV4Ri3klqF
cXqUqV/QdJunG5si5wOdHBijQRxpMLoFCjfM8joY+Ow=
`protect END_PROTECTED