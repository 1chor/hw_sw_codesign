-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
EorAW7imaSna7ufdEV9H9rrxjbwByTEmHY1faJUfqCvgb9gngl99XNqo9aKmYJhQ
EgoFLOzalcztRIR1m3V0iD35maNKuwu+JS0dKJwlrNQqMSfW0nwaFlN6lzRcvcsg
n6oaNlvWwph9VN2rhVLXGM9Lor4bwmtRwrraPh+wBI4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 98328)

`protect DATA_BLOCK
6jj2q04UMYsffCssZqGPtRtdGe4ji5G1HibYF9dK7yi+Absg7p95kA8xuw/sG+AT
CgaNguTjcM2Ry/b36ia/zmqYlDl0MrVPo8Hrxdi4Sy0a+laubrSOnNxyuHkR90e+
AbWLZaGPUcm39Q1U/xeNZEIx0Yy82GA2fT1PBJKoWXfQ4Mq6rrjwa4kaccU1e5Sh
VUGy6CDmyJGfkCSZHqv1IQyTf+ltgOPjEwwNgIG1A3X+A0EEjTO6u/++3uFfehhN
112M5uEEJl9eNEZSPJ3LY6+yiNWrUSTvkOq63lk3IauXemm/R3Ub4Syr+aOtn2ze
70KcKhvJhX26xbCMTaChNHKPVWAkJbuvzlfa/NxZQOJNNnNJA2OheEu3Z9UaWpKt
PNGmj6NqFPVGZuuEvjTn0jeggybXYBqzZ0KmcpsGW10rjAqEXB4BkJ5gCsh5/GLE
Bh0sNYlTpikpbYCFnYCXFpavd7S69h8tX6/zbQtvub9+CQWHD7FeY3bfTrRvpQ/u
hGTt7G3g8X9wl4naB6rtzS5idoXx1LIS3b3XGLJvYn0AEDq5m1gTb7Q+37izKPQ9
lS0eRyulUbFZwLgw3ztw/a/o2aEJ8H7KuSGwEK33gHuvDFxIGpE2/b3jldjGjbu3
tMZmHb9agsVAokepbmiQAl8pafME/AyKDYx+LcbCrgfzT0oOsj0qMbF8p0irkcRa
/qIdWgPy6aj/X8XsNusqk4qZqS0Kd2tsRDDnPJ9qy2ZzGSHBHlQd9bj8mDKuqNZF
eVVYdFNrnD6xrcV9pNJeQNbWXy35t/6mGaSNtVj2n7hUUt8o3rIKqQWVELNNgg/U
HvC9kRzaF4V10oAN4dlGUZUypRw5iAfc20Z3gV0T9SdoCbU/p8PjBuJeLlKU0fFb
kPgUMHqDnpPpiq8GGJcqUzeYkpq0ZBRgb+V3ZCMfEnOXETPqEyL34qBb3ArV1f9W
8JCgav8loStdrnMjww2j5uG+xmbdC2blZE97fAVfZiuLed9QMnipaqYwlAROCsRK
ypqFS02SUbqvmFVYSQErp18N4a2uUNMrJaqntm59F7l1NIfLwop1xMzipsHcuehz
WvKAVbnwN6jFhkvPCEz0FZZL2r1BstNCyD4ekLSvp3Ypbhbgzu9jmoRzuv1jiEKK
jcYt56DLpxYQ/9mHJgHNBPGeWF+V9XzrMj6pYR/ONDxlh9XNdN3/JENZtVo1jr6j
HGgN0Lhnc3je5gUJ/8tGQxj9/hR0zN82Gyfqi8b/le7ezG/xpLt//9xP5n9VNg8w
IalDDhMx0AGg1vq9Eg9/lmcd5AjISp8g9r4fQsR9u7hxl4qlbzJGxHTLNNVJdWW+
hzRfATPtMHY6JXuBguq3uOt87zt9mO78e2kCpYf9mTko5/CEi7PEJvqXfJqQF5S+
nBpdqKJbi+SglvkejiWOSpnhWSd289142c7qouWtSw+Ux/7/fAa3tvwVTWdYbHGA
m+30O9rHa7S38H7sxJ3bu6zpHxelYPz1DI8JWmneij9sFvu9NcraYrFJRz4cnGWd
+yMPeWYBvl9clYeL4Dv+qDhaWquQtntYXaGmKVh1LKzoeYQRbotnKCgRIwZcP4TS
4shXpse/YOyKdvIPT8f8x3kCutSd04r902D5e4Xft9lxa7M+c1MjCHyDwES5j6HS
euhwhZ5QQvmr2yeowQBc0N9qpaT1fJ7vWh0XRWssqtt1xV9sweURImjG38Kdcjhw
5LMh+AYfjlKZ+MYxge5o4lpJaOFiWpbX+Nic4BQshpUfXUuz2LNIHlA/nQFPWYDo
uvgy8BozNjqJnet9XLr55r5679EiBzmfJSTP3Vd49Acq3LNCWyEYB2prJ/C56NMT
1Gusevvq035AKUjBAzGvyBZJm/Edd+xXg/3XNBJDFwVhKUZF2XxEL9+XyOQni/Eq
fd29epyQXnvFo7LFLvW4MbF0NIOJYQq0h4syDR0xptsqeSUM0d4CsIckEXGqOE+u
DxmUTkgTqi9ULtduQDc4WsZD6eH/LXcoyFD4heGdg3LcDSazJvb48ht4c8snOTuv
3qsfvL3I4MCZg7b0a6txmtk7hX9BBD9n0KvRLO4oXmoAWoHA8eS//NT4Ylu6rrUF
+E9yeetlGS2fy7T7kv2EWcCN+1Cfbg68ZYfdRdl6djwRnMrmzd98Hz/Pb6Ovc39J
wCkYrz9VT+XQNWegLssiSqvhFWZPETtKWCQUzGOczYNC6ztB6dJB2cMFYa9P+hcs
AS07q1ewwVrYHwCvSMKd17bEu9BfBSduxcbDaowkEIa6ydLDrPxvdkTQzsxHcdA0
R5zStNVqK4ZrqWzBoi3oWjsaigCuVb2BIYIO+3RobZkt5nXuCdbsWciTsdZl46ul
wFqeKSBUjzslqxAT11pfChDBot32kOfbxQyzcE8n9XP5NdZ6c0+ipFNFKcveamtr
zJwdbNPjlS/pf6TgvQ0/00avQKY/f8c9KxHQ6xdqj2xrcnsOofIZxohph7AWW0sk
nZXWxCNUXrAptREuSdI/B/uRgWqe2SHgL8q+jqMPZIpeUff5OLRJisLCoUigC+1A
P1JjAYWzGdHPbn23LL5D0/JVBZbA+Af0C1cLESOZWcgFqXmXSBbgCu0nJ8G6crAv
PiciEnR6bXc0MB0ZnYtxpBKouVl/NNf6W75OxtcKjVTWYfTNtsnNmqz4bQ309BV9
Ms7sNSblXneUUTLqQRu6V7aE+aqNcdf9O1PH57MIEejhizSlWhDFNKEJ8oYwqO8C
jtCt551QUpQwPp8Ywm7+5eSQqJSW1am1R5JMPEt31vTQdp0UuZVsWbRODqlrikKO
LbPK95CxYFIaZjbwpv2dCyC9Lqt34NLNdYIefBYo5/DQAjIP29F14RhMh7YgwvWM
tK4qb0CWR9nIt8aXyjzQJu2/XlM+2vbJN/s0OW3vq2eqOTue2urk0nxFN27Y/Twb
4xUBeMam50KL0FOcJZblyFnFaFQCNjuSfkAFKf33AR/mQzgX4uHg3UZ8X03HpCbq
nz+FOoi9cMhT0dJQPJibzSBmKta90B8MiWw6SXdIPzGKlwMcCVLj4CjBo6fkVS4t
uo0ewJfilfc7ablUDi51YtR0felAX/zulZ5YII/mA53vdXBDHJNXK7vhv74kNfUq
juZgCYlugTEMzsjp42WrboEfIP4l7WYEW92zjcNTqrOh+VDu5XNJDCUKY3JCnK6e
qQmXn6tMaSzhIWZR48QqFb4VFVIcJ1Fvy6jzO/hGOd/j1whuTe1rJGyHQG70ZtFw
IoLvfmhKC+WtPKT4sBdywm0ERZ5bv1nSLPJKzizXZsEjUAf46cUciKZWmFatuL3N
clUtKCeuQAVPjm3ZxuQ4CNznkeMLI4t990JktwkwysVVs7gN1U4me74KwXdbmKcp
WrYM6kghb+qzRmS0s7uOtjqeV4rUJCEYZYUDy6FHi4hmHGPNRcOAORgcxbiWp04Q
LtIgKBELeksmGNGbuIL0Z9W9r+ucLf9UwBFY8VD3IOtXgrfQT493xDEliSYplsvw
TV0befHBnooMWQGwx10xIzS/7Sg9flIHNtCp0EyGxIfzcaJSrOvoaCz0+lyf+ses
MLcbz1iWM/23f2lV1gpFEwd8Iv7wyclUdVu8P4Z0nCasmXBkPFWRc6MGa/Y+iqUM
h8qwc+6Y2+VfBgV8viRiDTRvTaZzjFN/7wySPZY+eD6TNpmZ+mnT9aEJ1d9pW3AB
XKIwYA8sXbHXHznP/TUi5hFA6Z+leqQtjOTh0aJOXp5OPjNjGwpzrL46cxqzVkcw
Vy+nTbp8pVZpKH+K7LMvVVscSSksSeFK7+ICTQBwN8VgtdUOse0/AAQdMAVWMdSc
46c4KOxCtkx1UmK5DWwcBNu0/OoJn5cPLJ1tRpjVb56QfXKmySb+WvxONCiFVxRZ
jh1XusbhY2XQH0zzKDvTZHjqdTwnlV/+8JDqKOF50ifU2IKuGnePnldl2aD1DwO/
sLxck4pearYUxfGE1Bpqky49dSn9EfeqJXanvYK4L3lZhPKyanOCTJ/bTmFaETdv
6V7wjWc/nj7RBEBtbTM5hd87c2UPcNN4KrXS2zdSnQ1S2O5M+PmsI5ePow+M8nka
AClGOIRjcY7c7xvrYtOteiv2RB+rVWSnwIdG+Mi+oCYmu9MQGfsaeA43rytejRXB
OsZRYsPx/Iv2hE1a/GED6ltQ1SZoENO9WAJXGUGbn1qo+TM3j7mm15auiOn8lkRW
Knzh0YDWWRqllPo5cvMkD0HtjhSEXQi0XOkRsb+RZit+5onzLzx6Iu68mJeSvy8E
3kllZIPngQQrX99Dx4Fn/BcW8uciAT36zgVtjUy27hAQm5d6lFFtGLEfFAoNg8Wf
4hGzKJRwv83Do65oEiLdeIMv6eIyk5GUuAbYVMGaLzOPmS+bs0e6XWGOduOYvhsf
1vTGFLcX3t0i34O1UaCVBqWzB+qbjDV9OaO3qUOJBSSrNLwd5eylj1OijBcMteNN
COD47Lpq0hnRWy9zoGPbhHjWjWyMNE4ZX+FVoJEivCI5YQBzRP59fVLopnEFwS3p
Rwct9BoMO2HLoW6uHbLNUmP2YZxR62BMqMXRgUvnc9RcEZbTQZeZLXj++3ObyvcY
zbyT52bCl4Y9AQzOs5Q9S5OLfQUik9LNziGXV6VyIXsZtAhwN7kyXkO0WOZi+BpP
PZ0lX5FvcM3DjQ0GLR0IEPyfbg+5QbtjNAijB0wL2RRU0wIbXg4Z9+28Q5GuL6OW
0A5iIoOJOVl1nzUsjmhpEf2C816vdFYCdMeEOCZO24GQjWGBRVdCx7suvybKHxx6
M1cbuN7GHJ1GbxpMCnVjCpZxlwm5K87UB7e3e8sfECsS2Gyu7XTPu8/S3mf6ULgC
a52CX3/Cp9lAmfKujEeMHcARVpG1wbND9crj6zfgKEZpBY/2b1HaYwGeXixvIBE7
k9665XqscK59H4sNbSqS6Cktw+/Zloh2MMMNf6qb48CiSEuLE29cul/weCUJ0Iki
6tpqh7NHYav+v/7gBMBqiV/Oz2h+JMyZ24LydMinZtfMbBtufzJvIfIwVigfQAlX
sryQo6rf6fAAMzv+c222JQfrYEWspuRkW7CknJw87diDB3OFe0sBMCBZpEemwF/V
AbIOdDZabguOkY9PK57ivc2faiKn+Nf9xCkCDmjgE9lmcH6agwpO/vlWI+Hpvuhy
WtkjhEwiAFfc02sLelChSZ6fuXTRfO+UAPglBKqOgizsaete7OemmcFUqe7qrAzf
qs6PokYTZsqeUBkwRTJSyJCP9xX61BKHJ2CBU1my2mQROISNxxMT5uLHvbkAl4I2
mVPa2fDOP7m0ZMT8pYyUoGwVEdbwvsJcHMbV3G8fBgptCJ8Jf6b+6bfG5ezzlgEC
/FZ/QY5XkkUkyzpA9cv8ryKyL+Oj/lkQvKPTDWOP+K8XnsW0dQKNWAFIUsqD7sO6
lmaw8U9jb4kV0BTET3iSLw896hv8Nyvac8dfHlQn6oZwo+Z4biA6v6X6GQM5eL5i
PlxmAe93ISPOXpws/xz46JQUS38Vofs6gDfepJWGHFj1lhcqDkvDO/FMgda3djpX
qSeEB03gDyQoJW2RrsLrwUxHlhtM//H9dLRsY4tjW3ZqTCHzCAV4tDfwNgJXmQeG
tXJDhLpu9xProl5oVIR3HzFJWq0FGeZGKhniZLyiWIhyAtD3I6NqF4Rn4QLyPMQW
co1KY861THE8gSylfEuoHdjOyTUTiIlqSKuVn6l0H3k1EpyP8lzg2LXTUrBffJTl
cNhO8oFT+5Br42gpO6rQGAqo66D/c4ztiYxtG9uhPivsXi36e9HuD3Z/rjMZBMjm
QbT0D5A3d7Ypq4qR7pLmoce9pzkIDC2+4tbkXalx4AEXh4I0gXHf9pr6NjeWzEbg
jet2vn+hRPKT/BPXZlQsdKyP0VhXl8a1Mf73xWlZnvYyNa/OL9/i5XN4hZRu1Vkx
GWMg0KfQoj8oCFuKZhb4yAO1VIKj9uBRr5zQFHfKpvcKm1pzNoaLavrgOvsqIUhH
aHIHOnLRNrN0AQWDfHba9RWq9yiQfIKoE4UmmPwd+9FfVZCADPcnPiX5cZXiiZHk
60Ox65IpQDmqrkGVRQOC/dK0Zr1BhEID6f2g0o/rcqj4BFPbxabhb5OPqaJPX24B
3rS+1rMGZ/ra9y/NKmGsrg225c0qkQSlEMU471DfudzU8AyA5Pft74SIhVGuw4it
djJBMjavheCrXEW8vZ+pqp2wl02K19PrqQ72jayZFNP+tCJo1r2EYQuExfN3Tida
x4VOir9aXZxTgR1QnBD2gAsn859+zarBbvL4iC6MccoU5eSN5Wh4pA5QVmRxgTEh
VpbgFEGF+gG/hifDB1DQewg6b26uw7YSpA5ydVWmLtA7zbrxKD4JUxzIkrRbjT6o
BKpvBWzXc1rRoPrrRAfxtF1DhNkYKhlYPekvmuquchvchaIW2xUX5uoYIPVrwPbw
eTki/79i3u5fI1YwwqOlUwXIkpfax6yWH3Y+b1Nax55GwFfXPpJ2+M7Hq1jTeghL
nELI6Rz6utPZhYCX41rSRDRheuf7Gfrjrn1edlXBR+VUXRD974kETwdj/VHqqD8k
6gERYeduSCB8wSt+oj+D3EF52SS+gzWX0UI3da23Aoj8nW3/0KPUfu8XrAkJyc1G
WWtuFqATwKZxuPwPOC/kcO8SJP4x896zDxE03eRKC7TanR1eNK0svJHaP1Or8kLe
xchq+sUdO5PwzgYrZJPwS5Xrg5aAjXhtGXlvHNjSJ7GwneC1xYijjeff6QCp5Wut
LnEMqtOGTGGBmfzZlLsHXdfjxG5xRw8ZwwQPJfw3C+3ZSw3FiJ8A4qbK+jJmT4DA
x+3lRKVRONaiP3+Zwa3p7j3ENbvToUXcY6wnmxz6rTMP66LvoMnjxxKXXDqvQ/C5
Tjwu6aA8MRIOvsxuR65ugFwPonehP57C1XWntQSHw6QHgvZcOgHcN+1wHfiF8igk
8vkUTl9AK+KQbNmvsgVMtW35zL/JoUbWGt2mlv/m5VxGLA085QnHMc/gAwbqQuDZ
DUK2ASjm0xddBuGdz1WSKWV43lzhGsK8B90dn4MTA/qCXh55p8bolzm0torRKzxn
3fa4IUwy48pOkir0HEoND1GCyoTh9gSVxbE/y+uim7lktjfoc7AdVZOd0+rbAPTn
lwu3uVf0lpIyIUW6J/+qSdCJT0Z3VFzkwiSSb7Xkdvp0R/+Tkhm9FR7ZEkZsoExm
eMH88ki6QFXdFeDs4Rl5lLlRkJJrhLGr+22aR6u4WbIWFzsblbc1M3VQL9RmwMh2
ntMI8Ao3/lJOLSp7xWrxO+0vLCSaTY2NDHoJg9Mr9WI7wZTevbENreo89DnlxBX1
qiCu/+qikvgQwT1nS0XkENhogMCeGU1aJTjl6OB1AW4Nm7mcgRXDjyMJxIH+O0bb
p39450eX9k4nptBWKDhYx4oY49l8AxubfxBDY/eJ9eyvAnxTfxX1pfIydPmHhQcW
KUIrCrKo/36Y5CANK8YdodkJuHefM3ZFgE4rttNQrWtctOt4akjp989Hq4/bZBla
7BacuyDHj+4accD5iV4KaL0DdXptVSbQwyDo4sEWCnGT9QGYZXGAvlVq8ercjRDv
vHoH8s9fQe6+uDsew3TN12CBw7KOspwoy5m2QFPzdb1RbTAzRe7MyaG3mqRY+DlQ
zgjzTQii9WvRhUm/C7S55pYo4cIbiBadtpcDvxH4f4U7BSQBtsysHYd6lS5I/SEM
UYhFCs1N42fYJCE5laAyPEnl2fdEQzpbe8mt/5hHhitwc7hvsugXWR33GCwwdUlX
MaVT+VgCKznpszce7Q4ZagBFD2WNNRzIf4a06THahJcbAhfM+/b38LISlaOtD/84
4ALVfMNLjxTg9o7D7oa/2Rl3T23vxTjluvXF6FcgYqLk/jyxsPDtqkMgWJppGopC
lwwIefRFCwg3112eAbk1h94cGdntBAW7DB+bpwT0ZFB9wpI3LhT4/G3EYoI9Cgyr
u4DLV3Gg5C7aYirD9E9cD/fYRh9aQYcmHxVq6WZbYvQ6tBVwSUY/VIuhl0FD2bMA
QWycDf5FxDLWHXEQT6hD33cy5hNPqvehQcsvQJY/jLjiowVVqekbCgYpnPdQiiGp
GZ/qyDHmEaaVMGYso4PBIKxv5kRfQjpDMgj09cMsGGjgGnK6/BiuW2aqDVvLU0ar
6AfBfhwMVDdFBBngtg1akV+pY+kYDn7Jt4MGdwGtPt+JLHj9OBpt00SaW5y1cCOg
tawkpZzVH5pV9iet4kiwAlxZYUKAgfpBLwwDBZy5dJ0SmzVm33KgpqApyXuI4qFF
7qXFcM1X3c3S4LBnnUmXd81QSzXf5bzGaRuR8VOjlaTLwp1rLF4L5Cs6Od+oD3SA
SVObQgLQ8cIe60C2K8UhFCyxbQUOnrY+doY6NISs3BS3JQzCBbpd32pJ9owxZzSE
HmR01BDcFENTqRIoIZi+Ohcm/saL+xbQ4HXcO92Npgrr4tI32Y8m+uyLD+FuDU29
POB6NboHvx+iBT1I8QaSPihtmtHUJChYnZZIg/38WkVqxe/5egkNpxrXgocAsEFt
I/QwFICx7QtcGLYnBBzHbnlfihSBawxWpWgH0tWkhzxxAM/v2Fg9cjKO9MlOEvQM
lWxD7n+NeENcplkzdCkT8vQ5ZkYyKxzw089gD6wk51oUrWTSN61owlf5sWWcSlXL
t2ugSZVayldEZivdnsRI307VYvhpupYJ/EqZVRyyQ8Z6XI3h5bDo/0CwHpeiJ6/S
JBNdY0jnbZt5MNZL7kFYJ45YUfc5IOf43k/GBteY6DVQZoCR+4DbcsRLOgNUDiPU
cYi4ZRnfrSjAphqMrjZdsjPCIYAvpN1vNzUG09G+qrXEYfdZr0amhCZ5lMQMkt64
iG33A3ltYdWLHVl2yHBwEtwA64YK/xr/eVLitzuuNdPDPiaVUdWhVBQAh8QHu7P9
azQmpCasUen3R8erYuetUFNdcq4mwF7efAAq5eGJyHNLs3YO1y3XAvx21w6/9T8u
oPvbI2ikEQuSy3+Y9gyeO2K7C/9r+23gmaHsb7nNK5O3Jg/6h1XNRGhNBYaT+YMB
NI0BRRN+zbITOfqKC+4Y6fO+q6MNWa9QNk69/ZjxppzUnDVikiwv/vRQAkdmj1+D
z45MeVyktjV0wX2M0Z7yUgGsA6vRWjXjaD9URXZUd9QWAYzm5NQGCfqSRtaOYcf6
SzKeAwVPIHYBWTjkPJEHsUCbt3s4qFmG2s9LdLxzwZ57jbrHFZt7hw0LuMiDMk8P
WL2PtODkPic6qwD+x2J1Et5+fgMOJseDhIe77fvjVgwo1QkXhVG+m8Vy0u/Yvxzs
ujcJuxxWlNgutnh/PNi2Q1HRpCOhno/zDOC4MS1JI2WekNrEcndnLC+6sKoL8JZb
s0XxpLqkiUHI4WLUriYi/suqLYfoOa75F4dJu/VEfmSdvOs5vZ7atz+Z3orlGfyb
YpElX7DG8nSXsm8etoXruRkdkx25Z3YV7ONz5QSdtSF18Q0t5jSHrrqYLZUCWXTR
ZaseZjqyvt9KBUi1TFfeEpT+Z+kEuCyBWV0oUyDvJmFxrMmWgW62xxyxPDkhwZDN
9SbO2F0dE8GHbHgCoZ6LqoeP+pVlQwFIE1oulR96827LVL5HXLCK5z0g9Z0Ea85X
kMExElADMbm9PSvEClIkzuV8/H6X5CV+Wh83FjhuNs5p6tRFZ0hr/SoOBIPQK21z
uq1TPpIl3xSFgkDAKl0KnWByn+IktKwRic8cMQfyzoHgIiNkPTxvThpWAhk8CInK
1J9JHBCMegp7JEy+TzI86q44x1px//FJ55x7G7FlR+pXBIc/2joTpkdH9X5IfviI
5Z6R/ousv5TaZ7ZdNhRVD19AOfBXY2bHvH5En+jC8xfkVB0PP2I9OJ+O2I0iKA1l
V5wO29zA2/WeIiZ8RyQut02LiaVGZ9vt6StJlL2kZBi5iRFpxoONKuSDDLlmoMtW
lMS6tPIKYXy9KZRSBEwFOp8+2DXrzmNkJTaZC8Z68Q9mHxJJuaPOzAHhxclLgcW0
CNAEnQB2heHZFKouUyHxOevs5fEVO8AmWAkduAsldt0DstyB7R7RufzV1ByuEciD
g/mLTEDK+xTmA9D7hOzh1QjmoU/HpCHyApTw9D6YJezNwwC1s/vqqWZZGJ/1UYU3
lj0cX4HWnkTq8IFjaLTrAsrUPKbwjLF14OYm365Fh8bfnEd3VZZOfCqfrsgDLOUQ
ykLLXXE8gkydovb4E2LSevCDvpy7wdHEQkUnkEoQdzW8CkRYCF/GAoryOK2YUVRA
no2mlRCuAu5Z8XPr7gTrHJBQexR+9lPo3+q2mtV14YnWn525PaqLI+U4SBJZWVO3
NIQdQt5XoRiNBGzDWGNSXKGZbtZvkJ0zRoNhNXVXOKhHaX/wwF5r+QPqzqv08fXf
OirEC4TAG/cfqHtahohx3wU9E8ORAB7Sxhfqdd7gW1L3G0rUQYg3fzMQSkQKxK5r
63X72yZboeA/mv9k/M96HAF5jXJhXJdZuEz63TKEzKU0Ij6uTwmxVCisn8RxsQ3k
ZpIfVptbSXoFa6NCsGiAR4IXNOWwICxBQQcHxZOTnuhUhvcdjjcJRPDYNCiCjYms
oXu1OEFy7YPPeEyICGwV0v8uwMgExOPQsS/43VArCFaSHGwkb2/YgltPTp44XLo8
cp6VEKtw5xYYIyuaWD4Efm0a01UFz0N9CINkFoutwE11Xun4Jym+uyi7w6jxrWsP
FivG6u+o+qK0Lq0JwNKXxF3akuO7j7U1IPyPR5JkvuMXxh7jBTq/8l0qsDWfnXSS
dG7NF+MPWKWWw8fESsN+4p6/jPK4F0MEL8YmnXGAiUbg8kABC26Y1y7+Rco0jAEd
eRaSazCjTHuqUM6iTWlsLj9gSpw8WqO8qyT2sgPuLFiqFqRvItkCLO5Wa8AJ2Mwj
Id97UbNOybLJ+Jjtl5W8uICLz1VbQXOQsr2Sl3PbzJdceTUl76n6mo0ofACV9GXL
90wKIL1x+eRI97TVIv8T6OlU2APLU1fr/qULZp/fdsKthHYXvaprODs2GYyklGcj
ZhJsNFwZM9pms8UERGzdHIBwrZdtaGYGT+JFOzhdnPP2WgAH6+0xgNtZanS+V10X
2le0jDLKgY8UbCq90hOeBnnzn+rEAQygBO/9z3N9+iS5irkkb0ljiM6K19NnnvY7
wsv653YR8Kxr4/tfv6aOVZGz4JtEw/TSBItrCYXYI44Ye8RfaKnwWotokQZIDUQE
LTMiMC13HSfmlXreLp5s8O+GcOr4c8cbmyiMZkF3sFzvki1CB7iZ1lblB2KhIOmW
LOT7eW/tLWCvR+6ovC5WWvVdDmjuZmBQXA8+3gAprTUCWIwFloR3XXgJCZCOHH4f
BDcQKkKYIwwWFSacl9poTlR3oylwtd1Sud8QcUGOAQPHxW8OlputD+r6v7/uP8b2
G7RRsg1lBo+YtRVUIlfN8+EK71Bdm7OBkvWe4EM6+qii7XUkmiFiEaY9xrsLZYxq
8ayWHH5KZ0gz4f3TgBEQxo78EzVrDuQi7k+19SFZgVFy0tLAuY4hRgm6JaOW2kkA
nLujkuOAHXDRyUYm80Ak5v2002bzbCViHyOXRu675vy25AqxKAJ16kiXACzW1zty
FaDxV9ZlHgNAAju3sT8iCtr8sxc7eexUSknOWku06M3wyvxdr/5NuvN0nO6vXzLt
vVxdniELl59NmtX9/+6bY/MPJRrVZPpHnub0xg8DmcCWa/tRp93+AW+alkz4TC/v
iv1AjjSkibMesvIQRSfecSH21jzlu4bIDp7Yv+taTowMKHQEvHs1bcXEX1QTKHKj
6RHUShR6722I7/u1IrH0+dUCrOu54e0smblBA4oLCITvmPggEyZDRkGGN5ZYpX8S
XasV5XdvPLyatrgwM4KNf3CDEt2JdQRuOjYkDjYDyXT1EJ/ydWUp3qbPTRt75BH9
4b43/+ASmLWF6SQpA+Edwv9VMEwL7TRlxvG5V+QGIbVMsWjsMUtdt4NV0ATQDu9J
XCUQgS6x1Jd5yphcyqBpB0ui0/8X4GtChC8ucD7qaeHXbQW6CF80wxnyGwNIs1tv
G56AyaXiXUcJNK5FpArACPsIkeXVoRAlq1lg1Ab9PNvcNTD7XcKU0xMPMaq7Eh6S
ChT5x1EnVeLzW4h1LylLHKokfE5xKI8N/zCtdmghH9aSb17/jOq9XLU0Jpi+iboM
YuceW/ttSwnp03zm4UKDUKbRMmbnqQvmGoJYfdr8g3Ut9TWLBkAs0aJCFoiheCp3
cHlghdp3Lvg28hBDSjtotkpuU7ZLzQONiLX1E4NLF0gYGoYdLyZFIO6fsRfBDt+N
MrC/TNc7C+pzYIhQsecW25bqBz37IXOkVlMIygei/gbjxwd66DOfiHJCsqZn/qPq
KUfgDzqmBQUkpL4pWM8sWq9ubVQRaNBdFlJdSbJx1eLyhw7n9glIkptxO6Eks+DD
p24c9ZQYV4mO++99RvBC+XAtz36wz+t+E4Mkj9rUdfX8TjoGHX1Awlko4MvL7bVq
0qZpeHbpFOL/PL779upewMgADae2SqO32vG33CppwrDCiPGrdCrCcX5atRGOynXC
vwg0aYJ/ptw3bUcixQL+z+XGj7MTUxaLrrmPdkxF8nMatfOAqlJw4U/v2IFhiNYN
qL/3HldGbo2KCmcqMLRSWBvK1ksGrd5SeYTrCNLjrImBncUmJ72hVf687gD4+4tn
EFoeuACTUWQb6Rtu+BXSTOy871jXXHw4Xe8mpuL8XXIetlfBYuRG8JdhyHAlqqBI
WBoz9feQwbpqHY+6mL4IzMrhsYASa5C+Frr8WEKOKdIOb9bfqWD3uzqniLVzK/Cf
0Q7yXeVEpJz9xubr4MMOan6yjxL3f/4FRNFC6x/JNpFlu+CD9yhGyLg6XQ2OZ8yB
DL04BwjBqxBxcqLUpakh6MZFExAo+GETnzSYZLlX56NPDSQnXAxYaqU4C/TPYPAH
pcCPueaRLiuip50M821ycBQgWZMTEKOwBlPKlpHK5mAwMGTBPUni6NrUoKieqCVo
MjuuDMtiAyldsz/6yVWy5yeT+0+Z/RPMz79TbRYEMmnOBbfDoaeKr++lUCSNaj4C
ymLOAWNBhfU7D0Z7X1AHHCpmCkfPeZZ1lxuwUf5DC4ajZSQ+1cCWFWXEGHX53ZJl
jAXOS2pv1a+YIOQtqCPAdDB/6sZqvZjt3SQSsf2B9+/u68trN8xuVyxrgPihp+Tz
QU8xiFV1OObk/gfGan+Wq4xZ3/YQkbLA5iRA9orHW/7hO9nxu01uYNAgidZp+Qez
e7opPtp+sryFR9adfDkJ2TVBcJPHz6VEpn3EP0S4xpAdw818OZMka+bF97yeIdGq
M7zsuI4l9/YqyU6UpYif/1pDSmLi2ogZ9xobg2ECtqUAnIdxmyqpLZIozYfoOOpW
XUJ97HMQtP6vuh15QnS0GOmHQiZP7dU3dP29IfZp4Jwhi76MRYnfkSLcPo1omv+v
QV0dMrCn+6bpwnqZNWJwGVuqBSQAwj0jWEToljwkcMwtIdMe0K+Jvn35EX/IutzY
t1/1J5fF6LdHq8m1315t3rQ5QSc91rv5xwwPwkWu9IgKGsNAinhGhZbmi8AGbV2e
r8cleRVvHj9L1pZodUImQ3Ca5gofWZwJUR+qe5/kuaxaf95sxqO3rDYrsBZwxWr8
ybZbGdA9iROh/6BDwxiqlnsvSMBOZXc/7w0V32oADFrOQ9xfXl6tC0WOBH2dNB3w
+DIP9AVmOnDewMq1eoMJco8vGnw2kfJ/Trha4YtwX0l1MCfYx1y+noCxFZT2OjTM
ObQzplbEYUIbUtPFLM5nX0ab+aOPGxJGCZqXxGb6rkJJa0QuJ+LIFxp3D79YCXIR
szJbGU95o0TQMQMFQpLGbPTzNXpRex2c9GajH/1dRr4/Y+UENuEW9l56UgSe+9NS
LNffhIhsOhjM6e2PDXpF7pzdLf5gl2zNr6p/FUms0xvBdJLBV+IwxPYjc2L73OQ7
Zn9cbn/mDVzEWdQxPG0Wyioke0/XIq6OsHaldEII+mIJxjVfFSMhMKV2Sxk9ufj8
TE4o3rfyjU4QT6cYSvXZer/X4/dS0ebDtzuhu/cO1FoAcZrYM1HC77Yjh32mqhHS
wbuK33ftg00J9TFGmpZn+ce3PBS9yYkqtKSiJLIH6KgDh5fS6x3j5KnbkRDGhJix
6FUP16xFxNY2fizVHXLPGizxI52VzxJzBFry52p1cswDSeriRjhCJiKoX/ACSGsp
7UZWAr5YIfxSIpfabtQ3t0LPM3du5jXNMd1Z/10h4tn98+dGNCdWhPOA66EOyGlF
jyOFeJHIQ+tcKcWA2WOIwGx9FuufzfAuFHfeNRXV96k7NPaarLDL2rikVP5vMR5l
jc2QcCmm81bCNl0DJwzTe+YDbPeSAAi3hwb64tmGqTUsBVONqLlhZ+abQHWPKAgZ
5+sy3qDdGfdE9bScyWGHob3YbLDHyQBeTmHVOT3cMWT5bqOUAcUmzmKuGKNn5Hp2
QYA8/0jhQdTirGM2ZPY88sioS9TtmIPPcgBTereQjaE2qTU2N4OJV6MDCZr98kwt
FmR8//OCdQep2dBaQUV/7z1KJ8YX2L6usXoy6kqcYYXy0uTTbF78BbddbUSSwt2C
OgKJte8NJr9SONXvrWZDaKJee5VpH63NFMiZT8gXmX2WXuu6B/1TgTdwQ2nvx8WP
FOSuwVd3oPbE3yHUmboJYhgcqr97sOwHom8zeQSUX3weN9PJTClRvuLqhAzJoBuM
F6L53d4z56FdlwDukdcGQIl1lF5zExBi+8mGTi/+BdOnae1Wg6KVj8FiyjuCfuyl
/zGoIk3X1ecr3BURxinN8G3sFvPn/MbWdlgZ05IZR9gsFx8/rpuy+flhO0NlTUEA
RSCBu4zqCtLLvNyeaWKuegwEp0QceZvGOCrtstoFlsiNHsIY4hUrK+J8llTq9f+1
RrLD9GeLdL3jqHAbQaBfa+rYbRjO5B3SzNA67y3x5dEMLeruGUfEA1RGldo/fCch
LNLXrvNRPDCHEAPO0LjucWW/ZNADqGQfA4+6EYaAJ9rreBEoGNARqgDEfryoBPyQ
djNhuWD0l4nM8IA3tWLgBPwFeAWKe730wOhppx3IxU/T943OZBCH8JtQzWZ/UnPN
G+uBRhosfGgeX9odXgjpQbG1DO/KmbW9GZeDji9Bbf+hRWQ3Qu1SSgsubl2NCb1G
gX5ehnOPXVtsZJ3l3dCGKRhU9sxFKjKwsQ2gynItv6p3mHTQJxMfPRYKW0wlJXqi
nmRS9DizigvINAlZeMofXfpUriWC8usszyz6OLm38B0MXkq7hinWII9X5eYX2AWQ
Zyia5som9b+g/EL71VRMYfYVXlz3s7/+07P7jOanxDr7DyOYTzXBMgxedGJ0CCzT
ytYx7IPKyBvu4VzVPVm8zJzs4yJ7hRe+KE1xg7H9jtAi6kAlJSix8G2Ni1/6xOkG
IEscEYLFEdPltAZfNMTooQui7yq3MSuoLym1tdwYcv2zceI9MNgPlwGF4QH/CyDG
I5RNlKltb8+s38pAxrMV7UmozCQfZ+ipR35PEm3PYtMARvBlXUi2/zxXpoADBrIc
kySDPHPAdsAFKz0ARJxX8RoMAajcVq3KWs2asg41tVYiY/NPDRJPE0awpBddWdi1
wUKeAY5kSoEV8/WKB2VPMc12BXUeQRIU++rxL7NUccXvJBa8JEaAMAjkiFvxvPmb
zpXLUg28d7o9HYJiOtz9RE8JG2w2MQqSI2oohDY4d7oUyVORywfOUsPo0N0RwYMr
t0S0ak2VV8W2rVCyEqkZ4tCE5cwjhZ7rKO/2dl18M1Uz7p0hTZMXEId8DgrzmpdG
HQZ7sbyUKqjPdebo2S4f9ND+M/mzs7qzrt1eWgJ4WB1CueM4Hf5xTmSOFwGAsBh7
9pFdX7nBOwNMbBbRmzWFHYffxMcDcEZr40kIilSd26d6iEGrKA8gWQnisTBjCGXC
raCEVUrexhjcMSLdLQJb57CV/hPMFAmORW3H6fRR4hswSa1l56gN/axvJkkZwBoz
gEh/9JyAMXNHYSBrVRfQTIX4i5NZIdVr9hvYa9WrNrwE1we2EPMVULm9mrYOuVJq
YWt39Zc7a8gCRb1X2pHN4lKOPwDKSpkI8Uevd5J2XH3uDTX7VIbzPs6g0H2FhBuA
ThXHfxoBCts6Vj+w4d/baVEBArJfnyf+mVLmf0fCBTEk7sk6+wZj3wQIH7W8jvuR
MNeD4vav18z/zBqvfQf14tLO1Y5wXChq4vMiRU4sknWASA9M8cznBfAseTAzz9dJ
zRt3JQ8cEuK4sty10wY0fZeSvxW7fb5fsBRZU68SDOayEyLtGfXI7ADGbxvSwt06
rRrD+RnCfvDsDeuuo6aYDAM2haXOfioOOwEIxQGKp3WjXh7VhA0sii/YKSlx8Ugx
TUYtxkAArxXYNt/C3ihkjCaGdOQWhopTac845OBy1k7ocXW8aWNJnqk7/gBuFdk0
jK7NPK9RDuusPGqsyFhRRzV4YLAO+W9pQKN1E6wGVC/V9GfOPW31rHLejK/ezlld
FE0SyunD3vnw+nj63xf1Som3OsznlN+3XvPKx3HOlkHzkYwIkxyvMR6QPGFKORZJ
ZTlGrAdyWmHafVLmhblAgqI8mnkt2p9dDMqIVbtvPOdiurpzPzgP4bokwOPhXWJL
/IZ/+tFZQhwL7Kgtgn2nY9S4KtXfNEptJD8BSNBmkLXyQGOcNFztbu6ooOBt4fmr
LQEgKNHYfe6JTjerkq5bxSQ+rdo49XL3s5U5PASPRLewXI3SFALJuEbKJZ5YtA1c
v+RJJjreei5stTsW8n4amOiBAlef+dUx3J0Uw7tuZ60txzne4viCoah0boS9DTqF
bfzDdT4sLwcpGVsiOI47t8g7YGDRjHKqF6qANVl49Yo7WDcaSVTfLKwwN3WTWhBC
E8E0gZOzNLuB7PLxwMGpziYC6Ir+jI2/zSWOqLgNSwfUwQL6XVhfC3lok4vCgAiv
ZsL0BJh5M/kWP3V4mKmBDam+Gn9DOsth1OrHn97vuSDILQkcT5DH+E50lcY0HK/N
IYFnTlMpPu1aMTb0zFvCIExSal4sFHVFutdQ1wAa0tQbynfn7dCxV7oF4DJHPZM1
67Ob6Zr53k4kTvCzAs6P+WBQdOrYrc1uIcCoZQwBzPcjCc8x0HFiCIafgyRksAeN
RDn7p2RTZrhep8NJRO5NUWTw5RQX1f/d7ETXk4Tjd8HPfGgkhl4QTYTwQz0oa5nV
DO5X++zmY08MDLSUZQ25GrN5hl9EtVXXrcmWfotmY1HJAX11YTjiAQxXVmI6N1qj
DzyIsiPPuVjBRDrF3lBCAX1Lb01FHtDe+S6MNc0wimo3AxRtn35KkDkpXek39ebK
1XuQo/hY9vPf44bI8uWBJYwZPxw+RpeyOyUL22SOTUkz5COJ4z8VHvxUrMJCN53/
ncrLkLNsGxRa7ttNybjfB1otNNId9J+CPEofmsJn5rHCQ8u9fSEnaAkasr4DTseI
tISU+47NppXb/3agxP7ZYZk2d/sq/QAqbMGwhFJSzkky6IzPgOIxf9Dhleruo8l7
tGQTWI3sLyTdmu7eErpmf2/6uBe6CqdtiOajA0DHhoXpldwJ0Ps4Dv5R89OkwTW+
QxxfZUykTMIWhWuvCUOgEDwSYrXPCYOcZr6jKfiHqrP0ySLvCo4YvyEgbuy38viF
CMtEjK6GqsRG6bP3tBFnCieLXYx4VPRH39IUXW+Dw0ZjWKh7mIvQqoBj0QyL6XL7
b3FNhkR9NaxCJugs9+Xul8efQWGT16box50xsGnZNbzBcB7bwnpJ328p+CriTflG
GWTI3F5cs8Ia8Jzg9r0jr1Ht8KjnY6zValOyjcbJYj0NaTgYexZp/TNuQALRkZsq
IRipMJ6uT8A9HboDo2u0VpGM5oklhzqytcGW6JtT5zp4IpL9PgduEkoPYi6PIYCq
99EVLRrFpSxrL+PgoYYhaa83g2lXTift0SE/gOb64biwXiFtQzGLhqp/tZEYwL2M
SctDhGRO1wGz1wPnMt1N2Fc/Y53Vx7lYUA3DoR8DM+PADkf2m0P9e1b1m9ap8Knp
x+lYYdmv8RR1RwWkFiattcNxfDskbMJsxkvggFL8Vdy6v4lPQSzAxwE5Hk/lpKeM
50Jev/yU0nNcnntP94FQIjws6ylGDJnMGKFSh41IQKlOYjqU/qpJag+JpwjwBoHY
EqJqA771W3YHH93hWbeg9buowRYoylr4Mx44BtZcBw22GQeJZj/4b46r1++Pj5lP
v9HCgYy2lwIj39BUUvXCTZAxVl6t7MK6HkspPYmcMFTFCkxyuZxYt+mfOVXRem6V
AbLjH2N0dJ4j1SuEz/OXsTk/S4rUvCRUTCqtpWKd+jhpR0dYedzMugS6BWyeQu1Y
oBxp8I/iNwJafe5G58Gg5tnseIo/ywLfNS5ntFf0OWlvCuh8ieNR7ru+L7/pu+ad
YvO5p4eFQb4fv8GW6prLYhxUwUUyK/4tofIvTfTB/Xm23NS7hx3/eQCvgBg1mxXR
IXqkRu8Kw8RLaylKzqDUMOM2yD6JWrCky+X1An3eucBC2SJP+cVdUsIKymDnCd7r
Wkv9MOcd7HwhW6qFav8WosrKuhBcnklgG3gmzj/MZUgvYJCrrC7Cu051SSDOZUOn
mvRjpfWYrADUY/X5u/fJofZhuAcDaYwqMy0532hn9ZfUCZPgl+mgFQBPWBOStHrp
yjHz3fgulEgU+qVLA0m5TsbfMMceCIitmDbNSwTs8UJplgfcYyhNoOCDL+IpIion
J1d0zw7lAUnO0CmPxeOFDgER3YB8C2wpe8vD0599sIjjNEwalLhtFUv2Zv0w8mDF
3ZNYD/YPldr5vFE0mU8PViWnNi4cWw1xR7YhcyAAaf7ruKEv5Zp6/OK2eKuFd+x1
2h5WUZPTVX2TCeICow6GJJfKE9gj+/Qp9u+02AkQs4WK/0i4l5i6hPe8MaaY6EKs
Z3SjypcZvFPUuifdxKD2a1n4XbANHE50TDdcXBTt/dOp96jqdl+XaXcI7Q8tSQMo
I1DidMW/RaminUg5uGf/4I40ZGcZBhZb9rFF4Sx+AjYKMJI2/LjYQt7AxC5tsy7z
+QpnDeT7e+1bQV1V0q2VPZbEWPclzFNb2V0RqhrAg9xachy9wTRa6hp5Z0IAs4k2
HCHrCY1OsL3XAYct4soi6Xh/HOtrXWXeFTzQWDyseX57FUxtyHIYnFc6IjNcTET2
5ZBsHeiNNyqgzcF8k6GfaAD1+RjOduG80mAr3JWehApvXbt4+skSi+GOplGXXBmi
Il5AwpniW1WQWD+OmVGB/ljfo2oua0Avebwy/A+5O+1AW6jqWltJ+lPGy1IQsDFM
0G13yZOs38MO0lT+KWrMiTEh20Mvciih9KInY7ELlh2MvvsTmPrZUSzCToXafA0A
/HeJ5be2BS9nbIoboNluA+Nc39fYfN9DuycwTVS99eWxaznecQRMuirKc/ECJpCg
E3xwzPxnyo60SSdJKA//no9AIZ8clVt/pHbA6PiKIEEzXpShCygkfgxZCVO1Qh/p
9dh14vTuZAZ+kCgc53ljuARb0SXXOGPrOgc8W1FXXziP3VJmLp6mj5hC9KUi/HWD
LV+o0gfjwpI5EAr/Sp3lqK666nPcREwsndIJeW/ZOpz6SCTOeuEfJtAAqsg5STs2
5w9k4N+tFHTiBQW7M1ieoew+wY0OF5/Ka1ZZbKCu/U0gJVHc3Zt3Tp7w+wc6m6Q5
1aCahBR5EeD4MGTQGun6MZ7yB2oOWWFen4Ma5Z6N5kwOdwea4DgHdmWSB8LlGvbd
gw4EK8UDFi5bPwzBZcwr0Svq+tfrs+olqK8Q3AeuFpOXgnn/OiuIVkDmXxUOSAKm
rW1Vms3M22tUbvtqQ3GxN1EkOMgJLnnXduXqFAAgbVCFBFVVAihLv6FZJHi8tHXd
9j5ajL9E6fr8EMG+syH2EDiPXzQt+KFn/vAMJX5JSeBJvh9vSibU+3q+DEakW84n
UQbqmHqzMlhhWfwuuXmG7NS/javPm4lr+ufC73N++WKoJuHuBeN2U0hc+z3CcjnI
jqjuZbGUUul2ZtxLheJHoXH/ipp20xOxYln/uaVHDGCrYMn59GF2+j+SKuhdm3wr
DO3MgWi55MlNU8aE+zXCTulcqWGnYvO31w1AsSWCrBqXepma2cz6KWvDIpLBP7ve
20eLUfRfgNXA1Tl2cQxSdkM2gPfMmFXiOG9nMOjUPjWS9s60WVOQ0FR1EPmFqleV
GBG4bsvc+W/Ukman3GKN93LHl0QteUgkzIXnQD6Tssn08b6w98DVVpueBSaaIh7q
x8ejlUHitAoIpseZ1EqdBUTEKAXCgV+ZPqNkeVZr01IBeEfOnyJEmFyW5954XVyI
QD8Sf/CWzrfqhZz1gqSSQFmU88KlpNQYI1kJKEV2nhQwlaNqTaOMwtkCJffQc2Xu
0kNWEXceF+G+uH9Wq1AB0Rdn0lB4toJhfHC62F6q6G6wP/QrI4qJs69JYeLokV1E
kCEMnIj74vqjpFr6aC7mw1mmns8Y2ZOtg2Gv6kITSu7RREerdrXq+TPy/sFKtnVE
vsfastEyLku7MY7mv0MdJKuOgxm047+xA1iBcL0xZHtA/zBjGtnO7J9Kjy0P51s9
HSUE2TCgUAd8+WwBUQrsZELNck8FGVEU+ZoxhMjWtGai0OnjYZXsjZOcG9tubwyO
Bwqdym9A83U+exhdeiwasPq8PMadkqiCtv2h93PEWWqITiriFsK6f6/hjd6eyli8
wRa2Se89FcWpJZEQT36heR24q8gdIdtU9qKK+OKU+qPjqru84hVXBMJBoLTk1O1n
tvyv5mWH7s7SIiK1Idw/AksUWWioZQRvxLLqAPqoh1eVxLhOa+jC5755NOSiBDXJ
Vb+2FHWCflbk9zzCFw4ZSNwDiHtYsKwRa7N5gOhczHF4M/9rsXenmlsvlyV4bT9s
2sfgG0sdUdbrVUAABOJRUz8q3Nn7eMiuLNfPMR9Qfx4c1TVOeE4Z4Ln2YuySVXlw
VXlwfX6K9yB2UkWwrOmHXI5nvpUiM1RMws/5EBXiyXeKWOutamPKokvTicM27i4r
pseLX8cdg48Goh/DJTwTSP2mpgj7OUJwmoJeWMMj/EQUqOj30vXUnKzgR9qlGwLR
tk+yaGmF6FmXj8bX6Gcnjmu4Sede0ALWnyJADxV5rsW38xQZiy4qT4LnOKWSeKCe
C+4GOwvRQ/WaNIyjC44m69Qm0S/E5cYC6eQ9AZZDjOlcOdj7syXKHmE/zVfu+/Mh
oUUuTdhPxppS+EVdDjj3T2mpB3Zfi4Y7q8sLGavxUdIzKfx4Giqewfa8fnMWSBcI
IJNKrneBW78Wh8p0MJZQkoom+qDjvK/si55nV3cAKLnTR7qkzDqkVf3h2eP0XCJr
5YZAhpdT67Hc6Vi9IrlBgPteXeTgCZra8A8xksyqTvZlPL080rK5oDq9Wsz1EiWa
8XVlaAt+tKmDhRiMEFTKDnxUX0la9wAMCjVOOIsi+qj/DVXgZHKEnjzmSidGnfye
QxlYHIOHOuOGwUvUebhM/bYEFrAq6H5Zd18ImQKpaxwbJOOe2Fu7VVzeWRhuhOpo
5bwmhVfy6E+Y5PiParNxXb4/atfcu5WZpi0Sq+TPKIqcQZ3TcIjbOqfteeoEL3aa
9loM5Z6FeIpKHCfgqMoUn1ua+3F4R5SQJXs+Ob3Ao4pAZ1CxVFFs4ctGD/vING9P
CcKjHW4n0zMc/H3mEANS5ps4J1hf53tvpwxQqZ+yuajjc/0X+q4s206ASEt5plGo
RhdWlh9cajizbZDjTydwiD/kv4IWMgAHr+n2uVoxRhCbfms72RAShOsise1VlZH5
oIPZw5LJEUAaYmEukIt9Hv4XyO5m+Uf6J/zYAnGOre88DU6I0OlPKATbFKD+CEQB
quKEnz0EhahJgmSV35Px5m15odtWb6SWfpJrwHzoBqg4tJD2YH199R6XuoUaxmZy
9Ffut9+4UFGDWj78RJeN+Vy85PMGp6inLBPxgcdrOvi4uMgUD5EbdFFbLTDgJ12I
K187TkC8ynXT7VuBqYkshVqo7EL2eSsE4U/zDwBV8ROUhnU54YEF+jfrLbQ7q20w
8wyTnZsYum21KTFd2zYcVtHgmEV5nLDwvDarJvopXSdgeItdTSZwYXqDv8UN+PCW
Bl1cBuII836ktnQX/gyNUBHEtHEFTMEiiqNXZi6IHPL0Q+cxK7opF02vbzIcqM63
Ax9a1+DR4LCUrerBOI3wVPdgSt5GDax3y19MVXvqU5OaD7DrSvLEIDoQd9wA9u1X
ESqjRB+MJkFcMakH+zyFJ4qmT/9K64B/0Gq0fYUYL7dpzI8VNJp39mG3ulDjvBdA
xULjYQyQEQpr5/Vl3PWTM+C5+euoo7sNomD0hleNR+4sMtVBIkKKeDO18gHQwAQF
py1LTZq0MGzdQ0wvUpVKE+fNogeZt/BPXheA7/hMDDgOPM4YCaMBtOUYYquRWNBU
d8stbJVtBtStGKda2KO0NfqK+972LyMj5oa37zdaRVYajtfgSHRuXE3SfDxLVvRd
HBqSDSiPHlmzKv/vikSfTFe9OGGIgiEz+r3ZvGH4zIa8Ys8vQ5c3dvWERDGvRwSX
mNJRTBjws3595+hvW6v+1JkIYAO2Uj+ynkoOfqzX7xDrphKUBDwZb7JPPIqStTXF
O8ICAmCKJ7iJgTp72u1kS3MUUJfTZatm1Xcfa3rTsdnLMKvuuqVAoxG0x6dd/4ry
Bwj2OSGLM4S9mMKkIuJ29XKAYrhudx+SEkCnze6f9cO+laPinYg8EiziXFsGzZuB
qOTAPEDCRuWHa6k1sCIpswusubeGXT7EjMsano76TkB+mZ3kPPHQe6a1E8FtMWQH
+7CUORgPyNPcD75fXp2N/C5TQS/M6l1/6jgtY/rQ72p7HvMkQ23uUW+UgiOOonzw
gZU1a1wk/AqPNZ5CNrGWXIHPrWZ5qI5gD8weedocAmjSAsSam1+KHB/LThpbDMhP
vWMNFR8FF8sqejoeMpyXbIKlVShdh5lJAMGNt08+5M5/Y5uV2JzFwF+mu0eLEOXn
gL0Uf+zo1sk4y7eN6xowjegyb8ORso+8Sx86LfRVZb3eq+7t+2zAvuMAaZo4DNJh
36NM7LCbUkkyOge43OEKdkZoK07+zDACMEQA+Cj8z7d/KaXoGtKDqeG2UeRZevu+
mqE9ELk1qrIuSVt1jiS/4Pj48/g4GQJwWSvbjH9JxuIMo9LfkTmdTl+HZbuj4I4A
KfxmG0bIqExMjoAM5GIF8aE++NUO1mB5cadOnqB2jRtJ0IPf0NkW6OzBkJ2kNfaD
ZCfGHb7r9lirZR2JpZA3DIFf+9F76T5zSWcEG9W8UW87g95fczc+rxwFwsFK9DhN
xYkcU+lKZKt9Q0x4KDZgnoBy/A51S693PHnqDrVJ5VATxPdFHZPm4bt8f1xt9xu5
Ij2hRqWTueA19MBh/NihmdAiZ3mWFxYcAxu8GlUskOvxfsSyuasfwxHjGnX0U1Oh
a0DWaivstXIegTECSQhCaWQF8mFEgWi05G1zpOVKBR+T711L2hqn4eNybcxu6KfN
Jn9/N3dnm6D02ESwh9rcTLUM7muba/xm/rxbWI2QgYSqEWsk2oKvvYUGX+EjJiqp
CkzI8WYX2rEynVfJDeIBt2QRLp/LOgB2+5uj4WyCxRdlg2QPuVsCmQFo79gKc1iu
bXJFb5va2/D/3N3jbdvgk74OhN2TtvW9VIUdFmqnWmSz927N2qvQGE7vaIcLIL2Y
3WkyzsArS/0Eozy1DatWFvJ9/fhW4in56gJrweOItrPZmlPCPb+iv9CUBA2ebx7I
RVd7P5skkVv1EBNob3LPWP4LYY4aIr6TWaMFiqtG6r0HlWrvY1+TaNnDWCm2MN5J
kkmiu2c6eO4pQ3JOy+tbslqWt+TSVVsQydh5FB8bXrwh11n6jV/OuBstlg32PHbP
HmMVaoTQqAymMjy52W+OzlP7nQJ6JH2r+HcRRsTesfL9h1GLJy3TY2hqIoUJ1Rri
NAGf4i0XQwfy2687Z4wd8EjQXHEotaXYlIiP88hbaELzdcMUfXtFuQsT2Gzfux+j
JYMI+/d965UVNv0DbNbiazj95La1YkWT7uIcFpkBZV9JbU/kGh0ZKbjRhl0Koknu
LbPz+exz4Oypz/C+7YlZA406HweZMWvmUjusqhqjoszv/I9r2gav4tVxMlwpqzMk
P8v9cxQQtrNlSZHnaEyQTPOhUHwWMzDTyaNkU2xzms7XGoEvzLee4kENZIPt2zYd
C7HBWwLCEnl74uoFe51n7lvBe8oP3TEYovblp23CJvnxXC0x45RLXG8rfSHCgV65
roKnEMRTbPc2TtZmtMmmZii4dcE4MynMrOItazH6O8RdP9jYlljjnBRNUZpHELxK
gYoHG5TTwWcC9YUwipL4Flrxj3uywA08eUYJSBzu5t19/UtMkI0IDRhhtH3jNcCu
MvJnI3JP/702ZUR6baT4u0KSijp8xhWkNX2hyvsgL8uZ1rFnWVgLrq0ALlorcx4c
d4+5KAqPwW7joYJJAtSemlq5xZkpmpa6cNfXrkqMn1tcuFZQLgCx9SaAzhtjTdzv
xhHhDWw1qhvB+HOa0VDEDeSsoZJtrBHD/c9z9KbyHieyHjURLg91e81aCmB8YQGE
gfTvP5ynfdSJVI2a9K/5N3TLVpvYjPybVe4KlafveNwSFGLXMlkgxsOkIHWs1k84
jnIJqHIMiqIEXaRHSB3stACP7dxESIXPa0DGcdCVUoRhcCU9XXA32pIaCyZ/9C6G
0YX2NdFr6vvIecWhbN9YvYDZYtJwPlKVA0KozljDHazepxjfaDaOTqqX3k2NX56M
CXV8VGmB+lnq1fP/nenuVfeZcyVRWqgiMvFImQ18RkU6MekuoSpmK0meURopGrXY
Z53LSdW+BPhO5JxaqBpeunQXuRhnOGXqy5b767vGnMlKm/PrWOXD2Mw8pcSVGYfB
+FpKeMdWKN0U4FM75GtCUrLf51bqbXnXTseZxt/pB/en0kvV6GJ8ICtlpSOSC5oh
vp1xcUEpGZVc0tjj4MK0VTeI1vTwfRgtEKpwG+YL3R5iMvHutQ06RbMSkoKiD0hw
l8hGaYuKocs1fd3bdUh/yWgYt74bRZIph5QUl7yyF+uwgVAqqwTY8aAqRA8FXHDc
yMEY+M35T3uZTN5DoGcmoSdmnNp9CccVCyEdghmW2uD4CFol7ZwoP4rXs7LlXPzJ
G2t0B58yzeYo9gFmSiy8UDM9eCNQeiIdlIASC+Ybt7bRy6KiW9FVkjYQUoMi1R35
6jEfCkdqpjMS1+wqW/rNYjO4W8ughurRB6ael5PZLTEFrlMHEfZMM183e/06napS
l6UbjCVxo/fhAkyf/b0NPXZJsZETPOwsTvcXa/EJZN4xDahBtEa2TtwqaQ2j7soV
O+yezYYZT5q9hdZz8xNyhj8oFtLSt3iKMiDQkc446ihfSwXvAAXVdwCrUz+dplZ9
h7oO/54MkYAizM7zb4CidRP7KLE7SKAwLX4SMYyIKRp830Xs+ROSLEbR/DxmJFr4
YtwJx78xBXo2NSdKHYDqVVQ7ARo9SNV/Kne56WCbCt5p6tdxSm0ArDhXaOlAJJz0
BrP63AiD6taJIpdeBFidnsfIlmENV2pV8LX8bBQpFewsNXT3K7zcuUlI/ks+m3NR
Ne0HJGt0TxhX6qhC2OzIvHgBo4neifWs09SLDXcYtUqLVWamm+gruT5V23DBSYFm
254oI7AvdkCpn32y14a+dHbvUk8CnNqA27dQd7bEOAC5Lu5JwBd0vF2ePu9KSphA
yJXETlCnou+3va7ZuChnIMo8Khny2sp9ykJd9vPDK+TCZezRnJbz1OVxHtV0pUB8
N1OsUT331cAmIsPf5gmME640ayJ+z6vv4bnM0OLLkM/P3N1fIAa5woJWSpx/IaAg
ueQ2ctac8jsfnndKrfi1LaMHA0+IS8+FHs4r1WnS7YGWTyAPlvh54v1V7kari5ka
mpWWdoi4K42yzpfwezbSgWtpj+FAlbb0YoYquURMCXZh4zBE7M63tn9XzCnlBE+A
tMwwL8z3vh8HRLH3VoI5Mwcc+0Hco2Z89/OUZoh94X6jMlrrz6DPUisS4AqXIxN1
BTZjde/OV3EzHs0Rys//y0GWNUKlfcUHMUQ7z1sPhAvaPWztb6mjmkAHjuFaZnAS
xv1c4KXZQNVKqj+J3S1qItcuXladkBdJ2T1erir2Yw//pYwAvDGe7p3Kc0hIbtJE
7ntYLPMEkr6wA8grD0sp+GpuEIB525iwmpDQhaLfN0xrV5BbTkzD6cez5JYvpkTe
yTa2W0z6Or4DbnMvtvBjmKiCnaqj0jIeyrDtvzkX4/5iSQDY6Ko3zYIaT+vK+QTn
j3JD81Yp+MGOVbYPksHxcOkNC/NTsHr0EXsISsVePDbgcuX0yeqKfxBtjcuw40Dh
TTNvQXektAJQZH4ttShF3rU7EQAucHfnhTIPm9P6+pALnFaCnUmXK5FmnqRgqWLt
O3yYnEL9GOmPmWA+ZF7B4BA2rGtyvVmY10I+7wTj1Iu2Jm1giz+JFeFK9iR69oDq
bVPkxlLQrP15XOK82BVFZ12ZWSyy4nf8I4GLfT/h7OreU+CPR7sYMhqykI1xZR9l
qXpCCia8Y3aIKgrUyIzyBjxAvp2xRPF5/wXBIku1keele14uF9W2+JBCKu0NLuxF
NyBPzF338XbVfCtd4G8CBKE4CUOniuvx+UlMeiizn6CQeASgFBKiX5kWSToGMuer
1G2rV2JgnrYkAFWJcNF7ykJnzupPkMz+sGz8EY/iDMze3AJU4MnZ/crEba2r01Xj
xaY5JPEYpa4JWGqZWfxMrVee9sjpW9+vszd4VsvogzKq0aQLxLnXN4llYnV6rhzB
deK5IBsKMAkSs6SeRt31rc/yJ/DHxt1p73cfBZPlShNtFF2JWZfmb/84i39zBhS+
JLIegg6F4bvddMhuupV32c8CW43PD3Nj/i8J3T7KHBfFbz0BQ/XhWyyIkZ0SwSXl
takj/rkG6SGBzaCx1yEd0ohxfpLh+QnAxGX598KF16JzePsvo5wVUk/z6tOqo3Wl
Yaz4Eab0uNSf/ankhrFISHM3p8LY7B8hn9J41N7ztTZPKuJW1GSlDQy16s97AM6E
WBEw9UoCak0Z/uzip95QmXp+icef/TlOkOgEs5RDfz9p/Hl/Pvanw5dOl+s992Ui
KGGIF7+wjoRmlBWwm2l9SHkTUl4ub8jOD1X5IG3ka4jQi4WTCZfAQJGBPdIulgN8
dJI1pON+x7fEJCo7UuNRYZYI33+Npb1sc1CufSl6ntf3PEr6dMViVkm3oDu9MVZU
3Hu6hNlFQ1+1UEBe70rHj0Fju6jTlo0IYqwnSAMDACrWPx14f7qGVcIr1HlSWbhK
WfaAmAiDpa8axYhA5T8Sgef+0Y/agMPO9LwUV4Ww08saFvCoNPOgGU2NYW3shy3a
kdGCHJ13++e7rxUsIkQR3mrpglQCKrKxpG5iCfKLhE8ijbJF/9dganPb+l0gseWW
SylCAQsi/g2Q5HbqmomQI7SlbPpV7h5jlN0wEptfT6ffL8CxPWENYuNUT8+7DgES
OynVEIiDAX/dOW3EJeLQJCflb9Ti7ek7oyYvHrdKsy+/nmS7t4J81/qOl/e/SfF9
kD1SqSQW19v1/lJSTRg3Aum65zKfsl3WCayeSLGLjicTEdAXtwsqgD83CPYhF9U3
VF2A06ORVlAQouYzEdmrQChbbXJc4ywzF9x3IzO0xJQKMEuCHATkpNi9T5044ai0
9NjKvi9Gjv2npN/xLQwd17XUKksp9Ur78/QWPFp055MFMdf+buG20c1bSaXO9eVY
5nMyR1Tw5A5uSygL6fz9Y7tbiycD3XLoLBAQqFrTKwMc4JKe4zR1PcV1WaKrBkRv
aEmLjFQk3SEdC6Mja7MSMaR0/sBjV3hfldJoi9xoP+WY2S5z/0aGZP7INFo0rwpf
g9TxMuJA8IYkDSQM6WsP2493fEmmiP87e8L4eIb5rHMEFS3PqcD9KQTAE0fZlQaH
4kFota2dWlAtSZbdfhL2O3QaYrmJyiraBzFXLdacgi4efimFr64a0Sh2QEpko9+1
b1XLf8UMQ7+zKdnDiO6SwwYogxsd8dv6d1ZIj0pJpBjKXGHMmfyShjJhq1d+u/Ft
G+Ix6Pyr4ahGEMr/ngsmfA/LxjO+cE3mIhmQ/zhG35GGlGzkZYNfW8h1OoFs3v16
XB0auVt57ZokNDimJcqVQPuMSskaJSFWTloj5ZgM7doquqzjRHTTDzOHlSRVCqhC
CDZKfqwTvo/os6wmGXYClmxZJK1Mo2M/NSmfzk+BA8zYFC8HzkbzfgVZy7u2c3jO
vYREAhRBqj3imOnUR0grSQn/7RmLJOIaVPmXLLO+I9hWSRhtMb9BCvN1xhSkesbx
LdUmnU127PH6OljbiUFt8SSjgaBzyZKLzobV+0HY/8OpoiXp1K91mlCmi3FsTvJw
9rBFSzBcLg6JRRpnzYqZDPYLP1mIyZIVziw6ymRtEbDcg+nTqEF2s9Y+QiKSLdTX
0jBmA18euiLv98raS1E2PDg2sOvux1GGuRg9RqgDcFy08PFJ+5tRgYBXUL/F90/l
jVUBSTtuyZPe1ih6gN9ImPiQZ1Vd7kLbfzx9gtogxkJSLVjO7qMcc2PZ1/vN9ApT
0i6qSUF4yMdi+FfCWhK71kWrPWi4Mr9AMCjUESloJqYmcvHgMZ7S1zyNuVwfWvy2
dD8ncBJjKjiRXCfYE1ljMCEJTbur70R4O8SnzWro+9BEycouFqnXHsnwRSftdfbJ
lbsa+Sr2CUN5D5v2kJNU/hcTQrgUJaBvqIDM1WcDpFYbcmuVEjuZrDfMXs59leH5
QH7xxAo/X3NI7Ombkep2KcfpNEmFBra7bVwecw5rgrNqWNmKVcrbyl3oOG8jetGA
Ti55JZTxYGPU3REq7/95GfE/KmQM0qwr0xxBdsfSouYxa5MTySQJ59xtrpg7gh+G
ONe+KYWbciLBAnTTGPMC5CEOb9pUXEtXaJpi6LTwvUEyZSfulpk2w90Tg22ZudJ6
aq53n5oBkJ1a/2mMCnJn3uqDE3kWr8fn1D1Q8BnQqvhCwVp3kKmlmIeZJjonY1CS
kig4ORGHV5ykVK5U8/c0iZ2Uy4bMKSOXn4pdfSn8I+6qSzkXQIkZdbSfJICaZqRa
fs+9UgzAZLJHrhwEF77vCsKE705pRFeYnnu0jIRs/8t1N27itcXpMkuYMyv39Pxk
fEEuec7IT1UVG3PMSn23Jzk3mKQpwXtqk0FegGUdt3SrWF9Q8xO8SfkwJfRE51vV
Tu9NwW80UeMS/BqYxUQ+vSC+DuxJZ97dkGe2HL352RVEm2KyCM80yknUvRmewxXI
3Jr6pMQTohR5W37k3x1Tj5Lt4V6/H4/yK2jEVhMTTGHbIXfNGeLX8t/GNbT98iTh
HIN0NELB1/GNHMU0l8aBdHj1dtUZihVeelvjwMIw/JiFlRKTpLvwmRcEedeemHTA
Ih3I0/GvVoZdztWMDH9XoNetfzY9UHFkjQoPx1uBYA3kXMA15BqHqQIbmpLW2siX
owP/HZrcLVaIfZXG9r6kPR9SwRxyoJwysgDyhdT9IJqcOM6oq2PvtiyBMmQgdZv5
vo6Ufwcl9tn04cMEg6kCQRPY1gxycZRkEFmqPEyIEDwBJ02AkrSBG+L2Ps1oGTM/
5pU3vxdDU9VWZwU+E7b2N0Nl6Lrb4O5vXglDqyWl6xd3bt+EaTgdO7gMcDaQRTSo
b0jQgzbuLL5HKtyZDxGVd4+R6g5KUVodeTHXbONbbafUYLA8lek3pOP5M0YiyH8y
nxuLCU14wd1w/oxexFM1LV/BpivNX513nZq3AIaAh6gvgIe8a9FJKYzLDc8qEeVt
7Vsv5qvVXQ1W6wL4Mt2gtSw6TIypRfkD0oVrbS0DrfTkEm7JlEueaEtXSQ2SyMNM
JOIaNbBKqY63uWuVfxLRcx8ocfdVgp8p650sdkkDEpaErlNs0LTJIu5MwdTrXxHu
hJWAbmW9/4HRxI38JBwNAzuoQgq2nEQ6a+lrOf8mWCpOg+JiX2H4qNw2d9+Dt458
ge3ZYoBTgEecDmDePUDzaZj791sctdvOqwG+G0zQMWxifOcf20Sk3dMk0aXgI+yF
JrzBPIeUrobju5Stff29Io+315MXZtPKcB2CW9CrRrwff9JQ1bTsehE3p4XZMeh+
mYWQv2QdRlSYoEIx1fO+lspPtp4vxqeHcYdksFeBzNIO8NlgCbxSetrpxDYvBSZ1
YDTSNjaYCVQwYbc4h70Gjpvr1F6IZ//02mxX83Xz4t7a1XAeB1lU4YYzvUbh4hWH
oNYFzDubtXgf+2+n9nyfcYJ1QBn7VE4V/HsKAstjmYMbZ92hSbSow3depqzVGPxJ
jHxChXKXLXx8qgR8EflbKmCdEBqEnYE0On06IXnAVesR3nMiwMk274murwSFhfry
Er4YGjEm/3pdnIXoFqaQudA4SDLs1QcaKS89F/f5eYQlGofV3SR/VJ5OSm2Ymlgp
vNK+NEec6umEC3uHYYQwR3qPtQKbqps5vujGQ94iD8XBouYbaTLPYlGMsa1NouyE
YoXkSf5oyjkSYS/UM2/QC14HSefjGIua77rTU9h9zrzryTso1vDkJg/gV8B5/dZ4
gF2UVwh6vdsRXQtQBC31UuZpsfbxKia8e1W1lJsgAytcFBmyTWyBsJd5V7Y221dm
jtkyUsdXIf4aq8q0BFZiQS9gWaWb4iBvQIOBvGPkm0/n8LoJOoipGVQdRjkWWq6J
NTJ/cuTbG06IHG9CXYQXVLah3SdkuVfYk5NFevEN0vxTBZVS+fJhPJJKjopXfeJW
F9zrUxSfzfXlLa1RsWeOgiKNmTD1xyxUwBRyiR9/WfYYVQrZrhz1oRTdwfYbWTOA
aXO2XOMD4u3l/xMayr0iQzLj9K9O+Kf/tqbVTib9sd3n7DU2xUYdIINOV5yJzLu1
4WmtT5iRyoepStWghZ6GyEvcSFtvM+fQ0K361FFciTi8cbt46yomxFmM5VxMXfT5
JnNhkh8+t5/trqDjKm1H0n+anmGtzjmx7ir4N/h9PSGvrqs3LUCzADhMxkVoLK2a
t1Xz8Pqn8UBptmZMCXHEDV4AuUoqYILO/6oP365h7hlt7f2pg25AYTbdBQCB8xsO
F2U5rjCwOxO/lEUcl4w4B+TaJ/1DMKsRUdKyI2eblzF0XA1DGiRL/Pzc7R/nsOgR
gi70EMKTkFdKFq+py1E4mXLcBE91ez1pcnmWAzFV/wv5WYhD/LkomWOt49qUwQLS
jy+MXcTEvuN05WlAh3y02CUzaZftCk1Bb7WHt6Do6zn8c6qSQQYqMHcy/pqwGtF2
TJp6OpuDmI4OdvQ0nlYsH0P38eNKN2wwCHY6t3oW7zvMysk0H9z3M/kTEA9aywPk
rVyXPfM61FfR0WdWbnF6e65IdIjGWGRtb/mpGvoMiVK5eZl8sOTnv3KbIC9VPxtK
eU9/yTq054V7bHsQs4JxzA5cn4PrEfKRx7qJZ/Yk+Ge0sLyx1+iqh9CoFxWCqsfo
XCE2olokKtbAO/Eo0YZVy9HFLt/97GfnRYMVwQg0h0hAZ/zuIgUq1V2Tg/Vzx4YV
as4LIILygn8IngNlxnoTf1V56jLERFLuNPrhfOPWLDNDvV5LkIsFu97JjINg0cwi
4AnlIbBgbvKGEh8+genqzsqLYKDVO66+/qEIWhRsD6Wm9zFPOd3zvdIdGGQI7gL5
D4Lfbp3+mM1Is0rmH5Wc2pDXpsS+4/gN1H6fQ+/EXgk42XlSqaMZ6gIiuYmPogbV
zyoiWNw1vI9TuPVNBKMSDm7DgeQS7LzVCnu9gH0OrFGVh2qY/vatsz+X1RbUwdXT
zIORiwjLTSWt16Jq/MatwXXz4GmshToijMsQcppcg/elwpPC9oTlVS9Xxtw+yaf8
f9+WTJq2bdq8FLCsHuk5ppbSLLX5kCJJMlxqoYY87/ViegrJLhleKFePN1bjv9XK
VaFK/tZNx1G+6oF+MsX1xT5x2Z7hvr2eYR/1w5K3T2ED2heXDb2sb2PHbj2s0lBE
L3fTiH8cmMX3c4E+FE16ac8ZvUcmjD5lLQ4ejSqACEl1I7fwkLoVSiT4FiOXxDvm
2c/ApsSJRqvuwu2KDadR+uZkGLfUvdqNN8uNo0etarsXo1xbc85K5xzLls/AVJ+R
aYyKd8d95A3CvmhMNjQyYcdZGtbaeQQ6JEhuoKBhWVdAx+J1VE6s5qdiEUksxExP
S6wZYRVGV54P9KjLAMebaKk1NexPevjHk1EgdSDsQwnESnxyOsyMSDw7d6xGVEe9
BB0oNOkIwJs7nZxpvaHIa3IUR99rHz7/PHO4n3LU5chOG8o54QHwMTc870Jftk/b
GoeDROmiJXQ+YevmW7GHnOZ5IVY9kSxoRzUkjlF9PPKgPAmtza0RelKWuiYE0uQT
YUBqujjHnyPypBWa+oL0m66J+ZY6t4e3JXEwfIj+cgdm9NJ6Etz8sLiNW/rNGs/M
UOy3CnlctdZGbDrnyXNgrxSb6e/uLHd7J9szYLXd75cJpqaKESM8nPoqCfy9dxig
9uTjBpr+KhS6oTuJ5r5ZUEsCeEVX7GlnBLbF9QfUBSlCVPr72GT67dQO1qFPVJY7
XNGJMg5TUyvicxOkDJ8hvt2NjSthXqFceT9XiRxRdS6rL2EMb6dsEegTWcvKSSEd
TRLjBAYFNJE+w5p5MfMKil8MbeO2tW9Ypr6KIQBlRWXYrPgDv9P1/3hH8MsVIXPL
iXdDMRjWs8mwOM0kCqkZ3r7Krag3//POELGPR5NbHbTeUY1HFq4mRp7y+leonCvi
S8zJZjxml4BRK9LI5znPCtuWAapBOqttFkxfqYihmRQfriBNFEGoxaQ4LepxKtw3
q6E58WHXSOJdOtFjRJSeub/543U53rv7pTaJbhU8ljulo/ByViN3UUgIZ/LpN+Ss
t9EIYqpFrdeE9gyBHTJoUAfxyfRVJEq5LBMXPnUF0HHDik9C3IMfOzQQQcjScRk/
9Zc6D0JHUoM1gm3BSNkGrmocnKQgPOHlM0Qi3U/qlQrblp+Flv1UQT9Df4H1ffs2
2NTkOJDnt0HYnAP+deOz3LVFAhvK45Re9Lsy2wcIUrSQG6Qgpimv9dqdEjwBRVrF
XvG70b69QllC8Zl4iJbSXyX9U1lFDv6f/YKquWxKqke8IZK5pOmTNwQiTVj4vpLc
fAPwg1/N7Kld9u1KCHlJwfuA6aU/zmYw/hDjXywbolDUnk5fHIOuEn02LOtYdHyS
8DofdYf+VFmqy8L1aReegyJoRCvcDQl7wypL2lQczA6LW8vwJfWfOLPU2J7PrzLh
VCJDQZ+wA3yWCKDID/tkjQMzohflb/Di4sRGWVzYjVP7zSyAniRnBEaWzvR1wk7X
CO2mNQxdCgXmybVWR6X0lY93uxfk96aTxNbPl9+gNzgAMysfOfuDlHl5fMFVj/bj
LZlix0E3O4XAUu2TvthyDjTFUJo60Nyd9INZ6uV58IpWaC88VHLCDJNfeZROGAA6
eZPi4UxS+Lc0B9pVml2/fszmsoDtRVM3tPj0zWUm5t25qYhU/4NFiPmt7UeOmW2O
c61D3UeI0GFn6iDAEhjuPJFxE47SLibIWvgpNekPEGhyHvLK63EU087JWCdnrRm9
KZ/Dn5WJCdCVmg8bRR+oB7ek356xUfvMOWLTovX4Sht6/kf6QUNI7ure3G2KOIYa
jYihRCfNzv9jwk0FN8MYbs27ZQ/dzmlkobx4TyrBl39EJx7S155OmRpQV/wKqnMR
u7Saxg502tOUnAo+yKyuSiQZWbCzHWlxwTwsZo0uS2Z+DKyk5BYfjd+MEMY70KQN
ivIarMW2i/0JjtDYlQAAETOU0DjfX6gAzTX5OzFy7vQ2Mt3BTXcl2U6UH0GEbesS
WjWQd5zdD0ADQAKRe+FYzhzIEeVOCFpdTKp1P9t9OyR5vzRLdy9fkqaCdVXlYQsO
ReifSYwBoeYlrmztXwS92Jdp3g7L1MJQhjY/goN8kAWTChB3LRCKvVGl2XeauqjG
Qb8SDXEdL5DhI0Kqdb90r1bVSMJE/zb2FasvbAHISz/wt5aTS3orWylPPg0jC/y6
A6XbPkSZFr8pOcFkOpZR6U7RdG9doRHV6CCcIOgeSXhaty6YqAcv8tINxuTkeX6n
o0NTNravafVnJPTjKBWR5CTZ7qjTFHXup43uEOVjFIvzp4jdkxxUAatfC9Sjgn2+
sqcv6ai5eVY1msVLlzoK7V5nKc8Lp+QTcuWGk9F9dP3n5qidMAGHPLCMB12M7HcH
9nuu1WoRCUSoVV+kdrKkP3NcUU1FT307Xbu5M2Rdiw+L4Q8IV0MereUY70PZWNrT
e3BdZOqNv3zHX//Jx0AsZf51ODJhUgNGY2C8m5QU8KXg/fWOGbLPy5k8nRa6cWLe
eJzuHJNTORnFMOYmb/lEaMaG5C7vOKGGZq5/Drf3FRFJBGO9j+5GRTBcp1OUXxDz
ubBRfsNIyF9TjOyc2UmlGWfgfAXFARw1XNYv2VlhOa3AUhmJBWT1WU7v1EzJDAvC
lutqBo3kurYtt1R20/uWBm+glPYdZrDoEvIBetPCzRTJhmlYfo0IUKWMwdR8gfJo
KA2IUWDrTByWPhpy0Xu/8uTPZWw5jT/eGZTy6yc4uyFOMQnbNnc7k85NIIbQhn2O
R9t1FCP753jU+wAB2G3s+vXu6RVc8EcUpFcJTxmeHUUvodTn1Ty8ORs4keT0feWW
NNf6+DrpoVTBpwWEmtggJBjRzJ8ydmOlT/Y9Yz++dVYv24q7sP5vXY/TNjtNqkvl
Ik4OFQBmP3Vn24jNqN8CtwWn1fmn4mEmB4GUl5PWkxc5ZHRYEaDKV872IRgoQPoX
rnz4NGLRuU7yvJnhoHuJ/hIoujfEiPmCLsArEa2KEBtAry4rsEFdBnGqwGZ9EmHY
fEiarJDhbaRUx+/2kuYUJEUw+I2FmQDXWIAJjryRDeFxIuYjFlYoK0SFUB9afYRr
yU/nYor2S61VWn8qNs/mOB+yP8oDWDv4eR/jXmYCinmpNm2aw5VSvatgQomXfdjn
UUaomkBKM3Qcnf+k42nz+4usG8kGgFvSLyiwcMe7OqtMz8DIj30NmlOEq+g4Z9QL
8ahN2BF4W0Q460TcwMd3DIvBRaYCmhDeF6ORDnO0yENnzbtG5NY52dNb+Y9UNUpU
lpbJSgRHUbvudl4OM1aJhfdadM5BwRZS+xi1e4oTLyRvNoVFzPWm1tcdNrwTE3YM
YVDpXymvwJEbRZ1+wKZHxrjUwx2xyW4Kd0+WFiVDVKqfBgV742MZyhxVzVyahjj+
qROTMyUWEecjaRGR1uToBX4CUX2KVwN4bXQL1uHfGaPr7VF2zHoy+/K03XKFDkmE
Nt7dmaicccxznz7SO+vzc1v9IcMF5YjZAj1HfDlb7+tU4eG/bcz3J5rHGb3QU5Ae
CT37QjSDPIZOjOzTB4m8JaZYBM6d5SfVX116RZkXGi57AAq6IelKW1SfSgJk3pt+
Y/cp2ww/LS4sNNKkowRVprk0ndz5erPpNQ28pXRUX3p0mp1GYsXzwgZkNuELXoLt
L0pID5R1ALnpqP8tZj8c7GlKBJ5IvOBoV17/BC2it944vCvyfz4iolKMoZgB3Wlk
Q9ul7L/a9/dhBxaj1lEXSR0uAM2No4st1zcwVZsdGIW9nYhTCRlGuiSpY7Wu9cRB
cAJBYbsRCo8XaHwB0van+8sVhA3Yfhz8DDLPxD4vijca/xfAdjSLKt+9qpaExnFE
tWDXu1FFVgsQ/xP67WYvNJQqHnTPEkIthf1NXkr1X059Uu0NoTRHhKxwsDE1/Pct
tSJBOOSWeZf8GbXAhYOaqsH0ASt5JIocuYbImAqNjfixfncVBYrXBFMepmtEmnn6
nVtFvmxBro5I68ZPaoMmqfCiR7myQ6qL3NVr34oAj4NLjvjOJp/4KQWhK6bhGD7j
GH3J4fLVIhBh5onXp4WX5YfJ412hVq5XOXd6vvuXjdJn9jQYbCG2etdSCyQwC/rl
z5/gif7/hhVgRhnLvv9VlAOvtcsO16y5zV7eY1w14Y8LMXx2ZH2B4rMFYXg9RWGH
nMipkA/2NbztyuVxwCqRZGJnWZjpF5Ja/EsVjPoRwf9PxhXG32K8aj+1I6AYtjqJ
vw7YifwEAvgAPa2K2sqTd8/3jHhLqZ7hbLT7p5/t4/BODjoQ+ZiJHIZ8IoZuc/o3
DrFvfUH3u6148TQkDiHHSf4eHXhBMPFXKTSMuo2nZRZgFrXwzodmhc+LKzxlDmy2
QB8YAcEWv0CQi+HP5iroLFoaM/hKo6kQ4Roi8SWIRsBctYgEdK4IHIyh4MuxBn4u
0IHX8/paH7GB1wfOxsZDgU/3oqw55x29srk4dB08SjN9CRnUuKR3U70DKH4+p3s3
WXi6bAGS/7ug3lizA2wilfwuTYcWIaSUk2W/3NbCh9BzbxlCrYYjRrExMxLOp3s4
NNvmJFoAIvVt/bcAKnCmBKjfdyB/J11UDIokW8lA6ekMzIny6ickcBENm6IoAZyH
d/R1WPpHFcpfPFquivj9t1aIWjosSrHOJCVOWIS0uDe0l7t9RTMaupiLDoS6i5ey
38UQoelFa5yQXZawS6yOAOO/MJqD9rWYqeKxAqibd+aZG6LXHBT5aHumAkdeJQvJ
3SWaMAJOX5CWvpPNdhUOZOVc1I4ppcVq075qexW9rPafjPYGKx0aq/d2fUD+m7is
PK6DtufyTwFIPJVGaeR9VB2RYy3UmqahyCD0JfAxDr/Uq7vK2g3Ewc+47BZ8cRkb
XuJ9/k5fr07ZMbdZZBRavnrs72yiV+vsA57TyD3BqmXFFCYNuoLzFSDBsL46jfvJ
vOWS5cwVcUAJlMFTZC8sQ06xtbK1p321kM6ZxOdXAAhFqIpmsFXSqfmNiMMks+yB
yiqkZvJ/7TSeZ3HfkivmqGLw5wvt3LwZUz6sAgY66mYJ/JdyiCxFRWAGHOWcV4Cs
ciImKPjyp5u/lmlI/MuoC+pWr89ERCeDOLqMxM8/nJZvEN+jVMSradzsvZgDApoi
wQcuJV/Nut1GezeGorNhPdMnDUDUjyfhNMEBVJSD7j14Pd+pGEa04gZjLq5F602x
RBwJvz8rSUjfPcnokf0l+bm50vU/LOrOSRFEu64gFQPtjOXtnQ9uAnY0hOMncsNR
co7QJMQ3bpkA6yiPmSs/0DYbpm+diWoSdPFOtI8PbJSLANpRV6vqgETOta+NgdsZ
VBpOJw7D0+BBlBwLdwUsWARr+anddcTmjOsZMZnSSzE2C+SI7i0JBuKostYGsddi
tQWcKET2nN9dlYZzp+g7Rdp9dvMdQZuCffLoqovhbK/AEnfsv5xHjyiZkvB+Wwco
UQFpTblRs7ikduQsuw7J6aZhKyAF1Ad8/mU1Xvd9iRhogaOiiHB/H1b3xpmk9UY2
sMH81vcCZe5ZiFC3l3hP/rkLvMFQGcxm+nOt3VFvEu789CMrnnwPDFEvcjGOaxka
XDXrBfATCptiAfQgiXGRYnTQIHxE06sypB0rmiyV01Z4fJZyiRTZvCc82887DVum
6EljNrPbimizDgtZ9tUvdGCZuW1k/mqbBfoAP6zMC2LDuIG8xKEKXVNYGXRaBNSB
VtT90Esqln4heJWsVCtMUAERJBnLCdn4JueIB35SsbU8PgPQ5TCNHOfAmBqYX+zM
5Cy7UwATmsEgixi6HX/1pc8t0OjGf4JQ5zPFhzpdRIXABsukcjWJz0ilT6PiVt9n
nCUI+rtfWCes1gUc541Q7boyon/I4mWbkldMvB8ca0kq6fR7Aqli/X1QyaJFD/sj
1TbONjOvF6mTN5WMr2C884OpSUHUIkj9xlVaExMw/eslr0GlbJmTqvqwwNfne+iN
GLZdMnG1Gsjt5yxIGxYqa/zdRlhER7A5WITx7AknyIpHKxbIaYfMJuYc60FnTBTr
xpbrSYtl+hUBdbBJjGehTX1yPlYJnDF41BdZLOyzFy2rlM7yfImDJdWHUthu16Et
38p8PubiGBoGyQ316UFvwkpF/Ay9O/q/BHGeWNyPzTetfHgA76vyb4JR0ijggpZn
VJrSHGzl/Hx0R9rs24dmwKPAQP4Vcs+v3SwZnzq1fbBjNSW9J6ZiTSpUT+RF71zs
itABkkClxQ11+LgWbmQwQDd75n9evCroNLWqxguzw26eJL3JDszjwgmq58ONlp96
XILieRT+56CJOFYKwEk60Ix1NlfFbBiH08QSiiXkjBtP+iWXPK/JCpPiXTQKAZZs
BojWv8D0UtL2sNt+EPZhor+Wocj55pKMtTIS1cycJQwd3yYIMJDqrRavthnK828y
kY+CWP3uuQs2kqLtaMzM+IQ+NyJzniaSk2zL0nJ7phGcdBhaAm0/GAZpQrtUZ8pg
brIVheo0wwtzHkNwVXB4clcKGkuB56Lj4erA9EFkdD3lcSdQOPvHFxZtCAjMjjCl
/4Van4uRMzDYOGwwi5RRSdkem3f6JlPtDcpyx6WqwxvlXNXPQEOZd/BwdT9zeR2p
/p/b//oM/y0Js2KQVy5PWUqYCWWcr8gMb8OhcQDM+DlJKC7WqFzopfrXT0iXGxhp
q+TckSq9JmytUE3WTdMNHmSgJfGFpfx0uCsQPcYLkis1m1GJPgPU/GMMzVTwpppv
8GhUKRgqhn+WTAP7Wtnz2JNaX90PUWp/nEsHfH7/7zZjlWdNwBDkpK68NN751wca
HtFeHHRn4YUYFW1ZV2xfX/LPbhADnMJokY4eg8PYNm7nRkzWM1H1623Q6HFpu0e7
lU80loMrLVmecWxocT/v2YrY2xTQDj9cFCcfHqg/NbmjhdDgutmz8mPLnB/FRKh+
bCuzRyJY+FkDfZbQSiRIXGQeGU13lCqIn8R/xVzvybNDYmhaVv6yC5s5A1EG6WsL
iVUYhHCuNm4gvVZyfA8r6uRvBcg/G+9FxpGn0V84+Q6nAQMXMfq1kaM103z5WKVd
m1j2AwQxr9Bv6EOt3lyTQwAWquP0eZoGB7fGMcHi8UFxHlepzFPvz21VuRxmjo1p
uDXkn9m5jeZe5HdHlbpxTlXMEC1EksdsN4mPtJqQJrWVJOPeBAM6FP0R+uLTFN0p
uvHiq0FoMmX3XINlTqkd1E/qaicO26dvBq9hH7BBcZhIfYnObBqrhXYdFzJFXu9Z
bJAW2HiK5M4r2dvPjyzIpVYoIquFQgLlMW6XKARHoa6kcXHQXwLqX2uTKPFT17nr
CRG4son064H3SYb2HGudS6j2LH3wOCsJhqiWzfujvvPKJwagt1nHTtXYv1Uvxrq+
EsXBMWnSW7Xcn9e21gKXvoEb/99fyAHsymmSAGmzHbqmYWvpBU8ZfSzhLXLV2tQO
nMx73IHZqgURCO164JMsNBg2syGtmrrjp2vYLY/CQJGd41jPy2IlYuvzmERhv7K+
lp9DBbSDfqb6hjhRwgCSk//cKfjGkzX8qYLGFoqe43+f8U45my1RRNJLxi5/HtCO
xXsgdwLOeIQIE/OtU8Rgr42LsUS0q2f2pSUmIQ9XmrNb/WRlCqmKR4LqswgSzKsT
9El/DGUjWlpUX12D4dx6daRHKKYISwRO5Mod1IsqdA7PvUqtudRFdSU+AR0gMzmy
2dXbDaUgaMJrfKYnUBcPqmlG+6R7YcU8nSpusINaw3Gq4BcqFgBGz9RtHEHrebwm
vUSf1gjQ1IvG3MegC3IaWVE3pTI5S6RAmuuPHqcidKFgzwdlv8MVWkuAGIr2kiSy
CMyqciJLHuC2skZY6wksd20CylpSSZmvm6LbIJ1ypOHlsnITnPa8EMCHIHkyxkq/
71bDZFv1n7F56sU6XoLxgCFNq+GgcN6hOQF5yTZTIPC0rIltXdT3jn1eLCGmQydE
JHMNNzbF1iB1d46OtcARPxFgj6yW5N+CP6Pho0zV6hemWP5YUMy2k1Lk6Xnqq6U0
ZfTT1Uaoal0S/+MU8TdlFWOVvvf2NOabGOWWg9o9vWyLsISxnHhgkRS4KzttSAhq
0ZzCxRDOl8Q4qRU+nQuyrvnGAXMTqehmxW700M5qpoBhQKm8cSFT0WczKv4vvz1q
YSEk7i+zgsnKvAGHgxeudgxX0syWj2+WWmWORKpwB7Lmvd+xPc4mz9qLuysmeeJx
UrG1eV5806xBDPLRcY0zKilOzO6VzXU3um0UyinIvNDawqxX/qu1MYoRCKgCYCpz
9MaFnE7T8Uh+TxqM2kxRMhRX92LaNyvGPrbEfmGJyuIRRsgcRDDUjteJtTZWgOxj
Z+KTbIrze60LtblE6xhtRZ9D2AxzvYq+qQXEGM2bvXHAcZxS9hYEqIvbcXgo7kze
PmZymatBtL13F1oNEGiT+v65W6nUvKWLY+hay3UmI1k4NYhIfwmxd023xFPzDi05
Tc5qAyaLck0CYRIf8AsPTrns/V7z+ahACayvG6j7fZbwVwUnSmZjmS8v8sLCVu99
eYV+TdctkjG3bdmj1d/Z5sbn+S4SQsEk+9YF/+8VY+4RCGv9MSbryFfSlPASLxHj
XktQwYVeiKtkDnXBgOHXHJqbF0Ws42guV3OhNqCJG+w0YcYksvYEvblMzujSoss9
I/80HFMRTP2siYwRczhoYiOxBbAG0JgcCY8GRbdgXwcEoNL9E8oPou1mdk324doS
w8mM2nD2VNV998J36rlDpsD0dP3t8vaIKddm4zeNLpGgGLE6yTZmCIqwgy/dyiqt
F1AcxXSqUJRxvvPfeprLJTKNMcDh7QLxrfIzWAPW1t6D2tc0K/i1EyH2WilawIlv
HY1ps2Q5bwlY4QVORCo6vjxCDjal6BdgfzXHOwGNXYmEsti7Ugt7KyhOLx+kXiTL
2DC7FLRJ6VkzEVGFvcuSnuseicgBcW76px2wmxeq59Cz7cdgJELc/ZO/M7qFRE3x
JBTffJBqyAnXxuvwKhhFzyAxHYpMC53+qZLVu9yZ6rXi7hW2qdR3JKywUlkPz3nl
QkQ0Z0WZSH39viHqOt/wbpoLenV02TSXdZuLJBYXhxjrKTNf86LK3EjIcGWQ920T
BZKkAj7Cqnoxt+RRBnC5pxIcbsQA5PpjrPmEw5lGUhWjho5jnXUqyqmEFOArX5+E
Qq5ZYS2BAlkYvvCsaYQ9Fp7dRuXcr1QSzw3xno833SzkDklH6vt7wkwU0xqEjXQB
E7t0jYqnyJYHaMCVsG+G1K7IMdV8mJ5hRLnzxpzRC3tQbQ13r9DxPeH86dnUpYQd
JzyCGHdXw3dUP62PLjTJHc5Am7A7Zs4cPG5W6+xX36NFqPPElJVhF2KEMoAlqmOO
FCngSRHn/rZc6ojrAkAMd4+Ob3X9PGcaQ6KWsK+SUQmCBBU6zNCqRI4HzWBh0nRi
iXPpZzf8CK27FRqF93rQUIIMPEmlQRijQeQHBK/IMwyhOCVUQ+PejyMJ2ZfaVfVq
Qx1FMIXxg+eNsKn8qRmmL5VHH796NGX/La72C5HRslu+hWFn0cKrF+p7fY3VZAN6
4tcnEc3Q2hD0pENXd+1ZA56/bcGgtpqpm3hMx0iySG+gc+ZMbH20aMaAtcFEctA/
znHQ0/xR2gqTom6Z7gFKVh0hqTDLXwt1hUj/t3FCVGq8gcC8K2k5G27/Dj66nyFK
VgNokvhsabvEcGIonYyTXBbiFQ/iIKs2B6Lr6cWkYchsAFxoyvSK9EhW9bnpK1h3
dS29C5YB3xEElimFBOQmJ4H9I9+ViRPP3azWAbAXQvXa0RTAy1833QtVw037f/xj
HzbYgIsTqKA+doB9q44TBpsFZTzVWJGZuPSNj1JHTz3rpeCVOpYiyjg/HIkm5d+e
Hxzt6ZDUkYxVjpGtgSV7yxEDIrXH/hkFZ6V8sdO/rbYT96PO4+5Ey2Tej5tzBJ/K
yB0c9rkVxzCSm358lb7pelkUiNCz6a4QW/kS2IKRSBcQ3w6c/WThREKg8WUy+cvf
yxEM8zFwojZ87yTxvaxuGUSXKKVqNWLv++Hfv+9BWO/lBimKI4wA4snejwn2cw4f
BnJIh9pK3x7fz6vMIq1eTbKaubco1NwUrJoa7DhpMihrb8t4FuNAmbIQ95nggJjj
IUF05Tj+YI5A2hDCzDNyg5OPQYC8sgSkZxIB7FhOciFPs2FNjpzsZjautdHaH1L2
boz/8HqxMT8tGUyPtxzEGuTvEnE32fP5yQj0scsg5Y0O5l/YF244o/nzvyXIEn96
ert4RPDi5lIYJzA5ZmsRH7bPw08FIj//DBI4JLtl2PCVUHaK9a2xv7pSh7abb+p5
w/z/IBJUIGBUslxnaV8PYe+AAH0F1dEXfZagHe10dnbZXEbhvOy7ZNRgHLHoPa9a
YzfZoU8nahtwQ9Em538ZyZQifjk6rwiTo6jxiVdDu0N96FEGu2BbIPvqpjS9WjyF
BpRq+r6YA2Wim7/f5zkRzbIjduljznXz85eXoGh1okFQe3JU0BVUFtq4GOivhaNs
x9q18o6DkdXRQi42U8HzxXVkFfTB36nw+Bh+Cieq7lX/Te09QLBwNij2jdJ9ecPV
Y48QlitIhXgQbFUJbeSGb3kq1madUJB6djGjLulA2wl7PSMY5n6EHzKoWQUjRHo5
PJ2QHfjx487p3ukfHQYqJRQ89NRn5hQIai4/lZjKqCVTVF+cBXi5f9R11hAJxQro
RPECr29SbHsu54GS1G654IVNKRcd7o/oZdGivsYBFb7zSOMkJqi9kG4i7V4g+oFT
B1M8ObAdOtDgmzI0uHqrGYV2IadlUvBcc9qsLh8GROBms0PSiYAL3pl4Zo/jAhhi
66jKK1t5DOKB5lRWFvc9yHEL2JRSP9xrhL0Mv/vlTqkXjvC8/5ld+Xob+Jfczfuk
4tZS3Z2cCbxEkWxvnoPR1aZOEB/s00arJzjMHxFMeEhcdlRMZZgb21Yj0L4TP0U3
FeMXYeqHS2ngMRq/X7uNH/sOqxTCMvhqA3yKR2px1x3VBSz1dH3kwNjQ0VTbIvUb
Y8KlkWnWJaSdDRUAluhMq9c2k/fAWABCCIYTBFXDmp8onN8cYcSI2f2pcv0Iop1w
e3rw3WxVnYj1Gbr8mMyS7MdrNAbIKHB2a07wLMKpoT05qDl3wQI7GLnrooXAuFoX
BORIziEDo+CZwGKEcv/aQQfRUtplVLVuqbsSiky5j4hWLTRNgTnazuwBx97OWePY
MG7I4LvugwcHJEnY7BfHAGZfoC01hzyh5wJJf4xxD+9EzwbgOlzRDcFXdwWtytxa
pL4HpgIoHWKDQ7hmu8wk7BNdkQbrs0FsEO33HIa1nMsMTP6xKc3bdjVQgZal0yBA
rlLmVFmLQ3WH6a3WbevDnn153852hkQYflI9Zrz/FrDNoTbzgVi124LqSnAdfV2U
9F5/BRpsHSHMMpnDmD+ZIwXUs5XJ95J+shBbBKMtpsKI1Z3qvqiHq1HyMfFKxxM9
d7J6bfP1P+86TFgCAfgoTYSrx+cDkKTStIiD6R4G6eXSwkawTDqgJtGIv8S8NwGo
zMQpdySngRL9m3isyHYLNZFx07SVnUqvOW43ZTkaJFvRwwmgrAiwaAwHiQ4ZkIfm
ej1mtmgX4gELAWRG0xv+tzI9LZYvjuN7B5+IXAKUgY9KNxoCIO+aZhH59yKehNmZ
4XQMSn2dxeEPA2Pdef/T9p0Ekcc62dmQO3btdZptx63ovRRE66dql9Uvmnu5ZCj/
JgTXR28fRAYvDEbWFFAOMLMDXM+WEk8zenOKsYOymyKn/0qaIgNONdAMx0WjIVTp
/we+I02oHCKsgyPf4+1i0VywdCV6vLGCFShoTgIGfPVGszkOm0rVk8d2Nmla7Scv
PJVQhgZpx0sjRrybXERZPcLL7ZFO5U5ykvi8Z6RiKM4zSIBmoVsJH4W7EEoMJ/CM
bTcN6/9dLz5sDuHdGZPkz5/iIJCsg26lFZbKcBnIykJXn6oQoaMKfLDBkJULvky1
TM7bnqPa8aisv4XZ0DfWVU4fv1pXe9keXVqj0RLPRHfWnExd+RLZUp72p0Ea8zUF
VCd/Gff2JPqrTnukuNdVLlrdm1lLZntPLI3zHLoeEYDIymdEvjr8bzTNuSgbsDLv
F2BpnXZJ/BPltlZ5mk17nRtfJ8KlUaLDg1dLd9bITN3wh5fBK0bsfGbBaOSom/QN
Xf7CHITBZLU2tEhEaRCam0Ctoqi2+FyYiT9ZYf7RaHgGPO9jlOKioYKyuYNerpmN
lDqZE4mzkFlEmCsxW9k8Ntozzr4waInsw7KuWkoKSgrS10yq9sIcr7r22x+IXLG9
nc6Bh2bIKoUo3ouqwxsbef8PDV323jcIW4BmaFYe80VREMclCRGFbZOkiqWmNujQ
6PcWIPAzpcy+YHpjDQfcX4RRDP2sDH3eKCWFuHZaNx1IqUOQwvEK8+TAjCOcJwX6
ZzBR9HxSldyvvRrDapFkFMvKtqzqnNIJl2MhrmHEKp/aAIoEPxbnhFz1guuhtoQD
CK8/KiCYPsnpG5iYfzSs0wU/QFIv3XfonC3kbDF6TGh3x3DpUbq4JpgcRmg/Pv3Z
PNedVjvAXZTbkWOpAWz0zkwWNQvB2GjjznMrNxwvlVvh8rd70LNtQX5D9Hkh9hgr
A6kb9FnfF6ipZyLHqMaaTHPBNm9BJ2/cLUfKulMjlwzpaBl54RUBHb3WvHK4Oy31
atXy7ZuIdQZHDXp3fspbWsgrkmTkocK3wngrMnb38D7t71wzjsz2CtN3K+JjAI3O
zmvyKwmzIVXGHMSpPBMq5frF7EI/9lI2BOrGqqXjAfqtmrvvjRFN/yAHjIaJcrYL
aTG1a7oWI1aIpQGe139jTeTRFrYWADOg9FwAvMpLwoJzSG8YMMdx0p7/DkWEfldX
rbvs0bfVBRF4nVcUKwaPwLq2YqG+27wkKdpMfTtQbDd7pCB1SCGYyeSA6fhyg5Ot
7WPJtqAPlDKv1X4mt6nVSQTEhG4OcLdcCmN13x9wLxN+S3GI2zre5ux+upxdlDvo
PR3bwT2LpyPr7q+h3g9seDTZl9GkSccaU+8FvF+xQgnmc3Xm4ir1wJ4JIGENQpIr
rmbLEuV/bK4fI33MIJiw+7V4kf+iFS4j1aNqiKpBdIAFpREITSMRrzGUbLn+XeMa
9D23o7+wWy4ZsQiwlhOsXHBnk7Y0mSPWbL1gps90OBSBFsrNE9DparYci+hM84vU
MO+FbYc3RGGSZsW/o4aW6GWOmX4mexlE9fj4o9UdkZpDgns2tuXXq5+3i3eEU53C
4w10uWSIgH4WEDP68BbeENShSx7rUaofWQA+MzX5QlwZMrBfQBniFbohhCJ1gLCx
FwGUxje2wQhi5l/oryJp7BTJ/2xg0m0+N/8IJ55qdu5MBmVhT4Rnrl10Xk9AkexU
uRG/5Gxe09aLLA1hv2XRksSdV8ObTV1JdLJNcIfbnZ+6s7w4lKH9EJSTXXweQO73
Tz0m0AttWjVrtua2fujynqsvnd1meEgBzzR0FC1obfK+BKqbHO/nUPwbc6yp6778
6awQvTDEXF8jvVN7SYeLpd0Sw517T1ytcenKQRTG/F6Y8+k3wudxKTYOIJVDPCev
tIf4SuawcoL0xRpG4NtGRpqFEYage4y/K5fhpBk0FXVRnjljeiz5ONcLxQ3BqeF4
fI7euYTnKn8jeSgj0xw4qKuifcEeb7vWy4tbkBGQ+q5WQSaiUkL9T97M66ZIt83k
0YJHS4z55FvGacY7L9nCGcIxPAntxx2WwdAdLow6kNz/9hLMmLTqtYezLizelPwH
E3EEWaEYfV/yE8sodA3+TzapcJ2KsFZ4eM9tQEJD4gObVe1eaCw883El3XE2f/hS
FNiMugFpfTe+VdjkernvcGFTjgRMkOonBF2+4skCBEjqupyPjffG8Wu4uteiRoG3
8XsQuOA0olk8NTVsgi3OjxZ3m4QX2+xaF+Se8eKx4fbCUbckHcagBTpMJn1AnbyM
dXIadQfrwYuyQJXDPWEahPtn32JwPuL35JjJI0gsGwhsYaYV6IlZBPNCbnmvgiCw
0HigvKcNqALs9Bzkw1FyQJDBQzFXv9W+6LBNvz5lFiDUsBus6knzq/HBMRHrE89j
2H7xCx3c1E1lTOFsvy4Wy3x9SngBDJgLDIm6IUDEveUotiugL6i8rUtSe7dpqWeQ
b7ewI6qh+GcuUYNwLbI89ba3d4cJ8MYzijYVehi2numSf7jp4aokE8DkRD5BljX2
UPmpK0i7ZLgGzClrROu6RmXNJTFVQb59nZvgVw3i9mC7NPRmBOTu0YTSd3kZL5zG
zFxFfXXAS0GpjN6iQkluAW8kjygy+R3CgPOgm0l2L2P5SqXYJmwjrGZbGje+nt70
hSycSrngyPWedhSreTSbfWMYqkbWZ2CXuYe22NP66y1P+YDt3os8HiAjn+6WrGwD
IWA/lfBgrJBmix6b5b+bbs26hDXweN7EJHWpPwMnPneV4VT3lMe2p+Q46klzThAw
OtOeWmZ8Oo0Q8PO58qoCs4f7wd92Xd2tFTp8JHQHyYiw5NZA6Uj2DxOFBSmxI6/g
o8efjsu07ZlosZV0cokDA17+nnrFBrXxQGvpJ7eJL+suxclKm1IfQ4spAEFaS6lU
iRgZzcUeWrQ+RWuv9nHz2qKY3o973ubWxyM81UNg4ZeYVHCF+6XSiismcZGcGzHf
g3tjW6OEzmjN+5OmN7K5cmmP7dsBVxqFbo9PC49uc8h83SFtMsaT9nwSHlBeWMH4
NyIYiQkkLu/vTFKUlgzXyp0gx5mr+P8h8XN8pwh5jqrLLHkPfrvP9HyAM/NePsrH
sXFwFBJSYzAzwEQM6RsQ5IKkTSaqNEULAWK8WHXZWG26wEw3U+ai8vH0LYPqJjo4
uBcRCTwGo7Y6Uz+dkFMlNud5LRgIg6/7EKLM7WA7MVKJFOZLeLvwj36JnMNc/qTy
/eEwQzjlkoT2NRaYaL/XriDz6hnBQeS4wbTATXEWXuz3nTb9ZRoSyUwmh1nUdxu1
kgIUNc+qefT3uLa1F8EeSRG2Jy5PsDrHkbB1uFPe+19oPQk5bdKnk5KqJ7k2Bos9
dUuw8lw1fA1brrlwE5eN4U9/aLbhT6oZfFIWvb8/L8xoZwGZ9187OZL3z7kdXRFp
OINyYDFtvIN2qSsd7II1ZXWvbaf6BAKwS7BVar1EljAAnDjXNZ9kS3sxKVDswt3F
AJLKFIQd9oimCKs4F9ctfH8T9QJBdDeqz8U7K1Vnr6OXjS9kjDIQWKJlpBXkRsqN
Zk6KqKnS/MPJKhqoWmfk+/EzXg3bmmOFJeMKN6xrwSEyA2sOOtPLliRx/NVORKWn
Y5w0XM2oQCRyn7fgrftfbrsy2aJBPDr8akVPKXz5TFa6/uUl75BUGM2ekK8P/lA/
FZ+SLi64NYs7JplQgXIZ6zEqIkLo7gKhBULlX1fmloBhtIXbSLx3uVtxurROB5FO
KfehZcrnytMpqYbaTlnEW6YhqNQbVPqhi+bCjNhzCC4ZnTHPuPK4rPHhZpp4Pq3+
H/kydyjmmAssqbizvWLUAh91JfVr8tScJCBkyasX8P5t5xs4tUsmTo0ciNCpH5Sw
7jrwHtPs5UVfCrRgJiBTFSu6yqtloQWJvxDOx/XvKzY8U/UmsymrMrIA+RQAm9pg
FN9DugZACx6/Qa/Fnnyf3LOecfnqzEQ3Z1BuXKDm1HTrTDNE7P6Mdjems8JsgYJz
XXfxwdU9goG7LjNqgXwfKleJ06qzgbs5EhxQX1HzL7Ro+Rm05kHp3NKu4uYgJ1Ad
SON4tlDOOisrfjewc00i55clO6P/BYUOJ9d5epWdJJjBBnyzVHQo4S1N2Ovkwgis
X8b9KUljKuOVJBE901drLOzik+635ZJQB5cNS64tYSDoslN6u9uEM5Mg49BVBy0l
ZTwkbLIIsgK4M66p9xWMgO63q3ISD9bPQxiORVxoh4J79AJD8Y6VTroCQ1bXr3IE
UdWe6WwyvzNL8UVRcvpKINkJXMibeqVm+eEjWTnurH2bRxQgtI3whks2hczFm89R
tJzUf1ruLf5t4fqwoTbwTP3aV8YI/QqPjEwV/e6zjgwq9zmBdbDi8wRxHFw5+Kw/
Bk+FAOZRd3m0LKpqGkhZ11lVlkta4w5HadBcnC4/PfbtwE3Ep8srTQrDqxyzn6Af
P4M8RgytBUAtXzO7O/88jlbYu/nE38Ovr5oP7hFGkpGCzloe079FC3qvrtyuwcVJ
PI6UX14O2ufAKc7FX0Z+C3GtiV8YJ514YGr+PniCdZp73VLmB4Eyaw1TPsIofgpj
Pr/HzxYl42WEFo+iEsM+3XQKYsX5XUICe93tQ5cuX8/yxg3jmEuOqOg+Yb0+CN9v
AB2cxYG82urq2fdcnoAdc2vQYpaO7L2xFmfDmftQ3TG1ZaV6ZtcFk/ObFRrV4lW0
rW0AySgz+1GJBO6J//SjK6/2AP7SKt5UKfhGyt+mQu3vJ+C5WvBjb/MDYszVOSyp
gQgpE54KGK2TGwccf60KEP5ZQR+ovfXSG7G1gWWxNankn2fcgiydeT5TjktQyj9X
grmis/2dgJYC8TM0boKqDpG9+4J8L53LzKiXSP5NDR0cSa1sbVHHQkYCcDeDjl0E
6OKy5Ivzlvjy/JLyFv4qq1IYbQJ9g74FPWOfU2BgB5FyHfkVv7JOQdyDGKZRMHUr
EbpDcEA3mWfA8UR4ThGn/rKg5KvjEPs3PVQ5Vnys5Cn52IVzCFZ/8VMcdktvyNPi
usEEYOYfNshlqMyNuBCLmh499Om+NJtzxZNDO22NKw6gKZ7NznguTderPsL9lxU2
ah+NOxTd7+S1ZOJ8dxe2v1RM3BdcCWBbulkhdbRpJIOSruS/K5XKOg1G7JcQRqJF
rZTXYESyw8HgLPKxQcSoO3XGzsC+eSPNWEXTIadtpq3N3QZJ1EA0+tV01cAvP5e4
Bgezpz4Hfq9iqXqeJdKXIeziyQRhHURkL1Mv7ZInSEIbpiu+ZiZz0EewZ1ZKa5Hf
7TKy7zPuEbDnB8nMArZ57CVXeQwO2wbpMCcKGnwmiTZkhRzTaQkGbqJDspx4d7au
8mH4ft/AJbH9SlHi3FWoyYGMKkdC/nawZVnk/UGVt2Vfyv5XIzSzd87Pe0oavrIn
0jT8t1diY1UV8ptSY/N0a7xvNB6Z/M+NSoIE1+UCPGxozVX3yGdzLBGsx4X3b1dY
aYVp62cFMLULtU5UdmxFxQp4seaX45t2+WE1QPjkfgsdIXjrF8cW9up7OL3il/Bo
rtx/duprxqVD+B3N8NJgziewshp9xytBrTpafB64Af7vuuxnuHA5gc970oGO+ovz
durNm9FX30H3gM/ApJP+8KzNaUtQyiKx8FOSNsg+U7HuZ/Tp0JEBaLLe9V5u5f1r
2WJsLKhVpep6W3AtSC1ldKuQ60aV1hL0KiLHgubaIhlnDJ2ptHnPv3K+9+4ThOeo
H8leBMazPxY+HnypOKYZHkMG2jBnBJb5uaqqdqjC/F7z87tSIcsf9msOlp5gVv5V
TCw9b6xXog7Y/esyL5776jwCVy/tyb4CkYhaptXtaELKuSTeN+fsg5StxL/Co+gP
d/sC3HiH61rAc7x8KE9Xq6pUAaUmGaM7LzENSJ+Ni18qzuq4FHFLemtYslCjyeBU
uJpGO9ibFlTmiVtg8f55wsIIMTC16xZyhIn8O+bMHtkoVbM+02Q+V8jOl/sHTgfn
bYvK3YKMoJn5KyAg+s3WCnKL2U5MoAEqUE+Gi13h0nzOAqgvPJC8UXc8IxqSxY3O
VR4cEypiiuoWZQFoW2XEiOpQwbJfxlZuLgAGgNPOstc5LrXl4pr+S6XQChGGJkLg
lpr2VAt4HsCfOrkLHZJxC4UUrKQo35V8JZvSPiLA7LqrNQEvltyB+gZapPWU9sYP
T5Rep3p1nSrm680P0yEBHQHIwoZM430iH8iJI1QRqKawgRLJpLTvYCFsP2ZmlHmx
73EU3iXtE42Qe47bNQ2qfL+oAcrDsd5Z1k+qCXCF60SMlIsv7KxrKz+0cJBahvYS
8lyftAg/J52biYFHiHSBB87CzUGEGyhTk+HsWyUu43p9+Cx7wfdAdGdNDTnAds0U
a2vXi2qlWlECbnYhty9WT3PoxX21Xvg9jrOAcz0kUtWQxlSOOFhPMfJ8cAN76DRL
V5UTjjDaLLJvqZd8q1aCA/FcXW2JENMMI6vS53eDIlW5Z3pkJbrc2czJ2clTf0NV
D5md63Hnp7deO09qGEXHyRAeuza1bDqW5MoEbFd1oWCpBoFwIAdiA+1LqJS+yWZd
uTH+qTuhba+XZUy1ZzOuWjhYdoE4TjCWQLO9Ztx5bjsYod/Swjw0CUxGY+hvXAmu
8onOvAqU4KIzG2VUaGu81fjNewNdM/ITJ0hcUqTSqMbwrWjJSLEPludEWshUfpRv
uan2EyTqYBXP2u1lD7JY0+olvlXgmUxH4QVshMlg/jhD1UyalBLuoBMNyAG+8vzU
8u7hb/hkeMIhaJbr0OQ8+Wo/7AIEp6DrZ7RJYBNmHV3FQengVLschNWb6yYZnpz+
rHquADMh4Ot0yvm9i4x9oixjlFuIOQcgqGr0Hwqga53rqnbbATVppMlfygHcKTay
5kRggNN0DRp9ve9QXO6Y3SJPLgWXOAiWzdMlCb+eWIIWK2w7Sp26dSuBzXvlUySn
x1E2xQNrRGrdpguB6q18ACTIXR6s5Tadkz7izBgTFhVMaCu1/ClGF/u0LZ87jqyz
JrErGoEyGRRzD0ElGyQwyBA4CYtmQkPpF+lcYlF8mWucXdjrtHoljaqvgWiklaFw
brXwukgZX2a6wHbsUMZz6IrWqWApXBBny7gDOuaVq+KHILobPKoNGRXo/y0zymrG
PrIG6K6uz4I5hMqjWGlpiHVd5e8DTa4MUmkvN8xnenRmZ3xuSFzHUd8IEZW60luE
JfyzG/pezYf9/0LEDfHAM+Yi4uqoII/gb2JJcEGNzwdYBmwnQvXQ92oPvFJM+4mC
/8xoSo7ePeWN3/4e8HlfCq38Lu71SrXd06oI97bfl5jWz4riMcFNt6G7Haxg8kUQ
oUv1AocuCmQrRiq0Jveytz2hSJurqS6m4pnTHHbEiySyoUxcNctATX6m/IvZ3O+P
cJjKv8ebR+ZT5Gg/Zg8WHZs9JiprtBLn6jwewyVoA/xQDl1x95DCSa3EiEneXmuR
K741XQUpjDWLZRf2ewjNX4GBVkKoYLqtUvgYIN5ByIdwX+Xi7yCUaZl/Y53ymgcP
5groJzfypJ2fGMG2iW+GPELULv6IYyEjPyIYE49rYjJwf1whhWyBeBZ3sRDeQUTH
ti83lEg4zPJKs+uFcTQg5lcNvpdn/avqaIFTSL1frnhxmQqwIVAOSMjF+rhzaAAX
4ahNq+5HZc2AQj5JONmu8S1XN/4vY/geSiScLLTxhugnzF4YAJbj7xD6QQz0urlO
2l4WgRd+0ze17pxMMlhGE3zaHBzgSqHhpbzEnEAzFK3k0MAF9QM5uoB+CE5k7Srs
0aC928QgZU5J9ryECx5yqFUp5ZcXsblz0vdhbk4qStBQlDW0GOQayQdmQ3wmj1wq
34gZmNUycywn/ps4PUAumpfdu0IMBGE6nVgzROzd8QZgaR2577fnwLA4X/8oWtVP
UVOdXhQiqogoCJhwk0XX4dTo5ikuhhLIzj90DFErIZe4CXxilNWArUfgz1t0sLI8
zvF5HlGeftt6hZ1Q0HRYN6+EpSuJbtINEg+Cg0cD3EDBFFszQg6QyB888KL11fP5
C9Q79UdCqUEo7MQX+RKqPwjfSlUKDULXyUHNX9blKudeMx4O7uCVzECTgPrdFn4g
ulA3XoK/2EcSxinoR3qYmhBd8EWJkfhnfArZ+alrrbetzfCapLlD5hGbTKzVMsm/
ID0ccSEjAVYKuP4NavcaBUHFpMYsIW7rAejV3LN97e/ObPTJOA8VdwGOc0k5WDMR
CNiLpi7TvRFQKDfclGP+KPfKKt/Pn4l+oXwj9SKjJCloKy+ihSn9L7rzXCEinOb1
bfAnK5knrmaDRgiYBxuLV5uthU1UExwQMEPfB6JkrRK3AZI6+feib2NgOv0FFVfF
KGxpOqIxANK84CgQA+1gW5WWfIRnGHQMLQAzrIvsofNhraupGcE9hhF/XrlHlqV9
wNVx3YDEhFQSQg12pOVNGfDV/ueiCtiq97Kch5pqZviqSuECbEIkHnIm5tKasnIW
OkOBi2kDspLUNxT6fULZxh5sk3MsNau3kDG2Ld3UjPnmu8rAdTu82dk7MQDLuUA0
7Eqd1vuGK2plu0sjKmf57GByUQfsjyZwwUOkINsSSGUFm89/cG87Yn1ZWIr8EcfB
QVyR+TqSBCM3W4+0Z4Mqb2YOUiV0DmzE5qyaIDCOwhf8kKvLXhidOmIn/IKkXRre
jJsOQ4VjrsA+Ghu9Cr2bN+G133ZV7mOBsKyX3hpYQNUpfvMO8HrvdYsjG5mKnIyF
/vAa6+MWXPrhLrNSP/fRxFMxRPwodIgzrOyzLRPZYMiFLbarBAH2JKctVRsxj+sM
cIVslLxUK05FdDSK2YqY5lrU359qBd2O9HoUQE1UKLckav+EGOtRSwGu46d8bVNF
qWN1Zm/ngxbn14NITNdnN8sAZeuGzpQ+D/Djhpza6v1fk/55pv+uW4pMaj6r50dg
NZfu4ClcXh0zRhut76co2V6cn3VjOyae5Z9tdY55hVP4OFkI5iRyagMdGE7+dDak
Q5BkFGPpfFujG2HsM1GBUFJBRhQLrzm52yq0NinicdmJNiO/7Du1Xgi3oBtpm69C
XinHpOzu7xJ2V6U4wrzzE7CkhEsknJGl+7nSwofqUkocBAHMNR5VEkeYe89aqSeU
yjJUvvTzVpFxjKyCtvaNT9ICC6zHCr4/tX590OPowThNFIct1sqZuZQXvf9g5Wmm
NrfmySbBokBhjAYVQKiKJiF3O99DujUnFGWeFpsEIoPFINSI4l7g+txUiVB/4lNb
Kn67PpxoQZ+uDzQto7XUDJP8MEzW66ziucLiBynAzw905DmpaLnAod5DdZPhX8mq
w/PU7TgRNPtakG//iPGYO2aZYcz0X8k/yOPqyOGjwdsnGlkFMhGXIumdfkj3tnZG
ZQPsbe/71zelAAeauGcu6Mc72bXp8gqnktcN1TWlb942b2CnQs38Tputl1ug9rpq
IFbbirxMubLYFS9vxahlHpHHrjXvzesIAs5TcqdMsCKqi5ziP3DTNGdXE9dod1Co
rQw0fmcrCHEA3fxFx7Dm/GZEb9g6lcuYAmuPjeqN6FvfaxObFeH6A+WtTlN31r7X
zBuMsPjOlgEBcHtxuPg4N50MrVKa1p8syLjZYgzkmWpZrqAMxNkmVgZ61P1AwM/1
zdX6FMf/H1jmCL13HTb0MZI//WoxGEl0dOaB3Ng9TQ42asUPllvfwcCS9x3WQvrZ
UXMeFn2RLdRTutd8kFxMlXqwU5BPvLajySFC5cLZ4u76i0DpVQnHrDf8G9IBvCVC
GBzzsaYvd4Jqtk64jouKUwcoRnkHWJ7KVU/o9EX5Ik8rxx3Zci9d2AeL7xyPD914
X6r0zxwqtAy4xClJIFa9qFdXjVsBpuolfqF51w1O+ydIsN9BGRZ8nuoBm9KvRRX5
FXV1kFRoRB9gmfGDF7kMnnTe7HpgJlmFGtAf7ZHzdZFmhSLvQkjNbhQpeUCOTdyL
zAzapBvMYE8c+0Sy9j0K1ubCNGxk0o9/IOiveNcgLKY4n0Vj0ARTLWxBBmd0Yyvb
qj3m9/f/kGC2r1Z+ONJQbCmCyFWTtpg3YRyDAN6SRGpl39ZUUq+kHsWOVo6vC9sQ
6IOCIBXAsEOBHof7Ak0cmMzcu0fJsGjzV6we1xdzqg5YpaNS2hNdKFRt7bXajO/H
fPma+idByN+bnR3O4rqAh1WLodEKsmPyeIG5gPhWdir+tiy8YRqDDa0Vn202dE5c
9m0/Y6VPTIQNQ71KYvUen73Fj8gZ1BhlPmWqVXhUGvE3387NyU8WQGmzXyIicj4m
O3KTC6AbHaJkZoYHnNISC7LPNszOcrgmOYDPVXmHR3lOcgDyT4u+yg1N8aT1H0eS
AAHxQzoolzR7nrx5t9XIJHDfkjZkolqMt+V9BwLNg9FXn1JUh9oAbtu5hagm/ls0
Olqr8iBs30dhKDq/N8fpT4/rxa+8tY6PNW0rgHebNn6+I8IN3WCkThgnvjzIK3H8
IxnQYg2OL7mbQfOLzAwP4JjuA2M3Qhc4rFI0IuY1CnWDjILas0vGvCLscriFCdd7
0RJ3z7PKFJusiJ1HzhgO48hooXZ+QsZYWMATOrZz/1kcsoJ1f+z3U40IitDS6pwP
LppQtRBrqwoDoNNRqKxhHOZyonKEkEM/PpNDFWChVKj6ESx445HRZ3XB2/ftm4jk
iJFzVRqaCT1ob+t5emLItIti2cPnp68SU6g3N+FhqstQ2e0FUgAEVVFM+ZTNjWwz
Yr9b+5T8DHn0gPGCMgPGfGLxpBKdsBTZiyUp39ngL/e912EzMj/bNjJdwHDP6SHO
fe9QtdpS4tSgJgH7AEoDTAvW+666l9f6pT4XS6wCIh6dSzT6msaWdxI9Frw9UIWA
lv9yw9tQDIfNTtovLhei/DKHrzxHXxPZcpg++5NNDCfI5WyA1gp2vvUVH/OMZdX8
0tVNkwPyEm2ZKwt8d6kdU+j/rH+y5lm3cHZxUllEO54mkmHmsrbzE+KfO8afAVSb
DQSM9rBQn6ZA1eudUJ3KiLtYBycZ9P3mVmSjpHR+ndEE5pUS1wg0WT//bfz9ZbM4
+MguHmROYZYePX5KdXyei3/rHwYD8XUhy2Kvveb94A5z4o3ELGyP9GM58NgoD0kC
1qQk6fbe4du0318eNFZokiY2sgNKTgwLEG4j/ntdsbyKeAUwehTgl/lgdkw9TBMm
D2xUMXry6d3Zcfq1Vijb+hfWdEAE2EpdaM9PmIlyD974AvyvDYH0cYPibV0gEDwz
cLF7NPdI7aup14C7V5GovksgTtSrfTRlTC0KiAykldnUKsAGMN3wMeh+6BQkXZK+
z8pTp5KCzoTAYkFmJX9V7uPkAXEvIt8IshOyvWOPz/f4Ty9ASWbc4/q/nHcdWb81
N5L1QC3x3EukvIWJo3XuH+SKxAkaCR24czlOhAknuRRZKSB7TzuW4KjccQkSwV/a
dDaK8jSBdMxWztXHBcqJh7+rLdZFRN6gKniTOsZlA2bep2VZi+g2z/77sQmxZEdT
DsGUgA3wRO9oCtLOJ2PYpf5gImQkyxEKbS69INPDJt2tVl8+/N/yHPp9+1XmHhpz
J1f80xNMfYJc7TMcnbmQRfDcoIdnAYT4g1cE0AvjCWPvvPH3UcieWvHT+C/47heh
O4RUOQRBo4Amy3wweLoYSf90mgzEz69qcjF4gvmWdFSfdEW/gU8uTG2235s2Dvte
gYwkLRmVmchGK6UXx2MZeB1b88EUXHWy4uvrU2jFY6Edj6dxZSKGc90QGpP8DtWf
VG1UgFUOOFOJ97K3v59PZoADtd4U659vBJOonKKdnW2grwyXa9nbFjz3hseIo7/L
EZaxr6oWQ3YycN/Zpsrvi1HbFTsA5RYNiqG08MDRxX0Abh3YJvKngNmIT9ePtsbR
+6MlRD7wYKulLSgHM+g9NES2qQWJI9EeizRHw+m3azjo05+AbN2dEi+ZoLonybJY
YsCR0yJ6DmN8O9yA1wOHJCR2Qcb8Phn4luhbHX84zWBVBtvtuC2/ZukF9HhckjPS
OSmjPYvq3CmbyUlgeP9FjdBAIrGcq/2OxEfLf4miq1qkwWncGX7prAIMHFhtYbGR
LG0JKwUwfuHfhgNlUKPMob1zjMRDd8kR22yDaZhiyp9EKCPz3XHWxfEuXR88sNyg
TbQC4phWpXD6M7QCSbEj/10RbaM1ux+CjkJ1K+noJNdXkGeWUQwunyGBJT9su4qU
B+D979QPh0vmc92ZR3X2nsd3sKS0/4+nwQyfCGdaOk6qx5vHFn7Z0ZSubTgESbZ1
Y98F9OuKqXLJKajAolHJN7h6pKfvsls8RL+HOuKShQClPqje6cuB4dmEGegqsfBk
ZzsRd/OXxHPcRSFJat0Zf4b7wfbG3eCHXNIY6tbDNbqoYQg4sgDaTyzJSLTfvHv+
mOEOyDVKaAvMgqxIPi6Izd2TI2Am7aAvPDLRGHfIz3iSfuhSoPeFbu94/euTYdEF
SphqJnkafwAoX1g0yADLp77fEWV792SPWNUPGTPHAlAjJFiD8EzduEarz7vRdgOY
62Jty6H1G8AlRXlkU16qM0bTg8Oxnczv6rxGu8quHKLpXXZiiL/5eLjZvs0W+NTm
bQ/L0LXd0G5pO0l/mAvSrI+7rJRhUUj5ncSdQEEHC8JhY/CH5AlDDnLxGae8+zqM
dYMGVTc4Tn4pxHRt9vB6fRjnMpZoNB4D54PziuCkJclbe5rnBA6jFdj/EXjLadxg
BJ6B88dubWSpR7H/YRfYgLawGezQQGSguhE/4cwWucStbfR1t/bQKqeqd+LeV6Rp
UmDhqz4G9lx0EXCLXQ6cW/paYeTGhxUv1oFOtKuEJlGGK9J2xIxWZ8zWM2cRryYU
3QAGuH0ndINbo58gVNZtsWJ6c55I9RauhiW6jJQq3SrXBuTocV3/WwzNeTuW//Nn
is/BSZlFqtY69zlOur8KGsREBYGx4krcyMGwQzLvUEl6qzbd5CR8RHFVcjl2kfvb
U22gVeTuuiNibXfUdQrJlaLCta/P7homsHFJEckF1uJfcD6+T8LROC72Uk/8gKSg
Uy9HM9oejSItKtS/I/Y0fc4OiBAgrYzzzwGF2nlCUGQcX020IkKkv5YaQpi9PeoD
vRaHC2TK3f3g1asgRK0evleOg2HZbqXg9M1NPGvfiPmJj7x+1u6mcI5W+oYQ/Wow
aL5/dT1ulsJ6tPx2mNyUJOZzIpWlTKkDxi4SxSP0l+3RmpaRjmSpe0nkuCAsJMY/
QR70qM0JjMYiFerTV6r/oR+276S6kCLCmGBLRcybL/oLusaxGtH9l+UiveLIEXaG
iZn4OooKOX9bix1Kvc84H3LD9u4JBqy7kfXvkBFnf7pQpt9+W6HxlpXbq06jVqsA
xuYwdFhjozBXN8mqyJ7EW+DDmQ61vJTXsiAAU9LA5kpMqkXxbzsB6VaeA+IvmJXw
i9ehdZCUt+qIHwbJ3YF96FIB2YsRBsghnBym09JtgdqWcz3djaFQar7zqZAGq04V
zoNFztdlEAkn56yoOJZMNAudWY/g/T1Q7thYx9iPVcMRzfduyg6I2YsXLwwDrImU
ZEAoW+1y6NHzUJF6/6oO5dKYI4Yu5N5Z2owZkQDwCp3xzn4vyyhwbtRhHZyTKC02
28roJteNDu4zrU9IP0FpCBW+0PryVpwdejpwiv188DKIvNGW41LcFnB5PQpYQWmY
zWpd8GUgSrn/S9FAFvz2Cqtuz7hSk5+JLovbHALY0D1VSDv6zA5rZelTYR/H+Ii+
AVOdDlxFrategabjxPfiBoU24W7wZ2yfGgBoXzhbDgueGuDallssOtfAN9DT8Dcq
BCE8a0yy9xQglEJI3YPMmt6D71NgMfBlIN5BJEo0V0/mxRB47I+EKyREVB+P12PZ
jz1PY5Go8fmIJVWwOH7tFmjoFzdds1C1BGBjRvdd5aazAuPZwmgwSUaFOBFCIQUj
0ZaL9ELkWxRLCqptIPxARqex2Byo0NZ1RPmi1l4QzqdQ7mTn0Kr7yFTouFGCX2rx
OvCatGSjs1obSbTadRG/TYqeFrBryQRPwkt/DtHb/jEDt3Vm2P+/YXCRhTKW4Fft
wD/buL+Hz3d1adsqdkf0LSrisn8toBfMv0JAlX9EkHPnG/tPjiufm9VFHSpqMmdc
5kB2EKSt7pE0IVjgDXmi5E7USIpjTRzpmuMaLFs2ag7qi0PF/NdcPClQQfnsWHax
1Yugpq5KY7iBLjF348Tg9URFwcO67IkmeDyGKeGctJ+7CLt9Wn/npSLNmrS6UMKP
slBbRl5amD1SOAU6uQc2pDzQDe7naCPYPHV+IdnP70Tjj2uy+ZSUVxAIGgXl6XAh
UODtSTuPxqrV3yuYxDoFHxwfMHIp0LJ/KwXiBkkVFzoyqy94r/Dhda6jJHEAQ+ej
mRxE75mM2sAvxFXqv8iEZn1fWG7bt/POI66uG+cecKaiq/WX0XZQ8CSWxgkzG8Y0
OPkYWHHEV2MjWaStlRVWukf9nk37PDCj8fUR03v1CwZjMSYQ7zF6/uXOGZolxu/P
gVgw/7bAavwATGxEmDxZGaWOE1Lva1+drLtJ2jjx73qdoHdNBWqhE2Z9aFyhOPVH
+QKLuomY36fAzl4W1a480WuAAK+VggQIl6i5dtjtdBtyCVU5pBmQN8UPy42dq7pR
t5mfT1qnsDIB7rkp2krBh3OtqCw2FiS1r5r8p/tASUSvdEi05zglYbWj1sp73PZr
kXvm9Kj3A1ZhacQLrYG9mjp5gpex/JxdsVGQZY68cKT7P8+W5Vt52itUD8kyij72
MZ3iEt0YLRZVuLpA8DWKaW3eJADe7lfdYxV6WB6NRdkTNHOXzmVclPTVS2caw+yX
inUE0FXjr3AcduNVltFJe8n7rq/vNBF0VqDrQL4b9RhLqOsuwNtL2nDU6ERGhrd7
R6XY5fHMdIoLCQ4cW+LTVBFI1HoLqzegtRSMMAVBWVRuEfdNGkhHr9oNp2TtN9Nc
PjA6lrD2i3eSADoL/QMhVIIx5XlU5PrbdT68emlsM6MS8NiCvymzUXDo4G1LEA6p
kO6vqQJjIpDFmctkQpz1TB9v5J4YLzxnaVERpcMUG77M6b3s65/HeKMk+weG7zFG
C7Sc+Z4aS4NOUF5X0WkoeWl2mmllbgjeP5cBcST5zbeE0J8dt+LKkpS9x1CTWvOx
8UqWg0OZRon7+0qWKQutq7s/fqFwmYJ3B33+x7GgJUkiJ50bF1bV/UrjdtqsAWyy
hMTDKsSU5lFXRViYqgYsGMvZy6KE9hjBOQr1AhjK7MvqhQIcw0v5dMO2RPI0Ic8Z
7OFy2428X4Te1Z4PAzhlzzE5Jxpbye3enMAe9XoWcqmFTo6OKVGXx21tiIolWog8
80AIWZUmNWaubF04K/UQqBKT5pDdtZdGHpAbsNiYbI0eM/whKIMZpLQwiyh0eu83
lwG1OBXUyJca+u2TyXMTwha1ZPJjMYF6r8/bxqjQna8rteT4FyRcuFXry2P52M6L
qS1PWbvcME04Amr3bUt0sCUO1IIo2aijop1sDHrI6TMd1wbsnWfQF7KQKFuyCjMx
laLd0IEreDnpS4YrDBtD79btm4DrhQR3/Ue/FgmeGVyyP5jRr/IE5O9HGV4QBFSm
GmyP6SBs3epH5J1G//Oza3yAZPLniZOBOxZgNNZL8Xn2bwokGDGT7n2kFwoU1W+6
2z+3LH1NzpSfVoJ13LTHs3QnDh+lsPBvyVvqTZVMCVlj0ML+VgdCtrs/9i/uRU8J
cgGJKzEFAVagJBEaSlWu2UpH+Aa/C+9ju6D1OmQXtqpTn/auxwJpGvkioY9V1q8r
6vCySc7uu1n3A+VeYBVEMhY+Cb3Yyd574+ZDJ/u4rczNp5r9f6SHXfH2+/mfbYSN
JlvBFZ8q3aTWeS6kk1AuxevEsmuXzw07zXeTAsZNPVVjodMQK0zrQSfJwmEADaLy
E1zUAo9kaje3LIWbjo7kg2h70RIrOK0kMFbf4gfqiob1aTfAZERz4F0zCz9nQbWE
2E2KkV3QQidV24/LP7JxODBwx90lxiwsCbwAPhSH2WezUHDm4Oo11E/+YkI5MOad
11ab0RDiW2E/e9WPqIAqR50pZuKC5i7e4XVb1skMfokMcj1KM5kphPbCJRP055N4
L5iNeLFVPY2qVRLZ9M32fllkXDeS+2ditCugZ+K/mvdrc2ICkZ1edmUfjCtSbUju
8vyrlxHpALi6Q7RBJRESlVd5R3zznSA1YaJ9CFrbTMsaOB5lpSyfVRr2ZE1m4OSL
PDNscag7DlK5raa4XLWy8YkR4qHVrLmtQovuhjnpMcV6dnbPcjW4G3BkHOw0N5up
X11D2PCwpTRAPMiecLmUdQq/C4rRzgdPqoNOfuCI1a540W6F2ZwO7kMrKdKcCZVm
e22T8xgUgv0iEPcPwy1rkZ6vT35oIsBrVK3JWlRryOgiynjm4eQpe6aHso4mS5UX
m7EL5ZIU/1fS6cbbinBiU9+3Ofqjwucr4mE81hOA72MgpyBfs5Rks8ZDsPaGOGr4
ZojJ/OeTN/4NkhQsBx41gLoaC1ruh/U4iyHh791hMov2q98039tK9M6z3q87DsVF
F32Myb5TTN2DaFTJyQywSokPHvkUbbXEhn3bAVc1ZZltvso2dbvPToHDDOTfSy4Y
JH82GAySvXiDuQrvsYMUrODe4hCjCAd/yhnby/Rhe4bmIS02jJeZb7wHCuielI/D
D5eg4nNd0uCqKfpBsx0yLO6MTKxuh1D8UZrq7krnP8bV1FkbxUqKnOxHBnoohXVl
h17Ur9RnaJe5pyDaEvN0miL9Ri53ZXFrsdacnecJafd6XmSnKzcFd7Xrna5qakDM
oPq/4yhfqYC3UmQhlWS6PZYUyqUMis1ET0dKyATlV2y9t/sCFT7kbaMmLL56GwBP
bHz+seAzrE+g9hSMTJn4twN/fLhAVvef+LVXL2Ksy+UC8xk4i7J+hHzbnQhe5UGT
WD5PmYGNZIxhCx4QFd9JMV8A8t4kK3Gy58A4RmV5LwwfaOxDDkW8KWuGXPVP/juQ
ELyT/8OocvrFXfl3uQxFdfP4c3gouC9bAlC/N8OwjfSMPeJtRAwOUeqWS0hTzBNR
fER8iV7hKQb/WqM/khxpdKfqc4ZnI8RBfk7JTkPixlw1TeTrA6cEVSMNF+jCxQCo
6PCWvrXHmIuHBZ/k+ryjJL0kng7/Rbc78lSyQfSjpzzRLtZeGXptecRJukGcd3Dn
zI7wASs3I/HtsVbwELdKqnpcSoo4OGyU0z2Anh+WTApxEW/aU+w6QMBqQtppj1Ik
2RcTEHWUE85q+ARum3vjwKn1dDlfAPVPT4WsRJSj+FZdOTnR7GUdvAnjAQLhbpMT
sKCfOtbffJTMuYGGqXuOH7rt51PozGp0cSiAbVHxSZB5rx08WBTHtp1dUGPygBGM
2/sSQuzvI8egZZ2fOWLIpd8tvMbXspRbjwwo+ulO8Gtp8SsLpbLSvPS8VzSU+/QG
doAm0nVKObfAZ4GhZXnP9EcDf7/1aGRPUrlx8iMZ33ukk3sRlmIRF1bbWb7Thryl
k4Ct2M4xTBGBoCWDwHcrQIYJGTkA5Tk117WLUl8/SaegwLn5lXxxShFAKT43R9c5
E5ekqm6m3fZGCNdm4G6HtNsj/N45uYGQ97VhxFNmuj8SB1awkBEtosTW3CZNec92
sKuDraJBXt7ejS9czsXUosvD8nmcTp2SmsaUjk6+06CG/vrPC171IzafDsfXjlOu
Cwd3QvQLPNXzHFotppyHZI34WEJ55THmL5AaBauxVFBDcDpagorAKwQBU7o4FsiP
zCawQr/EU2HMyYxjd9LAMV8b3nHZ9i9+AWImzQh4pBwqj6y/H5ynuXN7VR7y5Un1
YoIsUrWGy8iJfEPWQazXQddtPp3ErgE5rcu+pTyCgVTjLadmbya8MmHwn/esjQZh
VcIx85n6gkB5+BDkZ5h0TRaUeYbP+8XWmVL5NOF4wUXFDEfRe+tNqRjuvvUf/5S5
JyEC4XHT6m9As3rIRiCcblXzYb8Bv3O1bmGIAI/xC70anif/kj62ZCEeIuLhgmoE
NX2b1hCtgb+JiySURavnFJGdA0NE65Tkf7fWcKSeRTbRqgezM2fWwyrb3U4oiM6+
nBND4QXr32y4urni4CpINuFQgRUZixtHZuGxYVX/ew/3RgVrquqMfeVtFe5QD0OJ
o3Poy6EAy22qm72M2nmucVH+wbjj7jTy+BzfZLKDZwFcIEUwRWCcXDW7B2NAxqVL
ODYcmp+Od2Y/IhLCBdvrrTwfXycihM25EIsVGoKj6ZWAv0dM1RVUFJYMFSwsuCvZ
qqVtYZJV5NvfKpAP1jMpo1Ww3p0tgAmu7VON5MsLs5CjJkAz5j4vaW/LDlJI0NAQ
2OmscUH3HKxyJfnhldBsMA8LXrLtwbojMlL9TzT087cde+Nx/7RnlX5azMV1uKiZ
kTuZntbG2G+cnPIwf5H8gwXQKBaeC8A/WKUJnt2hd54xR0lWML0lqpH5H9GTVsyW
sxsELDsAjKcjknVOKYpL0bgFp1rlCw5SMd9EeNH7QRTWYYzwdTEK82/gw56k9tPU
2LYINycy+6FvQukpLGKIN+ugQLbx1zq5rbrCl268epvM6uyy06jfdiz8bFCI4i07
g3ih3qKbOfRs14wgnNwBXOsUupiFtY1L9/1BlR7Tldl8vLZLQvjJagcyUzSIIkAl
JUoPqH504a9X3JAOOGlDnsAMy+tznMS5qvPvIESQm9uivrH8myzfPO0IkIkFIh4+
hPFUQQsLqFDajZQcNLlznHl3XbH5Tcpf6DovLbwpqYyHHSkUZP+FtBYTnRnOuuJd
P7qp/eW85Y2aioOr7MduU3tLYk+WI4UF0BCEQAo8FEpSctV1TxdECnATES+rAm9+
pcdG+JHwX/YXYwj+K+ALnGpurB2qp9+FPpBnsv8xiKom4jwgtSpG5n5nrqkGaihs
p+hRSrX2+R4W4AAVXfhBruvi0pUnDg2IfzZ8w1JNEvTtzy1zNeXe6/etLzQ8isEi
ZSHpO3hbJyUZCEz1hQSVbRDkBCYTtu+3CabGXKjd/I8HXdykbXtZcj8mYea7BxsT
HeKnnPsHpeECzGjZVTjNlPpyM4IxZUa6W1jdNDvXbrDWWRQCDp1ivIDW16H4LkQl
lCRkP30mVTasLBSNwaemJnnGFpiVZnronhWAvd1czuzuLOB18z/7kSwuhxhT/tkE
N9NqDP3WwQdTbIBRjF7elF3cBICNR9v4oDVRfW+bW3UOIp7m5Ye6GRcxjBk/jaOS
K65w0WMtvxNViNgzRT+Tcz6xhTaMx4rmbKRONCdOitxeG1K8JvcbjeUriBV1Wrk2
vxju6W7LKp4/YBzglbVZhRS2S3MuzJgj2NdnhtpmnnSNmIcVu6p9dpc71f0UNTU0
X/nZfVqr8adoXCauDR6m1ZQfPxlyYZvA/EZkrhybSEHgIYlYGLNTWofqTsqPbxcc
0qutnZc5XRWBLgTF+AWsaoZeGxhVxo4A/YXr+LoqGnSv4hbxD4gJriN2BgUbTh0I
4PfLMUaxZKI4YL4DCMH4w5OlnssDPlRV135ULaS+2ap8mGnFePrTK2AP1nrbZrEY
9vmQ93Uts5ck0u9hDNCGNZOeDHkSwHEnbOaZPQT9lrJYHcgMR8SMPA2rqJV6NLA2
WPM9P8D58uXpT2UEdg9EP+g3ZfzTxgpSligr0ZvzE9JiuADzy9knUjAL5EusJR4J
uDeFCFloiis9XxX2e1wYlM/cLimeF30uSoI602CdHYQp/w0lCySkn2wBTvgq5ife
Ul0IGEN92gnE8owNTqLEp6nbnNO+KIePSqpYH1xDt5LnLJ+kdMmjiaKwwqvk/I69
ccZOPp9auE2sXToi+G7Cx32qW51LGIlZa229FwebgXK/ztcSX04nBXfGK3IvWXX/
EQU71stm4oMx+A4RdMNJKbRX5wNVKkdOaE3OvpIiG33/c/EVlTPa5AYew2ZBuO/L
IqJ/fk0gAy8YuYPtwMdCfPLLQSz443h2wBSynLieRwlwaeZvB+MwhKRuU1Xe89tE
i85tq/KrkCE9bhoN4lee5uPHZn5zR0F4CJ9LL0p6Qg/oQcs4DYKF5gzKRlV7HSiJ
dFmSMss+aVgfztn6Id8268kd4ajo5yShYQ7qpQ5+lWCynGHqxCdDZNL9Hr99hGwr
QWwxr6aVPMUfTAE2Zg1rYIKjNAWABdxn3Owl7l8pWfJAhHANB37aeeluBUZU7FcK
eDbj6eL3tVuM6ogAqmW0UiFLm9a+2jDuTvMf8vwXxpDaVGiAH4ZhIAerqa4Jg0Lc
6iLPfudO5u6z0ntuf/323nYVh3JsmPiq2zuRFeA226+zdgZdrBD1zMV1s9xSF5Hy
3Y3FYLBcAVYTmWXPH6BbqingD0nSfIWJXS9PFe8mcUTZI8aX0raOg4oyhd+vwnsG
YmuQg7U+K7mFBPq5i6uXGsU0Hdr4A5uCZ0jrzLXL3+qlZWGabJ7X0FAD6hl6MXvG
lvfqijlukDhH9zrLhL/ezxb2RROSz0TJ7M/VLjnUWG3lHMHV8R4OwfAspzawn65F
qp5ajztZuBG1ammfrSXGHsq8hAn4EnSsXVmQ86bYzQv/EnyRZXly6ea4B9jPuSWh
5VRb1YDb5u4m5TX0owtRM9xIGdNxSSqmrgjtUanQaX3h+vT/0xw40NdIghRXQ56/
JsJLmhds0CzcXhppNpodxsRF893SHsHy85UpsyYgsVubgiYQuKEENzF3yUcdLPWD
vZeIf/+EqJajFq2PrWFo0Bs7zUtm6AVlK5nr2keROi+Rlg8NZkQMZHvd+9ziRUSN
yTNuaUiXXaJsXknHvy5P02UvBMAynUQoGuwQJJGbBynuFVCILyWH8WZ9J2dhaeE+
dkYgFB50LBEZYIWQ/hCnmjnYiS76BxF/svw5jkyL9+d8LVyHnUXekrmoLfnY0bQt
kMiwofMNNzAHlfSD64iw+FUBDCgMiwh808Ll2lmwxe7Lo7mrT4ctyJD3cNAISANG
IU8IWXYTWftuzON9720NN3E12gaGWaSJDSswd2xACPd2a7PCb/1ZYJsmI7Djks2w
tsoRb0DQw+YYAg02+zRkUtX452yAfWC7N24LoMD/ilBzTPYFtwfBrjHANWRvv76M
K/gINpDgr//Wzgj8ZPUzznY12kym8TiiAKNovxQ3DvNSKLibu4youBbm9o1RBT2b
vJ6URxTa19ywK2FSfpPRNdkoth1Q+nn2byFcE6NgbY09VfL4ghaowa08NoNdSYuR
kuy5oWRhKmk3Gm9gY0IQRVjRHJ30A5xeXr/2IHMv8pZsM6HG5muy8YmL1V/XWurV
kpWyI0e6P4LlZp1wVGl54WupWXbcz1ofEccRp70Y8AvbpHYZwt0cBxDMCvcXihn2
XM5qyV/CWiEJoLdvf2qeghg3GUG8UYV8D0NNLG0t2bkoWuMUM6LjPnwndg0mAQxK
i22vhkyh86gTvNOQ7vsoKe4GH33OmT7aoFYBwQcitCT9WgCI2fM5thIsEpjRbcQ4
eQja/+SGx0hnfVKFrDZnOiLgN3nPFlN6VenDT5eysd6yufm7kDzziyjETxwOBMmY
sJCMQCUIem4MSG9E+sFelDsfJYOP5lGhozjdx3JuOveUSHeEUbox6me5LW9icja1
zJMNaBCmbZqb2WIwdbOYR6d2p1HpvtV3anCmPL3DEgQr7vb3xTG2cgmoJeLVsI2E
zDMyqbvbeNWIJMYdG30gcRBtqO8i/xW4zCls/KBIR3D1CFOZ2172HDcL2Yi1ERNS
Vnzk30RMxX6rDPK+cTVEqedFaVWOSF0iZp31YwjO1+DIPJDAZxfDH5I4/by3iW59
PrWDvVAB0S4p2jc1gxhJaGB4jYVf8MUTQPBuCfm6eICxzjxdnab/hlrwYnKpabtr
9NfBQgaHMradkMPsbwRb/yeiyOdTo4shYaHWONeoHEeQdCunUnkBERY37H7s5rCs
jlCZ8MD7wM5fyIaT0PGm0Wa4MwDLqRyvJxe15wlYs8BruzeRjIW5lOGAPvcVA6uY
1AItxvL8NIhmJluUrqpiYjua1+vBQrEmLor1Nc4qiweqH8r6h64f7b74SWcbo4nI
61NE8dfLFGnE3noO/mOS4o+Zd0uJqJcPwu7XmKlIOO8Mc8kY7AIAFsMPy0LFnVnE
uhm1sEBEi9L7WjU4iG8FKDPz/mJAuVDRRF65hHlcLtnsn2jMYCO/YgcVlTkXGKcB
4OfE4RrY/6+Xxse8b9L9ziUkr6JDnbTF5L8ybGW21AiSw+KlX7wAFvUI7d6I4RJB
QOdpuwv9aIjSr6VNJIdCuyV0FuEMJtg+fg+ieobJDrYEwSXNlFAuNEyipCkMCEzW
8iQlYyniIV7bpj1nmzNP8Y3mCL583mL3vF630zfyz8w9CaESovhJcn8iCY+wRc1U
VbTCdeSilUvXWjCSvLG9WbtMaIax/WPnx87q0ZxXgNmMufXi5rVg7G2ZR5GkCkeu
0US7100eGPVM7R84qM/r9cMAEdnUG2IPXaTYgDbxyoqAY/Y9xeL6VcsETKK8ONWN
sJ6KgB4oCPYBHI4rGOgFEWted7R06x3eDhw+rjjwkUhd20pBeNHsLtvMdB/ez126
Kc+ybfeu+Xgu3haR1wYEXvnD2vbKcJ7y7M5dKJAAWgX8EdFcmcN3LT28DWulaQbZ
I4ke3PEdYfEgj+4oU8typ/HhhSGHFCbrKieIv7aIOE2sjz+z+2qMrf8nOrm6/poE
Rav1Khpel1Jc2aBRoT6EA3bCmABofylPxN4eqeq32qRVlEESDbQtqG9koQhR0+Ej
fOUG9NUq2DkM5U0ZadyWLWWmlBe6vUxJ/0eu18+ugxhwBQE260uzsUTOTnvBZoT5
N+5ajXTD2TQLyiNFY0WZ0CK0Q/DmswxZczt8VLaBHkzimpi8/5SKv7Nw13wD2V3w
LaROHM68XXigEcugdICbJb6Fj+kUadykGicEFZjKjXuZyyhOYbPqzNzKoVw0uoxg
ixNWmsSC+WR5kAiKALjUiQjLAERJay/dAwiZR+sHlPqtl4ECWhC//1xOgZsWgPrh
Ok6vvs7aAKjXXCVzRf9TPxd42NWLDZCjs+MtvUWoNti7W+bNG888MBolE53frg+g
qX9erEtf9HvA8kPHGupyDpc/Wyfp0853I8aleEoJmlx0D5lNZwB2bNtQage87UgX
Ser/72A2veW8SAd/xSuc1UBQtgyyTglmH0T0aqJfFzgtAcnrNnK0RmVo/pshWjmY
p0MHSecxrdo2UCmPUJxoZ4+lB59VZzfsFXWEq2VgZXhOQ+Uy0OqiF8ALG5y7Irzb
2ksiN5+q1MGE52tEe4+uqHwdKEa5QCJs0n8HR0lCAGEP/0f0eVbYHmciv6PmllZl
0Qph4Q/YrJURDVeULdoN7kEVTT+EON+hAOeaK9Xg/dkLW/rMEn84uItjIB/PbFXj
mt96HWJfcYd3SnkJRoxR9ZyzGd4c+X9RGgRs2mHQhbcPIq/TYn1nTJKdqvJcG21y
RctyoGTQoN19qx+fMY6TSYYd4w9z1gx+FgXHXBaE49zT3q+S+5OnQX13ssWj3dvs
RFn/94UfrGaSljlZr/fqhaYv2g83ok28JJ8Qu1fOM6tRHlscdeY1SxMWyv8lvwBB
30QcBfAkqqtO9FgzLoJZ1PaUovgKWs6ZohsDACGhGX2rufWLUVPgoRruSGTNeDkl
WhiBKK8Jrnl7chvJkWwKnU9QjZ8B3Ti6jNa/Ua97NYURvK/7vZ7lrEICMFi0sHya
/TqYupaxzp/CMlKJzULBBLhksti6YZP5Ohgtd96+EbPPZz5/yWR/49NCKZs63ECz
STIF6dfOMiqV5/3/jd/U8xUqum2TmVe+JWE/TR4AVbhe2pecRNvDjXKxX5uVBD/w
E+Oy96aBod/Sne2I+AN7Cul041hokqkYIyiel4B086NrIQTffM+wx7EovhkBgI0C
ozbiIHZrIhCrBQ32NhYR8DMVNfX3+AJrwpZY3XlTXG747e0OqoqsnB65vbi6VEI7
L71gjAfZDwvvaKF+da5MeSHo+lh3NyX8g3vYx/508XmE96W1N90+fAHgQV2udU+2
Hoty1f9bDscui/PKLr/F/FxkXtsgELHKQHiSYN1hfJ25kuH0YUQiei+SH+Vtf3wW
S6+c9AMNoS8nubD2sW6oGnSEW/CgyrZucFF3wtH+4q/ehPlMPTWvIoCA3JnPysBr
/zwvQj2UTgR3pstCBSvVnRdH1Fu1OISvJLhLbrtspbmI22A8LupN8ZBiqlOfEBaR
ltXEkHIakj0tzotXmnL1dy+osCED47PC+oPfQycCa8tI1jKiZ+sUzM8BBRoVEewo
EdMpSq1DMRsLbEtwJf6ysjEssx3SwBuTu6fz9p6EpBRmktwwvFungdR8uImxaFFI
2Bn/54eswmx0+W1xu5qvUxXF+rQRCzDq2wycQM5jzQBbh042uihnmW2eufSGvA3l
fZ2PdEhh08oeDxERPvTO6p/eb0pKXIoFSsZn6tChC9oxiqA+9FfA8fqmTlag4eC3
6Dx3kTsq7rXFTljnGgnLlZnJC2UeqNZAWfag8RbD9l555CEfwOYIsN8z8MXEESn4
81kU4HVsG/hUCmbfBQMATso1PWxHQYYfvUo5JrDPDjlxUTnkdhpVnv90mZ1eO9cb
9L5iLX84LH0H1grDXcSuEr+K3XNIshm4AMj264fyM4nIKWww93lHY9XevOTRPZCK
2qYXFQQZcZgNCIFWWogGPAOH2ANI93H9yIzdnRUoxmG+F1B2AoVps5vqTsBLkQOW
yhtl/fF4h2d7nUJE74DXnYL/DNq5vdFKMq1z8ipZQWCyt8HYKMV6CXcNe345gf6k
u5LSKmAz1JHKl6yJ6IjBS9jX3FPpoUjHwQVnmshnlFGbRW93bDA83G2IhBlP5zYF
jEybG8JQ1UKpAbFHAYqY8cLZNzxyghGNSzXm134R3mrG0jiDcnCiL2kItnK01xpF
3UujJd+grgrce2k2JI7WbF1v018+X45nb4De0YC8bwT7cGTJO/FpkXfTGN6xlZrO
56dR/CC0J5pUaqXyXcAWnWtUte49kYLZ8XhvLyfC90toXewqqCQirmjpgT+M1yVS
CGwxOwaOiwNgOasnVJsvKgREvbmPMY16wHdtajKyu6JwXt2cCxEnuq2gc/EO2QU9
uvWm22mCdNaC+eO1kWeW/6LPlDKYbcw/V9g+uBMcDJv1W/M3VpM1bSS7ByzqhV2I
8gNod2kX3v5bglAjbjIPStwRbO0TzGcDRpCTeAh1jK8BViE1CE4uWKlw9hf5Hx6X
66zMBuDreeKK5YvBNgCJ75Z+nejH0w/GuaEJAcLjVKAhFPzOMWkukx956egyxbeS
L6AXxt1hUQcqL/t5MsifGYisKf5CzxOxEGlHviAQRGK6pfsjJydI0ieqo/u6pCqL
qfZUzOuxaOKTM9kHVwuwwfYquCCOfxRqQSpshz7SfKacwtW6sh5+24212ZxaQrhg
+9+2WPDWO33fOt1ggYTclK03H83pXCA2B2FsDlcyYbjXzZNBlQUlOiJQBX1Wo4ls
CMgLwSzrDxYnx9OfmoRP3fq4P2zlYcI3skPHApXqyVf2mfAnC9mktKh17/U+TqAZ
bNhxb1msqy0+rB7PJmPAHzeSBzwQG5xd8UWvb0XPMjm3YfFEnzMj3OX93vFRl7TL
ZLqVAGBLxb7NfafxgpvSdNj+3yiPg776qORVP1ngWGlK7JgZdUI2wlJF01RQlQ//
xpm0aZ/TrdSQeJJAh/aGyEINQSDBextH65adUEe5ggXGA1hD4x+HRthanb3YMuH/
s86XQU6LqZ0gwt+ZZ88w75Gki8gSCFla3Ly7VXTPar2GzApdVXUhcsNqRhES8XLL
L8csdBkxA+x3v90sW+7aqyFslRF1lc8l1cyd5zSM3K9FnpTyNHKkX2ZzDrnvileN
cEubnc4sG99aehCHE+eK6/CTMmrrAxQP7Kq1Bcq5enMo6mFn6s5V8kJC5g0hFlKc
DHW5RXxrOtisnoy9GD1Gmol3mdUF0wxdDSLdb+mVpJxhQhS8BqhUiL1n+O5dt1mY
eSN8v6GXwAaBbTNQ1aOjkk4NteAWgoCN2GvYLFJpd5GIjttyxz8n0HXugLTAigkD
nCTgoTrG95sJIHitgOZ1ZSq1SqFFrqpLBbHccLD565mSbIJEc/2aiTalq14o4HBj
QTmacXxDce6qywiwiD5RcJ0Qj7+e0dPl9BIp9HEGQjAZkqwJ0gEsdtQAQdglNsfO
+u0rzlqFjFCfsUku8BzWZeHDszVIzkZbhJzXczlqMm7nMbX+OsjeHBcel4DMlXhm
dSZjwQRDxTcdnf8pLz74eRdbmVMw3mAYrPPHGtGktOnONKr55nn2j+uMLtP4Z8ej
ceJ863k/xWic8hMV+f6utKhUXyo0q7vktywYE7rsk7VIK5QQNb2fyc7Bn2mio6j4
EUY8+lIQM60h2NgbKtjDNXOMWZ+9zOuRNtfCdma9Uu4v85LY0ppN8S/iVLcdQWUh
twokcCHOlMTTpRDlv3y0LI+9+2uavoIBKDFQQ6Stps1myiDEr0q0BYWFZYBfoYxP
Bn862nSvTbbZrKrOYpcpYrZEHBx3NL8Q1wn8AKHgP+TN96DYT6KjVItD0ha5D/po
3rOYn6B8zStt7aRi5zvP8bFWOQXfDTmxSeIUhOCpjNiWPNB69OBxvpJ09bs28vka
jbOEgn/wbgBXDaNUSZyFobF7v6/EcGtNqLEbcW5cA9LosX0pBGHbVSRFQtB+QIGv
Uzi2/WdOMQX4yWCFLyTycZc/3IedcZBLiRP96X7B0soJwuyDL3zRc+6IyxlC63HG
Wa39O8MLbK3EZWJbr29+vBY8wiUjUKIDJmJ0M2SxFz9GRBcd9xzUB1G3bliuoUHw
g5TyOCxh+97y8ji3IJS+aei3NvfmdeRbx8GZAfo+u7gDgwd1gi0An8mQkepUlKwp
bhrKtmW+1FprZSMFfDz4IpLvaU+5ZxGgA8jKfGgCX71lRi9lrEU5U7v8K4eX0t6S
AR6Dx/ekjuHzpRFhCzTHHmGKCZfrHBDwmX9Dbqy2c1KVcNL8/EEpcOKFbb2CWRYv
6+OAIjdXtReAd4uzS3FE7Cy8YkfKEHY6SDQWmc7YpTeqlXY9ZK5VwWpVO+RII5jX
j2C2tlZ2UUY7JW2utEUS/ZGlnltvQzDykB/1vKVNMBOKmDONG1gRrwdNF/p7r6Xc
6pnMWSj3TBRYVkoDA+hFusxPn/eu/7/cl3uA4zU8bc0G8Br35aF0wAuKS455C8EO
5bA5n4FmBZ5eyc+urFuTi+f3JqALSHeVkWsH9b7G24j2gsVrBfu3NBv/NF+NlqaN
xZg5SBWnf6Gc2OHfg7iWifRcr9oQ428dt/HXDx9G+rQXd+sGg8DpULQ3AKk0yyTx
vvz2VmEC7NKvAAqSiFwyYA7dYLxuxSvrVrhQmXXBKy1v0wjlj+pJxv2Brh/MRV0q
v7c74qXyI0ma1qdAE9z6FqGqAyj7QScPIAO3sk5r/K51QMirLUYRjdTGcdCRf6qQ
KPZZ6LUFdIdr9TfBc5OXYM8cT+15uvxMvoPf6yPhEC7UGrbxjfX3xBzJtJJyzzmE
ex2ER0BRhADwA0hKzggM+X75wYQVpTwy8yyuCfkyfNjl8n+xTrBZ940I02+MzI/Y
agw9zO5oYRptG4BVssfYw4ctDkjtI5Ljhux2Ix60u/y4SUD7Evw9IwbOTPcPvZXp
kv8O5/9XG9St5UdciPWIo2tqz0NItXqqnu6VWJUxYjTqe4sqb9WtWq3VTuciZL/Z
QHZwGX0VUv224+LObB/RExlqEbgQ+O+zFY3xh5RTO30udKtrYgnSVGXLJmogCvss
Wo/xvGyvYwphEw8sP5JFHTmWBRcoMCis7QdrPi9HC4mk4A2lAfnyfXL5XY5+8HRI
0079SK/mz6dc7BBICSxnX8uSiV7HDosLS6M/bM5FO6Xdww4UJFSgvMH77sHyIuNc
cRkjSJbI+wHpFhwcYTTAbwSzSBYEfK4pg91ra+6/KNdNgM6PkgbabIZSS5jbTDZS
rmiIa0e67oNsmwWK6QbYIzFzR0O4P0xoQ6jKh0mUlBDBDB6B3dxEsf917m6VvPGN
6ekR/LFaA2xQcv4KLAQrU3onstrLNr2FxH8qwDbhE4qIi0vdslHtG86sPum86Med
iNTqgZR4WdssXKlkm1Vi3+mP7tW1VCUKSjP8iq/SKMJvk+y1b/PDTCHV8mLCCCyx
HwEr1DYQOdqcEQOzUBOvyQWdFfzG9PeU8E5P6H7kiht0eNNK58rx91UdKsPDs7S1
qKcM9TpXzOePfje1OiLRIyr7hS9MS6xbYSd4IGaNQuxysaQVQR8BEkKsqIlbOqJt
FjkiyYTkwTzO2G7Oq4rQ/JzIEf2fLLQFhhVIAftX3E+9Bw8anHDyyHTOxwnDvrW0
rDL1UANvilQR9FUzZJ/t9d3C6iUgM82djtybIf0B0sWuTCpbDHHcHOcgF7w1ANPA
STYdU/34O7QwFMP5ytPdL2xNBTw4EPKZImcXfnZl3JbiE4QLrv57CpJ92jrp57iV
NV6FWZTZJLdDoPyeFCKqVFYxlpqhH2cWJvKBfraaOvgi/s+5T4w4SIgoUd7yS+is
o2uDPjwSSStzZ8uSmb5iV9zfwtdEEJeFhVCE+ueFJbQcou/Jrg9Cq6SE/qfAKRs0
IT8i1ij2kJUmlhzCkesgNIodN5HbzoMtvrU/VDhK+cSiPDG+ofb6ckYEnp0vMvrO
Pi6TpHiF397VM0wonJwbvOXXue4HShbVHgccVrugQgJHph1e6S2Qo7At/OMdI7w7
g27wvBlK1vvFwesnDCkWH38PSowMOwMH/g/lG79k8x7PQoWUPGzy68KplAGQ3CXq
Ck730uvfHFeEAd0l1aLrTm98OFsLpp8qWKWtvyME94RkJoQ+JBg0Vg2a0GcyzFS5
vgo6X3V6nc2dx74tKI6+csRRw6hceJF3Zeuq+oaD1GVQ84xHfyEKtvdkFgyYpqKk
8+PvX6j6R2m47EzXK9/0KmSCYV4cNwptra/SuO+ZgMmv1ZB6IroPqLPuU9K3mTyg
nBEP0DYa0wmDWxPQVxge1QvTSsSuSPwztUHaiRjQhvzEQcNxQm8Fz7m/L0z0i8g9
u8NFU3SUuLkyGwbBlUfSaF5+BxZ3zpTmE35u8R1zWQrwfKFzGgVTUedoMq+jhel6
8T2Y1kgn1vqbA8JJFi8uL4FhNeMcK+I2TQrKNsRQWvROArOzZtok0AR0YyATNXi+
XJs849Sd+Ny71hTHFJrAL5xEJSbmbV/7X/C59j0uyg5BwX2u+dU137zujMZDmPUJ
9RQnDAMt4FcpVOF092Xa4oflapIlGDoAzTH782Ap8ugQQJDSXJ39b7ndBTMtejon
2ZkV2nnv0h1ndEHqcDW8huYByTOAVVFKWynTMYSSTOO5JZBUzKffq/29MLXZBIm5
MU7g03qGdGsFEyDjP2dFkaF338IDIZJ6TjJTCNzYoXsM7L6cpH0OYfHTpnfs0N1B
+SzGyaIFOp3z4a0OOfgtbEO2hyCirifBuG3Ai9757aDPeQb5odXGydCtZ6eIXoSF
b5IAAUH2evZWfPy5G08AcxCUqJYX5Cw73FA6vgOBKVtRGa0j7IXvbw7W97w+TSKZ
zQuOa5mRrSnD6oqZRkMxwe7EIF5ZesWQwWWH7hOYKCh+n3xA2XsPjFCpHUhhQpss
0+aPB3LbpdKEVlaZBMGsPUgprP5pQUpAZkYUQvgKbUiW1JFWug3CFAszOuMxpQsK
cXcn/m7VpCoMJRIPrLkNpn2fXCuWmMUTRdld7SQXiCfAib0eAwahIpZbYqh074Gd
34kYluO+yJcx1hNDnHyAVbBUdnmMePYqwd4gyMU6k6t4Vu6FwMly+cSjNVzGkm9T
idsu88bueaAUB51tcH9f/WVHJWgko01q9qzmOuKmU9SzvRbqNJGwtePhARXn+99c
b1o9x85jAFtkW+MJrT21Nx4bfvjWT8A01A3Oie2by9zJ177JdCPO1Z4nIVOShrVG
kksCUddlLQpkikl/A4TSywz2FcP2S6E2TBi2aqXm5yiKOR0SG/UsPhFbRqyWiuzo
slsXElrsL8cwcW2j7dIYEurNnT6bDX/JIuVnUJHlhd7fKTI+QhJtqGvsArqT1ESs
rsDNvi8mltmyOZTFnBQCpGSwak7mQKUHSmuY0A+O42QLYxc+dYTnGQ6FyO3zRlHo
BAxu+6lDfNpFF/Vv7zHqyTAMpmpYs90T6rNLV5jV8oMJwwQdyCcSSso+Yi7sSOHf
TikEZpe5BvgK4NbHoxvqVm6sqfQrICKoSr3asnUQTwF8vd/ETqRLFoWDcUuqsa4A
ptPyJjd6InYtkUjyqd1+bUF+pvauxDcsCgcULNH5cHV62L6QJINB5fNiRckBJ7Fx
Ndi9afC0B5kNOCteDjNTVP4WX8RZA93tLPi++k5ERL3XgXS84lT5gFOIg9M91luK
M2ClYSryB1rIRt+EhfZTjhSJCKFUS99DBdOOYOdF2eR9V+j8BrnIxLM82Bb7gJ5E
0RVKytapqtrQBX+bpu81RgAEIgj+kL37bnTkWmb21iVOE2BMwv/Ti844uuXexCH3
DZEzd72DeaS0xbllFQy70/7A+PNN4YP8DDQTN97jx9hudAKVV6OiNABHR6ZyollT
qH89cv267S+QKgGvTF5hjTOYRavqa1JCDIy+AyYdF5TL2R531xOVxJOiU7rYLZqQ
eJADfD1UJkIZSqextqihA0px1jjbYYC5XN/8mEua0gRig5PkzUaNdZXbmkRahX9s
YM01gK2iiKkv5o9Iz9YJ3OOvrZ/toL0LaEBYB9l4YAR3ZSX3WsjL4+aUOmWDynCi
8fXuL7djATmAMYvt6v39KLD0BPV7h6UyuS36DgSD8Y+d1dI8U2Txeml7euX3sGS4
Qtm3S10cOf95e6mY0zCEXUT4iYphTQIxeUBZMdcQ8D1GL9fUCOOgkAKlOytks1pL
3CQdOJ8FyEYVyzIY0zyQqUNcTKTH5xJP54iD4VDSUvmIX90kQUShBpP43C3U19Ne
0W1+e2Y42WorTHX4s1M2LBfNB4qFmzlnw4svcgFOvh9IxswBOTK0JhX5osVGYwWW
NSHaMLiXxscer4MT3QLGDQqJnY+YX2IXdkMeMw0QcGLXTxOHhi1nl091yQfuBU6Z
up3jUnDErZyks33Leh937beabdk9CZMU9X9GF2l5KH512N8EKloCKd0Z/LU3EctZ
vpXIvptOPHTm5lNIJHuebKwHFzGiPyUpEqsr2DSv8INzC8GISbU/mJ3IEOruKQG9
2n5jrBizGMZoZVlmW3gYSIt6r8c/28HUOc1CWBgFiFr1Cv+P4YakZT3dHYdyLSzp
Ft76MKEOoJTwIQSCPEcvE4BN0BfoXhAHNKb19x5mRZzax/NEHUX7bNF/FSh7Cn7K
qn/NepNK6G6CeK+H6sEaQwBkbK5xiICyBt/RmW4nR3/LHhf73E73A+TOx2EWWV/S
9KvK3T3d+w3W0HI9vCvYcpa+tNSYccVS6OXW6JZeRzEyKtMFMikVnldrdtHcFJtR
LFIP0WyINSOAO0OlhSEjcP7w7cHtt0zx5M+6aAyfp2OXxMmjR2OiBTGEsElIkEpL
InTQzV6Bv0ketof8YRYoNEHYYePBaahFyXtBAbNNRy0alytBUZZIX20Z0H5wQB3v
UhtP0p1K/N6cQnZn04yDYkFDm/UNdxbcPiWxJyXH0K38OGw/QM/6za7kin5P+dQk
rb0wGY7LLcUONFeLF73bRKXIcBijfP79kUGqMXyqW/OwjH8Df1JU0TjORX7N5JkU
i6XWHF6aUTSaTjnThGxFN/pxQLg6hQg5D/NWMfikEFLtir8gOuqmHODSkgdzi07m
s0YUoEBcBj2doDoo9JVH2h3BMXRSJ4LGKMQ6GoGrMJJEoTAuReJFFQexEOS+LgWg
0n0o9eKpCk8sbUQNmppGoq2bedSDzm8Y+n5haMmjkdnzSha6PDfvUpqlihUnkk7R
cEN0UcmIqAZx/XiixSpUEFFamXKCJWt8FAxC+2wnzgiM4UvouUKrHOIyPqxSPD6O
Urt6LJ41zdAWedBBVRpsY0LuLkwjDubL7uhSlJ2BpRj6RdkkUmHTNruwPfUBnC6l
4JscjVXxYwImuOiR+430u97xeZ4SXw8vMHZ9aVwOYa4H0+AO2wXg/bzUB5KzvpaU
dnFIf6x7QGk0EW/SCpk6uJ0QC3V6GP9N24Jwq8MLBJvGPn5r3VjndqIoUdKiQwNJ
a1nSgfmmg2Ri5yTf+YAE/MmKNbtYjcq9lJEM5FBPbyY1tZtzRKUZ7PY6ZEj8S4k8
C5/d7mtVdoKYWRhhfSHjlVzPInivI1Q/3rTCr9pnAdDimSWXkUP3NCQpAbewNsig
jiC77mqfPAIDCRVzncovVz0wspkpqmskOihLcD2Q9JF2ZC8HfthIEjrMq2021zPw
1sDOrAix3UOd5zYv2EXz50Fz/sprqv+HLJ+rVotaquG89E/wjXo1HgjbeziRIhzg
oQH6ddkYuoIxKAYVjT3ul0rka8TR+OBgQp1hUP8qlTfhIOiAOomWsUWG1hmqbmyw
JTWS/kQqTgeixjqV7hiBhLcY4HstA+AxfTYRSLzxaJUhFR1G0+kQMkFSdD8/cZp+
onVlys2F6b3eU+Aymp9L5+F/89pAkQimPogyw9EdlciWI2V+b9dcb8EdtJhG2D6M
kSbjUs7BrTL4IzQxQDMYX2Psd4zg0P5u1kd6sbK56yjQuT9eHq2JmhpJH8PdYmDO
rkJKXUbNZB7GbH5d1TNLW7nNBEpxxRhp5jJemkpv5b3DbI6XPZKE/LvCQlAdWxHE
EDBBcQMdBRLInj35JPeX8fDe1iQcQ1cGmH6c3yMdIkG7mkVDK++UDBz0N11CqUaU
3uWcfXJRG6BwrKK+xZAyEUwJ+WxC54AkuwEFn/xWxKeyYerbI8O4Pb3Z+1bWOr8Z
OS2FIgSY5UFzzAnwwDyAl237x/tYFpMp/Qqp6aOOy7l6aOrVsNfPOHHDISBP/KPe
UyNc4+9wezRVDLRnI0oGxoyt1SihBF5lGbkhmh4M6wxI4FyuP4phPkvmFF+X/qs5
jNxzxsYPn7G2TDsZZFPMrpP2SeMysRRNskPeJ9DwTIiOv1OZPOoyz7Oxn5aE8jGU
YW2kNimMhFel1mM1lExXdO/hBkDksAkWDHNtcSQGSAP4KcWfIlC8Kbk574e8GZot
vNbbuO17zwqmKwgLQFiOEFeKnt/xLR8dzH18XR4tr3NiAapXx5tUHiXkoKPt2Gcb
EucjQfQBOYD8XJTYPfgj9Eg5GI0VFKqnnTnsCYH6mBjz2zIzQPEGDAUN/MRIdhQD
5sZOyjEtidF2Fa4UYXvGSrwMJICPT3H7u0wJpitaE1BLb9Rvz1/lwVsNT35UZCZ8
nUAZTh6Vw3vcORDMGJLhPdl3188TytGRCMn6B6goBXyG4N8Xh+xABZuDKLrgVkox
6MprEqp2DUoyw9mhVXEm0XxPIawHJakdTrt6efGG9h43KQIGD//aUvfl/tK5BQg3
T36ZAvo5GzcYjZi4TvOQmBqc1Fe5m+ZJvDkl41cY9jVAMs5W8Xor5tI0tLC3kpsW
mf6Zn1f+RfwPvgBDi3e7TnS2iMAJcwo4O6zpgTRqLv9uIUlUeY5tFF5IVWovwOX2
jUUodBTtspbCKezy5hDHxZxZAgIvW+Q923IQGYLaQdvmrFfxf/XAH5j033gV4nET
z5WrWFgk0iG4HRHUEsdOwq6TUBKURdnuYTzyTZI5R6irOBxErTSOcJwml1dNzA0a
5kka6LqFc0KDZFdpKJtK6DbGlgiciBEO//7IUSku3+Cag6t0oe4W7+eG5/dyvQfq
iyNpDrbLrJ83+OdhZk91Fr+2nFzMsMxeeoDcOaJwDGt4eqKP96rj4qYIag4ktsta
g9fvz8UPhJxA0Y29DaOfuNx+rscYpOTmL1iJowZPMbJC5rAf1QIUnTMEIepSrGOX
dHyY82QVnoZqzcnvbTKYsRD3/u1NKCnAq0Bv/Mx3de7uLoG7EeoOG9FgL8f2fV1K
m1LrkMk9O45ht0be7D1huyhQjZUwcAIWj9/PDp3HsOA1nVYXVWdvfS1Hsl8KglWU
YiIEScC1Ap3LiMo0eGwN9PkqLGL1pAcLErjnC76S1t6XQ2haAfcLj0uZOxXx9GkD
v7nJ+k4MPXNW5a7n25VLsGcDShowGK9Nolmmhv5E7uhGxEJd12lX0QXCWR5U4/Po
+8FlYMde3CDJ2uM4MjYUupVyRD/nNS16gfVtcc1B3iWoYvpSCEv84teu+xAYEn1U
ATZwe/mvfNhQrbmLa5Pyc4N38jbqEcc/W/djW0LLLojMrltDwgzGLrUw+Brk3fee
x3YLIhOY94Mqq4tkQnPL3vH30rDNnVeHkq8FdQd8z8nI+aXkMkvSYH9votTP+jiq
GwHi/5G+xvXo2Zj/K6i5wqFq2HlxHlNqBJkhbayshkhjfjnTes40E/3hzz2DI+8u
bVnCE+7wHmozX60JTURT8lXDlgsUmvRpngyeTfGvCqEUiNmtfUbe/9wbqpD7DxpG
a11/Rj/osNbdYWvB3dhOwswhysijrS61ubf/W35tqvuVOFE4rvOcwyg8PuvIum+k
krM2Fxgg4W++pMRewIYFIi+w7rwMjBAKzra2x1HaBJICpdIoBBfFMKcmfCvQvuRZ
RUpDeLYMVf0K3kwUPHAIrx/EBm9uDCcjcPw+Vh5mcFjhffEqdYx153x2pJ8uhl8S
NHX+GhBQDvl3TQ0JChlqftHvcp3stymYmKY/mTzEfz1CF+PUNUPR88FzIyY9gipG
yJp/QhlBQcxHgqDNT0d/jz1oC1vfi8nBKlNeDA8YAOuXrVf9XKzLk1ZzpgkGJsA0
mXj6HfqJfByF2IwP3B6FZqCKzFxLhsqupp00wMFONW4BJYD0iLgqqKq16Ln/7p63
iL1zt3zJ5F19brg3U3ULFppQukD0WwpNswmm1AXqlHxJp4lO6X292jEznt0TDXDI
XxG+RyZQ4PoRhPFUwjPmhDqFgzmPTnR+eqQX6a1w4M73fEXj0sYpZb84ISsEaPK9
RSl9TOYgSiaqqG+3iXfWL9fvyFoPlHtFbv7b8POPcI2/Dx3JH/MEFW2jlO3lChiN
Kldpx84ZBR8APzKgPVTQ0MLsiqhZqN0ulMVVQ2nARoWan02UdI59zFt09Tcwsdnu
H+3Hn6H76k+UGCom427lWrtpGTJ+rGxQdRdf8dIylIBCOJTwYIljKrc5m3V9ePdu
e1YHRJWyt2yFpbMODUwN8t3WJjbsRH9t+kPLq+Lv9CfZd8WKFbAaawJO02kl0SBP
jslNclea9KgCyo4xL8A0DLKONlMW4dkF7BCopcbkqPUtcgDbNHN8EoKOhbzqdu10
/bROsOVEKkFmIZPwe4h4ifFf599WMHClxvRXDK7GUFDyMOYK+trCgmp8zh40UH+y
WdBm1NwYphnPRkIK0p2fW+BehReKqJOqRuGru8n0Fv6TQXaLpKkd8hucPJb8715p
KXmTNiN8CR3mTQNs2sK071r1tXLu2LFBarO4PENXjPTq+SYj9ZKSjy/Vrd/wIvyN
C47oQHfUhkWcDoN78bazaZc3Ak1qYPhJKnb/azQPeoOtc97tiS9Jd/ZhcqcG4NTO
GdU6we+vCwEGy4MKMhsjD/gBu3NxRUlLnI9L3F/W/Hz2/JFoxrbAvNs2/BLeZVFj
OUR5sdHFgipBGILnXYrRu0/YLyDwvCCaIIpUS4kw2IlqQy0gPI6JK+UZdQd+nUnp
nxuVM8NvlKgao6AwnFGvGrHO7/fWltnueT3X+vrKKRQPammSSyol11JC9Ggfi34w
KDCHW7vFGnqFcaCm/X+vwP2Y1lcVaAkP8ZMxfqJG6Z7uy7Zlctu1eQC5fTqpYnmR
YhEI/R2zXLN8++svjYv9ykEcWY6ctvmha2i+D5sMg6z+TbsGuVhPhlhtDCT3v9lU
B2mwRzziFn7xUbd8LRK9/MkJ31MgYRmsCaGUn4VcQ9wG+1Awh7V0W8G3vQSiFjdK
6Ekc2JXuSj6yD1nbkmlZkPiGK5JKJ0MkWlKsO03nh8vbqvvzTzpqflGf4IJpLUTh
020WxUooGmiscVEbnSKdXaJXa8cCdrznuywE7xv6NotgaKZ9OtOfYX8TV74oongT
jGKsAv1aNT8XtSeBVklzkvxz4sTNxroy+PPF9enNg6J5AW9HB7MfPAMQBNXF4LQ6
WxY1+wycgM+93WBkVxdMM93Lin15q4OSArW1O6u+oAOV2Heak2KkoEEaUp+8W3P4
9XQoi+cyuC5Hm7SHgnwXzX5Ape2SUDrgx4hwFN98eC6cztTprM292hjmZYXA0kTz
srfecF/ifFnnfJRNWJZiPyVSBXih5OMtaE1O1IdoHcrOeOcUNceXga5iWF5/RUZq
NoWYvZif2bFEBTgL8K4sRN8bXpA3jikl4e2JNJlzTONZr5eqF7BSpkGEckKQYKUQ
lmXlrMlxFGd30N1euLHV5lIeYUiiIjSz6Z8magEQzszGLEbs7r5biALtRoY19jUT
HX8EcM/8a2YCd1UycKmKOHAnyJeB9FA3RnO9+V5AAS2lFimux43h8pEQleiqiTEM
WEJwU5MFrDLXgIq9tSfYYwvAIQh8M6fywSAXN4YXtHHuYSNmT7arnlbfBTfCsnLf
Euch87ozqdE8MPTRt0iiJGtqTJ/XjgqtDbN1kVLcUXiIBkqgedSYk0MNFTmWEMOS
2hB2xsjG+rniw/MuigfOyJ6hB01+oapEfPoBB8M4o/ZzpT3VpkeLwYX09nicYTui
q8mgdXaMFSnyz2odMCOWdckp7VPjvxfXX9NxEoYH4ZpZQ7IFsVFpMw0CDkJ9Nqaq
ZPBYXMLzRjWDSHfC1AXs022jMLukjy/78mYxwa/1D+Gigb9Wm8eaTOFHAo88po6s
XMS2vunO240JF8WIVgMjz/mCbEkZl6UfYzdIebjgqqK779oL5HjZb4Z/GjIDuvIN
f9UnkUTnqUDTQ2Um2N5sx715MATNGV3YmB9ZL31ZJUVKzHW++rhYWeGv0Non+Iq0
TRjHNEO6CI3Be1du3LY/eHTP6ZfgFmAXAQQXmA6rg/R4VgrYmfS0VETsg5Qh/Xzy
IHsQBLgkDNuytU/Vso15wEraCym9S9uKz6Um4MyylrOCFIXoZ1Rrr7XjLmYiuVxi
wd+7ZFJqhXLyflP9/sHEiSv9SQM/j5qiV64q8drsOVLQvIMYXvtiYMNGXFDzfX/z
QnixtHF4pKHEo5tcbWZb+tshRjcbixFXaAzcu1PifWM68p0aLofJEQ27akF2Buew
dN/kADp3GXFWJFFHZHvI8htZuugOhCioCGoAvMRsqBjE/hJXSP2TkuQXsnjgbVR/
Ny6C5yc8IMl22BhEdr5Q/1DYZDO9j5V8a6TCDttTv0qzD6AmVOohRngV5gXEY9sl
ZJM+ZlMBJNHFFRpRIUrZIJHOQaAq5X2+qDV223zUDvgu6ZK4LEkET8/KNoDa9lzT
KkZQYBhAiFDocfNPdR3O4m/YpbHvNxV+JbOhkFTBrAcVdIitltqM7FTQkopL9LnA
Kzeip57OCj1SUAeyH0HryYX0KI1ELSpQB0TzU7tZ3I0/6xLu73FUno6geq1rHweF
Ffce/p6X43qTVG8/NMC6OCL5CGxXu8RMm85f7V2P4ez7xPOiP+A0UfiBdCRyJdlz
HvPs44ZC4jhXo9FUe1B1FNxBdF2XWUTLJCxDW6+1F6Jtu01+ypCtupylq18Uo4SQ
Qab4JaxKqxhbVKuZpvBoL9a2T/x91pl1b1JD04VUHrMRzmgPzJ6c2vf+7zoZqWsI
fkvF3Z58K0b/ki3VAofsYrd6TvFGP6uf+0z65w2Z6oOttIDdasI4zzN5WaNY2Lt4
YKkhj6XC5t9JuhHGSmdPjAGNRXHEWZb0g9koemInGBF4QcZctRY2uimHp23cAHku
ZaISJJHMbpmOSVdyR6A8Bo3OyqsOgwunlWZFsmCBISKCyxLUvO8SdXhmHK54GQaD
1Czf1VUBa4aeynVLEUEdbjsrg/Aj/8ZMcMn3uDlA5YSSd0GvDJr2VDX8cGiC8tD0
tOkcfw2kAoySA7f4AvtelUwx5qHtCT++dpqnn+qIb1WhN2rZJtgzn2RmpLsQGnLV
YOjy8h9PiniGmtpL+qwqnFsmafHh3PUHiS6dyez0dmShHMoFuhNKz2dJ0buMMYl9
LHCLGWBNYU8NE30w6JpONGv9mT6oJT6tYp8Fs99lJhgeJE66xztUe/whqFIqoHzb
xYyF0AowP2YwGEA4VWWUu8GcVm61MMf7VQiYaD0m8Qdwl0/yefKfv9RLgRzd2TzW
q5Z6Vtyld/q0/H4e1sVjczmtS587HxvLGhLyx3G1LzI+HoBd3jOWzfXXMGb/k6Qg
GWPkyGb8sKODASJxgR3NHOmXfnCO6uR9/m1wO6RZHwMIoUtqUGlSH808hRuPT//i
880fw8d23sUsE2BD/BHJOjvZuRnqwSsw24Pq//qyZESsMdX7VeMQoH7d9dNfi+V/
0UaEwE+6OdqhtJe6cmnkg7QD/SvvjJ/GXHOBaPlA5sHk4+35pk+keE1EEcYLr2p3
sC8Ts6Z8J3V5jJH//uroBSW3RcaPwfGeRC4GUIE8bGsscCq3cSO9kQFKMiOeaz9C
oLCbZyLO1ybhHH8FK+5pCGE+JjX2jiWTNAH1bDJxmWXurfJYX+W/wuh+t+t9R/yy
DhyvD28uWysvkbZvUE3MoFHafnhnEWK0Rykri3rY+iVLgmuS4p2ah0+M57OkqKnh
gbzOD1GzlhEFrPK0NlECI24lopNoBnUyrMoxkB7zY+NgGn5eLdCZdzgqJbRSaQA0
z1sEaxkN871RaGnFLNLto1riNEptlRYht2eE9Dns6FlqzggwXsX/5gEz5opMxH/Y
3fmDb4ovtm4YydeYE9hHL4XaB6PCU74bqT/K3Y8NPTIptPNlvAJL+5AHxZXAAjo2
GVPBUjLoVhDSTx+kjldhQbKrUMbOYlpoG18odRD7XTwfokj7GpwgJsPJMYeCa/OS
YPXoqa7wP6R2z0fGm07ytNi5Z00y67FEur9h9TdnrQ2/49tZG0hk1XHJ6LEGyfpX
oRK8Kdz30qQyjyFACIvdBaxtupMzQWpfu17JAgucArvwKgbeNFvT4vMFw0t21S17
4T4/I5nYhkR00vZgVkgEfBHd1BlDXp6e4CGf8DBtYLZRKYtfJ40OP+sJ25SukUdV
IfzIQ7DjxNrtyfB3XbuVMI85LGdheaM9HVTrSs3+JJaYYl13Ox7Jlr51rcwzirgP
joSOLDKjeVsEIgawZYcsrNeAnlnX9HwTgFyzx0Axiw4MUe9X6b5aHOq2tFK/9Bjm
jIexAtuH7wp7ALgshDLbtc/3qTKR6bvracHla56xvEYHWLLHtyhJbIwZlofupMj9
5/6pEyxxkftmVD+C53I+w9IeBQjvAOgMew4i2/P97p2+azyJzB7s0k17jLWmj1p1
POgX+C2REjWcEnr+Ieeox9dsPnG79qgt1O/gJBmo25aB47RgAqh1lNt8/hvCvbeV
ppEgBwS2enaCrYM7V6qWkZTgvuhhrt+02Va9pGFQ57i8ziv8fpI+xLECAJXPNCFI
sHoNqlG3b0K1BNChq7leZ8MZtUeTsk73I/xpo4RUyYhMwj0y3QFNJpa43CgqiBxq
32LKVjXTGn4QOEbLvCoJMYuMyC1ilzMkZxhJXW1cOS+Q6Vz1dcjbzwTQ/5oQNVQi
ym6PQvp15aig8H1KWG2fw6n0H4MAGl2YGqsC80faZwTyprwVeuIJjMgVnV7XRt2s
vg+fxjv5FO9VO4WDIZnws1HPTjduxIXWHW/4ny+zjmVD6PZX85cNekLmgDLvqTuc
6IRgfBknxaXjSRth52Cl3KNoxrkVxNyVDMx0TdrpLtSfm92kCHprSuTVdk9EZyDW
z4mb2NtTnauudSuBmt4Yu6LtJmruggMhfhaRigc2ATb5xs9aTLyX3sLkVeZ0XJkS
y6O4b4gOjx7kcce6DRV7u4G/+WJLHToEo9wGqOYfU72nE3Moc5Ela7QHuUzRfe/d
5MdpBMd7PDrbYjRKYQC69BQo3t0op97exNTDHoOSdGeuFufeK9lH+164SB9zDgu8
SoZaDX7qvfqidCrA/GGOr4XZzEu0n7gAU1ozC5i9n9nRG5621EHNgEUQ3bx8hOKn
mXI3mmYFiEGOukwcMMIQ3B+l7A9iwxzkUo3BUCa+DVrcdchttdFp+dsIWPZkJ3u7
tK3y8CRt8ANNCW3gikzKZE1z5Rhil1MhkNoUIi0Y/11uDJKTYJpT7HyOms/eDR7+
y6PsWp2JnFpUhbuR7wIZy66OJ4GP4PA9xaZJ2Ht8gM2C4NB/GoiVLwrfu9OWa2Vy
JScVjy7YI/pfVUpBbRpqBSdQKxNV7RUbWfx3+WoHy4w8USE4nfllEueQqc9q0DaG
YV9QycjpBw0P+OGXiqW1waCBCXc0tBB2+CNSShZL/AZJ33Qm7L4VllXXU7HvjeYK
qMKkRiPB2S7i/RV3XemGaoU86NcQop3JZdkEtCEcub9Lac+D9zvhOK1gToMNFtwn
N04Y46r5AMJyJNgYwmeD5ii/qJo6oNEhsXKe9R+GD5vtM3knTXvsUhAYHunRAYm1
RB8KdQU5ZzwEHahvF//fVXwUGQrRCEzHAR/YOPKwHiIpefge5hD/xCG0o+JolTCX
WmuMaO9vVyt4BE4wUkgKN9873trWQ/Dayp3UW+EefGg8TYjs0BWMD8Wt/vKjq6MR
0LbszfktK93jNz8bCOMvflk0WzAHu/XmFpLercbaEDLiUovrS49WodBnJLhSK2RT
sfUxy9HbPo2zDevK5Zb51Lm4aN8Kta6yHeiZA80EMi/njj5xlyWTSeBU9ZlM1hRz
rd5GRrL/Wuhyu0zia9dUtKtph3cfQmVuhTYLAXTPVBSKrMCvWmMGhY3DFgOyQ1R5
exVeFWIiXOcleiQEnTB9AG99A3qyyxivNyCR0TvqtN0n4/eFzHv9+kQIVIY9onpo
fcsXVJb7cFqrBfab4NNeyXc/+wgsHz17a+qhhmkfp94Uamp4FhoSbJdln+SerKyt
67U/TXrNKShTESTr3iBpdVtWIuWzaq1puR6t8vvrmVWWCgg2Df0Myz9gT5o3Az/K
P0oADCzuFYRwfg9uJ776uOiLx8GBR95fShwaA+5jaZS5ldQL8N46WwG/6fpgY+P3
6ur7b+rXD+70eQgTP7usrQeiuvNqcs9mBB07QSA++3AeMakOtq2x0Qz9pMqsfHj5
PTiaMUViwQFyJZliF3lg7Vg5FmGVlRcxfkFwoFhCIag8faZpjCKNwttdnOzTAfEp
qLPOjmrAogmy2WtJAmK2xxCyXM8OahWZVV6ZjsPWq0/QFy/nP9mmG5GgVIzvSx4u
kr4ynLy738DXPgDy50ONylx/nb0uK+h6VWA8eVR/15ricr3dGZa6Y56EtHQ2OgEx
qGX6tpfP6p7zR/oqWoKHh1xCvWmDRPEwEAJI1JVVqEFdyg2YcGm42Gd8YuO4sCeq
m7QmDxBUw70ldGjXXpjbN+3Y7ubueI6ukQ3eXmX1UkMKetRcaj6GVoVzSbdE/swB
fLCVeRfmGNE5gId0qD9rL+kEX/OfGf0Z0Ba+V6eZUsxnv2wj6kdCNOH89nmcFCp9
M5kGAPevDDNzRMiE/ZIzelCE31CK5Y9++FsnPc7uikGbzUphqs06v4e8XuxE3UzZ
Cr8a3GdwCDQUPyPxy8K0k/bYFQou9ge2+5BGBFMog+eo7uGNOulKnVWTt+DcoqmU
Ah+O67Dc7gkjx6M1uEN3YPnqmYyRQDiI7kBonM4sYLxyzRkmk307dEfdVfUu6sG6
2GGth15DWQxHMirpqhpQFQvGTwOjicLWOTmFBIkiKdzxHT5StAPHV9U2w2Sxf378
8nEH0+WXNS86OCci+NxZZy0wq1cba3Ge6JnvRHByTx+aSUTAP78nTWTNWIzJbgEc
xukau+wNGPXW0b5EhY8ETdOhf3ytKp+t08zb8QInXut+QBJqGFMP8szwAuHRkVOj
y6FNk8fL4Pe9sAEJhSQRqpy6j8myjzJK4sfIctYjfbwSZSDs1rslzrI5kLkKrk3x
42tWUulWCLKIxgISvRh9cbJgzv1qYyk+cSAsB0MhfnQMdDjgbTnS8EdP8Dl4CDIO
OFleR4FqVJgT5Ka/Lc0VP32l/lUB8uo1LT6Y4qXyTuO9vTLO3pl8h+7/aWWXNscl
HB969TLQce4KaTnln9qGENhnYGotHYT+BEaVbuCaVsYIlzYNUZMtd3bR5htO6QF3
jlSBNKY2IXMxzN9ZXN0vV4kIGdL8ebTQYssQI8y4NzsDmjanstOqQRRIh5SAmPgU
lY6xn5tIv9kfRkhrt/Aykt53lv3eVWRGSqf7WSewvkTBQ9XspKqilpX08Y/+Ai+j
nWPrU/Gn8OVmW5Z+Fq9K3T3fGBT3DR3csf5CLdryUse5TlQIZdlCUNddrZ05dqkm
iFJnZF+Yn5adu0K3vhsPu9OoEojW8S4Xi3bEsJgHBvoEj9rQI6FNgfa3chzXuff5
IXF+FT0D2I3mYqzBvVEqItSn8V0qNW3olATlJGCSWlJaq9WSeYMB29Z86Sk6kyv8
DVHlUdr5Aky63XfDaRrXv6rIC9ELw62Utt4JumxTbmuBA2c6TT+JwJXq/Df4Pyd/
2HELBZ5rtItp3OBOpDYPKtS8jlTr8hCeXjDwsuOYSvsTpBeCuvYpm9RWjM4EahYl
pKTMk6ZNj+4v/4LLbfHLkgqUfz+VphlC7jKKh/19Hiqif9mAAgmxyYn2nuCLyhMA
czmAlEMkeniUZkxfocF9imDHko1f6x8uFl144m7wDcAsica/0750ccFhE/Wl5Xh6
m+qaz3ZUhLl7sRIMpqsbDTI+dl90TIYKBnbgDgD87CqIxtuaE8963iGnEVNw9Z9M
IxF0ZkVfAN1hry9tvBrzOsyWgXXIX41Tlh3aj4Ehje/x76saEQ1MwSMKevIf2PO/
vA9SJvJ9jeB9z/bdI312abyl/pxiRQ7mGSwKNRB6rLRRUuUfMRHlqmDO5ViuL/n8
vxXPl41bhvK/sdk0Ei0/nZ2BOcf8OuRgv+HTNxFbwNgLJB84NaptASsC3Qt61ZLy
BxGG1BX9+pNNen8Sbtpmabe8iOwl97sJJZnNVDL7YBXo1lUE8+nUd/7IAgd1048E
rO7gjw9ivZPVzH94XQB9mD45gaHsXnu3LXl5NfKjBP/wF432eT6wrhOvQ02/u7bZ
5Oglomh6qwwXEcfN2H+XBb2n2GF1Qk6MgFra+m/VzMaIF8Z0Lj/q+LqQ6Q4aYSMo
FBH3Bh8zCChylV8bUvbqZV+w6bY+iJQcNEINxuDkzL8+oJsM1V/PZMAf9gSwPoyk
320E7O6IaO74rTjMg41ENS1JepyYXQBqdzRSdiDov1fuWWPmUcoVtEAkw3sY5Mdg
WuUcUNJ5xUiyEAchbCDZO3mOdSQKEl9eBzdDJypxNSyxZVCfHzY+ethWBDrkSo1o
e2HeiHaLQNz9HNT3CUjKzW6lIsoZrl9A6aLMViFiCLOKXp+hN8qBn34VNqg4KQeE
nWTQn3k9q6gcC/29wccRk2eLFK2ls1uUSbxdlZkF6bRwS6ZX1JBKmOmnGlsvfRNF
a9cf+rV+ApFM2cV1HaEapzz5KH7ia6XjZjODVoPuI7o8WmdWWOjySbUlsHNZqwnU
vRkt37ZZpQuTJZnTiRvHGphp24ZBeOBq3zqCdlO7mfZr4dJwDF+cPikMww+da7DV
onMVttglREIOpRKGB2se0x1me3QwTLyByrHrRaEKhVIoH0cbs5rWI35cPANtmS4G
/K1sIQkV6QjrX7q+bPxI8Dfbb2pKQxsv8aod/V7FJNLbEz0aGprpa+l8WJaFbTr1
pT487MEw7qLKlqJZLCWOmLYd2PLOEpRI9Rcwsh9gcNsdpLuhbrTrWKFe3bJFH56K
wE4Hgoge6rJ2MkxIerzhnYd2Ox4VwGqRo+Rts3nKzHfxPM7my7CccpzZFIVErd0N
AdP8wcEQIIqmxKcwXn92+5kVw5Nk6C8ySpE76CI4ReJk2eoQ3PgzWBxUfj+irygX
dlE31inUUVEHYxq9U//PU8XOUx0uLLzfuOEcjXw/j2bjzNx5xcM28s5FKdq6qZm7
HlAErHFUpxiaAKIAhmDHONezoN8hZOb+5CfqZUtMptGPGLfsrOwotpa1OxPIWknt
VPMzehFsxkxS9q/wHKDASpSUAT/YMZC2IkfuY/MJW1x+5HueMiAEU0eWI8390EqQ
XKmwQqMfcCSXB9aIsMKXKz3NJIyvrsA4NCN2YygUd0Uk0A+aIe/IjMCF8NUoDBcK
m6J5Y3vef2ZJ5fG0hqmoVE6JxGon8XQwo1Auus8CyknRnbbv2y5/gm27/kc49i3S
kWMw/7OJQF5iTDlpfwNWSz/Q15btOEyQKgxRb0+Cj5nHpl5lTzyWrn2SrypfwJsN
jZNWtIE6mzOdQ33yvCRFJ1JnFoGxiYckpUp1phSJAmw+IfKzOfpAqS9c4AmhuKnV
zjaePksmrk3adEwIk2fwKd5rDSOd2/5dBZVrFtCgZPRflia/S3AOpZh738g7ckiH
/lfKzZSl/wjvwuKmeauysWe89AHNO17rLtuwhxG/nSfU+U7eLI18P/q5LfoASv4u
YjEReNGCjIZn0Q5uHZSh8rsyn441hmCftByuHUVbHw0UvZpR6MV9i3seNV4FFbDt
WZMtg+cjs92bviP5TGvcmYHsoQGlGo94pHZCPW2Z3iIJs9cZUAoRvt8Ukhqvfswh
Ckt008vuyIcgMsIc163pS/ZgHDaqZJrGyNUPQPSAqys1K5H4tl3cmagA0c1+vyMD
teJPiuer9sLzX5i05cq28/IUVYWgwNTfPZ1BA6PmzNyiqviJyplaL1OEZNa/N1AV
garv6EXuI0Ec8RBh3HVZWiCgymyl8b6JkO8ylJwkXSFLWoI8yX2PhlHaIBY0KCkt
N/2pE9KIBH96L72qLk7fqY1tCSWszVFBqvBaBqmhwQGBboComCo1+Bc5qCp2v5BG
/UFymGYAhQezdPu1bXAHpaakgpiXm/mrKMnOnAj2xazqxLiXllxLKN7ZPYcAzev5
cgy/TRCbABOx2K3OKT630A/8lWr08KxpsjI0JNLsVx6r2PqqGyrxokeulPaL0PvB
Tf8uZTYCo4I0C+W2SeQ+d6a6rUFhBcxIvpRLV5940UL8sOuzQ934jj6mIsny9oUu
hFVYEVDokaXhgmzs190Wj6U26yWwvisctYoW3elgO4g2jG+nFYu1heDHUwY6BEV3
73an0aHy6Sm+247Qtd/VXCn8ssq7caxM9XNOl4P+Zsvz+B1QGEyVzEvKFUjt6+eN
zJKKpNGOKJ3roTlDxmfgDEJH1owQGUogABmpsD1lORp8YebwIqXkXRwCVWpvhD9p
lKmh8xZvwqNSo60TIIZv8YznQBNvu0/E4eqGlE5/Rn0dm4hoQYeya6Xd05Wi47z9
XYIUm1XhOxdhD5DEvrn864T+5acAbI6AbNnvYEgST8DF/u/B+3/mV6KkOH9ie4S/
Hfxj4NXiLHm8q10C4EUYcdugz/fbFygV9YVwTUNHKONk9VCIZeoiymNLPOkhbpma
FeIJtTyV0h/WLNHn92fUEg/JoE2ajfTSE1ZdFLOfZVbNrYyy8xFRb/oNmkh4n/jX
G+wFsUZrlq6itq9YHvsQ6Bomzhgj/Mml/JQFeaeQtTbsSTBeEDIvaJ5yOegpF7LW
PMkQ/EkMuwIJ3MN7JCykhTw2NBamLyOBuzlXmx55UBBLbvw5xsYXwBp7r+KuGGbB
ee4/jWrr73FEs4XHbKSSZJ0tcJnqLgkW5VItEWlgUwFa9+ZY8jyOhoOW1Wp/Wnm/
e19p3FH4nhWnbnB3BmzbQCjoQqUF6Mxaj2s94wxV4q0xXbBJgwzD5L1cha02QSrV
VtLi9EECqDaXwq7pB9A8HiMG7Tf4by6QSPOeta+7blSleWIchAC11dJdLNy99VV1
IEyCXA2IW45NxZ1eu/+yY6TdvZO7qkF2PRmR9nR5cN8ItOPAcpgHvVVXXrJqFlgF
TgoalvOxICWKmB48LgP2Btd6bl1HyjLecgXHNttysZ+3xTZf1Xm0B5tm3lHnHL5e
SDsAgzMiS5h1mrKafRW4hGVDtYUO2c+DRnLoxKKkWqAqHWNCYljDASKm5HR76yRX
Nhwo/9iyHRTwvHhFnQVNdzu7B7G0cFswIn5s0YIpTppmW3CllIx8FnDm024U0fBN
QzQeXzszL/slDGgefLsXo54Gib5anU1xAn8+YM9KyzQ0vtHB831BEesOIiXyqwL3
Kgxy7QbihTtg+Ki3ks6z2lI7cyIh4NTFIxtpIpVcEIsmt+g282TKL8APFFE5iRK6
0g0qwVbzOcD+3MMiTW0IVYN6UMElvQdUu1mLP+6kE6DJSeWcfCVfBYygpxCfK/9Q
gX7BesXLUQnQGtyedVhW8rAUnWoE6bSG40CZ+tQEUglwavQ8eAhtO+n5ad3o5b+v
VKSlx0VOz2+x+YitC6P9Wvyrai8YJu1M1Nv06OjuwKqMAvqR29bJDLX9NC9W+4RO
ttOwAud+aCN7LhWoBuiEqglugrFpdnBZ7TJyB6P1gyjecCZ64pETN+ESJcxMqUeJ
ZRZV49Zilo/UFnjXO/kXzi+yYtH1HFECVCDhrPN8XQ7qqrYtksXkAKFiUDRiUDV7
EbYgtnBox5REPKoBrTb+QRF70BqCQejno95yN6PvOu9fSET3AvkZsw93xqVqXGp3
FN3SHflcIElg8PDKbvWzQCehRRA1GXH4Xg/Dk/3PJ4t/xNo3Sc6H794CZx3jEmQ5
JT0uXIfe1rW/XBWOklWevY9QtL41QfNhVtYezjuD3RrXc1/tJppCtrmKghlHCTWz
dRdE73rlf3djn0hLGp4i9WX10iB0FR9S8Qz/CeYrqCN+qB6TiGCg6oAoL8NfgMtF
23t0ZN0t9qWlRg8kr+55EPhnVPhPlp88wPZOkfHSSHFkjXtR7P/ahgvIbm3bhp1M
RDXxe/+/e4od72Tti6PZbvIHEUVdDNcTNHP8IXiwdB6AhURb2eYqkvqQ1afdkvxn
xnQkYuJbXpxUQtjXhxaj3l4UIHs3I2IWPE5gPozrjN7CINjepdYKzkLAw3dQRXYh
WzpqaswM5iDmbCTVVh2BetYQ+PyBIt+4M+UumCfEUA6Iw28dRFA60pChwnJPX1XV
zsVsPhvi7VyyKKDMdnbTSvnyl07TR1WmfAbMYWXgsawy13Pm05vXhM1Zqe7ji+YV
dLX23bwKhGA7bwfLzQ/Is7NjRdIl9IEyJ23e6IGYSBDeIuJLKUSwXHlXZV/cbpmv
PyCjontwiW3Yrpz9fMbibmqcrOPv1hjRV8BoQxpC5yBUyzZD50zG595iELocFzS9
cXjNl1vWvW9BgJZTKnKGHHnsw2gC/ms+xlP0YGKCyjOe/IP3kSZvfwm8mY7bZ0pH
3ksaxG+4/pctmMlNAukdgsZONk47h4Zx1om1vtbXWDkwL6woevelklmgbXuQ6Hh/
fhgeYrCq2+z+fKVXZijKZX9YynK9BHKAkoJbN89SpNtqiNXjiVYae4GW3f1ku3r+
jiplTkJQnlystOEEdUAxdMDzItFiJlJCgRTms/bfMKJnrV5TukqSihxBN4R7PyPN
0G9IAeX0b3fqJnc2YIaUhc3PHwjVl7dFCv0LqR10flcYV//aMBMZiJ7EdbSofxLu
HgQ9hUzcs2abgUi5GZ/k0m8UK3P5AST4gnhRBc6ZTioQMq97rIHm9kMawfQfmBam
qNhHztrUODqNkOH6dTNxwK/9kOqTEEgh7a4sTkO31E2MK5FOo4snwdDH5eruV3NM
x5dgq8tYvZm7X+LkVLL8m1mUCBjzQ5BpvsYU+AMgB48QjchKFxqf8O9Dr2bkGHI8
KtRgSmY/k2zMvVSdr2wjgAE0J4UYd8MLs2I4+sVzrQBnl3yqWKxxNMoR1YRJwswh
SMzdSLont4WnvGDvzsDnSAsk6UTjfjHxD2ourCSdE4KbTikKyEvuXwa699HroUJQ
6aq5sTzcAUZumkfD+787tpLS71rZv/9rZqtWxr5FGABMgi5aQtEcQWHn8jhKDSTC
HOB7y6mbK3mkqEEs43fgf9CwaCFGvA2fWt/xTAEL8SCYZSAscp2euS2C+E/npogY
8TeDkVz4rkNLJv+JCDShWhmZxhFjeRPslstrXMZogBM1gdtKvbOCX/hayu89QDEw
8oseM29jOcwxpOU0QQ5P1qmasN3y6R0XZIL0k32HQKIFYNy8DyDTCBOYej2/s0hv
8TYSxoUlC0EP8RharJ1a0UR90uHfnzmvJlEqxx9TSoZKJNVzYSGycqQ7REjR6UBe
8e5rUhgPaknlL/sfnJ8/F7H8UtpG6l4EMHxRdMnWNuH+CVpRYorC74RsiNLZywZ/
41G+6PExZuOLCFh6OEL1PycMZiPEYX6sPn8/Khjg47sRK9gKw/vFceWfBw0Pr+/q
Qt8WLLU9lyxGEvg2OvohImFKnEAo6tpXQNzBemFLVEQFKaO2eWNO/Fyd9VORxG7x
ixpF3hrjCyac+2p0KmX0CDNEgNNLHy3x9TlgDUYywto4jZDB9p37LHLJtaCMJKVN
8QS2IBnFIg/WfOuNublblDzkwD//NsCuvLe5boGjSWSMdE0uHPjMMu4GY4ETMSK3
LICXlcwRa7FpVMXlAgwrUqYkcdxLDrb5utXA98vtDhabhpBNDLOrQlc876Yli2WI
BwpQU4ytAntraASP/3qaDRqXYnGCl6rGol1MA/2mSn3+HtB0gs/KMwx92XCQ54gW
UGmRTH48wVNa0CtKFGCRF4YDs1W6yXGB2PZ1/C713uDsJ2DJOMuBlXEhezyO+SaP
+bDya7glO2doOcarOCyGAYwZAPPg+aU4myiTg1wi4y86OT/e5A6zunFz6to0Lz2E
UnzT1jotExOLl8wD172sjia/kNXorqnMRQ4bkEonuV6zQSTtMKi8+Lk9Bm+Hu4I0
GnMOsIbvZATGKuyZx327FFnwCTZSPZYw1JO8QALOBztnesql0+q2G4xaaYpWIoVJ
ABqb2PbBVzm2EYtKT0rWr9lLhPG1iCvOCbwDZeOhk/KaLMyQdoXz0yIZo8u7Qtx8
lRUX7ttpNZxal+JgXLlA762fhDgTLIpxLY56YGAM5KbgKG9r4L0QdWtcLAawgdGM
bCYr6rN+SN9Espgb06jUwUDl2VqLY6B9EwKxiIh3zNs95V6aQy1E70NFj3CdpAip
xhs8dJPFY5m7cGySx/qzS40RPcZ97sa/+P8I+0Ta44f6k0H5Sp+WzVITRQgYm9lE
69NYUmeNWK+pde7tXp8eF5x/s0DmaBz+LE9gOGyJCMFFSwhqFt0pdmNx7JShr9Rd
76WFZKiIARSJdaqdjFeqO5DPRgYNYmhSEs1KFe/v7bWNp6xPMUseZuQqbxDurVdR
Qn1o2T/JnX/Dfdif22CPdiwYpQhdCClN/+BQUPqEiVxm0IRtP2i0MIAirXTOToVA
N0hDMqPDoTVReF2qjGl6NhlevWlEDwR8+hEPLFQr38jyApusE1rqxGNz8cNx+Wd9
zi6iBML5qMhktnbboBE6CXQXW8QZUdcKGYyB6gw9d9Ky/ew0gmYs2U2uHNPkZ3eB
bAodJjcUxix4FbvwapK3BisgiDEEE7RE8Iy5E3lRF8yrsdxOuusJsS4t4msWT/3k
BnvsOg8Y60HP95yGHIM9GW4Zg/IjGO5B4idbZguhRO4UF6cSIvqULXRrO2zCcu4H
+R2fhBhVXFtq2sw/96N/MYRPEEaq3PsWrvM1Z0fHpY38FySi5nDUzar9/DyXGhvo
7oYcEzrdpLUCRVkJ9OpklH4IHQRgwIWUWEna0Wyhrd0oHaxDJJbiK/WAI6+uL3r9
cTvInnwuWOcMRz7n5hMZ4vWivo9LV9VTQpvRLvHOA5heefYSCbXhLSqYdEafzFMd
1lluKec4ZRPVreoxUpAKzOdHIM0i/yzN5bMThjnEGC2sedjkkNVI/5KIG0sadafP
qywUTqXs5wnO+Cxq+H6S6+XiVOHWClt7OKeq4QZhmFxrH1QSlHgfP9G8Pnx6FCgF
ED21lUhfU9tg3dQl0pYmrW6QKxZ8QmpVtUweHjxSO/SpbQAMQSZtq4KYLoNR/AJq
lFLSdOhe/p3EPgpx6BJzPtyAV9by06Q+uhjxOysIFwH1UDTvU7UkxCPZRHGFY6fn
2UVBbehqibjSKLAAW7uNPsfKUOMyX2W8ZVG9dmyf433A0ktmWsIqdVkhCwut+mUr
oY2WtwB31KR9dBbUrZ29oWR0PUjUrlPBPAgBwXtlVlbsCfSn8ePc1zB2L3KU8cAE
rSZlw+7Pg9cxSKSe0EKdO2DUdXfqDuOdjOaJAkYfUBmBUHLo2wiFkpr6gufXHqC3
1oLCZrLH438bmBWPfehT/oSE41zk5/qlggD9YAKXm+rLCiKsDhZLZE2ASiGODED0
TmaRZamyN6PbKzVX4SO1tfByqCMYe0GgNlsH5TF6f8sxlUlEPeA5aevAv1hJUAo/
udev61crVyaGcksNnaseY6Vsmpu7EGKr78UzXJBacUA50VMg/o4Q8p2PNh9N78JS
8730R0y4hy1f4LAURP6Fyjmc7ehktmVdUNzF97sHzYHSWBOhG8XBRYYnKEje/VSR
3kqea1UtYpc+fRnBEeYt36c54DBmFkDe8r/8czqjv/E+EVjxyf9EVSAfNZlKnfVA
NVCXgt9em8sOU8AaZP46X79YY/77BNO/1jhu3aS6+YsLnDQ9eLswXxWfe14sd0yA
zEFVT4JtDfy4HDkqGQzYj2ek7VEEzgA0CPHDSzZ37Z+xsvF7yWwTsearSONMf76k
um4zuDixwfvm/OM0HftCAAzj15tnv41EX9OQgrapyUy7WSuODRb1wPfNIo89bv5m
Qq+zkO4BzVhY8SYYSayaItKMn5zxUlhNouKVjEbSelK6znGvt29EIZO+Q6ngWE1A
6p09WCJTC6qKAWvz9SNmk4mAH6nqbKDpImX6rGHN5J9P5lEZubflb8co3Q13+cmR
wB5LXhBKRqs/jOdghj3bqPzqtOKuvNULJcBIHxrD+brMmD8+P1t/S+vrtYxvoPQM
TasTaBg2oez//91RZ0aPWruhjIjbZIXHnUTSZLNv9xOUG/cGI5I8vDDzuOPqO/Lr
/l+/Zvo0OKoqUZyly5ZJzAx0eMG/r6cTSH7H/j5smj174snlkp+b5DeBtdeUIfYc
8YDNAx8wwoxD7SqlVQJPPm7w9iBtkwTOie5yMDXACDpGqj+RcOgRgiD65/DjmP/8
yXN/Ysz/QycZwiPevhMCiCH/xoe4i81HtiQ+yDo2xoEKRt2pG2iKXC/GLJa2owXX
nodqpItckaUb8/kcHgURAJ5ipMKfi0EQMWNU/4bgmkF/FUOFONbpHrtkjDUa968c
bVftggJyiH3e10EDvbcgipChBqOsY/s4gv2vjS5/2R8yaiUcHJRe8pIM+u80DejO
9LI2XDTz9t3pKqiHyLsAu5xFCZQp5vx1uGI/Hs5b4BODM8uvNebl1YPmGc9vdEBF
NcKvOTNV5lwMNFNe7GuEhDEsXOMtjmBro8dx9yg27H6i9Sd2fK8FzSvJ5B9IbEkt
/GtMtHNV+FwRQgpqmytaVwUMkhxl0skhXIypSWclXCuUGtV0cqfZ6GnWvnIILYd/
4B5rZ6qlUEAti/YlN3z/dHdv7ZJnggCBMfVmis4o0UKen5bvUnIHrJ5Sl7hrF4eB
qdofTUTdSymhKD+ia1D8KJzML7f0SUjeVnB/DOmIBmnhkK/gT+XHVnNXRyDG2qYH
W4n3BBOkv/z16bqFX7vltPeS+KXpiSRZ7ox79akN1ckEwFUw0Rkp1HeOlyCF23E3
9ylzIc01zmHmErkxHXpXqbnkv+TbWe9d1kwN0U/BgixEWHs7zo4J22VP3C/fP809
9A+X/ooMV9Qv52doa9dyR5/Q1FclneJ9+tq28Z7TvV2ntHtcQsBP+jTRGI+uBJEV
SsMM95O9WIO0IULfEE+gJrzoOHC1UtCtr9IOyu06KXGZ/kxIDtNb5OkUMPR83ybq
5b9mvF7uAn6NMOW4ANo2IJOxUIb3+qQVL50nBeI9lF0MCa37Ao6YikSm/DJpNS1/
cQ/Bbcverz4eYeSHzvpSq1aFs3K1yTTMlnuyyZ1Jp1vRu6LyZ5eWDqHbEyzRFltA
9PB1MIk2NxmZWGo24C9HEaLktYP7D44E4tmWk1/g5ds17crgI8pKcNzNzQpL2af3
ReJrTve8Gqmrp0WA8Q1naaggG2BMSaN8fC9Av/JMllr/Wvab5/tFUdLE0TmZWl1F
o72u1O7Ee0iEQ6yPcFAnjQrrY1HCzUZwadBa/BmE6wpok/jw4MUIaPr+0m/9yTAB
aSD4n0E70Ms5xxwQ2+dxDMCS7Q43mfh7DoM8uxCBwMxZAbumpmA60pxIqqmCiuF1
oUutmtWSmg35rWT7rPjf3dHduXYVDmSpXpf/Ahd/Xvrr5ZmzwoxPkKv8rVraM8qU
PNFe6k/pEnqU6Cn19aVXqFYDYz6ddRoZ7Ad50iSX5reERIpQr7qCLmmtDsulBhws
gtn177RFKTNI4Z+/OdSFBlLdnYXGmc9ywTt5i3S3H78FqabWwEXRp2aeFeManySj
Wmvu7QvM4kgOXCtB0DiSOf19V29i0TFoyRZKrFJTi0AgH0GjMDylpZqd+tLHfM5d
/g0p0jCvcPeGu7dKlbibxJBxIZBdsdNF0cb2Oy3SCjy5WWuIkCAVhxC73gH0dss5
0F21Fz57rfWtOAdFk8wnkAhvKVioDtQX3lSFGdg9JHGsXl7P9rTkwet9JaVsjN8M
YUxvLcn8BuePxBHpTHm0+rkwsv1J5quxt6Ejeaj7fzadZ/lpTv7rSC8nWqve9MF9
Ucih8SyIDTriSQK3qiM5iDU9C7bRfjoxVncWDPJHmroXqTAZsh14BVPDQQ94KIrt
lhbj7uoWxWkJZIhKp/PB1keceB9yEgs934HWiEjWYchkVQaXFsc04ssEvUbKH+c/
XOpoZBnNzcVaXiBo+9RB3TOlHcQTvONF/QvNoIr+n23RF4fxW6mWQUD7dtj7FzxB
JeR2FSvGW8zyvNYR9gn2mDteaweOplm1e/o+8ZrWEtWtlXmjakDz/3EcZok0e9Gh
jiVbh2RwhrhOR1f2JsuH5rj4KEUbLPSg4qMfDzt4yW3oJceekwiT1q3jvWWsjAiM
4mkAt4pgqLadDfXaTJELMmJsXAUamH4OkT/9hFNrHwXqehZaONu3Fc7VrmUzu9mN
pDHhuIB85bN4gtrexN3d2YIV/thJoH+uws/OIEkGEKnu1cfJNxMRIi7xPDzaZmVT
ykpWEOujdxvBOiMo6sH1IRXUqbBMDHiVoQEQ80b1zrBa7vQI9kCaD81OuJ80BtKY
GxnqrisGRCd4GYNVJbo59sXqaS1EUBvN+OAClebKXl/+G/FV7gSPB1+OsFgmokKm
iZnIsMzPldfYuro7uD34d06ihr0zMeihZzvsYeMwkMJvs3r+gWCj8wms8m8t1jjy
lXH0GjjdZfJULO2aD/2xzO7bRYpZvavOV6WOhRjiwMiTuFsABPO1mi9pXwE9brUc
iapGrXt3HYvFb6yLgbmdjP7tDj8HVAnIwLG5/1el4M5kqJ3NXYuQznlrvy8xhMGd
ZpLDdQTADaeW3zqe8sfAuAMyWpMSllXLG0+dNaHTjHJy2/WM7OADJaWXtry5snNd
FdSIh282brcRKoyoEIQOlZ9WtGFrG89DHw9YTJxt0EPI1c2y0yxvcvrbr65JduNk
PaN6vZTyMtJUeUeTZ9hMuBsi0sKmRdfwZkPkZigQprE1nzDf5WoJGSWUPmGfGDh+
20Xm8JDC5MDGa1+7dWbal/mBwvhzqd/6donOSAMTjKBHcdzNDE4Yqc5piB1Tqxy1
l4QZYuA6iv5GgXvNQ5KmKDBhLSE6YFBaC9yE4LTrz0D6nwPb+ieWq/u5eDwblvTH
F5TaaDhd21Pm5M5TJ7PPGmWLsOppa3sK9nX8sNtr7xQlEuEj6l61DYvoYUB2gM9j
SdAy1Fs+Sbd5onPH+ZHOeLF0goi0dXgbrTfpu49AvKHWbJyk7stfCQxhJuTmmwJN
g1RgpBVpBbckKMKB1IBmXdzvhC3vZKpQn6ZgrBNQT3iXegjo4VThrEdtj/pFpyKr
q9+uinhiHflR18Ez2122y/xmD6r37rGNShpth1fbDikk3acZGCuvjZpH3zvw7uus
ESiyXIiYnVSaICJcD1BDN26JG8/t4QGgi6ju3JpmNwiMAf9mnoMPNHYA3iltvgIL
EjnquVCNQc10ZqHuSPIuMOXdrbfIQ+o9UNqZq7/HycRTmj93aEWip5zvF1NGebzT
8BsUBK0cRnkf/UJwDqbvdlyU0+IMWoIbkoJQkOxJ9Hj/4M5VhvE1BSvaX7c7010e
mXKbPHAOsQ94wD5CRMriHlTbGnn6Qj8Y1BTUGPZgM7bbnObwFfeln6xII9qS3gH1
kFVgfGibb0Ig0bzoy1uVdDWsGjIDAUa219HyIF3tG4kFHss9FarRZVRfQ61H48OP
O4hmJXmqZ7UL5qe5zimfqp7FWS1aHxHR5H488zi8MmFLUve5IghNqYkzj6Tcz8N6
OReyWhbd/TkiwcH/H3T3cwhU74wHqKKElTzPJmNEW1TYks2jqQMBv1lFMf2mKGvO
OeqZnpTPbaQFynPcJi/xpZvEBuIlgnSt4UWhVC9j9FiRoSNjZ+1ZPERtZFJ0bTtB
aWX5t5XcI9YtQPLnBhFkrmcM59WjjWVO6nlEzP69zNC7O19cR/RQ8fM5u6U1O0Ip
WX8caKcQfL3aAV5QsXrGakqIQXmhoaJ1mCGFpPvoB2ytnp23uLTo0XVpeCK1dggB
cZTUjG6w6CGtn9/5WFzCv2h6cWiAIgfomv5b+beOeFPLceszk50Bf8xAtxbIlBFR
naZTfAmMKf9l7csk4KmK9vv99YjXcC7cMMSeqwy6Olbzeqn7uWkMmyJQTlbN1Nl7
C+GZtJGHnB9iWfsZxytininz0nfNbSZgFMmdcmsx07NzDYTNZ2G5GWHN1jaPFCAA
lC6lMDOFcctFnV56MKqUxiK+xQOb8Akk8+Kqy311atn2afU6vwvW+BPZznhUsKC+
9KYmvbLvOpv1vGxNjaECC2Pc0HlU3hRzvjrivxq91nnXroo9SHqP9VP4MSIk4uJR
YLvzpUabizVKfXQWD8PHfHQHoGubJCSaGWjxFNXVW0B5naKF3hckVs9rTBDAjLf6
gxm20F9KaA8GfFRcB8Wt8tbCzyrCDfpd8UvU19/pkaCXe+RgPu+w3gq9LfTcREg8
F1EC+yVsXe/iwDaXcdJ2zR1It0PHyMqtkwQtqUMFDJsoHEdPHhqk1gyttehHYDP6
pAlLKVxEZB0ZHZRqGzv5fhAXyNkElNxGQ0c7v9aXX+UtmEbSVAxNd1KK/KeK1KTe
BWmgqwPxqEoFUl2Htok1L/kvzDgVihjS2NuRnnfBLsmDgg4rKUnz0f52RqBI5jBe
/eBk0CYow1yizeOweOwarkvH/6RsYXhy4YcFaCA8gi6qc2ym0qnw6YS2sSZsHqFB
caNhcV5YscBxDXwFiI9gki6au3FGHhS0pqv4uud8pnFa/w2jSrC/GrJ1CdTW7xPa
AV5SAg5OSeUj15tqRSFmLdHvCUnNgRgA7jl9OVxkKsuKCVsetWwXnfOGSeoB7E9D
0KgSlbY0dhuqhmPWuTPgrsbc95q4PyitrZepRtYPhyW+XzLddZO7KDJtpp1W4hEK
iAghEFEeP2EiPzEQG9eK41ciKtn2jBsKQbLzT+mA5oqwGxF1sjlqnKEbn9KIdcwY
rLQ+UGU/IL1Qr/8kmk7jSVdXqG0XELA3083wMQWw1+QcKcrt1utTCeNUON3/Z9nu
mYlR9Ap/Ej+rXerNb1vo71QWgZ7lTUELGi9+AgLWr2EWS6/vNrfElfDpKOHo8wXG
bbDB4rDRC0swr93WS9mlgWord2tSzB7nW27qA0V6qKNtJHqXM1+7KBHxTXvIsH1L
FvqGBsXCRnVZHS02JV/EKSTVA+KLzvbbFWGwjdnMwQYqYOZ3oIPDjFGqbWP5G60H
yZAgfRAbpuIwhdcjxaQwUUlOGjRzpDRq9Nt9tPOckJHczqlhomcWJNikV2DNf4yJ
Ylb5WGRYxksYF8xMbVZDKAKaOfu8J8xW0dGKeCnQ26Kn2ALLsxvm8SY8kdy5pCsZ
RM5tjS+740egoCI1kVynjE0vpthK+ywWiZwlO1JW1XRfk3iFHckMBJDZVntvlhet
u4OiM3dII+oES0qjWgdE4IYCFb4IPf6KCaypdmUHLvGgO0OFyCjvnZiyX//Vl7FP
nh6eZHeh7WrndyswlUmebgPow4pFv2ZDJENNAMvOnv13lJogEQwO2JN10vxr9VUs
vXikk6bR+D5irB+p41u60A14toVZlVfgLft2yvcFXRHDxYF+Wfq8t4OsjugIh4eo
57gNoYGwPP3//9dJCHMRjZ6BSTykGh6fmsrBrEgW1dabIjTyNmeuZBdu2/pChk7A
eut9NUphw2jQNbT3iKhgpdW1DFrJO3TICr3TQap6cAJY/9G938xCG4X6aE05/2he
ro45cF7hQGhMu6LvkwLNBRoOLiTcMUep/u5cCZGZWZn4kcsQNikWai41sVFZTgfH
6KIB0m9mm9FKPrAZvvX2j2Q4xM6aK+El1ZB0Y3e8mEL+H/p13s4I+G6sIBYtLSu+
PZx7drHvMnkFSvEAebtaMFk+Dtre4KtzCP6z/GagE9+DcxZoPy0y/S5M90+Yodu/
kWruNHsCrUFvz+9VAhqoLg6adoNxQxy/x/v/bobvyip1vyeqB/IvmgZ7Cmr4psW3
CxPZ0byYnyU2ot3WCnZpdG94Og8Zt/ZMw/Dy69kyM5cm1WsUX5mOdpN9d9ltGh3P
HSjkC5rgboFIzu/isDHuIMYC3uviTQGRnXL6VhbCAIItpaZiXDmgbdS17pZmEAbf
Nrpjvjbd4Mw++a7CpdEK/hJHeRtWat0IIYUI8A3MVMUBmmYrnW4lDuGItbqHcsYt
evR8cN7C437Zv+q7olOI3veVBYnguU9vyCij6zL0hm5vXd0hw+LAHQ9L0MvfObBT
4IUU+a+3vplHZvQUK7eV8VfPgprSchOv08L6o7TUKwcIIR+m4vCj2wIbVgmOm6bZ
wGUJ425Kn+KR7/mvKao6wzR0ehoH7oUCMISy77PXoCYHxrelV94isePdYp9ssNyT
4AheM4kFg+0YCg4lQuazQfm7xV9NSXrw9aaQd8qs0iSftDmjBavpO4RAAGyNejtc
FVwB9BCfIRDJb8yPtphe2cmcspJD+oziw04r7K9j2NfEF6yIscJP9iV1PSWfw5xN
feq1199B16SR8a6Urvg3knbtD0RufIMMNa64n0rHryUGVoPDJTpePCgUlA8HtHxS
IX08C3AODM8OgpZBfeBmJLRli3GfzLMcj2gPN5o1AZoVMHKJVCLpJMffs90TJYJR
l6T/T/2X4HjKs7wpQgMshxzrlihrdKsI3Oo2vzhZC/+SGS2KZhsnsz2e9HtrBc6B
lSlmksEb5aL1WaXJ7zk0zRKN8JNPid6NG5qBWwa3pjBCOi2HehTmngtNAeZoPQfA
PnC6fZFbwk7qfOcjFEcrQUh5uCpSOlYoeEtVSqycJFdPH53Dm8QmqIzUEl1uSRAx
A9Zc+28KKfS1iyxJRXPz5mRrBC3DbmOY7yfeVGZ5RWEVcStuRfK3VvWY+vc3+8F5
22Q2ixW7J+o01Tqk033PYl5oGzFvxA6haiwQUFFqEKc0lwp6pmxMzcVLcnMiMRHi
5/zvlNgL/uXIjpyNonmR8OfDZZ4J1HKzbQ9gzDruh6T8UFCEI6Z5VeZcGdhlpwDV
BjbofeL781EBItIFoUy7aDSfYaPjZsFmOPpSmbDjzf0WpjSn2xo8mtXsYJSdjhJ9
JPPZ3rVMxtadyhrWvp6tzXQ8GLio+CnxCJY8AgubvtOsNHd/foa6LXAwbrimtpH/
YqgCJtF6tg6VwuikH+UvUmw6hWAVlMQhNV+D/ivgqj3xwTHx7YKIkiwm2ElMyaas
DkgI0pMgeJL52n6RXyN0f2j7j2cUJFp4sS/OoleeDZua2Tad9KbABkFzVyJ8OuUR
fy+4FJRvaTkSoFLLu/01FV4+u+S9NlAVYM79RZXKOUjNBgVesya1tUMGcWWFk0JR
pZQu7bUJ79E9l0OOca6uFICfBCqUwOOmO2ROSlIiGpeTlRuux64JeArh122sTOBn
rk3zOnpOprTLfoeLY09oRkbAEPDbANO6gD0HVY7xQQLKJW4WBwEGfGgbq80vO9Ok
8kFSPLPzs6elQdxMn0W4A/puwiLI+Lurvnhf90SLxW0aDM9yW93ru8kFDi9NROgL
9TW8EI4WdqsHlG2WltaEJ7HjSideYj5q8xSRh8XO3JoaR+WrwBQPqkRQVPOmS9Ad
8twunoWAx35XdS+nmS1ViCTsgmYm+hcry+6xLWw5gVg2XFgLvyuglD4OEWw2gevj
t8M6s/l9KI1x7CMG4xAiZur9fNti9OTLyLgGTRnF6m6CmwMEUiMS8ZZmuqyUceXo
Ts7ov92WxfOwGEEI6CNQXwV+mLE40Z9RERE1F4Oho/MVFmDzBxpicU0Dnk0n8DBN
dxLr+armu535nl2oufBkGJ8cmBcLUaw5dRhZtYcWj00JayiNcHpspVZ3/ewnUt6X
o5hwZ+GPrJugleyBputTtL9wnQPWNrmkecS3nW5m4YTS3mnj7vuDlCwNGDRFPBNi
rHbEh1jLfKG6KWqFsI7ivn1LGCOHpbkh6uCmNVfx5jd8zV0UAtwuVcaDsjL+kpC3
OoNAawbjuXlzFFlO+Fwn28Xm/FQsECqVZSOFAWKNemQgysvdFWPQ1EpqNL8EhTca
0Tnzn4c8UWDlsCeCRozwMNJlfebm9k6hs/WB2YgvBlWwrhC7e2KXH05bczoMMQsl
JjPMb/lI2FkrWS7ZCvygmXjnJ6VE0pyiySBa3wkwOGKgBLAam5Hk1DvHXMRD9X0n
PezN+gl+100OwxKLkqnb00VfiI4999Ats/Sc4enFdW+s/PnJcVa5knGkECnqSOp/
Sg7SRc9R3px07C6zBZMPeUym/jg9PXGN3fMuoFzyNzDVx9Gq5tlA7h0JVB+dAwqv
zlhjFylweLpMASewEkG8pNyl1BpiGqBZ7pu0btM13cWqURuUXFZIZSPEv2TLVTX7
99lTs5jzdjZimwTL7SXgZFQq10xRWAVP6EMjkeShqa19RYERCepfttWfQpO95nSz
QRD3dCbvik3pJUWR8wpBDm62hpkgtZfus5R4XYAjsLy98aVawDVaR450yLnfabep
I4/vNDm7gckd7Npn/gkfF90L3tHAFTfS6f6N6rBirG+tbbCCrDejviR5EjP81Hqe
GtngRMSWNbE0sPwEXKf62KtMUR2e+dnlBAUEcIIdsjT05t45LUV8LFMky6FV4RfS
XclcZahznsnPy+N68JksJUY2FmzXUZcODd9cl9xNFFQzzE5X0vJXhgifVtmk004H
x3zfEL7nRNvqIV77NZZ7TQHl20vxRi+RI5wwS8Vlo7936hhp44YSd2+jGS0xW5yu
E3J8yp34suKgtYoVWuAkb59hldUdvv2gwfbJFw/00xHjJNse/J9DlqphuNFQ1oQD
QWVOsjr0K7+LYCecPZnZRzt/UzBSLXvJOJvO/vZDldSr9zAHVvu7lTAGua5u5uxz
S9aLJaDqtieKwI8kfCuYtPuajumW+C8ydOulG5ZSpniT2NvoPU7WqDjQ8WMIyh/Y
7wDKol/3j6pdn8JAYHxfviqe3MRDlLP49SE7Ze9TmyYg0RhmLRJ8xNX9531rTXs+
oAmisQDiybWgmkqSaO1utbUH8ITw9HZ0FIquZJfXA8Xzl9Q3Kekd5uPxkZiVJBqQ
QOlpJzdjAd7A89PXYdySSXTacphjhYiovQmxbJXap+88KAcs9l9y7vmw5b81AD2B
mxep7pq0UptbkesI9xAaYQP4IgDhdcFV9ikRABWiMRL3kHIAi+zB136+zZm2bcwd
7fkeD+H1NfUgIE/EfwJi3E0gP1FMYJ9KngLwyvJf9wEDL072U9WssjP32Ofyqcp8
+xh3qAqjRVDik3gRw4ce4EBJa6FLPCLKNY10WVqE3aqrddQ7Lny0PgWtQz9vBmu5
pbgk22zUckRWV3N0nO2T4PpB85M1XArhwf9IurfLqDWPgB1fDcjJfRZ64F0LD+eO
E7Z1ouPC5egsTjzXyooHJCCZRWeAGvvPbZGUdV9y172JCcS/QRvNSyGQW6v6OMR7
pnzW+b6wKOjIUp6hdTXgHowMzrpsMINKZnUb+WgiOiBqcxLOF4OueA4WqGGHTOuY
VJzCsMQ674HS/uarJe7G7FaAczo0p3nceL6BR48dvFyOutkSJ0yLsJNKUaaQU3AA
L7WI2MP7tg/jRAsjkZgM9wYmRfUbd712WOcQmt8XZUhh93PL3rPq1I64CDClKkWE
jvrVQigHwC352J99iFA+EKZONrTPlmVD17ZBn+eyR/3QfsGsv7qgqiarlM12S88I
qkcMvAUmMDd2ba2G5l4W8MbeDa0fBMVeUhksEAsd8Nje0mlcJqtMUFAPXP25OQQy
B1OqvVAhl87cqK3ZDBqjGchYK+UEkUZvxop8w/t5pC8QYEbEJ7WA7m28qSDv8Vbo
Mgt5oUSIItgUh1bgNyGzOAvZWwG8Ca8qHqs2xbfA62aWR5L6zKERuIIhD3qbaGCd
Y8Q2ZKzevarGZplGixf1KtZRjFqy9B/6tI49ewbNyyreAkgxFIaUiGYo2T+zSOzv
U7iVu4d7wqXOkNjUb3pCWdAXuZ5PGyjBlsVxr7O/0T4AwjVP2lv+bCcf6QuAcIpf
vUI+jt8uw7cMKri9wBzuJOg6T8dCHdPKwbiCwEeXgV9W5sKaMasoEuKQ5NIsXh71
2MQNC7EZko+07uxY94K5cxS/YbR1YweNPrV/FXBf7xIguszaBZgv7Y/yRHv8USGo
Zr+rDfTtmYekfuuaRHZcPg/83kppJcKLXDUMCOsurcmCV3t2nDeu9czHkLYU+mpF
JPr9T0fZ07wxVC0Cwnj961kMAnniAEGORg8mohlPewhyWUiq4TA6t6EihrAs1nw4
6ovUOXgWah14vAfgcn2KHduYocruvv9nyh1kGVCDzhQxK7xQ8WlMzpPmzpZIjhSz
8b7VcNiEk0hN59jGJv5mwQrR0IQM2URiM44cI6IvX5U+FocALSi34d9ktQqtVtUv
mzH1zwgDkKo/0CiwC2RXeo2YibmheKXEdRQTg4itWR0fzqk0VUJWicp8Aqca0+AQ
nkQsZlUT6wgxzU/r8A3LetLF6KLRrEbXuUB3BflmXFOBpoHMxWzjW5ZdYDmCweAW
vuPkGvZVxqhejv3KOcaP29oUN9iYIX8sCOiMXOnMWmRjOBYDsgj8khDotS3n8sJQ
buFP0uP5o+BTKpsaM8nDaiqx8VyYCFyfFqf1juhPH1NDM1YZ+oCZY/bA9FX4PAe7
gax2INiuH6nC8e+vR5y/Ggs5hW1zQoSGDJkT6Evkby8wI9I6XsjzxuGqApVF8gHO
tCrbn7mFu8SQBndLQiQlzLGbUhuiehVHXKchQmHiQ3IGPyf5ubv8WmnL8IfbMemR
qYm2VzJuQaG6ly6Lpb4LHrLx+l5TUFkgPIxjXWxT7gTT7GDPfQJueu+auRybXabf
SSs3TTqxgvGEJeeqmWu/gDJH6VmMzEMlEw4juY1EWxZfsTI/guDAIPHxkaUv2qEr
kcSm7Y4fH+PWAuzX+bWMrluIyaTCrmRaMaxsmcjkooS64+aZ/UVCZU6cyX8XjLVn
Z10PQ2LRAOH1wmKBkWOd9kzinp9l8GVN0xtVdDpeV1NTn1wGuY4yZS6635z9xrBp
HN7QJtPkHWm1SZo0tq90RFV7TVns2TCX19nqXrmSDQNadygSxSGfEPrZ4RRGhwus
7Ax8ryRy0GY3QWRxo4IwMkTB0ixq0srulkBtnhFTHGmZTpWOY93PW7yp6vDSZdBI
PyPjTIVMR6mZ9eD3eoT0sK6rf7KKSFn3dGFe/UKgTEKMlVdtpJYpbWE4dvTfwgbk
lD6b9CJctYucYU8Tt8Qg5wDRrTgqPcaOxKT1m9PgaXP4NRbXbT4u4lTNw/yAmOi0
QiDwsFKTlZPt6XjNHFxWe0d8SZv52HewFnrtmVWHGmukt87+FaUV7Nc/K99cm0tU
DTp4L1fDI58spUQzfSk7LPee0/mxzv1v1ddl2HmVxsPW+92y9hkzzN3Oqfyfz1E0
8kbdbMrHela9hLUgBFN20Yn2t76plmIWNjzL9eGdea4N3ghwPefQr8fZlkNkpHQ9
Tc4wPpID3YM2Gq5s91BQbL64zXbzCFDABsV2+TcgSyyHk0vA5aOm7b+Clu/fn0Q2
AvD7YtJ0ZR1Qgn1i/vSSAO3KAmxo/ffi+o8scoEIxGryxMurMr4pz0VgW9e9FlSz
0cf2kREa5bYtGju+9Bw7pns4vDyI7/K9+UHnBB/rGkhf+ahNRO4I9EGp6NSXs1tJ
rBRh2yP9rqnh1JHPoWp55qG+SFBSnBkbEEWO26ChbuhZq2Wm2YI0mCr7AsVSZjsU
EPFR2amSXdV29yBQ8fJfI/zbFrTuq/yGxihGDOQgCvTHprXYhFAWsYcvoz9K5A4t
BR64shSPTBgPPDO4W5TTu/V4BtKzJKbFMJ0savPGHwoUC20J62/2ufbOoIRTprUp
+vTfYS2B9wPAdZBEE1TWRaIuqkUtcj9ox713fPuLPTiLM/G3ygJAsbz5Ffx7cJzy
7mLHg1iLlj74VAqzyIrryazI2xwFwVuL8o0/jOnhwF3Dmb0u1yfYLZBvrql5Ppv7
M6nHhCp+VLlFr02tCYo0edhLH6jjHNX4MwFQE2rZUZZ5mrSKFTeoiPrl6LSFeeF5
Ra6K/fzWo2pJJV3bimwn+s4H3X85nD0D+K9NaIk5LaYnqVhyJxucWJnfLCC1WF1E
ekzSIFLakDbP20DMMSGQKUfAh9tthnT3J2Jj6U94zzKj8EcGWJSfPnGr6m75SnN0
dOH3JglpmGYd9Srbwfn5Jz5hwhl3vysEmFJn+yj+p6XHaNmj0GCiM5s+rVS46bss
onYjvhQLpLnUtQ1DMSR4N9pk3UUPd6rIKasblG1eRUReTEsgpao3AExwJAt9AJtS
7nbGkw63C+KblGoN0QMqx+PuH1stuPKpeTD/6zMY7HybePUS10yiLDoRsPFnmdwg
AGjuWXLWJxZhkZMo6fgD5L5Elv5DoY0ci55JwMA84hzWDk58qS8ta2wdm0OxwFkN
h0/KXLR13kPrZNWCGdw/c7GEnuYrt9kDV5g3sbx76r/AZNr74pDn6YhuX22z5AuD
P3qhnUcRhI50j4Ii9RINHIIlClx073CEJSfweCw/0yT79Hlrihx+wTXIrR12W3Pk
dyAgKB6JRjYJ05eT/yFUflI3W5/Prbi0/wiOJK+kCYD9aPW/POSIL5WcSoz8clml
hAxlSsMNrUhsW5rxIGlewbiloYGu8WZgVmAl3OL45qkKP1AA4oEJPqgfkiGYc2TR
qKqf3xNTs9f2V51b99ekleg1+ErkpuRekjgOm6nKCgw3fiUDOnvhYHX9sVfKp/3M
IBzjWfYtosI/u0d6zrL6PO4ogiohWjIya5OHrJIgqmLKVr5vgMWz17dTcBuvq6jB
YD6Bwf+cxZSoxbU8JEvU9Xgr0vHjFTvATYQwc2UHigmqRXtlhr7GCmyMnD7kjMoy
r9rxwD8OKd4QkcOhRKBmtBrOkakCVfFhutWkSqCtJxeazv2bLv9j7gTIURx4Zj7a
fgbzKLiAHlJUH8fmevszO1E66AThB6ImTncMpB9WEiNKd4i13gVHUhXiVCStlkGG
z81Ou8DxAF7tCzPfV1wqliupFUqDK2rYj69PnO6Jabt8DlC4PE5nOmYtIeU80+ID
HzTP+TweSEN0sqN2M914r7TshezrtgGpP6iE7lOlLRvSxnQvrsbntw9uW3y10V8B
rE8ZH9aNODice/jBMrI62gf8nQT2yuG6JUnuT7pdYwumllpSB2wJqsI9QuagqOFD
zsf1qw+LHl3Nts0ooZmwx4OS1dCxqL4EaF9LhW6bZPDTlFDTmuOABIKL1bSrHS0L
8COsIkXJY2E0fhoS52EjEJB7LmxBbkTqEblc2AIG/ZMuEVRKwZ3lTsBXMQTuoQe2
ecN3ahuNzgNZno+jHc0oPcdHwnzuoFVBcleYhB673P8r7fJy1n4zdqTzwyUDXTGM
XQixfzk6ong1hC9YT8/Zkje+hxpWYvNKJZKjKrXrrrDEnXqL5kZjh10L2p2ouPCs
FfY0AlolS6S/WZ3rMMsTVsiyFSCnhR91TPTRl/5FYBRwJabzd8OKrk01PAJzgcuv
dyb2rPhVuH5slFEUZxz/V5JBO0sdXESHiM+gAamuMhtMq8pZCzGS+3khgzmAez0l
uBvdY80n9rHw8UOz7xhvFnDdSSaVxquY6HS/nsidhFWpHJMHJl2H/j1toCQiNe7i
H0VUYCztxIZn7ISkjexGy6w/NOW/5B7epKbCB6gUHsItm3qXKh/vUbBJGxq6LGXn
nS0emadGYRaqixaATlisPjYWrjWjjRzpUSRX18uwmzLgQQY0Ap/cWbJAGvDPyqAh
2kI8J+R/JCTQYHXl59AqBb5fpEBbEfANrA1D9TOl+NGquB1235nawC05kXo0Pmof
TVBbvxlcwqZ3sR3iVzPO3ASDO8tfvk/rAB2AsjcfCOxBjwi6kwodwH5JWthhywAF
qsnrJ6Zi9x84FrUHdoZEhjYL2BblmMMJQVLX3W6EH5Yfd4i7hcLR3wJBGbPVGqDl
zX+0C3OqesVjNsNwd3+taMnaPAaMvQb+U41wu6m03IjrE4WRCwxOAXsXReTKJW09
U02mPeb8MBbRh1Ijn/V7j70v2xIZKbuZhAHDubtuFMP1Io5+tnUs0l2z3sNv8YTQ
Y5gmg0JSWNn8qObXawp8FpaKztz6jJ4WD7atBhd/ZU7xxvaFeQCbwji+5RgoZM59
J6YCayFb0+/yINTT6wwqrfmJ4vXUapw/TuNvWAYAiU9fIUt/4Uw60k+QRu+27K7z
/1UOc9+a5b7r9YjnS2qJ3UFWsJnAdZhhvxGgPEKYBda/5FSMzWKqS42ATB37e1Ph
bzivMwloO5fvhJiR2G72mKbZBzxDTYCVo/Bf4PX9uBREjhqmyvwTOG/eKjiXZYnE
/Kb75y+WqKEK0bpSN4Qd8Zhj8caRM69c5zz9BF48eRJWRjy5WJuQ0z91LO7En0ih
vL7AnaV4/5IpRPSkuEp4QPYYSculqi7nrxdiBZUbisTVozJ+eSDu03B4Qb/8jDHh
jyddvcnrB8ty0uXBboJjJ+ohCSI/1PNeOOtS6BCNJPXczSMaVSQyIgCLNMUfFtUP
2zt7ADCx/xnDU2ftOLq1o64hSGp5gi/YCGN1Nf/d3RLE95Qihw3OOhk6kuzzrq8f
qO4fLxkUPacM+dTouqSmZ/dEJ/pz1D5JJTVQWH4lL12cKM1kMSlYETiz4hMnDQeq
d4tX9sM4BUgGkLSjvox0RVHQLf/2h5tl68NDPsPiId93fLorZq9XZEAs2w663GVg
4s894rYDJ6J0ENrUs227Id0uzIN0D0Cz7xDIJVk8Le5dJ6FjClkOwea0h5RB2/yR
IENgPRk5drUWXCEd1+CQ4cWvqFnYIlZyQtPvt1yQFDOvyyoaZyMOQyTHJ0d2vz3t
OuQW2CoEAVwckDHcvILbusyHQW3mUd9Thjw3QW+lJuBJVqtTDG9g4glhtafz/29H
I1/WIyUPhS1AW+Ly7KsB79dlpowegQF/VuytOzhZkWfMyDgW0LisaohcXN/zFERr
0UjEmDkYqFCWqeBCr/1QstTBVEu5Sp0hElM7hq/HmxxxZatNkDdH0h4mSHL14aa3
ffRF1IoqinpPgshpM1VijcjaiNHZPUG9J2KFaNi7ACeE3jIO/WmEOUPhdsb1TB/7
22kvBiDAvy6qzsGnHzsPuMeWy/k22/+ovkk5C6z9Il6kvJv37g4jFuJqNqRMdbdM
Ht0n9HopoqXgXGrG74NZ7sdgZokv3jis/EUunKy9GS3VbuLttbR9nPdQaDi6SMm5
Cw0Az9/hW4QYMOCiAxdZc/lwUzCJn2scxwttVIJ6xyfhfENITPP8Zi27Ygw438rJ
lfTmD1wsdwgQH0Cx8DbeUkcw/eYLa2bd//64fi3QqBEESaBwG3zGf3dhptYS+fBe
OrnppWKbXEzDkxV+MJiyWYdL3PwhikrhBM5+ZhFayytAcuNoOAFTeNNFcp1m8Wc0
76/8RCM09igpwewYr0c2ruHr25PNI4XnXKo2aD/xqMqdpxsIXvlM+HjWts7BL3TG
l31U9LIjSSqrMkXUQpBlcImglcNn5p/wB9tbSyD/Gf3LpvHNeVStPiLMuojRwMJn
NiP1iZPBvmv8xmMAuFu4I/oSvAl/xBYFtlbQTz/TbvZGM2Wz3kkyNhEFgScXEAKh
/1yU7Q4ADZAHqT1S4FNes8GvEHh4avmsG2py5t62qFqLdYaiFUhjDVTrYSLFfFBT
Sn/ZUAfRMRw0gBXmCQHXdw8cyIBfECZ7QgiCQM3QFi8inXVGWTi81b2pnz6SUYLb
SKXTjz2GnL1MZ/LYg81epRFbsCbF3gXZ4ITm3n16TATy1OLcB9QYBteA1fcRlUro
a9Z9/tgp7sjC8EM5+sRS7il1LZgv6vh6H0rWkrHZX65WRB0R5VSj/HM07U8iIUhs
2YxwhE69rqICXmI+VhsnwdqxF8qj0d/JMq1TmMvTT9cHyUv4hN6Bu2l4Q/hMkzdt
fn6R/WqeiztM0Pq9DZy3e5beBGUNEkjNnXnqD0f3ePcacTNyF74xq6zmWnorh1Dd
Mxoh1jy5UTaNDZSkM0UgGDIh1FFPObj1WLI5u2yLyHu7efXegvHL0aQBIVXLeJrg
6mnknttU1TE2OkqyZ10sp8dz13FqZ51/TW+9Bjg/8lEj+yAQ/22uRu9dCyB8h+pB
Cmg9D0rEAo7yex/dQokE/f71ryJVBsip+aM4lOyfCs5GtzWl2eycdVjWbxie9wXl
7XM+7IWSll0TkRsy5KnA5rQlV+oMglySZSsA9PTArbM4Cbb7nHra7MdpIyYp8Qr5
TEV0WyqShzRI6sW6IoFk6nrK3aIE221J5uoyafMqTIIyJV/WuscYr0x7tTiNkRON
n8bE7rv5qBZiPfnODiZ5b3HgQzQTkfFmCeQK6nlKC48b7V4Fl0F5HNlDmQxMT4lG
up+MSetXxJaabgW3FQm0E1+CacZxwqd+iTqcUP1wkNkO3767pmvG2uDz/+g4zkUX
O0Xw8BytYvxOMzqoryHDDE8pEw+LSXv0Vd7BxVYJPw3UiZ47gWHvG7jeAmTT5rZF
FcXey23BPFLzGySdtgcC7/nsWw3qVbv33z01psafDxunU+/sC1kQlUMSX2uJKkUL
XUuEBrpjtSFsZpmMTQbUqZv4IBAAZYjcY+8qu6jxYDRI0ZVd/SS3u9NGMfPZ562b
HOuUfntRldds74RxH/cI23ZRqBhEKwcfcpDKyWnmcMpj1vHeH6CzQlO5Wg/26yjC
glwEsEOMp2xWRqLtQrhqMtoHLW0SJB7/ozzkL3oHGXJM6DFxo/YrKVGr70+oERgJ
Uc6vP7UcTeEH4dP07qaPMB1k+f6JmKp3pKhlUrW+4yeyNnI2LRWIgMPZPblOPMGt
xuZ7YdrJL8VbQxPjBq/TDqgwg119eqb1dq3OaqTHg/CWUVjNUuqZm6wKShKR7Rx9
HvXTT7jl8VfH8da1lpIDQYLv6NFr4dPT2zjA5CgEZTekArKaT/ugmKnCAubXKEit
ElcQ9ZClhvpZWfiBk13hyzhkJ00NPDZ/LBoLWvK8JlXd/UA0AfyK6BV7Ksjml883
veLd0Th+iRuYCITGd5qzq0M4JpXKgNxe5CxzIOLf5IPfmfpUG6wuUqlyjs29xeKP
b0NtA4yq0qx74ceQxDpNqK4ystsK8NFtq76JjsUcrXVe3lB0Q849LCAln08pbqOl
sXEppgx7DmPEeQPbTNZkQ4guOnCl6KN7WrEN8DS2XkinEU6WofvN8VHxN5jSwbzd
X97fIRpPqU2yqKvcLLiZkJep/cQq+dimjcoXz76RJu4GyGurFWlQtSgArDu8Uify
hoRk8givdOlDEmhFs+5ptFcGfi57dFVVEONDYxJ3nkV0KuFffzCyISntntuDxLow
MOQn3RCRclBzOuKzsMFmHB2c8WGUzMNYkFmnfAf1hbw8wGv9d5O3DOP8KVFeza/a
HQH1F6bbgJpmtdAAJkoZq2BLrt6A6ydruG/dWNYxEjGZ2MpOEiJLBiSDjWHuA+Ny
PZOEPfKqnPC9pKl/DPtuW+OAg0jgjEMesQW83BxZYpPdQ+2xQlegEy/iP/Gppjeg
V/lY5BCP+2HJxGULUVaz8qr6wwcpym+qA5e5SpQEg/HUrY0JvEcIPjBPeIu35VJ1
cHjqLcyYOaAw9UOcbZ0xQZZzL0OpK1jv7g48fIZ74NooziZcz+TVPAfLyv/dysO7
5YGzYo//PxJmB5gBhF2g6610d88hmCCwdKWn9gJ3DgxvrCWJPTg+TzW7hhQj8Nje
h0itlYRMS2z0EMCTYM9z+LhslDr39CVBF1yhbDAi3FTREUO6rcbrRmIt9fCoSCB8
r1joChDAKhLHtuQIsG7yUwVFCg7lQwZBuyjhsvi8MyII5VrIxnKz6t29If0iBL3b
rHanj85nAyFuKFFaU5FtjMtr7WXMuO7PzKOIg12E4znwBWEAWMoLEUijzhFg0BtS
iNtcZR/hgYblB064SzrleslBmfWod+tgoL+lU2KCj2S4K/TYwmhpNMxrXlZ+NqQa
AwtUmp6zbO6DUGtPw8j6rpAb1zGFAzBnbBgo2KludHiQmQk+kUIdJQJy9MMWBJbL
bt924UT6YPr7ZrFa067Iol9X8uli2sVKdYBH2y0WBxYTBg5N+vR5eIwyMuML4nFh
JV4Gp+GOJpDMzKVjQyqqYvj22mD0hXcsfnXowSwysa4ah7lQTtkU36CypEuxk0QL
c9eLtPV91k4UOjZYWVLavtv77j9Q8xJajrVDgcrkQ/sThmSahNEdbtI2yll3OJWw
RRPp2emjfXoRINr/SdJBHaKr82k4BEJLzkvO70sSHtJIx/pbhgnLDM8l65aU3Wou
oLq91utJwgefDHpNq63c+RxowQiO/3tvZ2HWA+Q/eo6ff3O6Dua0mSEWi0ZImge8
ytN03ThKSuW2o6qg0C5oaRtbcxKR8R5/s7TA2Ho+yohnaugnG3l4gEumXLft1cE8
KI4IbNGe8u4P3kocy/IG3uZYvxt0vfq6vePgEcU+LZi6bIAKVwHJzDLKu5f2zmAH
umedkQlQ7Ly2ib70b6e/euzLNwEM/rY5XbsLCQPHII3+Lcm+4x7rO6EjX9lMv9KE
8f5j5eelZdyYZ03fg1hzABvwqCjwMb1v3NutWAW++jbwEvA/cVoDMAmN3FQHDZNT
+l1RvtXjLQKQFxocao63zGF1tSeOqJYBLXAsVzGPIIDsa09jrPuBxyPiLRlOdYG2
0TqqTNZVSzA5jF6Faw2Lb7s16ve6kgmiYhgAh6/F/g+1C//UY+r1OHNeRVHVw2bQ
j7J/IdNzcmT/tCUs6r6GWNnzNtEr9aEJKNcclmNRTSLTqhLSWzDCwa7yNfCCzsMB
xKwetk3AHhO+Jc3NWjn1tX61vN0nM/jXYWxKugOGcqbWg9FRC94KHSQm+Av0DxKH
6pnRNprlX57a1UjKPLZaX9GeaDPsLk4bQphpUQmwa10XGPkW7FG64xExZXVUwuIR
KTHjmAL8pZYSkT00GQIBR9Qkil6Qv522UGArthyrb/eFntE+cEKIsxQwwk9ZhZs1
N1soLD9ROvuhgKBeUo65ctVLK6/N7P/IBjt3ghPc3vS9TOraRXdDoMaA4FuWIiZT
SBatyOdc+Zq4PqPva+XXhs2xV/LGlHwxjwTOHdnfvjAm/rwWWTG5Lq4baXWn0aIq
yfp2wPRR55klIfouHtl38FyJBXt0j8U5ZcLFxSedTpMBoChqSOr+SnnjFb1vtrL+
R/K1ZnEk6/fAQDaTpMx3+JeZJT0cOwc1LVngdjs/LDobS/g19ohTQESQH/v+NBH7
qdF6L4ULtHSzMPshrjxXZxhIwc90wXatjpR/I7K8fYktXIg6GTj2getBZjQiOJii
OZNe7McbiXWrDD2tv9OVJhEYoD2tqB0WiFEs/RBsRisbinjDALZu8Qpbc9j2PK3n
rFndZBTZeBxKHe7iC4njCKTfoAotWpMAHNf/K2R5mBIWqO3SbI8D/A/Rt79OU7PV
D1AT6ENcdFOVnEOyqPJ7y4xpfX/z2hJwP9yvWEP4OHuMZCfFWgM7gE7aApR7vmzX
DQoifU7VkLPJH4FKaPsFHd0l8HqjQ7ZD2S1PEHnpZs16RG9GLNOxiniw0DCrOWBZ
y5ZFs31Im8ycUrwny6Gg8SUxlDjOk6iQC5+pqSboGoAXdVFxO4mFdqbHtw+P5uB7
E/3LYqQqwPhGLXj3V/Zk9mvX+POTEy1lCCOVtNdZUxgrzxCViSRU4UHC4DUc/n4U
o7Of7ygSXaErmQCTdcocQIPkMVNsJP6U+2LcwGDDy+lNtgC8Dzmk68VrOvivtjRF
gh5Qa3rk2b9W6WnIyk4zBAkILWYsrNZ0GOVvoAdRh0nTWmMxrEITpyPkOCFEKKuM
Hp4bC6qAh4JW0CFbc3K1EVgJxEEZHNOkBYskTbwT6gUKD97mga+67RHNqh40a2sG
0kUT7jS7bqNO/s1dOe4E4EyZK8JSXIQ0yoXKY/rPzUAR2HwA/VJ4NqOuNiFEl7Ay
lHJTURWY2jOc+9/ATH4DKB2pIWaRUVRrXaBDhujU89FS7tPQKn1ZBEw9hnOUKN/4
kXLbPV2c1jRkDF34tVuUTUV/8WAs0xxwMp338zXL+7bxwEHQGR54MozMCm+gTz1X
wj5gW6duv3kfX1L/vtN1UYvSyNucVKi+/pETAelhPAFeNRKDJcBLj6tGbvw0AqDe
tmzny1StAO5zf2+Wg5Oi+Seg2zrh0+HvypldDd9Om7BEYT0GW9chZbD6ZMl5/rKi
QfZsP0g14pmZZW2a/aa4e7GUYTwDSO7XeVCdpGAmlj1UuQf4abFea05/AtAiTwaV
pH/iTFc4IFhRL+RgOeUmKOCVqK713qvmxoAhGDZNSfInX0ej2pouu9OwcXZeMfRM
RtcHyCg3lxyoh6+1ZhJdt87YzsU6F32wQ4mMTmKY3XOW9kCfYKOgGT39OZKaaCW+
wvRNPWIvwuJ46XFzycTHg4ooi38UyA8Xdnsfg3gGvndRbcnk3bVZAqoLdoyW3pW1
bNN9V18JvkAXQTa/sGXN+7YReiUxv2NuZV8PRdyeyKVvux8KX6s3fhmK8HKzoVdi
KvrABVdLP4jLwF9w7VgK7zMrfIXPR+F4jn4ywreWJL1uvVG6FDVpMkjOCAFbK2g7
UfGB7cqKp0bEXG+yYSbpFM/0JtpIsTS3b0+BbcxYK9PBJdiHvvLd7zprBznHkF0z
TClfuuYVmOxtLu8OpxoVtesXGBA3Pq0iVDg/v9u8TMVKdnOqrXxQh4dq5CeRa5Mg
C8IHEUZgThSBvbvN/Rk3TKNvtKcPoKCsbzLlsPnQs7AYLrrz1eOgQasHVICHdeL1
IgC9ClH0uIHqCbVDSxtjvO/X96a4FOQhvj7c4WFYLw+xnDxulqA8jBVllosQjN9U
7KqdUFSKJs9Ruc9LegHl4/NrHl/ukAR1np+/oGm4t4OaBGn2KFGVxV4SbANcPJBy
tnIPXWDv48NT6SoRqyCYg+k/LcUUDW3Bbpzbsce35flOxu6+H8G1LQ9csH12Stnt
vemWeGocUuikfCSabXzdpdiPgB1p0cxPOsHdCX3cROWsDkHOOU8niD/1CHWKUQ/a
28eQa+J09SWeZU2PZDH2DYH50nRoFfUkTtSd3T6TDbbaJtXwQsevzG/EsgE1//TO
KZu3VHx0jSeMg+mKWFriRqiUFU3QxFaLHBttB52YyrCgWa+vOyOAyEBwVzQGl1lg
bJTeFY+TzQVTbHGK0AuDfnnoDBefahuM4Y12cflv0IWRAuAAH/6YY9iqYhEDCleq
cks+9nsdIj6fs3oBYy7RXOeDHKaM9nLmrCvm9tBFfI3AVhH0lVx1dLZbgbBBGM+w
DB8TJNWGmXVnaRAVup5Wddv+pYOJFYjGS7JY9T4WI//s/NhxDZRUSRjayl/js8YO
qr+KH8aCMG6fQTC6opj0FdZg6ddH+WvX4tTpG5baNS3kElEa9vXvstJgkndq3giQ
urBk27uQgD4GnsDyZ073CrhSp84wyKDqdD/GQrbm4TlZZ6CcL67EkoNYsBTmvhwD
1vucBz59BOQP6P35nI3gaxiRPXm5op+yB041X76ZWVfFNW7/3cnCDXxhI9ZCFsr0
KiovGc2dTohNBNBqQ5u4SVRcQbzJvs22mmvLV+1IXvHv3tiAkbNej2dDDRQAH4MK
scqzgo1P00s26iB8pi9RdWExhBGcOoUL6KP8fDxWVDHNokVWKSv1TBbd8ZEnK+MJ
0teTiKZtM0xOR9rivyCZu1Kzh7VgyYcYahjRJkzmo9SwAxx+seCp0pA2PzdNK6A/
K6qtPfbsBT+cBLMm8Dk1DNF1j5reZlFKFRsq9IYW0KTctET16vJGiCFC5skIe8eY
tmyBwOb8OIxVyZiZoN+47uyPk64xecCt3xryptPVgCnZYf9k3AooXv8CI8LV66HE
u/fqW6EwJ464jvvyCY6ipdLkqnBHAP1p4eyDr/AgM2iCDCW36j56Je5YDTq0z7Os
HGopz54yBM4ga7BmqMopEZrFFui0+kvzuUeP72sLyg80uKqoSUeLdfKblsq/Y2Qe
F1ojRZHjNHaHqxnkRg5rInTAy6WjkU1deQVRbUan8uTr3+uL+gpgLf6jgtNAwLgS
mL04S/Oa7XTsiZGvIMswsuVFI40KqmeSPF2iyGDdrLJPq3091aBH49RXpomfSaoF
nBtr4wCeAQFLvuq5kVZpV8Cz+AbNMsfvu3LYXPu3B/KWOaXG2QTpNBfvmxUyXbRj
eD7D+k1X/CkxFo0QmbuvIWf5K/W/9QxNeWM/oG+FyZsWD6Tw8J97fjxxLl4TxsUi
J4DE0lVpWV4a+o42LNrb+wSh8POVkRcFU/VNubZpiqab5O8kJ2NwSZytYy3ymcJL
HFipN/8W2bEr064zYWud7kyvDW4gdIsUyf364+JQi3gRzObxIupS574EuBJ1Z0mY
uALBr5WoXsoC2Duu183OQ5YAYu0mjSN2xkhLdJpBHH5dtvM4korFEE677XtLHdaQ
TEDGZ/+b5yKSfIu2YvSbvxjUtIiezrKO1zgsTDjkqiF3UtFR7tJ8+5HDutbRnpv1
X14Fn4fl07q2+dr2jA31PbLsLFMiDVsfQvvaxmXmMBR/4PXFzzar8mMtr30sXMKQ
g06N8JntjAWTPXynB4ppvdcCsmTaRoVXZVrE9c3ABcaqT5PpPKvoB01OUJirvbHt
j64G6WMT2PCJQJa89m8B9UIW1h7OACE2IlV8ruh9cvPVTywtwh8y0PDdwqdtjbsz
dnBnBxi0NwYv+TNiRsk89Kf3PngfkTnj0w5TZn3a46o7jQDZsm0W+Cd8pOzE3Owl
IR9uSIQEJFHI91C+oFC4f9dq1eF21jWzjYv1M0++o8zJ4oNsnLVbfPfYB0H6xUOq
4j095COx+6hqq36Pk0QgtWSociF+Hw+LhUK6l7FugkvV2hNjlyQVZnTlwo8PVcT0
EA/F7Cer1NP4zDkBiE21T/81N0EnaqSr5NcF3ooEYDiS1vSmE4Wf9GmMniAyVebS
B/FKYT9h9M1O1/8dLwMHjA0XmeuP31kNRcRGo13g2tWQdAfmdqNWhOj3T+nw/PSD
xhRmweZkPLQlXJyKkcxGIlh49Ex2SIX0wuXvoE0MsKNt//iYfdH63Eh8trmFDBg3
F52/DrGTMw5vxr2i6ecEFdUa0EOTA8B9VwE8s7hM1ixoeLkQ30DgZjD/K96SqmAa
IPABGf89yvQ9AlQlS59uHDFZUwRAPQ9PuR2WsUco0ZXZaaykek9k9TTS/BKWvjet
96wupeRxlBxF+eqBKo+UQeKlm/+CpRkcUX0FYy0b6d8XCzePnPQuCVABHKXWLoPK
/MdW+LzcpwSv4I+hXqY2qRYN+KGfVdIH0RO4I3n8owrCovyN4O0ffpyAliegLjn0
yqaVv8VKctr1tC+S4uvhSDnPQlGTUs5ziRXJine6oAT46AoYbJFQ2baYCBATM6zy
Ngwrf8kYb2beH0NLt5qBcElBkDFIaWylom9NB8Q7i3DJ0jQBg35srE40qyycxqFL
cdW9+70ud37o33I2LtZk9j0N9QSCHFN1rd0+61/dSbc2iRpl9TN9p5p4euw9tgdN
kZ94+MLWEsvkWIPKuM7uYUNENovLjN+3SOXT2t6doL8a4cZCcToya8nc8erQPVr6
JXsKORbyaX7EFBh6+rckfcKtAuy6ySTAEk4M0H8E2ilSig+K5U6Tg7dTsFlfOkAA
wQYH9tLgNqReui9Ps2cKOTnfHYPPZ2hXmH6ZH3+yrNFO2Ptu8Ms6lAZeKQyIwGfq
xGXymCntEjALawEyKC9PFLmtMtEh4nbSvdc5LU5QNFqtMYpTLpy69inwWmeSkUvn
SMc6N15V3D3GUnXgEGxb82EWouspOtK/EfEPdsQm9Xyw1OTB2LsCWtyrCdSTGVKN
QKjQ+CC7hHLRBZXGM+keQ40fUjKqmASwW+Ri/FmYmaOBiPi3jy8faQSLsjYD5vY4
vSixlrch3x0BaTis8kqhMbgcoSqyM4fEJnsOsz/fRT4uJRlcNXqc+78CuVnM+0kW
S00ghfCqfW3r1aBA55jZPE9DG1idIwnihnjbQX6dWNcisPqOLC/VzhO6RUJbzxan
tJV0tptSrhhUgSyGAIYP5mz9X8GlnqqDqOSFs+6S4NgrZMdFpPqQtgZ4OCb/5CR7
CCjT7psrLMVP+pOOa8ynt3lEWbo64Nx3tic5QprAIJgX9gn497sBpWP92MgurJk/
azUYcoFQ4nqvq/+umW614j/bJkoYcUB4C4WbfSVi9XpAfTmnmEJVzObLYI5f4ZOr
ihbhteKIT0SbcqqziAmpEvzOMUx57VriCfLqbYxcstIxV/PJhdSPYpP1KJRf54Fz
RQXZ3BwnEnZgci7iyCcuxti53nPRR4VXemwhf2EN2KD1COIi1OUR3of2TwJeX02X
aRqETVpGwcyorCKbWdZXjjqFTFIz4z7Qo1US/v1otzdicX6jMTLaHbBiI08GGG57
J5VL/qnew5orzelebpz/2UWndkhSzaaNZLwzjwdv5ylrwldLDqQedYZmdwzA7NRT
6lBEI30RtYFD4FpA2zLHv8X6qDHnTA9xYRQKfMM8Z+X5EGZJYHYVs8nTlqf+EfiP
HWkc2eS4bGmqbmk2N9sfF8Fh/olFLUb4CE1ozDsh4mK0x0INJP2EF6GBRvs4KDuQ
sf+w5OWETCgyRZVgILUZ2m24UWURutPtGyoPVir26Lj6DS8Rwxr1UD5nzOHdSiQ2
nnpEwMy0VEenS5/Z87++XOVEMQPQ4HzC41PAMxRZHGnD6zKGYoGT+97MpamBrKtk
j+5A/hvwHFNzCy8Q3nVti7UyB+Hz3KlyKzPFxbKjM699AdpgEu69gb/8QHYBg0GC
O8OP+Yx9BNTLwfw0s+VQ9jnU10UqahmmHN6olsFNKBUhftEHMYiEGUIv1UKuW4u5
3TksOr3ET8aMjp2ei0tsiSCNOiGJYnpn40XqlRQLO2PTjaAREnr/hXknXkd9lYsO
glM1wHykiMUSjP3UDygiwWSd3xCy7wOdukODLEApSnocqwNDvniLkgbiA6rqS3hP
OwI4s5dWioi6Tx36NJ4EUcHDol64v9s61uIR6ZheV2HdRASlLLA61dpMJ6MK4bPk
8zi7v0vHC5nhATcDlbx7lQRBa2Xjf1gbprXj1sI0Cx1DvOXaFB4xXjrHXd+919kJ
JpbZBIzDYYtVit82WMb72wV4O5FUDGNMS+bSEomz/WbEbpv2PahV+4ZngqEUkUA8
hqistFvUg4sR5gsTUU5G+jE1X+0hMQe7Vl0FA2jzcLthOjr9Va8ibwP/HaEIlicG
AYQjwgNEtsG0BfJHHnYh4RkzgK4wu77BSA0Mg1ASgruhuq3xd1zlNHvwygXc6mlJ
o4u4MN9NFtrRS6BMM6acOjYpNK8NRBIt0Thv89reti0ewvlGteYqKIRUDgiojkTR
QL4Tl2nidD0EDfn5AkM+/jJj8wo37XPasiMLIESjzP5ngyFVPs83hWy/92u4cJBz
AS96/h1iWmRmVY9C5hzP/fS+4oeSxbt2Fk8VKDRxAIjj2+kvIVGp5RCeUmesXT5E
b/QmwJg+C2kKNY0OfDDCsXvCRRl3b8qT2psjqxuYbO0Ak42yblnBUNLlgkodEOfg
zPOjpeyq61PHU5QPNqwDq1DAmyZTyTEQi8bXPslbNsV3eRVzGCqi+M+7u7pPmsQP
6/cuzG8j+dXN47y1bBIUNqW4WVMGxXH8zoe7SzwFja0m5yGPg6G0zOacrCuVMYQl
lv8yrH6FGHHY6gYITDm+jpBb+KiQEMy6OUeq6s7i2ye3XlV8VUpgJ3k3/7PzfjJ3
7aeC/H9sbHvwlWGkDYBJSAT0URkLzUMcxYUJ0fdlqSSKeBdURHscWHpPPTIE8I+S
JXA6Ss/6X4jEwMXsubMq6AwQySnO8/ydRt6HRgyy8T/D03YXZPzWAIE9Tu/PUia4
wuA8vp3X627Bhbhr7zI+5Ynqju/Qen3pBQXjqKeFDmML3/WRkdDMbc1nzliCFzLl
CRq/WCRp4Dgexvz94g+ektJ0We7tkfj+Zcsso7TFomRvAjlHY+Jq7fT5KFR6GSGl
rcDvKncfinZNcniLIDWDZ/scopKG6zEw8DreqDqUSm4yYy3IWRLDIg2H1UFXmxac
FaFmPuL3blGJKA+LQmrQVW+Dw7u94hwCJhPm1VjcHipyJ/8wW3fipkOWanq3FgU8
MjwpSHipMW7kAGvm94Bb9Zs59K4No49KQqugjiErgDnOS/lio/8Uy7esWvo6mZfn
x20vZ0+8bMIH9DVrFw5+4Ho54U8cwdA+9nwyWEeJW/ZJgRJr/7NAcPaP6q0ARyjg
C9AVG1ZgfBZQueZpLyX5MsY8tHCpz3pyfNXajQU07mgyptsydmO/EUne1GQz8KDP
nipQ87CyZ0kJFGXe+EfvpBSIR2tlm5esENw5tY1ZtCLn76AwXkee6bCKW1OM4GjW
hAz6pIO0OjEa63YLiBHK2PBZM+96MEQXWmA9WTPZW92ky+6dxKwjudwQGH1PLeOa
iofvbe8z6MbfpZ8cgbAMYFGwZ2kP/4h5CSQHqGNLFhE9/Ep5Q+ium+f507yTMwYa
OcJBJnXw2N/YOKCVb4JhPWrjXeh0WgKKn4WVkw58VOFfrOSbxL+lmKHvawKspp4H
xq7RnCtIZD8++wNyiQND0nj1Y+tx1J1HbomkHSBu9yLvJG9BGsORNFijjIwXEfZX
WdtinUaFTcaUFsZwNiyIX6X6pYNmejtgmHiFWdGA9nqNH/8RT8udt8KTvsCKdMOD
CvYNmDqDBWuwcNB6EWmuumNIdQZeByY/b0eeynz3jMbW0ifju3mHRncqdePGGOVf
ohuY5ytMpA5I7OLNCMXLIjpn780ALvxMnVJOv88bROidlAgpG2ey1hHJPVzs4vSH
PZ6eIHuOphBjPe7qohY13hUKuM7ekD5FJN84sPlyY6CZmS6G6+xcn1ZZH5awYurj
vmFQ7YktxZNyy5krgZ3bXUf+sekZqxAN5bMbFgE07KoXIBymLKV4YZOe5aQ9fBa5
HAC8EFXhEnLvOW+bZK03eV2Go7a7b/oOIACuAnLTqy0DGLge/gVdlZbQDK1zx5zb
xnxQ0gEp11/1quKch78aemzRKSXo2AOFowZw6QhSsSLWiqhe+jqh0JOaVLbtl6uV
LrailsT+YANh6ikkS8XhHCHouzvVzC2pDP4MQfzBy2WnchrizC0dJnZwDzLMMYQY
29gMeuyiL0ekCoFYAhswR/yK4fh/9y0Wi5xDQhO6+EmXPBrRsWWRVOm1kkgx6cy3
nRwgIXvT5dcCYEEBVv86RsLmTiiA4YU58Q35zng/krapej2jSrn0HfqPmE1snQJE
m4fVNXr130CGgB1Hu7LMw8uLfzEh4MwBS1ATCirD+zLfTLjdj+CY8+KCCPHaU2jy
y9emI/v0fGgPVAHe3nIgvuZJn1L3Wfmni3wgKMAgzYAGl6vyqYeFhfv0NGO5QtJ7
3wrwM6q5sckkCEfP4uANiSqIiw/u8iL5eiuli5AiyC8mUeAHr0/p/JMh01Kvndvr
NAEheqYKZ9Na5Cktn2u6gfUq8WRJVlavWqFnIOYsws1ABp4tJBQwPEM0BhdNe+AN
tveB8k1MEj1+DlSjWeuWRbNGuq2UOp3XvZHAvWc6qE9tXV6wfPNBM2Rv27lyM8jH
5+3vrcTAGkI9eKkH4Fr4WqoC4RHPHLfdOso4a9gdExZzqcTwXNLqTAuAsRi/5I2U
Mjf9P3l/aB3E2ar18BygIXCscrAKKWSHfWALPvvWBPzeBrzBFi6IDFQ24HsmDdNH
Dp2auGItN9zvB9kRGijhXenNSxqYTyXUc5MoRgzuVRv6xbJS68wsmOV3xlmqtH9Q
lEd1AN0Y1efB1xeQSPOnT9rxJsx5vCp75IdNt9goyiLso/xvFhFMPugF9Zn5ihTE
vUYWwgNVUTNtXB+yXNMaeasNZMlrqDylACbOikYpiTwQNbuSZBaFig93jO6rOrjl
qfudRuHCNVz0h7FDroMNuwFSUHHe6TsRcOn26EY529MmZfebEVT7LodG1RZDQNuY
Kxqyo52+qm11K1UF4zbLQWcv/emrx6p8QBREYHlZGvMbP3vXiQWYj2Z+ccwiX+PP
k4OE2S20cBTx2h/UniQKsMwNV+mbs2FEdnC34/tSMbbapWfVuL1LVKw3RyBPlHI+
QwRRtKD366MLeG5pSjPIYpK0hM54bcBDJydgof0csdj5/MyD3sARfrpx5hKd66gb
WKD1dingpMKkOmDLv92DpmsueeNaI4SZMiQTO4BGVjNq0hvFNeBVNrdLNJMKeHD3
6NFT5RMzfYjVMJai7k/j2lRopI9+BAPcRJgc8XRGXKY+K5UZzcSL0GNr0BML1bRD
tBuWT9XsVRibiDYbjKtKQKI4c65mba9exca2GAje+b8XzLmcvP06hMtl3Z0RUiVe
31N5xwbAsvpw1B5MTbcYSqVTUrh022/wC8rovvM+XyaZvrQV1zrmNeNbRSBD0QdI
lhiLQdDUZesbbBWukdQIIdUxdwH7pBc+9j1HCQyNqXVRxUUkCL+ggb7MHqUcb5JV
gH+pdiwuTNjDXWQOIuaViizi60zvs/AfwW+gOM75+IrBlj1DmmydifpRZBH7IVij
vo15/8xdKBA2y9SwKqc6xgq4ySFl5xCvTp0Li3RPt1LhGTdcpTWd+pVKGtL5mNLh
yPJL1B26U9s0KK5546YzXwp2CRaulCVXeK69IUqQtY1I+izDxmKzaIgPtBx7FZET
kGTi8iEmygxG8kyfoHi9X1JOfGYW0stDd18iQE+1pra1EY9gwUTIT1AtSc1eCgc3
zDxArytzRqrGeg4AYFfnprl75XAfqcrSE2nSLmeDnuh3PukCzEhftjkXse7Cjgp3
wNpHw6yc0wt3yhUbTSJ9u8XxLHeOKdUzRYheWd6vtNSwsw6sBe+9A2LOvkwNodKR
orO4Kux6z0E9wRlx8hpLJu9Rr6f2nbvH8XjWMFrheOqfL++1YRwOCuzAsS6NQPdk
oVX3cwT2WmbR6/W1r8j0H+P/G9YwD9BVUI2CC+2KoH5MSsocRMYH7dP0560rst/A
9uKmULqZd2dPOWtrK5lfaK9fSEqDhQ2wOspAoBvFRFR+KkavzMfe6qZw6BlXLE8r
zXOvBtCbHm50ON0S6cg9bJLq5a4RC3lvcCz3TGUugmASF9KYebeli+pVR5QbMBbk
2bUPqOD4vjFbfSCGGo0qROeb7S68CZOQzdxDEo3ilNgtyq0AMbxulL9pjWmX0jru
HaMRmQtDhCaNuHgxohoIAaRLr6ePUDbkVQMBnLGbrmxgfeGBjX0R7ycdhdiRwp3g
pkZTIm87miX5M+rpBInqLBcWqFh2wiKF/zilniaGSzwFhh4fE1LqrlcZa5Q26DOa
vZrTKhfcjwAId6U54/zlanateaWyAuCvwdxyDCAOmdSfCJulGlEPY9SPI/guruR+
gWD6lvMswLbU6M9TdVfYLRB0BHdSS/YTKTR6EN74Ed15BDTF4c5fC2Y2dPW8+20V
JLJ+mqAhx00AYJ2izHZrZEUnq9+bdCVfHzihlrNy2NUbRwdW2ZbWeJMh8eLYy3It
1z8U8J3SYKvbOyMHa2/NEhegzvi80eVg9JK+5FpIAbU2tJM0579YSZnG+mkB74+g
t1l+NKwkakrV41wOUksENQWhrTMMPsxPrhUlDbfv1T390ZAv+cqYMofIPJFTzOVL
XyQyvG6B5IBOKT95ND4TrPO1EnnllESj4lEWwRpff0C9dTsv6uVdqcS3aNvdQiiN
1TQFVTHi2oa84BeP7e41ShWiCaKL9r+mhd5jqVkh+czdCxDpxIKT/+5wRG4DRJ6l
oYoF4TNPVwzldsF3WhVdqzXEd/ZIAJSCVRDzamomwfHcT+p5ZgX4uI23asVBd18+
WT91eKtAd9CNp/aVaOHfxC9wD15qFknheRQOofZ41BXO5jrca40/hQxaykbGfHrg
dJXTkzatrgsBa+gJ9MrERD66BQzpSfvEm62sC8DCZqL/q2DYceyumcUt4shWbuSz
iWgfZLFXCDHLHqSjFx9NPzHJl66DGPTlThZsD+JAZUTmCrlAfOrVK4oG/w1NKFNz
vrxtRULrO95/Kzka+Ka0Mfcl5aTSP1bwXSnA5yJWcZQj1ODNH3S3ZAZCimfCORUB
1gXNnNeaPA6jFoScGuLjzceJFLDRLs0B4LKeijEmLHQ6xxWVf4No2Bbqe5Bcvj56
XwGkhe2EVsW+hQQrKHByjMUDJ64DyXr3OWM1UT1BLbiIcv0C41wD7qdpm4snth03
smoWIR2mGszNFGNaTGqESJhQ7haTqqWtWmRNf+jZ0iuVOqtWznauLEHXe2p3bM4Y
vB7dGlwWKRjRL9zDkx1vzf1UNSGOmjyRBUG2Kyn/VabGgZvf3fvJOt2uWrDawTA5
mvnBY0Za8NJID/N659oUdHEXYvb3FH27XT0uNNepQ7cz1lVyOXI+j677arbOiW/M
McpRATtVkYuXKDGEHaVBjovRQYPsxpGfnikf9ZweB2g8vwBDD7nKyMiED/ASuwxd
7GDZEqE4E2N2V3vMPC2LLEu4YOWXEPYak3gWxMA1ZqrD7f9t3NToxV7EkUSF4qyh
a6Kj0zG4LYTIsCRobZSAv8tBDEcHE8kLPXOQ6Wu7m6CExn49XD9KB6hK+AFFQnCi
HEFg5AptQVzxfHVFVC426GxfKwJIpTX5W0jHFhYaQdPyo7rjIe6OTXV0VkCIM1kX
gidlz2ahLAoL7Omc23aelq4oMCIN0qDVdchEVatkGfw5/6e7W3e2dl2l0Ifeutb0
F66TzZ9VQRPhQAtPZ9oIGk4ycADSf8pwj1A6mzi7V7qqEqukr1M5BCIScQob/iL0
2+RrIO8zYOlJHS6RKMhK8r+Ipyj8/WM5VSl5ALmMQLbt0vntC0xLmOCcjnW+Pr21
dj9QbiJE0k2qchDpk/Q8Po6szPh40pYBMN8BX6g45ZhevrBoyQrIPHNqWHOM0GMQ
cCBqifDPYqED6aAfDD9DF2/jAtNVxfD0PHSXvySBDyDFmYAkTi9M8NztZ2jbfx+z
ivC48XE8RmIrcjZLreGoGUV9AtdT2gzMgRuQ3DyEt9FlB2vk9IscYRZY54Wdx8N6
RIRqzLReUETCYo2JIdakl1i8SAhA9DoBzvGwDKwTk1DhmuG2Yi6zwqmbPgB33Rgi
xIg6NmvxUGL9CaceC/LOb8pOH1pH0AF/MBETpX0dPMRO5FkYVowE8LineTtu2Z3d
i3R0AxXTMxm1OOMEv9O8Ga0yUz76PxapEFGmmpgR07zm0JQBswHkKJFOYIIbmCBG
mjGJzJCVlMU643Ca3jBzz53ywgeU59GQdU8BYVLzT7B6SA7cYHJ7hyXfLVjsrmB5
16C9TaaIIRtrUz7LRrJ4BbjIu1sMk7Z24Dz1VvDEp7DY4L8+AIX4SqUA6Sod8fCj
ai2ZiXgoFwVVsACoizWDKiBi85vPepv2UJb6dr6FCDTeBCshsnWpZWv+RSJJ/HsD
ASAq0a0m2M+ba3F+5MmiW8uTL+OYate486TveuOG0hXvMciUyPzxkNa+ua3TaR6O
OY/xXj5D1GzKgGTTahKTQrLkq8Ue8K7iGAX283E2PCQJfUxXIMl5CLRtLfBTu9ZS
GnxvjSzesSPXZhelSu/SfXl9T8h3HU28UIW+e5xk4iVvPHO0x5Qr+Pe/y6F2gWJa
Dv0sfIsrR2m1NF0y3o4ZfOFJdnYP08XsxfiB4djEUFzfLTqpin0mqCK7VOmBvQaL
lGicyvoLUaRRHbyCVPeIQKmuR3G56sg4NylLq17WocDgKCGjLApDgjAcI19iEzyU
eq+VVOF1ViCTso38ZcC2oHUmfAh9iqqbEL4vJMOOQ2JLA8QM06Rp3lSBMlmjbw8y
HBubBdQwyZHyZNKqTVpYRSytjIa7d5IWWIkvRfkYKUWJTrvaKsFPCvVMl9nx8jQv
ihBnY7d1u69MKB0DwaKBG7q1crSD9HswFSYuRiWWJgiH+UzvTIX2wHeC3AZFCuEL
6YgrpBj+9v2vOfEg/Gxn5Nj2z64LXlWLR1wIfHOEcoqnwE5DfLb3wWH/YlMqylHK
MsrjbrnlGcSswvjHLJjfCGcrCaVDIX4F41F2w7Yi4iVdC9z04IfKcD72jHchhYWV
UqTnKBMuggYhH2ICxN3NOI2uKFBeWjRTzNlXbrzU2VkyE2i1ccHIl8VEcOe9I2f4
vYVHQ5Wj7NlEpGf475enjjabivBcwn2nodz/pY7WIwTvCEnBdj45mFxATB/Ra0iQ
yoZ+loj6OGTRoyBqWQgdR4Bx+ULYuHFvKP4mf/nKK/ttSTseL6hAXQhaLLGG/wtR
294TC5H0IoFYBAVgXaHziDiDkOna4Ceq+HEXYdMbygWXbIdAMTy1uEJqO2yVHJPs
R2/MjgSeIKzz+xa+XDiof1Fw5zqo76MHOQMOGXmGv6fftVwmfYSXNENQKy+iTPSJ
uva3l7fuEvMAfE2scxuXqXHfBypHQrkyw7BMgfngn5URCZy+6BsF8QawhH1FyRlZ
wx60+WGSHe9kWKCEZaXblRzAOnsUbercHdg8MNA9tUwO3xR+xwPgr+Wz41iGB/K2
hpZjXCQtNqwkCXAOQ+N65S6J7RZT2/ufrVzpoDHwnxPPUDotSxgVyOTSSP4fyVVl
eYXTK+nVzOF5xLs7LwLS4HIx4OZP8OhZBPEvybu4WfudnPn34S7jBnnJdLdq5XYQ
axGpjCe3jxHARxXKQorwymMSki00TAVfleIgbr59MWhWtHYS/RN2ESuMNv9/W208
hev77pTmZxyg5AzCW6EyTChUCL/VcjWCZkcHuSgYM8r7Vp//tD6PP1TLxp+G3cqq
BWZDW+cMDBSnbhlB2FZpd0IIzLx6m4y6qbgqe3sfRHGInEQxry0wqSuozG+e9c6J
bsbUC80c1ETDYoeP4XqJLz5ky6+/hOWP6wXdPotqC6TNQTKjhsMiPD2gsm3bpJYc
r5uE5M05tMpbBkaklmo+mp3fZNn/G3vvZpFtYATk0KwFi1k7/BB7qfwGk2zfUAGK
scnpbf/2pj9bDHhasOHT4KnJM0fG1KJ7+TQ1BHklYeC8U0xskJd4IUOFAQxfIOQJ
wJaw1cHpn3x3Y0PStMdDHKm8DJbj1IUnCqJReM2oQgZQFaM6tMa2sYTSeBSN5i+Z
wz1TkQ84GxJASsx5+oFeo8TMqBlhDyL1IOSvvjcWKxuEtj5J3zQEzirEAxmwncBk
GZGUTB/BVgrOxHW7krSEAs5Ht+iZLkWsHkn3vPyuQUb0OEGZPC2RM6cni8rVMoMT
k6or2QOjh5S9RyEgptOpzaHLTVKmL5/Klcyq8C6E8wlJKpkIdbWaGE2scSTVyziV
ELfgac2jwNJvnRnQKb2TFqcSDUfzi4GvchsQSrHxolJ2HFFq2hIlM3qNh1u1gr5k
GJ11TFbh2NBCMLJGJOO2SGfelWYUVTFELeKhtwOtu2Z8D86BCczzKroZXHkwh1/w
AETra6kJaPNPAXRwJnaACXb3TQWGPrOfCUu8lHG0RAJV0v3CbOJ117veFoVMR6eU
Nqi8GWszZQfyltobw3S1jmC2w8DDLyzN7VkU/zjqzhlhSQi92/uYhr2ws7jBXMDU
nJAFDDondjJH2FlUnlIX276wXCSDffdjD4aE6bJ7XPRzPCyoQEM2mnPCdzTOKkcf
gI+sRsSqJT8BMrhlhSZKxzlUZOvNiZSyySLQzv/+PYVnGOAGvX5bXkOR/oxQjpIZ
Fk7M0+TTtmN61/Lpx13Y3U/V4v8DPPju/dkYsPEmm1U1pVt6YUOAOl0Ya3mLnn5i
5D3jE8Xdp1DN5yblTwgGz2vstBYY6TOfd+J0w8riTG+Uy5j2V9uekFDbkQPhMS/l
bYJ3WD61nplRtm9GaVdngDgpIynUC8XrdgTutnDsd/f9Vh8m7g1xwdR3A8H51MLR
E72SYbnM1qisk+P5hxm+QsmGD1jV4r4zXkE5/BNp/YjyqPHfwwsMitPmYl1O+KDx
XA+brnnMdw5fr5X103vS2c5utCrswPlIejRkz7cvyUsX8H3xIPN9tOrO3pZtNlMi
vNrjIHzEOzN1pdoIFKGJD/5xufkB/ZOlwrEfR5O1dapP0cb2gr5RioGmsryw6HRj
Ei2GzpY9xcwfIZlDJu13BIJgHnDxWIT4RSCd8MYGYGJ3sNfBpmXq4RaxYwC7eMSN
8KEf/0VPxYA/OhiahsR87/kRs2H1bn5jl3PTCMqMcNqPo9hbIIgnHNaY2WEqWawH
g/qii/ieXovwhVt9+R4mDouNCpI4H92b33erZvJwGEN69GoI+A0Q2LyUNReRTQ6n
KTN08C7F2p6OCE4fvKzSVMq37EifvbpCfJHCE4j588GBy0wjZmcot9zdWVuux8uK
a7vAfJ4h1TNbODxEEoyyv5ykF5ECR3qBA35IQq/KhjaiXZJOHhIHZwwKJiy7QsiJ
IdfxTvn3Dj+9HoqAh3NNshG4E+mkbUcumaZyC7XL7kRyw502Az3WkAQHsJNX+N1I
q8vkFKg6nPtzlH5WA9+xB8K4dZ5PNKsMkFjBp5hmAEOsv8PK+pmY4MJR/7uWAOx6
QKqIR21LZA4h+vgPw8CZMBStTqg4Ght9BadDx/zZUKAO7Z/+dT19U4jOYuLluAcA
wJBMRyho4WXEJaujC7R134FZhKnrrf1ctcBSQGqSDat0YaLGVXRREebmYOP9Da52
UnG82kUp59GKtXd21C4yxTwGUmMYYhm/O2C9KdKZipCyeXPuIfO/bbow9yq0UV30
gjL3n/cQH0E4KIYKWxSn1wSCh3XYPnuavQj8bl8b9B032txlGoeB3H6Qeh+OhLnu
sgFkpRxKftdn15juPE4jG+KeA/goWVt4pi6BfPCCEQaf0U2am41lFQfTj4+FUepn
sbSdcwLikSdL9GymF5hwQb8zQbBnlITkC6pdvJbkcaujuZO3JMXqaMnZgq0y3MGj
oh3JQjw0fgvUNeWuTaJYEUJFFM2KEcIr1eTGJJTvH1tZ+zTEZMDrNG2kW1Qs02gf
1xTl7LqFuMBS+W4Tuw3+tyMFXI7CH7I64aiSkKfu9pRwbrRZu/51nXwl8SjP6OY3
t6UeymE9Dz1wj5WVXhRNvaQv8XWcCmjR8TxNcnPiJtBzYkPEEjLOvPNDbTcraVoe
wyvrAA+Fm+evDvwwXZkKvv0MkeeLk2aQqzv/WlCvL/8Sy7dHJ52CuiXFa31nooaw
H0pdOOqNTWOgddJkocb3BkMjaNILkHv5JJIYLjZJPrtz0LaDJLsGxHfKGuXn11wc
+OBnCLF7y++XrMSgg5j+1BEOTpxz9O5Fx0i5cHFLkFbXP9OZv1+r/MTJDsxjMyQm
MIsFE+zkU5no/dBIf96x3qu7kTZz/K71G3lBYMUBQ7VvnaXTYIj4WM6jOa9K0YQJ
HRPKkHn7u/3ocePkZKbzllmwO5lKQX1OEbcwtVP0Euusce3LP4NqL7ZvAc0H/qPD
f/xeqhMIgzWATX15DgzZ3pYDffMmccvLmDG1q1DIzr4JlttsUZj9w/WZN8MEeodd
9/bowMuo/FCyEJsnrW5wKUaYmhyDopX4DJI91Fpjl5bhfIX/GeOZ2icIZVeJeMNR
BCr7VZxqdysCA0xg2zivjzSZiW2peklfsa2uNlsKckK8pIXL2ncMSqsYbRZb9NTH
TTuE4qUZi/pJLAUs1NwV2v2JufAtrUTYxL4PxmzR/gr7ucrEphfotQsYvNym2Byh
MqaWA3jkrRmSJaBt/FUtHVLiUNuCyE0OlGEuNQCG475c8TBl06lWRHg1JcDQqTGs
44vUdY/SUd/vr8X/9w91qhHDFnoJq5DXCKuRkEY/UdMrQU7X2OyoczVesgShJDKN
SfXC/czKqkyaOmLSOTlwpQo2eNw/EPry2YHLoViQHiueMXVeY4vT/r3vKALlBEg1
tC8YI/wc7dHD4Q02ywMlqwkw10QB6MphHzmkOPw3rATuMnzMcGIYYG2zDd2WFURl
cbsVzMuQMtkPUb6iNgt79botwMYBpnpyrWm6F0r3Zx/TiOPuSm50M60raFLWFIPk
Q2d3BpTLJiYSgJLfiY0se3LmsD8kF42UB9CszpESeQQHcuLJMHmgKCu3KAqlzpCj
tlbeNEITdXhUaXomBKN8sYvpTmWI70zPINOxgBRH6viHOmY6vThB93b9WXtX0WfE
5n3PmzTPGUbZKj9XKqVhqiBJestnA206tXG7XYXdiVPfzz5CpHr3J59q4l1Rho0Q
gFfq5nTPHLsusLUIN/I+saTY4jBnKS+l0hPFk/T9riTvxcgKi8OyHq9oJLBahRho
hbu8BtVAy8yB9n+NA1tltw8zFPSp/P+oqKNzhUsmexciSa8Q8JTqPQjXNfJ3fOEH
HAOKlDcB94QT7ZH1e7kW/TXNQiay4o9fY82XDFIKMVQuHINZQBhWr4Pqof97q/sh
Aihe69eFIZxJ/n42DuUDrhMrEpIav0zkGOZ4oQFk83Knl2u+fizt+8zot2CT4hGo
bfkim/GgKHU3IifWWCxxaRy3D0eHMrjQv3hBYoej+eSKaWoXgChMSOBslCi16pEk
`protect END_PROTECTED