-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
cL/mKdquQMRYZyLY2MkC7luZbe2psLS+1bDn6xZ3csTy5ktFKnSO0OiLMQ9GwODQ
DAlvCoAQQIEU4XJEtxmLbB7Zz6fdObzsSRXat4Ch8HNqI2s9F5DPmIVEPzUE+973
pc8P2n27R1Kq/jbLz4r2jW7Lxp6FBVvmcgTsJvWTVVhMCONtPUPo1Q==
--pragma protect end_key_block
--pragma protect digest_block
p4W9wk01hrR41hTQ/mISqPIm9Ms=
--pragma protect end_digest_block
--pragma protect data_block
O9NLmPQGsqr/3jl1nmvp7nPPx1rVeQTeT/cW/O0QqAFL3YjBAvNEdzS7xSHF1yC0
HsiYZDtwh1I0NwKDvCYgUcMEJcONjNgtYfukiZcS9ZSZaRSOvQygKL4BxA4r5eHX
aL+xnREt47xqTbdjQk2STLeZeDrmLKyRuvriNVJcG26eOSspO/XM2PiEJXp6MonE
YelcH2lMbj2g5W1BygWUctxM8CXepQSEd7PfgsJRUBAnRSTuL4O4KqMNTnHtkTzH
+LznraeHrdHV3a6J2bLXeywgvWH5+blSaJ+wxqda/f5xVU5h6m8iLd4iHhjo74S7
yUJjr0iW8cwYfqjXS4ZrKv8tJT9zyxv7VwV+XnbS3uM5+EC/Yk5redDqSMpNaaO7
e/K1uz7DvC0TzGIKHSTkGb4+lx7A8hLK0nAeVp2lRLfHapf0f1+dDxzUsVMZVUNs
EMFP929wm/nHy7s1GH/9jiHxSUoJN8Ff2P1h2wtnAcaVMf/sABZPd/4KjlDl//OD
JXhUL/N/4T4hYT7vrVSTpgPWURNrdJrbUaO/sRK3FbOZzGa3+RwPO3AEun8sjsX4
yX82HI3TRZJrO1A7qZaM7B1lpLfzPX5t5vdHN6WrLttbFM6ZjulnhHikhwpInXYB
I62lKvJ6vF2+Ey4FrSCQwyn4ZMPcHwHUjy9eM0KSpHA3U0IDe0bxEi/7dHcyXfuR
3rSPuPXcmWQ/EtR8HK32Z1aJkW2WzmVFBA8JQrlbLJZbDJ/Idg8w7DO8Sb4O0JzK
XQFa0c9g+3GgFxhqUs7lqBF7AdBH6TAfzhD+lQvBbPk5XLrdjzeSR+8imDwZcdei
Qz6tzMjlkvnDBtEROjP09cERkQQvT7iFMOUSpENP8kNDOxIf+K5j1Pn5AZ9ABDbB
sBte4ule01t/IZnACKyeEqI3/LVOKhqP6uaxiqSIdJeF42+0XvrAaCIOclMlrQfh
TAy/siWcSUlRC4MN3OFqjJrhnVdWo7EYKnNquz+j1/U2Wgl8HJXuX0edvAK+XkjV
BbQuYrC6FyS79k2JcrQuHIV9fUwciqnetJ2RxenuBjcDCRpOr7BSuzzncB30nO+8
q9jpBzsL3M1f6+IZYuqC4VSE5mJhkjNspiraib19dhqw+tdPkZ0OiZdGNzWXC4gW
5f9UyfVJBN6Md9psnD5cXr4qD06sC0uttHhxhLblCymBkEjgPKMQ2/HsperrqgxM
jNFHasvXblyIDrrYqIIm1XuGPFFhbKpV+Yo/jisfe0ck4telyZD/8JQZuVPrgwGe
ZpImElA3YbDnnyf82eEeBJY6zS9K5Xh7g3mJ79RxBQzTYOxzro0O7qzQKkVITh8c
lQsP5ihbGh4eeQDh1O8qJi8hXYpWXgHJlsJXPXu3NPYIq75ASAMkLuys1kGvppR3
Y7tiV6MuhW/iDP9n+yRILxCIvdh7htpm9J9NcpLruZXT0XQZpElEepxMYatEj5S/
sAzq4fZBPcF/t+u9hYxTwRSJUqVUcJmTfZcaKaOuOB3e8ED11vyb6sxSP3mg7SYV
5SAmTcDb0CgdLXpMUXZJQskcY5AymV8t7ClWw0R4dt53yXRXJ07HYotGYFmQEcnL
0INFeNpZzJzw/AyQtxmRrbfL/2Le8LNU5V/aJUNKioU9cc/WwyJ1M3D1vPC5kROX
kd510YM68hfrolXb4J6AcOhL0AHwEmmn0N74Ro//ZjJW211umB9X4SogKxkJWRuZ
fhkSZNKXpzQ/z4Z8dYAqyzlMdcviDpEMuyYzluOseyUwn1x+uobhpLlbcta38w7E
8kChZjFbBCe4RJOyjDAnN9+nEtntkqBBiTQ15Vw1XC1Wpr7+h3MfPNLkPCL9ADdl
hWYTZou8dQfTvpiJ/HOGNIhajN52fW3T93Ez7tJbd0uvZDjI+uiom16tvU63/0K/
7emViupcabQ4G330Rogc9mXvdMj7QXbYd8ns6FrwWzzq0S22CIJfhnJ8awHqRW4i
v+BzJoM5bEcskvWgOeVJQthsA5KTBSupQSPkADp5daY9NFa9npTJzto9FrJzzbfG
SukF+64/5o/MH1tKVmWhXJ3fHR9a7S6HfWV+swqfqGx7k1teYjgf4pDbrMx2fx+3
sND1sAUQif4RJ7auhQvjwJTMc+IJmx95Eeq1aIrOiolxn45tXttBhqm5T5jSIR7G
h1vD787mbkLzkkBBPyDqFyNZr1bDUahwY66PgUUSA+GeEdon1Y1SdDEo+cQJ/IFH
rqz3An9OF+by2fI6KawL4QBpzhjtMqIP10DerobZ9Lv6GmHthRCpkT3+uj2f0Gav
xQupXAhZW+faP+n9OjaGLcayoiBL/HSKqNhzIri3crVal4hY4NFrARqevdDHko2i
bmqC4c04ZSjFgVInqFWhY/uHmjpAzYg0ddFkrugW1sL+T8YkodXPTHmhSnaIGCKB
NpRTvHvNx7ovqfHhK0hPt0/ioR24g8G2lxTC9qLiLi013PLFUgmzDnfed+OVMw9J
Fy6awhogRss9eTsJsWSNRCtf3I/50heAH+YcUCwD0Y/TurridYid/i1+nHXZV1ii
PK7GXYvgcBqZa9XHGaLJqezemzKzlyiX9BQAQbRgZ0e6DkAHMZ7M5P8H7VEU8R2+
5tJ+TfxEQh+yvb+gmxwj4NYEeUVM4UGy8kypffGQAvujyLTXxuuqOe4uNbz+M6n+
QE8RVnLIJZTd7eKUFY5ZrEcEtrW22wW/HXgBi1vB2aXaKnOIw6cO1aT5/o8gW+9S
zqHcgYYBjqRYHr0CScGwfnBlMQJbpcAAb6rDBYBnQd7xIblv9wex0QJ0fLwT7ezq
oi7L1fRV7Dc9Ah89Wcz4v+L+KSR/cv0IkwQYOMfn2jMJecPVQuvW7kzubjq1NPye
C32kmBZW4TPr4cAbpiRtw0Szgl62x65h6h9wy+mwyTvLtaskbvhaPZWLZxbcv7tt
LEvp8g4rvFx/8udBr5cTwlMy3evdfdC+iG3S7ngoUsRKPzqB/SejiHtMU1mM8JKG
GiytsdTLXVBqoR8O30Li/Fy/Qv9WjseRN79Qo211ptk4ge12jRRu01Cb1T3HcVmw
vRbGLpkhfW7j380fZnFUfrTNSZDvpYMj8lRhJANmm61bXtmfVo2Gc8WcDiy00kA5
pSu9TbjhwirHnadNto68kGKIb/4F+dUiLJv5ibckrXDdCoTvA6+pMA8IkCU/Tl1+
IVC2JJHeCdJbq6Wzg1cvVCalpT96PzZiT/EEGnkhmmhR7sLvcqPs9ltoMktpjcSE
PgN+2LDe9dHXonvf+b6rqc2R0X5CmF0ujZebLKo0t3Kba1PVtczl8MYxtDdrQtQC
9mMasZZpDuN/8TRBFgPAerAgWcgv97Ab36c+2mg8vIgM3s208bV4yJowUJ7fQV7e
J09JiKkePsjvnbactBObi8rI6S0aNMrHOfDQFCDQvfBVmonpoPZtd7nE/cTLitix
v6ClTPN/69EJy09Tvmgq9Jjidg7lSPaxn4AoPKB/KMo417pdkMCuXTEzIul5+9sl
+eP+FGIbBLxOCJ1tnRZYphoCMJcBiiFvyyAHqF67hwrynbRW9BTM4KA1lWYbNHp4
fB/8d0h8FUJyQau0dSxk+I/MQE9FKx37V2yUcP6IZOQd+H0WIl8GK2DPy84+xRRP
y7tmz0baT1749sZ4mMaRy7jLJejQu6/3uLdrJaKKiiZg4q95a5MDuJEkwBmUKuMU
ZMdqWj0MTkY78qXIfDYK6iHfNIQILoHIGPuh5spafT2TNfTdJBNXUcUMwEVrgGum
bmyBdsg3adbpTu1YeckReQUxK0K4Su3WOIwzjEdIErMkyLUwwJorI64o1Z0xw9Bh
rXYIeLuhtFgzPykkxw+C7081QqEblAgr2FuF2p4NDALiUSS5aoQ6JaLTSqL4oJLj
VxSDtNTZtfZv3CCLCwaQEzs59gEyNKn0YR3bODZY/u218U67H5cO5xurtmvVlKl0
sSHKWCg4YgNCANqCA3MbrKMhWIAQG2O/r6A/bpinwcB6zlDa/Ru/ay/mwz0iLI1U
8e/8HtU5axQnygJ3OSF4PYBkIA3VUp8WmmaKfWXqGDa9lumByuyW5Oni21f5UKHx
Tx8TCE54IdIN3z1psnXXmE+/tjGfBFSgkE3RtSPIiWY+ey+3lYzAvxGn2vq/pJZx
/M08s6g05n3WyMM4kgx4W+1YWxo4VCzSDcYAi9Nzl58ikmWw3s0ZmaVvbZUO5yV+
vOkes+S4YtIaPm/Z76112xScm8TGIuUP2NI2SKaZxN9kGPSaZsaMo0rezceRaazq
kxTxcOtDQxhQVZDPU0xmm2yfW+9ngU3ogbGzbu6drUHKGSO/v1iTB1ID5iDMtuwC
5xDqrsmKMd1LE15ijeMa41vITIaDz725own5j+cvK7flJtgM7vnUIakIue/7i8JU
QpJTx/Afm9Pzwb6Dw5rIyL2aGnG29icq1e+kWC0hHTfRP2toX/M+KfEjH+BoYRkt
5rfyrY/WEZQAhc7n9EqAMe/pxsfp0jdGm1AFpYmN2Tqvakr2w0IorQueygCqAi6a
6FdR6jpg5UMo5d//A9s9oAEWK6nVI7G8qJmmhyder0/GW9Uy8vx39NGMvOWcdNVR
DdRFhy1GR6OezSX5kpN2aPGi/OTSw6igy9I/r6Vj61Wk6ESF7RQR8uh0/zK1lSeI
ya4tZs98FIH/dRugldSXqzRI06KkdfiX9Da55Hbqc/VLjALaaAQKsY1gpcYkGf6G
vUPyq0dHJJ3LqMVAA5oYlqRX+r2II2V0YRwwX/OLp0E4wT9lY/FhIivyJXQOBQVp
ruFtickiyZpqh2GUEAHiMDZZZGBOg+0ic1fSMjqvAAkNh4F8tR97+bH6eCiOjAzO
Pm21cjtYW9YyVuL7alXwvaHJhrww/kSg8+BWTnC4nQtJkt35Wu4ILUtnJLFTm5WL
nAEiIxdZmfz21y9C1bzIOQOtfbPSZxHtFuLKnlLnmuZIxic4YoAbt7Vw34AJP6Vq
4JOUd4y3pA008Mam+6CarORE5rVn4uCzo58Rg85q5j9zb1Qlnm/0QAHCfFvbwFo7
diEZwjuaiHFnA4isYlWS8TNnjZQf65lxWqDQ9HF9f4qwjhWuEiZGSavhsQdVusEp
WFa8X6rN4gRHRG2Sa5ghdE35GUekBJNXVz0HarT1C6mB436uKRIHOSWufcXvEhyM
tBDE4XNbiP3SYKB52/tb/eKQlAgEege0UXjLvoejAioNN0xNQ+yA9n99yYRhGOin
TxsoIkY/DexXW/Sfz7z/NRPlL0iJ1/xe4f3qiy/xQDhbKdW2hu8XTYJ1LlHzetCn
72/ucUkSxCaPFvu3wWNs6BqQ4zWuaI3bH6+6d68iAWWK6HUSXDwVzbLNKu35E5ub
ot5ZXHm7iRUCyNX6NAb/7Yw4041V5Uhx/yUVVKM2Y8uB9zqvQ6vXpkiFCGSO3JMB
MslVczZPH5AwgOKoDXzcCmLr6mEr/PRUeawOn2a48+U3rp9DYQC5fgF7jSGXjmN8
wM5GrwmhcGsPaas+LnoSq6G1E2bPjc/x3FBcKuLydLrW1Rx0u5/Ty0WO0B2bM0oT
p1CkK40MfdhXtqA/pN/sLm+h+uj+M17Z69t0iRVpU4WgBA0f3B1BY2KvZWXV1a39
hatFLQSUwQ1q/cKlbpFX3DTZYAo0w8/8xYzTEqx5ejtA+w/Bqg4Pgz4V5UPbpwb4
1SjtuOwNgKrLjp8tBCyA8n860hagt+5W9QzNex4nM5/evd/4Hbb13jyYIDUS6vYu
Ej7wyWoVfDxlnkm17rE6057pysiHeMAmr8tlhSWPqvbI8kkIv2vJ1cT+F48O9AmH
UDCOkqB+a8JzoZ9OBYGJZC8ZhAlEqh/+13lACkgfUtaUW7HI7z5iqR4l7nZrk3EF
5mMGKhF2mFMqPBNRoix4NMfQ9JK/z8Gd25m08Rdf8vYTGrQNhI9drhHrwUb9qFOn
xcl80n6yhxlE45kXOfff0AVgE1AVD6hzI4Q9QkCFzUT1KAnGTieLfu93wT45h+gD
2RE5gmsiwsgmOWKbrOeJsqviAtb4DzaOWbLOwLv4OzVffI6Q43QvQHT5LcCt7mIT
8l1MldsQXnWJLfYzF/qqEqQMN5n9EFPCNgyCAEww3faZYExU8ZZX5uIVl8DK8SlA
w/ZWQ7GpEnHurgLD8gOkZBiKdahu7XkcVVlezXFnyand3MLg8OhCsxe/g/ZYrxO6
rEquIlAHWXQpvDYiQNLBq24AqIC+UEvrY7WSs0TdP0NLiE1O4mrJbtaS41DKjsB1
NBSCEpnZN2IoLrC1NuPOU4eP+rTGay2ROqC0T61Pmtc8y65UrSsAVOp9qP46rMze
puNQzEXjXTAQdjL7kF11s2GdwiY1GS4Utuvi7c2LpshDkWEEvwmg1vrzOFNrS+nb
NektOEDCaIbA80i0VgIdupAqIlnzmznCPD3FpNyD0MW7CPJdGtPBzj9YyJBPDOIv
eOU3LYNkvJT3QS9nSXdZ0wyuQ3VVfQajXRnzPrYSqUqvVuJBCijiF7GbwutLjcEu
5RqVjDHnUS5UCwo1uyJK77ZXbppdiWVe72ueiNdtl1fojktR2p5qiuMhKoW7QINo
5sRjrRErcLxtHfI5u88Xo4y4YS2Iz600v9FGVCOQsqw6fP/FsITOSwH73rTlwU/V
DpaNFxPsQTR/yNGeoWPMmXkmpM7zsyEgvtYAnprCQU6DFBnb2cg3ZEBcHgQApNRZ
VOkAahX/lnR/RPNBABN+DzEITGx8zAXSAOY1/tZpjsYEN1/ZcjDgqYlk2tXqTj7j
h5JWxjdqmK0OoJ1Lesq4nPOHJX+vkFH3dETWTt8OTyqhNj899z3epQmT+uDPJPpI
bnASUIQCZye3qZvXxVczc1teTYswFm5+qzGF8OVOO8oQE/k3IQj+lkClkLQxNBRy
zL8n+/trlNupjTbuss919mbWkmIri3cbKh+AWyBQxVQDei2tzmd1ysdxp24J8gMg
UeE8SlMkgLaUy3OyGhW5ldlQ4LtFjPpgoO81FzAbJhbEas4j9y616Y2IJs2B6s4s
ScLU+io/HwI9gmVXJF1yu3QO76g1+tiP6ck9KWyjRUMoh8YvLhDVpLB2fHZ8E2Z3
IYg7lQJo83eC5h2O5fouSJxADI+kpvW4VQrC1NUTr1nR3TeSscjs2KOtQ+i2a73J
C396Ph2r7FlReKKDx1KW4gJ/XqpWPElxU4bdZNj1qd7wciiqvNg245aXIkUAU5Z3
/acoWSwIqjQ/hDgwW0OdeyBHutofeKQBLJ4Vl0/hkt2aMSB/aFlMVs8fqkaPW4a7
KVQ5v+/J9N0t+mOf5eFOfp5DIxajMg8to5fMZQem8R0XbOVPuGZHA/oOyUIJF47v
xd3l/h6wTlx/zN/kP5VgpGXA6OEjeoPnVUKJqOHnhVArcuqpU7VcuvJVDu9OToYh
WX2M6202r8fkZyiXTu0V6TuXPW83QLVwk3nEPeRZeNVTAmYCJXqmBXhD9n1dLawJ
sYaGXrHyGaH2E1zd9SASv9PyrXwItfV369gXehG4Rhp1LVToCg2hcjvz17uUkXau
LDHIDrbEK/QhRzJ9mnCFv5JaAooOyWWQkp/R500F93DII8GJkPR9iL8wZpGjilUd
N1qvZZcC8g05mDpb5MHfA+RvNcNTiIOrpeS2aTHrB9nhP06qkmbEnvfFkuC1+RJb
HUC9BoqtSv2xlsLEn79q0c0/8ZGKCUBaoHhDGmbU4XNv7WCXKEfsxpJLsnQ+iSMh
tGKpWAC2lftEzX69ztw73KhsoH2nPp2NhoGNHkKZvA4jx5Ntg834MgYE+8EFSpC0
MH8CEfijYI4vU/Zv3seHa776wcYPJjFekHYZKl0RstcBAo2UBNcSyf+zm8VYGX7X
4kIW6v0EQuL26ryVp3dLnP/xIHybWUb8a28rz4w54701GXWV91lrp0ztb6qOTa9S
ajZxHXOsocrpfHI81BcPomnk364aT5smIHV6dUk9Rv2/J5wwYa3x2+qEGs1qA81l
h7UZN0WII5iBQoequ9qBndOU3U86nL4k6noT4geQP/rYc+AsYs+SsOOfCw1zcKzW
+CuiWPcd9h6OVu2pT8dmrTIOJV2oUUdFKqz543fR7opN4R+fvQHfee+QZ1HPB9qf
oYkEyJofIEwYefGuv7tYiybvTewcHdpKZM7D+J/x7EC0ZXx8h20wONBQQFfCHOlw
QMnkmE1MpizPm793jOrQkb7+NVBy6Qh12U0OA2RTc3PXwg1l1qZIF/q5iMRVw4V5
sDkbNjMu+qwf3nBXOErwoh0y7XbBg4yEY4jjCxfrRVHi6nb6d+6aYItK4dsH079R
ohzovwUrjfWra+PfzQVXsvY1O+caZjX4eAYK2qkOzhnrV2EC/4hLn2/P2R/edaF1
7EZN8cpHjO68QDEdl36edV7QcpwopBE10+vBXkc+mwT2oV4sjnmZVnJ/jJTZRXPF
r9r9fAEPvGOrYPQ+jWmFOxX8DYeJWO/FJYDibaozqFWbAjXMaxZJApsD06qFSkJt
0t4WnUUQdcSXT9hlaO6XV+e49lrnSAUTdkbYNPHXVJvTKekGc6rkAY+lHOB553ll
feC7Jq/7biaPIDAwDRVQtkTo7N2NKS0c2F8tuWOyBRrI79qGKuJN9xHtVAJvVDug
QCRiS2sS3I5BYujSu673s0oJel80TKpqq4NrH3wL0+ErpwcVzdMTH1mue2BkwotW
YC9GCynRfu54I1QRHgWpTTnJJ5uBbM5JYrL72G8tGnlqZtZn0RMItHTlAYeqyiTC
snE/YLVa1kcT/LW89oJjz5tvyu+Akoqu/jmmxFNapi3KO7F6/fLGL28eRP8vydZT
3LaHYIDwxCpsmURXYaIhj+/FBpZ5PjMnMFAzMe0eT2NYSGi9Lvh5R4macNi5uiiE
HL1UPqKkdeOOHGOH36fADrOhbLuH6xyErgaQXgJxJXjcFPcyuF9OVAl0oYrc5A7u
DJoW9IcZLMjg+GktL9SSLo+KsQp6py6FyqALB6KCyOsEfV5B5E57gA6Jv7cXBshn
R64YiYXnV9WSMZs9zK/ydUYeLoMMIFT2D7kH/Tju5vfr+XRf24ikeYlmg+BX587C
yzdn4vb0RExNpspx9XAzoPo6w6nXHrAUbQoLAGUIqWbfXkz6jfUsh4igTRSpIIpQ
cIroPs9Ggb3C3xhXvBr5yA43lQPoT3sqXvLbi20vF1wceplh7WFsmZHf6u7Az2SB
4zWy31kw0UTwfKX9KVA5axxQyWromIdYNiKNVX625ydkQV2eEBwYh0j1rzZ6FfCF
c4gBnj8eLLXuBKBtb/AVeMA3D++7O2Uo2h1YbsAPzudXkdr17hbG8sbU63gYXaDt
2SlqiXz5Qksfn5nBtldYdU5/taHN+2vn3PwwUsd2cCafZFC+PU/N2m/jgaUGjmJ7
1rruGSmRQDQE2NX1e5mBWdIRP2Eidk/xiIAQTMxS1KI6AdRE4dHQIfQyrvoNjppA
nzynKot3Rj4HgQd1JKRxsPjzgdfAT1T0/cTtG+B9NvYXYLln0CFW7KmnSgidzTQh
2R4TZnHh01idTMzvJnl+WA96Tqs/G2CAqe3JPO/cBTO1WYC2VuFu2iJjnLHlpCKm
CgJ9rZjVf8HnMJH2ku9Pr/P+LoAau+soKHuhDzrYlk1ax7xvwqocHeznz/PKP8VR
gXDf1OcrUI5KVPCRk8GKwkfFbq3WP9lYhmDtLbUhrrxOBiX0F0+DieFblsW4qeHH
qpcCkhBpX7mUKqeG7eCA7ivs4ch1t7ijhG4gZQwEWZuo9gQqT7aXeJq1V99D54yQ
Et3Qtb/xcyRFQJnddSFEW81cMzJTjo5ei+z7XnAGpNPdfMT2ajGUgyNre4ZYJSFW
qrCsTr1o5WZJLBmuZRRatZUfHSDqbL9Ara77ZzpuhRwj5/gcC01uIWqWh7xbTSMk
8qi0GLuuWF4tWJfXKaTQVYXD/Lf52aMhYsnUiKN0JKz7efQW/tpuJ+SCzNw17X7S
enMyhbuXBRLG29bBHhG7zqxnSfyRODrCACxa7E/xhubH3R0lGlC65KFl/N2efde1
8+mS2IIBY3PlJPvexp1u2R41X/6jnXgjCQqr8Krie0dlBekwP4giDxauv0P4pmFZ
PaZC8e+9KGCGWukMs1VlcAfMrdhQ65cuvRfBp6C8Tr/Jz7CYJ+LE2Zyy8eXJ3Oo4
lZpQWdk0h9W72Pj2EzgGbfuWXk6/Gvdy7hnbsHXZ90aNDWi7BsfrofO90Urp0o5G
V4hZ4GDvPj24z4gDgvD9cjBBiEkfiQuatDBL36w0hmRvBEqkNt7siJPfmPznO2N0
J2BHeBSlaUcD/Q8HJICgYny2vc2gl+4Qh1Sh8yMvBg+fIOwHwmsTn1gq1YJa92aU
sITGgg0zNqRMLnam24TGHuyJdnphI91R1Et3eV3/rMKz6ppsaWh31Ym4AFpHyO29
1bWu+Z0JV43jZsrh6KiwJB5IPENonGc9wyXR+8yYpndB9IP8PYdGw1g2OXtcg2T9
Qc6elalK78mkJUbiH/v8567D6mgHL0Ql3yDeN51sa2Xalunvs4wlSWO/sgklMi4P
/ZiAcNxroCqCAbaWPqvAVN2qQ+vNCqo2VdMZe+3vfhyjmDhjUC1lv16qzgI7y+2z
u0VTz3NA1Urx2bNPsbBb5ITdoir1tBZCJkvATShSkLQcSqnMS0B7SE3J6e/mUA3v
8fxd9xs64qMPNIogV4hqdDfXBSuuyu4n0ukphEFFFudfIqtNJJIHLFRhBqmCtTp1
Z9ZMf4Z2REPby+Nw/n2sT6SQkktas3JVHeaytsadoXkrdLK5GQyd2sZzLRS6h96p
QfcOkCAv4nAXso9jucwzbDW8VL0Npy6q2CD8RlJtKKUJoLUKTn6R9HNcj5h++Exh
lFLcpKD2OWeBE/WHbjpXtZ0EIhHn0yEQ9Uv5W2k8co9uql2xI/wCEuWc9bClQuHo
A816DvxhFegVBUklAzuo9GfmU2s1fbgbnnUISTj2WNrveTazC9aq0WFPFpGGBoao
+zNUaNzC8k13onYQBmL9vFyyQ6epbJpD6TA/CWBdGInUO9zo4EAOm3MXmv/7ac1A
k+ebq4x1MrdNwAHEs2Nyf6Q3bRtdYixQkBiU/yLbCN7TDcvbMyXpzffjgOwYHEHS
gI4eYfjsLDKmkNYxKfHsxstr0nTeuvSERy4lI2yR0X6SkF73sJO7cVe+I+fdErTE

--pragma protect end_data_block
--pragma protect digest_block
gcBhmwLQJ4gKWtnllmuF8K2tdOU=
--pragma protect end_digest_block
--pragma protect end_protected
