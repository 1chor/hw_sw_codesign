-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
pKazWZVbgIVOlEhiLDRQqtj+dLQe4M3sFSEQRkQ/VJxezOP3EM82ZGvI2Qh1XNZU
sclchBSmn7NA3GikPhQz1/3BHzI7s73kIKZbKl5WSxLvcy3I/YGxdi+4J7hkJQIv
VhGLBEW/y3HInSxMI2R19/01SBMxhIXIkRzTpUJllilIu4v7WRsxmQ==
--pragma protect end_key_block
--pragma protect digest_block
qsR0bB08JnogtfQqQOHT5Dh9qno=
--pragma protect end_digest_block
--pragma protect data_block
fCUHcyXm3eXH0E/Bt7Chj3NfGtDQoeTqQFpXTBtNxfJ2MNj9HAUxVXxKuLRMKJkt
7XLv7Zx3IbQ/mPZnE7Y70hpVvkaxOlIpZcO0xyIeMLsjYeEHLwsN3zgc+6vVmxay
oanXJu//nf109OUL5sqBsHhi80dK9l3JlEl6V3vFZLoCBNxZoEtYrZBMjuXWop/o
bppg7JN4qQiS6q3cnlo1qOJoXcsbw+840PlZsVhpsjJd0ATRVU2LP+/aOeDxEu2O
luS60IRPWR6bi+gEmzciDX1dbVCqrblgiAeaTAfy3tYDs62rziccL7vQ+j087vSn
Fr9BZZ6sJNIdwKiQgssJ08eIOXn4jEdY+d+UBe+huhV7knwGE2wsjWF2KK3b1Ula
AfRrlUFdq+f3ulQ22hGGp0vCzO07diXycIICOE7sRFzPUVgvEHqAOdPkt3pUExNt
s0BtCYFnDqGywiKI2d+e8rIS/gm0xWhv0vEU1wG2YfobDAytZOUS2QrjnNgvoFO4
MoD4bC7pxR/SuFIJN9tNlp/A4zpLkDLsmMY/vTSnGeFrl/IkzhsDvyh9oL+EShJs
7YyOsfhCfR4wzJwQb4D3TprpsaK7dfYb8VH3VmvVGI4x2WNQC4X7KzIH26CG52FC
Qo/Md8DKxC/78Exg+SzX/oqsZT7vHgpnR8tyA4aJSW5TrYbWABA/uHtUvFjBRy6H
oSiSIyCiC5eYMeyrsPlOdqP2C0kv83wFHir/XL5U0G5N1nVty/e9s8Z6WAtY5nTG
oylvzh5lxADfPMwPcRKR5bAJMKD/pUTDTB3wMx+PPFBfV/Louq+747L7qGO05LFE
C/HZQdoiKgQ8E2zLpD7VVegOXP+6Ktot9teM7fTWTAYFhCkBaHh5Cp4ArtKc9SkZ
tz20NW2xut4L8Al65t8hR+TKH8oKV/a21NG14K8K1SkGhbvF0GYDSglb6HKiKSyo
gSFnR3uUeLf0h2QRjrO2kbuXU5dv6IehokpAgayXPNkgCxPb7EA/vkUFqpSrO6tf
hgiSIIdnAUrJkBeIR9HOWeR7q4Kgw38bGeWgHfBq0z3r8eE4bwbucpuVj2m+fST4
Qcrd77zj1RVO4rM81ajyfjvzURSjFM6lNYCtoIRCg3/e0wBrDp+/d+RqkeVjmGBg
YxrOkahv7lNyInJuIiIkauCNtGtKxDMrg/832P9TX7QEzjN7ohhEtN5WcoRAFLbX
xpSwL4ZkXRYDnRyQxwzM0OES18UrzMTMut6DEPmMb0mR/zQRmOYp8CZw6c0y4Chs
vQtLi6SHeneRTP5MEybZLpLNOyEhWH8HO4rcOUV+xKVPGVF1/QJNscxtUIRdzAPm
PylqYlrRPzah3l2WqPAMqj6wR2/b7DFLlbWSWbv1qYid+2S5BiRuY1PenTypcR4c
qiquFXs0g1TLdeE6ME2U6pvcQxFoBJqVDp4lFDUO8EuKMkoURQYT0/h/roQ/H5Za
1pVg7I90HTMBO6TtGwXvKxrcSZnp0az36sRLMetd5KTEzTIZv45ZRMlVTb1VxfjU
4iVa/aMM5tilEF1Sq0SLBlsvvJiEXSc7fabghX1kW3vLQvnqbckcNLwpvcaxwM/m
JSgnyqfIx12YLJdq4DKoP+YLrrQT5xGBMhe6lgX7wfdN2i71zVkI+rahbZuRUMUK
Gtimb3cSSz9ZWXx/nCQfaeE9BQDbRB5oZZesJZ1AMJ/8xhK6kimS3cKziDJNhvZD
/apRYkhGvRpTf2GmIXRGcRFDUb0kmsTI/SXxFJK5f6nA8pO1z1bDbUppXkWco73c
gyLMDkpQNkVFumu+ntFSKOldx2mrZlQvNHJJU2a7+9EpmEZRPwbNabsVh0LvRg+Y
0uEXbf4qkjZfQJtBMlJKM6k8z0Qui7/spniLdz2fWuObGMuLw+sdtURHrMZg6LhO
630aBdpJYZm06jXqhaxZyavV5JapdRKDhXf4Nnum9ndHMiIvZj/sZVwyPIqSSRxb
patltxoUQvEaBxoG0CE3gdAjzzoVsfFxhUOM4KDEwzVZiPHF1WNx/pWQH7941ZyT
49sSclEhRESwfdJ1cvLEim0WHgWjAUVFxOtizS40GQSlYvcyF8su0OzaaBtCaXeE
WDbLLl/Tw5IAHJV5QC3zAdvcUACbr0LkhsQmw6H8RfYbXM2c3fxwjQB5x6F/417/
hE0vnqeDqoUmBB78aWHAZEa/P4kW2qLHF+5P0a0wtBQo4dFYjlhTKZG8rhltQYYs
2HBQKiXPSmSk9uhqBQksPTSHttLRD84tV/p5uLd4rBJnidWrACYUsaa+++XdTSUk
s9TA58rZFc4Xj7JA2EiSZBx/a7alJmv9EiIGbJFbftir2FqrKm+UJGWME1bDi/rE
+xo9zpsCuAeTK07jTdarxQ/RSt1+CPRSkj2QRjVHckq+ZIbCP0mvZ7rPU2/LhBJm
dusv1jDC64OllhIFAQRjbXJj/ibQ20H/ZeIshW6nzWyHgT2IVFiX9nPQZBscDv/L
UbYQ9JH/X9LsYCo5l3cpLzW1StEYAW6pue0Iir698mvjsp6GHwfsLzhGZD/sUxUP
BZcaVAvK3vMGH+XQSD0AV5hVcXThSPNHhM2SaS9PjC9MOq74XGImg4TC+153Gmdi
kgkyUmX1/W8CVO3BC9pAmEZMMnD/ykhwlNIbgRQPLAm9oxSuEbvVKzhSO0pDWaJD
WezTE/BxXEX5b0+TnH37RmD1C2C4ImsAbjKKFo54QDb/wABuEzJUPW/nmwDOeYAl
HxTqhsUglCjbi3Iw8a/BhnyQsB9NRwVmBsOsdQZdEgCzDDFCqtIc6FjkLRjFW+bi
rc5dy6c/qAdwGt1H7vN/+2DlvGsRAF8svk7JBWTF4IrTJu0dv3oSZ9i0h2GaT77U
9DzwH+r6FG8Op1BhYwIdNpJ0kfQTcO8HevsF1l8HxzMMsBNUMO7qNZVdQY0bR1TI
SHmN7lsgsR98YPX2HLT69Vwgkt4+iK2UUshxbjoKizvVMrXwMT2ygJdHLiz1rCDi
6yz+ESuekonWWtyXQHhR1Di3HKH6H+FxDvOuy0LZY02ZkrBf7lCYrgqS4JalaiZW
EFrVL4Na+l7skQHaH7vTNjQCbPj2Bxh1wwzRsMXsNZllGNsifmJxDepy/hpVKQMT
owhnivjxsHfT4f127qHNG2bX46s+EYPmMRmE12GJezVyaSqOkM+2cdM1xVtBRIwh
tuLyxa5bkUu72OwLc+oXDMAP/7kPkhv0X69vtOMxUYeHkYlVwof1Lwv1J1gS9z1b
YpNJekKKlj25i4OWto71GKHeYoxl3t3q1OjgWl+iHAu+pw9N0qvtKkvCvWaRwrIe
NBn/1TTQmgXOw8BOSRw3PJdPUhC+Q0bes88GF+8SVA+WkiJJCD6XK2vYGOY5/PcT
A2QzY3boeKIZj4rN2bFIDBrfh/QrrgAqTbVUACRAaJlMs5c1QK/UbccTaLUwimug
8+cWvZ7scG4W+mWATY66qtcuBSqo3lYSqGVRwLw9fFhSjncb2CGEz4cW6OHUUt21
j337Llm4oNf+kY2vCjZWiU2CsZPwBvi7oFWvhzfV0FJNJ8z93v0YHiMnrENNDbBq
2oRiyUFOlEDGSrHU0j8NbFf6hZqHaxY9wncMvN5FITONFokhPrOCDxdNv/2NnxX/
5MdmKE/yXxQvpAAHOM/XhaFT4fRzGVrnUYNOOwdhRtEeF7peqAykS2gpRXfCBsmo
pIXgI2Ss3zSmnHM3VZoMfnOb2zrYuHlzvV5EQAgWjHfcUbU8Tun6//0Q+M4IGIY4
gitW2043Eoq3D0zfsb3zs4Xz42cOBEo9FEZq9Fm7QYMBT9ca6we+L7tLP8Le+oPo
c7b3AotJFNBVSFKb8V9A/nRci1Hab6/qsc4p1UxC2yNok08j1yfgAjRSIFbIIJWf
s95tVHMJjmAlVjUELKi963WnwDZuHmy52eMH/gTNbmt5iMVE/EKdJxKsbzLODIye
ilxdgCk0xEPd5a8xmVx5MEuv20VwJFqzNwk0QZJGWMh50px8wkJ6/Oz8IONaXl1Z
L5yyFQeARRjjPG/RyRPR1U6J69Tkbhh9ZETlJ44bLzntrNqZeCtCcUpJoLn5LpeX
YVbV6jnIaaCAAMrm4Gsxs2wRl3pNjz2nTxonETY/zdEbwT0EL0jZ4y3ZrNMiY8Vk
n4dPKr4au06skRBhwwgukUxrOUEwMaxQYo/15BU++9mLUN3TfCpGNG2Uu6SGJ7wK
mTRVwe1Gns8gJQKBlUKUN5NvfCaqwVlknaHe21Ad4UjpUfMtJIYM1HdaQGxHgHkv
uDzHUixIF+qdu6zHA79QzvhxZxupruY/fATaktjUssQ/iqI13tt4hXmI9KZCjnqu
KyFbkOHXPeC5N13sP7DbAqwirPI0Fw3OsB7ffcGQ4lJ5xzccZ+ka1ZfQF4USnBcl
TVok0WOuwvb/DYs3bqihx62QHQJ3Rex39lTYHSr8VzctpYwkN39kB4TAVRmbRoLl
5aOpaQwdVhqYS1pnO/K8KNwV7bRnwhaSBbzCTIYCm1VIab2eD6G5l0cg9LEDw8rN
wpu/HMEYZOEDNudx8RztN99Z8HkvIMoIVxZQc16QZrzipcilxOwGn0YsKBrbkpjs
5lqOCk86pyTNYvD9xCFDHvqPzCV55rsGamwJ8lpMorRRficfJ5Wr7vcEU1WbRkXY
SKIxeuklVggF/HceTvEt9uT8BhIp4SZOEJfXSTtknTMDx58UxY2P0/WngpxKup5H
DxbuJaW4uQFPUkJ9ZSB/u0UfOf6ouLO6sLwBrBxJHXhLGdZHZEMdNMOzvhelCN/f
15VS70pnvc70jvGjQnIYCQDPR0D0KuGHdQwTrOQZJBwDrTrlg8Xu9LNFei4Es2Tt
WuMN8x8FWfpF4EOFl1Cc+GA/3kyuXkpSM9mv/EFvpQjksCoDXKk7zuR44fT9jxVz
TKLNj2qxLhsF4EuC6NkfAy90SflQZ6XAjW2UZhvhkqoLw7AMLkxsGk0xrl3a+Cwt
yIM9Utnb3e8qS4FIpzXdpOM3Z2yNjPYpUAkebcZJaYFUfuO5vu7z3LZcasDhwYLc
osK614MHZ/s3EBNpGBD7V94R5KYgfCiJG4+l1r4PDSYUkwNbEzQqjBsJIMgLCvyU
o5SgxXqXJqLyInXfSBRj7aWxEkASYGI4Tqr0FNkM3p3yAI/lT2gjhJzFMYPWjaVv
M9LahxCAcH2HgJNy6fMHAhXme0EiE8mczuqXFnE4gH0mEg3bMtNOTk3knedWTYu3
LB/H8v7yqEeqmKIrk8HXGewIlUTFnS0WC67K6wdJCDi+HbxoJZRTJruF+HQi1K9m
u3sichGGqBZ/2snS2WWoFtJS3Ok10ym79bWMuKeORq1Ixwty7Yk5CTFRKkhgndFi
Pm5iUSgEoEnQMKIkjwMZHstM2T0LVy7E/S++wPIlvw8gZZ8HvqUNHrmP/CmFO3ZK
3wcQu+/FO+LyUyZaoUWxtR8169EhqU588yYDwZgFuIEvYvaGu4C3RLDMOdV486Qe
mlUfh8oNX9wGga1GYN0vJTohOHitg4fFzkARABJBLXL83/Ypr5Kf2MEk4QvDXbf8
25v2/zVM1xnEGzO6RKmLj4z7lWWbAYkhG2I6SWrnB0YG7SbBNl67mMGDP2I8miZL
KC29ekz9c/AW2bAYTHF9YOkkoSz7/RXj0Sf/hQxJ2W9GeVoes1tOr3FdUMhgLsUe
a7jm4LwH0Rulj2rvMrukMPbqmDvFfUV3yqZl+gb0rDOAVghuIFAc705KzLjqZ4oe
LR0/GDzuqSj7wQSwC33xC50P6uqyMVENVXiq8OQYc0YkERh9Z7JxockrMa0qxoH8
biV6R6X8mESeWps0GAySmUQB8YVRe9GqaJyVj/A1TP+N5ku5xze3sCYLXjCQNkMh
om0Cj/YQSG3y11Ltxvi+9oh+lm1zFnmcIqxlgA+0emojmkVEs7prxEPR35YqvMbM
94oHPAXbaToF6Id5dHtN/uddip1B63++ZjXR5Tdfkl9HNeLaLakNd73wGl/34EyV
5eUIvZCpWo/b7P8tUwbzSEtjAe4VMdaiRYcTVRbfCiW1P/qHsWf8N/H6A9dtTRhr
JUMpc8tbCN2QWF2HkK7kw0/2Hg7sTPIgdVPtpdjcLSsJ9iFAmD6upFWvi9BxIPoG
GMgIWZrTTWx/FR9weZkR1yYMcsG7AFccvWv8TuLC/DXotdnpQ7uLELigr/egI7pn
TrjAeOqMxcRFDCdVDh00s9M2Ysqk71Bk4DMQf2uTdvuvGrJs7ebvAGOU26RPUtIE
29+l+hsFUZHXD0GZsp67fedOv5B+nelmAkv6Ke7QnkYyrpeDRqHVp4+t8bcw58qj
n5VUEQxmBIkbw884/roBY+AGrqafKdl3zcnBVoFlg+BaqsC8NsBOMPpomSrB0RP8
lFPUS3CBXFtfE+WItbJ8B4ldaZfACDI0nZs/iRftlvbxZnguvKOuKePHX6fzHvLA
U/EcRs6tjN6mtt67KflDywIM34eLfHJHuW5CyLIPGfYWIu4/pAQLYWyHLPbsZ8ni
rbixk+BRUHrl9sL2eCXvGZYLHX0RRFlq3U19+xx5RhhV1g8ByvQNdouKHAXDk064
aazWC/Duc5cjSOOY6aum8jsITyvTRuBvoXkFAuPk4HeFBggoWjhTqxzapSd8Yc5r
Q5BHwzoMLaXlkcWVJMtPHKJe/eO/m/Pp22mROCDMnoxmbCTSL+wVzHvlwrNVTYdc
JTHbGs4iR8xvBWj6irnsVabDfuD86aXylMitlqQdAIMfxRrHnRH3AIhyr/hwKdqr
FprFC8oBUindkQmfxEs7dy/11CZmpcatC9TsPbgtH9HtTNyffIjgiYT8TRUx/nY8
Woi5kJg46woBkl4HByudF6lN38uf90ZX8T9EVOFi0LAmwKK01lF1WnmbSkNzll3p
KEDrhYiQyIL9NT5c5Wk8zIA+SfElYIb9spPEnY6g/09yzgGBgb8xhrrRXWrAo5sy
DNhTt8rmy27E/znENmqbp0shgiuPqU9I9+9BMn1YYW0Wv2Bb7qmzLY0BDvuQoNHX
xk1LZ/hyImXdf5765dmnwRELWDctcv/9+F8w+6//tKSXf3mOSAXk0EFK9ot+2Y2W
kIKVWoagyhlkNh9RvEbIe3wHsYapRxN17evqvoRyi+8N9LtRc53Npi/AagfTssgp
sqcrqcS3I12KFZ3XGCZG2aqHrBO4gMBPD5Pcnsp755WpCfpag7iv+LNMNTqbCoAj
xlEj5vj4pwho8dJJr22Gp4bqE5XsEsttcxrDGeZbe0toLffWErVCQwFakiphddPI
OKJkaRRH03+46X+TdVjVmIrDRAjU1NgBeHWMHg58a9c/AI+X6vPchP2VmSPm2wT5
3LthtRh1BmxosyHihQNLEnUX0PqiMSLORQKsxeHW1gHPLTOfe+KtMReMi2Nze1df
sBTQsPI6gU5WAm3j6fJaGzR2AlbzA72+sWK+/O2TL/sGuISgqa1lD6wm4croxRih
fDhUL4usQRLVCHdwtdoALwSA66iAqOGQSWAi6Rv2TeQCzy/CHO7ZtZYEmSlPvw5i
4Ufbu5ONOQtU4eqDGB7k+21rLWGoYHuPeI+tKTuWE0VUEevclnxz8QsTHNWYjgoL
9fMDU28ywcODAeTTwry5S9w3RzXVkWkKGsU3hD9JXyJsFKVIBD26CJJD/7HXgzuU
7ptskWhzkMJePvcMT7wDcP1ZXl8FLlT/OtFgNMq5Dg9OJa5kiYwY2e1SrTC6GSYN
vY/hn3KcI1ZfkrBIfdYPR+/ybw7ec+pmoc8X8BoDvhysnfmOoTOCDwBs2E/RBPNx
9poEek9vHIZFfKsmCCmSiElKY6Wl7qwOLkYOEViNRmySlwvjg/gSk/9ygc1g5ymo
sqhUdlZQBO0TuVezq6t1roGeFCN5AnqHpTVNkmuUZCfXet5ylxmvUddIhGSZalz5
N31+bTmZuQbmzee3hOnpXnYcAs8vNb7+x4rJ+XYe+hRzgdcAwTuV4BSQU/yYajrb
7o+pujjyhXJFLOBTgcnZRhpGjSjRkUZy2C7ULB3TXeDOnRLlLTCMezr+peI+WtZl
o30jT1lm1ekBM0rp/Kc7+am4FDpdSnO/MmIS2ePgGfHFxXe19L+et5GTfcJnXedQ
Xll3zw465P6FVf9wypaMGLIT7edNK2rC68wbmpVBd6jUebkp7brNHk+ip778Twbn
zGlrG3HhPpV4h3xJ0qaOP/K14N6R/OmcG4mc9+eNeHlxy1ULybw62Z/reL+TE8A9
DnpUBP6Apgh8qiXTRWcgRI5ekeeHK5iVUMAoT8xA5mOm4HIWRKu2Sa3jZkBoG+wP
f72hFfhRLw1X2X7qLVT3IGJjI+its7AaKyfZPgUUvcHU21bIoW27zHY0I413HGTV
5BlkX8ZGZ1f+Sr/a+TAxPHiAYyRBVENYGEIPHElDfNBvgyjMadzX601BlHgP6tql
rS+8NflFpNgDVoXUbmOyELoa3hh1NGccO1FjmY2snD5BQZqZCJhfUvaSUQPpcIlK
LMjmq+5xT89rFzd0aS5bU/ZiJY0IkuSBGZXUZrmUYvW6vlAlzblGcpUwXPui9FFc
Ni2j7RtYp6gdBwR1ot3A0gsLNKGR2bCqlqLLzH7Gp++EARVHQEbhd541vpS4sWq6
OG9D4syyiOtpXE8nrdShFv3yHROuwITT6YJtgrvqX5vZZh2a/YYoCEXi3YuBwvZZ
NfuDXSI6q35vDOkQ+EiSxBZKrdVopt8Kn8KuoeD9z532ZEdqmW0TM8aeudmRyKDo
DWYXnXzVSvo2sXDDHOQ3zoY7pFttK5w054PvX+UOukf0TAqRpdwnbD4oNR3e8P9W
b8YhJEv8ZZRNohovSQzE0H632ZWOaaHNUi7z2TSv3GqoRFCMowRde1XAD6QG3P34
btffdoL0v0QWNsK/bfs2s/zMWyTRLycuXuMqxB5nPB/v9TAWspLSVuelkvUQgEzE
OOZAHvFl21B3iSMESXIh5P/gFW2eTjshMjeaTuOEL6N8tJo4DirEJxpjRiQs9sFx
qxzB6/7WqgfhFm0DHuWaMd44kzco52/L1o2vZvGxFUfQ6RgywY1Ya1YXo5ag1XZ/
GN3SNbyp6ExPSOyiWUmjIz741uoUG4oxuH/+2mEbrvPsw87SnD3qxKEy4wmudbIp
fUNDEW+ejlHmZ429QPWetU+f4olX3JfWEyYN0Tnzel1Vc2wTan6f5tIl01rkEEcW
3NNgo2Br38i+yWjxC637nXSCTfomwTGkrfL0CG3vRBoqt98Fu+Q8tcDHpEOryv58
rthNIMZNDL7ifqunHVA7vWDrt7dLRsq25GIKBZyjpcfeeu/dApReemee8OxyAyTN
b1kdYft/IgkntywOGjj+oyhcZr3lPQIROx3V1+z47xpkSfucsKnKx+O7VZlJ3upd
uy6et3TRh9l69vHP+D1rwEwW84+gBrQflgAS0BZzbodG4OtVgmadRfydThoHe8VI
6VTTxICxRwZge+9U3AgAwE3j+YdlP5EdJXZvmzoEU35p4D4LUMs2QiXmnzXaazYc
Douw24MCZ2QS8kL8DKEAzD3pmqvyGy2IgctYvWJRAsY60Zvjc6wb8ItfYHHnCw5s
QFQEFbae7mgar5sak9YyiBm43iE7j5LUYQBgJVQO/CJBrlgDQ+aRevoAg7c09RCA
KdzVOmdetuM/8QaqTrHwZ8PS+U5ze1XRUCkFJYDAYyO4oU4exiyFz2KUa/JqueXF
DKWGwsHl9oCHyUCCMf4szPVQuFL1AjlrKhpaW2ITz2vjhVICUI72rwmsjEzttNhC
St3BKPiTsNh6B7j1kyU5n4nA3J7AbN9dZaCZDgN+r9ZAsaTWyPm8o3WL+AKQVG+0
fBZn9OkaagrvE8kvQSZuXaB5R5c8vQ06/I10j9nVKPvjCURFinRvu1HCcdq7btos
RKzD7aoAcMK5Pf/6f4fyFJhXaeoI6SwjQdCAZO793rwx5NInXHiGf8NCFGvYhAd4
+u/1JDPw0qABVDWaBXbysbhogM+pyQDy+J3QCryClsAkE09YtOHLu0avV1HEOMnF
FrWXne8yON/yFvDUtMV3AaF3AX3+sZDRx6zWwZybIR7aKL9uAJZVxsm+RuNhASYd
qtP5hoQsy3lm5hUBoCUhsZ03bLXTLnIx2srKxiZQBFIukWl4ZUNUirSIq1xLR7gz
nvG/xgX3wPy2pCi7K6+rRteG93CQ/QteWL4UCEpwkTCcsAFgDrkylvpIjVhA/R1V
YraOnXrHEwW6I9m++vTs5PrvJhxXDEfBYuiYSso5o9So9hVHyqlcukx3Tko2A5oc
uWxvGKYbbqiBA57CqYCm8qbJQ+3EP6m7cjFU9xI4qvoSVtsLiqRYhFCS6fCFARj+
BOz1iqtmXk3bpPmF7sq9FZr1lfIcFrf+JWC/yI2+qDk4x6GLLfMjY8vOIzdtk6AN
GscnVVaBUQxV9E8ZyZvvYaz1WKsFzSiRGypAyjH0u4rbQahVHCz6zQPqQOHONpC0
+YwsWbC5v1EEaMx2jfXO58xJXSCzFkGnIhxsyq/IGOmUuuBUa7pdQGS9lS4p5Pq4
KXDAvvPFtprIUHYMT8j17uyadAQ8+gUrlyGb4r3fnn0f4vXbJ/NGugSVkeZ6rFGU
u0wuEDrlRhB1/48DOJ/O4c/K1lLIiTAscTHbVKfm+cGW8pHZbXEjjqxNeGOeQW/v
uGLZQhNNUaAuKT/MBZbbtsLEitkFlC/dn7QCSBwTracx7M8V24yLTl+2yp6Rvm3I
+TzwPFDr4U9O6pKBYXYbJJeffLTFgv6vPax4kFiSY5s2AMWBINGWQB4254raR5Fj
Tw475GZTvR2TAukfsjdWY1HMCQ2i3ejQgm/5dWRjBJmv92fljeF84zraASjICMAR
xBn5vtuR+B882iAyi50aMM/hb/TPEaXvrCYWM25jSOw+heGoI7RRpgarq7o3Swmq
JFJZIII59fFjjKV6TrRCAAM9WZL6fJtJ5I3abthywrkclho3ltsNqee0O4D42ecF
PumVH1j5wcJx7y6eIoJnDb3JPuKSZt4/MWJII8qfieflWP654uGbN1loSj/CNwNp
fUdqmdN/LY9E07gNEN1ET+LUrjkpkNh3DrrBuU257LGQHCFsHM1QCpsvE8uTrSd4
rrT0K/Tp2yIng9feon/LnDt1xiQgjtp5z/qmEySyb/L/8I7XKh5ahVBmJAZ1KW3i
I2KoqZjzeCiVlsiwDw0BV6o5OxfD6dMfhPvswxiNhkTj21kQwwC1j1rSr5F1IVjN
aPG2RhkQ/FLhOCNyTpjQlSgu5YT798A1GFyW3flU0yE7kPM3/fvW/tm5Dax2naAr
HFUqmmol4PmxG5RnbolrOIxRwRtWSXzdDBM2uOBAZT372u/Dx3rFxKMeQYL20odN
BxIkdszUaxCI4bIDU/IWBHDWmEiYHmoAOF3ecbrEftOC0yXYEhrRQD1ZY/Elkhzu
0RHQSU6ZXVkBT4NZdXS5ag62gVtpAMgPxGRC8hjfaTgbCsJma4k7nTpLnN7b+88o
bId01vK7AKzlSU4lRXCfydGq/0xj2cAQi+ijgFhFN/G407k1bdLGgxUNc0FEor+5
Kyk3Bo6jRwcSUCSsmgMtbD3IRX8eQhFHd6r1IogqpWzQ0vAot705Q4DTS8nYLmEv
Sw+DubgiEVXsRy6Q5jVKhE8fTUB1nMwEpjOCLXCNZqcmKE7RpwZXrdh3kj+F6eqB
VHOZKyeWDuXg4T1/8agqeE29eMpbqgdCEq3pL1H2P2zqTUfDN9sVWxtHVtf2KQme
elMFSk1EdMvAAoYiZa++/URRa9uXLUiOPaJwDrjxoJ41XzWsmej62V7Y53EbVdH4
KnzOAeRyQakpB7HDSvOFXkZ3jHMbXbyyElD3p0DCjS4BbOw4IjVcocNe0nH37aci
5VQk3PL69HCai9fip2SPzB+AwTILurGiWECB7y7JLzo3pFby0XCixPxgiXmUPP51
6zgZqJQDSdNz2ooDb5l/cJQsGZc7MoPGcX6L/Wyf5QV8qoX1YgKkxlwwyhoHlc/U
o/vbDta92hDJCawH9T3yVTb9z56QEVcsZ00KXI7vrHkHAwq6fF8HZXAD1rB6T/9H
WX6cR8LbwpemCd0rGudolyocHU+NBwAZCLSifN6Z7xs6t6VZer68XBU3hVt1WC33
9FRl1CPjcTWk7L3AVZJ2AXs0sMkCY/q2U3C/QHKEzZwKYep9BnTe5M7zGzBfTV84
6x2XTNJliFNzGUroCLjU8wD2uuuPI4rSkbrfv2kbiQ95arv/uf6JUeki/hgnALmU
VpWhD6KN2m0LMAGwtIqv6hUlxa2VMkzXeJ4n4cHtEB0GPO3LFptz0vYerwSzdag8
jhneNHDej+AMRJZ+HUqaKlpkY7B049Q6ijsNuPUE981928MIOd5tQE4MY8t48Bxc
5NgDFwWYFemUNdgZxYleVKf6DZN1tFP3Nh2foF+islqEcwHxhebSyFsPAbgZgXh0
O1MPen1I3XYgFwmhUOQXDEz6l1W46vGhHYzNLNnbOXu59pDbsMXy+ea4XmxU+Gn2
cpBf2VTQ+bEeezcx01SwU6HQaZaE7WJ8qW4Scu33z0nJ9xUo3zzONpNBAG9hHY7J
Mwy1ASJOkuSoGlon+vscF8Z5yH8Ux0n/XEUB90ktmqUtr7Z4Y+rnf92XISAclCZH
mY6mAKzntfFt8zaS9BisheV/9MG4caVJTkMOuWjALJcIjw5KpUwNu8wICSXAIPQM
SEow3m6SDBFmU9+yfBUcJeAR+rSf00uT+zgHgSAg6tlhwP9JsD+MD49IB5DreIPq
vAe221BI9NWZOgfSGtFnFmbd6s74NyOe8XmZ0NFoenZwRpXbW2gbUBvf4Tdk0UZy
s58iMJiNOA0GEpPDzl1uUxZ/cq4P+aFCJe/L+Pd0K36SAj1AbzJcuxydmDpcXUPs
r/ccUbmupp75uCYLGbuSr0D2F+8Ub4w/djuW9bXU2quHSmfISsCqAlZ9t7zwEyiB
w1FblbOh2DiG2ZgHQkMxLwzTiuPV3ydKSeENlTJgQAiqU9ujiuaZLNIjI/SA2Ko9
K8PQglp32CKrJ1Qv4QbvrFlXXoXiCq3x1+USRHywyQkjgAQD88yaHy0DV8+52PEH
xOO2FTGlSx8TaDeQ+Vsyr5qwx5b5hX1YL/JgSJka+Xw5Lx8uMQqPwnPKFjWxI/Ep
82kx/adFv5gp+nQI1QJmbUu+BjTMFHB5tWwexXn3YwY3bhy/OBjOkIlh7StdYpcn
T5SEVxQg/GjHIQIL07SV+4E+tY3myGO8votsUJ+F83oYNtpbts5Le3mNwmHW43w9
t8fVxD67oBJLjRWk9lNMCarFYdgTHlc8/7THtUwrrR6zAqyMDaSRiqkYYnDbZxLE
DMzAGrE3ihwSTg4FoBptMPN+sTd33ii2JfuQjsb6IU1ahtYOWJPanWXKH59A1OhU
j9yJEJ3zGjEwMas0wv8rbGJ/uJUmV+rBi7GMB11y0Aw9B/eAHhhOyhMKY2s7b4rB
UZ7T0pRomB6OhmLBx3nw9xkMxt6/OX+IenSe2r3XuxBb+oLYFVp+8dYxsGmcMzWS
wZfPiLxlcjKiFfwCzt5VRvrxh70bIf9dhsLB8VlBWBEKr02cNbgTRZzdD6gDH90h
t5PUEbHTb45TsD2C/FJPg2AZ5Bfa9I/g0LQyCexBFY5oVV/Jxax3Ady16U0BYyGj
7/ZkcNZ7vD6dvrC7r/COAOtUNBbwKG95yIkqOQOOJYhqrw9xV8+YbkvmSUqWyzVy
PzUMSNj/s5LdolrZIElFFIcUxEn+E1dRL4xE6MQo8UBqvyvfKKBcKG9FsqBhYyzN
tre2ubxnM+wcq9Cz9YVvXQvifsbcmvY0D9lm8kKY31TznFLBbseJu84cjXxG8hUB
blK7b5HDRfWlmRp2Xt17HWY1xyATA6XI+GHl8hl06pcn2xGeTQ1e7QcS3P7ErHKR
kft8Qv5xh/fv/aetsYclNYWEsCMAC9PZU/GrIM0kYBEIdlTmAR9Q7+xWfCNUOWvO
Q8U59fmRZiLLf1iPdpiVZEHNtz9qGKvsHyA1I72a1hI7hIRfGUg25tEOKra21nXu
71abn5sZ23QQ5sDpvxBldJSoyUmmEjUAkmheDqZTlA4+2Aj3/Pd5h8oLib1qc3k8
JA83FtrV7BOlajF/6TEmr2CKBayznZoh+yO5hC0ttGCnBK5H5luHrBDRvsRcWuBb
S36JCyfPCyY/UdRXIA1D8P88I6O7y7+sHMXAUm3lQEUeY4rPbBIGbzKGwwChseVP
wwwGqf1FKya3G+AtA8rcyrMeOMY9PO6JI5RMup9K9Iews+D54uWvp+IJejYthZ8/
oQOmruLYbl1UAoTcUE3oF2BjJJrmv0Db4+WOlMTnTGzPpBM7Mtxtg8SF94pfu/ys
z+EUnuPdUierOJG+NrZFjQ7GemVyi5ocyKD6ZdUV3N/KyShBRiqvUf86xY43Vdnc
4hO6NtLKTePV9mSq5IRSM07vunBSPEm4zu7/uY46zGZxo0B+f4vLslsQd6WHMLE5
q2LgzEQLTX6AoEqqXdPwlqzpQB8uXQL09vzy4WHcuvwba0IaJtfQzYCVs3bwQNTk
MgCHAe1EXAdo55n6mcb+zlIhQCA3ZREb5/QsTtDh6aF7DXBSdYPI8VQHTX4K1HRL
64EV7di6qdWrZNQW0UymVVAy/Wa6Vyld7XO4rtGNtkMlusVL9h4Zwib9O8+OL35O
mfYLMC6017u+aeHghS13sbmKXRzIAjnv8E34qbQ4f6J6UiWzlI8u1JhXPFGax+Jj
6mkfnJP137315DO4nHVllWs1w+ME7zzI2P1ZxhykK9BofrbfHnryD+vMhRiPzRmZ
v3sScqvXBz5dAFVBdw0rlrTsN2nI8CJLVw2oX7ZmxAq5n2FN9M742mOEh/FD6Asw
+PljbZorbYODXlRVvOdw/C7ZjSo+mvjNbjqf/8LPUcPNHNmsz5VO0mGQ3XC34/xB
BenMNNwiDMqvzHjsZAmI53s4d8k94mtc4xyQZno1koMBfXyQ5VOTc+EC2xlIq4YC
O92uguSb7OVNwoOlmytas0eG/qClH2H/LLu5Dipjlf7vxY6cVmu0tlzIxVUDWK6A
yTAY0eaCY6NK0ea46/Spq3hZDuyokE1hDr7Mh5dYLNK/m3MhMv3uuEVlgOUnvBeS
CaqrXApBvLzogOCOyV3SfdbVY38bUVJh40gWNbCoyXp18G8d+9GHTIyFO5Nta/AH
EJOO7jR7JsaKiPcdM9AQmxrOmv+Oypa6BTjNlxsleRubMX2RMUc5YutrvEbnS14S
IkCX5OKl9jX0SCL3r2xxDwqFk9bxSp1okM1zR4MvRpRFJY5YNlUwIXqUkqgkRXui
XzPQZr4IXk96VnySqT4WoPbSV9HPfZVimEyZoY/Yrsu+yJvFPsfyIG81yAWhH4GV
nMdRCzg+j1R6hbEjlhmpfNdUYrwHhZZ2TwgkAZJDhpytoaX1eK7d2b6aB40zPbJ3
yc+NM8KsMCWQXi1BYTMM6VKt/cUDP2uXYhtS7MfjFHhpXebPUhlqfwJ5CviCzLnL
0I1cvXtgdOfFlk/Y18w5Lo/kb2xwtAEMdCLMTcyiMjjH/56WdBz0QZBxWoix69tV
e7MdSSNWlwpsHL/IB17sJYXSUoWh8t5QuuulnX21zpMZHq+Oc6P9+IIgwG849eED
TX7k6oV00Q2QYMswwdvMTa/6WsJQrfAvoni9YBWyAioRNZnIPqn+cGTTDxpNZVFI
MDIH8uh82RvASooKAS7EG5WdPztOxLBhbT5Xd2scQVWRvrwL978p3fE9vgE6pWSL
KWZn78Piwp90tx4pO+zhwwR2FldH5o6W/W1bRU965BbxQbxLzOsMCxe6vrZ2lgMI
TFn/SJLGjh9HVAdRowTM3JDsoCNmx7hiDzBF4rqk40qtr4QkozdkwxWRqEQirWpz
ypupXrVAyEyzyhNn5oftPJRSYLoIblzWZtu3Brsx0Cmedq09KuwUTspOPh/GXtcR
JSNw4ah5G4InxvRRIgsx/X8DMjcavY/jdArr6RKP8iJyezL1DcwV5z7ks1yfLTHD
bMZ/gVCi+gab8Pr6K6ccgg+fB4Ig77jHYW/6bjBRG8Bqdhr510fXofZfO5T1dqZ2
tMeaMzpVMy43rLXwAsZGXipmN1v/slyneTgKN9nSQh6BKQdvDxpTaIExMoy2VwdJ
v6/e080OSM6bj9OIuA9K6d4NZgajTg3sZ35+STH0aHVKWvADq+AN2Xw14/Fro1SO
rI0EwO021dzCcq2tyvbKGkQScN/f3a4ND0wsGteIEN0FxjvJNW1f259N/OIfAo4l
4qhXy7JUgQbVs9jBgRG9ZeN8LPXe8Hq2uzj6r617i0PJIF1rBCr9oCzJjq08YuOk
aVW4ik5RMvuT2/0KukyzacuHXe0ASY8ewBeISjJp2fz4DP0QhV0nc+y48Y7ZJ1Wz
XxbTPg9nG57aVXXIySOyAvBNuxB8xLqqcbmdLmGXPDdtg5oBcTPRC+w21BiYgWTm
A5oAwcuMmBP7egRc9OMCvUVRvIsQWYJstA5eHH59JK0loyTIqdU+dsO1OtpYhnnJ
VmJ98AYU8jRDdettlpRCHJ0Xq+YSXI09VhVYSadxPYdydGB+O7R5JGEHGZH7etUd
H6CFbNaOAnKOQJQ1rCvOmoofhkkDWNqR5jDRa42f8a5WPbvFt93yG/KmYfuQ7+WL
jdp0lL36yMEdXGcIugGEIBMFrdimsUXPr9p6ElJwq0p95DqqpRbAc4VRPDcu30sU
XnMGWNxvj3qjr4ld69nRgyeT1xcNpzw0GdomPD/N8S8WcrZbsreHDu/PHot0lQZT
fVNhpPtGg7Nb57ZpsVgeDCNHU2wYu4CYXYGE/yq+BplqSQAk/pS2FR1LFvS87CI7
b1wZfEIirtU733ZTmm18KULWz/3e+iQ2NDxbgOrNORwSq60diwSBOBUvBOFZ1JK7
l9aoi/1CpwtZh1WYtkuQN7bCRpWcLO7WH+/y5D770N6MCybMhM+fyObF03ikO2/M
e2WVsBLDnroBMY/a8XnvV/ykTQws8eDEtHLNPdh2LiwUguL47ss8/cmS/WcjuXv9
sczxB5KnoHYUqonVa/2lOKJ/XfLJdnqsFebV+YA7JATNBlrYGvPpfpmTBKCqL/TR
nZJ1i2xWn61th5XWaKpYh1sKtQI4Ct2DpcTKSQP00lBh2EC+hqwR/EvAi+ystos7
duXDPnlMLC45oSiyae/+t78TJk/rw2RYy08QuLyto5NP3jCWywDp+tgFMaJKvcfE
bABE5vOHSxbhAxBqpN3dGN072Hx6KBxpuLyZcVnlCbdmm33g7wwG44nhb50MN5E0
vsPsV9DjgmnIExr7DmjkhJF9mfl79YlRztLZ8gJ3CCu/K4X8m19cXw0vSRG769cO
0F3YNCnmD9ELyYN5MXpmpzusona5GfFzHG+bgEul8Y0aRRXt7oQPGjjv9tvtjIs4
B0O4HDdpGLZY9O8nlBJMbHrIO7BJg8zB8kPHCE0LQi9DVAmxG1XuRn4Snatk01sy
c2vczU8xvHl3syJyD/J03z3xrHKOgPBxVmblimy6fbjC3vPESj65wE0QK5UgjIcJ
MyL3zLo22MIz3crHW3nWeDARKO8Ckem0pDJ4irzjBsYk9h3u8dQIlDV7HXVHTm/l
2k/jktLzwKHkeoMS8NG5zkZwX+cq/bbn/9W831VAVvre84SqFRV4+wgctUkOUqhO
S+Mo7xVdYjPmrwCj+ShLaEsPXzegyrwNA0Y8qivZEP44e0h/2PV0JZQbQc5z61Md
2iCl3WiW83V8OFGalC4QgKopIoHDSmywF8QFFcZIUJEbqvcSEFFlRbyakCMpgACc
vH+Gzt1vYlGdWxyoK/BS3Moy4iDkksDZQsmTN/9tkb2izZM/8FWCP5bT51Y6183H
RF+w8iMiVW+8u0az58Y1SpfOwP61littjAS4K8y8C4jHNlrg9k5qJ7T48Aodz+E0
8G1yvUJU/xdSCbnM5/boWAjXWTVdqC6zFQATo09LH6LoSeyBc/2hxS4IQMUPgdX+
eUAEtscIAFdBb4NdTmWUex4pdQ6ry345S0jwSGJ9VNkcFWkLvxJc3toD3Yffpjlf
F9UoT47iz6haOcaZAdYleUPfxNygyY+ilGMyZz47PjhWfN1hhgVOaiLqZHrf24Px
5dU9Y2fIbVOxullPTQCCf3vnfIcHai01n0PhWOsmErW18BiT53WbmHaigl2j21dc
sCcWhJPrg0IXg7YEOs1ZpQORKlXNPSy4TnDTDC2COWgI8m8s/FE9FRq2d4rhgmyg
XCLbcYH/s3e8caMfn6tUlwC/XK8ow4eRZHZuv2XoR0IU2lc4UaccP6O7e7CbD8lS
39JCCWnn1+Ui7Fi3/f+9Mq0l8mSrPTjP5QLtkOxhJux2ZCJGDvC/MvmAI0s471lc
ldtthjVEHixmSz2789SL79/VAMiaV3K5R9PAiuohvj7yFhMCsdcqomAJN71i0VBf
rP1RDbJbWWa/ny0hpC9Q5I7UGmzRCBd+YNVjgSAXfeqfpyo4u+KPRVotSWc/Q2iT
TYY4ATXWZZ4U37rniQsQqLHB9I/IDLa5L3rySvckZjji/ITj2qMw7RWIoNM/Hbg3
duZdpCVf+8UB+6WYjLsXLsQ2cYvseBGR7SqdX5hUZwzV8E4F2RU6DPLNjPm+h4wl
L1J3ghwaVLCwM3Jl8uCDsPgJA29qd4I2l1myfPCDLig1g9GO3h+1GItHDTDHZ2ok
vU7nzT2sxQ7XA5UGAGJGk6zFnaB26mKrmbwvu/6KRDo9KvlQOuI/UBqhqrK4iQZC
IUfhs/qDdDXswEhtofr5MOSOThqH3Dm9wN4icG1bp0a7DKBfs3UK6FIm8mooN2VA
o2uihwiz+QPXQNyrllNUd/4tgKeKaZxDMbN08dyJa+iKZ7CQc7SIEAJ82XHHHjHG
IkHn4c61J1Fz143kav+RC6GxA9Az5/gqua7JGUJx0NRa/BVZtDWU37iEmdpARn4O
FKSsDBI+OMaUxC23I9V8XRNWt5xI8cZjA0XyW5sRpCxhA/aM40F9kaBK1JIxYfGM
hlcvs00trQpc43I42ahkh0EcqYc6W275nZnhh2bQDG45b5S+qSICLYYxsWrWMcby
sk204IZPxsO0zWuh/8zGYIMcVGJk3HJtNmAB65Rp93PLG0IL1lCvKqLsLUH4bVQ6
GEhkKu7f4zok3xKhqYXPcNs7yJW2paKPPsZYgUdypTBKPEV+wJ2NHaCXaLa6udAG
GpM9aASccWz7kABxGZL+RsbpgiD1N6X5ptvA2gx8+HQTBgH8DpjrfaVWVc2ffrPL
ljvLCSx5CoTLxnJVdVITUeh8kwHD70XHWGmbrkAuYsjjKdhyrc7BixjROrs37lgk
kPB2X648YRyFcIPRGxni3IaFyBZdNFC28yqN2LXhbNUy9CsyAuPaq2TfdC5yAgZp
23mDa9rgwVbz+pcjlGOawo0BS5aLGDm5RPzfVCNzyu/ewzpwoQ0xTWOPjSNkgB1y
wb4RLw7tBkf9w+Zsw2a5459tl3LNepWWDbRuhS9KUEPtMZVb2bMmREOCuLK0Z8WL
z8+sU9rNFcuLUd0FtlpGEDs/RUirtDA5PElYWuJ86E8zZd79POIwOck6T/LTdFOx
6uQ5z4zPcSsZ16MxDk+XYHGvLJM5/Ix7aIBv20WDMAI2BRBtWw1ShUZqvuZ4IOTH
Hdor3RhfEsEUNacwidABAUdbAAuEGxe6dtTEc+4787/d66L9M2ysoNuGYybsJ7x1
JFmfdXStLXIqbwO3F9eFgoNq+XXJ9r6yHZ0IR3emQQiBO5DaUhBGL2tSJsJxsZJC
qCk73jI1FOiHQauZDRShvgjsRJxaIkxepQ967Wd2HFVlfYpOz3oG9uKU818EIg1y
odZELns7ETSxFHmopb8mJh6KwOLZFTX4zNrnWUHo9SWmQE57DqySO6Fxb0t7Vy2D
QfbYM4LcfYS17NVYSFHai6D3xRjBGBgbvsswx8F3As6cNZPQ+u05B66KEtYAOvbS
N5aB5gf0ExPA4Sd0zhzbvzHEo0emz/T+774x0aOKUmIotBdL9i6wt+Qj4q7oUJL0
5ks+I+8OjbpPWYE2OSF1jPlV9pPCcDR/3wDY6AKlGELnjq2FFpeeEhGYrnG02Pwv
fnN+j10Dw++sVd+0eC/Ua3ZAysGmN666WERq4uBFigeHcLdLuDoHbOXdQYrersMB
HirqWsP+/dXtDxPLn0f2HaPb0j14l/5MZ4/i4BGSFK27qGdBtTFR6/WjlU/Nwej7
JTx4sOGFRJ/rhEiISpuvC9wSxGOzE4WdufH05eMqWElq2ZJHDznYwoY5/m7v5I4w
EKzkNkDKXoSMkxMZUPPnOFE1Eyg7+LPBNRpLe9ZE/7SfXnpxB/T5iARSzK4yDkLm
a8sWnh80AadjEVbvK5+a3yisBfIUYQEoxKG5NGDSh45PHmVRow+JUriJ6wbC3SYj
5OoOxjLreVYgDY/kRMuiJo6FWU4aCgwOoWOWObbbsnmG24rsP54Uy2FK9vVkyZJt
Cr/bw+scMaZwO3XqpCu20gjb8v8KVfbzLNfYDZhF0oc5yGaXKS2aSEogaEF/T7Qe
cb7GvlpcbGX7BqB2Kw1kIBO62WfRzrPoxZ0oUVuMhMaE9qTeXa3FRlH6K+/0280y
FCk+/kt338oasZLMOFR/7agkVfVPPjoml5rZUDH+Z+31LjtLPn7dhYIv5aC159Kg
GroiIFd+zU8R3S1/tkgoOFFUyJaRWwOfFWx+BvY6AnoQFyURRgKKfENP9yjhLtaD
cCTx/yLg6rYXJMhHwhZM9Si8H/v3NUIQh2j7zQy9RtlrKlibKfsbV8lypJmRSvUi
o2IwXli83wtRak5378rTvwrSv87jHA3whcoJCHtTqIIh5QJQiSeeFECDB8I0WJV3
Ea9q/ABZelN1mLF74H3g2L30SAzsbrBP+4QkSA77Hm7JXikWdndCCW2imWQ8SiBV
RAfe7/pd7a28TOwgWPoJlG0Y1jfgk8EMcAPA0a/EqDF8auEqwluLN4fgQb5H+p7F
OlNe9juioad/5bqXH/+AMyGFx9tPWwqrEQ7pi/rMdiucYR5k60b2gnEvm8fukOiQ
PRJi7gTcivrPMi50B3wcKAE8MbQTYF2/66Tcr9Eo/gZHQr5hfT+Xq/mPZY1msOWa
41dmd1PyvbnSUS1exI+y2JB+++U0og1PbU2Hot8Pw6tTneh4Yn/h0LMcVwGRraUz
hkLSq6E5ijFc+z9jg4fcj+z5j6leXLZvC+w2LTT21Et6BUpzL8KVJocyaG1S5twE
O72WRrVjscupOwFQ1wn6BxEalFf2bCKTTLMJeZ3sVVTAAVyPYfectW0zroF2K+Fl
FOHZmjIRTeHpY8E0SUJmCd4HYCJqrIo6+YnWHELQATPn4G4ie8BflUYNabmJe8rM
h13lhWe0gBVayTksRIgKr/nt6djijzDX9H5Jw+bGSyDzFTK37hy3Vz8gXl7mq8N+
OqjuRhD9V+8uQWLVezdQ3OcFfUXs2zYatbiJaGAKMBCVaL7bI8iYyCh0sdW72fj5
px1atMqAQyjhYtr8a7xLxk9F515CpeEXKWaQEljuL3gE9KpFax6wV2aplwjnHKk4
oUMZhJ6t+WJRmD/r4kfDHaixppUmvcAJM4SYwml8uoPNMmpyGCXpv2az0gxH5pGX
VD8sSn0D3QYY4mMRkQCg5BxIB78+tblgcwDC4kAXR5HNhrDy/q8zTA2y/VR25XTi
J36gyjBQOLU52WyRKOOEwoTmqHG0IJA6/iOMVKdBUsUr0TL5KvZpsAD+nztmFUKF
6xqfdfZfIOlG/DoNJoRqmR7KrwX5d0IsEr95GyF840B/nuPbCtry7IgBSaf+hj8I
FmJIgkuvDcODjIIUTpXeTA0Gvwf39QWGGSfiply0cCjchcEU5ZPjiEbYUJcRcWK+
onkZUYqZrYhU0fpHFcdGtI+azSTnf8D4yuOM7avZ+KI2sHn8aeGmrZk1NXxBq7zG
67DJYjOX//dlDiHA6dBT6kiBcjlL0TyQKfeScMWar3ytqd/OV9UGWFtPzztpblP+
sFyNkfxfXZoHpOjYIaG9dymHQ0rAfO1OBAF+NSbFUpBCLqF6usjexqCX5vjjGT9b
5AxxpzCt2WBabv0dczFEkkhM+IR1aGkT6roqd5xf8xMWnk+l2P80KYiHFyoZM8ex
Yy9LfObpIPECe4CT2W4LMGvsTWBes95OeEzWagARoUouDsBgWKMng/bmAKay8hHS
cVyV5XBjlIc7yz3sM1W+EQ+DHgxC0vlnd/6DrrblVXGKs4AyV/F1izyVjhVBhUTs
CktU+5pE+LnyZIyzLQcp8SlR0nD1DRyS2aeU74DtrX+rtLNqXcjrYt98FtOxV99m
7zWFvAoyvzjNulRj1eYE7tbuFlJumNJDxgg3aHJ2/JRDDVbuQsUEg/jB9rIvAKcm
aRSwplAFjcHwTQ+0UU9hE06cOwHd6FXUVWutAFEYMjFQFv/kVvVqGW6etDef4Sny
enFsGXDWuV6QmqZkdFSXZz2evHzL4VpeeiJKu839HJBV6/3EVdUIyiNgPVKTvN0B
WOQLs0JQ2asp8k64yRlDC0Hr0uGOzZ4Tl45zwf27tV2wudpBLEV9YcgXL+MCfjmx
5Lp9q9HMBRSv+E9zwoiPyO8W1lL2+oVlSas99jFx1QhfJ/5MMCsvniJg6n+KBd7L
whHdm8D9giTawW922n3T41pfwvGEvg71Mv8PcOSFN8p60b5T00e/UbmOL/YEEr8x
g+GD+6OOGZW+ieP02+oIj3og2ROfggKqqwfkBOve2hxpbGjEbbRh7JibozGU6/WV
Ym7wkSSl/ARM5zXgHg9/neEzz41NtGraQq6bA8iC5E/hvHCGc6cvBFFEacbA8U2r
zcJQabPkJsU4XVdtB0zZv/HKLALmcPEMhuB+FvaY0Flsq8otQDe/pS0iUe2wbtts
mSs7f1pRw8BXgk2T4Za99K8BO0dizkTMca5ebmbnHCvrTmi39Y7C9E0zk3v0FHt/
Y9GllPnon1kB+hahOu1iwqWBrl620YCxixBSTIHbtHIR5KUXvl9lu9Sth+Ry/WxH
+jzEwJz6qJI9gKJkb19vMIlkFyaPCi4xKcM82zGiy9Q5ogSjqgxE0UIVCuhf8t0P
3LLyOsQApQtDjP3qocsdVDjf96PCv9aG6kpE586HcDJOKfLehtgcUW7OP5h/iXZ0
7x0ybgpKRCJuadXFcagjdSVSUk5M56rcE32xRkeAiDRxDuaxrv5vfEvD3fN7mEPw
uEj+El5WoSNUvhp33hEsRoo4nkPEVE1VrcuVaQ2KiUpXk0ouRz6dMml70DeWOogy
wKDVEyQ0Muiy43A6lar6gmPO1lwQG3cxskrxFogie8Jpy1lC2n57lrOTpO0fOR3Q
7HOHObw5e58uTtvEfsqA2lORRd1pVAfkaT3lmHWjJ/noi1NSfQpzDzQ0D8G7BY2/
Cmm0zVASFoO90svu0SGd5iVrM4+T01cACBmmfD43m8wMSBICaYR7tdDIEyPMLhO/
+jU1TPtWmU3YjHfTtUpWL7wjqxm/obnLTV6W5OgWZRRAtIDb+QYcqY6CdfJ8WGTt
YSVZTkPuipyM9CVALVcTLW9qrl3sWOiSgZfcu00ey4bW+ArSum0Oz1wGj5TVzJY6
m9MEYG8iyoQTTUqXz7UsOk2agLCUn+OQREio/IndGvj1cn07ZW7dC33OGL27v+rr
Y8+TKd6dXxa8yU66ZZ8Q4B39vMt4fOQw2yhpr+jqXLaZdg4CGe1CPLJQ6qKMZ8HY
VO6965M8i9CpWmMd4XLvZhuY9e6v+uwfWSSp28InVI98YcBnmGg4KiVHpZGgWf8q
BBvJLuMk/xt+a0OMOwi9ssQUS/71hCFE3Pff+mCIfBusH2HtdQAU0DUtSE5qYNRZ
cu19TERBGogpIcw8xvTEO0uJr4qz4aigkz7O4lFjMbM/6/toNmYEXvEPIcKcPqKY
dWyxDjGV6CUR0fUG2oMU3s6eahdkx8SOlMpt7L2aptgNb0M8QZhoZaNkv0diHQxh
qj+5p/6Wd/uBqLI/UfJWU5Cxnkx0Lc4HGIthcSvlHpPINCbDgzEFtHgK63Hlny+2
7K4KiSYNXvvEXV6H0RQMCe4Qob0Zh9/4E9rzj2UMhMQJYsfTpdYUmY0FWQo0aXEF
h05xE3uSwTi02BrmgLNwlceiAa5v95mgpMWhV1L6KyrQYE4gwtOTuplKFENu8wIb
9Ckpvp1PnoEBRkYuBxwGhAm0sPRFl+60kNN337Eq6c9cyFlPaQPR1J63PDzy8qM4
mNdU3g1bVs3LgxjdswG2AUindCmCzfqpBDOa15GGKyIjiiN2Eug339aWNw5SkOKz
G0QXBI2iLKX1jnnKBHD3Hbws6KCjqZyXcgvKAmm11k5VyNf6JOK5dc8TXFo0dsEZ
jxA4Et8wppjHe38cEnG4sIhd0nZWCZVl1O0gr9Zyir4bDr/KwpHW/8s0Bm1VJxvw
Zkiz7GtF1e4F38R6Jj+gogONsiceJfoIyPesTt7OgxVyd+IgdtkDxaMtVA5cxEwk
l4sDnaSz0+y0bIGZCHxv/GfEXcuqs9XGvakMX1WMDNQCfpGZoFUTxfTYlbBWBYMM
T44OVmKfltjqFo3aHZ9xiz1k2Ctlw9YwLjdnN8FA/0ga8Ck7P/ztxwwX9Qz3Mi9A
EoQsXqLxidjWL83+xovnjcADK9ro2JzPmfeLOisMoSkcfrJ0uGU+q4UJYffGCyWk
gYe7/cA8O0nZWs0iwu/ZyR4vGWHRTMScUgNPvV0YUF+lPxxA5ybK2rdCs1twHy91
2pjbxN503lJKSVKSt1dNMdZqg3kaJqPSr6UIU4vNEMIHc7ANQVCTj4qttwQOxYUt
9VhKOfeIde39mx0a4YmRXHwO7Y8pXbKw9f7urpjVN9/rfjAa4s821XV3LgaC4rO7
TrKhOy/LNPCje+U1lSMZJ4gZX0a/mhpA49lhuYE5PgRVPIM4JUhL5ZVGKsgwQq64
DUUCQgV1vNDMJpj73yCIGvRbhA/GY/MbXExdyX4ckri7zWIHzwXaDdOA+VB4HqzG
Edy01enh5/JremjSNiZ+wTNd+Ui17pPQlyO4GM2y9bxtK3YMOraHgk1xtzNaW6Rp
U7Ft5BCYoaLIY+oj3rIhExpBypK29WCdyGqVD7ncin5hsmzacfUEwp9PeSHItOMU
7dAJGkgF1adkyrgsEeL0E7CKKPB780qC66V7V7b9hf9/7Ugq3aUOYy8JSydJlfzE
xJpb1EdpdHhaQG7ycrTNhaBG7ZNTkTzfwqKC6iWkwr1QSx+8ATDTr7Zj2ac6Uhvf
4dzeJ1kYfOpM65cpXxDXptk251uU52ftcihAtPLIUy3Gdn9s3GXWRh2CkqnFrrkn
HSPoNany5CSW4E47lcTWcYW94LFRa2cpHJK8bISVEiLSOQz/yKYflPKEVLmxYsaG
2JotEGcKu7VNi9buyxcQcSQ0ZbQSaJ6/ZSMZhncGUdL2OK0S2+o4CVhgpgrz6aPX
5xLVrzj7jNshy6Enxb6PODOkBlR53w/IvigS6Y4Lgu0cY67yGOFSnDNZwozV+y1I
dl2fyVfnxSYoZszNBFepdrD4rUzWxneiNRKzwGDEsynm0AXMirPhWEHK1uE8LIoC
eeX9+A6vj6MPuf0EnldD31NkJojxJUCvZQE4QDj1w003IFUjEuZG7QCbtsYfJ0AT
45rVkegqas2emmw3KFzvIGnlpBOs0KWWxx6r8Veg1I89957LYQLDx4584kiE8uOL
Grt8ZISwCW3kqydHkOaiuL1ZxKu8vJLZ7bHmdUMj1JL1gLAj0buv7FB6SX1oanU0
kcR2A3fV738oBfQibh3jBMEKvPqD0G9+WAG8uX8b5Qi0M8y2MEMKSRZ8l0GnuOM1
a8/gYf18JZX/cEXcvGkdqOQxt9ONDOHlQ/OkypGaMlGARhN09jS+YR3wuT1sWWtV
GS45xXN+43CgKcxNN5N2PR4poBFdYPYQJQ1NNx/YVZVmdvcCWOenckNVfD35h8of
KSaluG0ZTm38H0RPn7+Bp4KBmzwCFH3bJvjOqkhBjl2nMRheGGML/R9eWZIc1zZU
mZmQZnWLp+1F65BGn83Q482VmolKRURiThUa3LWeVgGIX3epUa1ON73CBvis8Wy8
3WIY7484kFHRjSTu+SK3AwHTcVaLXA6OTzGzyCGPENm2tRucmzXDbEMFhN2KG34K
sksFXyYA1AzahdBE1ys1664RhVcm10uBcEAjVm37qNFf3XzkFBpr+IvFM0KBsSXy
hlAuWesdciDy3gHB7n59sT/uFnOIOlyoUAOGDIJ1yb7TDJlBzoAdqXuLKAiglsPB
r1mgTPj/OBfEdY/ABCVoxubW0Xj8RMBfw3yLE8SDxmoF5oAGDvly7GmjUVX2MM5e
4kGyepbmLhC8ki0exQTmqjmUolBa/v4BmthPLBL5+WJF+Jjfn0iGVmA4BxIQQBuG
vJj1LarlEroDE2F3UVi5LBs5sRsNzl/GCbbC4SnuWp0gZm55qCys7js+E0kftigh
ihv62r8fbPnTXZZxIizWn5R+EoUKGYxHJGGh5vaVZbtNpm00OCrhVhNrr14JyQu1
UDhCFsefVaIPeCvlucFqhtAlA1bQr2IshDNkIQFoqQp9UDCbiGAgndmBrQYt8gox
f8apt6F48ZbmK2cx2i3Rc2GqTR5nVmSTEuV8GZ9IgGKYDMI13F2DnOtxwmqe7lcJ
nBj2IKxgf723NhEDgPcX+78EvX21e6rVqRE3x8siMMzREuDWLAd+Jj14Lu5tpf/U
u67glXw62umSbEnCesXU4luxFuLCTVcmJuEli05753oosqtJUK6Dszb1wncQirC/
H5obdmpJ0Ohhs4bUFYJrsjVlryppRMm/CjRLC/Roa9yfOJ8vxocbyRBd/txwpyOP
zNvkwJesARx55t1heRDtAFaN470K90m22oxlCLzzOH+U93y92aNXCaUeuebodLks
ZR0X288rKKcpzfSk+WXrKR2xa15lJjAgB7mogQp6N8QBTuIlA8BI5iGT6JFtisYh
zGP2Grot/7zyoqlSj9UqFRsBUFNxbX2jeR6cJ7zlQl3oU1nyKNO7iIq9GwUJ59wC
I1ICe2b70XsmGFQzkl7xTT2Kf4hYecRsHw9zhjSwWWj+VA4MExxKPQy0E5BgAz7K
3KlkM/aWB6PMcYB7zRVlIq6AteES8JEWWWafS3zhsXwi2jVO8vmtiTMij5mD7H4X
oXltluhvZsj1yTves7fzZNbNWl0tJFnphWqlpdK3TQi25hz/+mAQNHcLgFpvp4SX
9/TAMN/8vXyo7BZ3NYLm7UbrDW0EhuNbZU2sZuPIPp8S0UO4Tmr+YwlJ9BeWidW4
NEreqS8nxGErtLz8J+P3+Yji+Hi9YRjFnkGRJwEr4p2ImC3KQIsK1X5qOjVoeBnO
2k+70h5Pvfkluaog0XV1jynVFktQYOhXQ4clrMF+R3lqLMrX6UE3rRYSnqLKDqr7
f0E1pnjJV4Nv68Gv6PLx6cptmi52omDwm8A7APxfo6nvUFxOGMmzD/e/rFWp5BnG
Bd1kr24vIvrwmEYySHYkuWzRk4ShGnngBFnKU0HoB5xmABNbwI1Ev7V9eH9+mr26
A81ab5DSvvN2+MKDUHdIHJSyo87lsNkHPbaOvEcuBcTxYVK+GX3KCsIfNAYPkRG5
iyNeug0VC+9VmFPBASO5r1uIEfOqmDgRVlssSzEDhqFsqnAvWnvdsVBsRNgWrODW
LTSHasBEh9GFzp0odZHnAU5gQJxYcXxPYezagd2zXXQKXEBd6+GalIIB0Y6Oi5QY
oZJXjwVpHjzRUi1kyHeV++RFiYFPUsBKuhCfpOUKO149Cz/mDEeeKDek6e/cBbd9
ZEaVEdXxkt68SpEizOeqmERxJoEEaENyjGnyQFKn3MBXn2nl9fWHUL5UFUDRNCOr
xLCa7qcPHrbS2YmmASsE+wr4yHaK+9ZyKZpQJj7/5PqJJnVYMfZPzH6X7DgaRq/k
1S8ByU115JdpSHIHra5otWuwdyILBeGNVwSrDJ0dSV7vaQi1GL5hGkvBdS4IZ7GA
iw4XnpvFEoXXyfFZ78Y0L5txPncqCVcF0guP4nvC/cpxKOvQt94FnsurHoJeWXFM
nwKBYOlH2Wp1CmDpUuqwNYXPNpHRZn6zbgrGeKNNkZFGGoE3lxQzzP3vdSwEFtj0
QTEKQin7NtbVmk5I86OszGAi1lwcUWwYTIHE/Mt0dZ90xgBP/5f6DdmMZXPWm9rU
gIpL+xjdrD+n6GWv8Ybs7yTxwP90d//Aw0leORPmcBWVgZIy+BaVaqfGgUIyQYW3
C3ZtpNwLqQB3dfebDJUM4lOziP/EzT11b5iZLBQOS2XnmXE0bnsVZipbDxBCg4g4
FEtrsBaqUsc9MvHUA+TfgWpy/1+MSCmF6/u/98ehtbeC6mdFs0yNEFeTIH0GroWz
k2ib/H29tHLeqwr2H/uF5sgXusoUunkqnsrl6NVATq3A4hvbVsZYpWhiATTT0Vo3
+To8PajCtJ2++EoKqJ5ZMXiCi3phNjVwyWpjv609qxIcbk++Axd6jotJL4FV6k25
EYi3yiEKt1ihuYPf6JFOvIxhVfPDLVC5kMbj3BRgLTNSoTOP8SsGPR1xpyRSzl7Z
uKcagMOF8LR01jNmSOPTnSDdCXSAvZU6yN1jazu4TdTElR7ril68cv+nW+4ZxT/T
V3EdZTWCx5iiaeiCKX7Tyg8AhKWheUGbjQ7IJfyBr/LWzsIhRRiIzmTldq//q1Js
h35BAtqk86vgsRkGoQimgCnpKmVD4PCdjom/dfmwJ6T7/xPkPnTiirfBioelvVa9
2ScmGtFfN3k4X3R9+auP8Lp+3l6/L/dAFjjGxciCIJp087pcaT5EK/eM1FCX/ijc
2WB4vMansYAY5WbWFK2srkP1zbi0ZlNtPAYldQf7YbZK311xhLv59KTKuHvfIi46
kHOz0gX176BT0LcTh5UzWBG1MSzhS+YYdAv7tFoF4Hw5wQQvTRAlR3dWRamfqnQR
e4dmA2oB/pWk5aAX9FNbJM9P0Jh1nvinaiKOkI5lDUFwrJaCuEWs3OZvOqNDpKEP
w876lB1hcnrFCapIGVzO4cP6k/pDoAkm4hHJuGkSq40UWn7+SQFbb3JOzHud4/Bu
vSCVkRp5u4PjRPsH5J+cyyZA3RcVbowIZj7DNnkXHUDYniME1+xJuD9zMRBtvwBx
8R0k+ftHqJ0XBV9a3t/a+xgh7hrU7k7+flUBwB6Syklje+BOFaBgeZyK1waAmg69
GpUKP7541ZQEWjaDHwEQF9YCr4nG8c/vQ3iW0V0ePl6sEf9/EofU9E+OIOM76cl1
tqtSvkvKe8B9sZ3rSZh3/QefWuR3Xf48HAKO5KhO8LGCWVvBnD/tBCEUqMxlIji0
s+fwQV61nG0dMKLzTdynM5dqtp/+4rRZ1WJWyuNa17qqU3fC4FmG6Y7qyMErK5Jz
kzYaot0+3guG2Gw7GNaBy6xHRIZ9EXC0t7z7FRz/Ynvb58uSr+CUsZ2b23hfuJJY
PG52FF22J6SoEGfggFuGcv4XzaVIj/N6L7kXde8tAnuh55g6wu5VITGOBHtCH2td
ZPj4l8uhHQBLLLOMeGAJpLKEp31OEXj430mMtuP4tYrBACuJRJnr0r0/ZKsemK1P
JXx8kW6+g4SlofLCAGGuU4v/s8byqk3Q91J6IpOZElrv76YtWLeqX/lD8PkxUbyh
f5waM7JTfc7ls7r6MxWa5bJPP9rlW3Xy63coMju8JY11TIq5TCuQNVrc165iEOcF
BHGL2y6BJ+wnvGxgzfp7nnMC40qpb0Nv8PCevO59wSJ3eHYMie59Gdi06GvMApeD
tkSn3UaGvL1SFyz/08WfGlMpaNKveoweoyCuO84wTvxisOZkMlPSYxxJKi6I7OM0
sDV4GXrYAMv19MxrMpS18TYdPT2dVbGwkITB51k9DMBcg3MIJJLSHYIOpocpkhED
SLh4INUG8bl5qOwYg34E3lduiLsmOwe5KvlE60qyALAliFnQg782EUsgrS6pgyzP
IfLdiD49WpRLOgPAdpoapaFeBI5XLGv0LIa9LrOsaN8U8mmQ4qvhuIz5iNqOAPwi
GW3pnBmpo/O+jtVgyUTBDz9MyjmJxqRv3ZaaJiVoWmX40cDZUsH3aV6RAtCVXZF0
oaB9a1qxAClCIPopz94hL5jg0zNdgsGjuivD8LqUtQ9ZZ8geFgY6Y2S42YLmlYd/
YJd83NDGsmGelWBQdEx0iv59xYiwH0anDbDnjnX5xuK3QijhKBF0TL08pqs3UgHQ
+rIuNX6RMwXHYQMLQKnoQQV6TNrUS9pHhqX3Ylkco/ev75K2GHa3iOjplHhd1Zxn
gqKhyzr6ki9uUxd6Wl89Lr5NJT9v3M8kAi+fES1jHRjk2iO+c+43+9TcSrzutd8o
ynrI9rhfE03gdz2RgZwWWvILn2k61wbpei0CJ0921Y5gSNJt0FxNNLqQ5Hdu6p44
l9SX7qmX8ifiAWp7bT2T37X9gpEVnQb0qZ5YSNZf/qWhEhPlRiabMYs4uLnnorss
bJt2/2gePvEYojbkw5YX2Zwd9EdE2hvL8pTwOKosJxgftTo3QUVu9YRg77pqq+Rz
LWIb8ImDOvTYiGET3mQ4Hplb6zhuZh0Ho2Va/PV4qHMGgZRKkVQMqvCBCX+qbT5b
7Ec+tyGWkoljQxS865MdPT06roCd2GzzLHW/cvQ4ZGlbYIO3axPjH+g2w9/6iqEM
SbHGOSbszRpjVxJ2wVUPwWvwTgTVnR9cUc9XB03KascpofVehiTDLM/nNBjXRPNd
FdTZ1iXUX8cZxMg3svbByLbCOd7m18iuZqwF9/j5RtQXMCl9UtlV+d4UXoalWZj6
waN5JwSS5n3MqKkPcUaCF1qXuENp7d8XMEerXUlo4prlP7EcOR9ign75Q5g9Oj8n
z0ytFTlvrqIk0t3rft8lXz9KkdVVG8Cm1Jl5xQhNpP+N8QXUIWkJG4Y1Zf/dlQuJ
/kEo12wCndegK53R4HIeIN6PC05Jptjk9EENmBq4yxItHWFTWZqM5yS8p0aL6wq5
Uecbkn1Jfi39TJmDZSHzMEsAILL9GTSu3UNs+wuBVtLruU9EamKslc2aRoqRz7FT
mhmaZcIhYe+q1GPkzecQcpixRviNbXgIA6MNXPHMNBvsOJ21slt6PMBEjwkwtS29
ml3u51ogsZsh9cfluuMPVy9Q/8EkhNh746Cb4PBlhgoDYi+1FsdLRoLOXYwvVpYU
YbCpUmQGZXbAl+Haha5nq6e2DJWnnLkaKqLvbAMaBLb2VawihfQsL9ITln9ymeb8
0xI8ITzjgfl9y+qePNzFbDACUHEW+rA1wbVL41Psti2/TvJAyXw7tnLhJgxBSVY5
18Z0GnLf09RICjaB+zsRKiSfxCZeIQwz/u8MhglVapuwscAKSOXbKY8vyp/7eoJr
clWTPuFdxJsYl+NIz283AotbFqyDaEpEpVD9UgqPm0DghiO4R6zgpP7LmKnu4EaW
Xufo3jwtCf+SEOWoQA9QJ5ikFfddfPHUTb537jIDbN3id87Acg8C5db9d7r5kkeY
MCZ6BQOpoR41FrAmnA0KBKrQ1YJXT5TqubO92zAXcYJsb9IWmpYFOdAZI8SdCBPO
J4hrsER5Y9T1YPi8Tb4z+CIqoYeAYXonIWNLNKYvxgM6e8IqOBJfxKvmKgXvCMHv
NogmAuUe4mq1SZDtNpWVCxXqOILGZrKddJBA+7UWP3/yuiH7iqrN/NRjpy/a9ckK
CaVUjGX6L/549Q0Jbt2PPZlc2SuEZCR6/tXckm472lOVlTYJ3OLsiljo8TeEbByt
ZFLQyWefhhH2P8jm30nY/MdBSO1QM5aNFA/OzmlQg6blFsF60GAVyqO7bH2dA8GK
1w/flG/7Gnrzy4GXiwfTM7Invh7YDvpWKp/TNp5gtQO8CtCxysGFph5aaLAnubyv
M2pYfVGfampfJEcAKuM9XR92wvsuX/YseOezDG1gdQo4+lrCig/VHfVn4JUWqWq9
edk/3WdwlBRryyeY7I165y+ikIeHIczUtAzg+/8dq06F3ldryfASIetd8y1kBLS0
07undeiQr+Hy3QVdipZCnz9nWopNhaL9OSVuXnak123EL/L5rm4zymfIArBjGg9M
BzWWbUlEzjWUohUTI5IDqVAlHhm/iAm7Lyt1kIlxa9hMHVVpBo1nlg//WopWtajI
Y8c0MtnB1eBeEEgIg19f+LcrLm+GLugP5+uMowKziEV2vUHMGoT7vQOZAnfCReRv
pcxHos0+6B4iCukoNDdEIoWPuk6P5axH03QduEbaNhw0D/pvDnf5I5FzvpFsgnVp
Xgj3HEVB4jIGhW4eYU2kFs51laezYu0pyg/f/QOTLJWzd6SbUn4tOcAb81+pEbYp
ICNMnHsJg8pojmiy2th/x51FHwLbkx0JnGD2yKk8Ig4+xQ407cIwaXYqjBJqIsjU
nbHm+OC5/Azisv4eDPBSwFgMfKFZigWIaI/1beJEQvbkju1/frwdavGOmgHVJlCe
aHLl9cbSOQWM0H+Dy0VsMLaCcMDmd/vbWBE8sA3zLs9pFMoe1JCgV0vgbACgJXhB
UwmGrWP9SilNEzzC8sOj7NlzVW42Q59r7OLBS/0Kw/YuBrd/6GGOyZyQG1YgVQe1
MfrlSYM+Eu9XBNkUGt9OjyXbAnqO/WlJZohl4bDM/n/N1EhLMk4U0vvflM7q6fF7
5A+gyUpFKqxpDzs9T0HvxW3C9qFKljgjsZWINFXQWMhVDcRWGIhe1o6XCpzjWPhm
07Lme9QMb7kJGkO8u2mzQFAau4oOU1eeOBdb6N/ooKbjFrhvHLif/0S6M7b8U2ss
hh3/jAFVB3K1wOC7zFlcaqYI4cDiqTPDm7C7jeAFb4oExz577nGN3D5THZIlK5Sk
u1xiGrI59NcAFHdvti1LEWhA6+0XmIToswpRN8/4NPkiq3rAvYKVHwMcVG+xt930
CCC317+h92AMypOiYiUuopUeQvDUt6z7OBR0+ePy78e2dpoQ7WBNF4boCQsa3Ic+
+A7EIh+BPQ2HcoISy5XgkQ9jVezTQ97Ns1OHG1DQ/miIJbH9j1KiITjqiNh71dYO
4qOGDw2MCS0pvwHT4giWixhpLplZ40EJCPLsEV4tmvpb9q9EMrcCAVjw929/7pNS
KTNWbFimXgMqbXOsc8nDobuTc6sWMLMYgG4mDBNQFw7k0Cm+3dZthkIkdQegcf9o
qG4vhEHQhCKJVObwPl41nQ3IaCrCETtuFt8x7KS4tQ+TnSrBt0/w1pXZAh0UyZjX
UUPv6k0y2ZE4cQBuAq8ySU6oFvvQLzjEgTdsw9AznxEuC+tdYTBaZeG0+1MzabrD
osdKDE9ZA35ouLRfZrUs2PY7g2MkEvsgKktI7z9dSy8Brd7kZHPTLr7m/RmRiXrK
JewNaOflairVz+Xl+AGs/rEtV4zkFjyHtwaa5fAPqrTbA+p2+0wWA5lX1IBD+Nt/
PF/g+0uMN8NNr0+pBc+b8mJw0AU5Eze1sR73ZT98puiReBLXNHnDMxf8vZ/IrpR4
zF0Cf3joVNmu8eMCxh3rbXENeqWK7ZU2HKGmHEFi/x3oAIQGH7W6xTNUw7EnQBe8
tDvQXjeXeWHKkd7GthoFKPd1IAwjh6YwO0UdIt+iUy1UyIS8CbkuOzDN61oDK9W0
tax1oRVzRnQzB8wYGk0Y0lqYOCGyD2dV5OGflQxOlXuvP3QCxMFxBgeOkMcAAa4p
JJVC2BJb/ZLKvo2aRfg/f3HnAUVbI5BYcjDex9zrfs/YdyCHv00EGRv7/TeagOrE
O7muXA62zRIA0GjjvESh7+gzvZUUnE8/585CoGlxLeK1vTUoBEbA1VPDWfWKMSOd
gYfeh3yT/WdAZ4XNmfcJAN9o6XaL/dKRQ7POkfc9lKfaedJh+WnOVs3EqZBucHfL
yci8PpBvfOXvXd8QP42gtloFmQsIMf6BZFAz8VGTIRZh2FbZWRttCpsr38whuuLi
b009xPYoJBnUdG87FQ0/Q75WW9sUz+7GCO2nXKBTJSZXmMnvE+Eo4nG/hvrCJwAF
mc2aCEbgO9nvIgY6mv67Zd0p6JeA6syafh0Cazn6z9jRFm9qjggjkBJaCyyEwQft
m/v6gCAt4A9m66OZBhhiuucaNddSSvohH0ICQcHi4zFHP9ybDM3Ansor5aCO4QUx
ETRMnB9W8TCXuz3FKtudfQ8xE5sfo4Yd9CsNan3TYiMSYRfDYbzzt/AkwDcK+xFV
Lr0PpVuUzOArmbM/tlgb3BAHh3HrKFLzxNV6wnOSiaBVw0q3ZT9QkVY4Ipiylt+O
udNN8Jmo2RVA2Ul5HVJd5O7OSmdf/gd8pOGudWFJI5tUFuss6VJH8/ktA2VrwQHv
89oBX7UVl4eI2y0R1wxXUW7aH/sV9TmmZb5XBKch6bIi5PZbQZIizgm5jZEd8pYa
/6cZbpG5lD19SjP1U+Yteukihque/mQHCBf6+WBnmN7nDts0lBlUw+qLesp+XOKE
ZEsr90e+q5Z5S9pd62perth7mbFUoXlPbwABRmY3VIg3hiWSN+k5Z+rif1GmFd6W
XqpxbRDlvlz3OHz6osXQlk8YA4Bo+ZfWdxf7Z97CaF+dQb+q3WkAGtndQ+hoXobZ
dreqUwBarbGsWV4W6FIf4/UG/M2/wpZSnGxldn/VmwMrYZEYiKj1Qwnt9sioxvGK
cwBtZHj0Sw/s7jbDOgni4a41eU1e6hIT5WRuqlM2wOfvAAMxhau5Gb/BcleisU4p
eu2yjlvPMfPpegBzlJGLOGMbvNVBfpoTYCEEINCtkLAdvRkMw/I7vy4IDi0pSKFF
4VVqNNGnMbXWRpTiba1yEEb7f0+ijhaA7adT1eI2e9z+3YxFhyRU0bWlzjtrbRSN
ct38M4HsnyGbc6qVMl+x+5Gb4JAaHr/ugsh6MdGmicCcLjVXvUMB9ocjVim8Cwu2
b8mb/TOf1dksOUNaWTvfUn+QYW9vcAwnYyHf9PJvM8YwXxIktXGjwNLdNbGShvj0
BVN3AkfqvnSrDuu0P3k17TxAHyTHoChwNsXUGJ0XxWARe74gKGXY0p3rSUFrSQLR
wmTU+I+M6WuSYxcfbXMaN4ALOQhrcOnYdDcgp+/OUUJ0DCtIWftzZbCv3riO+dUF
YmemLHL9+qUkLwrjgzL7pBk8NvalrRv9P8E0FAOoDP1PjEvg211DDyoMLyaHGQWh
Txi0Tm8k8unEcSo4lH8JIKAYJNbX4g2dWBvNoRqwnwe1D8XiflE2gjPtulxs9Zv0
6S83yBERNUHQHbu0HpRfPA5KN/Yg1w0QjbEsIZtfhsP3Itc88qiy1kFtUwz0PHS0
x+kmT5//sFt/vV9Ic+fjW3eAt3IcIua0dy4GN0LTfPSim9yc4q+cTqlU9wHpCDJF
9wtOq72rqUi7kjHAAcX5IaIdjVNdRq8WBL2dgcQd/qO6iOw1tXxKPgMyXrEn6LO7
f4lLKSo/RcbivGSaSpCIFNjQ6LHUX/yuR5W0IKz1KybDacC7DOxfIAB6FoTl6bmT
hCAwV40XmjKTD4N5p4wecC7zKtxBSrsd3oMxdrMz5Tp4AEp09SubsHxPAEOdqwYs
LFpPKOXYQWnLasS4ntRYaOcHGLlJyfmNYQG2IuMCuvG09i3iYqR4su26Jepya3sG
P5rB0+Zzk/sKavz30IRnT1pXzyH0kPUgkJjdBKjfzRuxnwDhmE9i9tSx0Rh3j2hs
j5oThYJV4QU77Wru8B4KMK7bO0HibP0QXhCG2pr58suCYM4ID6dGbrdqPoGzh2j6
dfDxdsgi6CkvTR2mxPbL3C+lRkDLZBRuZkDhIm4Dpn6b3fgwjy4qlBetcbBes8A2
QwL/ODtJ1gZuYJO5Nmu0o4IEWK+jR59J9ZnWi74BlBceYxzTq2GZ1L3W9DKtzzwo
5g8tn4j5SuEQ3kBsYH2q2BmOJXVcgIgVqyDm6o+khxZPOOA0iTjqQ20VlJrwFrt1
S1olWKERQLK6E4OYOTM5t0C+jwTm+jo9R2sYK+QN0Ha7VSg2j0nr4cguPIhmu78+
EJZwHa5/vUDVwGkehV6sDhgXg0B/PcciGzfkhFLPW3FRiWj3yHO7L8EsZ9bmf6nT
dBIMGIcd7ZISR8QRwLp6E7/7pMMOG6Jr9ksfBySNKv3jJhVMYSM4p3p7oQP3rpPj
UVjbe7Wld6CsX6pSfrA74ALhDidHsK0fh3txczQoDWJaKctghZiCcwLdsdl4nTRI
PROKACifNn2ikHSxtkXPFf3cPx+MYAm4XlyMV7kgoFH3QEOglskFpX1/Kdoi8KB0
2MK+BRuFjJeV/veBX43ThU0FjxLHi6j7D5/S5LDs9JXshN7zTJYcMBYTl4yZFu+T
E5dp+v61tPoOEBizWAvf2kMRWzXN/HeDcAwv1rfuY6+ANnHN1ybpEwR0mwvS6nMX
8yC7rhijsV/VwgXjTGL+Iww3Et9qGDGtClaGVE0/CSbDcoxRgWQ0/xTkdf5BgRLb
ZTwkkj9A7rhTnhqR4cRKMd5+IJbChXROzptI9OlmcInfFQF4nY5/yW4Xm2dKOBiX
7ctYmhXe8Aop0pYNZ075eQGYWe4dOOwNJOEIzVFEprpHHj6/waOHFH7wGKEYX1iN
dN3Bj5Qwpb979saNxNxaXZePbLWkqYLEP5J7qHmte2KjxNjkU0Lxg21oeKBFlTEs
cp6W/GhLi4J5g3poBHP4DTKFKebaaqfYRm0Y+6zi8rfGJfUNBuehZLKDUIKN+1Iu
dupYWPPXLPw0RISu4oi5I040At5aqD8JpUNMDa4CtprWNB/9iZ5tkTaq/8LBxdSb
MG3k9+QjvAd6RmGXoAjoiOvm5FFYmkySF6nQyAbqcNeSzl7REMEIECGLkyOeBzmg
c3ycw7Xse9UpjRcAW2H8CmUDo5rwjYobh3NwTwUaP2+wHiunI0Rxfs7egIKcM0CV
l7iQSXYARlvwXPevvPuSKslPh8RJ4TyA9vXEFYgomIetl2mOaxP6xB/QrKmojjD2
3iF/2faMvdcwhoqgg2az+1bqJiPXk+VogOqtJUHIz3wVX0k8jqjikeBrBKXGSo0H
Qmr1SELQcLLP+chR6lI2ZobpV6wjnQegDV4CRh+IjFp/ckhoSosm0W6lyjcWFwFP
+uItbAncaL9F2sZoWWmQlFKYFZ89sXDfssJJ8MlTcsZ9/YCORB8JwgiVf7Kihz37
SsH5UhaFvW8TueJt6kYsCKVwY6AoEd6B5fgl4tJ4c6hoo2/BuvBVZ0NgJFOMlNX0
TLK957dgAUEroryqv4Qk1t1dg8APhom+UufNNRPlyoZVoJ3l0wqG63xVSXmbPseg
K+6QrcTATINM2+1gaDd5M7ZGaj0QYnM8Nwp/WBH4BhaK0XVBx9B9Sz7ISvlcvBmm
3DZbJVqDDVbp/6jHUNwy+hWQcUfi3SyO4bz2ETr2NMwkILHpfSHsF0ILy3xZ5pof
u3MVL3qKuBumZU/B4pc7FJuUJtCLWCPYAHI8de79+o317oTOaMhLFntSKkU4aCAI
CD2o1aGi2eiwmU5RdDU1CN1dzZIAIqR4PbP5ATQSgUZfI9j2tl7C1g1bo2XWdh1C
Ot65Kb4XpRphdoZko+LKUu3QZgQfcRaUJVA+w6/JEfuqeUdbxv8XyWoqwroZ/UK8
unTprvT9QL31f7wNaWUcDvXBI6gs8AdFg47FRZEwGNZjb22VnvcBSaHwdh6Kv/ih
LZMm9AA5EzrJtkexKC1evuGhd5l+4hHfGGZFeBI/ggRWM6oeOqOzLHcZpewEjYGB
85VUkSFAlzlRUK+L9ojQNT+RxkIIe7VVkO2gCSV+BQzrzzERIw9aWPX4Ema6GMvZ
5oT5w0wXSLtZ9NNM32LbG7aHj2Q1QMSq1TEd4dSOVjiZrtxi5pFJHtVYwtBsZ9aL
2dVWojc8lMsMrHf1a8xqiqlrTu0ag1mq8lA3r6Hcbt1IDB81LQw8t0wDdSAtVpoq
hwcOUtXdNPrnNfSnNHZUYuC2dQy0gPMLIcNNzH7DZ1RcurlZrm/+ahC1zcK4nlAb
8bazSoFZn4qgIuEPuzJ2tTjFGvbq2+tpIS2OSdBB8W+gcnBhSYFFgNZ+ZvLd3l4+
w5e8eOfsce7W8INc29QTJVz1OW03ZwAt8R8gzU9+TXfTP0oQMpNSqZpIK2LGLHTT
iBH2G/Pu6+5w8H2OuuA6vx6dRYCXCcl584CH0XOuxNPCkB024EwwAPU2DzeMLiJV
9Xy+pYEMeyER9klv1b26zd1cqQ49pmDKFSG9XT8+94IudunhFiuy9MEQZBDfvh0P
pWMtwJjk+KQaMGJg8sLddCXRIKexca+94bDRocKLJliqW0y1jTNTvs8amGqhw0g1
n92jgmqBk1yWrnQ7tnnMOKfXF4u1vyU0zvOjaUsJcEidSLP37a6MaTKw3wStk4xQ
EvXeO4FwHzarYFU/RSQrNK4EH9ANgfotJB1KcRFp6uPk2p2VsSOXr4jP1gQa5Qbx
I7LxNiwze2M7yGoqeL66oHluuHdIxw7kMzGWBeqbDt1GSztiXC6vZva2pI/irpbh
2P1n+HjSTSinv46NR/U6sEh30WSyicdDtVbXVOl3nycntOy/krScfxdt+xTXABum
+zouUU/pgj2tYXF9+WCa7fU+uOm3PpN61fDffJrnWwxnXlwyrO7cN8xTN3GqE+m6
WvEAzlamClHBwKaD5nycV85qUjaf/PIlo7QdcmuLjVItgMonmXMXPLIfYRJzOsIb
AX7NXLSjL6O5lzcJGo03600GHYoaVUK8sj4wVBCwc1CbhhGz8q89gwmYDOmXQv94
LxeZ1BSbqZGa8/KBSNn9/hIpeCvCKToWG8+FMAOK1hF38FeC4VGvMsei63JuJ2Of
cxEUJCR5CId4GLX2SW1YjKe1ztTY5pzWhoTTi8zdsxUfmX56kGF1mmzLM3MPycQ7
mAKG9jvms7r3VGOhuGBWLbWrfkjvz+DLhX9fP5gsZpEIhqCEE6r0A6W2whvtz2VB
OaVI9xe2iIFmaSeFghusG+1WxxvMVFOOM9NDIIECwCcYBX+8F1Ca5U+vmKHNKcuE
MNSdgVNEHw6Bps062bEAkkf/7548x2ueDfFL3cLHWh/CHKwmOeUewqoWQ2qY84N0
BI6un8ms/+fGLhXHAlZxZa0OYR/g4Uog82rt85JTR/RyHZvoHkxypQnxleCPrLEf
appkONCxpEBeWQS0cDWQF2F40wfK49evKouoaxyGa0j11lQ2a7hD3dEUPWHUycu9
As9DClhJ2x1NA8lHTWbDteluRU6chndLPfqk68NAjAKM9QV0G45ZciOwsHnm+JXH
pT92cZIUCsbmQ77M4cxiQhgPV25FzjNNgCloIBbFW7QoiTHUCqiyKUucksJ5GACP
lobQAYJX1Ujifk99l523YO5C2GDZOHwdiqG+4MTpJsW231DFXOZGuCEnKUhS2YRM
mVFPUdtInFHOvPQE6raWdiN3L3w/YWQw+W6rP6PvDkAuXbRbcGMcfCOMZJogpaVZ
bxAX/xIc31MbO0u4kSyDFRbNGRm7BTFJoEZz/6t7nBpkq5kDhGXxj3ujLC4+bKuv
UxCf5A/PVSjQchFjMO8uzord94ScJWUYfMjNSe4cuqLg4sLNEZyXNKQN11TKBi4U
0LMDee1qZGW/ar59qQ+6IxrMPgxLBips8IdeRYgVUo1EB1bwLuL9eN/3Jn2xyHWi
Lwlb2ZR9uPC4eKj/cG+ZeL2RL2uu85kUeU7ZoadzgLqE4oGAKtoZn0Xu3Uiir92o
uIzl+MfFDsC776BullP//w/2xGLZwifuIb79j5l7nj0WyhLaccjIFjZmn+5H/8Ew
/s2Cywrmx1hY1okPsX6conufybItZj+Ed/GGS5mA1L4NGwm0ngBAq3N+KXwUnHoq
KAr8zEPddvQUVSaoKdDfYCX38BI4cT/MFiWt30KuUjEiVDaBw4vLuifZq2E8HPeq
332jnPZ1eWzGNOGzje6eXoXFaV7MOUrm+0qYPtmwsAnS1Qzng92HBMMUxc7FMoHw
j4mCXI6XAAkQmivBbsCVDrv8XaMQCa1Mi4h5vWKsCD9DFuYXKSsD+U7B+QFVqCjo
dQCcpHlYorjIqwJ7Y2MfWkMKoOZrXleXZZ5HbaR17yYiAh50hKNdHi5kDgovdCmA
/S76jjkdUcm5W9ek3cujWR+Wz6YgxulWVEErTM14GC3zSgTOD7+jJXf5tugncRWZ
Su2A2cuzn0Xe+EDkNGi7WK37Qp/PF/iB63ckmMP0IRk2wVntpMX54/m2vnlWzkYW
7NFIhtAx4n2J1Gb6tVQ7hpOPUuKHltA2rz5LTWqoQ8gMAwvIEQYcw+ftEhkGjoZ+
XzDL27V94HuJxHWkRe0Wgki4vYl3WsefLo1r6V7tOwKR2iYlGNOAXZofnIYZWRBv
2gyTgIJNZQQwL0S3+5oEGxSyp37dZza64qEjslBr0Ic71vrxLF4dUI+gic2aplMa
vcnjheGQvNvDQ8aE5Yer9YThTGOfPdMVMiYep69mdX9kh19mjJO3OzXv8MqCdo+6
oPxJsY7Tfc2Egkh42rO/THHMw6Y5iYWobHaYmwFv+PGZ8AtQvB2NrFO1DxyaMst+
x9jolz6ZHNEdwcGkOPJVrKCob/nzWtBI9mYwUeKqrnHc4pUJD9DUVi3D9ok1Rpsl
JHf/WqTVNwjzq57vJxDBIiaFCgVciuktx94Un+iXCzBXCQ1jqhHW8WXL0fnIxsL5
fTzl40ZGDt/i3iczFk2e68uDne26QnyMMpRyjq22M+eaTNkVW6mZKyXo+PQ48bLB
EmE/asQEnGPqhw639CMxNZBb0EvwK0IUDuUcanCBg3yNOcAO8FFBU9aWq8g80BN8
8kI7HjscV7EGBwYwMSuSGNY6Uu07reo3XX04zXz6G2MAh0sFncVRak1cs2x/cIe8
CdrUFrtRkeowpFcs0ynDumTpr9K1o8VlKLEKttHcJdg8+9ahmgDckQs9wTBP8CSc
DW77pJH9oMWAN+Ny/IgVdRCrITi0lxBjd1B+6BA8J9cUkw9sm99GzHjGGG5ZmEBn
/4x6TY+8HZZTpEPgKtJt4ezrzIbRyTCimXaqgBEPDRBE6hGwkQL/QOgaDFn3J/yA
QERyiOfGzs/PR+z55KFg53pqpKQ/xE7VWswP1wYnryXYff0IhMEIWBGqeNWKJUUz
FnshzRncYfDpvigChJn5bp8MESItXV1WeQ+0NQGtQjr6grgOt5KNviLfecHDT8Jo
TaylanfWlZVERoFAOXQp+6ZpODEZBjzxJx4O9Qr6/EiE592d0P57Yq0kzU8ynWqX
fEdI6HrdUV9RR9jR8d+vJJuZfBCkwghaYV717imSjyFRHcrMR7awWIiPZIdPmoVj
sbH4saZCddIssW+ifpn3SYxr7mp1vjEjNpmLt1ubWulB5X77YkM/AjUDfiMAdjne
X+98ix7LtLoYywxTQzQWA92DIXEtqbMRbjq7w7iAsX01EH+fpVHG/UBAt1tsIhQ/
fYv0o4ikcXlos+S3EjtlCile7aXqvSiiB23oHkODrZ5JBZyHgmn1R3kc+HAe1Ylq
t0+XmsU3a41noe8GyTwm63lV6gfcnJKftzLR72ZHUeCIFDWolq2u33s+I0YWSTyu
zjqrn285d3NBO8+BR8fX6EyCiwX3NbV93NPD04e4SKpJKtPqGPFXDrSufpb9wyyJ
c2Boun7lc5yeRU+4cfGSGhUAS+5iEbVYJEsaY2Zp5ULaersroLpqa/jVFTkl3w1h
UPxf6K6b/1vjHWDxb2ugb9xmlM5OvpWGOTvPTH6PY8n7ya2+4Mgc7YVhQLLtUAML
xWtQo0ss49oEt/CpaT7LUKytyz1Buh6ZBFIHhZSP6kU7LqCSDcZI/3xXPKfcy9Rd
zwGLuHil5GgGVcgJAsfg3Ine+h+zRmy9y2GHDvggfQ3mQn9nsWBdQbSs0gSsoi5J
RpNZp6/fUmjHE5QcrJ7wOrQsAOtodbrRkRn+XnzDkm9zVaNNCHGl36HiYb6NwCht
/NHEC2TEu87GQJvg60Bw0JifAmkChoD7jAcC305votYl4tZy/ICejwg6/qYun+zS
XZM0kcTeUPta8L1u1cdpYH9YLuEQfSRusIEZpBXeJkh4FYN9klqGpjY7l6CbAAig
JvuxNVtOyoR05XZ6LgzLjK/KtWs3dIxa5rGnNG1/qcFMSWqYw2LNx8uUgXOJ/yYR
JnSTr73pFY/6Ks8NU9sYz7N210rx/hcVh75q+YyFmetVT2dM2jvqpR5yaz/g5HwC
doKHxjvz9ufudzPfD3tHPMO4LJeOxIraov+bA7ymFsScMd2pDmlIF2HC8yFZN/wY
8BWJzkFzVZZu3Dst1f+SU4fJswTDO81vEn0kqqfBFPl5ZhcH8XnP8tN557tb7Y28
IZJY19gytFHxscdGmjQyu6hRKwmsvsk3m1kUs6LLQUyirNIJNz06H6YOuKe3I31G
VIFG7IPMiiM8VPtQr+wxB7zr+60C89yyZxkv4f0Cn3EJFTMpLIwmb2MJEjN3aS18
iKCbsCAoBUK5V786Pr6jFBW2x3EIPd0k1YN7d07lq8mdhs9ZKpbfvpj816T+1TsW
BQOo0mt1wkqbohs5xqd9iYuyWhkz4fd3HU4joL+vN8r5Vziea0TJG9mp4bX+6dn0
MdyfBnLlctqxhsximgxtUkjjd4Gg6woYOY8+wkwYJxXYkDsBAvnxYsregyLrtadG
rdvgAmD7h8I+LE+JjuP5DBa0/NOuyXMTSYUMcz/QScgJbJJteRFcLU1ljzOkb8O4
hmwLOxb97JYOSetKq/zKExB3JX6yfegz9fjZHv+ZazEEvzVryPixIrvWtBOUJ1Sv
tZ7pklidJ+brfpXqLsvH63XpwZtFPn3rn8qseSII+A183kW8Lm/IN58aPVxiS15c
RTunnYldGLUNCQwfImvTYZQYS1i7spIAEB6+V9fLpaGM8ibWX8SZ2LaEW1oY10qI
Vp0Mg2rXnuQdaLr7v59fVQWbX2XT0jPGoD8P0niJz1ZiGIAYsKYHDHaqb1Lsq0wT
wSKER+40iF39trngEDi+2e0M1jMxLIIM7GxBYivkgin29ToLn3cEDUUZ/Dt5FhQs
C7Ye5Yjn0RFXKSajT5E3rvSj9et1ZUb6cSeuW5i7ZBYROXnJTmpGHpRy6ksLubHK
Hr1XXAYel6JBl0YHKXoxCF9cLA5OXcl3ts0z5ShUIcAWx0VUd30XhCV+CTv3p6mH
mQ47ANW/DcpO0mVcE4zwjza3Y/moZJtD3VoMsm2b3Aq1Hc2wzqzvxz6FlaFjmXIY
Rq/v0Hc4nmAjZLgYM/rnxbp4wGifg/ha9jGS11ndJoAuKs+iLpZbMlYOKw1M8vrL
Bm7aupUO+pTYlCa4ZRQXjh7x/Aq31C9y+8KtgV9USrjdX3T9waKb+D2vqjbya4Rd
Yoxdm4mbzg7Gv3h6LxekzKVxLJSTfd6C7/mvf7h/rKNf+N8YfL+vbVLQYDYF1jSe
Bt6ENMbtQsk87+wnnOUoyqqGnlU9SB3FrNh+VpoPuLAH61Zsutr2ThEmnJLelZ8J
x+I0wYwfYZr0kpWtdxKcZqL9I31SZWIT4qgFtDwXrLZ3SfNiS6E5d+GX1myvot9j
2iIfTGU2QW7jVNRFlrGaPjLT0quK+6deYLSfG39E+iIZWKnA2UJtNUQqTOTo3ena
5iJoSWmGw6PEXwaC1rA6s0pzGEG2EXjnSti80U+Rr58A/cij6zA9UvYsFkWGSf2M
DJxRjzdAHWdW5AtyrjHaU6xC8DWKErjUwZkvNlTwVAjsvAwThNxbqDrFYHG5wkf/
onuY5shVxoHYdRtYr/mfsO+4LgsbAg9f2Uu1A92WdWS8Z0VwcRiRl16Ip+JbUgWU
i/F2gEr0LR2WZ4ElrYgEOqImEKFRe2lJY/3qiJ+n1CKFooBT0UzBJ2MDyDjsmnpZ
jD7sTDz4g+2czW3BCXhlU2Hk8E0/y17QN0TCKJ9PjuGwcLMFuPskUIWY7BSCeFFP
i+Z0H0MPW9Ww2NYaMMDEeb9rldUnFXhCqvlQ+QYFPZuOC4so1gs6tTCCm3RG4cCu
rxiGDDUXz+iiE22Yt7TnyRJd0OLg1ShjlqhMTycAYmxP4DmTdZXSFEFZkHLvzHik
VBvw7Y2FsLwGXy7J6TAqOb+ttN7StxKD/t4gQJ9++mUCt44Ekl3tjcQmoWZe31Xi
AS6Ye1W5qkSGkDGzuZawkpAzY7H2gh8orDJ1rI3+ZCc14B59K5A/QLhQkkf+HuN6
/z7/raT7BHbs8r8GOyH4pHmIdsdiTLiYJwad6QZ6ZpdCjKyG4HY1mLrsSYvBWmhh
vs6w0oNQwIOD2lxXoxO38b1njr7bkfR3MmzfxHWq/g49i4tJjgaOYpGBAl1bxCvX
XJErXQZeSnMWcR1GH05UDgDBGHQI4Uxutc59Hk1mqbrMXK7bXmVhsglyvhK9vuC8
bGplvKD8+kUBu2Z69+7C/w1F8HchjKlinu6/UNNxSFJE7LHTu5yPU/3ybDsQRkRy
YclW8mCdFKZbpnxMacTxqw2fkJYYJbV/qY1n6akOQrEBu+GwGOGkD2fxbXZlaawY
mrW1XBiXaU8lB5zYAJ4rNN2aUTkpaDaYwFiYRxD46CahsRB2V9wvO0tVRcVXtyeM
V0EPSUCqA9zIf6ECi3II/h7T5A+Y8qcvBF/yDWuCFAGiqgfJUc6jtlwrI4VlBBRF
UhUanrGBfnY2vPEp0UuBGPE/DZyAW/V9iGpUEDIrFWtTx86fdyNY35H1aAxHrHQo
Y3d/0pIH2eZIGURcjkf7tP0wPLhYRadS5ycB2JDB9yiVKvl79bqrbSaE3Ry6pflD
2h7OZf4NLUT7c8PXzuUK/N7hAUkbsHP4+7DmszWq5YotBHx2ReI4YVfPIgFG5H6b
pqe08jAXMUAtEt9X74eumFLdmRgs5Jm5WH/gK312mKu2yNV3qnQ6sR8cjd8exDHN
SsmgH1hWY00u1BjDWG82xRGjyh+adxZ8CTVy6lFPmY/Q16OyjoN9ZKiWaEAi3anO
w2aFo20rkMWAoRyNFBRzZ0K567wmDmNYpeH6D9RQSOlqFRm5K7gN24laCe5lLjEj
iKfOD2n+MUPFptXMYWQEY78Z0WjPKvGE+nG2ziEtJ/mBOqLCeKZh/jtIdMIC9H/w
NpuTN+34YbpJ3uQvuxh+J02VhxevIFC6RWMjeJuPeiz8PjqmealJtRml9s+Rtgd1
YPbIBR4I+Q4BqPNBW8XkPQKl+2y+IvDJtFeMyltWLqTYVus3VcnJZ6rQkn+PGbPd
nYRf5xzHG88MUu2CPSLydsn3MxFMBC233iEZuuMHPmcm5cETkjW5RYuvts5628XE
kiTJfywDRh8GEn2369kJOlaUzB/0O31PmqqgOuWg35WqMZhkUvtN5czZ+BLf3otF
qcR7om79VRdQJ//5vbURgK3snq7NWyp6iwbYkHUtYZOV8Xb1WglrKgEqqW2y//He
f/vRiybY4ijDNbuHdEYGvlxa1iKe438YmMF8kjBnUYvSK331ly3XjkQrpN07tKds
vXU/X0b9XTfIAN2G8cQr2/NZMP8rflwySFEGdu/UuMAlbSxlPzjxKzUSUStBAJy4
gR91/HSvCvSsDbsESUXKY/kxPz0ADIhnlPcT+3ALreKPayNItWk3mgt0Ws+0bfP9
H3X5TawRx+iwYlQMzt9Y2J35P+Mw5dN70jpO5iquRyFfSMKFz0E4RV4/LeLEuR1P
2Yj2pa530qFhNlWbTwhydRpDg7VZWoaB8OyO/HkXzxlCJtnE6dlv7bqG6QymbUzK
RgZwjXSo4H9KzUqa6KbA4h/1/mwpprE7NV0/ygpwaLcArLxy6lvhfBkbyL22zOig
zfQDjCdfD2nMrj5BmbWuP4LRfHyCBCusPf9+K0UMLeA+sDCPSe6/HbSAIx1mMowa
ni28ZdZLxuzpKFiBUX1gcS1vhk/Q6niD3H0oE8iDvFHefrL9QToHbeNnxcqrtKcu
xcmWQabD4rzD9k7CaFV41SHK35AJLpf/zBnk/nWMXKUS7RwZ7Hgv2tB5ocLsTdfQ
9UGEHDmVxKIJkfA9pqFF3EV85XcGOzf5rWWOTmIBQM/KKdMNEMg6/fB3uMrk2QfZ
HWORceLxcTbAxKJ9/ZCoUsD5HFJjEqGLaEcz9UgcdAgiqg9+kpFy5qvmBsWce6lM
7kobf7ekY0pH/2cUZ5FZYTyMkbnoBeoEgJaZAkPiXWge4NR2D+4+wv51RayPAkC9
65fsz+prc4MYsqL/WQDNf5b9xwRMKA8fgzqauHdUd/E2zwXXS+5SPPFzdTQMXqFV
OArHSCiEra+dQzn++/vPvXxj/qcXWlH7TNuR+7hqmvlXl2PJtco2PHjPnSzL887i
6SEi/kXdIBiwZt406jDP2Uc7Z1q0c91VLKl32kLsfSNhq9XW3V7czn/skp7Rs5wS
NcclriTDCGCpFh678izyvI1IttjmbgfwrdSC3FeU9Xc+w88YHDaCVpVPBIHGxNgJ
feZMB/YDOiR25wjVDIpceWvqSmlr+QC/AMY1bemcUIi+J8CDRyy+z3gxrRNsqafV
iGVs07/OUHAbzxpmI9n1AhrFuTegPQoGpw/zACW/L+0TaF9OZ7OR3jwbK2sBQWL1
kBe6eNWfxKJsT8v+SM63mQQpZdmAV1BVIYUJoCwcEHB75ov0ZwucXaoMBJm1HDJj
7OXPAdPwagaGciWAGA5q7X4530YpGADNeVIIyaZx7hp7Poej9IAQxeGXQ6GN1jw7
4P7kUD/fACkwzr7uDp7yTGlH7FYj5VUEl1SSDj78um5VG4ICxOL2RX6/JcWZeQTb
PcLVz+dJxBlbiim9Mnmxfz48FcSyq0b9NV2f+SS0lxqllMPQguLSXbOsgwKXxQcF
iurrGNAmE71pjugjl1kVq0139v05LcpyWO009BODaM48CswGZcSfMLlooEdX71kz
D2McCjoEFPVD5B91ifxcuij4FuVJ9A9jKUFoAadJLc3BIWo9mQqAvl2w/RF58llc
jFQr2VH87WIBc2tegAo0JBRdf/1hyxrwDa1YzuRT3Yp8EIXJDp8qlXk9ea+HZFGg
kfkQ568UiJAKES28GiElqBf875/SKpUwlGk9tXCnmODwchtnd6zWgZQHr2Qf/9Du
Tps4zZwQ8l0g58RKZZk3XpucrmijuTm9wVpb46k0T/C20njCsipm38OxtA3wQjG2
8W+OwzjlPVYIWxKuYKKgxFQMlCGanUmZJvt3DwV/JRgBcjZr+kIXHhd1cUZvVJBC
VNe0xSN377SNAJounEiSKfmwFvXnwYjv7/fvoD5DaZGLj3OZKrNLifubQaufPoEy
yfYeHG7zrPBzbKBMKtd402jxPzHSqU/vPBytpRvx/iptIi1AifiCJUUthULB2evk
pOkd13VRZ36/UBQ4O8Nq2pi6KMKQKN0Zht8DOQBuF5v7aw+UhyLatVziA0TExhkx
HZ72PLb3GWovXkx+4J6bSaBjqB9MLx9sRAYJLT+VeHIB/zj8E1YcqfxR1FUWGefh
atmGcIyWYizjVdBYJUa9qoQyT/2pRtGWbXuWm/ADPI9NLOkzyHzW4QdP11CfgN7T
cKadaxVTUfv0AbEufQ/jprw3PhicMjxoca+3XfQt9cWeuR33YN8WJrVUP2cnWjQZ
4XWJiUYoY1/cuQJXLs9OCLcgDSvq3WgB2LX0T1fU8XoP5+qjC2tq9MjGd7esbu7R
/Qd25BbYdlcdjwjlNMP0nQ1GtWRqBzbypGejKXiIqqAVi/jIzrIW1a4t5osDh1RZ
Y1dHQf95fkdpTB/Trvq2mhK1ivJiZ+3CqAkwMjysLnEuJzaMN+msdUGkngJaA5l+
HEV5Y6YY2doUbOK668i9UF4FdPHV5sq6rZTfJT6xecWfKREdhgnl/CIdptbheIkx
2wLly2e8oLrFnZYhKAD3MLJZze4K4JpTtbCvfjXkpkpRZ/+mYTF+aiTaLqYI7IBo
kBEtEWZUpAzyWlUtmM0xNYG1buQ6PwgDj7bzj8vsYPm4f7MsX/Qy0F3WUjfRJjEh
J2T61vDJXYap5kzzZV7ieLKT2WeQyxtT2hY+o7H4Nmvf0MNTIdY2MlWHuA5DLflL
73+ciDrZYKeylrBrjiwpCuemG2vztd/olvc6R0h762hxGo7FaEly3dgo5BwWMQe5
ZcR7d++aT1456KmPPfCcO5KE3oO72CSz3DHinnZtRTbsfcdlFggA5/n8vabaIE4A
/9ruLTSecyMDoTKdlyG5KQbv4aMN8A1soPuyjHSw9hBibAKOvn4EzpOK2dQckHBg
hs1YTpsGl22MyeiT+uh3K08ep2YMGSjiQcqntuOEL5jJxhIlXlotFW0hYnBnVF9/
wqHfeiIeBtmrJ6if85spK2iIJ9qv2pw+gfMxZSE8dLmEQAxfdomQv5YPFwzjMg/r
iMnZac0kC3gy1CBbT+AwSZBVHTzwXKwi9FtJWq7MYSKzQiBVOiL5GN3uoDFFq9jr
n06OJtYWrQTatBGvj9Kv4Nr3ZQBKMxICw/d0hs1a37mc3u0rs42/li47PMTZXiT9
4+x199wI0An8LclkZfZ6JZYrJXGfjjcu1doUzH2dTKxnD8uaj2XOFW1DEzT4E/Ik
cRm406sFJgHqBmnn3p1uOAAy7P+d1bjLn3ratmAYjnoYp4FKmuAeq6wPVUDQlOH1
+KNqx2FEKH/nuQ9j9nNDGEYQwOa9PItbMDFv7CRBJonW5eG6djt/+0Z2bYzJFfNS
faofomfshJd2yxV+uU0nf+db3P0ZtYobwztt4mJVmbZcIM/09OSsHAwYLWFioVDD
3Lpyqzy/RMahvzWQgE1fH2dkukxZgXOHkfb1L0KnjYuH/eIKKQISLwlUUkgTdp/p
mKBY6XL/FKD5JbXSwl20PB1Qa5DLYsaJTyE0Fg6WyvPtkW92iftngHzOXIwYMnpU
mbB027KE0yRMh+/ihTEKjwScL8/R4WoI+nvVzdRrfJ9doY1WB6rLZa2NefTbTUHP
Q8uxLFw7NDRiXyLQhVS14sS/8ZykCaTm6g68DJdYtuAhFPaKfmNQPLmpLJRxXPZU
uvwEXabjOD8n907pEAF1JcpD+aSrhU8muFC109aEPXcH8YfF0U4IFucy3w/5QQ/6
hQSjVkp9LPsGsb/8UMAHvYsHIvQEiqKqHbLZQMwh7ZZogbOUjCcy3P6Ejf+3/89I
lQKl2HDr4UGbetajeGjF4g3Fw++x6S7Sgtg46XY2FytMN16VO6HWMC1iM0eOjFqD
jQo7Ej90HabiterzyFapsQPN/psMlXhbFML2XjTZtS6zwlHxsVJxTweZYVbhoucn
2p5+86eAUx8ab+aT2XsMPHBmJs9I/4FKyt6kA8Cqv71eK+x8MTBAb4n6jmU3YNbW
eoZpPM8jmtqKa7uE0NK2oVE8lDRSRQuihU3WX33Y128NRyqi3sbUUrS6uhe2kBbr
mHktYJPQcl8cBWdAg0oXlcviq+foyCmxqaPirCOj0FstF4dW82WWSVGNca2/UKVm
0PYf20flasK8NWa800Iy1WCTjy92ahaoOdYT8CsEMalu0hfYHVnObw2RZP+Uqre5
NT5KB9hSJNdSZXqeMZUdlcP8uczqn72JI3kZUEH5caLR64jaix3GUDz82DCRq0wz
YsqU5gtytwOTv5FI/DraTfyijnAvDzQE+R4XUYiee5U6Vt7wi3uGv+NvqZGbnLdN
owhEdsXLoRlzuaxihlGpJkwqtpN0hLc5PMcQnIBwi93cJZnw6gPlOhQew79Z5CMQ
QnDPNjJT9nS5bGqVIBMAYSOFkrm/jVvmz7P4feqm6JepAM0lZkPYWdHuT0PoRMFZ
52twnovzruIB1MHq5Qtaw0YcSuaaBDOvf52qf7ew4T5XRXXYznp/vMwsZ5AetkHc
3dTkW47vcoS4gAEVwmNFYcOJ1sbrjEmunTO9Z+Fd0B0MZ4LOUlmmGqgSAxvXdMYy
x6gEqUaZtiJG83sCKmZNDynYEggX1YgwkQaC0Wi6YIjI4SUrJm0Cny9AdChSSV3B
pGbYqbhCqc4mbRIVFLR/ybUz3AwGcHBGqUVo55syjv0wUf2ASCmqgG9561Lk3F6g
cUQWHRm7nCHfSw6lZjUHIQpsYYG9xcxOC8CpYj+MDIGuAr84w7HEGLo52IzoA0pP
se6Z3Uv4iLYJmLjbmeDk3TiAOfgsZ/0zG8lkM0srkwIv7QlOSAz5XZpVQ+UD6RxC
YondRBPhZgR87vl0t21e1jxucm4P3pTXkxNNkjme/Jayt/tnuBGN4sDFc6iiOrli
uXsT3ulwn8SQYoSQ8Im6KiW34WmRSE7DnQsdlexo+Gjy5bo13XoKLJpbXP8n3tOp
luSYCiZOTWM1JTbxlycRSwBxeRJHftWUdPe/OpicYB8kHnjoJX7GZJTPV1TKEa4e
sccCN1TyK1w/l8Uf0NSFu9cakXpK0Q/cXDn/Zog4BlFOR0uiWm4uBBtzkYuTResm
eBo5WB7L0skY0Xzb50N6xFbRPoB2/xUohjUHc9sEeLyRln9STEijq3iL4MVSQDci
e35kO5y7a4Ws6QC/DuiXv4bhXUK9WA0UTFI/IHeQOn/nMFONfRPA5pJ8xZmVHA0e
DFE26I2O4KkEe//AMXTKr23FDuC1VKo5843PRNurLlaN5diHoA3NiGkhDS0tdbFP
PkET2dPWVmYqyNES495Xkj5t4BEqvkNgWPdjxiPEGSS3OGr0pVE6etMA8ay8rQDy
85zo6cnWejvgZ92CXgxl5Y7YCtITxJRy4cboLEMJIVIHE5jSzb5whTMOCOxDcOoN
nbJfKTtQPWPSLRl3vebJ+DhlH6BJKOJ+Kd9uyaPBFuS7Ma1LMUmSpEOSQEAkL4hy
p9tdXTRcrHwphXEbdPTOxJh6GQlpiE9xGFaEKm7Wniuu3LW359wTF9W9UTRH0Gc0
uXS5XggZWV28ogcYnGiJaFh/ULnAWLaEC3Y4uyvPj3gszvFIUHNNVwat+EllPbN2
7Rt5O0S8Zjh8TOhb4/Gi+B8H3nEtYzkWX86QkLeMv9IF1C89LO/YM0O/RYFSZ6FX
3R+OKf7P3HTgVAPD/CeEqJ0zMINFCAATw4CGjiCRCzs/xBfYsPOrcyOPQlybOk5m
rLO1WaUlODndKZXf0UEbcDNLkPhXaD3e980ig6wakWa703lTPGjHFXMKg0l5LqCr
h34iODxK8oyYXJ4xHanWOjBOM1NK6ZElAVShdEUpblz9vZzLP+HwS97sH7F3pbbw
kaOuYXoiCKpZP1q3xag05jnD/ttVsnMkckZU5DhggyYVEUEGHlq9yfesJhOaR8xj
BDh+u4PJw/5zID7uJbiGBzy0pnTG+dsevcw1ui3Vb+ZVawNBxJvYIPRbPC3g3eaJ
6XlErD/0T6rlRfJLSEhTZFvQijGA9/3RVauH0HvTac7Dc6Ozu7YBLKbzqdupiupx
RS5V+ROPrRnV/nuwt7PjTe2HS9akV5Qgmc4nNNXsh3DmFBpOmlxUs0QKqs0PInJ5
ovk4Rr6yheIYc/p3bJR6tQuBhUAJffz1Qj9uPEcLNo3FyUii4jobgCgvDaWM87Pk
LiVQ6HVn/KKVBX0326fh4o+WVLIgS4keI7tjgdwbmLb0zDYtkoxLDpTPBaE6JUz+
RpX1kKGowvfMHR9AaUK3xLk0/KY1MeWfDjvSvEUYsr7aHANy9eF32FDX3fH1cvSP
pf8E4tKJCtBbie6wB79wWoRrgemU3bjazJvF8Uh5CJq5tjYM2YQS7wc25gPiF+l2
r5LZSGEY+styvDtwV8hAVxRaT8XaP1mR4nn1FjB5I3JI4DarnT918lzUYV0dL+aY
c0b3a5rmOlPU3UrqXMsT+1Lq+XKMRQJ00VOCqzX4V1BYAbYGciEORhmABM2GjC5T
0TMPfgi5L+yKZbLVE6IEryauu4QUbZRtTQqh2/ikaewpaw/PTHR27xsVFB+aBWu7
/7sXJ3qUDFiaR/Ngl9wAfDQOGiiRGQnFcniFmh9xkyvMX2Xdc79W9KvVwBhBnUE5
rEQialWnCIrxcCQDIXqf4BnGV2DKvtkCa86ovHReo4LtOevsG7mq1MxAH6ZaWeIK
IiMVn8AxbVVJqsqhA2gcPgsg0sfeQlP6rSb9csRhMJQU3OoZ6lpIXoizNiaIlL8P
MXHeiqaqgnOFSm//TtTIKuqM/ZWd43np9pEMdhzJv5iu2c/OMQBClLHVQhg9TqZa
QR2IUigrtqFQ/qgEqaXnx+Hxwh85ddqtgyAEMaUR7xGcv4WMYWH66PWrDzBRC13E
D0aOCyDmp14D6ZcwzN2BqWZU209IjTLtZPC1OIzCLvDuqZqJ/n9AQrHG7O9HUWHx
FtyNcSY/PVAUh00BubaRzVY7aqkYYlcdf7y66GeUu9UELjAq9V05yztY97XGXt5I
qWsDgyrfdAvR/DGmQOPpBGryOg5mtn1RpbzcMh2lEvShzeixF0JT2JMAh/CtI/tc
h1AB05yVT+1ANvBua1lsiOuJfn3FwwhpHu21ngwOJs7fUnrqdNFtTxrPlHUxcTVy
avCWVITSKq/SFjg9h+eLVB58lM3XA/ehlEjL5Wm41c7TmhVtDffiklzsFGVfSMd0
ioRbh42VrV0zHmPAq3/nsUmcj1HLTTPnq2CpDNx4W+f7pOJzFtvcfpjBs7xdOE2Y
LjnjVVLJ3egSGOC1lnZ6QEDFRkwJOVdFOO8bpemHfESGWI8Q8PayT5GAilWQXcWi
EfQicIevE6IIJhsEWsUpQC/4D3YSQ0oiLk3G0CZf9Ju8hcOTg2k2XFxWVPOIbdZU
qbbNNlCbeL6yw2Mz8ocYbA==
--pragma protect end_data_block
--pragma protect digest_block
C6vW7g+p6UgNZYhF8UCXqA1pujU=
--pragma protect end_digest_block
--pragma protect end_protected
