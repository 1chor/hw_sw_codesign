-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
CQdHisS3/4cRH1eBxMEXHXJSM5BE/IZ6R4Uqz9wfNxNHxT3p+lGJ3wDvCHHHjqCl
PpAMmvjL6kE/i+EsApKuxzyrE1kHsa77iY28zkB3BHnsbjIg8A6nnF4j3W6DUdZI
Y3dyytDEjRSf63BpdXw7d9im9UUHVMu0/oNvNvylg6Ngc+v3hmeJxg==
--pragma protect end_key_block
--pragma protect digest_block
sZKY1Gx9NbjDL22qhVstJRh/Xqk=
--pragma protect end_digest_block
--pragma protect data_block
Dq+p6ABIYk6gOEewpb6kbqitpdMvUVujcjxLimsxLsD9GYVHtP9+9BBc/ePfQaAA
ORIk+qbrV4AF6nG2NnN57DdrxZ8pCKq//5W3uKesRZN4DmAKlViKupCTdDxfi7hP
HubcgeZ+BdRAlyelYcIYQsDEvu4efUqxo2mSvZpN3KZIJGFPQMQMm4gxeqyaEjoR
lWAiKyCj23JyIs7s9k+y2uVhs3qS3RmmuQOjgLqJREHId+CN7FIy1LxdTb81t1or
ommidvGTdUUWpJ5CVUTdJWAdBQwPWV3TGfi4BlLgqiXR/l+UFzxEfqWi+3MwOk3R
3wMZu3RK0y1bI9DZeIjh0ZihEl/bBSTvYzdgysOeFh/0RxCuxcEoKVEIeEFU/GPW
rocT0NNac2swpTPXE9Q41S+YUEXdNbknw7y0OFkKvLlcheSpQprSbSktFMViG4eH
1GGZyv7Qr9BNDDJHKkb3HyNuEElNRM7LaOeMBba35by/6H+bBOHYsHlqGm252T36
C175VVhmKmJ01jVXvOSILChl9ni8puGdS4FWwa4IDUa1RubJCs8GK7+ClriH1nGE
V84ARFcms1pXTuZWe4jx+NtF8dghVkHUsY3KfEnSrBiNPRHOOmfuw8139dEn8TLw
q7tWte7fXt+lbeVVdoFPje/fFJxIpaDV6m2UHVki/xZVBb8QzwqLpUrsldDisRZQ
pOhpq2lyloab7hj3MH9MIcpJ5F1iIC+ugXSTgJBkZGhSbok5D039EoOMoKWJPldV
5vpSeyD26o+1jheqAAUXac4xHgOGM0BAe+KXe+5QMD91e+3piZQWHNcxAqBhDypj
nJeVYtTMeFiXvwgiCCxFowwFBg1xFBHUHyS2O2YTKCYTgDaqLo5xxhi3qIU5jaeo
ACHSHoULH02jsk5YuGl/mSRL1v7M2CEVw2iyO2lBvYdtgdzic2E3IOxtVbg9r3o0
qNwsXGBMzh3AHcH3+srD8N1JpILv+FYtSu809csNpCvhp1kuEfwIAa70S3XzhbSw
WDnC1qS+GCXeZza7KC9xje1H7HgwKA4crgPDd4QMp54Tteo7C4+rqLQM9V+acp4+
8EW6fV7+yl5STqaUpG8QSJz3KoQ6JP5qPJjWKd9zFjgrLDRACcA82zqOZFVMJmMD
B9tSwCzUCyHht5CbV85QGQA6WN6w9LKI2rmqdaZQsHNaHx6zQofjFfYLznArU6fN
CFm2cgEd7e5eTN+rCgxHI9IHldOncz1FoeS1inlaKBsHcP3gCeW6ZquqA96AxUIo
ib8lbS4k/0amKYVld6YCuHLVaCVw0sWUe3Zrt7pObUeQuszQoj+M4yXdXWiAu7G0
v4jZ3yHNlShQxty09E4XP2Ur/w1ZpFQKNI3P993dhR8fJ5OkMaVmo5bXDvKQBRb7
tV5bImQwPZE6ZwsUvjZC+9FBxM0c8HPJftczLyUCzy3dN5GP15QJ08yVCr1SyJ+b
ZGQipWSVmL0eQuvjw/A5Dn6y7JepLtgjqcRQlnCZJ2cfYdatfmxHdaFm7KnLhvKr
7mLBR5RK0P+Olvw/BL0SLjnlpJrdDdjLRv4hSNeGi2IK1lBdiUcI46UBmuo+mO8v
ksgx2ShkrOjbHqsYVfuaJPvLFL0EAYblIOh2b14HsJCgFVBR7sP/GS5CFIK7ds0t
IMio3Tnzr/6I3DqtcE6ZTwJMf6Z37hBYQB7kAGi4oS4YttGHL8foyyWDDPzfFT0s
YRANDz3ugUSk7hmGR2yczsoWGw1o2pIiq65vjmwAyPWKs9f6hvJF3kBPPi/PxsW9
Mh9/5KfQZYEAfXViEdzaHR+I+9azkdE2GBrDvcEwDI15tNaHp1rgDFylSolcb/HX
gvdWKV2VWZ6TBFyMnwkOS09iQUnAstpOGXELusMgDjo2rwnl5Moxi9XchstD2Wtx
2ucef/5tIB/DwwycRQItC+46l5L7inQL4I53DGhpyBQl6zo+k54p3WPi/zUftqFI
G58TwWpw4ymW7hHNaPQO9b/Vk1/XiysYWSPCRDxUHacqFGDYQccGeqDTvkdpYtno
M5VR1+jLhYVl32XKOHuUgCbXvkWSPOmi7g4MpBBDj+9d9Q8g1N6lC2j1TENlZiR6
0XZo66glG025TiowVvQEO5BriPoWWkUTPkhqb845kcRoWY8CPBbHXcFJ9J22yujr
a/R1hmrIb3Jxu9DTI3ivtC69zeZBF5QTXbWhb8cuPmGbZh5SWr/hZPMIdpGo/T1i
9v7oXQSgq+ZtnDDi8gmX3P6LdOEMurO8DjkzBHHT3FszVHrZQDsvY6FerSSj6CEl
nJUACYvAKCOzEJV+2/Dgx47Wcv9TyYtyQdXzbCEFzThlTJZVqXBRT9XadH/RdSfi
cNp/uU9B2j4qCd2k3rCX3O2Tg7CWf2VrBYUmnCe8H5JfnBDXz/WEKNy5+jpHLHDd
DhwAloQ1Y0W7kAt310rYs/ta0KiOrUaeKiermIvW3Sz3TyZqnVf6vv7tt7N9dcJo
wh/05Fke0B2xNmgeLW7927U66fcuQJb3FzywnqKYpGktqPJxAoKhkYfPnvfBNe6V
KB5wDa1PITHFP8khgCKeXFjxpajVUvJ1awOF0hfU4lRs0gpU0IuATxElxHlF7FxG
xJySA/X1iFX/zpdKql12C5U3bK1sgldG5RnbHEMCdc8qL5LLoYDmOSWrfFKYbKrg
iqbFauylTh6bPX5xnS5/++k7srOoqc8CY6+UhPG2ZBhqntdSn1FW8f6xxFRdQ6A5
y1P5Ii56d0+kmtRw8kV6eDvEIbulP1iZ/0AWnfCi0xUUKMkxDh11CjVHvfMoQ/0D
Gmuw2LfYuiNn7y8CyQuJWjTjnJH2FMvwRID4IGEJY7GaM/Ad/WL8zdXqhvIavh1X
zQgt/4lfqQSaiJbSG/z54Aj63J2qp98g5ofX9BT4OFS2qxAQDw56lnrSbSd7B1Sq
fsytRrbY48bH7na4sgbJnaYPmH70nmdP+FrrYrKvP8Jv6JMoE8jOPWB+SkuI1F/P
0viwRMakH9DSGU68rhPE8LCJW9lCw2CGKMUE/UwfMoYqUMMflAyJXwu1jKH2VmkD
WxVBZg4cSwBCU9jTccNWtUProMg/p8hxr2+1eez3nyFkKrMWnyNQIv5VPjE+GjXN
9/5W6eVjlfasXooqG70bEeBz2qyeOH5tuPptBBul4spfBwOzQIFgMN/wmPRwj3uE
QsOu29Lc0JKl0l+0dM3qytKcRMg4fk7vBvxZwta4ynSUQafrtUkYnk/rpvfl3w1M
OS2QXxZ++IfqLC9p8SW6jHfjT1Z3UWYLnEege4luY/ho/w3/F4Vx19l6kitkeJcp
YFWuoM360+GzkKdHOF8AOQ/ha8R/s4lAuzPd40lNvdMeNR7VEqK7BZ6GdC3lNML8
9LX3VO0rqu2n12fhV0V40VlWHV8ZZmHVuCxMcucPx7KZnen09AVsskHeQOAXfAz+
lVO7j8kMRoCYxTFCK3/tDXIjc5awBkpgjQskVPXJhcDiX9sKqCr0+0D05yqfnL+x
4VuEa6WrNr1ZEJ5Ac70cwuRRA1phV8eWpz5/VUYFIhhL1LHDodZjSW/UKupSQZHW
bwV3P7g/zUNwZ6FuCc660EgQPHwBv6jasqBLRvy2+VG/0U8oVwPmcKIEX3KxT/n1
CKDBawQC9VckgrMbm0fippeYMpBiRODUIQmgr7z8px48KcpNsv9xQ4v23q7EymDa
iHbc6wzfRzdONfTPNHhlsHpk3jAzFDFP/D10E1FWugsuovOMWnE06e+lUWc3wKVS
LN3mxJXErYhw6ab0JIB7vU9rxv2/dWPEtGCcb+Ab2qDRSEK72ijPHpJV978mZxJI
YPjsfpG6lIp7WjdqwLEIdsBxZ3+45+T97tVXcWTnwrNWR2aLsovv4Q8SRyoB2KmU
7m3y4b5NoCnDTBzl4em/b/G50c3OiXkNoAIop7z7/3ryzTliReMt2OLzbsOwKFY3
m1L2E36vClNKuZJDH0Sj814Zb/mK6N0fggBiAdJc7YmqO9ctmbm8CqQ3qqXQju+u
+aiytN552NW8DZQuHj35wY28SKnLxf4fZSrrJNmrKrhOGCp5VLBWSekhhoUXw/Wn
8WHVrDqmo00ds3IJibyVPOALAwr9nx8jo7UK/VGFcX6ttAp8PuT3ITstKqG0xROC
fAyQZi4+vrybzUiQyf7dYTzCt/fPaUlDwKxNQlVp8WDi3gctHh0D8XrCFubXlm4q
mOLkACDWOdgE5EnjW1obNY/JbbOtduGbIpIWa6Wj0hKSAGv0DO3RCOJkyyrFg7nI
fNnBcvn5HBqG6jiJUpXx4lAz0aNYqllbgn6QRD941T3ATI0tH2/XBWqLxqmTpW3T
IgQJTK7JFSGD931TBc2TEiyuUlhU6WeRBytzZ+r93/gpKeIzxSY0VE6noMi3hVzW
O+XxGbHLamsP/mqNemE35VnQucsaFmxc6Z3I0WoCHR5GESqrtp6+Gc3oowCEMN9R
1UXW//mRlOlybRNVXuNC4X3Zquvcv4Bh1y52UJ/4N954DcOZ8X+WtC3+jugY4/jN
wO+uGG4a5vvNKbriRmsFenj3Wgkq5vUtOHStTj9OjRH3kzLEC+tegyk/HtTIV1Jl
1Brj9W+DNOgHXlvukHBpzu5RDTgxzkfHcg8+a/yGR6AJzGLaQhL6PDbMSG5lf4Zo
rtHm2WjQqm6hHRGol+G8VWpne1u/+lg5y3rY1vcFcUitcRDd9sNTAeBGO8XcE9lN
fF1+inrCIS7nQnv/BkjjlQkvKZbzZOWDPhDELooj8Z0kry3++VPQmd7XzGrX1xlD
PSdhg57ScZ2pPcvXO9QdAebnW+XXFaEe2x+gz1aNw/v3/TBYc89RS5flkZ979A+J
MjuOGlKb0vzQ8lgTgC0Lyf9w0WZjAZPo5AdBTybj8+DFjsyyuGs+fTKO+uLD4tc6
u2KlJhoeQf5C1n4dtlTF75Ax/ts9dNgsm69IHfz4Xpl9qD+w9fwahyYsmH36HwFH
leiXy1BiR7sF3HDCtLor9CB6/ixtSA9QSEUIDwgeYbyq1Tnm3nkRsfkacDX93UEx
3/cIelNR0Fu7O+hW4H/Q0lI1frgBd293ANmTS1qQYTITsBedYAjri3moz+GO/9QA
q9N8MC4DSFs3MjEsfBLuTevV1XGxNEmpAEsD0syloaTN7gym2gjYtKPxWtcfGzK0
ZbJNC3tX6EiPUnDKkq4RpsdF9R/vJajsgo9p14PEim4pB78CYoFoSYZK8pJ+f4P0
xFh/w5oca2mZtDu7P/EbS2VawCfnHIslBrPCOEGysF+Uuv9GqK6XSeAgjjY2LRze
eu5StjZ3p01+8tbYFM4u+b7uu5Yterh4gov6FvSi6g1TLHjyX6QVYubNR+Q5CGl8
nKmgFmfXwQ/vAnS6T3dI1qwC/vRT04Wn2KO9y+CMplbsni/5MuNpT8Wt4WhYmkfX
dP3x9KwTWXxVoe+n4EwWP2E+lwdw83NWiazO7VMqWETMzFkWp1BU1/49WRx+ZKGl
ocsutxyphBfkvh9mlZbXhRzmkpLkQ2l5bkI8FtkQf7+LWMqtJimjOVRnYD847kN1
b2KGaCjaFKNPlv0qzMybYAAaxmceHv8Q1QN94WEPOtIEaHM+df3UUI4V5y0n7SCy
D/rBirs9JEbFGpXC8uL6WWsOAfpAqlPqYhdRPRwXiuaC5htioc2cavbOs4KKlHSr
pIC5IookKUareoH7zQYxZIxP0iXN/lGClM1hPZ1BW95FQKDHQ0gULrg4Zu7Uzay0
N5NgpY09ZqCHvqnaqHh4vkofos9vSUiJrjK+IA7bLiuUKy0wSSZAEBtnKYGRDK36
KKOPKwvjokEmiE7VSmY20AmzRJ+dKCNpi5T4M5/TI7jpZITsV816h3DL00orXccG
+JYUdLC12QB0ZprdKcFXvpDEJ6QPGPNMrOAbftmNqGfsExrOA68FjdNaCn5zl7gq
M3nMZU2jcFqzmaW6y4pNmMqzYvQgfFq44hHiG5n3IvI6r8OTiIwpk+Eo5ow53em8
brTlNSa2RSQpNXMfKAKV01pp+2NYV3HA7Z4tfTTs38OBYAW5J0Q6CMsoXjyRyj69
1TlWMqfGZHhJnzU+2jg6do+0oxE9R1Pft6Q8NxMulYSOLv+oANCf/8rMrW3mOCXV
716NTKtCEtBzrprt+HDGI5bN1XJr0j9MttsB29K3sSQfxGX53uOFxZZo690d1790
9VHZc5XXWwP9opZF3esYONhnULfG7JVeLZNyumEc3cWYI3uQvCGp+uAFd3sKUhoH
X4N9L8HtmAmL3z9qq1fHGi5gEfS2MsZdUTsuHLSxKPzqMbd1mSvM5fimEFhrODpa
uQnTHe21IX5aCF0pKhzWJCxwMJsrpvZ5QGZWk+kXOGkx8WtvT96x8pIvYsFEiO9Y
Wa3moEyPnXkTtfS2fwtJbE9El9DiZuK6TtSb0+B7yQ1awBBZiu10NezDlaJos23W
wrLknJGDq4cAJtsNTxeSZyNoSmokOcJ8ny4+3I5ArQRZ54YceCT5llJ9iVOeiLF5
F55DCU5zPw0z3L0f2sqC9q5Ent7LGxb+j5s0XG+98uGyhheM8fqgVpjwS7v31R3C
insV3tRiVDzJTRgF2S5fBM0NsLFS4IWYFJcTlDkoEE1k7ZNi2oiTYqIMMqb3njVO
myv4/6+kInmYPMjf0N1YLU7eVh96YJWPFdJGyb81jFzR1SFlibPCwQrgyCTLYQv2
QEBEUKdvsPA7KOf6CQIonUu99QmKgOU4L8h2PNVhe5gQ1t4yYRfgzLgfsM7gXZPf
dsylJr7GtYML3DmIZrfss3G5GsgC0iEWVG0n1eOa1cPwaMbVQLnPfGz8ojIXQvoB
LdtduzZTZFTT2WapYB+RIhnPwzp7viVTorMub29huVydT8ce0+SBxytl9KAfKkuD
p00/j3Pl4DBqKYB1e2reeZQ1nPjOgKy1Mbm4+z7xpa1RZMJOfQko7ze1vQHA5207
mZ9rRF3ZumSpI5yC1mwTg8KX6+wvP4ZfNHStfcOVYS7c5sf3RvOufEJ3Mp8BzoNi
RkZ1Oesei/buMRr+mwUpR62VGRiacEoyY8rgx5PRFkuS9Eg6IbJkcfxfyTEa06Eg
/QID5pkboQZKeBmgSkfmd/L7BYipSlMqJTdefRghEuL2FZAfVz1hd8uCgJ9V3Icq
Ao8c7jwRaPw9kFuCf96bVGnzKOBhRrLFwKUse+Yp4seQ29ErUYaC5IDCTGW0oEKi
zjBlLJpHJYZjXXS/ZV+Mx69FMZr0LFOAQy3phgEWmGt7TNP0XA/gFOGkqcNYtErf
MRJ1W1uH6+8r0s/fE0CGQl0SVyjee7gZlGfl+b21thSNhPEGcBLvUzdHrTLafKyN
nbthCLMQb8PlIfGpS2djVjz0F/oQZ3j5iv1Bhv+dxkb9QccLOZKoHtZxGP1IHUKN
7de24HEqGeCvY2oRdXNFV1AljOnDhjJC1dHUCXMuaBKKLpmFp/o1EKo4vJiRDoNs
+pljv3F/qUnKwugE+eDZRLOUUfQreq1U8HOYkeACy/jqVGosoAE4kdnKZLE/k97s
OGQo0/drIBGnhWXQX32zBLkhJasuihr7QzUs4+ujJ8a4q/YsNL9hro9sawvKKFpb
xJu6AD2KS4arcAD47YnKhAmSHZbVWMBSteIyg/ZIdysdjg+W1LYjwD5A8Gv8oVgF
GGsNVLk62Q35rV7aXD83SD7yZ85PL1eruiHWuUesKWGQgB7jmNiW5PqKDixoqZNx
bcFGjFD3VgoZS/e0KPSfxHgx3c4QQRh8pZnzkZbvxzjWnZz5yoEc3afzPZ5oJ2Sw
LDlnAAbdvMp8cc/jzPkjWLuPGsiwLYMXnjBQ7geYx36B4A9ijErwDUlQpGSppztH
gWlSAP3Zzd3/cELFr6GF9s6OQQiHoyVx+7T0/LzJXwIUBVuhe4wUgcE3GgJcdmcH
6rKSxj852zzSzYf5oFmjKzcagsAxRTLrZoKwvPMHt8o1MVoe7HjUJiJrOxqHLAen
EN4iyE/x9K8dTLn20TFBWc5nk9DMhd6MrQpa0VLkhz3x6DjG9gFNAwEdeuYDMf2b
F9Hq+ssdzRYb+YC0eSDgv9uRDZ15lpUUngc9SgECmkhbPK3nLwhbui36vjit1L8p
JNGp5FbVlgb5/EDwm82jAytqHOXV7DYZ5j6ayvUyXvFmvBZ2kqCRjKs0gUaSuMbr
o9y2aJ6r/b+Y7U+T9xmoasV6RLoyr+9M8x6jszvZBB/Mpgvk1+JPL5NHpyHZCrZT
YlV1ujj8k23/ws/2N7PYnkq6qM/HAZFI7rPjOAgqaZgAgPDt9uNv0oHYrmekcrXX
bYSLGVuS7Ad6o1FcfiAKGSocSmdB3Dq6L7gMsHO5xXpUeQsShow6cJqowjFGMPFt
N71VUefue4P787eL0gnk0n1C/X0XdsYMG1xN/mGRDorBNIXsseOtzNq7BwTgxT6z
t5RNSD+JykvAdxHhw5qMsLKfy9ubV62wIeDdGRjBbb0fe3arTRDIbhMLFQgwYkmM
o+Vv2RKq4fvtQjw6Dxjzw8TMPEBGnhx/J6tORn9f99FcvwVTCQvcxtJ9VX9tECqW
e5Uk+vCX1dv7jdpm2o1Bb+Mr/l1xdvaUrt9gcre7ArQqwnKKDxlyUXHMA7luwqRW
A5ILyiobL2pR3tahVVjxRU7CQ7IOs29iDozPSsiLqnx1iqsuI/vMVkXp3bEd04QT
OGr0+Jmcz6BckBAKYfhuzW3d4H3eZUPco35vld0hqh4S1xNI9vY73oeNN8PhICq3
YOrsl95F63e2GRZC8tLIWCxOkOiR7S/ZBSo1z82XTNSn3+mmWcFf+JD4wRAuhRSz
ZPw5tGrc43P4HKio7h07FnyC1Ak8yQ/KBLQULEF6VChl1Hazyoo6FyBouNr5A76Q
3wYEFslxvOhL3dX8T3tKr75XT/upOoKOh/9an21glAt5WaQfBVuLEXZ0YGjOFEt6
y64kikn/H+UQoNGwHsDJSgwTxahmodLbLLoyYjchEXNsvTFEJYX+tKnHgzD/RRTm
DFYVopBez6i/dUkSl8WnKikeROWV0tYu3VR1hcb98Px3XNtbIlZw4gFNkqmZF35T
I1wYip0FOIlfvrFL/mgKbc/e0CEhnFh1pQP9BbvZBc+GSm1ZSXPGNLbN0kQ5gV0U
/kn5ImfM/FgGQ9C/8NM4jHKXowhqqOJxhE8fI2JNpCIQFLX6lpMP1zuRmLqCFsGK
DydIlgi5meWcxeqLZDUgFAbmR6lPwKp3uAB7s8OzUYTklzY0q5rzUOaCtpVSSjVE
IDzIVvncFSzMfRe5eNE2dH0KaLh3VyMsur0ehpA5fLsdwq6LkLABAoJYDIwn+34O
3ZKUzV+cOs73vTJBFzXGOwLKHwo2LDqOCxmpDyL20BmxtisEtVspiO54h7mb0iag
26TLk6iRIwn14JTv5x2eymYPkjIerMK3wevxcRuQxpadOjaFntbV3FKX5Po2x8Te
Rk8iNLcqhEZNi1eDjK4pwSfTBTtYJ9Rb/q49+GTCOLk/APxGvOQzt4fsikVUaKjT
Q/rhiODj9aWW5j4C6Jd0AynZ1WqHUjopo6DHcxQGLbj5ECg2f7dlZCJZ/9QA/tgW
YTN4UgtZBPTeaeruaYGj71yTHImc1xXFT0f3borHJoW6/zSQjvih9c+2ucz93J70
DQya44+FIfa29b+BLg7haHiRo7+lpaV78Rllf3vMH7TAqUOLByNQIC+ZaBKPiJBt
BgI/7fXtUFiKc0g/rfnEUTbiwRX6nrcL280ZdlgyHL1djQlgZ5yXUOiIqdPe5mnG
0ly3s6/P7FwIPvFuenzusoHmjy643FAbaGO9aJjTfVuHL7/Tk+++yGbSOV66oHYX
CbT7HP2kpUaq+JroWBD0kRRzVF7zj0defCu0C8MQXb1LAZJgfZfwlQht+Fk0gjsr
X76/ceEFrnRaxy7HCBlzfFr+nxWY6yldOvRf6VsfycYDbdJALJqic8d13mPGB5s8
GNV9MTJhzlD1t8QeaVvHZxbXNz9hJrw0NNYx4hnmFTztF2GlsbS0UZpo4cCteKVE
uRWjs7rn8+fSTWb6pKjbQzXR8OCkPOkUnkmwto3z/QCgNAx7fw18yDgA0EgeNUzo
vJVNy30a//IxaSCigVslY/3Pm30jGJjdID4DII9vpDKHnBwENMucx4Wnl/vCU1Vq
3SoBedn/OWg1EleWV+ZNPIz8mkyw6xyRYWgJKKuY7pN3yeED56UYQYtNn6MfIuaX
10/e7toTF2iPzL3cbjBHwK2qYIVjYqIUEzvzBTYFKohbrFiKZ3dzdAPds/co+/sX
m8LUwbUJfIFW3EnOlOv9X2e2q1emw0MxOij5hZSEPsLc1W7dYIINHIz7nikacNRZ
AI8VJY9C9kgsn23QCvS2i47RjeQ8JJs3S27RL5NqnkgAq2fAEwnADIxHcfOU9pt9
sofBh5KBtyyV0ogFMq/KRwtfhABUEnQpqKjxZnTagn2OjQQdiOfOrRBHL2wRKH6x
ID1jUiT/PX7qNyFFJpQ5yAr/nX092yfXQli5qH9isFrBZ/3vydP0mAClSAmD9oaP
hEX0sv8/umyJs/UUmHZ1xhUvaJbzta3h9X4h6+6Hem7lXZkd/Bpe538KdndfNRMT
SgrtUYui70wGTBOQ2ZsiYdKcNbf82Kl102SE/vt9Bj2y5UhqE/yRBkLj5TQjvlCt
KeLFCQcw8vZR+BdfPc9R5k8sSZ6QTp6npHPu7vBH2ElJkOizHPKBjBfgH2m2opKq
+dhjCl7Es4EK4ZDriPm+ezwJO4pytc/tSwCTysiW12q+paRIJy8ZEjHAAjswc/ap
pTMhAgDScel5wQrKF/SYHA05uurCK5W/ezY52y4j19sBLISlKImyMQET8lnnuyt+
6GJQqbjVwGPWc2x2nfkRHq0qYRkVHC8YrkI1Mr3lr5aIdm3L+AEiirBNGMsef9iZ
yW7IGSUuIW0+Sc+W3hWm9Nco45RzHpYRGqd9yFFZw1OCnVycKM6Q+t5cjg7rP3Ps
cGTD6drPb+i2T/12+Qe2n5O9V1cWqFb58NFgimnwQCvYHxoMeUkEwd68Ki2Vke3U
9ERhapPyOisVo3N3N4hFUvRnQx+9A+X5hPdWwMGdcQBvviB492ENhm0kuKrR5Zmk
f7hc8RT5yPWdX97yPqEk2O+G7gLAl7ghu1Nx7S/lQAT0m03u46vi5qlBqS8ZAUzl
HBFt/N3XXsucloHoyHnryITgtNY8jWfG8EzllT+/WOcAg3wDf/99hGErnzhUD20E
QofpkoB3SpDM5P3wg7THk+9myaPqMTsqOCTono8LF8iZ6jGo8HrkOEnuE4+FP5js
BpPsq8LmuWX+Xmgk+rsboptbrf16PzkWSljzEF+BZioXcZ4fETqZ7o7pGfFfPI5L
Z1tJ+mXPueEZpvNDidcrTGTzY6D+ljcix4+v1/6/QCPMoBjm8twwLweiO+PmliEG
iQ2fekifvCj8XTTNtHz1Ft0dQ1eYph6KAQjyDRncR6z41GHsEfz6hqVh8t66aQdG
ugQnr6Fv2xn1xeZwjz6asrazmAQyk5D9HSR56LXCRjG4aunaRJgr9MI7vEhbIgcq
yFNuQvdOVcDqzVngEOPBHo2X3nFjSEV3HvHWBJpmS4YCVRTuUMEAC8RLO+YPBtkI
AoIv52eu1sIWHUdYQYhWQz6OO94FgWIA4Thg1QJcU/n9pbK1jgcY2cCP6o7Az3fk
lO6RISdRz+gfVx/qLRAncY9pea+EDjkksX5VF8EyhT37Nb/zmHZUuECHS45muMpW
FkXTgHykceHQ0EccI40TbBw58Ngk/2BjvymArSBCXhHh9dodtnOtpR6p7tBmiKZb
bXLSvnMnkekpeS9dElMPteDKei3XGY/1K3Ia57hwiSKk5MGhJk9nPQ/CD038Ftp8
R/wXiriNvhzOFgX+opgXSXNI3Yb+2xXDkMYdPd00vfcUH8Ph9P/Xq8vYsYW+UNIQ
2Erio7vIn0BhpXjVBgzV3dxZyyns3Qf3xG3hyj3huNLuYYrKXLuxxlF1bAEidsJ8
gHhpn+YAtTDrRru2p9Bt4qQ0yHGOf+tg15jXffqLSxN5fEJPu047ln73jOj/sCJa
I/UGMfFBVnjpPk0VlVythvXSb/ZD2vo7g1oS6CuNzoxN09odWiAmRABiwqxq9txy
NzKWMEzyQFrC66CvCMw49NxC5+eBGvZQ8X8YvknbqjI1aBhuxvHvGZyX64RyNJxV
OZtllSKJsTA865YmWAgWKK5OT/FR6YwZC1bWrg5oOOce1WcVqCpx0x1d4AE4vrrd
X1oIWA0/wDbt+Nuul3HHueuomAAAWNjhSrCxaNjDgssB3OzGVkOXp/FUJ0HQM+bK
fkiD5YVu55kBw87Kpiu82MeDiKPXYRg1/xEb1zzWifb9TOd8052QWM823dQco976
lZxhdYYlzxAio23Cq621H5U0p/c47tOmCey4aOAbNTs7tZJp25798rzTX6Tceg1r
lb9BYPNi7BVcXmMNtrqx1Kuyvqc6QBper9fOtXxsGTcWg08K0UbOvPfOTHOqNItD
nfwLJGcnHR2FNYmT7HwaemuCYz/xQ5D7J1M4pHXlJ5P9f4Xo2hczLtvNlT08zkk6
5etryy9RwSg1bgtkNtsBGh4aoRuS5eMLnP3/gTRWHaEs9Jh857oqguz2OlndDtay
pIv+FCyEWUeaLrPfC7boyHXstYsTQWFz7lYtjNrbzTNhDzQTroCbiPJebZ3OlASg
dRqljocrvbnEirjNoZ2jWJzpn7cUS66pFBkF0p2dQUn7H1bFmbxn3O0GTdduPQ5E
eY9dMcaySgOM7AQI6I14zPrrCg6h2XOY/VpLEMUsxTpB+pm0/uUxqcHT0CojaSrK
cJpxSzSnAYgZcK3kBBWt2FMwehGXn9ib6EcJKwJSbXYtMru+E8rzCB/OSGzyoPYS
No6KufH/clz5S5U/SjrPuCVeIdFsU27ej5UMm01iDJ/1mjp9b2F76QW4hD+5hDQ1
KOY5Ddq5s3wo3sLX1YbMqoNfrE6ODmL0uFlVuj+uPg1okkeZSJrKJTbsxniSOIXj
68gHJlY/u7z+pNHRmA+1HRe2P3UphDwpcJWfD6GRoFfHHI9ZWOL1qZZTf3gCNw25
dWTjY0j8jNiMBVvOEnQW0OWY4FI5FLQdqkwLF/+ALYMlzAWp+N5IeW8kRS83NNL2
6W/nySpHiBM2DYHF9LozXK/FGXJAhGCULE4XvH/C9jjS4huUZ0WkwrRuTyCfsRPq
5jMgasVczgPMSc1srDzU5XcFIfDkMXggX6cdTqRDMq5Dmp++8GjlJ3XvF2IS+ZlH
ey3p9gw0Gi9m9WYuyHGk7Y1BhDGZP/qu10Bhn+CP5efFa2eCteTJ8qlMQzLiFrdj
4+8OOuRReGa9Phhv7U8w4eJ+YlJj+StSOXk1QiSXPyQ/z5q6Hi8NtO5IN6r4pi3M
WBFT4A5r3M3SpjKyQj11J/MJR8ANWlUlSRGvemU+AvBuhVI+NankvNK94EaKXJi5
75MOBj4UZQqM2IvRNpmF3Bf5Vq6kBaD1Odt3ObSGR4usiIShwM5vCQfOuazIsdB1
OepwsnyF7QaE0ingtwazHV3SEGZ99KGRJAh5NdFLJjczopYU9P/JAAS8ddrKSxr/
2GZUW+tyQYglSldh1r38VH5bxzGH3UPVF3tX2uRCNoocPuJJ3hL3zZy2xyjpvcz7
BH/uAsF7Z+Us0bnq0pINUHAO2nSdeDwCAfJJp0rzEbrG3wiF3iB8tny49Dl8NsLm
rDWMkrImznyGlUg/oAsQi6dqSxhZX7Qaw8YZfd/HyBf3lbcshryecrFhWI42KlL+
cK7Oe85DoxQJeNG9rjic2JaxJr+Q9rym2Qk3vT/RbuncfiYYhHodgH74nund/w/9
cuq2wCqZ/ag+yLbbMY2K29ZvkMfZgU8AqZwjQNtj+aHUWVegPeinvEkwnl6r/spP
GXBE4wLJ9kZBcIjt++KnlT0Cb7f7QgzCcG//svdFe+0tyiH97J4s6o4ROzjCbY8e
W60ToSjnVoKTCU8WsWD5UJ8cvxnMuBL7W86k/HAshm0gi/6keAwP3x5Kc2UUbDCj
mRUtgnGU9t5d/McQQ5mVogli8uvAdV/0H10bmZh6bykB6r1de7W8+KDiq37iGPcD
I35SSoeSbc7mTDnjqGGq6DJQiIrmpEjIl60DtvcgBbBCof05vOrm3UwL9sci8X/S
poh+2sCTqmd84YXSqMectGNxWUKfQwD3ra2g9fcDYQLdUmtLGgKqTCS2TkBl5QRP
A682fN6l55YO2DItsfXT8ry7YRV4Vm3e8YBB/XibG0JvbqmXQa3DgL/+R1Y0+Phe
YJhJf0KjBc2PtaZvnANc0CEs3Bd4QMrPRAWqE5kCYP9SRRWQ4Azg6RuM4lde4wYL
U8w37von2W4XPSkYOWJ6vvFheRz7hGtmAUhy15yJxopa4NqFwwGmtEqrsacSSvP5
dBykrx28rQ89LmnUTJzRS4SQszc87kSEP8IeTQnNoXMQaey7IHW46yebVwpFqeS6
d5mOxrqqDA8lTWsZ/2v0VDox//uU3rSdXmi5OLaANvnKMD9f5TUig3Gb3BsTOP9P
y2sU/bAEDuS8xQmyUNgSNFckJYZrxR+aQ/DSE2Yn5x5YADLIY1jcOc/UjIrInmnq
pZJwFo1IjRAUsx7zm5ENWU34qEq428qO7hxUWF4Lw9tnbplbwKa4T+RA3sYgCxkL
H7PVAMjmeS4i8UBifYAYBxSY5fvlzstKFD3y4ZyrX16+kR5n7zCC8AkwuIjNO4vd
RM+Nit9UnFnajMzS8VmzRFyIpAHS4dLFpAGarnF7vBbtz/KL5uFlWEMt4etM0xIx
qGbiRShbXeTtXvfnYUchkT+jrZD/8ma7kV2gKM81FG6O2e+/RN/GQpxa9wZvKRK0
zDUTjceaWHANJ1XuQ5rY+KeZ8oWRP8iVdBN23Y+qJHUQngZOS3SFOfzxqw8bzCPC
gW2KyrSNAoUVpFt0mep1ffzey+w8KZ6BOGsljDBMWMGZEQ6sE8ZLnVDzwkKFMCtO
SjJ+iKniknrWtjhMMOK5DxPg64FRhcJQ9z7SNGmem4tnSMR0fZoufcVqvmHt1+KH
k6jqimmI7+AG+WNyI6I2zKX+6KIPDXA0vggPrgAdzkXqPvhzN1c6iAqWApnJIk9M
id68g8aUgt08sZct0N6rk5t0dwtR7PprrmYXjERQ5Jqjz5LJthzPA8RxjIWWWM4D
BsC/7FzI3MFIZhmwRxIBWguCwWCmy03UsrHceC1PUMuwFuHJa3ZwySuf0h/QpmF9
FZ1dR7ZhkHhYtttB/imvuKRLef7y2Z6i3fbcvvOtpsPhG0lYz3rxgrUKVyLzwaBQ
0QOz/OAe0f948a6rNod5weQhgNYhkSw1O+gcqcqWz3hy9aFTaGYWTopQwYVGKZSY
SLr+wS+MgOdGgJlnAV4v+FUZIWEowL0naz7GSAHGw1/q7762Bx8WMKavePE9hTHh
kzQSE8yQq1FFL7wWmMWe1NEcnYuAYaYylBw10UsCR6KbnM2RzjcQfjKCL50MBZy6
Js90of+xYpqVhMMSR8+RarzedMUTVQVIgNrHdcoYzKhth2OhhBZexdjikVWPDs59
/ItGHEi45j3yzaI6hR4DQcDF/GG+KTeEwje3w9lkog+7Dxd+Cy9kYiPJ5Uto3304
gvTMG1PkClRqm+h2V65efAzCahNLcSg4JnmyDwRZ3DkA6FJephl7vrjemm6v1Qv2
nKK9DGUnl8v2XA6tLmKXJ9W5K4efDh+C8DDJp7qkc0JKPgYflxYxtE7WLcTo4IiU
qhXMN1bBS4paBX2UKNK12ogtyXheHux9boNe2ibeNAdh92ih7wSVx4nx2ojwj600
vD+6xAmT1cqdD0WlQDhu9aeVf52aWJ1Rnn6VdY2m9wtaxxM2FXLT8Ydvyi9JDjfc
1D1BNnrLOpSVW+y8MCCe9Z8VlstbZ0NCJgX3up+TJWpkWXR9QqC57kaOx6o7boRz
EB/oeOT9+zeqOTauFaf3+VZN4qpuzb5ZrrZ9rA2MTlVEQpJgZoQPJvopVKXAExO+
8+D+s+SBd1rDU5hzbeikvM3FtXO2lT0fuZ1XnG+FXeG0SM7BDXJxU69eQj02cLsu
v57inQNOgdzPrjRZyPn0tGAiGHg7hB7tlg0XGYGZG0m/CmvHNSn1ag+oa6vk3zDn
eP33X86tFqylpk4vvfPmga26CesnbFgXQQelIvmV0H1ceMOXTDaM0szzentkrDcL
2i0Xfneac4QYo0ynOpYc0pfwJp2WmSADTshI9XnfpkPsu/I4YO/a3rS0XWJuTrpH
wJWO0rJH+vh2PgOQfbqWtAteO+h9XhP2VRkxlXx1uriUOm2/O9FVogceWVYE1dUM
TJh8ii9/tpxm0qAbJrx/ZWOlm4D275YKHzHLcbezB+z+fSLq9RnfmuC7b85W9ZEX
pLjHAJEZaelVbWW9o71q/6Cvzgi0Tv09HRFkWh29dUYamA7SE1nIFsJc09kdpZWp
PlNuq1VJyCn2KQaDDKH0wktL9yIoGINauV1e3yS0c2PGr8SpiQ/2bjvIny6J6bQZ
ktamk4Uoh1QJ2h2qtiV8kQCQ1VdBb92Dwm3QJ3quMbvNYd5CxW9vk8jClfG8rEzC
9CB2v55A4u5slrDsH1WOoePHsTI9lM7XgJS50pS2E9Y+ZZ/VThQpvOzqKHiFTkFS
fSrGDYI/4+GJgC79CGC4YjzBjQb6GFOw3wiy/pw74h2TjFbVg47ZafQsKg2/+0nr
OARrGj98FIc5qrb7RlhVK0sABquMCJDs0NA3H69UNqWGl6dnQXw4aunMruuvzNdB
h4CU6IA/ngdbzdlRp8MMuGJT3Cv6Vetd/t3PokjRWcjLAlpGtqHepC9TCyC+16ic
6f63PwqCAG5SJVUQpdXcl28vaQ0rzF5FmQqgorpxT2MbQbV2r4ICnk6td6ShosMH
HFzMxyos7iO1kCH0Jl/38E6ZdwN0ZRqG+Uscrzfbt+cF4SuGyInvcJyKDDFroXaK
DGaEJkH1HxVDZ8s3faizcsvDq1IjJctteTqg3TCRSFnM8j88S1U+roS4JwVICidB
6ll/mRzkMU9WJnJTlupRr2Vc7KCcIZu8N/vwnU0G0HGHAWwrcftlD5qpArSOr9FE
Ewg2fkgYSilhacRtYXjGk5jcvSdANTZSaPLVyuSR2STMQlXjWgqKww8artOEmOKq
yGKLSW1UP4kTZcb42DzWOCjZfUWCLsCNPmMxH4ix27SQcK1caVUuPETWEVmqsoU2
lQXWmkeJvAFqQi+x1geN8Ok+P7FFAjlv+w/xOd5EfJf4NFnxBCfHfEzXojMWlMwM
/F6ZBM4sfd8tky8vzb4HmTr3XOuCzBduElh/WRevQjc41ovfoHZfX/3WeH5LJN+V
v+vSoFWyEQ/nuquIj7sfmlnL2IitiScu7o3DqrqnOEEJijnzUN3imeN+/CPGML6X
d8TbvJQQAV4vGBIZ/e3oVt15uqejOJpRmP3cgA9hWDJO2WN/jmAZAoFE4oh25qI2
6zsZXp+oXX7rFLbKY5kACak1UEFSdfrjIeVag+agzawdKjpCvKLZnYlz7LEt6Byq
HcEg2YZ/E/hErghbBqxtUq/k9/Vawer1Vv0q/iMmzL2yacXgrSsiLr7tx1zYCi+z
lDNdxLeIMdbiQptpPBjr6IubiYMZkerBtUBRQ9H695oBx3sl+7CFokhMjYYoJZql
9DW4ruOdGIVYEwjv0n32NYCkv1OJcRNJWaK/9wGKQPbCDfm5yXy8hlTEVq/g3qWd
d5nMSU62Upg1YJbszwVyICc8p5bRFtbQz2KTAwTfI+6skQ6qNhF+UxcQQ+Ek2ESJ
sdMmPq8QNBVms4KCJSFodoYr5eAAdRfID66m2FPptYkC0g63UimzOcuMHr1mXybE
KMcfH0277GTrwI91grfwhqO9jMc9IPQrdsJv6EFC9GC7b0oyQ0U5slSzx4nNMTBs
qaHxoVqWdx0Ub6WiQg33Ce85SbVa+TMyXcx9d56TM8BkQibuTp3LbWbNWdiAWJu+
PBLqbVDboCXX49Am9h+RD2wtcJR73Fx/F9Q1ym+9iFdw7JYKQlQIAR4pN6JWChqw
stz7qnNPA9a1XT1RtJKq2g3BHUhmXf16sLFzehiLbVVQQn55iHXWX+wOPissiGiy
WPivQglNw+ZDD9Q4Tfds7rl3k3I0Cq3wkPuxQGDncf/1oLniCRUtL+AhZ0JBo9bC
Tfvs7g8ZgKr/QxRzM7IphMFHaI0rWKBybOxDb23MtpukGjQajNaQ4wSz2uYPKiNu
n61RqhXTaoASlTjyGGJg9JooDC4thACrEq/tewSXoQpCEKXHAZ0nRyAn3PyfRaAx
C9iy4tHyHHytr64Mc2Zgi6mbhCSS6NgO2k0zdJbxXQWly8PcQ9HJBHnewi36bv6c
EQvm2L0IrU0sfcf69/SpyYhf1jECaHQVJWNlVfDkffGUlIsVkugiMG7EbpoL3YPu
SD2ToL5WL47NrUsIsurlIJ3F8bo5CSHxC4WCFVf3OXNHC6Qt+o5k05g0UgAtHEIM
fM4JvL6mSJCutg2YRRIKtiUF0QxujR7HgJPy0dxGvjhWh5JS/LvzOQhEF4ssa4uT
xLlzYAc84LFeGqTGCCA92Vuq7jOKgsetSJD3WJhBOh52iEp0YLoJy7xgRjE5ETVn
BQ87+gYlqHiIUyzc8RN+sXL4wTbncsmUFHKMfVuI2mVwoSAbtynGyBzmM1XcT9R6
yLGx9sNevsSkCfJ/aN8eQb9WneHCJO9uHcWj20T8oUkAzZ+jYN+VCa8awng3P0xw
jNtzgUooURLRbkYFYEi88amRvDeO9mpNzORQ7RJPixNx1mDCYN84X6HtOZo8LFbs
rmLb3nDR1+iP+DdDzu13DGi6n9/lUK0+f1Yaw1Q1g8rXRYnD2nR+L+ewb9pRnMQQ
Rmg8A3hX/B8cI81Xmk75GeBpSQT2MblXD7Zm+pt+umorVcfIMqg5jgEy4LrwBFb4
4CjYYFkCPOz+kOYfqvDi6vOfpqo8E4AqJoGnmsUKG2L5x/mIXq8WacGtu+K4Urbk
YGtZcE0BD5UtFdmqU0B2eJ1fGJ0+3Do6ULsUXKXvE1LLpRl2mU5TU3G+4WRmTWZZ
3P4QuoXENzikPMhU9zu53XO6dik2E6XY2q0pb32cFcmUrnGygdHb/mfn5pEyC6nf
lP3EMoyBK6FPaVexxhSgeL2PKL8tvjftbm3sTifyjlKYNgTlFlfTu7BIgGoN1x6H
P17iDeQaWhwHxNw5OqYmN06iA/7LvJGzKAmSF3SAiPe5NBZkMC0BYwAZWDboUusA
hXnK8y9G5qKeqV3bZKyvXZO0T0V+uwRL7WFDHSEH3mEiyb6TyYfhFeF+CavqVqvN
Y8l6+0YASDvkMYljm6wwYbvWiAKjTPq7+L7l2nfIbPkjAzScoUwnX1eveApAe8qr
5ic1bVFCtre4+HYGD3bZn3XK3UkpAjz6sXNtrSabPcnEoQScp8O1l/CXHqjlXyDt
6ClOOSFDMgDgubm9DVWqySmWRBMNkhzGZBFQv220J0MhOXdEsWvEiUZhg58BETNh
eb/HpGJkewFIThMEs7NWqUxp5zS1flkEgNKJgMVQEwp9fwXT9aJOdXLQYJ99KTtW
GVxEGaqkrHieRuLHz943HhrLF3HD8wjp/lMeyW9dh5dvf6VYz/85YrCpk3HJaGB5
BKK2J3NrBoefHxYPErHCJL3NyYjbrT0oEhCAEZhGCHe0w9pcI5mCRmZlYfmbjpsJ
divbKJakuK8xyhfzBUAV/qYv1YJ5eOkT1zRFNVgYtytNAvIZv1BtbTw3VsFMUYbK
ATvL+eyEEr97/1nxacWwNBBDGtdX6cPKGYpDsaMDobvm05U1Lzbqf9WI7FBMV3t4
BBFA0TUa2LgLXN+Ys2WF349bjnJ8roXxWjXsl72B3fARahXkmpBFL7NhrrhLdhbj
J2uIOem7ADpiu2LnPHnTc6d65b44tgWBQja16es3KAYEFcFdVckKgI536gXqoKtu
TqbKgpu1rBTQCMsUohNxRlKGdz5N4+Ztk9uQQAxbPoXoHfttNMRdwh9vQRkZgiBZ
wJuB1Q8BtFoV9hWbaABLq4+wDuPVGi/r8KEmA8CZ6kVGCI9N7iESceALDAdVR79C
O4UYP5Jtgb53mS/2iQPj28EBTVtoP6mkNGCUQJIB6hLsOX4mko2kGrZUe47V/18i
181WiCTrAWHSv7jBuZqXLkXGXXe5/Dl9i7farWcQrH64apym0g1nq+/B90O42b5V
F9wk9ghNVSgirV74QAOCZBwKuOfoeBXeqDlRCqvzKoJYLbuekjN4AticgtO+I9Ph
z9t2iw6r3LXvHN3srVaHaKQ2M1zHd9fiWA0l7aqWxcx3/QCzU0/mafl6ecimrDIp
TVf/j8mhmAD6ZxlTFZNTdGGuONy7UbQBosSBSh7yDEGpGN5Rd17TN+b8YhbnF08G
9qL+i2j1O0sBs92maIODkLRbk7oUjcLjC3cN1hqW3e2zMWHjJNIYroPg6YShDh/Z
GpOfJ62vtnSU2r7Aq2FjvGJk27LHntfdikNDCjTdjyCbnMK4peF1UA5fWSp2t4u4
RMULRk7N17aMQ6y6Yads13JvJnyrNEslPSRzSM2D0XBzIpDQ1Gls/5L/SqLvGgQ8
arlGxGQS5tIPWf/8ZH9L8qeoBr/xkLhIWy9Jud6fk+RI9lTKqIwD9u7IY0ar2iCZ
XtMHohOjCwBK3nJb3ZaraoQQoT7pl4MgTnIZZTMqOmUZYseQ5nxHpSbWCeGab4sZ
Sj4jcVk/w4R5LTjAMWsjO0vYHA43YAFWHOG1F6A+emi1O5pPhvmOwDytXx3V79PJ
/fSjtLXkCz1lwszUzEHjmuaObv5bsNb7hrIsBUAAfcsdVYvSSISCbE7wPathHvuz
tawi1krzKpt+IUOOuVnlUWeSoNghAIBJkbSy7/XsO35iwI46cAVjQEZMcsjvt8bL
tiahSwUxgswGYHi1goNYaleQrJANJCO1KIvBMOF2B6TD8puD3M0dv/yQ+s+TXOrh
sKPDkQLuAKfrnXAOTW+HZSFGX63WkVEN92w1YiiewAN5QK+vzNKxam2t+RxYRSf5
OlqMfIPhf5iJznimg97bUZ4w2iMmyUE2XdVcLkwRpdh6EuxayNZ99ob5J2KbJ0tl
0t2BH/ks4AyaM4YsX9p84FyLM16MvNOQW3TM1+yS0+u0LcqhqzgbOS/lEeVvsKeZ
pHQYLyQv49mFQ7wfperhOXnDCEkx9nY7XEhco6AqVllX5TA1ma2S2xM3LLtzU3RZ
4HjAFGvA5nRQChlxyG4BXMyZphtzwCnMmNG+Bq37fea4zyy+I8Bs6h9aUK8p6NhI
lrOAAdkb3lh+ID7KuN9S4y0TjeQ5osh8vXig+m6a0ym2/u92dIYKx1uwUqw7bwu5
64+8iaR4QYUDSPJSPus+qCxbIAdlp8vlZGIOw4I08cmu0a+ky+7XLADi6GXZorIx
pfNDYoFx1x5mZPatx3B3b4v0j4Z9WaQut7nGWQGPrXpPQLd2K3XFI0YPD3si8ixK
NmbeeLtg9dC+KeOhiDAcQXeKorcA6ieQSShdoxrnPMZkF3yFvxWkhDmBZ6nP2gqX
YehgfWBrEcYRjU1jt+KAVjm6XqzCQWFspWlaagNoMqdHSicQE6E66xOq3s4yIVH+
75GPZ36YZhJTpy3v13qNO7z6fVouCjyJpT755lzq6Ekdr8L3AVoQjdiN6UftaCjH
AShCFjMpKSWU/DyrhrmzPB8iTnuq1M46z9dv6D7tjiDfwsNlIYHhNtqJZZusKdl7
yj2TrQ80YZ70QLfRnpcwI+Tdf9krT+OmT+UeaTuZoZwnvjDehq/d2wGaL2DgTIrQ
ru+r7yDHDJW/7v26rveFmX4UseSkKxA1yIKt6pZn+uQ8A+hCduJckp2H2Rm3mFEG
eCXvndwAyCRPUhBb3cj2Om+go4ljplS2eIPM47Kq73ceh9WfwS6GlZULNA73mXre
Rp/2TO5k/YEz/hWZa4wveaP3ny1uNyWVadv3oxXshlPy+g4RIFdox0OOlPZ4HWGM
gI86NYhPkOZmMe/L25z6nU0KfQtcQBQUyFQH+pg8G9RcnYcHTAEjdVZ9nb9n2aP/
DPjDFmi0+QxwxZhlWGj4fExovF7g2C+Gd3PbNkWKYg2mn/hEkSWCTdjTd2kdC/rg
3kd4wpK4M/Q4CuH7rSAi5ky058nWs9FOWYqLJ625ePUWd2DkG1mATdRpUpQOI5/P
JCsRGDR0Skf4R3WbvFXVIdpdbvuB3f9JbDFBnqwzkbloJyBzZCB/sASTus8M7Fwc
OAR128BsH8HO+UVkRJshS9NciBbvIZxHr9ZA/ZECVWrLEPC6gkGVSeig/EyFwSZR
pXt4PrcVwUU1j36g+Rc8kavjD7W6Dp7qh2zbw2T8Iq+UjZaqXIWce1zL++acdNmM
dUAOqjS3OLH4ie/CyCzu2mOLFwB3H5Uc6CCsF9L3U428jSTkBJFg4b9nwWbLBuSH
M+Waah7pODjvVdAponhGPlypvOAsv+gsyjXShdNxHho5upnerox8DMyf8jBKgADk
u2B8r7b+12Ljah5lr6HeBMUhzzMq2iERi+JH5NZF99bVL7/E48Jq3XZDxdFJCyqh
MVWDAGy44g3nWjSIkHRW30tly5igBVJEg7Kfwwbnpj9wYKK4VmsifaGjHGWCBD1h
BHnZZ3XvD3gcx+ZdsnXEuHqdV83OQI0EhlpWUHCmaF/XAHrfbHkb7EAGq5xJDOMx
aEo71M8HpAieu0yI4qcNi6Tr2+JH09xiTWoHcDajRbFowdqZLIfqWMHt1Gwe/lxH
i+40oiG9b2UTYFNIwgBwXBWnUyFhouPmgZ+2gD4KyktkVAoBdVdZjeB2F/b6ikTL
kI/yg6iC0PpeeTAnXllv7QGZxxH5nIfDOvwsw6ucj4dR3VIh0z8lTGhtKkqTt8bu
ufXs3YRifiJlvgZBQUbfKsio/+YnWrOd0d51KQi4ra0uQNpOgrMMxyW7Jp4vfitZ
RUT6hjvXkzC3Gu6CzvJ7rA5uFKMTNaMdUDnMl8Yet/Nv6UyP6RYVFfZJdtgSxPiM
49N8WSYmj8Yp6NxYwzcLTld/qgEkPXXUdPBFL6gAjrvh+5PhHeT3sx+6kHK6jQiz
pQWpGvzMwMgiV7BBlCBpcf/IjSr5/5PA76b2iikDHs9paDpWqmHAO6dZ5Ekmq33+
SMJYv/Oo0mxA+w5jrZYyYop7EEZTxLfBU8U+kkz81Qmgz519ZBTXsSx58evhVWD6
jBNReBpFZCL5Obn+N+oXvsF+udCoLzDad4Vp2iJWC0kIXhGS8HlGc4YOWOqDdeoi
JXmvt9EIGVDpJ1j6ovy4tqYGFpncaNENQWVvrfmb17pctd5SLBZccOnlmxVUHnj6
EHRpskFGpKiDghatGu+CyUfEhoezeGB0LEmO2ylhZXTAfVomhY5v17gUORNDtfgN
EKD255CeI3zeuO8heMehwmaqU4bczmiSCP86w6l9I8TlQAFkOdR7DYOLQY7Bvx7y
rRgxHpwbjp2HwrxFhqPg6+g1IIRlNGKAaZahWWqm51JkWR2Lkrc9iLqcN12pYlE3
E7suOG9aCCVd7gJPU4bwz61IZARbUC4wpdypPqNXEFVtRqfsGFNLGramr3+oGyu5
vK76dDtVFrEe6iFT56QEW7r4lgWOo+wJw7+oR/5R/Z6vVgqRPOR5cBYDhEmDzeyp
qyLu/aHpryH1xF7uqeQnbGUIREmJK5c8uXi6NyDYdjQ/aDoHrfP1QxPsIdnJcQNj
LB+mro6GBLrRGS3tKeN0ilXbRqePcFRi/VmoOPlnzwLZKtzKJrjO28UBnozhWsML
3whyIIFDQRVMZHtDDlLA7aeE0l92mGSbZ7nhAXMgXR1DH6pGJiJhE21i45KR93Zc
RIoqP8EIKvWRgnakpqh/Jo17K2RcPTI1RZgGUdhuJArAOzmEgzTAzh7aHX6dtOwm
H/08GdC6n/0/ZSRrnsspEVSrYfyFokaksAzEykr2SPKaOU9dMZ5v7hAYNEY0hZVn
rxTg2VAmOQMomi8m5WE7OMT/ZqOigjOYuFoQ8aofq7dKY6p0t9zKCe2Mleq2CrAG
p97Uwy9DK/K+lKrXgAuM7Rw3KreOkXNxJLiH7cE1jrhptGsk7lSzfAv31PlqH0GM
2ajuXGyeYr71dZ+LCO6+preYoBtqISu2UH7QXf0kwvbQ8ps3E4d+a7lA4lQFOaZp
tABT4V7faC4jxr+zt+yIITuBEsq3UjF9pHkzuIOq09qLpyuXla5+KaLFw7BHOCQV
W6IFnjaDtjFs3JTyFgpCQQBRR0yN15FFQYW2XD9USiepMnriEYs4b/g5CH2FUZTw
+vsslI5koEBhc76cuI9iH7pNqcs7g9W1+mt7itux7gDYpTmH1yHWa1caHh2ipO69
H1RPspwCPtVW//ug+dckzVLiiB1/lBL+GRGjFF/5rSsQHlBEpwXx2iLbSQWQYGBG
roBzrwNFDAHJy9mHQ5QrF+3g0D436UhS9+zW2R0m6BeW0bSRGTI2k5QEZzn8FVWe
qib7ZmYFg3MxFYATcmgQPRTROuSU8BBG52GmGLZ0VveDAFxaz5ZM1ywyTzGpCwdX
dRTp6DJO0T6uXcnw4+4VNq9EMQQyd+LE/Dm3rnbJVpvs6Qj8mma49gVz2EvhpJdF
yyNs5cDR4zA4vsynSF4c6qgtrKKPKKrh5drt6BB4XUads0nOzuV1odx5G0tTpZDV
Cy/+tcXlpPSw3OkyKmVN5rdW5AJgDIcvfBSbEq6H84lCAsBOJa1Yje+i6xe4Rs3k
iWPhChA+om+MCz1hDMmvNNQtW16dNklUSLZ5mzPBlxaadfzdbx4siVv3QBgxbANT
jttSU6rDkNxC+vEFERUlclW80ZwzXV5Znmfy9ZBa6bQANBIC37OTPwTvDJniRX2t
xfk1Jy+XXWOCuIXNSCmlAo2NfAn+QWdlEIhuOuwnCPrhK+IvkzblRDlXZOkg8/IN
BcJuH75QKYfcxwRYeSOjzCxZd9mes5lt7mzzXIdcnSMaGFhgIvWKcoVFh2+pc3Ou
OK1sL2VjTmJVPbjEAcCbTMvmdHGINpYTW/xoAR3ZQUueXIG7SopREHV+rqiUvlcX
0ufkHJpMomHbHXIUyjyPokrV+bAEQsQ6xgl48zTbDqDUm+WQjt/0cSEwxxeOKud9
SSoA+u7/7R6rsl3yT2rZqVKtdZ//etDBxj0F6P8OAollSfvNv5sbZE72in3AQ2Ai
LzK7Kwqq3aO9LE7G093bJVZKhbeJEHgI92titDt8TkhTFm0tYZoDZOzQUqp4gFwM
1aMeR5cdNdaVkMbOZ5ksYGRxRufaiNig3vT5QFSCmMKfUVsYB3wYkseLPEbFNxCQ
im+cAiIBiGD6+3EPQbJFvt4rJateKJX76NnroZSuIYtnQpiNjrIjnLIvI/HakWL0
1uvJLayvx4fZZs48vaEvYTDbCLp5ih9OWOUG2KCagaZ36w3oD6MkwwZRYb6H4MuN
JSQqe2gUKAAIIoAfgjE82XHMRQdyuVyNGlEMhj6uaqF4Xky8Z7HJqT9Oddj9svC/
+ELoJuTBo8n0ZXSoduEeZ0VO6yHokufYcmj/9LulfuoYYmoTkbxeoKHoAFjfdsCT
lOJOg6Jv3d5xLX1gvNHW+6s1KV3ayimOr1iZ/H/WntBgZ93HOb1WHub6NEi57Grd
GhpaSaKfoFmN5ThvrUkdxMxJgcKWlZrTHxN8x37IVegWB8XG5QkdrvRfLrLJBgxt
1yedREnFiF6Pb0eAPjMekw+A1BkgeXetxW8oK/s3CP5s/LvKXRWusveI5vy/IXTL
GfMGz+yV2ifVz46pJbdAvbuFDgSAEH0rGN2K1ecgO5dN+eOyohDIlWucKOMIVx2g
AMuG4lMwG9ubXc6wY0giui+NAfOovN/QpLF3V9AIKJKPPmjmut0L69lHPGTHkNHB
No56MjAbh4sRWybND4ANI6SHge/YxYTl5hLEswiWuzIF+90q05jJmsTUFX8Bm9AA
oKj+kmx8IQMdLWVwdQlujDtauiPtdbWIiME2phPaS5vBWbAyUOB1peLiBtJuFh8B
1Nj6ixo4xHT3+yYvhpFR2kz1Z7eMGHOx2ezzeaIkbyaijTSxBd8qllwqSiP61shy
DfKR1MTxYaBGPJCDtouj3XxWEp8gp1NX9Le9tcpAeS1tjM+wChzbmyuMBwLahS1P
jK388v3iKld/Ohs36P/xdxQpIJlUsOnzT+7sshDTzpgo6a6v3e/ceQZrcD4ZZZfo
7wT9mvvg+8kuwRUBqx+3PLxrYHr4TfdUJx9+QdbHLdrNphJnjO+HYRClxvrYRcf2
/S7nSL9e5u8noJ4obHpGQwF1JwExuyPv2urCfll49FxzGVQ7WeRq7hoeMiCADmEP
HShpWOfQd8QQazU3h/pyD7dnxHrhYlQ92qytJnRX6PNd8xYCoyImTClXwbf+KTXv
nJ/MsqHYBcTyqxc5U1Vp8tGdHmZOj6rScAeZLmNtMKrliIrmd5ceO3FfTVaqyEwq
0bc2AE6BoxIc9zbT4N/fJUkTZ8jSdqNmDw1Eges+ZLURJfGVS7AogwqzaxRnrfKg
UBNySox8ZxUl40s8LeezPfVD+z1Drlr5nrCzmJFfmsmkMIP+k5sLuofybSv2dWw0
3dmA7xNRG/5LFtPqI3HCVuaZOmmgm3vv/Ty/d/FHjvqTqSC/1oUs+8I4h5yJI0V8
qbH+miDVkPKxEj1VOiWlJhNTGP7aeKlAHBijVzpd1+HTr7e58OnxZS49ABFMq2aO
1D87lAglrgk/lrBiw5ZPj8XP825l1Qz7SLCVoADx6/7cOuKDGpXxsNbvmK3Qnm23
TkUjO8e/mFpsSo2JCkQRYKdEarnE9GOwkte+1FDeJLJFeOdNPFLFKf2ECd5ttyaZ
KRoNRs5vicmU7vpKKtRXn1+kQ+1nA7KFAyTvn79MpKjlyc6PYb2XEXRJQNc1jHy/
vOPLalM3A/Rv37rU9Xyg8M8k0WQdXz9QWyTdtfmjsP4PjcEHl51RSNfarAMa1tjY
W6ar3XfHI3bdAZFAj+4fcS2fv3D1ZAQwfN/XV/hXqPuSIdxoxP26VHSrJ4vghzvz
0KUrythS5Q1w77uLSPTpOlkaDQd+X/oTcpjV8dPJgz/OioAbS7wSqqvYcJWwxNSb
N19ghnxZJsb10zQEc6JWh5NWkCLc0H+Wf+8fmkZ1nHGQle+ZB1G5I5GwflkxaJ5H
c6sG5mZj2ptpbqFbSZcVPwFVfLog1MMrmJzYy2sbQ1gQ+2vFRS1wlt1GUUSqR1/M
A84Daw4U34kNVnDg9R8eOxa0Q3CB6JsQUbM9CUG31M/DHvCj/bSpaTTYYWHISv51
2Vusc5zfbIXGpcl8luxVTIrbdlmCHDwdvh+iEFc+r2i6zhnMtaNve0XWJyf+7wPi
DI28hLLGlY5eCTIR2tyrG3IkbaAykbJ8/4mTWTp0pNuQ8RivazQ2Iuw2oqzIax//
QWzuBzgVuCGDxCfLnLO//J84r8D4Gffa/8F/wquR2pxn02pbpeh0T7efI3bzQJE0
/VMfrMvb4AZZus5r0QeLOfzkjAeJroDg6KDhQX4/wLWV5Sow9lOPfYPy2aCPuRX4
LuCrCbwYkjyfz2eJ3IpjnuMUJXnfZ3hr8X5cMU40G0EI/5KR0h5YoGuit6x7oeTL
whxcMnqAA9H2P21HfzxoXvgonUwVn1n/GwNncizHOQEYGUuRnH8rDncqPwll2eoX
UjlogQumg5SFPnZEljKWSGvgQcFAInHmWmXMBLqpBRPzFyPIFbot/VscTyihk7vZ
lJ9s/Ju4fv3zxrz6/oCOEXCwZWJNRm71ZfeEbtg46G/Sae0SJuG33IMs2hcNqj5k
LUqHdOhkuF/YOYyUiBZfGs/9WZh8/ayoo7ceJLdFslqipDyU5/giPBig66rwe0Fi
IxmV0FdVsIzSp0uQ72ufWZu9toeh/nk/0oCUcFIKnAsYIDsCpheBavHqP+aAOF2e
3BYrH6LNEfexQAgpDFmNeq1PHxSQESFSyOr5YQSLN93x2uB6530IuH+Im0uq8PCM
RivZbmjbgDn1OedtnIoxePCGonKtdz+lRFKAPZHnXAx1msRVCXVVyrY8SJITAVwk
/+hrfus9TTj9n3xAbdn6tve+44Qfo1BAdbVlN3tXoMLh0/81WTqZq/h/ozOsYI8Y
GxW3NEleZoM0pKV8CTC0aQJE5NkjYlbI+IN3gyOv4X6jgCcsVzUXuHqFo09VBJut
1vbuJBcTATgkod0OpRV6Ol0jeSjU2P/ecdC8pujZimdkV39vG0nlEB9F8Evt8wat
FmeSqdOCaF3Qk+ZwtRjEsRJzyxg4TqND18zCRyc/VOsCRpSFh8V71r38R8NTYB14
ol2zsviArCGcdA78jFYpfXNFB79pzVX1x7vhYNDfqtf1JfBusmLR3MXN3Kup5aR2
PJKkdocfen1wcklvZCkqHccsdqdSKk8HUAitlmPwyw3FjGLOsSQ4s336zbGfF4Oo
uKSM89uq/yeBxj03ap2uM9avEqeY2e4G/QxEcQ7i/0rLB3go2oBKRertJwyjYGWj
QP8ycFQd6mgM8bKgxiqyc/rke9YTumEIYRS+3vzUEXrrBL7Qh0KwPLU+uzNZTfvf
+rfvp0ErIfAyX1+rockjM45QV1p0M23Irjjf9+UpljijJlKyFbXUIYiivVZI/Paf
G/LReKqEbd6EG6oGdKmVnqPV5dElAUhXKK9yY8lu8v5WfQlRKotJKkme5xcKo/R4
Id11rqkrgEmJZ6sD7Xc+RBN4Myp4dmrUfkz0RDrun806E7fP+Gw6tgyHJnpfkZbm
cgfXzbGMk1E72IMWlXeQUCcLE5220QDX03KygQhV0WKWhVObgp8DkrmzkUhgX3hm
PME5IvE3Thk0DiyprTK9xB4007SpoIWvrw5ygyzD+Lfv3tlrI+OSxcBnxhpKEg+L
J/px+zQ66CSK6ZpGf5jzk7l8DXZXvL5xXHTHCkyer2UiQvQLptpQliT+QdSSmnVp
qCMPUygjqzIBOk8V+h5uwIo4gNH5pGzT/tMPn7QmqSfRjsG6Z9jqvr3NT0RPbo11
KzpvuRuN8rC6il/9XRVzdiWP3k6ZmKpmpALdHRsCQrBkfG7eA3OJ3YaYKxL8Rwja
30lMqV9DXVRttDs7R8hE3aFMUSCIgZ82gwFW0XLOk9CWnmjChNS3wntM/VxWpmjT
ChxmkxM7v8sG4UOYu/+ZH24EXDp2RyzH4+kjfcMNhXHxxlfXBCtC7JmIp+h5MnPX
R9MwGyahmROu8kZ9OG1hH6ynzRGUk4jGBNTYaq6wKI12cFmhZiZU2Q6cTlCoNZe8
cuVHRGFfvioqmC2TjbUDKui9Uuf5uYynbYxn+BajlTbr271pGRukW6HbjVxACNJA
K/uhDCRUdsWv7zArn82QwBeHJIr/2ll7an4wf/wq+SGqbiviprBymKmVRmmhJ5hc
ApZiafveBDC+pe/NSIzedu395KD7o4SMZtRmpkE8JSUCdDuabTmrEVLghYnU6jOA
Dp4CtVgTzHO6V2UuxiJJn8b1wVHrAnE03A+I03u4ot43SW7gPwFwAOlA+suT2OjH
YD5rCwk9WUSVakVT7HJYpJyF+ICJI6sKuUAf4maA9bjEWLZaVv7rq1GrQe1IyQrO
ez+q5KX9ip8KlCw+hQ1wZQLvg7aLRXsmEgxtKDH9/8MAx3AdgIW6I++2pAL/qas9
ldx4ujUlQqGrzKLbyaZBHK1wUQcgokSJYDFJANEDhXrGG0FADCNCgvedSWmKoYnb
DUxMG+WDKY4K2Q1ebSKigkupoSBpA0QYX7xoGkHboBJ78eVjUuWieazqjais5soL
iZeTJNTm7oScvK6xyGEfRzM38HmjvH7P/w+jY4TU5+X7ILS3d9ES+zU8CeKzwoig
QU28YaKZmzuA7wJLkJALTLa6GPf3X8ncHyjxHd6U2n+gwzSX/17fU7BBe04aGoDu
ez9FS4ZmeFumEfEVdVCMmij8NHfNY3rmD0OfRGFSk3P48KB/Y4AbIHozke50IoxM
/SoPsbM3D2rlo5tefn5oK+/WFJt/PHc0e+yfPxhsuPBPBRm1IjARBZ6Hx6yDo8i7
tBCwM8+iDc3p1ntHwiTcbyyCNq9BMWs38506gtPdq5Gn9A9TJ7Nj9HAZwNv7Nugg
OPGWaWOJlfsEzQiaRhSRzPGsAmzq9wWYfBKUJqe8lBcfxNG42tbb/AAEZxdkd2fT
AUR36D8l039uOIwuWJD46OBgIFtiXRD4QhChgqbzkojJMZqoLjDbLajrPpB/YJJy
F7WcFNufk6UKw0Ox5mZkPnHxgwvYVMe0kTgD4KrY4yMvfgFCZqEmGvgouA81UHdo
IQJ8gfFPspoAEPMdYR4fKCdyxARpAeBK0qSvHzK/bKFAzR54mZewEuDQD00PuKkP
xs/Xb09M6lzDaxSKiPHSSoNRo8PocbB5DNMi+9e4L19SkI0YXg4R229xs9g8EKJW
xDmJ+2g3uxZ/smvNcClU4Oe0HsCyWbHBAyjXXNImaXfHhjbRgUiMZONAAyU1V/9p
Qb48RfpK+IctjviPb7CgF1ChG2TCKkzViokD1+YOyxN5BWar7u6j4QNfYbGWd0f2
QbZunaVr/3Be1OO86rTkR2VC+kgkOdj6kYBdcKVzKxyl4FT0SN3DDamolyCsRxJ0
IOJomSaiRBBYEIZdXQ2cKeE1Ll5j63XqxVuBWfqrDx1O5VITri2INmkJujCCLYyv
x95tF0UYwXgxhqVBathSzE2wbVDpWCt81RWIW2vfLGVuZQEecBFWrZLwxJDRvYHk
O6caIecR5LJkBlqDMehLBtnVs1Pg+g9OLme25YxDWBouKpH2h5C8ydPfewU80oLp
a5WxgS3tL1Kb3WSGXhRC6sqDLi51RiRtHvbomi4T2WD5Dpy3K+hK+UPPMbjvpYGF
xA+dHTfI6dZSUcN4Lmkcas6zzKLldCzWLHrXcfahrEDhEPBkgI3tXEtEbh9ldxMu
vU3LdwE++VwXbeMkLM05NaAzeMGE5HfFmtbzrlGp7Ubq4zKwgN2smOnrIaG6BG7r
8W/xkaWB5HunT+hi13p6Z9UnSJuUIMZMn7yx0VZ8DugxU59M1/pdWJFLWAkGHh2P
gcHOzngoNptd6Epane1haguNJRAW36Qz+tUc3+S5zaaqWJck3b8C251ug1rLD80b
khjlqBijqYZh+Z65S8Yvj0irH3IC+mfQdd+WZzMvQqxMNWhP8c5JWq55BMHpUut9
5OFPbN2+VSnUCEckT4dyBpNTyHX7YqksSo/MgQTwSVlyTRKgPNqRieh5xo/EbfxK
HajMU3MCMCy9M/cAZa+RJCcajrQQlRfmd+g02znX6/HNisefQbvZ4BEiQD3t8I1G
pbtRdXtdmfM/s37T42w8j1egiYAShIBl9VpagT5ySB2kgohOGf5PF1E+GfxPvBy/
V3ICUGZlEnJpXJ+x6lGtUx9feN773BCZhEK2MMhBobFoWGSIARcBxRdOIKt+JkRP
ThohkV+YDmV3oPycedyYCmMsVXd6g4kpWm67WoOJEpskv2leGbPpOru55xd1klzX
XzGoJeEZWO04S6ORXmheMPjMF+E5JvKphnQrRpCwPV0vTPgoZMMPVlLUjpNwYWFw
kDDHdq6bjZC+CNyD9y5ghKe4qKopRbcN341nRDM6MZAh2+L+RkxIIlm7Zz+A5No9
9bCZswDp5826BqF4hxu5n6WTS9VppH4ncMSS/XqqGPy4nq/HgDvqkfgKsmF8KQz1
VSWfZaWDYo3NNO/3ZUR1t2pilBQDNiavCB2Elq8cjTh9QPA2/jq8qY7Ls8T3ffZq
/IcVJc/BtL4jS1K+vEG7tiVC1FoSnPjAMI4PLWLLDtfjZ7VOxxnLdcm6c02Dz9j6
YkNbhYRstPvKmRio8Sjk8sVwn2czC83v0jXUhnVodRo3xfYujWROuii8PzxTQpSX
ckuG43IK26br8PYy2/Oqcs74nepr52hQyAE3Ad+xHqGmau0VkuyRDFwY+ShsPD+K
fZXEmO//r/99TFGtcDl+EWE7AnH25vLag0Y6JpFk14wXEeAbQ8Pi3kAnLf+toph2
ImZ+qdo8O18C0cfGY0yNEnDZq5KEzYxqCpM+6xrKsp7Wwu4HsXORoUz1c8McB6Hm
9RIrSyiiHIq+EhJ0BB2Gc2+4TYOwT1ir/YzL+HIX3tsA0buHdEdQqa068wGA3k1M
emND2Avo7xJ2ulpHPo15o141mFfXricEPv+U02fQLWvx0l7sTegwr53hdjr7whNn
5xSNI1q3ebmBhIBoJWr044XmxP6aEJDaE+KuvEI2sMLFTrLNlJLTbej0eWLd0YzO
SaZT+CxgaN6caK3ATcI+bOT0Hk/0toswgKk3p29YxmfEVEL18NGP5gQpVQ5eYbMu
OY/D7YyBY10jXSzZooEK/FpzEdrlbuN1xNGIYTzexmzvmcqyBnMQF1kVpVxl6sNu
gtwlWPoS2XE2Q97TiSkPhVm2Wnez+0rNdpXxnAHoHelKQh0VboNTWmxp5piuzktW
DwIqVMfM5s0vu5wu8bSoXHvNpOqVhtoY9sdEsTqbqUevMcOVv8NVqOr+WK3DSAd2
nMzqOqWqojtggFDMbfSWiGimro5z6MTClalXMQgH/1AzxQU2nPMV46uvpeYkTR8H
ZKI6zSns06GssigKP24KXPdvsGPPmMBEYItSC2wcOgus13Yy3yY57tdSg5ykp2pf
JQM+EDMxGGRwQKx2Jz8DYn2VWJMdzktliPk4thMGBMribmhC/maTsIgaIPdt4WKy
4KnCq2FR+QpG8OCHHlUfFPoNnWUifEKwQlLRanxwZf+1AAy7Rklqv3WuBBEOA5K/
V0KCo4xVGCYj+QWm79SgsBjpukyqh5iPP8P/IVX8RwN5boN9Hbr44WLTY7qTkM4L
JxW0s00VcF1aXVkZTnttx7ngicnhyIYYKlxNJ/UmKW0WCSJVJ/BEtL60e/g0BvJO
LINaUmbHI1m6jR2HRl4VwoM/AG+IjuTYTN2ZidANYF+GgtW/Wbl6qWd51ZYPsWb/
Y7Ywu75p7ZMz55S8SO+ilXE+yJg7UtY30nFQGhXYo5m+8Ia0KgfIhPiG3qflS8VN
3cAafeUkJ+GKq0gqAvI1mz5/UfbAmFvBgGolYtDd3NBzMod6D8hJXYxuvgNRjcQx
+o3OCHymerFa+fPiyHlSSnQuL4THqfmOTmW0uPvQxO8HG41dTfUOu1fBhXm2IXNp
TTfdpt2fm60AMURDULFxJML6OlGKPAbbNxNs0R5+Uk4Ow0CzTy/aeIxU8ek5nxHk
fhZXDhnCuxvATtuiQ6op70Ih7UAePcFn+/eqVO/GrT7S1HJku8RDA7rKwbzWINgW
MNVVzqf8yH/ZwnjQuSxxcdIe1kYCRnwBzlSCmAZsWAf9MSILLutHUUOB68HBsnOD
0Uafc0+VrHiDwcfRH3yckmMY/zHlZ/G4H7a/kaZicmVnRRu7YIWHCcO4Jd0v4oOW
+AIoqVhmUhRhKFXDl2dWCg95EQhaXoehe1vUQUOAwulbLFTeU5jcrDOVcySPpd8G
nN6k0DONoaS1T6CMeG+sq6l+OSQupM8VIFR/uT8UaqcOgXpvns32fZjy93Kql5Zl
3zX/YYyKibw9guIh01hW+4GxqKqSCwZKvDKzUOVSVWqLA/cCw2C6lz7wzyUq+vCJ
dB/irf+n/zyXGcbwh5fMdwVDc2JigC0zQb8kmyGC6RMIxdkqTYcWGOLcaAZD/Ref
liQZ2IzrI1ZhLTNPZQgjI0xkr2R4mAvLoY1xe741Ic0gk/8csXB0JJeTWALoCvfO
Zg1+QX08a7T9V27AQsBhL+0N6/P3LfZI/O3xgY75ejQHvrECBvPYR6TBvUyDQWGe
Jj1OkP86cu9WY5SUwv3ya3eSARb0J9r68AW4p68i8HBhUdZDoTqvciawkus8lFm1
DrZwftEibMcRG8u2x3MLzU07XcF39FO/PN1Nh8M7HvLjxE8iySEmmNY7o1ylTp2c
HGwhmo1vSPwV1BfKAm0XdxR/yOZ7xL+82xeQDgDuEslWKZoA3C6qqlKUJt3ENABg
+sNTuUt1i41SCTQdZUXbIchhpzV9WRc7hJ64IgJsW32Y2Gu+ebMYK3uX4SUstzvP
esvz/JIe5icFWYX9jvfscpBuNWo2d7ClbLenpBnIfbHlqD/T0bIgNJ7vU2n6Ob5I
MximVwztaWaBpDWmzT1SutxijxliSTH16XS2fSHWXACF0XWz/tIEuVPW0qo8nzsK
2drgI92YcxaqoKBYMn1u4dpBQ8zaBUM/h175S1xyri0LFufUdrRIwG39k5YL+G4y
hqsfIrv7wtkuRTqa3872HQGQH9BTZEsfreKBl1Ym9aAw5as5u2r7wKLTQbA4AZjX
BDZvuVIGqJ+5AZv/zigAm23PbZ5n9AgvrHrstfx2WA+nAEdFCl2bb3Ggz1Ts0e27
ddNJ8Bo/wbt0G6gKsr2mBnM0BgY5BKRxnkvEUTPq4Uk1RAW8e1vwgbg13tEFP8m0
Cn+gyoDzknEe27yGscNZN8u7nTSPwk6JDy+k0FbUHCuV6X9mHrJw+ZvzW8rVZ+0L
ekiNLxcrLHex3eRqybzh9bAb49YS3niugc/ISviv+xjfPhYwaXKbNfq3j8zHhyE3
jo43JgnITKMbFoBPsL1ljNiUBWYVNk3hjFpkTDut5dBjTwEhqhxPXjyUMcu/8xcq
s2AdrLYQU8LNwFDa54ZD22JoqFcSkzS3yvUYVW/d99dhwlfYFgbg0W2Ywf2EQzLC
d2eD8CLwbtlSmdxoy31fu4t2eZYV3GocjstZNv0xYuybaV1s7ldeyyfafSL5AGLI
tAHIiWGPw8fQ629dkphB5jr8feLLaptA6yOQO79FBt1Z1VeoZos+4LMvbpsKq8F6
x769JULRHAeKICD0mkQjd9CoZa/Yfz5XIaI7nCSZDsoPsOwkMNqx9U13b0ZwvAeg
WrcSdDlHqe9KCCn/k8g6ilcheAd1941l7tKAjwUerb7qOay6AhYvgd3akHGxVkTW
QdMtp4cZaPg97xB8bwEj6SP3iB7oBjIY2rlPy4MXr1mjtxsF+4UINBtQwoW2h38w
4G+5bUOKpw67RhygmFXnkub2oOzJyvqMohVhAxyJJM/1zsbUEQ9x7X8epgKbbzqw
u+fGgroebaN+5XfiRyWN0IXzkOJDaWY0zliWFha4+69abE7p/QQxyoGRYNZ5CRnq
qyfwUSScDwCMcvL/w6kV7IcrD7l5LL3RvMMe6a/eDrdI7B/q4LHndyCLJFGPwQVR
OcU2fPk6tTAyPOtZelDj6kh/St5/by4hYiXNL9LDiqwJimIZALHKNjhCAmbRLslt
Nkv2EfnsTngaHT4MxgJvo2IJdkmK3kr+D98iuyMOr6MH3r0vHsSoxUAbzdf33G7H
c60aUaSUYhpQ/WilHw/BlQ==
--pragma protect end_data_block
--pragma protect digest_block
jGH+NpgB4ciBGq5l8xGoJU7RQIc=
--pragma protect end_digest_block
--pragma protect end_protected
