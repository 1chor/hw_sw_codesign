-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
uFwlHSheMk6ltmM5r7c9CzPAzuUHzI9tzJ0b5ZVXaqe7OP1QOfNRGlTo+B/vYTfP
Or33cSFbOEM5YGPQSDA2U7+AeSbfN7DqFVGabKe3dFcrrap6cCghLprWARf7Cm1B
ro+6WQX1ZnUk9B8dHcrEoJThj8Nl202gtL5aGfpakm/V2s4Cw//7aw==
--pragma protect end_key_block
--pragma protect digest_block
WwnrUPneWV/gXmtKQP4MaR7xpFs=
--pragma protect end_digest_block
--pragma protect data_block
OYDiLJuXbwcRySuiVAua/Xp+BwjJ/PuhHl/8UKfXM9nJhX59BSiNM+hgOHUwxqi0
vcDula6OaOXIhQDT9smKocorB+OpGcsrG1uegeoabUNeAEsyYfoJmguqA2Xh2HzP
Ou9h2/mnzZT5lqm8wL2CZCAculJspdmLDpuWBAfh2peo+93fINX44RgmZ/TeoI46
BfbcO7uZnV80nJLN1SIK+ufa5HKAUlJNjevh0PDsmBt0c4Aad9TFiy3/pLj53LVQ
fCmg3ECZrIDJ3uLZMFklMEl7syeFJ+CvnxTan9MbmuuHMljXpvsgcpEgnGq4siIz
Diq9EBgJ/d0off2XsYWOkesLQR1p5vfFXuY4/j2/rM9fhUPUubSmrLpiOZ1JEt2G
EVbIYH71ktEXflQlMRXrV3DL5vy01OkAXKsWlyl10hdMJC97K3yIS/wTjScRCyGD
MmVa07XShYyqynd+cIOMEDP5KdLMUrx2VrIUfiF9s6UJ0wA99aUbZOSys3U3Ldkb
XQYtwyLJOg52BEdH5hARCpGw0Y3SsZShn7dC4Ke1ZHXd7StxLphhiwzhhfXBavO+
x30IvvXyhoNdqoD5G52Eky+YHxBoJrBUXhQksdqZifUVeyVixfTzcGLTeV5IG+9K
Ntny+TqZ2OLx1aM5BBeCeYbgkmfUNERtk43/ksjbUkML1pt81bEn/3Jrap+rX+EZ
uNY9MqTxheI1SxvapWmO1tFcbDSfgVjsqbBOLTwMGvqk3xIFkrCq3kpjXVIP422I
3PiFEHDAD9NsRJWptpcoS6aYVkXQHDQjvBQ3LBsZKY446ZatXb1JIv9h60KwSRMU
o1RXg3s4kOj3xvzIpOc+t8wcENv4wgkqftUHDFtjXYPTLy8+SowiwclK/vynSGV1
hS9NpCu+CF5UFJHAGt8dKFBbH4dKBpNCU5dVwK+GsJTX5tJcv5y0uorHq5MsB+9H
fbDBIi8ilA07PcF/o+z+Y25moZmntqAZzOdX4wxRRxPz7CFa1PlqSa7t8Di4hLk7
dcVIFrTnImV5DzgxJhKJxGa+IyEsWczwuIOMeXhNCds01APAjMBUr3tHvjetVXR6
GVZNY4DFwNa9rNuykltwoSARELCj0QWPE8DEyYQY/DTtp8LZ13LMirerBUyxmNTU
9GJYfCat54kqPmnDR8yUWJ01zxvJIQUlakdHxEr2vrAYuixuidcnonRxrUWMl9E1
RdDNA68tNrPH8O4SAvKquQoBhijjnn1iFBuFpx/gEWTluf/9HWHBfdmo3MBlh24s
2ljLlY3HoAEgojT/RVD0W7xfhRAKPp5wJosIr2JQw2B/IonEvLumfuv1L9MJqkaU
/Yg7g7GhLfiAQqlHnYoEMQttuBpDM0XK9DLxhoFqd8JSV7lT2UA7DDRIZReCy2xX
+1ctYAtWEsOzVFtrKA6bvo9jknGUPanFkR/unAh8h+VNxuRGFHHFeih6RrdObI9p
/CRY/yun4I66UkSEYvvINvQ5o0qoTvpzvSKLcp+SCwATPZhN01HvFmQBjd6S/7ls
iqd1lXGQdR53K/vcVeotHPmOk2284Nu8OcUy3BgTNiafdV4pJ2Nm/hXxXMXbtSa/
+67vzytrkZuYtLVfSc8jOnT/uVRoee+lKNXxI2/DxkIEQnSvYQPMOrJ63ob5evRv
W6YriU1n9Vthv5jBqnTaHqq2xLKmT12iMJE608OiniOW8E6SdaqjiyERF8Nn7DFc
B2cajmLkwQ1PeoVysxH8+TutYsZKT0JeylzO2CrTNJiJqCf/7iHfejChD7PRUQUU
kqDB4318kHqnv1S4taupkjdnEPmejCx0dFfScga3ApGnfqHghVFa0qj50n9M35cG
ZbRdi5S4e2ar9jkO4JhCDXipkSc2DndXJeWfOwrV9/T1JJLZnJrL4cC9ewY9RalV
F8Pp4rvXPOyny2nJxRHpdu5W+kUqnVKKcJghiT5fU3i7uZEaIadqv33VYJ247J12
VoMMSZCBnJFvNEqg4FOOiqWpQJV6I7DZoPg5CrrWWn9VZ2aL4lQEywEUciQ6LebO
ZLDvQesQIG2JdH2UuJ1KGMt3FaxOdBOjUELEk5y9nReO4BxfTBi99Ae/7+x2/y2I
re9A8RhGZ8Ntf1/q8QtjtGNSF8UYcS2v2R7ykB3k9AKPUNKdPWQaihmvN7lWiozM
SD2rvteBHexb9Vi7Ic9zxG8YKEX0vvX+U9LKUH2nolys+E9zf/Tw2IkI3w0gsWUy
wBx3uRr7uR5KJxqZ9768BkAihBDvI9QBE1v3OLUvcwGweMm91IbxLh8yEm4B+Odu
uSHo8seb5SKFamValXSn/xZkOewTbi8E6cUAl2vWcUSqae9VaLh5+3jBz97T/LK0
1fMU/qYk9d+Q72j3QvZJ+qhLTCM1gPjcWOglNyPcyFA3BZpivjouRrOtIYrJc//B
OJmue6ITuQcGlQZZCioQ6hJwCy3b5LWHbnnGpWqRy9DgUNsLwEZjtACZsEfAZnPK
B8QO1aGHZwvchkBOmwBhmhRL5/TPbJp0MrTpwu2lGCt7t76dkOMuvUFdInWXwrH5
SalT2Dw4QisDGFXFQlXIZSh6UmV63kM4TQVukDy8NjKTRQgO25TGcGnUzy/kSQeN
ctxdTr1NoUzn0LwAs5t3wEv4x4zrxgOLUNj5jZQKck26oSKBNqjMXrzLHItAfgKq
iU9WJ0YznT+iftiJhCyH5x04qGQBH45FC5IJMgGCo0jQ8qRXc3yC3nbQePJd1wIa
RReiRqKYExNdhauvx5m3vjbZ9QYhza8of+eUt4Hp/5aACXxd9VE3e922opy6PvhW
Vw5vB803WN1zllux3HMlYiuGXA333cbwi89sWNCwuZPpI8iab+GiWUX0rY3gaX4J
xlU8KdUCaVMakzw9E1T71p77VLtbWkQi3BJCOLahFn+ZzLkBu9T5GfQmqlFWgJIS
NjEU/9neT37FXn+TaPnBR+/wTOFpPKYysHr0aSk7dAQLqgeWdcaInf0gRVc5ef0I
x81uy2HrjWLgtMpfzwKFRbki0ykPAgnqfshTIsmLxhF06iGskWE/ER2/rDXGuKLO
oGvCKenI2RSheYMKSbxQsb/agEJBX0hFkRyyibzg5PqIazpDAhjCp+kR+ffinGTF
9yEqCKiUtBLTe+4ek+1CyfQgXH1UbP3gqGwK6g3KTeZXAsS8p0Q5oZ/GU/Ky0TnL
dy9w7EdNh4HgfwP3pGYQDEzkwSLq2Nr7i7EzvV7vvd12SX+xTrf6sxQ1D2ORttcO
uxkk0z32crxhqGeG3hPKso1z5Wy2Io3gdxNHGM9H8R28lL4iPxjBLpFHRIbjYcu8
4/sSJYoKtksGw2fdxGZ/+9fonkXxXyzFkhaK4EOPuez8YENLyHIVxf/ZGl1e2ih1
3ohnZiA7YQLC/LWraJfE87Gk4J5ZqXNVQR8LIgIvr7YAL1qM4QvJJyAW2I884O35
b44wDeXRJpmcm3DLFjJxyWIZgxb0zJLWX5nWwXfGbAONsU/USS66WmlIvGmVAVbT
PF5H86SY1H8Lpu7oqz5giO5h8ZIdFT0g0UOMhS/vMMqbfbrJMhgs9Bsu9yU27aP6
oSQpM059/yg+eMt0Lh6pFOhXAzBzQ9+MECWBWG7J411ZUHVWffqLmQz41lnsayE1
FXuCOjilo631k0MI3/S1y2S5pO3i8pj6xEN0vdQ90KOWJHXxtRdExIBDnkzzLTjI
iIrPAXNQl4dOqSRNCMTqLLL8xMOneiGuFWsT/VxwFGmR3ktO+ducVvOZYC1qjwN1
IZhKnLGnLFGURRku5nEjgWuzZynM1z1mRx+ImX6lyeSprFOCqN7kqCZGSXw90/mJ
FZ4Vjjx78cscaF67hIZY85lR+NEjjivDJ4VEoUTXUnmdSlVdiFNFdLOZVuCrUOe1
n2E9ZppVfq6AWl+LRanJi3DoT6j6jM7wZkbS4+3t66pjS5utmHj1J4MfNJf68/KF
+z1OwiWieIj/vR2dy/8WTf9j8St3jgZCcDAwpp3kxDzm5E0ov4q9nVOKLtcWeVhW
P4D2xAv3j8/NSd3u4L417bjQN6gsmE7gw5N3cY/McAbL+EKJvziL1NFKAb6EsJZS
GHBR7adHy9iWMdNh/0BjsAyG1pTZwgr7bwGtglbzGL5PENrl4LL9bissNbIrobDN
a8PKB2cpCRJcysUrBdA+DYaTZnHRCIh8WvopHmOFVngTMclZvV91TGIGjB1muIYI
kGcabeAwKn6o+5Bw8L2Wy56WJDM2MyMqKWsAATNosSKd4C0G/qI36w8bCfFJpgiL
niNHksC6m59Y3Bfuaypbr+3q0J9w53R+6uu+JrSO9SV03QuwkNGDbaBA9QC60gCG
89LHvjRhSP9qwmjgXBR6DJt/cIdtFG5/xW1fiGb0vZ/gi6jQtmAm+u3+aljArd4Y
JwSeuhtlDu9B0hlohj0GmMY3j2BGOvoUeoEABNGshLXMU0X0LSzo1ovBrcutesbB
ej0ijSFd2cnQQHnywy05mrXNnet+eD3hUSfImOQEAzEwmR21/66vpx6GokNRUrQh
h9jE6+Zfprprt+NToPXp5dlFh4EuRs3oVHBBmlN6rkV+HaPZXxVEpy+QBlYiwts3
WOM8a4D1NnrBqbnAeaeQ/atuYcai7PdOHZCAKayFM2sUpZ6ZbFDfKTPnwfE+EvJF
HCuXecg+/hr4/EBxDXGJcgjvxSng7GpLftd3Tsk2i93nsohnD+wAa+RdvvR8Dytu
b9cqxUggvEbD2ki0/VimCr1X+I3cMb2ZGL9z92SL15QogckUiaPWS99O+8YM9C0a
FYmmPZbTup9wtVJzMoe2Lk4ndMCQ7sjzMSqA0cV8BsXi7Qy+op+eWrRCUL3vbgF7
H31xeQZcoRj4OdmdmgA/Ra0ezOSnRvE4qLDBbWzyes2U8NeC9Z/ub7DFcUGJ/xcC
e0GXCRBoOt/tti345pTNA+EbfaHB+E4bZOAP2So+CIzuLs559zRQFXPEsWcE4Ldr
FaNgRt5Dh9BlnMlS3QQTF0Ehz6ZzIeX1LJkUtCWzFfmp1h1mZX5E8FpWGSQNAJwD
Q4u33rGJqpzodftVyErOcwbt7p192cksVwYMIr+EnL9657PjFYfzuqS7RMKzXtSz
eH+BO07Zftyd/TMnMTJRTW1CuquZXNM3VfFyCnXpVCzQMiHHzgY7CtyUXtrc7Q9u
yrBIMay04umX8Tj9TB4yjZfZeCxYEbyF+JmlggWzSt/AohIves5b8TvsI0/xEJLB
q6bpGYsIaGdowDkBh2weTrRyc3IH/uVkzGaSdnK4gaKu4QRaySuIbGodtNOQVMfN
bDIumxSwFcNjqDS2V7iiW3EhuT15Yq6BfScnXfCSHCDCmrmxzh28oUgrKHUlgE/M
z1Y0HlCMcW9zs18KvqwxwL2gbW/5pi+vgIpqVt9wzzQLaaRFvf8viJGYuWg2a1HE
n1aAPr6jvExlI6TzRiClLSkWbEAczOTt8RCtlly+N0WnINpFyXjzOBTmq/z1KO15
HN2hDmH36E6upWLkJkx88Kw6TIC/mzE9rYUyLq8UwHKS4H154seG1LwWaqvAFgQt
3hxVU7JVIWQkzsiIzYTRPfZVUlGz12gJy+KLb1azxNsFR2SFOONMz//kB07aW/wn
Bt/zAQQ6b9KG7lwRJVgTWVO4siSyuLxp+gl1Hu9S1FMDYdM4P9fmQ2Dpoz62Geuu
fEIyt1LaKgJGfdvvuuwOk5egG2upBjzOJ+Y9Kx1AYj3rcjmXvJtJhzZ6JQ5Iv5d3
RNDdN9vrwEQ46HDb4wKayFPES7m7wwoihIXrisKtOpDeUMEmDZnRzZKSK5VRh0X/
ZX5X5ZLC63V7Cg4DwJRe51I0IlNU83AASz5ojE6275wIefK3KH90tPclibBNTzYx
mcQPR5n9ALb6dvMMmPKym0Nlcs65MJMk4UQ9efMkF4aQ54pp4JAtzoUOgsqTk++A
7kRFUkG3386UESLxl/JrnVw+Bn83mJFCNCh3Y1NkN6OHx94i39mNRnZAi7QQD9yF
hqVpS/6uF8ftcaxjZTuN3WyFF3Wyjo5VgmT75P402+Ku3sqa8Nrdoyn1XbALTU+C
OfCLE44Mb/fZ2fE05fCNKqt5WL6BlA/l81tPxyioLVF4rktbw2qVAOR3a6aVMAtk
BaseMsxi20Ebq+in6nXjlVn6R5NVZcN/B1cktz+8Pys9UTfVDbDmjgRQh0ui6X9q
xBuOTit0BOa/29ZNbxQM+dPbRfXGpJkC1/oV+g4Q5N7qJ1KgbhWSal3GfafI/ScX
VuJt+pTP1ik+43kU2fumvXfyRhIijK7EOxprTX6pIc9MMSRDaDuxxaIJp1BPPApY
ntEWDh4Djylge90Vx5q5CkEKgmccH0g0HAsBYG1ityYb+/dbR33KIllCyM+cMjR7
LA1yCiyEXMN2VXqXhjbVPbc4+BJdw2P/J5TQBYFqzZylWSgXLhXewBzcrjBOLDkC
iaLhMQtCTsrVrVEikkQ6j12ujkWvKeadGxk2ingxEED3DYtF13bxquh1yvprShl4
ZuxV4OGHBiI2VpaFg4gPX/T7AWa2RAlRYZM8YzzEOkZLBjAsqMg2aU/AUTB8gIfB
BrRnsAQncyEqCSYUfNlrzBo33ZZPape5/TA7vYsLtIkw/VLwUzDqLb6cJIvKXNjH
3YuI2akRgXbHQJ4kMHI20G2jlQY871TxdIUK7cLKNq7mKKe30/RU7Id7tFYxxQ8w
Y1dkzshIM0Y874rPx1tN9aunK3jG85vhIub0dbyp94UgkSFNHI0E+f/c0kl/Owte
AXOzptq8QHW0JM+xLeIhqnuWtkFnn0DIIeXTrCScNHIlarHcZ1w/JT0R07kDAIu5
3Evghv3lfANMsGLD11CZOESSPUNUAWxaeSNggusvWOVr8oLxGYcLYzzUfurfkfQD
t3a5c4ExoD5QXdDYIwhRoqXVFCnfPAOANHYuYe73iUPOGbGnMAjmRHMn0WjhR8Wl
OkbURiQ097LfSJNvp1vbVApBGiIvlmdtvN6zBfNAD+Sa400y2+YGgi1+/LZZJXoP
i1OzC68zk7zHGXqcLtKryCU0LJRLYJjtt+XbtqySet8cFaEOw4BiqABwOjHQ0pEX
Do/40S8ckTkauIsbIAgEGZQU7BCIaZPyAu5q0apvJMTIfACFCJrO+HuZwxXAwi8g
xJPDs+OhA8SgAhV6rZyzKgVJBbUzVeF22NekDakHa+/g3qkvarGsk8+qS2+3ut13
juCoZNlbJt9C/qf7cm1QooI35VBU8qqIXd4lLP1c/JJ5iAN0l+SVBBmxWbvdWSS6
iLGQQwbg8nKvaAzjp7z5xbGPAjOGEK9PgW3NAM9RJWg4ALKWbu3B+IE/Qg84zfti
WKwOvYHDJli6nuhIbBBj9gbLXlU32/sf+sa6mTnifuERph1ErfU1gE8ltw2x+UYY
YP4ZKmWmWCqL+QvIZYPSCdchrN83eHRmUQmyGr3iO++D4SB2vncKUvVTRS1NYCPh
z4eoFOsvxVEzVr3+93aslzhwz10qqAFB7fIFAm6i333CgC+fLM/MFu3u0WQyCaY9
M/sNcALlztrVzIYAwoQFwOtBUtwyDkOjU14bhJQdRxwwommTci0adDVxG/bfu2rr
GOBW9auig6U/0jFjqOEXF/0vwZvcjTHUJrcBEDI1xyeTx594Bw9MVz7feb2kXU4l
FrNjfBuIwRAuLTRIq5SdJyKQqTZcXNpNyrB0gJiCJgJ+QX3yjrL8/Y8KKEJ/TFnu
05J91ZOxNKYgXdvmTzXULGgQwueylEJPOAFyMKOxSUpV01wxXpsbblVvGJoYRApY
UtC/5RwSNRlD+UR7dzxE7usrLyt4W/lAgvp/uMJA5q02WdrkQcC+ZjwLvw99Oamh
aVRJToa6u5/is7J0rnSoeGHa5xBwl0/KWzw+RyXSA9/amb/EVbN7CMEdvavOIHjb
Vs0AV2bBqO5c2diPAn5NQUCY7iMt7/WI8FlFViipJzKY2S5JZPbSR4tsZBHFJ+0y
J9VNCGMWb7abSkSKYV1mdCJKh9hB6vLm5JhkmZECILGGcpxlLzeCmIqWRx3NNv//
21+06j9k2atFnYxM6oRTOppeKSKheNSGRjdIen+OBvXUIUDOrFZnTm9laOclS3ls
AVkF7wnnirOJDN+wXL0DmA9B0/s6XgrQWmKevPG8BCybjgQGTE3XlInjpmAynzJA
8907TKtkbIKfZ0NPgZGF3wul2vN2Q+VsjJfI+rX90lB2uB45EIK67uocf0UjcON8
YWzvVhFfVGvbomORXtHDC8yIxhzAcHvB1DQYA7mb+WpGuQX1wT/6nnWLyvrSFrJJ
4swwMsyiFQ9zfDuAmbfJ1ZsWzZ1IzfrS3N//gkuj+HPJtC/B4fWGCuon7tKMO8+F
Eotq0JvPFUWDv5X8yYokIOHB3o0r9C/V2JwtUS5Id1iDq2O/qKUatKx9qzmEYIHH
uLaNqz/ga1JQuZhGiwbiR8LMngQED18jXtv1HtgeIGUkz188nDzkw9+ekyBqXoTk
ko5ADBWLbR2CwjipIpHWJCaZAh03uZShlbPk/RwJTYRaC7192F8K4yZeiNBz/2bK
dmMzOLPB0zHb5OmXuzOnzqz7eYANn5Zjpz1lOsIStcM92Ijl4i9ETUGKgHZIPk2N
+uCRqF128kul7Td+zT/lLXU1egXbgWyp8Bam3q5rBoR1dp6cxf/n2oQpSyDje8hx
9kJPVG34enJv9rkUhwnj9e0eOCyUuLEXCRfV6BLeBNoWqzzr9oQ/h3fN/8EroIen
UR1+f8cDgt3ftvFgH8K+VEgloZNdW6PLjXhznbtDWXBoQcZ6REUWKkhLZTP7q8ol
XQuGPxMoIaB2i+pgW86Y5rTAHJVwWRdpNHGNKHzYozPZEnIPSF9T9iQY1dIWGTm1
QhErix3SC0HAyLSb4sdGKeL6Dc0m1BNdvuIKmvutIXD+zfilgw3nMZjFGW+vWAba
BXthV11SGBLLm27nCT9BeVu1yHiP3Qo8iNj2fdLPO2NS2oGP3qdWpq4J5rrv0DkD
fmJ1aqmDOGIgAbAeY0LumswPiB6vhdXWcmj5Pht9HIVYUccj39aIaqDwv/NiKwx2
k7I+3w9EHRIgmR3SZKA+R3HmwlGGWf2XuaTTDdeEpYRWI4iXEwLz+cEt44fKso97
gf9IL7OcoHNqWnrum5Rn1bppR8plm2dOGzYayJUeo2yCokYzrWcO2AxPcrTzxKrs
d3q8cB3OypLxSkJjvm5ThECcGeBM4xrciHIM1sVLl1Hyc0dagEgTV7Ow1TrYlPdk
oUffA6LcmQ/EzlbaFOiLGo1V+CZ8NhuwPVRGb5XVnd67j86ureRmvWse8fgQaUva
jyY0eSyQ+/tbSwXs0rwfEwuMg50kb6mSF9w5yq5HmDd8vatvS7y4fxn6PcTCR0Eb
NLqS/Al9rNT6u0eM411N2ZWklXW0AMIN/4B+usk8c9qZJnpiBCqYm5159NFX8F+9
8huxOhpELcioligQCe9lumpXLFBq8InTrJvv0OnPOMIPI8Jiv62J2h1ryla6BrGL
VyK3Ehud+gXacWZejkplsNC8r5Z+pR3/KW1YFfyP7AG3tdwhPLVvoZ8Ts5iUevcs
BnUCKg83gv9r2DOXkIX13kB0b3iAjJAoOwW9dg5YWuwSLiRJLesCw8Ox+RBKqPcr
rGdxp6iAm8j16vTLI47gPJ2oznQgo633NMT3t1mBAOfms34xqyuwJS1W2KMAVvIp
NpRZbWkktm+rPYa+uEOaI6cV7mmd06g5bfj62D1h5OvhJkYErnNGAiLkNfSDxamf
NK4ybP7F7bmpxF0BPWKt2QKbctgYzQhTbNQZCAJSJVaXjYTsJeXtmZrHqcso58Oh
CyBe9SLunw7dSZ/iVenD9a1WjPzVXOLJqHqXDv1ocq2jlxYn1ZIZNVw1Py9pGbPJ
tOAQf8/oFsECwe5Qmto+w7BZIXvZQ2AkkktXn8NVlEXnVzOEK5aqnbpPwkGzDWYb
7fin2++/MGPxfXtFex75vhLYFPi9o8HGZDvZZ02rv8cwH/feCmLSysOu4YNNC7z2
9ADBhW6rXhOABZg7WL0dpBJl4A7O8Ikekq4Js/EwO6HuVUvlnqYfNiule4h7Z+lg
d7i3mP553qWYnryVYWOQpRIN6RexMLvVf99csKTZLGt5YODMGrnokwPCwqOrjGpl
Q2DIHYSUAmrvHd5qnkvy3FoChHHN1ceFRu8h1fAQ+WgToOH7SOElHXMWPxBsHrfq
ijHoqYHdSmo/kLTK+32DP9mQSbNq63PexUWq+NIMFtyiZtz9qQcjCalsy6p3jeJT
Z/RrDE4lMVFh5fJhsarLcdfe1ynt0qEeIxJz06R6VevuMHtKIbKFHZSrKwYVZpr3
CFmxFNNOGCPXgLr1BZRlSiW7jlx3i2INilXKd3Gd1hZp0yH5hBL/GYxGTcZ/auLz
4YkwXL91NKykVVEBzdk1auGI0sJ43FCiqVr7/AuP/1uchHSjR5VlbTeKLZz8B82T
u07LmIUNuSupIK1S8d38CPF0JbTkCOxUAnlvOS85TtJnyzW1ifie0uDIFw7T+1rG
TWzQe94cAMTbNzXahDj/tqZ5lcl1MsU6eChDrztnPMh47yfBY/aA4OiFZiBdaXdx
ad7rDFcJbfhNKpUGFGIFT91Y9JJpymMN5WFZnzF9GaknJHjNU4AVH5Sexws+YgXt
w+l3OOv4Sg4d1NR9jsv3Pset5mt13/F1nZVV2ckHYLIYhc7zMfBK9BADw53V8Q1e
FTM32I9H3HSauoWjvHikaPymfBQw6ZG6gcy7C/sGS8UjPJ85fZBbDHUmI/ghboFL
ErjEQwi8xgX7W33cPsWfSfqK0jLTjywCZjTvvmmkbzSeei5LY2RqrzuzkkWPuPYk
YYkLgqgzxYGzmZIM9gOfzTABCVwEqJ38KjgjVG0umC+o2AzG46Jgkdxy9/Uaig4r
iHzkzC9Fw3o0G9lXzUoMT3v2AdwnbpxuBIdk7pPNMAh93tIvZCxux+7tVsyN99x2
bNoXdxZA5DnLu4cK8AfoHKM/cfpUOygzk3MNoYXs3DHEwbL9LYqMFp4ya0LViyxy
btlSjM+qqrjjHvVwu4t3j7zpOn1xu9BHlMGFzODnR6IiT4nyPn8jYh8Cbr6OD+cW
DVRcLYzyG17pD2AuwmJbdjITFXjqBDN5r7oB7TqfGszYtJ4ZSRWNuyV+9lIe0xN5
k97R1csGYGWwpVYAPetnJ52PNxStge3Nvxtrdma/Fk4gTfH3X52cQlKj8h6n+Fd9
EmO5/f/1bc/EUpZtEVAO78c3chtyeHSMy7mhevJ+SZbU45NpVz+zAtCR4jvSMcCZ
DS55l+5N2UTVbbM+ewRxurPjJ8aloejWJh3b0SucSInFbaBa/6S2QsOzzBw3+S8m
dfuj5LJIxQMjhfhejoHs820DNvmE5G/dqRpqHJQTrskJnVjBpdaMb9QC5bV1o5FY
PXwva4CYTLKBDJ5Xmk15TOylsM5dWGio1HiICVBopOVHh9WtSC9AejpnQqTOwsUv
BjI8eGoj/eccSUZIwzoNxRARtjINI6XLyAOXteZVjs/S+QN3bK9RbIE4iutDxPJ3
SS37czxvyK8OFnVoxj+wduQs/E+Ug112R7ejuz9mizmneZ2jK1lKHcg9isVDenj1
TcRapf05Hh1G1lO3vhfF7psGYNkShmGA7+44qf4Kewi/YZfAs7N1KWgmKQ7XutZ1
Sp+9V8ydc5E9AsyU1/ddFX65bgmClqlLsmY8eFsm92CACmuGHtQaADMy8B55HTjh
VdedOwTFuV9X6+GML04zoQKzExKNKy9ztaIjhZ8GlZ+NdNjWnE84mwrgbVP7saa8
yiWxVBzGWbygFS9IOKVlmrFM40Vai86/aZFenAh1aZRy03ViHAu+bxwPfdON2NWM
c3FJBQE9a2umu5kaKlFBm8O6ntfc5oDODunLAZg71jLCdcRyQHFExinJyc+rYgvh
PbZYU3HdNgI+eOxuy9h51Cq8PhCPKwqNKlWfAyhjHAEbsc+uv/ccJSndFn7OGswL
Ki3g5+tkb6T0WEjNaH7L12zdOYpc3mamYPAKcZJSsM5KNNu2hpUXmFnOpn6FkrWD
IfBQ++src4J5l9axeqO6HZVAjhHClzV3zOyXY92Tm0QRzfIYTBDRSQ/9OaYBNG2N
wqslapMA0TCIKiETX11r2dC/Iv/xhhWjq2Hs/ApO8dhplhCwkBENVwahh5Rdz39L
/Pa9ZKDPDUOMs9yaZPxIdgJyzCt2kwv2xE4gm91QXmR2EUCwpRL2NAjEmf9AIsd9
5rgmc/NXkhghcumtShDoQRBp/6d2ZMy2UGWSqqPxAIQMs8/FdgYxpa9ybRjlSxx4
xZWtyNKTfdcRM4PRFfVAVd5puid86DXYgliNVjL66Sv6coftWnnGrsnJkh3hJ9qE
Cm1azbuCDG+bucnB5qMD84nxTPYQsgaOjo6wspvK0ok5B9GnYvrcfREMt+Pjo+IQ
vOTYqHTf38sUymI2Yg1otfBPOonasSTnqJH5gNIDW7dh2xPspJ5OoQ8hU6Lph/u6
5GIcrOZgM7BDT8XnvJZcbwuGHpw0p1jgUQl5B+2aAO/0PnKJKlg8b6RmGHWibPEI
qLgCCzzs230WXq2zc3PlGbGW2XkqlA/AemCy+l731p/s5he7kUZOUTDUdnFaxrdf
dyUxFocy3X2PaE6UlNERO5Muf+G9PFTHHfJI/ESQbzXRzejFKNxRsrh3Rs74++Bi
0/8cjfogeqTRFNZYLgd1L3yMT/04acDSptkpvkt9Ll81eH6lBXq8jexDB4XdgCtc
hSwaJuaSYal0ZXoJZvDDnPedlWcm7Y0Kxtzop8CD5SxWNkW+AdGZmB6wXLmgcllM
UQ4ojH0xXWSF5YL8QQgLWeKlIhJmRIYJg190KkGo11pN+zo4AZBeDxpAVXgYHw2M
ngeUZKItUq+UDoZopTdoUeYH8xl0R2ki7hHELEOd8v4fctkdFLfbIuC5gJyp4YgI
GPb7WPJIxt1aiDuw0nXPbaixijxuY2yDmevSccoFH2tkPnqDX1PduVkXKxeJA+gz
BsWql2wOOiCQVRW3fZ2MJGMu/lNSOULiKh6SV0OGURn/9NdlwsZ3916ApPkhGZcW
XIw8SONR6WADW5p/CO8cMcqXGjfuoCQe/h0+TCtQWfWMvms6FMJwzMZxUzu0tamU
lbo+kJ6I8ubWG21rFO6VmCwCSvui4sznMZy77GPfVvct8mtPtNzp7olnE18j+cou
YZ22ltnWdGPKmts/TBFx+me3P/Wh9vXZrNQpTk9OEl7xgp0fi6gIP0oXU0LWxNsP
Yo1QUb1L0YA5EjlCfFiVJcJv2lMcsTyuTGeETfz65R0grHX2wYoO9/5EtGSlv3eF
lOQPeZQbrIZPnILLCkpynOU8QL0uCAuGMQObjsCtLQxNiLodFHFHKtXLBB0isSt0
mnp9mndbTZR1ttIYXLT16jvT5l+pkJXHOO3eVShP1DCqRJtGDu/kkZnnyzPknHf6
pZLo5C9jbEwEfxPx4mNZpDL3DgSyDvPZGtCuDsDx5i0SzXBZoMAIwipz7csQHMSk
q12HtUA2YWp3rqMrGg/ZIzMS+hPzIYF3hrAZ3WV7Ng7kGLkFl14fiJN59SsEw1Pg
29EM2Vr0iow3oeI2SKzN58DX9KBwK+wIXh5p3Zoi504XigfiGsiyh0vJn0/34CMA
q21kNUvRH2qjC5CIODxyUf2Gu+Nm1QeTJbuj57Xjb8ZgaO9oCsta0/tLMamDms4I
+RavMwlEDGXqZOfm7CiGRwKPYHijAlhh5DMIHYcws+44N/I11b2jeKfLs4+gmIRp
++ktnfr3NilK7N3LJowmnxlGHIqx5zyEXMz/yAVNlIRDuz5GKqGyaYZJPQ7DZx8i
a3j7zxUaqq5jNGEM4v9d2SHuDgDRVQKhPvDQoNqFUxpu2c7qIyPFhQMJzpBFTPvU
AJQlS51mTNKE2LdrMqQ1GzriSwmyHGva73md+/KWr+fONn1dk04elq8CzEb05ony
c7VoZVSeDirlCMhMtukVo45nvyhxNNqzWvzshyDrEvmhJSU78I7wus7Ua5ekcmhZ
30BIxzKtKjy49UPbgBeM+RpUFqwrBMLMsWHF8tai34Noj7HhsaZB7/Ov5gMR8G8f
hW0RcfLo6KngrODyFsYQmL/cSdrptlw8bZagXANg2gGxzExL8tQqbhE4/eGzaQOv
mdXLEV4TzeHqZXGQUTgfcLi5PAA4zTWkvqO2W9DM/zEW1IpOTc14Xyq2yv0vz+zn
m7qEHHXSi3NLmAImwGH8IeaaRXPwuXvnzCTitSX5bsu5lSzvpWL94hsjmNH4mjs2
bFbwcnBUQJba9XblypVW80bq30eX22gyJSbJhL5Hs0CELKRRxwRedTBckCxWdoZk
vqol6QCJfPEUDQpxbb4OEl1+S+YC/VnSxjmVHsMAJq+66BNSw7U1ZfBGTFMC/71r
f0ZI4mObln2miSNF8+FuOLX+TX7bokCXYYrz671rvG/AkWSbcOyRXLTWJkCWT7yC
fOMLuPXL8yl10Mn4QGCywwCPfZviJDnr7YIwa/2b8DOiW02SuLqSp6B9UG8sCjCz
AHFciLNHMi7jHX+IUZtw6r29fpOqUoWTfoth1+3VcAVrwLTlCCBWSbvDiC14lxhQ
3Rdv2QqShQnvW0c+1H3kJ1SOICsSJbZtWvovl+zpP+7ywj1V57dPlMbd5GWri0yo
I9zXTyis9sSCcQtr5b2oW96Baps1i2rX6ugOjpB8nvIv9EODGBvXRBnlC2J3Nkgd
vvMxzc4alkSGhxCReWw4idj5G8UckGiXhzAPjiMGImCIjqgqPjL6dcfhHGyMH0Kv
v8JFaDNmaLKRz6HJrbYTYqXmnG5lgnJxFVyRwTD2jnLHj7wc9T9ydsckft2Zd+iP
XRIKJtiy5PAKs6TB4Z4q4PaEoOKcETCu/ZEDZF2bnX0NnIcqwS826RLtlmts2vtO
/CNNk+S6HzFPu3lEkZ3O3GzcBmrCaKq0acq5eMC6qcS+nVFduKW32aBq+4ZnguS5
D9LkL/HColaRNCbNPJ/XQ1xFkGVLi1ffV6hXOuRsfy5MVQROf+9yIJWvMsKnaDr7
46D+EgD7LHBM3MvEUUJKhZ4YytDjyzU1Ym84kIISrDJI66Gt9rGyJueQmaGtppWq
UF73QXYWgeXOIRwtMJY9jZbszcTOuRqaLsWzbJY/Gtn7rhaEGog+6ouzfOgseJJU
cva1BdTLxmT/kzvf6lfuWEgml/+ZZC0SeBd8Wz6x2D6Td+g4yeKiMVs/VxHA+WCk
szDBRQ+aeVzAwM1rNi/0uXor536+DG9vKg4M6XCmfUOYCiy356/WFLj1cgax+oxq
vLoe9GvtoWEUGL+QHWEwUCILCEtTqParvVr9oo3jmx0u6+3gZXqTIc88JK1TgptM
K+IcNUdB9wTbIhfmIrdLUQpQKL2apms2e68ttSrtUnmUWsOtmxm4d1hiv6jJ2qrC
nilVTCQ/WVfHMMt+WYnmhDqRqYCYrWVfelnTnGrEI2hFeh6H+mydPU23hR7aMzfO
wP3x88CkUz+B/zV4s2x4dDaPs3QcJkP3R6FchRNbGiUBvKQmuuG8ssMxOU4bucI4
ek88sBgp060+egyG2HTdiaxn8WNEkERG7ngY+6BjZpIOCUaXbn8Ith6TyCe4H2yC
y5zkEpbYWbbpvO+zcJTfjWg1H3fIwiMsjOxqFq++sT2KgkLt2afdhhPCHvfJXy3D
ua3eyw/5daKzRkIaB5AqMT/71hcbpaJbnrvkFWP9wjZfbLFM8mjD6vuHkrKQ98E9
cjjfEpSZdtyujv7A+/DhsbHkK8aFpqcdau/erDTpEKpi1r4OFGM7q9G2IprgrDye
DwQK7dIGz9tvAogxmhFH5WRauT1YrqVEx7uUXot5Q2R4QBqZoqvGejQ8TPtjYrnO
2EeYiqFkmD46FbJoDzxF8cFQ1vub2dy4537cz4AYaC0oE38yrTd0MORzO05mXKPg
8mELGpqecETWTRXvAiWKeMHiQ7YD7cqhxrr7JMlSRQTmI27JGi1vZzerjTr1J0W3
SNiRhByUB8xJxqklVeBFqzonqNS3yn6p8+ou4yJ/c09BOokmww9HR066BiNmrh+G
iR6pyCSSskTLeMA5nop5dQkkBJev0bp8ycjoquGOI7VqRn/8IGg5yggRR8EQPltR
8LQuH4rppNM7Tr25gRNQBlMxfIz2Q58SoF3Dv2gPPzQLXC9wwTcLES+x2AcEtcKw
ibzLY/s3cLTuVeSW8xjJkWbAeX9pnmeKN8JCQ1TVj7o6z2cs0dMG31e8Zt2gt0eE
N/qb/rQFVNJiUe+ocXTfhEfbaLqccwj068j+xDz+MDE8tkghQezw/I0wD+ZbpasA
Q0UUMTQwYaoIo3oZoeLeDz8sEWw/hKbzJU8/DpaplqSGx8rPnn/f5DpvZSZ7aeX4
Q5IanqAe2aXFtM8iK1u1jETmkkn3ioYqGE3qKnMEF85mNEQyDTil5k6JO1mYA6r+
/LO0K89l6IGWtP0axktxckd2w0EPnWs+6unfJiLBt2iLGrva6pHCdVry3O97qriT
dJfk0AOMDyUMvLvLn9sQK/V/xU3p2x6VRwqZbkVS4SufZ6saHEejC/3/GxytDbtx
1cmEZ7cVQbEiGZDHEdColm96pLJRCZS6nmgqYKaB3FbXctuvA0vol6rcupEwJ/ol
fBGfL8wHoex7vvk3tLjdv4/3UiavLOS9POwOjo4QG6EfqaSxy6Xj0OOhNkCZ1tHC
wGgrZXvoXw5XrCpfyZnstp26nXjh08yRBK8JeaLdE4VtaELdHYM3/vP47FrkGWfD
deQFGuaew+wOetTIO4g/j5+LpmyeMFkxE5y4fDfIi0XNeLcIeGJoTUlYwaPji1tV
ePqaR/Hpq2IlpGWRewrAgCpC/tdGZsdm9K7u74+gSqVXAoNmyaHJV3zw7+3htAGk
q4eMb8ughfesJp0ncKkN3eFeUGEeVUfGs55x0DodNc1LpZjCEsqjOMEy2g+hCff+
lMq/ZoL7O04EsjStAgbBj040aeAYPTosBSeuPxATLCiZA+/kaXIChIPHPX3GYgrr
ty9QNwT+yZqw9uhSyubumUjbxSODpxuOnyUvS6tTj8fGrfQ/uiqImDWblhXYDsJV
YyPGjNLWy/W3v6pFB1DGXs7NP+1RHy6izKyIl3lTMOALe3LWL4JLhmIgUzpHfE3i
jHCHUpy8MSJlQeCIJok9J5b22JHRlGX9YLHSn7uHhxBmAbt6veoDC3P7NG49Sgws
/RnKuuu34WfzpLgE7qItxD1HFAeSTL+/iSKd2UoNNnbhP+pC6JUc6fLPee1SsA28
blDxHxDb4Jo+SRw5gnsg64vySBzthgojxxe+6niV5Ht+KLHAziUEdgJK0GQAjOIB
HpZ0c9HcQnXq7R3BpT9+EcqfvIJdUWCCmbTg/4dHuhs1I/b+mDJtiVESYrnkcjPu
ScDifYmSPNUvqjZ4kp4U3Efh7K5XMuqXPJU0uGWVTtW/IS6TmZg9mY30RtEzciL8
TSa/XI4IPqO7YPwhTMQcPnmuiX58ejDSbJ+iU0WJCSmyaC1V/8e2STTYA+gfjx77
Kzc8SfITZx14GZEaIa2IT0qN2Av1T51sl+7nwZmplrlCLFMmtUOjeqLhGu3YVcpq
oKKx9e/UytMjk4AQwZiw012JpVsxacatskMqC2jO/jXH3SY7vykltr8iQURWjLFu
IMERHFpaRwpTqVtC+3hf+g7n0MLwdVPxP5O6+0OooZj5MvPWnn4V1JYj5qi5wgpQ
LixreZ4MKALh48KP8umrpfmSjDVMQq/bQ2vd5Ly5YHfgQ45KHGoM424sy9JqVGV5
syQBcBMhAolT1jtmW0gRx1vKhWpo8AE+vdnN9WZSQcowDnDhBZkyhAKhn4R8N4f+
pUHO9Olr+92wsDJjQiev1BhECV/TAanYsC9QyAkLL48QHXssWGh+BGrq08QHofTm
sSLgqpu8goQ6HXllt0yp1Krxfqx6NdTVonW5dNlWGK99Z7qWOp6BQv0FgSRx1ULl
eoQxbGz+coztzmxmO2j+I2kBxSO1EZshMi4C+nCw9jtiC8OQEdV2130NwRmNpfo3
mNJdKjjN4YhtOyVYKMFZIUeWvZn2JMRJGPCw4CM0Hx4X3rWh1Ro08yBI01ePx1qk
dwPUpr82Kh3AkkjKw9QRDaY2OHTqEwyAN0VXP24EtENkuwXjEC3uVhHYtAcRveZz
THdN7x2go5VkN3b+aiUszAEy2xBapSAm9i4AQ7bUAW/KC5jp4H4qpUDCOg0wZ77Y
e4U51k3uU5+FODMV/y6YXjKFCA9oSjbJrlkB4aXNJs1xDmDVpXQ9GHivnAvvCgpH
9je3a2MyfUJGdJmGeiId1Gi2WkZIaEnC2kByUB9/ZDt6Ub4zQhFX9Yqvk/sTIAsq
2ivqf8DjUSTUbszAhw5uc5SSWA4qeQ/N9HBOnkH8pcDQO4Oz3e2F7ILSE19GD/Uc
0f7W0wP8RyPOvqRCKq/K8vYSGCNyNmDBNZ8sdXMIkCQnan2vKHwR+DGU/FmytZ8G
7NzoIhLWsWUEhwE2V/awp9SSo5smHwpgOoGG7BNjQJrwssU2aqLxVSBi5AxTbFsU
BEKLZwb9U/I36UZdL1SdUXzve3dvqN2cFwOUxmDm7ZgFtl6kY2lJ+G/vhBdFLZv4
01I4243C0iy6kyjBaK+9NQmgC/WRq6TxyOymt9oXB+b3UVR2eg/nD+wRbIsSXquD
nyIzYZgS8EmfM6ZX7Wd5AV68pJCeLxn0Lh51te1/i5jJacLzhNVGySTtg/mJiSGy
WvTFiGt9WZR1wtpXBb6gW/f2gQl8j5VZg7MXY7tlT5IfypjufwVio76bScDqFOVa
kiD+Icanum47t85C4AKZwJNHJTD42gsEHl8O1rMJutwF9osFQRUTTb40X/NXqGa5
G9JrC8NM/LdzbNT+0z2T236GSAFD/81b8ce+7WPalo+PbA+jeZyGP/u8kyn+gp9/
P2C9FTeXqUsbdDPqg3aNs8+VBQnJYsmak8F6331g4tmbjwr6OACkTqxwxHAGLgAy
Q7++68mxQejSJzZ6b4ONSesOVUvGONYPYwoz6+ePtfnY86S0JXDVSJxauCmVJSAK
JUy5B591VYdEtqsXdlxXyAhnHYNtSG+8l2RraEjgukKRqVtGubmSdILYnPPzPUVx
p3NGTyeHDkIMxySruIe9rI6gWWVdy28sky+guiCCDl2iVGnuOw5dc9ebcu/emxT8
NvXUdo/aw4I0k8DA9jGCxqxP5jKDZn2fDRMa7VGcp817p21occzXdhDd2G1W78Vi
TpTXstZn37/xOAUzWXRKHsobZEQ9/RxU92tivgOM1ZQ8So5JUqsvAaAPCt5NCVUT
U1WvVBpliBpbEGJ7n+CD8qFHczFf7TZ4P/l5Gm4Z6d8sOUIvZfuI3IL/BiZrorJn
naBQ1wWeWjo77kfVTxZN5XSzHghgD9sVew1kuaR4fdMTYyYlTJ8H7SMyi6hcHq4D
dPho3CLxxrkipM7luVqRbeavCHXjJRgHhBRUGtEmahZAA64DuGlYgIpAITgWuUep
PNUcK/u5/jpepZ6ObsQl/Uie44EsTjgQtqv6HE7ONon45XLG2B+Dv3A1m76YMf9P
hZZk16qsNkAQu3jqf5BkLsNCaC2hQf77SEwbWYVvB/4D563KjTPyYP5g1reqn6CO
6IsGbx373ldyHZhWPRTXfgwF1Vpimx1Ju8YUTaWo+I277gtvARWTGJIenSVrm0fM
ZlvKC3TQH4/UBpBXGmGq0mIZoxEHVFIrgQ8R1TM8fMNViZH580MaYrMmE8m0opJm
ezM1APx4+Im+b3Xq+QVYSr15WX+u3H2omhPuATVZOXfu+kHRgaP17Aa7oyXZaFko
x9TivHXZP4iCJ/OqQqV8gZMPpdKEkJmigphom8NDwY5UxOp6v8nvoBtia7W+irNT
BQVRTPjf50uiEj0zLT2IkIIRpikfuUQwLL00vwFyP2Fob7QU+JmgD4mAVmtou7OU
69CmVkJSaBC6n3lrxVTQnW9PZKCs9sfB+lvNZpzhkYLV+2EL8gWdGPzw77QR9AjD
6YDZ2xPx55PeTRDTh3hbCOhFMBzX8SH3ANqx8pNAbR/I8nIz678azdf5RiiIY9H8
zQw9gFbj443FymJ6WWs2YeytNChzKTh+t+Y0i4+UTSUh7BsTA2ZWh11pEnca33Fp
l1CmLoXoAf0/EFYoeG2g8JLfydQGUJJyPbOtEgn8Llmw5v9ITCAuHGD4JA8O/B2k
xyHD8niLRpu+aGD5V692YLzKDFJMJnP7dyp+8e5FdWnizUkhbPXeNbXAHTAyvgrm
RE47DgGzBgf0WZ/EODrjltSLWMIq5Sn7x76sE2sjrjHpLGOexq5hvKlwjXI2RVs6
KCcI2XGb9N/7/2P+oOS6NUHIhwv/vF5GalAp2qG1gMrFv2Q3KY0PP42x8JkRzvLe
10x3rZ5C4W+LhkBgOHFmP+Px607cRnF6G8AlHAMNKlM9/tdHVAiFMVOlO95OhDV/
cLBbkWwuihEnhwQATLlHc/LQeGqpiKcXlMurD9jspa2oPQdybbIMao/gRcrOF4t6
ceUjRKpoOwnDI3JxxwoSnM2MU2OJi77y8IX58EVCniDUyTsCxE8XusIgCX2Qpq2A
S0YSLbSQMMfSEsuRhvh5XFlMHiu+rVyGs5OiLvKKCW4Ms1PXYFGa9g6BuhG7wedi
rMius8ER9Bsz707lRcOWbl52txHO+Ch+z63Gc8S5I5cfLsOJS4VUtwAIM7zJOLfk
gxB66lDGE/dtcmHNUWQ9Vqj3S25Q5nkEUlqy4vgMbH5ZhXMV+gyNH+t2Bm2qLPZ6
b/IU11jvkJfbkKQXwR3QC1cDEou9osWauV1LmfTAgz3oW1eKjtnF6gU6GsoApLIf
IXVF652URj9L3nij9wr6wNI6mdF7R+32G6vvqeqllTpeYwLIF3BpaDh2kY51e/82
2Uvnfgx5s4/UoUndsefVDPEOoKryhKlUa2vZ6ciDFb6ytQqQoBtcYCOgiXQmwsA6
qWKcLvWGsfg3GoOj2tnzxb/h2DuPD0M/iqbMGYOFofEv8tBcggJaKTkIs1nvwuZH
7DJqvdLHU/o7IDcnOnUo9AEIh3qCDlyLA0AXD8pig4Nvm/kkTJ8ky6Usgdr0YvnK
eP/r3ozq70IXD6oelkfZEjCSIlZpxDJI+X9V3n6G+63bRlokqUVEVyNCuF+SGxGb
iQkh5OD7rK+uYRBUk/0FkqMLdWDYV5PsYIph4qQLeuxCf+FyJ2/BWqkNThM1x87F
uD5zQcpj0HxSXRPgb9MvX7zqr/lLROe6Ma0kjZoLCGTMNbSedVdLtA78O+XBTFtm
lLK/x5M8mo29c8kbz24HDPaHB02hg/TaZfBlA7B/06Bskc+SywjUV1oQx0g9mgXh
m4k/jXO9Yj9wRZ9LdWuhM1ktCSpvTpXrFRGk48X0K6aPw8EpiCsFQffPAc/0L5dt
z1QvG2L33S2tuiCrXl0Xe0TcT3pQV0jLrWGdnUGTx80OXS8ddqACKk6QUi5xQie3
xlwn+aGFs2fSfPwW4Sv2PXGMWLdG2TL8yM3Fvff52IYfY7Y2eETfTnbIqaOWUP61
r1FnnXmiW5CIAClEmriFX0RzSGcdDEFE4I2z7/QAxfGjZ0GXirdAPtQ7CA/KlIgs
yVwpbNUNDbR7YCViOw7p+xXRWbaESG7X1eSdnOxEg8UsJr8jKLu3RgcBI4sgXsv3
RgxdTrs8ti4hz4AH93CDrKOeRizpB0MEDD+qL0FH2Si0kMZBwTZ8hd+orHUOsy1L
/AKoqaeZ35Y7B8g/3Z9mBZkMkq3RXJbzf7QmjAFiM8puR4/8zM4tAdJKRs6Jn2DC
IDd7b2thCnkOkuOwY/fuvGCKrwGikB2cV00YPe/7DjcX1axxpMLIRduXzyJcTof1
HyxyjuzWfwH7Uv1g+pruIoQQYUV9jdkIf/VHSWzuvxZZqxx/OBt00F21Vo1zU7FY
LpEkxdsbDgtI+o0N5wbTw9TbJrtv+QmBAWn8nmSYPg3qthw3aHgZLI5hl4GVPRb5
e3E7ca0nnYLjb0m5fbln8DB4NpieRLQ1V4ubZigw2WIfrmPBwUJgBNmBx8px++it
7wF92u175wiz2LRwQ5nAk+d5SzfMGNjT74sI12QRk02/ZGTt9yM6gw6yFsofrKFG
j43X06WyJHCpxxztYnGateSS0Fakh8cdf4EC6oR6iyLsqFJH4/THRCLyjaFuiP+w
/Pjdx2oWia6YmFweUlzxF4cubyswXhuqqV90Hai1fBOafoaONQsquPulDvhr7XA5
7msjrHn0AakptAo6FWajQ8E6WPep4CJ1fNlJFmu03aWMtMzH/+m/rnefr9BZD0ra
+iveF6ZE23F1TCWgJEYKEUGOnJaZXGp/K1NmoK2+RypwJ7QKqUFYaQiTPZY/4XwS
k0OOoU7QR4zCYQ97IxGLhNUd+13/9dmXfi6WiyMlM0aR+LidTVgIb22QktGvVpXd
1eIFf5KJ8DwrsKfHgFpaFv1NlOdCmb0HSDmoax9/33UPRLWHHhHBK/lKvqQXwFKB
UcF9CYqXvsIu2BomMGJQKEBHfFda3tT9egvloG1nsG3sgv4rwFa19AVrbx5m6i7I
+Cl6EV3p87qQozIq3rRAS0PjVDICdwqdx7xkkfLCEznDiceTPEreU7pQkICxVbiK
V3Lxex77wFTmieZ1nQhHp8jX/VZWOmT6qY3ICmvo7bqKStQFTiKBOnUJQJ77Nqmy
Ygm3g+hr6lefkZTn9IU2X9CCocu2AmPTHtyh8HGIcQtseiqaB5TOHNu/3CUm6qiU
ExFr4RxCQYQwcjbBY0IfWkWlJJg0NN99Mhe7ewBFpEcPCBw9iGmAFM6yN3aeZwIY
toMgzKEjouaHWlRwMjD834ihPrL8hkb0w0oeKV+YRo4uXebMqVLx0XXlfYPwSi2N
VnYnny64iqlr6/z/TzhVA/PIrNq5pZ9hF4nz41ip36ttwr2phG+WZJTd5cceXiTB
1zYoZf08e/sCT/+75eXZc0cluadTczyifHeCAP6nPidOx8Ly8bJoMU203TaCpI6D
lLAYYmU+6I//DCjX9m6hQO7w6X5416elA1sdoHdpSICTyNYDWUYrByLmqj1vfu9s
NEyA9F/hr52TRsmPDz7V03i7FdJGu0uWbpb1DtM0vMmstlpb5r8ZRr1GyiZoVIS+
g/uVHPvAPtRcrUJ3Udf1h999w+RldErvneftA5AkxhrQpw9ae6c57iMT/0pt2gJ3
GF7tiu8PkD7jRRkSEcCq9Y+UdkMfNpvKaQH0uXelnJ7ycPZ4/bCf26KI7dBxJu8l
noH3Ze8APKoVYkz8XbGsY/yAIXJORx7J1M+Zp38wK0WoFnIxo5frv8GahipMg59w
qM5vBkMJhCFUhZLaDbERoV5TD5bXSp83wK0c7cnB6gn00HnhDv8wvLbJ9+JoPMTu
T9rxEG2xt4rF1zYCMPg9/aNPG1dD0mfE6NqniZJAUkHW6TH+lc3fx/stCYCHsW2q
pFaXOZvtUNiGi4i0VeqN6cOzXCEBKuzDUlThkwDs3teWGSkhYQ+W0BKham1oqLV7
6u+WdnEvgMXv8ZZqsPGD/oeKJ1pty0oZJ5zm/GqRACOOYGlWT0/ctGNVMlhyOj+v
Wb360YBmJL6EUOKuDBr+4e1sIVRLUpK5UOkOA83aj/lrBiyNQSnXNmxB3rQS8N73
lsyCB2u5FcfHVE4AK8rq3HMrQt5GgCwCsJ3k69Wxok9tB0qmkj7NBuyFDMCpqhFo
8/PiQrJv/mdd8YZDrFeHwqWypxYEoTQDCKBhEvSTRpT2r03w50mKqmEqIwLv7yVe
uTgJ5L4yzqMnlpzfcmNEDqyQVLAH61nwxDL0ZH2dwkFT3U0ckbcp59ScQ06xl01O
ocMnb1VyhKuuJMYel9nhTUb49xBWPmSljIaUdBUOKj6JKkTE/c7XyIKHkHzI30fD
NOaDcFisGROHDJIxX0d/WDJ0xZPgQHy2aptldja/UnoWW6V3cl4+QCYEGD7GLbp4
7X5xR3ctgoQ+vE/qNR69GoZvoz3VbyUjd+OuJZ4w3lV7VdL+Z/J4wUNIUn933XK4
8Le0B7Le5O6Tc9PDJowjNLjvGihopTh11+j7V4GK1VAJW78HVOnt06NNDmuL6eL4
rEwbd/HpS+QFT74rb4auZB83f00HkEtvTzvWolWZsIlu4V0074UiheFFaMzzuByx
ioNzmF9NVD3dMZIpqraMjSPS/o28udbZc5NndX/ovMbeCv2e4mA5s/gnU7eDFwoq
NGCwjnXAFIIZSejH2K6JNlOrc7oQ4O1gx2I/x3zHCR3/M+xfPZQxCW2XL089SqOz
ZyBeH8PgR6aZRPgkllLRBp5V4XpgMgM72nkQQ1VdP3C45s8Ov5lIAO4mfTpK4aSI
QatGviSyoEYSNrIpERc3Tr1mD/04e7B1BLBOmEY3IBBR39CD3XKHAFa3P0nf7zub
EAvJ6vR4uT5MoAPXAloe6fS4DRp4CXcoEVRBzg7DeYooH1D3kp57P2cT6JoKFoVC
p/Hk/A/n6lhuM5EMGmAr5ZPCqT1xlyw3sJ7qdFGSgxVkAv0fnRfqSuPWqyD8KBIM
72f+dc3jaYPmk6I8elC1UaCms2ykJX8cOgi4OwWoVuAZKpPz7VOU9+qr8nj+xGgg
nWQxOQ4XVrBtg15rTnjmN3RssnHH9iBKqy6cA9aIf67SilpnK9H2sij3W9ZfnikD
5p+qWBzk71v4GqwSi9DmD/Ko8Lcmp49VIfcB0QSS1tIO3RN1Mwb7tsT48Qi2o5kR
k1IqoLDCUfLe9TYweWHfX/AsZa+zsYby4o8ML3JHH7JRJCkW5Xj7DTxMRv4gzd+b
vXIrIOSwYy2zFVdjzM39HeKqrLQAuAS6wpBBIuXrg0lGvzFeouAWzUrPeAqi+X0z
VDlBgtoGUMR1SYMYJ7J3Dfmv2sNJgk2FJogB4+lcylw3ZqkCKZr0s3nSi7iKvHtN
SBftv3P+FGlvi4lXyjlNBQyNyc7P+HYziol6uuWVAvXxfOSeMCpN+DL8oYnXVKxc
UxKNj/QTZuygIFk+KQltw0Gaa8f/SmclDcKCwNmKJSdsiS/RrOIkJ2GxU/Ll+rmz
660rDtbUoPjON/upPvwUfy19clvBf9mdTyIOwRIQ1iDvWqijNQCV8NPrMuNPvbYf
BdpanaEZRFhQQdqra9hhkVQf0d9eErb1s1NNVO+1UvF3RUrp7sBF/pHdg7T4kcyk
Puy49DXG3QzTjwqzafYfhNHBL/7jqt/Yeapo+9lrz23RD6cRDevu4nvqND5KgNW4
0XcAIFjzaIlwMwaVbbuZn8W+4sO1eCnptKQC6G08T+KkItAAPqdLmS9Z9U44DY7f
TR8zkYIrFlDqQSjhH8U3eY7FS/UuWSYDSAZ15x0jfNqIcx9VVwlrV1YJ5jdnaGct
CmCkSYyQopnNJjQrgX2zceEUJts5ZNC3O2sNOK6A1Y4MEqA4KvmL0a9uPrFga7wV
7rWnKpHVpnNUkzXDdjuA6iC2PP2mcXyWckZIs1OOXde5v5zmB1uOxI0vYwDpWrMt
OQpi2mad8fmUru9FYwH32vzbKz7Zy60ir0EcdtXW9FN0fytWNzrToWMa0V4TRVIN
a4BQqwAb9tmHPGDgN+059Ofa9sq4/Z8YUW9vWNrReOkKPfJyxCauHECMkfUZLUYo
3IYzChXNkZDSr+bIjZ9kq8ZAYoPO4IReLX7hFUMtvzc7CSerStqJrPE/vhpFXJw5
sjAnFKiy+mkTHSGnRj4y2byEr5jod4FDLrF177F+XTFOKHAfKKQamqyNLb+2+NE5
GNFIDurpWFDX4lBZQFQkTi49bXywB+x9nSBIPV/osTXlgMC3rx+yDira87fG073J
nOGpaZEcbiYxcvEQ4DQzD/KNylAOWCM5NdBSOdYLWYyGR1srF8A6eGClyq2zoZ5N
SOXpPLnjtDfFyvab0qzcrCe9AAbtJe7uqHPGoo16NoALZpZK2l/djpcWIoGms44i
f/rgj8KBH0wiD/3fst4QOlC0L9NyM4LBULLDTbpViaFSZyn2rJ/lPX9v59+bdg9i
p/VK2dCAG695TAZWj+7+rqq2RLVZFM2gKglP+e5uyZyBPQhnBNmMswG58+FcO4as
MFbbaBzmFMOYlC1hHfTZqVhjFd4EukwZWok2h79Wz0WtG3ws3oXURGbw51C0eKmX
RoMlv1PZwWW3rY22SXR61m4v9rZHrEfYuxYuj/8xfYEFglpljasLF4GDYGCoEFEu
53caA7DDTdjdzADTLAnZ4M2gwOZi6gZzdPSenc7oAlhG2rEi/yi7wluK0qpHr3+H
ZZ8JDkjdLePwleQfVU+GjsCnMQ+sMXRCCfRxetnRgjv7jw+PxntsxJivKJi48ZHg
z8pt7u8kOHRmk/YoLQBCGPzOENWilT5PTlBjiwUWCF/IDM/L4vXBWyDsy7SQ4ngh
0mQ7OjaI36D99J1IfCUWgsrmFYiNRPPaS+xd7ijEA2R1uzsILjAy2gISGxarbsIC
WFWUw48VexpmgL0iF8dXl6qeba9efKvj94t4zINplTdnFQ2Gp/tsoVX7E1LK0lSY
ciWAiZlS9OKViiVqxxx6soJyrG+ZAZBND7ZBnQG/YLh0JxBvt5Iii46I4N+SjE8O
aG120HM7N9jSaYNNbJiCazPJze2FGwrqyuIwjjvvreEzrXgzDBFpGqXJb1e4x5SE
GnWtaCjbbITC/3vaLxsLHi6lXYduEsuVLtqGbJ49VarSIwI1ML+d+RPCneHNj+Gb
Z0a47boRCZZGI3u8DxYWAM7QhMw3EKUWbU4DhmnT6SN5xdZxMt1IAMSLQME/LTge
LyzrPUDk5cKmkD9/1+mmuQc+IZL2xerpLx/aZqDP7O+w0Lc/ezDOS2J+QQ4HXenA
8LmH6W1ZREHkFYzU/sfc3PoNL0Ts140PC8v1xdDqqFqXPSaxv9WZ1cSnYxdzHuLX
10x2pPRAZWkEuUArx25quVlrhkglF/zK/aYXRFZI1nJ6ZQYY8WDj36W1p1vnXuc4
Ovo26akz0Hf3wDm8JEcX2WHE/GJrhhA0c21C+UJrQFp0l6R0Gbwa8Vd30Ufvntk8
9R5UqvPqAmLT+1vbcW2Shxj0pDmVXuf7x54kc589DYjuwyUyKcZYp6U7lGoXfz/w
slLQrzYVZw+M/Nrxp7n8tgBiELPoaZT08dPMD247tKKB77QVbiKrfK+lRguSLJKz
is9IOXtll2sr0xNhMZu5MKzfpkuxQLSECmWIReGIB5LPZB0qGecJbJ18jw+y6e4o
PUcWc9eJWI7lYN1n2vxZ+8csst1zqdJQfIZFHlOxuW/Iwg88vsWxcLxT7WBN5yn6
KmEONEFZJCWzTZ9GCzCe7wHJWxC3OTPAQjnmeHY9MR7N0AUEuE9O/KWTScutl+uX
+VxQKFCFrT7bPfaQnxzPqevPhpVeDu4CzQtaDLDo+EureQsbirMBpDQHe/gsfsNw
Mbii8fi2Brmm2Ts3xMHPDq39JT4AH+Ehu57elCa/Kjw6a6T8VMr9ksz1q3blW91z
dxLPOKV304yhZ5oj6WOlVfkjWk9XfEuqnO4k9paLWXNS68MiB5A00RBQ/q/ictZU
J8f4SfFqH8XziZ9Plxl4nC93mwZLU7sb91pKCs0abyw9Lbxk8WX2Zk7HW64HhuEw
Gk1bjpAsWJV/dbmLruHgrVjnf5DV/d0fnAFytLMG2xmrJ/wzwSZ846nT2WPru+Em
DcBJy6mHS/lP5tmsbVWpE5c7uavc3BDf5Enb1CREynOm/x30Nn6bx2AKSLpwNC7S
xTTVOsLccY+TBZ4Z7dEOF4NxjvE2d25V544sYlml4OFC+NO0YoaN46xo63sFFhLW
FTxfYSd5btAh2qvZzabVXGfkUe2YrLTTKFIL3LZtUTyTqTLa3W5Rj59qw3LnDtZJ
dtGwCaXV1viqeVaPcZstrzKDq7xF90qwneeHsRbc+Jmi84JyenNnedB+Hk3J9idE
nbKNxZYBnikiokGC7k8zW9C79smMb5S36GlICgJKcDkc3/wZb9OQn/H0x51BPKlb
OtZ6oyZtwsAp0thrP8n87++Kn/w+GVbBptmdqYHctDpY8AhplPdflawNfRQBB89U
L5vYkGd+iL4DH2xbQlK+FMJoZd6lbvtbPt0j17TTJrwEaNyi+w0kzRYkoIYUJ8s0
F5FamBSTnUqakAcYJtTWHr06k7uSwUUs5LoGj9Rc3jxwT8NmkoHMzXkdZBG5DHPc
YqvtRYdgdw0vV4rCR/qZjyt8A7QnRGD9Zgo93qQZ0K6xX2ZwPYdMMtBfJkByLVaQ
Y7SfgL76lc4ne+agx468Bq+wMolyd7Zeu853HflmIbnUXPW1+93hcZ9c5d6s0+41
qDwNmoH827/4fb2Vw/e1LPowN4gzwwrhAoXUIxIx32S958Kkf4yeL3TXMhpvZ+wj
AYboIQpGquY1+ef/dO0bLScaG24VEbZRVHPyslYNyGohFqpo+J1SCy8bpjGGdEZM
abcv3HR+EsCi+G7wg2rstiGesui/f6dRf+/rke3GcT4DHLXI037q+HSJ9hIm+BvZ
SfViO2vpfn5MkYhevBXc08jcDdsDnx/P/YTHw/Gde2s2TZak06fSw71ANGWcAuFs
PB98Pik4Sa+meGsBOT89NENe3Bg7th5n0UDVHhehK8coXADHWLwF6rw+mrSEcjN/
GEoe4tsy1Q43xaOfdnSmCWCDx+4oFtGzMBhF91qhb7XWtv/jb3qJRLga5sui0dDW
dbXtbG/SCm5dUz3qH9xMbPKVCXECY1d0oA7LqB8UQYxVIb/avJFAmzWfMwG/5nFc
uP+ImFVOkx14boaAZ0zxVllbHTRZQpTKkp24Ls1FxowB+cpLJ7PfpnLpiyaigUmG
SPlFj4mBztdqpEoAS6ekpzTGCbuqpU6mCq1fHn3cyUxdS8++HW93gmZyGh4/Q/Hk
5HU5dqpBOP58PZTxmLym0ksXalQE6x0zkY2SgjhzA6fQ7cNHpjIILQgWfOCy/XHs
6tvo7Q+Y1wk3XdKaLV0ZDSGgpMNFW3lZwlADHxIJq2OPYGUlNp7eap8brHJkbF2+
cGieyqdjVX2LnRPQNBk1Bh2axhFJgT9siofEySCnO2opARgAI/bGmyjTbQH9Ghif
+16mtVsN/k0MmGnEAgO7aN42+iU13gQyG7M7n5nvDFMtwhxoMMkiAqUG/DFveIQx
/1n2xAF7ZQI/3FvfPnwvFNG6nRCOAaQsNstU8rMsKI9oepN0z6dajkWZyGuurshj
QgsaLo8gYuNFwtQ9Z7uJqXYBt4gpj49L2ORjBx9tJz4LDeQIGexAIlrCooMP+pCM
wfahyPnsoDVjSjo0yftq8RuBwgOrpiYs5nnDGYiFOeB2lISM3CWaT6P3scTbcv1+
jr2Fwgrk2CNDhGGTwyjzeT0NUVNrz7edkZBg3YMHfvf9s8D3GVvGEMWpfCXGXJMH
XRkqCRiH4CQzc7pnNE54mQnkac63CnbSqlIgbf+65dgWa+ujtt7hHqqUei85W2im
e383jLajH4wPRF39NNGKrWy17Tqgc8SGmVCZt+2m3LcJKqdJZtUu/i+GYq6GuLn0
I1pnq19nCFurvzG4UHdYSsNdF5yFGkQWcQBJFlBJ4BrjgaDUOIlu+6EJkAIy3l2l
EVEbINo0rbG2vQgOkjIdozaAzacKP/vhyw0iB4rkjiIG5Jvn1vVeSKvyrQlRVJTX
ah9s2WE9bXBOV+1Y0nKv363yHGDzewkdOrm3JTH6Cj3yG8ztwfBmhb50G2VxRjF4
0UoIxGSDKatDFDbPxc7tMX84FrNyJimHfrWQ4mHgj8G3El5RdCBXr4m8HkpcfPBb
wpLFvljVBEtYYwd6a9dre5Pia7LozcDTIuxlqm8LHKgvc/Q+Sby3l+2mTRHM2ano
VDjiuIpEIWAIrJV8AyS6yxPu/EDG8kPu4+SJjnaBtj1FuprMTnq37+PkQCcvnjyk
GQoFfc0/ASIdhRnD7fWOxg/hd8GS/ABePXauIicxEUGaUU/zWjJ13Pzw6525pXM8
c89rL0Jjf2Z3uw1/z4giCflzLbHjv01D1GwgRZIpzf4LNbDrA93E2x+alnex5WlR
lClto8+89XuxwpJCnrFuY2qEcqkWcjozTcjaTElKBf5bxIknQNeRmMAqiCWoxRfw
dGe8MYySqBSVzEkUo3Mh+aub0aoULnmHA8yKTPmaWQEbDdHcbtILhCEfal57Hxuk
iUrOqkpo4EU8GHEVQn4A6krP4YNtM+JoVSTOSN0osDyMeN63zYxoWfM05SAuldII
Bx2H0pPj/60ebYNpNifMYTro0/qCLt+0gQgdtDAK2V12Z4hsMdht6kL1AZ+iCYoM
/HzoK8k1Zf82QRLsxI67iBy6rdM4APgs8FnVkDFySjM/vCfxhMtSjicIguKVeCW9
oP2cmvu9QfShLF54gZe3G8/sK5d+H80vhb/JHY6lgQUdphpbAqAWfpx5Th+800Cv
cnaR7xQNDHFFUj0OZ4x+wVG5xk/SUwqqc8LmHay1+dmIMjp4bDojdWy3/yjzV5F6
2Mo2f9Ns14t8SfrnibPZT6l6OPrVV4htdXf4uModgt59YzjZ8f4Ak5so+MlF3SwF
YpEvZyffQzMrAbRTrO9g2gPYdwfbH77Syt8bwKMujP28pF5k1IAyqIdWEr3T0Rvy
cJu7/9b4xPG8HcDeGo//wm4WF/zWyLVel9IkksKciF6A1QplwLdnzXbKUrO1YbFJ
XYlD4ypyMkjr4YzfmjOGlON7sXm6ToaZw+TrN+lT3TijnEulFm41dR417nFBdOBS
2PZ+3Ayv/iaBVX4InqsTl01XsB0dHv1k/z3SogiP3msqcJcpPzZvGBOITJYW5EW5
8V2qb34+c1xAJ4mWP/xUhoxicF1gVzk0Fu3IckykKX9ZV9DgpHhehxRx406WhxXR
2t9MA6mjCzxfQgmPDH/089t74C4FblGJ8/jq5FU85f5KDdFbScfVKElqQBV4MzlO
uo08PBsqF8OCafrp+Ol+Vgg/+dFIZha7FPOwTe/ySXr6ZQx9KLIEc2kRj4pOK9uT
wztieqg02KbyiwYAdqYqwoLU9epQZGJjnYkix471RiZ4v59Zb7ytk6WKXCRTo72v
iqfxnx2nnrfvBpchOzgqCCopsC0CoPikw2HxKhRMZKXW6fgg+607T6op9pIbUP5n
Nyh6xe2NRodtx86iUGScbjw3fosMcGIASBdxIXqXHAhaqHZLTWI4G3p4M4WnD00K
BXRLwys3JVIjVDGPyVNUx4UYDroCmvwUcisEpd/Z4Pp7T2yr6NuwCjkExznBqRJj
ZdtKoroihBnF3GJq+FHjOpsiqthQmwD5g9UKGoXDVg94TmhSiT97/McV5E7nSc2x
LByM76AE9ROpfhg7u1ZcRk8OWxWHJN9eqgVchfCIUU8g0BxPjAtYP/XNrMmpRFMV
desDYeC5Rf9goGVqHbMS+SCp9oeQbM2cax8zxjorzN96YiaPJWGqaN8FSxnLc8Uw
KnSSWmK4rSO3KxAh+PbBff0G34iXhUNkzcyNvLGaAaSWof5Tr9h3WKi1KoCL4SCx
Z7JrpCq8s1sHEc1YSslCFY3Egc/zkVtI0/mpqR/HNeeIPfPFM1jrNhKILpu3ylyy
PQYUrlL15av2xHJ6MPy19bqeFaL81URFDpsREj84yNVRHPLxe0eZ5PWjh5zjB79S
m3ttBh0l3bEfa8eknmt2PEF0nUoIcSKayIeh/vN/z0L6hwT+J6qBCjAkJ6I7Dtoi
aJgNMiuImdRyJJ9Yc4Yrej/vXqJ+ers7qHQ2y1ThlCBqbklHYWxeCx1peLJ0wpDV
lynkdT7O+rWTdxhoDa7zGy+zprbijJmuTKRjd/Fd3IpyaRZZYvXoWJ0og0qNM90F
YLfouGWoxyXIi7GF+1V3plx16bqdvCbC05O8/2AU3bT8r4KJKKZVih3rL8QE9QS0
+Yh97WQ2M/0wiZ11CXG319BPvl0N45pcm+4g6m2/JTj12HgwIMe7j8dPmvj/bb+j
RLMgoFY+gFOspjMFaS3bXvtYSNwSHe1djpTTxA2kC02nE8Ekoiokc7sKJYUx8lAA
TqoLPu05lIw21NrOnLDM/e9ltLZ/L7flKfQU8JnbpTF3ryrwuRTUA1US+8/fguEW
75xvtWloa3lENGeWxzsmPQuFOd1TvokZPBAVCkPwfaBkGqUZfev1QnYgx/OtG896
woc0/BidSuHNCgi3MoRRrmjhGk4iSEhJFd3mBv4RPVX8usd4oKuVGvyt4Vp60qVI
wbiNNPOWSJNQmLzD7hfwk0lJNVBk3P1E6IezJDOQ/1/zNbiTuV7B1KwP8hfkqCbh
16Dr/TDXuR/9JKhDHpfrkM6qmmQpjcQUvlB6r7lheo2a39WfTeeZmG4i8GI3k5tB
vg52TaYRX5NEfDSEIopGqW0o+AhajBh6QO3Xy83FQLPR8zAL383j5lA7tdZjXAO4
u4pyBnmZNx3aKoBT+e1vHmuyTDszxWPQ5cvbx2luDDhK/e1MBUD/iyIHuUkLJ+b3
a6SQPHQ4LKrhfZjo2yMnEYtxPkKNJRlJ9STmBRKh1UXANJnUxmiugLt4HVib3t24
yd8tnbEWiKNokdE7AmfmQUlyKNuzfYEohjknGGMQn99G/TJdg3ucCknsT5sLe6Js
LqmdeIVuoySRsAJywIR94D538iZWRm0sydqoZav+GV9R1/4jUcXe+cBjOfsVtThw
rE3TR+I+a7e3XfD9ASWTGnYRpRB2g9WovGwJ3KqHsGywa+Xp94rM8x/YvvkWMqY2
5F3HAfvuaF/GLlS0yNJhrzTTDSeQTO5jA9RgUza3n5oJO1/VKdEB4eQfB9UYw1iD
wvj4kQ28zCooFa3bYbQB3Cv2iWoIdHWbEiGV1h3kZWcLmoRGQLOPJ8cx6MZwpFo+
eytyaYU4tdM+lBs/B9dsQBNg/CVbVbstKYI6VukSu/IkZjHuNgTfKd35mC24giSS
dPK2eWMQqrwu6RskdHDu6AjgkIRHHlo8XUYt5LRc7AqtHbaC/k8Hc+R26gsHaIt/
t6miqjYABloQ2i1pKy+fbVbJD0vgD6r3Qc6NDp0VFaJevLQa454SfLXVdvxZl6D6
ZWcLc3WqCFWshtrq2Cx6EHuys54ns5GdIUUdJKfvg9pwDVz41kVeamO2W0xVq0di
bbwmISY5Bwa52fKHgXHKKB3nLyEWN9DPk03sko5ujN9nza5Zl302UpOea+v6Iw9d
bfglkAkeqUcDSXIIGUpTwJm/7jp2I5wSJPi15dGQzGbCsfKEm06az9dZWstKVKzy
prFoy3NeKnr5rGC7hapSxIXbn0uvfHPrvXmqgJdE+EawatrIG6DvMUGPWBJjMhZu
3ku7ubWfCp0v2BqwUnSCZ3CcHRcVu5W7/tIvdBnkgZqu4eXlcXtCgnAd9QY3/jaN
KY+wUoa4X2O+ewph5lEGWdGGOvH3WEj2Ly4H5RBqeV24K8zNHxSPx3BCpNqM73yT
0nl+cIEtlbb3La5P/TwTqUf/l6uQ2IyHSsaDM6cRdG3PGa3Xno7nJ7zx+jqmpP8i
k20YzbPmIwuqZljafcq8gCnshJZcVfrDGvam6CJ62sIqyu+W1ZppB1gXgUCLHiHT
r47B8eUyTlbOpu0pO13Vji0/xarhQOUt5Pp6n7U74U0i6mzgg2zKB8cn1U14iqRh
zQTkF7eqw3pDDErczIyuDwGVRicv9QEIl9/K5t5p6BiiKcCCxbQpbPRMCCAEJahM
TnLGnsrlwsk4MbtE8GCOe0HqkaA3z+KNzGS2Ho+hNsFUjmGd5JtnRHrJNkciMWgX
/nDC27zu+JCETU8RRF1Zdm3wzb9P6rhNqJ/VyV5HLQoN/czybtLBjpgv+221ilpT
X8S7xNsJVByQe+xgidEFG9pIyCd0n6ZX39GhJCy40dtv0Qt7L09W8208aniXX4Qb
a4aPATIVoOAOGlkagzdKaH4+q2n0cj4OkF1GdKUUzIMrCPhwF8aCm48Xm6OqGaOa
YJtfjWEbUCD6HaEUrOONxrQNYDZ6kJOdJsS+T26nbGEvgD3jdJgLlqcogfbn9i/U
1FM9BiBaEepiZLxk00m5y8cqtm8fVuKGtZ6rmwzQ12c+VPysyPoGxiCySohpQHMY
Aj9MfQsGMAcTVs64GoS9ttCnMt06APwTyIu30lMjIPZNXMwB2Qcxw0Y9aMN8xnOv
JNEsJ0ZDFTSfcmk+eZmcn/idw2j0VvfobUKofPQUxmd/JHZq9bkzaWd9r+7BYDFP
g9yVUTPYazroR4pYsPxsfc0ANJZIqXbDZSzx+txpORroqH9fJqeCWrxXpuVxBBLP
IfkcgB592/a4A59T0Ef7+nEk2vp+e2BXK6Vy3+adWQKYbWePEXrGi00cOYiOu3xo
PPS0/aIiB+oPTpcjxlcf+A7Wri7onO+KwySWkID7hI1Qss/HHKNg3EreiIEHRMay
P+IcbWddLT4AbyFgyxDx2LZNofE6w8737atlHFgu8awo1dIELZR3+fhuKtR21OGl
KbXMHWKFJWtOATx+2sFZf8tNUMn0oTW2mSNIk09fNgpdwP2/Cxn0CiD4E08Y5Bl8
u4O1Pb7gHaAgQmEOyfZADvB8FB56FGWqIBJJaBjxawTsSFjXlnTwuXFkixq+76yv
0u5hf/8UQPfd94wDVPZ/J67S0zh/iQHDwGkF2Le6ZtDofumJf90/P98gZZkgy/0v
PB9vZdGFYB9sJeDKmfxkDy0pBMHDCG0QYHZUP4AYWvfWrl/5l43iaOhAUPpvwL4Z
PRYszay3m5lPIHK7o/ouVvjpCMGV54/uvCTf31i6/QgUhhYMRdtIVlRwyeIB0VuO
/ZcdgiHJf2IgxoGjcJfX4F54pN6VVnIfsn6EP8lBBptYnzankkpdNthzoz9S/r3f
bW1TdUlp4tNUnKcMCB7beY7w7Y7HisovKocJ3y2GFAdLYH2zognA69Y5ewS215R/
YEBWO+o0LwJZxLQy6zdsbfZnoT9/LVk5a2g2FxGn366obCAoAZ9Z3HgC+jUYVzwA
kJ+OrNOGJJZQZZTwXZLP49IATmOc42XgCUa8EhCYn104lakkqOv9NR7RB36+3xG8
HokfcKOWAbDlN9qdaVIfa9iJblsyUWR9YVY9HaSpp88ISur8bnxWYJ0r/Ple9BU/
Ierm7MkZI257mC5S9TIoiiZDVYWFtxo9BfT0afQYaRd7IlEaCEyTuFBR1VCXFpl1
43KH2aeAdpysWCuAfiq3ip6YWCaMh0MW5cr70XjOq5S8a5vHCkYamNdoe7ESqbvq
bE003PSpF8h7bbXqgcDZLGvmpKZEoSHSOa9T+XqBVO2Z3ZNbPDnorHIbI09GfiXh
mZdPm4X8lbie1NeJND3+TVBlOiHTORzaYXdKivsG31jW3lzYmkHIORwG7jBRTLHj
M4vh7PNqrhlomW8YWok36mtYP4398/55XzASiwYTl0rGArVBL+zBI6DM+t/pjRFb
EZVts5vCKyN6fvGiEqal/v6WXMkAtYF6o7VgHAT1LbltGtGM2nYBBthaXHvR0/2F
5nkoz85hSbPWkNjy6+hvxjsn20BNVeBe9Yx1TVNtXt6ka4PSPeCxbKXt9CMI5a3y
ILLlFSzKpYSI2XiyvTyWYBRA7RAW/IadUqpiZNc5dItsOeHLasavvu2eHJijnE6R
2OfpsassDOMCJNbP40CBUNERVEs+bGHnSq0du5QF68aSbA6P/KE1U5pp6Vh4U2fP
9OEqhNg0PDZ45NWL+0K3wuEqcQbAWYph5OO8LwOZ1/SP+8pZUIt04ejvOBbzZDJT
acKBRu2b+NpXbCf7EREjb1smQYfTa5ksZMWKbnMybnf174BiC64Cbl6KMqT0xb3a
MqO/p/250ZIhFk7AuSHREXIOeEwVD3O2tPt2MD1O8Ov29PftcG2zYE85KjxsH6WF
LxAF3W6eEOA4ufYHT0PKnfQqi0z35eDI7CIkWc/klu8wAZHU4zEnFcwsfFWIGDqi
11VrTTUpf538QOebyYdhATgGBHkH5qB7M8FnpdGuIyAH1v8vJFRGxvH09HLp/bVF
2MvXfInor5mf9CQMhwdKsGgkSVTVzaKlmBsEC4ZLwwm5N5Vxq3P10FdvNdfVyfkh
S1+97dKGPTUq/UyhUxZfnRawo75b5gL97S3zu7ygxmDCpV1/JxPcLszusNIU3wAH
QDWcjSB6HfKkgSVj2ysZLK931r+c17K1WT9Bi4cDN7ezcsOeR8ooAjY8WorRAeD7
mcu/qYvJuatQWI//aKN+SDWD0oc5z0/uLTyKoM60eUD4zDDoK36nsA7j0eH085TK
vIhWRXaWpqPsEH5cKYlVfhR55Eio01nGo5alzvxjQOL8UkhCLH/t8ya1pVwriIfK
gZDNfR9gY/e4wPA55shui5OE1jjuqNRZjT3IXAtILyWK6mW0uFXfB4TLYl83msQB
3trv14hMSioEfETQNbcNBX82YOOj6IGeqtkjXfjutafTWTBegrAwyx5i/jnBKIoj
NDobRUoSX9YMDGP/bg/W1qX8F9HTZJpQhempuzKm28EOqNMTD6gFbFcdy6eN3pDO
RAWC4UCtfEOsyzQuRyHusjcKjfxNtNdsO826/RaJAWtJuA7Judtmee38NzdFx7ys
4Gbn1TTuPdlqR5OglN7WAyrdwkxcCnORLmOA2kr9DhwLmKjkPvZGPVFcD5GsG6VJ
PaeSfq26ODr2p8CkTPbQn1FnQC320cTRmyXXL8zcRQ6IM1pZSElB1NnNfXnucL6f
a7ZQZxx3HW5UjzCeMT8CkY6O2uARqO7ZCqiBCx67oApKh/6vf2DTRbz+7Hl6NUv+
cJHKC6gQ0zjidIdvkI4iHFgBHVr5xXMwKifl64jJ/7pLl0PaK0zllJimouEMkHdF
eu3o7SKIucXwl4q9DF0rw1Vaofwtu1WTCbiW5+sPu+7Ku08rS3IScfiDulOUd/kB
NvPTaOjYWNIuqEe5ZhFW71Sye9wUUjqXApG2fVNFM/FXyMQwq3zWj22bxWGJkgHh
6RTsB7G9df+gvaB/8JP/qhZFfL6rwHz7xZuLQru2UmpPc+UJqHEsQMJsIhoTlVT9
GX5CPHFQpmlo2aNtLJSWRV8HEfCzNXZbZzL53dKdqKXPQ3deNGrqcLIJ8tVWJRI2
FTgorxN0AU1a0//LA6NdEvFX+qJiA/AE/t89HL84rf0Y8m66kzokrGxljPgdhL+Q
8+2ef07++NwhNIaIt/V4Dz+oIOzecQdRTb+Ed1OdJao4x1g6c9q7hP7gZwAuFdvM
NAcvGVsc/YJ9L+CukIQ3Gs0XxkmfWewiK3qV2f9gCg0jLnXJuF3FJfUfm/iax5yk
jzlffdKZMNcfbiGDTABMtyE5N+45pw9GjsBPCg15K3XQ8lEXF/++Bclja5nufHRS
C8MtAVXreSF2DrMxWFZHBAmFlLA6RnqK4jXNDu4geo72CSnRya6hBWdxGc/YZPYR
J7DVrI4ZmGqmf9LMoEzS7EyI0WbnnqqtXES2AKZGmfivkQoKKYBhwrLtt1EILp0J
6dbT/KkbwVayC2Fm7q0ILd1eCy1wWZJn2qvj9KhgIDmkaDLniJYd3DCA/Ynyo/xe
iDrL1xC5TmTjvXb1zwdhB0BED99oxTtiHSnVw2BSMq1i+C1PX6KfsgrPMPzDiAwM
Ze2dryERoTm//xNo+CYUJsJTL0U/CQG5wnuODkMaR8qNKXQyyllu7RH+7PIYLA+h
5aKlaJQZD5g+RQVDI1pDVSb0iqJWF7gJ+tjRpxa1qev9HF9Sm1+uV5jGdbw/eYNt
8ldNQ3Pn6VGbKWB6xPB0nAlKeWr6wc+wym9lFm1rQNtqxjuk+4HsIrCMdZ/fFzfe
yWFHXUzp8HA00SP0gEvhK92jW4UDJxTS369mcXAoZJkIMmVWrT3odMo6W77qr5LX
BUAJ7v5S9KRT8rWzLcO0UggYskN/h6KYkxOtFD8c8+buHIGFoezUxJJtVUN0C/7n
efQV0qpe4DUXxW9Nha9dZyYgDQqo1P93T0yn3FtFXOldRWWIigkE0C1WjXPuHD5v
yye6ysREoYXMaRdGv337nfcssxht7xGjh2fMeClNcfYo3yHctnnua3/8hQNgbBKp
0RyTfwTHFxeKFr3qQ5kkKt51gn4ahNI8cnBlbXPJ6crQmg7FWFaMfTXUxCc+x1RX
aoi9mQbJ2dmwoJQ9ZJhZBc53xLcm1LgpIQA4B2SPxIUyRo+b/H0vKdMxpBC1e6lg
PsxhiXBdwXv4/JxoVULqzh9XPnGj6132PgcU8coMFZej7SIlR8gGZumdPcGNNiGN
a58sl/3yF2XixEh10mkDrKkMQtrjpj0ZdKMI7uagr63/g2BqoPj9fhXTTJY88nDy
GQAfVAqJGpE9aEn8YlSJwxpoEsP9ClW4+2trDYDoastmuYsWBCzh6yGLQpu70z5M
zZ1Sl7DDnWcmeIFKvFVcAnc8iarbVc4kY4CoFml2hpBnn9x9eKFnRPdKQEw2f4oj
vhUbO5bNgl7gFbrEIzGAyyPnleJ60Wtq3j9m3E7cE1Ghy3winIDVfhGXhFnKUq/L
JnOUUbNj7VpOwfFLHQoe18HiRzvghghby/SI/uRt+NtT49F4ICH3ErxPi0cPB8bI
ujkYHRNMZzFjZb++kmqiDE4UGOcxbuAG5y4kUK+v5rFCqT26VR3zWgTI9+57wegv
vBFmjoJxhtQbLEtDc+L0/Cp6ltDbzMuoY2/vNiVYSkoX1E3RPpkU0zbh3nL6mrT8
SSgZ6Qh720qQaIvvW2GqEUuswlk1MOWU35BhdDzSHAe8uL6OJfDj/gTItcu2h77x
cVH41v4vmM8iXHzkcLS10WCUKJEaXgC+flHWHe1akU+KOdQZa3W363EKsUVths5I
am5oYpyNsR5tZk+Q+40/poZvhkAZykFOzWwH+oynMmkMbCqNhiSm1Byt77Y/B/o5
m6oNMxFeRQrlEhl/N7XmIYcxd5QsI29ZkYU7jzOYsS2UQrnuTWwn9Wtj2XpMT3Q2
ahmNY2g3CxM5uHIcEwByrI3AFx02y+2rqsgSOY1Lv45K9zMv+WasphuhxmKYJl+W
tkPQeWXlG8xkeRduNShbwPhlD7dx7IyKF3wV13phs0OBcHgxeFpfbviS+r1XlBgN
C3WgzkM+vDDgW5MURwkl8WU+WrfpRqv3O87IfTJiH8aPBCHtQiwafPvkr1k4sht3
Ss+b8elcRcCK36c+R0hUHmG90Fbl9qDT8Ah+cY5j/LxfKr8Qhhn929JBjc4byEEe
SW41DVixf3mmIdx3VrZYlS8/tZF6xObICJJCDEDSr/3xEEUgdAzvV4TKKUvf8wt7
Im2PTY4bN2907lG/+IszNPJciPyXThiEP4yPXqttipPBlZYudDOyRpCf8qrc/xiG
imI4nulVv4ccB/3wId8PFup5fWrhXaORqVDNMdEC2iJE7iX1A5xbHQNOFDhZjHEw
i9qkeuRu1T64V5jtJFKzbRQZqpIPJoNLsSiObb1kJlGblsiBcEULRliBCzzUsRVV
9jIUt1gvCPWaGiCd4vSBVCLWNW1rgeqycRTsPVwzpslZZUmgX38uY8U0DGVFHz2x
ZKo7mF9V4etwlmYOR69wrU+ToHR7/hPfk2jOkNz4XD5Mf4Cmae6X93Iptg28VirF
JR8XbmJSt8jgREJU3+hImYjcULuij0AcGib1KqDI5sr0ih+CiQMFrcu92kKWBKjG
n+8KIRlKbLzqfeGFGny0rIlpIg3W77JqIQwXuRjx5gJ7Dd56jtC114+xwRcktqaj
7K75TtW+Uxj65BSqs/drFTt0EpzklfBWLhEzCVBLqJWm6UfwSiRfnYjpBzPrjv4Y
w6sxxGo9oe0zqNXk3Mnbvu1hmkR2QWgNhRfIsx1jVwVHSvPB6Ty4goadw4cmv3ff
2gl4xhBqSHxYXi963xmHG4CF+ttKH83wJqlHy38ZtIND7/oJYAMEjzBEOwtQQrmu
PdK9Khw+tyjiL6EWWC97D7RAXWHqlGRhbvSVhqqVNZAM9HPioyTW82gujPjQnIet
cJMJi/nwoWFt/mSutySCaotqSm65rowYdkfBdboKptVgzTejwCUPF9p4unaedJlH
TpovgvNrUauPkRhtUq35qSLQhyLiV7KzckNDJoSyrhEHuPLqmw0G89sbxsQOOscD
et5ojCxe2887DoQ3Z4X0HDlij+I2QXPZeQc5i1BBKA6zI3dRnbOOS2ceAnsrWkLT
JqOWMOHwtmPibrTwPXMHoHtEsqoinN2QibDvnk+wHok4ASF9bdpr7Hmw7QJ6ip4a
cFg2Pu3BEVCpDd3soIPZ4thdF41+c9sGP6k0uRv9EqvGlotxXlgDee4ccMidPknO
VTr9OqsJ/Jn+kph1HDHNUMC3JJbhfzMZ0ZkAV7kCm4iLcMpmjE/NCf3isYxm+VbK
Ui9tlHRi9DEVn3XsQJl/DcPprS7Lz5EKcVE89D+uytVxeglb0o7fvL5HYXLvwkpb
p9BVlaqlXWfey/4VswJ+tUxpJure06Nyhxmg6NEMmXDSAl72P4qq0ja3n4mOawaM
6C8ySkCf1Qw8mLs1xoKehSi8Zs543VwOcaZmFQ9Y1JvbizO+rBg/JSFTUi+t6aw5
xXk1RAI+nclExR8kFmmipyxig1M96A5MHEFCLSu/ml+wD0bg/1Mh+VNIyrUQ+QNh
ty/2X5eiXVGVUIgMkjl5NPQ9d/ltYuMHJ86IffZJytpVJkKhYDnO7Y5Pdh7oa57r
tkVKeYCuXhqb07gYVRw3zcnaPuXh3LPhwyvQi2KRbc2sEecJS+pyKHOzHq0oyVHW
mNexp7MJieTHaDY4XkeBiaePdHTunzn1ttqHdq8nxQXwwJvlfhO2LoHxUEkOzEvx
/Fpxut+Jw0/QSJgB4+/hPw8iCaF4ZWKLrOaS+Qpd9ztg+aKlVGsfEl0Ndct7+sBh
aIEN+hEXL+QUBBwBza5GlkRS249q7shispQnhGjxFqsHjIzwk0Ifbnit3XI9d8um
l0r88LE1PUdIRzjnOa3MFo2TCaQnK57+WMs6tMfWLTGa3pXduVigNaP3JrV01L+o
L22H1Ube6amSewH+Rz8YWDa4d19fXvHBl/9ZtRitGvoqGpBvDxIUwaAmbYALYr5S
bwQ1LlI7xAvtkGf2DAjJYywZ9QmyoSi2BGg+QcShnELRlblzbLCaNeaHcxeqL4Dw
nEbDxyLUcroRpOpGolPcA4HMwrPGSgEqFI3CztiN+vFh2XFWUuZF1bBF5tnsAFOW
GT2uD3CQlD4CB2upvM2IMhbP26TgUpp2oFJR/apO/heu080P25Rzlt061AQmCFb4
ONYj+S4Bx9FAx2QFJ9KnwkZmjFXMGz25OjqrVlkA/yvIKdkd/fP8ia7S990ZfVjy
GwPyzz1B5PJX5/vPHZmv8KCPH+zh3GLsb+gMZfOYV/zzSKTmdT51Azrr3mnaMmQ4
MT+LxhXAWd9sWFUdoBTIrsQop0FkLjUo4iukQeICIjAwDQrPxVSlgwTNL4BW+BS+
h19scDYlwEi6ZGGZYRsilPAKlHAgyscEiSR9DyDF/NmpZot1bZ6HBi1dFGDd2R8B
EgUgwBdDDyBNTCCSc8f7E5C6cmBI9cIAe7vhu5EUkyVCAQhW8iGIRHsNUGyC3Yw+
ZACi8mWGSvS5X+QQQW+1wDeIKr2rFXqPrzxm4J8aSl93jloCV8ibAfq9IFjYN9mG
01BTyzFraf6WzgbDZ3MprCqZA7qQtXJqRhbdT1VAsMbgPZO9r8h/zgM4jaDXjQ8x
6dXywI146EDL1q2t5yfSxIt2S4iTkhL2zvx4OUukBBIGVRet6f1fLxgycv7PkuGA
yN8sfoXGlUA+pjUYoZs/I8xJknX/Iw5jfsId9b4HxeTkwKeNTVQUR6xHXWeGmnYj
jjPd61RX/0hq6Ssjt8ex1fofv9DeT2nm/1Yp6qrORS1m7r2mGiiAIgGWg2WVR1NG
LM3ukWHMPV/Jh8Kv80dyW/DdVw1s9RGOufaCchy4OhTGMpI8w9mJYru7KhESWBI9
nDsLhIvJLeq60NHMjXOXNZUz26IYtW8/EyJgvSN/i6sUQQ+H8gAGDLO5jE76bTeI
Y8x6Yr6Eb0w0jUNFOPrm/VAc/KVnAlKUrUHCrQrLIscb9LoFFvzgP1kUusk2Jf2f
ORnaevqaov2XLHTDaAIaF6MUvRhafDPJ18zbVYNmKG0qQj83LVihUyE+539FsgJ3
u4moA7LKzl/EUvUBm4lFVNg08ljQQiz7CIBM8oI4ua33rVzqWsE1MzXd1On8f5TI
dZ5rcD4GOE3vw9WVLvZM7z7Xl8bcFFoP6LQ1G/HOICw2haNVSE0vRRzjba7Npc7h
8ORudLNVU+WoIzXW7alUu+4mS497eInSV4KuDzzG0gick3CMNwMzYXHELJ3yUY9x
Sh05ZGGEakjYgahJEqeK2OmrH+o2vOibeACj2pRFcaceC9Pvjnm8BxHQ/tcM4Rrs
DEuCnTxHT0l0jUB8E3T00N05oRmH0QoLOhMnLnI7uI7b9NywnUOv6j9NREp2HKr6
oNcG2lei6X3qbnHzqPivNAdXC6eBzO8DFmv8WB1E89JMiFiVlUQNgioZ41/XbH1j
nTV1lVEkuYb/epXe2J45OIm2dPsBD0FYJAXalHSneEL4vvFNf5dfU9Wma2JGoQ9j
eHnhxnzhmsS/7vyY44LH3S8lr+bTrlDP7KKl5V3N583LtESUQXXJnDdUY0ztTows
qNKf9HtyAGqOjjOlpb8vyaYtp6m6YOs2eNDNGxu8AELRZBFM3qmuxv4F05m2gdKe
r0ITjyZXhyef1wHH9bXyLP3yEf9WuywwU2XIEP36MFw6UnKp5vWtDjwMkCtQ+FgF
VkebT+2a7w928uxZZWlsKL4AWhl1YSBLkmoObYLWQwnVkA6zStGXEhoHbjIh8enU
3bA5zISulXCFWnBzLp6vBTZePQcDDkSN3s5OqpZW4X8kVXQIq+m3LAjYhx7UPk8F
si4LgxUFlsCM+og2LvnBgrdzNrTTHZwHtcTUf4IMB1QBwd1/mpnZ9vVuKRBWGRhu
u57f+vH0MhSTIsERKoP6R3BJQW5LC+GhKqCxIFWp+8YARLWUBeu4YhgOf3LeoFRY
sqNiZTbIrnnmFMQK/bxquHusamhn482wzwQsYC2ILZZY6tcOIE9cTgYdj44xtLLd
QpgGnCmqh3r52hSJehtJa5WDuRIC5ncnXVU9CGk1mor3FDrx7J1ntDoVZvsSAwct
epCAEqrHWVHpWgXF+msDMJFUVf62K24pvmpw3XCG68wn7xPmpFT/qbsKHOoajAjT
NvTIN7ZBMBZjvDoOsamDQstHzS0pQPYaGwnFjn1cXoBiliwq8DTDbFwHj91gsgQa
BsmF3Gf7qxPIDQs1ZbxOMhwts7Ya3xelaAhTYfLCggviogFSWlI54s7mrXjr/ock
iWLvmmvrVPDruWKYSPW33CnyuH5tkXu5QoANbE0avMkgVOWKTs0yXPGVArE/x/qh
lZYvjrqWTcUBkJdPqNqZDTlEMVobKLMYG+zVz7GNZ9OEQjIFAN5rryOIQzd7lXkb
+6kKPvWTMEGrosEzMmwKDWg50OrCVG+KUkE0inFxGlowMTK+6Y6cgoQCSIIDe0tU
CpoK2mysvH4+ptffVKQOibAfOKVDDqBR5pbUob2spZCP2bMruUzxajCczVq0joPt
+Ba5lYFMoJY9xWqaVj4KBNadwLl+qf83kDf2NgpF/QaQiISPPOLOTmyef0N4KfNq
2f3zBAoRRXu2Hi5CFrRq2SfaUxDCjGaXjjYKGx7Q/vjPu8J2MtJIEonQ9sRVwaCS
GqYPP+AN68uYW58aUvhy7eKTf0+LGkjawp59p39RodfxBzIsCdc1QCsVz8SxWIcO
IArZaYpaM8fSZSjjIN7tEee6Wn/q73sFst4gU6GG1v+ZQJNrPvDuDyHAg86vqI73
0dDCWX2zMUjj5enkr7fcXTQUp8r7S0N8Tne/WEdV0aPCvkR4d8Z7ULg5WVEc+Zrz
uKNEhQAzSFOG3USABBbtiDvEwf16Y9DrXlBmc0Hq3dB4Am4DuG+yHnnJ93/O3o5E
t6Wf30PGeDZTvdnYmOjrnGAUS1XqAqEbbgwYHof5WuJ80D4nVlVB9PGT1fR7dhGu
sq0iww0djh7akffFeX3x7ON7wBlQ49pqpHmEJogHAd/6aB5uXJAk2aX4NVbxnJc7
aHg0eD+a9C39ar9iMh3hynSuFM5E0+01Bx2h8PVlSMyGdai1eKHWKNQd+FIdXUm3
LE6VNCKlDNyMwww749TuCrpv1wk0JCxbn0AuM50jVT1D+cTJFpQAIW2oGicLo9mK
lXZgePd3iCeJQtPrPPG4T3Dz3xQ51S8cDV78qoWc88rda8YWbd0N/w45bt+O3gXE
MNbW8Ell0WC0G6auewrJoAdFEiKcmORznqDNjSLq9J4vlKN8S/HIQnSGLh2J/5NE
Ozm+fU0secbLkBFF/1KtuNOM+H1J/QnIVFqY55C9sMRFXTIeMeHQLwgqtIi8N4im
0XNRwCX/9Gk5OU5LaN9uG6yS2TiF7CuSSQiqvol1VT0ejYWBwjQuXHlMduk72udf
tOC40Ym9HPuas9ZkkNqedf2ZhpDvyh6n/CKsz/g5bzc9LWJ4uZ3599+b8lEjNNC+
BYCYA0lJpGzk8YLAzqANAHa5R/VY895V/eA24Pj5cy4TlJNz+dnFVHirOu6J1dnh
pX+f6ztcoEi+pIVeGSHDPYh5w7Q4MePvatLdYYu7rcujJc0eRL820wYnQyoi3xrh
K23rjD7QjJxNG5aNglgeWMhwqAhcoTCZlZgSQmyfFay1kA2JTG2yBUW517hYnTrY
uVRDizUQ4KUM4VlEv+4MAV8p+z1fAYf9m9uvKxZTVDv9YC8QGnVpRQItq0RLeNaF
PNEj/gbPGwf4CLTEmnP7kjZY1KmJeFjdSXOXrHWvahMXNfA9GAsmOMkbYXjNsSl/
8fgjeSoKQOJS9keo2VFazhJuAnFyXqFvPhduFED2rMC9dUz9yMTaE0rfbHjcG4CK
8oIVYrmB2muSNC7PICJrJmj0btq2oFt+kY4BqRVHVeT2JGhW0xUUuzIq0YcIvdmf
FmyNSW+eRyMTPoMDuQ/GA+9bcTILBvIfXUc32zbLOpvzIPyj0wRSK854Fz8nsTBW
ApAftzytT/c/IYAGiMCgTwj5TaeOqsBlhuIyvqLajtBAR3GN7xUY8xpzPDgtAK5S
mllu2oiAvm8wLsWHN696MGTIdN/G2bZtsxb8+G1JvPIFQW1ICyoXn8i9Tmbigqx0
90jNNcaFKubmviuDagmRAkeC5EK7gNwrf3z90ulHELk4qam75Mi0p1WrO61lQiYQ
MJ3KppikARZNDN9WHMMyEilOw70E42gut7HTnw/NkHZVS/31RjZBhczuq9rPiNyt
nuamHTRTznSM5OdjQ7AFzNrVNOQ8y+PvSwyUOo9vKYQ3B3NoYa5NnKpdGmN/1XR4
RSZC44pMnF+IXcOzdQmQB0JTv9oYv9cJEqVlXjEhKG+MfHt7GWNq3bpoMEJDlQMG
aZHrEJPaGfII/u+mrJBgxxzBwVb70EOXgPVXZ1tCf+uSfIhb/4URwAh2zofIbcR+
lYqLZcjWsMwKIRYOWHPjq4n/xqBy2aRZ414rz2dAbYvh5v4FI5lmcr0ZBRptRAvR
Y7JTEckepzY8eFYaXjIOQDCxJr1F1WrD5syUcjczTkIF9kv1+RNKmHlnTasmaLvM
t24uxaTShu2fHiwsxgLTdm4NeNZGST2sDdqmkSLUquItKiHbfKqvbvGUgRoP5P7E
Y1zzKFHnbGonN0wb8s5gn8iwY1RJVG5R+kWLB5MiV9NLKm63IlmIBEOGnUUzs/aW
TGkl1gLlLdpzz0uXw/KFE1o8Er13hKvS2aVZuSUzSzoN18xqZyuaY9lsXLXbacS4
fY1Tc4Lbph2lvNEQ4hpErpqtqCA9QcWkWgQ9iwPr8wVa1EqbnJz4r3TGJjkGvjyl
ZZD8W9W/S+0BJSyeUDxF1eTO8MEjJBlmc/869HBD5ifrtRoZ1x4tj1ifKzr3ycyW
qQBSmC/Yp1xspEr5yGXN7DI3Sqm+4Yf/I76p2HEpcQYKRxzoLwX+WRm4xA/69eH5
GzUwEI44uV/WsPRJ7wg4+cSZcRiAriq7TcD7jBjeQE6NwNFf3znie+xgOk4V/Ro6
k8syXRrFhZdyXfFyijSCYGGTe/+Qx//Z+Mi45XTrPcrv/TWCUkqQ1Q1rjx7NYUBk
dXrYsmanAq/cmbrS6mW/TGmHpfSIVI1/2K2s+ycH61nzWyJi13LLDynyiN7coiHQ
ZOL8HrvhQtjGSr2rWtVVW9/iO910YgV2Zof/76tz1Urn3LombU0OSB6IwRZWvb/7
4HmEsRcj4RpNkNmdNyc+wVSMpUeKVfeC/BDJMlFvoMK6PsXhKmdIBcgh68eTJWOm
loZjLfhO7G/5n2xmhjeWbFFM53XZSVcl4jJyPzikHr9esQIF0BEbbVCrdOOahZT3
FKgkSAZ4+o6mI6tcXQi0vkL7eKIreSNHhutspxxi9TWlNVWBdJrOVE+Uy1oj+tgj
XCFA0JKmTgBfLDGB4ts+yo9hm7/nWqQb6W+MET8XHP2eW0FIHA0EaGOx4gkAtMGE
vSOHmw4L+tVDTvOw/NavSmhETY06dxd9lG44PS8Ch5nI8+E7IEOoaFtW8pZMIKdF
BA8YOAIrdFOaqcr8eRs7h/94Bf73WRnKjTzrTaVxN7zYeQI4d4ur+jnEIP19o4VM
KFufPYzAWlPcTlQCueOZ7hB8GflvH4FcmyO5W2hQJAr6dD8UWfE5ik/ku8VJD5tq
3dbLmZBssklO9WOQ/v6p8x+B96sc1TNWuYM8yNeqU2Aylz7dmLDKb/rmF1etjskp
jONn0sPISScnbFkJWum3EToNFCRaq5ZzTNwwSmdHgLOdrG662B7AQ9XKtl5fqK5l
Fj3+eupw2jvvA56IJ4GIwOxxlxCujrAeVJ8MXqVA2Ym9OnNRIZdcqIYfukFa6P+3
uFIw8BoP+AEFQ94i3/DpOcW2wCPffwckwlQHOY/HKQEyKFXfVdAM4Hl3WeECBBR7
PI/AYJP9l8Uz4YMmPjj7jAv3keZnT+J8ZpkMpjj/pK7LoCmsHDzXA8TUNchSUcsY
eaGgep8xCUjsxzxPqEj9GzCkYeseUDyv0lsBvjqbRj1VtqZfc6ovk0fudHZWFuM9
ZmYOgZVHWujRrurA8kADaGOtnF9Gb5nIaPJmTJAbDag8c33AgkSvrN8hCQiEVFWH
U+SwQroRudl3t2i89hrnKXAFKCYoDT3m8xryFjhOS7XHkL4/BOwqghtm1iCAZhU4
VyKKQo6OBj26+Ld+711nnFPM8jnXKq8nhe793/ie3YJkHMbVrGOULM5U0V45edGe
bLuCOyPMcd1Ft06ZQNFTAm2XNU/hosp2+Zj7LXJ5LqlJcArRIKphOqNkwDRm+4QX
oiSa2wLTlDG3ewfrId6oRcMizOmz0gKQSMeF/+xf7wvAhgbjaB/aILE6Gh7cjITZ
c3UsnChOhddwh61Fyqgpcabm8dy1IACwLB0PRBELUGewl9ij2nwFhXK7smC3Xc9L
+KNjGVFbLJRmWjBzb0AjrQ3oJ5kZzBdIKeEdMSUSOJI9kKqxdqL0av3s4uC4nKmj
IGy51tjVFTvArDqe8fERIW29x721sSP6skYPBsFcPI8h/R6rZU1bbJPRlADpfii5
/QMOXzPQ9KaQFLJht3bQ4dksNGWdtlZlecYIJouUC3atRqY2PylqQK33RQ8No4vw
VyAYijA3SSI1NvrPEmtM2Juwu6LZ3a8cY0ho2S4BMmSz8wtqrdo1vA0z+wdZGnNg
+A0n0TSouEB3jOJ0mZb7CgFhHuaqOa3ts8jRrEkaS9174mSpv1IErXgupz+0CpZR
k+lJveIYRC8o2aCdo5FEEWYdFmvJ+Zrwo0kvQdXKb/tmIi5Id6kMZJsiYP56MxVS
IjJTq7gpGffTBZzwdVu8AlWVVNNZKT4jWbD6M7FgRebDiPLyVCJMAL7bz/DeLlfJ
jjSKG5WqyklLXmnPO7w3CxRJERTBTzA01mwX3AGkLcEtHAIdyR8HJF4Lwuf+RJ4a
zLI0cKYHSQrxmTZNHJK2a7Au7GFwdpoRd98ERr7jkcIVhKINaUltTIoe0nx2tISK
NSth+FKNWFInSm5OcvMy3rF+vR9Y+VQsnZYDxiJ6ycdikW66yFnv0BkaK0S3nnuO
dp5XbWDzSxsUraE3dZVo9FYuocSLaTx0KtkpWJNMBYX9vYRXJ6Iheu/Mp/ItIrVS
gOhx9WJMC9dMvEgbj7AAi7skB1nUASisceArnSeOmPmKeiFDNmlF4kW+ovn/Ope1
2k93HF6u/dDX/2538gIgXr+DrWwNLk6oq+NJWSIkSuvDpv/Ouwmo4k1mBnxEYK9B
Tc5trjIWuIfmnPa3/UJeg8HXXusgcAaoK6G0EwUfMRQxhwRpqw9QvKFE97jIv82/
jJvvqg0SSBy+OvhBxUu7Vsqwo1W25MeGBMCiYguubJcevXqRNau7Xzo4nXlufqKz
udduwGSEK0Y0KSvXPspE3rQVXJDxFebarr9aLsobUAm5WEbCc9C2z5UUVrPHsnug
Vp/rDTbqLbXGsRDQpRUuKChoGWJ7N/ynqucPa8D4ZPnBAztJMWuyafdarSNvYHD2
wl3yLvghh6Y6lsY2/EP3qYxw8a5Zd/9N6pTrJxlcNL+2v5cZGor3KEHoZO2RJ6ta
H60tPjmHBGNMnq0eHJX3F7UY1hMZfwLS3TU0ApPyBHI0xkrWrU2MopgNRppHaK7D
nFOD24+aNx4q1o7wjZ72T5q1N5N+GX3uLVX8O+dThEr+b5IrAiJFv4qJEKQm/h4j
Ji8Wy5uFiYckIq1Bio0PDIQzQzNuz0pDV6iI4d0RLG0Dp1FyGLuMBlEjV2W01J7i
ULW7CtMX3WeF8mD2WxOrM4/ho8zRKNpNQufPxPk0IJkWDdxJNx0uedfWbtktCUpP
nMLYG8Abrd6C8WYMIX/pJ4iliZntK8aNiOr3yZ2WvoWbG7f8Okb46k+gdfA6GKEi
yOSLNJZHh4Q24O8y7RApZq3jjCXiXG1ueE9bztnsQkkBigxXMahFrRPkaH/q3rHr
8gu5qDbsFAQouiC5R8Ajf/qNbNZYjRElpMsYA/D1p8BWaGQxJZXL81RWDgicknah
kuWVWaUXqgi/dDIGPzdUoLlrAGcX/5jr72VvZ7KAbzT6wACnin2+thDcujWmgNDH
g6+hnzkHf6Zypa97B28GO0YL0RE+O11b5TaX+IRKApmO4IR+4nOLsR79nInX1o4G
blhk+ItDypf0qFbkgt3LYOk287piPC9Lkpv+CIUsumSJsz013a/olZkwB794RX7c
SpSK8GQBvAumrIAb/kK6ETfcz8LNbKxJjZdcbLaxQ8VxHozhP3Ba32lwjrzOIOSy
DOsWkwu+LW7Hs4f/NrcMgkqC52+9GVs1+knxknhxX4gLljy2bNIeaCxam0WSVPPu
fl6YY1rwmjLnPhv3yZ38RDsSNEy/2mbHZ02gdgLDqvz3s8Q31PObivn11b2Er8lh
cnIA+wzxTSjLEQY8/SDqW0h09JzNTifN+aYH0Z7os2BJBLE3JqBBaH2DTUQgYrB1
5D8o0b9ViPn5EJYzRmwS3fqk3rFj7x2sh3hJ36kLnD72ZzTViiPFpcDC7LAIZzap
cg2P73kvMlhlx1y8rezKUVKX5IT4B6Sux7ICScgZFeJaD1XuoY84VLGetGICytEe
RM4WZU+LcJ+bjVsQums5OnY6Ta/JUuMUOO4DAM7Ol3Fq4QByZbwr9rDCafz/DAmm
JbYnCv0x70SJyyrcGP8Wy54bhjWpQBjp3VZ01vjuWaDdLqMCjDtedzJ+K6Xr5fGZ
KR6urNQrGydI9vXrYcMPLoJLgiB4jCbSgc6eoiZTYG97trrhPW3ZXuFUM4OBtxwB
oP0tNHltDOWtA6iKwUyVRAm279B0aNUPqU5S5aUxtm7xBtzazpuab8m/vQSfz9XA
E9R8RfIEGdJnamas9ItpdsM3UPYLB0Fei53P2RAHiL+TJ47xFMzTpLpxZh9LuxRw
wa6AS77H1n8nRm9XEjTuN+YnPdJhkhmlogceDkzz9ycctq6R5igUzmO1zynJVQ33
seaQltM5Wc4MqNft4OpzeWgveQb1DPgRr2pjjiMiVe7vGw93Kj4nxPxRKT/bCjD9
vezAPLmmcgAwNCkn3GeUws2uHOG+JQ+78nEYHB6pbyhZpEWDw6I/6EjEshV4Z0xy
hbi42d2v1f96Lz812sDV+tVFNX70VJ+UIfDp0A3IJGK/GeUupRiNfpCDB39Om0lR
8Pyvcy8MRlZzAKGPGC/OHvxTV0c6CRvKkhyIKlkXFovQr6kdaYib/IHU9Z6Qlpey
ANnuQlP1nfifqmqVnwC3MhgeCIMw/MDbSgYa71mTG5q/eK2yxbj5bA5HYNh8uXDz
IB0iJErDACyfTeBC1hmSDFXm0N0NOW/WLu3UenLhRiJVfC0ZpceQSgF99KjklMdP
Z+dHLa3OhFmPYst/xeYM5KnCpMdBxpXJRC35xN2JWKGozKazCy/kjRv3GtolU/Lu
4fuF66xZvyufDBDCMbgOupm5gftsyPDqKU4QQA4zGVmyxATyMV4WfLtr4wMX66TO
KhvUa4D14wZZrFAZ0CC8ncaYJhAyE8n17uEPhMx5kXqJDmzRRtwCgiwhiXEeUUdc
PhXwWFkxDS9RwGByA5EzD9kj9Z3cOZhhSKm/Ud5OSjq/vnRR4mnLQf5zQx779VB0
e3FJ62KEXI1ny8rhCEGGgnmJ0PEE4rz8sBmtiwC5M396esH/YKrm6xlII+I2VXkU
t8EF2xm8vTJPJdPlbBD2juhUE/w7j47OwzoL2QaPuufe11fZz+puS482fgvM92gK
w1WzBC4hCO4qHZBUViuoOgUVLotfprJSsbBChCaQhElp/Lf8SBu6JmYn1qAUeYO0
XOer+9ipUKAKLY3ZJDJPA/gGNBFwY3jqpYn78FP6pWE4FMMY7QWnyCrxOMR3miyn
U8Lxp6bRmVMyNi92OwuJ5I90YmF1KEuR5uHvdYxufzYvl8lYdnovxgy2Jdgx3hC8
6PknxH1Xd7SyHg9t3qFbxl0yODnDOm/RPWfAxqRmtwXvR6xZfcEWvQtvmY7Ni80N
nxBOmmKGYgg5TxBSGprSUaQ5V1yzSZ+sWWB3C/ZYteTX7sJJep3zJJQJmrabjPNq
ttLPJqdbAFrvsLWD/NRTpr1/KKhD5ytzoxkp2RNRKjx5vIXSl1j8vq8hW2LpeKSu
EXLq0Wy82Ay3/Y07fM0YynwwYvu7UYTGZmK+ZKJHalU95mSWpfrKbPf3rOaspCLO
ZDvMODyeyv2oQOO9pNjqfWRCIYAimyR+tumpx5uDRw9+oiAY7fYA/y12eIvy1Lye
aQXcwXj73N4QSx92+zdoBRnl30LjNpdTAHku5L6Ruq1Se5ZXUOVBuwmNqshXKbe0
uVW6AfZrdTS4PBi62q0MLFB/Z9GYlXWJwznql71mpKHHZPOXAydnHnc0yrt21l1r
TaWYCIt/ntw0vhhY17PaR/gngmNvylyvZIhaK8+vqZ0VuHGuNAc2JsrIYVy7ycdP
DKl61kg3lDnK6lW8MVndP6ros/Lm2m/4cX4VADk1rrwNDFzQP3JILPPTb0jUvKIQ
l0impxXkHVhbsZ13VBr2SEOMo93eTwV+Oox5klJD9brZR/QfA8/EAphYheKED0KL
V955EHtsXXSfPhCBiL7iLz8uDO94JUywdxE4G8Ce9/l32uoI13k+SB51uvmk/dpK
u/ZUimvSVh6TcEawZbsEN/LmX30MIYWgojXL+zfQvqK7+A8amtIOb1aXf48H5P5K
zltvnPs4JDRpVx5DKqWN1XzOfX5vBzLTsGR/snOxWASgiZIZedR2+DQt63gQv1ZM
HN6HJmTXoSny3B2Qjl4F1YHgjGsfHSUOSN8fOC1qzxZHPKRRuAFtYLFoeCdeXt/D
Y9FluU5p7FnXmKBbHR2qeyE3YRPhDZctoK1OQ6ZlHggRYlKtUicxtHAX2zB0Zkc+
RqNJ70O6T92yw0tf9BMF/10EiJL9fQNKwjekP3atghIk5CAxcPNcVxKOm+JvBpIr
YLyAnbmbBI4BAwOPWngsUHjHUQIiHaCERM2XOK6Tbi2drmHbS8fM6g6risOh5pXo
MkwPEr3YqvglqHt0cPKxYfKa2YZEJPIseJFmZzFhCpkyviftDUzZkK11NK+MFgJz
b8OkynBlzmtBWD2zcYjAZGaX+MPegVh99oOhCo7e4pbDURavdASAwySrp6AoNQZn
6ILjEF4UEymS0r6sTq+ntW/CXBWqCGs5rk9vQIUf6aZGpdX82HP+PJ0s2wAeRt7a
3Vab0/5/Vq2oATN6FuOcr59EUEWytFfCE1Sj94h9yFrjgJZW9qkIlGErOgeIwBKU
BLkroeQcRP3ROHqGE1aK+tqKpyc7mWjJ7rle1Fdv2AZOIyK8qWVsqCXyi/C3T4gM
2zsWful8xKfEBwKrY8aZ+7lVhzW7DQTKhTE+b5gJthf+vaUvjYFUeyZbLJMNpsJ0
021gV0OA+as0IEuBIR3kMn9Kg/fqswAsw/rv1rJ90FuXI2uXQdmUdbbxYyIj1/jE
Rud8AgQxA6RvUBktIYiHWlOQx0CjWKxnCALIAHMXs4wSS/AL1O/6yZZFBhYRM9ra
9KDIVn7QpLn5uVsD5wAnHo0mGlfkbKOpr7KV2Ch24p9rMx96CR3EVczVjiajbhIm
iC1GbkbKFPV0/1jwhMlT3Z/PXm2hYy3BZT3r+iTTdhLlX3K93LcyyYTE+KnTTWQ+
QgpJi2WbysycU/kqNsja9q5wFj3EbjtRP/aj+YERtzXiu2XUz79jd7nCupUps1ij
gjUt9Ewt2uBmZlVl2mo9+l69E8yrRsR9CuHsRbzWn0+AyPUR6Ww0SXMHqRgobROo
8RATfOVkSrWpBD5ev8P0/DWnIJjadIBG9Y1fvxoeGXOeTPMbRXuCZSyd60zn0iwc
fEKDr2FNjx6429k9o7CzrpU4BgM1Ng9FAoBLI5w9QuWjHyYp8HLLz5o1K9NMK1jl
C+AFcJmtuPZvCbF29L5qNQ7TstZ9vZSUS+4gAo/iLl8beGrF0oZUcnkdzGJ6ilt/
1c46LG4YPVmHVxgDQSqYFSxXWNm6m4Zm50UTJzJBx8iT73nDmm9ICLQO3Ph6aM6F
ofb8sB+/cMAWiQyf+QkToj9ZC+EzoSBNTCR3NbWge4kpp3Xgys8eFeJiNg0SJy7n
hGgVfzTGQAe9LVugoXb5rV+F1Di38I52bMdPGzIBDBwUeTYjd4PiuHpn+VMwhT2c
VCyiXmg94sTrtmtzPwQbro1+KS2bVxFINeLTMzP9GcQdmAfBA9xk16Or5tceBlBm
fKMwqPzCdEDvSppkzH5Qqfb8fFdkTUHfsbafZBTVmV5uRKf4LOTuIaqwAWts/2yN
V4BSsf+2SxetzocpbTIcoewryvW4NiYi7dbDGJ6u+/4+3ye705HDxhui24uaeK5J
IKqRPJsUVwRxg6JGUDcBp1s6ExAAE438dmyt6xqEIbiAXWlaKKQ/OWC+M+ygpSg9
x585hAHxSHNu+tYWVkzyrh7pT7WJ3SoTOl4sNQJsHYJXS08l+EowHNcw0C9CnJKw
v3VEaiyew4mzr8Fn3BysziADnY+dfIkeq3gCaucNp9JWcW24IbPYtBEIUeAL1a/u
yTh0zyeuAEPYmoUXKJxGCaybb4V/MsGr0o7MVY04fadjdZddHOdJQhivbanXcmlt
bgBjel0v7gTCTahut1/U9RpYwxkfMb+Jihv0s3pvuS4WYNXSX7g2Puxz8TxE7f5w
tq86/x6Ddf0XiinpRG0X9aMBnYY3yyTlvfEdoPqpwW5DI1KyDvFve/c3siNjjYzP
HfRKHCptL+3MmptDqjsV452rVBnsoAzXL32hRxathY6U+oxappMuh9v02gEK23Ez
TSyQ4cXPkdZjfJN6lXE5h00O7n92JFmkbzwOCTsenUz+vjHZk4v8hTsd0hKYCl+0
Naw4/Kv4HMaZV+/ZWHNRRlrnmyCeC3hhs/gWqQdtVE6shfsIHb+8717VO4kz3ltq
0KWs+z3B/tOuViZUg8k3sZfLFZ6EzR7A7IH2i5K2/Hv91GiQhSVh5tzambeH74A1
GVUPxujiz1DcMe+l8cOihB3RR7J/Aa7VfBsqfjTBbX2cfURntkfRE4lnlS1vViDk
4xz6kHGgIUCE1DNS/MjQYG+Kr22TEX2GxU04lGq+AhV2SLW8ALojfgkYRTPgbgIn
t01km4t+W22+dHpVs8ximU72+Kr0R7t0u9CWgrxv8IhqOqmImy804eGdDSP96Fyn
YJeF/mPYvIWns6qfglc+4qNKHrWACX+SzXJAamnaD9zM1o9k/NK9A2kWKnD6XS3v
+4qN51sEj8QXGguXvEW88uTkt/hW9mJnF+ew0LiDPzzWPWnwgLGbgW1ln+AFWg92
hk0tF7Xtsz4pV2ItkL1o7RPE392NTrbQGnHujoVsaPaCCnYyw8JX2pIsecZrZLXu
69+EG+24REvfQKJlfVk1Tp+9Q9oLrCmE0BmHGhUrSGvK7EWoCfchXq5+xaqEUJJ7
AQUKgEzpZ+x7XL6fUWRFy5Xv7b9b5Oq4SlbPi8mCoWE/hMivUUOVnZdx1Z/rNht2
iktN18anuSu+QH1OE/2lj678Ye4V7y8fkIIrH/w5FdqUy5wU0diNl5ASsD+wtoTd
rrbUZWu7KRbal6yJq8Nv2QpCAxFjSMnbmTiyBjxlhuL4hoaQqWNsFzumYvopVuvL
uNNY+pbc2VH9rTsRyBwvy+5lP6RlbXIY8TPs8TeWVlpL+XETmnz5v3xy1OPFRhwl
HnuL2zAkHdOoQMl0kLX4tAX2emtGCTN8RJaK4WdzYS5M4ZyFGjlwwTXa4c5aEVAA
bBAzKXyV6miWlrhsAopEcLfUfU85U6nmrlSYSoVcTMB8uEey6FZOZOYFHecGG5RU
0O/JQCu3xyhXCbqLFq0/XV5qQBZ79GDbpApAokr7A6+asLfesF/phId5gcQCwBw3
aSqFiRJaDvl1tigUVSky1uSxcBcxpRGiRLX17GHXWfmPCKSHp+/iX8MDO4izFWXF
NOQzuio5986cNm2zk2mLgwjEBhP35260bY2rDgHzgT0y8RwPiXMxi72Ns1fT1fxj
DWoL1HtfFoF4B57ZhLKiD6VjmXL7pHoiRDpmt+PaVdfPj6ozTuFIygFsY81az3C0
nURlvUODhCdnFbjlOJfJxZTYTShIs2mpijyc224Qk8Qy1GP5W4jcksqraP2Inn1I
J5dc1gv040eiBzcLBe6EFHOMliH2gtu2oEg258E46SB/sHnbsaiJVAZGyFHwfBjg
EqTo8CX5vnCJbAobQIAD6evv3UrsF7unYcxsVbC+C99E+9rejLMJiT15a6BKNRPP
YwTY10WyRktAZwQLlQbRLQFi89jENS/UgILpzTHivSwAqA4tgLsQC4W+eiUC0nXI
t8fEp8UsKGmggpRTkomzfPOfiRGpc0cpotbBfF7m+qM6wbzvbiUzovK24FFdnYkm
B/vGgegW77h8ByZksU3SGtt81lDMoyX+puanY9wwGxmJaG3kzgmfo/9yAhtBDF5s
Xvv6HC2q9tLNXs2Y1KARNJhC834pWRP1PoDhdXAlMyARtjM56EjFg8RfYlvTfglq
Z2rAGLnxrY8bIoIDD2/QdF3xuUpOkPMsLqwSAToyXJ8JDNw5aEyZ7WQHPwPhAYFZ
VVP11JSIv1Y+DssNimnHPxT91MErJEa9fHJWd0y6B5inqMv7Gk8NhIDV/pM5fkqV
evXRnCVdSpW56LpSUHO/RRCMTa+2hfQpEix4TPwYxrqPwR5ad0eQsiYhOeQz6w8l
q18zysSfXWIHHgK2vKpiOPdRx1kiAvgaEMAu/WjCAVmMvTaPZr8u1a0HekqoI3Fn
zxREcuiGQSpm6ZuhQKaC/TBYW2Xk9X/vyAn3yO700UL4ZslIbcgbt6fnDjkYOaOC
L6KmBu58Lec/nd8QDIezOETGNTGfQvAtsdKvZF9+Rl1+ldFNz95QfrfHalRhYhA8
fV7SSlqhtKLr03mTyp+7JjwhHrCNbbwhPhY/TauJiuc2MBKeQD9w/xUSo4TQ8it2
oroBN9RACpux10tBXESc8BCFS2srgYdoKhGphdbUag66AckF9CGkRdA++xc1KqH4
iNpLahEYoVwD1kMOvkixNNVEhl5krwuvba8fbhgwqwVCSkJ2/uih8w6jqulMpBQD
djk1eZjFmgNW7XvuFZGRjyleSLepbrESBhRF1bRajkDrGoJFaRjLA+k7ZdRSN1YR
t0LVoUKBK5wtOxk7dOugybdMYW2oLIIo4n2vnHl6ufnd9oGew3GI6od2X9/boujU
vXH3sJqArEBR7muwGmuWDQiBjiDEYusA2AQr8Vch8y53A+nd9eg4WgcyA61IU/c/
bkWaBapbsu2dDfTrLWI7riiAjZwMD9QdF5aVQOZI3Nt9JLcTHb0DiGIpkVh5oCfw
b+jBe+DjQ11tyDRAYxFzrNIZYvb1wPF/GBRtiyOj4P7AYt4zcfyHPNVgeoJO7od0
wbr6XZGPfE1rsUec/TzNktQczD8vMmLjoa9b2izVoxfXIxcXsOeXvjHG80FhebKl
/WvRSVpzF6qtKXRWE/KSx0WJVAB8UMMj9hc3rP3NXqnrXJuCaSNLC1pZT7N/NSs3
2HXYXZ+k3WrT788WGl1/tIgeO4Yjwog9P0EtG5nzmC0feePcO2cn2inrtKbjnoIE
MPsz42wUffx0ZphocX1+LJJtiSo8XjQfjQns0YGiwOOMU4bYkmOxUdO9mnVTgvqv
Q4Jwb6KOYuNFY1i7l0Kv8OMH8D/ALuSjJAnUPxBq3ZEQuNoOYDQ10Hwu2rVvS2lF
7gimPoYj1TLaKyINCmOf9kqWT3QRRG3jAhmITiboyRGJJKLW8JMC0w2Z2YLlzld6
ITFP/8QifHIM1QdRP5hgCSS8/z4ZcRPxanwLS8CQjE+sa2Pu7hLfKvhLJhWlTFrO
AOg9Le7pGYGAMqtXGoIX98dNal6/Ic+whuFwVaHlgGPrLHKAPlOHJA3rBYjvwrA3
jQAtuHkQ5wLQIRFls/GJ8bQH/kFrgpUhTeEfDOwOabyEjxHUrll51awBIAct9fWw
bwFiGHqiQD8Kf141vjWFZhAoTfc+JMwWtT/Kzl1TR8OgwGCCEW9tUeAt46zh+G0d
3u6fUqJfgxWdmdgseh9r9pJWSUcIn9SShheNqLiUHvhMOtX7KmrvjLfEdKcabt6c
ZhAGjEq0e3ekTVOPxry12MtwRNtIF7lmhi3Q5DuKwP6kwrOPhrqKnh5K6j9tXIq0
R4HdjGbODHtY18glf1eKfg+JgPD8TCaMPgR4Je9siep7TzMqaDTl0gzOfE+/nLnj
3ScvRlKOKuIUvs4NbGwOZ322g++6JipAl3+CWg67zqCaZ8icxa0N5wUB3nbaqpRl
DAFyO6sP9BG13JUPly7gGH5P1IqIlfE9Q81vC+l5kIRlvQM29e7WEMlWL1RCINpR
yBx2WfSGIpa4qv5qvhE5mSwVshBLe3SHGcXNaydLkitkVeClg3gn35YQDJNIqJne
FJZ8hj3kdekJAjfysTAlkGPFhi1zxufGMVb8bLgG5e9LLLXkw+QwYzXC8g/fyoro
8F4SkDTgMkHHykYLBaDPO8hkVJktFqYj2YlkuWNJcF/fB/8FhoHseImDBAP1vhOa
TY0Zu/8kfGqYq47EU+Sy8ntzg0GZ1VikXjnbYWvkcWiZFiINhAkWWyGBuAX9BsLX
A5eKsaqACygmAaE6xK4L3MVi+aVP2KmzPiq7RnFPK2uC3hoJtuaq44C9Cvls0xgL
+tHzvSLqFVB01uP+TUbM9dGsYWvlNAPxvByZOb0bXet3m+CuXSsLn0zBLXxU8j2L
V3WNbQTdkcwR0x6h++pSovG+i0PamMdDBjjC/35O9B+Ruhxlb0XN+JLGjwORYa+8
wRnRhf5PRGBKafek1eCxrMPAaUP0ct9bkgKocuC5CUhQTod6JCfqcwCUNQJEhE5s
5RlLU+qYz/opMVdkBjag/J9VJLQcGe6fuQZTyeT1clTXBOFOXGXnUEPvrLtmryYy
qaDOdz7CozhjF7LVnmaWRmI/IlSFXg7EfTjoFlbbKu4jSaRLH3Gp9JgpUgVOsc0V
yCDDfpG5hPa+VwfDG2pV7l6aRW5Cwo8XqL4splQe6WvDmuMJ9uIfmcBk5pveV/wG
U3/J2pilF1Vc+7ghQda8aKlMiKfu6vP/xozuPXKVcLHGRNcSPzqsbXjTTirXJ/aN
pvR5bYIsG65vejIbAR4vREFbfYw0YU+Aw5RmV17uEW6HxCZgm8+wesu/iAR9T9YI
EEZEQy9i66GW23+zPrdSuAT5lc7pw3uGJClkVE86eU1NGwT7H3eyP0t0eKTsiJXh
7/B6gpSpe8pEZC83dcZlwbKceb09W2rlaWidBwoHnrgH4UewDOATfErn+HNrsv8G
KHs5yvgE/5OsCvDQrUkw/F+LNeKevAowivZaYvodROWDJXdsKQCHhGFpkUspjt9i
26EhafVbk05wIlofJfEg43JgpXm1o9hgJlaSPQRtH9T7Cm0uWym70c7mqQLEFnL2
DuqhlY3VmqQlkzHK8t1Q8OesFMQ1TEjKfLAVkkkZ3D1l0Cw5pmgbxqMfZPpv6TNi
zmgZukxd04rA6Hk33/Vwnu0/wSa1S3rrv3mRQ8FiWbZGyX2dpA0Iz0Bo1dLP3Gn0
Y7cEr3RxFtjeaUciNdBWeNFvyTSpZh8ATe1ez3bm0gwpxZPC1K2X9TBWYxrkQ7lo
9THbmwprB28qW6bpuSD/iRY30V2Ajw/aac3XgI2lk8evR0nsqElQUMRLjpdnYqgA
ZQsfLb35fH4cYIPavKdPosThskkMVxqi7fvXVKkAxKSm+4Zzr5pzpHbApxQHx//6
qwxFLIgW8lG6GhmKcNjZworJHwO3JXtkcR0Gg1Jn5B+0qeNjheYRamoAakEc1WsR
1QHOc8bvOPd5X+xENUWPn01hLJ9+o7fnRnWm2QlgTYBWhgX7W+8GH3VVDIW5IbCL
xAvufFlpivePKCofMtanklxmbaYSA1hbV9P3B5bQn09Pgm0mxnOWx/+IVXG1QZTe
7fN/a/cYhaL/RbSVvjGQ5QFIFcyvvLc5MdlTvSi3bkC17b9N+IR1fuM3IhIHLlxc
Crvb+9f3sWjvxsYoFcALx6oDtuMQcZ+PhSTyfAOmeEhBlo4T0H8ZPIyU+jadrTvb
ASwvUtX8Y/cWOZfSqqLG8b55bzOQhEX3xwU4JYEJbT/1wv6XV7ScIzs3RWLRc5O1
OJ4fIakilMXPwGrAF9Z+rPn65DGWcNuMOrcQA21N3XsuXEXhIo9k6KAtBZFFwF97
vC70STRcjwb5exW0wfMbYmGVi+Ts68zRVC8tu/Dn3KGdvTT2cCosIK4iqKFWCryX
9PIzrwl/rRgQengjQSFIUDTQXLftsJe4y0ib5Mxe4CF5EjYInZAW4L9xO/eCO2Zb
gn314RaiG+iGdueod6DJdisFoqVSnjH/DxIK2leV7/OCJl2im9fWI9QB09W0/WmY
ydhiVUVg1LGizOZ8TgPvnggi57xXLYihRhsVusBG0h6KG0AR2/ZxhAf2bNNa25mg
8459knFHTeg0cB+FMw//mYURMKTWQCXVlMtipKaTRUEhEWPqiAsBC1yUccFGTsER
6jdb49nmWXiWb7c4n7McsTIx+C+sKuBDzdGd1C6uWM9Gk1wjIg+1MYOMymxQ0nhg
zqViR/ouP16oKoFCNF3fchXDqoS5jTiGV/AOzcHpxbD0ZiRdHmAJ1tzuFCPGvWqc
B5hi9sxMjuFc7fYL40He0ctZoW1OBwGXr3TdDQiP7H+Ta2Glicx4fzXKQ05F1efu
R+QWwFotygfFER71h2pta9SNBKfpdC+SVF2B0lgiHTu9623MBdH5YE/ivOERBsYY
1tCpG4Gmu12ycb8esC69U7jm/zOqTydYLozSOAWtddtjk9ijeiR6OeyLzZphUiJQ
vmoY1OgH605mkbwO38DEo7iCYHByOwJWXobysq0xT/6gftz61Y0NW7KLLgpCngJi
V7oFwKj8tGMj5V+hzRS6Fx24M1dLGWpVwLA7+8Z7Prm7rlSE8PzKcAwJIhhRhrQI
Wer/7MYKRhBLny8732VYninDDVguyIbRPEUYJU/lf6gFwTcgTkZnZohfZ9qOEUP3
kuVna0wheNYfitP+8s5cITCBFp7zL/r6g0R2csCCb6nRu5xbcQgIH3mpPPm4DZ/Y
Ld1elE6TcyhjsA7W/0/jhzOQUJKMBYPhC+AXHXavswV+4YUff7qE+/WBJPJj/bNz
slOQZQAIg1u/zjJddUomZphzJsGmba/blRovVBCAObQaDgbCVdF8BeX0OoS2GJdl
mZ/oXfoOHhiJ3okd0MDYboyzAM5oecSqElkqTOsShvbTgTiedQlP33QQdAwnqR3I
AHWw08nITXEVIOkg1vU/AuYQSApUPfBDyS/tVsaBqbwvzod6ASwV4YQ2jwyxkM+m
rQb/qS9P56gMhf9R44ULoviXL85+FuKPPqAhDZMf/7dbl8uQnKxDcKtVf2IWclgB
qvJJ2iwJcXGc5s8PHZRQC9IFmDAHJNsFSaMXhKfXgLsc0s5OgQ6dJG/iWRVjpO6K
OfGbvYVdtmmPAsApPOPDhE6rwbaSYzxZUJfyn/C7IO3uOZ0DTG5jS31GyVSQEnMF
NEtmGZFPLmHdpY5ZOJPYDx3v1rWEzm8PFaSh893KW73Rfyv56/1qXZuuyues9a3W
mGiFOkkEiU/xvPU11WqAayF0EdU2GMwPYpTh+u3f4Bhw37sru+ab19jCIhpVPvuJ
k5YpqMEJVGlcn9xT7DggDwfn2wX8TenHMgdUDp0kGBqeOZpEqyZi9QSfEss2kc0d
5hq636oilvgDIx+FPRQ96a/9rFashS6TYGCrCZhQ+aeJszPOivqFOtrfjpFsM82Y
4d9GqDpUgrlvBE1Dmfn6E9ymMMvEnj544aNOZLjt3+o6QQj0C+Sgoo6QfK87YeGa
saMwE68LGyObB0lX8pS4oMhm6Iv7OsKaEk0B0N6Ozte6MLIJGEIJdY4fg7nRDs0o
twAnoKdCHY6LO2rnRX+gfeoIKSBaXG7783ZFwLOflaNHgAyy4Bgw/dJ4wrFLYS4L
xAFj7zoUt2OHWUqpvOfVoQid50m7qHK+O90ME3vllAAL+zsB7OvxAV4m3DxFD5G5
WvRagUsqLDqnHAN3QL6oigBnA4pIIk/L8nfhCqDK2GyIsu7GOtV08Ufr2HFuuOuj
JhReSnTSKX4jKZeaYnHaw1+uMrqgjvovdFx5viiVDC07APEGdg16Na3g6piZy3hk
FDqv/EwqQGyvCpniSoXFk+2Z3GQEhYcBWP2ApedAvZSKMUwVzqCfTvZYSrpC1hxz
Nc66jvJQ1hTU7xooRQC515E9FBAAXfJkp52tj37YVxUjpIPr1IWhzYLgwuUxGK4L
mnQVLcsecYWyL5GcrPuSzt/6n2BK0J0f3tHhxhbz/lakvRvGXmjoJLa7da5HTYBR
g8don+lkqbVxDG+tPUt5YzqGdl70/8x5wYioeVdoPPP/NwbbsrXv/oVtXMaok7EB
HL9CPqllt9CwepdG2RjiLmgdJPki24zBDswTzavu80nK+M3DKvIw/PgUo6HvVitx
WGAe59QLjQ48OhE0UCyREz1RjulxgaDzXgX7fdz4ZceqsNu7gNxjeBSh4jVgQZTZ
giyDuvG/iXJEZ+m5FQCaVmhtrl3Adphfauq1P3wb0n4Xwj42Y3Y4k2rvm5hXWthQ
TgB90rNbiSM7VcETNRwLOn3aSSKGt3Un2B2A5vNGZ/p82bPGZ1qeToSg/Gvn2Ggn
rWbIBYBjCzL40v81bCSb5kQihSpZ2dQ70YfYXrnzwnlJk0Wlk3xAFUwz8K38Lkyt
CXAUh/xw36Kpw5bHwF1n9l7dXHuwAEk/ZsfQjLa8Mx4dpJfoogtT10ERnoHg1GhN
XSdG7OnPMjj6ylK7tBD0qxIlWg4CD+MBTBfREVJlBJJLXiIGvNsYwEk5vZEgk7dp
YY96/g0EufBgC71J3uM93PbrcSarLIMnsDN6MU9tkXJWJshXXCFPgbd9NTPQDHaQ
N9VAnEVIwwSTVK3aUoM7hFyU1kW5Q98/+kyHVRWVVA2Q4pnJ7xYkUY4Uy2poyKc4
bpUaIMugoB8EU5QXS6/Jv0O8FOf4l4vFDLUpBteyL8JbTlYozyQxvjhHjw8i9kHb
a3lg9hmp8uVrv6BiK4RXSvcoCfbwDPqvL9xBTpsTfW8fc6X/pTwooAnp/t+4WHzV
+nK+GUdQo1gNNMtpkaHFMo9KJHE7b42J/2LzsQkThwKhlIA09w5j/YR1P5RoQ/gZ
bW7xloykGsnvWMYMcuFrBS9akFkvSwaDcOAP6n955QQsHCrlfD4FVOwA8pcdIjAS
IN+HYE2QUruH1BiP4PMJq1s0OcdZBzG7ERGK6QrtYWD5u+X9zJCl4di90JkaeFvh
5ujv4zKub7Gk12HJ3esyQe4L8BrG3+s3hYScaF/rSt+5O27cL7RL22x1PIKW11zJ
BFJ3HXf40tTPDP6JrybBS9tlj5GJ7TneDJlxa5JBnh2ZiaQi9iUnOFXOdRARUSkG
45VWaHNDmaSd0pxhMB5MZGedxMV5NMumMBlqlVdYwCrOzKXqQifahCtCiZU2i4UD
Rx7Ry2Ld2jL2fldLQGYqcbpMeFYo0JrKi9IVlcVG3gNiJFvWRrHQ3lMr3QoMuwXW
52NufRPT6RC5pEzCi7cMIqkUqvAb7RFhXXs2B90XUcq8ST+Btk46bBH2fT9rvUIb
tFL13G9NCeAtGNPxolzcEuoeiK76vBfiNAewklNGezHqvXl4j0UXoWSnXJvPBaPC
VDQpRMMcE8czS9ZOn1Y2bkskaymgJpJqU/VZ6WmoGyJUFes2db7lJTbRFd/k0VHe
4BHA85potGuMATatWaN1hbKJScUrmVt3HaOdujPB+iZju4bIV9r4RXOKWaK6AkMd
yxCxsuN3DBN4V8f0eMGYZajMrmh8yi+G8ucKY2na5sorvcHPKn4VsczdSVT1nee0
mN925p6jZ6aENxW89+2OHovFQgLEF43Js4aJaVptf3H4XvzE7U5cMRHW6Q4oeehO
YEto5cYHM9Qt+IAuoIeGfO2/mEjD5wztNR6T4w30XFhHdvGBPP/6X0U/Hyu5l5m6
kWUs439uKkq/Eg1n87zrupRbAUsI09+EsGQVYSoolaw4iCQ02h9mbisZyIAfYnpf
KJ4e6ymEubILs+9JbCkh3Efx1S7FTVxSyPE8S1Cz6uZBfjcSZHa47nNMEghFedy7
EvMwzH3O4BmNQm6gAYLMA7ijBOcAcWzAXmqafwseX6HRghjqNAGee/y/eQyyKZcd
PyIg9tM1L4+rdcUyX4et2k6MfFisMJvTbU4HFu3hCQplDy0yFmdoEPXrqPxCB/uS
z1tITVscMHKH88e9h+XWJLJxytaq/9JKnPwtAet+Uk5xJjH1RjzLRv/Na7EKFicV
svmlI0EP5B0a/GF76Lf4YvYxyYSIewukw8Ateqg3Zsl3JyiKkCkJvt79GgQZVzZt
vOV7KbL46NPJr1K7UyKKgBfEAo05sMVdxHR0iKAoFar+6FH5pm+GNwMihTqEBLHA
6a1yfskZ3Vb1njXVLRO4Yt2S5wvVWnkVqwneYEvJoM4AYGJqiKPmCaZpU+jDmas0
eQlVMDMXLYhbYMAK2sUA4jar5POQRWKEViGrRT7lwhfKBQ4np7vrSyBl9kOWieLN
bPocO+k0Z4ZJQniCvVB0TttaFZOL1pA8nzsWJdFSTFi0myxo1ESX0wVGduiMFEE7
YSLV9FyvA8SrQtgLE59DPVBBC0GC2VaQcfuQXb6Z8JpLJr6NjDvfkXVPbrKpSlQ8
QM15yaOBuEEG68HzcSuoBAFVSeNMkjwbmhkwSuICX0kXQM6uX0VVZ2SQP8qAvxQE
Fbbl8GDlwWbfTfEwtkYTqZSB+A81/KDeiMVVLoCUppEpfFBLYOEgCbCzSsmAFYCZ
g/7L5xuhJVgNnTI0dMgsPvFVLllOZ1iLKpV4Yxuoqeq9gL02MU+N/ekNPqgt7EIP
o9tH08VXXe+SA8mZWbHmLPKg3EPRT9+9KjnIxm0kJsqJ3bOnPQ3E3z+ETP21k++p
y9jtXlMHZUhO0GHLKcmRqNXqBzM5wrYs/MJRR/91WQRW+d21hyJJ28e56B5+FDVL
KvWQxFI8sXP8ttOgjRnnbwDvYEtoUWWRdSaU1VTGm3b5L70EptZYpnZp2FPGJMZm
1Yt6OKa1vdEn1/WD5jI0X0eFxM/qkfaNcTJ3JZbKZsmOc2yaVHAjyqnDxlTdzZdY
IMWXJ/+uC8vz1AqRfosuaZEjLasIoMFyWM2U8yRsRei8s6wfxOJgc7u7ldvJu7T7
IAyPvvpj2T+Atu7C2l07KjL/ftQCmKsuHYXDDMGOBpa5OzEahnkQLSI7hGoBcShc
ptdFR0rUsUldXsFkEpFev2l/f6bwojICLMCCNyY4KEvMXtPlrHWSj6YLjSZv71EI
M8rNmk0RqSzdpMb+b9iB9JruezXRYtkJiZnpx7Gem+RzpmaNAe5yaQxc6WB1hISz
DPC6Vbud7E/v0CLC/RNxKS9b6IZsThxkJDj5AWzSI8Anj3jFimzibBCbpp5KC3pr
0658D5zqhm217ldmvwf++qlcRCzVK97t0GbTCc2MJGTB7MwA8lHVXjfqUSK8JR1s
vHChxHjs4GyNuqdMhBHSDItbALiG/cvPVGaB/3tDK9zArYXOEY7SskyPPbeCn846
SgwztevljC0DficuoBYoo/d4bIT2EVAkesiEkyYmB2LC126sEnlmUxyfRnsZcExM
g+J8aDm8RC5ecKHl2z6nHu4WQPZjJCQ9W/Bnp8rgzASyw63D+yZIpc+qPZ3onA+1
5BgEa8qknYLuPJjmb+Tpq+wcuEm84WaiiWI3YPPxPqgdeRNywPZEsg2mAkOdrolT
P7uLo+dlcbCB4Wv7LWaMfPuyoO8RcuPkiRNSELGo98FyTJSg8Wkd8WYhZsg0irh2
QGHXtFfg3F56onY3DEm9XOFaoxubMe2wXIuLmqxtu+yibYhGh8eGE3AxaqWsq8ex
WEMiDxhFi/skfN36N8ULHmy6b975V5RSvVVCpr2tGZ4bh0n4usRkyHp8+0KGRlJv
W83D15FC0uwgIqvHz8qi1l8X9jdOGJz9ZKfZ2cWGCxiKalamSwOOIfb+ifPEdCFT
hT8Kp4G8wS+27BYylNl93LMSBlGe4VWlskunquO9RPSdDcmVS3wMYuhFLjobBXMr
z++Y+OHFhVJ2QxlyYgqR4svo2DnV+z6Ij9ZxYxdgWa8un1hwX4ISfYAiPJxDqKot
kA5cWTEgCI1TI2OMDDrhzQnikkfkc8HHluunXS96iMeeMLCjNNZ6mMknoHTa/5aA
VTytxoX55SYwYGEjUu49gfPdX9CwDXhvQFawDG/z1sJ6RMF9Qzc87nQ3Y6LEfzI3
480g4oTsfvflnC/RqCj8zKiH2kjkjAnwDHfkqDQQuq9LXaa4xKjGXgf8YJpQ0+39
20aSU6shOhASrhswzIUZ+nVTMWpH2vxOn7CyeB9b4Kf9WvajZi4/5GX4uqSszA4A
liQrfDKPD8ZFP1c/ux9Fn9UkpSjtPmzG3Olmg8btgYQDJZ8j3AI+6uPy1UnndHvN
/r3/z7iyMzSNB0lPbYvfYhjtRt77dSSsWHCo+eA6Q+7sX2Gqqle/1jo9rrEPHoiI
jjZ1PNGhhl6am0ZQc9YtCpvLDavDm6X1jM7/LLkKEsk98HIJ/tWSbPOACUOCWbuk
cWc4XYsrwsvKEsuLZz7CvDQpjfdkV7MEgsG1q4p2uKVxhiWWO63dZokV8yJ0+QzG
xgVLfnB3v7a1QRGX3qn+6DEszxLm1HBKkZZ8Pf4Hfq8BT8H0myrFM0IYaoL26cX1
FePdl258m9mPHZ0Loj+4yWw+mAE2Ntn22V+2bEWonsgTOgN7pDA7/HkwTWmrFEaG
jRgPJlg8azb2OMD+KAT6CUhWbryDJWk1Eor/xQh7muRvuUPMP9YuNpfdrec3M/DE
KlQvERIYTM4i99nv8F3JCnT10va+aEBjMtIAkxLE2RqkgZzTKOghdS16MItD8psh
/HB86+dS1yAFM7AZsWrhKIJl8f4XTLWXem1t0S/kWsQ1Wxd8ryh6rL42ztcTytDg
9EgmWWgLJWqvtTh5lk37k2UjhJmU0Fy97nJE341p3qEh/XvfooEH4xRNRquwXNgh
D0fMZ+k824ug2wPW4yDDNcrKt1nNhFKBQ72fHEehhV4nPZNprA6yHUwAGhkjL1bM
f1nw/1GFQlzilos4AP3oLam8TTd6jyzaUQDVvce9ejPs9ARLcEewPFvO4GBmN4pH
SouRROyvV8o88h3riMkfv6s1HSOZAK6FUeCm7yAXqoKVU5wMLOAfmncCVETB5DiQ
zQTv8Yw9+WvaCCXJZg8y7fkvIF2BXHcx7AcKmmR9ADaSo4I82a6RV+kY/cIX8K8Y
3G8lsMIMfvaMxZCwpJ0Iim/sB8n4gCZEmHDTOiUU2psvZpydzkyL8w0Z7IhsziAW
xAFvqtE2g4XOeMhMPoakHx1fnkePCG5HEUqjk5Fd7FbWYet54AuqEni3ZNYp3xRC
AaGwG13VrsFASnrea1FTgPa3sBkiiWiJxChXnoDmfq5k9Bl812iEDumsTLqEQa4X
3fw/Z9oXDV3QCMq7YPhs3fxaDj4v0AP5C+XvMgI+snEnEXwc9GGTaFDnZpkFWSln
AdqOiwPMJsz0QLRviaU6Z0G3UDEu8vhRIF9F83MlXA7OuMYOrEvt6klEC2cO+x/q
USk2kDE7xZe9kt9x+DyQaxhFh41O3OMZxefvF7mD9Te8drMG3JkeXeGug6SZRlPM
qHJNMgxiVNpUarosshNdKrXBHrNreKBvOEcWwybuANR21RC7M2dQhZs8j77LumVK
Tp5IXZ+E8nCxFegQ5W8NxoMi7ZL9Z2UXqw4hiZMoSRQ682vr8FRFbK66hu6k4jWs
9QFuBrW3Id8fRPhOHWmjf6z21UGDbtAzpteVhwyP7ZJrJs2+2I7hN+cfqtSFu+MW
8mbD7Fz1qyiJZcHDIETFw2obctii8OPYRU2GiuiuxWiPnHMEFReJGHpWhfJFEb1A
l12FoAebruWcZly9rSATiRWFTmC3eGL6ATBA1mJnbfRQ0RaoKn3eexLQS0gEpYOw
ryFBXePFQ8DuuCsozI8tNf7NJ16mfze9a1brIU6ljUdOMlqV5IzqxQ8q+BsRKnJu
UGA/e9Vfl3kgm+ud5+/yXz2upNzhaQZ7NPkQeycgVjN8BGKLBvoyFDU4i3v02to6
cp2YNaPr/FGw5DbEtN1Ck3y+vEyM8GsHLX5osTxqJSbpzkg7v4KESgc/fWo5vIlh
ygYuGlBRu+hz2rTf8zmGi3AxC2fLdeCTq0wy+j7vKUmzk2fFdQeoaLflhHAlLkCz
UBD2geGmfql7lTbw/XiSsqRMV4nsTfaQbBud20Oi05ggfjc09/03uqyFrQj+ivdK
DQ8e1QWThlFedBjJvgRLErcH4aSNf2sppGuL8zpV5OklEfIOD7/xG87t+S8SRKpB
8RGNGtIvE52LIr70Uupj6/j2Yl+F++uidVwgnnReEmYwccN1SLiFZ288q4wvcSA5
O56mEwuNFqDyuznsZU9gEFXGvUBy9BvMVbq9axvAQ/DKFxitgxCKBxObc1kzvINN
gdSulzjO7zVzqS9EyH5MDwA4VnvdsNAIO7vUpcIgfUgginVduawCSU2GMQH40vm9
oRccQm28MqL6RIwwRJX7dhzLaB+s6atttA/nc7TUZu9HJDFFjSWfALRuaQgn//GP
NokfErR4QF0QqBUciiQL+rADrun1nUYSo1W9NRCXBIINgbXdoo6B6/OUbWARrbu0
PQpmKBYxDYLZhSRD0vIfcGbg6iuoQxu2K3G0ikATRKRlhAjh9+KkTBfLHZIzort3
QePEFT1yv8VpGnlQFikGVBKD7QKWvXOI6b6VePRBBz4R2oOC1KRIeWBVRx9XZEAj
eQM4HOpiwA+htHDvNL7aCJ793kaDStBfIUB3vqBU8sfuC5chdTAs78LNQFVH0+6n
Xzkn5MGu2CHPw8k+UzI6zIo7ASZWz+bq+d+D6kxwpGi8oQUcdpGaJTOBBGc05NqD
nqJPkZYnwCk0n85u63TPVXSJXByHA1YNq2WPjTUUPkJWCwyzvxfCZ0TuZMQ8LT2/
+/90ET5b1v1wuafUcxUTminr9GPhHtN7UJWc9EYacRUvhEBW8PASQElHZf380EPj
Tv8vj157A9eunxJKCdvk6hKflri3pqhtaXpuMwyMX+7nkj/EQcGadtrwsYIWDRBL
ktFZhuUsSutR3SeetTLg3GR9N+D46Iwd7n43J/3ZY7srNGg5CerIg2K6r5+I8Z7v
tjsGyqL/d298Vps77RhyPKgFIze9KEvMJEELwP31jeHobaK4SzPAwovQUgqrJBGf
ZQ181pAINqiyzko9xRQohZdRjJ76iK/RdOmYIRjMjJzd/HEQfjqCbJBmVX1aV58F
RJX9GghzKdIipKSssDJUei69vc+B8pwms6BwAiJi56CcSRH0hcYtfmDuCvm1p7Hh
YPz9LxjM4LnuzTmoViNjm0MbttHywNKkc/qSNhqcsFdzTaSbpc7os5snP9Yidgks
TVtyuJerGQsVhGRi6tpLA2ejepqVneCMfkpBXY4W0xSj8mcBSY32+EFTeXWdbXZm
ptQmmWvUEaVsc4TnQ9Pe+XdGemmG/ly7YFf2N/nDkcKm9unft1Gl4D2RcbES/D62
htgNKvNwnsFmoJOh13cD0OF7lwlEW733bZgwxQOwnOcdFIKSh3kQ2hrbZFO1lQvq
kox+Agd3FGT6pz8F2me6zCm49V4AucWQZEsT40VNzo07F04syqydEAnHWAMLbV9Q
CSnA1/ar/u0ByL1cwC+pFzSiNtA4N85Bf7oBCvzVk/vhC5+2+oinhIDgtwHBBiR9
AumNI6AeJzuTnN0kcGMnMYw9iFZNqVhDaqetd13jkIt9DHjNCMQqnUd/7JmKuCVj
Rh+fM+1QuTKjkb0WrvIXhOgDPsorXEThWdShW3EdlUyDhJUQEH7ZK1XuR5XZ1RP7
9r+5b89PSiOd+eKGoiEug0Tfun6xAoG0i5BewA0QqlLTNjdUq0+/Fzd2w9IjX0HW
aQQOFLIekmRuKPSGt5PRJ6WUNsQ65PqippHmAS8GE7GJkSh7zbCBbMVvjdK+3qWd
X+npy5kNW1i2ExcDavEcySHA9qGb+Cm3fNPD0TJD3f6YzpvUon7o/Ap7fn7QtQsJ
odFr4gjXVkqFsAKMpjglOHVhXay6C3fv4FJVtvjSJ/MZHWpiINN0L+EaG6KhxF7u
F6O0tB+spPDgIdEf8GtqMohmaepU64R9bRZCqHGz88VNr2JilgIDmS+e8JsPBloi
yO6ddbsZL/rI4rcT9iY/9qq8P6rK0VyhvzD7iBlPFD682ygMDgscu5LjvWwinARo
hIYaV7aw9YT2L+nKN5DDV077maTXFHaUIFIrjJRIhjJxjTPtRBEly0ANaDFylM/a
LM+WycMEgfq5Y96v3RnCH7yx7DiHHoxJg32HsXfeGPte8q2K1pH/BhP9M+RSzdLI
nXzaHiErLUhWj3jzf5WOjcHBRc5NKr25xHJ+iI6jiIoQQ5jkSLkx4ffVmEJypNqh
/Cixijrm3M6bI0v0XCPlJ0uqHuYjepM8QC0NPH8YYfKSl/UYW7aKUzK+irIfBW04
d+6gK94Zqdg6+pV8X4BlMbLXQQqSTfDFgfvndOOzbkxjsLIRXlRY0d4a4Extivft
9qYdiyxsKaRTCfqt7P0+FqcU9r3IRGjdin1FDsIp5WzcsRyRDqTw4v+XwZReCXUJ
hgL2nDRJHc1gJJm3mP1XvMOU8hfsg+tjn/eNvANmdnZKMtcky5v7DKO3+F09aBw+
XfOdyP+aNNsZkaTRFSh7zxmtVaW4LGUxucn7SI/JjEgd5K8+lB9zIxom0JBXF65B
xSApZe5d8bNm5pplJQKlhBjVsf4ojfH2Sa4PStBHBMCd3LxFT1tZ8cO2Q2Z+QBul
tL9zhGfIWnXKtQiI4B8nSBjV2C9LHwb5fKkNe85ZAhcphLG/wFRiywPR8yTErD40
DIKm3XNDPm0qW+ZFR1du0HWCh8f5/vP4J7AggUYZGRqORrX8X8DoPP1FtpNCHRpa
WvfUvZ+4YoTP9LUhN9ZjAp+jolFqL1qTpaz1f/5dyb+Q2e6+AzSpBt0frUXCwYnB
Zr4mO9S4F7OrSNAVcD97xuyiI7m09J1u2cBaBPECqrq29EMWMf+5leUVJJ0cqsD0
Gj5lQ7hLdHJwziypd6ynvW7wbrl83c7L/vcvGOVwFlIoDZMRKsLFlfYJDobzPGYq
GXo52d5dyuVVyeBn75m1a69rFI+0mbetJW2yTllS7JmU4Wb+uzVfpcWviG3soBkp
GjHJyeRr9WfEtKZWDkaG+WDwBGouRs6i2uo599o5PxrB1degoLTkbUqV7tOcIvFb
opiCSRtOp0HC88sC0wFW2u+c1to35DvbA/OCKsoWEdKVq6m6YcCclRn/edrDitRC
6svMFWqKH3tevgCqtAJhXlmynZefPiR0bLa04JI4cJjE1tXI3UuJeVrYd+cjRBXf
bwdHfKf8qa4xb8ztpJHFZeJXZPMEqHjoFzwJkKvCa8SVMSDq0HRX2Ub7Bfm9AQ38
vM9QUHliTuyQhrqZ1ofSBjbEAZXhiztsJiipIUJ+ynzFbE9DWzyZfC6MjkpbyyT8
6JZFG7HSxGd8Qw0o/VJNkcRd2iIF2IRIb0W4vRAo9A32Q5Dx+qUWufJPVXLHfQvn
rySVo0CgHv+k6ZQbYYQqw/hqGkHjju5rH6V0QYEAhmtV+cht3EfBNCaFpwz/z4C/
3k47uoCXGkWwoRSO+2IZqRl82akYzCkLrrT+NWf9DbGzXkPW/PJW36y4TQClQBFv
AIzD480OgaH/EKM3p68C/fNI82S0ZpUwQCLHfl5CT6VZvAqTZBRk5hgKcXY7fT4T
Ia2OOn/PmuzwOo/YTn/0NGmXOAwUdddKx6kGAw//q/xrhMRPthXFakpIDlJqlBG+
wF2mwSPom847VxfngNxCTmSlTejYnvLr+nZF1eEp8B+WtuzE+WKnH3NYCYOedcD7
zH/skALDHaYEXH7/hArMTsrhTNo5Cgpr7BXH4rUWeAEpjla1+GPkZNLA1emQyTpG
UdDirhfkO3b5Z/PYWUCpbTpsFwSOywn5QCVcM4QDXUPAul7vTGi1URqB985W+7Sz
y6Nktrf6KEytK36Ikqtkvy3WQKhQy0zvmr93JqfQXA/um4m+JC5aeK9L7fUzqIHP
IJQ0lwpXyJpeEliU1rYw9WtLqushMYUQC8EcdDMLpcjtjtA+CMjHOJmEfU9BAV4T
eDPIKV68lhgQY/o4QsX8WDRZ+UlDOLbSzP70ESpuSkW9ai8fdBlmOiq9jry5BbjX
Fz7c9Uk1tntdSL8oJFe62VN2uAJbbdsfSHuRO3tZy/+fqpQMPzg3HBPgInL8SBxr
24mz72sipRoCShFKmWBQ7+EkjolhS/j2VQMPXvwPonCFsZbO4xMTeTm7JfXB+CQc
amvRWJGV1Fd4218QjrWtYwxITDOzFIShCmm/cwKPtvi4CNZEHggSqKPvBoP4IM6K
AOfsHNuupSjp5suwnuOcL48U4GzBeS1LneoMDrgs+AKx/BrCee1uoDW5H04b54Ba
bt9xQBhbQOdJOMBKNoqj9uOEDGBsf/hnvFFWr0wXIUUAiRiuNN4RnV1wyyBit/8a
JNTHBH/R6AXkd9zTxYEp5uij0VujQ/vpcjHKQBKw+I64O66Ky5Ra9CFrT8Z52jCR
5kaOxv8R6BprBVifmvEfEXEW3t2uUZqzW5heYTt0AxrNEA/HxtBzFTmXGhYIGhw4
qoqGlnErcvDE9wrUbLkrNX/9RUUrotdFIEGxMg6UnMhBcRQYuCfYTUB2KRcOrkuO
+0OOkJ9bkNZNkal1DiHNt0PZ54g0wj9iZUhnNgCdkOalOVLR488Tv3VaMifGRDIZ
KdiDZ3+CBNY7Eam26aauW7ZkUTLfTddh1KN1lrtQwly87kxuKNF6zJ20EtWkp0q7
UurS+dw3vs3ZdoADJH78ZRso2b+pBuT/6Gk+wf94hl0c67lncGftN2Kjbs6Njc8A
hyX8oWpLHyXci9Ko90LGUodjTbKO5G3t7gfHUVVDwmUhQUKOmg7/rggdwGW1TJwd
XcVSNCa63LJvvjT/VdVkIus9o71niW9RECPIPISbDmwCLeG4nynyPnAMy63U5GDc
34ZNN1XvJAUbqXyNaU5BHDGg1TOtcHlIGeIoKr9LSXFj8zlLiILA1goIYwQftMSF
3gxpVonozqZl4VbzLCIRgxkYg1fG8UiE7jTUd4PVowgUolrwzLGHM7vePXhk++57
O8kOgu5cYDKpP/N0zOtlQsDOiYmB8ujnrFb07HplEQyyNNRz0KQXzCskNxvViaIU
wfXld6tFBoFnWfEDATVIgalSdsgv6Dky7CdlHanviIbT2as59O0rEiO2vIHz9ZF6
gMWCqCrY6UnFjmzgxip2gw8KAFcl1xKXJWZy03Ora/0nCbTeq3ioYBAfW+xOYsZs
VJf9uPSQ1E57e0qG4Ts04WVO4WkDexYV2RSjL96ZhG7mFgoWr+QtfDrhl2v/Nkn/
WCa/6k4zv5Gh6+vD4s3Ne/llj1M3NxvYAS5iT4Jmu+w7XP+3fSQrJuC5Zu62vRI5
awq27PYbfo7XzDY/90I+FE4JIMviLIdDtceiufjWZ19m9N/IZl6dB9TZA3cch66k
6k8BGHCynCGmIuzoJfDlbVSbkJza6PUyLnkT2HPZe6sIed5ZVextd768AqKZ7MAi
Ns4H18YZTZsaf915Q9Ue5B+P4AuAYJGau3eRQP+d1BWMKCGtrh1B772UgPqhN1bU
ltmJDAYMsDbJN9SzmNYl7gIAkAR6KeNUyDnR6BeEit0u7juLqWJ7GEPVR7rUm63V
KoHk3jNertVt64fHZbgTdFNreuP5bKL+KeVRdEtYwdA8PNCtY/6RNuLmhfM2gO8Q
4XlSBMg4n9LD+eIgBmKrHcE9NaqpxHOcm9uFOJMtL7/lMPAyRPr+P0v8C4qyuFGk
sKJtGvBcN6cDIaOlMDM6iih4qWzSd7UwjK9Suxktug9RsizqPl/0aThJbkZNettB
Kky7GbDAQ8Pl6MYXbwGDNyw3KQ+qm3vyT79aBdLpRLXVpyBnfRS9cG5Ap1cPQhOh
79p5QlxkDL93A1LtCSd6Mx4MFtoRMoK2bSxlb4LuxgBMcs6+WzZemtZyTZQkL/vq
vaxn6HxpdnTUvKtm/2vGIMPwIMK4JMSLZqmzALBfw8yGEqWsrToY6LxrtRpOrNM5
Ei+qWcldT6NSYujNVqnLrMGPRn73bqAS/C5pXQda69TZodny1zYwFpFO7fG/lc+R
UhJpT6qnfaDEpmSmu9LLgQpaLrUfMeHODllhbaivZ9hpUS35dphhFViIo0GrvtU0
PzEDxrnaFhcAOneTNhxhje9bEbTLHahHtI+ewTb6a2XTAp9CGmvO18NnL/p6D5M8
Q6qNqj/0q/+0UPDxTDLDOZscQLxseYC+FoT5zw1srQtD4pkrS7lt8gtVfgf8rGUM
Jmc2ZSQ3hmV3qFOT3xOCoCycNNmwrDweZb1NYDmItlB8ILN+0oG0SzTpUqTqZxdl
fG6UD43r1QNXFc/L5vMj7ZLVctNWpVHf4HrOGLEMwfpg20laPNU3uFTfr/x3CwR+
gomqZaYMLuhfrv/C3PWH8Jua1aEh8bC40wmk8DDqJv6umEQSgwS744Qcyd7WEKyV
Ue2jglDF00/ILtnmjItNzR6sPZFECc/TbdBtcbQ1kWfLVTbMnDUUcGClkfrDB+YU
kzyT/ACMKoKm8kih4TnsDFjS1Zc0qC29APl+GfbPdlaNqHBpoOM7Ri2gfw7YyS3/
AXxQeqn1Sb60VTOexmK6zGobWheMwTHAJLZPMv4gURzUym6vlCIVPoLoxNcHeX/f
aonzU2f2N1HT7U6rMBXlKrlUBSWuqR1RYqf0mzLk3ioV+mU1MMGiKpmxdWJ9zqkc
pKeJvLPBKiR62yIOKLSyPYTgWX/ozF0zR/76UdWOc13kYzRVU4f2E8mH79ipkFWa
7J03RoFM1H+Ett+BPkBV2bmTUGumPuoSl3swzG8zUV5RFUgPWKcwRM06oy/TZloK
EaTICs3XrYAh9IJVYXmFsfesGq2zLv/GNRFtqX6owEdG4cSz1jKl68A8rrwdjvmO
AtHlijvOARsc4M1j5HBcqoE/rI3v2WjACLBPlG8s/xvM3JkNm9fvBmswb01zoot2
joXZ4SbYts0LdRdxI7+OmGf4uTqVI5Eshi5mScGc7sfBuiHa2TDmLBl6KGcNqGMb
twYZ4CyXOVqhed2APfaARbZjY8OdlMf9zDA+JR4RvZuuI8h6gQ623bn2OfRz8ara
G8RK4N5hb5Vo9PUymiyDxxLiSB2iUxFaVQLn1h8P4yHmJioXUTyphpJdKwFg3StU
BT1lYiFzpMqm4TCuYlJTz8wl8dj9QCbl4JERLF1eysojT0S/gOSnkwzjecTShM88
g1TWP9YdBfszCwsLqKbJ9WUl6eCed4W44I8wi7dUE5tULOVSSMlC2zrYvD174P/C
4kuPI5t7i0q7FR0rlBh3ckXXBg9EqJYUV5MHvAHA3C2SggdcjTB0b6Nzprv3IQl2
1V9zs5dXcRHajITbX2vDNObp/wTuJYk+i8cmmBl8z8GatFLgn41Qd//s3cphebsW
IS87L17N2bg1CXK8flrCsH5KMRKf4sDHMXGPzRPpICGizXwENFbaa7FrOPNZDAeK
Y/IiIdcBPJWxQNvakNiYcpNG05EZOodXmpJHWCqOSP+CzacCTazef/rJo48GyLft
QJsWrqfFUDvc8bzVuQ7k9PsgEPHZ68kU153xTjHTJ+XwDvEYCUXeU8V1wkYEigGe
TAEwWpo3dSiTBUbqJkNCjan15riQdpD4HCrFy59WGsT99v3ja2v4Irpk42mTAeYV
S+h49L/eDXjC2qGTfEB0mGGoilZn93zQeMlx5dfJeQH72EKvuGe6D8BF04KcvNSu
w0zpji6ZAdPyOCfulw65ImXXcl0QB5pnjNFNE+Uuv7Q6vGyqtwZC2hiFAYGP2kT9
4/J9ff4GOC3fP7AkxkAF8ejGJhim7lj4CCsiMbsmrnu4rWz4WVymFtlu1Ba3/Ov3
ol88ytWWsLEL/iXAZFVG5WmDnMLWj9DINVQ1S9z0SkbEIOziKyAPOrPokj7S9l8d
nHMOgPxgP11ndcSvXTm2HwNtGNSXaTkG5SKDxmUgSER/7aALCG+EvE0DhcWS62aJ
yCTI4nIeRBuN6LS9iPKRF9dJyK/AWgFjb8gcXs/ChjFSCvE+oWSKMVCDHyn14Ryl
DZh5ysZxxBlmoDymG3f7qdOQ4kDiMEQ82/3yqfNHA4X/qBk/5jN0ljOgv1x/iPO1
v9EeZp20vl0+TIeEFSm/aL7LWXJH372OFaIunESVa53Tfwr4pKBMltpM/gan3aBc
fpv+z3iPCk5D6aayEO0p2USjP6Ybd0uCh3Oa4e69y0urnvhtPz+qZSGVRSp+HJ2r
4M5K8SDc/rVmYK8OeHmiezW3uhTEOGOGEo6OLO4PYutnJ9UcmzL9rvsHRZZU7q88
+VyIcogK3niJo7hZsW0MPVvOsj5ZOMWAzSlOJeLJnQ3NIzSkGMRjFv6L6TUbnXc0
8s+q5ZhRc2UMFWzbM0d7Go5tYdWko8JhQQm9unF+YkBIwAzgGvdfp20iHEbe172B
WAkUV6zNPjqmovmOOYTOYGh/gi835EePZUo1v/4BGNV0k9RsP/MroPzWC2ub/lbt
B2g/tnkIBsl6Ybn92oPmA9/h4xmRI5oU/ThGeRd8CRd+gemGfBnToLjtihWGEpfV
P4H1b6uoO4rTrWAx9OkYKXn4+W5brTUv/eHP/0nWF72BcJEdRblARW2iIw/rYIM3
XcsMJeTZXan3UA/5B2qQ5n+rGc/Ggijho5//ToZ+Zg9Gi8h7YzqYC3Cn8FFQ3+vj
AQ5eDfzV2/j8/SmJqF3s44B6/95jj2kN0vlSoFjwyIvNHBBxJErTylApafwdghPd
+qTyW/5wko69fLdqDXGQmYA/dvR5D9jwj6jv+riTHYkvCoYKBKi2hjA5UXbQ714I
HUs7qUvKAYf0kEp/AZV697v7uo23UjsJMFhlmT5MK9m73oj9DyQubpo62kGtvfGy
immTyBPCRgVJE3TXpujhw0OZmQiqDsxm7izFkokPTPMatYPeORzn0a3TjEUO9J8B
yTQXEasWySRuCTmrntPszYorfBW/MlWqe+3iYEWJtiZ/AWD2VxyyQG/lnv7VkHzw
ZqETKxjS6Iyl4YxtWhH4lQMJfm47q8THldAofg2KzM7yMobRrZea8uszJ3LT9pbW
srbqp3q61IkOqZVWeRYE4QuZE0HfSqFaTSfkRzXG4XWMM0Tza2gBlcxn0QEdvJv1
FRIwSUcyM/kKsZ6f54lc5nb6+awigEhK9HwY8/Lu7uuOF/fVTHMsxgtBlhb/YzLp
tOkkbS9lS+E+5HmhvkKz/BECTfN8lmmoNv5sCQV33ugqHXoovycDbRD/Bd+KEjWD
cFnYLHcYKJ/+IZ17e2vNEPI2f3RuGd42A3dvXCcimmKFfLb8aLqzi5CPp54bYkI/
hF34/rpyDbJClNxDMImkhs14TWmzvy0N+zuCtuh8HVqcVdlt/thvfZail1Q++maY
BmJCAsa1i3ZusKzHujq9NR82l6a25qqPaYmfyyhBScPFByOGTEYPJ49MnHSbwdyM
6cgfUmEH7NtnG+27MpRmX60trdorF6Vsivjbc1W33n650cw5yIFDWTvraICQ9idJ
FaXc2pODAyMXP8OwoH4jQRsegeZ/aSHgsqhJWaLcmmHacDKBXk4GD5SsBrtDZPGV
27WjwX7sr/Mt0Zh/SXJmfbwQRWL+urdwEZH8Pg/gk7V83b+yIBdjRUOmeiWQA5PB
ZsEQbES1ox/NMAN5pW5Wpe0Hcsxdq5dL4wGSWo8+Umr5Z9jMkvHvNpHhjbBTlWnb
EfeMM9kvWTisxegk3uX+Hcjgp5Wyg5fYGWnWDr3purbswEfxbc0ZfIVK2dSSAd8E
U2RvwdVysshb+5SKvVDHp1aXPZpyR5TK/3uKDphoMkX40knjo4Ky+7c9WK15fmfK
z2kY4gbMxiG4cnzbxbd3BWSxQSkMRFQ30PsmhLJO2xle3wXVbbsJI8e0xsb5MNly
gPARTe8Efy/262CKWvbr490Fn8YJvFR462ZBOyccdcYNeVy/zgvS1Jo2PInN9jvx
vn5oyy/m2DhMB7Y3uN5V1AfZtU1cCxDHlAFZKkONQLxKdISh5MiepOo/V2eV5W8h
sVGj8S6X0MtixLHcKPO1pbmRWbo2BL3rJ1qwQbI1AeghNr3e57pj9xAz8nrVcYnM
7upT5j6rwIewVAorceU08RoNVSMOPXu1Hr4PKGDNnDbPD/xfe2sFgAN10gA6Ushv
oo5y/oHnASH/y1ePMnpnUM0PtVzUaS5GRb9khnxdLjhnS6TT/CbGyVO49KdLucHQ
4xMoMzLRgE7ftZ1hlcy/dGe/ph8So8wg2C0Liz4H6RV28DlieLUnubGaUcYLOVVu
QIUg0hPEcJ5XywHkGPyuAlF8Fmvqcxo6Iik82ILmbIfbqnPZn8TpZvB9wPgXAlL1
mzA915EeFRiVM6Qslbz0Cbmf6AV09yF3tt3o9t7RJ3DnLtIfaxMbcOTJvlZUl3qK
hZoi34BFtm2DFWtvv6WJ50SmmxpxA7whE+omPgoytli4sNS23FZOUbzD1k9F+qTj
QU6hhtZuUajTZMbr8j1dPq/RFS/GRBfp3K4wqG/BxzB/wQ2yXWA1Y/Qfa16cYzFU
NTf39OG7Ug3qDuMev0E41RhFIRxcSLoiHOkKd88ZkT4+ThC/YjIstLajfxOPnLex
pcS10WYwdIRvq23bN6iEvjtPnHYg/riOyBVltemVh6x85yoyE4go1nn6fwXNwGhS
nDZyDdYyUleRf3d6Z91QNHwsE31/fhfyL2hhSH4ul8/yel92FI7e95L1pgnWJeaz
mrhxrz485vGiTOrPTdpr1omlKqMfwjlYg1l2WX2lKL4+jaQaz02TptTx+4eNDTeq
FhgU/nUeC6kxw1CN92Ihno+HLWHyG0xy9/XfSzOUbvndGzo/fujxN4vg44xbfhgr
6yOwuugB7wEgLmRFNyy67WBfGxeWDMqwT44f4zJXMtc/053hxEBNRwp9Wm3KVzmR
0DDY0+Mj+omRmfTuShhyGdoZKW66mQmAW6aUSnqb0+wdPHI779chvcYHJ7kPOKuN
qKgmgWusS1YcZupUpb+WA7tWBqsN0bkwsi3pESA2p9FiD61cYDEisQzWq3+kGDnY
hLyn6IzgovTJP62vv+lg20UFUmuO5MSMYCz1lBFA+NyMvBJuiUQJsTdHbTU/YvKC
WJQp7SaC1WEpq/a/dgQPt+cdjfRmtnaXR2bnzeDv6621/8c45HXlMnCXrj2yarI6
8fH/uZMirgEL0ekByTbfRSQ+tj6w1XSjH5DBqwarB8ozLAkL4IAJpZKDUbOFiKvp
LTypwfmaVDfpq79SFrKB8ywiGzi1Lo9v0DptXVSsjW+Yx54+tMFheZepgdiZZbnh
WpWkL0IgIW2HcaoohIfrk7SIZm5nQqddSmsnE4KSBuFV7xV6NXWzzHYfSNmj7uUR
sSBE0Mfpf4zKPtDsS7CIUI3rRyDV8spJPC7UYHfWM7ssSRJWGB3/Nql1l5egtior
p3B9piBKo13BN4EJne5jjYumY4Xa+sWBJG3Dc35ZTeWpqG+bL/huJix0KLT7ApvC
668Uli5x0761/S4Qb5S51jO7QKQFRjEVR/weX7g2LoERogGyg6jdr3+2+7kIG7Po
BoIp6eQp70AzSkUgR93nTw2J5yAECsobCOjFsKuNjNqDDBcOQ+U/EgNqLMJQhKqJ
VCUlS+vOdg9es9P8Q+89LbvMXDTg8kV+1K1XSyfcTLbAb8rUYS/NZgEqSLRC1A7Q
+5551MQQ0dLu5Q3JkHUqGrgf3AXpgw2vxanJZ0DK+ECdFSe3MtnzqXVNcdoq9QG+
WMsd5+ciOlTRK9+DhDjQUn/eM/n6Qr1DD70QrWPQ/VhhMSDeUK89EkjIY0BgFA+K
gC3jA3Td893h8sFk1BJrh0EAquTMiT2wxxl9KE7WW/fYoGjN8qXOwHFSzgQvUkdQ
DjWLVZfyZAZRyF1GHz1tBgs+5XexHr2gKjt1zgA4KMuOPqI6XqkV0n1okwif0TQE
N14VZf5OBtQaUHpzbXcy4pLvOIyoDCyqU593/7JTWIPUFc4rz79uYX4NhQCbXH5H
HNif6+qexzLgCLlcICSkCE7kqA93N+6owyYY9T/F8LCh1NyUTg8fx0+xPtTECEXg
K9na7KOfS0e5Imy/wY9NWmR49KNAu4gjfQgOjOJFFSuASnk61PQa/LsUGJutwfNG
ctZA9oxo7dsRB72kMa/C0E8snyBPrlmT+uWLEag690B+SVyqYCC+/r7veeDdRnx5
SHyKG3Y55J2sAKM8Ae50VVADKDaOxNO2X0ljNdzsorhMb32IL45tgMLnn70GhT1N
J1LMpRQ8W9160pv7bVc2rZwHstpKvs4DuSXF0R2Mz2070PnFpv7IxaS/I5vQg0F2
rhUVyU3kwtSpv0BAMNfPS4gwrqqc/LC83VVnXpDnz343OXxqQ3W0NLXizT4TN5DB
s15diOvYJH454sCSVY5i13/IAXRdtjwOHQiG7XtMjea4mGNcZvXnYyoCSBAe31hM
ot7dAiqNTGgqM0tbyTLikpnHYPfxsTEG9GDqUR/N+uQVC59Lts1Hv6+uSDvyMSW9
6AlfwVUdGZXc8ManTKGXLBPl6dafHHbX1JzDONgoa+WaQ35ZfT+3ToPWNXnRCX7q
p18MjHbclRBDUdckjfFGfsgbr2MBc6tnfK+wu4INLv9lfEKN/6V6cRgvJ2gkwSAE
0pyYNCaT5a8fFl2vU1bQpm7sNLysTNgwXaEnVPkLwne9WK/CKS86r+/ZHzt5Q7DI
ZwyHkHDLLo83U4Pw8cTxXWPo3y3uM9U+d+3iqmRYUwApQygnfL4eMIpwjhzkzfWC
XAN8uAgD0mHdJMEOmyZWPEqXtyGfrr4zTvtMGtaNSTgV1U1ToZoyqI3qDCOlPWbn
Aw4WvaLYvt/ngQPpCBAq771tJzdfv0RmbFEvuvlPDrmSFM8rIZ8U81N+3fRKVpja
IyOUnw7815dE41GrKsOI6JtmQZnVp8kbqrjxA54TN8qz81l/ihvU34ffEtfSbiBA
ImAP9p6JhffjRsZ1vwPydxlsb9Nxxb1PAssK7RcElvz82vYi1iSXRWMTTGmHkcPA
VsEo6TVxELgkVqeVl3x+SFfyTJi8B8ALvzMuwoNUGoqM4tGmsjQyQWkOUAK5WUCh
mvlFQ0krqY8IE2POyP9q1AXesMbhMED18KQBq0891dkeVIjQLF7dw5MGK5zEmbwk
7gD++NvJEsycwfn6D1R/rYvyZY8SyqtPSSkjBrG7kAxpWy/bhlYm0UigPcMhwSnd
EDar8PBbhAOXJAmIuHnyaVIQqBhBe8oKM+dYaDynWlm1YDKIhjeqlR5x7/LpYRDM
z8J345hLYJ/TZ2ZHQlBKv04S8V7vN0Jai9U0dyq/s4ymYycoyzqRH5vJ6ip2mbVr
gUs27CATGtt1Pe0GtKEl7IzldbwvBAxg9PTQlpmflyXl7Zx7oeMH26nYgggEFZyG
kCLsDowkZofIRIW+MessoGOdxpNi+BChWPYz3+S4ZvEah/yT8+E+1tKKnjkZq51t
0xiwgzk380Fx0AZWo3pEmua3YVGyqZM3rlDlUKAbqmXW0goCOqKunwNe4KVshfGc
L3oU4WJwDCofBJXG8eeawo5q8GhCS2EXE0V7yhTiku+HWTD16L0XR70HUXTfZRY2
WksiP8G9BtBQPDXpGc+s4FWKgQriCa+c0ByMTIBs9RNdj2wxP68LImQBviup7FPt
wZT447+L88BrOvMeCFkoayb5lnGUVc7f8XZh+T7JG6UAmjXkvlVeYErp6Qzq7rLJ
xHooLNx1jW1kRU6jHbcKiX/JfubLxhF+Abec2xd6FuaKNINjPFBFp7odixTTZ/wX
ZJuh3AC3JTBkuBYpL+QHqZtB/jjKKnhDM3pCSxdPi+49EowakGnssfztCO24HWI7
GD73uX25TL4LgMk0PlZWXuBfVIDesXiFI/2c7qMPZWdQTNRBdt5LkiUCusgfmNyK
RLM36f6loS6DXN8yZDLWy5NJSj9Zkr2GqcG1b8Rv4B12JlcrB6wjb+uhrHK+foV2
MB2cpgG52lkegrVz19kXEqNuVe/gJ3qnUL1IkRtOS4i7duiiXKPCchRRSHp78GVB
XYU1Gb2UuhxALLJnQh+uyiRmUMZCemiDrNc1Xh5tBeb3MJN/3IBYDx48tzacIy9K
3FtWphm77X8y/NlaZS2UwtpqERCWmMJSJSGhXxKZ9GYbdQTCGGCbauT5sDCVdZwE
4Najgc0HoqKEfZ01ZzJ7h8Yp54wP9r4WEZi+sXJARzHvG/tFCST+AxX7Ecb44FYY
qhhiXe1OKdwZKbez7x5K8q2YIVXqGL/9LvZe85eZziUktTEBQZnZ5SAcB/DQ9YcE
aLuddABPeMPJBbHh0OFQ5pq2NepD7CVge/mvLPIhKJow2XahytGMz+ZTBkeTP5m8
iIBTy6IvwI7TMLIbn88ZYmIbSLP2oXLstWqLc9kvZ8KL9408fFVo2er+ivu9mlSS
1YFJvXjelihSzAfnWuTvpKUzxEtpFVdE86CemXE1ON8CjXygzEn9IERAe27D64iO
xxbSbuP+wYcVt1RWcycadlqiyovJ38mlR+Hf2arhzTfZ3TiAEaahMyGEksEXvITH
lejHRnhO3CM4woSNGgODZio3mF4G3IO5a90rFq8f0VfUT2VPsEqSW3DZsYu+PS2U
WaS+CJRa783QYID/88IpcTBkRIGGNHblmZPF6g03XdcfTvIcnf51dSzkrK0N0syb
6gj8j8GlMbJ7xrOrTH0dxR/jrcACmB281FaijOY3KWjSdQSxtxaksAJwYOY3NPbD
7aer9AsGqwmHX54tk4o5rOkLzjJSOBOznoQpUg4bJtkI2lyuTzp/veRqZcR8kDA2
NynVCZeaer1hrEETQ/nJwvGwF1XjkpaZ6WJCUIqVXd6juMWX1WYZdvat7ps4ASXr
GT3AH1Ww5IZMj9YouvhjWX9S/kEyxD/coZ0409nuVbY3DkXGC7FFkPLiCFz7X+3r
qDbNSa4vE7lImyQ+gMvI5RJL5VGRiLGD9zhgS2D6YezkXl9GXYqHHeoFh0c5iS9Z
8+C8c38rFm6JgDXt3XBcdmyy57cKCMxyFylHRtk1cM08WzLy4O8+glH+5reOosAT
/+XfvKMotQrwAY0BdatdsxLF5yNPcSDLnlLtwLQOcwk06KEKnqc44eiW8zyzoBz4
8kRXpvCPf12D9UI7yyX1NGuPh2fN6k5WzSGWX/pvVY4a82zALhaFdddreds4XhBV
phmtHN9sZ3F0AWBq4PH9lbQEJ3pnuFWFxasxL1/Pb9NnwI0OZZEkFFw5Hgm3F4E3
QvqC6z1m3RoAUOaf23mN94PWt+m//u8BR4O3Y6w06CS4Op33f2pldbPjpqS9MJxK
MLk0zM1Gr+sFxTL5uB7by3/DWypS9P5UI2cLvQiEP396WgBGzghFkkNeo+37nPoG
9w/iYYlx3srLpr4X+bPuKVNMT7aI/lHeEU6XlOKtheDozoBIpi5Tg+0wOu+knFLw
+lRsVQIQTN9hX/HnGSAkDih65yMO8znl+aGw3GzYYfS7Q0SANsnyQAGpO2erkB0t
z4lqGP+uSy38YiMDzoJSZKLlglwfLktOw2ftjwGlU5+JoI5rhF4HCjMVFtTbUCdG
ksYB7te5D4Df4u7/pqsAhKhCfOjQsx6mQ4ydvUOlZngv+fBC3/JMDJaJudkB7To6
jDfswdm1Kt8TGTXjPIVoZeHjZ+0HKdET/L4LPRlFf3iQpyYtlXnAWUydHu2dND+K
z0zZHly6EMbgg/Brxpn69eTSH72mAOBJxv3f9wrQbRgqM3tOrDF8zAWZKGfRU6zj
ol8o0zhOy4SRC88DiPWvHY/RnuX23IaqToW8/Nei/VaV2Tftl5nGipxMZOMWBP02
QLphSPDCJl1bI38jPv5CquXG1aBFsG9bhCjK7VYKaSFO81n06oZBI+9PpqzONKhW
OsLTAa7TxdyFb7L0onRS23gXQQUr0Z4kQD8UWTBnwiJMTf5qjZNAiEBS2rfbPPx3
dEzX6x/f8QPR/Z05m12qtp1R9/t2z5F6rpF6jFo+RA07Gi9QM4IlnmwL3n2YpZpJ
Yfyt4l3oEtTzpLYlr/2DCqCZBwoymdOmkrqjntf8I/qN1duvbMZTKStFbC+TeGc9
4iSCpgkPMB0GQ4Xyh/4zOdKgPG62sa3XgV/ztuAXGaQPivjMTgm0nNKl/sDWKdvL
XCVZQ2rdQk8lSpNTNGsrNm86JQKYLjBC4ZqG3nHdc63a99ZUbRas+TuOZWFCbupA
5SFM4PXbW5FCxQ7Pr1Af1AuyLbKtDYxb7lrfv4EVqxdul0F1oCdBJiypS+Py1iSf
dBJml7JoHKur76W+kqB5a9sUKmTRSObVmhdgZzX1DbNqTGq79U0z3OiiHJyROgqE
lu82NRlvw3JbioD7/kFpwgFa+QmPB5yoLkqEtXqpv/h6WleRVRrYbdMwAFBodKxP
YW3wdxnxK7T2SIH8z7xDU2lFuPSsJ5jAtKHzN0GYJBAH084twT7CwA8i9SgOUuTa
cQhHDv0juZlxg/g5wc2bjw57DGd8lnCcPrvl5CE5doqB91qJ5DFkFwEHh7wKl/yW
eVxnLeiVY9lrqchZliI/G3VgX7IZfWHn6pwjcjJrHIFU8/38thFexCm6/o8W9tE/
xWhTQHQlnnYSruoGfKEQGzq9NK6EBSeP/t98cH/PLEuP37ssvvDqAnlKL8Jj6S02
ra//9Ofp6UX+dPd8I/GRaqvkZ7BYNkb9MgNxVnMxg7CRxFFJY+JuM5anVFs1WTc+
+JhCgy+hxfAf7KPyIHFIjdVjv5542uXAsZ8AC/cELEvFtVdpNr1OI08dtE1uYLJi
rG0xO7JsCXvNXjy3ekXJJR+vEmoN4WSoi+3Px2lTBgWM6RaHT5puz7C8YBvTlkns
r8Xc/RtaOTI1YaIvi/PgIdClO6+kFCeu3J2xgW4Y+JOWSavYqalBFX/9eU93XHZh
aQ0l7ZBmFILihKYB3eKfkF/paPQViurvnOc1xYWQlKiq/q1qPFGXC/MEYe39ugdY
4M/B1tcdxHhpvv5EmQqFIpmH+4JKVPLBzR87wXLtLfVJ3rbUgI3tXKipK6eM97we
BPG5Qgef4Od/vEa/JqHUuDUX2oyun+fyqLk3wqDPAfumY/FxKDFlpizYjAYKzYyU
I4olXh2+fLs/N9f+Xv+5G1H0E6i1zbmb4pPYp9qstHMv1HXMatLw8i8l/WL/EJY7
3Fjjdrr4hR6vyJ8qcc1AM1/fYD3wx4nj2Ido3iDMAvGO8NkTUaubGyraiDzROwed
b9B/xTqWAy0ZIKFvzuGZJFAip9HKoOVeUjg3ZhdwaqemFJElc5gidEo6YvbTxM0B
84389WqkHIEl4Cyw+wNfSeayMuSifHq4QUIW4QaIykdumea1SJTDA5EIYFYBBj93
vhNkJYpRPyfZvFGt5jA9tfLCEdwApqzuMHL5mvniVTV7/3qcqwY3+3BDc6No20td
Ne1n+eDBv0f0RsnrH9Iyc7CtZ8kQ0aqk3KnC7JRm3Qclrg8jRGXYQtomLjNMrn/T
PaKMjmYLak89YGz3GSxiD+dKAm1YO3XwrVLTphpmuH0OrhZCLw13Cb7OmSsWu/N/
l+ctSKU1X9+8ejZUsM9SDkv6OPKzMbzy1PKBJNRZt/4m+lBA2/+kiIpcHeCkZJEY
uNzEMnxvfRmJkxDqfPRzAe+zsA6Giw0D4kikqJZwLww/whv1kKePQitNJJ+7793i
JaKRiWe05+6GMRpQ5IsiqAXsAeFcOgShD/ge9wEUWDBQijPRjMq/0vKvwhaIZl3G
tYy+KoPSKYDqvmVQxL3IwcMiJsJ1ZEDdFhRolJSUdlvUbOp3YeJxjhd3x+2HRQbK
2Y6qsVkqIvSZQJLgVYPwFAFUVkxddsQCTO5XnCV+Dpv6x3km1rE6r2ad/esuzx6F
G4wm1oQOSkvr/bOVfd01+P8n5FrSFBqwo7VLc8LAaHLtiaefHs+4AJ/q5mzAlu9X
mqygIYe/JqO0vNpGomMTbwN103cDBR8/I6JLSDzV5d6w74TJVyPQI00jePHSikuu
2Pj4hm/vLgtWyeO5pssyYq4VbnjCDRs8tScwxNNoeyjVnzDtzOxl1JRp1PJATbA9
2zb/htThtTIwgrSwHlqfTwor6/RrV/o9uXlbHtKqzYR9rCB5yIWNG0sAINF95Et4
6rVbbhdNFMRikYak/uEF2f9oYOAZIXMYyRwq68j4vMK6m5rRWf27kYYtDSv2r3r1
DcpjfW3gP0X2WP1D3mJziSl37+PiaCl6az6U9Tfyrl6bIwqDpEb7TbmvBllLyAEM
nfu/q6gOX9T6Hms3eDxpC4Xb1bfyL5rVvH3IMOMUeCJ8jt9WSIHa3/n6xG3hwH6Z
+HhByII1fsYAjsP13UiufMMa+iJ6ixEmbDUAZRxwfUXlki1oGeLmmo9OE9QheCkI
YJwxgqZNHBrJMScvaJ3ECl9HxBombCjtmBtpF5AJQA6sero1aeZP0GuYSZw81rgF
H9vTK+ByoR06GrT5J0suEtbHRZfl60USp9AxXD85EAwDRQWcG1JZs8DPe8fum4zV
U9GIGJqxjXSGQd5gmhh8JO14rh6/n3degp9qh2/JbMsohSEqVENhkCpppeMCnW+t
b57XztIlkHvdP7Q7LxS9yDnSRqjt6TJFlm4zKdR7vpnn4omc5gYc0+klNY9WJOCy
p+SaWeT0UPbvosXG1FQKwLhns//LDCest/R8DZCixtZ4XEKx1VsWfnol/hpaNjaj
Zjb/MXUhdbvPMasGxmrtrBSe+yynCJ6kT+qwUGocIc2vZNZMU3zvvBluyo14SJK7
oTzWmCOrxpynSMkMuhoSJuFo8ckD/+tHmqAr4k166yrkG3V+8NgWw0XE0xZuzd4U
2a4Ocyv2r6uSyg91jmeIW3D89AYjw+a9rl8YD48sJTjlUTGrlF6F+p9V8s3lWIjz
XDaLWT0RSReITopMO/q7lUSviJhomLHfaSTtotVadSIGklmLLYiqVH4wm4rnAExy
zFf5QVjS2g57wNWWIWj+xPF7zGmP6Z1RQniQBNr1gEGYfIobDkW53Wmit/ca9K69
itPAiyFQ3JZNMZZNXzSn0iWoaOdyXHRQMv/8x1aFsIdJQ2dVCZmx9MXRg9/6MbBS
R4mhbWjz9ID6SSOvqJUubEWzit6pxTz9jz+bPWDQI6Mp2/Sp2ouQyLb5vFqMcZI2
fEYYu8tTo14CdVUfidHrlA6ylWqu4bGwBqYZzKN+PKMz7BVWto5TgsjMxtTovs2e
fv/j54kcsQ3ah2ZOf0e+VM7xj5l2eUIdU9B+DJtpPfiKJa064d28uGR9irvBE/Ga
XnxzUzcs0rPiJ5CnLhmKCvROV3NFMCixsLUmiwmJNZUnjox5Z5BQmY24hJvCdTmS
+Oqshyge6urpWLZgwXBoj6yoSuhUzFhdfYRzyPmXm0KbFvYGpLwwAln4QQ/7p6c/
K0flyqyUxlMrDqDln9Mv2/J0QHI+cg2HWEqdDagKr8RSPk0GAqzxQFhD8ZVH6cA9
YCoZqU65778MMbdTXVNo0ti4vDclbvyX524Hq0VyMSX1wfQJpC93i0PiouXM30fI
zcUyEdcgfM2cBP8kLLU/TM+REyb2azqhYu3A9yyW8BgCHBmtqwkWGQWoWJX12qQS
ICVIQcs66IPvhqrIL35SNk2Yb5Y9IZqcWjqhhk/GHBKhPJCzaJLQGZZU0F9LdeuT
BTyv8fWowqf3xxs+b0mipRNTzW+axdTPenlBuvCXRwIBn84tWV2bMLFiLNOS3o4d
BmndLshVPT9fxlpD28jeGDyVQzIJ4NPTVx0efjWxYV81FT0rGuaIo4sufx4sZVl+
KVeMVy4zlvAV9c3Bli100BN14WXqFi+Xd+A0Q67UL63aUnmWfwJx4zMzgcWCQnVC
MSc8DTIPkDKZ2gNBkaW93RvF5oLUqj8B+H/cH/tkxH3qYtFzuPxXuIrrN3k3xESz
Y1WoY1G7Qh72Ir0NYqqCYkU4yhCBXED/mYTGsohF3Q0A1Ku7PsaToaEltNuh9qOt
h5YFO5xPcZZfQ/pxS2Zd9Vo6ZyQqyZJsxwVjjA2CION+NbXu3OubGP3QEPfbO1AT
zqX5erxRW3QDbqMWSgiY2n0FZuwyc0olmPJOyVwxz3pPKR0vmV4kyjkXJjQp7LCF
QTmUgqUZ+EOgXPthFXpro+Dq3ar6fu4eypTdvKeDJNiNmiq+xzGYqgn6FNylpBcy
r8wrqJIo+8A17EgNDQ3aDOBanBs0m1od+Mcon74IEkmX3fOujNKbDF2GLYQvWK/k
WDsOZeSXaS0sTBKHr5sftAhT7vY/YQNlFFYv1uWlZ/2/qPBUgB5i3NtCVPI8RHM+
4mMom+gaooQz3glytnhfGaBMVl2hMgoNrCfnkn9e6BPht2zzRW16WDaYmjLDTnMd
KN3Y79C7L0CAmACZ5Ax39SerdpJkNkuQs3bFfQ5X30KWNa3W5f11gm6SryufwJS/
xR96ZHXcF0eIeZRAfJe38cYKwkdujhWIem9yMEY6Bdnpu+TAkW64yiPoTWwTSa5s
VHTdiKjMjxVjvPHeOeuUeyIO0sPJ0A32Kf+/gsWKfTIwfS1WE4T8xYBXwDA+yZeQ
7g8Wxvy6CWgnN+TtEgcTctgJTT/1pxQlV633Ufwc+NdNBIKollBCm9DEfFiAdcON
3mJxl1rxPx0XXfSSvTtulWO7+hC+OQn3Yvhaj8nhCgzFeVKNYId8gHrZdYZzTLrp
s/XoY2cz7rACY+OgVn2Z9kBoujiJjsUDfxK5E3zoHfBe6l3V9QKlKJlDBZhoK1xQ
6PzWH22kgBem9sQDMHz8K8mw6pdnENYW03QblpvPOOfQq/RND+Ed+lL7BQmkuyHJ
ll02mZOEF2s6fFqvRYffM5/ixLWrh8M66G02KnLLF+DLBWlyPI9ib81gzBTNPmo3
WiMuD6pF68rxVMQ0fORB8r+fjhItYnH8CRE5krr6VEwKmWNFj8Tf7RWcZyrqBCGO
LVYZ/IL0T4kGa7VaVpEf4Ko9tnZ0A65Pd6TeUpitU6eWtowBH8VwZZnRKe9ZLyV/
xdyUOcht7T47dO16Tjy2Mg3HSKt2iEP9Vf8Trx4gOWW+XWW9WO6/8oQAjyXx16Bf
YEcebl5ttHj+lsmrGTGWD1V1XjRJv+zNJo7By7ujmqWlK1rnDFs5UnApp0WdA3HM
E9LyLep2dW0EIMifvon86sQoMJcLLAe0tJz5lVVZ8J3OShtJrwbQ6VIphKdo2aen
ua8r6P860sj7iAFlCIOhmZMvjPAvX80fA/3YtEaLLMTKqsDPa1Ujv3AfCL+4gJn0
ZxzOptLUajFWksW7nQuoJzYJugly0XpbnIKM4+YkS+Evdq2EC+wqA3fZ/EODtMo0
VIdegvzsGPyn8/rXCtVVwmFDJGxb1MJsOfi4UfdQwFbwQE6ZdLQ+7pWHd3gj1GUh
FbyoNSz+AATKJihPOsDZOR0QBNYvPx8ODtSOuoc5aSZCcreTBLIdxkHjMfjtHFVI
LeSUuVYSFOjZ9Mr1RO0oyfDlND//0Tmpv4sBn8OHrBMEhLO8TFhNjXTEOftei84L
8Thp/5QYl+PZoum7lU7u6Jn13aj5uOKdKO09MP68XohsT3SVPzfIeJJIfvWObamu
M9NfnXs75B7XCXLQgMMimpK/JjACZDUkeY1xs7rSwELJhUq8trUG+5FImYvUV6Bl
4zGewU8RQl4udpYWBN8H6AzZOJuUijqlA+d0sQ6e7lB82/6uRtBbSA8TcUOEocht
QVF7+mI/GR+cTdgode4XKPaMOX1gawemxIYYEyrvWRBB6fPuLPdmGS5/JgCirkA9
muyTQH14Q8bQtM8aF76ACpINGb87nmEhR4kOTEb2ZSleffUAnF1R121RufZYx9iX
9VmENm0Uxu6aFbUrvcs6IrFZuIxm8eicze1SOuY8pVFoqNG0UT6NSL1h/IDAP5P+
jmOM7Gs0Oas0VepOZw+EvCHU6Eavrxsza9Ov0P93oG4SAAkMWnquJoyLghDaK+yT
d0IB/+YPRw7vq0Uv5YP6iiL0wFIn/7WVcvLHghcbucD70bgYx5aQ5BPsM0ke4A5I
nGRpJ+wY59gCi5ZvU1DnUNbbL4kDiF8TwOot4OuhtoG0ii+70qtrZcxwuWNmhEPy
Dw9bLmBzwTCKL7zurzmg/KEwTclkhPc6Hc2Zmc2aHyekubSH7+dfoV9eTwU1Dmoi
Ij+nFohSmE7yE1dyHIiEKkWR0EWxLRXEW37vr+bADyuFGd13BPD6WQQD9ScLPKBI
YQbaNjecoEUMWVjjUBmqMRrLilHZeuVkG95HnLigPameCZ8tK/amASO5XlrgaWuM
cIbilbMwHsSqMAF5c23R9dPbxANVpLMsCeTitFRbjsPz7nqj6WwEvqzb4O2sq0sL
4W+ZJ+DwKGfpA0UIjLm/S1BkxMrKwLdcEy353oHEd/eOVC/jesgU7uoyA3xQmSkF
ckXnsw2+fVJKEXAk1+kwq1Z7SMuDYoAy5V3y2/93wmJEq77MBzU8snDAFuUtitWW
Yix3831mtyiemPaJzGQv2R1TtGIlUCChS/O0CthHUZTjngilYd3bHX6evdSyh3qP
xVyoLuTlRRvdtWd3kneRRNo0jNwfzfuLQfYDUlKxPi2h6g6RmTp1dn982ucIo/Ns
TleC+0JzpjmB/IcJxo5CJUkkk+FOO3BbSuhv7wmKFxW6lyfTa0TfpLKgQLsh94qB
LxCGdfxwFc//92g1Laz2SIhRhlgDMXLkcnK01xKMMT1mkDD3CiUkg+q3c5QXlXHd
RJFsW7SCBRaTzDpC/nNvKy6maKJmMHwGE3n66TW0npCeQrAjJJGMmDF2lYQkrpf4
+7N44QyTWylAdbrswHF+kITxD2Qeh1dFGElVcgivbQ0VryEF6I64TtpsGCW+/TPI
alX05VstPG9hDnLQ9QBHa8HE5pMDpB9pBhPxQ1pPnH4U4ZyG2U0I+MQ0GJNIOq5M
fZggRIu5QE3fFHxfu9fVFSQSggsUAh3RIO2gf5wAnC+gleUFtTXwri3MPj1WWUQx
wX9hE7PVWNQjByncrGiz4i+uG2NnHH9Qhf8zk8xej35XPKlNGJTOMbCxZIg20LGw
BhCe9N76t96ySa6oWqjMJfvsAA+2dI1DUSvVwJasNRl0BSoXsWgTJBssqfg1VJ7v
5P10U3gR6l8THpG5TSlVbavMbKZ601QIgJ5sITwBt77xU/vNT86kzGjxPtJbN/vh
kT6x2/xveOPfVHhy/c5h1U9J5toChrQsiDSbsr47ngd3frv6+DilmE8xH1semuhn
nV8jFeqio1ZYAEmw1c7KQEsZmRMUEvZPysNbQVgHJyztsuVhiCyofHk3aZI7nOHd
BpKkbVHeXiFAFDKV9dkH1JAl2lYumnybn1LJMg9RGG1eqIMXn9fpvyB0tspnareu
QlhqY8Sh03b9ftQk2UG+JohbaH/iLVfXFNHKrbaMUVA92s47Sxp6f+pjL3Xt++QX
zeAtC0Fdn9kEg+zQIMJb9MPG1QtRW0X/dnNUSfyGRY0lmc77ZSyu1tgJO3USa0Ne
BX3km8oeYHyCqeQk3vMXALf0N0xcv9dqkFHD3RydJc58vb7i58coHjeEpYa+IIlf
EmSEZKbGdu2ph5UWvms/QDpi8RiqtjBLZiJNwzxDBh01ty6xZSq8xGSOJ3jlNHUj
hekmKKLYXbDOxOlArmLkqrFbMWTjQM265AbewB3U/mRtVLSoN0nfYqTtZup3low/
b+Pp7VPdBkZ+DvbyITHPSA7ufIgWVSEACXV3eL17j1dzqYXh+0jflCfU86z2FOAg
6UszGFD9lxACh+RjSX6/b6rpu9YsyHVd7sm2XrvX26KOiOcSutx2evhdcuwFSTqJ
RNrcDBIUR1OHVsrNkOWDW8LEa6Btly8pGG6CKBm/gsTBoSF/c5EPCx1jJo1E4ZAK
CTeIKJ+a2q82DIpcpUB6Vji44bjsvDAevJjG+2GsN5zf+5Zh2EgDAlh/l296SpgK
z1w7AZTPt5ZMHWIAGK86KD4BscoAUbBXzIqEoUke4PuGlNtovHQcOZd5onJbbqj8
GjyfeJdgCnva5/OaYu8RgN0I78YlwnRcuZGH3HAM6CWoMZ5/y/JTc2edacumCWHY
GasRfovba5XtynGAZE9ShxVss8qCRnldlcJhLJVd2y6goQinwaWFm4NVmeCBlFAq
1wOcJsFssZTWKFHDKFevVZJgI5KxRucwjtouEWwWzQCq1s6BOxf0vrq/uoF4k28n
Ni4kPAYAJyGE893JNuwVWgru3V9eoBZA9m96AUYf1PFYb7nJQIM8YacWPCBveeuk
RaTmVgswqw65NzzIKkB1F1avR0aiq9jICRp/IjVRkCkpnhUXdXrWZgnfUS+eMt61
aLDakAu9p45/DSXBdMLSGS+b713WFfvA4yGUWAvgPLwvAocX49bTdkWQhaFUYx/I
0ka0lg9G2vQk8NVz/usfmr6Afg4RljnsTjG2vEMpzXyfMuhCIcjMQ5forxhbkR9i
VGD8cgF9YjAWNI6MHC3cHJwwELVB2MFh/P9E4nMYo2XhS4SxK8CVeTCK6GUKjlAC
TjTc44/8xakp0WsGor0pCxAL3ClimRf1H5BpWp26nlf//cqae+l+UBONzLVgeIKt
x+lX9FAm/xRlU+ZOG/ZXFLhkpQPFyAZt9Nck9yhFYOBoBqWuGNYLzwaGykcJ3lQ0
OQy1kVQfk7dZlZR5eBs3nhThNPxCc9exBLkgPGxyQpb4qWzTMMsqAH2Tb+/iruAB
oT/kq9BQSNs7KdEH3rll6V6g+7Khln6GFFQC5Hr75AMGQJDjrdjUM+LmtH3FOpde
9b4D2MdGgkKY3OpoceHfM/b+y83ZXDamHq7VxtXPS5xkODAy+XabSHsdu7XMMjT8
sR8FkBrgjn+s6M6ft5A769qH5AfjvF/BkO9GHHeNhOtyXDCPJRO1r3ShHYWS7uca
zOmRZiRvbR/ifrtiT+MSsmQHaxsN5we9GQX7bcQKZLLsWdrradr2vg8azYEYjcGa
ylkclzw08IuXIsu7RNIM2evVNS9kZJ3nGMTkVTF/+/EkgXYCUmnwor0ahgk1aDTp
IuCINfA8sMWnvJUa3bqT6z9y60NJod9qS4QHdxEx7VvWcDOgavxk+9r9YQ5p378b
Vb7KypfIBu5+gplWiljsaJZI6+P6+hFqu/jttdrMzZuAuwncvT0SYB0qo/0I9XNw
pkDpJFqmnkqUDZTHU3uTq8bbhNTpmy9GFtm2k7Ggs7XlMIzeRv+7PtRh8NXkRf/E
cMqlijGixkIwJU2XvS3wdU6MsecJtvWzXKmSQJ2X9F2yk9UtjhduCcLZWMXhdmsl
5YValO48KMP2qKSMCJQLw61/eAZaNDdWfbmCtYfbimp7Bg+wOzC4P2FhkE92CHEy
AXn76DHaL89U3JsSFRivMwT7vJMsOfQIB9pASvsA6Gv7VbAi+mZu8Xjm4EX0tVAl
fIM3pN0aKPQdwQlXCbd3qTQg9H9yll9IAu6gnq11k9iYv/ji1tmqHOjc4s19EqQL
F/pASgf8oRoit/Brt1+uZvPoZ3xm+MnkRifoccFFn+xkbHiU+MwG+u5PaoMYflxo
3gqppXVlVSC0vwcF+QnI8uVKQVKTOPBZ45EgROGaxoi7+PyabJnWOyi4wVidzmnc
znJCsm5R1C7xzuVlQAlFpozMCJY8mbtHmwRtQDWYGMGKgS+giA9GqYgBE54BM3y/
JfNdPU67abbLpfyZbhwSDspwOWlyz5IrztLftsz7T1RCrAUx/rP0QFB6kxmPlfZ1
ByNVRK5gvwYqCVAUtFZ/8Xc1X1qRTCtgJ1iBBRgeQymOJtgZua7BQhenYXkgDwbp
6LRmPNFrM19hpdqFdvbSsZCD3G0/Mai3IUY+gk0DYOIFfgKbz4OvNyUW9oSSVssC
kI5qeft9hDTdwdHFPrv1gHWEVHbV5VxTaLndz4Qiy0iyGIVB6gy9nlpdaU7+SZ5g
f9mALwXwQRzC7uYLgChgPKefEEzXF/EcddmWAgb2a/D9ufBXqi3jv2huQ5i0FtSc
M5Xt6aElQTrBdlDfcNpTKmwcOkkdb6J5YYyeSmHV4r63h9iUidjPJlbXa+QVOSLu
VkY69KAGvpRlXH20xFunmZabyZICKI5LkWNk8YMJ2igWvxMwQKlDQPO2Y9e3+EtP
7JhQChL1gmDatPYgtuJe2iHC2hzXWhHm67QaijVKCrWZU+iT+IhXDtWjYhoqNhdh
yJs+eaHdYno0utMUUpuDmcBX2Oz7Z3od48h1oRWUBuLPi0hWfSEX8F9Ki0CR1w5h
8gSFz8AuAe8sx3dRkihQnt25fffLQRKw3rP5yFknJsd++2E8Lg8DUN5kwvXxnzD8
aKxTqJ3tMVLG5Zbk5AMUfmzOLto8z+kCOtEYWWBtTn/3x6Gy+gwCm3afXsaSHpNB
tLQ+CkFG6wBb4oZzfPztL9OqKHC4bIN6EQx3+cZGpDRN1hxNd6wuWEXwgq5wXwTS
S5CxyM8avSAncSZVxHo9gRnw2equ6ugEmQ4FDUXq0kqy5aHUK8hYoSKQWcCRkq2l
breFLqQ1/yuKf1oCj8chH9LdYXYix1eL5omdtYLZ4Y+HpK8a2VahBKXPg8nt+kb+
2aOW+8mLEhoSNmtKehNVjiEKLAZFtnpUdSwCTrcl/eTWOoB/iKkMwoW7Mt7zArn8
ssYNvfRCw+RAKpDCrPQ9Ar8ymowet9MkWVSOqGJR/BnS4BLOqBfAfEsCkuUN8hqL
1KxCjpR+N78AbUqKFtNqgyH24JggZmK7EGHnDc4KIyQr7jzuyVNnte0syhJE4vcu
hG5jc/3vXaI7Wer3tzClHTjsZ8EXaA1WhgcbmPVd++7iGkYy2WtCaUfvXNOGscUu
/I/bcs8Pia73UzUIA9++hot3vkmQ6cpnvsirXVsfW3ItKB+aWczEsWMNbTkj8+vC
+OA/airBXEsOXpbO98n5dSTnq2nm0SsSpWgG1EdfIkdb4zDQ7SxKYEL/6m6Zgf1Q
xG1tvspdywOS9nqUv5wvqxTft5NKwq6DQcImHDjaWJo5e1afHeMxaR59FR1Kej3c
cLjsEJslVSkeTFaz1nDLEXqBvufRxdasWrIRkwx0Um779DKk9/e3KmaQr0KTaI68
nsB/30H8GobJ/9kJ+e5KQVLZESRHzxTH7sIt3sDy6gU5PRtL3h7qjs3ifyknOuTJ
nuqVf4QvKtfRARHhPfoEmSqeiSAVJjrhurS32EjtYrqr0cK2KZKvYUI1FAwXeySI
x9d8jpxkYJahqOrVOKKRlCiJQTJQV2exgZvhp5eHmjeLb6+excCPnW1XUqQK3I7c
zHJlrAk8anMb8ec6pS+5FLnnLuWfLwyQL0qEF9ijBFgCb+y68IkGaD+AvFC7wdRm
G0mvx9mvAalqqUNY/QXzYsq25adVj50hebv866FLbm+LR7ajzExx9OpvzkkiyEwI
Rh160dCZLZn3Vj+SJoK7HeVeYoOIXH4wMdZC8Y+asQHrfOf15yotDlv8nkcikgjK
WOFK0ib1Pz+nmc0TLyPfIurqP/i4Bo8nKHD5MQEEGy1TDcFnq9H/0f7PCJc4jCs5
3mM3aF+fMFDLGprIXAUlxnZPVfGIVV9Od7JfRNfzxYcgdcE2Yh5cKOkRDPRZhKeQ
chLEKOq1BWCVhe0jSP9C7TyqDH9O/Z0ALUQAnxhEcE6nORk3dpUJVs0u86ivtelk
9PSftw/1ekpwAhSgDttiDqAiQcfxq7DSZOFQIsvgjj58s+3GYR6UnVx0LSo7tArL
+NIAxlD5vZPYCbjFBuiW9ba6KQFuo+jKP2ndv2V0p4TlzcV2CXngnkZ2qbSVON75
kXhzuZKznNg9WNg6UrnZhFIuFLCc+OU+hyrm9h6nWeEvaLykbEUFwmoI/MX9OAdO
xptfqZo4CnSRUqI8Rw8FDQV1rxGkn8RBuYg3eUGDPxHYW9QU6/eirSzdp9/0d/pG
E7JaK+4cNSJEuQvH8cKTKmLKvCECkfMnWX+j8VOcfv+Rmunc1WTAP/QhSRke3ntn
0QXyofywv+pZY/vrzYd5nVwIt2B9Uvq6F8HBkLrD4SVMYz95ok+zf4kkyPGuwndc
OnJ0P2c0waI/YiZ4X7tG+IdNqpYjgpzbU4Oz7CdS80LBfKH9k4IFp7JH+jmvmEfW
XUfqZaIxgeIHRE2NQTtcBdEI1tuTOIxUMnyrHbSRXyfcRfRWLTvj/w0o5PIJ6qug
OYaIzCuJzQIqJGlmrxSIYML5sSPRz6+gQe0DS7Pkk0HW2Qxwx4svT7mYY7pAcn05
yS21hKHaMUS5DyNJlr9dXMvdPfMCFVcdoZMbIGzkZntlvuAbHazQ4KDu6CVuQ0GS
CSRXEOT8ohg7v6k4tsjkyxjCn5MDaMRcnVX0MzAuE5Wnm6CM5MQqB0JAvXVrRfVC
ZMj5Lw4mIhoPjO+L4+CgU5xuz0xhdMYtZGNvkV5GNYsIFfNtQUEaWVBwoFOi2xJW
MNpY5ZcypCUIZrY1vcIXE2kOSc7o8AWQRoGIPsw9+3bYoOoN/nsoiFy+/Pwu3K4J
iIumeYTYW+HD7SKz5mJN4Hb3Kk2KxODjnwgaYdcobKlPeP4gfJDwxTwT8vFesF9E
6ovWF2aoNMssdJqG6c5xuw5vp6/3Dt+7Uo75G1lUtGMggsrZvhX5ZQmC5V/1AkMM
6o1ILLmxx8cQEJF3bpJbKjIN2Q3bpTdifBJL7GuNmhr4/3NKHWWeurYbdVVidfGl
1VpzSYyeSsbhA1WXYI/Cdhx+k0SrbXmmDswBR3r7cjvAJ+wXs+miWCwLUL4x6adt
q1ltLeeMEEVbGcwvjFe7nixJ4ETWMXowP1BPTuAk8s7+qsuN2v3uhC+qKAO5lq0o
tWGLGUtGPWgdaHo6uNQ/jVtv3CR57HsBt2h3OQ6Y91B+Y7dtLP0ZE67QNhMczIaQ
l/p6cl3vM3wJUGJMZEFRLUqaRKSt14t3a57knaKh/XikefTpW8rdctTeKyKGnOr1
75hHBhq1q01/JugeUWaQHZ32ab+dVd3zrjCPIQUFL7tROW+rsG9v2cV953K14LcL
ufElp53pRWVwllrJW9FiwUDM8QQ8MVYlWop+u2h6u6yvAu0hbixCWk5DdRATyiap
FUrI3sEbGNC6c5aCHD7f1O/pR9S5ZPICOfUaIAazKAybsiD/h4I0WciFPmZ0aajh
XV20+99t22vp4x8TxKX7zk8vH0Y1kThlXkaPfKB+hSNWlAG0ZA4faxMGDHCAGSZs
G8gTCNbIClNSUWroFy0veMu4Z2NziK6NaityxH2E2H8cKxq7FDtMFnYLgIHujtZx
3jStBUyxrjgUGdThbdeqZK4Hh0Rvz1dhmyamZlhIPrRUjSGhrjNhGXPc8RfvoUxb
m2U+B6tE1bymEvTZY9TiB1fewoFru2/twLFBqhoUjoNSKTUHCy1j1B4JS0XuNSTE
UGeENv7RLL6ZaAsfqIt/6DVUBog5w8lJsR7J2dKr+qQyos3Ohwc685N0olCo+NI1
35m361jZ3UBICmG2T9OK7b9fQV+GY6W8D3F+h7yUuojxCoP6HwHQnTKkGW21vwPU
BrIUEsTcUrMGjsUuxT+pJPbuqtrUeyn3lcLRSwZ1Cn59moHEG2Qpa/Jy7XmWtajc
GKRFjcHvhq1S2qS9IFFYkhSNgHcK80BRqQoNV3+MpQEpibH+s7mJrzjTu05qx2mW
HPYxpP61G52Y0jf0F1GH0XWb0ZCs/ZEJPk+/aSOi7/1ZU2PVObO4s07J/KHT4LSs
MpZCzheW7sKNe38JhtGOBNUIELemVgZLCFC+YyVu53/gJBp3Cvae0p0dV5sM9aLn
Fngr9CPIMw5+xI7OVm6Vy82HTxwtZRe3CpLFIS98lHSRWDP+qqqkrhqki0p+0u/W
mR4f5Zdb5nxuZZe8YHszYbA3lHsbYODDqtcrp7CL/ehb+pNNIDkmd8cOatClAncj
wK9Mrpq8vd75Zx1WADd7yazFEpnLj1D4/XE+xOpWQCSPskBlu8+xN8mDnyYm+EnD
F3qfnTs2B5CW6HbS3YlPkb2xUMwvYosMAM9ZAHfFrWWdwP7AcLr6uIWkR/oLlFWT
0fqfXw3lQVENvlALiO/LyRTaygmDpCN/lSP/DVbwER7mI13IM63YYUmH95OYIlNm
cfKhJ4/1vq/yUVG0I0BhZdjdyWWKFspzjFZD56GB2VwebkaKG5utc4qvQtlKNoUW
p7mpjUfY2FqmjBV1KoyB5KLZh+ZgNvDZOGEG9gXUGVT1nu1AbuEiofj9semwZy4S
ASln7SuCrpSxIJHJlC/bUlINlvDcHk6Xa1+7zd/C77dkgC/y6w5d9ZJVNGDJ29+X
ymZbZ/SQgv2YswrzpGhUEB+bijBolIwJExtGjPy97TpTOtPxLRErDrYpzvXGa4Bi
wgbAav0bvnv4x52Tb4KH6fjQyTHwNXe156KTl8cumegKGP5j1a970BUqP8TmE45K
k6mOyfbRMKoDn20Q55MrcuqfPlZEkHuCoov+Xx2KT0yaPPOlvsaS6jOuYmsD5h9o
6x1/jyZh9/9i/Hh5XbD2TlFXl7aJ6pWCwtcNyCol3HZXyA+msdDc5zne4CduXEUT
K8Eel93axpl48nPvHMLgK6tel3Vl6ptsbiHrKI8RpCXGSVeFf69gnjFGCO5yYMKb
8xPffcPP0f7ELg8Cu5xb+o0fKwLM28fIv+tRr9wJ9jc/63GmrpDx96tHRXQWzwfw
ybuxnRIlZ8+Cu0ERFBTVquFq2pcTDy98qP7LwJZVbGLVF6KOIMlPGzVd+HwVvjZX
4eVzX/qyLlHnZXxeynwElxv+SvoWe46Ds5tytTC6sPwVWW5hjokqtZdtnLKYBefv
SbB0qKspk1CXC/yrXDLarnU8AISb6VTG/wZFcR/CBJ0eJfsDSYug0y6Gsf4k4YfL
TKfj2J/nt2lwKO3pNLpAYCnZ+4DZBviFIekLiBFaIdBtvhnEdQ1yLQJi9AJROw6n
7YL9ZGmJVNW/iIt+GkMGkmTLYcBZr3RrEa5SY88imD1kxYtYEKhOHeMhruCG0zZo
K47Nfv/dAndFKuieQDGwIv4E3doyk00q9fiDIbjPLDX5KgL8CJMJsn+4TB2hVJEI
nvjBlF6+yBw7NWE6DUKpw/SRNbXzggmYDny0kOPsvo92ZJ5NqXj1ljw0+jaAeIjz
LL9bGyxpXTx15yGhspH9PR/iGS0t4QLxSPdFbMlVDc2hP0nnsEatiarwlQ2wiOKy
wi6sfAyMZKkUKOPIosK2wfNIxfJFXe3rciVbcSnvelKkI+pQVFhbTdbLeQUQWALM
Z5jDP9georGM+iC+TWSoC0SbkEdhSg7e9s+ZN+NZO9dvJmSakoREtmmbTsWoMtkq
AR0iPRg6+B2Ndkjdxxf45QnT9Tox4bL1IAQFu/a7njfSfAiu9kTvOHYo94VoEgwL
Ww9ewa/EAiQX5d4cm6lCEQTbcDhz7oXp6KKz4noOB8oOcm0Gskca/b8Kw4Q2Ot0V
Mob9QfOJWBfBUMpp4tcAce2KzGVxmenrXlWIwv2iseiT5s2lmuWQ6Um8oI/BLNlO
KrpQApRfWxVHpPXuIjx5p5WCLyTXcaF2MhunysPHWiRV8exl8qniZNMQCauSYHPf
4xlFC+TAo31M3YlD6YQuuW/04jJ4AG45W+AEFxO+sGSlSJvVonIMWlaA7mhuvH6m
03Ro3hca9f8+5H7MYWcmj1bjH8T7AxnL5DNqtp3/p2YKJguaFsb01scV90wI/drr
P+iGNF8n4FgIesgbFrW6lmL5XEuidyBgoL23P2ufxjfMzWv7a9c4tg2RZftqW/Vw
DLYfAaP4tmM18Ux31bz0gpJr7rOujSu5RBif5IWMFqGqSPJlWlagznRG7PfPAI5U
6gy+gb2RcImnqHdRbzNtGlOiYNWFKKIaQtJq79ivYDik7jRf5oSFWdjvp3pwmqqB
LIOeyrkdaMiurf1HQK+oW+XSoIXZ5UiHGJ5G7SR/gr1xMzXLjl0px6+HIucwTAPZ
NIE1uYBQ4Aic5ULSMrFz3ZdjZxBNkREkDcy5DNs8vut5Aaw44/g6BIsNpGAQ9Ck+
RarBF0h7FYc1gE1KntbgNcHQWIieMbBYYEUFMoVkwj1Ib7sapDOvL1r85PqB06nr
n41eN6uHd4ZJGiYTv1cXdiywIOt0YGy503UWUycOnF+U3VRg+XttMXeaLrOB4U3l
WfqqBdtUW8gnBXh/8Y/wy/+VhSmajt3j/0cRFYa7yMEDU+uH6tubF98sbiS4fTHN
CFKCWJzKZjzvtXRtr3Yu0lssp/1phzdRk5zZyzFz22sXBDAhBIxyZ6wdAfM7jKpO
nzMtFT2D9wMZ0lmkcpd1xtlMWPvZ0z+3h4g7YViFQW6hsrwiVFboNbqwcVUcvMkD
twoB/v6WijpjM3AlLXO76NGoBs0fCoL+A6OVPUTrJW66xJHM0c5dBAS5pBaT6HCX
EqUpYUkSziSDMjbvvEckvehbMB3ErK/e5nggnOqsQPNAZBlu+kjg4CakGG8hmfHA
3ABlQ532bM+Kn4zXng1ZyMGgGCfL5wwOqlYzctSJoX6byEYXAihXvG+1MuU+vUQh
jL9u576puqTrrBC2UG9mMplh1nwXZ3SD9N9DEJt769cFsTrcmSEP1HElqIszLJad
yZn1UiMOEXbMxYHfuYMvzBYrdn0i6mEOjJy+I/FG7Z96o2VNHLGZ1CPsFF88Hay/
xNk55qbzaA6WVtvrxY4oWRRDB9w4sZAtS3a8XUoIbRhYGM+vEeftpaO/B88MBRUF
s8EOIhHtYtfn1iKeaeSDe1suGs+IxsCf1zxmDGVAWAQicRuDEztV8HNCuvqwCpy7
Pr0GzAUFxFaRHP2jRhWZ6bTAfMCRrTku4O76iMx4Qwn+CrlJvl5hmWcsslQQVec6
oeDxoN0ubZHq8qWfYqqxQ+a05TmecBP1QBb0XkkPPVdNYcGRReJlYtBDDIFIczvj
FuR9Q+quarPSY8lJbMgn/TbuxREdSJ8k4BPA0TvL2udnMKI9nxrhrAmMvjNWcbX2
RBfktSX0JAn7xcfsbpIo6C9ihrOC9fbOkJ9rqTK6Eq5yjbKGpgjNdTQ2fPxFpDQA
A9XeRZpJ7no+WsGJaPTf5sLHy5Bt7ZOjXFeqN0gBWLzX3NowPiX2z7n+fkH2J9LJ
9ggmnEtFBdeURLF6ac3FJMrrUAWrZyI8T6piODW9ORMIGs/C38lF3g86Zzxycbwd
AjztQQfkQwQbxAFMgOAX/CnURRA0ibnZPuvsIBPt+s9hDl66MzkVpQhUlnn8ZdqX
e5YGbO174QF8ZTstYxi9nC+DTxUoAH50VDU6Ch62071k50qLNdLzIyRUaQn0pecO
+/mCm14aZjI0kVs0SlSLg/S6wJXG/hwoI5aHnBEr1PTztARhcZ0nRBPFXabWhgQn
NNcGrje2KcM76iWXGgaCStDDTJ2zOoxVHkkkph1uskX1U6spMKnL0aSDSrm5YjaD
bAYXJz3dk8mpE5KccP8KDv60/USJ+2BzgVeudItqJPSquqVPj6JD4hd3zK7UQ4Zl
ZU9EI728blZsaXyOtilKyyRk/UAt/xZOh92XrpBoAvTlGRyCAeH+Pr/XaCZfnIf3
QrmlbtMUpR6hVDAJMCsK4cQj2skjytZxf7hDsM5Bqq+abPuDhtHlJyLqP5eyTirO
YoYPAq6/SfwRDbw2CqOqvuuyR+ZeG+QMuPRkQtTKac4GF2kefIQMOrGA6NfGbfGV
5xvCLsl21QkdGy4/DYItOzDy+8DZMlT/DKaqGtZjW9PtvBjxE9Gek+L5AKQ35QaX
LINzidK6UDaM/p7/xJgtU7t6mG6L4jZlepU0ZJ+l8MUghO4StJhfZfCEoisKDRlZ
4WegfSgEY4TkpGEIJGyYirCNLDmZnxPD8C+Hml6RaN91lZIFiidIFqvAfea9dmzu
0oL67FC/Q4FkEJEcm3PSB6HQcJN6eXEypnVb5BA2vDWT2C9jROYMDsLfSdfc2h68
mHnWSN/CuWDqgE/sGaKyXf+PhfW+t/seFmlNz9NzIfzCRrJms/NOzfFWfz5chMoB
ZI1JBHEVNfLFBJBEDZ8YC7AYe544aev+Pzk+YgyWGmPKRB6H/l7a6F/sbaHT2qBY
moFcoMBUnmPglw8BSeeXEkshR7NETXQvZgYtBiLwTdrv+ydZdyzmycrE5X/rxVdG
pgVP142sMfXn1imqsB/VgMs1HQcus/hKyg67d63c6L9/HF1Ql3J+a9ZKZZpyIqST
ISa3XaDKTdb9Gge3qbtYtfOj3spEdIFfgvUyoUjP62t4FB52xBr76Do5MzzBjW7R
gQIObWLUU9iZjQXyKgUoQgvrXiVRHOxTRZxg9yqqxgZ/HR9W022dqZcegCXEcilm
sPFz1ev3LInVIaMw7CpfGQHAv/QMapEpijTBuxlSQtZHbALpq/Y7zPXWKRG7ncj4
JFRc8eGLOjoy+E0V1nVyM6kIIdEIkUzvdJmmczs4htodQnosMjKUjCJhUbIGgAJR
SWLfCwjdnlhf3CjfgxF9k3msHEphFJLmMZMZk7rRqqhX4adGIrxjrGrHo3K16zFG
kW09W8aIdw8qAUEuFn2Okn5lQWayX1zwdf6NXPwNczpI1aT4ra7Y1NfARXSP8QOb
6gnLmFS+vgmLO3YOc4ORd+i9GkXIfn+9yxoWmNLTl9ALxwoT3b3Ddg+4FwzAitxq
ROpj4jU1bRcEYDpRIWZBemGTnuE7LOGgkMO7iZxYOfmLLSX1dMmZVsz4ZHiSlODn
8uDT/UpL3Nc5Dqv3YBNxEZybzpD0vGTxsNHtIlrb+TdQ9hJThDnDGRKXgomeyaLu
y2W99q1QlrZbJ8nKRckRlvU+1l1ipIsA2q3+idVkrhASMIQFaW3SIgsJ4EzUdY57
l1pp82YeQFfoGpVe4sg3gT3MQ0BoevjotJncMllq2vXKJHktpPzHmp0lCjmvY1X/
DETXWPwZ1WSwuKyn+OvgA8RrvJqJFx68YzTzRS5J0pAh/gWyodyYJttNGpXyEZOM
6AYMeIW+cn2Gwe77P5rGJMIYO0FUTqo3My9E+aH3A+AGetWE/LUVHsPzDAuVn5j1
ruGNK8uGwmHeb3Sag4/oyva7k5xbqQoECAY+ImBubm5Nv/JulA3vu5VIPL97gvsi
haCFTvyz5hdGZKH0VYUImFMVd1tB3jalnK5hdVnyNd+BlqhOyUWkVgjk95E444xT
jzzOFYuSoHJHhQlmeF8OQJrT6s0SHeKp2GKO/Cgs392F3MYA0J7MMTj1ichpB4gs
nzg3IV7BctC72QPXFx1RLCngtQJn1nWivCJuDhTWzuqWmSj5p/A9XsCXKxpk34nO
UkNV4TNRCcfX4IeUjnE7PIAief7yVNIVoRA1vxeRN71jrRFMOacnA+BzOjPAzJGG
m7BPVWm/qu5CWGRb/XD1ncgqhHYHynfA8YMYIV8GxOs312sROBSAhnOOYGud6ttB
/w8Znpry5Cx1R2CinCmbkYvtKOU4hszlxoI/fegLQqUuTBbCUnDuOYgHkIPj9wYU
fCOpkuPWLAc+1iEyN8uWd/hJFgFxhhzGjge6SMIudfoWA68DAXJw99ntiFY8Kz1j
HFxpHw0O4a92fOCZppzKYeSMxEGuFjJGHpE/tGQUI+9v3rN/U4TIZQ+kR8RKrdzh
BakpD5/hpgH0wZmoWrsZh7ChQF0KQLGZza/5jNuO07cM5C0MibBQUxjOv9f5c/KZ
3hzTSsZV2YMsRLjZzx2QZ0JIiXojJgPIXiNG6X+vSllWPnLE5hzAUXSSUTSC1Vuw
t2oGGJCwU+g2Izf0WNNZRLf39JsU6pg25F0YtRrvy8hig+RL0vbrYQihuyo/jvZY
ehq5bjb20sfbzWo7VAgYE3Bpf8jxwQnqrikOUPG/1+bE2dFo69l9OXXDlyaQnG9A
6HU+mi+ZohDQnZ/hu9S94Uo6BFQ4f3iEFlXYxS1UrWhY0ZR5X8o3lvuCp94PTLZI
+xf2Sy1chQuQJipTdMbhVaal6FyJAMo8ZaqSOHow9/CCqbxdqOWmCj9gW9Xtnq9W
TAxPuTKetwK6pu4bbEpmRMRriVELzmsz7P6gAharJoCAGz3TjcdkYQQusuVxkSVn
jgtTL9wURQCHjbljZI2TtzUdz4qlrbC4AqkuPHln2jFM3l+Znba0FY+BQicX88ie
jjRm7vFzzS7VP0kdOysULvFkPdqSrgQQ5ZHqNn1wMLN+f+hTwC7ssHRhNSAe1tyU
cv+/EBZ2btRjlYo+8YGsElqqXMscKQylydeGDsklEJ5TANOlyiw8PjXS7WN47J6/
+gVoMumfR1KEfwUCIIBtjduwtKhckIGh1M/XkfOWOzx93DAl1gPMaT74zTTEKMG4
5EaC6rCKks7sx2ZjtdipMVTprqr6NLVYCSSi2Z3HrU19nlUQ1cWR5z4eu2m3CgTi
fAdx6Oix3HrVSfMYByqoZDDXTMlAx52GuU5II+EM6sW8IG5hz/lYouEmff/NGCl+
Po5nkyItZB379YKCS1iVPpw+fPglYqFUCTbDjR5vUrN1c6TRTzjudgkfA682Q41L
L2M43rszHBPsvgwm78HjFWY6tpE3sczbNhv2qAMrGmF4EqH72UmCfqDcpTKAXBND
cgJyACdYeJmPK31WFTsKZFkiUWiWq4Jvx/23uDeB+yF2uwCdDSFiAhii2fOsDpi1
VLm/6V309iJGpcodaFu5bUtK4WzpNLNjRp/5dcxAPhhh9K92fTGGg3J7QRp9RBlb
D40/sWhKil/Iz8duIqtZ4wldX+nkK13tAS6+lIWj57BDjbxEPluioUCXBorN18nu
oZr2ytwDYJtJeYmyV8A8/LIIEa5RdANZpwJ+HPd69W5g5qvHfs00p0uBG9MfDPDM
5C3E+rCyFQC/Gt9UJIJy+mc/bmwBGWo9hL2jgbQdHfDUMbwzdhXOEK55YMr53PI4
oX+Ub1eUMq9f1OpDKUdo/UKNTeuX7ZG4BLX4f6RvU/PMOBnuJxY0V2lgUJGG4Zce
N4FHRlwO8B4g/asI8L+5CzuECnurfIdATRd3EXnzr4nFttgnjkGpipzIfhR+keV1
6Fi5j3DGDwQHdnVPIE30wco0ogaI/R4xgQxImtVgH70vWNmo8LPMZu+6C1A71NwZ
xmwYHcJ9Ult2cjK61IrrwFqEvJWLKyvqn+1hJULgCVrN8koXYTlfRBGSjUWBWbQU
yQk6xN6ysG90KC0Vt8ZJulUyRnuhRyZWC4oEbrs2zKUe5BJFh7CLl77tNuoDLxPB
htUGuvn1bFAX9hLF0Jjhazmdiy43S6axks6eiU0oiDFqlZrGinm+YRVIALhTbATW
GPv73XVIwkSfO25p8n9BCwg6QjQ9sZuviy9GYr6jSKE8Qb37lahVp030cKunhuiL
NctusDbl/XZYa36dFkZPgRCW/mAYXs2Jm+YVNq+HRcguCb75gEecpiKtj/OdAPhx
4r26IkX/yi6ebPJXhFeZY7dyjgGudSHIr7FUySwodluvpFjovdUSAhLzo7yPPvQ7
aPmSIlZkzCx5UcOptd9lk+Q1RAiMgiHscT3nJ86ErknjrsGhSBxDbOwum5k68+45
u1tU6tOmwzONlJ15uhCMI3p5iLgdMv8fQ25pWN3anRhLG8oneJELZ51P/cn6JJbX
ZnCO36n0Rk1r3+J9E1Sk7kkD3MDqgCTJIeK9Cr3SM9D9oI25bvC2c1c7oPulZ2Fb
qxqFXR+XZa/TB472D7p5Fxb9VitDMNHGOa+YQ3qsj9JUVZTJgNjyUZcvADkmlvfm
1tVAyaizULgX2eaP+kcMIEbnGjvqfi2Ky5LmDss69yAi+apeGcei+KNF2qFd+SZY
jOnIYBGoomivTCddLOQ+/OOB5Xbe2g14h1sQAkdxjtG5kcXee8zHbzrbp6wuPxI4
rPU5GWalf8bLKOpatb0bsf6oOR4adRZfpfvLWmoLzxj61Vnbjg4wkxAFEMW3Buha
madYM9fssQrflt8gSwKPsAOaLuDCuySoTW6fg/dLQqgY4sZ8RjDf1wf9CgP5ngit
ecHLodaXkphxIRwBHM5oVnc+RPOuFpgNoL8nW6phiY9iF9yJnEGa4JtlQcO22Pqk
2PofC0nMk0+rmEBJBGjcJ2kShq/SCypZ8XCLIDjWs1xrUfyw3KhgexTqGw6kgkF+
a5a657IhWenMNq91r+6RqgGfIAJDo32t01KcC3W+w2g5IqgKrvxLCnbeGn2pJlVI
uuuoOHBWUy7DeGZgr704/1ShLLDKDespot1gS4OlTEjPihWNYDk8DajaT3R62979
sr0aKn2UjkWhn79LYG4d3hI4cmborv510V7UlLLk00xKr0EGZESnHeP1Fnt5vtUc
NNK4Hhv6rdfY+5SfOkiN44pUlOs2QXKumhu4jXMXBoAeIOczW72gq8zr7evse3tm
hKijfH7i2y/x/WPw+rvGBk3Z0tKkFzIal0nOf60GcCM8iGrDk7J/2a6I2Dzd8u4Y
1LtZPMdx9FViw77WDeiF4nCeHtEt+WEt7HcuHqd6WDquNQiODrtTopUzksWV0pc2
FDTFJDxYLIv/ASBoHBJzBJE6/39+YUWv7NgAllTvGXKlM3CId0JlabocrljQtPsS
RfjBED7hwSjwtpCYpCoHY0h0c37m3/FpBtXZWimsmCTwJ11iH6g2rYBUfsNuQG4f
waLR4c2QKNkxg8weHmFFgr5ow0BuSGiA0r3BiAgUbiL3FVujKUnz6ow7dpm8pnpR
0oN4ENv+Yw6F9oRx0tPKqH6Gki+w9y5n0UWIamuUt0xkXo+KBzhX3cKb0/T4DoCt
7S640iQiW8MhuFZ7zSoF+2rndaXBSVPDIzeXHyRgZDf/H5ET8TBMWVckLjaX3kOh
uwoIDWOaoRsoizjTMlhsrEijjky3+zK4qjWZTwRZwkZQJkrl3fYdcyRa0Beecg3l
kHHYE0M5B1tO6UYerln/atwMGir2QvhHI0enRs9Y3aJGbtUADU+E+gABvimIt7fi
6/ruro2Jdzl60qCqt7PR8OyCRNpgyEms9A0h16ZZvJcM+wOZvS8vTUeDVLkqYx+f
YuofJ3SQ+11VYzqTI+FaRxryI8keCL7khufz7rr00gKJ6+BJ7nh81IQZB2CrUNkK
+hiVWylf2X3aBwFHYQtNz6QrY6eQKeY91BarqW/FhMk8Hmp+f55YnNbH21wz4l2m
WDO420T7+BnE0Ekbdd5XSE98aAO6ObMNa2kOHlU8YemZhjMgOTP3BBcDOmRc/+Ke
8tA9c4oqvT/0UQMr6KUz2t34y0NYMGS95v1krKLeu9i6bwJqnNOZgPEz0qnQ5t7B
Ps1VmGpDyK35pYDhXZYPnTnCICL/iZNhwtxyEIQihHgg2nt7cKn/3WjxE1J/CAsW
zzVu8Susc3VbYxbQ/KFVmW7AtKJ/ONORRgVNqICInaL75U5s0ItTXm6q914OeTsf
rjAFPDjLhS+CaWDNScq9IFAChl4TEQ32p337goBPWaYeI7SC54+I9VyU9lOmbmJU
zbjNlj8VsqweHqNveISfDSWXBtI2oeEbgykYyXlDFcu8WpHGRUhAvWVad1C5jtS4
3mvOju9R1HPTYkht3jpKklBsa/JdwkZkbg4pKksXq9vz4Z+rH4dXCu4GDm78b5+S
IRbOgqCOTcxWrNareK89DFL0SoKE627ucY71eyjctdTIb2nC3E6Yr7FF1Jaq7nUi
p+OYwdY2fex8QuxD1jcWUScMDhByWZ3TZFbKh5VECcg8l4wTh7Cg8ZTOpOUM/GfR
bKFn8aM9m91fxb0S9Jdx+7F5PR/utAhk3BjeuNe5fEOb0HhaxPvZ94EjxU5LU58H
flHW+scx7Zbw7EMC2VJr6QtVmYl++ZpheYLhHs6i8jsyAqJURU/OohwO6fUd/fZB
IsJags2u14EHAAsaFVXSBuTO7F/ng/XZTyzCzDybyu8PUjjnwNdjmisICj5YtQf6
q7nnD1t770DQ7GozRm+4KauYH3JeAPNwf7O/kgNtJDNnPfjAlHwhZr1/CnIr27Z0
RZi7Wk3RBQVbIDFFEtbFTVoF7MuVa05hqMmKADEJixPs3ipG3PVkueX/BkrxaycD
T+73iGlXDl4wfZ/n9ACe7RmsKBePnZLYS+l8fNJtqYcABadCaaUvN4i1Mg4Q5b0H
e6gWfUmTZIUZLOf74PMjY5YcPd/2GoQ7ArEGykI4nu+fqs65B3qTE0mhwJzY/EcB
s3JXg6AwlkPyz/0TrI1GdBWP7hxBPiKMdaUzpXYN3IbnlqoiST8RKOegvUbagoXO
4SvmV+fWzJ4O+uepmtQXlreEP9nvUf+48nZArxB98v8Jey0C/PDyCT4TM6WIAkFY
3hpqKM44hZgUg2qFeq7oJo5xGRUkRb3EMyuJj21+aEuGzWe3l+Q+kT9vUq7WWivj
8wLk1nP0me//2qXcOC0fjHF2FBfTZgIZsSCARAhCGZQU7U1pj7BGyvwX7ezbjctb
tYoydiV7KMcwaR2egKARZMmZ/mrwBeA3h26rC5+Oq76GUgSns9RLgE/RM88IimHh
gdwUAhUExLREocnJLCSMR66U0UM+MrasBK3oz14mpZMJcJ1ZE+9aapZCjIZzNoUs
WCTeJTZhXsb3dImjTxrcjykruYXnVcwZflzE5N1cIUFITtmW2JN25NsEsJhfdIv8
BCSYhUJquBmXmC7EA9hviZe0L3HbI76aDOw/kQL49djx4MYxkn0TexvfT15gQ+Yf
00SXft6JH4NUtLCzDyjj8PGkt4eW0SHeIF3t/SN8JiZHBCbIyAnH2hOEdcW8hMq4
cCET8tXWDCHF6cdutwcNWW4R73SeTtz+enzo3n8ZRXO6ddqsy9pX5aLahmh5l+Ou
c7ZzAXqfOz58sDyZwHoLv8Iwksg++AT41eyiKhYQzw3pa//i1RgHtCsoqdWmMC7w
HnKEeRmZdVe8VoVTtxPpvk9Rmskc+rWkxdYpouFtinrFAEpVaMIunSUMY9jXIJIR
E7FBhLfzgtL5tUVUpuSxRWiaR6xIBsRBw8eTABZ//hSzZazJuWjofEfe9hBD1F+3
x/EFk1uoLdTNWz6fy+r6E1RF2KFpf508xPh0ZEfel0DOmrqJJlCw7zl2R+Lkb7qf
8djl8V/kCTne4q7rqrh2a6B0D2AeoDEg786pgi69/DtfiCLhQBqz2LyOJPAD9XXW
MfDTuhc2QwnU/7Z00LONajN+rCMnwefOQAvj6fGCGoIznm8u8YS2b0scMNNwfsTn
LJw62ZI9FxDQYXy5OpecYfzi+OY5fZokqk7FG++RoNqtYpHWjFbAgdp3/8C40f7w
lrg2/hmjW58rFKOsm/kaTjb1inHhc496cumLODoeu4q/Y5nkDlOmlwnrjTTlijZi
4yGzzLKBBrygrDe5Van7IRQeaMmCRx7yIvDdkMafy1/3bQxkJRSQdOyN3lak6ILa
lzftQGFFymLR2RvTatwDU9xNm0wvvz4CPGI1Glbk2BeJ8Bh3hQk4tWqYIxzRovZ6
hyzd5YB+jC8TEmEK7wLCpgSqGZ2Aagw52MfOY2onp5D75Tl9dsfpjScbG/qt8BEv
1Q394JpggW0R1BOOLBDEgr0klofyz+aRJ7MK5HZhuWKtH5or8OC/hsybsY0zkJ6T
DZ7SdGuY2a2BsGk7Ritfo4kEjg6MWClwU+L4NPAO7pjKZZWys+4qUTV9UNvi4zTA
fOShduO8THTV6PBsihgFRkD5kMkI6jG13cC/Hx3lteQv8jWj+H7VY4ZjohX3fx38
X8+tzEsWEJZflIKxnTRLr/wZjHkCk4csS2gqTPDVSHdgUVbgm4dKmsdmNXgUEfjH
dC5yYJ+FbImNDIjqbTGGxeQAaQiaYXhka7L9a5AtvJtJGmV1/9hfnuKlO+NejqgD
miNoopBrw4MzoAAigl/zJ/jqeequpaHhliWsmd3g5dBzMjV53HpXEGNsbZn30OJa
JUqaCMH0E1EURd4ZmQXiA45AuqZIq1bh6gbAgzOl1ZF/ZIXzVsnrtfo0CEKVXI8W
K/nBgGcC3vkEykxedt5qEEcc2fhBMkQhhfBEhhRWeia2eHOKr9ERJMtLXnmXxd45
SLpriIVt320jOmsNq8W2HJ8us9wB64VVuEoyGgqLyUBLxU+9m6iKPX1HCdlYdXhW
K1DwThcEAGDcQToXJk/7mSlsvU4CsmHjbGhvlzxwYyu686qpaop8nFVs+F9RVtGq
jXiIb38V3bIxr4OXM7Xs2lC1TKuXgdnragUQGoPt4IL3HXvkyaYCFNTFgb3t8zDo
hQ8JzBBr1Zycwt4/GQtNBgXHd5BE2d4apWV9Ae+51CaEdHbhDD6JDJnHXXCUahNh
sfmmO7KSsrpaGpRVtSwDUJOIQYwZaZSKDsXlPuy0cSA6S+D0vec4UUQ8yRYccwMC
jjmCGbkQgTE8x9hfb19OyMPAt602WybGs6LkIr0P74ZTccqzBiLeqvoFahA2Ydv2
5W4dVK8Z8KjAFLKtJYswYn9HpQhwOBXFV5jPwXlYmV5DDPfkOj2F6YgN1fZ6hOl6
CrGPd/zXqg+4afTglQiyFwqiycj6oaNEZlwKAB3ckfXBkzGw97jSIOsbHK3wwVmc
d3iUydZY5AElO9x7+hKPlGQJw9Ujtseo6dpnARXsB5bZ8AM3KA1MkglIkdR0y+xa
ls8LDOi9/zIGXBpgAB7Uo2n6huwCz6h+FceF16J4/MGNSjdBNSCTwQVKgeqrttfI
R8yukKKraTU6XRPEESYDxvdKvw5IbrrIkdAu+KspVJ7SIo2WIvsSm2CUSgEyObo1
DK6MYQvQ6dYnct+Y+jePqK/e5HjLg7DlfjJluKv4/syD5pTZQ1yWQVJltjg0tMPl
u1ACavx8GRRYZTUBE3SSl2Bc6xUlxZRYk8CT8+0Ct8rWS/H0OLR62U0bom3ESZld
ao6MRWtT/ACD2juFYmHeAtNUzRY64FSLW1UWK2CDuNS4J0UgSyQyB147StMx/nvB
+Y/X23ldXNX8359kT2JIfEfqFeQ6mPt2EbAa6TTSOfrIM9/F7Js7mrOQ9Co5y1Y3
0dmrMmqgSlso1v9eeX/KA9ywoqWmK1MA2pbwfgMESXgUEsWgHQQ5ZIqbQXDFO4bs
Cw3bEkGCMgoTAcIgCOUjxa3YHug1gd7CJnTUS/enX4sXvS+WQrpEgzoABFqCFKeq
4vqtiUazkIqZNTgH4C89N8CM17PlE1jv8Xoh/MRlkAbaYCDbR+Da4fYuhmQ++eec
IgZDpP0IDtXfaeIPs8QDaaKuztqrlB6IqFdOuCRgd2z8JvhwGUNah+WGlDj8GXPw
YIrC6LW+WP/CNdMz5mF2GqYm0W3cRerkj2r9cIsiH4yViRT9S1hjIeurbqYLkNe8
HGkkkChxT8hTA3TxPbxkYFpP27BRY47qCFsELmKkyR0iZQtG4/PZ/dROdWsOL/nQ
6OkVS0HnZliu+m1PKy6YptivFTqKBr2vkNY+mSX/aiZncL/yUKqPARSME1G0a+Pw
qUtSPeyYuT4nMECqMjmipgcMbXGeFpkpCNI9Lh1YM/BqMJW44Uc1iw2850C8wr34
ZNNRBMDvXujrK6bjtfBbCpNtS3CYVJVtO3rp+xkAVKVdCc3XtS2ZhfvYK7w6qT6n
EYNCm5tHY9+63Plaw/UqNFHKJKdbQ2prC1dtzRaZCazqlf5hV6lS6dCa64/lnobM
9UUxqDmgG1YHm8JQqnlQGdJoDttjQ2PRBAiokxpVbNPDl6eG3CSdNSQea8bpfOI6
t7EwuoNl7EFSiy1hew042XUz3QbPcyvX4sESdilgV7hxlZ8kItYhC6oItXeBv9Tf
qzneOH80Iy9Nu14+NnIyxewdBeZ+CV5ztz6OqSrdXRw4lZq0uymA1Icdmy+7+a4m
j3B+z/GrzclcLz56bNh7HMrLoamruBlYfTedWpHsbZLncEG1GixWEPbj/av6a5mI
kjnguHMft1v708dI8iqAwqu9IMr/lYnVAoG6wUc+Wr/Tt0tywzKbLQe1GpbljKuq
7zLwGpJ5vzbnKIg2fl2rMlK1jtDietr+eBx6B/NMmYMOfzmE7FU9TkPjre9UFFsm
pLCZz7tKjh1kooYTPA75bAZQ5YJiV/sZmGkfS3wRvnr0ZdB0N9lpcNCiYFMYQcYw
EGGqQ5lNvCEr5edU1EWQGny/ZQ9ZRYvCSlwuhFI/EySyHph5LqJ4Bmva2DvTalf9
Npc4M8A2pL1Q1c0zX/vfGoJ+ctk/LqMf2JA9WeLyFtzQo5JT6wPIpxv6E0vbO/ba
kNjqzQi9Ba31sjy3BN9aAW76ErvaCun0+CuJXMDGNdyvvOPfP8l+88c7t1BzoHYS
TQvj0n/LibXGnCDH9IJHbIuEEyqW66Z3F/g93keXY9jhhYBv57qLpgY0ASIDvQHY
DN56ya+WenRkFpczO6SGJs5mQFzrFMUL4lJO4VGR+F3GSRtmK8dGfzxblZdDXDt0
MD1DMc0QsMe8bfQ4UPeBvg4AI91JqcKU2PcHuUwJ9H2ti3q01rEfWORhrXzr5a5L
Lf9n3LZ/KfdfAIZIYzG8Gpe6T7x99T58IiDTAf54NzUqVHg0M6jdy5NhJDMkhHLu
R0Gz0vMpu9zBWKG2oyKizMwrSGIjgItZZYzhrkfsC8iAWmu+B1e+L0U5PzD0kcHi
LoLthVan6ACY7QIZyYNdiA3Tx4FDILTLdb52/pKJEhH9GMV/SnK4nuGZp8AFH6AP
HbHF9gOlkPSvJZDBeESwuNwDFiAa3fg5tLOTqcEE0UkMDz0P+svscV4wiGr/PMCM
+5Uw/JAWtUa/sFjP80gsVpO9HqU+Gmhsqa3db5xsuRwjc43G5XvOXzgA+u3F9eWE
FOwxavHc9Hc9BTstjyyS08FOZUoGLrlSIjG/EnyPZwsm47Dw0Y85yRO1c5MJfCtV
3HQ4jQrIxmGqozdh1n9HBamEf32dTjZgUDCJsWa7nWh0lx1Ggu6XFUjTAL+Z5KiH
7u2sxAX5GUwiy4tI1TU+ds7/VHltzqAEV3LPI9J5mzOUPUV5zjUDtptXqByYwYHs
ChkZxhwEV8tEjRrpxHUHOjB/2HZ3qnoX4hLHK1XPD8idoHlbX9TehvkWOYRnjeVh
bLyYMGuF69Fx5Ei7KGZeVCuoOd1jdvzwZJuu5Sv+TrAJAqoElk0F8LJKM1413yv2
oGkCwltJyo5zCt5Vw5Fr2IGvKLycUvbLnxP1FGJstynh3qfsofiatCN0nVThGKeW
Wwngyv/aibPyzpkMV2bTa0zEN95MDH18aiIrT2E0keuuZGdHj46T2UcsfD/1fpSW
Pxjk4XxBwVTpzG5ovVH8FZcatN7aRj6wZqqqgAZrC5uaTtP+JuS8VIlDHh5Hk2kR
AJPdfo/Ai8DLPVpSx9H+clIuRUZrB/jfd64+/VhFJXs9B5IEixUgIe2PITCzH+DH
pU1rCKLcfCeB6rElzHCW/psV0o/LU65lDb3U/Qgab8J0Pt3yiadJUNmiTXSJOhk5
3DZyzGzFTrYkf1JsNolZ5lodN73QXzOMD22j8mPWrQt93wWOlLXdo6TncS+jpemV
2KN4QDmw6lpl3X4f5aVGPptiLPWXoJg7WY4hcngzT4qfNhMirn0jcydJqEvH5Y9k
YqDACf7urAAVGkgTyYejBZoBL87CPaJbBZ6zWVG8WMvNpR8Xynffu11xieDMzJQ7
LVT2uwTrHxf0WkjLkZnMXAv+nZcwGkgjFUCM8TSPHaDrijbPyDNsj3RyiJ0Le4BO
bSiDP1TwlLPiXGo5K9jhBUiCneBxySy/iesPbPX+om9aLB2+2jgTzifbW7aCyFD3
ncZtS4MBVyZHKVmozrevvDNIcY/Ei0rFtFL9phef6+QK/QmWlI87YsEabFn9Ee4V
5Yo3kNA2hvA07vathMcE5maiMOQn2RqVJsapjJVFQ57mSaECij2ST5ijojv90psu
FTz+CgnSgU+yWGDzzLfXDNz8DCLJHmHrI6VfhUrzJFfNucKeUcqSPi3VsiOewq8j
kUu1MPvV6+bRUKiL59i/aoYKz5P3TbxuCLO2eBEvzFndpcCAyh52VVvFF9Mr3OBq
yXrwKzIHGssaL5O51PWe4LH20AUDlLNONyRrqb4+R2e9B5HCcZWeoutkquK4PQ5U
SvOhnFwstoZbH5NxNWd0/TDJlMk4aCHdXYSQh6Xw99lSgYbLKANuUZNTRvsmR07x
mb2kcEseZB2qiKtHuXUdlu4LU+DrfLRCYS/+3gmQW1rwdnL+E7al9wq71kQbJDdP
T4O/rMrY000bnbYOTvGXPfJgOuvk1J3A6WWxgaTHzPIQeJVBX69twXaB+AVtQTVr
CgFCLid8CYambP+2yLjEHukf8NgK4qaJ4Y2cn159/kSyxV8kHFte7iMyR4HBkDbo
iYFO38RLZRX+yTgs4lqNYc9NmtIwkcVZdCqA5pGTOpVTt54q9RDQNihhERq5Y2wK
ghduBla6yV4l8m5DxJpLHuHIllKj4KDnGXvYnimqhl258mhNmTYCxdEoj4DmCzqP
IrRU2M3JgGquJs92bEBy/NlqreaSpmt7LZ1Yx+YXt6DSlEvMDAPSZH94YL1hvSb+
a+6M3yQkIKeYUZi92iFUgMsV/XbXUC4B42D5LM/maSfxlA4fkgBAHOL3DuI1BV3W
tjFirD02OMDWvvyDFB/PuDTLTvQnoOauX62nmIkWaIUFhD8VW/C+YY8lkAExdRI/
U4HVEmLZv+J2ukZbOJuULyYnh6rATtUVW/flKjW5pEmr9w5yaoxvlBWNhbDKIrC0
62rOJdShOcxzd8Ih4txYfechoBQ/tx2gpquejJVlgbtRNs8CWrYhc3ygYmwVoNCJ
8ZWJV4EUwuJ6ThYYIZuQ5zJ+yeX0YRo1p0l8pc1d+5/NtmsS22qq5dwAnqCtWN+I
Sae4tYCDDV38ca7cclk00wSXUiYYco7LXYy/3RAAgipmB3octZfFyXC7bioyCiWu
5cQVIakIymdGluwzf3wXsfjT8Syvo7Hs5fQpUcfim1XJ5n0Dxhhc4rAkwfBPez7S
M3h3xin+2Ejox0QKVA2tq9Fv3L2o9+zJ70t7oiFqQUkNy0DI4DPfBvf8kEk4CvxD
dWeTtaTgPS5vIt9WAXxF+wswnhLgXBAimaL21KNuUZ4jsQjeRPhScamFa03zrPqw
ZQu2w0qQRZ6JauosYfhX5bbavIxouJkU8Xs+I4VXSgtMmL7nA3mGlTdxAoSsDMkC
pTKirnAOV663Oi7d5vFOC5e3eE6RJMYktjP4waL7b2fi5SYAIuoSkqDyOrPhuBdE
oJ8AVncgEo8tFr92w2XIlJzmw3UTxn6T4sZ2CpfYFzHJV32vRw1h8oxrs0A6E2Ip
/Xj1VcKl/KRsXSmdAwLhwjFwxzi0k1PYp8iiCrDzfxZmRs4P9k1tOAX9WJL2mcm+
TNzUWCAqh5HEr2N9DeBi5nwtI1EcofJ7A/NQjtmRHT1DOKsEu3iTvbOQp4NXwfwi
2pPLo0FwVJU8dB1rToCkvVlT66Vqiq4+t62r6GtAfrrcEG/H6eDBshI48FeAPwOd
UQn+aqRH0DRJ4pmZyRqVlKLOOMDDfSDp0OBOzZ6Whgomy/VnJA3zaav6glzRh4OR
f4f7qxNFppyKeD0DuVCF5A9+83tTu5Oatf9nnF16h1qbBRmf6SeFAwiZJQZ8mU6X
EKV8mMX2S0a2pWdvafdnbyeoc7fEz96PMEjYJy95Uq7cEtFknaGLn0Xl9iXOw6ca
uRJ8idoh6gJQpD+wRjjURCna7nvT+Ha+6pFEBo1eFTrlUqbhSgxRuvlN4zsCPj53
1O13D0kArx30SVav0Ln9j1OIvUilmQykSeC+31nLmmzZwUCnSyRrwdMBB15BNy8r
szlwu/i8PcDnccKj+fn/5AVhv/wJ7h5rLHlHsICl3Edibx/2NGAwxtRfX+3yezX2
aDNtpFUkDpGDs3hPFl89Sv/aQX3+zO+SUl9zUNamss6JQlqX3HjStHMnP25adW6n
kfLGJbL8IJhEY/q2R22AO3+qUT6IFy0QKrzmMKEcK6nVRAl+scnd/wS53daCbpSK
QKQtesOd+xxFwn/pjgDerJDaeC0k4EfBexNMnmIDy+fieGJJo77HdTJm2EGaeLk8
xgxqfb4qBcgAfcopob4O7iVk5pA+Q3t0GyCOtfzBXFCw7Zg/8YrduHQui1Ye7Hb7
YzU9P0J5P2m77pxhV/XVoD/C8ziugAIJs4uBhir6gOuylRQKdLycK9Zc+IIooEhh
1L0hlCGHmLQtKR5iDglL+bqMkClXBi9tj1hEwf4dUMB/CGgAFIK5h1u9gwEj0KMs
0qaq8crsrvu61WPxyE4kYwppk8Rn/E8zQLCGQX5+2HCdD2oDxor2Kk8GYg92TV2t
y50HBEswMPUdGPH5Se9LWGgOPkZGX86qOe8lbKuqiNJdMci7DA8KqRH71JvDWTgz
2fq3+spPGXSz+eW6yIueD/ickQWZaOgrQ7VT4GndCyhtZM7JlJ2ll0GozL4xVuVp
ZCNCBAn39/oJmLFwt4Usm1SpJ2Bw4+ObXwvcURxFcsC/y1gSSXu/bQU8bU7e2e8Z
Mc5u1YSs2TwolmYqjV9QoNWbCmBeGS+t+QxLqGN+cExcMfNHN0P3GhV1bUchTwi+
pYo+cU3MaT3SawdDEMO5BoCEnmm18eYMIn+Vp+AgLP1E+koXOeUXmmC8lpcYn7PP
Fbm16F5munwiu44eakoHnhfXhNS38lWP9sQsxFcGyvtLqCwpIxH1mOMKIGTYTikH
fjTke1i1ynig8f2lUgh5heOthM9IPWSsmhNkgTxNOa5txd+4VIRJOLMh76PXJrXy
oBtbvgqP+MBgVra21hJ9AF8gquYy/Dn4AXhFZrfTrUilievi7S17EsYpZ5fziqsi
Zxq12tw5tHO0x+Tm4gnwF/nxQIN77XlZJo/Nt06IBxlew4HxrzeW79gPuvNI8KFB
CtCNFWlE0gQbQqXg1eVLnkfwNwu6rbg+G2UgHlEAk6f3+y5UL0oGRO0Xuz1/0mE7
uL5KpSVII3n36dVmhwW8RxZeGBp7U9eCnDL9zPO06QR9uMJab/P4d0UgXwn3HqYE
f0Z1ET5Bmsm6OUWPQtlEfHwU3lcfIVKyhd0qzTK2MRv0yWmrwVpt/1kKtaNjXI0d
fWQlNtZFR+WChE6wus7UTsFVdABV6OyvFM7YAEuRhaHfsHfHH+MHdC1atO2QNvod
XR82U7lICLEVER3lfefn3SRJ1gn3vPwPKecAJ4I+eUi5Ly8OVrP4DqI2aCU7kWyy
91XVNFC3jbXBxzpGP9BIEBsWKJDukabAgZRUSPUyz33GhsvbycpNh+INmu70y4/R
kbwHknvYjhjwfA+waXQXnKN23YtxUggoOQ/HnddI7oT5t2TuGRpEBlpYtWVh8cU3
nSt/0nMAkfTlwVy37dGXf8nnmNhuk1U8YdSqozajsm6H2ybWySI8KqjiFzQisfC6
TsJ35veYZbOCnUJ5t6LLz3RjkxbO4lVMBRTuHlRdvNEiFnrGc2v7imVHK7ieVEu9
iTXHj9TYBdaJdMYRqQNXrfLdx0DkLzoiCvlhvQo9EYsE3Kx9UtlB2xpo59ZUcLCe
7YPehVDKDLodwR1XER4RCi0r7cxa/b+1wKdEs6JoJfyybYFFklcb8glRlwUrW9Sa
dZOHybozkLk212zxOEwlhH+RmIQ5lxFpk7bFtTR6zlZzg/VKlVBzYN+1q5TLiBXY
m46WauoAMGgHna0A7sz+eUVkK9ULC+gR9O135eY2GPnxdhqOWUvh9Hg7iRLlypYl
oRu3gzyEALhOhPkq4VZs6iJPyEFEaVEb+GzSdupP9f6dh5RzVPuT0XkBZt5hoIpa
czKstUINh4paaJHfm82QgxFv675AEuaSA0AGdg04zKGRykacxvlcfFvQpo5uH59+
9ZEXxsjN2IRtRFN2USWDz+xgECsqF2qzAd7/yk9F7rU3Ma9CS1hZ7YQ3a/2FcDWG
zbQgoOaBfkleVrxqWB4aAW6P3HUypnaa8lKXif0QM/KrRz62+RAsl1w7bdBVZUwc
TuCcZavprrphPwmzMffxoP5E0vlE4/VdlRwfuZKgyozzQO+WRsFTOIwjnVo3LOVa
zz427mMbGa+c3t13OQ1tbBzNRpbMc5oYgH7HcaTlhv1HZro19kT+P1L0cXvCR8DI
7AyxjK3dtMfm3TMDIF6m2evZl+uZyTKsSItZS6XIJ9E6PVEi3Z2tFXRNbyvwu0E4
0MrmCm+6O2jozFEOkhR8sp3evLPeYQrWo2pnJzxtYXBrimOboN9AVgeYoP+ahjoM
kmTPRGfISfVy8UY04AVm0ttkusdcj2TfsijVy/yJOV7EbiwG3xI4kbYxKOhgTfJw
ow6E0L23FbHceras74MQEzT3uxGTqnVy5t37sJWuHZDD28arbMdQXgaNxsVZUxDB
XY4M/eXM3dX/UBDb0AP/hxu0rPwkbsuXXsXYJo3HvqK2SxPzW4Nv1l1aiqah4K/4
ult8wuRdZQM+Wm8GOEUNFSbJ5YXoeHehp7+PA1imCnwRE4LKUE1sfWHKt3U0/PTQ
N2LMQoXHtIlRO1r9msxvYbsrKSxN3u48MZerou3++WqsglUSWLQqgIjgNHOLnulB
YQdlQZ2NpoWJ10XQ3gdq02ofZ+iNpboPMYYGL4mkO1hz9DJ8UBo/I1FGa+oCoV/M
RKLn/HBIh5YJCzuHHALjdPIeEljfeOslhi65vOIbOwitJGV8ZmBe22shsKenjoz2
RXqdaP71yV/JPh5ksAjSGbXFVd+e/OZO3PtQ/xhgMtiKR/G5g0cGRDvL4jR0VmxT
CgRM332IUteAQ3cnVMc8aqZIORk5jPNurSfAE+uUPVVAaLSHnLlHLpJvvMIfxpa1
/S/xFLBkokFEl34O6JNRRIFXDF0zbNyoscSMqb5xAInBTeOxSZi8Pa1a1ldzWv5N
cWCuS5BDoqUDMF88oBPY6o0kNbbAwyX2zvZcId8ZXebhJjWK4YVoqBii11RSWbRO
aimDCHqw/TVogX6LjM90s5yCWDzZssGW4sAYA/uNew15s1oXUXqAXqOZ7KdQarSY
PHFWoKDO5q5D5xHNr7gKuit7ZBcxRTeHjg64XsbnsRa4KNwxH9fw6tOWUeGHbXKG
/bLfsHN7QW4lgIO8vVlw/qlSoJ4tTf59+XiQS0g6f8oLk6vzkE+q2aDr25KxptY7
wgK8UAHB6ZJm4Pdtg5aS3zRMK4Hv07XC9pAoIzqOi2tNNto79PHAybtJtwCTs3S4
yAaXBYRk9YfeF4FUQ8CXFTG2S9atNxB7v5jUYrGLf28VethMplbJinWR353l9wBw
bY3Gsc6Tq5ar/5pUz3RfBagT9bzlX8dgV8B2eHGau9no8QUFBqMhtvjbOnOw5snC
L0f3y0k8Jg/k0apUNwOL77scJMfBEf2XSPR2uZbCbeVsJEbRtMNeH/MjOLItm2LG
iNXsI8dd00v+/T+baA+BSn5MjQnTbRyu0SN9EWUA9y6yQjfao21rCczSTaoGT6i2
wjS7mAz5MrvznTE4M7WVA4NVff1e4h4L7LGtc2b89Aw1Sv8hR5FZrPbZQAryF/oo
GCNftFETi328w+ITLkEXzsYGqW/zbQXlxH0g4SfMjK4mrMXYX75ed1QqnLlOu904
S0XpYmHHRw93RH8FCGTXsHJgjKK6lrSKZz+ywAx+WOlDzAU3TkZ6SXfOfCNcxroz
qpdsZA5wP+tTLhH4eYkT4XIfd9MJzlFtdW+blLompmiWeiA9Di91Q/FI8BqAJ6RH
rA5uB0h1VbyxM9wf8nmN935jRdQ9jf0+q4vfd2i50H1rgbbG8vLSznMWZkMD3rsa
r2lJyKaDWyM4J+yg6iPi43WV7rIejaBSUP3UX7Ky2VdMIfwCwDbO7rlTGRLbvSd2
OmSzg3K26cF3WBsEzOpteJb+DAsBtEK2ww8YM5uzKgNunLsqglZhFHxHXNBbiygy
eTWrSJbrzb74nkITiWsuIjReDepNz5c/P8okG5RsD0FmWXL94ax0W/mQSmvzaGad
tYkyMHhSyR3Jy8hgUCFgmsn1Vf5nSB/YXzcNuG0Uir2VhEAlSn4MKHp0CVZX2CtW
kd16s+6UEXCNXOkT4JXCO953h3OI7TCIkv/W0gbaS+Na7krZV0DJeT378RwdYGoR
Bqma9+MKcuimNzqk3YJAIaZh1lOFimPhjuDPSRf65uceKvJpnw+kGKTqYSxulkbJ
Agt9svZLF2GDJJda4/j2QwuUkVdDJRYwvOhVLxAaGFwxFkFP3ogUqrsMgZpbAvJD
THmxu8ax/FWP/7P2qhT76rck5ghy5yFk0CtEHKmR8nZhBHikGLvt9ozQreeGbwtz
BUKIxB3n+X1FIJH254yI4o1tOb1bI3YyQMxZ0bgATLfPt2NRMO9JrC9YPN8L8lkB
MUT8XsuOqDD0YRy6iDli99KJ+yEIg/Z0lAOYzdo3Naf8fnXlx3Mhn1qaa6tfNcnd
oTNx+62nd1GGoalZGiAjBHKn7uOQSq7S/BNE64nBGRku5ABhDTDmQe+P0L/9PCWk
bZGfS5dlwNchz5sWgujgee/DYgCOSISZacdn4ZZkOYrcYqG4dhcJbHVC4HTomVl5
Xj9PvE7iIUvUVa7NS462BRzy6hVLp2emyUmU1GAhELabr3+8b2Csoksd25t+pr9v
EGLKMPjLd1QKxEhTlon1YCR5ZqBOHSILyPNL/S4vnrHIwGTJ1xBmxT8BuvFrp/4P
YK1XLuLu70huLzwnwoK7uZ0cRgKRdPUyBRf8vc1v22vX+2QK4EkTx6TrqjdQIAGD
2AYvlbOw5Us8fICG7e9wAz4elM1jfMB778D9QdHKN0TlSR36aFKuqg6oXrliTarG
CcIOgnsmDY3TZbxSNhzR12uerJ0muCCuD09Xeir27tyZeXlHHT3FhBlWJtS5Knex
kTyxryYwBI/hWnwCPJDWETFxWZcsteCEqj0h37NIC/aTgzFmGV73KpH77f2ovnRP
qIa63ZBz4hMI3O3iQInWh95v8gi224P2SZBfJjDM/pCw0vvRdTxAuKqX0ls4oHmP
MZiEd1G0nvB9Z0fkBw5f9CoSEkC1fP2WBwyDt3nN3b1OFMZegj9vgqFo8ZLe0BjT
atxF8VL2wcaQF5ByXXY8iyurLNFA14n6odSvFL2IOBPHV+PL1bMqTLqbzoU8ExeL
UZHU6e1B6DtMmCbhZtIZPOkYyzd9FJ5JoQ3N+3CTy42r+UUOgIrKsif6rkTcBx8+
aUqzCYv7SCbexfxkk64gawRi2HUKqT8oFa/4bkEdhMCkAAkUTdbKAZG+V8lxtiGy
q0Ta/9SH68j3ONBnwT5d2bhXwBRed/08Zv3PR2m8/yD7uFf8E6Qoj8kfDRat9YIj
uZfRZCDT5klibSWVww4H13hLY2d+DTPy8hb4LcpFx5vTyVWhXX4FZKvXXXDg1ARe
3awmtyN9iIYiywq+ffG5C5tFoJYFXSrLstLvh/UvlrCFNu09VJgjp9ALpjPbG+18
Z2C5+jq72QJrp5uxifGVtcQfqdEBT8mds99fkJgYhGXPgldY13aibgEclzwm9Msy
RyGydy9JNixZRB69P1agnOZQSe7dzfJNPRb+OMbW76S34Ppi/qjgy/vNcuddFHeA
Gh1HbCQAM3lgKyxt+DYXynJJcFj1kD/mAOw0AxkuFaKtKscFaxgqoOFufTSWgs0I
vlS9dDBR7Up65cyKq3/mdoiy1HpQB2KGQSkqYhkQyH2bTMQTF4LmW4JL2ixjl+qJ
hS8TtYMrI7p6MrvRbDqoEIYn+7ZBopZTGp9E1OPPasAm4ap0JnWCtIRL6rDMPeh+
QXGCqigssARoUBVtTFVmxfRy0IjdMQaYLsvYGDk/7+HLxlgZa2IGyhAifZJb8PcG
u0zRnJPrYjK+cpLC4Udq8az4GI54ZAp0+UGv1Vqa18RcgsAro2ct5ciHS88nps/4
o8dq5sevx9mIRjijg0y44PMCX7C43cfXQu1F5MVvCqMwgwllcLWazDYyko2OJ5tm
HLdlkAEalyr6KeZE2Up9midWifm4ad1LfTO1C0PFA7KIpXcmwZYn1fURjrbmqhop
3JjWzCreTYS49OLY8fupBw/EINM7J1I9pEgHnMNDQzExL5qspg+LhPHu6x8O+eDT
xuxwVS+zAoocN6CX95ilWe6D/oKLw/qaEyJ7v+eqVKcWjafrEYWK7mUuUj0sMlsq
T3PRtAaaQpRQDt+6datBoa7v9bQ+lWNq22w4PyyLeI1gkAArq6j/b60TN/2AeA05
4Ldicyx8VEZt3AWDgytSeOsLt0/jf0gah7Vs73SQk8WifzZTXdyhRm1pGf/v/Y4M
NICQlXkUuLcTY0Vv4/8SHUcWCw8SgTqP5Kw0+9GiUn83eoJIv2unByQTiv4OoIAj
RwiEJAuubTF1+FRLm4zEKT0J0YutEvN+XKKo9eb5Xc1CEQhc29rwTtqwDmthVrMb
1R1A8MsY0gwUNCZ6QN6eHqZ3ie0hOD6clgZsvWUb9GdMDvY2hjPiRm8v4qFsxiWL
6HkIvqNHx52JQ8w+2WjuZeQCzKU6mCsCv7bHpeuH7L6c0jUmxOK2rpqAH32xhu+0
pBZ0pWl7lIzSoi8qhuDEKvOr2KfW5Ks2SeU41ZNxxCjo1RDl3HF0dZSIsuTxl2nH
0nnllznaqINH9VeWjHchE4ILbpLO+0jWGs3/vyutk0gX2GIfkK1BTmP/MvAX4oK1
zVPp1dKuNCKdbDGXc2Gifqv/5RYX0g4ajUny12zT58UBKexMW2Aglmdn3MnSJwrX
PS8jMO4Sn2ij/LVaGkBC0Hc60kW4KYEjMcxxottwsVzks782DsHQa/wC2OQJyPGW
AEGF57xCizQyN5eY+oAu1MefYi4w09/youIG1CXLYgCaVc4ulp48u6/kmFs1yR3A
uamwbScg0e1EyL5+DOnrr9u1iNaSPDBp1FQhjCdx4FKbT5f6gH38UFuHMmmOwOBj
miqIAQYBMWZRlcCZQlEb97zQfLgZ7QhugBMe+BmSnx6YjpiSWMSF+SZbtSNai2nj
/NCE2LD38QU4rqpmPS4Sg56xAHwmKDJuBlhlzfyqWtJbYFzbVYdVi0CvvnhbnSeT
7kyfAHwAGRljwdQ41Bf5xBLyM8Z6SNUs8BURB71QkEfQOmiqgbXsZeC5ohbu4eJN
GIBWDLWYC3nBF/KbXt7jv2SXk1NyF8sS+VmkE2LWP7O6fT4X21FMh8IbhyFqW0fX
h9FUj2xYY3voZacnNby1gjOtiCNXEgM8Pz51V0S7FErBWt6ttiirbrnC+baUwwzF
bBb6RJ8Gole8MSiLSLwPZHLhJLJgPZH7tzMzCjkf+1SVbY8Qj0C+hq9jQ0b5bWv1
sDYFyGO6vmYUlCntCpdsLaIGBy80gJrPpamv6hUcagfO5RHrEgWLgg2LIhMvf1dD
2qVqKhJO0HRJCFxrVl0Qts2grW+KYkpH0FBnWfsyqcy5RBYQ3Tn3xmMcjAojD2i/
geBYPyHK4VNkuSIT5awAe99yl3m+wThGwNEtFA2afjQnDajIz0I6TeDSocRXkOKY
o5appY41Dh1fCwv/ZVgt0PH7pq9JY5KYZ+MwUPNnLlCUj8wsiImz95lL6otCW21o
8SBXTJ9G+rXFKJdx4clkdDfkB3/CVEgWLJPkj4uyodHEuI1UQ6Vlq+FTPTON4s+E
CtajFsXnqTsJw5xjw1rBo9EQ06FWYmz2fO9Dssp8wXT/8GCeykQg+RcFUUobnaK+
lXyg4wL3PeIFde1Spqz/GG92+7Is2LMc+0s1qNNDfY3si4tmY2FtKe+nEkfzj299
vn6YdZ0crWLGlXq9udP3EaFWEQek+VfOV42A/UNZOJx3d0npzFfD/78jkcKEPNxl
f2hTnvVDJ8ZxKdkY6txVEMUNzMs7zAB6spIE/g/N8+P7mEQ0XD9GSeMX+hOUW0lU
9HTtQpkhIeissO2yd/84+3kC5KbJPrTCT8P6LQRP8DkqM0vS8tDwkpW+hfHfHjgZ
jUfYpLcX5J22RXzTt++YNIf4zhTSEaOENos/u8CyPuN4CGsf6a3m+7ajhnP2vu+Q
Y8saygapuFw7Gu3eBINOjrhUkN53dypb4FMZFJdMevV+o/7/JxbIzBy2X9lm+4y+
Bgk9P1IDWQKLr9WutsQKj2r8M9QeDOCGIMAe9lLpT0SgcTdF4+gD+jLkHcdQeegu
8uATwQRutza8DqnMjflzgSX7JTa2XVi7aXs0g7SQlOLzELr/gp9Ebqr5L3GykCN7
aqa7BCOHR5Nkt+67v2AP0M2kvEc3Tni46eyWNM8rATrWInixjMwZcaXowyqzxhUU
F69w8LsumjFvnWEUr4o9r7swc5fL0/VR4KzxjgL+UJUCj5mKECJnVdXqfc4x+9Jb
faAuF345m/iF3dILwC6xu57zRS+dGlStlFXz+TuVR50uH6SSM9K6qvAGVGtm/qb2
r7AReqUDDxGih4K+uaOEP9c0iWoFGNGAnupcjRkNoCRv/lMMi+WeLlPMkK7WT/2y
drkZjXGGivHYR7XU9A//eaEvzOHsq1qZutPTewVhHK++T/M5FtTEx2McITqc6DBS
/hhjNUt8ag2mjS0hIJtBBHMGl2m82FZKE/yi4XXok4GXPip0p5M+w+1W2GSuk4y8
BUd+zjeosmPbiH4+mKstrnvZLJrC4OuPa0W3pjq7VvzF8Y/JcxnDkntbcA+5DYwF
iEHkr8Ayp3Oh/rFvVNDewoaEqYNd8wGFZ+VZgquCznjbfVz8i6gq2A7AuyJxsrvS
iV64pg8PtOT+Q8SLCe9gB5e7I3+t7zY2A81hWPRZLCgg9hq5QNpRZO8Y2dOf1fwv
qy5yHet6A4ADgL0wv4pXZB9ZSCQWaZto2eDIatWzqtyayN/LlEpiZ1gB4Xamcwv0
ufuO0UvndoxAl6cF0LAspjwTy3v3npl+gW8Lvok2A2HTqektgona5be2SQvdxDE8
lh+Q7OomAdyNnF4fxHy+ppESfRLNMZBtVb2si/j0n9Exec3+LjZusrbH1NSCy/mF
Z9oZAHF2mOqpfbJ+TEVSrSrFtEJd0hi/dIWXXvkOV8enJ+WfwdCGl+PmqgfO2iy7
7LIbgxnha+WrEUh75NYoJKXw7Oze+38QikGxd+2677RhWI/GVT6Btd4lMPFwQCDu
LP/iJJVzECDo4sbtdT8CWy5EATSSnP+nrUPLlpG4r3OY7Ct5VQh7NXgi1Udw5nd1
d2O3YSoEZvypZgtpW8W3bVRMliT+uzxVEK9GzvjFXlZd5HTIE12P+zzAnbrjwN8/
iDw4vmDaOv/5pvH/tG1mDur5B7adMf5GLKQS8xJakfTQrPfT6W1yFuaos6YPKLab
ox9O3wRI2ec7BfAsL9185jgnBDEInXstORWpJU1qShyZPGvwixmyM5usNOrj9X+O
8jWk3RmxhSjzWjweO18rNH571bewGgVgqfPn5v7kN05NMKxYusJ7UkLFeini5YT6
qkADb7qL7yzQv64Hoyuupipvh8zaqLtiF1zBC57FaSOiUbHTAaSbggj5v3J+kqvH
B7Xp7JCrOkr+tAK6IGDSJ4khQAipkJGFDzdYuiighUfHUlDU/tB6DylSdLmGxWO4
KcT5ESh1jmidqXdSRobSaRyhBpSI9cz1+y9F5hIrxv37eqbwkVdJyvwnHKRsDTNL
x4vo+hgKTPNsFhmBmIeR3XUtqbq8WbuHgCQNFvJBKsNSRr3J6a62DfwaB4JmM8qx
KD+vazP7aaQCnsVCIEPdhYbgQ3GpxUJBLQ+uRWJ21C4QHRVQT2lyGJMVtkoc/HcX
2xG3wLrnLdPKHBBKgALUrWuEY8jo807GYCX1/GlAX53baGsVe5DoCSNccIUkdNl+
6kBOjCd1Ho3ZFuX4IUkc6CsEoWMSD4IPItnKRYeplvv4evWCm6TqbEWM8ka16oKm
8TwLtT62ESRDVix04hUWOjmL92ZsDPztdT0CH9hnZYqroOj2AYhmddCNUZ27oziB
56bggtFA1qRMHANqLbPQmOvhn6fEeJ/bEPMSy8hPvg+bMbbSaYgs28VQrdUwOgXZ
xIfZiT/NF11zhJ/lFm+jINvj1Fayzj/If7wWKaWfTPGB5+EWsBXnqBVA6HUIlS5l
pDDlJDqugEgyyuE1ZYH/9mDfX+gRAXyZDroTtvRVSIeHh8OtI69MSVgMTzaJuqe/
r2mWmushx6sDKVLJBJS9OGvftDFlw9bkxsASQeEIVfTwBvcSsLfxxSkSxiy4LIWm
9Hrk/mh5MmnNVD7x4yBfVT2SLBFpInpFlWs4+sqBDsR8a8VdN5lZso7Zo7HSaiji
EHu6bGoES2f7QimMkHlevesI7kR8sYHWCFefRhrX2SJQr+zodys/kwKIlcGKLeBS
SByjo7K+wmYYzUl3VADC7W+bIUL4gnXmXQ+9yEyT/jrzcW10darF4enbeCGgA5J1
nO1In8YiN89unTCNVP2RN1F/Cg522J/88rBwXix5SBk6k2OjCmCjDyqO34J8txqQ
g6znnXqRd3/qnN2GzShXJBJcKNnIz0WKe06SobXsvigxzQWEB+8bD0OIbFiQfBqp
7j/pwNveXrAdVCA/UVazLlDgGBU+MHKY9hgvg/UPTRMs+OnPecWqOrCRz0kYH2RU
vfWdChHebw3yp4J74w1NEM9ROcM8T2D6c5pAhscyT7VaXfCwZsSTmIVQXV51kfi2
c0RPForjC2QxfwFv5KGMX8GKB3mJuBOZSSG1Ks4QJojKElfePN9ydnrzGPLyNPJG
0RlJS7OPikhWXqwZH5LFUNMGj3P+iVMVG4FLZ+lAi3Pt+SHtnDKJAqo5UxlBYXZC
CimvNGyoAfSJWWD6AEwl8omeR/Az17PjQQ7l5JJwqYlOY4Knv0HdXyTD/FPrhrQl
AD7b4dBkolZ8CLcfYI0PYh8ebDM14jjl6W56RY3LQqz1ANwig4p0DOAaRcGjMuYW
DB6cZ6+XIdcNN/8Frl9EaUIZHv0ET2vFGGZWCtWDcxCA9b0nyq86VFT405AfChnD
gBaR1C+OdjHswRm3AMyY70snQyjTxbXlgy7cZ/sPvAsrc+DQL53/zBdhv66g+iOy
xXGudOwivUQ/mTyw8W4YICquojQMZ8StcOyBWu6ehIXtX/USkXb5bOWW9ef0iveJ
kmbL3aqHZYpdvl2BvA1Q5QQTcSFmCf6J1Q9DcxHx0v9O+2rUzgqr07LeGKjV3swu
1Kg7N4VgpCCTHAxUVUFXkYDWYiFCpaDATYM/y50m+MdmdUf8vgcnoZAg42sAsaYQ
xz4Lt1yZo0gCOf2X6H/eqz6Cq+6anQCBjrInZOI8QoqPMasJIAE81AXqGiKmzdlW
ITj0nBfgwHA/Z0v6cPbdhhNKsOO2ki0ZKHyvjGxchZRt8xEnUQ5MkY1RgliUUf4g
ZOxNyx9SkcYM5+lo6Um7OcoaVs9Rjjp/xZkAkkUHR37PN3PYv/sB6kGbBhyzjdbs
j/O9rDDYOq/MtbBrYQjv1baeWs71M/4/n54DaFAeRLHN4o+zg49eR8OSOiHp6uwo
acvIDHNaIxHQRI3WaazhRoeUloZpCopWr7ME50RagrVTHF0mazPvMIG6RlsWMi0b
DBn+QtV3qBWhN1zqjxsMngIiwKUBDkZCAKkPPPjqFsC19UVlUg/U5LvWnWkFknxi
RcLt611/fUOvyZgqj2iTItFjGRiXonExVPBVq6OgOpfqnMUcyAuWJzWDQ8RIv3yP
+mtSQf21BxnGJ9Gvs72ewUOes4fQAksTOzIgZ9d7QcIIKJZoVS6F3iXaLpXvBWas
Vev6grs5td8DUSmbrrB4Pgrte8ilxvTHcEN/yYpMMQIP0EEFFN45uBsWjd31MsHn
ZNAP2TtdEbuSUUxSYXSCFzrbtTrUndh+el7FNrrmJBeyCpibqoVMru4OwwoQaal5
oWX3hXOS41Q077L/3bcnuIROKLNC61yE/F9rkeDOhw33tiBuN3IjdUMZTGh+82RV
21Ucx+2083tuHIJ/1RqazSdJbWe8UUG3E6Eocq9psEP+iIZCdmHVa6vmUEEUZgQW
nu94dp8z+096WFS1ZsCIMOwJeEuBmELqijWXPzT/Grpp+uaHgkGL8BWdE48NVCVs
+8ba9Gky8tS7l3q9ap5k8EIwBeu3zGVm4R73r2rUReGkdktZOkWuB8PRHgNJ+06y
I3lO/7iA72sOeDcU0IulTBW7HW3v3nN3A0pe8MDWBJEd4p+oyxAfeZngC8oIYvTd
nwYqr8XcghFvZreQsoXQ1me+1hC3uOykya3uqNPOC92lszUhifQnq4HcKKJnJUMF
4MG8MnoAy6CGDXB8w0DTUksFKzNISms4R6I3zKSWcgBvMMTvh85c6tPnamE/VaNR
3mKlghpo2zH04FFwPp5BDtpLN+bAW+VSJ9r7K7QUf9l5RHs6z3RClc/a9R+Mgqif
+OnuFKaJAbmea5/H/of4U+wQYkabYuCyYqSLOlUmsqHFygqrhRdLFXIL+ETfaxMa
6cwQlyXTzX8rOiPz7GyXb6HMyXMJ7GfGpr25Q1gkwAA9YPYdBNYoc8GzeMPZJRTZ
pe7R7bZH/ICafMhy2JGWYj/FwsG6ATQk9dXnpIlBiOw8zncj4BhlsXuBQrfvUPDE
Ruo4U1j8FX8Noe8jVuGM3sMV5jsJN39qVZBLGxvP4tgXzWs6gBbhUar6IeXnkxDA
ydAaoSl6jbZvAB/CNIm5SMi35GZwF7iyTUKm7MtyzBS0omCGQv1tvvzckf/JLf/n
/YCjyHY42uxpbj/pXZDm6xzL1ecbI51Wd1YwmR567vhenSYIIEEdjgM2MDnfTe6C
R5W/XkYm12Iem1hE1weqFUh6W1fD6bi1kclmsppVFItpvDif6KNBvrGS2LMuj7TP
mGqz5RJdDth+YtZl5nxgFj+vaA1CiGtx7aGfVNxNCXaKFl6krw0qBJdydywJiKXC
rl96oLu9Y3XNBoty6ez16RlieiMPuKO4QvIAIr88ozRbGVdTsOE9coKbL7qvzapp
6HkCcO/gOJQJzdDk+dCKxGkPx3xWmajJZUQBbzN312gzgJ07jsd13JpP2oQYc7xA
Tjoje+rcWxl0P7hZl4uPfPwKerBhFtOZ1hXpE9QVmD0fSRz99n3VrIqq/hyrJE4i
zlAo3yVOt2e8xaA4jLKkhpLpcZMgKYXu5+7L8RZ0S472/EwfqkxRlO2SYoLyhLJT
D4iMwcMTqZHQkUKm+wYlHbM3+FGyCKuEqTwkXA7RHRbXCl9EDtFvr37V9guChtOD
UkdFULpm/rhf5YXL90uYPfi44h2lm7BqJWx3h3/D1oT0XtAa3sX/BxK0/jyS05H5
Z6ZPfz0zoVf9X7KYPLjDatjzfvyi/+WZInlwe1MsR5KtRaO+w9Tu1+ZTY5ejmr7m
JfaM4Zqfl12Dzrs9unEnaHYzH71wC9ta8g8ZTc87JR2gP51pNrhCkuvdzBkO9ZJY
4EesgYrWQEQGk8XTWh6az10UPQKWoMtMSXeTUVIQa90Q6w3E+9ch+vNKi6PNX6Gb
9KmcyKSxydUBETNqPApN4QxEbouB+CaGs34hlEBWJZMEw9ADvvpRq0qxsHYZZJVQ
c18cnjnisZCSzTJu9tzZsgZmXKZyEVxcjY9/AexvWa/Jub222194eyR+oTwCcDzP
fz7k/l1kKAv26E767Dghu3UYgM2Dk786HcesxrVL6x9SevlLScCRKKkZL2zsWT59
XiaFoOf7l02tQpuANbA1I3kNz8J1Lh+PLJmUOigyk0uyTW9n+Z9IM8RdJZBoxPM+
uhThg/1v7Oopat4ZDiG35bV21AspeSQ+9j1oCvpoAmjKN9XmZs6GXijuhO2+GU+Q
6i8fMKwgKcSHOKd9Ot1enS5eu8lyqHjj0bedbiZXZghzbDVIlPmZcwsWs5O/chr+
ZUD3ImatPUs21CvPCWrOqU56LyyVIc5z076W+A43erxm2WWlZO/pQMYbgm5bNpTC
0bCL+DnrcIQqP98W/TP9Qk3mByvoNC0I4gVxlbg4XsLY8gdqXyVOEJ8JOjixAsDf
Wc5hkinjgRBcjrdhP0ibJvjUmWDSwqIu6Xzbzzr1dOiyLibk1eNGZcWMYvgevVGy
76gsg1fduxXIq+9xvjolzcNtMoJtH93LK43cTMqp+wVxE/C5z2hk4My0ZOf7iwSe
RRWydMQ4ckkjxXafh16ob/zX8mirBBtuHEXqJVPnPuoD8p+h+UtkOlBUEWhypKlA
hdOdyhpUiicZfjCkUJVKABTf3GLCKmI8BfTqUOM10BmoceSZbjABxVEplBsGnZ2t
eFLKXOO+1UsFD+MjXurMpV5vh4UfyD7nvaBfABc0ylG1y00v4FgJbluSLmK1TONj
Ne/3lgtV7ER3uKbXFM4qsBuvfPb1XoBsrmHyQVyVo7e2TN9h4rZTnFJkORMPnFwN
G4y9Aj16TN6lMjXYR66waive1HvRhjJ8IaqXeKrAxhUwpkB4qdbuKFwjiOfF4p0q
0/ZUUPcwraxYXLO5JiqmvkHUUBumg1jO0iEMuWrVZuFfqbRdV9D2k0lsiUyotqJS
l0egkrjbNuzbuaYJhEq8SbrQbRN6lQt4ny2IHGyOf47o8cu0aSbCQ/84A5yF/8eX
ZBaRjVdf0YwGY0yqmisPgod7LR3LWutHiI0APW+LWPI83D9ao8W9ATPckzmWQAp4
4CQxkpvVQcKrMYH1uAx00u1oNHreyD366z6n8pVJteUPFzb0YoFVyqbnsD1wAZ66
5hooU/BB3ulDNpX3o3ysrToMsWIu5+hF+mRb7Z+IaFCBQAo1rT08Sx9SQ38Ofbio
QFyQtBhcGmFcixjIV95JcYEF9dUcXKEz7LJb1l3PyYwcYKCgKyMqdaqm7IiZgM/z
7JOMspD4nnKt7/MjyHupxjxJhP1GZq0C8WU8lkwWLDT81trIK1eXWe4wTK8Hrapg
AOqJq59okrhie1DNctYHLOkg+8NfnXUezx5Pqk9SrEwVQnv0tHrQbx0TSIjqyuIR
D+X/OQitcVfdtIRsMVIBT+dV+ELLlazi0XMdPPhSWX9/LQ5p5TGJwRQ2biePLR7q
if4mqVwhAAPltV+ibwKYKVEDItrI/rWi49RHl0x8107pWAgsq+yuL0SF54jsTSst
Sbr5Y+ZVxocgxK1/sbCTf8BEyQHS3P9atYNuh3ev5bYKyBpjEfFS12EXq4O4P6d6
tomYByr7PHWBoh96G8x4W9FZNppGWIjcyTRFl+nXvG6YUOa7wcTnTFB+M+9fAX4I
JkBfT+3KOxq6iDn9TmyAtova7x+cp0UCdpnPHiJfdTuxewfkPlC9hfEAUnEBjH8Z
rPLHjK+KQCpllzCSUnzx4Qv7wcVlcgKTHq+sCa3xqQ9q7dAK/BNkpfpL+bF6ZgZt
C5d16nMPyjHbzisC9BAeH2cQZEgSyUHo5FyEYBhhKKL0Iyb1xN2rx9SjZhqBvDB0
A3EuhHqb7DbSSXeOkQXnpJgqCInpe5MMSg3C7zL0M492fafVgsDssNOO4bgOerLy
SdjWkjKLN3fMyAtbhIbmzdVsWyrv8JisETZI2jHeYXnrXY/bUjrJUqHdic2f0/Ab
P11EXtU639HOabhq+70lv4c60H2jGMEDMc6cIg8XJOFeoQd2Zx5/dp7FJkMzWXMc
bwUGQwgKxd5aiFr5p36ogloX1HOUrSb8uoChPKHykoQT+VHc9rn2iovx1RPl88tX
Aaig9by8YPWjhrg9uvF+6mceSFZmkBgspGOvf8sA8gI4TSQgP2Y/Lxx3oF4CAIoE
n18NiCM4mqWHouV3QHIK9LB7k7gJu3l4awrTabVEBUPeZW617soxoJgxB8aEjQ8J
/vu79UcMXKyNZtRUoIX4vkTxLCBe7HcsLWJuOPFQnZ6cVqecy8Y0bcae0qcEUbZ6
lKxrPXPZBsck2yOuOSPHxiBqAdlaynJBSapx+F2FjZHAffCqBkfe+FpIeLiHFyLW
nF/hSIT7CRvcnMsiXGR6wJYy2odBttr0t9As4vNshuzCtgpYbQ+eGAeFDqiSofIO
HceJvmPcl4t8PrmTM4JoOZlx0DH4h3aJwKI2jNcVe/tY/10FZjeh+KGWc3LPQnSn
Jq86GJXN0wBA5uWJqZZ8Y9aqviMOVVo5V4J4Crqfsx1TTuI9FVeQc7LsKrsasN4o
oUXmW2Z1NPos/qjN+hWCovu3vPBl/SCtboD3AOkbSdgPCxV2JAL4omgDtbgP1qRU
+ZPBtHoCPDc7X5I+F3grxAZW6hO73B/Ffg7gSfj8qNe3hYDPuVF3wGOxLMLryGn2
+YuplSALQpNnqCF98Pcfe3+xXLs71u5JP5tfmz7lOvw0u3HpZpnmJylS/tBSn3Ao
E8THBBupEU340Y8zYJTdUK/g7boNCxin9VmzFEkzCnQxGXQP7WJ8U6U0735jmoTJ
/c3XQztknxmETvYfhQKsdRnygVz9bn/qmvv5wZQNOq394EiSgE99cjA5uaetoRnL
cMJK3XUsNgM2HNSSiTXd38aNLETkutSGuazbUlMn5IR62LUGS5oMGGyMZqiBk+gM
EHw2QvKGlRvyDe9BL69vwtLu2Afi1BstBHo31lPNZQwDM6PAdpUV1eQRv/X9v2Nb
6LlX/GX+JyeXEjIvEBRVlVIh1psmISImrKk5xy96qevINYe647MhslJHl5lI9v7Y
mmbxrrB9DIxU/k2fNTJtMrZmbxOI+19nfotThppobIIvFo8y9sN/v16zx1KR4RpY
GqpZobxhuhUPWCPhWFMCyFE6D6tHt/YhX+sZNGL2dYzBQemNf2XgyNfAY/wLDyZ9
xU06tlRtE1DURgr3KNrhInPsOs+FnuHmmsyUZY3k52qiZdL96+OW2+aPkcp34Lsg
iWAqNwjpNN7bgpM+I4XDgxGM1/l5a+3kHrSBUXGyA3FXUE9HOkS3XJQTcvDrTPTC
FL+Nl3Dm6h6zFhPYMT/NAzPNeVjLRcPvTLuPwP9JgoM8TS19VXKeN2cT9NVEGd5z
yRCN8Po6ajKlJG+Umm5mPH6N/GjtEQV4dV5yMZnZSBcOdWb2UoIixK8Zr/JXSQzw
nUfpN9/oRMkKVLAX/gMqwoERy35oejtQpH0gO9PRJ9ofVlZdmJpzKSOgQG8OMu85
TK543qW16SWQgrReP4bS8MkVht3xbucUHT/4hnykPu9iRZ9BXAk5QqOLdh/6TKIx
oxPjIP5zVb2WwjJmN1WICIxPvW14F7QfM+lwmHFUBBCRk/XLAnsI8FutDosqgCuF
I5fg0r/KZed7/3KhEFxwd3Sin4fW1txSNYOdTjdwEU98KG7KrZcUe53h5q/XhpHR
iyu9RQNCi0p/K2tKN3Vnrbrj0a9qkRFRdFb094qLkfge9ae2oqRQAu0q+UGuUs6n
kD8rsKNjVLwVCs6sK0s8TyfTAK6UuOpw870SLQWSrNKRrtxscR8K7sPPvO/nn/Ap
rXigw6OwRldubK4rXHpgt8b04hdmtMsubRtx06QiPsdlGSKM+bIdhbCDngZ3+BQA
W5FrvtgeOJFtQMPuY7NE9/BH++N+DyNeo0eTHeLkUc9d2eZ1F+uRSYi4lFj0E2Qh
gScfOgoZJsW+IWMKJxOop35ydASEluMjfzTyfAgtFDeHpRYj2lwCkh+xd2fMeYO4
hjEVOG0rybwmaENxYnGor50RQBCVCaRkH+KQGuw30n4pw7rjWCKoKGMGMx73oKwa
qE0lh8pVkUgYcenvkYIXOAGli59myf+t+xsDr8vJ50l88MPOQAmZ9NEdQcEF3lLU
dOooijW1ciVNSxa+4h6pj9kbc0LnA+lf+7Lfwb4FodwGQPdvWZVOQUodHDu8FTSj
fNZymV5EqXzdiqafLYORiO6qfnRsB9dXuX2+ldWWPU3kru/Kl9R32pEszr1c4ML8
7nzf3lRzzVLE53c+DBwVwlWo4QadiugyIQzAN+WFcaetL3XUTxaiMkxm71PW6Dme
ispuNVJFi3et6e6nyxBXtvI1CTo+V1oLBv+SfmOgyM3aJllyEHCsyt6Q+E9cECDl
OSKwHuMMsLxZOdrEz/7EhBZMSi1STrKR7WLhY19gNCq4dJeQHaqLHRdoCqnc7Yha
QManPuAAFZVwZeUFWIwBvCs5K9BEhHJuJgLDXH5tKX/nQlEvRaH1XmY6UviDZRif
BJs+lnhFzeW9W3JwsvWE/TpLbOT67u/SiHgUk0a/oCfPuhzwU2Ug0OuD10AK3chr
sJIigcC2kYvfZsInDJrDdHt2Y3cbrWN3I2Xi03c74EjEk2EzbIqiJ5K4iy4kM6lT
lKxIDkA30uclb+rWzo9siJuH4PJc+YJuKyLLxN1kfQSedeciliCtisl5OuBGFL8k
nFWYFFnzu0BYcuATNSAplqYmPwwZ8CIaAMEndaiyvCFEqGrz9HREA97gV9GcS7yT
laPm6lQ4ofho4fbMW+ihIktE12GEiFviUecsC33c+VmquNyzZv/GBK9m20A0gdUa
twM6N8JoOnPdqLCmlODSedQRANfpL6hxXxvk8p9cQPxMxZWkiGPQcR6IXTlCBeul
lWUkJ7m80c1F3m261+sDBs2muAQR3JkKt3bXg/q83DK9ZkmfR9z8yKq/LqXO83cw
Du4nG6OtjliIofRgkct/awL21J5WK8yc7ConTQ6z4aRZO47tkp8f0G9c4mrhyAee
X1UqKMU/+dqmQRfom+I8yc05eNXLDieL+WCuy+qJQrjeK/DvKVp/TTLKbgotvo9Y
2Zp20IEQokeS/FDR10/TzdUo1pXu+w6xJ51SoKSktlbt0uVOUaU3Zi677FoXO8Zd
Czqtlaz4pKq7hse5DvNv9pjJQZX628/nTp9T9DW8VHXgIIg1lr9lHWbH4kPI20Bi
z/0yKRo/yMoUrq0LJpfwT2zNyuqiSfrDNC0uueqlEr24wQgjYKDkOq6CDlegit8Q
j+Ro2Tcy/nMcGLLwjYJyVek9jtEX1xAXbHu5Dq+fpZW0kTmJeR3zVF8iX2sFkJzP
EhnxKTMyjtiNncZxz0lZmegs4TuW7g8R0XQXNuBosuXo3twKznSAmEAXW1D2eAbF
ETmmGmTadaZCGMTvYjFK3lUT2HcsIPB29nABSnntfcMdSy10gsz21RzJe09V7ZFi
Ihc5PsG82zSDuc7vm4fDMBq7v/DVRYA5DSAVm1k1wR9wiHLLltc/5PVjelyA4ZZ+
rB5qKoHT6odISMv3ayYXmGyuOhwPCxkoUa0z5td/QzFHhj4JD7OGx6ZOyzbNmqtW
4TLv2oqozWv4zOvR23A1oa4ZL/wPnNbCnMINrdREE2mMNKLkiEKRt23+63yA00JN
mmVNVUAfacblknVM+BAdxuib/s4TBJ7+1d1W2ncnLqg2UIJWv8BySaPkNsqXdLWp
hfHiuQXlonpfR1GzXIzM5GhtzAZl1mWtbtKR7g2QVxJKA42oZ/+hkZdvHqEYYdTe
3k++8QeLokZwuVvlOpFCNzsAUehONNUA6onjqmTrAqwp7ExiXOrExmLqqoJrTRap
HNsNX71U9p49joY6/u4yOdCoTzkQTXr7gPsg7jMVMpTZmsyJ1/tKw4ncq+ls7e2u
VynRgKTX1pk3Kb2oAz+kyDki9WwY7RCvpL3IeV3GyVG0jVzSXV+Qc1CVHHyqK8Up
Hs/Ezasi75NZyhRkW0sl+N4SX+KMXtpGIiH41Ci+L01H5+aqkKfa/xpYvj6lGst/
R5KQKcloUPvFrxEy75Z8/4sMCJ6TYnNXEJ/jn1z0X3LXZH9KN6Ncp9pWkEvoEfC0
3PvTn2myZTVg+Fgp3aD5eNxiNgMJrdx75Qg0KCpogYlj0b6k/EElLrVGBoe/vUSx
gm82drL/cshw1jLffl6bSLRi3w3AzhM8ST7avh0H6T07Rxz6IkrMlL1YKLVj3hvL
1acFnt46zX20gsCobMlk2h9xh7jKKr/juySoUahRsKYlmMpaEnqL7F2uvEfmr3P2
j6XAwsY0OTUYRlFiijJKBVKhveHM22M1zkDw62GwcGDGr1uBxTh8q8vUWGl+uhjk
bb2YV+Ky0o8SPH/XO0jlBwdfSBWdpR62j2M1HxuyBEbE7H2VDhEwpKpY+yqtOuww
bPygz8Vk3FSD1fzenDfJYNrybcvw5ISLVCmrQvKy00X12vo0HpMsalYFRSMzcbor
iKv/CaA4FD+c8nxJhliKhRIQ5MxVD9CSvs/PIczbNM8cVhd3ymb1HAX0Haezi3to
1fT+IutUTHIDmSA03XTxqm6s3Lm+nCgM+DxF60LVxeTgr40Dwxjte9Mw+rpIjYFW
WhsoRwv88MXOuiQGoKgOnTTjsoH8cNjTTZsQWpuTytOtmsdS+eD/VuD7UWHzi7J4
zV7Xl9SJisFfQu5jMg4pIKylUg2dgkRMznyN0Guyq0dTBvB4Pdipz1RWThVPLVJT
hAMmMxh8RNC7xvxWWnZnrZsCoa/IEM0/vkWuIyv/GnWCHBhLFpk3THIxd4O5c9sr
lbABaUAd18m5DziJBmo3EgxEwMQb4ZmuBmv/SCK+O8DsEoX2v4vDfC2BBygA/23U
Iy7H+B7RDsfIE85XtpIoZOL1sxnkHtZH5Gu2+uxS9XZvY6pL07pA6Dd1fl/LJMWj
SQxrYhaJD7KKrfliT71Bs+BYeOGOw6vA083DIOKxUU6gXValFWAKn+X2jpxQYVkB
N3gULZ1j8KJY2Guok1Ehjoz9ny/fzZzWDtPC6aA7f/SEZJvzb1a85qx4O+og/GVK
5jO8fb6ZcLu6nfx9eVqJpR6HGRVBZ1JPR7Req1Du0XxDse9Tl1IZg4FpjZk5WSSh
BXhwcgx83PvmNV4PDNAVZgfbpzDE4yEzU+E8YAhONGYk82UXyOXrmWwLKb17E2OW
VGgYS+fZ/2yboB4Ym0Z45+IXlLePAuYdHFynM/v2YvdcuzcTTPHSNmIDBjsK+k0E
T6AXvLCiRLxjP0dXMg9eXyBj8g+6tB2KWDpG4mk5npy+5HxGc0w0BaZTJnQXYLBX
B9s8HAD6SUjs9nq0JYzBaX0EJdj7rKXisNJ/bfvl9Oq7RDl2Jh6MqXwkk0vb5RfZ
LmFoQn7rviWxAWHXs+7pGG/ZZoxoL4yqJoIzDgZibYqokcEivtbs8GSQDa+eM3jt
jeSgAiOuJky9U+p2NUZr4dI5m5XyiLeGmgzxxytTs+0ByRFw6HWHm0jfud2kx+qa
Gt0V9bDzG2tkhgJ/dasj/McTxqNSpEMXtv5WsNDSiprQOptohmbzzQ89UYrhKTyP
gv27lGPvXFXdgS4bJQVSdSvK0k/gGVrYmBQGZiY18WoZvx8ruGIscppu4yR38Zm0
kFeuU4qBAW6y3y5MQ/55FUc/ZwoJGMq0JbmPQ6JTtt1yTm+zAcIOJVmIHwqlBO+g
7ufWI7neVcX5gsASZXczBzWjsjwm8b4yE77g4fCgI0a9OWnDSW4a741BrqVU7REM
ocAn+xp+jIMrGsXE80kA79Blp2rALwXpGSibQ3uLyMjYt7Mhk5bzth/ZJco2knQb
gtNSKv2umEaKvu59WLfd1Q/eFuY028qlvBpGYtevVzFnLLpqyZZsx+WZzifOKoGk
xKMM8nHHQVUDTQ9l/Zbzjhv/jtlKOov9J2GxBorQjQrK9ufXxIKHVlGgLx/9xRf0
2SC72OoK2pwlWwUmK64pitGbsrH6ikgvi57xU+RoFuH6K4t/zqGxcASo/kIa2pwr
ppCfR2kST+X43aNpYmGRvB4yrrjFahYpllfj2+toZKDuYmJ3tJLLTWbllrSjg1Zt
b+looXd2Vxr2sKZAdhi+IllY+kwmI/8wk2ow7TnSzA3ButRanjzvqCEfC3KsUsO3
iFW0vpR8ENYBO1SP5IHAl1C3aPglu7qgAcI6olx+9oXUgTFXVytdj9BkYNElgNz+
J5bVpnb0CS4tzuxvFNupyApgFjjkgMidRYiKsHJ79jq9C2w3BbutBD3lsQvdiZvC
TBiFNZNLKktcxG599V4O0t2C6dr23oZfI0o0t26U6gdfV4DwmOcpRSB8QRhnTCEF
VCSFiaKSK6x6FveXe9fEdYVU1iuHGoexjNjQtemQEnS1uW/Gywj01suhmj+A8QWu
GQT+tRNThMwzJXJbSY6gDpxNmWtQePpK5AsUn2F+igGnpUV0iAFyHlaFQXilWaLb
Qq9zgsqSqDNifDHNLZjymrmT4OY0YnSCOUSHJFAj78GR8syoRQ11FQJrd/AiNpTc
WE1iE6pS/+flqh+kRTlxKWoI/hRoG8PFIj9navwtdZpsZML8HdZ2IfxoZ3Se9PL5
780CdNpDFFJgEU7GXRpkX5gd9QXxoQ/xuq804MLWSEL3ddq41CANvexbwSGh79+h
0n1k91W2b8odWdusgPYOYJq1Z+4E5oNQo0NkrS3dpCmMSr+DxExixnNz3gnwRBNc
4bJ0+ExFqH701p7+Qzv7lg132rt1Khba+Y6gRRHEKerCD4vw6UaHBvSS42FDMk8A
GmphVusrqUZhUPKMcDVzL4ObZ13+l/GQgPhRz3RFRerKkMojfOCvW3j5WaRNUcwI
St0vj9WUbnPnBQemeTc3s5DQUn98Y7ZNOFxk+SyK2ZU3TXF4KI08vDaEVaURqBAL
NlFPk3Pez4gUO9fwNR4TdOs7TRHJ7Zf8wSCM33UCO7sigl+wgCMlbOtNK37ZiRgo
oRKX1pl6R3JMtKrxW/17QtxMzq+FJL3uw83E3KBSu4uvTedEuQgbYUk18ThwAjBu
uvNaiYMypP1JzOkgnviHX3cpewhCEeXgy7rMfLbHn5E+jEK7KISPS55srUllZL+Q
V0Jn0G2C6K6yWVAu2Q/8MVpsbgtMyipcHivOZ0oq/oiqaBrQ2dmK6RgOIqW9P7Ra
E89sRCHeXIWpZGXx5OQJRw0ZaGS6ooQFAKqTy7938P+g4VXYoVlomUsqykMUhAQh
QV1l5Q/h5KoF9MnKm7jBWtW45zn7kVLBDbteqznr162EhVj5prEBEf/UKn3Af5ML
FczVCMe6K5FOblVoxqE/vVK3boze0JZWjIqSiGd1YK/fDUMVr6vLKcEIaHE1QGoe
9B2UwNpMXvZ487DM/d4dPcpoudijMQX4LU8Ob7NydPvVUGlRA9JzCc3qvcAKCUHg
IMZamhB8T7fsh2MItvFDosjPk1/eyoRgXio/pS75PmwApqzFH4ymPU9yMDszTKkN
k+eCd0UUgL+S1EVo25J/G/hLngKbu7mO4NhDkBnPsww5qq9App/vieFfGuJtkdHL
GuZyiZudVZbuQDViNYPZSGGFBsY8+UwHKXWeMLl7qIhnoKSPXggo3db7DBFsR0a2
3YR0+lrIerquvGFaMB+bz5RV5/XquIbAnbBJ4Joxs9As8aTSx1hPb7cPvkjubsa/
jThU7nuDOaZ3yH20aa165Mf4o75zNOM9Gg7IheZg0jfC4yBoR4HWZuFM1KwdjDGU
D3zpVr5LUMBxrAZplHwxthUXn0oY0MnpEKIXjIhsLlKEezohPIh9K6t88F6kqsyE
YcLd1Og23yQux0C2XqdjTtrVcEGvAc0suJIhBq6F+UtYwZNNmVwTiYPIvsam6jQQ
TKtUcxSbpdhgU3zOfH4f/4tskPM69KTeXGchh9F5QLudF/P3b13k2lxOnqq/CpXJ
pVXCckI1yYiFUK+EAzYGdYgXgd4Oo8LBZDqLMU10RUg8YK3hgAL6uXfh1SwoYBh5
9FtpduD31OFHO96LxtFsfyqydRdq3qUt7XSSdagn+uY4V1C4fmmopkV/YFv8vZ7v
gTwBQ6d/NsVPSPwwHQrNB61O99RCYPtkPz7xSOEmt10nl6kpTk1NLIFfoMomxuGo
rvBXjGdQeuQL0nuD1cTVZQxnBDAmTR+MKkHzQKAY1Q98cCfPGyzxDx1gVR+pK7am
N47eLuX7w7xEtOHidi4PWpqx7UV+BkAsRWF5XGS0nBT348LJl1ZMZ0v68sC7V+wq
zkypMbL/8dO1Rmens2attswE0f38zqYAoxVpCJrBEvkE8TmsnMaBV0ozbPRUkkAo
ntgSRkzV2xcgNrJSabaYtSMDMlgSKiT2hgC584iQly6YiRTwRzrDjfEWPe/kzFq+
1wURWMKgbkEdDyzcZC8TrbZvzhDQbppVEZooU0WVr3ZrjidXrqZJJW1CagwTwekU
0F9vlVGun44nJIMVYA0xe4otD1TQFFukW719IJ67vjgUJBP4J/DnexhBgGLrfoUq
a0qCensPa8LmIFVPYVmnR5gViKpvT2C0SG912UM/7lSNxalyA/TEyrn5xB82At/H
n5FelZHgYP0TwLDU0LghMgdgv6eoFhfMb6cr8Cnm06zaoluHAehRdSUvVgfwAOhQ
fi5v6QkJLmOQ9WY5QXsEsT+hfzkzeDY1Ui5yHIJO3axtPn5eJSoHdfNvkt9hGncW
gtpCzqC/PXlZGt7lRY2hS53jHD80TepaunhPGM6a9mI47a9jZshro2VMfj1K4VBl
nJriyOAlLLnPbOgfjlPuHnbRexkjzCX5Xy3rM3wgjBY75tFnHpHJ5XuponZjbwdc
sANUxT6yQX6mt29smdSmQElu51FPH3KBTUTerFyqvuDk0vT3cwZx/iCRRBZ7Zf0x
+RISarF7Mt0XvWDCnyqygss4nSCtAYOCmejSCqWOc58px7+zMc7F+iffdvJeptZD
i8Va4lqRScZqyDMA70sSJK8B8KtbB40yVP/Te1fAlql+Au6NumeAiwpzJaYZrHiy
iIQCsmK3jmvBzxgSXEJyyt2RVaOw/vcUwn+QVoL+8p2LF6EN2/zTrmm/eD8qVXBI
aj/OnS5KFni9HmzA5CaCLbh5JTNFmN/bDkyBpArh9B+VjtjkwIsGXsEIBkLa6e9D
TvmVpbGWbLgQ5eRTxplFDkBu98GnFRyriKM6DyLhQyQE61hIKi3rfKPf2vkwPPa1
OzoHSbcun1DmqACg7Td7e15A2ccBJ3F6FRwVyzmHszpEjSP7mTr4SjOtU59RT41G
e43VcL0QiYU4VfoOSsRujxP75QecO3ValkL5CroHTuSm4avWcSSNapCSryFTe1HQ
0EPKXFkEvmAgz6ObTq5w4sNXTTG7AN8C3o2tfCpwzEIt21I8t2URM2jHeVYr8rDc
feFipoLZYzs/e2RIXcxoisuaAz9E6c4MpNPXO0R2SkWGSc1HeReLdMET5FfOqZSy
2fEEG2erJtOecH98BY5bCea2VDuYbr9Z6ycdvByWm9ET0TxYz/pFAiW1QJGx7gKS
/75LQHwDKVsxvcR4SpOzE6GAdsNp7OJoUCHz1tpt6QQLlDWpbISC4QnrBeM8ympD
eVNUfQIMqWNwuSGjz8rZ090US0T+N8ElsXcVbG1dlL5MvpziV3IDvuL1jWMak2Qb
BYKm6602XFT2txflQG0h5oOAvBDuRom5IJNhwsmm1DnPAefVmRJ6O4kB2nXrwCB+
x7HHqLQDStyy940HRvEEO9p7KJqQK9pqbsvCujkan66md0JI4c3vlZEQrSW98mHO
FSmAVV27M5LxzUiOA5Z1Ujl27cqL5Z2pVEXYoPZxPyClx/zxabyKabOOtO63KrXd
NudrqBVc2qfnESzrAtbT7Y7OhnZdAiMZy5KlsHnfRZYH5dqH4W0mzxBk+5O/rsLQ
qZCjCIlZxIVktlE+IfmhoHKDuKyprDp6STifeYTA78BPIDk7GxPPrjLh2+LhOKtX
Qz5Q0G1CC4kC/dl5MOcEfH0tduW0KHo7krHjiEhFTLDmc8WhF6kkjv9k/48jXG7N
2xZmAWcYt8Lrj4btXUF0ossdZUqugUe8yv9k+q8UzZOJK0bbgQ09b2xoKwQ94Rr9
Q7B2BGHDIaVug40ebTdKfstRMiccoC6xVe3OhpgiwDmYpByAIUgUA/T6FRMVPCcZ
qrKkjtpaMnqu1xA5FNv2TMi/GC0rXQ8tpKh83MxKKueKJcMo3JbJ/tsaW6j6IcPN
GU+WDvCc8gafA/WAL5phHrpXiEXhaNRYBJhtilUNCm3/kCfCCQlfDFfEItphcj87
Cf+Vo+Bx3/7Ux/bU8xOi8fbcqR9BeehEtHJJ8ZcTbh1ALvk9SFAVtYxl2nXIXOfQ
EZ3HRHqUqKAWCeYpYqWwjUbzM+P8hMzRolpQLn+vfdmk4OM1byZPdUvDv/7G3HOJ
E0W16XhstDS8i5qezuITF6wsbW4G6Q5RNNnUr+d9CPfmhfOw4/lbrKl2rR/J7bsW
XjRG8ajdsksHKAdpvQ1Wg11/jk9/PMWJjp/1+JptydClsNK6upkVcttoJV9QPkgt
xLnODq56WayABFp4qauRGkqIAcuOnrOt6M8w4zFlUwCmusZWicM45/plEagbqIaI
JCq9Zjwv0CwqeciGjDBoy0Awkv5mxAPMGXPanoq7BBufkLFlnWxKQLJC6+2k7o6Y
MCC5qP0SLCFOVoIakfiwXO1lXbQYJ/4ees+l1POWlJT/7Gjuqaig4Vr4iyNLumfr
7FVlwb17eBIGMgySkisLkkH2NWnGaiDrurrsKLrBrWEjDf393oO98X2esJTgNIhw
ltFNp1PAw85DMltA6jozjuF8QHH/huSe+jB3b5/VcGVbk/DiSuqkut93NFaWleeN
2/VdqEJKvLkVycLzTUOAIncODfwNBm2QAtx9AInqoSvjrLsL0w7xR+CUaZu348Fw
JKmbRVMB1R8PkjVW7eAWHVdnZjgNnLR28V5TC2x5N9aAlci3FkUqyW67FXO5FEeB
OKP0qAOjqqKx+HfGz85rucCA6Xt6F3C7h57Qejuk88JrUsYSr+ledV0UlJl94QEF
TMmKHTAByg20zPijSeoCLppGF+beHHKXUbzglUzPvJ9x3BafFTd4lTYGLpWYzE0P
yWhkmK4gXZkAlkkb6rTpeceL3BR1MNFZK8dXqbo1sJ8XK+C6rdBziBxPIHdfq47J
xEk1r+WR2zLOtj6Mevf61EXkrI9W8qyi3//syw/yV9MCiUHj22GC7rHcQtfWM+Yu
COUfVbsG8CzzJXVBFGrQywzQcp9yvlLX+WJE7IVBJ13BCrzGhsju03Kh34YbS6k6
chg55VxKxzhCODa6q1XhjFG74Jxh0ruS1JZvkXTZviSMDMncVohoGlu81MRH+ZYi
fAhx6g5uOJFmG60vogSufQEHVmQYryww5I1nfQpdakSqz4ncGipNzUtl1LK4KReB
JZax6BpmQEM0ePfuLtCNkRhm09j3BCHPDnBiwfgEZofwHeL56+S6IRrDLH33ojGn
JzB7KuG+Zbs5RsOTCQ9OIPy8KWICXnzXa8xGi9DhpyY39+yfl+/xFjycLYu54uac
eIUEzMTDUqKoku3tIG/rD5mKHLnP1wlOKA3MqyHqgm4S//ee3PWPJpOUMRk96hz3
xrjCdz5So17Zgl6u3QecpK6BRgOey+ofoxulBV3749GHEnvVJdKCAUu/j4T4ZxoF
uL1I0KzGbjv4Xe6oDMg8jW86HMxZSRLDJ6x1pcKfTTOplxoQnv59wSfSktRCaPYs
8k46HO8cj7m38rZVeoMckm+JYzraOt8qb4jTeYAd9WE9TBfzqv5iEZFhGQ8Ha+BF
fk3OR70THMmOh3AOWrP5XUCaQyzApdWN/Z1rz5mVEV6gpHN4nW9jxVISWGHZswAk
pEO3Rq8Zu3jsyTMavir3ZHIEptZOdpcnckPqsiSd0iCpuoynYCvfQ8CeH7f/eSsz
1UkD2qf0Buj4EofuKpn4ydMS1uC2+NkOgS3hOP+FtErEmMmEdK0AK5vI4DWKG0lB
VRLjG3nKRwqluxh6JHKJAhUUKxuxGF9gEQNw1qx50KoclVE8zxlC6xafxMdLYd7C
YyMr062mrwiQ2kVsyxoc65ksginC0gvdZvICcq3qJvX0yUgL+jULoI2KCiFQO8NB
8xfUXTkk1FjOISsL9eBC3QCPzGFjzP6kBv6v3ebob5Gxsn9QemwfuXzcAQV749cx
+TKNQ7HzEn48hN2bvL8w9WPbS05XwOXoUJJZs5c7j3jyQNZxJp8wRkmGJE/D2wy1
/mB5/gapSEZGh4M+R4vpG5dYlPib+tkbxgPTIJ9xoMIP6V/O6MOMFmgT1Cd1wHSj
8axwEZ/Mo5KqkfNQ0nze2SOBzBZI0cgcYcSQ0emXkgY5SK57t6C9rhISRB5P37G8
0+V5pHGM2JrDNzgrrYJMMteeREkywemB31+as/NgO07Y6txLAr8h636b1ASUHFj0
trFwP9GODMI/8JESeTjLxSuQKTECqmOXWH9mCSQAaGeTGtVlo6RonX6A9iJQQB28
S3EnA25rfAO2jawDLm9l04CsWf3l8uTLroCw8/j1TcYpGgzZlqTzSGCoQtuIizAC
20f/ihP9tnKkC7ytFPggFnvrHBlZVpR1FlOqLVxgMHPRRdDIKQY61h/pb5nBcUeL
YNun5JAEPw32tnCipEM8rxXmLEdiIIFgc1JD9tfquGaV3wF/RDrWp4WaJIbpSDHr
oV5n/2uAPy+6ERIn8TlkKdG5wqBhquvZMqe6YtVZy8OjuJMtMdohSkbKiqkvDzPR
xvrSatPEzGEnGwswidc7kZmOgwRjUqgKUUur9nD47AIoIFFgk01oISwcutUhE1kD
kafN2KpLDHpg1NPx9WxRyv/U8K029hbsEYXMYZpJCthHxoVzUXjaxLTEyC5BkT+2
N/9ysCfEJdWZLhvN6MGqtdveJMrHxF1JaJOR/DMXF/AccKMutSXubLs/ZRGZY9dn
Mk3asL5KkfBhzYg3M8Tv5CozKEGaRwW6GClKMnEx21H3kL77DtNzG5MoUH7NxwLd
vyJdTrBEA7TD1iNKAYuz1Byxy19FArVZ8vRTZ1LGRJyOXfp1/FgzCy+in7z5jjEr
Vyym27u60DldzAOvjhSo7ASQ1UAa3BpfhBzxpvqJhqruL9lz+DoqS/lnRHqekxIb
t9YY1Owt+W9KQ3i5mtFADvnI9IsgMC6Wc3fqPeroZjHs07wWyXNNvGxOdlggH2ZH
pvVa3xweUvroM9muaC5YllU0qVeDpGOSIl2krRIQIeD6Rbg93EHbynwdlBJbQ+CB
WH2nljmB2y/2VS7FoHpZMjsm8pUQr25ufP5iOoxXzYBtv5E5Wo5oZSDIsRyM9Exm
1lb1JvHG33oitVCWfphn75hjBXpKPP2bfraaNn/8qPcG/HR+IBqMZhAXIJWe2Kro
/olJMMSnhD+pmc6dV2IJnqX7723+slMdxxiEgxZJnXdCHl+2ayBucMgtNA3hTNJ3
rx77tZS9Wfxz2dwCta/cofQRZJM+EpsEbhCT4iGxfBdttdZGQzUxhZxFixwPLumA
JuTYZFxZXuqcPCfAD1/u7GZYkfBoVKXO2HRDRkotZgP8UpknMrDOTnO+59pNhjU7
0ztx2clRFcLHYxyDGThmWf2QPtciu8mVcgbIi37dQukBNoxPZqu7Gp9/eRWpJLqO
+3L3kBsx1uqyv7wyfI6rYkFhkV0v7QP7x9qd4CJr1HQXL3IompdPjHRzmkn9BGkt
xmFsaENCv2WY9Y667G84GjFHGksQ0nzu7kA6l4dad4A/96zOb+/sAdRnLeGP3MXx
ykS0oXTdyZ3SXaBUQdxKTggFL0nV0U16QZLiB1tthCdXjj9+2H1lRDN9dpgkcJ7z
nZRA7kXKMRYNjTSxrjdrrrh2mdvKyxbHrAIUHivOx295U4C+zCeBW3m+KLMLJlto
2CeGkgEg3eih4p1KcedgT2+yx3WxbePMK6larlgZDwIts71zo3fL/Hf9fSEZ+1fv
WbQ/P9OEVrwO30vmdBZRTge+tEcW1e/1vw8VTR9tTkIAyBR4r0k1vNODa8j5yCZ9
Fpqnz08eqjHF9G4UF9azksPvkKysciEgSDvocWe59wsvqTNbVvBRLnEQQVL08EQV
yMoaP6MAyN7nRKO38HmrEJGRJB41z+/FAFoAnW/k3JAF1gLrSerXyWzKhCJbcjUQ
DlVhNDWkEyzaAvRzLDiSJ2j+YaXU+vsYOGkIUvC3yDJNaZg0oqGyonk/5Hv1Vu0K
LjTCTkCU5y2t2nGDaPyh9HWd/hjYqkeTrTasZOTGh2OrKFzLrqJsaR2n3311vAfw
QKbdM0+hHDP8ATd/HblPS5M1dXf9mSp+cHdDtqyEY+BWyXxDCLQHPI7yECxb/qT7
mLu8ICdf4BocpysDyueF5aMvJSkjGo94Q5GV4Rc19aaO/Laa2uKugM+Z1w4IW0kV
/9+Cw1Wj2MdDWWEqDBc0DeeqVA0Nr9LaMQ+LSBWxTb3Dd+OGUlSwcL4YNNdZW1/y
u97BhI8d0LvcCSr6w94T3YVLwsCElloh01mpvCPb0u+mm0QkLt6fr2gjRjVutm1s
AxwExdd4hAAUpFXjvx8xuoFV8+u+n7uhy6Ma/tj2PGaciVN7CD86Y7hbpT6sgyFh
GCyJQ7NwEMsjKq4sv3qKjOfHDWLy9WKLXtuonLxH56/sXLlEytUBftOAaaLRBlhB
3b3AuvDKTrlptumfIy2GUGYH0SNEQBvx5SCM/WZwV2/uiE30v7UAnWpVaf4zE0lh
hUROBDlQEtGHgigNoqF81mwlj5fgOv9RGBXobeW0RBdRYdTUTKoHf+EIbxc7s2jS
TSosIlzeQYAXOTYkJNnl2ioJm4d52zIhSbs+YcQLqtN5U/rhus/GpYzv/tOLnbDR
hUsqXyOnwKZB+qEawgyLboy9+Z7IzUbYbI9ywgeM80v5lMJlic65pz1RfMUMsolP
0qriuiijQh6G3qag1dT3a/U2wpGoYu96SEb+6G4kFJmlWCIavdbEI1UDnCch1MFg
f0kacoH4Xm2e65aA720uTRwnnrcESAsYpuSIis/givCQxsHAAICyu7SM4eE1sp2H
BVnmyAz9EAVIrOtXsnXXPvjvgfKV3/olVY6TZ03xua41/yxq+E6GSJspPlKMRmM0
0yQXdtAkzvjZfn69EurZ/pyHvB8iI9SfkS69aLi+Xo/HcP1xQW0lMu5hBRinhGfZ
KOaYxULUt9b3W0MWg2/hHPaHJhKx4zOaeml1UaGL4NVKA0tn1rOddZUUXwScIqws
rAUskJgTzXhMtMlz9gPGk5bcudjd4XZBLTf9ft3+leqO83SwWDbEnj+FLaLiyCm1
317bEWmIZK4ChCyVOethMH1QZsComlkoo/cF3c3klCC00UKY4tew8VunXf9ky67x
yUb8XyTE1fCsfe3ro9DXvryJZD9L8Zk0GiNI03gmsYYyb+kptookGWCAvgye93kN
u921t3glv5YGL1dqIXwymjmta6cYZfnSdxxziEJy4krWtlwuK0qtkqXZG3a7VVF5
yfTG9K4Fm2tJufDtHSKj15YGar2KAZECApL1cT60bkFJPjjnhlaU6OKj7ZKtrj1a
ZbToS4DH8D32L1APltimsku02Cxp/eNe5rsg5P2iPa7wK/xC8fCqVUi7+rs1vXdT
v3Bl9wptN+14ymHBDBNPkX/HGPxcvcw5osoS3bBT9+eztIeboMw++Mj1wGuQc+Yx
qA4dGAOpeSCdsZ1Lo5+ICwftNo6WVg3xAGDWluqur/RqFzGr2AbFQhp3BvUC9iyj
RSasYUiCsz3RFmCCqBE97CEjbVNlQWUtJMHApFq7VvdER4tPQn5zuWTfOy+5ZaG8
4abTOb35AJS/hRxt90XKAm0JYXpmKWjAcM70GdOn1EYabDJzyy5z8gkwUehCE7/V
FUyIwd5KSQBdCUogjr5sqQggPHvrzsUBDmodCUx8PprXVAY+XXDTI/8pCZGH6Sg0
0lZf7lUJWKuFF3Z1d6x85bozD5nkLrSSrhb63V9fI7wBBVYiKqaXfrDwIsyWByGx
md+i73LQ1ahBFbGYNPKSgGyQ43FVwid7K/u2rd6NCXRgRi8o/moth5lEQ6nGD8je
zB44x9zX+y1sqorHc3+xoO6UVK+4t81srlljX9Whgs7kRVvkPxRZvxX4QCz9qz6U
RWr9UHnNIziz+hnvuSykcGZ3ntu0s90vbAGgewjlFGfvP9QY3O1lJyAf2JA/K7ct
A28F2E1g5Pv8ZR4WhApNzgQRUL+yPo2uO0gvph/8Ns9dIL5JwKywBz1sb6mws1aF
ftfI7CdW3nW/iZdeHvk+2iw7eEYA2ZRE/qEun5qQXVca86F10oXro9+sndLxuuwn
DHa1Gv7bIdM9FYQLxRnQmfZW2xQiKd5V/loRc0V1H4dZaZvhelBk1dii437Pfy+E
IzQD2Zb+m8JpFzNimTz4xmz3teXCyAe2/eGb1Lm15jK24+COCPPIXUJinTsorR+7
iaPMAvhhsroNTze6DuXwppzG4b/VlEQfj/TJKSfpuowVt97S8Um/wfnX5jc+dvBx
rl8q5z+N6oeIKP0hFANBcOZxezc75ed45JfTyoEwv9N0LHsBJ+HDEXG2ES8TO3oY
yR5Vo1fFiCWR3SfbU8R4/kjcmt4kQQdLkYKLXLHyU4yXEnsUxLkXGN9DPFGYIfNX
FFaYS0r6k75iQpqQt1j+Q3RBLZdUIqm/R709FJuuHi8Mqh6F8OoTgmYyAMFD53oV
jcpFC1tkJqr2U1fZbbx+ftUxWHdQC2wG1xe43p1ciNT1KHJLS795YO2bpLp93PXB
o1TOnkPdIpzmodXW0aXtXud6dzSIaQctdzC2zjBnK1IH3YjC/1M2my6EnmEDGjaq
PjR78BVI0dY8mHoErhYBlkXxKNJ1c6YgaeTav9ulJplP20Hc2Snv34a/Gc+jhNEK
5MhPScAgrdaL9bApw/aS4TnTCQ8stwSO4FyeUmq8KlC3zkDEkNF2JCeDgNCjSBTv
NDOaXgVQe7yAH4FELGJIY0dbJIx6V0k3m0ZznvzJSXQ74D5dQwQEoSwtLY43NQ3t
sCyPbxHnXR/grqVS5mmIj9D82x9dbJhaeDWTIhdUioy0WO3V4UCBvV328E4xD2y7
v7ShOA+UkbKITcEpSSQ/IbuliY+M4RRFyJ3uKND+sHyBFmwo8dCTEl1MQmOzthbH
WmL7nel7TCwe6uP2uHFpsuKx6/UxLejgwht3QVVqcFwxslBVJpd95ZY/pG1mlNNX
vmWxzvoXDOKm7jAAVwg1Evve8N0ZFF82/fKhdSQ4g3Bg357T7sY2RaggvrBtxSQd
EKLug7p9AVVvxSpn7CMKVDfNZBuNtbLrjmYfgXMjNTUsMy+aIwKgzxLZXQ071Ln5
WYAcJmla9g/GqhaFD+i7hghBCzKvphXO2BJ1/0lToXz2qM1mXYBBaNSo8JMGWT3K
dDowjyPqCssBP/+Wq+YWnSUQKoE83UQb6FG++kLUerxS+Pq0EzmDc4vQPyiEMKEY
UkEhKyI82jtlyxSdcFLmnkmZLcjn9TrxkCX3WQLp3T+diRxWnBP0n5VxG6nNc/sn
nXvSVO/0epuulD4qrj24MFKUnTAlb7mxAYBOQTFYR8njDFm2ibZB2mhP8q/zsaLu
1iE0EEjcQG3AoEUQHUdq8ssD/YzvXeW3ZlbWpgI2fcfvHbhykjZAbZSzDQQos7e8
Kly8t1aThQU6y4bWoaXCmHSxdZwhiex5wBV4H0OKEOkMr58VFTaNN+PRuoS2Uh8H
ZISrOxW90yFnE23/YFv93oSyqOJNCJ+BEPhIaDDiJWXISm2RWtCYFy0iUeNkgovd
awjhgtArKN6r5pR7wHXCfndPwJmKsrttE40/fXdNvtvz5MA1t3RDU0ZiZ6IyuDeA
kOaxuFEg8LyxpysTAlNwWS54pB0oVqA6J6lC/GVSaOO//jTeHREIj4lIbq+5eM5y
QYKhewpt3BaZHEZB/6Zqa0lWU9Q1TglyMLF74kgTlAP5I4V9txoFxWDuVxRkTAeR
5A9KAR6R0OgtZHonxkGkyv1HzIp8W7Kbt3L3yRoXLx4wjXAh5pMFTYMO2Htdyc2Y
4ZulTzkF3F4vL/XDbiVDtgJq0W3fPgWVKQf4gj11dMpC52awGOGljLryB3xSr0eZ
tDRfTj85jzt2+cAJ0fCTwreEENd08635Y0z0SPmYLs+s5AxCHeQ6jqqtI53ysksv
xIHqyS67TzsWKWVOd7atnXl2LvdCib0rIk0eo+IfEVdemf5E6g4jp+B3kQlTBooE
Xm8yqDWuxBnSubBYL6PfKPTmp8gB6VkPCTmp+H26m+fIlHpCUN+ZMZLymYuwqE/k
2o7iojhLQYVfHVcLx5hZ9KOjS72vuwlPWhGq9aX4IoFNZq7Xhnv/L0lnYC3OiZFH
n9mBlgJ2+UKxEsZ21YSjUrxRB6LEZc4Ap4dj80ZbyRzwbhjMDTVonJX7oO7Y8+Ra
YaORKx8t+6PYjAxTTrwhuf8Xt6ddzCQ+scHdQAzbEt5x8sUz3NGze00gbZyYUFvp
QGCUxoMxz4Xx6Nh7lg2YcPntjeyRBd+aix+20ui2viCzaBqs65QWkWwIwl5Ehvix
xCRwIylx1wu6xQLMrNZKccKw6sdoV+lqIbmH5JWULX+zA53QQ6bnU20Y4t3b0qAY
MumknmUO9luyCzV/Qk1TtdntdnBzWNWGyPRBh3MRyEMCtVqFm9ETVr6aKnT6mQ4h
CteGj//i59SJEYhkpw+8mlp6AlPX703sj+g/gT9dQg4pcoldfMweKCrSlNMV4prB
2GtInvGB09lfnWdVxOZrvZ+jrBhMbbJFNoUri4F3/M2vml+UFRb7kl1LHYdKFoK0
x/KdrlNr3VQcnaSRLpAIkPa5S1T3qD6NZiLVx35YmtL7IxFXGI3ds3eAvGjj/Rcg
G1zFd/KKJtzmPDNJW3kJzyIYePPGmNgN1HAWlsEvpqlksijtwy3aXhw9FwPqCWqp
OEo00NkdxQHUWHW9a/6iv4pFV0l1VWfYz99BtF/RrZ7KXj5abFKsYNx8pPxc53pA
h1Mnm64/k8zFEre2UfP3OyXCTQYY0DIDI4UDHwmWrwPUBUMQG/8krgMOM4ZPebUT
NI+7SvweBGq7EC7fY/6ncfCjStrj+TJPtoiw+SBksWzaGc5fl7Hp9xd9eqhBzFNs
QazbNKChCGtN4if6KTTr/5RL6U6DGzOYNCdsYLMq/Hp04SWK2hOn5gNklH0/MY6r
zMV/6EeRGEe1VUHBFAZCR7sZXXRe2/nFa51PTYdVeIeJyIvh/Ohc3dqJSU+lntpl
JshE69cDh+lhzImdhnwyHr9UnNMtelYPiq4RLWm7H8ZD88IdIibxgdZy4oSmY7gJ
pbrXV+zwBxvFIUiwMiZ8YZKvs9jrJId5z1DIH/et4dZs18d0FZ4csCAtd4xuUt8d
CJQod415sF8OPF8JQbQW6Vg8jNellVkdgPm/YnX9eMlPa+iKCvhVWm/eoB9bLO4r
m9UX/5js29DpGLXri3HfmgOXke+nJS3LT05TwXJIuqoVHYkgbwK5/GcMOrf/vXiq
GtYjAmF09zEXs48+TXPdWrbfMiEvpQBtrCGMGK9Pha6JBGIDRR/jtSjCTqZYldXg
EhfdAy1PVC6ojIbj3dJpmI2QklfDpD7atQu8SZcW8Y2g4TSRe/OooCxrHbKZeFIL
PI3TdV2Sbb7R6tECqn6M0MlXT1uMKKcfBIVNx7gS8Bqawr87bbK2t92qRn0b6ty4
EUP334R6YPWl7G9QhPTPAbkzNOgm3abkmfpQ3y6ZG9rmEWFrmBdwVjqCW7ij5WAf
Gz86Az6lLb4OGmYYv9sI/LBKp7ye96S2joDGBFoYLW7UmNi3A+8VrkCdi7jwpVYV
+0Xm7dbWfuKMmxOxGx230d34CdNbE5qyf4WkWImKNmBD/lMhIJ72yiG197K4b1jy
tTRlMe6tbX6XE7Od5i6MRA+Tyrj1JHzciIVJ0bBFcpykq6ao+0XDSioylKPV5dRB
7vtSfnbW/FqVCvsass4AOt04kV1+un9/jROmhrdpxDbIE8awxsR508s3R8IbKk6y
5grIexsFQvZQxF3Ri2RJ0kHKXMSq4Q7GqBH0g3HNQpiFGYDBQUWv1BYCnPh5GOmC
pOj3F9a4xFxxr3LRt4/1XfQHuI9dOO6S21JyUajMwfvPppVsjR+4LggOzcpJNW5i
x6K6ROcVkdGzZL/FxXhWj+nigA6nJWhE1gbWRzpKwmSIRPe8V8YQmFquhh31QgeD
wiaJ1lJ0VWSyr8D2CZT+NqxLMzYCzqIDG4TCx/V41ruTNGKC37Aq8EBWfl7VxCzc
6uql78m7DF6loIJ6rikheeCacaErvdQdwmebnX6mnX6BHOtmvanO98lsgGroJRBY
1+vw5PonHkFqxiS5A003xDvKkcxxCI88V06BqJ9r1IBdpUJljX3MaCMIgue8GAHJ
bn1ymiF4RdSpRRFu/H8pwAbu601YN/tQocgWGDag8COsc4twgb6BX+stQTioE7ee
w0vwz8K9dH3j7ZK3N+4l8BkHU4E8kxzQPuuIsWn37mmcZCZFlfNXf6DBnp5PvNcR
f3jwMc+1t1EWLOyG6tiWnG5NiJK0lEYL5U9rByglZIy779udGUAWTFFbSjUUAV8x
ziY12f8JVxlVujU61XGXQGEAZ9afZHn23Uy+Tq26j/DNlxK/mBLcmf5yw+vRT7qY
O16xfM65n9sux7G6pmE2LlSBsoLDArkfRDB8C7vaTHtdCuIsQZ/7d+5YGwmsb84f
qXniHZNPBRt+FEcwQGV3xqpTcbJTd1MjgZCyi0NY7jaO2s3KkWuf+iVZIXxXNfou
tumWmOQrZbjiPvytkzFu7WlrV34aXCYd0wUvfUBbg2Ku90jikomLihbm9GtNgbS8
dGdcWdTZHiKs6/LD3yw3xUVFjvkmEjgqg+XEPFDrbBPtpOeq0hJR9ZZitSdFRUNs
LHp6+DQArPj2ICi2IHvQKI9rfFpw5i4Svymu5LDsIZILXxwiD1s3xmYfcSvA6DuU
Q71FSXfD65g2/83OAy/Ryse1tERYjnUSy2Q4s6qUwUDCYQskexn/ZtjMyYPhQZBA
eAUzvWj+mORuCl2Bv9emb1/B2l0rrKabQpB8gKxesWxWfb4kcY5c+0fLD5E50Ld+
egifKMUzCgHGuLXeh8NbgIB0iyRzjLjfCRgNg6UCcspcPs0Cf1mY2eAZiaVEQUtj
pu4teM1DtwhYDwonbgDnQYm+PPm77JsAXj4yEvcpaBTahgMbjGmlyayVakoPSfYJ
CbrHb7+9LUbDsZyylZZA7YYfJISQGvykmpEvUqnQgMZLF3tvQh4TL7l1tN9ffv8j
NyIrRuUXWeHdUL0UHMLRNe3tUOmxG5cvUnRSERf81MXMP1fIj9BxLzcMeUWQUcwX
yz31zaPcinOWj0m4M4JI2skhixbewVczt3J7TP7hQfHizFfY1w5lMmuwFFMKq/hM
S7YoGtbtz5LebF3a1lZ+/KFv3Y3/2YEL5HLNg0FMzyBqC+RsYpjsFrAMYmk9aAFq
VhOg8o2nq4HTPM1MdSnAKdz/3Qo3HYtq89o8Zzv/v0/nvKjzLt4NP5bZ9H9ON/ZI
M7ccxoLydRxIdKmQBlJPLv2EIy8jnVwrUMPR7Vop6Xc4Axwu+1BzVB/EGeWl/LhJ
+rC5uMSUYqELx+PSOnezVuq8zAS6Gi4ZyGlQKMgxb3+pYnM2zsq8aMAukmi7bOCm
/QNlStQS26bO1jrRH5pugt7K0WRnG37qGurm8JP9cX4Ub3DW3M7KOviWVljJsPG6
M7h0lWBrRw40Fkn+f0Fob/RvK8A3M5/nUiCVR5IDE4L42oKSc4YBrmG/tTOqXbjY
sXsg5s7TGCHYIW1p0mA8EoSKzueFF4ywVfKzzY/74jnDRIwK+pUzyybjLXooE/dG
swTpuE4eXs4MR1H6mJ/8S3cQbRuG5ywtw6xklNAPu+uPgMbDvwc4UgjWn/bcGsDA
NhvNopKPITUBB2jLUrI4ChBhLqq9ssbADoDuhhDK8ZfQ+9nWiCTfXkiksOMPwjcV
Qaecrw4UyDT2ukEWcqYBvQm4alyGnFXu6KEVm3A+G0LSPFUvVBLGHAD3qIxGwZGt
8zJHsi2gYo9ftNwTuQ8i6ymxl4skgycKzCFaSKryikAl4TWP3FOSb5ul+eOae79D
6EJQhTxNtGkgZCwJtMRvrhJ9mqcT/ZLl/SQPLc2ZEVrFvxwFLDSmFPHbrzPz7bhU
9hhZlni0V75vYhQiv4j7Qb0SjXH5+8jE6zIgvW3jWJW9nk2BU1truYcykSS1PaQv
ciHAXjS309dVihzCGUhMmpt3kDtlZLleLpXe+s8vCwmbhgwHuccsFmlaVMm4OQJk
KjxnBLUULob9qC3ql8ZMbjoSWX0sTMFl6u4sS0UgmK01FV+/ZwMz3MongKeMpEmu
UxF9uG5U27bF2l/CpjJPEGIMFm812pTYEe7hKUzRRprAEtlgHERBUqq3E5x8zVZ+
yTQJJkur0iwyHQwjrBHa4MAaXb26boPaacqI86TMdZvlDI3g62TjVnKOItKZedOS
GgSz/HZApJNqShsopIGNghcjrQVC4YzTJen+0d1GBfeJlY/NwZHx5iIJ7p4+d5VT
yxJhSn1+Xb9vZgiUEFzw08H1w2OKhFIbEKTSGcksk8l7Buyx01aEq7q7r0xoocen
H5xreOou1X3oHxP3ISjadUvSLKOFREXVlwaxWnOrI6PTaTgODBqzLEk6P64d+4Or
JSs/TAYNmzhgHzkDcNzh3L8slYT+SD19C7z6tGUFB5HxldxYHj55hgeaxj2lLSS7
0HfchPM34MnVhPHqBO6AkcEXV7KlhMx0CIjiuh4P3aB84UIlSZRKz/LnzNNwcrFx
j4N97qXKGu2DfJAQr0s3gGFCIonBTQJeAUQizWdNnVpB7PGVa4izc+82JGFEmnzI
NJO/pjaam78Gh8yPGioUoqI0zDUuw8hf1gaMdVkiutuWxh8uKxfJ1xbPibGiLMxz
VkoLEDvj9R5RCQvspr1VIf7hP4mD+FqQe0Veb6ekvHvQXFSbKjXb8XpGozcib7il
XdvZu4AkmFYTl+L4NcpuNrqMuYxA1ezvxXglm8z475i8lOl5rYWNqvOWCNI68NfR
HmdgUFDjLA7jPW67qBj8B9P9AT18OqUUbbj4VDfyQu89QEExUetIVW3TIsS7PgM/
amIWmEuidGWFCc7eI1LSlo7Ov5s2E9c97EIwsWQEAm/r1udddHjQ0GWOvscShYY2
O/okR79/pm05FuZMTwOMW2AB8dSlBqw0J2qUpIEcNZ7jtLkZg+7kRO0SoA5WV86O
Y61Vlqrvm4xkGPe21hhf5kqotJ6slYH4MAkQFInKiZuTRnaPwiaQz+kdL/4M6xhB
PKrqnRA/ifGj5YlveiC9kPNTQXeCd5F97MKjBfXdAiy2FUfb4LfTppPxUCdSZ+J3
cFCl5dXAPRdXU4j7fuYeR2K97eHWzlf0m9bGdj7Sb6QlGi8GclRqiBzlbbzRLyb6
qW8Cg2Gu3sVp2W9fAbLPqy7A0MItL8BsWOupsap2OlzieQ8A32mlBUmghXRiVwEO
Mx2jgA14MMhQNnv2cs3XrBSBcbLMp8xHGtHnqpJIYzXXbvymQ+rIdIj7NhKuxKQT
dlR6B7AtPwkYVf5k5Ri4Ygc4iidt4MIEqhnin8qhR0+kdBTo9NhvGast82+z5jDL
tzkx7ELvp28SqUAHQdfJ5vQOwPH+aDWXLLFbusWSPb8Z+dvZbuUqUrLmRwKF012p
bxfz6iR7fJaKQAZLL0OryxATBcixHNKXnEVjF8gcKgiKyXSFw4QgTdpgjeuKzxvz
k479Z/qRnP2RgL2oiL0B9M7fuiTkvaeRyQOsea3h3nyLUyWmg3vLMq9wngzXV7MN
ZvYHJHreJaoqPa2GpugEC6uunMIdAsJEG5Baf8NXri994NXmHKqXK6jZD0jd2YJ0
fs4L8tU8vkwuq6lknB5ZVS3x5ZimnpVQNBpAy6EqNZTVr7LbejCWs2JBcSkEUJws
qIteenBpAJT+lVHEx9sb0iLXBF3HGhac9Cw4U7Qd31W9IKAjSg/Yd+tIoMe9OQNU
WDbObZv+a75W2ooz8AOqvZPnIXyQegj3Gb4+9/m0HN3lfFbRajRJTO1JyEwD+p9H
Z+JA+ROz8h4VvRC26UUSy2W16yfA4ByJgdAG7mdSOyl4wciYfRSJXBG/po9Ojw4Q
KLn/JbrlMmgi0KN9EwIaoffZF9I0uSmXbmjRVrsM66nntsCRFBJ6uBpaUBJOP25l
MmmGHyBEc7aI287M23P4FQ==
--pragma protect end_data_block
--pragma protect digest_block
hIwhpnAQSOm66Na8o4V8KF0yUT4=
--pragma protect end_digest_block
--pragma protect end_protected
