-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
N7ZiDhZ+v+FFPVnuS9mdxTo8K5P5+IOW/TI5JZIP2W1XEN4Q6EkmueAJtP3OCM68
iFaG1Ig5DhpBO7Jjka33OrKSqNmCaZPHO9a5lv0ba9tK/mVtYDMeoxd2cJ2rNLAe
MlUCM0MmyLetkWjsR+ywlNkgnHXbK9Xo/VK68r7COAM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 39354)

`protect DATA_BLOCK
agcRmCrhlLQhPJsoFGQNvTuA2bW5Diho2OgEqbNVwRK0wxB8EJa53mXyFkYZezje
xtjl5MmwPFawO2Mqjgked85FF+CllKz/Vb+CF7hKdw43mY9KGEL3zZMeiEMM+hv5
qhTIM+gldrGXkm5tcMn3xxCuaPo782sOWpbKOeVjjGc1rQQCVgMslKzbB08D3DJ4
ZVut8eYQ9Je07ewxaY06YkBelXbdXiTZJ9ja7fjtLS9cnM6abXwZvv/Bfl+cPPFq
AQ264U2EBGKRuhGwBIe+MZfHTyq4Kya+f3wFskaVkt0awpRErm1tfJW+1UucRd6Q
Sz2AzkIdfbU3bTS19Yfzoz6lXfLpmKUdMqXsFTE1vUJYxwxwVBQCMNKdF1Ch0aYw
CwRhhAHarMPwh5SeyfEEqX/WYHzgD9NJhTwc1hgxjeYReAXJAQG/DECndArpNtpT
VtjWoTRhAbfIdckXn/yClnfkzqxmQGLhnXhkkNdtQk2zrnL3O+Qf9NpZ2ZX4Z93Z
jZBoZFJJGFtQvjRAGXqDdjWD0hEQWi5uvt7RgynRY5f0BsSJ9siAnDZ3/bWKr1u0
HWHimLM17UkN36BOgcEKke1+ONZoLeToVpjyWhBft1jqmhzKG66mP69IzPY9rg1x
L1GJ4MckAify9J6zAKT6Vdp8iQSgC76pjPpKF0xQfNMBjD12VovuhXnRHuDb0vxf
0RI4dHu+EbQKfOLm8UPYkuZQle5ETQmssgOg+leabVvdEAQIzXVnAxztIMcfynk7
8E9QeCuOhmXfd3+79WqTuILL5OCW9KHKGFh4XUxoq4KagvK6eVN3PLRc3mYvqP1P
npeii7s17BXbxpWnBwjjlKCWeDOLMF+86FzGE2bbFc1+alSBYyrSgM5Lf0xUGYur
7OmM2oW6A/b1OeTCybOX/H2bVlyRMVEg0JWZ4omdpgF71zYIMpLCQk/Y3dUglM9n
DsmAcXv0A4lVyajBvYnehPBSohq/ehrfeK9t0CfG7ISdxzcwMjgq0LYZKt4909FK
z7lb8Azwh9E5j415btYd0S6mC3/KjzU9p7Cvp9daRRNcyuX5+7FGNecHeJzAeK1I
bAnuwKbl9nUiXMW0bT90ITob3WGFCcvlVXZMHKmJCr/goU4sujwiGTW49KlEor2V
WOZ8QyccupnRpdBzf3lYUvOm5sNg+pxIvnQPIDy1QsPb7paqqbH6bdg5JpAxHHlf
NKA6fBMM5kyokvkRqp1XfsIRJcceVxj4bpSoMRIwFl007FT4jHlFqN+6/7X98RDd
9aUsk4wc799I/FCvlzR/+H83sDj/UxLnaGdIo7+DI2/CIiqR//FHXR75eBXsAZ13
6W2FrFRqQeC6V+UlLwppHJ66Q4vVpRgTiepmrstFYHkLHVVE8qpZElBCl8gb0h1i
DjlXsw6MAxqAZaBThPBbApTT56NlJGRC0qSdXaCueQWQQsQVXSUJ5aLRc2avvVSY
kJNESlIP5AnWNCIxClCp7aGcaiDLE9fIDTvXAlentVQX6TOF9LiVkScWu/naNciX
xWrB2JHhcPuRGzLNS7IVKXKlgmCOZTetvdj2ZKeTzAHLC/WIah4apJUUlgkrtfbN
v78bHcorgbPrIuqIdiq7OQxiCGCYIS39hT5Ojr6tyJiQlKQ6JHZej73DgRJK5DLt
+zIRUcomLjvi8fhwKtq9NdRNdrmpgGXhovY31vd93IFZg+Qbi6H9MbjzhX/8/Q7B
UtLTK5Y1EYRn1Wcdi9hLXsslcAfKjXPPzyWWqdPNTw5ctbW65A38E+9POq2kkRYr
Eys/9ZD6R8PGes7j+fIyd42Xkl42VO0VNWdS1uTpVvrwZ1lcKu248o3WysXmOUAI
fWPdf8vP0CWREOMMo5LEb9Ze77KCisxZGUlI6hRli354qCcvVZSNHi+wcbgD/Igq
syhIW63JqCN47V4Bb5/Bcsmqfi4P66nidHDaDnlNrK/FOek8wiYkaPOq8mSSTnWe
6SbEt6ztWWoWy6x8Q9/wT86wVNyj7zXFTP92u0pAonhTxcU+1pm0N7RoX+Kb3ECC
+9Xcz68c/BQa8o0+XnFYDn4HSdHtlzisU4+9rS/jRGZEr4jbhdYd5uzQY9uznbm5
qSdN+Bh6wlwLAERIr5+DLquz/s3aWhHBWtAAad+tZx+1BkbSPH+KeoUeMrM4ykzD
o7I1cxUk2wB3J7DmoYFGa+o1VHg0thpdrNm+uO+3zN+yah5N0+hw2l0D8rf2zSG6
sekdRvnW0QLNl9mItRG0MnueMsZ3DJ/BT//Fk/1ezPBfZkCFyAURpAmUouXV10QH
eNISev7umq8BbfUZ+R1316594lymk4wWeGkUmngG/rp87YZKqBFqjJH+Qf5gXqZP
c7WU6uNS1x7sNh7b/9GYfzrV5ef8i1i802V2xDHkyR+9sVZmncbMbfMjFtpTATi5
k6RREx2JFCJKn5H/LOVTCAkOuEFOhKbOcHxu+VN4zQnP8N/XWV+cotOU8I7IrlHY
mC+NaVK17wp+cFOGLVlVLJZH0tBWoVmIsDZzjIb6UILcD9WCDgKaiKAeTOxxHwBc
OxMyom/mfpshFEx837bV2pSMcgre2ezPByfFYVjJPOPozDAnT8MtrNlULsaqrKGT
BndBSRCTlgyEJecdBJZOOQHq7qW1iz6WrSDxlMcQaSwjTDJOFr/B/S+vexv6GYyw
aP6bNSJPNaCLoTtHkeKDzqghqEVEojz5PYZvVBrM6XUhuYMggUTBW4GFAb4spiby
n5sQeTl57sSaGSu+JIFVlr2RxUrBMYz4vX5TYz9h+2nPepD+YVEI35WIbi1PO6V0
VPc68YTJt1pHIrQYL0brOe6eGkWUyC+1L5jHKen4hRaNhGW194vNdl9G61dxzHCQ
hrBv2AMIhK/ugaO7UULNxMxfm3+eq2hzNmYZL3VFdFER0+ljkqJuBp2wNWJVEAIL
1E4r2Grae2duNUVIXO/t7pcAgWsan1jQafECcx63RieiDnttXB1+OI+DA6Q/Bju/
GrAjhzLvTZZnbWKRbjwj89P6lobU7CnEObgYmnJF4/keHchvmYiEAtk5BjCjDYO6
8Z9Gs3ZUwbtUZyixF8Sr+T6gjOViikd7MkyDTXRunu1owJwamUzqvYXwzDgcrRm8
rjoMcK0eV1j2hOyxmyAVqYE8ZGRfVDEeFbXYfggTh8S1OjG3fDRaSY9GUAFDQgDC
XWgs+byZTMaSv+cA35bRrQ0nDZFl2WlqyBVrWOUtOlQPEOYpTrbhMHuArTESVWIp
0szK2WEKHfzL+PTnHgpWifki5dSIVMKeid/5N1TegN+h6K4KxzrbitZHJNJF8ezX
/EuriEJwAHBQj6G27joIQ87VyM/zTaOhLh5y9E+q71co8MR0FhtqX/aDMFCyfAQ4
473Rtzz/lPTmTdK8CBA46AZJA3bZx5+N4YHaRDq6UOkFD0qeUuBokhF/gCeCSPvP
XnKmltRjAER0hkA3hUZPX6NYpGw+W2MME8i5tOVhJlvMUsHQ+7SAtescVLO1RXiz
5rmS4cnqDQO0me8xmZPr2CcRml2laClJpNwliGbL3N0PDw1yxkF4pc9MA2myusBJ
XkPdwFimYStI5tk4hZc09czPiLLho+hz6KccxkUJGcyJZ9aKbh0kLH5q93nUNUkM
rLII+PqIS2KtQk5IyN/oPynxLnzUxE7yqolQFO7beFg/6LgaN1Ez4ZREKOL0qRAo
Hc4EVSQ7sQYcavyddE4EOGNwQF3FCwIKWEWEOVIVH66EQu+KVPo1a831XkqaGKJN
5HUGh7kOmm+ydIVNPsKNmkyKwdG/9NamoY3TYgiB29oGjOa0O6RMzW/SsSF1mZz1
iDhXAx4xGoPnewikUJJhxQSrQv/GKOzfNVvMbhWUtlcZiw/IQdt3KreTPKb59YRP
GZuBjR0tKIPbpjIN7yPSgFHg5lABixr00BkLRwM3HD+8pXDcIbm78JTkTpAULGEW
qufzp3a5Gi6W3sNibCmAO1tkdocaVTEjtOEsGlnTJY+wsS9bV1iRDXTutJlluWqR
61K2PHcqQkjBNf1mAsbNscvDwBG1s2xaIoeLNv2wDda6O+iqy7Jt8wNhx0Rx8Cvc
kV+FKCGaRAYuWWEzugg0HwJnP4VurJ9K12LewOUD0YZceWrrBHXiA6VrniC51O95
2NQ6ppFwhouMqN1emgLULmWazI4e69P50stmIWccMf5S7adkiV4GOMKlZaBkGNX2
BQ3PgGlXi18U0ayr/Zhkw8QZa6lx1mtULw2Hauu2rwVEiYoyuAqOTXmMOEhHkwSl
7twpKXLkrV4ESQKWMjvZx+LjnK0pY74lG3RoB1WMoO1OOrQUui3UownTpHTlA217
1m5I8lzc+b70S3qzvxmAHEtgupluktb0H7f7SYFJsykE1rAWpcwj/ReW9ns9DGX6
kfNXDPbTfRfrgHqpzGESPvnDKln7NrIK31x2WgB3LNNKG5TPOq0GdV3OrXMKhGln
L26XAXRNzcNUjePMPdkqpZ56jViXJ0KGSeSdp6YcjkoBG/NeLgeVEdS07xv9sZ/j
NDgFjZN3hlIKBPwcB7Vf52o/+ayPxjOJQM8ij/VMRmGuogHkM/EEG7YlUAKi1tuK
2u/VhfNn+ebHLj7uL/NrWjyLxs8MrtHjA0TaNBGmhGNsFMfOH6ziQyA94tA4X4Ql
+pEPhfse0TOKpiAyD5svzAoOcMmdj0qcaip/d3fqd5CP02k+A7XUOoMgTpzpqUn8
52f13S7NNH2aYGLJhNG+WiA7BtCJWNvbSGkKM8hrU1WeH2o0LTqaqWj4Ju8nIkC9
UyKc1E0UhkBKvs3sg7NLqmUS60pvp2kFFqT/xqgSrdDerClrvN8BI/Wsri6s81nV
yFRC3roVaATtuzORp2arUWpRXVWZH7Zi4wHLVUautOV+b2GXCJhOzUwSqALBFR69
q193KCSboaQBJHF190hRoc0aE8W910JErUIFtQHbXAZcExFO5rsqf5NeViY3D7t/
rMIjUqCM4SI8stMf5iDT32IXwO75PgVTehBvGyn0uY2kyMjVbQXcQMws8CHDh1Eg
SlcVB/GBGo0zIDwYpArwx8szgHYcxC//96D+1aQsil/g8G3uHc0Xw04yjTe3Aa97
x3bU22J6qEDBr4JCeJSry97SgFrzlzs1cAZsyZBHU/X6tq+PbBuIoIOlhUPTxkd1
bMHgIRefsh+bSMV97czo2JSlepPSizSwLUi9yAU57ZwJUVLOPjHPMffezVrTurNK
CfTWujm2ak5K4JkPuLWA+8yOR7iKHso6IX+tXmajMYzePfr4WmMccvSDutbObGnv
BcaDn14avlxXH03loowrHk9P2eAp+ryKvUjDmR8rLvJ5JFLDFrH9zTi8ncpmmo3Q
mdTeKVkLe/RCcyo09ZBY952FqLvmZEABduGqHJ0i5lRFFrNL2SYgaHXlbN2sBU77
m18opzvIVt7D9SAOWvnw8MbF3RzOpyCNLTAc5WhpTPgh79jsquAyTqGSe9nDVtYd
Oq1Dnq4fGjRG+RUFWpinTYoO4tSjjJad5+4KvM2o0orYDdiLeiwWPFHXv4bF/heq
Y8YOL0Jmd8i5edLmLg/qB+/uK+jilnOG6QkW7sB9ljvAoysBYpvk3OwYZKB0m3a8
H31LXonaS9jw8lUU9BxWSp6/CPYtyLuccUiOFyToFCxlflMcGTReZ2LWd6/7671m
4vkt6N2cN9WsiKsDQn0zTFiFLm6lmnmt3VnFu28Dwm9HmFn1zm46Iqbf3fHOx0ZX
Lvt2O9yCsBkDTMngww0ElIJfh9c84X3kOn54I5K2EKefRcB1DO3ACkUid2USAohZ
11L3LsQHLfC5hI3xH3IpJTzGBWi5daFo65pH45b5mFczzbZu2FpKrgjMvsJAl+2L
CXn3iMTfsv37nkigojqWZYHrXkALQecIhTgG/wWVL4cr+zwFxwelapdvCOy+xMgl
oMqgifSCnP2SMMU2pPDoLmyVdv0ZNO+vOVggrKzsOGfm9WwEP30mqrrb3WBvnoQB
4UPpkLVRNevTH49H9C68olatUQVBHm/NIXEJcPfMKOCJxD+NZddH2CORn3OJwpPO
Uu2UYj8PW8nVrScwUaU4Fa0f2FBLUWXHI2602VE7TFojrs6DFgLtjRtvg3GKkl7e
mGQEy9iwg6TyLE6LC72Ya155kY9bMYiw52VnlljxP6I12DtqreTla/QiqTQmJn0F
NhV/yjGyli1xOsFmdOdHmRYA+vAd79pcCrukPFrXmMkacCsJ+JeAkRQ23Egm2Eom
3LsnxHcfx9BT5aOMzY36oB3ER0UmcPBk8eoVPs8sbrFQ7j84tH750+q1GwPhKQ6/
yzqVoZjK6y6y5iS6W4HmLQwKjVICj/q+UaeNIT9sr6jszHVlqOlLVuxj6/YRvXPY
bcs3qmTmgdB8JF0U+nIpjHbgUezixsNh5ALwJDSs2zcgTRvOikFPULlG8Pk6o5Ld
emNS61HYQ/EGtaiUov5MBrNv8ruMrUQSSHdvmFckf/hmsZmwUwWhc3o+q84rJBOb
DZREBfdT+URvzzuuX7UYER/Yaxn11bEG0BaTY1umidAsMqQh6Rg67wmlDPiw35sW
0OrGLjqGCDoe0JPGh/0+Y59Dg/SJ3EjeCidrbJZszwCnRGK2+bv3xn3wMegyGcoT
rObquCDf04qdgRldN8hqLW2rvAj9Q+hPgM68N1OWqcUOJzNmSisWCkeyDYs2WzAr
QkNxch2d+FLp+0OGdikqzwWQQtgNfxTq5/EQJB0QsR2HPELF15ehMoQsPI2Ujjcy
pc+eZzGMSaAEQGi7m/yZhNnwru3y5h0prj0RvDM/MfSnZRpsjhcikf/gB9VjkLDE
rEo3Rb3sJCWyTWA8XyhTnCOyBjCE4Bz6hLoRlKBi1xaok11Cq1rgHOIYmLnHO0zr
HgrjNGrwOV1FCxswUXptnqVBmuaH4Ck9Cdg+Mw8XoV6fKc724tEllohh5slubzS1
uPf8B1VwDIV9MP5eSgiZHNljrWHnk4jb5SPbem6ifYkyORNQfY6zHQMXqVmSoGU0
DeH5jYbQsUGJVtgYJSmFx1UtW4Fysw3DFwpw+SC7CU4j8N3q2AMXEPi2ge22f3DB
pxqDjh65ergRQM34OoEP/LK7LZh9EZ5D2wjbqFd9yoia3qcgi6qwUSX2TaCn3mzO
MkVglXe9w9KakHTetOL/CbARFbcM4FfekOtcbTEcmhA46w7pII2XU7xaWKLgSiRs
kcpyDlooeNkCjQxJHGojxGCRmaUxBUv4a2DEfI+ftTbb8dSAIneuHDFSlBwlQiar
doYRWQPdizmZNihW5Xpm4T/pKf1nleD+C1XNuc7Bl5n+aJ9Y/m0+eQCFHE3TL4Pf
G2JUckm82xe+fwyV83jC1/ELATM4S1rPpOAt3j4OOwMAbykeX8+0ayFPytZYsIlT
cuU6cDX5aZ9hxHKp18zioGTuzx+Rn8t5it+a4Z0k0K4/L8iiQTd0/ROdBdVwe/Dz
fNg4WFRxSMvx2nSn4X0bQ2RNj2RasUarheFP4/U7azF9+k/s/l7WbjCSCy64nOrq
PupSFAciDnIzMPJ6e3IVQ8067a1t/JvJ2rV1wSX+iFDgv6w2u/3S2VGnMS9MBCbw
cDoIvefzRX89JrjgHybwCXXr0SMX1Hsy9B+07EAGR90oxlsw4KGCp/qZE7DHJvlv
+GtuVRlfebPpE+ltPBv6SrIgilyEBK1RBT4FLE938JFMJsunNBdl94TWO1w1dhqs
ysjlPt2KHdF8ZW5jnzyEeXeJHzf6Edm0j5dmNKnEnRpY8Q43/qeyckQePM5TffL6
6Q5EzaOQB8zFgcPcm/Xo3bdNRs5aJUp+8nsPqkqqsJ3lyRfnNiKohbNnl3LAZwBQ
hYIGu1e9itBidBDhb/ysY/dgY1SPdqBwaWsf6lF1JDmxrhZbz1wglh9mkL3KuWgt
CCwWHHAHxIlaHBiAe58f1Cc6bfcsxwRaoZadijcCd4hg11L+/tDv66wJC1u0JYZy
P5U0s0yxyZe/GVBqErZWavMV1gguRLRmk+DSK7NzIv1gj5JMoa14fI+KSioWfCvN
5RaA5gVRCjBAyKkGacRCPDzZnp5/IVmkQK1M9QB4UyeTTh7rRgtqoiFzNWkOQ2dF
1dOyw2rCg/jEQX3pkpi+r5xcEwfUUemSKs4zh+01XYSDrRaaQIGCun0IYK1j6dHn
DbsR9pbmAk9J0UF9L2wqx/zoL18uvsmL1PgcGB1L2j0QsWRPYEFNXLF8w4PrNdV1
E0MFOTTz4pWcNdU9lXpUKbyaxRReKwVinWA4JmINISDg63jKJWPduOPieX+1MF30
rAPPm1/p/+z3Hn7gopu+Cyy+xyfVRnmsrklIhrdxAjpHNqkeW5aWUiI4UyixaMqJ
ZpQX/ZEHrTrna9ve5LlpgUlk8gz/uID1EmD4yBvzwexfvfdT6UfrQLAw1TgHldkv
oEkWyhTXPk2zdtOm1leFyiZz4cx7Pj3bVhgYZrudm2LdQlYMEq8ILtjwKXK3atio
LCmJLLkYRoeT30U6Mt/stwXMC3dFZ+Ut30hFnd0O6uEy6jRZU9zTZ0L4UFJlfgzx
6Yf9mzY2uIhS3ykfHCicb2WfVcMKuH4oXs9SfMANbZveT6IJEXYwn6mNVW3ZqlYJ
I+a8DLedCv2dW5bHmi9Wka5oFfQsLz+v0/SpdCLeDJYQYlDJFabUdzihaLl4sAXi
HZj0PCt5aZg/qOlvz0b27Cv7otqmS4FXegQxeRxFItL0Zx6U9WFQPXS/faf2S9da
+ro5IrPFfzsqKlyO7EWOonOqIMkBYk3FEZ/5VxjHbkJb0i409xescc/nvMOL/cAX
tAV9iC3mC8pUF9lIiXe7xGX1PzfdMjOJihQMhn0ntN/YkjNadXQ7IUirl87ovklB
DiM7qN6onpKLLNrU786RpnVZqwScwg0Ihtb26H8VwTTdZ21nDi5VGRGJI7T1ZyBp
O34gc1zHcCoW0RQC1ORnYcI1OSRYIPn1L3LYv7KPtKFU+HQAYq3U4NqGFkH33duT
XXEnRACoDYTXY+cQ+C1FPt/pZM9aY9Kw80WjeQuEnD92k+o7D1nGfXO9oFFG2K+y
KDWdfL/jk1PsaoJvAjrKUJ37aBk9w7L9SEoVk6GrBbqrPap59VtIOdnV5bWwKA4W
lTimKS2YKa95+zW8XCbfBGSPw3sfYa0gQHDRUjRpOadKltsJ6JpgEUWMb+kM6hsd
EzQfYaK1/73jvLgMANQkc+Esw41MlO1tFKDQvliOR7F7zJB8JqlccWCFKB5u6L5C
3TXFkc31SgFuuqGWdTCD1ud3TCBEbdER6OsG0bem4lpQ+TXOrCG0SC/swgLxhLgs
wAk4wJTQuuVv/89KUTh/7SfJe9l+cbxayEREFM235FpwtogiS+DDNeUGwzpStuqW
L6HZn4UFzTzGBBtd7ciUVa8YsRnffoBDbVtH7geWiQ8rtvI13hYYvFH+PCIS48WJ
1HTDKpwbNzK8DPAEuDoAC8yrtKk68CQF5z7OvTIlN2v0avbqi2S0DfdgHJLaVFpe
ZEegU/n1OtjHljHp6oKXEl3Nz1nqY5IrLCqZxv8KeOQ7l0AbD9XYsl1WJqn5uaOk
nThFw819wIDGImQKHlPu1r7QEg/yAjK3BF/TksC4P6MF/u52qlWdnGu+D8zt8YkZ
/yNYYDzjtn5SF3PS2feL03c5cyFYbnowJuamyoDDGpRNMNVTC/B138zCDo3bIj23
ND8nUk+fjzrui/H43P+j8HU0UIIXC5Pr62Rih/qnEJdWgWqAYa3s+BQtGJH4HtRX
1WcPxae5OD3e+HAXGwYT7wOI9clBX3RIxpOSyYAwLdfK32WenvnjiRP/ouSX1qSE
qb67/YgUfdqUN6iFxM5TPs80PZDs1CxjFXBJ6g+/86jaOvbct9SlGmDl0JvkhUya
pZSReho3oVcNdnhFqKH2nnYERAVKeXrPd9rlhTMytfsp7/C+/I4POtbQ7Y7aVebo
AD/07j6fmacOIEkCHW9xpfaNtut7ZNF6JyT2S9844eigIMgZtFnZaSTmDTxqDcjP
Np8/U3yNAwBE7gW++yH1ujYzUt/IxNzh4dSCQAQVn30E2nkSu8NeoBUkdWYw99gi
dB+0tqXv+0muQc2pfF4803TLDOZuNfDl3+PT3Pv17U96B1hjnE7JnSOJ1Hg4Y8Lw
Ve37jFwBD6fN0mX6aZ0gJaPxK4zf7Gx7N1DI11j9LG90CWQ4JxiL06R+WB3saso1
wxhXWsWH4NpAPss4bWDv0PvwShkVUOm+v5H2qrx0F13Pt/2gFyeggEwdUY2ppzJT
ZCQSYVcE/9B5FcPvEiVULnT3fcfk1XaG68R5DD38jpsUeoFD5mO38nxDsBW7og8t
nIzwc9US0OwW0GlUSpPdNJHHdpTsceqNcBI7R//P5iI98D+glwB+5u/O2LQXRqs9
7yhevsVbqdhkqwdBqMTPLNlcRtgy/3LJmkWU7IXird7SppO4mhzsG432olWIopuN
MRwqt3iyGk/2R6E9677OYN2S9UxvdG6jXyvRpfPcwX2IY1Lwps0rml/6vthlwPvO
1FyFdbfxlZlu4cYidpC/iezLqlE6Tm8sHI1eE8MM5403a4Fsw7XiJRCda49yitgV
q9Gj2aqeAujKDysa/MZASsMfFUP0L9DMhL+g4FTGFFRvHv684RjAn7PrXwE/DNw9
fJTQDctoE10N1PeeK85u2ufEAUXKpZeLF7JMC8iv5yb8KSnmrq26vMafAmVg+/yE
xObV9jbuqDa9LnULINOfGVBSy2HEjkKa4gUabaw02IvyxXnSjXN7vhvaWczBvaiv
reo/E3sdQYGiS7q01CdgxQOqJ+eD0EyaqMJG/cE9i8yNCIof/1xI63a+V5IZ9fQp
cQwtHWmK6LRExmOLPIdH70huU2/yPMhJZGaojl/FLMIRS59HF9kxH5yTVJh9Kc6w
QuNnuiQMV5qoGse6LD/mhBOSFIYzxZM04hKtDSQZixgNGkGqG4T8YKUG4bDR/BLt
JKwj1v6BW19YIKR8PTIjZt5RAtLjo47sDlpk6hagTHKU6W0Ba13JMQyLvGNbV7+i
nRAQ8D9CJSBVZVgs5hTaIt6funv5IKJAhZ++esgkPNBB7uzDd0gCuYxIHr8Zyf96
fPouOCpZ7/y/cqvp5oJ539SZM51w9qglreTcFuscpo+9/KJBvGQKu/AjqIOJkKHN
PyMWVt9I8oDi76hGC3ormTBPS8m0sFNXW8Bv2U27bhkuzlOMNU9XvmdZlTCf49bU
f+VaX97zlNm16MbUHm0zg8PUhN5HwvQCnXnqaUIkeuCeqt/jF/koZ3r78DOCAw3n
ONsxZBCB6lo8bBR9MXeYmMy0CbbfI735XyU4nvt5wP6tOFPRHiyKT2xHETfN6Wl1
ELdLiS3HrskSiTNtY4xeF/fSkhRi0SGWwK1JApT3y4TvSI1cDf4nJ15foSUdK5Qt
8y5Wc+VPGQbb1u+zH6b4XbT3qroJUiVqYbFJdJt3pxlfcIjNJSGM6ar7WTtVcs8S
bzRlpDkN3H7YjLGhFPs0B33f3IRkB3eAcG40VZtIXde6Zh3hxnBEOICcF+1kG9OV
BdAsfN3RxUgE9jyvvqeyWDiYxa9ZWLirh42I7wMk7guGm9ZKmXGPBPg9brqf3kS/
bHT0YYGt3cRFnAdOMg38NdNdFjEvA6aTu3p6B034MANAJpeXQXlxK6OoUvEhd21F
DAi0wcFkakjdsCnWep3MVmChiqxjSXZIGRiI/c/uBXx/PJF1qLm9y82EJ+ytK9q7
3Nl+OTiJ8f+Sx9cvVvWyJXyDi1/aBda+G8YwoUsRABXvP/5h3mtY7qblfVgdg5a9
51Sz9cSaSSrRzJWSJHvXtTWUt+x4qoqPnrLqGJWgs7XM6bKyhBjX8AHEwHN2hb1c
HhMUo8oOGTgCoOzBrnxaet5VwLgFifALS0V4J5C/bNjLW8AYoqPGznt+XwLsObkX
wR1dc5WIP4uRHqFc8TCI/2JPSXGpwUzdNCCGe3lSUrhZxqfrTSeDckvtsMDxgcdz
uDJ1OF3ksDl0DlCkuH+wijO25RoyFW+Ki7dZIsWJZIUGE3bcCvJZHAA3MwuM+i/X
bhYfTEyNqVzLZF9WykCZF+xzFq40d2HluQm/csbKqGJz2KqBGBbSMt+ctedk8Ghj
xwi2aWcLylupMMlwNLrWyZOSN3h6Gw0e6046o9KmEFjQ7RK8INIr8aiTq8Hl49jP
K3lhlgyDy++GvCE7s0w2voHbL19bZ8Pt4YDBswV7YycsebEtW4RonjjLGgiqgd6m
fllPeiQHEE/sR8DwWVsBhiIm90OAWlFJav0VjejnKBmLxNbRbOLbvQE5PtHeKTPH
1szE3/nLP4ZFQ2J2ReNGvH+0A0FJQYMeNmpU8hvcEAkF47clM0GrqqlJIkgo8fKu
AJloZQGnjkXlYFH0Eg0f3CzO+HV4/6SC+QdD4i/2VHqcMVOhjKi2gz821cAjfpfZ
UloNc/VHLCxUFq8HXmt52qYpGz3DVzTGMFWnntcYQRFt3sMJUsNflLr9lH07V2MN
1dCFtl04nJ1cTZCmeOth81jlouodGuHASL05+RbyUinmqOVbXDE35CpO1LftKZce
xniOuz/fZ0r5eU8vzH9Ej1ND5J9WaxpWSJdYRhnpPqnaOCTU05uqRHC7nhJFjgn6
oOYN9rESXBmU/bLPzRV04VFJRD9IoPEKhZQo+c9fez3CJakSH+FnZjlbwmLS0jQe
vj7b8TKBOUNB8ho74w76Io/y/xDs0qyM84IdKip5l8MJvkNEdNFi4Ke6w51fDX/a
n/Ujnyxf10Q0v3BbgN/Nrk67MBLoeJfHZ/UXmyyC1ZirOFSNweQWTho/b+0+Ziuh
kHh1Rl+1u87CPeEaHIGm/EnjyjKToUFdqvyadIjCLpD6tJJPLbCviggc/Tz5EJoe
9NyQM7W0rhoGL5gGglbiMNMWXS7jujSRnGc/rdXnlorJC/D1DqJTUTgWk96GuZgN
iQr97ZKUZLe08uY5E03DdJwWKnx1cqoRp3PTw5qvHUimIJLzAf9xVBws9zMePhlt
IvbYHN6gHAeMFBPv5qbkcjb3UKMQaNLFBfpx54kMBGW/xc0+ZbwgmHuOGYTLRhgb
DbwNBuYx+982nchVCNPo0Mjh8/FaUhvJNRRDdZE8EH0Sp0nFKbn+n+8aodA5U+Xj
Dw+0c3J3ORnBacqc6pQC0jAuiJmdITQne2tQK7MDt3gOuXv+1ItvZQcWQErxz73y
pJc0Z+ky7LfCGsiDhb6SKmG2uw9DC0yRIH6pcGFIEi64EDfaC02pJ1dDkw0dHq5V
HcFDS1lgZaI/4MN1xBuTBy8CLQZ3zE9EsiZZ9EErZARB0Lo+KPtYhg/HIYz2o5mF
xdptoSmYSsjfR2QFUAtSbzirz8P87Ats88MlIBbtYy+GMh/FlDH9e214R1bJBpBU
C/sOFewls4tyu1D1zV3BWoqbZaobuvSomAJ+6RSDpTslwJSbdsWiMr68flXDmcHI
VJDob023iHRkKnWsHjk0AIhF/NZa10cZvHBZjNMToAx9GXKr9weyTIBWyj35DDDF
BLFbOLXAir6kUZf4Ei0MAPucPgIth9osZQ5umLYWjRhgFxS3BsZLsleXBoX6FC4m
+ocsXkmvNvdXQ9SO+gg1vHc1rPq/tjGPbQLlxW3Xn9Kjcp6F0njIeIJM2xBBI3xm
p8mQ3Y58XXk7dMx+HekFFgUFmbpSPwa9DKOSq4I9c/TGJZamhkkiU7o8IBCBxiL2
csxfeThkjWx+fT1VrFoGNRa1cN3Kep926VvN+ucRLcPQI8E+doyVX36HiRw5d8S5
JqWX5noC+ojN4V90WBclfJIjmw80SfAk9BU4fHiv+AY2kAwo0xG6y1oXC/524Ij8
vPRNJ2HphNWZW53i7LpGru7LoRKXbl8xuQPIqYwItiDn/xlCygkjyTeKpj3qf9MU
gbIHnu3VC6AivfGgWyzmG5FyKLRat8vPaP8xDne3zSrfxxETw90Q113PwIUqQ1ui
uSnmIfD3QC5gM74Yaay06zdId5ZrJ/P5pSL2rrcQsD67kUTsOGEdFvcBrrgdidZ2
XPUl5oYnLtP9clzqTmLwE2w3np0QKSmDEo3sQVsGBTLQ20vMvvyUEZHEuZJnkGQn
mrWPSilX2FB0/aaMS2Jx7j2gkXC0oqI/oDsrWFvtnxO4/6mnDSlkDUOls48J5KWx
SYZH57aYkIrRF7D9hCNuvWTzIAQWCYV7b/RX0UYF+dR04mhDQFdg8/4S2hlAVKI0
afUS/vLA2lIBN/xNn79iPa3STEQ2JA0SWuTB31EyjT8Lrrc0+uqMaaLu7nwC5EVX
SjKnNbE1lNTSGa6pmPpW1NEm39DXfjVvFcnuvEZroGZmCrdTim3qDkOjXFbUerya
bZ3+VZCECeQ9WmDi8WCb352yl+q2mRd6iVKcYYgpkVQer7tGpYTHf1Z6/uVvwmIp
Xc5e+IoOb1TFAbaPLUasjWlWmjUPEnWVzuWZoBTF7RG+HNh1fhOVlRBtPJ0P5wX8
ZaE0XoZyvWEFfdUD9u/CNU0+f2WsWVQ3F8jaY/ETvPGdJ9vloBKYKQdO6e1s3R+j
mj/AeV363CU4vWZZFBxZhYKyHXvTvcnrwkZNm5WiABnvr5Q1ZTJ0hj5yeNfd2YDH
VpWZR7978Qn2qIWV2yNyZyg7u3o9QwU1kevZUXdeVsgPzM8BD6Iu5PFG4AdH8o7Z
ChyAqrWGmkdW3TVRcmsHrP5NL6eZa3RYDEevxamKctGpsWYmTBcmsXaFeMKOnxLU
hS1cDtYgCSSDaZwGyHYpQA+flVMyLxaGqB3P9I1GZ+utskmlbrL1+EKWctsoxWgK
AuHHzcv+Hv++rpRwLDdNUjEkg7i3mqqOsmzORPA/+FuZzuT7E1p+MtEJYQsVDcDZ
l8N1yOOFK5FRv71Kk3bZCabqwzHZT4WD6nsRSkD+QjHGDtRlitLboGZNuad3xRvl
NP4fK2pF8jpMJbbLO7cUhQxCVbV4RXUlaWAB3IBN6XiXySNLr/VFgrOSsMS22EE2
04S8YVuXnOLitvFGsT6qH4ItpDIrDlVr/MUGqNO9Qx0knMvogi1eQjmCfvmy5ceW
pQu3S9ykalXfiEKs8axbykn4XMbEdhd2wiIHw7rKD0+xi5jjcWsY1SsvM7ClK6F8
rrRVBX1dbiXM87qMxRBp0N+Cy8wq/l4ArS5dSJiqKS/ezY7nM5LMMS5lMJdyet+u
Z20KZ29q0CzRy4IfDdvMSskLgVzBuF1IgeirZzfA4LJXI2kZjNFCfZOaZApG7b5C
4nPqCQvrmEyqDE6jt3+9V+UcaUdIzb/4tTn/J5UeQsICxseANuJNnzNexhBxzd6T
rJF0JFvyp3xmmBeFGTYknmg6Li1PTxf7+ufG+XdG4wqM2rbRRaxFJXPXPa7XmGTi
ipJUI8SAzn1KaxPMr5a04nk/p/I4KcHevIlipQsaZt3Bu+8KktwIt9i7mdwyFiFx
mjHGfKj4RrvQOjx5auGPzA6IFZHg6VxlW3R9E5l7ohI1brjU1av8hi0uGWHuIQ7O
r5Ctavi3SPbRnGOPd7OmtDqShIYDwFoADoa8HfHjd0zZKpucQsdKtHdJ4mZ+E+z6
ZwsRnQSUlSEbLnLngZbxUFgnKyme+xpaqw24uQo+qrlbqHsesIene7WMj/2euqso
IYNRAfe5gt4qJN25NcMMD/0qfzEUEPBO5ehJ2vVqXv9lNveaj7R2rYRS6Dc0uX4s
dzggiOy8i6hTsUW2E5xjMCFjw7jDLs0Isp8Xf8DfgT2/sJ/JvvL0bcBNC5Y1+6XY
7fwT2El1gB9kqZNpdXYQl0fXNt9NVKOHJPC18ALqqSKr8XN/Z8JxyL+2BCWd+3yC
8mtsA50GQR7Xlb7iEPE+v2c9gwwAcDcz0zsHFKY8mGENZk3VTzuxQnRts28rmmG8
dMHq1wq/UWbydQleZv5oD2RJ6cwbM3IP56ety756BJbu/xfYWT0Om1F5paGqHeem
hFWkbkaxiJUe7Dt/i/CNcqTuBw0gOdyB3UoupRJKtDjOmJeQucL8bZV4N3YLRM2i
vv1Aq5bmMh21woQ0PixFwp0hDgU8b+Zn4/BxYRIwWddCnQFdanJM7yLP23sfpawi
e8QehEJgzfUJMTYRoxyoYDW5cFPCHBU41cIdTpxjDTcp+SoyoL+AoTmTn13PAPsu
XPu91BsBNqqtv7/Tw+Veg4IyNMB8QJAkYO6rr73Rvbwq2QgplPJGhNk7SSy57Wgv
Jtwt0P8zSlPPasD1n1J3vXvxwRg7IUnkqMQVJm6jrC+v3VMCyHbhDHUSk47rUlXD
BM5CWWSGS/equXF6TiJBA30fcQ54V00frUrY4FBBpOKVn9h89/DTd7qQ7jFFlfe9
1iwb4N1oiVK7M4oDPaeL4sCGuXZwaj5pvFtnQwfcCe/gR6JEviq3e++Wb9W99LOs
p3SL2m2pJXISFOU8Iz5/WsXy2dbl2eFfZiTZ6TtVOBKvRCmfAK74Kgjnpim6sfZx
oNoz9rcQVYF3+Y4iZ0nZAe2KqYGSVP8TdxX/F0FtoX0R9vbgb4fvuPGxomp8pk0N
fvmUApDwdekroRKIxgMSwn/iUH3OQLbDc9cWsPFrAuK7K6SXlk6jak3rgceMhv87
bzWDJHdf/f0NWdltCrhdQNPh4QvhCjaFHn1t1TbBG4T2y8tOCufFakmFXdY1u8Rt
6zhCfU+JVlj2trkkH1MiTrSZtpGP2PvPHFDtAZ5hYPVEkGwLU0e3DJfCosBiGymv
VvOO9RxUlpUB3PdCLDMyPr1/6Hc8ZWr7kqMwuH4IvuwErh7mdy4bWJYGMYciv+q5
HQi9UhXzQif+3x3tNQ9ALnnXlNREEb232PixkrZz+f9wcnyawzEQUs9rN4E0N9Xl
eNuQE13VqB+EQmlWkfMOADp6oyYljtI/AAJhsvm4CfPrda123vjt4cHCjOgqize8
mOVjYxSljhOwpFXUPO8avgnm8acxWjUcRjvQTXMtkp8wj3b+1qme8kzziMLHQvDO
oDDxuVuGS+PE49bu1MAMlG0b+/czLWsxsdQYJ0Em1xCqzqybC/ITFaI9gTKQgkAF
gWisLeQfb8hRStwyFNlbyAH1qxTGcndQhj7e5jPym2CLvSzJGPdIb1xbKVffZOwe
ezDqGBtop6qAtuOSf0V+HEjrxyXTHvKIGB2vAcmuZ1ZQR84VpeZgw4V50cBWcV0n
2DT1IYt30uvdWj3qUmC0h1jfgu822g9h18mtexzGRNxsapqWIt79zz1KoUu0L3DM
Uw1+sicGMc7ZvLQtmzZLNwpYLoHX0RUcwAAyhmVkvo03uAuZruwrlPietwWzZA28
ZFHs5Ffkd/e2FEFWmmogLgM/lClz++6YucqHvf6VDqRpx8PLvWHXi1bigrzyrWEb
Ah97BWo90oHm2xWuvGd30LHQsEL1Hmsiqp4GvJEe8I8nZNUeCQuFiQQkeX7JvZEP
rvm6Dm2S7m8n0cdROAj0+4K68WWjV9hmJVaF+gg0UWD99RSXJevOHgB/Ij43BweK
TxjdvYSKbBGJJBW5xriJwekeVnM/TiJoDay4cvvP2UXP002Jpwl6r9izLcPvcuTl
MquLQWtYsEGSojuwWTdSJd28/d6Kz7YIUKelth28OP7Qt1oRbLVKLJWY7/ddttDB
OyyaeXRG36o8Fhv+yHj1CCD4F6AT75kyIMB61MQDgk/LCzBb4CKUq6mjh0a34Q2x
dEtdAj52qZLpNldAT6LREFo54PwifcAlWGi5od1KkMlJDMRGKG6astTToCvbQiaQ
Nm7JGomfU6NmVR0ebCBvtZYKDwbe3JtTDDirui27FhCsntYh8046zmk7Xj+xsShu
vEteIjrGYQc/oCHzykqwRa+LVUOEBxnJ2jju0bDIyqSiiw7f2yNSIKwofq81U5En
IvN4CEX931S7mVQx/LEsY2TIwrlS+Qmv/g4T91+RMJDzwe1XXCIi2YjpTuyXnVyk
NmbwW4/OZQjShK8ZsqtIAt0Y5KTZ08Qc5HP4TMM2h+r1ObhTcN0vX9C0UTUcnjrE
Icint7S9pWiZyHMgE4WNLZGPNjdL94Fq3wPh4ioLjwkMpCJav87b44XqnoEV/MrC
JtVdCKkZ76XqvxjjwrjBuE/5G+se5Yk5KcbCwq8nySEuzBRUQ35mCUAXNpBSiy+X
DvSV5OfbcsLphOK1nqY+pHQgGXvCCmevtDHQnoKsz6JHoxlNwlgnVBH5PHWXWMkz
rCTlTeGQ2NrHXgn0+byOdIXxTCYOG/inVa3rdJ1ti5y3dwIX0RiExCNHcasV/yn9
vTsiq61+eGaYA/WHA1UBjzS4ipbEklLTeLdgq0CrtCIiLkh1yDbc/8WHRS80I88u
2FqXeVw0c74IX5L4iy2HeR/nvIVjJ9Yoh5CHYpOEEBydHiAHUkCrr1l44848FKzx
7+i1M7QLDBflmrNLN2/2iDk7/D6rPsUjLgD0RhvxBAazujCaf5EkgiR0No+JxgFu
Im3mim6unDRhS7acRBUswCNKFlAIIUItko9ttT9bxOcTP0PQHBLD5YRqgL2yaE2a
6vT3xvRx9CY2wZFzcxviqprYc6fFIYr1o+z9mETSNpRpNdZhQwyDz34CGhsWdqys
dRJM82iZllBMeOS0Lid5/sIhLl33Wst8ZQ5moMcc3ksl3hHMD5P8MMYkNOi4BFYO
Wat5PJbMjpQ+ruTHKYkVE8W6arymo8bK3yphnEc5qwORXP+V5yMuQU4vU2codmVz
BEbR0d1y4m/Ayy8EUEr4Po54lM17+iUKVpYE9oYEze03oO18TO2DA2PfCmIB2GOx
xlH27d4ZLgW1MZfFLohdwskdFb5vPN9PvndNN+/5jtZIJWnojywUri4AUQRqQy5/
XszsQ2G/7s3h8SmKH3vUI0AtuyQAe33OHfvw1GNOrhEHv4QMGnqc2/yQDr+ODKPy
mCu64tUyksIgSKGVoEQB5cuXQP+7IH+nc+Cu6YpZFighxXWDLzdxa8lmHvXf2k7o
s1bcJ9gRPACApxF42L2oDc3FPcDrGG+Ri520Q6cOrK1NBmyAiVG3+R9cvBEVSbLz
jPvlLpj2FejTbzPJWSNpbLqKrx4+dQ7llrKKuUN6PNShKIkp6XNHpZSHdMjvY3So
g5lwAGpGhhloaeTQ4OgKvSqqoUwA2ewu0NL1QIIcCYkZdH9/NCf1djiedLn71ipP
4C3iBmG3alELj/gbpbgOO6X7EoLqkCieyU4CzFAOr96hDzkOVcu+Y1dIDYocvt+d
twpppitNn9wc6BniTVOHZbumXr5bcGhEiF5lZN57/QG0yAZD70R1Pah0mL5Nov0f
nntZ/tCycYcLrHJe9yDe49IWBTe787o5ZBiKs6DcjnpWbMP3zeIu84yptn8im09F
VomQ2lsX4NbjWPjdiRw4IRVrAI8c7PSzEqVDjm4Wed4rgjiPosYa8CKkq41MSgJ6
S/vVDlRf011lE406d7ChWUA4EMsqbG7KxYv1ZTfm8HARgWsAXMFyMZOs6pJLtJp2
PCslo9FWk4KXIRbOuqVSIhm0vH90CLXG5oSaNWa0kyWsE1fRnCtWbJnuHTDFmnf1
YGIs93oAqBRl30kZcofiVzowT0ZdhSw8IGciOhoqdo/T2QNBrWnsN6Oo/LFA9WQ4
IMuPqhLolibgoBAo2WqNWfGNIM3giv8fGb27AUelCaEOYNQFe3SteNTCm7uBEdWe
IG4RjGTNkpLvQp+LITIJQqlo9gsIIkUJkIu2myEpPOkiia262BQ03HLFqKfuo7sz
iHG7MmMCL+2zwpf/u83Q8r/gbUz8sZIIHDOCAFwFGvOs4S/P7SobLVC8y/VgNMVO
ahksuQcCUcpcQwsihMzWCkgdyvaBId8TGcch2Df3zqzBwam7mI+DrBFih2Nw5I7Z
3/cQ7nrByZirb6yH5um/eT71F2swe99vutUgc5JOxCARpQC6xIFeEIVM9sInh6kn
r4N8OOqxQABvs+LCelYh/pe0YHsrl97QTAfHCHmkpiKYsIxjSiqbl+zxOwcsV1cX
fFqgwx2NeGz8p0EuiJO+CddyU26ojiBM+iC5sGReU70clRr02RZJbIaYzl4jqlQi
hztYLThefcK/qlW/1m31CAPRBli++LwB6O0yiN0Z2m53hSS68suFnWkU7LvEuAx9
1nNUv87TdL8B2hyElS7+pujuHaDEDOAev6alkW5/9jKGLEx1JE4P0xI5s3t9+qrE
05Wg/sliElShw7p4ftvm51+2qrlYxWQz3F5wwMNRCveL6SA+aGW84hYCj4eIipjO
wOZFSBt252SpX/F17qMXyC90kKmsW7W5xEzs/fpD1NqLUsBVq1HnUBXmO/FeOHqb
qs4sddpeDivYGWzghSS6CEF6qRZTJ//N4LyMoSQ1qXOQ7lnxqTBcAKS2p6kEwG65
Ipu1iIy0uz3GfWngbwj5H5ZBM2lzUHVOCR8q+9afriI1K7Zu7wHsnRLWJ7LDl3YK
ldLs96DU2kTW6MI8nUGfEpi6v37JUCN2dC8NUHa8IauIe6BSZNPKXPmuJXNULPLF
jdZq/ezamrer4QNCS0Jj4elY2ZTP6ZdFWekpbYv7xYM8vTuwAlEQAnyXNnsTDLKa
pc9T5uvankjE3pOCTcvXicHM4vPAmsCF3HIv5H1rYhxRCVhomfucfT7TpUhpi92e
2HZ6Zl4Ddfd7s6LMbKbd4k9YfHKh2kjlFD/W1PR0TrrddBAt2+KdiGcGvpOXHfTc
LpKqFk1fSo50PxmqX3ElEv3vnb7GDH5FyhuwE0kN8u8LkrqEx3tdZMu2ZAXC9O7d
l8HTRky4S7h+uUEhCSSd3Y1xvsUof7pNGBbpeUkm0kF0ajYcTu7MXOLFlIGw91zd
LS2hXs5dLAzVChHm4J1gmhAjyT0a5DzKu1HxNY5aNd878r2pVkWSIaUr7vNBKMip
6L1Cp8bBSEKCKVKILayPIqTl1P1lF61nYfeVKMfhdtTGBvW6CCLNWAgJTvE264BR
iu4f1zgTIkhaJ8UQtgH4lHBbJCFqdC0aQdtSFtAFNYSKt1vG7HdZnkG1YGCKgUZk
LM/aS8WJXKJ1dOn5NE2v7gcpoYgpqUs1nWmP2418Q+j3LPg9WbSmleSYO4OwJFYX
HkpJCYWV8K+pX0Qp6fbohClUl4i+SeJvJf1udbtGo6ReAUz2Z2c4kQkf5KO/307v
Teak8JtJHJ0FMCsvsNY5goHIiy3cAZdcTtZsR09MprXWKr0pF9mABU29siaTjbd3
275h2b3RknR8NkRJOGQ7VZ1J7WA9Xv9KLgwXqyROymfpIzudrLlHm89Go3B5t4iQ
HFQRwaqQU/QxFose6+V4ik94tO8vqkMXfxAhS2saFiFSmH345gibuUFWBjbfC3Y1
Qg9pI/7LZDreVnZ5Hd1S1LWZPK43Lv+OL+gOLXEBQ9QfkZRMbYHea4r538Ul6CMe
i8As2z6MLwdPPUo6OrNi5F9l0BZBnDklZkAqnHICW/jeMWDo3T0PG8N2AFU2sMU/
11TEXmBxCG2pFucpLKHWHhDtPfyS1TTaZ9Mf7rQk7shNLqnIDHqqkzstaT94+mpb
ogMI1BpHfvs2z+1iH4bpt0uJVmvLzWW+ffjX5Di0nM/ZkGAo5lgsCsdFalrmZngL
1Avl+M1QV4XF7JkrTpENyA6qOZxIWstoJx8CYCXSYeF61p7c/3BI0p4KxSzBBoKL
u0UsEF7HVB0PChMmXXEBBQKyxYH9D/QN+93yCbD0sBYLN6gzkmxNkIxMHe10sC6M
QwirWA2Tg3OMmaVNQqTgHmkZTh8T46sJN2gupg183pf4ZqRcwWt7eFYvUu9RCbUO
lOHrKdztzKvHmOl+ULYjELrbxvDj93xCAj2Kyrxg/0Ck0syKl/juyOGMcyjC7Jw7
G4fei5U4tNt06UKoHWhp5F9kg9PKXasEsKfWEA235oJsyvtgi7NLZsA+g2suIOpb
HgcU4aAuxb/hj/O0fyh1hArEu6qr3CEJ5drl3jUBy+Wm61+qE5qOynqALhoJxZkQ
Ini+0mJET91LNl8jDu95JoDqhgoVzbkrstiBNqc7pqjN8jub+ePvu9fJlyv3Z2Hs
h89nqNerz1E9cXlkZ8ao/9C+4WH/6ZspqAxzh8JD20WXMkiLOUi0zwfb2USfkqV5
MqR3XvwUe8WknEQaogCSQFtr06DVgn0SGI7TZdBzITIHS0VpnUIAJUFFHgVE15Yr
bO3v6kugKNpOW+jqzkCWuuPuboqomgU/CebONwlRMV6wNrCTk3SzKXSg9pXNs3mx
Pd4w8Z7tYpydxHfHrImrpqPQDMfqwTZuNv1zmN4vhw+tvODB3nFB2Bg8E88fh5ri
VFPDyq8DwKuBIXdDEXXGwv0XzfawZ0yve0L5KBf/tV1DN0fFgj1IeY34QxAdY7qL
hXVy0uLDaFFLFt3P0my13BD6NBmvHXVHsvUxsqerpvsZfI51H5I3IMyZUWSZCSvT
iAu564dBmh/pE7OsENoD2C8ExK5msotDHKm0GmMk8Ahp4r4DrkhPKIhemxSr5ZSo
ETn8mH2KrkwYJxL0iTu9e0759nNCDHfcnfb0y98acUaxfKtAvLxW4iH+b7hNzTv+
TIUfo88EPWcv9p4NqsYxj+gQKUX/hLOuRI/OfphvSNsxGIh1mhuObrSMztE8bV6g
9ZOLKBjyZgPxvjjZ0JmgQrnNvcxtryJtS91yZoa6CzHsY8rd3puwPR+/K16ASOJ3
Zr4tSAjI9QYgzkKWDYTq/tP6rFndOXt9fPUBnEv3gQrp9Jmg7uG0U3xcXXY0++vt
ZzOUQg6tWMz/t902G/X4A9PGR2oWs6PZME3JINJHL2wXiYZKFjUtIXGAnVoyJN80
ZtNS+sDF+48/Ra4vgsbl0YKA3A8RltaD1CInidoXSZPP4DFWe3pxVMTWYyBG6e05
mBauaS7UdSAZ3Gnc1zvCU3UKU4S7onV/JPuU3X2lXIH5zCYFN+7fBFSZUK+rUPjK
YZV/JeIJm5vYK9O4MXhGdI8bLIIXKp043o2bFLFRgK4YF5b1zKbd1hRIMoWLYtAf
eKoUc0doMBKj0mee0HcBplTAuufiEnOkaonERoPRwYi478wPOKuSlkE7y6GkoLpI
pKPpIlxjR9qKU6ewbHqYwan/Rgxn4QDsnSngzuaO63abqZJ6RpqY1L3n6C4N4wfK
e6Xy0q5kAQQvw8Bhr3dI7gJeGZ20YtbRL+lC+5brewcCZf2DFdyA5zSZuTqsnBiK
72LoiKTDI+dhinpHhvLE1wtwBZpm22XMPq63xFINQfnJ92hbF+t4ddIQK4O9SOvW
15qGUmRh2tdrM/S2fssrYcXL2f3J0kAiV4ETZg9xDnjwQ/Ri+qsJzdEqZuT3/aHl
Ed8pmvGlEef5pH2FYFY2UQbECewCK9UxbvLbaiY7aAxcpnLvBR1O+QbYNgP8VxjN
/bKB+m4ZlONUTEGqpotAhN4/RBxXFZxaqA1RIzMmWB45wbaEmPmGvLAoj5VKoCdo
i1BNKyO1MqFlBa3pst66iv9bR3i44HMZJYm/crQHrzskFr/DKl7l2eyr3r81hs0g
PtwK4Vlt+kMXV+V+8cQeB2wTPNTPhjgwlOl/C6Dhb2fAT63bgOD77pzQpcajLe2v
0/bkPyASuHEBFJ1Zh+lbFINI0VokTHeoxhWuGR+MY6TJmzHJwPwfi0MPMTR+Tqhs
BRSNPekBbHH0W01okdlvXSUXlGVXirTs7av/smdRyRlqkM6gd2Awv0sQ6lqMDt2i
PFoZHFCZo2eu80xj7LyN6Xzfe+nx99iwJiQtZQWLRtiNRm6BEViJLt8O3qSac73M
ws5KgqQHjMXqWlG2NUQuaR0apQL92CY1TUNTnf38qte2yaGeXLRSfi3kFy6dx1in
LU7/XTT3f+WNgc3UzoZD7q+MI65Sj4IixU5FuwdkvLW7ZKbsrO4G9t2DwWOhgV1B
T9kOoaNzocwTaAGghhAUqohSLHFFnePKUtQH9vjP2mG3qKXE5hL8fsAllNhN6Lni
M4NEjYqy9GMsxx/fGXqyK+2QkmsYV55LYW0kjPaOhytfFfPTC43n/fOU/NT0nDB2
DR1umMssPupTV2GTeXpEEppXQjtfcpSEWnocQd53O+sWhDqWpulXM/TKNf9enT2y
OSH7/Jnu7FpjUl1uzjIEkkImk65aZm+4rW1HgEhDr49pTYrdRQRksvxbYsuAKkMs
cOqfEGpznW1VnWgo/b2q1eu31s4bQbnJiuWSjj6AfLt+uUqzG+QycNvWy10mG8H5
4+vVRLekiICG+LAaN2vxjKBcwbTwKF2lGcz/jt2xVBJTlGvd8o5H+COiY+aXhM1h
KAcqyM1lnWBJDGqCMDlByhyE6hbul5CpymKY20gdoKSVq1Z88p+G3kcuIhfctEDr
AeIpIw7jfEDvQ5jwIfvVUMCEIag5XOwNR5GYnUAuC2bIjHVCpRT4u3VRsXmZkJKS
gX0sS9f+R6nsY5MLw1ad3N9u19WgQFjCK0IojomBYqi0woNHAQE3sfr0Ijg4kEXe
4uFX1DeXPCoRgwXGIE6tJFDuOiQ5zNGSyihtK62CE0ZOjTCiPNEzkbSudwPLL9/Z
Wb/PPz7QtTIJwZfioxFbMsdSJG0FZAEzzm+HWbbk1h+19O6vX3niWB5mmz4c8Gyg
r/swfwsUiwaD+7q9kMxe1gLwy+/JbaRT6q0DnGzkKZcN9QoSGIt5A0Wwys5udTgx
rlpDskvywBQJpebQnZM0F15OxsYqBflvkji9JY+hAh/3bhbhljd0KjGyN3odOMCt
nAqB8CALJUNhTcFHAnNglsCZtH91GOsfLwWbnh1T7eAF+b4kVsW2+2HYxn9aV/ry
ncwIt4XcuFIQdLIBJwAXOk0mqyzVXGWJxc9BD3InatENmaktA3AtC3FK2Fv0E4FS
GxpdEoP9Tnr0OuNCBdq+3V2pdd/e7/D8nEm3MHoXCBzkLT4ax2al8nkQDSTdPG9C
ILulG5maF44sZjvqLZwVp75VOKTHGi+Wa8keZuS4v033yELdt62eb8edh4v8yajE
YuZUaw0NdFHMBCdPFD0s6EBE3Ca/VZdjvEoIr7C0R4jGxZ9/qjgOPlDtpK0A3oWZ
sg+Ks1q76Xtl8M90LYJV+qZ3H6ccKZC7PltuLracCDN37U5juocuFv9Ey5hHA8Tg
k5YMQqOA6exk1uAU2qZNJBpAlJUCtLAWizFLhj2KxzK+RYnhd6NcSI+RlG3V9PIG
B1eOuEWugZG2qhxYCYDwAsfLQOm3r0+9HiV1Bv5FDEvNm4/fv3gKTuO7duhLYWWf
mNnfbK4gk94+JrPThBxajKxyHljrDoc6cN2EjVz0UaW6ZpP+d1Bq57+9ia6htvms
W70wFrePKYiK6pVuC59cv6tiJsmers6XijvGJ+774hSgoNeGrQsTmIWItL4MHeer
RBAhY9sSE5yoNvX/AaL93B2Ye3HPq6DJhMN1WEUi2md/H5R3bz3cERnZG3mh9T2/
bpJnL1UOV8NJdNzBMcL3N59nl9Zr2eJ4yuq3oQGoWGpHnDTCyXNiKu51dW2/l8Fp
vweUf2MhMMtuuxXBMtmB/rILaH30+4K86+iqyHpq66vSFcKRecr3L2nrFF/h2CfP
7LSwFMiEvaVp0TnhHIcop/sa79tgwleWe03KN6uru3QXekno2LG5AH+obG8oGQm5
BZIROoW9pwNk/YWnTmv64T7EfZNMIbh+luhpX9sZeTsOw7urqb9tP3KGukRwwe7H
RQJGBaA8LxdQA9LkCvjTLF9ZRJhYfPTL2JDWXeKDvukjkYHn+XMOyqsXnUWEASUl
WtAKX9aBVEF5RqnUDi7dJ35jrm/h8nI4vHTi00WxxL4pDXuaQCgazaxzEx8WLwIh
NMaR1K3hy/3xvNKs7zaKh6dAcocVmGSK1aKaEcUJZzrZ+tAroJxe6XHNSgPT0Hdp
EGYeYDXnjOlQbT3uwDOB+s7fDeUWmOCnKSg9T4dBRgqlz0k4sVZds1OYsiQ0QxCT
IqQ1vLXeS6uiCEZeF9onrFcyt4MkC/xn1T6B4jVr4zaa+IcZZ2Wqg3/jIpASyfEb
KrNnrAE9ZMEoF5d0gnP9T4H9DtEdVo8NDOe60SKYav0GB2cKHgYeA9R4D6K04C13
S43Xv1VpPvEKyouHgJ2Um9xHOo3x2jSpufYGBiByh7yoNSxGRW9XLu0JkYIqbAZ6
nABiovuYBiL6KCaO0lhFJFoXm9vQkeMdpyk8mEln3xjoehFjbyfrSZ1ymoEUTu3u
0kxCsO4fvN/myE5KGLwZce79bHyIuDEzx0/f6KZ4jfNaQFMrYaNSrKs92jpJTO4F
cn6Hk1+HNjmsM4DMF6gHmkbM8Ep7T0jlhjhhEPp2CR1c5D8PD7Nqhmy4CZJLWS4S
1OGiUW+InJhPQRn1n8zv8pdhPwCF/7qaL9Kt6M2FWA8Brl8pWdArSfMLzjDLIMRV
esSfLVnv7PbcovC/cUPL6m9cjlijKYpZXee1BUC4/aXGuNac2zLhdD1ypzxxsvbC
xv9gdTgeKbubgHRlRzd6VDZV4g/ervBuZmWRohAYNfJYBaOS3Lh2q9SGyxXytCjD
TefcjBykO1K2Bo4aYka0AV0iPq8aiQok7xL6eZyHqsIVRReLMb/tPmNQ6SLQJ1q4
Q5fWQugzJY7gqZ1/3BbsP+UmpNSWUfcI+JQ9+KbJxOHDaz3mtMWyois9Bw9zNbCt
VgnmnXbqMQpnTpZXeK2LghMbrAc7uxWluSGrbopt7roXcEKK/Mvn+FjwvDbx9aH1
tvKboZJE2Dw/FUwUuP2c3xz8syrnuT8eS75Jk31ECkwI+2EIpa9A9H98iDeUelDd
aCA/iF/KNjmyqNRrlmBB23O/5mhia24/SzjLLj1EKLXRInb7eczdbuFdfX8fXWJr
IotCBul+XJWeL38R8gY9ET2ceM9PA337iSXsovFNAmNm9UfFdtsSqtCek9vKr1kK
SMCh8BJ9PmfYIG4O1/rf0t6QA8gK89nbUnaCEAAb/hmtx5y/YIg/yc6obEMyLsTM
/KnagY7DShTRj56/Ie8v1esr3VtBQ+cGUJI7Ps9jGndziaOmH1jeoYDJNQGKMUUK
ADiuj2hsJBwrSgfkZg7WooTbRZ4IuDx7ijGkc7fvIWhHehekkDyX1dWbTs7lIj7O
PVqluW4tx92ldNP73g4ODOnqloKALOmMLo+r8gPDks9PUZ97rT/NdZHSDDaDIXNd
xNv+1ev8wzevc2WLu9G0AqtkWLWylOyBOjZhUHmsxsfqiyxgpBMhPiNV0kiyiblw
AEF2J3B8sdFr9XGID+bF7HCgS3goXwjVemlvFeOn2Nq1c9jIx7vI1vvc+j8QJgwW
xEx1pOtdETMU1SD0YXA4+Ej6I5g9kcIdeWufkS3kTaafI3z2AOJINGYZKtaauW4g
rrEPyyagUzETdYq8SlsCAXNvEHqgQ824Z1VzMpNOVqGofXdXNoAAdTH2rtX5nJ4b
60w/bIJm0DJV2fdQI3GerHyRNAGQ7ofKUiO5WRBTd30v+CGf4JdSeW4ZEDzJi4c3
xXqEY1ahypYvhE0qjscn9aNtlQM99cjErDYldZC3E7EKzHYlRdsB9OtEYqjhQULE
cAU94dp9nX8YK9zbJ5xl3GVHNNLpBqQYk3yAsGgiSo5eWzeoT33N5z6YW1SWKfI/
EJkKzD8WvdOjWvHGDtxERSl0bBF/UkOLIz4B9UlbbUptxJENTEsr2emnUQoaIi/t
43ERa8ciaczboc0ifctolsjTyQc9yhgs1JQTWc8E+LZosNtT8qhOBdzdCLe4Kitj
fLvCxxjO3DLqGqcX1t6a/pMRcPaOPLbQ0DSOlDjLrIPxiXzSNquvi/rEb0EuqhTE
Y7CcLcI8emNb/wE0U5osPx9sSKaG+sWS9bGhZTWttTTRCrkblDdNrNxfr+MJXueZ
/nyZ/WU2uOAQ9z3QBMpPZVuKay0xloe1mBzvmGnXv4qhIhQHbZxDvEYjt/nbJ25T
yjC4y+XoebSl5AIuA/MEyihX5gTbGow9I4HAjKlWdUE+19EDCHPc68avz93ZOmvH
UNn6Bphd2GhhWBqo8aFEmNb+tfif7lMdLgNel2v7T8eSxiQv9Mu40uv6uEonOsNk
psSUCMY0UAjfEBTy7rB2RzyvHwkrSpmYcYi3H/HfCwQDT4fPKbq20bc39ZNekuI2
ChUIuda86fJA1pYhOdgCNcQdtjPlthHrlCwS1vc3J7GGdcJDktnaj+tgXEJgSdyK
RDigIdUs5qyO+mgIK0GFcmOk/x5Y22Dlun66Q7oyKBMKFNf0ns7YogjLmLmf0dPG
84TPbAPf1XDuHDi/93Q+ba1wENKL+i/h46QBBb2W9yzWIgC3wIn9gDA5mSDVnnlw
yYXz6QGfgKgJZHJmwnrKvbWy5kJ1swASFrJN6VzlYlj85uBuGZbQmygUznySascu
5Vqqc+MWh6AwA9yEyXUhCH2c+j5bC18ukTqrMptIE167QUmk+Tu+BP0znUx4XJGW
qcy3KvlLeSME8wpeU8r/jjFi+q2EluE9efiB5SDbK3NOEmzH2Qk/yDbLYmp9fpgx
TTvARcCnL3+JVrBkAgZ/Fvw1p/yohoXz+/rmVOg0nArDIDIpdXXL2VMv0oHn7kZq
KT+wVOPCGaXSY+B9uo5QvasTzkYtraMpoLUyAKuUwGUdWh7dfbe6TGwH40QUgK+t
V8K6S4iB1Ro2nDTSvxtRIVyzr4viJt9kAKTozHM+stBZjonEpniAkKUGpeg4L/os
cOVolMqaqgt37IsKehyUaU9d2U7mhpEflTfnsdcVjAqa5U4dhwKJLWQj5760FzxN
5yN2Gsd1eTnn5NJ6qfS+tk7ZlG4iBWApQghZO3gvJTK3LIgTcmgpA5jQCFpQooFe
Vn5UygMGn+Y8Kun9WrdzlunEadYoIUH1rmPNvtdE4qGKgDS2rxJbZDi/llrpNlrS
o++1OjK+rqsythiGIKP8ILQT+EupiemTw7ovt7ViMmD+0udhQzEU5wCF5Ht0ubYd
UEO9X9e7b0q6c8feJXkbSpEMlUtkQz795g+/OTrQshmsOux43Qa0crMaGCNpfpCw
eV045LeBq3nrWcOQHpP2/B+cxT1zC8uhWvR1T0Dj/FxsGUBXc0RFFuuxxe4Gq3y7
z+aHuZuuG+A5TZ+9CeUxyc0oJz6tqUIPPn2oDIObQGLI5sUrmdNxVrd7v+tEVYOq
pT57jHNiI6AgLG1Ti5nVm9q1hGc2/A2Q+K57zsP+zKBu/nyHz+JKcmN4PRBJQt3r
Ja1UsVvyAIqYsI81qJEG9DaGT3eJX2mzlyUvkH4ApbwRRMIZsVVeYLDUKkPjbw54
+Q64bW+W33iVFINngNyFiq1lhX0wYX3Yj+5iWQ0W75/h/skXNBcfPDIFH2QVtU0T
O5ogy4BkX5rovugZOHPNK/70ryxxXd8SPp2x1U6fTwZNDnXvLh7bPOT0PkzMmPHi
nL2UgvvgAXD/lV24E63h0+/u3KwAA9mx+vKQAxEJTpzRfgfKNg0Z6/VFRd15+dl9
wQNf8UI3ncPFm+19kiYtsXkC4Jf8OhdtK/mF4URMD442diLJghGr0YTL5fYc9UQe
stL3zG+LW1XrgMy4/m1VrAVtdoEecyvTn1ERsREiGzRyQqMiQZW+sdMpX1da93uL
aEk3c8UCJwpmGULFO2rg4apoZOKpQBYa18zC08llNbkb5GlMZpGQcwz/ca299rRA
KssYNP3h1QqUaaIVQv2w56my8GkHidwwPbNlHeFJ11SdBuJxFGTtUDMfgKsEMbdk
TzDyZ/QBQnyqnj79O6vm9HauAFVekwCOQzl0KbkZoCkkD2xK74ZcazS9gKUSNs99
WvosyTM5RTM3r44Fhoum077FFAisE1YN9UkR+GzX7xGWasAO2tG196PkB34y9byL
07F07d4ZtI0GbfpTB3A+T8ybs5tOuqsTQxi1xk1ATgtBSe9KoFn+nyfKB/MhiLrB
GCRm87poOG6NqrwW+l5InkLHUBse+IJ12RB+5/QVav5aJPEAQjLt98NxL96Cf2oE
5DCJpIImXXy6cCCv90fd6IEOK4O3G41+1ykEaye2IyXsNsGqVSkYJxHfnc4Xt71f
2BUPdIXuDkxngmmL5faUDDOXkJAdaSu7dYZGLxFbk9pUAle3VYmPyOsW/+qNyfJh
9Tat1/LmhKSVOmp/A+Xnf+Ot1oRU3q6DJYBleUFI7/bVQ735ithDmPq/zzgmwTS3
TqOtuIFEIu3svqKGJcUt1y6oOy5GRDrPu5uMqfM7wMNIL0JQmjh4ThMwYIDIGbPx
t4oItepQr0KE4+QFfB6hZ48/WnmTF7SwWVR+kQjf0LP8CJKhnfN9t+fB167sNQqd
lW8fImLz/wPq2KpzDKnyzkGg6/AHY5MFNfaQZzp/mJAGw5v/MjSFPc3H9zYJphMm
NZIKwsaaKv3DidJBYtQW0Iv4qn1N1JCuWkC8LNuMZQUHTurqiLeAHpshONveKd3e
7cPStQ05oFuRxnyYN4ZjvD8MWUatnOsHvQ8A+HhqehRel7iHHjwDk7scnaDLoXEG
4HaCdz/NRqajbUiG1RUFTrNj5gFzouNsHZO/rRtxMxYGt2F1TZM56exvJGzTvpCJ
8/CYOl57OOdDFYc8eGy4HcKpHTFdW4X7LqL7ofeX/THhCln7Xpnmtpcc0fIANXqM
vVwju7JL+gB/TktHEx8+tciItaz0ZQkyD68pEIQY3Z0MGRPjJWRr2Dguh5bIHn/r
3Vlc2O58zimMGAKxjq/TWlplNRDs/BmZMpHQ80GSE2zfr8U8MR519nZLf6BdE2Rt
t3CksPi4eP4E72fRhWRzi/7AKLcfgK4QgE14rbvkIM5fXKNTSLKF9fBNfA8mAejz
iHaQHEFpwK39qrTA7TLXLBo9UUki8vBt5+NuZeqoJU3A9JCD8bxug7FNHTsFHmNl
z4O5gC94jdDPHSxolrbm14Mzs/v3XLtWo8pVQfE9GnbFceLI/HElmOvMHwROC95t
nLncxvgxms1GtPT2wBwn02MOlHs2mb129oQlSXX+25K/R6IhTv9ONBWFkF0F45HY
Oc8E6LsrldsQay4LEJTwNS/T43KSAQAgEw/Ccwx8aNbBpGtAz4plu8POl3L9cIkl
iZ2zicZLE6x68ivcJCnlvzJw/ZkSlJJIlUnj9JlodGNInTB5O2s7vOlcuD0wCzCZ
pJtkziNzMALr6/+VvOnXh6nGfo0ehlY5N8z5FRTJF4HJyC90OnBIjFXfqtPCqNCb
w7AWRIrYHOYhPv1jK1jXvSQYfENs2Rtmbxl0U9Nf6dI6FjxgETLp633vS3tw1iqH
tmIZPRakjtkEA8+WSmSGzePGcgJI99zLyoFiAfrgQZfj4sLjez4to+GNPv0oueDC
cFrA1mV7hmLgnTgKno8Iyp88dABVUtSwR2O7GQa0kaY4vdtYmvW/+z1UlwXubznL
pSgxNfMjh5BZDhZ+CRlYtCQJIZVY81PTQ2JyVd9g/mqPyItvvKrGxkeXShyH1zm+
JLmd37YxUM5SOVYsbUdpdcvN2bTZHLEOSWQx56JP9UEI3s0HCHqQrKclqt5aOUKf
pL7HuVIj4joRox4mLgAVAgUFENw6DowFENX16uW/XZle9fzaguZbbi2mnr9yU3aa
gi4KTGGxtQ9TSuS43bPaVR/4shAJwuI80QQxAJ6xArISlB8tA3zsGK6y83+CH4FV
k2bWdMNjRB2nyTAnzf4twY5EhPkw9m9wQm00tpOCrpfEvGBsG7ffHTRYbFNEcrE+
bFdZZSJvFep2cXWw/mOBbtY0DfpJbXXdlSVFOSV74tIGwi0hnCRASRgIyio4dIv6
rKutTjNALbZF2RNQEQuDqttzS+HRYBmgwCuGrQciYRZt6xRlIUFPHA7UAsLA/gdX
1Cfk5nMjHJ6zG5S6ogmZnXR139OTDx+NfM5gJLfNcj794s7NjQGMIT6MGDGZdJ32
QF3SHpIRCBkMu1XMAt5AePxLpASUqgKrQb+1d89SJb3wHAP8s7IX1rT3w5Ftxjh0
mC1G01EkoQ3Omo/E1HkMacVmnr+PdXg+K/AJWd1ck9D+rQKU6X/aCd6pVOuGxOvC
/2znlAAytaeq+tF2IyoIpuTx78aKl2SPNPwSq17A0RHLYPXDVK4PToQLqihJ58YJ
/3IR4Pthxx5vcFZblqtVc1U2YPE78w1YduRPsqHawjdDb5idjHj62ADQt6vifWiB
OOVrbyCWZoOJdG6Sootmm2G2gj0belFMbrjtFQOveAVq/WjFg55NZZEz+lvZtUGg
f4lkdiOWYEDBj0W0PJ4qm6G2nXraEdMdTK4ZKTws+QgPu1FXJY21/IXAZmZI+KYa
hDCMCaiiaWH0XXDfN19xLjcPlG3+aMGxj52fn7uIgchVPhO5bppGPUMALbR0lOAN
Iv/aXe11oISZQLtL438ZSRkaM4wAQXvAvDmEMNkRv4jOl550C/018EyiU5lIkDqi
f7sr9x69iK8XjmR08pXa63KE88qjosl458o7rdyGLeeiRei1Ve5rDPLdUbHH+dIw
MjbzfyW+wYLj32M9jL6CK0bNBPS2VtkdXz7317P+TLuR39rWYBzMhANKJElPhoDN
6PlM7aX/d0cwHcd/FLyAHMl5WQ/1NbXifUqZo6As+BVGJV+2E/FVfW8869+NvsY4
DFUJrOcB5NAkl1WD12b8G2syIUocobeVw4DnCZBMtG3E75sGhyNsyUdEgDW4ckLf
2rx8DXCPcnTkb6Cl/cbh3hUl8uhy36TYF56jwB0fDUQ/tW7BfelEqJNzcxNrsHM8
ld7uZQ/wZuD74dCC488bCG/ZyIAC7drjQg0ON9GVVon9ztHDQlVWUg5h/bJnifFI
mlxTjn+410rBZqY2+D9qUhdNpMjfOYKJ0oeXKRAiVbZRg5/BoiTRj8dJHNWWGl6t
WfUGl6VYA0Y5XdQXi0K4kN5QR+pEgQbXTBoXpwtVMKvNWyEHIxFJvNwb+gLKr1BR
IOVnv4bCSUti9mVK90cfQTcWu99hxxyXrwtE1D0MHVkgraVC9pmTMpo9do29b63S
OTSHozRQrjGyijLp3N4my+uzj7IQ/Pjo3H9E2udqmSrfZ0kixHcI+V+4sJxsJdEs
b4upooJuimoZuJ7OJCg6NQDfWs4h1E0bZsLvdPWFxo6tNXldaAZirU2OxTmG62Ro
oBaJAKdKHv/LdSPzd1cCvyiJN85ngYWoyzfhAFZbsDUxu74ZIUOsjLKaZTX87NJB
sTXiNiDMuWqT0HXe4Nh0tUHbcMcPlNZ4/ebmTqwNKP5bOTbATXukYN74DsIFZpV8
gODiShdUGGwuel+t1Co8RLW7P5Vn8p1aXY1w8hxOFA87r0JZ723bW0MgNEGm+Xhi
q11Tpw0dVKwgNFjvUsXVb1sSXQmx0dJ5FRr7SeZs+5Ou953AB4qxfki9xZ9W7oV/
LRqBMvc0XPUTgDegs59TIaYvXaCMQGbg8xzFO3kmwRL3WUpB+uoXyX1IuNypXDuG
GN3amOSR+ikUW0fgYP1KOfD7SjgIxcj6mMvaQi4oACEu2TuRwPTjpst8+m8H7zLF
eTjStDAoQNBSaGYwYBVfBFud4gDRWq+qZgQ6PKh+8ZnwwNYHgxyiL8H1dxC2Z7ej
d9Y442DU64UEhA0OEVKRp1HOGqpgMX6/XWWOz2Fj8hbeQgJDHbdWLEzpb933rk3n
jaA5CZorKAb3nuAaJYo+j5Ut5o6TIB5n0t6waYym9a98R8BpO3I6TiZ1ia6YNl3Q
FIZZ+0GsRJmzcX2207ozbZoXZ1k5nycZ9cGVDUWAkGhavJcMiS5eqpQe5hlyFOnW
tFcDVkt2mOx0E6aOfVTS1le2S0cLmTm1j/9A4jYMcJmFlEB38zd1izytPyZxEBLO
cv5P9b/59PbIsdNsw30S4htegZuJMKo98xU2Nb2ckuleeDoVSZzpLk+tC5rYA80f
Wi+zHIa6D6SZ12W9WLtnvXmBwfs7BrrKTcu7zzs9UAi6cYyGx/zmSx75aCfYaUju
RP6Wqog6aYhQbaec1hHYu7w7LG7qC0uQfZdOt9fWjuQuBm3EGkoFYWmCkH9VfOXI
drVmgpI1xszgzGALvCLRZiLPKC6tNO3EsB2KJRwjd6xlOvVp+4KV3l/7GW+TL2NH
c6bQ/WYu9RG8TFJMY7SNNliStdHQVlGI3x8uwYJtc+EUrV9q3YQFL0W2FKeL66+x
3CBNet/47rY4jywD/GG6y6JCdjF74wpmZJO7+s8pZ1Xl+I1e7cBXAGAtSfLoUFsq
j1/bFp+u2o2hZFGpj5n+0G5zJkMQW0oC0dFpsJ5RTLRQ92wy4mHVW54v+YTEyND1
cTQQOwCmjxQ5xLpZ6Gq1NnpT+stkQ3NBGm9yAtHuVpEGy1og02Ep7ZEw58FfFA4x
vTewaKm9pFRHtoxjUbtkVSQDvhG6JBVg6kgtbLRn2y+3mDceNQ+qpEohm9wcY7Wx
2ciHLUfE1OCJRHJ+4k3/MgCKE63jOTpRMelJ+L7iTzzWbUd1vhd3oUJScs+z7Hbw
WKhO/dsFePFaWhe6LH+G4o1L/d/aTeT65w++9IEog4Qvonusq018lXWnOAxmJpsu
bSwlgJr1eP+hRXvF63ocHv/Ru+ddMFvtRiPrmyDHcgi0ThbxMphS0PdigZvME0u+
0Jt21uFjI8tTWtSHbg9ullWFUbJy7TuJU1m58szzemF1DUJyj2RA/WtFUaqPh7EV
pgbUY7DLXon7S/zd7L+Z0EPEfH0VNfkHryn7wo76DAXuAcyOPy+1aHCefp5RuICZ
xRQapLiyVW6d9ZRwpS183UU6JGeb+zuSG3hy8UuiXBuil/LYQ4YP5bvfp7nKsyzT
XAEDC9RPTLbRtNvpnoTMkJUZkh2NYEA1i7BXmMaSQ2RmaQFtGv13fJVLfkBMFeDz
6iyEBOKT6ksEGTXXORqNlelD26GudjNlPCIE13aE/ieubR58QdKdkhIZgF9VPuna
T8VSWOZZp2ze/raQGuxiPImOEp7lc+79cfopNqZiejKQR+48DzMm2cFr480HU9wf
ETIGu/Io91h3LFC08SP1J2hWERZuihxvJ4+346caaD8zRDmjlzecVgEA+VvQXEJ5
LOFkGUcXLvF2v2hsFCSbZ/RnJ5ppGu42/f6dAHvTExmh0VZQLXsnqRkXZjhhe11W
kmZYk+DPQWMSQpFBBfkdAJCLdtv8la4ENXaDFQmXef8LmugR0dXVUNwhqrk7/cqf
jSlFWCuYWHyHSYJB5QTSocDiaNU8S9btHDy/L4WtgS53Dq8uTJgcUIlivkef9bWm
dlK/7IezPEM/vMByDJK9PI0ui6Pgxs/Tde6KYy0a+HAXC569RoZ+9+HN3gDPD+FO
ewUCitsqTM4eS55mQaP6nnpU7z/4bEiX2WhJSlQT1VugBihA7a53aN+YULYeYzhI
RKfVk0vlDnB1RvnUJQT0UyHgEBUzZQHPpD5FM9TAsh0jR9D1wwdh7lou5mbNqrLH
FpTYPVhT4N2dCSr96e3w/TvWP66KzQNkGGAb1M02H3eqei6EqyMzdGa+FFmdjLe0
3Ib152kBUoEHl2nInH4NO1swtcZ4ris93Rp6ELwp3WFHSVk/0ywhSQtHfDUl2QLm
3PBtBPFh7sjH7uG3eqqVsn3PhwM3P3pveb2nq9E7kRAPz3DDzEPQtbAkINoRajSj
J/wbqToR7ts0e7H6D6/IxQT8KBhY5sih99GC575bFpZFO8OC+EVsFB1dq/935FQl
656CHBeersKwyEJDViDuFDTxst46j1y16vlaoT94LgSe6mHRnWBW3OnPMPAbnyCR
BKqwb15DX+SqERgRXDdv2wT55d+am0rGKjtQY2wxY4hYCH+3ojpGHCa7eOgf2k0j
cu+J+koJjS3nRi/8AytPb6hlUFG+GS3FeS445H4VdZptPKOe9PUi84KPj22TgMJw
fXVgBrY5MEpo6e+qmJvj3Cq8lcugtMOQWKKDkgedo7Wj5PuQ6QbFpfT4dthbthyc
rpDgvEy3kr1gx7+CU/CMTci8Bs4zcVPXSQcp6DW7pLMeZoruezRUsVJ9Z1aJniq3
sjv0PjUrq6dRlRvQa418AGKJ97Fgt0cPe6cvFNR9NjvNw6KSH57sw/0jeTpZHNI4
J40rEi3V/NDXpOrVWyfOW2nvqsm/PBWcAddJq3oOHdUvLUAFRGOU3WDqVOJQrLvv
q9tBK6Enddk3E32JUrAc9ivFDxtK8H7QV2vNQY7e0EIp8h0w50NeDj7+OhUNmzWf
wtgBF+F5vaV5s3OuipnyUwRhYtMrPxbZllb53GkBX8jjMObR0KWJJmcUMIB+WJxx
XHXf4VV9y1MpgIwqeJao1bwg9NZwTyitpWBW41w8PflHNz+L3s6bkQD12IGG0Xxy
7pBzOHoR870AiTbHIWulY/jlYRO8ONiiBfkOnJb3Dl9TZ4jjK0lC9OOH9JVJKJhz
lgn2EG2NLParKGgHrBq0EkWj0fDWOaCnfygMwRUwhamNf6kYtGtqG40l4Z29R7Ob
8xiVSxU7980e0EWQqaDNXbSo76j3D6+mfdGAQocfud6i1vGXDNMZKDRt6AjC2Rwm
YWc9K7i9NwDsc6PJnYPzmHFSdD1gFxuSxt1uzD/E1qJfLFKYPpt24rGlgy5Gui5K
pVkXFrQoJnVMyPLFHhiXtjhPybS+A8rpFYPw3IXODchTBXYw9WtKPEilB5fONo6n
bX1nFhzf+4ET6eJWr36kxOa7wsfoFlABIdrkdyupokHWUp6fs+vLbnptfbk6TIfz
hgCw6x9uqM5Q3cnCharj6tqD0oBB6aqv8dJT0x33/ywuQA5SZMm9yrmf1ypRVDke
bOTnESznYZqtMM7VTkZAGD+jqsDeaN98tniTAfiigs0u1mWW3iG6O634Sh6mKCNg
ucAKmZGzUTMDz4y/SkQX2uote88AGy4Cv1dqbwEg/8EemIHHoACg1meJ6GYtD7H1
tG+i6FvVgYggx9mklZ5UPIAnJqsxFZQL2SoLAMo54TrsSWc01iJKrbAAm1EJHRnc
dH8eA18xhwQrTSMZCyuqRBgIhnKoVtCEz05PhWZqxjQOo+HJeWUgrAW6qPp3hKfo
G528AohOBJ0eiw6pfqGlzyH857pyAc481WExWFDmO8KOvVJtJO10g2YpGpQQHQPA
96aP7uDfSbTVH/kVmI3+TLa2tQ5fUQSCNlnaGdrdMy2cIav1tcQ/KlvS86c79EiJ
TETwmrY22rC0j5Q88C12pZaOBkb6UglsHbBmZ2L2SuGrbkH7orrob7TPh8G507pC
a26Qb0PdWr3TYWn9rimjPjulr4qjfdKrARRRFHOOoduLMuVAm0bvwhQArkZgZoRy
xRgyyM9TfvaHiERWMqnz39xc+R66aszTfVCFPQcdxBpwd7qRwMtTLbAQMTP+trYt
250q/RB/24BSEs0hSvyTA0GQnHBVW/qXidn0fG7n7OZfP3yWwKUpBlT/t742+wLf
4QIBXSLcVwk2KtM6rNRy1axsRL/lLSgRxjvWM3WoKACaqFmX56d7wE2CjjMrLaRY
G06IiWWH5cWLoA1CqT9L26ozwwuvu0d1vQ2eiUTiFKKgqiWw6ayX4vdry43jWwwv
DzMYxC7/EyTnUr/SFt4cOY7SFNkfalzp0kTtoTjdsr43BabkI37NamPbVWjxA4ak
+9E/jcRHBiYGxOjEV72JnlK/Nq27chbH/iRLJBxXShFTuh6VlOjSj/AxJeEjOQWq
LhHrmvehFDG2+QAW0pc4b8Ka1mE235FuKDi2IEJtCsJt8UVFBHyedx0lvTxypJMb
tuT32H4rmwcAkgWs7jZ6YCAx7IZ77lfyUSpdAblYa/fKtEffnTmf0C2dWLtwY9Df
154ZByjjLuNmMiXKJmNguatiZEQoEDw8nClZmkK6uddF9rpFO94TvtSD0cMBCFod
o1+wUAZ8srs5M8wdvKFD3JeZ77nf40cMoTK2Hv9sNAzjxBS+KdGlMxrMNeGv9XpQ
ixDMUOoxFxje0LntMWvHOo3Z4hFwDC5mnqm+yWOJkao5tNogyrnwaeVS2Sa6DH7F
JW7Wp3yQ1WQKhnZ3iS2NfhSwB6oue2fFeeb2pnYJQ3LcpRXnWvQSVMyFS/Qu96sd
M6Smr7anfcJxS9NdeaGp86T7lEh1jxCjWxEjZtwr1JojNSIlF1K2GffJs2yRt/Ko
jeL5Mejyw8FXQjjWjjj5/8JJqArznx/yboWcRk4c3qChzQmbC3TpeftptLfG/vy3
CpZtb+3uq/hNj0uUOCBdnNuNShZNcKmBvBeonmswAdhL/pyTnou8dTlkZBqoFqbo
MPIsFsrz8hf3QEdqDNZN2fjJC7tljoALQZY9R+GtZTMPosl09WCsWUracYm5Cn+T
Q9aUUr28k4Lpyjrlu/3Brb91WjsKn5MfqHH8WLZ6ekA8dBxtVZvr/2lIEmqh8ASl
iJWGLZSp3co+BFkAgUy1AFWcRp7RyuBdv5aLWgowPuIrjlDn2sfYUsr7alKkLXF3
Yke9JDpt7J0k6ThnX6i62kOyv2NaNiKvkPUMZ+fxm8aHtwFZxhnAMbNoOVUqCaMm
PsbDI6It7z+5+XxmMXqUqhROW3rygynTv3rY9ulSzx8Znsu9Q0/ce3/sXCQynRoa
DHdUGiC5euc0Lmn3VTsxiyojUJg1b2AxRZ2dn1Yw/8N6iEiDSzjfJkLJwZ47XWPV
eU0rwzkFh74in8m17YSviVD06lXFxs+zvCxG1dO5UEz09WeMeGyYKU1KzSvRfoos
5V+YmMnSoIXXSGRH59UrKEwg8K/F573vgKwZTx9ubuKLeqcSpwaZrWYq7uZXO+vZ
3b5GopP1Y4MoqlP5r4ZMNMIToGKA1/gvIaOKYUKyDpIb5poIDh9q7+J1G86MxhRO
CxpPQ5dFJ3vJgeUkYtF2mbwQ/Pq8b7jDCrEO9vt6sFNH1fNeRRisxyUCYorPbUpv
tL9lIUvAAZaM1BRwQ0LHFZGi0vcBSZY6/pDoGRKXjcYSzZ22cbdA39Ihc+tcB6tq
DjlY6lFgcGDcj26n3K75ifKMFOkVhfE5pJ00XjeljU5Gdlh4o7elayX69NUc3Cm7
J8jGNqKUBn2YMlZQTDPT5ZCmIkS2ALZHcUuUA/2ZSuwXCUTqLa+dwv0sEk+zU5Th
+7SV3/q02Uf8JDIELhhnmooVPfT4alghsif6qKHtuDPS6Gqy/z8GSovJP65ftyns
PyOuvA8v7+Roe0tUb4A2Cp2J3SctDxNidz6t7b9KbxFw3R7yJgEVtTKuGA3QIsR0
iWHjxMmbaU0w9thWmp1JHpa1X+Yi+yCqq2dIiFR+g2VRxPy4sAVOM0YawZ8kOHfY
3ALFjRAuAEF4UTG8DOJMCgK9gPZDQ30DlSG0egdSv6ZbGO+4X78YevRvlRz+Exvu
6xn8AQrTptrg101a+z2TqEZGiIlqxHQYmuWcmf0BvNIomPfx9Yh8IwpwQIXMKe+V
cBxM2hnKDe7tEDUUWsx22YLaTVJYw99gCRu6QZifc+/rszRi6sS9j5hG737NIqqV
QWZXyOAddkkksHjjUrDVEmv4xyiPFerLX2040Xe9H0T0Lkkwy7Cw8O7RMKaUzWd1
vl9e+mOS+KEgoybqE7YtbWGDjzQH8QXvjFTRO6pkWUpPe0TBWTr6LWm3k8HAnZwc
JK+x8NSNx2t1clLq3KeELyAutL754SbpcB6Dv0hqJifKlvjmJ1CDKsILzHKT+Cti
FGmnplK1eYB2DK6NX/NbpS883qWNITmeHEpo7VbgdlnpmNj7rzbiWCxLJvBL+GSW
PsOjcL3bQWJ9yMCW3Vt9tEWI6P6g/spaZsRStRSnldth2BMy/coPTUYUL41QzNgY
9FG9AaMSdDlfO/Bi3NlVUpUI3z8JuUd9SB3/LIp4fviXwL/Bdz9N6V3dKKeHUw6S
T9l4uowLa8u+i8WIchNO3CNRTFm29mYeud4RZrijvlZoDCxpA8cn+XraKNEfLWPT
MxUoOK65VauTXPlFVmAqYHeD6FJ1msFM2H5k6WMJvX+XnNr4HlK9ZEusrpT7mciu
lVZF658KJn5+wYfpnX/N5TIMLTNh/eSvY37BB5SCxg/Iw0VNHG0P2R5LR11h4dNR
XbHuqD5omGEyEsiPu3sIyIIuRsaBjY/fuCNE9V9opG1JAbWnzTJ4545gjKZNtkev
9LTr2xDj5iykyEQJ7YVn1oCqd7PM2SdeQBTA9fRsbQUIk7+eTqq2U75+fHv5+KXj
cd4gv5MAr0Xn+oNp5/xO3BOohUMkpnio5K6AxQTgi9D8hF7i2HPZFJiS4vtsevZc
Mb8v+624BxR4UPtgWZ1PXxAdfKLJkv+a5bce2prZ7mXKWh397PFTjghyX9eu7Yum
MQvBiUGBzKB25R3mI/OPs71ymkpLfj22TbmPu5ZWxuVjnTR5n/wPzrNXI3VroVbZ
zdrzxGlnC+HLUoMzOXZwCLHdyWluVcqIWL2U+prpHKUyskHUV1DTDC5FGD+WDZB6
GoI34M+Gw5208sZEju2txufAzuZO43m/UwjBL1fJyW7og8XGfS9H/XWyQJczyKKA
pJwEXMgtCtVWZ+UJ88+8y8BitzcBtn+DLp8CFDLg1LNEl2raqSzOymltG/T24gXR
EnF9EzV3Zbbx1zimBKVYuB9KUndeuXIRbv3KXsbo7VIU9ercUdGwxv+RGAa0ooa6
SuOgT8CDQnYXKIul1z/DU+u+Kf6iahDvLo2rxW7N1FcFBusZsH1eQGxiPkoKtRx7
p1/V2K7127n6GJUFgqJCoQlHAc236xCtqqNvATMVjl9pr6RSOpa4iFRfRv0xQT0A
Ksk/kB1HQlbkFPSTjPgTAkNSfzn/Z8x2YJ/38HyCSutdtUHRGnSL+u5xBxoY22dD
zZzgqD2csDj+k6fBfcjaJeQeS7LXgcj81gcz+YbdLzGudqw7AHRWeZhG0p4GE9Xa
9V3XT4U+Hcpr2Ux//dRq1H5YGAqFubjy8fg+/u0BTEhilZiLSrQhBS4WDdhYmuh6
5dFiqNY/niZ2eFjYUGwnHfnOmQXnb15f0Ij/PFM9zN9CLKtn68UVLBnaC3++QDIU
/gdNWiDd4GpSvYMzOA9j6wQnfGam7XqQsTd0gpNXPcetPZWrZ3hAp9DmSNQWZsGv
pqbSmcROLG3GVU1KPyITpT1SL36rmGvvs7m0OCiyE99XEFLGju81JwWWD63EPC13
whmlbIMC8djK0jpvF6436DRbamcFUp6CQ9rr+9Cua0DeSzNjyZvsSucbk+tOj2x6
qZgqbYR9S4xMV9Ljot16qKrn1HbFyCN/vG8WuSNhlxxcQZSEDOvIXimrTjasoGox
a524xoJEGqE8XKfwg3PBCGSjeW80xx79TznVz8JBZYA4qhZdzb+fflQOBT3TheSY
nQlL526bn9VobTVs4Ucv/V7ac6WCM3/4aODL0nSJi/KcyE3rX+KoAZOKJ/3gzGz4
Nl2V8lkJHFiZsNQEwxjF1e5yUP9jg+FTfoglxpRPlwh3Y74K7zMqFcsQpTqqz80t
SCUog3fvHMLmFoeaXBavv3FfEBUt3/RY8lRsSWtB/PPy0PZAybufHl4qHydJ7EYW
O3sCAJWrRhUM5+/y+qm21X6UdlS3kP8ACk+RhpT5XerKlyFc8k/PutQloGHmVAue
AoaBKk+a2hJB0TC+iavwxDjnlFz1Wapa9Sr9kRWAfid70iXzNv6txQjK2COwKMK5
IZgSaRCmTv9SkBwqJELvyB4lS9PW08DioLuXlgkq9WeDe6BmTn784N9mjJJCVcRQ
eeHoLEluuaHapo6Zc1MoZ3RHm9JSrGlSIUvYSeCutkNMEZ3Fpaz4tKwE+e6Xq7lE
jY/0tGYRQS8QTymJXxx13zGpITU8bdfCH438mxOwxp0GqRaFHr10h7sSALvenDXJ
a6GolqDnh38TMktQCERHwVIyQ6E1ep3G2jBiJpxzbO8NG4hK0YXOlpcznZncLhp8
ImYEfcOJkFTPPOKeSVYdP7Etc/iRaqNiuGIQA/zbKG57IqjxEBQIX0ZAWGtQR1vt
KpfWugdtwT7hKmoz06T+FvcSAHB/PEW3iLHWP6LF2cgvFtro0IRJmRa4xXJLvo9Z
2VxOkqtQw6BDdETmKKTA+PWSxwTFUH8uOmaACSgOv3I+4rMfcBcVl+ajJwRKoOW5
EzVXfNISF2q++29lZjK7/R+CvYfQ3G8pcKLu7W/1AGGTaN6PN1LR8I6kX0igEiEp
EJx2lJ8MKrB8SqkggC3SO4BnN0iJ/7PWje7dj5iUucNf6dzD3FKZG1yDFjO+pN9B
5x3rsk6pvaZDwtqquq73qJC4dJjb4txFPhE1WPye24ucKvLNQzGVgT+T4YsaYQKf
Q8V9Xsu3YhVJIxEvl3s/6dEhbtweArgKuNgz9UKs8ZYIFSRU/ric9N7omv1BOBLi
bh624sCs5Tv4X+u8ifo/O+IvHmgmaZ54Oi4XoCvWKoq9c4ol58M59dvnXGdzwPiG
TIn5J0/6hkf2BAdSPq1xBHp1LapBOT67kxaqP6SIymUaTgq3DSIgThCOQBzINP/0
7cT6qP5h/kCMPsV8u2g+CatxwhUVYEM9XiRPqAXO+C3InAqOltGh+4XDo1mYzROe
vtU/5tn3csTmp9FCelvxefpKYczGCv/C+O6a2+CzCctmOS0MYOXyp/x55hVmhzZg
3E3NexmQBwd5X7zh2Rtqdcf2lzw4SBb8Ik5t0H2PJysYgbvX99Dv76WkZImJ/qo+
cRVfJkbHXdc/J2FK+ZA3OxUL9KJb9CU1MPb20KMaN4LwbUYgPqYqeG4W03REgQJt
Q1cB2iyQ65o26foYPRI+kYxjJTRXaMdUehIoEyFJS8nnBaD3h4XUEpVU45ldi+Yc
WWuej4OSC13rY5FPE1rBc7wRAEQWrAU/2CntVQnu51JNAAvNvKjVfgaeG2wKT0b1
BhEsCZHJNWRAb+nPVQABR2IaybmTErmiBMq3JeE/KaAuCzQOxM3CaMQdS+3gtfJJ
U3erlgNW4aMrDY0H5oaUm0eGtLTEDTvZPY1TSY7bsxCxxfdfd1orQzGYzHvBUoZ4
HFOrxJtS6s9Siahhhgyck0aKHKxOkwBWmttVJ7IMGxKQY7NcjyBd230BzaZ2VJl7
adoa8f3j62ongMnXbfsRSi1OA4mTb9W84LDwbcVGBwzje71Gp1AXRVJtq9G79ioY
eks5YSivW0kPQjXtMDqr6ikLwnDGHyEQSiqIjSHeS94Ua+u2Gyz6BaxLpqucBJ9E
VtKprLBDLzJfxFm7AFdDI2+d7r/SQRsFVz8Utz9T8ysKiynHpC6yp7I8f3peZ+KK
nCyXcsVS9TkAs3B3yELhpX8Yu227n/osP3V0i4DW1293P0JRmNItaVI/myIm1LyN
+94VX3eq/1q+xPOrl30QWVufavRaorrH7yt2ZghydPU7I3uyTFcVGElAJRdoiqm2
G5LnWwpqWN+gCF19Gaeb0fbg3uOIRHhZwdVvfAYnCegnIRdyZgR7PHWCq1tdbawV
bayLLlVv862XdLhFZA9KY5hM5d2DPp8cMpjdRM6DHlHZNqBpJLBfkpw8TBfW/F2s
a0N0PFiF/lbPJFS/WlITo/GkHW5nJescwJPpGioGEIG7HGBLSkU3NDC8+K2Ndu1t
Skd9heuJ6R0w2qI1tN9yWxjfo80TZkIqw5Xn8u48YvVf9mtXFDUsN01Ti2O40+6r
4iqKVeyf+cNhPdjlOX+FLCkNAmU/JQdc+ELuTN8KiVRnvWCJAG+Uu0b2/1nz4t8O
EsPMK2ohsCuuimy/XIZ0pqZMkfD0MXG9Kkypxdl7ilFP66ebX3paKxU7L+uPllU9
6CfqBfgnSdiw0R8TUjGrBiZIAytvfwYmxkwRQKWNIpFSpKATUzV6MwzrBYlhq9uw
zTz9331eQINgkCy1YJMFufbVlwIxRWLeH/zo1BZzDw+U0VyexyJSt2pYppoOMKYb
skaKDqgl9eFr5yiql0RoQ8xgGPC5CW5GPz7G1cpyNQb+LVqQozRO608+Ue9aN7H5
GXhF6Ez2EbRbHAiZ8uwSh6u6qUWHEIjYBFKnoKBBYq8+u3InwsPwyfK7sUkwAOBZ
wW8ae/KHEqZK5rNJ/B7a5sezo0MWSTGieFEgiqz5Lq0qZAcUJmceMSHJnvmy9vGl
RgXVKhnq4lqR6ERxqwA7irw6yq+yeGAimP0AeDnZoNm6VJ0UX+sNjZ0Bb7+4kijp
nhTWSuNyuHXIh0pEnfAvFG38TzNOcCwAGw+m2pQOOuK+UZ2JAw3/10w8qf8WvXG0
wegMk6ft3qqk2JvKr1YnuVWY4y/miEsFXXvmq4oPL0RtflZYIugi5/nGzPQ5M5hj
AeitRKTIdqASPU7vEYrjnCScC+CEv5FtdwwC22vqA5it39DSM8V7/kEcIg6avMQR
GAm82la9iyLTXErF2sn32jWCvUcNGomfhFkz4TkOT/iQJbqsREmMOGHC7XJvo5bT
1IsTre5xx9Ji+4xu8tlFuzCPcqC9ZQHpJVDbf2Ej0kouT7T5GE0Df4e7kne1/9jJ
eevQT4E8jbyFP9zO/Di0OfSdeu3QLudzA0bb9WCQrSuOINjCjhv+BKikmBxCQVP2
Ybjh/kzD+0b/B5eCXQyO0Q5Z6OAaIRzshpnzgs53NehH9cS+63yZL2Lm939dq29f
2HzPzNCQxHMaKFDqLTlYiikCJKPE//EyXlZsOe/oaiv7RI/WpAnP+id70Y1wjwbI
yHiV1YhgLwVhbeAgwenAiJF/nCj7B5VC22Ps4vhv0FTIR8RO5IAFBuk8nYqnwT2m
BRFCoA8fT1o4W040kaSqBaKINirGHmo3gp8TDvIkqM7wRQx+LkwtBS2+QKUCWxPo
2zp6JHxNLeZEdxnMubgC9trt00z9F3icYrlN3+47G56I799Qf7PjsxXE3m/U0DRq
B+dpRVDKPzdqR43uSsQNKW7chz4Q+cn2PXxQbxwc9rKhv9LAMcVvreuvCdtYyblO
eaRaVoy+DTWVBJwwZMyoJ7iYJ/JJzyu+sqNHA4bJvPTPrpOqRPM7SXd1NvJZ/NpE
dxoGW07SHNeenKbz4pWGJG5OWLtYynHh0Xh0B+dn9u5zUy/9+xr7Bku3sY/wuQO6
pO2h7XsMojnrIfLEgWBxT7JZRjsWVssEsVr462yuIZEfv3AbVLtHZiTPgKvchm23
6G0HDRJd0r0bjYoy6QU2Dt6ywm/Vll/nINoO6MUsEKbg8SQ0hI2M61wzGcxl6Gjh
1fZsasO0VAshSJBmo09sQiFuG/GTwKdigr2KqBF0GnAiF1Fv6Rb0tAQ6vFOxvZKw
x2h3sGq9tFrjnj5dOen2advxn9crghJKr4TGR7zuS4Ry6tqN1yOh6tegwY6tnOYc
r0lahG3hvyYFShtQQsch2sRbkqaIFp+QE1fi/rpD0TpeoOPKhPlpch/35i7CUPcb
5mLpaN2ndJhzjMDv0guLCGkjKoOfS7TMNkjOjT/dE57xCnCHReYItbQSdKe7ib2j
K8xqrCmQTyFC/5NDLThS6frl5TtuLHDUP/siRLVesN70yjsUfgGgiBNv+EqpRIHr
mjDSjXC2lOEaQSYmS/6/SUQkJ9fXXaNlGb195TRPDauZ8qAKerHCzZQZZ67YdOzp
XtDz7BSsjLVrYXy1OWjpuCr+te6IS/NwGXhdWekqnl6k8VnSGL5sViYnv+1cJou9
aJgTmBm5rleLJu8y+qBK7opHSwyisnUkJJYABafgLicfdS7c9tjjpTes58vBmaBz
D9JZHRRZ3vpjTKQOQ+ha3+z1ivYue6zriszh5yZEayCCssD81UWyZGkoB3msGOQi
Hb51tWc4VBai18VGQjf4jEQmjC7rTvlYjGmSTp7zOuLfhdrYgkRb2rwkVacY4jzw
35kzg2Xf6sdGXHgsoMa3UBh7GA4oOKFLhJ1s/IETu++uY9p+/6aJcDCqey8AbI+F
hSOVdIl9uULsJhVoj0LFNEdZ6CUrDDbo25BUC22qFdoVGkCtu1dLe/S17zLI1vWj
k59l87MrA7csqhSkyC1fq6FtmodGbYoqN3lIx1b/XhcKsFPALxSWEnWHcD0lnucT
5ftca6g/rC9LDBUik1jLDs6/5S/0ck/f6ASuYtEV34moaXvKbggdbaS6sriAO9+I
AqxTJB1VvhrGymZ0ng99lx9gkgDRkkHC6O9rt7/GVmKNm/Ao0JTiSSRA8cD4tnav
IgyWnEoRMb8hUwfuboKK+xgWhVYWTzRigaPbMNsKPsWYJL3Rkjz10zHV1ctaImWI
1o6s3tL4/Ms2bRY5A7vEpz5IUYoXLzdENL1GzZ/5rqOZ6wmOZcuZfjd1QLP/NnWV
/o5WeQmgSS9BwiocqAq0R0NvbaX5j6JANz7H29BBbsbPzvHeaL2P9kLxZTaIHPZE
XFpRVRsnSpkf6eGgl2TERLKJ3b9fhEmu7UWzVllHjmwibJrxf8hO74VEeQGLVPn0
jVb0SUyIXVkFHuk5ZigD0RIL43L98t8EXrx3UCvfOixuYSlqcO2llfw75qNDUua+
HQwrl3BxMhrZHITHn11WGNx3uIm3Gsw4GZXJCsciTjanGdEPwfAxyLfmsJGpdqIb
T5cezG04LkfJDPrTWZQWodfPkKQPcVxPTqeA7pxO17A92TX0IU4/buMJUkzRSiEy
opuVn+l/BTVcHJaKkA7TCyAnux90NwtE2lY7vc5J0qASMy3WkbP45CIxW/lNEIY+
7+w8c505Ep1Sp2TDTCn+t2kctGuFBzb+kM2JTssWFYbmSBE2STGSH3QLbnF/Gki+
5mNkQ20qf1jJ60d1tuSMtPhtWkgpcAKavN0N4ORVx4IgMgodEhRrqDMMgqh+USbm
zpqsmOsaG6kBXsfVTvM7XfkS7G6WELmUi4W5NoPf+J7Au/nrs9+IrHMdnyWpQbeo
pjurRKAQRqT9haMMFImXkjNnX2zKQFolpMi002I9zh/gVr3HvxcdhfmBx5fMqQS/
QMeGq3gO5K60Yod6TboIAQ4tKZ5Ya2WXfQ4DTqkIpWGxcPOU4YUIPaXpN2fWzlth
iP9jCSPuY9I+l6u0R+BQK4+swqDx0/0iYOdEU2gKiHY5RpfwhvGklAgfQo+WsL8K
W9JNVgHs4dtQ6qrqRqdMJ/RnRWS2yasoMK53h9AAnghbvI8Dp3JSInO1f3dkReni
gwSg3bJsZmjKEMr7hfPAWFHo1Fb7tdpH3P3D0N/i9I68a9uMqvZzctO8T2h1SAW4
uUXCyzbpq2AQaHHctbsHNlBvvRPPG9xoLxzEyMrgLdPL5BHLY8POv2s1KG1aR+sA
TdweXb46YNMFzxAck7Yzv674r29unxVP0zhxPX110ka6+IHpuDiB1F+y421KbY1c
LJ1sIpX9KxcR94428pJsZ+zNjOtiqDIeE2O/drYZLVPgp8ekOM1xFJtpQqQNF4am
Y0Q5czFu00sj4nxqso94Rtkx/jlh8sTasDqEygl4N9IEYc9ZnA2+cLZIEZmX9KLA
uRb3Bio2VyEnfeb0rtkmr0t/7ZUed14hVQ8WaBoZZzYZWaH0NZnx89WOKdUXhYVs
KXmjfCtvZTECuqZQF55iRXrc+PojjiBH9ZRVdCb+101ZY6Ydn/t4txySVaeH+Fni
M98Kag/lODjZCT2Z98ZtQWawiRBYFgGCvgq6H3RRnSUCPAwuLjrAQJtOzS9pnQZc
nS5eZGtUADIXQ8pH/+wx49FGn6Evbmj31TwF4u+K9Y1KMUZATjvbK8DYaLHiY63c
FY4pZql8Ci/HDcc+hBXlyJ1L7k1UD/VE6L++m8sBx8I8UwxUPsWpc4Kyd97kFzDC
A/L+2URqrYRvVUI4ONboRDMn0jfRFJi/W3SLIhPortilHs7C9JoB1DIFVafiblzx
tMvm/5W/reYUlnCWOG/MvL7RonH6S/trrYnDS0pa5WUOesW+xy7JPOdtFKxNtCt0
tUS2hn75rtRzaPJry9ntMj9MeaLYHjaXDjb9AY3ZJYCSyqMfVUV2p2j+eIbg+rbO
il8pCgcVngZ1RP10ujYGkZm08wwyjNEGQYvZ0PuNOxNBXoZFwzxxoGuYnryL1LPj
1ro3Po0Dmn+o1Mk6BrOxh2tKeOnsg1OL0DvXsMvsOabho1zWZzn+PUIl3F2LfN8d
p2PrhEe1xGhwR8DUrx019LyNLt1AlUTf+sB8RanA5bFH1RhxkdEZRpjmST2Ua7fk
XKLAgHqyhaaAYZnmZU3QWY+LJK/47gKqp/Jh15fWMCH7h9K1gYuW2stimXCNqaTM
lVJ+pcg00kKJwH5K//GLiy9VQC8OOmx/gRHThlISLrysAvDBz+nOYJcF3hFwVIim
jgQMomhk0e3zFLHZ5my7uQcqiC4LEPC/DL32sXfH2fWvxbhw7a2BFYxckxOEdYjO
uCowKmegmUMJUvWHLL6Bm3JCT1z+0gvg/K9Gy9+7GL3k8KWd3CiwETco9KGUMAnh
/9KVxXbUkwNjo3Zh05w42igeNW11cobkIICEXArVGAqnYTVdKHuzaq57eKzoKqc9
G1etjyhP/CQl6sYVH5ttnshIqQIj32mfx0AeVBv/kz4sg7PjKIvAH0+qJfzeQLjN
uirfzlbE1VXJh3AWOFp5OlFHxzIJ5F2LKTRfUC9nbOLVxlXcDZPpLjTLPv0nbO6p
7gb968y2gr5QJUxucwXPE0940J9c8bv1fVkDgeuflIK/ydruDVyGSWALUYq75ynx
+K0wymJmM+1d8lmoThvRldoAQO2CICQCuW9EebWj8jXABhImkmSFkWrsKh/hedsP
oF6epx566TQxsLnBQq4u8EWVGWupBzSGJjEIDloNE+3tu2rnv2m/s/CQjfiLcRHJ
5kNharnlebAUscuJOS6zV0tt9rOQaJP3e1WWwo0kwvlXYoN2oPLITNEoYOolBI6q
6olmpZi6j+CC6eVwq1SmIQnRz/OGZEH9kPjxjsoiez97xmG6ry3GD3MgZsO7GGz0
8DM2tuHK9GMGWJQ8yDKfzvKWzVu+4NHUzCBFu1Ps0g8zAj07KyxzOl0J7UuMojz8
qUh1gBGlNnXxF5wD/wKFVIEk88r8EAhYjA/m0REWlT8KvwUhmjJPL5aU/gzkImIG
LXSmQqTDe5fBKmY72f3XTXLopuKmRn8lV0/6u312peQ9PvWuLcdPmMH5ptcnbu89
oO+2YWn45KIjjlVyYFGaiiSXOtQFEl2iL7CCTTukntXNU/MTy7NYMoIpP9yQYx0w
4+tE4T8ksbyTiWatkNai94/uWVNUYnQzmyg7MVR06etyxUkuF6eR99rSGyXnl245
h9tzQRqg9H/qk2wTuqrCOWoVjvZARbbyjcrvMocEnpwt8FJ4BPLHfHlRPn5+ZFKo
04q44Sj65ZOYTGOMGXrujwf8Fw9Q7PPTrzQGz1uT3+vEopnEF3e3MOBKWW6lS1Kt
A31Q4/tTNepoyN9BS1Xh7MyBkZO+amJkIZJ3eR+z4PYh89JKLs64EtF6zCq6H5kr
EpqK5An1wfrQwttOHBWK/560YqQchqk8VWatCaMXoCigWwbhEP0Fw/U/QlOTHMYD
Blqxa8oXqjm0y5F3eFfe4fUCeaO2uo7aoh1DuUc3lyJgX+lKnf1+tn3DjRx207h7
INahdxT7Qs7zi3QUQgyQjPLzLLaBd1RfgaYWpNPqtc6n854n3yDtBtGn41VNzeFh
368Q1RzMR0h6FekqjxCjrcnpITAdm2v9g5dhAo3xy+sdaeYUpY3ma9sEYHVvJdiY
SaHRNHQlTDafj6UMoLsS23yMjZwfBmPE0baR0FFGnR8XiWGwCscIVyEAYql2X0Pm
Fz1gaP9xHz1yXkWtgfnHKpIDyIiF0ks22nsL4S8qqD5V3CgKBxfEPplqqQqMDOMp
iT+hileMpqbCAlY4wuQRu1GVlUw94lAVN+0BvQCGpVUvDBU4ykoxJIzCojLccUVQ
tlZxhfCWpnW6eR+iurfeA/OyvNiHU5YEkMkpxqs5fTZNf6uDh73yzYUWdTAfHliT
cuYgJTN89H96NWN795lYxzVy9qa+yRSavWb3RSu9UGU6xPf4CPSpXhELnKRNBk6q
glowKg+izPlIGETLgdF0fkIeg8BfXRmmewXoKwWX4nI0Ds46jSvC7u87KJg8VtU9
7dwSsDuW9hYRL6qz0IQhlr1d4T8jJau0qnQR5jtAGjWB28LzaLXh1qrXJ/1kaEcl
/saVBX8iRI6OhqLUA4ZyNXtKu/fhF/Be5XymJGFZryVN6h+vgDVnCDLDWVuWkAuF
fDgYj0nqxM8DkcvIB9LGunvlLRXNZb8c12+mxXkmPmi16GOohdTR6zt4wtpSoE27
hTt98y6QZGnCoZloKSlic3ksSDwrz92wl+59h7jsl6xPzU2Beqb0/sdfGd8Y6Hux
ZtqT18JZjeZC2X9ZVWr94K/ENF5fzaGgVrMjzVRe2bA2GTHsKwVQ+3ZVsFMBPZB7
8gco0Faw353tOz3RKobEE4HgMk1XHQBgNIZrthB+Ag8FfqewFM/1yIzAS3DtGbmj
0TMcETeluvX30K2+dveD7XlFc0VoI5MpapcaoPH0Nm3G6wsXex5zI/BduaTWHDT9
CMxSQlVXVPwxY03gw8VDhiTDRcXcFx2GN6nVlHxVvMTaJb0N3NWtzKUKfM5k1KZe
mng3/E16jJgdjHF8w91+5G1C+u8FdrZZDVwkV3Ba5IzYsGDRz+3L99AV7V+8E7Ql
wzuFvuOghiwXz/tKsbLdQpDSQ1ugND2pW9TcgMJuV5/ofkxTMRto32fhXLSWoM8/
OeGoPjC33dlVclr8K2rvyUA5nk3qzcIWbyzuJ+HRdw3CMWhC3xwY7kUQ3Rk2qdhV
uK4z6r2x0E4Rixj1LOfAFj+H95YP8RItrBHVw44c0HxreSBBLoQT3qd5PXLKuHIj
mRGtUN+Jywe12f56rRMrakBehWuVbDl4sqe1nWDu5r7on9qcaIa9Nh8yxA0dLiaZ
IKNDkKAg80B6B3NebS65b5BI8a3aTbWMA9VHODRpkXLoh4f4IlCiaVDX9JZe2ya5
D4cYIPhUW/d5hnOkbSYzaw4TnBEZV2r2L2SDjZ9dHhM6WbkbNVbUnKZynmcnNSCS
ZiE5yXYQFMn8NSXnvceAehKrLHlu1YE94rp7rZoC8S+pvNxu64lyS8/5MB6UrkpI
IDM5FMoAkz69dPTNZPor+j9C6qhqLCvY63TSa9J+pjTe+GZEp4oXfMFysE1bp0Xf
IghX/B6RRUrXZuTB9gHe1l4M9EjyachLUOf2RmKRADq3d6lWmQUKkfP8dM9GAODo
9+fymq/Pkp6fpIZGYTbUjZFQYS1jLjgJeRGzxQHRy+Qh5NwWjC9DJQnQ8Ggq8Wd+
quaIUJeL46UfIcCg7KKK5KOJPcGCOTe2NeCKSaUnT00rxo5hFFLO2coHnhnYZ1eR
ahXFMvu0EAldQLioze5uv1VCAVqPrZWqLUkNP/+QsyVg9K8eFFc0uuVT9oa7+vtv
hnkAowX3ygTtQhkSSdWDXcMhETqHKmGEhJhBeWcfoi4IatgIU/VO6gg8u8aE704O
5S4mbUYFIUO+YghOuNQfz8ptxV/NgKWJA0W4vc23BVufFUVcsFqQVBSF9bkGnsJs
Jv+ftf6jr93Qre+seM3oL10f/yslthgOSKrXircx0V7PN+tOiDNR+vFIzk1n8Sfo
RRq/QLy2qM1+ZAdSdlEShOsNTg1IDP9hLL03aRtGHCQDeGwpRQvf0EMP+3p0I8yx
/zNL7qea4uAG7rUa48ZAugykn06l27ocOROpdZrL2YF/jMRzOfPU/R0Nh+PpCQFv
bNcdIjp0loim3BsxQj4ugVdXkE3mov3ihB3iRgrUmXSpvTO7750OfxHl9nfaL6Fy
FWzDf9oLT5K32N6/HsHaUWM8Un5BHD8WVXeVVNY+s5BACgXrnBDQxaGYJKayV9Tn
bgqgNa6cJ5uzU/gcbCn+At4v5NeFRjGN7WBtCrJYcTr8/ucytIz/jF/064eagspO
eoMj6yQOpeNcVExyaStiWCi7p5X8Iqc/ZZGzCQ8RDUBuCvJZXdo85E6kTQYX16Y+
0meSkNOGjMH8Fiq77G8/C8XnSLP4aDcC22tRC896sYT46l18hx2gow1NB8p5N0lQ
NxiIoMRwcCn4l8SouQbW0fqCJb17QiD67q2QhOFhUF12NLaN0HVkgMKuDjebLuV0
HdN3DM86hsH+CU00Jrg78xIpHdaBhcAEd+lgcbDe/BA0yI7aKG+YxuKpWnTx+2tl
A5ae7M/0Wi8UEqSKzyxpjnWubqabA8UkLEXVVwifOMdyR1FyHxNTpmjiPWSY+cGH
tbVLoPygO7PiVCLTw1BPllmwycSzQvN5ABuOFObkaRQ7dhBZbkgfMeKx2XOoV6f2
39DdxIzta3dbqsOIY0wB8q0yPyWGntg8HKyHZR1Y/T+0Q5+rIObqkvaiIKSqCJwt
nmyIJrtZLZy4QN6RM9BrkrirerOh5kMEE/RC85B6U8+UnkVJqfFAMbjEdr8VKgGS
NPuquVk02RiQu1MA79g6TRnWxNfWGwc1RguOU8Kf3BUOcGlXf7gQMyE/FRXHNbHk
w9g3eWKFE7Da5U3BeE+VyQ==
`protect END_PROTECTED