-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NPS/vvROXFap0y1lDehYDvP3ZcSuKVeGx7e9iDvTOE/BX091aQzk9XuwGmqflsLSIhv+mgAmDT54
WdX8VRPsKFj0UyxCjorycAMp7fmiG+ouzS3GB4UqUPTFwl1Txqyiz9hbIohiWYsCOtX10rR70B1R
FuAWElvKTwEl/qFCakimStsZvMFE98QDaK7/2FjUZbONTgZI0M9RfJW66P1SSsiNrcK8fZpBdNmc
5ok6d3DQ9JHR1+mw9w6D/E09WXV7xlwPNQb5Ym5NgnBWxjP53Rb9oq6w8U7m4tNPYb7bbw2gPfR8
05NT67FbpxvDIQhN9e9ajp+UMvT6fz9JahWVCw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
Iet3BniegKkZxPueejKWSFskDqCLzLdi3KEydXHK9pljx5nSv8+he1rCL67qlhLaM1YIyWzGpUxw
CNvy01eDIGFCNObNtck3In2KIWAHCKMbeTmYouK4mMxyQEHQdBNcxCRNCvXpJwXs9uENTL1qX15p
i0KchMK7g2ixAdyvDmPO7BlER88ztEmGLgJKCm5MGPzvUsOZcBpi3oqkDfLRTDxXaR2HfWHndobV
65tv+JAf6JEgSQ6K1s3GqvHdLEpH7uG79ZOX2mTsoqTc/MpeeFEExmVAVYv8giMc2zVRTgHmYKoe
6IZWlBAofRm4m5VjJraRNXs0psqeo52QgwwpGswHagOJP2YXqi9xDv8KVPRSeAP5OGpJ5wdAdLRV
rZTkBUkSJUR+Yl5FuTS8IoteVWoXPtTwQxGbvlAHjcsy/BxH0I4mAh4YGxoOwC5sfXo+K0mXj96f
yOKYYtrB/C5v8NvmjQCXzkXM1OVWvFVwto6hG2qsL2nFWMXMxygHVQydlY+vDxJZ1jx89ZFPeJ2m
o/qb7mtcUmPzVaAVU00bAXusPAm6hz6EZr7JWS8X+E0vGCuraN0F8dqv3wT5vUO/2vYM6r6Hqh1E
XznwUtdbDtSatEevFX4qRZ1Q14H2ZlAxpuuMwGiMqQH7afVfvDzPZ7R2fmE+q+kH8zVnDp3InGrF
yRt10qb8AZWKbeDf1KMsABQTBFFY41mexriSii9QK/jwXyffL3ic5Po+uWTE+iY4jPxb7T9F8Zq4
ZEGPSZVaAYfG5opvVp2rrLdzrHNsLI/rhrBiLkqRzKMsSjYF4EAKfMiz0IMjZAx40Iq+ADXDoRM2
3y8UEv9l1IHpYwSD4gX0YVGOVi9gJu1vYSMQQvXA+lx7YSWN8xuqLM2Lgx4fYVn49EF/eHrGnOPJ
RhxMmNU31VEdi9XKb9BA4yPf+VZQsD0zqBg6Iq59YgcDm89qpNcyiooSw0kUcRBCDsL/zzojtEmn
ZSjNQGCuyv0+GxLPSIUjKk/OMSa6juAjyzlmM2Jfcm6CU4cTsrALpNhYUsg+8JQ9YUWupJ7ZOCkr
JytoeUnfGobmKSpnscwlY2m3nGPQXA1APxVEi4I4qPhhEj4xqEESfYEZL7Ozfd9FutqMN9p5Y/0J
Hu4OOZ3nWa1/EJrgyzObFPvuDZH7cEeC9twjm4P2c1XCUjBKdO/txINsXM1CIm7rRt5SWwimboam
FcnKhjdXoghH3geDx57ZEGwxIkdJUnRu1DBh7V/690MrKU3yk9agnHjK5uIgbrKR+s8y7254aExO
jFhDggl9QZp7uz8tIa84gM4oPqgq05tN3D9I2uaalK+2ia1YVQJnf3OOugvxrg+KykqA2tHWRdhC
nzSvIDH4pYDkqZRVlXQmBk4A+l72QMW2q4GtsisS4jxhJvY5z1WdD4laaoH87cyHhfAgCBuJ9kg/
iMVz6quiIx5XIxJk+p29LDodrog1ckZrhqsK8dRTjjv1jEqWUdIqUAIsP6yts5YvuZZM2VSeu/Zm
rUmM5XodPP7Cv11E83XNL27M7z/CUxgHKs4Jnwx6eQYdYt1ZSzN8lCjDzT7aO6L03NcIvygr8rfE
3YzSZs/dLKBszhOC5PfsrlZsUVwRgcNX7Ybde6iKelBtSxQZUKjayxFzVnUKe0F2CcFhQRBSdx4B
Qz72CPUf3T1vq/EZq7+Kix/HA4GemrSgNxt1N0GaON4BynzQz+X2nlfDdxj28WEOIygbwcJz7p9Z
h/S06A5vblfhZi/PqLltOAF186HN3KZEU22elu/N7xWlklfXxLNJlIhd7fy2Vn3QY+kSUSRECvuT
IL0XbgTfa0qKcl5VgpIE/iw+AITBt90aUPos45bwb/6q3AyVZo54eMEBH5Uko1C5ac4weIMpEBd5
3bpSgXZ6o0+DaOqnWjsKwWaUyl2zN7iDlw51bLvATG5IcxBEB0EbuL6xVOhux6FeTSOFfN4dQvtk
2nF2o57gcvQ/FiLzH2nX8LhFYnIIv4kawhFz5wE58ianEMBUM9nESNyxLBxrCMjLoGY3CxvqLVoJ
w3OwvMiq1cbDuPl3cdusZqhEcQ+Y4eMdCvkwU7XpZZG+DD+WsqE7lXcUnnDXwdgAeRheYmBEDLKz
cQGSZi48WHqrtQ8DvAKHOZmFmjEShr0Nkhzc3koE7CVzfgz9LDO1c3BVKI9l9upBwyQ7QHFS7A/X
aELcs/f6PcRhgnmJFNs10A0H/gVE/TIvORwcH0+mtWd4md5MggQA9doUwPHGgflLAe1+FssAUUy/
zI5b37rLJufSLGeQH5d2qrxFwCxLgGXL7b3vxta9KHTxy0WpUCvjmDjcQtc9eDlkodBGg/pSm/j+
wRJnOnI1GDTf0ttXZKlKS4MzMwkAJ+TuuVNYtie1lGLBj0MclOJj4TkIn9pSbvevYq0coH/+tByj
R04zbIE8E6o+cVbWjVwhzGPYmB6+OiXpef8FXnMcAbES+AV14iuMsKogaJEKtlfJjpFTyY8M61qp
Z359Kt2Plk0jFmoxXnMIDA+Ze91X+hbVNC9Q+lLxBbVdSxXLBeabTJyYt7Y0JiHq9yvjrDJYR58N
taancwxfOabMhuS/5GzW06BDtJvB0FSju0hiLSB+LbL5gCPKoixc8EtXFJQu7oAeTTPtiOZ7oYUh
7CIBNHRzif+2u740p4atKWHOQfSkIuOOYwMB7AvdTYuNelbzAliZAWCZLCilMOemyZNkEz8z6cZi
7zvL/kYZI2bS9fWtuOQKo9Rn35XUCc5cfE+UnsSV0gGPkPyJItsAeCJfFr0M5bwhRcpjSdwCpTTS
at6+tVWur3FlTDDChZvaEvDm1nI6QzG4kuJohTAmSo7ugrNrB6/NnlEAmcKAQw6mhH64ZW44pGm/
BqiRCYxhaD3jeAC3cRXIJ24Qu6Rdn+l2KtCjaHtmoil7mRIT6FLCRU4HgTrROpKb2B3zcN7mveEo
MdrIIjs/co3VZ7M3O3LbkBjOtLjf0SC3cKZZckN65dmMOG6ssNf/7BhVdHXnb/nKnzAvszfE/IWN
lPHkOVHUfr5ZEZMXlp+ClFwkQ1KT9SxMAKzJFwRvmbghTrQ3OZibeX/WwyRrkyDQD+7AoMieYPUn
Dym5T5CXvVrQp54OFCaqxLTcvgqLt7iIcZyG/BUOJman3iiyMZx1a7QSljBrwEsoS0vV2l4zziw8
NwIHNkt4vlxMKQkqef+v/j07xd/ik5D2WaZi8aEtkF9TZDFmHQ3RjXZJm72rFkrdQE2di58ISFIP
pGCyxdqHg+QjHIvZsO1qyWR7CCIY5EjRyEYE5jLJbCEwalb0LFoaYWOA84mBosrIIPmc/jpqp/rs
ZN9wpTUDBdi3n1zhkhz8/HWTGzR3V4I530GWVcfKKnULBZWFUeSN9VNmZ5bdlEOLnd87kt8WQghh
TttWVQSVrrIolhAC5T5ok1EuSnRnPNfATFSR9jX/xqlcbpAxtT5vmYshruiLyiZk3DqRII0t3jar
5T6y0oDaxegVgeKFuj6pKn5bQmsI15FXlKLe1yFdSXyyW/LiMfJCLd1bvyvV4s3rDR4Usip2TY1A
nxvpva7F2KRk45uCny+9wcM4bUgygCDpM6kSoF25PXY9Tm/DCtmmdKmiblx99by/t8kOv1sjmjUP
8tvO0QrLhI8d9V05VYR60OrzZUZl+aUwRSJ6kXqEOlF8RhQPIJU6ih+jMEO54azD8G8F+wb6rXpG
Mhg7wtxJ/TEIlBepsRBGN2u4ZtI8m1gI0/LbLvqM3BN3AvixZgYPm3UkMtDJ+VOl9lAl20QXX6le
EaCbo+knNk7qKknP9HVvt6iPgglUw5IMJ3WU+NsOqJ6OUjkP6lOyp9oiZB0xJdOQLeYSAuJVK1Om
v7u8eCUTeVcFqAGSePQx+6YGR/+DLX+fw6OQKE+6aasrtjQYmiylsEDdzE1tEGpXD5uKsmLl3n36
RK85iTLJhd67HLrDAZu47o17qxGBLzwfU89v7wtHeNSg9YcoZC/s/+kRFOD3tOQkBjguFiPQvU3f
2dUDJoa8JEyLh2oDuHVa6qSIqEcYwz8fKf6Yq/1jFKlb3u0P3M+6ttyb6ogyOvk2EBiKy68uwL4r
OMtud1pk2rZGnzZrvvOFopsCWXV9Z/Yx9lQlrEK6S7+jNsQ6iCpIOwMgHIcNIPcEt4i0aMG1x1C3
eognzMKhy9bEJRGlyvMzoRakaQaHRMX8D0KAeTKMZudrqB/tif8l1oEUQUkOv0HJ2IaMgAXKompd
n59GiVdj0mPPClxJsHK8aqvpsvBsEv5v2fJV/Q8L10j1H6ZwbqAsReV+MQ9327/Zd4Rh2mQlaO+w
nLOHQz4W1paXc65YH/NZtcn6PjX9qlUbC8F0n9unWU+8W5bdRFiSLeAlj0WyCcCdK9r4X163jRnQ
6c8/32+PH439BwqTVhk6EaFqB6E59kmusyEVWJiXfyuLMLrxVm1VpeWGyL/LOoDclg+RBQr290P+
hCgZq97x60FPJ2+BB1Ro8blImTTw6Ac+vGWCE9uaxktBhR/GRsUDn0FydnMoFtl7Jp0WsRw6euAD
tJfKi374TyjOEpJT3j6YyWF0utYM8g6Yt78LhMS7QpgPMd8axbfXe++8mzAXjQS7Ss/8PTYEZZ76
rEh2mqbrXRyiLFclDosv/xG58Utghrukk5+F44aQAO3g4eygYz6wcopaD9x3JTAxeCFbPhu09Hf+
srVFB3ptDdXZubMYoE0ISp3RsB5D2q0BJ3TXyE6pQxJnT0hv9/8DbnRJMIDR345lMGbf6q6oDgXw
pTR1hjixTyEJL/PbRnEsmvyCNmVYFrgyfCvOcLIj6vXjM1bXsyibj2D5Xdzhzasv+U4Nv1+dD3g4
GxcaPV/382THJe47EF6avRz9w8Qp2jF3zwYIKrnTRAhfKu1WESgCQqrbljg5V6e+7hTmFb+Kbw5c
VlG9x0oSOInA+Q3J0RcNRpCkOnjxMPFowRLa4Dlto4jFG2CLIHliO3Qh81nnS5BImQAzjRLJEXYh
DTtEb+XyU3Q16cL3hMMkmOYbnULWDYqoCic2FZf4t4Op1V9suDTc8Olwybtg10tHFVOl4/cjJPWF
5O2GPdQVLD4fDdf25TRaFpA+xdv8W2AE2DTDsroSXfIP6FpkjCr7VmS/5KwfZKrhtHjkz/Vm+des
UVV/dTpImky5XH1Y2W/ZlStDcscvD0O81ZQqQeM8IWOaddztqNYJHpy8Bc/OgL840B3GuaCfZwDo
nsxWt5zBqFlRK3huxl8H3DVfEPWNV7rHGF9weUu8zGSpDzsuAgMBdyGKozju7Ri8HjRDjahXMH7k
3g6hIEsYfpHr8z3ccuBN+E16BhoyqNSKNwZToHVMfcRKKK2TE+66CvenI1ufcAe9ZmGoNZxl+gwk
09HuIapirZhIY6wJ2I8/KDNwHgya42s0St0hDMnlimHTxcOOckgC2tYrtlwWv0+tnNGcNor04xOl
RXyA6dMDWZelxhD2oZf7pZZHfTlJwzkYSSbTPClWERhq8XoDG9cNQRVYWgC7GKF9D+wEGQd0BJ+x
Vy4S5Ws6UIYMvKwGjATyCPwPS7vWv3xQjIQoHpH+9Lb/fjmGDvi78xr8EBW/OLE9UQtcX9EGN4kh
QGQMZNdkpIP0Rwv+aRejkbVli90O7eOvQf7nCW3bFnN1tuXQxFPAzR+eGw0k+3edLdqy524US7Ua
B9jSS4iZqQp9sQvbgkkzRF9uYQ9u2IviXJd/MyD8GN/f7cx6/DEoI39zMk/JU7W9ia6Ln5KXTMLs
/nCtG38IyD68JYpVodVRrsmYmZKFHFTAB359tHDHPEM+8QzWeLXPQDpp4S6fsBisJ0FTLxxZ6/FE
+o29I7lH8g8BNZw8dCvrwLHZzmCcFZIg0Sa84WBqT1H4pvd9yYALm7TBWQDi7G4be2GwGpUbHDT4
3E0pTAVGiYJ+8xc57KKtanJIEXR+0C4Krlx0Lmzy1YXx5D/hf70sOxdEKkd5WCJM+Fezm2sYP8bz
w6WxzhmE9uStzaFIOwsr1i5x1pUJHpSqk4XowgGmllNq9ti3ieCIYlT3Pnv6qt1mLwNfu86Fr7BL
4+Na5CWNB4i7omuobD0P0CVKEpGkPZZ9rp6gDx/E0oq1988LPmKxqBzu7x9J0Y6vF6tJ/kFObfRK
hyhzl0pqOffvBYHSLLPdi7JDDPF0fImW1OHAKOwXj1w8CACucjJhO/opZMatKx4KhZwh7VfMD8cj
tdtNun6SxXi0TMBeny/FdHm/h1s7O6uw78oW3ugDsfsD7y8Ua9ieXphS+P6cZl4yShmi2PObkHI7
qENJPGeHpB5RE3z3+QYh5/3oavSVBCU3WSek8cu4XrfqsBUS7Vp1nP2t+6hnKsdYLeNfkr1SFfWz
6CGkEsiyM+Pdg1EJWiexHD+eyY7dscLaUEQPpWg7zWHjwpltti/wPtTOYuq+H3bpoZVVA3aGejHP
GMkX+b6KGBfDO7wyIPfdrRX5tB4U4bYeuF2h0pFG0Y0lXlgqr7ndsJp16VqWMjpBGdtxIdqH4+zW
IvDmrds1qGxuB6bDtDkNOXvzggkvgvly1NnNpOy3UB5DBiD+ml72nfu6wkmDC/3YE2j6Gwc5aRhZ
sA6lds5bIbxGFG9HywRwt33htE+6luoyKYXwXCesbXAGyR8FOU1hYphFqMSgkp1Y/3CPb3s7KzYb
6Z6eS+FUNEf46lsHErddLsew1eHiRK7/8IWQ6ZjGHGsqkC6GAPuOrQRlydsP97gJIV//C3CPYyia
FJlnz3Zg0EZvjb4V7YNDAaSn2oEDpobP1M8SJBxk5amFULY0wkXqXy4Nv2JzXr4PySYzh9vpVbMa
Z1benbTH7O/+8JyPGV9/xJDapjd+LUzBYv7tWIWPqqmy8SokJrD8lbRau4OMx05JzSNdzkawEVoW
iE4E1C6WrEJ26hIn/2MYaApaOTOo/muaf8gef5M211164TPRZFgka8cw8h2sNLdspA9+4TAwkAzK
EYclH0kLKXxX6wue3vK3yCerY/OJw25B+3mij01NXLt7KEFzDVYUcdL8+QqT+UZzTYdpFpLfRpyj
pq5xL9oZpKbaYmCgZw14xtzwfLWcZsu4E+Y5i/AMF1z/G4kDdaJxui16Ym6QwxMrprCTEAVo+6fz
2d9MFjamDBNQNCJzQmOgKGSK8O3QobGRztyhEvA3/hWLnN4Xk6qj8iDCRHu1gA3HCaz6JnBDRg/e
p2Q/NtYVddXTRPGTlh//zfQYeY/7gXwHe4sH4m/te/EDU4EmxqXVJ6i/nZ+Zc/7Z203zHtftoTYA
nAPN9EeRE46CYR+pFSNbo+Py6VXASo6HpwGfanwCfwHO6Id5VnSXHwF4bBVu8ArAsKFuDnTP5gTD
QoTyO9LyYTssuf0wcYAeDVm7KBPZk02erx5+PfnOb8VUzSHTwBk5cLCCr+AjZ4edVUV8fT877LGx
9Hhe14UcDI+y8k+VGfSmfqqj0s2o8OA8cj2rBuTPdlAXVFEt8k/wRTnhSAAliVWLRZgmwcT3noJV
XZnm9brcpxOGkRKbgHaoMQTHs2JXmosjX6QJdlwUIM4uYJCtiY4W9AHY2heB4bnTkzupiE4Q6yw3
vijnzIu+MyhKLzjzVdo0oPyZ0GcTbwYVukttdwAPafTYpQC8JQXGPr8KG9TYV+B9d8JAgDTsg4db
v36XQ80n3x+dB2D8RXkiUTI7D6Hel2sj0WRwAv+huPqUKJ9Zq8/JZzly64YR5nJaBQn5254O8u1h
dBmWA7mQGPBm5W/00La7GFr1xeBcPO5MwddskAiTuDnQQ2LD0SWOdg5BFj3MulwjhnNpAGYRQ9be
9t6YMhBflrQf5QjAT1pTWRhsu+mSkgNgkjW/VDiRzAOgPb02NF6M0DP53IUr3FV1HYDtvDYJwAuj
eTxi8ACemCg/87NPyFzkYtji+W2g0bWUl3KZWRPF98gLvl2KuasUgm+8Nx2nTfotyXtc2y2ddV3X
BfAG4nKhMtMu9Ld/To1qdv60+/nsvFDLumHp/9I6f91N7Bdp7E6v9uH4rX+fncNUrrTlgAH5Cr5v
lBu3MWjHT2v/BVKtc+0DdKoNyWNwLwqpVnhaOtSU/hTrJOEpxVnslVr5epaXOTXvo6RaHDpTU28H
swmigcxDJvWmc8kL0JgFdtwzPuLUuUShc1YjWn6xEA3YZt7S+v7JBkIpwkDLuVpGPkPy8HFjNr4m
HIAosMNGaospLBg9gMyzAbh0CI3p7kpYVZ3Q0tSIUSfietCSxq08GxaBecCyOCThlFu4ppQwerkW
7Tz8YUickhjwNXUXGu4RzHWpAMXJ2zZ6g+JQO4L8eTfsnSWN1H1jER6j3IpDSZji8TBc+Pf59Yem
7iEbN2NyvLuiGfeM+TDxf16h5f/wSjW/XF3gKN8fc79K8rMsdShx14UU8BSHB1toaZHQgbQv2vuP
t8TodyMHKl/m8R3uAySSOWZrQqxEQTOsXUH92jd5sQl6Mf9m6iVVozGBRJIgZf1qQ6TFgndIPPkm
TtGjKPc8wpyhepDLjXg8xFdfkiezET6MQ7y/V9dHtWo4flMNTD8qkoXys1qDXadgy6oIQGyNBwL7
75JMuVb+oBiuznDyr5xautbOY/4v7YDSSO2llXIxnkMUDXAG5iI3SDRiOvZzjuaFLqAE6Cl+Urv2
ynGeAeyaGJbQuJ+2cfNjNy5cSa687GjzFfMWpimsYTZ1vkZkf0VWUtxwVR/Y3eh1pqop307s1T9d
ev0E9d4Ztx08PifPVOV8BrjOqdLBVWP+m+Oh7cBYGrg4MqpNaizpv8mmLQeQADYcQW7MLJcgMWae
JufzZ2bp7SdY/hSfj61FFmrip1qO4//Rpmai3WmaK5JS2FAPhovbMlxgA/eOMVmkHkVOv+Yx45zT
bUj9BjlqtpinJ9TUTXWDwWuwgilLIY5sPOZpcLX2/DE2BSE1w5m/acadreot5Gs/Il7ilzX+44Fx
PGFGSC5vSH3TbH5Npy3lNze2u+QPzH2XSh8I2ZQ5l/ZULbMgUknZW73zMAtdNbLV3AvsO+1q10IK
iFRmQYsghFDy+Qws+ayIVN9sVP/GAWcW6G1IhWudpE1IlB06LV57n88LvVeQX65M2LO4ZtpJ2Sie
MaL0ukfcdEOFZ6QRHqIGCGKaCm7qyuYQjZ4fiz0Kp7lYtQqvsV95iQH4vTUTv0IL+4J1NusV4h9T
sM9JweOuAEXvF+st7uJoNFPV821LWO566wrNcklVo03+33x1rFgkWocpp9ZJ/LEQd4hygtT2JvhP
XJhuIV/5BKxUP1f40UYFKLV+k+gEOv/+dLbcnir140cfTYd6CEVvGumOtIiDl15/7Y2tF887Vu56
bmLt/mvyu8W4+PKaEaAXNOB3tlYOuwkUzL3nwLVrRrQ8ssxroUSMiSg73m/XvfaXHPcIvl7JWdpN
qa/YB1qVI+UPP+uKkio/uF+4juJ910F0qNASTYvLGSJXmfIzGiPBYRfVw7yQ/LB/P45yPrwQ1GsO
GBdmmQKYstlH38I7reQm151G0OYacJsBBDcUss4j2ed/QckiSAuPPw9KlNPVRJaDJ9spqnwaCSnN
S3TM+RB4TAbONFxFi3Ag8Pqkv1ZcofU3QiUfLVHQOPtM1reypZKmh91ftnEs0fn2cFLij43alsGr
VSnGcgNEw/ySy67T9ADVgJiRj9pLvfq9+9XGzJpJBqUGLcEPu6ifSlWzz3TFhp8YMJjPXVZfXI3k
b8dJClDpkK6sDTe+5JCK3JliCJwrROCfPnFvvGuim4olGg8WirGxWjtsICk4S9v3RSL2atvjtnhS
Y6N6WSnLw6V8qOrYCoOoQSC9cevArF9SzDe7xp3XIpp/KpP2m9snglfCIpLpgBEWd6sEDg+Qz6Gi
XhJ8bErW4dJRomMToIJO4PP1TEUSW5CH6bPJ9xYOMrDFMniQb17IdX5UKKGmvCn6bFzc8iNUQWrK
ap6VXCdWGRJSWpk7dLEntFGwKrGjsCJDK/vL9Q+7Ulcp9iATc7/Ni54fhY2R74a+VulLog9a73E7
Dz8optPscI/NaWrGdwEFTv7SbGPn67Cm9bJFXwLUUhucRGJhqUsG4mI29O++wMO+OscqmiGU02cS
UTfutwp8ZKsNcSb6W+iNss2KdkKVTtndFyxYYJ7ZHEgwQvSA8+pD/3kJDYRSARA5ZXUxNrxz+Z5Q
e47J022BTCfpej2/BadKtEAs5cLJEOkudrBLg5s2Gkupy0u1mzBfexjLwhQfx2Gtw7pF+mJJoA6d
aCZlh/m7DPY3QGILrfTTKdrMYy45ScrNiATCNbF3dbBhE8OH7VDL/2grhw/2LC2J8jxO6iC0b9LY
kKrwwZfV6udhKCRN/q3W9B9N6ciTgOYIWo9eiG7fG7U1mA0KsI1bpcx41QwGW6Ks5nqs+YKX+Slw
fj9hV0MUebFCBnes+ZRu3pIXswtyKaDqdjkrHXd4LR1lY0+xTHX9zdlSVPLzsNicaM1Zu5+GkKhH
V1Oly0UeJdeQ8UAkAjBuo7q1zM8U2ehfBWJQlgqsRWuzglLfzrF0ud46GhOkptH6RwteW/kXHz68
8sYmnthKXQCu9vEX6sMEPVq0DVmAe+TZ2jF84JR/C1Vh3gybO2UpwHBrnZuTzq5Qs3+ueR2estFJ
1xQfTT1oe+JVRqwGdUpEIW+OZB18YcGvLfcYuR4hDnewfh4FbUIM+16oAtTrxvMaKGvpyMXSZEPK
rkR/ygdvcvjBlXGxWUMVlhSQuuWx+lRK1i493kyja5/bsFfV3etENcwTrf+UvQb/YkW8+4tDDeu/
cttijLuxwy79bbaXD8Rv+K9hu+tACuzr5VkzwnQq5iC7Ru1dWhZD54AbWQ4PF0qFiAjas9t0QeVn
7thSQNC2NAO7evR8Z++g7Y3OUdmdoODhBSizqntLaYeqCO5p/SGiikTwIBxLLQ4MCzCMQeIEr7Or
Hi6WRpV0UbBgyKGEzt6axgTCEfkKA+mth360MY19HZzTdTTpWnRmyPRw+OpPmGl7L0C2D4Dok7qb
VsV1zjRUDXGmKOuoAp7Gux8lYKENHVXqzRJz41t7ijs0NeZSfiend0LeMbJTX8guMyZ7CL+FrnEE
UQpaQGiqgWEwQky+/Q393gqApyDyOj6+xQrWdfR75HvdF9MpIkcdSxKxhta+2nx7nQ7Rme6V8ZfQ
V4cVCIrJjdztVwfgY6dhM4OjISUw62uHoV8hBtfWlsyfwsPbIQKVIylLLSDE3JI3KwL4lgwEphG2
Ku13GCbloyqKBXEdzpu2mHtQut1jkKAt4QZ8CCDkrFZOFHLScal7Mvr2OIK76cIUr0HiX7CKXtvI
jIiFvQ8YFQw4LvjproOFB9dV44vxtUi/2gI1Dz5jgzphLiUO68PuxukMEykM4ZxiaPftetHUg6aB
ERwlXSDcZsZ8hffwzWBmci0WlX55gghg9OLt6LvZtNa+5QgvkOJEvH4rdvCrm6q5ov9ExZy6i7T0
oGYDjmWgp9Ge2QwE2PR+HEzmqMAl24iw/pvPWxTq3/9dx46zyoDolnbbWA/pojHI2p0PoVfNcQsR
nKr6jVOLOwi/FuJq2zq9JZ+aHAsM9nHlkzBHNKlPQgPuI4ll3YTyLSJLMKNLhO6HWeM8DpcBOEhn
YLtigmM1cDL8JYY8sLQI6HDtZfU0lgOTMVgdOc8LE8kvrwsF/naZsHlMTnjJiGIYxQlb2Uq4KOly
jaUTR5tgYel5igpgvFiYf5ADQ2gAnLNGdUGhty/iy4KHF/li2IoXJIzFbUuHrrHz995nffsTqh5a
7SvODPXjMurSSjgRlwWAX69m2ZoluXh8BdbKErRJysYPqGrmv4f9/u4V8Z13egPX1kcFvK1FuFbW
i+potOYceM0wa3o6nqYanJfrIX53POSBUT9qOPgQ4/bIpWspF4bQpRrJKWr5cVQw153niEPROeJb
aV60/vEc/yn996XjqG+jHdLJSLdd7+RJkTlEawz1UTZoUqCmRPCtIiu6A/q4KX4GUIYYtegbFRH4
evJMYKA1uYyYKwlVnLQA2yxMVo8+/ixkHNVyeq63oEMKD0sR5UVTrirRfaVprewu7PgK5FmpSEQX
pIBOqAZa+xOG1gQ9d+mpZ07oVN3KONyz+KkBS+3chYzm3cv6esbCK+a31qupxnDMGmagrgeBYjkM
sjCQlLW+67Lrf/JkVMvBAAj/iZTMNCmUnXykwt4XLVD2mopYs16g1ksqO3komfgBojrsRiOhUqPn
dbS+oEaM81Gk9KovvRlKo0B7Nb+rdYMCZEOR3TVGgzQqWOul77X3bks7W4qsl2HnGPQrTio/sWOK
5jG4gH9NixicsGhw8FnlyN4dripcryQRn9p4ffcdORzDNxyDz0oumrrN0eloy2T8PT9xxVJpsn8q
14gLW5baxr7jiuX54wcw7rQym+blZjFZqXKyTznEmejfC+dmOjd3I/ecyll2L5sMx/noS/zuQIqu
Km9R/8xbh2giq/dmQowvdGBdzBGrh7/Tpvdx3h5Twb5t/DgbP5MPHidXi8oEWU6brLIc9Zo/Q8q4
T7Zu9qeab9KT9CixuXbigedIc1UC3VujqzdWZaSKVZxK4DlS76P6+ZBqTbgDxbiiQJ1XSybtE27V
unKjRv1HvF1oj+alboeb5wQbRKM0LcTU4jy25f4Noy8NBEEADfBXFAC1XBYMkwMvNgW1RpH4TVz7
06uwtIRbLTeOGZfSyp24XqHNhRe3c3nGw3HRNY6wurXZtLGKiULTdx6bg1Zma7GqsKQz9MwkBUJU
jrSWpswt9fUx48xi4Eac3zILfBx7rZCNtfJyNg7/ISabs5xzPYz7FOdSzJDFCRxEHCQ/Xp5XSi8B
lbkk4FliudVpwEsYatu3BD58XK2eDlEGKZA/HkqJzbdnk6xq5VLrgozhW2fryMcCfLuea2YmFPJX
9PJS/iYyq6VM6IPGWUgG63WuxQ1n4vrNs9dn6QKytZJTECWYN8/uQw18lECMNIAzdxPzmY8vlUqz
R0pVLtHEzD3v/h6ntB/8FtfgnYh9p3tiw9alg0vaPiyR+hTDrb1+CjJeQ2ngRXVEv99DVwUQek8F
KtulVXi7Y8o/ntPkzQqsjtPhu8BLxoCugZOqsjZFbmAqC0IUbMe/wG04qC5u7lxbHjAxMjpwKoAs
X6KJlPx8JF66+gn72Q3P+39iyruE25El4UWOe4yE9wftFi4TlCAAKoafIvqNWuPYOMbn/s5BNLVq
x2cTGbowl7Hm1pyyijWnDgwaqUi/TeNCsiXL8K1/ttRYUkzuIxil/Fe+s7E4hsjwM/Pc2PvZEHZ8
aep4flWGDGw8BSh5FbQAzTE9pmMXbyJoOkOTN0v6CzIOIHU10dpWOAC5hwHnH/dJ2sqbITtgYkce
5dcZVRBp7VgnADUIbieCBGB2uRk36vagFVszbThfI7tCYeB80igZqFDV9wp7/3fKMYaoYiS6xvR4
w+dDEkZnKMiuGcABb1Pr4XFrVdUefHa3OaiWflJqxZ5dfrUTfgDMETiwWhVyUOGc0d426gfVHt8k
zlm1svl/5zlz8O0iOCQ2Zuha3DwlyJ76/+VFs2dASDPKDPD08Vp62bFiiCOGqw5IWWHLVfV1qejM
vQelkcw2CA66ETu9Y7/IwO3HM2nrIBDjxvPIYGqev7P8MBj4qTwQ4pH4euj+iZRUaZr3PmUjqA84
2nFnU0C4icBqfaR97GdJPEFiFklIoR8Ym1S4oss43Y2iIt4+2JCXh4evmXRp0fGJhR7HCCTmDLHn
rdxjuYydpmN2QI0nB0nRARBz5A==
`protect end_protected
