-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fy0Zorh9UucW4CuVh+ntptncupPAdkcGwPItOv+XY9dAUlrUAZPhRiV/S959biu2LzQa+h8gukOQ
HOkf4KlqtWhSpgnJkreXT3lBEyAp98vDOgdTRVZL1KrmEqh+IZQWsoELTJL7i2I4DErJFb91HWn0
Ja9GCwmk5cP5rvoFD5n7hwka4LBehudUHHCowPr13LaGpKHrjjcs4OpO//L/Z4GitdsVI4ea65QW
ECHSkJVLhCTzCcvWaHiFLsngJ3HbUFzKLQnfqpCXOnJoamBbJGjCZ7CK1tX7Tf/GShPtvnlsNJB8
B7SrDHwn7p5tVVBnEzU7O+LWKDD3IcBWZ/p7Ow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7440)
`protect data_block
xIZSCVwNGcutfRmEUO/ijyLzLza9nfWflJET7OkuwyDc7DMFIwynppvlcCAWuiF8lT1LYlkAspWr
lr9ECl9DIwvgTs3X3De3WfcTRHLb2GjWo5xqycW5JNzG8vCbgyieb4ILNYT3CZqsp78Yl1mVSv2R
VYZNEWIGD5PlZvZtHNK4ocBRAVEjssWEEPL0Pc8aPkL/veGZC3efya+SdNZWXmfbd05lwynGZf85
cdfnz+4HLiMAZdqR+vZk63O/J8f9hh+1d6UqczX9fjO3/upBqxeHzEZMLfvryq+PSHNWHrD3Q5hM
zEEW7SLIIYSIUA9zjkhgDvcYzktcl/ZxWbx85G9ntWGTS+fL0ss3beQvl6zjJUmA48SI3I72crXH
rEtM8yGse+KP/VHqunWyn0+Xn8i2/YH1TP8XWBXdheIoBSFTxNxhMysxFeAAdQbrpqQdLls0wXMD
ydY4ndfTSouqrob0ANSvOcJ0zlkLuxuE9ViXV6Frf0GlygRCGiLrblecCJ3NMK1IvLdPaoC8uwgk
RABjDyxFw91098mku33pNAtAq+3d/mXJBkcUZyo7bvxy051XPGuAfyFf8R8M79BRBaprjbMi+fVX
K6sM+8F3knu448tZy/IjeHqcY8KJAofHIkEgFeQIKLFtNKIG+y9eoNGOQD0EqbUWy1sGyZxtqGnj
Ve+J20CwiHZA+9wXtS9pJcjGXI/ULULPAFvJWXEQCP1Ce6NFiRuTtPhgklWcWT4AbcvypdUd3P1C
lU0V+RHiaqobSj0USWzdAwyOHJM9mO7/lZxH1S5NGDEjmC4mVYh7qPVN5l68lizsbxH6Php8vwN6
X9tnAdwuEEPYvfj13RIHKmOOUtgkmTyOEXQvvKOyc1cKv4KFAMMlxrqqx2hJhmO90ip4q0J2tlUE
vJTl8fBr5vPjZiHH3MoBQQ1eGpLtHBDKSPQ4E1KAOHoT9w8LG0JGmRyakXBTiGSBa08RiT5gP5Qo
7hcSiN6OJWhnieKhg49X8q4Yfv6gB2vkTU0mcyOmwWNEAyoG28z7Fse6KWTjU9mR4LZy0CqYnJEp
l42hCkuKNgXkBmbt5DlU4xuBttw+8gMc6td+vK084wU58OvyzSrUwQqEuNfwMxwAK/R6yfaks1IT
y/xJ6epEADwWS+Jz3T1gJm+IEtZdL8rqePzGuFOzR01XpsFAVB+502w4YeiM6AEF9F7Gv7Y1xUpf
S5mGODtjF0O2We6hY1VJtaoHgHLmWjeZf0Eb2P1Ku7x+zmxygqRSN7iiZU2BC6q7GeEZaoaimXZV
aJTGkfhffqxhXfkZgYQvXhaOytdMCR1U6FZjSxU7X6RQQQRMEdO4ONQAfF0FoUSECwvwMDSVauyj
+DfGYfnwcv5woiTwBvjx7ZIPn949kAOz6XF0E8Ez4AGauOkhtunEf0SnvQaYxfpXsKddQn/vTAed
b6kyvK0eCED5mSevf/dP39UOT4VfG9BWF6Gb1btI99qWfvTj4XDzkoUwB57wwjoYqperLEaeusEW
I+IkJC0sL6mYvMSAAA/9me9X/OYFT+F9idECxmfc0rSsuxbirg3VdDxGAJ8Ffbzv+hb3xvRdzdIL
KGW51nBvzWaxs1OmjZjCBK29n8aE8gF1KB+Ho0MAsJWT5P1unn5+wJwXSTUUvm0jOEryhW+AmmlS
VMqR6BY8u/xf/J1qUSd2n9iKkpc7hI10kmCrsuAIAYG3JI+3uKDIgyGBZsUUTXqvrs2n9PG9NLKO
TkqKM7liy50n0RfkH0tJOATuU93tWLxDNoPXIhLOhKvsEeD/YMGAvFBfQ2hg4ASYsWSaxAagEeg1
dLpO8IlCY74jwlHEXByy5Np4RDeshGArm9qHmgTxpZC2kE5q/A5Kqr/XNm+cjWfZ6evYd805q0Ss
J9l6PGduxxn0qv/Zn9HZTRLUZtvEZE1mykkAg73e44/1803sK55gwgq3Kq8AbMxtI3IrnDwxwAbu
Ye9iqr8hHhxGE4T0Bl2S/VuvXsphCDfycUWPPqCD4Y3gSEtth5evkCYGctea5FO5EbHeeVLrzk6K
OeERDcnsYhc+H8380xEWWE/2kB6BWKD1ayBlp4NDxHiS8UNSejDJu5wTJuys3O8WY5kOMl4AFkxD
/jmxbUi2O+PXRdejrv2hW7+XvkAX9mzY9Gvop8lvJhNKkTiQcmlGPvscNeA1sgp8dKqz9nNbm/XX
LPpOASLaLroGLGY/VI+C5C0AiUN7tTPwaz7vBxmlEGEBwYCNbp7cuNXxlCkD549yhDPXmYmMcKUT
IA18H60iXEuwVXfXfgqnBvn4rPYxylNucr51v08hHJhAdljYXmm82SVxU77DfweiciLDleR9h0le
j9lvOjTsvGOLK1iu6g+w+NdMB8imtId4cy+frep3muQUuAhMMBx+STXZfOo0fmOgWEwcBlBWrze1
ha/GzermW7Dn3ZwevvnG9a4xUgzDpMT3YET8NiHgmPTUV8sMlGR/avXiNYVUqtlVW3sCs7O2jp58
hUMNM3BWc2spbIsRa51hlew/eHHDh3oQ1jF6ZS9LjWZ1J308WupLTeTNTFmEGUoeJ3MPus0o7zvN
vktEN6pGlDEZl41O2RhureHfMtDSbsEvFDTflfx/u4YImYKP0/2k1TBrs3ShNEZTknK5Q7TjYZSh
Umvmrg/bu8cKPjKdbt0yh0QNIcmm87XPWxtDBBK6xLr2zGq2rkkWaRI2vGfgo9M5jHXGm9DVQNHz
WtTq1Y0vfvATPsOdzz8G+K1Ueum4HKA0wokimv8cwHLM/gjanlVe8lsqC/r910FJzusj5+R8CkK0
+ZsycAJl7Pd8hNtKuIkZ/MtArn3J7L5KrghrPSXsewDbWbrfNdvmaPcHUzEAiiY2xtdfEt2Atzn7
rzg2bZWJi9GJOZWVNMi+up13A8unAur+10HbHaCaOU9bZYF2SkgOCkpUgAsnZ6qcaXcEzW8Gegep
H4Ad9TXKc4fHp+Qpp0RkBdobIi7ybTsbxTpkxNPngzrLiOo/vJrBH/dWRcz3m7BCbo8FAuMFwg4v
E3ivNnL50S4B4+cJa2mBzQ+5Vuqg4PWgMjhzRZID6aaPALOEODjLaBzJcL8nWKI27pYqUOjO4jSa
LttexLj6LWmWkI4Y8NGYVi76XeoFMy31/S84pS2+9BxgcRj7n3BVhoM/8RqWL5d304GZ1ppQeaP8
XNm26F6igRROjP/iKufx8GQ87G3HPdxr4E7J+WPG0eMolCBl0cU1CufqeImojaUPbyiULZfSEplK
BEjeaf4KHJx2iHCUQkGdWWVQ1x7TmXFhR5YOg27LM9NHozd5sNC1VEOBTxxoKNp2jokRPH1grpom
gP5ivFd1/02RBwBziJq/MuY266ZPG6es8/tXQ6l+tTNYM8mwNCZ14+ww1V5xLABTQs3a444JGza2
KveBP7gmblf5RDDKBp4jc4/phaHZ4ZiGCNLajZpCNrizaW2+zT5WAai/fUFeSuYEq5A6c3yvG1TZ
flgxZQnKwbGa4XJ0xjGA5btILy/ZuHN7hmNnaDWjMyhpJwlCtDvDw3jy0qHgjmbkoQaPVqmd9ok0
fTFjlcJRg2cRWFx31ohTTKIsNUrFZcMAwnMQzrt2YGr4fnJW0LLbI+ZVWL1WLLsvohhacB6il8kX
6aGx6/SODKOuxOxBk0dcJMHIizK0feeRriz1T7ykq+EFqjRinunJA/ZpZVfwcKJNBMgMfGNgTbW0
Am7zNXJTF58yw2EU2uaFqhrzuloCujhsAUd7DCLxJ9tS8VA3V2F8zILbWkYfUlL53YSWpVHvIS6+
SQzmLOCLqob08L0zAtmn/kqOdHz3gkXVdWwqNHh99DKREnmsAhNHJ18ZQqyxtYoMqDv86IfBVK2b
vAAVqmWjV4s0W5qMlH7abEpH8R0sgIGOmHC5ML7fb4AUJ2Opi2FWwhOsRDBQvY+l3PrSVgStPEv7
BQFMQUAKPLThaYK3G9tLLFcusOxSlw+LPydSVRUEsf41q87tTrbe+M9xkY8ndYpW4R9TcWrSgkbc
oVgDqSC3fbhcoUIC0U/ZXCsuz5lGxpoBbOnSCAqdcOsT21/ZXH+vmKiUfueShCajlirRMsMkBVu+
OGOLzLJapm9BoqNY0Eayi0fJQ0oz+PRO4CKFxuOI18Xc1owrQCECaGjM/p1SvP0T1+DMmqK8UrSg
VfumI4IZ6LCp4RxbLrN9iPhVvPB29gy9TNLPww1Du4HVrTzvoleiCYxyWDlvu1bWFHEvz4F6iGj4
nVPVlpBaWVa7OaDFEiHOAI8nifOxOaC4vzKN0JuYUYLF4BKNR4M5BSrBJLqEL+EF4d0y+K2qXDTj
O+06grU1ptgT8d5skP6lvgR2StGgNothni1nqFrI51I36BFy6CA0YpoZw7fovmqPyBsn2wyAkB+Q
MlcZr2AcWkXdZE6JGCIJTBY/CumOzs7ZvGln/O2VXlcULP4h5QPztPn7M6J+Qbv4JIOBv4dSzJNd
kDOn1yxSXeZ1FJg1/Y0xuTnvPdOyYxq63BApOwVr5b5/V6tZeOf5II+eNdT+PAC7iNKylVHlvsBj
/4Vzysw6Hmh4E6mqXej9nq2uAzMEYyJIIjL7wCYYf17oijXLhytwaBttooNQoAUcKXV6Le2jOgcw
vOQX340E5YriwiIvZvm1SBlL6C7/820xMnC8Ph/ssP2XgoEXx5uuucwBwO6xEg+mWr/CI0PY/xZO
qxI6wESe+OFjACagsjSRIMUfkDFPTkKlx3avI+OKo5dyt3z9c51czuMlOC8kX7NuRB5aDesSOJE5
7xyp49vDJscYeSkBrGzY9Q1dh5ffUwNXVOTmM8IPlVgQIt5pczdwM6ZPOS2EJbCGGJM49572aYet
eTLzCko99A0BNTKSyeYxD9yyOc24n/9VfHmm4EOmEdRAQQvLKqk2wyJZ7k7rE/vfqpEqTltaGFom
sV/wayEMoBwuUWGoS/AQoh2LlsfFSrzGJowXTHfkCWfU99Z4m6nQnrXL2RtAYktDKXLnQ6a3diF8
/htImQnUl+71nlWuo+Q71geomJLF8GzvDyQckpXUekzcoqk8Su61Rqa2rFzOoHRvcDTr7/jHAYQ7
VOdSlKiPTdlSDKCTp23CzZbW/Sg+tCpjP+ADPVoas353qvS3UNsj0phmnkwKtlZJZZA0ZMJ899Vg
pMNPSiraJhfA0IiqBnahZEHcNGgU+RHvdVsgWh2HgmoBW5jogMmPyxA+kVot5jsh/2dXnzXct9Sm
O/1Qr8g2rM6A6EWvOvM+h8c4YlFtuI6qOpeHmErzbffmAaHupdnelNPUE0oIGI/rMhNDilAC+RTM
6wOuoYYFmCE8D8E4gpmbPQuASCsyPJrkhTxeOkcz2V74cvG/oiTms7Q/2H3YOhLVSNpg3hpdAg6V
8QGia9i85jziDdpF2bZWP2Oqt9VvUdQRV9G1iDi+BkHJESUm7m5PO6wWI0kt8zQlyPBpVp8bV6XM
oKUzeJtE7p4jM0XRWifgOGHBOFvJcxg72DTy34lrOqPlC/MjzYsY83bp0MOXARKcc7x3dwZI4jF/
2uZTbNdvKMuAr6R9GqOCxBbK1wcpa98P05KBiVHndxX9+lN1sO1QVQTR8EXala1yJqUG4iiMrxIz
eAw7SHMI/+o/p5NXKcSgYeh87udoS8Qfybr+T86sIBxC7uM71Koe+/7JhyBFGP5IvDO5BrliutZq
T5fPZ561XUd04U3W5SHaASN2hlC3Y2Wgf73bGJ5q03i+66PKmuZB5E7ftdr2MWexEA53Qz0o+x/f
fh52no41U3O/VnD+4thABS5Lw8rI4vqpc3Pbvo/CtehhITf+twZ3KFgJBrERpOwmSZkbKW/w/rnl
mLrfgYob2hiI1JkqEJFqWloK8XmB2v01rMG3Ml8OuOcvqt8qtfcqeakMHSeTSNa+ZnDTJxsBIHQC
Vy55UkStAxwXa4w79XdIlAdV+rFpSzTJ1YdRSpObAVnepM+gwXk63uphyDTHlboqw5suvGlUbhBV
tW2HCvRgla00nSUZaHqIFq1ugOUwD9Lg//JknfY0HceoIyFVSZVwvZbxSxXxctrV/8mRbWo+6FCw
qPv5x8rcKeUhACR+r3YAFbvW26LltL64yZjZW2YBJ9k9YqoOxd87r+NmZJHSzbtwv32kPXVqyqS9
J9lH4eW1kvrjYpxtpBpyWK1FuRXoxjabwn4sLoKOqhxtjvlTX1vBcN6NGHGhIPuBb90KdaeTDjZI
f6t4PFnwV8rfH+ZTfEttjm29KsfxuDmaZIm1LmXPEYGpm/PZ3C3ASyNuihKxZB0qMrbhbi1EYqL5
J4h+MXWhZl8W/+yYvC+gS9/v1LdD5sXlHBZzdtMgQTluS/688+MVg2zXoizc22iUtVPgCnuncE2I
KcbkZLbxcTvtELemH6tI4olJuOJmnfPz2rQBfbuAPcT51hrhHQ8yrfacEYFA9dtqb1AokP6ZtrZ2
wFN3jPt6LkZWeJ2eMN+2D7whz9P+U0rojP/Y0u4Drlc54vLroB+3zQMXpxDdn+QUKdUPfKnr9zjO
NEhC5lb22KCatE2LmNlXRXa/M9B3rnmsegInWQiA2uh6mcR9ia+TUCw4WaS9qt1mCnJphWbgQmfF
u2La/7Vnphs2m1DvjER6wFimMgj2+im63GExEbjUMipHJToaEv9vYrYJLqEUSO7PI/kY4t2oG7cl
lcxSmNSslmJejec3lTT6774d1Os7AkeUC0WvPrZOegCqotNNoquLCbvFnQk/02bImN1VILeUkQBc
a/YS1eD177/Ag7x4U9KSvlmLtSU4OhirTbL4+DHvRhB+mAjHVc5Pbmglm6h8Mi/FU/nAczKi7bC0
dU2q58vQi+jj4fI00WY8XMjTGGa2oMfaLb2e85aW0RW2CvzIK4XWD27bIotQaSezzeOwxTAEjAh3
pbo4ZdVIiXgGbKy4wN4DVz3fYCEJgGkSOIy7PjheuAmuLWrCoamZIGC1+ZknuzOOnjsGxuFReh1Y
GuT5DoFEUhe9zjm09DZQxwrkWsGH5GIJxdnxx5Zll4eABEMudiwNGOuS53v+sWDWeCHtIpO4r3N0
T5iQO7/R75DYq9vkSlJIiAXIRS+DvbTA1dcB3XYTVHFh21aUaZqQMyAeMBAevH+st++3UOUJVk9K
YdVV+tFdD0dBj11yBwSjva149UhjCPVlNL+wdxieDkbxFSSPr1XgDq6X1qsmMMdJSjp1tUq1cLJR
wypwXYFAOiDhQQUGNq8AUG15ajrVDsZfTLFOOEuRwovHunclOrr5G/9l/wBi0++a/vAUdaqMbQkH
rZO6mV1cQs4/ikYwJ4KTpa49C6sLZFk4W3r2GprmGm+oF+1BzxpXDtuykdeFTbP3KeTw41CuZ5XE
4DXEQVDRoH39X2SG4WWz4T9esGm9FbpXDI+EeYpsaLZTaMkvxxX9YM3cu6UammZjsFbUon+smIjY
hHEfFekbbCXnL5D6bwX7CAn6ol8wLoPCk3u7t4ijLtNGWSdhhxZHcIriIQxGxNwb/Z8cF21A0c8z
8usLUlxQhLhVabETwWQq/F+o89HC8M/Fj/oXrFgGu6cNPPIikF3ZExUN+/3AQQC6++sin9eSUFkt
fDuZfE/aRxCWjfh4zDzMhMoCfXeEWLdQ/1+/Jlp7/6fxCRfeaC1YXOCDEXaqSiu7v9gU7NLCZXVS
sdYxyaGuhX/n0Mh4vnw0ph1XMgWyboBR25C5+r/3Rsu6HNKeDqhldL98wIfzD0gy0g2wvb+2Ij+s
oqlFpowfpSpy5p4VajwYgAzNo1FNiJYgSzv4kk35CgDZHIi1kTgK7zyHmWiSuCAtyEHxqVCULvsR
h5OcS6fw7oFFt4DVpTAPN891xAUw5//y8zuA9ARhg+9x9BIym0C2vMo7rG4ZaOGbWUbG2Rrc9jcm
7s/7W+YqBpE8UaGE92O9I4WiRFAo4fYacmoxasOk0qB2r7a+W2Hc9lAucYSWb8d7Px6DKl0nUJ8m
ICROaEMWWNU3p/FTOF+t/rjV8FuMah/zL+9AQEYVngqX0YU8E9xIEGXXtcYc1nAL46DpwMFg9IJ5
6a7oSVV3iKcGfHA0nNHaXjIFiNMcxjkdRCe/7KzK1P4iGhJ1jKuitfuUhYHKiT7jQGHdcVsYYyiI
1baHxvWSBUc0oqiedSTtD8QaqCN1eBwg3uF8HnethO31EnWr+tlfg6g7seSQ6BG4tvaCc0wSNGxm
TRHMrvSQ3ffrwdxp0pLyX0zG0Xc9hnFNqxx1qS5JwVmKW6YNu1l6dmQboVkdVwLGga9R2TF2jKy5
n0GXk+p1eyQSCTB3+gvEUI/OX8PsCjv/z/e4uqbdTRpQMUSxP6CC5mXmC8kywf5qf0RLZkBoBD06
kbGT13N1Quc+ifQf9tg+2Gd35CqC2+5xdICkqWVXonubK2cFJpaLk4oriKRLlApC6bRvKBTC3cuY
5GmFBGnMGqNQ1hZEDWL3B3pd+SnZnrALK8zwsSIzT3IKdjVdlwA0h4Cm+vZ3TeQizk7/x29Snt5f
gvI4QxneSoNmGP2nU4Aaw5Faj5fbZBUsVvS2pf6DEub7MJOBYuAE+ho+/41IPbJqDJENpESnEtP9
vyFYaJgu7spbSUy5oj8lcKR0+6vDis5ikh4Y3UifyW+xjqBcnKs2+gWfWx25GYsJrFFZf2TPRnrL
P5K9y9929ncYYokjYdrw9VddAVvoCLA2NQYyC0YANon8K7nAn1ndijjZpEy2zupJwhz2DUWdLzWk
vIUimQvMgbpvCxhMyRIVOzqJWl0LxG9DuMVlqlHHJM36MvY6zKHkOHruSPVVV0Ys5Imn8tB2uCGR
jpbE/cbEbLdX6ZIZQfkihtn4UI0m1WWAFRXdqhio5isNP0HMeDk2OM3rcfjg68R8hOGvqkUub/kP
wAM41DIjKYVhU9BeZJ5m8YVFHU3HqqlcEX2E4cLKjiinWy/Ddh9R8PfmWSGkTcLmjPDCKenO2Iip
giJ9+neVYZdVrBXd4rjIneVuVtZzDGXnLp3xH9wD5w9Xu3A5ZzNmVTGA7/YG8rwXkhWgYC9D/7Mx
mDPSVkOMWmFQjmXHz3yhbOL8J/ymutij5IBPOSOrRuFLhBXfchN+b7Sd6ZJn7YY74dyvldj8ZGZn
7BwevDNp8ZtFn8E7TdpUV7xPh9vVvuTpgFxIuGXl89syeOYwnxPZtYt0pW0X3dMHzDgOt4+a2bAI
Q7haP+NQ5k1F3UH81np1TlYiWuhU2JyriJhzG8mHq9UeYMJfeXBZN4BI91H0QvpsRysXvQN96UEX
D83zdnxKEz9okJ6A+FU1T6N7+aFRyiIA/3/U/qdxuWq2bNlZRR+4nCYaGZD/V0stvvXwla66YRun
Yz3SJWksjZpoooFN7pN8t2F++i+lUWrIhof01Y74eESSr+q1+U33T1Yo1FcCwRh7kkoVjREMybRg
Ayu9EBWQk8wCFGnTQykYgJQrs56v1yaqnMfR4IDrPSde7rQ7MHUisKjISnWhECriBt8EI6o/+1gc
ID4qAwdi5cvyjpAWrmcuCJ8HtQyVYYItuJo0eMDMTZVUFyeiI3BrZNNICfG157QBtkKqmsCKjHZ/
U5tO1mbWF8nsvspJOV/ku4EYwZaWmvmh3+EMoMMduVp29dOx5m235hnHLHcMAxLKKFIHgdMSp4dI
nhgad6rDW2i4I9ilIWhBiWcClv1d7KdmxVRmf2HSB3jCgzZ44/ZEOgX19HOY6iOQ2K4pyReqSmcU
oeHiXc5kH/drBf6vXkNIQDtVlKOruhdf7UXPbsidJeA4TA85IMMcHT8g3HExEoWQAgXSEPzlaZsM
mq6c/X6gGHECh8f9Mij6uEYv16/GnBpI1h1Y6TjyUVTveBrrbt4zR61tMejT2/Ovj7BieaxUgKuT
Ry1KGtsetf8gqOY42ZeSGI5AnrFVgeWzE2kOHDcY
`protect end_protected
