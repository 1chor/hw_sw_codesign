-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
7F9fowa7moyYemocuP6IilyDpg1EWpJJinanlfgTH2nVTIOBxrUJTTmcNpgb2WDg
amPHXN2b61wOodRcynI8cPA1Y4lnacL/B9o804komcXYDH8fPJg8u8E1QmHsdNH5
KArGPWHZExGyU38vRrY7vpMkMYh3J7Ew/q8I4EHmeEUVZzptNIdnqQ==
--pragma protect end_key_block
--pragma protect digest_block
9MebkJzoQqi6JtyCrpBSYc2Link=
--pragma protect end_digest_block
--pragma protect data_block
aIJdvTXJaxx0XP5YBmvGsU9D1J7xxHwsmdfQmzsc5NbQ5yKQ4uoKAdPdv1oasP6F
/NO/3d95BO7sW35Qk9qEYnDYTJsUqsd42DgUoGwQCwOXQC0ShFiwKL8E9zMPRgxt
xMxMOLSk6UEc0e/EYFe1kb8z+rDsLg7mYFPoMCDJ8yZXU9Dzyftnxlw7WLCEBsC/
fu5+Qx0uD1ns22PHtqsWNExwhECk2JE5OO+Jp+UD4yZjnpATXI12tFm96QAtrTIu
5nyG/C9Njlfku6vnZOj7pwqkvQs/eCcOCF1fQbqmpqmd7cLq2Pgt00n2vRdmln0w
TmT3FT3qYW0t0o/uKYBjh39yze9sIwBoQcvjj6XLlVaJi/lb/v6BQoc/e8hxegTC
9hDZKgNpR2psQSlJLeqPyQ6RJCYS3a3UpYxz2qbTNchCoLqHYSLthSDkbaPa4rIH
Fp2XHqrPoP32rAv2AozbAbcxy66WDdbFSSDPlhkt4FaGyjam2v+tvLVkAzWNxOb0
0/3BSNA93ciHDgSpcx1piMS0Ac7VBH0bnT3G9fcZmykjVwN1hVxpc8BCXk15L0Bv
knGxWjCNERypVjxOHOhgr0/OTqEXhKwDrjZl6s4TjHxK1YJONm3pFIcX/HuTWOIz
4eDenjv7swp20R0V4YwKrUbkRRr62kTJd+BnRqM0cdXgvjLQMqEN9IkpcL0vDoPL
xYSQNr+dbupeWYV+j5ud7e3e8q5ETFMVKMar2jkF5qJCZ1PX0jggJ39WDO/+dTEF
Zn+liQTC9WLwGLF2RZ+ol81hZifcuhXo1cgM5KPh900Wai+pAjErZzBlRXZ9iNy9
v6P2X9i+6M5qAd7PxEJB9jcRANdykROcAgGuRmd8guk9v4Ifd/5Td4DA8XG6x5Wi
CldF7q6SW5r5wlN/c3nH3otEiLvCZYTLl4XG+YKJPyO6wX1GtWXwcTOuJNSd8cAQ
8023ZeVeiLcUMW/S7MaDnunhT/pv98iFaEwFYbdmgczfTqTxHJX0daobzomZKtFJ
CZkWoaHCsrPtqJfw8dAPIc4IjAyJNmWTqD3ldJXP4WLLW8GBBEIgkPLF2FalY3uK
A5/dK5HWhGlbkoL6wgY0Q7O7KVaElQIuUAUFRtPpM4k8zSw5d8Q7/RfS0wM1wGaw
MKIoJ7cLENMN4weJB3Cb+GUiKc8E5n6EbYdk4ouAgeb1pGtCyA3RjbBqLoWaYgY9
mueTFHERm/MAU9nTI8FAFN9MGGJRL3SkTkzx4XtfNC9Ah8Lxx7HjgX/K3223r6HZ
nMtgejrY6PUUoEN7qRGcd1cORxNqMyiEioEaQKeAwNPPr6qtQ7eLwb5vl6PNrA60
K4l/DCNLqrJJAyeN+uQ+OHPFvfQuB13QcHWM9x8Y0yPLZcn/H500o8xNvkPlN+Dw
qGkvtvTyb/O05FqzwoFSJw0q/Izho30ecQD4ikoBk+8Bqh/zN3n+6OJ8Put60gIB
lwop+4xwugsVxQxiKttyyRbDDUNA/XYzrNsrV8PpqsXCzdxhZnNRG0L7Jv5moXkc
ZywUc3C5qvA0Vyw9V35RFQcp+Z2uCiLUpRYUTHvahCEUXbmpTezBwhyjpu37qUzC
ju/hYKlERN9xnQa+rtj/Qq30EblMFynZBjobl0oBnEktSrbXNq7i5MVLomQlutel
8oFkBt8OGKGYaQE1qtIgBIJa3FNw5i8W18tKAiipGvey1uzZTNE29NnZc7TaZR92
7evL3oU/6o7EkZ+AzoEwUsXToM/VSheXUJL0kht9ZWNa3vIsitBZTfJk/WyKyWSK
W0th8zvFz83dFK0oHjp3hU5wqF10E7yjfQnf3V6spzuKWGBiLQIfUxfXj8NtH5Ph
+3vKBMGFS5roncBcKT4hAb9rxVch0Ub7hlSGqUvyuHF+gca/Xd2fytrDt+XGhpuB
hFTKFQmWEVG8wbKli0hyGAWRiEgmej2d0h3hygf5hF3Q26CmIIICqU3BgE3zE/wZ
hoQjd/0nYe1V4j7mp5+ltGcxM2km8T9jpceQ9u/V632NDjTrhuModmZ7Jjweom0s
VG1P3C5Ck81Yq64jxpFT4HssljlJyg8rcqW3IG2+JOS0VL6lWb8nyB6QVRiK4GNp
xQJJV8sFk/Z7us2f4KCs/np5is3tgiZpaycM+cIjW97gJhobEt2/abCnCY2SoAPd
pX4OzjDxhoTdL/x7UgGiBJ5/MAlUUDow4Ha2MGVNe2M+SKpPgGpGO8/lFtbu8lHO
aWovULXZnnCNMU0X5PITFVGu7DAtgYfzk0PUQUXWxd2mR8AZVhY/SXlUmZPyPu/3
VhXcSbPDjEIpFRZPKmMTxy8jkZIUOvCR7mMkxbEv+J4m6MQli5HUPWalYnL29vsk
FKlPnZjnbFLcAVDI7Gt8HlSGwMAi0/nnhcB/OQ/c+Vm7isTMT8r8hzy1ELfOFolw
hySUI1P4+utOc+6ZOhc0PKlEEODoh2VpMC26p4KBwfpfvIjXLDgbUWTYsebZAnpw
g9lfar+jL9LzhLOXUoxRaSlVNKOddqU6FJBpFAStNLE/SE+q7t1wmaD7EfPv1Egb
Q7mBp0rz2AWVZC5A8lXNE4PkPYBQ6aHIwyqgRfTgdh5Up9asHbe/4NWDz0Wq0pb6
nhLGJKwjwdZH9+T4UXXRLK3ft75mZtI+T5YYJi9SAU0ImBCTDg3jLr8LI5F7uLhe
UtQQlyIix2r1xAfh+h7INOa0NOHXHstB+6UF5o2CQI/uCdQH/jOYKlmToMn3Z92w
DcKB43S2UpJcl2++NOn8ThyQ076O9rDn6vZheSmmigvw9/9tPkUerzFThss2P2CX
BxVxWcTGnYmFODSdV1XvyWpID7gVbq2pqR+T0ps/32a3nc3KAJuTtN3fIhB9nAcf
a0UPK2fCV5mWowt7tKHg9n0nhLNSijBiHJXB96Az/9avhRvTcWRp+hpeKeyIvmZl
JN+5tkT5pQX1uHR5ogbsBPAUR2zHFJnDECA/l1J36afsMG6A7cyZhxwxWcimGY0t
HXkZMaWWYOD4HHzELAuZiR6Q+bWOy3rls7O+l+wqijtt0ZMhYcfdDqpjk25RH+sA
RbndRjv3YPWTwvX6LCeZip8P2CU3pzVKnihYrRmwwEDBXmOaUQ6Wdx8Z3KAQ29LA
eVjd/TGH9xmmaqw9qHlrSHL7o4wcYlTMDWKfh2nnb37dOxfZJz2uqYb7EiCiyLMn
+hrBdPV7QapnyBFoNjwA5jrhPmaNmz4t31gm9mZpDFyG8hAyr23qSYVGeal53Dpz
87EftULKiL4S4oZ1sDdZe0H7FMoXa1xgptNJcJdLJQklLRe8BCU9k6u8acktT7A6
rl/6YmwC/fSUClGjpAF2o9WYKEBT7dsyKEn/BvJAYU953cqt2xGSbpllsP7re9CO
cK3krlnDgQxosBfUcZwlvN3FuiPEBX1d8JbJqmhde+Y0xSgmCMCRyXYQPKpkhHcz
SPcRNAzusFRKDdZQlQr6BDoIaLsGI8GquO0MLXJW9ddfU2kX0Z9A/s11UFbRmxC/
OfGCuneSkeqDCNjgCESl9o35+THpeApjKHYfkSj2wQuvt5yG/ZRVyfHxibuk91ek
hNaVJJ4EwX/3fsv/q9TiKmU9PMcAnF6XUbnT+zNcALqPqhquBF/UJakVNQh5qHmj
ffKpXfpU0YlkdrOVahAOB/AeEUjcpDNq56UOWC9sdcWqneK3fxwAHN9H8bathPIb
P4Ll6f9TGSBPiCmFe/Xyne0WCp/pdLDksvoK0cAPO4NXfh23sOIDmy2+fygEl1Xc
ss834y5Pj0ANlisPIepzN1HMsuvg/xVS+VzSZ3A7OE35NuDEke+MIvrgYBnTYfNW
N/HDOtBQ/Qc1VJy9zGFR86qxXF17BbzR84uZf1FTyDeK6TiuJwDAZub44i5a/dRd
v6EEd6kc/dzT+yJS03TXCzn+qcDwGn/i1GMUWSBOjSnvnj+xHlxeG6yBBP1OkMnK
HFBb4mdE4JTvd7i4LvKyCX8Mau8TszBOc0xLwH8Ri6l/Kxx2KHKXR5ZgcajCTiXu
EPSa9fwlibPPm/Oqa8US7SblAu0WLnDNM2vOpLtNKU29Cm+nVdc/3i3tnimXuhto
8pIKDhWxjixJqC/UqiRLpIE2UDo1wBD/50GkZRBRXF9SB/X04EyJ8UtUM+0L1y6x
CYpAdwqMwD8kQHySZuQYKZuC2BU+WBNXzPCG2wbhIaAqEZBYqFchxRSMioC8aN11
EJAnbpgNrZ1qDTdCp33LMezTa9yTNBY+bAuRcQuByjBiaBWN+j/76QnTOqg3b0MQ
HNIWWsUqM/I0zrV3dFGiN8ySMMLVqI+9u1oZQKqXPvS0qnVzK0Z8fTyuJBrLDfa8
TyXQnKn6Mj3kserJfdDmkmgVrweyXhxSPDmG5oKDBbO8T7D5hYoynxTO5iy5V0iw
752+N576Qa82JW0BCK475sdXRxsC7SLVrK8AvS2Y9wGhiLyqprXuCH3DsvbKiwLj
1ThS4ydCKI658b55qCYlFpxfvRWim0waFT7WiT65A7f1UzRHa0kdfTB2co4ovQxS
3fANVoPOnhVl5VwMeDSwRp3LsG34KqNgriht2LZswOOgGw0lhoxq4nCiAPXtHONa
pbD3G6yw/AQ0Z3X5oo//Jv7gJWBoyCxgaI6HKxb7LmjNQTanJPQcRvn5w7K2dJoU
GHRPBqYXdz/6Gqmu092gD06lZEGPGfoVW62PWcM+Ve5YBcODANBGY2pfT65ngjN3
19YOBnXS7EnLmkAmbRDAalBUAe0PQybvXmV/LHKKLeAb6YUAI+M8zDx8wIiY4/d6
+gYT5t5MUXnSKsrM1Z+HHbySwtRuLMHUaUBCigLPiWRYMhL9jFA4H6agk5Nl0+9A
1z5Qq4mouBGXXqEzpR7+6winez5zyZjcYndjdTUHLmaX5IhPEVAGp/sJkcgxLsGt
r98rjMEIUJwYAvdwwyRF2sGjP5X6NXvLqPGL1Ooz+O+/CJn2B1yfzrypZVEvnIiS
NWTDzXTvj1wehgrvBdYIttUCOlpgiXrV5EGdy+f4F2erIrEQyWv7xblpwxpUAyO2
++r+XrqOpv9ed5A2cJMbwYCgmy7lF4AseHku12p8AayziqnFeLiK420K53vc2rBm
tIUf3TsaLIMqiZ6PuFggMhVFqVACvLZK+oZreWpQAFRF1DKrku0fg/upjozUCfyq
N/AMNE/4qIt6YKfJRRRkFBRQm5USnfdVW5ZMnNPSgwAGO1/3F8A0VSrNiLUBxB2r
xGtneqzx4cgUCTzLEJeDBwC06iSSsFAm3mlKSfQyDuNRZquO79/4sTYf98BguV6H
cVI0nEPuFCvPiLElzyt6ROvy4SaVvpZ/v1XvCQ60acEpWrMBr0QtN7uWc3zzA4z3
rBaNQPkXkQh/UnezLwCrnkpEbgRFRzVVWRq2E6SrEYnZLVg1bNXwEedrSpMmgFxs
1E/tgBZI0KWET3vFsicSEAM2+39jSoK5ATRp7HuHzPNzc3cF7ggJ4umcziimQPBk
6DlIQuAwyYDZIGx+J2ihAz2lVnXmA85U5qoe/F/a3WwxvX/behgjsWgJxqF5/JIt
/XbYVuD7t/PLGN8/fJvaJ2ClZ1qCkgW7ChIpwKH+Dsh5Wg3se5GNgWsYtyajB15E
ur6MXvs2kZaPkwkIMmB1pbcXLw0WZ9JzxFwRY3GOtpD/74Y/Qs3vs23Abv5NNJgG
sCTso88r+kd2KYS8OUvn9k0762ASRL6NWCwHTPGmo6YZXvnI9Vmo8pVzk9dSBMpd
692yx3E8DVryFw6IbtcHvS0C0Nw1h9Imp1P9d8y3QWaD7C7rcjzn01UDdo5dCsHj
lK/z2kbbLCr7Mp5pkuMt2KniIuGVnZB1VkAbzaeSrmtYdbx+Tle1bj/qoxT+frYI
4X2IeKi7dBz8XZvaK7LCOodtkv1qw5W8hX2kgKfvcyNFP5TaEYXdqX1Xwll3roc/
1dmRo3whXQspyCKaUH8d0wm1nTt9PJ4yV/qgJdX8NMDv8T5BRt6GPJs+zuzA9/sN
Sp4FwGrQqM7JZ9eaxS0ThMW9YxbH885eFrdR+9jIzfcJMutBos1BMssIPq9cMYT1
QE7znQkUIBu2I68f0F70ArnXAuSYC+BHHIe8ASm2RJKSVU6P5A0rX5L7k61kUDgl
0ALglxkscQbzy65TGgXh21kcIgOfqXWZFnNcsIvrK3RTkrU3pTSMXum3zMNQ/bWm
UThPCoWqYXQMiKd91GckyacwxPNtNSGf2OXrt5fzL5laQRHhqI0l3+SQSrLHc3aQ
AKBxMnNsKLrETeP37NWQlbWzsYqheVu/Bj//Q/MZgYAE6khnNkpAEDZ1RTmkmxi2
wR3za4WLzzXLTnkVmpF/LrQ2h7HsW9a5D4AzgkozxISVGGVXXGqtVsXKvbOkXBl0
y0YRUkxt3CR3oXvkPW3hQX5bCfTRbxwoqULmlbgGt1TkOIJgTRxt3UyOZvN3Gnz+
IfCoXFSRwmOHGy76P+AcK43t+4Qg1rIHN//miXBJm+cxCZbF/y+wiebTEAzkwdLZ
0ivzR3sExBxjcDJe4KnvW0+urSKU2zsY6xxxt6UAO5gcKOigVVS+fefGpKVwxYDi
aJTCiturf0dP2iK1lv/mdVINMiHSIH2PKsZBotoB/ywYkXMOiSv60OZiZzFGHgwx
z5kbuGuIR0Qd21dU8fPVLiUSOf/ePYlfJSOrKgdusqe/g5YBDIy/sgeKEJnKHOQ0
S3zY8rZG+BAuZVw/kuiiSXEW7moXO40EuDKThXVjSAsLisox+vVbNNkuj/kgp0ly
xyKr810S9admfa+AoqjWHyJJ+BZKl/UHXGFDPXB2dmjE6nTx21cTdltdBiPeNzPz
lEB7FvoUDNL8cKu6DkoEFRkaNqG8HOnggCavI1R18I3F7a29L50Qhmbp8wsyW9jn
+OntHLFD1XQkTb23qmp0XqG+D74NcxtJT6NW2UmiKoMktoBnWqfpE7trb0L8A9Ak
wBs17/mafEhiRJ0fgG/OivZTJEf9SS8QlVCPeg94sF6WzJWud7I+Vc9tJqhJR2/u
xiKRV57Th/tDUerTFfyPn2kyJopE+Qi8nyLrNRqFSu+eOkDhgheYbDkRd/QbXtcr
UezZk7I/h0pTi3opZZ6lCno9MYFuOogP8no22g2yJIiAY81ynWuSZqCS1v32TLf4
ndVOnI/NOoYNUPIA4xvs07DpRRNk2dAjcoQLzcxndKmDKihnHIyGl930f1lYtlRn
6QG1v68MPgKTNta6ZOuUWhH9qpaypTOv9eBwVIo342fePC0wNT5AcJXCFdNI93JT
1h1dXNAj44SXruaA6irV0SvHdIO/b6000bUxuadLg5yWujVwlF0+OtWfnpYWQevY
M536cFUeQtJzTniubTuY/LKYOJ74+CryZ7dtv5ZBWerHFcZxllKOuNGVTlNMzNmw
V17vc2OUNo9ZLnUW/sdMwspuj3G6OxiMlB/y2lr/t+m+TXzQ84DldlIiBZXB6OM/
WrGlIBJf8LDjchu1wX3CQnWWF6pfXv1Xj7ZumBP9H0Gd2ZS1YEDnl247a+XLiPSN
mVOtGgnQKWulI0omBaWCtE21OxkQ5bmxtw/OCvXGSz4lzc5/R0PD4SbQXuuMKKs6
nPX3vQoC2E2W8eK7uRlBwNVtZL8VEPk3EKeIclQOAjQz8EShyP8vVszqTKXpfMSD
NYiMWHqHSVkKphnaGHtYBBE7YPhToRQ//We7+9LK8MXyQy+aJ4DAREwi9ecMOGA5
PWauvj8EIK90w0JwyjHyFhv+dSydt5AAc3UQ2g8Svfn6wnqHbnx/Ql4+/NmAQgcB
3axAsuYaubzkA7I7fVib5GTtsHzsTi3rg/exwJZT7FuzzVySFXRBCmabNDabmo0Y
b6ZnekPoEI9OWTHzoPKxNc/i1kVuPBEx0ROwlLRu+VdII3WmcTJvD17lefAsJDkS
9qBvVPOEwmaGeR4B0Hz4GsSfGKRC84gKuuXxw+MBZfqul//XD1Rpvc93jVvfHj/D
CWppjVU8CKCTBILNRq9CGo4LUtTF9aNW47i7rmh83AGR/8B08ALhZFHlgC+auDRl
SjKNyWtvme6kXdr8uo+VMJrVgizS/Oe4XrIv5Ry7cjpkRZcar0BOxv+c/MBsDkU9
NaiSsn8CCfU3DZK7Q0PvzllPtU7PW3phJdf8yxP34gZ6vndIcAosvhLsW9+sWIji
jc6FitevoGxgDR2NfRmZB8QpN0m79nA6Uj1EpGgRT2j2xYAm+wkjG4JS3bwWha8L
k9D9CS0E+EBkq6yVASjn823053lTpxCiykJD72KCBWipZ91YgDQ+cEVjnJTZsCrA
QWX3L4JOg+ulx0YCONmbK773RCFUhQy/JPcnf/491k23fuajBUIzbIJr2uAo8n/P
Ac12FvHhVbVWbaOScrrC4gUfc8+zaAt30cIpqKPW99PMm4oDpdVLd6x63trDx52h
Ib1AnqTSXiIywzyUcEo8Qm1YQYX4imCNJ7XIeCDu5hlnr1q7IXeDd9xBKg31FkEz
MTVE2IcBm7UZ2ntMwAYW4P5L3uKhwaYqimfNpSjZvcxL3DHxAJBtMK1/SDkmsCuK
24K08i8z0EMoyi2tiyr7lhZgOiKbHxwBGH2XF4zqIQrmNZ0R0Ih51G/742d+x9Gz
tiyudH3VOwfQHcPBEEpo6W7RrgP+Xonw9tE01gWSbHgUTEvh47butlWjiMMtx13m
Os45uukYIkgJjTcnzMy4NWrSWNWKnZ1ybCElCBfrOY7+a+LhX6mo1t12hiZyZtmi
Zky73PlsFig7iMszromdbtR6P7+eG/0Hob+cWtMv1l4lL5twhIoYFD3/QG6A+1kN
bVlx1YLM1RMpt01K7SA6haUAoBso2+3BiRfkwHzD5kl7NrsZiJ7lBcUFysF7pcaN
Os926BSjteO85S1vXR8mYQ==
--pragma protect end_data_block
--pragma protect digest_block
Wqa4FfHybsYMFiW42NMOS7JZuW4=
--pragma protect end_digest_block
--pragma protect end_protected
