-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Jo+jwVnH9RNVSNHxvojP5b0ZjEvouLhar8h58puevkhrj+AWNYGAEz9DwwDAbvcD
iR58th9K/tBCS6U8fWp+R1q8N5BotdKxNrbfcDhAjXqU6CdBr09AWi7xr0IHleWM
MvBFdVhg3IufNLvgSV8X3ip6Umz1yyRFooPIbuSQZrw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6048)
`protect data_block
vogIjsHBnxcS9OhxG3Edyvm3mwTNJZLwVWovXITSDhEt73LMTXdgmEBlZrXXY5UB
E0uKh87vwQwMcGNoDDfhg1tzxsXInoCQew01IjIvFBjJb6rkhGWO/L0Na1J7Kt8l
iJuJVSGWMH0fl6TgJCDbIP+rGinOMELkL8zniUMjf4sEA5RiG0flA2u9eZOQozOk
QGxS5lRT0jxwJ4+5TKfm7OF0yICHIL72t1ILQGRu1Rv+/M8O39F8zdG2Yr2yrrs7
wnf4adexMeHspZPFk/qF2DzTcG+DPy//+h5Tb/pP1TcO33xN+Euwd+8MV1Asl9eO
tlwdftC71kWz2mPFuuFiVzmx8NyIWTTlMkZ4ZgD/FkZq43qHlF5ybwB2Q04p2uSw
EL1CT6wZEHbFdVBXiHTa9T/txxf0Vk8lvFbaJJpI36U/kBmBPvMolPLrJgjsOU8+
wGUE/B1sz7813Poi04QM4NsnUv9tqCpuQ9okWKBHZAqB52ni9nSMvTbtyfGnvBMu
YyuytqC2tqjUK4sOewe6kunSWU6QdO3Bs+UxbK9+7/OFhPb14sdXnvP+bDZMeH2O
rEPzSNBE9lZtQM9EtQku345SBzW8kWSI3UbX3oQ1WG8ub7GsxG7Z8fOjsdZeR7BQ
5S6tuYkM4Etwf3Zmj9cg4vk50qQHiG2OISaIjQTeZQMhdsIVX2Qwn6gAsfmUkMjl
bDz4401haNZP+ebljjFL2o+yqmp8/FhnFj6QqOAmWgdkDHi9RjX/QKcr71WAv63w
6hZIaddgKe36La4Y3SrHXPTa+r9FM6K/Jix0PfLOLniGMFtGnnjAL4sKwPUS3e9W
x1QKcKCY+Nj/dYB2Tu60lzQse3onc1DbcEggrMN1sTAD2KKu1txqoZhCvdBjvEXA
JHIhgYFC+E3NFOBe3HpihyxhyFtshcCJzLm766enAsULkCgoH5y65XJwjJ2XZr2s
fePjp8Mnfq5Gktz1O/Jevelz6L+yUnCblzB4o7ghKpyyGl4sprBkoowk4t+JFVxg
APlGkMi3VTmGAFrGM0cKQ3HcUrbfKuk2w1/bjuCKorHOOujfGxMRzEhz8WBV8v0v
mzDc55V0uQW9f4TGI1W7gP8dKkuyBIKLdnhBpoce/zc6ipLQ7xcloIb9tTPL/0UX
Mya6ZCepTcDY1cq7OcXMNoKhWcjDqBTzR75Qd8XcxuY3/BpoT3XkX6eK9HRJMv2+
xoeE9Ayw+l3+8yN4QQSIcR1oNBV9sPfIBLgP2vU8jAeaqRV8u4ZCgBuoj/2jvvx/
0tWDDtMeesd15uH3MFXdsAeei94/wBunG4z+OWexmQ9t7SaD8vWfLJByWYj50tlw
ACtAVhb4J8L/7tdc5QHm216oySpJOEIV5l3GRHGQYx2UMEuu4Gn3zMgTVj0qBMCF
+0HV3znQLeMBFiRmuVD6OBekhISaK9LcLAWVktGE6bbhDf/nL/9RgZk5AHgjEEhP
69ABuxtHBZB8nWbg+SFkDqoozCHfx1yHFvcvquXTqQCzyYcfXRL4i5bDPOGVsqCH
Hwd6rzUUQRbTAiwRaDYtEWQAA/bdgo8URg7V2NPjxJhyZyB/ppylcl+/oMwgc9D+
H/VqiCh/PaNxz3RyxJRmJ40NVQZof1R1V0sze7K8fDPOV7qQaEicjVdGJQXxdFIU
sYI0DzB6kLhEjQwYoyN8uTPgskG9lC5/FGkbx2Bal+BvQJFBgX3rp1m4e7emcXtV
VlXYD+PV3ZlCUWbV2y6eaKmwq4nNKjKU2EuCZl7RVTMYSGo5/glFhhOtnSYFpSJR
r9UynGy5+CDPpsweMAYHf/3xzUE2Qq3TVggXzABuMoqwNULofVb5jeyLbnTWfeAq
st7INtUqe/joGLx+iD2c9gKYfIt2sy9sOTyFCMW1w3Ne80oCdnSehPKkDJVIFFLk
D5kmk/dDCJTiHweo/y1ZPX2EDmr5Llbq/Xks4/X2iXKyCq5rLST/lzxDg/jcnUvg
V5DhuMNOpPoTKAy1dnBRNgXmp5aUdt1P04bH/epvvZD6WyKEC8pGIDmLhurJmC4Q
M9vzB1G6t0ggKhfBUMap1VvsWLhogZfxnzmMtkiNpLMO1ROPHKOdYa6oPImoh+Dq
xNdvCB/kmTDusQNm0tbABNUH8TYoz6LMXTx+n1GLKJwPTGDDKxxNhlm4+GxjK71y
MXCSfkc1C1ZT/mSMbHSLoQf6M2UKuQw7y8NJ+Hi9Mt2odiLs13YgDfIcX5kWBbdz
LbDw5v8njQFEYGn+VgwEE10mTBaBI3g4FeBeJkuM1xiyo5R2rLDsRmXQByRZp+6D
9QMrJ5ENdmjSrpi5zgpI5p9DxEjJopgyEYAzseMtmoqpRWu3sxIn6KWPTX3Iuchl
7rVDlWaWc8Rh3rZgzSJ4nRONf9ZmUgrk99pBysEF6j9RU9my/mM6s7/qFMVG0a0j
7ZBJFfMgIdYnAzgYPxmVLaW1hm8aZRbydixN2Z/IJM+WA0D4I4iWEb3Loc69ibU+
d3x5eTyNzGzqomNr1fibDGs8HQwlD0ZDsQZFgIWDbXRkKkfPJNCumHxzVV4W4gYX
d0ZRVtWqAA6gyc+9+J74hluRnjI8dkyYYgkvFzx/XedBDvpNOsKLWh8Vsp6lA8fj
memCSnSZjf24xw662W+U3bYWDkZT8GXaH7/RpUaPcvFkTVP2Wv3dRXpRQysSw7rQ
SOfrO1sc9Ku9QSZggOKirhmKFfzU9GtK1LGh/4SH4Rlw4DoblU7rcXdRYu2hxAP5
OEUuLLTH0ysjyDm0KTKtX+lA6kTe4QukDn2hDijfS8ojV4OKtMkoInjcb0un1EHq
zkDVuau+FrloZ+nNnlKkhjDJ3mvAFEBGR/TPNwGnLzd1mhEA7hyw1F1HPXHK9uOY
gMZV3Ov1ok5DWBMgSptU490eWR6naMIxbAC4f/6fo32A1DbVAT70TojgoRhAjwS8
B7fGSZc4YEDjLJXhbDnm+85fhoGwi0gtmCN8s5x5Nshp67OMvrtV+JyuuDsGKRDf
owv74CniOayiT2uI7XJKgdrEzGfeKdrO2iItTBD1YlkpBzt1YPtSM2RJxQGHDJo4
3CUvHks99DpkaWB1uvlYtSQtD+6NckaCWjgtJz+jiadhxnau3Z5Tz+CZWuFed0kX
6+/HE1H4QvgjlgJQK6jGh3RTCQ4SydROayJglTrUp8VUrxKj73TFAMTXeKFzwYkb
h365c+h3ISMmeHsP5Y1rJCueFAx3XwatxaELIoKvfCrrIhSmeXWVscBnSGVkqceT
sZgzoisp7L+13Nh29zh15ms9MpYaIszsnpC7NnLAZTJ8jqAetlJBtoEbZ1Pw3D3L
coYXL1H/GwROMtzaZjRPPIIn4hyciC2eaWYYSlErMKTRSytPSO/hv5PKum/rRgi+
HuIzciBJnhJDoXuGk2+LZSWzMbd2AQenWvICIPU9rQayPQgKZEL/S7K6TUnlNP4x
S9sPuuemWEkoIqgcp82tAdSuJMgMdX6dxJ4YXizubvp6FwCYnMOLNSKmrtZYCFm0
L8CsRr7p/GCYoJAIcYq9Dll8MO3+JVobFjBslflGGuqfMOqR424lRpFDhwS+mm2t
BIt5x+FG39G3cYRPbByOVYJJoqZ+HFtzkSWfFjIgkhDzozrFzMgYNbCJlLCOouWM
IQ3DXQ/JWU28ZkG5UjcQLLVbFXKeQSyn6NE+yQSBPxR94Gaq4BaceSWTCeAZBVP8
aZgw6cHdFa6gFL8BBJatT9MvHJIdzt9KrbqHUIEw/uy6jM/Sro3KTbyBljz39rFJ
1K46R/ALLqjxUucY5PZAKUaKbBMh/5St4P65zNDKPRwjbui4iKO4iTxrjgPqUQC1
UDaXyU/jLSNFQ6a3BqtPmjooXloZZDLDuGt1ZxWCxj67aBmz2xuM2yB3hcSgl4l5
F2YL/qBa9HTEEC0RnMT2VAlVMYPuFch81oTXZxZrmORS33VJC0oB8gXckIqs7WbC
rhn4SyEMtsHzI3/i6150q8CuplX0ntNhg//WH/emyHi2SBbWAG2r7OXP2Vx90zRO
PeNk/eJqgFYN+GAWF9yTdG1LC3t4PYwt4cJmndjbZa5FnwrGQY8iXB+eDkPGvxso
a79U6kxZgncYO1e0SEQ1Qg3d5CRzR2ryp+p5tLxS7eQtBXu1rJytoLqaJ473+CvF
0Y3pW4d6yb8Ul7e4PEdCF9mJsjFURgkc4JUjFrLPvQoTujaA1fstSx7mUUTBGvlF
ZTfUmDKaeBLfaO9Dy/je3ye/c7vzdFQADow96RYGf1pQqqzIatIISMNNNTQRK7bQ
fqQfMZsRERT3ZdHchztnLQYASmPLt1s0ey9+6hIzeUX9xJ9HVVx2kJM0hHDQ2OS8
7ngHK1IX9SvONMsRQRzssGYGPWECYc1QBhK1+4nJg0FfxuCDv8NRBLcOyNmcA9pj
1QuU0qwt1y24uUuU6EHE2DaXCHMxicf8FsyyxVbfyNkXdmgo/mbP4Hu/J+7R9EnZ
XMssJ2tE/FQ9YRBoE3a3PqgXMhZAZefVijJqMR07c7JK4jKdBdNq8prRkYt4P83V
I2mS+0EBPbxINeELk7OCIh6V0YsGYLakXP9k4r3o5lo/kMd1qgxNdUsSuJxRQszc
Mr6ajGNwgJwTmwVR5VXvLd+LN5n9cVA2hZ/YBFze/TPK1osqDe1tdEWGfJpx9VvS
oklkMrfe+gcx/24pB2/DWUHmz2d7VFiqIjYXYh9/ptPeIRMa65wSJVjdtyxT7VA7
5yOkgUb67qreszBna1VrDSzlB3MCaeM257WvQgi4vJGb6e1JDz+k8B9FOAfavGPM
OHgmFmgwMBFIYpio31yoDiDQc9Fa4K7OxkUODo78G8Xru2sbEbC+csKvmIcaZNuS
tW43Mm+omwpZXHF6AA84T/ag2orvkJnE2/5tBQEuH0bp1WOTTGz9DR5xEkvdAQdo
zajeTRfCEh1V/OkdgyKo7OOqW7IaRGTXLb4zqRlPyi9sI7GgSkeyFgd+ilZSbdeq
q+x/MvfCBTkaiNO87ICiBav78P0VSo49FMGvzJLWZxNO9pKymJZvc3AQBjVxuTo8
AEzz1Lo8kp54H1x3ROKHGTOuU4YN/rUjjFl0g9l3c8jFjtyrQ3EATl+fgMwKHsHW
GwuEsEUN4NtCqHJ6zRqSztO1Xssbyt3XO/7xaeeuP+B1OrshR7xpcihKMx86NcPQ
cpA6NwZV+CEVN9UVzilIhmONhqAwNI4u4PzbCrYHvLfeGHfqy4V7EXa/MapNYQuY
7Z5nWQWW8SG2kr4a1VqbCkEp0TulmSDcape3NVXW/gmZu5cs/L+afuGE545zWxQ6
CztIehBR9pI8AkOdp6rRksA6BljJ/WhcVgqpJZDZAbSq0X6gorec9eBMOQaKkIGM
USXzQLZPjWTdA8TW70tJkMZAAVVzM3BJCBDfOyWxn5/5hmcLxr3VWOuuWN7/KFJD
3BIv6/ykA8OdUl8aA7AnIjstFYza3PWz3NKI8kYnCD+4XHQbbTvZLWZaq5t1Ql3y
dTxgqSstLyyI6nYnQIZAGweJnyPqXkB7cfGWvmfZvUstO4pUUIRYWN8gquWl2cH4
/F98jycjTus6A8hwKb2hOUpgtugUoo8+Ddt7cgWYO/24vAr5u3vHG68mW4dugUuM
gp9P4UN9dqCGQACRTbl8/oDG+siYunmcdW1WnfMbXAHm+Quu9cFGISM7PFwn05tm
YlEwfuDAbN8W9VEeywcZhB+h2WdMKuf6gr+SrLbPmNVNJLPuA9EtUZxMS4PEKAV8
A5Z5w7is7o0Cej9pOjG9dKCvVrZj89gvJhuonlkySILMyikf3cGDXPjoqAcIPK9s
4y45byHOki3adsbw6Jf0I6i/MkgxIJi96BcqUCUJn7bITrrMevz8Dj5INtmJlqb0
pmpm7bjBqdty0OQlGvSWpmtzTesqTY3gk9j0T0qnpLZVapS6rbZdaOLMRyTrrDkV
NeU27mn5O6mH1M6lFGEOeKK0Lt9m5iezUcCbyHLaQwDtqP3AoDHTGYNGAPunFpTS
y4YAvjFnXoegHSNFSdlLZGCUeDckKXTBXoOuxaIbVqyXI9xPuloHFbZH9x58NNns
BNEMH0+IOMU4Dv9eW/haMOK73f/Gzmfa1WH9AwKNLy///JXLIq/YK+HVRGyeLnPE
Gj1hPl07rySIwfVsNmbjJXUB+gbS5eu1Dlnyn/CDn7tyVHOgo5iWlwd2gfNQyl2d
V45WqFqv/LZcV1W8SO85oEzTeUaPrFEC5Yheao1JpYa1OY9mj5uRzMJxpJXrPn6E
wWOJRMDHCyYtNh9lIxQsepNZXzfEU8GqiGYMAdwXFaBEQGmi++A4bZAKguC0VMQe
u4FEIdN/tzmWu6ZRuqK0b5EqBH8+nxB27kamoUqLmJ9tINFa5qBkQK4DZEZlusZH
Lt5Wy5hBuTnQ5o9+ndAVbBFw0VHQlDdWMuiNdkA639W/bu+jWxRfZtOr9Nk+U0jG
jgrgtI7TeMYm6aa0Ro44CbWm0wrwmkRtA8G/eQA98VgAFqIimWuzC8vZB3USXyI0
HzOBLAsmFMNiMoy/6u2JiB0imnBal8agWbcve7uPXyBsYz1pLh5uNE+4RM+3l1FE
9uXOvI6t8vO7FJC6JdV48qnREARuJcB4loYmiiuDHYB+HvPMGeC60VbBNYTZcRwX
MysiE5g1AZS2V9GKRubejPOiaxhVYRFXSBH56DStPbZ47CiyKhr23d8nPxYbMeVT
IsdBUCGaHCxYbT98lOMj2B/iQ8QHAhUE2ficDNp+ktacwqCUfViT0H5UcY1tvMbH
qh3gYJAMbpkuOa4gvzS+v8konKvGVceeUMTu18B1O1/+a5KQbVvU1uRrxogqTK3m
ngbTYi2LNjyh/6rAjTTDw6+tHALqrIIW8Nh9odvOAj3TGXggKXDcN5DmQJhnCLWK
qfhqO5iA9HWHAyLu3zMXfSQ7SFbRDfFfdJ36Rd2tSjI4w9tuHilnirHsGsRqSeI3
8l31Tcahi4aQlbvlzp7AUSsy7Q0wcAyPekJp7yjMKTM/efr/1HBQE7LxSLIHCo9+
suLkfCdDaLK/1Up8JNl5smgGv4thivnWIYhEyV55onHNQ8y2XVYssCqpWQa8fuAH
G4Cmo8HkKM9D0o1HwhyyY5bDg7AIf7Z1O96iFLneiSVPKtZtRca1V9Mgxap+IkfD
pYkBOBWU8mcs2CiikWxXM1VsIsllFWcPxosvqV2i1rV7xmhxqW3weadPqNTWGwza
uRXegzEsujpQ/el5E7qyiVntcJyrlE9CEIWL6hGFgI3ryXl/bqA0lkpVp+SFPLOm
fP3I6ErVQQrHpsNqvsQPUytKjLsVIhbIrsfXPksMYiUdpK9BIQbkzDgmTl8MmGbL
cWdqbCj7xg1XnRmlKOeWJyuOyHOJ+bif+0dCBuLlXZzzoSfdyhhUUTOPIE/429td
eJiu3r8DnQMgdVZYlhkaA/gK8sXzAZ7+SynkFJtGxk6iKF815KmBhr5NkE8WVLsM
cyBSDqNQy9AIBtf/EtdQV5jeEzyClAweZWzLQjzcD2AbyKbf+cKYA6QPl2S3HHW0
L3nKYM3pXC7fV/ofJwpeCw+MyfG9cpuJJn54/TZSGknPRItneyZfi7qV1iKxHr8x
zKzfAGYarUoOcmz2CH/QldJR5qnudC+D7EGrzQIo/OPLLTBtZsFSRfgtLmqjfWm2
JTfHJKzTEMHlxwjZL4JZanzHb8/XNfBQCJuobesJ65j3v0sJ1CTe8b/luzGZWHFG
unJzCQhpuq23xy/vcXG26IJJvtBeoxPbAfWmRMKWpbnph43YHqYoyNcYLOKY4DAD
BtiBBIe4Qn2aUwpNoDLZ21zgjdgC0VyiI3DsDDq8ZQFk80gORq8mCAXXo+XDPCHm
qawlK+Z6I78pHzxhMEYme0VSi76RonaywFc1JPae4x1D/ovW2WxugV5gEhseivI7
gG0wTBTH6yAvFaP7NydTn5bR6a3VZzHf10zBsuOseZn/Oc47IF2T537yclUWKZ7D
E1m30UM57MaJtxYKUx6MkfX4/2QjeEBqjZYemPcKfvrk5rJkBYAwMSk5fcRFJ3Uu
`protect end_protected
