-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
iTP4nWNBbibPhdt++BLUL4RkGLFcQDSane4WjG3DzY2XgYdiR1JZwdXLGlu1/70q
hkRzULf7WzSgeMXC2gtt3j5QCgdgcxRxEiS8bmAXdWf6jFiA8aI3gc9gGQnTuVP/
zpKtC6xfkg+WsSaRSzWh1krKCqIJV0t8Kn2MOPB9nDA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5104)
`protect data_block
vNzgcCB/TUedaWKg7JGlrtgSf25jOCsAkyd1KqbXmkrrFSt9D9IOw606OMSbimwQ
AM7L0Z3bIg/msZUWc6nad5QIVhEP+hI2MFZq55fMYgYysh2RRFfmOGiU3gXB8t60
/muYUrQhCxUE2SAnuG9LzhGVU1RKHZew/4lPAzn0qQWBJGWqgv++3ta/ejQA86RX
D5TJZMOLkRjzynF7f6wvpOvuMLvr/jmPQA11DKQ3MqDvooYHSoquqmV2lpK0Ef8B
0fDf41LquLRRAO4Elwpqjg+bdOyGsOu7ks2e1+4Qmw7T5qfBCKmtZsWhdYI1TNiO
NigGXm4e1GaoCtEQBd9jQFKdLHvtzPqf87dH4eJaEGCCH+rvO1L/01bxEyJnAnxj
4hLiEb9Nh8Pnc3YiEFfL+XqwiOZe6wQota0Z9/o/4xAmT5IF4uO9npdxvYBSjApr
WIKIGzOwPstCQvwAnrKXg75eALqb00yau0s7q0odxXerz01wNu68tJkAawPYKSqq
KYlgVmAODxJCoQcDEFn1forH4sDc9amHuFKWcJ+q9mzUO+hhw387nLS4db7iyHWz
xKAnx3PwBLGJRrqk9lXZcJXcmNQjwKtLjDUixrdTS502O9TbnAKbkfXj5Bt4sdgk
uW4cYaL+F/LbI3q2h+KjpTZIAsgxfAS66t6eZEGX+t4uFh1kTlRs134Z0UM0qxbp
IFbS7PAWApvQEj3flXb6yGwWuPKQbgO0d58VKDLSkal/vXJJMD79MabVIt+jWs9N
QA7ICsRCoNY46VKFqDYFpYQ44+AO/IJeDdNtDXgz0vo+u93jSnYD4kepyehhJhgr
065Bb0We0dGNZbukfJ95I7iFvKikrOh6qf8yglOUzzuSQRASFzno6bd8GLLHGW5f
ZS5aESrzGSYPWTjeG8p40KNlWqYeJfovXhIq+Km++C6HkXMiVV2kXv0KuVEWLIEP
XsEIvZNR2Bz6yPpJroMmZGNEDp4OQyI8ClyxpJRhsXRvF2lM8VRq+4bwsXYzOXtM
bw57BClsuPGOtdPkh+1C3ojjSs0GTE6rSBYORO3aCBZ/YjVZiXU0NbhcmlomdcGM
ywPGJ8BURHYNo5Uk5d9OJ3kAZZcu6ZeGWnN0A42RpwkocRV7HV7kJ5NPZwIxEo6m
l3hEn+D7gSBky7KKukAnO4IOKXFANAN67frXsCydOLgim1VYLszN0O2s7S89x5zP
HudbERtfRb1+rR43BBWuN/Gqs9pgJP2OERwRZ+Ib06Nrwf0lo5MnqLSqQM7t3V8I
Ec5tslYRywB6pxgRBHrr2S3q3P91RlXLVzPRMSTNqhy36dUy5KaNeMFT5YkJPKEU
5lLvtIZb7iZwjc4LE0glTEPktBOXLF6is4BeqitrFNvIOPOedSs8/eQK7rv83VmF
GswyvAt6G9kLBDB63VHGlaDJxT6n4nRAaZE7edZSbsgKtQN0RQpHNxfUmJ2dj8iS
4ekctOcWaDZIrBvdZtcpv3sKPshlAKtpyiE9EWTLuNelNPcgazOuL+qqKwt040st
omzutoLR2uyWaj5tktPVi11outXM6As1mx2SDquZXzvCqw9gmIOFQ9vg7/aVMBBd
xWE/urbsN1tFLsrpJcNBuJN0Qqv9PXGRMZCk5VyrwJsPJva/wEfPdbxvO57xMd+L
VtE0LMObiJwh8TM31NbwVCN2e5Pd+P+m9P66lR0wOvN2wpii1mAelZpFQ4GlYoir
PPR8T061bzsVg0mcwbFkOH4+0mZVIqGzoIrZYP8AG0oJ+S3YhlxYICy/OscMltGx
5PmbresU4/owqXIZW9kQS3rjxkCqMTxnCa779TwMdA67GsdboM/MT0uOwS6CZb6Y
56pw62+iCc4HH9iBb+EYSCKphoAlOGaMXWtOYMHy3ogPiQMpvzaczwoT5sGP5o57
BBHI10heOxJB4IVq7bup7DjB+urfBMtvWTQLVdnmn7YgyIuhnyaZYcSgiNWkDR/d
bQWepo/XmEWSMiYhR/XcD0IZNKx//0chCphAxfgfYgcdmiy73dhTISpEqPYEa8DB
2MAJGE42cPXpVGZDDm74u/WIGw50227/XZAmYv23Fbq6QtBcXK9mYm3EHYdtMB7Y
QlTMj+PdZS6lIz9asY0oqSKOo26pYeEePrpKseIla3ZfX0JeVgOSKS6u0f6tm3qB
I89WbzAQWg3ic23sgeyEQEo1jJGQwxbeAzT4zSG+x3X5d8rLrsHXB3peZQ7FcBkG
isVrcxRiC3ZudsBx0cVGAbaBWK6tGkgiG7ZKODofTXglzTPf7QSZmka44ROe5scV
7T/d5gm+P6DeVPR4QaF40H/mvFMQVY/uIyiQTJWuo7jCAbUWmI2zlftMfAAQ0Whd
IeJ0pAlNO/Ii7WPDzLT2wn4LM4JPxpzkxB8mLQmOiXG/PdzpI3vNA2M+GGBBEIpd
6djqxqc07ijQhNqlJeLPe37iqkyM75BPvtqCzhveiKKGH+GDI5gwmq7nNUtFOpKe
m4SWR9BtudDZxPlO0hz2KcnLKVgNWFTrKTcQZNby8/KOCfwzPa7zpXpBS/6j9oN+
q6SFoEP46E9rnTXZ6omw0Qs0H7yxXizzIIrKyqA8kvMn3uXtLc9j+OoOukPJzk3e
PL4bVkdSysSxOkUJj1mghTb6zBpYRmXR6NXGn2hNmJwNxgtpelchPTCQ2lgHDQIZ
XScmQv9whsDxfoK8VgodJhMyykRt2h9KNoPHTXX6Ejm6xoXNp2OODDYc4KHo6CYX
6KkWZ7Y+Hm3+huTqN8OT33U9VJrOLwe2f5nRDS/D3WG8+8mt2r7wckIZ/tr3TPde
LIbhJ3oNKe22ak3HQnSTD/+kPmgAFFkF8PajNvKKak02ct+6xoou+KOIFQTsTfa3
oCY3uCfJzHuXT3bFC1IiKeuIaeDV9kqulw3xSUD29R7AwYs2Cq5KLRhlDkTPimVU
uG4+WLGY5XFO7ZgU7ec0Kx0tPOEyQ/wsR/bojhKcJFNMfvLdJYSgQPakwL+HdOBP
PBAk5kM6l0GS2eSfyxojenMiXrItz57Y3Cdvl1BhqdBfY5+HC8x6Nz3rMXQL5UVU
hvM0EkWU6F3XtkHe/xAm84XbGwQRzlGcjXgHGzPiuKZ/LbVjrrSXXdfb4giZIGUP
S7/SQ4sr1XzqnNPZRDp+q75KBp1zg2G9zmi9w5xuUv66J5iVv3Ws6/Yb7FN3G6tj
6aecXRe50WmYMag99kJvItsBGwNC48ub5MquM34vb04l7sHuGRN3VeMLBLdVHvVC
Nuj0nueU1FPcsHpNKFg57xuLVBDY44aRwc0hOoX5zC/Ek8gWdYjuUPSwgP//L6gK
b2wxizUp9QTC/stYXB2sqQrmvTw/3JRUNyTWosTHsdpQ+hWNPgGDlzcDc48dQl+4
+VknARxKnRhUnNpURGD5zVxEHk3/M/+XoRXSOz+wwZ+1bNv0FyuOY7aZ2hV0tD8B
1QyOEWv3X/dps+d6Fcy8tVQpJfqF7DjClWfoYZgb8RFh6kM1O1O0Mv7NKRo/ytuW
QRGcNa1OnDi2SOvDKAAq75/3F2DUitzXfOZD4+C682EY3YtKWZadk+c1umGs52EM
P3YMXq3tAgtBKjlODCO1XcNqa7zrTticp8fQbtxU3S5ctWfNogOPZbDJM98VID68
lCLOYWpq77+98u/ujzoJXu4bao7E/I4mMWcxijpi0EkDeKF0St6zBMWouod+tNXH
M88hL4q88LQ5L/Mh04bGMwvpTE6jLiV66qW2p26drBFw3KgjULeHI01z+nefbPMq
z7m85qt4YjtObCGmyqR/2GbAAwHgBke+JhhumeR2K1KnAEuhLsOTzYonhc2IimVV
8DGOqDNzygczEU/YFwTP+dD42YgocnAvkho4xQbhqjmcyKDkYI3nizdxk69mWb22
n1fBKxLsmrOP/UCSR7F38674HFke7uhcNH1o1919Pp3diiWGVjH+/p7MCdX3tjid
l6nsgRWbtVGQJog54mwQ3MDkD96fqXVH8ulfMYhJaa2e3GjwNF94FNEJu0h8R0I0
szZtZ7kirwyMNU8ZnqAK1MqzUgCZzpuzt9o82gl8lNrqqIdvWdFTRcygLbcCZxJu
dSMjFqdcj3ZYErd+vc8DO2Ad7SrhC+zEp7mU43wuOgYr/F+p3QM8I6YQGMfSOKSS
yP5E4yF+YBBI2YpKg4OlY4J3xeJJuT0LwrPh9jGhQxoAdx6XCgrN/jedsVdJo6X7
gMqordhuihP22AxDbVU/B8MDRxAQX7QJIHt4A/cifcyF4c2tQC/3deu0kLZCHfbK
lsurZNXdStmUAVn3aB4C36iUFb+BlkdksgfV6TPAM0Ap/UArcwnphZp1DFI9mxjI
hsNBk43P5iWNQb7ZNc84l/B8uPtQAy9iXXJNMcdkdk+u8sxWqX5lLMcx/1vBGPIT
8zVOHXcCcj9GSi3pAngTVN7YAvpqe35et7ClhM327WsZV9kA4yqqtW9nJ06/kJqm
mgRSy35H8IOPdy3rVO6Sln64dvbFz7SB1DmZq3Sm4kKGvUF2sPLHqN9bmguM8Zm6
7UJ+bbfKzW93nLsFB1IBa0qFIpyIABEINcEBZpMp533X6obID7OMz9/fTP8B1qlz
EcnxzNl/ND16imiCXv5TIrPBLMvwOpi/zeCRoyOc6wOBcXINvX0Ik20IKVlv9C6D
i3dzznZm7EA/Mn8dMJ1vUD1S/RaECJwsFxoKJLjzeWr3zLqURw7bTIoCogEGN/s3
orO7Sq5M2Dj7zWFOb2mmjkhOnr7EFuYMMcuYIE9kE98aKdthEBD+1V5at6CCvdcW
JqQH8bfcxzQ5PNLD+EidkI2VBkB4PMI1OrloXQqsY9ANHXz8CM9JIe3Akj+L2aYR
A6bSBLu59nQhegqyEbZuGDz04D3x8CV1OTlcnakXEFrzMsjjeWf0VlTJgBv9nFvj
tPYanvq0+WwrC58Xx1wEhBbcBYPi3hhgr/v1F895XJvSOBzWabHCmvESsYEuUEHK
Fq5bM6CzHs+D3+ZtkGFRu5Df0BewRFLdKm3AJr4ny3a58XffWNmWgx3YdMm7ySya
pB2USDlqyRtcEzjX/4dsjzPeNLQFxqJ5GMBxo7uc4ZKxXx+fjImCwh6qujzIlgDw
ua5T5hmcDHjc0pJ83x/lLZpLAnec54Oi8Ovi6Q2lGlNqaDVyiQtG9QcqWgVVKEqy
fzcnLPJmtFLn1ADdCkkiJbra86RiTrnGneANZvoLQU5VgFhLppZC+9CVOv+bmbCI
Shb9Fj0v9a0sEIlY6Kh0ymCeu7OzztcZjsVqGs+tPmJ6eiVINGFuRhjGfYVUDE5D
LrCbo4GFqHn1aDV8Ppo20G499AM5SEfVvYn0PR3cYj/qnpaf3czZQE/6cJiddcE7
30KhUbD7UDcUkJGvYjKfxVxqLOsw2dmkDtrU9pGIjEiypmpZVYkB1JwLJV0oD7Q+
CQ7neamDQHmvXrwmdMAIoH220eYsXEPJaf8fK5wnPnp9wvH1gyKV8f6kCE/6KZFt
z1+hAX2dc05u+UrOPr4Osfvj61WZelsAdYKN6twqjB/eIaz39oobGe+eWjJy/Yqf
smrFwyS4BGqu5gcVcTnHSvNdNzoXPmpzSOkKAzx6TIiUpb6o0/CIqi+ohgT89lfj
VTUO2ZKX8Uo5R7iElnuXqltRmhUqk5GAn/k+5Wc6bEZq9dF99B7Fj6sM3brlZaOo
ggVx43Y0KfaANQX8dtsSP2kxhun9PNNwypqSfR3AKsEbQ/nmqQZeUJU/aAw4QZao
KPwhx79KkfRB8HhWuKA3b3mJ0QgIWPEdRl4dCmZSDnOWAcVDn69uj5+M/eLFoo+1
BbyGJQFKmY2fjltOQv4VgqWL20C8gIltbO4zFYOc03yMkLf05xoAvknyvEt+qJoZ
6OIDBP5z++4M1HGUB969mBhet9DAZxkNNtuGOECZb5APW2qYx+JhPiB59XCX4UBX
FQUdiGursS+DzKm6kQWLvN9cKv1YzH4E7gFtUlzj3sI2kpdZ/3yoDx6ecPRegbb1
Yqy6L5R6ION65E3sinhsVEHsQ3jv3oWXu8Qa1whkSY2UTXTE38YhMHRTv4xW9GZJ
1w90DkxY2WiZ7vEL9FmdAeTx2vAXAwias/KjpvX5LjlIgTpnx6XdI0VAUt3h5MRr
zMM1ldUkc/TbtGAgtLTuifmX8FOBZG+n0TcdztLQNQqNO1CHwkBscQc11YUmsDie
ialv8xRUm/Z44TiEGnn+MscU0Gw9dcuPtj+p3RXAMGUklMjwUwsotxIV10T5FHnD
D39TI82VZOM6ygJXjKR3m6sAQg5G25NLY9QC30J2HTtionDcCX+pbLZjhDq4lnvl
hH9vedG3nMvbub1D3rDi01dlanyRF/LRJoPX8A5BX+gM+onvtCS6jHMy2aQp1Q93
yVT0bQOXmkd7NR79dGpUCn6PNQvucTPBVHXjboRiPQbozxmJhzIRIau7p6PpNebr
Gxrzb6V5MaoiOJea8sSzm4e9SjH1sT8jJ6unu3nz2mYonqopbYGtd5RfydeRwPlN
tNrND4+ImNOhmadNoN3Iod/8jGKK6hK0sFYHnom+raFlqhfYh431ZdazGQmwqnpo
F05l1wwp6qDpxpXt4Aw2d9nc0QJ5AHWLo2N1wZ+07toJIdCDqZXeI4AOopZ0UTUM
T+fvqtJrElusEOE/ZYgE0iYTBUCEfPowE/CgFbzEoo4NtHf0qA/8tMtw7AopDDr1
y/5Efa4lrxr5cFPY5ltXb6WLz12og5nxR9qPGwWUR4gcytGqzqYGp9SwoHhkqy5I
JXz6YmmKbZl8rnPOHKb2uA==
`protect end_protected
