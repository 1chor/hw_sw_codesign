-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
nVj0+IWoODq+4kWdVJAtCUS05G5LTAzIfvWxyfqUNcUHx3NghH4EiWSZojLwBgYL
xltecE9hbEip3gqtsSxVtK3IS38hNQ/CqUxKLv0p2tAFTvYAzHjv1WIZ/R6Y0JGg
6YCSwZHLDOUD2SaZ5zKlV+n/qT58io2qoL1LTv5SgUY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 2888)

`protect DATA_BLOCK
yAECwgaI+rCbJa+gHPGo9tL4PWcfzWAI2f6Ron1L99RbAaVUme0zGqto6Fb5jrop
zw3rcBp6tMOcCa+dHZklvhLTy3vDlMBNuAPf5ct+FN1j1a3CrVSX6QXgMzbwUVKd
a8TYSWrJR92qr+oDka6AS0xt82eqROfuD7RoC8fqYUXNTyKGg3r0JRlS4fHrenrB
oobviW+ykK/qhSF/6XSTOoQYVso7QbiAflMWt7RTZW6kyH0ttRN6wv2DfhqhNqRF
m4Uamqs1W+Pd451XhGNZy2hWtrxwQYUX644DayZOrOW4JhprdZZaiTHTuHaOJYjl
TXJrZqP1g/4IQt4i+8FlsZBlzL5kvsW9y24IIPiGzpdPLhMJwysP5nTJpB1k277z
H/A+BHHbPDxv9+eCiFU5oQxqE2ktYN3BwHlBIfbH01UrPzm9YBFxCFmkrYQef+0O
Za9cWkCI+seGqtIA3YNoqdsGOB9NThdbYSw0SS951SIE1UK1BdxaqaLYrTYGqNsS
VYSC8AXrbglH08659CLgp8HxCYMIiKlW0V7yTqs3OETrvzlkTnZB5EkYl7on4mOj
5n6c0JntenZNMtsKQ+9gAqdC00YesguGSjz+WRBjcPtiHeQ28tr0zVTw20PDLbby
vgtR7aVJ2SNMtt2FdqzMH+UHnIKvrwS1ypiWsP+zq7Gl6kjSpvWFvkMbycuaZuDr
IT8k2AEepQXMw5QO9YbtqldZKP3zxy8Bl+jEU7mCoaM5TntkfWKLYKTAm/6xiS3j
VdcWf1bkc7t04Db7oXHQB/Ra5gsZG8puRnC1mosTOibtidU6pYnMKN6SE2hGJmMD
ehQ+eomuUImxKu30Pl2bBE4yCVB6vEgbu5ILj8GZkqSIfy5xh6eZhcewISMjXpZN
pWA9VpSV4YQNVJF/gtTtID1/h4FpZ/4UjFizxNBs2YqXVwb75VGgvZzCSrr2yYwL
WncnpHrRwViUbkEVq19JEVUiQjWM182DwyzkvMTnp3bgCQvN9mwp2vtOQ0qlGcJj
+mWYy/7eUWEYXJ80mPXVHr//J9tbv8bY3qVqi7UOTrtv6LeiYJmOrIyNd0OP4M1t
XC5mqos//VjsSnIbmbEsMm5D0wWOrqUzfP28zb/lzTY1OBuUjy4LQXQlPKkSWNSa
7nJGjskH/gUQhAw+wAF3914QkHXXErDjTHsIVqOnHgzoRduQLDi2tRNhsahQSN56
fOyUSFcChIoLHbccP7IYPloLdmnCiXB5UYmbYn6LZsJHLcm3leIawKeRCZUKTpYw
FC3cMygJimAcj0bXiIC7CA7XzspNTfz8Wxd295g+oUcBjjxVngJHEiNxjWcVUVkD
Pmy9lI/OXB7017r5NqHoq4fqCUsBbeHjU0D8JUMMmT3155MNnjyFaW4klIxKzy93
WB3yWVa1Z9egBeqY/HVCkB80lXtkPCYwe6suK02GUNsK1swwzeScA9kRnf041nZ5
95LV9n7K5MMjVYcbqIdLIlfaNiH+hhPiFWypLY4AWxUfuTgnShkbZ3tnq1er3664
r5HsnpTeZPG7fq3/6wCjCdssb9rgrlUeNpnRP7CD9jCszHS9OWUAV6A1DRjcfR7w
3yv9luJk09oRQWqf8Qwyq6lPH4xU9H4SQYfHS5TBXzie3ET7lo4dL91uDyOG/8hv
hNrhGSWDLPxHEG3h6vFDM5qMU5+DFDE5RQp8yHGSCxowDeOtOvKofnIuUhQ6S5V/
HI/SPzLhE38frz9lD6hiQsjFX68/13FcbwbHMjuVQsADm52tbBZPl8pJuol4WwEA
T0Ci/LR7An+cZi/e4LI22WiBRbWwX1cq5aMmf3TmAHCZNCFSaY8hVpqfgVJbz+Q0
VfdUIvc4+RD+MVurXPMdhLXKBwlViKKZyBFwweV4U7l7k2043ACQpH+X56W+RMOE
gmkA8Q6u2ZY7mTwXbiYsEHFYBNuRzf7Ak1oeCIdyavERzRHWDol1r1SdXlxuvZNe
kWECkZB9KCi8C6k9xPfpKxq0urxcFgWFbM2Rp8EEKG578CAS/iZvdO50r8xhAovd
i/Pvv3UH8cqL2xkwpo+dqvjdfIe5jUN2xjdAqP0vGLvJn+iOY3nvAaj413QveO29
j3R14SBbt/LgVt+zkHIJqak4e83TtI1dHULBo6QcgAlknWCARegV0Fz9ZqWjlwni
3ghiul8g3KKtdJj+kC8C90YOXvL4xXfGvLJ1jRa8Ssg8h7H+Z07FwQrw/QX9xpvn
TZWZZ4XXZtE8qSGcUfA66zuu8vftAt/A6myZbhdUw8T4QEUmjqtr9Kq7vaVDbK8Q
8RQrJokt2skB69yQFJnzWoaEYTUzn7aYcDiTyJr6/R0VdD/dc/YBAfpE/NBnoGEL
XXYq70t0qP1FYWZ8egFSrTy3EMc2+7XGS6h+Iw2oGpNrTRdWlbsFRGvW1cpUO+iI
Z7/HiPCt/XYAP5px/QHhIYJEIv2m7n3qJLNSm9CRQUtWBxRXp72n3vvCd7Q9swm3
9/CA2voyPSV9wZLvcDjs4p1AfwjAWb/G8/FSxKgxbZNwsfBl6ZrF46ZXIpJOcfNl
v7wWQGDFvNg9Pso5FhodDxk5WQ9EMHMrIaFfRR1GDRk9Wzh7rVzrN8TVv4H0LXqg
LTufYnb6Hd5Lsc1iB+RYKZwU/YNJMkXA+S+aeV93NqhXsM16f2PGaavlH4r0p737
JpaqS+teiRtF5rws7eY+ItvmKYcgc77YwOjfKFQODA9V7RgP/FzOP888G6NqFQul
Obu0Ccbib+9UsqU0Qq2SIgG92AOXSRpRJhmOubclVZq1kmm3HJGpBrGx1YYR4iTs
RWKvwYq7oL9wSWBCNDlv0rvVB4JceN7siIrmm/ZZ104Utjlm1QYTrFKl5k0UH86G
T9n1h0ZwD7JwuenjxabRdogKaFxczzfdfZA3FOs3PuuCAN1WAgZPApsEe+mDPgIW
HSJoivtBipJ2o0jOXOE+WBEcM3CCydZeqHX55sCIMOpmDA6PG1yyjs543KG5905z
yAvE+kQtWLbnhGTNQLYjwwhO/XwwGop4nytO3vwSRqwW7kbaKIYsQZS1vSx7kDSI
i9IYBqw+I41NW2miaTMD8LZyaxTDf7hxhGAqxIkrl+uNdSGmv6RGmm9E6Nou79W1
+m94UPSNQR4pTJAylG+z/bmI9T7sTee8nH7lrJlYuYxOyJszPux0iNP7TQLQndy/
yeuY4kdvkov6rOKxKq8pjs4VFHoJeuJ6JTzdAAjRp9fl3cLqlZR51hUj3Z8N//7A
G7qbKG+867zaPaRpfKmsCeZcwKSUIDvIZGwpCKQur8EMZ197r1fPpeVDmcqqxwiH
4Rb6IFbpuLZ8rhXZs0t78R5sUz4Ac9U8YKsEcZwF0b+g8bWP84KAV69aYOMZ/q0Q
tslljX61P8avvkRSJseHT0R1+oFkbqDl33wqUT/OxR9BpGBclQOo66qZpZGWGDeR
TzhL5skR9arq8/171dZ+1nq8rmqRfiO01KDKn26fSYeJci24McP1BOpYgv58ufHo
0QaPkZAhTs1VpTVtAqgR2BqAMbtqrxdahbKZuqEVSyb8Bp8A8xL/D4CZ9YXcme40
YomQSPEzSPOWQuwbuDVPDVblB7PFiyfpjuqF9ObJiwxUM9bonTlKkSjqodeudNN+
MdwlPqxmZENz704VWObfaiU7CNPK/9+lKTNYObv2dQLUsj26rTDAuJChVFHYB+wx
LjVZlDEshayjoM6+WghdqDIUy4HeRBRdO7hj6yxqF07SLqHOPL4VcsBK+yPQOmec
A8xnnAgLHCvhGKDXYUukkjy6vIK+V6nw/8uTq6lc0yUZVbL0+GGYI9Hxvtr4bQ1e
KhSPN/g/3n+ccnNPY71KS+IXNLQYopVDW2XwldBcx2Y=
`protect END_PROTECTED