-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xu3Q6JxE95KEzbuOYOat3MilkoXQKcEx0SF0QEjQTUebpKxg6bINf60XUz23rbldQxMxU52IbIyS
b0YpDZUJ+Ww/A0x1RBM8D6X53B5b702vVQPrsKHYCWH/o9Q+YjnqBKzt5xImTprng2pbWeJTcA40
zNRpj+IEJB1/K9sLJJvYpod+9rJUfy2asPNt9S7SfiVtZOEbtp7VZbmyN5IM3Tbz0NO06atVRxdU
8eXALVUFOTAh9XeS5Q21nPCLq19D9gtlXb65Mg4V1HoL0GDHLN21M1vZCE5BRyHNeFfPex4l0E/v
8/kpE3JVK/veRRnxPVdukptTFZATXLTTyD+p7w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8624)
`protect data_block
a2cUtAYWMb5AuNanYWD38dH5IPXQ/XGeSvgDnfnNRy2cwRSFH3P8Y9M2Vh6ry12q5NO9UyUaS00X
DJ0ITj54w92fqJN2VWYY64oZeLHRg+55WHVGneKWXW3jcqeqQ43CmRfXlgKeYSWpzUXHNrkYxhdn
mUi8PvdRkJBiGgFy5uZj+srtb5rSsoF9ZhLGmBVZeKvE8Qtm4i9io5OYBVTzdWBP/QXOlG1GX4EK
hFISY6ECUUIVM8lJImlM/tLvgtB1xWId4bQtbWtbaYIPV3X+Zv9NTIvCQPQ69TgqtttcULbkO8N9
anAJ2Pua8bXVfJKLiOMzgfQtpOD7oVCTweDqNlXaCmCGCKWKkXgLnmcamLLA0wJ1iqXpv3gd6dT4
h1hATXGAbAiQB190sdgy/uwYe1OSQFuAGs2zENry1m+/ozzk1qwCbKpXknUJljgKmrx18bJZ9b6F
FUE64nJT9Y0HaFwww0Z0PWODC5oUheIJvvgM2OUDSxORsF9CdZdDyuu2ltUOtaqdi6sG3TyjwoWU
5mfEA0mxFWYhkxngpd/VxGkufrMb3F7vbUjW9Z9BluPg6mGHieDogqQSZcnMOInab6JBSdBcKmYU
ghpa58y8nfsA5TL7a2a8iiwcoM1q6DawS+TaZ24b9o30+T0MCZAr5bQQYOrNUhldwUgSRf6bHqdt
LvRGy/Tb701rcbWQZNFvWnxBGmR19j77mXRC8V36t6rFu4DWup2Z3YRBlUK6uXSdtdg9+AKh7hKd
DK2VxQu8nkyyCh4ZMDHdxDy3VjaGr+zqCzsAN9+lE/ySXs9fLpZFhBQ4TSMIdeebH0b+mb3kzPug
9TYju3zQeTkOTARO3vLS9D1Cii+K+uwCfmknsX7YeeNlcEEJQ+DP3G3n0Ajzz5r0e6THYfRa75LZ
4SfyFvjHytN2EhtGk3+z1JheHJuHCpVX6ydDVEY4Pzjj1m4vGKbVXcaMqwBzVzHGmFtisQtYf7Qe
tp+3LXW01Y7vmoCkRs2zJP7xtibWYeSSw+zXN/FLLnQ5m8nhSJcaFSOAxtZieVuVlZ/nFVpVvtvK
KK0jFaEIvvDW0qIZ4cf1pl4Ebs2CtCRFe5aEnjhugeiVAFxs3k/kFhlNcyh9Xw+6r/vba6Mpc5uB
yhGR+r7NA7sfewFgSfjR7iK11bSsrCU0yLPankjvIqeF42NOCThhMD0ce8tcrzojWfmYSncqYhV0
5LvvPp5RsFR1v2uhQjR9oNZ2phoGDe138yKmm4zpVwnOJzLYv/+czMBvPn4gObBZ29m2y9McZvA0
ewxliQ0HWRQ+GayJM/jYuPN19jjRGxBYk0gMSiNBT9NPsU+GtgJCTx16V80g9/al4tUxnX2IrExs
23SkWpkvE2jc6tiHMa4/uKd1al5Ef+yfNP3dtd+71cdrSjNbYwDl/6oH7FVmRodcL2Qg0tSxU4e8
ofJrTh/Q57WfOTl+vEP/YnK2chLu/2ZDnDzXkkWMZk0uLbNCo4FQDOYzV8mLcQW70RhdF+VhZE4c
F0Cp8dzIRoynFB8V8Dzt10iFMj/GNa7nyppPSR02SO50QXe7ddn1HI/Jfo34xMh0h08uozQ/f/yt
pT/ZnDRldY+ivpge2B2mCniK/6fDT1y5QDklqgh9OxDCB8ST4KdQuNl/qcPNz62Jy7NYJXfVKcso
C7BaaOndcArPkDhaTddmO+fvCo9L1+tyk7zzo8qQXnUXBBAoQTk9HiU9RWInUlaXM5mCHyMftcc+
nqgIQk6ARmaxl3ZdNXAra9uIpVXzBYnOEWS4pPvJyBF8vrm94JK7NTSXykvML4xapcRdAhCr/OoP
Zc62cdpStMVzvUHemL9M5DzreKPz7mQRyXTzcWehSFfWQqTW9ZgJjV9hI0FieDDTXxgGBvyuoURn
etbJhC2S2VHlL+qdGriSSJesOITA5HGKQ5OSjmsZaaUisjr6mB+lJCAZZyaJiIlhxOTyli3DHIhV
iL16OqBJz/F8fbPPYxeJ7vr80Z3/BKZKyXpE964gVtNH+K5lN5TDI610G6NQAARCI/nxVv2TZLiG
GA0J82AJQWrpGSLXsuLwuNVjwk4itmgvckrfQG1DCN6v+VYKiLAlsMfZYTOg6hO/zRAEXTycIzWh
BgN0ybElH4D+j3HkoRrvLatbGfH9OQqoMrPQPpfsby9dks5hRcdCgnYgJeLp8LLEkTYIKJRmQp3i
gS/z/g/OGZKB4uhrIvNVwPqRhkh31Kt5if/mMQc5QRbro50WnHB5pHukc9pU5xaXhgMk40Y8r5yn
mKGM+iaA5UorGwrTfVoqTh6ENtMCcAgccFuEjpcFstWhon47ZaopC+N2bHY4W2j0fmw3NnPeMU2w
r4EK3pFJgG/W1cV28WQW+l90MOMQNlSGN9uhalnqRFzzdYAD4uOnmCPsFQa6WCH1vrB1VtnLwQ5i
lkUShOwC5+LHNgDLh2PmHVH2hJea8jtmy+OQW7D5yWLZ/OMtKdJLYB1ysbZrZVXBQclfqJhKK0id
rdd5aHqbfTx5J9dPE4cE8E9HRjKX+Tsj3qY7S8RzWFnYZ263aJpkPX2pbwltdJfP5Qf7PWEwycSt
fKGt2ZrICnH2IQUal3v3Wav/cfW1vQuwU1T8/b3YirSdbEkAJrV/AN6kKd1i84cR7NChEoFbwOZ5
ijBtm9Pd846l31+EPijVbnDbkQoXxVWXJ+LDAGYs9rT4cF7z4b9exhvNVDjPMUWQHhfr5Wxyl6cG
wlTbYJLF9eMVb/je+hXfX3ypaU9+yoD30AJJbKRoiwnj100ZyNLFU4PC3MuosYcVtgngPPt7okUx
KMd8kQ7dUFKk2kYeAxR4eE3Uik2hsVzp/lZtsR+15Mibi9Qbo/QFN2cFYo+llRHamT/l6E+DIxHt
b89pcUdvM6UiHWxhD1L4jlWGWCKciyuVobT9iOUen7aaWGi4ZGIRvCJ0qwJtSLPTTSaTjdrrg4ds
zunj7O6nG155i+jYocACjB7LQEm7o9EreM1hWFNQg9BKlTzu+RvoqpUdUllXy/4J3bqn1yxGdCYM
m18WuIn1qMYv3LSQr+uClb0PkcXWDUMxhNlKKXsSX7wTXYo4nIhUgRCWIhPhi2rPstDQDgku+FEu
NPZnIhNhA5PvwPsL+cW4de6j0/ZbLvUh+hmRsn1u0Bw9LQTjLutWAZXfCEGJHsvy2yqF3lOdmTpQ
JtEoczApInqqJUvgmGJq3U/8+4WMt2IX5pa+ggTZ3fneBOuC28oOrNBpnPYF6gymK8PM1RmMTOdu
22jLqVyrdmj53/Z5tbdcCzKe7cXVJ7Ae2rrlxjUgo4zcoOUxX2b6BK9xlKlcj/I12TP9YbDZp00q
3OaBsCPq9+Uyu8fWfUx7MUc93Lo6hDPPDdAF7vbnaAW1vI6POpL7ZgyRrxDkH2w8C9IsT1AErWU3
PmAqgp5MnAYxWk/6Gq4TpchKCnbwBWB6rmFmSrz7E6Q24L3XlZra4T4gFnTtWrpO5GCzCEyMnibI
e4i2Gz3sJQsOeVegM974BEbDApgjxSssWaJkVdYPH3diPaxcm0jhO7wGtWWTSwKW7rBqcUOHRB92
X/ne0ADFo6uIJOLZTTQFfy45/IctyX6zRitdhiZRSnxvmZHNXrF6CgLQVbp0p/I+cpHqrRQaARCD
EVoNoCvYhiF7heOt3FG1YqH1UnQ6p8ktXY048YQHa3y3eZCtuAv9fGbySQePraAMnXSt5IdDLEW9
TV+KuM7xhvYMd14F/x+zMq2B3d8bBrd9KoCzJ59PkK3CU6x6+2JnzxWO8lLCp0I8MC3ZyXI/rVBy
3C39r9C1A4Fh1Z8KyH8IqCzMdRDi9M+qG4f1t9UiXVEBNH+TNvUdd2iMeyutIXVwfkdxL80J+ILj
Y2o0khwLlseATIWPB+SoZtoFWJu1AH1D03GtnuN/7xAx4gjxErqayR2Ijh/1RDyfc3b5q4TsaB0c
b1Qd0vTfR/w6+BF7D1jDQZ+bp6FsXbLXS16iKRVSdHB3ijewgYJ51YpH+4ak28RM9fhBG72dVwKk
+LMwhwbLGqfItdK9pEJByCx5wmEvGZ3u03osRAP0x6txreejzlohVqQRTRyUevTxi7E31q2ETzmk
aMBTbIizNuvjkQNQsMEKyu7X83CaXNhXQQlbRSDXmycdOsutuU5fTnK7GddpCrxyk+nXSPdNdA9C
T1xU9vOPYLzjSmRRAJLphHDUPLVpx2ayI+vMSOnR+YEiSh2kNuB6GuhQMYyl/c3UTcu/RBXarfq1
rAV8tI95q9U2hp68NcTSoUMWw6aCO10sQa1qG2+yQjnWzAd9TXa/X9qT3SxjVE3kPYtP1OnCDLEM
/6Up3yMUU8o33OhUbbnnSSEreQ2lvpNeHskk6y1Ath1lzB3j/cDH0J4atUaxaiPl9Zb7EFDaphCH
XoXp+v/QFwp+jIsrfTXGfHvkY+f+09BFWptRKZs0oz/AQcFmWdnQG0cymoJYe9nLtIE01k41sfQW
r2REIApjZreHxP5GyfZJZS5SEUfexjXPdlrqXLrbNffPAUbiFPnDsTJxv5lISpUr1uXn+5pWLynZ
7QT9OfeDTRMmT9ornZ9qTXmtDPIEE4VyZS6uqoavIHZkfDhG0ryjEXYpx2/LdOS2k1ZHt3s79mQ5
EvS3AbRpEHAw9+p8CWWo32+GlrukMfJb62NwyvZa0w7Mbql3D8S70n4LPffbtMrtxGfrgkKhEGcb
6t8f8FHMU8FeLS+zMngxltKqzszG1BaGaLf0Gx5CQ+CkbIly2MJsZj9IFCW3H2nbuMWKXEX89HYt
gRkVT8cSGY00ujtuEsl++tcyj7uMSs0O12IdwkZH2SXnXuo5r0Zlij3e+MMEkutFONl0f9lcKET+
asr+B2bDAsdMuc3+ucS2qU6z7zN6IjZQddAkvBRiyuQ9Qs1fvoxURFlExdBpQnTeeYy1sAvEIuzV
MQw8Zh9HFRJ6l9w97hKMZccdRAmN3w5UdS6OMKmJ2PcPe4tGpTmUc46of/izLf743xQb+KRhkV/J
ODKET2Juo9BtgoV5FLJ+ofF6cQgYhv6tbnPCbP4wLVgFIQXi1oUXtS6zaNcwUJN6VXwFLvGM8ipE
9LlnaNXOAtsRzyd5LAg7lc6kQNuF3MLuHlWEvZQ0VXItUO73M1WqfJ3Oipk47N+n498pdeRaywQQ
nx5m2qXY1XIseeyteRf3qew5tORpOU/bAE+yPoqZ23zH+pQ8gI6ZvY42d36dsBFr74F7LQ3cLK+J
RT9e/5eTy8E5AtriUMdAML8qniKairzVBHr/3X2YREsZLlqwVWVeJp8mHvyhjUTDHNLvsc4YQAzV
xao7Af6mck2VFNANQi9XOhbd17cJ9WEWrM0W7Zw6NwrjbjRf5jh5FrqllDsA03yhoH1GKucPJgr1
juMm9nE2VA7vLyRMLuHR33+VGS2YZGxQAJsT/hv50wXgW0OD9sjXGqYpwi9wTV9RrN6RbVM+4mDp
qIsUqHFXUP25yzFAzTtX/GG9mbZGNuHki1Pxc1Hz5CnX2x+9sB5KImFXzWrW6raXz/f7Vj5WVNAj
RUgwedt3EEcCsayVCxEQ0ILJL9UmLT4QLheemX4fMWOKNT1SDkzFrJLARvRajYjFPrP924fHZV0t
VBO+kuy/tyLNOpvWC8zZseiyLBPg53VHyTKvOh9ZwboUHjEBYEpbx1s2W/VJGfmBMdgPlqjZFcZN
hj5O5UeaSmQdztKUac9pMZ58MWnoBov22JA+CcfxcWk9XGjgXeOJ0E5htkFkXLXpR1ywduAw9aZ4
PMoDZqf0Fizrw6FnKKqJPz7oWcKAG2v/SDB0+HkJGqc2d4guNZNgF6Xnzsp1Uve0U59X+zfw36h+
4p8qMaM2UWdz2MRb1qxD4OdlM4HuMcNrO3WoCQrJzoAluOyCOKa8R276GYwDGrcEurYQT+8VBFLt
65Ykq3oYn4FQ+v4t6pkwP1RW8uGacJvGoILQoWKGze7usNcEOuu8SKmwj7b5jus/oI9QrVLz0asR
0j4ujRmQi3BAlEj84P5MicTW6s0h6Hwg3WgXGCyy4jegbo5scxaip07A6vTAqB0Iv3rLZ1R4qPdK
TKsmLWzQh/2TvazuRKLYJXGT03IxNHIUX44Afot5LQQ4bO2zWe0xD2EZTmBs6Ap00Z8YD+FyxOT1
GJ3qK1L2k32ENsGYbMfT5f9X4GJq9PT5mzGnDjJ54QrYhZCxGbMvh6HMUNhYp5KR0tpTcACIH6lh
pTptBRK3ApijWRkI6G0W8LQUSBMmuvMwAhLanE9Nrvj4E0y5Oq8ftSbPICA00xUgUcx9443CPSCC
Dns7sXVJ23dqokItGQoG3EecHUIXc+MackYdUO6CEnP/dHZZVmDixAAh2oOxCJl1glrMbmrhkxjF
cYS+ZYIqyOzsX/RBuRfd92avN+R1b1LC+asdLmcLFHRU5EAEfs7+1Rx4wHsjaO0+Uf0Fm7kBFLhm
Az+qAKPwUb9sl58VHsgncWIkt33YRtywNsHbBzwPU2zYOBLUlQRNE7QOQ7dfIPkCTmu87LD158ah
rd4TpUP4BhGVBIg7g/Z9qzND8oLEp2ZidUw6XRBPg4B/6qEz0KTovT0dpf2RaawALYDrM7ojRKZm
FaesJ+JbBLNpxfCA3/Or8BUqjMybH4s+TbSx1ux9/iZPjxjcSIQC/wBy2j+hAs3frW4WHYa8HHe8
mQ+2/b+/RnzpGRsGsyLE2Y0yrhfmYqFDpAwAZsW3GFq6YRCmcaT9d6U2CH9IloUUybnwAJSLdNP1
Mq/k29gL2GmgeWBdoYphLGau4Yu9/3lQMVw3oSw33fozbPbaz1Zx9iUnvrX814qmtSqk0exLbHEM
XVU3qpS5QqpBQB6JYCOe87scvYKH6cnjfJSlgH/ZinzONLiQJVL31Uiv7hiWNd2iqqGTodOKl7ZK
hnQ43TssFIchzEP8ipvNSX/7qawpSflNstZrAaj14XiQf4nrjzrcIqMjZZqTso8guU+NiS5L8vSB
IOFOzevgFDcky2U3JZIWkICG40C5QQwOVnn9nDJEHJExLOyB/rmT3wBmOHobV1Fob2w1MdBFcsu5
voX0XlmqbYCny8+AkDG8kJlS968QVWSfPlFW8g+oMiVb0RgCcHExZQyOBSCNTjUPJlSf7cUhkx47
RH0q9jNE3wavMx0Oo8MisdpKl/7TtTcGSMjCVmUUHzA8WDaPUahq0hit5QWlROxj2y2tkuDE2Hjd
CPNDQ9yZpHsJUvAt+cPTUSMta7IJYh7zAMOFBLJ1DJJUbZ6fr+FD74DeXCdex9U0cb5EdONlz1ni
lPUDYreCk+I6K78Rvjq02JvYmvEOiA0TzjAkUU75VCFV558/BHerfvzasH21K2Xx266VAsSRUAxA
DqBaq6QrhnGd6faZHymX6xjzm9pn3JvCCPnUir7gM8D/7uG2M3xzWOTyD5HcBHJ2wbOrQ7ZKHu0O
6AyVaDU9wRahpDTbfE1N03Scw3cenZsS0IrReh7aZwt4eMLX96XfyqK6zU5xPFgrpb2J7B8nQQLh
YwiB7NdjtpkVRBukl7AZsv5R20LXRu1xBgZplZs+HfQGF6/I4zTXjGeeo5mnUW6l3JnMjqQi3zu9
iOmmmHAe/SZjQ3tU7QuWpa2mHJDILl3kTonl/GaboA9Z8PS8L2lkITvtXpeyoIOO7UUdDX13Wgwb
JR/6/s8aqdNDMDwd9DnbkHiv2WWRIT26NAXey382X3fzIpcxb7/5rD4pvouSOJBuEoRjyPxk1sSE
MZcIOp6ob5/G+GUxZXN25wmBj8Z7yQtwvqUpgoot6ok5s90lPFetoZOwnyAw9BerPCr2vHDzvKu6
NfPZME+6XCuM8OK02ErUHhJrDHoEk3BmVJ8I3TdL5bUza0WZ1u/by1oO9uSgX9FrrTOfnWqG1eh3
+fIoHbQaisZvUDdDsLDDpa0ZRdmYQ+xWFkROXSiAT/W6cpTa/trIO8LhvDuimcJyIy2jpjqKDlPO
bBj7BqVmKAN5yOPvWHKj8z+TpRdyxkqjwz967VnnD/XCo50eQDbhH+dQjvd25Vxp5uvBdcTbT8JK
FlIAUthctVpQJPT2LLx42WGoU9j8Ys8NIjoYiPYfDbywG+jiwubEXFI4JJTGyQpVps6RrbbdqiCu
rhIO9M2x0re8aCrbDPY0EgRa3hMZ0MYwE5MmXzb0TMJylkwjjtgmCgPi4f9IBAHBqjeQrrU0HVLB
7qLGZVABD9/fQxPilrV7bL2/Gcs2FdSq+ZKADlDHLX2KFyoqI8fzMm+b7cLKUrkhVa6rsRf6LPfq
8Pcby4RYFlhvWbFGbIa3FqRDLmJmXjM46V8eYRqzP1AE3ssx3XEeiezSGpah5BYhfmG3ThJcu/Sa
Uk71a/tJ+/mpO0Pg1rB71l5DIbG+ZXem/H9Elbcg2+xZEYY+22TTbsREZSE3ESDLd+6amm4xw527
525sLBIaHD9RQ00VHMBHe3mi41a80cfb2WshdJ3lfph6wDe80SyVFSAQSb7nUYYeXt936Gxnh1uS
Ow6XEcfV9X0XGHihFLhmLtf2FZnFVLQgnFOCpJYxHb1G0jFOg9BNOxWQwUqoSGi4wy6FHY/op4+5
DcpGgnxu1dWj/e4EIIH3e3iNfH9ONL2E1HyVUqDbSJA57WcSbPymD+Q1GhwMJ8sFayx9G9gzrN7I
iybJa6nISx5ZFtkR5MijDp2PfsuB5Cm/hnCrk9KHn0kWvjC0rZWmzzNOnw3TZPrMlKqpwfOKqlmq
HLgDIGUP+eCiqz+c0ovhk2bHy9cRuouILZYG+tfedtWnIDqL6fAblUWYjLA0S1vK0zYQwezkjIm0
oHqfYDolx2DfJR89dpkigzacC+mpyBdrBBXURDOjcqU/JBVidGlGd2GkvYdW8IctWuuRlHVS57Xb
AcDdZcLSF4j7K+vS4w4fRMn1bhcYWPGOTIcEGGs5/Ijnx/iPVGcYW5+OkSutJPdHDbzs7KPAzy3f
cRRwNhSUfRxN+l42iaj398puufKvEConR50QHvt/qjo59sJOZKb+3qUcPmdOHZrbCpEGU4hraMJv
NYcZpUk3EAGEnCFT3og4DPWB4EvM0hjDRk4E4dHwCEeyPxP7ClN4OkgyRZ+xsudsfti/JMLDMkjf
rA7u9uO8sfHLpskMqOYnvGoILXyC/eiP6q2e7da1oQ5OfK7IVh1foFbjD2E01wgZ1WmdydCRSHY4
WSAQ6Wxo8wU1DmEjrsEDKLHSDC8L4bBx/ojJQ+4A5Vg0ZEs41VZQ5aTiAy9Y2G5D/CtLAK/eJns+
KMWInsxhckmMcXSzWLWxEErR8sVf/yX6MNKIm9JnXjkdFON13RrsrNiDgm7y5zGrHIg844GQFo9O
uqD4dVtsDkMJ9zXJNPka57WIuaZzcGpwpVkFXAWawt3s4SkPCxTVFzDfcnntHqwbR6gD+dNyYjRb
W5J9qrwSgicuvif4Mj0jc3w6XBTZzJjVhWHeihVId9yWyLjh3ma/Sx1Uuz7v832VrbVbZYc/DcMc
Ri//zBIk/6oiaMnIHdHt1eJ+5HWW2M27GoV30/UiODYNFGKXsDqE/LFpGP8M9jTy8tfVRlWxKrzl
FPhl7asKfDWEUYRa3VCTAwHIIlmGPmzYlYfrZ0KWgqJz6VJM8zPRl6S+kGoUoCd4r3dt+jcIPWMw
Fy3UHqeGiIUw4IFp55FET76MuSUKLUn4WjzrqxbMDwifPyv4SRNB4gXfTAeiGtKmSDRPljl0HCXY
zpihp2QQfUY81Jw13klybMNhvVxEBrWrBh1Xw6+2gVv5zMAW3I5i4ziyE/5gyvMT1+s/pJHgQZsJ
hLidDP0rWKxLH2psV+74S/PsDf88dxRPr8IdLhuMG1tJBCuA2FJj/NswXi5z+5LPM0p8+MlWTV5p
xAC+MYZb3GTMjmDwcSiuFjv74COFt9PB66KYu7zYRi+TF5RIJw1uFh+SuPwYzNevxvonHtUyYjW1
B+cva+mvDk6GPEgo2jMSDUly9qYwh1F3WggIbiKcEb/7kEw0xqx/OWb1368lWUlco4FjaEyfmaFa
dKDB14QDi9uK+1bOqaWgSRlqS3hqVnorg65ZcN32aYbmqhgdycMSbZV11Yklc73JqrAuADrCnndR
2JpufbwwKJua5rSuEdaYqGDKd2Ma3tWtJz4M+w0OLllhiy7jcKMSIalIUQVJidTTrZTAeQzJTiN1
JXq/HbfscRS9N+xmQ2sHBBQnVlUJp7VobvEFToNP4S57wI47I69QYL3eo2RGfBJMJJrbTHVnaRm6
DfHjzHSicrvaO8yuio+ZcXOOs4Mb/+tCMooQs4JI1eu6R3jRez+NJZLuLGo+ikctpyjnE8X3FZW9
QdfytdJpkjTgXejF7P25O1HgDvuP2Bz3WDpNcKlHUv/LHfjbOR0+9moT+ZlMh75xuYbAiDs4zOQL
78R+qgL/HPL+8BQ+Y8uQ/qYb205Ka7lHgbdfe/enp5pGM+kyDdo3fRL0MKiuFQTKZohJjMtUm0BM
Rmunw4LODAIeop9Wn9Tg3S9knCB5YJVB+CF6f9QKhACeB9TvAuhUiftYQ2rn/B3v118rSDK75spu
DJ0Y7Q+38u7HG5CxIvdm0fdyOBEUT6QvjpQJkCnTyHmh06JZ9JSEEIpJO2TVROG+Gi5pxspKpsmO
hR/to//+9wpjJZZzzRtjLAkItN7RROr+uc7q5OxgPFsWpx40/pwFubZAgDj9hD6lQypTuqNHBsWR
eBb8Mya8CZllngc46YTCt0BIW5coP826hGQcSprlJeXgv8kkoTknQaRtrs05czoVdvd7xmYwt0lb
MDT7W4rIPcLXG2aYvwa/Qu48QMGbuvAusQNTAAWAXBKtQc74IxbKkHr1HaG75eU31JCua7yAHLcc
1i9IbIatnmJCTquol93+KWmyZJZTvBI6NwSVr1BgBlPC9Jeumfyx6pRwYZ/LD4G7KBxAtd/MxRIx
/fX1GOp9T2rooCw9Y4dFoHNLzczj6iy57MEwPiUI1b3akMtDb4x2GQzTmEKaR0lxilki1JndEnV+
/AuW61bjHJbtLbBhHAQBcwyIaL4Mzcuy1LXRJiRgI7SthC9860KKtmzy5iNFXKf+xSmNJFw4Z2VW
fLLmyPtYUrF1TVg6f3QxWSaoKzDFTx8p+LS/4zn0vBjyy3BCnXv5mZnV5tjIVYCOEWdeWQH5WpRN
pMcKoPnImGbfTuZWAn6sx/1JONB8ijiMJtGG72hE0lDlQIMemntM7iYGaj/Nn2xseJ51n4yoPVO/
oTDzhI+xaglj62y2UhH0TYvvAAa3qXTndM1vJGyE8z4ibzLPRNPpolKBgSKiXwF25HkaY2MF6NBk
XL3XwFe9D8t1sL+xV1HclZYMy360ADE7tFcsWqc8WfXL4OSP/GVG7EfSCfDKdnTG1r8/CORRKLTu
pZ5TT1REL55zclTa0Cj2h21MGW93aczxPqrRDYrc8xlqGItbuaI8y9ZyO362Mqy/FMlgtTs+uzx9
G2zxtGTMg1+KQsC89+K9UnU=
`protect end_protected
