-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
X8uiQIhCX5gY4mtw+i/+WwjK4Tvmc1/6N9TWdY+F5uEKTo2qzPbtp/hMbmAhZcTh
Oi7OSSXVEOL2g2H8FFFLf9eQBoiSVabBBw5gwPteQSmvp5lNMR1E5XpMlfSGwUBE
0ZnXyAnDAJD38JJKM43PcYxPcVpz9THdqNkn6SCtlkQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 121968)
`protect data_block
VPlrUIuwmZGY2Cgx0WOcUXxS2414SPw2o8vE+EfwI+/JhO8Kdfv1zAnizOg671hC
qLmgD5qgGKTT+nTw6enYQUxmY7+HGRV6M8OlOIzUuwooZuw1ZmjfumPb+OfCxSVz
msa6jhIWlkuG9JCRLvpIDUy6DLItk5793lR/gf6YehG24FIN+dPHPIWzfGlavmpb
HTlvPn0BZODc/5fhxCMxj+LqY5ks9SsU/z7yvh5u9W3MBG+GD70wHDdYtqm25Zkf
eKxaYYr/UrEV6nHPxQnuT/z3356IAuIl71mZ5ZaJxr0tBEyVnLPSi4hhCIIyV95M
fI8E9OGW3JopGdnrW30KHIgzWMHdMdncgQSBx/RYmanjT5QnEhkQE5gYrOcylCw9
vdy0sbc1HA9L69fPzq+5U93lehCzMyfzOHXGBxXxG+YJP2qXHTQCP4PkvRZ23fp+
lLLCbrj5xxBODPph+SRU07oHA2D1VWZWm0EOEZEw5lH//KU7c5wbw+pOFcvSpZwM
H0/4o6lcFtDiJAhUGe4P6hoTs9JjQKMP35HpE3Muc5gmFVq5hSPXLVbzDkg9I/K0
nAua/1J/+nkxUvXc3e+AgSeNisl1aQrKocjqNwmk8oz/jemF+PFv93gdQbBqXl6a
uHOKaXe+SPVHDyZCxTVk7LEoHAB6HWVaOxcZbiUL8k1LAIQ193saCbp6KltRJwSS
qabMzRW7BFIWSfT3waOb1GlalKQjFUla0T/ydFpzWeNbs/9SLUi01dWztf1iaB7z
Hv9bmC0A8sEahHd5Z3/sBUGxG+efhLBfc/qjlpxKUjdvanxoRD0apnFCh56e2Sm4
BwSO58/MZr7yYTPIbNusEi/5nHFKnoZQr0TtH79ySXcvLfl+hn/mAuE/jrzfj/Wa
SEucs7WLWOQ+SMsR32Iv38sXf4tlF2C33pKKIgqziD3/OAbmIN9x3S2NQxkM28iL
FleJp3fX9vqeUOMx58ZUGUSl0SdpPyNN7Ps5FJ73V6kz/7DnfMoFbrBv/SLheUyQ
o8047UjbvRMKQOeDkvKCL1uwQdxb83kOlE9BqLZg8kdjzSIHcEIEXKGdcZHDvRqm
Fb9qZZpNMEYveLxC+Fp5Dn6lGV0Ll8fixD0lsRcNdmdIESn82nYq9vN6iINvmjdq
lIyZ2wadDdE7rsFkuvu4pTKx2jkaL8IUOq3BF6UbFjIhrOGBGH+8bv91SCswi0+e
WKKkdhyMmfWjC3L2+BFVJxIc4oRJY4xFp2ijGATVcM5Q2QJ4HlrtV4oYPNl7kgIy
fWET4oUxygflwedbBATV+7WBVRVQ94wL0gB+64sxRszJyoF8JpTboJBsmCfomM2b
Ky9rCTPboNrTZhPFADL0sW+i3gC/zTJYyKFLCwELnTtoh6B1fUns9bGasMyTS7NI
5Fmp8YyUU41QLPCQZ35KeU0obcJ16sC6DArxhdQyxFj29B+B98u2YAieXg9mz0jI
9xv/MMRve22hNJujN1syyflWuFlLrn2ORlPbzZkBok9ADfxgc1MMn1CM1c0u1iRB
SYJi4KFE9XiVsmUjWpOYCdeNhpwZYROX7KAzM82J6I/FwJayEmYWtStM8o1kwKK8
f3o3okc554KkThXdiY496oCSuhIfjmU7R825tcmqNl7BYIklaD/Yfmw23RqoOnc5
8c8ArRaAX3RZ6qoI5YJ6Qa6zEJc/VUVqmobtZGquFSyf5F1NlQEbVeKXz1h/Clbh
07D0Sgz6vP3rSHRTIlnKdQ/fZ8tVs4Sxt5u9Y4rZT4Nxx79duKUE8q4/m1ZOh/rb
M+J+9GULpwLh7upTiaEXWm08KYh148uvZxcTmI9ZPpJ7ouXMRu+tju/gleF7dv5r
HxIZkZQtHuxIDipqOucgJKfLXVIHscKczYyuHFbMiy0kEboDT9hjRl4NSEckVJ0r
sdTI7dqo+V8Bn7+HOA+7fRSyOt9NQM5B1G8UEic911I3iPu+F+RiaC3PV2wC8K8i
voXqtlxJgb8lbXKl0M7x+d1GBPfv0+jLBqjXjhk0Vr78ZIJ/pACsDkzTe0KEQbaH
cY3/bdrn5qduHTJnFateGRoGxm7CKfPhZkRt892+6XV6ez+UL34LIJaeG+3VT9hu
P5TOcv6v1urR9svYBgKGVyhbTji7ZkufhTyi3+EdXr9F4NCF3zzlYw8wK8qLZ4QX
pvkAXqfCmlbaPZFxfPtJohwdCyHW2sK+022ggSQgwJ6VNNgq7pDOK+hyYZRo2W9i
mWsnGkhPaJn01bvmcIEzd21Fo7OHwX8tn1EzEoXh4K/4K1hDSlGNodyzIgxg92WS
ieJKWLh/DFiq+sUgmmpGFfVGKpKDMlwsvgcHadew/2cCAzm8fEQKUv+UMGHqjTsa
I+QfKQRThaFS54k1n85W47hTc1C9xHS3NmFI1eXe0M8a3MYbJkJXV4CIcQudbo/K
z1a5k51HOrftM+BtSHnZb24UjgZMJfJORCUm6q5F7zrjBjNVqqcb6C5upI4DPH/0
ujEJGCNEBUz5uUeggOzG10qwc7Oh5JE6oNZ5x3SCw2tDkNWCm66zPI/um1aI8rP8
clHQ6F5E11ApnNaP+jtsKP7VLxBON/rvhrEkj+SMvHOQkGJq+TWz1FyRSkRTH5D+
HzXKfAbWhVNbWVaVVaokloxo3yEMKE+0K81rQfSNwTSiGlvg0gUGZurtFQugZYHz
Z1plDTedivaQcqWqWSHP6yhCGdkOorxEFjLyeGINSKpevuuZDSZMxGOOfEjtf3P9
xMOqr6umU0+uA3sXzKa4rb+5GY/HGVCi6PQAKvtijKpGTbWVT7tNRt89sQDdfVS3
k/SoYY6BM7gB01mlp6kezYXGozmIWYV0lDfSL4KMUFLSvOGdiBLFtnJFconMds8Q
onk+FBkiQU8pXpvHgpXY6SWszv6PSv9N6s0GrlBiEbh7tVJe7CsiedHLRhvd0AjR
t4cMtPtyKTqL/jKY8QFb4YQTSQMdTm2xkrQHhlh/HOwBpmRytfO5mb8vH/S49zch
Mk/PVHhk4GQc9BTBE1rctC08/7GlQTcCknOIgpWruALWImmBVFuyXHxB22lEeUjc
LRu9DyWIPjImEFGQl30w7qgtyoe4JTSnv/aRzPQXLs1NhFEE5G/yr+80RpxnJ9xs
UTB8M9SrsUVnjbb8m3vSpNr3aMcwv13Cxvt6iT89ZsDG8nv93PhVb+p5bSZV5kex
yz5EYTAi13FAl8TU1ryOvaa9+zU3aOo5zZCOolvuOK8mAkoyPCtViFJJcRXcxwtI
BpW6Sx3WeqTaXhP2j61SpRxk++d3wwIflvggxq6Sdtf3iZ8wPES7f6F5VzP8MlRG
2oMi0U1pCXg60pvT4V0hrzyrXzGqHOd+V628hS3AZwdAbUhmnLTK/Nn4bXQ5AvOy
y1l8wnHV8ipP+tcadDVnNDaC2Q2rt08CsXxsSYDfM/SICd/9OG1XgSj+V8eUSlLj
Ct29x2DpOXeu8VnxxcYgQPrMmZ03TG/rRmcVYFuFpDyXq68v+artepPaFy1fU59r
P3YJNCgj50Vak+zBuX2h/GhkjhYNX19uyiaoqOoKKd5lRzaHNnPf+FUwmSjegiL7
/C68kYSO5PDmgXrzXeyMf3PpHb6TzeNrKFddU4FBsRQJNvVQqefXkfSMEOjSA9cp
Tv2bPA+86pNxtSgBcAQ3QGRWYRMeJmhwczv5Ockfwt8P9ZCAOajEOy6W61khsu/c
Y4rn/bpVvaFAlouVd+UBGY76sdYA8mgA4qi7ms+YuJ7uDkPRVnI86eJCL3JERMmh
aoZQeDkn/m4X2NTxP4Jx/3oy2BBPO8QKN+Su9BMBtskMkdUusj5UjZq9X84aC8b6
ztiUk6hXMbBa3Aysk1TuoJYE7Hc5AoTUH8KK9WOgul+EOXZxd+Qfr8JtrAdGIQgL
ZgyWEjwnanb2gS/I/NlGErzLaHFabINKXaPArFNQ+HwIPqVvJeJIRHnl3nz4jWfx
+qdaoR/fhJcL4NWQoLBV8/vCdbQO0EXjnEwkWCcDT0g4/9TjdEyR5GZ75dHgx0+c
TXL8/uVZVvHbzMDQ/2Xrx6GGGFby/3BVencoxFz5yS+JCWPBKkB7Zcw97cCS7WE3
hIEZiigoc/HN1lT7b8hoCjiL1IPnCReZmfR6H5Esk7F1sAQxbmXVzjFLmc4iJTiV
KfIeaULhH+vlPwX3WHzHArbph9h/mHVogxd4dUVIcDCFyHMQ91zzjqWY4u0xnT55
9HsNfAv5Oe3rdVp8b6NF4pbXrUQ+L91t+xdk6pmFofyw3Wuzg0to8IqpOm/i2EaQ
MiacfwPWb8qRfOuvfWJeOSEvbawH56qWn7W2dBVkDqMpQ0XQWPGS+N4XOq+JMmnY
j5SpKQKyeB22vE03JiJefcPjKMgLnje9T+HFP/YC5Rp4V4d8oeg5q3YwCSx8oz9t
OXzlnS9KF7Z6sqJ6e5qNdgIro5tbBy0LX463eW9fzXrmQcwRcLITOMf4AiPeId1g
tJGu6X82NsJA/2k1xbAlUlP2Fd7CSB/XdkGIK6gZvm87rW7z6V/6IwGmLJUrgIk3
EN2IfTpx9j/UWbqjyi5SpgUZfM6l9zJcnNOJG1qX9pjqYyGEgpvlhAKmjf3oTmxQ
m19lpdCp6KHIsc2zv/IVyVJcfTyzO7itU5Ysv/GH8M/VeeM+wNpN4ZdfuZ7FsNLe
a8dmkb5Z4Z04TPo4NACCc6RQNKURyHeVvNj8EeVlCS1HgDXzZlpYSB2g2xj0zVt4
mqu+j07HJ8YZV7LUZIHkgTKJFsdLnUfyCFFnEjBcxOBh6JyBmFvJ28Re0FiZ/K2L
Y1TmyQl0HYrIJm2oRnzv14BEX52a32NE7Qh+8cuCeu3jyxcgJp9x8Ag/JebdiKMT
xzyub1h7PexsmUtgm+6/LRVAFoV2fse4Ooaa+YVLnVgDwA6U1X7l9WKjy2Me7Tcm
aoan+do9vnLqnhd9N24Z5ttIyPYD2aFpdMcpEy7yZuoBG+awLXE25d2D2WnDyJ5W
TM4ftVAkBBuY2TKS/YrZbjjekBLP8oM0mC4WlFSkAGh98p0T73lnNKiezagCYnNA
w7NjFSQ1RssVmYh3svTC08+PwNmcnXGR99FmfR6KEtl985i+jl+lUfIkZYgwKfB3
MHFn8clYcdvS/gSYyhlTvukDAhjCYanz87QYoYozEX0ccjIlK8vP9dS9ht6wCALa
kmbNy3/LqHyQhAkZ4/Vy6sqS+XWhCZlz91ufQl4k67HG2bmOn2G97SO2FZU0TNSq
Uh406Xink5Jp575Vi2znl4uvwIzVrvltVfIOMj1u2q1EMEspQ3cNpgBQRze1+neS
JrLfyG14YWIuVPOcwvXDagUXnu4vHh+n0ggGfRO8eIOzUhjb7W0oQZLVLu372P2I
whblHlagSsJPKUxcJ9RF/hEjtJGXNc5wvfbs2r9vZpFlscd7hqmy/wOKnPTtYgpX
7odBUcQpvsoZk0fKXBYbP4NreJoWFRwLEQjStUXPceMR0j7JLxViXSQokd4OVI/Q
xyv1vLYHDS1vrl22CA2uzNFTEZ90DgHVc6MnpQArPugiOGPigNKN2teYl1gnjMbf
Si04bxUANNNKzTtjxhe4jZKIQGSv6jnPvjPCykX96XK7ErvPS6qIx1K1wHVdVdQ3
1AEasp7DE+IC7epicknjHi1LKW1+Oowl4gAYA15L12jIRjhexLtEmqiokTLWJgwl
a4gn6T78A+3JWCSEALbDLh1MRwfaXJpgvxKJUYASagXUKVwTad2Z+adYCnbYGHAP
+WjOdV/Oau5BzcyTUNM4DKYB1Vj6IZsVziQpBS7kaH5nRqw4zDcpaGiNnHpK/w7x
/vzBiiyHZjlu9xt/IV8Holbmrp2aa9SG5hnlGTLeMkrvp6j6pBjbN541u4au+egI
DQ008cqa4R8urdABHzT/44x7QXcsAMv5HwAWlB5NrpFJkTzBg3zNq4PR+nochXfZ
H4J4aw6fgMaEHrz4BRD9sl5K4i86v6B7TW0lUUwJ6n6lNs/FoKcK1E9Jt1UOEr5U
tUxrnf6jdsVD2tQUWjFQ2u/eyIZw/eFah+n68Q/g+4DCBbRVxs0aJWazZWtmozpW
3Rg29eR6baRzJHPD4aRf24mBJgtcizs1YobGLiskShuvVlgFaENETVUMftV2fhpt
mc7nc1siAJMRjbzMVYZbT8Ag/zDnuuHYJq1UcM78kqeWFAOx4qcBe51TAo/yQPgF
VLQ5H6VuNJ9ImhNYkng6gwz6+0i1vrK/TTJMRWpDG2/pbuWkmyE9J57AmxMdD30T
N3NVvaw+MUBtn/0qGS0Pn275BOWjQqfXiEKFpnZsB0VQ/+4xjdyTaHZOk+No7YGI
7enTCUno8SgjeUDrkZhaoIINXEr/KNbZ+a6hGaZqNWkNb7+pMlLeGbJssI2Zcz+M
QvP4xPXeyekvYKLNypMMuzMSlYRMUvkNqSbecMmALz1OZOcCWJ/kheDpHiZCELGZ
lfZu643p/OKAjgRr0GzVd5DbRw6iIuGQkenHB1PIDOBreIMhLf0iujxc3jFiCspL
+FJrK8L15TE5Sm3HHk5s8neXjtGzz520vt+5U2ilpiGNCwXplBfAevKoGj8ph8Ga
i3Xoelp30bPNQtf4uB9mLdQYIC7SBzVa0Fj+cdLCLVpMSKI9pRBOs5PxD5/iAtnu
pi39igni2Fwbw5Rruw+oFUyneztm+8EZFoFivrQvqJCTYmKUiQQOW34omOY7Se9W
6aFlSp0lC+wnBiD7hWt5UoU25wluegHO4HqBbqjrzo6IpOEjEjrUsE//Y12iyXLu
IkdOmtGPgu++gBsWVWjwG8GWBIKXGe4te0iNCO5VhHjoFiUt9uAlUxQiC+RaiHiD
B5xjARsKd9wvajP/Z4CDZP7Vym7MtNPnjWNEae/pZ4lzAcVdIEE3oJNfs573qTht
UTrJSxDyR3H2IGduNTwhL6jI7eUVMaH4zIwqK3OJ0ku6w96KQqIKeVm7KHpPgyY8
trOJT0UU3BYc3L/inEF888LkStdKpoQMHO7493RxoE+iQYcU7UK3cgBMAkUDnlEp
NIUw+xW34vyCcLqZGpDTEAdOAKA/45qze/tuOoVk91Tb5N2Zefk+IhnK6EHVyfZs
ryi/UhROeUW8+mpdqmr2ARlTL2XAHL1TTb6qOyOxS82Sw0wml59I1UJD1IMjHoWN
WHfLhLPCcHj6+IGIJ0gQ7s2cMmw0R5/f85wpxHZdsbEGWnSHnPkrVvK3zVbE4xAG
vN0lRTkaoK7o9gWqgTAIDc3tKJVZioisgRn3ppj9eHWLYPdSrGzyf+K0aWQthp7y
SYnTlp4rylMZsbbmnE59nW/EXFe8+4RVWx9T3ZrujYfeDWOYg7kZGmmAf7YO7uNA
nzayVvoXNKsPEY0xrQpZn3QzjqVdfasBCWempG8vUXWLZKb57iyQC1tzBpqGL+Xz
w1KptWGhnOUSNCYvi5Nt5gy/T8idTjGuoUKDJpxyPIvh24+UdQVTUk3cjYlyVEbY
a8jFteigvx0AVCuMYowdgUT8b0x0pOxDElGujYX14/ufFYIR85uvBHA+cKThcS8g
bS4j+JbFo9n+I/kL1KB2aV9elIbeU4+BoYtbJBn+VCL7FkvVkXA1rWzILmLi6o1Z
q+JCG/8bdDd4nZkjkDbhoFfBA3pCPn3/h1mv1RvagDQTakjtXc1b3y7ZspiKhP/T
SIf0/3odO7aaikjcQIZCuVW3WhmRPS7634Aul09fhBi2atYBi+2+GNeI2KHAU4gZ
tjrzPgxX9EVmd2bWnX5LPt3w3n1L+RIlObBP7hWGEZm7glMdLYhegNYeMAKqusHm
+mSxL+VdJbquBl9LG7Fq5vLckdik9PvL1Y/1ZTA1ziRf7Z+3jiNgn0SmlJL9kWSQ
X2auvEHvJDCvYNdhE2ebdw+cXnBF4mtfjlum9wKLUeXnDJjtzvar4/JhhLr7gdAY
5C3KBV6oxJqBPKO8X3qP0ABtNnQGtKvpHViXqhlP0SMw+FMv6ggduMXyiyS9CFJi
vheEGDaCl26GuBewcuezHPzjl0EzfX38HHM8L9OYpNwWlm2G9nDrQgGA32MwyeFl
Enqyoffl/yu2uzIW8rBDdofMAYhZvbIMlbbyjO1MGmVPjcQl766mU49mWpHumIfg
cR3tik4AaK6qe2SwxOfx8mHZZrIEX2SrB9EivpKdDm6Cnz2kCGXCq9Q8dWcDrG0Y
wwG2uU8kLDbaxxqt3C4Knzx0FZ2PzBtMeMtRLuhltzPEiYuNUUTqV4o1fUb7vi39
t/cQbuOMr5SpimqoxH07YycV1NtsSO0SEO2cJgV0I+Zc2GRNej59TbEzq2a7CYPa
Ytr/FRGGNriAGq6VVnmAKRT6I8qeOgXVj6WkOePnZ/G3e4cgapooa7IxypV++Dul
38kyzSPhU7s8jNu5cNryC1HirzG33+al0QIHa3lNGTbA2BtG1bvAs64S01fVHgWG
Wcae1UXtG2zgunDxBNLYnkWD+HtYTT4AeQxZv7HSTlbnKvWA4NNXiVwObpyBSV6a
8OGaqAIWBtbmmNUpoz/Z365MzbOSKvG5oQLBxLdU8/SVwGEzceFeL2syJhsPgRaP
JNevmyIzTaYDS/oZO2H2gsxMSCZ0bjs2H2BLvPHMbFbxFhCD9vsvSW133lM96kCv
1SAmBGmeNTxCUNo3UghHkp82zwopPLjdnF7dYGUNhqQ2IT5q/H87F1xqVOxz7e7u
MvYcEIF28lWpK0+YKg5zGwzyj2KOZYXwkc8xNUI5i0chgssWBrilZJhk/z96t+nH
ILdTfDNtIbt2B77ShN+fA/qzmqwYNCZ0xgnEctC8rU5Fi8QhfvT99qnGFBM6hhim
apjteMZGLwi7Xrkpl5rOHdAU0W34XJ/ZNsZjwNtwaZOuW4xnkyir4rQYc0kSlQdk
j4bXgABlCRbHkdat0dOVS/MI5b5VvzZyTHWyu0d6vyhrJSjjzI91wcxxJssEa4fu
XpYDbn+UTcRYtpa3I90GMG85fF9Cjq/yCIVg2O55GziEPgBW8GgIeJaHiw1b0+xU
yaVuQ3l6DFbDEZNuVNQqDGg1BAOEPTKrsNXKMOnjRPaBlD1tqocUGdTlBPMG3dVC
0NEh4rRfNGKDXVidVGaE+UvKFyx2y0Xhj/J2ykAzGPBt3eUIpGisMEKA+adx2lz1
rDUxoNlYov4s7DJvDuDWUcOv4sr3EjWkosbB/RhrLO1qSDQwxCbgrLu8ahPokY2W
tfJa+EWVuNz4Zf5Vr+s1+dgg/8VvPXg6UVpP9F6uBGIQAVdiP4W2QXiSCXnB9fYN
P8K+WNWToJHo/E2FKj+W70sXpm5LEz6vMJzJ/K7iJxtlSnQgUX1r67lbn0Dy35gs
rvcM8/DO+I3uLuL5TvdEsj6iOOlhhFkLLTvufZY2maGLPXTOm6C7VEsVKOxotXF7
S3KSILOSxHDGodgu+H2fL6ZK6/zj76LHqb8hSzWi6ZmJkl87pheZyVwWZUQGqWEx
Jvu27SelCU+Ly+6Ryr7WP1fFEFtUIonEDKrXZwz3xKwESSoa/cX8chlnQNR12keh
RdK2R4h/tQxD5Mh+e+vTSSWyUFnsVnKtMNuyozkyjERNjizIY3qrXH9DiPYRZ6AV
crdZTfogzeP6ctuYi3UnPGu3Wn3P94zXJ+CyFRYq4DJI2Ju8WB9xNj+mgcFeW21Z
WzUdYwtkp/fEiZCS9Z/txnczPuL6ICi59B2tjPZqFRjb4sHJIYiaQYnrdq37cmq6
hd1RL+jZTKscEtDcbkpcsTbT498ypIpbM7krnXiNLclSKTMk8reYgtV/INxElX9a
v+cEGVbSgRGLvX88iY82ShqWVI9XpcYj61krx/bs+x48Flx9+h8F6FQMbB0V4hTI
cPAFPubGul0hOSEA1wzdXVirAp6jdqLgRFDKGPO/QbcPLqqZVridcDSanI2L0ADd
ScIX4pBA6GpXP2tBYsLltiWh+t4TGRFbiLfLfgs7MiE2o9ICWwT0Xs80znIKloda
jyHl1q0HjSclS0BHxMqTLFGm+2AquLLdxiV7TYML73Q5fzM8O6J/qCgSz13sY6Zg
hAi49C42Z3Y7a7hZnEpqc1AXnDMgAWbtNRzlfDhiUgX2wv7mCnMpAdsiOqGZr1OC
V11T87tKw83J7CSX/bM1RjIhstvB60/U8KPS0+TTFxcJH+u4D1/+ygyKtdZvPa2W
d78X2hGA6WLWF209MMFepLoassBpx++habk18AYAlM+RtEEq6Jlrouyb79ZOdwYT
Zti9jYSDVni0BLn/0SEsIP/PHyclsdXb4gP1bY4X0KZ0IsqteUS9Eu/4wrYNUuD+
Msk0RfXRlzEmEu7Fuh7JfabjeBSVzUMfgyeywYgdvxNdY8+F/QwrHvEGTydjw7l5
9uXTWS0AEfUpJVY2+st/GSMPycXF/x9rQL8RXCfCma6MhIPCWGZp3k+BJb3iLxT+
ETf3IZ0JaR0WsqIHP48m9ooVvBUxYWTJei2vjxlsqXGyiTFebn7EnwmEMTfZANph
A/zhKJWdXwLCyQUg94MscPgJiYIoesVGS6BhYOixRvb4Yf7g+K4b9i/vnHzDkfYl
bbhKKIJI9GVSR/B0sQUpgvWwbZMEdDWu8SiKJfmZV0cFiM4oHMwYkryHenvq/NQS
6aVxZiJ9dryB+uk1qzvsyXIY85QGWLJVIeGBSQGdMGkV9ZbzBKict1RcDQERIdI/
/sGIzuKIi3zv+WQi0Y0uON1xiZDNMADxzYPtZ4b0P0CYRO3FxIQp80XwfBg3JWZC
rpOEsQWbvFvYWTf05gIAr6eWpu5RXAYdCXpV6UIu41CPsjRAZAfDYu78OAoEK4YQ
hbNfmmsS55cR0jykzDP+F+HjGeTF2mKIbuDlCKw73FHdhORy+/XuXCVl2UZ0576z
yH/tNocqI0adaFjPUIXfpmnCY7i9tmeMQx9K5uCVXwasXbQW1hPVYwbg83AoYplD
kTOGMYvKaMuacMVBT2VHNbocY7SINMwBfXWQ4MXRqAJk8b+LIa463mOnYd+sPA6m
vcqmsBUwNfJKNwNWx9UdoFx+xh315g0OVwRbjJkDRnv9m/RLRTUKrnf2ZCDhrAxW
b1g2j4LhWJ+2iUMa8uS1foiOF1ZFbvc9TZ9uEEJLj82gPxCZE0uLy/eJoMdgbJut
GO5iYd47q523obqmydNeVybu1bEktR/zIrSJ2eK5h3B92SWTGM+7AP6ZCrc01ZO+
7PTcAIjA8xOy4Sr/lCY24DhN0DVkkSFauTuXxbFMOr/0tqSKAlEOWrC99Mwka2Q5
ykPUWyEZGAJMA6Ev5JaYjZOQm1NrTjO2vCb4unXL4UteWBW7yO2d9G8F8dX7KEQU
FfHVYdrP3ARyKj9BoQitxxEzqcSYMyvmTFyyFDkZNFUu52rqCyJTv+n+s2DYrOep
aXnNucBL1uVMbhgX9imhGwIMSEutXAkGroJDVxv1fAkhndURMIgIQdB2jyKXD5+x
7QynWTfOsdDL39rIJE2NDKghvF4DMNwqWqfwuatFlQhGvlL/qDykVteL3MUYTKLB
BjPIc+Tbqh1yQ0vXFQkXgQkuswi+HVZaDZCdTuyWOWvKJNh53RqOw3YcunkGkp3H
qV4Z0LOh+cGglCCEIs57bJMSKDGEoiD8Z+PrSuqGm6+SfMDbqJmGJz7HkTWLFnWi
znzTZXwCT6cPS1ri/ocbDJ2yq9WImR0u0k6Yy6ZdXUUK1AaJUyAyQoMeD/NzI5Jn
Bp4xqdtpvwa+BaXEMGgKjFAao+Rccyi7HH4CB5tBCGezH3cP1czPnuqTFe0x8/+j
+ZbsMZqX9bN33af2oQ/z08jsqxXAEmAlkO4kuwifPxfPPII2HldYoVsMUfhXtXVh
09ClEedHdOF4ddXAdRRD2rDLKkKKOj6fYJBZOifxlrZM/X5UCAhQTWkCSJs6JUl1
dxBv2Ns+UMXugvVz9fz/sdXY3uyAqUhV7vI/lcmqjoHGiJ9DvLA81hMKfOTve0B/
6HfSfoy1C8GBlRpVpi0yvRo75doSqoB3OQ0qbkE5bWGMhKwN3vXB+V9OUyoxmARU
6QKwLRTDHA//utvdwSCeXTtT6UklSvCQllX6bx2xTRagdlbYl58wh3KFUczEv2q2
RF930LJK6GNUb/M7kr59Ek0+YgX0vRVq0nLjJDXZMJEansdsTrMT/p94J3OIEMU7
+jYsDPClB6urbNZDR7VUYdsrC7pQedGU2/+uhPhd73tAldTfV9mC8s0qrO4utt9G
BIprzSaG6F5DzDNNEHQ3hlA3VWsN1ifNZ/O6Dkze1c/dxsu/R+Dvyd1I2q0Db2fv
cQHXw8gP+WtFqqFEpcszoccPntnWRk8YGsEdMeADFdaxkvV0Gs5r3pJCwV6RxFCQ
QrF3aRE9FM93yDTP398fAV3vVi9yFMjvsTpFp+VJzejBGaHsppPf1O6JNTORVIE7
BxkM8XZf9R4iZPpsa/Et0EyhJYbxWsd93JL3rrw7ZRjFSwxM9xXsElZ4EA0SMsdP
ly60U7Pv0NIHxzHdOQUASATeMFQUlvPDUXcjHrT9FW5l9ZJjMEUfHjG6BHYPMr4W
aM6GGZ8I9cHbymwosiawDgZ7oCXoqh9uobsOSHogDmoLAzkR3KYwQ/f+BYp6PkHB
zUnIxpEFkzJdTiwVYQdvhVRxd0GQ3v7j0+uffMSA220hSpdJbzoIqlBIbEoDaMOk
4APkxh64byHt07lE9adegyvesaZWaR/xNv2gvMB6a8YmMzyaR0l/1E2GVmyHgJuH
0FqF7c5RxznLkqXveRtGRpMNuNI2ogjoJyPGPJwpJeM/0DlUNebgPiwInx65faii
Ia9rjh9vWc30nRHN5ugCbG6gJBlbYiEXpVobikGO8ZmJR7kwtqxy+s1UXkZqZBbw
i0APCTQiIP9fMKx/2NY5b/J77wLTl7TlgvPE2PJK1znsguFevi+yrN0Nrbo1Zz5Q
f+HuDZ3wpfI5eqo4cR4RwAeK7pCDQ4R45alPlnmS1f2tY4/vzJBpb1eBIwdLsn7j
VPEfo8EqXWoE8bLo02CpB4xWyn+yH70P49c15RUb4c0Bq+y2DsbU1AGrKI37KdQa
zHlrbbjXR6YhgD7lvkM9+W6suHf5zSO3oz2iuBwhznc+ztlq3/Gkvf4ApE+p5UeB
GkuSw2qjz1gr5/aTgFiXmqbLS8gfWuBDPUf7vtMGxad8A6l/EXm9EQDavFrcv7kl
kzzr/BqBkrUorZwdsWffEDwl5Uva5SnhxqYGz07lfHMUNQi1qYvMrmFWHtMDV7rx
N7jW/QRByQQKkuihwetOlQUggkhQHOILv3/yqkG3QFVvbLJXWzFfz4VMVRCOrrn8
9uXIcMkwJjwR+1C5RzzCuL0Q4tNsvRGD6hOGAJHGLL4i0oqsgnOtWZuK9TEIrRx0
BYXUpfBcrk5f50F0BFE9osdwMpX8Py3J8cAmuUDmHmxFT/Z2XFCswHIe/IYUXQE4
qe12l9x+7Nqg27Lc+2t9jABZWIW9PAz/eehaIALwoP0ypT0xmFktf0ppII298FLl
j1snFNB6qOWcBg5Mqta+F0ZjVYMmJIMNbEmXCTZoF7giqj+0YhA+hYUn+dCSMY/a
XLMKO151vArZLcs/OJawidAKkWMWzMWZncCYrCoE14wjeP+/fX143jjXdlyXyvv7
PqqaCbTVdlF06oUhisCbb4AF3vjTgxvP9eoM6KaoclQ6Oo06hm2P4hLQl5Awx3zF
AGrG71hr6qYnDRjkPlZbHWqMaE4f9RNmJ/KvjtkaofjAGhsp9zgVnGK0qRS4YNgx
k/GhVt2GwCte8kwKWEIvxpXIpE04Vx1rVa//wvFUmerFyDkPDADMW5Q0kor+XNgn
TM3QaOikRc1C+/7HJZsH8D6+V2UXcYGsA7Oo5OfiEF2Zsd5vSiwXBIIKRnzZOLE8
/3r4Z75b+3dYus9ExbmZ7Fz97mvMI5/NX0L8CZqEHUqGZZ2j9o0civiwq0Mkd4d6
dXvVXP+w8Yo2YoikPwhxrIzDfVCD7QA+HTgQj2XlXsIn8lDYhmdB6UR4l0kk5xPp
kZI7+ZnrM+Pu/jfN2XK2BIZ1Hd3WCV2ZaqLWKRLJj1deeC6bXXw5jPsZLqL6tWoQ
SWSzdvG1Gm4kKf9d2PZK4ty3GyIvaldhvTlMSTE7R8GtBTUJnMaLhYmDubhNj0+A
OthKSC7mDn8qox0AzrGZTbvYxgPiyPNTBUy0SPDHYHeAR1RkCT9RnuF7FhpC4H3t
e57M0vNUBsAX50m+5cumeqaDogxPJJemb62N3/yANzIL9WJZNwPEhwabUXZvtRM5
TzHmmExK8wmvyDzGF3elcrCYLki6CV2RnlbBc8XcGrA8nozhPWf1Kg9omGsdttwt
hlwuvuOS3LX0MRsLasor5psa1ZSVaTageMyhvnJBGcjzjZrk6ETHp06BJEBxANxY
1F1vNUwOL53om5iSAOL4EszLdtEfGjpF1wcLfRYvSVs1lKEShBuMdSQa6idARv/t
zyxOF1gioHJV87yWudT9QnZ19qyavyeddXIQ/Ny17vYMHCCQIQXPomN4WXwbu48Q
oB8Pmutfu6wyouGYzTy57rsmryRkW3Lx9BPa6442Pcqmfl6vsg4Irz+mJ15Gjeqs
LgQ1dUjMYrKV+IWQR6a+KzENsnWLDQabiveIpryOJWjsMJVJC4JZFajrOY8Vqc5h
hvWX9ZsNlK05V0swkdIWFxXqbBF5YbHqf1kfNQhDuR4aHmwKcyMG0M0z3KCXqhdi
5WPWSjv5cZqK1LwQQQnSLAxK7AtIjOaeeVccBnvssc8VxgZBfEeF3Riu6TzhXMtY
lfiUJ27QhWwF6nVVxyd8259EoDtEPt1CO7ZL8klrJeRaZlhnntScSVX5Eupkj/f5
4//7vo74/raTwilRB0/g6fPRBY3LUHjmmdtIY1D+r7a3NLX1+bp8WOl7QKMUACgH
hYZHx1ot8RDE1jYT3T5ir4ZFFdLIejilBEa9GPFI/Az7whV6My5WD9b+QlnY+9DT
hYBxMWA7pA7c06N4xz8boMSI1Un7FcOab4Lo795jBy9g6cH7opPufpZIE9E5kM8q
MW16gjF8GMKvoRKMl+hZEzRTGZCrVHx2x5RGOIg7UhlxIygUQQq+zCwKlhjj0+T1
D5t31kJvWPZdpG0ENSrB3B9VCJEkyXqS9a8LA6ckLz5shzp4SmzxZEFguFi2Bh4K
GUgZR0NgMaF48S7iDRaTvilyxxkMZMvEMwxbm2EsvcKktF3PikUbcuygSOeC/nUJ
XlcpfCMB/2iaYVF65PoAmTtraljYG/Gpf9HfO8iynLKC4fFBK6KqV3uuBmM16jFe
yXmC+17nVjvqzdQ0SE0rThqeV6LwCUqSjtseu0JIioJ/F8kiMxxY6nnDqINM1eh4
UvEpidAv6TZ3LnZuiei4Rb1icbzoqYhxqcl+CgHwj9yMzS/9D/3fGHG2DD/nXYZH
8EPd457wHTqNm+XIpj/bC2W6yE+lEJNkvv/5TfydJeM+1iMa5lm8ufHesE1F+ipJ
xP3JtNBv4TtQWVMGDSsyZTlkHEcKhBYUCdipmqEHnKgxaDXKvBBXacGwIqLtqnt/
iKFiMlr7jBnvuVlUqMR4M9NMTOTxxGjLnLAbKlBFjeicGA143oZEJ1QsXx+hHNPD
ESdHJ7/b0SImUaUcEbxqzNNkj/y6aQt/hgbcGhtj4Zgz1Rrqc4xw+gord25nlhqe
9bv5/veBLnblm6TPbooix5FO+vl1wJskjravERO7CUjRPdOTLaG9Dbu3tn62eB7x
u+Pb70KAYdTJQuG9xtlRQoqrbpccxVPOVbX6WhInAdAzqKvQfI+frs1sCaBlrAew
yqj6K3EmfSk2MID7QjNysDIpIqlsQztiuHO2O4JLiZhEIDtpMIjSDXfg/8tzdeb6
XalrBdJzyKKsemsVKOg7ztPXm4pNJ64jayfsTZGwt80GtlKynYEfwTYvgMxhpVQ4
GdOS9HN39EqLfVjdCXOP68JOEoooqNVze7exN3fcNKuVKhNrPhtI/lXZOKYxL33G
auoG+Rgn822vneVccj6th7erWVVPt3SVOcKNJS+2nb8D/Z5E1XwSnjf1yzhfDp8B
rUsv9ilgc6cJ5mj0KbO3ddJF1yxDcf7kfIoAJ9Il0pT3tilAVZMhRHVIxS+BMzFf
walIzExUvuE/Qktv72NMJahVfZcDUCAXG0hZV36/GCc8NwuER7NwdivkbN5iCehr
3f814SqZicSXXr327CTu9kK2hX9muts/GNa7n1/6fPPu1rdzPAAuiY/dD0dXFU2M
bNzka0UmYXoi4Iwke9MUT0GJ3JAQKFQanankMDYyWCvs7r/0r9t4em+OfE7fUJLL
XvKCPXPDLWSqxjf9e7D/rr+W4TjVbAkOG3YKDiuzxCH8j65rtOVxCQBWAcWSYJWL
wdm7/CIp64DNVwQmHxUmrOQLTEpGp0CC94qMzZSumXc0Wx20/xc/c0jQDgi9JZBI
PNS+tBqMsLL2ntLzII1UTkxEKKF/UHjJe/eXOL0FASUILu5otyiMu7r1qH20WG80
g3ESttCdKUAMO6hZvFJMDTgDuCXKFe7kn1LSiOH+OnZCM92UFE3UtwWVaAImbsP1
AZXd4HFJbyhAHmdwYTWmlN5K5AUxUV8DnxssbQ7YKIcCPcWG9FOOY1JU5X95qP1q
b72XlRe9BUaQ5rrESs+qsjvcDN4dsUTaxV1+VM52xfeBLynhjTSsfX/VjGIhhG0O
X+MASHqCyhJ4lK+QZf/fMXg3xKeTOrgeSrUrp/+4WcCafwitxH9T/bCdGY8RdsJO
cvanSmgvuqQ41hxTNe3eGbcVae+tDu03Ca2TFHnXAHsTiNH/CAiZNjnfxNXt+mql
N5RVhmZn7JDwpUwY9GVHiQ7XiNfDM7uLGIfzdhb1TXq/IKW3oFUDAoYD6cZX76wG
BVBpAG0wIHLvGHLDSMNn4mqSpNhV9aunsYu9gDBrJPnECRGLeiv0XC8s6a6ha9Me
9vIquxu69E1uJLZbrPWrxwIJfHQMyOYhHuaSEgqq2iJHAwBiyekaljAq9yxJEeJR
t/wujz0QMyeNYo0t7nf2c4h4dOcr9vZO24DGmBS1Xb43O7B39iGPl3Jblc+9QnNb
/HnwZtvP2lGT75Qz6Lc2TxWSOcIYvWRA1xfK0x3WA60UP6AOgTEvo/UZQfuQxuUf
OWbk/P7g30mg4LT8nwB7TATt3ipd6aQruhT0t2lA5N9Ybc14LmmIjWDaU9RTswLd
+x1nylNcjEPAW5yNp9ssnuY348dzr+lck84gwPnaun9IB8J2lfLkj0eNDyl0mAju
d3wEa0rQU3+hU+Cac29nXITUj2WzJGPUYdRmgvoBl2bc+M+BDAtyh367nsm6JDBV
crOHyLG6jRL2hVhjXzW5jABUn+5H4a4fEBDsolpvgbNMTof/XQciUot/ttDxefJ2
lUUOrL4QB049xuvnGYSAsBjn5d8DOVxSNmEvrjFUGJeKYOYHnSrbJg+b9cH4/g7R
riBRuBly7Wt7FtaeMvV/0xt8hMyQo9lzZo66K+olwqID595suEL2s6DxBIo/qR2/
asuh0Drf36AduwHlgouPYPTAbMIOy0oDaupsxK2WSFYZsKpAQXDDbjGsJvtG7saa
gdNnsZjJKCCRjpDj/G1tQOkUmRutGJrENs7XzfK6897HiQ/jkpG5GVT1M8sFrv/O
kv66Nd/SnJJD9DtbyTKA/+Kwape48G2LdFsRkhHym/KNXWdvXo8yNk8EaagnZeoM
b0hG4cohG96D/ErUmZQ672+CQG7E80X6ArWMH2LbDZmBAsVpr6XCS7a5ZTGk7uRI
/3WPu1+4rORQ/S6CSmU0dzRl+wU7sMidqpV9OJzGvtpvWgJC2CI5FNSz3JPkXedA
ng8s5/SgShkU05Mbkk2zm0v3687ALMxAir7gqLEeJd3Z1IwIjUAscGb7OFFhuTZ8
vGed+gYlo7DZmnixCJF2OEX0n8z/t/Oc93NeBuHXrt89fgxyMwUBR26Gx4FxuSs6
PsYXo8XdwWyto6cKPP3zZvvr6oTr0S6Ei5CWYb/ZaYGQTXKnt/agCUpZVkGslHaf
J/hBiFDJtBTn0gc9UpWSIr9d4gjVE14hQhPvNlUQfGlWTei6cfuEy7tAqin8hOQ2
sx3xi8DFQDMlnC806Oq/jq6NXoRxvZG+eykbSxfSOU+Z5aXWqn61VwFmZeVh3VgX
lmmvFrkMN8W8FkwG2DXzP7kvKtPSrodVn+EtdsScNlnN2lOmdbQ6cgj68jkaLWMz
EDHeWzhKQlocpa/YGI49mzZw0YLN4ude+kHO56t0RmnD3PbBbPlmXMdoJ182EGEu
a3wKwfjU8NTCaeEhLRcmAa/jWz3srY6livbhgYtm/Uz9PL5cQm46W1TE5DOnwq0A
9pAC5lQqzNYn3IGn3Wg7U8EjMgD9I9o2s2EQreRcOkYP8GQbHUfVbekTdaNM4fDZ
4QCsGBWIkM+yxUL9WLCMXnHeGNLarOBzuFnhfPXMZpmGoUhKYBoSG97TLp+iJlBf
sxd2/0a/HTkCWeWtSqMDcKAQrmWA6Fv0M99erwjBYsWvCj7yjnPqlQQqooky6L0X
eKkLm69qU7cy+IfbkoIqfh439zqnygwgDJ1qVnrFq2ahxgLVEUGIUTyo36PJLhv6
3LXVWx3FxtSH4X1LkHDjC4FaaMm4JWwlDeyg8+Fegw41ljxra/PAfecKB6Zx1lkW
1ow5mWNXCyI/uGhNxbiYsYkE/n48kHsrX27y0sUTFXZauQEcCVIWTaLqxVFqv9wu
/ZwFZSJiqWjJ22gGgV/P7JsG+K/DcCLoOIP1Of0VHZsD8W1Vyfb+CXhHpPDYauIP
qNOIj6ZttNHCwyZimAFI//EFe2BHTOJD9wW9osfMlT2PyvGGn6HVo3WG+ZJTKDW/
fnUa/0Sh2ATQBXaMtj5aBkFNr/S18BjiOOftfkuCAh+IOFus+pjtXwPU0qIEiIkU
PR7uLUbN2xcCGtSqTgaePRS+LQpByma5yTeD80LtivpFYGaBV2pjP+9uWd7smywM
b54JSI0TkSqqSHoEMoAC3/Qs7ZjVLzS9kOzPh9Vl+cHo+7oV0ebjltvWEBZ9y4qI
86HDb9IUVLJjNQ9OZQYy69tvxnsA8Jqs8RMAEKCKXO0+oPSlNdq+fqP4wVwryr/y
h6aeNdFePF2EkyiJEWJJxNutvLkDxtdXnlRBLp0O5K/x6DsrCKnYlAb3QepONu91
At7CuZ3LVf04Y6faVtJBDLG7bojYzF0OxJ5tT1degOPCYd3s3FbtA7+uKxuWOVWa
wG+6407Tkf3GIcPm6aAlnMj/NCTQ526zuVEfslafFBKqy0D7/RBA/npfx+GLDoTt
TjdALPrmuwh8xULKePs0NW4UVrTdxbamft4MRMuCIyn+Y/jMawCCp+e2Fe3vJj0W
p0yfrvJ8ixf5jQJwZGebLSbS+ffCHNu3i/3cnQdoEeFeF66IdY0nfwpKtjcpg7XK
MBZLYGu9cx5fmaZAyLY8Myed8NPTGN1/rXAfI+PrhX2qt1rnJO1RSYU08r9PNuoC
n5Id16TK0EwgE/ePikY28P0HKeapyrXZ37sCqje5mNZPN8QUcthW9ExqghD5QPy3
/1mvbasI49L0wJFKKUdcLuCWfVHbGIFWPphN/9QIyj+yXvCckPLG+NbB/017buoz
017URBZryZ8ENuDGMsza+SSxwAurBx3PeCrZCOJ6uvOHMfko1+Zh63WVm3yVr4Zt
s2L2CkrZhMRzFXpTaSdNJU+hSHEm1Wt1uMKlHkjPhvsjOGKzV4HtcWpCBFrYtIYU
JvFoaK97+gi5z8NAgruW5MJljw4TB2q3llTmxcyGs1brHsXtvvWYCRuInuzSJ80F
dz3t6BNELCoqgVRNjE0lbSGXTBAy5luYWFN1RDJyirHPmX6H0bKJG5xhPBUCu5my
43jsXbLN/YV45gU/91MgrTK2K3XIw2Tq9SLIZIX+EyKcQv6PweJYCZnYJiZSIz0j
LMaXXx1hZw5wjLfQjPI8IC6wZRzbuLV5lrT9PTEVsK1p1dY7g0UjK2pPu2VUAtpk
4qutA7FiZe9xf4+SYWBRJ73ngTnHysWKh5h9cOef1mrc/9aacik953NPuu16WL3j
kuJggxDSfWo3gADM+LOZfITHF2GW92eFFQasTX01OSZDQFjUd3QNiH42uYViQXGA
I6g0iJbLML1xXithlUnyXmvUO2vRfIviNdr2H/aWw+8eKFhC6qUS88K0RBfQZcAI
A4QtWUTdqoc3ynifuf20TSbMzOvrowb08r5xI8erOYOdsx20pmAglOR8ZMtF8wwm
PXEKuw/rI8B5EZJje+9I44L1f7LX+phusRHBu9PF+hcYLrOQ+V7cNfrLofReBVPw
XSmrDAdg9A6wXiHoE9iNQPtqIEoai8EaCeo+MdVlLwtJLug6EllJnjY/0OkdISyj
h9JHnpJbRbzip8BXhxb960P0dta0rQGT+6HRGm2qylQ9IbpkTcHlpP437cBSew0l
X7ZqtciwT+L6WsVzeIhIU/b476jI4pPR5JKwbtLeO2HOi4kF7hUBOgrdprihbXmz
tGINSDpw1d3E6RSaWSVv1QyhgTBFLKDNH67Nj0rjHaaH/um27PI3bKiJ5bMTRnBU
+aSw7mI9Xj0bt1mwFwni1yNQPWs8Hsc6Sss4yaoCJKZsMcaOm3R20yce7yEm1lP6
S5rm7TqAB1JckUa3oWFkyjO4ubu3UmmFyASPSi2NeD6Jt3j4qA/aFCm3uZ+43E8l
weZdKHwMYmI0clD92j2SrqBr/a9+lUk6kNdZqERAGh0yKYtwDMYJrIJ1jPSVkuIm
9Nca9TW/3tjKKVHcd7kOFszrorhXkb3R4LLn+XCI7R9XpC8mxdo8BBGjBLyWiTJ4
eVn6nx9wbRUsrvC96E2UnVuLyKo7hRIG1n2lnYnFtrzOYID6THla/9HMMz3qQ52L
mWs7o3GU4cDhsyyyXI5jx69Yhu3rl7pOqbaPxTm5T74wsoIpp5GcI9AkJwQcQF4A
dO3A3wUUbVycSN+I0Vv+PgQYSbsAjs5ru7kuuIJiovtHLHlQb0Py796NcmxIWliK
+aHc5P++VZuzmFlvZ6fQ03AyvVvHnHdawqNVksk+cf4cDexp0MmniopyDV6980oi
MzVhTWGIDj2pVPo+Pts9BWDW/G0Mx0oJK0QG6D87oxmoQMeupeEIAQ75KWqJSX3m
UhsV6r42KU3vrklmLuwGkP7Oun6Vt+vYIfoWWk8eZotO3MWAHSiOvGQ4ffXHNA9p
HX1jKOAcMCe1CX26li4ZVhSZiXQ9vCnUcyAA8WYlqgX9jft6zWegTc/nALyYIADr
zO5saF5+cnzKQ09Tu8bwwPgOYAFHENhzszuck//Y650Qh6VONTtPBeI54mGj3tCh
FMTHqfo7a+CblBx5+fmp1A4/zzQjvzxS8E90f4yOISqVDmdhFT6mAypVINgjm8Cr
nPo3ha22fgKJ8cArnPCFDCO03SA33YNPZBFY3BvrQWsqjHsDdTYKqbcxVwmIcGzn
DSrVCUzOLVvsQeDDEtAhRF97cHUg/7VJp3okoNEtmYJb4pAEf+W8C/MrKd1yTBFy
0U0obw9a1lUlxfUqjkOpmb/0d3I9wsJsiISLdQIhFiASPQdj3gmU9drnlbcRlxXN
QdDk2vhGhIHoGWfwyFd3xp6+twr0NyzOXavnYlA4eObiIqQjYqNcYIiZBt/klAt7
JLy6fFeeJvj/AJh6SOfszzMgmfaHEIAgUWSedvjkgL25roerKMf+tnwR9JyIaEbA
lBIYzMfIsn1zE6FmI4ksAQTb9FMbcYcEkpJbCbdcpsz/g+0DsIb3mb5nGo29/nJX
pqHyBJKR/ONlNw9UYIelIJlY+5aj0FARowNvtKTgOMxH0BuEWK5vOxlVMJ4Qlfx1
WhI98+HZaJtE/xYIZnlTw14CsXX+rArq6h3375Vpa4atEjU0VCui4VvVTCY7vLqC
5wdiWej7YUU+Px0aMhhODGHPdxYTipkUDSpNcvFa6oTkayFFx+qhvlsYgmO3NvXd
azAQPVFOaxO3GbmfuHp3fSptHxyiehTwe7MuifOJ/vkegYNGQtKwDgl8qYsv9Qgh
ZGXTOMjZASPaqpOsFenhULCokabk/WJ0mljJ8bhngEgKNndRSy92/b/ZDUqveGy/
jK4YLQnndFVD2qbVZHNqEXuzUVQRh9d7F3drl8tEIpWtECWOYfGs7WiOO6QEjiz/
81ZTzf0WzsVTUOSWoTyR0e3ZOS08TAeNLXJfEOu24YsmZWEIUYg/tNDkpyrNe8iQ
AuFfNhnH71TRRxrPMJbdX/Mz4VaO0bMcurLdH4UnBfRcpBUmA1/dOvdx6h1Dq5QG
0aH/4vcAH85O8gUjiSta1JS+LSyqXRKwxxrdrP4KNjWr7Zq9RySWFxg6bsZ1iqRO
TY7RbgM7lXsZs7Q77N8LIvFxjPEiH0p5W/ixOZaUrl2WLxP8Hpju6YlDETfcze26
uGH+CfQDDK1P8EDXdwDdeFllWrAWQRBjdNENZI14+Ro+ZkvSdt8q5jMewT+cH8Bz
3uKq4sGlG9dDpHO6DT3or/K8ttTT9pHQnb4YAg/V7l7YKm1t3mmMcDuvl7T91dwG
AJYHeK1iw3uno2nNiy9+W832bQmEQM7sR/SGd2Gs8FXQ0dcO6+nM0hS4YiPmiej+
93qEYi9CG7tA71qOgRqBXUm2vJ5IuxiQjkVyGFozzVjVLxYn+ciB9t/ZkgV/N3MO
h8MA/In/4XXOy1YQdn/XgcwCnWd9TmZq/MSCI05fkNFMiRmaIxNE5EKz2/m4ks8e
jWpQBex12lp1+xv5RfpTKZLhmMlzIL5frX1Mh5tZzyxjgjAazbOLdYX2vZi3WKLY
HTlyP5ZwDLuIoaB3qC0odC8N8XDHB7BcTEeLX3OVFGEhKfTswbZhzon2Owmfpamm
+gQPehu8fxBd0r/eCU4i7v+aRjS9+mGrFtonSH39xIGJwzP6cXarLD1lrdfppfpf
bcjQ624RqwqumBwxJne2R+iK+1FNnNPAfJT6SmDrW9bCtdZms4GXwa0FKiqFXLGe
VONoSzH5NXm6zrKro8MiO/IzVkHfR6zz5dhTlr/CMGl9TS7oQB28NgFPoouzs5VG
+wkahB/Trl/uS2dw9HfTi6JMIt2Y1nsLz05lr9HCy0lCDeUVLe2DjlUrqGcX+0P4
BVsrc9kIMBy73aaHXP8PHysmH8ss+UOt1lP2FWNV6gHX1W7tYtZ8MiZo71FwuP4N
i8mYIb2+WuKkE7g4zbip8XNQx0WgAs6F+s+yBuf1BOQNEgttMGbe2XJlWCmCuVXT
DgD5qjnzLN6Of47LPYAOmgpVJcqazXUSWfhTkfEV8l9mPq8Z1b7rh4YdcaTwfIv5
242EaOXRFSnX3VN6oNp6q/rKXAzAZPMMVWI86e7RvJg5SSK+VW1OdG+HCwWkX57i
W0p8YS4RlVFa+Yb//yEe70pP9o5NEmN1vwyVl+AFBJZF/bADcktShzVl9iNiYAMT
8OtDhVFHTE3zbhOwUOa+go0YZM58TomrVNph0usnUF1ySYeVmK7XYilIqTPlwpHv
7FUJrGO+tHM0Ui+zZIlaE9YWTyFvuEDnYQO8GxiklmbFUuwdAFPUvKYyAz/o11RS
DEp7CmTP/bvDkDqck4cDo9q05dhEBQpYOGxyZUAaG+P8QiauuS15RL3hcbfzsoQq
tSb0AiFvAYrohKzSCDzkctYykikUXBNBvHt8P0hFkiARfYNeljG50zpSKxW2QxHK
pmG6n72LbylQtL3MpzEdpkpeL7d7EG1AlkmcuKCbbEPAEt2tfHqwU3CiexKo0KGP
E47u5i6PdxURCww3EfCNFg+JYJrfoTIPMhtjDb+cdOU16sl+Yr6e2BF/BAcW7Dhe
bUweOsD0YjM1Ma8JCZNfLQUnYxGxxPF/3bNZus+tgLUFbhpitNfvIogiOphVOvpq
XxA+MLuMbg+0s7h+2xcY1yeZsG3iBhJWtElXLcjmIO/49pGQ5NOptEE6p3ezAWsd
kYIKXtcUjIhpTasHSpU9muy/3RhkyMzCxGPpFfcsAu/qTd6hAv4p5vbX8ceHMzqb
4l/b3jYjPcY50pUOxztzZS99ZS4RMfjwA5MLG32PuzglNhSPLHD1MFqZrZ7YaZ4h
huXieLba0P/CI/ruBmi4rI1vyMiQq91406vJW5qJulB1q+ToYC4ZwjJKbaTBOFzK
xyTQHjQZit33wpDh9m8M+hBw6tmHHqua2Ovy5xSn3/yeaWXIpTkE66g9xNU9B/BF
sDMtZC41i7o+KTclR3XKRLu/QT8EvgkaqGhxM/jlr7xU1ThANytzi1PaWYjaRo0p
DTb2e7OGRhsz2VaDa9zYFJb+3nfhIGo29hayEqlFgwGeqIjBMxOGvtebp5pabHe+
xH6ie73xUzjenY4s2NwauYmqs5QmTpsc139TBotn96CEQ8cp8HqiJ7Q5sOammSFy
5IdPN2MOlMXUGx42ccNP9I9PRIg3hsZY2sKMxBfKb8qRMOIUTqizBsGy/pH8x1FF
R+b1VSWD7N4czd7wVMuhd8CKESgU+9wVaSUtVtgIuO+e3gbkq6KyPG0X6Vvqudjm
3qg6zzAE8czAkGdMOGoRl16i1fFpvYdNjcDE0WoTo4XDulLKoJyXIA/johjixCfx
y7ijJ6cUBN5YUd20HZepxvJUCLdEHhMXG+FL4l5vLkMMKt95MOnVImmFhJcgQQEd
iZ5H0EsjJF9oCRKUZJW9cu8q2Ec/iRXs+LTmNyUSfDZY5D/a/Y14yDNXwB4hgbzk
o1AY+r8Q9MGWUI3Fi1kQfCuvF+yzQqXtpfpXXQBBX/LZN3nnPQCe2ZN3PdjzYV5F
nYrR2pgkFKLt860sl8ClvGSL0wL70hUlmxyvnbWj2a6vMAVQFKpxEl5vPkQ1pJlU
jGa+M+sr5Q1ewz3oEIkEnyxegL8+0gh0pzSM3ed5um+nOv+8pOlZpoZVlpZd02tK
40b0+UMA1eGZg3sdW1Ci5ZgfUYPZdfwZZqszi3Pn7mtxs5qFh2P96HKnRhQRvX5X
iAoDy12I1XfF4BoerWGdAgSQ5SVzV8dhjqQWq77qm6BK/wLeQ10V7WqrQcVF3fsJ
1I4Wjb+ckgvhLzaiX4GLoPyCw/9w/vBX2Ksxse5b84ntPV/hpisMsSXcs5TaAnED
yBdRLfInv2yJRe1oVHRWzYmDXlxKzpbS8mwJyUZr5FrNxX+WgpkPYOwm53aPJLyJ
hu/XzO1lPYqxUgEZX3ztbdR64CWnExF0O9uWRxeYVNzNYyDZhpQy25FmKBTj6jkg
0GLkvVOwOL0hfvgx3M/qdLYYi7JTeFBUS6OdX4oI+sUlSjh6av2hsQCyN+pKIUY+
wNLlNitkCjFum+ceXU8XhU23BYnmJ7/MBj0lbiMoz5gpF/fJyMH+BJ5Ox/ngQD3R
igYWU8AMliSDPC6lo6aQ6s57Nnq9Gbv2yaoBCvgZpEYfD7UKg1RzZbEeWazpPfbq
ENu6bMZoOCkDM16D7RMAoUM7BsZIjNKmiMkDWSOT5EweHjqHxwxP6VjusR6DUF8I
kSjIIvLfr2LolW5vX7CzJzI4g5LX04AjkIxc1zB+2zdUNYImgyX1Teub6NczwrjB
s6Th3PjL4BpvNwL1LYLnc9YBe3XZF1+aoOMQ8LkddwmJLmsomnhya+aCzQMCB0Or
vNEWem0YXplLlrdXzeaM6Lt9ts4YIv8snnO0Sxx5N3yyjFNhOZ84Cn0RiwIeElZ9
J3wYI2jZS5A93pk/12/Nl5VKPlkkcl++6aJP6ofxBIdOrrj+pbHKPadnJ/Ujy9fx
D5/irGhPLnaP6/ziSgyYhQXXWMpgo4758FR8rCNkz02yvebLdypPE0ZoXZgBdzwa
BuvM+ooDwopbg9/TSouOR9mX2FGKGqBEkv4xvov3jvbHsq/r4mls4+MMzF0YIUju
wMoDB0P1hdeVFL0kwUqjlCOhwkL77vCS9OV/uYxMfvNmbAhk+LMCfTTbD8moY5lI
aduhUciik9TTowBy3+3xTUHn/RF2CGoV6P3I3/9bsTAmx5h/zTt4EuZrnA8eRTnJ
Y8nULK1TQZT9nthtAU20tffXSdkZPMyB25/tEEjinL9rOA32g88N8mkL3or03QIi
ANZCydrElcR+WDbqxrqqhLCv7pKZSPeqDo8FESEZZuSoDdf3TInS5DxH9f5sKuct
Qy+bty0gWCNL9jGOxiDmXoIiTMTqLln+dprkXAXqSDOMnxVS+iUWdF3FpCBtOha9
3+4eSft1Z/C7Oy44ortGVnEPzmqqgEQpxBR3iKzllp8atWnzKPOqw6Yo9035Kh10
Lk802qlUpqGCilyKjD/MtNyHY9HByL67R4X/JjU98fS+FGo7/v4cYprlQUYA/igW
lZGFTTxMTfIkVRXpVzlqudA+6w+iEeUqt5tvSV9zWuhPJtjAt7Csh8MXoFAk5ZNf
x4M8zrVou+9v8P6MR3OGrOtqEDV7g30SLygee5YH7droBPmiibcBQ/Xc7toIAI97
JB8Cu+MfKBS2D3F0uQbSOQokX1WgXPfJ6OnAptY5dFDuSCnaZW9IlqINK5adYg8j
W0hf/6Sf7iSz311bl3+apj+NoelZw+lnAYxzk5n1dtRifkClyZrxPSOm/WFXeVUP
Ttz+GvA5eiyNPbchzj46VhoG6At2yGgUNfZUdaJ3Yqo2XixKlEIuQFJNenCKCZI+
oY1kwe4JrjdIwNszh8bnO7feK/AVLBM5DVY2OIAF0WwcH5+3bs8hLNQcpm8SBLZg
cjmqPdCw7iaszRKFOmlA/A7PBoupSlFkBJO7AJX9Ls+IkyUxZKeZgzbjz4J8Jc/F
wXJlUXCVdof7kgqbPS1nBxQodMTSYK1Q/ZtY4LwBWLPd3d6JQDWqnvUUVUbQAYlv
J0rPzcAdc+LCmjbVdBVxUw07V7U5AvoyGR0AaR/kRr6xZfHb2w9Gox6AOGDzrq7c
ARYgZEFEgInhiWxd5elSYeO0yPtsuSd4CWeGISFSV++uDAbXL8FBSt/Cv+VnYFmG
QHL5VMk8T8jCPrcOKXjmrXjJZOhJPTvjgWg+Zj6FJLsstCta/ctO7jglU+EBogZt
kJL0Yuxiiq/gw6qeMNgurL1reuNYL5yYxh0hx6oWQa8go0xxnDSVYj5BqYROzTKo
MhmiUDhHup+Out0uA7tx94rFxXXwD8CcOVmxgQBP2NaUajlirT4rA13zBSGdIAII
Tc4j8h4m/TG8fCh9YUSkcg4gAUIaqQaLnfMi+WWVt2RTByEGsltq2q/r2Pzh9GEh
p/eYJZf368QJYVRk2KmqD+up6KbimbVFW7soDW14tChWKbMkDHehR+9sFXjnTLV9
agr8mVw3ktQqlvbF+4QK07aN3X9uXt3urKDsVmckYLweQoSPhXQPx1xtvK0PraIN
FZXGKiBZhgNkh6wcvSN4s1DdX2qGHIRL6ucDr5l04gWgOjCdLHjFnPDSEav/IGxY
ljtT1TUJGcsUTa9swV5dFgw0xpi1Ntmo+i9ukBJjB/k4Ek3jzRxM6P5uquKSncuQ
Xw34IZNHw6mZKuJkz5Gvd8AKEEiP0g4C5qtnvJhv4POzhFYr+2CB1zMiX6xaeTe6
fnaQ4HGu9fyPBId0xhNYU6WGXwsfTz3fE39X099++qDHDJd+lR/FtPKXqxl7+4r6
/d5dPcw59V/DdJf0sDZh1wvyx80RP6bczaH3EhiseUR9Do7ZLyKJtXAfDFvvTERK
aNv4/JycTVwev8mD8O7/etTn+t06pvasthXH4l5VtD3vsIyUeGxdwcSvBdjIdRkM
tDXRBxlvDcCF7UHAWj5zhuftkt/CECAtO+qiz4bAG/FHhftYWsBp7mmppdFPAd10
RQ6PvAjK6b9buFGbeelegS4v6rBKllB0bDbKE3T7JjmISOdLbUEkw9IFA5LCLUoe
ODdP2QKCeUGWNyFO4Tw8Utz3medENNg8I3u8vKrWwpcNVWzE8/B2XHcO9Mx5dWUY
3yIpaD6HQXdJAqMlt98+nqIiLG/EID/pckatF3p0yz44ZUIy4yNs4hs9SItqOUsB
podhMqHx7V3xB0KQ5fQ65a2rPX2Qk3Aeq+CFiICTaifct++QUyiSqXR2tlHGooez
yPqXXLbClDKe3B7pWJJMmWJm+PcyYNlt/aRYOpFpNSZXqIxyEhJRIP0YgJzDDDRU
D3vjNq2hN7FFgZgWyGAXp5/o/GhqYcsB6+mvsXgpUy4gpxwa+LRL7t+QGEL/FiaN
KhO0O3DTYAht78Xit8pfAyoH5HKg3CXI8MAEPNGQn1upMiBOrxy64qgONs9TfDBe
zqYE/L+FRbkSvyFOy4IGgSnovnPb9i+chM9D1o6FEkGviub1ATkm9CDVwK02QZMR
vrD1pKZ9TUoe+jxIlGPT1hWG1fh/vLRjBGeY/vgoYgwJ+yfxtQgxAa851UKMmCjT
Hi0q+GCfnsmYGe6gMJyQIWqDxRo6cFWC8gstRI4g5rl/NhMJ3OSe1Klm1/BvOsfp
A97Fbh0zWPPJbv+Oq9HBYc7HccFOCbA5N9W8BBCwUIfRsbXYFnn1cOAeA4uCQ3rs
sYX6cC83oEjjhP/CF+gdD9cWOerpES1sZDav0ma8BJsQC6Dl5qdjPFMHWWoOD86N
lzLDR5nDQNm/APY0NpT6x7jGsMWi35ba29jV7BnL/qXmDQt5ZXKIAq58ZG+xTVvs
f12oKjbMtFBmTgDBSJqUcOPbXOYToOhTPfyf8Ds0/VMhu2nKeYAFFUDOTBXvE2hf
QtyU1tzSPVkr/KNVTb52bjahe0F4ok3E4HQ0z68H2eaiBFYgGlti4yuW1DDzRSgZ
rS8+O7AvyhCUdp+cnkn8h5V+GguxkFY1504u+8x0n+SL71P3brelse8yxVLbIB9I
ojx7CHNVhVXZf+/Hv1Py60X5GkgHID98KETpjLiWJCu6TpwT0xLBOMQV+hLVx/p+
By298AUSNzfKeBVr5Li7CGDn/YRgFeUGQTY1yDdIA5fiWTpe57DHKFYMhYiNPn/s
Po2BSX4wfhtA6eqVYYjI4C4xD1vQvin2HoIVLP4pEtMR6fKgytgAwlx6bCGlgVvl
eBpXcPPBO0oDv7gS7s5XnFXDI8IzObfPdBY248ARhOshhd4yyv45bTcMUvDjuiNV
endpOU1Fy+aTHtX5/OnxrkS1WlGGpJaKTa7wj+DZnhnXRlpbBoRHy8thSyGc3Q+w
/InCgHzt3By89lFcYGR46fjBxeDWjTd2RcYB75pe7Vih3Id9+MM27lFIstM7C3Vo
H5WM78IQkFda9l+EMbkRBDBOulwWsPAe2lxSjpuxTXKCxOm6jL2JyVrGKDJG8nHB
NMsa5qPW34NBrXdC50v6yPP6l3OYPfaivvmtkdC7PFgwowpZSUGqL0NWVf9BJJPW
sMBGNGHiGYAwx/7Rj1m4deO0XGpCqH9FyWHjupbyQyEa2AixmGvYV1Z0+3Ms12ys
To6XMnllUPp/8HazM5womyQsjiAa1916C1P3BOYzxBq1U9cpHr3HgW4bPpVs2Dnl
u9rbf/xpr6+yBKusMOIjmiMr3IevI5qiOoTLRgnsuItLB7LatpLfWIchwhmQoYUG
AM49RvShkTti6KDcg5Kg6TpJ7G7cqY+U9o9TJCZPP3wi63VZM2nEGJmM9mTdFhIm
CFqsrl/Qg5qGw6Kd5K1hg1Rk0ALrQgoRMhJoR39LuJqvarx8TuWU2KQDcamKYxyp
VTq5e9oTaH1lBMZ8q81O1B3EfTMnvkwpPUB2yyQKY5ukGCap3WV85lNUs1QivS43
tX6iuh5yraj/sARNwHd3sxF1dKxnSE++mr2CKj9G+szQDFWn4uueP5QK/wM08CVM
o9KYKZcVSsHyPLRRlcNGr41Yt6n/26A7KUrUwN0THZ698JZB2Q3FRmzuWugoe3SO
obZ9b6n/BfbGyprxau6n2dljqpmxDvd2xWYipwPoxCHE7ZWb/Ojpbev4fExjhhp+
FEZSdW2vp/hjvK1L8VJSHZCJRikqwE2bQv0Iac0SCOO3KZn3qiUPdUjHhoy/x+dw
cA5JTiqwc5cyLsGdhjSmaDMM/g5JXyQ2RC4hLwQawa0Pn+pRVtnpm6qcdOwguBiu
8E9aQTcaNM/C2/SZfUpmormHoRI0o5YWhRTgSaYjkAH9XNLnDBquO2AGKpkczlMU
jfaPuVM0/Xg2XGeFb1sMa4IhJOPVSUnnZsqnqfUpVLNJ0hn1B/wEyfFHCPK1rjv1
tYs+wA1zltykEV3/8tupjnhXLUI5pa9B/iRrXloaBg1kZC2aEjZxnZubKHhUW3Gd
Ugo7cE3kidfAfTiVfogWDA9XiRi637KIOHeGq+3/DS7/KH4rqB9H9gDp+ysUAMq5
8S7Px/8r4vq2qhHU66rx+mcwdxC6GX+yais8oHQgJOLBSZ0v0+p3fGYN+h4x+j2B
3ju+p1jHAfFJ9ZlFLt2GNBNdcsD0Q9avq8SgdVziDeTBrFZoNKk5JggKw7Age/G7
nG87C6CFhYaCv6BdvEXBVo+wV01RtuC4b3D1zJZH/4hY98NxLhJyO+Io7C7y/Rhq
w0Uqidt6BYRejSBAruSH+poFpPAUdP95cO+VsqcdCDz50nBKpDVzidQgo4PkXQpS
EY7V4pviI0jSmmw+zfdEsGsj1cZex0R6AUWCDvfss8JYMlfgoPGH3vAEIedVvjeV
K+xiMXdT/7M1VEkANRkwi+e3UpxVSnxLIqVucWhzVpkloAE6LzHga/awuqKCojEC
MPh8+bLYvf7VDmwf5v1rn1AF4B1m2V0EcsVrw/bbcEs2T+deYow+LsXHnaUsiIzY
RJICoWmAs6CIO7fwendTo4ncSSuNhhPHxVmYTHd7un4nYJYJat5yZBlXFz6WX23/
L/prlPUXyo+G5v7hb1dtEq3D1yd3dfW03UdspWdyWGc38zs+r3GzQGahuv6NPaMs
f0DeW042cYyqTAl/yprUn7An+qAKDFSoTO4C5LjKb7ebEs+3IUYjycaQWsgTfy86
qWpiApiIeHilGgc6TgKqXP2tsx79EmUTJvE36EOeta5LcIbK0VlnaUNrLAwtzWtF
cdenU0wMRJYnt6p24hIMIDdjhBvEk7Wm/wA2POexQ0Nh40Gw0gZKdMO5MLZnXstF
YAGWVnXXClzWp2yxdaJFA44XDvWG4A83YExho3FOCfc8tturWPWYscND0HmwD21g
txYINia9W+0brnv9XfFz7s5SxEWOESp3SCuPDi201rQQ6FNjz31zm8oMc0FaaLSn
u6OXoopPkVq4l3enwN4D2f7HIIrXd7Uu347JuRwxEK17fPmYWazslL+IbJJNAkHX
OszXIkw6ZveHn3ES7i7i5LOqXga+/nPwPAavZjWhU+9i7TgprMuH1q5MXN9GdnxN
1UQBszdq8OFQOPaNWboKKxas6Tb+wRxbnStK1O8CA5CT3RB/orQXuWqZhgLD6c0p
4dEAvShaP4TzuGpYWYzTuOvlXNIwJ1aVt50bmlpc5U5m9zq32aefwW5hT3PgxxCd
xjn29cRhpzWx5qzR/GRZF0mAyCrVK0Qet1NUckvk9HtUaNEkOXa/nqayf+96pP19
tbFhc7r7onog206CUScpKsvLBgfheycRK3Pfa53dlaXfmoMpKW24B/tGupsKwLi/
hFY6/GxmvS+xNWlXjkdvVfbmQgs4ZEj8hmomuc4DhzyYuk1xUtdH1ZFdUo4hPEXp
EC2OTZx4ZNeG50cchcT1iJwZRhDMVfqjzo6NAgGwT2tRWGxVNpF7gFgDc0M5dyyl
oPVObQL8EmQSV1sxvYpWSbbWfsL6HyLLILsuuGNCqKY+gs+djanOik+Iu9/AnZnz
534skNAPaD8jdfZg3k7dLCtE7tuAbnKlxwTRAcfdMRjNDs9KQSEm7El1uqHwInSe
SqbGwpUj3kFbBHRJFAoqaWFu97EvbSVyjbVp9G/RE76x6E/aqvnptJUEoVgOic1E
4CdedoA691WSHF+fpPpVpwopqiFQrNKh/YuncMw99C0QW8dAE4iek+fdD+22lUz2
F+4W3zkA8k8tEeASz7NQ+uQYCuz/g1XM4yXbChaJRI3lYcZswg+Tz2g/OrfLtd4h
j4WURSC7xxPoud2zw3yzNKqImTYZg8cFe2Nmql7aJH6MgbKUGXje+m6iG195pLNm
Vf/HjJP6KBPBaDmvzpUm2M6vFPriixUpm0gSdWUWRC7O2IJPOlZnPED1l+0rxVPB
4A8Tg2JLa4TN67t4GoEtnAhvhjp7PjgltQtP6JLJCD05I1Ick+mknkAH9sUBjtOC
mCx5+TEeWkPdYNcdIJTYKe6z/vxRLxeC7SqCENBARFhkjuCwJKcme3zue7ltSAGo
FZStODeD6xVWA3JHkxv9WP6HJKcp4Whmk9tEKAoZqQLmoCkv2NlRWUVlBEJfZiR9
QEaCb+RAmW2CMaDlEIuariDt4oi+w4pcWzNN27BSEWrR2QvCjI2Sxu3wdLgngUEI
muFEcyFia62pn+I/gyw3P2PmOVuFWaCllU0uGpGz2XZOYZP3fBv2MfwUqW1BzWcm
fnbnolzP5tlUBvcNRoIeRCHrEJ6NTtBnONFkwLge/ZWJii1CmURyafkc88g1FLki
/MDaTxnQcoACJPImfQCB13VB+n4uXGYRDjLImgE6Fk3FSElVvP7epn0NtKBX6ZQw
3VN5KIBVP55Pp5zgSKMrKgchgzXVkQouq1cgMcLERGg1ny1u1WTYuBV/EAEMGgwX
Vn03eUFHleiZb1TsB+Vx7y/mNlnK/+LdRa0xfDP4sWzw14CsULjKa5M/Bwaa80r8
bYQRsj9xfXhR5oIUwmwcEIl00e+eHgB/r0cTw97fdLTCI9qkJtpy/O/4iulOY+QE
EJLOP84lOiRVE2b9TcGbH5o+2sqUlb96Jc6iVvysUSFqglsPNFw9x47giSFnVH8O
es51LpUKDqWd0tY2Lrh0zncOqShvfCQc2p82iQYLpSTla3JvE63+i37djBQSiHVx
+b/RQ7mg9ZojgP6KZ6OhGEQB95StuGe6w15IH/tSflnT8PO6xYagHyAFv2xDRx20
RBIqDgg+cmWN45MyPJ5v6M6dwV3bkPekJCdOdPEjg8tcu9dI709V2GQqUkvOMeQD
j1rfZureUqSlNJWGoxtB9XzBbTcad7JrSNHA7OWyvqTeZ5kV9fSFAwQHU0xXxFrL
5J0a987lN0OzJyHtLtHIC2br6aSxgWoP/oh0i47KOtuBJIpiDvcW0fj2W6YE9qp1
PV+hDBhhDqQ3YVVo1lSJW63llJFlXFi+121z7WMmBsV/bkVm/W5fJdY/+bjOKnKP
5OfQ96g8yrsVvUBbV08mK1k+vR7HSemXMwCDgqM0EpQgckY19W4x4w1/XdM0eevZ
ao0NU786H+LAe7PIWhLs+wJAlMGYcr5+rtovWgziHVsk0HKDTgZ8CGwTUuW0k6z2
kO1xzK8ViZ1QR5p8ySE46ee5XffB5Kg57vs73OsPOTPeQoorhB69kDxi5C1mdtb4
ALSj2b2x2C1QvXZahsBamANMuy3kJswRtjrOpqy2A06bQqao49AZgnyhslQ3xhIZ
16VfhwoSrkv8VVyPyhXOaRzdOfkIVG2y91x3aJT1Jz8BSzXBg1EEWPUyKXI8w+t+
G3RqSGCmWnS6OPdKSa9plW+5RfwSPEnTwHoi9Red5vNO/nqZQu8kk7+VjwnEs+Po
hh/yawQ04j1cslRjfoa/2rq2+JTGqHc235CSpQ98kdtDgqwBJp225d4W5EG98Eh1
udfk2XF71aINKoXTnapuZxYE/ozpCKd3y6ZUbOqSqyUP2YhcEIGN6jbjgNWvNKTP
z4Y7onc+zKzaZ9QxT+tco/PbInygLDrzogD5olpWQRoWK65HWpVs0GlYJIm6HEXI
rhG8vC9IthB+oYh8UlubydegVHpcmeTMmcp5JwCJz5YTezqvAHZS7KOAcFpAnhIF
85CbIk5zRzfEpJgeTzV19XaXUZlyws2XkUNOJpZqpW4bKWx5MNK71/YB2xvKIeFG
eHGMSV7Z2QNuVtXmQgoCE8O1PiQFUnjQE+aX+S5NeLOVLjxGZZj95AF+LYEIk88s
I1nYDNxDYxDP4R0BTSJUqeRpAU6s4K9hkqA0ZK3Ann2flySrylmIpr0voEyylolM
pDVrVZWgnCFP6c8SswjG4+01DDlaDLoNjEYCUvjC/AB3uyVeKutXWpoDZsGt/eFE
D939WgcInT0On9uE/LYTfTglGJIZwAlKynh1DUkB1Xtz3k+WnpsW7mz+Fw0mrXkJ
DdZ4uOjrKAKmimDVKZLXFuoxJNk9JVQx0Bd3Xjg2lzU2r9ghIlWVcQNoIZi7MKlM
Kl/UgA5ifqsuQ/b2p7oA4Cy1cFysZmiWzy5p6Adu3GLJW5TFQUos2+6m0bhslYFs
h+OL6Cuc5jo5maWjmbpXWOb8OKgLOWp9pjZ879Q6hFND8cWnw4ZviHLOQVIiLNau
NkX6rZG8z7kCNaBgnhMbKwOZwqz5XYb/zdMAZwD1/3ho5HS+uajub0ebMTb0BC4s
twhZxYbjDdxLOMaNFPpMRU8aA5Ey65ovQU4rcdGDMVq1VzamiqetX6fbGZXVUmtX
JJl4AR3/jWx7Zng/myKZuZCG9BdRkXBH5JTrhDwDg96hLbLSHXad+yPdUWWrMF4s
Yt+HlFML9b9G5+04EyURK5ghnmSuwjI6CNokioP+xV6R+Lajam6BrUeTd2cNAKwx
MZ4wyzzRznkGz1JwhkAPfUTrhUDAHSyI6AEy62C3C3MLfQvZtnVf3DfdT/2Ic0n7
VXILLk+ya+aUaltw8yNpAesL9VzmnsY61DoQlFrp3blFBI89/itAgzTbkIG840nJ
Dx5f7O9hOhfntQz8aGTXKYBpWK9gw/yolvCR3gT1reYMUgD47Vh1F+ItvSF80LtC
yrvd+Fs6kslAaePfAz409xLoWwoRLdwFISpoHitrTIjN6gFa7V+a090x6si3BMzG
MZcUfosK24jIAxnpLR82KXVS+wou2nLIt2eR7apgWwhgnUB5tDA4Teu0ayiJwkAk
/t3MDTyfmbtGiU8lLYOKTwOo5B14VFJpybyz0AA9WyPrj4KtWEiQ8xt8jRbnlm00
oC+gEMQ4M6CL6xEiNFkNNUYQ7KlRM7NXuS5cIM9YnWcR2hlg1VNv6PD+sjT/VNd+
Zdx3N64lX2+mNug0HHY9yeMg4QW+AO+4gcJUEVf9Js6OLcz3zEkj7piiv47YH3Rf
H+vnZFEMHtKESQhqoBdsqgmuRiwDZdPGAT87wHTrsQCE5/CDmO/BUTIDcU9/kngY
UXSVInYv6ldySeHhi7JMaLb+laIKFMS6RfD1UkepQGlJ+Um7hhOsDMm6Jjv1JGd9
HfF/OYPpzbTHNe4pv8SvCRZ11evJ/hFflbw4zKUn2H2BNFh3zRAA8STzlWje/XFC
Mc4H4/GBMWVArFgazYzlz4Rbt9J8iwUDAeQN02XK5O8zOZjy6IRCLby78e3lKYQQ
CaD/l7LkdNm3/BQQehF07GNG58hvm0FL7lxVUe5CH9EoB98nBUP0g0w8o99ql9U1
EDkC1/XJCmvLRwKcYtCv7/z9a8/aCC3ejNMYU3bf0kRNsmgSP7CtOpXNCrP6QYgo
QcawxY1R7y+Hy94KmvO0Uyn0F8/A43KmGiXZZUKqpL1VqHlEBIyjc8L5e/+dy5Dm
CaT6Y5FeVJppPpigq1C5PxWXh8Z7EA6M+COvwKzDTkCDONl4H9SCmtg1YPQmmcNF
MmKZsrXezQLZMgJnnd7eWtRYkd+fPxEeH9si/T+WzmzAfmCxbsDeOnGz9xbyQ46Q
qRVNmmuCO5ZuQyj+psI88zsScUmKwYJelpBaSekAcAbbqGefsvQaX3ZV8QnSHjPL
QfnShQsvSORT+GsmPwIufeQrYiKO8qmILHnfqIjFU6nxpl7I0KIhODrVee7Tj//O
G8vGWcW6LFx3lOD/Wdct1aU+/7CR0oUhebaIxvqYBaUFm4zh3DniGnnswRczSPTd
4hG5PQNFuXgaWmYCrFTXW1l1g0UewgP1k67vrgxiB/EQrLKrcf0gjIBzmd9UusWB
FzUABfRSdWy5D5pjt5gIRNH2MECfp/otb7q2XtFiaTTt0RR4wA3UViZY/afd/Aoc
uBI+ddPojF6n3ZbTKoH5ufE/VKI6y0cgifbF2ZNnSFVYDoNhy17eo/ilcC1kscPR
ct594Q+freE2l6xfEGg9ei1RjieTJyaZY13wDoMXkwLVaSW3eoa/2va/1ZidOb4r
WBPyT8mP2FEAtTYvUnEqc1eV5z5ykPOW2Gp9XrYuQrcFtt9Wun/ryyVkFiZG8KXA
QKaj3FGRGBk6qSM5iNKiJsUo71n/MY1xA7zShTDc1FcYCQcTOoAAOGAA3nIt8k0j
u2uJ4vei8+Zm5LBLQNOJzOo252zOAtxXQSr8M9pMNtLPPTBtK3h4hEUfwv7/YF7Z
Scuhyvqn4DPt5mXSl9d3+UzIuJ0A8D0TbrzMVBILz8S7kCqRuxlrysCc6TbPE2KE
DOVV509cP3x4jhwB+rPQKnMS0Txe21Bgn9RHV1GK+AIEruHOTGLNK1kuv3Npyu5m
gXL/rJ8M/KErEp23Y74EXpDc1Tj3+B3463UayhVLNU+B0RKiW0DpM9NndtYJ7aLS
gsXurwi7dRQVJ+pWeLwwsriRoygPEHGBsj1djvkna/oWxxrMhayqF7dW9fUE+nkH
rV+7tqeiOqlOI94Bt0bfoRkAhQtC+6EBUZtY3Rf20gtXc3kNWGup08wIdBuFevhp
JTKMVD22x0w9kp1Pb45uS/Pn7fVqIRMYJKGkv7i2GrdgG1Lt5Jnls7uLGam8VGrk
ZzrF0noELPfoII3kWKl5dWZfwyHe+Kwi6BeBtlIX7E0BsxV0NYexI8SZD8nuQOSQ
S1LUDguwHiMgl319Xtmlo6xiKD4pc5FYnlbcSgBgM6LU2hxGme9dGFQhluepvV+h
deY+JZ55S9ExLuHuiBCEXIVFst0IVVnzAaGEzXx0PhR/ONOn5YtTgyts0QxpqWzl
9VRrd2udGmCbGTXArjUE+t3OY2B3mYeHp1sMLNGAareMuy6FCy70cRD4wbmfJGcG
yDY5vSZZEswPSIXTUAmR3K0utmYn/OjPyGo8e7J8S0HpNN8p8zdDT/zUct7xD0x6
2ASs/81tCswVABSY1qOWwTrEADwooJomVtfIyf1L7pllVkhe19j3Nr0BKob+FRJ1
kLE2LeRay8jok2s+JB44B25xBHhdUVbzLQHjixY2Rx3oTcoDY/y/siwPmj+/JMzp
sTnBVXSZ9KgyyItjbQSxZy+hxht/dyXer88v+8KxD1EvU7TvTRLLFMfgoMJEpGzB
EEap6pzAqcXvx+geSBHq4Dn+ohyOXamaC4uU1ly9iXqaaTde6lTk373oKo74v/uH
yn5de6/XWkE8SNKKyO9Uzw5kl0Ov+fYSKSVGfZhIRXRAzv+kUNkdL8jj6r5MS7r2
7Z2l1weX68pMzqRmbeSEcN7y2V3LSMXOHLJE09qGEsY8YTFXuAS8cC/ycRI/BnKo
IMSYOV3uH4UWzQ8+1E8gycnMc0IlcKXzKWz8CuSkTxJHIFbTL+wf/Jm8MOumNycw
MeYOS1YwIyQwLtgnejwRO38WPqedQMfJJBjS1XhDyPa0r+k1qcJEuyAiabu9zkM3
WS+S+mP7mI4u5dTfFinMowkmufbTFxvcRI5IgQAXIktb6EUh44nKsa8WdhkRxxF4
1nEE6cIRDPow4Htw+GnuN+wtf4nAteTmldyyP65ivXHlsCFgijWvxmnKAgE5efKH
IGY8kqlVqUKSavcYRYKvaTJ1ztXbxwRvCuvcs6+oTx7wymcW7TzM7ewR9uPtgYSc
6uphSfuLcdsPsPaJI/ykkeEZTT4ijxP1tv4iGgpiACPHmJCrBbVoTnOIO/QLmzPr
AiNc4gRe8rNuHzpP3g6we2CnRENwrPNsPuyJnb+j1rlx5HRxqNwiwHT0p9uSbePN
4y5cLVtdfewfKFDXHlKty2E6Z+p67Mrbt0nKcQr5D7DkcUkxYvDhi3z7JA6nqXAv
wtAr9228OMso6rcmtlHDQo1+fy2/P0PTTHyGG9BD+ALEzdJrfJdHFnYiWjdHJW6t
18kKxNJUOtmAqKW1Sk8sE0cB5s4jse5bLKWXAl9RrQor/UCUcS++rp1ogUp7rYcY
tA6DWd3nfae/vnuaSN8lys0suFkqNu8HO8Kt2Ch/3javFynMr9wEHFvnBQLVNXuo
TX+EwqZyVpvTuaNQ+4WVNTkWBxm9pPJwdpo6+NtoZTBHOVGd+z9GRVP4LJkCuNv1
4EE+8FEyEu2cP08qebEIn4wL4MMn40hfMCwxj3bbar76DoyaZhhIj6FZsNJvxVcq
uOYRscxUpOXBFMkj5BQYoQ6VBlK+K7AWJnHKZlDcbOllUQ868hYPmrd2NHoaNCF+
BWHQMdLkLQscN0bpMDPN3laDZaIxrjsUGbCJoldp7R3cz822NkOholA2z7I3UUCR
NCEPiH6gbmPC4Kypd838VM5kxF94ReZCiLqZayslreHMAAHENFvKpKabdQfzK73W
8I254/ZRPZkVqUH95zwQ63ko++jfOR4ojCyEzaX3vJKVcgcKsSxVjyzNRB7s4ruj
3odPNyr3nLjgETV65W4pW7X1BEeu2TCmmGHTsfkD1CBA1E9P0ypwXkztoE/2Lyfn
AZ9APETYWI3EINzo7sGXZRQSaQ4cM17AKrV97uHWRhTaRX2pLCxpj3Q6i2nJ4Fj1
678s952atVfZXGbkJmCEio9Y1+QGvK+k2ZWM9lW0/89ffbK8Sq37frKPqRKbtLLm
6j63PgjyqGwyRt5zfzOjDQaNj5rd6lCH43WVYvjQ28IPYPk9Zt9WQhiV4iepOxHo
8RsXEZkHpOF/RWIgeggtu6IqOoqBHLdjK5/TZsEPs8DdZniL8AtXwePoADjH2uXP
ULHmSRw8rQfRq5giKasYAFEju8IZg6At4mX3HH5rraf8+Ow6lCkgh3AVROp59JKD
1sA0yJs4upn8S76qNWaBUIu4p9Zz0SfQ6PDvlcMx/Bes1w/BQVtgGRQvALt39hCE
CNTk4TakR/g99fyUahWSqjtZzuJ4jvAH/Q7O6A4JC3jU+lHMyv5CEWLvBgGXMD81
5/8wAg9Z7bOcaRmdU4n57mlmzWY8D5qHWwae+EWICJTv1bL3JHC/nBhSJpWo/BdV
p9ovxJr6NoHprADOx6vG21Zk9II/7HEveBMmUWhXhGa99rFefRSO3N+CB3pKM1Gi
FVbmcZgHyt2ulzlrvm1bBIVSJjVbiQX6H1NgOeQbVpUidBvC5/t7Mxaacui24ZEC
BD7U74zJUNw4d3Um2qFD92iyur3Tao/1HEP4sbWnm5ZGI/noTwTw7t5356/O0dDE
VyLuNX9smH2V25nK30rfC4CLyffGG+o0kNgoVWCABIIZV4qN3oswToeOdjA4lB2Q
nktG4PpkFc+eFKWbRCM43T7mQLnpnbww7vzbMIPCxpsNJjqpmQMNwa6F472aTlph
x2WBRLndomPjkL5/5fbFW+BDlo5fh1e4OHVBFBg7oklwe+xIWVj93P7P3NOspDF2
vyt/VZ/W4KKgOT9NKHFhdGpKzHNhsTLe1DgCpYS7AZyNO38KM7pn3f0yxpfS6x1Q
YF5HPwir8/7TshJG1K21JDBgrDd48IjqpWi3sQKpL8RdFVOL4K2x9mJrHE/4b05P
g+6jP1i0d4+izcJazv4z2kNzMu21bisHxGzQlDH91raeYbqvSqlHVRXiNm9sncvN
943EfNdlQ31ytsnhV1Ge3b1sGYkg3Dw6fOr2gKbcyAiOOOkMG/QuYhk/qq+IjsEq
G/MsKnKK+PUz1cXJGhPFTFPcDqNs6l8jLWa0Uy/stL+0B+3maGv5nAviqA93bcFh
oucWlwbGZe+QpSm+bjx0em/suqIPo6IYlFWoNsPHjIa2roR53Ouvokr/rSKDAgWY
UDi2mqVo84d3V9cBKxC8X+KDmnAKzcvi5ghjJCCbMIgv5KZADMuH5/biKgzi8Lhy
4FkIhp5AaaHoSi+MEImmaz9Jk/OjsIdpQPDyjp2h8A9jeUbURvLY5AP4HOq1phR4
7X8w4BUkjb56BdkRYdekhOarT//loR3QGuxdINIVLxbKD1bwvQFOK8Nkh3qYITBP
GOWzmL8GImg7aQ46zw6bOCpOn/kushTF+1bjvDVXLXHopLppQIotYDKw1pNeC96a
Lz3NxQ1hHW5I5ivBMkJko8IrI2qjMBFTf0HqrKZr6cv5AZbYb5uEi43fL7HJ0G9X
EzKbTHX+UOpUNn0i/SoGFqbIgBhDPeI4iTC3TJnWI3T0ebAUbrJEskl+Ht0hVjIj
Mkv7KOvVAK9G5O10puzcty5b95gK2P7ncKbo/oTpYkTfQe6h5OXc+FP/qLE1l8G5
h9HumrdE+wuS3TNPxGSwZZvOHXFdAEjZRJG0K/55vPtStumCZNqMp5IdBoPt86Ol
S2VBugeLj5ll/fzJzl9kOskBbErpw0d7UcKoahT+z8U0U1YrX7OOFipEYsG/QgKb
FwPDivYQFZlNXqE65AJtEmFiI2m2eEGL4unPiu6AwaBqNm+J6UNYclJCX6PrEW1Z
o7s7KzImgvhgxwYjZhNzBxepgf+JjuNIBz/8dU/WuXJijDiuAEWqbRmHMD3gSTuR
3RqYkj88iIejX9zxlhGDFQ51SmvYqrJzukZn8pucTnevHeR9HB+V68wZ5Fura2xi
5cYlE1zGx8hFFSnsLyhH+e7KaAV5K1psCEQQs6Uq5vB+Ka1eRM8zoFo5VjWQYFig
D794iXZUSq79N3tGpxqdMxW7ZkUHMlxim39Zq8nu1uAeSuIuR4RGLwBEUaTI3aht
QWf10xZvoJ4B2GdyTw2bFTWqtY/sjohgMdRBIpeh0oRcrfqevvf36jen+TOlK+oK
OjP+Zj1wCaHMclaOGCbg8urzrD46X7QoS+GzptbQEQ/yyD0PvThTxogPyDKQ0J2g
lBuRQcjQWIRKkFx0F5WcvBfmxOD5TlJsfAflq+1n6kGsNAco8G6YcDU41EnuX5f1
1MVAlViAjwJIECISDeX+GXMgOzoXiWIwgswgNtR1sBsAJ5dWWsyJRmCafpxUpFwq
gxbJD/tPdkv57A6hEKWmfxqM2o66LKeODZjyiil8++zHmnJt+707DJ9carxbexlc
LenOIvkQgO2QaQMOCAdpBGxVoYgxH1NFNRLFozoSFqtbzy16KiGw89/+eUJUtHqN
zx9ZP1+H3Av48OF/r6u/cTjqSG7ezMDrd3A4rx6L6NoDw6th2NaENTx0grjtmmwT
mVETYbbzqPHKj2OHnF36hNvx195yA3CS87/GpdjjaPrm4fKbR/oVmsxenElQw2L7
UQOcyAovBi2O9Nk1YgAAqfFMTLdxyVkQLxAyAD8ncjla8UwSlcuJABR7bb6aCwH1
2EqC7F0oNy0pHD04NJCVyTm+3wvXO0uiyRtqlidM3LmlpBohjPZQxFVfB8hzHhCN
TF40eC6+JPWOhlyfz4RHJDFY2U2MeRsN4Xsp+cwxHfeMbhq+JNQbifFCuqp4FC9a
i9jOAir5JLV2QxzRkE6r94GHVo16NwPB6eItDG1f/mmQysLcHsN5VeE4SnD80j79
VnwPAvI+CRRJMCI6oG+UY98FVyto1E77ev7TLT3uwFWtt41mp1d9oHWffueihNA0
VGWivmt4iEJHX6rY26Bryve03R+Fc39eE0Ynjn3Ao286ntAM9Stbqe9gVqm7EvPA
BYWEMOEyYXWr9OBXU/xQxqLi+gT23EP3Nlzwj/IU9zQMiSUcaHbxGcX4OgxV7jKl
cR7xrk1pMc1CdCUaji7K+O0oSxLxRJshQ4jE+ZixYBeAPBZxdI61KmrBnWIG1LIq
fGh6yoEew8a9F7vX5WnVy7bbdznzvlovDZ5LhcM6YmdwwpBXnpvjSRHRMNwJ6z3E
G+uKVSrRWFx94JuJm/AECk60LUIGEmAftK8Q68tCGh5JSJNlYSYYGSMuOFXf7V9s
PXTlqjDMFxTK99Vbmti9JF5V38OcioJpRaheqqwCzFlYREwQmb4bvV6MTKFCZTuN
/oA0U/N+DNuPBfl5CeUqwAPehZb28hJYEibnZCaXpnQTZmdSWChB4awpCbTWhQyQ
79s7QH5ujYfCHDFBI92WbSPNigH3o8JwpejV4s1GZ4lpVk3w3Ww2b+aOrQMqG5ko
h/2QNDPw6RdfP3w8AFYYE4mpsTz+7/FnZ0lDKGD0DCm4P57AJEuSUCZQCHrkZNI9
WY9rJIr6Abymi1Uf1UUkEa22ZjD4S2q/UU9ITm7GxL7V81YrJxAenYRZvDarHuSk
teOWkJBxUILYFyyXq4co4dBguD8NbcC6H5hwvTfl4JnfJvEpx4bU1FVO+Faxg1Hf
he7W4I91CSpoYC+6IBfxu0PRT1MCiS6TYXIcAJrikNEDL2KBmq9i/DN63EA3zc4D
UJ+OeIO9g6m5R9XteefLa+3tKqH03DAR+80eJN4EnAmH3fA8eQ8MW58MEPgQ9BDe
+y7Rdrnov2XEk4+na4c5EAu/QlAVF5JEGtwACPQxcN+Vl68LTByZZE36J7Ly+8bb
80uPXDifYTjxffMcWSCVz1TykkVGB83dTyaSnfye45+r08KhFEvLlmtaTb+hY2lc
FkLLoNmhl4Cokvl4WiiA18bpfFbfsa1Yc9VW5On+HCNiPma41hxxsAK7gZlxoQzw
XFwbrkURdP4nX+WyjdPceXxi7N1t4Vx2yNABBvw07dU6OfwyxSOpY2AW6Jo9Lt1D
sbpO4JN7Aglh56dL6uiat8C90anYD0J2BbeZ/lBV1nNwi2UxboJJTddBfwrADjXj
lscPfecrzyse/ydRBGVO5h6MRNiQBWUDVdD2t75eimdC0Gu3GJfZfC4cg2mYXFo5
NVG1TgGhMSAu5lrMyXiXlhkb59jAZ6wnLbpqADGyUt18VgbB2QH/8ipxUUjsA0Nq
SXrcDXGUUM1mszdIO7GwpZqra9TKHnf+n/WQDCc6Nen/Eu4Tvb2NTNDYnaIsJ8QH
y9ZSYK90FGfNykgARYYXGwRQeWN5zH92W1bxugHHI4ZF2Of/sMIeq7u8zW3iep4v
23tkVp9KVObKTXleFmPUlb6/hjXIP+K9SkBaAZ88QP1sydoMwrPKxfVV8h7nl/wa
g62kkubKjRCAZsu8K1mOdR/egzTgqFgfUjqBOrsqFCgAPSfD3aDVRXArnu76146o
NZaErrVBQUp4OLOc8jmFbO9/uJ+uliVCUtmqdFqg5DwPqQf9RDg3OLLlOaAM4w/7
hbE9Y2rcVheq39H+bqKdgFOnIdOEYh8PaOMxighsFkQszUa1yh+u00XDCdrzBtaN
PI2PyfcRH4xWBO2QCY7liAMAN/rSpig1KKjBlDbjbse6jssqLZj9I4BL02mb8AGT
AdosnE0YCxqg1+AZT+v9ogkTmoCLDiB3o4lSToQ2yiKS3t2voeY5HaQAisBZUlVn
GqGlGSKkoagpSCZ1UCQXoU2E8IgxAfUeMRYuPI++45MDflUoDxrB7JgIk6TjadJP
aP9F7qbDLyPKgF14bu6vYylDPP07/bNIM8TxJLB/39fuYjCShqSdO8AhiO/1jJJL
g7vguz1hGBwIho8Ha67aH5CDb1PC4ZUWn687YPpUop7cZFuAJYPpBQaxIYuzcpbM
Bcn3cVY9wG+9Rsk+9wMB7G5qNEu4FueUSYA12BlQCjkvU/NEqUTMCwaXJTPAhQgE
y5jJ+Mqs6R1CCdx7gUKvg+kJ9znvdnh9Uzfpgww4WAh3EBqFQ1D2ZCFPa01Qy6D/
SFziM7oEz7zRbHwvYEk6x7iAoGfOUAMRtA59pTqaad0ZoqzHr3ZHgTndcHoITEdr
DLRoi9UbE7/tm46tCP+csdpnucL+wuY2wohOkWKxa1TTBDAtuULxQDXzBpHLuCdY
cY0pC9oB0BQ/BOzzCNWnQNWB+pRaBzz2NyM+IeeQEgys2vPXqkKsFXVMlZC4SXpj
u7iy68sjAOafo4B9QkNPeRfCELIEcIuQdfY8ghqJfIkDBGMcOLIO+kUswzhsQBky
gT/+AQ6ryZGbdle9oNk3V5QA7Hy3ISpboGBw9liHh95jS6WXiCbRcGKCfG5lu8Vw
ttDNmILCWo0UnE0Na1EaxGPrsp7qqaMZ/6joZs/Crm0EyaYoWG335D7SIerVql/D
4AIOQZnNvVTWOA2rGDj3xmLFVF8mi4D0lnYOEmPPVUMsB4DkmTwvG+8PduoscJlI
w8b/mE05x4oljExh12938WcSvA4TqDAoEH5YXeloQd5gsiPEv1giJlDUvnSTQbv8
nfjxYCdhvxx4TpUeFWcWf8xQ9XmOj5M1JIF/sOX6HyMIicbK/eCfP7rujOC0Imh+
TogKjcdNk6X0sdbWTzJD7KLKFo7GPv3uLrhgIaNd11lohSgxLolqbT7dwq/IrIry
9aR+OFpvA0CkgoS4wKJthpzmEotXPJHjwZXu37ZagX0ujn+kBzqW8G0lINor3qXy
ZzSUZ550ALAulcilXC3Su8QktTA//JwJZPoBlWRMj3za8WO8TZaVTvOCEhLShCk1
sQlLkGzs6J3RQTLbzovrDnYf4RZsE0Der0vPc3HDfn/ILDLqPDJfHIK04vlyePE0
2Tk89a5qhLqhLBPHbGttNGNgnSuQVEVaYStRvvuvs4IKdwa9Pj3SisI8xeZ2WbWM
hF+p2yUW4NIG/VbNGJ5dhxaw7DOd1hz7ZRETGataaP+QRa/q5j6/d5Z2IBO0gNBN
zOCHkIzFtfDfyfpfWAH+9kKfFjHePV/4pt8spnqNsiZ9S9ncjDMY6WolmydUjk6D
imzMFyNo6vroi9oVQZNnMhDO8IX10jqRezEvY7xC8X6U0kbnZzyCvwRL2Hfsa//4
U1ZVCekabPGHKHxrgv47flxlfKWuYdhMT6y4gkhJTDaRMmquganpUrouZhljRb+M
93RPugBan90/eNX1t/CT82TNW5YRtNc/cPB9HGUCChDa6cX5DKRP/FKBipzImI6O
M9FKhz20gNeWHLw+Xw5Wjl2A9N1g3JmeE6zQFr8piMGLpwgbIoNROjpDxrvozLPc
Cwvi0LKC3fnDUJHB6+d2fvvYsw8b8bCbmV7pruY30DKbMFdz5WUk718/TXz9iAu/
4ByhkdXyIHWf03r+OTVL24/8LnmYLbzNYKXFQS/X/4YrcEXKGRgtSZHxGU0Vj9F9
nS4rEFFV0yfUzIt2zCzJeRa4IDeXAg1H6WxWlYIPvy7d4pBVuuzOb6nA5pXw8EzY
gvqvz4Z5wW5Dr3w7gZ5DXPd9cysnXHtX7yKZVQwUzm90fov0RnRF8Uj+ZHwBIIO6
exyIfdgvH/Utk+sDwOfl0m7e3RxtEmaY9cqKTpEux7jVNRkSRNBfFHA1VxFnvh0T
7BoD4b9VOgNaUeKiSjEnY/rWZZfJhTp0L6ioCAHVuabkjPVcLCuDrdceCFJDlP4X
ylrJaQrQ3cOn4hO+y0o16Mslv3JAn1HK9S8QWJ0LrklJircOPLUBXkpEwAvE4jp7
LenO0XiZjI/OWl2HGqm1W3Gpl6KKHzzVacxnEZ/8/lmlQZK8KaqRr3egQ33ICx8M
Up8W4lUWcGuWxmHIYjunooEWGXXjITtki0w3hEBeK9ORvbcIF3phg+B+0g9veh6S
yeYms+cHhs/+O21rd0zJfDXgoaBtmX1y0eI2/Udkpzsq2SecQMothKDoDMm5PPBb
qL+wV/z6i2HjwBwAvIuC08IlyJHMU3Vj3h7yZJTJ0WO9GkHbagkWCJ4e3yPr+Ksm
ad8hTCmn1bZp+FfLgkg6YjkmQt5BWLDlufk+1IhSqh18QnRNjjtdgoQ3PRoQj+zn
zRx5egNyPZPS/l+Jqty2b/KjYUMjzblWGVJBsOj9kOfZMKr7cZDr73wHjlmvBEby
RPDI7/20MR7cxK1qtL2RJrxoQlrBgO/4Y/emNcbecVe5wMRh4h9d8XUJV81ldg62
lRUAsPaiaia4NVr7FHWcbuyp56BwvX5cD5dsYlDELQit4c0xUJP8rWiy8IezeRIX
49t/23sGMK0NahA19mw5eddgsYCSoTXeH530+poYdYgNagw1ukaHk62e+rQPL1xE
K11C4EYhjBempQxdqVDbdgh8lOvjw63OR1msbd1VSBx3IzVowbEqp8qlLjqvzpZd
ekVDCauvvUnDq8J2VZ7rmKOOBTpZ6ZqMUBFEi4rk+6+MfE/jWMDDoivtLscBkwpO
sTP8d6TwN3qT2Qx29fI601Zo2SyovehMpjtHpCpI1BY08eYua2H/ZCZkBIJnbfLh
lNDXFIkS8xUUyt2HYttDDKy8cd3LnU9AwQ8l63HXKZr+TLYf0bOuuUPy+xh3HuPj
cMRatu9QTVcu1uwdxnDZTLXI1sAjt5ZFrii7+buYBVzZ27MTmUi7E9spY4pIVmZH
YVTBqt6VIq7spxuHAa4Ks+C5EgwlNgyltqOFCyuZJi7qFVF2ZCz0Dqn3lC/N/x+t
SRFx2a2RveOoDppgkH/EeXhOBlZNWOP23F0gUfdy1uD+yQma9FJ1bWaZG3bX5qpz
trU4vIWPOxmWkkJnZSYt2b/Do5SUVFTu0oRiAq+htjg8e9rA/s/POhoRyUF+a7ik
FMgxNhTeWfwh/tsFUvrseSO2IfT6fPEz0pYno5tldGUseXR9W7vHGr75/kfh5h1S
6jphr0k9p29KzqL4C/C/jKCnb+ZFzB8+dqCROQXflWQgGzikgGk2yuApCQseMb9y
wQPoL2DRSwlqL9caNzJjo2cDWr9AhqN2/J1wcNFPf4T0bzrT1WnRHUnOhQht1JNr
uBhCSvrLmfK9T4QXk9f24ntrL70qRej6bt9YxtM+IjeV8rcXBZNAmSrVgHT/W9WL
GbzmvHiRuxYU2pq6oU8jTwoXT/tonmctm3FxxztTtzxydho3o30dUcZ1WBgMZuHo
tK8JEV0coEhk+qbIQrdVQnZHp0p/LqcWZqwB3Nh9dBmkPhgtFSn2pVqTIswbRgeo
Ot7DqPkhLpj7xSZHxqs/5lWLqHhNj25hFllYTvG5zBGuIRo8ikgqj1dSqBzA3k19
AfRQh/aOx1SEeptNBjvBKeryboyT4cEcpVkyBOBzt3GWbQz9hQt1LJWg8+wunPsp
p+EV/Oz2kw3eQKMLSZTPlgY7yh8vJ3ZQfxbBNxODsSpHmTfmVv1B+FEsv7INd0OS
ORk99xS6loaa8DjlJ8kvbjENSbOuCnlhokGLEurrBlAzUrACt69UkFpaJET98BXF
izXdQkSP9XZN281LViIGxl1GWleooLlbnyAZYJRl7UNdDenvkr5YjkCRm5KCIr2h
1E8iKsTHbf1hlVbWLKY4nCBwOCdAVOkm8kDFaAh1IbHiCEwYr5ryUpLux2azdF1j
JJ6UBiCxGpsAnpyOB4/iGVz+JhLjqrzgziOErF9EqfVBk9HBc/YVW9l0MxMP7vp6
GFuKTwI26abbWfLK2nrsE6AxSsRF9410NqO+tVLKOXbzyTCTS/QTDBfol03Du0J3
yJRP0GnuYK8DxPR+iKUU50GJQvlVGZmdfGOvbBmGz3/Lzo7+XQ90IfPb1UJFKlbw
/EbGbNR5NbxEPMBNK7iuK65ZyX0wBRU8hjRYTe/4bek61+5zGN1exmTc485Y/Aih
m0rVjITaB0s9zSLLe9+iwVRgY2GiDPDMuTGaEAYOhw4z3elUPWqSZK8Hs9gyZWMk
U0YryQf8jW9SHWjKtSOhJ0pYdqP8D58uS8UIyHkbwN+l6pXrYvPfXjYvBnLTsnvu
wALBNGlrGjaoo6JOEq59u0tr+8ShpAdeDsK69Pxk5J1lHrt8Rqj7y/3hN25R0Jh2
zOq4PEY1SSYV0dWP2+c6pM2FyRMswNZvMfJLlPVDWS+zWSxFpicUG+nksJJ7afzR
IZzcm7lbESHT6uWCy854k/xgpChDqvERWIpuSjvZfHTvpa+8WL2tuQaD+KVwgiKd
Cmcin1v1jNQ4f/XMmlo2BfBr+BoEQXoK1SFMsHclstRc9rcVZlDvCk15kkGLuD8k
ootGOaDSGIrt7/FyeiCWkO5X03/FiphkgQ/p53D+McpRa9fF4jNOkd2n5IRPULfW
8j3NHt44v1zFuZm1cqNw/XRDk/33N6Oiv8nEbWtVSb3nZb2rJ2jCQF7hHDZ3P9BX
Pf/CcrDORgm9a79fewOC4yhbmiYr5EzJlw+7ItxXfZHyljUNs8v8Rbt7T/LXDsw0
YXGRRj7nzbsHM+6RNIqpem/0TXuKvNJnT1lzB4AiFfmPEvj8Xm2/1kiu/HVK0k2E
RGiW3fmcvzbMZ2UIbbfxEFDIXP4U74lJH2YVyDpfPpaNAk8U7V7Vy8BKavyJOKS4
MBMED2zAghzscupHfEjeo609Fvj7Un/iXrLAXbBIOVqOqUvhkMWdLB7GSM+Oljhx
NFn6HIykwPdUX8VwtGFcslEFnpzfDkW9rY68fDtLOvq96nma60Efy7TPaSF25kZZ
LXeeetkN3q8FVVoMYbGyIaxgvTZMCBm0uyNg0c/4Qzx6x2u85LNL3llQfgFEq0au
YyTITj1llfFuRhkx5cgf6JdpYSRnItko7s8xgqSdkK3ux6lWxcipCRkT9haq3rfb
ccKC2Z7DdCXtbPyB4k+n+5VwT8M7tleG5s42bNGWFgGT/RXPQJwxRuUb9dDnrNmV
lGlo/YNrDFWEHiXsWqFxpNX7Mykmv/KIIUPrAT2UHorHQcCJqww6OUCgq/gvNxWP
GV0QHR0dy3N2ErjOS1tQWPSXqmnrYJFBOjVLhx9hp2clHObpQS6I00RNt9eh1DQW
o4WDHOrCzS4GAcgRt4/rvemhayrqNBFp5+8Jx4hTYFOCWWVjIeq5YHDqNGp5pBFv
U5atHdXvEqTrRmg7h9Lm82MrYlvSqVRmkFyJIM0QXElF8d3CqDmIlgrVk991hyJC
wP6mSQLvFTLvoxWiTul9WC/ot8TNGa+CmGpVkmXiAzw2BvmrKLJefS+3BnXUuuTT
L+0J3jkT9e8aN3d/V5jPtsZ/8rwqzmO3M1h2+vZVLKIaxpsqFNDhBI+fBfqlF9SK
E1oAfUQ9nmbLrr8GLZlyC6+eIrt09cpju2yMou4abd/O01u2XM+JvwRtMShKpi7e
r85Fu72ZJOke0JTLuvedpe2W1wn45DBChlxGqtOtKNvToFm6PyRi+paJQ62/qOK0
eXJaTF/bGrYS04ckVXmvA8aCUBxld1lQjy3PZdRuNLvsFEaIRdGlHqyeUJpIvZ8Y
dwz+/5bRMsdxBaz2GZatx591x1YovCXvWXmqWIYAIHiPabWh1/HpIpM9U4axMb8a
tmAUy08AAF5M2kYbqMdwQMBEoHwgRnyXffes3rvsI39VZpLtAVPc86bKEpSiRRsi
QrIJ/jQkS2NDQWbwtGW+xyv924Vzyeur8WlNmqaSCpILxHSAc1uUmywOTop53IcQ
tcnNDfcKhGZhUiFJj+g6Vjb8uEE7U3TwXkwkv3Bnbu+UxSVz3AzOKVi8cE6ZS9EM
WoL6syGFzIhxD1tGHjf84Hb/5GcdpofmcCp395Mc49AssLkc8aLvzAxm+I6s/itg
vbWmajoIMpcmVc2QA6EBglBUYwOVrTuCLevPMwSg5G2oq9T3Zi1JSEvFzsKhU0yr
xSeg0kPc+eryXRd12YOH6AkbJ2bwPNv/FzovY4xlpzjHGaLLRGGNe6L+Vc3PgSw6
W7polnkxA3Xg6G8LUCjbA8WzSGiHMAbTDDylXt88HcPX+c/B9MWJHJOJMTVcEO5y
JmfoDSj7VRHQjF7r4fuCGahM6TwJm+AMUfjRqXVDTkomdvVWnswOKRpijsj7BkVQ
d/uvtM/vK/T4cLXvCaXvYjhKqN6qd4a6846iVO8Q0zA5rGj3AMPRwB5YrAjONNgX
nYd3w3zy65StGEywYgCOfmQP8EvQWgrE8kMZLbh22XA/hkBX3bnVD+UOIT3xrdOr
LznCRFD7YifYk0WUMrB6dZn+zaYekZ9eNqopcFGwDt6S2G07Le1ahDSFWiCiWtWJ
e0QktJLOrYNnkHCi+1v4WqQniGuqdL7RdOsDtEMh7TOkWNptwNwx0y3semoTbDSa
ObZLzLGfCKv9sj5blq/l/3ZRye5BoRWsc7en7EvcocTKeOo8LM6U8n26qbYj+SYE
VHdeJd/IQ/TCx3Hb+ms67E6pTUGDcQEzsIzOhYwLiXoHc27OHf3q0JFjvXe2GCN1
WGMbt58jL69eg+IRBdlGwXuYCB2klO9uQhgueaASzuczkQRm2srPzHhzvHtXoaQN
iSvdgo+IZUn5Cw7z1yg4SQ1I1Z8yVeGLhjSrJW8woli+qnMSKrdgE+yYPYYwb74m
uyNB0j302Jaf3WAVbSJUn+xY/hAxpZ7Sbe2j2grQ2JJxJWZXnFNIpDaig/yLetMu
hLNdyAePowlCisTV0qYI/WNy/E/m0wreo+jyPeSgysVrGc9Mw1I7rucvFi3K+0st
WrMLmh0/ZzvoPfx8H/fy2S97zicoN4w4hbTpcAA9Ev/VlreKBUpP4zhRGg2cEM94
DjkrJ9jB2fy/bmFxGMd6T/8pfKVtz+W03jkAt8AHNp4TzWw8V1pMmXu/sQnsy7X9
qw04jMVha4FvixBPhU19d5prUhoKAhNQIvcz84hJavRExRosBXg5Nuo+zu9aM8KB
yIog/5mDoDKjbsuZd2m8ToFwsce11kHSvJ+4zi2Cs/7DxTwDXdMjJjXh+/ZRvvWp
4r1JI5RWCldAoLQM4T2n2GBLbBuPjTocwIjlvbRJN1ypSekDGqc52GzMeatX5E/9
BlYmresZ03tQjq6t2NzE26WlqpFJXa5BKfRRSSTcPb2vVUMgtRMiViyjCCYUDWRq
eTIWq3jLg+dyTRaBgVC+DHSpzdzKYDvAZt/zY5xjEBBpYlomm2vz8K9I2PuJqzTl
Xz9/DcCyL9vRlGvWmKln55KPzsAUPHJxuCvy+SZGJLTzz8Dl+bojOZWGy5ux0ck0
pRHhRZjnWKkmuulFreCffMbZqnq7EleXMEiPcmUmurj0jq+YmxIPai/dGkB2z2O5
TwEMgAWchsHff8wHKt9ZdIB6/1+0MaH+L+TjuAyh4RJ5vwKFdzRovOQFSh53nhLs
RpACtErwXOUsVd/psbjFMJC6NeZJZKMLYfqgfaLr/8yW3IYFTK8+reZCmfUWpChW
FQNb+fEcBZDHvHUxtyk5pi0QYTc9wnj5iZQTWsUpbPTzjW2+FhitOjLVCtfEdBd2
eLssZZoJ+NGpAmT7Ol13wKWgTbQtnRUUxUQKgOhTp93gWLj8Xvs8qSyf6h4E1+z4
t+w6OD4R+/pCjrtJnwFGBlxD06OHL6BgTgEVd2Wj3UsHJgM/EKKS8bRpbTrfvH4G
uJhHQA5IImLz+iLhSiZdvxhgLmBUlm4wLEK21Bu4dn6wH6UYqGiRgZCYB5WCT3J1
Wily7P7wqMv3OZ0bFu6MfssTVQBlisBlgLiRaPvQdIa+FrGrWt0nKxd+5eXRZqXV
UjrZtWkrHGYgAZSInPbfO2g4v5EF4aYlsh9vMK7rjFB9X8SOkqRsaRmLU1NtDa5o
SbrsW2TVgm1eaudjU5VInp7T4QAeKg/CCWJpcTj6fWjteEJWxtcESCc6tkQyVp6y
YTCFIi7cpdlRpf+AM2oxMIGMiysqhEi0yikYQA0HRYCHPc5qY2pRy8fLZFRID3LJ
Fu68sr3JYLy5V38R9+LRuznioTHP1L0IwrgwkCxrmblP1xHbzMtnXAZSmCBM7TmR
38xZKN1MmjOS6tGcV4/70su0Q6ROwbCNKN8VaCHdQmkCvrq1AYgy/0zt4jNjgu1H
/4r96nGYOe0tLYu+TXCOq90fZTubcwozmQjiNZJm0T56To74wXmvHkS0mJjtE4Yg
k+zMIIaaRWusJQ3iXVQJ/70DtoR+BaGX7Sa6HIYQtZL+1yoeyPvPxdGyJRswVoK/
L9+Q09hcWccAKNCwy4sA/GIOHeOEDiBvbJcT4VEtIodyl1kPobzuHLxuHacMaEda
w/hFJJmP4gZZ8K6tBBun1ydmcTqA0sO562cDJ+9MIuXXXl9TV0r//rf5bmvlxRoX
2pnORGyoC+e1WEttiyXBwo7H4OC1++1xpei3sYfSuRCxfagpWEjC5WJp+OS0ijUO
o+kCB/INiKZGTPiL4wOKn9Fh/EGDX6eIdg1LAasnG79iTSR17WCcfxO0Pieg6fmD
uzCWh7REFMlDNtDGaX1hldvykN3zgaqj9nSD3UJC3pkaEbwTTMjnKt+2xm7aG9Fe
0JuZDdlBm8s/nLzBQ4qIWpSscp8jqYX+wyzKb9nZvX9duCI22PS4az8+u7WlR95j
vnslKVte/5X2uGFDXAxmTqx/l/w8xdQV+4LLIlh0/gN+LkpjvJ508tKdTju69PGc
cqXOazmPkhx7Q3lb04baDguYUBpoRunZxq6okWgI+5tgaB+4edhWl0ytNdQhPadr
0x7IxcwfdCbPnMwdGd01Eko+ZovzS39O85M/ub0/+88FjPVEz5QMtIJxT5Ube2un
p1uVTx9Df1rBzBEw1oO1GREFa+k5rbplJBvuVj78d5wdfattAI4C5090bN6q0yNl
4nbarqSx5U9TS0FngzlTmm5F8kmz1E8q8oaZDKkZILUdBFzSyHRS/ZYJiClOTtmP
smU3OEWsnkEY/AV2vpGReANU3XyYhhSoGmBvI5JmAaIps3veO8cmpeEVIDjzPthW
139cp1PpFsnPGX+NZeIRhUEDjPX0oR+aJj4R2LQ7YojnxhXQeA+zAmIDY7B/WsZx
z2dq9O+mjSILjRrdIfXE9iUQouLl8sslKlsIl1RsvQYac+PnopqAbu2UUFxCUmfC
LVh7LskaawbtjpEq7MhOSlkEVFzxjf0s9rGE6f/0/v+uAm8Z4GsWJmDc5Bde4wS6
FGe81c6EZjt6s13FvHorhtW1MIx92N+jn59bkpZrg5qi3d6CdNkTBMoLJPe60eEN
991kQ9L5WPjHq2PERMrydgnTUI/YreUH11jdMqFYwfVw0baZhKOQXDlkfDssSIQL
nFyfbYH/ILh+eQHhCsSyM4XFOsT1LQWLOyiKDF/29NCio7sb+lRu+i0L6In/loO1
MkEumnytgPW06GNvYA7PTNCxmfxnjvYEojNExukSsUYEHEQBpQ1Er9VHWP9OjHT+
hhAW8/+pkj0AGjEu6qdQ8MPm41kY0JNHqCMS4WMg3a7H4RMIk95bwHpLxMUK9LlG
uSG3XP1RlsWi3Fs2bUabqv7fvz6ztBAbDI7yd17X413c0+ShqozyGpuNbwIrHCBv
muH2Bl/LICgrnKcqfZ5KmodQauC1h/tVNpi0c77aH+++EZ87PCs3G6tGyEeCY9iY
m8H+PYKRaDYArqbp2rJpbwYiWGqS8/22DmVFu3ntUAj6aUNYDQfSf54zSnGt27WZ
wDVHRkhtMZpftHRw+XIWxSid8G3qf2aSXwDYEZHCK3Zz89RpY6LcYggDDJrg4JRV
1fazK1UWeGkuOpKTBYzBduLgs87arEZhpljLdtqUo2eg67iqIfq6soONWR/BY7d1
JfToK3iq6rcgK9ENqobGSPJMhv55Tss58qkF2+lGWOTkxxaowwfSWNvDBMNdHabX
PqWmklcTg4AEOe5fZQ6LoPcIrgMlAxTWTtokhQ6EcjHSkdVyQvAYiOcxiFgex8O0
Zpb+tpvinvTm6ssNKQuMv0MVYk+3BmCsJCOKpVpzXJaDFE6MWHD3XPEx0g/VD46f
S4MWn1ZNl2DJguOQ/P3PcQo/iyxKlo16Vj3ildFjiZlQDkMPqsLs9IhDjdQAtg/S
qmwrTYN6K+X5Na6jgTSp0LlN2IWcZ+XT1lV1/A3GVOpHwnEmtKn+rquF5t0X3Yzr
5tqEHo4QdpQZQXmyVViArmmWAj5LJvi0Lcbm/vRehmovqO8X/b4OIY8NPrD9WmpV
FJ/gjSeA+XiPFgwQZB91PGN/y2hfwqUnrREHfUHWWGyLpRD8cKf9iJFc+5xirKsm
gWhEv/bo7sBsurIO8my5gRguW324foh1SSqOFuOCO34xe2Jk+5jdcDCAW2G7rS4Y
3IElTiGHMnT+CErJEI4VhJ5WGxf960H7WON7jtepGutsRVQmzl2okMHzuyEW2q2p
wPwBVliWwgO8EDF3VbDD2CT0h4b3LZ8MN0Fd7SjU+sACWggGoobfgoVZ9J6amZ2f
kWlrjAhyYcbgaGfsbUNY1fB1p7JTM33LTz6Zk8r3Uu1OBOuvJELJK/XdtVQNVYPf
RRVBTpEEistuDT1Z1FaSZTDgDTTtz95N2HVTsde0Dk6GWbfMm63nibIznQCVdAAK
l//dG8N0zfu+rEgyAPrkDnRYKrED2fDyLCdWq6b05osCDVk+8b6gn0a/jMqguxZW
lf6wFLKEaZP9+qfsKyNWRAh+/7rfKQISuG3H3ZvX0YgigS88DCT9SILhCy8OnF2x
WJ0ebVc7dTfK+ZcH3P+vRfGv324IaXhZ3uHZfFW2rEQklcDeCNvyHkfUzNEvp/ml
2bnsicxVtTGWoORJ1q1qL3izcn+x/b/k1teQkdJDHfYHgTv6Kfc+LFsC6WpanQsE
QZTv3jRHBKqCtJsNFXPX/eQPZJBEr//hixTHEa9gnRFWw0+65x0Zlh2axQbE8J2f
9wZg2QNsIy3YX4m/xOsTZHWHr0aBPzA31U2mmvxeIavqZPGHDuaH2cRWjZ4BqejG
560Lm7oFZ6En+6dcP9JglVxL6DXg2sIqM4YIt2LEMjwADhnVwz8sMN/DZSrOBibo
lHcszVdAar13cLN8S0Ipqbs7s0l5qtebtutR44cbj6aw2TAk0Lg80z4fixAIUXmu
ifqhu0HwRzt/omcS255OfDJLC2TZNEodCgLEkqwINp6CwoVX4Cmk0O/fzsJo99La
EUtJypuyC0n0+FJh0RMHV/ekVWrkbGVA82ZB6KdFTE+MM5InwvDAiGF2Bns+QFZK
ZvtcVjLL0LFc3PpmNkBwOtu8sqKEtAiOQZsvMFBIy6g8U9nZZLk6jJcc2+zekiNl
oHZ/6m26A32iamIKyYaxF4pdKwAJ7ZPwSidccvSqd2zJ9ascOnXjuoB+68vsOLMP
33DrFWszbiUaubaB+n6MEVSDOea2l2W24M16bQi/R9oYWuBg9dfp+UbB3Vei2mzH
B0iH7pUxNc8mXaaI8Xj0Kz4Tgo+SxwmKR1UK+0GSpuGohX1mYqoMxjcR3mLWM7xo
VXgPsTs8jsoulJIBfIoRArughXVzHvO/OLKTzAL6dTYNqQ1WqrvP67xR16pY/izD
JBlrQIhdU6+aya5PPyqVwZxc4fJYUJpZ1qgtrTT5GsOvN5Vt5SrMxdK78YkHLAtf
/JjM+nhrinb8uwRKSb0Yhb6VtjDYw9MBvy8IKI+Tb1IfO/6vSdZ3aTwT6jM8XUZq
p1O1BHwuO/XmNdAIgCP0xDMr9p1vUgm1TvygSzz9zz69FJJwGOVQz70EdumToJ/K
HE6friXACQ7sWnBS2s0qwimuoG10hPo3BU5zLV1SHjKfGECrQSJgv6JiP6Fa3R6m
IiIRwwkVpQSjzKKbKtP+Lvb/OKkpmnPmcUtsqnVUM5hJSVfTKPJ2WGAJR+H6BXeD
WMyBfEbXnPgZVIOmmFlKS96kggqFEIG4k1mHF59QEvjfAaQ+u4J2/yZL59WO41Gw
qDi55By3rDGTM+ptiDo+fH1OAuvRqDSjzJ1nNKWn/eWzJGBGZFFWEZsWEXvjUKa8
cFgfJtmc0UAHGffNuDWrhSCSCvGVieMGvKvp9nqRbNrDkCQnIswsR91iskF6N0a7
V2mRde7wqcjGetWioO6hK715Gr2FQfe8+sccqU3SfvsA10Vl+M1hikGP08NRXorg
imB3NEcNM35xaRz+jtYMO5d2STL8ExYTV/fzHtYPGHpiMefim2Q+eDrB2DSX8ZSn
G+cDlO79s2DXvmiQMM7ca1064nrFsavRYo06fBQwgfag+PBX3tUMYiKKXib1CTNW
J7VTCp49j2/ar/iwwkYZ11iM7l4iO0mu42p/hN5GnFoZv9dSOX5EQjeYPrI9UXRu
XvmyESnaMmVNEb+tW/cvy2j8BzhTAEx3f7YZhQv7lzfC0BGR0Wb0k5JFf3CrC4Mt
eIBTzbJv7WT09Iz8ceU0PGWDE0/Uv3zCjKdszey0LleRQ3r9lHGKzJYC/reMjHOd
YxpXZvy0gplc/5a9a+FDcLaMPgMRoj2gJq/gzWT9Mpr0cT3SMr5WlK86NNmqQ4Q2
24YvkxX+0h1Je/bdjESWMRNYwF6iOMuDHF282/umtQotb/yfdnjHmvKybRMvAFfN
2TLk4kUUXKH8QpqLZDh/gVhRpARkZoxyUzVR6mfCZlHY2mfrtef2hzhcURaSfdlQ
HFtYatbCSTavJgJl4S1mdy31Lak23KkhcwnB2r9iaDdegEyQ4sxjM5casbXhl8jy
8w0/aBQcpwkWNpoVkEnD1DzLRtxFs/yu2gIkB7PyAqjzu80jmbncl7BNXrqyhOjb
o95gRrFRivxFDtV5Zc6YoYnQIu+fRK25ulldS7Z867RLaeVXK5cmo2w9VTrN6Tu8
iOf4TPSwcNWP3vyyO3xK3A4dt2l5afzSNBFvOrT6m1oW8uMd4Wx+/jnqnGmRHQ4w
jPmJS51Q1BCyTOfQ7CqN8dWxwoOc2t9/kqiAdmsOGaEWs6qARjtro8AWvzDfl4uY
rFSAOa6tDTfBhnxhjQ1yIz30Bjcch23Ncz8zYVE0llCdYJN3jtZHQ0N7yYEpYUOz
/ZpAJwf1u1fHOMfq+q+hckGTN0+NQKv74rPJ+G8tIJxBvFUSEdAPcrpccQfrVY+a
hV7t8cM8JCLWBt/ZPU+5YGUFOdtzO31bZY1srFg59OVJxe4NW1+L/UizuHX5rC2V
dvgeG66ozAJEiatZrx7W8YQQD1FFN6ak4tYBSwL8/aiuyGQYHrZTwCq/hsvVhWKB
VDnuxowzCNvbLsqGHE+rNeYZsJ5Vj3QEBh7BfqGNZoLXEKgZB/dvWdvYjsq33nLI
1NQrrpz7zyJiS5MEwFhCsOHcvBSnodg+sEYnC0HBrX5Ki8X26Ndvi3LrU8U6NXkn
EbUD9OZwNcb6R0hdyefPanavz/W63Tyq+IEHixqaSKMeezcxtPa0ha7w02NQ2F31
1L+czAYyix9Db2yIFaHpXRMPgf6EvOBEr5qZ2/AASu1F2NpFzx5klU5dP9g64tNK
JiclFhRGGvig92YLutKqtEo/T4zGWloK7qKhZrhjbxOM88+jxjbseMuJw1u3wqT/
b9BYuEzFKAi0yUJ65cJRFIT57x971eSF2Veuhcbi8IVCFrqVeB/88FBPnP+LYLnL
mab4T0sCfzBl1E5e7B5jHRuUvu57PfFX8K0lWEKw0hfOn2DqHYOZLEizMStA5KMs
UZC2h5s4oEZcGf0Dm4ZNataiB+BaWsKj0WIk2vWvuUZP1x+bZRF97VnRF0CrgGl2
jH9srPIfmPpsREF6dFGotfVTokuVhhvCQ/RSMUbWuQJ4A8hFjogCyt1HaH8/wPXd
hfV5ORkIvOgttZt2s2ROwThTGDRGtebaRK34jWo+sKKVG+a0U43zWAL8IMhKQBF+
KShlMFC7KJlv8XAMpNS1rrfXp04PR7ohJUMpZHyQwKFedujxFtcqHsHyKX+rftdy
lo3Y0YR9xrez/wXO2kLYqLHzUhwpO+abUiTCnj1vZNKlCQe0m32Uc3c6ahdv4b9X
nZaWnz1tcNdenwGoY+YFC6Q6HmGkHL+dQ+exvdT9AVFje4uXw6K6ZU2a0rFN7+6H
Ef6nT/fLbXDM+QTZVpLVw6G9wxbhG4PfHnX4vXA1zJA/eXf4AmFj2FuIjO/dl6xS
9Bz4XylLX6gK2MSNKSCdJEuuqhE6rRmscVCNcPAZ05VFlOhx1JGRuZZes5/scdka
IMhvQyxEn6tdJZL60nBpVQB168ATtC30C5q/gUDUNZyrDE88trCkcM1Ikjbb6JnH
CJNinRMflxPXBX9gI2elPWTv+sYAFdz0N2mv7EKtSEw2aaqUGJGtu9IVk20PvADr
KuQTb1Z5pNVsxP9lFq1xqyuWzcBtX57NVswS3cVIgv/KToMhsNVjnCrerL5jM2JU
r8EuFOCzsB5bX4upiN/gvRu7Ddfa6DHe0Xpwcat7dIvb0PrY7yBOBgcicbBADunY
K0Ehp+WV4JFrHOn20l50GVuh2IcS0LfMOEQZLaF4KbZqpLIkvI6Hz0mFVenud2VI
V42ntRNFWDtssNWs7J7QjhuGX/uW9rUuBGRVH/zpfWYBBMpnBkv3p83eq6kjVwE0
0hH1gLNILyYQaTZI8MWzcsapO6F8q93EDU1Wo+lJbAyOhwYrEejQCu0MovE784QG
gcCbMdmsE36VHI9tIFPwVMjJZlmlc14sV/sCEhxHhXeMFpsIbztgwEHnsYv4lDnm
+8BQ0VyT4yXtshNdyKnwooJi/5lUyMEfh/jCKvnSIRKBzz4w9pYsBqsyD3KBxI6x
spUNY4wFxIJ13vcy6eJ6PdGBuWZf4xFiqyVo+AVjfxvQl8+D2xU+YrOtpz3mzxAN
//mWaYjjqiVaKCc38mK7kPyYfsE2sy0yhVrhULAMpuifPhOUkMWMwJxcu9jyW507
VGQYyuF5ZHo1z/XvsG7ix2Z5wpZtfxvIWo/i39I5ZmGJgylFC3qcOQyIKlhKVxoi
dKMhIkOpYin6bop+/LeyJqgfnsyU0zZES674fJk43H9r1Oi7C3DmWya3g6Eb9CWa
CdZ58t0SEZvtvL3u55SDoPagcsFm0onmtw2sGPYNN/ruPmSrCWO5ej8lZIJo5bzS
XOA8aNbVfIzZovJ6N+MIF71jE9/W2aKjzMUbkawBoXARTInzCOQjyhdRNS+9TEWS
FW1DLjEnE6r2sT6aTuLhSwsTUYnoAXHMsGQLLNnh6YviwJvRAV5aMLD7nmcICwZD
ecW5Ksk5vSucB8ANjdrC3uKu34FUdwItejD6vuOpZTreWUwmDnPbzFnHUXWtj8wK
4Fp4qgKvfr4HXzgY1li3MZpm9V/Kbx1yhzPSnrJcRESF1I9ovTREjteI1STGXcor
BKACW55y1g+Y/YHvx7XMmQsmnm4eZxbM3Mgl2CG6N+4vrezKWdMTy7y+nfxKosNF
LY5OKfw7kl3ptdlNOE3E3gexFi5++aTZaOEV8QE62He21A70TTQUhBeyrPqouhC0
1O27fwlxprWPpnl8RTQfNWWpE/deYnmG6wzr0w+ZTiD4h4facGKS2iyLjp/cr9uV
atfouAd4OFWHzEgq9cHo1wTPcqirL8RE2dlf3fqsdoHE7EySV1i1nQBFC7D5K/Yk
R/uR2Kv/GbUJMQfIQ46bAGoxkphWHbKp0NEzNnfdo3mOovUy1Spi6emIA2IRhJeY
9tmMU3krRbOxPCbSWM2X+iytbOZGkRVyT4nIVlboBKPyvHx0ipplaX9VL49i9IN4
LAye+VDUFbw739ezZZnhF/p8rY3O2dfpjmZE90f4pq0d7+czJhMSYVThzwoHhqpm
70qBEPFY0bwAZ2P42wIWWMXzzSXV+2RzHclh7onU51Z0seUHVCXsH5Glq6vIeQ1E
1lLjj79DIPoge8BDCc9wD2Dx7xmpRQpHzJyZTkK1HO9yylNqljypOhoub8L4SIWP
LmggYJwgIkGJFKu65wFwvRg35QqbiOZ1gaZS72i5LGiFq5YF1tYxl/ftJwM4i+uV
OWEo5KeFNZvQI9Z/yiMREWjBvV7h8zKAtK8rYapNyRqOcKONXmibSiWGB8KySni5
ovhCMTvOKU1eRWMxvb2n2r9ZqhGzyUobyQzJJ3QKqMyPq47EgsnLLwqaJ2ShzfSR
S7eJXiJH2GT09u8c+OnwoVNwItrz1qhGAdcnUeDX51r1Puj8wun4DybLeLzV/uVW
+ExeUJjWGvQxmJNqonVknOP4jCADgxHsrKTxusXaXWGLMzzr0/NgMIWR7K4Qb+nn
J2r1MOsR9ufrLm4BeqRHfAG4P5A8ih1VBqCcj+2CPpCec6v8AjBhQvR90qewFl9H
K7WFnT5HcISRypfJ3GrB1Pw59o+Z3AiyRK/g7A0KkkvxuJepQmrhaEq9wob2/9mh
uKgGrrHsUbEiM33t2xYYumWAlN204IwAEJL/fv7iylw9k1cthxurcul5LrDACE/O
I40J2UDjXWLTmbYXi6OS9JkXLU1hyRJfk9maDQRQO0b3WfJxjKJsvlg6byMXXarb
fFjZ8V4SkmhJrabg4TgeOY9Hg4hMzwabOnXBaSWvV+8Qe0Ln6J1bcVXoUA7+XQXz
3wAHE7YoZlnCc/LQh8sjwh1pI/XUhmGiTc2Dw9CMiYyNtBb0oaLqnZ1Zohzaur/s
6vGRExbLv+j4pRJlP0rJNKTuup9xkZ7GPuyLfifKEe2J9NELWWEaDPixepuU1bzB
XLQpxU26VguZrgOkqdpb36Cfbp/R+rPAFyN1PrNEjDQtrIIDrELZCFEoubHAWOcK
K7GD6Mel4LHResIm9lztadgR/XHBAqd2s/Dtb5yoo6EhTnhrw/isOLbKOAGiVegY
BfDLYej7o1hxWDrbH7eozHWY9IhcYL/tW/4Y4VMxKDO1R0L1U8y6UzG5oM6QUWSO
Al377LnescEht9U4FT/6UTvxmn4ZHSYQejqTAZGKAXtsgatGhouBvQ9tSXEMe7BK
UOcVQGFuRoDJKGdyWEW8PsUekh+FGgJc30vY1Onsh8pjJqW+TJZRJvxNjgNMy1ZN
Sek8IKbjgoa9i/zarMWd1bHYTJ9oI3nvU7CrBWbzr9X4hWrLLE9G4xihMoKdqwYV
A4eqcM21KzrOz/2555doiT4nCR8phnmj0g1hk21qq99Er9/oGiTbpT4ayolUCS0y
IAm+BPRwr9V8LTsIHFlLuwxhnkMOTxPSFA/p93LHctAEBdJHCMSIkYAWT5wQSa1i
xxj2c2jR1CmFdzbH20j+zWBYh2Z/puG73j7sKqnfJPyrwWp60seQ/CkgKJx24J4t
farpyw68SeuyxiV9GZ6MkaFpvpAShBtZYU+XuOtJs/bGJH5CR5iNzII5ZbSOU1dp
NGuVHX4W/cbhFayFxkw+zC0z4fJ6MCrl+0IzLP0ar/DOp0wKwsfwMMH+0xXEIJpj
WESO5XTI4j2+AsU6GYiT5udtI8w4LEYCjsn4BrxZq2++/kfYAhPW/e5kQDiKikJ+
uMaDFQyODanmc3vQIvAdmhklhlLzIrbPIOd78ZJbUaNEj3Nt15MR8nWeEQH1t3nu
2+rS4x0o9Mb7RbnTkuZXccMix4ypT3ZN/B2UITgRaDyroHs7PuL9Awib8Rsxx/zN
cEsgBQDA0sGl0yYcRIF/3noKr/482uEpLPUZt3oSTGLbmtawqzljXMwy3Kaiylc3
s3aC5bLOwOESp249uIkB53NUYwJo31DZJ3qM4puEd2lLyc1q0J2BUkHPjpdtXoX2
8Dg2GFfT9vlbNsIC33X0K3lU9oWTCPqIItzAXe6QDNAD4J5uZkidIwQpL+pqzCef
f6IKu71PUkLRckR7iKBi4gvJmxHU5C1nE8Qxs5ivbllyhkvbh9wBOkpTYIKq9DeJ
zK1F9AsiLwnpU1Ri0QDPrxRtpakMaPAvemMvu3btcHMp2M8RKgyf5OMsaU4w2tPB
7igtU3Y1sUEmeDrnbnZGLlp0Ok0mpnlGgc/XX2iNq4leKOli9iKob9aWGt0HbOhm
D2zit8+xPwVNswfXBfykcOSiDC59413Wh4xc17M6Kfr8ekM9fUqODr2ax+1QiUam
VvsLSGCZAgk85qOjGLblhRl4TjqQlMFJn88wxqcBD4EyN/RCRDlCU4S6T0y6H6lQ
ikRWwps8X2Pb73qyYlvkQ/Dw6HdJrFj9ThC9d7QWuyyJbBfn6h5q9SFffWPNd8N/
oUJh9mCBERstsYXWjA2RnmxAHQ54qUpd5SqVpBWK1ARQdnqRxJ4cChTgUaAy8tV5
WE/xi4kwMZ2aHLPumEjOO7cRBC43BkmdxQ9uSOjxKKhD/DB7IEIDH35wAuYoAiS0
NpyYIKbbO0a6IQLWmifQ1TijnUZYdMZ/0cqgBKTQFEc0eaY26laCmTsvdqDqzpeM
uoAedfRZHvGznd1hVhu1TbQOCewNtIc0QO6NT9ZKkI7GUX/ql3gXsDOzYU/GzfJx
0Bzg4sgAMmOxf1q9nT0p39U0H4VC78GyE3l3HReYzKr5Abn58JzKh/NUy208kGFi
hfsFLgQ5jkUnyd3B6AX/rzlin4El/gUQ1FkWog2xqhsp6Y1sFCxGSZUYu8lqzJbU
3i+ljfWEekUCnJi7ljCS4J2xN7cTKkrSJr/TeyJcsCU5imj76XJYiJE6ZmRb1dQ2
ylEGkRMB08znIJ9M6pej7yUSuG41r9HTzQW3d4Pkf4jUpTe/jVjVX6BNHAM4Za5G
ux7DxdM8ziU3u+Xm6FXD8S+HTGKRfhDpfGzgoFzrx0MyI4nQJuoGH9hv9cLssGmE
NF8w8pPezNlQO66m4v6caMMmmFuBFXqDt8q0vfvxYgxhcXKn5jJxzIG5/HjFygLI
e1kEBHnoMxZjcwZMjwiwpJrelGIn/+FlqrQvUHxXsXfpz27+7fPYxg/LIgyphorq
6GB1w96CZ6Io4T837g8LRpfs+Ue2h7LIRR5AvxaF6H4d4xt21tVXEewuQ+PqYh+7
bWzNWePTA6QALIxq2rIZTm5wsu+zn6jX68fsroP5eRE2kuwToYkIzWKWNiQw3x9H
CUVCfyy15ZPV4Ogx2knYWBdJ+rttc/lBoDAvQhrvH8sOa+tYc1EHW7sjXAFSyuGV
LYHtQUU7h3j4miGKtgQbPk9j3+7KMvg1Q9i7OZw0P+AYuXEzjttuEznW3zwQmdUm
jInn6O4MGJYU4d3m5jY7BPDTfpMAquZMUt250rs2gCRxF2OD0FrJGeenHdk237FU
bYDWm9LbZS21DHOsuUcyY8DMm4CUR5jVmaNlDGiTwo+eoyXamq6fMrl6SPI0vqRg
sCQ4WFY+jTs1B74+AkgpYwaIXA5aQBbwmYfwlYhQdmtrCP5EZrnlXKZPg0ztysD/
c/N4qKg2H+Nl9MJZzd0HrJ4j7B5CyRn5bT+vgWrpbzd3GrfBBCIHXVE8RbhhKb9A
CNv0QIx6iGH86o1NJ0CzQgfVJvgL1TYrp6pnY6AqzonapyR71teVboLMPENv5mI4
UUepgvdID/TIPn4fM8qRRg5vsihNl5S/NiLC4GuMAOhaqsfPZZEL3iefzIGzmMVs
WLjXEw9HDKwsfnlQ27beiUboYRhp5GiNn3hl2VdzcVWu0zL8sv2LIrWXK9/8+Ru9
HTvRqoI/4M9/ooNlJJmHO296TLQw8P5mROvSauRaAGFhKSGLNhEnaxRIoqPNhqe0
36emTSnZHNuucUC+dtZ+fAjunXXsJzk3s5gedbb8uawj1TiyV+7uhYZjUWZvXeMS
h5leHIhDh66osBYUID4AQdyJzzO8C6uw4HTeFjlAkqU4+FhAQ9+CHnsmb1L8pp54
1yqzYx1Odnj4G3rpyk1AI3jY1uDTFkRy7fy+DeXtEryhM6uq5dqPH/QEQR/d09T4
kaHNs6spJLieGd5Cub6hXNlvp8zHPhohT5lqMxyLs3HVEv18t5CiFRmHpBAZ/XG9
X7dQvp9NuQDPGYvU2l9eiMsNKHBB49J5pwXSQdy8JFBAowXwKUSQvnRh7YV9n45h
6m25ntNRU5/jsV2SPfrrREejIsjs27OrYkAsuBU6j2mAnkV1UAwo62uZEXQG9xgO
7ontA63wCX++zUcqEfAUUjCxXDshkTFMbN5bWDiqx1RjyDeNwU/Ne9P+vaA+qxPs
D1jTKjRmwUD++A3j1WrvpSz6y4lOTGivFfaBcjo7b1KtPfx0mH8TpzJ50svUN99v
4kUXZVFSJZoKKvnQ+a1AnPkhEgSopihtyERbDVyQ+I+I8SlKmcJk36WZp9+lN5GW
bwVK/B6UsUmUc7MiE4TJqCbjEbC/LnEZJH/mDLsrCMbQQ+mR5+lfIiSQ4/Sz+PF6
nOTBfu5ffiw3yiUO40J7yPj5/Sw+unMZTTJdPGtLalTLqpjgOGV+SCEhO0kopOW0
mBUUrwTBY6Nrs2yDma7qYchC7hJjnQqnn+aQl99rT1Iv1AZNBz3mtLC4fE0W7Mko
Xmxo789dffvNtiIofjAu+pdvmFCOm+7hijuOh9XVlT75hhb3PCHSj1Nk2Aiauy19
xQ1bNFkByLOyjkYOUBpJZ9z+Ya/EsNv8LD68alKP2iLmoI2CvbIw74hH8thn9/7Z
JkZLpGOG7nRDyt6BBX10Ekc5M99J7IlXfWS59+kdAXX1dIYCuFdrRLkVM2ZmHY1c
hQW/CbRc4v5zyu1nTLmSin0M9bGaKYUvl9mtPJMw3iN6aPNURpcU6q+kWj2mgLF0
E95pL9i/748379mWMNyd6smrP2kJAr0IiMfbNL9cX+hioLh/OGzxCyIMitMh3SMI
/I4Bw8eLLWpYL59AOHJ+Hmu5oI0SrpIqLjtLNWLuy1KjMzZvjWgw7vmfxEOUFW4X
QXX8F1nKvW5rIglirK28OGUjO2ZuEWkfEeorLV3X9uRWDoxYXQwfyV+YWqJsXdB8
eKXZu7UUkQnmWsG2dAV0s/P80qkrUkHKG2CzB7JZenRzQMu8B2r32+BW53u4hDD/
aBO4853WD8ZN0i68RPokpAjwWi+4qbUuPDBasrzjQagrqIZ5LaxsfDFd9AXXCs72
T51ByvZ9ROtXEWM09N1XAit9XCRkFh2j7VJmoFXlvTAtHWvEqoy9XjXt2AguFz7y
6tbwENuv5uS6z16oHVq2WTsJo7LUgnRrrwjYouFxiP9NysriZK36WP2HPWrrUDgi
Lt20Tiejc2wyYJq6uQ2no+uOR1KAN3voZOLC7i1zn2uVuH7DYkXwm1pkH+dREWY5
ARXNahQMo/eNXKoU706awUdbjkhfjBoWNP94/RtHXAnJEEsqjaGNl1gc5mv5cYea
6RYYreKUvEXyDtp7Y9GopTXWmj+CCGt6FejzYfUpYztavqXZDB9Z/Zia99o53BTb
MwdMEQ8Xm9lrqzpnWL2y0oxPsbAH+oYkionoxg0Yc8uoV94cwnWFCm6SadhAEGY8
MRsV3oVWd390+lywvblqsADiFR02BwouYLfYQwABc9CYqGhnGWju+LrPkL+pM+JS
kmG4XbmJ3A9CAm4bGMxpiO8eZDeQ1/BwFmay2586ll9b7QBdPg8ZMP2XJtinHUyN
+dIm4kl+X2q8ARXhViX6yqUqvbHz+JDlA+YXsAnyXlSNTA4xDsOKg2An0+i5bjBR
JHwWaDOExfaEn2jD/WYEr3j3C/nzK/2DyhK9ei7E6L4OQqe0oiD7gs2o2KrRP4O0
Fg0VQXahgQbTE07NFKGG+7fyyN/IwsfF1w0Cx0j5frT6TJR3Hn+0aSdhXxYGFIK4
tL4MbCm062LKL9UEmhPjcbGSoXUKJ4e51c2a1VZdv9PqbbcwDQ3iLWoc/DldmHka
CWJaxm/AXHVyK1asNmI66IC9YBhJJJOPVMbktkAEZPWQZhLZ04R+2yZi1Nj6cWHi
kSG84ijTKGJPm88RlGekjQoH+X3KQEBw+0fvaGltwzRXOM/nQ+xzmR1W7VCZTjRn
edwWC6hs2OoawBO2y2uavHCBugpKaEwF9DTjHfvHVhIzu+ozr+6sZoql4EBR/Np2
ty4zYjk1Ei30dpgsYDLOVw/lIQnwikfYCLkM6R0FRsbn/QPOqh+ZQkgl56uE6GbZ
YP27NfIq1rYcRDPhcZW40FC8JfgkVsYlD+f0rQhk59XdX85RgNF7Z4BLnnQR7o0n
WzekUreGSLzMnMDfGNspPDYYw5L5EqtUBcHBLWwNc92tCmbm26u2Rg8sA3NJ//wr
6jXRK870wV0F2YZcNmCWU4ZnpamhkpbTNwqGyw7v+4nSYSgYDGqnMcY3PxomDxxt
ZIc06al+Rxyi18JK74HkEX+vIco20MOwqs/vD+Boj1N1GW00ej8e9dZPs7qbZDtc
XkZBZD8iLN5BJOyHqvqnQzQeU5O8vvWF8hRvui28gphJ69QRQqRzWciQhYIycAnU
AhR+xeor/qg+8SWuMqzEnrf4szeS3zxg9WThR4EubTYsJaAbX0kMoK9CcaNBVcA1
4z7j3vlc7d3D1aZM+Qm311l1OcIgQcC/yaoNN05TGLJe/x/6DM2lmZTzUf/55BqZ
V00eNgl4fKYBTegXxrH55ZZ04YXF8vp1niwgted65vKBB7xx7eY9/PXCtge4Q11o
X+WDAvFHh/cZ1JYLw1oNmWWPURCKsQ9/PxyyoezTmAkzhEOD6b8QbP8KM4cl88A+
COyvqo10wzsaNOBiYRtGrOMc+rFSmAoqnBtD19QVRdnItfUk8pwPytPBSAJXx6Ul
xIbM92tYR0pMmVqQSXAU28V44OCJs0sBd0l7riBkFqwv4SRIT2nbxwzk6fk+DCTC
vRay8+P43m2Hzd3aPm1mX6+rIrkVFS8lS0MXkG0gfjL4QtgkEVDZ+UoVjzxBWoVN
pu0GUs0i4rZD6XLWE/hND4HF6SNDLdU7UJJL0NkesuU16JAMjd6wsCCqi8sQtsji
0xQcr7coMLST3jxi7/oquyDJfQWq0VTyRzx/3JUrOckmWLJodIWIXFxLpKTVs5BA
Elt78DbL/7jzPxOjxnwynWBpEuop/1xTFDXg6xKzyVS94TlHZ9LVwdMg9WKlomJ6
bU/InMKOeclmWzkL+3TUEq++26XQmjWXGWFpB4KcGWpdg/eQXhEYSWyJgkz1ER8Y
OQDXEGlgQOfOZBbHatxSW+1Vig6WSV+N0WmllkyCR0QLTzN+8fJKneCsJH7xpRlP
y8rUA3ZxblwtFFnaKIjC9gjZby6zbt8BYbqW0ojIsmQ7vrSwaVXSd//Tkm/fHX4S
ntmFTdahA6weHJT3HsO2dhqmWY+9xvClNOo9BPTtyNM/IT+tYfIEGbhw6wRTW6c5
ccQ4jd/DaxCbW+eGU++4En8jgugAg52Itaj0DjGWlRi/6xEdpW/h6v4blYxU6IOR
K0OwHZQmuZsZD7wKWIiLqU0zDE56aMhR2j6itD/E9fW2vRtD/8/P22x1UtOESp/q
kHCv7EBa6FBam1fA5Yn0aqR8BA9Q0SzVTDIVXBCfluAyFjQEER//Kx9VpkPajq1X
bVT0DdDhASvhrmOE2fNBnVFe69MWD4oQ9RGmXXf0ByfIiQHbGrwOtw0Rji0nMDwe
LY+GWPbXI34LJav1ehZFln75evgl30nbSZ19qFeex022uq7Zz3h6bKTOXGK0qvGU
oHnDGnKvQALM2+XIdr/9cRMU2jOjI4ZcVhztRSV9ONzozrCHplCZZwyB9tYgpCwj
JgQ+AHb1uSG4Y5E2GJO+GMurUjAkSFNsoq7ly9RTrRzNI5Rti8ZZ8hhrGKlHcT3B
HvI6nktvVUjyd6GyZneNbpNQeQ7pILu2L9pysHFxgLnK9BHdXI5CGr/odhpFHImV
Pl1BtTBEXU1aeiIDz0Wp3RX7UG0rU4LghZQXg/zMOlNRN+NKTZ1UUA9L5jFIPYuk
sotfWmZxuhaL94nBQQ8grEhquJVQLFVzHxkhaITmUzRtneNDkySMuCPjAiRgRmWk
fdPI2Wn3+Cw2l41kCsG2nvPeS9xnAnuKTp6XFycLdSmJtum02neupUDhtNmLlLXk
ttZL3My7e87gJG2I41ZT9sANr0Jonl20Zz+ADNLe874xW1IjP1H2uKWc4F8S7dQV
jCgaKOmOPJKWUyYCkCh+zTKEGBOuktI+XvgW/FnGWhyMwjUrR+lrEyTMvx47OTcX
2POxFb8Xp7oQ5jjTzQR2mSwOyoheTIHroq0k7MFEMoZvlGRO3qT+winc7QOahfxo
GKRJi+HjzfrGVyGPXwm0xCiIZw0t4gj4oU0kWe0P1mo2bYQlS0mMiYLGMCILB+BL
6k2qEg6Xw8KA01rd/Gbsc7EzUAbXH3LGhWcTn0hFXA241b7QGZV/Dxrp9ds+rVqu
fcw1NhnFOQ2lWEl0m7buHQh7p9DFUnjX7fj8yLl7fBQCTyUxbydna8o5OJHXiiLy
19aa1wAnbZoYJghO358puXDkS2z/HWAbp6TDQnnaZt3ARZC2MgkgovcR5BBRQ+I9
VRtj0fwa3YnZhTUTMHzminKh2FstZgT7GTYIdiPvhSRIwS86lJ/lkXEKWdoJeS55
LMN9bhU9ST20M4F7mobJJte3V7fldn3MM0GTLks/m4KGJt5LqYqR4ISVftznJ9ZD
1PtVCernvj7KFfEDyjDrv4tQZu+HUjcvQHtZBoenvSANB1UVIXs6WIBQqzFtulxg
uOXgJEPQpOkL6Q/lrN4sbblxnKi94VNa8oa/Q9vbR0tbdXcGApYayekU3RE/T9zI
FFLoBkFvcbSZSY7El9v/UGrzG+9JwJB2c+aTZHaIBsw5Q6oX5/zoh607X+uxbx4C
WQ4IlU2GYJrNR42u3wHw4duIshc9wnJc9WwJk2agdaK7bNokhMQok5Euu86TxRYy
Kk4d/AOsPDU1SPW89uElgGBHCLV/9jYWs+YEA8I22FVBZp3LuzEOWFSDLmj1zJBq
J33J7lcBV2hKv0RNEPoT2ag5u7anfYHe2Yyngb12YrjU+m6H7VO+C0QXmSoxVGFC
mipTvM9UTreEFwZW9PWG2s/ZU5A+p4Eul01Pgkkf8SyIQRoBSvo3+wQ5Fic4gxEy
05epk1j6J8Y6xQ5ZxloAephzuOmeFqi1yKybncIuot5nV3uo0YRI1M6drYghdnmz
TrLyyjH6HejbjHTk//1BVLSmnxBBnr/mMC2NeC//vOA1Hkb9PHUipFWqPc/PhMW3
s51mGLM2eVdmbPuOGaBKnLb1WFj2LvNA3S+osQQj/Mrx6grIxw7vYNdnwNv4i/Y2
BMhtU2+Tykp2BNp4FVIpEJjC4hkeW0/dDMoKxaqGR3qrrPphrPcNUnUg+szOwxkl
ICkQQT9Ekz9o5nvfDKq9jn49ZXeD5+p7133Il5SWY1gczCWBOwHCgUzx/lYRzykC
ZCJVH9E5F1VzmEdxrifLLMSf1b0OxyXeNdlpqu/G+n/edHQrinaLw3iy+arbGQJS
Fylyq3VUQ1Lgac5MarXL7OY4mIrDUf+dWaUDIk/ewdtoUj1+I6lGm+ncIO5w7kx/
X41Y9He1RZTWSGffrNOXibYNAke3z8E7VsRL1gZG0WPTFJHO1Aask1d4Fw0XADBM
d72g9WQNLXTSrhsu3n3T1gTojEa31U3dS0Jz/j1okGZJ+6WaVtGoWAmE3a0rL9Pf
fFOBlOiVTnRH55TZrSsR6jCi6u551PTSJybytql2Ot7v9f8VsjcwwWQmiNdkI3bq
thq5a41BeaTu7i21iKAvv+YpmPVtNQmM8FKuCbSK00kIVq4uyQ6E22iUMG8kPHZC
NlZ72kchPRSUaRX3/St7uFtpTyMaJl5XCF9inMsuOM6NjL+/TiKz4W44jPmtUVrm
22zeaVCy6coC+s0LUOxzt4A4DeFh8bMa1x4+UpvsghFZocnsusI2e/gR2Fp0Q2Rl
cKUCTpXaBLF6Aj+fljbS7pLs1q+OJacjg0SpM4SWh/rbxhLLXB/agHz65wvWydf0
Rsx/pHSPL+HSn0V7J99gDFW/zwJIwW7EQXpvbcB2mtpSBLQyfe4DKFxy9FiqaZGb
ARk6RDv2teWGOxF4kqTvPcyzsMSGfKhQTsSW2rxiee4YaAmJiRuJ241n5LyVCE1b
bHPqCYVh/ulIT0+XVIlS+q5pFw35W69/erhSlu8OxfPs0XjfQjJqlSYYFCYSMvLe
WvLD7tsY2AXnWoxUKLSKTGeweQYtyvQF1jF26/84oMEcxiD6c93rbk9RaAp7PZ5D
nQfsVzzTlBmOH4WWSyfjN3hXgsIbu2HLK4+QzTEz3pR3ahbL0zJlCWFBrn4NEx3p
hyFCH4D4+IBkTyEk/12oOgPf7oqiqvUgxsXxFFG1Og0h2F+XCfp4QIMW6zq1jFR+
YtKxPHYIdOJe7MekbgfT5MWcgMOP6w+MjYyo9q2zi5q6HGOniC2aW84rYsKFtBT2
N13isS/c0/5a6upmMozhFg/WwuuF+JQs7EGfKAlMlsDTaC/EP8ZWJUbmjlwIuf5X
ocd1dKMKSSTEyDdTB9UNJqWpsuapltXrwyboRq3hToZXqu4F+8WdgeBs+ZRFK3w1
VMuYpyrI6IhwKnZeWF+ml0/bz5tWIl4uMN7ULX8vUouABc4a4qVpnLpwXDhuIlei
y8RwrvcirN4jFgy5lVRnSTCFYx+yLxgPLH1+g4V59vukwlfUDoY7guztbw2edPDT
Q4rzLc4zPcrSMw4cZFmY9Td1iJwSP7mG0GoDM57Mvg7nAYl4I66ah1Oh06dXV3T7
pEbpxR+KVOhsakwTdj/GDlkcUKo7Z2sADvP89ISIW+rCr3GXoKCUeOxKV9s4kadv
rrsvKUlJWoNfaOROppkv0nDZf1huJU2YA8ut6OPXFxoUsg0CwBGxgHAH255qdRte
1Yhcrqtvy8KZ3nEIsUDSAtzgTJzPhpwEtvfsmkNO0i2rhk3pzYvrhV/jK0KrtSBn
UNfNpKnvcX8OVtUkoFSkyLktM8vihpzRvW1SEfnRBZyKPa8m6QDbUwwLNSBucRTj
PDcZSSO1BHlc9VJ50ydrYk0KDQ9FcxASq2b2r9B//A2GOKfXycKHVxoBPgsHo+mA
/0reSntPwn4/jfE/UjOZfzSoGP7fKr93QWT2poBeepIX+RE+DfQ9cREmn7f7uIk5
OuvR7LSBaKvHHteRl0yZbg5AS0pQ1OhUXO1UH1VDPhkliSfVgsyAFCfsBoMi1LhJ
cu0UMvxGmTpzTl8iBGBk4RwLLA1zpV4ckOtQN7CI/JNUKoMO6L3Ncg5ReDnC/PaQ
CFJAc1RALiZllwvaGt4lme4B798X5/QzeA07vPadFRKcRMh7ik5zd7co0yYcVlD1
mdinMjipawia30tsBUXgTMXAr/T/9f4LA00iHf0uxToYnnJBmWZPDLf2rE4Q3AuH
bp2Ks1bMFmcmH4fY6AhA5OFCTryeBbnpWBobhSlRyj9Nq8VK6uNs7TglwNzlfMf9
jPHrwS4Q84UdQY58yyOuj2Krb1XDAqWCsljudul3stZNPYmKXryYi7QYNQuE/0Nv
NTFFTx/YheOEmyULtovBqwSxz3EM9EJw2gkySDzyZRllhRRqiFizA/hBdYtcwXGM
fJO1M7pnql+8cKzXEPSE3US16x9/ff8GEKAvTWp3mC+clOPd5Z52TYlzZwnTOqks
i0S8bxstAHQWPa3KILVky9+xv5buqBA1JB98RiYdIEuZAeym4eWYstKRA+DPkTbO
xJmeM54tv4qIFUx4iIbGeWU6h/EphVRlt3RYLLVqkur6US1mltwDsa/kOlhfbBaX
PmGbYHiLfX/op2QKXcSGowLEpBrTImSPSxWwOQrr8TNXTZbBLbK2Tl41uirg3fyI
aa/3AVJWyuwjndTuxKpTbfTk2g1qm+HDPwu1sCROqQ1oGbFeOgERKc7rkFimXvnE
UehOytOW+Uteb+UKyLlNEvuWN6UESJmQ9J2xu50hl/cwt4K8UeaWKKvVHq9aV2m7
OKLq5ZyQxzpATnpqvA1dunr2sINaP2RQcbwDLV/5hmkIzFqGrRJJJVyns0E2Cr8d
AS0YdSv4TZAQwIQ6iwn7Af5uoCxbi96Rhj/a9lP8hV/bnr9SV/9IElsyI/RN2I53
7IRFJE8wdfCR4DQ/5pg6gIlD4kiwBv2tFquE8pWKO+WGYwTCBD2IiBbdRkqJrbPJ
KfIx5S8zsviEyK+e/zd5BQjkD7xnAgy90UG2n+Vx2n8n+TzLTzrb6VjsaWj1HDB9
bT/t56FXYiUVkEywL0p2wbHrnBW/5anWt4p3ZSMMAvwsAHbVl9PnD4SkFUbGuYKv
rldiHGSenNtoC2wxRW4oVo0d0d12jSzYKIc+pnLg3plakR0FpWx4N8V8w9+wM0sZ
oV1HFR9DnJL+ofW1t/XO6C9vmw1vuC5anFtk+QIrk51pC4jITGeLEEbbMkdHUWH2
N6WqqWVsRJod2za0/qDPkbAI4wyw0EqhTJASXKfjWrjpPTpXBE7u8FJQth6fEgNP
7vwAEM+6uZzITHBA7DNX2yVZcRkzvOIed8B1xAVW69fOcsMlIO7TjNDhNOJk1cRx
PyeoYiMVjx468XutLmYDE/peBAxgvYJYVoU1n/LZ7GRFbMcsnDI1XhgF/9VqziVs
I9f/HxbgmpsC84s0GPkiEICGqRTCwU55wLDdRPp/lykrQkL4L3sEX4eYXX5MWX9B
AJpEyPJsVIX1UuLYD3Bjmlh8zObK+bFeUORY/tdvDWYDpa4pme5SRdhWO1X3jRmD
HTXfSi+ojGfGA1Ju3zeOP+wDsTq1X+NLPeWB6eXHDE5iwu/ZHaCIATlVjjKjLEyV
6sZSpErxurpIoklkn3nTHaWYnLsiqb7SFjqn6T/R4gYUl2Skh555nfGLDNZPlQcv
sq4EY5gO42z+oIP8/q//zE7Dm26NBth73WuHOFdMPPVHCxAVcCw9hjlxJZDJsvgO
kazkssY5jKHL5cIqS1I1UqTS8PduOmWxCI+lmsqCVTnpPFE75fLMDsq6B09osBML
+FDfm0Fj57/p1casgaOBXvPQbCfQlJVBfq9xrw5HbQxzviReeHCJmNEvr3url8pp
parhrqNULY4c+bEKuaydEW0TBty7zZb1ygaUoCqyakA6IaNPil1Evb0CDyN0Vfzi
CUPubQTljFO+HNBXJoQkasmik0taO9sRnLLRvHR3sThihwiEIgCBbHIDcB6rO+JK
1oGKLEVyYY1AWZqT2RY37fzjpCB61+jgGBFXhXQHrR2oN3lNYyXA2snUI3HXrrmy
zNmfaxf4qgMfBpb4YtUq0Kv7EEwKW+NWxnB3OeDzXk3QXrKrp1AqZU40nUiUnTJp
L8vn5IlXT6NkGc500rZgPSlHkJmyVeb6KU8XVV9Sn8tNuvgOFQ6xpkZj+cHRyqm7
KzWNxrRqR0Q+k+SGZTAkAnwXEXXPIvyj9fnDB3dotMLEw8FG/X7IxU4dHxSGAwHA
qMjZfSelmTGGK4jTY9gXJT16XFq3VtT0c0JpGeXAdSJZMig8N/09rXoZJ0Qh/nZ6
gVPZuuIRBY45DLo/AqUb7cGb5l74N6mNqFGZMzIbET1NBcQ5vYK0710BXckXzCMQ
lvn+Z72Cym64l4er+PxNgYRqgU93ffsHainZUzAZkmZ0ds2A2NuY5tx45bbm/zJZ
/uC6b6fptrR0tVphmxWvu/EdxaiTEEwpHOPW4QkYst++3KupCoC2fu78+MyD0kVK
fzjVErEX9vcioDEaum/AZ99OTzUESSg8e1/r563qiKgp+GDHW4F4yST6TQHOD4XJ
KiFCbQbhlp10zsTMeKAosqAsnKtLDiXLUKMKZRkjXp1IavWGjLHeRbjx8OsBxJGA
o/lZMYIuJMPv4kLp9aEmbgiQd5IQ86AVLvjW1BjfuPZ/eFnUR7+Pn68pgIf2NGXw
R0o3iROjX2pwrCQ4ifRheShabVwF1qTxoCbeV082IIl6oydHeRJ6BAI5+yMYok1Q
NocZOCdVpKufsFUY7WRMnIi1QTS2OxN3qKNkQ4ahmdN1S7GAF/Xsuw19wPKSYGXN
+G/q3FAdVeWpYuGnncuwjfrPE5CGaJqHZPHUJdQ9R1TrbUgztNvTsVj6MqXSk0V1
a4GaI3PpCuNP69OU0MamFx2eZB74EKNqQGmHRzbpKipf5OzC22zU/zAkbSuUQDwy
YZ+y9OI5ja83QbnOZXmFhhQ4U7/Mh4pX6kfIBfW4PTWL2nSHXg/tM/02hW+SfVbK
xL8zfRqWUA8y8y/L0iITLgDnsB12xdXjbYGNrkqY6bsz77R4zKtHb3nXhYs2clyz
oJQiDatUnwVtkm9sYPLe2IESCiZParmFnYrEu79eZNRGS9GZXsPQ7Zg23qgj/smF
pPYNM6JNbSRrLJH1LjN7Qr2uBBDo2jxYOWQZOJRwbenD3LNuSlyqBO9qEA2qoUOC
5NbnNqNlum5LqTKmJGXsuhLjctlFF8kJfzJYjXKLtILUIjbpPYL34N3aFp2ybmSu
S+xFqr1q1iPthjDHGd5A1jK/IKfU29VBXY5OZEFl/pwbre5NMQScmRSSd/tXPwn/
TDxlCq00aIjX8Dt5pna2X6OCuSgNdOmQqSBVstpqG65clHj6OTDNLCPyoxtj3WjE
pkl73vzk0lXXgNa9vm01oAnD0Yf5H2c4C6Znw7ANF7PF8Jt9cIjxW1MZfmNYhvAx
/3wnZ6rYiKD7Si/LbTIJV3w+AArcSVMptJLWFVUfzpl3LVh2oqvpUEQrxu3K3UHO
Y1xWs8gKXuzSiRthDigeKCfpMNQ19H1ivbGzjb7/rdA4S1o05VtiQn/gfqMKwDBh
OGOFl3KBKFGzEFDZ9STDuY5B2fDnya0rTNf3/1AAf9u2WYPhm/qp1NNaAwpXW55k
y2UnGrtJXrXHu+l5tqx+ikIgrV6js7IoPYgNuI/KANOAEDBn4GoCyLbXP9AM+C8Y
TLlJ8Ohnv9eJNfe/I0SLYORoTRUJVe35QkFtcM3bjYdv/bs80I9NAvFc+f1nK7LT
32TXGzNagJ4Hf+RgfL8n9HZjF/tEmoSpi3gKN3h8rz9WRnbpZ6YTxfuREOdTPyNu
jwqsE7bCByZARMP3rMxeW1CiUswY++iDdoiBkCT6Km6wcwzu4k09HKsHiGGhGWR0
rQ717XUqas4TTbjr1XhmkWx4BuVRINxA4shBWd5CgxTJbWIQ05TmebvpIjzDBy2j
oGaKW8Ov/hgAuDimZ3LGi/4cvniFxQeMBNNJ3/R3d7lJlYItdei1yq48VdBGiucU
eLhbKvN4g53UJu0uxFb8B+EjzxPN3uO54JTLQCSgz3D76UIvNCcxfYakNPD8cJF6
sJ3qBFhpCwyLNH+ioR395xfNlokT4ynBTt/GBqCyAl+KawXAKttNWwNp1yCBz6WU
pED/XsqItKa7HFUUtIIop/pqY/YGocwg7lzzKLN57Rx0ew1L6Oe3qXRL9pBZeOzA
V1vIIp3LIbPxv9f0Ftv544AkXa+vr4N0IYLaxklvB8Sm7nI/b4pUUiZSJWD9f+6I
JBaG0+2gDcYT8bl16I6SCLeF7RTmXJ0pQipYNu0FugNDcTpboJJrLHjtgz+r9asX
sVhe7cqTZI9cXrqG7dFBA9fwNAMo0SX1t/xpgoKVotwh/g39mGenTuhF3z4PJcp5
sTD1epM1vNKWvE4+dk1sZqNsESe/igIDiisOzruVQWBxF7QL7dboHzX83pcTMCM4
XK/QICt1BZuuS8Vp8PD1bQvrNveXNGq+os4o07kMrs3IavMlVnoAQS4Bfy7zy+wX
to3q2zwQotHNDliff54Bawnh9rNnuVyGneqwU+ZXlwhW/Zgj5athxNJKlOUIMQCK
ttRYyp2IophxzvJ9sn4sV+bAZs11JpDQMGlK+YyeWb3xNS6EpmtJ2uiosrOTYZ2f
HJumYYdazLjd6EtvlsHcg3jcWqApLJHr8Nav4JHlnpW4KgiPe8geNAGV3wvEXFwR
ovgtABA0YR6z46HvPOjoZmENrYna9aRr6cOpRvHdiZNQaBcD0AKwZ83YiYsAtPiA
WTPuphiS3ZxcphOOa5L3bfTGEe2QNLo7ok+Mn2EFanRr8hBk1Y3feana634ySt9u
qvq6xGkdFraLCTdnD8rf97MSVlAu7FUCudqdo0ziN1/2MPGPqUHqWTKoIhc6zO1o
M/3tZvBQl/p00BbfoncJ6fFVykVDGMR5Aj7+V9nr04mOePYvCHQQ9OcOBBH/7vvB
Nfp6At43ZFKJb/iU6TyknN/zyj8DCMjWLmTuqWe11eCRrKt67fs3T5ET8ZqSmQjH
FCoUf4hze4E9TFdMrtFEtYlvqjxUFe3vPBZ7VCE5fcn1ZJcNFYAZ1TfUqpnTFuVr
1DJM1pxORqdCirddvLg/YkjbWJRMedzBOa8sSrRCxnHcto86gwHIslHFbS1yv9pY
ip9jY6MdF0caqI2Rudok2COKKExZuhfLI8Zdscfm70/YcYWvkEtelyrY/wUe19nM
MMpSl98eb17eThht+V3JqdwFTexwIhVEnt/8QiKItTl77f81kk/cJvgH4JENp5fZ
E8Ys3K1mi791of7HJqU4GJCvg7soiXfZJQAuW6Msv3u+j1TT8Hh8hrluVRLPysZ1
yaBoDNSlR8aUOHgkxDWcw61mFc3/5iddR0xeVYA6ooV/zICoZacnrjqd9P4FaebM
HFqTvE12Ib9D/8+WT9jOsyzCUV77Oa1g/DW622r2nQ7Kl2Oa8XtERA0XmB0w1+PQ
kREbLwIzMBNhek2W75il7sMP/dqH6sebAqAfljIuUPu8iksmjMB3hDFSDhl6xgev
hUuDX26bSi9brEvUeDXN3pQCPCgDKhKalvK5S7GAmB0aVIMFlZuDUmmRLHXREjpq
I1fe/L9C30kNkxmxek4cDgDYT5dPgEFGCR+ioSVNmZ+3Ng4ugEgUTvWKLq7bnm8j
xnfBoq4fACs5cEyAqtGV79m4REHFDnzqwxYk+RcG6TlUcBCNoqVKf8Sf3a0nA/CA
vfuyKcv0sfNbuY1eHIireyuVUcH9dg6FN99q7299k9C83Lhm0+s3TBKoOKEMQUrC
Jlv6UAlOpC4AHTr0MbbaIjiTuof8VbQJs1poSaKicaA08Aq+hJQD1W+6FM+8BSkh
ehX0zLiEkn2E+dt8tht+P6QK6roC/3kSLStMdGoNVRwwKSo9IgQnLXnjQ50RWqrH
kaNyqIEiIrhR8gw8NfEmi3oXURUyr4FDJDN731ryrMfJEmIII9cy3BMnmD46F+uc
xyLuJ/5Gxzn2YfrsRycLNJ3Z7qNKV2ZDfNs+8zFy9yrfbdOeZLOizz/Kpx2MCmZM
IzRFggq6FAXHDq9s/2Fo4L2361pTBOGV/AuINEr0tEDgp5V+w2og5yyVY3JRPQVc
k1stQPvKaCm8Xxa/gGAwvPJSu8HQrglXBReYHVGh7yp6z9x9iYDXfhATiZH1K48y
sH1G93NRjRN5VwKw512RAq5RB2ORSAZDyKI+nkeI070qVe/c2OIqszGo4g/rbF0m
a9zywpljmdS3XgTFt3N4pE8F85VEMVUtlydQ1LlGg6n8Iy2RKt5JsSnYHxQzQ3S9
JU7LsAtYuXJR9mFjETyvFux4v9og2jhSR0kzoTtm6m71IocXz6bJQWgCFXYWavtD
eZFPx5P74Ew7Z5ksqm6zBuvoNFv67zz9+a3nDyG9z/sWvuNqwRHrFkvpPDqGkQQ+
KVw+KekPHcIRw722gqDQ0YKbmiQYUS2d2J5jCIBKTeXp56Km1vzwuLDsQEblfAhK
Q1Qbc+ZaDxrigpP4A8LoDHqIv/pEkpTFJ2Gxi9kCT75ETAGczIChuuHlcCYL1Kff
Hv1QJ1f6mTAnHDQZoiNqvtLK7Z72gdw89BE2toYZcj4Zr9jBzlbYrlipjn8jR/OA
VB3n7NAJZL+ijtdkhCC870MnaJIsEYQdOID6p82BySCxd/l3eCTfenHbRDrO2OCn
UWH/fX7k/Dkk6lVc4AuTOYQkoPTn8ISksZ+TxhXoWLDGgRcwodGG3rJjqE/QISdt
mZb3fMh0wgDakyJ1a2qDWmym6w9g+3dXdrHrHNflQsVaDMxAlFcS8i7gY63KGPY2
YpPhRnIki8wharGZ9QZ6eD1iuVITCwWNRC6cGAoX1d7V8bKiWkjPPmf9/+H0pqte
8L27XF85nzLgFd6S+JOLyAEWJE6KIbLg4XEHoHAOlDQ11fdEDAd/5YI2uaP+7lM2
CQXQBDMlN087ep+3iOzc5YtLJHKDWtFm6+ztoSD1OYS0GRCA1DWemrqG2tAtkfFp
ycr9s0r6vWr/p7LUQcDkZOhVfAg0rNRiqwZK6pYEukXuGzzwifvrRePQn46dJwmD
K0ktSaF1QwsGnXuRwxi1pk0dywkxXh2R/efZi/OzN0b7as8jaacuFIsn/v907UuJ
ND5jBFTNwYgYe+qpprMa30CFiJhTJOlOQJ+ufqIndAtMrSztNNPavibfMDgUkPhh
3yC7Ko3V8AQcHmPYL/58gGlvGMG+jZIg13CUSxw3+zPZs769wkdYLE26jbbQzUlA
njk+w8Twdi8nhf0wYgGo7VZE1UQUmy+t1iQu4dAlSVlOju62+/uthCbVKbmaQS85
pBAK0xil8Bu/9YNKYppMgz9clQzK5qbsmMeXvHPdwK6+Zk+g4vkdcDujZoSmPGGl
I1J7PdFxFd76oBw6yaRwUlYQEw9X0KzBv/OKQatMztGBI/eeetsJfiZtUZHGFvqI
idR8EgWk1fDmm4FjDporCvX8wKL0dd3csOPK9fLS/UKS4jjW8r3p+2Ydz40bGKc2
kUXgsM8zUlc9iiuBqsEPuQcr37iAO6kbQ7roXYg9GlX0f9tyeonyvDraF4G9o1JF
ex/AeeOwS4qXhnDRBE2PfsjOsIinRNLswbd4au5pphvKha0rBl+VxCKdzqFnL+EG
yzCiTZlaqOU3Xk7LOFO4yn7UsQpBHqDrgxv+egzm3u4VlleBQdPXs+HpupNmLG6H
tmUGUY3H7XoI0n1flUOHoDZwPn5NDcAZS55su29l5fjdQvubsRF3Z6vH+ijpnbZA
+HtTpvJwZWcmBoX9o1GeyB9FjIt7L8hSd7bmxx2ScA/H66TJnvhzsEHs5yHPbPLO
1s71U0cCIVtdAcUZeYXLGRC8mvQTldMW9dMr4Y+1y1806B+ERxBDgfC+X7n4MVLz
rY//LhAXHDVU4i4PAwSDZ1iqvvsUDNNcTWDaO/VL2ldhzP23YHaqVftB0fIEu3M5
grPuxfZlsO/O1x3emdcjOCKEjXEFV8jxQMXoaY2aZ5+Gp/eEwvEIX0E3usEbfF7T
SqQtMZgklbTSMNj/HSfgAADhlaTvTOe2mF4998lJg5YvhXEW2A4iB7a6XSA6CsH+
S41HFBYMDL8uvV8E8XEoFjxFOOtbzuC9C/ooT8H23GgyyQ8kiVkCV2Ufbj8wfJRY
wtmJijrgX1rKHu4zWLh4v4UY7fFp3IDjPDQviFME8CEJbD7fNJoFOBU+6YmAz20j
1wzhf5k61uIroeEe/16l5WJY+y/pAJSSCFnqpRl7eBA//Y+Ur+mLDq8iwU8A/1jP
ZMyT23MAuRSVP/DY4zcVWJos1spumiCPO2QzTWIOKeoSDNlsqst1YYU1D0hrm2M/
a5feWKD9YMJ8roukmOyJvFo39kvY7kqE6sJaEVZgXsAT5Cwad7EnjLyaR8i8qP0z
xrr35bCkwDNl5WwoHPZmx05cvmgRUEw/e+AKRJgGFHBZqsC0ZoXTvBanDco025//
bu1e0jeEDpZaRRMb3cCtsgVGWENKdcwWn7WKZ4Zpt8RMGKQNxaH/+Cnj2Zph14If
qMkwprOwnHtQEAVEW2U8UQLDaxN8C9PJYIfjF5v4aE0x4vfRxFhBborpS4MhQQU2
nmXXBXLIawf1sNRIqJjr3y0Y7BWJrwcA5V7+bopaZye+iiEpozAhe8BUXPPwBCzE
3iiAPZ/KQSr6AWZkHFgOE+cvIwjliAEBU7xRInVC0e8nlgfewJhbNZZxRAGie09m
Iad4HSw+UxuIMqDoKnpHxATumi4R19iFx6IJZZEBPkQwAMpQMUo1oJhmD98Jf2HN
IbBnU9o73b6sxuUo4dYMseuI0+24M4TYl0FzI4ZWMDZrA5GsgPtkPeYMXK/H/3Zd
/ZrHXqvCaRg8PN9KPW4Sj6460mCihnKZUG86GFNpiZtybPeAScGC290z5beDpBXd
MVHZFCFjmzNL3Hv5yNb4msY3W7zaT8SIf333s6o2Mt3ucQHZK6x3hhnbfm1xdyPw
Fyc7Mc+0meTTUElIHL5Co5SSUY65pCg5sODY5ZQ2EHBFIWmtu905OsZwPYO+PrlF
qp6h8rA66MyYVrCZsSU8YMpd79BG9PeWK3vSIHYgl1urB9JgAtCIWXIxaBtAaorm
8ruKkQIwROviOp/lBFOLvC1x4Qm1IPTKoH1imRw3WhKXgqYNKltWgfDwfyG0EF4P
MpjaCMTBMVCcOaD8l/cs/pe3MdfoC6Zh4WwqDviy7yZlk/kRkm8olGWyNEkG3mXu
jC3b5LVtnfS1m1nrI6fEHSdtWgpC/SX30G9PQOBfb8JhFQTbvu+rwMP8r7387Zb+
y2cjR2fwRQIWx7Cev8ReUBE0ivD2N3exAgCTS1HgxfA32hzt1OnhZW5eYu4HeaeX
rzECkKyhY8T83KLzztgMxquzOVG5KiY4jdl0EO3Tbm/1j/iceCXAzyg5e8Pofj0G
rtEannksliWrxKYFabA05VkJzxC9siPYHDyh7S7vRs5RKlMh3PGtXK4qg3Q2FZBB
O2BrzfRhof/LDGEL/n3AUTYXXnxlnHmdzXEieDg9SHQ3Wec1KJfX22snHL/JXQ91
R2i56cXjE37uqzL2qynJWaFTcFP+OozbQAsoRNIjRuAkMy7C41vVCkHyJQkpCRU3
pkrFySUPOArIUTRf31Mpw+oLm1y4f67V4qWICiQn3DbXeKWbGBMNXkL+iHA7Ayqa
SUvWFt0ntA6i4jj6kFK1VGAger4kdXmrAmnGyFlr8HTT+I+NJiGWjxenERaFpf1x
cjXrssmC8Tfrq5G7tYOu1qVUPOu2sQdwzIcNq2+F762UlFosyHbYAenlQL9/ACJW
nF8W4iBO8UgcPxy8FAZqU57fQQEO5iMPhXrt3W4pI7pXti2Jgdeyuf6UQR+tIb97
VfvFprK+O+deUYY0xtS7Lwz5C8xdf8EzRjN0wZY2uMRjuzVUqMulyG5VN2qvFJL3
1ksM7KE7ntFApvTsImtwKlCf6jefHNMqa7zrinLOfDC5mhkfqA0dnaHyyUlJVtDm
Qc6wIltQeXnro75TGN+gB9EzExcUFWqxM4qf3369WQ91eJH1Ztzn1t9rUIDhPFmX
MaVgmJc6P5Q0HNTTOOkk7tUX415jmLrFJcU+PwnXGhi40rga+hZZ+lcxmsrsgiNZ
X0LOFJGNCAVx24gSLmvzEd0oYAnb7pYQ5olMWrYTv9m/EcmC+lFyj4MDH05PmeHE
suARiarnHJixU9rYLeDTQYsWs9LOxI4AM1Y4Jhl90VRDWjGQs82vF0ykvMEtYawK
XJOo/V+gpJDAzCuLFxv1fWgrLj1Lnw4S5Ig2mZ0fWqrje8SoWnISi3FV1kk67GnW
W6Neph/vHr5StczAw8dgCnc3ZWy0iM8HWrr1SG9dbfdUq63MCy8dq/8ENGeeVnw6
T9M59LTrB5akqt6r0gBA55yX/K73vD79femoH2PgcW+YFEXdE7HQlcp63kDseDm3
JXFAgAA+mQ/LBUHfTD4fcJPRRLYXx+nO69h/eh25VCcyMsgnZVQDMrsvsMsQ3rTL
jP+zFH+4ofIX9+4JPxRKKCOzAuV0HMRZaXLfoGjITYOP+12upCW2pBdRoD2jAduf
wKcqeKjs4ql3v4nYf5xYX4QPqP0hlyNA6A0t0MYCV98HBRgB3hx9+gEQm4vqvDaD
sXOEhSWgzAkr0FfwlBRoD7Zmv/c+X042no9BmddqrrTcTlZ7XJWuzrV3ymdzI00A
x3MTWG+5Dq3hxfDg3B6nrIKA/d7m0NLPu01F9lXleZYn+j68nx/2xV+Q4h5405PG
bmlg5hBbWjKYcpoHdp4ciX6yA8I+HHAGVIDJGbEmRNC+T1+U60IBnSLqWMuW6SvK
AzsMr8LXacqE2Et0/fZ1CCxhiF6u1I3GArhiCStsGE1nZ2gl18QjtGkGKtijWHmb
0mapV2AKjDqq4GT+QJTJnsvy1fsL+bwzJQg7IpzVcLcDcOKofFdA8YxsnybcPKNu
U8pQtQzLD9uQIhza246uf2ZsQ+sC6pR7rWo5Z4Bfy4DQ9lszc+KHba2sYGtFT6WW
26J6prJpsqiFpXjb4RNTsuTCoztBlaca3+o9tj9tKB6jRfDrWbu7rfDqEFURkC1C
YzgpitMWLG3rhSTXZOJ4Bqz8vHBekVs0amYRxFsHi/p1Bey69xzz2AEbXRjIAc4m
46x2jL9Bqc6lsE+doPAqo3hEgW+V2jPBb6LpB8rcRHv6NkXK+peowoLE01DLVoRR
iukpCwBNHLVSzUvHx1P8GazCem8Esr1a5M1YGp5E1V/tpYn3AnDMiQfpWiAi0iMm
2Tcl8bzyS/+90dLaVBy/Br4wQw7lPG78zjpCr4c1dzimDoG4wgIlXIyNI3ar3u58
HaU/v4ScmsB+kqt2z4Qo1MAnqlP9bnN6AHkFdFYaGKeNfGaCJN088ST7loHe5GV7
0mVCLbSZ85L8qGOlGujaEfgxTd0J3spN/EUo+HQ+31bBagMOqaY1ZvPDd1cAI7Ln
GgbrY9IrGgJkncWtg25YC191yvZy7yEGOAh9KBdPqvbpbJfky5oHROIuDRnmI30j
+0G9UM35PdpBrCj2BpzbNUuhtqYwgJPxTcOoySxFznoHrN8exCCBevj5dRZxF1ut
TbYY3fjgzTco6YOYP79GjZEeeyuV6yFb2c7XMCs72pKo5bUALtAHC+SkqgEBtjET
lkhYWe8a54Y2a9WPxoOGXIBkVIkRvT+7jmoELNmjWPp+qGQ4ghJWnX2h4lKXfsYf
cThph30TyEmKphWuRYF2ENlw1trtMAkqWqQ1wEtGmux//Yc2vcK9a7Eab76vJdUA
rod6UtwoJrS11k1BwoM/wqv1PLvTQOPKtXYiM/H8uFx2x1dQ5U6eVfEqDfLg3C2n
LF8/KRNuftBJdaQQbE1NQeBMVbd/nSilQ3z+ou5qXhwGbQlXwauxeZPqpP3Ea5fX
a3uwydF1uj5QM8itqkjup0iPVN0Lmc+36ZNj6CDMLWLj57eNrGdpvXrwcyTv0bJv
WTBTynwkHvdnumXt67hbt/TnAO14+mjom+/B89Bq4JEDUEhRKNTM7Ny2+RMHVv/H
YKIkImnH2aWH3DGa4B9fwc2P4CIPVs5NagNGM3qH+0VBYVlQ/dx/R9rrD6gFh54H
g87vXvx7tvY+HDAJrjfxahR5xP5c2Waz+f9ElVg7zOhXPfLl54XE3zo0kNTaurW9
afkFpBEAmysbSqsSLgfUWXmHxf/7dT/dRC7nlByLcx//7FGWi6vuo8xcp8NxkWRw
2WpUtmBPl1blaJjxNNST/oZOwupAptRomiwhBvxnuNHvbzUaxR163jg4M/2WfclS
a9q5Gmqz5nA8NkLSJonRj5+CsspMWfwgnqtIxYi1XQdzDskH+MNHqs9QKwgy2HeV
mmPD47Obf2dCJ6kJUjoj1x6TYxt5m1lWGNODxI1nje3eGzjdz51WyhDQYmrBt/Ih
m0q7A1F1+calYu2Jp34x2kf/5lvWB+dPug/Uc0OZX5eG3zNR+NXNDcWM7vfDoC3f
yl+ZQNM2PxHu1Kdnmaw6UKm6NNv03skSIv6gkxeH1paRoAjHBPDzz81PPUzsH55O
GPFTwqUrfiTi6Rmggv/BsIeoLNpOSRyCJpCgJjazdE6mqqJLjOBi3atVte6hfFME
fcJXpsRE2Sgv+4MenAamWkQYVL6UYik1+moDyb5T4FUYQyM0gjdXtJzfNUlAFyYZ
sI62SsxcDlO++4Zrsng41F6qbveMK8LKCD3gDiB6iVd3Wuv6TBzjfVbHMw0t7oRm
+hnwPHPDo1jEMItOcirZdF6FzSTV7unLXWEb7Ee0JJl2QE4hj+KXFCdw0+G8/9DY
zN80Go0e2+CqFhCL9Y376EvBp3XuOp3RZzQRhQjSd3xoDZbHxuj8uSYTVULmXKxv
a5u3SVRGna+5Q0gGWsL9peJF7Lc9/LTTqEkk3kiu75SwQXYTzx7SDyki3TTvvHUN
IBxypxOSQzKk8GTwXK/sYYPPsddGblzxWpAMwn8Y3bUUq/bfaOl7RY8hbsK6De2v
leDlXD9ElF2WdX6V6eIWM9arUWQwpOZbW2bDiEcVHMjFuN0TOWv7k4anUtH/FjlF
CyNfAwYZEZeZaYH1Wo8WXx1EKe6/qiQOwjufleLEBXNnn/oVVD2Z+qgPT0hG13gz
EFnvsQkXOOmmM/EpQEKfkqEdVFDHR7plilrAyyQzrvNj16FmubnltEnQqiGVj4+R
kxxkwBL8XJGAuhRrVKq2rmzSXQsYHNa1UhhsK3wMtquaU6RKsoxpuOIJOil0NFCH
DLdTxlr+FyUIcx91zzgv83erj3IDfQ97n/NblrZhary4PQvlpmqOPwL62SFtj0jn
vfkodObDkrHvYaJSEoRsXHMVNqnBbwbfw41PXz8fIAfrrfYgFfpc/qicP+lH1HQj
hUW+mFnbd6D1X0v4aCaGEXYfER5XavDQNFTwTJMMnlrhbGkAdtbJr+7innpBnCyG
1IzXH59146rwL9l1M1hX0SAXoee3soNMb5arr+/477wMWsYO/rrAceL0it4bWVir
7DbQ89jWKmVMjRoQYtofDj1dEtO6m/HlSKFPicwWYwqDKZA/rMctHg9ViRvoU1M8
JF6S3kX9dSj4LKgeDwojqvM2b2bXXfSd2X49DJcJzCkQGj2qkB+2fYIWddM9NqpW
mFbg9feZtWhru3H9Bjggn5hVnad3zy3tUkNF8Pr2t+M+tPRK82IoVBT2luVfPa3a
uPsZXHnVkySOfO6ZP/mNF2kFtK6IxamMTgHXUsrJ3agcJelvFyZLetudm1eVGpOX
1Uy67noUS6AAMKzAEt8DGjJPXH3MDGdbZ9OV5De+JGbkg+EMNnZjZfc6+inKcaGO
VIcSaoW5yY1ChFacOsU4EMSgy95I8raA92nNMim8wL++ETKoLBkKfRXrLB0O3uJi
cantORIg/4Ou9NO/hERcOtGORteOm6mh6sBgvKI6PZUFE0HKQ/4spYrjO3Ou2Mv5
5HC3rWeJ8Gap37EMRgK+ujyQUM2gyn/SjU9kkOJx3MtPr/eLgOyAoYGA4xtwe9IJ
DNrhzmq6nF6c4DTWLigBDDOtueclB+qU7Y6gvHgWoZo5mr9ClGLFuyaMDC1WOshT
5LgSAR3GR4W94EJuUU83C0zinzc6m3JgMYbSXbcj3etrwOY0vxYR18O447VAEhgz
MxA3e5Mv7Uk7hO92BXecEcgJMBPHNc04I9kiN5lt4pndMUfaCZAmAlAqEsvaJD+N
o0yY3MC3EtdRJgHozpnotXAKTmbXOctQgDM8ayR/VPUzb7MrZpThVS7D3LUaogt3
Hf25rOq7GyN9t72X7I/38tCZdH1wG6maN1iZyxQUKBlb6RnfuCxrWbNx+JM7wr7/
VoUfLfmDxwtgI8uek8iDqFBWCaThAi5F3bnU+DCrDTTaPLIVknCQ5fSwXH40Yl3y
CyMpkn/H69zqvw/RxmyjsrcdPh7Gv3LI26jt2Szmohlnpr6rZXL5NODcsOOFuhg/
NWDejw0YvolZWz9KiHnnlPoFImVqy0dIgT52dQFVB8TXxzYyJ30zbfVzkjnKBhNf
ilbIeKDI6RwX9k1jyRAdIOWLpXRh116jUQ2uVNvYko1LrrNBujfdIy9w8JcTRFF8
ehLnj0b35W78fjoAeW/tkKxvIngASJDkHdMmrIy9IWlRYwASy5QF8Ze9Yqk7dtnJ
gqAfeHz1PfkFe8HJdwK8F1Ggd5hHvFQkaCVXi/AENPbYmONqIroEbv1bDh0Jh00Q
hlSAWl42E9RR/uzdNu12rSkFqB8asHLE57NDqoKCfpWm4NZ3+GJU+ldbuXbQf0EW
GzOD6Et44AXoKR2wV7Lf79Np+zQUwix5aYmGy8iTR18vFxPdmold8Ht0b6HmQJA1
v8qeiLoK7+wWaS0Ah4Z4/WtGXki5Nc3CaXOfM8eYF2NeYUr9z6q1KWWRurB+oGUf
1tUG9bGN8uLVsc9gtmwpK/JobljC+fKUl98esXJ9EvhOvAy/2SxpjTcvNV88lfZx
MdZBVqswdHLpBdekkjbizL0yfVlxJ8fia4PwKvTJDBHaedE33Dd98H9p6x/BooZM
LHEOY3e8R0x+UAMGsj34f+ZROXbHuiYNh7S58NNHYILUBpFQhnkzrRYoFmpdjs/Y
ptHoo/Zfx15vyJPQNp/scFHCeZuT70YjM4vgKRduv/mZlwnwZqdzfs0sPyjJ3kjx
dP5XSxqbg9WVAUZelL3GxWNY629rdeRzi34Ah2gvPFwGx6nDJKd8Z2Lxrvsnn+NE
ap1RxWxmEN2KPghqZ0exnma/uo2wx5kSdx6t0YJCk1gU37+R8BwGLjutsBmWgwIQ
9M0GrortI7I88/M+TECYk1HxKwdNz5ybY+q7PMkVpANVQJwSFHLpuTB3uOTVHg+X
m4n+WmDXKq0Jmk4KMLr5BqRF08ZJa5V2yGUHRkjcRnaiGExwrAPj3ZBlxLXfW0KO
dLObc66pI8d5s4gAGed+odxS3x3Dna1GOxox1/BbZiyukOaZCtbuEXrBKniSMSJb
cDVYxov9FfJbMCnSTtF/ZtWt7Tf2uPdVdQpS61VNUtTrkzyoSVJZV1S4it8m3u/m
w5f8waqv1SU4EQpI6rqB14MWicDNK1N2otdIKAMc3xKmWPUudzKWCffdPOjxMMQ2
3H6QP9G9IW7IOpBoWeJnGer5Ndgtcbn1XAfHIAkNCHRh6OSPwoseql/WEHjr12Cf
zuj6lq9zZzxPuDXxyFCDS9XkamoWqkLcPhS6+v2iHSt19LpA1Iqu/VzM9Cvq5yqi
gt13H2jWwu5HWlNDqThHoV5qyBHGZons/M2R0F6f2hc+WsC8Z0db/hboVMmuaAAI
urf66fiOr0lMsF+cMErmoTmvPRvC0PZ8SBruynw0PaC4U8uCfLl+Q+w/yfNqKFN6
6kARXH+r/BJBFhBEJD9cWXoddF8zn5fthinBIfcgVk9FwcVsixZPWFkuaK5h3VTJ
TTJ7KmD4xVrI7HM9S4/Oxlj5t5VfMc4bW6MEkkMEJrcqAvrKMlE6mXSEFul5Wc/a
bxFUJUXGBX82l9FjupR1hmyd1w4Aw0KQRjp0GdkYtWCh0fKC2iiXFjtylADn9qbo
qkLgfqIljmk/ORwWa1NUhb0mVmyW4KFpsFAI3RvSViO1Jic25kIHD6dXtw384vPy
rv9Ili5oNJHSSryvtMIe/VQqh+/K6DcQJRjgBXyKf0Y3yFE2Ozwz50OZbXKKBlWf
yJfm4ra/KHPIajplVIFqZIMPFldSJC3wM6zGhZoPUKkB6r7+cpDOE52Ovh3vbdRM
IC7lVTg2HTVoe8QNtM7mPSfx+QzBeRCd5gV0s1aVv0Sg7Ft2vcJWJJlaKx8FX7UR
D9JF3CdmLiIxwivOf/pNl7Keg5cIxfMctHxq9UlbaUSdYu/+Tqbc9nCyEEnPUVwA
9uvGdo7PRkbUPgn21b+mYeBPheE9XXfHBlPb9i2/8zCOCLp+vzwQaHVBVWdbSADl
UAiGoJGSoi+KIZL8oX3UZC/WzRxgKeLXQUFRxPztIybZN4gl9jKPkV346EmEM1Un
lAJ/WE6rmGHc8/yaEachjq4zZRpKOtwNeggnLC+sW2vJ5ILfVZpr4KD13ClX5v8f
ZEOAkucKon7BSRnR8wj2+77y7UXLhdUq/g3qDmmrznbr4DRULqOSTxRmF37YJUt5
hkvsUuotp0IGvqrzcAmgRe6IgAR4M9Fhck0h5Te5Eu5cPXnfsBaPfbVCrwXkpgUr
kle+uDCZgn9IqZ2w0HUZPS8C9IaAX5eD/A7tu+zInDBhtBJl6VjqPvMm0lLEw2VR
nsj/sC1k/L9UdetgW1iZWtVmgbxjZxGfy9QG7Mlvx1v/TdENpbhaKN/30MC/Kbnx
5c5Dt3+Evp2lqRZzB9GCIJGTg1Byg/bS3Mh6faju2GN0ZjmAauoFKZrwysXgPlDm
a59itT+05hvSZNonA5p6XR5tKLWDM4hl6V394TDPKfzWXXlPxb4Cfkw3jSvPej5J
Yi/UmBr6CYz9JWtgI31Lrj7LtxUDiaX6kc6Bu5AjFYfoaL/fEm3hLrsa5nxz6JvB
ZqEbBTsQSbjykMsvTzR7lM+aITXyEN5dXj+/X6bZwZQdI/qmcEYJzrgRe46Uiw7+
Pg2SPV5Xn6An5J8lAmBT6fb2IdgfE4v5wcTfQW9O++UZQT/oTvRe26rvePHl5X8f
BL6GpzLcaTrktxj0uQPwrHnjIFt0bP/7OCeCtJ6ctRFqqvC0IeI6vTird7b6QeRs
zpnZJ+xff2ZQ+ohBwXu3UUtYSjLVwlKSlaq9qQcOQqG2zoC2acYkpFXD2Ch+xVzi
F+MJGLpk0pIWMINuy+xWx8jxktFrdwLvrjyC97QqSNR8q3DxPce1OHnCnSlr+9Yf
Xm4O6Chnw7HxJkj45hZz6wYKpoxN89+NAOdviDlcQbhNlBvt6cQw3+mvQKLqYuTe
pXVKIq4eO64CQstVOsA/jwkm/LSTP4BYmrdIil5QNXO+gph5/ZON7gF+mKWPpADA
m9RNYSP3sjeUtrIVfDwPKnxhEL/riJkVhYzhs3GVZnBGEzvXNuFghof38HP42W75
8Dm6dptkfePbv0z/+KI+OT4lKOn7VyBEAOaoKUq+92q4eJFXvYDxl40xKXuznl6h
cTpmtyR0ikuHzcxnxRf61xFUWlXpfoDnASfw3wvZu+vh/C9esIXeK4R1Efp/uNQV
5FIs5RICF4ym+oZ/jL+hq421oxIvVbTNgLHqBJZ+L9q/Zo2bLj0o3FBrX9z72TUC
1Cb+w5yN7/RoHGy1noBZth/vF0lV1RzL2smqdKdv19kOnkxjIr4ggac+BRZua7Tx
H2FyyPHo4he7uyG3jC+GMWmfIfG4/6cX9Gjl2J/TiNfckKL0zRs7kQyEPHJ16DMQ
nx0J408n6/utkoO+1wyZcJ1uOwo/IUJ4TiJM633TZslqruQSOgRrEoXJNdk60q/R
QF2pAgx9qaoPMADJWltZbJzZMVRLbXQOtgw4lh6rK8tnTK73TO7zYyyzb4+bgCHD
G73W35+pSB/bPrIk3CkN2rUxmhgTPffz9WFHylf8F+eXhZOXZ0mDPrjt3wX8xxpE
lX2j6otw8H0Ves6EhgreR//EbVkPIWBcHPRFQa2g3lnpj5dbl9Al8WiNINTTYwWI
5IDccQSu1aOd8KSzPE4ZscvKzkGXPit2Kj2Q6g5Tt9BYrSaBSrKho46uZ0BNz8gr
AgsezfSxJEZE2Kx85CjN3+55a/akCtx75V0lYnZJOZ23K0pAA57N7254CYUOMaZK
wHFUw5S4m1fFinqM5g+1wfqscGEKiLUSyJYRCX9Ri5UEurM0yK8NOpku4JcxKwXT
uS6T9zgDmLQuxbYZ0SLsvV3IZ3lrOxBtEyZJEb99rOVe8L572PXzbG1M1HwUn+Hv
cFbYdiBEmW9clMjebpadDkz+kQ/P9gqKOBDjH+3Aoi9T2IHcOcZDJkCC+ot2OLOn
DchCi+jfeqfrvVjr9rIknNZkSrbK9uPEl1cUVb+zcuMuYGQ0NCh6PB2HOlOAOGCf
qgCv8c8eCcVXkHl6z1IVHLh7rf4GZLQ5HrRu7JxDj9sIy4Z8PY9HDOhtIp11/aZG
qdDr4gUgh8E2Iq88RuVhWtfIpLWbb88+JoWjy8TnQuMNYdiy5bF/mBNzr3oXcHn7
523UJf+svXKJkrh8VU/N6BDkGnzs2XlXkmded5Imxn2DN1U9dQOKKcj9Pfa6JnUJ
UAGSvtzCVCuQzfXSnRv5vLRS/CFy6/gGhvS2JD+onYh5iBJ/Oo28MWPV51rHpxhF
gwWHBkA3zX+4vq3C1QobQeSlWkIKkWMNpBOsK2yk4JTaGK7TLvsrhlb0hh9vn8FY
SaWnG1fhUZAiImFSRkPO3utIQYJOx/0WFdzj2D0M4JqDaDtT1nh86C2w7juBhVG8
NumZY+fHZDr+26x6LBmYqqCus2L70TLuA/OGgSw+AZ5bxlLNZUvZDs/Xr2C6NtlN
Ko6Z+z1OU9fVv2Q+FQ/4CSWKs5q/VlJ56P3gxEJGH6BUM5uU9/7GRhOis8tgHlp/
Kvx63gE1fXeZAlel7+T6W/nsBG3Ydtw8z5FAvrtZ5cdxg8Mu6PZE7OkxnGw8xMP5
f5C8N1NWFZyYbLp4jVv2/ca9VDAweiwmAdD05HtZi2mmg0NhcGWJh4g0QCufUvIJ
CcfBL4mK8e5XxZILfRZi6r4vYENvrBEyZnreGlOwbMk0Bh8yDFtZ7P0rlc51nwAY
TyEqZTLeLSLDwueGB3pLq9nLdG0JsNy45DwqDjyW8H9SuX2HFtBF6axO2hPE6wDj
LwebsyFVrJotGBbCWdw8aZGEYJHX2ZCSPjMlBnWYHfxFo3ie0G4fUO6eEgXmCbvo
famNbGOrdm454ijdC5AteaQ/apILej9s5C6XRZXlbfO/+fJwDulu2Os2crfcGnTy
Si2o51mhn2M9r6gx6Y9+8PTJZ19RcFo43G+NcKONKSHc5Yt+p5+yq+6/ymQ/NZFi
Or+ZLLjKdaXzopeOReVP7f89U3syzjUNYpmLDGG+ftrXr9GHzh+a85D0qMXJf6Ee
r5itRVnSnL9UZ9LSDjqmwvu124ajQQt/SIOc+kFj3m6a0M/1B0qqyeXUnoEkfCT8
twhUOIOvQ1E63uZ6JunovhXa9ekC+crgWC+9hUgjz5LHZbWreM6lQPdgzBN5FOFr
KSl1j6saz45+2DIcHRLL5GFc10cz4iuSPsyJihZ6gkBnKzSD+ZAwS9n2bYeXNqvm
nqjgFDQ/2FPrKmyeE1rCg4L/z1ds3I+qlB1EovIJFhpBLs6W360YgAqhfik4ewRp
S2rRBuxyBVo5m6S1QIigMOR/OVOR/x4TvRKGIWhYL0QHE4bM/nx9vALKjKYpzoxl
XxmWJNWFVCy6ZdwFl8lT313Phci5AdvRUm9QczzRzA+o8bjaRaLkH/AIeYHjkwhg
pwtB6UVAenFfDLMCXkNXpXXQGdBU0ObVeGYxA/elLQKXCwvOfeX5rNyeC8e1gz0y
cHEbLApR2pJxhSMZchOukSWlEFQi3Y517b/VzKMoXUaStjontXyOBMN1AMCUsoMV
fMjEVsosbFUcl47e8Lfw3NN12k5GlNBmBAm9ifwnDEm585hrBilZW71t4N+/86WJ
2wQHVuDhJ3oDg4+QqfybS4JcTE8LzR+l7KCy9WEmOWfqNyYW2nzQJqDa8bson498
w6qBn/2dEprctXYNIfStZMSMflVDDyyRkdDCUjb2KR+W/C+N5yrAMxAjmIPRHB4N
BHcjg7NWMfLarQetF7xms5RHEj8x4+CP1/+APN6nPHkbWlGGLDzT2Bv0+XbrI/H2
CEBK57QGMYskXGoQXmXXlDWfClpbYxUVzvXSOIRTYRlsAaNklmPZZ3LJZDGQk/nU
2OacUFw7Gf7PycDX6vi0thtRCraErUOPS2GBT2dRzGnEszPfk95hoycpGAUUm3nM
b/KiUk4qjgjozKQVGysmImD1+0DxZaTcXXtDYL/1fRE6ESY5/OLAJqrzd0az3BmY
G+xhdiYyVoKWDN+tZRKsxYbNYtnpZj+UuNgbAgmOr9rGkyzA+FY39XQuUOxmcoY1
+usLDg9YCm62Awxxc/VNTVyiYSUd0XJBU1ZEaPC6UfL9k/1ZRrB2Y0sjLACHPWjb
Tb2Jgw6wv372da7HTVVSIzVHh5xWIoPIMFHLtFMt0CVWt7wtTRvkzup4Nv3A/MRI
+aMNc41uFgwfoKwzZo/QgnnS7Othzg0oKLBUL9GT9pNnFzwfCVQZkmiiOtzCbphS
tVPHCgQrVTJBte8qJJ8rnUkCLndxdcxSnGm5BQZhrycOhei2KXafdonQ7hWZjZ5I
XYOR2NrRny0IC13fcnEtJycXfws1tGM7P2q4uJMzzF5QVTQ8Hir1Lf3poQzviXIR
jPwwdEir6cG0wTnUVQSyTX+30d2+WwPHLsbnKsdFvD8uoEeFRZlHG1fty2HDfQN4
uTKg8ujZ4CMCc4mOFtfbvbO3r+bLVk8aNooNo1OriNYpujvkyGwSgIg8IDGcQhrf
e+wA1Nq8pxhmHGyhfewQF0AZqRTpE3/IcCqOwolrIUkhiUmplatOvKDeMzh0WkcV
zdf4Mv7WXiBbmzT7ZwmhEio5RwGE/alrvm7jdyom0ho0eSzuiqXrpRofXLQFS2LU
Y+9RZE+qtNo+unROwAi3u30DdhxbSpw24BaNDMnPEqsV/89+5Z54qHUWH8cTpvVG
2xYsgPxX+VRLqFaytReD0JSmlpodzrFpnynoTQhANNf5TROaYvJGmYSOThLrCHby
bpLYxbMBPLm7k1dbJ13Wrj5oHnLC5tsK201TVIjDPkIHgNxMZo3J/QHWcme8Io4I
QDo0FTUEMiJB8uO3j2ANlfpuXMr2iGjBrc30lCS/94shTPWFUyzeSLAR0pHfgsfD
EFNDjgLc8GKEcLbm5evgCbIkHN1a3zGwQEaO+CE3/mYyEreosMxUoG5gd2vsDnkH
x84ATJtWowXzpZndGSKMZOGSkHinEg/G+4udQrP/iD1DIrDbaKY8rPjYpNtg3P4L
6P48nEuluirieUmLh32AqgRzrfurGRnAhG4IOUj5ZGQ8jIEU9hZ4FVST7qVY1nsE
r+AyeyOPj8BQ/aZgvg7a6oUSzQROJzUrI6aDTJ/uMz+28fjklTeAoTkktPe4kpdR
5vXH0D/9Wz70NgcPham2q4Aq5DpikSPa35cVNk7JZYFUF1DU5qrok64RG3jnlx8+
CdlRbDQ9a9tqZ2fER20crup6RpqVuK9FTfkppW/vExLAL0YphwZXYqAz/HXm3Dw6
0RBnm/qQcd08gPlsLIy6HSvLrIN07pKnoUv+KIahqEaqWEylb2ue/qcRREV6hNnp
QsmBwD2e7fSjXy10Z+sNiflJ9z/UrzyStKBC/XBihSYNLlP53h2vC3J0RZ1xhUhU
bYtADBJwcXb7Dd84akrxdwT16y+vA4/l2/NsJapvb5d5B3ekQya0OYes+350+J1H
tkGCH+UC3f1biYkAXcruG0bykIV4yfUhM1HZy1EtOqT6aCjHDgLh8BROMZneuJZk
+xyiMPxS4SkSBtcuECX+SVrW5AQEdYNpI1gfn6F7VJaJSvRfnb9BpcArVh04P8je
bF2VvTWkjFLeiDOR/eEe2B1SgfOGj1cTvZuq+y6JDuwDj30Xa+GnvZ210V2C6ele
dtwDzZwrO4AwSx/0rsE8mdsOO1XGT6e55bpMX8rRb3XROQ/QfEL3ivj2I6xP4ybf
9h3tB3uTu3CCy1o97N1HU4VHxWsyCKpeTdAiYM9tCxMjAtwSMdv67GGBiZrLzWA/
4IwsYKDbbVu5GkHkDA4kz1zJQ/mpSN03D/SaOnpSMzxxFe0RADqfA8pAsGIFngSB
hYveBJXmT5BkHwRIVaj3g67YBXUmWGFbwSU/UlIswIuzm4KIEns8Hs72sSqc/Jpc
pCH2MC7tAHPCi78mOTsm7m9RNffyIELv2Tyiwk1mkP9mL40w6LTti7SfluoNaxiP
GCXvwFL9nwMk4TM6OBCGWRoAiX22yV9N8Ws7OCROyJ0iI7gcKKSdU+czEfwOiMJe
54AmcPQwQDgk1KMRIYme0m8Z4lY/olhwjlgTXLmmjqkd1zeQkqX4tlL2K3a0tCYM
CcPXUWaumhPBKwZ9cYIIuCfZs4sv0DjREUTnpF5acxVbbQMKFsm9cASDU0gVrLzG
k3l8dq3n2PpyUIds66SCvk6jydWb6d1F6WX/axLxUm8Qc4cwYtNq9MMheHQTFn3N
cP3RC2UnqbSjXhhQ33colUP6sC5+IiC2oml+rclMX+/Lk6zlRyDIo3HCs9SdxiNy
zE4x8+E3orsVup4S4lFlbFzj4NTgv2mXvbPKsedQbsQO5YwHC6X7UXiSfhRP0fxg
FfzpobsUdI+6vXmltWw9qCKW17gnHfGP4giuTW5uwsc8zPMYck6k6BuIQkSe5pTh
ynsOitcw+stPp1SpLV94u60aicptc7K1lgQKlywZ9avFz350NaqzrURar2H9nMRM
PnjhiQzU2UDMrTEXL7EacDfNOCQuNsstwDaqNJRyLho8gAiPEMyS8PYAJIXWvDm8
sWNE7MHj1zbYLkIQfamTswlOIZg0hsG6iXOqcVyH+9jZ5wcTkrvOH4a/uwAQq3N/
gjP29Ktr5QMlQhLFG9wrg80gWgbA/JbcMSkx7Qmhtc3GZm9hF32vOVHzaL4PxWP3
y1R82J30nzOmlm3t3uKiNsmr2zx+83WWN0gYliifDK8ZQm+Ii5x22ANQLohP8yqs
DsH246S+LpN5AFseAfCJCcdn/I5vgyNhsDM+nWkKCbPcbAKP6UEFNfa66YtHTL0b
tbAwqK4k9s3jO0BwmJUjXDDNCWWcNvcM7fVCVy641KGvUgCYWYkPDA+ScvLEx2jT
yp9VW28GeavF0cfj+owSZVsy/JAvPPvIwhTH1I83EBSZiUncFKN+i4APNjRfEKUE
9tgkj12cpEQqZYdT8gmg/+pgjOwQlgyyhqPwM54qtOfzfpar3XgmlKNa6XwWp2eZ
7vW4xaZUZiYCPn4zZHZRO3n9cEL0ld8AbcLoTpQNshO9qmyswekQb6ZlYBUyCvq+
RbvoXZZnfsjg9m9T4P6cWbiPZtJjDUPuU+Ha9n7EIIQZcYPgODmd2n819GsYxHwG
8Ew5usoBz9RFqd4n92NXETiI0k9MrcW/FUWrHDigUXD/eXiqrpNI0/BlzUsrfwZc
9/JkrbAy0c704SP/AhOVbGOKHYKgzVoB4PvFmPT6HfXxasjQ42DH54FqS1I2eX3t
XRdJ/S1BbLdmrIyv5MLXAKoaF2ewCdSk7MNKVCvvAR2fxtDOVDfyibybjKOebaDa
FcN0EwbChtHKMKZrpmWABafLOZcBxP34GJL6xpZRICD88nqqybRAdzteK7qIe7aA
u0+OsER2cNSTTBLnmahD2znsoCfubVJGp4kKn6epiqGJzdRVCZgRaMj/g7OglnIo
8IzeAOUU1n2AsLRUnltq6AeRNwt96L/FUIQQO/B/6XlUxiAH12M18+RWqq/YFZ+J
hUzX0F63Es8mLQIuLYiBu6n+x1IXbg37nTNB0FZ6KWyIdxVawchEgC3OEo3ht9rG
y7t7znn+RUXMmeSE3aFGJe0kA1jNwzzMq7PNbcJGCC2bSmlo3zkhf9ckJggekJyJ
ODNRm8nbR1FCfqO05ytPKrRVJL88sgifwuZY3EVIldfJ11ghOIfuFmgARwWTaWz+
xKaRo6W5F9n/tP/kmEmP93V8aEYNYEBw7u95N3+d+wtiIJzN2G0e/FBLzddW6Nkr
0+kCJx/Px+CmZYNfFzGcZMCYSUHeIyqvT4SYiv9eHQ3dGXPxtL8zhXXXdepl4xI9
hSlvGK2vy22+juHKSvlKbH8lo70lvdTmcHW3CGO6fG1/Bd+4+pgpXRmDjMrjrqmi
jg2D8PG6xYhEQI2/HIRRFpiGPtbyUQ73Cis5QAAtVNwyme+FIDZ27jtSV9Cuqdld
sEikL4KawmLGecs17tX6pKC7IvQw8tHE4oBa6kuBnXjCdkQPSlFmyzC64KdAUc5V
7qo6N3TWrAfcRBuvMLn342r/dn2tnV4RFx7/tfd76IoYY2fO7VtAL3cbLcxepTnK
JYZi0rV1QkPqA76NlvLA1jdUeH/Llk5o4ttvot7BEoawyQasUhLIF2Qnqo/CsVoc
lG9HMspivBiI+yfyIX+j51ISj/6C2bnE9da7f1V3CVbjNVTZFlEcpPQobssybFUz
fsrbeKNxvp4/XrhZDhJ1HeD5ClrJ0KgPqtGnCSSYTw6GYOi1DEXRSNd1WBpabKAf
f30MKZ56RzCGLFu3YbqNp8uOGTYrjsQLpt2ZIC1etNTyKH3seHnLMM8SqvHGgcpv
Wm0VYRR/QzT9lrx4l0YIyFOXwvKb6appzNCQMdeelYL+7LyV7vMqkehHfj8yjDKD
fLSRtj2Kx46tpqfAS6V27N9GS+JNTjB0EuTR0+kQoYcqXno7gf5wVmhVtMTlGLps
ikfk0hdUU2RmvxOnhvkNnVLJiL0PjxvIrr0O07RWYf4ENMNFFtGiPhxN37GvSnki
KDHB0xeW8OCn67HY9pL2o+vMPi/Oyyge8NgNMMTzSoBFUyX0V9OXUmHM6DLPcSDp
fXJOekstis34nH5BcZGM1SuP7QFlNTgd3Z8yN+kWuFMKspUKC6CCqtlqS0APV+eC
uhx5Bfas05GU+b+Wx82O+iGriO7+ScY+dySQ+E1VungY++8hB5CVZSiWdBU1LKTi
n4edLhXqcxid4ldkBGZUQUlPtniX6b/1NluWgL/daJkPveWcPCFN3ypmAajmdKeK
T+gDEm4BNsZ0Vbb6xy6+fMRpsdvBB75dxQg9N+XssLUfZi6n8TxQBaxfdq0ZFsYm
I2/jqnLoc5r3HgE93kVhQSzn7/xIut5czHIaksgXCpYT1pOw+LMP81tQQSLuxet7
FIIStfcD9tbCN3j3+D+HiIo0kAeceCVGXpOchjtKXZgt38IzsUDwuOg709/Yygst
93G/jGFOCVYwQLivW4GoMxTK460Qym1kqut3FezLqlBEqeXFfiZnx+jbRwmd0uUn
DTK1N7WqWjKzRqCiDtTWMSPFb5A7mmBYHuyPpEnZia9fCw23xsEs901B9S5G4j36
YOogphnL7omDtwGmZVZ7+IKr4v2iK+fnqY00acMIucFPWD3BVoJjGi20MFbVvUG1
TapElxfyIWPro9P9Y1qErcB2z+J+ldAhkrpeVFTAYMEODBmfk+ubJOxkZV53Adyn
vv8fCYHehK8T5tvDo5xa+CTp6sA+UVE0IQ4/T/4UraUSq/HYSNIt/azIfTUg+IXI
b1Pe835PE1kA5vOT8NsoXo70dgUulaw3lfSy8lWuNErjj95y0K33DaxJSaJaMXO5
QOZVaX4tC23ydvsKNlBU9J0lzcUOTDS0gFVLgcjC7eBsqlExOwzpP5vsa3NFnkUd
62OZW8KlIG3vWnfspWGtzQMPm7XtWXerMLrvjge25tBoS0ilhRzSWHfH7VDWxUFC
1ZbDR/Cuv+HS/xYuX65RYyCEujmBZfolK1TrppJRzsJqvQXGt7LWTKDmPZ9PS8PF
bGj5f/C/4pn6MFs3Ww8pizBLQkLOx1grFTkIf3wYSi9VFNI6Ddk6iLtt/slG0NPD
lDA/cI17+GKzqtrdg5NK0/RXbutWUAlMxMY+Ferc3GcF1Ufk9hxRPmMQth2FeYoa
+lBx9ZGBAtkEuhDfwcpOfFHBAISDVVJK3TsDP35Uy68GOli5vxT9M9IeHmmjdR+H
JRX/CKVjLbpoCr4J2n7U4BFrX28ozuvSnJae6TzIVMUc5lxiy7gktb5BnzxJwbsa
rI4LXTG8mDzj47ubB+le3IxF1UFJM3tjUBrFfh417NBRBQCoxlXBvyflgYHAjMbT
ozJPFFh6A8k0PpR/g17aa35azqdrLbRyoObF/uY325/9Q3w8u3R3uQBBwa+U6cDQ
GZDMEcws8wvaJsOC7UGANJSScVeZkov0Mb/fnX3IJvsClBLtjaKvxqDhYiPi+Ymv
sjMAn7duhDFOShiSTKCtwM7dLRwFhr57PyV56nRIGUr9QFdj2VY71NpZr0/aEsw3
rc064LI6EcThhz61f7MqQbzj1MEYwk4LWalBDi50/lirgtK2aXC0GSzonDk+61Jc
Gn/+xboLjdeHyfRhTN7lhfPQsbdOMezwVtv7rmv+iwxgZWYqCxOL7q/W+kpFAAOP
gqNSNfKaRu4qnr5VVHYwvZRSQDchfFHfugJcyHqyhKSHFP10gZrP2dJD1jSlhZdi
3n352yf6ZriNDZp1j/Cwm9xEj75jbG8Pk6O3xweG+gwhEjK8nvs4ooMVfZmKtDBR
C93TdygF8ZwCumAK5tAtP7zunw0wBOgJeG5moetTqR915uPzbKTaxPd3S8VrA7iD
brRqDxaEE/MblWAGPVNZ+FJvQ9mcY+VrDR1FyyPrILotuzQmpeZ6/7JKF6X5IWBU
iuGhC+AvnZUr6XcAisw4135WIQwoX3YE19zQET7rIvEMlmmH4X26qLWUKlCiHEe9
79RfPI5odFnyJ0Lqlc7KIkS44Y+XX3Wdv67AJXoES/mYiiXfKXOh5C5wJ4k78vsP
lJqVjrleZRgxdp3ewj6vcgwfa6NzMIvuzxwpWhbVyKqVBRslV51w3mkhSWWjip95
otZE6ox8cMBw0y6f9sS0g66fX82Vxre26vubGy9Hz1JAo35qnj2K4Yiw9WeFZgVI
Ux7hDlp6G46GNv5zQi1ehdHQhGYLis8kLNo4jo0gDBDcMIJMszJq5h+MEMktKpWM
qBo+VCrPJJdleK93WgZUvUnBx7B+dGL62eUtXH/X1SC5ae2sPieDKUGuf0kb2fpj
mWpdQxzut7nMG2usCp567xRUz2d1WMlDfjslcok3kgLamrS/Aaqc8tyeFWkdPkua
4UgxFgFsXhLlQJnMIhLNRUZXl3qusYx+QbunP0Z4lmMHHnFaJ3+nNumj7gSSbZeh
OTbjYX4cSSceyfRa5LsFC8okK6Hyv2koyo6u7N6TqzT2S5IxchY4tLVEWcqnK7hb
maRtGL9ezge5hq/wjgqnIvjI9QQUPzYU+s1TyDsljqOfudiyAiPOevRl5RqWctuF
yN6ZTU1W7SJdNQh949FOEMpKGwAQI5LkG8WajDNJXdFF6s5tp3sj2Zdx4bD9cvlr
0fTOpfIqIjWvfQ8P00HX9ypdyXSTisHxkYW88j8w9D9Wlf7ltwL07I6zk1CzTNyI
AkWEdU595WEsMzswYI+nv4IFZkxzSE+1zn/cWuRKxqZ5vBymQYvfHAYg1Q0m+x+b
peWUr96aGcmTFCrWLpQdMAfQswh9i0iBPUXGEB0B4IF56WA8W7zr6jJeiWL/WRRx
gfzXNkkaH4QnjVdraoO/9G8pA8YzzRFM7nXVMyCjz+HypjVowMRhlCM5EBOlhN2x
sx069k2UWSg6iMvBgQufj/kvj+RtoFS59dSZVDbWEdK+c6rFMTQDZ0jftMoJShJf
wcn/HdQqug6EV3KoWNeL85YCjaIiHhx2ATKi/X8ygCOV8Ym6BMWDjutyyIKgoJB9
wYkqcBKY7vuTRcwT/vWU1/ueZvQhHGz9NowhlymhdZL9Q32l3KwDYscfRfxPDHhR
ZMjkN4U/dCSnTKXkSGtAq6xsTrjzxSTZXIKqTV3kIbVg8/G64yV7fnPhqdmro0p4
e5J6mcU6ub+clniSRUUkyf9JEHlH1bbfwfSauEryZM3qibkYOXC7sr502A1MLIgo
I//h6WivGqBQ8LrzBQTtnzWF04D7ba7fWNHwYHKK+LH6VfMW4/J1vS1gDjuFo8to
KEQcojNyfaz5BpkCcC8qEoj1UWljT+280aRWNVl7mqI5DGtgi5fSBqFW2GC7q5CX
PQ7jTR6jO5Io1Eq+lOWwb+F5NiLPqWF2IkxDscZTKoH+yEEagLPCXblwpl/GPagC
dQTA1XAnWwaZF17n/GuOic1TgXAFQNhdHEYR1dEhjsaO6g3GmuQi7s5FChyxI1oQ
Z+CzzJdZZ6xieykiKHarQoOeJKkdj0gg7mKF4NsH7rm8Xc0tzuqUjJedCm41jopx
G3fBcIrNj8WYWe5p/pIHxY6lCgrOZDfa7ZCNVq8od7E82sd5LHHy+MpWlnPjyHGW
KNnJ2jEVli6tL6esgMlcVOX+ko3Hd0k91QfZVb5QhSdpWD8BkPtk3WHcN9H5DwMt
DVdccMs0GxqWXgv/NqrdKrQgxs5hDcLrSck6kGdHJBuO9ZbeJ4+RHcvr6Lh1cw8B
DeiM/L/1jCdwzrE9SHrj6m7hoSYuA1UcH8UmXLtRl9iUWHD0St5aO8cSQrEP3ryp
7iJwo5JoejvOehC2n0hE0ThawpoTJwEEbki42mC5+xWGUpG5wIAJsBuPY7tKsbZY
B4bWVYIogBIx7rw/f09bXmP5/EG9lbYw7eRNi5vlsnWxZL2bf0TJbUQRps4mSTcl
8I51ExOB/QEFbljVdzYj4zJb/eoU9W8HRX8oitjngWUvyf6OUCaMlX2S57nlQYh0
HGbY6DklAgNztqA2pD8OiaM1az9SZYcMyPhmFiSNeQbD2ShschviGaWzj03q1oNj
KDXpw3lGZ7EMDt1eeYXbMvbMqsHRdyFm86xo6WHsVqA7aAVccVs7LZ44RiV5cDeD
avy/6F8EKJa+yJvAoi4tU6Y+6NjxwUwh1LqNDL6YIhBHwsqoTkFdwB2rLnNorQJr
gcFk03XkxAXsT0WZVHZmJel1W29tDIMIcE2/kRqmS76GaFXf3F5kjlpYWiH+ajxL
g4iUREvSfw2KwV36jpTL8UCuwJEL2bFYjf2E21JZOB5E22MPAghYryGL/9H0pQnM
ZzGBoHHHrSO+fBUBhQRrrfJyrFjwholkXErGOqUz1caEIB6Voni7HF9DjmOlhllv
0PRuCQxu842RMBMQtTWPejD/X81LjdGeyr4PEoew2Df5oSqPeDPkhPhbbXbroIGS
5oOa7o+G8WJ3EXVJPdbNIfO7SFTHdZ2JOnoHNg8V0YEWQb4oMi2J0WNiFUUT72q+
SZcDaqjJuxW7Teh7+Zhgqj8ct/olvpzAiNcB3EL/mZw82G+SgbNSix9oFQukXnXU
9qRpFyzQRN6F2Su4QHj3NUoenViG3eMhRBjEFdQBUa3WXw0ChzMufXu7ox9Ex+tP
vJqpIQ6bE773I3gCnyY34U1ohR8Z87q7DZ0mYaE6YBaRbpigGKp+8EJWZIVJM84R
/7Tj0BV3JjvPG0h8EuNAPUBISrMvQ4a3HrrHT6EBmllFvZuIKCjHifHoCCcI++bI
UQ4QflFr3C0QXHSS9eQ8wGVAIPQGjFVwravYTYF+qBdFONaoLlJgX7BkFnh1QKyD
2BZQwKSI02fO400P92EpwSmjPIekIiGrzLj0UsPx0SboRmEH6ZHZvdRMVuBILtmj
dvZ25kKOTvNl4lmq1OlMfGQfaagwInQ/CVuwBX4NGmracYmkoTTvgmvp1kW3oJSm
Kqol3OOHbnt+56XQEq5aKWaOCIcGPW0V4J++CemY5wDiB8fxRKVved7g9CCZExH4
Z1nYOGCgfrV0sDbPkDJhIHlWBOKls2smu8GLABnvnGB7x1ugRIeKU4FjAl2uI2kP
WQWkEt0oINCjoYKA5xBzvvy1HN/4ykiuXkU2Jj0Vsb79q9Zidsv5SEM8HUCyzK9k
+Bk22vmemxtJy8S4GU+bnGypC98/tqV90Y9LDABtmEw2OGMcGdXJ6aGVWRW6kQfb
4owz9l0w/36+wanYWDBSHurWoAoMzwi9LijadsltXtrcYYIlolC7/6sg9JtRRW8m
2JUT9M+ZLQSHfLg4SJh0IuIwQz8uiyjOO0NurpqihhNPqXwKDweA0hS2Z9lt2xg+
TQRazGrmHCFe0PF2PNFBMQIvwJLB6ZBYPvkcg2B2FUHykdMr06KSx4giY00IKd1j
srXRxl0EW1Rq2PBVKHMEZI8FUFFQ3ODHURKsnHDQIyGhrfpj9KHZWdEtzMHXTBuX
KkfAPNyyMKrEvw/aztG37B7QULcHHLi9V6cJHAG2uZteTjFLbdgGnSuLfeSbxTZH
IzExHwclHJkX6nreul5RjihMDI+TeXz30wQ1OrGmtQwnQk3sj1Mw3V6wfbgmm+SN
PFn6JPRZvnBU5ytuXrlre5nHUTVteU/QBF/y1luTANE5LNOa47IwOTrI7xsvoGcN
qOENJ71W4wULWu+i+gyuns1TC1Nlf++6g/OfAkvKJafRCETc97TT9D+3jGsPeF4c
Wx/b67Vt9IVD+fcPwyyHT+6adat/C6FxymMzDnoFOmcoL+M1OjcZkm7ilmMaN7Oj
S6entXZ4ObfErBYqJ0o9a2AJgvQo8FDVQMptmfvB7bwZQgHnkmrkWbLQbGZGvNRj
EsABy1fzUYVBZdtCE63bmJuvqbPfaIisS7r6h2taGWf9rZMIZJ2aJFYDoUEEUOK7
7xzBPM1dEutgpHUNNZmpu1/kGW6AHbBhxI6DgFj/x8DBD+czxBLDBfA96YgRJOKu
aYW78hkzhjLEtBpoCJlGvH41EFEuoEt4ybFhHjr7ZaUhkfKrL49d2jOQQ2guwZbm
qn98fWbTJrCoLOWHJVsj++7kEzH+huBgA9sbCnstyvbzyYjZtep5lC/eZcrWaPbt
ZRNBzhcBvMzu0W0yKaP/ZOamyWicSM9oKWFkjsyGU81TYw129wg0MGOtVz50wsI4
vy8aHjHXxWg6XHNGKhTK9x9jEFsp7LKhzNV4fchpZmpVbv6NLdoOq8ntnqKYDf1S
dJFZogtfs0DXGrhciyqYqJG0JjFFQ02wG+R4WvbZ1MHPEsQOdpwE1ilJV6cxcWHG
PXm6c60oYADeyPOzc3HtsygRz1lqIG5F3+QjNVovh0oyByrAIbtwK3ujkXibMjYi
3OE5/8xavPnbzOxgk4X0HG1Qk2jv4sxdaMJWOK4SNuKsiujQTF5CB8nSSOfeH3gU
72veH78JP9qrbmgYxwKKNUiTBS+QJlkQc+26sJs2Dp3iJQsqvZq3L110oFNSNHjN
MKPq/G0VQLvRzmHfHQzdCO/AMJgvxP3iHkGkwnOmJX8ZnrZCnDWhjLAh+ZFIdKwQ
bJ/7ZaIK4ZRvS2VpRwqsgYpsJVrVNgMBvrwSpRxhT2UjbtQFSnEqI4LYnZCQv2n1
KHdr4VdCL5fOYsw1jgYsI6vOxjy18CW3KBNyCSKNZ/nb1QkmBMsvX2IPOA6kbSm8
rU2xwwuj7NdQnVRYD/5+Yhv+va3ltb6PDpJ4OUku4dF8mO2ormxGYrKLxOJGOhHt
leR42GEqgSclmHBjg0TRpJuzXUw/LamWbnVtgi6CcZBKBxmxhINd47xk6oSUfHnA
9tDLo/qjbK1IJq/KDVxtfmCSduypw6wwXOygGy+1yL/minUyiS9tdkB9NCmI0Ibj
EYr0DBl7A1qeHdyfUm9bn+Lo6fSjhUs5PR+9dw4Z/JUPGQwbQWOpTbY0EuzefQ4k
2ndCu7olsf1DtYvr24shxhO/ir7icF8l2oEHirL0XlJaGAS1LSIMul3QHrnXErYR
0MtB9pTBrk/hu769S7pb+6houwaDMnzLmrfG/j5aN1OSTkeLT01RZsb0q6MXubzP
SMArnDMDB9d2GVcce67MHjPRwNx/bYEflfat6VtBLXQc5p6xyFt6r3Cu7eFcm18j
7+9h62baAN962qxDV/PyIachdNb8g5xgEJn3IUn90ReW2gG4Ve0kE4nUyvFGFEFA
bYOpI0P6AE753zbv5phf8touiUim9VsGwuGokAmAKFs6gxcgtJ6w0V2MwlQVjdO3
3aCsHOMt0ip+o1XP13SRr45s8K1vWo+fWbzk4oStMzXoxS0rBr2857UbGrcYD2wo
LVqgw/LA7p9dHRNMeAhYMbj/lLTx7JBVINl5vbx/wN+YnjR2VFKdrWr20Mtpys0+
rATAENuCEj+wCiNlhF/cBkyXTpCmquimsh83DLobt96+KfXxc3PTv/wF43Fm2oEI
lS9N3nzebZPLcu2D4twew/XYV8Wj+XagaKubMf2lzUNGecoo52hkS7kL3KTnjBao
P4/xXI2hSUvaCnwJaSo00kvMul7ccfJUHNPtCOqZGKZpsc5DsioMkmIiTtR6LUDS
xrMe/SRq1n8E7Vr5laJvH4Bcou03w7BSu7GP4+S+nmUPQFq5ScM9zkirjRfPEghQ
MOe2kEas1Xld9DlelQncdLxYxNzhwC5yj1By9xXwHZCyWfkOKAvHSNVxiA69IQtY
eL1usCpX69U0KawwzxEgRZ3E2cy9IsAWGN/6PIOZ6anb/49rCGT1kJvNszO7iad1
Az/f6tCONu325GwwtuAvk0cuTJvUudpLuOrcZftoTzTrvVUY+oqRG+vifjhm/eXg
xr4mlw1KFWdKyEQ9RqCHm4LvDlKgL31YcqzXVc3IdLom/O5QgniJsDtyNE+1LTE/
cLbtUgnSdXzJ1AwPKorxPDsawk482Yo4Vr3LJ6acBGBmXcFrpPwl0qabnQ8BaRiA
HYO4Vi7Tuys3JYSu7xmKQw+N0e2R8mAfCKwwTTkVQUIwvEOEZvDf/VduiqsH6ekS
tMhPSuWXwG+VigVXg53/zzqyRfo7jLJPO1ezgK/GK/vb4hpkxI7nsCkSpuuTlnOD
Q0Hb8MqVprbokSvCz2YGAdjEToVBi44GvA+amzQluXeYkfsVPeA8sQouUeFmtzXn
vVoLY5yf5X4paqOpH0jmeV3eyHNuVawlv5nJ79kkcl36Qfb9PsW9v6JlWS7XrxKF
A1IJ7bPROACxG//W3n9PWnk8xiVpmkX0M9OTu3gf98z6tRQDCCDuPoWAH17Ygqtw
NU7AxtaakPygemRcmA/BSO0106aULpBCVzMv2S21SSdhE7S+7ZnZOwBotZZcP4Km
Ivybzu91OuqqM40v3V88HjwTLBjQBgSHimhWre+k4Gimspgs8zdJ/hwwd7UKx7rk
iamFN/vnWfj0Gk6Ry4Psndi7+E+angmNoQOhjgwL46VF9kiDPGmHFj4QLtHGeAzG
RtMrp3hQrjqNiBxjsoXQBVRSboCFxICOgpZxKl+hg7BPHixjMABWDvdxzTVfmIAW
48+F1j0ThAf4hn7RG1YCny60dtRRqXWvTI8lSq+87SXFKz7Uj8hjIlCFr4cbmVnm
a6L4rBh+P3xBEBCd9ZkniWjYl5ZdBihseHp+a0rDpipzdZFnZXMTRPeM+IAPpRlO
MmS/f0BY8N2ns/iPeGJb1glk05YikL8VzO+mtfZZk7qjvVeu9m/22MbbZ6lZ15LR
25SnDAL+Vb/qcIHJ8EiV09W48BM9Uny4XUsY9Hb0Ad6jDm7g5dI3bKjR1Fv8IfxI
Dw3HxqzTWNuRBXXHEAkvZUgvEJCM5oEK6K3C7h2yRwXKp2dJzIglBXf5SVNTIqmQ
DUwARp4mPug6kvy/SGBa/f/w1UBMN6rQxkoRhLFtoedMq8gBsPMQnhFRZqAFvBy7
yJ9hte3i25q+UudWfeBgQHqfbx+nX5QY4n5mGfh9HmpN5gcnnQNArqq1wpuO2/LQ
pCyN/eTH6952TJgRiuHl9iw8IiMwgYPF55Vg4qk8TiwHKax9blOX4+v81GYe4xmX
ZPg9D3Klccyv06dhNAY5/a9oZDSc5dtxmbieTAt5I0++e9mUjUv4MJ3IW2n0YFLH
sKn6j9glmzIXcPr5vfnWaEf3j6l/CfQpV8YwELXF7VM4/sU8SJqs2PfrTl2Y3RXv
RW5Z1tUcY5p4+CKwAoIAyk2OxrqdEcfab5Z2waXrtfQV6qInmVhi/s1GW/pqo9ea
7WvwHKZ3wn0Wo+sS0miD1dKatzZiOy3ck1s25foct0le+QzCaSghCmTyF5GfMHZ/
HviNBmkVSlB3lrylYfB+AoKrCGIWVnt+ps78UlSMfOWh81nf4wJeLIDdWn4SpL+2
NRBawRw5ap2AdTxE+LqpfM1LLCAxtBx7Wi2FLV099QVLyVfbSg/fW4VZaw9CpBII
KWWS8ofRSXQws4Q4fBRSSY7PEMynGehRoVgIQW2knxLKoxNy+zZYrEivodpqJXHo
QytEFm31OsDCdXi4PrG7qHCjW4khoA342W0Hs8v8U2jbqhfH5U6uAxhKwu3ivp9e
BS69aysPuVQTZPvi2HzTCggudenW9GnrymDJq+8DXSMOEfBfPwv91qU3ueeIyUTZ
uDIzqDZsoEOHJGS+/yRNlXGPLqoV4Ck2rW2kXwhDNd5bpF6jX9823ug2XojkYRsF
yo5Fg91Q1EdzaROaLeyjKTFUPWK2RU2YxwT1zxjAjP6kuMDaZGBKrPcNc1miVH9c
YA55hHsQJzz4CuwZXoUXce4dev7qbYDvzoOhUQEykIfPsFbyp1QUI5S/Gq8512pT
CjXqibWSG3dAQYI+F1wnfpVjuou9oyKa19ADwaABbiO/RLkMPCFik6UlVozzriYM
ERCqxqNdchUF/85yfXjy5uSEXKo+zqPyTPGJAct55m3AsFb7m8hvS7zKSiu+AWNr
ZereQXoFD+iE3r3LjtYvVmIcLJZKqwhUp6fg+vPYgGaYXNpwMr0fFdFwc2Z9LrWO
/24UjFIq0jfMaqbeV6OMqCyyqKlGDLJ1/DixviyDpwIDmsWEUF/bR4QIL/Yh+jUt
nQKFRH+1fiavszPddRtwIHvw2FmYZcbW/0/Crj+k6gbT4El8INU5S6PyGD94lL+h
jCVD/P16enbOHRYyOc8/d0W7RWpYzfdTljtGkQirVkPzXfx5xyWo1QwcB/Cv4HfB
K5/HKz9fCIEjt+ByZnQJP5hUwPkMDwnWkz202FvnW0WG56GLinaB/yjARFqWdT4j
ZIaFmkdBENB8I6ANU3pUhHi5AY9fBbbd4NsLjs/eIDpACprXatasVpi8iRkmQnYL
2yQDVav5tGU57Pd2pAu0XSTnjlPByvMRjpqP55ndo/rmpqiRKVdf1TeRAbHZAKX8
WoV0fnn5SeverTcZEINS9Q1dKQTJmHtmqZgJyGdvE0Q1G51Qqc+n1ZsE49x8QSrm
Jlh0hoXZzEyy0VnPw/u7XC+Mbb0pnTdnnBqrfUGNNmc9xtaMNA5MZknwnMK91aB6
tltFAx4Q6vIWkPWN+TtjXbeXc/Q/zeUHRpHXGPg3+WJ6KmIWeY+8Cby9mupWdVUn
mH5j4/qqDimW0dNlsnzhYEULu/ui9423q0VcZ5SJU0vGec3OMnjerwYTGb1I071b
IWUon/ibKc0EU9NtBPFA6vjvujZTgweH64qERzgOblVoPb55yu/7ZF0XpdaNW5DS
zgIEuGkaeCbvVEfnjcdsigC1M2Dz0ycwUHSRiEWrc8VDAEhBI1FUQp3NhFoNkswe
LXMXp6faBpc89QuBOKcx4PluvpQipz0a5pTTm7g8wYp0QUDAnW2ANN18L2cJPBKp
Ytfz9AEWXTc0LgbTe/HNsXJUFNbRrcv2R2mqJEi5WgIxqBqku35svYnrc6r4tagS
ee3S7i5yIoKBjcrJym7DXZD0DfW78ovkzFTRmEOzAbDYDBACvTN2hhP1j8e7eai/
Do5BBmM0g6e6Fis6sdyvudmmvX5QDPF3AxiGXnmhS6OlJiRCC8rLtpQJvaiIXFTC
KC5EypPZYk2xKjv5VM9AQCJMTyraQ2YHrqry8EpGxWoUi2EcZSHFvTcYjI3eDzdX
ZzZXYVXR+msfg2XSNjViSDpiiiZUjhZd9//Tf9BK5f5wMtEjuqAhdaLRGyd1hnwI
PvcUCAcLxgaGfYdTu+smMIEvavunX2jKb2wZodfZYsFp4gVZ1S0MTwewyp1UuI0N
oZMQYxQTzdYM/9obB3Xkmz+UKDExQAArVWq4ekDOArhm1GpSKjSxH/K9txgt4hZG
89EKW0Y2ifFcqDfdSAIKdSdml+Q2r7T9SFeb+dGCoSCZhlfANiLVrbPUjnnKPIvH
WkDohbRcR1RBAnGiQlb/aVsxgdjjcit5HMrSSkSg8OqOxpUrAYvAN4dQrhouVE28
qhPCjzDn2Dp2iPr+zwhZEHpKWB++aGW+6UmvnyalHEyyUfZGvF7xpHHXeAQ+btvR
mbTR9ToKpeMBElaGDNl8zasi72dGpGVQE22OuFj6YxK4zIknfJycO8zR2yrwJlvY
1XnrY227duPVHqpsncxPbO3NhVQBymEyRE6z/Zk2PzMCdwZ624iYyUaTPpJkKDow
3RFtmSjZGxe9EnEsS+JQYwOUS8/NEctrmZqvEhI30EAv9C7hzIoNrZoi6KwAD3ey
08fkbxYlQjvXhyMkFScXnHMorij5fy50tP6Ck/SoAd7H7GR290k+OMD1HDo+lmGj
HdcKdRMc3u4giCa4dE8Dl8HK0QJWOS/St6TNpJPBDk6TRkAlWcGFW5jVXZbOqZ1b
5KZs7kP+kRRA5bMaa4afZXV1wtzNc6TYir+yuN8Cfwkrf/v3PvcTckKxLQReWU4K
znFyftwv5YBdgEcevBhAkk0KYbZbKzLKuLb6l26+LNDwr25Jl9dDLA6z5py0YeN9
Lt12jNDOWHzk8mGlY6pSNHo165DYNT168jaWXwbXZDDOLfBTygmwbskxweX8Q76Y
/BXzDGmw3cJvg9rat8Mc0ErkFax4Uj8R2OH9qqWXWfzYsqdpHEiczzy26GcNtywz
4bBugQkU33Sq4ayl6bHAXIRK/xbxFCohGJ016RiNufd2+whGtSodsVQjRGaPEZpE
ibSDWUYDzAFqiFYS0iSNAk5XXzgEN2kYLDndA2BIwujiHGW0gZEQNLO4sjFUdWMq
k0BqqkLXzk9MXfHO5aHv1FkpLjfrK9jYZlTFUXPJA3Fi6jbjpCew7ZaYVr69Bxz/
102zJCSD29uzJuMkukqDemVAQ+jPx6ezIDzQSKuKr6rUkRy8Jis/GdXRIWZI/aqe
kZeGcuru0GWbsE1guLraNLRjOx7lnGQArgIgxzwdCMKQ4RcUY4KQN6DbCx0EXHs7
Se8cXplaIwvHmgkmx6kw3HQ7193GxSwl4pyQQISLtjLd8WpcDkZ7cV9yQqOSKT0o
pPO3iZCXbmqhC3ixg+y/CV+SkxCSFkHE4PuKSH2Ck4MArqkwby6bQuaZpwbvej+U
Gg9CLe4hNEYqXNvhbeX8P145NjRbEr2HxOrDqrBncjeKGWitswyG96yJZPzUar64
TyD3Jcx3YpaQ2E5kAhsPJpjZuvHQ+yo4/xrHd5lSi9Zi9Bu1yeTGAxz7MtD2wCEE
qzul1ee6m371DQCt/xp89SZnolihC4c9A+94z0UVoZrO+HIIjeDKyGbvMPQWRiY5
p+wV5Nq6T8bDlZ0PlWi9rRmvaCRF1SRTzbb2Ddq35l6UlEuhAF1uhwaBdD+ygvMc
va5Ok+dbggRoOQe9OADunE2ylnxq66yt/0PSWhL+c5y3Y91FSXYmtA5MwmWWwBOI
BApEoV1kKT7ldGTzkrgKq+rvNUVvT20guEMJofOUuCmmgvPWBZL6BQ2GUQV8QDBY
5JzN49QWSAy35ysOCnbYZOwPCmDzos4pAL8Dzc5zraJeCpkR6VcKuUJeeszHG25f
SEOT2V8W4jIe3COmgxrHrkFB5gMaa9fFN2SIPsImvv8U19YZkI4kGwutA6IhDQEg
9BPY/P4yOMtdNtb+waEoC8FA53cG6V95r+hhKZd23DgSpA780PZLX4EoMUyg7aKD
r7fqYniSMH2LR/2R6gEw2UE3rGerszSw0Aa0tkyOqNj8yQ4sZtCEUfnvdG9SHjde
kq0Gs5o7qUKUKsJkBn32aAOQWEO3rc7LsPlaXabFUTaR6M0Uo9UrpRyaD0a3FSLc
foI+JrpcG7hfWwesDjp7zAbNuoCe+9TK4rocAQwr5z7cCeyxv7P3Tl7C5pxgWFu5
jksYATmLzrX/yfUlgtp5gmnnB4wMMtOZ2I6sbcgR3waJmSnXGBSe82wihbk26AEg
cZj2Tl8QY6VyuK45tmoC83JZHrxKSx9PqGeNEISOijQPj41vMzTU4EUBm3EL5aQO
Twqyf7ctAhky1naiZgtnWfBZ7Rruw7y9N7dfREAr10LqDzo0ldQLH+hSNhGcoZnn
y3QKxkJwYwYYSBFxL9E2wrNmLUDyCEQbtnPIwCaaO37lYFMTHff9+W8eRzvgF/CA
ZekKL9viGRtQOH4TTJq0HKen8xl39YbdtI75ZPf7N9OC1qbntof/he/OegfwORF3
jx6D9mdHxCO22e/eAmWDUILdloMuMI8z3xOvRUYLBzZWV5kZYlRGuOFSRjAbJ7Id
EtixYZn6AnazEkewGhQDY39no5snoXkPydz5YeFJyY3vrWYrj64Yk6zX22Lu1sIm
dcVugjejJqUYuhby5sp1emYd96kg+qbyJn+XA8tneXQVHMlOZJHNM3t7/d5+s2eZ
NnrvXL1O3yTZgO5uC04IPKxanYg0OK0y+Y1LXonNYFYYTPrpyob0HgE/ij3npUAi
PPyxgbAzd5jBdXAdg4muEi5JigJncCIBkRh+T+PcHhT908ZCxGhIACBLNajceY/1
QfCT/Ssp9HD9koCTUnboW569Y2tyInhpg5Fqjo3nmah83wcq5CY+rS2lt49J9xi4
FDeEOOj0TnGhB86CTjLfiO1zCxx7KR1fjKgPeB476BShOMlwzc7fy6wl5I8j5Ckc
OLJYKfaGcpbxJgXngAqtF9hcGiOah2pexD514DzhbBXoepJlLlZQZG8C8LCvremx
Sj5dmuvUvrA4Tihi5O+ezWOBcJDDyXEo4bLGaBAtjIqi55duDxfOdrlf5YlavZmn
8J2ZEAKNTHEiRohrHW/wsc32bQNVMSI5OxnJZJb/H+cTO+1WCC0jdp9LSHY81OLH
pHD/F2AW/TjCuFIv/pIxuOiAcFvX99V7tghCnD/yQzWrAnOIyMcU0OaAH0TnoFYO
bA53el6MduINvO6tMwQMA623tl+WNdkZbjvOTfEE6/Rkd+0O3WqrfWboT7g3cSFo
8MK72DGuO9zPgBhMzCcvO/2g/07NJUXIda0KvzLI+0ZsRQwa+f0k778WGJt4yw1y
+f0hUGB8v/pQQDZ1K4Vojrche13FDGPEzJl771q7eHNzNoptBL/rsPTr8vk/qQNB
x3ppvHJV8aS7S/iX/Qy0Bf/WxyppksBVLopchsh9XvWtykVLzLMkPQHRYEmMmKrX
CH+HkJPZGvqTa5xFjx1yfH1BHyzFsBOsGTs1lTO9+8KXTXDt1RgdLqT9WdXsjIGs
dETALuOt/EnRXRJFHmmtW2ied3/LSxSlVuQO2LiHoATQ2fyk1RaqMBMJcSpKsF3S
GA8FrSCRIJXSZlEGQjEDBa4XhsiUsK9vCdw4oIcMGYYLRC6QgHut+YMhR5GVNNMe
auBr3gzhFPZ65KGErR4oXoA/7kJBK75TB+V/avBAHklwYcBAZN8SQY5VIeUvwPXA
uL60lkm1WaiA7Zuv/jYlzeXO70qJ1/kSpWg4tuaCs7J8QGAdGjNHC5S8/IYJ7TsX
HmJ+SM8uPHdTKAeCq3YP7m0PURtXC1JwrplJnAFlUMi0fbKeYTiEzFL0z6AQ7vyI
NRGfYeN3rcnr/8PQzIzx9fKGmEoFGLDt75xyiuVX742kTg4BNlLG/Mi0vPL8qYBH
glqH9TPuu1EQohY/lbaofheBnYMWBIIK81LpuSpMpjJcvmFxLcnM7bCcL7WDx2OL
fF1W7eW7M0bwJ55WUVNskC+ORGHRxWhG0wNdURYtRNgSlF6JSo+b0ZTeor0RyNJy
uklEg3abdDvjCoChsB8oJ+0/z/d/6tTxnT2++FQvEYohrVKAV7mCt3xISQ0kad3X
gJQLsM2Q4erm9/fTBQi+xjwTNV3HXgeCjiK9m4GclnDyKU2lDFkU0xiIRBPS8GbF
z33p2RPQfo7II3ue0+TIn3Jd6MNqouqdGuri9rCFC+7OdP9XzjkoYvzhkZ+ojVo7
YaL8goMY4DW2YGTm54nTgnb+DbqTTq1CITCRckExAPv4rRjY2nGuOPS3IOx37hG/
ahvV+OxObFM3G90ovm/ikvf53YBw+T1oJY5BiSnV1OU8Lx253EUXlIl+iEsEDM9l
dtojE17zvqR5+XVKIN3pZv/p2kwqxoM6/ZtTU9d+syUUhbDQ0d3zrRxaCQeijFFR
gvYsTGA9v0Z3FEsNvschQJIT6/LpSTGkeo1Ti8olLwG8fmqFWHy6kcXRu51mJMmV
7g/ak9oEl0cDvw3p6eo7rGJda/vwNlIXK4wmBWwZGViwXW7NOS/Mp6b9s29gPnVx
spAAFLLuXRY85ipOqDZGpiuCbkEM5Ly32uR2KMHSIW9WvwG0mn8J82CSB3Lq+jPG
8Fmy9Set7HnUbKQY/hx+qXfMROp2Qnj9CmuPYes2qOQykHl/9R2ze9zsoDIzHRW1
K5xmadUF5ysK4ki8++Iomn0jkptLasDNh/6/5x3HBV46jD2PCVZhA3cvCvTZh26f
j3GPI67RaEhOBmnI/MLZpn39DFROfjOceabZsHM3wsvr2ZU5e4T/1rr4puym5KBN
hGlK1631WfOKLGhA0K5u530ttc4KHCLrqqwPc3BKCYGocL+QaM3/4jIbOehjlg3E
jNJvj73Q2xX79cdbzC5aLDHBj3G3b31RRhypWa9LKcJ0rBtepRGGnydLKvBQY1PO
YL1MmWB7pwcQpuAAcoXqQi16z17s4UqotS8yvyHrkxYDt+tzpXsyEKrqu63cRew3
Otv8FXkIE35Azmisz+BHxj+NtbGh3tsVfYspcfvN2uQaMQP5KM1WrtqVIPNwqjRY
QN9rxeOsPT2xcPxqD6jhU6E5sxpY2rwcXcYrOOkqTsXyoc9gnbvSq6IPm9MiJ5YF
ZSZKGme45SKJINRsWljS920AkIBC1VEqzX3KPUjEkRwNGw6OAJ6V+ixeBOVUAAds
Ikn9l0sZoFHEgyn8epD6bMB4JSl75D4TAFfAel/tvoCEk7XWp9a3KrEFfFyevMvf
hRYFWfFV2IFQXrI5dP/TA2Kc0lvWC7qd4I1/v7VCoRZsHwskBbjcBEjyOynKve+e
k+s+99PvJF28m0bsaWI2yL5u6WbQ8TgQm+tkhv5dzGRS6POBVmc2skwJ54DxrKQy
EkDNoi+PPZemniKidLeaUvxQL29llEDQfqtkbSX7SqCFEFNi1n140TTklzZ683D/
gNJbyq6ZxpZ9bk+05zKfdGtNT/oeUM25d/NDrQtohRRDl8jlejO80YIaIJRAGopn
zXRhXd+rSAm2I6JgoKcnD59qgLhGLz0k018wXRiEuK4f6RgUnM8RmAS2O00ryk6Q
lkxI2vKGDFBdOp9KgGKCCUP70N1ZiAlfJUBkxSVyMhl41uSC7UmDabJhG5hBr61I
l471KVt0cyb5sElKrq9cFIhgGwAbKubn9EgIgtL8AfJMaNebXbVqHl63idJUPlSh
pNhesiwQL9fyl3ooHWBAIYvjwxY4o0dmkCGi0Imn+d+8dxE3ejn1buuBDOEbfj8/
XjILCoU2X42GGZ63NjQKgatvLskcLQZM/k207JWz3Cq0ZCY+R4uqz00xKAmToi2A
+RTVhWBMmoeZq/K4Gek2eBbQwOaSmPdTWUrHSXzwOhqyNhBOt3ZwvI6gZnJ8rOi3
hFGn+ivN5cdmS5N9KwlIS3FonW2qmq/RI8aFtqLbo6lkJK9XSEt5Mrevdf4VczF2
3aAGeoSf2Mfp+bchXkY6rRJvbjpPa2KiSENFj2o3snl1Ev23Ah7+ZBfti7ikiH2Q
ebqscIIpbGc3+9ywUL5T4e/yGwjIXOgn9NquKWzHvr3vy4e2EpVXt9bdo+rp/dbF
d7sRxc9KWIBEREpuExZJAEYSR3p2GHZN2KCJb8Hj8eMGylR3T48je1WM+MPC48RZ
60Fe0qVVtyYAa/J3+T1cf9zxS92My48WbaZKB5t26tyPi7tNrJfRhg8Er2pGPee/
46U91XYq3v5TtYpqLMfG6uJC9VeUvbou81qWc4XgDVwuIDjHZF2m+rXPqDD5oSD2
LtJkMDKaa0h2MOp7hY9UTRlrfxCcYXp0a34lts48OBGV/AZCZUaZiCXX4O+FVZH8
POY7NPxIki6M2qVuv8+P4foW4uk1pDSn612n0DlXEVJBkSdLvMV6MLaxw1h0HR62
CXgb6d/0nGt8hrO+Hp8GPQF7qvLO/J8ckqyAAHInLAoyoKfseR7EJ7aC15mFKsan
IeZdU/5IAFBpCEr3x3MSPGH1xbvmLjwuYmkh5I8ypy97SfWg+x5F+LejSkllgPMZ
sB3nVB9cAFtBCdWeUT+hdBMFm/WkhDcmmmGthqZrezpPiBXbEB7t6IhT4Crwnrch
hLdVKu18kH9YTKCQEtDHrdM1si+l3coOFKd0M65wrK/komZgJvPn+PFC0U8r+IBk
7bBXuHt3YAl5ay/4PSTthEuLmSmzZS/UJuNPiUcOInMBOTi5cAjG/AUQI4dbRsZY
MuJYnp1ArwotZ6yinVSR9zX9ZDokta7vPue+3W+tBx+Tp10OWG3OIt2tvo+cNjDp
f2+HPpkaO7Hb9UcL0vdDE9sZgw0CUBY5vj0z7TBORlRqwS0a2SMToEthrZzg4KVm
g56SjI3wN0wqG2DckpmZNaOMhYNZv20wjzVfZBBsIBk9o8c/xYiuNryUpQfJsalw
EcmlD2HnQGR98N4j1UI4IwjeTnkrB8OzxS7JuIJggd55+fp6HwQG7gh6ieAJdkv0
LaLoN4GRHlmv6N8tx7Gz2jMKBf7VwDW1kOrxvWSG66xqJvFtDjEwHdF9HMEdRhG0
rWYI55j5lPDIr95FOrWYBwc7C2LzvvshenwFXdj1AuhHFQs46OcIodKXX1jl7jsc
YgaqBiw3qzeQTGGKv6+YIiWaCBiFZvPyqBwg6ALW0tAbRHIsWkSiZ6+PkZE9kByg
pYHCuFFbbZXDnsThBpu1RfG/1T9tGv98LcCOeynZ5+C1rlidf5VQb8uEY8d17bYT
MjKfiX0XcaUlEq/58WdFW2eU3FKNqzjIyGDjx0LNJV4xcWyTgnvDv8AxqhGaQ1A3
4AFgUJUc1fnKB6+tsMaKEtX6KylTKwd3CfIde2kI0oDdrv1LOsaAfVLHlX1OsAEK
tRXf3tf9UrWx2LpYxEyh/gJvQlagGF9IQ4XNKi8xcQS2lzExU8+WJJxmLQgVq3FN
mWiRfPzpmvZRMDo5Qa3HleB6DShHGlkPFejC8dVGkSTU/kapTNE2kogLARb5mD85
XTopt5pbI9skJvviauoTGlA+gBn+ASSX0crhY0qfaDDbP+caud9JwmxPy9yYPfzT
EnwHbLMXs/niw2Ul5zh02Xdbb79vJoo7Q2Kv17Le5cuSggWIO2BqU0Ru+UCZwiUB
5P/9wbQkaIQpToi8y8PWrHx3W32miUwHMgi8GUsKEL9FkB8Bewvy7eRVT01cCpm/
/NsbgMKvCbks4njKfJ1Rzbp3tkhikCn4zUvQ8VrB9971cAYW6rCSlVSFbWL5/Nse
6ou1XwK+YBgylo0jch/AuE4QHncBwjAZ+JQOTZOlxyj+eit1kElBgWuAcklG6Id4
EjrTECvJPO0UPtNJwKolsudnOYphG46UeSnf6H7Jq1nXB4IligIT7ckA0qvHD7Hu
akrlwXLYEGKf3iNS3i9DWLQNbLUlVmmqVlI39OUC9+DEXev6HeYAFNZve+D+vG5s
2Nut+XT6cjc136yzIM/I2zDO3AOuUEIN/2Y9nO8NSlcmN45KOoPkFBOFo03sJzVj
SC1fFEsTa1tbsJuUp0cuzBpRhuk+3hENdxGVNo/bZTaSaokswb2drBaTur6UYmvq
YAyoaQtYAtxSKbFz9/sEjvzbtaa1bdfPUKE3Yh3N0kEz4KRVA+tArrsjG4A3IH1F
HkpvOgtioAMDWXCKBPja7FKYB/RERswsoAyg8NfwVn8Uw98eM3bIKatA2VFjUHu2
qhVIYPIILiPc+mesKKUP0fR5Fou7LrrP35V/UkB6FIIq19o3BCTMDjlcKIvCgxAD
1aGDKYA8kkJzVWtWH4f1KSOH+L6w0Gqck2R16XvmOtboYxPyc8IuoGPVFVnfp1fZ
nT8nkwfhcJRrp+d/OcsfwZhwDv51smIu+WT7z0Sm48T0c7j+gzdjq3VMNvNuuxUf
ldvE1zbnqw/soyb1m9BRhrasipEnhgmlVTEa/bpxiY/cdV2RzkEP7gw0F9q3EXYv
dfZVC18t2BNrLRRHcTqk47ocMIsTPWtVkzofIf3mqCktljZ94QiA5w8hskaAnuCt
uQVKK/54q+u8kq6CujHbLJ/3MmvxkEAFaprPnM6WIzTXGsBQAaZxVmb1WP5V8zGc
ffc7bEEQeThFjW5+u3vNw5EHhrdlsfdwnnz/UzvE0C8G6N/JBIp+PK2GpMA1wKkP
nzEOWATrcHjRViq3hbJ0zbV4JEnkToHjI+A/IiIF1A0giWfzUvAhKHBy0HdyICix
++oQlsnUkThp1AZ1tzp43WJR0OWm0zq42cfWVRSCDcC7nAzhNrjfYRKmmdV62j8X
LH3TDATPyTWrnjE8V8mqMbpcMUAshl2K/1LPGcPzdvvO3CVDHqRo9hL6MJHUpt1r
jg0zS8o74znAr1eMVTg8ZdUoweYu4EufpotOT4xjP7vjHCPdk1+C+VNpsmDkOLiv
mQR5N+vYIJOuI9CtlJ7o99g5fu286+RIERkIr4a5OqEHR3Ox+xM1TiUNUHshSh1b
pUqWpEjjhxG0x/pU4VdH2RYEOApgKWYzMalCNZmAmwtcPkWubyOKTD1s7mqt8Psa
lruTaXF2QzHncX0MSoubFo1zgUR2Q4dPubZYhn0264UALQQpy3nPYgp3P0DI8Oso
R7kayEOnE+eV0HlR/kNEXEkfa2qc+5Hx07XGgk4UMjbTF47Mj7L+UNHx6eqGb39p
+gbuJtXEttqXDdIWxhWx7H/rnOMDcrBguf2BMtPI8yxtKnngOMVY4LfEJAj4Xnql
/6323/as6k+/zGoJksOgHdgaEOAWFhCcWS9otMaqsdizMo+3ohAA2CAYs26x4kvi
j4AZSgw6njWTFbTAGHRBCazRJ4omBfPr1Si9w5N2qM64HtgUklwpeSO/XIlYuLjK
JEPAVW47rKS4p8zdLnYw8BGTeLl86TASFQvxIzBltzAC7T/+eXlptrsaHX49gata
yaA0c7QoWeN779J9HMnW5ejjrBDBxI+1+SvNIEKP9x81gymj0ybPLxB/I26Lj6lG
jUsVluVPL2cPQtzeiUfkl4nvVz7ofom00cIjgvHYO3y/qY5wi33HGAsvqrZlLcA5
1zGqRwPX+P7v+8o3/1dOs3dp3z/63H3jBFYM1Dsv12QX+kUBLNEuHQ9D4IYlAOMp
UuPH4LQr7whPAugLRlnD8lj7vUMXmYS0QrsGDd6bP6h2YUpyl3S/rQOqaDz8D6Hj
kyPHzmeplVTfPDIHPvmozyQ5Ytffm1KPckdC7A8WUjVhcPQuHDAAQ9F+a6/i4K1S
+wgl8rbqx4MSw314kOkGlCYpreRawuX4KNm7dSoHl7Y/KVPOUPvPHyIGmuNGziJY
63CvyfdBxbv43CKITsG/xqtYDRIEqFwf1LCZj1z8So96EifZOadi3ZB+65R7zhx2
lCSzx0HnJrAQv0l2+iw4OEAtTPb4bFB5kmFHDXP1iqSZQtjqKpvN0QcHgqsWgZG0
jgiVe659PyZmawbPVxCA4BY01EUxdZZQoYvq/Zsj2X9/EIgFQOlSbhUtkk1F3ffD
2l0jOp/XhjiVpwWViym3FQ1i2MXan72CjGDUyboxCEK/Ugz1vww3e3ixk1U3cN7l
Zp3e0bepzsq5BhbVWveqKjvILsrsWLr/lWj7BxYo2598gxRmrUtL6Y0cC30+pnhD
pXSPtOkoSq4qWEMEX/NiScXr/Suc78noigX32o7Kzb7rZGPo8xfhCpNoidZlMO+A
e+I34mXFPyObRETw29xtIbJGLYhrwgVsLp4voXs/NvXljqi5KSjwHceJNAT+0kuU
ZNSwEpetpUW5JX2Yg2ypjI+pMWx/buzp8B8BLmRJPqsuVzTBzZJws8/huvktuP3/
of6lnFchXv06Kz+TeIMH8UhkabW0UjiNqR8Yovwsu/7p41gtQc6tcNn/h9bFlJkt
vMwyCAij3XmgTobk3ygAeqJ4MaeaHbmXHBRZXfAwrCM1wO0t2RvwlbCGV2067enH
bobNvj0cPtSm//WeK8Q/HZ825Dv/uzMCyWyQTVSpgysTxxVVshtO6mEVInnkf2PR
FD0VF5lu9Winii0yo5P9G9/qkPWUdq/bBgrqmD69+unY4LK/BsZL3yWcx06U1Lxr
V/+/n9iZaiqL05VsAyJz+rKYmfbDcrGTl3OI5+dFwg7atnSGCqPFkLVnjnmdVoFX
oBfhJSykMeOgmCNwqviGuoRs91Onx+AhXqwCE00236NIc07r8eS80tWkRjTwzRUM
Z7Eu/zj0MFbKjnCCMHao/2kuAk+Ix0bp1iefsNH9jdKXZUdDlezxfCCZlNrF+knK
L7BPVVGm+buwKb7vM87RESaukQ4ehz1cyvLKA5dZeOsKwjBk3BBrg5WNGavYR49I
rMCSHsCvXNAGHCJbziSKL2SNnPFnv7KHfW9ujWyPxAE240Gw2V3K6ra6R558VqRB
M0ucGGGmh7eeKxQPGd8OD+6GfsuqOodiscbRNizyFiV/8KekVPkLGIq3VNjxxwxy
3FdtGWhREo255D2GR3ttZgAsR4cDYJoL8hP/t8/Maux5HHJhTHXNGTGOwyO8Hmhi
CafVCpXajqqaeIe4HmYDC3jSgGJHXPaQWyMEEl0v1+C2gI00tkx3N3z/NlRv8LqP
yK5cBkHq+gkzl1pGlcAmA76OK1Uhuy8tMbJeTRl9DlZr5BYKIFcrCrKs9Xu8foO7
2qdTKcZ0rHHqnZR86sRYLdtyr1PDlSTJAe2h8vZRz0mXFnbYu4/y61FaLrJ7+PsA
nKri2DpbmpHg4TI0x+t9KOX9z0ckRJQJsyli3aiisd2N6FE4kV70Vn1COPssDzpL
ZLw9i94pTLCvN2YD3yesJoiaBF2WM6dUds/tsHV4dslI5MJHVUxGTewQi8MFQh8V
NQwRBmcxtgTFACPUP4hwpRPTPfIGwzPh+0YUZym0mzlhTAfW19McjPRRwHUNHQNS
JrdWOMOkwyGeJRrxhzmNek2lsMU68skyJujOZ8UU6Wh/CIlX2B7h70krAVrSvpAg
vV5lk8aidC0RP15PfSDZOPYCtybLyRt42QEkKrl6G3wVc0ZUrn3KqNzKEKKZe2Fd
R3Rs7Qrn9QjLHvqFoYpWIEM6par9nZ0TFCGEKPL2IAUD0aexn0aGpUsT0SaRg7hu
ygM2KBNKjPiCObmMO5DgJWcSWxxtMB5DxRPPTyKaWbXLxbUj2ENPXE49Izo4i/5h
xQI7PvI6k2lg6h0d+w1zHoMP3iJxVx81xH6bRigOBO2fMBToRK1oFbaM3oq4UNHx
RRtKYnWg99IXpesVAJNfZcMTm4x4o9r8g90ro85rbbsdBxQxBHBJtjf+tCWB/NZ7
PdkCVaQPuJOo+oF8VrhP67kuvEgIy715du/s0Q7s2mvdJKIbSOAndwnroZw/1rXV
0khBZuvAFvhYZwNBmAoxkF7dfTLB6RxmAH7Ia0aQIVxhvpB54J1KEb1N6yO+6VDU
NIFviKNAfpdq1gIavzBmcIKi38+tRl7bxVQ8YS5EyIaigC0dBK6IQMbxZsjBqA9e
gQr1PJJjfiyucEJ6d/ng+8gujCn1AyWpHNmjN6asrK+ssLyzMxQLt+9cDq+Lgv6w
Ziw3A3mtSy6/A22RBsjjiY/BI/TuKN5nthOmef6wzDIAkPrRGz0TI5T0byDCLytf
AOkUlNaystASa5M2moPL7kHIYdhNL8c1USarAZ2P5IyaqvELJt77yQBA2jYDvoyT
/Gg00CpRnKZ3VSanvf2Kui/JvEC88F6zEd39kwNINfX2G62oNPWcgtuy0o4p5IBa
sa8EBimCZl8qHHUqniozBSs0RTKgqLouNuK6p4DeNpzZdlY2E+BuvN0yMBSFmjsQ
DSXr6gQZgrm/vF7dugwNtyYQXRd2WPyQgWd6RI3Hgl3XETnVy7my4OqVZQGe3i/d
tAnhBUmnuCKicDdTeDjWtE0ABqabehVRO4Iohs5V56kDSfaAT/nwmQs52r0UBGz6
udei/8SNK00xsbXu7qJUm1snv67YTThuYYJE655PhlP85qm1W8wc0SoluEYpRwxQ
pThgBxEeEl980EfwNPITayjO4DlJzCkcgqh8ObdHJMYFnM96yVSzlDzf0hHrLHiY
+NQROXH6f7MKZqI64axXotnKyumFtXBHBGdkBo3gSj9lQ9UCwWcb/NDw6CRyH49u
Pb6TGZAvVEwGM3ihUD4XFs94xPH+qSGP+0gMAPM3lCjoIuzl+MaRKDwGPxgt5ssW
jGDrCif2PS83ibsp13XIZ7UhI/JwXDUYNRxcFT/U0eCfCgVfyJR8eaTIUjkTt3eF
XL0JhReDfYVTSKi1xXaONe4lgBS6+fw3c793P1Ze6cTbm2BRMP6eQqFJzPApJzIX
ntXQ8eq2Gow36NqlBny3cZmA7ZB0+XZHsiu0tiAVmfkM6wR/KBzZpA3sf3X1DA7q
K0d5rVl3hNKh3Lvgve3kuMTAkhIaMoKQg9KYZU6GEnR2QwjjRZVizgtRtMdIWypB
ZINVIObmAR9K/GDui7sp3n5F4W+UwcSXAiIyWNsmDt3hHfkXq99V6LX7qiteqvOq
3eY965yidldjeBQfO7CLxaY5eOTjBjsIhXcYQnH3MSgh9wZOwWQhky0gSak4Fke5
xOt72DWz9M32xFYynYQVebTfE17Ft5TstdQciKU0LoDUxVmDrqFFy/KQww70Oo+P
Pv99n62T8wnfO8r+GhZ7W+KKeIptO81+7iTJixX6qKPEjOMbF96NHl2G4qDJFDMh
I/jEaJ6FWaewlbH7uvz02l+QA3FZADzW+OUQqnqfm4RNSzPT0A4gxY57GZrCxh/8
T5cMEiSbLdN8j3+ODvDA77ulCEuUNLaD/78FLQMlbmSkb1n/JqL4WROzPn9XSv3X
0r5xlV04CoxQvUiHVDtM3pmZpYkeM6FLAV2WkQva+Sjrcms+pcgst6pcMo7u6bFV
iMe62R28rpUv/OAKoKHRC6M48rIKtnIpayjoOdM9zX7uUQswnkyU/OjsDLO5j4Ah
Bsx2q6hQB0zRN3RCERk0OnbikEGogfzA/w1qjK06B/tLYSbLcd29c+aItUYxYrIk
NXjDvlRfMfE645MIVGUozJPFwapXPaqxPtB6ruJn7DcZpAqQ5+fCApfyclBEx+i6
qscCvOqFhZeAya/T9shZ1WqlSD+T2CLh64w3Zw6kBUAJlN3sSpshzYSwW4DOFEv6
azUmH7lgsmjAeydF3Za9CpH9oRzJ1e7eDN3IJxPU1Jb5OiPjlKl0ovuj+AQ57r0m
9c3SHwcP6SjKc84OKGWOEyQRokoU1V07Z/oIRLOvDWQdJvgavlAUWVi6JDS/mZSy
FzH7PiZh9rnsLtJe71e2mXhaV+89gd5UXFsAubM+XhSCuz8okPwuSBk6mdbv6Izg
vXZ4WM0b8IanRSBzlau1V80Yv2CHRiayUJLh1akC2eG1hMkpeuYQ3TfiE40X9xYW
Qdn4NT5FkxikBRBTqMzSqWngAubvidSlzk8jwIFiroZH+6BdXFRGuJJgOVwlhOR0
v2LvcXo7WYhWJj3Pyr+pbtkMdqiac/nFmaxJ2c4P2h1UAJbX2FeYpRv0SYw9qn4S
ZXTUzr78C2aP8UC+Wg110ZY7YOhak85KXvDncdVyK8qwvMGdJ8VgwbsGzsH/xjdp
8D/PDfVjqOg3STOChVOl0HE4zZOpGzaj+RbcrLiQQS90+UZs85VYAN3xSzGuw2Rv
7lfoEMhqXpNaRVOPBpOjoYdNel8TqIynduBY35HBOTZsBSW2QHM29MJ4RlUTMKlH
QuualLutTafRXflgpQkA39iyWPOuWv0ib5A4h84ENKsLFea4/Qwf4MQwwQtri7al
oUJ0MI/HSmE4P+9TAGCameyHQqluxyY1NwrsWh0i2o/Jm0R1clQxuRoRgzMOyNiD
YUfQT2KTY+/rPwwUaJX0rM7u5IPKMYsa49sUvdKZxKT6FuPG+h2PToaGprlhVaIu
BKe1IMx/rYXndXzNJmYwvYwr8AbcW2FxnMe9E0e2o46pS6/cmLIzUayvqeyledoV
TnmpTScpKokchrjv7kj2vpFbA+O0QVdSfoGun1c5sWCDi86WNnC/NWTaCfFzEmIA
ga/VMSbRsLHHQSwW0JXKntGaWZlklnE6RkIForUS3S6lM+bWoZt/8nFgvCswrwki
Kgyq4hl2dBSSaRGnjcgaWir0c95t2/+r/BuOV4y6If3Lc44rFi+EmHhXk+8BwR4j
nvw1QacIASuCLBLDOuNZdHrFn7yFFtNQS13tbGMcFfE4yNwFftrRuuxH6zg4noDP
yIH/2soyU3nX1ntx+Qe9L0HIST+yPtaxR9yKpNXYxarls9ksWJAGYo9jULgkXu1U
Twqy+VieUv8lFsRhc0qvq5jTeIK3eCgH4o2DMvC5YoS6QX1tR/i2vPEC9KVv/+7e
e+NRGEBsfsKy1I6tYWcqC5duVhm+Nc5OQoKUh9IwIaMTqxrFSQ0hE7AcfLgUx9XM
RbHWze4p6DfpyhmH8QEhffW+N1QVdusCkmS8vj9Ltz0vgDPRtJn0srqJPVexnp+B
jhxAo7uFFCj5+HvJny8kwt40jnyP4wQl3ObUIqiD8jkYUtyF9FXD7HS17I95w7Rr
csKqN+2OoYV732o3CGJ3GMHkRcBxPC+O+DVWxEXSiMwjN/QF88oRnX9nE3Aqalni
5O2tTiZqqJMpGo3Gy2wphWoJr3V/eLnL/orlND678IXkli/RPWlatF7GcNs5IyY0
ygAj5wTqF13v1kk0LhaxvaJjcRG2S29HESVsXoXfG0wjD5dioxovdOTK9CmWDVgw
jY9YsQa8x0BSNrb2aJKix1r+srZPa9Luy1HfQIhpmiieCKQvd0mbJr4zamrNHhBn
kI2CGIRKNo+EJAqk5+EZlDDGVbXJSoFUCLyCRxSJ1Y0KCl2CfEKBpdZdZ76m2sbT
FHC6tyEfs8SULwGxtwwWCpn2ar6Atg47HiFh7hBpa+CyfCH0dPAQiVyIs5OXmNxg
7Q0zgNjrhDwOHuXUWo0tntjju33XGGouJ7x6ZPr3671422dO/VDJiWXb69i1dKuB
dY+fDUZXyFAT1wjGzJ40epu7gprpnZ5YuUNv8UWWDuRewyKj1ovwBWwy8qvUoEEy
Nq2tZmmOv/trJefL9st3e0/fCqrhUkoAu4zSlmIuVmeJwt8OTIpPiI+s6h4YDv8i
ECFfpyY1BmHx5cUeNhR9RbzvAWn6eCnVIiD5TEDET9pHL9zj8YA+91PgPsJGeudv
OgoNwMjpHLPKpefa5KzHnZj1fMPqyA9uI/IgAiv3vHPBp64sI6fDKKBa3zIwdG2p
0S85V4cCOHrz9zxzRHcIXL05hmGU55Vx8hHTM+90ex0XRUA/4WjS+6Ea5iDZPki7
jSqZxKQiUAyQEc+vv4RJTowUV2oNES1+p5KXrjJLaaif4K2LzXoWVy0ewsJV2wVQ
rEoQetpIC5FTp45uihVyLm/vVoqqg+UMhdRm3ZKwPpD9wNcu2L+qXM1ZSS/GJhVb
PFWK1K6QzfSXuOcTeMfZFMZWCxWHF7XRVbhklrTl2MrQpuFK6FVDoY3Q6LNxTOIz
mKCdyMK/cHQr2NK0WW68INUi1nSeirgppr7iwgevgRwxzIyv1G+XvSbRxXaqx0U+
zYqjBBcM0K1zcAwgSvzS20itIrpeuHSDRWE1/0crb9oDqpWXnRrsCc9TJJoFP7Ia
64nrqvBnbk73pVoqGRihSXjlHcHMFFyER+5smOESK90w4IEyLCJXhqNpAXRGOkp0
uOD1Vcu9ieDL/PmUMD04ZewubvIJXY8RcYr0icp7SRFbJ7X77zjnzy6m2ivWJ2YX
ie0dB34aXb2U1RH4t9Ry/uHEGGvNZcR3qZ+pQ14QvEtmB1k5d1w5S7CXgmMN+ucN
A8nn97RF926xNk5d3GdbZb514g3tLbq45ikgjiQ9nyaYYEedJMX6Y1fnrPhIpRv5
CzK1c3dLx9HRk2Clp6T4/hyuuUGH7J61f3I6YMK9FIui+gGCHIzINZZglo04JALU
kisP1Vo0eEV+hD2rrShFlxDtdiMulOKAtnTngLft1pk1/sci5zsiauvJNOpHfd6S
CEHOT1510tZ2G4teeDioJeUbKZmdoz9JlZvA2gftv8vLr+Ex6xXY5WYuP0NLQEu8
SpjqRVp+WJa3gSQK4evHMljfTQzHZ/hHFPUJaCZ6GKZkuWdAGthRGJCSHBgXOegu
vdz09yyU8cCE5qlf7876OLfNncR9ppH8qv50MBqpAHYeG+WK5DW5DumQLrUnB5fp
3tbphSqOSLYD5klo6BCE1SWKpiTHfy8ArYq7f+kA4rUZtFFKLVmd0Yka7JDIjnEa
75Qp3pjPPrn/RHzBBmsTw7JzgSSPsRLv8dUo8Lllx0jCTShlZ0ma6P3qyz2KODk2
vJDKlxMy6G7zCbeR2bHg0O9ih9CL24DYvLFcqD+qnFecEk3hN438PrWFNsQE0M03
JffAEOoCfO45gUc3d1AUkIovoiuGAnRX1fX521yiYnx8PZsNM8UcNfuZVGbuGaFH
GWZB86QtUAux0RWvW3iT1EJcuFyjKKjzUT2+eFvcKEVPYGfdy5euQ+Bz0BM+i65g
xjizuNc28P5gr2lrUfm/zZ9z6tHIix3kn5kc1KNKzI3v/9mLHDhIr02kGubIobBa
BXT2YpDwU+XIQij31QnKUg9A0bQx5xKB6i2ZO/l1lehWIuALgPikPmkTePcFZTDR
L1X8kovYdIF9HaRUSSQCiiXzVKHCgy12zCxKItIc0TPDdOyv2/oFRua+QfiDFegD
qv/Ri3xKHwYwtsaztpx0I7jTmq9dMGLUGcE6ApP12yj2GoceBlO/BtrDp1SDHlLz
8yIgF6tIh9/FeeCTK6jt14d7eTQlAjQZ3Z4Rbe29VvK3qmkXq6K2i+ElOIXvOCgG
5hxUmaO3bHwS2/EMtlbDmMKUmzRpYvkL/MANZxNSk6naRc6HBel1rnX6xqAzUxCy
vDsrT+d+F5k5dJHrVUdqCpwdf1z4QH6FiG9xLd+ZURx7Czoi/NmTU7mxQn5fdMhu
CcTlM7SJYtBzgP1sdw9uRnnv36L+WrCq2CyRdr1YX9jm4AH1NutlC2h2sIU60wl/
nH6aQS+StBv+BeoWXeNNahIdZiFRl8KkrxiNrrEqcn9UN6acVmw0KNRnM1Zvp8OJ
R8JpOIn5blQNmj2hFl8uPrkVTCuRPVmPrt61yMW/dQNekiFyKxovEpRLHtiWDJw1
o6f/ErgYNkxpeqsCCGLzSmMLTmTdHYWT/4b4ye1YgSNBWdFV5xQggMre2EJ+P1I3
kO9h4gqm0/A1BBbgnUkPptK7gDX+JbrZQ3KKJ7mQ1I3/E6BEm0EdokSYBh0JVt2k
yda1MOtLALb5DDBhTIq767CrBWWKVaNLElQKRhL6MfrMLx4fGhvtOXDR4qGvowc9
ZY7RGaWsYsuq45pqU3s4swiWeti7j3DVGbOCxtx5C0Gh66v+cTAioAWvQRD4yhu5
DtBnx5Ra5x2wpwTF9hhK8wDAQzADE6ZH8D9Up1TQ+hTr8XB+zJMwBB5k5TJZ/1H4
lhIKL3vPFe9jY9prO8c0amVjeS9ae+6yz67QzcUUNORsaRuYPYHYENgk7M9ZtQO5
NwZ+eCFzN1YlFPvki/THeYpU8LiY58yt1d7/kb9tswdAMNvCUFiUDzDDFL2ngeae
iNWHeC3ppNtxsTc4iywb20Jaca1zYeCS7rDSwV6UKQFXdE+SpUf38Hmu4xe6XPed
fgA1NI7+rX1pxA6W5g48vn/zQS2PmYYiYre6dPcOUwD7jhmdQeUwvu+VU0Z869Ns
hCBWITsuh6c5pyWwSEUoHtWPJJZeztAISJJ5/kCIbXV8TxQbEIxZ4DArrvxX/305
CMkyuBAkZLi5Sf1EPwd665su7B6e3zMIXP753DibjCoyyJgGn2iD3jKeRYQmvpPJ
yJ4XVgUKezBYeFoKM9DtzE8yIC+KZgbSIKaQZt2GQ8URhygScJXxQYE1XfuoXaaa
+TKVEMDADAhIy1gTGEkg94U9SvcwD8EJiN7wPfET/NWjE5VBwdRp3rzwo7lltvX/
/QRFJesakd9rozR+cCdlSkJSBzB1+vGTV0TM/1sPbKHuT+tPE6Il3ovU3hw6Jnr7
EQZKgTyatgrY/xN8HaiS43HOXnZrRMmthLT+IqOyb1zC8k4v9QCdxMjdDsQqOpnw
5TXhOq802FBRAqQdH6LC2NUJJGAPXEv32B6b9HEwakDcp/EGr3nAYsW+HqYkzC1D
0Xdkh8l5PtVZ73kX7ELoalM0Zam1Td8T3zAYKwpgjK+Jx04VPYulMTpV7DtP3QPQ
EH60iHK9tKGDyWV4Omn5WwPjdUZcqWelbjHcfIQILc9PQ8VwzMJ7UbwoSVKe6pnN
7dy2NG/6HDQRZuAY5IC0ULDklapiEb5NYZPOWBsp2jx4/gX3g22XOMShRUvRb53K
eJFAwhlJz1TabCLeKIiaCGNk96uuN8bd8onqAyE+mU/olFo2IoQ7Oz2DFaoeQ50k
emUelaXoN3Os/iIfzaguidcElcgBbVVCkZv3ZmShiyZYHiDfvYhaP9MzUHjztPKI
Kk6UaptYCF+tTKsejE6pISXvzdRbH3qbow3TSPa7qII9Fg3eCV2RCf4eTSC5wDIV
9KKuaZAw3Mu8cRXcPNtddgcsOEVqejsLtLuRLzBnwRES7rQYQPVZ9nVVFUJYXZj7
9kr0A69Qk2ObJ0BqJzd/ncrhwlou4ClP1pt0pbSApXJFS02FuSg4ZfxfuXkOFDOI
RBQrd5jovYYiHN/5xJJRykdX2kyy3VYb8IniiyHHsauMgsYdnCvnVkXz0ofda+46
lRMmcEdKoQTrFvtWtVUP2qjsEdZCGBBTHFavkVnLoCV6PdqIb6RIHl0DvwmEq1jy
D3vPcXITrqGKtCdSoZoiGFwLQYiQmwpHVvnlQ96dUOm57hqEQFVJoYofU2qCAO6w
IvlE1Gj4DYxGbjfhEax9h6OO0ZmpaB8NFxX1I7TslhYoE3PSN1J/RSrivKbJtvVJ
+wzyu8W94QBoToQFO2ThnM56xiVxHZdNS7La2fQrJocz8WsnKz0ae2LcHxOX4+Vu
lprVCqAFTT8//t2Fd6KYcnnZ3tllq655MF8Jaa8mGtLPXFV7NV/sgb49Gc4mCpR3
c+E8x+8vScGVD0NqnPMJnA2BeIQdleWueGHGtPT3JzOoAysWxuWHVWNIPMfBFU2V
nQQvQZ22xTo/hKw8LjhcnSuw6N8WGTHBG8j44Ks/ku04R8+kvqll40STf6KR9Ako
nGs15w1zx3MYXDQELRdUyieo3BHXlkDuwVkojofNCUFwoJNT0UvYCr1TrvFOeyB0
s8jlx7FxuGz5eqnJm6fkS6eLf3/Buq09mjm1mQO5vSZXXj4uXMLq7FLvRx+UZ5zY
FWh+Sqcy/xXMB8buBw+0gEkAigwQHGTr1ExaWIoZAAEKzH+LwaAj6BR2UDGJgNDI
y0+CO3I5q2L/WZ+n9pu0ltsA+BJicZ6GM3qS8n0LcgTq15WCmz/K4jB55EI7YCdj
8PWkeonYxeKgUih/Pv7PMiq/h+AHKl/JhkTW9hQRJTVIBWCgw8NC8vnkrI/zKOpf
zgnJEQ8tvr4AAVpf2hrwvs2uz49iQqtZhXtLohD7wXFJSx2/NVOaJZKAAAbh3CMP
WCpqmLZZHvVVBeGFcUh6lK/XQ9oFoWJcvyaa6ZekYpC+omBwEHev27pemftEktC5
BGisLYdfL/t9rGNLp6iZIzQ06okdBoIrhpsVOHWm0SjqRhF/R+SydbsvthqZAFSA
z3oIfv8niMtcvNhWhmgSM8VIgzk914J5fUUY2l9He1HOikYYKfwTMK717VOUGXyq
fktvoHOd5yHJ+zC/B8j0F06Iw9f/XAMxwKPg4LgHVGIXKJMR7QiSCET6iUUxz+hI
jBs2/TmetMN+pvnNPqIk0oQmwmoQ3a2+hzwjMYg1+wClRR49hM89EJ111q+c5EwO
dycrGmdk99p7I4E591A0iJHqLPwE4lWTSPYA4yP0LbxbqDCQjQ1L6jnSSKuJOlvN
3T92EzSDhlbFQ1Lqo3F1f6z0oKAcTkCEvTCFBy2Rp5CuN8NBaLp80msDtolexGZe
OySctYPkg/F6S0bKP+yHQGi+L8MSZVg+KGbmAXb5pyJufFlAwXdzbfmzU3WyM6qx
ycfut5M2MXVOF50EnCJFzAFcYIg8g7UvGgxkK71TVdJFRHIknwDEyC5BGSWTvrGF
aEU0065ZcUun1bLQwVYX4KT4B3LbXYbB3mNbZgecRog+5AyZJHXUOX2il325cxRw
yEkIlXgv7EbIzj0OZoIo7zpeC6EYgIXBgsIpU3cP8mzIYJ+0wwWcCgoI9BX3uYVF
Cn2SLGBWOEZVnTwGJj0dKQuaZO3LMGU/3EYspvcK8r7aB3Nb7wg58sE8Cc38IVky
P3CNwNkdtfVnIG3drlppDoPMN8UzRH00qodHLpthzohpfHu7Disjk+zK2pjB2Yri
CBW5mJ9wkzRwf9b1+Kq+VV007IGlCdJtRSJPrUxBRy4MKg7WrTuZgM7i/je5Lm0g
xcmF5ujA8UdyEdiifddAtp65/PiBDLnO6ppu2uLBQNtB0Oj3xc9SRQBSCftkdDF+
Ey4pdYL0jRzaNNbQYfr8TK3eGfqcwyx4bCi6B9HSTT1MURk0hzf+KECZVbQLhYZ+
mNTSNri/oTqpl4mwigYfqqFBi+Q4lxar2YSZ0k/MeMJWDkxOFNtZHxvdaevdHKHb
caoEuQV4NPIBPS0Cp3x3WPm1B1SC8vUFOwzQR4n5HNjIL4495VCfSGVVjm4Uas7q
LuMe1yd8Qu5Ccv3pIWpojI0v5B15R1lVnMpl1twiwDTBcpa5HWYJAGzCwjrUjI8U
f06VuIYnqDu8iLjBsyHdnLKlGveyhwhhifnPsa84K3drP59c110ZnhCOcWiFnj/a
JpkBWU1byU5AkKZScMsEUNLaLKhd1mjVkqolQZeoTP1XGHH+pw/mT40oS+h6g1AH
T13BJjwVVNY6wb9Gf+mMrNNhdyTxFaNR3YW3oxkhExK6h3+l+9U20YnAv1WjoCm+
7nBjdiEX94H/04KtOoI3x4VfKc6KSz/ivnNGYCRmWIkcIKtkYVZ+XaEq7IKlgIZh
2aig/UsHxuXQs3pv/x5ga1rQt8LyqAIWau4AjCKomJ1E32G1+ANObDpDI0R3MEDO
bG7lFHMEdjbJr4csY7dd4USu11jhAJQHscpH9mXMNlJyEsjoLlBZ4RhzKawj7OEY
v/mjBmlBMo7SY48KYVtLiVMpeV7QM2XVjk9nKcIIWOaMAtafedPq+QG2sfWfpaZt
gkR1cLAyhBRWQl3ZraL2PbvFYg3zGdhyN92D/vnl9cFDV5gxPQ8pqX+FTmI0pszm
tv2IJL7DnXUmS86+en9PSLulDnjbvfY01VOicO7CLrOffF5L69dctDlXKhvYhWyg
FfJXLv5Z4wN981RE+OITKNKMJxaA8cJyc4TwJa1cpBpjyhThm5fCtsaN5ywK6xBj
3X4wcD4IIPrJDhrNTFyNVKi12mLM2r+Rb2QxiHopENBtR9Ei5VGdwlZK7XriXWOK
anpPM+9fmAES8sEuAe2pxmJ1K1KbCjJnJ0VRLVBdRrPIMO/LTGWk21saN4DDjgxN
/S7B8tgBCMQBMm8+62xDcnxUdxYYW51WOLFt9LgRyBQHLEkinu29txEZfHDaksY+
nbe5WvTpytbds2ZeQ1LDViy1IvW+Yml4r4tS07Gb04ZToRXumGEs9esjmDS2HlXp
tEGi7quUu3udxkb7cVqmcP8+mIdc+QZdyE/hQrbB6X5YOdeIjyEQ7pWZArnG+DZP
F2m/WtPxLPWAoQUMH3ekjdjrFuY02UODNyFSoB3Pz2Kifh9iusaJFFykz7+XyaRR
1iiYZf6AqNre5fBNumrw3tisfzUPAZOz2i2dKdnG96Aydzv3VDIQ9KMrhkFK1z0+
9KEngQWt7PAOpB9jcbT39aFELMZrjI/LWWu5MLgmrs788507GPOCxltrWyfHfSlQ
mN1s6DBbGzA0RSWpiRf4QVZrWLxRey0ED29O3BndV/9ZsGLWtLoB7rmOMLYcatri
XRvCbIisdoG79hFhht5sEZWIX4MKN/ETL3MzQMZGebKrd8rI/naWxC/rYXJFfTv4
VDNlN7AS6xdd61CW+Q/B4l5W9OMbKHn65SJeQszSDD31GJc/wrm1KyQAlYr7IsRQ
eXb5/QjQgWD6phRNlhq2PTtNSTWCzHGBViabYrUDHXkBF1q8n0rdg0EaZoWYuKRY
TzlbqDiYrf2Tw4I+K2I6eio4NYoy4ohL/s0F/wrblbduC10uQcRAEKQVLLxFeItx
y6UvGffDlo7zTLeAwEw9Zqs/OhdgbHxMkm1ucAwvnEChTYLq52MdUVoxkiB7dFC1
9MrwJCfrkWfz/q7Qjxy/CntYmah53mn4ulctpl6PARvuPjC+c9H0vtOFnjA4LSCP
WihYuTqDkOKSuchiEs7cCCPUvaQf6pOKnXZ7uuQEG/FOFK4rRED5dx7hqN/8B2NY
Z4gSjrFxFnADFiqJgNZwFach35MfD8kYY+Pbxu0yOqkzuT9s5AbQE5W1+a8dC3ru
u+QjjuR7+IXP/4ImV7ulZj/kW1U/VMEll6UH/SWwINZR1LoTl6Uw2CE1DAfnIsjn
c410my1yWd3u26imvQk3jNF2+1lfiBUn5Lhqm/v+Pgv6uyikNRigJai7ocRnX1v0
aFmyuX6tMLgSCrbpVwVG1llLDQqQ3xCKPqkdDHDDhYzwKtNCYIg+JRuviPwocCbN
I5dNgYzV0vi+d6l3CdssJJG1AAtEXJqm6m68UeqqgGcBcAeHFBiia8xUXrBAaluC
DRJzCVbN3VzKunO13DzXlOQhrTjyaAsT7vKTrU5l5cPWMLOaeFvbpbhcRmxyITYD
ckznIK/lfSwglcqf/PyGBosxZOfAjRq6+wXPk3RYLPqQUCV/5G7kkFs2MPDmTm7A
hZCA+yXf71yICVupyYr3AGaaxxJWfNpB3xmcfQPMhpt6GNFj4LI9EgbSakUBcnKR
C5skFTTNnvOSAo68tErW7t1ywl6Ks6XKu6Z3bf4wGKdE5mokSeT/NgOzOD+qD/I7
7q7GO8kI8Yuz0V8Fw0YBCjqoG/TucN1yjXRlV3QRXuNRl45PtDmf0JHwv9rMWbP5
r0y1aXKC/OyUnLUfTN8QxtXCAgdRnj2qAajDbs0SIU3mbSVLL23rvEjtizMsp5BE
3mQ4CLzMkZBJJ06ZA3EHC3kf1OoUr2+hGw79e/kYIGDLK9fckRatJ08MEM7HZT4r
TB3o/WynikflnxfMDmGajl9fdlTWuYEigXv3QziTXGXWP+oHvzuVI7WpqpOEwwKt
xVEbtNlZ+TilsaWkxn67YvRExFMCM2PeScUNhpXypER3VyXbMZWVoXb1j0qbb+oE
ZO2QMc6he9H0M91FM2NN3WFmiAsKND/uH3gT2f5vcbCg4gxT0TaRck7eHm6MpsOX
A+1C6fTZ0yjQ9EfdeyUft49pl9+kH7ZXxbnaTdoOUivxYzoldme4Qq6p0b0lSZPo
gXDYphVvhtav+OH1HSL37Wi4FkWdqg4SHK2ptzTDsb+trHCB1ShT9iDoO6qsxdYx
QYkzTW+yKNlyyoFMHirkZQNtHtKRswarNF/+D4SJl3IYUpNEg1yfdNNyvfEpQQq8
fZgjIdPqU2htiIphgUE1wLPBEOX5xksJixlYOdtfvXFQhg2MyryB3jqo6E8nu2w6
QWeVseNT6V7t327ttScEv+w9psRBf305CUYxTVeUcW7UpFOf9o9FjUHl3nfmen/+
buFeX3cJqS0eswrhyTnYSahWsO98AyenyVOPvoEHztl6/AvyxGmhqmPrx9bEFUvB
MvJJ6zmcFkxu5rbX2rHzJah2pvekmdLpXNjQSfXsyba4l0hg9qQ/ZflvISnXy2sd
Vri0kqyxytWpD/nymHXQsld0gclsnCj3a6dOfqyUNZNHsUUtXS+LyOLVP1sYX8bp
2BzQCqYCZ5mbqOMjTSSQD0dmys5qvgyvTx/ssTAcUPH1agK0fGqWHnlNnq2h3A3T
6/dtGNUjxhv1WO9ttO5XEr/NtBfwhM36WAWV9qSVeUSSFUZuXmEdAxUS7a62Csv/
6pOK4jp44V+cu4+b6XO9v9pqgmWQVNfldcIQiTdmKb3GS8cQuq0dYspGKCE7TKpn
lCHkPK3vIGAEokW7hTiSt57vGv9WGV4bcO4jSMqfQnMfmXAcU+r9juDqlECQHb4v
LTbljtA7XLKJVtr8kseIAKMatKOxSmbU1Nj9wu2gjpXTW2LetShyB5uuvkjrmECD
EO2BHftfif0WAslNUONcwRWObtH7heMzv2PKeAeRyTTCQ0/XzL8FeqN9DRYEuA6c
+WVEmdKmsJvF/WmctkAWf75TTqQlcjFQ+7YMo+s7v+JpCk16JlHRAekd5tpF7Sij
Rx98uIuTQP45jYVrlGd1P4lT3iHuz+BlsFS7XznYK+ZNRiuZ+zLrBzke70t3byRD
VgRlUV4yAlJsvhvbNR7hrP9gxQAPer67vFwHVXEU9Nv0w+m18sZf7KoxAQNLHJnQ
gHQj/SyK7E3164DYYvCubgLbyB2eXqKv8/p/K4qzPJWIWiEXZgK7bfp9OsjfCndm
7YXaRxeE3RJPupptnSQWoAWgaR8JezK91hzRj4KdMqj3a1VdOxCjiSpQtaHelEXk
ewOw8MYL+4nQD2Mk0NGQ+O1bJ7zwieaJQ9aYy9+KUTIBJuDu9LXnrs4VHYPXrkq2
TwTEBoEC+ozokfJ1t6mVWFZWICS5X1dgm3TF6FpmxHLp18Cd99FKxdOv29/zKrCW
BqWTcjyhFUE48fWYEoDFtnquSBjvK3cLQFfEoYb32vwcaMFCCsF/grNFe706XwDA
C09z46aFqaoxymIvNGemgeMO9GZ10fH9/x9v1wLr1oiPrXtu1PyRB5wauSmQ4O58
IIEJVeMLtE0tJWHzsc6+bWXSb2i9CeDIs21w4fCyWmIMlp8DlurTNwu/7uuEKiTW
g/lRBd6wfzmI5hOhJVhHobXtwl0O4hI7+OQ0CyF+K5dd8AaPLN6/wTx1GArLMfmj
NSL9wDa2YvgJAgeomckUXix2N37WZAaO+4uLTaFBO2kTt0t9IOqVq9GYXLn4GDgC
6qWtUjNjuJHL3U9RF0XEM1WkyTgZY+l/sUgTCILByZe7MDlP+GrHKBlboO+gtHG8
GMdBQcunv9VMBLdrkgwxsXoTuLwAQaNFxyToPvg/RBDBdNMHz+OQ4+HEo9b5MQpk
rPzMDipZYjVsT0NyVMYyu9JtfiUIsjR5JLicdA0jp/FAHfsWBj1fK+CPRq1vJSG6
+FwSFSOJLMGah1RDsT7BROL4UzlhWxYYoZuBN7iIF/0wug9RsusYlayyYXcjZGg/
1tq3wuPSmVNawlckTWetHXBsIKpermZirinsmEgVfL3CDDs0+D3zfCMEfSMLwLVp
Po3qL8w9wG2yzv7ScQAmjwJhuQxZn0aWoZYV3X+OeVypFRD7bJrlwJqRdCJ8ipRr
DF16vsHgzTUINPGY0+vl6Ug4qAH2j3iSzjOFDxU/hQ90pwKcCpbtm0p2RJBrqb6D
dlyRepmt90nHGc+7dRrejHVUZxNDOhLsngnx5xkaL0dhWKYinn8tgAkd1ZTm6uOn
LJqNahr3a7KNq/3dlnplHIxGIxEKw/wW26yL7PWZJyHuRO6b5gB4SevlmqT6MG+g
YHBgHVvFpsj/Q/On0cSRkX3eTAd4pNezosys8JqgXNDX5Ztc1nS6sF4nXeE3NjmJ
dap3QuEgY0xO0KNQi1e+z9kErzFZ2kp26ojfKusE0y0aJEISUxDo4CujHORt2VG4
wOROKaFj3IyodlIrd6MWFjIe2amu8yOv+lCOpDYw+bkw4rmvA5pFVRNGeA49aF1L
P7RFOAMjaHHwcgUT3JVPaoYc8ECkINeYCCFw1qTcgTaqwou2icIPBcB5NGXEgULB
S4KJUng8tsrtwZLs8rEOwvwlwVeDyhQlJ2nI35IElLDTllsezDzrg0BAUF92Yk0x
Cd4BUymEjA4q6pIvean8DTUrBNnQjZhOaW1s8H15Yt9EhQGFGXnnnhPnN13Yc+m7
/2tJtvz9LoKaoZ+lwGSmkn6NtTfG+CLm0AoRH+1ugc0uF5wpSVKHbvns9bsay67S
lI1aW/E6u2QgezdqZW2heuSfRqb1D8k8TUIEJk3QO+EyWlY4ZuPO+Ol2aBDiiuoM
4KbWo1Cwx2iISe5PpdH2PVcwuY1/TL6jB8r/RHyMow8DMekWwYsVKwlZSOUNS59O
T4MSpu/yZe39I9+Os58/ACILbPdZl6CniEnUQJHHIKPJD3TaJW+ZneTyfJv0ancd
bCB35+L5MyCl8sjzIPgGQ79wdwTU/pFKWTRVLKey02IpzOCnoR4b47WJuFhi4unS
djUYXLDGbIrEOP0WlDNNc74i7I9mv6NZjTThYZY7vTEAVILudxL3lQPJ6McvWi9n
UKW2VPwggnTnE1I+053ou7ry+VUwMsvw5DiJ5QhhkidcaqGiyckCOWzQb30iPD/Y
W4f8ntyj6Vav4QT+7WssiTFzjYhfE3v+tY25omI2Jny3hZniIEhP7jhI+8JzsxYa
EgsrGaWn3Dd2GdUCxRrFMbEK6VHMYDjLhobTUPlZdQF2uOsw1/qFJ30zByLmMLuB
04GZWokRk86E1dVZGCHNxQ5cwaKG/4rKo74SRa+nTnHOffmqi+bfzrJ6AZEf8PAh
fprdvAatV09vsDQgwaJksPkGyzBQyPNPmiebzmNmGw0vrRdeeYSoaBVTytiQQ+1K
4PjsHQHDYPs+Ec53JB124ZB0MHxCXEg0PucWMol3Od0pYVbiJDR1vTtke3uThorJ
ukSYt4aw6E0h7f77joFDvClHSkckxU2CjqeVNTjIcPBDoJqz2faQBE0uh1xBj8PA
R4pEtCrgs44LkBPhGweO+7CzYyr7/flCgQ1WNvbtge3pMFnQUBGt/g3Lek/fICgv
NhEWt0PoRTgmotbVIKqol5JYy3AEZQVEjJjlBGs+VyE/cmTVE0A8TD2V7EIsAQWd
KHw9PE34aTZLbR4kl5J2TjgkiN4cmTZOasiF10yOiCTcanY3UBijJaARXVi5Mm4Z
HFB9Ba//EDwj/zpDw8NEznrbUZGysSpxFnLeofOFGERmwDaCHA16XoRfWIhCsYWC
+IvdwqcMTdXIqaXUD85Pf4KowNQW/qnPQ/PjUqsav/qHmttcxD9WiXBL7Xoe4FEQ
+LpPrdJLcWR4VDjrGiU1wVcFOHc/Zawp3aiW3GjFZ1gmHrHlx8zy4u39iVBJfk76
SmF9UrXXMDtFTvAUsF1MxDCq0Ew3Qpm2r490wes353Mp6h8KJSmIyyrYA89s5TLI
LMPDF3wvWeikEyeB0CZaK73GASfuFP1tOk9UqcFN/btBScIog2cbIXR8/TM1Cg11
Op0IJf5ZB8GoEmbPSdf/kvZJF7uMfl6mrfAuHeh3vX/Am89UxeEmWI6O1msKdM6m
yrPrXLmm+vI5nqpI+s+yZXBZv9QP8y0ZCCPEGNIILfTfOd+8zfgdnN4ylFKw4CPI
fRc5ul8jeExBNWDXU7COEdfwUdk4Hlu3OAe0Jn7f0Z0qXaLA1+wQbUGLwIr4rAkS
X+wBGldKIWUT3RbFIP6XTDQRjF4Xond/qfDWatRYeVcwJaGRz0iBFK9BgOwl/xFf
m3+sr/gDxjqPeQj2z9Ay9BezNPHhVbnLejiMqxbdpZYGP54InE4A24LdDlT+4j94
yLbF8YuZT3lJdx7p599TJNYElsae9M+mfVRmu0MAMA6yzuoInSNmJql4M/pYTuW4
Tt7p175c7HhvNh1pU2HZUOzm/hjkjHMw+YvCMEKDE917IFm+DWcz1SkfKg7KSMxO
LAAOiag2FUyFPXC2UoPw3iU2uW5dKLtWLJDd3PuMjP6+8lJUyN1iiHHkNHVtKDA9
4s4CmU0HzfEPUZRKpC/BbWm/1POcPPCgF0lfzQvDL6ClmMubjla//zUbm45BUYXb
4894aS4QWrBF7Q/YDsfyCLUn9s5piaT/yH18yasVySg/P/zcWoFtUyStXwUA7gtK
+AgAl6mzLlVQVD/GDDuBOd8/+2udrYKUbgTIiz/YIg7UG17sUrlTMzX7KUZgynaU
z2G028JJW+2xP1m9QkmX00cZ+rCOnGI7T9FbwRpKDtnTshASJgFWOIHbMzAUcmay
s7yHbDuturVzKVSkcwia73fT/bX6eu82U5g1Z3sy+Uqvp1PgbtIdxb988SPeRYFz
6+ttsEskWDY5LvYLuB01c8+ikSG5xk0uMu36m09wRbp1nvzXg+J2lioTp3/Rqvrp
PwQXMbuwDAz89iOPTH9eiVUXsHXr73gZIgb3DxX4SkV95FQ1aPDvKXnNXwlXKqmR
qQx/PrC6sSIfpJ0zbcjKmCHwUBr8/G55/rpe3DScTGX3bDCUREGqivyqr28N+WBt
TPlk1k3nZsr6vYH8dBW6bfli1jrZ+RHabKO9yrb9EyeilklXA7A9afmDoH7f6UHX
pXzooDhE9gIcnfgTtnLfwgi/qTSlgsFaZkAruFOg2s2+EszbxtC8kk6XUV04+Mm3
WCeeC5IYAR17bsbB9IRIL4vsVPHmx97h/Okoo+Htuly0kNbh/HpMecPg1g1k+hH7
sUyZqeXZVjN/lv6Aquj5KquJxupeDo9r7SxVvry9opPXXcKnscmt0rq5NUwMkdfE
Ol7Zj8DJ6261M1ZTlQHQZl3Bibr67uA2oJFugOPGhNydqd5yp98IJVHLd7MaIipB
BLGtrUcSmi3bpwepgHjWDRMKtnEum/3C3Y+HCA8srWmeM3rNuCc8dhGeeugEiGbz
1j9dJ1JgHDAU4VkG5ecfwJD9lD69K+9OrWTHj6u2oAS8NjZmt0pq163IWr4Fb/+E
AlajDPkfVe9mDBbHBkzIY2BFg7hQRCiMDUnOw32GeDAT7y145bm2BkvncLAAbQ3F
gvqZ4NHCi4KGlWGLPdMRVwNPmFG2z7zLK4u66sji2NX5aLyMA2cEgXRm6OscpJs/
dogUlajb3pzqpJLWrImXjmiVFsvKUhZBGmt4u+keXORlOyi5SOcqrpxk3+BYYimo
BncDqQ3RBNiHD7k0zfuGRI9oscW+q8/Q0eVgDQzc+Kjs6CQ0po6oTscDkD5XhkT9
rzcT5g+x9feQ0tAOECNcMT+NoChwnaorI21k/jbTfcePgCu3n8GZqMfyjxbSfZta
CDr1MjvRzhb+AjuR6pdKSbJXc7QUD8ixxvw83JpNLEmuKOaukLdolK/Ib9qzpOa3
w2Mj2gYhAU++o6N7TadnCBj7znnb0gh4k22tHD0xrcpmVpSdUM11RfygiLTlZVAk
6pLRrPdutCpqKoFaN2MEvLhyotwlVwm0i04Y9TxQrzVyNPyLvBv07xIK4uT5WHWe
9CtliMrwfefCNhEhvkCK4hcPyMAXa+lFtQX7hpb8TB6z3YE+f/IwwNuhvup+I9jW
qvTYfJsH/naS4pdnGFrYDc7F0JKCON94JisnGEhZ+1YzIQRfCf5CJo7xvLD4XY/Y
cmmtJphyPMerTdtL0r7QKP8ZUOA0cYVEuy45URK7hVqMJlVd1G2BZDK/AG5W0jtV
sx4efBD+DhE3vX6UPiI+h2kFvQqi9tbZVRqQYUG8vDJWk0nI8Req0WPnFa/4KhSX
q6z/yqZGhp4ViZEBQMJROpMDMq8C5ntkwYkLMTV2tkqfiyP4Ct5bPVFexC9AsmnR
5g4AzGFIcxhnqKNtZ6c7cDjU13RCZw3/xxoOLKtR7NS23fQ1wymccA0mMd8byEWN
FbtDXbM3AhBIFwLPGOwF1J1nFiOy95K5fV+8UoeAr2qRmf9YNSEBTiz6uf/hoP81
Yu4yZG7vPtGSD43Npvsvkc+fV8wmHjyRZe1vjjYQlUJ6IsUJ9OU/yW54U/tosqks
LT1HiVLK8ENDhwTECf4G0NU62NoOw7w2NbFOVHP8mUyR9fU1IWRdL0ObJj7tPTPQ
GnVD1hAHd8gZLUBzUcUjfzm/+QFMewuUbnZFhZKBaigdICbHXq3Hd4VAmKQ+4tVx
Z5/Eo5jrJD0aZBvF4YyGYu81tLibtolUN3NyqJF8IrbZKgUdPcsROjLQGjANmnRx
HtpaB3J6P660JmnyrxQHuBT48ElRWSpJZd+nIuWGSLaDxxlHL3LX7WIYTPq28/+y
gemR4yF9Ac52P5Jx7bTYSLvWUsVquzIiMdTdl/yOLNPNR3ec2q68arWNLsw5OY9X
sxwDoR+e8wmqYIXoPWHz7yiRwqG4QcHcspK+ONjmj7AADVLdH6RgnOWKQ62U5Nrj
dXASwIv4afDFNsSawI9diLF4o0+VizJ42bj4vd24hSKmZ9sCNb1oDd+TRae1FG1d
6n+dPmgD8wy3wayx8l0/gHdANTlw2PLdVdSQe9uoeqAFFtrHpyWBLYZqELVFAZuY
hLHhj5nbUVATvL0VngG9we404MCkrog1RKWJZn1ayKgmLKXNA4iZijmqqoqZQSBN
IrjVXxpFA9joeuIYURjYo4R2HGryy4gTOW/ZDp3dAlilBPQFx5YmOl7hL0CicJ0U
zlyIx49AH/aYQ86mfbGhSweyZspzc68S4i94P7DdKk4zDrzPiEJeNorD9uAc72iq
OTJpra0B8i1ElR6taiu8BZngg3LHrNxNtg1Y9F37f5XBVQUx3Sj2Fb2fn97KldQx
rOs7aZsY9IgXJshl2LC2Yg7OsloATgUxfpjtSHDkDSdMiFg97nt5fgtq7jeigAqD
OWR1RAlEcxw+GIRMMsh4ZL/6Fjn7q4Z0bL4cIid43cQQ589m4j4gnxfSh6rmXGBf
FbsVfZu3cslWjvYiM7ESqWEWH46h+0hlUx4d6n1vZjW/HYg+rNp9y0s9zj5ptEkX
QSH88BBgzm3e5OOR8T0nXRmnzHUGnqtgKh2Bpfhx4+5dAFHgW5t2mgesjNlvQvPh
SIgWm/2se3JxkwAFF/jUJ1+eAOV0JnqJtCYZl/ix79z8vz1zMs8mrrw3N1ZahvKV
uEZBKUEA1jSMegUAL7tDlP8Sxu00QJKuiulPFOr0BQc2MvdfWVCMwsnOadJJjdAx
qakOgo9gE4Cfj9KoyIbve4vFcp+1Dc8y3TOXpGjgDjLyNYp+szaGkBCYAhUaWjWb
EOgjldlVRJ9BvJ13ZsBDdezubFrHmuNZf/3H3XtZU4K8asJRp8zu72A5fF4rV7b+
QHawXsxJiZRrDcdTbr48bModTkzQWp2da0jRw3+xKQCe+bvA3GXzFbrh8ZpsAGVN
EqQ/oS0EWTodccqIXEU19xp1uyTSNZ1EBeTG6F6zADMV0tc1F2S9NV0frO17EbBD
9brFBQRcCym9qhOvhwNR16EkXo7t2yOWSTWiNG8rbIqYBMJcKkkIDgJgdah+rY0k
Dg5gEduDN1ytfnkk+xbgkMHcAITuPMiVtsvz7tN/T/FYrlVH4plN4u2IGnpvQuUp
yKrsOMN3bPycML/0ZNxIZAT28+FQIrgewX4bCP8OA+34exTnbQeEv1Pxskv3ilTi
k16ps4zhWJ+gYV1crO4Gy0YXPAmX/dG0qGWIvBKmHHs5l6n/vpZ4B487PH5bEePo
CApoBTWMpxtHdiNUMsc7L4b3PVk3zPRY8ctym6kAMcq1nDPbjhM/qU6TwhUCa1Vp
mCP3msHP58ZpnX9VWHJkGvWeinzo2Ofd7933WJ0xUTe5vbr8S4m+xB5PylQxgez7
0Vcwi5c2Lue1evGzrYwSsuc1YL3atww02Vje8xccerPn/8WGkA6D94C5Ce/KYEL6
FyTB4rGdUZ9/uqdxxWvtioyS35CxJcGJpPpfuAc97U3ALoi2U/oHbPXRKyOSrB3R
ICRhwt7eDgJKdeISKPrnhzYFgSypo7YuYaMBh7bHE5D1OwETcY+DUwARgWA9fNaa
nxEzhX8XcwvOi/CS01HPt/p6GOjZmUriH2LFOqvPovbvCFMLoAhCNt4kA5Q2AYuL
K0g1MuWpVELLJjl6e3eLcpmgpeoQS+vuzoo06q7SHAmBIejc8tKTdsHDge6kGHYo
oksNf2EGThMna5+AkB1M06EX0y//CPnVnfNRwt11sROzCGFJXwbHIQvo0aWHqXdW
0FmRegoNds/XwcbsUfUNl4252ORv64NrkAePDaDldjLQ9fDlToAU7JY+gZ56o4G5
rcxTQ/Uwb0jjwMXN2qKRnwSKSPrwZtKTBz2NHewH1vCRpY7s/jebMeDCa4wi6hho
2kfGR/GoVoRm/ECPEDGZOpSfJxdKbEAxlrEJ7RvHAT2UBdEFSYcReuKd/yq7kLGK
tF7DM4Uf5N1bFxsx7Ih9qwNMn7i40pZoIOuQPCjJqL2whkJWivbLjyK43fGs1QeB
GZmbL9yDjF6vOj3jDCu9DQpnY1YCayF6K4aLOMoeGHFrnJ/6AE4MgQ44RnT3gEFT
DJNoLE+jtNAmLIBU0gb4iJgbcOuH7pCD0CvvqxtbrmLRdlgTXs2ydqiVTafjLioh
Mu5HvlHx7iQjeiQV7TC3nL/2oP8lpkflOH14DN7xwLms1gzoENmaLrzA5EggniTO
onF3lnIR7oXDT4FI4xul3kudMog+tD/Cxl+u6lulmmfpfzj4WCjk3szq73KWNJg9
fFeydYvsisSU4odFHTRlEyjYIK9s2GqBHmjlJIt7gti7wnFSvb0N7lnrQbXDBwam
1AP6/P1udzXqR4yQvhUxNe6QXYIdlN8H3w6Un6TBlvmtpz/1Kf8I8i8aKNJngEDs
jdV7U94iYjWvekn8aPe60eOrISGReIir6lQYjxRSsJaOQ0x9sMZy6Ydn58ePVpbT
oxcKdPCzy0zdcZ71DFRe5jb43HwWx0sP5nlKBQC35zDQZ5PRT3hj+Rb/eIsmps2h
rUbWvNEVYB9MwTFTM3/jlwjpcI7PX8zZMBO4rFiSYptUfsVx3MRXcM3s2miH7tqM
XSpAyobjkfFeXh/OcDKx+Qu/h1S7Id1zsZOvirJMzihlLhNeiE/VmM50xRvgv+6Z
HCQcSJEITLIOcQis+0zj+O955+iFC0R5FBk77FoSSpZXr35uS5QXtKxR5zeo3n7O
jsB6duPD39gVP7fyaAa29HrIdvE72X423yY0EOI6uwAoUv9nk8ZlGgHkxcPVePDL
joXgSLlZ8+03rFSaW93TvJVlhcjtCSPrRnNTmaclZIE2747hc3+KPgc+XQBQxFJh
I6lQNS1tNyEEtD7rRyTusX/65UV6NdaFMfsZbysoBmDzMw7pyttBAHhWGW128u3i
RNItnt+7qEAomcZFkRAn8+lwA+iOpWyebcDPGg7WaAd3etIebmdK/5So5ME/MlFL
V1qmfB2ACl+iRbUqRzS8zYjiFzu1x4Ba/ZrDjjf3/iDADTckRjjxe7kOuXEb4Og+
8AEHb282vMYjFTKR2m0F8zf74xcE9Vwz+/WuHqqYD8Kx/14+C55NvqhyorccniFu
+5xb4Qf+xp+dYdCEcXluJrplXDIi+1VJeqg+m/cLApCZEEHtWKHcVhA7zuQZmkz/
N1hutJ2zvtlLHmIUJ/s9rluu/qJaYT/fMC+fscWmGiivGgGs+xAIJJH2YLOWv1fi
3mXDj1XAHI/n3l/Xek8KrbMMLmg3OWIB+VRuxCcYEJtuj8ojrQufFrMqS0FHl3bB
Ca905it+jZ0qBWOwCuneykGYHmiWDi2evMZ8fmG3FOTj7hI8NdQqrdlTXJnVVPRn
2FDG4rlJLSx2DP+Dj0KjEvSuht2cy/lIhuraFTN2am8WNVD7fLR0up3BvBmRVcH2
YBENkRmKc5lWlg1OkNXPMLCrxESsR8ZChU0H+1522XzmaNE4ZqD19677O9bYkRI4
DgL0FubVwAkTHKnLCYWEAEN4dbv9cBM7dQFS8lPZhpWjM/wIfX+OUGxJNrhU7wDD
kEuegmD6EIFPyUu4TAH0MxkLgkrn5VxeLBkpgqcrggIVjGYVWHh1CStMxMaCgKMm
i0XU+wGmy8COhX99gVlB/7e6uxHHYPliIYT3t10vTBttoZnBvfoYultpdI1V2JDv
cj05GnLRvMXXtNJGzlnPnWJvvmuTlRz70v962t0Meh8OPgoqBTnuYECeCATfD9lV
QVj+0psXT/vBaibxfI7JsjI0yN/zFBn+bCuYTjsOyPUcVCau80+bjnkurajeem9p
oemuYLk0MnU3rjFM2kaHrMbQ2xxH/1yiCZAk0ECoxZXrYpiVj0U9J6ateaNlKlxG
THpBrx8cFoevPimCAyU60m6NUFisil/TBk0T90L2IPEsM6XZbQonk42gGb+9zvq9
OvM2lH0+LZjfDRxzhJwYKVF/JQ4vJEOREyMT+I16onSisKBnWWVhvQNE/r+CQYwZ
ENf4AEldMPNXfHcBSbzP1P+0UHPg6wv6LPMcNaAC0paN2co07Q3YAgsr7KeUQUU4
g4DyM8PIjBjluPZF+c6ru4DnrNWiob47+iLHZCp82m+aZx+hCwwMWc/4GfBf36lt
4+gy4H0TsryN29xEJ0dJtB9b/RlrQerQ5ZUk1qxJp35amUK1ji/imQQsC9Wp6SUB
xWp8I+XaTILsAH1Yf2rqR0KOZAbhltvF4/ULGBeJTX9LkTQuugvgQdTZYNUpiJx/
f/8EL5CpH1w6SaH6M2TvW6TA1jvSYMP2xMYqlFykGoQ3b4Rx1v6/rJUrHrv53zt8
H2PtYxbx0FPEQXfbNoTTpJ40fdZ7Z2SYNV8lDVehq5rhS2aNDN23SsEpSF+gz8gP
nFNtXU+bce0TtOVellhqqqIxmLnJuRszHhOUJcrUalXmmQQ+9RbJBLcYzTwdQu+j
8b4RSo59MlI9p4UwOwo6BRkKoG38ikfizPW3H01UyqhkBCcVptykU47+6dRXEqqD
7xOOBKbZ4bPp8AoPMrdLaCOFOLWh4HnPY7/Ujpje7UP6x7f4uJ/vAIx4pheGlTVB
755s6hkt8JlwRmAbFP54xSd95hTOswwxZDoTrRR8VUgK3n017EwqbE7JRXOcKvcf
agQNdNF5yQsQEtaEaFDhe6GNFbIidreDFlGkLZGIXNqL+BLLSK9q09PLgeLAupH6
BtoD6I66fVDsPt+e06J95YPgTjKXatyCppVzENsp3P+7BU+T4n7l1FHRy4hYJE8N
TBp6z78E8y+GI1que9PqWsZ5DN2T+/grsQ6Gl/pAWXAa9zMtyciu17DFyv7yI3/W
Ddfm5AdZst6B7JnWxu945XcL65uLVY9PblGiMk797p4MAlZHcU6cl0nuZKkq53Hm
f3lnA/lKcrDVx4SBphOA2S0FV7L0+HUMzYdhv6EMknpwKboPGlIRAeVvelFlDGtE
hBTK+/Z9MXgGCkdi1XwmY1xO13Xf6BYPu3aPWHq8+w/oxL5i2nYhunzFYnptElnB
65Q8JlkdnFUDNvkWnWorpAcuW0n67Jef+dxIRwkuKGqxlRwgRYD7YLlYei5jTao1
rNaqcQt75JyUSjpxm/0+CH6ZToYgQMP+IwjA20kEPCN09RZGci0QobCP/TVQYtT4
dPcIjDbd0wn+rcKfjDWFLoIKNX4oc9WQdUTnJLjPeYZGNmRcOXQIIRNsHSQpC0H5
NAnn2p6NW13H8ehQPV7g6ZJei6I01nPcY5dIhBJgqCWgZJimqTdPK0b+fFjSlTIi
bi1xtkE2qWF4JOcyuC3SmjeNv4MDAZywT1Gx3h+UkUeyIXBvZnkelXHmCl0DY3a/
CTyxnqnI+NI1CqdT/wD7aGo+R+oZZAaVSj+78Y1Fa+h7afRRvxJzFHWzdHSHJCnX
S8+fRWmCOyj8R0L//6x4FhBFuz/e0lSYmitCgZt8MN29y4KXeaBcVVTZvkhhabxj
orWrKOqFCNeufNxP41KiLC/4CZA4ZGDkNr8I0OA0jS51KvZelBlRtmPUGqgteJqS
DDg3TpZBvKKIiLSrME5T5i14f1WUNDNpc66GHv3gEfSwngQZw09qPWh3gTMo9olj
c294lggLRoCUCm9P38zHspt5XtNFSCBkeUleN5aVOb0sjZdTnEERcC2A/BZvViWN
mlTwIFWHg/gMdI8x5+TWE1zsZqUZk41wIrgRTmeyz1SWCqE9//S6NJAdNT4YmvKX
gujAA1g+iXHOrnnaiEmZdR0g2jReTj/n+DXBXehq/nhfNJ6tQyrZwHvjPy3A+/U7
0aUIEk/YfxdU22O1o4/McDvGoba3U5o4MhSN1OTxJ/kWuXPgIxsBhEIawFiPNOIQ
GhBPb1auf7Jx+DQSSN5CPkDDCFi+DNmSN1Crp9LekMCS70PPDGNFzWk6XZi+1n6J
xfaTXrVzijR9be7E1ds5Tb9IAmFyiqcEQUyivFSQPNkrDPJsByuPsRimEWvWwUfv
Zo06w/p1XHgN8QhBsdZKCC6f7aVjWfJC8AYkY+gdjndVfEjmXIAEWwVj3GqXrIb0
B8wM6Dog3xt0SXH9RBQ38wOwatTRV8yFc0uwqnSKivAgN8+9hjRHvaNM06mmUgUs
SChnZyvKXVgbXwqeK7BsuyhzQm1CYwFPSqUdZlaR0WRG/icoDNLcktufC2sgBhC6
LFmIc1iYEsB9GaSg4gQfQ4x029wLJQmA19V2WNqL3IpfOMPsKtAIYYPjBbFfxydT
mGAFH1RFIHJTYV6MCB+L+UqgoTeS4VFVYZefe6TgPW5UmQ3FcDh/2o7B9Vl8EY5d
iek5RwqsWAlDewDxABuhOyNfnCR7QJ8E6NvabMskyDIdmZbLAtMt4IdSleLYIw7Q
Wb7ARbGc7/Gr/qizmmtBwTHaHgiOnpFu4nIgNT06HLraBcX4cWMtqleXdtrNbqs2
XctzVr6t2QzwF6CQfbH+o5UbmgN2W7WlcT55YsZU71qYHlUY1gqRBCzjqf0JPf2m
kOyEmT39FV4nfl/DPahboBvyr7r895t1ViJiVgM7VbTWthTcBPIF9FnK/ZZVfpfq
nEmgx/tuHm22DEnH4ub8at1kN/0m0iu6Exsy7ZwakwYcIPuRwxkPwa2mZfKR/JrV
ey1mzantQAhPb6Ohh52mIFxaf2XeUk1/KW5SSich9BLk30OvNBEllBbrC/rRPe7j
XySnJfzHxQdEkAtUWQSx1IRtWrGAX3cwJdDrXRB7saUVhnEBblx1Y1HuaFrvhw/v
SWZo21ehKjbGM1xUaG/dYc5zHQrMHuWPSvvGVtZwmlO2lm635QqZxQAXAr2f+Gp6
0nSC5/PHN5BtbfCdKIqfI+dJLubC0m+muajJuxcyvUX7N2yEmTZ/mKaCyO/nlRHK
P9r3+nrkivveHyplBhHtDyt9yVwfJkjfLDDNl+wiZ0lkgFt3R9KZEsaoAucBwyxg
woVI2G9b/tQVp2FK49i1mxr2kNzVVlvkBqNXmnC9SjHrSGwO/EZWWSL/AwlreN80
cLg/MlhDUMMlSMl/e1pFFIK4aamu8t/xl63N92GmcFMiktALrtFrWszx5ZxO37VK
m4aOjDwxQnDKr8pQqJqI2/Dh7jGhq9wnam4p0he4lLqVvK9KX0pl65RdLf9ohy92
q2D43jnCN9MRwxDBoTKkwmQp7Yeecmwen3T36VBlQzSWve5+TrBHdp9bMy+GABLp
mB/3rKiJCk4yIpywrC3CJzvdBmgy43SqyDsR3bwwu9QVxLyBXSt5Nr6u5vgHTIH+
R83gs0Ps7zo80+M4T8IWjmt7k2geS6nO/T/n88ROVNG5adDQSoD+c4+esfQ6PN8F
j54MS6a9cduSheSpLT5mjQcnvf50UocGVAwGyQP7J8EoNK+OdoEn+AeoriZT3/wf
Dtdsf4ye4d/6eWw4vVJMgZPAfBXeuxO1yYiMHDIBF23oc4h6sUDLoD7XDO2cwzwr
cqR8at5luySWjsC8LLJ9nurMklq5O2rawmng9MxAv9Nu6l0k4+AzK6gMDxaCCsRQ
L9lfzSvo6W0oZ3BHj+TA9XJYnTPHZ1CKm62qpe5Z4DXzrmHubjad9QQP+/0ZLmxO
L7IJpbqoiZDPZmKYT8UDUlGmY5Y+mVzBeJoaXoH72o82miLNJdIjdERuZDcqBnRB
sfM4wIhvW6UY/DSwgFtrkGm7QTMa7FvnCUw2H7gT7fRYRGiD5ah5pQoWECsDf2cs
mnphWKa5stw6Xpji66yv2YjPZCpfyYUDMIKL388my7UEFxofNg9nbiV53YaWWEqP
gJNCqbMZculbJAX8JczgyQK2WF6vOinpXtfn0jcE8Gm7xNywg1/yzA6St3NTIU6B
t7s0Sm4/jGN0+d/LcLYt1MplHmn+TuzS/+OBvZ+uOdcpz7O7w7+7ralNnXiEKLZ3
Z53CygSuZyAkKXf6gX/lRFD2+H7/Z5tRzJhyMjOxeLP+eB486m/i+XX4uvKjbnhz
R+/F1AxzQoA0mzqBBRV/Q3zJMCoWUv7l0gQUEimgCiSUU5994AIA/q4cyy1uq1P+
O0jbNwyBd2+U25xAgvdJ4BLC9TOJdoj2+RGaj0bt1GhBGFiRsgNCeM9ljtD749YA
Qx5GJwLFSmPz7G8/3a4UjoAnAuHb6NwsnChjNqwYXTug8pW/tzVgXxqgxnk8bjdP
rK7iouIlfkZXMsSy8V/dcTk7WoalMXVFEZZEj98yjpisPR5ZIxqMHDOTJZ20TYA6
zkJ+KTKpktCI3SNyVSoylLz/Idjb7ZqMAZXkWaFuoeD+JhfKCU7p0dDf8YKjTw5n
alcRmxCjwgc7dkJwBKNC9ICEDMErbTb6mIEPArLU3FF5yjvmf1fxkTUiVzDqUCVk
Ab+zJzs98RQkWQ73ZTkb9/ihO+5sUqA4VzgBUIULSEyGsqWvwNzjxG+gDUbwTIjE
un4VV82hLjokyZFSZ2kYhEDKtiar+eVV1SQu6OuNmCXUstaJXi3XcsE/qYf6m82R
DroXeKp/qPnLSSI3g74eXYKjr+xEBIiXsu1tsS15bF2ZHCNFnf4MTfhLLcJDJ4hi
AS/OyCqb93Fk6/+st4dvjW+e130+u+Uq5R6rMbDbqKlm3TGbf0afozXfese2cpPE
pZjz/kVd4h34EW25mE6uu6loue+mO8l7hL6wyT4MpqBoStsk9MbKmIZZDKIat0tO
hWCm3AnLLMd+67iqouz3q//ZweFkdvnTohGBTsaGSP0+sjqwdNV6uuzX9db7KtEC
eoBlH34+6HnkuqmI0M7aXljc0c8vg6kfrZRHDqTZC6k0fT4KP+mW5sOAtOS+Y7ou
A9O5JwKLskESSlcqRtG2c5zdfBPBWRcqtmoIV48PQlH7YHgXyB84bgfUOxp245x+
qF9jv85fBbnF8rHRd2q6b4t/fZlLQ0xYmAlCmsUJKVVXJqJJIAcqcZon7nGgPuWT
sT4ErhlLpvsGp40MMVEflPu3IZNF+eaQ9O0HHEK7Jb50cz0RaQ+0dTb3f5f/j8vN
ZhcBpfzmYjp6DOfQp+0jlodddLSN9g5rsvt5TNFC0cI1RbFhdzeDxC2FuRc0Sosa
+zPvL+Va6MVapikqpCeCQryplwN7leypXwKCXmn9tTFRxXaVfHGtQ+UNmRFPkf1o
1PV8FGOQauQDV0Xvzu6Dg14wQnsD6TF8rxPvobpSvZolORvfzs6p6veuvuonfBDX
cJCGpVHq1jbyZHW41rAALdxMvsrvHJTqAsIGQiEDw4xpUJ7v9Kq6b+wQlHWZW72C
NQhNH9hu1u2QquLIe7h9RvB2t5C3kKg9k4K198GlpPtlCifcLkyaoqWZev9Bb5GJ
oDvq037tcQBq+iDpIGJbd4/Q8Bp4HAQNx/nko7Z8h8P7ouYPlKISrPWqbOoCZxLS
Xe18ZtxgKvt58hNOlMpQWyFaMuwdSIjqbsuH2I8hVl9UGKK39yaeaJ5weJDNnOXs
e1UbrdQP52iyE4ub4bCU7xDeve786NAFOx+2+hDR7jQQ+bwI5CJUBeGpCiFICaDB
uBAUjR+G67qOZWpCAKbLtnNOUYdvLVbf2agZLpkox9FowVCJhM3gFDj8KbARXBtd
7JGI+CYRKZHXyRSXzH5cS8/ZMVj7jmXget5Ivjg5UsXVUVGzdOa1cJexxvNk4BkA
bxup+ff74eZbsWqJyeNt5uMZ86IPFAI9GdxAVbTTzbnBwGHWwbYycdLkNlybLjSP
aqhl6Oz79Mj4TRDh56GM2fKRoZYeF4w3VaWQVr8lw5O8igxWHbpY5AqkC49XPHlo
ao2Wwdfj22o9VTeWkLc4apXkd5st1BGZfwkcR94nKvDXVCn0957AeuBPxnSq6AIv
tytuDnJmQy7CyJwMeXzA2OMO8b2anqRUisuuqe+OpBSJ2FLyX1Tm+pzGygrB5ByV
BqBykeZ9H0JIQTmO9z9Jdzsm3m0cmQPS6OJ67bQrp1iK0TJduKmua/U35Z6XhaJo
UKrDQUIrGqu65s41UfnmfAtT6BvlW4tQLswNSlC6UaQULVW5kWmLQOMMgvzIIi5i
TcSej32XIeXWkoczQeEqEDJ3wdQYkEPrmejD9wbLCfxSTM/B+ui4bvaOY0ENZJRb
k+TD5v8iIrmVOOK29vlW507EFzaqYtyD4/jmL1hvBBwo6wuRGPqL+RGY9vJG1HbZ
4EHzzO12jyEMZxhurZ+2S+e7kfhb3D6kCfsbjzXcWo+rgsoZ4I1PELuNeqwkFtI9
6WUKBcAh1ZbzM7n1iCTJRvu2xcUM78L+waPDvkgUFZgI2k1Gz8pUILzuBwTE+LNu
G5Hg/VKWTuhRlL6AdViBRhD/OLG+piOeQnxndNaUXZ7jZ2TSwLCQfrd4m0DQnxfy
Sm4ur06XT+RVJkkJAlleg81sanj5wNON8kBSXj4ZEpH5oEFhWRbE+1gYSKo5UbOs
XZSBXaUakA/hMI0KYwKiV89c2/MdD0FdnfzsAgUOXfeu5v3HzQK0X8fesJ4MyYSi
rFGoOfiQb3DyLEMPSfzblYkO62QT9kOGVkS0Xf8Xh9IVl4Hdf9zTkW36dehtF30/
i941ynL4zvkr6EJkGtfy+0SYsn281mWuYtXqbwY2ipSHT4x1dhVvmr1ifhqUQ+TB
oacWCMFWBnIcobfRxTvq5Qv7MpVrCA1ak3vns0ZSAOxdKCKWtsoPw06WtSCIP2gS
ISJzSiE1OiPeiDxFnofkXo6BIxwiGyKeCXcogPYJVIIJAfil7yhshDYb4aKE3g5p
eK12gHXzx4MBYkf0d/XE3/FqPnvzNfxtpaH7RxYf0k49bg/a9cOmsJ4a62pL2rPR
XOTyS1TQ1dP1sWFvvWzGVQ7afU4VWthNGhP21UPPt04rC9840ndPJ8Eyt3Gbpo40
MKtHanh6w0w1FmGXWIkmD1XP29RfmS8j3YDIhkR0G6zn+kQ7+lM2x+onS7NLz4Nb
4AEqswK/MLQSYMEC6rukFkI5WHS5VKdUUMezfxMkDG6P8+GH1Akr+lEHS4xVlDUu
a+vGbeNcqrHCnpFFArju0Y/8NC5npLL7VDadbNQrwQ9CW0SJAIb7L5ZD3lFdidBl
pdkgywKQW3aKvU5nPuxWnQQu1eu+0UyW87SDloGyg1H4sZ+VcPZhYKM9GUCbGkYa
FfJqYn4eL0YhtAYoUd7dsK7Ipl0csbyxk59JftYuTnzLiJ1xSSRuLLzTKI3C9l5u
sCPTFortAxkwOEX8WWY+aNjnqixN1/E0v0AFlGT32WaE7+4R7W1rGOzJpqo/NRwX
Y45rxoNb5tnKtiLjzCE2Is2kSKy2SHeW3rCkqPK/81HzmF3bLJCKDYMA/ZJ9bVBE
rHwACIquXmAM2nyQ39FL5zQEJgPmY515oXYW7qfg9OT0mK95a+rqFY1poiElwdN9
vvVEBHuUfl6b5N5a0Rl6ND7To/wrlR4MFREuDj1m/3r2kclEaInk6aV/51AoWYqM
3jjORQZbSv3xKq7eBv7iouo9gabR1wkevlpnbPVYST82NwqkwyC0REyZCh9mL6Nw
Dnxqi6lbzG7q7HW4P9On660YwZnGIHburSfs9p33FB6FNZnnHZT/MU/i6fc2PEfV
81uQqFtRovhB6/z5Co275padDdb+VY0+D7GAIB6rlKf//V/MQxnjAg6owG78pfcG
kGi1HRtgOGmGJs/z57MF6Id4WcpTZEeOyGj9VvYLrLRe5QQ/yRRBloikSvawVwQX
tRukIC6jZkL9u7iHuN9OlqPKWSue1P3pA4gBcMoxsW7i6hbi3jOYCUqksKwPp6xx
Z2hmiyoohbV3qtFguIwgnkg6iuNEYw4f+uNLqqNI6Cuww0PtxGdANAMYOlPzy+O6
Dc7Dvm99D/DcKyhCv+ca2EgJPmYYBbGqh+eSLGBLQJigATG8ux8JL/Eq0T9LeQZu
U6i9E2WAPJnXfx7O7AZ51qp7LaUqlQOjyk6jjGMiopjJMKaoTyXF+RTPnrrAhwG0
ygbXjKCuWNwxhw1EQITC/krLSHbMsI5Z4/kG547IowO8JCezJldueyTG8xZ6LGLK
HPhmip3pesbxMQEJl5onHBRFOjStZqb9JcBLp53pl2ddtqlPU/DAENK0X3O/IqHq
BK2FphDYN55eyRE8chVxVL+d8LcllEHv6kFFsyyhWFKBNHLJxxy1tp9KTrlkrzGE
ZgWIlmYNXlpc0v+GX3nmkPuaTPQSq5hvR0mRxGJ6hzWzfJiqzFbzdFSQicNfb0bw
kbIp/LlsWpECN7miJW2WISaPPXqw97lRSMkHCMrHXaSU5xFyAeOnYoeXfgLO4LAj
69vxrotPWXTwKayLlEMfjbrHRDGs+/7WuVvlJlIDtaBTzMqq2Vndj+VZZNSgdNnI
KJe3fqnMclQjiy4TbZw16SuypyRi+APiYX4XMHHUZgHkfNkhufnutbNJw96EyjSG
dngpvqU1ld8gdjP/E9NVEuGd1YnyowozxqhTmt4WA/CETXf1kp+Jvnruf/wKvUYO
40zHwJ9JX2o9jA7sFVVrGd6n5gyRNWTL+VZzt2MlvXngm9Ehk0+vC5zYo+K64aB5
eLNcUI492mKLjFVY11Z0gUhARp+gddAV3miQoybJMxGBiSMtI6l+zv10J5hfilZg
yQjPWBMVOOsQVAaFmv8P/DujzvV4WTnbmSBsB3TtC5s/h+myWaNGtTx4bASBOoPI
wW+BB6z6QaZVBoadcvAUDdvcvwF0Sn1Na6Fkrek6GTBw6tWkftc76twOsxTRvV2A
4sS4ZrvRJy8Dd+9OoXwOC/P8l42427g9MG8CG/ajP8nLX+s3iq14iu9JnIgwr3l3
GcYnSacVY8eXo6/Q/SSLzkoGlKftBLqeK9zmuDepHMPG6Ck151JLIf0bzCWb8OY6
aptkc7r5qMuQE9nrlWX20b7nz1fIPrQCriCFPkLbzQ2gkBrNW2uqdPRrULY/L9XO
i/kg7qayIywgiRnAjKfZRZZXyGlEIiSYAWCzx1/wNqQWGRHoD6KHycs5a7E94TQY
82fhOBmtpqKFo+Jp3XdFp9IsGrGvUs36vc7nhvhANsVsIQiimN8BoVrBZLTkJRQP
9UdWEIHLXLrB+4nCw2NxjcXwA8w8BxxVO3yVGDGQD6npsYMpXvH6SWv84tsNm8w2
2FOl51+zQyks3KEWV4iVfa4F7ZaWlTBsCFM9vDz98GskpVQ4z10oRLgGrh5MVT1H
m0WnRwngSjYEa/z196ojchHqO1BeKpla1GTp7wPRoa2H5pmYFHBew302lKLRlmta
rOkhwrzVfrV7MiGPdYVHSL/7p/Uet/jacORvbES7pdDkmY6rtZ5dEOmxN2lrjfIA
rcy+PFd4sJCli3/eoMJJ+f4B+63zwkdhf07v3qR14L5wfmBcyaa8gCTCpDhjXDqR
4e0Ff2WjSFc4vfUwxkuVU0KbJ4dNCSHOMs5FrnJXhIlVI+ymfky+HB6BuiB6CihX
opM8EKYSSfEd24CWbPkEn3QQf+JvvaRVYNVbadSa0RycioNT7TizJiDroOEO+0XN
0avB4hkb5G7Wl5tlaIZjKlBZRmWQNZoc1jKcZA70b8P8GqSuMnIvnS/xrs87HQRb
R0nENAfwKfa3KIQ3Jvb81wlISKuPCmeYdaAez/aQ2KEyLOLb1TiNH2Vo2P0H+Uck
/kvIbe9YxC/D3lVquqyXPyFLgTpzmc4DkOvmjCYEVHCBWPP03c8/ZnGhyfH2+sQH
0OByFwAOy4lc9NXsH2jJxZgS1XyJAsQuk4WEWNnA+HgKpkD1WncAxQ3jIPg3JOGH
DLa6nMN1BFesuzI7FGrNBKd/rOkkl+rKc7t3Zj/CzjHPnMThxo7MCs3kqyE/H2bs
/iCZU+TH0d+baYxCdKUNVkKPI3sjLdu3+1eOsnmWGXrJUoaEcbco0kB5XunQ2qDz
1qOIJ8eXwXYw+FRVxwxQEeg5nIM/GOOVb+zQDVM7Weq4u/5CfRp1ok4TKosjxDpY
4CC4Jn4MfEgFeiO4FijdeyyYcIIgo4H9iwsNKwX7cWe2hXU4wAOCkYMKuc6Bm7Un
0XGLnWwYKViho9jtqUyF/lLWqnRK+LgAV2NhJf/PUrOelKiLCPYKynrpb4+Pyouy
BWoZM8KfeZ0FetrP1sAOLYPWW4maKciKKMWCPKjWj8xavVx2KRJuELw6mFkyN9h5
dTDc1KTJ98cLDaEqgA3dac//hQjvzjFPICDvW7zBOHPlnzTSJ0/mm5o1dJ3Tx9hN
tOu43Gh/q66MXuyluCbhXOwTc+glTXSirRfX5q2X+UANO0cAxeLRwSKZLcicrSYi
+busuSEfCimDz+gxcfMECP8+7zpPPvEGNFoR7FFO7JpgqxBsFueBm92dq2KCy/Vl
hSUz1jTi3Qty1+tbJ0tlIc9f9tgkkP8SW/SRbdb10OPZ7E+Q0VnvTiar13CSnYAK
sRNGLLIKFp4o/Ue2NAYMMbojL9ONhJrOiLkfe3AcwnA3kDODGdb/F4l/FFnrsZ8c
QRYAbIrXWlunTSmDvin0JtJVpI1okQQxnFNHBY89QM4O/j41Zyadx4susbcPVhzb
Iv1yaFo05ACwuQ8ub2aDnXwOekl7L19O3cl3dYT1dINC95rSoEQa/iDjhorgIV4U
4+dpOM3ZdjGu986HOqpUrWrX0R4KSX4Emw4P8BXlxYzs7RVwkJELU03S/Gk0SJO/
YpFAK0xW2KqOnpoIX9c175575F4SS3SR6PN08L9MIG708fYNKbFly3G13txOkePo
jFs9YhIU2nMpOj1EQlEDUfSaIKu8y388qnSGzXBQm9pAT7Gmp8oRseOxSZEcno4N
IG8jDAsuw2lZg/5snAyZqrOehls/c8Z3itgEo8tEqem4vR+ag4FtI99VTo22m0mp
0OTSF4Lol87MTv0mcsPZlQKyLLvF5KiFKfRglp8L2fi3qBH0ilDkDz2qXmr24Roc
XQpDIUidG+efFyfBnSXgQftMoNZCSLQ14gdVb726WXbm5nKJIR1ZSqtuRj6b1jHU
jzRfwveZP44sYzjqZScumjUAxMJFCYCriRXpNlr2mdyY7s9n6HoEFTD3JLwqVfz3
XO1XeC1MdwbX+hc4gK/pAAuxXpijE0MW/IrZF8UNUKZXTCpYoJEPdatV1MQXuJ6i
l2a7BQe9KZzbLobz76F7CkghRHxDmGjzRt9j/MTo15hBl/XlQeCYgbN3ERwJrVbN
2gjBtaHxrPh14WktqLEEuCmsf2nfcWhbcu4TjPXcWfZ3Yf8aPxbuhnCKi+9VIYh9
w5t/SU3flrSZm2plGXNcGctQ30t0TDDAs0m9+RyM2QcBS9dDoIGMaEKk/rLMyC0F
DIFadlPwyxs/exNXfmEzUs42nVzXiCS3VHELX7RCd4nnPH7Ib0CJx2zHKHRp9gKu
drdeCZGhMT0ANPYI4O+HJFMT/C1q1F73QMGl3cvgyDw7e5SNVAU3Hc10YSm0FgNe
uMIheCp/SBV10aBfC1ewbqM4qKl5AgB+az4vmZVu/YxHheQEQFBD1J/kWjPExgOx
PbF43izZwb+IZemIXw7yonEx8K6HV/YvXuIujxSovpgjLXw7yr9I8Efow4ZkuRYb
HZ5Wbt55e+DUXgNO+B+AANxDwVcB9NEVHYLKAImtieOrqmlDbMg8S6HXklxCkN5e
HtaoHEbGfTplU24Qmz7RBDuL64JDQexSDtRNLIjbbb4F20OeBpng3bNDdKoa6ViH
J9Q4P6i5eum9nBF2vi2ncKrt/YwxMeZ0AywjBA88FXNjS1Ya1kVbBOZp0BtE+9S5
TflW3oiqyaYOzRdu73geMD7VN2Y+jaaweqmQXW15BoUCDPMviL8WwcaESZVmoomq
L9GiRj/ukWlsimVKTTT9xgl/Z0FSqi3DtiwlldQC8ftH4nR3+qPW5wKfngoTqIOz
DbrkYI6AFDGD5HDNwuvm526WjRboWNAqg0/8osXnhSV7nFIvH/R8g637BB3TmEso
X5PpbH/TUAdB1rXB5ksXb3aJXVbCGyZsitfS+oJbEoeiDMh3FvBsSE0QX1+5wmIW
LKtt9lIgWL3UGHFDwQn6Mm3roKhHaruF9Sro81hIsh81ZFYR6/lfweNrOoxalApb
JkosFr2gV7BoEs6DwhrPZmECcb6PKiV/WPi7SQqWM2uzzHfoGy67UBtEjhcCB15I
oVraDFDtrjLc/LWmJ/aSaP0uaOMmrtn5KYpoS15C9WqMaf87JBd0cp5PZ/KYDi5L
CKjaK4N966/C8V2UnN9ld4WxQF0MtQc3XBMY3eYOiOPUrgC7HjjORD3QXmJBix61
sZOU0dQNlJb0ZwnO9h1IgRJokSKpnfMheAZpPAv/Dvupxsr48J4fosxqBZuhwwBN
hp/iz8SA3VoDYmxhhrWe7eBsy+JzBtvl8+YLZMy4MDeS9CGb4h8hND7JoCdEKtsp
XUlp7QZUKtj1OCbXRd1v+9PhuF4DlGv+8B3FETQj+fEcp3Dju91D9JrmlkhlJkbS
HYN7045/5HB4xpcLo/aocp3jGbYZ42lq0FQftLuxYDX/S78ueDO9qiqNNRCFUpRp
QQrDTd+qLkSmsGpPlezniwj4x2CzD/O+v3kYeajWI2fxzU0cNDgbThhWQhuKp4tY
AfDr6kcfWeFSFbm1sODjS/uaYSXqRJGzAfT2IuVJb3Y+j45dLHa+qSUD7y+Di4eC
Vn7vyhdbVhUxCq3+LFCZHCvsFUQKJwc5+MY6CN/DRT9c+HSxBTZf//ApELIf1ISN
+g6thlvriOT6yVxHQuOzwKVUZXfp1LwOHKJW4ybh5meaERVyvlVMlwZ0/Pt7gYt+
8HNNui8GPOXl5HkC3xx4j/P5SM/lCpwZXi9dWFVMEZLwXi3352h3NCm0wDQ+5+z5
yV2bMRJY20EZnfcmKJvOu9ETeREnxfShg+vXXL3MufqcqsRUDNU82RSiLIgQChR1
QGpXIWvUwvjcp9JdFLgpzjqA46wy287jOHFfPFhKBU8dQCEWdhlJA8FFZUCJehAG
+janDKNfBDITjWc273+aEpXV99WKM77y6qSKNXJvReesf21weuN9Y/paXpyjoQKN
v9Ow/Lt6P4wWWPJ2/hmhob5iwBrOVKWhr2eJXbpBj048dEKoacLSEXACyrTiQovp
Id6kjwAak+XmLZYHERmZ05P08hQSt2l7k3Pn6wugEoDzFaVAniEJlWU1ALrE6EHy
Dj3R6ht58c1bsSxZ+SSzik7pgY2Jo1vmLuQ1Jcpt/Om4gE60hIHijBspAXZbAjvh
1VBT1P43IZxlLr0ijVZqEdIBgEPBbUvHObgeDHdEZUkCV6gzxPxq+Cifx+KuRpRb
IQ8Qp4YmCFe+tZIx0b/G/pv8tlt9dIAdlcVuVJrAVB5AfISperSd+hR/2sT9w63X
ytdrg3fL/OSgCqzqdV00wajceh+uri1EfQtVY4HJUolXAfpcvUoyK4J+ikafP0lI
BUZ1nU1vwhKgEDJgTRGPqT7oaZRGskPA+8F3RIVeJLkRnkCxqPphQyfAtmrywrQK
ItevflUIPAvfkgnNGt6b3zgotzyaVQat+b2ye1l2Fs6bzPynMI3VGnWQ6/LQy7Qn
I4UHI5G2nIz8s13G/r2a86pk8OODbKUsYrnsRzZ8FKy/n/JCvRSbHVEaDyzNhUe2
ttebVcd/m3DTpRdUlvbkemfseAIck/0ZPkdJeQBguAtpCRzGkfz00Kf2D9WnMY0K
rvPW+235LIsyjz6oFlSxUtUv6GmTq7Yn4vvkXll1Nqt4gj1o8//kKXNAXwIBROLj
Hi0tFQmzbq3HBmotXrwXXhgIfsjper3Dz0H7gl2i25Ag64bxhoNnPO1+Ieh0whDM
AdOzvbOKxvrW+XpYHxv/2+dCqFNn/cA/L+1GRn72o6mmcK64/95uOilmxg+gQnzi
uKRuF6Qg1u2xyjXwRWTiHbQsb+3iwv9BTNLzkOzlr0/bJSSm+K+eSnexsnZZ8P7V
cGYuUFioXwF4ngZqgBrkfM9cr3lc9UTq15PehVKlSZVawQx1cnxASkahO2oBrtIv
K1+YdAgT1ccd6y/vWeG08C0Er1T90gSzxDibK5QgLIDN+L7pDZkAKFnZ0z5XMdeN
A9Y+v2tI/jdZAOdkZkwEIY9vRTXD1DpDUMGDLY1uyeoJTesXHvDxM7DYiNYduwJH
F7GWNhTWJeSGg3xbKBAbtiN9N68FJk/izYHPl23yLkfKdH2bc+FM09rIOgbdx6Le
cE8CTROUVTzidKyQuuFwWbUoDJRhGB54VPo0WtIMVICxgTyQYxJZ+DlVS1f7PzRy
9JfglVPMxQSY/Y8NjgfHEfjWEhTHIVSjWux/ca8mdH37bHnjkW5jp2iVJulqpigy
W8NwdZU5RvYl0kn2F4LHNy5+vJSeeqiNEehQWX2CarBIP/Tc6k2LYPgjjsCLHz0e
gEBfiumVNT2yyRO4DFo3p6m4JQ/xS+jWKhCKW2nKagioqoIvgr12fqP6ngmIP3A9
e5r7s8N3xaw5e1rX6Sx7z6fwncLHxbtMMrwuFyfSjTFJrmXxJw2GMdxHIh9RKfot
+AIyq55gEtINTKztOU5ptmV5XO/BW1ZieAhG3SK5P1PQm94541q/NXQLIT46JO5C
i2nHw7iJVXswdaSsCt+ofjSbOVH8TBhZ6N3oeb9OXi5MOd+fB+pqwSDgJwVwXcS8
Q//8DWoGD2sk7rtxSJrv+MA2e5MycXzSMHUMrEMSubSVGAYNpOkSeYZaaky++HuP
ph+jrxc2oDFd3iqUXmzVUrX5EkwQe+TBbvg2tiZ3rQ/dNrxkN4YZd1fT2S/xU45j
uEy4RT3liS20FFX8o4iNwPkSNPct+UWCCeW27ZEBl+ugC8EB2l1kB3aSJ6PZaI2m
MfJdJHVu3vlEFUQtTKSIOir9lz2xhcoBGVfDyiktWHp2Z23zZAsPPcSfJAthjoyi
OjX72B/a7DBk/yZoJDf0cHgT2eR3MW7tCegM/bYpqzZSPqLr6xDXamqp8fmAOZ45
Aw/uA/eMnSJU4wGOmGGupaIXJKc+FsoxRCj9d0J9Nyn+1v963931aGrupl6QsE8q
2iICTw+H8xfmPEWTDSy1KZHaVPXtxTOnwoXQUdC3iMSF+r8BsNJ8r3CamnVPZxnQ
7FJT0HOZfBvGR22v1sx6gQxJ7/q3+xi1arSKZxWNbyWtH9PdCsCHvm+j2r2Jg5ih
241hoXHaiDgbZthgbThG2+SQtfrvkIPyWilP/MGl5vXlfHZw0IuRjZ1jfI49Vq6D
398G+2nKBdpvmqy4HfJJ5BVPMsKlulbKo5WX+uQ8IzMLpfpiifZ1nX3cfAcNTEqj
JaWTk41slnnCs1iri8jUbWZD1zWsCfV612Sk0+juANFvvEak/XrIi3bK8ZyNCy1g
rgnt5Ortwc38jFi0SzuLbyeERDeHnl06OXbeEaKfcRrLS5k4++ThUssaTzRTRErz
WATZeWSnrob7yAFO2FHjfh5PtyYtfMvRlXRKT/xVruiHQ5jhL3NLi6lHGOpAszmK
6Un1s/r/NRNWfkI0VdWMRAsnzHBZbF04h+4OiOubuBIDXHQxm8CKdID0yH/QQdiz
iIFahdmHFUoOLHSDM0Mh8FXqMkoE92bngXPcjgstmn+nBGzulvJ5pCnm9P8siivR
uFwPTogKqznEwBoDMOZ4D7/9EZ4K93aJKXZbpHf2hVASNGM11Jh9fXenDXalQqNx
TCbV6ggmxrUM1N4CO0cn7r3u6Cl7NNXX3ICo64pIlqkT1e82sAMXSHEyEAe6COsj
++M7heCvlzcRMoUKrpL8665JaNzCRBLnx9oX0OqGBkAGEi0JSoah/A4Nfckgd7wG
qbuks/tie3C9p+3eLSf8dcYCw7ZrZZEctuOCjabxYveZ2XIwVDBJMdv5LbjFJrWd
pKE060JC8pQluBsc7n+5RjueGEjWViUs6lDRWA+7iphIDx8WouuelhZTU6KigmMV
e7Grkr7RhHxQwgg/IaezdpS7EIkyKo5YpvoDdjvL+45HpbSt6Gini1OEpw5bDx8I
nT3GXNNqFmc96iaIs1RRLG1nSLUztSfdqtaPl/5/JE9kC3IU0ClVnx1k58Glv+TZ
Ie2P9At64OSqqz5oZWBtXlvpVwpPu46HljgpAjR8vvQBa9/F90kkN/jI/yq4bBfh
VF6iqNomWrtr9z9ZyHksMnt+3Oif0DTHJesTRotx6ONGnCTZMRjY05l2iZ6ynM3A
lrnyKKBHi++TnIxZIPWF1dM058tSuRXxHmpo1PVuDvt26ekn/gzRYLKigJC3bRT/
NWEBv6Fh0Aeg6AVnEI6oL2D4oq8QAmowxTSQPkTOl36GqDbs7G7u2VNbV9+0LYC+
dQF5zAfuHF00a9EtcgBtMf83mwjUVJdk96qoPTaZtpktq1j4nyBYeMKrMWoWdGoE
O4MViYQGfsHaLdVjA0aM5ef2QOeFgQgjvWAmyUjiz9IiPtAdq87JtUbf56XFfbAZ
f9uCluIAKwS6YuoB+7WJJ++kHIBSp6jdE83+vjBdxYiICl3di8AuWZ6nhUbqKRtC
IVvKuGmiAxiDqpE7qAH3JaMB1Xe4ka8uk8253WQ/49dz5QwFEAI6h3rl0OxT9/3A
kh4mXR6OkDMLZ8kJ9gXvnIfx363HoaKAuG/LkrDfnEFK3ds7HFqHK6ETcNI+CTQT
MA1GtJ9TSL1B1VrGGEahaml30O1Qze5vV9+h3h/H/L/okWfRPV5Q8vXnyHQdHJTu
fK3TUJPUbcT8Lo0KXj0PDRtzEmOTZIc7t6eVKXib6lW8WidlkSWOo6npEq2BsHga
wyh4dj7YvEhdRPtk3aZr9Q4iVUBICNQxpMgUGO8MzMouvhUsblbstmSAhr8NgxMa
w6z28rCKkLBOg21Y4SlME75z/HTTe4+skQ21+LIgNVlqenOoesAZw/F/2jXN781g
MvEvR11jeqTRtcbH81jPuTNVdF1q2g96qglDOFpEsQD0kumtvf9xLnqr46gtc4Rp
B1b9xz2bD4xsPmCwPeQjWfknLKA+13PZZFLEkGmYDZkptOTXlwE3lqwVbcoBklT2
NFklyuyJkPFcs/U4lRH3EVoijN3m4QOrnTqO8V1OAfSQ8kZ0Zi/JVUo/LIM0MZT3
wv88JtQfGE1qGp2afQJQWfDwtl9yfTc82drY7OzR2sKjqfsG7zt+jURvtHsODw47
vcNOGGuuf5+XHyjVcPpOS9n4ImGG6eBkKpFhiBWoVf1ggi00lRU/XbL0yq7apSjw
SC3C1OMND3koXDdFdo3yKf4v599W/Sw9vDp8ivc//8J99v7CPnhMF2Ncieq7TdO2
cf9XQMIz5r5HCMf3tYWR+4Vf2mgyiFkA9XN3NYhC+y253thdiV9tfQyVb1kC2iJK
n47j6OuPQ9HQaXKlp3VBRCPWeD78A/pdGE1ediLzQMNDxOlf3uFp4fzr0NC/nDaj
qbCz3y3DGos4qTpVN6NDmsVdu+7mIFMybqwF1K4ou6uo7k99cAfmuNAUV9Gq2hdV
IJUaViu9b/VdmnEJ/sgPmLXEJkNgfnlhLyTjbTW4R7sW/oQc2YUPhR916szIeTzL
13SeKkbKftgikCgCkX9DLBd9/t9aNlR3jgoBSn2FfYUHKmsS1AI1fwbi7LaObMdo
wgoPfx0CbD2Vh6T+fasaDbgiXGJRe31qwCzbZucOYsJvlaZaqs0KM3gbxWt8jqwt
krb4v67tKPu0VWe0/NUSd1bVRas7fL1zvD8Z5EZ7fndJ4UH+a32RS6jR7WOI3hM3
zi0+4+y/+tD7AV1qFMzHVBu9ZI4DDoD5kUK64nYHI13A+DyOCmRqn/JTNvb/xWX3
RoH1h9axDcuV+lvX9thoAygfo54Q/gRS3PGQeXSZZR/0GPmYxND0Ne3UToJz9GnN
BObB6Y7whoPWzNBXZljj0w59Hl017JLcRdOUz+deWixIawtC3iqLwtOi/iKXDY22
DJhAC2CZl++gX+ViTUvIA1TQ5SRTT2x3pj8N6wyBMTXXoDuoqlXeAcKnVktgpwsP
GUecEeJb3+N1OgXtBleZ62xBvvjg2+F9xQwjAAh2M/W3pApZnGsAOvThgq22Ss3Q
BkqHQGYL2mjSdzN46ithNz9vFCRUUfDQzA5L/m4TKcyIKn0p2D3TE9GlOjFoYizN
P1ruUdOb+B9HmNg+yVlIWSdQQX2NDy5BzoaQTeUO9lsy64Tku8QpK4nEiqOKcxbY
IVkMP3/h7/F7vjIVEexg68TPK9DDwNqO6vYZ6k4a23WboXhFUfInnWGUHxYvHoKQ
LvEFfVAPP7dCN5dlkeiGuq9qfrtLAzWUIrnzBAx8lC+nqrQzJ2Q4LlpftgAZzL5X
dwYa1l726QDK7TVmRwxigsVVYNh5Ilm/xGvLI1QDCPHh+u3d2iQWbW+3JSYlExvm
nrRnUKhKS5MhYO70HGXoUYlrbnqvMx2oi19+/PYNBnM21BKZm6zGqdcVEf5tgCC4
VOadppPzu1SIEKiQFen9qb6u5EvywLgIxarN5iTvDqOmbaMTfhPThuuupdOJTjds
aO9LGe4ZmqUn71ubwoMzlRhP++1nrX3MmBMJuaG27I/sli9aq1VUAFxxYgMfG0pk
gKxOri1nfrjxuDrlMuvEKwVtyLtChmdh9kiOxw3vdLUfJdkHxlxV5V7bCw28HKnW
qlfiAiO1MI/NVdjFZ3ku8ZnuSz1WR3nfJsTKjNYhFzAdlmanaprlIu+NYzSll7Io
w0745ujHMRc7iGJeojT9Sa+x6UJX0/0K51QHb6SFx443chpJn20+MWhnh2Y3zcTh
D61kRqLg/KQ8RoPhstiewzQcDJb200mboHwS1gml/D9Xncpgty8aPJBTV77riMFu
Vpt3AyYJJKJwYbMl9ZEjt1p65z1O/ASJ9Xy3TUU2FNmg25nperF1MlQtzPFF8FuT
e1eh6bP3RoZ/HVLAhrLa1NG+QMIt0qC3LxFgfFScHODVrY/5yaXM+al22Tr3OqVg
3fZAMjyBgC3mGv5VmXqm3CXBlMwqerSj5RK5g5fzGeh6fBykhKh0wsHGZgXeMlrM
DEj0WSp6xkYFPIvPOwrZ5qvxDtvosRyAqRvX9Fi2KfQ8UNF17ZccZUvfs5gL3zjg
2zNpnUJU1yFBCiutO+3w6hPS0Vf/GhNDRM19Vwpys35pnZPPCTSIRSV+eqxgl/45
UbFELD1Y9LUF/XjIzZNnJ/Lk/RvVhEfnAwj08oBNMcN255coOLi1LnOJh0mOIHsh
+ONhbsP4kPMSC/3A4LR1HSKM9+ZJYtlkV+AEQV3W4XjjtirPRTBH1EWn7xSqD8kv
+sMitSdLAHIx6brdNpYzfxE1OGgZbCv931UImTlG4aewhlYU8jkGatcKUYaZvm9z
PlXt0TTygTZQzfry0daaLHrAkqr6/ZpFcw6m+MESfbKSL3T39ihAXso/MjKW9oXE
R+EzTnrAE3q28c/XYn4U4wcQpgxspjwoJdXzTaE7y7/ZAmC32aOAXSrf8+8gWE6Z
/2/rjwUw5ZnCzABo6RMPBDtklm8YNtSNzMtYP7RqQ2Kqi8k6pGSSYyS1/ykhsQsg
orBQkBXa+TMmMmYOzBTSl5VlbgJVboebi2bzUtu5NDHHk+xx+RRhYBCFGMmcQc3Z
1EoMVM9pyolZLwymPGbEdRGTEbc2A8lJMwOjTc8h0nyPr6YQ2MY0cK6xe8XzwK3t
AIp5d8XqQmKcyCbjJInKCff7z61mEYGKTZxGkUD3yFPF00VSfCgz9cDdlUz7Mw5f
r5uGRPzkLFWJ9Af/DsnhSQSdj8TA4McCFSJlFF0bPwLtyTU91MVQFNMc7vk19FT8
Q68IL9CdhLRg2+LJXzr7IsIrGIkCXNzMlcfq+A78/9Z8uV0ALny0kSzHcWPUzK+Z
EOvCZa4sd2KxTip8MtGIX0idzOPmpeQ3uzzHF6/uuyMlATqjbqioA2zShajm1E58
F39NE5qiOtgB0x1v+3ITlFC4A9ZxKB/dr9JOcCDpfwFLaNfL+eMpbGBcG4f3S1Xc
SBYRUW60gaUr2oCWsOXnGIjeMPt1hkNM7n1ZjSAcGVGZOfeYCOf1hfiekc/VeUzu
JDMFsPbV+ODRU9KE9EENthOZ0nrnBgmQBzSIlV8J2Xl4rFn2HvMlorI+hnk46cK9
Qzo+LJzXaNKF9eER6Xk0FUGHTXL+sVcNL5zYawLAfV+vXAwti6A/uoNLidNoaCV7
ghq622YyJgYa5oScxzAxyVSCGqbJmlGPdHpVNPqfRwOIeeD6+wdpLl+PBYbfCS13
wdymHJYK79x2xJdNQQUqikkSmSuL2ZjMeF7570HLKkf++v4VK5nwYeC9u6Ktpmzs
+ZQhvhXOSuO8imhiZ9D27GIo1/WNF/w3uHXUgXxzOo5XgjNx0qeeezj807kTZiTO
UitvyipIIz1xw2FpVUW9ziKkkwTWCV0CHHoTZJ5TJC/WAv2Qr/MW61nN+FY7OVLa
i0XRAXzbxj1sXAK5BKXLCPdwnzPYM9Vm4RqPMtwy0EGAalMGZAZYjQGqgtY+p+lb
11zcVDL/bg8rNkpDLNKZ/uo/bIzbexW2H1uVAqAzJHHWmxThn3VUzg7VCd0qjNMB
x8FLx+YW5bo65sATUmnFbp4GKf9MCgt8Ucq4rs4O0ItFDclnpX/n9iGsR/5R1S1d
f27h45ALDRXKiZAObAMjG8V5tNbRQdwHp46Rms3pdHddjGBHAaQwu+d0uZvNG7Qn
0tx7HaTrUWOP52GN82XQFNKwr+O9+rgrVEodHYj+giZ//hcwptMoefqY7snCO0Em
J/PtOFTi5Csg8s60LLHoFseeE+sCRMWxu3c4hrbDP3usqiUTyG0ntwpXVccdLeDU
fY8LnvgAPZwDlB1Ic6oNUzBEepbpjik3xvT4twY93aaNBQ3z1xJJpLvf/iaKBGM0
1IAQlK8tNDQxtlTkaj1O74VLOLC5UA5TvYT4C0ktMnVuybVwpfkCTaF9Qkiv8YPL
fhLZJSelJhzFDElpjSWfgYVwVQCDay8H4xnf2Qa1ZXfWOG+ptO/LnQ2DUe6pGnXO
`protect end_protected
