-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
iLOKm/4QGjp9qu8gRWso9jKNJjJ5x2H9XjK20JQ3eDpJYw+0eEnjK6thMdnR4zsn
uvn6xgAyva/LQ8P87WdqP38/8k2009ikoh1JXoqAwDPAD1bgAZsqF1F1iCZcqWZ8
la+S6o0EdvFm56pINeK8fx5IS/kDZQl5yygKrHXWQO4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6096)
`protect data_block
MWwJN/IbOZyAJyAEqyGIiewhWmfjlMOnGW9BiEDlNVoLgVLNT6GYG1RgJcIKhb56
zQrHE8ky3VOoRj8XBJ2ZSq7LL1T7ugDHJkpjGaeqd3joCLZehtGHorTVykMKW+7G
bk4H1I16+/K4iV7PmsRhbNLCcROfmjpqWTNrs3ojVuA3Vx3lQ75Zyi6a7R5Cu/Tr
/LLxwL9lO4+2Pm1ozfr+zZECIN8FRkdNZES6a+3e5MdB7SKNzGRfnAUWAxFYXVcv
Mjm0nf0pw+Io9XcB9JyGCYW1Z1li//avOBAdj+KCsKAM5XpjrUijxWp5Ecxzg3rz
t9p/JmMYdGDEGHo/XjD9l3QIBNdtwoYJrXvr+OKDydtEN/Cky/P7GgrxswiITwlN
XypiAMBysT9qX3UX4pek3vFT1yCkizsZq9Z+W6YfYG9oLnfU12GnQP9ilhCPWHV/
ndAGJ4vy2mozbONj+wnz5fbR8aXGcgbRV5eVyUA2cGIcYt2oiJ7z+9BHisCptZzB
VhBRtTn5V189eampNbWNa+fTN2gxeP3ejE1aQtkIst/9mVAeajJfWrs3tzxEE/k0
fEcxxGu/tLXOlvOaI+ylqP5oGvQIbgbah1UEHfQ6RDv5ZtaZn9q7cbvIOH/iSZel
1dmjCJixz7tVxCp4XM0nPPcEmNNyy3LLF4ZA8b9a57z2A/y5kc7ZVxU66SwQm52U
z7Mjn/9WOP77FSpopSrNVu2jAkNMmTG81bS4WBez9GORMmqjjnQYFGITn5lP5IMy
VzTu0qefiphs0i+xPm8mB89/HmpbFzx1jec6NKhJ2grhuI5uCbcDRMrs2mlcX2Du
R0nWJli1DJMKLG7qwBClPROodvYYkvTWwgeAf9bMtn03sgJDlCZ9Wy/eoCD/wDr8
0KplGELWvpaPUIykX3lVtCXJ+9RKtA5QRJEbRNG98WcV02ZMsx51tO30A3pSxsLH
DyUay/EPWAnabAQxvWqhnqt7LCe8aTMwwNEiujF9LZZZql9M30bqF5YaPrrW9PoU
P95gkmu+a2DUu+tSBDN5nmWna5stXNXCwbamtauFmXw5FgoLHgqHx6r04IlMWWae
H8WNVeOkTslpENVStTXcK29UMLuhEBIJJzNTCzdHWAQxm0TOxVRj1Eg8+GxA6XXI
mNaoWYq2g7j/peG/YGAiQldC2v6Rbojtqu01/5p6Ges5cWy6U9Yx2F0E0cVhXIIF
TyMeUfDLpVsHmw6M/pbEAa+AyO+1MD/3oDxFHU8tRa8Y8ZazxA8GwfPvDMAJJK0x
CmyekicAV521v7K5yQED09tj6iFuE+JqBHJVdCOaGUrj5JE0fqEezR2q4njU/MWu
wDJ6dIgkhFuk50Nh+sz2tGFP+6gXzXA3QABPYXc/Yu6k0Kul5UfSfjaD9W48NKox
tvwu2D6JQ0fiyWJA2mThu4r1HZ+3+f6B6ylPhSsC6ANgsS5ds2jox/BV12u6fv18
miBe5dlUelNM3uHisC5C+1taZsH+103buhs6S9hyZ/qFmcMo2ls92YBR90ZY0weA
SqLbX1H13a3Vkx3bPBrou95W9iPnY5I7MSP6oHNiGlIumPKoLgOJjAmRTDntuIsv
CGOe/D4QaMNKWlCLtVGnK1nFZFXrYhTxtS+yn/MODQ1IiWp3Ld8dJt7dwM2GgFT+
2Nw5jz8XTdMejEm2jo3Rj1+AmSB1R1goaBRDzJMw/jqg51INNzTU5cldKXrxawlt
v+eg76mfuUTLYFmatzbix+4v9ok1iw0NYpKgsOq+dt8956mK3zEJT5bAlT2YxlDQ
mfL73J1AoYw1hdY0OqV1U7SyhaQKnV7DIuPhrCftGsjL3uvm42p764OU1ReCk1qs
LmbNkPiDxn56pg6w/tqCjYTaNVah7Sd74+rkysun723YnJNlfZfdGPwqRoORvKrE
PGw7RjZ7jfg1DrTlRGDmqOCj4V8aWCC7kMkMXNqQpZaV4G1TngxsTBRBVJJCl4ek
qFLjefDOpwxeXFeyWgPu21Wh4dFpnOWogaOkigjHvO4VIfMDaLeFBmHpPCRllio1
fAYGfV4v3ok767xCvsPx+OsQBg87/2GxuoD9X1PQCH3Ot6WzpitZb2wYWNU4pzli
YyA+5uoBGd8k4AzVd4R/vToyMbvu68Uj/zCksbCRVNeeqm0kNDf9RTIDa9+36vcS
nZRZJUyQPDd9Ob+vUhiBQVcaS0CX7rrh86FehFtPopOUNTvHcdVyZmtq9yO2Wphs
ebV7Ih2g2dW9TcBaGeY6HDOY09m1SWq7KOY3gqaO4dNLcEofgV6HW27zYwzNF4Y5
2BzJvMoLSJBMuyH8jM+UM1eqFWk7rQd3832jFiXD1QQJDxRPh2ktI/JNx+M27KXo
Qcg1PGjvRQLVKUXRcdkr5DJlhbUxKKLYDTsf+xXbzqbR0w1rsPR2KOn/x5vOHXfS
A73QY1I/xGKCwhYkCr8k8TsfytRLtyKLExVIS7tz2FhqWWeeoGFpZueKmhBKfcQL
eKMmRLWKesmYUiiWr1AYE4OATCRZfIJLCpyneNuCLgF/uRUJOg444NmC5XTVrgq9
mp8zUEMFDCKZflOzGt/TM1xeOD6cO8J/ILxNYn0J8VzQU8ChLB5IJgqOMJ4teoBP
+pUQyNxL13shhtNBZqGvsFGK1S8N1/Rwe/mnu3f5wIRd8rm40iZX8LKawT/Bkyo6
zwfPYYMYn4CrhhwZ6Bp8zkNSOaeMLRJL+3SFEM5x4YXT1GSjwwSs0kQmlPzGA7X8
hcZmWT6hO1s3LwGB7QeHS0qF+LiYfMvhJcQperNWCASODB1uYkx1mJc5LZ0tseG7
jCdwOggcguE6bxonSRcFqOrGNHUzgvG0MfxdB+EO9PZuVPERnfN6/GjypyRvQdbi
bw2U/3IlSZQkNAjbT5r0waUPhbQwERuqBlcyj0HW1/PwzJtWMYb2uP1pDhBPIuVI
reWywcARo4Xdj0r2e8u2AAvs+YMXrLx/KWhQQwwy0gwMy1lP/aMCtK5kWJbCsFfe
FfHhnFq/KNS2serammSasRfoK2ivS77FsjZ2IPyX2ddgh16i4Nl4E1otwL++pjgZ
/3yQaQBVZ1bg7sgblXBK4CxovaLTklMSjKMnf9xXk5SlTqWLTMNRIpvrdbjOaBvS
ZcnrmpR4qrPQj0KvPgRGNGc1X0S++u1DeGEq5U/Zh1iQU0f8LFkTRCJ68HGsBWhX
kAjdvMz7VcZ4qBEU/QCjdNhh4xRA/w3gJWLv12nV3c4May9nzxfh8V+9htwN39OH
/k8TJ4woAP/GBcVCzrC7mpLarxhodG+HA6sMIV7m7ein9QvWX0uv2xWGxAheIBpz
xs7wXvZhkoRYsSviiEcGf8aYxFm/+GVr+Bv9Tyy/qr0mTOmQSFvYFDOafRdPXKZq
Gi/DgmNYDhZCLnayxpFwz/qev+6/ITFAXMOLr9h/tjLo+ay8eUYtNmCTrSouU5Jg
vcplkF05WGzAHaChRU7mZ6oXQ8+MHl/piZkAC/9ZeNvjTml4tG6ooAZXUiUh1zWu
A9YUErF8JFNbDjpIJeZTJK6IHKV59ioNeCNxCU1biC0CCuOhsbmFVv0pR1r2jes6
I5pr5aXT3NtIwNryn52Rr9/gj7hgeNi3KK/MvX97KWg4jyLfy7neG1KBGAr8RBpp
CHpjyipwiDDuFXiuHKSNbj+ArJp7VfIYEIz6HTsiYYQXn/aAMX0gXXPR8ESDDIjA
/1kbb1n0R860gwbtU2zIzRT0ognxNcTzBUfnrk+YsumIwZfFn1eaPKNSrEJmuCeD
+rV5TFvh42FAjvzxnPogrTcK5nNWVJcRmxvliE1scDwe5a04f0vyP75ye+o+zQzv
+e00LWEHgta3v6GVzdiL3hw2FOVAzPK+5ATCD6vMsEh0uxgCtZ2QWkXEXRYxwMUk
0HPEDEONeHG77AvZiPlWJxJqspmauUG6HrRRetb70M28zWoSfm99nYvoX8yt6+vl
9r0HE6vAgbFmRAbxeCD48lRqZZDxxS1omR0StEylSlE0Qo0Ewpw8hiqQEweswLd2
mZZoYwTr/fSSG8BQY3mKc5ukfb+Thl59m4g5l4vUw1VCYMy3EEMpur6Spj3cMl96
F3h67FumzKG3J73xb9ID3AGBAyUue8bgUhi1fxK873FEHptOUaKNdrDHY6ioiUJp
bZSE4pqNHmlyOxVUbeVqYGMMxWVOHqTbnbZ5hv97gfYt5PD1HdNDBl5mZwreqJdV
b4UpV4pnBdX/kP8mGrxlrxi//sztUSUxOTpSFC1pw1Tk0lN/7zuANDhePXoHiu1k
M8BNNEQUnQ+nfjKMu9xqprbeMkhOKwjR7/3S99q+re0xQWwgqQWNQ8zVCAKcNbL7
3woTJeCTvDBX8viWmXGaWYD5CSljCUdobZNMCu/yMrxWmD32z4YGejC/yITRwnxx
Wj+BFkAHnqOt0uUDFWIwpA45gq9V9YrsPuBF8p4+jPAEhrx+begKHD2XJ3q/UyoV
2KB/qcbA4szbth/iwUxD0l+EnZgL+FvgwkmLvJkmfPGsnrx2NNRD7e6v5X2IcE4e
x2LEYjfuuMucn0BFE9++96+q1o3ahWndtQXhwQ5e0JKkM6tQYNCRYaI7RSWn+W5T
z1ewYdPp58f6m0kp2Iq72lqtzkNF6zylqDTlTG5/sHFYTqm5OdlKZjhTrYNn2Td8
k+Zc0xfMruB9fiS3LG61B1vr0hwtSXWsryx+pX3azlCL/GaTkXXUjHKDWWQyuR//
yGab4geEp3v/01FhIiqX3nFziI1Ech+oDqOFDwgzTdjlnGzD43OdY2MFVHzWAh+H
ZtYZXaNRwN8UwatgX0tBU8vB8ygHHAPxsGMnbDGvUhFLzu5iDxzbqwNV42Cp6p0o
EqaOxdGLV1Lc64ZJk3B9ty7PNl0JDYz/T+MmaOlcsPlf/bJ7hTGMAf5A6WULszRc
c3Naqbm2hGvgd0x2DLn3Oi8DiVT5b19Id3YurAk7jda8xazOfLRsz86AUSpA3GQy
EC28gpHDxxsGcS7t/M9gyB5KEZbKD4FNL6LWHPlArp1DG5bAcYGOFaaMZaNyyvhb
LNln5P1bKFmF3mKrIZrVQu9g2BB+S2slShnmjijqyvn/DMDoS+2+nwoFyGVc2Rr8
pHTPKIW1G7Wi7AuS8+0BHi4zyGvVCnGYC91UJZlbxATIiE6HcBum08Ul4LLxFkT3
KfyJdK6v+/xLFeF/Td4YXeW+8h8iBuc+y+GDzNVIRu9jzFoqO+2Sitl2BdP8rBmx
dGnE+dCymgn8JFEuLF00nwMSSo7/40cRVY5NlBEDCegJBdPCw8rIi7Y6Qqfu5tkr
pZs/NvTLx2qG4I/Dwlp3S8A8Bk1iUDE2mXennR9las/fMvFN3C+EEaWBUVDRI40Y
DNfuFFILZ6ILPuYi8tOwY3qcoWE+oxV9/cwOxa1mg1XTgdRDgSEzM8ToFBLrylNg
l7Ni4MSven2q3NmrrYwpfpSCM0FXds3gH9kaAPWCu50+HKJPCniikXWePWa3whwo
IR3ZjyQI7zGB+vSuhDm2ycCRsjd9pgx54Z0MvSaW6ANQ4G0yDGHVXUWJ0S7rx1p9
SqgkIqikGGg6KkVt9Yt26Rs0n2k97OxQrg0Z93Za00hwU8eP/J9Q3XjuoyaujKQr
41BO88cUZkZH8Q9LaCmGED+xR1OUCFgG2a5ad6HGpaRbi0O6h6PRwqCA5/BiUPEq
w2ZRTajjjbGDqwIhVCnP3+fHkTD+54u4nqDUBckzdpnse5dZgIc5QwGPsd3Y/NMf
mc9TW2uoZaOjeEKUNgba0gy+jeK/db9a2PDjiqn30Fxn3JI+kpGOAoyLwUhdlxpU
eVABR11ke8lXtx4Iyb3XveHzoTvWT9ngD5QiyCcTiWnjUWsk7T0BA42AZl+4lICT
zBwjDoRKPXFKEy3nkBycJPpigQ6Y2sG5sUJR9YH3G0q0E+lU0Ocuwt48zSq8QBmm
J9lmbuNoi1AfpacLdCA3Iu1vcommnIB6vkqkAmkfaqHqaDV15LdvxMDBVbM2iS2g
lEMnxRJ0IdlOoNImcmDt4TeUG6orvUxGAVl4jwv5EB/7Mm6rPU8zzNLsk2vTiWK5
A4XvAv8b21iza6Su2MTkFLzx1TyycZp61HtckjVQZqMoVl2OdK9OWzG6KTQjK+n/
3I6lItmvyDD0O2JhP+5UjYQrjWWhQH6KmJGarVh/DytI4It5v1m6ts3rv60LOTXq
CeNbp1gy6u612u71mT5XM0NkcwVb7hX/ZaYQAXdCT8v7vvZFsVe2SUvcW9jjby4+
z7M6WI3XpCeGWa2G7579qxqwGoeMIFIEehBDuhAA5HDiBr7KTHXZ26Pq9ezW4/F5
bZR/5Ohk0VwnpqJsw8BGfSfEyPEQ07RFJxbZ676MZB9lqkdn/GwdDiWQUFKY88cN
6dSEqXvQPuQUCCpvz6vqCsFtKIAyJZJ//NVERgXh2wPT7M1Eo8NHSQK78K1nt5iJ
S5d3S3z3NXjJimQU6WEr9/RUWQhoIOF3COJkWiiq7V3nadaozUimbCx5acMrkTkF
sgn+IHRZtNLykgAo+y05zCrorcLFpCh/n6pVOFXJMMU76HTqBfv0XgUc1u34crNc
A5fU0WMH5pH8op46NEhR63gfzF1OuNRwwBT4zQnOT5jZZkrfmfD7WS3yfhOvApKw
V9kHciE7TSaglN41GAXb1D0hjEWiLCd9J/C3Io75CieFvm3vHnqzoznHT9nrlZtX
vxLBLgJtNZAaAJaf9zPN318gLUJiqF8UazAKj8JbE8YW0Uhjp7FZ0gdxoQV56mkV
0ojr+BNxkGdN1MAXAoNmpyvRi1/pjA5YSvtK6qGF+FhievA6G9ccedyna4d+COn5
vSB0ECRd7gO45eLsG7kc2Y0yscOzdwp4pJB0IzrCALbKXzJwQPEAPFLMfjNG+jiN
BxoTicWv6BtBJ39bKvvFXpUP/zqZsUyEMbdP1fXCikd/Zmz5ghcmOf8OUdpFbIku
o/Rtq9HLe1UDTt9jAxhgQll5ux/dysAjMUMHe4aluGy+yn37G96JwFu+grqhjsKi
Kv48iSsBV0j0mMdkICPDwADtGvXfG4YAs4DVZhpEo0z1VU2mkn5hLNhcPsTGH58E
l31j8LlWOXtSD5MJ8SnsxYHl9w14EeOFCIuuUfttT7noOqtb7J5ZTv8A65/IksOf
B92b01Ioh2EfdvS1MlyxwK4ASV/niM3UEyO6EFhj9fLlM8efZyshur4FjoWM+KN+
kT/H9fW4KQ4LX1NTKiFxwgORWT0UN/B2kI0hd1EjBvW99/n4Is+0IcsaRquifD72
9WmdfdcClClK3Ov6vdWDW7E88yUfGLWMGz9ubKpHKPa/dHaCgm7W7tCBqjLmZm3t
1SrMsic5gCClg1SgNK1i7SnXpy8loDwQvyCW0V2HBx7JoMWILNV+hzw8SI1iaZhh
hN8S9EzFFBY+W64n7sOisn4DUohFyULq185gJiIA6HydEoeXGC3SwABAlGg/OfwO
zNJyv7SkxLTZDfMv6xEDUR3jACvQB4CB2Y0z+QJk4ncWu26JdjAFAgBhPDu5PC+a
CNFvuRtLyx0NcTCM7SBU4p8/IsnC3GP3nHQcK1V9Myi+BWaBNaYJuaNZQBGr1K3F
HSP1jBXvOpLn7EO+lEEIiee11nfiuOQ/95bHnxd4kllcCPz6u0pab82R9Sukxw10
dAzN2PvK8n3Kw1jG6auivhWmz3IHEIQvoRgsk/z4ZzLtdtHOdgweJEY12/5rzxC/
t4T+wrBGvXAPr5w31QxbCWMbFV82CHZo2fe/qBtcdtzq81Lhi9QD1i4W4iE/WgUr
mLp63FbWqSYn3pNPjXifiufBhLXr8B4qIbG29JlggkSbE+Iq4x0tkhIIPXcHR0Ld
5Gd8I0KtMGlD5TOzNhvSksmJhj6v2YMGLFFoaAYxm1SWbNmai391i/O7IbdLb3fD
T4zDeaG/UuglBTIt/KK8FK65ZTpe2jho6XjJOkuDEYDHVSy867hcbIYi8qS/6GZe
p0ql0lYcHoOIH6Y0SmOBo/ZIZUkwjpLkVkLKNBSyezoPCZW0qt93DIt3iTix7Vua
JRE44EZv2EczE7LksPkA3RPqkKFcvH4rAUXA5vlHbjkkT985RlWkEMeYtHkak9dj
`protect end_protected
