-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
iEbdIsFy3lsBtkxI+DVR33oWHlzjXJLQexc0CSyA+6Rt7OWz+nlNd5ZAgYNHWgmw
ymsfVD1MWS8hg/axq801ZDviJ+RJhmIpB4WocdySo9NO8G/2/366oqnUJRiDb15N
sKUajQz8zFPpZXpSeRJiWxz5wyikBWuJjf2I0LC1DgNy1tSi8vbZag==
--pragma protect end_key_block
--pragma protect digest_block
RuL5OKG0LH45RLy74RzG8PUAAOQ=
--pragma protect end_digest_block
--pragma protect data_block
JJjh2ex5scGY1wlm2xVQ9pdCC+jOxWFZkGWYY0JedKYDnB35LRDQXCaPIxKqof5U
48HcnqPVY1nmpq8CJ4FQT2wSReJOoxuQvaUgzV4uSa3T0hbiCrIQ2r2ATdjmFUvh
7q2ycPRkotfgAbOyNoIWHuFI2RTecKiOakr6m4HCWbp86gcLMvVAfOMbo/XmjBiK
HYFEM0imrcXzYRV4Rd5z2KFLDqNE6Bc8xG4xUBt2flXvGKFH0FFOW9pEoEwSPbRY
hkMw11U28YvcyY+OSrtaqkoMyVrbm88GaZ9Xu5mvVCoUW5NxDJjLJNCJDkywlTIr
yvQk3VSxVER/xBcAma/Uyca3+qpJpRTLjYJMcmRAWVquP7LECrmktRqgPRRr9fkb
ubDzzamqy1A7Brci2zigmtNRRCo5SJENU5p631CBOsxwxHzoopWpEiIMaXY61kQR
WaDU1AI9pETON5eHetYH5QiyGGwB3zUy8hNMtnNOHfuN2zrEAgP1tS2c/LX9ngYC
hV8tfsiMKwnmYUAzXTS/Ksu0Fo1tMjtv6yjOIA/3U7yXad6MC7JIwLrlA4n/QSB7
WZpa/maEB/Gea0TJIcwkMyRy3MuSlizMcjLUMz64KwGp7PGwUcJ8562YpHZBIV3/
e3Ql3x29H8uveW0Uu8pbIivwhpR6MsXSzcbOADrkoC6irG1GjyBkrnI00foo23Ix
rl2wo/zllNebHk0wcIIZEdXLlcX9DcdNzFX7hG7Hc0Nfd1ha6rwtTjxpmXKm1mIb
VJNnNs9XndE2jBZow2Sf7OppmSyzsKBMGfktX10OzvyJLTEh8IT1jCjHMVuSFFy4
Sq31ISHsymFtHuzmqxOpptQXhdG/1EiSF+6Jdhf2ogqXU9QjuX4cGB2zBS0msGjC
f10OKgDNvqRY8lYKo4ogcKGY+CJKBI7KQxN2QTMKWY7f53Mu6IET80as6y/JfQ+e
4pb5xmpaqbLG549KtLw0tnXGGmv6BJs/qjkcmNdkhtxxoTGcS9PXZYCTR59uYIA9
ak6MiD6Do0agf5wTD6S6yE4G3eaEhaUXCPWuqL1WdeSmf5uXR0IxlgVjE7sVS9Vb
5mM2GpK10AKdA/uI0MObaaZto2a5KaiMFR+rq6MAOmFk4jS7jj9kVxT+BLcG2skm
JDbyBCBwW7NWr6Sx61tzVBouydI21u4U5sNGEvS4reVhQ8mu+e2+ttaCBnZdwniO
jhRs63gwRkvWpf+msGgE/SZ29YGj4M3iUFADpiQBUja7u68p0w0L9RTHxT2joy3x
XGrOHKPsamKbyNSx0Vrb84k3yn1/YvzXSNM0MfdMOv+B+MZDnZfMTSLSl0rGBD6O
4iTdBm3U23UMro9D/ARiphcm9WnEAugxWhGGrh+XpPz6iW19OxSqPAoD+u48Kd6L
vhQnUE9TDESG6ZhKCXxz2wjPIMVdQKLnBNEdFYGcBJTsVwJqJeBbfi19c2DH0ksl
fMyaJPN5gh4rq1+Qz+BmT8xa1hMDO3FZ0YTDnZVGu3BuXGerClI4dUTS599GyyrV
ybA5/pPAwmq+cEqqjOAtLC6ZzUgRgrfsBGpz2QCAwvuA5IUwgYsOARNzfTfgAnNR
5MqDUukdFKWMYkzgCc3ZragWQQjz993G0IfAkkVE15c9nao8IWm0Ex+PBXUPjNZh
RN9KivAEI4ZieeMHoWp7ejmQastJFRAfWQCNBmnSJiMTLlMqa4bR0L8bZ9A8k+mQ
vHj0DsVYzn4E61Wobi50jpINl9JgIsWXLW7pAs6lNRLtWv6T0hA/ggWRtrliUznz
I/owph8rC5ANKx2RPlQckhkSjHhhyxzeSMjzdDzEEhy8y+3L31BwQZCr6B22LhpR
Mfxu264ZGH/pdpH5xH4zaNHm7QTtbbg78yv5/WjCGleRIuONXMHuKi5lfMi0XOuk
WFDk7AezHPJ0abYgg0KAoliZqbdvC2bta7LyVqB8G5KfEhW9YdntuOid7S1ijUbd
hQxOVZhfR2oo25OD59uKhB8YT6VA1MekTRsmQWwaorXQgS/urYF2lQJsVQhvgr7S
PfIIkPTC2M4Sw0saE3wTHUqeB3zS89hWybchWti9vHPBOqOgYr0U9MPsCYoBWncr
hNCw5ljZzEUipk2eqokgJOP/QxkgnvuJdvQ6sR2JdMEwkl1CQzcRUgXZbyL8lu7H
+zYXh5mlmxmk7qPWxJlsfH9J05tjSlhH79LVb90ZNdr4yGwKQzhoOP81UsoPdKMl
UfbKwlTfw0SuheD4CeJbnPLJEpOmPdrZLQCF6wLtiY/CEKwjNyvt3IC7C8KlrekH
Q8yqH228HlP55GfXZFtMnTGrHKjbiA3zRMn/jMgB1ydMl9+0fplsGOYXpCcl7kEX
OZeLnagV3B5e6UYieO7cTFZ1qr0q/knASOzFkhKRMI2G6SMHB74Ti7ydQuKtv3nM
yizOk1zCLmMOllad84ZV17DM0BXouNNN5vmb/amnUlkxIO94pqYHEXWk1VhEtBJ2
z4SeIZsmKv8LfE6bAEGn+avL4GO08SYlMDeEzIA/co3zq5/gf+vNJg5g18NGoDal
R5Y/ppeWPpS4VFEY/gkDnQd65geQcBr7Gz0KiD5cDf1upnYdqgnVnEEuX7BJdp3/
beHqDvcaQhtB/C1CoOyXk2CX0l2/z5QqXtVzCjtFnYmUG9LYhr8IipktrD6GMDhW
cnhMnpHRRdO9vwL0cdkbIqkLs0av6nr42lwNJBT6dUPba7rYarHniklxFArm6EZv
qEcYLO6CXkOtvLe9CFkVs/N/vwXBz/ulpS8cZ8dO20fYW4IA40CKnIy9/SoDi+94
AIVZkvlq48OKgo5VBLd6oYRlMfauIOJ4CLVG3+DaCplFzy/lDnxyhyOVemZ1lkL4
X00ran4eylyMzA8jcMvDF4fGTz72THbax+mab2FCJxDCN1Rab3+0bUZoLBlPw6lX
fbWfbRjl8Rme+FR2EceHMfQIN//a61nHhAXDEPh/nRna6TYCbSQZswGdTHA9IyxC
K4Ej/CBsHkMZrQzOq2eTjSXzY5j+FcaZpTHU1D+HZC6JMKCPJ4PgFmBinF9iYT+b
A0D7raVnrorRXBPWQH8ua1iaMc8fXwDdxNymEwDF9tFkCRmyiViPXjYOozKa+Uj8
8Go59nnvl6qRKYQHj+H3FRzuz8hSSYNmk23WHLbCsNyMeY2iXI0s+68tLZ9VILBJ
TLFG1o53N30Rj/5cnjWTZrMhzVapi0Y5RPVK4b1Ro8uZaDL0CPhuv0lRSy6CUoU7
aU6vqwPjtt3RvISeQsrUL0dD1UMdk1kn+AJZ4uagJrBKT1w+gInn2dG1ISeb1F6o
H5eHwaHzI5HEfJ6h+jUm6CqStlQ0bRPf8BnxAs0YgjEnIZqEA05V6zVqvLO4ni+q
EjwqCNgR0IpoiOp8VfZFgY+cvpd7PQQDbiQBc52UClXWzv1Wg1LtId0jHhN2LnZ/
DHs5mOd9eW0F/PxLROPcrap430oWlgNOOdNVv6m1qSqNkEyvcw1hebIvvuEfDe2l
dcb7EGpyEzfCfiVkgIUzu+eKqvGiUPwngWr0inqbQxTcb0C3BjbErxYygqcORhgR
IkAjg3d4IArENumxBRwzCZjKx9AKb2fqg0COsmonrb5SP15B+rPcnK7bgfh8Epz1
vu5wDFpQrWiObCgzNZ57O93v0BEZ0s+3Y5lDIGyJo09k2ogQFcEWe39vgr80bJ+W
naZG1WM/2A0voP0YQ0pLmn/LcOgy98ESiGc8g+AEXssj69clpVan7tLGLteEYYPA
eevfpcWz+Z6g/Yuz/N8rL2MPmgUD5QDLR/cIErza+i4hdz44wvcqO/o90gjmMku/
WO2mcMpY4Q1Q1xXQu+Ttf3hUFg4DM9ghlvIazmsG711mYeizu7DmlGz87nvK/9PC
pBiLX3x+qe/6rRWMrmNqiUL6xCIeIRt3Y4zk6FVmAlXos2ZZexznJ9L/1M5NfMa5
Jx99svwW761wezKPRkcJ9qqekD4jZMcXojufViAVPeWAN+g3SCCdW85FY/se6E3U
iA+bRkGLHPDgtele6qIJgAx+MTbZivzs3oeyRHCrTzEyh3+rM7belHR3X6IRCv4r
h/sC2pogg3bbR+WABC7ZGVlgHiKwPmbMZ0c4QoWc6XxJLB1WG2c1YwupAnFULUrA
vJf8YvM6A/cbZjy4qp5e4M/ZwW3JLfYku5W9/4nckqLRu9te7dQ0LMkFtE0TyoQa
mmc+lH269C0htelJC0A8I1fwx9u8pQ7P5qLo6BpiKow+GzrlXXZBXo5HrkOpYid8
HqcZPU8RpzDjFRDRW1Fh4gWCbM53/MXjP5F2EulNTucpMuRsAIWN24upuCQXeRwg
osqNPlOn67SdLqHsu8QERAmLgIoTnZjGdrWWUQf9KumZXMgDrS68MAd1fWWK1fFN
rKNPbIeutWhgVd16w7BBrtH0PnJg6JR7Lg+j9hHUufOf71jAzee5AuAtL139zfCz
ioABunubv3/AZ2TkYvL4WKOUPBO7P59kwePKQYlYnDnqlcaYi7y4195VnYDXwELL
mm7RW0IT59/Cws+q1TVn5zho/+O7a2UwKRHi3b9ZDS/EYpjjbQU7byONXTbSfE7c
13jsXZY2EvWf9RR4a+AYBlnosrMlw/1lOIT3G87zVnKeyTlErkxa7tfjAlldtGIr
kT9zuLrWMYgM+NOnTaW/wdb4z4pRqYl5V/buHd0RGqQH9NwcujRzkcyqSOSPom70
Z69dBujONwlSYZEUMej8XqF9WrgG0LkplyjQHNDREeBLzNXGrzk+uT76tG7yitgN
1OfnZliqYcMPvc3EmMcLQNaoWyqB39M65MbUysxSN2prFBs/wbuH7iq8M5Nv0kr+
lp5DsQus0qI+f6aW/JJeLMm0kObfCBTfmrJzYQObZBENWShky2egk1NvYgHZfePc
LMlpZvp+6vgBrvhuMuKA78c+zXtJ6WeMmGXFoKkS8J91YM8j4O0THodiG21UJAN7
uZingrhj/ybc0hKmfnmq4MZYTMAoebZNmXjcTB+Jt/a4uATYehIhhkH6f1TilRFf
3nibjyZdVWvyENCBt7i1WRLBNQ9L9AV0RPSVL7bbcvupnDahSjMvTHEdzLF9JnWe
xDsk8GSD3rPZl0QyxfDcJdnrH4V1xMY0FNvBcjtsdFrngJGf/aUdFca4/0ST9C5u
eK6kyBx6CUQafEblyLIPeGFfCPojtprd/VGA9rp4tmYHnjhHbXTWA6+48eRLSS+w
VeoyNCTHioAeetRV0aBfEeC6VmlNSeYUJ0jO0NTdSi5zqFQnuz6eT7FSPEG6+QGM
wonY832rE5pYnAAcR7oMYtQX3FKxP6Rq2l5IFSCPQAekJGG+PL9j77qT4goWMsub
sF37ISatQsL6CTXzhZl14vdx6D0aVZ8PkrAUTdiIARSRcUDKb2Np0eYb+FdOnK7p
NuWQPAoBg5YzMaO9okDBDHozFQRnUm/BJ7V2torEqPRcdj26jM/5epeuqLrlnOOT
0W3FxU4v61UHe5fdFDhl6A0PL2+FQZrkCXHO0QdK51Twg1bSEPWzrlB3NGa4tFAo
dFwOqzIocIm6+f92/cDvEoJe/h8hZ2HOqyrNh9SZzSjKnHxBF6Op4Z1JsMy+h9Cj
u1gyFA9MWr5o8Yc1w+4dhoVSyUq34K71i+TwHm0uoQbi8Js1wrRhErlaGL83lJMx
XlEmmfv+FQ/AMJv8RBuDph3yrdb/DooakJcpSRLHoMN97MxCC26rSKQngW5fkBXM
NilXv0m8j3tf50RyG5vEK1lwrw9HRmM3vNx7oLTPMWVYEfUa/xIQuqZhCTTXcvtP
msOEClLMJ9YG+/0aI7tD1Acupmwblif3OVPgof53QFvNAUHioQ1688R6r1NQmhlR
yrVXO6myabsfipXHUaENC4axWZwHdNHlanlfsvl9spVYz5SZhjwez8mz33kIcCVB
Ez/MdMxv6mtFm+nmuz6SdiJzvyM0pUY+KKd177YfLR4F/qPuPsxW2AYSht15H4+W
h1o8w3hHmsErHI0vUQkf9m9GcuSUDiF0WpP5L657qSbzSfK86y4UKdwXl6mLY0SJ
DuC7pfJNqaFqWJp+90FnQRVeHUBfqTnr8WlgqsxzpzmA+Vn3AL3xSnWbho49ahRK
yTsmxaVGpdfYrFFKguFe90f/Q57zGEqD6dyF7nggwHE1FloLDFPvvmUYE6Jm0Wde
UK7n22cwhAHB/kgsyGyoyF2Jpow6oJ0ENrSwcgBSi7/HtAqgEPTvOUblkGOHaOmR
PppR0xy6mGB/KQbIX9kxY60mLRqOn/zloPe2WhLK2A4o7omRegS/kq+5K7eQzNbZ
Sq1CN/FuMDbT3WLuoKiO0WoXGic+7JvS8M8KVPu2oHzlSigCNF0eCNfxynY+l7CC
2v1D4DqslytqYWy6/rFv9sKle7staOY/VrKPeqOP5k25EBKRerm19oDbM/h/MDTY
sJ0EsJh+bwSx6yVaTBsD8rDMdkbX/g9p96KIY1rjBPzCJxlqBIlbHxXrXtIOx6lK
Xn/Gwc4K9CZ4asoRPGX7t40yLttYErxd6TDLaVs2986Hic2ey+mwFaoTpTVMfkNV
vYw5o3zDrqEkS0co0He93atFybH4buksbaN3z/waPRoSp4VhYMSnDql5XM14Tl/o
ey95wJmwRN7LIsIx92cLvf30lzAYnSsrDumOHXdT6hGQNTikSCJCdA97CHlCWc8d
1BRN/ZSv8/iK2UylOVG125nbKAmM/RzsSv7hYLm+bfMdkw4MkvSKWh4qMpbxa4ev
l+mbK59U2IyhBFfZB6IAqnKKH5TfjiTZM13t0zka/EY6YnmViq4c9ooyF/iRuvxa
QFoGh0+e51kf0GnIOd/oYu7dqmstfADKDmMkOYjLWTJ5o22bSVGHOY9cihFB+zi+
3xoyU/u70O3u6QtAqYm/R6xKneFpPOXul1INabGdWGhY0esAP/QztGXPnGxYkJhf
759rLMI7HOqJhtJw4pDV9AAq+GjUbuH9UQUNo99008aXUoQ+23rIr/M6oWELoXkV
bEIyLvmjb3ngLPnXs19rYFOekVhm9uN89PisedhL6mELNJivjugwFL4bal4/bZ2v
mtuFq3d5hK+jicuoC4bNSBg9QWZD6FmQBFuNfgbBgYSDZEu24zxGHe57TAnPSvpg
bTEg3+UY8Lqx23CX7vKVmrX7QMTSNPMXdhPCe638gbfB8Vl/gGOLTv2eRTA9Vndv
gKbiKL7oaX7xMAvz6FaoE4EbaRF25Ix0XSy/yJ/BhA5ofhcTAjIEK+xGr62yG6Ia
1zxwBH9u0BfRoRbgkylvrP4DHpHBYfYY6gKH31eqA4dtSaCNNPGxjGRQskDtuoIu
rIbliXKo07kz4SievCYegyla7KJaKjY3ZS5mmpRCNH9m4GTBhxBvdzlD3juHrWB3
0UiG5YlqKH4hRAz0jP0jYnSnVwDald8pqPcnPRtAgLB6WJVkiO8OLhwfTuzgFPE6
/EeiPXVxEPnDDM5ke3fInIOZaNY+UuLNSPzp4fOzRRaoOLVIHf0uF9l5/ovJTN7s
rCEHfSSvXZc8pRC34CknmZw/Uv0ovz2G7qNI055KXPpDhIuCIqtwXwyNvZfJOLHm
KG2XJEgG5uRz2qiH3TqQ3MZOBKhUdouvs1fXHM4rX+qlzRvIikSUPLmoggK4tAxh
R13he2/XkL7DPJUk9gYkxSpFpLlJVwRZcIygx6+YCluc6nsUmU5J9Cs+4tf7r6oi
SiaQ/dIxaj0EOziaFxq2KXZH3YbxKyEPcXWieZMMSC7Gb/LzrbZEx5j5hTdppM2s
e/cvACQmQ2uMY2AvHeYE6ZNivMgloAKxol+0ZBqwPSMh/8yLtZtKL+4HUv9Jbwsd
hsPF5GLX9gT77Jnyp90ptSIWTNJi3IeQd2gl8bLVowECI1KU0sWLi0RfBWmcw48a
/UGOq6eBWfhKvohPmvxhq2WW//UB/doLX95aoH4kRe3pGDo1sMfylw3BQ2QCO9yT
ih0btoshuGJBNMyO70YNWgzBT4BqtFU6n+96smcyjGx5XEVdk4UjxW/QZH2RIjYg
EXmAaOfI78Na+73WV/Gx2g0bsFPKijHGVpt93EL0dhryJz6ujO85a2zOR++rHZKV
pndxXVRcZD+oAV11s22ByRNxRLPOw4Fzdq7p5KS5suJRepKBsBvrS9svIiEEisYa
alQ2rCjhX+GzzLXnfeiTqJoLzqbhabl9CCo2sjN6lS8niW33bl/AEKWf6BEnsSUn
o57V5u2gqwGsuEstZRrbSVTQq20qHjVXuy8BwjYG+uaQXes1Ccdj2NDR5d4aFPSs
SWYybmtQo0oV3lKX7hpfSaFY3AAffb45mVQhsUTVAoQAm86rmqeLdYUDfD/YkGYv
6iKc59tRW1Plba+pANFuMXVa30PZSCiVGY31VhYvFtJWWTJzb98J3bpjwwHI20v8
qjm8bs8HxQdJHtDPb3cZViC0hG6KPcnsaYyA4j+0SkoyzzRrEGN6si0c4wIAa6Fv
K2YLU5CAaDoWiP2dxUmETkcNHi5V5G6vTJ8gBgHdEdxlZs+kyWg3zJLWfTfqN9Lk
24RH8OkPP9/KjZULZz2a2/fG5XX6cduIUKOIi+VbeDWhkZTv8iml0AyVyMkISJtX
XfdB1w8fQcDbrXq16MxG+VcPuF/9KTS0CmqNCc6UzSwzG7Z5FfIh4j9Jc3zbHO4V
168Fkcxw35EWhGiEwqfrrjhKiXSsP8luFwPpPMzqoRONsFy/amWr893OGwxaRkSd
KYocQo6lKuSx8lx5qRU0EPEvhxGCeKhk5cq7IMMW7LNrYhWmFVllETYDsVCz4FVF
sFZw1W1jQvb7PJET8IA+rA5OWQb2lE0NEL7SfEeaJav/E203cQPCLO+wF0/zIFvu
Md3Fuft4GUYj/fU9B6+ELjl7ifupLwgrq87u7CS4IKEt1c891u8hfaQoajEBNDk0
GBMvTX8exQEeM5dwHGw9DEzKKBVxuZ/uF732baqE75AAXrWxbkBCZAxAqRqrUFJP
LtQyawHFVCDrjjTer2dKGRorQM+7oSgPefa0VL6sQS+G1v3GQ6smQOb7LGm9eBaK
Q+FmM1adzl+fHZheTPxqK/GI7Qwi8wkcoIwblSdvP+o3o+soMcaL+MJMaB9yxNCw
gi7zmhDuI3EJNfP+upci2iFHgwOU1CabmtOwZZON6Ih4gxCwzTHS1mNSrgFkafD1
Ll+Sca/cNzCEBC20pO5ADAWFDz88tHdFIrVYGIPQF1x5skuiMUfa1fKeMvCz/x2l
6ox1e0jEiblSyy08Hym+MMZXrpDKsCgMINdxOB3Z7iS51SmJMgG6ykGRZqNipzzw
XLo7aILWOY5XaYIOkCRVJzJHiV/MPeMk/xucXO3KQreW63OENYgeSu+BDIBjPBK0
O8wO6vpztUKxjpcqCSHu8BEYFmVuyjmLnbBLTykohhayllInTCogG1Z5FtNIiZ6t
5AYmdGOaysZbV1BkZ6RI4wNHLv+r/e+let2hRKH8/CSj5bSxrJ6ZZeEcuC7hW/Ju
ItuQr86PgYYrumU6wdyPCgRCXHgAjg2c+domlZ+7nseomEVS5CNFNCQMHbFjGlGz
GqTKG79YrMXDjfUHcv0V2eauMvE1t0Yys2TdBAaDn4YbPhfmGQBbqGlLw969Dyy9
LKaMPLAR+iVohAoj9i8vWporDBoA/or9/XW7t7IM7v1YkPYSIpAfXIBFgS52mOf+
7AAU11lAZg6vA5hLf6Ne6TyY6XD4ae1k59klj1PU7FLEYBEYb3iPjPRyh1Ab+mbR
QhPkm+y17JeCCjbl1DrSw1duSczhYtyvUlWdRUeBA0ONLtF/Q1uLs9XJUvjTTj4G
o9D5TCOsy7rDKpKdLqTZmGvIeO04OHWOWH4RHia9vNns+8dkWPeVczVpCUZaOOWE
FtCerFlaet+/rhjQOyudwmmUEQyeW9sUWEhQMgSluOF3JTwUETQFMoSMuvDTsAiq
1anb9gXSdDDISIpkaJTHZOD7iTRZw8HFTFV//8qKbZNtixMCWqWt8xd4nqa89qUM
J6Lh8bLVZ2uBVqY+iefTFPpFk/jATZKZrL0Up6UQxXA0TJNMccpIh1AEkk4BKDg1
NgrKJkBWwFSRqb+e4AQpR6zZXqy/WFLi1m3skkCtDdq1IvVQSp4Ht0SIq1bKNa/7
vCTVfjpE/lA6JyDoyN0RXXX9Pqp4IOO4eqDRGLJOsqVfsicE2znLy43llPGp2rtX
BEVwSCjrHXYgGZdw3aBW3B8rB8gXPGRoMpZAOhrxt0X226MIXQqw0s+Lvylc2+jt
mHmTju26M9BQamfAryrlUC70yVDUHQqLls2Uc627oqdmqDnxrnWqGJre75rIhGOC
mFdkWEMo/Z+KmOpNjv/+S9ZVGcr2CMaleG1vtYAeebTqIAry0y/PRbk/P+tvyS+C
D7WKf1ArHW5E+uWJvQtqczBMMAiqaXAbjhgm04U6AluupNxeEtNe6JHbgBUUUjpS
ozOvs1bMIQxa1i6Jy+tIl8N7NKHkxW+Mr4/B5j1kvF9MHwPG3ui1jf3r1mBVdkvN
1NAxqQqSbuSSspyciSlzOhmsN1SQHqsMerXOu6e2DIurapBMx6hCKeJRdtCgCWeI
0SzyEJiYcgtsm4KoUTyD+VEYKCqdjTU8teXN9gLlAfkDMqnooqc8EvNSGFEXTX56
AGf+LHGGj9nfrurtbsxkoj9mp0ML/IRhE1aMD5TODtSS9nzlyctuz/Ipqb5jvdc6
gmJY20/XFjpMwGofIZ+udc9+1w60txXF35gYCJTh2dg4JHtvY9xh81cNormbwVY2
XgykfZMZGAbf3yfVa3OM4njB1kZWhhhYPabFb+HRvqczH1TDjH3jkia5wodwHK+/
IH7+pTBbrMEmOIDjI/ScNA2zTnBnr5c9P4CpWE4sWQdanW3iNGPT9q9s1vYOk2Bc
pDBe1EBPuUu0Yre2VZ8FMa1FvoXTvszAappet+sZ93QMewHCvLlo4oCWmd77sJIQ
FMaD1XEYdYbyvDAHbsC/arkiPNcZ8RwA1mSd5Y5SRj45s16M5mnQLn0f/2Q1nkc0
KJFpKDaAqgmuBbNp1lvYCUXVXqfnDbcE3avnRDvAyUFX7SK0p3Fu4umxGSBhfp7d
E59/PbLTls6AcPP/2STBK0VS4JLdm+y5Bj8/Nc/4aaDyGYCgYf0lSprTDezF1E+M
Mb3ZF1hz0twtVqlexoM8R2vv5/97YONw+PkQ0IqIa/xKEGJ9wI3S7GXoifOCLwM1
08ptDzfg0y2svmiyppyRvQz+HHVQO3RXZmb/eUwH8Gq16Zo3R9s58fBdAZWikrV6
SdnMGJm9Q6Qts2E5UqpyHgGBWNi95zxgiyZA8NHFHGmITv34DH08YIWyH0rZsECN
vQYnbAwCDVl560lc5qtGHOD0RfPU9PhvpkYmHf/2nEqIivfokIDNPUfgHlEdOgHR
V7c08Y0jJA0DOcrsfJ47RNs2e8fYpU/rmpVVWA625OVdP0w3RgG7K1CyLPUp/Jaw
IjiHRnO2h/Mbs6BySVCSWbbjlkPCXGbSeBBL0izPxo7vkyXQIeCqf2xZjTjYvx8T
N3Elhus1a2FH19f9WzjV6+yZZvnZq0SP7IWK+oyZr/n+adifKfSliEvjHhPSTrSF
jSct63NYhs4WmbaMaBw3q3rnSNLukVRFT2KzroEhPrsCncs+qHlVLVgIL6++rgdm
4rCkmrw1xfV4vTfKTHxOHMI+C4St1tjGULueaBT25qpEyT0uPMfdxz3U/NxPAiBW
/BT9ssIgg3SeWTghKXlz0MmTuIK9aM7dH24JxlTD4BvtUNefENDtdpk7nJRZGktm
l5fE/PMHp+lYVt6ZXVrwHfhrzCphEEiaOcpEfc5lletCuOJ3b5o4BUTZXRS11FFc
apFTu4ZZUCOPoyit9yunnCxcCYaWyPdgaTfSscgjixPt7fU44MuED35jojb/E8Xq
qOFfvuLLtmpWrq3yCX/X3euhr/ClTnGwPDQYO6BH2TtC/1jXAcWM3TKR5a6vdo3+
jqRbpYA8tDL9yJrB7HmT8cI8vscf7WNnPgsRgtYVGzOrr5+BMYA8ugm60HG9/yAR
Z6wrJ5WeY8/vnPjVSSqGHIR+JDCOAlOpdY2eIb3eIKuRgXPswfoasUW3e0rLp8pz
7trZTe+xl3SYYqFj5cCX3nQadZrWkQZua/3kWPlidx0fD1cKwfdaUpNQ2lbcmqpC
RRoxKDqKoG+DQ7EO59sJlnsgXLsjE2/7Afge2pK8khXTsESy7IdN6jpGHSC7eu0N
6YjQtcjHmmaPsMxQiHcmd0rZno0F6Lk9n+7dxp8RUera9UNVjeW79jdlsAaZVDqV
DeG1OTvq5ORiMMlH0X2F6akPuUhyAMytf73HXSFqgxUYtk7l4p6BsXx0EkqxTRnD
M7ieN3WjhHEWRZcQ599gsO8BWYoLfCuRq4INE55eEjrLOApaySwAY29U7ZFruIC9
7FHHebzbf03OoHzVCU5QYlnLb0ZKXQyN2dzAFmpLiNMQoGa8Exw6NA2kolY6yzIE
vrMbkKDsokrZiULsk0aHqUXK1kGmm6MIzjyOelZVxPdJxbUupr5WZopraXG1ePIx
a9xOTaYNR/2GlVuXsdieBIHBYDbao8KtLuDCUAFUtpKfB2WDjVl3zS0VtiH2loWk
NJ/Uc89rozGYoNKjw+MdAnMgF5XRgcIXQguFD/seN74iFeipc0Osz8x5AMwL987Q
o3Zcce0bcZZhy7JrK3vAad8/ZOCv3Izat2c547GhRP7t8Q4k0vsvH/pyPNLtNlU6
fg28VBzEpimn6o5y4aFU20instFvBO0gDKymIbvhrJQYIofDr+AwXJqen6leIueK
PhUHEGMXEBxYVM0g1/ewN1xtA+yVjO8bmEYI32OUI2V33Ize3dO9pcjIeyPAco9Y
fGcK4ZJFI8+totYoOALl2QwZ0vNqQaffxRCnaQVC8ZQ1ioSibIw9x9HUOrlwhj4r
HotX/xks6Pxjl/8eg0eZfAwGT5a1nocqV0pOstmxDXhUCxaUDJ/Qzh5sH5cZuL4b
30Kt0SfM2Bc/WEhCJgLzuIkdvlvol+jojioGtSnIB1Y6cMg3sJqnnWfgA3Pn4pT9
F+RjIxR6xXfVj8R8mMFt3UvTLIyvCmNToKItguzkbDvunR2YhFU9MPmif2c9xcBb
aqLzepsESOssIHJTPrfPnsHVpz67llV+x7KrLw9JnToMhqQgQ3snTEnU4wzI/WVL
1UYeRUmb2nF8PyapNzJkLw2xup7zyXRI+s9JV8mc1bjqcL+JzLq5Fse/4aRUqZy7
0g/uc1nh6ij+iVbcKeXD9rv3BEMotcqG9O8V6N42qhbZs4WSdQqGC/esGQjL28+o
f/ck/229r9ZOTCbBOiD3ARUXQw6ztZglpC2bMvvNjIrj2RbKL05ZOsMG7GovhjkC
p2cWtGeMwpl8vZW5Tqs68wq/qaWpjpJ+XY4ve9BZPxk//VoKVsw3nHHMACgn+mnC
82IlfKSSGWoGrBR63LipTJkIuA8q8PjBXWDuZML7lFxoIR6GV5UHY7DH4Oa1ezFF
xNYXGllcGfXH+TBELoQxRK8WXjfne/SUK6BUkWDaRAPRQ1OP8rG8voLlhZkP7pxn
PoZvSA0GCIWc6GFIptgGP0yBIEu7Mk/nQZ/9oSMstegARmrfaXsAIKv1boJlMO2M
H2sKzV3ctOXfJpt5fR9on5CyZl983OQ+Sa/ZT7YiBHHEa30f3JwqpTOOA17ymaNW
Vm6bQIe3OTYhGJ0G3gpP19nQs1IZiViZ9779neNgyEMdHhFSgli3OJGmQWqJJC5K
q6F0yJgDvT7IiBMR6Peg/UKXpcg70pXi5fYa3eUa5h/KyHAQvARInBS5JzQsqtQf
dsZebfAbHkgMnb1Ijehx4uvHrVoPHe+d6bcJ5Wktjn0+h6bbnJmSVR1z8Ry/AT2q
tvLoqvFd77IDFUF7Evycecs09cxe5UOuKA/wpArBLnW7CI0wcrQm4RhOrcoizjTX
vnOzzzio75b4KJl1y4l2qsVSmI4dackCg4MJ6aR5rkB9Ma+suI2xix525GkQgC/7
HkusAYZuox3Fq7skYZ0+Y2+9QHAX19CCBkNSCEIfEGaU8WEM9DskMjgtorvrorBK
HxlcCseo+Ub1/a7GNmdPu6dGyHggMRRSm7lv3NxZ2XLxqGxBSh7QyrW+0aJW5veR
MD4jB6bRzSjsQW5kPUoBJJzukaEmEzUVRcX0YOOV+3yGB/8vxYjHY8FJzGGh/8+6
fYoO2BALh9j3khp3P77Df20eAidrWj7oo3S02q/yqGviWv+Eva5FlwGih4QRr5eY
X+9ELDe9e6kjjYz4v14ztM25rfI0B2jmrLCQaYmqIF3GDpHrrQBJ71LEb6w8SoKH
kax7xEelZjqws1WQvYVQtw+7is8zycKcv5MT1iTo+gzzRGoWN+y+2+aqCo8Yy6O0
56Wa2dp4OnvvauHHDQGi9wP5h78SdX3IIwxsFy1HWqHVQn15MVbEcnDm6gGWa8V9
9zijMRvzOftw62THPwVEdZtE+oPVUYKAEGMryrHepUjrAatfooD94CEp9V9m/Gw7
NgY8x1RxGbcf2G432qgmvq+mGeJHIdd5v1wTMvv+nJS83B8JHKn8CTo9DbhTQVpI
UkZzIJuQJlw7Dft6hIt22lk++WXTJSP1Q3PNIZ1TngvqcsbdE+hg/uIYU+A4jRib
5CelXi5HocRoi2sU7CjphwIgGYHkPTPUe0zpmcC3LecZHPTxOqwVrQU7U2JZ/GJp
CEWH9eDjS6XiQmuy2MQo+Wd1OfrS+Hq9kOkXckw5VS4eJiQkn3q5QsS+adVO9e2A
dAcGiCeQ/6FHKVgCiluJJzovkAAfoTg+bBXm5EuwbS3nbShCR7PHhRTOQj3UNoTK
c/7TVo4sEmINrnWN6XjVlCo+Vyiq8EXs1ERSl/wgZ2h2jTT9epLYs40FAPrzg5Zf
ms8crJtiIIg1rYyOmlb+CM7kkEcQosz68/yKPyWY53SER3Dlkg0mNAMU8Orap79+
U1MDDd8dflbXDtrgMM4UJ+SGU/Mj8XACqSdgCC8VP6MjoN4kmvYatNZXexROTB/1
g46NUvqV51BsIE5rNozX1nb06nCp48E2rSLeeNEsZtfozY0PmVBqeffHN3e/Cu9v
vpO89D/dr/MWZBMuQkNpBdiw+gnk8K0S+eYe0tTZtfOUfSgGabCs5Sw4eN1I+GVC
wlnSJ1GBBGqA7uvHPSMdQTWfsnzbBbiemTIm30CmQ5MV/HPLWQUpi7mg/NqG8EOZ
7qZQTorLNRMOyrYAGL1XQbPWNrpuOI0VvjFdW6zwNeioFyuVHJggj96KVbAH92OR
YUVmO51Hv5RsuANrz+sB1A6jRo0hgbhATcl0cRrcG7aozIw7A8HcZMKz64658ScF
PJao/Sbqk3DhWOxsm/EPFHl4gzilwmRAGWeybypns4SHNNgF+vlY7xlN5LbHmSEg
8Vg8AQihkrXHS856HzkiiTk+/L/mAyF0WTUYN51LsL08iet08i5RVY1MCDyQmFUT
iAfc5+i8qrPJSwSnvzrxon99saeR8PhlqeKVMxcB6hzt04TUMOH8xDQzCsWDWhoQ
uN9k3hMc0OvAdDucIJOiFLgSIksYKSQLbwXUBpqVSIrQxzVfgBbgmxqYhgtVdYvk
6BzdFBAUnYL9oW3ooGnNFmcufFDE68Zp1T9kq/aWbrwy3COsgTa5o1kZqOmjWmRk
aJxAm1cPnNq0+wEVUdzsabPNfNQyG81MEBm84t1jK+lqQUXKyaOnAR9NX48kMNbC
Tb0jtDsGI49+GY5Z1HKXuUrAg5+YfYgyiO7p9GvCckV0zomuxfOofPnFvMai4h9P
/dkFjZC4tKUtqimk5QPG77ZQbcJz5sL3aUd6RjtWq5YbUWM62XV27l5Vcrc08GHN
4L8+/ovYTNkdae5upvU+Pmbyq+D91XlFaxqv5+hc5eGF4EMShes0stxueBlGyP+E
DMBZh93/CO7C6R+0TSGuRERmmfQhlsAeQLDf0fBjS0SqTgZNdYp99Hu2ijaUMjmp
ygYxKiVONpf7vdoUWC0+Sq/wK4DaoAvqD/63fIIZplGb1sqMWVIPZLE9N8Tot91A
piO/Z0TiovKXMmM9j9dSzNPAMaih71xHWmtCCznFv/481F3LMxTumL5EiLYTQRWt
t8tBM+sGNzZ1qaiGpfnVVEMrHB++yUr/zKBDV+FC0/FBVhJ7csvP5LSvY4d8qkM+
RZqA84HvWVkS84CvjuECrh9+Zh/AQAXf+nya/LoCcodVL5HnJMOxCNH/Xw2aKUSZ
qd2yH1wJEtb5yd5mVs/LqjyXKDhciLNYdin2wIzXltCluSfsgPz7Ub/MQ2ragZki
LpalZAHEAQWTkzBEUmtUXlLsCNzcGxyrl0EwCzbiHQkuZV+SCRPh5LiQeNJpG+3B
vfyj63tD+aIfPSxPsCrjXcWpie37Z65Z77MHZyGot8B1MvISdnv6HICI4Ducbffb
mnttRNkxlY2O5TN9RE13f5wqD6h26lLT/jACDL2TOvIVi40ae5uhJcp75I6Wf/bu
8GomJiM1cXrf38p0dM0qbNc4s6OAAuy4cWLuCS6OBAFFD+MecEjj+ajKDI5sgPHi
NwsPyv/Z+wOV+0UpfDRNryqUP2OUcDvP40U7iPtCAD32N90oIJUBopS7HDUUar/e
h2T39wdq6+TPkmSZ+yN869ezUCguGWKdhPcgA2CKFEIyB7jbDHwbfU+pdtHQCW5S
oAgmURpx3HjMjtS4RprNAePBwIjG6a85itsZz4TgyYhTL4QSRSSn0ML7DtTo1g8Q
VeGkL8ItPTMNuhIxZsE4be6tdIRtDcW6A+qH2c1OKKMSF5qEgeiyZu47rfxOD9Be
XnEM01yLDrD/+VlktGli4rRWX70tIhGvy2DdemykvPEx36gy6NqQuf0ODy6th3xY
0v18nO3mdAdmVPH7E52DW1CjFzJd3r18emoR2yflyC0J9yU8wTimNY+nXq76MNpY
cTiMpfYMWe5VOB2gjyXXUFKHgdgc3IRGz9mIicyAmJBeVYok6bwIVQWMf+fNLI6G
jdrb2VizZJlrpoVNrx9ApweCK4Yx1CgwOpdB9Avj0oEt7WkOYPpoPdr1KmyKs2ik
3k+hLBUi1GlZ+DqnGNRdS4hcDqd7DZJWjHAdjA5SfXurZ007uHxe0+YbWvTtKYM5
T8Nvq1l/B3Jnz+SBsQ8eWBJt1n2LmBRZvsW+k49XpDdb8lfDZU2THXzlcQx8kW7k
pco3pKKZkxQ+iKtNq6DvH94mVenGMTvhe0Qsvndt87fzsV8vDF93ufG0n4lS3jT2
KmCw3M3RpPUouF+KjgA7Wa2X1GESwewQKB2MRVGmp8kCJcXiZYfBmW1VkpXAktnU
xeOEsj56DbOrbsaqi0Tm1gAfAQWitGMCFP2DV6uaJAPvX+7udlytito2BRfU+Cqe
Sl8E+Pn9PnVWpnrdUBDl7o1PD6IKaJ9GPun0do0OEF1DrBwJfuhzZ8sS4RVAvv+0
5WeSp3tAkMbTBvTELJvWpz6uMlnPnxJedP400FNJDlzVKYAvGtPBPWs8qbgLTGqQ
2k0CQmLP+5JWRJt0EN2BVlTGh8MVjhQolMQy9ZBSpLOraeD2b0YzNLrl0Q5obbFd
R2ZGvl+Lo2EMVi66echO1sapw+/T1XoyIXSPS6oqjfdYfU9HaT7wQJqFiwzi24A6
mRqhLuR6kw8YGtnqX6GzhqiuLpzC1nE+oX6W9hI65L/TlczwaZgpNTKhqOQXyg6d
r5QmPHtqBaIJXWKkYqG3BrpPjq268ZI47lxHQFnxP64wwyCwlr7AzW6C40Puloxs
bEPA8nxgl/GOp5fqCVym/zmZoyh+zIxMx4tytaf9dDSYeFUImLH+Lj6RTeXJY2/+
+/Y8p1yeXxV+PWVcWrwjZfidI7jFzvk1xRTeNDXnkQHTPjktbk8lxuO4+56XuIVl
mDEDNAPmO27xLsBGJ53dIkFXdzTxBtXBfxVpRQRvRhNd+nkP+zQzhW/2rbbO/8gd
lF2h/ipcHCfzFVCoVyUzDO5sDcXK+/7+obm8dZvylNohzcjZMLdePCrFwNCr5jLf
MkzyX6y63E7uKU6vjmChZS1XamOu839EDl+KGvy9FUteTzVXsFKGRsVvaaX3im6w
dPQ19Pv0zcO+WiqInUcNTNEaEKGAB1HiccHXv0gz0WrCQulcaEjM1ql804t5+HA9
xKaHDB2yRfZuzhWJjvKDqtMtcQBJ2RfQUJDx0DVQVoWH9liHCElhPIU+n/ryKVMd
eF4oRsfHLZdiCxCLImVQ0mhRdt5Wbj7RVNpqsULei3tUw4xZVgRLkHkrEoGlqPv6
FNRRk5cpB59HHZOd8H4nRNJI5DeIedlFxBQX1Xfmzmevvus611d19En6eGg3i8WE
GAe7E9ETKMA2Zil5VNts3QaHoJzA6qO3BQO9Lo2QHk4wa2zuFh7IRJUbec7WP57N
F0swVECK3sGLOCRiWXVnwVkgta02pax2pWHeVpMjwZ6qABQ5eg5SZrAqNhoeoBTu
riG+mxZaVXqa5EpXEtELsEwU+cXIRxKzUDi+YwGHoJ7QjWgUFYKIXyUS/kO92XOB
OIK3ZFIcf5I2DcChiyFr56XlPauLxLxS4uRsxNVelgSskKydof1DpHA7OeDqyQlA
EOpFKEdzqE9D2B8IrSD2Kk+VlCCVjhuU0WzeIyg9w7RySyw30epDHL2xU3hMIzA5
A4/4dxtGnASknMx59FRe/MG4J15CYndU9tBXKC2Qh+X5wrwaq10Fl9q4ITCh/LQl
3KINrgC21DxDUTAdP20z3ClGd8qRLc7CP74zjZ+zJyvyg4GtdoS4NZtSGdxj1d74
S3RnmU9IrqcIstsyvFp4HS57CS35sIJEbe/M30QS2i7znlesgNsKJy+LcwBk0Q37
5lrpocvISY5hCSU8mzZOGMPVohpWU8UHFd8cMb0GKENh4lmJTK4uR0+YbV2t6z96
+8ShoLgjXl5Swc1DQzVBIxWLXOyJJw54V+YxcVqqQvaEf1V5QzDcxbSybWrNg39G
MvVd+ce3WXGj5mUA4aDU0QM+ZAJpk+FB/jGQbZcrKlrbLsKuHP844I5WzUsVXTK+
jXGp9Y/1Z7Puv12bcL/oZWLOO4lO0G85/A+k6giQCYcXSWCaB3INcmyf1NH9T+vV
JK7pVJXDpEs2uW9K8I17XeOt/n1tdVmMl7dGdpjcDHedJaAp00DGLcEZuCkLmv09
pWpN/3GS4Y0sKZugafLeWTdLvFD+qu6r761xX+ikNI6C8v3Gal3S5G+gl32oKSfB
SHrcBLORf4eGj/LAbCYJHTfVG6cE/+El0eSUdJRMawnHdrn+J2B4N7RMOscO4j4o
exoI5rQYqYXpazWdBEA2yAq5oevdeAOa8EVSCqo0JF+AFhJjb232a37tB73+FAHr
HvwHwJa8IOZiUh7KTl4hvsqwmFp6k9duleSoyeOQYsilSOP5CPJbI92Ns1MAOtPp
MDP9KTDaH7ZKBl7Pc+wLfVzga59ypLgd/HeWUCkAiauvDyElZOd0qY8xHDG39oMq
1E7deVfVYYdT14GAvYlc7kREgipzEibmH1jdATaXrh19N8k39LkoPY9gNT5t53BW
2ZmdCguTDJKjGd1GzGzMf73o3bdgdtCaLa6Q8rXObVNDmaF/V33m/M19E2Q9XK1E
M8FmPYIPPx8v842i2VjriLa6LX6g6OGNP+p2st7y/AZgNL9GUEHevQpJXO/f5IFp
uS+VVNZV0wZcv6YxO3R4Nm6VGTCCzHWBqhAaXAxnO9KCClT+5SgTQ5V7kegITpGS
R2+orIeQ6lit7RD80fcnZXTI/WtDRVdu+e/iDFuKzlxp7gjiqMhvN4ZF+uemAbvX
j/3Cu1BrDMWjDq3ziP0zr+e5Bp8tKs1SwsD7QnlM1GVwDkusUkf7MXQFtbaMkXNR
Tv5ERr4i7YvJfsY6ZZQbd+oVqBUN/Vo3glTTdfXs7q9mevTP+eBM9rN+kQndNd9U
6folRRTl31XM17aQuD6qvSwzcnDT1VfusG5YR4rLYJddZk99ga0aLVc3gdz1RSHe
YaByQBHOM7lzwFCxeHGrNBsaD01OghLU3+5W5fRJPrqa7uEGZlbJSK6hmy0yLfAY
5IPZke0d36BYK+mdmF+hXSrRkcdytzZ2JdBaPIJmnzUYR8bsvSdF7mKAwK7kzxB1
gjgHzg3xO/vqcYkMKuOLHaNEV/Sgo6Cg4uO1deNH6EsyHEr6aYt1wvvtyte/QkgU
yhmcOvqFfsJ8MqEH1wh44IKZJ3IJX3lQc502Zw6ht7JIylcKLGPQyvKe7ua68qG8
VIbofFmIcCfU0PoxpeudhssJgx8P7R8Z/XxCnWzrSR5itj4nuM4WsdKgHXCLGjbb
aaQ8INaxY7VEKvyZudAF4sSsO5mlJ6VNI9I7Yb2wbaTLDEh3h4mvrhQmicI1Oa+V
TEkrbF2IfFDR8Ca6Z/vPGXbX+bWHeWfq6tleHR2F6f7bTpgoxm2UEvIsDAme8IyM
Bgo5jWenal6VZgefjdnULJpdROi/3qlzFZlj4/wwVCypuLx9a3iEF0KeFbQQ0jVi
q8ttoC5prd68P76THxYI0aulcwlXzAwErdWTL7eAgjumLa/PQnp8pYetOxUq6J1S
/PEm6F2HD10Cr1u3vJXWMHcRD+Xvu5rvQ+LfvVWDc0DIhwJ4vzTF21VGmh2DNChB
KqH9EvddAmK0Ld+gydC5JKCgsMSuGShoexjKpHFYA4Zq+XB9bQlKGyk5qVOAU139
uwWzm121WbHzb60mDAHjSaj9j8Fl4fmGHsyzxl4nZ/yT6Z/Hb9tkhTZJycphNqyw
jWP6V3F5mJga9e8tVplmJncZtTMN4TB26oGdnm89u3OJgEaoxhNIzPty4dp+EkmS
wnXK9wR1EfgUeJjBgT9ea6V0Ao8YzR97rnCBVTLzGs/4euXOrVGxP0/jM8oGCu0q
lx2p1BqgFypJTPW8Td6sk68zcCowH+Vf7QKdFQ+FoArKsq7p9Iyjdz4VPL0S/1KF
O1Np/XaKo6Zfe+cVncSLyw+QOYswKSuETaiOnKUPvIrlrdr91Jw0eYDI+tibvlVK
rmB+N7BCxl7L7y1urTX07OKj9W54GqftuF2ulnXrDls53yfNYpcqgBPWxcKsgNry
BxRQd/UFFNF8bLel+J0qHmzG7pScQkp26qipZ8rnLnWwHnay5HzFq2ARHywsrgqF
sXCeBUYIHVQ+eLO9NfvchM8OQbUL8Y2patwY8S092rZWH2XtJTMs3fnMxQMpg0w9
KxPHhGcCRmtYv3XW+eInV85D70pcibFERfeMSKJc0j7SrPq0Bpw50GtLA346Ih+T
lGRAlzZG+K5CKJ0bffhrQEkPvGgEh671GDHY9w3Edv7uFQGLIZkbzyGhIkajGC7z
VRSZGxgMVEhvEH+9cxKyZNUmNVrsyVTe6sJ3VRk4HnxeXE5mtDgoLQAi9DsISp6h
9LYlMvDWG8KJfV0rF04g747SkhEZBIDwEHqIzQUR/rgUMnGe4fW/934r2SKlbPV0
iYcIiOCRuZttbcZdoga+TUopoOd1Ei7seH1fqxsPG8wiaHS1i8IkzQG7CIlvdL7R
5uUwZEJf/ZDxPF+MMNdPtBjxHedrzOO2E4EIvantJ4rXEETy/2M6W8QvdMizZaGx
FumJs5DLDJNe4fcdq7gbS+UZxG/Aj1s8B7CChDGPeNbOofVASx4jUUB6z/yX4zld
jCh9DoxSGJL+Q023KbUBtNJucs2TanBBPiHTCMEuzSXUP9ewg9X6ktKJFwtsi/Y1
2Q8ne0cVCuN/o3jq+B27giA5Uih+d4dJyere0kPCc4J7NgrGI+UI/i39ur6zzNoZ
XTANV9A5VV9U/QKNP1lyJHcZdrC3o/V+0oPYwTJ3fcDQWE52tx0iITMnLl08HU+l
ghjDBQmq3yiioUAqWxF5PygcI5G8mIsdG2ZhNhSu/e8CyWAs6ZCLWxI/e/ldv3uA
FgruGhmDyC1aK3mvlMnZ/2+l076pXa9AlB5eOnMsqd48A+yASrPIu77rP/eGuWDm
fZk/FGEVgDqb+6e2q1FuXsfCM/hzKSi1VASKqgr6GjhzB+kpkL/eOr4q7OKW5CG7
7vEq2+//UH7cgJJDrQJYlahhm9rSaOxVgA9QCJFLlzspNbu98aN90kLEKVs8x1Uq
vhhx7BOKteHqW3rxedRh6wkWKrrdBHtDmk7lli7jV/rK6kDAihom9Ck6BDx7utvc
KFGpel4rdK926hL1h/hs5uRncG1N1+ME1F5RRPHe3oLif39y3RgrEwUQlM48qsjH
368U++X99caqtsY0GuJ6VBVnynCKlGYD+OgMH2hSLmwMox2PDXl3ZO92vYRKr4Cf
cQ7finS4No/I6oTZYmcp6ozIi0SJHXOAhVbSklXBa9J+CbdLWYjqytPQr0sWbrXm
5qNyuneVntMR/B2fdU86ga8sko1EYP7iO+xyspwYCJ4AzJCku31BHlgBaxDErz68
JZPSKsayB6BHk0KL9gSGNQ0d+be86uiAunHoFt0YOWx+53nBJ1Pn5r87ppHs3YcC
8an3t5UAWHxJiuLUe88Hs0y789eUjK3MfoRnxwFMm8h9utt4uY6SVHEi0oocvXHq
jt7F+LX9ZHB0cG8L6BxezioI3ylysCYAeCIKsC1wfFfVAnH0U7JLMTWe1KC++1qc
+E/xd8Gqi/tg+rSzDQmeFty/IrfZUOD4jZM0oSXvM+uz/UCaUdRU6X/E5UXc2MaZ
n6hYUm+D7GYCsezGsDv+sPwfVTGNpdR+Hlx1Iidl2bh5k0hbYDsIWASTZ/wHEzVu
xYirlyYK0sRiysHVvotC3gHCEGINoAQ5ZcR42HgEL8A+VaOOvDzyqwW500zl+SuJ
jYszEOAFClT+kAU6eDCr8VSHIDaFB0AfTWPz2cflOdpQTUcxdXRDa/buNFYbQlAG
C3omjHkfqxsPWEPbBf9qjREbo0DKvRq1V/nAoNhwfyMpFKerFdqudXlqx8rHcFyk
LCrZnAMBQj+eKNDslVtFvAh4Wa+z9zWFLBAgNGuhNs/qWLWySO3YCYJ7L0tHoRZo
vbR1cozc5cduyBje+6SMzOyDjBYf0ajLoyS9qQNhFYMoh2x7Vz61m3mBDTCVCl6y
hRs7xiUp9mvoR0phfaMW7ajz+CM3JdHJ7yAx6riWlRkENTZy6I0YcqJV9ZTB1A0j
vpK45Wzy60xU+Qdz1RMXE3tVdePvCcb9HW4Go2Q9eyFtQLM1SanAnRTeHeyD2OjF
nsXGXJKnToOpre92CqsPrYSP2mJQ/84J2ZeR6FNeLlUvsySUYY3VBXlqgIn4kXpm
mQOdwXm7PJqsLWjnX7efFui58PAJbnCLXbYoZhjwxia6XV/D1fRU817dZmjKHzdJ
UC9WeK1WblsuNmbibwyQ0w6JZ4NFsePUI2hLf5pOH85veSMLGBSpkQLPbgjYGL8s
abtk6Qxc27f+uaGRizJDNTBX2s8N9xcV8MvIAU0/pEZHcPRO4fthUNRvkH+8rNh0
1e2RcjgyB3NvmExmpq41F0McRD2QeNOxErtCxhpHjQqQo1baS/rfIoS51kEIvUT2
7/ogLQ/FbxC6zWn8Zz45/yOZHDJ+WcGwkD+VAco5QGznDaYYTf+bniOIrCsNH1bK
uY3J3iRY72r1kpKOkZ7Viwd5iEWxT7lhanZWdtbNk56U0PhjMVgETu9QGaB1HEuW
PHZ108ER1me5wvlaW6vtGJlAJu9rwsn81J01ZfZADQvJ/wMfiFPiJ0JU1jzKLilv
yFW9Lzrc1N0MVucJO5cNiTDR8TwAer3PxF4HNqhS9cQdlvmuRyFiTJWIwC6WOh/5
45LKODi2Q/jpr1Tes1EBPEEHPD66rhy2L+UFew1k0K2CexUPjvxt56/Ltw5xnqFN
ql4b3JAHITBvwlWrPAttw4uN+Rpnh9l82dIPEdsA4aWAUTa4nkcZY7+LntbNzLfN
hBPePWsTPsddWdz6DWV+W2PILi+drCEjW40XY++tzLl+VA8/JoPJ4/bdRnjTS6UZ
7k9DjrrrGAsQJteueGiaaTpApYbRs+yv6SefXy57Vloq7k/YG4o8m6+KAteSqgex
1GdrNZ0puKmAe7c/REAocYrUWUuqT3lOao4tI8GiUacw8ipA+s6oFH3QugtnTKli
/UPyPXQnYcucv9y//MzD2Tiyb+JuMWxEHpa6SJShqTPBquzSAFuiUkqEHc70Eh1o
BXj/Co6IwadpI7W6PUH7xdk+Rt8Lc/vJ6JkagCBrLqtDRre8q8pZucwfZApzlCAL
c7zWE7NGn6G9Aj7N4yTi3DX94IcC7h0x4dEIweU8DUn9BxcvnpWsONR4kEh5UQwp
k8MWNIg7XSQgy+LzEjvn1NiBAeu7icfMlOxHrU+86N3e+PQklAjijcvcysQRtGQ9
wzdIeTHwcA3v9aGR0AxGSKFZCV3KtjpP/mjzmUjgr0qYwEhv4kdQYz2w78F4VRGA
ZQ6ELBMP+z82g7w/jqmdXG8iUdrTz0HOYzPt61bggule71ZXd0UT3wi3rwK/p+L+
KuwhfHyU56AsxYC+Rk8h79pnfDUiLKmaLXhvlGqmASuZfG0I/sAGiLZDpHasCQGW
vIuDWs88DLtaFNxfkNGTT+FYgOduOhu9gvtpDHdIyMeKgDlBU087M9VZGYWAX1SB
nJsLOeb8kG//zzNP0CKzZx4+Znko9a31hcjTxEW58cMfcnKLFSEn4hgAWUUV91EK
aAuZDUis4VB4aYNo9MMnKABZCTOhu9zTY7w9dor0mKNemgu/Flfj1RhK1KCVkZnk
yUVsdalviOBZBTUI6omNPcIvB1MQ1xndUcqiSapvQfdTAf/E0O+0p42wapeJyBcH
BV8ldXCdCG4gYpyaxsRYF3iJegnds14ISr5ykOU3Pgp12lezArFWIXTv10Ki2xa3
yhoEKwQk/hsWAYy4XAnVoYM0FIl07d0Bv3x+MOu0BOR5f144h3s1/8YuK7PB3mlI
PFtdex/QiHzioa02fGJiEnLX2VsVIsqIa8L5A2RrTnk4zH8p/fnA64ETKOyA4KJQ
xg13ltGuW1VXNhELAwGy7YUh/+DA6fIdpWTS5i1lwmy38Dg4A3o2MvbGrVKShaWl
bdb0G5sNVgiGbDXt2spcqTGpBy+kExwlKpCTGJBsodubPcraiu4yeHqtfM5LdQBy
AV+0eQXYX3vw+kSyMDILmT0Wp6yl9yq5QoVewy3uL2yhog9RtogpqTXHo6ReBfh0
1yiv84aeTLv7xmGafAPyrMzZ7Snj5pmM18sai0mLSZWLyrNhwJw8trGMlvNWYYN3
1pmTRqoLDMhi51kUYfqXYU+xZVETMj6Cck3HiW4EMJo0XWgthn7anXZCc7YEXPAm
mvDvSWjIO6xFWsBCJqoGEicxH1yPyqS/d0+cwfYC8Jgv4j+kIeSXCVcqwXj6E/z1
89NHcIf9pXKXOf+WtXsLGbuYAC+AglDamDg2VTsdBhu1x+Ummqs9VeMmDEjb3PJf
GmkcsYcVT0jHbC7Ip5VX2kAySgfPD0NCweP3RC1OTevUJtH10NhrbYSgDbs7ZnmY
Lbquj4hbXEqUScQvPOk3jrYemXnnFMHMoqwfnlWYq3YWZPohIcl1BjGZAkC0vM1o
ZAdp5JJe01TLEjCTdj3YllLSSAQgY7DbyvF2DCPSmz+M3IDfZdAh0fc23JJ7CJA5
nT1eueSO6vq4uR9zJFVl2Y01aOV6n2Ml0wzgAAd2ndWBHkkihvyMHnN02kxNrY6e
L3tuSv8HeEeFY4AN1wbGd0MJQCHYe2sA1HTPfptjYYODN4XWWzaARKzgatJSlce6
ATdv2YgaRNqc4JZTWdGHkOwoCKiI+pC1IJuTRUf7XuuZx6dBAN3511xhBS3LGtCN
sAovXxkGv4vKXIozVn+iyZz8QQrqtE9ojzZLsyttp6Dc+yR6D4Dw15B/Qd6kkdbZ
oWM0NwZpjgFEG6rWex7X4ESDjPzvOis4U01EjcPM5h0OyYI4kHOMrdZMGifloq/B
vQRk3WxeepVEb4ARl1+YhMHMy/DecjjdAXxs6ksAbsuc1QgD+PcJfy7Jh2t70evA
GObK4qj2pAbafVgeydQuV2cAjG1JDx5ko90eSrvuB63Px9IUhaDBx7VD6r1QBQld
n+1rJIUPpu9k9t5lzwltCr4KBpyDSra61E+ceNSjVwrkz9ADEjawQib+PBjgx9I/
JVxeZVOv1ZhZ+EMTbnR/aAAivhQgLhmAkcYrBC/C0KPj2sAZDWWZ1QnQypvHRrp1
XnCS31xX4hEcSw2GA5UpCx8f2iZDuTeaih6Q8MaCEfNMMFeC8Fc40sxid8oQWM/O
+SjqcRm84kI0kmgKReLqLgJtoRJ1AHIMeYKdm8VapFwJ1PlynrjqiVbbS6rtuMAk
fYWp18/01uugkHANheH5wj6ef1AXBpoKyU+c/27jqPEhH4U2XSue9IC9/yMHwftz
GEh8MO0sxyIuqVCeZckDvdITmVcruXX0MDt6emQg7N2zDWMEPM69Qzz/pBhSW+Xr
sO35xZ1llf18YrB109f1fGwKDJ3Dx45Xsy1z8VtjiOLfKdDz4O8yqriknacyEZeg
CPvj0dMVDZ7Sm+7KqhXeFJDQwcXr0Sw55Z4wq2A/U4CnxqYkb4qZZlK+mkb2adB4
HB2fZ9hJqWTl/D/2sJRzoyBHlD/rxi4R1Se/OXjkphPKEJqVtRw6CO4E5QEiDMmB
4SpEIoCJzqSgzXI49eIZaMukNc2VkFLc/bhcloFIunK3gZdqmrf789dFeaVms63w
UvvkrBpwcFpDRbzt9nQJNoWD/ok/dJC4+OeYpj6uHOKJ3QmXjlUbXP38/36Beiac
G6Xa1JcZOuGR+BNwx+blupi2Yi37MTedF4LBQ+u5R7pJTl0xJdo7Jl0FbESSqgGu
QyWoYUiL6NrqN5uzl06vy2pnT10/RK1G7JPiYlonl7mzpgbTWkD+y/KSgIrBEQV1
rZ2cBCeKsz9dajMieZu0mp48Q1WSx3z4KAqsowd2yEz4Cv/JwWIYCWhfGkZfFT9d
saKPs7rcFLTw8Y06y9jqc5iB8Lag3jnfjnd0Nca7ZSkEoG30U/xgxUifIE9mt9RA
z2bTjg6fR+xHNhVlN0JocUnzLuULh+6WqbVtXq/o4TgUTbRXvQiFn+Ds/gq7LNw7
bJepoaXJeWq7MBpuHZiJvSVhr/olKhyphbbgHCOtgT8S+gIu6gJEX2S7ZqwCK3Up
9S3vEjRCLgCy1kQlNFaTiAUesafv0m2IzNVq3E27VWDaNeMqDOAgts6B/ZvvoF7L
dSBL+LWVRvc3rM8WgULq1VEjcy8P2vkM6ZdLCTYjPJqfb4cRXbhLGlLggQf/zE2B
Gkyph4f1EhtenQt4enWAUVeJ0AGgCcv9HZoHqlNEZ1S3N0frWi7So2tCkHJ3hEdY
IBcfvtpcKf8U1mCKrT41jwce9THlv9Qk8V5UldYVHyAOGe85ujdWJi6kjax31v76
l0mk6KDu+tcD0byrDbbj0ZffvcW3BxzzXBxYPcFDxCu7hWaAFR99WxNGJKV0AP1q
7GXByhtlTn2TaYabhjUOdrgRh8xHNWapoFpwDlBOMc+1zfCb9MIAIpzyyWj057G5
5UVjYqfSm9/ipBTz6b88IOekcnDjksAWhsHmHBhur3n7o9xNcKDUHBDoXi2vR6JS
709i1vc+qitMm4lemJc9jPArMWcK6KuaQO1rT+6vjHd+lWJWlFcp5yvYqTu84AeF
28pjxZvUoUXDnL5wZuEjS3ifQBuwB3T3W9nHoyoHeLoJC3euHyE7Q/IFVlHnpski
iO8Vx1nz62NCO3jQgLo5lPujuZ2WA0XIRE/2oGPK+JADOG1sdpKzRITQszP+aCdm
WAg9Uy6u9+fqP9XRk8WZUAgm/xBGP16N9HKG3vfX4mE+niPtK0Ddp0wMxNwvHgXU
MauMQav/i2KNs7wS4Q6rstaBUV1INDJD5xWoW/dtQb1Y/7VKccxXDo1ue88EHzqa
cfSo6f0aG5B0lApDSPdaTPk6za119acq1dwzJGj9IcUNvH5YpINPgF9GnNNSYWIV
brvZzOGtJc9Pxh+xS315SW1vcRAo8UpldSwTB/OJms42bhAvCnJb6Y+uW8IBoQT1
3QudkLVy1L7xTCrg0o5MUjz9v4dqF5iwg6IqDQN/IKzm8ucKJiNhpiAaGpo/7ni5
5ghzjdo7x7skmWGDRncQZzJgHe+U6/BymY8VJIzF3ic2flwlbT9BwqnkRllTqRXd
oLz78AHdKIWYXx9oU4w9wTfZA57CZFAaguvsguVg8Axb5AJNhzbQ/AHMlWzVQ48N
u0sjcul85Jgs3294EKk+v/r3VJGN6OnBkjg5jpCBdIjAQjdg3ozrRi7hnPKfdbEa
3qJghOfdu357aMqlG2qLHJaPdA0Np2dN2uN2UB9A0H+pwdiMQ1EfB0+soPRWTANU
ytdsZDW6NcWm6Iw8FNDy7eg58MJ6rdC/MNivbHUFxZkN32+hg60Zoi3pm4Emvk3s
hpcFPgh3J6GdNAEq9YW93v7VARxy/Gc6UBf/S1KhH3SIsdisFUDpCaVBNTySq/TY
ftBwvldOr0glSG6xO9kAsUNGweHnttCetetrZnRCN5jkzM0OYopEHtYtRoGj1Vj8
rhwAHzkDgbdxI0OAqdDQH9O6TbI+dk8MAT3ymLRgZiMil7uOjBni09JLYhhEMws1
7k1o460jNRQ7RQJbl+ltFltzMwnT+waCnlbXRfuSxjx8MrIHyUUgHd3jyx8OSdOZ
h6vnKjgG/mliWQy9e23slcLu89EfgR1gfXtZ0rQzKXZJKAacQbA831IgR+G4D046
TaQZNBDHkIFsZIClSYybm6/PyIXBhI7jQoqvdCs9+zACmLtBjRFZPNS4OGpfBgdS
+bQPVJ7O5Fjbgr5agBWB6X4NkCflNPfoI1XYnwi0cEacAgG7irfbqiaDZ0AoyFS6
PoFhCjOg97nFA8reYZp5ZqL7Cl6Qu8irPS9/EARLa1beg+3QjZS09pfa6w8FH7Ux
5OQT3E4PPWZZBehxvoiSwO38jKoz/f37XRZW5xlJV0H3QRztdGJQ5PslKmrsxJE0
HwpCZGwci3ndozsOFMg6clxyORkIMCfaumSTLbIdTgxUUmPQhyGX+RtyJhLX7694
72SrPH4rQNmJ7tkIPH8uC3TWEe4YMG18kuaDsyhLvWHCY9AkaHzqsEwyQb71VxZz
O8Ngzv/4IGzoVlxxotCxQHPbZY9ZdYJJpTLt69o6IKPG/C+hCtKgCRLXXRJbZbPW
WioAJ7Zm2mEtJG5H2LQXhQAPiL3HA7hZZzRybIM1qJzlC8NZAhTakN74yaXyjq+s
TeX/IA2rDOgiuqQ0AwdbAAiGZV4o/E0Fb9bNTi7ddOhbW6El5XqD9OlOH6Pn8Cdk
s/PKpP7VGQusyy4Sv14bv6Vutg1WcFLOZ1onEx1ePEyTX1ePY+vlG672kARR/6BG
7D7cLJqTlFvPhHob86gvj254eeg1zE/tYxSRvBdqtrB4MYxsugNAeK/X+muUeeyM
D/KmxlsRMI/F9HBtXPS6tr5qbGK+oRSXTwtZlVyPNOCxcAcUhrWrCgS1+Rc841go
sRQJi2M520BG+sfVfPIujuPnsDOQT1oSPmes7UHieMNWpp5zScwY3Xdk66ddl16A
1SstZT4xxv9WC9hab1kVtmodK5qwoy6rCK773UhZ6IQyqivgSTMFddu0FzfjAQam
qnzWDmAoBFQVf0dT1khPSaNP5gyg0vM9PHWKEmkb98W6vf3bjf2I62DiNS8LMiUS
1IFw4l+E4f9GfeNV+DA+Bc3Un06Z9YAWoQowYgYC9bLXDvdxaeDStWO484A2dBSZ
+TZLfkHTzwNp3VzPSHDTrz4riWA7+76ImH4z21QHVzk6DX1x5prp1o8LpcANKzyJ
WtJRGnzqd/8jXnzqphor08nuSVytyKNY3GJyM+FwsmJbFhcJyHr2N3K4PtHpNk1N
6mJbMl2cSQE0cu9f3tDiFvtQwJtBKzr0v5R+wQEeSG8P0JaTlgcEZDw34RrGBti2
ksMGRkxGZ14PiGW+wh8axnM1Gb2ZLBD0mTqRb6uK9jtfwlZ0TmWubsYUS6q26jFC
fD7f/6vG6M7hlrorWOufEZvR6IzeggxByBB9izDW+Jjb+rBISghizqniwAUtJk4h
vXe2yd/6ih8FkjO8TjiIMJxAo5eZbESHx2qa0g5zKWbW6ASG+brQQ1+4WOGJSOfK
50gL6WvNJbhTyijpvHVpCjFiZDQhvXnjaHmWdYP8Ic9c4pFlLcijSnB/bdMCClCp
f+L3tO2eLS7ONDQHIx1xacr8IoAMWBrRX0AqAWvH//T7BE9OpcG7Djpz/PfmaIfl
L4TGh3KpKL0US+dRnLQ9WlDWNJ9E02JhSltgX3kJx7hf0cw4h8ibuOYr2JjSxtuG
CdZcrivXIiPuub4gIY9HoWpiKKGHbl2h7IUR4PvI2IM30RW5SuCgElv9R8UlacTd
apanaTrYdZS0fOjHZ4UNJrtsbqPfoFOskVYaGRMXuXZMfZs7gfJzmrru/xYktPac
2DYqKK2UEjdzvXObGw2x2/5mA8AWHN0rJvH6fQocDrYCRu1yOBtlb7SSbAyKLHdm
OWtMMTEugSrJ74FO8WOl4E4tc+l3TvhabKHXTqVo8riV+ZOyKGy00UWm7lzyznD1
Yg1/jh3iL47LJBT65kACKhLb5F0ZRS1b0kYNls7T8JBLvOYg2qUuMDbzqXR6+/cR
ZIUiXKlhQYV1kDVmgudpWhkEAWoYJe7YICWs4C891Aw7nwp8bdV96qT9xKeKD2Fu
9ax4xIwAAbFG9epk9bznZOXADxGyAIoNxkO2aposlQHqslCjRGHpII2LCoqM9y+n
nGRg5m8t3KrB7ZREZZq9Xru9ExucqamkBrBu9tQ//9IOHL/MW79aIT9o2MaUjyJI
wdF33pP/wMFYNYcPOV7+1Qh3IgUvZdj3+k60gAn+Hplrc6g9Xs1kHrMYUU/f2BJg
q/x6mYdOQ/Kjplxo2fLrbEgUmu8RSSrKZGZcGd55qvjCjzr+Myta5auH8Wfp1+ON
UNVDqTDV5j00SCsB8LBSEIXtWNRoWloWM+KY7oJQvlks18HzRco7xdE+w2kFR+WZ
f9BckNMrSW8LLdSfOO/sCdujLtExp23wlBB77fNnwHCWrEz02tHn5LYI7ztJJsZJ
/ugUQPpGCwvcvn+xHr/WUVMrZmmG5lZKf55vylROtoRY8W5a1RZ4k5CZTAgj95Jz
atCnDUmvZEPU2vRuBoANxRBULbn3o4hXfTgcdJdX5lTidwi8adrMFIscSzHU+Lki
fDHVBDxmyw30nVsZu1JBz+ulZNG4gz8SD57Efhaumyra0Y38d2A8HFV9biShkCJI
Eb+3+HX2A2BMG/QZjWzWDkGIYi3lHLiJAfdY8OTZBeeUmJFk/WpuwYJIDpLAYxXP
w3yQQNvhWQGWG33W+JIalA5ow+KPb+H2d+g4LUYqAR7uBLoobRNGnEV0J2OIq6U6
g8zv855UTuO7qtxejnXXVG+pZZ1JeMYHfpf917myA7EESrxiVJSMo72r5NxsLBvx
ILCQ/v6CE3ONMi++kt2t9IrWo9+T+wY3RkvVUGjSyGyxLh/+RBA5MLXPZFCaziJ4
gEpOBWNUtaavwVk2f/Nk9vgY8gQlEaawiWwn7e+Cbdcxsry4x9g8vN04Sq7MuzeW
r5VVbt7M6b62lqGBfnrCJay4Sp754whut4h8sxglMCJ9OzoD/x+psHu3lSWWg5nV
pG+TwPNjsZL7L7QHkA8ykt5vOzqQE72bSJ5e68l4gKzlkRlBPBDwAH3M4CKSJIE/
G5hklfDL6vPmLmIBy7hMfpjg68QIfpPoYX4jTWclqqNPcT5jDcfjDxSqsRrgSWfW
UjxA4yXGCO86DxeEycjPD+o1DspJicPb1cobyoT43b6on5VFJmOU3PoSfGQjlyHm
cLoKnvCqTO8u3ayzXDWKWaTeZZDV6Kakj4QLIA8eSQgmBuzvvnVh0iv/wQiVM9gU
oZomy+DDBff9FbLJ8+XxbIOKmC50+KBY9QzOAbrhXpfNlblmfbn5xEJ5RkG9v1Qc
QI744XDw/qhEjMfyPaRUrgyaJUrY4zHXYH4lxingZ4bsB6M04+CtMLUF6hQkZjj1
xWVDx0e5Y+0IH3/awchf6sRRoo+tB1DNJljjjFLb4KGZgMLLiz02lun4x3rT7znY
l5I11YBVUzrCj+zUUOEH0cL1Ezh+d3KmwnhN7C58qyfpOQaqmq8V9YOdIF98yvbd
jCLGcYpww6AfH2cPviDbX6JhqdxXINE5GdA4jMAj4X2eN3668E2kcdh7/NS9AbI+
pvYWdvt6n8uk8sYU3IirB8m/QL3m6jfl9wtNiAdR6LqS26lyxBjMyVXfq4M1ODaT
MXPGC2NXxODgH7IFxmEu78W0Kw9WNVpOqlT5R2dDJsoQbHQT7g00smDPYMjNSVtd
tPtzh9ZLA9Ji6Wkc+B+huvb39C5DBcykQahXJYWO2JAljRlVMKqgrlkvn9hx0abD
j4BrSp5TVKnfGel6Dsvr16BUjr7/F7kzjm9uuBQM3UvJjmeNUA8qnZ0ko1m4q/F0
NR53WW6ux5qnSFOrrYHlhhnaT0RU8jIYJBCLmRgBbs+22rG4GGo0cHLhrZGzUaKZ
SeDgg/8RK7ICgZQDKhwq+JhwYNHrZN5GYyHbpejW7kFjEWReJR7m9w4RIM5UDI4L
iKdFcjVVCJF+XYtu+aLftkj85yvxtKgVx6d9nrcur4mDhCFqGQ0ctynPBlz7S442
jwhOsSquCnaz19ILF6muxDIz2bZys+UPeYqWJiUZsXtHdLPfUm6M98eQZ61RGWrY
M8UJkEyqPVVMWX0Mm59v4ae/htNCBm6s/sYndlQylzjnJs1gpXLjA6IltA3FTYPe
cGtiMIVgiuwTIZJnYIAt4wjjmgeA7D3wW59l9TF4vm4leFdUtOCvOYy9eiPE0eYZ
Ifx1EXivdB/apH3wipnvmZKmZsbiDshDVG8h70tohwxu0GRlcuQzlWtS+4z4Ja/b
36X3XeNUqS/iKppjchG3NRPcvqWPVeOuZl4YD6a03BDrVMJzurePDQTw9/XbSsKo
cJQYsCHHmFj0xD/4aa9wJJO+xMOSVYguW5+Fac9+thzT2p6HX6Zr2gv6gsK9p6No
KviHN6YUFzgNQhYcS2S2VDPfKxQnQGqyh3l88d7XdJ1UVy1gkR15CRLj6Ub1opHM
5r/Cje8Y8YkH2uEMYlsh2Z3T/xgx+t+KkUaJk0cN+4n9ACmjL7Q2yn1TEWGkPwop
tU/cApnRqfSr8o1CR8vnnm27sQU/xhke8jwNoFkESj3uwBJk88oKile/9wcssO5W
VD6KQixL3g34yMDpb42dPTWRBi5Lp+bYzMZ231eTOV1aOwiUxc2JsMMOF4GaVKUO
VRPjVjPrGIAnEhnh2bq/0Eh927TiipkJtayEPbq2z0MF1+TAw47CFziOwdvFTXDc
PTw06riPyC9mwFdPNl6DUg7KJ50ppSBIEyFMCpISDr7sH+XMzX/6A7ztVXw8hTYL
MaSVMV3uXWeFxOQeo5hgnmybdTR8NFw1l3hmlrDd6Q4KsW8gR+Orv/gN3hDCscmP
GbV6g48Y0RiuA7YPaustecdKo7GCl62CKWN7qwyRVLVCjUaWub8Y1l/dq8bMRsrm
lczrDVRJhWrqrjS2l+oKazF1XnrWLx/CzAOOkj4I2/PRvhbyB/jHiCi5CLgXvw6P
JvzK8CgO0Ry/FUXl7V4wrkZngZYwytSvmKl9eKKr2hS+xhql6NrJfwjDcR8JeEb4
rH36qpRVaEnP2CSnqJA8fnD6bajOtE3UJgAcB7XArjzQMWoa8IKQX2YZoA3hkbz7
kGWYQv63HXyXpzAnui5NHpGQ8GIsH7eeT673vg5itDjqsm7g6NJG/5x3ljzdNPB1
luv9+Pbhcv6ejeGTPR7Y8aDo+mCYO2+ngAMAqzWhg/BIJW01gx5bj3ZyOlredCxP
lVLRrbtnTWHENrjqA4nztPdittf6RA2jKPkTL0jFGClFgy49JEZfVNt9wYxkHVHk
npM6u+Lqo99qzBuA8sjkTN68v2VaIAhMh7c6yCx+pJd20BUBOSPQqLqHbIHfeOl6
kEuTCgGUSbC9GWXI2TwwOs+7TotzzuL9R3HOtRL4AIz4bwNGWj4Yud7i3mpbqnJS
4L4TXhvvm8h5foe2a4pS4gNNWo8VItb6CuhzZHAPsoAwipvmnO1mA9Bui1T0ys/d
WA3sV20OBkiBWRQgE2RkiBEnJbNGr/pMOYMBQ9yBlf0kJORx34qR5i5jKxOQdj3C
JtMN3w5PA+NpRqdHhIMj4CeMaSrdkE5R0LjpjB8CiPiKrBbsP8GfsSaPxTQ0KQWD
D1Rt1828kvVWaUqizkYI0VP675K2i9GOuqet9wGVmbp865cefLjsavpvFe31dJC6
+kDQv6cHp2XZZx/SbyBeOU2VIPzunJtUuID51iwkvrTc4kOyV1yY6b7NkXE2x0St
UUnu6n0vCh2f78rnfgwZ7Ho4/6nLNelzEkQCBrAhk/65CCY2bfVDqxsCZAalm3Oc
gIsFBHw6In3mp8mOdjLKfzF4qyDzFDWEYm32vsf40ZRC2f1QVzn/Ijp4CUBT+IHz
LElKI1jjVlmVRcjVAv9696Gw3RQsqxB93b2v1/K8b2SUPiCQGrlZIz3wevwoJuCa
lbRdpIW5XNHpKpPksO9W5E5URA2oAK+rU6+9nAKtgAowjXm0ibJFEF7SSbkbiud4
U4T0j4LJouVYDu06ZNZW+Q5kT0Pu23oveyDq79iLk5aFAPGQSncRVeogt126pv70
aTYye5MNxnQ7knCFu380dOac6PubtkfNMiYU/Bfb6qQI2LYo8pjFTfrb4ZUOQ2lM
7h2ptjpbaqcOej8SgPLQAubfagBzBqnQkaxO4Fz3aLTaPcEZamSe0/1DvANm4ShZ
t4a2AfvLAw4br9N+PsupVOOoqItqJVniVgi07/npbKf7xYB5ZfGz8ENw4y9p3kuv
/nfuL8qWGP6DhYhJHvSXibU+eCLxs1sHQF4GEf7f/3htn1MaWJjV3ZOPvmg9Opoz
1nXOBzmSgRh0vwH28fkmJnH1PFRFfEjE8u4MdnlyXshIRFCRjPYNjI4UPr8LKACU
zrteDPTIgLn/kvRE5wJ7IHp4R0m/Yjn92bkt1AeGPdHZnzY/4I3/VcVjQZrYYIje
PUy+1iU+mWSk3BqrPcTcuyTcHxXffBINSfXexYZ9tL+837G+NwxPWNFPRfmSLpnV
5r2fgv31j/h9KMS2JqaJtZsmqsNrwy4r/BIZJtad+kVChDBkoZvMFdbSbpyQ1GW9
Lx73RBHt9e0hXOyn43koKohs4w3acWLJl+YTtPnCaDd8zIYsa8i5jAiJ5B5rE/+Z
yz7qWjg5SqzVjjACjExyl780gM/8pzmmi5DQCzQqirnxxFlMVIxJ2Z41lpsz8b+L
R/SX0x74JoPfnqhNc2zHnoz9Hnw8IuP7YxEJ+l/FI09UMn1Tki4oFCI1jg02MGM8
GqeMYhV71lK205V1Ud8V3wFt2q2LCYbWLmPGb5b0QgJFM1mFOnSLtIcxaY7zUNMB
Otm9stDH55DykZHYJ090m1CWSBTjfRml2J4X/ENLlOwbkZyefgFWurWv5dXA97iv
IpaRdWcmM0qR6FIuH6ya9dNAheNri177i3tIEDKXFYMsHUD2Y2FpSasRFN2DA0Kd
ZKI/IdWcCxAAWgjdAXv/QqRimYWKXJkwI3GUZ7JDX6MgXPjLB0sbDlIdHlJiSuOK
TNX/fAl8oAiWSV7Jy3Q2ihxBgRaY1p2jmj3rNvMlcFy2SN/3taqzBPcL0pE4lfpN
6Gsp4apk9srPYpRdxnAhKI9QJapJSuEz1dDk/EP9Dc9+pntTDhUV+c9XpXTrNym6
aDV3+Nq6UP55FbpFhhMGn/g16VzR1FIgGQEN/1/TXPZHd782o8YBOI0puhRUMuAz
AjW8m7ZTq9OGa+Qf1dxYo9fAbDqpAe0uKfjMZ0OVZyZ7fdWB10eepbKm/4ok40AH
nwE6gzTYHYK0QdnF2MPJzI7yLh7NS42X3eq5D0+risjhj4bSTCfiND2WdGxs/qLW
FQXFRHgehOpOJobgZxf9kyc/ODu4RVPkMR8Sca8Cnijqn6UxXIjJv4epeyXyrXkB
4DRglrtveuhbFoixpmzKoZfLz3dSGZDtAp2Q3fk2I38crqwtod5AKPvv5gNOwY+Z
BHXobSJq7KyCCc2J9CwqhVjjzr+ClsPVOEdOu1kcPB3pboO0rIsjQWkuxGxuaZvM
cyeS+zk4DHjhHPuu1GeRwJEwj5RmJQSTgvbSzYTL/aRAfNuVI9xf2iIO80Id4ZGM
vxItu72RLzimik941jrKrbg//NdV+Lg8I55mqaxmfXtFaY+wdYU99S6b7t3zTjII
sRRurHSOvG42np5CbrujBoappYAgQwxPxd3arwrQhCdBXfZdMsEluHP88zDYuq6Z
e7SK3SiRM9pj4WlnTRxdQRMen8i2b1OTdqTxqtzjK9XJs+Mu6Vq1Mv2LrnCtFrJ2
QezOVKG1P8PkCzNSs90rYQuKkE4VdTBKyE0qDaQs5ljiDO2SjJ2qpb9PpBzXKCv0
C6iCmPQjMYPIoqaMHQ4aWZgz0s9xfLmQJFaceTOCnf/W6zo4vfUD298JdnLmf52k
Us5jfHTh27s/yYP5XK//mPrQSkVnFXTg0UOiNtcVDsQ2Hk+iTclUOa9zUEEPmBah
gPkplB+8WHnNBiFVo7k5CmgA0WTCAxcvPgyw1H+2rED5MBgIRXO7VvhP+NMAzJrN
e38cYJMJxItb4E+UP+tkofa3jG69qUwlaHMJuhnQ9bPe/yZwxbZ6jLjHme99H4m7
/dD3ys1Cn6n8rG6MyyIJrVL83to3nOXX0h/asPwkKcgaMD/tVvuM3RpTJatT7DgZ
5s+rqpkioeB1KhOcNk591jVS9u37bhH3evVnQZlDCY43vd5aEd2kkjSY0FBWFSUP
XBKhgLWUujU8NzwjYfJMNzVxzMcOsEYnkeYRhUesTZqv9YnfJi2Ym0EqTl7vDLuk
r8EMR5z/dekuBAoZdFb4UPpbaavMgoG2ph6rMWParScW2dnzXF3vGJ/+Tt1eJuRB
J3WjvbSuH1OM3QwcIq6VeJzKXaPoh9PB2teCFiN/N3BM2q9UkB8dh+C1iQe/3oo9
FRnh27XGJIm4tXwXIzdOPC6HYR4llurru2UsY32iSCT8ZHakglfVpXtN5se2YQB1
bXPds2mFMmtMhKYUN3TRXeqoZhpZxNz716V0RdklKY0D2MI6nWFObUB7y1RzxjJe
tEH+CyYG7WQDCF9fFbMQe0Js2R0j/HkvmmdvAfYZAnChLYfV/fgoSzBwkC8u6Cix
VnQQQEe0+WTuQeRtbL/e+Ga8iCaaXSI0ZyNtiQhpE3mcUb4imh9FXXUB6BzfJlrt
ksfA1R803aDcmBiyqlgCsXtHlI/8sT50fFxxjM4Ox0kW077+sqB68Wm+jN5vNobk
9q1CCF5DvP7d4qmzIL8+0pCCeVEPN/j7GKD8scWO3dTc+799PuCZVsu6CSZFZuud
M/sCmt24esUCwTFnELIg+/UhwnQGJDT2aGmd/UagyjEQjUM2T2DSKtAirBMdWm+D
z8faoEhZMORwgaX1k+VvSnkieBjaGpzROrhHAUx8+TUNRjtthuxJC0SJ7wLXyfDX
0FkbmEzjEnoHbLPrYFZZj1ogA5qMw5iLC89TD/E2A2avU15hKRt7oppe9I13c2Wh
Idp5IMdMnKvoTJQAfDvoyQwWtIrXJ7LaH1fnP3wQA7Er7NoRccAbWgA9uunK+NYM
ZKWlu0Kz/v3vI4kJJPh0r8Bir8X2r2gmRvJf1I6QT3o5CgmQGmoanJbkakmOuTf5
INcAUx2HoL6HpHhhdRx+PorwIfvNAKLe+3KsrcVs+2pTEhFKRLpaTPxTggkZ9T1+
QZ+X/ZPfna//WnRNj1aWggjVIW5AaG427U562LImipNNOJPaHAUMxZMA5MkNeNsI
nzgI8brJXXLK3gkkFVy9F0RNksOBSM9iiUkkLtnxlRUz/8l4BDmqHG905L1FQFvC
1O9m5eNQbuBb6RPFMK1eRliy02kNn9teyztqf4pR9kdC4l8UKIgWmy5s199plEA4
a0f2p7Rg6wCiWSdO80D35nuCfP0HbqoJs5mLvkK/prSAyqPb+Y/u0btR9/qvj7m8
ERVPoR4rtKxWy30MA4INAyCs4zJH2VaW7xtQFqznzqKIcBo5bOrgXM0Z7r+teQPR
4Q/ExyzCd/GNDLx2s2gLrAFGL9XQpDPFtRTmn+04buRwWjhG62Dr5yPGz4vqpmZS
DX7FcxkvGx7a/d5Ec92MlqdAHaWQ7vPTkDlLyu77iDU33be9CjRbL+soiVZr2cgg
wFJhkpQG89ihX7o9RA2AGk3tXgdtWkXmwleqO5P8SDAj7F83C1nXehlS/Ia0O1Do
qLoiM1ZlYxSM1JdOBNwQYB97bS0VJMKFSNyD59Wjb4Uwo113S0H/dAwCglah8IP4
Neqpu0GemLvMBqRTefPbRJ3Qqw5zmINRBVaNfk1NiZ1Twxt5GJad9kDN3bq521ew
/XccO2A7IxfnW+yF32CJcFby0D+zsmqktLKumBgT4xmHa4yAGmjxt8eq/5gsDrGk
rkf5i+5zHZ6Y04roL+dmDAuVaj1Hm6/++BgCUY2Qu6AnTok/rQILxahsDsRRvDEC
DTjKCOpPYAFp8oNsIp5YBbMeiS0JY6iRKfpekgsyI6wHIXdh8j3+2OC0r6FCwFwE
LBydK/2aVUyxYqJufOEDs80YTrnClTgqh0ztDK+NxxdzYG16OB7nmeEVOa/qdTpg
O4pDx6hx64UjUsl2l6Pv5Yc6hJeMQ17/tbPnJV53gsB6xsIoJBUqZjE2oSbXo5mF
OZ59vlx792mwUUYc41a2r+ePd7Jqh0L2yRakFhB3eWR4CLCf05lt8H3FjOEqOy5Q
FeTWCG+t9a3LYmiCQdvTRDcr/I4q9x/s1oJWIc72ost5qIj+5ZXWw1kGmOHXGSBP
+OuTRgiFg09xZRehXiZWS99hKtoZuh9TqZ03i0GTxWFsf05lOO3hOGfLeVzluqKq
YmYZbX7GWJrc+CzI+gFg2LFJNrQHoS2diPZmM+PjI9PCPTvtXfOh/LEFrSAyaS0M
u4XMVgCbfa8yAfOg9zFZgXatnBhudUjj9uE3amh0G2SAP4onZbx81YBZnmp0772m
msZHym8a+9/nYG1ahpOgpYohVcjvVciSzIb3TQIS78LD5Lt1NB6hOYotKoQKHy1P
b+F96z6EUiz9YK9VvEyWEkpHoekNi1+by3hP3V+rKYI6D5Szpf9KAbR0maytXCrp
lZ+UNdfDGP/asuUCtu+zqs/VFhzLIXLvxvifE2Xpoq8wyMwrnzJ+XlfaD0Of3/gX
av+0HYuEHMenQHc7mNQ604ZWHm8IVyaa/y2xHKv/hKhGDodUR6TQFcGmQf97URUT
PVo8rml45o/dHKd46iwyDOfTseZAglgx31IecdvY2T8/QCYw6Y5Pk3dDm8hISBil
Pm48Nby2l0m6v05SXHJ6S+Kw4uz6ISLnmB9GrK9UP9iVBw+/9hxblxiY3f9WcMCh
w3TCnXHGqcjucbKUpoLsqqErNmIHDZ5j3Fs2psSxjro3w52wjkjzcXlWjqrQgdIs
gScSBgBCnQi1iGWa+G/t9YfXv7uwCTaANP8q7uX9hnYdK+uXwP0eaqFbDMfl6PEx
DQiUueAtGAjNFh7cGR30orSOoOgtILIzfRAwp6vhdPHNUtYZCBa2cjQC95w9L4gp
hu35mj/w2FbVGCQFPtkeaXO5gSm6qOiM97rONGcjFOOLEpA9ZW53RLwiFIYMCyri
aCV2Hl6KQzB3sWBZM59t2cZFtyhWDl+J2Cjl66Cmn1Jkb/Z0akSc89MyB9d5TvSE
wjLwnFCiVbST9/MQl+76B8p+6hxt2EfNKCuYYgiOS/m/mccrSuHKdzZkhs7t1E0y
YRIK3NIOzBpcO3MoyB8cDasX4UNpswi0zhy2pJn8WMpmk+HrB2ryIhU71pJnET7A
nI4hRFrokwVGHYwiaWzWFUm0/0TK/Ig2+2HAd4dlnfzLqWYMH9Z1PqJ4REcdlOj2
0eaQe3SUXYep4qzdr4DMZ0PGyKaSlWfW6lnZm+xWMq4/Zc3RKRXOJBO28NmXYiC6
y80pH6hRoNt5OaF3NGEugjY/l0kGeHSO8mmG3CmLBggs6v9YwWFjJFCoF0jXiEG5
FlNC6QVop/DQxeDkD/Kdiqrm54ThLlZWn0v9OXhULmP7To+ibC0LEF/R1Vwq3H+7
m0CF4bE5Mia6ryVMPlQ24EzSnGJVo253JFZJaSz9ti1/Z+T1+ZB2VXDPOw68JC7q
8agLaF3yxpjmpb2xn8WPkr8CGgOcw6oVBVTjYYuqZV1C0i4kTAo86J6PbTS1LeTK
69+9zJBIMatXsDICPclwotne4UvKHy60OgbNSzv4P4LQT34qyNCRLVK3ePOmT6PW
ZpPvPJav4AkqvaKfsVMDtvKYCwBx3BTos4StNvZccLMr+pflB5H4si1UjmU1r8NG
ghe4Dsc603dNW/on7r/CjD7G5QDBr+HJLjZdUoRSwO23mnLgOeoiPpyaFvMfeeRW
IYWNHkqIXufJdU9N0WTRlR2bLFqVK8TOg9y6gcC5ibrZzbrOl20FJcjeKxJ29MTx
1h6jNYYejalWeMXjBkai/mKP1mvl3vupBWR8IlyAqENPThiy0Z/Woxwf0877wl0T
rr3VraKfj4vInti78MgZ5B/6bbJdQEMp3Hb3/eQcGBau3SONZ6wwHDHC1X1pJJ7M
CuU7DSpjB/JB0rqv3WU4Rz0Sx9269vKPVCIE83j7TgKfzb/vSzQkydEuoAkgC4Ep
gsuadHGHo94nEI4UAIj+UgsppRsADFggpPXhoOoJMiDAtiLuLtFuCYrQ7+JaEUaI
Dsb4L/QUWHpbhDeKmH6hfUUdUxnxRbaNlCfo5MD3KIYo5QAWWSCk9z3WwSFEcaLp
wSfr8o4xerW62+ErJLkGFmkFzQBx2gy+AMhlQD0S9PMdvbzggDtNLVW4Stp8qnJ9
1f1ODd0oLiovbUJ7EedwHsOrr1xsc7H3/Y4dZu++3rqjApzLwLUMdaOFF3Z4TLcI
+fjGx3sqigl2BeFOaaplu4YwEeswL/0XbiYXD/QiC8zfpQr7WDIwF0s0ERlgFWcI
4ndlL82g2dRWKq9vKSNvHSKuYahO6cb/+EbGVHmjToUu0A+X0mL82pmrGBSSGQLk
Y1UN/4MYn29cvydaeqIdGRgyyuc7TOP1ESjzsgaLyWTyizi/aUy3gjV+zNSm3cV1
SOEZ5o4mvrERYV0/mUiBgcRUSwdWz1GALSgzKg9YeVvZmE4z7BJQUaqviLZzdgM1
6ZplshtD6vpYp5BYOFVJh2fklDOKksBY76RVXD2MPL8QxK8T9HN7dcXfSk+qbYda
Np3l6Zc12xE1g5mtj/6tt2lyc8y7l0LdkW+wV+TlftxBxCUDJBbUcmSZgYaCeglZ
MEHbi19SQnJEBsdSI4kpY60xSnwonxV3yxtkvL53K57KvZa5lZoT86okQaAt6q6a
FPUJvpBsgDgncmyP6Rgq/8nhyHRbK9rfaZ0s2Ikf6QCogx+Dc1pLI6D/uagi99O/
yYKAIIMbQGLuSTXjcpg73R/SoiLRWobp1jfyroRBBpmy+vwCJBG34KR1zpZyp35d
IWZBoo3S2jLdjIOoGRAcl0t2mncNRTZ+Iu9BoJVv/WVhj03GM3kixUzjQm7qGSL7
M5aZUXePJSI5i5u+log3BK6x4MBhlZ3EAyRhZ9DEpa/QgD5X85DMcPgoqxvfxZm4
HP5thv2AL/wOlIe/+lUC6y03rDQIRY+bQYob7wusrCT+tWN6zvJ9jxwVobS/P1t5
iVLqdbTMd+jjRREyFfwjw9KgIQZOl/36g7lcEIe8Q4v2Zw18f9O5gepKjyBA1ye1
74M89+pyxFexP8RTJ6tWdqtCU3s4gC7tq2lxTSE7ieIHAcNQbJDrI1BUqXRlXyoZ
09OtGz9qs9/nSopTaxufF0pAS8XkIwAthME2FeC8ptaBTqAOu0NtgadikdR0kF5f
o73FCihwCO+a+wPmMDk6Oh+eSpRYert6rRKuyb2a0StujT2Vsir61Hl5GXZX/Pin
0sXuL3D5p/dSHH2r4tYO2CNySgeWZ/SQ3Q6Auk1PEVoinBO9rADxQo8rG/VEkckT
9FUSMSCc8Fk5T54a+7MTPQQNnrLHL8RzOmbRcA3lxeRQS+v083tRJnWbF+CvsuQN
scfVL5J6VXGWc/D0MTgsRPFgy2WuvEdPLnCs1M1nzOQbWEom7ROL+GVSFJrHNrBW
wjZ4zGIlBT7AYJVvhXIBo6mEwWMHgjSCarrZSsJUl3iMg9fDNTqIBPozRCCU6VwX
coPisuSyWKas4J3eW0D3vp56HTHDCRT5S1/IehY0CWDB+45trBjgGGG1+4g/P022
Ir9BdC360rvwp/frEB9I+U2eTsXm6TmhQkW9FMMa5ZqZXGR1DlC4F/YOJDRDsbFc
uskGi+AHjf98JltCUEOq9GT7oCKZGwcSOshDM3tKi03haM42mPvS26NYwgkL+vE0
4OgwXHjOzRudA1Rhutxj15hUsMPqj/3cYEsoGwKnpHbVNISEInrjbDh2jIF1/frR
9JTLgzaKyiKZBceRI7FisStP3p7UCvVqBlBl9VzmKO3+iwEFEEM9xAZQKJHtbFeg
2PAWyksWIabBt1u48RK987hSqMe3kwdWzrCv7XqKb+WcD53jE0YZ7g0tm2h0PH9e
nAC4OkRUdlj84EuJRXYA6nkFK0Rv0WkCMWdcVtiRnnQgTf8b+qR7+x0zXPs3WzPJ
irZh2uLkHNZxCeiZUEishfbUT6n5gh+iKSQM6VEpTsAeNP7B+3WYVR+bn/9jC1L+
PbHZioQRek0ojaQMJHhCzEGjEt89Y3lIjNuko+MIdD1Pb7kPgebcLgKClTbuMI/4
+CJIkqidQeciOgiCBSAjWkH2tKPpuFnOX792A3cT6aAYAf1CqB39WJwZqY/5GcTI
bKxtjaqA5cyx+vXDGunUpTvjOl2bALLRU673N7Y3sS4gCE9DmaimBraaXjPIBm5n
8tDTOdr9aV65o57V2pmO0onHe6RaRuOgznvrhp2an8cDa6aYutU3ZX5nUz4ctqjv
R1XPDEG7LXcFOlLJo7/sJ40ZbHZjTypxfpyDVSfYECLUykVA4A1vxGW1PMtKvrZU
5C+g4TCF3gPUBnYpmB93cQv6rWuV6Qhw1wxuRzvviX7DJHIYfI5sHMs+TQMluoTw
CAJn3PizxVI1AQskwXXZRIGs7bCv6A72P4QSMLtpivt5yYFMPccofsILpIWLyHYa
DPvxRrltPyzB752pkqqi4IgCffDb7gMzXjaYDpaLQTFXOLrNjEWkAAq3D7cT721B
afgBHPZ/KCq5g/GpdVT7NxR41Wv7BQe5cnw00ZnVIRbIcBWiiGLT2zdlw5YaROxS
w00TmEdS0z3hKWtOXheNgcpIqpQzyvPfARyrzy4y/jQkrYy+lWD8vg2PpsPRw7kQ
Bvbdd1UG1oBfvLRfC6veq8N9+tcFeY7fzxvQG2/N1jH33Kcj4p54puznvfNDbML3
9o9PcqgDorCPz01Bvs5CXhK21Fi+h8fMDMf+AibM51/EIGj1uIvfolh8/PrxRRRQ
hbr7RLqmM0zVUqsS6P9kCEB22yrPfnKkDOt1YJS2hWGtjTl/ryzIsTLr9M8TsYgX
ILYPej1XNh3l2hFEH+JqFbbgCg6ODhkQo3Hv/dMU3xFdJurENnZ0JWdDEZfc6azH
EYCRiX+Dd22Y2RqOmfvSsQ4AwR/7n61mFR+0otu75tyw6rdXVPSrPo6c4jMOScPP
WO0gvNtcq1nqJ8YLt28ddc5LdI0keigU58OzhzuZk4ekZcBYpupXAbFQ2vkadhNS
friq4ZCaDfe6F0lkHWmeIKb9p5rZ7bDwC8Y6SWCzMTNeC7QrxXvr9BGUEbV4zFuc
8ZtwhKy9NQAekUkXBb1ewFgX8xDGZyIEGtds07Ah9wEUY5HhJ9fDr4WXA3B9XksO
R75nfSXu/tFKTLBoQO7kozNbW3JBzCBfs8oMVYvrsXq0HiCAdGZRDjifTRfgd1vP
pCaoshJBtuumN0bPSIzp1BbK1Z3yab00jSa0KVFokqKU4+RZqxe/WlZaigW7PKyU
hDfEF+7V3dX1K9LdTBzsNyPiL3hRN+bfV7b+r4t/fTIaiNTje3s/22qVMwKqyBDJ
Dqr5pTjyyK1X2wgT69TNMErdeYh7Ga54bHI0iivwR2E97Q2vax3Jl/YrEk3ZM2cw
bgBpgQsCivYGvsXS46+PHySNbIoGnYDUenI+vdXHWXU+1b7Jgf4iMBpDmyZOL9jm
eTsqnn37Xh8OM00FYYRMIh7C7OM/U6wJejXeFSXszmzj7QIeA3NT9KRcRVOS+JcP
hWi2rFWq/jP2PaIGFLuuaYcIDkn5PPetVZZAtKutoa7Ah2jQ085O9X+hlN7/subI
pz3z1bBI4qlTaQ5ITMlrdyX64Kwurfpwc+D8/rJLzAOPdEnNmg20g3brk43S+MFe
pFH2hSTzvbCJc9IWAQ2tYanSqC/MrWph4pj594TaESdyNyg/5PqrqSmiQHMwY5r0
P+55QUWjVaEQghBVE45SV1XteBAcZa4nrkRXxU2nPiMI0z+j0bHCRgFTw5NZ6oXh
/iBaLA6fhn9uF+a2IDgVmmVmwPYvAE1ZFyhGiu55p9wY0Fb36YgmbcEOBSXcoea4
KjY/rUcx5lVUbxI/l4pzMuziWVBccA1SXFGEoYjTDyA3pRfPaMB6E1uUqctqXtcK
ZChJ52GReeF+5RjN8DCJBqjZoKytg0VaLu8pRvdCQz7JNKXMVa6jy6s8lT63XySS
1n4/vnQDTZ45cFxultyphQGSyqnPOP9fixrdOXBfqqbaWrLzmuwRQwzHuAnbvAut
KXIAzP2VcxHdlHcmWEB/0YTQtFySY1Y9mxbvYrzX56sy1iZmUsP6vqf5mxgbkChf
LVgaWiAtVLIiZDFT5MaobqjXwS4S5TZCf2w7ZVI0J3iLWxKrAs5tKumWmsdvHzaR
PyYaqyVhpRUXbzkXvDzW/w1PyJgL2ksJgupFSbRCi20LY4LgdxzhYLcK68LyGfDi
jYJMBXGZf0yp3XbsN5ZPcDJtS0FFtpmbidWBqJuSyPCf5Z0eyr+3CHum+Bb6Bl3F
yH5qibrrNPgd9pOC+2bj2PUGV8cS8pUiBxs4dbDLrLbAVbLAKoxY5nIvSBp5SEwN
fZpJNJqgeBJl1SO7T7Sr2BHW2jk9PxxFKXxkQJniRA9ctcueSjFuk7qqwmC/4xTh
bKmwqaDyGAP5ZZwzvClX0UHklQuX2fOZ+3NgQlyPlkclhiCbRBsL1It5VTvhIHb0
DVG3IsbUVBGFa4PpzKEyqfXI36sIvIVLETWhP8iqmgyQxQ9R0wAXjnKyL5PYVScr
JfWuup61cIDoZ0N/etT4vaVFyBRrHj26SvUL8RDrej4ipYtfru8TkW6v65ElrN9Y
QVcURh5OkZn2PuPFoA7NtJ6ycj6ufFwlph7TnT621KToY7MOr4t2vC3qKpmeR+jE
v6SzYh54bmIVMGXILwW/M1ObHD50eDAhX2ige70dKBmMWPdS4RZOQIgiApencQTn
8tI8mbMGo8WmtB+qeogj3OOY0AYAmlNu5dLfFCUSVguWh3ufeQoGqOWqb6orR3Hk
rPgv6OAq9/MkPw9IFcTuHerIT1ZcbIrOzpm2spCRvrnug3eMEEevnIPGZbCBNEG8
ShKShUmAJ3tIYnk/lbEebaCeZu4YW/VqJM0vIkO9vIuyoYWa8xwKNOyWDqr4Rtkh
ia16EMyhRgDBfatL3TbfolR1xyAY+ddDSLWDQx6I6tK56XnAbBdPuvqjHYJPIAvc
mSY6NktcAfR9YcPmy9UkmD2VHs1WECDuZN2fpEiNF9AEzKLHhNuwwQUVZDHMbyrP
fEXaFRliVn5BJMv58DqjDP95vQhmEYd7+hzqYBN2pdGwyUHyC5bE2W1WlxEmMYvx
d6YtQmWkUOcTxdnYG/rWa/3B8hoqqRMabZnL734tyjBTOKl5VxKFkDlwnjDPUusM
+4XkeBKYUq/B46c9BU7rQA8xQePI8oPycG21qPju81fu7yJeG29JQyq7wX8qTn8i
ELvt+tt4OVruqojul7Ip/jtwspyw0f1Dl7mBg/q5pHe3Jsm4M2cmfaULWX9G/qQ1
fjB1PEykoh/KBaDNnqQ1pTaxleChDAbiXZsvmqiqpi6waMrij8x3sjyKs17o/evW
h92s2SmgBBkijCIURQPDp9gW8OEDZQQwGbuBNqXw66FasGH11uU9RTRFStCF50Sl
P4KU5rpdgEP9kYHc+HMgCggtv7+cnVMonM2CpMZjNNaUQfs4KqFoifjjhgK5sN45
iCSWcDN9nDLNJSclML9LMgjqDKiLuOHLnfNDucWDyDVcLpLSXB7FpYNXRH6XLo4z
+xW8sEGRtRJZLt9L/yWn6/TsvYo64Wvpd/YWIzFQzzsDZWQpgS6m/3KOpcgZe1eM
YrtxMrG1vgJ1a0lMQ3LXobs6lhGzn/eJEXiooySatVM3SYZHkhyykxKcYxsXoZ57
EsOlFcAl0OFBV4zXqo81d1JHNN5NAUyw7FrT476JnXgnbkjynN8vIF7imkAynA4F
lVGZB+wLF/Hx5zYV5CBboLBUBt6yd7+kcFrkYKCehZf95OGCZdQOUJQk56IGJgXm
K5ui5zCbqdJz3nD8/WiouO8FcYUk+T4Rc8xRUI0aw1M2XB2U87knno51NjEjlnE3
Hwbf6kvlpF4n2sVitWuSuaMlsouyrgBTF5bmZAQKItMLNTHrcYSXq5sOA//fFJdy
ZwmoS7JrvlDdteR2CZo/sBjbMAsIXK+B17Y0sMWmgzQEq2kFOoF2a/m9kmGVKRvT
Aydx5rhtuV2BxCVKPZc8xnp4gynSU9/IAXqO7fNekbp8YGTxOjZqT7vP/QbF4SgE
MbPClC6nKpYJvMHeohumV5nPh3jctGPmfgjmKsWrUrNbLbSV4AV8tFU37HgZoPLz
TbfqaHduZ0yYItnQd0S0hs79sEzH2SOb7Qy0ok8CdWYkBIDx9p4TD56aqGTw+FJt
/4vOedJgRGILB7Zegm0jsJub6e7ZusnRF7IHlQyU0vCQTE6rHI3+ITYFXNgTQyMa
0511ehluMyxpWyVpNa9/clwp+58F0uXyeh4q0sQThlMk4KQAXdWyii/gYylPZ5MS
75fFQTdp4nSKUgNLjMu4U3D+dVuPC2ri0QisqaGU7B/QcsB9SZvhF3GfCn0mVETY
2C9ujUqXE7fktiOhUbsU3WHhC/fK5D3D96QgIilaeKco5G+LqYMQ5hOSviLHZTTd
k79VQ1tihTv/GfQHNOkgPkUVG57Fd6Ib+oaDlSh9eAnFeuqimxK1IyzwvqNoh2RS
ybrrSyIbF1rfR+4KVH8zS3DEn7NAmUkOjX7G3B50mSTXguuilJDz1Jou+VyOupn5
ZzdCsbyAVfblroZS/Rm1NEVtLwzxlTv+Vg2IA0cqfjw5t7fwgYHQvjVdEiU3KlAS
5gtkh/lKqixSkgTvaJ+n21rYbjP5tcuGgOOn2xQ4qgBNiD8q/BcTkYUmJeniJlTr
meiqi9au4w/dwybtHoBqgiFth3tAhSszjkgkhML5ORTc2NNm8nXixUS1A1dG7SZH
g6Dm5/dpQGd7GICLlTQ3LpSwDtYBbjNYtztmM70+bE+vEoagXjQWxchzcrcnosJT
4AdcCDq03R6ENuarmQZr5WqQl0oMs2iTwXHcmqbvr9mvzr3SFoZ814SJBPWmalN9
Nuf/7fdnu3lkmYGHvs/OicndGz4O8bpyRIeECCPmnSMTCbwS2gfpjRsFNACWrDHt
mxYgn/YeSwpdrWOZ2o5Qx+w6q3V3tpAgnNPwdo0n1roNkqq6uo5sCLxu1/s6yb1V
lNag+cAY5+HfC/OZ5FpqQvAPiKVBEEDNjB0ubwRFihZb3bnuuGYqDt6jYEgKD3iR
Yh0MOnpvGzBhZ7yjdiGQx0Sb6TqKISiTwqWKAF8cPyphvOdqfu8lPM/fAi05FUbm
rPTTSrHRQLgWDqQkzipPiXnCBRKgKzYKr/bv08DNIV56J61d3m1NC12G5uBo1T/X
o+0nJ8tAAvsOv5OPNkLLvkyMXKnpwSPPg6DrZApSpdJOUQhBWO4/br/gtjwThQO6
foKJmFU15WqVW50/kr/x4qCVyJBHu37EEmnchXRp5xRflhJEb+ollMa2/UkQVw2d
PpsTsBTaR33woMzx7SljGuBWZNS+4rhbBOCaNTuuVDpsOpUp8Fz+mb3BWfzxgX/1
3y4kLXO6QflZTSLtALq2eHk6Dgnjz0/jfEKFqL+2pCbhJG4mB3DdqXunRXA6S/MY
s6ZSFCw5nDV7sSB1sJqMqRHPN2lGYRqXKqcGH4iuQQAMnZtxLOyZsiGzDdBol0BY
EMmFTp8hnN4jrzcBw39I8KQw6I/lAj2/E+tbXQvZlV37vx1qeEln+GWPHivCdelY
mDbvZW53hFVDK3hTLB1tDZs49oVT/TmLDXYyZ+iRzRxEdBIibHE3qUrJKn9iyEio
QYvENvYZx0CVKY3ZJ3LrXaxgjsjxdrgKqNWphPL/z/ovPG8k8aLRokm/kbq/2YSV
Q9saaI/3S6DtR4ZKcdCgcRwEzVEibZkDDHQV0HpYcM84KTNc5zqM57F5X5qj+sgg
I+5ZppJNJ6Y8IgL5Si7mH3k6Za4ugHZlzaB7v8ajl2tARce/ecWh9sLvWTf3sfFC
89ALpIyRUg4dkMzHyfyjqrpjjHANRyLPTb/XzcrPSbCbK9fZBVdZmUoQApGe+QFt
/z8JQCUBiNQ2w43xFygBse7xapA/lHfNj8hUP4+TkKtDecNaJeEazGZ2Qu1lSA5u
XT9nk67++PUGqjdL2icKVeOYjf68/D4LqXxelPlnrl+Qrqe11opXf1MIoUhDvkD6
/NmLCncTynt0zaVZ33PoenmHpdHALjRzgNj2mMO7kQzHk3q59i7sdsT+AGeCk7jy
k8WhH1+h1mw4CZOR+STvelBNAKPy339Bqyc+m4MjfhCCqnp/he1FceBEK0bf3eeP
Y2bf2c6MZG8eJeQLpVrwE8zjkph0RcSVMumLWV3j8Rr6b03CSHdHfCoCGsN/7acs
U/ABxUGU2qXBQqohK+g7WHoMguSNHdI7xCU84usetytpaGrOSvAMF6//4oyqCTIl
syU32IPwB9HQKZXWLYVn/c8IcB74G5HtR2497ZK5mmyzC9sPRQvr06GsZMRvG8V6
LuPaIe6wOcHUQAPcipPb3P6M7e5xFtx0LOO1eaRWoaWOrnvfjQJ1Qd/numhx1ftC
DZYgvRimtTZE+bw6apldXsX1c6zzjL3WYWW0YHQL330D22U4nEPDgyw8TAr/gkWp
zsFC8xt+AMXlWyIBmBNfDR92kViId1wnI2oeSoI9AFnvUilalmIVwWtZLrdYf9qx
aOJeRLxUoFjtIOTWjIlG3ZJ8nzwyLyZLdEPBHD78r0bIo7H7Llz1/FBUv0ys6dBh
++u2AzBgP4N4+ICqu7PAkQKs9e37gc4L5jyPtaZdJPsyJajIRiQ1K0/zzheAP9SB
4z7TxpISdcQEnJRsSHnpCrmKyODtJxDUPcHwZf2Tr7p0S7/8xGaGWCn6QXgYOSKT
58WhsLCnek5NpkPDtBo8hJT0SW4t1yfIrCyAafhDFE8RMH1IE1BB+/Ly5kYjY89z
/7bkkcUF7PPsxiCH32KSxmlVC9xlc5XPY4Ez/V8M9d8lKDVBcQMLsvbSgBOJVaXB
0q27b8mN6BixymeQW4SbfFBsfxwtJ9KxtFeNfi+HSD8XCdyYvlCVwgbqfnkoJd4B
qGOeWK6t6gDD2zsi42IQZcq2Xzqhzr5Su2EBz7BKBa53nByFVSeeGYSsMTAi27yx
+4rxJSJD1p2OwxOOOKUR2fcWMy/CDvpTsBMwIOcDWSoooYb1WUJrSyhaNmNJq/zr
B2q6x90VadUcx05FUMcqyAzU2ZwobDQZpkAlu6fh3oYjaUsVdsoooZtI1uOzs4Gv
BziP2LdkQUfCR9IgSxwFmWbfqMmvpvwUPJ5MCU2X9S05AEonXf8F8lgQK/VDC8/d
MPVTEFgfGfV8xHs4eJwhCFV9jlqdJcf4Qr1S8x+sDCIpLpNwWoW4Pu4hv4FKA7N3
THXDoI9clbNGk50ijheP7wgAndalA/pQhnJOwaOfESs2Grshly/bZz7oclazIaCt
dzwXDt35/CHG3ApB2deNNuZL0Fyc2PExoCRUaJDBNmyNWIVPdMzcFsQsHER39KFe
AMPnmOk+7/H23Li/7fi58cHMizHazSeOnJC37Uz8yxCRurEP93MiD7fqVUd2I9wL
ADXbS/gBBpIH6zDZ8EU6Nb0LTCItXdRNu31dVHHZULmcjKBXjjn3GxsJcrj0Bvlr
QJbWtpEPl9HvQ5H3hCIBAjBdBWHUWMewsn8kxowzQdsDjrpcOM95EqjY89mms2Aa
Mb0QmGE/DBS5yzeGdW11YX/ZZ+RCU33kW+4Ppev72UnZ6wVhtbcXGKYMjADo0Uy6
c6P7PqH9pE80wPKVQdBVIf9yl9Ks8auTX8FN74PYad1sLPxPsGIZkNTpiMXyoabb
4ATrKfk4XXBniWqdjLaSID7dxe+VfXxzfPUDz8y3BktTnefZ+FMwUrsdMA3wFXLq
8+5JH/V+UlRZIBEt28EL0XTW+z6GJ+XzM5D4FRZ/Oxo3PGGD6K65rOQ1FDidKVH4
1c/MUuQb4w6/wUw/DA9934wAL8jYSGBYAM+jNN7q2zZ3pgWRtvNjKfDEIw6r4p9L
/IaTo0KU38+DefFSRVjmtcaNLnpM2EqpNbbfvtxbkGkJdFmLRNoxKY0lOWJzNZ91
n2QuYSJNetl8KXgIWDatMZ45XbtBI4WVl1XXSuFC6AeJp6FFFTFCUbcCcA80L/Jx
yNCQK7/vEYn6uSZZP68bc0af+/RqIgX2huafeA44tNLrsSWleALOeglSkaQy2IkE
l7B/1JycqLHf2/96zxLzY+PJ9/D3bXCg6BjXa8vnVETo00CffdsqeI/Z/hptlYIU
9Fos9oMszdrNhHCCYOq1kNGaPYKYHgjEY4eSir+7ikvMmF7ua9GRQ386zO9Da9/7
Zz/MXhhmEsWkv/dswn7E/F0akR9S7l+8cUDc2U8afZooJncc0q1tg72ntRBpbLH0
f9bhjt3uK+kKe9gww9o5wUimikKSRrh+5zrlOlFsoSCDWsfHe2Ri7eSN0zP35jg0
muUYvfcd9rxdffiIwvbc/iIq7g04Nd/yxjTrYKGAhpX1soD3rSPlY+udmkKq2w7B
jwOVUiYKojpftIhj9p7SexcfHscolMHbapVFJBMxnXOBlJjZ8JOiI3Cb/2gjZwjo
M/36HZq5o0fipLlT5VyTzPaszCixBQwkOhtrlAoLNQuaH+x/I7xoPcyNZByCaDK6
v/0icI64u7rPG3bkDTwC8aFcPSDYlXQLLioieV9z1iSe75vO1QgXkt0oEFdxo8BJ
R8tyJWp81h0zSpyct1WsJz4vOL3ZZxzwNSuA9H0xe6j4yMW6wNK87eD4VsnIOq28
5XXqKq1CrpzZ6mqtCD55ont/g8QwqvIhJEVic2dxQgeisiakjkXBVakgdw7nuQY3
si0ZvQeuLZ9otY6jgMFw9zuRLhYfozmI6JhUWFf+ATPowLFl8ROFSZVm9KOU3b1h
/WaJ1DfCajXPySx2/VQI6ZKxph0EWOJzxLSmGvtE6Kpjk5wEr9pjaTJXm4YhLApn
6lchdF5b0xUovDPAXDaOFalv/JxpRK1hyYG9a9Fg6WX7rM60eP8ns6+KSt2wCehK
0ggW+Z4q5bnMkoLebu/Pa2NvA5v5jhincabi9ZxjebC/bWvPuxzyNY29xmcTyTQn
SMxbfxxwgGNwwfiTSUmrHZqkVWqJ2S/7BQ1kyto+rpMdxR1wZftGdCFVdYIRa//E
jRNlWpPByVyWP/9iPP3NsMSHItvUVaeV+lRBI0Rb2S70U0MqxUDbsMCroRZD7DNQ
FYR4/DcNODo/XODbgf4vpNks48huhtwSILWUiUPtrHmdn8iSHJlqAVFIw95XvITL
7sb159OSwFNev/LTMJMC1sPd2wtEO/KjQJh7jMB8I3UDPE8PkVRiHLDvgjlukjqG
h6/RziwvER3moYJMsSmm9LjcSw4jixzBklo8Juogpj5VOoFgbzq61ggiHc/bKljD
jUdT8MNXqvmz4ExMS8rzXBfTCh2Y/y9BuANJOya1n/HlJBR+fOPJDb8juEXclS3t
ZTwp0G+uUvK6sVEd8JD0ThElrC+pMwXZPCfjmGQxD3riwAmCyl8zpNgPY8UjPM2A
2zGNIbtVE85EmMRNlgIk65uADJnchvjnngpo4h2wpGoJkjdM+6Sd2OQUrCJZhKbo
GckW3drLlUO0VPEqnH8NEGA+QTVMGnFJD6Fq9kpc/QWhoTTRV8g8XaCo8UkQ4Zqv
k/iqHJF6v5P7qT/5xHaQHYw9KcKLYryNdBr3517uUOhcVomvIt9LV1lj2+Ilo2/g
tyHgO5e0TtXqtvbyq1VKAKJhP/0Sbhaavd8J8N13/iSJeBCvqTa1AnkwzAKYIS0R
x62bmFaKHNfrbOGfUfFqKFrYzXSdy9CF3KKd2a3VEs/qLxJKrvT1INYewrRHWJxp
0bwUeKd6KBOFxLpwrDhB2qKsurqSLXrm21FUDwYWeYs5lGaLJfYumIzbXNulEGlg
K9wnUl/n0dFs/IbmrWq1UZT4O0Ic/8yma2YJ8Eueeryb4yVCpQXcKCmC9vTCasVG
X3rxgtQywEJfGxPTz5TvxWGkpAUEeyR671UF/pwKeefQpBl1jhYkEgf/vMX7UvrR
Tjna/hErICrfK3GbkCP7nuixeVX7CrlmhoyxLXlLRHPuof/tHcS0JGSQJ1xKt2cp
ph4Xey6k5tU08S2YxQB6yPVyvWQ6stzckMa3jH+hpkFgf0tx16if2+zNCExQbWzq
SYJPlbga7gE62JdY3BCUQxPrHOcE3ZRkG0CCc8yTrvkQAtmbAF1BuAXC6xV/1MsL
BksVWPaTNytNNoUe95+5z3AAzWI6+r1MUh0tmILkh9RjMBuR2PMK2rnen9c/VnEM
1mPD7m11s5JePu9taEGlpLhaP3ePdwoLXGmmjvFh6xtfA5KryOSBpLcPwzJ4sK4W
DgLZFm3lfDw/zTJrdHTUTu3N6PNqs9OF2Gaj+1OJ55JMB8QUT2t1yYJ5RMijU3RA
hW8Ierm+Z4OHKORSwBKa9u3n4Wmz5M97zVxzND4o7W1rQua8jn3j+cp9S31vjz8S
taZlMn6xn685C+Yx8remQrCjAdnfbgOX0Kow1CFpI+QiEgTw11NqSgQF0SGR4khT
z1LZjnrYcFqcwQTQj9IjwEvXhG0XZ9Rpo9waOoAa0TV149lAbgviIp/t7ihSZIBc
zLUBBMEYepiqMe79WSuBp264/qgKiq5ySzxCabqcPNwhJQCwJFDkhUXL+9LHWUVy
3hN2uxLv21yzgWoFR6dQhpJPIxUkz/54u+4S6YchQceUubsbEfN5t0s5t75cdAuF
I2QvctgKFe99g2UMnRs7m+HPnoxIiImvF6uvRyRKZ3B/UrgaZyHhHrqyy1zIDJzg
ptP64b+B82+GRF6DJEQFwhfAYXU593SvNFZOf82tl1VIkvwoFDax0dstnJw5dVx8
5gApGkSBtYZK9vGJXOR88IVryS8GexHxNVpj5peDiHdJgQwdeq3xxPrQ9/9CR4oc
x9MChEpJPB2RPFDdpEBjINVn+YQoS0YyBa5nAcPD5OFryFZDa/PgvLCNGKRWjr43
xBsaReCpoxGc593N/QUd4Jivp/n/VXGGug7iPrtui382w6BlbjIZBEZVKFf8shkl
9YQ4RTe0/8wGwamIMWm/CpP52Ul8giE0c+SS2/lCmJqAiBqZTgSxcmJsE3ZQqdF4
5ugFqQ4xOQgvoQAdrl+qW24bbZPI8lWR+o9325iAeMhTouRI0aTsJvapyWS5EqGZ
mLysWwKU6fT0JE5ihYYrbU3aZZgygqeoYNrcXnaVLkeCjvTTYXSbtlCy6Ydp9AIL
NgZNLTkosPXUuASlhwFEViHsVZFWuAvWgpwFI9dg763CBgQw2O2Szl2kV0iWeLh4
KUjWqI8P0bTNNx5OSfmXp6hnwdQpRCh1A5LWdYPc7wh0NfGRORV1gxcJXVJf5d20
DeMHiSF//ANqAqAixPYt+ybqIsRUEK6AUT0YvelsnJtdRkPP5HiWuiw1pOUHf782
vUGvGMGUp8eOO2KDgRIRJD5I8XCqZ/2LGG9lj+mD13LHhJDINon9FP1pN5Q7QcNa
8UTj8u9Gh6BiqpSXxl6qrj2zUXrX15DBKTj/Yv1FrTHVwu88dOx8L2H3zyb6FYbc
c0zUSk3QccjmHO5Db0QmMbfWXNpjd52AwOl6wuxavB3+B3o+v3MBaJM/o0b46ebi
lwjf0z9vkFiTfT9edbLWVPmL9yId61qfa78P7cBDUKl6nmtn1FAVhrsBUE7BIgIl
q30dZVlZVe3r6TbN7ZpqDq6RmgO6E3aILwZG6qW+z7FUaQF5OxIoopcwdku1TLLM
tE1iY8x0hpINUQhmtkUUBjoveV2C8dRzkcLtRSa3+v/if/zxgF6XTud08YMUaqPB
QfGPZYLUTQnsBnSscXtS7Kjm19xNz4vouaTc8aXgY2Yh58YjVsoUeJrRrSLPt6A6
nS3HOBR4zCn1HCm9U/BP3Pty9ngqzkAsbTDFckKgJn2rO/UuSNYnOqTfOAjPRw2c
Nrp9edC9F9yuGN6kJPffBVp/Xndjczbrw6sCUSw0AMxKuPXwhUva93DCfqBAykT/
lrIiJ7MSF7zzA9YeLaCo6a0FqYZb5dHresApUT/2R/S6wAPQSKxFxlqjLBpPBfH6
wfv/BhkmUX6ciQHTt2yIAv4hMg5q+EDfsG55l4Vp3OLjCwmoKH0/E9MTBzANk+Xt
ivAmD9y96toGfJs0rD/2hRPViD0jW859dQyntI0+RjHaxRgneFRNOiJYwCnGkhSJ
wUcfNvohOxbfPrZlSsAJQME/sh4bgWtvUs5WYfEuClfSBMr2y9gg7I69KUC8SE6N
CLTTQV5G+56YgrUhHEKzehw3KAm6T/ei3uS0+rV3a75f6BDxyf15ch5f92RQP4e/
cbbcJvT9Mht4auzzj3oaog4bXjVA3ppaGwZtXPhSNg3BTifDH1Bkq83F5+/DmCaj
QhzSAgXvmXsl/WUUaERVH9a6PjXYW3195o9ztb47SywBA4AzxtvB+TuPKsnnz6A+
tKCoZhbIXkaZMDMNqm+m03afLNQgyYYZ+pTKbOx6beyYpnTfclrLJzhgUsRaUoF/
7Pg30+oOE4O1tCF7guDaH1rWpcsRtX5J+TFPRG71tANRy6ui2icRBueFqNxpN7S8
rLNtvenaZO0m4Uv4U0t6s9ADKo5XaT8iUrTGsAGJfXaK095QXd7MixgeR5mnu1yJ
kbzilkurJooJiprM5CICWWPr3BhanyEXiEDQGF2AKQsntsWBLy3tAnA39kglO/2r
sLzqgOOQWmYMMkT/+qP7kVmnTnkINN0c3Om01/fq8kuRYJolYeTbfkQVEhUb68mu
7a6qcxRCLZeqwcnBvs6Y6aHp9oRNkgdg3fn+u7coe9Tpo33tpT8decTDpiB+VoRA
6dVW/ScS7fUQp0IVXvJYOcOE/MNar8bUwj1/NUFwlghIPc/DmajpVJxXS4FJxNte
vZyysBb+pdyRY/Tk+uyvx+LgirIeXt0MINMaKKDSyd99UzV4U+FMdpgRMAmBykQi
z/m8rrF4mZ7CnVCQPyg0KSvr0WEx1/SQRrF56RQRtZL+NqiemdIIV9pNbiFp8keR
4r1kqWyOpgEfQDQTgnECe4IIpKiT4J/6fcSc1YDHFPVEJqxnsRBIFArvMKISg7Ph
b+H4rONPxeBRqbftpuRziei6+j0cDML5swht5Ps8rGM3uyNIUkdovbmuvEcbmsiv
13vxtMf++vG2Oyb7KgFM29a5EukznH4hngZ5BxV6zaRN1dNrwQOhCrVTtpHrjUjv
2/v+wo9YUNi1Mm21u/DMvI8M8v43VRVUywVrg0rODz7Z7v8QHiELywlT7rB8fZa9
Cl8FS6ds+Jwa5kWoBGIaghQefWYaMqxu657mk/dxwKHE5k0qPQQh5lXVp4dbTPIM
AANJrw47RR4kBKsK6WE3S3mppVcHTIqlD7mueMXFtSaxifojgO/GPIrtxsshJLwk
7Mru5nsavNMXe21Qa4TeQd3lX5ES0POHSdHYm2ogCskw+rIdKGRfd//ur5VyhUe7
p1OAaooPlinvvK1SSoioAOqUJKow1L+YKjN6acmo6xVR8jMA+Ki65ADKw8//qNis
PAuW7GuomRYrXHHN7KkYdNvek7D+4S8r8+LSiaLSCQVg8JzARQtJzPfLhxsnkNIf
GNCM3To8FXFbv9TyNu0+i9r6qRse7bHROhYJzWflA9HDR0UoCpA3T15jpv76nO/m
JrJEkXClFIBX4JuqOtXyDZwALQn36alKrHwnqvlu2O9cpgJUu5hHUsDSB7llHwt3
TknJO8XG+dMCT8fCPkGRy/5FiTt2uQjwHo/HZwZkpNfruG3dKVodYdHBjR8BVIPM
y/EzZb3KYRmvI2N8T0yJKhoKNBTVEISzSvqqWoPD67vY2zy0P3GPV+C5ElMb5CXu
2yrq9Nl9iWyQ/yTmAT2nR9LyPz8fZ+L16tlqV8J22X4viYBNd4pHVRMjjDPT0pUd
aAdFP16dlQoNVGacFGX0JhcKs9sLnr+20kxcozED2uCi7rqe1V0Z4JHevrxwC0Cg
a9wGtjVCZ7iCnzKzoJNXVAUzojvvbWiXcKxufWTgh0DJDQa019tajaMhAWMr0w0l
hgjACAqKyBZ5Rq9GWWDb3yrnkyI2mpt3LMFEyn6/Fn2PYjdPT0RCymgiT4a+v/yL
xjwDKj+1HfncRwfPed3rlzNMyM+zZ0jzkcbwppO52QB6nrLSpaFsHDFcmtprwZmb
Zve+g5r1jXTWp672jAASU3yj/DbPC6dTPqdht7idYSBMon0EMuYMtob2rs1g+VI6
h7vYw3S+cJaHxGRCkRezn2bdXuYxXEH8d9Vr2M/MaTJDXiCkwfg03aW4Moa47tTv
2f9r+DBWI5E5KiRyhp14H4lUZOnZqGk+GgT27W7YLeQKq+qxaf5P+UHxJQs+056Y
2J5R/6ALFz0kBK6X7eTCXwXQcs/5JMprVZffIebYw7wKOwMvR+s3dv65i5MkYays
W5yesHZrG6K+YHvKjVNYrWiVw+Uykiq/WPHCr2NSq4BwurCndOXZk6ehVM+U5pGN
oohF2N+03IFzr9xsEyB7SaGU3NnFTU4w5PogYBFJhSGu7ZCc9XLZdkzHX3c53foY
42HKxL0WtO2hy7O7zNZqGMQfQET6PwVlxtSvtBoTUah/3+0TCFHgxZZb/IJX5bEg
iCCkcT4nu4SKjpJChyAytMNmwa8w98lx6KRA8W13wH9xenBg+VATw6jANluCZMP4
ueODc1RJ1UPcU4Xkc3qJiFZfmSlB2YQlaPs6tW7wIE+Q165xyd/C3b4prYYOJwRa
CoZTJjOIcbJqNtp/sYFlxxgZW4g9ORAvUQ969g8V1DzSDeMm93MnMKd+YhssKXFO
PgfDA4CTkq48QtCovnf1fWaanTeNUsvdEY0mWf0epTvZcGD5/JXPrrRk1aeA/305
Iv5HeMhyWM4wCOp9ObLv7u5oYfID9Tjgt0/bcyakRXRhqfGPgp/VW8zJcT4uzPTU
qf4Q+DDw+Cvdv8seUvljwYxEbJLOyrJ52dSQa9O9OnqkCPvGICLUOlsJWioYG6Yz
roN5zftSnBisDihEVyoOWhbCfw8+isgYzsk1mlcIB2Ovc9lzBaCURQtobyFCvTqA
vKKjzRaLZ4y15vh18ARIS89eYUDS9kjhyfqPkiZRbN/dVcUqLpTFOH8UwU4sHhok
WJeMjgJ9HaCJo8kymKntNKv4rJb08sbUBccO6TmW3YXeJor6iDvhxytUcccGYu3d
61bxwGlMLdRdUIgm3x1k3vIsZvSzf8VQqMWrktjBSPkLt3sHkcOaPZTI4VsMXLuL
9oOllfg32vPGZLJ2vDIpsxLXIzYKdAW4DKZP6D/CGI/B4AT4E52hRkXGRw0KTmu4
AvfTvhg5908EZfrw16YH67s5edT8kJluVzi5AHfR0yiqH5OS+CMh8XxlD/9LxJZ8
ny4xuUWRPBDcNk6UWi5oegiDJecjt6O5B4630Zg4Bcl10fpkJ1naP7b8o0FrFcCX
UbcvIpc0iQfMEQsYyIyrh3Dolr+RBx/sDB6Q/rKSWSw7WZxGDEl7ONXAMG9Th6N+
S1uerTj/8VQUiJKsCz0HOKXE0/DHCI+x8dq2Qd4PJEZ5uWSkRGrGXyyGgrCOE456
AoZcAe7arLlDxEDjs1tAXYWT7PvmuXa0318tN/WbIdpPSFgrtVNvhOQzUyb5Z2lu
2CX7erTLhPrYGXlwKUx+ahKPlh4xWQZNDBKIb6fSkLcsAZpoFWBvgDF9dUZ6VqmX
XZ00U5Rv5AeKvHKFLqdy6um13oxZGP6S9Ch0KCJEufPldTnnAaKpNh0m7LqFY9Ul
GgYPf0QYVQQ3enjy7bOob6TedrQWOM8lFBHzgLHX3UMK1XTIdC+fO7jxritZSHW0
PwiOy+zkmJtWYyEpN/KSsdn/wEkarCfGk7U3r2hmrBA7U8FmTXumBbacn1KrBs++
nFSXjW90WZj2s1u+DJBlj1pIWl/6OstYxNXckwbeauL4qRlADMTiJS66hgePne0O
R2kCRMBxvIriSf6tNziTRN7YKdQVAleHy/YvRF5/97BbvDLxKrysePPluqHdydEp
P3coloEZmCjCelDLNHYxtpwmF/LX9ZJqsdFdoK40YR7bFMCE0d29ZXDrO2GJlGaW
IcMGTODc9+bCEE1esxhdiOtg6T/1/nIxw4048yoi0GBp9CkyeOJi2N84xtQw0SpO
145B7dYV2KCYqRkLfxoze+3rgfgRU337Sz3zvODAGrvxHKUqyviJX0Jyhb1ereph
spw3p4i+xYDLVNxGGUhtrghI6Eqbn1VnBiCN46ugSEDrJ+xV1J51CDq86MAy/hoa
PkY0FyELoFcouyGOrXsaRDYOcZloD5LdMGPb/ItUyd/OBjDNhmrGalyMsMGJ7R7v
c+aMjq7vb0yPQ7WnAHTO0kb3EFMqml6clwNgspbsRDi7++sbvTZhybPQgzhaZkDW
X6xphnqIipVI186rtlLtdpsDDIm52Awu/uK47Y6cTjPiQ/xgBwJ4tuvpxi8Wi4RH
FqKkIFxR0H87EZAvSQzvlBIEIpu8OBYDLYCIfhmclgwiZOGFX0GkN3Ni6wvET+e2
bfYi0QzD/yY1sFMn12wVwg4xytr9EjKQm1xIHU5wjF/eEER8fWFTcV76zR3WNzno
+uZJ8sGqn+oMUsTUDhMK9DGCnoA/fKbCiVO4zQPxSQK0qXQC9b7bYp3gJmQ3eEDW
J7dYjsKEAwd461vDNcUfnBo2ajeBN5/M+/AM1Te0zpfM/yFeChY0iPVjsXg/BOvb
yxkc7RdUQXMv8V541j5zgJhvHMOoAkrFFLXVbTlT0uc14zZhQLbrNcSUJrTePxqB
KboGv6FYJvO397qwCZSCkCM4RWNq8IhPI5yWSGPkUs+s5KiXdzqBQaL5zhQ1ZaRH
W3HOUvnugmSES+lO3txBSW3Rs7BDJim+B49MBqjGvJaXXejmns0/bWYKAJ7uAraV
6mYpYJEITE89ckdLzlIPcVQRFiIRiNlWrJPJlz8KPR4sOzN4LXkictfIcotHd1NW
Bd221s/N6zsqNc3OmpcR/EP2zqUa9xj44kDL8Ug8Olj3nqkgggz5ANTT/qe7q5iU
iMdklWTGB+lq6mGEsivxEA8v8yDLlcuD1NikcSwBMooqqjEx5vavTrMFRMrFTN4+
Gs3xrlo9yS2xUInKh6SKZyYGmbJ4NKxQRUTL1oe9wJpfRbCuVZp770pILpDs8/TP
5rfMYZl/hfXqQIWpPooljVQaIfK9y/467eE6e4mM1DeLOKZCdjOomIWQJdSjdL1A
VQdb1eQpFOfF79rDNmLKi6tUPa54UMi7xsjr8DfWbRtCcFo0Iy5sB+ids3Vg0ZIG
DoaJc5UHNxRSPo4I870iPKQwZbzgCrDxjG/5iTpEiGHr8mk/XK4BskjQkNGC1vHB
WbE0ilUU4JP33nvW1VfHvgPnJGW+BJGHoy2hZgPCX24BAKB65lHseqd+F5juppAp
8WBC4js/tZdrM9M66kHhO4mxZ/PoEVKF0Jvh3PoH7Nq2C86f3nxgeLSvwahTAcrz
CEH9omVBKAXvWiJ0QUK+rvkMzvkH0kd/HpCyDLzgFU+G0Zgu1bqjVgS0wFxqid1k
eylN7LEYAbJGH8u0aG4BL3XCi2Fu5diKGtuxua0R7rnh6UrkLBba+40MVGYAxyVA
VX0vlB4OxBiiaD52/2a/y1RzE8++euuCBSl2zmqAGmTpK5cgm6Jhsb8YA6ChGCW5
lmZ4blbafOp1ztvlYddZi0VoJBQQLBDpEAPCpRPmvTwRfCOhEKXMjxsV9TDRNmH/
FdZiYIPyYDw5hX4TGP40zXS7e0GYjn6ENPqnrGmHK0rtwoylxgGnTuKAXrG+VeGk
5gAqKCzHp2gQPLW0sy4hXzl+FlwQ66vq5oLkT5IvgDo6+dHTqS7jzbAE0UaObkkj
BueXeJdHWKWrjxr8bXxssmx7usEXVNX9EeuotCPQDqT3lwvMsY6hrjibWLJK3Hbn
A8sf9zBojjCnos7WUouECOqLfPAmTea4NiyBC6XUgLA5mB1wxuySRTXKe8e3zvyZ
A4I6Ow1KEoAP0SqUl8p5slbnDpcxEbEeJBLbOKor+1U3rw/Hspr+q97v5IYcPIyA
kkYCDmpKAcMuwLF1sroy+Wa0RsdfL5RwGc3DbWsRfFtqIBdaIdFK84OQqhcYUF07
kOmfwqyEKgyO3RkCB1lSDcdyQ8whBJ2w4SzZHltYvypg8kynTtt3m1/mBO0XvxYJ
s6MHnysEYsjnGgyONeIKO2l32YXOTWK8MQyxHcM+TIH9F4HbutkoIEW72MRg7yvl
QGdv+D7aztp0UlDJ/g9Bykpf+vPiX6ntY0UGNkfpTTqwNbDl78kaLe5+h131X04/
bndg0KwEEEpjymC6tdxZo5hrtyQ1iR3eLxrEVGMHOCFHenZDznpIQtflttjS4V1L
JA0QED1JhrMXUgSu124SgjVyFlNqKZXEt41kpO+nj/NWjDo/iIqbQnL0N2CpWNG2
2MSWuhIx+F+iPFVFroASmcXAr5mXWUwmm/xeo2kVjYy3MUhzmQq8U9ykLlSc0eLw
7/DsrUxPUzEIURYm8pgGeU3XvCCDA2ss5JlTkubKA68Uwc6agiuBz3IhO8UXqcaX
ll/NxmctmCL2ZTBS1MgN21TuxPxTDcbGAx+FTv2PJjh20fgKQtEOymiIjofJmwrs
6Ot1SJ1Nq4Csaks6A/rkRlVXhP7Ky/pFt7G06S9ib0pmCuT/hBeJZ9RFefccB1EG
B18Mc2VsES6vKo9GDY8FhtL1upeM/jASi2+9FVkhDoby5tpOgNg7QpgOVz41eklW
P4Wqd9u3hLZvDqNYXkSK9GyRZsku+jT10tE0l0NBBRXkXm6Z/WStCflfXKBOxWAo
X8jEXc1hIRedzmI9obYLHJ5Z/XCwfW7xbfmGuYCm3iT8ScycZDPwjOF6sWdr8WBt
v9T0p/7X4z/e7pdLm0ZGIXScU3PnEZiBYj/o8BVZRrI+D3XPOKwkgWAOfgCV7dgv
hOWk/MDiGmG7fhYp9tKbPlvkBx+8UzuxOSQio+H5Tg2Gi+O1lE1pIHWSTU9xP+hA
dpaUOc/Q+x9Dbyk1doLqk6SPKms5YBg/7pY7FV54J9g+o87iSeUiKfBWYJcYDfBx
LcU0oilFW6Ct4mZAtsK4/FMs+emd0kF28g4fRKhZkLHfM7PIKsiQlff3d4AJdRSN
3zbha8VIjVyhBV9Zh7q9dg9n9K0O/fSAOFtIm3wE8kvLMKFnKGKubl2h9mdjAdXP
lhfAhRV8zwlHJZyrEdNflLONsN3BjIGfkwX6zMAjixZobfgOg8e2cDWq2BsHgRRp
X6Iiqm7vOWecjRmUrB/nOPrHOLM/0LHPlWKGQlZQ2xSCPWYg5asiuGnz7PLBW4iN
HOmn1RPKf3TZ+3jg8N+FqN8uw+d+QFWCFBGkd8/qVDUMH708RAM/5UUvyTbPVyZv
1SQL+fd5rrZ7bLkN17M125JxKjd29SrNCyK4Uf27uEjdHKL0frJXWSUVwQZPiL8z
cur+BMBbFJnT/+hHS4ThoYzf8nIIJiJ81nM6JsdodK/Vdv53q/ISx2Guig16JOW3
v9U5UWGP6d/MMGeWCeWFn9m07OtQDOGAyA9pQ87ycplnYU23qsdG4idt3CzPJgpE
OIZ6uyaboR2R3fhLQk/xSo49cDBWBb9Y4HDOY8CeRdYb8rymUBnhH1nny1afyyzQ
zejNxqY2eSTvWaufWJW3wphBTrY78rg9HJLg6XLMPGwkII3POVuMVlF0zfM3ZTQw
U87sjv78yyqh+am00kPmARyOtBqMt8GsWo/xONwCoGI7nNmReSJYEc9J+G/ysnlp
3CNPZwqGGjxwiNMcgXr8qnuWQHjp8y96t4V9iqyMRHnUE1lxmPyQ6JTCX8hEMb21
4jCkCG15R3/qDGeWKz1axoStKNFNyT6QhkPEu3WlTSTUyyb0vK+y4ehc5faXwgAk
nEF0YhmkKW7MSrPjTxu4NwNzeSW3E5eMjbBUMlp71b+Xl4pNpyzqY3megsdpzx4k
VnEPrs3qN+0DLLuduLYDHauL5O5gytAVe9flKnQ80wDRTIZdzMwEOHLn+BpE1sC0
tooPf7EVt0Y1Hy2Bk3CT4YIX3mgjAMM2xLg1lQh4N9tX7Iqx+F3NjbDrPcEtxwZA
GJQFYB4XSucYPKFqk9lS7ygULjJqtnOZl/9k4e8Xzw5yWayqy4aAVGQ6nFe9lhKb
JYFia/JF7kUHiR/QtEVOCZS/ted3q63AUkAZbdVbGU/kpB1rO0tJnSX7b1UF1hRj
mNZU9hFTEhvk1Sw0TedmZ1Ng0tHJx2SHkgpg950r7eCLXE4b4fmFvL0IQafE6UcC
9w/c7jka0FLXbvDSF2aua+hTyH36kDR/iWLuPU7a1v8MR0CXf+wNSASKqlnKa80V
og1TDlDb1Z6FwGFTO1jy2i1K4XPZeLiFTXSNXBRJhLeIBGUoNhExNQPNNQw7QSIG
EPv52I/zxCKODdDjp6ysk3+kQ3qtm6cHnUmPcGRB9GNV44OaoZZ04q3RGHoEzsJ2
PrwAQyoWnMoBwzXHOl6954C4O3nFqSVwxCrPgDryBGrtbvPI8T006EYB+FVt2bSJ
tVrqzhj4AGBNN9yHWbbIVnHM/9DByJCeqLcqw2hMSMdYpN3cNDYgjuevdnuaxcyQ
IaXeAt6DmFrl0kA4LNrm1VDjU0ZrbnlCJBhzty4iiFrY+G5rf0AaXub3KoEaEm9i
gc9Md2OAnWVwQJDl0y1j3D0e3DieYg/4c0s/T0OzkkG6EdXg5ZlHREUmh3micnDa
rZvqkm5UfAUsEwxQ1DwReWJK/F8G7bPy/KCj3F0Rk9Ry61f7gfk3XxifZtXk7l4B
FzBg11U2luNa2d7M1luzK9LrxNyKzAPZB7XyNCNq7aF6l/KRgghbprOAZTNT1Lu5
xDck8pb5v7d3wCZU/gYzwO+d6xMuZCTXypUQ+P6K0UBqMktZ8wcML6jWFZIV+wk7
aVJNlJFFgwgBHnn6t1qW65bter/I5XXgeWg3Soo/btNI/mFPyvF0TU5zSgy3CZCr
4b1g5bdW6yCVt48xGZKX7xT2nSwZMEyHTU5TKM8mzCbuVNTGVApy0Gcj/JRXeL6/
ojnlBCzdNUxDIYoYQQPMipuezB1NXmYTJKRZtJogGbrrxNPkANctQXkK6ZZFfEQV
HBcxTrC1cMqZg9hm2ZePL8Hu6fHyWD5jOofHbeny0Qjh9UgXWnIjL0nD5pKqSzYD
b4Hnbcvarl1QUNzCFb5CAlQKUua7SERuLfD/vZq0I6s4erb7jFfrwa4hdOMQOzeM
/iRFPx8UUfHzOl6cmH0/plCly3XABQCnoHCfqF9emI5cAh9+SGeoHiYmVdKKlZsF
ddsQTA4Nq4EWGMpPjj3vNR/L6+MxdbbyoJXZJiIXHtzIY7bDcw3qOMHvZUGAaFoc
1ROTRIL8nYhX/bCzrcAAFlb72f+mbW5kBF16wgvETyWyv9WjRi5OuDNlO1jRBe/o
//FiolJMusMjtaSd3uWnj9fTKezB3lWiwOkV8h7yluTOUbVVqUBNnoQnXfg6TzyE
HzuegCQW2xHv3RVh5DbTyc8wvAMBh5gxQ2VWpCtqIcwj0Yt1Kg7J3PfKc3xwe/3H
IQUO0eet47ZI0gD0mBW52gQ+iY1YZILxIVnxqJBgJyg4YpxpNHauC0VDhNnj9qZx
shy7b1czCFIris7h+FV+7iWHR43SCfV36HJ6J0G1S39XiwQ3NMTQlm+Bi2LBPZd9
2xcxWHpeM+JOQmVQ4H9v2ivxwBQDrjZ3yt7HlqyQ9rWgnBoEyi13ScrE+6x9mSfh
ewWY2AW5zhtLgG91zawwIySEKoKVCi3a0VuXu2AwyEaoLQazwGsSFAJBOAlhy+5s
oAOzema1htjPZBgdfHa1AQJIDkLqiv1gtksTlnor2Qe1eHsY1J5KOi35W8PrV2Nn
cb/arPUkKslQdgsIPNvmHoEhnvXW3IV3aYQ/Qv7mtyf+SvGFF/aoJzvFIy4kTpNn
Ep5GKjsr5NcRO2USdEB8DMb6YtloMgYmoX/owZ8YwgpGgtWIpv2EyVNZxCyj/IzY
SxF3ncIy075WZ7xSFZA1xp3RCdWMP19lN60WwrsRHYJwwRXYA1hVc9uQPYl1ji7z
hrTf3QvAgUcOdA5HiZxoy3AEU8j22PYNOxrfSbD4+SnWVwa26Eondv/I6eJ186QZ
pdx/A08Dl/tg4ymcixHvCaXVtveJHC10HobStMxN9/bjw2qBTIXyraxBHrRz4Wsc
jn3ff+NSqeM7nES2HUoNK5cYtvHAfmYDBlVph3zq7jo2Z0Gdf5pxAxzaFtkgryuj
t5sfw2lKFzVaFsKMO1gRho9LKT7hgdwuqNE9bPd9udp1xoVgaKPFqPqGOXA4iQCw
VLClnjNT2kJFrRIYfz7pR4vkjEBb4J/Lw7h2UGVzFoAHMnxLxyCNk5LrrcuQosua
W/MTgClogdhEQ2W+olM1OorLfDGhhUX2bSQue4W18R57FdnqXLt6l3rXlT2dSDSS
c80M55OqGCwOmg/JUfiSbbwTV+co7FCpGTD15XfWvRk3NBOi0GCTs1xozE98FOet
Avt0HEiZvVJ+BCPF8P2tW4n37Wb3pjSr8XpgWMPv0IfHT38DhKCXl4IedEYcJVuq
U68fn71HXsIePq5gF0C8dF9+87ZgN/BduV4d9m87P4eiSmoYxKRICyRlO8Bvkg8c
VYFXu+rAdfWA3IShoWqX7piizDheCXnk6mbDmVy9TMjBZiQqRaq0G5NZaPa1zxZY
szzgz9vUsIyS92HDeKTt3kCrAmb52gGIHpMPLcE9s+xUijGKh6ZqwoNZHrwTVSDT
thTFvg6fWu43LAB0YEf/ZbzjlwbfAy2gILN9OOR76WVhDp6uYb6p3iaDQvqcVFBz
wWwHwFFXCIXw6YyFEqf2RupH1ZMdjoYqehYR4WEg0ZTHHqAjrG2Iz4+smGTKYBXr
6oi7bljIVC7Kqejn9SnGyD+4dLtFP9A3/9m0q+geJtHCKKNscp53rV9oevhooRux
FWiP5ciirYFirhD6uvA3mHK5HIiy5tK+Jmsyc50In6BsNKSAgKeKQBPKbICjRcg8
k3Ie7RPUxfnkQ/Y90dN4bwqg+0n6VkHCb8c7DOIax9KgSw8ERESLmrVzjaNJ1qBp
Ra2+A7tFDn6sdbJLXInMItH/PMfnPP5TQsNsAb5CNDc=
--pragma protect end_data_block
--pragma protect digest_block
dgGwPUSuhHDslvSwdCEOjvdGDJ8=
--pragma protect end_digest_block
--pragma protect end_protected
