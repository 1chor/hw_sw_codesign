-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vswlzUD6Ht9T5cWvKzzfU2nlUkI9mog2OIH0yG1xlNfLjH7JBhPYUD5eriM84e4KLKGL4rfO5j+Q
ufp0Wr8kNSC5M3t4WbgJvkYpCntNlGEKhX52/jZBDvrsbW/dA4Vrwgp6eDcCNU0/bjVKBnuOyW3m
feJvZIJMyB7evOKi5+dOD/02iUHkvJvHP1gnq9F0Ao1i4iMEHbdUETAwu3Fyyzidw0eYnAtjJju7
5qL2Z6xuVvnOzUUOHwSexJqLQQljE3Ao9BUPoV2ySx/RRmqQouNDBgwYak3ZGKJtgk5RG1zHGHBO
ryiDCK7/0RrudlY2qohoxakB1HyeGf59rM3hgQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 29232)
`protect data_block
8N4UugbcVsYWJF5UKtLtP0FUtzw75EbFJHvFnNjafbYrvHqcMWIclHIADVbfjhV6eOR1ZUxlg3hP
3dABiY4CJcdOedDKwkP91Z7RZOPLtAtsJiVj5aJE1jZFgtx27aVwp6XGAKnKJ56vX6dGuMI1aOQq
FjaKg95ZldeJzjDNUbnkt28nt5emJ6vjY9AgLkE/DCwa40ylKOTlVB6i+t+QEsyymPRxaVFZTELh
83KDcwB+rIOp5iCL6GJFtmmyT5NxbZvzomyeXRtwAs+kd09wYPGZvcQNqfzOAEAUY9vn1QsPRtdE
E0ZqE70soMvVsBcIr1sViz8PXrjxWiSzjBSu5E2L045SvlRFt3+wA890CHXhe4wViDxfqQXzi36V
+Hf5c/rFbycWw7BGpKqTSxSnMHinSSmpbZoGbpQCKl2EmTif02YWDtMS7fhycwxiRn4MV0FfQRV2
U3Pdg/k6QX//55BYRKos7vNecgBj2VjzE4np0oNXJwhBGHbbpniwUODUVZOFy86j3Y5TNRo0pqvR
vOargmSoMSjuvDRX2Ecv1u1WRXjO6Nkwn/jUbbJVA67rv7QRHKTsSGvfjKC0dg+WZpbHp77yz8N/
/bSR1f6btkg38NxDT7PyU9VxJyHXQlW/WUaXkp6CLqtzXzxjR/xglrMcc7FVIbyTQZ4k4broLkJ4
2Wzi4XiSteUc24DOX1DLIeAM6jv60sx29J/DWi8L9BOBLnUnSSA0tH+pTKZRahmAZmyJSNxUi8lA
hobWSifZiFIEDqr58cATYXSE9AJDxa46GW0Q4P36627SaQFyLQm08PZPXJMf/azd6mGTNGgT6xPI
xWp6quqRxdiRxmsyQIIz63XVAOp1xTwuahbI+qqI/XJMU0J/VoQ1HdzZ36cXauIuP3Z5pIHx/Q+s
89P8CqeIY0E/wEyRKokdEESds3W47HU1waRfakB/ewe3sHda07C1oWujfjnSd+WmPX7TvpszznpW
aBZMVh0f+1WNvcojBUy5wDe1tspg2XJ5Fqpce2RqTKUQQLXT4PFsgHI6TgYKLeRLTMyNU6Kp4vmO
ncNn6368IwSBosbanX8L2pLiDTDNKWYfna6t2mme6dVicxstE1XE5hic1VnWolXp2f5BzpZdOvEZ
sE0VjWGHK8TkSxMA0Fc2mTlcERc840u+9KT95v2RFkXFiz4TGTsFjFH99wNGqAAik23Pj1njHqL3
OoDKckXZN2q8eXC+rno6H+ZKTjv3jCZDAJN1pInVdIPwKRAxkz9fXXiUhQb8a9jVPYwNzgSVjeiN
rWl9ZHjxnLmA7z5o4tcGurmj/7sJQDrMaleuRlJie2G1kDLSvHyleqUB0HbrCByUEF+8c/eHDVH7
ws3+P9zgJyJEvQHwEuP3MejS1Gq5iQdIC5xJ0XWqlHTmFqzBI7lkXo+SLrwFuclEh8b4AfX5WaHU
Bmyef8z2AtMyoH1jUF1Mvpvx9Wu6SsikIS36Lq9aBWS78cInc2X7KvwUhvg5SgYD2v94B7sJ5JcX
Z+sbj3+p1f3ykHxFt+1ZYEGJ0JOx7HOe++4GMZ5jeivwh7yhyCLeI6MwxcHnCdlURv/3Yw2Ks41b
wAvoyQmIeFp5CIjWKkJQFXahH6qCHFIhKWuIXJjUbeyV1xKDAUUQK7NKWwPYEaF7OZhAT52mjjnZ
T0gojTXI+WLLWc9KXQGqm/jkBRsW0uuyOXYi5Z7YhzUmMRTVuuqgw18kOaPGy1k3dph2lnueWryN
aPy+SLNR+JYbbUvuHkkGQku+VytQu1+8WDnImYscCKl2IfgDOc6HiQExQ79+O6V3Rb2yoMCcktvA
z0HuILga0BQI/Py3GWgf8fF/DaJ3I8w1UKT7M3EtXGcsniUcvZnXuENkGoD3ldR6wKzO99QeMe6+
qhluGQ9yFsygxH8m8GapgBJNQp8hWn1K0+ccr2H02BxCXtNQqupUYmm7bMi7QzRCtA885e2jKF4m
zUqS+fUg9+pYxiByxAA9B9Xvvxr9DZsTq3myJLUeHOHLo01QSpKTw+NzHrdRzI17AxODRdKUnfSc
u3MtKe0D3hX5EPvmz5gcHvgNOyLxUl0oeyHZoxMsIBIrVDj2LMVLsyTTrmCDXzNRESv+c+IHXFnd
0iFzV6dlD91EDtqcvn7tXsDSE1mpFAdoOS79WD/Rhz2RLjHT2G4dmjff1shKWVXzV2n1X8o43H2/
+Tw+GaRyc4ljlq+qIlZk8GFF5vPd+jAd/3PB/UClzznkjOJzpvn4tZbEnbr1J20CtxbZt6t42p1n
2oYM/fs2kjXkl9JgWraHSxBzqLi80yWjqHxD5u73QZrdTfNILsxdCzTBPl9mLttOvjD6dqvOzkbb
JoZFDOgU8+4IB/I+BWodD+R6WbpIPRpouX3s6iXkQrIn3ZrXikHAWFgllWCwUbPug98jgQm8NoW6
jyHWIn3X6n3yFORAeqhlk4Fk2pQxHk1UIPdQ9/SaGr1OUNYaYawE22xVKmxMT9b0oREWaERy33g2
ZXl4GEIycJr5ByMYCvYWFF50GxG4U55u1iBmYYjFzLkuWGhiVZY4jqtptBiu8Um3miPf5pJs2F9h
OxFtStGMJkMHPjd1efCkw0PCYHd69qotCez4tx4pxWHRRUQzU75R1Y4ZtQpOiS6VM3NiZSoHJSHV
OmK+6E35AEVOM0c0RjYpKtpCgxzOhOgOo6mg6sO7OS3TapGv2z69ILdxIbnD6+d1UfcI5JY4h4OU
OQ2wreQuRSBb8nWpCbEh2yW7TtG5iUVPsrDfN/T0fxRBGGtUqvcfOsVptvPG28/+eydrRSzZk020
2e7SR/YiGr52VpL2j8FBh53TqsQJrdvhWI1HSIXx0ntefSczfnYdCuXUVdKIAl/pfMJKG6UAn5jp
4ewuNqH0FRSNsUQObb/qPHKVX1M+Bp/uMbin6tI9tVJcdIi4tBSSz3NJ0Uqw4+FmkltPbwIP/+Vi
4qwOIfnmhpdoAl0W0f4EDQcla25qeseu97EcFlIs1JAnkg0eKyYb8RKaYiYDCQMGHTQJhSWaLMhc
th8aLPNsaqeagN8O9a+dAbrSVqkvBm1rdxznHK2z1exc+NpxpB1st8Psr5tW+dTP32D07PykS1WW
Qq7Cttz9RHgo1cGM1QtO7DKemAa5RD1Aopnakfu3XIOTxT0cL0USoy5oH1f20kDaKtVPFEiuNeI8
rX4/C25h7K5zDIGJVaF5On6bbEalX9J3LWjA7NUYySQdSRp7WhxTO3Ow8fYa4Qy3FJMslgIKOjlH
pW76seaFCqh6YHrJtpaJzy3okWWC+zLtbYEsqT5/T9P/ELMNN7ywdz7rBk7rD+KXx08dMfDGr+kd
CppPXdm0DABcCMoaW4po+imKhcedCVsTzuMPdbqq5RvkfYheQ5m1ufceRIdI2F9xiA5A3qsCJ/s3
iMEnYwflFWP8xhYxwVwlLWLE/FHULL/ukRO9StAwetMr5RF0mmKQHLf9zyF68tPdmtGIV6/dvhHe
vipEH5bCMcV14mHbeuHgN3n2RZW6xp9K89PK0f/nN9Gmt/iceZgUOwnUyeABNRHRDEtIC+veQczo
wesewuQ4UzKKTAR7NXlbw/HxtB5uu5ZW1FPEF+myxZymGEo/dx61cOEltJDt3CCxfzhZKrylOFgp
33f8mA0VfAzqzVvx9fwRB/lz5l39VoyiWi72HHd9r5quDj5eN8oIOc1O0rDehgwjGmdyRWpurOct
evOMjZQXQ34PrTOMYybQSGvbJ0aq3L0H2mYUMw2Vna6o+wcuJ++VYPK4dZNp067xy7Czcke3dcr8
iW5FTHVPiMwsuBXbtCaMDqItF2duQh8w8Q2G/Pmde+7Xndnngp1YuMEBHf2yCXx24HjvaRWolsIm
nsm6+igSOHnzIubUpH8xbpkOTWs5dSbka+JUR59L/tgXbFi2X2kku5RuNysdIYDCgSMm6uCRqtPv
6mo9pMaqyEUfG8k6P5RNyUnjIHxoGl8I4MFkWuezbBAQFrRgszHbk4yL9K9onb7GpLlcMjznvQu7
YEZSnuk3VOHZtPPsZPnasvBORwvCp+iiIAHMNuNIEn36vkknBApPdFKUy6iLrZVnT337moJ6JifA
74iD3Q63HpD3+Kyt4EoESrg/ulSXYiFUtpswOUdP/umDuEo14GMyvV9YbPuYnql91VcvvSbthFwK
+8A5NNtJecrgGlKN3srmyuFM5SfqNsK90v1rTPx1TAsxNO/CrKIFdVw+jHyR9BmBr2fycDWGEYi1
tFTcsYE/v7kNBTeS6lbPNzdlQIVT4z9qqxT8arAHQfuEvWZIYENhNSk54EwoJrLq0CFxc2GeYxuP
52E4TckiA4+bQxkh8ZJOMIGJhMLfXb8OilgXPoZ3lfujbr1UiioJedLNRVzQJaiuH53dLjq4dPmL
VnBJP86zIUPdDBrmpINPjoz/M2/Uyp5fAdBJBDHzFOM/aKsyzEuhNDJrfvbYjTDRMuXrSFW3rkek
EmQypkxHI8PSiEgFIX4M0AQwc9AS4o/kbnJ+wWtwphgy3ru6pqSRye4warUBNJDWz9lW4YonGD0z
OkgIL8+q5iov7iukXXxxTlUtD4ldZsS2s/JyrDqU4mmItNPytNN6bTmT1PP+wdUkwoROEb0uoaDp
7smN4bD7dLTZRWqseQveQqaK/sDfmNWcAZVlGHGZyMGImPqxvsSai7e3hw0GWoQ7M/oyXhW3TXuO
Cs6o+JhFbvHOhPtUx8RH3qr/wCTIA8EBSbkvx97Kx8GkvsYGd501+nEUlFMj3pNVUw+yUq1QnLoD
adCIYsMzk65LKJCSy8YpdVrv22RhLDAdTh7usMmiqYxi3fhjKP3nMMYspL6pmMF2e4tnOSgnSJrD
nygYhm/PneHAc4g3oqXZW3Tiu1AyasEgruDhuUoB5gmuOKTKnaLoMiBXgI0F0EyZqaK7jyXS69Zg
YYWCkFpcy4EFlggthYc6haKBamPekin35IbqOS/Ma8MfH41rRAxVlZT5jRwVZZG4GyAn3ZKhp8+P
+zToiXht3HiTfoMouD61ZMtVKPjI7WsyDWhP0xtV5vCa796812G/oCNrCHc2S5C+NqZq2bgtp2wM
B72CnpGSzgwAWHqd7cJLRlgIQjdhn+kEFbrgTnBSJsXfqdOKG+q9bR+1yuSdR8REySuXKkSzE/Xs
ZpDA/zfAbtIUkfevbKCZcT8wXnYhlb5LAbXll5A49UFUoaAZrKIdILP9u9CYwW5VKZjQuPru9ADx
6Uz0FUBuTz+3h/EZy5U1kofBE6jNjaOn5Z5eH5QpWBELrV0y2TYJKAt7aEugVbbWgMXs+vnZtU5T
CNQ7M3XSss6YAT2rOeBvZPQKRIo9DMBDmYuVN1wXXPtnxRGIsbxaSRWL33mH+FYuESTzf4Q6yp21
ogCfJhjpzQnAPJhGkUi7t50WP2AlSv7mU2/u+DgcqrXK4ldLdyzjIvsKZ3QNl0as9RgH5BizT85L
0qHlcNvZWp+xq+M42pFJz8X5N4C09+L6fDLqwY/8Rdol0uVsc8npZ+PQd9EQrDJ88Esojl/tLSML
Zb1xLU6v/+HfzZ1+I7njwPkccXvTnYE19D+4aHF2QNQNyVk1Ioh+fKlJE9lW3F9HV60c1qsjOo2f
I6Fob/dJc9/FDb2UXO0s8toMTAk/T6UqgE+VBjmfo11DVtCj5tJZ9bZ67TfyrnFH+t20vvGOsW4O
7N1rFTpdUfHOosG3oEZd+W+sKlt82hjSndjAPpFohTeJVosVM68JDgQUB9ExbbrRd4szsE7McDK2
brHREb8zeJKxCuWx3h26fGf+5+wBm0PDLkC/qSI7GbtAxTxrx+9DKJYWhTnkoRdVL1oGLqtFVvDo
6VUgyLwO8h4n2pNjGmQvJayEPMNEeACxoQkiMLXls65Gjkt/31+uLOgTF19sghviMn3uA2Iai/cc
HlToV9Ksj6VPe/HEBToyS195S8pmsgNVwmUcls9q8TUKuAFzzwMavL+lUSh60zWmkr+JRcLwB0cN
Div53KoRWIo869Md8G1NmzbzF384PS4qNuQJD/yjJHeQMuPI832YNrw1Htsf1T1w/cSTM4SptGQD
s28Tznrexch8y7cVsHo4s4TZer4IBep0QIcPnCp/WA/XccLH/tgvnV0dHM1LwWq+qDsHtKX2SHxP
3StZnlEdTVLwjRA96HJqyhDYA+jYydNKbQFruIcrkdkyxJHLx7/A+IjEoow7t+EhDIZunWwxxjN0
LMXFPfBljLcmMxU2ewO6bdBVf+HWjcUOB6VS49VmkS6akBlq7aA714Vr9frQP8jX2OvfSUiJRaTc
n33CPDcGC6Lwg5ut0s+kg3m6GAfbY4VMCqVu3IOZW/udha7c8sL0kGHKe7NjnNGs12YE9wHoxsYi
WcRRWrv7PjZ9zzCIXD8Cb3lMFG98Y/nb04BB5Me+YvJGEP4HOHbW5COTzUArUI5E4OMRR9he/kwE
1AcPqbrNNfk7ipmlK9v4f2muWRRyLn1G3zgYiCrnkPwjxwPxguId/u8hTMUZ523Ol+b0iTwtzKMV
viyHx4KtyMgWJ3ZTDwc7GILoqEteJbMiSh81OASpGTNj3m76DnaU/T0g8bsuM0a1t0K3C9RdDRnN
TpMuSGHp+4MEKjpjMGeuX1x2HxDWzeZ9NXAAE7qTen+ivPzqdmJrPw9V35F+wc6/t4PSaQ0aTZhy
pI/6cw42gUqeT1spw7FpEy5CnweHpec/b8k0FPAj66FsKYOjXPms9OGqLSxUH1tE9BG61bF0H3qs
GPsSk4lE9M0/KDwoN50wyGMIm7PfYThDjwOmSH39flNqGjaaPK449s3yMkrBapm6McuXTjfZjrey
YCOpTcMye7tByXSq59xVxgtmxpacDDsA1eRrnvo7b3daZDrfXpHjIRIQN4z4y/kyxtWsEyuTEJXs
GlhJc+zZ+ymF6frsRHH9Jc7dLFQLaeMrV72riEWVeIGR0AaCkRszEu09Sd0k0gKxgXe0UTnEXli9
Wedekps8VVzcS70PFPVLVyNoSjnmkXaaaEvzCAoB9rSZ5LK5yl1H7+r0QB0qwU2EbBAFpPFVVPyl
vW0ux7qd8qJYc43u7lppYQQaKMokp0ywpGC/DJApCplzRHsc0paO8Dv+mkq2XcoERhK4gyWTcdXp
KP6OQg7XqJ54+zxZeVjWU6L6V/IBT3ndcLYrBcbfH3caUSpal44ehbWJdtPObb2bAC0QPTtEOYmW
h3lL2f0qGZX42O3/7fDMIOCK93OaRx0qwI/nKiEcr2ZOQjR+zXYDCknTKK5UVWnWdD85UW5ZLxO6
lQdLSMd8E96iDth4f4kux24ye/+qJCVk8C5/9mt8WAAitFjfIxXqxxEZ09TN8JJvZneytT4UKReU
b5PCDmKlfvnm0SDJ2mDu97k3mDJAid0boMXBAuv1nK/TZgwC1qclTB4LdepASdqBbRqvW1XGpYIh
9HurVvjghDzuukwzhVDgntJZOzfK190bBOl831BknxCX35T42W5+DLyXTRLRaLI/BKbieOsrIIMG
UZqeszFZJS0oWpMSCZQh/cFWjU/xmIqUICUjbLPdgSUerkw3G2zU9gu6Hf19oPdfkguJcYO1BOKt
8FW0/ZMalj22YJG0em62d7/kv9dLb6LllL8RH27nzbLP0BIuDgDGkVBO9VwCC+GDs6R/2AQbIaa3
1Y+/MZACtUZBbNvm/eFFpPyPcDi3TNDdHX04gJurlZBZEdnJeEU9vtR+/Et+MBC1dups8EvWaP00
QkDmYS/MN2dTtajQh0YRdrvsiPOOW2zdOgUWhnIGKQCV8UyNxGyDRlBBLjV0Wpai7Cxepi4a1FNY
DIkB+LCua6OgKo1i2w2IO9pF0QJccktEqK8xq3u3uBb8W25erjGFnfxyZA6PJnoPQMoZDFTZ5IIS
pd6Do81yv3UlOXFdrsbKqEevY4hJYcp6w3xuVZ/RNTjQfPCuMLU8BQeZXjXfJQgZrTY/6unZTRPY
VYNI3o9F3XOj2RNvBYb5lQ0k9rXCPxaLqsVVrCXtzFiq3D/nZ705SAkL2FB8giLv6P1RHn8QnWSu
fP58alsglh0elXOtNlDHqZ7/XPn5rrXF+GU0fWqp5hZz0YzR0QnItMgCg2MsqA9YMWvglWWBJYLc
ajjmSngeSL4R4wSVb+LIgCfw+iJ7+ZzGQYi5rP2TvOdTzKd28+qcx5paDmOsfVAG8V0g/3zxfsjC
f7/5KLEoO9XRrOvp263TOedXWu4r/cbWPDOtgW3tWAIgPR3ktX/GX9HkBH9w+OhtXwUXHasfCe0z
WFLQCpR+9m3yvlWsMx8JonnNZpMEVsZWGz0pk4DOYFFZ29zSBVIx0SNbRq6TymKsnQkWavLfJrEW
DkAm9wmVMm0zuFNmdq/ctekC8r2vVkDw9EJXfVazt5ZyXcgQGiQd5csd212CgyIqUjCUzqZp2PsJ
GjhQuHgBeBEoTLZbRdtU0VLvCmCVPA5yn/TwQsxsBUw8e/Xz4bMnlGQ7A4qkdM/x0jowcDcxyYh8
9A1D8Q/UIDopH7e26jEto0rSZll5eaoOGAoPCnEAVAlQeoP7sBb4fiySHJXXV6wqilGn4FIjy5mP
qxnjtyh6VFMtUaJ3nvj4/1mVSai6ORh5KSczInJUT+occqV3EFLeTY+7Q+QmlCkCJKij3QKqsIWT
2Vm1mZtlaFfQQnzGdvMFIRltP10PQnMPWuacv4YCnw0zCTu3Gi6Dgd84aMmGIka5hsknvgQzbRfw
79gKTZQ1OAczTkvuvwYufylnOWIE67g+Fr9CEX9aQcreQ1O4stjnK05KNnMmeH1y1deHVBG+nIE1
pG/XMafXYYXLNazp8pYQXCdF3Vt1Tub1LrLk/AgO6L4CUGhFOSIiaR7G7biaHlXhW/eIKhIO0UWH
MX89jLQv1WRk3e1J8B1Q8yeTYTDnJFnGErnjIbL8xp9WYVkSD+7rNvoBEGgdpQOowLq4zA7mhNVE
Bqe2QU6vBIUucEDgjkvQIjw4Wsn592EwVxXTP4RowLw0ew7AdS/aucpD/DyaAyq6MJxEl2th4bw+
gK0bqBVVwr8uxy2a3Nen06s55MsY4nDtSk4d3GMq7ryzH3RsZVFLmJqTSn8ZWifGMQTSXqz6l3OW
G+6nqraP+Ue5Kwzeou5KGc8VUtkv+2yZc1XOXZ8FY+WO+egrQWcjvKqQ0wDOdJYVCxuqGC0ylglT
YF6SELilnvIBL0q2UYQdvR1rwD9MYRankr1a+4NzfJVL/QJb3Zy7mh/BIbWbB8qL2UlEna3vDq2/
k31BkOJpwpvzCME8datlhykoov8vgeEzSxqUY15BtY2nvmS6HLqA2m4p4unRIcc8N8Gkaoh/5KuZ
k7EikJAgID5lg2v/fpKIwppFveWa+GJYQBFez9tglGGDzmJCjI18ldwbq1Vms5n4DFq62cIBzYMK
8CjW5yzF8WQESchzebcaj+yD9gUSB6toyUvbqHCrTIxVezOToAYvlO9eTXy6VRnT1pui7T/Ja3SM
TDjN4v3h8kbxDZFw4YARUzhJGMd2ihTAHnujCffkitW9lh6huccPhR67Xq1Ci2H2RJ8sCtpi6BTG
kWb7H3Z4zws0OAo7kWPuJa/2qYBzP1BdBzOrcVhQfy47C9pnf7bona2EVqO9eVNg0t5Kr+CQyChs
6GJK89ovpCJXDfA1OSU4W0nzfb4qqjtkPSvt4X8lWBJxFDn3ZgA4YZ+8d+JV+p5u9J1Yw+cCjQ4n
bawCJxsB2LRP8rZwYQF7qbPAVi3/2eag0Q9+1q6o1YTJusiNnMe/qWmMXY3hiHxEYBVBZA7+a9t0
DMrY2Qs+ptJTvBvw1+0Px+bnF6flvAa82DVRUhHk0j47FkfuKXjn8Wr1bxBFSiqd+K6cD4iLuGvL
QsNOdQ73uT8VRjxmetZMhBewFXe/5Go3YTdp2SuHPvQNBDVqre6HjUDx9xZpux/kf+50CAojJN1t
lKJ9+16BZewShRCti+3xLGBlx6bmoxpQTPnpM0VqWkVL1spXn1AdHF8CbysHR2W3dfCL60wG2df+
mS3F+jdcfnxtwm5zN+Wwvc29pNS+2ZrGPWAir0BzdHdAy7Wev8P8MpM2i1DURoxJdi88jq3NmemT
x9zkied/rmdzXzNZ4dhguubgF8w2BooqbQi4H9T8rYiyPR9D/rIwJWUoh+DD7sdMHmeji/24iUYR
Hqu7HWRA25niSYL88wpi2P+dGBRf20//kYojuh5G3Q0KhCrTNwz4Q/Ty9bkozYxdT2AvPf/hpyHS
BwW6SmOwQ0u5EwQHJEqNhdwSXQa4snJwnkSRk42NbLBbQM5u6t56+Q0Tzf0CONtzuaA/cHtJKaKi
SrF8CkvFQY8OwWsI4j/o5WKaR1eEoZYvRUYg5jmVCaVYdWVDCSj8xzsUtggtW4+i2I37xWKJAuAl
o3X8QVaFMy/+Npb4KTh1QUnQ18jRsz1R5ac1tmz35Bs9RCXmPqnwO2lAuX4ygL1VN2Zaynuv2YXO
74MCDBdsn2dHsLsUingiEs9XjVWrJUaTiDNscUUo7r1XSRLvpAR+fQqjeFbjk/mn90304UgJjrmG
XuxCpHm+LNZ5w8kR40WhAy/JYiqYlB4mCh9yfYtYbl/s5YKDZOOY4xykpN5nJL4ja0kpEqsDH7eq
d9oqY3d4aHEWreeYSUTFOu5OrevmJhBax9wx6cMMimkwjjqWPJvvrKJEj2WW7IY9+lS+id4PfKAG
CTE4I9X3lJhzxvyyTLbDPZhb2YujQMEL9wI/oNGWct2UKKZ4kX9dyYNWbKZ5RlwwTOTH71UKre/m
I56NlGDxN4wIT0IakQzI5q6X6gbHNXjvifarswxFQ3gs6aKlivyWOFRjmv/NPNxkZ+efdQ9pnJyT
RRCYjchl5KTyphyDvoR3lCGBRnNPRAhrtm6LslhL6RnGGCCROP+g9s37NG06LisncwyvKcLDNweV
igpH+Xacs6oLMiYweDtY03HSiWwhNHXYY7/NVjv/kzWEdqpFHZNnaCkmdBE0WLw97VbKvh7OqaIK
NpjC00yIR/p1mSI6WJVsTcUlsu30pwMxK+/CHCl+AgsF7eV2KK7ZcDom57H7EP3962a6FDuTLH13
Iq0l3fxbse8PrD6xNQvavvc3LiYz9Z0mwrXUqhHsNh/7vphHiKsG+ZrA+RlaD64OgaUtduWLpOax
ckDNlVzQuiCT4Y8Cbl5iL2EPlfL1cSqVDz5BoGp10J/x+RSMTaxMENUd+r8+/1mpxMvvG1yZtmZD
HtFihX+JHsGr3ajnOgMIC7YUkB9BAkIs2U/6USAt3XCd1VnTTgaKU9SCruvFgumUxtuN4lg7rw4T
2o1ebXhBiRJ6ZyCFGjR4rCIFGOPg7YHq5pDFoUdkyZutJm7AXYvhXFNVOJSrCJ9qDwx3bsEoY5ub
PVi7na/DfYEP30iOYIQU3cXwJqWrabGk64B64tRqWXv8Xjuk+3WQutdZUGeOO5+15AgmEqq/qJuC
cva+6nF/16V5flufUfTGGYrML9MgiJznvACgW/4nZ42JlX0UtIV2uCjJbzYB/maKPn8lom4xOw9f
mVe7rPQigT+C+A7iEMiSP6yGL0UkNMsNMbp7cb5HTs/mMAEVHgiv5xqFFX9k3dyg95+0WOSeK+hC
ccnYAiyKGcPH2qnpX9ufNlFC0Alt6bVQ8m2GRenRSLvySPVvkag14VEGVl4h3LLAm84ER2ATRyx/
mUQvMhCyoS3B/ssULlwIuwe56Zln83lnpIEjC4TwGhyAqkdqoLrTcxKq5rlFLiBQYma8H17IsVIv
7R1tjk++By6HeDZb+xjWRItWc7RKyHoAqBb7GsuCZwSflLd0nem1FYBGs4oqHBk0T13pSGdoXGzK
oMJEUD74/py51vpYwbEQyZA1M7AiR/Ao0AYVd3YMhoa0rJZqnXnrs/SUAZxBPyrMEKH7wxwqXYli
olNZ/BsZeGq2lthOao6krG4Z/7sCrBXcXsEmnx+TyDuekNrm+iQccs+8WDp8wgsPYe0Eid+SxTTy
Lu8815YtCaIC/AOMYmCVWC6b3AIY5Jj1lkZMygK8IS+geesG9g6zH9eMCAGfccNRfO4Xsuq3K1+S
4um3ZPj+nFzadOOYTEUs+rQoCkVfMhWF4z0w3W5+MD3FoRevBXAthMod3lI6ImdaWvW82yXoYrYh
cUm8HLDm+0oZAKh6GCbAWzOFgzG84dHeokvpgssyKjFdvtYQa3y9PVzLpVjEQfFe83iTdCLirfEn
+X3B14Pj7gh/cDv2Jx6+S5QOg6pwQPVyDdbO3QzHMD8HX7st6tNU7yPiTMeRIvRNBeT95DXHl/sG
QyWGbtu+UsCLjLofc49SMcbof67VTwKlhqPH5+ZtrtDJnB04INqNTel56uDEktjRMob8jRdehyFO
0ZJB3dYSX7Q9pDgzbrTfOvBc3FmzoNtYQijHp37dzFjcz0sr87L19Xlj0k3DedR3ZQs2oFQhpgwZ
1LNNNysvv1qrZOYNvQc6J4wDGb64qm47hoP85vW+PoTDr9mZsmiPwzqdZh6+7L59EZ/xwjziCT0F
1uS2EO6bBI9JrpLil8LZylZAEVPeWYzsCmp2Xzj2YY6TX9ETJXI04fQCVg55YO9FQUxk8MqZxG1u
+vmJkAV6A9Y8UDVDS/MqX2gRYgXK+pwkjG6b+h/+C4Dufs8p4UuKLLcngQMQ6FY4dZxPHJk5CO1a
TAjBMEh9dCQz9FhUUghPM65qA1g6VHTpomqzDenVa1RsNVDN/JewfBmYV+7StdPjV8j8kH9IuBWj
C732YMVbriyYrcOQQ1wc9MiJ5RxX5sqAnHgRZRLKgV5gFUqylNYI8KyZOT2u5wwrq8RZZQ/bA13U
Vg5MrYFl5zpf4jbKPTObctc7QeXyfdEbS75ZXJZNXRrWkIp1xXSpOXIeFXc0NYC3yKgG6jkEOsd/
5MIX8weyAYxTGsgQ5IsEfLRliyLWjD13AwTYUIhE+XOinh+hXb9mkLM6jzMxhlyuQecPOeQbkTaT
GIRJMSzwAKBwwh5CdwNUljq9CsRhq/qVGvf6MR0sGXpHfPIHglO4IU36yVy9Mecb/MzAzDpVQs82
KEP1miE9qQPxsffyhZStiBAwznHxSYVy+KEENOtfZzbwGHu/tbZClVXIiSsy6NSH8TmbLz3aXg3L
7TREQKQiTY5MztvhCLfRKPZFLRBg7hqfGxeLKaneWBq7LtXIjcoxlugcpBPsZZpzgmRnvhhjeo8p
Ev6gSmn9ydiNWd2+4KoKEcdh0uifoMk4/AV/dGKYw1iAnThfn85T9vdZJ/z+yzolevps/NXVCrqK
MB4HYa12XFwDs6m+HO56siRl6PfIMorFA1bdxoAKbz29bgvEah9PZ84SnN5/dvNI0XumqGNg3IDn
mGRXsfY6LHMGToebA66i9Ejlqf38htyHmxhie/tCV7asZNZU776jpDzJPKY9FRax/WOx0XXLR9Ah
e86R5KEWcuTf3F6XvU8DA9WV1ohqc3V9RVvJD3psxogxhFaCGRhrRtvt/bU3/R/W3ANsjYxT8xM7
QbwZpERmOvIgfEoo/VsKg1S1uRQcHXbIa1C2goG99xPOsdaKNAyQLHwsIAf5pmFnvayErFtsu3cM
8f4uuHq0A28BRDwktOpyCF7QCQ2xEggjnp5FAA+T/BY9rRETQhzvLEI3DwE+eYIXSflKYOXV5wjA
QqtRhPqbNOVXwXVZ6SHdheX3AA6PzRoBqWHzMIlHq6WHhvuER4Y10KqVCngks6DfQvaPBeTAfpfh
TuKIgw++m6azm3/r9WtiL+QombHMfMRzelfAobefSSqH65Os95951ResgYjeFB5u97pmCxVVbucb
18KF/48t0Q1ZPeKW1ZYDXx5Zt26erWOj3RZNNFuxZ3DCBDKYPaA6R3DNtb5py7X2tMAo6jqbsYg1
zdhPLujRUrLXAkOOojlk1bY1japumr3JKusrYoI3a4SzAXOPW62vR2ZZoK/o2C8AG/K+5TzN6x5v
Ei0+4fefr0MFZQmdON+PpxkWUEtYibTTDEyo2JkYblj1CPHJ/pkvw4tp0Z/BOOWIt7n1SXYFlPuT
1GM4uhBQMD2kvQM2Z85ZndFnw5fDWHHl1HajdfKLkaXvEZvV+ycAsiTcDb044/qnmvHzPc0P1qZm
XF6ruQyi1PImBlOFpCMrf1sbNJkeHvKrge7x0MTKA0QgT0fTWieW3r6QwsSr7u0ZPsohxsdzUCz+
boQ/0DLsLbBDcvy0Z8cAq9Y0SKL1Fv558Hznlh5ah2jLA5IjDjdKxgix10uA6eBUgBO4PbeGr91U
OjcUsrWwnnj2DJri/sGhRpQhbH2DnE6ya94cZhyOEHqgNxo7lepo0DZlS79S/5lYJo6R3wNaoyAw
fwBsM9SH4lJSQ2ODtnC9OO3VvrzFhxVvDeYleap/LRhnC4tBV3EwiQwT5vUb6tb3lm9e+cYyk6Hl
u/4mdkk2vTuRl043Pxsncg6zssxogkqgHYy8+UnS2CDxMU3ZW287FE1UeTZUbqAyNOZwtwM+pEs0
hnbGEgp2zR8YpAONqAHUbP23idqAcm0CFMrOhl07daHCozXetRvPDmWbQwf/2N+cy/J0p5/XPyXV
UgQmedDpMGXTfLE0r2JuBrLrUBvv4YNnL+SUgQPVll8jZpKutgpVkOsBycbFsvOD8yqSr9xMpEem
7YmM+hYfqnZcjI7m5iufjtKx94KbtTvn12BAL0FkhFZvkaDQqBZxxf1/MeuYyi6nSbDPn166g5Gl
Do+91LuM0MOKjFLMTzaZcJHabgc0HEoac10ooSNytiIsuXnq28/2zrM6ppAc7VkXUBVG7hX0qZIY
IZjFMEb8lkeT8DglD56mV3+qjd1hl+xPwDLMmtawf+pi1wwo8KDZh6cqo6pciDqyVtJ5glFTmeL0
qRhZ2BR2ZmlniEFw/Ee3QjM7f7ppffPYLg3VXpkn3Hw7DAa+V/4oVYbsoYKQoIOfHnCY1h1s7R+t
fkPzIFo+cKQKuhT07YtnqTSTmwHHPf/o0PP/6WtDzYXdGy+e28mGK41cKNQtTlIkTDXaVMnPANPs
7TqBC256X57l03wm9QfyYRDlpvBo4AqzFfmWcBP8JF7I8F5Kdmzq59o/7rr9b1Fupz6+rHsSif8k
BRxXz+z7Ng07LJ5L40XgtYwjImFieSf7Xf7Xfuti452/neblkoDSn6j5csvlJ25VsdBl/LQLFnVi
UkVqjD7/2zGvuNMOEl78ZY13qoRNUzGpAzVTF3np98XB/rfwEwDL3NuqpiE6ckqK/F1Y3oWCLOMd
DFH4xMSpcon14AZ4F2Ttac8U+t2MiuC2yo9xuL125c0TnXZEjVJupJzA4ERgiarXh5axLUse54ju
nN9GQKmA2S0BXyHrquLwteZvmHGztn+yd/baH1BLuKq7iAqpEOzt6/oQ1uOfomBtEjTHKMky+2Ew
hpZGr+vpDzdFKSjDUkEj4GCu/M6+d2vBpF1WSZuLzsx/euTHXvO2aoHFAVoamen9JzmrryAGSU91
ZlaSjM2JVNJsFUg4CmUm3eJ+qHhux7b32QXegNoiwHxlMo6i4h9ltNAj3B041R59UyaF3aBu6Z4g
xKWOpbGxrsJej9utetV8pNerTJpv4BwdR7PwRwuotyqsVlCuerC0V7OfM0pMXwD51zrBFayUloff
IgJ5exOQBJy0DESnGpAoqogsx6s6aT8haMTS8QoQQpVJTeg27lCR4LRB46L6Bj1LVEftPpHwzEQG
cLitwxgBsfhWc019BTmy+JJ+RzlHi7h372f28dMie5On/O0e5dwGQvDvk8E4hj+ue3Cd1Vs5La9U
G/hWlIF8sProygg1vYDXtsZZkewrJ4pK1U/ct4WeaZQTPpyGk6gAP6G+dNYBBgLvOfm3BrQ1Ymk6
e9ZV2uVJs4W8JC3zQDB81erFTwg7Co0BOEtgjKivuJH2NRj9S3zw4bl288WT+tiIQx+g+GuzPCXN
AEkQTpK/bpF5sGv1/GkqtCpT8dYjtnZteb5qvgnvuVdmG4WVm0mrE1QRNKYcWhgeFWpYFGZCSbz8
BGP3M28JFAwxy5G5zLmnWQRfZUB1dkLux14Y6azX9C2WI3zOzerHe1Q1ql3rn2ssDxJSU/UsXpHm
4pCz8KHBrvhS83ilkFlvwoT32o3YLAMfMfL7Z1/ZTGp9G773jIMxVb4C7vz+WzvG8PiJSwIKuWK5
VvGB9KFlOIsVUCbWB24/Ux/3Z6AqeP06L17qVfW928pqmFNp+vi39XS2qoK25E9BsQDBw8lioA6e
sLwLEnDSDMTkNXpZZm1UgiMsMAVb0ygZlh6l7LCgKqtMQcE2d5qg3eFO3ZOn59TVDYuLdahf7qbk
8FjZ0fXcBQQZou/JdpgeA1AFwqMLW94kSbVPogGN0wdZhQV4Yj89NEr7KqvE8LX1xPLfNLtlX4SH
eufXJorTmpN0Mqk2T044tewTD6q8mOoXU0jQU41KsuRP406sLdWmuwFxE06Q26kc57KkYip5ahkY
fawTE+PuCyLbYouHq1QLcnLP6sAF2dGb7METgJI2F/fWYHwUIxcroAMhTglkZ8oq15VvpcjsWDS7
rbbUSrRa6wMTh+GWK2eEh6E+F43GGM02NYn0g8aH/8sKBGuKy+3/9rQF+HA+V+yXUtcIlBwWnB1T
khdyGjnoXUxOqafkDp2nfanuZMDNlmCxvSBzq91k/7A8/eBvQJpMIrydCDpEsCDMoIrGKOtYvLwB
DB2nDHhEj5Zg9iGB1a+kPjpH3IiwxRkXRSER4p6fE2k15wnqvgpc+TnFJEB8rpEh4ehuihlrF3DH
8ObxHlplJOuvn6tsFVhmPvZklqXbXx+IIzhuTNZ7mkFwZ2zcwrTOFVghsGSxdUgkIBYIog4hK3PY
2yqjNxxSBrx4iJgeaAwhdLTiN7OW4xWN8RI5HQ4jYVvarWVklU2GZnhNyosM6i/PBHPm5MKmqBqD
burq6QGGx5DptMI2iU+qIAEurhUljK0nUjgtndiMpsNZ62vvmLXKQIsIrunwDqmLRTHhvEdd2THS
/ycLlM2rIqRXetw9NzLGp5V0lDbil0JOhpSfqNi1ZiGaYeN2WraqyMzAkxuAG701O59kmCyfY2Yr
qczXsQ12WvFtq7sOYL90uCtcE0yCh0x+ZvswkFQtBc/nqBIkRoLDUHWg94xPy3Pu+5QgOwRIs+s1
O2yLUUp4kh+Y8dxs09xDPEo4DJ5wxWv+eDPEh2qjGE0t+vzfR73pslKqaskqiJTXtvuePq9WFKSD
Jku/rd9cttWLJLziJFz1nDTg/3c32+WsIhIQflbMlEbISv7oeI7qegrthX1TGNcm4sdc7s6wVM0k
uS+gXDam3Vb7P6Br0qjDL4e+CaaPIafyYWkfCJ5qFuY3A/H+e2vQ9TGvRTCD49mGfxRgmmYb+29c
zEPoOVaoWtOQ3KwBqY1+WLScrrRpx/nw37d5DamKpU/fCY5aB3x55oqDoTJ3rzplQpnRRPJJeBL/
nLlC8eY1J3CV5ntQopsrUxnM5EvrONLbw+NAh4oq4S1Mg/HO/QzJ1T/mf//xl3pgfk3law1OVEIe
FFeTgcRgx2Pnkko/S3X4c6lTwn0To7IyAHlqPsj87MnR0zzLLoW/HpsNdmy8wPmw/rO5OueCr6cT
Yc6G7RjNnCItI41X2SHRW11QlGb3w6LjBNkJRfsxQKpeG0UUQwhkIrQemWZZ0k7Z+t8Ql2g9P0U1
hix25wmTnyiFAM0vX9zA7Qy3mu0iXP/0Abw8yV1S/SN4amySF4LzZr7c26XO1UPFD46VeYLJvwFl
xHDRx5BOineE3+/guRRFOmDGccYs0zua5h+HeWjbmFkAvqsPl520ShWdyEsXjlqUmJXiBYVXEQP5
LFdjdCBvhdugTm4ejl2OryxbN8qS+PAxry2Ykwn8RumgSdRNbLUCRQxv1zMaV7Qfz6anaegln/ud
vYFmAva+IP6WLrHRJY1ppDGvyTC37Krfe4A2puI93AagG9sHSeYjCq389KRoYolNrc6hsZj0MD3y
KxSHRnbYhBkwPNcviMLm+3P+okGBZ/VjqskEIfK+TQvZx/Co44RTYn3tlVsWii/oRjowFRvLg6o1
UjYJvYBI7YT/YhTOILFWFf2zcm83qWtW8zj8Tfv5SeSTr4zN7nFLProolg+rSed/+vSh1KQlzEgE
5RXp3+yluTg9gEHFeZ1JjQc2EKUTw1cpBJbmUga59VVopBgS3lEnN0W2caUGXU/WaJ4UkiqZn42Z
JIQEaRfzRfHuHTOfWDWyrZPZVW9JIou1MFykGqWW1y2KjnE10J9g9k0IVvBvcWBzszH+jONiE4Aq
7PSpIrs34/MGYPBIcL7Uc9gh8ORo2yfdNwqRDsstkeLb/zpfsmPBIYih1LGohiBCq8nUhOsRAnkN
ocn45awhma3h1q2nvJS7u3QTGayCwhUYfxZvBPqjNa9+Lutme5OmikG5iBzt9JvEd5Pga1pS1EOq
w/hsU8gLwNEgV5Er5AerpYOjzdLhbgBRjZiYQYcv6+LgjDrVzrfzcglzQ15zEjQQk1BQI77qjdGa
Ns/el99/KnQbW/qLiZPEb5c/luuSXpgFw1m6qF216P8FHPwCQjnjYS6HLOJE+18BkCjyJ+QFj3Dz
OtzOsJX9zPA2rvOeWRiHZFH2KGaU/LJuPm5VTMyQgTH/ENYUqs52ZGEm1e0RqfBm70FaryCCQd8z
nPn2ZVS0WWh8kyeQ7LmvAibtx7mmjaLzJ7O64jfZvLOk8wv/KP+m6LxSpZ37yagaUfm0oRQRwnDJ
Ei/lgA0FZtevepsCL8NjGP/B73fo/OCZOBmQRzCUBYCeqRtFykq9IacQrJBabpB3ouePEfStmu3P
8zNZJ82iM++jo6jS7L6hq6FjRLVj+a2gYvE4amOsZ1W04bCJDE4w1BUpleAs81gbxFG5YMc5mrDp
lH3Bh+d8o/Gik2PTn1JLFOdPPs8kjSoubR0ibzpS/vKWpxWcb4H8PrlvvpWNHlAyKjEGuechjRjr
K5UIP5ugGiPLX8//OzKq8Y0A+zUZCtvJCNeSq80oiKTfJZaIPJQxivKYywxsXuSxLaJiexk7Gy6E
WNUp3xiuri44qJXJvHr7aZ6E3LTViiYQ7ICR8EbDLm2NmsdgULCxS/TRqpfLkiQU3HRLclxdTMXB
0bw94aSHc6t0mxld4zra9YpCgQlh3WGmJNh+qRNm8p6tBcIn0jUpUDz2b15o34K4VgsWdDb/nRzh
N7DyTqGpwOlJMK5A/H3BvFmnwvjihfl0td3U3soSgjdxWVHSzNyUD1DvWZyAeicDCmbHuA/yMrOn
hqHOo6wKZvOMxBinJTWalM5ExS+Za1LFSs/oQk1Zw8erXI6BTnYmA550IsfebjV8gIA0ZtPKqYsy
DHeEnJYiGn4+r73XL4C/SRD5mB1tKofOubI/BXKQ+zaRZYIA0BWxt+x2XahH7hO8stD1RIJcbUMM
MfV9GZMqiBYAwuYchZT+l6dvw0G9/o+NsH//eKGUwwY8TS2XwckQ71g43DJmXnfwJK3lDUlO9YPy
RX85j3I5E94xTX3rCSqf6k1Yal/OUFPuCt+NMQD/5KFMv42940xKLCfiXvEGeUXnK+v7pwve52FM
/3/Aj6wwf2EZpQt4dELMVe51tzD76RcZcZBl+/i7tUgKsO+bmacctzXPNsrszY/ihXAdRpCZ0eXE
Fo2Yw0mU2Xo4EAzMbbPwz4CFMmnZlKTEf2GzydJ7MOpeTTRB0jB17TD8h2kPFn5ggFS2OZrNLvuc
8ESt+V8li/W/QvKiI4A9Od7NOhPwPyFtkKrx/Fu3Z++rcmFBS9CwFt9ke9Z08AP5LPeaekKKqkmn
sosCr7WScTV+txWDL+ALXk1I8GmEtuyRfuJSzi/0+tcdb8Ftqb4dgWn7lULZnFWb1xVGWfEDBLXh
iXxyfqrlW7JwWHSlu9/aMGI52YZTlzHPTJS7rE+2e/eIvZUj3vNQuLReGhlyCYATdEoodC6e7Lhq
HWARkBsSRGzURqHQsvtWL4m5xEwsB/qW8Sd0UOn5qFdv9W/Tzf0+EnqZy4l4ktP61CrqYCYePvmi
JjMDHJu8JJY/lh93mL1ZFyb5Mq4f1s9RuaHQOuPXv4yHTdr2+UiZopPvsmYjTvFEwtaae8f5Xt+6
49ETF9gWFCJj+lmnJa+0XNeTrDWBWBFKGQwwxx0tyg7dD1c03iYuFb+O0CyYJpsRtOMD1cU++FDv
wkfv5CBALUp5zIAKihpj7VH1B+uPrS0yDTsjnyo5/x9iR/n2V5FaCfV9iuiuZJX6GcXVt+hH7PXl
HHAbdr4K5JSlv81uB86WFlC0VTBwwbX1mDAzJxaIHyBxYBIUCCqypBBNeoKBq0cvthDoX1mY4efW
iqiEksjFZ54K+vk/CSdi9Lw0j5DcqswiggoxTRO3chg83GAGFafJkCpGeU+eM6tk5wapb7Qpn4oT
89HLdRsN0qfvq6tXCdf0ECABoBg++Xg3vrvrnm7IHt2L+eq2Xff/uPfHG/Ml1MzUbwInw4s8bLgD
sPK/rmh00J+YI/JQEj9pylqMjm+EustE3nee3Zs4fcp/XbSpGtASbSk4YWwrDl6f3mXmTLr+eVX9
I6oA1ez4aUQt/lGAtAgW6khu5TOd50X/K975GsGyz3/kqHUSlHgFmgYY9jD6XT1Y9xj4Qez4pFNU
wYR88Ho0Lr22bOYQRKGYNgil4mKqWk9LnS1+EeeiUnQxcvHeOcZERa1kpqUhSGZmx7lOMztEVV9E
YJumNE4Afc+4QG8RkTPeSYvyculbrhi4NTpJISzxON9EMGnfHjNUEYZ98tYoVE8r7ZBDnaTqiV/z
410dxbRb4arhZbTON5u81OjCvk9pqFxKwyxaWor/0Z7fNhk7fnB/fDdvJnhjV3CeiGg9Y1uuH+Dq
08+8wRbvzwU3gyuimSHq1YvIu92nGIBNFt/LqTJ4SorgnwMarRotKgR9XJQXcqJGythigv1smKnD
ELQXyrJvb4cuTvcJksGXLGqof+SFpkJBQIDbnh8kPCAByxRLW/YYDoUquWi8Psez29NwKhyFDrQA
I2ZOrdTGwgwNa8OLapBV4yQNlrmTII7XJbMxda/18uSuIqFZtp2qLHsRc4ahLRFVrkBuVjPwrKtV
Rda04P7JPW6KCrESyvTeEXJqRCaUvlWJObjkwrPVqYkgnIWcPvHQd1Dnr9hBr80qOPfLfetnBQTJ
Mm9d6lOMLsb+00RzHGcXUw0UlJdwrnhRGOQgt/tHYkRUxtXmtU45WlWzqG/U4crQ0xF8qlARx4UI
YKRjAO7f++/Lk0/o5cevAZ75OBMJWaKR5qz0Rsj/2wFO5P7gXhq+4Skxm6yS2jPQEnDt93gWlL/6
QeLxMb5ZVG4p6CR/wQXl299tBL6frWWNcYwVh/a7FvxKe8sEZy5yCDS6ul8dPqle/vpXqdMYnJ9n
cNrzDX5tFopVT/MHl5tzHB3AtSo6/y/T78SkZRYXz3KeG0eQyhlvYfWP0R8xCHezQfPaoe0lbyZT
2a5zKMRrUf7899kLx8vSlrNO7wPaAbrvf0Z+lnHEHNWnxKZmEIckKb85a+l4e0kkHqSCX+QhKeyJ
a2DAKObPuJfLTNqJ0WnKHDmETmJHakMyG3Tk1u69geQxkTUf41wz3vACqrGxkH0RbHGMy1yF6W6D
PCj6awNLlp/izg55vOFfPH/UcMCLXS4N/hQg4Ka/5Ki228pCGRU83MG1VoXGNnMmudf1I7/fqjDE
KHkNTeBod3ruKq5YZ3cyQGx/gG9h63L0oUn3kAeOGMkBSrLAmaO7Z+7G48XZZH1GKGCJw8Ed93dB
jrFjvya9jVrkmTqbuv0udIScgJuFgt2YLdxLEGdpSxavS3tWWQM+qbkYV7YMbM0vVts3Tqirur0K
/M2Dpm2XwvomDAkHGnWwbi2FhMnhddYNqwDLFoj8hAKqX6NA+3bgy0tJOmD3kzCQaanu5ryjGEPP
MvnD2cBGnCwD2K9PLQqparvJriOWAhUS7I540bWvUbzI1N/HgcIcUY3R3Nlycj8aPOVq6D3l2LSX
cC/NbYo5oXPgzvwK++aZQM0SacU8sn3pWqT/RtySvAygi8jdsZo7E7KsssiwhuQDEelK1+sfiedZ
GOHjmnYQINad/NiTzK4PwOp7nNblU5TEvziP8hMAVhpORLEdoAETi5gxij3pteAYbSxpEElsdhBk
XCN7DQxuxdWOoGShLGD+Mh/k1GGs/CtBsSAUfb5vlUbyLCu0QZ0WyaMDvGHkfXuFZdA9b9d/9BXM
QLpa3dsl2ydo/+tlyyDZCzyanofve8pPvmcTLEyR+PV3EG0txyTrdnkRvSTHUs03VGiGuiMQA9rH
saAPCE/gss84+4U7tPNr3KmVRHE3W4fd4BLW6kQcZSJoahRSz8c6zoxelRwgvl0Stut1IL7G0Y+W
5cYcIlNdjJq84EMD7PS9yZY4s8HRfULJ2F5b8YRgdQaipdXc8U5HWyjdyT02k3aASXPbj7scwB6L
kcl93cM+uiRMMIFKlBc2ev39SABDHaWVH7YRVvpVVAwSXvq8K2To2/oCqNv37o1blV4jsNx4BuYU
AfrHrzsAMQlb+M4aujFhlhXFLP16jxs1mEPED7yRH6RwFh4UhEsPtlpcurjq2khKp8Ys+ncQbJee
mToP5jqWEyPs7J0YBMwLRE7t4JvlJ0JNME8x7e2Y+6NZoQoFdfMkCe7zQiFGkEMLU4FlAk7mqKt0
tEAgLjlxOt/axC3f+hc9+E/vtPXyR8GH+3taDOx+pFBIltr49Vp37JdhIaKX5igwhpJ9N2XXjyoY
On74a7GYnxSbqmXLbQXf7taGlu12HcUHjqGIa2PODXIe0BEOggwsy1B9glGA4q9aqV9gC8y14ZEv
ONP3E4xelMxOtwlvvb/3nStPElt//X0/kYAgFWszkr13pJbuSc9WdFosA9rG4SAK0CnI+rcjkYWA
lyFZ23iDFCK3fBDZQ8jEmKa2yJyH93gLRxl3t24GzpJdy8PZunEti43fqLbg445r6BU6K+uOt85H
cEGf/H4wpmKDdr8NwTEo7YqKq0ALVhiuQH5G9+msXRyIDSzZVWncbfPHDd5U404PnXPCLwGFT9lP
p//eY/AosWkACIy1MxBX4U8jM1M0VBxUDn7tsygVDZUWUnVHC5sd1yEX8ORe1zFnPriuMH5zFEjv
NwOSJh5rAvWq5I9UsONNd+3ubFUdrJKyppki7dP+Vc/8B/0RYVAMf4VuaTQ5uqOkDVX1koN5AJdO
G2CSU+MzhPPg59lLR18B+eEUeD6yv2BUrMTmZUtrxr5dZy1rzyPF+1DPcUTqZxeUy72xFLdyLkT/
JgTg4G2EAnoWeh4Rd1UjmKiWssR3AwDeEpaCQ4Q49DTIlOL0FpWH+ug5HIYBjKOv+9pOiGHTGYX9
ZNk7UPHaeMAXCfMxcx1VjHR6cIdg4M6o6kLsVHQegE6GOETa+o7L5DkVbTvRUTIP63llOyK1KDCc
08zCBQ+1MWaOMh3MOU/HTgEcYZvVLEUJPCx5G+iHDn2tT3jePpgZFNkIfOUtFfkmin3gzHRvgtyJ
7EpkGRiICTm1JuEyMpbylkB4b0u/uhQJqbc4qJLaGP5EAn3QwNpoovB1/SDf/NpI1TuxDU3df4C3
NT+mVW7w/91Zsv4+1vtm0U3OZmqAJuubm0xfhUQA6+IwtotfMWHVeVQJGatK+811WUoViaVK1pRP
9w6yr+iNqCZV18yLnLqOG0TVRQaQxlgY5MoN8F0ud32CBI/h36Ey/e+0Aws9NUn2x4oA/5EdwU7b
0YuYUOP5YLzt98o2uDsczrqrXHpEBi5cbTegXwVbQLXEyLqbBZ3RQRSybL2LKCbbIBebBdfwA22N
Ftamsjri8/GZOy5TiI1s1Beh1BRbxEaZGcNuBa5/3QT0bijG1LIWK8gIFZBB0MvUKKNWV5glE+Xi
E1RRqzkcZS0mppH3uzyypWt9NbfwtbHJebB37o1qZtjR30qFha0V9r1pyuKpVG+b//alB13Pg3p9
WiLY/5+6UqjwG3xMTN5pNjvUc4v/hGNFwd2D+ZPgAjQRMySop8XKUWvY4n3s/QTv5IBxe5lXXjyF
AXUYKYF9Q9xQ5RdNCL84Gq2apDrh8MxdOjSOZGjEvv4bCf6m44ud7pZX5DBc55ibUaTGjVNXlDuZ
jIFyhUWysHnxarzgF8gJTRpA+B6cQmK8CIi9bJZfHFA6GvIbia0APeK41l+dNzPN+KszF0DKQJLg
cfzZJKfpGFhBDz3epR1pmjiqm+/31W4WXv7W+DASFdHJAPEK57Hjoyk02JWzL6JDKz4MRbdB2poO
YSxFhTcHNqfPQsoCZUCMpwJfVWM7lPoB/pJPu/mNIt4TQ5o0QVgFawHiDptzuyYhzI/PmXsbmJ5G
O1DFVvbGG/aXYRb5L/4ZNB+LcG3uJfomm/7RNVidTVHJuxH5osnJazGWqpTDtvQGj4da5vAJZCVJ
nV8vcaEwzjv0Y6ZxVPtaADqa9EeWHukLbVd4lstCCgNXqOvQnr1We47IFfYv1qTP+dpcMUttyN+/
0IFPXLj7JrGoAZNqNX+yL8R3+M3DIMiE+hqLGjk43i8oxYteEMqGTHyLoN5urwfWCuZyCAe4/efQ
SqMnonX9ss+6ZxNqHyOZoj+H68h3SCj1O7+0TiJt5P3cKgXbH4dJWd+AGrfPbvPOJkICGcU1LgNM
2n8hLhXQdeGa3hymuZ1NSYAMdN9d6QQUta+b4FGbn1dDmlD9m6PCY7vGnnLsKaVryYdZ0Enmj8/C
mySNQmoO1+wscso4o9ulqDKPNChHVKdT8HVf87/l1Oaee7a8dfXVHKxygUgaeBgH5h451Wr8G8bK
M8Ue1cJDtdyfZjBIUqQwKXAjSl3VhExVGw6UmORZNSelegf2HeII3xtGbLQQo2oM42J/DSOfONGa
2o/6396dUCTY+RBCahBqfRk9Vz5mvCOHo7ZZo3/Yy5zUfUTnfTtOq84mCKUH50iYsoyOnscSM01I
bkAVjqhGafrnjAXO9XT2rL2YGpkK9HjSRGAy6DgcmJsDW3P9LgfFan4L4Cv7uo0hQpmARzqNLAK4
ljY3DkXUB3/q1RR+R6/LnnthxFC4Z6M+eYQQzejQsdztb/FiQVqF52kAKxJGXf1p10zigZusJVHo
bAN5pldkBNGC5eRpBSI6YDXmms+tNKXZdyvaeojWook30w1Nty2onRKCTJKff/LGs6Lgct4pC/iY
glBDi/9RcmkpUAtW73U78TipqUD8vkKx1d0s/wl6PDio+fNXy063WWqBWAQFVBX0IQBni+ccwvwl
pr/UtEWCh7WZapIlaEbaeGhrZKKqHfexL1n7WVnYticDk1xuPc4QqvtvqyXGqt+3gIns3xzCcPZu
LGmPbtv9oBNyyselTrOs91F9xpXoiYs8xNzMOfRjzsQU1BoVPMTeVGHlBwIDs7WipC1kNrj3ukgS
mGLtStJGic1krevcwqyC9+y7TQFDkwvZXZT7aTKOsjxuboIctUrMVrM8rerwDdxxv/vvFQgW6SyN
jPQYOrwDZIXCId5yu1tKCXCOC1tvzWcAMFkSrydjZdmzJZGp94bdJ+QMQ0exZEh0zf/5v5jWD/Bl
MONbJRauE+RrAhQHQ3GCxUmQ5iso3dCBpgZg+oJoHR6y7UQo7fVmyWUJOtFgxCrhwaadWLaBAew7
7FqmPNr1QJ00LWdiEykZc/J1QXmsZ1hjSIf5NtEMT+YuIcLZEm2i0bADVQd8ZDkQKsRiSLJCTcK9
IeKM/YCV1vZ2rpCObtwAHKKrpnT10DbdegdhBm7Wvi5rusvuGFzedWqj7MnnUto4lZEfNs4nqCmV
6hoQzOX9iOyzp7h1EwjsveP77pSu0lFtJAREbnLpCCSrAcGcwXC4EAJ4gF0NIccQhDGfFkiXApjn
RkVRmlB9qByYOA/1Kk/40aqXSJKCovJlMPNUSRSy7f0nQNpcqy7oQiT3Og87ngocjwHIA+B4AqCB
VHv95M4BIfOJ75Ek9cPbVbd6GAiJFFxWG9U3Uo6qXTsCAPmTmzOAig0UsD96KkzMLNG0t+O9sI+d
uvJ0knE4WlQ31gvMC4K91h3rCVEbwFZo/+2a9Ct57PWrr6KQtxFNDA1RuNKmpEPi1aKe6x+TRevS
FALw6vfuxr4VilT0iUY5suVM+pf55QBvX8xWgnGyyYCRrPN28OKkoIuUMeyLbDI5yT4bjkcVcCem
KcS88G5MNwD00I8MBEgKKgbkbKQjgFR4pI6A2/ifd/SPLM7e23u2f7C/e41BDqApw5fdg0CyCMbq
/gXVYHg04jOB1Ypetc7SaGs2UvTTsFz+xoNW5ay7XMsHypCJhQpCEB4H4ovyTSDSTgJAktdyQNHR
bGCwNc5UWSrDteb8Ka5MVIorf4b7O+55Xg18ypNrzPDO+IRUybSMqlP6H3I6tKcgpzJC5FMiCqMM
pc211z9Nqo5awkfomftm1gQHECkxUyG7YUbhB3fKX0TqDpZwG1tqsugnXd/+DJI5MCF+f9Orltr9
FGUDnLjg/GadcKvhsE++/n6pL/pZWp902ZzLQDDgK3KmKubY7rMzHLgQLd8dw3v771wfVoLv79gL
+QVRI1pmnyn66B+x5Ew5vlhnlj0UY9CaXL9iMLmC1+HKs7Ax2zG+m21A0Td6Gvi2Vodwy3RfP2ma
GV/+quzcd0iuJnZD4PlQ48+FAGNQslc9+ZoLXaJZcEimYR4U8PMr7fbgrt7DwMS05h9jppvG5toJ
vsaX5ndfn0gF3iBPMITIF2F51D6ugs5GogWk4QKlgHP1rx606gK4ZJoejkThbg3ynHPPNH+NgemZ
gDGvgpkKK78XrFk3u2DK8GsUp+ZIjFaKb38n3A9cIIdCWR/eWuNZa7TReuI3f13LstMY8GeJHN0n
NIzYstyO1qzoNv8HvMx98aMNvTpAou1JO8XVroGVYAaIZdkLar1oqmqL+KLDrehSJmmuTACyCx9u
uNkTXjTyhRkMIGaqe2l46OC9wf3r6MhIwLr3zMj2rS96zHt4Fa5yHmLL5Z6KQYzzI0HzPaAbVwYK
lEWy4sObBvMU0RA0a8DEqsehY4dfHHykzlai93u4uLOJ5q1qErXNghAzbaRmVf1/eswrfzfOaYCA
FERbgAOzuCrarEU9a42A0pBpa8BRQW10/uIk5kTNRPFrrNoi4n4VfUKJTdoOLFGsqHg4dqhPFiE7
4bAdAJZCbkw3ncuNHvKs9VJwJduSY6cH9LUe5HTDxUEeugGqIo+BA84AechAjEUfK6/Go4cmMcVZ
glt0p8v0j5+YO8mEzEPQl0ly+TJBsOGOsG5VeDHAq3l8bby/avETnUfT1+b+hMZi84Gygfii8qT/
yh0wavRqJZMcHUekYCmKfCBCnaVVw8zkkC8QmoZL0jTJV9cS2uUEDNz1K4I14Gvol6L/C0qRsjir
vdXsrFtQEzSladStH4MUKyuCF5VOuWitFcKpf5/3fbNd9DTyQaqNmqvT/9OpSTYX82IE0Z6zw0mE
OMyICSfAPRmZOpokRqqBCDkAe5SmmrhjtV30FqHPKs8XfFz0VsroUiN1+1maG4ZBHzoH6mlLkX+C
bp+VPN6rejYshYAxXQSHlQ9/aJVywHKEdMjxOEWBnj0eEQ3tgZAmsdK+oQJ1wUcAVGhZGxWViIAv
UasJ8N2iq8OKZ5yk6HANtA4+k9/lx9+mH9RW3gi5cvr2tcJOgfeH2Xkxr92k4NRatSIC3fYm501O
1TKIksE1kGQ8KzhIRVCyBOXTxp/FJ/UZSYdsMLVWJGtbWvdYpaTfQcZ90qQ2Ghoqk9PxaG4NnE7p
3yNcr63XihLdZO81iYHRJOX/AriqK1/u7F7xqOxrQ/wtjLRsxU8raDoTT029CD3Ok2DTUAI6whY0
Vabo7ncJuDRKzpI9wmxSk1qGHi6/6tn7uEzbvjrVySfRopV/bxRJEna5C8kNNp6a6CgycrHESKRI
dRmGgXyrbzVLkkMoC03cuRoL3VBhpLJ5QNhnaOkEJ8coRPnB6P1BrSXjHKuxFxQsDQawVPbPyq6L
VrdHI2WhbRINYrZ6RnbzRHw8m7BdomOUerx1cE5YWWw8hx8WQm3kQqHBTZStWSG2FORXABOxi22S
d4f3150IOPD8CLKiqAvDBQC2RJvKW5rjV4GOy4sy7ALcPIYAn9cfXs2S6iZL/22uOBs38VsDCyC7
GvVZHYKVxcWxo7p8l3csoG/pTKmEjMUNuU66EOilUH+ularKIlv7+HBzBbLbnO7EQAJamwK+90WN
KRyUoOtluUwHyn2+szTMvn9Zl77xyuwBpmzJ10Dm1YddZtFd4kWvTw/TubA5JK8dPd786hKatXVQ
NOARPgsNP5gpk90bOb1GCx5BENeAnNZPOe5mGJ5nKKI4+jPcR/szExcpKmesXVpn/pxY51O6BW7d
jO2vsZliFBCpJ0lmpIhOJ3ty6ADdsN89pO8wO8xZsDdhF0pSiYSrW+qWwj7EOCWyJBVH7Ri6dtHP
XwdWaRp2rRzwNfl5+kMKUIk8mXcNyVTBNQHrERdBjrGzZfSaBO8q6wd7lYUn42uuFAPE8nz4/HM5
cPSHpL3xRbcwNUowkffBcfthSaC7g833hwL+XBezNpQmDMLzBPnQedowFtl+bKAzEWW4aCEamFAL
SY0Itk3bA93TB3YUdjpI8Oy308wd0hRYctgLmhnK5C980/uLpPbfF/Dxoc2Esvk/ImvYL32OYzEo
/xhDR30ZQKDnxcJlSiJM5K/QwcU5NWSfe2fahb1zFow+UqQh3W2SG/tZ2x5CJ8fM4xD3q+DsJor+
qrMq1eRg7802feJvKAlw9wrE0yPfydn0UhdGCP06FewVXVe5AuIzRciHCpgCT+BpqOitfd3kYEit
tnYO8I4MRtJWNGY4fxmH9e2AUD/QZBDupZBYPAWMwz1R0IqmqysQ51gEbeIuTfU07IEAAJwq64WT
ZVeMBPXvI4XB8Xks2FQkzIZr1p+3hiriFm7Ck1BTbr0NQ3bPjVQilCSB7RUWeTvRwH2mlgVNf6ex
NDvbcejt0TMkMRnQWi6i5V6bwAGlTI3hg+bvXhLjm+SQa6V1EZu2ZovpxCIRTqx49QRN28yckRcM
9cAtpBPWJWew2ajqzBlFQ4/GmyHPNfTJGAE4XtspwWFuDlkE7TAe/ZsXF2GKSIXV63CJvxCOIQ09
7L5jTcQM/2ZdSCo6nX1BFjOIuercLeofsyzHgCq5IhcqwW5A0zZMNUzj+sBzQUCjvXI3K2CKWfQk
7ys/mwI+Es6ZxE2AtLSNcLFyW6VFK+ZMMTKiKSJnVKwO/MpifkLA9gxENc2HH8ws/mqZHHdEifbN
mwC/JgzN6tPUfi/ZEzsyLJqbIAtEaAdnpmPEBUVKIvItXH31Ru0M7OjtixOPcLVUo4+NYiWc4ZOH
nt/oUzMsTrJhNNVCrWF74F064vxVziZgAiaNTyyWDxwvXQFKFM6CDnnY7Pg1wZ9mfJUzvteOGUS9
RmmYVaQpiUxrNZ7za2JGNqFKdO77SBxivshBT1PNm2x7v1Scs23VbAQv6CBnO9Yk9HjNrFIfWwgZ
vXV4Skw9PTAn8Heklpi7083tOapQC5A0Hc61SbLCKOelBlz68V8lHGe7F0sSlWqTs9VdVF7hS2Ay
yyJ9WrLefCvBLM4mupxliJg4olKNcBksRMCocBzdGweanyjV1ZuXThArwFZw9JxdtHTDd7aNCwH0
H6rJl4GRL53xXQuZqOVwi2Ho7kQxmILOoIUhKRB0ElxEeZn3NHR7LbFWdjr6O+GPu9ivXsWe/3yC
6nm0gTeXqUKeGvmt/Y/MClSt8dxavetH/FKoUthvUyLjaaOr6DLOdTyT2fclu3vt1XezRATcEast
Sn0zwbPabAA50QaJ1FRWwQh///u0GyCsyjfOmrS+ltO7rJrMRQ+LwUgiwc862MlDA0NeSV2lP5F4
x/dfVYmlyKHSqF0xy/pJCVhlM1FhxeBR1+H7kccyKecARW4Nuyd47/SNcVT3fYgl9KCRRnRdnRZy
OBBLSN+vB7ohbWIUHP/YZpNTHvVm9sB/EShJgyPwdWk81Bapt7NcyOhutwzln79Kf6R4Y6NypZgL
81rT+0Y4Dbt9zUNq0HQ9Z8whzNhAZO1sjUwJxgDX89nPecY6K+n7FngzTxe8IH2eUrUTOSPrDQAI
71mxAChOJy0RWVwdYkx5hN91aF/S0wc7aXTKp62qillxNmaGeo7+HdoN+EZeNMeG2yYZH4fXZVXQ
n1RQR/oDCV4jxk2LPCJgIVcngDLg1qgFOtNrGujHQb2KLv+8nbznZkN7cQI5mAoak4FWuxj1jEv8
boGXQe+o9j4aMTv9+5P7/uZz7nWPIhKMFJQ7bn6XDvIe8YGec9foksmtcgJhhl/jzLtM4yt9pYtw
a3yL7GOSHvLxRWLVt5HuDQEwmDAq/gUHt6Gm72Fa2qoZIXI3fVXYfQ+uQnrxmNOODibs7yQc+I8W
UumYJXDB9NtzdJsa8st7idnql4ONjttTvIaK5+4cRNWQoRtGv/qSpwWJxOQMExEita9gl8vQyst6
WRJFKIHDyGTILR/Txnr9KegZPOxqYVoaKSptVS/0Wqy1QkW/MWO5T4GjmworB7qGbKNZ6GNT7sXC
6zyW8tfv2qNBWb/5RV8muYFD0IUVVLF+H/IY8T+g7xtz19qdnr7Q3xmnYYWwxaeIREEDkBYUTpln
57QcNIx6hz6cJoW9VQlSyStickyMCGUdG9LXTYVYAIiycT5FRBjtTPYvBPf/BPXJAHFeo4JPr8Ru
RLtV1Vv0VcT9ezxlFfnwDrxa9s1m4G54cBlA5Oaz6JwwTks6Z99uDTHBXZ9uVuwJrvrFvWQGgCZ/
LL6Gyf/ljy19mTg2fPzy24lRK0V5LzWlzAtA+HZW8bQ9wGJE/lXx6OjZJvZX0t1+oHhb5NU0bPbU
bSah6R21i5X88nXtivGwI8Fdncdn5BMxuSMY+/pa/lecYxt8f4Sy5lmqDTUhW4lnqIlwAgJCzOg0
ZIrpgnnmYm9RzIEJ3xGPeWhvXI46DlAAXzIEEJXp7PPQCNnFWau0rCyixveKew0ATL27J9ic2T0w
cpTU2s8XT9jvzNy6amFRQeUUWEmDB/fenfne4H1dWbJKR4fhNe3/g4dYz2S0lcf4HIip7LI3xZEI
8BuDWLW5qr3XyBNYaY99OonSu0b+zwNta/0OIwGuwacazDlyZFYQlrvZwzG79IXSHG9rqZkf6ela
FAwnD8y4FJRbmysbCMxG3lGaFszIHFK08LEyCbfK8h65f0la7vNiit8HpgQ8A1a2BsDWHZ5Dmt40
6uN0b1naSpx7aacAN15C6H4vSuD1RPUZrq7LzYZ65plcD929QlCrcTA37F3iv53SJ6zbnSq1FYmC
Ul1dDiBadELZsH/SRJ8JsZ5ftyNKQYL6ZCU5bGxb5Y9hlWHhoN2aSOInXp/VbWAM3hNCHzAzOqHg
8tiL7iK4544FoO6xSqlZbp0sjwsVRmzjDvlKnJubnD9d4dR6FmOu9I37weUGD0kKoBWWjKSyc3Q1
MO2JfyJ0csCvZKyrgpyzOik8LkO3IqQBYkG6pv7YwFKWG6dl41R0e1d2E6H041ZAv8EKs61sfpGM
/ByLVOgR79KoymY+nK/JSH6jpbAbl+Ejy7gESg4bVMMuKPJlhH/Bv4c4ihXjdgiajvk6qGy4aarX
d2oIKVutzhN1C6HVNssgeScc6LBdwNc72T6SLNKHLQTBfBdBuXDHOXjTmTcg4PqwInteu/74+e+o
smb71aUqTQ6ixjlOjznoCREF6yWef8qkI+EBdlO4//Cfg5ovZzCw06IGQwQFw37MJwzjFDh9OqXs
eDhQ50izPR1abpU0DyxwN4rlGX2F2RC7ECrk8MrV5LIo9BFzdCWKs8PTxsI6y1lS001qhA6SLsfd
aCak26oxOs6DAzsdgNpFnkex650jqAXuQjsw+QoHacZ4a1z+Wl7lZdInIL93ywLhiIHy3+rSJoqq
mCtoofOD55cI2mfb0WnUR7Ne4ge3U/4f8AWpunR/ppDJbO7UwVjld7gT0gt8IVzGGeSCjL/VzinX
7pPUJ/bwPqrtZpo4cFqTCzzzDUfviHbLs5S1rmk/+ywGSeWR5SZXTU3UxrS/B8Ch6905UuEngH6b
y/OUqL+Jf8QkCH6o5VtdJ88dqQGOcerkp5EyLyIaCoW0EUhusWPkV+3uZ6ae9my6ouWfuLNw7yvT
RZskNT5UNYfCksTD7sZxJU92u0g05nowa+NPd4rRRFwTj4gj6jBQLAaCsmmRKvz22rkCccncq4MZ
GgLxU+k3z30GqAv2hNk4aajECNyDm3lNkoJayJIt1c/QelmldeCpuCWw/TB5nSu1v4QleLGCQr+j
fTHujKPEolXt/LMyVBD0xVmiprUNL+OuyKCuqVKkqKzhXpR2Eo0UKl0Gvu8b8odGmvr3y4tnSDAw
eo1Kw3nRz5K4+QVfuLhphBxSypme2HQqpWxs8RuT4VJoBspmuMeeLNKlzvjqGHfU2CC+/9m0WALg
zBgMeE7T+jLs/uLFAblO5OCzGPYzS+O2KHIne38RN8Ut5pCr3IJ0lJh1ooGPNoIlbHDZF2wzK1lj
8WdloPBLUzmhISzp0Nq/Khbuob+d2nX+6+fj5Kg1L7Ss7vSALQQvAuPF0vzo5URptAS4+X39MknT
ZgZo5Wio0ZxXsUZYvEqLZayeOk5Auz/X4cUhwVWFlcvMVqNwzLAdAmN/wiyTjSmyUUq7N6e9P4JL
BeE/kpVifK5xVeeFs1OtA6ywZmoIsRKZcK5/LgnLL1+PTRBvCcZ+pz9D7J/2zzHhsR94S2C9iN4H
eVvZjj8nwCAFJN+WKcnfnQZUttKYmGmzD8TSEBPyMZLx2WVkB3UovAoLkrXM1rpl2G0wuRQ07/dU
aJAGnWyYpkbsMt3XUSWDuw/oh7QGnvFZFW7TrSLTf3uRL7aOBx8+ahqX3xZ0SebP6ZuyWFcq0XAD
f2MYVuDfBIXuQbycB0H3Apt3dOJtW4mvfysB8ZAH6BXedTemT1pmx5A9iVvx9Rgr2i8+y/wz+/Ph
dIn7KowIfpqUGcUMpCfzQpQ60psSzHIQFuH44L+Z/xih9ZPkacIHjFOLpYcCGePC59kELxHUT1E+
f3yqXOB77DwGOPrtwj1QbvPyw0rvB80yRAjAcGDP/YWpMP0f6tticEmiu6/B+eEq8BzYliDGd91k
ZNqESkuqCDScLG+GTisb6OStSJRKhubcDIq1IE0vVv41F4RGIqkZPoFSu1BzNOR5veKPoZtfQhi+
lUUNgAbClVHqkhM99CujLHkdJY0RxjHIKpy0sEvIqgN35qpawUYcdIfP/nLD/wt5R5Q0j76APq6M
u/0Tp5ce/vj4EhcGgePyaGIRpdBd5l0JVvdNh9ljOcGXKGTsEkpmLR+brCS4LlvcK3abLMDzRuWq
B/IBqYM0z0Zht8ywpcpbL8MAHRork5VoLgC3hiLWlt4oSl0BruNTwheR0XjjRTiF2+sLryEdOyvl
sJ1Oz9tRyzDjbGAB6CCWoclXHlm23bTVZz5gleW3iBf6KDvy21UfSCaOipGRV5Ntpi+VXnzSShTI
6QmtfYT8T+eAsgQ3R9U85a3i33J/7fDtCbdDTnygY/sBiUyzYg4Osdw0eUzPgjLRcW5grNmIsa05
cruj+VFhQCkxWrTErlb+qG+3W1lPu3/tAaSUuFg1zLDyAzjMMG1fAqpryEAcYBIPqb1SkGX3hNTF
MAN8UMRNCQj+YNkV/ZOyrX5LskbU0M349UU6rbb7fAXIPn0qFsB45eFYDtDCx6znPiUytvqPc9Ph
WJu81GZ5ZLoq0dVHtqmBurgebf2y1/1rVJVPhjIWkI0v3oIjVguv+sSmZEZqLg0twaLsQDXkHrHZ
cUMSSAQONyi8mFkf64ewCT1dlsetUufxwew7tkztX23G8gaRdsvImki5WcnKH6GWgCVU90cbzgzv
L+yYjE7mXvSZdfVGQ03N3zRSTR7T9/ekjRnghJYRiFrvXgaIyITdfxyMWYTAMOBEFFY8W9Thh8yG
tVfh4tgQZXAnuJO/8EAzV1fYqeaDuRFGoseiImdYD628K2EtGm1erC+ZFtQXTBBrPp3fsLT1BbfS
+/cbK/b4mcyyUX3p1ikIj1HacpkNIPeANiVmeTfBVFsN73lDDI95vA3ryGi77U5YgEzHRBx8PLd5
axaxn4MVWfh/HGsHUG1WI6+4IxJsP8BoLm3yVjtqd7xzFSb6Ljsv0VBB9fTLEAWMqm+niOXsld8o
zx3LDpHPstMTrHfeTWUjBdxp3SbAkdPYC8zuux1dafrY94liZhIy6xOVlgvHCTEjE3JcMlH1xqAg
NTor/V8eKQZRHpZf/i5xF9tuJjalbMDRfN3U+A0PfbJ6RmywaUb2P3llu2QipRzJEXZFSlVGGe3+
DV063Ba5E7W4wgQdoxPcoengTwraL6/SjxUQ+shZ3bPMpg53ARRKKM2j4P7rpbDtbrip2FOXDFb7
+QjK1PFKi5I5vN+q18JVybyeHEbgMjW4YHkBlD1wwEpoAv3/cscVHeTu9gT1KpbhaEex47jLOXuc
wEllkcxTF6lokaUw0yjqf45M0DNVVIpvhdgTCVN2R3HDlQ71zl/SnqeKy+jbGq0m4pZW5Xb3fkfo
UcZ8Cuil7IQRgs/Y5nczkCwXwey/NepZfB9Qr1PIAd8DL+z9kjuXJmxFhCsy0K01wJ4qoIKAbhEN
cbp88AfGsFCczTz0SIWG+I3EI2Jsan79a1vDZFlkPza1qidEcQ6lEd6Tbhb5A1wvXuy1D11GW8rK
tJUlknIyph1hfPqhEt8TpU0CsNVUNb4Hvl8xPRTV2E/5bIcx9uTi5mHcvFP5xWjlgTnl+pQR91E4
WaisxfL69hjszAgqpNEsmQkNHc/yKocczgXsguT78fIXdrHaqTyF8Ly5V88R7sj8kD2guPsM5L5/
tGO0484PzJc6a/nqOpVlCHMTBKynCuPcpciLP0+aEn8o2nqlya27UNMM/G57G7VY5ECZutg4njZy
uu8acO8xQvYYkOyxEH84PHGly1bCWb7UAi0Xd4dYhvcZRZOEtdzrRIABYGfVyyHE3lnx7nr9R/ik
scJ0e2UAiKZ6nvVhjM9OYtgqYAu3B6YaPUoJPi+2ZVo9R+xLtC3v7SQMrtBeXFPDGqhf5b9SxOm/
lngwuLh7D2nYptvTaMXdTc2u/sKWkGZSdM9Uf6FHqgxJOU94U2kDVgPjEJ3hy14XXdRFOKYvnUbI
RjOKFTVmsBegp8BVVDmGVJywh5ZIsS2JWaWwtHePlaVBa6MNa8Uo1GszxJT7tOyBGzkFVY/IX3Dl
0qmPKI/LT2VkH8bSH+qhXHL6I6QrYyTO9MPTwFNyFpDyFfUF/oqIWo0NmQapYvwBOb6eqHK/XTVF
Hf5FV+4fujaT778rlhUBiPZ11KssMt1LIj3p9VOn+JDb5+X/L8lExAGlJfzLVT3kMRmbDem9zBPv
OThDDx9peowVaFeAucGteDFwIGpi4/2jik/OjCWd3ksi21qMgr5Kg479+/HM8Fj1xs0GLXUn+keJ
K+pYKumJLvdfkgVfD04VMRVPf/Y76EjUXAZS7j8NKppf4ZabvmG54PidP9jwy9Df534JijzeVvwn
7BSiGI+wRiThnQz4AC6ncoDG8mYc+MpKf7omSIa3EF0qZmMY2U+muLeqp+YpSLEioRkV6Gy3Neew
+5kTyTtEGLCH5Nn7HHlhBL4MRY1WiMoUsstgLDpZe3k7GQqmYTgnFB18E77GvfmQGVWMmDbeD6yX
aR6PaIld+jw/27Gqe2kKA17vn0H+94ZfpVBDe65SolNeE7ergU0i6W1l3WhGchI3rpIOoXUPDo1j
igtmI4zRFunj8jRIgE/pSTpTPNsnZMj8ycgozY27+TI+HHht08sycDY3tiFchdhVnq5FCBnwUxga
iSFZJ/Cu2ZuyLyitvAP339cKt1gyAOGWaJNnEdRspos7pnSBPwUaVU35CgD80TqJdW8pWeXz9sMm
OT31IdaC5bhi9k86f54ebjMsJmESvoKNP2HRffgKF4go0k8jpPd8tDEdkQkOBSl7bDZG2wFo6Keg
JE77TH0NLPYiDqUn03wrcf4gWWjuSM4cVNnwAGHQ4jPDDSBCAJwUmCFT22W/M1gKaZx2gSLmB2ay
GS9P4hfMz7RdUqFcHBTjudt68SOWkw3LXYINEODTyIIADzF7QInCDoE+9hFFoBDK4foe/CA/Y3W3
WHzFAk9y35xledWcoH3IrVLdiwsORVDzDft/az4x78Y/iR1mL74lQd7fc/x6RjAvMJJFyBbtsCEZ
2OifqLx4jx41Jd2qwghIHxrxUfuOZEZ6B0hFxe++mdPcTlJb1xy/bPNAc7OwS1XmAiyRGtpJzywb
mYwn8WYsMVUXJqf0c4YbZhr9W5ah316zORquDBHMZ2vXvnv/3q7MO2VR07kiE85w7z+AVI3rSdQv
KMjHANP/Y7Ojza26gWh0aQxgfW6DUtkbw7ji6Qdr+62CRKMiQYKJUInn1VGEvdrHD1DNhUb8fc93
wKsy2xHJCFjwEoTZ1XUxJgWnyOoU9ZMEBIpqEs94M6wB7+QKqpV+yS1tjaOZ94v88vQxgZWeXzDM
rl0JTyPxO1JSE+/l2PItGY+puVy8nEKevFwws8fE1HEomNdY6itpz/Pql0/9RYO7sk6EFDButBoE
wMY0U6ZHvapHGFFTFx3ISwhs+fsyPyu2DKa7S1OpVEPZD0XArNurfY9cGS+HUQTY2BYMKEJmcq5V
/DAb3kNf5I+QPt18qIqvar1tyRGrVFL/76ZgcQ3eQqxj0Ubba6sSlf26BaC5iPcp/V9Rd1GYF9cb
nEZd5H/G6FlO1wK5mSRcsYdOUMZfaMttEFX/IwbxSuJ21kBU2HO2knXoDPkihm5Q/opcneoROS3s
DlPGQR2RfZL1v/AP0PuEd85yZx5KOrsRh+PWz4asj9mCqQQiE2CFrkhhfSCAU0crS0Mt+dpCZC/d
iP+po1qGN2z/L0JbIqPISEg2OzJ8gBVDNkSsuus49gWbtEW2m7bGMxsJMfnGEA1KcHGYXRQ5N1CO
ixgXG6UU6sCgWxt4TTidHwEGMoClXDsuVdx/Y4vMfRQnXgr5Gg5V/Qu5aAhfPrtPmUSOuCslpKNR
+fI3BQKBpyioPtUbBXY6VQqIeg/5Y8kA6XcS/Rjm6P8ZOCSVHVLy9Hnw/cVXcpyhmyAK74Qf2A8K
1n97R9QU9x1bgeoSAy2G4FlhkhJQiomBpJksac0Z5U/UHUHdxNatwyhsye/SVpQFS5M2gwnjohOD
tDlgB6h6Yhsvv4Nsn3Fghl0KEkAklK9PKrL8oaBl6ODkocuzPk/SMgZgQ56QJ3OgEQ8sxR0AklBk
ssTKeT52XIWSzM3UNMW/W706l1kmTn/bEvJgxRGH0H1qYStIPlywXUs3RU9qaNJ2Z74RqfTe+yif
Tv0qokRtGAl/0JDjXrc+uq1Vk6sWC9OJASVLrO4JZLVwgNoZBbrqzdZNYSA9RohsyVejOkZGX3xm
ETAK00Fz6VPfbiFVPZiVNrrFIsUVZA5ynzvMUAh7TsCZyGj6BlDAiqIUKOQtVdDPJJCtpGw0xa9I
aL2zhBgryboBJ7u/u2WX2BuyGRVpSRQt9NNPT2uxEwV5LF/2nCQsfP+pk6ddho032sGtteaBL8Fq
VCIrzKpyNdCG0BzHdg4KF9D0miGz0KgkaW5WCO8pmugMDLBIHdieSUNbQhzMSqlcyN8cMgnxWkbK
i9YwRmmQJJkz6f4GsNzUxNOQ+Ipzvdf9a5f2+UwvlosWOzO+vF6cCWoVqaeqpKNTEgGXhoBmeAF9
4gHZVhJZc8k4SaOO6y7FWDx5eDn1lkjuccJ78EChEoU8TJootGteHRE916vVFR2rBfHRi8fqf6HG
egLfZpNL1YCDMF9CZ2cRCmrGoor8a5LtTsApMf+nPQfUXP9VMUVC0ZFVFcIfDWqFDFWnjNxNl0Y0
1J68kz+xN9mCxuX1uwmvyDg59TpMnISWjrryo7yfv6o0o0sARIOziyUwnUi92z/orlXiCcnzlFny
ILJ8+71qzP7UWfEzW/WGn3Bzgr145FSM7zVYr71yU+cgOmiWpRq1sKFsQzC/xk+hFwDj7GJ2oWop
iR1T3sP9Cf+zZhSP38sgLwqaBCbmcc6biolSxNq/3vT9iDjA0zZ1xTkEU+P+MgCl3cFACuau5Cpp
je/lIkHqXQvy2TblCuOJ/rPEOXtkQhFZzVuBKxJ5sbW88APMYUOWEoIlozI93nCUeb6lBEz3faHi
sahR+dJku5wJaiJRxa3mOaw2/t8HGik9/c7IvShgWenh3Rd0Nvf7oFUJfL+TrHtcMrPk5aym0Kj9
U7uHpvF/U8U7qmNtKt/Y4YRpU3Kg0AMXENa6BTAvT6FjzaNwDz+ydfoAzWuACodh7L4XvwdA9SQv
kBHkc10am1lxbl+zloe0G4ro2H4Bpbz7/0ziAqPcin6O6NvHC2sgl6ipZSb51pJ9izgSDUHZPAzj
oS5KRZGcu3TJ1HgDuR4Ee4K6qYfHETYvokXn4mOb93DUA5S0J2UzhdmXsOguQsH0Lv75Qrh/birE
3aIULWZNnNwrVeJNQHRkzPdBWRrWfPdAfHATGnXQ39Rt4PZpB7S02+bpsO3yRXzAw4klBPXg14Qo
858nk7F3nTC+TV2FZI5SkEbHCclyuHpyZeSTfHJSQuji3K6T+/Yz1mczLSJ1j5UMqIlouQz66PPN
HJdNPZJi8O37cLtohPVpmS07qN27f3y9p2uLcT0L9BWJ3HlY65kgyGWW2jUWlYEBKKXfJQqEcnSt
geacpGdcp4rbtiPz/ES63yDjWMB4qPsS5N69EA1Ix13wEem0YnIS126OZe1AbBLioO52962UNCIt
BQ0J1cbait7wZqRCpPWw6po9eZEAp7ZMh9/bw3B9Bfejv9cWuuBKMXCAeu35YFHZ
`protect end_protected
