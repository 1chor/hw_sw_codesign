-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
IhLg1EpWA8uIZB3qcNICr6w5aoirti/EKZdCiPpE7ALl+LidqtCx4fm0cISFtUES
vmwFBcLDwZOKnOQGaUmkEaE1aIJn6/P6q+m4svdTQJHRNX92ifY6wjY/SlvCwYvu
x8ehQy46jgUYz2NanmQePA5EOdwzqaXX62TTnIU1BlY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6624)
`protect data_block
4BLg8+gJJ7kAMKgerEd3H1wszW9kfZeYRuPTJWad9hLu5mis16VLVspymw21jhW/
3KjyvnfAhF2TZ8eDpoP4G8ud4gb1pd60q1eAwhfME8o7D+C4++sJhmWcKKvjraa+
dNWeMLXikyBQMIy21+O0JLyN/hJ1HmVvFzOCNSwOj/dl+DjfdZFF5Vh3mloatknE
G8LCdwgGACDHSlKXNUJteEpIE5MN//cYEEcMEkGRG7H3EoopJcLLAQ4MyAt7ZEc4
J2Lh2A2qXOukktP3J/OMYxyl5TlWkMxKOd5WVltAZKnI/BpgZLeh5T1weILyNxim
Vpl3/yMpVxAvCCU53LVm44e81bOmyo7qKiTluHns55qMUvAbUIetJmF2VLBP9HFG
2ZPdZ+E9RsWCjXCi1uky5C45ABTZIOtJky1BXbNgfW0UemOEc/tMqX58wXDNYXzL
q5VmTX7o7FHR8DmCsPI+robaGyT/9ptGEncvzv0T8CW3B/jMHgLZ/fTPIsuanLnr
c/IOcNZCzNhxMqS2CFx0rzpU4Stfdv17n+V+EqC5Y9HCV9qKnt0kcoS3lfCGSg/M
jlrdk0gYTfLrpv/wcHmE3Xn/YeE7QdKr7d2vm4StmZ/aExXH37IY7rHJe/SCQCbz
P4hMYuV+VP5l98mo5C+8Fdm0AHmkV0kQYUWUmxT2d3THfo7JKvzdHEgEbTBKsGsj
Xo3dHpQRoJUZrdkNuCISpgVI57Htl0RLm1mktFh8npFi2wXh6tIVtk5PCbiNyRDD
VaggDO/0yGH4yL2t+amz2bGFX6+17X9/n8uvDq20huyGQvqxENYR0cUA6VyImeJw
vpRKmf4bbJEx7zgPIQgjlGpiRdcuqED+xuJKRY4mSPh/2lAgmQvG0vlJpAokjlHK
dO5MKY9M1gMLoLxZgFGV6xrpe8BrQkQ+mRg0ouB1qRS/kX/yoAzy4rPAqtFVTypv
lUet896oSX6Kkwhnm5SFa81e/WVM2OR9K3/xgaM9KFseS5vB2MVZc8D6hq/r8vWr
/0SF0wutBAtqxnxeObSh82M1tyBxee/ThSasX+c1XqWHUU8ek5JFYB/dP6jiYfzS
yYhaC6fGdDSWBS4eg+JqQw+HOr00CsQ5Oj1MfingoqVW0zeReKJPL0hIxv7JNuY+
6eu/PwTznRKRM8xk+0AUUUP45UAdyyERKZOIJ+NfnMcGxO795FmbN7rYuoLiOQy7
x1eRAyKJf2Y4G37XormW+B/1/LrM6ND/Le6i9lsBi0F6S3YVOsPcRZ1UcmReZ1iP
wjyUeWFzdIiR9KugAsk14stHcHL51pVfYXWECr1ZAhIcoOh9tPr4cDiqEmwSwvYU
w76QuBz/rf9oAObeG5eLDxx23VpCblx0kGhKQaL8KhJvwokuzDtZf/G9OsSYl3OH
J4AQ12Ko+zGsfHsO6r/qz1O9pyi/xacsrdaf2F5LNXHN9CWrU5geM+n7WLsrEBVL
VmAbjl1/wKWKuF/SjrQ982AB6HCV9/AS6xeaq6UeO4k9K7nUMhP/n2RdRKGkLhqX
AXMV6QLj0krmHNaasCTUdXm/lDuEhRCmX1IHE1L4dahxh4OQGDtgblbRdbCDcldw
9PSU6KusNw9aXhPNKxRHxzBoS2+UkO1xSxrzwVhDYEKO/Q8DnrVtFc0RNhgeycwo
CJtC5LIybWnEZTSwK16hTkD77i1NGsvybA/Y/D6mDfLQaUJRg3+CqTtgFs+1LwJ7
i0ziOtz+lAeQ5PYCQGhLb27juIs8D+Kf4TmAVyc2Rzi5JmIompBKvuiNXHuMdaX6
qRpr+O28vqx0nKoeMOcjVSuAgfj5B1tdyiBU5l+HhvfwuvjdXc5oGsUHJ0UoBwQO
pyeBziAyuCCNdkW4I74ao0G3YrdCCildPsELXQom0VPoqwkLbZMr7e9p/g7lRMD9
7K+104PvTsYJm613h9c3p8JqtRUCsbiNdV4xHaqLNxu4HkRcAe3lbzZFiNgdekiU
porgnpVR6Wn+WRsBFMXvOvGMmcVAg95ZxSC14xRJbCgQ0DVK8eGloD6YNb9/Ze4T
p6EKMFm9wF/ajAMdwlJLpo9YfrvXnv7DIxTdChja+LcJzkRugKgRO0KqDVl9dH1E
muIO/Q/YFI0Vimd6KEda77Zl4ss+BpHeqUnB1/uI0sksTMvVQgSRenQrhoMe77FD
84MSHpa0cxMm8qkoucXwa7XX1lzfPjohc2obpYM3i37QjOVDvl41ceu/yeMHlljj
zCV4Wj9QyVMV3Py78Ii9s9H752Pk7XoXrYNhxjJvbH1h4m67+xkzcpW/8YPB9xId
i5SpQwRk+mgr4ynF9j5N+rwKbI07+RbBVrKaeSaoGV3bdr8g124TFa+T1XILiF54
WOgP7XCMp8kCaeJtEg6hIkBqgUIloroqNQW9+rlUAgC9tTc5lq7Lf6uhYJbYss2Q
vWq5wvs4IP+JI3k8Sl+swzu6ieOXdW3l4t8TmmgNA0TedrldeaCERTTCOuINWPII
U7XlifP1S13w1HbmP6jLTVhEsLnqFCoOF+aFJTX1/3LfrBcoH43mzsYEyaMkFXkI
bVHD2JzR9iGKGPdlUNgwvJKHYbcWjLiMusKlML/JDM6JYksLrOXaHg5B4aPBr9hi
c64dS1uRNKFlKu97XgUlquOGXjUQ0nfzMyhb8sqfO7a8Gn2sAQWA5hGAmsRjqHMc
9uo+oDLUqsNrBndt4Gdd2czFaELEs0nVuwrElwqcrYA1W3VY7exzMP2ioOIQsKFT
CQ7KxXpqq1wI0Varr7/OHOy2uO86ms2u4fPcogwmPFl23WA77b0yNr4S/fc56QPc
XK9VKwTKdriHjzBW3eyUik47Mx6x9stlkfcMLoKLpnvWg3kSpFL91SCmSFF1rRZo
N99CcZpZuGHIII70bZzoviQBLnOXShdt0Py1ykzKY6u5b7Vc0vhWGlpLH3+WhGCU
AbYDlcQ/wErmpzprJeECMsAzNLeDFbpkUA2hFI7b2y3G69iz6RrgowTWOia0koiR
dowxxrxssYB7Zt1RpYYg4w1VDpt07VUBYk7c6fkI+Mh0zwmsJo4jKS1S2FbDRHYX
udBj3EYzLQ/BWlfLXoFIm11COhDGfiR0a/BLmxspT+1IO0maVTZ73dGiKW7OMH3y
vo6/h3qeeDhBXw8rcoeb5OPMU68E7QT4CwXhi//UZFFfqnupCTscJ/60HEyR4muX
1xC9qZxZaZBpburkGOK3bNpp8FOdryqMVdROv7RR6jnuKBLikNWxPR32m3Yc5MFf
CD1BgrjP/+9fUgCJ442ie47dc37320ekwT6FHVUjnkmmEQGi80mgNxYJT2/Cu+Jy
SCSj4r43sGn0oBrH2914jy2wplYznGB3HIuHpDrfqz+ONKG/TueHEX7YsZQCvjDY
kOuoxYGjrmMB5xHmCB7As2idL1FKXtKtsP1X4PpnVo0/Cbqhpop3u9xNQlVFAClo
w/Nug1qlzwcoI7vw6vaoYJBrU44E/IvyGrYrfOsuo8JZ6181KeJP1Q5/x96Rw4Su
RQ/whFhzpYxag0L+gHzzpbpTCJvBqCwMOCU9CRJleqD1KGjxO2u2NXxd92w46mkK
4VIi0moCrceh+CKAJ2yJMCHnl9P4XF80kRPO3oofNbgIzpnA1n0RCFEntRj0ulgY
zKGvw/EDXXzU0QkxVZWmNlVgAIG19AMz77G0+HybhZYOIsHGlFfqFikq6mDKBeXL
6EXvw/mJG4+eDCh2rEpQuTjpHQfd+aaLg30jYtZwJ8w+3qeoaNHBSF2+hO2nUA2r
lwogITb3oju17RJ2zPDDK+gar3nei5yFL+aXcuccv/D5wp0OORh2RMwMAD7WigC9
E0AOrF3BF8MAFwdI1t0N2gmiIO2Nh7DESZwx99Ymh37lT7YcMMNkHMj4PqTTLuSj
YwG3PyR6tRnfIYw5DhQvBVq8KhCdVrhXDBSYAXLdlfnDqEovyy29iiPE3U9WNovE
RmCRx10IN9vVmo0jERbwsidUqczhyrCQjCRU7REE8ZgGo+5Ty5PTdmxiTU8SbUiw
cNENJdSQ4g6/SHrjP9TVhNGPXmVNDl0z/1ZoL+Z7h2JtJOqmYgsaAWR5mPrTeHjk
6iHCv0ZVj1t5QA0ddty9b27JrhnqPLZGX8cL3QRdcb1vpgNe90qNq8Q0fvdF4/zk
zi3NVcZcIStf4ABC4INKusHKmLNadukN0OksS/xB7vu79O4XKSTAf8Zif6reteBn
pYOKlJlumjysdXqzkAeWiG0TUq25nd8NvzCo4ALG4sk3fl5PTRZyG9CaSasgaPuB
3XKJoxQs6M9Ck81OAx8mD3OsFdKmXVVXVoNUfH1DCeI3xTaGZguNP/PefvjVUzgb
vvyBsiWDEEk5Pe+tuoegwDofiCW8UMX0kQOR4lRl1cHMDZ39/TpOveyXiM8Bld3c
wmnjc22vaTdmOCBxOO7p+esvrcvqAXVdCmiHEl9GgEdq+ircd5NSQqsFiOhhP0E4
e5IdDv8bV3xI8sEjOFfFRgE6R31oxfKUtROOpbL1DtZJZ004loVC+CmGbKcrfMfl
GmxXEPkj3JEPkiSFxN7Mjz2Go/d5ASZQZOMZnE9oPYaf6+4LKZv849BR5fLELvCA
Ujl/IMqISao8yLZzNE7lH6epfQKxBN3in6TVE72O4MZwxyVijkc9YpRClzTMvfX0
NUewZc2CVhN6NLactTwFGCrQy4U62pJQHGjM7DHDeNFAockiqnS8qroEe9vlhE3n
JHA0JineuWrE0JrSqqknWXnt72Hl8Ag6M7AGMWbvTdJPerduCJNgDhjvs1AEtuAE
iTUg0J7CTYIIN7Tb6fukBONK3K7J+OMxOiW0hqxyZ1Vc1vbSeCYwGvUv7NkN2YqI
SfzcRdldYWkEqB1Dbo5T9KS3vSHj5Ma3IS5pADgBXipoxUU4OmNhDt4ButMESBzK
NSf6IjHtfxpBzu6MsCIR6NqxKAKxujECkcYrco4iTkqFGg9OqzYDmO0eJECtClZf
ho8R5XoOc2/eq/fGxNyPGJgHYfbuuTQCsAxYKvMaQf3DonDcSll4bhlmfnQhSxMQ
Lw5c8jamX5MfoSqlrfutfXOYH6Xi271ZceuJy6eypO6NIvOZfbh67KqX32V9eLh6
QF+GoThs0R3dfM7rF4SItwstA8x9oxUXPS7e2e2tYQzrg8dGPeFZOw1x83RwKbHj
XIUNxjjf1H8G7FwyyrsrmjHekmPtNwwVL5gnlOX+CMAEb8rg5mmlFW89bhcem4kx
PHnOE9oLPYvqD2xON87tCSQFSCONl7sydd82RquKa2gUOJCwD6oSe2xUZHtN2sKl
GIw7bmbRQvyqRg9ZDUtaGPYpg6m+GZNW/aLvQgobNosuAP3gg10J28AtHCpg++N9
mAAqq1Gs1o8EgiQi9z+GrYbapbGrhqT2d0Fe5t+6JBHyHHzH07ztHXbFJl7EXWM6
uxW95ZFZUmtIee5mEj+xoYEUVK7o3R+Xgg3yWeEd4xCu7Ik2yCADfK4X9fwl8plD
xIVrOGrEuT/8p0lyUF1uUKh9B9Kgm1J0f09lFFUbhbKTsE/i0BqOcKHmnbn6BB/j
2lNPoBGnxuOISRlv01oGuyvWosSxFor2yKroYnJ8ymfBurWveLNhk13JDZGEpwIY
FXtYYYzIiFdlM4oPiDH/L2YX9ljemawi450MJQtMIWdmfvCYviOj0oicLtw92JU0
ys7W6M1/+BjFTMugQC72I/IwWXwkJzdJHM2uq5BnRYAiIo6zw2UwcUAIsfQvIdBl
wxrjKn2mdh79uAnw3o2Escf9SvVyT9kJYrIHfqiCYt4vhK/w768c1Y44T2oCwGQp
DZHqSOuN05ddvZ/T1CBxHlMkzG+15HoLS8Yvw5fszSgb+rSTkIztjdzKAlth5ucy
z40N5KRbIenjKqB6pf2YDO9XIdCzLJcFz+1kcma9yMORkUCBIpVUgp9Nj2pvjHvk
MlZmBkhrNP2Tmluluy3Hw59nllKY14D2P5WOmZ2Uol4ekr3SyyFzFbJc8Xvx4y//
B2yPCkzpXRALCsQmKNk9VxEG1STAoD3EpAI2SLok0Y2JBdex8RSQcJNm7TH6kBmh
koGCt9cRyB7UgR+biFkYEjisbLikRaXCLXzeTPZmj+ZWh3hlpXgrnwZC93qCMyQo
+nbdiyMJFvBjqC9nxjgagCzyQ9zz0/Mb4OW35SbrdJesouxaYyBB/2EfcByJD70F
GXlYUWK5cH+8SdbdRXRUm9mWy7xeBneHlleFPW7O9EOUSL7AEMywCfOzkV1x/Y4G
Kln64AwPYiyhfNTv5v7kpiseRn1Qdr7jw4o9wJd0TUrCnYR8yGhYlbnY0ps+FJYl
BN3K9g8MoJt3Vj2aMSGNwoAEzYrOgDaTuctaUPl/SfyYcGXFkR3N7Jrbvt781Jmz
UuDw0uoTB9XSm+Dlg/eJn5WgfSX0dpFis88xQ8XB+dwq+axPkyCQ+j90rvWiUWxz
eYtXbzJ5xh2MXJn4YFe7Xk9RzyYnCya1zEQNhrZQXPnsAAg+3txAIeeW8WT2Q/ex
Ayr+DkkvIfS5XihzugrC1lBRr6fabQdqvUYmV/cP1kqQlBV1MO2epirXY9BHXoIR
tGg5vpUTTo5xg5AwUklzjTU7h/QDVdqOuupL/ktW2jJYWLBW6mA1lec33dYgpv7u
s6Tu04Bu1RkQIW6S5S6nc+O1pA51H1UN6oopwYtC10d5BdNDkE2Jvh/8Lq3ZiNbR
iocM6W5llGPJ6SvuAAMS4mJQb42N6WrOhgwgLaVCXHN6iqrTZS+ABOHGhgkjwKcz
GTiYObXAF9sK+tSaFUHGHcGxucnNHe/QJgjDpi5iDliX7a9B1s4N6U/il4hFQqoJ
g0JTer9V/MtLTCv2wkvguwTDRwaX0GzkFH6l3iRplF77A9QUgJiTjBCYoTRWTTN9
I4FPLjOiXvOD32EcNHs5I2npcPP26MY450p6DBltGFouvu3+NA3rPFNgkJCFN7pp
U50iHNBeFxgR27qX9AoA/GNnnZaZ+WIbUuGbBzTCNydrmb2ltJtz16aywNBYMeTN
071fSm+ElBjmwjUxg0aAD6y0ITqTUPBqlltF63MWKgJ3yBPQZ5N/fmrTSKd16Ciq
/YpeaC31/CYw3Ryj58P9SWSqIAjiwUOU1jdWUTxodpxnpdbx25mrVZFvmoRZWcbc
AQYHEzVfyhu43U4dWyCKaM3He1ywbNBfJOO8ub0H3M37e079xEVD28JM/oAKQfUn
YBua2FGq/cnHEt36w43vhLYQfAP8ZqtOkWRGCfNJgkoDvjgqOB6qul8fYvorT4O3
Yclvl7uDhNB2ZTBZgRtageB9w2DlL7Mb3DldURMNBW8szKxKnJ31nJmY0Oey9M+W
nhCR+v48ARcJuUcOSRU5slRzd2FvjB4prq7UIU7tLWGaGPFa1qkGQ5BzoiVL0Gz8
mOwUicZQ7iyJq71PCWQGs0rO8s9d6fQ9Q6vGgEnQACz+jtt6ZbFkHnUo/r4cjqlk
goMUKcrX6HPtuYJRhzil+u5MYT3yNVuGDTs4cuMrOB5uL6oCVWJZaaeCtpKN4Fdt
GUtprs9IKnMH7c0e5rrYB2amxGpdzqDOuSNRpHNp7weXU0ZFNDU9pZSmZgFeY2/5
yV2LeFZj3elq1yPqw7DiaXuyJR4bVj0ISWl4pFbC/SG25n72lKLrHtoZPsP4o7Ym
WsE9wWY5RPgdJdBhixJX6YbADG5DC2hXfgZrpJN12L9Em3PFa+9nAUwy6zrCjLCr
H7LVmOT20GP2d3I0rIV3KFSAGyVhFGxNgpVY7DB+SNYjV4F0p7P0wPDri2D4C8cf
RNoFp+2o09NBARAA6yZZgptDve7zSl4ZlI6DvkLQkV564xNRdlOrZ1t3OTWDRGGx
qUYEcksNeDlj07SggGOxblnUBsYnOc0WCqKWe8R3rrnBfaNJd4qg7ATtYGWbhPyq
7930Rjbk0rzIoGOUAzwWBvkkiCuB36U72ZCDe4gdwBhhFuofNANdHj87eREwNcQy
FoihvDDHiBAZ+3WH2AGnIJm8IbxVWYVOuK8fPm4+phwKe8lNLC53iTNjRGmg4bxj
ARieVT0dCuickSj9Cq6W0BqR0ddApq/syLyViGBDKBX7w3eGmfqXpAljwUKyYuon
IszoaG/fkPhCjQg7c+5nEnYJbKb6qC5OA+KusinEyw5nW0xG00GH7fVJvMNuDTgy
1oxKU2S9Szt3CU5Cs+PN5tsP21YWp6ui4/UD2X3YtrIXoXLjEqmx3Uw5I1+k63L4
ud4uQiI6W6OZn1Y00k4tAYNMu3wMn6DlPlUS5BIdfD1uRLwIiPYei75utc0Q2uRY
dv2yCp0wMEhGj+AuTTbqr7gG6MgpOxBICp14TsrkC1/jB9E7Hj1SKhWaCYzVH8RW
BvC/547aQ5t1Awz/DhXRKiPfXS1XgXmhldPZMKGthdR+oGJDTcgUmJ1m40+2avI+
taVf5Rbw/gVwcff5T6lW5B9NSd6g17vJoXyP22w9nH3zZPhblAtNC5OCbmTlGSAZ
ehGMhXeWlgzYFJhQh4L/GXcQE5bDiokfwn/Fjpg/6ye88yUjzvNXgMZ4czillrBB
qNHkXbQV+ef6mPTSrCRDZR1yza431+LqSbIUKKi2j36AQFKdQN3CxrLd6hEHvefJ
zguTJ/QTgBnSGQ2XpF5Q5Xme6M1KInYWtn5Pq/fpqd6WoJZx7UAGPSZw+g6B5fCu
H4o6hDWRvNGswvTtWne3ocmbvFUeSL9W6WaWAH6gU8vmxa/XXTBM/eQ/+Yjp6Qt6
O6CdKb4PIbGCAswRD1QURHnEJXcyAwo70dPIc9h9KSTuC0gY9acT7EJCiicUAMFY
`protect end_protected
