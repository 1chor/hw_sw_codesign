-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kxjp76xt+UNISviVXyqa9+bmXHEIrnzXlILx/WtJnqRRgF9clLrmDsp7HgSu5Poic/C43h8Xv5Np
M5LdX0mIaTdLmKjI6CB9zfF2VMFYXeIx8PX+Pb/RmiGuX2XlIbSbsQiQI7VeKVqoXxUMTkM5OPMF
V68RlwKFoB9y9DW0wQ6C3974K4rNIbTd0sccz9AVNzzg/P9+ujR3sZRtK4CC9Mic3OYxDy+Rd+vB
y39Qw6IWaeUB+bHoRwrZkPR2xhCbcwT78WPj1VUU4vjaKoAZD8lGoVp9v4ejsjvBu/Q3GJrFChxQ
zwUzXUJ142qFWRVGQPKIuBrOFpBAaXn8HMLnfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6048)
`protect data_block
Sx8gBnlsUjauxBWyeR7LtN5VoJGNiS+3dZKt3DeOmEija90VMkyuYSIjBqgLJbwz5UGnilRlTQ7H
H/1t2hNoWL72vjdep7wsGEwQSUO/P06zLB8cRv4Sh63JdhO7UMGKvf+2Sl1aTnr5r24qOjs3H3p1
+ULSca4HjJ+1NnHQUH6+Aop/1IR2UMQehfhoSb79SwAEPyzCmQzMos2FC5NQe+3ferBro+g0Gno1
xE3Fbn5iGYBLlMYV0HGh7b3zZing/Z6eiT4sOi/HLcf831/uLe0XeguMHD8NvOBf45jBJ1X5pDUX
+RlCgELlUBUyq+EL/1llCNU31LPLTHtdz85DPfYmPyXR6AIRleT1+Bmr6t//iBj9JRBuYM+/dXmd
95E9uKWF4rCDj/knd7Ret9vA6VZD2JK66xjuKZOwQECFhHNb0EIgGgLpXaiWW6yjK7q1FWHdkU3t
u5hcNy8P2/8ZHxwBdzkC1paCH6ueEaYaAxMrfD/kd2YLJ0W1CQADCAZ0zvp5jOfjh8l2Afv6XaIA
UYWVRRd2boew0Rm3h9A2NpewcrDjdRlsLnEfG/+XEkwjRPgVnj6zwQ4dFjXeF+4AgTIg4fF/+6m2
apVfvp7mfMOoWEPEjrBCf0jHLTSp+i91HH+fWLmgDj2zwxxT5Yg0WU5SP8nbua9AKDBSTEoG/dEZ
q332UYrNP38FKOWNcBQgDU0BJgksmFxJCGf9WX/H8Q0oQ6ZOi5EZkOLLyyPNGEHlgFQTp0pFrmT/
/XsXzg2GUaDSpKTrkggV/rPlQQfLVsivBcmr3+0BZa3SeZuv3c9OYLExqEOrg3AlTckYwWu7nteN
S006AnijzfI3xAbda0NLAVisjYp+ZpGjYAcitUnHNPmotU/OEWU59XaINNZKVpGmRTNiZlNwlOlY
ZwJgmYk8KbuuIqDb2del7QZZzu48LGq2plvtYN+Yuu4mI6zbdZkT3RFGCOGV758nZsuBkjJEqNDb
3+cNkg9eK+xVFTLernGhpfeyfGshSzwfo7wbR8e/cpwgXbSNdsXf8P/0PkBMZglrHOwrGJLOsI67
tYWKqkGytZ5WK1OV0l3PSJ0BAtB6iWb4GUnB2Ir6vz4TAtF18rlTIndoC5AIniyTt3pNWwVa3mpt
A/qy8SsohLxHweXGz0C61VXFDUOsXe4veTwsPpwD8vVDUWIXw83hNfynYKDx26gj/+Z/oiqpnX5G
nzWaSjosFC0Aop+fREdo5eLML4pyNb3bFGqaGOocFxGyS+w9myhFZ/j75pY6SlOGHpNF+3U5Lxqm
VrPyveKtu0ASKlizvAv2JzGYXgFmdYAW2BtlTPdIkmhC74Licuk8MiBDzRNjzB1YbVvVifwhJVUq
Eb23Vvyr75AH2WAJmf+7gnDnUjUKEYJcIbx7Jq8VZdfumjnFSVIC3smygzyjJlNusRhi33QQKbJ9
Ss8/HPfK08vhkqAlc1F4Q9rc3aiBepQ957D0gyEJSsYc81qg0afYAjnOYMSaYN2x+RjroncxM46r
dWfEBtl7eTWuxfidWH9KL+DTiC5n0D1BtOXjLQMUljUeVOt//59s361D8M4IRfd/UAG5LYkkT6Pt
E4+3LiINSMTdk0nIV91YieSnS9CbtcMfWnFyKKVjsIkHZgisTc7pQB7nqOnbKt9mwaBL05yv2H3P
cjGvkCTI5VphP8pMaR3te6kjkXvMuVXqJaJdorOtMeaEmpEgSmZ8oAH8H4s03YBZvgp8w2e0H9Dd
ba3fPGvr4gSPMIU6z1pJe6MeYkBJnZi8cniKHjcZs/ihUMP8KZfrUv0N6W3F5mQrVcjPHK+LgVAb
flCoaQUheRV/s+8hRsLQm5QuWTyVNDO7bV5DgpWkxDRTqKo7NM995MMZSYAQBk1VzbJfmNG8pJK7
3b5cJf2nGQwlucHN5mxtxw7pGthHLRikLFIaDexZx8DSZi+zmpn3EJy5zPlUdcy0+DAClf3Li/dU
3TwzINREdLunHcculdtq+M1Pr7II9vYY9cqTMXI5RvVITRLAPpru/8DSjVynXfZgP+4ms3EC+Wc3
F2TA8jImylcmS4yf6SZ9cGV88v1vMsUu9E6E6jVOQkiz14CgnMYG6+jIORSn+IIAFrfHhgOXhLql
GRVqZsxOG3nlApSaBeY9PIXNcBVa8LZoBgq93f9EZeFYzXoY1rTLw1KW1BO9C9G5pS3liBd8LRPM
E7FFE5QYNyA1jiHONtI634cX3TYd2z+wc0d36KyGZazTTJT03BINRhRKQgLWILYE95n1+g3M0hrH
0s4wZ4nftsTkvCv7EWts8SkkmTRghc/4co+EKu1K28jzvTkm1cekZZ+H3vVu7yyoeDjeLT/Oe1ev
c1yjDE5H63jg3GoAm0ZZNEbMSK4CX4r4a66urT3ChASZzG2xBhLEJyfHzMu2pj3dN6nC0UW2bynH
IlDf6tkg19oiRQKmjl3Q2O61bcam/+GP5YvYWkjGYFJ+8UIy8xQS1fpAvuOwK0uaPFoRY2d/KqrO
FcRoxsnF7IXcrJKbi8P/qDPiXyUE64S997LPB+c+joESrRRWFPYBICmrjvx7ecKLrGfgNaCX3A9E
bjNqatsAOUhWUM8CWo91gBkA3iYTSJjZyxA3fJV2a/C7bQutwnrhyeAmGDNJZ3T+sje4GVcdqldd
ScnupzbgJAqBamTfH2gj+ACzdmvvM9nWVDvLfSmN+H88NIqv3ndVOA6TXkJwswzudHF4Uc23Sbco
MkCGIuSahJL/fctIu9prvkzALb5pZqmTPtHtLl44khKOW74IWz5qEsqxs3cTW5hxno3jmD9bj6AL
SNj4mP/Yb4h/MyoQk1hlP4bxG8c05FlngoXcPOVH+QuWHKR0BI5bzgXpHCpqpmMPRTEqd2t7jVuE
FEiO3u4rwSUsLNW+WPxj1oqUSc2Jx4JtncGdqDZAjqY2ZiDKo0XVz6ZF/asAoif8JKy+4LTyqqG8
OtIDTsp1HrSA/nWif6ZwzA4q67AM/3xl249UlRe7v7YbNSaQ3mild62msnTKtuPwmMikN3qg9i4q
wrGq4/MupvB/7XqC37qdjpC8pjGIpw5jwpjWY/qIdxsxdQhvE5dtevLyI5JlOdLXQfeUqDC8lFCd
cDYsZ1gRTZUWMAEBGIdRGUGgPxNrD5JWDy0SDd7imcHbOhE9Ylf6OAcmI63mQF6Df7V7BSp6U9yN
/x2Df49oQfFBPJJJA6yDyxMfsFliWT9L16tTVXFh9YYJvyeaS14ZC5vAMr8V6aCzVTXokjCZ844J
cQb/v+FkJTPWaRxg/SVp1WLwG2vxztIxyWpjr1KezcHl9yrfHNdxqm9qmxL2jQsojU24114OWe4J
afI5uv7oZI+E0vfnp2u6l14BJ+a/IN3YvTK4thcsQbvVOpmC1cBzjDK1Gojrpjh8SCeO7hOdXaRS
6GxQUJmfWXODJyYWiCNO0XQeEFGYXQDgsHoHOdG5NNLPZ7Qfh0ps0tWCuEU2WKNC1jujomLNE6Q6
qCzUeaSPPLncP0uUUZfPBX2SkxRvzQeozfZCvfR+VV47bJdfT3FlGbH4oee4oTKTX47Wi8LTe3pA
9abYxuKy84yG4rMIV6giJj6d5SdCKwhFka5Y19csn6QzKoJA8c9RmkuVX3S5FC036usIuekGhup2
VN8PJL6oKrVhHdJ4IcY3vhmXPh1YlW++tsujGjHEHU2hYB8pB8DouZvmpVZAV6uRQGEuAEEgwTaw
oDj87G43CIKxN61hmLLsBt4wSOE5Ds7YhWHL8oZ4B84zalG6dlERQx3jSZqqb6XYyhPJJVdDhvNx
5FdYpuIAFfe2t36THkvvs7NZTdPpUIDB55kFniAHZO9MdFEJsj38GdTVdJ+jpw8E00a+WhEe+WGy
0p6Dm9gv0npLI0A4kRmluZNJ0jlVMLr6I96QXzPlSzqcsAw+VMsEG+IeqxTBz5Kx4ypk/hxIjufV
P7Pdnpjf6TNomuwNp93Y7g3Oqp/jtQP5MQPQcX2tPvyR/MaGXeLnhIUv2O4XTxkOih+pvs46uGdO
V4H0btWfSu5p3reVmsdkNpd74lWjmkkM07DHnyGwKG5L7zAMCBBCJgreVo5s8H841XxB6RU29quh
ivjpmaH4rN9uM75qaWNVOTYNgjVQxOzhJB7YK5zcNKe96TQ9p3TUdQjzt5J0f6h6qAvkaQkuQH1B
DrgApcibC+9x9XRQbyQtKRTPIKWSKX6hr2smAdU+gekVSGaR2yGkojohTERdZWOKYb06G1u47ana
wBr5xPTu7aZgBTjcw+DjOJUrjK+yAu6+1qBeS5hCbrvQF+rZ3xH90b+8hx6B2sLTWZMGverPbBtj
aP579QgRErheRSbobC27lc+yfrR662VbnitgKhplZtzVSQDBOzlsRAAjuQWasx+q8+T8Rl/DQfkP
XGqkm4FDIVGNzHqNQoej8xqq/tXqEOnH09ZkxhFfxVfVhcXlNHImf+TGAxBwMbNnJD7M3h1cctWv
DToeWheSySUztIv2oGuV6WUdwU54zXcido8K5GPDfo4oyJBOtxZQXR3LgGV+cvL0hzKlVry/hVZp
L1M0FuQADW1YL3ygKfS7D00uixN4Q+k3BfVd6dLyr/lsFeRocaHhW5U27goAPnMXjYO5oAjYykE6
8aMNnP2KqKXoqOvB48qb4P6eHp30gIK/iKt7470BeiiuovHcZ0n0u2f/nKWAEgY1C07mXMx8Xl5r
rLN4qCFqcG/B3PQYCU9JUecBdkkkzvW5pyNmyvc0qps60FGKPAS+rQ1z/1oojU03qjJq8qX896NG
wgIaiaZ1S7nyA4+QisUTMnyybGXmSuVjmDyYtjKeI9CZnVVGSWENJ5HwRuMrRTi4fWGm/Fc6dOp6
748IGHtwKdYz4UuTwKuqQNR5a0cAWUuxq7XhtLFUm3tZLkk16cuuVIjyuJ9kVspEQAbilawjQ+mB
XgC37a2epHbIUU/InzYKrEA22lJarTXXE/ph4svcjNDlxElTKnZ8P5hA7RkQyk0waNhxnXMIS/Vs
spOaMVC3LArO7g7x0fNkLV//cMzyBx7TlwZc23wGd4FIrTpZUE3THIntOeRvuhUveW0Mz37NAPhB
/fiich3euvX9DslsHdR3xc3g/Ok13XsziJ5vY+mHYKi2Nh4EKkiFPplFQOszpcdjeUlmYialE9ny
vxdl8wGYVnHUqxhByahHIXx2k1AkcMW749CMHpwFPuja00ogIBqFAvipCxQk+R3QI+JIxqieRVs8
aDw7+apIXJJ26vAReixNafUZEmwIvPdiBqqwQalPPnMMx4wbz0NyhjPIHxkaWvx92Z467Ugqb59X
3B5q66KEBSdibggrfigggwSYWrRc8neGN3vKk4ZkDdxgItFODssFxU7kzJvaC+8Vx0dWrUVutJjc
jY7fMWsx1aSjSCZA+FjdUfEoxwUNgGvWfj4ZvbJ80kPRYujL5QdHr9X8SbN3KTRHC32dbbbE7lzB
JgT5f5W/UQXiWRF1zfuNOwEGUxGpo2saDvtzdOlfEDgrFLDNRSt+RXIzAtBmRgdicdrqIggwgk4W
3vDFDZZYecnKn7MqgBNJZQHFA2i5vIVB6AI9/b70ormFJhRId5Zi0EUIsFbc8a4d2ovEC2bs1orv
EJ6M5cRMeBElXAx+Czql9fFF32kAxi4WDelj4n3VZESoom26OwqfQqUhTmECaJJzUMboPCoQN191
KZ61kCekyqfh8X98h/vCbD4pkX2A6OPsP/L7aWEu0uPHG2+GhxyJBmfg5jWJWs05cGUUWDPzs8/m
StvjtHNgwHlu5kQN2xV5BDGIN9+h9edNpKPq0eTM6V4HfFdjKLo5iT1sm/DUkUQcckEbJTlecZhV
Y4AEoRaGvpsAragXZMO3xdgnJ/A3vc6Qc/oSyyb7Du7uvn3m+nmQ78t5Pp1UnU6FuJPEvfI/X344
LRAAx/AUlTa6Z6G+2A5D7ao6GkN8bgutf9MEEBzc33c5C83aEia1BGemqOV0qwpas8pbHMoAuVXh
wvs1DK3W9u5fqvY09GhCFcfT3JJo22HSHiQHbmH6/v6uFGkWqjUC74wfNb9w46sB198wFC5dmbXD
W5M+kbNQOLB0WDbcxqRiPVp/sOzkSkmnHOwE/F9Hpvcx9XdydaRs0pO3kpe+2Uple898PrHfoJqf
BTdRUnsZQ+kAGRzpK6BdhA1NYLOS+n5eFPpespsikn8jYylSI7moOrQdldclvOuxggPcp8clJLvE
tIx70DMACrXGB7xIvALYyYzXmBSgI4wraHej4w/1cr9UUGg3iM9xmTkF9ORs+MJgyQ9otr6BQFTG
0+3AJZAW+wiq0OJ14hBzIp/GGucRPGLUr4hPBHKD2U50Xl3H6aIvSys1ss1h29R/yl9M3dWiC5ZV
7lP0802Khga4bN56VOATlFXH6XWE143R+ApVBXrhD0cky2X9NBSAcpEQzg5JrFb+hOoB5lrr/tUx
zBqGXbivReedUbF8uPYPXR8db1CIMGCvsDtCGjjNwV2H+y611UVZvW9ZKujxc17fkELqtEhMwQes
CMVymn2ofujKN+aLYFtGpCifOZXYwgymwabWSAYDPlcBfFzOM8vEwtrJ5Nqe6rKyRB+vH9mqbErM
GYgvwNMv0fmzfufauWdnFf2UxPWAoSdTJgCr090IKXpNRgmxlDYJgLhC5PRo+yCbfV5Ioun8qF0c
1iAt5nAR5DKundtBdUjRgxtOSeDGY7VVMwxzVXzHJT2yuqZTv8JwdtyPZK4UPB/zimloAk66B0X8
EVuMUViw2aMfXkyOVkVtY5cXYo13i3kS+BUhod4nmJw3znWBLU0TYSgNvJEHQCOPUs3s2K6Gqb7/
T9Q0aUkPh3W0yz/OIu/eHlnvtwgO9fLO+XvaOHuax/e8Wtpm5TNJpFDhzbFelZmJSy/f2HsF30kH
6P/2Xaj0yc2Vj3SVT+0ICLauDiuH/75aiEXBGH4MJSIwWbogVeZyRngxCADw8sJRQoL+vO63ZY90
inOrLq+eqCBL7ZMFfsQ2hqJEqNwQ6LFSOzBvyL2ONwT4DGlRCzRAmB95P2ZkFzbA5bdRqaPgjLfa
ZcOQfWxPA4rdvIfwpkeSj8BYsDFP6ZbNEujgpcCCKpimHkl3DnuiDF38DUgLvzJIA/ddqvX3wPxo
jTnfn4EqshCCkmn/vmpnHXn/Iclft02+U5GNjcqVoz3zpEArWqiFJdyd4lST3tjJWUt4YBhS74Dl
HcoKhEV1kQd4fYgQ8hZHe07nwg56ogIqmTr3HT0m0lnR02ljRn1XjSG8PT08DtLqIqGUTVZe1j1g
YlM/E/W+tudzRNMFPOzujRKrbQW0TXpraqIKUDnz3PjUL6z9OX2CJh3XCktQ0dHpyRu4EJ1YFb3+
PTLMEhOZsbLq1i8jOZ3PlH6KIYFVNKo8WxhPsM7bvQxo6OzSbO+1qM2Do+D5FfgHoZaMsxrLIhHd
x8dJPpW3GGPFGjjMq0dd8lpZDfHp6CZrY+GIPQNrTt0yIkgjhG5rXbUrGJen2Oc2Hbnjjbrd82OU
4ADXVvViXRWBu++gm4k74+dfZRzpYnQBuDPP5yfpeM/8N0FjRyuPJpA0eARQiCOaBB3rc21QQDbt
iEvsYi0Ipu5LORkOeXgz29+ugMkLW5ywgO6WAiuCZomuwhK+XrH64I6xztpU6homTS++Md1G5WCt
ZLAOiaVfGbCIyRqQnNQ57ZJfa0YKbG6k8/S/1rC3+yTZEq7kL7pS/lHFl8bkhZhAIefMUTZ8qF4Q
x4xjgIOo22FRzIk40OhXT3PcFHahw7XE0KXGoA54g6+yX0wyR24pWVf5krtC1DJ+dOcGDo0mQKLg
P54wVnkRm4crac/Q3t+wxQ68NHDWl3bpP4sbQbV0S4BkpcPq+FF3EdjwtNmYct6ZUOIPS79G4nhA
nKS56Qx/ohrhkrjnRqNOg9pt4b+VnliTVUJX9NjyiiYd+7QRHU9vAfOskxMGwqZ3N207UtUSS3Uo
OIJeh8KBhOfP+969LZyQvtm0dDudb9VVmuJDkXQojFeI+3P8gVnvXTh+j0tOP8Kn1ReoRmxQxo85
RsbtgR4V
`protect end_protected
