-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BkloG4f5Snu84970AQ9mqFxWTbZbJFeDp94IrA4x/g0Rk7CHItN7XYCq9x/Y/soy
D+5tVc4CPhRGwFFry8ST5hM4cY+zveZxzwGxcN9piZnHDPNCMaqNvbw/ZTvqWpGp
Eq8aWdh7YqSbAo/1GOWgs8xAMlrQQ6A/kiBJPuPz1uMs+U/ADXEckA==
--pragma protect end_key_block
--pragma protect digest_block
4hfoWx3uMLMoZXdXF3gDYeJIb5I=
--pragma protect end_digest_block
--pragma protect data_block
A2/59jTZ5UwiCCHDEHAdr4sNWkIMtqyNPDR4P4DFTFC724ufCj8mYBqO2vwiEO2U
BEwVLHgs7bjQS6myWzKaMTp+3h34/velj13m36eJYJ7PBtdE4nCdYdB2NVe6g3+U
oJ0eZ1uNZo+R3U+Xf+/nvOab44nXlAM79BVsCjqdM57TZ5OI0Hkw+XvFSam4w+/E
+hZG22GD06NVaNlhLOEARFa0Ep2QGMFGruX+A/fBI+9z1uHslgP+FyAII/ywBXrO
8EBWkUsgqaVBlLUMw2yNUTZo5d9wL0KS5imxw14Sy4IET8B+lfo/Pu6fQo6vegCO
MGD4oL802Q+sl/TIB/tRS/F8jQCdy9dVJialF+x5TtpB8MXhbg/pi9atVM5peWgl
6Gufa79VkB3NCoc4WaIOnTUqKU3fQ7HbEIamLjgKOigmcUZPL/LtKZ4K0vxv0xXi
x1a8iww2QouMRcUCi1U7AjjG9WNInvZyE4aEbUh9gpDxnQFWugRG6/MgDxPZmSIb
BgthRSjfroBeEy7hs1A8H73JvW2/d5vurYe3wznYG6qCwyiJrEkJqv3OBxymN00P
yDXIM8d2ZlnlVBDwF0+3QaYIePTSkXFr1I6tKNbDHwo5oxopxoQhDyc7AyK4s6Vu
P3LmfQS0bF0BKTuXTBePozITWt+q7Bq66vbijhvOMT+K8wBWmElX74zOaNyaLeP9
YljijSOyjU23GRSN3nQOT2qN3FUAuPdrrRr14/gqnoN6V+mogQTbXU4g8DPZLjaT
+iFfz3WCaZ6WgM4TfEfStlO8hMotxitSS6PDYBC55t5kN5e1OFrzQ6cds9zdzHas
fJvdHzPQu9l+1AUGeWrQyZrzt3wEWupvw5En+gjyWirX9SJSsKfgAul+smgL/gHi
+6XqTdnuWi0XqurBt2UceOfZ8J6k4Q9La89wkTU/TRlC+bVw8H9966CVmbEF5gzT
i6AXUXr1k4fP1H8w12L+DnGEcaaFbAayKWSUz9UohhkhVElsbOYuyOKDL2XcdTcy
yfc4RSIwwlMNXKFY5aSbQneBcPCxoUSMLOfcSVpqyJkxeCj4yvRXzBfzoVTp7ufC
rBcwgSRbqLEC5CD9wBmyZ9KZ6l8pqbaRj742GoCo9vy5SbnoTIP+IJ5ObIqy48rI
c/TyuCCsXW4b8Et5HcziCJwxvv9SDKlqmGVkn4tg3jjBRS5qaasUZqz2kW/dBMtd
THMfft+kpaA/UC+E3sXpfZFvs5YKJ9iwsoMBR8JDNxCnFaSr/a+bTIWG0pJXWD9Z
JSRDekMMq/NFyMoPItS+WxIzyP7i8vt5cl1tTz9lkci8z2caVCBfKlRHJpmVR8lH
FcbBuzRSuRgmPa8YNU0srOxN1iYZWd8hCVpPeXgESPfpuASop1OQ5DmYIdsKEk2z
VAYKDsWEC47dBpvzdWo5MT8vwYAc+rC71qyc28v6BwjegbCiLTlgSpJWBz2Kq6bG
NAegnvB6i8s8MGzupl61KLnb8Au/kx6P0rEX6RFdnfuH0ZxGkm7kHnBA9rDCE9BQ
2Peuebtv9uQsbVFwZrPRLzemAA8O63AAkisH0qZIc7hGiHi8EkgjmETjREdolyt+
VAW0vyHKihkxO3CESDVMGN2ws6dtoAqFYJ8KYYCZOcYAbTxCxMezXmLSAsDWmJhY
QrUaHr1z85TaY2+BjVo0+D61yDvQ1EmidSt3OuxSDdoW8XPEFVNWfJzdMK9XaeKF
1Q0e55WJLxUQIvUfW5W945FmNJA2QJOvvxRz2BRRuoFGbYmtBixisWh3Z1HaYhkn
ayxa5HwKmUyMyX6SL1t5k0p3adm8fOkCFjM4uWwDSp5QN9emoy7o2MyvK491sIZo
WrtFPChU9++rbu0fyU8fsMuYQJTbpBc8W16uPY/0ihBOHTf9r0s+EghBnrIRXqRC
toUtps3HocaKhH2lLdNjqTdnA7iguXW/j7NieNl/QhqU0zcp+kkWJBEHYBTr+ntX
7ZnkmlQfM06DqHfakK85nYY17MG6wIqGDCehiCG0zsQCM540TyiUsXbw9MzSYCSC
HZt0M9hQDsluV40AgyiuN4bSgneeCmRR3Ju40xBsyRVNeT9Tpr+COUvcStFxYQH3
LCs2aXFpMQ11mpup2R5QVK/dqNMaKYFZxw1WFOJrQBltWiy82CRG8SjM51JyCVEJ
xjDScbNDbxwOSKNLvFpmeNhSx4hOx44msfzCad9Vml9JZ8KM5SsiPojkTPaoay6j
K1M0PoDvcGKPxCmgWIVRBdbUQg6msx+PhnnCfU9rg9Cxg0YsF81B9TwnCOEcmXtw
7ABiNlrSnIv4J36EwKSMc4wZozx4NRpt9lzTCMz0HGfaeqSTEsWL7cGIr4FZY01y
SMwOk9sV+JEldYEOul6xA01NOe9iDER493IsM43gnSsquHC9RViOvVXTapVjCHk6
aDUER7ArbF7xb/bv/1ZGdn+tGnOzfcVcQdIc1WnpEFE/AMijiSxU3sTcq2q2G+Eg
+QL+hIkczRR5vPFupeLvIlzEFeBr3txJ8C46KOGF58SRYGcXL9ITVPPC2CKJHxZn
Y5tAguyOewtiTVIYQyc7JSglGa4nH7Z/vByzsP7mOIR3aQV/EuakZMD8CdST1J7E
bQz3cwOsOXE+JRRWdUSGfmbLkfTmciQvGFg9ep8Q/ALmhzjdtmDfLzJjyYLHYjLg
j4RoB4cRBhYjRBBYc4evQtEppS9xp+GeF/T3/V9XQaibjqDZtxcCMOSYU5kwdDYF
PeAAA/csB4Sz+TDsVbQEC3sSwc2ZIcPi70SYP0OjtDHNQCA/V0rvsYPZ5OQ1dPwg
iP7xeVyEkD+aIdUhNai3q9WzMSdAN2cKIJebZN5dqRTmEm6VmMYwv/gOiegLn+on
TgZhdAdJbUGcnT99i42yabogIyJ3ZuP9aMoenCeEIcAycSnNrh49BirULCn4rXFZ
2Ox6By6NhV5m26uFkct/uVTEj6Qm4asJukapzZDsG2eAv2zTS78Wwc6kv4KLqkzv
5vBy1VHC2jDWA+fnK6SwGbdJY4AlARwbfFgTB1tQF9Bhbtfq5nTQMIvowggltaIi
N9Ky2JE8EBoELuimy8sBo3qFlrJjA0wWC0JUdRThpo8trsQVv18WJTpogbI8QKE5
qZPeBXnW+2rhHyIiGPd/83KKeTeUXjdYyANbBgezaUnD+be0Qsbq6aWM4Jgv4Ohb
j7rL4leu2TBxrSZ96Ybo19dAaJQQ8vHVtPWbah/PjgjvnCEw36LDJL2poRiB23TY
xlPq9bNAmcGfO5DfxJTDNA6OaSpAocnoJ/FP8cB5m/voZIW9PsWGp6qgtZSXQLye
13DMCxCUFonsn1cfo8YjbdAs7qUY2lC1QMI6ThcJpJ+TkBUIGNV7cjtk0wuWKZyK
NwyCUOjuOU29G/7ous03NgkCdfKhG/WDtcvlC+GRTKl1vkKxf9urhWNQ/Hfbm0wq
eOkHrn/JeXzPPD2ZsQC33FyjlVPsFOCQFk1C5Xsa8DFcdA3ZtGAml557bTlnxi+u
qCP98TAzOGit+BejTJEeCLU6TxfTYLuiRD4US3JGAxKqQfsErPC6Wj/uVb6DhKcL
FuMN92ouJiNe3vCZqTUGX8SpXB+WhwWcgIJia4nkzKQArVxIhYCZgodJyevU8oia
mWnaMU3pBBe17B1mfOJFYpgfuYzD74fKUVLKVAOS1aZoT0t5F89V6ZSq4/aYIBDr
8ST0Eu+mL7/5X2Qq4Sc91QLvr2GIrfJOBVSfrJ4woxNH/n+u+efzrhO8MUFnY5Gf
i2j7ratvZesdtVpPboBiVhE+ViUf0rD1wUwjIV8T0AU3O90esTEdnCb6IRCI1Vkm
ZEFkhyO0xjWovM9ki1OQnId+T2dwN7mE9nsPealym13DoVwX1BmtP/6hWMLKxl1G
MeH2OZYvvE8TzRW4wtAL7Ehuu5UPW6pg6QVcy3uF4fJb5WrxN7Z/X8NVkVx1eDzm
gWHy8J5ZLR3/y16Ehd88lZQja0L3UrkrtZoyGKImL8VyUfyY5LLRKFTU9AHYrtec
JmBeDaHe3IkG4EPIq2if66EOZSXwBHlhIJ8vUxrxPrptdHbMMRz5w1ZlKqeK5Ck0
YV8v1dqCVPLEmE8ojlpZ64RuGKxOMmtEvt5JersjRqTMpwTS7K7gGnzz3jS+ZQp+
EAlxlB7NeSkXEb7pLl2HzvfTYRKRBYlZrmzPgCy6V5rv9TECX6mHRzmjdWPX2kjj
U7WgFGs3WstFptOjIofKK5DwR0TFmV5QsyoK8xwMrhMFF7RxZOxgLjc6SOfxdjHP
Hxm+VAAtKFIFtaKB0PLVXiDEGpV5ShvnAZEYjSgFI4rRO+hEeOvl+4WUePyNJRMz
avAJ2YMxBDkE1yCxe6d4xoSuoFtw8q8YoxLqypGn997yMc0TeyQeY/64R21Oimnx
QMZl2v1B5Wy3ZwKjlTBH+Wjx1Yy0Hq3/Eu4YzwvSBtm9ZKOq7Cv4sfAOQ5hoOabb
aBEMyjZYx8q+hgFlQ3SOYSLGAvx7qusJWsnM1dTug+JcMDl6Vt0O8++s6qbHOxqB
bUqSj/EP/mAxg5RgCK05qajHcRWS+tFyvjVVlEtI1B0Fsk39XJgKhfSv/UB9jnSE
LrxtfTzOHA1ZNB9Im12sPRIHGzFtCMWP4hScZ9d8m3nBjMHA+o89XWOt7eWofapM
yQ2c0JslMDOuN/8/rH0KK7xrni+1WByy3sfThQvyFQpT+zqJuB1GeCsMZqDkv4JO
BqECC+dTaW7bBq9LIAF4gl9ujG7OtuL86Yt4/qpkDWshjWL0Ta3BizCzns2S4hwS
vuUd/Qrn+moVliuTcYn9JDx/rtjzC+P5vFstvGHTFWsJC/e8S3Ex03slBvZBrPfh
g1mjm0hBCv+Rzd1us9k1ei1T9VvA44b/FAfeBhwfxfVw+y8fMTqThwMrLNKny8QF
3MDRQiNgixB9HkLRYWGhYUF7tfMedc9f1KzD4/KQLTAAzujEujQaJh8JsvEZrXcl
QdIHJdauvS4hfnyZ6unPD1fXUAyztQotnVHtZyNkmQVdX1sxjjj2NlUJtgs3zppq
cBDy5+LBz5uzATvyXkuSZW9GCeDvZlyp3tL68CtopxDSQPu9I6elyq6CzKycSFba
xv4MQvaHP0Mm71nVtwlww1ePptcCtig0KHz7sw0xGGVnTYu43B/6bwYc4A6yZTjk
fKxNw3cSS94FJGeAKUvRPeBIuMVoD0l/QbxXQGfCPol4ELFvYe6k1nyNC2LhXcBj
V9BecXAv6BPAgH8n0TZDqnClsGX4kcmYKlmFCzfuOo1yW+gBKu5j/JLRVncLlm3w
nBsFTnw7ztwBuZ0SYSj59z8MdZClItnuv4W8XndxJuXpSVi/88z+OF9Y2PhgXtfK
MGKQL2ZFQGLGJhI1UMKL/u0qj3rnv+VoT8cUeBbXPsMOChilzPNJmDQqULzT/0Ff
0jpgNeVUs3wq7FubY0pu6zSUztEdSibFCQULzS2Z/aVvAie5QRl/Fk/ZO3WAfdEx
1ihMq9YphZAHRqqPrAir7C5Szc7U0Di5k3CkjhcYyfwR/v5MHbou7Hj9iS+a5Ixd
iNzFMMJ60yVB/SQx8kba1YEqcu2ZB5AzQrs7OwAIdewhbMCReV72dBabfZNsvAfN
qPS51/E8obHKOZqVaPCQXfKremk/Qu9vYwzX2SOqlqkH8NygWNZPxtAjQawMnKbK
HgE1woqDU3aus4PmVUrh972UfYdhDigoKIOBMTiD6GwWFUAQPBhd9xl4vMvruLx/
afcEwWT5IUJCQ+sadkbavyt0ze6RbJOykbUpZl4IjJ0HOpLPZPEC9sdnTn7Ffagx
DgdBL/9brkmeoCF5kcvHyifuTuEL9DtCMb7y4dzWZHoj8OVkIJ26H+8IYO2kiu6s
lk/UvMjK6S9NriwH95u96gyr+7735f4nv2M1big8B2VWcOxtx7Ex6NCCY0ZBbYYE
MLKz6MBlZDnPQN++/dEECccuHiidwyqRQMBUOcxQR15nz3Cgy53ewqeAPv72sbdk
uhiJUPFVcuhH9vaalYnk/rbkgp7YZV7X1vzTSnNDaEaFbLz1Ibh4MSSTsI79GQet
ynBQJVT/7BAOn7VwYgRL2PlLYHZw215U9JLJE+swKI9x8MbnUsqSTrfEydkvvccE
xrhNJMyMjv/nXR3iYgevjiwav+Lh1Fke0gRvKiIRrEtAfS+U3g6O8onktClgw4x3
+GfgR3zR+gpmlpCKk8stTZ/h2+cC9lxH6FFmCul4amxwaXyURw+eL11s0qc96/hQ
yppQOG5rQJ6JXVeg8tV42O5/feqce88ahCOcuyuHOmMktD50GxTMIxV/Dr9DvXcG
5qfEkEAhmXTwBNWPn3lz3qHXDDIpfvLsUDhG+oar+dLjS4AlR8KAOjeg7ssCOhzH
fXH3nsSw+ZxTNSH9pyUJ5w7q9ZwxuXiHG6Ml3rc+Lwhl7JUjMx0a0TVEjIoacN4G
Hm8eindKCUDULi0bPnVn9VX62MsIPJ/B6CQicEpBccvmsyg8T1Feuts18PymM1SM
TmC7o3mxDgLZjPWQ4ZKwQS9S4CsVQcU8T8F+chatTIx9hDamXASB4QrCSxw5/Gfc
hFogXP9knwRptUdwS+fXrTGQLqKGmmsl6EiSkpg9yJ7OfjS/59OaiEvhjn1Lbxwe
vcHm+fA48b6+0bzVoeo3Zp3tYutMrphqosmnvPOwvfVmPYs1Yf7ynLBZXXp+mV7+
ppLKWJvS5F93PYSD2b+8+kcx5yecZTjsC3U1rIeTclzDg8mYM8TItMPZXi5mvzT9
uCEQ3sEmGGUnEu/8G0vbBbTdpDL41hwSc3CyH9B5RQ3jHVW4x9TC0LlPTOWpC4HT
py7iyxkmmKfPa1KTwRgudn9PiKb2RYh0C5yQG/5JYw7p/L7gS3nYSmj6u9uV9zkd
7mMDvTsmTAMJEFLJ1rN4IuAiHEou9XELZMbBP8rnJRBQbVWR2aSwuzsE/qgQ9JBs
CmCyp0lZ9/l5oYjDWz09+5sdqBhhJ1JSxUsOVqA/XRHa0OFBprWYLCwWD7Bn7Svl
mdQjVCCcXUvoHn1sJtCY2iS95qHzruSuNcAtTV0neryQtt8EbzydXSZs1BKb/4LC
1WoNFavgTXF5T9x05Q9+NM6oZpyFrfhBMYk+eUpjadATNYy56TKa1TCmu2dYHlFz
uJIDa3Fa8ADjPwRHL9lyYEOu6ViWeV2OY1o5hSqwJ9DE4KQH4UB1c3nNH/+Www9M
wP44+Kce+wdRKrPHTR2tpO8q1iOhurlQFjjhFq1WrFCYepzK0gK/erLnJixMpSTQ
wqmYNfjC5blh6paErKPJ79Tcdb51INsKw+jLvP+5I1X/1LKmzXYHZJPhtpuhQa8E
M9qCElG8gajb+C8WotEU0jjfH/hE5PcqI1/NatEv5YoNuAyHcsHPig7SHBky5oGE
7rTxuyHTpBa+5/S+r9h168o6DYI+JYkdQYXsrM9Gew0DR2uTcoBW4Yph08dvy0ve
XV7B0DZEzVAq3gM4gki1C1dMhOHKtTr71fxq6eiahFdx0U+a4CnTsqC6lEIhFrVB
k65SOko99CGqbOpM5GhEuUpuUFiBrn81iqqJYfa0F3R6TlXRLu9RUlcEp2fU3fE6
BuY1VlpRfYPg7xDGnVQVdJkKVksMfXKEfcvRIAtMM0MnFEjzdlZdCyp7UnNZR92l
U3dxK/E2xBmFFjbCWeuwrdSdldOjS8vgUfj5rryWPzB8vfWl9YQI4Sw6w75/ChY/
AcaWIBZ+TLiu41UC/85yvZAl+aCaBqIptjK60QtriImqOirSLrgVT6blTHAHfPOb
vVIP6BpQg9HzJdqHhj78FRpyauAKk1lYso9GeCS5KrZPp9mt1Hc05uCi8GCkPjgg
bobCHrUaUSsZuvkszsONbsTqyVD8ERrSAEM0lz53Gc8Hm+e+ooXy53Hj3hBYTFL+
4lKAFCNqvnojWyeHfiEUqyi58tQrP3SIVKyZpsIZMr4PqAgUo1drezykDgcLKwq2
uZaZ/xYI5XaKSBHNMCjXbFrb65LU9he/qwnmSbalIzBW3FeGW8ZfnorZPoWfYG9f
qF3ScCUfLk/dFnCl/9kTn7oVKO3pmbLDj8Sl6ogPYHfYYNUaVpYzD0vJpOLGSExf
tucPYbU37nATqNJRIOIYLk8wrshNi2anr+8fn2firuSE2EGffSjhz0W9t/aP0yPY
d10HCeqxDW4IVNxU5oO41FTC2q15lZU03nFLWe13pQ4GjrOxSP/RRZhnsSi9imqQ
yQKO/bfYq39hC/ylI3MNahIjNEmWk88OKg5ezr3h+OGu8TL+4kQx0zhNCNQScGKB
pZQXkR9pNj1sHRhWIyAQ9TmyG9uxP4QIncddAQTm6/W6QsnvFjoqA//2a/l1xoPu
kaeTaWlRzyoc7HPkq90CSXxJmNXNfUza1AtxPpOTRW0r/qNSxViT40ml45XzuIhY
Gf0GJIgefsrF/tpFU9awOVtRolBbi3U+NTaoBdMNgRZnm1tN5zUkv1OonIPm3Bv0
ncz3zX546wQUmwYPU5SO+KPWKsFiaigp8EM4T573ZU4JRdffiiZ7XIhtz77zd6rP
9zCWFR/evxGEUpv9mDaQplVmrR6JI1EvwmuMLN2zvsBpreAtQWd54jGwURYBSIgK
ujfzLuMwDf/27LEGVkVgxXraB8qjpjllIcdtb5+ympLBsKNOUqXZ+iTN+btvvp/Q
nBw3qXh9SYTWtskFcOnqvgRlWiWHN95fVKdIvoi7by/QRJg+3B2+RnL9nRGwxxvl
ad+F6Z3V9kizY+qEV9unoyFZ1sorUJzr0KXQpfFr2TEaaYsMF09mAwmjD9bFWMgd
fumjhGNJskHqBmVbNIDy+mkV47y+ICELoR2FTKbk5YTwOuYXc1/3B8QV39scRqOh
g/ghld8PW6nMEtBueDE5Q7TxeFCSas+2dE+lLeVDV9NPmAMa9DeU+AEClzfufoiJ
KKkUxcXq5zO95C5wKvqIzgaV0ASzEprUeitAOqoepaJ2h79LcXIINktuRoMuzYwg
RtWsm5W2vcfmy0CdABy37iDQxvacHgeOuPG5xVKvgLW65/MVA3lofxm+MPSvxaEg
MgYiBzUVo8RsB2xYkUQmWmMYWFMgm54Vte0+9yYei19FDiruPJ8dwYtg5IP7TPFL
D8ehG+cNkh0zSIvpg8FBDu0zMR0xqEeDo54nW8LRIAzAtDcfUvrsLD/7voErVnEM
IlAW7VnBx8yAQcuGHcSenI38bXV1cczxGKTBmR63PA3gEXVe0zFPw/cNXb5LO5NY
gBnTQNyKyWsiqgFRNsB7KuEXjEcqVr2IlFDNnSi5+utQwSWU1HyQBXZVYtsCok2F
IYR3LMBZYlV0XTfBBMtKWXOkSO8qqtSEysazyJSXuOVbmbXEpLw0GtzwONhfXDRP
I8LXUkynV1PKgSVpT2qry3B0RMUgTdi0ywzMED4MypaW/+q14MbZgpzE0bC5SMEX
3GJdPemYg7lNaNGw/kIQZ+1NGaBT8SJ/exAI/Crf1iBB+ZX88qauCldGhthISRT5
F4/VkoguVgYtP59U/gkxWCd8/OhOFioX91Z+on6ihn3XlD0UU/aHl/Dkl/bcOk8X
3m45xV21vFftXqqtSP3FVIKW+qZposEsoD/SKmFD8hZiYlpIbmGtITnLH9idy8AY
x8cY6hiaAsyI84L/ziRG7xH+WfvedHUaTezzBCRM+L4/SOW4YGkY1Y9AKu65xjHW
wx4sfEoTSRvMzJ0uYPxRFPF5LaqP7l81nyR7K/qtUqLF4Da7kEbWsOwWONe7SApM
7L3WtaG8nESUlgZ6dAFahG5sWMxLCgRXsB4wQ3rOlFlRdaXLtDF0h8s9GRTDQjXQ
cNLk9Nq59laavC7atln3b2Bhyb6CzG42eXjXtqUtUjvYtKI00Ps5GNEI8wM2OryX
t0ECKJUg4PsyDUdrp+Pun8o6ggn72bQVavJJzET+Ii9ZOuW3D8PXgyMjG62HpwZk
6hJajBoicNMGTBYQZUtXrnko5uu51epX3n2C5pGH7jRIwTOxve+uqNCtQaJUtpiL
04OtuH3pxNQWK452arR99nH2eVFGZ15w+jo7sL33GhWhbwUnIrio/bguyen17H3n
uJfx5eDtRRknf6E6UMqhC4s4o5T4xD5FED77HefqDOYWDTxYajZns9cI0gwrDt+h
t1Sd7aFA8OAk6ET9sRSNVlGJeeyaJRr7COOLwUWHjR8XYRVZBbGWEHGAYuFZ/6W4
8A7BygjakYgklxt4+78uQRJ0d0aHcyZcKeLp8UFPRGPuNpYlri2CAhOG1ue0rFeo
eP7JFp3DKaR3BXmhDEXz/I0hxQOVmL7e3TsB4cMSqZ8mCZMLSmUvqvYI6zcK2K7r
YMfyW6B4CtcYqWsDs1TsvlM7Aa84voKuVUmY6yHlf2+11cpLqakQjhLxIovVpJzq
l0w/lsawG6L+XzdNpZECmJqyIUR+dx8/2FWhiePKVUAJlBoCkAEHOw3j0UJSqbV9
9tlf2EfaIDdryEonWj0U1lseNmLeNy+Vm/yhlWhlMQHlVNHZ2gpF14eY51/sNpuy
avfCyHTt+sKiSy/A+CXAav1ocxpbdCxtJEcOLSaULQf/hiWa4kbTVTh44LbQ+X6K
9hfVVqPu+ME8l9EV9acoxabRcnGj7taNgYunqXduO87ZtoptQL3n+Hc6Xfe81OVs
aYQNPcMzVzTSp20PEL3N1xSDkdn1Vfqd57mbus+MsMXMWgt7DlD/XNrM2R32O0tO
EwutJdS26UfM1ZwhBeeBvo5QjaYDNoBgPRIy1M8l8TnGZ3EOn1Ew2KApOAD3yhEK
fTXJQ9RcczpjEHtvsNJvj+wu+o4l0Mss8eYbP8nRdjt4bmr3AunslD1ZiI6VE8PN
+iX8y6rg6aFVB1p8hc3FvbPiOuRHpNeixSCDiVl31XUPPH8UQ0wnPUwhC3bsuvXg
O0FQI73XocxkIT3oysPMHJoxTzRz7Pwp2wGMRXqfh3FWMhpzqXCEOws6tdot1rQA
rgAAYEeqXr7XJxv6ch0NIfpWX7P134U5W91QLYyO6GuFNLIlOxG12cXOgpjySGM2
yBEa0fT1/G72TpDNY43gYqhAL5rNxY+IMnOSvpjydg7vTIvU5WeS1tP8HITrK2h7
8oiurRFe9qnKIekpCzE/EhNRVXbpsI3IVVFLPayKYLFUQ5nYQbS2V6JBnk0KNdN1
W67Zxbtj6aRMF8QwMRg91kShZtdwNKNLviGzRvAgNqbOgB4DS9tDK0o7DzlRSAUe
lolZEU3zgcKZGGNUAk6Uxrw9DnN6+eqWcvhAIVNZ5KS99CepiDh7xrvimjLTnfzG
JW30MRPmcy1pzioJXMHY0Pvyf4eHAOjvDeCwIzpKrGtEe3PFwKZYsfuWKznWXR1G
ddKwFLkflxa/k2cntn0lqEbmYUAXRk2f9wuOVHKCGF6xpHlgCZNooFFIU+dETDtS
xCV2awaJrBwp9Ye1WhqtA9sq4qxz/jismO8eYxANlz8ccg2RoX0G/zNd2notRzL0
VglaUTlMposwbPR8XrrYfIkIHrTV2Ey4eeyeieBf3Mrii9yVovyXnL6BjgzfzClx
FRMnfbP5jJauh490gJIuWAVYScvSXqZYWxM8YyY0oQ8BKU/zmMxQx0VBIz5XtW7z
T3h1hFPtr3omVbysbcxspoXCAevMWN48LxFeN46iBvw+xZ8a8tHHKzfPi6AHuLU7
vNmr7B5HHRVJ6ec8jn01u5LJSdwQe8U5qT7pKU14qlBplpV9Oq6Fsu5WTfjO00zZ
p+xEJU8P5S6vUpNxCB7ul5KtsEndma6s2X3cWk+3gBLrex9vR1GRamUkSoMFCjiT
O8hIUV2s7CX7RPdwqto9sbLmjOSClUZv0cifOttP0MtVXZzQwTPebBqRbXu4Ph9t
tH23zqQ0QFtI2W8IEGCL2Ixw2207MXwtWDrZ5MwXTumKYXXQm50pboaIgzxf+r99
z0b7UnEm7k8H1t57EkJAQ2xCM1WblwpVyrxDyraHki5p6AjyvsLgPxvVYH9fu9Qy
JezgYc+ehDtMBv1LhwIn+7/3bJi+4G1srxV+i8+0KKf2em4CqvDgJLJJ3EmOJqWt
+mLJ340t+A4F+w8kW2MPaozKzsXy1YlJ73gAnTnfhjZSRmOl4VNEbnIuhjiEFQGA
O/G96XduWglRxlYL6BsS6WBMytq8fvutVka2Fl/KPiXTvJLp3IPHJOd32dY86ggq
+/l0V7cZ05dclDSv9+rIZjKTovVPmV/M4MeDxpOlyw+GJnaodB8CwDWFMAHs0rnw
GGR4PrL2TmEsxah0rmfoIK6MAB5Eg1AprQJOlnGFtqQIV8w3JzHsSDETxNg3+A35
/2icF9QkzQEqxy5lpQGaSrtDTCdjS7PI+YjMRMvPa2HbbOy3x0Ll/36uE6dy08Sr
/syvIzkbhPnotEpAbZPEhjIhzL6SI2epvfDV9vbxnXis0RbNWmrT2VtWlMoM0CPH
g1UWX6KBwhkpoONv8qJTFH4JSODH7/SceFxmdlc7Jrrn9ph6ViBCjQgmGe29ViXA
KS/LEVAVbnXMRvrw5RU1Ay8uXFxbY7VCHSrSaA3GRV7oXbmIfQXESzpSNt8q1t8r
PzBiBYKH5jk/IGIetakYA3JIWrr07JCfBEs6QK2m6P5MA9Kd0+DanFF9ZpHIVlNz
mrdWADxOUPCUXsalkOPR3+glhFWdOHlspS1Mtd7nxwjazJRd9NIMKlWBbA3ewTBv
UucIANjmAe7Cju2Jbl3ycsqYmdRqomncynb0E7IKOJgCdHkah8JCkvLYEcg2lMBO
iKDl4p3k5lvScJP/gTz82RoDwNT3PhwHXGNEFeTZOpNdHLxXT+87UUYDo4fybch1
slSPHT8k7L8pOMGZCV2MKXet5lIpHMDOipcii05ig2jBS2e5t9oRkjdW/fAWCd05
SBQKACBvPkIcCc3/OW/wTsP+isN7Y8r6ZTOI3qIUfZAvcYfw3bGoyYFbISGfZanS
uzmbZDmYOhEyVJVM4c3eyDfBXJkVjxs5p1sF5o1CEtKUgkHmcpRIqMJzGDUycu15
3Eob/YNIkJFq4VfOVnvcpZhfcT/YaPPE68VSSpxzPrDD193CutxSNBLiGpl4o4m8
0MDnADRIu490KupXjM2fKy8YsGp3xC6yYQpBYnj2854eQM7RWI9qsPK2FD+vSHaB
+Er9XkZoSOJLXPNYetabdfc+04AWx1S9fbMI4zNtGIZTEZibXDfqgsPKb9M6MPEg
q2TndSTwUxjmB0cFamRh6TncTgAP4osEoulexwmpB1yIG3iOKG3R4WuDKdTrTFsu
pFti0+fVr1GqvDa/FmfoIKTS0iOiOOGHXUDMPFqLglVkxMsMW7PcxRm1lyflsvCr
MG6nLMZiC48ZCbXCXs6PlJArU7CMRYLS8U3s1UXVyQf0wl6Bgc12Q4403AV9B8d4
Y93MassFGLkWc9kBdZVFrhPpnn+dAYHlqwyznDwOWpGVus+K4OAijLGhgmlIapT5
oy3rZKtWoyJEs5MAs/Fa/KdO1PH1Q+d6AElrKVZXN2zsJVOZl3kJpHndzmZnJR4R
FtScUZ5+AhtxCRtof/huQYo1B1fSnQuCBkcfSl0emJ2fHo2808HAG2OpxZTcTUlu
EQeDVQ4rsqy64d1iZh0A05nJJD6Rpjv7Plgg82gZr/NUTvEyxofRN7SesaVGZauD
/5I9duoCPjIIudAldLh8nKC0gJyjexat8Tpgxfv3WTB78zeUdAic3XbL/7H50vp1
bNVq95o1Nbi8OVYLOrNan42+8rKsXL5latEG6QSYYwN+eC/D7osFW7LbU0p09kuo
S7FRC+MmfabUexXCo9JPmVGJl8pDBOz8hwZuVBrqdFym0NlOMPZKbl9uSdoQF6nd
reSzxryF4RVNPovZEEBX8J81xMoghZxra6PQNsuVkvPQY7L35zXqdOX00PXjhAvt
PPSQcbG0L3Fxlc8XvYNKiFMeWHGwYRsPLl2/UDX648gDmo9Q0YTs91ZC2KVXHDTC
q1ZS+2ZI1s5/p9BJklQNYxLKiLovPf0xwH1GLfxI0O2zDzodXpyb6pPu9XCMyvaw
Y05XFc0bTK9FZ1hdss12BZjlkFL1JqzJKiZNl90nJ9fX24s1B44pUts6M8XgIn5X
HdSH8rzhW0RO7iBNxZuOWgVJ+8YfctroJF8AgKEzJL3MyZWVlCc18yR5EYFHtgbW
G0lI74sbamEdU1QrLZQu1aREZIDh9EptSD2Tegeb22U9XYp50pFvBv6I96Jq9aL9
Ar6b2eivyopOsBEtAZmtnn+Y7sRGI76OJWrRzpIcm0oeAlxcnDt95LzmdV2mMk8U
9/y/M5fv4NJ0epkIJzuK2SxmKuVutoTTB/4u/25Rk3qcWHtxPedVFco+L3XfL5Gy
fEw7zDqn3uc/E+C/lLly/0mB2KGHrAL7QTCqiqzrA/OI773E1yecgnGmMrOGHum6
Yl/do0tU5bL4r22teMAqQGhKHPrE+HWmupAzZCT8jEJAR3vZBvs6S7zYKG80AFP9
lbqddRbLsqW0NPbpvzvLtNE8/rtutMz4Ze62bwZ8RQmicSCITYB6n//bxroibQma
T72cFtoEtZSAJMxaDnyAMbPFZxs+fMjPSJFwjNZuP6goovUQA2V0A1DWE54ossYp
h4hEBZKXBIZALP0LIjyWFGim/kXHjpF0AwRFJ4j+MC1yleQaWAElcio8TBxa4W9w
9TknRxTdrbp5QyIU8wYIseLvfinPTUatt4WLvZ5rIiDpJBHxK79jwDCvANFvdLGk
qsl4yO/8WsLIKLoNfYCnDcSWNLU9YXYR0Xu2nmJB1ZAsv5xs3AukUxeov1zVZ7E5
YoQpzGwpC528OrbDfGIKaisL7cyeD5GbPmRoy3cQmM+3yGMgcnem8OY+MjtAiTDs
ttOJl0703xJutineRoKKB/kQQwMAIZmgxOmsneexZs4IuADOmyGdyxTxjiuP00+5
gPIhAPNplBGN84lVODdwHlc72h6nTelYsef3s9Dcj2Yw8VrD3BLVn/CLa6SvJOGK
gTwLfi5wPdV0HAMIG184WsprKhL0Y03EPzMQIJ6oRCQaJonVD/8pU8kcIkstkzR2
7INX9BE8jY2fzR/W4O+qvyIG1L41mTd3SPrY1YIM4hR5LC2B8ri0Jj8L+6XrcGva
8GSQ9UXDRwYRWxz5UA+Qv91h5i1cDwesBjY9MLmRai9qQOnuR0QLFx/sIbTudnUy
URL1G/ui63kL6uv3dVmP4OKVvdATbn3NM01fsk/H1av8NjDdN+MPCG9RjBVSGqdk
s+WSpGKzReMt8YA6GDnnmiiXBULWjW+7CDBRbY2gB5DvrevZ69EIq8JMkB8VkU/e
JPBSa36W1QTrT7dUPKwqopUoY+LQn0LNLtfTaDXO7JtzcHB4+sqVdOoQJIkjxOx7
B6VomGqnS7kcgOh7pnNX7mqveBk10kWI1qz3iRDUs8iN3f5DW1GiHPYVg8djmht3
qaNNHYQD8HtE+/h1uE++5izd2vYX0rPn0UPWjVFG1I6Nj/FguGEFf0wqEH0YLrLF
XVItYJ32A+A8mtlHvBf3UrpqiVzPSpZLifUNmeXfq9eXEPuVDxqs3Y2iV+Qck0+/
zWEMIVGLUf4369Fd/RciiEp5oqDKwdMe9pC52c95jlqHkRY3baHnLiLYdwowQwx3
Xzt8kNubTp+/yuct+al/gPUJoaYTLcyS5YRWSYkD8jyGS4jhtEaMUAC013/2+GyV
+/RFrXyErwjzLoRVNeSbb9q2GvbsNs6bjco/ZnXPE1w8IwwbBI9nm0HSHStYifMO
UGaEF2+8yHDqwmTo4rsWRWMqPH9BrSIyMjBXbcjtn8Ti9VnUh6o7cdUKXsGWaNgs
+MwhbXkwCtxIl3NMca52597/LRHrsfBrDpk+c8ArZHUzJGwlvc4uuKkNY7uMkC5E
QckUruAPZLWYNdHwXrO3YZJ8jvTW/CbKkd9BoG3lM2w18lhl1O0WY6TFp3esKldt
MNMLBqlu17+8fa4oJQkosGoT9IQ2UTzmZ/8SUs5xzjZ+ENFlDgIqvpNKutHE7vjG
u3lKCyN7X+nzjnXvmByzW/C5yZ3qYoNE21cItN6ImC6stcvccB+/BuAymhdTJWsz
IlgYUROE48rbSjvJW9bEdWc1D5w8YT0Hq3w7Y8ocLS2gA2bczNw+VMOhqVlrBSOR
xJN4dIsKvkBqnmAmlqir3VNEw4PUbDOL9FsRnNX0AygylRX5nsmb7pElePfVNv4B
YC/E4inGWIpGG7KFFjHVaThVD0A+QZn8gvfmOZG9fVj/nWVpd8SywAAIY0NVwtr4
UfB8hEw2Q4u0hm1ckUugtwBgRUMZvAuavE9UyMtDyKs46qcIYxWW7N00JrjtRf8B
KGT5egsratphH/ZxnLvPF0+ZhBKnToQqlZFjZko8S4k/m+KK9JfDARu9LqZDIjjm
+hlX+kNFR38mAByT2LYujz+KK4rNB8WACB5coXROc3+EZOmVSMZ2Ej7GRvh5MF9Q
g9/hXxAcDBwdpVhHq+f2Ms/CC2S8UYH0RR96ssDzwr3GZa86skWpq21O012R9UD2
JCvzHIxzA01V1+P4ivs32C9C6UyUaV7iUo9kydAspZlcDzVLJQZgaJF+peDU6NQs
oQGgM08KToD+0M7b0490PwEMTjsBfVxf5wbYGL4gdBsQWqR58sfVPDrcng8YLLC3
tbO0gPINMsWqAPNwdb7W6LRO8sly+C9li/5NRmxssKQXxIsGrENYPX7xxpq5faN0
Rg/K9NB/UaEDDz62lrwm2ilcia0eCTxX1NXmbsErLNiEzehYu3lpAl9J02uto8iw
nFa3HPAqsxIPbNSYjuU/Zz8OZKEPfDlG9my+6A321sL3IaNGCiPqk3xYMP+diBwf
kUSQcO4wYuRhaZ24fOgg0/lC27XnGqPMjI9/A0NfjffSiToawuRI3On4I4NbqTza
2nYrmAJQUtvNAGmCni2WOYDFcmJrlj4WcqshiOPt4ee3Tq3CXoZlfPDQpHDxFEgm
8pcJWNg1To8UJKvrZen3yjN66qFUIZ9+dDYIb42jp/UOL1YCeA1Dq82ElGJ1ny7q
e8QQNYv6Kq4tpdcGuNbkfuvrcLRGigT0aVGKHVo8xErlMFIHdO8OKTwVPbF7K2wO
QigeD62MAXN+KdsNui0QS+3d4Tg0eN4GAFwpEgfj0PC2oHjfpIkUPhu0UZMAFMVt
UGHR6FSzNOmoDJxYsIqVyEwE8wXFEiie5OEOnK5s9R63vFTiMa/TKANhuHUw2T03
TvuK7WK69OGugtRTT+ghlA48FCrHrLnPLYNcQDo7B48azmeuZ1ovML12XIA6seWD
rkIioE9+KqHDr+/Uxt4Y+iMjmg63l4LqTKRT6AvdayFAq54uV5uAO+bo6XA735WC
02h7DNZ6Q1cV/gcZeYoKGMIGdRKq4sNuoWodURSUUTASI+qlEqdkugLSxOM4I0o9
cZrnw23Omtr944Kq72xAW4R2cpMJNMHvUeKUbGMjSbYy/nf4PLSzTbP8cGhx0Wjo
XMyvV4LOS9LrE4bd/QJGDm0KPxNcnt8gK+ZhWcEPezqWNyCU0kzhDtLGnVK5FuNA
jqErUvnZPj97YZkerbe/E4zzZcG3rgjUq7QHrB9kC7sDlX2ykFR7tsrX797FpsbF
yGZts9e4FiJGbLRKZWnz1BILoQm4BjbKx7I8oufPDuigV+g65VM8CbWVIlTOKj1X
lNjvTn8eI6pNdAP5Z9Z5XP0bDCEMTg7l5UmOjcuNovBG8/IKkv2+LI4KqtY7TFuO
wGm/p5L3Gonfj9LX9F2TOVvxXJt8eesvSI4dQAZ1Ych5kqlJDBgCTraRq6T9QRG+
HMCbwOOVkAoNGaHlbK0CHb8ww56xk8oNqpMx7gvMJxEEA78OsfEZ6ZEpPSP1PYqc
jLemeRSRlciGdDZe54WNXTid+w+AJUUiEpzjXwC8rjY9T1jbgvCMTkwA/PTy+XVZ
vKDO6liSzVT2/3NYpe4Gb6TVdpD/eFNMG10wDoEcKONGOzCEU4wuOip632GVYBc9
U5yGEILeTPoyoicW3UrS6xN6QM5WRTONvIbWR30JeCVndFgDalX8rc/Est8m+elT
p7DYQO0g8dKieUPUs8vTp/zFUsry8TyE8Y0K95Z/YhTxILo/oo0vJfSMmGiGBZ9W
e63c5a39+K/JNF02Je+x9Yb8aBhcOHQF2hBRwcD9YtpvyOVEQLK/pgj7/SZFsRAi
y3cfGSPWDiWwQs5ZIuEdo/waXegT0P/d0NNiSo6GrdCNV2P83aduqYwsEMDvUM7V
IyidqC0YxnndJSaMN+rUAQdBNWmMvlbrfkSAqvurOmuPb5jbgfKtbQvN0+AC0TPi
tpJp0mZaq6i0qY7qJqWuLrPbt0GCWVWKOrft4RgmqFnzzRiKE3eXxU/+WLehVoOB
4JLMkMWXrc4ZPywizpI2iUjjywpC8XATSlc+oGj9u/YybIoVUHp+42Jj5VBY51bq
gWY+guOCDZrO9hZLGdoEeJJ/I1weZ1zlyTLz+aShAslAFSn5EEMGpvuTvifQqnjY
Uuhgm8RMxY1BuSL+4MIiYQO2U+RYePqNrZIptL2fXCfcPXdXK8CbkumOHQKy9Lhc
b8mGWMAxJLBu3nk0FIxf8wqhJnhidI3jTK+Za38SAAD5hXyH0lZYLnlTrYYGOFtN
Ayn9avKojsnhtGm0/ycCUhe3VvmDR9aD0XZnN3o1lvix8S0zQtPlyATI40DnQqZb
vbhhK+HH0+coapDxmzucq7650V8J2DzjIKUsoBsH6hayBRrmp7QKLJJn+nxvIl77
JKkVMmV4P7rduEF2a+QEFOWyztWprID2ynxC4xGUlk6SFPRIQlbXBpKtrBjRDk27
n0U+z6uUL0LOTfE/MXAmcb+AHcO5y8wZ6FvvWu+MpqOaRwdlGTtREJc//pxOfWFf
/DzyyjLchnb/iEbegwGjFIbs6p35y8UbNfWBv4LNxV/z7Wr9oXxXonuyjAQDL/gq
zSI8qD/P1skaDFGCeB5XLr7tP/0M6Dco+dX1h/ZBLZcNfzFx8eMfPDlU6HpO2pL2
GPZeV6eAi4QWPFZK+swGeoxmTno4q82RI7bUNkdt91iPafVBUaUH3D27ZiDlS3Qi
oGOBBbSlcFcLK7mMpjf6xBlDWD4Vd26pxifPsA+mR20WGI29cufMc6R0/X8dicUz
oZoXkO6OHWPT2t6+R5DieDdwD+SR4xJJjwpf1/3HAOJLOhTuPSAo7i7mE8zEbYm9
AwJ0pi4OEea/9BHUnyx5Ht4brqfbzXtdHrc9wmeQVJjQ91VxvHyGYHd1T7GMBUeT
xBE/jR9b4DTx//uFK4W2qZjWRz8thxjpykcQvkN1+ErzDoxc1vlaeRz6jc4E8HSZ
zQ3MmeWRQ2KBvGr8/HFS2bsnKRgQbmNj2IBtZyyPNdZc9G9DZkwjuSfb/Kv+6uJu
iSwbPR6kziAITwxEWjFzfdl/WRYFss+DJ55mA2kjUNchsoNV3L67D9a6URRMNNan
g/sk0Q1qOZaAvqUtfPApjZ9i270g4CG4FdVXFjldARxF65hhMvVeEfYXFWau6X/U
Iu9M6sH6RUeCXU78cVkLGBEjHVzoM5ucucjWoiUI8GWXiXc65Q/b/mkmgwQrRMFY
OUg8kxv8aSfPa9qISrU8O9P6AJNDXal0K+DkameRRaq+b8/bOjgqpV34/LiK4Sy7
mwOTeF0V05vu9/EYNPd+UiJ2zomeCEbjookjmm8BLzI9QLkMKc/qguHwVWIQ+mxw
LGj7dTmges98FtyIl865viPuTN20SOW9derCo7aTFKZwLqYDYPz5d0bgLxpE7Cx4
E2ghS9qTTFOcXI2/lr8kFkXa6wYGGALJtnUXJRIZvLlPEgxogAGhcKqlzGSmCXy6
sgW6bGqVJ3s+zIgKcoOlQUlepua214cex7mzXikUCx1cJyCESI6AFyMgqYJT5/dN
gKPLtDbBlsWtyUDB2gNcHJ97aw73mkK1FVyGN4vNl7ve+QBMjusriwh9g3tzqDat
Snyjwneut/LaT2TMSclcbLfF09wuwHNoSRQHS4Qs7WYML/YAz0KiKqmAnzU9Vlky
ZlkiUtJBcX6Uzzh77vw82i+ppfljZelRzkU7yoy+0RZwZvdBIoKx3tml+0IgjrsU
SPs2GhWeejDt8ET+FcW+LcKxo4ob/jVJtSzIEoHtS2ZJ4GrCMXQjBTCawfV4thKi
M5bQ5YHYu/YZvrEZhVOQknW7OR+/54S7+4APckjDtM1fEmXMxLbsaHkquYnqUK+u
/ESsa18sLpPMdGOoH6aKrSnJK8kn2FXgpNDrmoCva+kqBGBoQqDE2m6PR4qsObRK
j159Yv7iqM5npC8AMIZRKpqH4kHxhsA29JWl+YTHCCQfQgtEL/iRXn3L83cDZ2zM
9fF89T06JP/h4iVwKRf7NzXFCxSd6HMroKS7/asMltDgRYC0nBp3cuRvf0k8zJ6W
RNm4CG89HsUzlMU/C4a2kmC+B/vlbWSN7KKpZk5xlgjoZF5sW2gzoyLvOowaXoV9
UGk7Y2CDKw7so5NvPIRCijvD+vD+w2vUlnnqnLYwmI0wvkJWy6MSV1JbGJnCA0+3
Kvg19jlmO6bWTgh/9KQRjTPNHyPPiDokOqmzZKhT+rF965zq5alshme30q3A/hKr
RXW6T/D5TuuG1p+jVyZQ/puphntdSc7CgPPf2ayDGRuMow1FqHGX0cPcs4+PvzyV
G96cPy9xY897dL1b2do4Lgt+Yl4SC6cwEQJobfM+GdhrLhkTk4u2reTqOA4KBE2u
td4hLKxpWKlv5NKDgNvStRlWcnBAlVy+K1+hkX5T3YTgHIjxYAkd6teAD6oo4hEm
tFJrKGQCw5/1Z/QNys/XAtyEeVpgcKdwbnww0yxvHWHhBhIKE9teFotuSokrw3Jf
gR1nKbDGrY7Dkc95bfFMVJu7mCz41p6M4iohdVo39WvdpPoWAUO9Q/UQ3dWYQpsb
w7up6gfpdz80rTSWJ8VjHdWiPyAYIcL61Qzur/ViaILyuSLbNnc+ab+/RiOCT74Q
Q/eBk9YPEP+l9ZZqQinW7IVt3g37dM+29MWKQFSLaaZplU39JqFJisN2cxzgRC7D
r13oTHM2UPUdYl39FFqMdxyXJ/pD1ee5DqSgxhnCiVXiUbVAbcyuEKlnk3HEkxkv
HCCp6SvDE35ny1i8Y5H95WPTHNLF18Q2Fel5100ToGb7WICVWZTKVJwjGGVhQbaH
NWBk2B9veCVhIJ/ikcS88T6HiaVZVeLXiXsr6Q0ALtSCHo2ec7Q7+pyQQCns8ZMS
KS0I1ALxDF+g5ZYH//NDuYjI3/PykBhOSFY+YEcs/l031++He+hCzZ9HqZOwemlG
qd5RAgUjs65aX+UVy0tFiK6o/PbQQ32QyX/OtIN9XS6kSlHpTPoQNBShS+yU/xYc
a/xzyTgW6AqVK+jEfNSUsGk6RpK+A2NIC1PWTiuBxRD6OqyfjIqtN7zicu1KG5CR
fvG6g+voGJkNA4UOHKnZDLpJXAM1OpsJXWB3rN8YFS8RVNJEd5It1rUJIIB2psMQ
wOrnw23s4NnDcPw54FnFXMQFdqXJoZDFEnRLz9LnzzLIo9m/8X3O5gmGqO0h+jKi
gMejlGj6pQmcWd6G70CdNgG5siKmTlXO9h5EW3C6gK0XVOAUO24NYt8vJCxp8RQF
xu9UrG1DwqVlpI8ZJdEUtd1nlqqdXETsbX3BsBMtZFf45DG0SnLF69Ma+WV2X7z5
p4TfiCjOHt1rm4iEvmOmqGK1qDxzfC3t+0BiYKZv0Z4Z5yUkKMPsBsE6KlXZNE3u
XdRZc/vYKr9ZJ/KDIOVwFrVK+3fKwQlpSg61R9nC6p6aVbvonJr/thV07FDeqbG6
x2Qji1GL92VANk7bhw0oBhf4Zn5MDJ/bpDqTOPrJOqbTMSzEWF2kOavQKQT+lT+i
ZtBIGRnPwJvkBv3r5GRYSvbh4+SvsZlHp4Z+goJJGSHKNYi4TDix535EMrHa+LIq
5/ZH7HtXi3xzlr9B45V9Is6acdEjHFJzIzKHlzhMWE2laaNNMKdodLUU6KxtQxK3
aCReZwgrGkvsJAkXkaYN1gWBTTfjS7bdK+LRab7gEGD4BKYVOIr0c8ZKCcY/WV+C
e/mUdbAHmEVi8f/lV0n+1L1yPaFbYVOHHwrm1b0zccz/sflM+uosLUf7lj7Hvtxg
yZHGcLefFj1lKyFxuIddGmCFrOwylETOX7xZK0iEorK4RmwLajb8QGJi4fIjF5Gi
FGCs9v+Mh2kRCCbz1Mek72MaxsKG7rwNrTkD8xPlAB4NUJ9Y0JvzG1zM2rHDbmCL
RCSCH4fpPfFN8hJj1/QvCB9uO2Az9DyhDPY6dNBHjTqYWax1o5VUGQWRe2vdYdVL
SyaGL+31kcq3p/swREjIOkMgnO+PGXpajMkl/pepCoEfvw4bYrYNTn0K9q7yKPZ1
o3y8ShZGB3oM9wrvEOh78A+LmHKqAuNrV0PK8+s/Vo2EWhzme+sm8YkyXuPNo1Rl
jMjr6xioAZUjjEtBQcBuWSKHZAFL2f1x4Ia+y+XLbCoglFUTRfkgs5DJJMvO0Dxe
3i8jcQa6bC9JgtqBuVjiH0u8cb/r0fYSG5tkP3Gym35KrL6KqP2wOas1ueM9SGdf
VM+5RmgBQuPvZA4DxbLPRzJDMN3BsJbPkYEl7AZYIgaJ1yJxRxO9awCqFnKTiDIZ
4AXCtvIHO/67HSrPxOqkJKZCC9HcsUtfzqYYBz75mNv16UhNu0UEtAWVpe5q6zv1
b3MR3Sp4AoTFfcQYk79CvtOaMmTIJNKmlzbcWNy4B4eKH1pDorypQiDd9xMx7BMt
sh99xycTt+ozWTGO/nkUYT5i6/OqihuV9JOCE+4Y0hXMvHZ5rdUUi30zvXoW1iKm
QYh4Zx0SiEoHGNdSFnIw20lJp9bJsBH3CYj4VBX15pseQvlPXkfln9AM34Kma5j9
hQ6muqowwAE57Um0YquztLSANwAWByhTH/27aT0qV6hnyh/kb2S50akc/ciGGmce
W3olLQCmEsJPfAYkxZghYiO4XyyTLcGF2hf0avkCztahnBTPo//3wYEtKS//QXDR
X2RV2U1yVvdpnMKBbkDSwPP5E49NFaW34v2E6jnYvvHYJqNF7+5UAOnQvLBmq7yD
YNgSgrteBpoYiHVGIRSm3y471RT3mXGG/PrbP77ArqgpZXS+nTcbGStw+ogtEGDw
ynyUD61cuuS31+WEbtXB2FXl1oY4Dw/vwbhD8MPFnTc2VzYOd+LuOcOe8QOBOTWX
0IbR9lhqz1qpl46koUSCIvRCO6b7e9L2TDvht+e+a8IlBcKJEpkCdT2Iu1u0Rzy/
980iQrYSnCWWaJzEobFoZbEl3reFK/3sgkINReSDHpES/UEbB640l47sMwrIgoJI
QaLWC3KUMp5v887q87P/LLF+oU4lUWf7BmWctO0bPWBJb1AZMoTeBJX8Z3GSirq0
/ZD0KSFHpPmozIDvRc7nEKcWVnTDzGvekpycnBy2fwKV0xZWusx6nQoEgi7LZR6s
2ChA6P2No0elbSwerJJvI3su8Wm3ITWNEFC9kLPLU5ZoIQU6w05fKhz2NoH8NP8Y
1OXFx9ZNe9GnAzvUPkr6mVJzLQ/qtu/exifTWGCrGNKjrRCRkOyaFmo9MPHoZgGw
f7LjihLZRNRTjb2b0luiz+nRe8UiwaipLlxjEJg/SG+q98n/P84jwnHHwKuJb7Dw
XXPUxJpwv7KfKMgZEQ45ziUtFlL1tw0XMBOh6U/6h5h09rmwejlb/6gwOuyUmWsq
4TrfOmU7cXve9yYZulX27OCc1kTVwSKtSFyn4JY9JN0Lno7UBpv5055aGl57xL7+
XTMxoXxpalEg630ioFbFRsuWtarUpnwdKysJUjiiCKJXRdVU0tVGVcWgD/Dfp6TF
B3nB8/jp20yN0PcdomADeffwhQBleqL3hKflp2q8eq72ZwtdnQ9d5Er2CHhljNMl
p5GYc7MUgn2alodAy+dK48i47umQFOSwCuqBFlQk+AZaC5c4wavVIpbJyEePXt7T
KDmoP4qiC7xLj7wVVuwK5nF3JPbxQ3TiA/zcNmvLZNpUJHelkNYjbMP2JRG6UR0O
+BPWap5HxhIrZxkfEJp6ODLwdatnxq3WW3mQJUvZFIzr1Zv/10ou9IMfz9eBiU3p
KD/x/Z5Rw2aqNi3dqnYFBij+n46RAOrMdI5YK8py2PQrSHBz5sKBA1T1GzygIRlo
NCbTv6q/rIO+GiLMXrY7+Hh+VSh0TRKqz3huFzKYu3uav0CS+qn4W41OAP4RPoUn
sdzHRKscLoIjVrBVjuAfaEz8ScMTvuYepZnjGDYu1JaDquMGOepME/34P7TC7Sp5
IaJH+plyju/mqoDEgFjC0qIYnRncL7ORAJTmW/ptq/ZoeodOdA60274lOCWc3pQ9
g+LARc64vtQiXzzf3cwB4nAhdm7crWH/LEvwO5hfekMXWt9QQLzWP8wGqTRKOqcC
4th+KBcQOQvfhccS8f9FZm+YUNpjdatmC+a3NsuQ/p2LpT2Oc3o1ovW7DX2knrT9
J4oHSIQwgtw2pdg91QXwwxMN8qUEOOdYyeGT0X9ekUWy4V4u82XXoiaJeK3JTXST
y2D4Gnns6cFBpZFdLv4axWjXtQMMWGb+VAzfAOBdvzIxuaNkdGyxzyqdaUZMpNn7
8BSCjs0yGoYJ9Y5Lh+ZYpB7UFaBKl6Fg24T6doQYriKGQ1pHiSnhkzfEOli78zg/
49I2xKHZNXKhHEf9lg+GiKy0QGXxnIQEyf0xryAmsmS5f0T/o6BxEQrzj7d5YOnb
uKIC8QKc5qc9rDPSERpgIxh3s2dkUIvFap+fDkehO9dwF0CuQTR7eX/+V9D5AZNW
12Ygud04yn6/W8A6I2YIivvB423+ft8HnnCPCBRIlQVxu6WJXKE+AJoeHjClhE6Y
m9Zj3a4bVISkAQXO3Hhj783BWI67mEpF73t/a+AdWlnarj0dIApispT7rKTtip02
N8KRqJeAiEuomRzefsx285QfWkB9pC75xzxcKlMQu2fBlF32Lb/CF4/tMY4KNEHS
ntXc3Y7qdHjB8guQ0oOh9842CjxPUwfNvJLY1OS2s3+4G4pOJuTz9UYGf6Zo7UWG
xzcYNSzuPWJ1McLgw1/fi6vzRUWObDQ2JbaauTlh7xr1JQ198O4uW0UVVcSsevQE
7NFeMlD+jnMQ39x37cok/RCsSJdu2mcsk6XiYsYiGEmu/U9GN8JGke/goyRiObOP
nsTbY4m6hk742gku4csmAWFmoYcyFwYtuw4lTJv2hKNg368YEhKPN0OsywL3C+7i
5+yw9aORM4GHe+ZlQCT9oL8oaZC7ZkoQKSLI3DS475VYZyaUp52Vvdmf9sOr5tac
q+ley7+t/wkCLPcAf2VDEvfhToPSBTxaP7grSX7eNtwfVjBEfpLV7mrhXBnqBdhJ
IkcdQHr7EknlfWCTKHeaqUkb/6snQ7oxuuVa3gIqOdHX2SOHBuA+/gPApvDgfUYA
tWGI938RPG9BrVXzp2H3jBEHAOHL9VVCFFPeb5CeFt0U9M9nRQhfZGU/QYAPbcYU
Be9m0HQ2e7P25CxpbbTikvIwuulTmstnbM2mEM+8F05jJTYGQXSgBx9HXoYkZXc2
ig/2nulRD5x/EOHmC1nA+xkb+6G07vSt0bsyWfcKQDp4sUo8mAQPrFF54ELFYYYj
QS3fosb0GSLxgO74M8X7d9zEQIAi3xw8X0I8u3C1k1LhcgfEAbdbh48HkO6nQsFX
ofJm8bfyE6lW3N+qwPVJgNMDSuBtrtEs5aoYr6kLY57QhcJmHxzf2y7F1U+24me9
+D/wLSRuKnWevwpuTPKQ7f/hso797rc8AE1Yk4/pZGlbfUlnWAY3KryRGl8+yixZ
xFb29mtBkY76t2s1ziWaOib4tYC+rxXHXfjh/xyYaJea8F03DXo4mrl1VvyAn9XQ
+s3H/2Bp3qG2mtq/5qmsaxEbc+x4ud98tP9V4XL080JAAHr7mM8OTzKrOd/k8/YU
bf3UF9ZJckMvHfwlQvObGnqOn5QY+9bU1YLzInGNQ+zaG2CrhX+2fDiFQA9Oi+c/
NxPl363wScFh6pzHzxJhF63ykwrQ5//kclLiQPTf0+DQm7rZKvBWxGSryVXVndCq
cuAzAJ3HVXwKn64PvecUXuwsoRL2rKiEDyK0EiKlI33eUsLnuUhuI8NrL+06JRIP
xoDtfXvGkhCmw6vHXslPVCTws5TN69+Rp4rFw/aEa4dkvME66E/mAqRmdMhZC+g1
x57zWq9tsqbDSEm+Xgk94uStO/1LCGzeVUMliMbrtbEUXv1F4ATmFsY7tbWQmnf6
ZNH8lWBWAkeItjGZxWxVpH+1NZfZoM3pjyJJ7Djg/BCXtmrCr72eZmDu2qU45GVc
SXyur2zSPbqHogBM+DXN3SW6zS7E4qyJrP7uM3WjyBFssu68LVpGnDOiBw1y5+hV
YGNt0n0r3zrDMa2LmGv8jutE9KyW3Ylf6ajk9yk3bM518wyRWN9MxPSJRUf8uaNa
Rdhrbu8bb5zPCdzmqCvZMvTZPdKdFjTcfEIBdjQJAK3NCx1pwZ0nYfEEFq1ebvoF
T8tWAEnZSgDj5DZMu50f1o3hSR2OtyN/xXq3HX7briC4g2kghGnnuZzoLM0XOPhx
8FqGxijLPeHM3hY1ikiBQCWrQUuygG/bZpD9PSr01Z6SYIyQnaXHqDpfjKxV4v1l
GtKcx1Mh/pnAr65RHkfY+Y2M381QSwZYOf7KYNbVosWIRbS25DGh9DwRafhAjw+C
zEI+WwMZER2KxKBXTvV53oBc7aH9H/QIKtReewIsz5HCBKETl4yllxoBKhMMe/xG
TEfAxA+U0WXkia1xqD8gyPdiTH8U4dOKbGcv+0ZtgWf6WAnETmVgbvj5UlI16YzG
fVjpa2aEyfStrltHBD/8zGwRysvZWsIM7ipVEJWqbJAKXgeePElnbvjAnIZs+wBT
7nMiuOB5hfH3Gk4UoGP+xNkcqcsMzPleCq3SamhCqR9MMjGT8jx/4S8n/vSpQsYc
RlA+Tzbdd2QlE7BD1uBdwDx5I92S/S77HaR33xVjfd1/siut1wPcJ/E+bQr5cep4
cIHbLRMmX/bQd6AjsTt8b1hUnOoBqD9Gsf8y51Jo0g1Z5o9nSqTS38if/RObkP/5
vF6FAtI2bTVx0cOog9RUDPLO0UmZan36TSToo2Bn5zXeSuFwDpzYIbi2+tWmClft
gkAHtmnQA8WFTz5Okfn8lV2/XdPlQfw0jRi3Sl3SeCXpILWdV4qJNk8eYFb9OSTR
/DYcId2mA77SD+utAVWbSLTjbAJXS2UifNSc4m6DnVtFQJ5KsHRitJfHwBj0N2Gv
sxvnPAHEoiAv2oVPWHnoPfNITFrnY+0ovn5sM5iV2rnmod2T4bEgwl7dsE/mDNtf
jM2OTnxMxw09oXG+GYy0yv/1NbIeSUpuUkWaQOFA6GWqmJNCBh/vnujhnd1z5NIa
hZyBZU6k2BzbtSAUlZrnE5ELh9OrCbm4gBIL07GodCtZJxF1TyD9/Lqf+HyqGJmM
P6hmPzw6RYPDGZRgEKrFENeh64Bot/FkiXciiszonG+ST2TOip7gXtpnhDKJkvH7
OR3poqueyYdRfISDQkyvY5S+oYF4Bxk++aXxUrI7L4P9OPLlDVFlxvxYvF4mWA6z
P83RYIpI7MUo7jwleGn9wfI4DmZRMK+RD2/EzAEJrD75GylCGkbOGZe4OGReCuFf
hqVsBLqTSscXU7MdYjUOMHrM4ngA1N4WrxEQUlLvwb423NJ6UBhonRRgS1eoJXGL
oaQUb9mq9I/qXMRxvi2fdasXG702oJBienin6C10sepHgE6trc11u/SQvRYxsUxM
PDRRon4BScvdSDtmZB0oyKBjtHuI9LCHSgz5Uo2Xq64eTZsw2D7mwsSeEj4IQJNT
/+Yt/nPegdDjFWL+43Ao1rs7bC8UIDMPb/Tky98i6mVggRsSRw03X4wjxiRR9i7m
IQSbhN4Mmk7fKKUeINhjI3OuP6h4svJD4UOm2z+A6isSgcFcuezMdck4c/3d2Tlm
zYU0uIQRfAeD8EqFabGmtVjfyBQRNrCBmcvHkPmsrk1lplL832hTDPgfLDU7fClZ
Cv4SSNNR1WLPzcb+8vq0cb5meVAAgnTkqxksSaRK2JBlr+55zahBx0D4fEUvFDpt
+x7NL+Q8N4ac4evVc25/l0n6QBJqsTJrI47gv+A5pKwPk9Gd06iZe0ro372X5eW5
CefRCH7DcBdFNFj3oYz5mFlew75sgvK5v7L2USZ7zmzy5L2VQ6/erGnxUp9x1rcK
YMkeZ+ubkw8nQ8Q9hnnL0eHv+4TaQ+X6m1wNddqFY20X+hVP/cW/xbjq2fcPIfyT
xJwALyNZgAQs4cb5jysnj5J2Z0TC0MIMQwlRQYliaYlWh0jQ+YIR2dw/VqhgdJ00
m7Urbt75Rh/3LZO8Rb9eJYblEgYqowo/d9UIjL2MIPDhUsaPRhNh9ttXen0Vd80s
8T3H2N6whkcLNx/qgfV28a/Q7FxV4njRND5elZ/jxH6uFxpVQPrcSxl7EuhatLeR
k9gx76OPwR0TcLWCEPQEo2IZ9KJUDG/MKjUbx909t5ggC4Ogfo8nT2vwTWh0VDY6
LyCiqFeDWqv7O0E9tL5I3D+YG4BKyZwwd7nsQIhfDzQZIar09QgctBF5xreUrXOf
xshwxfqOdgN0iHKb7qFQQ3k1gzOKK6TtUr8YWhU0AsrS30v1tqYm6GSTQUxVAR1A
AAXjwGeYon8leq4V4ul7bbyM9gw+Ks8q5ppDTN/jHrfcinu2nlwAoTKxfr1DtyOW
MK3fnS8JNwz3vjlMBTp3Aq/7xc15XtF/BXH7D6GNwyzCnG3AFEHat+dGvmghx3a7
WqfLSzFxT61wwPg8y9nA4Canxe40b74GtnXUtCK+qlDYCAxvLQdzQ7g5Q2NaFlyo
nJzTYTnDj+ap8k+VxKgSaSiC0D4TZXdzt/9xHRTrpSTDgqzTd1Nbq0SUp4JFZFBH
MbF8Sxmqi30Kni1agIflR8OZ/BHaogM6X0abY4qCbj9//ipLxjN9UNO2Bv+RY72B
0Qgo1QTKeN56KzlUJygbehTFvV7FZ+FCTm/cWkLjeHBlb8jLvxPmyiDOAXHxqOR1
CLrRckbP16hl28dHpzK5hhQXpkD/zn2IqoNHv9ML48SxHmgkleS8EVoEXBVmtnbD
r5MlNACHU0cRjABhBAYhNsO57s4SO8Cwf2sFt8SwfQWlBA4Ydq/c9zUrazCg4yea
AY2Ql9zugqwp9Y+CaRJlAROXZbBnVHvmykKnVaVzmYastY7Tiu3WduYU5ZjqISHs
HlZ2KPT5+Ut9CjRtgJRM8Gcj009T8rdpXJFCUAgDRtuVRV0yLiKDnMAltrd7c1Wl
8Wykfwg+1IAEj2IGtGbenVzYzDFHtDWtlHCXTdBE8rONofAOFvuoBorj4NU+qOEC
luVW6dF9/7hunbLDeUfCB7iQB0zXRKGS92h6ZZuCYCfTL3hZlskYNQ6iybSvNuqF
iYmanJfmMXZuAJdbtl5iQPmFVZUd/v44hYX4EY+PbAUOAPXAivznTwErDP2hsF8g
B4/C0ncFJQ12Ouaxdap4Y8sgGlCJfxLzusBpaKJJUttS1cSS/9NF8Risu/cus+Bz
jrc+XsiNKcqxj1niXdq4rXzNvekJOxDIdefHv9PJBa2crZmkIcSqouy7HeDlIacm
Aaq1eoIu1QkX1fRYlEp9S6LdgVAz001Dm3PDijsuhKChZSjEaoISUBfqrySYQ6mH
kyZFDdFOlK+ELHRUxOTMizgghW+1Nr/TSeq5+VgYegpmWGc6tQ+cDogwYbQ1VL4b
wzuh0ngoSBEfz7uZvXQjm4oeV4FnBO08sec9/eUBXQajPJU+hm/Nt+5XhbTkT1LA
UxaHrHaVccdxA0nIrCLxaEURVKq7BlgdHPY1J0yg8i2wfevnEj6I4VRIp53TnqLy
G23PtvbrlpfjjxgwSZc3t8DycxSQJrGehIDK+m2XhtGLKxa6aGEmNwsTA6cL0WQz
Kc9Zx3abpnNxlzgwhWPGcHfA1UqwsE8hU3NtcXBN+aJqS17opTloWIrfB1/Db33h
PCQ3EsoYRVfn6C6fxRpp4kKmKaFgmcRb7NKh3o4zlWiWKgXw4r4G3XzwrFpxPMqC
b5nm+9ESYvLQMpkoRUuw1HY8eitcUvyxgSChaCicHu37Po7Ir6l+wIzZy4r7P7NP
VOhnJ6i+YNre4oZ0lAMpU6r0kD+WJmVhAWgTBM5+VbV2yo0tf5Y9zITVj9tKbnDN
YVNRH/H1hao+e8MiPb81JgePlPkU+OTb6YrFpdMHRbfGQfVPNTZQbGjKjxf2G2ws
MoXP+4Bs+zCUDQ0Z8U/F+7dSNODW2C0oBUyw4ppLCJZW5Li0R64B3d0i+MkARWrk
hbNCgtswblmETa3GxdcsMll/WyNTmkodc3p4ZQ2SQBXAI6V+6jQVNYZQHBE8/a9R
KJlSRHJtNA4Db0/9iql8StJXH7qiEEfuuWZWhRffZ4QjrAVQDxYBJrlEZuzfafh9
ozlecWPELbTTM10VjAKS74RqyvS26rEPRnTZXEB5t0EkO8JtgoMC6iy2VCTDiRBs
THKJC8NeUV1NeVv7KGBE+/WEGjsi4ud+NEjKd1X9ExIWyZYu7vL4hBCOCmYQYQY2
k9XReVKrQSm0MsDjR+pLeKA+wewUbEDlLx5fnN+dohi3dlCnCG+LeG5EZ+IylOji
z2/ZdtphWKWSNx8oMD5HdDneuM4EPu/nHq2H2ffzYy8NxSIFbsKKfhmy0VLWsfJb
7xefAFVQZZ5TNktSZWoVoxPI6u4slu/6IwvSuralgqx1gRWzkFtVdjMXEgSSyqZi
P7XLssG64LTAYOVn9F7Oeiwn6kr8sAZM9nepv+57Y2jrJpqfuEZNQrsEkyMcDStZ
X0u6vuw/L+bASLOP9DYuonxXGLrFImdKBRDSXLRBs82djWAvcTey4X7mGWAPa8//
NqsQhfTyamg98C0t8QBDUat6PMe8XSk+LLbYfwkrkj2fWxtJFeQLxIesgUIcsfbm
2pYFbfkS9p55ev7uFP4w9QefW7FXdoUKzh+y5FcBOU+N+arl6XsJdakQ1FJE97rU
Jf+xWeesuNlzSrYe3zAOwjhgChjc3g1MK0kkSSa3qoZMOmqtm8S4REbqAMBZwcsY
1YY+8ru5xsrvKavlVgIBUWr8Wdp3fCdqz/RUwhJnmEF4wsP/+CEJO6C0MnjmGmpb
LGE0FeqyFLcnf+fycuCm+rbnR2Z1XCvuXIVshFPlIpNHrITopxCXEo6JpjUxzgSz
/V/3EGIZtMdSfS91q7VoD2qkp+jZrtLJmI8VVuduCx2qJzxEs/2j65TA/3zfl31H
tBm+YOuTE5fMLds7KntlBWDLMgCbetW51CUzUD6hmmprVuEqZot3ItQ3EQpyqYys
ofc/UDV+tsXCQV4tdM976izszrlKn8Q2uIjziXm/a06g15p4+ceFpaPxDinVa2g8
sr4AtUHIRJA12hOveHA2T7OmQ4IBbweBZdfR6jmL7cGC0jzOYGCi+nimmB9TolDx
VFBK12CN5RI6H+brtZGS2QkY4BT3YqsQy2qa76ek3NN2tKvWF/SXX/ClUwbkloRZ
MMUOMTknk9uqD4itNBNlXAdajWzOvUR0rXaItkmZ1IK2ba2z3h+9nnex0Vieq/WW
Q0thij9XrRQ+qo2EvZxY126S6YYmyokAWguk1b/18YL8xP9zueYx8wb9byZKOpfW
T+0NC6ZK27rMyougFOy5OONCI5VyFh0SEhoB6wYPDJgz04aGkSozJ8qIfPpbVscZ
Db69t7LYh1Wp0Oelevu2VlImMXMb+Wam4o6iJdqiWekx6nQgGbN8mKN62B4i/WL1
teBEgaNStEETPQAjtY81uGVdor4s1W32vC34ehE/Ef9jFbSfGdPvE0jwNmiVDXXS
TsMKxcDbLurG875l+JlJYpGs2soIaIp089DEPUul8+YpMjWxkL85BB66NRKu8hX2
3VjWJoSQWjNj7rD/kQc57L+nHJaUcB7jxU8BF1ZS707ryDonI3dr2DFEN8j4I/kd
APyxHeZNrWy7IBXVex3WonI8WVVyB15UAqX7sCqLVaN9FfwI/jeCYLmxQLr9Lj3U
QNYK8MGaXgMs9xy8Zp+HIuf9koXUA17LStoy2nmR/musgHHU3ky0NL7vMblEuqEx
tJIoZ222WSZRm9kjYjys7vDgBaNR5yDG0HTBN/QrAsPXxwZIcaEo//hnilC54K88
9wDKzj7Eb97LS8oWXoD0iCP+2nduVi/mLNnnkY6VPNVs6bzvLHuXANme3ZEc3Aca
HzY6P+my9AMX/ScMPufxTA4yOaDah8QkZDsiwKO+nxlBNL+1lrRFGh4/WE6astS5
DeaYjB/gUKkcQJnu+q1qLt6so1Ep7uPBc64lbrtZ//OMTkMjnp38PXtXuRzwf8xe
gTY2HX6r7VxOdpI8e9oq+6vJqEmZfyvNNe3+NcUfIEoalIL0rGT0R579NirLizPJ
riWqyEs0AqwW6In7UbnHOqQcyF2Y6OsNzoEzoC8SG+sFiG3nxH+d/us5yaafRT2v
F7TEEzgrqSSW98illo0b1VuVMyXTLN3LmrZSb0YxSU6Exa5zbVUL/Im3eEJNlAHP
y9DXgGMFDS46eA2gaRqIX+fo4cLostRJFAXYhB3Lp8ZZgITWEIV1KpcbhwnunF3o
nZIA05iby7LZZjCqswAMZ3iQoqR6mTa7XCm0JoPd0JaPFigixCgNN/fHP6Zy4gV1
kifwWf1sCq1cgAC3XjrZaa4nOaBYefERezTzaGmasx9s6OjZ1CHE6WTFrpBaz5BO
LKRLKD0KDQMvbqsFFexJfG0F6Vtd7WaABQAT7y8PtonlkM+cQ7jPbenx+l9cBAva
ypkU6Kq+iZhwzmhZXb+SPdOq4GbF3Y1Y+VjVkpOBo9D98OEL72iOl7/E4Fx9a7eP
8XfPBO45FRYzz7f6605tjDr1lktaAKeL7GmsFUzPKfZ/DGY1iRcQ5Xcxpc/R9pzW
8k0Eaq/1UOYShjAOEf2FJyMr7RMxtRrdQuPQiRYhEWBChInd44mgMz2l0J4/poNP
O/8BX33ctWVm7p659jBz/ya662OxkqwvuYovyenQB94f45OTTM10UHqcWIfwUSNe
ewHJkKgm/MYww8sJQ/8giJqCJtYAlxDkWvE27NMT+BklXPZ5M6Grjzk00dsBqGFP
KiKqC3UqZ9PtqlWgc3VGxkh9iISSqiwiwXvE4Wu1JtIKUCVpVANWohXt+rmVjg4r
6ikXsx68PIfZ/2llzAysyPdHS2TI9II9MG5g7lCfp9djuzjodJz9RZWJc5k+Ij0G
viu4A6lkhDjbKU9M2f9XxSNmKsfFEkYFtDzWgmw9y9GTWysOhstyEeCfQvWDYaWd
QOVftO+4v4AbplvgEXTTB/IPVD/fR/xJmrotLeWkMDcQvtH0fimvvGP3pT8v8VhM
IJvzCRcts96llQBaBbLeNUnCcZSFc3TSf70eqVGyH2PrAJUSVuGacKSogUZ2kMYC
tJKQRkEbRmye/BwmSaIkSh7z8iv/sKm2IU2SicU8w4tuiG+Nd+zk9ro0+xCgEIZS
WbKlUicaVYDxXiavlEpc63Uq8kpXv13R9bgWpKhaaw1ZsLtURkwxmId7VYuKanPO
y2lW84ATC9ZOZaFhZ3p8aratXrdEvsWayPpmw/bk8gTC45XgtnqqTpmscySMtPLL
Q5rukjv21BNwv1aYyan8BqflkVP03vNiyjjCBAvYdnQfixtMN86EZCzs1MSItCq6
fQMTcoz+IWqMOezBLY7zlrhr/63eZvjHZbdkVBF7qJOwp7paB9FcLzDecTKAi/Hm
GAsmBIJVLx5pMbaeqPbcrxn9+j/eLl/apL8OvI4z4HJptqT0oni0/UJPfdhl4yIY
0UypAMJ5W8qBjvtLJCk97hojIeADQSQ9TExX9+Ozkjw2brEiRgVfv+ozWZpqzlOF
MGsTghrCCmU4sMK9sw1FEqZenUCOZX+uYLfCa3sQ789/2oCGJDVA1oGuLqpNX8AY
jNqfAxCthvxeOv9UGN/4aLWmliQfULe+kL6yy0k89MLPZBh4VM9vEIHQw/exmama
LPDcoyppR1X50ai8ZzwSm7LewZyBPilFKxwacBNDzlYarwezJ3Jr2+Yhl1c/Krvg
iefoWZtftMRXGd8P84zzIKuJ3YC7O8D152rKWJUjy1SIPlZ3dS/fCrjCWAzkpSDK
zEsj1LIPCr2Uz/oB13w6RnGm0/4kQpg/aMkU4HBIkzoupC/Xof9+D/XBiSAA6VLj
NSCgKXsfZqeJz2FiGGzQ7tE3kxwRAuVx4nQMr1ccqwB84uZvIKQa7QTOvz4X/O+H
F/XhQ5Hj1lvPSZa0czYcEGhevRYTENw5Ov5A6kZB4TmG3b2gHrHzR4ohN4mrN6WZ
Y2XQQRTYHlShDrgDGqLuZeiIttPeb9blkR7cnKBPH/XxlpUvAXt/8vhvAOJwFCOE
OWFY0oe6M2LxkLjBBcn5fwg6Unr9TNnxRyAs+fVpN6lcx63D3+ZIXaVwEzKxZPg3
rSGOOUCqcW/+xEUZiP47jQdsHCOR6mSwFR1e53qgsKLfAmgv3zSfEjiDrMldjTBU
2YS3sfHXKp8noEkHO9C1Y9+0xzD0DoXtBNdl562328hTAFR93rVfKxb0/w1LQI9T
nBF6sZwTda7tuVazZoXYoUy9UQj+69V2f2aRCGohtpDUdnLVgYMP9muyojJZ2piB
Xmrpt4RXq2fqnPT/6KrYd29lfirfBv2wdTSzK3vppU8cgZksPHv2CcZLDdjzL0O2
IH7wy9gUUejcMSJEHnfeVslvETFvuBXYLMyaQf0TLSg4qCbTFrWuFPZ2QuXOo37n
Uqgtu7VE00YlXUT+RXXndvtYDqrSwSOAs+6t7SNdpJ6qHcve1HXnuEurm5NOkkMc
MnWXK9x9jXfyRhcduZMXh0IAv+zAC1eczLkdjgxarWwYO2N4ShARMpvphTGFhv8v
dd0X3k6zc4k/+wCR+iT6DjDJftDnZCDtr20FSePmUsJQN8LMy7G+v/YY35MGyVgg
gmBKakPUOVKhMNDo4v6W2LLmq6yAHZ6xTmgc8/tA0cIf+q/m04/LJkGkhFC8Loqa
Y3zRzyGc+dBaMzkqtKoU80F233Z8jk5LZm1LuhDHEuiQ4GRB99UEtpasYULmMjXx
zI5qJH4F+1q4VOLMX8rxEWNh0zTsJfeROk+Xj7HZHdxa5EYriJ9XlPyBkWtQrpNC
lBhzIq0DkvhPfQrQbF6iPPzs7xd69G6LRIhv6Z261kAP/DLuUYFsv0zU0aycyLbV
hQHhvHAcodTAiBPyHAvE3/biymPSjCUPfVkVbE2WepohTNOIMhjOiE07e323Ur8W
BmMRweSnGEfhjpYg4gqBIFuPV0mm3D+9ttGNVvRJFiGEZExNoAi7qghB1GoLdpe7
PlPghzK4rp8zU4PTzCFklTZQj8UuZXWisJHPBdirljjy0I8pWwea6mB+x5hhOw+H
QcogXHGkrJLQXRtSy00XGoe5XCuitRV/hXS57sUc5bvVA4WypNCHpLZqCgObAJ11
0RMWJWvgnxq1r9Hrk+d2qMmj/zmAJxLQHeMDssgI1oB+vd2OAbxdk7hXO9+0a5O5
7vXYjJ6v06SC4b/SPZlmggwi7a8SGKiRgLdB2G4dsoEGPNZN1nAHQ/0KJ9NKboqA
y5WQQVDQi43Q4Lju+tsXVXDkG8D/Sw93wdUPt6e4Q0hRcuEgnPVpLPk0NMqWJnxI
N7OQGQ036VXxibUFLOLzrrkqBbbWOwgdrWP8BcZenwzZMI0PklXiDoBEr7kRIi1k
NABIFHkiW8veEKiU1/NGyLi9jkgIg5wbk5eSgsZ3wHFcbPjfdP2KzoZViS5zrpka
6OAgT5n4F43c/Ycc2EEwK3ScGGLvHmEIKNnt3PBjEWq2Aq+QDcEN9w5ctQVPwiJB
Fjys/iGN+aryMRCEG0eJ/zkVTh5Denqk4dsqZ1FaZZcUvqJnjAVimeOn/K8POe74
IVKfBmWAoMfQmJc/H9OyZGRgxfGHp6IXn5kbH4SVQjU/6vZLoFVlYlnGAZ4E/dWN
8dqKrIgc953gNnOr1CNJ+xnAQgX9isUFw1K9LqpQCFSOjzTNYbFAWpJV5q7VImG8
1jJPUyN/UbJM2Rp/aTS9mugKFUqUeYrBI3CR/KzpSLzObMjY7WaOqWY7eeM8RuGR
NOmbLN04QcuUWorE4wls9Ovrf7Yzl8y+C+TJH25bdqEwV6qzVNWy14yVgryWtdte
l2sz1RhhST4k1Pv2pT0A3OtjDrLuUSwYixENZwmXZxD52J0TqQIk7ofqRDubxOxT
V9cvcXUGRuLGkJbI5PgdYoLnCgTCSZOo7Ycj5xd3o34e7bOHm13tdk8KUPewBnsA
PQ7/aM2ZCM8OsIwZmLtcfKqV1XSNHhT8utybFbDdj4/Ob0sR6w6YYCSz63W9y5Ww
zXKYW/vgo5bYw6srl8p6un0l+Ti8VYV/HEjdkM6x1n/6ZCbfq/xcCnPLJKwYf3dA
9T5it2nobPqvaDqTmjlOseGoSBQjCIyU/LcXy9hn8UrzecFRxi5q1Uvlp64byY2Y
87WqIxnuLF+sIsvyvkVDtLbJwivgSh+w9UK9v2lI1c0HLLQFUspya1isIWP2K8Cj
6SECt9IBQLKHmmkcOJTeNMCcMjpsbKi+8fFZwtWDMBHlwASoNx55zXctOhy++2q7
Eg29rP1GcH4jjn4ltAlCnivRmk/hXq8DolSeC3grogeCqJA7TpIywc9XrmOzPbzA
qTXV2flSsaetZvWsGxON6otqCMkpNJG03mc3fyVM1DV3Gr1y613NbqVLydotczyz
2HGmMUzRWfJQFoHw7IAVASQJPbIYlW3ZfEwgX8oxYW/QTsLRFmEejKYs3NGBqAkc
ecvi8n7BKKyoEO0fx/UGxLjZn77UbLysxsCw+tq1KTTBWCzB9xTTn9uucpSg0I4t
sYZRvQ7GkqPW4InGgBSYIAY7/+uEJIW64lSdj/siAihkh7Ljft2RPv7L5JfR9hG5
80310oxswNW1zJpH/63aK2jwcj9USNPgQVSTawGtYaIWdLBvRSjS3/UOSu10dg99
BCyNpuiY6WJuQoRouCOUiuG6evq4I61HH25SHa0hFEAgr+TspCFkRNl559EklS3h
xtA7KgmwAwaazCJIQEWAf+3yfwAbrJ/Piv18dlv/V5Uxz3cYUXsKVC72lS1dFSPo
wXeQ5Uu2piaOW/cx+Z/ooRtz5TSwApwLArnlxZTkvYaN/Q73fcOEmS0UVCtGNZNu
PupEox2xLF5OQORUMyUI6wXgCGDFxCZotf2++UsHkyHcMWHRCjPtVRv+/toO4muo
HfN4/q5PNW2dH4psq/RASFKTur0REsa6aMdHOFFu7RtaCWh6zyNEVn5cE9x/w3Os
uJ/2U+MT6+tVBK4bpnU47i75q8w2IBuDtdONkVQ6JHLlN5ayM29mNUJmTkEeOKih
Y8WWG4K4Uy+jmNhqiL3DCU20069sLUZeSpX2tf634Sao1IUntU4wyCPSXRyCFMmV
p2tgamOBDBYV8uoDxXY4r5W2p286Tc0wHeyNvJmIFXTgUO2QkhV2uugbSeMtksef
N0qhWoqE2Y5QfsDLexKflELXdT2I4oi2l7hxrqAI5oKwmzqAPkI1Tp6DPrbLOD+0
OnrXfuZiOb8J5i1hFn69l8HpD2ENTmOpQDU3Nr7/HuRfWkiVWWYTdgKR7AdLmP/n
7rjLV77QlZodkoAEc/KFe1yp8y4BOJO/21RTF8/+ta/XIuWyGV886ACZWZjVJ5lS
+sR+30gPHQ9K6a/mfQN01xFEcWr9WSdMO4UpGEiGsga7BlpH3LK2d9ZBDiGGuwSK
Id6xzTTy0mzYNO6M8eIVYkxG1UQt0wQ1Wa4lJ8mJBb50La0/Dsf9HFwMGQu68P+h
fXBnEqde+SJcJMyFtrbEWQ2rimZBdDTyM858MvpamUnKysd6uOKS/puOTT0bKECp
vCGDxj6C6Iamm18fzr++iqJJFe9kgsouugVdlrYBB92/lpMTcnyCwMZLpfIvbOxI
h2RcTwuOWurMCuPgJ/JpNCJ/ossPAopJ/pnPsgLXlBvFSTslJBIsbP9m8RiDjcKk
Xz0riuff1vmE/RtCW0J9/52/9dk4IOZ7U8EbR99cm8ofTq22S9Fm/xqtbFWiwTup
dccm8f1aKPZ/fR3qKdjcKVAsC+PfySfLm5aZXvjvhU6GittNYePpil56/HhGFHU1
qbLAdKmg0knh+I5VKA9x5iHcgToM5f99ofa/1Cb9tDg2KJuJyLD6zemiyhyRVtVR
dfra2KNLvn8cwqIQfw2Q4GJl4gDhwSCTMBlo9q6GuqbhN1l0lkaULkMP7lwWyCx2
nbaQ947OkcqiAX15Vp//bkGNc/bnAg6BM53X+KPJhAhjsAY4bK7a8LEW9AKsx8Me
8kVbjnx3u4I+fJLATPkdDtxoMk4qi20wE9fXYtuCUBu6TZZD5R9oTf7vtyx2knYh
5vN1SEWPtUqQ8pEn/04qFyTnvQpWhvZFk5qJaxrXzZFsfnla7zpltY3q3E34yQND
FXRtBqJIAeYNlU6lTwJ4/rTPd170jEJjxmaQaLNvyem6f0VTPTigDyTT17/iMlbf
/yjUxM3qHP02/1sbL03k66Fx3HwgKmgzWsiNoshvw1p2iQAJyMF0PUR/E1oXiwjD
wKaHBZY6QbFHYuEiaUxRo9OjJE/ORUWTlbEZn628LSGdyMAi4gQ4FI0algnAYCQo
K9K3ehYexBbckZxDjmKLKSqqHqBf3++ohvePAsKiJYeBdYLdFRCkUfdEy1iARLBT
Y1K0vhY82yHbRofp6u0PHIkL43VRti7B00pggKY3FsDQvOTydVUbgh5stkLbJ94R
B8cf/xxc4qL/eJvSt6NZyhr5/nO7LPQ9YTTQNNy2evww3nBFcEbEh5X28ygfkXBG
yi89tVldGGgFgAkYSB0l1HuOazVleUlRKHFZo+ePmWw/IeFRiS6kqzIN3V3RgVPe
7FEhNcivbsIt7O1i0zTttF2Nf07/xcZ+HIF9/Y+7tau3ahZy9TKfMj34nQKWhN4F
BcKS5kI5NMalw9QZZlzzvKlc/V8zh1ZjEIndhhBLZEXuTPAzDiQYWo2he3It5aeA
UZmGdfWfRc767nsQ2uY/3qHGy3fe40APtjXtYgnxwjjTCQy0ASZdN/yFEz40SI5D

--pragma protect end_data_block
--pragma protect digest_block
zarFnb7Jez0Ok2Q9pYhWl2lo++k=
--pragma protect end_digest_block
--pragma protect end_protected
