-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
jUvgoLPLnJ64qbm5uds4mYjtebHMYXRzjen96NS5FZ1Bashh/UJtB+k865PSwEww
tbbmt6OPqtq3NHGjQokGmbsMMfHEA60HAmF8RWERn0KNC4MqRWXHFf8z1RrNaVwc
leYXYxe4+9kKo+/3P2zoi2avQZBEoC81SyOlR9oI16w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9664)
`protect data_block
nsnLYBU367dxnmmO8onCajfNQnmDhexOwBQS22WQGHz7qEHoTTxqhDZ9r4uGztz0
1xRMrLdUjcJhWAs60g4w702nvTfCGhv8yIHaCVTGkxvJqNGIgcyBkVBjH8L/9QjR
c1LypfM3Dw0M8kHJZz25l4kU3Fox1b/n+mO4MOjWYHqoo5CfR6y2JTqiRBzzLRQR
/bJWyLxP2lrPB3HUba4Yot2jfjs+wOC2vkHLyeKkKyxXl4fMmaTmcwqSsTy0xWKH
Z4FtA/cuRLnyE6xUaTFY/uwDZRUoS+lSpiCDt28XtVtEDhBcKLQuEt4Z1NixqJXW
n2GhLSkaZbh9+oGjtMp0XhncoolJNfO8/pU6OhkJBETX9jQeRh9f2yU0b/5cr8vJ
PrM68/dtALUI3VT+UIXwGwwebgJec8k+DTYL2qCJabF5sXlRhTxv4yLna6ZphovQ
dB61Guu9NTm78LdFfb+MS8wueBDxVSwlMHPEHzjp7QyHFQq7p+oRkB4aCaXLJy++
yUSGlpxURQ032vD+J4uxW8Xyr+5PpuqY5P5kETAqSbyT5Pf/CJDKTZH3+F6MHlEn
edJZAXXFiDRXk9j0NqbeMuB7XuWOIwJwUmOp/NLw95MUOL84HGlpuXduP3M5qSHP
BSDgU9h/rX4GXdLu92gK/xyTpWgo28zV9Wp5JMhMyTgh2TASH2CsojYfGqkMVKUb
k+ZSsOIPcoeF5qkjHAk20ic3fcJdiJOpI7yYpTbefakb7xR0ZgafYEdcQ94xb7fU
GcQQPa/L1Zu26igK6cazvy+f4VHRbD/MSOm/wHF6DTHW0EwcgG1zwHUCGsqjdkok
9/REus3/dq0SYoQwsDW07NtcyyThG9lJnuX0ZGJs6EBbX+6EROh/Yi1iOTOQh+eU
buqnDpwlMje5YVhhMVBLHLWLeBkH9DzI0T49oeejpcuBnGZ4Osx25so3AMPkhBs6
xofWVSVgbCnz7LUA3W5rFe2vvEwnfnHoONLY8iIJh+WP7hBvF21u2v+Q7ey0zoMS
Kf/GLVV9egV1p1UqajQ5rGh4gt7+DSLy8VdIyk9kDFW50qps9t4s/RaeMUGZH1Mf
6n/FS3Ff/V36rGfhR6fqsR3SGz9Mi8/AvlkoIj2Rcme88O4st/9YoQC72qbNPOT6
q/ojQw1XcKraUc3a323vxZns3CsYhmFOo9XxWiciizuXLgkGbGbWTXfMSwSyTh4n
XhQ2n/w6ZNk7pYkZiZhbfuS+Dk9QBVr6SKAF99Xi/iCcjBtMBi+/BREm5eTs49fU
8QAhFWjul4skFpca19j+HeMVqmWXzQ+Nz4emfdk8nMWRIVIctrHwfBvbIRVjFMPg
0yYiO6pHiP33tKNXz/xqK6ZnLYNuqF3TT2akZh8rKcj7Io9EgO9MCnoqkHp03VS4
YC9Rd0Ww7IpGbPMio6O5GToywCrHYLyt1P7okB995fy1A/TWLCGQj1LYk7xBMF77
nSAuP+dEitUeDgeTF9SktoOSOYsNqKuTZc4mM2f7tF0pln7GZddM+ctEjTVDJfZg
o8K7YrHZBV6aljU68LT1YO2N5SDU8uS6v06PwM3BQBeySxDEWhxypmDAs/XC7HNv
fAEWEX9GINJgGAMGAydvVgVSWjmJVIh3zdx6h+nVfrjfzNuMBexJF6e2DWj6iLC7
shh2fwKumlGpHDrCcUhu5BhvIOFTZGShPER9ssoAlERPzFwvaqB7YaYz1fl4eZ3N
verHjanOFn272nqta4ZDC1DoibqSTGvUn6dC4DyT76Bq5QYivp1r5E68vnXqGf5L
9YroBYxwbZqvfqhoxb1XN9QckE9B8TAvCJjKxX7/+JMu+5r0UallJfeP7TQpxPUx
oM1uAXhVRn8qOinZ8c5O6GS/xuPgFboHKetjzxY5cHTrYeTrR+b7PuoBr0UY0mQ+
9XZoj9t2vIs0LW7IkaM8mVkVb7j9+fa+eRDQG24Jv98EjuU4fU9fBpStAl6ts4sL
C++ZckUV0q+gBk10FhQvscJmmit/CmJY4JRkc2KKfLwzbeFvx2s9hETT3cEvdPWS
DHEqXQgpbkA2Va+62k1/k+rIt2lnXMOgxdMzMKsK1WdAywsvVzqEw479MECOs+Ck
/g+WN4NO84g4VncQqV3I7SBIuHVSkm0ejA9odKNK3yadY8QApUMBBOK41lP2mn+g
yy9zW3vaIRCbe0pt7Gb1Vg5WJFZDrdwxzQpWGuiJLdRiU8cl2d/98QQL2qQSv49H
Le6X4hw5u3GXfbAu/+mzLS0KBibx1QcGeEzHB7POwZh9uUsjDm/oO3mIMggS7co3
GgM5s4xYq/r0rY4HcpisK41+nIZePwZH5zzy057FdkxNlEIQtDyPOqfWp6FaStcp
uuwjq7KLTO+x9RkDdrDUyNBFuBYpNFoMNQpldS7UXJ4ZwfU/PcNA4RdoCQOFzuxO
y8wLQYgL9e4E/59Dg63rnUrMNQUKudUmtlp5j67OzCGeIgI+QwzgnlCi3UNncBcL
7Hjv3ZB8mhhXBQrv50AUhIb+px+7ApnfsBxWkQ89ySI5bsPnBLfIBtUDfDjtBoeP
c+B9FQyxBAm6jeiZhq4xRCowa5DHfvmZYusxQQpGe0oKigomMHHHT8IXstA+raZL
xWFjgMqq6hQykj0Evvf0xinhOSQLWjnlSzj7xaPqVGu/tVxI7bURq1jz5CJIIpHB
XUuhy95S7r7T3PiI3Z8BXrGMvQjNv7Vo47C9yvH1AnUFsNlyV0PorOusqmf2fLpB
x4FriqzrqncmUcmRQtDG7pys6DbG+W3x/TVOe/aYb8fCs/whoKHxG3310wMdcE6L
Bw86Cwmsup7wliTa704HZe+YxYUszsyf1fRbVa4LLG9KQ6LqLhc/2FFScIKQsILe
WAUbcFOj1j0OSc09Q7nt0Yh2aY9okzIbXXrfomS9ftCKiFFXWe+GkyXgXqfT7/1K
agKxak8ES3WpKXfk0AzF+yAIFntJ8iWPmotGQtzXlk61aGiYUoRHgMLGi+xLrKTZ
8Xg6c+ypSG2+6aHCQKe6UMl2pvZPHDffly162LAb6LeBhpQL0c7U569mTNDDG0F3
2It0DHnDMF28o9mZlcG6FeaEBTiW/G450yk8Nu+Qlnqrorld/yRqPLICa5zkjxGo
E4g8gRXz+Yc01C6LPALbcTjRXC4eugLmzxPumAjMvDdCY37YtNM0/CDY4FfzA4Tf
wKKV7a+q4jUu19DI1Ux4vo7ZlaPhpC6a50TMu/8IQyZ8w45lRouzuNGZGPw20t72
D0TNysVoo2XkAB26LFu3DgMeJ+rEIvWj1jmEcEPs99h1cVMi6eMnQq+5o2Dgr6+F
+ApF7ilYkLYye0W3Xrpk3dr0Chz3EQbUqz6ZFRWUK60nVMEyf3vEMV94i3rA9KJL
DDMLsXHF7h3QXe/DzK+LHYxBZuxFX2AuwPXRut6Tpc3Q2kopWr29Ptrhz+dUp+hS
eqU+ucFdiufcmtxkaewsA3OgNApP0ZMLbVsDZH2/Q6qqqdtHWplyN8NN9iJhmfLy
XFo+h6I6mJU3US09NyCwIhBmA+JAlyPRj/kCx6dIrLnVz/edXnB67ZupHeq10w1c
DgWwU1Xlo58mtDpvDYYCWLHF1cX62IR6Y0Rh2Vg+M0FtoTkH1zuGDlBjAchZfiaz
LPJ1Fz4IVABBpLuuWM2gZKOEFbpmPXXdfG+Xr/p9N8u1rGHhapLhFOSS04wIu2Ui
yZWdYu16l99hBdS0ygVN+m3EG6QHMafLdvXShF0BTHUcsqkTqPQKZGXh4DfpWrmG
s/ZyI4V1LLMhEPAPey5jcd+MyWGcPp/e1aaemsnDCBtmy350I+POL7kxEJYqrgJc
eGx9pwqbzfEzVzjAkWMm/gnL9p2ENKpbEAXSd+MQQWoSD3v4Nsx2mr+W8yJhWJH0
oSBTAGvWhS2bT7SpS5enUWiRTaIP/dBKbQ8D0laisK7Z0eEZiQM+gSILVSD0GzUj
9GhNXB99FIIk1G37UwYICBRfbbSiuZdeoh0NojqFQ65ZQ8c+fWAoZCB2qk8EY7wA
gNbHb3nTPYFzAkNeB9bLGNftAm2BQmcjuvyxYv8K6MzC1yq3gms/mr4D2DylWEvr
krIlmEhTix92AU/U5xRZCcIxrDK+bF0u2GYSBCHBikmwloeP0oylRjw2nBzagIdg
uOSpCIc5sqbcnsKC2K4u8sTSn8xYghDUzNpRmo+sgRj7EqIxrrLFAsOMZsIqoYZm
HI9ak41evb2nG2qIjY73rsCWAzSf1TpAXDFHn6Mo2WNOFObNC2sAHzgmWrYjQmra
n2DxL3mGlOnxC1lCs9DggOyhjeMk4TbfYvCidE5tGdpmKJxDcumGpGNUbjR6PcX4
/9tD9ITweCJVlfH8p+0GGBytcAz/vrLnuelF7OZ6dKWMckpYYvZBeJTZzxSzsL6p
whz0F+0konXmO5t2kwCAkIMsTNBDbquVqRbPcHCf4xgTxNWpU7+SFL5kRS08QnBV
VAEWhUG+rJ25lBTspnGJSuchsHjFKs2oboP/SpWVbvTPZmT70JfuamcO47MSknor
27D4dtmzz9I92uJlnpTGH8EsloXMAtnfFOCWv1unB3RzjhAr0xo/1Z7Kf7IXitOG
ig8FX1c/GVDVpb1G5BRAdk/3JBXDNU1PXZbFBpcuYCJXoIZdb9NdO4waPwWzmbHQ
/y6xWXziWfCHnSOLUVb4Y4SZcRRykXsyE8SUiN3/Ly3skd27ZhSPD0B/8pGyWdDW
i8nr7jIeVp0xRk9AJJf/yL85CGfYjIx6CVGACxh1MPMPzcRGqmG4lzlXJOaMYSin
PxVhfk4+Bss0sjdMRdV1Cq8zdGzo8DD4sZ6sZMk9JM0JX1V2n3LUSD3djEW24EDM
9fnvNHDqLXWowMhlojrpaiPiy3YQOXceK8mdNyyXS2dlNYsYpmJ+nP1wv20BfN1d
SwxEMd6qxKdth68PglFMIC8fQRSYuFPFfmavoyzhCnOzut0lRYRBiXWabrN1O/nq
iR5OT0z48rKGrMh9j9DUGy6xpNcJIYrwQOJoEazAKwKOgWHeq21aC5XSeqkb/AJn
9/E1XKvvADyy4QMZ+QQNhnubd8vosM7wAvWZJJPfh+JfQrs7C3CoxPcFtK+FpJB6
Ye8pm/LVE+dNl6RFdqiuyVGTWvjndmbbrd1TNTb4BXAKGi0ZdQoZYPVpCoEgoHDg
p8hKe5jgJP48aoa4zyh1jC2LnzwLV+KWrc1CPdYc3IetMpvXObo/dBRUwLyjJf+m
o6LzyzVrcHO1URctMHA9Dk+8ZEBgXCZDDnzMxFAuPUC4TXV08yZpGNTfQglZCoxd
IzJOdwrsZKgvMqteTMhRF/SgBYndBYJoPAvZkd5u4x4rIeM6W//W3/PxCPKAjtgX
Een+TDJxS9Tcd4rtCnyfrIjQ+zRdHVO4X7WkD6Z78LONYTZUuUQVLt5UVDoSsWdv
R2YpdEy4Gl69kNFv7Qevnv3LqEPEXN1GCInqcyUiLqaUQ/B3QgJdbSIAgvAB4cZW
0uZisbfbs9izYA3pxuhvcFDXvBGuQVvgGZEbP4TAqNVidtv2j2g6Qou+BMOS4gGJ
4kbIb3yi3gHNGv5KjH4mFvlGEgOgy7MwxFeiDkNPA/bFJ/+epciuVspJEpCb/IdX
MD8kbiFVjp+bfplCYIrYMbHbE8bjufPh7iKg4777vVQHlaAqBB0Mh5jhl4l+R6L+
/BWdtQrzt1W82EyQVrzugi7kXFG4AwcqEvqo3jEBz5lyi+YuwfzkDtY2cq6ehMUp
Nk4q4FGMiAdOd3mJpchuJiAP5XaSZsu7mxHF67Y09vAuAouEQ5gaVjufpoMLNcUS
55GbZxLsUBsNlLrriMpMyXAcwj+NQ2OMO9h47VbfOgVN1rtKWYmUSlORPIKlMsU1
c/tB89DMptLaphzdwO1R/QB7qqFw/k5T7hljHtcVtPQNfz9INy/ZFNPUYb6iLnSl
P2MWDFDHbhD78AW6aJwHp/LyqunBkDVLyk/7xoxJQLbYBhvW5nz3ZofMnW9d40wm
VPzWRIxhwmkYC+Ur1zhzVP3oONBLAboEh/Um1maSRZn8j0emMpoY01YfkSoZc8yH
g2gt3+DcRR5Sp2SJEgfkE5BXPp65o5aN2gMyN3gpZtkHDA8ZVN5JsPCtXl1vOoDX
kSNTZzZz4EVFJXWiR9Ho/sZ7gPPbuepMuU1kZAQSLm6hYip2Sa3snG2gbTRNj83G
c0/Rao10pJJr3Zea7xWyS+D60UJlxIvDbkd7lBgRfOfN2kZc5icmZozKu3wBODE7
W/hIyzAyYyQ4dqShcUN3xTa3lEtwPfPnMXsFMJkNt6r2mwoUrnfx0Zp3Xdq1EKX3
JXSD/j2y8wS8XfTJjRqc/qgjjeqiy7ui5OvcuHMaVgNTBr4es1V/i5TR/owSSYcH
T229rfBnyX5bRP9Vq9tpC1xMozqA+pJrPOPGkh3bPSqQZvrlvQKtCWr5ns7lzR1Q
jLM3uRtNZ4J68pMnENTxcwjx128aYnoi66FCLB5Mq3kGN4Li/4H2ltnPVxOHG3Yk
YZowGVSC7bpR0NaYGQ+DiKDUDoQHmW80qdwz5E/X/vqG7sIsaR21JpgAod0GT8IS
RG6QaYUQMjSezNzlM+eN3es8Q4dGMwYvC3eL/yNoDKB3L47t3A+CsXdqIToBJScf
8Xgj4bj4CmmXtIK7z4q9Tsiwe7R1nUW4t+dFpY3WGsO89VBNLbzcD+4h8XlOfa2Z
/a3J2FxohfZooMxrQrfeNrHuE3UmoYytBcUmbABg7SGJCs5q61r9Ry0UkkSoMZsz
LO6PBKe1j47ju6fusNLjRR3iG5VRsXspoTqCGvXvZpWQDOPvPIcG71n8P3sWLpdU
yNtFHa8bdtbP5aFRIDtyUx4yh2up9YvE1TEdM98e4jZpFP+8kMC9aCAQBpQn1DiQ
6aRSz1onffvXfTLcbAxEHSoRyFWmBY2wYv+OfQTT7KdW6PSKwHc56NM24s/yLFPS
0bHCctTcpcx1xiS+wGBAd2MRg05eYeFdONdahiD1fROgbQhWZ+pZsnQvm/ZX7jlK
ZBCX8xNTzYNcpsQcBwX9pjTJSU0SFmJ/AkpHktc1WErVvFtJTtgZvIMSOk9Awa95
KmcZunh5aQrLuQInjrJ0iSNe8vGnPZkpNWjGR+3ZAflQokSk0wnvxz2GvXGLe5NB
nCghEA8tmDY3UW6/2IG9LYJo1x/t69BRQSkfp3eLjiHoRVC97YF+O5XoGACo9PWx
DRnq3JjgpyjPzPP5F9+GdxoI6KZRdMd42GvkbNgxVsx6m9a6QUfIhEMZdYmNXhHQ
50AkIMrTR18Ub4oZYK/uwpG4PXWApoY3eXwZZiiYmLozmko/RX0IJAHzvoOkwIEg
3oIr35UquhYczBntHA1Seek/+N2ZmFwXKigcv51q2AICgfpmBt5Xnz4JRJopHDq5
62NLwqhjqU8PmYKX02AbjmJBrTcYzJrH6Ui4e2xHpCAsXrDZM8O+KsJTqCSV9blx
mT31rw2DXW0pENCycI0bcSvfqDNreUt6YPheIU9dArn1/2hN6cbODRuTRLFQ9dUC
f55CoWUIF2Tahf843v/YvPKSY0zkCpNtr7XcSvgjRQfwE4azhrfq0ysVHqJ84D7K
RbFCREfDyL+fQFdQQiI7XGj0WrdRjSKttbVBX4GQ6fpbqyZKvkLZxQLROgYEEvNW
o8TzrPfeur4aWOj1Jkl1sOeWSdyhz/oBdxDreFxt4vkP2ZN0tB8+2g7bM7dj499C
rLL67qvU5Z3kXLdKPN2F3DssiV5JDTFPL8riURsaNikj5QF0Dw4EE9/X6kOBiki4
PhT9mBSZpFwWXV6z5tO4R6iDYqILyWujG7WURlhqgUqW1vH/AccyDK3Y+g3Zd88C
7C+z+sd99AhHUUmXiN88aBTMtTOMaslYyQcg0w8lTb67StdIgVXu7Zcb624a4Z9D
RxfoxLvJTx5gsrZXNMnWxQydAUzmXDXuTrZeoJRl9JDR6fpSwFfB+lcNqZIEMs4i
ljc3n7pQuX0/Idzz/IAyYo+JxXu/0U6/PQ7EASV9TD6IwCJBiAuvRKVSXCo6TjeY
CbkzjcS9gQw31iuY6zAMGLnNGZGa1f28AafgwwvqhOuMKKjGlS+KAp2sZG7nQEF9
n8a0QZs4yvWbF2OGSgyQjXl0im7vp6QHlDVS0ubk2mNYsazj1ds9NuAu7y6zQEny
gQHFzAxdqpJi9rj6jx/0ljhpNUdKbPwu/OEg3b2zCUDceV4W+gyjE21O/jJyUC1i
sdxBOTadHz7jbOLhmcUEkqKRNQFfRU0pk1Ya8fyMG5OeSB0hhgLsbBanR8DXEmd7
l5fQXV04Qfm8fGQ/lwr4HsD8Byov6yI41nIhyMQXyboKOm74We9bAia5Fdb37UER
4QEdP0xf9/pcYZaeuae98jtpole2K6vU6lYCrQjkyujogWxRwgPFCf2R46bsKSzJ
tzQ8l2CFxgSO7Q6QxlbfSvL2mKIbcJCkLY86VJxdoyUmQuJVMlUzMHBiqlJ7Cn26
FBX5s/JqZmG4bFECIOKCNHPBZVJDut1XcQwwscHcisqMRurmXbTVC9FAHQQhxsfG
O+lzubCZdW54whR/9QSbYfWFt1pa9meCX870U4bSfDb2HoGBEcuHgJMOKNCYADZy
3MxNo7/7scJo0wTcNVfevSt8F1HjC9TvXX1XmSrecN51f2LIvClYvS/iJuCbChnE
6UMLj01jpWdfpp/8UStlGYnjEAeKCuMhuEBI60VOgC3nGEJXBZT1b9lgci8M31mq
x1JAbk3IgQG42SXZDWK1JhKg5ZJBf8Fa8kucywIphmhyZ4wm/jYb0JeQFfL2Wgui
soO/69mLfpD6DdcYhl5VjDeeFFkwrBRsjDF7/w6Rq9/9gZiFsVM3jVLwa8xYEKUT
AcGw7R8vXFKWJJD9GTfR1tdJrmKFqR54zXWD4BOx7NjqO7jjkm8J1aof8ok78PHL
kxgbIhIJORhuNHGVMNZzsWojBh0wgu56rlzfWkZZnFwoL/HCqw90RrheXgZqn3K6
+Omg0RC19mQ1CUSCHm6v+wLWW8Gpjm8sbK+ufWacjaCikIOtUsdE+DZGAY4UDvRP
zhx+liYAb2UvjxSukzTxIXLSFo96lrmlZun6tzTfHJRRhoNSdRKAIdnJyFO+3IiO
aqbciexX7y5qd9bap5uOAxGD4g+N1QtcEMegrQxN+mwLRORyFxV4UnewZuNSGU8A
oe3pZYC8x6vWq5phIVmoS/VKET7TtHUZq7w5aUyRQhsMYaUuj2yF8FMuwI8gzkHM
RvXoNKwJzZNp2bA5oQcLLjslhATe20l4vvcKgG07Cza9dlCGcqn3jx/65h0pT8m6
5C+x3y0bYaPmJbW3doyHwnyRuidh8eEVrxT0ZqbeqlgZaHoPdqJEKXumibWga0aj
K/2caNbOZpTFbb/lYZAtDFXdf/adM+QC1L9yQE4y+lmY+OXU3oXNLg96ipUn7ifq
iHEDE5gtkZ8nTDiKiWFdCrozF6/7BnxDFpk5yAatQZl/TAFI584OcCgwINXueVW/
VFkaxyl9N8/iliWh5wj/Sp21ZmWP6WZV9LbBdg9KTDNrgyMi0U4LQJ7wwikRts7X
yhM0/4Xdf+is1xKt5ClYa8ipLQHT19jSFMXbIU0TkjLZXLRGO+njdi60auCG47sQ
GFL5KQMTkx8QNeK3NWk+8EmWWC5GMXltYPHMHoJ4LJYUXZDBtZLbwrYLNqbJiVo3
IwKGjry6iCBCx5O8iMsn8UIITChBmZDPprKXdAN7lfDVX4air8tYOGVBnmWQMxa7
E1gqGa1/8yx/Wn0Yh9y6R+RxZcbVyDrQWO/m9yPPpIorYGc+rdFjaiZZlg5LtNdl
IDgRD2eSKcegZ00etpeA1o564Dy+BQF+2M9+ZG6HRh6tUkspS/8j4cAJBwJDZ22n
50AasbdFMAh4cNTzkAXEFnLOo3xfz8zR6Y2/9cS3sTRrJa+mF9pgZPJIZzIzxlh4
6yOpg19msxcCg+zeasGj/H1FudJgyklH6fgcmoMFT+MNoZsCcTahPA7IF+tTy4D0
KJS2wCjaF9ujraxxTZWSBEYmNJUtbwvzC74fYu0aov6APJpAY70uoxl9FJCKcWfR
H/feziRepzX6hRgjUv0ur2JEjm/GVaJcuffRYTGy0a+qu2eHEC66NVz+/bchzryA
rSgbAQyXRcRxLzhqZXv4GAKqNAQttGmYt6pPcxV9fcO4YyMhTEK2r+AtW6Dqqq4Q
Zwi00BfcA93ZiqMGkGSi+ywGkdGYxqBQoMJbSN3jmHbY/hYd33g/euxfIIVVLNGG
LcadQjOWkT+G0F99faRQuWSwEr/wXtiSocl+j8RB3rJKbsMZWcZuL/i1FLTxBBVq
mdc3L13g5tY0F4afBdtpTqqHqmbh+yt+G2LWKfDl8KFz+7jScZJyzV0kL+y7srNc
sk4xAOgE+FIrKj52Z8KMpwVOifZv65NVy9Xj991bcY/1VKb+80HjgJb5BQZt6aZz
Yq0vZ0kwyCXOQPuWWSFGThAu7tQE94/bmb2eRDni5yW9S1YQQo47X6pKWiNR3gbZ
F0NydY5zL0dBPIyr0lITP42sWlPfr565VC4FNT3BVX0tSZNU9nfGhD0bSEtUGAy8
CyjmFV5sbnuqV6TT2joQ2e3GZave73jh6YGOyrd/de1PgywSv+nw0frOsI8xGdzh
WeCqPBQPCJJuSAvdtVbTkjFdle6QuLl20y+3ROLMFgeJpFbCZ2zfd5mjqwEyUOw5
knT2XLVTLO5jA+dToAFHT++nRMvtRXT7WJPsfn9A3k2GKLeplQal2RRak0Fjtpoy
K4wutNy02WKFuf2PcGzN4Ce/7onM3jwn90QFvUHNzor1L9vwH3+oUDr60vzrVw4C
qy0r26KoHbsAe9tMGv79a2h8GiKIC5Yc0JmiwfYPq6G/EPX166AZ9gBESEOVn4Bm
83Mf/KkTLvVPSxR4+JQyR6DRpQdBA4XOZVUCrqMc73cbFQ5fW4InczQk+ADXbMwC
DqG2KJGh237MCOfSWvdBdAwOwC5utihhkBQMWIdOVhKgJ2Q85xzjXBPFuc+yco7S
ivMi1JUNJVQ0UityEl5tpOZujtkWJQN4jyN3XKohwuPck3oqbSFHBzuVnLF9Ks4u
wdKu08FrLOGHHQekGZL1A2DHmFM9RTkrVf1PJ3fLROzEUHo2BYoQCqcmMJZHO56g
hJYyt6X/dDKL8/hUeYRh2CuqTj7yCtw4oFfmiIAYigBvxAsQ0AX+zFVzs66T7Fue
QaLRCCyNBDw7TDFGjs9d6KmR+k3W7I/wWq/AxF1vHWzE+hZDGdSDjh67wg08kIml
4A9SeeFlC+rBd6AJE3EYjh3n/z4+CQpjinkFG01ywyUJx7+kMrxXDuj01Y+8yCbI
NKsuByLL0IahoCeeHZxVpKNvR1Hs11nL1j67GGQkrw8Yv7uER/2sXHWAQWk423Hb
VdoCg8a4XYN5H+tHd3tg2Kt0STPcq/t+E6bs5HBo4vqkOe272gvNWX+CMTepYHTd
ayqFDOjd7clTd4gP/iAOntooDBrYQ0BWQIuHiMlSxoPdTAu2/Dk1+1K/URUQw+eQ
Qk7RUfKR3ECLSggehUROEVChmbbLq7EE3MFY9sf/JgGjUJTlmJ1soofCC0fcxjV0
QnEoRBU5w6lWFJz8Uo4Yk6MhBgQgk3TlznU4wXmCc29qVMrsXssLFhjEiG3iLLP3
0QdB5Dv4/JFpEas6kG6VuG07bScqTajwBBcsApzv+p6B1tPmer8HIqS8w94en1k6
1Xa/fuwMCObsTL1MpZCh1hhVcJ6zH7+a7KVuuEXRbF24GwMDQr8VoF1qSkklfByh
fbqCIvtTvQzrbKNgOykbMOzLrINn6vOe2+lQpGB2CTZkTwrKZ1W0B4k0EWLrs7hM
f3sczBK93dO8aoaJeS/qDOX0snAgc6gKbq8R0OEiWRm8g1Cjl5GNQHClSEhnny4C
9T/ZwaozcXjHQa2S90iTnmzW6O33iTmxas7Z/fdCNCvme/HzR1x53Gz0F7Ij8pON
di0GbuRfPkeTqpKWmCvy6AozCJl8/lqe+vXA7zcgD6SvF0Bb2gN1xAHAQ3c/G/o5
QJOyE9mH7SGAGL+CfLL0Nxco5MoyBAkMwZ3QLFN2tBMYLX87BUqIwBYI4Nhb01mp
bsE6EGprKSmbXlc4jM2oDJHWH0lEiVODdOuppOCNQgaetckttCnccoLu83SB4pPO
M/Pfc+/pofJCCBHUnGLHqK4cCbSnKmiBeOto8/gCnS1TTWW00KeST3ckQcDpWhuC
wneFOi7NlGVo5XXNLS1W3O70daJ2cH3H4xBS+c1DcT3pncbdwyHu+ZeHA6+e5uDx
L6a75SW3eRTKnVXkZVWesYL892MT1VD3Phv9Xq/F7eC/k5nybY5fRtiZdNLmgPcY
R2BhqRjhmNorK5YG8OoJjM36JFIVn6zDmhlDRwjb3eUdtuTgeHoj9AFf8W8kth/X
6OesQSGiC9m8hEAfd58ahoAavfTYMg2F3Hl3jUrPw3J1PsMeWcVgS08HzAGS0l8S
U/vT191v90tuc9nMN6ta3Qg4sVeo1Z+S5VQuCy5jbTVfYJcX4u5ry4Z2S/3dA+PP
wjljlPOXypflq6+gEQPM4PoyTIGWrZmIVzco2Aurz5MUriOUvcN01ewXWpH0seRE
2U/W8DVugOHEjpaueCFwAknhS2wsP4/y5mLTkffvOYa9hN7GEeqA58X9huGQgtX9
boF8qVFDtezTZAgfCCrxlnVydGybhK9ceFVv7HJBn8xRxlQ5DDnEVRLAh9ObHbwI
kzs6QG46FZt/v1IjbGjtm0BwPul0NX/gV0+0640HIzrqRKhZZhNdHulSzB0+IZ3u
jN8zXQEqlrcp/dG1vSWs3A==
`protect end_protected
