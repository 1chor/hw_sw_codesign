-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
uoUQ8HSNXhAEDmXZljFacxPTQ/LyAYmEg/HmmDE6VF++3BOoondJarx4nuij2lw2
KR+qORW6ZY3t3omX16UsV3IGW0iDxpIVuVArax5Qnr0ZomGyV8+7lPkG4WRYoT3K
bgA/tEdFqmUzEspkf8y6+cTCFUL1rTLX2D9OUJ5H41Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 49792)
`protect data_block
0711Ru2HMHq6OUq3Il2ptjuT+0k+YndWYMOpSya/O1kLxl5jJcw9MEf6zitkQ23q
FMi3BsVoNeWlV5NU/XkMdpWZ75yyld2DLMyE2DiOi0dv5/rfIQXEvR0H6PyQwNfc
/0JMqSabLMkNQBxmZEN+oonmA1x7rDw2Yu85lYPIKXPfXX721V2fLJjeVLTG43py
62qtof0bprmZ696bj7Aw/aH6kLGrzb4NRRLc6u7BD/ghFgUgpBDLRiyXvze5lsV8
WzQcOnXaou3JOGuZIQ8lgFYnFH/P06r+dtmyNLIy7UbF92e3ZpmNGKFoKgOBHjvb
pb3HBVaEPgladdjc9BItjan2jL83EigrNgBQr0UJ6hW6SnDxTGTlD6DB6as38kzu
G6Dxo9wgw2iojOTH22/ShL3mkMQIf7vbF+01ndhnIEsV4LPuIEFEEq04EwNjItSV
O8zfR3fpIM4bCTqSJM6Nj5tSHit4rc4Gw3H25OBSk97PSrR7GMD5ZqUU7W/7kAxl
pxsfy0brUsG2nsvRkpr2I3wfFQkDyJRrSi0NMpfsO8e7NThuY7w9gxbn+CxYX9Ks
Cv5zm7a+7pX+aee3jUeLW06f2DQBxDRZW7IcpEekTOODlR32k731YYE1/J+7H1B6
MJZy5iWbgzh/tHLmme/m4UUmcbeV1feyV3ldnLOJ1bceGFuAhWx4NBmvY9w8OdxT
asvhdbsPzXCzPEw3fMGVMib18sErySE9xZ7TQlSM2Mb4qyaEoETUEacNP7YWekZQ
s+Fr/vPO2w8jVflSPyid1kNppLiTQmha2ukxOl99Jz3/se4Msh130gJ4xXz3pVOY
0o7XoXcax+LdFYJDitV+2XL2oRWH+Fn3x7+Xq4tMU/6mJS5pOEwG1UGhRfnVAjMC
ooBjwzjOmyNxNtqyFoj8PTPAcvARdDyspEDmweijjT5I9SBS75e2sQrZ0CuVIzPd
sP9fCoOIQNRjkLrVzK1wfVTXZjn3D1oMGDdSxjr8wyXKcuADwnEojeLo7OKuIO2N
8F685JqCrK+e12r/ktNuyGXCZ1TL+8jiF3gmMBewAiQTXrBYC3Vp24rt+n7AFS7u
s4VYQMd+pJPo3R12aH1H+S2kxza+RnxzGclwz7RW0/zMUcpClC7blDTHm+LLmFah
idlwfeGEt2aLArvPqJ+nYbjC8NZXU+WyVMU/ED+xd/r1p3raKp/Fzx1DQ+0D72A8
XBojvYbO10ENhomalj40oSKZOB18Qf3bNfepNwfZ/RMCXNGDUfxEC1sj+3rgakSQ
wX/JS79Iok3pLkQ3csvc+B+XkE9sJVjq+umzpUSqSsdo22dfnTbP2JkaixONit8q
+9DVdYriJAZLgssZTrrZKOKTCF1cqgGtNfWCCRwgcXj87SCOZMYtOW29f7cbZScb
bZvxcZ3sbSZNgZ1lgW47fJ+Gy26Szm7t9zDrM5gdqdcG6XT4oER+P+XFb7IjQWLt
mckvuoxOLraHPbV715TDZqxJVxSYUqabRu7dkCqv1MOLlzgS8ZkRGLGISu94Hfl+
8FKEQLWw3g9YcWqosCdUJB0IWsc0vqDjlJEqEbfwblRIHzTFyl0fRVpE5W0soE5u
tBD1g5tdUBmHINsldojb4YoektJ+M6MbyqU8InNqGmxqrMiHm+SmHxG5BYP2Q4DN
4xoxWVB6d06+hxtyIADWS3+G/3NejpZ1Hg4I/P1KfND5u9lb6uvOMjnRAQ4zfspY
zVhHFP/SCFDhSgm1rV7oORge/rCkHeZAnblP+i2y26Q2VR+bPL8bzkdz37StPBNI
dt4hE5miSSvji5VY3NJuRb6SCOdzVoIIdRTjzsp+l+yciSDE7yfNFWFATVqY8osM
NMEyTpisWFeDMQjWmTQCbEqeLY/NQd1Ibj3Zw6AWQ8xM+Re8MoiHBsr5NUe0+Rqe
BW2chng6+0Y+g6/H/IinbYLn5cYR4Vi1IMc6Zzd0zHYrYJUQJdlC5v2VNbutM7T2
ZWIOIEYZzuvI+xX4i6roNBHy2ctVDLPDPA9UDlUkBytGjTKeCC420IhLmYuDyM5r
1THUl6PVFeHPicCs47oSVY8sNnYYs/TmK0mpXmDLoMi26J9atvkldB2dmC7/I8VA
FQScS8A8aoNUDAzz+X8dTuGjU2UjtILQxZSkX2HzwXfI4YnDv6leFki7NLcgXFLQ
lvaBYxNyIrV874hszfpEiGKpS+GPnxM/+C0sH2mklBWUb3trFRUSktamJEv6iMiL
vW+990MBcjQvdDL0+DoUllMKXYYWasTpWgoswuRv6YNba/h0bwwEBHNqGFYZSWyI
ZuLEio9ZtHFxVGdh1w3Rh4w2GcCWN3aWAxzzz76Fo8jI6LsmyUJe7I/dhAXf9LWC
blb1+Luf4Q9i38Ln1K3bcFHCVHDxtubK1wC4J22oSJBh7ZuvPEKqQ1vjUHoq67Nt
OctxUmkgo+kstfT2ODXE/fHxj+kjIPzmDx3W+dkg1s6o9M7+ENHo+Sptuhr2ULKG
RNYYTagJ9+ourn7Q7VchmfpKg9sDW07iFxt6bIhuVqTxtpjmcArh3tU5NtclyzEb
uWuw9r3yWZ5W+623IBRCdfTTrTQV4HaDjJdKjOEe6gezGIyzS3JykpUyDOicvr1+
RogP85o0GMqr/o2cRWS8DaEWrjaqtXDGRyZUuO0BPx/zh4mLqAapsflTJe8PTcUS
JWlioaQvCgj6JgOIlmf6BEToxl21nZ43uYsephp8Vha0ObCqs3YB1VqGBbhE/m6r
1mqfsUO11c4jdcQJJRujJOBB5RsM7lH1u+tL5kR90QzG99RVtH8qT4HOF3ISsPaF
ccJUp9BdbTKypMpGMl9TYRYHrRc1vKA6Z3NLYwxkPw9XDx22dmhoKcQcucXkUx6X
Ad23ja7qEuuK5FmqBDmYOqADWROejbAGJwHwkc4lyi1k5aMz8KgNdzWLFBXpOToq
wXe/kaPIxpnfO1ixl69W3Zup0BMfXqlNPdsU1uXYyRmksk4CCzT+xlrrGD+tPZgF
qrJc6rtw/ZRrfIgUhFZw2Ej6tKmPwUi9OEZC+JiKYpYwVFWc8/1M5n1cPiyvrunm
104uFYiMoaQ5nrd6piNzcy6vejuSfUnfglZxrjzRsntKlShL0Qc4PQxIu6Gkc+XC
UutR/p+mJT6GpU+zZguP1agKf1IMZWLIpxNbEdHpjJpRyV9JUIyG80a7xruQAmSk
u9Ddp26V+v3ck97y1RcAnTMjDRMZJ02awStTRNOCJ+kXmnQ34ugEweP5PtXgmF4E
zqTsjUFTKJMDUbWwdA1ZdJTerehEnbLlme3CClmoW767+MYx7eeP+MQDFVsB05kw
tYb6ScjZS1z3+96YOWswv6m1h0rc/mf6ZrQ2LRxttXP+TmWKoggCisiiK392QWvO
pxXAsV+bu1AFmkdkTJF35mNX1XgOvT/jnp+0CpKvadpMDrdJNOwhfMjrTwknarLq
8gxJzxG1w+6HU3FirODboOwvgEFrYj3LcSXASvpTgxwSsR/8Lx50Z692jZzYTT6n
Ctnnle6FVyquHqP59i/qTU5wMSaFM9XbgqyVPtUUnsGax4kovzv6zbPOErzlHifa
r2Zx13ecVDI8TMwNrS4Cn1iuc1I3oImpB9kv/yWkf7zXxDGZNLMZDqxSy1+RkXOI
MaPobgnoSZVsYfEeWNeotQ9vEX6S1IPqUKTcWJHLvf8UkxZPVbbqs0gnA8BdLdxM
YoJuLZmxM+X37ssqK4pszd62JofdTaVWZiyvjERweXSMzbPxsg0k7TXEkAs42A82
WTutg8T3vNaMTOltZwNzDbXiqSLtL1NwG1y5lmRhA6LSQAszVZGJjVZcLi3eYRy0
kfH1bafm/TRF47ugVczABQHUO9xMLeDibK6vWk/7ITWow4TasnG0AU7X2+J0FA5n
7bOF1eBm1TNTExcjkY6gXl9+/F8IazOwyRa69Dw5vEgicZd2q1ww/gS4cFaLKs0B
+LFTR1DioSg4y3+QSVvhgl31dUV/MluAnPCNoRkxnNkhNKqxsZdFS4tA2V+13Cnu
sSXUv8Brm8dtCyp13e1AMUz9t2Vfkyrbq61TsREWezBfu3VKgq+LnDuV5eQV1lYt
wMy/KiAjEiFGvXoHIWenXIjMJZ3YSM3rEW6dfmL7E28VyEqSByIm/EthXXxM/hDJ
mTze8zIRAFu0B4QDQJWhUCNyMKbwVXq3A1VnmxROJHV9SEuSAe/YNAqcSCJZcAJg
TlgCKscxMdd2id7FewJYR2dCDMjeEg/r2MIdtsnkzKDXa42AYLKGlkHrajvEy8fM
DuKJuBDhOoublohZ91QPjHGdTFP1wUIMmPsydr7xr4RFDAyX6itnIMnrAdcuuSp6
A9h6vEWLNi46TdoN3kHzRWSRcL5h8ylevUjEYhE0p6ferorCO07Ii8Pk+7vNEDu4
Bw+XtWJP68qgoVWL6Krf1k50wfMzU32snhIzuWWAWBMuBo1COFPUEt2InSX/x51A
rXMCKrN4or9BVU8xaLV09tfIQF4VLH08ForRn88YnHDsEtg1A17Bv8w0/6hGxAW6
5o/Qq2gKSpNoL0lhHHyYuU8FozZHRFBpEsI2LCluRVLkzUEgjLpwSSg4oDM++JWE
n+0aAzq4aTgFuiF1hgwPRBIFQ/uiaYDcqaZD3yHnQaeNJqZZOgv+o+EgMx2My6ib
O/QW87NBSBfEkR9Cq2aaSGR9sxNdNH2CCiDTPbWF87WDUY5thF9a8jcFk5k4Hbg4
pBxgw3CxsVjlvfOInmehQngh9GtdUWNgtiOw28cnEauLfVv95+etKnXZdznkGZWe
Ax8x3RnhdS1oVkxs0xJPyNDZwn/+MKbxEqd/Jz5zYEqWQnV8jFpWT+/Z4K+rjsk9
X8VmPBycQMcaxu01CCxJEuDbMq+Gpfo58TJC2gf5Ypuxtxv/+Y44xSTuCEzxbNYE
Dn3d/gHcb04WXC04aSG6JXY42YO2vb2w5/69oEQXOjx3XYXPL1Ez/qj4MTLxGEZa
a2ZPY0WvNhU0n+Qqx4aD7mrEhTlfioj/CGvVkbX7cUzzw/HNTWjZ20Zhs+/YF3QU
0DDCzpQVW1R2dsoN/awGlpe1qG4lA+YJEA6AA9rNM6IEdcnxFmXSFjaiONeyYCrf
fC7BbyCBdBVlkS/uB89DE85mLmTi8DwF6QxM4bT2HtwVw2HF7kUXOgeaQnWInY2K
xw1iFOIipHK7liUAZYirv9jF0xvQ2Paa8oKlXcxL11yy5qrvHcTy8q5PT9ghItgN
rl8zwIauv9XYMnh5TUMfz1eLVTfw6G3Myy1WKjgtA2vGcQ/r5EIApx9fXCzOzk7N
5710hoNemcHQlP8XD21635nwpFwWS5kmHxaoA3uLSc9gw9CCxLMtdivf6B16mhKs
1DRYBJu2XO9h31f60gemNa8Rpqh6BfOe9lfEc0TJ0Y2wdk0HrdxnH+KDUCElPmBS
fYx00zgMofMzsIlHezxjIZkj4glDIi56rdMqgAQrDnV16u34IkGrHozHzbaacBf6
tNyY2uxRwjT+3TkxxxKJjQTgosHiOdHRw+vpUs9DCJvhloOq1CCBFRzSDxAaBSvz
SWRHgU08uybZT96GUuIDIFfHdbP6aU/vjOKQXV2DU9I2eMs3lrvROSQlN8DwWIkP
27kTFlhMsJkcbSsBC4wIpKFEJabjyRxWGLxXMrLMdLcPkB11lNXZ3ob7yLyYnz6s
sCAayKHAHMEZnZ3nBnnDLzozl90+X5P7mwRZJu461/1kOb/vIv1vx/r9Rf80yECo
u5zScdv+reIhefjckUc0QlV8pK5jScH7jqbSxZLVwWTGcMwoV1PbQLKN8r9syBSx
+c7A9hi1PM+ZE6bLisaP16KGjolYyG+LQQqqYzr4n9q0jfiao8ikLdPzDSspnPKP
9C7kTPhFX8AIw2zT7stfQxdiYcGN2hW2MtyXeAOLd4aSGtphZ6QjlmSi/zsiJXOH
YNIvV4vTQoxFh6GuPx7VRMN9759mm2kHLY1vJrwZUNSa2RQF5w2948JPIRa9RG3o
lRHqBisoLU80Tt+f3VoPUjEIZgjD8V1aN0GuMVtrgmsr0xXFGQQv5v6xcwynRcyQ
CuAkBZ5Hr7Rp6gaVd4nPHcPmv4m667QYlwg9sILFCNsoGFXQrty4IKNMxNxnrLPw
H1kH3K97KwTcpLOr8H8YJLV76EJLvaWlU94GuJKSosUKn19gp1k+NsWIF4a/g5Dv
mXN7XvaXR4GuKYviXFDYktTVEfLFz0Oygwf58CB1fKvvUWxsmR0nxB0N41smOax/
6XsM/8S9gHS8bmpO3JZIbKKnC8T9vI58LiE4NtygbYynP3p+MRGOXdoh0oXPa95C
oxZi82HUztHDKneGjUkqAGAghwldNRW+RBzFTWiLHjltOEGf1aKVfH7Nl5WExINg
2EdHDpwAZBy+6UJbwGBETac/0ZJSvrAbMPjQ7FexYw6p4TODcj0k0vmBmzwzExD7
jt9V/WT3hBxze+1YJVWWpU2dSUfn75+pp0ZSgKkm+hFBPwkvYdYlHn8Xg9wRgRD2
G9lmWPusQZXHY+jJEKvxtpDfh8yJdSfJYJ3+UB+ppsbx5xw8G33EncJzJbKiBErg
jleTweczDe4ILDLXEQ1KXnB1Ybyf4MF7DvV3Pqa9bXbw5oHtD7+ONC4BcYOtUTY0
uym8Pv1enqYkPTJznEd1g7LBivqcrDDOmZSMbIrQ+aQmtQYc4p4epZJGRz56GyM/
Kw7ZH2Zr7o/+sTez86b5lCWkAQ2kYBnk5hi9p1foefbmoflhbUCxCOp1qhT/ZEdn
XAKEZuu3VbKeJ/38lVwXikJzWfLh7G6cYzx8e9/FGCQ18xL9O+va6HUhmoa616Gg
RZwNi4H0YDKbpwfN1gAELBL23ZvF0kLBk5/jfRCgvouat8GMqc1IfqFLmk/3L5/p
D/Vu4LD41olsc8B9zOS2T8CI+jMxiUuo3zFAjgDMltCq9BCCxpwqXbQFKyXBt5FS
xM+h4yEr8e5pHhhU4dtIpfH4lRi8AtKRzwrCF3BJBmaXJg3UY0HO8S+mP2fXJEAA
MXLuGtmVKu7F4QTH31clQby52maDHm9JLtvH5kW6P8mVNhYyIpk24eLXaN8yc0mM
YmBkCcESk+5IbsZWmVS76A3rH7MAjd9fi2P+g/rXE1Csl8fDOin+gXymw7pFC81d
1cMkL7rM7M3YVxDgzIw87d351UmN3GC8mmHdpoeVx4hCA9h2Y8+pjIIgdzQzl9P7
jV1MksomKY4z9PTP2XHKUrAqdVmmWnAo6D6VjAxpNx8PSBsHYPpXOy54M/VlqbAk
aZN/Xy1yfND+EIzGTYbMPHFmkO1pXxSWwI71nrBj4Di6kwdvMtXsyG2K7lUvwtXZ
3yyeJcQEDE+bOHXxq4EpL6HWbHhjc9smiMDLvJQZABsqC/+HuzCGo+OLz0/hIVOY
5evaG3XuUL3iYIGMfOUMGqKzaTz1WVKnx3tffZ4w0qhTexQT5KM48m7Uq1TC9wv3
Xpvx84roTGTN+HrTPoZ+ttmyshvKyxoUUwaVNR2cqeGGbGDyYzpd4tS0ZtzcdU+j
JdHdNkf3nA54twXuxWdc1RKdoaV0NS6gj92anjd0aX51zC3NMycdMMsYljW/hCyI
3SqeqmHnoQZBb5aSm+er/ESOm5ws/h3l0vE9NDHMlLHUYeCS1pTJVIpiwsfkF/XM
VUEq4tGPfm6DUcmCiEU6Q9m1JMM4oB4LTYzHTGid1REg/fFFh2DAaM4nrHCM5jYn
9EW8/ygpAwMWxOWZrCHx4w00zCBtuKqxZO6LDliu4p7x0M3VPWmWVYGS/IZvobFn
/VvuYjEG9iqZhIwc3zJ8YQcE3EFtRBuRPJOtBOgKUUxCfP8Bc7Aot//7Lprfn4KM
YHfF3/Gg81uGVosHXOoERaZypXkWsg+s5sXZH0cPKy+1znuVkmul/f2I2UiJoxkg
vu5MrVTyxBZsWuIL3jd5TnkbiEGPBgUDZlrpJHnQAZVUtFLamBdnu9Y/sSxgV7ke
EdZGFjR7yxduDUz3mpsQNFrhQqQVIsxwFrvlu0aRi/8mKvLiIk8dsLdUDtZgqP8A
yTCbgbuqGyGhyGjRNnHD2j2pIJztOcWmqkuVb1vfLBJRAxl1sk9BGbTSF0y4CITE
uiB6s85tph0/1OCq8UDlg9Bdyfi+vrUWwuW2lU3AIV2ehclCRP6hf+3j8QZeJ811
Kv5R2o8+2BxhStHjRTzVG8b54OMhArsaCmwWNImMRZ/3VoWJ++rGP5AjbtCs8bTI
TsdF/kLVUAEAPiT2XlDlffc5lsRjJaEFi+BY4VNsHSHgIIuhMjLruJC7hoDq99rt
K+O7nhZrMjEqFI3tnapR3P05MLY9+iiAdUIOaegV5prQ7E8HpD7opgsqX0XqCLxN
Ev4AxYn1hCgkU7+u4t2BtrOu2aBIV05jQ/otUq67ATwdkZRaePq0u2wtq5RConn3
OveTEZdChegqeAEg8A7QB4fdlc93+lwbl+oNM9X6xnqE+01c5E10iAUptMcqm4H0
d/XTZCdEvG5SAnwOnXd33/pwcpIMBRdjpBk8W0ljowSdhqcEWW9koWJyxHK5TkWq
ckrPhwXnpcT58ecBPqdssWpxEl7uf3wSWmxVDeF0lLCSzxAkaH+7PCatv2HUClSz
tj+iwnQnsYrUVbMNXtFVKcEXH7DNQMsT3DMoX0Fq41aTaHQNSR5ZwKOauz2yqjzy
IkILnjLovy8kdcrHBiUkGmKWNTgw3h7yrXYeSnfngGxia4l6TahNCzBAt6F5iqqX
ksidwgGCjNbE5uCsgKWkCSK/FS2zbDOVXSwL22c+eVp6el6U05K+3pmRg74szf8T
QeAyAAEtk3XB2nVDk2NJQ6A94QUTv0J4ujB/NxtYcRkE9ov5COsLe/5L6RbuvHra
BlQM8CsEHrfb/5QNmhHrMhaj1V8VI3l2ZcXWn1xD/3UQ4enujrL4zrfnX5Ej6tdz
3rxG0OYaSnalqqu6nc11ihPWOQq2nFQmojmtrSsxfzuPulpv4Po6ez3rFzyIgwvu
t/5N2GNDlGpaunWxcOwWuHh+oOlTt8ZQcRhNLprzyEwFiSrNAqEGfl9sxQw2gK8J
zVMUcJ5LcKjofQAcFyBtC4SIPzzlfOO5TxO0PSoQjINPegXRLAmKI/8YHaGeqQN9
+EgPmPyaZwjBBLKRzIfwpaql7e2qcJkqhi8kJ5AEtf9e+woy4joPw5ruuFf2VO95
Jh6zcHfAz1lAPuRUDyxiVRzeQwv8V71wPnbk1q7ePdywnT5nQEBWB+hOZd0BvK+L
8S07QyYeotUons/vf4hcLkf4xc8IU558LaStSaicp1dXrqVKX2UCiLpkoNZ/wcYr
fKe/NYtiVuA0rrAZuVybUNoWXNBtRb1R8jqYF/zWSN97Nox+XXA3e22Y9JL9Pkv6
6kBtcDapRFhPdaZEx/St9PyNXRWr4htT75s0MHzu1oXR0ITc1jiX+DtQo58/LBpz
QrOMZzXhTjFSbQoIFkGUsmzWidrbWuTUHj4XioW36oa5WfPSzWd+ulEjnoEu52Us
DB9vzewAIC6StDnJ3P9XEzvxsB6vzuwtO8QfJrTG2lRc3FfG7X32gd8swIhxbEy1
UdX6RcljoFsm7osMJKq7tlgo60faGBYWXWfxod6MVu1a/DPuYIoG9Bo3uBsVr4x6
8jAzLCC+wUsROTxb4ETU7jLTzvEcH84hw4MbOTEghCwL1QQ+LyYn/nO7/8i++VtZ
idSn8n/yKWrRjNJpMvICmwbvyxKD0CLBfVGb+frhLC9frJdmDOSqAXyREGJ18Ror
zxBTGouN8pPM3ZEl2PvENlTUJsPwV4OfCKKdOcjT4ibchrGNrmPTcs7TmsqCQXkk
omG7o9Ei2X85gwx/Un1UVZRT7iAmdFZmdF0gTcM2zbMkiMDr6FmV4W7yGYm205yH
WBLT7H6tT0Tek2lmIldRZCzbcfBae9b1B2D2yRQYpnRgQ34b2X5Xk6YVyw/IGB4h
+vyrtHQPLZKy47UsffgQOrpUXqKLhfGpHTc8oqYaqLoHal9hoXveS2/LodCB33l+
ni5kT6Wz34/rIYZ7RpIXhxTdGnuUATl97M+KZ3c/qd+y5PhcuZSgaPPOxSLKAHh/
/g/RyZCEEH4mw2z2NPzp8rP+1ihIQpIf8MolqZTI5XIACCYrt1G/0wnJo8fYeXLb
y/Edc/0pj58fW68P8Q8qSMbeB2bv/WDPM4l9BSp9F3EL46XC7ZNUlCaQx1bF1TYF
l6yrK/Uefg6wqTKtY0eXbvr6jVwyl0oCNI/REPl+L50LlR4fr5aMvRdb7dUJotf9
gyaXzJqfQ1hh3vjEP+MenbeTbNM1ZMFtxXy5fWD5YY6fY5r/hGiZC4nCPVbJNQ7z
VV74emlvcm3Xj53lU+RxTWrqG9CDP83l+hWwQkliNrKUfzEErVa2qd7/1P55pP0i
3H+eJmqNcC2XwXTGLPx7k2lQ4oqkWJv9yMlyYiBgCfwljHRrdZYcr8gYf2RNyEE7
7Mz73XjmK5Gl2vkqpElySddyDI1rta5kCkJ66ALmZakDJDz16jT1vJPwxa2x3EyO
Ickz3FzRpCyXo7z2Ao/DaVFIqA3XI4aQFoBHQNApUwf4grc54LL41mYWZRhaVLC4
YqEsUtM1i6P4CP7tCfi4j5FTiDMe5MrwxgF0KOJ35us3LymKBnJMsXfhQUrI/Due
XDzTx36J9wLvmSz8471jI7/NAZYzQcZ99TtXes3TnFkGQqVIDmcrIqGI3jMI4kYQ
9RomKaHUzQHoGCH3/DjvWVyFgQtfHuX4ekmmqsj/NS2BZ8K4QV3nWzeuXlu4SmN3
AYkGfqODdClG0aCi0kryyRw3Dup4MsgDNEIQ3U1ygymk1l6Apsq22otAc683trSQ
LczHq2yVFa2jtBrFH5tDNQDAq7hESqOoGpW8wSHDJmf6R5MJgI6cowiOkYs33cN+
rkSvo4mdGhHsWl3KLLrTBaGjuBpN1PsO2/ZuaMEiGqfFXQSaXpO8i3T5nfPfl/nE
NcIeTVGMHRWQEPZnwIi+dTgSdOwhsp5CPi+bS2rar+YFpC38gwd+UHUQtRzm6985
qi6eesUbKTc4KHkhyWy6QGuATxOjqm8x/PyQ54SmRYgqrxdTF3OtxFFwNne6EJ0j
DSpRKUAa2iLqW0+tyW8CZZkinSSFMso3dufT5j1f8Ak/aOUirC2vyudB+pa7Zqb+
kFPB27ZkeeNEoRCrD5oYYNQPKaCeYq53pQqIXBjovvqXte3aGfGuOFI6VubzQ/wX
3+YF0FRfkVCpm5UEdjPDmPKUKrZhQiqgqG3zYTsRcA4qIDGiT3w2qd9JLglAHmRe
Kxw8zcbged6YNB3rjMPotblOCsFkS3tqRk8JeHtBLwJtDSMXrxCg8FeP299Dmcvp
KLDcrzuJdkVTbMgmCfjOPoAMg++C+AY+fqu66QgQKpPgCJXrTMPRuzLP70RPsXOT
GFNT97HKznw0OVaMgZt/BMwdLxepqHAqmIaelWS2VcjfoDDvKIU6vdHKMdZPazVB
r8QmDw3Jv6Z/K7fc8RWKRdNQ2ke8NSy42cSOeA2t1oji1ch/brUiJJSuM5HPxP+Z
50TxFe/BKC4+QPayFW0nN4J341irLwKsFbRNQ2plmsGICAC9UQb2vUfrBuS5VqiN
kjyNzTedW6/lsrgqoi7UJwVDf4ie6jiSQAWwmd7FlpIzGrUMxULan5bRSi1rT1Xs
hXOaBd9wpcjF+TeuiinjSaw8PwOkYxmTRXw3zGyUEpTJiEGpPVO4pt7RuUurgoK/
oSjj+AcnaYxrazXSTsulKQx4CF+Q4KTMn/TLHJFu0hfc9rkSqN3gim1xyRTz5DEo
e14mFx8faPmckPuxzWbB1bWcMX+34EUe1Z90nsX5mQvalTy7PYXB0316U6wh9gmR
/hbRtNRJvfD6t7dFkdCICJkHP3LGdlVZVi9IqMcSk/xAoDFNyJZyHv04Lz7u3qQ/
/vjIB8z8JeBsalK3T5l/gfoG7xXlS9pIBFdkPeujioQA9KT2cQGxFF727etGFJQc
tPj4+BfDEd9aqtt8TY5mZ6HNk8ZjknH5Jd9KgZYw60GDoHEkRTktmx0NjeFudMq4
PtbAfMNPnH9ku2zx6A5D/jWKKfKCLmOYhQLSYxYmTcidvGrCu0WiCQKl5frrHF6R
uUHgNhmCY3SYOw7V07rmzjeS54SQsUrDMZw89gxYqWdTiqJ5zEMmKjJPU4u8IT1f
PdzAb6ucZEhkCNdvfzBaW3Id0NLqHiwjLgkBvb3Co6ovqgVET3dW8ExU8+PIVGL3
p2+YmyfiO9l9qrFJnZqZ+Vd6J41Zs7KGlMtT1kKcjN2f88AtmidV9uLpVt82F511
AteKEraRoIu0/lD2tEuFnSl+CqKx7Z2dwS0kT5oZJdViisRy2lcjcBDiPKdU/67a
XM21gTdS9EgjDPSevPqBA3XEzc1da3RQPOTbp4t/p3azwlHxrqvQTLZhH65JoPj9
NANgoFWNVSo+cKEZyYYbxKF0Liw3JJHe8x5NjChdRgzzBrv7mnlxlaA1xND2QFBO
xJifemeJ4ZjsRqNsCiTYQFA3prMSNF/LQnYWSsQwj8J2OI8Gmt/2FzMc7BHk4INL
DzEtbjMl7bh2/xO/eLp2kwvXNDI5IuLsQI7TK31gWumwZxSJV49yi+zEKVAKRHyb
05u6f3gBr/0fYBjiM7ASC/DQddgFN3BMjdYPsHtDpas/1URrXNTaRLkdqjaxbY9X
DPtFb7Jd8gEFJT7dYEXy+Ql6fervKPFOaKusljTj7XhmzlrnmQwmNyZOzzj7USvl
ItewUjcA9/ECV9sxrEzfVXAqjm6hlMT2j2Cll9P89U6FtKHbwN+zkJa7WXkBGmhe
63smHlQUKqEqjrkW370gC0YuTIEkgpY1dbo2aAwObJhUkRJXJDTBqPIiz9dZE00V
rfDGby8JbxjSSgjxdrwMihrUqp6rYFeYICd0y5t+rhwlw82NePPbRuWhZMDMCEWk
LEQgepMKcaUEjjPTXURb1Ao0US4VwLnOi7qvcrFLRzp3gbH3lsNMEPsEx7+zGi37
gnT3lujec846ZLnLWvDwaq1zEHBOMSxU1NfQqKLkIDJ2uEtDQwCOA/bqKftTux1C
a+yHH3YjD+PROoIrDMfjg6nHcXQ5lTBr48xr+JRj+Az6M87nZaFOh2KuYsvDlRkj
7MPMPtLpTFSEezD/8QZhkn9UnjVWvlK7G1Bsm6pkfdnUu2AudldkMQAc5D7f0v5K
1c6Obn4FCRbl9+x9RWYlgeFNgTG3uxNKyITCQ+nzh162e7vC9KL6Ynh8+JROOfoc
gI5KsrYlxKIhCs+N3hgnhVH3gUqZ9147Dso4l9omwEHTbErTZIXTuXMmZdPMVQMH
j0ydhvLOLTqP26iY0hxPct27tp8d3D5he44LK5spT6wKN5FCMFKxsFUSs9+oK3UL
IQvAnlB22qwNv7hVqidjqdqf62CZKqyKSS4Sp/fttLEba+n4Kuds93gSmgx5UVb2
eS+oAIlOfXOL/A5vTOD1RGaGauCwjodLjUlKb56cabCVCdfF2QNrINHzVkY/s39C
NBCHSqaPQaOYbk+MEn5irTUTm+5d1NarBfeT2nvaVx02X+fdJqgdt65jCMALeJ46
ZSsKCwecQBRnGW0VkQngSrMrKPwrgSinwEMAZRz/5gzQSaNAjhDQMiL9SzNmBEHc
l/0+f/ghAKq5eZy7w4bldMWc1TbI0+pr7gY5fcjXFBbq9W7nzwcm/Lx1/NnwjdX7
W3m+bfnPJxGvhK7t5g0fSzAO3MtEmREb99dnv9hhaUG3Aas80OyrjdjGuLwMx88S
KCeXE6bQE+9MdzVQ02jUlsRv0vfFfOi4pVZuKXm6OEg+9MNINLEzHXoZcAumW+V0
NeCWWvJZ6taPKRF5I1d/WIuevUpw4z426mP+GRvSW7cS0NIJykPEraOGP2hi/42h
4FFiwTceAdx4S6oa46qM4PQH73bK96fGknYdE8gpGHMaBoHIS5aWrNwoaC+OfWMq
WTVpwdkIpYzzrX0J37y7m8wg0sxndIT8N2tkCq/gTmUXNGzz7cLEY3pUz09+WDAT
d2quidAiIEr7YBKKlW4KL9eQHkft860ftm3YMbw9oUEnAnknRGr0mnmQXu1Pfogb
6u4IyAU3sfDKoDJ9bAF6wj5kIvs6oppzPliC9RIaWcdheoB3VVa4uYFUhzp0A2C0
SdwZnnqMnSdctNuF+Ji+n0WUBTNylOvxlj1igWy/XAxthtHbDAEEaeaVj9ArcdFK
Koyde8uFDMcfCdABa2YQL+rjcPBIVuEIAaxpnd7pefxD8BBTt5eIQKtnahlJh2Cp
9I1ZR6G7pQl1Yp5WQj5LA9Kye3yjbbypdxDBzmugaPQqV9gVaPSI+ECvlRDLsYKN
zU3uvZ6h4cAZPTit8JPlOFKz3IpQl3dmlROeAFby6t/H+81oOwOXPJJDno/nxWuH
xaLidhen+LxFP3jbQnWkF5TBdKA3sTKK5y6FPLnibo/c2Many/011U7mwsPEbGF4
iyA6FHCIFPI4f2cUeN66AsJIfa0J7LFmsY8ZaXk29irBXIqf0zC37G1r1c2L66Q+
ZshGa0vP6efn3Ed6C/T2hu0rDabjnQ+RL5br+hZJexnPb7CPpkcv0FWUflPVoRpp
i2uPDgshldQtMomSqDQQyGoE44+bSarmTFBVNRYoppKPheS3MHfBz1M9VxZHrkDB
YV0mXNVtM+NdnaDeW77OJvXfvRQd01MlCYFH4Wb2AGPtMHf+qigQnfT4WmxSGS6x
YWlhINqOzjRjvcivCUgwY44Q617GHrepsjewZLd7+B+MbNVQl4mafVTw0mB8zX7j
stAF7WVIMUGCATL1J4GpIGvtR/lTWlHg47afmBFtudECozqP+MvGgw4wcqQw5wTO
0MdwEroXzrqQ6OiHzvU0x24pjtpHVHOgRtnu4/eLxCpWwMLojrBzsVqItG0BAR5i
p5pEzPU0SV9tOXn2qSkRA0GErKWP2oOyoT+oRYJnFHE4ppCXd4haDC8ts5dELp/2
1MXmqG7k9kVMVQMy93DalXIFPvAZl7MedZq3rpR/1jRbkXVF5vh3HiBUj4dN0H+/
covXkMYgS42JdECcnfvXHw2WRA39IS7VAkgWLMXgXSK5wsAt6S7b8fs6D5cjUUif
XfurhKmq4SLREkM91K6hdacc1xBqXQdOcRGdaC1ti8NWQ3o/pM65M+XuxbkQ4py+
RcIV5Hnp1bJeRoctozFD1Gz0Jhr4kvrD3vuOPGVwBJR74TqOPbYv5HiHLuH11N72
fXyhFifJRKgQEQyV3r3U5ibGFEgZwPTPN3sAjStvquF5Itk8OtGbIJlnlnoVbKU9
VZg41ViirhRzd0l52XXvnzBQlX1glMGzkqmFYdhS2AppMrM/DzaV9cAadr3l4u96
vJNORXHZ5io83LQfB91R6Q1sUBeVW+L+boNTKnWeLwZbMZR0tob1fXE+eNSPopHs
IBND6k5M5m9dPifETxnm1y0sbPfrSRnZZzW1Ve369U86RaeEs32uzu0p8Px5DoIX
uJnG/wsZO3syslOdJOIdAXaiA7/azAEmqu7iPkEy5vlE/Rc0mLZ1U7Por4FGYiG4
gBe4olyvZTt0Pt5HGKErxoeCfsu/+3KUXGrZqhY7PlZchl0BZ+ING/B/xe1tiYta
nDSTyq23+1bEEzna5CmMCssszo54xM988Nu/nnR+d2HW6CrrK+EjNDWGYePhoyni
u/86FIxJEuzVfCWyiTjcu6urtUzLuukMH48HYdnGSG2Y3GiS0GjyK4A4tEzOzUjR
vjlB3X+a9mbU3M3UFEfRrpv/aZvu4siLRXCr/fnQENSfAfpMvcVHdYcrB5VeVQ6h
wPjAubr4euaGZV9tVoCrCCapLI1W2+n+z7pVE2FMEj84PC/ZrsjBwh6rz0wio8In
N2oyNPI7UI78GWExphy8h4X0NubBtBfIaesJSTZJ+IQX4epUvNvwNQcHJ/POiou0
IAK1AjWPGDGwhWYyONTyCm9cwbocz0UlSpFJfUfjPTKoaZ/hat54/B/Hvz+C6OeQ
EONZb8yd5F7diWjft71HLC/Jsgtg0lafxVY2jKssIX5X/J9tjANRjpDI2nWxkhtl
zqcJP9FI2pybsNq8/ogyut5IfwyeVDHbp6MbR7OZo3n154NVyMejC6B02fo6pWFe
4ASlfJWUbYRYf/2rtREqKBRbI5y7/iQBvd4meowFJtU5VxqclO0dtvPQHU2BU+Ea
t5WjQvIpg/8ZNZyMQt98NdlimEQKvIFtl3+HYepeSJl+j7T9I1qzQOmUmuwxMs7j
jas2HQcb+vRANajamloXBX4saiOqPUmcfMeEiyKbYJKQO408JHyj5XLFSdM61g9q
OYP4dHrogxV+4zGIQnIvtxhxQ63bKxb3qcPVh26V635jcAW4IX541jZgdRolyovG
EIpciUZthogm2UOD20NcHOw8CKnX/9bX/sMxq/OMTKfTUf995OgnG+XvBMZAOKhn
1ktV0SLVM62GLyf4mQK5uDMkZf7Wc8zPDAB52GKM9KJ3Tbamy9ZqYz9Ka6u7pPtv
u5YlkcgMEBLAxFwcJYim+/JLKtqLJq7zzJqsF7PQrDR+bUuu2R+/sAwBu/L6es65
kNeNSnKOCdwXVIRn2dqmGcjIw+2STeb+FpHMT6fsZ8rlrf/vjLccuslp6W2A6nTF
2fbd3LgHh5T134+DjU40NxtnPpMaWexOvpu9ToIzVBJgVVhfC9Tb+rqGvVQP655Y
eRM3vQfBsLFUSSGsUvcrFopkGXSQSlWTOwZ+MHP37WHc/jidq2PeM3JEvYEBut/s
uEncJhrJKxwtkFoWKEzNvvtH9bSBcXc+KzQcK5P/oL0P/omD5a9OuxXK9cyQeBdL
Re0J/HfqsbO3VkT9wL1ZTiCx0Dx0EqC99gUtgnBBAVVKbMp/Emw0BiISBaQX8A4z
jOiuGMW43qMKuFHBPhNDTNogOuOQN1TUvf8jUMMDOEPDihOJ3aMGwetbsmdM22jO
l4+3RJWtermtM/DP8xuPBnzpDdeoF7oKa3NM8feup5zkMxIDqjlXdH19saA4rs4z
TbCipbbKm645jgmoMhsC2saOaj6GQOTlAK5ddx3VsOC8VP2DLYnOPIFUHflNeX/f
nELsDhbd3hP5g2wjeLScYiYwO/a7FWn459P3Vz43/eZcSXb61pA/PQwV9uYFuFCt
yN/P1om2JTyeu4eI1i3588Djin7hr9H8ykfyBl1+QsSyj4zqP6w1xspN3MZzL1We
+zRDGlWNdy6v0GteGEpo6Ox1Glq3tVpOhBblD3OdA9TpkXzPTA/DlK5MDYe0fj7E
nKZNbQKb6j1AiZuOBK/uyJ00/SCQHCfMA0cgzQkH7LvT+yz5FOJEWFGpOgDxt+uF
GwqJEHuXsjl/QrlVJKWKlNixy3Ccp8GxqMm4q8ZEQVsjHMupwAFCJLxbKfW/7CAl
XHryJAXY1ZOgTg+Zq/AAABWt2aSNizANpusBwmu+ovcFzIg2xWWIJnQs6WDGU9r+
U3ZK+4nqiAJMRPHNEpoemM6bUBobbUzSSJSDOkPT5stT1nClrTfGxuv7QJx9YfWR
EGRMRMKp+Qr5VeTNUJXbRbcrGFqvsK9LK1MLFfgq71K3RJ4dcGq1SLw3E1gVz6tZ
sn+9PnYoOb1dGvlCDb5LPYTcvrUzrHi6DlzNuVXHwDthzT+xs47ziWn+NkAJ658V
K0CZr6LE4Uxoe40n0OFjdVL+uTfdQAwUvnayucQxWNqsxRwPI8cvlmeVB0L8NZCn
g3BBciMe91J6bg9c9NeE8h5vhOdahu2sHKfa2bQsUz11p1MKdPb02WbbnOEet3yn
4qcnP610c+bDAz0hBK6ml50pdXJlAYS5C6UtP2kJnucp/zxxgLQ4qo62HFxwUZBp
B2WwS5JpOuwsE26UmtwP0b1ajf2sPOdC/N1KyOWbh+HrUeHehp4vzm9lzT+VZfh+
9Ib0aBxcqLXsmcZZxqaUmAMcbm4Ep+LtLUuMyrD9BeMmUcBJ5CnS0LL1pVSxsj5j
4eK3+N/CGUZPLCd5ruk7zYzj5g0YaIzObnnlRa8vR2ufJFTNYMcsjXsK/9IbKHby
I8tkdrfL2aWqZThQaLrNbWM/kzXLZrbnhza9pEFMQ/hzeKulUUGPLkm2xYrRDTPl
0JD8UrNhTfoPxGqHzkjOykGsr2KMlmvbQQUFGIaxZol/F/tAwjgRY16uLyHWBYbo
+AyruzGZIXfHaspEdNF8dYP4R/xADYW0tdCd88eQh/8lZTMzMgKAzhaVHRfYufQQ
ycBbMBSMVbFjsaYg90mXmIh8f+PDAGxnT2yLqAOOoeLhtDKiACC4iI8Zn0IZSG8L
trkKNx+L85O/uy97W76o16itWO7ORyW70Kg1F+9wrXRGD5xdbYGPEXeTb3+pQ5ik
zFVom7p32Ly6hlB+NUYm0QKcaPQAB2LQTNLWA1/CvE57WO4ch6rRAEA/gypmHDbj
QFPUe8+M18sB69675XbhXgklBVNhaF7L9bX0XDx1QqaLGRqGgJSbmf/iGsoCu4r0
kUXvEFPUcJyJn2Y4A4KHFuhbBXioELtMmv5qL4d7ruSOPTBe21Ycv003UXen8s/h
pdWDWV/aFSLNnHC3L59jrgXGGsDDlI3jNi4hOBM+e+QDDE6oeQZrU/v41lBhrZ89
OaMUjHy02uZJqWYj62FcPEw5OyBDjcRv/iyJqMi/prnApVAmWXDSgQf1VlkxW9Eb
lMY6feB5cZyMSjw544JpOTwUGjRbv354V3oPN3mcxUhshuCZ8kleLa4UP0KxBEG/
mfLwJPIbhvTYbKr6H+0a1/83MJQUvPBiK9t9/LIPOLqVGsn0aFnScAlc5o1qNePt
lr42yI915ShE96dPESf3vkjGVdzsh3/NlMksipBT2k1Lws7ve+XNRlhTM79+Ra+M
v/Uo6giYbzTYU5L9Mt1rLqiwFJuyieidKP5hwJitQ2bPXeSI+nNsroqsBieYRc4N
WlIhRIyPs4j2g0pf4IY5wgDl3FTLaO98bmvvEMbu7H6e8j4o+j6sDlOgqOxrA65j
pA3qeV6sLOVfltHCX7+54flRXPhOi2qxAyxOJIXi2O1dBadBUDnjoz5ZoxbUzvcE
j6/mZJl/Voy6lPKSRuTsAL2hnFQIJRpu3cZSmwpDf2Nu6VSTb12LQehztDMFojN3
FkBPRjdZekOh/oK9UqAT+WfAyoMHOV/AWjlYQWIPcLHWnFgRzAdPGHO9dJyDgV9O
A1uYuMkZk3cU20zLV3woOC1yJsEeefnOVmd1DMyNGbe69yv0kNKt3IOPqUFkzG44
0ydRGS3B2/+dLy+nJfLSoZ/g1ro0CDLuXmiSKsPO7prM60+DR5Tj3LHyVIv0a4Nn
PpzqkJAoEXcqxAhmFlqi2EfgvaiQ9vEr6AHk2SwRz4U1KOaoaadh6TqoYEDnzeCk
IT+cr+NqU/6tdJoXj4vvEpbbR7DdI4Rm+SOrPC5Za7LpGT2hvWYLS2ril5pWnJf7
NLsS2L2dH9aejGFZjvV0iITy4ORgxLkOxPf3N18WTPpCHuHMaHzlpDQZbFjBLVFF
99L1+aeVZ3Obt4UYD0dBQIKBf6+4jiWJSpFmGWv+Iqgun4EXCKdldyx2Vkwignrt
0N0gd6wqfmvX1PgccJJfd64QcU78xD8YqQb3HQkjHyVqErkvOO2x6j6UIN4FGweR
wqSI8V9NUP9lSfHi0zZeKdfO79R6OyEzWSd4VVYlVC/GLhhaQPrC9koyvIwxK3cJ
O/RevsWJxk8TEfQkc9cTNT0R0ZdPa4UK853DKYH2A4N35HWoq/lzx1YCUOZ3jPFE
Nb2ug8U8Vfprj/yHplLptSAKiK9Gr6vu7TsJm+CvW4wRCytcDeW8nwl+0NWbw15g
FBdbIIIBE41I+PyFoDciC3T5mc71WdSQKeUKtL3+ypnUs4pZ2g0qP5/MVSnBDebx
eBlxsCkWtPXeN+7tSIzFmIMzkg76FD5HOLnU5g/dUVfEX86F28ubIJxPITQ8QR3S
vNSlobDhLAs5erWcfElmjeNeU6YBX2DmJnE0OtbFHt14/Q5UGVj7gbYWTH3QaJcO
kVxoqFLHvmZLRtygPDmcu4IuqizFUsSkUDqDNVsDaZRxEYtGjAAXHfgBDxMVvpFG
wL+pYbA8Bp4wvdB+zdV8aDd/ta73SA5+nohvrb+IlROquMgzlFjQ/tN90Vjda0C8
H05ey229lFllvCdKDTx2YzMOCwooodvDATak+eNxrt/3rAMnR8kpqGE6OI4xyuC5
FdteA6+sIWeszCatXY79SN25yEt4Ww41p4Bnt/7kvB3eFlAiLwyVVa0s0sfbW4PD
fuobuOuTc4gTmUjpxs1F8ZN2+D6HvO+Q4Mmk230FroFyc5PkeU7m2gVDTPdkKf2t
EASf1CMv78lpOcHs5Ns44zjzLdF7wHraUPFZy9C5MJiob5CjQ1f1FcW8AHHCJqsV
OH+HsTbeFQ41iGVPnLsVvGMYnTDsszMSqPRsU4y08XyW18v8AIRzc+76YrgTReak
HrcmoMX1H0SmTJkHN4tq3yozUijpx9Xw252OH4+KgfZ/9d6MZ79tfW89emnyYFFb
IHtaCKUgUuzEDF4iQlLBE3OpBja7oweWW8S44C+RfGOiw+oNueNf7uxj25ma6zll
PRp/3P90Hy1LSPLtMJa8gwa6Bj35/Wdzwdicm/kvRY0ThcA8MCI1YE4IVAxYptzR
wRdCD3V+bp3/h9/Fwi9Qmlfx6xaaaoEyijzN14fjN1TWGZ4LZy1l11daAfWY3Yzt
Lfdnkm3A4XjxBWTAS2sg6YpqltjqLxncgDeLtUFXlIXNzOguSMdrtLkoyXkhim4F
U3A0UbY3M4ZbYLx2DB4gSddW8JOw/xwPYfcz6hABzY9QQXA5PqAWbWTLM+fjh9X5
bk3a/wKvcoNmbwWS19/bI82ilAIyPp4B20e2JenH8S2D76Y+zaSy8xlRe5AFpwP3
ASK+y+C8N2tx9CI0v86xN2Gq0HMd0RGltWwt6qluMVNyukijqiLoGYbFrYnJD0ij
HiojtMKKoWocElD1pQSmDHUoiYhtmZwTxOvxGsVthNzks6MzAJh6vvmVALpZ7wis
j4SzNVO4giMsKcXcxt+WEAnq2GWfS2J5POABBziIxEO1FX9DraLnhjLZNvn0mbN2
CAtItx0XY5aom6CcaST+rB3Nv0HmoJJxs8IoWX8lHGct2GOkfjAdGU/brL6c7WQV
z/52mHVPKYhTGxs9Q6jzhs4PG9pqESggMZ9wKl+cdVLCFAxRJw/Kc7Yo9Go6jLgf
4wLMLgUGVQbdqR4qVdYJzfLZAIyGwS2HYcbxJeX5oQtiXUb5joxYKU6d52AOjmpW
UKFIhrQzva6ZIk4oZqfFnMaLDsZ90d/U3a1dARzlP+MqmbxHUtYuC5K3HFKlcz7B
c4e3BBSaO/aXnS6MsbJDPiLf6dfE5FRM1qPBYjOiCTOpjfANYDJzeu8MiQt0U0fG
9HU11OwTtu/yKz4EVkykeIBpH0rWY8WJZvBeOsC2s15iXfNshzMh4czXReUluYdh
2BYjA1KA6dtYpzGoTveGI93CDAVPBv3GnzjxGK2N6B9tgbF67aqI6KMXC9LEjpkF
8Adqh2GBf772K2ZZ+/IP2Skk6/SOPmFlE7JHrAozyO3nQpF5xinEjQMUjD2sG+W1
ZYI+xY/LzVA/1rdFK6M5m6pT2HzjKaoJDl1nvt4+MZqdgElfCAq0VcN7mBhgx4dq
/v/1md0XeFsmOwtyc2fNqneTC6wI8slGWfpsONgzPpmpYWSXLilGlsuEXVums6pS
nfzn1D0G02b96KtU1zdmMDX/HVi94/vnSxTHNGuNCuoHEpbmd3/rGFrTnQ3HUpS9
PrU6JGs0+6xZMDqytaB8B+RJQ2yqLjgNCA4xio8TBMFJW69rLKHZe6Ze7R8KlPSa
QotNDhr4Xh2aYs4EMUzxyrIoaBywx2UWYzV76wJ1KeGof4ReD2vFYrany3IQtjZh
CRnPSS9mBk8v6qLjR4my8+plAZQyzaoXk+uAn892KzocOmOSDqUYgWAP5gDwXTGM
T/7M7G1aVleh2+LnWbloO1svbDUOyzI5rCb6F4RgXZdpZ1t23ihCMXt8pZT9whtf
C4bg/QwJqm8PP2Bz4uYxhJ3mSvU2NTSM9AqrjjgItjsOp7DIMPGBJUzytnfR8QX1
seeGSvJZxy/OPkStMgfh+PkVdOaSrX7rtF+pDr8Nd9moQSG1qQcOgzLgOjQ//BOn
RF4UfrcehMZlnOUh1Hnmnk1wZ7vv8ssBicsleLXhRUAoZZWHEEGztucX8VXqfuFS
rdFZOuOgici4+r5sj+ODFNQhOTFcTAAq5Hyd1voLFsCytDoMvZHGoG7bgqo8D/1V
s0hbU7DvO0Gep/48H1N7/BKq7EKI4QuI3EmKIHiZqxanzhMJUvqcP2xu4NKRV50+
/oNR8y+iF/aaZ+pcoQIVIlahKOC5jk1f7g266oXporFzja9VVjzaJVm4+n1mOp6d
MhohH01HhM5uiIDfLMoD5IMBTi/19pjREsr+iyV1qZNgWWNZE1qHq5U/OHbx24Z0
jEPmFHNOOnb0zKkPlLif8MKSEpW2h18gKeymukJmQTqprzkHNf8m+QH0oNceeL+X
1r5IcxOPxsMZVbZDGMmWVFp57xSf+odpl03h5qKkoW+Tx6NUbDgBIH0NTY+dZlHS
2q+aXZSzI6ud4YaUSfQmtvGuD2qlMdwNC8OPW86UWBbzYrTr1kMverLh+sS+dvXH
1uKRORPSHBcNNGqdo2abIMGrYHeZK5UhUPVjWax+VTX+Fzhqd6bHJvI+PQQLGawq
PbRiJXq4BDfAiZ6orXpSbbC97J6//Ii/196CO2bNS/CRaCi1hbgxZQHZTt6Vsl32
EAqL8nHFYUt2nqxG7VGEjJSVDmDNOjZohinLPyopTRG3hqHUDID2QcSI9QxtyX74
Uhgs4WY6dARpY4AwnTx/A4WkGYNtt3bWpIUPVedabzliVn60dpaz+2xEJXIhJjF0
1iaLMeAprBfIm3kTiAogDthU0xG+v9/njuO2zUaPqrYQZ1S7eGwU9rnnq2VeUJw9
Od50bUGm7aHHrywhGsgXBKH7F3eYdhbUAliASYyGWe6MIvoCMXLpT5bBpA9LWrF0
PvQx0vDf+eZX2Y4w4IL4hSWmZQU4tx0Tjkl6rqrKZOpQtHLOaWPDD3BeswYc2pHY
Xu9SzdOvyQJYjIK8nELFSHKGpZTFSA0sXO3szfwQd2xHJ18dRxuFXcb3RqMsrBja
opfhzbVIk+t/LQ2gkRcZ1ZUzAVEnfFtOTnVv6YbPLvbMr0kqgqLHqdaqqV0PG9J/
cCmhQk1RmGOUFYt7D+XQIiwlZfoN1U2ZjbXlKDPJCo2BCc+4JXriTe4WAprnSRnI
JmkByLoTo6IPot7zBcU0QwAirkq4aGKGDyxH5PEuHMQ6e+l4KRphDLYIJvimZod9
LCsgjdC85Vv2b0dajtYF62+4akYdDa6nOAKE8HhbbrA1jtQnF3snZyEBowTo/Luh
0bqk+WwyUY2TEj4k9ZrHE8eiok5lX/47CebS9tCYSeiuxsMLiuQXGm2uxngVW5Aa
V++9wJWeAKpRApSflg7tRnILgzIn4n9QIP8uXqt1tMoEv7AkUWrbfahZqeIIbKyA
KkxMhu3HXQD+BaJ2vfYB0mBoO8KDNFN1fykO6MchuzDYksj378hmd9T936EwmNWJ
47A4G+xpnsDPQRs3NtjywnDi9KsXcrb0M6GkR4XDjRgCs3kdeHQCQZEK1+IVBtXp
CzwtNXbVREd6LK1LejDW94P7YqKqp/eUFo/mExNe5W4m4M6stAQGEJNNylHBYkh7
0wDXXvOxunV2U7N1/wICNk/vV7iT28uMXYaa7bC/WcCqTvmXX/nU3M7gb43JnCO7
ILVU2sXliNYd13rMhGTnQ3EwRszQTqMeI//b+iLSZ9tZu+SdCTHL2YbW3+YizneB
A1skmYPlCushj3wNLjDw5ReCi+MY4TxIr0F70nwTl59oQeLlRl08+4353h/GnZsc
Jp/5FiDxlo7JMudjQ5SSDCmTfZX8HDJBuqwzCrouB8wJAK66j6be866BPSLDxLdb
C/Zzg80Ho3VthfcU40AlfSd+An5oZR5lBPNsB5Jgi/p32STgpAok0O7ZUFh/B14S
AkyEyXkVs9as1FLAaKLDWutaXzXTYoR49dywXaelhWlKi4ptjOtiUVh5CZy2e4FS
pmH2/5IPPECF1Y7MwamsSTi1/GoDOSQUXn7f/kr+C6COGEYwl0iGqva7v/RrNKzp
8zzEAV8W7JyLkcLOhYhp5rBlD5eLh3GMdUkOXs2SsUmqkr8TA0qyIpgPflYZ+Dro
m221rpyzLfDEqQSRkiBUhONWaO5GhWnx/FYkqMwfzetIkMx2IVtP4BEtyU210pQV
dz1ixtnRtRUVwgtzsGTiViXcFWwStXmdJulJQiXGRyw4i2Y5vcDeiovmP+ieuUM6
oS4ZvGZ3/Iyb6xTtRlVBvxMIszP50L+SRXTY80eJY7l3b7Yl0sAuhj7p9pihdB+e
l6LGBklHyeq2ivil40Of15UXG493BHyOup59h59ToMMwShSgrAMgg5V6irx+cK1t
9gLzYm26XkGz7VEqC4kHIwnjKZbRx3RZc9s40Yw2kefRuYBaUbJD22FDh2zqyvH0
EeoCZrOmLmhY9pHbZM3dzg1RG8KXZ73wG0SHRgg8+oqYEuY6CtWYOy7kHB1EePVU
Ziy/6dJ9+n8+M4Nx1GnFnXF8qx8fLSTX+qt77X2M0oJ/CAix2B+0ajp3qYCqWqQQ
pMZpRrnX0U+fEqwie10th61HvGY8TFTzlsRQuvoVHUOpFkbbgoC6A5uWdfNa8ceN
liyvwVhbU2Xbbsmba9evV2/Nxf44s5OiKsm+lsXsABj+H3cF8JKm1QP+kbZgmSLL
0pnyESOSlH+Wb8Ceo+GN4YDM6lb8SaRhydEYPleYHNaAiZdMXMkZ+HXkPfRn355/
/rzyvfefvkucyz+FXt8nRfkv1vJzRgCgJ6VATYq/9mF2b068vBRKomlKzZsZ4BIJ
xDpye/D4yf9etwARGmi3BRo/PZBejHfXad3YaqoD0JPcSxf1ElGLE0Gf0oQM3/3o
igRuXLF+KpbH1ebZrQvHhtFf3zEsdYyw2LxrTtUlYHi303ga6MFj3p/5iCBDg3pP
BhLtxAbiqCOQ8yWj9tZAOQJDxijDSZYPTN8h6CcSClAizpwMEjZcTDTWlx+66gvO
qd2ivENiFGBerNt4jbNqxU41ee2j/2guR0SgthPx4k8kKe7xOG0KRdgxPzF0H6D8
zOhGEFXusmXnG2t6INk73liknGrj/+rTNXduVfpXQ6sCj/p/F5jA1zvwQmK111Fz
VjatyZGoIRi6U2I5u/VyLTg6vBM3UAFvSRWhbdegwv/UT1fbHqx2HymfoE2N+FBe
+5wOSvgLMBgy+eIfrIad4O6jmMk4mVNgcUArHViFFaZyXdIb3IoPaMk8usZMyCdt
SrQQHtthf+Oe2cm5hJ/dvxpcYnzndMAwRkym9NTscKFxuNDvehi0bMyMKUG9txUe
CfnOcQPC3jeHJl+Nq6bamI/gL07W2Yu0i7Y+U2qpkDh1oFehANyQwknxMKqUDv3Z
OL+/xYg/hb6mCxfbtvhMzo4JSWG8ZPq0vrEXd21BzSV7JH6hHuOpMwOxHeUfb5H+
rM6e75n5OhISB6oIdAj1WiVWk3+Pnr4SIa9JxH/fVILrRzXn3meV4QpUPeRYT8E2
DOLjMAC8OPDjMK8wsFa4b97LIY49dgbIpFKUN5nTS0pnBagrlt5USp04v4oAHt4d
zzX7CKLjH54j7Ahn87170Ak82y/VeLj4ScxDBeOx9IQj+35gadMtdgswgHgOhtYR
p2dEY2Y/MYwSQbTE0EFTbmKIpe/FHFxRdR5HGsbCzKdkT0weNXG70lwzyHw2dcYl
X4mdY5dm8HQbIblUWOSmpvB/UnbvIqe/5zFkfqkHcGYxIUs05aGvaW6T4wHzTIZQ
GzcSeqny/BZfbNDlBZxf2idL4hO0ADvXL2LiucZtvja+KbapRVwgXnhCNsuMS00P
1347Mckf/WrNMNn8rUZyTNRQ7V4BIU7j7+BNaWXLERTPe3f9HqiW+aHXmi6sk4s3
lus/OCeZ0ins/Djl1ApVshjsfR584932thaT6qeClYqk3UrPgieKWI2JsPzrDtr7
VHykum0j5xUr2oy1q0+rWAw/8mqMVa3LuAaCiOfGKEKn+wfnRFLnh81jOGKRfzrg
AbA8zAeNThCKp+EFQgYTazsXnoCvbexvTa+wp5nRVh8QVk2N6PWaUsWEsQKH12fp
VOYqnxwS8txv7ifiJ0u31LAlZTtgvdGiaI2by09L4awd3pvqbm/Xt/ANArQ5aRZP
gKbeLllsUZTzo2zoyIphc0HXHLCnqsBjgbuaIUE+tVvDzKGD0JAuWaAu3C6Saaf8
AF2jCNiWIqZVlO7UzL6Zn3oFikfq/DpriIkZ0WBcv/tx6uH6MUjvhA0RtaJmBPAU
ZN2cdmhW3baDY5HQOQUiljZy16alEApFPU6PfB8S6Z9GDtvbDr0B4Ytswf0JQ+QP
O+7a1TKTB3vj5oo0lt9MIPArG3xXA+EoHihuXfusad7hlkeMA9Tgu0gFrLAyw+je
tlQkcLKB7gyEdPGrnkKjxqteiApEzKaOeVYkK1ZvR27FFM7A/hgmc/2TsL0qUK62
xMAYVqB8Qt9gwF1/OqsotAb0rARvWpBADNAIGox4n9vNS6EA+2LhXetz4VHmSeeI
WgE/+kXyzxF8nJDKqYNiha7M7dDNpuXOEIfkQGp5nkbOC1CMHEvQuOWZBj8ewZ9y
jnYQ0po4769wpoflMZB3v1TV5VgmrEZC6K6qGHRSqapLOD9mBRxr6H2uCbsnG1Py
9Iyj2j6qfWRS5DAOx8+kFx12onL/kaWuWznzvouqlWJAEsx79ZKdd6oQ8pk1pPWx
RlSEZe34dmaU8+XcAQCEXSdhGH/z+zpIkDw/dpzL6K5ar1I72aPRSnDU14o9jJP+
1aitDrhsrDrrrWMKyjtuJIBy4pQ7KZFinGZhCRBXrYG1BhkT93EO6LzZ2YtQOnjt
0W1lxa+6VjhHFPZ7yK0BFIGQXQ2DqSakcr4odzap3XC4tvMrBssGKWkVPZrQBjVa
XmTvvbSFvMNKAupnowAcP4DyKR3MsNInmgHMz3LDKomXaS/dMJQ4XTG1bBOWMVGC
Advj/+QlBNu+g4huIEIQTKEF9/+SoM6zcJwHAExO1mx6f3gAp6iMWWq9+erDIlQr
FDINb5btqP11f+LnPA8nKe3+wwUzucVmqmh1yeVCK42H9EopsIQ6cobLzIm61iRP
UmBk2PQDOEkDgTN3u2yIZ7rLJOmIgMwrBT6pYBVcygHNAtc8U9sTY6ShLOcAZRB3
Wil/N3JQEE43DiV+OyIMxec35piBLLAqWgx2Mtn0/IozsRF4PIuYiFkxGFZXHYy0
UIR+XQlWgV90eWi9iCvZDWvsbzvF2olX9NFaVgMsmrcjKVDXmOrSp2dhYrlkl0uO
ggW+jaoGHeBlI1e+HDsZjHCujF1JbStDMd20Preguiw5rh4CtXLrONn74RXUuDWy
71RvFrW7G7smg5eU3SrEi2Y9XabebQGCQIctxT3USdY1j2btN0ZXnWgFbYzfMy/2
wZAmhVg0wl7Y9XVjsDbVN5Unr2n62RfiUG17fQzN2ccWv5B/3KGmO/a4cb0eJzLy
dXhQDQWm5jIlthaJgtaqevxh2My1tuY6Qr8tVWO6prnXij+8LRVeb1ej4Cuu9L2p
kvtj3fE3T4Jakb+KRwpGN2M3ahP+se861N1g5sARiVvwTdkR9J1aoYDS24+SfvcR
IAp4i0R4BjPF7NeGw/X9KyTzSqWhCVxgVgP4mokLGpuuYyERAZXta8406baqkZlL
TQPzXsfkbQ6EqKwePDdVBG/A0ty8iDsAbAwp112Hqvx0HUu/Z+/zjq2LJinFNOMk
69tWFajvg1q0tKdquhvS4rTLjjMZlwQIu9IehxP4IonTkO/HXbHBeSH2Um4cMKex
4BZ1evt8CeUniH4eg0O7VOFnO4x6x1k1A6B4T3c4gtp0cKPt9SG2TbbC0HQ+C9Ea
9IcQh/85yqf1nI3wMNPAhATub2ajESVLpJlPFuTEcLqlxGL5IHBrsoM8abXBjXkD
Lnalo1+iASX7dEHK9KSF6PfNi7sN45TKcW+kW5gZD62F00PDBrM29K8H2w8PXqSA
tOOznsW8Z7Bgn5q0KJfrgdBNHu7ArVRpdwOqmBWjTSFVL1Yyz3VYJuExN3gQo0Yq
gPKTo47pW77ZzTVN6rQi68Gkyl9HUnlIeqkF4Ii/0sLlA8Ye6UU9RVRgb8Lp28I2
QA94Q2BmC/b/Yt8wJ47xxq/x4H+XNSUKq5SXUOjID9RzrmPVbFCRju0gM3J8ccVd
0omatbcjsgB/wvTx8rgt7mSwWe881nT6fnTz4Fxm9LD+9Ul77ycq076ZQT0OSa7H
llun7ngPJWmQ++7zh6DAknzzFdVkckDCIb93LGZQRV6+gScPojvMwy6Lzpd11LWh
9Ev2SG6MA2CukZ9ZKqQI0Hl65tyv+L7g8c2dCGeKmnOyLOhiyatFyF1BhZQFd+Mj
/AedW/vT6VvROiAaypDNwu6Tb5OVQiFWtRoYCzBLuT6EP5LDzlBbFK/n+9e4WYsr
CPkP+toOvTZKObfL53q/T/4TJkAifxMgBAkbFNdFoDDiWSDu+S1a1j/OuLPvYD5e
gl8eCVSHleVY42Giy361gyfB3rysD8KZouGNPqhFfCNRBfg/FpxKTlu8XvBd/LG0
LqgF8248b9ld8VFIoBwHpYGzQi4v4hSgtf+YLKCU3sD+OOXW3FwPf4L5l2dBDKHk
PRXyIRpLL1wCUUwXP5gJ1iS9Q4IVa+zcHrUh7z/RgmwLQgLB9lDiejgwOkwI0wIu
z+CSkEWqeyj1loBqQApneg+ltigWDtku2/kyqINEb1TwKYc/HVFHmsI53pq8wt4u
E/pEDPCZksb4bVoSuXsnHNVmxCPxzat0NqFLC/lKxitUHW9OKKw0NU1e7D/yzNHX
VrPu4NvOu4PUzvDsvKOfjOu1SeePNuvbTvu3R/FQ+KdStilBtqOyUhc/xe1oT0C9
xu5gDAerYao9Dj4mQkkewTMRG/StD691R6MKrgA/77cAUc/TaTtRNc58UT09dHPJ
Qngar8GstbTTRoEEW84x0xcGTKgbi1pfc3J4zAEFt6qucscRRf0LFegp/lTCsCcZ
cCSZX2M2xD7adNeLcRRpSzhYIbLRx/PVlMyQKc8fYcVMP6VDTaSa52oG2j0TlmDW
2mPWYKpRhVOBi+bPW7BtDqwCcd0aSkp9NIzQMYaR+ICEus6D08mXwELRS7rQH8/A
HKkbXk6XQtpR+qJXfNxTYK+VX3x836T1B44qfQeQMLdtjZAS4dUsHMVnJQiKxP9k
29tyvuTeUWmdUtGji8McomUjmt9KFNUaB19Ih1qGdCMMDHmgg2jEQC8AoTc+jMMl
b6f/+48SpjjVlJo5AqvRe/8ldilU5Usbp+EBl0B/alJRNpkUSI50ljt808XcK/GK
q+UYoT6EmvaUml5q7cf52BvGV0d2Vevorbpd4fKvdNcaU6vPK21N+Dd8nxKUSBlp
dsfjtRFVnZHCBD5XAuu0l2hHm38WAX/HOW85wPpLmtZ8bb9jXyCrk11pd78hY621
ICF1JS8+vcZXePKLzTXGXeYo5KJGfESVxWOziqyS3+9fBPGWMPSI+ToFx5OUb5rZ
al0HYwPeckxc/m6ZrAPplpIAQRC+Kc+Z3HBd7S/E7q0FlEvYBR0JBDi5Ywz5YUQ3
uMuA88nHTCM+XBC3z90Ud9lasCAH3j1cbMlDBGT269C4RP8utRhlIt/7nvVdH40i
eNnYCB46FZS52IMkIAeKBFKvjAIihANXqiHGtlFwhSA1QdexXoCRC1BZC0cxDFHH
s+oWHu33a1SUQp+9BD/uOaXH7l0s0tgWQZLgjTAif2k9M1usVdMBcP+YuSD/sQB3
LAxg4XwbMsv02rsLkLa/O50ahzgLsSNv2oqTG5HRHg8lfwwz4jdWliFiUZ56Ho4Y
0fRLxw4tEqLJe5eWtmUii38nmv8ho88ytIyN3Aw+j4cKewmeRxMSiTxffT8ZS89z
rmiDdhUHgTKMNwhlcUPpiZLMtObm5UUNgcIiY2rvnu58+f/Pwtd0J0YN16x1WvRI
roY09t33uM6eXwMLXidc2cSilvgzqPqbj+j/P7oJdWuQ4+7f9AHKZ0gCjUi/sWrQ
CGhrgdQvhA0Or3aBhjZojK4v/teiaereNjTv/62IQRoxEf477Jv72E30nIzOHLAK
doopH7n5qsV2kyAYMUxZw0S9FtO0vaisdvIGW3KEEjjGEHiorewvI3YZCXnThPjF
jB250/6vM/Eft9ot6v533s9oUaT0uyrJ3i8+aLlzCi/bD88o+TXFBiL7UQrgLIcg
AgPyL0m4MoNsk/Pc8FFhbXShltNgdrugABT7DK/lB7VC4jRta7jJ7SxvukjXJuJO
0i1dujuFIR1oUnHZ3tEngGfYnZK7Gi3X4YKHNoqRNWxnIhF5E8jBTyf12YvWTjEM
xtZSExwGrW+8eKjG2KlkIPKsVFj5XdGwqGUOzito6ADnivECbsR8m28mlkmfbYRS
7IhnWLin/Xksbth6fny8AWTOyZrFZJjBI9ZS1rtSupRQIXz/+PGPYnbVsu4WJMM5
vCJ9MxtYfgtJAcplIg7Uz0Oar/s0HCSD7ibFp4WUPvhUZc8MYVvTcOpW3XsKFbQl
sj5nYswX7KsNR6mzI3ibnJG9FGeleYt2VNGgPovbjPycrhdAjQai/W9G6KFXjzxZ
JfCBTD3YaeNPbjd5PSKt6IwUOtxO9ky4UBtPkZaKafPnZaHc/iIor4Vmv4vEqci4
HRVvCksc3n3ckwzgUcg0lFF5lb5u9bXS6pYmErdEibJ3evzFt4ZVQHoC/XWKJnT7
R3Dmq3hIqVSXRqiX8tKXd16GoJ9E2QNPxUuz0pODaqTHAHLayPaSXhlxr/zo9l3s
6N3yRLr9+KMRXvs3X5DLsLiNAkrRWu8usJBxBgwRpabYwfiKQJVJuLezYDerlzKh
M4+0UmAIsNB7ysIHNIl3QxpSgk5vvTbWjA8a4ECxLwdsbCwZzmcLnd0Bh4Yec+cz
i/J+g9ZeV3Q7E5VVY5vCEB3hEd3okaOQUI4oXiAV8PNpbeVg2qtYEJV9Bbog6xuR
nSIYt84cR6B29RWZKnjF1cgdHECRbtb4m7h5mAxK0eZcRKhNtXAWt2+R0fGwXYrk
e8UPQBTqg37BG6r+hnUU3kMGM0hfLbDm6AsrxcAOSmK/txAT+xkt5B+CiDpWSjcQ
f4CCTgK23STMUXCZgMW1wr9L4zxLNsaRgTjGjjrx8yVSvfYePLHdBLJu4b82Hahj
W/EEflU97ZeKJwTEO3OJkb2chKahj5adBWUSyzmxtgN6wDaPIZ42qxKdM7HQlFcJ
dEngukfaH9CId94VLp59Xj3qllbSx2lIulxIiUW21LYRk8eMy8PG7P2HvZhkiGYU
jJvcxbF+Ws3S5jQaJFyzbJ3s/7AFf8sRvrKSe+loIl75BTk3CiTpbb9plhOKEMZs
rppU5oYF3ITUFotFA4+Xmjmh2kqUs4yBaMlNTCF94xbUnTTD5lbFgXtINMNn/WtI
HseyC6sy7cOxwBw69LvY+AKNK0YDLT6V4oSbrWm8j2CzeOEH1cxE4bmgihNXdvyY
vtsl0EMQ3pkfXJHXt5+9P5AhKNat47LwyD4kYuAmNXnDUNHvvZSQ0M6IEGbCFXh1
DcQ5GZSjpVQZylFnn5ylPuZZ7OJocAv+INMWZK28vSGiEBgPPQVpKctjK09zvKIv
28LIcZH+Xsvi24I4wJhY4oS4q9coezCC5ky1+ngsOTBsYtdSvoHfW7DKrPAnbsl1
cWjmyjRVH7jqhHtdb5+dBHb3FMOaa+/KZ9jYxr1wvcU+YTbuiMj12XmoD0fCFWHP
HPCJy+tiMNBo8R1RSouV13cRsUtJJI5LdIgHgSIHlLrXnMHH+WXahucsWKLVmr/q
QvJo9qjP+2fw9CH2dK5acET5JxaEODYvZUjGgH/iDIDuF27vxQi0xfoeOGrqAkii
9bPnzIWiYDu4hqTDYnscgh7OteBPdc1KLcz/6dJCQI+0UDtxJtXAIKITuiejHCO1
zdShDfDKe0sOapgIjf6QSg7qL+NyNF9goEBSctQpJf8/wsJL2G8ZmraG2sDEummW
iBKkDtHmKb7EmWNE85V7RWQqHQ1qqafx+cB8R04NOr6d5S2PywFCRSqUhhbWrLEi
6deM97E5gkAoRmo3m1z4OFaXtYhS5o4rUu1nuwdQcXHWtZ5VHipCnoCs9KlBdz7E
YLcr4YBHJs620sZSR7wCKpyOlnJ8Aifw0pAEP3x0NBCIMJfLdH/+8jQ+PIURBaGd
9p3qE0XuRi7cyYG+rGNcVL0z9oQyoFo4ja9Rwav0/7DCS5Zt/Qq/5o8fs2AmcfQe
6mNlbsezkqFM8CTYqpELk0EYOE+sKEthOTP+ElG2sgZglo4vCoEPHuus0zFTk5Wy
Bmbs4qaA2yUm0sFpCWQ+wdBz4Hz2dhXXngUY/QgOC1RnjvYuorvg7h19pTLUdXVU
G9KeSV39M0pEqntcKXFiG+aGT9Mpy0xLpHg1K/9cF6qb66v+eiLg5p9mUY8SYjtu
wZKl5MxezVPwWNcTgkwHfj2RmiggoK5a4U/h6pcb8AYM1eGaOgBCPJejLYPPRXYQ
QPztyJJoqtjEc+PTdGfybjiX+8TkLNYP476elZ7Jt0WEl5gDk1IyWNY598j5W1cL
B2ap8hC7JW9J3DqkhVALbEO9idIEXp8tIpUipl30+r1KAQCW6QPHXsdEo7xb43WF
IVDe97cE34uRQ9G4jXUkenVDmwZyC7L+xEJckvx/8iAgOtDuw3+fpCtsCmcsOl55
fj+J2jB1bu2uzY7sEWE3pGRq9sj/d1qvHQdE3NvjOvIyOetkrVRax7P16lMw3r+A
OTs6BeM2N1lCQ2p07kw9ByMZK+Zw1SWRaBtuDs1uou2sFqkw+vmawPK6nX6SPB7B
JRn7BCAcV6mKZubqPw7DhI/G+tM8QBpPPEIgO2vmE+kP/Ywe0EXnnjBCXQph/tym
q3XhBXZoptJQiurUMtK9qzNOuMOJdNjV7cCAjWfoz7okA2vVeIwjq24EZUNzSwoC
WhFk9UtL3A/RFPb0Uwzyos5tttn2G22sfyyP6VPdFkIsR0wcgZvCpcZh52aoftvJ
BHD2qsVnVwOzkGQVE1qf2FlA/rdjwiZj+dNrispgC197BtxugQgh4d+GRMLp4Lcs
InU743KLgrdzGENWZ9ug6WLiJuhbWZqEfcvoYNVj0xEdmdozZyBtcdhDrV29YOc0
Vtnu2zFMG5Z+1RBqn+i2KzhJGIXWZfoPBnOOlI33unmJG1oWnFEq3uVvWt2Xz05S
oPDhZ0sOqQeruRbUUC/COjrHCTgv1f7QOR5Q65fDZ72F/w7D8sd1GXppm+27N/r8
o8+Cvmy8lKns1CV0cP9WvM5hXHbpk8RFt2K6ARgNR0XZFLRlL4EOsluPKIXgqY1T
m38+yBIKEOJE4pWPc/eRZWJSGAGbuRuuCIyQLj9hD5A0btVoWyaEmLq5D3ARV+S0
cjClbB3etsYdc14uAAezcKxWWqvFT1HfZxTHy68++SvXX3xg81Paft5UTc05sLYr
2E83J390j/T/ww9VbYLENng4nLW9Q+A1EkYZ/MCWV1oUGa5hvYr+ZMU5gGXkybk2
8pKFsW6SfACvmZpnM+ofS4aMLXlR5SVzAcfgmujg+uG2wuBhjNsF2fk6tXg+lWGl
eBsz4uuXc66opkJE5eM9qSosdihS3K1MX/N0aP07XgXlbpTbRb9FRGG6+W0mQTRC
96U0wpfAJs/CeOxw1yQmzOIPjOwy9CdNlNnt4KXSOkxzSCuk9LYMMRYMZloZYzBs
P0I8mku/E36fTwkYHihEzIXBU1p7wsGEH9MweW9wpF3nl0asYr4UfLb5Cm/c1ySJ
YqHMiIQCg/O+BRqwVjnAkMIipIBeU1g3R+akqD2XMRN4+EfZTowBXa/hhiamfK2r
EN41hwccQ1qUnltJBphr08oHB90xMEnv9Di+DKdUSVUNf49soUolhYoYA4024AOK
m0lz6EQBy5ML8zAAUgdWfHAJhnelfH8qjCLSA664OHuPS9uw5t6xaIaNM6O+wyHF
cfjKvxWFqhjOdPYgtJLauQqEIE9OB1UAeEizS+h/32myMOzs0sm5rQXybiIWCYQh
VRyNIIHcObvneMlNN8wZaHmu7D4fuPOeWMnpZh3Wvq0Y3QummsOcr3Ybg+SHrOo5
/hOXhn9e3dznvS0Xir+NqUvXeWALWLf9QDwrIIOFQyszkabH8KGzk8cXof3av982
+mKYg3I6gtXRcqbi9LmhFw8/w7L0gHN9zBEWoc2fxnyBQAUebjIhGdMRnt0Mz/hk
hW7Li783uoHApr199aeFylQUlkAm7tkF80B3rS3wGbsm3cif/oH1bU/uq5ZA7S5g
UtHp8zQgDw/12ggYg3QzRmgxEtpf1PRGvzYW696wLAC+nfjYezg/5XpqbG4EK/j7
VFgMqL4wWn0ta2GHVsqBCEOTCHDvAUu5iOe9sPr9myXjVilOGijgmfX/bKb2y1C4
3NNQbXqmR1FNRVgsOUwCzw2xuDtUmx5neRwiYTpngC1ZRajmeMZU+ccaKjlrF4xX
iK2TrsPsycNwC6byHA7B/T/uyl0LJFI7Mmv+/htx9gBxjsdEZJxNxogfKpiuyGFx
BFnRqHRYJmnWg/Gw3PvVfd7Oq6VLUBjUGSFJZwLJ2G+e8AyU14RgvVx70HuB5qb6
16XVqJYYNRZeIx1Jgu3CeRJhS8FZgT5tTxY/cM/PcYK1jezHNW5cO+OhIuAAMg5P
wGnAUjJcyFiVTcYnNCCbBccYQ8zXkaA+ioXA8WuFl8295YWqx3ptT880kAfAqfof
Ob+xq3mp7ldP81JY0pyi9syJIoelQQ+fBJlJ5H8kX+cNiF5dFOX8b+4bUyWTYyNF
HNOx6vCS8JVQ+2u1RqILu0P/PMxCH9AgbAHy0hFPrryCiF+WsqAlXrul2Qxm9WkO
31fVb9Tf3pjc23ARFQ+EwK4hIBeak5ktMGTIRiv3nzaZNvQvs+5nLqm5+Jcu8l9j
0+2iDmv3sKRr4hKjjFOSi3ChFJAd+kCH7HuHetsBKDAIVWQQ8RfFyfLWlqpki/cP
5KJfVMeTgeVhkrUzVpHr5MbHRzs37iIuyNldIfUIBXAk/PO4ZK/x0vrUgy2ugpKs
FrkkDxd51bmG3cyLcxpFayFRTR4IFWFy19OL92wzFPwhCEii++HGL5yVo0TlcIY+
Hvqrf0idSkN6ckJFQZ73tcb2LoqSlXm9TJuxZHlh0lTUN9H9slcqq6kJK5M04Zmw
kvyhpPIfx7BvyivYF9KMf6CCTBlDaiOlSRbBnOSg6f+INEIJqH1ZvOxQh9GLNPH+
PJEU/d7jo1TwIa0roCvV+AuQbIGU/bwjmkqjb+34gyimC+dz78BxgSFKaGSKRN65
OESqg3ypNl8ysuUwkz1PNk/0JRthKOTzNS1kMo4Y3TCV1+kADKRlWOIeI/lxrBR3
qc/lHd/+JG5c4JH2QJZ41Mis6rojXHHHHnlaVpn3UWfPtXbxtMAJUTgYJxzgoXqo
wEtXN8Ga8Mmzkudbn/VMNLfuLpJvYGwzWdPFPv8kbIzkl2G8CL5w2Z6ZOGzQV7Ly
e6tMVi+NK9iUdl6FS3/+2FVDGwCya5TkufS8tcP1ivtxonXf66DoaCh0FFRD1n17
LWKS5efWWdcWHun/kAVloFKrWAyzZBfZXO5ntW78UbktZBlXjdgr7e4AG8A4EYOH
u8lDxLhrAH+R6O1g+jchMUcqWXrt+QYEPjEAgiTGvhoIhgtkbsFNODE/FZ3MrIcS
agFbADZSbLx/1o5AsgIipYsziTT2xVa4IUWEKIKN6ij4YHvr4ZEspm6xNHxHyzN0
T60YNDIDnNI38Bg9XO5qDQwsFQdhRPYMZHIqbDUmVQvCfSTL5xj5MAJ2Lp9+UlvZ
H6PAnND4F4nQvnaj6h0RHRBcazuv6hGLRtP7AreudNCw03suKjR66BX5/Z15vPN1
sJNFkm5qBYt5KLtnRi3Ua9uIYjQka5JUACaSd4nugDTgsohLgODAWkM8kmiVSOuk
BpVspwSqVVQ2r7ePZjRTCztXFKwzV0DH5tzqXssRoDnX2q6DeWuMgYWuHZtvxy4t
c3xxnHjrypQKExBnNOVHgJBscQ8cXXgtoMbjN3lzhoeu0fA5oAKfOPaRdB7RH/1w
qwNmuFdWXhmAiJBBm5rQ7gthjMZKKlCwTemWLCWkqps5nmP5Kz3vypScIkj9bybC
9ecUriU7O3fW/NgYvWNvc2BRFcn7Q1K7PAiDUumM8cPeiDXro857KyI5CDP5Be/a
ZeTSUYRvnAjoogeyFBT/4W2ra/JQi65I3anrVoQDTTWbc/0XKCe0soWIkfQN5VjP
l524dQ8E+xwBnqec1NB5waJTSH99nxzbHSrovCU5R+1f5AvtGBpBQ+LEJzY/edE7
lqU3NEj3PUpod5WA4opmUbVtxzhO3eQGvCKyGcGrvTxnH3d2QRgcroOxbzubuF4C
uf7eDnfC6rlI3p9ldPrgq/OkY4H1ik4a9PblXQKgO6IgQKRgXg5Mc98q722HNIMV
CcvBCmr7FWv3fk27J4FKDxkafmoLaZeMuyL2jSdjCowV8puHyXne12ZPNjurEQ0f
a98wazyhpVcM4TRB8WU8mIIeovzHX0SxpPoszccU6GLZYk8QqBQzLsqKjfZ28ZGF
RRg0EPdl6wbQmBQ32YLIHbZlNlDKzaJhKmG0ssLDw9fD1UncIS4K2VQlbX8LE2fb
fL49VfxoNH/weux/qBzdY/hQL9IN4+9o+LZrCRB62cojhiVZZ/6ODKGpXd7oG0Eu
HdIGK+BMMwc7NInDyg72YqxYJmhlLFvMjqsQ8u+9zNvfF3o3Z53kR5TfyG2rS805
TQmKPholzYzf4CsCpZrl/lZZ3dxNS9cgJpC4LCMNhUoQg4RH0nZ8gD5DAGKl4yM4
lpxMXNjMLvkRQrzrVcY7CHMleYg6uOH5jy87kfxC4v8EzhsPE77EozHA3QoYwiLZ
IgbULhsGazyrfCXTlguBW1vUOXPAS5ZIwVo4E5Fi2SOXzBotGjbhuu9VBG+3pszf
L7cHb4lkJmuoKhkfUOAs+beqynKz6MxUxNuvdmjvq7x9QmFA0eHGnt7LFwegLpQ7
q/761gweunoshEaqT2ksyCfefMXgN78f0b5LZdyKns+QdyzNPLDZIDa/vN/TLibX
mL7Rdu8AvqLL7AMudEX0+zJmIwsROPwS31m81MnzrPFb+IouiH2pl+4U1Rz3OaaT
wm6M1n9BAE9B45IsI0EiS4LOSysq8EWlI1wJPWsbXK64SfVUKOmm+AX6gSMxot/8
0sg/wQkSJ+6UNEYSoOBOUVtRqHIOuE/Tku7vy6bt7iqX2I+tSYHvIyH83XOICtch
7zvaq2Kte70XZQS3b0Xo6lhCZmD0SV1VaNJobVIZqLr3//R33AzeInJ5a8t0GvIH
/UFJ2tu3LoULRcZ52IlRpcL6ptZI30YbGoUfIHx/UJjzmKGqGnBo21VheFdERuoJ
1a2khWDgDPxM9vRDmJOMeIi7DLsB3GB6+r75UOq31n/WOxai8CpVPThPZR//quIk
piUkFrBRxGtzD2JaSeOIfO3p3kaJsL49ZEcYZANEncWvdIKjJDbSEtKOh2Jt1yN5
i/z7wCYwG/fFLvr5rpXyTf1sYAWcs5EEiVpaZhlR/+y7PSNdC4MaxoU5gXB0LDC9
9UhMGr907/ez/gtyJWA04+X7yiVCOZ09tONyE61qZmVznv4gMujWqMQBwOVZCA8g
80w4Hscq5yrbiQy5tDMyC7/+XATEDoi1RpufnQpJI1BQvFh9fi/BHresAR2AjBvE
zXOmDZV4HXLBaBBAUsSv5eodggP01qptgNOByK4H7640VwNcg4kxIVKeRp98deP/
1vMHVHw5jjizAQYnJjF2t2lhdmSZBx5mIbBh6lUJBLE1SgIFodwoogCV3npSAaJb
t74UrUQCiVtAHU2OhM4c0ZdW4LS0FA46kDu/1rugtLidCDaphku7NlmihRP4JaC8
MB+93ogxRWxkccIHaUlrkJvsBJiY6vhTVpCawz6muKlOahvTidZds+WL6nFvVKZx
2csUJ6wbblNI6Qe9LO58CiLGbKnlCj4z4FXruzPB36XEP9TrXpv+tMinJXFdBHfn
wFZu11aaUfzhuTRF7lqUCJo8xQo+rZl3fpIS92rwK+zfO+8ok/gptBAy4r2KlMXC
F84C1X6qNQG4gNe3Qeq3Xe7glMQ4YJlArdMlXfCpi+XgUDx0v7Pg61pB8Duux6Tm
FnuznEjySk1tX7L1S/d7c65sQK1xz3x9M05c03fAv3gzKAcNMsQXYH3xG+16GjzN
EdC1ppHOMa92FINo955YZWDqtCeytg/YEdJhQ2yhWWqLrxiu8ufE6wBuelxgHwyV
SxAuqXTyGma8QL4bu4txth57BR/wq2nYwFa2aL3nvUascmPygeb0l5s4Y7Yl7kfj
h6jqM1+iqOCTw0UbKHv/KmVWpCrJk2TUbE5KgYRTRxJagnO1oK+IAcS6um6ktthF
PbmfvimOZP30xwg/wg4Kfk15wjQKSWJV2KevDkmjxAkvzmMR13ctFa/sKHd6zOMj
VA7USN9tUJvTvuCGmu2ibwhKerymEGqZ9c2R++mTN/+4wzcHd9bspwERDVQj3FWF
oyUmpOguJWQzSi9uAourp6x/yCseM5kMjTpHyjF63dUlCZQVJ6tvPur5Csj2N7Jr
jM6KURCoYzsUDOvl9vdgtTvQ9GcYBTgI+OyYFxJVBZM3IKLrNsCgyUIm69aG5iGo
A8t0IwCZnNvx1TRrSJIJqtSi+NBoFXsUfb0rsUofKUWNNKuqtvVaxou8mO061tab
MYR7KDeK3ySCZSQW9k+U+ed+lrDj06LHWTnFIt6WsPpE3+TsrAU6WbfjELLpjVu9
lv8OjubHD/+dGMzNE5lnzWgnH14Me1bUD+6KUkkIz+vwAb4Qp3Vt3TRCl4EzCM2o
ip3equHHgNeBrXYprJ5EMXaQBVcZFuACffc6LhcggJya/htIQ48t8YynsC7Dk6eP
MmJMwI3hGWem0BZZcbsL1n7a263TK1wKRwcauqfT4DfDIcjzkB/d96P2dphxxQfb
gU1rHfUT/7VWj+wXhIq0ndelhNtPo5KSPOLh9fuZf+cqPnwYNgd42N29WmZptxq1
OO4KAPok0M2rLRvwP/egnbUwPpsPnk6kpNvV48rqglu6kxxFI07wb1BocWn4ZCvG
FoCjnMtGLDg6wTF6JpJVqVGxg5XGQhSjesuznaIqGK4LU8ybJlX7bDj0yuk1v/If
Z32bFCLGCnRn7iP+4MMwkpo4uivCieb7id9zgDrIkm1R78HCs3uf52XNSER9b6am
IeClbtcfarMEp8YNvx5I3meeAsW2tfHyJODCCoq0u7lbF93ly5YQcgQB5yXpNRDg
3LPkcyNyLdoD+NrE+Kjr5IJEwZBYIPC1XJAZ0v6VKVrjJvqmTZVL6DeRubh8lMTz
/+hbcd6OAy67q6abyKnNuTQTvtC1k87Q1iSJoNyFA1KKmkc9F/fJWrRw3C4F4sqz
K4Vn+iBEvExmUsthIpOHRhcRIGpzxIguzqQurItZpPTRj1hBv6wj/rKT9CbbxlpJ
SZgUJRZp4SvbOFo/CD9oYVTKErRr40VozMxv1edoyxspuuLidwYOVDE0fmwYgCys
DypJxBnR+gTeE7vSuHHgBYVFibqOpjB5XTJjAwR8tyB2x1GOfQr7UOOO169S29jj
gH4j8aj+UPyd8USt+ybf0JU0DgvH8LCwv+sPT9jBVmvmqgkj/9FzZNCAmGxYvCjP
iqj+pmk4cUcF0Veg6MAQoZkj9IgF5AcCeydcsb0ZDXZ5OEZ/nPSbRYWYjE9zZLDi
yLF7W1bFgSgHpOwEs+et1xmhqzckVfLTYpZFS/IYJY1sZzXJ4Hh4KcaStJIctpFh
x8ZwaWulnEZfD4nsjsbkOYy1ptA9t7hB342xrQvFemyHQxmlRx7H3IMxFyPjhlIQ
R8A8SCeT5XwwIum4Tt//gFgjzQjkZUfmuzQkGXqz89JUmM5dtdtuk4P9b528EFMv
tmoVwV3nIf7fYdOIBaT5Ns+S7t3/CHlSHMGlnw7pwdK3Lxb5qvF8sbTonG0G9YmY
hDIQ94AFMN9XeFmuWN+ibrIzVDbPTagDiTdl9YwSlAjYudXJQ6ZSkNIdzX7OLYOv
0+DvQuUxPrnHVIvTmVRBACSYQx9DRLimhI5po8//K+RebyUqChbTwKu8sMUPrfXO
imCAd3iSwS8ZfRE8CHXgHy9lY1OYp2OiJw+b1OAp5ZvzzVOxlzbBmDaffAXLhxq2
T6bKmVb8D3Ld37vbTgvwdUyJ19uOEPdC5v4dAUI7MeqbJPj5AUiL/uXRLml0CX5o
/jirR5T6OPJtbbwZaMlgMVCZqLy8WmX1DIrufqCcFReJP/u+lDKmQEFANABROTMU
pVOQ1A+B6PHuEUh21V4QNAPcmCQMT3tqfhC+Nm10imW2s99jlUeqkyfwmS5RHaE7
TT1gR8XMgZRFV8z6meyQdtMAnU/TeoDsuoZwgRZj4AJ7CLGjCge47fIlCy2Zic/6
PGvYiBPjUCsIEMtVsqf0Xuhcb1S1QONfy0l/APTWoXt9gee6MpL7Er1KrIZl3to5
CZDoBceo1jgtg/a5+spTYCYW+vnd7UPB3vOVUg9BZJwd39PNo6VP1+uk+tauMkwZ
WMuNmCohTDx5b1Wi2qNIQUlBeKCTNGbV8QPcVZxFVczWyNZMMTt8GVDwzufI0Gs9
lcj6E+FAiVJ+xF3RgV+jvQ1k6lN7u+vdFAIXxnBFWEmsPDW2NrarG9ACy1VGjFE1
DGG3/7FgPLcwLHW95o4tZqXG+g5b89DdNwxkZHX5oteyGacabyG7UAVXigFROCjh
SLf/qB5DvoWT/rS51+W7zgwcag+6R46HMWp0Bdk8dbaaN9BW9ShHPn+P/19q5cNz
XJ5VdE6Zo98f4scSIPpuibAAuvO7NC08Si9qFGkKZLI/OKof06MrxRWVHHsMzmZr
zetYWIiBIynRkRfIwCUpw7L5cDn8WA7r3JQxf9TnCNcI5ZZ5AgWKZ2u5CWDZqXtC
UDAZDeBWzakiz8f2W7LcZxSt5itgU36irpwsVrBxocJCUJXALzdH/tA2t2zR+vID
JDqXItyhatMVPJVtIsRYTU6FTryoUPLgWQn1pnRTfrzRdZwP3dFuBBkDxKO1iyaC
8bcvB1Iky+64MbNk6cU0fTVGit2jydLGH54jfnGno2v2QsTWnWheWqbAQrM02dLq
Ny7g+cA0mUTzo549tzJaPyFgFjOqn999xK8vp8IfHnVp+xIKe5eU60aMn22QBpX3
tMUFck/PVlBOt53fwaXQcijh2npU8Sh2U9lFVhqOPGqkWhyLcvkU1B027hziDt1A
ZwbYFywZRHUpS/tD78nwe5Fx4HLLNt6j0hqjPreLl94xkcUo8tJCkZCEb9O4/CFr
SHIUi993q63gHZn53Vs/JZoiYs/XRDyCzepQhFeGXV/lczDfFSlsETWzYiPplvWE
6AvafTN3j3/+duheFr7iii68AUOcYinCVJO3lUFG4zouQ6yja0kvjAFGJS/v6sBx
uZaG7dODy1cTEeAncRYwnqG6+6pNtSdIfufUjHVKXHdoLFjX4Oir57cbL9hv9X3s
3G+B256gcqDUFqIZ7JNrWquU54q3PZvm7K2pbDqVQGdFP1dF/J19pUXrZjJ+2e6L
JdgIRVFx3PCtY1TN87FdVSSH2OvnPJZgIJrNFEKDPV/KeErAdhDHzFYBmhvSQL9l
Ol6sCFibxLRzcFoKhLyfk7cZN8UdmbXFjb5HM9v88EmoDX3zxYJ6JxVdiT570744
PNK31sIV55xLiTJI86kWbalz8Ef+U6qtWZiA+TD9LMPLQZKLGcsqhghjnGwD1zcS
K1Wk8TpExewlanlPRTiCt8zayMNJUA4tk8QT7s6Rh1+7OXzn8ZowuyGQ8b0JdN+x
WUjhI3N1s8w4/r7PAAFZ9wXOnvDXYk1JSFNbd9txzB0NtWRRQhZ9rWUoTrJMfgEa
OEoGHLgGpq4nMD7gkv3zzqs3WoZQQ90dNhAeS5jZHc4UkUMH9zsMeup/kYzhUAc1
qHXpjMqmHyJwfPDBxjIvfZjJ6/JaF+R90Dp9QLlOBGk8QWqDogOi6yszAMzY38Pj
iZ0Lqy1uzPMtrNjgIB2NNSPhImYbGYI69t3/LbS7lQQAJbp7LfVgoG+/rXTBvhx7
WkgpjvIouk/NC28Ce5pxBsm78Y3UXdmmEwZI4LbD+c1tTyWWiMmv1Q6a3+q3IOZG
ooYLOwjwBGhXFYbZqbc1wu6goa8TXxoMIQabMiIRTPd0fNTgN4AphuvTggUlkSNL
EfHIU3m3A/0EXSFhhqICwuS9TxJBrwK0iAN5Ilc3RgWXHDJNjeeNkR4mZD9l9MNp
5DT6KAFsNpZaf8IJXXe1hVXIn3oU2Q3fSf6da7Vkj/IVpQdSihvwtzPuMcpkkAVb
HBG8g/kv/BzD75zTZgxT6u9aMHgr5r1WyQ+k6BNXUh0Q1k0bgPuky5dWVlL2lqzU
95GFfL06jwCM8zeJAeb6PJMbLFA0I/a2CPQjvtzE41lxkyj3B+R5KVSquwz7WtN6
K+xydH5hIxFhbSWT6p6Y7adEe2ocTPKQEhV0dVWZiJDOesat/Vx9Tn+UZ749tYAC
Uis7VhPfabnDWYfwGEs0UX68nNCkyZ0sXNTqFjzd5QG7EJc0pdAuFLDI7cAKng7i
16qUV/YYKUVEe5ztdJer3K7AQmGoviWkqzqLk/ywsHI8tgoz3ebnOachdS09DALn
PSXPU7bxAB73MN2JUqF4HGsZ/6OxIL0GTLhQuzl/NqOVioukdLZbqV0lHIVB2aj1
+98WliBhWxKUCrAMnxraMO0wyu2gZiP2kFj2kX2ICwaVqwPTqxSh3Ll9dQFQK3hz
DwCe+pbfjPjJ2obPZkezr70Tt043VbglQs8zwusG90Gbh3nZIl3fnoBj8Wp1nwCQ
oSUEL6o5WDkBIUyhpXyUa4DcqoUYo8oULXC9WBwj2tBmCLObW8fdUbRDyALEtDSJ
NO+PJhPvVzT7ZCq/ofmynaHJ55IqOHfXFGu2zyS3I/OSwI7rpVHDlLiuR/xit+RZ
AoRurOeFAio8Z1ESzFtx8pQIuGJMGQkY3QWUVr7B+5vV9LMGsVlqpxQr2fWSUA8a
L0kBNHCNBfxfpCpjeYIXAf+9yGKlHHtoAk6xAJFt1nHnSG6oKlewQANKZKpfplfs
/BHlRjOd7bfbw+l9kLzP3mTWtQqVg1/XqVY11NZI9cQkMIogZ/6hyLQ3LkFwuh0w
mMJgU45oLVvijMHVR1gPCPBCq1pqyIsnvZv/pKpvfq9fKmNU7K/Mk2JF+JtJ2j0R
me10y6czzr4Cr2HLoS8GfuDxmUwFFA9wyYTz/F2UAwAR/aqXswx4rOKfU6Oghhcs
PBVXk+0Ym37aXblkOYz+glAHgesrmJP0bHBK4mzy4qbmIEZYzWpbmv7TznZYYuyo
ewZFz1ZwjDR69TR7QG0oUzTx8dMBMOo55mkobajpfhqjv5k9EneIJ4RBbWBrRGXH
xn4/+rNBwSFatkGC//4Mrt1Plxg6Q9Rj1owYU2HeQTla0NuGqMsJQ+coctFt7+8L
IqRLZ9H7HrE2kUDuD1Dly1yBq9TazBpjRmQhKhPO+O1Bf3Wi2dSMASf3lD9X64oE
IFErdO5LzXeSOC4n/+GZ4cJODkeIZPxg8p3PKFK3PLuKS5EmBFyB/IzqfWwM9Fvk
r7gtNDH1tsnUm2VyQyza6iqycOl/IgTKRxkJAYNM/AdL82PGa22d9gHveX/MvivK
7BfsHcXX+q3YhqhzXVv9JvjbSUnMCw6/v0dg6bBs+L/ksJHiS9pexN1aaZcD+aGj
ZGBGLX5XqIrGoY3zQRD8VzRt1pr4Fzn6uPIQNcYVUJUfode29NavzaJZX/fKVL7q
G23PlrKMXJ+abeJC8H/M5bKacXr5GZ6nzmmLu5RtQfNYBE8ZeIdPc5x3H2B/ziSW
sWz2pnq7xwW+LUgtpLptPGNeYSJSQclrI+CRto3594Y9QqRo7U9J0PiHKoqdYt06
zQ7uWnwZ8I7UsujrbmYuBL+NAYgxut4ZY3UboKxfcb+LZPVKrC5CSCCCl1Syagpw
+shGPZPZTcQhAF4fP949NWL9j3yHGhWxX99ScW3FB249qqdZJjr2ov5yr9tOZdbf
NBU7LbffNHKZIKMaINMOzC8tluObgZRGUOxDk++BftZYFs+r1gzDmDJwBXdc0Po4
XrA2h56haPIkbsFuH0YRJkKoMks/8Vx+Meoa3Q92dPfrtWeI/RNMbtdB1K6F1RFA
MvAEWTwkowBRp7fex+SPGiqC5IkGdq98acPNwFn/X5hnAwt5253OsnZP6nDZ79Vy
pbjbLOl5Iwgw0olbMLvd3hpuQ16bp2JBlIRqpC/GJOX3NicRFHE0a+FkS172P3e3
LKKMeuRGaiB24XC+DIbREDsiFtdW5V94lyY50Bg0bCd8d7os/kqOq468Zhe8rcF1
i0EZBb2OWcEaaxb/GHrQGgbKAN2RwbmluA6XmdApJViPyudibwRJu00nSgxFfDpM
c2LwVHHNyJ3z83AHTlqvTbIG1PvRIcRq2YtDojINj1pg3nNdVH+NwE6k+pHqfule
SFWeqAPT96bArCq3QT2RVV20q0CdntaKGBeYkMSJiarBnF9jlYebsqOjv3c3rYjw
Rtnka/yQWJtdnU8aDGlz/6WJkesvcFn8ooOe6aWHn6faenO+akeVJxaCrVcMJEu0
WVp2lPokcOBzFoy4v5xTTagMBdnjG7mI3HXFMSPOtzIeiFDiDtad8BOcjMcJqWJJ
9KqkZQDCsn930CwVWnF43yOKNdRTniXU3czR91lClt7UfENR26p3W+YU0ineov2T
uuMWL9ltzebT6Gnh85wTwp8gVuo1PfbZFj3a4A6+id96LK/H/GXgC20f1HOwQ98m
wia75e33lnRCjpqq0ekUU8VdfScr/j2Fec7w3WRU0jgodA179AYStLu31QiHpc3t
XAlOvy/g0qfnWxjUl76lQRYqQ1KXvAnnj1QtAX8pPOB34oCVtQyfiJFJyau5Ta3a
0kJPG4N6+7cFF6xogS+YtU75624BzDa9Sq7ggg5VketmaDj36VIybAGo2PBYOgD/
GmtV0u4OsIUxyMjMZOEyP6sk4Ovm5nYTxfWlZVFzyLndvO/W5q18B6gYkIaRC26k
6KSwkutmOvwDRcigg22fJPf8YRhmMfvuQBHGNykKHAhIk+XxkOvZNR3Tumyt7x9f
6dZfC7JVCkHlXFo3RHEStCLS/03YgRXOfNNEvw5QNalL/fkxhW5I5FY68HaGvWqz
hnqdjSMeDk+6DcyjYsnc13ZAdwW3egPpiYO1oLY3RJHPRT73XHPe8Gx571usRjoe
ng48cslLM8QMBMqjLrT3uledt3/RtghAe8fWrLecj+9o6caNYqek2S7kDWrUDqaW
aSHTf+rVZ6mUoNM3bA8BmMbGSRStxXJZdaAkGaMUJj7lw3cuR4D0+hf8N3r22AU6
btnnyO3PK3Tqqs+t+CPTTVqC7p82ZXeyCGgOuaXmjK3RU9ba0TjgCQlOou2zwDxq
mM98Cz2KdllPWwNZCc1Rxg57jTF2AT0ukh544aXZpTjdVHEyXNnWQpEQniLFyKwg
wZyEpRvVYjOz+3p8YrbgKoTsJhqVHC1ndqO3KapfZ3kIcBuTT0ZPVRRh+fY3rUma
c0uvkMIWHLf1sPMSzfFVsrfT5xxfjCtw7BHf0X0MQ17TVz43n9OSoLDYKAY0Qxvr
OkfQSbkXIfLa18AufEXo42lQEuKZTfaNzRRnvdw0uSuk1K2UCmBck6E1Is53oqjw
TIkw5xxg/U8nZF8W1S4MMTAG1BxNtBiLbtWdaqhYHSmEmIKuLadqS0jNP6zNR3eO
kFLnkYcriJ45WT8QbFX940yvQ6REjVR/hZm6eltnueeG4xxFeagRNO0bPzve7nzQ
O8+gDYxnB54XirzvMdzFn2yMKGjdgM/n5mIs7VHbnlf8ntxMTomtGtQwjemVX37S
sSsojTAFyNWqLew9xTEuC3UWZdrLQHGNPNj+aS0O1F+qz/NWpAKapLPjdUDdmIaz
9N3SYNlkpFR4mZbzC2s209rGYyvRi2tqzYOcTEctBhF3mKrinu8nMDPOMimDdwRW
2awMpcZ0+mKus0OQvEPi6Y8q2lIkj/XdW4Eo0vTs0/+4S9dxZOpCOzu+Akl3LZss
RkWL7/nZBAUmF2IRnlgozRztGNgz2F1+XjYhDp65dfzf15B5eBHbDhyPstYnO4yZ
iB9wCB5aeRVdPCOhaC4b/gbn/g5snvMfg5ynrwATqf382wA4C+dpFI6SlSS3fUHW
u2r15+H6zR+VsgfGobdM5nPcXB29CI3G6KnAciOETcvJythgqahSn+O/Z16qe2k4
3uGnb2SuFgSGfXhusld+u7z292xOtx5r9QTufLjD3GgBahKm4Ng9myW5WnrvpJA9
rOhZXmNiD/oZYDGKHb8awpovrd//t5fa1iklF4YzeeZsgFfvj4hz7Ei6f8CWMh86
WGRRZh0becFr99m41a+DoEeW9eV6H9uBr5M6fxUbzOSdpFoNOSSkIznvQ7lYJEp7
v6kEtQbdp839dPxhPLWveuO21AiyHFPe3w10tbcwRAnBNok3pOfPOyaEi7sao6Gz
e1+Z+hxqQ1UFOm+xXtpOWflqcZk7BcKYNJc8WuEyQZBZl7EBM1kaAmtcV7aY49WQ
baHdMKAaGUU9uFObVNIZDj90ifYrd36/cFco68YGU1DSxq2fd0FDBhNt5ta6YnLg
TS96HaNf5XIPSPBctNy6H2nYh0+ht1PqoEH/GcMWG0Xm/LANpVv9x8Gw8sxXkzhR
t05vSkfmn0ZBcHBBxDMODjWkWDoO+OvXfa4Wy3C3p/VaTU5WXJ7TV1ChTu5vxy0Q
Df6PFZR9aebauTJCiWRhWgBMZYncH72DgkFHiC36j9U0strFenf8OvHYmA0GWHgT
mDEQdPHbhGX+y2riE406TRaOgy5EUBFJslBkN2GPZmcJeY61cBeOwPEapEcxxc2H
VO+vwjO9jGsk76yDmGdG7JmVmtpxe0csFg2Mp28EYjLOtmcs+rZkXp0jPL86GxZ1
cgpqs9PS+uce0h4Q+7mDt2CH3bsGAlT5y07adaz0WZu16OeKbH4dvB5QJMkfE7Eg
2mfYlzKOepMVc2hhYB+qjOI7WHyc8z99K4uemc6xGkwJxkLgJPkLiBS+Xftbz2Sl
xdiyWjw6uka9LsK4cGlRM9aW7iITlOd6uLOnZ2oFn1PuFuVmJG0kVfXSAm0OIQij
2TTWpKsTUu6QBo7gb6MwNS8WrhWVTWzG0i6lj0o0joPLldQLuUZOehE75I43Qza2
aDznuFYg+20WvtCi7LUyN1OhjHhGBxIr874+VYFJRrY5ptgAXirMccsePTRX86nB
Xe7+ErfdqAJH9DtKc75Hjd8bXcjDUwZmdG0k6iJU1EJf0HZZpKD3LAQIl1C4xFfv
NxUyPITDBKrT0/rLvIyoC3mE+ZU2arUX5G300Mf4f1TRet8IQjM19ngPwIrLbu1K
Hj7N/6rxRB+Kb7iWW+bxJ1OADFds+Rzh4c6cqP/ZV3IrzvkYKxxZE1r4KPE7k1lQ
9msXdTxCJi3iTuG4bMB65BmpZvw3bFluz5nCr51BRXR4aOCUdS+wHDjGztwSZHyk
hp9AkKWn+5zg38g7jsK/2MkdIAqeNzlTnPJpMxQ4mEtm9YeRoDeiAKEaJdVf2Uwu
XBHGc2xnTWHPxpNdesUN5qBgtO1tFcFHrJIzbgDKeEZM+MtHZBMz7EpgwrPiURPg
+h0PPP0lJuEMFob3/mQ977I9v5VsBf7ZBe7JKrnJaUKHyHEefXrlvcciGYsqAf9J
NwutRvQsAzrdV9MJyFdUcm0jGeU0cE5gEvS7w76ZrMjLLuceX/fFvgeCIFESyADO
9+wcNu0QzbCN/ne0ourHolIkDVwtQ3GqU43uLzbzLFCFOpLumkraUgbp0v2ynMEs
Xj35Pc5SdtxgTk0RlEi2LQlDLgfMd38XODDHsfIEflOsLoxrJkaL1I9CAiyU3v8m
j8YKy1KPL+kkpRsGn9nKlmuKvPlYTp8n1pV/9usPGyFc7j1uZjg+runiniZKPzPu
cmvxdx41K+OvhljFy7XKb/yxK28z9eQwif+hHKwQN69v/BGGqC4s+avwjBykhN2s
PwugYzcgcwIxINFMgFVl4O6rhmqpu+BdLRh3IR4CaZV4/piwYKB2thQ5GzuPQ+xn
9G61e5z9sW4pNoFP+oGLqhoMKcEFeXnZIXGMJsmHw7mavsrP8D+RgMf/yVq1vlmU
wJ0leI1IrL4fb3XetHjPg/IFQdHI0oohN79zZYFgVmW/m1hzxl4JC0OoS0M7e8Tt
DB808SPRfDUo4EUoRQoq95A8c7YrN13BKZsF5aighlF9aCtEEGHPdCGDfZQS+BKG
6+3+FqaDieHCo7M0eTvQ0C9oiCjYuhOkhLqFZ21XcZXPyRQpLXZjTE/gmDOVy7MS
aHhUNL8F1uRei3zmtZ4l0yzBmomP38MGo4GxNcIyEeMCKaeZgvr9cDrlN/UGLsE0
gsU9rcRiibN+b5P3DWHxBVzgEi6g/N1kol3hxeItr8a3LtkD5dP54nI+RA9agzdv
qi5/qoW5/NHwWjrrKjOpa0w5bkhMj5alEYHEZ1Syn4nJpCtYvC1JBvl6tP6TcbTa
KRK4vVd8UX/RgEQoOtEcEky3T8V8QR0l1aa59n4fjNOxH8XHFW/vI8XFfoGpLPC2
2qgQZmZHGO0hmQhDYT2uGaZna/hn8vJ/uacBaIEFD26B9ypy571EWw+XurWeDy0w
Fu6BPhHq/4QcYQBUE6TaWfCz/mRCeAsQhSY39iz0zmdmzkzpuoph7Hjg8Qelthl0
DJtPYHS5G2RZ9zzM4NgEHI0MUPZfRxv9TxwMjaF747q8KGSRmoQc+S/x6OdJoNG4
i1jn40yUdRMubqWGD8hlMN+fBPKxyLpnZlKD5xdQZB+CfYjJQ+glBJCV4MtuMQe9
9YxU73DscZbjD3Y6VHz3y0yWe7Uur46BcD70izkZC8ghrzsq4Ms8tBNUcfV1EiZY
QLfmF2bCb/FapLJY/AgD6LlTL5KVvkKpstIN0kOhORbCa5sI6uuoU9OZTXCKWlNM
bFQY/itxHSW45CIegfQblImu9Mstebq3A3nOXcZCf0x+LXWFXAQ9qeF0Cdz0emHK
AJFGilsQBIF3832WcFkANk54NiGLOvH+rQkcKblhSapasEQ0Sgf/D5jx8xVeatn8
tFYh/RgYZ8gG2ZUYHBIn0Y2QvE62PtnJtmExHdcY7QOe3mY7L1fO1cXKtcMNX8Ud
J/g7iG36jcDmDFTuYMhw3ikLF9mF+O04wCg5y23GnVIHWRbvmekX6KjxSCKwA7x+
2H4uT+BYAKq8KiYNt9MtonmsRA3tGvxgHeEjzQF50aJtjK52Do0/Ko0YgwLX+3Yu
UXjY6LLlfdwPdH2hFgYraEfoxSNgPwc8J4ptBsI+7yOdiWlCuUqtl67MPHpo7caS
Kzwx2IyodpP783VdDwXZx7QYnIMwu/sKL80hwWPG6CFUK2v0j8aUE8ZFN+FkP81z
0/6T+bl/rP5q+r9SbNzoSV2C2IGT20yZ1a3Cy/GXTLu3CN/NYliGRgFgsfkp9OEZ
axbRPUqbqczmYaGwShJKxTgciK/CMcxS5aO8ReiZU83DEWi7Shhvg+aAigMV7ozY
nzky6qvgxwriGY8iCpwa0M+qerRsJYx5NMh/l7/tXG5ycV0+lI7WZGqvkTA5t2v3
9VSnMS8UtPkqZVUMf3bpb2c0ao2PYNl+f49Y6vmkSExwYTzJuFXlOZST3k+swKiX
htkKa65Wk2jY6FFf5cGONJnmDKzuBq9Ca9Va1Y3qI0EkpCNgHdrJEjwg09egCy+p
FoOrXz5TnGDW8QjLmD2l/hemXZZcftBTVE+YUUU0e2V44tkP2vXQMlfUmA880yIU
Pm4nMhCX8WcZJo3KqhzPbVdnX89csFHJNdE5I4zPXpW+CWi0M3RF+SteJI/HTPBh
Qds4H6dGH7SihkBjOxsCmLt9RBKPLf7sCyoAYAxOmRuUE9A517/NwvVNLNWf7bel
znBp+eGnIN4w8bNbd0CXSprI0e94fyCDemsYm7lSa9ajkEpSNSBvGMRRVLSau6s6
UmkfbWiJmYmgwcfmY07LLSfUTK6CnySykLr9t3+ClxsnKRA9nF7JKeIDP1Y56IX1
lvB5q9iEJOYC4TFNvyRMk0/43EiymQcIOykcOtdbgq9WFlhChTGfOkcOp2qZmtnL
wdWGG2C8Mtyw2jiHNZCvCqXBsIsTVqcaI8JogQRYBrKfymv1FMxS/ZhvjZiv+DHI
bUIkqU8YviEhsJnHtn+X5eH9hMj8rOGKdGE68/3W15wEVt5pTKtEvV65zbnMn1ZO
f54MutDLcfWlFsUR4irJpsUd4yuPXRP8vdRgiIyLIxvVPvJvHlkhBRxP6u0og7hJ
vBEEQ8sY2tMyBRLOj5KTvbK7cNikenzFa0C1Tvl4PxQXgZIVsiMGxSWUumF154h/
DOGwGic/4uWHReH0i/dV8jl09PU/oj1bihoxQhKHQ+SyphaYZoGfrae8ePrTYIv0
Rl+ToLVJ6TrcRoAwpa9QiNLwUU6ngikoW9HL+9D8FRU0GdnSJQP93yjeJFDE7P1w
yhCxbI8/o6FyLKFDhycK4ddoY46Q8deS8t/Xp3zFCXd5cDJp92/q5DrceeM6hULf
unDi/2QTWfds6ykAb8OTU8hz996EBC4+DzrnQ1GgU49Lt77YmNyQRfqxh3Qu8VKB
JNZlIYQCFNyDgrbZ2ShJQ8H3v0+2AfX/wxa+FpKy4bhxR64pXaWIs+sMN7WaOGQa
P+KyMIXpcmL5gwUgphNL41jO1aHXGTm92GWVUntEvaYYnaKbbjm+TZ0gTZLEukGd
XBB8m9LBXfGn8aGZri3Df0UKJtLHstjZctL+ysGr5DAu6t/oueSapZuF+IFt3Ysx
IZ2VaPgalv04gPLvyZqJ/cu38Em8OJAOseT5nEkN2f6piPhh8BVaYhQo5GRmXaoC
2WWHBctQWHYUIJAWM1HVkB3Ptey1bEOLFfOa1qUxfukW/5uAFF/o4ksZ39hUlMcP
dcnRh6Fixis2Lb/jSAdvf1mWMQQbMQsHOAYayI5+IoC+F7j8fjEpAevhqN74Q2AI
JBOcO54/7UM0z8H9mvHmU6UZhJlN9D3WeGqcDVs7utgcEPdRpc3P5mzAQWRS271l
YNfaQS+UQH7l8T0VNre9ReHZ2EfdqfbvHsTQcSrqM3/FuTHUjnB1QCajRJgUUD7J
wCsYCQbwvKpY3KqaqW/9g3lexIZPzg2JR15GpKvZwgwKwWyOmCH61cfbAUPO1wV7
30WrFSA2/EUuuTKEQNfKPnnoin2A6noTgqIdWie8+OSxGHMXP3pUmtrF+MbX4jQs
OglaSwGIRozyGGz51K3f4ir8OHb3j4tAFhOm2D0iLCXryTIB7eEb2qNtnlXVKscg
6etCHZKerDg+WnxgDjiSat7hxLk249FoMj6hMrKjIIoMemLZVSsE7UK52JEx+PEb
GG2ztvThv7LUyfC+7M+w33HiygU+52MvwziSvsgn8fTCB+AWh+pRdnKQZKb4ww2g
FmoGMg+DLIw4mlEKHE0UOqfU4n7fd9GLATs2CH8XBbkL4NIh3vFgea449QFu0i1f
iyZLEDnfehpuSnjQl804okrLLFukZAX8YRSF8KqGSK8Amb/mG06pIYlRo2uqDvCA
hNx9MDNSzA24e6EEzizeXO0oCZcEFWG5MgyNVLwWcsOhFQ/rtS8bMCVo1k6diier
se4fm2QTpefwtdJ99ajIzCN/a2aHdfVlv/VTrUeZVM+t9nAVA1ie5sdi4D4807a4
JAQO2NMrxy2bJXVczCvs1huQfR4Ndkf6eUtjg/n5nuDGkBjPE88uXSGE/vUbuPt9
cnET6TWFxkmVGSHIGdywbJy5UH0rVdQ+c50HARqw/yBWbothdP9fyPOWRXnCazKF
PnskPJCEerBKGA417IVeTqkepaCWI0Jpr9YLi93qLvIwlmjQrmSFPYFZqexTl9vl
MGrKDfh4E6GPwEPW1/4BCHGEkZPk/W+sVyvD4VgVuVFpPkLw5IfREfnenrF9sFzG
uOMPXBqH09nJjbGD0rGmVSaVVrrT6DAVPti0/zJlIbb9nUImTj7VEp8SfC19DY5B
VUv+wn68h9X9RaNj++R/sawONVEHS5a2DwD1ykf7L8LyriS4Lm6vs2qAlZxUwpEw
ikErdurOfTVgZ0TZL7d06RkFtQnOMtrjz6Z0wBwUId9oOs9Mc1BREeGz9GTsS0ef
SSliYnH8fsaVafZZv9Mp3WPjTWLy7KjlMk5H4Sl8xWbt/8CvtY7ckMB/T3GCB3Zi
Cc+5VYPy//H6ZNWWHndfz52/1HTYZoi/saw0EvEFuSWY1odejW9oQ21Tk5ZKNJgh
TscqGfFrBvwLEK6KHNj7YbXO+DkOlG2QkxuXrQRDBKh7cwQSwJv+Wbbrdqg2Pzsn
J78klKpcyGnsIUObi9sRpKSd306DUoMVPXWBp6LJAOzQOIUEW8ytd0pq1/l0OC08
AMPqjxaHEisrMGf0kdw/W0sYYpxqy+2u8d0bysTWIDKyJ1LHDeZFmwvEWucMBaKs
v58qIueWFeu2aZutD96QuI5vriGPC2PuZ6oTlsjfBhJ5sg6k3YyaDjmLgo+RTW/k
xynzpnGGi9ywShwmtrCYdNH3X/Mxfh61sHWTWIYGbndoA2X6pmrLg2IAYvZ0CL+I
1PkezDgadFjkwboueZBx7x0sIpLUbsqDaJXPOPEQFZ6eNljL3Q+1yDxDYl0USfQj
ptmZ22ZLx2wFLK6hTmVDXognVoHrXKPb6B2Jw0lkK8QZKe+2N2/2opiZg2KVIpE+
eQsLIsqN75UTEweQ12VS/PXMoqRL9jhPYlHF/GkIZ3BDfvspcrQW9ldGFVXTH2UO
klKwz762+0tbA7z3vS0AEh+893aQ6Xv/hh4QR2E/D4/DSKUakzrcUzMDdN8iVSMX
EP2Uq6uSYMAbXlvlMNAdjJ6IKht63RmlIzFSYHgjoYjRPbrZApkbKzfNSmDru3sc
LYoaP7Bo3vMoXcIvc4BIzxqL/CUhBJR4dDW4MCxHfrQ1IFL6xUSnCnGjdGLwfgex
3GPpi9zehv2G9w9GECH5e78wX8OwLFg+Ow66sj7LRYXhu5wlSMOuKpTpkCqergJp
g/vSPn87LnkMrcCy06rLgewVYzreZ09CWENE39U/7EYjTRbvRRCQ1tsgu0xzcjtv
70uKJKDbaqSKva/UEiM/+EFVtTNBLmymE2FLOtJzojVSh5X48NuR5GvZm4Xq7Tsh
4SJi+GE0Kgh0nFk7nTSn9p216Cx5D0iW5e387p+b4MKW+hyWJfZQopyamK0+/MG5
06iVoOzyEJEnZ1mLK9wu3N+GJjjcwEPhPMvvAysqNC6YraKTaEwqQTPm0d6KP64w
bRgTDxcBwUJf2uMiO2WRgU3q0odq/x3iE3jeBoXuEJIMjVIAe9WZ2JhGDkFh9RUX
E7+bxp768J8dY2Xjz3ef+R8v7m0ArRDnxcRg0WUJkLGM8XZN1AVwVRJpCVvUl+5V
NMqqMMcv3Ivth4DPhEyb88BbFVsDX/zkLDGBpSwdoEWXhhYpSBmgdg7b0J0aW9pP
JmLUzvMpbH3L+7eFrE0rPhl25zfCUV2I/29rUTmK1pvWRCNL9qfWJiy6rpf7l6aT
1vsZpCxTv6XvM57C5zEmmXM3FFllPBj1BoITMpyKmvF2FlU89OicyK0QHJNFuZdw
J2ISpn0p/JrBo3KxZ4N5CfywpeY3tm+llAJNxfmmenlNBdXtQvihQRlfrEhiqKhS
OOOF5a3nX48AFeh5hu4W7s4jJOHfU1RtUMZQw2kJv/BkES0IbdwwmK+8UUdkBR3/
jwDSf+M+INftNRRB/yFXsXSO17TIk9JIwSt3/8plU6I6hpATu4t6rkd+qZNViS8b
anUdTzjL8RUTdajRmwiXcGc/CFXWSaRtrwGsvConFICa98HVeq/81xnnJJVeb17T
SHuTdzAOfepxzQUtCpsz3u0f+WemZjBSKx8BwYSHV5CSpuU03GPFdwcacSvaPiyc
LGMLOwGlBKOFRQDGEzZLVphgv09xxjcon6z06nrqtBh0dxxIyqgajHhGTIgBfV9I
o6omxsZwyydXpXGU6u8DnejShc/myC78ZNtWEYowpymhfCl1mGdTuz0MAY3oaNf+
EGhLBbRWiGf6lLC2I9dTwmBSH0a/OzroclmWF+A9/83+AwvjtXVGevR+iF+18IsV
V+7BVYPJ2UM9RwBXXdv7H1ZzCY6sdXbZW2NK14KtYneZJwZ54HL91pEdrE++Ztuo
upDLhRiX2yk7fyKnC4ic/G82rNXelc/SkfPGB31UN1h5IuDIP7t0Vw8zt/pk1/Ov
+mxELKHNycvdsQ8r/Coa7LVZfzla5xKn66QodFnAn9fuVk87yaJSrDyB+QjTY7X1
f8iShPu9g0RoMbL15hBnDzZy2Dpi4QuvjtMWGN0aOVRICn49WPMMQ3pPTANWXJhC
KIvdYl1/KCI6FjiKiAGymtAqbTlTPoHcPsRZsg1g+OqNzJPWwuLaZ6/RqEOFSRd+
vfCjW1XAedYZtDIN1WppGyyt4jt4zP5y/h0qLYPdvK/MGC5gLD+TNaLY+XiAf2qq
+r0uckyN8uM8Ig1Sa9FOimMK97Bg3vZ5Yxe9ufWgYOwYTqNp5Z5Sf6jPUZL897FD
LdrpIjy5R5Q8KNdB/MQ/drmo8JWehwMhULq7Wt8nJjVRBp2NV3R+6a8tZGr5Z1mf
h3T2SN1mIclXiviythkPpCoSutmwXTWVZgTWSwaM5x+DfvB4dWxqPkucx9tIMjL9
YcPpkMxBsF0FK5wVtHkAdAIH7mah6SFAHm2iouZBe8fOvmGNMWZUUIsDkzpQIu/K
+o8CdBtnjAEAAed9r35aqmzR9r+oLpDL65JQejewR8iweg77zwxjsJF8QJtG7emA
L6GTqullLWKBA6XbFlpsAy07JroX6wH/hLogZba+5vSdKXoojN7fs7lKQTb6Y3VU
t48VtM9PQNMqqJtAVzcgvfSfIwraE5ngLgvyfqCBHlhPEWc1SAZy8DyXR0wcY9YQ
fuae8bAp5DXteyDMEN/+0SAEt/+p1zFrPbWePxNq73woHV2Vzz93fE2lUwNmS4s2
5N2nUcRdQs5Yi3skaxTTUxgJfZ4vb1W6p24Y/Xr6P2ROhmXuRDNr08EPpepw/xo5
kZcdIXgz3iT2WMy7Dv+empL1fFbt0Bfqm3TsnPfub4nO4T6Y0DmauoVXFK3D0St9
sWlBEiv/mHVRstuLHoEMC31c8RsetJhD+XneN1O4n4Z59Zs4qQMH6v/7qQ5NXilw
YE9RGSsvzE+CAgYFyeeMqND2NWQj32m770qD13m5aTN5sFtxaQoRnNv0aZlj2sZi
Elcnyew+wojD1eVHeG370XMjCMSnOJhhlCfkQxbF9wKna/rzFCotdKShcepOA6Qg
DSPDsM5ZvmHKvojOSSzHVnFsmZeRHVyh5wZFdI+L49bXaO4pMCpBJD80hB0ekOi3
W+m1j4m2y21Cn0Dzb725R/dlyjdQ5nsVPaBZBRGz60R2EyIuC00weRYJiwU9XYO3
0kfONRFm21pbw5Y6+OoftQ8qS49rnU+fkgM9P7LGhhVitbCXJ4ZSkTUx7FNxyYQr
751lsx7B9YAa3w6oVjF+21ZkkiVY68hY6KqKeFzgkrhaWW7JVi67agRgmyfpFNuk
kWvluoPd+NaX/JTU1m9RcVx4XnBgcCQtC1K+0gWmpBlSho35doq9i1Ak7tO8j1J1
c7d46nQdhXrlg6oIQAFzZAWNIKHgmhXWOYWl+pP+oCZi5WeHkewBOVEFMwKHYPhJ
2illZlh2OWBpWGLBhs/ufJm2dUmHV2UWybJ80skgXb/9rSI+qx+gQ4gCmEQ2hbWZ
qbRtOYAyrI/AOfTd+12Xne9kg6WfTsBxWzsOVEhfqzx5G+cpT6yceGQhKyQZC7rd
pvGHk4n/UQQnnHzPA1YF05omRxE7aa3mb35egTQPp9z2B1NcaUUEV7KckzNiFzfB
AU7qHb0kCZ5n7CB6ud397/NsALHSafKYLfCVpwM7D9JIprsLbLMq3yptoEOKqKZo
zVUvNPxV/8nWc4glHNo6duOxAT3vnz6YqT4PHxeU2vdBblcuMltjkMk0tgB8t7Dz
zI0TeQ1TwhapfV0jI3Fz3l+XGF+cQ4W+0sJP5clkNqH3djenuBUTEZzmnsncsW26
jCEzH7ODusSfbJUVBRygYG5hzmBVEkL2E5SGNpyTpspYEt37iBttpVgKEGBubaH6
iZ+J9yeZsatTzcDSw+QXiJjcRXjCZH9jIjFY8OEeV7D4AGFwhyP7fToYbyaSHvLX
vlKxWlFJMtA0bMXw2Mwhv8jaAKu14awuwt9Ho81qUEbW7mKS+bgoJhxrFrvyU+kK
NhC37RwHl9mOOl6FICKnJAVheGPUfSiZTkHOJ1bT6lA9bsWNMRy5SEOiYe6YLpQd
rrrecaag/ilvdK3Jpq1Y6gCGWgXi1jt4NqXgpWvhaHTg+qodnKSa56Ty26VreyXe
Lav7Wr0p3yY6vUbvNo0PPr7jacxLgmnn1l1Uh+9gfcsJQTyLMTYD/pm/ZTvisvCJ
VI3XlarhWlLn+jp2w2MMnksofAKvHs4jGsTjXzFK8aerNXAdINCHDT3Iie9f+v9Y
C8e88JkS6nZG2jUzEpyJJILHhVw7iqaLYcBD06I5+KJvO/e04AiduCFsZAIhsrJj
AA8zlAsB1KH92BSe2gDi9yECe71A8/O0BJEGJQ7/tMPfq9WllByqXTxWdkL4LSk4
MQYGBfuHOO0XF17BpK0JomVIQw5YZW1QEP21aB9PyJ4vkEAzd8doYEJtFINopn+X
o2a1BhcqOoNqotEudaxdhw8kKJMOfcN1d1TCOuHdtfPyGv/a/smlU/d+/ZMkCl7S
1Lgfan2tJdEPdDxgF9F+qKLF3eGJLz2VSRveloAq8I0DnCjm9rohIkWNLRZIg/pe
YMZM1ip1ZNnnL5dFbLM5hN6dhPIr19FfrnS3bwy1ppXWzVc6KOiCbytpiEywc1fn
Kq8kNdQfK3gac0Rg/i+rF4oQf4JP+Nm3ZcACXP22kvGQGNCPKvqImgWjvNcmI/b2
VYu2iPx5sqoL71Wz80XTmvz1lr+pn7aeyCr3dd373u0Og2p6LU4+51xb2m9YB+Ex
o7k8Tt2saosgUkuccXM8jsXoNOhBuKX4w6gcYspbXcCu5YXz6bS6RokaXzMzfqNY
1wS7sPdG4HPuazTRoqEgM+A1ZJON9Gl+d0sreJhSmNJFDgprM9yvxeu4qOFqSJjP
ArM4ztlI/EBawbnlmxOXONpQ46BAw6o3MAOoRW3CMtA3nWD4h3fein7isuHhzZfo
93fiExoVb8mtiZRz4gVtAL3qtyaKL6D+Pb90kxF2NNp+jaTGkxp2IMOBcpieoEoO
85/Krq6rQO24RRQDkcdWm28A6S722+o7IwgmvtqBlYowKQNNyX6m3ViMVkVOKIMD
g8tfWq+vneqZDYYK4+wWMabtSbFM+dQWN4lfa20GxzJVuzVV1PlP2tG6pSxfFHdt
aCnsUD1jKYP46/JuJ2JyecnljvIC7kZBLSyfACE+UBtr2VOOf/hBg55nV+Cs5fOz
WtqGDCiXDqj+bS2d4PMjLHW+dlgde1ZTsqHM6Q24MtMz/eDtnkNizkG1xhQkvTk4
z4exMqgtRKdRmN/wocJiJFJu07uWiOyPeGHAlUj7+SujY3nAc6CfC+q1bJk2RBy7
UXhN5KyVJNtz9DBfTPNuRmydqXX6+hKtvUO0b/yPT5QVJh3Nmu4j1/KPLQvsi0GK
vPbVYBiGRBDY7RGE008I8OhC9QhkxxdGofF69U0urw8H1l4b1JvkbtngW31oXL3C
uwy9FAeUAxEfY45rFFw4spETJhs8ztrcSHw4CvZFkPkILAksu8IHL+cbI/FMADna
Dmf6L2F8eeXMkHpUOa/cstJPBRCb/DzKSjxXnyVGbNmLbLEcLaoXMh8WnPiwfALv
T6ahU54alcR4Lnh4WtBNrHXTEKguh5/OqsENyzWbo1lXaSy4atjV2XPfldJMJDmM
alsLiU5g5td+AwuM4x6FgC4NIDqBrTtgbekG+uxsXIVnCiCgYWYYuwOokkraYLxI
5Txpn45wah7vgH2g+SYjkXBbINCiWfDAs2aThOta7wzK3xwnJCpapTzRy+rhCO7E
sDDlik5IerBjFRY12PjdH1xqrO78ZWRqUt5BeJgDnyQTREJ5+z2M0GRAU+M1kCZd
AMNFfBiqWa+AboGwG2dYlceN7XTyvGwIL3/zLSALsV1Oq84vT6WTn/HSVAKN0obv
L1d8FMW/p5YRqkhFsp56YVgDVBLtcbWYB891ENxJ80SpI5ARMDBy+1NRj1waLy91
KXvlOoI1evjTSIkLg4wViALRj5si7knV+RT02Bhb2kKJK2NCYDWUlHXXyuMC4t2O
dvqt9FRt10/u2ZUwyE/vRBGPOpsi7pUAT5jVS2n9AVTlNaMRoSgsVURFHLsRFylY
65mFHX+x6URK5wCmwu0dzXjlUrrOVpqKSgO79Mump3KLOx7uXbRYbNDXIAzv0tm+
XGmfZOdniv5G6kduv6dfBJRy7CpkVl0G5tiPJ4wNu8WFwUhmM2oABSIoVR6VapCq
KQvDotN6JOYIl8JByF3gAZjnf3J85VlP15cdfXT4Ot4dBDOj0w5TwTLr7FiTiFdK
nqr8XlLg4nNHadBFWcEvz3WFusG76akrbWkGC/R01mh6mw/mG6rRYm2sXvsBYlhC
LMD/NKtcxhnsKaFvX6SbGQSnGyU3QyDZwytBUlj6Ss5Rzap/22+GVF1YTSePdhUZ
kaaX8ojwMWoobeI98UwJc/a/7c979/MZ8Ezce9RNJyGZel8pUF2zYG5+J0DCXhvg
LbLoCPrvObG2MH5ZtsWs4oJ81lT+OBq+F745VxDcD9ylx/oBQuThe+6reyZaFZeh
6hgqQ0clSPOD9wJTQXeP5dA9UPr6Ci3yBxp/VzsQ3f08qp/I28ZvfH8sxe7HQ0XT
Uk1VCirQA56satGPFpVWfm1YjD5T9+ZMXoDr7l1mfh07I3CqB8GGGhhRwOOegbXq
NBCDYqXFIrtUp0KJ0Pv1dJN/KqOZAQdvrej/fqtE/eFnXlmrmSgCw7Qf4+x8rHI5
7xquoKyNrjeqPpGLCjmxJdR82ylwIrxrL6PrBCyFY02JO+9kiMbBlcF3VYsUgLEN
9i/SEgS6Mbh/HMMkGmnzYL1564s6btrpLgjso8Y7Zh4Xh2bPRSKCtBYQdjIOR563
kaJB/aJcaM0LStchCv5mSHlb+xRb89xgu8SH576fF8PmC8Ubvdq+e5A4eICh2e/9
BQ8DOycUh3EfprrW0SAx1W8Dp5Pkr3YWHapS7TJwVISw5eQ9WzETrQ2JENevQTXh
5wznypns+O/ri0SP9H/QhG7J87umHayPmBqDGQrFrAJ5O1faJRs0sfw7lC7oq4CJ
rF8PS0rYuUVCH4FQnoDq4Oc8CpEF3NznE1S611AYeFSdI9yfv08zbf/ArAztCJIk
o6q/kBhMtPxzy16D1PyNAm78W2lLU0vBHQr3aY4zeP5ytgRUQhIpXOTQ0wYMDCUS
YBc/f/Mo3PoGfGsXxITTI2GFIkZrk3srxH7IlmEQbg04zOjJXLNqBWFBTbKMrH4C
wri5GmHeqeCi9nadO88pVBy1xTDgKlhCkrDABjvvk4uiqNA5KA9uGTgoYdMf7sRl
DO7csWu6dAYNq/4d57bve1ydZU2tH5Q5mHsDqCPtQm5suuy0ZaW/bry6wJxqunhg
KPnSqlFktrfekkaCB7r5bdZDWu06a57U2MDc8OFl0VRtwdZwyMMeZm4yW6nN6U5x
mD97U1wE/EYkEneOoKk3D9sAjzAtjhqNruQG6UM/i4S05qAMzGB5xeBQUDPOtVjZ
fOxyxVXdq7oV7KO9ue9A8JQ88LHtwLueZOpqu6tFhLVn27JLINZ6oLyRp5KoOcM5
J3OKZnZf8foMxGcH2uJ2QpIzywC3GseZnN8tDzoZDwO0eEC6Nh/csVufjNuPi2za
39yt8B6QH6DR8ksgUgNENyjoDSCpEMv3J4VIvTtywEIOH4S1DTAUgQX0R2AHMdab
11LIrUFApjzLhsFtobqwuAUbeFnlYhDJBh2hwy67ZbKXmMflA5ZuaX+Cgs07bVrs
PMe9Itt5DyV5PtxLMWz19W/OX5o6UA7ROu2r2C6gq749FR8LPx/YqwX1jMF/d8OY
ZAWjAWxSeNf4Bo93fEXYJXxOgcA1YN7J/3K+0EZgh8V1Y4nXtgu8CtPV7KQIhyjS
C4FrORQiGoeUACilRbyhq52J1SM/ifBLh5Mq8NjVk/QFhD1PrBcXx1hB5/L5fcYD
NOldAbeDSA+M+GqsCM8U7qWAJCkAIyQUdZZN0cNrqx29udOlYELY5Cjcy+Tjg2Mp
llKeJQvVcPw4wJCL+YmUIxjJIWkDpWsqidlDdUIrLD44VeuhHrQl/dx1ASAZaef7
dBb25iTRFRo+ICVEh2uEZb5BziG2agmFENYTQy3aO3uDEFy5PCnvcq6gzigHa8Bb
jiK/npUDbaM51ULsQCnLDWuk/gtjMPj5tO7dCMjabnEtXCz0aXqB3IZOHv09714g
xnHuKcVJtv3pOt3JnW0FbO9w38IzYuFxfqGyls+HchhAct9tHcUra1xRoQcED+4+
CjDQTaiGnjKW3WdzRT2wlFVPtUhrR1SZHR4Eznbu9pr/ngNkhtisZXNccAKwM+m+
0nVXzCmjgapO9pLcbUv8m50GggCYIMtdXzIcTstRJQHd64PDWcLZXrrajY1ZaVTZ
s2RLE1W6EXiUlbdubHZmiFjfvKM62xL+MU0zFuqVV9GYFK7VltRudnyxcXar5XzD
F10g4uJp0aBhObBwMoYt8nHYQjEpiA6xPuO4YcordUhCoQKIXnPfAVwG1pXdTBIf
Iy0xND8PIAt8sRC53z6f2DWKfFcBMXvKKS61W+HkFA71kgGHxnpnimmdQrEzinD+
YQa8YGcIIgUSv59zVqVPAfN628UFqkaRek8vKoQ2Qih5veIO6x7vVcC3V8pfYD9Q
Dzg1ZqKwRAX5Cg/F/OhzeJUCq6z0E5EqFCed9chwWi0ZrU5J+7rdbh27IUrlV2kK
ddJKaS66/e1H83WoHwUHEDcZqN3StgFrTjBbOowS2kaz2/olW7FhTST88fylyxSz
+ATqVa9cJZjI8MLDRq4cLW7gPuVRHv2JQMB8gcBhv6351hk/R4s71vOvS4YQZWUW
6b5JpQhfeLbf8NVS5tM3u9KuVrNytUtpd/REG49MuEXVHb1hPyCeH+8tuxlc3eyP
RLaYojx4rQM9zzZoCOzbMnRWkPnfTQHo1xoZQhgMNHK4pWDo8faSvzVZgCumW4Ui
VlHkpBP0G+JI9NM6ygBOxqvk698bXRRphZsRn4WDYbsnIXO75FCci5Dt6Cw3h0w4
E1+HSjKUE+HfEs8f9x3o8SKcyuttOo4jydMTIZfS3IMzTiHyu8firIlYDNXfBiL/
awMqUgiMktxd+3AWvOD4TH5+WZndMtcn7JAE5izrLV18yug+qHUzypQreZOi81GR
FLV8QXnrgoauk1cURfYvN53bofaT5UMYP3w9CvpUcU6E+UlAD2xCM9QPazxImbbu
NTNT3ZHahDZ+fnYeWzXf2SHs2W+chfZVnPrVIDcp3sRIDD+D0RXNTZDB7w3+30eT
NnT2ciWTrqB/0OGh/9G1fNnL5EEF/e9e9topqbE41Q9KhLNkIIuK1Avm29ZD2/T8
eJY9so5eFlPSfVkZDBqbaUHZoOYI117L8w2E4WAULKaNjwr0YMitAwotH7yOesQf
vEaPm/r707TFNV081NnJQ5TqqJewpQvZivKXYxc5kReb+GFyYfIG/xbato3wxhP+
CD2CcLdJSaGsfYFEufGuaCzEuYL+OEbO1ywSwnsCeDAFkgpZHxBmUAnBtotaQmz3
AIDVOmwEmQ9mjXWyF7H80+OMGZVA+rReT/vOrGKw/hsm8vMtWhQXGqsQyabXWCkv
Yebnxwo+3C55uX9hiFMnrzzycpGOZ1VOo9o6Pz//0J7/cDdgOdjoh8YWASgSMIIZ
3MvMRiIZvaXAhBinhWn8k1OXqviNqipLRgHi5VQ89qzDFrnkCP4dJUG6oJ3vhsFI
i4xWRQGvSelZHi9JMXXyCu6iSnDuMcLKqFIWcvWCdxSNkiYhYcPiR3d3EiVObawa
XKjjwpYdI7mZqzfnVc/th7eAxj3bEJwWPDJoIPs9Oa/9jA3Pjo4H4b+ykAITc5la
8RWChhjdfwgo5f0DceNjaobgmeovXEoSN/4JAx1H1XfppQVYm4okjpvRvt/sMFN7
zIoLTyigf1lOMLubP2j42rNgYa0eKXkODwvBYuMb/EOUbVkXZGc4H5CfZ4JmD8WB
83p36/eTHH9cVu+xOiz0L4F9ybjE7M2qDj3aZPUylTdEqfx6mjOsbIOvmQJ8T7/7
rNzT6Aov1PQ+mEz3HK3p4ac0pDM8i/fivgjHs2wekrjdGKsPfNXw99qcJX6Fy9dm
N2ShwYjgelSWqTLgg2Ax5s/7qj6/8BxsYS7n6oaUaRXHX6TYA1bI5e7IvcVgVXXZ
Mv+JwG3O9JYgeRrVcVPx1SaQlIPCgqf2E2BzOjLDH6rZNun0WiIuSuFeSayyobGd
jxobAIaoa/EK0QL5poq3cHgMDvgtDnhtIbb+1jYN/AwiupdqIPmqXdAY2sEIeHZt
ZnUP1VkPDNXYhzyGPMt2+q9+27h//4WB+2l162+TS/wIw2AxvJ9O2stRf526qfTz
xYsukxHZ5mUkr5eLo+rVcQIDiAMnZqQmM/BDQk7LRP5BtSsI5N2ETnXvJwRkK6GG
9IgZ+ztPv+Uk7ghdsK6aXsKVZjtYq/DJnViMZoZVsxU1/uS7HPZj8J72Dz6Y2v2y
1Z+9SMj8bPG8xqkXPQJXDCznBSPitPxW+0vSjqnAZiFdf2+ezJfrUu6qjvuIV7Jf
1i8Z5KKOTXNAxB/riCEo+mcIaHbXQxOJzZ4vkuQEus2Q1ZlnK58OnUHw2vynd1Mc
6orVZDKy7vpgI4I4+4G8SpCjO8DhYf4Za0QBbKoBPKk8qtFKqc/fjn9uJNQJjgkK
ich5s96P0+eWhlJKfgUZlkz0jjhB1bb6EMlDur1lVqMAWo5IxmgB/sCoKSChgEMP
SNsrYjYPJoUknAWu4VCEsHcqPoQ6rAtGZLMY5muTA7NogGcP6lIzVt1c+M0iXefR
2dz0eTeYiikxHZ5+Qjg7Nanq6hFWGLU3U7YmTP+a5A2yWdW4yxh+/7VeY7daNWxd
tQIKl/ClGaBTIweUlCfFGEK5ImAuw9TfZGqNzNMenSunZkjE/54xY/5YNotUHlBX
5SrxGx4wGHhCmqbfjwJtZ3WmzwwwQ08Bj3I1qIfLTQDGO7lLKjLld4EyAP8hpCJ6
tlafctCnwOghXiVT+dr6nRxKfZbRGg1ICsaj9gQThwsiYH4wM0qXLbrALTF67EQT
fkHB2i+iwJtnPvcuSrjQX3nKkvQRmvy6cS5jW8r6OReiLbdcuvjklme/c2g6sC0Z
S4ZMsDm38LdKFmUY7QkOBwRO0DjIcRRLbof5wVKVyclulML7vHBobRbAW6v/3hqp
z5sZzLB5ShRzc5hmGQbtRYcuUyals9gC2hESodr7YQa0348M0ymaWFWsjcJUKQ3A
pc8hGuqeUaIqZn6hvc+MsQQOtFIyBqZi7vV+aHlTCTOl/d4pAJDcBGqyckpb/8rR
iVG80qw26fyO7hu+RXPc4AJwlf7S2UIcpR/oFjxkpdUT+ZyVRDxw67MF5RyIQwrR
S5p2nRdjlIDNGccM/XgmUYrmkC89+A6gvpgYeO7pKSrDcVW38EinFCyZHYN8a7od
GmX5wzJe3XEWA5w1AyHkVz5J7Wb9NU5mb4HPzHdTau4GAit5P1CVEHuc2vs4/7jy
lqLBCrEcjjiwU0sg3ZRWDgtUSyeBXEq9UoViJeDMt5fBKcclSyDPLKgo/k6Roj74
Cluk1VKt45gOuE3WXkIp4vT2pXkRIA00MdIspvOflrCf5LRIejUlkaDnuEB/ipY5
tgcjowF6CtHlpPoUX+suflzpj9XFIej0d5mpodqX/YVS4jvTZt0tOV6GdeMTGFsE
Vaggar0IxOG2/UnGlD1sy+vpU8yqGhWwNKKXlA2YQffpro62TGtD0J2X0uwn8s0l
Nd59jv371o+G9EulDXzy9KjLqpkcFVK0fHN4sjDE1+gpnetSNb5Hci3YJqIhKZ85
eyHFdkrwMyA3dpEL57xsBtCZoY4z+1Yh97splEPVg3j1zyGWqMA3KVd965171H5p
VWrEO3XowL14xWAQBf9ZZWHL5rfHc2kP9mnJ7s1z2FcWNwVvp/EBNMwlZ2+mfomv
BoCHLF0XuePiVqwhIZZxhpD1TbozyJpQSnNfKcIit8DvcvnAW24L8vbRk8Nph0e4
GrSD5HT9YnWqXwIB10LizZS97tPdtC3kYwua+2/38KNDGy+f5SIrDrnmGy68HgSA
4stQ4Hm7uTQ8F5/1+vSBC8+xhVHxVcHRKcC/ZNtE485DdnRv6XSn7HmPk0dip4dw
sG8ZVACofUhyd3TK8ry8mzpcu49HOCF4YrruBZEBm2xgYZLG7s3kPvThk+8wb1Vr
HhYsf59LwPzza7nVO9cHE/C1UzMLbSCtrVgUGMHg85UDHzqL0IyyiAtLKNvIIhjN
Oa/bDAKzt8HxZ1S0fBinNXB5oSI3cxg/EFYPsVzfBkHrdTmnK6wPcHu6dpa2Ojwt
V/v1e6lsDSmK/3qBXaSKxEdcpMT3DUxb4EBPXjHUlfAKHvaf9XRHJdjkALWyeaPr
zPifrWkaSGLc5zzhf13aScHkNK+od7A5JG6nzprlXp9/JXhFN7tcJKAAV0tI3ljk
yzlq8BuiXCA7YK/Rr2hympkU4AjJBpD1hrrPX9U/glvIoyy70NLXn0BMOmNPD/K4
41VIFkoYdKJDVZ9w+ra1ZriEzf1rbzoC5eusrbLq6tCoufb7PB31V/Q35IFNC0CP
+bbi4OvY9uL/fWIaOB4cf6SsumfyAifdIc5ITfYeOtsFlIve3Y8X6jR3Cmf2ph13
SlFtfh9g3SjNz9zILnGzYEPP114y+X5wBsQh9HmGtOugZLO0BC/aUqQ1Dr5wF/tP
wqA6OcHoXSiQ6zI2E9+aQJwu0Zt/rio/FA/gm+v932gyGEd5pWnq1LQYn+Nnb4QJ
QuuBsBhNJOnp8iZ4m5A1Jksb0FIYdz/jUw94sQpZecyxjgs9zmwYqXhVyUgeQNvy
JmToQCQjsQNuNHwi/czAy0E2S4ofuHbfKWuHb2Z9z6DIgBuHqrvH8Z8heMo5nMjr
8ZLEFF/S2Q8tciy9fhmjLTv+JUFcjBZkX8cgqs3CPCGqlAbLx2WumaJbGyvcV1hi
/gAxmnIQroWCS6pIxVtmdXNVsg2XorvgbV54TO/2av733B4aMg7rR6KG6nHVHK+e
3efVzbMqIC69Cn7rejtvxdooVJJD74djeyHJDfDzWXWXIu3kjwEO4RlRCI8qSwuE
XXXl9gOxONmiiu/KnYRD9gE1gIH6xjvnZGpePHC1/uCv1MK6jbi/hrNvOAzzwdq9
cdAeHRpYAwkFaEx6Szdy8LzGZSi7GV3HzZLA6CTznFSgk49EyakXTU0slAiPKi4i
CXncO0Os5S4zDPlAs/nDC8UFCvkwqliNM2JLroWapRLmTiLba8Z61N3wPgsYzi7Z
NIKDgmvD4L1/dZ4eOcpdQvxInOSFBrCsqBTxOJA79KsuZO546ScDpjRoNiJvOT+9
VAP9gd3iOBBGQJnQlsOelbPbrAo1CgYS2WgM++4kQBbcNa0CZMOgPxhdlJRa5ihw
XfS6mhklA9Yor2Qh5x5Ll66vyYIcVTgIUv/xvhKqLp42vyJxBYhb6R38S0tsFkvR
nHhMdS/ofzs0sMEMUu02jQ==
`protect end_protected
