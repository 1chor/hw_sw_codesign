-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
X/HYbARTxZls7l1RV+WWQldNZusxY2ikqsopreu+4EGnBgLmk9cqbmSUUhkyxaxt
JoMJbOGPAp4TOpjqya5+F4lOUsVkq85Orqn6UQG8aYBA/5R5yxzg9a7Q+v+5DRWB
diAxJVX+B3OaCSj6Lrff9P9hgosXBSK9f0Cr0kZqTc4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 52256)

`protect DATA_BLOCK
BU64JZPcHklHwSpCzOfZ1MuFsFfbHNQvyGPcJTXwdMggwSuwl9HT7uT+dNg6BBOv
ariacQv5buddR8Vf/d4s2OD6xJNZpycsEWWDc797/TQjIK7A9SI5PaSmt3n3qFpk
T8maxBstFlGcq/QhTEn4mAA+Lnctgy1gTpS6z/hhhHH91gMSONXta0MuwjJo9IEC
nnMcxYfaF1nE9Mz/IqR95PcSxbEHUQjxdi584qiRYVEzyfdGfgHZuL26lo2nsfuR
FQKHH8qrd63dntX5xOiwX+0JtVu3ySnge1CGN/MlWUafGaiZVP8hanQfsJAhhXpK
Nbk7i/d9fN0BYIaXTz6ggolwS17rVeMItNMnz2pQ25MbvcHBRiLhzan1ihmmwsQS
wVOFYJJpKcJ4jXLizZ7tphnx4+hRS/EMdfwzbRzGsJ7q06uFvgyffnb1fk8KeElk
shRB9lp4SKxTHr5edp2loRweML51cIn/nNSn57zeisMYmdLDV/P9YYsPzSgDaHLM
eTIsvcxxnh66SdlUDkOKTwKPZgOkZxSgz1RVJ8NaImmruQj0+gVIhON3p8KCqVuP
1rOVRO22u9HdEbuQn/NhQBd9cJPgP+kdLHEtNelAxuYOZpUJ5wcgoUkrn7tRSl0l
eh40bAcsRCl1CC7gnxrYNGRHmYpYFzTvLvhZ63HFj7SmUo2igdATUEYR1D82qu9x
dyePj78eefiB3dn49DX0tekPPQvbLQ1X2u6nQ8fyOdSeHNQOeNzBcIqMHpTUlrF/
zi0HeXWy0LCIXq2Z65voDcS0T2h2XA/yt+zLGb67SdGEO/TTq/RNyG6UgL2DrM3Y
6oAgGKu3olEJe/5EcUMsir6C98hZxj+HTPXAnIwrsqWFqOxeHU3xqqcFFZiq967a
XPX0kJH/eh/PJreznpFrvEl5lAGk24rPNs+pNyPHCb/bTJUkkj/d5Q32QyYS1ORw
m5Z2AfTBrmk5HS2xKwOR/h6TJTJMs0hVgOaceG9N772fvBPGVYOCFxH37vrJQPyb
unS8eKCurMHK69sRb1L8jZHNrOdHVV5+SR1tmN9VReSLx0JlA8Bj7lR1LrMCQtFB
avgqqN5yi5+gRODl7HV934ptGPHudpMMDlL67lC2zhkJGd20mkqMemtX5SpJeGMT
+Y/AxpPxuvjjn0vqZVoOhRu9b/WXTfRDOud5q/kw85wK/c/x+9DvjTv66p/9ebdk
TnR4nf84vdLZ2knUdBFIf8otCjH5nr8h2FoR0uTt7UZhei1P2oPzbF42KIkmlSHm
orz7MttpIe3saN55BaVtqwcGUWyqQpsbYK1y+VBH7G0loFrdPyDIHvQRb79ZvvBG
fzdUjukRvu99xj5x7ptacoikG9MjVnyTWOO+DggFufNunDdZnwjr/7pIt3MtZZC1
jEp1w9y1LwpU5+eZwrKuEoFIKbwncPWzARP1pVOOB1YHuMjPDfZzq19vD03/TLq4
XnkMDLGFT0tVEQ9tGFSNPgJA096/aTL7C/lTIODaK5Ts/mrJxZxZT5f6jy8a+45G
8VB2Pnrmsj2BLNhvL9y6TTWddqTZ1Dvkx89/XS6m+Q6giWBJ8XoOmPttkzncwp9+
femEWYL2gHFApuWLH3DG92YI3pQHxg2j3b5Nrdzph/Ef/X1X/FfOMXxPrEqkBv1t
N1H0T7IJ0MXcdRBWZWs3Ki0A10TVTyDpG2AtugM0cqBcMOkNXbv6nt+2Qy0gjZMm
3CQNMSvTc7PmECnvWyqfXIrMC2cAk7CPb0uhWRqiqS0UcnvBO3pg1kBBMhHRtB9W
mfnfMp3xZgETfa5YHjWv39QocCNt2lQ78Dl0dsaDiWhbwzGtlVzuYL7H4Dntxm/B
loe8FoCkhcR0Eo/3ArwgUNsyYZ2e3z1AQr8m9g6J4zFSh6qnU+KgQmgtvKtm08Jp
yNDArVQTJD1kSnicI74928U+J/pbpRH0sC2Wr/i4bXM32uk3jXwXJdZ9xSIMIAqd
bVqw5ZC1oXbl6fUN4/wofUBhwfB0FUJYHq3J4YJQ/lgr6lF0aG+AhLvsxCa+Xki8
OMed50rxkenBFiptlGwhIgifnkgknWQe4IBiY82mQ3FI1y2rm3fsIFwlPEXUM4FY
mTmCsZu53h5b1oOCr8EIC+6xXLUkZMWbUHJxo8S6t3eRSzf/9sSjfenA/90rQ/CA
GMjyiBVWRPsrIT04V2OIwqW2X7VrbbbsfYLQMmyskvkLxJOVN9RcpLR2szk5JT7F
RJRK87ornb7XDfKiWkEL2ouM230utde7XHr/q1F8tUvWC8dfNcpK1Sf6VD83nB5A
DywIpF+gF+Rj1QQCOWOBac5/357gipM9tkls76Zll1QKiHnDHPY84U7FQH+HJ5w2
rlEHm4tnj4Sak8PwV01QGYahw+MvtE1fcVvM1N5vnsEoXuj6X/blS5eTYKTyEu5N
89C2KIO2fWSrksorQiK+DPoqjMFxjrlzegxVwK8mVVRBlsnQbSYZEwg1ALrSbM/W
P4kEFNUUZcWIfB4qQuxQFBK3rcpxjeMilqLGoy5A/7eb7NLIO5ep8MoX0Wn/Pj+Z
g0/0P8sbIlvktnE5GvYUZXUXcXgtpU1i5qLU5gAZBqRv5JxS/dJLp89CUqnRqpni
9AnPzM19xeDJu1qkrjab6Ivkg0W0EQ+evi6cnhDYT1w37Ibi+xyNyldeRFxBWX46
6cyvtagePUTJNttEsTNU1VIFeFfQBJEaXJsEwncYibJSrZ58VZko4BrtaddXCkxu
nc19sMJot4UbFrn+vnW0kqwoxd94LJG2htE/eO8C6vHbsHvdx/0UQOprcVeNkFnH
y4JmEDe0mjaivBtXJq/62uS48a/5rhyxSP0HYEM2HfeLjNq8nhxNEb3Ca2aY5Lu/
u/znhE9oJOZvwRv6wJFw9NyLKL4ITLK8eUzWLQZBY2gA1zPJTkbrR4Bph5MrCwZ8
zyAB3HMKWQiwoMb30rHyqVxOKvv8uOj5fuI8scaHEav4JF17puvQwvHnU/WxBD9W
f7lsMjfONxyMHZjcQyPzrj+pzySa82YGSL3UvquH9ZfqlHUNUcDTftfH4fB8wUhZ
CVCaxqUlQ6PObUh+5zt9FbGtMyGxdPcR77FiuNEusExMKmrWaTx0lZrF63u5OoJn
D96J/LizCeG+4ZAkvbAQKQMfW/bUu9grIh+TuBuRmDbS1Ht8U7sItxV0k2u0IsTl
/Khq6wHO044IC0mFgpxSsYhSru3/KCwBxxQ1IpIsofL5frcYrttQxsJG6i+y70Ay
nido8muHMCpFs+pMzAwzyAqEOtWqfOhg/4GkS9xxaXjvhMg7aXhahi1RbQjQz+kM
AqKl2t7YnlTqdSRQ69TCeMhcOyWGUxy7ldr5u6gswJ2Lv61qu15xVne2YnbKavQm
9fgvnlLO6wVlPjWxezH2lAgiUDJTpEsJpA3lCcOV3n7tGpVcWoILkXjcv0B5P7TU
lkvjk592M/DFbnuS7r30gDuRdnUahtm4MuP/ms2vRWSN00nY5jzwXSrhBaXToBwM
1zzpeJ0NeX1h9iMvQq6O7/ebf9f7DBQqCIUmnxSA3xqjbFeuneDGkNUdiw4MgjJd
jr9T7vKhO1wBlHfhDpnAhrVOngmvoFkAnw5HxLzRtSjtdHEoO21T+qL05vBa0qf1
+uF8Wo6oIoM3QGO9mMpdC4FgCgD9NNRu8aqDHY7//7NI4VHaCzgA5j+FpWiWedtt
hFn90eSSYeC0iJgZff7panZKFOyfQ1dcgpky4N6AVtFP/aDX2Hp4XKRIMV3/gFKR
OvV7Lxx3MbmzdNMsMjF/2tAGjE4vC6/s4GiCrIuFwnr4GQt76dNHJgFsrOKwKIjD
yQH4SQGR1UZvRUZ0TVhBldUauE6rJaAtN1UkQXDUHvCtYq8JRexBZzlKWYL7v2HT
OuPK8bOzWcGYZgttY5wGbv2PYluycHGwNcFq5Th+7LSXpw9Fv28QAA1lG3DB40nW
UToIbbq41PGIJMD485dzvfYFIwehmZGhyE4LaUjnR5APkEZUif2vvNwsGI56UzOw
KoehjDg5CCjBcGuQoLt7hCjb20SLW+t9Wq9TyGkqzGwNfhvi7C/CK0MNwjx+wi52
PGudhpuI+107Bc7NTFyjv8lT/0GPghtm5BGLAXmmyK6VhmctqhBhj2o1JaYbUrQZ
jXyTsrPOXP0iccicXOcR0h0FEjv0adIjfl4N5Mdbq9Xa1ZhRj9675uAu1Mfub6SZ
abouXGti00ySFTZ/ciZQEKRbpvmZCnOuUhu5fZ2p+Yo2pamNNf57AzR5Yvwwwsad
bZAomtdzEnK7cYgkb+2KnEqFd4IHszerh2/l4mkVnN1tLa1j+mGKiSw+J+Px9mFl
AQ3NQgaKUBeqm7LlOlagylvVwqQo1KVzFzN1wUkVrLy1lZ41h58a9aPKjI13TrqO
Wq53mp+LLlQVo3MQpaLbZtwI9+MKrzdARyHip7VEsSmK3NNCFweuwIPhX+fayuxP
6HG9hv2yMMO+Wc8jzM0RwPVjywxxe6jMBqNppJLMrardtWGccd/mZsfnuH7iLdYA
ZTyz+QF/hxIjZOEeiBeXl4aCQxWRmzgsLniKrT6lTtJM27Vz4WbiXethHGGFXgWe
DUYfSzOt1pK+YdDlD5p10UhbCbh5W4HVnBV5S34uZENolPGC9mjXFn2Edc/NGF2P
sU9RY6bw1hl4gs4k536Mh1yGtP69LJXWJKbpVfohnD6iw3WahBt9i9RhGczmy2/2
SE2lxIHf/exScRymZcDyT3UlM85E4oi7QQ9lSX1z+qNLS68TQd9DkJOLigMVvVeA
GG15m0rX1tiNgtPnAXNlvN9/xIWgo5IWuSpr3iqMSqKo9b57zK6Dof9cxgf2thro
WIX0Y3AC9Zp/kdzoba3Sm3DM35Uinfonha0KhNldT8CzScCrbeF9pZ/NrfFSvM8s
ntrQWhx6pd6PQ/G3k052c0BgvEOZLbSX6z74vZi/e/JCrZviZSugE9u2DAK4YJ0K
TESZle8M8CIG0x+gBqQNWBshwXKj2Ef4CRNZsufdA0nEhPV9SZsC8XnATh587dDB
h3i24sgG8CP1CJVD1vvxNFc+1V0XCx/079IP9XEkJ88EAE5BYoYeIMwP4WO/Kzih
f99Gf+H+gipW8NtVZQwhUm2VNkYVmZOZf4lPB8c1nh8gfqYhBRoORF1aXRzxsGA2
BnHGscpLuxg+hbMow70SyTjqelbHerbN3D+mgUBGjNq0re3vsH0XXZHj9rDhR+/d
M+BeVu7FjRzInEMZiLOO4hnBeiCLNMPvgRoMEAwF5aDGDHTb5ThoISmVbOq3/Kz7
Z173PmB1Nh2fGq6bcr0MCK6SeauGQkA1ZX/ogvchy6i1usb+6HBZu5DtJTjCqTAT
RX3WsgxYNHXz8bLzVvyHQ8Iq2Hr0i/uj9hC9Yo+2epRsCbO8jmr8N9VhTZ+GVGdV
PubDgFWi2fH0EILJ2R9kDNezwlF90KOA9toHtDUFIJBBaRCTt6MndOed/xY3gZDB
wYh6MiUhnLdoxtODsqD7EFJZ6UH9PHGuYkoOLCL9KAB5ejcawLsJMHJO1iHS4UYj
UnlcD4u44EZ5J41OmhmfTb27hKovqIRSzb9YoogZtFob986si79KsHJZK8XdU9o6
kMq5Civc3IT+FtaTFAJr5zdzARGx0jc0WZswLdJnK9uwAmxn0+Rw8nBBsfA8kvYg
eBSCG5XdigxBEGRYvZUg081sbKfskJlyALl7f7CbjNAxkd+sft+AX8uHBoGHylT1
S0gNcgln0gnBGg/LdxVBd6WFJPI0osuG0NR+QmPC1/qMfmxTgnCTebFVrHyYKNqJ
8ouF0Teq6I49UXmg1sgaYDVWwjSmlCoBarDCyDXK78hREY28W3BmXQqpflHLFhAq
ng/I+uHaDRHbnBKFSnfX+Yenpl+p5zdy/h56sijwdyVvwneHdx8UBjvXZ2JFDR4c
TvbdZfm+bphA0VSDdbKxqegTBQbF8Yxy58Rz8w5p6jVXm6vEgO8Hvz/4QAPaFFF4
gVw66GHn1ctAdsQHTKPBiWVnSokmNsBOtjXQyZiYJc6jlmEPfRDnEKyvsx2XSjw/
9HN/0idp22RF9Em5JXdKbIx7ZsWcLG3Rlm+lwDggo0Ry+MJiH3rn4l08AZk4uBgb
/V1MrZHwOasEeJKE0mIaAYCardFaxeLSUxGt4153IUWsMyyz2LAD6yNf3MQLnuh1
JKu3ZoIVRS+5uZBiNLbybg8WivjMZIu9C5o/KOribMqUT66k+ZI3yJnqYI5/RxFz
u23MKH5sE5/BPDa22atWZtCBX1vqU9nFz59LkB4CGvDPMlfCxULzmI1h/Hj1UMct
ZZq6GnGXah+7qh3La3yQiFNTcz5JqnY+ULrnhhOorAQDPlRdW4zZzqsd3YmpYNVL
jju9Mq9QdePyVfv1DgoTbVJ/XO8vYLEmV/2ZIuup/pIWJsQAW9m+Ea3OQSmPc04O
0PHSPhCwvHh6Ygi7RXM//Ga9FBNZWh5nhaI3pjBPtg9mWtjiP5Je+lIa1P16nxvn
vE7/A3GPYIjQ8n43P4Rq86eXZhquKYiZmwsO733pFQKdU+ktEGjh4cCCIzZT2cJ+
RlLuFdtPD53JHghEtCqn/XtlCCKWfqcHSMANjF1dtiVAMkohXMf06c2tuXG2al82
0J+fxn9m9ijXkLqVXlzz8fbUyTKnjEzHRTxLCa39/1QiVwU1OrCP6BNB7lYXD13U
S1DUbnuBp/2jOhnlcUuyKwetOtedcF7USKxm2vCzypoEFLPb1STX34PYdEviuUH0
+URRA9qTw+nxoSRMKGTQJI21vxzaghuio/CM0ypUiHaU1itPKnK7Svi5k7nHBG6v
+dBLHwCy+064t/VWLoO6DsQJ0HvqkckUBp4Mh81aRyjxbU6MBsDGABX+qq8tqZEj
H/esAbvu0tKbO3i7g8CY34Z6JvoHyjGyD54nuvj0agZZyI++UhJY2LL6hrnYs13o
F46TrrPXcJaCnToMFT2E+yTbEdBfjTe8G3/vbLEtgLMUBW8iCUOuPECW04m1TODp
wmBxV0pqbMOMVzs1Om1FcP+3C4NxPSRDMVTSBq4h/cLDceoufIiC9j/3VTpEd7jR
tqj+ZQTdyZfXJ+sr6ZtkfiE8XXubruO0C1EA8iuqDYjvF3yOzt8yK3yCChQIFU4D
2o/rUkj7vPItKz/fb5YRfLOFMCWIHtM9SfEHfVwPraNYXGFBvWMOvpT2PGEKlUd2
5vCUu1uJrbh3I8nYNrcSeJARGPd2/MVOZ1lXzsnfUtFMevruSIpP3t7n6puvW45b
ud2argtF+zKb0OYrz7C2aSgDVDLm5fr+CgOpbh5JqMYyQX+xoL57kGaGRvLtjQ07
c2QE2BNF2Cj6LKN9hC8nbdGzGAZx8Cn34d65bg+pB2LbzYqTshGqD1vNg7SvUC1M
CY0ROH1Y7fKf+kJ6+J1n7KAUV+4yBPb80rT0nvcjvzXpGRGsfsR7ihSJDJsCFQmP
AgggyISHnv1qAfglENs3v/fxpVSJ/e1ojNqTCIt5+Mowc92PWvJ7zAXwMKgKOKfX
MryANMJbm0ZsRVMSrYecYIp+POkNEo2bJ/AOrCEO+BIvLeUm5HfbSWA0W5pA+bHD
9QSGZrzZBWINeLCJXNRn/qB6ai8ZfehrWm5UDLWP0vMx/UrTgQG22ycqoj8TmyUt
WP14+MBR0GwxpiTjEISNnrPNc64DtLhqBXUuRxwVooDkLTKaRBNd9CSKmA10DtcK
tCYI/6SGw0QSSrryXUsYgZbrT5LjEZl5Lr5vn3cyBRoqXSMLiLof2mSicEqOT/Sq
kiFltyyoMeeuFnwnqtns5UCIie9bPofV1tpL8iTfCYZQTY2WCS0vtwD3+CxH/rff
A4lxKZ8w97ZfEoGl3cAvMhUx177UJXPfrzdY0N7P/CCnyN7eUinZFULQSPc7CaK1
h4GpF320JQ5nzhZNwhtK/kwBSmpbedMsxIX2Gdzey8fYFFcf7ERhs0GyHw4+Zrex
RHJHjTex44BXfHXXc4C5xUX5iFULQ7l2KbZ2ufaFILkbp3++wwKZUdhM0FrBwKOS
l1X04xrNSg0bJcQmKzPAV5InvOHaEOnRvabfQYHyTUqs2Dw2KIPUC+yrr4jHQ5Wj
10U8Em+WDCtk+TGi3NKCYrmnSuBHy1e+Q4jxhdYG/LEBOVBKBN11DPfQJqWciFic
i7dgD9rWl9JtJlcxOG7zzSibx426iU3WItVqwDuNUzH2S24BJCjV7EDcxAXdR+4k
OF/NmGhSdKPn3UWO4FUy/G5aE5LoJUoOrxKhXAWXn2aKnH/Zn1TS8H1L3/6OpUkY
QZF82vk90wEH7Pv9BL78P5EiPfdMRGf/QWTNiqJZGJ0lN6jHXG6XI5yG0UC5IXp1
7rbcqJPzpbm6RnG/GYGfHt/+AF1CPYSwE04Q57PV1JUrUNuMAXRCqhG2+EMo01z3
nP2wpbqr9bTjimPWxPJc0BM4KfXlIdwdyVonuOu+zwY9Patlv6KS9SLHRJtNnM6/
sv3jkHN+WvWl8RlNmNsHR9QMFl5SwwhN79IuvPElt6Tl4jkki4znDgUFeGXSjl4x
YpqJr5Ew6Q32TFJCAiKWNlSiezApg7H6H/KaI3CWzlkHCo/iGSjHY3+jH9tavyME
JtW4d7gIo1bxpauP1uR+ZeDiy2V5EU3QlIfcx4exMwWm5UsU1GleFMXuSrxJE6u7
fZGEHPVm9Yms8/A0g5l4yDmI1nHsVIWDrRPUtIp9oprzZeouBQqp+w9RJGH46bnH
LxI1+26mlNYABW/jMEDhQ5kDAH9IQYaHEEV3d0ypULJpS/FrzrW/fNIlFDxd3nev
XLZDTIHkIQpXZ4Ud9Cgn8Ck8mGl9kTMuK0LbttY0w/MFlBJAmJb8HMOtPxilMmQr
wXL7nQHypj5KqhntzO7ET//qZjloeoh8SHXaQNOYTnG84ICalorvHyOU4wq95+dy
ED/WtHmyDhlnlFGCH5pDxVQffn/fUD2sCAGS7M+7COYrscurm1e/ObLDdm5HXRfe
YP7TsT7HOXxsdplqAlTi7tffrN61X7pcyfnLe57xAQgxWhZtIz0Slpck7Yt3cNqs
MxRjmSm/+UbxNF8YzN4RwXiyNqoilRXXzfC08rbn6FSyGZ/j8/2nto8k4cRsY3hP
GcI/5gvIm+5yYqRAgx9EQClr6KCIxLTX4O6oz8xAtvHVq32L3OxdSSEn3uiU+lXl
lcybZkGjdrbwY3Wvxu7lNpQK/oidgH/rphT7qzdIEXbbdimE0YxdBPFGholiQNDl
lc6j6Bx45lY92fh6smM0QbOIH2v1W2GtgueIk4dGXcwDmd15K5M3Y6Pjlf3u8QSz
OkPHkSDgmFgbRFXeVQVKnSFq0D9zj96ZDjvIJLxYkGXN7XRYA6mbd+sOkqF59bVy
KLVra1tQHkMjNOPETzldoKv8uZUisftiE4rlRb5gpC+dUPg8VxBPu9v0RVUNQrSA
8Jw7E8fzRScnMPBaWwcnXOOOU/DqFuvIlyUogvhkfMNQgJ86fLFgR1e8YaicsaMx
bVen9Hqh3g0SoE9TlvsfQaAsHilIzuI4Kr0ZVLvF7G1MzHTJITQfpqi0A2lCzwGP
pTt3FInRDWeIvMLqJavF4gt6ZNqUqP4oNlF2HwJoQZe/2MlpeOjCxJU19wzcrZuK
ax/6vErtSVSBR1CsTnDkCnVcwIGfUlXuzLjv1TNpXPb9bRJ9tjzoqfEbFr+3rkB6
uDKmWAZ+USkN2ZhQ6A1Gvy2KOfRT4hmKWf7GyAWAmv5oVZaFkyZGMhZuem/4dWMk
hCD7L8izqDwszOSiBt8Jb5N+3WEL3SziLDfdeyd3ylNunHHlflVm7RPA68H0SBaQ
wNF4gxoamsnkDe2Me8s6ZVzEpRBw2M4CECjeiG+4C2lkvwkLXw4jt/IiJ/19e7zY
9nd+PEvBJZaVoi1nMrYvc2bUry1+lcPzYwSpLYC7K4unp6sidM1oa3+HXRh6/njW
J8hkfihE2pT75IdFeg/LHpkdpdIIa5BHnbIkLcQALCq+qjaGUJ9Qz6wNRfAP1m6y
+cFKEIGpmvvQ0n3hBNwgbj9jxFCdmjFA4i1zFN55RR9cm++JvD4K1k28NXArbIYv
MqzFNRzcXts7XrKR54ev8gvhokYG7kVeIxrtk/T+L6XgAm6IpxAoSHsZ/jkjqpvh
Ez7b2iLUowuMRgJN+LxMapzajYdfY1quR1qeZY7o9/IeKDd6si2XpdBAdNpA1ny+
aJIC6gny49JDcFm5bWx+M00hvwS4U0zoYmvcncwVQ7C+uCkQW1+mwcUNtSh7Uajw
k+yfn+AYCGVuBs3bVLV2s671frsev0qRTbrnnm+J6ogWsf7IuqFs6em1BdNqeUGg
gLRLl7Hq4AkbpMb9dvb899w1zxuVjq4ClMjKJDX9Y1kBldH4QMKbnUFTXu9dxwaF
6JJ41oc1qfAfW7E6tP/Tk1xbxJB+5ot9dcQR4F4pMy9ql0+L0S1BepvZuRsUWFBT
0Gz002YHIti+V33r2RD73MdBnzcEQWaehK2qFD5FBggJ4WMHTrz6wsHoO2+YAW+L
EMDYmodE0q4FdmWDZJScRZzB/DbLkMNRRuOycF/BJKOKrVoqiXOpE0H5204phw1Y
wROA64n84flqwTwrKBq6kSMu3NxPKevFwAfQm1NC9HEmRKPUwmGnxiW1/y736tsi
AvmO2RJKlMylvA1qqvkI0DrqFNznbN6cFZR6mukK/qUDBvsdxpyLrD7igCR8nWq3
Cqhv/EXA8zyK9XDobZG3uRQXKGBLeDBigbI3uRNxEPgnqiveouErhYJuesmxxVZT
HYNfr7k9Pq1NxdPg17emlE5z3VjVAF09Vx1ygjecR0g5tXzMOxHaBaQlelF4Z9rp
YBhuZpfV2XHRAgt+Uu0aww0cvfnRuyWTmiVh1C1773DV2ZrTB7qLrvyWXCTjfbww
/qHE4/AdGQdRjRovrxinhge0xKEsuHWdIVwiSxBUFKQULDb7leZckoINieZh1DAV
roFWpWFEadKLNjAt6qg9hV9ZnOcAa3K1bWsgN+UKB46w60hRflme0twAjHx5viNT
kuXfOuWiwvqQjPXHzxY2qM5vnHBI4fQIMbHp5O9B0lb13GBXeDm5Gamq8L8Jy3/l
ee3NlHG673leJmZxWKziPd611GMIYohE+csHGRh2/6edQ+bezh0uGwduJMjc8vbG
Dd6AZSM5pZOeDwxANFTczo04roCe2wqDfAJNoJSHrj4CyNXryy0v+IISOZzrCCAY
aciOz7IgfuBcgyDWErP4luO37/q2f0jYrBeuZaCGpNuSb1LRMfCBMiEK/0PnDNNz
+lOzVXODViFVdNfdA2znXo4Pkm6Wp6EeFcrz6L8Z0nhp0jRfR0xA5W+YwvPWHjyk
guTksBSOdeJ8U8PWF2YRdRO6dcZsRl3IAsiQqtUmTY3NeWjn+sXetVchw2klDRlB
jMXpX+o4GkntyVS802y/CvcQnyZlm39GvHU0qrvAGaDUdAafbiesa5atzT6LFLa2
XyHmmlTmvM8fY4aEcIu1IIcnULL7SkFFP69aMdAbDVzWkRmIJlmv4ovzm3d+8HAM
hV6+3tz0qt7WfKk9BC3n2IZr52wo1SJ44MZZBJExSOmLToonAzyc00a2xyvd7kCq
J+IIiHCpUdTplcTSY33DvPJomBTqoI4um8krKc14X0fkbP60RLaBNYj06nD3iZZo
d9viG8K0x20Katyh+WoBo/iKshcRrGWofJkO/cDXWCwC/H5/mytrsX21HacPAkYs
xZQmUqoNfCyx/JtqzMerZdDftKGMA9az6cIcBfCemXBPSR2yJ3aHSw6C+jbbyUhT
TfyRKxLhOcOGOnnpmN1CTcUVaGIW5Dx+LPtlwr1WYp3wuSUWOUbgTz2i/cZSwse/
kIxvdpeQqeM5wvXZl2e7qlABSr0+XomBnGDKvXUGq1vHMoj01elIwFzW0tLwMgK9
lqYWAorWOwIkucFt0AI99cznA9NiSSqeBbT7HMwQck8djk5+nhvEMIx0wluvGJDl
aXZk7L5o7IqMUNoLrSbdh6xPk266GqMx3w2kvnn8HOis/Yd+rqxDFU7hVAspJq1l
iSmYx1PkIz7MCi60zE86dGyhjjykdUXeY0Jmk7deVrpO8m4k+1WlcIqgG4563GZK
3RGLFJlggl8spYz+Z2OcvF9YWt9OkhhBIo8HRSsrCPemyLN5GRGjI9fYFn0AVzxu
thCOktRBhGESptBmQn545iOZe8g8G0D1Ichg6cvEzs5P1Wfu95lxx3aiSF/QIx6t
cBf5ZC1q4YIwY+n4GiXUpqZbdEmwZAZv/Mz7XQUsw9tPhldJXs6C76hxy+RMk/4f
zLCdzfJWH9OJ3fy5ScGTcZQweDUVczI3sGkNZF9e9/ChcVpdLuHH2aE7/oSBttfQ
ZB9N6F8QO15ieb7orwQOobT5ciI41W7XsjEbj0ueVNUHJI+2SBuWRtY8ir2/WTqO
pP6ZCkE6K2xGd1DtXxd+tjR+xzoBct2H4IU19MuuWopETlXslJPIB5Jnz9gDKsK4
DSTiPjPbgN/ojBrhVz+ywWxXmWHGG69xbD6hhkoG70P3ZTyqOLhEcNy6nzJCMoUP
6ET++bSLaCfzX50UWoOStkoUM+Ett2O3578Oldp5k4b+AghUH/a+Kg4R/wCw6lvP
E3BYVpLfUIxBL0JB5rPvtrFIWTuY0VOGdxrNMFqQSYG/bdLgVpCvQxXJYbkbTEfl
50vcfGRv+f65ES+RdAS+pQFYbbruywQ7TX8nE6B5bJZ6ASoladc7JZkuRR5Fk0Rf
lFeOLMNv0HY/VtdojRGB2u2bRBaWm0LEmE140FEoCtHNFb30I+ZpHkSoVko9mvQ4
prPOfe6Pm9KQ3jKOhkt4+mI17H7jr60X4oKx3XzquZhl2LEv5GAnMANddsU5O75F
DQM1sLjcPXb+6NlCX+m6H5/l8b6Kw2kqXpe4BAm/Y1680zANoQzGaUpztg50O9ai
lc5/doDg3Jyg+lni5LvZauNkpK460NrjlsNRbbw2fQ5ggT0+lJ1ni7VGw3ihOfbx
djrCED5XWOmlAy1OAO2B4RmuNKlesPGw30Yw2tIZG9MKymijNKaJw6AVY3p44MV9
z8NDpe9s9gDrQAe44JmcmDiSD9vVB4eRrypzRlYiA8ionOM3G+cD8nGGczWIKOLz
JzAL/6vQjcE87kCaZgAcJp7TuARJ2927mIbuWZi0oFybyuRuhzkbCLSKS+bpEeCt
TQ2LZ4cJXd20lsgCAycwWU4nrDWmCFXKk19iPUlWn59ssd3t+4+fgYVaQ8+4O1sc
9Ys6sp7jACE05H8f8CJ7ZWWP/gO2a5lv0cg9X+mRt3GcmnCLnfHsidWW4TdScvQT
CGQKkafqVDHp0WmDHQbAuer1Jw9VF3xqhirWjo4ryTFSJJMN3jV8nClxpVIsUIPp
7gDMDh1BBRvPlGO+XfIMCnykZVozIiVUHw+eB+2fYffJkHarqarmQWtm+gIYYkJr
xf/wdaULrFei0R60CvfruRxODYL20NXC3/2JOkLioqcb6C6jrqsoDrW+Eme4l11y
wdwMLlYt6xzt8wQdCtPndjehbOe8Uq/3Y762hdjxGMRG13t6iMClUlHpGn8pLuEb
LDGHlcd+kB3nyW3G+6/L8yF/Y4dl3YTyeEAjMPfqR5u5Q0Lc3yCSPbHP3XRqhNFB
UTvSMWIdDsrgYE/xRJ+3ogvEtUbaRB+hMIh/pKmgZ187tgXG9/hQqapDngKKtEBl
BYil13aPGJ3AeN5mNaXzm0HWTZY7tXQJnpQk3A3GuGI0DB6ShgaDIdP/FzRUTHjN
lRpeIUoxGCKSbMmaSbWt+9bKn+z99DSoePUQs/W+GIKw8jyeG25F+02zhrbk0CoG
KldqkM+fR8GnJE8OvQ/jRWg++l+KfViKUb3Hp5mIHdBCdSjvAJ+pVjh+1FGQwfr/
MF75x5YT/umvFJQHvSNyrTORa9amx4J5ekWVkeIhsvKL+RTg3Bp2xR5WfP6xkg1y
ysDBQq6b53FmOqpPJm73tfzUxN5gU6WHdIM9807CL3rUpTdhaiHOYZ+NmeUL59DA
IU054fd3RVVWeENnNw07m9IKWnNzqjzls2k/5FuWH3CyDzPyo4yga7KtylV2513W
0R0j7MjhQ/HeSAl8ihow/2HmnZz+jKihqgcMv9odPDJfPKphgmsm849vI7SbKcjS
mmOWkOyDCuJ7D01IsqDn/KB4wOK86rBtma/j8l+wxQKXqw9ARXa2FSRafEBZR+YK
U0+OENC0c1W98nR2pmzVxjII/YM/453D76odkM9LaKgiEvY423b/Dqe6U1blSJhw
gwxzmE2w4cXch1HmGp5r4V59OIe5CCTJ8GkPBiRt1GeVGIhpxGmlSQxPSg8Qr6Jw
phdOr27sb1KR4H+rcYfLkkO+C1IgMWOgBJ3EXjVzPA20wb9J5ZfLSq56CO+HTQb3
Dxuz/B0sn6+wKyR4cBAwpw1E9K6p94wvJEBpzs23M+tH3OUCps+eRk3dQma65MBN
zwvXS0gkrEbKjgODQRuUj/rATlFV5xHqcEI10buaw2R57g1WLUpy84UEBxNSOVTe
Tk3yujZwDCrrKw9sp9ePP+w2XpRAQXJbO6BeYVxIxjiJG4FC6Ruh9Cc1j/A1Z/pT
NeunDiazpXELvqKT01bykJ4A8TGopmbPrrJFuhJWUmbj7D39itk0P1JDvH/HzYjg
A9QwJBifKwNOdj4kCbvQEKFdPuQn4lBDg5wtR5QBWncuGx2tOXpy4nDrDHVhz2ht
Ge/4DHDYxoOA9vc0yCCsntInUbFlDgoTYHX5g5l4VKsLnfFoMcX7PamX47qR2tSA
LeVz/uL3Sa4i9INFtgM1nBAXyTBwrm+d79DqhMM/nFec4piblRGNdo2q3HTVhiiA
Xe/Lj3mIbyfKt/frGxgOKstfojWsxIHeYGbYCLYst5tTJRLfrZHddUQhcp/mvtk/
tZdMpXT/qPNBMV7wQYxRlbkJENg0EI2EZRDB+QpIFPTJp0AlPcCsscauuN1QIPTl
xFYerWhq+3uwzgZeEPCixk1pfATS7WGcp38VK8FtrfInDIs9UpleTZb2k4r/LVzE
+T99LCeTJ0/LUoppoOQ1H5Sj0haVQ/nYp5TeGWKi8PxDcsLkX4BvmaY+yq66C+lr
C+K+a3DQNIbzkuvSVe6DX3CA2VtzNTKQApSmzmvydujy2OwOmOLzjycuXk5Q2R29
DiA0w1R50MfuboSz+bhcXMhSBEOxvj9t2qHAZS20Tf08HHbstWe2QLE/Q5QHw69J
oZ7pLqUH4myc3WOH9hEGHE0rEmnk+6PJCxg3naeXW4NBTWmUawCoU/ZgOWFugrmX
RYMEGbaBGyjIcYP/Eak0Q/5xj3BhsAEKLy1jt9Zh1Av92PXjWjezyFB+EbSDF9Qd
rjV98+2kKNjEykQ4J/Mhk2uVvVKDHwqkRoTQWlGRjbyqMQ+ILqgwj2gUwLUk60VL
3U+qICZlz8wPQJpeEwTMmrHZZv8J0loo6zb7BvTUMWE8TQjqVLV5K4VPRMbPV4t+
PA2YzE//pPKn68LIJ8bqYA2ZFP25bGWZ2Yrk+H67cxoDYkjMbInVr4LyBxKeqxVz
td4QCuQZZkcN1a2iNI+TdgRcR5/MylE4BbwwcNq5U7EBPHPk2gcgGyAsf7N3d+HT
cwUMKtaN5+cWrTasX3RKuQeG23IkkoCMbc5s0Ofm7HPScYMn8p/rVRltRn3zSwi3
+CKyuT131mRdbudHNJK+W+lDM1XNVJhbUuAJXxmpfzSUgayZWkjAlAi8i6XllYHQ
rCDrAyBiKuAbAzD7r1KRHWYymc6QHL9VKB33rjRi/b+6zj6TNmeFKGWEXrdUPk6d
AGHW6pDd4T1uzJ6ejO/biBk9CtmQSH2L2j8O/usZh/hebciNKIc7gpPmX/tkd7/C
v+XxKELGTjkkFvMhWCyMYULCQySTx9BbDFWsQVYXyYNwjb+r4GI4L4bQx2+ew2b1
Ms9niGjPvoBhCKmbi2b6p2Saw+sLRZYro/jtNMV6DXsA9kCKKNdwsD0bLDvpzVpm
rrWVmXxxupftmpilRP3eHTzjd4ms5gn8EL/DjYPoKt5Sm9uVqKrjNFEJKkqW6c7T
7NTl9uOSZLDN9tqOU70hzIRvLQC8M8dn4tDH/zFbejU5ZmNtS5iYS67MFGpZ6w0v
yVLOQSG27kzt0nZqfD09Bw8YGLtA4O02wzw1N6XCiYc+dsnOFId4w45hAucqSN9z
GlYJp6SzeVg3PmtToSE5FH5fFqR5tjd5DgErWLn2pWLK7/6QgazZZX7nx5QdhJWJ
I1bjuFpFKudP3/KiUEfbC3c28cXZ/AbvZhAiMILyAVjhwbFycC4OS9mmwKdkjYKy
IzOfIou5z+KYjL7CrXcEW74GvKytnTFcd/7qz8lLMtx7MsMrV9PEAfJiP4s9Fyy7
YbHjqKBqcqfHdV+Marf8BHJ/drqWGOgyM3nF3PkS5ryITO/S9+3gyRGb9GcKg5e6
0sA/KLG7tHx2cxLl4AAHdXdT3yiiGNt7vIT5MA1dUJaelL7IEJPd6FZ1RmhACiTi
N024yYsoVtu3/rRPA+jH0Ki19eC2lbxu/4NYE4HlnhKjriN6hjyCd+qcFju35Q+V
iuzMogG31QqQqojUeHG5Bq/dI1Ir0A96IhH39bNxiY8U0pZixB//yd+Njl9ek6Ll
0r6Lnc1oKBvhLe3/MGelg7oYob2Y13GUJkSoFH0u8b2qmVeVIT1RtvV5bbsrYRMB
mH+IF4LnYiYweKb30xA0/iUcMpV0TkG6HrfmZcXuWGE1tzOByFmv1st6/wDrjMLq
PVkR4tZEs4vpmr3pED3D0sbd0Rz9WVXv2Uts3vGPjcI7WpMtLs0nkK5lU58bOba4
Qkdjaj+ESTCxllGlxXt4RKoxuRrWdN9wUZmKMoDMstTGQmFl/6qimr97izJglUKe
b0VwvjaVh8WXoGDjzMCO5yHEFcfP5M5DCQwJFp9k8d+e2Qze/Rj1j0HYWUCCpGNM
ZJOKTfE5EaBUV1uqufBjEnV/PTngt54YuipUuGCeu5bnlZgMxewcOxCSru0WQj+P
sLigzeooP/+G32hWS8QN87Cqoo/ONWSIpr7l481MZaLJg89qHd3zsfaQjmsiWt3S
WfiAuBcWPXan46ndpFpIovdXpRuV7o6/m8PqugqtOB+dsqs21P6euXBVw4l+YaHW
bA2d4EqEFVpgrMi4b/lkhdt1Wq2zk0R9USnfddBidov2q9ndWBu+v0IhHIhvRk0W
NGZ8k5P0qqCVOK8BjpY8JvdBc+61k6bESHpqlr2v/CKthXK6xHq6sMiVg0mpjMC3
3QyS8w+LlIX3q138KaYpGkl5gZKr6/wjKjEd27Y7C5NT25YkMK9D4LXigzNwpPxl
Az9fVDRFVF5qxk9QtjsvPlfAHmUYoRJk+8KWnSCt2jeoGt2bYZ6IjJHYgEFrTmzo
YdAf8ItcriOlSBPYbYPMtGPFyro7dQFTuRxp5SZTvB1lqizEeNlAALlvjby76M7f
OPNaZ4ccze5zYPgb4zzdC3q7lvdAPZRJC4EeJ4ylSTypRDqWrFN2Ot4Hupr6M3bS
d6qAJE57KXjGsgmnCaiaE2awgT7C8lt0u17Gh8ZP7NavgGBKw0g3Rnr67kV24irB
AVbRd03XVZH0V+xQDDINgmaSIOhAL0QmnK49cVoszkzSCmBi6eOQNVOSCEVV1ASi
3YsJONlMkME3V1Mo890XYfeI5zV4bG8nYOb9hJNsKmxfAeV8Ge9dtYOFJ8qTZ73J
KmkrRS8/A87bYAYadh5Dd2uayRUPDr6Sv6KRa5WKKwszpA2SATYqtDMclJFcryP6
O420Y+4r+eAgNPOvTi2u9nwmHkADqx+xAXpRWaB8o7y8RjlX7riGYv4oFgH0RNqi
aLkIzr9lOKr+1VrurhnUZDN087tIxDT4KXk525r+9Nk2lIYYO+K9/O4o6PS73Qbl
tXdHqXJnmqujgm4S1WY62nooZcxtz8WhabyHVZmuYALBmHf+VR3Zyg26chaNuld8
yndBwrkRnNdQvGQT1RL65o2FAntLaTWFyDiIXqE/O0GPlFBmzG59t1CIq6lW0knF
Ee9pkPLWf87XMJPSNj2FwkRE+pM1bys0lZTdASOdIk3qZufU7FdJqfzp+QVzv29z
F2Qfw4w6sivVPkq02YDP5N8qjlN3dE+Lb+YARtXmMU5uvb3WHcyDzdcGNVD1orp+
0MO/ZwjDtWAdc+C+jDE8T2z7NqXpsdrVYvaEeeNLnEB+3EVL9idFRk3mLTC68kGD
n2JG5ew9s5UI0e1DdvatrhOGdrTER9NMD1w9FXEjeIHyojVOe5IMLbaI0XzbXjyV
l8F/HMPiY1ZyulnpqZJ4/VEaZb+5ido7ovtc2kYE8hn6wvQJNbl3g0K1KCrdgKt7
f8lZzpnLLSescFrTVbGTnFUx/te3FFIw6y3rD/lfw/Jy12Mv/i2D11t0dVIMNAR3
jwANs7ms/dVjewcnlznSIJYxUXIsYsTMEaw1TjEIGOBICe1caT2dMtT1CDXSRwDO
7WWn5TonepnWsnb2dfU7PrulrFNu6A41juvzmszlnuGVQbPI9LuZjQzK98WgFFbH
zCTj4qoPw4cRb8ekfFY+1IL6XB7PW4tduHlfjFGjJd3Sr6cdB4fKF6S6vG4hOBu9
v2cOB/cquFNR1R7X2oaL+W+lrY8p5T7txr5+rHA2DUH7T2mfBBMvrMRWs4QMInQe
VMl77mZZXWsuPjDt757o//R9CtUnm88M0b6IjWxJ+QnHL1WxyfPhpcqU4tb7+prz
Y5tJ2YIvDt8Z0ajWda99SibV10bPqnVzDJr6zC28O4M5+AWwtl1Ry/g20aPSZo9n
mCmzpaS5lDatRTJZ0EtbkCc29627CdZYUOId0NuOInj24qpStOiQmuS8kI3Bcz2j
0OYOh4iFeAyl3E/+vpacsDD6Y7e+/i4AJHf0qBxiaYwDtN4sfEpPXDw0LrqAi5WU
7PF0xZd14u7aejHFRS5Ekg04uhekSFozg8i2yLD3MI+uUSRUOrmK3CvNum0q8e51
3H1NaQb/NvbAyiDAiN4rZYZP7LD8Mfe9IUsTSgJfu6+R5gu7Cxc/S0VUnsG/DZOa
OIicx4zx1wI+rTwOSo8wjlSNNdEX3cBnYLk0z/Mr36LF+a1I+MYnxslabhhOwr0/
JrnOwlrD/2+IylMODrlpKCBUskPzJoQh9Zu8C7vo7vfOsorX3JWVCWTCyG2UW0GP
8bkm4slOWen23M4HHlF34niAn7yopGjYU5rJpK2jg/38bKlzYzMzyvNWhmYk0Uzi
hR40TYRdKS4f70u4yntglPl3W3XTUb4fMloaNxVXSyNAmYRogoMKZyxFZudstlPK
1e0PQDII4FLlCLArMXsIbJFuLPeWMfnzAveoeIxFu4BveHsYeobx75bXuXXh3sXr
ydryyVr9zVMKp0ieL0Qm2tUsxR0kMBtG+nDOaVj/vtXS3ZkiCgRW+BQrD//LN+0d
0IdKfnixI9D/MnNkDchrMlUnUOHzs8jqrEIg9gp2yO+WG4CQhxux3V1wLmSh9jW2
mWZ6n+KMzeFLd2rxfQh3QUf5NEg/O8LqEImsQblzRPA7yGLeGCjRfFL+btDXad8Z
omUJs1MqnyZKvPMoOjLlJhyOcPL+DnYAeX7CpQg19lnWFHktF6uO2o9daWD4+BYq
qfppVX7yHpXiqx7pvwKRre/vAktoGZn/BYIgJr+MdqldYaHmGAS61c08I9kcmAxl
dw38aGxWpo0FDT8eUAtqEn0226bSq/nCz8BuTpZevbtILtqmRT2cG75oUaTZBjan
tI5oYvocehpOxGSQjqHIfmx/IOqI4+ZPmpd9EsMD14Ss7JMSLD6AfN0lsnZkG9cg
V/HX3vBOX2VAhtEeG7CSMVmDhvrgB2t0nvMPVvfmp5yrSfV9mdRs2XqwtwRFu6Le
SK2YiTodlZ1WINdiExz4hi+dlZOihL7QzBBYIOMZIkXreY1VWwn8g6m+tCvTpw84
83FiJwM068oEj6HsoHaiBfnDRzMIrGslJ9bqXmKpbLHfPJA8CyDs8N1oWFf51qiD
N0bO91lifmDRqj0UrCnTjBN30a3MzKDkDfI+JZlmVDOGJjCt4kmaW0PHrRWlsJRl
ONG8sq8UaSIDp9u3abHHEnIEjC/qb7IOmBwjLc/3DDwZgiS+FKujtJkbpPkKnNET
hLQgOAzpcLWE4W0UY6vKQV07KlkmO6uWG3upSKFbx9Ss2di+JNof6mTpnOe5cPu4
IK9CLkH98nktTJKoGxJlxI4akhy8ln97fpB2NTCrIHbRSvo8aPtSeL6jOhN2JaC9
h44HMg6tapGVnp3a+JIEY5ph8dZRhGzYhMwx09xsFdyZ+RLlZnZzNlkdGRHLWsMY
OQ/hKPbN/98xe3BzjX4Z1HqdccSPsYtGNJmCQTLY7IrGAmjafhHWSpvmp9NhpPJG
ycKuSVa+eucwk+t/icXRqOhytrNDMEJq9vnL6Sz9x67Ty/mQrfLu50cPgcfx57qx
9hvg/qqyTooB2Qw97JafwN2U+hNjFHa8ALoJOc417pizxFXQAkBAH9JZAxcQoNKx
3Fdve+7K3A4eCaHFBj3aNstl7RuFHnbPUkM9EWQ+638/zuw9DCewTg6fYBBh9qTw
5rNkL3kxOvQIVpW9KFcugOTUzn+cZNamR8eYChccawpLnJOn8cYNZPI4UV4PF5Gj
Gi3MbbHO1HXpuUVThuul4iBofM1h3GNn43V9T1hE7tUUM1dyg6090hobcs7muP9e
s9dhrTkMRSjzvMQACdyF3ILJ+xui66M5s0qCKh/tLCC8QaBsRJOFzAvlDhGkClcD
30Eu8v94/xUMFRmxC8r+Et5EkSYVZcGpoYn3XvUize630rMhpCTcSNLye0DL40/L
j8lZ+FJxb48hXTNXemWTOBuZIQ4w7k/C+Cm9qY2Xxynxeo9P+gIyYrDCbHrl1zaa
JzHW2ze/zVZhGbqCDHat8YqahAIlpdS5ndxl3364OeohfibmYSBuIi1gBYA4PNGU
kkw/6/sl/q9naWGpUrCwGw9lEJkHrhCJbQZob9WYxh66OR2fuscftomgEqEr/7ZS
nFIF0+zO7n4PvANsfgNJmGJIou7WbUMlOqHzjcv3ZactpbFh9apGYgOb71rPYKtu
s8fA9m4Lyskn8GEi+vj1H86Y9OaopSmoEgjDK3Btuux6lT/fnBkkcBqa8CMCjv/Z
xb5CK358tml/Ww3gWKAJi0ObGL93RjL43b3FGpf4PWclsaPMqQcF9w1KnwcjVq/O
wk9zn2tI2cXEJrKrUqH0T4uoKvw0f+Y57CheqfcCi9Fq0QHj7Fq2k4/8kv57GfZm
v3Hpylg3dG1Ie5p2nhI8BBC+lqJYMxax4dtj0ejj1R8/hsaclFsI3nBUWALckqxO
ZKYgfR/OnyB4gzq4n106uaj0531c/O8mrdMpNA9kkyMH9FA+GAYiexpkw+i35Vvf
h9Dwxf1Vnw8xp6Ip427BwxT/DXFfM6no4BneGWCTGnG/Uq7IuLLgOV4J1OJy9GCY
SnnT5+51LenldQ6Ni5E2fEnM7ODnSbWYPalcQLTSDzc0LZ6nqeDc70vqoDEOoQxG
V16mCayNzoEjZ/ncreMw906kr98YpH1XFJxLbCa6m75+AY6+Ab/M34lx8DUk2OYm
KyjHQhJ6msFbjt/wtqhbPq0LgpKqpaIpTxCBFnLV28ZaxyuyRj3wcu495Y6v4JVY
vKDjoVAgyyD5kMf9Ng+Phoqw1PonH41w+nvu5d/jOdJ8bNa+bQaQIFTfZ4J9qMbn
gtWT0uXIIS9u97AUWSXUsba/ysQHaUbSswz5s9o0GJnMWAAXvmZPq9slxQWSfgxY
8b/QTZYWRG1uKInqaA8JcmwPzGNizWYZ0E1Tsu4Y0i+SmeW1+YFg7hOAvos2WUYG
8AEoHJg0R5Qp6MTjciRTzybrc0GKLemBohgVd5WmLxboI/WdysNeYacE7DO+PNvG
hd6uWQCzmsZDtIvo+2Ne3bmtIiaSGlqUoykaV7t8tY6GxzB3Ml+Vlv+6dtK1ycIS
D9I04rFaDX/fVtH8qSrQVW2w2T69AHCTQ2Rd9woMGliRTk2RsLOn+Q5nCmNb2ZH+
vYn9k7PatuYJ30T4wN6SLpMRhm7DVC6Ggsf5BZg3XAokFZURFplOahFyQcNSsHS1
1RZJMOIbWZsYMBM2JbmFIBXQy2NqGlwBRMPmDtaZHo18WeHmL/5RoYCSdf7fGMZQ
ZqayM/QMoPmwuaOePL85RqXBSpmdwSLDeyeYovKboPMvWijj6Ol+1X8Wm/wuQ9rP
e89k8mU2HWJJH0qz6vjrmSedeU888qWqZphsqKyYnhCLHQUeh834re3zlkw7C+Dw
luZJuIFGUqOvBl8bdkJ9b0wxJypYB6I5MteNOb1c/BIsKtsiRhAqSYSCGdesrkZ3
pxVga2pvdYNkVIbcad80bgeug71efAYU81KQV4h+RcoI53WvbFIqhpV2t85tRc54
Drz0AyuvtnaXFcTfgLtrCEIA3aDNf+v/9Hk9X5GIjJ0Wut/ibo6M3XXPF9xoqrmF
+XsswnXZqN1looz0fbi6nbWR78Z9sqlafNIIjuTby9aEbKUlRuJF4ptv4l47CoHD
cT3wH/MceQSkuliyGBIkffRncm3Fvw4iJ2IZPA36D8dcYgwhyrMugZrksm6hS/Jq
dnbSojEiqpMHcHmqyMm1kSaMMOktE0q2re6kPP0YXgvAhcmo5ZVDT1gE9JKSl4hH
JJr8inRAH0MJNEJiuijqihph/n53ttn6bFkNvcOQiXlkR2uz1P54l1hms3ecAxcI
TiYQ+CejxDARS67H9JvPyqGZsNInb2WnONj1W+G7zvxmy85QwVvtQDL7x9JSVr/P
MejRR7HTGaoz2vY22BzRecmpHMGSdTnSM8UIlIBA1srODvw0NBSaoiBmTGgYMuKV
Niog512khzJiBKYIt08E83hHHpqpPRC4n103C270+JOV6Xi+hhyezjBEc2oyiRj6
dYE5VxqZo+dY3avD/vBBX/dG4nrhNP30OUlKmEqApcNrtzs5yhv86imm7x8ZfnDd
InnkUuWM3F5C94hjPe4NGzHVudGfXRrs5MOxnPnlRxoDrzDJSkwdDj0FoYaKnC7o
UbuOm6rBmDBiwTG+Z9YfkSZ5EwZF6fljm4k03GmUoNnLtwcAiIklbjoEUalctVN+
+2UiDvZht6Ks2guTwE9g/EW2H4h6nWQ7MM1ChNSlNwDQVso/suQY5r6+AXrHVTKT
OSOqrXINGWbnHwh9u15r9FcpYt4JsGBXVhPItb+jExqwYrrsJHRmpZch8emoTUbh
rvloLczodW6MRDcY2/MWGUyuo35JSWiTmSrYoUr/M8wHLP6syNtCabCX37m4bCV7
Ezk2tw5KQraWMMERkKTmrS4ROydTHou3mZkmE2KzDSYxctkNHct55sPNKyAkBUNW
+TfYfn0pHd1RbFK+zFOchnCqS4D7DfVL47KupJoyKApLmJDlp385YONozfy6i2Hd
38bClT++wOjRkrTj37PGtjnYmOOY1JMN+7gPQQzS22B7MjGKf9zX6K/iUoZ//m4I
EV8RasRTHPmqlYdRQPRC3v6PrgwSDzaSOOotstBx64g0MGaoqeYwhVEaN3XS36Ad
Bqw4xTsXH6p8zuF0bHAdBL2DXLLg2RdbE9U8dzZ0buBuwuM3tR1hfiC+B9zuGFLY
tfmrGfLURutDxJ6aR5pz+2j2lljRITUMe/WQii0FmgBbeswP+mJnHJvGJSnJet6b
O4Fv8reai+7pRSKhTAj4U3oKG1X27zjjV0FGC38QrnO6YrPCc7gcYVexwpgmwVVs
hSyovuZIXe1BWco88WX5wXYDIe9DdQGMehmYkY+P5/Ei1puF72TISSa9yX97BPcn
+RgQG2bJ3YH833ou5NEAWPAuznWuR3NDL5/8rpgHkH7kveryJbBPyeeCbZpYSePU
I5CyBDrMMeNTrRlhvavOW/gwfFR781XaIDBasH3+PZsan5CX5vHWaTJGumPtUxyn
WW/Cv4ZIVtCqOokIypxvZUfP+9FSNd57ohqUIutgxOduaC26l5H0dkWc/w7eiDtm
Sza99ONMMuLgFN134BQAc8DAN2bCv2DXBhhKY5B0k8078TIiBuypVloO77AmEE8D
4dXikdA8VwPe8LwVXY7Ftmy863ODEj5KCFbfo9C/+nAaAhr7rQnVSq2sOIHQAL/G
xWMSXIwwizu5FbrNDPa28EQeovEE+U5+0xKTFvN962zhl9lrO0v/PZcRz7ssQo9J
w4Bw0mrkSDdUz6iAdG+5fhMm79KlI8dmO0eyH2Tdp3bYh4a9CQ7L+L80QDg4s4lX
eqTQx72YqXarbA4FC3JeKajn1WHQiX/c32g1o4anDFHAoGoGBggmxG9DhD3k2dQ2
BK4Vwlu8GCpwAP2X5Icsl5dMKW0lt7ibyMV+hvs+U/6JV4JIwRE/GcfWk28/EqJC
VMDW6o/C3CUrWWaij9sw3a8Fvn/nZVOBw/IEFkYLSWQzPjAfFpUOrjZ0yOMuLOR/
G0ky1J3dJb8sMDE03xVHq7V3EbsOryovR1uejo3G4dEfiIW5doNg9kV70lOIbu4H
dpZO447GFG3JxcqIihj44oHUmqcSDa/IfXngG4KH9cLmQQmmGKvwiXVn6Tcu9Cwb
eK79YF0DXq/RR0WwBh3Wvls2/eX3k0O87eWFZe6YXjUPdhySRc/nvN/sBTQn+9aK
yToAqbB6O8my9T3ZPzhMEBiLC/3tttY5bhU8nB8OWtO6zjB2BAlgXD4XWIMOU3jY
fODAfPUNJT9vmWoHZDVtGpr6e6aRxPpVauXbO+CWblNr+jV5xe5+34DlXycX0CvV
KYEgkko6gCTm3hh992meAp3cQC0FI9uVhUU+Jts7Q65Ks6Eo9AVWXde+zXEfJnfQ
E8SrIbJndS+6h7M7Z/c7YW0pNYL86o7cYq3Wj34l60BFhse0Xtv3xpXxz3BLxSXH
X9bnUZ2cw9AtFD6JFARZsEp/dZAgBDhNIjzweEVutcoRtxjB3DIgpGIB8wrA5l99
qdxdtYOfIl2TXYomfhA0w2JGPET862RILVuhvY4ktvHHR88iwIFDonxJM+Y++CHy
IPxuL5CutITsDIjRRfaVoYBHxKWnqJcNZVnswWwsdrBUCQ71wI34bWU62MDg880s
VyWWDlKmEHlQ3l4L81CFkzN8CRM1cg1GruLNdjSKgSm/AwIWyVAGr9bkMshZ62dK
PMXufuTkkfTuP5rV90QWiqVxpwKgNjJ3bxHqDaG0GZ+5LJDUAb/+VNnNb2JF/ERu
H05VtFRSVAO+vMiiAJ5yWjXpV1JNxfEAh6ZYwKj2taQ6wj+B95+twLIYpsmhxbej
krhRK1D/TRmDz6VFe1Z5wYuSkz/GdNolvVGsf3gpEsuGYauUKMcPk2rc13BgvmyI
lBasFVx3Kp8bGAgudTSEyr7aT4ejIsVFQDaY7QrPD6HlgH3qo/m94hTJjG7oLIfC
ZVQzQhLagKXPnOYZCx/3xRoVHJ+ZPjGrQb1ClpJmxqzsltvH4vn46Wxpbmn+ZIMi
uh8vYKnfQHEawZ8pCHsm3xCZ05lFP1/ous9FsPYBJTDhRG9hagzlty9DNbvAXXRk
SgEGhMAEGt9GKjvNgzW/kvZHhMhqzSL0bjfcyAp2BYJps6lYYXvG/w75aCJOtI4N
FvnFV49HRUvzRf4G8AQvlVpMP7rZGRAKQyCCKa0eivtLkwmdrkeKpH55bgvpyH5p
NJb64g0Wqp4U74U6yJ0L3dJn6KvoWkNbXlgYsMZMUH72u5aSDAXa7fzhVePnrh/k
fZt1X6z4q0nnk4MQia8FEDBzN8kKFT+79iTfqN7dbuS2vNW+94nIwrti0irIQ4x8
0pgOVZKF/1K427cINoJn9L4kVu342KEtiGLlsbHeSOW8us0jFCTEDfckeu6L44ny
T1+kSp8koUQFUyhEE+lIufgNCele8EPxuzdLePNKMEMA3tCXvXW0WxSQ5SELq9lq
z8qKvke3HZKEbE0CVoHxBDrKReJvo0/EZuXXQQPcInU4FjE52oY0kitMvSB3LHQV
gaOlXWcD37jXmdNT7snyD3ozHBKmuAxsnsA9rQhRP541U6dCBo5cSB/L9nZlymEQ
ZOGCSHEokSQkCYINaGJBCV/vfGbYBYddjbQ/+veqVTI+PyYcc6bP/6NP5p5DYIfG
5XRQDsqXZGb3KXtVYf+WMJqup6SynS27MKYWu8HqWMivyk9coOmCIA4D7i4BVF/2
4ynt0xCYzXaVHSi2vS7XcCktxZgc0xeD3COqMWbY33xQBPjwgNcEtxNep+prCrAR
PVn0E2Vi0wsgYzsLSsjw1HuZF5kRxAxO091HN+UjBirv2iJxNeY+IOM/84feNOc/
Yt6SZafTFVlfADNI7TweGZ6gXr8WDpcHX6aOCXQzA16U9jkfMdFjv9EV4STEKT7I
XbluHVnNDt046BJB7hUpwDjkZc93T1kYkPyr/2GWYpqm3NS+FJMZWilcA7PRPNOQ
oYdEWyM6fJHtM9diGEmL5kWleYnirLMc4pSHv7lR8CmIuV1P1Olc2SbMpdfgV2EH
HzvuD9QtZdyYOJ48YaqcDgGe2Xp5lNA9RKOUcC65kkfzR/vil1IjVpgHWbmWnAZS
sP57Mw0ImGjeT4kuB2O1JOVDQW+JZwQ4tbMXLkk0/yMwiwcIEpswd06hfzYi8UcC
T9/Cpu4LoEeZ6P/KtWexMHl79E1lf6LV2dttRYMKkSqTJhPSnkgvMmdP7MRvxiqz
31t8UABZABoEKwbtu8E4f7GZDXkaObqJzkxVTwcS78E5rbJCSbL9tlgRof5EW+2q
LS8AC/nsAU0SFw5y14ZUDP2FPIOKvGc9EoaUMQYhgyM4DtVVSbY/UhKuX1z9X3zW
xO9e8ftm/c9elW75w8aIL3db5q8rRIlpmwxsJ/xPXLqEaay18K1VjOvQZffXo9ms
SdzqQRaRzspmemyQCge0GApF/C0Q0k8XO97gAoKcDkW/ZwgTRr+IGPj3nYl29ZPp
nDhtG67mLuYr7hyQOCpXGQ1NiGZz0/HscFEKyo5CO6/pVR/U5S5tNDf1oC4GXcas
7/96HrzjQ4yKM725r5dWMhrvZWEtdqgd1WoYVTPWIsiBJ2TPBiTyo+v9wNAXKAdG
FLJr2rGrAElYq8VXrWUbInbs9RTIjOTK+Q7rk4E58A+liicM88Rf/CDX8F1Nsya2
KBVHg5VW3mL/HQcwKoyEIGzD6i+yLcPB/uj+nZVgFyu+AJtU3Bpv6UQFJgGlPeeH
wOSBYp4LNdrawWcv8xH2DqKw9RJSSMnjpw3pv563SS7x03N4htJE320ll7KM65pm
umLVyzoeb7qEw7u7l1i6NO6+QnmQIFD8QDdX6l+M8P02K0c/Nyh4q2XNYGiENFEN
cZIkAce16qFzmBMhsj4jjV/ZVzvR7DlAmmIFeJx9E1MNd2B87WKGE4c2y6zJLIiV
+r4v0haTWAmgdvddW6QLXozxnjcjt2iyj35p5/w08xc02SYwhlKJh9b/kBaKIOI2
xO5SFvHb7ysWMoHicVL3HZEuBDLK4n88lQLSHP2lHDJEIxkK9btjQ+Y0B6Kk4E8g
Wr38GWGX2YiuJCXOZ78F4vxBscPhS+7MU3TljtgLq9Hio9fFtuaYjnFjzaHFRRqD
Ks3MTuqpxtSCZ913cN3lPQUO/4l2WKJsUgN7WBR1hEZdX41x3zlEmOUGPyFjFW4P
71aTiMwttRtAPcmUxi3hzBbnK3yYVUN0trhBL/I35ESDXMNma+5/894ijU02zHCr
njb3O05gI4lPIe6NHt2PLszng6HMa1E20p6Xd45CbeSVR8h3VChvIFJZuVnmRczc
qdo9NdsA4sp2F/ad6JZE305CsieTQF1KX1KU+b/PgAmb2eI4flPhM2sb9a/JAGLM
RgpyfJYjtoh7mO6sP0dABxIgtSbFseIWVCyV0xLlxY8Vim9bFQdfZ2u1gGybAXf7
jWJFnswyLeW+EnMtDgnd7JsgUqKlsSFW0YnyauqzFkWqrdV3k/38SMJGGiIETa0I
e1f8pUBzmsCLGhAgsoOUqLCrLU0TKyb36Whou/PLkroU3pdtRz22D6SvpOGf/Icu
oG1l1+P0PZf8zwAnFU2drhsXF9KpES3WY9c2XGtOFH5Bn6P34r10WVJ7X2HUNAyE
lnNVkHH/F6ioIcgFOfCCX9gPZXAgjAP7fl8OUEKKMoHfCM3GtEK0gtTs9rxUQVUg
sUIyHxLAsWEHcoQeFXMJPGpy2+Fz8lSkwIazmzW41+LBIxRSlYz92//l7bBjcnXD
IXHVxGehBsBrjHvBVn1HzBwMM1YlE27gq3tKy9GP+vJJBs51exc1EnLWLQyejP+Y
GEDZ1JjX1RU0dK1NaqhEi9SadpUkhrDweZTaaRXmnI28ufQrbLJp6Y4AWKBEgDvc
Iy1JCKlDLQ7b9hv42mYT6kj6JHPWrlhJ0QhYGtn+hbOgdM6G5nI8hG7XNYl7yDaD
mJp6h7T6cn2B0yj2twumnEbnpcVDTBdweA52ho+snEY6NcMbr+8/MWN/di38fnL4
UakN4Wwyxkg/kk3+yewWwVG1+KMZMMHQc0OaSKwM4nYXsPzii8wRf2rrXtUumcyv
sTXMeZGssN750xhCqrmlY4c0iDD2yBSrjQ/efI0HZy8dMu0aJZ/xtiIIkT/b/KKD
g+JOk5VfiaPuTf2ml5QBiYlvsyf2sxZjl2DnWXD0EykeZXNW9CHnXyXkFlPwO+8k
SFs5BXQxK02nMPBypX+UhVW/P2MNZzwo3RPF5uz+JSkDXtQdcaDWKU/zdZoMPyJS
sKQ2Yqbmwfmh6ZfH2832X8GU5H792Lv5gUcwIwZNU8kuDvLz8ceEsPU7x/S2DiVO
VRTwC+TXrVHX5gFFnGecPcYwH4KY8JBqMzQ7R72cakBpVYg0YneV2JLtUabMqFQ7
MjYcr+HZkB6JIVkZCP4O8uGN41u8Fk6ygf8mMa8btYgTH3hLY1WfEZPiDJpPJ62J
UcUPOBoxa5MDqU/IZTJBN7SrIlTZv9KFTYydok480hTFNzxFqSLc5dJ1tu+ce7AY
8x1+taBOuTxOYe0RzyKG4VsNzlMW0ZnGUoc2iTR+SOglEwgHZA/b/GJl8dDuvHlj
obiFNmjB6dnbWX/u3cSQ3DbIwEaMwvCYS9iNtvDaBgTp+1apXAbGpYaiEe4Pnpn1
EJCMTMHVgyw0m441kCNrWZPEBfpLdleMx4dqi7IHdhDaUaHAT8LbRbVa16j2kGh/
U29Ny9gNNxkN4dqLmK+e+nEya3tZo75DXNonFkhRf9AQB9QxpOuEGQoVTl9yUILH
7QdY9ffwBRU5qe0tR1Whl7Bk//APCrvI3wM0xVp30a1nPdpALZIG1CTZynKXISI7
Hw2Iu6G5fA8YKsw7VYguOhG0ruuwE+wrgaTgpeofNBoqLiOaw65qXVLyr9gAX6A1
G9kY+b2FNVZN8SjJCdhAb8volJrfEIyQ6PdY/9CzF8MVeRW9qfXRxwOAE8ZkP8sw
Gjj7auduRSAUNEBV79vIJPJO/6YKVC2JnyDfYrMIogdvqyUoZOriAScSXeWjMUSV
IYJKcwU6GxLOkC8+Xg1vwqHU4ho6F7RKww7gySFffh37L+CJbLFwDFj42/oTFf62
Hmj0tHjwcBw5WdHO2eV5auNjnLxeaLGVX/IxKywXAQYzo/b2uqZHvLYk/wTc0loN
jXnOaaomLDcJvnN96Jx+oywLkiVlMSD75HjtwbwqFfHslQ7vtxSM1gVQpt7KRnQC
ZOmAWRExSzCUWouPIDhEW2Rgaok/we9ZdDln8df2VseU5Aas0ssOhdpXWkfyIj/i
RL+Nt2LGpgb2tAyt9DlrRfV32/ARja4yVo9UqQpF/DUOpSrZfp8iS/OSbryxM+T9
9m2o5w7HXGeIiSuXHtHOSQjEzlsVJ1LVjZ4AnLOzjvUwRn1PGQmvN0KeC2QdP8Zv
/bXs46hxZsJVKrjMXX+Zr1Z1haU6cd+gzMOoVLaIZV6FK9cfc5dw03No3zqf16Xv
Tg2619iHfjRDjtjHUb1lYYAdg1+g0X1bvhcPijmnzXMoZxH+s/T6fAIcSS6e4Vk9
LK0+gl392y76G2KTRIJh8iaKlDh5+S4FHv2b9aST7tJlVlsqdStUUvDRzjb9w1GZ
E/cXfJiRQRIiF7X2mypmnmjbWnoB4jbw2LPN5qMp0StwymbEVGbMdbxKJDdfdr3g
yDaDQ0XRJmsBeYh43wbJzZP4+nLZj42JBjzw3wLfHDQLTdjk7sDiCsxekjw6zvCG
e6YnTyxhj9xQtjcS5nQqKcBqCwNHdE0QUosilzohhm90u/pNzhfzUdcK0OovfYpw
39lWeuqyKuIROb4pCKKNlaklQMvHE/wJ3+QQgaulkhzoMgbmFc/fciLt9/G12Ayx
wYJ2KLuOacEuVEBglsI+LRkumF3kuCORtZ/SbPdsHH+NEIsEYPiRhJRX7DgZWuxH
OaSl8v5gIAWGoTe/mgWA1z8xT1CmUXM9Y+EetgF6tgcL9h41tfx6PiOUYYxHevnT
Yam9roBSK3Y8hxYCfd3upKH5INhUpOoIeH9jcF0OKrdUKR2akq4flLg41CDYFZqU
IAXXEA+UhwTJ2kSn5DkZiqViF53esvL20fq3w7yZaf44yTDNNZwPzpLvVEb9oXsa
9TWyGt9FK7+X68402J1iW1D4G6uncdx0lP8W1MW/3FkqOUza6zxNwuHkVo2vZQvF
gS+kVOp5+OE5VziQSy5uSNjn1SbSiQbI6tmaIWuACdvHuGEYfrRKQtGfw/Qb5KSz
l9yxINj3ewmRsBfRDasjCuJzAvcuR+Ow+dvbK6YVGapDb9Gnu3K6j5+dtsU3Dgp9
fx1EQZ+DhzEQFTwmqXbl09SLb8rVtvAdVkZTIxQkjDTJx2uxj12/THfsY1R/2c6p
8JxWP9T6LP4v+icSnbVRiO396+8hTCZYA4hrFcE1W0ILptiGFOqrHUS2p05iitd3
4JwPohgWHqmFvIPIveilsdrZzlAe38Iz2uyJ5vErd//rWd8Oh5LeH71ifxYMvJJ/
GD+25cABc8Vuc7IoWNUbE+P74uHg4XTop/olNUkypV+ac5YIUBV1AOQdYTPd13Vb
FtZhIqOJJwqu8trp+SNM8yuyOxp9nxaZbdWaBZqtpHHjzpLDrsNwFohHeQAXkJkp
XGC7Cb2ppbcS55zT4ONeAuF2R5arNNutXy3r8wA4dVcfFX8y3fHir4377vWvbSyI
mNrcKOhTGLRdsMkJo70+UrkZipRoNa44ABKFFCwRoiakj9qlDEOW3edQ2pO05dVT
MMT3u+mlgSO46DxvLIo347T9meQ8He6su36CmW21aRhIkWn5Dq7hRJB4Imyd+l+R
FpWVL/URK48IncCg8yoZpnUol1tvxb2ZRZmdXAf8+HTZ0moK3LHLYjj6Y2/D+dFs
DwvMc6mhSU5s6VNKrgQnMKGFnpK8hvccf170zFqwDwJY5NjB6XwxfG40GH1Qbi6+
xJRm92wzviyggDRtpyAEi/7DjsYzeZvElE/TYI+r9Uzr/vl6yl0Q2M7YdDBjQcg7
YMdk4k6STCNb3xkgE1mV/GLQoSuK20jT4+yGi2BI2KOYelrCOJcY5eDQ+QvgS2qq
TE/nb3pW45a7NdRRdaxC9HZ3vz7mEv4CUOU/aJ0OvgrIAmXVgKq3S0BLiNY3r+YU
moIk9BET8N9ROtpvAYDyg3bvUtkurv7WIjawvTCI0082rOWb5/5NKwQGGFFbtw8P
Fdkj/r3h4p72vecTZTrTQOwzXeDfbseq4yjSQ0UsxPNZZLSUN2CXJGaudAbkj/rG
FxQItfgAkQ84D2U1gvqGN6P2XsLsnVGT7TsqYwAVXmZvHiQzV4EcgktltayJMXQ4
KRbXyv6QvPQ2p8qzs8KH1+BQOnkz804F2+wwAKvDNM4LBWvsmGD9dbfwVR1J2Hcj
9Ki9sdW4D1UvJsT1wIp2ngbtnNplBElkDiht/qOUSpRqyBehteM9pswzpyAyxLKY
dowdBJsEybdSGY159x3dSR0FtEI9oudFLQSOYY56ds8o9FBvuttR+WMOweTOzqUM
XONDVwE/+SIk7qCKFMKXU9oW+6gE4pJo1hUpc7/K41Lc/63qSTXLSi65yr3/Nsku
SZMfFBsWhmhbcpfcbfyozuSrW21WL2nKJvWqmlAeQfNz1TZxXrM21BYWfDZ3y3io
63Y+OyF1kYnP7sfKNHxNCCX2EeyUPmitt17RB+YTp3ohXiMDvDY2p3e7rb1J9VDp
VmfdaYZ35X4sfpX87cmcFxJ8e1pB9AFnJ9UkYdmzFDocmJg4WM029abbXpW+iwyZ
xjyNEY8tMf7pShouADA13ynQ5kgW+hO81IgCC5Kd4rCHq/4cRxIqCnJAfxuRM5gJ
5jhvcKzwKIa9UpQRnxNiYEhAvF0H4yJhSKJtV9MQY8rXotko6mq/wwQE2Ps86SWu
o7gCXT3XyIbiW7NOPJHKCW3j8JkVipOcgcy8ynv8QzcPqV+4idJihVGXnDT9U59e
WmPG7pxvNGxZ+AV3zoh9uNcD2FF4AHGXL761gBy53vZwuZjkrWwJLdsL6Ryc8fF6
eHghIZvLpNh8LMqXQDzs+j8YGpzMyq/4Yj8YXPJudII7BRjmj37QvbfBRQPDbKPL
GhcUCAN79wDcYu5ntaXzLaTTGHvCRwH0rNfnNtJiqacAT3BDG9krVXBmQhtqYDEM
dc74Ikn4yqL3ShpbhFWkM+BmEDpGCmsjh/eslBOqdWEnnE2uAexbBYviKEFRSjAH
jWVckNbHo+KAUrbr34U8JsDaKO6/yYd1bbHQ11wktBm9iKR+X7H7DTQqwa+kJ3BG
GB5gLXpj8UPhPmedd8t73Zmk6fY35v9iol5YXqdoiRfC7e4+q8MQee28WAEMnDVm
OwWLdtJRTF5OUp28IKhfI74zWCBrqZiV38CDIsNqDNqMaXqLvjbqP83YuO58oiFl
9cpACdbbYPkONvKZOHxCRPp8wQCeHBXePcxaA+3UUNIVFeduhDzGveOzyQX2J5Pc
r+0n4OrHyLprEBwuaRC6vhdNTzAW4+cKpdMcC70MfQPyxz26o3WphjuSajProOq2
jgRKjkQ5BUsifHD1j3iaOcyibYEAy9GQSnNAz5C3qwo49DOaj1olyesb48PxaAYI
T9OL0oAd2MmkqwJf+RCQiuAnVN76mHuk+8VKHSLWw2NBPuMFWvKtZSoHML2TWla3
eCfSMS2OrgSa+hrHtmgHuYFOdmwjhTpPtGnVKv0hvwCE5NwzQx7BdBPMMsyeQ0ui
DPUdt3FpbiLDfjg8PrBqB+MbLTnu+XFwhAy4qwgnKXbBsUU6IndiK2EVaEf8ej+9
H0VcXIYOuKDd9+phJrJt3nG/rghnDDN3SwTNDKMpaoseCNM+92T7uCzdW8Uv0zKf
LZu+o6mdd0igC3WKVriU/J0wllu4OtSaZZ1sviQ4EvNGGWQFWkuS958U4qWiTdsz
TpotB2B/3wkSlstOddPIfYIYIPaOeIZvvPEvreQGrVuULXEbZdp85DL8TpdBNsgX
Sl0op0Umq4fw15B+cuhWNnJ6YcFQkCCyaXQJq2YCrcjCTogXSKZQRhQtf01cRz1Z
gVEmTWWsgE1oRY/4GUxWBtIKL/DlcfdoUuWjQqAma4ChKGe/3HBc1cY9iz2aTjAu
kp1FGQyV0LSGUsB7cQllXnXyx7WXoMiiG4IThTwKTJqqqw1APoU3+FW0nR5V9XW8
V14hjIyqBvzTAexENRfrqC0Wmjs4IR520zmUjT8bt13OR1nGzlFyMuxiUIbUCVbD
ECldR5l3VP85z95CvrbHc465tAYwRB3TRvKf6dlvRKl4p8rlWgiOsQ97GzGoMx/M
p7kt3quNft22cT78gvE2oAAR02KmBx43d9LBoJbTdoOzriEl14ndMDcg1HOlZ9fQ
a04KFwqzlOfb7cYw3Z1Ev1BkiVLko+VtPBrAKsSCknJx63Cvfdc8vVX9O+PEWdZn
kBpyTNvbKEnKx6qd9ZeX54uBNAU4YzM9KnfIjIB75/rtRL6SuLJYWtjd82J+w26X
gADAMu2Sukyrj80BjvP962l2mk+YWGUCTabqL5twKllc72O2EkXP3Ig2AHLPOkj4
//7O65FDtLX4qRk2OCbpb1GPDYSMAz+C6iqpBHP99JxIqhme8PvOc3f38CGkBlb2
ahiusl0hOSf0VMzu94NNVozZy0y+16ARO+C0aFKHCqGjpVqNjEZBx36va8RJD96a
IgpFeLjPV7dirhrizpKAh3xaIXjIQ1/ZkPPXQqPMS6Jcf5g5CLBr3s5zYKwyUFvw
YDllUbIIFb1Jemi7qk0jY5zTmFI9NKVwjMroy8+FkakBWSXzU7csFx80LNKvTodj
9mRnyNEGBuDVamSJ0JBDvxyvqPkMF7SLFeBT606YpXDXqjPwisxDHcENp63XW7cz
N0scSWJhE2vqbKXYcckgJN+kfBX//3RZQ+hBu9Oji3Fz4kERFM7ryi7cBwzQyKHK
XUVy1kLOoBpV0nhZSTFxJFpsV987rH21jyYJELE8hyp92aSi0x0JLT2CNHpxoZFC
rL2pO5QDmF16uWF7NXwPZIHs5uZiMJjhRTH/dv23o5WxzpX5Qi8LDq45c0Mooq2a
thb89izpQ5R93g+0NFBeDO4F2fUled7Mc2LPrGrqIvdeXOHnoT/cpXqnOnBvIDVB
qWd+Wjowh8XajTecPtfo94w+D/x32cbzKKUu8bANf2pqpDg1GA5crwxovSy4B+5S
i42tVOkNngqxhEGGIYmXH4l9e+CrfU6D3AIgRkLE1TmotknrKn66y1S6O018O6XA
/8TXTDxWmhmDci/wqmILjLIY02/+YZOGauNYtJp2HL/fPcrT7aTlG51SaK6NXe7u
0paabcaYl3mRoU2u2VoRCOqg5JGzImMZ4m/gtjXa+5ip9UQPjsphwkGTqWorOVLk
APbYoovZmapBQG3+VyPkuilwE9mDdWTXm7czDW2EVLaOtXMNs64MvoPy/Owt0n+5
DNbvjH35e7xqCrxI5+NKVdBtnD51NuQAi5L8KyLpggxQ+ZKdnJRM2Mk7mwt5cl3I
ABe69VnzPkR2/H151li9y3159FfN4wbt8p6afQbdm4HwgmDpwQJFAJWY7D6n71yo
jzH74rDesxMXI2iv33EfXP6WfJv/OV3M+MfQqlY5xih1OH5WjzqVDN28MEbBJer5
wA1UKGII+RIBvsAx1nPSD0P9ZdVFqEiJXBeme1KYqQRdwK7B5dPnC5y4M0mYo51G
xaZCDGQi6BIOvOYov+MGvslj1tfZw5bHjgI9Wc9zf9kZzs7Olt2lqGVyRjccZ0AO
OXGP2JcqqLtutP6HOJ5jWStcj4Hdo+W1SuGygFhW2QzTy66XcNQIM/BAGM3bacOu
0Idxe0AS/p7GNUt59BUPXq9khsmcfsR0JXySy8ebdJ41pfOZFw0l8kEhikuAJtq4
3AimSzjXm9VG7IZr8iJ3M5NoiCBixkchwKV6zjpw2uyAHZ2wKOiS8zoZXBMXkFZ2
UK//8DF5HS5CW+X4zrs3pdXFUBGMM+l9NDSEQH6xFfNgsM6cxXifiPBe+5xlXSBC
TZLf4rBknjhiScREtRXoTHcTuoMM7WpaOetXawJ2VsemAD54MDx6K1x2C6VNKM0q
o3bptjHLPzW7laiifc/IbotcC5amzlqoRGudLrI4z+YZhC+6HVXSGRf027xYpUZG
4I1q4uyj9s8J7US7G/qGR5ifsOQ6WoYAexSaQaqERE5L97aoloiDXrXyJv1O2jz3
SpM/OcQ93xS9smk1vRYK5bxrD+Omn70HMH2ceyX3yx8pk5IFDPTPuTOVYMuXMfv8
czGs5szWYmofTb35g+oBRX+UPos6DvoDVL8wyKejxVe4K6RHGW5WDTHOYNfRuz0j
PkCJ3Oiw6/rWDnvESzQS5pQ+3euUt1EElgWgR5etXOibeg1HismE63grUC/2ofCg
Q3a2W5Sk6j0cNW8WPYhN3cJPfLuA9xKEOiEQ91NUJVhncyNme1xKaUnN/iRbkkNE
nJkU+7bHZPMwLaVrAYe7gqsepMw2j3/1CMj19u7yISO8uzmiQZRb7tCtcfeljkxD
iPb0B5ABuUJHgIY8ONt3qyyZWWkwA00dl0i/ufRrtvBRqud/w44tu4+eyd3voRuu
vmHpnf0vC1i1QzfOBHu/OWu+EBke8nD9kXaIaXy62RjSX0zoh/aNWJ+R/DwHivkN
IFjXIwZOCbAv6bmMAPYWa+KUJxNRJDzn+7cN3K23xYl3Crn6FeXHtANeUr3PFXg4
oIcLmgfS4eQb+5ErBSmyKmdGkFS21PZTxlZDSCmX/ge4OzeTfhu+Go395FXS1ZML
38+JRcvZZC/xEnFmkARzZ93+semBI59lt5sHPuLz5BMefAcOjGNFpmewy1RuqT8+
zjtD08y0t6bthv88SDRrmuWsaY1KSuMSTkLi5thkL2Ca8qph/paXwUJs9NVUOxTw
nwU7eWRZKo/3xV7tv41DkVpXKNKnmj0i2Mkuc09ebAq7nqQin4hrUE0o2XOZH0+Z
EevhKCVG1LTFum7oqQXdQqPYb20+4NBrgU91uCXLlO/EeHRUNiJWsag7cT5WEftD
P5cZo9m5Wiw6/3Qs7mwl8gZAFuSFeOST7LGPJ4ztY8MKmVvmc0FkiyMquaxTkN/l
Acd/BT94YhUXn1S9UN1OyMZWte6chJP/fF/A6IAVKQHRoql5Pe1KOCawRN5hU2b/
jEBlsiRrMEE0KBRSHyj9uq7gHYoq3SWXM7cXsVi5r16tHkk30lp+5GkzAoSMQNxv
yPCld6FLdmNoiMmI1tD49crKMJ3gewj6929bl1Vx2c46iUOaa8czPmzSoQGhoJwV
/ZgZzFIHYdKa8NqVXgq5oGDGbx7qulqsimYp6dM2QK9KbOfN/IZO8x09/Qpe7V3W
KiBHcvdvU/d2d8pldaKFwYCZORmPhBAq+K7weQLj6vHgQcOQqRj5u2ZK8kGeYn/a
4QBfszpTbEbJtqZUOF4ay+aWE2z49dDrZG360kqS2h4WPwNtGgQYQR8DC4kdGMbk
QlRLmM60fD5+BgWV9yuZqeXKz/9PxrX+Efhoh49u+e1X8F5itpkbQwbXCnA/H1Fy
LOxp84UqQu+ICPdU653Qi9hz6buB3eX6tPlSS5V/6mIzB2w4j+rDp/681QlDS5aQ
MgHsunqCfGnPCyLbkycEU7OGZOQrgujIA2fz8+3VPQqA1GpzikjgNpv/u12AWx6N
6b2srgIzENmAK0lYolx1rIO/Wa1IF+5y1pSxJkN1SRMj+Xw/O62FdMtMuyifh6MS
JkBwXgjcLnrO+Iv/GLiXCmZ6OKK9Jay88ihf2R+T5dgaSK1XwkWIWYlVZFTI0crD
YWk+TACwWb4KshHGv+yw0b0y9GHqqgydyXEqiPvmsv2s/Wx9ij/SvrPfmK2ZVu5y
+5F5p3VqUb36pFI1LYsTPEugrhbo5XlQupkOrfcWujDE/wg+jUDXYSkt/K9dAJs1
07vPqcaBBPYPxuylbD0EIWpt6VSPW76wHAk/46PC93KfG8zQv9zAEkFfBJOB6RvF
sts7WCBCktgfKj8SNzzYbSpNQuiplVORAJ6+h2u9kPCo+rKeEcImcz0I01zpm9TD
161QeL7BdqGAhKbM5PetuHZN0Mw7bzZ2wOTjp8whhaPey/DbHAqa1ErS0t+gyyY8
SQLHR2GWfvkRPKmI5pszu92M7JfXos9iW1hTBslQyY67o/OKABFVlfooN4feL8EB
K2ROIkJzt1doxaZpwNXPM++v8mz1VXT0RbX4JuG/4L0iqIpjN3guaT9rllh+8gJZ
f75O+NsnciFiMtSPT1FhvRHbdR424PNkj5e/L1RH4hVzxAOOJEPJuvYahdyQGXGW
0vSyb9/YIQWuQlX0TqPDf08vWr9Cf/6We1C+1d1K2sW6FrRuG2jyV/Oxsn13T8OM
74qVY/GyvKSUKy2/oeHIie610+IahkPzrONp2TzOKhHEnlH7zqfBNEIFRoydROUF
sF5z7lI7TZr0No4WnumkMJnzcRITmnznrjSNrA98Nw3gOGIO/AcmYMHulqrLenli
4wYF3ODLhX/oDSzHXWG94/VfLAxASHNxoKbU2OW/r6c/xqO5F7E6TmaCnXKRJ3dE
jISVg5U6hKEo7WJtan3FWI9/LRvskiqaoKF5TbAzrus/k9mzPskOLsbUeyoxVNDG
mySE9IrmtYiB4K/1auGfWsGUAuR9T2msN+1bi92lCgX5ubZETM8ERsxbAhqDFVeE
1DT2CQHWYGQB+GQbxpYnJcmG/drWzQD1SRZcj5+N3mHWDIPS39GHxAAxKCoONNvl
TeRjCEIj47g64lMU0g9FfagV9PFx3LBRzNHhckmRj4echt5l/wEhc70s+iSIs1vy
/FjDi5Mlhj7XvClDaarhBgifsFumGFR+f/Xhs4bgPCg7o4f1T8s1ElJX8+/H15+B
UzbCgNilsx0Y6sDT3RYZrI9G1idZ091sDfZfpaJIPAKWwN127GrqbCcmfD0Zl2Hu
Y7qz6VNnVD2NqquqcUVY5PSOyiOT2BT0704L51CRnctX2vKLBZNFp6HmAcXLVYJq
MSqxjnE/83+gn5LCLD8VMI8sEVehPRkgoW/CZSgJi8aD8EnTjuNdfgtEoAujk683
2HhqXeYZdKzlQwGe7Aj3SRXJcL7fmKVBm/l6NNM1gdZSLrSTi94VL80SjyktonfJ
6MU0Z7Mp8cPUqFnNOu4YTFk/Kgjvlslp9WRY3FGJtBcT6P1bMpgc1KQ5hgvMiHQd
kulZaeYroycNt9Ke9Ty5fbdP7xLTxU7qjQvgjoKni1olHq6r4FNpdXaTaTXQpF88
c6e+nTNg/TlxN2grkQsWcxeq6bHhgfwM6Eh9yEAiJUZVsfAVArDo9jeTtLDpvVfJ
sidWHA8mMe2iiS9a7H2nm9K3fP15tAuruKbFocVs10mdfRppSXuqRdIx5F3Yjyz9
yCtHl6EAcn+Wf3Gi9yxHqjvstxpajLpFCRHngZqHG1EUcKcxmrNUF7S+7MGePjeG
LZZeeMFjdgmtxqhmTlA41QXuLJObrGimEoAaBNPCpDEBNPP1X23UawPsFm+GK2UY
/iG0fXiHi/Q+1QnbOT0CXEln8QmC+l5VWdWN8venJcx/PU7RAunKBoBvuCD7mg6K
1V9dMnvhDlWYn+EOKRXbgcMO3LfcNWbZFeUqDYt6NjpGgr+qdm4J8CjhY6/HJBAC
APAAcIVPLx1oe+I9R5xOcAXJbc3h85hFeOdo7/V+PCEU6LMIv4A+TF+yuGYdb6ic
n4ASqICU2I34uL5G32sHa+gfDkJp2Je/57oddbPwn0ivsn9p/6uEIBuzl9Sp5Ips
q6XjOCsCath68DKNYaFvdRtEyvZ+md6c3kpxWF135jBg4lxMU6ZHqeRNu6E/xjw8
RyjC5C1fLrYrLFoMCq1vr64DbFvOAhllX/tBDPLvraarMgd1EF819ssMnCdss5zM
ju+hrj1Tnrn6HsFEVdhqVnhcHnnEiKKyLBPCtXyKLofD0G4GVM6hGMvzakUEG4u+
AOVzxoLq/9fiIU/Ji00RkaVN+/mezctKF6w6//zhERRNiqFnatiZoefClQf0hPBh
6JjEl5jShbG04CnC78bSTT/aaejPQ9BGGki6pYQinTMEA+IXls/TgffnfcMsv+kK
I1LE7bIQ4QbCnQUgCsWckjsyio9/S6y1OgnTwgaC+O5ZCAp0rfLJN6+RYIBEv36N
7FDRVtuLZqzEjpgtUXjCrZB4SRqHQ6uqzRr1rCIjSXFVHxXOIV0/mOn0+xi2sR2/
clRQ2H5XPX3u/tOOzGA7QOEN0ZtsjYT7zXxVvybSA08uFcsSbBkvp4vYWjaOVLk3
ZBzInq5R857joODf+yo+PYG6Ra1/8XcM53AkxhtieLv76S8Q35gKZ7XhbR55eeZe
kbZSLu47kR0t3Ls8NmMi5jCCG0mEx7WdnFChRKEj5re7vj70AlD/d57TpuenOPu7
tQFsueattGPvRLll4gafztcjjNr18Em3FQB0PQvYrn0/xN1HP8f36G+L6/zrURSh
YFv5SiJ76ZLD1PV6o1JtwgF1uZpiQP96P8/0yWsMO+vXXjUojTJiI21xXriFP2oP
qWWa8KdBrsCNOXzpbpMeFMRTUu4rBiur2sfrGX4vheyqjlQEGI1mF07N2bCrAG1c
KFxkANmeB2UVJ3pRK3TZsw4MmvuFSTpuwosmxS3Pq+a8j/rwzNH8xkodMTyMXAc9
tJ3ePSYjLJeu3nkqqv/OptjHXxKvQo7ahYcTX5jBx2R4sGux5abt7ItM4AUaPBx7
r+/b1hl9vpfCb73Dl+rLJa/zjxGfI1cJMGL/6FF/BhFQIaOKrtUryW/aNrZja3bz
F8siloX7NUKvliuWwiMvsVijITgd4TK2uLhmupMtnGE8Jrk5YGO+aNJ+Bwqry96V
LXQyJK1iIIJeqohE39VcqGY0aFdUQO7lTSWc73XOnbiNU71jQ035nQlU+l/53n6x
KBKc6N6I4lLjoTOQ6YfFSkKCcQ7TAtKZbbIoDqFKyGfx97WWVv1cE+BH3JIMHiZj
33XTy9q9s+u1sv1yJVTKgsk7an7FnwuWNItWwc1pZYevcZgUlsHIzNBsdgbiJP59
rGrRWq9AabJr+7CNqz8lYEOEPFbXNSP8YrkuANxdHdWDJ+ncdhAg81sVzd6EjI26
qb8B7cn5Dz9Wx1a6tTpfNYh9OhlQigAuPyxC+WSvJbP0pmib2COkxyIlIBBDYxJk
pis4Va5UJqegWOc6MC8FZ0riIDR3kZyJDwxoNuzSgvFhcVptJ+FVMyavnhTCfJ/0
kQH6T+A7DcaKDLgokXshRT1nyQ5XGTEumH2CxGXnDWG5BqkVB60r/c9Uxts1tCvp
UYqPitkkyB/LDLCIA89ujJZ9dfhVPyw3zTeS4OUHesU+Meujs99iftRKdGlveIIB
kVQKQXidxoiJW9DSI6n0+gPN6JZ8Vks0/y41GbZmWdsfyxRM8JpDPQY9LohdzOMt
Nen8X4iSAJtGzqeKoY+U5UseSSw7e4uEyMy4DWMl2g6TbfKjBYBwtt8Sk1SbqigB
iwbq0geAwJtyfSftnZ3LOiQfF/FHscrjCs+mv0qdY69pE/wdbN1D6moRIGS4UxNd
upa3ZW11Ecl+ysWsFH9LBDvw+3/63dQV2U5fO0NsVmVzYJoRGK4mWgOk5VhljfY3
DP7CJVnncEQ0Gm4t+kbvci4hQleuTKVadxb9BLPms+riWGwWa7lhl4PGHLim6Qmy
Ob9at29NJWMMYl5QV6qnK4fwX+rBENNqZo7bywMxj9vyF3ExgJvT42nRZ3citgoy
FVdF1NB4FbWrijjSWlzoGkdNmTGGToXsSrC8v5IFN/sv1qO7mtDJqWE9/v+/9RX/
LbvUACrG8WzHjOt12o8ffR8SD6wNQhhNvfS+7qqIIDbosE5dWRRqZoWjo8bNSzcE
pFetxfL4WkJnTVbMSnRtD2jo3sykzSa56t2eG3njOZGQDipsjrDrTwoxrMdraOKf
9EFBAk7oDIXtHogPfO6FOLZFyKQ477LTU4OaXw3IT2n9GKODJyWwhE1xASK1VnMc
h/fAqgXMe5aUkgCd5aHGNoiJNXm9BUeffEBZmlAy19pfqc5P8fN4ulaiREDbXMoj
CVqGhuznU4aVkcUpvIjjFEesHPyi7RG2R9EpsEMWvNtL1tDKMSITW5u4iL8ssp7q
UeahnQv63oUFsOd8m84bMfxo9pIZ3cHoDgwWAjWoT3jaZgi9NgXGCkcmV2EKITdW
Of7b80G80GBuMRiIEji23CZ1tl9v/UCEBixfj5Anj995VSR/JcpreRmd8KaRWoKt
g/TSwvpqoScATteUI+J2zQX75heRJrzGSOj7h+U3/8Z7ldFz2eHRuax13GXv0gr/
LkMBE3QnHEL9YGIPwl+vLYb3zJsNg/xu7kFyFJC/7tA3VgGs5Ed5MLBVxikw1TBD
q6INLe+Oz/HBdlB6qLw86jq0VkFhww5LPk0uz3GSaPwvL5gisX+v29txbskVX9T/
DLhGrS4XTf/46zM7T6ajHSWoqW/47JyEH8Z+PoAEg/6pq9YN6hx6l+u+MDh6shSI
M52aspdlaRNq6h28xNlRk5MeVAfdxl4Yp0GSAOQSYH+5q8bd3OcfnCChg5pn1RpV
IKNk+bGLQyBTjwE6XD989xFhU3ljTuIgDSP2IN+kRxMDW10AgM2WZHhH7GIgOzlp
SjtSCgcJrnSMjrlBuFvyKFN1F6XRCl0X6sYA/4cMCYdr0mmc8MF0zDxwH1f+BF2K
ddc9mr2yhE2kXywbjTd499ShPPr2E8S7pTVo8mQnhhItcXWuBel5Qfkzwlbpn0/Z
AvrIeLfcwf+Zm6cYc6zAEd2N9t7mvlFD/EWrhsXK+UK7t3uv1hMzsQwsJ/XawXSh
UZ29GMWIlgDYzfY/epTrQebVakuu87Kdl9YaHY/8TVfBtVICKfNwEe2xzhBOR/AJ
hJNAvjSUUYpLDLkixJs5XOrzBBZX+TAnDzPz58TgHM+tI20/zqWa5axj+hlR2Isi
vBc3EgSrgk1/X4k+b5U9O2EVVOtX1So87Kr3D7cYFuEPOZe8/jVRenS5vm/7f/Gw
tlgVh7Hocbi97SvnJn3N4iGKHp+wgmsA2bQgcPX1ageDkehfKBy4z4ZU9gbUL2jq
mlMdI+/c+QEcrLGnrtpwXEmQEhVhcVdnLXSMQIzjn20feLY3T/ETpVR0b19aL14n
w7MsYhTAsr+YaJ9YStFw8e+L3mN55dhVfON69vd7yvkOWsWAA6hZn1bOHBLl6+5J
mwKVZzld4Wu99NMoZbibfpQOlBp5sPanWDyALt3rInt9R4Cjmmk9l9AAtvMSmIvj
l3EC3OvM0KYpKD7SZkMvi9jExNB230xaohQRkkv9zEuMJ4Ffp24phfYvCB8jgaTR
mMHDYKI+y0Od5N0B0Zb1DvEShrmir1q1m5mBsC7d90IUKFAe4fOToQkZJFcylukz
BEpmHZqN8q9ouKG/V7hOZ4wVoZdGiK03jvZ03XUT8SCdroAeJqyrI+CRhW/J6jSx
jIncsZgxrnohLW3YOGexMevQ64RIvKwXynJVN0V0pIeK/I8VA7YrJ/6C4eErQxgw
YGQxA3NF8h9dOsLVIOxTaIDKbCmAEUuAJZ/r7ma8+lOFi4PRDzEBTtJ00hW8xEet
JmuiOa6VTGAecEjL01gCvLW7ynrrl8PqJRKwoCJtvpkmPD2HzGmJggNBpxZqfxxx
ftElq71TgSc7e8U0yHKUsWPY2fiN7gDPT5ce/NWVPuLScB5Yfv5nF/4hXOHhtQJK
a/WQpudBTzT8ePxVV3QIJP2r9jN9u8alKVSJ2u30r1dv/e80s8eT5R0T9loIU25d
iqF7x2MhggRyzc5u3D6o5DVatY//XCcmgJezCpHhqEuKudcxFuxvQXGMqXyR655W
zRpbrHss82FZ9KBq1UlcuTSL4HDJU/Z7k6F15x3dPGlDWQjTAIZKI7E78BLDb4Lb
uWUB3ZEz1dS8lju1gvtMb3N828Xa2YegEQboCKpWxeCiZjTTpTB40idTrJkQ6j0e
9XFLyog+LGmp+eaf1n+OgNyUrvoDOgfbdsqaJWG+bCri2Oa7hhSHi7kxp1U1O87m
TzKGOnnJ0Dp1tQhlJiqhmJ78Loy+Hi7IHTSYacfMZCOky6+wBgVQIloLA8XgoBw7
5VeiPIBlDlh8Vzu1vkB7W++LnT5P656UTLkhn4N9uOzOy5tsjLN81bpd415tniUh
JfFJNCl8hELRJBMQOXYmvBnZIts4zCKc0Lb5gbPNEssXiYYf6sa5lc2HbohbbIKZ
EIg1h8BxSNmjLA6Ng7kCDJY1oTKqEzZFsd52OzbKlg04nA0mdxcjnkUY3pXhmiQz
/7cZFA28sJs/R/ZsbLTqvYf4S6OpABxzIHX1P6WS7B7fR0QCgJ6AAKRQsRBJGlBT
5S2luzkHAm4EVDJz5WyXZMUNMMBjQKAySObH97HCYYyoZdlMTALypI7WsvkDcrAO
nFtLLfk/3UJv8Uiatua7g9BqIQp+G4IvVFbexl5bGDU8iYo2qWPKkbIOL9O5oPDt
hTkVcQVzYEejUbxGCxxbBPny37GFsRpfFzcwjDaRa3t2m0dlJNNPq/eyvqzcHkLo
bh46B5ld46ykUq5cdjxbvN+xqrna+viZzmecTudkX8tI3n4zY5bHm5IHd9IsFByC
6/DfICN9ppA508AzQcNCmMjpRoYTyywL2WEY1tqKA8UMbUE+Px/Sm9AKEb6An0lv
LH09JYmpRJiR/eHyrKD+iI4qtyWoum4Q/gjTg636ibC+aqfTyn+MIgYUoDYjwmj9
QktO9FRHroc+IlBUucBvKyxGgHt0EaERKECUVwMMprzZNLQCBtV78pO2V8WeEJlb
WRKEvdbbvQD+gyjH9GaHoyBp70SBTIEMkvFahmhPXE/FhmCqYGROrjwBdQO9mm30
fsB0FdrvZYGPdCx10xTlvg/E95gJXP4sars+X0FV9qKAoNbu2gESr2FnWa0volEL
67yQGlzEReFHfxFGsfPgTfR/1pWYF6qSymUvnQzKyHelAd4q/GjTF3AcaqoCBIrg
u6roOOAFg+lvkEAYuWmN6fWpuJXtdKTCWYlcGQz1qc1l04O2aBmD6P1NPcbro3TA
9f34D2Sn66SIiKLrrmMiSiwGR9fBsC/8c4syqofbpqOxV+bsbnvh7MnRGa+OQxLs
z4Hjow0N3TNpnQV6xpW9N6kKgd5U+zOzSmikLO2Oz4uCpP8+VodnQMnyPOuP5bQ1
G1Prlly93uwaeGZ+RhuPxBN6RvWmwR57cvC2X/3wg8cT1K3LC6MeQw1jjZQAP8Qe
p2CGh9jCWEn3Bkm8QM0EQi+3uzgTfuVTUnydaDSqFrtKERiPojkUw9rv938VXuTY
mrsbsbk8X0Yl7dea8evbri7VKZMX6uF5H7DLn2Keqbk+O2xGAcg9aWVQk5fn3ERX
IKV5FCptljhqMruVj3ibifB95e9sG7jFTRlAvIN2F8vfDM2IkN3m6Ykz380gteHz
lmGyzBCMEHz8S/B6JmqOsfBnIHJJmgGVFxb/T3+InNsTuSgkwmPd7CBPJHhEhM8m
+7Q3ZiInJYpnehY4vm7dHFcrlcSAnXmcbs797nfVQzidamprwTWgneUPDNrMoWFb
je8okYX5XgpH4a0+0Oc0dkyUoyW7JGrHL0FkswQXBDKwkwnvOuciJSNjOCNkX7jv
SQ2C+iTZdGR3M5tFwFyCqJkRnHn/Q3pdNDg1GgCB4WZIYMNEYyv28bLn08uRUgVw
MQJ4a82wIhg0JJTRtqWSz1+ax30brZXw6JWmotMWtw7w9bi6o/5mcuxDXgBwUuWC
mjhc3ujFZ6dNZh842nbnaMPiHHpD9bnr4uS8o4IkEI+f6RjhcRsspj3CvTGI8so5
B18e3IzzvzI877UDlzDovZH63ddPJQy0goVNQaIjo698Hln4uBykaLm8hrs6+yGy
ecFbKcm+XD1Vd9I6QOtzmbHxHx/Odb8QL9v815mYRxrPV0K5ZbDSHKfj1+DBuSZ6
KvwDmbppSE6Qr6CmMyG4cQKRDuSbuC4lMqMK5u9I5THbmoCbfqqvzWqVdi5lbp8g
k8y/2yHKEu95zUJW/ULcJTmxg5s6xxN0JKJqQMsv4oRBx05aM9qFj3PCf1j5zA4Y
C9dWzApffBhDvt4Puy1ZiKoYHDL7fJVAQooNt6NQpi7agSagv4BZvEIGy3bY99w7
6GGjpAnpxQ3h7yCQM62FxEhCgOKXKqMcP7t1cG2JDMxJ3YgBouz1FzIXWk/AHodJ
02RlPGrJtcOhh93VPdEwmKV+qzxakAnmQ84c3RB+3vlZxkECoOLX7xG6HPjmjq3H
pRUWUvYr2vBRA4FD4HbGmVb5/r0luAJtELdzBw3nv0gRT53GYtmUDRBets51eT91
AgCh6HUs9/GWokHIut8yMeNX3UlZNc+z6Tk39gJyhJ3HzD7nmez137NwToRmITfY
xARtsBOZVGZNIaaKRWie2KC+zHyOE677piq7t0ICAv4W7GU3TFny0fw9flurT7y0
o//pGU8Ndcn8OTRTRtSclTEYqvhLtKRQhT7+MBsY8YKbr8l1vNuXkW067BHkTeUV
w6SezuoeKIgI39ZtmH7UrM0ogmSuTqb/Tf0fD9YfTLZk2hGtj9SKMngJZBfpzH7e
dOOC4EiWhwwJG0zlkPkhvC/C8UGO7qeG3FkPGUhyFLf8YscqNjuFKe9Af9BsaFyH
8vabkCo1NDjaIpxR2IpNWOMdcrnmQjZYcUiu1K99/5zK67cuSL14q9FMQHKr98JG
cAY9JICJ0nknyG5nDmvE/ShtjsZMdV2XGfsqKfARMCQdL4BOfVe7Bdf+JzFf/K9A
HCkhx04g0FusgqkoLZCOzpfOopuejYggGSssR2Gmy9FDZBR7tbAza+CnklsQ3X5G
iwqKxpkjv07R/mauRGB6pDDIMkWOh1Pv8dUDqCJou39XCNhaCbv//mnSVL20bxmg
kVNWxEyLfqdVO/1UYnQNqhQqrK17Ejl0TLncXcd4YnlI7ZUxfOSsiX/fMswgRRGk
akRArN7lu//xu//WHlJTiS4L0z3Zz3dfa/iSGl8br04wJ8V0nNuWB5TBNBPZrU8y
nqmslwFhq6HJWs3eE1/VhZOaX2yjDdoSiZxGof1cW5vOts/DuZao1vqHCxbb5B3P
ltsmWampxZsT7MHkdlN+pyRfBFkLfMeuhnnzDWfcDoxZiObIH8B9nEnYL1zLdxXF
8smqWW3LGUwe9NrYCGDsIr1y5ppqPvNYZZDuYb4VECAXf7bn3hFqZG8avRB1HlMF
1RUMjOY3SBcZ1of+UWAtq3zyGsDhjosZgIcHMBvaTczxSIi8t+ml0pHHmi/6hTTC
p/twPypm33jIWwa0zfqdnJQdacJ1yPJRZIBmsqOG+aVp4eGPYZzAgJxXYe+Pjpnu
/0LMfun04D4n55iMxvvn42MoTcNZFTM9bNQzRCS70AfKCGXjV06/gn871eCKqA3S
g8RY/izobDQC8CRxSiZqEkWzBzg50DuDe2tbBNvmy2C4fZMVSFarQN0yKy24ShpK
X6P/39vKHTZWC8zkt+rQ/y3y7GPFSuc6KglUgIqFYPTr6aUBpPyqU7SncFexOsvr
g3zWy2QVlwOwfpVBMKopWZ8t7RK+afLOBwft7WKsR7EptCEyqlMTQsoJfYM3UFb+
/d0e+8Pa48O3e9NPfcrAtNepUEo48s70t75xrVEAAc8pLCOqJR5itW1cWeihMyBu
rMt9qfbI61n5GNfjU9KI6hnTPIzKQ+UQTrxcvk+8Ow5/NkgIRGUHT5v4xePW5bMG
MFRg7Xeb+BoNmd2G8vrudNdZEeZJxGizIXqKqblH34GFjzQXOwFJkauMCbAmkSzg
UMvUtVccgicgoGBVxCzdsLKU/BvvmGx79YqRyCSWyEWQckABFPp0VugDi1xLBUsy
J/ey43Ma0WFJ5D9tkmj+1Qok22cI8TfYfZoBndNOjMPPP59KcQTj/h57qT08bJE0
nDyDdfNu4RXRJ3F2HjNRUiRghi71LmunWzR7LFFPS54VvjEuDuV9U5Xe8oadbN/h
5rtirnf6E2QXx8HH3X6gUkLjv3UJChcMMB226xGgD5corWDiw3iGfnLoYBlNMdzo
VrOxFWfChpjQkNpsonn6PzOieDmi05FQjHySlDj0CVx6Mtq21m2ga38LWPlVi6IS
SOgq0utAZ3S7Dy3Tr+Vsdrv0/XqStO9baRwbT+15rlCmYA79/PHDcWfpB8dC/Xt0
mHQEqoJDpsB1N6okNncPa73IK1hzp81xWx3T7oQ0C7F0y1j0BGNrQlbimdvGnsR5
ZBqV7pin4+CFBmnx2b9hnkr31TaQ5vKtGvrrSiw7ttT5JPsJx4TAxyzGjNe/KToD
dV16+razRIuQf9YHcT2568P2PJK65P/zunT/BJFjwW672xq/rk73Mfof1Pqwmu3L
PPr3Oa8Sxbn3Fq8ewh0Dy56K3ifNsSMu+xqwFZR9qV1VmJ6RAYqUJKvQcOaRq2wv
IPNyU+jzGrPZDftt6EQPwUysf30+m8Fd4wRCJ/39pXFktgZkg85CUw6EZ+XPwcly
KzB4qV4Ee+YiJg/EkeU+U3JR3c7KSjPhGcbcH35r8ZCf4BCHxGFU9lzpRb+IC+0N
5ewg2/lFrwqoobkJr2nBJ/voGbWX/qHQzDexsOmDjvbBoHDaGg8r+FocGcaGpkcj
z5Q9ul19o3vBasFrI14teVmKBhJ0glZicc94N3EV9F59apuD/bk58jMGBMibkp0s
ugQZXli58Pl1o+IneKXSx3aKBoBpB4aYfMmxNR6sY7bxpsTo18gmMAbLDq5nZSyv
VOCZGSpeUjrQxaT+8umk3UQkq0FRZygyNKnfwgVmDLTsi1N3hCsavZq5j+Sefub1
71Z3xY4LU9BrxDOhEnpb9ynwBDQUK21cOKAchdgN6hVhW6yIvJKVAmWDNP/e92/Z
pXLTHMe0PMG4XHuuDzNZ0+yAK0nHmEGBgnzR4w2Kt4wIKiOEzfb76G6PyATfq9TJ
0lYlApA7A4vHaM3up/5nVwrYfpsFax+S9XqGDVAnFa6bKuzdYy4DVHAAhJrdVYVC
M9J5LWdTowtrEl1bVhE+9zE96Uv7Yh1KI9XNwMG5qV9gB5VK/U2PtSNUvPQbUaC7
zfk963L7WVGc4IrY8GVRjffpAQN2Wv6yLsSPKme8+CUFJZFLh4Wtgokjh1iHgS+l
MrnblJy1AV57Esbxe5wAqUX4tzpB5dpkG9uwetgpLkf2a2Ef8ISZpJQzKnwkiTV4
j5oH2UOSufwZ92BnAUeI3dfg4aHRv0d9PLCDjkI1cT7mnZ3tHrnr3N2xR+YNucfU
raWCIEH1q73QYT1559jegfgv6UD79sDSRZ935yixZaYMXDiGDwDYwZ7B32Om2fJa
N8662UUB7sPY3Qo5B3ZjF+KIlLiZXmiWvtXLcLyjZul7SpiQN/B/qfu5Pr0MpqQi
6mJeQz40ty4fMVpeqSU+DkoJZjAWl9QhSwkEDW09AtTbVAm+cus+V6le69rFQA5X
1/DpJcPxKxHeVtPELkFul/VaAPAyo4I//kZe/gZ6vdSE7avq8VACiec3DS/Yg2/v
oXaK22c1N48HdKJILtSfbGTsj6bhoUjNw7awa7+A6kFKxnsNEN7PFZEwrEE0FLlp
dWnzjNbv5C4UVXOG6tAkmofNfMvm8b7T6LrirRZZGSOw22MhbyJivybQZvWITxOR
w1UzYbPpTkgQ/CVweKTUVJHyAdEj3lGhVgkxfj3jrtnQDLuKVz9t7jFFxCyymRC6
3qOMASpvS+xhHW8ByURAfnK63YBoUsH4RgcJR1Fcd6/8NIashgj7fWOGIzRb4snl
MDu210u8ma6i7PFDRgmtJx8d8anbossqk1ieKAxXN2dgHCXacNta8B+kNP9PvClA
D4oR/QdGDLIKGhZ95zJEi3SYUgxMNnfkMoQCSje0ghWsQiR9nyGJuk8XHdso5fZ4
xYInUt057pGnsHOFAaC421lH1Iv98EAwO5U2W4S4k8TfHGZFF8hMm5l5Xkm+qM8k
u1iI2UmxK+HzgZdC4oIGeEnFMxiIjr6kb1HlfrYztKks6su8CBHg6S5MbGn6qWSP
h0KrinW7mj7yeE/GfwqJfP3TlZWb9mzau04bpd1eWx4thQGNMnp7Xcv6QNjlBg/e
lrCackxO6SLY4OzKnNeFbLt6v2PCLY+MWaZOklG8EX2zXZIMg+9A5cq5bCvoU1Vj
EKlSHqQeIpCkUym6emeqlpHpd23mUDEzBRFAzBrj0/32wmqDMdmJTc6Sq44FacKw
VmYSEC3YYntuk7NfYwM3eHyvYs3RW4yls0F1uoze7bPZfAknUQxhx8C3P9++tICM
lusvjRRpykX+E8TJTG7FwkbVDzOsy6RPtWZeBr/J/wj3KF1MU5TvLZcFEhTwMscy
Wt+BqINsCWnPOGQAn2caFToHMUoXIfJSeS14zyWnXa0ej3iR0YfZ8dw5Hfdj904G
/SVLdtzwq7FahuC2ozBYub+aQs18BGpWTGN/01yGEk+tDwkYeMe8cu4mGf2wJTiQ
gOPI4BchvrzmyoMSeie1oEsmXqienRXWSZm1a+97AjvAS5RAr1sF0AQ1ql2BEenj
LRCxuQc03VCZEnXt1anvnQ99UNDV+jZ85zdYelxcxbYSCP/w9b05O7UYqHxlbQhv
HNZ8FEZBdPSFVjhguZpv3uy3D3GbUZvUknvO2NJehF0+h7NnD3S9e/fwy6RV0lUB
RNzImthxrlKJZSkUZwPsZd4/OTYIAyk/CGVkYDmky1ofiYq4Cr3P55ZrbiosnRfp
Fo6vtL7dGpr2nbZg8jfHk376iGN8Uat16Ia0xUUSbMmN5vwMO1mbxXmx+ThXWc1S
G0up46nRTcdGD8bmETJE3vNaSm230u2UrKfSLbqCXtTtg9rpNJHyOA9jisNFFrAL
tECTRADdnKcHnmcVrjYrv+lQhbL+dnuXsrC57EtvFytdM6Y1Na4Ka7ysHWSWLQge
J5Hl4KeGORVncRn0D+yFXbdWGFHNGVnsCArsgtkBdWJjVd+8tbQNC+RywNWFQwkc
Bp12YW/EPrIFgLHW+MstPD+AD5HMgTuZbBijpIQIUMp0iJX7zdaXHyeLxme8IgtF
dobfu+FZo+vnxNAKcMRkW+OHf0uoaLbFJDowNa0hT0o08V59i4BbIqckA6J9Emcz
RsguDtxA1d+24yWi7O+ANPeCE8WqzBsKBTUj5JeNTvW93p45OUtwQKhkQpqx0qUS
jH+0PRG1hRsjdjcfiQSvT6JM4UJyayG1fYfNrkl7Yt95qfFyPI7W6IIGXwVolzd3
fmBjNEO8f/G5RFlUvUPqP1Eg6RcCQBYPQQ5Hnh2NMYdELsmw5fMjt0AF5EW66azf
HjM1io6WQ6Q6a1enrKZrZxILuSfQvqQp3IGqCNAACyCLTCo84xxp2Ep/DNT/tcK5
WpOiADOu3yso9PlOyeaC49togCqjR28uPLv/9Zndy3uE0qkXeSfIzbbcPywgI3k/
N5LSD9WffTjtEom/u16BuV34XciA2JkW9ReOLM+yOyVZcJdZWYnwNuJpzeYFqe1P
GubT0eg0sW4QoTraT8Jq1X2O9pE3ceqA4HNUW/BKIPp/VYbBbIND7ucsTmhzxtJ7
iLLhT0yZlFBtpEAc+FYEVIA7AnKRzbtk96TNTij8V79jC5uM+Ml65cysRcIJ0J18
05v9snsADTQYE+24lN7br7ngAM3HlBCxsLBadGOTpE1L5dD0URV7gTuteR4iI71s
Q1Ix7kho1fR8fUHzUqJYVLZ4m+yDfL/zCjnqzCQ2QESa4E9NlmzZ5ucy8cAj4cms
gaOEU/bzKsmO5qPEGo0wk2b3Z3k0L0pBpBU/2x3GOaJ+9GocvyKlaRv8O9h2xogm
9mEU/2Im+4FBwH8ABEyqH/AHLiHeSfzZdjt20LIOJ6WHo7wjKz0jRP7ucAh+cBmG
IA2I8qSyhuGo9+YmSuCh6Ja2PV8DQQvYTZB4Zg5zGsyopAhhkkV93vBWpIr8QLwk
tpQu1CzFxfJ413S1N+fTb28Nw3SY7iXojaigJLeUNgRqK4vSH5rqkuPzBbaPu7tc
1LG+BeIxToLjKkA6YOh21q2VLow8kw73jsE1+qph88Jv4tHGmdCaz/P4TbJhMbjx
IFUTz0OnN+bMoJTY8IEEZolc23YrwUX3MGF5isNxG76FxpAvskkStqXCxpS5uXj9
EMIeiTzs6IAW+egC2LR8kL4jyLuG2PP2WzvrlS+pNopqMw4ZYx6G0VSYV9+GTOI2
rR3xNHs4dfbAfvAFVAmCpogvD7SiVMzS2LWQAQKvKLtDy+6OOo2AEKIQDwcEyJY0
H1tYnqt1oa934jdlZCl8d8F5GtQj2Or8BKNeVN6fH+WxEJbzGteMzfTnL1fBzcdv
dn5szSHsAR6+P8Dy8tkhrGcqF6plnC0IUboITCGFHDoxU+2jFbNLOAG3+P+xWLg+
Jo0BdSgLxaIuba4o9qDQ+T4ZY/6jQf2p0tRR1t766DuL0L3mSPVvXXrlUin69mIF
WDaFsYVFG83KA+zHyfWhGF2ovg7JKGhHInebNvyDMW5pf84NxST8xUPUdlG/eiW5
GrKw7EbfOYW73SCRFpF9jwdwLME2yhMlJmDnb1sRbOSGXol80j9kPkD23Zf0qmcJ
sw1IxqryFISgF0C2h/mNKrJmLg6WeSDpFxfNqOV2/ABtJCyN4fVEO3OwXXX2XHyf
GiZOi1zBFxIocpP0ULcyx7DQ1astO/TJKexgJgRMe03OflnwZls0lQOcI3P0rZrv
LyHFwWvqMb/o8Y/71j36KHxQo/9bq3JP5MYKKuOC4IFq1BGNnXF9ubZRJjtomLmb
+uZoClKC9N727BOR8A4+NbBuPibdZXnqim996QFAEoFWL4p9I1J1VsuaE7KZiQbZ
j2esDppPYhuHK46ETANe52CZBV74YvyuOG1blsKpUrznuFNhW+Pu4ekQ2DcsIfRq
0MwGuZKAD1pUh6ztagYgukRtIojAk1T3CCw4YY73YGbZhc9Weueo78fC/nXx0iFT
ZMrjdRO6smOmHe4vjWfUBYlZIL+mLtZAFHZe/A1MMJSo+KkEaPHkWVxZJMwS+e+S
U/M1MVoGNBuVl9Zh507n09K6+oyq/8RSr74BNH/RgGfbvBxq5Pusf7VyeCUyblhf
zOwsAyOZF+YEc/lAf10QkllSUOxPBW15KaArJ4WNCK9Bz4kj6ATvB00axODYg6l/
SVpUxSkSfFRawOeJ1x4rm7nsoWpftslC5HJW7l/WAVA05vg8zSStZx2imTb2pTGd
VhfC8vMQtiDmgxljuLYZVT7Bq6hQ/fZ2wF70bNwbnav6QfNJ+NAUJx2kZdBC0I9O
oCTBCCWLc72CBIZVNp3p4GfdcvDAiaRu2qVHlizixHSFCTkg2VpYJLeVykU/yaGy
OVnPrGE2QygI1REYn3x0msCAZfb9VyghnlShAKJz97dFLEWxUL1FZiRMq6A1ncD4
zMdLkzh/tXn2+Yy/dPhflSSBOpEQrllrXWJYgiaFUXF4SIzbafy3guatt3+/GL55
pC2tMJldB/PwjTKJ5hP+xTO7YETxdfCqdeNO5YHMq1hWnx+mSLN0SFmKsubrsXbl
rVAUmjlKkX2KPdlXjciJ3MXZ4D/Bc7/klY+arsnNfjfWF/TIz05ks0KVZwsOnt+t
h47L1hKZd7Yh6w/O3uYojeTrg7U2Tm8/6s7mFidaTOIQhzipAbknIb463eon5xF9
y3yILblvI4tVsn+Twl2bimEPf6tNG9b9VD3NfF8/pjjKeJJ0qxNyR3sSycu5fD/b
vmNWoTtWXcnBEBXDPhksO8o0QY5d/hNRJbb4XVgSLsj2R3h66eeAJecORQrHiuD5
dOnbw8iJ0f10uZFhFRaMF7cnYr6q5ewn2va5u89mLH7VC3hi1DIRvkSfSdm1Ag71
Vn+vlqZ+Sq4paodH+DY8WX905dgGzkYzm1aHxUWIXbUXX5YmSl+HWJWGh85nHloI
C7qrvKBSEkcxV/V4J69M3C2ZSN8VOydF3SyHj+B6zgIsQWWo6I9UOify63w8dQe0
r57mRm9bsY6+hjDP4qPwusbSxYLrIK6T2US3lrQnx+CTslNAZ8n+Z2ahIaWmkOkj
yCiSJDBdqtMZjkr/eogz8A+e+4K+U7krjQFLNdR7YYsLHKM2AkT47y4DfNAz5OUP
Jmd6NVeBQt6SeP3j07HQnJ1rOzvPIr3y26Y0OGWPatYZparO8TD3iNjTNV7DAffo
wd5Y9y046HoBUOmX5cC7pGVgFywF9gf6bRKScJSoAyEhLZqoJ3oG3f57mgbKumbb
f2gX6Ln7vlDGWSYlLvRwZha1490JvYQbfJf37hw0rimq7pxo+8rpWpGziBLSH6iF
V1VcNsYd+rlN+4ScCzCpkmsEl+Ckd3p9F+s8kEp2EAUrHLvlpN8Be8y90I7QEJxX
4JxxmWnPKL4TQJ5tUkXDR77wfExgYiLNS0BVCV1dvbfT3WnN8/Dl+to2H5GgjXlO
DlXY3kHOd2+8+SRC6CtFkUSRZje+GM7xGDxEWWxyxH2GmTfjBUibmtTc7bagSW6x
18LWT8kX1WdISRvSc41VYv9r0fVTCxjQZBuLvHX6dEFQB5/EnQewmc6B8JE8huds
n8jG2HMJC/o9v3khqXHhHa+9/0nP7nKr6GVfAvuupJz9WWI+zEO+yKWiAAG/Qg3e
YKaAVe7fUeyptRU/vEBZ5QZ68ap3mv/eP0dreifUkrF3zQqlBnpKavOyBH5XW9K7
fSPjdIgP0rKGtTnJ66x2WolQvfQE44xr+u9oyNQ8iI16Xee2yALVjKF4OIxubTYL
4VnUOJBzZnb5MKk0/s4m7b624sRV2qD+On4jQ8a6jufIRpHFO/arCBUNOrYjK55+
brifxZNgCrW+ObUygwsio9eJ9euOjauAj948VZU2I11vXXFAoXL8bNyBu6z1gowm
khit7a2sUR6jzz/1Kmpx0dnO9XE8+QZsRUQ/toGVUVLVuGdiFQVCwspE4fkLWTHg
Fe4EI+kYs+mfxH+fTVWBssPSY3SglHh5AF8H4hIy7Svuxn84DMK6Y3aoCGCOA68P
eyjG5LKfrUIbElSOwokkKsf+ZI+mda3gAmEH1n4dKULkOwTjTHuWHe1ebDvG1bMw
6AN8K8fG7pLpoaRuz03tjyDWHJeYeEjOwz4iMa5YQogaLOiEjU/qiH0Px4Ied+4E
IB4i9G+HRcfB6MEb6zOhBWPCfNtOiF4l/LZadsxrfvRucK5Z0eCAZoiblB/KUfoe
SBfpvSNSydzZcoSIpvRbsxKM+zv2EARp/sfJIV4lPWZezY4XMZrhLN3ft6I543xe
iAZaOp0U6Fx+zazyHAnFI4AsteA8uS9jWsuirlYYS4aq23WJIc/0hWx3O7vjuDkH
yThb6UWGjDN+pDTyythg0mscuBnyClrN8IHAYgnoGPcruS8rXUfTsO60IJF/Rbla
At88hhvASfa/oSGc4pFy0dtCOyKLrlgA7YXjtchjwCyPXTFt/uNQgROn5m68UuKW
EbYModycAhb5wNJBBeNSS2e9D/tVzHPaMxXMpUEUt2kwQMHAupUS3DJhkoEZ0sc9
bmiGsXAt6zbwXsTuJ3wWxHRRlG1dsYMA18iXX+KREL8gYfBUfkcf9TPqEM7MgGlO
AhY3O/LU84jsqdZOhJFtPsOXZhCrIKw+wp0e62TIV3R725qHPQ+hLNFHKIuhcr4A
k3JBPDGWd57nNlvB4UouxJPT9kl0D7YTowAHoJ1Hl66OwiULc8lujPXhXmcydSC/
Rc81/JUp+nAIMBw6yxZmBaS+k66dZuB1+wtSKikhcdZINN6QH/5SIl7Sn/B5my4R
WDZvJLOzJzPoAOuHsvyHtoFgP8ErwlE8MHbiymwq6r0HPd8AnrEbBvwPe5FUcMkl
DFB/QK7o9AD3GKyCaB+dsqDsaIGsXUfFn+Xg5HbHNKNQLIi/g7+XzE/kxwCZRLdl
ikGVTeqyRnUTB/Ty42BVeJRKKcJbQjYKzxW8t0OQnPKEc1GbTk+YRnaCBPHsHFYt
E6Mjyiyh3yjnqBntvp7V1hNOuaHllXRvEeDfvcyqBq63O7fdaHfFKJuLPzS+Cx2z
07j7TQyFUeAMOV7KXlexHZmDb2/2g2LfiJg7c/sJzYSqOWKJHACSk7182JkAE+BV
f1vUie81QzPRQ/Q7Mi9R7cNzpoZFTKqHaYVuNes02GT5nSFHWWSJV0MktWR+Yq7R
VAifJN1D7mVN0f983FbK1sm+hR4v1BD364jjlB+3D2BIuZialECjYMQobwEH80OE
Rn06s5AhOLgPgcG1BEjAEWoO1QzIqK2JlIcFmnD/7dIOeGSOSHJmnL85aiQM+o9z
tA0DBf+If8AF7GKstTWMniSFZmrCDn7Nz/W2t9PL6O859kF4UDXH7qmtZ5ZUkWmU
M63Pa9EI8IolkeS/G9vhDNIm9yVJEenlfITIghS6IrhrZTPWo1j17iEWGvbQzxum
4vYYuPI65jyQy11d1M4TlXkSurICdiwsRdZHS0TGEgpa5Fx0EYV5E/EKC3Vnn26w
aMchPn8lgO+WnIUvr7mYgDq20IFpIImn0kYe7bgd0aKdAhw/Z9LMXgUQ+SNFstwk
ecy6/FhJ2yh3YDhnb98nWYgq4LtA4zM5PI/VAVrYgdckDAh8D31AyHC1qBXPqVOL
brXmwVm8PLmUnA2m/wkOXwwDL+BNCcYNalSDlPl3jy/SvIPiYGGO/E5jKAhZan31
cxteKaWPEuKsKK7XF2e3vPTqs1X9hEgXYtFPelA5A/Wbur7ObDFpDGk6S4g/EyVA
OW3dt1cUFVEOY0TDsw4XTToTGt4KRc+75WaKt7slI1rA1/BUiLc7g9MCXe1YMMLm
/GSjqV+J+fq5vJIyKSZPCmybd7D3YxpZpePPKO1zwoKMM5CzDKoySMzgW0BrUXx9
+tx5UQeKvtdVQ8zWgFETegjnk7O0k4/38TIob6sXyNGyHf4cHSqMP4mhQ0NWhhC9
NFSx7NwI2WR9tuhvzvYmnEcSUfXQkuuC0RU1QzqXc9Jgr+S5jtD/qVPgxhDUE9SK
BDn8QfYTNQxIapUYfnUFk82CSG/ERWo5TIpeMZfAToztb0Bul+ZZphQVmy74+vyQ
ewS2C3RwCl16hts+tBD/pXxf9OUyLjz1T2rWnZ4kvzHw71MCoZJzGRajvrqX6q92
zBQhIdRvLNXwDAFlhDJDKBLk/LtEQVb1U0rbkeh1xlwD5/qxya65jGUBRavf2W1t
8YdxNVVbBtUGSdfUnrM9B4KEEOyik7lGvmJCU8Wla+7qCYja4dyhUJ2AkbEsZbbs
C0QyCxFrwTWWyBrbcChapO/hvd325w13y3Jm49k4X70Fhj7rCooIP2GXTHWXPpMh
RekYJDb2m9NoviWNZfFuj02/Rgf2UgOE1U1a8N9AE3IqMw3QV8sMOI+pPav29XmW
XICxUidGcK4peHvetzzbuHm4AooKQnPc+FfCIpSIJ/zvROPmEB74q/qvn6JkrSmR
dWBDHi9bVOAgPNpKj9lbtyq2tGzxWG39Puc5K1qVQR8gW9aHF8mHtFYF+H8L/tt9
YD0pQg1muJJt9Ua98pI7E7VqZfSGAnUUcHdx6cWmQWugPHB8nnismXF8EKrRQdJq
h1DVs3nVaCpvDqu/ztYfzJA+dbhXYlmQCQNUxckEGM+x+wiMj6rvRe0FPk6d38XI
BwHrRrxktbOkaLiCWz/7anX8PNTWGlg3AFU9JuvwYIy3dbmio+cgGDXS/lbFTOtW
CIxwhTWCJJ7ag+mnuQLZPffuS/CTt4o7vCS/TbVOY5p0AogbEZxoB6JSStZP1Wzm
n38CUqvA/hoEvG23vd+GTFURhmGUIj1pRk/b9moU0S0UgmQyiwn6ujkhbsSUROtG
0G329rB3ngu/zrKy3Mi9mFRTwRw4UKPZwz1OobpPHxS7PR2FOsABwswdUKSoba2a
XtcgUXzHN0uaQMd8hnd2EhSg0MtS+a97z5NSVlhvazZlXAum4FPUv/aWZsIp8Jb3
F9xoYZqVYgH1EkOzH6oaMg/DXmiirpjxkcLEDuwoHtlIufRBdvieO/8JuFNLPEdu
p6RSTNKYrsp7p9vaqWZd0hSnjvSdfydyNAvjADCtRdLtUrZ5UfKSsjUOahH5zA/Z
en36TBS8huY92uvv4703cVUyohRuiVEjd3J3yKPlunCk67rV5yOP0mj45+jDbhoC
ZiRKE/Jl8KA/A3MKs9QX6BikrgqWyWspmvhkr6x3l5w0UN3HckLz1YizAJVr5wAr
r1C37zUCDbPKph7rmlqXYUjLescLhGCeTO5gCH3mbO+NW4XvnqHuzm5upXZ9vslU
+tEKZf3e6iQckE9+tnzwbwAi7uIEfCeAzbMIc5D6H8anEgEL8zTemJPCgradKAEO
jcNjFemPRVbSCV+ib9fmw1fIbiJm+TuJlQhRRWobAfVfMxA/zc6HgR04bHzv0X7L
M6L1N3FzD/moKoHkjQx1a7Gs8FoMHSRTlsKEX1rUbhWMWykgpfeN+8JSoehB6Rtz
C7zbcAWXVDPPN9DzN81Y6G00tCvBB9xsgtAYEPnWYvdjjDmjN+4iQ11s1Mb8voaa
Vy3MogQ0mDSUazsz6XG2NMnlgb8sbEeCoJRsaSNecz87SapkNvGUmkAIQSCz6Poe
m0hSmyDCLxVNpHxsyyijsSHvjZqw2ZgZJi7Wd8JuYXeYu2rawRhMx/jTrLM/T4Om
U2ae8p9Kis/0EQ5NumyUOnPF4t21JE/34fY+HLH3pKFSJ3h+pUZD1uwmoJ69n/Yp
tW+ITje5LnRUfvVrMlfEJSgdlP+1rbT9sy7/f9Ohpq2Nv7V1RSByNhjaMai/SDaT
oKz7SsGdc/jR8Q00UHEz7nxSaht0bO//FNOqdG5zffb8sBIOxELvUaQ7Bq7o9bJ5
tfu7sSDrchDp6gLlysDTufBF4rqyUptPD1s6Se0V18xE/a5hMATCDDPWFBQmC5M7
mo3Y+Cp+dK5PVnOtPnvUqR17hnzM2uyAS6rXKt+6J73gnkzIjokG23TeFGY2S4WB
jh3ZCUr70SQ29nPLeq2o9IAMvSPIIMbhtaMIOzrh5NQd7QHLlsa/AoEYfNV24EC5
bGIlhkAl0yJO29z8jR+pPkEyeh0nMGXnVmOFLi4hIIF7RKaKjvvOrSVTiF8eNOnB
aozXPz5AzVSyppy0P8Yo/0E2tzfIkZwL6aJcQFHaQYRtPsxjDKeh3TdSygYKxLVm
OTAfmjbsXwttnR5dnBc1yI+a6Hsa1A/p/ys7lKt6aByLuJRSGQxYeg+jldAkE8a5
EFr1VGTqOJrcKXaRipAg7Kf7r0IE94xA6Snu2xCZ+H+QD5SQ2eGo24EEw3opj5hE
S8zL8XwjkkxeLeFSufjuq+2zb7y1vnYApTJ7ObyZc6O5nvl1aNW2gMaVTGsAPNRV
tk55YkbQgPuE5+AJ3trS+GOC+ZlMyxtxCQvb6iTsFvT2phRJfSiHEEw7bjsq43jT
c2YS39hfYxBmTjMdBK1mTtkKxg7llHWO2KqKi5+IygnivXRjKbEHwYi51MZI4Wnk
Re8cyx1zhCgFYV/G5M3BGU1rfbb8pHL5sY3yT2zv9tUiRo8L+mQPKgRR5i9JfN2/
UMoqXhIGe2ueRub4tfcZ+kXamvX4uInk/vxyTSdXlK7cgtXEsXNjSilHrFeEFeSz
kFLoraKxyBlfTG9T8sEFkorHgPGHtpGJ27adQ0QBMOMI2h05rHIxR0NEEvCefizB
B7p0SY5QhVJClGJ64Yyk265yp1QA89q3E6YnBhvuTb6UGdVfVesEySAKFSxVTc4E
876zJYvC8i5eLmb0L6mcPWVLw6F76WgutWUZgHSC8JSYBjoImk6yRNGQTISvV3Pi
IBfFkxhLJsaPz+5QAYyv+5mlHRbiI7CG3gnUwpv7CwJfTc51XHM88Ur9RdMJKCTK
zncTuEcvUipusuSFoTElDiJ7bH2ZBBrn5ZLsA0TNRaJYmdtCDk981FfZ2I2bMz6h
4ZtBobPxAOCzv9e6ZxLqWO7fodE5xLDbBMlFbyxN8Jepmig5Uv2F4YkTAD8V1W5d
jwhp7mzmSwvw0zFWc6EHNrwkdkS28mgn6S9SlsZBRZjNqjMuHonrzjdkBLnHH9e8
0LF0K6teG8YCoxd2kdlB19//W2LLzI9D7tgrN/haB2Vw4mx7XhaAzfAsfgyLBfKK
gINTU9mXV47YUeD2urDwCE3jMniOhaU7LeI/vr4BcPIrUBhDSWMlARy4GF0zfADn
BXARN85zKV0ba1VuB1OJMVXN94rmu/+UFkgA3NQKN12p5b4i3hcI68LLZGnT8mDD
AfnoPw8PSWeG0w3iygGGMab0+pFAeFjD6Uj79sXNWTdQki0FtBFQ3k2qzqOQGjd6
Xp4yyeSNmhpCqTm9+GzPNJjlL+BZof1CKBZYlWxznc0dniUK2jKKpssYVMbxULcA
5VaCNcb2GYM+IYpBxaJI0J1/p4VhhUUUZLGjElHd0jSWbYnDGDE/mfiFWe9djOtd
qE0ZQI6itW3QanCOsqVG51dVC2FHQYDf5pphWTW3axCOhTey7+/SUetxKLEFJi2k
DJUhzRvUVGpqDTTDn1wMLQgKFUFHY/sgOojcsGReIWbwsmu7K/5FT1LgFlr7UeWF
2R6tqm2J1mR1OGbR6PfeQyI6SP5MSaLeuJ+PWz0waPfXH5kL+0G0yIr+1j+e2LRH
LYyLpJ1Oz1u5qB5EjCNwoc52YsgHpRsm80saB78hOz130QcKxf8kk5d3cfhmZIuk
lrK0dUdbKIs0ywozMOaEfomfrZYhPUi1VOiKTZCalEqr40heIlF80Zax760hpdEa
682qD9FJ0b7zZe0mcbRFuBwaumdwqKh+CH9kzcE4isz3JXc9L3+kIU73JDcF6aPF
muJHiBgWXC+XEpO9IgboYPeJCPQmWwyIom6mfseSogrLGe7pnJPlYOH//N8znhz6
HRvPFrT1iiOeunqxweAX8Ra53lJUPJBHIvfjDTU5HNAHjn0qdLTNnLomQHFtWOEQ
rzIEW4j5dPc+73b9eS7mQ/iTrq8HRMtyGTm2OiTuiHib65xAOPhJJwgbFE0iNVMk
4zE3axmbWLG14lvtOYdBQJXQEI1vsZDJIA/7KxVjCu3mHcFuPczJWjLXoPBSMxLg
OY8v7k4JpRMyrrJfK923A1Sr7/shpDy7ruR1c+O4Vc+rVQNL4uwgqB904uG3e7Pa
0vWnOr6cO21eHFiQpqKwu6HJ2mBLqgaZm3O2/2WEBu9kXi28vhVRDkZKVyA3q5KA
k+ght2gXX3/4KYu+uKS7yv7B1+2Mq2hW0SYg5kTunvgYrhaoQga082lF1XS2gl8D
OM1ntfJy4rq2NiON5aQjwPx8azzl9F0gZnZg00v1kleMmbsgGRGyPA8q73R/2VJ1
73THdp2/smK/VzgmoBTRjPPmcyAeuJzk98KJNakScLfSfy67kqORn2kVDqkYKdS2
UGD9N291X4Geg2jhrDItW8N5SEv93cFgoFZk/EPg79mPcHBBtt4uav19ePgN456A
pbMVeeRoTPY6DgSEc/8ABBfuLipcxdcUcHiUMVrJo8RKWx1qfNNs6XHelly8S6NB
kiPIG7EpC42l8E9HmScOISmax2cUJFfTV5h6AgeOtKkkYg3kYouRyGIelz8MVf6t
bx5qlE3Kkfj+vZ09/RjVe5xO4NJXJp2Ar2kgcnpqCLbobuVPQ0hbZyecW4iia5Y4
INyYiJrU6Z4bPTpyoPhGPjCHbXsb1PzZzbfmlzF97BTo3lvnKiOklimNPCSTDW5A
gMyMXil6FegXHvnYaDh8/Zrnozw1Stv8uR97yhgE6efD1s7W47yP7iSxVCoVwBpY
NUlNbeMVMMCDApqmWRf1PIagmeD87FyU/1luukiMFCHTQdl7Qz3QaEnCPyK3xi4d
Vr//qKIwH5aRLmOby56zSUbZvuoCzwchUOwV9/MYWNEZ4cbM3mwcVZl9dGPw3ijT
9W32584inKoW0DudSjZbCFla43N7TiuNG892mVcpWVuhN0ph7Vje+0HQTc7DD9N/
Mpqh4vqngFPDRjCjRZDzHD3Ixe4OWOXcZjreCZTnyQlj9r0fwSKvIRQ7tQ7HaefE
YOZRgX1+KRUV9CgYZy/Hlx4L/aMhRYsJ+4EOh5GdjrA+HMTX65B6XojT4uKpRMsF
YcjS9JfEdcMH46zBBb1ee31CM3qHqV7KkzaSYRh4z971DsTc31ErUcKsxDGcc7x+
gnPqahux/LzHFJyIOAO5gOdI6YK3xS5nIPvbW9JVjELDyiCnW8qD64GwOh/Z/D1U
gB3Ppc6cojVf+FeKE68z4uw/fKGJYzIkls0OTOJVq/ffkjHtKBGzixPztYsylXlW
pUQsYacF1IhSZms9KtFvcs4Y8fPKK3QyeajGt60Zig5TRi0PYoUUfP0vKwRiCK/w
GqD7UY12aYjyvG/r041IBi8ouRzeVYwrU7bDBgbLh78DnLwpJ4lTIx55eYdMYswJ
sejpPso/Yc9J0Yy44CbpNdzo5kxFCGWBLfNnIUfZJOQQyoQB2U1wCBIAwI1hhE62
zXV0FOZVeVDEiLGbprowgk/gieIjXp0PXm2zXRU5rWCufNcz54S1VJppsLqYHA1f
71Zuu2CwCBGu6W5tAcXap85ZyrN5IiDeohnBOFpSfJlMAi3OW7mS6Z2421vILEc8
QBN7B8iZdTCVm9UyfC6w+oyonIVaS3B1k44kz9LGTMtwXyF81fF9lzYfK11L1gOq
YnT+rjlQtECkzOVVcBjJxJwyeaVUTjFQyQTvZnV5MFpUR/Cg4B13kleqjuTeLj2S
tvfjAZ7tWyeNIHVR/MwPYSIVE5/P1LkZ+pvlcs7Er23+pXXdCeWvOpy0uoaYROCP
wTcfYWuZ3zjeAAr5ZZ8NUxbU9EIdYr8xYAnNBSCslbNhhqBNDGYhPjTw+dxZj+f1
FoRPX7fKQlK/ypgwDC/HtHaBErFfidL2JP96SButCj6x36i2d3pvHfgOsB19/Ljg
aQXeuO70XaK7kZLOGjM3xih+uBLk1HPnUjz2CZKgkvW3WLvx3hCpr7xvBfAtofPb
xFWr0q2MzgIXl9R0Q608naA7kVR5bRhIXqTdXWArgEyVudNWpJ1oQNFY7ZbGSyhq
Mbd7ax6GsQ4pHhhxDYSfekKYeb/Bk2A9Muwb3c+jiEY7UHNMgTfV+Jr9E2gXUkn0
qrpMsmCkJBN2Ob+L/11rQ1TgMTUhQyrsG+TrQHwErKlXFRrNzyqgqXHan3nmGNYs
sRcCB6qUQMCic9dGj3pzS3tL486/NdFx18iriIfvLCeZ07QoL0wgEHGZG/cdZP8+
DMrDTXw6/50DWLUZbBJzHjXik71S1cWloYTW5cfa2oZog4PcUqF/MgcV+u/KZ0ak
jClbrquhPowyjnXILtFtAxtkfYxyVzi+9QnK2rDgbqeyc98LoSD/jypCCNVlIzQJ
S0R4ObaRtVms6fZYFjEmQg2bKxNcUWiR187AtAl0A1IBHTHYtkI0O7BDK1xMSUGu
KLeYfjfD1UZiJK3oAY/XKEPNJUVnrd3ygHvc/SoDNKNkjo+YnNUnwmeSIWra+PcQ
Yzk9g251cXgVGpK73Ro1j+ScdCR2RYx7fhXRHwIynZTXlT46rrpQGKFXjpKueXVs
a5yL44MUn5E67mXfwdfONstdKnRCx16HcOav8YK4896f1DxAcghA5EWa9S+RCQtA
EI7zxrYRPIK9Vs2c9ilEU21xx/CrK/K++ZH5fHJfA6XbPGDNOsyjsl7rLD86ENWn
qZsOwoVAQrx5dcpWygrDcPSxOl5m6KyIRfPdOYGg9VA/1zMS3OOU4ZxbQgy5KW4o
R7vYa4tfXkhKzHWlo2azxkg3AbCcYRwwvvqBqK41pOzwzfTJzoqctdP1ujuv1JQR
sILcoSsshBTsJIVCHCGVaZU9ha/39Mur0tsaqwLlhXIg19t8U8A7sX96YdxYxEG+
BSrnAbAehJlv4e4IMlXFwzerv1LltRKOB5rxnTdsMfohxa3wgO1gBdT5g3xBXY69
ega0tBpQSa5F3OeXZwrTcFvuNt4cQPGCsucc/PnxExJR98ZOYS/VtVVPFDU5guHg
NqoO5LbGLD2sD2kAywe3N6ws7bR3Jt1p65W4/c2V1neHKjOHH2ss6zRBzk+kZJkr
wHIuGubsE87t5n8wGeG5mf3hEZkApshLXGjzj7bUUlkgopWBul9/6buhJ0pxsvMh
U3lg76xFIPoYCZ7kAex4Qx9J2AwFWrC0V8hvJOGyaUYtRoVcpZQoF22dMF9RxZS/
E8W70qzp9PAyFDB02KAZVuem63tXbBwWddmpT2XSlFw2DuzOK+GBvC7whfCCoy1J
vrQyibppt1pU09qoCyZf+SK6gfqxaLAWg1ZpmFcthn7xc9fHYWqaiJt96JVilJtV
fA2jyladep45Qvk99QGfVpdnTrqa4iJRgZDz6arXUZeJBe114wvfupUCUxZ5wTF+
ym40g4u6cJ9XbRYxw8YiDVILif3ekt2Vn3idqp1GDaTLKJzJvJCR5ijXhukjcISQ
gPogHvNBLDpKIa0nDM1qBBFTKJ4Nt9wnUi+3xkZH3TcAtY0SOWa+XbD52vtcMi5w
RguHkwr38/j5VOeIlBV1xBtXfmVOAU1RANisa7UnxeDtMMNo7ZfeVneTegN3MYHl
0AHnIU+EcRrJjdA9yLLGjaDdDo8DycssLeg4WqPPTFhhK+zQBy2TJPHaVkC2rNlj
Uvpq8yE8Jq1CiE6iPp/xFJwXRJa2Kj5pmOH3hrieGPZnRK4qcdel259OtOCOWaTk
v8mTUlWLAiSjU4QM/XOun2XCoB+2lcxxNA/f8XucUl+PnFjxg49eGKuPSQlxJufD
A17Xrgpn9p5sly7l/tGHXqRpabr/wLtZ6iPt5rVF9m8a6CkvbZhKmLUQl+l7/90o
quyuDxL8Y1y/GEWxNnmVXzYVV1SdZTmUFMI6VWVbpd+Kur37483maxyJShOU56HX
hBlUYVrWXukogex1ydZ20KfR5NeHGSya1coNdtwaOB5w/RN3axxniIUygr6vRriN
NYlpdkci8QfOowxE4bmR1IR4z/4mCnAy/Y4ZPuEjFFZFEpJljhRy3Mj/fUJq6wGZ
MSK8Ue7OCLivYJyV3xm13NYAP3XJhgjoRw4d371L9WetkYu6yoGzvZaf5/9J/Sjo
3FSxVPnlIIPAPvqEN578MRBQGNSAeESLuAyYMMkDf+9FxG+lvNhiHuZWyVv9bm9R
H2dhcy3bgYPxvlZN7Um5szGsybcvdg/64FPv5G/+0Ht6aGlcQ43yYf88rbuJ9BvK
33BOp4yZIyN0ZJIIiXS+ETAu1fvnUa1XmptCmYxpRYiXbKitKo9jDCw8rjyCmTi6
Ul1N4A6RDcCJtvnIM3n3n5hMXBwFDb6J+zC4bie5uaKgxkQwRzcrsh64kbiZSM6b
IRlkne8tRB5ebP+fE2R56ejF1VExk1B954ZRvX2QbMlO4NN/R/sjgTwRN8Gixdax
tDA6LvzaMwHq8TDDK2xjBm/Z91SLD26YRvrerD5iizlWpocBOVr6imhsVptkaeuv
fpy3tq5F7BDwKVFTz+uRRugN8Op7bTyZKYUBX+JyWWxcJ0ii0jqcA5r0IR5NlG+E
5WluLfZp09zE1UMIb+sveCplfX2wpJsrZPv5Fh+t0tlbzF4CdUTGwkuDvqgnHJoA
DzYYG5i/AEr1ytp7/44JqlQtIv81bDTDlcFdo4ctmSieeiTLjsCnQTVajbV/Wp9u
OO4juCF4rz9ZunW6Bas5Qtg2M8GbGJfCVFIkEvnh7TQNT4l02zsumSDJwH4IepX/
awBax5IjfHjZnwBTZB8S6cZn4ObDi9+nryUNkDQ8IwSCTHSf+JsfGJ7ZXPmQZ/fE
bCdgDoOB1euna6qLok4s/SsuT5hoSiFdsj0IK6VpmdqucghJZyQpyPN3l65Q3YOY
DWbc3JrykUNNNz2iAM3phuwqfZSY0aYSnl8hKR16EosuIkJP6Jy9xZ3ROj7IuPZa
ZO93JTHuXVWVATH9czF97pdC5+g76j1ldgD9fdvuOxrqPSc20y8RSonkI0vAjbp4
3jStW5WF7HzLx3FyTFjufndDA4ldsdZgy0a9lvF1otaAgMa/Kau/vopqoWIK0lJg
j5j3MkzrI9inFhO3zV7QdjMt7lf6WhfvkzQNzrFGTKt0Ycr8EpX0r6IIk7jQBnym
1EBS9zGIOKJ6Pv62S/oqQ3A80+u8EdNSIP/QPWlub8NOJgWO96O/VdaDBQm4dwNQ
juKI1/7OvvVBs9WjFm5SYccGUJWFDX2WGgXVl8HOQhID3DNkv3VxsltOyAnx7WwR
8WZR36eZFBS6sRVYERk1IQOwEpYOTRLoFC4g/p3jxbfuaHRcp7slKQvp76USbCKr
7AfSMQN3XzBZ1k53UMXW+gRhQaA4LOIuNnHPhunolQbEgSwv4dOfhI9ZNLKtBMDP
2Ie4cUb38ItKJ1apbv7oPSrgjBNl+NP3REx/NYq3z/WD8cd7LCOzquIMXkOZlI2c
gHwR34deGLM0U5I0LeigiE+cOT1xt9CEyALOabtRYIlk3cNO4Bljxe9o4EtFR1kj
DlUkpaICl5v9XY9Ke0HIRhHckYApKwgPAZt8A5FSgaSw8FE5ww2LmOvqC46TSqG3
nUnYIfpKRszNj9owEC23XWGwCMUrzgkw4sXrGKQf1TMk9X24bdOXVm/AxcPiB8Ia
4596uKwLgCNQACpoIc/eYAysQbMuWeT73TEGK/tJseVbFLI+5/SMoIm0U1zV+nO3
Dbg8T46kLosElpFeNukdr+bPMP7uA2o7cs+Ag/zU7mOE1QY51rEr37oFrBoJQDhx
CcafLbVJFHq26tuSybs8/vleWTs6UX/x10kHmqz2lJjzBfOmZ7gxE897x8WdidAl
Vb2gyL3WwTc1jAYckNEaElXogzkAdnZhqsP6WPI1xpvQ3HLuAHT1E8DhH0wLjbrc
2hJWFR4QA8O9nVSFvpqahYSeSSW07jT4jhqTALiylTPZZzOsylWGjCwCeCwlPn+s
VMngJE3b7WV7+UqAYu6g0acaeE0/zwVClN3Yig3My27pLH3+S5gcFrpTBx3TWUm5
HopO6oc7N1LEomAq+mxn8R6HvXa+G0ol4TIefNIOiThUGV7dAVJs61KEErB0pVxk
O+CSNiE2gxlSuc3kclXsAX5DnNyM2egvHEvQ9O3aPdaMRwV183zqG//s1kGzaAeH
HW/G77bj1R+8EdpsnYFUtzIhRUHqDYJbLz91DMQqn4RMyZEk2fQtwHPG707Jgh3t
o2sJYk69fDz1UfNlAz/j98aLqA9UY6urOQwmFLpKROuBhwMl40I7iHXGzZE7bk57
snqmTamoo+KeFDagr6uxbY3XZ+l2Ky3NIwlbDgsU8Lnt7+V0TcjerlILMSu5jNbS
h2ShFEtuCZ/yUfw/qqdCYprzQx5MX8CBiwL2rz3q9Cqxh1l6Z25aw2jghVRU41g5
+7cKw85WkyFWfqDecjGq4iyK2v7Jqa/70YJlXX4I4z4XNym/ya9XS4kDhyq7khhC
xt69VXO9yLWO3+nJZn7dKOEnIiCyEbQt5RvpNWWayaJMVDY4cquOCn/f03IZv5Dw
N7+B62zN3awHOMbn+DJntlU2Y4Q3LL2AMO+N0ygZFDsTJYc4tlIS51Wx+6ZgJRVg
UcYRLY/tL8yfonqOkBQUVeH3iSmb2v13asVpTunv9kI0bM1oY8GtUWe7XXPXAIXt
1z7w3tB5vy3oAgpqkR5dCIPGFhTF109UxBbOicHUQ37Xor5w5WqNNjvisNQ4hdmr
AMZ5790aN3y5Lzv6meByQoLRJYXZ0fest2jtDUy+xm98MoCqBAwxXBhoem8iI3zR
AAYYVxibAg0BlYCBg/YAa9y6bF+RCk3TXGm0SGkzo60GiW4ebIMdrU/Ck7IhEKcJ
EpbbRSOaqKpva1BxAvvkTSSSJD9OlGpyCP2zhMLy4HDgF1bDQq9P8ZoNmCzaPWG8
C/Swlr5zK7r5EK8Aa5ClHzPpL70wazIEBKSZlouD5/b2QcUh1gdXdveZqJNNVEfB
Oo4XeN0/mXsOzZrcez79Mvwq9GJ551ryEfjDpWSQhSicD1sk595MtklwKUYeMiUD
F4cHE+B18Ibv/ldZwgZV8kh5m1rfwNIVIAo4cdLmMRO7M4eQUrao0ybBL5G9LnBV
qN3+V0sS+g2st5HGC43XueAq0/dP9dQ18iAj55N+Hs2AthtqRvnIn4kNUL4jEYnQ
vEM9F0pRaz0uHKGUYW5PvxUc5Y2vWiFkUT02NpMNgL8qML01k6JpGbMSpIhJhiBG
rOwTQ1ySIvBqkohkZBAzKM8KyJf+gEj48pEqB5XskkR/iUEokIzMMXtGt5dmbSNB
MVnH3N6zbDDJNZ21xMybSPIS1l2S3t/knS72imFx0YGqC0yi/h6z4fSgSYCLMQyK
swfzKZ8RvzUB1Aung3JPfTxUnANW4rxL/66LLaL9q0LZ7BDZM5RJoIUnbWwoAbFX
2bKHI5CGQhKO1vO9QEFfHcTrQEWRtAYtDupmwP5UXre/+WP48PdToa4xc+h6/gRZ
dD4X+2FcQxUs6KG5ENxl9B6PRAj6ICFGCTOjhxjQl4FGd51R7ql4M6UsCA+gsm6h
rG+mKiX9Mw1wp4BJy+jElofSQhGAprIwmsU4OanvaMGSThRRbp7J3kBj9U/scqvH
5RvTid7ZlulhOu/PG9FTagPrn2Fc4eQjrCvX72diGA6PFiIUbef3D3F5uQDk3g2u
+4uXHM8ezQpE1McYYn3N3TuIeF5WqNn/HNTbPT8MMbL5wyJ6XswBae1j2bAmJfvg
DYtqlpqLslnjb0LIyqlT+VCPKoTgbRBEVuLmUAZL7pw1YM/CUzbPum1cZYWhvg3Y
f5Im8KDqPh0WJDudfHZemxlBzhDulZIqj4Fp9k+Ttp+fUFEZk3MC3zcViyni+LP2
6S7+fEg2os/56fKFMNmqcicLBVc0hjbS2ZFZWByigSYYUm7pg0cRtOiIJELbz+En
sh7+IIKtaWv868oloNq2xg2Ne6VK7T7+Pj780tfdQPTluPfx1wS/Sd3Tyw85yvnO
7XExnmRzxJ6hgnEfs5d15lS6zjKAgUbYqfIjE+Rb87M0ecHADPjP1ToC+NAqEteV
57DMHiYLy4NwYQDj/IbG9+yqFANVdhmmkLaTqh7UWTXiNSjiPictew3iiTSZIGXk
xZUkgRCq0xuaWFo5q16jizXpB/y9U9CSWu6/7+LwJ9V3WkSrK86rJ+M/rdUGq3kl
OeNb8Awc2AmS61TuF/AHIrTzj/bblfWkqM15yFxKNsE5CdQUkFiHlvxy8ZPH/mt6
bh353xDA67FR9bHxnUXBWMHdiJIlwa799hVMMKjWdLthvSeOEKyGdzAhJLsSbIP0
5E1BmJFn/NHx+iYHMyIhiV6kAj1AgTO8fbbIu/MiY2qul1djlEuI/8qhVCJTLKhd
iynJKP3LrhkPAnYFqRAnhKGB6Q/znT/mJlDafKBvFm70MRWCJei7sj8RYgO/sqRX
udFX3stHcbOHHzJ4FFMneZxKUn35yjN2l+7f/rhkzo2dz5szF8CgXgtNNheqFmMr
rhcZSgacOFmZT+kdr9aWFiuN6suf17TzbodiLGRD0gqec8yhkHAsBc+M1ZrD1fs5
uOxsDqG04lTFzkz/u73RGhWf3vIHB9vyEHRqGhOGX8N3R/C6YsdmaejlUJ8Tibvp
azFCVKVgWyUUG67hS9daX9rsJcbK4jD1gaujFQZ2NEksmQ5utIaVtbLNqbZSlSm2
LuwRh7AuNczc/9wcGsgeJAwyLvmL7wIVxamPkS1hufCjec6NorLBOHFvLfqkymfl
EfZS+mHSKat57Et2TyF2bLkn2NFKDjxuAg0+yR7U1fDmK+Q5V7xhFIdKPYoKedcl
R3dQwsV3f3Nzoc1yF7SaQBBSx1gkLunllFckI4sMRoj8moaL8Ndr8nCybm9efrFw
CbZVErYAZCD/xLYDhpohKfrg3xDlFbKBINJdyprqHgsbWz5bGZiZsQQQiB5E/Uyn
srMhSxU0PpKIpQdMpGzseA==
`protect END_PROTECTED