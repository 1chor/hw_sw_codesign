-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
pMc/EaDjCQ6Y6jt978FL9m53Iy+758VJ6PJLR1tHBlChIK/6adoj3HxffTH8OEfW
yjhiCcSLgPaiV7PJVzbUtP8sepe1AxYywVE4MDW+lBVFPbgcIM1w/oebv+m6AM5e
+cMa3tjqfuTnxFWAimuTmgIPamgXZHksk8BD8mgRmCMwlcdvfT1/yQ==
--pragma protect end_key_block
--pragma protect digest_block
xdX0I3fpONnb7wsRo9NqXbzkqBI=
--pragma protect end_digest_block
--pragma protect data_block
Pd9H9FXxVduGSUOrrCT66DIg/1K5H4gePNIsdbzdelznSUU3bNpffytbMmEbFoep
2AvsTwXOLQ4vZpWKPKljCIy+1UY7L5stLrh3rZud0BBx9KV7kMWK4KZeDytchnEB
BYmQ8eRYunq2Vj+eIYXq/XCHC8Jgt6aSNNMMVLVjigURoSvL7Yda7NDmVDlJ1sZe
p8nC5vgGzDrKbIJRDzbW0bmfQwzcc3telUFiT3m7Hu5oBtDeJcyLu30kiiBZ0lIY
GwsVCzLC7Qw46m40IlvsIDk3ksBw268aWxunJL1DLdCseYx2LL0Y6s2tYTJvrbDD
MkSAL/MqvphMuCc69K7QI3sF9a0ZzarnmMMCeHyLsxsn9GxjVIjTpnj8o1NYFphG
PchrY93AO3t09mdmXtc7XronEBhyYf2MBepSyu/K+op2oMuJ7njx5RUws+XoGL20
pFEooOe0sKY0/kUiC0q8fJWHVYzxfAnjO0VaTuYiJdGW3o6SqFL5thyfcp35I66p
oTXk1sDs7gxATOk0WF2TbGADyHTUwZOAjMqfN6Wf4jIhnHI8sy3kDmNmfcX+n7Cb
kXvgUNnc1xdLLuk2n+q2vaFPbz4hpcyI7qiVoUdaWqnr9xkoSol59ijJXx2NJ8Yb
fe+uVAn/8n1qShQTGsvRvTOlHrAnx1KObHg0BhNT3wEzjkMwn8F7Wmlq7MxTPA/y
vhi4NMRxdvavfY1w9At8kwoOW4AOUqCfAh6JSHC0hXP6oLhNv3GgvU0wc1Xn4GYr
tpP02dsCWAMP4PNVsk/8Xxqu/n5oQcZw4sN3TdVjbyRv9eOCCvCj9tBXfMTz7L8J
wn17dhBtv0ejx/eH46UKku4bqwfgiTSScmGnl/pmzU8m18O4MKzniUY2ZA4qg1xJ
GVrDkHPNx8a+1DYoNmN68Ul1tlQXOXJw5T1TW7n5bSWDYp7KK+ZbI+niTiA3xQqx
cCxW+B/QalUr1UF+I0INyM+dwWHz3H+CdtH/46PokLKOWvlWlq4u+CGULky5LLi2
8ytp6L7vezYFoZgxAHEECjmKaJ029xwmkNHr+/xzagvZREushxosdXqrd7NHdNx6
t5lAviBy9E2uALpXFNzEAhBNlZU9xk+O9Wh3flAE9ykH3pQpE1sEfXLtUYRo1eFE
2MvStaagzyhl2u2+Qnm76e81XC7Sansa1s8oAuXkbxTePT+rp3Z9GWo0TkKbuT5G
+agzQuv2lkG5GY5cjwUUsF60HKnXYxsAsP1shpJNeeLMSIFBY4XuLNtHUsFbzpCp
7Gn+7yHkgblk0SUsfVGETPvMcP3E1IH2BzpJsMxpoLuIUhbSDx6m6dz35ajXRxbg
2BD1jfBKgokwhvksy9Po13sCeQ742IAyJeKnjsInkNUHZZrHOfgIz0luoXM2xzC6
khTiGRWquaCKF2LEilWujHE2Lx67nKY/LOGn5UEgOF+zmz9KmjUYmbzAcmDofYi2
1/xoomDXGMta8loiQYDfb9EGIxey64NEhq2bhIA5OYk7XKjTfhEVzyhziQ4zoeWA
zpsfHPBmuQ2ksG/HPgLBMh590rCHBqWXehZqoWE+GLiotKO5ZBxST6wTwOYKtWM7
2NTc5n2/HwdWNwi+SGquD+XXlUrjZ1PUAh+JEi42bsRCGlJBcZKS9WuPAcwKLUGc
QT3t0VcF3cabBpt8aTNZuunrFK5xYjJQ/pp/QDA1G+vhKgc8aFj6DKN4c6QwkQx/
nRf2JjoRClUKdV8YubqhE+WnK80oeKYONkDTEvoJsi4cw1lyDQOTy1cWvRAcoQHG
BEsgTo3HogxFjAYI9O1Q1V/yGuVU4KeCI+pWe4/F26XSvG09CXRKWwqWYmcqEtgw
jwHwneiw6Pz3b0KixXMZKdX/RUR8oTlKEqzF/oIEuir3xAKsk1krAyphgekYdNcv
zzP3focGnu8mGZYlksS3SWdRFXw59iLV3ZsbHMByRODquHsghMUIaOpDWPnkEfXq
eLgifAnQ+wLFgey/u8xlp4vVz0EpyoJSyIYYuBSsSbxteKh9RDx2nobOry7y6zgE
z6xM1ceqaZlEQmxD/eFF0p28IExqyMvVEBKwASdhN0OYtCXwmKJo+iWj1ca2WCRX
cvmTK0Ete5yJ6ve9Dhi8Q99CywqulM/Vo1d83eiCrciZ9lgr+P6H0IXCiHw6tHTB
38trJQH4fpY2SxOIDbSmj5uHOiLCoyB+/sDzkzk8oRwZFO6Y/CTX+E2FUjIy6urf
gusJVzBkCh14xouZ8v/M4+0caDljp57fg2zyqqhl98AwsZfQzRyd8G0cTW42x9Uv
EHHK6rK9m8z6bC/OW/yIRT4KZBtrlrJCZqP7zaGSk4yxHNTgTsqRAn4LhBfof2md
ZSe+bEOdzBicGVw7PpzEKiZ3CCpRAzxuMjCJQHO8f3qsJTz2obQwsEYjZx8vJ3D2
z7C9ktQbzRE8GDiBz7Og/rzqd/stUjET1HWAryhXoi/wRmkUzivOCg0BJszuYpzo
isdYysoHbh71Naln0ax9+9V7czpv4eU0TFUrsnlxIIN5M/wJutO4GrlmgGibRWhY
mNQhSZCk6Bh5wpqVx3TU4wgkm20QLrdXRjuOOiFwuhDQ886lHHdGnT4ecSUKBZAn
u2vlICaC6/IaRAcwsC4MoF4STVpqhCGSdJ6AUrZI28+EOAMRPAtOPiUvGZ5G0KWd
sSDwHQP9n6tZYtUg4disKQz4dcGANc/hUl/2nUmioLKYu+8gQvCbFGkDDxjM5ki5
zkDL0wPIjAj1xtBOhxoA+qOJnIqS/9LVTRyu8XsDf5xXz1DKEqXZH9dW6w8cOKIX
7pxosoZDcWm+c71cisOGKAAhPA3uymHXfzBnc2OiNHqBjiaR2apnHn+vup0LkWRk
7ec31eg3Dd7Ft7LOqZXL1g6+GHGDRftLHwiRx2uLE5IiWetQ8ldWdXMyYkqhHXtG
Jskj6nHQWboqxPK9RoCRNlDC4+xl86rqyOGifQHhr3pQfoSncipmZrk3piug/XFB
Vt9DGDcAQKUE0vjGbaPpY7OyQHOhVHontz9jSKNR7eL4j9ZMYDvvI4tV0iiwpIS3
XK9FFAA0Y1Clsz4tKc3zz8hnghkC1HzeVNYNABieR1563SUsroQe1QUEaCcXDcpS
/8W09O30Ps2hY2BODyAnczQd1HHkXRgHHNgCHJI3muzKT3WHJn1G/Esdo81L3HeO
uDftDCEjjd5z8rftJV/7yd61bTVbwF/TTDX1dk/3Vy5T9obj160OQGzDknICo4H2
JFxQDJo/Z8BkjcQj+kjVb5UfjDHo2+ZRytBEgYqPr836rNt5w6m6k5vyJhIf3jZF
DdnshoI5aB0iKKsIqg20hggkZnVVfwvUuWd5ajOY0h996pJSH584yQBf35A9vjkN
xvrPnCpKAYgXqDjN95cAHunnalBZeTNTv7etMe9t0rpjfTiX5r839O2rG2CpIxVR
MlRSty7d1KVu6vHqQjJ3cnF61O1AlERqXyV+6SuTshm/DPYmHqJJ/4DkTM8jXe/Q
Qyr54zag7YF8eyKaFGVbFml45KzNq7sxFHJMFzhh1W+9C/fRmM8Kta2LiN9cmdnc
QbV62QKkct5oA6nK/WETx1ZHxehIyD0j/kYneAunsteID3Fkm39n1LOCBwr84lMv
AWq0c2TxQSOl3tRRYpZ8eReEqko/sFIdHVuzC9nUrB+99SnCvs3aqqynLdlV/22Z
1FIynbR3YaBU2TFrMVZJGm40B8/k/CAEMaT6TcoFmBo6AqpA2EuQmIE3VY2FyLk6
D+cZoPO7ULYJ1B6iG+CQEjD4U8k4sFZUgkDo24ebT2qmBOrEkVJWTPnXSNG102gW
2FEuYP/7EGvfUSELTL0P2Mxtb26NbPc4JQ4dTvXwggm97nUosIWWeVofuV0vo7V7
gNtZsKeQU3Hw/d8L4mEBOVKouG06LvhIkmRaHeEIzoocDIDKWiSofPOHsTFSBkvk
R4eVKgS3n0/TwEKhTYj8FxuLdz7Vjrccrn32gxWAXgbUO12C1RUvOLyOUUBBEu9c
f5jX9V1DslYIQOQWqNg5saCwWpKpgJCTGu0X8Mnwq+e+5BHpvN/QabvBbgqEXMvo
6KDBxrjlIvmEsesg1Q0H/QhYEdCTZYZLGj49uu6FISh1bIYbabi47gmLLOSGFhP5
4lARjf3ZprgXmaapzqsJVbmVVAU+qtxWw2Ahb6Wgdi4GhVdsJt1eNfbXVhRDdq+V
NgjTFlwLbBwEbQhfmzq6iz0dcYCiYSQjsvCx8WbMjdwbfiXX5dTwE2QTXYriRRzC
8rybSP7PFAfNswlcQRmCPL1PS5G/J4PIxitTl1ea4T0N8oOpJbR5eausJEjltSAh
fXYhvW1sv98/S0Z0dNr8woq08/KkqLyhvZCMImsySCzY8eITs+U+mGrkYsovU/fl
fC587/n/HDfh7OwtSJ7xBgRHRlGSbY/rCiYJ53YiaQdYzXWedBkdPEkLFU3nHjbp
CpcLPOJP1FUg4nb2+FAn6qH8FaPqnhYmxojuWHWWaeJZN9frzamXaRpSOiwVNGZ8
2PDJ1Zamqx9KuqtM3LcghVkBgSt5RkbMdMDU9YOsqyfxY3uqQcGf5HWj6EMmnaXS
USHPknNtGUZYMxn+lIYgATRAT8Ffv81XFuEby9E7ekU+ZVItpmpjkKPUJNUhPE+u
G925W9tzG4cWjd4u1qRvXAyC9ITE9wjpqzBJ1vb79cfVApwpiT4w+Y/u2Jhf76KS
MLtMZTPYXaCx3Fjvm4WS7tzC5+8Y8e906sgq8WIKCXQUiYXRIdICRFYotPz0aHYl
yErZDfxYja6nQW7b51APqCc9FL+0l73enlbKplz5dCtp7GWtOjk607C57cvXCl9d
8zFoRBEpSsRsKqoCPfle16821lCdXEgnpixrRpfidgJ1p6KHhzC/bQuC/8A6gqeT
LQgGBZwejkCNo2wBWPl8Tz21miqe+Z8w/Wo8P+w83+JvchpSnjAqe9X/386ibnqv
Hs6G/XjKRUkofPAC3+CNehedbeF9ThvbP5o7+FZFmGTVobxWGDQFInjlG8e0Mzbb
Hmjebfi4FJ1LFzZ2isYVIbNEEMK+R/5pfpa4zniHgpqvGyV3yJ6PIRbabcE8+2hk
svbIGOI6miSUS2GSawF5enMmbH1OPhPHLcbr0vJjaUSEba+66Q8Xq3eapaMGI/Im
/iZSGHXHu4CHgvSPWu7MVgKuGyLO06HFav7Xirfoa+EmhB57TZiNds0WymMIfS/P
6dOpO7SQ3E6bnmFY6+E/C8K9KSHHSCD5x/YCxsszCodft+RvqbIuxSc9+ubbT55V
/2Hucm1ohTULNXtgLFbc1GX5Zuxm4uCg6uWnVGfPWY9JqDArliuDX0boBbe1EWpX
x3Grgv09siujL1Zs5rIzsb7likDM6j+2AUl47bTEfr5ii8js8SlQvni+AZlkZZjp
htKbECoimYxGu02jLgt8JMtuqi8h+6d2xb/STl69PM6FtukhGeUHqDG/cFvA6sWB
yeU+tCahOhrkOS9vltrBHpx0U9tJUI3nXcQ4QB/KIPzy8eBhh9cBXOnjBD6aX1Hc
OUFPvS5uu7z5wd8ab5OJb9ANcErDCTcVsKcnxEWtJ4vQDoaXoKkRABQ4oiSy+iyF
STMigZUg8EIdJkIcwK8PlX5NWMx+nb63uyvJiRPKXQF8oSTC0iqNAxEkSF/A9s5R
XfPfOzjTRitbdtOdtEVU0JRKlckggAEARAxL5vm8891P8sPtHXZHLMzxZx8LINAG
yExA4t5h5OpnmfMj804ZXo6718dox+TFOcH54ZurJQ6LdEo2pyDh7sG/4rTisRFS
Whr3tfYmRi0Fo8XUlCaq5cz/U7I5+0JimsRYZvBgs1gGuSt191n7k6+clmmNkvpM
AHYLKvrqSBsBmNqPvvb8XH2+2OUYouuuT93iMLCiAYMg19DIlRgt2bDJy5Z5hp4V
TmirefNE+VK2YjME1bSgnU6UEfVJfZfGxWiI3c7lg/f4jrIClD1omdFKaLxnZLz3
XPx3iArHIefI/u7MuKFZjhMbNkV4h/ColwS+tg0jXgeNATLPahkcg/NTXsYdRP3e
UB3PqlaZdPY26IM7YcsT/0qoGgTqjArpRgCpl9mefrLVMo2yVGWOCvhkrIcTajus
O+7XiDVDNQ/Pd0ogA9qP2PDeMY74zf1wlnqAHj0GCTeQ/H7ieVMHiuelHKY77+xC
8U4h+cToLIzkqvOcVtoq34opdZmzpMZqA7fglZEbJW8n20Wxim2U6mI92XKo9NrP
PsK9ZulwvvcG462Ny82Ovty46/p9nNgR9oi5dVodRuKGvGZ0yCKXwJW2dFRBcwM5
9mjWdvbg/8aJVzCaMzhxyH9rFF/Pgierx3hMp5mWYRSErpbyTpl6Gbl9qsBqVVpz
UX+yToZR1qXZLUeKiKsd/NoGBMOTStno7soE55rTc5GDYjQf/XmE09TUCRTOp684
lrrSOoreNceUKLDAGmgtAdewe711cqWM2JLS7ZMil+VtLhEjG1zBHKg5i3TGfEPT
GW+BeIsVTza7H1FjeqFcYJ6ILZ7KbdzJy08HEEEBeBUUZR7K8zYZkuTop1rzAh0i
xnM95EKnfkxTLOfAg5vG/twDUzXJ7gGRgcm1QMSaQYss1sPbo+d3TqZa2CkJ24WF
IdRk4B0Xsm/ViwbAxcc1dFuOXoDwN4rXgrSMAuyNkfXpvQnPX/g/p8l2N6DCvWa9
yDcaBmeYZO8yVk5t+IcZNtOJe+fS9xIzFij5FtB7L345uhoBQ1kqVacxCyEvwr4r
RbtDrph7cfarV/bw2cVkcop64o1bDX61OtpFi7OoAJcpMoOpaM9XPV/YyvS0KjnO
V0i+HbvCFHzLnpxF9z5twvonrV1l0cRFIQWXqe90gMOBLX54dYb/09Y65qdz/U7b
1nw2WWsy6TkNBS8Wr1SpVTJpSjUgN2j3OljKlzQjLRz4H5OrDy9cLeF+l60VCSDE
WYz4OLUy5Fs4rkXkb1VqOzk0YRt8Z2+a/sFDfHn5e73HxZJco4QRC5ZtpGsDt+tD
q4oTxf1jUGXx+T8HyEJxSIlMVHHNhfspvLbZv6GPAv68IMralOi7rS4s2RgGy9eT
r7Uzn+xTYpzUz0vrSH85QvnRbz6QgXv0Cz96d21mPpnAi8bSRccAouvD2hpT9lPR
UtYj2/GhYF09BQJumiW3IKbFjMDTjQQ8kt8v/HesF/7EWEATnUuVxJDh8/r4IN4n
kVLvIPfP3ku2OH9zvaBr34Xgbh3ZPVAf7AmYKYdi6jruomTOpbIR1NdFjNMIQqUQ
WWbPxEX29I+IEHefSwWSWIYaMZcvIU5h0jlbjQIVy8ggt7tcUTVUzxrf5CPZGWrt
s8CH1ZOtL7gWFHW1uxI1WIf0I0WUdal98Z1j8EMM7YmBq7e9GitHi/aYnoNiSNJS
t/JgE6w/dQUn+9nSt7og3ZsxMP2nrIzipO2jn6YFdyFRSAeBKbC5tMyvUvB/PD4i
iPPWN3TIdIkdTXlNZhSanAKofT8N4WRCP5mnQrLg3CPGZDPfa7PZ86vZ43HQaeoZ
FeyqCQNqZq4MnSgjcntWY3vktfPs+3N8Fb7Ya+UBXB0aa8YmchMv2bh37ptSTkHa
4NJciIo4R1z3Y9uat6qfmv7mXS5/ckJNyVMVqSP+JaaMqhH2gZY1pGCybVpd9xIl
7IkAMOP50dtE7WvuicUN0un9TEglYPwDMDVoffy4m3alLIHNmXXrs02KPoFOVFAx
ZOgtwc3vJmmX8Z2FmYShisQ91E04PD7Y7/lnNT9RbfSd4oWtmiFdbmKpRjHcUlOi
Lt9J+eBve7hDMIUJCBUfvnvIKkmHOuLS/ApYKXZx4VHCG5V/ZZW8t1om9TRIIG2b
K5Rz8FnwoeOHsFK80vDCjONw2rL3Ib+n5dj8v4UbYgk7u2DlI/oQ5Agw92BV04A+
AMvkrzjYLi9h6WnnfVF4YGcatWC4QEjgKoAVpLMS3yROX7eSGFQi3X2insaBz/yd
iIEin6MH7LfXIGHHBzhYBMbvyVZ5VjAoPuq2Vm4vRs1FiwXJSiQPAxt1O9rFbJE5
dzEiTHN28irRurAqLIJ49+W4NddvHkk4NvsOv6yogRYKWp25Qgj63oL30Hzelzz2
KPEMf5gqOSGNNJyLf8Cbn5wk6rg/NR/LY1snXXfLy+wWli6b+YYqkH3nSjTNWqM9
E7qVkubck5/U3CU2UdagucWjfeoeiF5aS9DzCTM6qjSzT4UHi1YEXnyLHax+TPIr
UEDgTm6Mfk20/FiHvGTQ9nE2/RE2w9ZMuyeiHJYo+E8d7h6o7brOMIUB/SFOC5ku
NeFTqsrOBOLyKaRxsqvoZml7QjwzXdcD6mXTA/J7H6x06S34J7F4W5hywbnYxNyq
fo8aLqS5OVg89DS43NaXsQSPDGcCbwCnP02d7SfoYEKzqa84iuNyPVlnOY5iylI/
yaCScRDT0X9LKCr6UJ602syUM11mj0fbQBpJWLmrkoDcMNbSUUVazlOzd2V3fm6S
F0Kg0KtRO4SbDN3YqHs0jedpTaYWQ5U+w2O68sGLSQlUQiA3etBlAc6o+yHGkbqE
B/IYTqAe+5WMnZS52KLBQNudkC0e5tMaUS7/0R0RjFjXpC6FCuvsPu2Eci1SnEfh
wOWVW7ZR5PQ6aQbkubPRcRoFTU7FW38CyyAlTLnCNMgDmTwP8ztxiy4vWc4ROCWF
vtGjNR3Uafbft/7q9pucM0tn3wrU0pWlFXrj2ynyZexJDzwxBXpiYcmLUfJd9CaH
jRrGum61Y77hv5NSlRd5pKOrTpQ+0zXieBeL/t1AEVAJA+U7gogt6cypk0XUUT2E
2vLVZICjQ3Qh/EJFXj1s8Yf6/Moz1O49gE12x8ueblYoyfYy2+Hax+fSM1n78P+u
cKzMWPzYxKPmJwvwJzF27NpNZcTj3JOzzneqD7b+q5S/ceg4Yd0YMhHglMhQzNJ1
69vlVUIhB5NEjyAusGTKQ5qumywXwXtDaZ56H+bWyY9xH8IxM+1doPC6Wo+K7IKw
sucOnz8hiBii+91tQ+QIvuEEgXMrpCkbBK3ayow6HtWd2upLOPRM382W27YuUBrD
xfW89gWDh2IQ0894hy1adlGN+yF19lHclbDSbTXBEM1TXFZK+ZT0xNnT6lCIbmD1
6ML31Ai/v1HeCXddpRx6dy27czzQktg0wkHrBVZNDtKjS1SSglA25SZYocVREuIQ
QWYS5Nj5sBLCes6DAP94YbBRVwYCE499ZQGNKfabknRoxKdOWHvqEY4SR6ZCyM8M
P/eLEt7PxD7Ip5Lo6+qjnUIWfs2Ev4OPoyiZOuhDyDhtWAnO4txle73dQzAqAV/h
VYDTepWswn4qvIYgBMaEPaktnNIyYLLr1cDFGvMhaysdYm0pWErKMn6K0L7HkWXB
aY1ChIwgYsWFFCUyRw3rTrQXz5q+CYV1N+kMVzAPkIzUkP+xAIlWA3HE72/DHbm8
1y8LZKOBnoxvYD0/7vIWYcIPgoUFXSSGTKptGVXbhWXsjEvHFsxsanMMuoppxXKf
DkkVdzu5p4koBiEoXxtCbCTF+5OgqB64JCiJZ4MFp9oR8AD7pPftbYB6pqoHtIPP
YPNgmuK9gnbYhK49/UXotGRM5V2iHDBR1QKvl5wOLeM+mguyi46Gd/R4/IY3lXQZ
LRmpxhuocULIBr2ZKFCAPZdThJPWip3qoMZO0/SdHvFTyReyBrmGzKFBCy8SwWjV
fsZFAz2Xw/fQzKLfAOh/DmMgQuC7RM40oXqYXzSx93PhDTDZ1DGHeo1Nl/2ozUyR
yyzooCu/lCa7cYXxyN5aMvRQ1ajfGPGEN4DH9bpwWToHDnnGwbl7tFb4c2SCtu4b
s/JeEZy1iPGHKKmWGBuKK/779i9Y98lxCn76xEYEcilnxXa5bxoORxt7lD3+vbQm
naFlWTt1AIVPvt5hzO8od+z9FMKrTzZHw6y3z3gfuI4nKzPQCcMP16fL5bYx+0ES
MuKWRv5xQdCA6LFI0bfy1lirEpMUeXWcx39F0l+U5hvNP/rQBUxjZUz5f/kmqLhb
Q9k5DGS5uqCTP5YNjQ7uYhpMCBaUm6rtBv7nnfn+R6YDfCO8t50UW3LSeu1uzYtF
rYKNGRW00vpon3TQlpRLGo2g0YyTpZZVYvhOfHw+OR4BgfKaPbCC9Wb6mnNBJBqR
+nvBquHgfhQNj5M1OeIkd9Tlny73aRa5fzRVsNWTqFUDbQaJA9h1p4rdycGtxh+Z
fgIBhykIe2wQHc/W601Lrrlw5J8+s20gscOt+6Pr4YTPReENGDy/4AfiHhkP7do+
6WXUIS6mFNHp9jDOpFWC9pqmAb+EmkfP06XcavzMECP8mHjjLTIraAMuyqO3yBaU
WJ56t8YVQ5LmuMdUHv1AYQTfMeCgA/+xNURPxkVZDiXie4ax5fHCxbfmqWWC6nOg
UM5HQafDN6RcmuZdDpRqb/sWv603oygprs2cu6sf3QvhnN/7t/VhRQokSPx7+JVG
WhjppmbcQgLKDnx7K4O8XTXlmvxXwd1BKlLC/QuTUfq+hQqtspWw1MhZkWN8n39V
2VCLwHbWBTVt3gQQQB4VTSQ1ppwipXOP45yKoQ0OWT/dP6YXU9Wuf0SU7OUF0svW
t8tbM1HDACLCSDMr3vxHScXgVcldhyN6+J1NxgszybnxaTqx4gm1hJwZ3hOTrtiO
USR7Mwr78iUwen6hnYxoy6JbdGeRraZgc2ILgbhQAC/gNku5thgiC88OLp6HUo9h
7O7Mz+ssjnEckRl0BiHVDPsgHOIeD8uzbvoOCMRq3/OdgO9UMtt0TAyP0Lzzz+O3
Fko6bPZc6JL2qFjVaztN5EwpIhS1zymXNPbMgkZZdlmGjZLp0sJaTDOVyJVaYTgS
6NduPWpa25umblrDaceI4p8kbadAy7K2Enh4wMdGyaZo8QErfX8caItZVC6+fxLA
A1XKwjxxQeQ1uS13nOiDc8qViUaR5XZEaBV7q/7PiF3UOE1xTs1A+zEUc8iRR/nV
WYr40e6+r1MS2AzU/hgmffvOeWXtexVXfdpE4EWd0WUwZ15jQNjnKTM5oj30Jj4t
7YXWCEuMaNfXRFJ61Bp9iWNQXfcE5kVZohh0038c6NbfTuVpj8kon6ZyaZCrPqWh
0HH9ZL97B7FeKFnoHFsw6B5tUtqW2IKnrzAmJYTgqDgdImpjY4lR5D1zR5elcnAl
+bYzrA4mIchvAk9ixVm+ewfHSJj6OAbncSNKk5anGeCWTC0j2T6iFJGE7EemSWt0
+sNAHGebWhDZoRDLBI6eAovgklnZ4KohcRPdhN/L+NnRX4N0xBrIcThEobImZY7y
Pwj4krXL6KLQJTmIH3G6F5AgeQPAGViAyRIgT/atA1wUPsBMd+9w2CGyUB99epD5
bBToGdxZvwWt8ufxYBQnpCx0NAMnFziQXyScDa0yUeiTvbtVm0wJ2bPzhmYeA5gj
aOoDB58gmn0sDIIriDHzd65O7ZOvQeeFrdkT9prKbg1KUblvTipLxXKCIIbVs/yp
49HD9DrBopko2QmQdOC4P0l3BTobBZOf9qs1FB+Im+K2ClF30HmSOHxHrzTqlFpa
GkmjXJcUQScpNOcN8EeobnCRCVnDXsRhvRSKJ2qHT6sySuYJlDwDm5Kibwsat3b7
66MKgK2538uh0BT381HpuDJpo7Tyq0vvCSIkgmvHeNOKWz9paDZ790OJgyJbbJFE
pRHjcybWQIlbE0CF9cbxiy7vnObR75ExnrQzE1uoHPyNI/HjWyKs+XZ5uB4gVDV7
DdV5f+6j0Kz5cNWiUv+/ZQMPSqEW6fu/LsswoVwhCqCG/ivoVUzvaO6V7biBfuZV
aj2Fkbvp2wcAepT07+XSSqHNoXjvkyLn9gJik5A8Is3JRhQca/Yl+i71nls4dsZP
FCBLTX52+UVMbv0O6ei+6S3O4PNDViAOY01Am9Og64jTtOzISzQGB3VlgQaqTBg4
Rb0fDhuAHfPOknvNk9l7UzLqUKFYZka6cGuJ05Yb9f6TTeLtgnR5e7l+WEk9GQsk
B2HtFmG/yjgdQqEhu4TnfZwgeS2oSSRUCTP5RIXRYRuxXIKZRv1ktIc9DtKPT62C
70ecDQobiCgXRX6AP+LALM01oGeA7ZjX3sZK7SKYp7ycVYrS5r9JNwhPxOPIcUKO
AYJS2fbvhrOMlhHvXtQ5Pdy9NGnVg5eXlUiazEFAfp21PrKD4AbwFJRHMEBkUudR
0tVKRybrif7iwZmTsWFKMnoN1dUvKa2Y2scOZwMj5P29F5utxeYzrQ13GwjNo5SL
4Y8/jO5CO5AuBbwtG02OPQ/LZZT4DxMy/6Leezx/ZmYDpQjIfDE8Qk0Vb/kXfQl+
q8kvPObJqzi9mW1pApfY6WdoznNswpl6BeQ5dWgxhilnN/WwfQmTQGKT6zutt1yE
pELwTbmVpAFD7EVucJfw+E5yKx+2Xj+YhORTbjNlPu0KO+J+BolNZMmzWH4O05o4
MAYm6gCy2yiNBatPhRQ0I9kgA02UJEzVqK49i9XSNGMK7J0XkurwRfylVnsnzr1y
GPUdSCUfqewlS1RkBrmitaraQlMJVMSYBp/fMcOalp5s3i6lBXb9/DMHlH/9ySak
Jk3yqjzb5o2qlO4tAvp3orM7yZfIDcRjAUN+/gQ4dwa2x+7OgabMY23pWugCbIhM
Qu4oRREYuQtOMrr2DfpOAEM+K2vowZWBtCdDjhNaaOBdABbwKABSZbtizACU/+ah
VbIL8uC3d5NyJ4FR9UkcX4MOBcPKlJt0VO9S30Kfzmh1INwPVRwDLs7uLq0m6Bhb
5ti7HDf/BYint0ynwlBJFgjGUXYKBT5f+F0TsOn1gFnE1S1VZyGmqHbLDVVVcYH4
0LY2mlZq9KQpZ6b/ApL22GORm8lX7ZdgYuRLzDJNvKuGChcUBoDKUSbjQfNb1zsh
f0UHPGxQv7h/v9QjR9MdbJGmz64TCNMCrKsEMtH2wgKWMnq8kD0uy+iTThSWWcDv
rsTFcW3Ln+cm+jZnq2SxCI0M4efi4o4KphRV3ZXUteHyA0wy23v5KBxi+sCkUw8s
PLKRaA9lzRkyyTt2oXyw9rdwVnvy8vosLelRNJ8nofSaVoEqmziZLFjB2cCfFxks
AEiDRBkQnHpc6UY4xKJGnt6mDz51PHkIURt8BFgIiCcTGcz5N2lGAoQWWKJTmSkJ
340cCoVCXUwGxSKSMOTcgH4NBEZjfCsbmZibA3fHY05eCtsWQFP5XmnxJSdYqHuM
byKeBP83yYY263n0bhmxrfFbMuoXOoObDhkv7uwj5r+jHUIvKxdoeGgbx1M9wu4L
c/2LlgTOmpgoExl8nyJRsnUaeIXmtJHCFnZSpeHgAGOxGReN5jwEstbVf3jP03LI
v+oZf4FMZVOaQ7lwum5fftxYRTtF81wtWX3hXupp12IFGBi+zCjbv5tLkNWktuQU
yojTV/2854pI6fkYGhBXDV50Jr8IjSBcOcUiPP/X/YU8LvsIzrxL35CjeVrGUqnx
Du4XtcApHT37FwDiURLRAnIUrC8UgZRlcZlg7Vs2M8a6ogVNCeJrzQmFnz5akGLi
inhxAP2y1q2OywAH5S2Q+i59F9obq8iR0wIHqhhX2Zb6AGGjQvUm8R/npRLc7H1Y
EbVVfgU8T2flfg/Mys4/8rZM4cgiQUlRY06+xrac36Tk9RcTYBeDb3jpQI/4BXOk
FneXS4h2KxQLIMxQcfnd7GBv49oXqqSq/q41C73nYkSNi4NTuHRWxtVlqasOdP2Q
cbRPagCSspK4YecVYVYDFmb5Kqi5wR22Noe9P0NrcbPSvvpapWs+MvM+Ih7IFu2a
P+28V2tuCxMzNS3p50vFxnFnLxlytde5BTqV1vhHKoucL7x25cZ9kGNMjaUzIh/F
SCbTZkjtB2oE617RDOSayZFNhMm5iJZqduwop9cXnMI9cDEiAcBNE/TuyTQ8N5nW
GQ1mx63E0R5CtPgsZjO+Le+Tfm9fjD/Y2cJ6aUeup19mgrIF2AL2sGccIiWN5b9g
aTDzWguT0eYLGRz77DvaXHbH9ro3HsIiWnVcWtO2YHRPy8KT2dy3nzuLbvD9bj0R
sMMfi+KschpdOcnslnad7cTkjnjYVuh7SXRsSNjK2jq0LVVA/jM+pezw/dKVx3jL
Sjbbtf4EFGSOM2ooDtYoOfGSEpfsdRALUPC8rAtl4pzKSW/mlRTOZIZmG6gWIW3W
djHq+rWgHm9CI3ZM/wmvbj1sbGS+Ha5ZT3xK8BBHFG7aqENzDbOvoAnUXZ7Cqvs3
Z3kc6He14zhN6BeoM0lDzPKZAjlZx52B3qelZv4DLducA1+Z3lP6Y/9pP4cTUIeX
8vCmDIrPQBWCvkatzyZM/FUUZi9DuE/A4wAJ5y/wkKCCqbWj5+6vDBPMSI/Zx6j0
XbnnshimKG2kuqWYlW7IqxqLXdG/PkFdyGKGiHuAt67OflB4UaUD3mkHe/UQ1vSC
Cugu3P8S6BSSIk/A+XOnZiZdRJDhK8kcW2jnPvChWAXZXFSVsKHPQBhifDkCFbTf
swcQbTC2yOo0gL2IGSGdDmNgle+8KwIGZiOolvVknZoPsPA1TeMzTonJKjxqNLcN
3jpXiNr4UebbK12USSJEa7G7AxwdrQ747LLxGPClkKwRAMtEzzdQ2dic5Q1wmcDR
K6SkOipk+YRfHRqKWItNwVXJmL+C/5lYHNtE2qal7vIuxMP0wR2kdMZRYssowKzA
50Zlqa2Um/pyy53lBKZw7hRNbO0jAU4tcoO9CYvMZGFnQnbniEkimZS3dM3Ni62Q
3NocINzyzRxNj7egzAqm9FnhknrAtW1jRw0SR5YC1cXRvG+rLW6oegDkX2VEg2KK
Mj7GX9VyS1R5dfHIVZcmb89pHuvG5EwmctDPQAYLTZRlw6Fn6Fyo4/NZ1z//4Y/F
i/54BAXjZ+HbCy4AcsWvnQiV4ef/dot5wppY7Ypm5peWlrTAi7q9a8B8e5oCJAlJ
FI8VrS+MAXrI3uMxE7u0eh9lHEmX3TW6/Ra00PDp6s/5Wb7YGOH9Q7645KFjkiCm
Decju5Vo8ZEmrLBVHEdEW8NGqnNq9GVyMoJM00KZosAx1JLiyhsctSwFzn4kpudM
rTeUk+Oj7qsQ+NuvjfzTWLea/4ZytXUC+V2L3tLab6iF3hxScGcZLkxCEFHD+Fj7
R+oQZ/fApPoOOYbBFIF/zseLRW/I2SIdrwINdtlSN7SUxkx1YbtmjXcW+fuSXCPA
Sx304GHAh2lNYP6MX50xYtgc+aDF5oMWY6XWc3YlNLi1EeH91LVDIXo1mvQf5QKo
BttQJgjIxmTnH25IbfHWTvUEr/QRi7Cjd2AqxTchlNoSAj3FjG844ScF8Gq9ZDwG
JV6ZeJwK+dymvEPEBBK5Wruc8X03cpaS/t9B2D/DZWau4/Ay0Wc7YaR2D/Pvns8r
53JSUWhGMCaAXCCtBBu7pbmuWt3FFtH2AFR19LznxMLZUxHQHmwT6k6KfsexF9Zl
2AL7Sl96FBI5oSG484HD+Hw2x/sQDyWj4eGwA9qSune6ljRPwU4dfAUmk1FZv6nq
rwR3JnYq78mcep/YQt76ni1w6e88xnUnVd5mTca7n6apMdFRMFksgXjBBWz9moFB
ktQAQiuL5z44JrT8ReZvY9hEjUCf+BRzSAWtTIVblZrbmmUgC2Q5YwcaQ18bb0/2
BBVyDu6iYorpqH52AGmHh3PGzNY8vBybyW+Dl2qyYMRTAC+beXPDGnpl38WcsLCO
w2mWaul4Q6KferbJkIegEynTscdXGUkvvKOGGvNndJqkP+WJ60Q1BsAelY0YAm+n
ci9I0IWj9DAwTBc1JzQvxlQo33ylOGoUOtSjHF4YMvCX6Sv4B1xIOgOzREuSMPTL
Vd++2f5cViDBC0ijsTQa3pDHY1vgLzGIkAQ1mW1XOnsUJsP6pzjIrKZibcUJJqOq
VO9ZJU8cWVOFIVjsQyxznYZbGI2v0fxoJQXSw3lPV1/xiFLmP9ajgFO35wi1j9iZ
7katopSBWYjSJSVO/A4HJt+1wo6viN0hF8T/E7idM++UtrQkekGs2kZ1BeXfbJxu
7k9990yP8/jVuhzyUawSXCtfB7M5/M/7g6uqDjSVRMAyMchgHjUoK+9PN6toKItw
N7ecyFzW06zV+luAzt+ZCydkQwaSQM/grBKZxuSOXhp7teJwgC0jyM48enIbvpG1
m3UHB5f3iSY6EcAjV9UolAdorJCwweUq25+NLXzRmYAejJwdJb0T77G7PciJt/y4
keNBC3kn7qzCy94X3C0dqKCVHECLennzjkLbnU2AdF98AVhMQs/gAfY0Ofq5m7JJ
qJQtagqKsOPQyXO6qR3/fph5eSfqs9RZq3ReRn8vefqeoQaDfyaYO3VIOwmZG4r3
oo5CvnR9U9wbYMcab9fc49DjNTee1fHcNMP7J3FAmVRVUUWdxg3ihsnZcqMiextF
OCupFA8mDjh0rHZjKs8rnRJXONGeHMDCckYXHktFyzHdI9lbyHNFbe6mR76/W66i
C4+8vyvQp+n9o6vRooc4fQQkXDOTJQz7/so2gqYPAQkOJ84orUa44FUhqSPOYTph
Zeb8I5FpwJROnKat/7tMGfzsIQ0Fm4NhwKd1i4tpbLJlxdPR9CO/CjBt2/btpZoG
yHebMDcqRHJ7BhaU3LXkZkbhNtVBP5ZUyezzUrAGBmhLmqElmUDVr/a1c+ejw5+u
0XbyBuxFy1WtzdxWeJs6HGh7yoHaWmJkm5YrnMdOu+U2EbK+Bd2U7bzGJXbMKeSh
QUaYAai3U+FTUxG/J7CZVuD2+V6B00vy6JHr/GDirPCEO28kHHztuAhre603pSZQ
WOPEATxiXFPG739Qe6Ya8U0PLTN+QPNtYHNdXbrGP5hfdpJ04nwhw7lB9F5AwJea
mKyT39WdQ4oeA+haJk+SacCJ4WZc9Cy3mmHPejk47+y6lewZ5VEt6t7lDjQGW/8J
241/DYfBn1suVz+zpWoQIQQI4OG1oL2h2HxmPc/3k7K9T0APa5yG2lbjamnoJy8n
XG9kG5O+6phj+CP0S7zlKW71UqHdfXAMXNDJ/lfUh+KtpLE10Woav22ww3jMcAN0
f6sUS6iicFCwTn1Vv3XMQFRAMybdj4cU4kr5y/O2f8d5ScjEFUkgVrjlWPpm7MjD
QEUTliEuxzjLRCK64qrfSa9OtUm2GGkT/40eQl2ma/yUUY5z2v6MAhVm23B7VprE
wpxWKLKx/K0DplnxP5SlFYmBnpUyeXGQ/NCz/GDEC+v+Zmtv+autTLeMsh2djqxO
RC6SzUXC03HgJQeEnx/1SrcrKAjUly7c/xJj5Jd4mnewDiTmYuezhA0+QnAXAm0l
Dv1SF0GNOrz1odYN7Syx+X8Hu6qZy9NAlmCF47XoR8URbiAaiZ1cbBkmUXBBzmOr
f4YUHC6FhUmJLUxOod7nBrt35IGVzFEpmUS0d7E4yBt7YaxkVJ/RiNW3lvsDY06z
D9Mf5Q9YsYTtDTMBuXh6iapTq0vbI4EoNvZmejG1kkD/glKN2mcGCiz4vVesTBU8
aUq5qh3IpTQAI8oD0X7pMogg/ckMyDsiK/bf/cjMX9leEFW3qt+F9tgyC7+YGSM8
Ka2oXR59H3YLW1vlgTbYLtX1GbNQFbPptpaPkruGoX25UXQTt9zESpL5kUc0L7pn
l/9JVbjgE4INnw3f1zUlac1iPYjuuRw3qksKz2TfTRxTp73LShne0oVb8Gek+JVR
tmp8PAMGR6fqZ57x3HqWRTEVTqAId3h8FNVMYVjNWzk5cN5zz/AqqVKCxA4yo2+R
fZsnup1SM5Mz0L9bzN98ZYrVa5ih9kNFw108+HNfeEHU15TmnV7wwl3LrBpjla71
lvs6yrhtWCyp6VImwM5+kTpg5NK13WjK3+o7XwfgtiYK78CLfYYg8mpt1bDk8hja
lggOvwaI/d2e0NXakoGL3JqMgujDGYm7XgxMToNoLOv+hNYJnCJNA/zz6yi0XCNZ
2C/GHauRL5FWfZRexw9xX/tQTkc6NwjGGgO0QuSF9TM4U0yVq7pWT/SCFjv1rI49
asl91YbfLJpCJZHGNP0U1yWIF6s7yZaiUnLuhp6lr5VsA4WOX2UMNpq8mMzpsmln
ICIBAZM8CWbebUBkmKtX6ZL7BgSxU43c9B5C2/Sa+HdQyj1GzhEsl31HDupeyWnf
0l+yejIhl/tl+lca0UcWA2Racnd3PY7YRSKZ+GYUjZTzR20kGfZOMECKBxGMd5aZ
/8x64/HZIXseBcB9hswtfHTEK8iyExKFjYGsPI0YHz4k+Dx2G2L6oSJoR0+fhrnO
IbXdbyj9S2SlrfW6FYACVj6eOhr8B/vlfZ+7FNmRg309OLp8swoSLGjAbD3k9rZ1
69DusI1hubXjShbKu4Ng4TxFWdxanGMkGQmEdm/0fxLoRyhDgQThNKcegYCLz+oK
khf432KYVhK3VOR96WCmn4LnmVgR2RU1QNimsgDeUjeyi/QRSgJnpwFgqwJV1nB7
ajjBA8aZPmHbz0Lv58LA3yfx2xujtuEcSdpItitaNS7gwRBRVtk0HXA83D8K1ptd
6HJylzIgXzTeCCcgIxDwj33dlNqYKNQjzsy3LnkM73USPlLXIdSWQw4Fma8loe5a
DP05NPsMStjHvqb4UwdMiQ7aAMpvCIvyNGn/gvvNfmS620RD+SdXPQ+5ylrDRf8V
JFkp7770OomVkMAIAwP+vFSRkaq3X9Ip061CML63zlZgVZIGplHlV6iBzULJ3K87
eTk1eJnkrohFs0CNowgn4kMYL4mjz0v0YLECA5veA6CWD7+mGilAbXwxGzhJKOMa
w8/B5Z7Kf0SERiLl41S2TYbrdxExtDqoW09zjfFjyO3slZIPo/GffRkjVLc69Kh2
2/XEATgxDffBWUIPIo7oCBUNIfckuZOOwQ6jAlaAmC/6sbuIf/+4XgyygOqs+bod
CsDBPF7Zg89cw+4dWVQktdNc0+B0bRhYy/bo36cNABSpflqpd9cBsMT/Zm5R737t
og1BaAHP9osXKFOBn795XbL9Au2pjE1uEKZ/5COuP0JqomrtY0EMM+CEfqpKi0Sx
l/89u7V0g75+YFSuDI6SyOPFFB/AEhN9ei9y83tmwS+M375YrzsQ5y15TL2nybL1
SZ0DzH58Auj0F4yGsSK9ij8YJmSNnWMmtv/To92Me9SVUM7rrXFjWppGfjzj9Kn9
CB/Bc4UhAwU9Uj9vqSQRg8BnA8PIcbAtNgSQFhA4GHY5/LyjdOzvsItajVPVm70i
DFnULCedTHvgCAzNmOEm+lBwy4XsrN0LBkw9JlokES1WUVeusgMdoWK9tMtOT44v
x2Y8t15wQnE2OQ39ww+mOs4ADcqEYX2tAOCvGbNC0eOI4uIY6p9u3tMvwSWqLwDn
91wFPA/fCt1asCeZ5qcbIGZwixj7Hgsi1KsfhvMLgY4uXqO3vcUxmPHEy/3wzFJ2
r+PpytgTdpSxseE6DvIAPVMmtlAkysXR50u50UsyOwQelfvAiMfgu8jVbZd1dfD8
bt7iAIkBKKg59iseAgYhkHtHRfCrDwKEcY6jyYUYO2oa20SqnKmrdLNzL1lDzIAb
4+kq+OeHilZUaJpKCNrik7hlTNQd42yvWuvuP+fwh2zcYCml6h7egbiVwhwaJPcT
bx+aQUZWP06qBBljIJirxERUnvMuT3rMjinB1HvZFMTOzelkkmq8yRVigHWyopYP
RJv0fBR5S4SgWbfnMeGQeQBUNmL02n8z5Kd78a20eRArC8dsnC4YQqOaZAY3DxB6
8hwkDXsidKZitNmgrKK1RbjXQ1h3LKO4+WN+F70dcNrb+mpWMrMgtBk4ZcKdF9Gg
Swymf82jEJbyY1tuapXFvzEwZ7hRYswJQYRwXpqSXeHg9IpMcSHpjnEeH0G9J0pM
8tskFaOuxJTHpxCQpUqIdLhYcFzAhCsFTBgtS0B0AMwOW3JFIib+mAmCryRX+/cZ
xFO4MthnOBhOLuoWOPfLjQR+pRr7K/9EZVN0ZgOi4konBkqMy+tWFUyvGdtoPsu6
hRSGqWd7jxxWqprL7XnA6ZjZepS0B+f54ebWNVcoK7xosij8OwLPFHvHFydJoJKV
bH+kUOCkO29HUPR6vlImbBAjMcthGi4i68Zepo1aR9Hz2NUoGISi/RRDmYNIeTAF
Z02Nrwk1vHqEipBzFt9Cr80aQWeDFy+xukLsrogQEt651O0xxRvkIgnnR3+veO3p
ocfTg0FX+owhztkdrmDRLAlVTHfWKlBXm55cE2ss1/in4axLEbBgmY9DIiq1VcOW
GZvPC+OENGDopx9p4D1XWZSM0yHwCy1B8lsXjLlhzcFfDLZHkYhrnP2rEiItQ2Oi
AwA6hcs17Y6ROiNKwPFviU96QeYdenLd+OY41K8nGj+B0ZCx2yyCNuegCMOq74+8
f5bkOeo4koeyt9/tKPvWXSXgxmwh9CZn8XTN2ZkwNafrp/Wl2ZeM5MWZ3+s1ZQYF
MPAeRXnz1RaAWhZrT2jkdl678+MMjqNSutkHQuynk3UTDSWF6gKChwjz8CdRJNtt
Dp2Q5riANk1nB6SbwXq2NgsR+p0eMfrWNLTK8+wn/GipUBLi7Iz8ZpIiIJf/a5yJ
KHxtVNdWJJOIZwRuTAdc8Q/Xnrgr9FjLX8zO+AHu0mUfX5smV5BPowPIlG5s2SLy
8muGSGWajqFyUl3wJ0BqUf667Oe+F42EftLAPoU8fy2IEUgI8teuw6xBCmZfbCwK
BrRniF1ZXK8J25xQWm8iZfH0X56GJJ/qzdnPBi3azCbdolJv/GMEKkD7KW5a1YHw
sscZ0sK9JTZxzGO9gtrB9kiHqsrr30cTMG+f10skS5Pq+KE36wotaWxiErbbphdU
FDXRQIXU78KiJNRBgbGoVjKizu8W9NBsWEA74Zs25P8ffDsdwCoSExgtRO6DFNOk
ByvDXyrwsYoA/Ci6G4sZ1AALSvuzUoSuFeGtWBI91y80Dc2iNpcrKwyLdKPqheSI
ryEud0EKCEWs+55atG097T305KyjSz81BkYFzSQuaS8Rj8r7npzw+8wwHUHjJnJi
hr/fhz5sZ+PsnhuNg1YzdwgTeNpHiOaUH9BUgFAM7FmibfOCUTuFsj79/UnLuQwc
8o0kcr7gLNeEbvJR1n7virNxkVmVc6zGARpsFdgKZQ+Se0yYr+kGidKyU9qMFzIn
YDGEHsS8uNIObVem0K4TfEmiqgPcrPYgPuw9PIGfng5kiRNMUNasACmznUweqI3Y
AVN7qkX/d8HivQp12TFgM0ES0o3LmLVORAEOzu+luBpKUz+oMMA8/iWTShklgtDK
utoVkPAqIzGGFWfPMVwD7J3XEOl6PYmd8d+XEj9ghrw6jQyxzZRol/A72g/INAzI
PsQlv7n6HCVH1NoiR9N8IK0GJFfu8oSzOw5ujs5MoYYZdCG4eiI6SK6LdhW6H4GK
QIEwHv3/11Upe1pZ5cTPEAJuEMdeQ2zK5wWXK90uPSKL6ELJPF5Coqmbjt04Mcjd
hQwiNudFuBgPIlfWOtvYrnU3N/wjZ2fk7vyq1+FbQmW+u/FjX/se0rEavivfs9de
CiS+q/Tji4GxIzSfkeQ/wWw5ojZDt9Vq1yffbQNCa4w+Kn75hKrBw+Al/b9sjhsB
WfmElCV4i4jGSzhaMI0/g3izsFLlu1ZxkV7jRLowyw2Z2w1s5LCEbbLXeaRSH17L
H1skJ4TiTBggvTHyQpvqZWhwZNB/0b33lxX0AcSvQ+e/NF6PSMG6ZsiFSJWcdYQK
ClobfG1B72m2R5gxX6TDIW5GSIaNQ+Z63Y7puS8+DsPXPILt5TIlP4ptQ/eUSRU1
vws817ZRl9aTw598aR/BXBCwjZu3B6wXLADHHv3LtYNp68UL1SXZjQgsUxh/B3Oa
ReKc7uIliulVlha3o7zx7Rf0cfLUiWJsRpr/Qlw8zJF4y0lqcPZMSfq70W+Tcnmr
R8GA14eNtBapQ2mZ5REI38HwUVyQg8CQ4UH7HHBYqFiUis+S3LaCFw6mAhU1h33L
dtSDvf2zm33epIc+O57lB38LikzVB+hIhwlRXltfiwb7Qkgs7FLhuFzka9AukiJB
Ny+YXjHIn4y3gft7ed+1s7n3a9xJt/SWOG24tLMTynCEYTZ34ssrJPeVwHbxa0Us
c8w8Cmt+oR7j1fEcRmqnFAz88AFHHY/PL2+HYn6j4wkAlDCiXQBLCKoNXBz5sh/K
fO8l/W80tQBkMtC9kua96fTuvxSy440NeafTd97bry21pioDGN2bxgTmfSpqdq4r
QjlKGcd4TyFBRqFHg9mOV7fMHXDzNyUWYEnIdowqyOdDaqbpqjER+kD4Vm6qkTsF
fyqL8L0IT/QAopB4xbFbUt/9M5uXCzlqvkGfaf3LS/+9yAuY7dn7mbttHkdgafDl
oK8sGBzlApV6MF0OJQK3F4MN8khTQPYgr1V8/dqG8xrHPNzMi4bxa3TWak+jSb7N
61zD7/Uyet2Is6LsJMKCVdHGewWrmUQ4pIisBaA9nYHCvgT2bPqJZ2GVZ4WyTcw3
anyKPKYVnMFp6X0f1S5PKTnW2nPBsoUF6KRX8G1D49ufpI/mdUFCioqxtN772P/A
hLNnTlD+0SjFGfjlU0E80N4T2g9/XlCeZqGc1ielhjHCy+nCiaNyfukQcwnBYOtW
H5YXFLlOc3mZWMHs/b3I7RrM4+Va2Qm5JmcXiVziYrulqeqCQBpwJ3F/qQR5jqBa
PXilVQ6/gmexxtCojZ9WZF7MavnLDGeQOb6cu/tLL0jmTYUulGBBDEXSrwKMPSsD
7TVl7Q7kFO0giurdr24lkZHugMiweWJqfbjbRXT6VuPOGISpMLtN8TUWc6ohwhb3
2IiRPBONpT9u2Hj6d9BMdblqNcz80Mdzi+glXSqExZVPh2UxYqY27fec5FPcDckV
pQfqDznlJy5tKbGCdgDtX8gqR7KoyKz2QXzxhYPpHBIruOzzAo0EldZkoL72oU/s
WddpywzqJVR0xX4Oecbf0JQN3KMZLJD4+A3UWkQkxvQUcW0DmDS+CbG41De2Ii2f
0YxfhavNqx14vMKGR0FQTv6aWfeXxtDhbtNsdXB9eiFLILQfslRsso69k0rCazj0
4XMXcuhE240qsJpX5Jt6o4CTithNBHijXb3KrcLQ0NAH0Tjmly8DEEvz2gbfyn2v
Vv7s4lBoZqdJiH5o31XWWWWd9UDmt8iv00AIPdp50DxZwioM7bbh8Pfi890ntEz3
Rg+yR22h5psGOsOdXVj1WhZXplQFnlmC2vOnDPwfnK5tcF9g49sRK90y36ja/4cJ
4Aml1Z0Lwfi9tzqK4QNQMRfNyBttwlXqB2FW3lEjolddJekP604RD/WfuPysHQNW
LZrms2qq0cvcXYFM7hUF8IcoedvBIec5N39eObHs4HuB5mha7wM/G2Tf7K8nrKOz
1RXCpRFkdDEQH4hX/TrzV9tHDl2zibsJCg8DjctpT49SyjLLOxTNjdIxzNhJKG8k
E6lNy0sPyfpFIpqnvXmbQETql5st3Czjod8XQLVeapGDWbfBst62b2y6wmgmL/vT
qkCkRKTy32mjQ/fyifpk9oFvop4k63JBI0Zqr7ZTSdrb5NjV0Ucofht+Xi+rhMlr
1JjFr/2O9Asbogyt31YW3Z7rRZRYIm/3wtPvseMsH8itNYWPmitcTTI4iRuA6cO6
DSfeMOLb38Li7tFh3wDUWtZWQF5g6a1VJHewJ3jUxJFk89f3j0aZl7FWB1warlmI
E5loMtcvkHGX9XFqQpZlWF3l/Q0o5BOZVETynybxMhxe8CvSnWC5D3XnZY0KnLJQ
hL5/uBnjElIjy29PNcTijZNSgTSrem4CX6Kaze1Cbz8yyNjWd7WczajJacXGdoBO
hEm7bhegpqoVK2WVC6oYtDtA+g23fDu4vKk/IZ8s8zfOjqXW90146Eb/rOQjk1XD
oYVnURslVMJFQQPggWttz5qWVKZb5lu6N9uok9Ezy54d/hdVTKLjLo8cQoBufobw
oLPFsXorMNH5U0Wf3eIuu/7PcFOindaSHQCW+MiAN/rLnwbXw3XdcvR9PwQNVfa6
1JnbPJ++pMuYpo8OchV10hCn2vCWe2GsKJX6Vh3eTXe2J3J/pXMeHFrEw/Ojcg0/
kRtVGj4Pr5DE4xFSmJgSY9arOzHsocJovHi/ax75ZIAF5ZI+d2iymlXCPptKl4nH
21XBSnlgjsKS7em+/cOxhCsE13v9xUMdvsjffBW3zDNu9QjDujLjT8MLCixZDMOa
sHXVq/qifQSZvI8k/O7fwllyW0X1O95RmNEE8bRO2CX0Pz+m5bIcV3hIKIbwFS7t
Aeas1sp92FnmhmPhmFTjpJBzzGZv0EDLNEftkOzbxcSyRSiJT4sZLfE5pzPuXQXj
BNJQJFbBwhOqHLKkVjWilPclD6gaC5l4RAKpXagJcucFAuhB+APtrC6R7at4p/Li
eqygqcpoTAruFz2EIvpvdQgVh8TFqOHoYktlYYt7ohlWrLcJUD+lF3JL08bUGUs2
wNp+VbwRqz8U+5Bw1be20r5HhnFM5VQezQm2AXT7DgTl4u4KluvdhDU/+kLNKOeQ
BxwuLqeFhZUWSiVq1w7Zxu3ZkOAks6kRuHEBwpj1I7sZGWZq6LHfZaJTm7R7ZDEI
4lKB33Ew5ysJoYp/vnna3jETAxuGgaoo1/iHXKU9iVsB218vNuUYfX91GbyuOezn
pG6rXkzSMxzmGn0pOB4KZUgT/6qcMcIbLCVikyoQmVT1wc7u0yPkkMFsbqg/Up1m
kGG6H147nJ7njv0mf6ENNTYv2EnkBP7vumcmcl4Wm8oqE7ZNRe8yn3uYLxvwt5vH
UZhqYtkANczzPp1ZM2RnjK0Vkxo4zq9gRO1xFpOo0zu/QC+/gEHqot8wWkV8QtMu
WiobNLqy6rRaYBe1SbclfVO72+zucwPxWSOywMfGpsTXN9vIhdjFJpPnu3hkkQci
7ke3RX3+Yno2aWLd4OS/4ju1jh6+4w8GExuwsY+Sj1NXp5Ws4bKWDyIQFBITEQ4e
fBAZH8e6jhL7gIZ5zZJzhLD7d8woPTAvpTJDOuCEURHVNL5KlRJHcRe4oxCt0dng
a07WY56DsGJ2hJSr0/jlK+uKbmlUW4L3k4lPFBZcxZJ/ubg1+U6i9PuB5b9PjqGU
SPxoN+LgoEhQP+t79Pj4a25RVtnGq74MLYQlNXbkH6FMC3teoB4XDElo7oUliG2n
F0zNyn41h9BCNJpi77DYg/AJSj0Ez1j/0Hya1Ryg5q/gHY7Hl087J/cKGknO9CRp
mNlX7/K8Xb1X1ac0PRI/m8inkTKimCoo5oRyV50j3tlvjOA1Ak/btEOkLZ1kJVNj
+ZINVC0Yj8Gc/1Vseht/BM3pRmzrP56EedQRxNEII+FjP9A6ok1LI3QmoFGy8WjG
WebczbacmLlBsG3RxolH6/gImM1bzOPahJ1LUCczxAzAyRRMIJmA/zZMQ4/WociG
heeOXq6g2YMuMazmv7GjlOuJbSnGs6lmWacHqVMgsDJCWDvZbwErajtbm8On71rH
xFL0pUwWgRbb6e7fx9WuVTBz/u7tCOqrupsFFOU5GJZbGRs9obgQzJDauSEKDRiR
57N3upapK09vhBm7slf/oQdXk7nYgvwAck2vSt+lB0ZlONHU3wxdGD1shWHjTEO7
WbtdZaukogpb/SivIFTO2KPiJ2tdt6s0OXNaKixK8swwECZQVl5M4t67SVrrRccU
dvHQaggV5mWwNBNpF2rhPFt2Xyu3Lgf5LVRsx0ykKr1pIouwK43pyU6oS4re6I45
NRVu5XDKoL3+C7P0w3LON6iBKs0hbYQdGJRsyYFibaKdeaRGuMtGSSmUA2ipB2fe
9F9EhnimMq9FNhfNeqUBz/a6xq+EeoaUvryu0yVfy/vb/A5HbWXkq3GICaewBUZr
NRjkxPxOhHr517qFAVamZ2IFctrKAJHVPfkbFlaNjg0hO5z2UdrAffKT9A8YyxfL
v9Kbvn7NyvhsCRhWzozFwvSph5TnThWsirhJe2O29+Ohnm2OkztXzHcoF8/Buda0
mFiJpZCPEZ9uVrSuQRp5nWSRv0f4fvTL4htOa+3x0IrYpOonqUW5J3M8kCyvkJWJ
v/WvYawYGjDPxvbOCvYg5Fe6DByr+lC7lby4QyM98ATQ3SnY4GaBTy8gzZuEg6yw
WDhN2A5K9DmmPPF1brBUs+xhK6ENO9staQyAHaBLRgY/dmoi8nkc6avbRWxdVFiB
JGAX1zMsvXDB1KPjQOcHmvsscgyGqW7CSQ6TNfB9+0mmtcIHfgbbkXlsFU3zp6qA
fHAFK79bhcNAkAIHy/Ao6P6rOiu8wzIzXE4y+h/k8OlUvia5OGk9n92uTEFmBZts
RYE9+4XfSq+CAYjLyt9U2Jl+CwJrwqqoea2c7FfLuKUCZ/jI445ingc4S6BKzHho
pX++0WVAKZuruEFKNB56jU6utyt+SiZkoacU9HiAnMX1BgqKcQbJRQVKgKbILey4
9yI5NEJ2AN1mIoemb3JmMWpwm0IhUCFvlHc9abx8ExrH1IMdqC7ovXGWpu1cQRrz
kAFcaY7dkdzcr2BkWCINdmXTrTEFEGU7OtGshozFnd/yOdFjRfVqmPRAI/HFxtrS
l0T36TfmxfLUwS7yhC/bve1vcQSLFk2m8BPlAS+BtjMBxE4aRpj/f3Y5wDgBcXkI
jrs+4njW6kMrC4qB+IhoISiUIU+/5ylJ5GEzoXkGN5NPFUWsJjQegIexMGFjZ/ne
rXohRwDmx+mG0ABw3Cp2+gEnsY91cJ8d0z/5G8ZJOBQP+C6ZsGtprD74ezxkO6xe
B+iwq2D4S/p1CnhlEQMQh22LWUO8itmm6RebVOcbFBm1WjZEhtSQEp8+7uaqJk/F
36h8QnaMqdSZl6IabMHGIpeDEE1ZDa7sMtCx+Q1TbGWGriM0CWyCT+zjwRcfGiSK
QCrSEb5VoZVR7Raxshyg19xvnIYN0vspmn+gTU3M/hhVOA261nc8Z0TJSi+6Nmpw
StZhTDNbfPgnOjfbNrikqvGb8gu8x7zSAohR+uNylnsXV+ze25UZozAmcJ18+bDk
zl5jNvP4gIp68DvMNo/aTIjoZV3vSYRLONr3R+DWn4kc4PqLJEtg4a9ne0HeMnY8
QpFoEsiIuS/I78ZG7cOWCUi4JG1jmMUF1denDcE9GTpzwMEdrji9QnKRdDjNmzpf
qyrR+yttXKOBRmVB5d0Wy1F06lttBS6vCweDoA34QDi80E5tYDUBAizpokIXbVyk
p6affwv6SHAxAjm/79vedbJ8RIG5iVmu+SszgwYuWfV2wEHmXO8hiPiytBrX0hqW
qIxP2TwVsMKMUx2HadI8O36affZN2MLmCrgXV8mNuJuJxAuzO2MN+q66vW2aJ/Kb
XqjsVPmznp8MBu7PpkzNBgBxoZGAokQV3AWyxY0mZOOEhV2FVWaye/YYlx4lHE0z
tvQKRkkBM3FfKriyT6X8j/TrPCjBgQHJBmMuayzYIvDSSEl1jwIMvLF0EoNwnW1I
mVI/80lHJeIBG6+VdmZg+CwG68dlctGg+Y1+FkDYOhC+WJ44sXp6J3WfApKWiWN1
71Xo0MgJ5z9A64o38F5yxAAV1hYifOeMrd/HmdGEXjgm5aAlWWUdR/t7chTY8Wpd
uOaAd48JZqtMFjokKFYxHnyqi1xgdZ4iMLQb9t0XaqiTXn9uvmsevVweAUYsUJSo
C0pHsJIy8YKYsdwnSk4EPnVV6TevFAxTUh2RCFFAcO7RliV2pxW9KfbCDTs0GsKs
QjkUlSplxS3hbSbHD9F8wd6YQUK1BHiFoYkcEROD6d+J05KwHPAtDnewrw+SeMe6
tZKeLbB7T4g7izmwx7jqO43IfS5ZxLY04hV5wu4IhXO3NkZGrKqSrVntAarJv0Hs
PqN1iUYqtcRn/7RRUWn/LQ77uwE28Ae24Vv0cYuAqPFtAaGWwPEP/H8dKKtYpPvX
OB7o0nOReOVhHx4XFAWLNDAw99H38dTZ7IsUt3yNQXeDbiZb2zBOCc7hO2mH1vMH
EgvVItwwZSFXSQ9r0Ar6YzfERIVlsAxImhW23jJAieLD7GVxbeS6yz9d08vUoFuR
KtGBGRa27kRYTGU1u5ViT7Www+isAq7xSr+7/D6RL/RSnubSLz5Hk474FQ2ilBI/
/MguunqvpmSIuwmP9xk/UxX3fwSWX51ypJwXhDOxwwg32C8mFgGOdQ4PsPSer91e
61P96mcF1nmR2zERmh8tk5mOjNYetePjmthGaCNNcBzbUaQC09Q8/UP8ewuG0BTG
HlGUjwVu9gbkTEAX89FaRLaP6Yiw7r5esX8jPOxxkhmfGqSAazAHz4s5S4mB1kAl
8Ek9pHEsIolroEfmwec9hRcaz5m0K61yknSFWUT4tFQZOpjPm6dVp7WZ9U29aKSI
TczSFg4sKzxkTSUY5AqI7UerHpKkm4H1jO9rtupdrk+esBLK+MZ6aO5eSl3kStSG
rFkiviatD3lEngADXagwjSep2QvT6mHqVDVtz89sMV+OYaFSCfXh45XKuJVsMIoY
oOulK57piMfytxprmLe4bux13VcXS/zzXaAjuY0Blq452D7AUndXuD7ib6OxmAJq
FKa+BRbc1GMo2Edh3KQfMmkrDUm/zNkQ1FvzsofrenKkxX/sylyUd8SEg9b4e8Kh
4QaKgk/0bsv/4Bf1m8GoHIQ2KpCRX17f9cv8RXPrrCwB0easLW+BLLRulZvX0U7m
ZRSI7RjROXzEDXzzyjK0Ud8FUm/FChgSTFW0jRguK+c+RIGp40vqJphjL+eUVfD6
rTHF4Wwk/SXuEjV6h9wXZnRi2XyU4avsOb8C13AekIZ70Saw0cXzwhzUvkbX+RUN
lBuReEJT6dRw6NW27ex0CxsawY2zF4seYiQEEE4+1E4uIGBGe3WEp5D22TT808Ta
+tMo2ZTxD9/r0D0SRQ8IWXa3jBggHejDyaFUBq7GZ+uap7fsvlWIgYl43wWAnflS
H1oC2NV/wOb2o0LyBRUrKjbSa2UuH5p19Eq9MnSIT+vJYrRHy4uOA11FU1sFJ4LE
Ve1elzUFvtZIYAt4dPDWP42AyMXAx+DMEj4QBC3x8EodOX3rnvyB8W0KkcmXKy9Z
FclzetsBkLxsGycUYUFvY0Vz8HQ/f7LzZTwkbV9NaTHIRwO60H8KTfPDN4r65w7+
mKuzTs26TA3CLBPk6tp7t07WsbAplXS/j1qIiRVI6nK9y6k6rQDfdrWnt0o1ctyx
sZraSr3KhAn/5v/Gqzwjn+Tzug0kD3FqbTxuyryQoWs1IL05ThVZ6SI9bjh+/Sin
/PKLSk3yrDGLgR4ZTgaViC7MU+oxePTDvFTx9kJZLSX7q0DTI2UJFwN+6ymvxnNh
pnRItD1wvp7LV9UmPdlhfNFfA13gZWDep0sStUB6psO9wMVyMKwrOhrSdiLyrFqg
fzuNApc5p58BbdE55NRwQ14xtrQUDnPoqvnNKi0meFo29diGg2mOVpZ2emYOrSUb
1IcGPsXHLC+TwjQf3TwZvEzCsR6znGAQP+m8bG7V5U+lRIpBwmSkP/HIxKgQEic+
dQTOUWkCHdHmbGvEp1v2vcIaf6R1FcgyGRnVhJpLnwRUQ7BDh1qWBvJjyNrIdyIC
ck36f8inzFISaJyZdiuL2IPbJaV44FuU+TBEWP0xuuBkLHYX4vzbde/vdzDI5OoP
oHSQggV4eDlLubol/0sF3X4N/23y5yK6vOPYUMWqOE1847FCie0kcZSMVm/eHGEb
p7N/318EGXHVW+AvfA7aJc0lgui9Dw6BlKWsfqe2tHp/FkVD8yoNFbldzpPPQpqy
PKEBi08G6I9B7LjXqa49z1AtUJKzEYivFRs2/Go1ndD7vO28f3nw9iFUfOcAT3lx
ggI05i0nAxT9Zk/H61JUGK1IeGw7XkcT4qjQkbqRoN6j4+rx4Nn+DTZHbEowyMKX
heiY5BRDeTAGokDSY9DkTgGwJfAfepYdH6W58Z4qtx1lA/fWTZ42TN1laVFVfYnr
soopsZtRppkilxn4Tm72Q568QkxtnDXDYiLJATL2bGy03hst310aPBHvFs3QcDx0
NLMZCYKQzg/hxMDWZaxb3jdV35CgqrSVFWLF7QEHEQzu4riVZpZbgKX/ETeUGh8v
E5Gu6fy4tRPnRG6KmvXFOcLT/SplIQLAu97MjGBOJcqRLiM0duAR5mFwh/VdpPhr
FC+gngKdw2CxTR3LCYldaOCGiNSBTYbmz+ECTKX8QI4L3Gewd8qjc+RT8OQDXvv4
YEEuHPHHhuUsF3VHIe3M/R+7Mv93eaFsp5+g/j6it+jT3Y6snY9rFWI0A6xr9Kc6
r3H0gpclOWOwy+Z5UxGggU92hiLF+r0UOCT2ICyIywobNo2KZ37d+rxEyAybZHzg
rVzfqbRglUpwrNIqA52rQgpA175vWJw/5/AjRVPoZ0bPxQUeL7Xkp9kUFJbSTfjB
UIMIKhMBNvZEknSNhVU234f2ikRU0BNp4VSAaSh0gX9ibbdCw0rB/qZyPJZPObVL
Kn1ch/IWVadj/kADzk9IP63Gvh8H2cnicAnaLIfP7X2Z+9IiF33SlDXrWm+XCsnZ
BrV3hKjx0znx9BdJlxzFyaypdcL14Fz1AZQNEZzoS7hszDx5MUB44Nw60yu02ygs
Ut+t/mcvBfkZvcrYBhwOZipLraPiiSizrqGVB9oY4HYYpV4Ogg7nwSenl4+EfjLW
3tl6b9gy/vYCREkltiL+XylTDdN/vWSn7FQDFZC+LvGI8nje7eaL4K6w2TqZsxTf
ai9ic60akwDEMYfK7Sgs7+NOuHDGqSEAAozv1ReISZBzmeJwwTwgFFwYb1esw/KC
jN6PH7dOA7jZnK+A++dWj35uw0rrOCkV4Lifr17We3+VuDDvk5m8AVJN4F+ktVTF
Hi2QAdYqGyyYsWA/qgGvqC8MnVH6SdrYrhcQeIERKfw4EGBfB6UGksR0DgQMkkJ0
WQv31/xwxGsoAXS61aBmGrv3zkeUuEpj+erPKiSasf/N1Spb/8jJH5Nvl3WqSsVR
omwDbIXc73BBTrknsRxjqrtoFwNw8efiL9ttBeuBUg7pgna5zmgN+gzZRSQZJ7Iy
c+VLP9KZyObVu6LI1rdS9kZ6X0rqaFmqgISvBI8OJncXwkeKQhoOBq/k7eB1JdIz
/MgBHXws/5aDF2oBPG1brTApCAh/QQ2Da0a64HMmKtIj3f3OJnqvao/66MXl0kL4
19IkMO6UYFPmJGc8AZhX17eurViWtO0mK0NCLBMfFp9dRCmbb5ZJTRTwljl4C7s/
ioZ8f+PShN5YJ+pf8JsdY4Y9fHOvCZ9Wu7DSe5s3zGwXLRmZ3nCa5RX3QnI0ldVg
G7gYCFUF6r4N5ClislqJvS2H+BScNfbBj9x4x1TGZAH5izqj+Q6rezC70Z6khK4Z
434gZL6Z2ROdHFgI8tgng/4Md+SeettuZWdXynr0ljoIil104IP27ikB79XaB7XL
COgCucpW3qb/wnUt8Q07LQmnUvNRiuVNXciH8pJQaLswasOppqRKbRXkAzsvSIoU
z4ihZVIsiLAa5Q2WeHXDuh4S72KwzVP1r/fVQwTuXMSm4ttVgInqwyB7uDXMJVdF
bWPmW+nbnLsNkY2/hUiMvF3akSyiA5oeshzL396XSSbkjnuCkCh+VdXO/9+mt9GH
ADj6qnZY95vLgJS1QeVWRHmf8oI1IrIvtVvkr0ymCK3CvykB1HYWCWwge2f3CEaz
FBetNYU0sVe7RsZ3YFkaNoPAgPpFcVPZb5EzzAtI35PQGN2lGI9MHc4ByGNmCaZC
Y7JjgEsanRrwg35Fx825VgLEnoRQOb5eIg7nU0YtPx6fl1z6tTGpBaX8+BWNuXIp
AT2xIbGHavbl2qUbbXacvftC2+5UXqpAbcI0E0DlZmLnCm1URJkuChXcXcBF2G2G
EM3mlj8TvkZakAitbKosRddNnyMTOzZWTIR2mBMDr4ybl4dVnn94k/hivm4ZdWR1
jnOz30B75ojOZA7VgdG7XBr+la2AGbb24ISFbfHe3lOcxdn9DCvQvJqCrOB/AQuv
P2ClqFfCgPIUujqsqS8npmvyABxVVPPIdeBlVenrf5EIaC1T+Ce9W+SpnNgVHVVw
xvnj6GA3Ph3BVdsmU3yyLMMKHFdhzgmJUVSejsLa1Psharegfo8fIcrhv/T9sJrs
Xtb7hScQV9vtRGOCYqInPA1gflUZeCH2edzirCHxwD1m7MHfxzuy7kZ6Fwg3DThN
fjx/fmWvSNUFYRRQQ+qM+2eX3RoRq3kyZkzaGOScsmGP3yE+vw7aMmPd9xnRTfmB
j8oWOmy7cYTSjto/ngvkg6Y9235CohdjSW32sttSgyMHt45zVk0uAFCy9/UC6rZX
1CvRTcCLE0vxzZXT9Jg/ElOg4oPUnYfPkOXgQ+Kk0v0c7MmNfGDhOWnv9kwSw/FK
LF1a/749yv6ooqV6p9zL4JZZqo0MadfeXsEk7Mz3QzQJ4HEx0mlajllI4alCHyGs
bICSMP4ItuUst61NeNr0iTQfW9cSKo3eyRY//3go4n9w0Qpcous32S5oAvdVd3ai
EzSeJOClHO2n/ynJTZ00Q+ArjMsRYY0ncBpQ6f38sq7B2ZIffzvsmOACkkCb7er+
iDS6rEyw4nN2WIAC3hTGyn9p83Is34jaPabDY2c4MUFQvUSFz0Ux54Iq/Wi/KJf4
1RQ4mzX0/pQyC23tZwnmfNBgBOWvi/waPklGUT+i7eFHq78tlkQHXWxX5V67Wvk9
7AADLXzM2cn3nzbnCe2cFH/mr+snHqAwIej+ENhVc8IHeAdqWUIQZ2PX4Ai1lgN1
vANvv1gXBC8f/idh5BL94wzajsbPHh4boghOv/SDSeuUD5grRVLmFvOioTdoVLMG
JeEz46C5eX/L3zPaQ2TtI6QVaGLmjxLurO2pToRFYf5EdqO4PnoyCNCLP3iyX6qG
HFJK/e9xxiNKP/IxUILeBeMGoHHraMhkZTed7LMcSYNlqxFRox4aCOy565MzOCjK
wCNlNS6IZQnytr3VD3xfOy6Epchm9tRVABViLuNfydnrPGmi8sw7I1hEFtk6eomr
7yIk7GAw9jx02TAfxalX5trheZSRpLL4slXuFhdPxGm7FgW/OksN8zEyYHMfMQr5
Asr/sNzXqKre+CVafeZ348711FaTZRswd1JRlvQqIKW4ToZL9Xz+avOh9QkZW8mC
GnzwT0d0TK/LKDHvLQkKEZbYpUOB1S/0eBmnZgmlpVphQVhGmja3vVApNc1zcsUJ
VJgPywKkcM88KpkHGumgZuL4g3nc9v8cl8OXxIpZemhjVwhRpGyqRESH3Re0iKdr
8NPiAO3caSpneTlccQ0X5fBpHQw5LzDNr+zIwGpAARfPtUTS9aIaIIrJRzA+R9We
6RIjLai/SeuIj5v9Q+KCy/gmJvfvsghgEUWinYFaSXoDt0QVgcKudjLanYJ+Eg2Z
9vjWtxXOgYnQOdwMtElL6C9DLpkKOkf6riXERDZCM2+eEqwtGaXuwfVf6Q2UO3QT
uo0xWx3I2Puqjb7l44249Iv1lturooBGKUXSLHZk+8g7RGf5458zyd4hnNoCAror
E261UIc8qMnSJ9uTQ0ozjEb2UkfBIYa6wApwj+IwR0d8NwwcxXACIHef1YH3xthe
+39hLOeFGmFWAeL71grND4NP0fEosh7BssfQp+FBNSW5oFhV3dSNztd1ZJRbsjEA
oCj1Y7nd96u4BOko30rzOX5h6aktRtQgqAb5sIyZymj7kkVov4zxDEVNya1/AUZ6
NYzB4V2NFgjmD8QYwdjjzFDoEwwK3Q8WCkwB5NcaQqmcNPnJYZWhaOKVCyR6vXRJ
nU/G4pFMPKfirAFRba2D7pk1ney3fmudXkunMm0Cb69/2QC+KWE4VCz1yV6nGouJ
hzWMrpF9YzBFjWp5jri6Hl22gbf3EzGi2bRH2LnSZ7VfJgtP+uYPL4oH221vQw6A
Htb2KO7P6bslQVPg/5EjP0DcNqrNRhGGdC+KZdYnxhJCbDEwJD+7Bd4sxnkQSyc1
493jY9Na5uEF4wq/dvDWtTHhxH8Mobw/XuUSmIOAuwGiI7U64H4kvo7eEF5coA7L
tReif9dENioCw2l/2Kkd2M4/LyFlo33hu7HKtF3f2U+MFM0T9IZfZH+L4PcKglWF
t6Hb7aQnPDkcLxYmUDF+XYK83SKFdrOpdNvGsgW6NBvVTl/ibmNbpamQeidLtFVy
/WC3Vman3RmMDh8gKNxvr0Myul8iYKIOAk4Z4ctTolKrJTiFcxLAYnRXVDL0+uNT
pISZmEa5nU63ftJOPxnmucoeF6BL7DbtYsQjVzovKgyoGxdNNO83K+4UsMjupYSg
7DNRpJl7rG4IhkE+E+DQhvKiIHLHLVZ0iA1Z/kC6lqdbuQsK28NazSMGnBfRUPo1
CT7Ko1zXd6XbhelhfiTCvek2CJGPM+l4d3dA9gBGnZQ3Bk5HOShwdDEiJVt9afu5
qAvo+5urIMW/ozN1W6Vets91Yj68E65iOpCUsgZ+Z/MuXiS1lnicaxYabCjyMu5Y
yYG2uUPZGPF9dhVcIpJcYHLK4TNXnjQqff3dhlXMXOjJyB2R8LjNqrNMoweZ9ele
jVAMkm6+2ou8YiBiEPiFckY0ekQXMJNGO2DuOH0Yk2ItqDXnWiz2awy1ah9+Frmp
hXl3QGT6xe+qap+eigKLurph6MNdmHI8FuwTv6WaJfPXdcNDzEEbRVV+QWjhOyN3
m19/ABZ9HsaP4KPSwTJ9jI6LD3zE4EeLutLvYLCyRTQjhF5YD/Nq6455T5eLeuji
9IFLnPHXyafzvts5Gr3ubbKhFCv2zg5N7bj2xhK1P+xRrzTyakHO2NdXMRgJaQ5H
qrRj0NMtmhbo5NxKU7VFpkhGNbSaKywa2TUW/fGOUcztqwmjsHsbX01+fkZnMpJs
L1WFnj8UmqKwUhHFFG3GMwqNcEuKwTnllupOL/+DC4mTFnR7J+GLq0E2hj0RblIs
7DO49VHXd/r/rq2sDQHMRf8a40keugnIIExHesZjtVUFLoOsqyWuw64UztsqC9tq
gdN+ymXmNl6yw7Yv2chf/JM/1U/IUm6Gdg6p6SU7NNLpo1pdx+V7gc9iBnV2r0hD
EtLYrEFNJ/ntNYtNwx5ZOT/5972kPBYrDc2peG1v2XvB0g/i1oWszbz/PoFjdHu8
WMwITXAb9U2GMfZ7RPG1OqoK776U4FZYcnwNLr65vN616OTUruUvZXjok+X2Isie
asG7zrrKjcED8B0P2q2RHhJ6ZSKyzd4jq8HmulwszvgQ3Wycq0PUc6o2i7HdZNi3
2J6iMnxRSWh6oOUJ2sK5lWMw5FWi4cO8GxtndxdPDHe7MzoXyXZjzYSxH5bIWvEJ
jXb1LD6aMFC8MFiJVBqMk7dtG3M/bhz5vV3iK0Ft3MuGGUOF4b7DkEkbFgtnWVRe
JGVJvey8OZFumJ3ll6sRAbYm7XHrK2+094mnHKm4YpylFUK26/woWBK/j6fF8yJ+
gJP5ulNfqoJrIWgdasew79TFq2wSFXHPkicEb7wO1sUmSlYPVrVe4Qpo0bWnOk4H
XedQq3YYMEK+3EobGsA+ZolwDz2wAWm8wGACxaXUkyDxZsRxEdMucgtcupi1w5QO
v9ZT8G5csqD/3c06hqIp4JLbkj1elF5l5sTGR1rse9DxuLBzD5SmJ6L1FGKNfu2O
wiYuH2p1hre2lHHECgCs3vv5R31MIBNZ1MXp78RG7RdnJIQilWW0HfnSG/j1lXKK
m8QZTyv6JK+KDAqhw/4BkWXF3uqhmP6memKKD5gZfitwuLByhUV8+LMNKRmCFkdt
j0QCZjDUtpyn1JXxicHe3TAm6l+eGS8iNBhbjFKYSJuJY+5Jpn61aYkbCcazwD8e
AL+Xjv+abcVM0CkRgukwb1WvKhyXuxrRpvOh8As7zt+gJ1/d+wBsgilxv8I2EyYJ
5QZS2zFRStYWjZZe4JcLnO3u4jJSihWyZGy3RJtYOT4yfeAU600QbC+wKKn50qGr
geqcK9DcDIgT4f+xIidKRqKPezGbZMLlrnLUmHlfmMpwXFttnc2NPa4k94iXTcwO
kPSX7jdmHZeno9FdG2DTtXWjJ1HoWPjUGjD5GqgTeKMcIv9n/GQ4qW6Jwb0nJCQL
O/xecElD4QNMkL5U4Z5nbXpDyiiJNlHn7gjuEQiUWPImggrXDe0Qt798OXXR+2mP
oNNxKTQ1cVAzf/fDdPLC/hP1OG5jhMOzg8Ydr4EkfBnVBM53DAxOvlIqP1k1pegN
1dmiiKocny9jpUPtZ5vdi3Hvn8LbQ+HzxPSwcodyeQP0KgGywqgk4oArz6TGRp/z
ge2EDFMwpdfPx3Xqw3ZH0T5at/KFlC/Yf+H/ZbFsgtVRaOnsxRNFxTy+FH6sPfEd
A/vWReb9EL19jV7dk5OnLhwJin29lyycKnPTRoRUxk/0XdPk/F9vbj3K3vBlUj7T
UHePF79qTW+8HEW5q4DrAXGI9jkm+LggsD+HtsR7uGu8skSVqLe7WnfUfD/Y2wF4
F1Es1jzuzv+PxHv0RwVKj7rX/ChzSM/dF6ppuGfaitQP17DMPt1Rntea0/v+xA4U
0CviM7XH2MYFRY7wNYET2MjBggRuWDlAqUoil4X4l7zRUJzfAs/McL+H6J8lkHwp
J/XJNevO88+7irdKJUtrmi2MKUeNcoT1sNGb+Nh4p0odBCO3gXDFHg+0GxLgDQQR
+Fy4jOUPsdcc/UwfYQtqc5sbMPaiz0pNjn+eFMpPS2hBrUMwWwS1C2oCHqnIFDWf
+1xfOrl5O+4vKeY8gc/f/R/x5BzvO9IK01pDhloeg6HCWqT8W3Qse3vhkeHBHOIc
lW28QOyld+Xs1Y89hVZ1hacW3ZUy8sTSqjhx6ur/NEl+eVn8CXhWJTbngAJrIjul
FNyvyS3Y8PYVam7GBH3u5yy/zhR2fB/9MVrtjDez3Vk48DaJl52vlPESFkb1PYze
Fonc7plZUth2fFxErVjJ07nkMArKlnGXbv5fhXI+aI/FyRkXdBeS+GXqNHagWUEg
CeuI1vn+bCh9tvB+EfIqEFBYLcWsUYZOY+24t/30AcXOWcm3tj4fPnzvt9i6jCWG
axN+ZnIhA1c/KhX5ZsoBHjlJ8Rzb/oK5gOq3ZpfNulRxZq4/3SgsSYUiMjqRkQxJ
6QXd8CULaWA9wzx+jmKzaagAkQV4e98DrweS8fbCQ8W3wN3tTvf2btTE46M31Y9L
HlGF6mRJHoeLUThNZPY6m87pJ05mBCr5sBCoFHjm+JdiScnVLTCodgSNeYeQExfq
oknAhYi6465O9w/dl/9FQSmNXfr9TRTNi2kuf6RT/t5EZJaTjgJgOhG3J3eGnmpK
PtpzX9+MaHyFkXPV2rM6d94Vzy0uXjRDNCGP22UHDY06blpjEPK7YKp+t7OkewsZ
20rDGD1DpqXvuBVk3RWkBLVtr14FegvofCMeI0kCDWCwxeEKCDEZi1IHf7uovkIp
K5/eAlZahaRY16YWoSzUTMChKXjy/hmEEtfpGlzzqxVAY7DLQaG8pc69c/2H4HL8
X3Gu5BI7/kCs/58UZcXbBkRKmeJ9YILexLeP+dogEZVAuQzxO8Xd/BJtI138ob0L
fLd8+2BVqDImQhALf1DqRqCl+jPtuxbj5Xn2W5lQ25XqhA0yq3NfZGrHP9xoHXH0
euz219MUuxg54tghtFdLS0uYUpCoxHwHvCJbbxUm0eCRtV+KMebgurpQtdMoR8uP
BXOX+ZfkZpDU8XNkbMrEh8w4Cd9hB8smOtV4pCC8qLFbD0aJaRj8DT9Uh2lS0qD7
yNGe6wWtqGjDW0I3YqBI78lnW9h3XuNjQs4BAvTTp0j9KAyhhU8X0Oo1pYmEnyoX
myXxRk/prxO9sY9+6if0ibuImUok2ei9V2cZ6GdH1vexZ/j5qciWZhueyK0/J3VS
B/SeAqI/+T+mM/lUZ9CRTz8xJ/ooQdeLoopnsonn8jITbNEuKuWsWJQNE62UZ+SB
q1TqxGmqjB8H/BjQwW+zjLR70y46uR/wyRIzYdCSdNPZNQAVVYhvXCjzZo4+hkE/
rhFDj4JbVID+jcbpdx+Uday4gwaPqZKbSKRSlGsx+pEc/nw+RrMceRQhjGF+PVzp
yYI2oleV2iI4P/XkJLQh+Qb/1cEXjbMBoBK/dk0iRYo/I1rPmASxulpEuPBRjp4O
EphwZBeQ/Mnqki3GVx4bVQD+77UCrsJq6iaq9N5EYCIoR7ID8v61PYykjJplOju1
JRxW8/9KufcBQblMl+l4gSoEYJJrnztm2tJ25rz75TdJs0wsxhtdcgpq2/gWVMCo
90vBevKF2VBslmPd8p0oNDnRIN5fNuf5wSgOgMLFGY4JejAukqBTnMvRGjm54GVa
Fs5hnbFlsu4puJPLYx3jJ0ftVQvyWycBZxYt/BTLLsFYulvZADwjXr9P2Szsqzrh
GSECz4pnbx2wZX2BpOG+DauyltYTrJqjOSanV6OkH7//AjjR1NJLrIWL9hzH85zS
/IgEGrFEuwf765ur3QXRqlK6O7kMxrF8Cbhb2OgDdyjz14JipW6TIsMoEG4GbKiv
YEkddo6dtsxhfaVCuYvj9WNGF+I8lUo6iJSOzxALyXB+hJ7U+GRSCJssl024SGUa
RIadsA6fHYOnTBXWIsMSVHG0WaSUD55jW1WpJEaktUfMCk1vArUqCnvhJBk8uJGL
wYDyWY5Bjq2LSuSGqxmqlbpU7q0LQWJmR/3uUTt5NXvXgRaUlCqCfTySDIpqPccu
9jlsW+WEp1ja1EY0scYxVcAPWpjFuWZNgV7t7AtIRnqLfgOjfq20e6RykGViw5xZ
WuFHk1szyZG6fGaOmR7RYSblnoTEyLFrqBrWCjyfhBczUtA0G13cT9nC+JEkpwR4
rH3Ec0jGjuUZI9hKzYAeESuDdr5L3PQrhjRJsIoP1NVP9s/A2m9Z+pPwItr2IqnW
vKaz6LDk0EgofsFNKC6TUCuaSVDEVgQTJ9bw/nPX/uxBbHdthQDBfPBFyYtFpM30
O+aUD99xHEyWR3JATL6RACKCNb6Xw0RM5luZYuG7VaZaY17DJy1/NK8Q7lwdschq
lP2VULK5zQAOY6uF41d57OgCpCXQkYy6h5rF2Ro1dk+MQvwkQTOdW6usZMIlJ+b+
9C57udvX8bhLtbfTDOErpGfCkIwvw55MtU/3+HCk1XhNEFbVgbUGA4FULgSnNV8n
umr5lRgYN5BW3fEb4Vw2KLAnwIApadbC/lpn0EB+SmShR/zU+XfAFtN43NFt8VkB
KI3E5DN8NUkcbte/I34ylpZi7fmxTSwY1NhuXWBeqPZ/Yh4yaZnQWvvUZIS3zFCQ
3ZGQr/g9IhV55E9JnFS1aZCY3zEHbqJxLWo6KZdBfVTAlHl3CRtnCIly/VeoBot4
qVq9i5eSVP8C3KJaRr6IaqJ3yT5cXOOCFIGz394O3abzfSg/EbAE4NPSJAw4iVcd
7p67pEV/TQ8UFlrgknLkN3bx2+Xx/9eQaxFeJACwhbumWEo7M8da3NWlFYZC4to3
1kKkmn/Kxf8LR8MM1TtN2Bx6YMu68HSaTkRDkdww08R7683mjbFY6RPw2Zb5c6hp
Q1FlzWHAotfogOGXMdqviImU/8Pey2J0B3d6zzwqhOYSW5ptBaehWSt81boIjo5w
417gwm9jTS/lehJ+AupftwD01RV1YzMp7Z8OcWbmWZT65WVPvW11jzTQsSoe14oH
o0+RnSjiy7uSLCqOqe0SOL3CpJAg6bo5cKStgRzPXCrVW7x0ZW5FRG1wEid/yA+7
QUCDaQsnBBF87rPifspTWLAyCIrdu1xHvkcQ0yWVHtQOAmYwVvA+klYDGVwsD8nW
glfmON0/QUxxjQskfVkIup8WhlZ/C23v7DR81kStI+ELvluZQ03ohAN3zBtmnVr1
LQF9WO8hXPlP3GwBmcNucyhztstoykAlKWEdmRfQZcrWOVSe1dsySm3wdTqUfYz0
a1hmfdYbNCH+lgW1a1ujYffY3e15s1GzZiufK7+SLTrIMo8dcIjpZGg84sO7jKLj
30xq03GiRr84hfaOth2nvpuOme27XmDxDjfbWoR50JV9nsOnhoMedFSYnZgw+8IU
BQ+kssgruiVaF+vE5VR+qTbdfSJJY+kR28+TmmqDwgafCa1wJtfvPHeQstwvCif1
OWRZJmVjEOfpgP0zLvRM0A6IBhPZqbOnnDoEu11cCmAi73/zXoqWFdTAuj/L36Qc
O2wY6bMheJie/ZEMs9szA5KO6BC9CgZc32nZLT82gXiTOSVG4ol8shMTrZJwGvyS
lpB/A0b8EHSxzIFA2pMnqSBwDXpaDqOBZwHoCtEOkf9i+Z4MfjlDLbN1LykULm9K
ZA97sFBuxhxN4EtWdovRiwiL+utUzV/taU3Z2YWdhMJxF0pho8cmYdnNKAhd9OJQ
eOPmlHM3c9KzccdOXyAJYMD2zfSvSJTweq/OZQ0oKZX70NaCiF3xJ2RouV5fyDS/
kgP/JGGnrIttXW3dEBwhz0Y8BQdd6q6c9kLBYanrNgSGOoPy8DSynOBKVohN0bb7
6aivkievqhZzkcf+DAU0PSEQGG4XMBC6t1mkyRtz0447DDYmvWe2sRtpiqJ4SBDo
u/VlbKvyuR2tXJ+fFoUmo1WY2jwiZgR9GxUfFk+5HmFDP5kBM1mALG27Z56OO/by
umtHIpp3F/Wne64Na7PNj+/KalxQsTQP641H4809PpOx0RduzQkiQBcZfjPfxdCS
SWtFg/ST2e/gkesVJJH7v3FEJA1Yr/qDtJ+mywzBJ64034qKlxNXD5o8dH8hbQtt
SowDQf3cmLq3RDOZrBY8NgPFLej+nNn4J9bl5doRPRQ3uubDNixJ3OovGbXt6rsP
YqKAOIKk912xxdvPChAEJwqWpBDsibn0RUac3uts0BizuGILQno+4kqrCqNRADeD
g6zDG4jeFyjCXolGZekYS3Ut/jhVAo6v7NiOhR0uCIgHj2vwLNBaHrUTS/uFYLGC
9A5vD1mTdZY/lmiASf7g5SL/keBAkWhAHAXoVqb4xthcfoNG1rrmbrcDi02j4v95
y9Za9Bj2nxUSmRgkMBCjkuDQfUywfocOvCKTAa+WFPYWUlfiftHbSEl2mmXK+Btl
xk9rzjuiA7fcm5Oqb4H+jrbgIekKg9IzJut8Qk1I9Eg0GUIoV2VSt1w0aXcIRbfS
5S45Z9STv8lraGZZK+7KUvZIOdNZrTekpPTmRH+o3HrKWJRSlbuje74kfv1dpdtW
jjB296qmjU5AmK2xtMRLpfod0pt0YOJuEn7qihEyybZBEO7PQlNdN85Gwgb3QFcZ
qGE4qgg+RUP8/ZwLIl/w4MaqI5oADqhLS6leS4FDdv40rAUM9sys3fOyjbAy5nR9
5oPV2by17YZpf7hvt5e+47eTEGBqoK2N8E8wzO+Wa6UlwuMRrOHERSaWVgLnshRf
PwmwaHWqtBRUaqMpmU3u92E65oG98C3cfmkFUESc28a6G9ybTeYy+MKqbWrIaDOZ
gOyATH0qlz0rGrE7PL5QZTK4ja9Tybd4ZOVxetJ51xNuPd8qtS/4kmhemaRY/VGL
BftlnmkmEPNe3uWCKPo7aHcl8E/zcgsidy0NkKmekWWHMYIsKvQ1Cxd/DU80KQhD
8EbGyqxa4VlJh8QyiKVUtDXiwC4ZcjUasH8JTY91bN0pWsboeomNFV2fSXoAIDrK
1UDNwhYelQbyJ61DZRm0b80mJIFRsSP0+3Tmzfge8JLWWmFfVdbQaeWlsxA0zezv
pY599Y8Q48jxRPlF/2zpd0uDuawEr5JjwBpw67dZWUUYqS/b1IcrVG1oM0zfiRR3
gKXDvidDFqTpsE/dBy2DhgaZD31qIhYKKFiUxpmedfnsFNzwhMQSOf95I+bh1Cxi
YyuymuOvPg+APXnG74Z/Zbq2k6fUJkOhfyohFW+0HZy/rU7LdGAXyhNrXj8sd7C+
tQqv8AOpuOVjVFDgtoakILa+fa6XN5Igewu+CYYgIkkeg/ShY2I/KfZUhoAA6dYJ
Ix08btk9ezQsve4SXc/+nyh+3AFN6riooWnQACRDHOc++hhzGFnT6oeA2N2oEZbR
p0831mMOcbqkZQpYJ2WYLBF8K5VZDvrHyLSwJBQTAlfE2xOuXwsDYW4eoaZwgVIx
o8/yb+Vj4gGjAn1GBwv67mCsAuRTimciZO4nAPpOW3PGMQsLuCQCF73puwdnDkSw
Fhqfwf767kg7LMWzgszYtjtGMbwKvFB6f0A6oCppZup8fY6du27IMIp21GwAShQd
zi16x18q4zAyzqA8nOYVTQn95mKBE0Q0W6IZgjtE0P5a3GPPueK6fi8OpXTNQj+q
pGHztl/BYdYjo4KfzWMTcZgvU2hfLu8ADIsuDIfgjEWfTurCpMgqyc8qJojPGbNP
izIN7lDphD1vedzI4WEalqntbeNkAzA/VbTyQf+K5jnDKHrkwpnDx5jAd05mkluG
jQUIeKEw23pW3RHIcsB87VR81spIRzo7PrNVkieC5D8istk4UItO8W2JTHB7Ncvx
U85YdKdonjyiZbBfRd9Rk8TwmBIzxUVIPb+aQtWIj6vUuTcCauYQYJeiJSSjmHS8
Ssxm1xZg0U5rH23y9mG72n+Fu/jbehusXHN5zlMXjd1VsMvzSxjdA/ZqMxi3sl+t
S492bYGnUnsOHL69+BPWGHc/VuJgfI+04Dc5OkvHcr80nHUpAjJohzw3pjg2qyn2
FI7SLADbRWTDVmcD+uzawSB9p/IpCtN1jz6KVDHndllbc11QJcx4TdI4ePQMZvae
ri17rwrvY0m7cXsHrNpeKc14JrRFQDVMPqPTu0yFpf17tauXy6qR8LAsmPF9EIfi
xB/GhGsMmNytm6SlEbzHzfMSyIedv5cxUvdtCqwFldHvnGrwwt5Q+nThguwbi9oz
gGqu75PGScH/Cx2KglFv+nm4G5hqff2BKFltEA+OtFqcO1V8TQFXamQWF2B/AHrL
1GhKXiJONMVCGcrjNqXWrQowvM8xH/LhlCmCHUtgC5ygYVoiI4g7luTQc7i7OISK
XW0b8dilBxSROkTD0opuR1xqn2sTsJODfQiGuDhJdN7a3NGr92Lr8eU9XhyR7qlA
aFzqCVzq7KbsorTakERDY5aYH/WxLKs16jgSP07Kmdk2N3dispIhgJ811q6m+SUC
e3yZKD7v58hZboeeOlBwslGQhAMEjPwuUDP7xXlZieJMAp12HLbpWuduLnwt5vTj
4iQ+Nm3cMxYIg82VftokStnXe22SkhDQ8dz0jDkGMvwgD7oUrD/pAaFGEsDyoKPu
86kcvg7VfC6VQlEWBAq7PAUEVVSEWao+8ClQ+RUYnXLYLcMNI+ZfLowWFN/V2+Y+
2FQsQntaNPnA40PMG20NgdNx1DhSLHFI/TXiyOePG7OxfKK9XWT3+9aORpBp7Vqn
xGAe9Zbs3RHHGhqnIIsiEwnhajbutQKYwC1z/zaPSHh1a6w1oiObCLaKcUFbFb4k
2dmcZQeL0W+YdUyu0hQ0bUbaD2JCYDYk2AQlcjlfzMrUp9SwQdljb3b2n9B0J70B
aQJIZpAfkTq4DvwRLHj7tJEpyzak3/bmoCP1j6viRSWbD4wDkjYaqNHhwAagsHZd
5hxDl9OMURnKePUphXOMCAnXr5Zf++7z3/0joNiDJCFpCoojn0w1iLhMvjFTaWX1
TN+6rbmOq+C/BajXSS9o8TC75ytWXr45hMXwEyT8e9Mlts7tbeSevJcg9GSelSpQ
0GPHKeOTbNWbd8/S9163wdiK6+ql2A+wI11LsmJM1LEh4kKp7CoroaU5cYsRlVA0
SpBb5HJk3G+ciM/bAsFS5ap5Bf3qu/C1vYdA2HYeMIXg+BFktUOBRH5oNepAwlTj
OFv3j7Im2L3FGgAeTEOJrs5hc3id5yJIBs/mlsIhi+7BMJBVxGB2eWQ36OFujz33
1Nza3VkLi4OJNdGzNvB4y2txOoHV+g9SqI20pzT+5BWSbAB1y40BbKVljh64FiiH
PxzPPhDaHqJU3bBrQotkL9Tq6aaY0z8JVJ+5ZCfKKuFS/oJ3JxP7hcPOyYsP2im/
yLirkvgr44HyM0I/e7gy2rOToRfGxnC2rxXiQ9mWBUTnqHzqR/0KYTwi6DRJCGSm
VhWUk08kv3VMYs2mwKShho+X9BHWMfiX/sVPprjHGnxXooVkJkQRa8Vw4BfVnGbB
00Paocbc4BWekWkzj95nIi4O/H1WfTJu5tqLxRIDOsCX264KV0hNXOagiqHBhT7M
yMhgkKhciqeTw+fGaiN85cTHTTrxGjTfPLURVeq0PRlSEQW2MuJFo4tOFNVQzSrU
za6jq0kYjeXxx/6TdL/kFZVkxlnbv5PxMaEPyKbR9JzrMjee/OgvdCDuNAjOG2TZ
MEFrHHsDG8E/wAI1jbKd/nvcQ3ogqM1cNWxNnYiRE5zibsOa7tJ4Cw8rxVx0jQIn
cC6dju5bWqY/lWA6Jmy8XJfBEq5Lp8L7u3gABMKsc92eph4Rsv7wAs7oqUEuYB7N
1Fo/7hprlgHBGgzI9nBA8bAgMZA9NIgZAm3+sXIXGy7HDhUc3x6UAyogFfhC8OpB
gU++DRwu10H6E/VZVgtrO/7IxfwvCjmckulbgZODdbrbl32hlnBP/13VpRtmb3r+
Lo45Wu36Hr3XVgVEI9zRJA/rutlHQzHIq49EXsklCgvXdDazTLlwIEiA46QnmYrq
yCyNaoNHatH/HPYpASX0PPEE0ilWVlCjb2X9eUSMxyNE1zuJMvjvLNl0ywzeCCyH
pyFsowLLKxMxJPJfNLiup04PHawUTXlQ6OUx8MJ1M3Mnq4c/zpV7gn7/AIDU6E0p
4WRcrfDTSsMthHFfrKpQcVYHdVR8a+/5rTWcXukNSYKk4e/I6otopU/JIvmuAMzL
te0VKjiwD48TsHbkycMYGAaPrXAOcw+clUssxnq7Y0sQFCRUZdbrzjUiJKrkM7RK
Wd99kNzgpwiSZNNjAv9a8mPCtleEh9AuEeRPa6iihSHQTjJzX87ZgFonApcl1nOF
Q1lHh5xtF/o1gH3iFmvt49f0MVwzniCdvNkCccngkS7q64fuW30WJJX9PVF9FAhp
mAu7g2U66DBkvy1Hlh2M7ha5xAtvokJXzKOHeho1SfxQXvSscwHkklCzD7JE3Xim
lmZjtFqj9QtU0m1bPOt2sNdNOmujjzanSorqIwfwiAdQ+mxbbOMoxg/yT5W1/mMd
PRUVsz2hxq3JuTcYj/Fua/2tGZthAUS4qx7UZcHYbzYDU4miVSllyoBdXfNNfttY
nbAUTF9qUVsAe9UOXRKRXkdWG4apg0iMWKnkOPWYUeGXafx+HPpXlFMSOQPxCqn8
UpgXLux7XL4Y95Ayj2Hb9iSbIqPFoYnQysru6AO5D0N/Ovx3xEmBqxc39Oc9dfqO
urU46z3ls12pnLQDu2IdgEOYASvvQj4oZ95/1HBjeTR76PEi9xuPbbB3i6xJE4+X
27HwLYaHGWJaqEFyIClt5aTJ6LMaidF/hxzMOq2FoLGST15lEAO22jRN+716TcwH
Ky06viDfEcudRgMkypSZUwT/6RCVeAGn37OL7cTE4l2x9GMS6+TYNMJ5TgnkWDdT
X8oK5dhVSjDe4XJrBGZwSxMZs3SSuuy6l1z3Vf42ZEt7TPJopvWYEfAihaC1IXmp
ud3LQ/eRQdNP0mTXxaOS0FZMSU2CTJQEFIXt+DyGis0QKTfLYEDKUwUz/g3dDLj5
Ej2BmxR5ChvDmkqrUkcU9DW9tIBfk+BnmTHD+nn+Bc55cQqNDIbIrBnMSPjMRMPh
nlkMBRdHiIGE+rRkdONTqlQbzRBekKcsZNSpdRPlrJeiqkZtbpwQkKEmGL89Vs5X
ZPT0H+/LazJQimvpZ88yEt/u0unxNag/Tf991MFo2Nz3C5zrFiIAwmSKIXvXu5MK
Tr72IB9JMPuJo9n+oop0SyO/VRfNGo5VAxWqkrttUJ7i3MXhb/fOMjCCw8tFdbUE
GDbOkZo+baLjdG3Pd6Bi1cZvRYFyaYMz7eboY1Q9EdTzHYDQDpiuEacMS7B/8Sj3
PUokjxcajDmNzuHHcg8RfuKAGKbORIDvfeKVZBUAEiU1lWFwz68QDETwHA/+qvWO
ZEV0Y5S6Vhsn61NTEcACKLrdNjkh7RmKcZavrUM9oP2ll4uU6Z8jk3RJY+c+YVmB
V2OYE5M6ypQhFbRRw86V8jYoFAq+NR2Lg/o1xx6hfb/SoMw0xM2O7DVws53POgp7
ecVQMAxCa0M8leEcaFIVK3KtP26J9xS9tfJPfdKy3R/gvQmX3c0P7ItcvIXIOmMV
ou1ZKm2ne8KUTawel56xafwuPV6lpxxDFhwg1QlZlivz6Dk0zJg1acrow38g4/3K
T010fBJGx7TKuElGliAIl3g6x/pr8OTRzu4jbNOHzPmaCNLRewB1zfZdRmGYXt/T
RzZF48hQygnqwrFho+9paV1PWwyrL1S5Guu8xsOGaAcHGLUTbE3TYMDS6WkTarkY
PYgEPIki9w36xuSjHbudMeNEY0lRtv5nDeoo7HSF+aqB8XWfXo08JmsqPIIC9XAk
uqT+ZO+ScN1nHxB6Rp5fuM+MprAAokwi0GQAI9MZX8L1cwffo2Cfj0OcFTGJX0Dv
EVNB4YEgThnYvH9sDWrgfP9CRjez4DYyrlqccNfYxtfFGBdZdnBbM5Ja0iGdS8Kb
zv+vBhExryQKVp8EfRiJUz0PP21SlkoLAu8Auc2Veu2SElx0raQwp/hTvtKZa7cO
SpkBTC3b3crMOAfPpnS0I5WjSA03QaMeVrJUzGgTvuapxas/AE/D+11apuADvmn4
gUXil2WngtB3v1M8bSMdUVkLVcRI6wzEHnWxl+WSnnTRuZXeY+5CVzThtPTMS6H9
EXu5CB/I7eVwdFQjAdClMd3rpCuyh/ZIfBjagDhddFSPzqY4mDQf66ZzOVnPkPme
qe00fO8hT3TDMBfhvWTfjgZK1/oVfVExYNtedoQsuKTL6kxMUYqyWe6gzziezpO+
7/+6Qaht/4jm4TfMU6x4RXOOnzA0t8SHQLjIkSDau5xyMvIPYp0gYDvFpXqPFAgU
6UPjd+Qx8rKM3d8uOj6kSVhgS0ffxHPzGuH8ngtLjTXFIUnAWMNhCkflfzSVnFK0
CkaJ6fm8imBu1LQfilzFI6m72FeU27rXXEptI9OciS8zSeAJsmm0risw/G93kDeZ
OKoLJmqnRQKEsevdW0gwPd8klLC1EyZxiRwI2qJ8fviFhHuXrxm55/hfK+VFrmcV
mcObsS3ZLCjHz1Sd9gsAnbxPidEy0POV22vmfi2pdXRDLnAWo4pPpmjya/srm1ah
MaW//+W9m891F7f+zermVmERGQtyu9sz/6NKlaP5XakFJib6Zl8TP/h/m5K1j5do
ei3hFrx3CRuO02hJcRtE0AplpO62nyObx1HuI4DwbYSP89kPPC5XM2aylgOs1F0M
PvxlSmX9vN9axplBx/8IhiE55awkv+1FcL2K4qFI7sLPQ1PqvI8db0eeAOJ7IlB9
/epVMLy4hMTEef6gbl02Gcujub4L9reOls9CAuNc+0gO0RgOcTxUTpZRdfGAo52a
53RYgfg2cQFac4LndGfE7uDgMd3vpF7Sz/LX3/w6d3fL0BijQNasC02IBmMnJZSS
B4bGpXfUdiOIkh9sTok0pbSVEK7tRTpfYOonrD/ikulZPVu6Qf1RFVI++ydkmzti
1AeI/ZTuRGBcZRMi/UKi7cyxv4XAEhn1E1Wm3CSdE6r+0AuZciEq9AYmuOJYXthn
giEX5Mr4gVNu2naM/ST7xvSvtAagEfT6RmxeDoUvw+xweqvOQ0ByfwyiXQM7lR3f
ys/jVxHIKNwNqD0wIgu/92Xvx6fR9ryPhOexTx28YHClJMyAIoOwW9rXal+lryZn
o5UBUzIB6Vo9bgoLhheLvOkM/Oy3jY+9TeUCfhRksYSzcJeNDfpdivOB6fUDFneN
niZio6k7pNfFNHJg+eBU+UUsu5NEjojHwDaitlhOnHUEarw2exjtWDO0ZRNbtziu
MgHh5zaL07HX0jaNZVf2yHOSgkmUWUmJ4mD9xwbjKFoZYoXfY82vMZEFgTMhPxm6
VAZfDQ6TNjM5LilGwU+L/RDRqk0sq+SOEVMUL/dY2rG2nTN6/igMrpUw/QVWjbZF
znZ2rDGoF3ZdAsA93YvNqCcJbEVRTlkpbBv5VCavBhijxaQ+bjSbonsqb7XrnS6B
CJFgWsHr5GFQn/qPgUQph6V5YNYghSKbbFU2ybYoY//uHlRB3so5t3H1D9vcj9Y3
4yEzPDWjJh7uIiU4gdVqz/GjKBc78+V9OcS6HxbOie9yrO57843pZ7ied6stn65A
vJ/37W4M5KkSnsL7Hvxm+eoicl7JbcA1TNPIrPymQAIDLZu49Wf71C9U1TE0lzk4
82lKW8tCG0g2MuPMqEhvuEQgzIsmkKZOwSq1mL6/zidQ7c6Uz7JpfBCXUV/W8Axs
38jMFZULImyxviNTajnM7Z4EnLeRlp59We3PojINF4zfWHSyv4oW/K0zGrats5nK
JBYSykqr6xctz4MKdDeZOdQmRmQSVI09U21UfGrE+5B9cPvc6UV9uA7JmgE+2vhe
XC/U2hQnJnLsOel0xAE8hFsGioJjNOSDDXrmq2tNPOVStMsFDYd+JXtwOx+Ado9W
Bpap2/tMunkYQKn3JLppv2DUCwS7OHAwEw8Gm05dg7WScsopZqcDfg4ITGjhHCSs
h7j5/CvAMK4Cp4lJgpkEFQjFpJDzYm4Uwv5eWuLOku2U7aWOWogpSjdIrvbMg+Ew
lLaab2uvv2ypGDXvnlOIGKhBxxjD9KdWydq43tPk8hUOkWNfU1T/L63G5adFM+S2
Leux/FSYMoHtwH/aJoK6e0KNR31QgcxHma/YNm7zdzXDAwVk0MnZmFqAXmVbBe1n
7qsAfmVewMBJ1PqG7wXpmY6bCdriAM88tpR9ohrc9ZjWL5O+SAWf0EmDXMcfxBpt
HggAnIq6A9SCcrfdHEuu0ObHPQ7lOy2/HFi4r2XHCaJpbw4fnNoP1mtRjEC4fsWn
JlTfAmuLYnqFwI1UIjGz3cXMz/Wuyb5RRyQV5LsAZtA2gCd7cdLxZWQDCVHVk/CC
sgp2ICcuXbqylVe3IQsESX93HE5IVQ6klCRo37O8XnUyoF8ONxj+Mq138Jqdd6Lp
vbymNVkMqN8BOPjwrXKnCZ5pxf6SuclwSswAG8NrabzQ1pw/zeyXJDK70vcuCR+s
045n8oelVdR1ptIc0U9wKzcb9KJNPYhis6unlU5wvV+GgUgg4Bi6epYBcCmGJzdo
jU9GiCjeaGjNxz6c9WsK6M84U8NuQxErFU9V6Phvf1mB4mXwNk/3tyqvf2o0T2ho
o2h7JmjC5J/4QC1MIq5IDOU7p+M/VrFJ2jlL7Tu3AVz8QUbajnOZLGis3WOqUJ4X
H/ZSP720UUcc/JU2iMqcYguJVWuQftRNiYK3AEIjttrvpSXND8d/bCDrU+d2mAHd
L6qSqg7ETuwahJPOA6Udtzo2UIouQ7FGj7/p9VGQK5z7FAWlbptlbMVD1iCIGBrn
9lTIBrSt/j2MW2A82doZkuWy9HO96TjVqEZ/OrmmYcZQaBUvqiuWI+1Fu3zgsKn2
kVFV1RCjTWvLWhNnPSFuddEMWu07YdfNTBDqTw8B+nqKTld5z0ts998VC/HPfDfr
lvz7xSEOzTQA/xKuDruoNQhTCY02N+ApYji9drqftVdhN5K44X15+K2lLrg2dxns
sMy44YQFaSROkNwoTnoy1y9v4DqQP45/nH23RQSjI5LWxygFlP7VdWZdbe6E6xTZ
/jhn3BtezdEz5c+/Yl0cS9qpKe6Q8fKq23T8WJtwfTM3k/U+oHoFBdUR5vzXL9hx
7bKaSaJndm5d3vKhUPOgrJ8vJqdbpvmbkXL+Ql4QpzrEbbKeAS/gWgvQTsVO3Ii0
YHaNeCRaCZPzJk72B5SHINbaoDvAUH6HAwkDKXg+YwPULzJf0lPG6vlkk5joGgz0
5vddxLVow9oEfGNtsXzdqfSV/1FoL3bpXyOLRDcVXwBROJRuPpCa9tEHZYIyGuIp
cTHHcSs7Ld3NZlwTRpQTccpgdHJMbvhyazUs5ZzYRYdkwWhKuJFvnAUJEHyd6Wsh
6T2k1fqwC9v82XMRnl22j0Do8a2SsAoSqsRzTfDpdO6v6X+TL2rF5ceO4WAHCDog
Eat3zUY+h3Ni5QFDQEJq99gOlOYqMbYurKSt6zK+WOmQWIfV9IvD0b1eHro809bN
EdVQ8xiwkc5v1huucs7BzxCY/w7gDGHI9nMCYkON8nWco/uCOZodbMaO6bqA+c7q
YxyEA7RTBVZEUIEOKMXcf33uhQGteF9hf9Ienboh5bD7vx90SvAJSbQqhigB4W2x
whb0L3EG3UuaDseNnPuLXPsZi/osv2DKTriuuPdAFw7ZZEGWMyleT6gfWA8YF49x
vCRZLe4SVLZdsbUT+ogOV3t9bcWHgIbhpcaMynddzlrHveKCx8tZBWgY6SYqBfZ4
z+xnG5XKR+tzbVo7HD6rkZcRKr22WZXDzLbrG7Yu0u/BSd0cGWNIz/A2JwS7HgCc
6Ut+jkuyMwtyNpguFPBrc5WHMnnJqR8XfFrAlAjcWOHR5cEJOWrwoWI36gPsIxQN
EY07ZZpD2zEQku1QOLgQ+wr/rqyihAxZJE4JsqjedP0TKOfpwoIF1K4cbRxZ3CuX
rqSCzma8XbH+kbPxHOQzveIl1dAPYv50Rtc5/zXQnBdou2o3rL0+FMbScMInYywK
LK3It8tMQe4raThmqQndLZcw8r7S7TLNqx7hp7iBVIG4KB4CSwfNMBqXqDj/p8ZD
11nZFU8HJb1/B2GlsKi1L3dq5bM+hHSEuD+T+NiqiSe/vuPRrQjrnQs4Ynv+aqdV
GxabYGTGDkPtMEFcFvUIc2H5g41TV6WZb+EcjcgB1t7pBijZGGlgewslMDQiEXsZ
VFT2YlA7ftNN9PVqRm4LS4+8CrSZOhEj1fxs+NMGZxCLl7eZto4TwLzb78vZHJWL
QZ2J0Twee3fgNfxI3v16PtUjgA/9afiVvjQc4rcvs98z5a48F8LOTNd+4bTgqHp1
KKAiIeD49e/ctSQN3cxWK7IpFOafbyHtvZ0QGHGeS/0jXu/Ay8SNVfFI5yFx+nAT
IVfNBWxjcSJkx6euyLQuQ73290F4Y/+d83xqb3CufLBZ/O9XpnlOfBSPQVX/+EEu
29pfum7V7yQYycv2VrUbKksbEQoU86G48V0JxxjJVieylCxSzDvlZ8tbm+P+MzBJ
17k0aWvi9B3moGwfJPRD9uQLsZ0Eru2c53kuGRKRjtH4Iq0BUyPuVTLE2ZLCrmZ+
bhBjJ8TyaETCxZuqtPNDN6jO5M7DFd5ju11qcZMw1hTiJFUhe8GJVqtUAqiDDFfv
9xjwjlq3jrF+yjyk+irQj5rYckjm2Eh8tBwz1BuKossJoKMh2vO4BUBqD9OSasMm
BtZ/mnm42jVbG9Ik9T5A9/v1rkj1u7/FQxVTpaVpwXzXXg8BXeO18RHSsPEP6P3s
baXbHfhgF1dPXhWwNpCIDXW0xiZgCasy9tN6stxBLfaMt4s7ej6enwJSDjqoDTZv
mL9drXCb4WjJwkbqnrOV90Q4HaaxNOCxWnUxgfmM3Qd4sexVCGsEw8iRVqJEknfy
PBwUvqjNWkg8kRN2/xPugz8UhqcHG0qEQL1wg/W2b4CEjXoHdPog9/xZi5zUGbMd
zTFVocMkwU3D4j1fKThfIWIJhBekLrynuEd7IPKK4GJqLX14iHRJwpICXaKvwLZQ
w3iy2u56NWYrx638Q2IP/LB4fLyF3vGRGScyNXa3nXqtNiiatka8DyNdK7n9HkaX
W76Ukj0MtuXH2HIT4hcrhwGBcyDUbxQSKR4Apaf29f7tomiZACOHj4pypdOFvtmw
+gWBW5EYx1qJHQE0wXELc0TxNGJUDVGLl7MG2R6IF0Db3RE4jCrtL4xLq65HXEZm
KYBAuZfcgsW0pK81s/S3sYWZxnl03C4Sa62SrjTL+6uW+Zg2suc0BTflAPfA/NGS
UajccuPoDLfjZfZVu9bAiGgz+TWBT89CfoyV7idT7eH7f67UAUkGbakf8TnKL6Rr
nf96WjW/Qn95fhXrM682+QLV1v42MgoHs9SgkqQ+leThoFAB2XCNS4m4S6ljgqTu
wWd6W+IRc5DItpuvW45E32fLo3W5+2grswYKR5GkX0PQZBswtpGeMtLgiP00tFak
0kS/TkjFR08nbqS0g7wSBN1K07WC6UPjOWAjXCYlUFcDGcwjTpewkCSAROwCzuO2
dUjJAe44ovquBB9VCcnLsVGQns0L+o5c3hc7hBU7FoJpaamYI+I4gf6DSLP1arXm
aUNKvjnptMHN2WPwYtzn2E/4U4aE/4BYK48MCXRtsMOKUSXK8FKoMaEZDblC2YSd
B+Evvq7DctgEFGjkzNG08HD5oBsrUG0rFawvVL9IXaA1JAFPVagYgOGgA0dhb3Ka
Rcg1LSGRuZr1ga/OVJYCR6rd4IlOvU/cz0btckxuRKryYLphl4J9r5KaEGtGF3vi
lzG1dyRzv2mDZp3uMNmAhYtfiSyjtUdAKQS+fHfHVNTzDAyV52tWc2mDP4NGgcib
jkvzcSKXX1NRcEu937hu1UkwuU4/xG00lIt2BGpGATsX6AUGaSthpCK0fjepFO7m
/FARrPjVoE3paMTm0G1diQdsijiHglHG8u1y+12Ba7v3+y/Uu7eBfiWy6MA9YhWl
5eH7vsXNtzDN2iS7gTgjz/OdiW+X9jPxEAdbUD99Q+JNh5GC0bGkSmlPH+eMru7g
rjG4Ck7q1n0gBGTyeJL0OCqyT7gMnlC3V2VKWFhMUYRJXIemtuYzvP1R9DVKFJP9
an/Zoe7v7Ybb6Y3qaxoS3s+LrAvQfeAvZXv55Tt/GIIzCfsBja2Kk0W7C7xueiei
KYnTtlYB16mOF8lL7qbxNzshsRkn3OaYadbRQoEKzuSgXCFR/2y+hT5JR6XEyMB9
/VqGbSfjbgv20NAdhzOpccBa1Vw2xlxEmXWaRGt8Z7u3XT0TPPZ++7xQ4vebBqPZ
2NtcnFuugyXSvj0IQfg7P85zIspWDrFiKmymqfPqIB7EzUQnQqVycpS/KxmSAMJf
QwXdzuBPNXe4uW27Sv13qo0WxeQzYWMLZAJoCJ5fEWO+0yLn4cURD315hMa0s9K1
uv9MdwRUFtjsL4W3KMhI5ge6Pm7C9gTJtD4NjbApH9dG2HBuunsj6K16bSkh1895
wd7tyGuw8AdV81AoPTNOf8fRNG6RImIZr3G83X8El/cK6HMB4Lf6LqJBtrsQo54A
RdLDLuacx/qEKjMY3KDD0r4aOc4i4VuOS5A23K/3EwPUcIkU6KPNcUYq5Y3BwD6F
SeaXzBx/82/yVD43HjoRCmrM771h0pHVFiBb8uxIFLNsFyJZz3i3BbheCZ063GwZ
eK+5b97E+imQJVNSZyJL+RmLT0lnEYIRAM/BbqzBFSVw3zcdQywIRXewg5skkYzA
yHNhD9E6jE9vEvw7L3YYcX/D0XL9496tdirhJamrOrsrHRCQMt29yLpyQtQaCP5E
cRzX/X0WhXFiWQ1T8UqukeKeC6HoCMrBgedQH1aPtEmmRotbfj6TdwVpERkrSyzq
cDdyJPFTtIuXF/FtEYE14DTO/VUGcKjNXcb0CLLe0zQku1rwTt6qcOocMYKBt/mN
2av48xQdqS2sYoiVdJRiZ+eg0k/49jfs2qsKY6XAWGeGae10E6YphyAoKltwMaLT
N1ti4/NZA/M7qIT27fEao+PD9D9ZeOFZfIXKoqHIOfaC5ll0QRhLIDO5HXKT+6ve
9iGIX+hEVyS2Ft9fqxK5y41TockrKl5zWS99IFcgkuOoSF+0wxqYgHFFqmzdXw/F
jM6X2iotgJAiTIBWgZOIKdeko6kFQH1NAGWtjP9ldzwUMr3A4/UA5LHWcSGJBOhx
iXy6tyGaElwrZblB8PR+P9WiUuDghryFA9JOaexyPUJGGyKQ70d5LCLmZlzZ+0GV
4V3BtmTiNp3X36ikk9WNarC/ky8iQdfiGligKT0uw1CKpzu7VfLPBRT7R7t4tEjX
rnd/2TO0NIyqykHzJB5fQZXBxKe4MRlyvJ8a5wNirHauqL4rDSNGTgzXZ0NDasr6
oa2D2hY5DE/VYzUt9BAymRnb+jaVP7D4ZDpjrVHSvPhpXAALlEtIVHhDya0UbJXB
FcQ0aYoTY71WQHrmF1/xrOrESSG8UxUbjMRraJAo8W0wKfqSQU5GHe/ztN1A4Wms
P7B746NJ/aL7aRAAJiAAbl5h3RZJXxhY30rYCQTL++zn29EhBccXLNYi85q4j9xe
SrogTgZY9+CNxKSN8yGKOPRwB3r/lSMEBAYV3hGSBCdDGnxgxaRcArvNXb9/CjyB
0eNvuqucSQk6ykRANaoc1hgs26w1JFF9LyYLaRSB0WYTMGSLoWYLPz12nJk8C/PC
M6hwAWzLoPkR3QwJSgNR49aP5oBNSpV5M1aKe9MC77KWSgSV5WAi6zgGcJv+89J8
CLmajZ67flJWHTLsf1HMBVYoho8+bDjGwpbEeAmBOTWq2/QQY5tzQm8xxLP1oApk
SuEiZNnBpsdMkEepg8NxNdOTnLxDzi4XEHAKUNjFswvwBVv1MYIa1WvUU52r/UQV
V4nRqWog1wQH1sO1/A8HHX+jci8kYcyDgO4t3EX+qysLzcCwECjN33oEtsBBe8iO
86g8VF0p8L605GU/6Xx2+cvQh9u6bmKkl83lfO95hl9KYjfiTacXgL2g6c1bSD9g
p4aZ11ccD8sstLRnnM6S5XmDYV4ox16dIMa5DWoQyx3FXMi2JTrSqplNuwGZCMPf
RZa6An+cEA6C8hDKbR79eIL2ykp00MXexbBNqf8dRYD2ADDUVyJtbV4fvrjwc2pD
cXXKXh1qMHKMjGdgSNmWuc2aP8C0zSh/hNeVnJH9c3nnEafG/tL/79V5O5KSmLyE
PEMtqFBE2Opq3BYh0qJqn8PJYy/1DaLUxBtgFZJNox+iTBWu43mR8gLWtFEX+1aM
+LbpaozAGt08vD2+kGlMlOEAxJGLgKWXrLnQFDT2qKX1OjsgKLAV4md5osDG4cZZ
poAVJWruNCfG9MxJC5QzucB08JaiKaHPyP7o3fFHGFFvoXXUMwgvlvzI5wrNQGwG
/8sZAS1TCgLbDFdT+2f16r8PQ1SdJ+xH3qXMV8cSzDEGAElKll8Ry/m2u1/pfJm+
Xh6ZQkCjExjkntGN46/vn2BYF55J1VA/q+oUOifLGUvfv82UILF1wkcUD+VE/jg2
W4j2hGPMow+bWddr58Gnz5bpOvnoNxScH8YQivbY1yaIpKg5923lqflBYUep8LFG
wlh7Q1Z9H7yof4V/lA6P5pzfLY6ZYYpQ/ATHHQ+Bx5FNTJrAU9km+IgBpcGOsRiS
E/zvelt+qjzwK/ogsJm9HBeAeFS0tinXZv8P1bZysf8xaJHsubbRriRgBuExPbPR
qDWczdjb87c0VAuJG58n9x7jycDKi19tmB2E08KypkAUHdGB+9iumUGykMOKRZYy
ytcwpMN1QOKGniiH69lAX59kRdirok6wiIjCmjYW8GEy4hj7TLb8tD1PhTR6EUj6
8ItoH8ZVukHU5GYJQWlvfxtLr8F11ISpTwW/5E1kGLoFbEXw3KAyhEAuspk3GDLO
51T6d9HPVIG6Jw5TNnYORvZo18XukdgtUjoWJVkybR4qjI+NGVXK5wB+w/d15oMQ
K5vVAqBvLy2Mti7RmIaGUeEeS2F96WmEtMPCbaGG3i9e8YeGxuznvmDBpWxfK+I1
Jb7jYVQpEWqbyg/zCLA2ULm7Vit3LqvAJHWxASxo9BC1pzyIu/JdsD+ijYfwQWT5
jRi0qPgcPPY1zcMrNXoBCbMcKD7aX+IJAj0g+Lb4wcUgYBGxlQxM3IkqdEb43Vld
lFPLAIQuZgraGuFS+d2lSkTJgVkduij3RddY2ZHJ/nll9AuHCXeeLBcy3b6hA6TU
OR5KDyFMyFEM4bO8BDWZ77Vw4Mt6K7gvapq37Y7AKAPMNbfuLH8kyyCNjIiOBUe/
xMoaexD8FN+Cfr4joarPNamlxuMjplL7EhrqWtxUVxLqJnwX7IHvjRt8VrQg69oz
z2bK6+uIzs5HcR2xraW6GRiGu8t1O5chWonkjSDg0WfJSnosJ2YCvKnGrkATjql1
OWxgfQ79qJ/w/cFr2uCx8DGMfIeFcgwrhqyWhn3I2vMl+JsbkkXzmWGXFwhxFv0F
23MucdfT4SK4YBZbVRcdlz80UBPV6p9vQABOHIPoItpH9hxtb3Nr72yFPM4zFhon
NlVf8UI3gSzK7pIX/EGopzhmaK/d80/xsNAAkcwLWahooUAwpZUDBps+0q7NCk0g
OfFnO1zrOdChuuueUdilvFr/3Dk3V1/4hv7VisOolgSNlxBdlVTQkSyyiEEutMfn
qp1Gzp4iyaUUEZOOurWexSrCC/1lnQ/0RdfLmmy0JBg3HQX0kHunkFzquP2mt7pj
jjkHcByeGfE3J+pfXLmLUcJ2Tny0fD4pxWRwkAwNPOemFqpaWRv8qqYTMvJnWDco
NBlkF3nRZj2AuvquRKVEHjnos48Di3QTNYf0T6Ym8rug5clFuEMLfD/484KFByCK
oMIXxX/Q+8SisXCRbLmO9WbTu9h5B5lYAVOH6uLZANMU3YMgqbhB+HYlxUubhsqJ
QBqz18iqBZ26W9jUFMQO9qobDjMikpCoHsUoFkRQxa56HiLoONmLAcfASkGpyqGk
vrI0oDU0SpEFk1LWqxU4ISRQyk2mNWYSg8C905uORAWuqxGAkmIcCTaL6DXrAJ6h
gsi3OJE4OLnMf7M7YaRXTGi5ppGsJnWTpF91if//4Yrek0oNq0RN00A5wMJXk4TA
Ik6XYWoLegM8qiEUIX/9JbKyea3QEB38coh4/ttPqKJXPuop3Maqsj0PkzFxAz9U
JVx7vh7jpQ6+je/dS7aP1RPiWp5ZCDxK6RN4AUbQSOsfWskI6Jl35FINe/hKbrjc
z+4ZG6dl+0dFlHkgfzH+u/pp8uiqsW4xX4ctYW7elvCp+/zQgf1j0hVR/zutUnBz
7zF9KThXB7ZAIzTV3WBoHwKAUcNrU24n0keVH6Z89fxwvTdLvwoBL7zs5/E8/A9Z
uYtnEoLzSs/c6AleS+GUxk0EbrBTIvfCV26JyKaZgo4U7zIrIgejcpXvMucBReOQ
amooCAfghC0aqvL4q37gJypeo0bKz/Qo99h1SSYsV4eqedNxzIy/ubtD4c2jjC09
43SweThmlbLWjGqIWTePdxjhcV5SbJZIu5xYGO0o0zbZimdE+ummHQONTBzLNi9M
xf4SCxNnVm9dOjyKj6GzKJIU9M/6btZnem2Jmq17a6nqUxJr306mjFFF3GHLhUeD
+q0y4Pv/J3JXunmmYrTRnvH1wfcSoeQFQ4Giv8F7jKFFiKT3zKn7RKZlJp+HBRiV
9nsNeW4KdVZdE89Rq6U/zdVYIM6nrHIUcpWYui7RkvyY6qw9oF8OmC/p3lTg6fBX
6VcWlGUJt8fd1g+WEFNvHP4g46HQZB6wetDYrFJSKhwJ/Fq4fICLdeTvLk1A1cVI
QIsxQ3qgR0iH2O6ohm9tfcldc4mJl02U6rY1LMFKQsQftrHzNvSi7HZiBlXu8tPK
B/sSP9++5Tp9Fkf7flpfYotXcicmKQLRSIw8+ilFtdH5Z++TxNN9xh1dk2ho+qkC
iDHP0cKp/f4qLC2S20uSI7v1j0cUfsGwa+qhgx+sIQvt09xTtXAfzOM5v8XdNqcj
MDt/tEGuHo0gaK120+Nh+DdslfpZrw5gOrakCkbfWrsYvB6fUMu7EILTZKNyja8j
1DwdllEqb1vnrfL+w+ncLmrgYlbXpiohhCs1LoQRyvlIAWdKEgHSgGES9yW2OCdK
Egab2fB4+vkq9pRWSIkqjA9yk0FjQ/jj3gi57N9iVLirbw6bElMRs+Zl90YD+XoB
iV7QOe8JuaXcI/8c016hg3nRnu2UQCmpyKS+0wLMXhrNj7Raoe0I+EEdKaRaW972
hboTbUG3pexCEWBjLKn5KLrrvQXIMxOHKqckn4Fq8aBBMfr8TwhR6KfPFWO74daV
/M9OafXxYAtEHOP6lViPhFnZ83PvCBUdxxq+O5wknEt3AUZPvcjsvhS9pxPIda57
OjfO52RbswN9wEqmRorUA3Vg9/BCblZcm+wQ0ckpN5pvxsltrN5Y29SqIUhrFmyj
a0UgiDKqc0Fg/W+gDxEJr+K5ZrOz/2QOwi9mHCK+F8WBbUkkUHQG5ANeBarDbQ1m
E1A0ns+m1S1EX9jeq31JkPeiEhHgk/MiiX0/V+oEgJinCznRHXlMRb+ksaZb/c0f
lXC6OqHXH/b8stZeK1RmaHdAlwsNuT2NnzT475VFuZN7z3p7UVBrO+Xfiie7Wc00
NrX6MG4MwQsCywYa5E7oxYA6wnn59g+6apyb5QflzNfN93S2L/ftdhjPBf4673Jj
Y9FuUky4RiYARcbJgEOn9+vGRBEngt3b4CTmZqqe3+DQ+GrR+P3INV3Mh4xNhdoN
+Jnkwja5YFn8s06abLju3SAd+znIMlmZcjEG0Py6SslEpLD29UoD6lmy/ZqUKSM8
RYPdWsEyQLEd/UrisvH4xiiOq6841ul/yEd/2oZnFvzl9nS9C1YBVbVfLp46vwFE
p2DLnksePbuVHIIXui09FuJ83pbRwr2R1lYksp/J7IXz9vEF2GG3Fm3ROFTFPnKR
yqmi9qWfZQk2fe8nzgTqDqbeN0uGKDexDupMepl93rEupxqqoDZytU77x39vN5JQ
UqsVSP8+P4V2h7qHW4B5cox/H4JHfk9RqobmHTB4OFqjZwcBF5V/nv3JlrDf/0tu
ZjiHBK/nG20Ic4CxjeeXZwa/UvJan3AI9h3ZLbu36PUKYZEQAmEBFt843JVHK4lT
y6p3S2Eimrc3DF/Y+UiWbJOmAZqYbBXAnuMQndmu62a1jRjeP+SzFqwsNbnfov/o
BS+PhhySf+fGGoOJEnodzK+XRmnxj5+0jBOstiJNVoPUlY8IauY4UVLUloERBAD2
Xx7fbibr9RxMAELEiAM2mA1cSU9TfKl+Q0zEI+pgK7ut0hVLrfsS3l6x8AjoH3eq
ABztNFS2XkmJFEgzl29wA9hT4y84Rn0cKnaE8Pc5WJWs65trWGvnwKOn9txF40bw
GT8KVsq/GLeCo+DeXALLSy1hCBgRB98RMHjRNyDyuqTLWw7gxeTmC1BOXy2UHi+4
TlxzZnwJgCvpHwQQA4csbbLKXZqh1aunBnY5bIjxapRjn6IGuZqysB4EGbweS+cX
6cS0Y2kdmCQN/jCUsnmemnEptaS0ePmktM3IcX6mvfZ0oEgYPzHx3KDKLjcV6Qfn
aymNzDk8TpZwwA41DvTEg3vsAq+7VIxm0Z1EKZdRCPa61yhaI0MmfzYsd0efF7JL
wVroH+LsNr8CsMx5Y8o2hDw29h5PUITyWeNrL2uri55U8GQiTgaI1VQ0UzTmjbwT
oxuAHRsc0Ig5f/gKIOI2fUCdYSHAa54Zr/JEd012n26jVgQucrF62Ie+H9TPeSic
J3kPQ9hm1pIWOo3EG5q78oZ4jybpVMZWi/owhp7gaxiSgnXADSlWbdu6QwhUSSbw
G2EoSzLiSxFNVYCd+ZZbSRl0tKd8I5Gm4mnntX+PDL5RR5lEFZKisl8t5xQ4vAF+
rctKCkzsuK+QlsnbIzIQC6EGcQ2jol79aVCWkXRyP4nj03mX9GbZjzSel8/zbu5G
XBKFGqAdRSrILpI1hmRkNP4Duk3uR5hcIMqvELUkCG20IqLlFiPPOvpp7Selkxd0
b+6Ge7WGyPsZFUO4YU2BkZuBsONmGtepBSdVpUg4hXkI9NZ3Qm+O8UrQj+IAm7J2
Hw1A/SFpf0RVZ6jtsR+kjJmgOsLFUT48DCumpg+mk2kxj4eRef00pwMNqADUrLJ6
M5s0LRZv/lgYC7IxOJPnlu5A3M5exZIhhWuPmIwHPVQ1U3rOhy2IM1TmOLEviKM0
FZ5OlgLAGsEg+oP7GCTDJgC0nbAqqUyNtvPBjuLWvFLv+r1rCXi8lG2ZrxOcMs49
b4XgKeRFCQfuwWL31lUwDdafzR6HLWV+Q69UINTCu2MbZV0LjyfQvUNdZBL/7N2u
16+7V4kVGQpIjOrD92hgaJn4qJRBHHyz9i2/XMPnbAZWHirne8a9RZRTxZJtlbfg
tTdM1kLLAHxWRgwKXO2t5qtwm8E+1Ug11d0jQXpvriCMDVzCmuYSfBmZC44mxKG7
7TAmK0uEJ3gO+7qmLEhE0gA1ejrb5t4P1CA9ODaXMQJF35epAN9qv34cuf3hPmmu
zbZ/E1ETNgCDOfoAO7dZlv8lLwofkXj9ukWbEN8KHVf3O6B/EVMB6JC2LTeZgYpv
2PstuP6Gp7hMGAxNJigUOxkLFxcU6h0DXTPm1mnpPFyxng4/DWgYd3dUvNUbaOhj
ffV/UfPoN7EDXCPkqMU9CyXxhnJFupAui7s3e9PsJ3Y88eM4ZKRJPiqSB8UBMc3J
U71mkLdLCWM8qWfqYpew3J2xoX7iH6DZD9ZtjA04BKUHnEapYBwi+y7eD5Jf7rdm
ibEc91smUilrz5oUVtwjR2wJdyE9DoStjLXONHIfTWEiCXMNtz/mC2D3IJ2dL5hb
JJ9NYTeQn2UYHjNI6SLMcD9Zkx/5kMcmUhhBhqwKdAwwlqsbO4NnOq/KBlSvaY7Y
2825ps+oPnNm3qQ9+Gt4r6bYQhEXKNqf8sR1CBNCQ+g5eZd2VwQALn1WuYVvQv8Z
gfdPw1mxWIL9vzUw+ldfee5/tTss4HZPyXXI2Nx+HY0gnANQTfX17dPBsdKHnDzM
dDH7vKBuGNNH/yZT2qida5LX1Z4bqGUg6w4P3GsUP5LC0ibFziUETgY0wtnu09uk
qX9mdpimTzx1YZEhzGP3cG+lR2IWEn2AbLEgivdbgO+cibQ1pX+etizPN2wfkH1U
w6GYZ0sbXANmufdIvb8wqLmYCbitwBI6/job2D5zOUjJQaesk3IiVzlpNyUggQND
5EbHYWgpCpRqr3CiYHY0o6zdQrHT3U/Bqc34Apf1GGmmv0nYpiG7TkNll10rOIAa
9bxMc+pb3OYkPxio7GsJSumCmtEXFIzGfUvM5q6jCCj9zSKYNr5Vlzr2A5ANVByH
6eF2QuBbYbYhJJhbnGorrRUqaCpfQeiBCHjUlzX74OLA2EsRy2SlXgKatppvKSPw
iuck017YXewek1xTLeqUIKv6U9GnUVfuFDDIrhagOe1219kjtU2sJ+jqwzldlPI5
NyZAnhLquzOJGxDwTbZuNlF6UndtM7fVX2j3aa99Crq+g/vSlz9RN3MXimLPgXXv
0nXNRmq5b1VdYHU4zrQMf2zNX50TlAvtyhNJfb3fNZJrpT8ZTH8+dT7ULdbdfVXP
oLiWAbbPWFuwWBMMOYPF4MzfavJJDc4czMcrciumMF1ywl4x3KWjhWRKPCo6761p
CPRZRnHrJ7vv3A0OKCq59lvHqg3ZDHT/XuVVlJ1aTeLjBDV0Qh1abGYUTSZZO3QX
5UWNfBVosPNX3kmhokaAv6I8vZFcJSacolsEQbwmjzujNjuYtF2o7BcEWS4cz6TC
I7bCD1VtEEEmIT91h2PUx8SoRnPCLbtlWR1Pna4eC/tJckbbYjELOIosUH1CY6ws
zHUAYPZtqjWIw/C6h121R8xDjpy1loQisKdic+drRXX/oK5dUyrsA8SWjkuMHASq
selJEpSwwlOuqmWbG3/YIjzx81pnoC/iqXCwmGFJ5C6iSijEcahrX/lFCtW8wSwz
fDRUdGC0lTj+frNDZGu6pqpUe2AT/9a/dy/jL14FbKwWA77EyFX3fDKweeGs+K9Q
U2lmxIRgTQP+Cmfi5J1yIy0DjKizQ6+V6KhXg+1lQYcz++U+bHOmhYXclwqrEyiV
EWe45GBs9vckez3wgEEgXOJoWcze5WEOGUHBRw/wZHPmmPSvHvBCABOQX9HmKukK
QyoUX+LHHxSyXmbqv7FPKW+dh4XJHFapUR7Ioc0l3S7qtyUmQJ9mLV0bmLpo6hYm
XkaTxYMBRO/CC7v4z+7C4+3TOPOaBxDkgEJ82TSsC8TNRDQFXCNHkvMb6EbN4UW8
XSkMv9GLONwJjvankEWVZDPR97UmIWF+FauITBJRJomLitH5yC6aRFQqKAJ+per0
sB+ESynyfMl8YjHVCzoMW/76pJunMkRWE10E7fjbWMABsf5wmE+VEG+RyLjqJ9/e
temamYiToQ0d0CzSaFiRR/eOMipAy1ElNWo8rJeJ/iNkVvv5NVIQbX1CKwLqlCkA
bk9FW/4UoNnYX0x9LCaUTGFfufr0CaCH4+lLohJio/7XrggLZajA59yGyUDWt7EL
UU8w1ZRxFTUyJ4SbRclEThbDMLUC81JNWeD34t565A5TXLMKyCSnLmy3ef9kO3la
np8Ku3GJy2BpPRMyVnqpoOugqgUDSwR77c2j6ANyB/pnQBWJGv3uD5XwL+fBvp7o
8WGcM2+lUkdjK62ePFsa/tZoJf1aDIUC/QrtcHSbQsbsjDDBUgGjnXTf5EYW+gEF
QfSLmplYpxh/ngDTUgC/mLsGM1iSbOHf7T1QmuqO7YsWvGp4sHHYtfHwjYrSV3cI
lc05upX6pE6O+wJyOj1ei4LIFnLw/yJ/1dbsdvdDS/VCNdnkqi5Upni6iPfJFiZv
hAytXRS6Eupsjiwz3UG9wIUY5uWT+TtfmporitFVGipSPD3LS1bu2VDxpYsiApfl
POAm+uRXDk3OvUxISTEtBeOxKj/9ZTYRy/+nUuqCHTg7GBDG9PXDss185U3WzCj8
QFJcH8wamVXScJyXZ1yLe+AZM44A5VV52AchZy6bPoN+bbp6OJLJaUqqcdNCFxAW
1H+dVY/TtZHb2Ftq1cLyrVfKaHHKWkOE1h5af6Ms2yRGXkzpMdBM3+GGWFmmKalv
2/U1pEMfTt0SdVaMLJ6+ZgsEdlvB4MKRoTKGHj7SVHCUwKZbSqkOEoZWw9YfSjej
wIDa5i0P0yFc4td45KpjFf5LJ4JFeXZgbYdaKkLYdzPS2q0vOHSqcskhBq5zwXTH
dJ2rn5JpCcvjwnQMcc+WK7OR7lzRj/xQVlRX+I+VNjZeRDi8B7LXiz8mPxaPoErn
6TMDsZ1r8ybtEdggCPSdzH/ay1s7g9dNZwg08/d77uBRjEwzFkQdpb/nDmblctbI
/Dyqgvyh/Vzj1qspceMQZeVkzYlej6LMrsggLGLWRaEzTj+8eUExcdy2tfswicCN
CGZfR+M2/xKlA2g3s2+/54oEjwNOVbHQV5IZQYvKrOQRVwcSm00DF5BFI72VUYoi
pW89pcNDrZJ99LwurnG+p3oydJuDripqtNzJSWYRpAhMh3omQofOZctkY6qJJavG
wI9cqfDPdvoSxj2zwxyQvrxECVro2gtBCHcDIbt0llVlk0I8eTsLl+vlQ4v8RrZw
g9b87rsFt5OBJp4wqqEbUNgyz3SaiP6dPemQXvNiTgQ/grKBcW5rZIsmGmDn+Oc2
baqIL19povEfRmYluwAJNpvtDT2mUnm8cksL2i4Tsia9qLLGiTMcNcrcgwWDjcto
wg12TNJa92m0lTHrC4w2V2lVHtnCR3R0ssFLDFHS+Yca2A0/SL1lLF13+yBKhtSm
mN2r4aokwiIJ4XnxiBMdWIz+iWRWXl+9gdVYXn8S5Nn/8H6tIObvtGihgOaJcyRU
c9iDMtSMK5idxMWjYxfPNcByd/p5Ro8DHLZVfikL5wzL06ZXaQKSsFLCDAE5sATQ
KCKH2/zJq+eB1TgXS6/jL7osRITjbe+XzXmbgDG2QwPdnMnEWO1bNuBN2KMK1x8r
5gPjM1sjIqtuJS+gVnpPKbYUF6cTyM4Xf8SnppoN3KY8mndOruqNI3UUVcF5piFA
kDvaMPPrUVMfQ8UAtXxk+/+ke15hlq+zih+dIq6p3RxVoDb1KYe43cX0Qkc6ZNGz
ziEWZW50xw/5NQsSeTlnK97JIRWnuraCoOHD9vcziyPJAoWdoJoUsC8dvzi1/vEo
s5XEO6JW6dufrwlYmcptkcnuuYUIWwNO7o4E/LmdQugnyvmg37ipgkSKqn/dBVgo
XkeU2jkAxfJuzPX5VzVHqyzAq7ZoZUIjLXdCyDbzh2+59Mp4GduJ3YbaZPL/LZT/
YUuX7CMODzWCf6ijSbXmdq+z0el3/JlYgSstNjMqZ1nvJaswajpjLbAvG40qnlBO
V/izn/Chnt7Vpjduqkgb5gT3nBAPAKyJ2WhHPz3c7Jm5KF/MzFlWH/X9jNsYmlwq
Mtcd1B2zayaHOAQNk0SWwE2svtt8K1BcTRlvlVQjNjC84dnIYr0IZuwWGGz+13cY
Q8LGHhqtVFeDRRgBCN0w90sLdrKG00x3B3YEdxkjcVBFiwgciPEjvtbUi9+8qp8I
OyZTTUS439e5xbBGap6XDgy46dUXntNqmt6KbgVOmdlMf8JshglXmyu8nNKoOwNQ
brN4yXWSQr+drOKs1o/SgWbpWsNhXEmDAUA1vtynwkLAdg6BNDLI8mB/HSoAtypP
8qA4hccmWqtiOrWZBOgARgsQFp3unkqRgrVaRb3uG8FQ30sXqTXT7BZtnYzcotya
qqtEYPzkh+ttr/wgPZAsZVgqGEg0Sc9q2kMsgAh6Bea7LF8ge935cGjput71ug8z
tOeQBWBiiAJ5Udtb0GUna16aPOhP2mslWArZLRql+45R3qgwmBWeRvJzxJknW0ci
HG2ltAhwUMQ/LnfyBbyi6Ls8jWWr8CAw8M0/OUIzBLEFmD7YwIbVEpPCmbseFXOY
4qZTbQf5Anck7h06IkDwwhwpuOJfryO9sMHQj/2sKEFh1oXldpSl1ET48rL8sVpp
87bQYc8mY7zi3u3n8TKTfX+L3AjvjJJGqthkab7Snl2w6OhPmUZcOTnKav5LGQLt
e0yvOjVC6qy6sYuXL58Wxz6fY349okADYCiptJs0ONPx4bxAgRNAyhKcrV7mpTmM
cVqqXHWyL546OYZs1OisO/3wSQazdrRcJ8uHJmuhyJ3epJkGyxdwKCTmxIvt5O35
ca4LbtQ9B4X1lbjRmbKDnTDXkOnmAwEf97WkG7fPNeHePBUU2iRxJV7ZeVLJQswU
Bq21QBOBhq1HF1JYxM6YDCPJdyfweaU8aVHR8Mv7ES0CnNXhxgKafrRahAR/kqhX
9QVT0JI6J/351t4KY67SWW0pDat0buWd8z8OKNZ0Vk95CRNV55LZl4jcE63IIag0
lPwHgBn041JuU7TV8+MgcOOLEy9J3UUhLDopBzH4VIa15e4ZnqJz7zka8DVGQmqr
1E3YPjgfgyKqA4RMqsCcfqRKgYC+vVuQa83gJyBfQuVV7HHE65shFTHIAyAlUtXE
PLmR5nZMpgRr+0jNCqxIZFbnKGnibdKqaUVJrFOaXVOw6VScpqVNSU0rVKkzEA6i
LGg/R8MyB+xlvO+YxFIwKxblEtLZF4oNsvMiXpmhugZqaCDr+ASGW35nmlom6aHo
5GI/r/G74o6df/Lh2igKjgoAFN1dMC16UfTtD9a5Bz9OvFSKMZViHfh7jjdesSXW
Ceh9BfX6CMjdQybFT2xui8oDrxBz7HZF/5kq+qAEcH1vsXSV17v7Rq8Zzng0tieD
CR8QKd1nLR8FO6gh2Nym619HdUT0KIg2g+z/PtN475aoVDeoOhEmiGtwO5bVjk09
dX9Yr1zqfkcznWttCOD8Eg9sW7bAod7VRgcavHmNRFAnHBtD1gIHpPMBLySFCrnf
4VxxJLVi0JURJsv0EVuf6KTKRerrw1FtvqiFyYCDX6kHaUH7DQdPqo/4WVnYOD2N
p1uTmNiTSk3Vls+NsfRCmcLnERO/eyltOHiNYu81WZn37u58MwhSiEmKcan1II/Q
3TbnqDIc/YgOReMV1SKOn706XBGaRcbJrU2MJJgLyMCNd5g6NTzJsfopjCE8an71
W9lJ9ALYILNApUxuM33SA3YdbMtko3zpDm+Hkv89pgCzPvP1YUFXWDwatnO99KeO
1F91/jemO2UGiwEc4pbbWzHYMXtYUk2myLz9knAgCixHNUp92wOV3FW44dOCzFT4
44Rumk4Z+q27Ia94lM6MAItI/oQCpJ0m5pNOZil7hdTjFEjzkO22zOCg3tF8U2I3
D3aJgUbX55ij1g1j5mx/HilohZmEEkYIaVD2Aj2t6Kj49KrM9amLZXXW9Hc+YD6C
kdWHdAdAqxvm7G7lKig852abOcPmz3ow4+wSu+8G2Xe/sjf9hFyT7hjTIdjN8kNQ
NGr4zvNbLq98Y2S3+gDLbhdiZfANHE/dTTNCOecG3fVm3HWbNVHAbTsUqCtOSspF
s27VNqfRBkGUjwzuveg9FNMLw0kHpmqIuWttRd8LWw/8/cZlJwB35hSGjeM+odkj
yi3J8NoplzPiISLHivpATFhPnJhO9m/jOl/vPRZxLlT7v3/1tORNxqnV6UYkYp7c
2LJcuT9LEMtrpLqdfSGWFs53TU/tG1TUqOHie3AMtl3RI2lFyvFxyCnwY/iX3XKs
9bq2YaWctThRRgzhyooMidbkqXn8K8Ln9bEEHg4OiX9CmUWNv+gfXITNCYzchwda
r4bfcs5o28pamNiWVOEQjwJ6VEfiofUF2wxu/y8mKCULCSf/RYUd9nUPHWTfOgyY
wJaQws++xFL9VYlc/Atyleno58XF27WU3wQbQ+DaxOv9/QEfHZbtaHgnpRLzT77W
QQAv0MmCf23m75DqrtdyJlK56Qh+LDbqfWoh+uHjzT6bM7CtVRne4MsswZwenaGY
U019W65jKoMmBmnlPiivZP3HWUB8YRQ/el/Cc5cNOwgDE665UNbPNMPI91tFIXEJ
SOC9WtNomQ1p50psNASQ5EiwckWP2l7xWVfwqdJicN/aieEwNcZbX8/yM/5b1sG1
purPo2uCG3g56s63cpq9EACjnMEnqxD+XPKs42ci+qZ6uv/9FNps0DPCO1ubFj9T
t2Awbdl7So1J66OZ7yXbRMZwuig2Z5Xx3buFVXGcZilMRa4uDtQv9l//bQzbz9zl
LEhtA/1IpSLvF6uKh4wqAlaa7JHJel3rnq8iRXacOZuGOQW8P8TCPRpfUXwZdhJk
yueZsJka4daR41cz4OFv5Y3sivb5EOkFKF98Y8gN0xb5UOO6ePc5KFZ5CwXPDAkb
BYGiEPXgIDgkToo5j8Rr5aVigHpg3V5ySNIjHJ2cWz4u3xWQlZYkNfHMuAQx4pq4
N0rSVDDWC27oKvROyw0RY3fvLE6g/p4GSMfHbeOFYqWv7okHzhX4twumz3qbweRA
oiikhm7PmH5PDbx5PXhvPLdQS9t4Fcrwqb2/ePhelf1FiBBetAr7fS98ZhaYqMSJ
QOP+aztTltYhU/7bM69tkDpazFCdog0E6u1l0+0S0QD4W4r34Sy8TGunsSDHYSnZ
fA4VHEmJUe1IvJJPLbHULJ8TLktXDuUG4fHYBulVgQybwuvbtrZd6U/ENP9tBP2K
RXPF+CFUs4z+8Df+HuTLht3rYhw3HOTNyp81E4AbIJUmTqCq7kS6dX2WGsS066Nk
4JQu7JiJmG4isYFs1Y2rRxCgzvQCvzve1S44qUZM3PGpgeu+Znw77fS75Ggp9mUs
kSOZyJCzJE5WQ8CYrHlriaQhVtPxiizSBNr/X7IOwzB2xxevSCRIoC4slBCfcDFN
bp8bRXKtyNSyNgs3Gk0UoAYJSMnb5GwdQ7aH2GkADasF95PLJuFlE11uVLBaWNnp
0MycIhhCqXAGUbLU1i1qOEFGa8udJfh6mgPruJvuSeoBvYwWyZ2voS/IEj+AwiAH
FcFofNIPWZN2ZQLufTr/qhUxkV/7GxChQOTeu3G98C85S8CJBS+CovxIQ52wBirn
5u9dz4JFxQYtTfGRlKBruY+PxwNHRfzDPp+Mqn2wwRgmA4EEP2JW4deSdkCzaHjp
LpgMe3Dwovgy29efKhkTaR+KY0nMg0tmfuAPY1+UjBgnFMrk0l6ioUbziWsAQbem
nSPqb6aRGU4mjnCZ5xne9fOXYyeYVuvMvGwkLPblrFiuCG3dKX60qhp1pn66lSGe
Cp8ITqHLs+Zfd4T86wkM2LqrpnU+c69kD2Nt3NWb7xPTWY15mLuDC0PjOu/fdMfo
BWJouFgSY+7AonQujLTRztbRtJkWkhsTaWHcZTQKYWivZAjTJGxNZKKET7RqGEGH
/FEV/ohSquifoBrX22VsJGLlOwUb548189gNS0jVzYE9xl3nyNn4Rcr/3K0GJK+W
1ANQB+yfXRHcz+s9bNo1g5Rm/h6KYkXlNAwC6Z92S0vu1SYPPNFEoSvg5+kgH8UE
X2357XGANqMJO9GT3URJiFhvbmhj12j9Irhbi3SMc/0Q8qKNt8QGYvOxI2Zd7AS2
2ZbwFxncssAacuzkJHAvOglUutb2LvsHFXkYFMpbddtSGIT4vz8vJ7NpE6h5EvfZ
V9dRPk7lmrtZjJA+/yjZ4R0WpTlRn6QxyFP/Klyz9obvSvo5lwF19hcKm6rLS5y9
ReouQNljOucbiw1MfeeD0aJ17NxryYDj+GSMKjErHW8nr++s5xUWBrG/wxoJ4kRe
PifsNEMjxF7boY6kQxA7CxLqUuws7zWVfs27gT6h5kz9G8zGpwF9azjwOcNJnjJA
sbLdAXdPAel/Vks77V/C5doCnY2yH5Gffb3dMYfXl4MqNF+yf/NHCEsBCduq3ZSQ
C07UMSHPE7oCrLKCiEw8HAoWQvaeeLPplXZh98vEuR6GjhbtH/Ib8fDFMZVauqRQ
YXV/DpuAtF1TIq4cRtanVyJywM7JgzRWntXFpcj/25niZCefZ7wCoR8OWWm29Ksx
/pAr+Si+cf/U9D80v5hoOvB0DokaoCUdmQPeiNU29ytkHqBtE0jHcMJFg8jKRqOe
7SNGNlbe/82TMozXHfT1nI5BHtIqrDETLVt7beKPJy3f72Ag5Ubo2sAI+H+sdKL4
YoGZlcU0sHzuBoc+8HZbJZQGpGBFuvnwtfx+H4N7Yx3YO0qVxxZXG45fyA6MInh3
8BvIV8qF8xiF2ULjGNh2TyDeHlMN/Nzy4KZIqw504iGowT1ZQknWSE4YU1e9Fia7
wEPxun4be2B3LRKqKqRj63iuoS22GOVzxE1N24Vh0kSjMV3lz1mQ7XLsYQPksC8N
ntIZicrd0pXswJuzjvAvvSUdbtQR0E0J9t2n8JZRutTxqnXHjR/u/3VX6H/poW1A
y7H1yqTI/krZ5CuwqYK8EAJNjPvWdWPPZCuonRUzmxNsYmG4LhiPUdNp13TKtcvM
mDK91ayM3bMtpBn3Rr/ZcYzNn6nb3mr4WUOOdbtd6LJRaiRsR6Jw+wwywzKmlGvV
ktgjN8a2R2KxvdC+vVlGgKKiO1evoL7pjmxwT5YCZVMn6xRP+zAIOEVajHtGYFLG
xXoI6gh3x/aISizwCJehIah9aj/aqg1TroeYZE18zFxY7JT8KFGKE5mTEMEPMwos
aJpz8wf8+nSk4TCMZFytl9HSCkcyTjLoK/3mOuor9ZUkJwV6vYFbMp2iAczeE0lY
jPBHjE1Q4B3goS9xAFyhd0k/kW9xdqfpArposjm29MDyF8LZvN4crnY7yGGn/r4C
+Ob/a/SzBDdqiNUxTIZ+7ciVA+OFZE/zl0wn+G4KkRyNoJT7BU4oH/o2PUfdTC1D
eSZ6X1BOiiJzGelRrQzM06ugooYZTCnUZI3MgOYURUA204+51zqWyZothKW0tOUG
dM7ZHnPkvbOAw0i3a0OiE9gKcrkdAkhlm1UA4qWjKaGaYq7PJQKJWvHYQz0RiP1+
cQoOoFxrzLf4cjKzpLFCROQpq6F2ycAukupNYyuOn3pClhss7OqzzV5SOOrISce4
EyzhGQIu2FYOV99uGNvjhXhZdJH5jbU9QDvCMT60FxhdetRHtOwEGQbYXSTvnYB+
kvcq/bhvObFMscUa7td09yJQ1oOxI8aS5WyfU6cfrTeGLhmbLduaArykN3LCozu4
5ezhP+D1LpzFQmUWc/WVyGECJaZZSxdk+U0VwSn5ofgxtvih7HxfeiJuQPcmLHhV
6Sv8Erp39S6dNiHZqaHJmno98ALb2bj6L2JhHflye9BQLItXAI4O+cNKrndI4ql6
FIFdDjxxRydV3SrRWjrGmThnh55gsySF0q7vCRsLuPlcVAwMiNVHa5Nn0yMz1mSe
do1V27xk9scaWpDhZdgsz0ZcUuELaAx2RH0UlXBkOTzHOzheW/oLYoV9OLJ2GhGi
9kuNZhS3UHaBJa1SEgeqolrXKwqkNVuzGrP+g0NF2d9aW20kxkDhutJi/8JBMQk9
oDCuGyaWa8AuBSONUemztju3CdkvAcYutIJK/2g2UHychhLHcY6p3O2xQxwWeU7t
Pn5WIwvg1byhVSoTFtr/lqaznPFXAKNO88RzJf36ltdi5vVnUcPL+g9BjbEKhrE8
XrY8yATDehEcBlzsz3kR7nBhphbtqy7OS+TfwHk5xuGD7SWPWzTN8YdhOIYrsujF
iPkZmV0qZphXs4gg4HFkEaIJJaTGSedQ7NFxojSEs3sDbd1KAUGOs57jpBctZSz0
j3CJmGFxQTIt5l0ajnafQyauHc4AVyXBUyo+b9LsQ0ovN0kqxxZISTLOD4DB7WEN
RUxKrEbqIaIfZjVDfDBebkVgOS/KaBRgdbLIxjbp47Y7vlY2t7gKR8PEF4eupGLr
slUtkuqcr4VRTzht0hNc1hXfeerBdpJmNPkoiOp8cUt07OaeIljbJElJFmnZ5sF+
MdcXQMV+7YSXqSOkTw6dsIN44QXFEpvC0wA6xkbMwwJmoZlF09SLuDievzb/NADh
hdPORc89E5Z8/I0oFOugNl4nxgul/hBosQKYw2eaAfKIgOeleJZFwGm9EEzC4XJT
jkh+6HGlGVgqWn38NwmZjNRZBAAJNGA9tQw0vgM6LCppSE6X2e5P5FpD+JaTFqbT
q5RL/W+b886jakf44HZJDiVdSkf4EGYdvKT10i+WMokwjTq+Ro+N4H0Nm83GSRZo
M1a3IFAVT3j8yxNykV6xIR0X9vdzlywkivXje7Vc93vaKzW9PV++BTOjwSd6eiv1
c24sVf54xyC+3q43iR+Yb7B2HSeC+SW/Rjs61FfaZ36LHlehFa82qIFL3bJ5LeAl
4JE9GGOlb4e+Jelo6bWg2jVLdxJYkqvXnGUswWmkSayzsgcfOTSqQDR2MoAMnGB3
nhFN2E3ZVQfBA5Oa7oA/90g/p5MYVOFDud7ZvX0QOzjpPv/r/YpW2/F/dIdprt/i
wNJ2Yaktjg3tRQkO/gDR82stE4KD0+DHGFKpm1urXB3aR7suTFuzI2M/kG/iFU5c
Zr19UK4D45EturV8ncJxDq9D6z95tyvWUgfTMMwNrPlviSRmBtuemk7o8IRAWjdu
uDfBQb1F4ejwUAUahRrzyQmVAcBsA2mvmYVp78QFas1nI7rjHFk8nPC27OkstSbi
7u0aXDUCt5kbIZLQFZvr8HYpLCaVAJ6K5K8vmysDzxKLM8FalGVTNzTvGV3KHQIq
L524SBqslR/s41NDsfYtdPMgfTL/Pe9SlIcaLJK7CqLc41GMzdqrvo7mFCxFXxih
ZqY6Yf5cBsEXiiIdE7cNnCGEHGa5bfaPgWcVlhD5pQe2v1hDYbziiyh0u/0wEtkQ
N2YEjtcTS5imV328uEeVlIfUobr30Qp9/fBPtwNVH2Rnbv5DciZVorJk4Dv6bE+8
x66VE28EyeJwpveVmAjPUtOr1luNhfnqGAv6/W9f5IeA0Qsirw/z9aHTfEuNbQ2W
53SjL/OgyLSgQh8r9WIj7oWH4QOMlCeAZGLwiGw5zMFoEcNDErW5ofmM76v/n9v4
4g396dd78uzwIjdn8W3bN0K9ndm+o/kUckJeCAekIhNc4HL2FzhnFC66qlaAGpVT
6/kFaxnreW/SbXMYUQyJh8/JSD5o78UrgPq7d+A+wIEIVw2yyTF57MkljF2l4lI8
hvJ0CBR3JYHGkeWGsOpnhuhFhi0dIfq2ICj9lXSWzsnifPA6PVMf/88gD0rwZvb4
WWL7OZ7En+SF//0x8ME18KJxc97+tvVWsPiIQMv+OdB5cxsgelwhITzYi/LqFwnq
VpMXbAcT5UsgZJKIWWdu/NLAp9S3yMR65IKUNGrRBAgj+fFLdwU4WYZDRHeNCMhw
oLkjiYq1qoQ779EwmPTjsZ3hy5HKUSNIyUAYjkXrEoHwp5+aAVdkZkBCDFQIBijr
H6tdtxnag3Q7HMPVDERjpVsIkaOHxiJvuOfdbnxG2PL3AEkrzifPGDzPoowYCGce
GZHxQX+Q5fDZ2CuOeACLrQ0VpBUp+rUtW5Am3k7P0RZw2wIk2iq7Ik8vLWFrOiAz
K2X6IZ16lmqY8JLHNk0sn1PT0a8w1tq+KDgJuKlMKkI3mZYiiPINeF4pWFySvS2K
eLtXrzkTy6aUCiKI/8M5wNGE30UGouO8KojCGNKpa1TjfWUF8stbUAyIUQVYhZ8I
4/LoMqHVZV/GyHr073eS3r3bGVn1RSr66KX3nKJHyJMjh1u2fjqbbXZJuKyYQIEl
2nbfz/lpFH1luMgj832uq5HZbKi6AjjfExkYZB4fIjKr9/rW4UeUb8VBkSxC57ws
91QvkmoWeVyAA4SdGfSdkRtSUf84/7tIx/YrcVXjDb9SIK7znT0LNKMXCqjGSot0
cGQm7FhjulPhWGqPS0146zM51xChwVz04J3hnf+1hEXb9lVuT7dIHp6UBAV5GpQj
bdVnmcYH6DjWD+u2AsH9wMZLqL1sI6Q0DOnksSjZAteQFCs+uE9XKLwzqTwHZUnn
6PMgpb09MhV/goUPvR4g6jpOFnFgRAtaRhycYR6KIqRUcm5NJdzdNkhcUyOVbgxR
7pwT1hTlqtOIsx9T3LbAXTKbwFohGdaB1K9Xld6Sy9ymT5qneYnV1NJQY8DraU2+
jXMfQ+kLNgSt2PDSg+CdQaH6+aJqRTD0x6ZbhBOYcp1RmsoAiq520y9MKZx4D4wR
GYSXb7Vtjo0p7Cp56jIMDWONt8h5sa15HTKgp4YpF+ck8ZTtofpsJRjvsN4o6EeY
R5/KhNeD9dFMybfwPT+qnLDSUYgA03X3JBR4u/qyG0aLReSSRAZKMZTnPpC+VSrS
9ICBiBKHNqfnq0n+9evwCJqsGns6hKkR5PEV7xlfPyiyclY8BLh/KkplSPPSd8P/
+Loj0qV2d4iqU6x1+SsWC37himsXKFXmHvGFK6ftyR+f015JVzqJ1J9gBhm4wYPP
Cm5txlvMeLdxc1bzXN8nkFPEwUhfOwtIzpSGpdIVtm3pPgtGoYWQah2R+KlwUwhS
4/3xvyaWCfo+njmefpkmsT8hZxQp7rmIXIvWCV6R7/Qt+LlSFuuFthMzwnwqcKDw
/6A+Y92KUv6tfo3IjntW6KNTR17V7mdyHInek6nWtBUSfGLZBtdP5WAHlfsractu
Dvv3CRZStuSsBPyFr+g1bFZAadwixqHzk2IfMaZIF8YROdmzkS1T6APdM5ToYfAJ
/s/zCGBwGlcPxKaDd+4uIomnAxlnjSpJciJZOrXtn3j74+PE7Xr8zGrrDVuKFem3
dGin4qZuE/SiOGi37Zd3kIzt+4FvyMbv2a0aLlDo74JkVFNlvt1Aq/GQIPTQiuOG
w/w2IfKeAiZfLmlA7iXNGB4+IwqVc+X3JRMNGz86JFRvzpTw2h53L5PThXbsmuqK
yiyY/9LRUA5YcoFEB3A6gQhzwtnMERnorWYlBwsMWSywwULZL4MPbCgfHoonwIDc
hCwSMiTq3d4c8W4O9nyKGlJx1z1RVKVzHuRYFpEV73+6SgCg5/vh1eGoCC3SnVp9
ACCLkgL6dJ67z2l0pWICPSqaQsaUz95p9iegS5vcnaXvJijPI1LPMJQu4qA5g72W
NqZOtuy35hxcH86aJF/vhGbwDso/5RKiZqQQGmTxgN6aUQhnQz+PpltWgsITXzEf
KmZZIubkE1x0V/tQPfutbo84MUuNSEZs24/HRfoBgA2e6/x2YwzPqDA4qShEpRAK
PwXcYDmt9Zn+DtRnppNKglUMIIhcZRIM2utZQ5SJIPaTD2lRciWtN2ed0lKwQbit
3DemUE03fwLwJnPfHSidAMmFJr9rxwUdOMbTMwI+mkJ2GHxIqprLnN0upz/+si0X
VfJ+hkPwlZBmCTJ3xSAI7mYYmVQrxOJ0NMG5mCsYDsNHT42yM5ErA8vtBvJ5tVVp
RgIDe9HU57hZjuIahZWkcmUiwvedBGZrRKSSXPtsx2Yx1S20ZpbY+JcT2Ijc3cnZ
qimGneK5pte5j2cWTxUSExvB5pF+xY1NMAI6hI4gWicz5TlhN5uU/8mQ5FP5Lzr3
oe5C/yZ0seXywd8cfa1+y3LAzSGqP9NiS4mkwjUU6xmn5569FkoYKEOe4eY48Flx
yurw+Y3oWRI4mrIzUm9HF2B9yhKMaxSRwj2EbX2ABHgBVFIUefDOlKYIkNWyXXy1
gkLA7IpOV+QuW/4ay9RjXjvhsIl1nNYW/WCSDenqBWIOOq/0tpIuTh25OcF8+ZKi
k6vBiUvL9p5LG8wFDLxeZnO8z052pBDJQt5VWYJjjT6Jcwc8ZmaVX8xwTUh9mAdQ
hivIj8IyrG+bdyamISHajUewfhU/nluomnA4gc0WowOF8NvnxNte/UnqxzHAR3ZY
K4xz7xVFR174MWYfgMlPRCDER7BcJrWYq8+4HiKeAY0r+piyYHX4jZTtUEvOGaAB
YcJ4LU0NRc2+NwLSFZcf6ZJQ5Y/HlGZsvZa5fe8qepT3TDl69aPxrJJ1tVJ5iwTc
31WREDe0VmedxiNZUAWC6u3+imERr7Z7FJWEJ+6kT1ZQ9ei9+L7aKbuGOgj9IkSd
TPCbFSeRky7RAhKDWA7NuXmsSUhKAa+mEQOQeaK7PQuD2FLkCrmnkWunIefuBWVu
/iIl0+ednC89aT6CMalNmGWSv/u0vMr2DO30tS8YT3NCLUryNf2wTBAiveod29OD
704YQMgMfFaAXfxV+9qkvfCCICBLvkHqLPibleCrqD+NX+Nws0xUrpVjEgtCEpCs
7OX+stXKNaK3cplxXU81cTz7F8+sJwZ0iCYxUnQ6Xv10TQaLLi9cATSkUI4sPO04
YxVD8B2C1vWYvGp8isq+MrUv6RCrhWK0nzVW/VtF0ONfBU6QUlqhh8AV6oGO7d7r
52pYbsBc7HStHavXEx2sLVT3VqmbHDkXF9wYCYkP7eOUnRCPBx8Z+is/TGS8yDvu
DGvpGzbiMnH0wNZssFT3BAEchku6Jh5fBelupVBUI2coSGt6kNajgd8Ik8HikHHt
XSA0jYZt3rQ/buXK0vzfRxc8PhigbaF9CIMt7wyCPDZKo3GwL13udVgsOVJMa5mm
GcQowybbdAg/dEJRIYvuOv3lMzKkdNxXnWlxHXTxiD/jtgqBxd+f+QVufxvzwGqW
ZXsVcs/rZ5S3V2WWHWCGTvXWsezrXi4/jrhaRqzTn2frNfpTxT4h+vxjpqCv3Mj+
56CKGmCFeXIGMjigyohCzAsaBGXY2g1c1FZqZZK8ul5dGHOlJT1Bvh8+HcL5Pbsa
UO9d/lov97+yg3o/wptvNMiuyQ2uIivqCONpPteKscQ2kho84k02XDkiwBI9fuUK
N2RcJqYzJRuoFn5v+z9T0jHqhcTGmsfrppQSasD9c7yYX3iyQHqx/WYXoz39QbIq
Q1BLlB8vGn6eRuik6Y0O1B/etg57jmTpD922NXYMJMO/1NltdSiEVYbWENFmAmfc
arSLBMnNrn+7sc569twQJ7WIThmcjsU9qISyoD78Fmy6AcO8TshHoOgiFDv8niCr
fz1WSPf3eW0y0/sJ6dgub1TbSuZgPKA3x/gzEWLMBDjA1U4wEA+ObDK3Drm3Aem7
FwZWaouG2H5LPCTjU6vJRvVh0ik49I1AwKtjzIaFb4i3pCagpk/ciXKfj2s23X2h
HMQMvcD/hietwmgr4wWTv1DwTyz8Rq/h8w29/FSzcm66AamZPa6MSiEGDYnnRc/p
v/TXSRCfx/WqsOr+m9kxwpWv8Bw3Yzk2QQWI26J4eOOP9syd8KD0jhR9/zQjg3CE
Apy0pCwP7GgF4gR0HMpvcc/RhOJp0zHH8Luw325R0B6hs6aW9M4HBs/cveTkyuqS
6WncZ2UNb1FubssbrESgoW6IUCbNsbWVCH1eYbQmNrDJ8MXBrIR6jVkkDaS0GjwM
GovyBWG6J7dnn7l/mGnNLWQUFmDBE1yg6qJXZ6r3D1763iQsn7HtZExkBCsAoSpJ
3Kdehya0DlI63lmVUrAya+ILVHdrK+qR39EerzzIsZpAU8oX5xZ11PRKe5ia1/Ft
Y++LBdPVlncqXMCc6c7NdYCukW1yJUmNKcMRNVRfEDoLKZlYnesXtcfMMn2kVfb6
KCvcWOqMOOdKiQhYAtL1C6eKOoBBvrt/jZ6QMSutnRaQ/VECY2THv3MOLJxrMLQ2
5WLTKu6Q+3NS4gN6Aur8eymZR6h+VXe6wlYocMDYY1YfPQtS0jmr49sP8zp3o1bt
7cY9M6k7YjKtlDkhhHCYK9d3jT53Yxz+muwcxl2gWAFwh9+VSemjhhKsc9AdSVu0
dkGtImpJMaqpkafFGWwjMK4yy00RLBgJBdFBLll5GjUAlS8BfZq3UJYUEFo/PiUL
8shC0teZJpznqCpLL6YGAgDnJv9EYO2SaeboJL8V9ISoSlY/TzgCy0no4ctV0sDM
PbiMEvYVK23CXAW+50rNx0ZvyoatJuF4/R8s7p741I9+bVRVUYEYyakLpjtBRGFx
UambZRBpNmnht388Q618Cw1M1WUBOOk46KOFkTIW+i2+BPWj5zT7fUaMtQlyOFPH
RSUeY2kWUgBffoaqO0PaUAYYtThPihcIG4hSL0jCKtteSqRmJ1kq2GZQkJr1Vlo8
hLupZzUpHCxWa4m43jO2le/ApJw2u+OWKPkbPVCmG6D2bJ7qCbHMgOfb6rdqeiaY
tnQDV7bFSMLe1XTzogOFWudVxT3diQWkPIQNH/4YI6Hz+WkqPQufyiXgRWBsIkJt
AoVVwBxtkWi3DneymEFY9u4hgC2wHa2MvXR94SANY7+OLC2L570BuZNStdiaOuNV
nEQM3ct1QkjxXXRPHu5OkQsvqJJt9eQ35x2aZPbVN/8pl0cTeDn9NQGbAqDTolsL
fNfWspVGDmKAEk0zT6rgKrG9EJP6He3yT8c9OO1YWgoIHr7NoPfKLIPhPToYu2eQ
x8GLtErKkxAlv52M3xNAHDXXocY0XL9f/KwHXZI92hljOFtBwE+NMGC4rWaR/Ebk
Omq8Qfd3Ff3APbQ2+RdeRX7nZXwqqHinC/IoRFnkCu6ij+5ec4MMneiRlx6hnypS
R8HxM8ma+AI/xZQaXLSdaADUBkYY4k1upWP8J+y1hZj9JZOVvRlmGE1aNlUxfQNQ
8XfZ4wJpgU2s3dl3r2EMpqT2SWUzru+48hvSOY4obGK2sDQlVcO2AxC4E1M8Y3uM
iqeEtzMps16sQVEYMbwveUjJH3N7imvmRTLk5P/sXW7dDqJBvKGRlvCApjD8I/bZ
V40UZ89yOh5cgbul7M50zFbk8cMmj6drIZ9Rb3XtW52KE45E17u0Ao8/WRpZrrZw
73m9EVaVDkkVWxQOL84m990dazkjpAJCF2zdyVAQbzxp8c0Ml/bcW/iAPJ0amnUB
lgyGjFMk8tu1RiPaq/776tXhxjfLAoB4bcsP2wNeJsnMtdOAfIJWqLxxZdp9aJze
+oyokRAcogdpq8LGd7ijVz7RK20NcbEDkBe2BtevFwjyq+GUzey8QELBB9Iwst+G
ADKjegjPGXnZ2TotwrjL23s4qFD7M6Xmq3Ze1WZfTQdMnxS7+8ZWHfJcji3KbvyR
22xEN+4YnlburXf2blziSqjXfGpX7ok41345kLfryQVBCOj72IaZRjSIVeTVKss8
ceHRHK8jffUvIiQ44HDpn5PDE8vzeNz3lx20LgWxl2fefpfGYzJoV52Y4XWm/rCC
1aXRf66k0DzFtitkOMHWDqm0WImvwjpxccbBPPKPg3m8IhyDZNPlNM5KXfy8gWSf
LPHl/zMXM3NbxG31zaPKLUJMQXyAqzYgOGEoSAO0TwL0raKesUv74J2a+HhbfR3M
lShks69Sb76JQMGGN4NX8da+o4Nd8VRHNkPlErMzWcmQvvFgqX1yewxtZGThbwc9
8P2ENpZVRplMCsWmnuiDb3tjzXBtzdGG3W41Nx5A9M3tkXpB/g7ZkfCr2zvqkBhc
NriyI7C/sGwYe8oMMPDb7KY7CrL3iamuXvObs6SHR1go0eHcvtSniyHgi2HxnFyq
ZOBZuedl+vdMiAqQwLy2T+d1JNCVismys5kDlGCAi3w/7AQAD1MT78iUIMrdPNfV
SpT5y8sc7iKtfhIPsZzGoXwxcGcezc63lpc7mBk6ZiSiKYHXDeMLOggEEiph4+s3
2oSz+ieMyPDnvbtGGhgqcxh2ULKhI43OZACtv8zVUhjfiSeGUVlOMu5qa2BfeL8j
xSUxb+upJpjDqLgMq9lCao3HX/xtCVRdUutzjQ7VWPd9mf16TEMiY/30Ixj1HdID
JqoWYMSQJl2+F7QKU7IfbJUoQ+qEMAsgziYw/S3O0Spz3wJ/jCW/9j4sM0LfPnb6
oydPZ5INp5R6QUIc+A6nt4fgS2h1S2akZvlq/6xgInNkpSKkwlYXGag0TONUlIzD
LwsUP/MUlv6nJjyM9G4K384WCGOodaSYNmdWcFD5TwB/qAiLHZni6f5E1y6CgVhM
4GHeqPcxZn0wOSKildr3mKWTYcZwXbU9T7erLtbZvFSrAhnMDqqw6X1qGmKKmJbS
Dptyb1REEBeeqMywZHBW6um/DBH6AOpLx7WVicyvDFu3mib1sDAn5lg56f91BKJS
bhWtEyyawGbI6TXbXA0jESlTjtCZK5or2SzGeSp8AvXAa4LijeOwj5yERTxFkvb/
kDwC6nc37VMnHxwniFBylGKVlLe14Vl/oo9O3EwuDQka1y9rX+5daHU1rW/pkvcx
MCXlBQ6Ix+XKfcWQQZfkIHJeyweCYVXZyfW3T1oSweJj4ohah5Y/Y5CBTJaHs2Vu
t5w+p8AKbv8cqrB6E3xyRQPgpQ+Rl3yGCV4H/EMJxS1TOfBURZhJu0mHimCrWXh0
uGnXIEnzP089kBdtJrq0s76OzKh+WroSuYsJ7xzl2sVTHelrWpLmDwgo8OT0J1Ts
Zh4nCoEtxM8haJejPVsDvEhsvzu/E1DB7U3Up5Qr/LsaLbGBrF4i8wAH0tElxv8x
gMusDTLWcJvNlA4wIoO7VnUQ3xqHcr7ZCoG48FYjxnEEYCzzi6bhFJo3l5fLr6ZL
FZj0DJKO1OGoXTU3G2O4huxNibRS8LAtRw94ulAcINaS5R/3RDsFojB5uUENrVov
piEH+XHB+bV+f4FA4LFMDQioGyFZIrS13MgpvQm5zCmeth21s4izIfdw1gseNve0
Tpf4ngGiuKQnVVIA+p3DsRW/tgQA3hvuTo9+rpqD4Xt+D21ubWgfZ+bY//mhDZl7
RbwgOrZz2es0x0U+JwYGcTiRPzfgQUm4LFJprStxOMiWBnSjvEoLBUW8OtDu0ban
dx0DRKJwkdPOnZCcUQqSoJD4ifTtGk1gJPZ47Lib7nKyNTuOYAYkGkmsdLuPTayq
Dp49k6D95KRnr7bkwBhfieTOlpSUBXx2qPRxvVAYGLWBnQLqHxwsADrVAyNnv7Am
kNnWdQWAgfRZTHmxyGmQOezsBv8aEF3LVUe7LI7Rw4ABJ8EZJiOfmekN1Y+NPjrt
R+RR6mrOiq+9P1VhVy7jAnYGdVvt1oh20bwTbet3ahJWGJIDyM3VCyOzrZ4V2XkT
POFoYcnPshMF0R6szmCO88G3g/ruGjcLj+PTKAiv7Sk0WPFSqMLGkzlkqx57QIbi
yCgR59Qj0Q2tjXDYLPrPON7JBvU5glfByHzO9UA9GEfW5AdiYt1zPVgK4iOXtnvq
GPUSSHnMu5gCQ9gmnFaHLMfhU/bjFhfjjTYuU6mKmemWH3U4PeXcyvVSLQG3EtoA
CLgnyqwsNaZF+MJ+H6WeT9efcMl8ug/PdghKXnaIrhz4gbHQnY7sdtO7a38RJ+ex
GP2COkxeHbXzh6U5UUrQN+CRA8Xuv1J4IpgdWZ5b8Y+W+hx8QmshnlKS9Xjx/ITt
bT9DP7FrjzOgc/Ydsu0Vmr0/4fQDzx4nrdi9esnSrQZSeJuLwSjG40IdX37LJ9bt
LiYKUY6uQvfFgNn4xYe38D0gBOceGigT5BmEYlKnVaFoDEMHxJWFSvVDVwp9vxYm
kWv8unRsQi8kcnR5aN53l80YRpe6W5GBG7kel7ZdtKIicNtGJeI8aBgk+yJ3ywtb
Q+EVnG5R7OQA7qbigCwOGp+/dkzxtxwpusr0mkLvrAUBsadCn7BhKh8Zn2pMNM7N
vFRMsBfxxMcWfODDtjMQ803c02cQLup9VAgqswCWWCYXyJjUsr+6NUJsmIf0KvdU
dtiok5AudHHq1IVaJt7g1I1piuPEWLETU5M3EKHc4Go3Nc48P25vQi0r0T8YPNrC
QUb4pDv3E0L1dz/ijK+rbBrmRgNLmzXMtdxnUuNvUOZoZnXdwASstYjK52Xsj/fA
fG0n2TzGm0p60+vcIguljm3gGt5EcQ9/Ws2AF00bLft1edlLLc2/AQWrjipilQ0w
yPo74UgWaATH/bCTMWSng6Ux6HwC5L6xVcTqey/e5GCorJ4MFG5qH0bxEMoh3PkJ
r8zqqFCBAsH6T3rCapQyCD2oCuSi5nR3lakDXcl9OU5ip9ChAMxSR8DQL6JZa097
I1eKQscuUvwtGEdX6yyUf9VicN4WKGUOCa9YXnY9xnr71042RMjodI9dgifY6evC
xZez2XN2FrRJJeRy3vKslzyCZjrSUQRW8VP0pTVfWTm4v9sYTCQjSLz0J2/wtyHz
KLWVSKCGxWSbBOYGt0FWpp8zeHgTWROgH/OBzXrllhZ9Lg/9GvWskmMzvp3gmBVh
BXocnuuvmF5yoNuHUyotxvrUzlwN733oTkoJVbQx/LN3EXLKSOhaGOQ6nGMdwb7j
hEBC1nIqH1knH7veB34FqLJJSGFB8/nP1pzXifNk0uBn6xlOKrCHzTYsshbNWmvS
s5pHHS1Fkbgh60sj9vcmIMsOG+dqyukboO9BujjUVassUi1T5r2vMcZRXtxC+3wo
FxSSqNvnx5/s484a9iG2XZXkQj+O4Wc2h5NaZPI+mdTSldolbdyBGc0hU4ZDaOm0
ng+HNW73IfFP6Io4nUxFPi9ZkJKTa90vzVvU/V5KqqnEyACMvP5fCRL4bceH/YGb
fKD1CpjZd3hAHYxYWc48JHLC5Xo036l4TT2rMHbbCy/DqF+JlcR/N3Eiymla8LrP
0OyiwK3ZQg1FCX2EKvCVtNAxl/fVW69WPblmhX7C/WiJGB0OaaWKCBqlN5ChogOf
X4EkiqATQdPSNmeKMaFkfFJhzKSQfC6D3Ou+ZhmT1hOL1Rl1be0NYJhgaASIdjBR
PmbX0lgbDvgUADmGCLItw+4z9debeXFavhLddpqSSEjYRXl+O7F2UFmU5KGpWP1U
3aCyefOZQVXf9Qsu7sgwkz0xm/5JQ7c9zUn8vF7aKRfI+4YhHnDipXVkMLBX07iS
JTjrz7k0haXjrAlJvvCTHw+CZ7+CvJwIK0s6jOrasrqkrWV1CeN5fRyCUBbM4q1y
gxYGal7prLxm696ru00B4zzPR6F2haBxnC0KcTvpHKX/zfSKMSb6wFynYHLoZy+N
K65D9Kqay9nqooRpod2g/Rlfxt4X0t+i+2rnJS7pha+pVibui6WD9gZUAXdfODm5
bSnG5OVe3+r6+LWzYKgKH5MwyNk6wsxoFf3HQhommgaKNls9zz31+p8mnvsUuIJ2
ewsgELsiQSRmW3SM1piTtDU5b8FT/XneDPttFfCR2e7iQuSOEd1XDzweuW5CmoAe
12sJhyBDNRYVYwKi7sw1w4JPKqZug3WmvBW2IFSd+qFDoVx7sPr34sgeawS1Dixd
il5YphW9zOsmBM3QcE/Y5UwueH9VUWoVduy9limEB4e6Ad7+KkLVRo/iPP/yDwp3
nKn4GjD3YmWEPeJEyp3AtsMqWoQCBGkYquEAyU4dsHSpErEf3XEhXC1m1vLRcXJ/
nePbGmdYfrdEEYFqV4zpU1nLs3/LuSoZxYvmRboalmn0Em9lzTNLirp+9XbWcTBm
0K2KzAve+T90IFW66ZOtMzH/zh0gm/dW4/gX/+2vJPF9P+tT3LleX3v+m7TJG5DH
UxunysAcK51ILP+GIckRB+E/PZs5+iGaRBrzGtYcp+9Zz1YvSxq+GvecJMOHGErh
DW5g7z9Pi4OE6tjU6eE57pJu+xVaqdQiq9ieARLlCoTN0GEttDvZfo1GK8HmZH3c
2AYV8SEuFrdvaaU3rjNrRHegANXiJNG+WuVQJBrM7LzRFtKm8clc2CmtmoEWuRE4
XW8Kxw25bizeCa6VUIVj0F91YVxeS89MC984I90pI3aBTyTUwjfV5F2c9lqxtzra
Banfft7aOR/EIWTOG53L2Ua25cWqa3HKignKl2E+d0oaRo4/MEZai9rgldZ1PMM/
dbsSSMKlbw5/x/vuYS3GA5quLqZG406oOUxsmp8KaZNx2NFfjBaY5K4OdwglO1YD
6zt8c+dX8Xtw6/d5bhvFEUxUE/n1ZN4Fn1ks7EVYIL3fhMRc+wWC8SDJBvcxug5P
hN7oLNFvqKL8daoyC6fsh53KUtEeP7ysHcyDpPZqJ/TQf7ZxJwRrKSpUF/QCQPXQ
+796zFLWeXAy5bUYpnglrbJs54d2YXCWWL2cCUwYmwr8OtPK3x3GheCAFE7YWqTv
CgBJNVivkjOxCyhyC1iOnYcRMkzwuj0lim9E4EAy2RZSfOoZIjA9w4nC0AnjTi8d
rwHaDMWuaiN6t+o1G0RT0Q8AIgsIPHTBeCxsuH3OSd2sOJJrHAvoZfhW4XMXb1Qv
Cbf041/rc1/YFQZq87S4xOEIQYM/5CLJBZKgM3D7FLNPWOEyM3L1Yh1Mmb8ZiBIe
b+i3htDXM3V3142A0hQaUCdcpl49JUO/9sGnnxHUU/sa/vhBeOsOhe66hHa254CW
3mFtso5jq6HOFT0UE0xcmxvI45eAwIh6+EmqC3vH3uxt79VC/gOQgWbNGKmSO7MY
xc6xGzDhVXGAuQ9B/MDRxihSDe9wpQ8uo/CeY5TXoFILnT1+zaLlq+SUCafzJHUd
Gy2ynvUJ2WvxuWd7yhPWuhcBtZrKgtthGq7sEiu4MJj95UC5BY91dEpfdvnrJTuS
7b4voTlDEM7qxh6l3mtW8+CquZDcBZxVuCLxVIB3Fki73GcYtWpHkZVWOUTMrGuA
GEh7XWsbADCMFXd1FHqOSjlHIDZnKgqA6iXF7TGJrNKhSKw3bTARLa5lAm4+vix9
L41PQJhll0xMdkm0Zu4NFG3xkzvmuURifjBG/KaWBCVdhKXrUgFmB1q3BC/IYNat
WarsA2hRXKDANPJ/c+tjZ23yOsPjhfi0ZIS3yB6uqeZf6GMYz823mGNHRIc+m8cq
7EcoKp2yoUDX9w+4qvgP3qhPA9rB8sNBqeGUtDw5IRiq73ULSf6RMaMnlsvtkW04
dYWmfqLUKmtGQu9N7YGEYLPpFdITAsIYU1SQMmJOBJCWpEAbXfXktMN4Uh8nHIrF
cQar08BHOz4K7Dedne9phNp1YQIM4Q/VfUZxcr7dxk6saGQt931Rm4v+ybMi4HON
M+cY9iIleM614SMfrwtev7zG1qZ27UqowTrvAes7JaMwI2fXP+xUM37+PFx68imF
hKzEeL7+fUPTm6YR5/OSJygoVXN5TXNVQ0efPPoNk/syNFrqrIob68ySsosOzzXe
4AUQENJ13Z/bbT/9DnfHcVxOGGKPb8QvdF3uFTqLNlY5FWg0ChjinPAqCen9zYzf
ih7/GBTi9YKtyLwnfeuyLlqHA92Kou3LsTYRBrQsgz+H+oF2KB07mWsu+kvHXLPs
N76R1YSZlWTNZzNQbzwTfkRWRhVm6KCzOinIH1c6fgHrRs7Jdb9gjrPYIOJzswbB
cH3Yr4HoudP9dttM1QKYL+GDlZQKYTSEMbDZDf336OCVo8r7zKmtRwesTYg+DxSB
hUrYyhv8Fy4O67WY8+lcNBFyl8sMzYN5Nz9+Dk45HIHr6HqA7jUbqr5k1NspkXYY
ruAmto/kLs7jQh/u1icdmt7Pi6FrL2Du8o8KvJ5uZkY/Iy+kz1hXYL6Bsx/Phq7L
+UnF/4gp7vHFE2Y1v3oCCaavhjpjU1vu7hhaNn9EulVQjMi4IXx4mRunFcE6blgU
v65kQKCuSXWRW3bHd7CvAPzPyEQEJ0LjRelVV0d4ga1+mKfCqP8xXt2m6YLL5/xK
/UT5HS4b3TYJTOWE2FRhMtA1xxcqwfiwlKVkECeGlgp3spq0+rfrIdKU3QQGI5+c
GJW5BJgNUPcPe+p++kaMM8C054nUZbjQ5PvCkJswGxUGHBIctZXIhFLwv6HyDsR9
HD/MMxX7n0N0Pw9dvsRwJVCutMvnZbgxq4kARl1jF195/YQzyehKCZZI03FInOk+
REhyTplelD9hqRV9INgOi1Kdyl++8GO2fjetrbD1PHMrzE+KW/koNv2LIDr8blJL
NXqfs0iCOqIQ1tjEaPVXw8nvCDvYMediP0yUVxweDJr1xI/3vWV4MTgjUUDDTGZB
KXt/BDP4db6DXhgTdJrdzgwmcgMRSWkBNPLTGTN4gRO8SzY0VoABkD2BcF+zysnt
3Sqs3hJmDCkiM3NrAy3NZzp2mNc9OkH3FaYFjd4ewYu2Kf6KOuRWxscDncWIuQ3y
HCDM3DKoxvlqc5SbDGEEs6kNBRFxqsNfhau0FSAUZClFw5dMcUGXtMGtyTfEn4rm
NcY3zenqE1fHJ+1faWAljP1V5CiIDlOKYhfrvKRpwS4V6N9YcqLmyTozmd9rQ6vz
YQofx1yY5uZqtPUi8++MQwY8Ls5zpJcY4Qoumv47Ss1ryj4I8EcdOmZGsCmEL2U1
3f/sn36DBAzBT+4YX/AYUP8o1jbT/dFpiJc/WPUPY7FkiuAgYYRsqBqm4CC2FMFk
kfFZyAjMLfVkscJi6qkWhTtXf/9WGggBrakSTRZ6qZoOn5/VyC05P/3Dj+Gvqno9
W5I1bs3MseplzrfTwU3ug7ny5X/lxfp/+lIlA59lalay5PSYfz8J7s7NOykuzp2z
80YzJa9d4Gjh1iuXNCoLZ4nMVTJva4jd7qSdgRtSofXtbyr0jDr8T1CcxBZ9maCo
jqJ7PKn8EAV0HogwZGhOciFJa807AurbCO3QmQW7otN7pV0GYlFgxKOT6at42X1L
oZN4ErHXEYF2aFlRT1ZgcO9LGjBOe3gKy5Xn4aT2lr+9HYf4NxhL9rJTHUkjafoV
jLJuG73WuKGrIIUcNpusHLOAC/km+7IdZriBLJ+TAmUmeFvOI74lLIOBZop69nIP
EtWicabmdADDGMKxtFMjjq3Zctpp0bGWSy3X+HUf4Oy1IvWwDjf2GpawNHca+G/f
O4LwbTj5JGDJbsQ7lFSvQ9qcxE/A3M2Kt5wAskUG2Jd7sf7P7KxkBOaaAoNKfGtD
NEd6E6rmO+dj58ypvj8xgKap2IGDCLvXGzbi9jSyzmD/qi0ZBNXy8bwgmMH0HI5Z
NQd+0ayGm7TaHmQmX4KV43EyCfBEe5X2aH5oODuU5IuE6VLEYD+NlB3BitSDrm5D
wmsso6s334CakauJ4bdp6jEolccn0dIah4IWo91cfrijh02qeDvxZCAj4ieni+fX
pZxS5NW+XM7BTYP8mJerSDzZt8z3d72TE5HYUcgLSUJ9HrhMW1Y607dVqO15MBJe
/l6Y+K8F+8TkAqmNM4Hvdy4jLbedHOg5Z2ml0CVEuE8Q9OzdvvXMzqQFba5opr09
AU9A5bUFlJqBwOL4fxAXNfI1L9KIP2D8QNHQqQNuw4WO/8Q/J36if2m8zmNrV0FJ
vBCyp7YRkpzWFaoIeIuXgUu9QZWgYwlgILY0MTXYb9uGAdm/St9AZaohTIqS0U0M
lC0hVqWohW/EItni5o3RYCviTkNK/4oTbFhjW4cWFvemipTz6/9UPp6rrd/V700b
uIQDjdgkY0r88FtFroiqT9ycfAXZ69cmSuYGXvKx9PKYQk650dZs0U3l7NMWn2gi
+YbqbZe2CfPIR1MiS2ED1JPL2HQPKTs5XCdmn0NNd2WiTPS6nGRtgs8bwDR8CNfw
Nv/XO/8G7wMW2FjBWmQiWDYQNpdbC2SQV2s+KSDkQRodNmWFh3JxbdvVYWegokV1
jx0cslBfi+AymzttAuin/lAjS6fushphPBqv/xW0KbqWvaMgkmwvKeboOThbgcId
Q08bvrefz7eYGaKc0/57Y9/mZozLXwJOgILNTH9ukLGZH7Q44p49WLpZGq9jAaaZ
xEJ4AiWptmtbLyaovwaUNDRIm/JMgz2/w9PerPfnfqkVllGsw15inZDPhvv9ClUu
ay7We2Zlm0DCCmzxq7KJOEkXjbJ2mnyjYBe5SzkDLhYjT+HEHhaXWUiMQcaWxZ7C
EyyA1qf+41kw2v8eOz4jmfSG4lsKQKHuTURjzjJUv7AqWOTLnJL66Evi0JzRVVge
wnbRkv632yTy1JroZ6No/BZJaY9oqCi/9DC6Tsj9Cy2OQ5XVJQTZ++aqgSAyd2OC
T1qieKso6wDYsJAs1YxEOX77uPABZXH3JbGOLGvQ7xg8FA1bayYvbnkNnunEow7U
8PYH1SHHitCrEzPUl9I4mudvlvTVDyH2VRfrFBTSDHp7tmTmd/txhkupi1vDG5RN
sjv0oaYZrn4ePSQYhEZA47onViQJP9O6GKTFppmBInicvY7FQQBJqcv+Z0lCLsxU
YaiMQYjnxYmMWVASS5UdtXQJJbL9YRAA80gyJY1Z34bICtLdTSBd0OtEA77EBLKH
OxxatDPYooazcGtziuOwlXIpkWxaNj08m0dlVhw7WmlKtYBgW5i/8JAIXaIqc+Co
PCOXaNw4nomXUa11nHa4avA8VXSTenpiTtp0/IQ72Jq7R78Ehv1yFYzHDhbYrLSG
Nu12B5BqOOIu9q7xOiuGAuma/dCN2oNWItGUh34CmbQJ9E6ValhaIa7eRUNlFDtm
TmYVLdOZn2HFC5/sTtKM226iJRq0dZWHfbpz5vreWNdS9fJS/sH79DydEoTzCvwh
KJKDE2yUnjzCOCOEJ/RTSLP9JyiBsomASwYRaQqdSr7y79VKj8na1Yk/ZDcTr05X
cxTyZyWjhy2ousfe3eUjBGovt6z9coXQDfvrq7Cbgm9Ie7BMeFYtWXve1ys7uV56
onRLrl+jLqoqsStup74Tqqs2vZChs9TdaHAYxYQEec3PljVual/sa76Rj899R243
Qnpon8ITK2f+c86V5ssr3CCDAmuxqHPbgKmoVgvBWcFxTqdzhjKjb+NFNfumrmU9
CtY78eFaLP+6oW1yIqgSF67aHzRFYp7wHKONpq76kLGiQqR70vowrQAYtPgyZYO3
TyomyZTDj0P8eo/PXIPsjAZm1jkphxkB0qyPSSzuWGTQbeWUprir9JPyXDitkRHF
mv/wMbhbRmJ7OeebURjiQ0LXbHtbZM2CZng8Pw4ZjwKILfE+ujVhDEv1WpvolKhC
HHx7xsyzEm2+JGcGpgJHDoaVlVJmAfy+0UOyPnjPFK9ancbAdFLwOdkGJSgCiPiP
D+C/HBZN8QDWfHn7fnKHiozGItZrRiSmlRwAehVyYsbNQQ3xdPYfmrE+fvkTYG2W
I0SGdb8sJyhdXfO0cQ2r8sXJBp2KTMFA7vqtaeN7k5PkDzqBMO4eZDS4RXMNp3/+
SPX1CRKjbsul2OWmVn/tVd2BjZEpG16+ns/iz0Ciw6QPomhvSpwV+EijeuRUVi9/
yWSUxOnzUAF1o96/9TJ5mi3orC1m734MMbCLqR9cTIDVIYOT9z9ItiEAkCKV8Rno
mIigOLR1tmI2bXaXHXlvhgML9kJmcvOESZu/jb0KOY00W+cT3Fpz7V7NW6LQDfOm
BlgxcS54erIRYgPtwH/sD8yDp/NIHTpb63w/cr8/doALOM18YZ8vSWJ9HdiLncgq
pRhvqjH4cj1ahM3uvswfhoE1AtaCibK1nFq0k1ZUo+v6z4dOlaI2GNY50ncoD6MM
bHs76z1YdszNKZWD1royub3+9wZDLx62zV5EZsfn8cgCL5AKdWyeL2QQhQ68nM3A
FkpoRWJW+t2aD8XAC7TwD1FAki3iSOjqNm7NHCSb9O2+MtKPkrEa/M16eaRbPu4m
tE+1uBtq1hVkd1XwUTgKXEe+bLeAHtyTFByzwywhy1BY2fKsktEOW88ls77L14XO
yP0n6fXyDIu0BpVI11xvQFp13Rr+b8fDFEQaV7wEa/61OtcABiKMcjjljZTFRKdL
YmHx4Z+S9MZY5cxZ4EPmg9JaGI7AiBecgexZmBbWl+3euwE4ZGWYIpfguYnNP0gV
sCCg20DajfkPXTtoKIDGF3CzZSLXH4RuOxMOmC4R0qbtZeZZ7EodCHydys+EmLRz
2+9NFjr9MbsImJr8Nv3jrggeyLUnKUjN9UhwxAgGFR4KccrbzfCMKmPmKMwpR9i2
5C1xYNftgdiQt6WM7XG91IGgQ0dEWWYACIzYMKfbVd78W3b0P6APJW9ZeWaIESWZ
sgcFZ1+ZfQIpDfHCBa5od0RlM3G8QFD4hq2COz5KtaRWKQbN9w8jqqos/Vi0r8/C
4tnC1FpKomDJPB9QtY+NaxIcI0ediStoP/Y9E/RxIgjx4En0DcmPmAeij3yKjTdO
2DjFULIH5HZL4bpY7TbJvEioONHQMBfXRum39pWtvjXmv9MiCdwG5Pj0yaQKJU+Q
TxIsEBN+GD3FwMPiOOZSDAVgUc/px0Yy+pn1rIxeFGhH8dC1wDtBrnYvXjjnz6f5
5XuxbNtX7JTnMqj0+qQPfkq2jmfb69T0ob4b/aMTlFKo/Jrr1exozH3Alwx/kR+o
8vYcdcAblhC0nly8glmHQaA2gLj3M4TAdq/JmgW54Lz0gUqy82kyhdtXexPdTVTa
Z73xsCCxcTLpXrJXhMhFWc1iPpUWT4l1W6lTMxuMQchxsJ/V+ZV9GDRYPY0ekO8l
oIMC0fNtgqm8A3tI4jvhj/uXl2UTzALlKMwdRtJMPQIwqNe1XtKAQg+V+2XjIYRQ
DkpH72LuZc7U9SqV1by/11MlNVaWZY4/e/V/mCuliVvbM2H/WLnGEf6X8ay4gFkP
obYbBqBL0rdeYavUgH7c6v7OIyJZr/bkHLBalymthPgFB6MDaZVP9fdTlnw2NpDz
4tOQhJNVA/LK04bBfy5nRLuGGRBY6EQ6ND1eu+H45LWxjSMkYFylSCxdaP4cmrVv
hNg83VIYLJFN9zjO9c7vVObXFlVqxb3QrcJOHolGKvMArL21P2hXEMiug0pFE94X
LVCxO+FgT5IBLacCLmlY8dMh0fJ8jhCChEPTM59SmszZX4wjpX1hIPuMc9ytCCUU
fd9zhcjz0lnWI7a5IAIQrrT1RCt1718JaWn28vr1wMd1hpzKD6zbErwB5SOORA2Z
KlTfGbHRdXfY4dU/B0ogirh1+P3VKdPnJV9n5qFwpwRANu5SL7MCLdnJw8mUMPNH
qm9hGw67min2FOqCxAH7QluODtZqGisSywneyPBeJf5Ho365sq9N3/gxmgETFI+B
B39CWAxqPwAiI6797Ye3NoycqjO3G+B/XKBdVcjLxMfJsPVzkfeM7Z2gUsQFXfYc
IVQvh13UYD0IsYne41dwxV1BFUBnb1qu54ewFlcoGhsYFVMd2L5S7JWHmtmZKD35
3ZAPki9dcGHssJr4G5tRaZs2tZKOv2YOlT7zscVgG3lqMgZwQgR2WCz4dOLawHLH
aZDTlmC1TMxZFgabVYUDRsoyqlGYGJa0zPvakZaVQX7BRkFWqmTfjP6khwr1ZPsI
qIXaunErF3ZLgQia8V/mI1zsXnPjNpGoMPnS+Sxg/Gvi1JY6G5X28HVr7JYqXA7E
cIweHqudAjXFN0knx06xFLeWKsW1JqsVOXTmVirLdpp+cDBXu8zwNuzS2ZtLBxTc
1BEojlhJCTtBwbvyEt82dVUT4R7EZ8NEsdVKbHAuuJ7v+yEHFm4ccpljjT4z9Fvr
29qkmN1UIz42fwX6TTatw3iaU74WilmMgCwQxYX+XxVf4/8qqSiieweOOFG8sEx6
arUGmXEN++K6YihRFFux4kKWZ01zCzPSKsiYuhmaCB3RYBoMJfT8IUqpAok+e2qn
J0KFy9BxF01diJayvT6DljxjOCAual7egpgLaQ83CsAQPrwrtV/gHYrkMKeg2v9W
CuVIhlWQGzx8sAscqmR0gyIE1mBizqOoBJIdHZJtPHyYekGoT9HIbn0IQGMiz1G8
j98aM1IEhhA6iQGzcTeA7sFD4cMfeil+UO2tk0czcxYTqfTW+8C3sz1R/Pvn3ZLK
UBW5wIkBaB7v9VFbSlPEeJYedDOSL3KHz3j3Vq7pK8xtXAxyRQzzdFQ2vsGG4Aar
i+u/ufjW5y75hcnh39ptKwcbBQH4VxuSt/5NJx3w97iOt0IeepUjebXfgQKw5gs7
7zJK3ioCxjqJklYombq/1zTfNj8IstPGkStRm8C+U5h8If1m3G3NZw3hzWFY5rQf
jdiPXUlr+a+PRr7R/aaDHn7J6ZaP7hpNpjMEJRxVSJunUwgSUpvLET3EdDwiiwza
avzmC9oG1bO4p9IR1LdbbxIZ9qVSpyHwRaS8yFKEAdkWW1nWUR+HYvqt8W9Hz8JC
X348WBqM1Ttif/b8Nw+AcGSnChinaUezXCG4GnMTA4wMR/b4se1c9NBYW+KxoY3O
gQUzeKZBdBeoG8jpyI0ya6utl3ptmv63TYvlKty+l69GTairD4D294DAIF+3Jtys
+BF1MtHvwqHp4b0MRXYA505t937d6g736o78lqGIfrHmF1tU+f2ugivzZ1qNjPN6
faNt7VtuEqvIWqH/r4d4jihetRbcu4fo5SMfrEsNwCGoK+Ghp3tNpU2XhVQk57WI
jj/Cy+QG4s16lQLoN7lgd7p0OhSa0AmIJ0G46HU7xtbtfGvPeC4vSfjq61MTVFO3
wfN7bnobzx5yy/b9UC4Ks3/hBlPY0z/ZQNE3Dm/JUxBipqXeVhzxHgTLtMmqmAwb
Sx9ufbyMXW7lFrXT16yuian1hDIQPJKFgGfA+auP6uFuafa9zlzH3z2E4JEP+k43
mxTidoFx3HXFJLbeteyk/Vw0dahgFD9zpgKRH9lMcHF4m+J5EPxOncZNBQLpCqCR
OIQzK3/8oiA2ziwB4PNiS/AfLdF7wDjOD627LvAgwZD0CV/F6oeMp0i6rL8rxjCw
c+yOzUvIGYmArB/8SaxDCkMAKzxbTJmcFET+3rOfOnc9yXtbuBzmz5yFaKJ2bJv8
SVaPcAjePUXAZ3knzpREmOYz4Rl/7eiONevdeU0nKV8fki+z6bMet2KDIOha11Co
Dr9ONpAetjXVs0oGT8Z+y2KW2m5zC6TzCR/5QDoeqeL9vdnv8t+KNqOmVhiDvDcS
R8N7vGKpNf1ZYa1GykAr/nDeGgf+X1YX6KL/rddRngR8bpPWvmJS3BM+wT5qE3FG
q5H78Auue1h6KzwKqkLvvnuB2NHv1IT3keY3rinPevWkBsKC4xvxEESCe99CEsCZ
oP7EEUyzgVJLZg7xcyt5GmRBv2Zyg3fBaBYGuXIiiSA0wbg1ySflkOs8CIMurJUN
44urO+7/312CLdFelS4dW8YFRK00b+2nPCy0v3AL/sd1rdlalPpQ5eujSefqnITx
GwuQPyNL5DPDvpLItVOIKm1sz9UlikCD+CravDYOobUBVHyAAsu+scyoJIWDIF4k
ezap2W4562PU1xJls24/cXH7smP0+RwnFRnkd/H/ofPX4Jg6pPIs1vLNSuvtpoVa
hJmFXlBP7wiw4n/ZejKEcpIuK5d1IK5klsHclahsTySuZFW7Q25qo+HTTy2Y+6yC
022IXJOCrhnfrhMff00XXxL6gFvI00foJhp9lMtHIHaJQo190mCqspwzKVEF3//H
aJcD9f90NcyQVGPIllzo74w1xw1THkR4MMe9MPgaRZgYTKoXh+m62RQ7zFDvbItr
n0u2ofAXYRjFgDw2rM4Oasj1SATN7VokVu3pltmfBKY/BScmXFIRy7qSN5kKMPtH
1xRolFiNlmt9OLF/vTLxWnprl9rhVc0Bdk8/mlxChed6M4lyVGjyefyZdhdqBmNU
vbKPbwqtgWhl1baH5PloGYjVlLB9rKXvveGQ7BW0K1gICYa0BOXSoCuwaKQOxiAE
qJvOW/c5W6P5HIJZq+2D8mRqvgVPlEfLWvfJpeLD3k+dMyP8hk9+q11fvERG/5BV
zfDUVtLzY49QnNjXjX6mmmze5ZFFli27/8O1P9aU76he5jGaIQl/CtFXw+N0nTtF
FGu6FzmujMfIXMe5cXnkIOq6aB7ndK4cXjwLQ+4y0cbwkVlBOw5Dh9tkpJ8w+qri
Cg4y6OHOV01tFXa7q+eFIgFUhjUOwEbs4szs3Npq6pubqN16kCNRtXJSYWTAE6kA
2VGBfjfVKICGmyix4LGNzabN47c9M8T8nyfYKTIIQO/9s5VcZ9IZqehnSHMOn0iL
G/9/mZupg0jziMhOsJRCJIFhIhuuYjkL9MD+lIYaFoHaViao9beiuGvG9N1yDPXT
CaMSrs7gIqIoDsdxhawRt1L6KKXLm5h9NJ00ZdDf3whY96jN3N0+xsU/p++pJOzU
mx8qDiRMxYsSnEn61g/iaekBCXTp3YYd8VkHcwwZwZ6B2pz+b7k4D9ynpNjf2HQt
jLmdwDsopu0E5BCLEHiYRUQRdJJ33I4kF8Z7uvZ00AudtAhqP+Wc3F6rJo8HCMLC
kG4jIPhLm9Z8jXKT1wasEketDPSTt0LVkQV+0aufU2McYZEQjCAAz4piYlhslKrC
cAbASW4LonOY4ePfvbKTy2OKD+ZkB0xTFKBJJIuXcG1gvlH9sbFHfM6BEcGEXuHC
1v+WnWXt7YNBOMCqM9jMJJbSDSic9VJP3bPr82Jen7L1GLjCIiX+9cQoIjSScuc6
SHTPAZv+KfbwCXG4FsuaS4VUyTsr1fIA6CX6Eg4TxMLP+TQP0O0WG8qGLvhjjWRm
apoCmxKjjN1lVrjLAbW37ewM1A3Y5Xd8UzzoEUqzbmsNCtwtHuYLPTpU4ek9+hiM
PMVMqQWeF15iAMPMPg+JQhl1Qn9ik2olnvX4kpsr+mpfE96+NlJG1fsY+ZzJEZgS
BowGPDHhejHLyjLWOiKluFUn4DBcORHUOf2A83IHMElqsLJeG3CcIUQ/rSUcAos6
xD93ndsDcD+3x7fhq/TcTsqMmnSHkB6TiwE7n6x3DN2E4HgIeFcEiXubncbhTCcZ
9tm4uBJgxz+lp9I3bTBZ6VjxIkz8Njjvz/lN84xZJJ8r7KVBwJM0Jd5NLMVuW8GE
tRC3R3/a/HW88v2LkXsJj5pZE5YrZ2Vmtr+3cZ/C3GZIvSI52ptVOcbmuIEHQkjH
rqzF3k4AhpiBYQDLG6VRoD9IEVpdXRpXFbeKq9gSuLnTAnDNIBBqw93amwySGSVp
rgMU4TxSKHyDIQi4G44xa0YK/q8jQyodOQQsKq8MQa9mIZ4P5f9TZEYb01GltVzy
9UXSNoOc8zv8vboRswaUAgp3uyk3F37nclJgCa8jU9zVXUMexT07Jg0w8EBHxD47
Q6uZCSXYp8bv/gg7OLVk6LtRt6dE5nd2aFisWvDdo+qZz6qaa8HjnfkPP/CbphMm
YLHjK1qAx8ZlSwOXSuO89EKKatXVmp1Uj+IQxt8m/eB7FLgMKJlg3v6lRlToNViU
tafFV3wJQyqoWmuMAue1i35ZMONm2Bkgzr8a5l6IdDop5l++zU0rvwHW7G/OTV4v
qz9ryAEgKsqDw1R1hdycVoxPQvdsyoP047HrJTiaegUqE8JOfY2aG8tGgDlgxdTo
daM4dAj2ultLahrtNFtx02YEqMtmfx9wpSUF7NwumMkj60nl8VUPV1OkzDuvrEqR
R/SMz4dkaXpDxJh0VeRxtG+ENoDuhrlUoS58lH8eKKxbdU+ieVPzC8jJyG8y5Br+
Tpvndod9o/aLNFlhTiSDaSWA10StFA3VlLAn6lNmwLpSoU3hDYF8spfj437ekZx7
DSZx8WDs/Ghe4tlZnvhizn4/GDnI7i3Zz4fbhGGEzZpdv04ErQe+TnpJaGbRZhIA
EC263bptyPwii3uosdH6UaSlirSWL9nR8rmvgLnBYKcyRomIF3Y17lRTRfI0ddP7
nQTW8IZFChunM4nipaAw8afbceQegmcCAJwTtTp8FyYBpAS0t0GTyh9O8o5HsV3k
eGfWUFfuovAgJKkvJz6Bkrg3kicpxQ67iR4cSomL8QsUJohKohlxf8y3ES/DNO9U
VO6E6Jx6igAq6ZBcX7vucfzZUbVEBPs10ujAfERJoyjgksq2R/zWIFUmOeFl3VYn
lTrizc24POLHh5a1jSoHJPsT6NTp96KUqkf2Sndx5dQhqLpq/4Xr1i5nSfrsp7zE
CUjt9fJdaKKcMdpzxVXWeqrlXgVtO9uV6ork4BLt1Pqn0NDg5SVJCUXzlXaDCUiI
okv0APjt4ZKsNpclQbyO5tAIdhQtW0BGOQkkgtvi3E/wqVEPPeZfcOYPbuBqQqak
vhPuqt9ik9drE8X/on27PURAx3Y38FliesFchEguy2e/v1cKTRLFgFSfGMIu6+oe
TIgQXDTCmEVJWRvM9i+106hcEAXVfgu8uC57h34WKmoxeUbdOBbd3OwSLWru1PZ3
8BUyqcereIHDFIpA1d4qjD6HWOpAc34ERiZ+pY/NzbexJTzKZC1KAVSw2OYtGAso
IhjFoxYCT9irxTEUYhTcwJn412mLyiGGPAunYqVAJL8VOcSYCsu0afOlKxOl4H0y
pHPCxeFzADfJDVYZ2hvL78Ikun1btuQdcG/6x/mBfKHMsfc5681ZY+A7eZJAUzOh
Gc5y5316dW8Jfi1/4ZVm2Gaf5bms+4SSZMX8CCSjl4g0z37E1dMheeRcovO5VDXu
/q5n6QX8/S8M/p8+sqilUPYvLfdjDhzJ1kyG2NvJ/fsURTSjUMGeyrosGtdliwEm
vW5nImLcm43EqE0ZOGceZiv9Xl9UKMHOl3AAVAaUDVK2lOFmQY0WR2wbEZOgePdl
+ao2lKgMfwK962T5SZvgT+Lf9Z5awjpVIbMzjz7xtUwUByc1wWIakjzGw8x5XEKX
PMUinHsP1AfxU++T1mStUUfFA8F1IqkNru8zeKGef8pn7FcC0j2uahTc1Sz5gCiG
1km9jKmIK8e96tjtFJ71iWv1IZgaDpcRF6lsHfV0t1ifuvLrnmdb/BzIMhwJHnXY
MCEBgbBHeQfNLJWs19Hvn/JjsBpJh+CcwejRhtKH9PITKwNHaw1/C1JGkwnZtYWJ
Vu4drq+UknF/OE6iKD3TCFQ3q0xIxau723SLm56sQlm7VqM7h6UU1LRFc4flm89S
WEAk1GrXHxfi/AP+t/plySAarVZkHXY0POiDmu1UxD5q/sq8I4pGxo1KnTFpNFqH
Vf6ON2hoM6ySjlQFHfscdsd9bF209w8dDTTXXBSS8AMl9vSNrFhChi0FIGmJgAi8
tQsA6ru9DF+Xe7vKQhiZ8vXQKUiww7vMKESERooCbAovuR7RAtGzRXUXYpq6Re0c
OZS4rPKQQL94FE5UFF/TszR/xftTVOS50yfwHfjVYsOOESD+nLgelDH8ywtc5uV5
CF89d7+dBpOm7xES/qGw5OKfFDbsaicfdQSFqtl0AunYSS6g+iI7YeY/XHf8sd73
75Ce5Jg1VVWdvcUjTOEtiMF+MengSN8N/Gb2sYESI2iuKuriXKqSSQnLukKuLjz4
bW6ESqlGam175jaiX7sE5ZiMR/LHXqA2/cc8k3V6wLnRTO8Xsnj0CeJH5iH56ofQ
VJDImS5r5OWpd+LtR0I/K/yE6LCQzXMwxokeks9msK+2eLFDGRs5Fufl59fzcqGv
kbTo2L+7n2Ha7N7wVoYGdlQO0/VcFYVQvl1J0679i+aVDMwnjjzMDe5ppeB8cDj8
yNC2h1d9ouknIyjZGQ+W/6nE/mL9DUxndybAJz26QbCXbTp6+TPvIFAvLk+CQEYk
oDaGhkbBnd5lxkGKM4j+DDCqjhHtsNAeOSerOR8zcX/lzaMRLt4NotMQesty28Tq
ZVBvtkQGl2W7YInpX9FhxU5OB+m8+oyK5QETUg6kHqADpWtdcnqy36+MceFyeSmo
pwmvUyY/vuGnt/WAwyC6QdkgyWyaJ29AMX07XVxyP6ZPaIXH9XFdMA54AXHVADJm
5cIovvASsSHA8h/5FRjUC4OqXey/exIBayMWXmcDFRGc7plLRxeNVHgX/sGhO61+
UG+7/GKZvGpPdIQx1kP8ACQHnlSG9+0k27RzJPLBy1isSFvvQd9QeETJjPt8m16+
QTqyA/+3ilNazj9bwjKQ7l+DUDzYwUdTGzEktqO/UKvmje/HWLVXaYbWok/zLuX/
UOGo0zNSxwuHuFXIiAdYhtsIfbIDyWtSoU/6K0Cf7Jqef+xypajPLR2AWaL9dZbL
WWdNXtjJaTagB6CCURdRCak+f7TBselcLWZIUoUBlkOqbWbgzM1Z1Xd41LKrAcq2
WH75xm6BJKXVGIGtFxbOnkEk+fFWOewu2y0vTE2tegRrS6PYC99c+69JB/24+zI3
uzKuWd/yVUWajO0E5i4CViMloOrvS5VgLVj4rWFt3rUgB2JdYaxBI9i659uldVpB
WjoaVY6tHDepPPudfHtTNttCk5eAKw/z1srahXZkHSk30HHQMRlhFf5w9EHzu4dN
pxOcNezL/FjoFDP0wJWwlGWYI89/n9JpitB70MagEc7Syn0L8Yy3vydy/7zoH8KK
d740EGuEsEbUDMVRiUg0D+ADox5H1PA+vxtTyX0uSJdticVhAl+SC+pUW6PklpGW
0CMNaeiO26HVYGJIbN5ITKObAoW4X7ObkjLCWB8BioD0gwFrl+WQCsBTQDjLR6TH
/G8MxgoUPJ/iSOKuaOOpKClnh2dPgCRIduSSsm/KocGjjjL7yZXJkNrwMGhPh3FW
7odwMC2dlP+C61blHZ/Mzu92xLamvvncwaxrlkRB79wCLLewjhGMXM3Is3k5o02K
BuigInSD14iIRHpKXY21KnRwKcf/LzEtWvBGbGfBRogHQldP5vkIVf6dhdkZPlaG
Ene/zqhnUO82sGh6+/AKp0jwfu/7CdNppsrzdPMTLzfOticj/VWReSiwWvNADSn0
KtAWDrcOBPacp7yz6K8mruhkLxNbON5M+qSiAzVhpcGs53d1PhdlTo7wNb7KXiu7
ZkKUDbdTdGDZqTj2n5htLlFqLL4AWhi8yitWTg8gZCEVDoRY1DKqVwsEJ502Hn19
mefVfMYmXoeYGIaEopWG5UNnCYvGZ0chcEE2Pk6JJaX1J7FpQchyC1NB3kHiDYXh
xQ7gxFVpsm+aEq7wTnY2HHXHvBr6OsQ/uLZl9dtjkmyQyRshlvhVvlMmp8O1/PnW
4/BhmoxQsJhm+uGlJ3oJ+9txUev4f2y9DqkeFCGBM2i/6+4pPQjVcBofnKGmyliB
IAQ76jOKFB9Vw4/mbIMb+q6XwxnOFIwCc7ovUGPMxPS/Bn+cnIe9J61Fnr1vP1ov
mxk6RVOJWaJ9GPZ6JBlgETq6tivRNEnU7dbrcKMA1KAMr4iDKypvE+WcywrDFt0+
zWjnHJO7NakAHi1B464jQxyF5O/G+com9D2e6P1Ng2tGicJA+kTZUNqyB4TAJhkE
hyKZ6AHcEpJ2r2iB4hNjgUjaP63/YyS28aOQYIwcivkTvK0LBrkBRkoRKA1zEnEW
5lSMG9ylWbJOJs/znhYj3AaZR7DS3iy0OUr2iVMZjr6VY+2zURiXBehZG6+ok3TD
EgLIvNLdJdRxR997T9Jt5KHJKRcHXYI+y6wH7GXUJEMNqWBtpjcFKXOOR7M5ZWHO
CsNBJx897gS0gnvmpxesgIZ35Tj2E5IK4O4s5QOW539v+jLENASzAbpXd60fiSvI
HYS5zShvMrWXuOqlto8XrWRLUTG/pCnIlirb2mt4ZJYBwxBxwMHNsskQbNCUb4B1
vopBCtLERIRaxvOAoAR8Vrc/gmcw8TLs/gE3lWVceDkWGIEXHFR8DK4wixw7IrQ4
Ohz3r5a35ieIWnEt/x+wEqQiQvh5WrhEkOZ2o0wqX6S8foJ2sQ6KuHgFCI3xvhKn
C/3LM9nrR9mJY7R33iSD1+UFEZQ7ZnhxHp8mjvy7bq/l729W8uZUaI/2gqs5S1LS
aN0Y+dUuUCCriYllk6ClZv+hdrTf0Ce14KIJtbDnK9FIl+E0d0o6yJP6vGBC5Z0i
boO2QzV8oBhyEzbFXEPM0NPNDV1/ESUYDhEANMO36kq0U6WNM57VfwQ1hR3wQS5y
8QNEqk/OFgKUYUYWX8dUg7/zCPdYxMcU6IiU7ufrFVxWZ9lq3LLl3yKUFXYlktdq
EzbRBa7SZUN0KHFEk0ImaVP3CrcRiqP+UJ3ZSuf4glV2xJ5yBa87pR1O8PmQcZDy
lbYw03lkUEaaQJ9eB5ZqAh3jMw0ZmRCpqM3HBiONqDl7pP6oW9ks08FtdtDhot9Q
R3PgSGs0AesatPffcvhqRrOt/Kg/PbMUpnRPZ61xAkVTp6LzJLheoWvQ4P1UQp9I
IAjkpoSMG7rQHhKL64KEf1zUPizaNxxpTi/IcxVWVm4ZaJLEaNsLmBaxu3Pyy4Km
F2oStheQUCcv/14Aib+Z2ahlfnnruyhKMnemTwZ4xKK4YUjbvLTkUc4/0Z6Sjexh
dGENJB29+9JPI1aE1i2Af+daHgO1dPn6aKSGXtrWJOWF7JZJGl+1G9yDwCp/ghG4
iZm7WxjOKcbU3We7uWFBHZKh8W5kFR6BGfQsWDReHgtri/6uAxdSiKaS9Zwhy90P
xnj1INvTNoX1uG9HEMAjJXMWMVRYW+osyYj9Xh/TJ2YlfwrdDPOVr/pXnRP/Y26N
whS65DobcVYJ8Mz2tCkJbSNkFoe1oF7OR9J0bvSo68h25pZuxZtPQogXezudw3B5
711Sfyus/X/yqQjc73iS1+cTNLdQZrUgCm3ROpGZYKxlgvbo8dR8o4aHnoqcjtPR
H+7+LSvWu/rNAtd4LvxvH5QaLNrvHJBjemxl4t1Wsj5JCmGNjRbHmkPIzTBjnUDq
iPx7FxVTwI4ygWh7/s8p1M2NBKnfosq8qNsHoBSX6U7lNroHTdICHsWbyNHd5qak
GXhR/j0rAhyrCMINRKoi2/ZaBt0cRVk/hDYZQkidC17jWTF1u27PZABub7Pk7A6S
w2mZAzD7BMLKFJCIATtYGEO8xOV+CK7yVBPV64xfRCL0akKxNPXXLVMef/yW/hTC
Jq60Bt5ic+cfFmJ2Ef6oGOqTasOuOgGvfofAo7PuD7BQX8N42bKpm3DyZYop7pE+
apKlEWlwzuxoGwlinWcZCTkQG/3t+9pQPm0k1qigrq2IOaDi19+iGZGrdv2JW2kw
eDt+dHIQXT0TBvs5hnBXpSdthm0oT/xcZMXikDn4iEz2WaWvrwgRp7YMjzOdDFe/
QI1voUDXCcIIW6GxJ4zHqaHmdw3b2DJBpFtczAGPaCj1Hu1lqcNV57ACybv5PO0g
ljWKf5H0v/6pG8sLREUotm0Fv0BZBXCFW6f4+RAKsLHTCjr5ytrtgbkI4C78SKOW
r5gVcFomJSCHYq8deJ2xA4DsC6vOtdyUoZBN3fhu2L/0V5gDHsoWQEpJdahfT2/S
WpVVHfaWESWimdJFZrmlvRU1ICDW0HvoprRNAZatAinkawDxo3p2qm335jsoI4TK
hWpcUq8jqceBPKj5w4WtADlQaP4IheeGHjzVUhgdLiOuoGixeyO2c8rOOo0Xg4nB
hnIx0REXnWVKyrd086iTP3hndTdz/SgK4Q77MtWwYtNbXN1vuJFgUYt1CaJcvEC4
OscNLZfXVSZLozCP7eRCyHpEc50mZcDgJbh8ySppL/mZK/grvjBOrFjI98hXBPxZ
3uFVGcCh3nhtZHKyHfZQ1DULx2/Y8w08thWdIIPu175OYfyAF9YmaSSxIjUYD9z4
WPQnCpczon9ytW85svxEsjTdfqwqHvpbai5xZom0PDdAfjvM4PcQ44tsGS6i435k
mnDfZMBeXT7kKr2B74vtK9Uanvts29lY0hBEJPY97JD12OQoxXlONHolKLCKoypI
AknyCWHY6h3t69+n6/jOdd1zp1xOoLO+busiw9Y/NutBURbYXUYbbKcA3PH4XkHM
6/VrWnmWe9PqjtPgajhvm2O5ZaK07eVjklu6katYEX2y1oIRGXRgdrtgTyduiGh0
sUd90XeHYn5G8jzGam7TH4RPlXGxQNWuDcwE7uh6SKpA2jqjk/ZN1X7xKkmtwj6p
bhXHcC63pLX+m9qwAa8cFMWZM9CjUB+O6qj1fgkk24AgNOcnsFWWrUmXvKNuVaV+
ahpzZORVuLU664WL32ZMKBSyC3wOlutQac7LchfS3G+bFXfNiSdN5881jhQkcWV6
AhZ8x7RRjZdYzr/QSNpY/GfXxgakuhC6PFlGeV2U7xbNDYJsm+XgbjZhDuiGgfeO
m18ShsPY2op8OEgmB/opadVZ8q/QGy1qmtYVByQtIVpScd5bpMeKbSyyk8PwwQuU
fPeZ0LzB6VES3dRAkc9ezn/G4Kv5x7Lio84zN46Z68W2NmeI3viqzIQkh7wMpYMr
B4XQedd6adzXG/ETPNDHb2Mav71DCdHZIiB97m79KerJRMO6vzGd/834hzVOTtwX
6ea3L3UMP+JR9li6bioFBnt9wC/yFlbO1YEty3Nbzq3Y9BtLBpO9yu26iVbfYXyz
rGkZ+7JxkE9vuO9M9Q4HpOPApH00GfnqFwktJUTVtRDSaJIkDhBGae2s3jDkUkQI
zRcPW8Lj4gTUsItXDhcn+eHxbc02f0OGbnt+nK+YvVOlyYt8HSSyo0MvC1nuTeya
dZJ4oywXzQcCxTPdbFTToGd3YZVHNfb46yuQMVwmPA7SFLmVtYHnlswxNRCgylHF
92L7oKb9+pdZlb7lV5CmyoKHJhMMmVV/0O4ENPcaJaRDQQfKS0U8NnNwC15pD8ug
KKSw93N2KYWeNHYiJW93DKJpkC7mXsuvhWIMHC6YDB0xdM1M26yP/dD/XCKbR2SC
Xb/Dxty/CWJrQLzVfEjErmv8JSg/CckOjz7fFGtorpF1+kyIwcge0O5WKWuQYD9l
St9DnVPdjJg9PIxO48PYlCkGAQFfFOW3d4gMbi5gdgsDsieZVDH1X7M05i5Sf4L+
uh7KfT/4nvgdOHjNBq0MWWmWAtKFDTpz808S/IdBAqBmdu/C7XqXUMQLHZC0dTQD
mNJGRLkw4qtKkpcvYZKD5XoDzOsrHUuCSU9Va/KYAKXZfg4T1y37vNYRELR2UKI3
/HEKF1lQVJWbNvwk7EVSPoj7kuMLBuc0Xpo+rJJEc2lIza5IrtdHsyuZ/r/DA0RB
etJSxoR7ep4IRsNlBgpK7v2Yr3EcFGBcUYm1WizC4dEagLdTQL1RE5BknSVZljzO
jSycrFxztBwJvDML+LvhmMZKhvyLDm5XKNkWlkkuyjrJ+pDfesCal/ctMmTHHUmy
btA1ZTRvn0xOKV9OG0bwq5TAyPmfug8w4w9dXNOz0mHrqa1AG1oJORj1Z5Zaui6B
aDJYzmaqUKP/PA2VANpbWvBlT817LmveypxfwayAApacXXft4cPuavV5K+XcRWzo
N29O+BPoNIRCFZ8WrX8Re/OnAvfoa1IBjCoDBcDdOxlFYZdGk0VgxeLtZy7b8dDQ
PRgC6MWDnKgcJHOWB5rBrfdBf6ApQfYZJmeRM3g6vFDMz8vOGq0TDwT1VyMoMzBX
MaoWA02D7PMXov0exqfkNvz5dgxXSsXwKY/8i50XeQ+e5qs4ncvnXrAeLwoZdblN
M9Hiv3AN9ttJcKjE8fMpYFnUgcYqGfScCbHPI12VwgZOKfI99uUzSGeLD2zFBX2e
Ad3udjRn8mNVhoqIAwLbzqgyuM91IZXbjdeYx7Y3MRtCBR6VdxG+qmvg4dzs2LuL
BtctN/ClHmOL2foU2F7tKWNS9mNljY7ia4D4/kutZi58FnNuXoNnsVKg4CV0I9MH
oLeUmHQK2GE2AP/osgjPavfuDQUd0b5qMWYfpzgTbphNkSiDSC1mscnhmQHWuhbJ
R2M0FaqDe/y+Xv786zWPQnuYO4uDUvG47f32Lj5lPoHpulWd+i4eLheAFBwsTmXM
C8t7ZGor524BKs4q1+D1KJ111GDMFyavID6RZF64Skt9OgcCX8FDbrsDwqLHwQkc
dC99ktqlK4AQnKDezpWFy8XEo98gclJKg+E/ClsWkYtfrn4CCkJWaDOt4BFlJzH4
9C0bLJVVPOY9BH/IxwGq1ez8mUkuhTB57crFheX1m94hNrKmvuZL/G5KWsqVVNRO
AJKUbDFc3qiGgJ17KkGlXFsOfpSu0aBtTFm2dnbQUGbgyxuPBaDMdOCFswzt7lEX
mj96KJAibAvFAZyXgj0BOpb0VFIK7gAGszKgXXXCA+jO/7aTjWVZikRYPZhUQIXm
Q2FxxpZfp+HZIIuWQGxEWqDVmD+r0fipS36SezxsgO9LSD8e4t69R5USmxOKO32q
V1BTPrjwI4yAR+EbPE03Gs2636QKdFvuk/rMErccz99IBmqF8r/GwlGWOKPml2gf
x4chuiux+vCERYCGKgaq99Obr8YjlDKWqwJPbGJpf7ZyuZJU/DzLdp8gcEmPt5hJ
J3w07HDAsUjmy+URA1ziYb4VdXqQFIwRH6Yz8I+LnIq2rElTOU79wwxbqPUTaqJW
vEfZVlXqXs2P0yFHjNYkVY+s1roR+Z3NG9OIG2SnXD4V5JF2dVnpVExwBy7CJw0r
V6WKpYqG6dWzEDOZp5Z/jnF4JkuC4dI8BDGOmnkVS1bo71JXSPoR/IjWQeRHIL8O
49VxSDpBnOFkptc5JhK5kbP9379G25JFq+bSdbKCgjQJ8bIQLPPEKhCqzHl51xtr
BfYUHV65poMKw3xDItcFxuDdL0g6sqhgqHfnP24FouylV7nczIw2YicApe2ovtre
S/y3j8bAhVrACPonOCmX7eq/aILf+zIE1YjRFcGsZjk0gcwNllB8Xp2Amiw1Zfvr
LRDOdnkO9O46zEMAPQrVwjq3I4v6z6zpMxdhsxm1moZzzzbc2X8NkfYTTRoRX5D4
0VqSJKWyNxZGgD99SN6EJaLigx3jPTDA4E1KbGxv3PYrvRuEM3CZXRB8DvgEagHT
1qEIhcITS33mqX5wR39ZGqBCGS+MHOyPC3f2Uina5BEk1IHSVejvwlb3ibqC1obS
fnpfFG3OdCRVVg8cFL9LP+XqlSupiBd6mSNi/J4xV0lXC7RqkZoMRG3LqZbhY/7j
MawnMSszQrbnPkPzRNB6t1GBjyEKpz6xYMndQ/BXNtQTR7xLSzLrzo8K7hCL/vW0
Yltw2TwKXbTNZtNwDzaoNzHugw20HBzmqE3Psvqhgs9ZDDrrfw3BiFnUg8k2EDqj
a1gjoeqgHweDNtjBhiejWE+0tWcwBkDF0LTLcTosl7CYy8m5eRND32Xr39zH6CBA
58iSa2UIC8SBQX1XMQ8MSaM9vw/7fAsYyWx0HFk/gTG84EEQA6pG9JvbdDuEX0+X
UZw4IKXHP3rBJjuA66CqFVuihD419rpuOPeBojBPwO9+uC5o7hW6kl++GrYuxtT/
FyxNy/97l7nYGBvCEWjQu3bIyEPFsQIjkwk90KCuSiBZAE8Ia5fXoptnITcLp2ln
T6BjWHVpfyvkNhl7CeR9p14mvV6KdIMbSc5F9G+YlOE2IFC97JJkTZRgTNfWf627
xHPybNxgi9J5mYpDgOh2LtudZDEgaHoMiazZ93AIq0N+0elGh7ttya9NbCxFlLAW
XoGVdxypLJyTYRZ3rsWa+hysZjRknGJnTMetehyYYjLK0CmrOy/0hlWPIPezu3IM
d7gen1kirsaiEUm0ViyulwX+L02vb/vsyGeT/fMS0q5YyGJC31gpvTvfCr6Hgc6S
OJmYDTrH4jAxj+ch4PcGkVtyr9S3F4HzBHZ0hrR+R6X2KCMZQIG7QcOlyLRcQ+P3
lzBOT/iwhRaHP3bJR7tbatp1ax7EJz7hrtKCMbWaCwthf0QP1w9lwJ9q1Uy64AaI
KE1Zk/UVug67yACu3y/t+DUctPBP2/7xrscR/quqwWkXCRXwHhmUnm8mIljoC6ui
TdYyWP3oSOiYui6j1KUKy+wqrQtLrDIAK+3lDB1E7q33l5zrLw/SkHQgl1ywqEIB
WmesbPTYhdRPxtIPwUV34R8eLPhs1zs8EGTS7IaudeKxe04f5ZmXLa7s3EKWaj9e
MgGM4BAEKVgcJyglPes9lw6gTM9+ILHIDDJua8JGwn8wzj914siFzC7gx24LuLnn
rwify9mXF7B/Yo8/p7v3ukj3b3XsV3zcASltFd0MOZVnX4VF73HG43VrCklGz1HS
nRjxJK8nP19XKLKyL1vpSqMvngJlghgRaztdv1p8uvyelUGODkmGdEQgihLyh2xs
4f+p4F20vW40WZ1fp8hPo2QeiYHzhIHIhtYqIzgRqU78hJoaRyVIbUFgjhb9aXxG
bENev/Er4c6lcYe6hJUFwRV3AQJ7bvz0oiKQDLEmuBgPYb/5bMrzn5JquhDxn3gP
wWwACP4kNT7qEhlGMRokPzgu2G7XUMFVBkRvFAk0cOa9mLRGtZYrHqxrX+opZwC9
srceL92aY2MoUfYvWMG2NB2r7XjC1LFNaX7WieKQWUp400k/WPHXUaQ3znjQex2b
2jokzjUiE6qgPkXZmgeREL93YLD+1hLp76yIuWLgNEqd+WThi8cKNaF/XY45O0pZ
hgGbNmVSshRkgmHxn2gKHnphMsz3zu5lYELG19DCYAx2WewePCRN/1Wi1tRC9txc
iGvi3LzrH6A3MWZVS7tGBjNewh1MV3VjnzwamTW2HdnHkB/mUW4jcA6+BO6HNOz3
FxHkoeVbyjmzC8aCVh8vemZdP7TilzNdL8YSqDaSynDWNGVrFk2o3F2D7PlsEIef
yeVyZv6C4QvhC9DRstvUMctMXPz+y4sFux4tD6UGwUo7MwRPOSE7KpvLe9tE9a44
xvbZoBT+c9z2aoHobd818iMwzcuS2Lqywjpn7iJ02nKBMkiaVC4WaGOxljRh+Zxq
tmfjJns5gbpuP7mwRY80iPobNhoCz8XbpQAUOqwBCEAJFadmzYd1Koe2akjGELgj
UqdA9mLDy0e1YUJBbmhQcBG4GTR/Lxk4nvWv7H5gfr42lBGSON5te+4IyaGlFVvW
Dj4BgFS2ATMi8OzL80kDPCQC64pCDS2tPeJT2O9iZfwEd+i78IN3b8qMg/f0TD7P
7kVpujIvIR1BgNB3y+yv0ZfgGAqfl4GlDWv2Cnftve3h9gHvx+1LK0xfm/6vSvbT
2CviPCV/2fZivHZXGMG3/imzA7wAjtAIBLgVXP9hxGDfYwD3JBdeuN4KlFyT/nIh
PK7ZmPyzGjgin0Eb7IUWPu1LFZqgkeqvxFX8c8yqhOqYROc4E7R3DhFHKb6DfjID
zHkUuasTDFPYtNuTerqMXBS3eNKOhVS5qGBeoQ8JTRuGwZDD/S5IhhtVXOS2AjN8
9omyFOtEWqSiNQGNb0UVZQRNLaDHyde2OapmkKGEd5k6RcUw+KD4KuiZbz52mdqc
Nud8J3tcZKqyEh4tVKQL67sKNiW08hdPpUhanSJ2z/X9QEubkn+MjpTw9wZcVVDw
0GfThCVp7LHQ9SOL/CYdpnbXR5Fh7jwwt6kjSDWxP9R6hVhyRYcPSYlx/iHX2LxT
dRYvQpAq3s7CBMNjVP+y0FfimhtEcwxNalP6Z4U2idH1k9NoJWvJTgfX9ur7KdbX
n2zpzSCc7H3E4N9PUkoH8eVOmrm3rQtO+Q0deJy5oLhFpwluYm3dYPILADq2t6iZ
8DUKNsMR4jVuq9w3uhfxBPxhDVftAQdMO9GNb8xu9AhdGjyUXkuzZ2WCHsjgsZGU
rSkw/cZqKFbmIcS9G++/3ftY68u+c7/jmc6SpJNyab2t+XYNarnvD3ONH8nu99b9
NHvcfudX8sYafnxkefZqyskLysI3ERZI7M8Gwstkp7JQzDWwlzL3lleLmEZMRZko
BsnUE8xOFQeDTyK8sebllaVupHRq0oonGIcDFmbv5vHBWIVnO4bPNf/WJZMOoz39
vkIT6cV+57jrRO2+14lhj8r0CdFLgdmwkT23pfvVul3N2Ac/hUVLwyVzYmb+c0Wp
jWYcbDdN6m57RH8qefW81QRhFkMSNtBpWpSsQJgdhzES1bslTR0lBCvZ97z6kiAu
561D1c/dCIKoNpjCxHrdrROkAQlgfGMqgjUQIlWCujJFg0XVKNLxyVriq1U+IQyy
75aBE2cAFsPKttHF7JW6qfO7JVto97iNZwE2JYEgrt4wtbb+fXrZbAKD7mhYCkkY
DogLhgax/WP/dmK8bqTtzj5nMJY7jsTH/R9ufe5XaVnDopGSp5tjft4xHswtOc87
pj0VPB9CEX907/9oGtJ/5RE0QiHiK6JTCb4w7/CAIKfiI4TD5FkYieuXKAMpLEZ7
n/jM3Ams89scbM9fKQhOngoxl82206NzHWQwL6McvKJiTe604hiA/tK1ntERIQZ9
5sRqQaNqSf4W5//CcLaNegwGFWlL94mQkvprViTFMM8lTlJRYE7zy7Xe5UdIfKBP
Jr8rninVCCvjmmOvGvCd/sEQjT9XyVg/VMgLDETZufcm0rx9E5ej8kzH+Qvj7lYt
0w4s51+EfVObtlThEE817YWgTb5AoKvVIVrwcf4H2PA0SC4iLZA7Fbq+jStkm/uD
2BaxgJUHNMlU9km0G9rN524eNH6dExyZsnb3y/wmNgQtTVdl9oN2Eh/W0O9Wzb9s
+2kaj+bCTlkCt5TwgoiMg+MjmkoJ5P1ucvWDgGmRRHFH80zLPdMbxRtGJdHsIY60
3BQqArCm9a3z+lErxN51ivL1tITrXbpKtn0kqMBKKJjZv2thc3NirLHdo65bPZdC
qHLJI/EaafgybqsRA6oOj1lUaNxykal4S3d9xLgFQXSD5RTOpdSRLe4Yo2BD3sZh
J2P5k7lW1wrqI+Akd/+RnqIjOYbMpOGwzE3oRiCEM1ZIFVJJKtzF1n9LcREreVYi
daBrba0F+/BmUvE2Ga3XyW/CFDPkDsHHC7qYSPL3icwugvEAlgYFsBPUZ84yy2Hd
AHcww31Wj/JuvdWCIw/Nsehe3oqU5rpwTw6Od6j8Bndis/F6TxS6TY+Tzcdj7N0C
RAdAXuH6RRwVoUCNKpb/M49h5Gui4dUx2Xf0P5UIt94dx7T4jd/t/cg+CiisCNxA
dhK/hK/okfGi/si37dbdzgrqjMxVRY0wSSfi4PP4WItmX5WiP6ovLWkUFNmB8xZf
7SXVXCMliJIoomF7Exu4xu9OjpwMcRX5iv1YC63vY7pLyQKG1SbkY2jKxR5s2e6S
oUFYHNSg17/zksctuM0VgOg7gwB6cW0LSbQLbUNiN88lzerkPYo2h7UuucMNOrC8
I5NLSftqljwhChiH4qhTXLP/m2Bzyagza0YoBWmt5288p6o4my9Yba+4o0svDo9f
XdT6pI9DVWPP+EYDbnwMPQnGbf86cBGT00wZKoRPhaoQZmLA7eMyrOCVuFrOHa84
J/5FHl3gKej61aQ5izcfZwpJnY601z28iiBASK+lzapGeGalpnX6jvYX0KwyoTJR
EsrfCnYHIlNZwn/FG7Yzvn6jlgZYDZ6MjjDjqnZcZp2/LC6cWHUkiEgWo7OEKLaX
aS27U7bgaKNkfOIkj0QSg515ipaXUyghEx94aUv0Ir5n46yeDQa9B+RRY/t9bv2P
qoiTP/RXm/sia5otjBMeHeiH4cGYZE4sv/AR4+EMm10yHrpcoXXK1PlR7DYfNkTf
4YQq2+xn5uE2lgn4lD9xwH9XmfcCgO9E0yvCFjrVBYSEbR80P1TlFC7gpkuXOJk/
EahRRbkclz0KCPtiPKDUA5QLiMUMoJGy6FJguyiIrF5HYoAPdSaoU5LrH5LNu/qO
zJVVshr9ILFDTW9Q+h8H9TGGp+38ZBUgN3Vjdjk19rlSk+ZxQZEo7rqVnTwt2T4V
n71VNBWwH9L7L3cUBSTyUcLllB6AExzjgQbFfqUBwbg1Ocr6mFRJE/nz5lkgzdjV
UkX8hUhZ0jS0RdlN/2CDHCSbjnoNurCWPTMFFT5LdMjavvOo09/cymfeq3zfbM3+
UK4w3Vebu4HY7yi/LCfU27TJL2PSlNAgaG0NWiAqADpKLMQJ4C5xpn4i1BBjfjdg
Xfpqu5Niboox6BW5i8ML8sjg5mUcHq9Ri4I+/s1AIddbqHOrP3Gy139TmexHjdsm
9aKjIlrdlh3mejxaS+V7fkn5Ah5eXFmiH+rCGuhjRW+Kq5413rcmsHsz8Zdn+SyS
giSX47clsYP2zS6n4rlt/8eEpYtDyQVTzq8NWcVfuqCAm7dtpVExmze6NIQdVdIM
f7C6naObmsEd/m0/b5niIVR6sETkHPDAHkNbSdZGXbdb2rAf5O8oiR0nx/ifGiNP
xx2L68qdon79NzbixvdBnPCfCu9GFVl5cPbXQEeC24ACo6hDnhnTkGwCt9hBCwUW
A7bxAN0YaQyFynNQU+i0touNK4anOSSzDDa4KzkMWOymrwOLAM6L+XABpN0qs1tT
/9KEtNxR913Zr11PzhpHRszDAmZufksSRmIYtA9KsdXR7pzJTga2FX06s8w/CtH0
q5WBkkOG8pyjGuz6ZCWjjcRQLG0dzeCp6E82GFm5Ec2SYxKJpj96kVOjY+7Odv1d
BfZ+2M16cZDWmDHnYlMMcmTEiG+ueRVC1AxGbKxUa1oKojyIHF7Ua/3k5H1KzIh7
CwMZ7eEFsdqYH01phVaqqCUAuOWuwbs3XbEwzpmc8h7MIaiaMq6Az3fDNlwMrGrM
u8rhIEsBoTsLbNAlz5XAS46eW2k9jcVfZJQFZPgnGFnfCOk79eLqhmnIV56fmxwn
KZSArXgnt1AMjQQb70aqEP68Ogwbi41njhlD6HVQq7xBvaQcTjIHBOBY8lVQ7Dk6
2Ny+DDX4hqepYnX+5VexWE/ApBzMn/RhBbltc0bUp4k5hCz8Z9cgFJMSvZQmUohV
oL1Yenrb3HWahK4Pz5jcDLKGAVoEjTDKeua/kgMrErmWleKudBaGxHARb1qWfhK/
B9uLW6GehIe9UC8GrUkGq03KJYlYnVpqTM1k/O3Z7vy1cMtyRrntLKSGM7fhiQ1B
rV5mS43W6Aif73kyXkqqr/+aObh9tcfqwmYDd1QF/WTEbxVvAXWlxLHMH1VHDp61
hsB9u5CcMAHRYFCpibA4r07BEMCP5mYN1GhQivYllTJNupNuJ5U2MV8SK8QECf0H
4A2LA2UeSIR0504aBOfPSuj/qKu2HLYUQOlsjcGlr16wP5YfuhcBEsOiAKfG0dqO
E6+iFuNAnu9q8kFygCWBBS8uEvqqj80AZJbN7ke9thq8WQhBn+eDfNV9By70SohV
QX5jvyiKkGin15G0NeXN6ckaZI0BCEy7YVdBpal3wgU9nOx2/NJkljON1oOqubE4
TXPSi3gDmpadNcZj3HLTwREefvO5jqtOzg8mKAm3jc1RVmwOIC1kkX7axX22CRBn
qPgRAEw7wm0apXWDarGYHvYjAVx9S7H74HUJ/sn9lmRu4G+mFOZbf352mmM3Oubo
vOs6zqhNSshKh1ElpW6sdFyLfuk7pvGeXDXIx0b3ETv/oNtfdY4hAO3FVJA1ahQn
0y4vMpEAT/hLn4k7GFprpyoDB8sXHEcrHSy3ziTf9VXcgaMLi8Dt8OO8Dby3UW12
Zt/0ksHrD3gDPQKE9GXjppcl1DwVeagO45nhDi7TJlUOiqdHizbQBYs/K0SMPSS2
8enN8G4U4Bq8z9eedwi6RXqnf1AFl8NruAvTV1TYhpvVrCSc8LPIAngQ7S9+jUfK
rG39XDGO/FJalJO4DmvUm1QeRsZesbzU5r5IQSqebjDOBLZM5XjbqSt9k1PfoQQ9
H2WAxmD9SDKpFM1DLJVy/P0sjjdTltl9xeeRutIRdZyUr2z8gcYZv1uH1AnNovZL
q759iCOopQtXFv20RXNw0p05dGwchyzTk+Io5drTlRQDwgh0y0vgzXgXeRHVaozQ
13wMPpeHRCxkSIsQv+M1mOJmonJcC5uOjF7WkdSn6ca6oYdKXW1G07pK4uK+0m8J
6xoAx4j8g4pgcsDpfMTmivLPTWcQraEoAw67KnXQaqoznFVrelRLTKaxs5oao0wu
duYZVESBZ1s+QWYbWXbyVCdOMyQ2BBY1lkQvl7C5EmKdw5ZULklQY1TaWHmH8P4R
rsPN+SpS5NEVe+odyW4OQ/Mo6npbra+0LYQnC1hAwH6wVeufABLrCM9ucsvJnTBZ
716TA25Vq+yFojCG2GduJhH7KF91j4TX/g871zLkMBQp+1xWHLtWcYDv5Yj8x/sl
WobgL5MYnbGWr5JYM8UEJz6YnhFPPo7on7Mzvl4li5gV1eE4WZx3kIbkhYUV4IPg
QiVkiNDs2V91RIDRdgujEXy6CwzzHrWLRMjYy/pgyfdkmhj6HKQZJyWy0tVZg9cf
9zJADOaVhvPOdw7u27pc1GDhMuZ1f0DOfupxdvcoR35LKUnt/dL5N52skhX6pEHp
cheKFw6KLpJgDGM1oEWZWuzL6Qb2Z0laZMrPQIQH2BzXdqzUl36ynL9Yf9UBXnTz
wTPViv+BW7Fca2T2kYCSAg2slCU/vF4jsBzlf0MaAP3YObLZh6lkUAKqTnzUtFnj
Lm1aioMDRvvXPqsBOwUua5NPkP8HghBkATyAzCENCOCnVXkOrwgQuG+8vkvlHAQi
s2EAsn3Wp38YG6QkrKpWPacyi+Xg+i7s/BFQE0b2MYLnWQUOB0wBdIPAGyCOaraH
D9stjBgSBWMjwiCrPVjcrEjyJrYTGTdnyBlGMd7AagPsViaBQ2V8TSMQ3/35jZgh
86NMWdrWvIpHGVWzPbBrg6MkTy0U+Wne811dOIqXCDTJZkSYvgpR3dLxmLwfM4SQ
5K2xP9CmVvwzQd04B8aLQfyDLGsgQ8/En+8o4g5/58R0Q3d2AmDu8e3H9CHzRaA7
F2WWngik1vOrQK/K8nl1lqc8KC/Qvqi8bOc+IuGBE6d8vz3f4ZarRqzEH1R0fU2v
HL5zNp9Cfz5lgKVEFD1rr93hhGmXxA+sCGo2gb53eHaBQ/EIQsNO/mA6FK6Pedyw
IpA3awWlJAL32hMNcq+9LwFhhjEBWr31Ak+DlCLp5/J1plNSsA3ZKKZ+q3RZKuK4
rEkddKZZK2ljsK4XVWZMX/pOrEsROdb4NHOPVpxpzQVc+z3Pt5FrGg7yISjfYhRj
Lsiy54+fKmNFzlkFdPf+hjKc4uxCMvKjrfctbV/tOi3kfvgFNALcpWOI/28EyOma
Hwa4OR3saXk9EjnkfNqLgPuQ5jvjyldDNjXFvl1GB+SEucl6B5Rx+nHGao3lA5nP
D/a+pb+g/Fj55MbHZHomqDgRaT+nffGXPw4o01JwjI+vRtKCfkiaXX33MzWLusCA
XlYv5tHDn14dFLo3RdLOkbud470S0zdhkNeIbBs0KJwfS2UPjQlOocfCxdWqWjd4
FB3njxWDOLDrA6oMfUCiFkzArtsiZpReK/jIvi3gOhMM8AzqEn4AlYqcOB92it/u
VJ82Mt6YT06irTnPVSyIYjNOeRdNVsg1w0rE8JgGTaOyFU6Va3IWdg9n4Ul4JiUu
C56Tpt1xKnq0zooeNM3s1Lv+2dZJl2O53orOI7Cc7bjoltJfxqroc4r/ut0OD0Ac
JO2LcnR6nNtVgxzi7aEdbLhC28L0F+UXsJIGrXb406U4tq19tMV5MXvjQL0BeH/I
jjw4hEutMFdhoskQLDOdN1rXSDH7B9uAWyt71I0uvpi8Lw63vL7hxcPEE2rspEIs
IxMRufSDC0BLrVHkEzqoMrhuyZJyIIM0rWlGPOSugCR++KajKqoWRFOfnfFjI+rs
dKJqgvtT8HiRNflT6FJmy8aHbcgH86xs4nKZ5fEyfNU1KhrcAFxgn7hnOggHLaWH
DHEFrj2xW401PL7O73wirXaKczHU/sEE4Z5z+un/Prc356zcz0zkYwwLh1i33HYL
aLf8m2uCsmrjdK93jjlA4JB7wI5zQMhhP7H6qSQTQYQt1hc9WnxdQafo7MSqO5OR
V/fupd3MVVgm+eI8gtNZ50SR1exQCGWldUDJijuyI5wOi9gRbagQzJI+U1c2wAKz
VjDrrMgAZoxOeFF2h2HQ9EeG3zJ+Dvf8+HgKjtbQD2a0awStnis9+cUWZbUHACcT
JRILBkQTD5fKMkogHQKke21OVKMwRH4FfAxr8KYq8QaeD0ttHScr1SME/rn72Q14
vHzz0m56mJMKw4YoZRfPyLMbhSVSn5hXc7dNCuTelt0K2wRgdu9ixpv+LqELcZ6Z
z1MJAQqp2gINZPjJXiFOmEpi+xV86oxkgt+aAnRHcdy0PR/0DRXpKeyBmd2Si3TV
TyCteDeNYY31ec2E5r0ciyUI38bXbDjJOaphKg7nR8gq70fkUQHZnLHve7xdMBG+
2nzyfiGNoESI2tVwN189pUQ/0qh7pXw7rRbOEE66v9R3SVeBvitf5H5xjDukuvY2
sNFVEA3+moU83zOR35Z8RuwRC4lqaxQPpQISniuPASpYnrTSccl4VybHpvxMGmDg
OlFFDyRUW3YNOBoTFuBokzAcPzocmPjT32fZBCEVS9M5Vdw0KXvNRLOo3JJ+UDwQ
oOGBFDKzpu55edO1GtEkfOcReJQNpmIKUBGfBNS3mi2fe5yESNsCyFaiayBo0trQ
5t4rE1dWlaEi0Y6Bf7d7HbHlpyDOrHtLAH87Vqi6kJxbnSYYsGcFA+P1BjrudGtG
nKEkllONGEOAsOPRXMODzdqWiPAxSh2yA/v6RpoZTOhjO/H67lztxjvIjjMhe6gt
0Hw/aXZ1wc+3g+3cu9J3BhjUX6Fu6n1C7Cp5xJSgqkrbmRbHaP6/7ao+g1no8HIb
o+U3wKbUalX4503AKCBWPCqhrqN1QT3+hWa6iALVevvi+J5+M1JN4l3bIrceL4LQ
4qSyGCScZDZMiEWEtKh7WNEoXbgfqmyipbLAVF3csG39Kp8Vf4zqtOoSLf8mHrhh
Pdml1YVcy30ozE3T6zdJlONECWuA52BYdPWstYzw0ygUjEkz8zKBGiEUKk7QeWjc
g0EX5IceLt2tbOn4+YJTp3Tt8UwWNY9Lk4awEaPqYt61MdvWW8tXHAv2q1wyIU6M
OnAwWCRHNWQwVGqiYJLPuOlU4EXq2DZfmFc8KGNeynewhB9z1zZcG9Sf9tGHJuji
sA53NTJWclb7133ynR/qMH5Z9klVPqCXC/9Z5Y9OtImxE61yCawBOmVi9lzWABgv
sJbqnBx74ZazrC1hP04/Kx1xjVUkw1LEUKYZQNkCPHSm/J9agBvYQMwdno/INgKR
KE1+GeFLgkgZH8Uu8Y+USjGhmHzWeUqxob/T8cACygO4GtrBv5uiJ3Zafh7N9Vs/
yzn8C2xigzBaypR3HNtUqTAoiJkAJ23vHQ0KtyziKpvae4PH51Ii9PqMYe60bxxG
Uge79HJzgVGLLwQ2CeWD3hSukqME4JLGXQmxDDf9Yii8l5zltMVN6/4DbJmVTFGS
0EvmHDY4ZHdpYYIZmdVPEt8RstKXWt8P5s01c9/xRp29CMVnP8imt0sEAPFj+qLp
LR/WNpHz6dch1sQz6ldxxDs36qOaUMwHCiPFXXfxHWgPu2h8PGB8j98jP5QHqEve
9xk3Y9TUCqyTai8CgUPgCSxKCh7ztPkAlxHDrUCL7yAVwTLQzgvcYxoL32djIyoQ
APQhj78ANY8EEOAURp9s4SzTLDN0txDuBGtCKvgZ97rGhhdICtuSL0EZz4TL9H93
+IEbOtkALqN0J1cn5Y+lo54MGuRwbbNt4VlDG90Cz83gNTDPndtudYOjR/n0oPW5
4lDIuHSv4X0UB3WnjMOaR6x7M9BAHpF/Cq1xjhOj1Cl+lYrW8h6qXrYvw6FVnvRz
KU1abV3c6fSKtrOSGhPOi1zXyGThflVWShkfwREFo3frrufK6vWRdDgY1fzS2ajt
mttUaBgKROFFmMBQTP379FvQnrTcHNI/pIHrFaKlMwjR2IGWlql6g8IMZn39QAGx
seT3mw8pN1YL2x/oyD9pLyvqduGxpM9w9aZAbMBtJijoVC0cA7fLfz0z/ycRp/Ic
zXcumF5l1o4J/aTrFS9mZz47SWL445sT6bYRQIdIzAKYbif0u7IIrtzjoV/fj9K8
RtIgVCFGEqrrCujW53tHPuMEo83GaRXxhDQZG3oK8WYyRArfSf0fCcVv18pgKEsg
S38mxSUAbWRm1kAkirVsJVGr3TlW2WGJNP5UVLrz4oZwuCfzG4ZyS5W/qj/0DF5y
ZM2ZfE4w7MOGJlCd4rggQp9ts/Ywemu3JvnftquKspJsaPCHbBeO0aFag4F60KnZ
PuHKPH4FN7sm6reN6ODEw82cB/iIKTlGJxIEdXqrNgubiLsfb6UZri1toPRBpzxg
7R+iFOiYXxG07geOAbBPnpo7fY38ZiT0qWHZTUbI7cOBTLr0AkhSR7YzT+G26d5c
f5DlgWVE4nz97jNXiJ9wP6Y6zB/jB+VxxqdeCWXHw1eU2f6SXT47i5sCkMwRnvXu
SnsxBP+c/aWtofCfBZ68C1CIb6X0FecdZmteZXGOlwqkOGIpAVUbEfhF5UJzzaNl
Y7Tk9Oj4tRYAkiKQ//m6bJesomP8ck5HEtV88o3bLk3J8IIrlPR2OiQOIWwi4a76
Xht4KVZ2KXkrTC08TYFxCvE1T9OFwOJ7k+kWkGfWWfidAcTFyZfsnJnCLyOdt1gm
GefFjlL3rbQEEU3Pb8aycKHpXc1mWnVrYlf5+iHElxvWnrE2uZPntLxTiCPyDGLH
cw1rUd0twdHwXP2QC30Ag2vAGvs1b8JqRFBUugLtJI13C8T5L7V75Z7oF8NmhJJT
hI5rc31YvfJ1QD5Mazz5oflOxvpglcJikGdods3/gzNqVHGwtynBBLR+jPQp5PP8
168jr77EwDXLPDh2qSDUBX0PVcSjwgcAV+DRQ6qCn5Ww6YhoNY3OCBzhStT98mMV
ztK7bcxm9JEF6MATeIeelkmlz5py0jUuiZnxJpVP+ogrey00WWd2DIvkZU0LTY9S
reXw9l7OPUyNsDfgTjHagxn+V5Fpcy/x7vb2hP8/U9flhkBlRXFfBHAS0oHEF94e
2a0XuHxu3aY1E48bp0Kokql8E7fgqWaUXcq6d7MKQuqBpe7txzJj/4KLt1mSAP/x
lBC5sEnoPEW0N6/Im5e8GxJSHU3qNzxs5Q4gQEqCKOkH2pXivmXoc8CJrzk/nVJN
yJzd4kP/nFLoqmlJUJz8GG1pmX/6ZVIdgtjTLi+f6lh1HpWy+Aa4No9yw2/DKVvH
insxls8HGY1E85hPE1oW8KrFzyxfJB7HcO76DYchdJt1pl/yvkYN+5BB8/SdhoYV
lPfks79bGc1dRVYqAqP0/sTfiAB2KUz7jkh4LA38CetR9WAwcXgw+3qR4JrxDn+a
Wx6O4sB5L1vPq2hS/Z0Nz7AIdXaszLGzsaoGq4a4Cf+ox3RpTto2MNoQ24TGUvmC
JnxIWXLuW+1TpVV1mnsC2yv1kd2he05YjznqnXBSvH9LU7feg49umBTESUGIHcV4
lP2wBhqnzOp2idNwiZ0ioxpxY0MgdpsMAkyN2lmMmd6KwAcKLCs8T1InQyPKm2jy
J4WAvOgpW2ySkABX3zljMC2g67HQZjG6uVRhZbPhfgkK+X+yLpLvjevoEvlUY+g9
LlAmyR1HZtkN3iig++qCZDPGAwplfio7CruqIHFTqWRpUqqaC+7kp7LnyZizvdi6
Ny6UajTmbuuI1Gmxc2G4hiY0lcwxjsDo407UYN+vg4dtJfKKssXoA3xFYKwXCMaW
J8MC8KReVWYERvdtWcomxqtJPCtbqlzZwXSyvFIM79C5lH3PaRXxhMMGbSDU3SYd
hCCydgOUVLwZmmpos+uwI1/opaStUIbTPN0dU88uPAXVjkpe+Dp1NoXz4QfJ6MN+
FVBgNWbNqRYTl1pgpLKVgCqWhjk7uz/MZwWgm4iA4P6n7awCPK6fdwQiZ89wHDZG
/0sGg4htkQsovz/5X5mkKpv7lB9XdNwoc3IGcTaNHKlIjaIa++M7+cGViGUvQJ40
KF0S+OSld11LlwAIhxyQBEJrbt8A20OJj2amoWYyly1VqrD+zaAXVvFpEJ5scUWl
/9vMTslaCz6DXuumBBfLmgJ1Yb+hKBZsm6CrMJ7h0BCW2/2P4Xndl6RHswjv1KBd
HX8dE26byzzLhmhl7/CukRFiqpovRf0kpLCnGsuvGHHB0sWrTMNjfIb/abbj0xoH
5LCfDRc+4YbV+E2semp1wNKipvemOTs8Zx1zu/fVwcDiGioYHRVl1dy4GwhcJEZO
9mgW+EBGRb8s3OtiRxGbtBxpOYMkVSeZB8xIQpYNVm0Fw7fVX7xoFfuDohEyXgcV
5ErQMQUT4lX2v9ejzqMEp5HjtCHgHmEvEANuWqtnNvDdyymQr6mW9ZL6/KJzLJAX
kjX1POyUOAFSpv2dePpEJTw6U3AdiI/fTQg00nqwbCPYmjfrGVGoqZnNmyUUZ32/
vZQHyojOttr16yFYtHgxXg/vc1WMCQq17y9neUGtmbopBqoXUcwNTttuL56xt/nJ
WVVcDFyOxDBKs3AcdnfTf8Q9e8t7Buo6bFxeo5Rxp9h9KzXiVJCfgG8C/Z4jCT0/
hEh98XixCO+jQ3tDJ6s2/xU9oRFqOHqTNh6UQHaVS2JY3TR+Mw/MxHx36fMLiTfn
oHhLez3ybYYtG5Plrg/B3mLlK2yf4pEY7wZHwxGDqtfmOr5+5RdEkQhQbRZviuzr
Tg6YfWcaYUY9UDW8x4frBfgwESiB/Jw+QaFz2K/vVTLfeQIuCuPgoNCRJkQvVARg
kSFYE2GlKjsIOoE1C4xuVCLXCLgjXgL9BDr8NIEixbBq+PwVZitTTwRm83DzsP0G
37WoTF5Wv3MbMAWx5uXXDaCaxcy1UbrWy+lqeaBiNi/JEfOKUgYndWYx1qkVmG1V
M5I+ObSw66iRpEW5osgso2LTUf2+pt9iemEsLfJxTgAOjl/HYi4goORXg9EW7Qmi
DP6BSTNdsQpr7xX707EMnZXAodBTCXt4Aotca4yyfTnhUyPzAbgiRZmzaUvHWWgD
1IkzdOQ/3Wog0fl4DjsLgFWr3j+NIpujpgwWj+i3SoaSrddvW2GY+rp8gB2AGzGi
80015dKw+c87F7aCOsA7e9xjX+uddrR1PON2djObelDUidz3pPFBndwrx5muvDhV
jAm4NmtrfY+4j3duDJ9Acrmp0Ios2mk3wotqn2yjLFm/+UpXmm9Qjl1P2du6N8v3
JvJduhMh395eVFcRGn2TSFiNsoAlnwfTRv8Me/l9sSR2xT+nb0vD2fwJnG20rXF9
8R7N2BCfLyTUDpvvwRVgqAzVpe+j75KArNb9w6cIKk8JlyLOnHWPigjRD7ucR1Pd
7PSryHL1v9gfvjzTnGj8MSDMzXgHCQIvqfRI2LotZL+2ZZ0NHBaPEiC6nWSi6kAL
XO6AVRvfTvOWBhfdXkhvK/NuF57T9qnmkzHIHzLZn8/NDhtm9iBU8yrITIDJPYLN
Pe2rvw3zE3+JgHdjbOsEocFuCjsgGheZn4KGCiqqTfRUxShEujFRqyKbEjDnvxMp
HQFKWCpv2By2YsDoPHET1ipxWnsDAB04YneNGt6/S46prxM/qa36OLI8dPnvFeNF
rrKre6CswscPIgfoCz96MAOd4e0jQqA6xuueLvPeLYmhxI/Y+VNIFH8EuGbYpHSF
rsOPD4xL1zJJNCbE0XuUCYZDDsjCVQllK4AOs5LFC8ZbKdBFqM5JuiatTIjuTl7I
myD1gAHkdk8nj/em6AklCbhUVIigEuZ2j1TCKnvIlB3mzdggcOGwA1srwFVGaBdb
44yiV7VjR9R3aJTiOCgKZXt/4FsI9RnWxdchUPkn+kg1Y1q1m9MjWJJKvjoekjRV
PNLLBNjbFDlitZ3c/S71gnZYziYNS9EB3+g1Z68549HU3bkgZmRMJXYgYL1tbgH4
VP866NJsydYu2awPknviNxM3bykynC/bKCKBEvvoe3DEOctjag9V6tFptqrvLRAY
INE0sy/t5UBE+JwtBX3nLXTNWvmrdaSodJyD8XVcZjbG9gZlkPC7rIOlWBAp6rUi
0D4tNc745QcmZRf7s4sdiUMO9vKZ8agKbcxmemhZsSIDHCMjvEW285HQYafja0+H
RcwV0EUUVckhweOYBq/onq2+gb096z2a5enJ+zImHbcgz2wRSPyWtAwUbdLUSoou
o+QSdRfXLAH+8OHbzAIUAiwdk47ptryJxUodwoZTxwurPmxfPhQYFiFNOKZ/eZlb
asvOTlXP5TjnB6ufjjxH0fF7DSqfQ/2FLbOfVVSmc0e5BWCSKw+X7NunjslYytee
E+qXXf2dfuiEEmShxZ7HnqKXD8Jbdbfr9TEj8n1lwpPYB0bf6rXyFwzEa28oee4g
7acZL+UVzWk1g8bW58xC+pHifdVnPC9KDocMU+xYEEVyu4P5wgtXa0pK6Yx9o6/I
C2pke5Tx7yDZvVt6DItxhzHLel7NtBp6/unBSdgyM2kuJOqaZ2oUMQOFiVr8bVuq
Lvwx7nTQyTyv4rP9jotJK6xmSeU9C4LJgoxbsis133bNjEgoRbN7mRwdSBQFyPWb
v5LMMt1uazcxnWc5atMaUmvKo5oPoIXxmwABHwM5Jr989zfPN7TILo3dVriRscYZ
YZj8q1A1BFBG5QgtyRjuAcKeKaGmVUmlSyls43BzE2o/bYUVJTOgZD1xkA0eqXsT
fC3lw5tKpucO4ok9Mi5Mg+wqUf0/cDp00T8oHoUm4WXCdE9Y6K6nwTms+evyJNx4
ime/8fYJlR7YexwUbZdxhV2JuePnL2zfD+DPJP4qRIPlye9qITj75JiUgZaaihfz
BFQgriHWMpinUSthPKuNquZm6K1O2nWQEcMXsK+ibaIdiWy+JjLPbgFhOWpfiJn1
JaeJWayFk92dIMC5zSZ4AnrdhPXJ43h0gynvoaUBnIyGp4dBeZcvrRVgyP+Du9YX
1taooO90cJ5DeZWVcyhjlChsk9OBFClDqiZ0fn0OOlQ2PD38EOM/aVuFbsK6+1By
mbOIklvmJhgBxOJSRVFU3xpwWFt0LDjW/7YC5kHtbSs8HOJ/UDn1S4VO7pzI7bWr
m8qaagpm25EYnTfCpt6gDCTC8kkTxXyh5DfE5VsIHw4ni8xmTauhkiNITlk1EKf2
+5KQ31euXRHLeR2oJb6GoAZZ/I+7YTyM80xqQP8a/x9G+m/jzoJAyiGGxlB8jNtF
UlYWqyj1iSxQSEfu/y9f2MFV/uS3i5AeaJx6OipNvxpaNAhDsQgmk7jC3l56jw+v
4Gdc/pZHhUs5Fm28uR1jJHuLv4SXc63CccsD6Xf3xmOt2u9BvZ7O+/v7/9GRRRMX
ueUT87jLbxS6NvAZxxC/7zJWo5ouiT1Eqaytavi/xAxS1hypzdo3cuuuOtsgGm2V
MKRtgQ8TnZikuJ7k2LDzhCIOce8KglsQxF6D3wkT0eakkgoQ4jeNurW7Fb+DxXyU
uP9oqCaZlRPMfkaaC0016R2RbUsdrTdPJiqBYb1cALpj96E4wvBuVpX55lxExNoz
9B5er4m1xZYbBYWmnzevWGVftxWu16nEpezX4BXaOWLDw9zqheGT8A2TPJdh4vyv
NkCKisjo5srW+7n0SBgqjaRI3SEFdAeyRCYVIPYoAe8LoP6LyO5KiPYo+tvbdMTA
VbuHj7L7sJUMsLeBwnt57Nk6Xu2dHvPaNV89sZmfpDJXYaUIxggDkIepXH0WYlYQ
7tGYZwDLemAxK0Cc7FyKpeXDdhibHq1QH7fjSi0tFZOsD7h8D/r++rZlUb3Uj5He
eM1kL1cJX/dvfAAozbLVucms9f5w2ECRkzAbfdA74QA5sb5x+YbECRIoowzCFt58
TPmLIN0Nkgi/WSR/YGom6tM+RrlYYJxUWxEOzwuh8Lpk8k7T2F7kyOz75NBELLH4
mReO1b0ib15dOFiTuGNwI7edslmElhZkKKvaxYQF3ScYqGrXBk76LbHYpJ8OdFuJ
4lbASXAmm1f0GQXpYa7XbTZXAkx7I+CnKgCIA8F4n6q416b/jT7y1Vsj2C2hCWH9
KicgwO7ixLsX8ajXeCgYbCDz23jQZPSsFGrq2cSSxhlMqW6Ogz7MgvhS7WsnjVtA
rh8fk4inCAMhcYUuS/YO74n4Mn26nqMtML7IjLTcvvrcpIU7VxXkrnMwzRUpKZET
5gv/pPi6hQbD4r5IuJSsbbD7bC5cw0+YLRIlvKQis9ZcyR/xVRus52CepArTWops
ASM5JYYbStkAEm7cH4402JSzz1jr8hJEBZcjVoM3E1vsLkuTKHgf1mAR6lGwbier
Vg0BOb0nU0yACYKqOacIrunOD0WKA/+Ef48C1Pvi4L0nHVQP/Anxz+7KZrOLneb6
R8k3acX2a+v3hRI5FJTa/xn/98FjDP4DirtF23iZFbViNMrCSDzLqfXOmolAltuG
UtJAXnJV6MWoWfmj8ytIuE5YSPYQ0w0EUnnNTh5UAokWSGsBh/jg4yDxgzaEqo9E
d/oVjVBSLnVmDIpZGxe1HpwpJ1B8TjLk2Zu7CAIb/TBbNvrr77ZjD11gRNacDGuk
rIQ1a5PpdoYV2tgI4WvzAacsX497DSftaAbHTmio6zMtJL33mRwiwpVamrDyNl5s
XcY0s0jcR69V3n5tljfT9vpCXSVe++XRl9Qbvu6mtkkkTN4IXKHdp8k5N6l5/PJ5
hUbRDYmkhvDWkaYR2WZekw5l6cOEQ9Ia+LrB0jPoikGAxDtaMzUeN7bRzqIPF1rJ
4IxwtBN6BzbGZS7tfp0Kz7YA9+Qrf8+1a5MTTB4PiMJHtNGL3QqyEGfIGg7mmcoT
X6BniqSP6etgpfAvi3ot7QGuP2wIor5F7VB4ynuBmP94XVLalmKnD3YR+mpUKDRe
c/TZOzZo5TLGAnntg81R+m8hjKPnN3OmLKF7U0neiHJf3UrrEFqZSx1xt2wpHTQx
06+UwQlZKpKXoj+Z7e6na2b64VDBqR0FlPzOKh6G62JQSY9HdIhyy7srfvJaAn4K
+cdA2TWpUPZPwMJWJUJq/TLxL1M8ouuA4PLTeWHJhtwuWH49MAhHOTU4AD+RTaEZ
kCy3N9sWSxn0Cfp9XLf/fD4HFn7hQ7ulxPn0rJRMI0pbxU7DU3z+/UJLiZwlB8hv
+wMXZZxpMYhjDSz+GEY6fwv3ElRwMScfarLsquTTA3+6d3C0asIH2ePvaAMPkstB
VFpWIdOVim2IBopUaJ1IKXHqY/jaLxpCtdi353hIWm9YKGNK17yLqfPPi5FsiLAd
dQQNggSwhy2unztMDCKRS4XKmOHEkD/gwEhGfNnD1SP0vabo1sOSU/bvZv9DWJ+J
gkS3PONpiqt6Zuq3y6SNhIMaUMGNHmA7uNb4OkdqcZL1DJfjN12vBRuNVIqObdtQ
G8VopBWnp+QsNSVcKsJO5oIozd7cBOEEWZx0rBHyTOpDsYOfQNtcOgLOqRdtchBT
WTYrIfsko8RVdYGVtWnVjy+FMrQvhcrTSmh7e6SJew3z6seykiXUAxhc9VwrdldB
b2rpgL89+Y644vnoNJZQukR917l/L/8MMZWjJqRVYWZfLsaw8TxKYj6wpLZcJN7N
IC1KK6DFsC8KNhvjcupDm1e3VIHQF4h2CgTqUC+HM4RBrRY2bZN3NXKB2/rJHvbp
/tV2OXLxV81ubuaDv5+IzpawuYIlqHTH/fymIZrNQmoiap+WL4VRgPFNBIfa95F4
ADA41ehrQimt4yA+ADEJV+23rR4MK7/7PlDlimi8BdGmXgAvq2YQvvHSzUSgWR6Q
ZwOJVZari1/IINQ6uzAn0RZwMEx3dGjOl0mCcse5yjBW4qF0m9V/7MRltR+nfxi5
HXDBl/7t1WfQI08iuh7lSjDKr3YxDMA/ZGprQiOnS0z1Y/+hkCoNd6WTQOhZtiVL
sechiVjQfgA/XxFXqRsiRn5b6zrRucEF8iXbyIG58RXhu73vikhFEZ7CFPsxal6z
lfbdlAURkPuGMwKPj3gRStRrX5mGhQhzb2m9t59qIgLAGN/D+Gn1xEvBtS7m6Llf
V+ujty+c7JLAMD9WJru8SZvsNuQjDfdsAmlrsvywOxKt/thbvXvYCXIQeccOx15f
N68nl/swULDzF4C30zWHxbtaeGq+B/8r72t6LQR5kP8wUxLI70pfq/5aqiDyREOo
Eja+tmHD3wpZ2TprQ84MLF8tJ70nZnBlr5Ai1c8kAKEFbU7dxKCZdhEbAeP47eGR
Xs7G+GjaQMqoM+SqkEhUzgR46Z/XxXaiz7Hxqh7IdCwgFAlJZMQxnWke7nsJMmTF
O8zE4BWsZ7aLsDmNQ3yHkh99fJRNHHh21g1AOMeNojLR6j0ToJiJqJuEoj2lJfya
bM+laC+Zibp/hhrqUC65Wm0mbntyR4Wb0ce2PbFpGEggS5l/GkR9y2ij4psskDKk
3yeg45eTFFeW4MsPiGJ1N8W3jCwDtJnK53jdGhv8fhN0HfDd/CXHdSg1ggSOZ3xZ
4mSBiQMkwNgijKQG3n0Gsuq4OeHGHxx3Pyf/DFmVWy22HdzGvmd3MchmpJ3xcy0Y
KraUPdO2wjITVqKFoaJs4EIxzJHWhpHZmqctP5bGKLS2YDiucmV7f84FfzcC0OFU
yy4hJhZIP77/vjCWf5lpcsLJwawZAFsWfaznfq3PwBKgHe1SYv5q0vLCkkOA5ePQ
AFUwvSOfnChPy9cG9PMvnrwM95V4EJ0C7epKvgyaID4JVorZU1hRTBwlVjMXJ05b
kUYIyIOKpoTmQ7iAgncSQcr3wf8LstJh9//yP3ww80OGc5Q7eZHh31LyWcKyxN2q
I5umF9+OF4NPDJwP0ONk6kZVQeWWaxKc+gz7rHITFxH3eYHzNJlU8xJ5tdbduylq
8FBafSQE0ZbxdHmiNHeid+IkiiJ3chM68/Q0xPCdqceS6eL3IDWeO5+01uelqoNv
Ke64iKsYQJp9Csfng9+vyc/Z9b+ILI2+HFwf5yaHZsA+TC6UMcqQ0b4CWIEQ+4Uq
E7juqJ0vD90q2mMNWVPGOclhDa5m1hk+CPsG/X+P3fYKNMoHq0QZCdsA3XrHhNqW
qU9NT+8NDXMiUCt9TCkDnRmVhCjJgyvvdvwQGl4wAsul166AYP4gISR2sEQF0YSQ
SxiTKO38VS+ZG9G+iWBY0qOwcxFIPyd+c9NWJMIlBdCvQvF37zbeO6QO0vzUeTpK
Fv2b3rzwZzN3a4TkMeFNxId2YpnsP0GGbAx8/oa3XdYQkH+X1sr5z1dGZAYAKCc7
0i8NrTIqO/khGALR3zN9A2TrzI4rgE12+IxMd8O+DVkN3hJ1Flt6wXFAPD7Fur6O
PF01IcHJTRcpPr/5lriohetrRlzdGWIXxZRq7OWR8oR0ul6HTMQ4KnGbfCXed8IX
5tZRXlUcIIJ8GCntuKLYVg7XmEoHPNUo3J2Ej6mvL2oDaGxsKzRucOxMJJz9eJ4P
mLted4KvzGw/NPQ5oJ48W2sK3t9hTBuy8gSiHvKjwWuQ3q6q6iST33m72wH3VvYU
mfzDtUfK3znZgClQa+wYqo0DcVTNnX2sDolDAmiRep+NsJmQHJpgjgDetwQMo+OV
SkizUlywWGZlIC8vkRkhD7y/JYsixGT1fRuy8g4CsOlRqRr1dGFkCQGju0zhR/fb
725ncJOuCAT8tA3IbVcsP+TFf7g2QvwAi5Sm3NtjRvmJLwyhhiROsmfw59ecO0lM
L2hgH/gKToVTdoaRlEP5f94YC2tsVfrx+hZ6u7omQRcUTRfphIVb60+AWDZeJ1vE
ybXNE3KzXiNyxwTICkF1nieq5ym3Fo3CAyoYCcYuWPlwuMss/Emyt7kWTkU7qrkD
E6wrbI4PX6yvDM6Y0HDtXOq0fEUF7HyJwWiNHtssuO+NldTX37lovtLDZYhRNbcp
iDu7fNaC+R+Zn9YtiqiaWC0SLqqi8flPFuptMjPUV9tDZ/7ei45RTkLkXhBiwHXX
Svm7ZE4oUxxjgCB+ql26hfQ+AZJN+Fe92VXkVRnloyVF8xdD20n5iRu+97vUXej0
gYMSxStRJbTghBq90Df9aNTdiqYx1PzDn83L8uSgsHe/HCL1oQl1VVw+Acd+m8DO
gPrJ6dMBl1cpUhVK6UT55ZwhiDkC8cf8zhpW9XgIn0BqJNYlOeogDT18zWrMcFLt
BSc2OhZt+8Y1fVxoqqxZc1Fp3EzHUy5qFG5jfJfypEqhx7agTicfTAOkuIXuCXfR
6C4Q5+/MdWgyUVb1NvHls4qbsPjmvBer1DsNwN4BLqOqTvNMpYM6h0+GbkcCLqkv
WzhNzu3CtCtQAsqhmPTvpXOEgga7MAljRMX6mGQi6PUEclp3hC2BZS6VhuUqcZ9h
ssoqJVSO3mE4X0h/rFaQNz3ja12cArPnU1yAj7URwkAZIplJqbcIB2kEvObZxzeS
XmYwSXT0gqgptEOPzUuXYc325x4TCon23mAzq3jRlLvMRtI2kE3YLxUEaI7BEMZ2
qv/pjXqy4wsz2DBNSVhfRan+/Td4l2rSu7PBU+GMO3PjeQ2neNIclIGVKIAPkQ56
2MfYDqxUiN2HsPsKTCpxDHipzP40JPPQVBVEkpfLy+jG2CGZO9X5wdYgjxZYuVQ3
OkzkfcdttigWHInBKEttnDteFATYChGN6iOobeNPlfOXOXSvJ0QarCRELctFYgfK
qTl5XfCiIuX+lcRz2GMhSYbIsi6XuzPWUkRAQEEhbzv3miIMMewvJDI8BS7yhSua
juPjT6J4d8jxFy7pKAjRX6/OnGsSSvovNzancPc4lagy65DElSBIt35wFnySENEv
MaxD0dzLaI+h8TS5YQ49CaYs/qUS58LCaqorPgHjR4Iw0QfP86dTX5oELzKrLr+8
rbZOqw1Z9KsiFx4a1FxGRoA7gHRtPpkO2DLzsOY7Yd6oy0JQUNUvLr8r9lNjiCsM
XTAc+vs9IFkyMDzZ2cChGUMfzTVUTRDOT15F+A2w5Xrmp19GaTZPfkwqTwfJSHUu
N2Q6n9ofKkDpin2i4hpwIcIozzHjmWI6jQ4c46nIoTEdV4eWWQoFJdGf9OKuDgoY
srTiCANJOd9SVPfe+y0d748x1AplzTXmbRL42MHpRNoECMMVTx3F7AhYZcAw0xTa
V7JYtQuDL26dHZazJ0sy6Vw0QKboPT8HV3Q5VifE9BvBOEWKrffslLUlPiTe2hyk
c5MZmV8DkbCQNk83P2bFaXzEyMabPdmnbglJU+0Z/zCihP2OEz5pc/A5r1fm8Aw2
+TZe57XbUPmaFhSBNi92ifybnyGn9iLyH1adZdRQ466EgcaI/Tlk8dDxvI+xJDi7
EUpK+3StUdQvNau4dcHuP6auI8ufoYfYyNKArCLiZBQHZylomEPcCAeqscJwTeUM
M+w9KH1kbUeh7jdfEuub1sSSNRll6jMLNzamN435l/CFFKmggjL7V7SfAgBNwj8m
kvb/mFGK63UAlvdILO4Z46y17B9Ln2Lii7J0hoaPTH/lsDPZRWXuTSO8fwhzFEkC
XfdM7AEV+HpTvsSjk99iu5wWKDM7DCRe6BHajpIWmXL7MSo6vi3VpPi2bRmgXOV0
EnWF8BdSbosufce11HMaB+AOmfW13hxNvubQ4J0IqMjur+8JKLwIbVqOMBv9BygF
QDOTOIFT00caX1qWcScLoFC84Tw72yAfRIUNCPhDLiY9U0fpbadX7RPIRmNEzbje
G4MKCCZ+Zjgs5kAajl5/27VUNGpwOt4I77U7lQjN+TMirFSMi1MgQbByYEnwVSdC
sAFdAUNGQ1CDsBW5hFnr024/XIvfGJ34ODaZFiqwJhTgliJjUi6EyAh/GW0lqaus
M7Z9nu2Wl5TEhqsFsa8Ak/y5ACNmJ/VjLggKy9FSMtAxCY+lxTRuwVjkQPmMIU79
ao9QsnCF568ZbViGtcxdfkbYT03fGDDTxmYgSw3+er847k7ihyJ9PpbnycBqlSBN
uBiTJUc8z+GbW5iDliJybEQHwvzsdSsUAMuywXejNSiocwob0ldthXNGV+tsYXqS
YlBdD2C0/sSW7L+wsubgln3nX2bdgtrGgtyHWElgFpvdeTXbsutY3dXaq4Zf1r3T
qSTa/KJ9veIMu/BFJSaqN0pI8wF5LOE2cLTPszbr1Y+U6uokobyYMKzss3aEqcun
eCzpGhvLBBCXCVv0eV5bgSSxwyGmhE4JXcJkz6VVkFrVZ7aHcJCvEs+jsEhNdxEM
R3LL120yRhDopszueNd4C8lhOEgK6zfYokU+9U6s3RMBHfOPFCUZE9HyPiSRUHlc
SO5lyfoASZFnU5FLtzZKNqHi60zM3ZiFMoThrMxVLvz+hZ7arCffRTiG/HJjY4qE
BbTHoz579zW/z80vmtPTQs2rKJ63JSiXehxkuLiJTihMFX6J+IJkYoK51Shk/8BH
Sm3JaUoebUWrFPCzmpEQzNmGzf0Tey9rmHLJEOMIH5h2JPp4LthQplnRatBlxZci
HBK3kTSDDkelw0jeswA3dLknN4UeqQiIsX8QPpdT24nGw1U3sKE+wVsNJmWN1/y5
vaIUzVtS1Ea+SOFTgEbmugTELQ8nqQ5VYquKn8u7uNI0ohlvkCW4pIhCKAwFfOC/
jkGVdHwJicgsB6fI5LjoL2ppE9eVlNVLejJGdaGE/o72XG77w8l1GhAEo9IUwfvP
S0Cp0KwkIiPoD0ds9+1YWxVlGeN2cHAwV61PTCOQZK8QsO7bh4+8U2gsj9+30ZHy
vqTT8vJxYcDzqDLFnlU8dr8+5x09oELHGr/zqgWKU60P19IDIm0tKb6f35wvWA3I
943mR4+XLbqvdeYbADh/NTXH6AcZBEB2TQJu81/yECzdlFKJTgH8mprkRlACKmNd
DcTafxjgP4Sjfh9Z+NfaBzE80b79oeE6+9vVkCkNGjusd6jRg9/1TZ8RgTHOTCyK
I93aG+p0AO/hzWoE0KPFDFXb+NbaYnSdG4gOtjqNW9hFa1ROqf2ihIXPBmE1SUCH
MgZ/IOI+bPYaC7bTfr151OOl4hsfjeth8Jj6HUwXYUI96YV8Wz/oof7ogmBSqzQ+
RlgWxtdJfh+A3MqV4AsuaqNlY5GZaH7kkxcTSl1uXBoFggtsvWoUuhJK2OR5pX3R
FLI5ZGAqtVifXwvpOP7Byq/hmEz1dbsaccCP5OEhmx15Ews35eJx2x0UeO3PWFYD
PiZ48fiSFhJf8PNBifANEj4k9HYLf+cUQbRM7ktZjuQuzgzNequE4+tiqPh/2b4K
qd8migFx2N7OrMyDU+O3u8Lyh32DiYirhubG97SxtBi1ruC3tu9wp/1vNmOKmmmF
po2BtpqXNHtVF6WBqky2iJEZuqwYmubJWYID+F1NgtvO5zc/4alDb+rbS9Cd57Ur
ryM9ViUTnXe7x5S7BUQ6t8whLaWotyJhn1S7Ga1Jje2BWWbHSIW7hZCCLZSN3o31
z69x+KoTWeKtEzvqNNOHbpRLcDPQArnSJ+Xng7GcKEytPNftQsPcaomZpNuurAmR
YQk6XsZ85F6twihWOb3cpZnNiW+QJYBjBUzEoDWyctceJWvatFcxLG5OkG51kjhv
aWwW1n/9ZfUBJzhhOEGsh6gZa/NQVa+naV3pcLI02uKdXQMWbamCSLIsGTxxGScr
n1GVP6cpMcEXtJwkBxsDfU2JGKx4ih5nNdxumIhA0HBa2rFGWVeXxMH6r6ILF2Vo
QquEIJ0NBAZ4ZHB48pNtlGIlkQX9Hi/R7fk5mjzPxI/qNxlEdDV3ABUbuP41wx9O
NBpOAqt/JqOuQShTWsX0F7DTtMV0CoP6rWp8OtXts31cJjiWx5Vliu+pnnqA4gpb
Sz0GIugIkDG/09y/anvuSBHxFW8q0D1E+k43kZ9ahrXowTxoTd3bh+l+AkOb7X9O
Bm03Fi/RYHUAEc6mdtQh1TUz8T7YD0FAfHQtsT21ruE/C0dxtJSO8sfnqzv8egR8
b3WGkwsV3tlz17t0kfthovdUop9kL3KtQs/lvFiooqb2UrXeiVWiOzPNfBFmOU75
WrDWdDhFkhN0/ZEeWTmLBfXs8n4u8BTgYrKHOK02ey5A3rqtVE50hGLn0rHNJeQl
Z/6m9ZEXJxVFVQu00wymjISeZr1O9HHNHaHldg++OQXravIUVOnK+Y7ShUXTg/la
nAb/tVw6987vn5UoAzPmgbLIBQYWOmjr/GseKXL6UjWA5FU/TMuwGwUaHZINSnB0
8sMAboioQ+lrpgOgciuDhhO1uJJMOMf8PyG183l/fgu9ratgGNDBpmWu5da83dMa
f0NCqeX+hZCgF7bHimYWSxNNet+Q6QB2hS9u7oz+/ZSkP5T74B9FASYK953BtsLJ
+PJsa70ZqkrrCXzfqqSjpsTK782ohBCIpjPTZIwTGMqI7MnHLC4AC8oRGthsh7We
dVhtRhife6etw5aSIukb7sQqLTouL4tI2StWAfM8L02CXCjjTf/htPT0Bu/zuRn5
pVHii6BBp51CI5XJ4UgOU1YJMs/0In6x2J2crMXwzdyurWy9CfJYY5DZ2OS1c3VE
L1nLiuFa1A50m1AqcHhmNwhpjZQ0E8rl23t78FDoGXsIBOreVoqyprkW7UNt/zUf
cvGWEaOp/CY6WuIW6HXA4Ys+GCdVe2tOmv87r65bZoxI1avYXOosIXhnv3wWYaNn
boJh3RpNejiIuLJ7oBcZqBltYy/OeHyMEMiaE7QThtlDxFOYUW2ajIWuQdFpwTKb
JyNKysc/DlzlpUiLibHRQH1J4OajIn8TiJF1ZjRP/Lyq8C8es768vZBuetaijtou
yEdpnnzqtjcXxHPPTjg4ngjPIOqaB7HRr9kfnzoYTM1zfqjSnZK+yrK/Jp49RY8S
bvu26ORF+HkeY0Z2kL7EFaLoDHSnniJ9UQJTvMEdP2KolNw+H3Iet6PgCawlxW3R
ESzqXKYP0wD21Hvt+DBI0AodADvc+He4HHSze3UVkbfvBwoG0x1+9Jompzi5AEZP
OCjhbyH6ui2kUdNic9bfaOIaMEn/N8HLnVhxYpUXJXZ19crQnFTtl4nzF/TI7n5t
1lxbEqH4fRyGLPWz2irU/cXLDMuImI9pQftz/RTzRtA5+sn7x6NiAHyX0P/pl+ul
MfQlpDri1q7nXm++LiCIO45KgDuczZznzR18mhXjxxNS4HBTC+Q+JG+ct0NsZ7fv
/OSi9F0OuRZyGcgtTdv3mtuKj/VDtYLUlYpzBayPkAzcesXmsErVwQ8D9Pof4+BC
xkO+b1nm139gmsaNbHEusP4/06yD/qhj2uV04gbFH5tcQXWIdNrKaPqScOh4ZTGN
6BG4faVmEJsQ5F7qtHLIyB3a1xWPBDMDI2KxBSl5vPYsQyPCscHGOv/TATbpWAgb
2S/tcNuIMG5fSxrUQf1OO3DMrLrjg9ljAZE5zDk7HLA56GIWLQvvG3tNa9Gpj3pd
hbfjRjWoVklY07G4RWJNUnKgFxBqKqZ8jdqXuT32f7ECaCPMMbBlg/cJe0V2F3Ez
wyA1rnkQtzOTzkFwKxtG5afgCpnvgFfLAgZPB5tcxJ8LfjPNVSF/Pq0+7BAJIjBl
DNc9NOMqjEMg/yVlFzYOlN3To/LB2iAXoFZcVt/bBW2/3GNv2Y0jomtxZ2WdvGpp
8Q5QjwsciGuGcbUnpajSPCZuH7/s/43w6Z8XBhIGl7tnzw3yfCySHhuGQdMScRyZ
HOHYGclzN2HN8IkMT8cd5ixYwCOgR/6Blz0Y/8Gt0oixbwCXDob7dWdkoR4tZ0yG
QZS1w9pjcwrOxQpAcc86vFoiQ1CTsDJxxy+WvcoX8LfQlyW+EsxBJl6PwQVw1iuN
uZxkDOzu12htrxFzEM6c5Q1HH98JjlefpXGftpDJHCXDj2vvHY6XQgjYRkD9E+gz
sjQvp/aszjMy6vtiuR3OWLXTqWYjeUcAY643jvex1kohPAx4O4QCKoVyOHct3FFo
AkLa2NhDnS2poWRmGgu8ZDdV7TvAISZjD7a7PmVAXHwdCaxO7BOjULStHl54T+YD
cK97y07zmOktD5NuEJPkmdnJlsDm7tmz5Mr3BS2/Jc/tUbTpIWifsVLa4wj3lWQk
siLsQcbvHHTII5Z2l0fwJbpGlYJgRO1LK16uKIF6B30SxXvIfQl2FQr251iLIZl9
2q0APJy47KwWAwgNzWk6j1kQJ/+nVvsMLZ9HqLcMZW/FddFlK7wFoEJU3fSVXXNM
WDYkiV1/d6+8OWhv+BrS/gsSejxRfCAzrzGBJWaSPK4SzcgaQffvsEAlo9jPYoQk
MsJ/Tol9/oh95EoxSc7tCVOCfk45zcA1ADybG3qrybxYdEA8I6TBJJpPdwQrIhDD
sG+aDE/wvV4qCdhXVfJB1mFp7H2sXsf7LzpA6b2W26PfHx6RuH+x3+O5d4FICyy7
MWDXfU/tajkdFjf25RNiTXKq3rtpuGW3IEow/j5/ImImTmGm7+h+ArIbavN9iENr
49DYEkuy9xwcvCBv2sE3innkuJMLVRKawQLaMHtrb69kiZoZqOFcf5hKZBu9zgSA
XseQ8jH1siTm+m8RnIjkFmpAIJd/jp9MFqiJV5xBJXLjoniEVg+9rs5lJiZMEF9n
9l58bcivZOm7PZ+CDE48MoWF0j6GS6tgmi+HXQlIgYdb4fI6EB39mM8Qfygh296V
bIdnY19WDvM6czmO5vXmlSdDkhvso9MUkNPzqn607zWLV6QxWpGEEHawNBNF23wz
ManMYT9A+9g2xmtFoAn/BTbSXAetFM8zOXlfG6kynet2Xr1pq1xqn7W3twf1wQTF
UqA80EjZxgkquUdqUAgmfZ2wRo646zt/q+kva7UekrmAn0/r4p2n0eL9IawfwFu/
hzRbkddyXEKyw1Dd6Peig1SyWzibhsTO+7HKl+kcM9oVPcvownCwdbZcuJOoVeZd
Q42JZHGqMcmveuhUxzBSNfcKkS4TxPC0+wG6Ua06MjX3Y8ZVz5vNHs58VOxhDjHs
ECx6S4dcbIqyX/rvI/qRrSQPwNWeL+lkWyLbcQSr+G10VGr/pCiv7UVER/Skn4Z5
3wrHBQyE80+G3ln0/1LDZYMsi0PqEkOCUTkslrq3+9za3g6iJc2NKvg/3MJaCvg1
AzZYG09aIJvTpsjXM3wAPrHH2b0mRit/46rjgexzQm4nHXLspw1kmNwxNsvjlyEw
5B0nQFkjNNZ3Z0gezd939BuIaLJVQ4wRu4htbImm6yaMgY2Tx9IXb8/BiGqnp1eR
uuE22lrBMLMuDZt+c6guADhkhggwRyyIqisvpUb6ssoXiLRFGJahrndQFypnmvUB
fGWRXQOcYtuoiWj753ne/WMgHagrSiVO8jPdA58HDJloRE/OZdJ8GO8Xv+hPmOwV
kflm+rOuzhwyT8DTM/pIqz3mms+IswsyxJ15FjcUy/sOiXvcKBvURnYefIJYM0yi
j+C7ZfPVKu5XFaiz/d3I4ZP6q2mGVn+43sBM7yyjWDM7ojlZca+NMzqwIPoZ2I2b
62zIXNrT44dhsTNuKQnJNAKHZzDXQyc++rEP6VJmrT2Yh1330PW9x6YB4cifaiKH
21XD00bodQw3RyXxzIQkw4yI3rCWQzOHXRpJLuqA7HAkpGUclAT/I5Rod5Idh7XO
aBKfgeLy5kzIsuIH9K3rYSuBctsrYibgEpPR22Lh9BKvFCWZdkMrCnGPSmBTNY+F
LXEZgLeTW8MJGyAx27J940Qiyhm6M1lUwgQZcAX/MPdr9PWARm8RxMglXcjS2DOE
XS9GCxvzcfR9psEJ4e2ZSVFjLpYz/q6yDsL3M2na5/F+4yfC0tSwjJwnptM5yjRJ
h51qvFto81HDX/eXjnQ3lgzybEPXMlelCI/ZL5xfn/hB0V88C449McEyIjeMrglJ
eQYRYTyzeoNEYuu57RifK63kJfWF2kbtdgI6BUORuJpIHd9Fj17Z6htQP0RaqAnl
2IletHfrdbm8Fb7w7N+ERaduJ7jsxGWY9LClcWXoSBz++I9k2rwlCudAPDy7NUOV
+l2ZqQP3wUNINPyX3EAy/hQQtpkVtxB+zq3MkPsudpKUje89H1RvnqkLj5jVVrC4
wzdidJwy+nt1ypKmpPdylj6yt63gBIDuIgZPlkHswFSh7CqOSXvsjoAfkJRpt+Xl
kjGxbgNYZbHM6A013N3p6P/beAwzz24RBk+as+ytF+0a9T4H5P92eX41xHQdwfsa
75RoIpCilfIbNzJ/xD8pZwvuyE4cAuzD4a2P1NnLu0Z6rwUgB55rYhM1itawiEPJ
GMO3NeiToO7YNeWJUuCdVsdpFlUIaeEo4mWlaT9euALh3iY7KDXMappPJ7S94rH0
PIGW4yqU5dlkqoiuRgYe+/OxkO2YjrFrjgNWO4GLmkWhXFPw1bjLYDIpSQ65zHWj
COgfgwjIKlO7oR0XgseUJ6mlb0iVatADz5H8rYfRQTYZJw4Wh9nVChO/Bdz863WI
ThUHt0RhFmjk7+VySt1yd1evuRoUg4Fr/BD5TSkK1vRvpGty7A/gZyAGYKFVzWFn
YLDCh+7iGSj7MNNn312eMqf4tY3i7nQd9kPxPW5jUXY6BCWn86kv90ELghN6nbOs
30vHUuubc2cQGQFSajYe9TDdmiXPvh0UlAm/YC8mQPaG7Dw1FUkj9zwonGXpHLWQ
xp4GYqf78f5ymkRSa7MBhSVtNoKAhBcdqJmkGUSFDP+IbzqlncCd4pLBxPG6sNge
nn2RYMr9PM24w5akVpIGGppJ7Rfl99k+nXJO6KthKD7se2dDdB+Fh4r4TScTuCxg
AwBZd6qhbSsfMf7WW71fJGZ9jLWPoEWF9NDuVUFTcv33Kh2EzY4oZ3TJkOAbdaT4
og3juWvap2LAa/Oa36qewW3xnJi0MoX+3JjejqCFADsyMlY/gwbPrZO2IMFKoMyl
shUIMd8OSw39m5mDwMkjKnirKnnPKH2qimTmbhqBaxpN+mvKYDLtH4OtQ79ktC34
D9mOjSMnLmrQmr3ClHiW5S8LN4dhQ6bsncMDt9WxmxQMS2ValPzpBfNp9LCiiSae
Pe24669ebWBqsArM9TBIJEOpXy3hzOiz92bMKT4xmv4WoVk5sUCKCk7Fn2mY2PYX
QBRD+QdDuJ5iJre8G5kiRVFn887PbK4FJSdaecjV31LBw7yJN8bg6H+sfrZBdUNy
z8XPnMNA6BPh2mtFRyZN3hrJTdC56w4hTaKiTQi9x90nW5GYOULM/V6jU4jGOCXS
y+ozspZb2hB7JAVYK+ZTPHVIX8fhXcWfNabCYgMBAFgiqKISeZwH0nZbuUpg2ZTL
ADCvY2Y0dba1bsaaCyPQf6QhYx8o2EG0wEd5lXJSGy/vJXLnSS4S3B5ESUiViZsq
D5V/CyVBumo0G0yMTYXjdHXB03fjLthPa0Uw7zrT46d3fVwhpoVoyKtI7yFKfkVR
DDyWh+ZsmpDaQEB+ZU2fUBdF7Oexh4LucYzibA07PFdCEfT1UDU3IsQVkQLdZhct
3PVd2UHa5rrrRG4kTzAN4OY3CZb9yiDWAuRjaaWa715LrWxF51YhInfRSMGfx5Lt
lj3ZXXU3DGnxE23sVGfPSsQAwU1B7fN9dmCj4BnWCv60PVKl6TZDwhHtOQ2IAfbf
V0plL/yh+XoencrVNiELKmX9SN1/hCqgB3Cb6w85a4w3SyDLa72ZEaijJDB35s7V
dLkHDewLrPV5KE1pz/JCF57U+VIhBabSwPua/lxI5Ohwao/W2+4l6Uz1GbBRyDJX
cPZUxbEvnULGy6TbsiFy10N/Pb78z6Ovc0NikrogikOUcBLo7vIp6rXaCOEqHSoZ
RRxd/iB4ScuGrzcbSy5ImE8RZHFxUD/UE/3dkTntp+nrMjSLYIebqz8u0M6TPEhH
p4weJ3WoV2+K2fk75I9ykalT/OeVoXYUjtG8h0K1yf4eU+vvqQURcRwT33BHAhTt
aWwLc4RYLrpTem8uswWD54mQM+82yjxhn2qaWuEkzDF7UlEh+NVbH0YUaeoOAswY
nFrhNtiGk4du1qSYBC3MpYXBTSBMIWzOju713bYQ2VPZ6AX7OGN3s0WgvtWEFxy+
OarWekRA8/wEdF6BISq6CpLUArtGvtrV1ikxZsupwWkIiBc0GYvQbcx+kKpxR1zO
rQBEc7nWyKEbRVDLsobu880ynChqC9WObYBao84m3heVmsdriq88ZcB5pMcvK5dT
7uPaWBqWA0wSoOGv9hK/YVpUpoYUB10egjS5+oGAX9oQ2GdBm6I7lAk5sLzXVs0C
RMgxnx30dEeZGTLkj7MngoauE5KVS3ZIhIIh6qXS6eFFklrdhFxoL69MWDGr/6RH
R2MENkTr6dS9rf0E+2glU61zUJsTDpT3j0HQ2pSXqnFoJTKXCJd441kRRhXjg4R3
fv/Wsyi8NcyCpQqAhu/g42VL8o5CPIqYhUvcEKl6fXOT3euvdagYlGIfbG6SAXfK
qOSHANWH1r0sYlBH9aJxD+TLLyHkH7RbZArNwYulHNELXO7BvqXb374sOlwvcZyf
w8Y7GMUbC9/BYAxi78YlKUqZw7nFVrMO0l5DATq6ZGzl8lcZ6v2z6b4+ABA9ig9L
gFTpEnGiIaR3yWpIRvUtUo4l+nJVLnx7NeSJlslcIWhHze2+Sy3i9cxqcAfpmJIo
bpgG5Qsq8cOMijJ+FGtkVAiBR+n8leVwY4w/DueE0T+aIQKregdecLmfXQG4CJ5R
cv9HvCl6bMbvs+USLlsc8AyZKK+aSOoNR94oZuacD6Fcl1YBTvwYx+BpJmAFZiMW
0YeqPXm53ROOT435FBzevKahclVh1cqeeCYSR/AWd58EAY0jpOM/YTeXjEr9njlp
555klcNlOxGywtBK7YF2s4s/lAzM47oG44XMtA/KSx5YjyHD/XgQZIQtfGPn3im2
gn8Vgj0ukn3+rHLzUw9l6WTevSeb9yvfJMX5kSuDv5E16Qr5DvAIeKOecEyFm0rK
36VOlKGKjR2V9zoig1UV9GOEs4TqhCv5BnsF/AapnGDA93OIZgjH1vmCs1EYYfND
HqkgIXzZwu6gH7x12njJ5LKpGDNnnNa6E9PcKB3i5s9L0nYL+cEPFAGqjg/2Jf4o
HGX6SPonYc0udV4f1pitt5moEvTq4Fj7I0liRhPs8HDKjf7q+XbpX/skMsVbNX5P
aVwVULGeoyV+t0fkZVEG17RZkvdzJ0uwPaO0bO5R7kqg6wRkeI/cXOPHYMsIyjrS
/SX5iseL+dM83cuT3t6zDu4vqfU4CaF9f2IUA0dNpETXyX7fPPJCXqRMlJEAkhXW
6Qd775efyraOvlvtBrWE7EMfhMMS1+Mnq9FsFJTABJFPgQVXE9Yux7MCL0ILka8L
eP0SVe8tctsW8prGUgRNiOubvic8+A79mqIFYkkhWMTqTUKAfUsngLoWOZS7dqlL
b8o3I8wJ0uQNaptPxNRLOiKgs0XYz65Ld+DBO1H9bPlR34APh6gdFH6CcSjDxmra
FdCqTNTxcliSgsuaL2o0QuE/DiFZgs+cMnirX2j35zVf4T/fk99+hHZ2nvGVFss3
MOxpN8bwBPcpUwzB758oGpk8SM5HOrUe2nKKaBPgamYmcty0AMIb5Y2MkKT0DEc+
spsUSeGHGwumuVuJs9sKL6kkrkVK/HNNzFw6V5DxZSusIUVWpF6eO7uKnTtIMRuz
ZdGaIiB/OxxgSvj+b7CSRXHpek0fJAsaDnFIgb/iUzmY9XJAfpnOkchCQUseDMwq
ZAfBIV7eHP0C4Xl1taS+XRjtwSyVulhFs9tLqK5yQPWvmI4b63qbW+xPkINhZMa4
J056HWmu71yUUNy2X+yJ8l0GhQ9b/dMobGl5cY4Zqfg6z3jnD39FQbliKiTlHS09
+RKl/pWdQIc5GTd/jWHil/wGg3WALNZupilEcKIz+osgIL6DktMMP7R/+pg+L38n
wOA1AO86DyW/iLFZvix/ePk5wcBMKNvytM/0dFc4/Qxu/tx2aUxVIz+MD8cxWYzE
cf32LPPlfmcqkbmsC3fVCgvhEy4BZsixhGsu7JgNtvei/YDL+DInfeP5Gb0ooHZo
9f1Aa1LuIFs0GZIk9kginVarR4wYdIr2/HXwe88/iBCelyhvzMxwuuUGLba4htYM
ffmnKquxrwXvaQ0FJpR9AciflDau+VxyDKpYVoNdV9n0gxDTsNyMpB2b/4Y3pu2A
A4h79f9u8M2a0J38dkrYrpal2QAbnIgn4gcnqR0xHPpe6FEkskxylbu+Jbewp0KE
D7EnDjL4DIgQRaTk5w3cgE58iHLjXpupEOy3NhXNVLvXEltcBxYS8VL/im7Vzqyz
LuYAcOnvvpGFdYByRWTCSTHEnUwK8BtHGiMv9gM0nlqTRH6fdX7IT91xcupDS034
BGFSLgnlgaerdOM54l7YFCV/vAONb2xOlTQfCt705Tas1vjpZrfEZ4KMBTvfpFOg
b58mq2YX+yTKcfa6Ikue12mqP+qf4F8gGcZnbHcObGQok3e8IkwREZYFvPRHgPoG
Z7/9uycxxmTD0gZ6Zp3r9CBlBrCjhL5lI4Z0Y74oCa7SGShI2eMyeHESaLOv+VOW
jAXXRd0VYXHxMYVOp6dbgi7abp459ndsjjff3hfmTdXZEzJE/xX6V3qQTW8rW0Du
E0PPuysA4n9L7cRBMIFw2GGLWWyEcFdO1spV4/je0MKg2w4rgJK4SpnUtO3IGa+o
nVrC9xBx6uSm7h2TZWVnV/7Mg6uRf3WVBTAFxCZ+72hYoWJtdfw1WFzo13cQqdDF
Uh5RGF/lqpWul7HeWTwxIM3l/jZc4U64AeUBAoBuEXMQm51M9Y3RXaNTY+2Lamyx
JRAhHEbxmlZOESXwPw7/3Oq0ClBSde7TG/aUPB/4vVVoFqA08ebjGfpNJlsP9vKu
38m4oFY3VrdOFpQ0mtMllEvNygMDuon9owDZAXcMaIdaXQq1ftmFh5Ag2q2uvvl3
Ujf9mzpIXKtd+8iM3FaJE+gWC2z2/99xNGAaw2vHHPLkxCL1Sxp1eTJ9s0BANrla
18QmJ5WfVtuhvh4hqEDqYB0jSMQQNepRvCsenVZOlyId401odSrKxwgVfdmltCv+
CeMpv/P5RQebbh5Vd56Ft+v+hMjicR5lzEtXOlRin9OmB3gc4x1AhXny81fy7ioV
BHUqvFd7WmtStuSngQxK6uHWTlrk/TxMl2Hz/GChw5vwih9awkN2gyfHCyTIdMBC
n4Rj9FRRGPnKiLQWgIlJ67M2FbZ11LverVh/uHpkT1ei0C/lPLg1/srRnYwzPUT4
SgRd9jU1eaguNKv84qsStMU8DpgHp+I+W7wrxxTcu6Ge94MEquac6aPYB/tjheme
oTP6DOQJjPkImnYp6rJQD736L0X0UOwQ8Ch19ZSUEUiDuc8paDcoml0NaB2MVqBH
jcIK0/nkCxnK5HTiERA+T1mnKl3SVeLmXhMHW58Wl93XOBTayqM2jmljq0/PDu/2
HC1tH7QiAQ2Rk1QoVjK/2K6+NexKeKsY8mwAMyFunjoAqMeqHk805aQ6by37p4yW
40zEWTu/Ox/Ha4bjbUhaxQpqf+XNRF4US3Q8OTQyHGDEhA1Z2kAmT4tSPc5sdsJQ
osw4E3/RIuCr8X5jWLqi1XJXxUVslIi7FbY2fCl0nbGm7LOeNu2eVehBmbkAdb40
WfZIGpg3YJLe10Sl0uIRDBDKHSWlnepoXetWpRNZk0yH0Uoc1YobElVSkqJBJwYr
bDhC15uCHFncWm4SltKuGEiaAUuZR9h2t7OEL7urbWh1m0oJXi5Km/WkVgdSIIgC
Zs9zhIAQTgqpnnC7jufpflDX0X2c3KCXC50I8+YDCtOKyCKmfw/9QtuetN9DSKaP
aBUewFKS3L9f9hQKr242Njl68ntNpkKN+PnaEwGKxKv3Jdgu/drvJB44DoQdIEM2
KQcejp6TFqYqMkjVd9GDBQCWLH61HRHB5PnZTsv/+lhlErZFS/+MXmuWM6gRoyMC
57cuy6F89mzfeu9qUbXncKYfq5lLrilelXOwCeV1KBpvyKpIEPUEX/PgHS+I5eCD
bHV3cT3EqkhZ7xEV7sf5qDM0ZOS+3rChXkTLDNZjsQBSKXw6ocuA3RV6fugKbc31
Iet61ucWRw71P8FCA5fph7GiZ3Q8OqmfJPXckUogBMTyfItujNAYtcMhcMjKNqkn
3kgTD07OLTxAZr6AiglA98Z9ZYEovFZNPG4vULVqgXSOMcFQVeEahILqlPH2IfXH
Sy+xVcO3+otm2IF/hbxcFgrVvFRlSqTfl7HUDoWRa7VkaeB71GppiPDGqEdkambG
IXdR3VlKukZX3PNm6rCoVsCeXZmVwGvTuRq5bjJ0DXwKE6PDOS27ymvz0hhAVD/m
rSUZ0an8pqIpXlF/PuejBH0TE4GziN0RIuQABZsXsPOqCp9uZvFtzAzTXJuUb6o0
qO9cTzMMca7LR/BkFNe86enHb/4ZJkb5SMvi9wpwA0jueK7fmGT5pGYlCD3Zjhnp
5+w6LMOs6bh/qS8EdIBxviuN5SQLRmDjJKijMZ9pcsTIF13Cqj1g0SRHbWfEFozY
XMj6/vTUG4BnmJeq3v2tsXbl6/mg+cfb6pFBo0cbcZTzjAyUq292jZNu9yWM/ntV
bfVGZ07aPGSFGCVGAd80ZtwZqa5x6Xdm3uq9K5w9x2vwROH7kLrbWRJeVoSUwdxX
D1sCIuXWWIOYFHZlWoMckyu/nvxEk4Rmzps6TtHGDwgnbVxa637A1QM0+ZoVBqTC
XsyPIK0/IYHQvcQxrPd6SrvSsCNqmaUvaRmHguP25fxMUE2JhfJwZ8eIhHa9hUbc
nwZxcNR4aC12r/0ttFt75uwwM3gEIs0LjLKQpMWr9tReCODop1cmh9oOOLt6HDyO
M64l3WXJZ8nnJv+Yb27IYfohkXFJr9bhxA8inAoa0fxpLhzOEjOuTA4zY/2kmuUJ
MA6aRb0h9yVkfZM9VWbFyhdkQFaOqw79sPrjRaVO/ZqJW8uVcLliyArMu99eoXM4
L98tzfx2iaXqn+c8jtGi3W0idpxoKqtIO/KhnTxLIqn1MhLaufuXLGG7qTaH3Rwv
mqHzOdFyUufyP9cO8sluMpGTpbFRNsBz+VNn6NAmA4sQ8RCVVJct/ridbWV1k6Ll
DiktYnCVb/7op/5ZJphzpNkAMW0B6tSAyeQwBzJkdz6oPmut/fDsmk9spw08wgmc
UAfXuLJf1vb32sROQGxV5EShQQEwChkcMTdSAre1SELK7Wi7k8uwPlUyoRYURHkj
/dhcQmGa0SG8th5kQnxd9C5PY6dx0uwPh+4IGq8ra+JOKQvqimdk5DoFHEr//E4O
68/WLUIHcuYoYMVoPmZDsnZIXdYCAkGR1y4cwuJLYULhYtd3p7hDKmIPhSEz9Gtm
YnGE+uUfNC+KDhmLfshPKt6wwVu7g6JCKz2vidToeFnRGSj9oo8DOtkKN0UAHWGu
9UJBKkRy6aKCNG53E9+cRJDwQShAXSd63RzEMvRUy4sVbyMOyxHAjz6/ZKTKwp1F
cS3c77EfmIKm3RQvT0cVAgMG9BUFNs1/RDfLE4y4K+1BVovDlik3dAIkP2UXcQIe
j7Sl0eJJvDeqiaAo7SYPWQfLVPnvbnF/oFnHJXE3zo5RbJdyWVsQMOuRdSvtPxhX
aVU41j6VqfqoGZNLDO+2aoqD4AccJbMQ44mLXk//1IVgDY7iK+0PngxWaEoVSP+K
2YgSC1gJTuq+h9b34wCRlCwg3uTPCEuctgk3qS/Vx9xcr+0Lprpc4+4a4l+2tE2J
qk39xArqrrC5dUStB2/rTzXAVC6+jk3eoYXJZy1+hKQ/FeXBHiYVmWr2Z1DSYZhc
/FqPkWcn0j6Fd0xXhNzsbPJDjEcC6MX+dSNipX4x97aO9T6RBsYjMoTzjrWvg5BP
u1ngtPCZAqhyvT8KR+SjPbH788g1Kdn4oKARFCTYz71Pt4w234CO3HDScy+MriHy
sIwBe81ieLdIlse0wf6ViJi5+khGClamTJp+ZFUXKC0OFgJAy5ikNZYWmhw7f2Af
de4WwPqmVpiNZHFpAiXyjgO6AGSxsWUreXW8TyF+AX9CZ+EP5lcgd4s3AaBh20Iu
WyzncyAg+UbFx/dHF4oRr+K+j/2Oi+1DgS/UkCzjRZVmPAqIiFqUE+QFObv2jY1N
8d9YAEL+RV3oD2Nbc5ziHJO/rPSRrRt5RqrBqM2xC7K9BNhtEBnZ6lwBToJk86Oz
Xqtpkkl9/WSb8cXITklPIQTHrR8TweF56mDgrngx3YdiMpOUIcmQHkj/QtZ743Af
si6iw/zV1+vnOQsME9YbF6jfrgBya8tFpXk0TFpf679sR+JG3UhxA36BodC//kky
vVef+k8gWn+UXDmNtV3rWmNTaQCc9J/qM9YhjZlIzZEo1KFyT3lMlhn/UMEowCny
T7BNkbF9f3F7FXhdSUvKdGx9gs4OArhUyOMNOKUtiFP9sPIINYcr3NY9eVpy/q+9
8iUb6VtvaH8rlFvGW/DqHBK6IroQYPfsBcxOxlZdaSQhnrxRMd+5C6fh4ALZfhch
xNlFm2XLe0plz+rxWL2J3cDz7Mkzckhd0LTmOAK7EduOLPDa11h6py0UBY/82yjq
gR0Eqd5cK8SbJEtYhvNFRvrZdTP55V+iCSjTm62EiuEZ+GNv9WNdPJNjwm5Tg0fk
7U/+JZMrthZUkOghshSpfqP4qmqK3d4iN68rVNLz1AvawnhCyh+N5biD2Pzk5fic
bxIx/xPx9WYvvxHeLr417MiKUvKIlNt3wfiu8Q6MDL9cEU5DXyu+aOOmcEn7BbVF
mR8Vkphwhsrh1DdlZrNgJHfh+C4OryxjPaGFFVe2v5Nykp7ULTEr03LTKfM6McDh
GwFJ6yTCCG5RJkvolgMr4CLua/kj/WDlL5rFmZ26s7UMnXhX1+QPlh+fMlL5IbsS
DVAA2ay49JbCASfriIxTHzQVxgF3Eemy+bjCTorePbdBy4ahHsNl9HvwvXra6JTu
S9YsHDeRPhQnoy1Blm+g/hreKf4ZC3+P/ju0Ui0BxZtAYRpEQJjLLF818c6YEEN3
1uKfJ2raoYGwtikK3hmZMOgqCC+vzM/dyiDFPkm3q4gUQm3WNiHUroLNcwMsWUiI
rUDs5UOecdJwyGZnh/ezRrOB8pYP12JqEY04jle01c/1nP2JKhFUCXhYe3QyOONl
3lKJEKHePb6Yjmhe9gpuyZwL3llSKBYQFrIMr/5toUL+qdJ05DeqwMdc6gJd/Fv/
cQu89RgOcPDiTtiH5XHzQU9dS+CvVC9uAgXfLxwFFCaaTKxsWL/oAr7mtiMlq4uc
GSMxxfhJjHo0sZw2zWeOGv0tgjDuuSQBtvzeeD1NARprACrDFIi+MMEn3EytQubm
F1JIgHXdhwIxbn8fR8oummJrL0IpIvF9Mi4zqGDW84/68D2XpuiUJeiYC+mToO6y
V+Vczj4VrODVRVLdPwIaOBKSlBycZmV7VS5mSSrUZSG8MIdnTVOUjiRJBopLIhYa
zhRdixCxnmI1e5gRqsteEEl5pRJ6ZVsiOpFxEXvsb4d8IsmiGemMHZ76zbQSlp4w
WlVo0JN56549RuX6kOB1y41FBu6i1kGda0P3gh2Ampg9rlKWJB8rvrZ/320iQO2Q
IqEu/f/YHvoF2dMgfkF05UR8ri2GLxmQ0ZOVNW2OkODBaOpMqBpc0KtWZlo5PVE2
6uUcawPhQ6swyQLhngabUeM7FDBeCStSxOmT+o78mbwrXS0cIpIfhb7mrEp2SwTK
/DJFEtu4KoTvWWOc2mbnO7zpNppurpRCXmjUzGzT7e5raYSWCZPr7vMm7ONL1j4f
/X7ZAcQww0BqOEBu3eVY3G8duFtb5Sohu5GQhWQDDhEscACEhb/5A4xMFJBq7hmY
iCYv15w77LpK38rFlWFNY/ivmSyMyhUrGQdoBRr4wxcYnI9r6A+sljE0hSd0wRMi
Q0u/OsZKYMItuVcQzo9o81pYYdIl/E8hMBTc/2p/YoUOlX6xcqJ3k+XyqN01Q9e8
9eVXjTqM1xiTWT1pcYVRShIoM2pQsp2XsayROk/S0/b8lS0onnaaEi7EAmKvXg9u
zxev2Tv48BoQmtYsp+69hHcFsNyY02FIXjML1xZsUdu/3wBPxhHvigjnt4boaNbW
eXtCFrBhqYlenB57xerutm/n2Vvjz8MZq3oTiWq0qgM0c2BGJNXTY1/iiHByOotb
OTHG2SHPLKkxZqrTfFO9YLBIwBlGj9Nh2Z3Uc0a2knwWZThlkeg6G9DmEjw+QbYR
cNun/L8OpP2gg4tTQr5UJQhtWMCzkuq3vIcVAXXkP1ntHJlnL2KnZVdPWkAudzh9
dhc3iGTCFiAEG8E3ixubNBZkZzXFcdYaC5AXwEqCdfQ1IvEzr98JdszdBijRFFC3
HynnXvF7iLKWxFY8UQ6+l+j8MS4u9qTNyItVIsLkIQyw+7E/HyW7Qbx8VMgBgQR4
eeMd8vELIuF2A0LJDOi73gvk5jtK+05y8TiOS8n3U3tjKgUWA2Gf5yvfDdVxlrJZ
mj6bRvmGXz/FecGg39K1cpMZB2+u6Hi2H/H60ZoSGeM+YBMKadiDCoh+n7iUIyvz
xc4pOmENW3R2kYp8yLspqRv5YFc/fSvXgwxTyBoKaHnKCUZmHFGO4IijjUxkzQw+
l7ERIVp/eSTQWmK7vXcaUXEVwxZC6v78zsYUrWu9GS4navPcbTFDJ+Vy391g6qHP
SW5TNvBHcAmUTVkkLKTNlOVblxAsJ59LW6Y1DZ0+e6A8Prpt2IPBfQPFVYYwA7qd
91BzDo8fxfCZ5nZ1niFj1tzc350qTDZVYoy+hx3DowNMvXNw84pg6FeO5AUNtyvy
5h8rvRx2i1qXmqJ+aVhvT4JdTHJ2h5cQRs2XOUMMH9/7ICYacSiYZSXBWli9PpgE
rS25HlvhPaKL6f7xEQNlkYttzUseI4UyqQVoqEitRIBA3BsANMeqqPQbup1Lc0e9
JNLE7WbVPp6aghki2Po58Mgcj23wjuME57lQ/p3yxAyd5pcbMWQwXOFmhMR9l0lU
1AtRP8gz1LaHzZhdj7bAU3in9VkMptId0D4BZbVFPnD4Iuhee5fsdgRijzypiqja
Kou7PWK0fogwmhBFZrbHV9nFm2z2hD619eyrOH50qYAFWqpvn2CRBGKMi7HiFmo5
AehXRdmGYTGijDIeci4N/1TBdpFTvs7SYp/MUXtGpbu1MlxvdGmlVNCeFg0Ps4iL
/iWrUgo9noiyL0NKpInvToj1Qhx3p4PL+6rVi8FAuvgQ4EjJq+05PKtn9CWZk0Rq
2W/NeEKhLu1Ypvk3IuxQjgDq41YMmdo0elxWqb5DHz/kIjxq+RXu+wSSFFQjMh0y
kU3dzMo6wx5sZ3YAIFeHR1Y8Y1wAoAddGy9DtgIHsFfoixQEC5maGtSQCYjnWa39
Q2uQO3WwlTz3AxaokTevkxwmcRT1hT0zEEzCcxL35NXHHRShQ7JNYYGJs05plrBS
o82GM6IMFJ8jZnbvr/+juuIbOHlHStkM999toBHm8PVBVbalnjOT0zc48dMuu7vk
eFJu53LDhdGD6RQ/qFHlDJAJGAhEXSiwLTTv4pRZXLjhY70UAlF1MRU/e5w8+gtg
k8jJKPV/cZUSRUNjHao+8kN7QNE+m7aOT1FxRqshL162wlq5LkLgO6HE9Y95ldXw
500g0sS1C18AmzV8KbN9x+O82nUDdMUWzzZTMg6oE7wjRQWLhWkVcGhHu/WhkG5S
deUIVE/fYrfFn7yl8bPXe3yLoYTSZ2sHUyEfU9X6SDiLfhD98nAn2wZF5Z97s5LS
QP2wleywmK+gXgVBfdRw0B92HY8z5qR+geJoz4u2LIGy3TS5YsiPVmk5div7sM0F
4N5UEvuqxq4drJv5+PGYuaUdNkkDGscUCWDPc/F3AiVeczU3FnFHaiv+oFldTVry
WZgdGu+RwQr06tdQpEVdmAch+oCwfrnLW/NvsZ6LUSkLw6gpqn/qFmoKb6Ho/nx8
dDbv5rY/RTqLpe+cRhMygmhOEZ06xyQHWuw7f2TrHEmR1rNsyrjxhkEnydFVMx+R
8LlOMcfxRo8zBFsR4HJmQqOIAy17md6Wt1+31ihmu3ApDIMs9JRLkuSgYJwbIrGW
i3btcRQ1atkKSDGdu+1BwEXFr0r7J5GWjuvk0fJ9LzJQ/IBoLcLxoIJzttHT0drR
di6HwFhf8WyqpkoSur7Afmp93dxIRSquQYDUP/nGPgJwvq1N5aaNPr1Mk4uijWfv
TpeJSR20vZT/g2OGwzlbj+c6R/pez/9lwetKsIqWlhLk70ZyZwYtU9j3t96phE65
1TgwznyMuSINdjvjuLiByGd1hvKBzvowAdjStFba6zH/cMlJYph1woiGamooKdnx
2uEh3dNWcEWYN1Vh6rZx0vLVwl5iBBhSUyQt2IeyomK1PPnyHB54c+66vg22RdFs
YaktcsmIQXsoIUOpHaFqs9Zy56KMpbHZM+616iG85CvBs5HUXxGXMmDyR/Mszkbq
eBrSSnXks68uyXymirRZh6iQmY+rpvVrKESbxWfBPdR0Fs79OlkwTkr85pz6PdoO
XIVm0MgMq6BhVaMPoGJycq5sLVh8dSlwuZdEqQ5uzcersGhQ+3jiAc92f52LHd1G
zBjvjr2kR5LDAquFTlxq2TFLDFdeGEaDm2hRWRXEk8rKx8nQQm5nD7KdtLv/n9U6
FPvqW6NUtuy8RSdyW+gEg7dQyGTSKBiTURAa/9OFJJ3fhbOszKcmn0XF1wHbXfzk
CXIn+uuCw+VbRB3nKS5zKJVq07HggFD0uc9kW+MJB0wsIrlFlYtQ2/MXieFE2hnw
CKeqZcTvGw/6YnItib8RKk3pHsmK2eGBtxDCyXAaZMZUt1u46O5PkgEXsgveCyeC
hOMCXovJB5LtKReRFlE5SjQTrtIKbxhZFsBtho67Ahry2ARGh1RXk3XsAP7W7G0u
zhc75Xkr0PqZsLPDaSgTzecuOPD5wHbPZAVIRHZF+TmJAgsOKGDzBmN/24q3/dSV
/aRZYoZTL5GMDBEifIhDdE5DoJ8+I4rHc1/kImgun57h3TszGzIbuMtdM1m6jmA+
uKvu6rNhACRTKAmK5swyM7zYm4MIejBDpegCpWwIiFTUoBf2AwOhhHF8S9ULC1Mg
vo1IycVjozEHebpVyT2/J9HCEnQGS8+6otkgK6g5yidXdF+8rMkePBStzXOdl3U+
GLCItwon+YtqEkCr1Tp0yDkNy4f+y14RuHvxKRRQp+E6HeSiLW6EWlgyo3awpQqN
bZeT3IRM1qxfYIH8IFctQEEKnjGbagq+fbd5C2PfIMb0U+XTxVa32dytua7ns9kD
O9TRXmVDjmTlZlpPgKlGStk1zs35Ja5JaqYAdf0JapkjVSbQzQhY4N47/NQfMjjd
8UfwFkrWgGOG4OjlA5Bw9Kf4C36C7tWL1lt2MQKvs7x8ni9RcejnzjS7tkb4TtPV
+iwejwdI81ZaKQqRqMT7WKuMuS2dPqhiBifZR2YDGPvADN9cdcdwi1yzdN3ckFcW
Os62WmH93oWbZJsJA7W26QExOgmS59UEUZ5G3fq9RS/W+0WY7K0muvNPulCpQTXz
4tPwuSSLqvqG0x5ECuuXWYteWOzrJXuhqf37qnT/+x6ucmR5+WXmRsOh/3OTRmem
hmmeLGdz/JULa9Lfz3eGE/jvViqGY8g8gtM31jVtPWT/pzpVhQ23rLC7MM3nSK08
r/Xmh6zFT6mr9Og+fIyXFqqEyRpMD/06aGMF99M1LUaupQfUIl9oYPCX60GOpeX+
7ssiaGwV7T6sRr3FDPV9MpAeATRZkApKmCDkXiHeOER5kfZ8NcTS8oYGdLICYbnj
G6ikfTwxhb53WT9+vw8zOohbRNU6OY3GwTW8JsjWiwfLAF3g66+cvZFxUW/2t4cd
Jj5meap69zBZyTOVH63Aimz8NRSowtKn/ateQRisRzViwkOK9W4/SkBknEOvnhYK
y6qUJNwSPPCuFMqCRt1/y7oyQC/qEU01cywUItjFSr9xko8AiPvfyDm6WV9g6LCz
Ej3uNjMf6eyBdpF2LggnDQKWRNEwuwBDFOkHGetw9Kh595e/hpfdcBeUu3PFrL9U
HZfGqNsVAmp8rif1fHwntCpKvjWYt+o/JrlnVEOOBrBGxAgph0Fnk6SCnwPeIk5d
JEYfbjZxeUhzVft5ROQn65/EDdcFwbZ/L+XPily6Riy/zavqxpfP4WtoLsXcTgZq
6AJoQbCIZ9VgJU2ML5c+5VG8es7USh6YR/sE2oQu88rlxc8xO8N94vp60UdC7nZl
p9KqI+4ceusgD0sAAJ9fa+O566G84AwztVNyfRjKt9suhFfMaAeHxkKLxlc6AraG
l6jclgIXhdNUgcGjnHWXU+RqsO8RhLZArQrFm2cmN+t6t3Kewebnx0nKnb244mby
SUKoHBV7awQT7dd7w7gKE9MneitjU53f+l1Y1Nlk/eZUH4RU5ncUABgT0AHgm3wU
z1gu0KTg3nZYHKKbCkMufgTf7tiRm2htxenG6lffGRFGjqiZWG7zqE+UuXXHAmcg
eZfEuCJ+SO5LPnZYu2tzakUF8i0NjTsA9mXLH2MrbgJu/D+HMa/3wAX7ne9lupPC
1MULT5eXgrv5MHTUZ2vpl0Wbp7T+XWzT8928YPugVJ9JAid/x+n6yxZbvDxCb0X9
us8+Sqb1xBgsStKWMVFVz+y+ENdep6/olfh0SO3UAs1uqMZrLtgiRT1YlKvn8OgV
cIlPo31KaEqq0l1fcDDvls7CxPOMl8xA39B0CWglgp9u8sicQ/1wOQCBrOczXgg4
o+Du81aBq0Brn3fTpxOFKD7NaWSAMlyJbBjKrFB+4eVGZArG5+/JE9pPIrVzqPbn
lhpBTuFoyc3SMpa65LxUjlpdHG5Ems9/lr6nqwUklZEafHc+GXv3bCJn9I4Jn61G
5C8ZX7dZpov54NTlcBYsOKmOxdYQ/3e0njk9h/n3m1/C6BU/LTEOzDrvPzp0UChL
RgKz+LwBFwb6LaoXsoFxG8mRc4oZPqvZ7oISn9DOydkwN6ouWe09vONXYD3LEH4Z
ufL3bI8cmhO80Ni0bLpO9t2OWkzxMAg8wBXOUZcN68uiCd5izRWDaNnvLh7j78R7
eXsaAPHbvXqk80XH60uIBTK0gc7l2STjNGuyTaDL3uOgoxeS7hRIO3B2hg+03Ky0
nndL5um7lVWUPOr2uMiY3hm7OlDVDxn+UMBGwE95SgOWhq8Fyt/A9gCbfpyTdJd2
aj6OenjLJb/yH82JkoIuo/pVf08/a+zd37eIu9ZOW9Vx7eG9TdfNap8Pp5YiYcYq
rNZeOaJNoMZEiecVPCRmgG2Gu3NTO1UyxzW6QkstqnWmEsv8EWiGzmKbAgMXYGJm
7DlPAqnLjDMy93VoJRAzbpIsmloDP9zSCslWfHJ8cYpryaR2ke9YGO6Tt7M3RQND
O+LzGdQWbQaBS5xZfmVrVfVeekJhNw+j33Jo4pGTES64//ICGP3AOqZaI1OxxKgT
nHiO0jlVGRtRugI1RKPhQO9FeWwAkopZ+Br2stmBCpUujFNdpd/fnxAu2HFwba57
kruEAUC/acbOsLnXRANTaUizhkf3a6idMk6AHq5SPY58NZBayrNB3J3KcLEU3vRn
mR9rd03DD7utcZz9ygR3y3MtrWnYT+i40LYtbgHmjPKzuIl7+XF3+8Ub0wGoeEir
CbRakA62/phQwsyVj7Q1ljlRijMdf3YKcib4OhjgrDQW4cGAd1rxVk701O2Fhdmf
3zsSVoIMtaHRZQL7N8dYfDUOtZTwgU4qc/AYHBG8kOh6lWUWsi4gv5GhUnm1DJ5j
vgoRh2M0xN7xQ6tegGGYyGHj5unjeW3xrsAQu9Wqdjmk5CW2Gy+0igBGng+ySABI
D032OhSfgNKULE2u8NsPLXd6TWM3WQmUzlJVMigQkfLMMGEJgFZ2iGJ5rguMkSUt
9rq8g9hskLYK3j9nvgJEZzKL0Cl2lvNpB3crWN1398rXLaXlsWcXzfgRfO/gPgsz
GvW6WNJ3XnsUl59UUMvt0nuns+zKbs4XBD8vAsl/wV3gUQ8yFlrzseur6Ko1a029
E4cmEs/bShlTqMqmVsUkbwY2VWZtXyU5FmEGDOabnfYAiRLwEJ1AF8MSE5A05SOm
sx3+6H7UAAMWABTqDEDqZgcxQ+G80kjFBk2MBSNaF+w1JJfX7FPfjpAj5YdhE0ZE
JpKPdpV/Da8nKNbTb2ajQob0U2WqkUS09ykvgEut6MxJKT9m85lEH6SYPYBPKqDY
4y06sYXh+nEmn/kQ+fQ8/9mOY+my3laUBTHjsn2wSmEuE0DxcK+Y1rgxyx9hEh4s
i2gC+VBAo6eeYNqZevghhoWuaP93BCxg+CW78wp2t5J0pJPE8IzRRbnOrLT+aD0m
5VdCpRAdwjevLSwhXTs+JHdeq7u9CHTMuTvkohq6dkfEVWAYXaYULHYLtGejIDfn
v+zgJ691q8HbvYidvIU1AbvDzv8++U9cAzXx/TpwSk4on25CUAR7DNqh5YjQOsaI
/a0EG99/dN0rytYscMOJosE0m7mj3HJD73xCTLATsylISsRMARrD9aLD01tqNIRE
iwNNdocVfWkeAHSS+qS9mp6Y7RY6r+luN/Z/nvz7/gyZVgtn7zq3B69MdEzR90rX
K5gBGoVqmVOrvVbTqw57NwbKApP19bs2yxdVz+R8SfLGqeexeD74MMNcVBQAxaNf
CaWNtR70i1Zc41qzsenvLr5BV4upLPsWXPJRCBnz93EVgCG83rMb2z+Ra7rd7RGz
DRr9CTe2UOq9BSkwrBZZjI4D23qZKbfR1KcoVkwJXZwpO6ZXo+8jGhmeXcbQHFTu
Y3wUWM02WKVigXZGg8aNEFN7NuRhDALHYR2Hi/jMKuRYX5k8zPsCzodIUoH2gSi+
Rqnq2Gx8ImmVT2reWRJLNDKF9G0ilm3KdEzWG/G0IoaSfb3LFyzQATHZ0+sRrmUf
DhMxV2qWi4nOgvqr7c2E4d76ZLYijszE1qdb3NVmzkDrvQwDSdnqtcupRzaZ4EPL
H+p9r+jYOUT5wAOwgHDu461ia41UiZq49cRAz+JIw02nwH8BTXZiXXkcB/iq3hEq
xoY0hh6usMPyAFBA56UIPPXnRs54/sHVLrOfk7mtRLEE14R9yMbITGkrUUE8Uw6F
pl/S2eNeJsLnSxZQVMbk+bfI2a1i3f62b0AezM4lLCnj+XgFDQsVZH+eCd8toynC
J8ET2bM99EXqQq2tJ6vpsCmT2kJFerjm2vwsD1ta3X/B16u9Qr7D6+ZAmqDhvHGt
m9jTaI1zA72crjklpNpK8cLEr4n5B1QAvFgH6Nq1WB9TyVLYy4DGvpPmLycdg1DO
bxogy82FXYKVr5h3wyasyLAY+eAxB37++XygS46d28VSJ5g0efi7I5pkURovfXib
OPY++OkXzvHBpHViPrg/DxpLP0RhzfHYsvEtceUmTIuY/WprPUak2LuzPpY2deqn
Lc9u/pNs5jTrnbBwZgm8gbA50mgHQnlCdkPVUcO36f8cwwI8isATgIqZkvLiJsU7
APApttKq7wA/n0PlbsIVr9aH6w4QVgVXy/0JQRDatrSLi/dbYJMOQDRJETqwe30K
uUN7SXS+R3xnK60C9UDfTFdwcEAFgSefP4Frjt3PhKXXWHx5UknZDat/aiDp+6eh
FFhYdszQWjxUPOLpdgLvXtPjybmwYdgIxDSMwxpRkaKjO4pDNQ7GHVLyKe/VsD71
XUatBPWse5D/k3fED1MMZ+zOJHivkxjScBYhPRtLscvVs4W1mbHq6Svtit0snoQ4
+po6Wjy516tjZUjCJhFVhSIOr7P+FVJSxkfz8AFSYqfVN54b2PkKy12dRY9tQTmE
Yq02Yji2eQFjfoPg2V0uRjay8ZkTYjUPAmuRR4CRR1yTTGKFsq3EfqObngc6gKBs
yUT10JAd8ui0pxRdtVB6ps5t2Mr7VVa0gDGy/f0JCOtn7I4Ii8zyxegnIER+ej6B
ZO+/k02tg0TBh/KwfEsAcsEc0/U+uCv0STfw6D3ZanJVtNVx5q8uY3pOmyG5VduX
DQJVJjRJRpQMdZfKFqJvK1fEVVftrQQdlFPC64veMar5mu2614xuLGHxEVJaKaOB
5aF9pTNHMTgZ6O6JUOVyqdT4eTSiXpZ6bqROV/AFylICxTFbpYhI3EpIXXImScMv
3hewJ3OeW8OMAoqSDyBmAf4WWZtQvl+THk0eZX9+gZxpQIzIuEF6dEXKUvRrSgP0
4YnMdo1iYjif3+8MthLmQs6jakaZO1O47DToC7KFj91l15VWfaZYfKEsc9D1Q1KF
/n6MRmBK1wDB2cLK/Xp1SgMRj7BSqSKeeYYbxD4zpU0zsBSsyQ0SaKbW/1zQj4Tn
+6npYPqeKYBRrm3BeANOfalhP+XSSY5axZYQW2811HfUKTGBCBDoMt+GZmGXVp4F
f5A5+CzPM62af5vnwRfAXiKegZp6DPFflc1UcLpaTqcO1YsRhTeC+IIyADaQ/zEW
IdjyzbQkzbY3ApZndmLJzrvUKXWe/44M1emBopR7XJyiwOhx9KCeKwvq4FS+3TjP
z+8dg87kNyJakORdSSrqdHXdsSy/fE9AzXFSgkhHymrJkWwuFytmtYTm1w48S198
DEJCnANXrZQt5PXacFKUxlfde3S7W0bmZHYB993hIIMwCVw5MLufuMG79MskYCg6
1a4k7e7D+iXLXu5RSY0H90BT8qAkNEkEO9sj8Yu+uDdQmycS61G/KCddfEAI+JXT
PrOA1gHdRWYZLkCanQBAqNhHYCESXVmYo0D2WaEaa8jEb5M006EpB6AeTNOy8qSF
TcHO4FgEWUZ7JHJqYZ0UNHvl5aqNP0ew8tUjvKH/8wTtl21Sn5tLu7bGyql4qZZI
2ynM5OnV0yoH1Kk148H5RqLcskuW+oglRI21fWN7Wy6PfHyM4xQxwUyK6RZ6To9c
t//1rfDppLQwGkBPc9pFkANuruWzrLjxCio6ka22x3f+BS1EY0JbuGYPnv1ukhwu
2xQajGBogbno2JtUd36eOKxwPc2/0zqLOj4sFxaDmRCQR0RglvIUWKjyW0xDyoTE
Nyli1EN3loBct2gIYGHOz0+wQk9NsBdZJfKcwR0N5bnB/F25HKbhELeiFJURwq/p
+xkLqJWQTJvzWiBUtkg0wSkShw3FvO2Ya9tk7ZEUSFSkTYYnzofWw22S99T+csEg
dOMwG7R3hrfT35D9ap/LESLzjUrfXBhHHyXQKTegCkIE8JxUM7IBdZV5LbR64AY3
IIXwNSM9rRvzxwSRX9uZ6UcL2gOO38c5vXlZJT7S0kVgKKWLEQ29uv+u6k3LW1ci
x9SgL7108H7d82ekrmysbYSZsI74YI4vMK3ViFaaXDegAv6UyqxHd/TyVeVSce7u
JRoGiuMdy8X8OLELfYRy8BRqtTH/mi70dudEsDKkqtsfKDQStsbD0VexL76FSu1h
BtqA9UHVDN4SnueJwmy8A9gykgnm1xWABRqmOL1TqB9TsVNJt0NUD5EsgOsYJbtu
4VWQkW9qbh7+cLFjAdGS8qwBsi8wB2ac/JgsCdCk3GXIDlkXQKb6wyguj8ZyJCSz
2wgXzdBMXc04kEcb3OuI0xPDFfVB7HD9z8KPLPeXyZsg+n+xQHA/MEM183tv4HZq
DZ90zTuKjtatPubhxboPNHiT9TloAVAca2Cob3DNbF2zxhTSnLSsFPW1mVGcg2ee
LYmo8fCIAENDXQzSKnJoccYJqdug/ZV5OdUnE9vnvIOjD6Y2HsQjfNsjCv9mKG0E
mYmuiZyo63asjn6EI8rs86sFoxVz3kc4roBZ7Cd6VClUCNEdSf7WhLYIhxKAWT/H
ARQDxJigUKh8oHUO6F7XUBMw8ub3opxUVzCHrOkmA7PFAzm7aLCsDoQq5aG4DM1m
0tOwJ+KkbWBNpN+pA2eZNwXx4E+xgwmIQl4fq7GjGlGMnBnXATqGhPAr6SL9C1fZ
6+uvinBj2hrSfhvfjpFvQhoEd4HxZjs+YH9dRd8HrGUcS4aHK0QGtSf/MMRS2p4c
occbfK6vP0xe9Xz7rYEGtnnoosS1neqOHoZiCIGnl0l+9H3k3HEZBGLDNaq+Pomk
NaYzqzUdMi6lEIfnFSAKCt1uTtZyC7194yCtjTtksGxEMKapkeNK1cs1FlPb6Bx+
U8syMhhKf+Q0VmKv/LUKzV3QcrYCGkVeI9HRTwXexPy7AdXAkLfd6487p0KQ4MOr
vrv5ArXDmJ7vpfnH1/CPjzVXesVYKhdHiqlZmkCTYpbnGwtqzDgl4NlaDbhleQS8
u5iVmbUi0XMXLV/29eaxpX3s47imvNeTaedEucToZE8+Mpv+PoNZgT0VprAGin8w
tE5+a8MhcYydKvwgSlVZyvsTL+LAdvnhHFet9GQwWl4T9eYYH1uPuUcogonJPP3Z
XuZVG2uAWSVEk2FL9lsFcp9fJNeU4JQ2kJR7tGfdzWELZTljsiMAInHRZX18B9DZ
UI1U1VEquhJfsD8aje7foRYIVlpFHzlOweavXTAMZNPSTs/iB66ZueZ8PuQ+5f3U
6NEcRwoVcz7gjWySl5o8R+K3JVOoC70UWqtMGnW2UMCJzBYQMaY5bLkeTeKnrC2h
MFA7u38qaQHf+FWwdBL0OZas4Kxkf0wKZ7cw259RTjqWiP7GfzIbHRSxAG0JL4Cy
85mU+u+S32hX5W76StoTTZaeRQCRPuiLf0SO9qjhxytdl+xiOzscF38ZK7VNiRWC
JVM5aDj+pFNjfeal4ku8A1PUsfNfqTN+juxbtqBAxAiBpss7yBC6UidJSyFfY7Xm
JNzSfriW8RbVQFYFec87Pl2DHQDu+/e/oDG+wmpclTsGS2OUf+ymYSmW8Ypc2rWl
prgpCzPtnnL+ltulUo5ybo82JK27J5f66xcJKIdkJoliVq5pvMfOHNU8jObdIGGe
j5sPCyvI/vXez3j7osH12+CjW1cx6auD9PDdkZVQIvyFa0HmENho9Am5WygZlptl
aJQCYA8qqmyYg1VENMtsJj8PGapTXXg22uenu+fWHYiR5HFbxrlUckiay8ZDwFtN
+GPkSJqShHttNRFLWY3HRaCdjfsAfCGxgTJK/fY3kvl+ofdl7I3lMxYfv3VhmwcT
cGqJ0szPgZOsyGvUf1WXiy8MH8NLuR+PjZX5ytO1F84I2da4qU2rJxMDRKacWi8X
LBCM+eNzThLs+R6Eir5rdxatDOgrR0FnH2auq0RcZ5WBgIjPPlyNaLqjvdoxqQG7
MBJIGbDRsfFXQxge2C2/MKMx/bvCb6PFteP6lF6zdxom1ixb+xNr+BSbcElqVvX3
wrMTZqhTK4E2lCQROZG6NY0Hr7gclRrbAsJLOT4P25fxkRaxLNJSAyVeP9IBM5we
IEP/jcbcZV4sE8Yl/lh5UsP+fxRWLMe/ULdX8GqRySCC6NgWNhRkisQY1DhoABxp
YxExRtbnlWqt6w1/t8MdUj6CpWfAJvU69gryzQqZjnMMrDxkrw4Bm7TnWGqOv2bs
Ug2SqBO9AhnSgdTKVk47/XAVaCllty4jwH9EtWAajm3VLmqfHifQ07YH5FH6Kvuk
SYzGjV1mWwJOCtbCECg697rAsJon/c9oElXi7U61xLMQ+2D3jcv9XAVt2PIYdedI
XlrNnKNK7aboeSE4d92vABQYl4tt9p5HR4VUmZVCRQLEiWgrWBNk5iiOeXd6Lbfx
of1Gp2Atjv0zUCPhPtT7CF+d+UKnSTOYMkvGBbVaoVDieLNDY00QzI3NIKtItWuM
YhJ+8eGbCN4CcTTX2ayMwq9FJO5yITVJCMQXOoyqc7PLMvVBhAIXHSBGkRXAyzwc
jdrXJeBIsyGyy7Uk9LPW919pQa58c/yBtutNCa8qOKC8t0qzJGsUGjJBI7JXDoG9
YyZ6/+UZhSTpjfAGzQ3L0I/K+8cwtCoxdhojtp4CJq8nSeIJx5FxpcwrDYZX3AUW
3FEGYCmOb8eLpFnpHUkhfuIpo8MJuzIap0M+LWWL3RMu/lG/Ow+w1nKr3B5/IYXC
+gwPRBV3dfcHFlF5a8ukpKdJmIuBo6r6dZCDnJ98jEUl0CuDZd+vtpJj1oszJ4tS
wECUfrGnTXlM4Zkpj6JFkGFz7eLFOqd6NMpXOFQVxXXQvyY6xT8Mq/GJ+GX0jKmh
tCkFiCHtBR90MwLFtC+X4sZpFuvTUQp0jq0pnKLAokeRrDxixJPtAiSDSM+lw7DQ
TUhUyvlw5ValEf6WWn6AGWuOXYJUbmmh92fj3JFAcLAKAfkn18LW+jTT8c9hXa78
xIf5hhrxhkFMcRSIKw5IpQeTeJHf5UY6qKDKF6azdo1ZNQga7o6xm5rWAFhiWe9L
7eN9jzjWCP1ZE/2FqMVgCtm/FEWy6p21xThuBw6SZLWzgBdaYi1TeOuLJxVslNSB
qJHPevY0ICtCkx7AuCIrCI6FxEqkvDez1QyTjJNO/azjN3V+NkETWt5sbF2RfnC8
om2KI4ad/5B8GvbS69cjd2hVQvxUfSstwjwEG8H8fLa5KtmgZrgOm8hiW+WuAPNt
7m1HcB+uB37udRG7Cy5CYImpWuE228/YYIkLAORwnlFFQrVbMSmVm0h1yRoaG6Ql
KY/5N5ILcWiL8dAyRKCqT1SUT/C/mu4lpgZ8zhrsrBs2teEJ/2ebaWBl7twGhONC
Dl4FFiVf8n0MwZKr46oZ95ZxFUa1Ba6+YA3JYSkX4krWH1oB54b+E42aFW9QE787
S5gs458vxkReQ3mC+ZfhN1Vy8LKHt0ZkZlK6URTc0G3Rl9cUvXnWnA8uvmG7lCRa
baLKUCngQBBjd25r8CrpJ78s3S3ZfMe7lOMPFNtgL4LxDquUM/NQBfIjdEeXvb13
7bXhgQZN8lAkQALNtQXFCda4W6Tu0uRcJPo9oPXKzFX9v/3V4T7mLFkO+8bNsdTO
90mRC5CRZNjnQzq7AvTBijFeHkIR21BQ1xXZrbpuJyBf3ad64y6L9isxX0qCe5+K
a8a53dQmYKwKgkfq4Utk18Jy+Bhu3mx1CvCme+p2X8GWYfroFoO3JX2/1WYTSjP0
HqibWM6SQCEjZLg6rEii9zi9gRpl+dke/255VtlsYyow2nATgwzuO/a58j6CK3XW
7/tUDmy8mvFt2hLJzEDq5r9DkHP6Yjk0fLmxga4IRXEbWNCdqNPozFy2EnYbaUcn
A0W/CBEUe0I6UZLOhXVhTpGheV4Pc3BkO6ZY/G35GVIH3P4gI1MB6jRuEVpUjYPX
vFHLh7ZoEy8UfmNUtpgX0QdmrETEIwYbRSt7K2omzy2FdJssxjp77SLVYVAqc10P
R+aXdge+cJwy3kd9trrqzBDP4eopdweuYJUzsrx+kj87ribUmUZTzXvVj7gb7kD+
xOA6niL8sbU08bZKnmW6CUezKzlKSNnTTPTMleIOfDU5PRTcY6QYo97iwTEBzPxD
vrX8L81GqyxjFJa91PGU3r+BdW1WdOLVs29XL6ymOv2TrjN1OMxPaC8WlBh/HX/g
NJJhdudiZqVSVfwLQALliO5IWyf8gMT//TDSmD6U1OXfUCDKfohyWuhkC67adPvb
9JyUzY81/WCWhryF7wX0l5RXAkuqxsd8IYO4Vb2arU9V8owciF+eXbdWOnEq3jtI
Xal9TwNb6txWZVukjWPZIrUL51uxNSYYtMb15CwCpw/OZf5kgMb/zsAS74fYxINy
JN5UABotQdhyDurvO70p44I6z0LZQc3cfqWMOxL/3ZPGRYqPbz1hftpB7Afv1ggR
CenfhUBwzbWZ/WjyhAi6nLOIyW+kql1dgzL6uG1JNcNt/gkyCrkfCN7WZHEf7xpV
ssDkbv1REauTifKkowCr5fbX1YXj3jwCNbCdhXxnHBdcgKHi5uknNx/jEHafhTCF
0LtqMW2Th1BPoBXP7rGNWq2AU4Njy1syifp/fvAq0xNlPufANhwp5sMqsidICxLv
flL4Wr27mhptMhmQEgruia1vfsQJfjLwzW5VhqRn+ycRUAK7IdlgjwrU7gr1GQXJ
jw0PPQlnPpIJnaikPFFEPllfauSayAba54xRVxKAi1pumYlipCtqwnG8O/KDNJtG
rIEuA8sz+6eeZ2hL/bx2a9uf+4CfussodzvB1Z9EKywvAkSyZnS7TpyT1nh6uRUj
XUzadv3u5X7DDRiePK5IDjpRzBSn7V3xA5qzn0xLW2FXmXW6098bmo8FJP1TUCCB
5+tFZhj/JCNX30CocOVq4vTAH21hH9kpEAOxqS76LQcnaziqXcEZ6CphJ9Sy6Mr4
PWtbL3pNwMZWpWUFZILyo14YLJMlwbHu6WLJCYEflDkB/QJNlQwLVlS+VEUuEthi
C2iIUX3yr4fHMOTy9BgRfwz1SgkV3+ty9RMIuCeLtse+N7nlSZGMGqarn7VQN4M8
qc5E4AJT3N+uJiedsxVDmBtnQJ7UkcjC1BDF/EVv0ITyX0tvKNtwjyeGj0SijOFa
NF8txc4144hRXg+1o1RicARKHuxbnReN5CxyM3ru6tDV/INoJjP333M8TU8sZukm
Enm6l56nLt00GZiq2tSC9B6VL0WPElcDnOyE9v2aKpts7omtQjn60fp5LSFxpza0
MU1eTdrDwWKTDc0Gi3kxM9P7IkUYGSHxTWsZ1thPRuXufcBX3nS/ZzIts1V6JWv5
UmxGTjgvAMYrT7iv8/ujD0OteWEuXsKm+vJfWKuVQTguRMHv8hfdAKa/hrA6RDm+
ZjnD/oh2ZJyy8oDMEfqZUrg9DRKH6CeJPa4Brkbksnzi9Auaxq5cINgo3g7ysofc
paoFJk8mNL9cMUn1sHI81BOQ5Qse2ROKCymdqVSdmxOPnpjvI/5vWWKjgLvM6Av/
4ZnVPq64ANqHAaUKOC/ZU97BmLwbl8UXeE974pbpiuETIo699gyZwhlMVIEXCSoT
e311sJ9WEmWp5xkRgzjdjm9p25betmFFyPw8/GC5A6H72tY4HnzlxDyPSJBb6PE4
l/lmED0rRZ4JX8D5Uumki3gOlLBtaJ4z3bH2iD+emPa2wgcs7tqri89mOaMKncfL
LJEHAp69DH7ozX7w9ebMV4FXYOPas7F875cdHPeNQ8anZrJ67vQxah1VqcfurfGT
O0dVdl5JGLPdh/2xWBOb8l9UxvEpmVhWWCm/mb6sBqVkbhrsZUZ6bd4cL8EjsYY9
+eI6VLVdpm0u0yY//nftP1mtkNYCJD9wQrMxT2iN5nPbb0StsqXuAcNRoSZ1rcBP
I+T7VMtpVGb2V0MTuiLQzgbY2DLcNRVLJ+M6jGLkLl3tVUFj/oFpBoA1ZT+4WP12
BdOcDeLurQHpOsAuTW5vntZ93aFHTJ8PmA9eG7Yucep/uIW0HcF/8HRhGg6Ifueu
JtfD5Va9968CjIxqKaR/dKTsB7hBtahnamlBC2a+2wJHbPzXu5Tqg9TnFWy3HY8l
5UaSFvw58q2Ilieus0QZLIkTLR4StkZi3DalAml+z5BGQ/HljIBA7uf8eaug/bsS
nA5vpNQjxOiDFjYvOdCzMaeFCAhx7Hqnr3filhMIHAK6isRnRwjmF2QB8TMCz4KO
yxy+szsCW9CVxmWf/sGwT8jskzydPL4EFLie4pFJ0R87pmfnSX9sSMBzzBZsyzvP
kupJ7FClxS2dx4wPs2rNB+sKu/Ev5C7njx/FDSVn1u4YW15LKUZwrQO2vxVJgP1A
TMCmOylBLnjuLwEdjVJFz0ZsdwQYISw954VdU8P7BO+gqCur6xpDhoKbCxgmZ+At
LIT5P1iLpZyRqprQJ2rttlcK7WK++fSpELfCuY5hPdgqcAi1mCmoP8jqYTfbzS9N
YOcT5OEVzG+aHJOoXZOmcBpRUhABmGTCdz+lkn3voFoQAG4yLRRBWpjNFSvB5FYj
CbmIgJRfuAkjDyw+wcXFNljQ5DJ4d3etuZQDwcPUV6GGJWZE85RMuBQptYRI9a6p
TU+QaMSgOB8fV6uUCSwGY0hFtRZdkxJtDqQ2Lew5ZTMHvU/zcqdFCXT2NFS4DGFh
OgW/AtQA4HmpVd3Ej4BwkWQCr7HYR+DycBLsAAG8n92q5c8ThYT6zG17+LGGJs+6
OCyaWMY/ZyyC+UCs4CkAq4g9psfOk/1kmktjpwzC7ac5UUwEYl/+vCge8xT5ZsbT
JR8nREN7vcREAOEDZZq8rl74YTDfpWEilzWs1TT/FDRdgV+pEltE09FidZNVSf9b
F9+fYVrXGTavEp4E2RUTxF3SXtSitYIKsAQC8M716LeSXrWUYTZ0Ti/VZZHDY2Y/
65k7/6zGBn2cdQ9DL5UvP74CeNmBDH+uBRBxy6RqVI3bJYEbEtUgyi+kvj0RaQDv
+9xhPHXGOHbo7RJ9Ur0is9Jvf1efnORHRQxfjZU+is0eamgCz4icmsNhOxsHTSAJ
ger5VmKJji9ZD4NyF9HdeCR1kV6eyoZXa17BoIY6hyOFmdkpcdm1H3PM18Knrzsk
AJOWKMfAYaBVLtXPeR5U5+ZMidx57nY9B/mYHFaGzU4zf5XPwNasd7MDRIGrSwY+
OTgJTf8OYi3adNlBZ1YRmQP4kNuWJfWCDdOyySoAvnKwKoQWuCeQT2m/KXIgFOWE
SPcvAVsVxVJz9DWcxNAu35bKFFIoEscElX2jHNUXRcAXi4tJnqWFgWLs6kmzuyZw
ZglWS1cp6hyHcPEwD/BHyD5ATiT9pF2mA8ejj3kPbGyMxSRkMFddQLVJ6Hc8JvNl
hZTO3RtFL13aTyk0kmZNCNXPpkT7dHakdFTl5IEH0C1rzV7GCByBWuf7hQFK+arO
Kr9T1DepB33xr6s1varmzA31rMN3z8tukdlQTqYpxxZc5qNqSoD0Z6L6x1R/an2U
WuVtLmMA3VS5OSYF2SGVh7ADw2gOTEB4ak595NZgO6wTni/L1S0lu01vA/eNStoX
lbaVY58OGdlmGltDhZPxKe214zBPEtfM/dMnx0bdGSIGS6KdkYFYEynxgunZReRX
/i2p0SUZgRqceGzt2VHeGrHEXUs0zlLNCootGCWcVxA4TjlieejpY3LjMSUFpIcR
xoVHdZZBsHnhLyrcXH74D+Bi2fupUu3GhcWhx2hMYPf/BbPSRYE53Uobze+DECWK
YVznkBtvh4jJSDIS3r9rYvEm24FFt133lOangJkMHdlko0CyXaYec3DxIAVxsk52
76faIqR8HADkhMVcbvIHNRR51DzVlJofp+Ryv17Qhi1hbsPdQRZn1t8XK/tdO2jD
2s1CjCoUtIsHgr0aCarfZMX/tpwvwx9h6hk4N4+0HtA2nBIWV4U6kcTu2rwMb/T8
ZvLvWx92ps9stuNnZPyJ9gI62ekikVkNBwXSdLN1YNdjP5w8pzZLUXwMYCs5GhEL
tPgkIZaglaYuUFsZz7ni6Gk4emCpnSsK/pr8JC2b9vFOsyrnF7HYsjvYiRZePjFK
mjCu4BmJpfqSvntkGEyweSQ/PpF5cm5dRTqiazhjJjI1r2z6CvR3o0MMbMk/UWxk
ZuZFCvUXQA8o+vpNYM7/lFp5cOxiXX9AdCx3UO5mmp/TC9tGPLw/aKQwc3MGWLtO
19HE3dEId7SAqy6od2J1GZRrcTL3psETjH+I3zDUvyfM/nhNmerUa7IKip5u5ARr
55kseM7AbVgEEUlnw7QGD8UU02SvCJy8dxZopmm7/VUnWpL798MFDWwSc21+Wekg
8GKRVL+Y1uw/Mc+ZNXnOB8eawypN7Ix0MaHnKIj2UMkoTo5vW0A7eBpgIIuWPDdg
/SJoVkyWLJyG8a9ep+WxGr918Z3LJttzUlc/eXmyLHU/Ynmv6y1yks+c71c43bX9
i6F3gs4pGmWv674Xp6BGRjyLtQKAmEZhD47fGVb9hzVVy1myqiZcziDCIAdjiKgm
hLbuyTFNZof9icC6a15R/WzBmGMq6eKLaoZBpYA7k4CLYiWTytPWTgRKWiGywFi0
6OK6lB8hpqJYJhnq+dbYWtNrOnOR0qYYWU/cjFmfi5VfdmlMhJ1Ghaqr2SEpEto8
wx/7IDLY3wU5yZETPNJNZ/85DWrGogoOPSmmuBK7G2gHhXmBGXOdF5AV3pqMKdyw
m+pLpPpLzTxRJbv69y/iLN4WqVFfhlb6V2ygb13V67Dsau3Ks3JbIRA2cO751TYo
uqKOAK7NdV0vQ2fWC2vBZn8a8u/inOmL9N1Zli8MLJawzKlr6emyIkq4Xnad7IzW
cRcBoR+lj/FVycSX9TEiDvcLuoQnKyzovA8cbPdcjvLTOuLABfADbjiRq5tG4pau
Zv7gDFTtrGhyHif21IZWeD3nT6S873a7tj+MnhkBEms1kKFkE8o2waPK3pR+5Vbt
RTRrEL9hbwdDo5/qEW35wMVfCOEB8IrhxVpJPnigLIE56w/TG5i9w6zXNxhmFfaM
5QnkPbiBXyICen7G1tWRjcXPCpXLgYB2k7SXOcLC4MVaZDA4Joz0T+1r+HP1efUb
mMFP93HhvoRu2r5gmC5Qjq2nGA2RgesQIsmDV6PSG+jDH4MY4NLjPyD+GdiG+/qS
6Aaq5QyQ14YY6Mr/W90KsZLYX3quP/AmPVaj/y9P8/l/vWAM5NswaeQsIVQP1olU
oFOCb210zF35P1t1HZIMqUXayD9EEtuQWf5YK0WC8kDWDwovTghmZZBoYuSN8QiJ
7VMhv3gxE3cM2Y9lpN2v05DUNs+ifcL/cMVuWX+6NORD3lruvfIz9V3DEK0cNx0F
bvliEprsOLebiolv3npeFzjMNy4cI6drEc2+ioQNYxNpHp5a0yOVzCb+8WIjYV5/
+H5MPIGUgJtv3nn+QgBaPAUVXywtsnv6qu0p+2SKXOdeTqu3atx6NK2OjGmXuai0
3pc9V7nIQtcEzOyCbPViC9GdoaFKlzbxVu9B9CevLbeJEg6WzZjXaN4U0JdbsR6R
uh/A+zeK/sysPj9KcubFHAKKnHwHqL+5BiujuYSJaPmlYV5LVUf3WGspFOgUCwJK
PS5gRMzSLfVL/vv/F/hvLzYjk/cdtjDpMPitmT68Qh/EMIljsxrlGL8NdTT7b9L8
SOrH0fYI9+4GeRg10g1jzYIMxZW/LQv99vSRARWqa1fKAROmTklybOSAREQ5wvrR
axbFhCBwl3fdUr5XwU2tTDWWARcIpcKsOGY9cuCyImxUaBL/VoWDRSsCJkiILVtk
3WDgktOxPwwWpo1pByTLTZmULAm7oamJwaYwJ+f3E21MH6OIWCWuZLGtWxlRey4e
Ex5OCOpcsF6OGRaazQeH3/iA8vgEmK0CZgOrlpAQnLBUviYwdNxu2kC9pNtuhNEo
Q45NBi4+4TDE+RCCrbFDDJOFlb9p5ILL+xk7uRxMraiuPqrQopCZ0EXpzgbxM/Nw
C7JutSHx8yZMPXbcCWhwoApMBlylcFqFvLOiloSdStSvqpj6BdXYeq5mxr8oURKc
ZRW+MXsnGejKGIo8CxrgtVyRp5S/qTRd412EdAEF/fk2aDnbmblUWWBwgMWuyNt1
NVqFQz1Mcdw6Gk4pMPcm7p8/KX/Fs8ZC5AgEaI3HuJT7TMVvtgzARGB3JGanLHQw
JPQvD1UpB+ts2pgnAbM5DE70u3pzLX78jh3q+fuVgmdChs+4tHdP7Rx1QQOvnY8q
07Afj7RW3IMCGbQTbSw1oGTfT0VP5zKP4z3B/YMZqjNyWewa9Rh+XFoNaX1vZQKx
xEuunhb86N3IAH4oHl1vXEna23a8amgzGEtN2MvYM25I0hRLMtUuH/mYJNaxs1So
xBDQKY87t3kU56FrD+oQdWH/B/Une75KZcbrQ0sfyw5gn7ZlMs03NkGDSkKfjWEf
4gYEk3i2tJWPTVVyeV3BOYTbEDge3NdQzgPMJwCzuosTh3gH7hgmVCuIOJd1jBha
iR6/E2KJZS7cj4pujvjrdRgxB6c/7fzGVYz6W4ysOHoc9AYNU8UWMuUEjiXTIhoq
fHJuYmDJzcP3mW+yuCQYWykpbHIypD+4b5oViZIMg5W1BOvn4NNr2UNupI2wwlkN
4cuK0OSm7/asYkHPBWs337/6GBCKD0YbxcNMWgJkPKcgyL9xqp741ECYowtoSazU
hNwNGWFTMfVvEeGPDkv1it7xdBdPuW7PZCQ/YmrXx8200jD0dA+UlSZfLbRKmxyH
1NYHt6qCGut64Tuhc6Y7/DyPR1qMsG2/aA0da8/2PuUQsrOGGrs0Uu1RHvTVERaZ
FaieHw0v93hyLTwc3y6ipgNXwlugAAu91oeaE+PsIvIKybd2GY+5q1TbclHsQabx
v2Sv4nyg5q5JuLY5pyb8+LSreU1uNmofdgPlr6bUt35onfzLkNDa8CMIILeLLiC+
igmTSgyyzBYllkBmMYhIwcN0PPRfbm+9vje/HPAyJkhRbdu3z3cJBiCsPndi3dkB
k5xI0jovBrkKqRoejQ+EBkudpPBO3qrw7qfpkKjrO0sds/BH1POWuN0E0TmaDY3N
G9Hg1QCs0nqxo0QDpuRSqC0a1cDOC9ItoIGdiHeqikQNqNnSSy/ZsrBpwqqtXNOz
/OjLv9FSW6LKgKMBf23mmfIHpKZ9We2cxRQDum3WEZFK97YNpduuo+/Cw9fpiW3m
gpmNscbwf7j4FT1IhoWRY9j6ND2KVM+EcZppz5nLkYFDf9A1on99BxwIubOMNILm
cfCCnWpAZhbHFkl+hPl3eaO+RHFOV3HXf0zOIu2vTehS06BzozvDmdi+o3v8EYIQ
p2N0Hb2kpZxK/PGjgFlX/meUf2qZAYtlvgDE0epeNMqAN/zaEiXEIjXCQ39BWHjT
ONn81uRyvipbigbrpZQT4zJ/u9PypQ4m8S1D7/YD0hvigzWbVx2Lk10QSb0A94BV
VrK02YGKr4D8HBeEXRMBkDlmmUu5BYwMMvwONIKuSMKD8UahnIE/cCzEv6rEF+x4
XbLsT6H3F8OqRN09WVBgmJUxYPSP0ZbBudyPA9y47MT0a2qgSsW7i/HQ0cyBjq9U
mWkKVLRiRxsWY0RBRXC0sskVAFqFKJ25vA88cKlqcQsnuCodqo2Ho1PHeC5go3/X
5+budU9Uy5ouieC8htbdN/eJwPu8Rq1QuaNX6wmC+7rX7OqArKrGLv9oJjA4XmBA
/36WRHqpL1RYz79ZqvPTWowUvluXuxdEkqg799agIzePQObK3IftUDSDVFzYFqKY
GOtpzjmwIiL0Et79/70l/rvaPZO5X7omonkRImHAKe0S9Yu9B+Cjlph2c9VoFFb3
6r8tVnRC97KI5so8vFsrMt8djc87cmhHmWbg5YLmX678fFSNWRo0gqZWsxfy6AGC
tUBtsPfskoEyj4/PdIrNQJ1d+0RceTJvxNXXAsv0PDn6pdfEITxg3iwKpagKD411
SaXqR22jhb9KTy1WXT2LBdtwrOb/gFut8VnCzFCdN/1YYdmyN+WHfR1B6Guvr+nS
SgpCYJSJmjvbgrjuTvvvRxCoE7rWwXJEQauWWN85vLgIXQ/ZR4vxlQT7nfygu0FO
gVvyRIB8m97wVlgo5enAGkwy8oQtM0hJv1acZYsrUxGO5PjW0f7yYyBhmQvKQHu3
5KEmHa+aBX7GwthUJ7clrhGP4g7s4Z6W+iZdmsJ75z6RiGk/IplR/B20G8MrM4/W
X+/V/ZH8pFH91o+JOumRvKKNr56AYIAMKzdNnJ89bqXly75tBkvaRxpyMUreUSXc
Go7iphudqvSdPDbiGIRQmeeTBhrI7BsJ79RGutfN6ddmc7azjKoULOZnhFez9Pq+
pYt8OrKVNyFeq4upN7mPcpbblsqx+dDzaPQ43buEQMf2zmrSPNV8E7S9TgtgcA0P
rDQMBudIq0LNkLiA8F4+3knOd9q7aZlHh+Uqn/rXFkKe3BVCFTTkMc8t+MfQ+3af
bdAe1evD1byHNip2FZeyQOHmfNyexKn5nBau7FC1bmg2aSHZ9oL9IllevvgcHUwy
4ZWq5ZphJi99kpbercijA/k7FUGnRGkiZIGP4xyvrz+0XEqN4H56LaYF9B4H70c7
6J42tx+DPNwtd7AfCZtWxZFIBbqtO3nAoaHevwYgpFPmEFZXmIDOHDBSlRNcLm9P
6AOThrg4X4+NBQRuc8kFDLj2NvnvRin0B/nUCLzcOyP1OBLMFlIzZm4AywbtHrwo
+o0gR11gIGqtg9aW7N8Crz5oDkQE/5WPmcARmNxuGfjJ5oMBVsdMJ6V1+aAB/II7
QstVFHdFZm8vaFaqRZuz5mp0JJEtNFEggrt585ynwVFTymtmzdiWSVZkD45ViMMR
9x9DiNTxwSmjwDpZhqaAtbKOFkzyC48Fc2WL8kMwJKlaF777SVucthvzedmknZd5
mEpqOUFZN+mUUMqmjckhutTys/hm20Klk+MJKoh8z9tXJtXw8i+5kDLYq6SV+tOT
SJkLd5XEdgmtdgkaHOT5xrqQAgAQDzEdtBogy7lKNYCiT9PPh4GWuy+ypAcMcDQX
qMJoPo3TXCisicqEO8CkGdqu0cLHtGmy9RxIkO86T5up5UxTeIKLw0IfYl26CyHA
jsy1kgSKEnG3/NhskNYxVtSTBmotUDgNB2d9hFlM+KICCZAOu4/M9OfPwc9voaJZ
N07LUSiK+6+Ne4SFHs7XzGp0Z+C8q5UoMHcU53mVVSifqA47dS4nJ/ajQfzSC/+J
ErqVPeqhc4WTTJYsmYueAleYHYOVNPpNuRUzr+kElkLwa7C/CbNusdyT5gxF5BKR
is2SOVyz5A64hjtUt9VVg3FB7+2aV4UIyhQyRqvXwrceUHM4eHsz/TeCOgbmLf5O
98ZMDXXHCEceT1QoMiW7jHBF7MRXsavmbibAS0YSSWq5fP8bYE1noxO9lg8slOrY
M2uwxcE3AKHC5SICi3VstyQGOOu/U52QUTWnmTGMHf0JQK4isZ35eJ48SFticmDB
29n+42E344iimKQZORNeNwHmTaVNMZjkw/SpQ/mZxaI5JE0hX6D/N5lR7/Nf7Pz0
SwULCJnF1bElFIiaxgTH13PDoQh6R9X/vmLQ43bAlMvlgJju+vBq2p23iL+qOIvB
iyEsLabyYuKd3ERo6gK/iBeSDtGjNLfv2WdGMmvCejIAglE6goutrfAd/Iq3f3c/
wHORbx9jJwI54RwEkhwlraDRi9xl8AGT5McVpoLu7OPzcpDr1spLIXynWeTTYv9V
biUYAZT22Qhd2Zhb3R/rHY3H8GIWKe5DyPJxybTEY7RjCXS9mRg5pPh8CDrmaLpI
UIrfkj42F0xaBGWWGdiPsFXSeHJh2ld+/qwhvlIQViufiQ1EjCmdS57DoEckfaaj
N0VCLgG2D7C6G+jkaQCF7eXgf21sejwnK8PxAlA/zYv4oGSAtv9K2VV0M5HxoD4U
q6dXVCxHoA7kKjzCfPr23pfifuM/SvJMhfMt88NPhD9B9v07nV7UjyPQRokxhSYQ
0puy6viCeslLCsXy8PAOsxsreG4R8JCTLqlYz/53Mk+6ucW7orNB27XSwYzQzFhu
skvmud+catpR37SwPqPrd57ptiFxR6BpTwuAICW49LR99KUYQLXaWFXhyahXZtUX
Lk7c34wqgxQDShSlhEuOS/W4bhwXTx93Eujm4Nkg3dr2J9dxUgWwSbCY0B/jO4fV
PfJNdEr/LXInfV1g8n5XkeyBVh3PD0srbIK6S+juvYg0bJo5llmzRp2dZCU/sdg9
mU/Id5BzllAYE7ZttfIUyvFvBhLn9geqZ0cRTHBRkDJjAdgkEwr+8apyd/5p/9xJ
fePS67i6a7eWnT9Ycv+24cmJvg6a0N9rE+/+55ew5Q+/2FK1eqDqu2rEayG4F/d6
cRoVEVFrr8po5RkUA3rYNsFrbT3tzM4N18ikQASSoogrbgER3/SAYQRsT82/H+5o
R+cffh2fci2+xoJ/p+xvRTZZS4HTpNGRrSuv01IXPO8R08Qn3rO/JflZHMmBPWaT
ETjY8tYO70zYHPuXp9HBv3XABvItzEatUy0I9nDN2IzDiL3FBOYLj+jrORxc0hIA
5i5FoZMftbHaw7EhEUsKjfHnAWAfudw7BnFDVxrOliYaB8hWIlzQKBfwhHstdCa2
aZtNqcbVShppFgcHIlBjSKM5XjE52G6CkP6UiRb2164DIMJP4IAksIsYQBiMspR3
Wvhh1q70BfApLHxJhaKiaesaVb3Fo7Uq1tQpHx3qrVfjwLBMWY6uLMOdkUuFJoOc
o4rf9PBkGuBjNS0Fc6HLkvEGAy2tJxI0pxOWFT3HP9zfsLMCBem+qndtEK8mxs2O
oMMPGvr2cYIfPPsHbY4mBnGNr4893rZ8cbc17T2cPFgQsfqu1sasiCtlaqQ2bOsS
gVn1mDOtQfQ1dy+4Rwj4cDELUh60+U6rGsg6R7anq8Ac17v9hAoVx3WdGPvuK5j9
Mo1QeKn+1taplEiQx8g75eTe/DNqkcnQcuaiz73H1UCobJREiUNpS/52n19558TK
XZnkV/QYNfKAp3gHSgldxIQYc4M31Btk+cqQUdtR35JeYVeXCY4heSMy+rKto4ws
I33lvfuaOupmUMmcduqrfrCApCYDOHqUPHjcPqDASuUUWsbXD5V43WOMiKPdN7Yb
qIgofr3i2b3LY9nR9uDnxWkAE4kYQH9FM2Qxwpvoi+DewCszSUcCThKiNxS3mLWu
6JqjG14miR9bV2fL7lQFcerF64bmUYNsNFOWFIaCXVs1VoOwe0MJyHB6k+CgSI59
OOOOOVAkg8cxrAymrCVQaYM2RwNuQnGqmTpQ7fgAoMPLJL4G35oh2E6GWnr6gvwI
itTe6Ftp538WvD94K9oZp6R6CXNC++O0jKQY8r9R+sSqScOaeZHx3LYMOb8PUJq5
tBCaHEP2AA7Qg18atrKsgoH3RQ9ES1KViwU3qWKMHA6muGyb/AECV/Qt4VNOnTYz
sl+rDYA6g8Ercmo619RSXLTwG9Bes0HIDY9SPlatjfPfVtQvnvgir7RCfCT58b71
Vr2cBJLdoFk2/+ekeJmllOxTg0ikX9kejwczYD7LKAP4e8LpyCCS2wNnjJJuJO63
kTsTnzZybPO2+Cb+YI/J+duzw+LwNnBnY0LghmrhPkKOJO5PVzVzDJwoRWXrgM3H
Y6ifXPpcoh5T7wvkRM87vYu89xZwwHb4xVtl6P6aAHtV4AOvctTZ+Uv/hA55izBM
H/gkP0GZo4t0dbQWC9G+y8OuMQA0Tb4HYN3g6AO3AUNJcUnSxSui2M94zjbhItBx
8Y9zKT3PgSHF9gK66iBXjXIKO7v2yDEPVBUuunA4KzaN+Yz9KhbXCvcm6pmqRkdd
ataeyQ99jqZ1J0fQhZDOoD62OeZoLx5kbNeZ92QNYYCfllo4EdmyFnfcqbI4+LmE
A4yQCFbVMElWMAuEImqL4TUHaMhavbge+9dOBCPnxBvmN1p8BKqmbNp1xkCy933l
Sa2aThQmgSLNXI7pcg0G/Oe3EClSTnNA2dFjfysef4snJZsonWMT4yAQYM8gLQA7
bOTAoBpUo3lYvFwvp1wK2j43QEoxgINam1QMXPkM7A8UaNAXpnLOGQQx9gmxIdEf
eAXCqU5/aI7ixUvCrKUp0ACvZ5LsiRm3E3V9Ea4pD/vWT496fm4rCblz3d4Psdrl
CORaDihmHN9NZ+sZ/nqqUMET0mrGi3FmHgWUBUTzgwQ6pYn8I32yS6jQY4oYSFD4
XY2k9bje4sasosFUWVLZJ3217S04BS7mYSyoxUzF75/Oc/PidLNGJSy9H+uMerZj
UsApXz0fiUA5EVkuIHv9eZhta+cfXx7XrzvCYZ6LgS/iXdjufwDd6Lw5FOpqxdXD
DbG28/bhtOnYFjiRX4+GTdMKIvYo9WG3xTqn/lvdRg4aGuSWUNe0FztsIFXKqA8K
aDzgT8bkshNToc8w8SWsfueTkx1my+cxbWOmCJhx/ulvF3Mou/cOcVK4m4yhIIXV
dlwmQO872sPxc0bUSuKrwaDh9AKN5/pEABiwiGgFKlinAXBM4myGAKb6WxY83g4j
9GfnFD/LVoGXSL9cYsL1IBt6JH1rM9MIE1Gc5ayzJm7YYaT7M/p2uDcTy0Kg1MQC
j8S3wIjgXG3v6+A5wS6/I2Y/mPhT+WjKdkqnSjvIdBwFKZRvFifTj8DC9QTtmrHs
SBUSLtsJsXA/kX1/gsiYOmbv4Wji9ML/qneM4ugOoM44IhvAosEv6xig7c5xyQ9i
tQ12v8poSjbviVOV2llT1PUIzTwMAREZp3Z/z6lY44K1MqVZjUYRBTwToFAgrL2R
62F1eaoxChXoI2kWwyjsx1sTjQZ4R4e5OPArJxkrtpDIlcEU98Lt6mQdPoCLYKAf
35v1c7fn6n8Ba2GJQyZ4ml8rNM9cfPaMqgIc6MkHmqvtVQG8qbdbLPP4Jaun1w2d
iu1cr+Ly+V1LAj50CcMCCyiGVfyqLW+CHJX7LZ1eLJj/p0yHow9K5hlpvHSWX/53
+EfFiLN4q5K5hWarixzqpIySm+V36kK7oX3ZtgU/S+qaVyIZWC4O0nliCvcM5VTl
eZNsSJeT/aPCI/jS0P6t38na5U4fu+YHQchyt5SsdP+OS2c8S6zQ+Y3tGwLd+Cbc
Odwk1SUbdsRRE2mMUNbGSLHxbOVLBFg5DQFd2wbOuLHXcw1beeRDJzDzGCf5/zwF
AewBovEIAIg/Luh6xkxky9abrexWERi8k6yF/u50lnuyAdtkYDIMT8P0XnOYda+R
Cw61e4gMuXQhLw3LpzEYHyBJ6z3fDjZs6upP7jytwXilh8/7u74WYb/sGo8eXuR8
S4AR42JFvoGv0dpPRJ89ElybkDuPt++WnIEgdOWk9VBZyEdtXVks8VAo2pTfzuG+
vsUaCZcvh35f88Sfvba1EtKsy+Rw2xqS4c/JhUgNHhVjEdFVrYgk4P2F6ve5z2cM
grFxYJkQkbhEomMO+M2rZfefw3oJnqbqPR1yddgNIsN8XcKd8rDQO4GrC9H15MC6
wXgYRGB5MmgR2EBxF1K/QZI5HTEGdxOQ3TGmUz7OG1f1bq7eqhRG/FATe5PVN0vy
BEUXDZ9BbYA4L+tiBSgsKXrxchYQmrNsEjJmhsnUPvt3JkEl1sz4B6NFaEgK2wkJ
4ez89sy2NcgAT2YD25rS9KLTCFk+PYh7k3jDV85z5z3scUIioyeraF0RbEiRyO6L
1fA9Px7jS0tVKnffMzgaas4xmZCkVUGN8o9wnQ1ASQES4ZZfREtZcATlxy5ceK2v
z0Hd6P1O3NN0yzqkQPIuZqLBF4Pay+RgPTFczxhHzmTUm+WwPzWi9Prn9ItiI1Bm
DoR7plUs+/xWVqqzdkUytbpPU2YZbGuZQwng7pZ4tcw27kV+Bt1G3H26TDnxk2iL
GdScDUvPxgSQ541LXt4i7y0v1c8f52RzCVHXn0Y6IamFZbka3Wb3oyDBt7xM1qTR
mLyYHKUx7PV9+/nh4s3yQEL93gcbg19BUNWtmmhg0U8HehJrx0BO56Dc80gozXn3
gkDBqCXtv4QOhpZop+a7hS1LBS/BD6DJSZMXLHNj8830pnye8o8kxcSu1U148z+x
f9cPfgfJnX+PyNWINX7YEkps6Hv5TyWcCHY+ykS7RPsc4JKOd8fRoEknflJb6Pt/
pkB9HJJyGSSW7MBHfHrmkpW66RsAX+NXonSSTD+Ao0kAXkfrlt5R+xBFFgBVMup5
yTRbEBNL1mFSazxHIz2CuwezS+mxl78cXN85ToYVPojYTzXsxGNrc83qRZuwtCmD
u6SSKSYY2U5zAAr6eCIQiQvrdy8buyvajzbnXh1ZeDJDkE//332GwkLCEDCvfGug
UY4RCMTXbme+W6uC2yL7tqRgyoF+Ntex80EwecmgDx4V3b78/oj/KCaEyNnbPUR7
4wpG8/aAoGJohXLp7m9BXObSJTP2kkWzokCAF46OyPGWLtViETwup3CQuDpzB5YL
nZXEY4VOnxKCTQmPupwOEqtxhCgc07BIQADafC8bY9G3jzAL//9QEiKDdqLQx3UU
akREIg8lSfgVUAU+cj4H4dB40opJAgHsV3Ij9X4SePcQmewgVvZeDXTparr09iKc
QL8pW+QfzwHgR8EeYyJZaNwH3WVUm5pbyvj+oG7xQC9Ir7W9dQSmaTznQ+DlxCEH
9eZo1K7cXec/nDyR0N5NjJI3QNuLuWtve4UsV2MdD59BXxmmGF4ijsEHLTFlPOLv
r3dK9pu/lRsLPfOfiF6y3UzuAGLGFoBi1CBxr3gp/p56q5+MTj5+WCigDcIV1K8K
vQja+WD8spa+vhj+jA1WTWh4u8QLsv4oQjJB1AXQRemdBcB2gSlK74OhP9rC8k5g
hs2GAC6AwTxh86PHzlRGyxgXrulcNuK2983Vl4aHM2jR4e+kpfHqrYsFiFATesVO
LDcMyo9bTtqdUHaH75zhhkPQOWOtndEjbnSykcFG4XsblJIEzjUKZ4Dfyfm+SzCr
8DlMch0PWgOeir9Qoqselro7XfBtASLYMf+r+tKJV261T/h8IQAF8SnkIS8u6BHP
0tMmB8aV4pVz9onTOAlXCBaETXL0fCRVtn0dDXiJ6oHNtffY0dpm22CUEoHpLKaQ
K6RcFZmyM7IgGrUH8TZQptaa7mb3hR1ZGjELANaV4gjacnrijdPj7Z8GkxDxwjee
xZFS7YiKMqPzqTprm6PXzlkOo/tJOaNyPboHy2++5XJWHmP5ogoyrEvcZlp/T8y7
uRyszCNbby7R3iusvmw2J3rJiP7vHePjgUYoOpAt386eYLPQLV+uCn16PZztKVtu
RQ2z4XzMoIovzjb8MFdjKEPOTBl+nQd5s0Gh1ijPWoQcI2rfzJdkYgrXVo91aZWJ
v1Hp0L6Xvf4rr2C4zTvaXwURpOXOoN7M7rJmb8xK07REAibcqAu3os9ffcBlNXJJ
i6HFpu0YcpxPIArw4qjIYK3pEbuauuavi3A6+xiTmNsqCiUF2KbuwuNj+BNztQm4
VNPvsVE3fqJFyt6A8yLSELIyBEY8dXKJpZq+uDcyfb8VnwQKtypfiIbI7BFWDVh/
4CBoaReOwb+9QmFHkQxYeVs4ipD2g0vJQgx4mHQADE4yng9NHySJG2cJr8MxGOpT
T3Rsr3fbVhkOxlQ0qle2osuC9rjvwDJhUJRiBxrYsVI/UndyWBc0yJtSQ49FoCoe
AwsDi8W9eO+PeB6nyCxalMSeMDQtoz3T+aQoo5Rvx6ZpGrCHVIFXt8iNr4ZbWcmL
WKBYqHh8FkulB+LFR2bZ06ADXp0n0SdzErtwmqvMaB6NXTE3RVwwK6icwEbX6qAu
awYTseJvPN/0cxOdYB2YJuj3SNkKGM5LY9lD/+7Kz9453OwQfj64Lps2BOBLRr6b
hVDqJ9PFV/5KpHJShMiqr6s1fpo2rYp6BbzQLpgQLo39cRA3XbHqVyEs/0wPf7oZ
tFKphwI8R+wl0deWsOcwDxfKbeVfpLJUgtsBzrZUQNAKP0HU90GnAalW81QnBrKw
0jo+hoM9V+RT/uLhpeglhvTzuIhkYVopZwBfUcGbcHh7TBP8VryfkSRioPZgoxvY
MtHzPU1Oi0uD6ERXaAPBvBNx10nJoRQpLAlYnDPH20Fybq3TYVddec6lLY7UJZTR
s+miFxdvtGPYJZ0omkJTWUIn0z/JMb9nJwVh/yXHoMY0fXeNozdEn3Dzd+tQUgYS
uQxD/IyhrIHucquRzaZ6Kyc7bbKLziqsLdTE/f6IquRvo2+oUqy4k6UTxPNb0Sz/
lyRGJ6aJbZSKSBs2bUDYaeG8hlJz9YBKvGigE8DvnYjxADUwfsHZe9xEOpgCOPra
ZpDVKR7bZ3hvR/i3zOjcb1wMKXLd2eToQKuCILqSTDkWyp0ICE6KJ8PWF2TzUET+
x0adnt+ZjxthEsUlRXjKBKH9Mkrhb/CFgeLR3Wy9hjug1sOQxB+FItLRzd/og/yo
HlXa0aw2f0DW8x0ssicAQDvxJKMRqvQQr2dz/JfXXBTD8P+Y1AANaCdClVK1QdHP
QfaNlU6Ll1B1JtHeqymZJkYqhJPj7kXackXexrsmzaeozTAsAb2Y3QuhCq1Ov+AT
aJ7csvJnZptZRbZsabYMsltvDpTqNx7CxMg+vw5V2bCq5OIX4AA/2j2fCGJzGvF2
BsXb+d04BsC+95esDTBJIcki/o9r7IUjAsqv/3uCAWqLZ4ZtS+B12ho+CVJGjxOT
szkn3dCYGPmN4ycvp3PiAeo0/TIQUzdMuJVo5pLSEIUt7t1LVx4+BnNyk14r7BI/
LnifJChWaX+EQlznSbdCBpr/LhqAq7EG/waUo8ffzGQ8MbYW5PKgkbD1my485pqa
AgODgRnckqVgpiITiyF9v57UXMt1OL8PaBJtXK5JS3v2s2SERUbu4UcGRiH/kFNN
Ny9gTJ8+zRdgW2KSxUHUZEWaaGzciMIKGOyp/yBIeGLfovGsBetHiRUAL+WHul3y
S9488jpa5VylvYk6OPos+15cK22Ikb+1WKHsgJBdvvYwgiZGMeiXzsX/WNcC9r4D
Y0msEoDDATpe5Qrw9LjDF8CBS5jqhj8GONbATMk7VXf20u1ul1lJoTNo7knQzZ8p
Y8j31XQxIPdthv8CCbcpFRt0SygCLE41fZ53ZwsfEfmBiNbvIgYvV8CH7qG2/1mp
/asl5FKvGzBH7RxiBX2FkscZxvnAK6uDWbxjSwG5QwfezB90dAhiMcgGt19gM9u3
m1VTiS9MLYuV7ADfhiGKUOOTMnD2sqgKO6VG9QUZ9egckUoQeo/njWQYzflKmm4e
NiYoghis8DWM1VsOucVHV7S+ffH08i5l20IbARsUEOA4GqH/E+2YGkvnQmjaha7f
3+uAKcly3hEUeSlpCV+37xrPz7G5iiNDmC5pp81a0AWh7vuxW4DpKg2Gd+yZvZpX
1s1V9JEqtetPpDHva/cXKmXk7Yx6FUgQThecyFxI2RuioRqH/E9KIoFSPVl+nj+T
9p7T5VP8wA8FN8wPNCoOhAH2eXBxv6SPlvbZ1yl8shCaQURk+GOyMEq/yfw42NyI
dzdVWi4GK6y8SBNNHoqokFggmgGWqUbnbcj9/dA1DV4Xif9Q4zZdVfHQL6HBWrvR
YdfN+9YZuqunwBI61qAFHPznXHufpEycMm6tCOtKP2B6xkSLTCru2GFFKTmCLXVj
S5oRGnbhzE0zUkYt74mAOmWAMPWsYBjChbYbhZVmMRQN57baG4/1j9ivF0p9pr9z
AbaK316M0aBwLenVOo9MaHaanvij+IorIkCLKKL00exop+qCJ2KZ7m91Aody/how
zmoPj6l1CffGLglw9cwdvNEEoVMuwimIKvB5DAeVJOL2ssGDE+JbIM746TnvJo/T
APNjYtKcasuE+x012u/ZpATwLYhXuD93sW0cfILiN4Rpwxl/W1zZRaPq26HdNFfS
2KeoRKS3fEwhl/TUXOj8I3I2FWlzKLXeLZPMYDW/i1v2/02pFO19EcBTFqN7A7p8
BWI40gElU2E/vxKw7EL0lBck1vTfe8ADlqZhTbXwRd5LmzSFAp0oXIWoBTeV0YJJ
n4BJtePbRNAL9VSq4iymkkj8EEk9Yd+MwfAEe7BV3a2VrOfGM6k/AwJ5JuPDigHh
tWlaIfHmtgI9xNut/EuvFLZ58pGZMDXl0MdWSpDsEaeKNVpJiHnb18xXnm66zhxK
N8Uhak5uNx7wErRdX5Qk8AVEcDdhGVUkNT1Wri7BZxWHSwd4jvm27dvbEcXhM/YV
B6T3+Vm8+/zKWlDZAwbyxq5KPjYGN2X/nFA7mTqL8eXy+kXqCHsCa8n+t1cXsGHK
fRSrw+Z0rDUUqDUacq7BxhvAJ29EdV7Af1CGcI5twUfzX2ZzFQbgjcJcHJKIYV2a
ciYOYLFaUUH2M4g6d1AdKIX/GpGLKk1ojhnAMesi+L26MhtYeyt3U5SaSSrXdvsc
BggX1vjCNbuKzEMt4i/tvx1Y88PystEBA7+TK4j2nnPQ9Owy2DJY3mwYG3hDMDYA
izdmUYPw1xkGt73tfJ1pW/ablH6boAP4gCLPt+4I0jD94b/jARhENlLfbh7I0W8q
C1oAWWLAasAd1vqXNlAzcU+/hhwU1tkkJAKonwq0x6Lh7HTzYlIfow+qYhNmsf+2
6AM8SPNyAVpn3YCbtMTkwEbk/vuo/JsT65GhhAbGc2U7uxW5gPDwxeyROUjLFitW
0SZ9BVQSCK7Ixf9Hk+kOIMTZUme/51BzvG2RXYVWlgPa4YqOz6+M36szbCQ3j/Rh
KD93eETzc/DkNslu7BIYPAF/kpCUWoIblMVnBwTnwmiJ/ybhbjVKC2I9ob5t8FQ5
m5ZvcQ8y7UH+oZ4g5MRpGMIEad/is+Y2fH2o3xjzATSid6i+6XNdf5wlpfkb3cV+
WM/mgP/W2nwcOjcTR/LDsDTr+4cyBfhxAoEle98FlVpMlmntItW9VaCexjJ7HUIe
o7zcqhx17brwgGfcMqv8/5a0ZVz8UojR49unThtjWegBL/LUMAJ4nLhgPerC5LTt
ALuWlpH3bqb0u0PsnJDKqOAQS6vkNOEoMQO2k9P7T3Hi+Jvd/1GYO34j0RYn72QP
lrAH0KCon7Pyp53m6nq12wuvwEFKp6tV7CrQmRDim61Z5q/RSFCQx235DbCVpfaH
ZdC9d9e/Bbq+IUqYzTFF/LbLDSIgOSmY5ZEZefX6Z/6JmExfV5vAVN8aI5SCtxk4
5QRRlQTHoiw0jh6BloVme2bJSpKct7ZswZRW0Y8/3S2cuDvyheUOahtTRQdp+Dqe
/edhPeOL7+aGCAlXVgiv79CGEp1jJuTFnmewhgZzl8ph59nJRvTcVZbIxc1u9pqs
IFZqkRe73Le/gWosAItL6pnCnxioQPYojiM9XB/bwZuGMz2LSwdqjMKWX/m86u0h
QhrtEOFkCsJT/axcppezqzwG5bWBIWj1Tw7GOEGL2nXr4wFdG27DF4Lb4FxP0pWn
4ySr4dJ5Ek7xjMI3aXpCgEWDpnbZtlxr/Fe1h82TiIJdMvPZD4u0H3tcX3WCDJzB
LcQ5nuISpQlYNv4vP40M8MQ+QR/w7+lcoibI+WVCeLxB9ATWCfvtU0L/AuFr0AQT
uxb9Vrbn98r5v8W+JboK3weCV8cpAJLdFEasAKqRZ80aw+OqcPn16eXdYzygRwP5
pj7EYfyNop4pzPY+4nthd0pG4StJujJFR2Rkedntm9lzOD6n4G9Pr+TxmnfsNHfN
AbKw7DMqmrNl9K5KDyZJCAZTWPA/HAY4TDyYqzaU6R+QRNsFxkTUEGA0Drnl2Fz/
N0VUUDMtZ1F4f2uWwovOsxkc1PwyyVQuYZ7jCnu3N8B2kmwo8CbCJCFli5uU8+rh
8DZDj4fNWd7lUGft2Cun5qpo6atIzwLW73ueTZq2SF4hAcwEFL+JIPlulxMhNXZ4
jWwvuhb9yRG0cRsgE+NwQCH360GdNrNf9JQckXBcxXFgK+Pl4fPNaJPyy5T+zfkX
RWzYjjU4LN5O6JtkaobFJy1/KFUZOnpDAgbCRoz1dn2APFa1c2qnYSH0NJ6r3TjT
G2nyyR/0Oa6kTghGgnG0BPlzepoxGmTyUiGPGhB+UN7HpN67HuBTeZtoz7VNgeR6
znyK+8Mho1M5vf98PePuE7KHYvedzK8eCzsJUTj1lL2pEurbLsuxxn4pncV3zwzc
UQL9TrOlyDqa5mDO0OCwHdP5WVa3QNFGLrpSKW1i2h9mE8xQ+xS1BLapeCrLY1TJ
m8/ixUUK+NKWxeh4EzKlXNiXPWB3b9XHDfiiRbIMIqYQ4b5TkiY6jEWmJSnypLPo
sekGVYlammkWZQO6CoXTyvdarPMi3LvW3VUu85mZ9PkqmGLR2Te9eUCSORIbLpXg
E7VVzKNCakh1PCDfqeHqHC1/2gGiSDtkVRs5phr0SL4Eq2Cxoka/+N6i4TNdcsMs
fiAFXtanB81WsiseW34IN8xATiZz2+KglZ68P6MvWDNmfsYVtffoa3mWoWsaAw6T
US9h6jHL7jAu1N630LOKYgrsJwUNKC/yBEhWGEHqUo/H6t567Xlb8lQm/nqKkSbW
OaxAxPJn/y4KbAe12Ak0pwQqjRjSzK5sJTD+XMqHvGEZ9ctTpgES30WJ7VrlEgpr
M8Ms/esNsQuA44kNdqb53WeWlxoHm9SF0aswWBriAvmYSFVvOW/ROZu04NIgsnz1
aQDx9+Mgz2uqj3yNG6bOs7cAQS5GLAciumvmkCRGdeazgqzqvzm6Z7D/seIyhCw3
6vLk5OK/yagKIDL/QiacC38DW2K+NkPElev9kNQ3O1COPkAQ3KxSPzZdxbDIjF5J
I2F6gPKXc0xctoRHeZqm/xb+ofTv+4THJykl078DICqYRvRaZPp9uxE2ZETqtaJ2
+klPNuwrwoytGkK3zAv3m/pDKaqZMAXg5SyIT0G9znQFgoC4xCU2p0WNJ62TuIBn
/jyo4APMy+KNoisyetuYdsEDhhCRQB6Bwi4ircNBYmYaQZJlRomLnumZ7g+ePHYC
Gd5swua8qwuT+tv/VE0dalxIgWf3glgiWsK5qFBtYTO0fweZSCWt5n01PHStlfdV
7GMPVIdMSPUoQMeKf+nWuQyNj6r4WOXqh6LdytwMZ9c1wsOndFLn2w+fAMJ8FkLI
UPxd826vsKYY7OQpXFcDyWaGd+DMXZjfxpmhm/Nd/qHCNgKUKhHhBp9Akh2exlg/
OYmaio+FnGzzilp1DVbWXfcGBc6CrhJtQM6trykTWLxOy6qdh2zY+L+u1tJYGShn
qYfIxF/DOJvaGuDETP/9CBt0QdaQwG6dKn87yLHHZHHj1dyf6jU/m949eW5Fby8M
VcqEeoB9DbJOc8bnclv2AvuO8sZoiABMziFs6/YN9An60XG+E26VAmTyTqmzsCPw
vhE5O4mxH9ggVWKDvvI+G95jePFJJnjlhXn6lqc9iFBTWI+k4+je/jZuaXg1KdVj
kq5H24wJC9Qm46RKhdtblcv3w+HiJsfxh9ES3CpF6KU7+eWUQ9ntuRSkS4F9xBId
55bMANEu1OVqq0eMOc/GFsaSqP+jL4gyXdk8pAjtgPfcNZ5NsurFvEiW5W3lj+JL
a286dJZb2cBGZUay6e8rXsN+s9dj3pVtxjyTp3A6ugcaPNK8KUyXS7J1jyCgjkQi
nY2wZ/6ReGyze6T9jHU0Um91oY/BuYfrahklPQnlJxjQjdC6sRUkU/Sp++EDmzSN
M7/Cw3stVx+lL9xfX+OIPXpmMXDwwHsu61gA9MY00ErZROHcQGgBpxnmsFFtOtwr
3hCoB3ySJ+br+SGtGK9I2NEFva4Q7cDZf0OEbAeirGwAEIHLsKjOn8eKzR67cUrM
KS6BREUzKd2MguetzrC3D4jUf2jnWmnfom7+ORTMJkJNpvA74bnLpBpG+GNTp3j2
unBFryw/99mMAyFJzR6Joa14vzYi0cmoa4sSQXd6m/SHZCeC7ebYuTubtvB5HHlK
gF9o8b+08MZON5Xw3zbH8oaaFAJ+hZmwiWtqucDK5CNy3PfIieD/vbxq9zTJEhbO
T8Un7yt+AfoIA/dYWMXTHvHQhh+ukIDKZRkjDNEclNi8n42D0Hj0WJGuCK++RH9h
ONjPROGxh4AtCgzG4FutNH7ahrbANrsERxhKmE1/WXzcWPuz7wZ3oLDSYySVRj3G
HcAZZzklj/CqrKbnqfGS6az6nRrgwkTPtelUCAO0OktYuipvDg0Zt9Z1sZYF0Bju
kAzI3w94p5ezBwB/q7jClq1YQXVpM6XWwXudsCWrnqmtEFf123SfzgXWx4heeVDy
1m+GUImHYfaBhDuXs1lPRq/FsmYMzKH1l8uqoGXujUOafX2xIHSZQ52OAfZYopzY
ITAO3D/qgxLfn9wDW4L6u+4wjJnuX1fRoyy9zYH5oA5yntv+TDi8YZN/1wVFbO+J
PeSyb4fWW03OWEmW2KmB1pKhICLRwx3TFdm8oK4mgBYY1Zey2eApPCES96Z7quAe
lr/s7IW1S6M+3RNfOus+o6Gh5OGg28bTivAuUbzRgU8oKdlmsTlRiLqSV0ZZsYfM
/fN/7+Z5CXfLe5xcK4TBDyuMdHo7q9yEZhWwOtUjoUmMh4rkirstZ3IkPMY1Plrs
mMxL0xctNOiPqZadgZVdrP01VgOXcinBMxO4X0qilT1q5DnB/CIcIe8fa2/hmIAy
qAUd7xRwiCKnelHFddlL9Fa3ijPsgeZkYHQ7FO6+W5m1zxxOgsbIZwxaFDlTnae0
vQR2c2+q1Lu566Xz9OVE8YhSVnOg3MRRnf8bYOYfd84XQ/Hb6PmMVWzeWBl1gkR0
ew9mNucW0YBdYhXyX5wBKKupDVtPQouFjgM2I/qtKzqpv+YAhWM7zAPFMbhD3vDz
xnyq+NwXxjsbFTmztHZOcJxPXTz3kvpqEpi2AYlhtOIsKnlnKILC279TlEpUAwN+
aOOio6HNNr3/4gsfYTFvYv50insF+oX+F7fytBCgPklBLaVvj1P23sQ+bYE2hGA+
cXiIPuXiS4KhkJnzsQcUEekUNFFMtaNgippmEQ1Io47fODTjLmD+j4Tob0kQZ8G9
1KYmZtA2b7A35xEVBx4appM6ClPE+NvrGkZxwvbojkWE5h5uKOjMI4oK4ojUcGL0
FI3g1WQiFkVyEcdhLQlSi6DsYdak05S/dS9yCXgxqwm71M0OltgnMREFUslw7Pbi
/qoufk8xoL2zFt/fhZLO+tyR76LRX+IXjMks7fSO1zMsEnXmGkwlo2Ar7HFCzJzV
W4kNQaJQ3PhhJQM/5c2EufxewEIkQf/otqXOr64AgNHUB2CTMIkYDbfdLtYmaFMm
PeA64ZBveJa478Z1NOyRgDZJLrDdDp+oSbB+XjpmqSUIK63w931bZcy8AL7banmQ
wzniQFMEgLHwvGkEdvqJKsKZw7OkMObHd7Mx0tsPQT2VCWVyLY7jt5+wP7mDrxL/
HoLdi0JhBeTTksyMwAiqmqfirLC4X9yK+5jL8rJaKZB1iMHxz3KgbPRqRDk/L+aU
j6pVUzg+6Oanvl7GQJelXaiSRyeVUHpPp7VGsjEvlhIGR2VL7osY64HVOEF3y0PP
eKHC0jy6m/HrzutsBSdBhtRDcQ/PKAWWzXpcwBx35fWr5jCa8XM6zP+ji6Cw8Awa
+vor+QkOu+698Kon6XnAs9mpT3JZ67c3u4H/YCRavLwfvdvCmpD6FI0aVqjRLLdu
tjP8szrEBDIwDPQm5d4Hh3DOtafru4a9spD0bfVAV3GUAEtzRmkFEeJb+PrPFrQd
yG9xIUVyKVcnX7RAPs+4r2JPAFEvXhAchabs1N0Pm/2zQfZbYATLP713Wz8+lnvl
6+XYXGBaK9poEEo6CbrRmndhx/GeGAlJY8J9RQL2IZCJoWxeQ+PE8+iT5WcEEcuW
3z5Mrz+cQZUM/FhC2Eg5eavFb2PBlyB9zxh8pXO5cx3WOgZuyRwPhviX0i66pgsl
QRkvYZowsZS7qONsDHuDbnJFtD+3enx8ijqq/a3DNMV7lggASIt1sdqp3j2tHSVo
0OUWHda+ojwQ1J6OsFrnnPSz9ISYNp92iTQNnGo5mRDihVw4xpN1BR+p6cCdlIhM
KJK8guko749tduoJR8VBLQe+gvrkqfENpOzuOQ4XPc+X9boHc3TmZ5BDrnKaQBec
GsHR6/gL3P98HxbSUznmq4fdlTWQYzViW1vIIaNO7TrqsvAuHVr/PI3PQTwqzzXC
NirK2vGofGUaben9eQ/OxrE2Bi7Asejf5uRSwb2re/+MOmYoc519poIdEaN6kHs8
dj/4j/fA1ED4SAgrjkRSW6y1Gixlo3RETG51vgbpgF0rSvO0rIfpSLgHM0VSrr2N
3BSirELpMzvRkfdX8sBfErD4G6x5XGLxLIaq4CmAQWd8mA1wnAF9uIJ7XnYveyFD
pKmTtbjKqfz9g6cPmbb1czhOPByigsQNZWbVNzD3bDgaQg7j/aTgvqQ5Aymmc7+w
OY25ZvoZ6L8xwxITEUNoiXbuZu1wvEBo0cMk6LLfT/TXJWgjCen5movHqxQtsnIS
BO50pW2kUcSCdD0eMpe25Majf1WWLYaaGQOjdXZX5csMamSkMG+m6sp7cX3WsG32
fQRijE4pJJlUZck8egCQJ89KZghAJy4V0uFcNrx4mdSHq3S7n1RrMnzlrI+/GbeL
s69PHV7XDQoR3ubqXHM539AP+ZOWTDEwKQk5//T42XkhB+iQheXz4yxmBA/hjoyl
+WItr/YhlIKFAj2X1z1g1dJ94lKm0tEfx/lgUUUIgLTPAx5sbiAOovfTYSq3ZR21
yVkmLBzIOfnUddwfjTpX3Jos/v4N0ToBFwNb9ElC0MeAOESf7f1SY9WJ/YAzUQKc
ISoMr2pJ1dMnKijwfpq98tHm/6bX8XA6NYDZHtYljJciJWQkn2ND6MQ06HkqSNYF
cuInHprSN/rSGiHBHweZ4xIaOMDphmXpidU8vmYoY5AKkDBf0zGD9SM6hZ7Ia4lf
1wmOzaVz5Gxdh86eofrZOT+JkGU6V3SJW2N6tsL5PX2nyjZ/66ySNngPRQfFi5Je
PMH2HsKYC3+ubuAaXpchxmmOKGWaKYeaWcZDsTARZceIiO5cjagLx1a6hsKwF5BR
BdWboL3VaL6m2kvNKj67xfUS+Hm1yGGDuw/yKCjocdiYO/7yvgnFCZcm961bN9UL
X7xM2Sozr4oYyhSFlgG/cJEfXOFYgtc+MWfzjJwWsOeC7lsFrEsurNnYPTDZbGMd
pVJTU2Bo7lIlHzqHtsD0B7zWtYmRT9tQf0NatBzSh7bwpxBSMiKqeodfevg04NsQ
8oYwxSARfIB0N/GvMEN3yq57vWUViCS/EsdxP9ifFGOqbcpxcTd/lcK4xCAEnA/3
eE2JXt9DQADH8ZWV07/UnCFdiWJG8xK5vzU8+/3rwPxTqG9vGpFQz51SWR8s07XF
JDXq6TZB8DaltAIjhx3ekElwG3bqcf9qpnacRT/kRmEN7uhO7AqHAl6bUPtPdnly
sGMdGXjQT+8iOlblfzxqXumBvGI2Kumt3H2Lx7bK8VbRk0kNr/H7rQ9ANhIdC0qx
j7OaQ92J7uaDrwktabrJktCgDivjzm4ENAruqX3tSnHO7U7HIMGqHKSmn2jjDaY0
ZQzg5Ieki27rFJOmLyBKxBbV5dxN8pt68dGnTwo3+euQr85nBLr5/2eqOCt8hEoB
7Kjde2BsQ23tbnIxfepOGc74smlyXZDGkv+f45MSQuDhK319hI1e8QeJlg60MoPL
sz3UKp6zb3QrBwcwgHyRxsUEmHb8Vfc+NB67ZZVBQyg+UevCmQMw2+xbmzgVQH+N
DvkwpyvuzlytayXRi3cGpui0Qyu2AJxDLJtSiRo/f6pQDKeOkqyqyr+BfQQIS0N0
II8zFC4P04iZZCnmz6JILrgNZggI5t+tX10NIoIqNnqkIQNnHwjnb8SC+hQuOyIi
O4NMu53hLVRNvYqxDFXbmv2QDuPv1f1bH6Ka5Kn9ftzNuf2dzi7euzNefWUuf62z
vVZEIOS9AZmdRIDB+40yB3iXhfaze+iqXq+GXpK3MrC/1mA/DytytjVmrrqW+LlT
1L3Ath5JhdMl/G+8lr2NtKgqVSAD5DifljLgS1piNIf6W9PxAQCPje5B6lrjvUtq
d4ItJaPqC1mt9xmumxdDfT0cF/C54b93N7BsILxOQMP/hrUiaSTfY0rf5wxxBQGN
ABb5wfvbrEXqi0r4WPeFid02vGt7Z7uVeGfqUfidng3qfrQeoCBebtJuQlkS7itB
ljAJiWYnODQGF8K56wlk8Gi4XPczwA8+cSEPsbuTS3lJc2+AkHKJ1v6hmOpfDCSn
dEBS9XJrsSKDl5sDo+qWEtqP2Zmm1pplCGIPSnJzf7vPq7MSLsvyqvJnbwDOqisP
XFuBnqFHiLZBV2Q8DZLqfY2gtVtVGwKec0MA2ae3gGMo3o6jA2iVBsIPvowxpfEp
nTuG0JkEYjpSINAke0dB9pc1IZNvFB6RMBS4nhPsCg2L9632x37Oia++rA3Xj+ki
8UN/ek7871obTmLKr9tvRqx0iWTWDoLVnHojk5VACMmVDZuolRl0kO3LiewItf/K
UrJT6eMuYeBpoGrxRJu6v826XY0bkfprfB4RaMQZZGoqsOBaSMVAUgg8EijZ7EBn
wxlv6x7Lb8sH4KPpsr8ZkCKwBxSbQLsfgXhrZIb/4zNR82UpKI0U1+PwRzqTBs5U
VgPNsGZnMwEqYIL7Q6kmILQcGif4+6YM9D/rJOB+3+pVFMmC+UrttNdX547g3pwV
CU80DCIpqo+Sx2UsA/1m3IxSv0xw4rm2JMmPRSaOmYixMJUDn5crC30A3w9TkMnN
CkBKyrldOHoO5XZt5F00g37vj9guHx8lRKkRMy2QskQ+qyPxhREdZ8AOinuP8Bp+
clkJr0v37BUiSpdXNaaRdeYQEUJbP8jCxvG8sqA9KhBr24yoHyNCY3Vur25R6q2z
7g/mLpSQCInPCDTZ2t0h8pWQ8kMbHMRZn7wb+vh+6yBTm98x8VinrqKlQVzgIL4c
DxFjIWnonmWBL0r0U2VXrrXQGdL0/LZO+gZIzodP6JZG++gqKKlnkETlkCuL8yGQ
ZIbK0ZKNaVORJo7hbeYzmLrxUOqLrleAO3Hns0SMPAqRiWPJzdXxhxSu4TcSfRb6
Lw4zEWmSER1BDyyfPIAD/kyr+9uCL2yLikEHQ1Ol9MhF9ekIbfF9EGl4BGXaN8YV
6WNySOKHqoGV9ikk/kCIznM7RN8QQgFnLmWt5EaZL189TAseLA82qvPCNLhY3bmq
jzXd2k0aZ7MV3xvCsrFMoVH1GspaZqf85bo2fW5//bTs/N57eOE2l4F7ERlV2Rlg
KY8F7QFCTrYvHUazsNa+gp0AGAVGPgyzZFFZhW8tp0Sjk21e+6UA5U/6duWVtnh4
WLZI+6eNaeiRhrtX/+yri0cNxboT/U6MfQNK+mJckT7LrlobdG1nh6KGGfj7cwgE
yno4QbKzuCGxLLSTKJqe6vHphAFKEQLJP8LPo+gqCwBI3CEq/VmiLmoI5GIUnsCg
XdYdYGlBJYwyEzjxf0m8bLf07Vo+ogv+ueR+QjKyjkOI2OZJKiV71Im/UeOOTIfW
HdL6aL+ONo/Us3BWp5Zicc5Gktl+SvRsOeqG+YLCtjbcns9cHhmI5HJ7ojegMT5N
/tYUy9/KcMve8YlzGyWqd90UjiWUvqDaCNzlPEkXvSkMf37Gyyf1OB9htwd+JKFi
U3Ph3NQe9sFHpsfItlR0uUCnVl8Benz2J2M8t3U5gGMZfqB+8SIbF59aoFG82frt
Kqp4KP/1GkB+X+JpHVbVQxZ4QZ/HU60tlpHDZk3NkCW74wbxMg+xVTfEadQ+Qmdw
+7lOXUeQ+Z40pWixjGxDElRnUI509vuB+bbFEkcVEcfcb5b3C18+hGfiAA4NSLQc
I8/vO5v+7XxF6rJe72javO2rWJxxOXBg6KuuTcq5jBQTae2U1m84HqzD79U2GfVr
r0pyd4mthX5dF7AxDvdc6iWBonS1vgjV0jueJTDxXZK7NSqBlI4vgwtFbn31xf8M
RhDcvTwrJGMDOOoqDZb8UIZWn8z4iQBOlBHuhaJpDGwjNMKX03WOxgqPT5G0ZHoV
Cm5NZInP8nhMpMZvrfCfFWGYTGUHojMihJAY3XlSudQmR00NfpwjDV6A+ylq5XyO
K6mRvHxgdLxL+n/qH2f+XkBujGIc/myQMu/oA6cqXPqtDqZcyjR8qKRV67f6+9F/
VaASI/ttRbVbb12r7g052IsR75NSIQmqSuAGRfhtxKWWoBBAx2ZXFztVMoJKq9+3
9eWNaUXlEdN5Fnq2+3+VetPA62WJukNrUkUpIl59DG5Sso9Q83Lji48/0eC7/r/3
tCqUPrGeMzwiMhhd4dadW0Uq72CpVEPNI63oVv44G8jTRgInoiGfuavePa1Xq001
ypEx69o8qjP1Cav/NUUGPKOM7C+G1T0sdLbKP3UHjMlkyYlT3ZrAD3I2ZflUyZoH
PEZnUvH1Czw5N4BvGOSby/mr1YUtqpP3R5pPsq5jEK8jL/F1f/CKWtQ5yVdznvPw
KNltV0mlEInqArPAXnhz4IfIaWBb/bcPm0pf9GqAYIuhMRd97WEbaR/nsBSiL7yq
pYb3/esbhGBXftQDGDvmwwluXYctAS2HRagtn789q0XeFnD2KydFh8MCJY+W+KOt
LurONaw7xUzxeyq6jvuS6H8FK5h97wNbLyG72VoqMBtEDVQYFpUw/EVPIR4RMgWt
mhlrc7sibKtd9nCoILE5uqLrOjtkzvW8O6O+dA8DzqeoPCp8kqmKganHJTy2znlV
20OqK28JVGjTvFO9C7+1kssZjh8JCdijTEa+WpyDQcGoTfmgM+vtaE+RitEu3AZV
1+zm9M7Q7kzZ/iYc6LiFvF/dNY6dpxHn/VjCz1anwghVqHQcJ4GiXy4eTmHLZ0ve
IaEi3kwpNMevm6IsghTyaNW/AMMwJ6TLIfJEa41Ddt+SlaYVLh/5QaVVktx7xkhe
YSQqKKlInRQK+yQc4kAcwc6kC/MdbcYoSr9Vpd1eqsreVEFujvzoHXw+BX0/LTxl
x9bQZ4SZ9M8omJagf2u3x6SfNFfplT0PyusY3lt4sV9YOe9JFfQVgYEZcK/4SrwP
eSinn6D9lP8fwFL10Bcw+NAzZ+jaGXPavxnM4YDGQHGdFTsPH0QYU5y2lTutgzmQ
LDNYQtHvSIczuUEuN2kQXG1M8CcX/SUCkXPheN8Z/JZQZU0H3UU6UBQhFhkbx5Up
+JLNmSJzSmbZ/x4h3rpQR7ZQEmf3sa/J9jdrUViP3dcf9zuma4rIxC1bZH3ygXYK
Jspd2nWeHGiwzMAnBUZgB4KibNn302c/Mg58L6tuzzT92xWaXC6pStB7tJLFlRWS
yH93XgUXYOqW148R9A1Re9a7nNrmSm+cd14ZgRT855Bp0oxUt/5RAZLvmsZoY7lx
yc6hGxH2J0tHJdxFBNLHnazQ+chpJu+kBpRhr/7npeKWT0DMAtMw6rkbu6lL2RU+
IwxWW8AnJphoYmRzytXnR/t0MUb7UXsOqqcbw17IP755/BbhpkpWBn5RT7ubIX+f
gARtmfNkT7tohfxIjKZ6OnahDKOm6bdLek9P3J5Oafr3NPP9aqhT/NFJaqvVzKOu
fJLuOH3fIAV5Hy/7BRwQ8VM/zLYdxbDwzd/ktrndYv9bFMZxlqs9mHWNcFkCi0ho
RZ8k8e1hr/BB6PTYA2haMj4psGEjW01HcK4g1V4KMmqdI7pBvz79tpqhAzxWa3R2
bSfxy4DZ3iIYxeCVzw+SieGOCqBX90mIdS0YomKQpnM7YSMdW6tToX4tHwhvBOOq
T1YZ9l44YXcw3+yDw+KN/+dc1mQigP8j/BowjLgzXuZKmeA2xMgXkFBonxa0qcHh
OgNLZ/AYamX+HqitADLojwb8rwaRikpwlMRRi/KrQlcqyx2RZCnFiEzKv3e6Yiuo
KOJ+dHiHXuwWcDpoHbFu8w/8KH3EWSKQe2EFAnAsNyeaIQD0Gq84AX0aIrQ826Es
gTtI6Ukwzrq6V8MwqvAtb9xliKxqJzcSVI4hL6ebYNc7nHj3t08Hd2hVW12l4rtv
dNzYBAffIt0/2ya8Z6C87lKRnnAUjwpgW5NODeoQbk2iKHuZtY3R/l99IV1upwS8
jB5fbNtuElIMIYaPmvgK3HmkOyh99Qsi0DBO3+4ROKjTpImz2B+JtubZ7TM7uxg7
EpolyFmC1eaRbwDuD9km+ePQMKsT3pfGEg1gX4SocJR4CEXp8tW9hSQffB9vdI4n
4wDrZOWV+EBriJrBJaUKfu9k/L9tFf4Juf8gP4XowbJQP9k2vl+uXIz6d4tUoKIP
L3GGvxjR0Z6PIIaI5fG/Ied6zXTrfR/3xtlTw786N0PdNpCWozbPy4/TvlVRL2U7
7GFPJTK5Pq39pY583BoUpoI/nwVD3C5FwASTh4ccGfWO0wW9EPl7yLw6hI/PWlvc
znlQlooGwwK0s0Gj6v+jl1NZcJgGiB68mD5BY9UZAyvzr2xezgKgnsgGzgBL5lxG
uaxsoS0YspK4AzZu+WrMBMNcNxgeZ7ASn1wb1HYfEKMLBR+n+/KBboczviEo5+we
UvH1ua00fjtm4avjoxLPRHnI0d61vZnyO8SHhToGgT2thJzrvgvQuzt/br3vTLrX
yX/s+HRyLrMWkaU5705viuxZ+KEw/lEtgYhRRG4IXRAO69qiJw+S5bX8lnKUo5RD
X9aXFgqIsCbhQUjUdlvluvSCKwZivVdvOmRO4oHfkUlGu3f2wrXu/lSdCPKwQPGW
oJzy71ewC3g1t3dk9rlD7Nff4HHKwc/mf6EutjHxHd36Q4kirlfPYrtD3oFce6xm
wp8+BqSkrVIfRXXygCBF6rLdgaK01dP0nMkeCsR9Gd4CSBYOMR5SE21yKTFh5pvT
IlyWP5tAx/ZYn41kglR203eVer6U6S3Evo1PTZgOSTk9v+WbUkJB5KGlkYe1E0Xs
jqVxGLQdywm5mb20I5sHpM3mEzx3qzqgNMaVvs7yd7QUjxjeUKgaTkusonS62ROi
GrAq2QvV6XIcjaRx3ERp9yTiR7h6P4dlzSmQ4H9vb3ff61XCNpM6TpZMIj/oMn3A
YBjeJi9hQKL6/Uncq+w2GoJeLRIRpzGO6SiIgU0gbhudPA2tv3i8RqoIHLETLn8y
YzHobjRf2V9havt1B8PlmPCeaFlfTFnVVtBmVRWf0dGvbkBSq340hMSCfjCnf32o
a3zkO09yDXzlMDk5u05XMz1l0VJKtufuTO0Xmmc6uX6/ofsrHQ+kfKx1L1k2LRu6
5aywS4CGFZJxY5khICnYAPtNkwweZQWJgPTCJ8ehYvoGERa0wd1rlzQLphBvuGmT
1356i+p8Bqc5yUP6SUlR8dKBDO7yA8giG2B+38pxwJZniQh3Ys+4itZxN3IsROEd
wsZLHeO7QBRmPpS6RgKMZGeGi63Uu2KnZbhkWy1JG60KWz21xsFvR3KJThJCJoUT
32tLwBzSQUVkhnppQqAFufykrLzRROHY5nbnboIyql8UD9u0SNg8J7xQGmqfHBTJ
8SyR9RtB+Q12QqWMVXcMwg8I9/VPf1FpzFKARfMy7u7VMIYYkX8RiQO93Y3xvnpp
OYRBTD6QWlJMZ6BUdsM6BxA7xX3JyEO5AcohoUJnb/6MbloU8SMK+/PeDBGv2vXS
hW/kfbGgdIjb6GjAmuuTJHT0+KTBAiJoYMM3m5xE40MN8/pMHPaSFvY9LPu+BwdH
SyOGABYJd2pvz7TV8drKFO95KO2ludnww4ekN2IQXmlLWZW6iB1ETFkDiW5EO1Q+
82EZHGmKmIKpywxO/SKMEPtIencjFjrM6VL+kncVH0CWGSXub93nVAENvxtyEhhc
tIc6i6+zvwbE5RbNuyWPLKZbd/kDbOe0Ob6888VBl7XdtqPpyCwbYXImNtLcwWqn
GXIRez5kww3sM3IG5TnHsXEHgWSI+kCkvjiVOhA0SfCFVOX3q73gaUDCr5YixBQo
SJLrx3uJRF/D3xx1NyWVd/wzrnC0rd+jEAw+pKIbjlbADIl1WZWttrrsmU4UQg0A
3Jo5qhVKyz4FHQ/ooeN0UZ7CN8ftBO5JCOKmFK5vOpE363n4ojio6RPhzUfvfrgE
P9nvb320cJRRhLGD1rV6JeThih4Srp0enLkbOc2cL50FutB+mVhgyr4S3OdTDIoQ
4E8wcBlhvFHiVDLhJ/bjCiI/3P9/Xq22Nw4F8qaaPem2Y06usnZEeQRGV3BNXvxO
7EsTdadWh6/inuplUsPI4+6sB0VhUW1V4+PAcXB/WqSPIFjmbytbgvLFLVSki3zc
9AWgkw5xUG9q014+iTSCBsiRH3+cxq90nyfAXXdAg8vcKORZuzZpQsAE2VRbapHL
fzJJzTfAgzsx0x4e0avIiv64pc4DSJwd4CUE+g4qPISaqod9/SmTrtl+80Xiqag4
vdvDk9+pvvSf/n32f3GnRNnGZgLXdcSQC3CLnqfuG8rJBlw5vu+Al2lmrd4fi9Y7
LG0atKwgY3Iq4xkUTdtdXGGut3DnsaPE9xpzOXCDJrVP3muAVpwJzvi2diXeRI8S
9rCBAnwW8cXPdt63XQKjRZgBySAvjlzI/g/v4BFDHoUJ6skx5opafOaud8D0Ss0u
npsmK/Q4MlC/eAsBiRk0pNJTF+Yqo/VZzDshQsIMAb72+o4wlnFeOmyvmDrtxVU2
QmlRgIngp5hbX5E9/HkOp9kgOfbSR9QmmHu2Li2+S7R1x94NdXWA9lpcybumhKbZ
drbdKNhre74ry0kGsAmAJSNagmEhJmODDoh/Eh/kSPkpE+7oJCTh93aX4XeUOKii
qjVrETQXR2JPuM+DH8LKDSo7cz8ZW4C2cJiYA7N3kP+qKc/b992xdWsl2FcYnyTp
D+8NkR2pct8m1rPte/OQTgQXg0TJEHM4TVSSjW9v6BK9cxvYYwhwB7pHZbuxfQUJ
x2cLpAZwTe4gxSb7NiQO5gmKs3K2y4l5dbGFaFfa46L0DkftXSXb8AiwrvNM0oKV
IsxR+JHlyuXlAUj/1wXksce2B++8ndMOaxxbp3bv+uPcuo4ksYPtSz489eYkb4fp
xXwHZ6gNXuqAIxDLCNcH5RF/RopqS0D0QauWmIoF9uG8cpr3bfLX14gTDRwpm7ia
C++c8CdvGK+1G8eEjBJ+2BcFWWM8PUurh++45EVSGu9mQOfd0FFCl+abq9ywKtJV
NNC8EoXhrtDt5dhJTDejdGkqDFvTxQRsilEh5VrdoN92R9AiKquaVFdNJKRy6v9y
nnpWJTpk8bqr1LRVpO9alajgbiH9CftBJ9+7sxuBLQtXNOc29dImSL1X7gK+sphU
e7wqcjvzNKsu/ClRVqYdnPMGV/HzBXWd4xRZwRtD4YOlLxnH3JRYc8gJIgFO8Jfa
bQvy6PSm9kzpka+uUqpNhyZxv2kiFNWWjdi7FzTjus3vDBifisfIRbouxTs/eyfy
r7D927yZ8lxPq3KpKBwA25C6zLebJgjILz8vleZFH4BCQcPdINeuwHwJZdgUW8SM
wYXsYwJ+6669kaKCkENT3QhP/LmvTUWCzqWkHUjuKDqgQZVF0Xim96PWUaFigQnx
8l12O+SbRPGp+EEksqJXUY1DT6o03yFAn1zE5fceA3XE89I2HSurHikhEVtZ8yh0
TqNd/+LRdjdG+IeBqf4aOc/BgH9KAv8EIX/dSKA0JgxXwN+jVumUVSlclI9+H0oh
Kj92YaX/W+nlpFOMJirU4o4FsYhySSeRB7wQlFLPCA6esIZZ0/8ClZ0i2DTFxlKK
HivyHkSwZjJ0plyuHetgcgc+T5zNfMmvjp09xgFkSzQjSWxCViIak5S/jEI2pFru
hfUQ0xbQxOm8kJocBL/TdEL03z52WCL8g7ERfgBYmXtlVDzBTSvw9iiNb0xXW+8N
5fTVixe13oWq993wSGxxqnSmljsA7VhmYRKQfHP41vsk1wZFxQaJHOiqHK+JdLKo
S1gEtxcsiEtELRevygh+8Ui0bx9l6axFSof14xHKqwSccrkhi1usC7k4mdPGZxle
sEcQ5NrUYjAeDXaFi/D9BAwUpFQ4WBE+rbOr1T8Xqdh/+IoaUimOwTFOGwFjccwY
4KCUxF8edfLZT9qJm1jlDFNrSz9JlNBKCbmzqPrHQEfy/Wb3Afn5mQJAhDYQ2bmb
eL3bh20OVx7Xmpm7kWDnsRGAyBEB1Lbg9J3OEOr4nrMI995c4QFABEASrnk/r0PF
i6wAF32Q6S0sRKVdPqp3oxZgwB903gT8LzPMv+HFAgy/ONDJda+0oUdB9U+V+qgM
7nABu0YmbVg0tT7nf7cX6sYeyL+tPL7l95oR/wGY728YUD9VhA6oID+FsuSJdSVY
NGmK9bE8PK23m2Muw1LnfCR/PyeT6Q9F/ASSA3rEtUbPYbrn2QBgpo0g6ZyKdTMC
O653e+Jk15/ZQgUwmGQdKJ8u9/bmMahW1fmj4y67+50z1j5CAKQmkiM68NShB9G/
6IeJBLjwq31IoidhfmtxpwvZE6IuruEgKTmSqY15LTPV72o/PuG7VRfP82/5bXRQ
IQne1QTi6Qzf9oiXNU+xAT1UD/UO191Wo4BkVz1jDBvyTXRLQBfqMaUtF5m1USYx
1jnSKFzuSN5VwPKx1qN62TSlQAxKCpYVpGr5rk+J5wxYdjne5aq4bhumoCIGpnc8
J283VOysB7zw8LxUJ3mf0G84xUATDMBc3Flvd8tb1jX9Yc6Fv5qQ+nN7B9usouhA
lLw89AGIY7Y9W7mQ0HMxQu9hkaYZLV8Pv6I1RqNROWhuHSQ3jC1ktKQWIXmliFob
RlSpynf4lHajyCXdr8rgDaaXoPEhL44LS2WAvNypX2lVkfb2WIetORgceRp7l+h5
9ah2wEjYQAiKbIjplMNUjWj6N5jNzIbQmtpWHQeS6Wxl+M8Id8jLWrlW+pUYO6XU
79tq29qCvo0NH3jxZw8CAplxFicPl7EHBubYqYRn4M4h32wc6EhFyXGZaVFgvsWl
Bjps3h1XoszjIgxF3ONNgFKBO0rPsNzoMboB2R510MdwrnjE+wYqtBoYu9vFF4p+
3A+3zu5K9RpKnxLbTHiZ0L4ANcyujYybs4fnPkOkIKWzKuISNeybLH5kqxViWbqA
PHmuzDg0+WBSOqkQ3kZHAdg8KA4ooo1iwql7MBeDoNILjiNnof1mDXRP2AZJ/dH4
4x4n2L7oCrbv8UK6GZnXkSMcrWtkMETFULlNop5YmfZMGDe5qgJQBosSSs0HJmtR
L5/CFI76YaWMqkYYJQVQ+Lr8tZmCNVbC6JREibp8LL+2xtNg1WWqz2VGSHJ6HRFL
Q4jSG2Uc8YLaZKJo4l6UlVE6GxzicZRf/AA/wCvBZjjSYjTdmDfXs7RkfUxwCmxG
QqnK+b2AZpRzBogdxI6LmKyRlCM+WXyYtChUOvnVnVAdtisyTBfTH6dRWa0oYlBE
Nvext29EJh4hjIG+O6ijysOnCzx19QRkZ5o8jpolI+oCRgrOVDkN4+PmWm+/ignu
1PrcB98ycayr9ZrTQ3QZeHtx7qqR6RxSU+c6BDWIdpaS+d/+z2vmHGyVPonAg9AK
2lCBQh3boBvFPt+uFCyqTJlE6ZMW+OYl5gK0nFKxVRaLozaapAy78CG/qkH0Odro
NHNnEv+pam7cL8n7Yw9sCOQKfe6rtAYVMs6f4up/qYziDKR9EGcfuQWtAviwCYib
IqmpiuEx/FYzQFQNJ7tymp9e6RENUloPj23xzlQ6CE7F7x+NKGc4SkZ7HC5JobbE
Rg6QzQAZvS2X4o9UFOKWw50ShmlLInt2d/9a4hBui2gE50dApXTv65DWduvKj5Z0
VsvUvmnjhiW99cr7NR/UpxgWz6CFZ0usSSeXdt3/Kfi1RrsNf3vaVFV1IPEvmZOg
cYySyBHYmHaLCTj7tFbOK43qD7pImLUG014yoFSfWjgFfW7H0jzmnNhcCWgg86dz
EQARKXr9fM5WHUJ9JePKfhY0TtXU0+0BqtgiYp+Nxr4QMwjtO++NattkXrfX4TuT
Wt2IlOTGplsoH7ISkBJAsuvQGomdU6M4iEenKhnEpi91oGg92EQm0f5ys77g61m1
BxKdXQkBksH3gD/1Ojl6Lrn6F3x0RApoLcb2qleEMyM2HK0lxavET57UkXBiIS6p
VbE7CxhJ8yqJsLlxRubFpS9+crzD6VP0jfYF0g+v7ZiemuyVb5vc5J2hKmOqtBUA
tR+Oi1qP3KIYFte8YRrBNz+kMQLLrq75xBTRIWYGa4YzVBlbR/gGZgEaa9m8ljxW
sxLKecVvCCbN7Zp1TN85VbxT12vbc0mNE0mp0nf1zPGjOH0U1GWRJ7PgBr974kvk
qCoRDtyyrmnViF8zTB8AVxGxK2/izJS75nXPawxuGURWBgfBUwcq9G1/cAiX/FlO
DPEkQyhtK/fmG55/BqCMprNeljIbawRdkigx+4I6/f6/wIP5bj+cAVKf7eV3PTcA
XmnaZrjSQ+CwLxuiR+fBDmGi+RqjbCPeeNbzYplY7URaBDc8qJkVy9eQ5UjLTbBt
VYUyO+tVTcDKtSsK9ggiImXniV48ZkVDN0eBCvZpb43cEiFQmH8i/sW/XAQoFHa+
iHo+9Ar8U4sVi2/dvu5byB5obkKePv4zPruW7pMi8H2lQ4zYaSDkpDvLSaLJan3s
6QTw12NwllEf/fRU5qAjm2tbf99E7zjpN5wn65pL5zNrIwYA00rkrXeRHtAlIqhI
lKMCnqN7BQXialSRdGqkpJol8VcQX3OIimIE1ejhj3Pc+dwqFbo5VPy2Z4028fuF
zPDJ/Kjbu9bgUxEA3yjwThIJu8rLo+t6NOXcwMD4Y7UUvsDOh+4Q5MfZjpH+KWvw
3Os6PWFNv1BVsA3WdCNtmC1QBRM217fOcexBon+9kOT+AbbZXYfBEI+Ky7Oca2Rs
wvzOFyWzB7eiczOb0NJmIK+dfbqExKLa86IXXc5nH7D39dGLqwLPzuooCxhiZmHg
Bp48T4ZXLR5IoDDX0n7riFI/37aBM9OdXlfwuigxe5n7U4Fy9Nn6so4ONifpqusF
9gVIi38If0fBZTeOGLTRAVvBjczRghlDu+R2+YVfZCA0WEDfLmP8c35cZ8hQ3wI1
gQDL6fYqF/ivYqW//lE/vIs2rWAvHgF+yAIcA/WFnTY3rxmRXRJVb5+1XellNJMl
byrTN6E+1XLbIomrV4B//3YIoYVQNshKIz9rGmEloiHXySfyF9CeboYfBlGzvpwa
8LCe6JtoZjPgIVr30kjvJ/7VfEBu+yjTAfjT6MRgIHqjyxj4Q3VUBlDi0KR26SE2
rXRf5u5kWYRFi2iDfdvg56cDIYt0pU0BvMYg1dwecLQbZDYqT1Sdfz2QO0CwiRiO
YxC8rGNDcDq1LBLOKEfVelqFRYOS7lyfi1dkcEIDU6+YuyXLOeLMvpN49Hf9l0Pm
le2GyDxyUvnxSvCgnhGS6H8qllLInofo8eqAkwSo2EPjsWADJdkEE9VqCNfeIcYG
3KK2MNDDn12V4/h3waVBmrxNPmeC+NuzVX8GMC08PtkaM2zKccKO36eQbX4NGBqy
oSww3cGWtKVc2dmI+sG3w0Kf0raLoW+d7U+qZXOatk6UtZeBpv+POABl0SnoD9iF
saf2tEulk98zsK9KwPO89RlkYiTCWmjDLgJyvER5+hDOPuCOifz3HfCX2DF+YaxI
HchMC4kazAgIH2/iRFZQVruIoRxIgSCRDwKV73tlzGP4WpAP7nXqIpvi1RQqSgle
hnM92bzdpLi513agEmGqm+KclNfwk0aGqsNdiW1xekDMvzeuLJcs8FYOokmOJWP1
aR0DdMa7JPWLFfjshE1I/h1cCQO9o5QJj+GVkTa7h/WIW/Cp3w+jDmQDuRS5IeNs
yTB5SE52sM0mt5wxaQmFbIWVlVP80QFOhUj281bQ+reHqKZBti007uCWnKLQocLR
4H1APyC9MML9AqWgcyTDYj45Fgv94GkXtYLqHG6QL67FdrXmWnYSxyMsx4ZRB/9y
s7zUW/64c7IBKawNt8x3PlfOTnsJyPOMP8bglsVQBaymlUDHjJVKsr0I/H1q1241
o40aVHuVmqykLhRfHL855YPWSlx7Gkg8c++K01eel68ie/D+1n+aL0r/flzYpp/R
S+QszSUXxv+FTwJPFg9YK+69I/gI1Mb3uUWhuRv3ewX+dNr+S3Di40Km8Cb+Ixjl
kr4ugJkE8yO2U4sjdiewuRvaYbOx3R032EFEZKpOv+FTeA8dNhaLRQLm1cYkpJDt
PGd/O88TW1QE/iZ1QyFGZUjFF5kk1U2OgnMjzvvyDgR7WT6puSVyRtq/vQYZJcfv
ThGfDLbcnrz18pp9OZDBzGzbW2uQNVoyS11kaUq9jGB3mIvhHUVr5YTHQs1OET6f
DWhYB8uGwvO6XoFOQxnG244cFazun63Ci0kOzViTToLRHSymmuLck3gv02S91azX
rPbseImjGkcBuU6Je7DTIsEC3kFhHyf8baH9HVejcfwQ5tqMT7DaIOR8AVez0ZZB
cFEiwuv5hfPocrvrOPq+eP9rdkKZKPBOapuT4Iz3/mz9s0cxSeMzYYllkbJGVvO5
DSFqmOaesgSn+AFRq3+VKlMwvoi0r/Q//qwnFeMIdETLIczxV4jJUeEcG6R4057r
N7V8FPztOo5A9CSyvrP2+xakR00vGQR8zboabn/vvoZf7/cGUvTNnUiGYFjFeLlQ
ZX9ruIrMpFlCG5ow5NURGy12sGD2KIT76KLudyQe2fqNnieW3b7hZ6z2bQ7jiE0y
iuIrQwyE0xAPGi0Sghu5MHmagEhZySybiDfW+GAjvtc2cj/dczdVb63YrGeXD207
zMu3/uyDBrO5rCfdCGJosv8Rnxl+k8t7nRtITaGAVXHfVal7r7mfGh4aWjEN7n+z
FHS8kcywM5zio+KWuH5deQiMEehh2yWUIIRZFpygtmd3ZolzecDRreoOefNPknbo
H9J1s1ncocAhKwnIHj10G40OFb3sVwFfYzTsSzhXlEBef4unnIvukk7pPxHPAYEE
jRYBykpRa1fF8sGuze9LH1ccNXHHz5b2SiTqf5S0ahEzztpHzkp5lBDobNDHJr9T
9Qt8GStORepPaOfF6zobGvMgPuk6xSAiKEoHC/wk1i/nFRNzpxgMpL2GfBxZmv7t
Ia5ZZ4oZU+Kfq5kxtsjahBEf1aiHRdCxQUxdaRKkpMNg7McrF0Lh39vnWrsYgWyR
vWcvMs2AJwJbciu00u3Wx8GUji8WnFvaM3sqHw0SVkexE7GFB3itu69naIcB3jlh
2y1FJIke6Mzbz3Tz9OSEg1cLscasd5lWgfoixFly4NfGNHK5UD7oaUCFjegQrlNu
VrQ1qW8dxFX8KbOmHp/nijP8QF4JMRXu9SjDE+C1hY9BAE/IyWjzQB1Ex9f8KwnZ
0luM7f2i1QV48HolunmeZfYREeihJJYtD00RWpkU5NLliSiRAMwmsei/dvUXuHeP
K9guCriwlK3ugX4vKgyPk2q35+SF/EBjBDKLluyygf5y3u8/2XZUEzrfKPkP9xJE
A6/wT4Q7FNP5/mK7UaSgQ5Oh37m4E1NL3priEQBFw1+LsoM5M506mXaYuRelqyA6
X+G7QEanKQfj1FERtKZAtR2uppbSKV+wubTbcy7gEkTAWg82SAQDpG7fhpn+acZu
/uH2ZZ93AjElR02PtO7OeGLOZjVbVujw9XkbRVQYFZQujdS48r/IzxepFxM7oNG1
HV0vVFUvLbDYHgcsexri3cxa1kWmzGBPXXZDTR7oQFch07VW/dtkNlrx7ECaGsK/
WRN7pWwUjWzFnRDQbSytWoFW5w+UknOw2W7nVxPTbVCkzftoys61W0WIPcpfgL5Z
d+eImHaBDW4tF85BrQEzZKqoJ911WtFVgIretb7lRCILIf6KNWzPUv++boj3w670
+ndPDEv3PVAeM+IMROyDMM33jhNyfHPR+Y2TALZ52jmQnhV6r2AiRDNdyJV6S5SG
AdCzkdHyyX9kXun8ThgsjAJflboDjRtj4XShxauXRTxwcHc4IFcgc7Q+9F2DOQRs
jNnge/4XA2nIXo8vB7HoMWQY4LWEEpJtQu7pFIF7lF8YzyTtGQsrQNwvTxrgKkDM
dxxeYGi5tkQFXEJIIt3UZI0t0Q9PIjh72KFJ6/X9aGayBYr7MNi7BO8ZW/dSpLzw
OBJUJ4GJGKwUlsRoYObxj1BU4vZzaG20cVyppv9XZFpy+L13vJ5VT5Rgh6y4BVqp
9qS8/UNjOsUAVkKodIOTOKUEE0mNiF/Y857VM8Rv5eWWr+LXCdb+0HOeN8cDlcNY
4bhdTtcyB4jpU4FqNRM8kYp0q9v+XnYTmk1SZp2tAjSADeunz/oYKbgSDDDB0ijm
vyhmhjewogu3QeTUCiANB+ijTufP+EsNTkjip8oFyzAi/GTilk6HOL+DVP50nq0A
FmZQZbbhaJQ2xqZp5xYAc5X9KNb6FSLW61IQ5brgWJvomZNez6vr/ooKSQVZBKn7
VZ9QM7PO0mEcQ01ZSOKrtVbRj4QhODvufMGxzirD0b4v+HoCETo94kU5LXv07pHO
WOfnqVHKbIRLyBS8FHQRSem3I+BLCsWUT8ngEFozaIEICEmewf+r5FudcHtsGEKX
cj5q6+c0PSaF2z65x42wPsTWp3IMcvg+GegYEu8tsNiPeYG9f312B7JQTUqYSohZ
eQfunXF6Y7uFb09DNDLhKgIvlN4Xeb2oXAPCkQGPsGtozxdD72koKwv77dl2uOsq
7Vo/0RXSS1UPzyjF6DRoqbQKtY8YRFmy4b1x7xwmWCBRmsDqMxeLQ8rdciDKiG8N
GU7gmX7zUVCIT3wYbPkshd9P+knMLvk7xE6HYY+FH0JDxFXXve0TGoW4cOZADKi1
IvscR0WPOyPvDSXm/XxPqCAAZw2eduEYEsA4n2h5lJazVdW+mOrsAKzygH1CSiEG
PkvsWelTRJeYZ9dmDYThaCh1/fcP0zn+P3slvwyHCxIxud9Lu4ckw1bDA2IcVJqc
v4hjou6RvtGKZdqe2hPrt0dwXhG70Yls9JKvi56q6MF5rTpfYtd6TgBrr5UtRhoj
TUc7SUG1EUJqekbOGlfFuk9uf73OX0bX/UAbbtJ1RaLOjqhvO1Aik+VmdaVg+A3S
lEeT8Ft1QY1fOA775jazrAbrXdOygkNsEAo3wUo8UQuk4GqbU8kgVN44cQGDnZ8Z
GgsUT4kEtdOJ+S52SOJcO/PrmC5JwiIL0nYN6L2dTWj2opCiD06ZDW24MK4JodQt
50YNc19syPiPACaUkIQhcsCg1v96TgCS79rGMsO3owPgLBn2G93mnjcWZxWFp/Nw
ayAFunOdwYox9XOm+FReqnJfj2JdeVpYVkmaIZDaxiYdb7Y4IQlcTx/CKy/+1ZzT
kKMIxjto+mLFrMhryhPR1Lt1iFBkUIKXPpeI+sppg0Eqm2fIACcpF3XbqNtBKFys
PXQR2LwzfiP7+83VFvSt3zrsD3peO8ukWYD49HkhwYCSX3D1YiXT/Sa3Du0LwuB9
u5A37FhX6gOn8yNRn7nfQWfA1ulWbXtZQQ4w5EkGU7iCdpve8a/sw75XDtK/VBBX
dMpxvXsvda0yQ5y57A9exyloVLmALU/uaPre/jFWRyRvlquOYmQ5LcOmhD0GeQnW
qrKa654jgXAtp95epfCCcSkJz42v8xmUMOoF4rXCvEjz6T82/4O88q2ofJopF/kq
woIaeyZoPfLPHd459L4C8WpuvKvAqkAgFIMaItGGKaBSzOt61Yz2Rdpo2otyCQU4
0m4D7XDlAdiB5gXCfKGEdWJL9l2ANT/YAhSPoXF1BWceIoIrUbMXUQ2ftfCDT9bB
womB31oOKLSqfgljyvvNHXmDgDbvsG/5RaP17vR39CRqFPaipcXGm0J1iGZbWeqo
SRYcgQsaFAR15+nNI57AhGOz4MzFH/vMSXgC+Txr8OOPjaQG1NAV04U2xCMc1Krg
UER3len6TQBtQtLT8odmW2BYYomWMewvhRAVoNyFYl8Y2ldDJWk0CzHsXpTf173+
URhjphaobQ3uCaFBEH/Y5DVyDLmnzDnH3mjcmfokc+fHDkmPeYD3a6EP+Z1MsGg3
loRtYosJzZ1zKJ/PFNjzTdL2BaEYWahMjTprzYgWOJDBHQ5SS/7Knf5jEJxXfBBd
JFvURRlkNueJTgMDXtfR+2I1fAvCER9PbUxlxEqeuUMsdZhPqK/ReEYB0Yko/L1y
5naGQMgEiNAqKX4OKpkTEBCITOPzqW1o2N6LVSGneHYUIg54kufO9OZGfsaNuHGs
J1gi9gCTMoxXWOMNr6uCjdD8fchqS8VDN+xB3Nh5AnrKdgK6I9ip+y0LM1zekHGh
vOC9ZVGfAtxQgp43Z+wLKFhsVWgR3hn9J6dpoItqPBCk9yelKVkqdAiLKanFo1JY
lITEDKHSpNeX1d3ev+mMiU0rNfwezaipIxapXk2YVs5k3cn8x1lVqCRIUXek+QcW
pMnfmOrrbKZTA87y9WWIPxl++oqbDwP43fM1vUhUzVgvv9F3MYbH4BNCJBonvRRD
HlbbHfzqtqpYkniSaxZuJ2Ml6dPWi2kgtgdV+PTGT2SXGzIf8OIhD+O1CqDJ/UDn
z6Swr7h4FI9tDRK3S67zWhOfOytRQ2O2xZ7RIJKR0srmfgwLawH2pkp0Gsj8cL3N
r1a8XiUWWKexCEcLloJGNi2oms/QumWkEgIMrHwb3ccNdMVtW0U4Ds3QXymSr1uw
bo9GAWt/sLm6TjYWEDTvXlyxAhAODvp0LZXulmtJhiauxZs8NAFZ57OiPy50rgpu
JRR/CxrA5bNvaHdwcczt1oi6Qep9LR2DdKokdqgnN9d+TGfrtAKvk9AiapsMubYW
Q9y8RDCmK7tRk7QILvHGlEOJO+wIyyomdUDwNLomN0Lbllpec766dsR/Rk0EiC5O
tJGAav8eOKw2acplPgi51I5pMf8qQNk7QSVCesL5mVQBMiUFDPx0s4j1BfeByLev
LNuQyeYH3z14PlmguftiiBITnpWsVNyDLJ9AynCSUIYwnGxt8xaJvkk4C1JVHBIM
CnKzQnLssvEXbJT2jcX007MhrgrR2ppypRuJAJN1/6ldlHxc0JhjvwWp34iBpgZq
9/zBCH1+a61av3jLbj+2sRHyqfwAB76O/8O5Lu1FDzgXIWISJMpPm3hPl9W27OHM
hIPJmOxuQ/hxiYAEqzuYxjRTLvSDzcAlG4BTz/YUIaxvNRxDCAKg+J4XwIJXwrlb
seLosHvTLW2OcGNIFmGTRhuvy/cbRc53o/hREr0N5KKEOYrEdlY0+5e3uEmsTVkY
B3RoYNCI9ptr75DT1+KAfA+bkUPfBVB7eg3FHgVJlaI/wnampl9MKAZ6jJGOi7Uz
63s2CZlOPgBCMNoX2qhM9WK6akPbzuXEw0+L8uXHeyVUhflS11uCDw8zZvOjyjZn
FcEGD1q8OEXb48zXhHiF07cjNqQ9UOyDwvNNe06DrD3A4A3Aw/gnRCK3bZso5yGC
q67hgBCFoOoEcU9sEsuxm0k64r38d3PIxT8u9hwzkfgoHAyJdpRNm5EyMZvWve5J
du/oTI8WmRckgh4zC9KIYkFVtdfqzzVV5deyt32k9bUvO49clujLLkLh3UZlqalU
GU0OuQ+YVOUS38Uy7kLNJ8mo75UU6l16JIM9f9MIypIiJH6sWtZxftHAzpg0ZFYb
TDFTyrH3F0ecnocj6aYo/Vc6L46ulPBjyY7s9b0oRnsIyK7sgbeu32z7nUmrisC/
ndDGsbxoXvZ8+v5fpnz62BKgD1txnJVJVsXQzaiAPe/zBYJ+qVieDbtNhBuX7hs9
U0uel0Ws9gbmL/6R6uJjkASDsPg0gxNOC2DnqCLGj+lEsCVzu1Qk893Cr7uPym7/
96yHMwaHQncFK643IpfRPm4WIF522uHXRoj6hbc7kSZ7RPgYJDE2ye6KKqAu3DvJ
s074YblxT9kpsazw5KJIYl3kzyPX31Ulvvg+VS6KT+h+B+VxlqMALxo3kTvxahGT
mprZP7z0jCpXvvdeyp4Bs+EWbqHSLSqqKEoCddGU/kmh1ASubySoXdrDcOp0y2Xz
3nmf9Or8lSMQUieuE1Ib2aAnGE/FxQADfdDQdV0r3q3jkkbSuG6JWVeGew1mXFXM
7t9/2whyxcSP5L1ipQtqFtVrQI1SGPoqiazSPiaTFITBidE1ApY0il8lITXGp84S
51jD7V4IplEEO9B1ra0hnYogiqW/T5zL7nwSnVKsMrNe8pR3FkQi0JJZHnETbxyI
pIjdYN/GfTalG94runiv3wE9CNk4onzMfUaYkzwETTXj7IMf8iBJMYUH/uCfujBd
PGSb7QBAz8DiI4wcxkvODhcJSn/IdWo0peX5w43Qx5BlV/6IKVJ00N++nsl7wP6w
fpCz+AqBgk0+FylC6Yt0RcKQdFCTam7aJ0tZr2Rt+Em+D2U9MtroT6vgNE1geNyh
v8gKh6yMi3ONptIbsx66rst9xG9XYIyIvNX4JVhKwGuUkUF41lQsSTKtyITfV3by
quZpxWkYCi3Vxvqf3Sj0Yjlq5mnQI+JN0TwG4JmoJoTBcM2yvTCCpAz50XaOYm88
72wf8QeWKV1YOB/57I2OjHD0zYwafbqCKeeyV8hOspUeZQAtwgy2c/PzLR1tibum
zhqNxaP+TsNBjw8Yn6NA19CqdX4GhqEr9elihAVMcbDOZz1D0JnWEXcK8720+xuh
QfefR7bePVEG+oGBJJ1VFVWsiVatqLlO8wKHTVUlFNpQOabeiM5nPkEBQ0rXiN1h
LHEbMMWN1PF/UwXrKGvWh51eeHGZgQ9GFr04Qt0no0cfs68LMs9t5kZTn2yRv0S6
UNwWhQbnRBrLBdHF8IU1a9wp/6K35SQMyscqqAZZQNbeh8aEzQjCuKtOzgNK4txZ
Ogpb6g1zsepSo4xkiuYDbF4Yc9wVLCGbtWkMEBV0b8nYfBiZJFP/gnHjAwYESuVI
mw1ALgq6cALVaPkrzQAQ8nE9OEXacj4GfMDdJ/sFkH80yjUh5UB3DTxjD5eummfZ
5nBUUgqOMMzTI+0gIaeLXg5bE94D+33pyW34K7SZRev7/50YHTF8IwLGNAeWmYXq
xE71ueUF96ZXpXlxx10ZlrPBPGTsGuto5zphPK6668xWqGBWmmLSDffHuoAsSB4S
TXRvYLa2ITaopCs0vsPCGlkDDe5Bzi9MvIrktAq6dAyptBcVsvO7BNUjxl/LBfvs
mwRyp0gM6/KGFD7y0o4qAj4AUROZVeyOBQFxU/OcRDMH3Iros1b7m5tCw3GG8B0o
Td3OOqTGBSl6csXRu5BVjgtmPBY6jJzTzsebdSh5OGt/cxMY5rHdtTf9q5Mkqckb
ev3GokclKu6oUeciFse70yvV6FOl+8Rh7y79UGuSGq0Ts0ilxamxyTjBI7poKV10
Pf4jvJ3Dlh8+WAvxGIV12L4Ywxt9olxkZ82GRgVpCTVblsb8RKwFmSOU7Dad+53K
Lt+h4xCoHg8AKxlp/0F8PyryESEdf17a4is30rfAGMuxCZI1d3ZS714qOlILEZ98
cagHkhjyT0okqfNDWxCQ1tjKZ6GM+uMabO9C25jvFiwk7ilYY5P9YAh++5MJVAS2
nfSWQhhaBHe+eMVYCDpQGisfEg80AyqsjKR42EoBqPbNl08VzYNxuaGg2OZ0ClCm
dvrDo5YweaoPN99dfIqIRi4HKlAoq0xiVg+q/1NAK0+MKaSkHv7CxqRHMWa9t2DA
KJI0LZ/StNYtKgZXwWiX4NWiTTYdSAL221NXWIdCjKCWrTQxrvLvvrRnOTAv22Bh
p5WMqL0rjWXhE7IdNBOebxnazdeNqDKe62GqrQdasqT91ZhkgeUNBkhF+CAuqreD
L7S1B7Yy3R5O1sbcjrxLkABjwEfw7Ou+sYnDAdedf/nuq8InSgy05hJqG2p30PXc
1BZHwl+KDwhX/SEzvI55cd5hp2PeWSYVKqr26wmaeavlkLhZ/y+6LjRgOP+gh7Af
semGMdk4Vn7Doy8BY7grFbcyEcYd6Sqc4Ho25A/yc6sWVb2F/RxMU6s17Q5gE+rZ
l9nZButMJUEGTCH5U+gbjR7/mqdWtcTeb0O9jLCcD5VVVGDVJ3/8EmQkIT/QVSFL
9we6OxVzQ1VWftCLFqIpxd9mWDCd4Q+JSY3Kfb5vIegIpOo2GrNO/edsphZd6efz
UisR5I2qSqOyv3oE7WfDa/D73FMauOX7KW517waWZOVBXio0CS7V84fugfYyJDjK
P3LdJ/eWzrF/5XoYpHDawLV980EF/5epgKJc5gKlcqtVgKJqbX3GLeZUCumUPMFl
/R9g8hmk5HlW7C1RZRvSMcKq0Tg6wwqpGryqZ+vuqvY4FurnXOp60KCvbjiH9RLg
cCO2I6EzjzFQ4F1wD4nA656OiRnND1dNGXfDeyq1oaimrVFoX+Ge7M/v6muG6H4c
SS0I7N2/tCJ1CRCEdBIST01mUWuuaRmsANe1XhhUa1jc2HQhoBef+h3EKF3mZkCX
57p7OC1aix9VNMrGgNqaHs7CWhPe8YQxdiTbioLEJFAL23EmNP3BO7i7CE3JAo1S
W4CZdZzr+7IwtAtnD80vlewVXLbPsKWWjagHADNQwJpQD27JenZ+1pKOEpYE+lmz
XvxMw+3AVyhosXvu/jdzZ2hY3UhoWGRwf0XYJ9W1Yn+JRW4jaaqdLTXYCPDvg78b
0I6A1chSTtrSWt7PjTFyEno7jjyqMkt1+sWPbO6YOcZ5mk46XkyUA96vNLwTBQxH
URigASDTmY4111P1xpuff7wJwAIGww1xnRhQ72RqxX+5hAex4spmxEFAVZ/wj35n
2zGPiVVvNEE+n/OukjaDPZJPqrp/iPybVYZvrgDLlYEcLEYa02/v555bIteZ9MYm
PesyQyVhuGtf5V6sa75Wp539GN9XI7H3qFYVBr4I3zfDJgScHI1cbBOGLbXqBORq
cd8OvH7SeC3/BZqJpijwj13uEDsgJZFCwYirRMgwlXS+YTc+APtzTzlI5787zpNU
WdvBH4W3CUcO1cCAX4H99ToOlLGeayssw4Yt7chKW2R06oWGFgMhKNmFA5KyWnFw
AccUCygXmT1ZA2TO2YKJwlNdJor8UPdIqBkfWOU71uhu1tIiuQbRclJUfpR7B+3P
yu1uhCCHBTpQtpw57hCXWeari57BAo9maisQWm37L9gcoyb0pCY2hmkI6RL0DpiK
cYyeI3nmx3pON/3fvYT6mjNFlgGQqYeWjFWmbJNVWj2n2EKBcsFBLoh5sumWA+sA
O+Iy4KYBzjmkxJ8wNqBMqc+fIOFYdbR0/HgbvN56bhNFjrDWMbcZS6asoXJb9wNu
LJ2+VfsRyS5KX+0Tbw3Ef4pkKkSZ3gVWfUNo9GA73KOFPhwSoU+jaUpu+B6NSAF1
pBo8HzdaacZqmcPE8kkwLkjxVrZ7mhG42oFE/x/Rs5CTGImSsZRmIRVol7Gv75yi
r2AgL6aI8sinkpZ8ZtZYQ3BEWojUkZroIbwJZLvTuiM1VY8qXu0XeKJuw9BB9BBW
nOHbllCXs5SNgqroAvPMQfeGdGcZlJ28ML034jCAAK4pYSDLMvKlRq0xwpBWquLm
ykRpzziWSRbXWRAjgHlriLJ1a+wbQl02RadlibkGSrHCTx7IWfDQRQ/YpucI6EuG
sx9+satVNpc3cwNRjiRpPwvlKqYgFRG0avZjqEu7Xg4CtkLCtlwyzHbOE9NkoI/R
uzJZ71VtstmcYUDPtK0lwdoDdvC/TIIBnh146I9pomOJ8nFJlwIIBzbkxKpuKv9s
IxEgqFcw/6GH7ExXFalOPyqkGBiEXDw5+9TW/H8b50u9LOgxwtuInYBjT4Ki06/6
JhVTN9lR3AEYNlFq2mZBvyZ/+1U7iJvQzBzPuKWdZuH28FMnDEfxbCRG+csE1qKT
KBhFpR2iV5VFPIaFsc4J3AbhAfCHg+xm+i7N2w+ja/rsFZocoRW2RrbYfGstFT4u
RBx85saO4K1hAi8PtUIpQMUrdQ1Qm8YVkHx7aoybAdKX/d/dUE9rMaWwMR+ZNCn3
1HcYeqk5UXTBUzrkW7M0LDiz+VWq7ZutgB2kP5VN64CefDA0D9i6pLo2aH04eqcj
Wdz2PU74Z5C3caQ52PPOD6HLm42jWVt1Ln0r7MNp8Szst1246qEgJ1SQLsA6siIe
AOHNhY/bW4c3eZ073IzdXsqoZV7Jr/M8IZ111AYi6AD7dBdxsXsDWFcyIdetJ7u6
JRZd2PgdJw34u0eOolT1JO3x5dGhbFHSw9shhLbgob6jb1mYGiUXNHhbfRBaZiO+
xqk9UK4zqiyJI314pTvMWSVDcP9TV1mzu9GghIESGazDldKx4AU3GfFU45HtT5A5
+jtd1r3QzhlJI8yayDEvTfce2exVkKd6tdB85FbbwI27hMcDIwmjs4lBEebdYR2c
Tj65soZIthw1LiG30C/wqm5dwuYREWSQ5duJn54uGKJrgZvziw0zM5K9tX1Kf4ln
+eENuA1FcGe+BLtrQJrgB9HD8Ge0b41ziddeZ0z27R+CG3+VhwkfDnDsoZBuXo6t
vOaLC/4HpHQmOKrjZCl4OTkah54YwrZwNiP9TBnEDfmU7ncuzmJL0AACxrB6j4YH
oSgCQHGnMTOWmkGkdbtdFUBGKRec93uUBy5intPVoOevu4ZVEGrKUoQ2v3LdNRUS
+0Sqol3qFybPQ3nlu/vQC8m10/J1Gkux+fh4zmCZbdanVgqTKmT26fe6nh7PeW8I
HuMXgkPxgwYAHx6ces9sBNhMvJPmw+mYdcrPu8U0gaIi3QmiBcnw0yuiS9/vznCP
h+pDrkUr6DLWbUk0deJNtIaB2jHId7GaEkAPIJogCBKCvyN6nQv1NxREGF7a8idy
8KGKlr2wiocdR/OuBTRnOLrcsV1CINRm7cMRJff8gOgsiX42usc4FK/aTbrNoNAH
uK6KdzfTU6ELYMt3rMOtwiGsWNPGeVwp0sJUvwLtwZNfPPr5a335Hai8ZXDDbATZ
LYTrfzULFVKNPbdieB7xa109wMkRyLlJfIpC2rR6Y/gGh+bPbe47TYiY/Hf2E6T0
a5FEwBafKVli64ZUU4EctypMTklIAet4KKzbYZjMBr7Na9luggcD1mZ6lDD6LThy
9hIrrssZQ3uxvR/eRiLzT5p4FPlS7IKNVezZjeikLcbhhdj35hdZJUMXyDEW7I0F
AIfIxWuLKOzsyuvaJ+YrcT4n9jUcG8w+uMjQCbepv+EAN6QGTir0DcPpRr/SQOYo
XfN3QHjrsMIrTlFwUrk9tz+pv2tRFzXjdo8B0Mv++I/i6Jb4PsG/BoMXevtma0Xe
ift/dpwTsNYl7T/CFwLPJYGShDSoFe4piECttYnU5uzi0zFxp7sm4VAjg+Ds02Nw
6odfD2pFp9XDlTJf0l+hodzjFUnCnC5S3UlLp/ioNXDdIB7g9gfdUr6bwZ06N9Vv
+tn/g+FsgVMR5OVjBTjauOl1/4mrG7w4ddsZh7rejfTBcKT8Qmf2Qj6GslkK67hx
ESx8nBZp4W9oIXCvyhXYWL1GABwfboRdN7k+x8ArXVreCDxduFRA3L5DVWKJXE5K
5HZF7sFejoOAiuVUJwa9F6wSbzDvsyOx66sbljfMx6iAibsIstEtxVi3IAACE8He
N9uoe+7KNVBBwQKacl1OMry/7PBJkyyF5KgFN/2p4eoeT+hxZ3/ZtQVd76oQFqD7
EbgRgpnr0ZOVW3gggeAP1vTk210taVD8PfkMz543N+t62w+l648dp5SejT3R9LpE
HVc9tbw4wTDBZQQr2/dfumSaI4dNHca/y978LiqA1prFoqEvaCPUL5pmqlr+mv2W
J3b2BaZRV6i2u9hXj2qpPkFxGbysenTAxk1sgKgjPkiL7i0Pgc0lW9WKGbmYrvBN
OODgo/trx4kU9iGeHjXAiTlUDKW2gAN6ztluqFgDivgSuDsF8U2Qaor1ENl9Qu/X
s7ZZH6iAWFBKczI0Ub2rwamBATaCi5BFq7gA76LMJp5T7xC88PYrN5x7j0u+EEOP
hOAUjCt/yCMOmFI1NQf8BgF1Q6HaXVBs3oqPsBp5ceN6SL12IGxsvt6XzA5NUyd8
bS9I8LzZTAs7IinnWMZoG6O/A7ZIL4loj/SSY6qZTUkCWTjk/gvy+4rQgKUdWdqX
ifxpcq6IANVqqdxSb3007OMszr4N8hDzr/oa0RikYsED0TbiLixrmsceSz2LGzcs
g6gYSiOeyKSNg2r3P9USckHZKOHP3qiafM2o/fS4hZUhiVg7f/nLR+u6mFYJ6vqG
NZoLaIZKc+ASAJ39bbpI8lR3jeLBMY6KVdnkmeJpYZZnRu0kSHlxV+CiZ97sjmOx
Qqi+f8iSk0nOU/5IpNLw02WyOZlApwvswdX/4v3ygkftRRIOL104ar3gDpwIEQnw
p7sP1jWkR0zZniCor57v170utwAumWl/r+rIghLkP0khZplnZvVsq2VLhHcJnWux
SKlpOa7w64pTf1mBLHtSukvPE8uNIzyOG0mD84bKyYJ/kcykoE5eDGeAbBAxR25p
f5CEmC19PsgxL6RlNCXwkAWeawFqQVat9ezc7IZ6vEgg3VPmGrLksTKjNw+8u4Ar
lk0K7yB7aVopOjs0MC8YAaM5T0f/YIJr6CNSZpgfuf5JPfNCb7/pxx8Xa32QY2+b
pc7e5Vk3yI/CH9hPbRvVuvQoI9Gvio5fvjJxyNhstlkTXJYJtEavr3S0YDpUZAi4
1kojdaoWFhKRbggSLF/Waf2prysII4bFTEzHNjY+CvEBe0hXtoGHmC0kD0V1uiUV
s+Aqlno81rFyBmHDpIY6/mIC7/VDC7X5BNvxUfirDolMyGe6nmnJHsMeDyZS79O6
4p6UPF02SOucx64T24yqzyVAtb3ByK945PQax/22PyKrURvnA4G4t1C5DaAYi4jp
rWsQI9bs5HKFlVQcIFRARJXq2BHbFITwk8kVSVTb/+HRNGjdhYLpR7fbdA/TYMK3
89pms08u8a1ZFPIsfWdKgsCTGLk+KoCuBoJ8t7ZsUkg8pDEkGuEuj6+W8WV9LRIy
U0SqTm0o0faDJxy1VxI5insBMqnSRvf6JyqrokavvW6RXltfSo9GyBx4e7mX0EAk
oij4OZkIkKZYaUcVYozCuzBcIJA+doGRfeC3tvEqAaT31hwTd37aIEWwOsHE6hUM
XhDpHsjUP6QpFnQJQCVnJPNUt0iMOQJhHltcwWC58OeLlkjbssMVv1tgJLqGUC36
bFw0gdU2v7Z0r60afsotWM8MrZpGhA7bO1uksf/N9n1zQMsiKQxGt1UbNwcGuDbO
DLZFOqAoLhJd+MIqRk0E+MisgYJ8SqlXzmaEFQwIDX+3DWoCcP7upEoHvu7mm/RL
q8XOZogwE/m6b5HW3LQzLUw+74HdpWTEoQyq/ayHZW8u+biiPE+iyvvpsU3ruSDc
sQCvLY5o+gUQSYK/dieY1QpmxFg99vGa48D9WQz/4TT6HhsGld1PipI9utFxN/44
cxsQwnlkzEDA6UEZuzoi3F4MWAXG1FLHM6SF7KPETD7gPp0cXUE2SKhVHsuanI7v
uk/KQ5MCRWMWzE+kFAM5l5qT8WYy40ZnCsdhucrgJtErvmFseZuFfu0YalOWXvf2
iPRfR3W1hZphJQUJKnncIL0fcGMRBT2UrRUClSS0vRvDD2tGRJBRVvG4UXgEsoMe
hyDbRXkcyu66oY6XIExpSbqSeyXYcPbfV9OA3W6Ia4mk8JXX7yEj9bArCxVX7Hox
6orVF7HsFId+mrv4FvOUMeuEeu4Y3NXhCPzp+LeUBhMAkvu9XgxSIL0NAr3oCYFO
9o7ZQfeF2LPWfsGLeEYJJKsr84lkgkpeSYd8TNewQYgEfHR+x8yVaqWWHDiNLeZ0
p6xiqVA8TzQKzJrRSVpZMjaIUKQeNOrl76nk7pIsJZcoVRi9jObQocMon1PNRURn
YfzVtsjJzxgnkiMHbv405rVno1dSo3EytzytXbYrFWL9X1lWv5oZCj/l4pYjuuE5
U2rxefmC5oAkHOo0JuP4lQvLA307pjlNNqcnPwmD+vcaMsDQj0vxX13r366StHsR
27q5ztQlrJ18I61bfNo1mxw3ofNbD/N0mx1YCYCwdCD8jWSIY4uKmD68tBM2I6jQ
Ap7szTgeNqGLZ1XvBGjhzzkisW/I19QMJQIhIUmCW1lLZYHSUaNpNSYDbdzQasuu
sQKy72A/55lIQ5K0/hFiFiKXuUMtGSZVg9OUCJQJ+kAld3u0tYmwsayk3WuETSnp
eUhwFda6twQ3S1BxZKYIBK3xt1Gn3aaM2dwKSFXbr8vjLYVqOW+s3oDfGzscp9bJ
ZUWh4a+WV9tzdsZSTpI0wp7O5CCQWDlKumXdFWcBDvUtjq7zPy6/83JfkbDl320z
N0R7Fvi/1m+AGkjjEAe76KuXIaf5GA16KPpj3ZdyNhtf6C64T/IKqVrsdf8g3uJh
GB3CVzpp3gXxv168zo/lQOGffDBaDPlDG6ZbmE4VAD0b3aJwQMxor63/bYvK9UkP
Qzl/yQUXgble6sITPG9fPxLB49+d4hYi2zeGLgmNnK1WOa5jxI9YhgdHTjFhkj43
I/XK4wGGLqxmmf3iGnR1r2hNCCBy/Q9LIecQtX2thIx5cYhhK6plRdvUYdW48Hmg
A+9xfBQ0znhqmP9CqOU5D+4L9e91s06EQYWCIQ1PuuPm1RhTNecy/WJ06xGA52xZ
HycIz2Z5/Uwdg++CaZdZFm7Et38waBidWrGJA1ShE3FEmUW3zsTZfcu84KKPtJ2L
MkK3MqrdqL3jm/b7aMVs9//io0fMRVrz9i5zW1yaamrzhsk9E+GgyLfa9oWZF+zt
NL58FD51qhWBRtcCQEpAtevPB95pEy7XEKIimywue4R3qIvrIt9Xp+aVMdan65dD
iXfRJ8PU2GmxcpPiKoRxLxhDZ2O2Len5pG2J5Bl7Sw9C8FBiTBuZHChDUtXCkiyL
nXelZpSpU1MJTMQfVtYJPUTviPDotxnGWHhZ6tMFJ+4RXOitA0MIFzMDeoFPw5GW
TfM91S1DjpN3KPDMyDRmj+/HBfZt+d5ZQgrNLMK26D3fpivOcp3cUBnKymYxsY1r
mcrHrl0ENLBqIJYdFY2UAWY3R9UaxA4klkberFxW01AmLEErE1Ylj4KQerD5P0Sk
NkRWIuyFkerioyyYwDx+hIZbIlxevV6OqGKGgtLJkubnLFooa7TsvOBjhVVkOn2C
RAjt4Yb/s3h16qpkNUOdsnqbO+xpSQwzK57B0ysnaVO0Nr/fwgOnlPWtSQXicRPE
hf3SHClT6PmmgyOswh+pYa32bMD8CB8TXjQbJusbIjh6Q85jYydweekvepkUAY9N
2V73XvlWnm2ioO2IqyCuKyxN5bTQS5rNV0Re/iOkzK1zeJ+cEnuXPgjXnt0X38y9
YmnIi3EggY3aHWSjQnht3dQHSlapt26e72tzlh/QSpdYrPdwmaZeP/MbRG+wWtIN
Xxj4K3ugdj3VN+jdvkJAgvz+tMn+Qe/ghLNaYfTGoREh2xyCLNnA9dhiJVRPuIXk
KOAh8JLi1+qALx57MrRAgYTkSedpzxWX55smf4wFQC0U6l1M62ILKVOgmnjClRka
34iCxApRL6xxPS90VkRWEWtCibzvIsPVMRsR/v9tek11fDb24y9KlNC+3b/zbnXK
S0zctBB+F+4btIwpyaXRswZl74L7jLwdHi/vH29ehG1N6hBcHW69ezlCat/XzEAl
gyDAN6cT38CH1rPsiP2NtVm+JAqwmzsg4MxZs9pccjASHtjd0j7gxQ6R2yuo0K8P
0Q3WFhffEh4jKisybRwFEwGU+TFT+bRTutrVTw7nmgmhXqWq0yg3l2yO090iIeub
z7VnOUftVCRe9KFG/cTPsQMkTYV1xIU0yZyYjuwlMlwTE+tynKbD7sHqufzU+6fB
e77nlX2HsvlDG2jk0M8BwPZZIXYVJJJymS8zNmpRQGOBqTCgx0a3aCnfwbb7Z49o
uDYpLaZy9Qm5tYGOfjG1iYB0s+cwqTjEVmiLLVL58ywrLbUiouNochkeWf3nL/wW
JM3ra8S62bQkzTm13tyHeao4cmPPDTuPSkjHNw2ORXOgntX16qIav0/k/Twvtm9A
wA58MpdPDmWTczJ13Nhr0B5AHlHDzMA1F5NnGSuzu/Wf+JxxKhFx17QADRGwUPsL
+6Ro+t8eLs5YXTz+5g1dguTBxPWKmSfZ8Euu9rx68Z0MpeB65DnFT+dhbx7Sv290
1KbTo+Nz/pBDX3Il6ykDC7uWdgMaArK3+y2u60bAXF2NLrcRLKDSGFXmENn/jK5a
8NtGmKiru2jhYhm6lKzrjSGb1BLlZ2yQg79TTQFU9EHgqtJ9UghNuZaTnH97AWwG
jVSTIf9HsXGu1pwti4AmWfj2E6jlM42MrwGaH0tk282t9rzFkxTAYdj585y1pXEj
4J3ukGtHo0vaFd1x+I+DznLfEWbX4meYKDR2LltkuHnGDiX7RFjDdnwJ/ouPCPh5
RZGMpg7gj09YvXwK03OCAAU+hV0ZCPakhGEfBW5sfJBW7DTR6WAqt1bPPaVaBZPh
BGvXbtqM8HhFwNVpjXsY9ju97nLxHUxJQcMLmEifv3vy0DCbM5x5QWOVxT+2f8H6
ruWGZCSMKdcCbTqwjjagPAzfIRuMFquoEDbdvOIMn4PnGmDrB5fjEBcw3v4CEapz
5gIIrveeHFWUw2BvSTQx+dcfzDil0H/4cZRVlUzmymYXoB1gdsXZsGI4RVNTAuDC
/H6AzR0sMN+Xx+FoE8efy8tJHDIUjMUGsP8nCjYuUBlv/UdCTeIi/dGQXCilMsMB
4EUY9PW37HG3y4sBntEZyDRQnbQnYTvx+h5gP8iUzJWz69VW+TrIrmY25gs7JTPc
AQiwiPAKjPhhJZdU8gT+XLvxQL+WWW+VDVgtGUFdHp0b76AQST1lSN84PGmqhF4x
bB2lXC4FGEo+Y89WlUfhRecfd9Z46JCh7CC8htnXQVZ4lBU4l8rZFS5w1U42VobE
UhKL+ca/Nr7sRlXKe6AJN4HmelJwAwisfr+3mX07yjmLTB/HGAc5LA9co5NfU02q
qXqFChtOBpcWhNSYivEYnvfNTEdExlrWU80lhMPVxfuNkklLJIVeTy8XovshVEQH
iqRo+jrdxBRiUOQ9SuBU5e42MWunT8XTW0og5Jk6khoHSJkOiFuzmkO93E5P1W/U
BI9JotKSYjnwHfqA57OfPHAvDbKu74mTwOsXXLc+zHcdGzdkcgc1oW3BhKT5gsJs
3JmMJUeWYKq0IgPVf0D4kifT86UvHk2O2NhUFQ+9jlnCM5KCYXwDjzL9SN0wHua1
W8g1hmCuGHH/fpR7wUx0D8ZwyWod/sagk6d2BDwX93kClszDSy+7Hb9SLOGXoBKZ
7dTmIy+Xn2PSshk575QmJd16ohg7Bvbk3+LryJckMo6jEWUeNqXJ70x2sRuH/gQa
o5wSL+zZ7ecS9z7qCQU1R3hlK2eUziXwa63fPfmgpshO0SB5z0/wRWkeuYvbS8GS
k8nqbu36KSwF9AoLwiTyfg9384gEwSdJUX6u8elTl0G7g4YppoTKFsHYz3FOpbrf
J0IuE9wB1nNZHWzouM5Ja2HwRk1bo1sO4yvos07sb2HFQFV88dckOvfoDA99Bo4R
0IdIb5KW0soqgHls7xgz4R1D17qgw7pAVidKD8knbkq5Gc3iBPo5RPG9RDOJEZWW
kPSRmczNgRtUiApY8o7W7S+LR/TARaRfLWaEtZYdcDs2JeaUzepjwjDbt5d+nabP
ZalkLICOncO4jsFoUuO1p4t/Y/QBJvQ/lwDAjIj5WUAGxp/CramJhvM4PHK7+wx6
TXY5OkmF7Mh69j58VNS5tZhwey1d1UqmHLIbfzdXYrXABJTb9826wfMaLHSx0TFM
ZIPaL5cFCRlAiStMA7y6yeIlKcbKigeaYaCOTFJUuP92NSpJ7wnU694uZTNe5oRO
lXQ4i/XOtKHIFBPJXmIQv6iKW1mE5IRO3MpDCsVrhKhEipNA7/Czj0OP0ga274dQ
OdUpXQIJadh/xN1jzn8ZOpbNXjHI0EEGQ116DldbxIyLdwvATPLPDZokrzamGOFL
t8wfnsFhmcLEz1NobNBGBUruhkaHcyb/LpTQM1MgMkHFjS/IIq22idBYH9rF+5zO
e6AhJyofwtSZxFaI7DVySCTGLNdeiCmv3RRz7LRkG0qqj/qX7FiYQED5BMhw7BTL
WRTxILqwzi8e0mnIvt+8t67O08LqYRipjzoUDr3f0laZmCvSinv9qFEGPPyWbO/H
pyMkBPvyr1AFUwerMQXv3v3I4/CJF9Ehv5PNEdt4WO3TBSWExCar62dLRqNBBMxk
jPcZHp/A38yPb+9AvIHudPiRhpTr5KCXuZ5aN37kADUz2SyDtwwjRJp/1lRD4TYC
f+q07JX9OR0m2nFB8SUL4Pgk/OypCifM/G975nNJXEtee5QpmtZs7g7panSRJ6Jb
rQ4TMm389U1lW4gSZYzRgKPt+hb01qly7XhA1LSSJSe2XhGACO6qUyNVhkpsq8Cb
prRZVeIqjT30EW4RY+Pw8WXCxR9YaS+NYS+wc5tyiSw2sj8RtjtlGxJXEDNE0PY1
nb35zT+2Ck12VKIHSyV0QSBCMkPoKAD86vVjaJ8WrcVPxiyvztEhkPLb/dLIosdv
Hr5jQSTSjDqVDMCksmaZLqHbKrNHON3kqHgjqIQiZx+eq+ZD01jIRd+TMjYGT54q
ThnonClrdAJ0q2qBmm0Svlma3vXq0w2KHLpk8vdZwH5GSFt3w/3i83MFlSnJRpFV
nDJ1MnapwA4EnL5Vr0rknNBg1PHIV/ZsVQR0yot3ukfKLC59sh8LN6LsgWqWfmRO
pyPLKCQDL9XGP7jxm6d6dkfGAAB+oFwod06Kqx64bLAUh/FsjMMN+WwhNZcoH2xK
R9OunmWEgBOwCOGp8dWOc+9eQH0FQEzW/QcNEKRbK73PNr4slBAAdG4QQbizr4wL
+bLceAjR332yRRLuz639FKgQIZkdfa6RHNAg9IPHu9Zv5UoynIERwJPGh9VmuJH9
uUJWBsz7+D7l4YkO5HG2O73gZoQb/mnzIaYVaTu1mTALU8VD8TcylF2KO+oxCpb9
5Laf2JcgFQUDtM0CfDJbqb2VVTF2yK6C4gtYRSLNPbk+6J3/5YFRyuFCXEfLhYy0
t1wUGbAdILe92oR2KPemorZbvBalHP/ZomA+cj6V7WYZEeP5dxmgWSBGtIqSkaEx
6HRIhI+Ar6vvItcjPK4oTptrUqNsx9Sx2VOzfZiSItgLYvHcLO4+oSl2YiWI1lZk
OWFsHHTxynaHPjqi6DyPnKv55sHMthQoxe6meIU4qOE5+tQ7K9t6n1c6NlYGFVPF
DJzpeJpdoUTL6J4cYJsZcyy8iTDP35HKYpSYSWX8qMyKeCGQqWDysGFaneuuOtgR
wCchGnCMHZM8Hkbdae6dxD65Lf2Yvwmox42YoSiMtYlelgo1cQK/p8O0SetjW7tA
6BkCk2cLAnJ6bhNOZzWlCXjdH2Ywj69gqz4Nn+TvcNnhv4EGDeCWs7li9xQr/SUm
1w9pjwIlt5fufWQ7e6NPsovOy2bCLCV1P7DkIKVuSENO1EVnWvrvwjT8Vx/FhBly
tbBfjg52l/7hWQkol+dXIiWWrDOFlbk+O3oSEo5UD4H3KyBoFmP7VBT9FIP44bHI
Mqd/jZPuLvp4NV3ivUTtc8e4uWjjRhE8X7ldcR5oCKfjAnLsu0921N522keASwKi
pfqNPcg+iiFKPd6ViNX0geL4U5mcc/yQ+RRRM4tLL13ooiPk4pMdWnl8I1+Ed7D2
bIa7MaZeVoI32TQI6byI0YC+vdyq38iScWys+DGs3A+Lyi5rAHsqepx32rYYEzZK
EGxXdLZ2maH7kWjaxQZSAt7My3fwbTb+Gj9fs27s8SUudkDdA0Br4a9FAbeIvzK9
pduveCiD5VEOciam3ookmCBbeIaHMt50nLXXLcGjfKID6RCMZMdyiqEh5OJ97xUU
Z3Uk2zSwBQ+qEqZCsjb6A8guU40e7m00Ph+Dnw5FoarIhRcn5fbwsjUoLmZLQd4C
cdmTkHbKvKGZNoYNxeZg69cXgZCAQku5sryTXLYmsDUoeu3ci9JfoXhc1NIcDMdn
jsDhvvv9o1TnvR4AgYu8hhIgMT5xd+1GZvS7TW2gpRo+q5pEiHtpgi/u5Wua3iHz
0RVahs7clsQIU/Xh9m5oMokHW5JPTFr2A63s3LxegaWMiO2UeUQEKQonB7aNC/I5
ep3i/2t7XaqCo615wFG8A4OJhPF8rm2gUXlHEUJlYRZReatId3YgKuYlc0AViqLc
cbFiW47v0Qij844sH5ll7wn4+yniUtLtiZfk+regM8Qj7qm/hKa0QrXaqAXab3o9
gC6/OhyAdLY0CtVZOMul9AMIJrFAio4y7umThEvU13/lnaZ9BYtqMIcoH9Sn7U4G
S4BrwWBNXP2BOz3y+S40A4VeZQJBe1pv5d6nA4YdAYD9RwwRwgQb7hMXNz6pVkDJ
P4HjKlXNiKrYpdPwjBUjh1aRXvgc7l7CRuFrGOC4Yh82Q7RlcENffUOqWlJRPFHT
DhINCP4MTiKWAOu1J2RSg4iZkBmZSRmluc8EFNDaLqCE65qYhxuy0LzaAsabo1b7
BfNsDBobQ1lhmU8nRdRwQxAWz9k/xFDu8Dryw2UMRFNUCtu3Pu5Q01pBY3hqjwn4
wro4bKjn5r8Xt5pe0GLpsD9D9NzXkaAvteU9m7hCDKmVrQe3H6pTcvJTbx+gPcor
LTNI+03i5MsT5ZBioCjSCtcxtfw6f7h1iDmRbc0x7GnMyFjKAXiPAmkDyKuOjNLm
TaAav6YgiWELfLX1RR7pSTKfumwsXCm/DkENYO/mlDQhvnVUSLcNe5vPyKvVo11o
d7DC94P9bmyPPX5y1ISA48sVeffomvWdwobjmTyFcnnDpwYizP/cZ4n0xdDi1hUo
fYHzBCLHk5GtUa55yea5Kubd42LB2erA1Z2ocx1Ii9ccu6BxA0v5SjLXNr0ZLD9J
I02GL+13t7K+ZzlobU/MC4SbtCCVL6GuwUEG7X7w917hZ15s7IcqUAXCHhm3Qefn
l7mZF8iFmXgDoCT5St3qRJ3We2ggL3Z5PPKGXJlnPqsdpKNHOCjL06L3cmtq4OQ3
9EasS3HpJlI4UXCCGQLidy0luBbwN6HxgepDC3l+SEQY0+222J/7CpUtpXzGtoWa
pa03HNuKvUJfIxGxqENj0sW22/cwQylxdzKrBnMOhCKSXmeeHs/I+Z2L+vaeGphm
JqSYNcDDdRzrIKCKPov9U6VYPAte9ZDFe4cDIb7V7nsxPhQhFKNlKUitaxpsR3Ne
1jfVyMRrlSb3ZV6xVCCnxPepcXf2kOvrwQXOzLNkUfQmRmQ8NFNqOYFLrijX6F5x
urRfKSz2WLtUHRvgP0KPFzzdu+EktvNuGAmXuysIkiqFAON1Kxkp9m7TPJpSG+I8
Zj6+ZxAt/R1DFBd3gHXgstbnvJ4TabeyUkb7vZC5JSklRvfSAndCTEq7eu4HxfSH
Zc1DaodFTOKZQvDq4YAv9Bgxtr4NjOuyfq6ITHBXE0u9y9f1H3LHVH3R61UjOLhT
UWxmLi2ACn+YI9+lqrDnvMSAkULeQe8SuescIGLF2FqHeLQ3+9p4qr0RiMrlrNic
+V3EjkKqNEgL4XalytCsHcjDAbXyeZzdGuYtRNPlub2HIwJAIlwJXq3MHITJbrhU
cV9GaazjbYgFPNCbzGX9BFsXDJ/rI2h/5ElebCavPhHNj8bXJAh0dybQPc4lvfvs
xBEm7Ub3xODm/ZQwSjmI1ZZsXLZmskDuyhT9YxpfNDkDbAYwxoIpIALB1O0Du5o4
f0SOSYqwp8E7jvPkZLxgKhx94IgrDMLzz2J+akgUrcGSY1+6SDh/Yr00zB3rMNMK
VeAplCZzfYQTOh94yEOh8X6wP9gmG3hHIgXNV1BvshpOpzDP2ISWZmR2vB6NrI6S
La2Aq8KadkjOL0ZIh2AkTEg+he861jAau8To5l/nE05FLsGzZO0CCBgvthRHbPE7
e894Wtbl/DmDWiweKdrUBjkDnAD63AR9BYzLW/ptZlEa6dU888Iw+/b309VRgnus
TFeh76SBXAN+GM1fSdl1BtMg3XDc7ZZps6WOJOiF3exmULMgP/TkvScMFFNq/NZY
f+koz3MGHdEDAoDx6FWKgQKmTHOhsOMw6jzqh+Zu59THL+vrj18pwbjaQRUR1Nfx
L4zHm24UIFjfvldkwjsH7F7wVylzwgy1nqGOQbGMzHG662RlNcJpDOkeb7s2AvP/
3pbx27s9nyvPUYpWVW+UEriMdBO9+Fvo27VwcHRpEaNd96MqqwbLUdgnFb4dPqrT
nVxQL5+sTgdBkQ0EcrjGFigqnx9Hd6wUmzXL2Kny04hoUSoG9OPGmUX0JAySCllL
Nv0SCbQr0Ch28qv0dmAGcp4Ar/MEBucxfeZD0ZpFF3o3imuKh7MC/NriPTCZ/J2r
ystlf0pE4BO0PbbdSJqmY66auHUY5FYKDoogfEJA/9DPHgmzzkcUI5bP/e+5pbl6
JIEzWX548T6zMmp4320ojfbwSqCqBSRG0NoBfkkYRRwWvJcVlfCtaApMCFgddiD7
Hawj/w68ZPBYvak7PnKGlYM3lGrLan7G6/sE9ST9vFWn7kPALyVXjfwWGL/5KL57
rb7LNbcW8dM+FdTZrVAkgoT/dfYy2yikpqvTM9a7fuqlPfH10BGxMMfzs/vX/A/f
zQLHniyZ+7X7Qk9cs6ViU3qN1AzLL/j9NgzFktHTGonzPbAIDqnA6/GQJvyDUGW2
wKBM+lwgk1IxhADw+sLk8lbp9J05SxGE8Xg6e73Kf2bQ794pOnU+3MkfIFwYv25U
r9kcKjdz1X38plwU46cLyebvK2mNklXJ6Q9Q4NEaPQnWy+6RpyU/a7EyyixnECWu
veQNtXcW5q4QgPLOTDdR46j/wrRMrFufRMp6gp4zU5GBUiqXLRdSCtI3fyaL3IKI
PW4pPHPDs7KAGhHoIcHubPJ+F4pxtwwir3sLx6Kr/lI8P8pTkyyJmG32N6aqFmaH
jolh/JzamILt4OhZ5Mdk2acViT1iSJ6mx1EsO/yC3NU0eD9eWJf9PyETG2cip0Zl
P5vx6FU6vOasomkOdLB2l062cLIKPz8pcFEePOf8oDSksJgm1zYZdWfbHvnfD3Xb
WDXFiayxFYcCw8yNqyRG9jNyhJlLSND+QY1yeGD5QGjMHmv20xH/1w9v8bItUiaL
W+0NifxwgHdnFxwYYecw4IyjlWgvD6N60enGTGNjOjy//0NF+e6VqnnrVbI+rcEn
xdrFGNERz8feu6z2pm3AoL3RyIt+oQPa4lkt928BnDcMZNiuayKVBkp4tKNc7pHC
zSiRRXuLl/g75sYKJg/ZiKznIRAzgiRPjnzIWmQQ/g83vRcl+PL2wq+bGRxPbZIW
vksMc+PcM4o1HQfqoAOTLVkCvE7f4NnH+K94Xn0dNhgwoWHSz0tgZDWy6wOmMuLE
2luaE7BtP7CNW+HaXCH4vXZHOvf3mD1WpMqeQsanJud1vwzPyoO8CQNyHG5DZleZ
z0Rssd/AH/7bRXawid1Gq+IZBi8OVGA9Ao3SuUL3BmFCWvXlT+uq38t9qIqzJUf8
LdbSqz05Tzkp1UzbYFRf9UjWBnQppg8Vei5EkSiEUSvwyNlkf1W7fxeX7uQOKvtz
JGimfF7x2mIyYK34sxISr7CvY83cUGVhuMlVKHDaC+OLTMedTlcwkJCULtjhqSyc
qIpA6XycjFAUKvKlcrm3u43dWGdmieV6eSfOcXvExvc4VvfrkBans23lGopIh3BO
kNi8BltQPacJKb4pd0cUtuNT4EvpwZ77zBEsnuz6ombewpbQnhIBxGlVzl8lD7EW
2tSI1L2E17+XoxcWjqc8YXeDYWvA4To4ZgFjaJmbdgY/simOup2lwR2QM5RcFNee
Uie1cCgdgYX07vKhNa7+KWN709wPbpYYYXQE/4qamuHWaAvT+E+PHV/27eHHmbA0
Fb4DE3Kh543B2pc8BGE8tQ0tzZxbRiWUMKCN4v3kS22om+LGGHaGaS9snBlyyHKn
YZ4ixwq4TcIV5rddj7SaPAVxl1dHwrUb+d6R99JHk3QrtoXW5Tcy4DjdQa7VeRs2
goa6riQF+UzcP2hLnJ+v9xFVrRxffPgP43LR4W3S81RIFtkmEyhLKBH5vOn2QmkD
7ptM4rmLACVuj931rX83q6/Hlp4H3yGcBHFEIEpcY+OIQMPprS+IxfA44MoVKrTT
woHA0YC8TCBH4y3peTrhuAeGeGurJf5Jqq1/eiQL7290ruUbU0n1W5bcaMK9dFDD
Ee3OQGW/iryBS2kuTVJ6Xi0Vpph0MSO9hpe2iHM1O+20EijfWFn6o56MoH+RL8Lp
INfLZVbmnNZiQ4ao8hpk/9/51ooOGJsDoWjln0TTm8HJ2U3ypCe0YPZSKc+JqqAm
o55PNQUkna5Bs/Gafzj+686j5BjpX8ZglvllyeFo4IwUgvMbZBOwWxtc0Eb5oTWW
QwiWPyp7Amqy4purha1PIKB9IdcDdU+NYAeZbWX+AHJeHM8Irdsotd1OKNFkxzfU
EZ9fwonim/JYpPHjWI1K3X81+NyyRq+hflXgC/kq/zinsehaayYif6fUz3WhL/yb
k7NacPeC1SI8Zh/gX1jsoSDl8JW7A35F9Bv/c1Y59NhhwEvElumkQOZYE6QjbJ7C
NM/5cLLqWOHbqbxobUENXylBniw0bM3FNisOiuPZmfefdzl3/4Pnb5FYT2hbh2tV
bwfrrqPTvqxcZvbB0+jX3PxYusbkAfImy1SwrZC84vxE+NBXVc3oSlwnQ1M+as5g
k9RcthkRfZ/Tsyv8I1cslYNHdssSJPZbZkGwgy62x/dWR7mlTryHrPqxOITu9ye+
/JwD7tRMQ9UWfkQRT0XcHkTtKgfhmuHPRWQ0CZtksbtnNGa0f6+ZQpYYhN++KjtB
hA4RnmR3VicTT03SLpiEihxFxyJqjv5KpZUTiAjNmoWwpxdMLqf+j/13KShKa5l5
oDOH8BygsZ+O173bSPDAvI2OOxra5rfZXoH10wt6lZqTeghhrMvBf7n2FzMdaHdt
hV3+rewvtsEdxSLwY9gSfVuNUkY06AIHS4SRj03xBsDluajVw2iMzzFrIojo6s8r
oT5lzU+itmM9OJcSoUMT281i1r+lMApAoy1OsC7YUhR/CejtDnk0+wDhdaRQYPdZ
odt1bWZoaJwfUz4lYSY98EZOqinDdVYn+MLo29YnK5HGAKdm1sFlBvL9nBwc/xX8
ebxu5PEH1o+eRu51J/eQiZWIFg34V+hy97JQi1+BrpgXrldX3fYCGT+9/MVuhyFP
JHenbE6KJhGW28Moqlc8xHIECJQgAgkqR2PbbXyh7oWse4Y8bT2peGY5h/MYpbpd
rea45ZdIZdtnh5Bu3l4erhcltCfjH704x5rLjFA7FNMPjkYJReLM2sd1NQTzzNPh
94ho8SNsj56+fbg2gTH+M389cjlOpdOb9nKLkSPI1Sfq3hXF+jtjlnKP5M1oV38t
Hy5CEmR+uPbPdYUDTpv66Su2cPa//5Kjmg8WhYGKQkUa4RhZ3lwRcr7fj7e3GB2T
w77QTnQSAkrFFmxCs1Kfb42UmzEczSibPn4RL7rfLuMRWU1isn5xwgUoDnsxztxs
bGm1Lgn+PHvwLVHpAMHor/M1HwDBRdoPcPk6/JIN8mOxFc/p8oa19v0rCBlJ2I/J
zOUWmShvVmErea91kkqO6Zor9pwUi+jm/pk14aH2vT2gwEB3beZJZLPU4jvzhZfm
3Xaxfc3Qz+Y4nYQ7zOrUpRXDNnQZDaYqXCnp9RYTg3Hq6W+P6mPePltNi0nr7Uq5
VoFQzSgAl4rbN5jXCOluhYqdU+mxFdA8y4aQmY275B+Pqgyxlpkx1fTgEJ4SwGW/
PLVhUPyaGDwmm+fovxhZppsj5omuWXkvnoIcQIYhKtjscdDohw3FMovYhmIxRCAm
rTmi1LMyfga+Ka6BdVZtbIeCBEZnuT+WIHT5r8ywH38nEP4rHNBUtAQIN2z/BVeA
vIC9zzaIvNLaIaDTP4/57X9qBcIwJhXqPLTg/uHXmMW8MbvlCrg70iLSlZ0PFRLC
8dNmTnzorySvxWO3rhJLiJVtix3UiceZ7m3BTYqrJLz30EVNjPeIXbQRmfif5J7V
0J0M1tIeN7BmNcV950d3vmu0y1gSo5WYWIoPrn5a+JX+WY44kMfLK+c3XTOYQlm9
kelubFYHYmcfJJBTgH4qibeTQAhp/u2djZWEgMh05SH2SQQ2VwpqWmbtSjaRJiBr
bGE8Fic2TTddHSkF/wvSbKiGhyAYffA9RU/QWcnOOAy2Pp/6rVEjH+lDva88uLEN
yhqRPXY1AwNQyFQU0D4S6XIn+xfR94IgQVFkwVjNZBUYmZ6su8QDPZu5Cdj/emBg
Q7S4WUN3nQKcWQ53jNBh+dW10eipXROxGpHgzMMa1kMObz5UVylHytzAP2Yg6JTj
tyOXP9sJ9tJGTyA8810roaZeIxe1l/+iMpm0vE5z+BI6lOR1QXuZhKq8v2x5RwC4
FV422UXG61lVZHYye20qRq4Dnuk4HDug4/9m4cXAChoV5DcgrSz/zlTycTxOL44o
C+v2S651o2FqRsy/+xHwWNYfxHr7lzZMUwWF0BA8htPMqhp2h0hC+bZXpHFaYZUA
4727nenpEp8auGAKY93v9KxM5lyuFXQJpuTse4nJGwxcZcRp/XKi0EpRBBL6T58q
Y2rAXqmwih3kw7qWrkIHCWkBnksuqLvCJyiGGOncqS0kFHGTwa9HBrmdFn4xGbKW
/80WP60CXGwzUPR5qXYgSZ/FOuCeeRn5O/y+BDL8kSpNlMGAAmLk9tuk90sv4Fzy
EBavK6SjaarRl+x9LS3w8MkUpNnJk8xMsHOSbG6KGzDXexU0IqmRghG4kOuNyfcK
qd0PzTX1HjgcI62wHn5P4+eqDKvnvlw9D0i0BnbteRuSHeuFH+2HCtrzXvwynNBx
8QdYqjkrS/WTtmDHgORtiQvInRpldGfNeS2eCi0UyS9vSq3O32oHdiS+CaJh5zjy
I7B10IynkI3R1M0P2EMgQvX6osvOr3BF3nr3kDt5awL3hJDbl9jpKRVNHWxyp2mh
MEIci+1tygTm9DpdZK3lCNjH4jjX79T8J2sy5l4WHr0/BuP1ZA/S7+PnJTxVqnsW
3/u2IuspQeRJSXl7vVZ8aVLY8hWELIg0xeFtpVG6Mb68VFjA9Z3a3J5kn3YDjFQZ
CPxgOAOxeSFzHJNE9WfX5vbZaon8mj3YyXOCoNTNtSwlfBH04MEAlcQwDX2aZuGP
b0LKnLMXQdylAiAtRChbH7fSPH59qBBPH7ukh3bxO9rUZXxVCKKSEXzOQfdYD8WE
Mhd5OrEMAi0huyQWgri5VUThSTOjs1zu9ix634QEc+/6WrJ0Jc5F8kA4bEzfH3hD
vz6O9ACCw47bV21frROcK8/RxRgwatUSK26DuM6uuus1JHcb23K3FCZsT3+lyICS
sp6xJs2zOmiramTxGpNMWPzcxLDuNiE0POERwkDOCdxElc0t44dtGB51/sOizel0
RQPCXg1I1u78Fkp9Rx5/4WGfYywbtb9iza5gUarVQHPAjjjlmzhRclPaiQzE5hSZ
sVlJw4BrZNvLUbtCAfna7L86T+o9vG3Et9Afh3nQkoU8PH7SZeKu5h43vVk6hYl8
5C5mwV5sHi3Bk/7IT5NQwwM53+SIMX3qA9thKKoB9p9B+eLpRmy9V5NYkPwBLlHJ
4jBI1OiZduskhw6fWIyXa3n91JQSmsblHhbxdtFoB+EqFXMAxoTqCMMEc7rNTX13
cekf1fkHaJWFZxNWlAuHiqN24FtE28QOQn7iiCwgcMPlWqv0kWzPMuVjoXJ6vmei
3oMjTpfIOs11IYNzAFeTFxvuqSBuhDKpsXiLjDIQRzf93OTpeLXExUFaHskQ1XJo
kK4qAQZcYdfZwqyTpwsDV6Hxpbqy+2CoT2DSzxB3cRV46fs28QMG07OurHIfBgg4
r0EHwE274PRm2D4yLP0PXa+a8yy+d9mRVUGXOjubJfzBL1q6z0+A1zk1b+qun5hB
gIGqORZYQVbtHuMyVegwwXvDc2dnbgG7SZycWgLg7okvoqdxoxcQ/DZ3LcTkcGHG
7OkTwUgDNlX85BlwmvJM5gX07UHEgHG/76mePTh6yb+zEvd8l8jE5WgIsxoxpsua
dJrUbVahHrK102fj5AFzyOMKzzrnCwi442yhbPdqdwsgG2VD6moQ995VTNekjp8S
mC84pIhebHE4KcPv2oHG87daU6xuXFu0T9Ig1TA6ARJuG4lLIh2IA5iiXrh2cKAh
DHB7prS0Qx5T5mI2aOPq6fmW38GQey9syjYAHisu4M/R8v8puib2hIev3k30yeNU
hEo/ii76ODzkOlO1eFvVEP5pteNaO/OMR1KPKUGoJEOi5NjT0DV/WPtpHOWfeN8q
59oGg+yyzCh+9ILRCa4A5yxVygFcmCJZJYJFTSLBk5qgR4SPoluE42Pwt4S6SthN
4CR7WvJFZEaD17eD76mG5jUDhjyFw2ANzmpfOTJutpN05B5z2FuDN7YvWg0bkeSx
xzMeopPJ+IBaXV+OFbzidpH2DwMbcL4IPnU6EbuSrBFIFjxY5ATj7j30CbfBakmt
pkHXrrWmW7vhxtvjNrUVMCme1kJkdAkMTKCHZZd6Kmwx0+29JeNlyuS5vEE+HLpU
bmYTksT/DXiPFrh61hHTkh827L/3NDTajGVThMBJIZI2DYDvYECXHx61A4vj+6Xx
CMxN2BqK1+/FE1tMM4/jW8e5VDItg659y/ScIc1wdSiCui6Z5yJ4BnGySiQCHgKN
Vy9XkDc7A1uD6tas9H/criJ7nFVe/9yXlZGmHdocEXkF8xhvtZyDEJ7hiPEjuxcQ
7ktL78KD9XlR0pOfiEq20NFiELZmtb0/bqghM1TXiAf/n0DSrcgcG2PN0GFneGz3
/Ijqi3IxcNISiyFu3XPeFnVGkgGnCfKPq5qstuoJVK+fdng2nurJVyLmpnHVzOhf
LZ9psjtmKQ1s2q+9t0RzTB4pzRS28qdc4LvLkMeMYnwhR66xM5RicqgVa2PlW9/4
kOZ+1KCly/LCLjSJLu7JNSB93TGjNFwGmwFaU1wH/zFGbzFjThkXMSDpHLSXB+Z6
Tm+Rvteb7pECi68pGyKavrYamvDqRSk0KVZ5IRdKzSo+QNHuDCZUFJUeYp8SOjhc
tT85lHAy/ew4ytHZMgVk9i6Mobv3Erh2Jg2tnnD2bnTDddIEhuhPJzPt4CsKwIKp
0TY1+7sKAyzOYujEJTCWmFF70o80d6PhdjGMKxtp+oa2aOMZ0ucUmE8rn+t1qmDT
wWZ94y1uspmKm5wUjEU/baFawwTy7cvGaNKiIDCLiCd58bj+shfL7ZVj6yq6IX8G
76WURKmLZ1RKQ+Qvc83eIH5AMUYYx9E23fP74/0CCVDCyddwAzZJvZBesh3qbxIY
OzAzCuakMdCWZiF/J+RGzIp3j+EEHvuE2Y92qZvvbixsYMNpVK+JJ+Kf5yG6cgIC
JTTMIitrHtm/fH/1tj8WkDjyfxR0z5DFxW4t/ELeK6G/rOHzXHNmYuJD44Labkyg
QjJuyk14zatL4TWpRa2S2nEq+IlzAcYOVhQWiZ7OadfbcVN3b1xr5lDkmoXtQ4Po
fHN3wMrrqK/HA/ec9GeIgU+9746JBxQqaAOrCLUCjoJ+7N7EKdpJHyf02jNdyWf6
rBvXmGgB27PHFgnduq9SfcuS1gGJEijVVIssqDhskywKPhDhLD2VireNTWLno9Ey
9bhZyBAZeVu8D4vYt4EmlgHorIyo5ohgsx08shvY80zwnpoQymilTD2h6fklqJgx
pb5cy6/W0MFv4ARQPyty4fsf/U5ZxOzSDnudG/pKf1pIBXcbkCvvUCmJA2eoyKDJ
mCzbCOUTSAfwpvUgaKN4FfKmxvrHtnLU3hBFT9Sj0gsJo6VZDBEV5RRVQ5IWC9Ig
oxiNhVKOlZbD+XZqBy1IPoYNuLHg3xJgIVgPDUPBoDcXQN810ZRQ6yOgf/JY/Iw6
srCxw2BoejJgLoCuGi4b2n9spO8fz6Y8QNk+2e6jJaIUaETWCWK96ov08GQcLC9S
Zmrl9w5TmoY2vZze2KxSJ3engKo1g9/BFyeRONFfRIOFjUsSoUBZ6LM7mFm071HG
XzubdcyzqZCnMaavL/x+1T4eKiTMg9cG92Mu1uyeHlT+rYaY3APtTkpMNcwFFe5E
6zFeP2gyExhaY/67kejpOaVdHk6u6uUSYpnky/71kALz1v3WltYgCSkJtm6nsxr1
F4kBSxN+Gq8jrZwBrlQ8xV9LKKmGag5BnJFcpvM0Yd6/55D1m2Am3Dj3DXGoOo8h
1rdBgzCqqVDFK+98trC+uG9Ly0mgegeK9q1pzPlG77CzaE3kxX04UoNoeJ1CqDAn
89FvNEek9vYp/7gpFTkNfwC1/IXfdYwmBme9h5a+nXOVpcFC86bIe5De8MPt3e+0
oWgPHPaBxSHoEElALiCXj56X84OaiCuPMNGHit9yUDO7ih1VxlwdF0lZPSECo/9R
P/MvEozT7uUSsqKE8hAnyfkJMqHRH6atCDmpFkTBDkl6UeOX2W8EeAOIvSG6iNB0
y+OM0FV9fJEKsW8tRjeA5LRfUmrCLCxNZjqA8acMEEHIOAjZUC/RMZYz4lZ+L1cd
otrlu3D3NtGC0y/ozpeS0gqZ1NLXcD3qg0fw0DOme+EznB65ZOHVaV8zmvrASNwc
x0rdphB67pfO5aoTX7lEK4kBpNLV499Um+mXfL7s+T+57O7AglNkCSSyjWWVzM1p
kif9298BV86ZjarsOxQHnN1ecG6NnNRAkVbAuFfUopsBh70uLGhrHGnUsxX/dCRY
4bKSeqyVxsSfnzO+VlKyaWwOMeMHpOlgkKIb/wytKpJThAgOJ9oRkzr7kSAHAg6U
idrym0Bqz14SOYp48iNDRtdUO3LNedUrHs34P3mNsacPazwjRhi+87PgJBwxx3Mz
CPOdzugiV7I7lSfQ/Qkna6Jo6pqcm6hVYD1r9D5WlMU/XNYgJl3ZpCsQ2bsuSrNx
Y1Y9ZZeAZOONvBYHJuYMw/UhllifS2ahyt0Gdj0kYb43Q9AoIBM5M8TjTP5qgS6I
fGqYd+3cwbkNJ8z7tIxMQq9lRGE4gaMk5ntvc0RuFOeiX4l/4yu1fiA/NPdVSPoc
IG4wYFtfDmihBHXDjPWzdubr/WaqV89wjEubkfQCBZ8h6OM8uoD9nlfooNMqj+d6
Nrv+FfYIq61IWEyQGrGTEKrXiG/vBhnAuFP9SfJ23Bub0tM+8BzrM3vqObwUIQkx
5H/jbAHkLtSUuk0AiSU75JgWwx6Mk7EVUuBYj6//PK/X0yf75mKdDdvVShPwTEBn
HUCBGomKMUDCo44kdlLKgvYeqHCo6GXvYh+c6w28OBI9zzasm7I4UMU41kSnx473
Tttt0j3apMBEXqabN24i75MUgt/9uCbqPXDicwjCwMF5cv3WaaCGz3c/Oc4pHgHA
55EcLcGmnIIHJiqpPfblYziWSzEsNgbIFrQmyHyBriieZZgQxP1+gNshiA+zF4h4
Zu+vSVB+uMYQ2skm9EEDWvnkYh+puXQl095kBMdeSQltRoYHW6lChGrjhRs3f3Vz
3VYlJKPRjMqamVHJz3OeCr+HDxBuB3BwWpkke3W8skcW5082biG7xNfKVDFsTfNN
m4ykXZbvyTX84K67nlyRUG5rKI1vaKanp4jSa0cXffqrPSdzWePh5NI4GlYfIBe9
/bpJXEhqCX8tn1TmL6gKR/EkgnnM0Lm7SWCH7FfR/747iSU25V/OeB/re3vAQGpA
uLklmXxxaYadLeu7/ScCoEQPygo4W2xWA9EH/Ng0f81ywN4BHm/KnOI6e4sDkYn4
zmbl51TWBI5LQwoYpU0vi2suo4LAq9hxatKP5dtzwl5Z7byIkim9ixff+8UjCyjH
hR4Nv6iip7ycdjX8CJbq+89BugpLCzbRg8JvrLsC1YmbgtTvQvKO95YD23avE3XM
I3K/4TkVYTJk3cO7k/eblqu10xnR/UoeaY6Gjhglp2oJdcwAuYRRjsJEvH542BY5
ZF4Y7/yWov/vGGFJDG3/oFwCddD4/DpIskgR5PCrH65t5Mc2sKpXi6mluOq3X+Pd
49fapS6LeqAnuq+WTR7I9f9L66oAM8Aw7easpUV5SGZKFYRGOWe2vEUKzAXrCYIM
YzRxmEVKwYaXF2XSg9wyWMEuq+aG+/jhiJPR8AkTFD/vapi+PXtRFUy767fAha7v
eywOya14A1Q4SbAJu+xd56x8J+iLvLTDw2fOLoXM2Hx6gKZCVJczb8RJ3GKmayG5
5FEdMzd2UQhNfKhqxbkHssjVNNgx3hnPfFicZUpgwl8dxPZcp9wOZnhqZXb08WWF
BDh6sfXL7m+wsKHf3s3D0+5YVbfmf3LxD/tn09p6r+deLNDq2bWBDsyaZRg/h6d2
hJl1wZAd0mOU0qKlu/WiYKgLgVzXNBkUN49o9NrVpGYSb5DHohS818fz3LgkwA0i
favmcyk864P+qjOuVfpJF34IWi+V1auZ6iaUQSCqBFKWG7ooep9jBQRYUnnPd5wo
5jJ7CFTJE7zfazzK954PRF0F6A12NgE5swy/RLjl6z+YOTeFIPMqoLwGqf0RtzXt
sXRjER4f/gKgSKZSJvJewA1NYxwwG020sLFLstyyOmQgESHG/ldw0ZyBAP6RvYdq
F8seExwvyTHKPq8bhLcb4qXnP9DuvOwc93PR3uAlrKnWim8h0LwO+rjLC6EmqOU+
JP1qu53bilhjO4V8kLXPxrb7nzg+8IuhmfUwrDABZdBK2ORHQOlabqgt8fmgWgHl
Y/j4z0rLSwVwplnxus9Lk2Qjq1NrGFkz6+NLe32FWQi/AoKbWPWWxeBap0X+Y35J
Kx026hPWYt06lbSH/FPoSaYaFIawFI3qFw5Byp1PozQg5vtZG5k7uvXDs7ByOiku
vyrOKM97K+1EcFdMn9/jqjqjfuRTGkYMwpC6dJAfYwhtkD/06oL4nISQubf3OW8i
JaaOAy+ZyCUDQwkNPQSGKgVniyjLggdauVNxjDvqiZKoqomMY8dskIY9TYagPhE/
PAM+NDj2TcUQ67D+SGLh4Ki2rWKBDmnrqE4CtqQ47G+GbPbhRm28nKti8YpXuSBJ
aMYJEO+lUFYPulhiR0ZRWRfolGq1KGaqHWq/IE6jdKb87VVUWoy9tf4d1ctmBW7G
Sg105sDyYNW/GMHl+wXWrmxu7pk76RG7i/hnSutVaAoSkG6MKyj9cU4QpqlKOP84
s0poOWjzFkALCC7Xkkm8fQTJemGIDWxP+M3XwzzO6zjc1OG7xDvtP5PoZBuZp8cq
060ATJ33dBe4I8RXqv1nC1ta5Ex2GxoYkLSxoX/19I7GTgAR0bF1+S0tUw9vSTMf
mM15I7sWYsVBC/36laewOUxPC9D5NNFkIUze69ESdT0MN1O/JIdkk20+U7uhpuiE
iZ90iC8+75FKePxwyUVUVRWlPROsoxNFmPX1YpTkV2nPmoETh+AzEgpzFPxKOfwe
QFFybrM8qYZqkeT4dg8iYx8HQ5NiffxYp08wBZFdXqWUi+hQn28qpotx9gUTILnD
DGEix4z6eNa/R2s3DU5wmKkpLj5UDm2J3+XE9ZTPS38p/188jPtT5D1bZfMsh5TF
BaNJlU2vxmfjpL1WNb2giozd3lhIOw7JgQ2awAOkGVwlJR7gwmVgr5Qq18zYS3st
33tPH2MqzWJwxONH60vpfbOFDrqRyibRWekfn3qSzaeDPENZBjpzZY8xM/tlO7We
Z8m/IL3Ja+236Kry8ppSkExdBVUdSiDygTBHqZC8Duws9rSRC7C8JZ8keEmPPXJs
XnLO3/3kSusBUWCCwRgJCJQgzHxpWISXzMGGXyyST8ii7RhMLXlcwJubc735+Ye2
ziDUjKuBLcPX2Rg8ryd9wZtu2Tcq5DJlo7DRQ3Oz8Jzba3i/ifKRLSg1z+Cpu9R9
GjmXGhZbawuHwbULuQHPZfEQf+N9V5Y9oxuwIk171A/XEqzCxV33+ectmLlXTabP
ORHxovhqhJwwonFggyaUOJq7MPzgroHAqwbo9Y6wjJf+FcQs9YZfHY2at/1VuEGc
2JmhMpnk+IpnuZb6jAMoI8PRwwZu17KQ+mjZXylcqclnpz9OA5wwj0ZLYKfJFRud
maHw4nupyc0OnX3M+6msBlhEbBx+31jTRTufUxqzZVV6DSvmjqxPTEJfZpz0jXRm
bS+1N3aGIzf/HZBkwDanmEZIS+RaMS5g+E9hlAukmfBQtq0ImTjw4rtd1BSDdFm2
rhoRNMsIYYDjQD1su+r3gZkJwcsHuonMwwEbZ5DZoJyAMWh6GEac9UNORtsn0wP+
aW8G2nSgYC0hLSyVh2ApUqFQ/4U9EwTdHBbU7cURgwQGol8GghY2kVsv6nCN3VWs
ll/Xe813Xl6CKz7DS9KG/u5aTqFi4i62H/ikWn4LzBKQoviNPJG2ige4w7nvPMnN
WiHkxdp3/3zF+txsRculY95KDTzcC6iXG7UcQ2WrZ8h+k7dsAI404eqQfZBBWQQJ
s9Zqgzc1qkEKqR6Mw+JMRLCunDwKd3XqxHbAvqJsDo/ebvb+AaH/ENUhCnmDtukI
DV/Cetf4R+be5+3bQxIV46DqK0f8T5Ph6E5iW0Ide5LH+PTsv3vIWCEVpJHMUrNC
+kHk9OlLgENAoZPmq/YhpciFveWk9T3YTYh67bG1cCS7poUR+K1F72IEgn30QmTN
FJHQwqcnYsRf2ak2LEBKJS4Lo6XQjdAfsKPrSQ/+j53UbAOIpYmkVoDBzsfI5jle
Yiw0qZq6X7CtPk5nln1UsZd4K8+s8AanTaZQpTFK1Tfw73QVThx87a83rr1gzwL8
cnornqGHtnsmV3yPPyU9MpbTmGUcQBbt7F0z2AxQGL4abmreaODLVTyEaOTcr0WL
l2NjIbr8lxBqN1UYp5TOydec8q+nsAIbq05fSP5oP67i3JC50G2XDek1oRN69LDs
69c3oPokoU85Bn+ri2kXVNihtL5ZPaW+RGJVUj3PRpNUjXPZCd+yuwvP4Uz6TR7F
OttiVpxVf58Ys7RO9BZrCTwkUfBPXeH87k7CWi5281iucTGXFndvK76u/fHL7aSm
KbhCllAuZmMhjeIa5i5P31tGtqG1NdMttas0nYlN/SBiYvpgrFimljhDHHATBuF+
8L1hkVt+cNe1qlOFXeY9WG6NW0tRR058cxScctVL5WJTVHkn/MBGgYi8KumUf8sg
wiEXOZm8v3zgE/GpJX7Jkj6i0ikAVBX9wF6RteWbiVDGWBp449FzzK57y5pNEndE
kyHWkZrl8MPstgvlg7wWAaOMjVVuwSrOk+NjklqiA292UGPMQW5ArN8M9/391D53
jnin3zDLjxvmM1YVt2WiiTcpKyq0fmKXW+l7i8440ntI68qpIiitMZAzH0ms6uxn
q9d7DJTavOUjbofIFV2u24siriQ52JYCXyn2D1UOsw1blb5xQql9H9kTqMY2z8ry
1M9r1633OzT/0SUkeEQb15lOa9JYRy/rM3egLZnKWs+5pjz6IIYc28NCI6SJLmHo
C6POny5eXwts2HTdBv0fnam9U0REY9mElHmkj46p1CBMpsUqCB9Z/+SGB33YO8Vv
8NIRmRQzifMFaJmAJekg39QwZIy9+Nqcqi6oRJOBOs4troMQ7rTvyUwG+CE3KVFS
jB0gimcyi108OeKShLy6E+/QGpBxqi1NHVg1t3kV1mhC70c+YruoF8DukXm8/L9i
5rXh1VRTDPNIJyea1cgHC8pQqfjSRUe/U6Ptpofz4+rHLZmspbWspIIHv/V+40MM
5QqbsF01qyAWrdF/cLSYZYRdQtIRiejZ678JJhob9l+uLMO8XJ99m+bQjVclTt1p
5BqtfdvnREPMxAFTvXYM5cNRqzt5Qe1zn2tKSfwnn3R4kwF0xKue0KfL2cVRAjwt
hugyCZHkvFOX2XGLpPdRDy0qHeUOhlhdMLNI6rd+amtyAJoA7XJYCOOWnS9V9HfZ
vRrdMzaH9UIMa6qeX9+LBG4plraQVC4jpxwksqMRPjfyqr2yEaQL7JwiWV2Dm5m8
IrDmOTIGRC19eF8SUoC4rt5OSEElJxvBXHGHE/rpbhzF23NWzZdSECSlR7uY1yAK
ygCW3I47XOinZCtZSrGtzBeNbbLu7t1gTDF8ZQ1JxNYVyWE4T+AJr+L8e5vyrtJA
qaRV2UU5hb/DoQvHrVzpWrEjWAml8La16YoU7JHm8nfSogaN81zjDNpuzclqJpsL
LteJ0jIPrHkr7EX1q9fwpyNLmFkOozSAdeJYIVfA4CqYtFrNzno5fzeHiozhcHle
0vgjAZUsAgho/GlafKSAt3XrPpIH60h3x3epxBainuuzk+nL/AcOXE13L5oGIM7l
6SXPAltznXJKlVdAvZYcZ9NeGzAmKE8usu2w3Gs02GtXDd1dP3XeyjmaGzJd9VUY
GhiPnHOxT2SoAaLSkS1ZuuPHenObTdGeTJFUdLAXma4LbUZ60dF+Sa19ga7SGcMd
CBxwQ3MPbDCiz631KoLlTzY59suWKaIdJ/ofA8c1CV3F+iqsy1ibNP1Q/bnitPVM
lFlDguhBjWnNkrpNmz2sBrugw9NwYwVVwmMjZvclGz3O+FHDnLkZZuw1WwjBkxgG
p9pSm9BBK6yF4FW2CVXT/4PGcPFS7GFdpJy0l00GrUEp9iuw1+a2Sbs2jjdfExbF
SvOornW9WJwvOveOOqrl8Tcszzi+h9V6iLssr0HDt5vekc1Sh22DeAWkwwGKp2S5
5IMLqs0wfOogH4g2eSca/j29pwmt9MhJd0S7FFoC9YZG2CdJt7iArUxy+473KSGb
wFoXZ0yKLGwOuET3PXcY0m3XNsmdFZH/Q2xrbBhREC2rm1+ZGQoD6iYTXDdtI2Nh
n0uahugr1Gks8X/gkbIbwRgYPMNN/cxdxayQeNdH3Z1eB2vMt3txQWezmWnUmeWp
ftQJ5aR0Q8RLann+ZqYFpQmiPaywqDrx2XL/VP5ubNKUi1M7Up27gE6F8j2uVMIh
qO5gkzCbxBMZH1dLCLJ1E5tisn0EpAYHFUXlDs+ya7ZhbdPafgrz+ePIYohNUcwS
LirE6jjb3PAHvaHd4kAfRSYxPp+bw8dH44qkFLygUMYEGv3gIG0HyHlvqHJKy1vN
D/FGyKoFLzzSy8VWkvb3qmKWD1UjMuqTrZGKe5SITQzQAn/g6H8L0up6F16MjiKy
AeukimPGFrP8wwQV19qY0/6IbKDUcqF3BPCGqCtomaLADTlgOvAiwUtL7mJ8yYt6
tPU5gSmg59taehDf8e+btnsUKTCW/RDEsL4KcATkO/gKG+KflcgM9dg9VfC4sPjP
ObgzUpqrPaUPjFeWTn3lF8DS/LOHAJDFe8f5meCfrZ/epampR8YQ+Onzu/9y4fak
0bAGxcsywLAVMOreQPzx7Hlz2NIAhlp+XYI5HR5oLqfMSIdqqg7o+FX8TJU7rwJR
pl6uQwzcRfsvZy75PjSQajM7OeL/bpKpO2NKx32zV7Y1S6zkDamDIqCZLlJz4Z7f
0onXd0OoKvZtAiL9WM1uyVvcD1bIFYb0sq0UPv61KvsMfd8Ve3C7o9rHg5177XH4
zyN9wWoXRdtFqIivfo3U/mZnNTi+/+i90+fyHmPgWWACpSvO+yzhW24yNXpogW9A
Fi8sbv4n1NXmFd+SWDKQ91AGjpuG+IT06Fl55kclla4AcQij73EX7/60VKG0aCMF
qyboBxn1SrdfM3v67ucR2T4MYgYFE0rmzDrNuYhtlZ5LwRaxREpt8tklTlgvuJVh
en123Wtl/Vf7PNRCiD9NUS+d8IihJrGLu4aLpIYi541oTsZwN8cBPPzph3x29saU
2dk5dGUk+xsZwklQtTvqXEd7cQuMFvxJZrxdK6M3QtOzQQ7q4ilUnKaKsg47dHv+
ytCoEBJtXs279e8fcB1MsDUSA8U3DYM5jL2cATGPmMjwxRkjyrWOWiIpvrPeKrh1
NuIwsJFqlAq0CQQI55ZoISMLiyRLL2WvXoan7rS+DxAw1lqGY1NM6aLbuvo8j9Nd
W9eklb7xLqVIFV+5sC0ndbsz0R8f5p0OnWKZJMZqmQP8iG03Ip1zQBzqZDDQA9jO
PE5QQx3XUokuO+FJ+xaWsfs7lG4TFgTdJA+lXNBLSmCH3LQ7q3/Tp2HSvSKdgf9S
yzatfn/MN8+yd+OVjNAPB9tSNhBpN2ZoZXC8sSYWKH/g+ZXSyvLP/gQpgwcUldH5
8tLzbVGj0jUjQ0xP0kLn88DTND4usXI5FRnK5QBc6ysrdXssRbzIq2W1lwbsLjWs
eHSDB8tdOP9oixw+nxyD1h4kcyRtxPLQfBTQQgT4dVFWvYXcq+Put2l5jKkppkGB
jvcaRKO1lcdvQ8sC+8IVrSSLVpgT22rjQbDqt1W1EnIAF5aH22f37j1pAxB6qK5T
Bpem9v53+l/zL4zY06o4esOWSAEhP8llYQjk8x6xvUKGxYj4pQJRswm0dGvbmAuv
n8OsB1uu81NqTIj/zmpVLVY7yun3l4KDQ1GLy/x3rO8/+it8iArCSPtxs0OND4Kx
UBOPjQzZOPRJCE9pXQPRY52M4daFpjwL8EyWC0MvWYSWQvUxutiYBSna5s4TRTqK
V8C+6fjAAaB1+wqt5pYMQzIif2ZayFP/wza3CqQ7Cb40jWB1xZM+AKij7wz+O6iT
77rXrjiosvRCyibIDlnojrHhZ+tDkMZ5TKEEHtvWCXnU/FSYqn1t9G9+h/YdaTdG
KO/VJK6IF1PFeeMYppjylCkbhFOqfKQmPx9SaS588pOvX51BguvWi8stIWPY57MW
0t/6+1AdtZa6vLX35rv1vSm1H/rmC3epKzw55OPCsZ5k7lOUYvs7d9vq6iY+NLH6
zjcJcS9fBci0bPeXDUs5NZHEhr5jNaJEWR8YFNi4w61oq4QDHF3ZlfmUxWpwCVdQ
x+wNsru1gzPnsD8HEYadUQeUWp+PaWpwZEfHIUfKta0ixkhEPSXFpS0u/wY8Mhbe
Rq54cbKb+T0Uz5Hfd4JpBoJ4IAln9/G/RP63J6qS2v+9cDfnIJNDCM0nWiZtSYsT
V9QRr5YvBamiUiHJW/TpGmE2Mfh+oPEHK0lfF6wem6rlprkLjlVSt/cqHzSa9KxK
uwsHKzLx1zAXJbO0es8HSvniQfbyRtxgzQgfX73HIC1NwjH1qPZtGB7CzdOtV2o5
gffYWsBvxqRjQFzWSwrQMCiWraxLj5+rHavvw4936XIfuR2mZSJGc+iMyKWyfdf+
glxI0MrfncySl4G2XnADVlkwJAz73R2M4eADPe6nN1BYETZGGuCjQRggGcADCyBN
NC5kFFXrgFQMcHR/PbnASec0vjlIpzRiYT2EevQXNg+ScztzjsubtdrSPz+oCG4w
ABVcHqHU19i/gItC/0kOdoVeZjDIA91Vf448W+F+VgpmeqsnvUqYyboHJyD+uyhS
DOGNN4QF/usC5QxHKkzsd0vqlm7JaH/YWs3Sgg1Kk4sG5t69hY9ovbZRISwFWiOD
h1M54ACePYkTxupa6irajJsXmu3+AH+rv3rW1AiPf9VAtJslXgbR4CdOE8K5Uzg7
pzMkITA2h7b5TlOb+222gdHiFiMtNn8qeYOrWygDrAkX0zVt6kJPyvgIMYI2sHAy
OUj5q3nqmVDyDejDfTrTKEGVKDNGpGHpMxxJbkWgnH9Y9HKWj4C/u3q8Gydfn/dj
w4cRGJYK9VfLsipMBT6dRtj7YdC25lIXaD9O/+hmilH3GPCMNOoFztMAqdWV+bdD
Eqzc9Rgm6MLazdysrIwaZvkuoMiAyhiohdtOlpd/0IK8GNC5vhpvGeL8D8vy6YhA
4WtcfT/vHks5v4v+wEHS0+ayYGuaEalbj4RWNy45VZWWUJDdyhUkMnUOXfg7Pnhn
QxGARyRWWCahiq/N7xN8a19vLQzYF9lvA/Ufvt+IPZIQL+Xw7roxZv9KrOJaIn6/
jLpUw0ma0pjn5AfNOTXQbaxGFwPHSf1+xipR1lhi/njzYPvPSd2FhV63Pm1CONSX
TJhFBqqvdvu0R4O4wrgOa/U/xBT0nHxidNoW85xtPWDv+cLBaCi0Xt2FnhZ1G3Wh
Sbv1f6WQaxXlyc7OI80oRfaiONKvg3WqxSF+tw1XPqCmI3c10YYRPzI4QKl9o4Hw
7jLl+sN2G6kuMxKlhZT5a5VVN1jEGLEVK8XrpQ8p59BI4gbURvm1OdNZyktOV5l0
hVG2x0fzdWZ0czmCY5/IQ89ye6lNBLCnopS2MFC8lPXDK/0wRx1dbEjKQlD1B+pQ
Vc55iu4L5lXQtf6z/GjFYW8+xp+Aq6j4Mo7QKHPU5FnA4axJiOAVWhAbo85jdzye
Q5ROCmWlvThr6WrBsnYZZnS7GUzaVWLwhvjEhkPUDLfbC+ArVOkhNsRuaYtq+wkz
t2m1yfaf35h3P2HWQxMyhUNjsCwAJrAX97M5v9MVizXXVuMxdj6Y/zUmm/NqWEXn
a0z244EF4MbYUPLlWmPU38FLONjrxLoB4Yx1C+xW2Fz3QRch2keyduggOLxGByRY
Hez0le6+HSSGlm31zPsnrHYM4w4cXQdSSWHwLc9rWoi8PqVY3ICEODrr/A8i2IAa
bC6GYRAw0q4YQ0buAaiecCyWgqaN4v0BuvPUjZw2yYPWxFL0MmRbSz4veQUU3OSu
HtfbZ2dZThglKsNwiObK1MmvAbGygc803L6OhEolR9EdkQSp0vJ8pZMcmPQm2agU
qqOOKkdKksh9vA3A/ORIls9AHt6O+nhAdJHi2JwnVuKB/ZCfApTTLvLT3Dzk2Ysc
nswW372pVpXP31uMPIqffmBTXVMW/94XB8AbWEEXu1+LnjTA1iDIAmjdAiF0igQm
AqnM67vh+1zqben+x5WJPOWEGC1ZP0oIg2DH2hZB0waCvRwTArh3r+OW6U5PCkaE
Eqi6nVMn6ucaV/H9yRAN7/KFCf6D0nBPoyRtsrw7WzGu57LpwCiGL4Bq67C8I08l
KRUC8oWQvFpdHlIG0xyx27GBAXXhGop26/gZoNygNw6RYLVQmHQnuNHlmgWkpHrp
FEk4fH794/TfjqTqDYvBWAG6yHhOUFMTO0b5WXqrRGiShdcyYnnuxOlDi1qWIdFw
t2D/Vk/NvnjPp0VaupRXCmavJKXLhVK6WZUPyTbU72sqD2bSBLd0emFxbyDTAvF0
b80nupVDHirtKYvGMEZgI9TKtuB87oNf3+FOkImEO+gEJK2JHSkP+uXVpcKlR28z
JkVkkQ3IrKZRZc8S51HBDbuZVyXxkaBvuxlVYkpO4d4DUKF57KmV8okP60GU67D1
f5NpuwCMm+SsteA5w7aiFJSKA/9E+mBYyllTwQWTg4LYkWf5E9L0DnEviqJa59Fc
whEmt52/Y4BXcrbWsunK0FZsx9bNFAXve3GNVPs4gI6TCWrnQYg0tfRfQNX8htPb
TtRh9nLv0AGfcXrgg64PYgU8AXt0nnGDeJiyUeRS/gscnynsGatpGoEEA3fa6+QG
4omWYfDsCbZH/GLCiSMW0ZpwjYtvhQQyiKa9cQJ9axwvYdbZ2oNwJAYf+QwC0aX2
9RVapabui4JPSy/AUpCJyWcrhRcm+QG98zZqwF0hjKIHnTG1CmCfiFfrLSVR9jM9
nGoI7quZ2qcen9hyPpx6CZvuUToKyEbqrvQGS9C1jFqWeOUvejL5puZdUGlmTyzU
PQFjrCiR9g3G6ZvF+0qAlEinozDuMcjrNvGzi1wGQ6VD7TxINOwJn+PP6U4zjXi2
KVzKabIFADXst+sLS+MuuFzCABgKHbuV85r2G5SaiFM8y7d5l0jxcY1m+veGpCFR
+GwG20xOv5bMgcK1rouTsKYGudG2G+4tdE6mefzcJYtL02PjYV1D4ENhUXpe8xV8
59K2czg5DztB0RtrsmNg3pSFIm2e1sgBQZgh4MZ0PcR55qj+KDhEuq6qQvDmEil3
7GC26IQ0sujV98WBUDziwxteu7QsDhdII8p1qik6PUif7nRYCnHczHq5D9g0H2ea
ZP0Xs5EXrBzA2ypus+i+I5AOKntD0PcoP3mXiRYBT833an5gIATC9O8l78ORmG92
lbuDVcYB8iRXFUIRkHAEK2pgS1ZISBeISyg4zI8bwB+MWV/3XKKegHAObeoYZiOP
V6liyiuAV2l3m03bBX4Nu0NAbfeZBXSHAmyhb5tlnIidtv1Zw1mGGbOV2TKTKCTF
+GENyivZpzvn9wSVdtNtQyzgXAz10WFNIJDx8u6ho+vPlZ+5E7ole1OdH7Kw4c1R
Dfkp2RuIqlXg7p3mGMf+Tkx3W1dXvRRpyyq8xat7CU/t1ShkiJF1qqlI/BbaBk0F
/eqy+JSPuAeT91iyWypOuWkcs6u+fZLo/ZbCeEjqdUIoLlFduZd35a33zImmCP1F
7z0EuP0YLsR175Sc7q0rFCRJsP1leGrufBLzHypCuTdF20AgbiSY5kbthhWR81iK
D+U9mRzVhtaqYi5A08Pl5D0fdZYeWLrK4sJGiaJSR4RWAAZbAQQKGX+KBprlZvq0
j0AoPuevlWnmr/H9CaFSgN2lkWd5vmETz5KjsNbCwY7otXdxDWHAaVJ8UmUr+0sN
ToJKRlzE451uVX0U60j5iU4Nc+KG+FDasb2yHY0Zrnz4iRfld1df77q5FIApRho1
ggS8VbwDdtw8y00wIgvBjkIuwe4l/aqv/EbNYPeo1FAYa45xMKsUXnMHXF5g1Cp4
dKDQu1UWz98No8NU6+SZGJaalgF22aQZeO0Q69OVMkaLWAriK7m/oh6WiPDkUhuE
5CRppwE/GiGtfgmbyyqu4uTgDTPjKEFwDT5JndvS2SDzKyJ6Y9HDA+cCY68dp9Yg
w7vDQ3JgsDl/V+gq8u3EPBjKbAyFBca7YmEBQZ8w925AlYx+9oSAJ32tqlep26/+
/88cOTvpM0MWdp+ATwx5LpRCX5YaGV99S3RyQ0N3P0Jlfon7hu+uGym8kAvOGZbU
D2Fdyscb/9klpAwR8MYpkpy5oJn7E61SHZ1c/RhhmxabeDO4BjO+8lNqaqoZ30v+
UZLy85q11zQbWP3XCuBodk18ZDHowjsYuPwUWPvH6hL2i5vlGFNQiZoHVsMgkKJI
ObX4AwqFmSxK/20nq0TlCYTaC5VbbT5DMONeOy+5BZ0sysDxmEDO559OCNU3HXvt
wDdJCtm9IJ191vVUHbUJeYWLwXH2mlbxUwIKOq1g0dQxKoh+NctqqYNEWQLv8qti
M31GCRWO9I0HEFs9dScThSPF8DSUxVTlvliSF9eLwB9kA63MTXG2s2UZXnz+CGCd
ggENEFjZjwSL2m/VnAfVYaU1SJqmUPJRp1mS0tPxA8bwveq7PeOes3NOhd9fOBnK
iFe4JdjrOUfWJ62sDDh/XJUDEQg1v6sbRsXbyx11hgmaeuV/xdWyIgWRJJDVO5Bc
XQOrbWMTpMZHvaDjQ+e53AitHpGkb3QSdGay3QgG8CAMa7pnv1W0HBXNprGwuegu
PZXhWDq7SzYKk9VjFCONQcu1ZHcLERqnSkn5V3u2SEnViHr11/Ut6Z0yB45H2xLh
BJ6MfLy3jY2smJiaMun0tTlcWEsH7dp7NQ3GfTj2i95V4mfJto8Zl6OkFLFO0F/W
EceW+1nf1Kzhsk6ewmffbTHl/+qvIs71CNDmjCDcBdu2JCc7hcJsRYklFqxubywg
883tD77KcNEQG9nHASnR8ExgVp2EBCPa8Nz6utSXDO2eQ5wTWf7QK44SsKwt+IDG
n2pV2goB+2KVW7ZbGT45nQmPmoQAgtPQXH+rcTTM+XId7qBk6oFMxwf2aJ3vLWsg
+0cwSgshXLy+YG1iMSJ5qKPoxc+wlgb+UARKfCUWbjurshB/61lDpjM/aMYlJUsh
Y0DflgBbvxx07sduNNUtz/2hbdgOXOqitG39/gjyCzMiwQjBSwC55PvcvzMjmVTE
WAUJYG6HXFOIxbgfSSWFZvfcMxSxMiDXcpWkDNgU/TMsq1g60KEa0lgWHJwITR3C
hnouMm4Ltf+BCdP7YMIwy+HznajrNCx3ncD3qx5X9HJT5N60L5lQRIP4CU8k3GXQ
tc3a5ocB71Lmp+/sCteIxi/zWhUcLrv0gtiE3SXk2V4TUapKPg74lo+lXr369yPt
3Pe2BkSBbt6VQPdEIbMaR3rl10Me1ZxkJQsXJzpzPY9VCSaRIQnK6+RNuO7xgohA
1SEPH6liG28y6fKY/lUNCSXjvIPqyEICA3GpmwMFyeWhw+j+ir8wVbkN4AsP+uRU
VQpgJ+4nRQ8JcRblfHNynlvsL5pG6Ls00bpbnJZN0fQBxTNuVqhec/5D+NFnz8uv
2XEkHn3E4IKApgqIrrq5bozSqChpReE3EslU1MKyGxtwDuW+NtUQYWhwLAdGQZdr
BE904RiMZbJe9faSEKX+kbyqlDPIHGOCxzLG3S0Pn0yVCjO/PdV8Gr1NjwekdI2S
7ZR11VBA/AW91dw80WYfLFK3iG0jishRWLkiMkwlGOwItCakZtrRr9zhhcg9vo5C
Z7cXqWRGyERJ9+S+vpx34zapedLLUQQK+2BB7RS0sJZWtg46z+o6dBjLiGGvp599
zLK2SpjLv3e0T6gQCdXFRyf7tJZ+fOzlpmzzLxW7do4TKPaC2jAb8IYSC3xHwapc
xtMFz6BmzAaFBKu5HqRYjMp/NJN8i6BYrUhsWqfAVAcHFGI3Xhp1S4aPdp+Q4uc5
R3SW88GfEcVHKVgLxMV8NlVSvGBaBDe8PGg6JHtGe0tK5gA0VFdCIrXg6Uqqzxos
CR29ndojm7UTtu2plgfObpVZma+dlfwsmJnd7uqvXY17lc1HCGnbgb0pNcgiMYSn
rbhYH1x385KdImaUVqFw0qk+zg90Xy3IvYqMYfE1P9OKfQB3Mgl+XHfCyZPHiezl
VQ1PDZqj/9s4A4FtvQfLT/W9H50y686l/7UhdWOJj4jIfjT/22O1saWZpE8wvomV
tVshnsgOaVQYQ26dd4SEDLLmSuigO0JuNOjuZiwvgivjDgvOy6VlIz+SSDd52XJW
gidiLUdVGtegbcQh0BPeNh4FzMb/VmzAFM6N/v69KJyFB5HXTiOGvNG96f0zEuGD
m/gnppaV6exOWxfmzSQfi2tRXxnMXlO3vECLkimdcfqSmZXzuvsZfnDDmYPSdAah
l0V7jQYnfuBksErr8+TceCgi0uPkljWMbk++g1vuxF8jVrUUGQY0fa2sd2fxxJ0S
LkL11YDQyKn7E6Z1kyFc7gt6fKH4Ni9ASp/+8+On37RS0w4uStjR2ei/yDSj5XX7
ymcts5cjlSFO0ytXucle+LH8Ggm8A9PI2cE0bNsvt8vdd94OTfiWUjaEg1rwRt1n
bH5fb8hvnZEeCvvmteLUC6jlJENFpgtdX15eH/xB2W9PPFBOqVOAhlk5i2PQPZqe
Hk/9V8iMRp7RWUvdUMoJBsW185FHUIjtlciMEGX+I7jylV511iPJ9k8bVLrwwXZh
mcDYA8D/UD1JIIeslyhnVoiotq7whA6Dg7QM+8KmbK0FGWdEMMGyggmt7wWrENOR
KTma+H82GMwKTcOr4RWvlKpuo1E6IU3z+tDjSs2NtLBkIOGJ+z+UPxmjyaR8Q5qF
AvXosycbg/fVeFMx+tYEVWxdrbSFdCEpZM4ZQjpitb6Oors7tzktXphQ6mUvWcA5
wIdDrZdCmSuI2F73Dt/x3VPVLhLBpOGCC+OxIzsh4SvgQsp3QZwLu4UGzayQ38qh
OkDyzBtt7Keajg/riwkVTM5Tqxv8F0h6T8Dsl/JGwOywkSZh38LHV91qKPcH1bjT
/3oJh/s6+voNt0KdHRJ+aLSNRHFrCnr/InvkBKsf2xQ6t8a9XbQloZ1jdPO7j4PA
FHJh1iTAKdOzviXQMIeDPdz+BV9aCtedrXSjZCe/6QbG1ABpNocewiqbAkLa2Ty7
31/N0IV7ylhsIYsiOZB54cZvls+fY0vbj/vyLBQpbdmrvbka1pOzGaAhhKuMDVxl
wAGEFhEW1vVCOrHPlimZqqaG6M7K04fhyhq+ttI+ZQ5NXlF60L41i6nHB2tJGozd
2Nei0Jdd+xEKbTdM3cArut2C6NTvIR65x3/rJZY6wiWhCRMfMfv/8/c4S/kL8Q2T
2JnFM6t5li5SK9tT8be2F4URPhoyow2RDtsY566VbyOQv4ayPAW4fFmEsYSKJSJ+
S0U9NKJUqiRateGE7X/XVxI8MnVzXdlTlWMm3PX3uUbecIg4QLlp5ZN7Ph9ZqJGL
SSpI/Y22vTdobmopDYFDFGz0mtN0/IBL0UdCQFpTJ8gtlLeIsH9eh13GQnJhMBit
IVII+ZwBmbyaROrhmooF5OmIUmlau8YM0iSfWJdsRMKNabmFsnL8Mrytpo1fggyK
jgqHD4t88yEXhrEd+DvOYtj0HvOB7z7PRYX9beBGmrG/28J6n9pQraadht98zfF/
eXzCQVMGPkYKG3UrC9BgScjBbX+ck5jxx2TvedBrq0b1nIgokG7k47KEKkmfSc/N
vSf6Fyl4ZO9DqXxXtnBugQLf01X/Fs6Q6uGtnczZCbhzwtTAD3cjgsvcFBYBeG2o
ol01xUtAi1QykJGOlYrOOakTHzERvxr1d2UqLSQorfE0NhCgVCXJd7GOkvSE1/Wv
/mIaGunllC+e59nStRH+1VPUk63yEpveqsS4YBWmkJ2tZy7cuRfOwgAofzsC6jBt
kKUoac0S8EWZlyHE3NJcWxOCrsWuz+Z6dE0Vor/dv1DImob20b6EDEMz7QOXtqY1
NTb+zZUk0jGYSxO5QZSbgfhEoxDv/piPW84Hm6Z6ZrL0eKuJgUPnWjgtWhqajkoZ
4xSrw2tGCKmbanCUkvIFrS3BW707ztl2f9vivUP29qtis1FcgC4jdYMvBNNp57GP
s0mE7+WL7hMGCmBHnqoh+ixORb5sbphKySW8oOCINeWdew5EnKBO7EAuIXyDFSxV
yWtDGdymgGqvJOkxVmXVCJ+EQlgVS16IVvlElQtkIvU0+oiIgaYdluuAeD6v4xz9
x2jCGfDD62KGBLqRyHZKOSiQ7NHJ8C+aBw5W8Jro3bSwQjcGjiSsFEez9CQbkeJ7
ePK4DbojM1NN4BzlXnjgFVdAOCoIWnrPEbS1y1+iMJsrcTu5+eZV/0OmbpcqFMQG
fuubr3nPdIf6+Oahzqe33mweZVs39G68nhpj59TexADPCDB62Ppp22Bh4C4fObsw
QdfTkvKfoaVZFe+3NsVqZi2q4K3nk9yDQN4iZWaMOkmeP/tfS0Cy84EVsn93KiFg
Sqgw8EPDoqlLGwDh8NPb5bux5RK8WhnAVTzN7YqAT+eXi4XGJp0bfB3TXGoCx55i
LLBdGaWfZ8mD9VuKiy57Bsm5q7naNqv34NFB1Z/Kw0tIZw1uVCQliLdGH59Ilykm
9djKv5qQO3w6KM0OB/fVDweqyQg3nxXG++t/NAHoB+s2BmGUBEcy63bG3zKLXWxv
wJntnHpHzJd/0Lv7YSTZLeyJGVOhKquLIx9UIIS7KYO+8/NhlAL/z3yS5yY7/cPJ
8etYiPpoAT8oj0/3v087GZvQ16rt2T6I/uAUmQ+sjmVsZB8TqgcezbndLjByGi3y
f2gzJUvvquQC9Wi2vz2rCUsygmfzV2KA7/7w8nY3Y8HXUeQfUHnnomHPB+kW1EEk
domNshUw/QQS2IBv7G4kiMEw5OEhB+55dd0awRj1+m8COnX4e2BebKjdqvj27xzO
CeTD2x16ediDk6inrbNcEWWyKkca+Vrvdr6qPo6y6tmYcvfYqqoJJXWUdA91Snvi
u3WBED/l8sAk9JTa3qLeQCvkb+LHrCOdK3IG+ke9dsN7tDsalknNBy9p32gH2Hp2
mPK+AlKUKifdW56PFOLNmH1pn0TbHOrDjb/ZMryq8/+HGbkxIJgb7AqlOxHnObmJ
uZ7XgEBJ7WmskpopFL7xDaQnPcw2oE2XgNcml5lEIMFKei3VKlk8xgxTUxQjPcJA
cop0M0W6s8uX2YcefNnuaggp/mzn1wgKjWEfwXu9sbil0mqgpsfuL1fRZ7CcPSJ5
xpVil46PxWyI14x/xCSRcXFRO4Z2ZbqWhIdcE2R5NTVIoQPYOEDNjF1c6SFziUL9
kfnRCTXvXilwX6bB7LOXsrTu3ooPtlbEbFgtDibTt2BbHiJ6bcJXFP1oktQXRYVx
Qf/kNpJIDVblsWV0NwyFT0qQCvliVy9CrQTIxmF7a2idhoRG6YtVtnoBta7f08pA
rCPFgw8xN7ptM9fXWeCJ9kMIZiZHMo7ugvTMKGlRTzAAcPrdzEQXL0pylDQc1pwX
a5i3ZG3IcgYXG4XHCfDi0PKButQp6bCJAeJKtiN8NLKeq4Q03zZFDm0Znufv0J3t
1Gn3McUrvCF8gpvDjH8ngxkhE/7hP3/aN88h1NM0LRc94s+vb2wtRVvSQLvmVsam
wc57K1wnxNchRrvwDRo9veZdnyxaQ0ihiMVw02geoY67SrITK62EtXSW1Act/MFk
V1tiQ4XqwuwcZ93b5gzSu6FhrsMy5AHOTvorZ7YpeyLS7LMRVBGO8OjYjOM6HwOg
ZwKDFMvEfilBA/ofWYtB5Lg5Aihq37TUQNIiuSEP7ALldS79cc23oh7IqA+bDQxJ
41Ytepi9I2YI6pJAXPxx2+8shraomV9KCR+yAsy6CKyJewXWYyoK+YKB7US3CdV+
PpzN9EaYois0J9L0xC6dp3kC0kPpn9iogF2+VK5I6DnKyrD90oDsp0h6Lot7Azvd
xB1zni1f2tcbkmX6tmAdafPJMDgTB4Kbv7DXlv7NLZiVdjZ/ccKIy9XpdNhpNiDg
ZvIMdYmi5iKpipFeuPWM4Qr1ztN+j2U/TCP+NfvltYw9a0icapMmm/jcQ6c1Tw5V
235Dmeb20PlS2Mp4venTG+ONBSiiHEOi64wqz7qq2emhwpnEoYgPAcipkgOCnlil
HPOOw6vLt33ra264OTsupGuMZSNm/G4J2naivaJLaJ+YnMSmlxKLqEFLOgJqxavk
eQtlO0uIOodE07hqD2l5qor9bgBE+Fg9JcxAhDuiVa8CmKCvkVcV2OJ9V4fzwu4B
7HWYljIqupHCieYDjINJdF1SBuzqFZdb9r0Y3w+KyZreDoKexPgFnGchdkgn4wWt
3RSCao+WoZHqmdyFYWWlNHyixcX5mF++IA5BN/5R53E+ZwBfDxiajdkfOYWqnr0T
BSqEa2lME65P+rMQkt8Tvp8How9FXXiN2ghxZlFnUMxayfOEUq8gPgaH+Z8wge5i
d1/ldXUSRSQKMWgLI+yvu+zr+6IBp0YE6Qw+BZ97UtQ+DcbgDnHNhLJwFpLmoZGp
I3EFC3+2VaBwbPDWBDoiXPwMbGiArT3sULdBEEdjV6SdrAdtQE1HkufqZmcl7Zy4
Dz+Qiv9bJjtpYVTLNiTodQ0rybMm9iCGNBwGPT5qQeUCrNWi58RIFv5Qcu7KWR4S
FruXY9ijHDTaIf3IbIvfP01pysmUrPb9+t/7pRIeXD1AWyHpQOx9nPp5kVprX9d/
iJYEfrxiG2cL5qJ0yTteuPFTMxNIj9cXL5SW1FOV6lhtebWONVdIkNOuq7PUCE6X
R6ttbWFDGvMMIR49pDCTd3VX2Z/fFq+fC/djddm35Faa5E6SXfh6fnqaln16JPVR
ex02Ee6pv2Ml0sO4wG+mG/MqZ2aTFQsm2PyeWw3R/j9D2B0ZyZCadp18k/F4Bp4k
CILXHUJ6BP/Lj94zgW42qevH4Mse6c4zDgSiOn28fItUpQQBLj/Q7w6E4077GZfF
KYmPtrEUV6jhotkoUFToNo2HYWMVjxJnB0tg3Fwyjrr47MQKSSxWT3vG+WtksO5u
3MIt3mH1NVdcp/iqVYfBM+dmMGB2+qoLK7QozNNpoFzVscjhwGJ5QsUzMOaJat3I
JIhA6przOVRDml3BhZ2QC4y12dHB0Zh03wunU1QrYgsh/2FeqMpPBlT/U9mEi5Ui
FOFxEkxj7Q7lE5Vf6AzbzyexIXk02Vp1jXGF+0xCjftVy4C5X+I5Do8iwBujN/Go
zhT5sy46gvUTQKe3u+/nI7mjEQP8lcdD0eC2nn6P9cSL5IR/43Gf2EVx5DPLB5YN
j1+gWj38p3tf+bZNKZCm/QgFlKKl9u9IfQ4f3wsJJKlP28z5XX+gTXLO94dwIQMa
XkqXPuxPJgDaTGQQDUK7WQYXB3oAywLip3/zR7VHsVlI2gmgAln8F2AouJN8b89K
ABWv4TQ6PhPTlAiztqrRP1MADDZk2v1PEVq0azDYmIP6IJKgvXlUtZv2WQLcfWXb
8LySr+ad3ql5Gjf21U56uPY/gCRBjtJtn0i0hMz9K/XVsoVGC7GZ8FyoHy9/L5Be
yOmRWuIRt9zJNtlWlb9jX5MdDGQ1k4RVRoB4ygYHMyjHxzgx6GRlofWeWW5cA0PC
ngnKoVkLv19WFS7l9qj1nvjb+BWXZEyKbvLvvkL8GLulX02BIcpqJsTSHEjCEayi
BD/UDfAxH1Eu9BDpYyE7Y853sIwVqBlgb28t+VErph82dNPhipu33G73Av8bvGYi
XV8azzksjhL3HUIiaT3oOTXMgVbb+PgDEP4HekAVSRXhSPkhxHy+h7DPm/4JeCjG
IU7NsnTQmUfUI6QgF7nUb6Tg1lrXlb1x/lC99/fFBmSYPHxo3iDvAnMG3MGa9dgG
nfyRibDp/iZ1SA+7Mxwl0NKuf5BB8zzOUsKf3j4IhE954eW7rEwEeGwxof5BoZXE
KyN7lkf80G7z10MUCmxKF2jDvqLGTJtyFQBPSKQaikmk7TncLMtGxONVGj10Ek0M
kUFA81DF7nQfU2uk7u8tPav4jNcHMycJUFz1asMT5VfsqGi2kdo7UpakT7JGT2GB
XBeip0TBS3QPuuJ/fdPJlHtzuvhTkMY1zHdcGmSwuhAYL2rwh5GjrQr2pKjFbgBq
g4pkgYHO3GDmzD0haTS0ebzKGSdUMWMggQe7h4UKQS+N5dZEVpagq3w1/WyKjbAC
S7Sgu06N4TcTXSunyeqX9i+vD0EHWXHWauC8TWMOp/Z9v1guW1s2+Bs2Y8E8nroT
OSfNNKk1P0bh5evzJumxwSuKRyrbG35lNbBnEmQFDqpfwbOAjvS5xLWeOnNngeHg
X2EUQeLe6DD3CdCF2K7lWvjk8VV/HXj+Fg9GNZsVaokOMIKJNPLPBdjq4dlhZ/BN
DyYQWUqCvanJ6St5xYoXuiVV9Mv74Eg+MjFt9diI4ZrSfVldVPpp5WkJace3AEtN
N1TJuAkcAwT8Wxnz2NiSZ3GORfSXw/WGQilTD8+ODFEB6IITuxuBQONskKE7G5Xf
nC8Hqyyqnvwnz6p1T2hra09HzwarnPqLcZwGWDkXSJFgAfEEhx1uM7RGpwldEcyR
XhCm+181Rpq1D2k/wiImAvGWp9BKhsx+5TqmJshIBWf01ZJtiAKoodfc3FJ+S3uX
3fku0Vbr0RqC7fg5oNoK1SuT33xMOhq9yG9/c6QcxLeOytAAguNLE8Pio5UCwJDi
GqX8M/d9Iuo11J/XZSBffr64iPkQqgW8lstcvQNMtG4GuIg3dcMvog12p2M2vxOD
keNnKF1XvOiNRnIrYBM31/r6oVjRgfxKMLMVCVzGcf9EuuGJn9XV2hgzJ/QzQoWq
GiXBJaoZO40lw7rxa3V2JYfm2rdbM61c95FU9jUUGdeR4YsQIkWbmkYU6vzY0CSe
vfVo2SaGt9ZFRvoARQksMt4/902rGeu8/VbUsvP6Lw+8D7+pG0hilDeHjkaPUiJt
3FsIoa98R1SV/kjWgUC5aZ6tnzhE9/qEV7xcO3oVlbUDkoqt36osNT8bdPpCU0VT
hH6hdwgz8Cmlo8Xz24XMRAxeIr4jDwR0YD8H6iSZeFDVEL+Pyy/s03gaH5LZKivv
wZvGAHYqOJqqOtA8+2gnY+1XjLwqziKjymEGUr/p9x8qsfhF4DaJ9x2VIZddfoqV
MlJs3CAPJx3Uz1HHpZzHAe8wq49MFiEoRIM4bOu2iXtUKQUK/tB3Is0souNB92FG
HnWmaKFbgQHk+ylRqG6A8FWgGncAjTPETKApcv+AE3M3ozN/wtmk6eb1X/Roda3a
MYMDjdjEDQaxXq96oTvqycTwYEW76w2tEQbRA1/X1+rJxp9xOGS8CVPVLUv9tobT
gHlqJSzXUhk5XEgUmS4inOFTy2qimYFF6fB+R9eC0Zjbytc18tLNQSYMoJ/S1ODX
jtpRDfr69HEmEKymiRVEc/TaLzXvG1kexQvw8vDn2xiAQQ+w48L2ezWQIoaXg0q1
RjjTg7ZMZQz1wgdqXWKKelx3CHilCy+8ZKG3jIqQgc2zEbfoOEOgoyXhAYX7Mmzj
JIFwX7iybgmfujUYb2iTiVUNrsvbRSmFlnOHrVcXFi15AyahxH2+WVDytUZMNMfF
zYD4GBpda6oC9auiXo1Gqm5lP/w2maus/tb2QdYwPkSAkNPh07q4gzfyyekgvWbx
NbdwV4XXZ9UB5gAyPjB/9uI7B0lJNyPaBhVtKSvPuH1ofx97+/wqJ+QQSMz/k0pk
jJqd/cjnf4Kenw5vbUiW1YEMXt1aEaAatXvSDwgMZqXiGFEIWHDha3djV6coNLj6
dqm1PfhZ5SQi3JFZm6vDDz5qmVbgn7GbDycQ68ujZSgtKBCRVoe1miPx4nEM1Puk
1Xewya6qyG5um+FFpvyKEsHGX//tUBQsloqqUodY3GWxj/QgXjMWwV3gkgv+0q61
USXGhsMRwdlkRwG1rTGZyStuHDb26P/Opg9I2taDCQA0RQ5Dy1QmtHsTrs4YacgE
3YWpA0doLDoigWJaSfvlhMtTmLl5BZLW0fSvtkHd/jaZNSk8n/ahc9JTpF6IXXdm
OFeBbFzZY915Y2MmpGOB8yIlxaWo0SoOuzwn3E5Jv/+ZyNJEh6VvrPNCCLrSbOxe
UnO+retzr4LR/PIgm5J6KxOFrT660AxNaLgR92PBELjnn7l54zd5WJrzMOD6fe/U
GvnHhQOfM5Mt53lQkFnu0n4QUWeG/1J6NnF0dM/8eYkBD2J5HN3knHQYc50V367w
NgpZXuvby76TfkK9cWlN5QV4vj0E+TLKHqqcfZYXTZjVrrlBm9sZVB99FDyXcbSq
Y4Qkn4+6pWxA0pKBIX7d3fwrZgkcyacgb9OqnhhJiTT9HAefCp5NkP7oM0x/e/NO
El3RY3Lf7FtfGwMJ/fysz6rsMh221VqJSePHbCGUXVqoq6tOoqTlHkD0m3sc3R+O
DVptLu65QE/LjQ0sYXPw9XlIH6rlSEWAXUCZrtLwM2ja2Nt0SR3tnvaLr+UQeUny
jQ7DzKfCSao7kRPs/4qruzF4UJuZRAPZYRQueA+Tk5XnzbH5yHb6Q5ClJgAknbBC
kcz+F1medXRKW0FcSw3D0q68buOEQYUE6d9REpMgJSJ8ISWbr21YAqpxiMnwO0gK
EvLHMR+qXU4LsfBGkKLEjpa+OMxZ200SdotC056C+hB8YqkNbx8ydYYeq6PN3kYS
vY+oh0cmed3LTskKkWVUB2/gR/SFwowQcoL0cB67o2be+DgLoEdkf5I5WBBMsmqq
ovZl+EGZeDf6qleDmP3776Rh9m7B4DuOud4JUQmY2aDqaf1Veq6DLL3seml4Uo6i
XXTVpiFHving8Iild4Gw8HxJ8/knsBnGhyxlx0OxdDs944vkCtqm05PuYKRFNYw7
TYApMkd7FylKByu8JxTJtDWjLEoBDdB4DU2mDKOGJVpiLMLjzXBi8kT546rOVx1K
E+mlWkxwcJdMEo5iToN7V7BEVMfbKwlIl5iPmebfMr/ExM0fQlz1sJOpo7t1+7He
wvAegZYHIHfw1CDiA6bnC8sa8IUCv21d8X9FC3kcloJ3OlXyYPDKwpLezb3b211r
xfKgvAYIsMeGpS133U+hIjawITmRV/mKWGkJ4zuDxZ8SskrgO2GghIluqz+XkRUE
TxKfK54Rs3ZlOTTU8VoIBlgrzwpOxVE5vLIsIZWmi6lAUH2UGaYEXHmYBbH8dkw9
aHSiR2RAl0mMewR7QkaEZ8WbjawakkTddagXIIA6JxPArW8Jq0FRXad0XlsGPy1q
tKUO3tjpYZEvS+KEJ9cbkZ+ovotoG11X/VqNbBLAu7ad7r3IUc8FkTqypyNaRrNN
1IVVVZjtnI1eiX6Nxye/7b/yAoOV5Yqwe3aqVa4Q3EVRrNxSOY3vRtetjeqWD4V7
5hnwWbSaaLcaIKRBITujLxyUcQLvwmBPGqrrZ19ETDdi6Jwu4Fj9O0iR9OARAHbG
LuwHHcAUxa8iynh2UlTbTHflQrDOfsstxlL6NQNAH9tB2ri2U+VBhQBxdGFgIsAp
9Zkk8UIkTQvccv+fHQrwiJH+jKOKR99u1S9OTTnBfyA1yQ3AXGzEy7KmEDObRay1
LMGkofkw1LwanmNxF/nmOlmxQiaHgEa7dv1V3Qq5GT/QFGEU7bCaP8/45IjNrJjs
gmBFMCf6YNLuaGwvo8NjaEQ31EH+xtFVXpdujJHV+16n4ORW/KP789R+/7tS4qhG
VDiohe8CP7WhVdMHDMUR3PySZ6C+lc0VW3uXD0KFQXvfaiVq9Ur8XlEWX1PXi378
MV1vGcqRmEMpTHATi/qlu+p2BV17JSJXYGCloWeo0G5SKvz+k4La50kG5anB9EI/
uFSeI7Uoo6KtZnZdc2+tjDUwGUCFikU6z5hyE0EidvxyQHVDAjNL5imVIisK6WNn
7fmQ9MeoRihe2UdqyXN5k6Pa1kVZhZPwstbfeIcAPBtjOXIQ8ruX2BGsAh6CixVE
HFiQn6OsqCrjQopZ3qRglUT+XUIdlgkyeOy1EA8N2zbDBBnNOj858dUWE4JiUHry
PtQap8YRi110sadJkzpoeIKeG1w8hTB2BIufHzaF2Hwg9aeAJlI8nDsFlREzNmES
XpWD4AcXhyWNCLDMSFlwuiYe2FiSbxFtZH4unDpnwfye+gatIQkJuGjmmQLCZaMS
zlzyIN53rgT9lO6qfchQwwAp7pPifdR+fmIWYV9qIF8OsOSU4GhjYQU3exGEUoY8
e1xOrjJtNKGZu2TjGQL3S+/BmWUh2ZmdecgK2TEdlaXS2wF/dANMY/MMFbJZLgGK
tdqViO4bh0ivmveXOv2xSBYC7lmoYXsNOTB1y3IrETgLF3e5pxQwzO805+FV8pws
iK0E4G7/E9EQOiN9jjzyIak/grCsuA/pmBKGuN685WfyDACWf0lLlwrrtnfquJfe
0pc+iv1rXuhmNqZsSD2OiWByQwe935rdvQZ3EfDnMCxeBf0nG6BHQ5oqEPYUod2A
apvr92l3GWjRev1xJgadt26PhJuW/wOyjuRaR50dffDFiAthpQA1cOEDxSpebaSH
4SgxVlj1VwryKVFo+uydvwzh9tIzndWS1mEDC0F1/a9dhsi+ksM5HaNgVF7YazaF
OH62VBp2S5KckR7aTlmNQ0wt6YIGGikhu/ipRntbn3Aj/QjGyegfgM9sC5T/o7+7
AweMkTS59Feelb4yQIGKwdSZjeV9oN7PoFrztcpGomoOCWHlNKIb38z2V5hI6EH5
V5XUZdVig0PLoQmNshj0NV923+2lEurXohIfNMkoMhSLHcEbkWZf1lkaNYdIL+ia
8dez7HwuqES4M5Lr6seAFH3jE+/xb0unZtYfW9jK9KTq5kk3HmAKD+VQOLPeRpMt
UNWjXlBJyHDpZPpTzMDtCjqWODYdKj4kUoUTk2+CnMOyfQhssWm/rsoZc5Ung/6y
qgurNLaudLCp2lBY/IEDwlkczaiG4N9xjIO9JMabT2y9YABhxqxeWgd/8yTcxfm+
TEZnJJSrvdNWuBVLLRsLhRfBX6yi2BcZNgPACHU7iamsjqR4Uwm0ayHmLuzgzJsp
7aaQNlr3CNFZ19GyWMm+FDjfPgwLSZPKH5D1L3SGSeVruKbzITDqMkLO7wZU09Y2
vGiF0Mp8XvgvZjKKiBYSRsMZormqhFp1HqGcVaiWvRIs1JJIPdKJQnGarcJI45rP
iBfFio9CcwRQzpdNxLQA0mFcdl3NOUPBQamw7osEPj8mvPVwuU4pV4Zu25AVyl0b
yKYWrTk9hj9IBztuaevWMuKVsC4teBN3RRTmv86F/0YpcFdbIiYnwksmJZRfgNIy
KHi2Po1qEP5pznV9pU1uSKU4PDiMiFSpkRDMo/hmTs9NMQh3SJX/HbtoDdEk4dhc
ZqBKpyQsmwHD2iB8eml2FAPDMEBEGvXun4lMQJ8lvTKUElDr/O8TnO3lNz4w6Bjf
G7Vd6Xj69U3be068FE3DmrYlXAiTRvQ/l4gBrAPoCAk4lO8D18iK3maJp7J9Slwg
LWPhXvMM0cQBiHZANuilWqxShzweijsG/05bLWfx6rrbAsxUVX8b3En8U7pQxSS3
1+OXLe4yegiCgKEKO6ykLFJJn7Ge0rJPPoNz/6oBKeTgqpPCE2IQ4UR9LUWCco/G
aLSyYib4hO5KikrqXPvdaeBF5C4/6vfMcFnQRvOWcExOjj9e6sem8wSorG4kz8rI
m4M2RPs4QpDJmkbPGFnGKHARQQ7WvKKjdxChQMdWr6MBj54We2X6j72kPj7tNgof
y/xW35p5O69LVNNxFt1fyVq+/aqP4x32rIw3bRbCSN8I7a4OSm6y0JWNMqlQJ3K+
fPIwl1FjVkzI0Tc2YDHOalCU6Bd7K1BGbwJqBVwnsTlkzJMQQOGd0kG8gnmLX9BQ
JlzCrQcwaL2nYSDzST4G5oO1Dcdb2db1nE6YJ/NDLHXt13XVQUPRXCU1CCZh9eOB
CpSOSw/waGAHaVBRWZZTQewSGi32cjmhxzvQcDJG+99wwqYYDy1wf6W8h2xYIYpP
xJl3s+VHjZyLuQEZ8ag4QPob/MOGpumRh1owE7TUG16bHoPYL7ChWy9wbocSHgJY
eGiRdgO4Zwd6vr9GuLIHVNWqpxL3ctz3AUoKU0G1qJG6JvC6Rgk97kHKxEy1sH5k
EsAL/70dinW6Shb5B8SzapvV4lYTnGVWFe6gBjLEiYPjj+6/AS2KLxEUDmTmN6gi
0RYyaWMq39Nxe3VuETe3qUYJGYLyYlg7jsDju5TgKLOGwR0LezUYYP7puGGITgzG
SVmg6rRVzjaxAAujyLUZPvhchAv4jiuRkK5ytTOmOvGri97PyhQtI0vm7T4w2Tjw
gLO+RWblAueXOOPJdIRvnOsNrNgANJij9AECoNwJMbA5+oQRTdYn24Dd8vNadY+Z
386rY9SEyU1pPLbp+HJHAMWGInU7TI7M6pTuJOv+fzeoOJKvbr9wog2spc3ID5ns
hfx4sHSbKYNAzwv5tKMc4qh6RyRjtEt4wXu/ndUwRcoYXXGkSOd5WvwjwgLOsF7y
f5eHjEN+e6aW5KIJzbggrhGgRIISbJokkmqCPHXe6ZkFmdepDcW2Ebrl77TR1p3C
mBMANfAwB/JHBveOcXiq6DYrIavJqrmo0Ev6Rz81vpx3ytPLHB96JtX25VlxuTCF
KC0qN8oqNi8UCOHBseMP9VtF2kZyVGUAZG+jAhvcy4M6Wc9HRUv7m1pQUG8tLXdI
zHF/s8nZDqB8DYlllExcdcg1pXAQQpCZD9FDumLNyMep99oarBbXWM3XWfLcKCGn
pgs6eqst1wcIuqn/gK4sq5rAu5zDNGIm/FuuWHSDTeoCo8IOGweQn6c6kBwnUwOu
XPiu08GR1xPu9qaIbxJhEQQ69iAhF6ou+U8xx81V/BeVfcXePzfl/CqgwcB9aWVP
EXbEArRi9ZbnTmdL/OBWfVs/X/PBeasr1ZngCnDf/MA/xEUii5vQxXlqQwQPHwsA
3fFJGJ0rh85P2eC7I/VOAr63BYg1Z6Q60YeIcntvHhOyvWqqhIfwsJtbQtzspq6H
NWEolqymTULTVxKjJtL1NSg6V6koJB6p3AOOsKFtDun+bD8xfk/vxmd9ZAprQrgJ
N3tHCKLkF1Oi/YDIHdf7BXdJgqI78KU1LhF0uscOdUhq0MXBNoUhAnf8EiL5JBpJ
CkrlnHRxVCa5OQDQR7hqNaNv9ay+KTSWIDmq3QYwqHb/E+UYB8/m557G0QB2zLgP
iMau0No2BtDEVMGWsT1DYqMOIO/D66xsALARNqoyslB3p57aW8lZcBTsxbxbZnI/
mM2M/4EymiN9o94rjjxeJXKYVD3zwQow+uINUHBBnw8T5x2ObclxrvyXFphTR5hB
YFROVtUqWRRy68o626di9AuUBciMuo1pw7CfteQzrkzURy9IKUShxqruTdqTGD8a
5pJN77HPaikbjfelSC1ngOTgNUtpvyt2DfHPAQzXczOVfXzJIn9vVrP4UQUwpnGB
dTmOm/AyJa5ddxdzNy7hHmQAxlB/RcOkjYkxXZ6w/dx6vg9FlIFeet9+eO87FvDl
LfslNmCI1v2EL27kSQjF5lCy/42v7UnOXhENExwXG9xqn0tKHTipaK55wNHCfqiV
361nJKkQc7hxN+cN6WCv+UCUGT15XzFFLWIVT4RSNuVjRsU3RW4YSPzSgZrjP8tC
8DYfXwIAkoD12ZFqH3N42wLUd3pUrsos14fWHE7yo8o1Nz8O0rp9PUZpxfZCcl92
npPccm3GvIuqPk+hDI4e0skbp5a5AsQVhxQoM1MOnlvdNtBZyZrpCM0Z01P9iict
nM0LPfyrwoLO+uB25ogeGCjor6HhOc4yaXfmoOKqzA0f6y1uibrj71HqWAULmMuk
KuQs2axGi9yb+6sYbdd2awSI0YLWAtfKjoeRXS7TwVQymXjckhZhgx8UNpfNg+OH
8+cq3QTi+L1aWdeERVyRxgXaHJQdDtslSlAha/nYzwREAcAS4iMhJqLuBkkNy8Mw
pZIrhOijBdnzvMMOuT2qBH10pGs/0VF+Emo3R+4tdygb6T8/b7SVkSS76p2PLGVA
tclCOewgELIY/nXC01G+NIEkJDxissc3JOnFctNU6Gxpev/7jnf44MnC8zAai1zg
D01IxFSzjZ++Qp8EiqycSHV+sndiaZncWM4Ni4VP0lxrl20/SOJVyNf68qZs83nj
apbvXQM23u5jkdA9gPuvaJzky38R8UXqKrBJXB2yW1WUZ8gr0K+W9Kw3Pf/SxBfl
0HYsKAKakM6WlpZc6BIUaZIWa07H6rMaRdy4QceC7MclMRxhPQvC47HjNN0i1A16
9jBvgj/N1dIfGN3GyciZdkndyJh0vxaO+awexu94xHrjX/hedJmQwCkPh1dq8b5Y
uZqe/kFouh8GdHkP6EvbuOr6VsAp86zjOpubMVtFezyuGOyZAZZN/mf1QxWrDYz1
50wA/rb+yctkYxfDdn1lYPAoXtmgmMMgR6ei7tEyhwAi92B3yzU0bI0wUw8TYIi5
uRWTaVSUQq8QJpqVwxuFJ9So97BtuIKszK56w/u98HB4hZoYZxkLp+bCzZVjjztF
vIpyX8TpqYfAkog3e03zcwwI4Q1THZTYSeoCwqV53vWh/Uj7VgWt/RLkOy3R7ui3
nMwY9ydz/fCM/arxk6FkxbiciDCq++EZ6Ic8kz8gWL+qpNIbUseI2/O2iOHPiFyo
3vzMb89DEsCgnieUmtoHQzqg57hU3VtOrRtCeZtiqYHlY+33kMBN/h7c+i0aYAC+
CcF9viQWNQ2YkX3o64T/oPxYkX7vEgaFeFiZkNaSbmarW59eMAs3+XFqxiKiJU6K
05ZQvRrRppC3UI3MgF5Ap1IV43PG4fdOvrzXQ0b5O4LRVv0FsXnaEIUcMQV+7O96
ApHiMki9Satv8jH71F7BNbif8CourJtIfSHBfwVMdTzgL0tJ5qvASz+u0EWXmQxE
TMfRMsyFwz9JQkPJOqQmRLX8aSq0yx5nPcJB5JLKkml5rqM3jOCaCFvg+jvPvGwR
m217yadQqQNyVLddebFxDdMtCDjP1DdtCj5Q79hTzXGJj8zcyxcXNotrUHDxCSRY
G0OMUizXwz2ucLVypGdv/w==
--pragma protect end_data_block
--pragma protect digest_block
a/4WyQtiF3hPez/QB5cDSJwPMFQ=
--pragma protect end_digest_block
--pragma protect end_protected
