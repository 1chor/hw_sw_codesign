-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
JqO5+mvd9jQ/3O5Ag3exfdz9ckXB5tpxLzF4noZdwxaBAHE0mS4VjIDfq4SllVTx
W4JP7D9cKbo6+RdtgkzAFIXIkfjvM6jptSN/RspP53D9fepODqRG2YGMfEu31bKK
Cjq9r5ZXuD/uN+k8x1Y/QSxx9ixbZILsudwTVf9Uzwg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 14220)

`protect DATA_BLOCK
bg/wF7YMxXtGEU0swYG9gfu3MRpSICURZRpR+z/YN4ru0t3C8OqQ6L42Epmu8Vtf
ltblmEp47LOtkUQxROOiS8njxWFWGYN//nDSzMOZyH+whXMdrXObiuCOjxm7wkMy
QVl7lFiuH1CZfsgMepBxJG7V031c2ENZL9cdEzSYPwJX9uY5bqfxjWXyAulkz7Lb
slw2j3voEm+/+BOHtn5KnT7iPz+Pbgth1DQmF9B/KU5IfDAnJtS1l+gXS5v5boH/
FRW8KcgCWhc/vLNenet7E11rwrcEX/cFfHwz5uawYx7v5WE2+kkvjZSf/nklEiDc
Cz1RwzhMo8T5jiinsM0h9dDG0M3VvN3k5ctD5Vp1BWl9jhi/u4WccivCYWJmNQlB
FwpGGZrYd591TdEJHVuJlfbSuQRrNu4yopArh4MwyBiLS9XjlaQj6MFhyfpB1k/r
jJmlrIM6ZXCFnRwaLVnDMAbcF9wT/0d0z6uSHDvqT7FanILtsdJskAMylm1pR4XE
JpaOtwMMp5tQ7KP2aYX736J3PmmZ22Oi681+O0ruL0HAnMgitjzDfEP8FYmDGq0I
NrTvGyo8t0td+VIATPDk8X40inTVXApszgxJOxcypxoQOuOue8oF2QYBPhyXKeLk
QtJYMK6x0Jhl45cmyC90lwsbtY2zueO3Ob8+I0nfe68VMsI0BDi/xaxKl3r+DhR9
Q9aIh0yEj6PCWeUEMPvsONBubMA7k06HF4+fm3ZW4oeVio5MDd2MS+AsoKfHV3R8
X9IYcrWzK1BzDXOa949L2Gq9sANVUadicuBKOs9PjgRjsr9OCIjgtMxV2F52ZDf0
FCg67aGvqbMaZ/1qXwYx10KCGLiVYeuuJMtX2O4RG0+nQmKIyYshY5qFsfAkbxLN
0L5rh/z3ev+xrLDoO8lsKhZswzu6T+rIRrxCXHy1NkXRiDHKi4Xtr/vPs9oPEI6A
Af55u6hSd8fCE9SZR9dEtzhYB4eMY3eG3SwygBT1TsllLkbw0GNQcEXFbUfdS6Ny
mSUu+LbHK3iWImszlQT2wzRgu2Yoq4iFJn/fxbS1sgHPDRhRQ4oC1AHZuMoOFYA0
iVxqd+GLa06pVZs6JWWP8pVv2NN2y0CsFDa4/ZSJd+V5/VIZKjg2/6/z6Hvwqbqu
uL2dKsaowCiWyx/1qz8YVsdH/AYqxW8uf6/vCA3g1js0SJiuhYgv9bNe/AIrUUVd
gIYg76M3fvON8PbnS3lY1+g/lUkUp0b8wTt+uDh4Y/6OoT/0OeE7A0CJ4l0vN//A
YPdqtU/pmgkn8m/oe0VR/cV71+qm9oMmhxtWKoTB02eVv0xsdoGrgxIXezBL1EsE
OVjXgyBH0ZTUgoX2XUfRw/qUaiKCOlGkxg1pEAKBRs+hpz0DPQrfqS7sEhq1spPm
BB6+5XjgSK4S6mKDwi3gltqAuJ0Kdr0UaLxujm5ehPWEnFEgD/1twjK4b0RJKwmt
ufDUZU+DQ4mjia4FO/lVQDecx14zChDmuWUw4Bh0ft4U5df9f+ci/zAE/0RRmyr0
UT+khIxbDFSAQ1WRv5CVsIjGZAmy08wI6DoCUznE4bYlC+Z0jBS9kAExvizMhO0e
hS1E3V+xHBvVtMA5IwQcQVsoEmecCiB16QQJvsaGRoLmcju4b8w3N6fISh0l2Kc2
dty68REmtUqW0BCdJ9Fal8bmljny8WO7AYCTj1WzremrpT9jmA/dmS8bsZ/9WaAP
Mg6Itf7lnCQ41+OHjTHhxF6WyL2dvIzzm4UQ6G/chEM2Wj+m2chtO/PD38mGPS4A
ESoDJbHp6Q/T7t75i2VwuUq50Oc2sUGPYhlFe8CBcbXr/Uz7RT9710xA+3+kJxvF
CROyHl9PdNM6OOSkJklkZvHeoDE6mCDxriv9g8aG3YAKi1C3Km4y1lWgaINJFtcf
L+ph6Ax+MoEcQtlyaZ4hWlsS/a+rwkH9vGeO4rn7MGiwB7z9pyLCkj7aTa6hYoXF
BznDCCKBQEot5MtwGBVyANeFIJwmpWvtfF8xYJ7MMk3r/ppLF5q/Zw/6qYeVhw/6
yF2v0KIBoT3WMf+/ClBHMRqvKA/jTEakA8pAIYGPQbc8H1xLAotaExEFJh/w8wLQ
Uhv1Pka+MnM4scgEOY2EPFyXbtOdmr1xhSgC7Rw+37LJeCcdB9d/ufqfAogei2gx
roYB29xdhqyfuvidfsHyic3fmroWGAQHDXgqg+4mozZfcv85TKDrxgxfD+r7aWVA
ppPEqBXlG8Py7v+fxL6ob3wIOgxrf4d59zRBRxpI19BCzXxcJTbckikr1e/mHFFN
X/Jf2+z4jDIrXs5JUYBASCrJXYxfa0W9gCuwlLTH0L4omwJvHMzdPYJGTZrsp2on
QVwL4RyofEXUAtJ2BaEJWW3Im58lZgr/Ykk9SFYxFR9I/oQLYsicHjOoofX5anWl
QI/BEv/ZDn5aQv9ocWSPTN5pSkgsAWz3zsEx2a9Q2Iequd3J3+mBGM6K3ft9tEDx
pseLACiV0fKEVQKGcPYukuZ9npvu4XgD6MCuTJvgLdNt4YcD6eaf0Nmyasd8iQLX
oJP5bftJOnPzx1noB7c8SCEwpG6ChSJdxzZQkNGFeMf/lP371/E0F5KGKZpnE+gO
M5V420HP2Yei2JHACdVrWAqGDMeeNu2DXFzFiBsFyvr04wrsNM9JVrZKV3BK8ZkN
TTekaOprUWoo18IL1cLoXuI/HsQ+9C/e2pW23TC1nLHejEUFurdhKn9kKe8sAiku
jc8ou67dLMqgZh0t6IrkiZGVQPfHtzIy7C0rMI5IJh9iOoDi5m+fg5Dx0qwyPw7b
epNQbsF6GsRHljT+byWlx8a/dkKCpMUugYkbjqtovEMJc/pldRmBfXk1r8mf7TPg
C3/px1wFyRPhRp5i96KeD3MHvjtRP+d0hzi6lo7OiaZuvoeV6fG1Z5ORUUYjdGSP
vubR5t1pC8RbzXmCSqYEW4LpVpBAQJB6BPu6g4OxtPwexZfgf9jj7NuskLHHRTDI
Tpui92NFAof9sH27wr6YVLFWTaQ+zGue8TdULcCmh/+jGrE7D7GUHgDXzrZA49IH
3l27pHIFkbndwcXaCU87IPn62widS42urw8zFoV+xjSkACJ4OvQXCfwjl5hoMyVE
/N8sUXz/xIM/KGihe7UlytACI4A61keSj4HeM4TnotENvAp4FUA3Oszm4w2H2hhM
CLTbZyZboutYY+ys0jgAz9cRkUqdcwxFv4GjfDl4qxZ3UMy+25XzeFJkMESwK7W2
OkV5yDqNNrWAk/X9jt/KlirzEqZY8CIWLxg7iywq6JXocA7fwt/8I7kPDdA7fABb
aeqlUb449NYJDEkcvnzOuaf6GjEDmYV3H2703Rn1n/RvF+XnmF0Sk0UWl9l10ZCV
olbcdQ+TtoPtlW7p7tX4gOIDRTh7CQsx3GsHVyfwWd6PjsK4VFufeaXFBnjEOrbj
NzgejfpgL3QGEHY7aPJXoVXmlLc1sSP5JyEWdqKBi3SoPFRKM3BAp8DWs/N65+bP
dbUNc6y6P19/lJgElugMb3jGk5WiXMtog2ONCsAuZyXJm6fgZib5CarFbJB7HlyF
tjc5bF0UVihON8cMb9zOeJzDcl3B8WNh9l+/9sSIfIsmBjHbcaV2PDMvy3MFnlPE
yelD+Q50UG+4O1WQENiB+9RiFOPN9NHw4nb3ZXaRHnLJp+a/XJ6twW8+NfXzWSVi
ome8BeX6c1Bc8ocg9oBZv3VeDgiFcmAS0VOs7xihIy3r4uiDaRXb7kvwdSmyYFAy
QV0xVIQMH8hlsKBXn5PHvdFnIAE0LQy4EEbvigIVows4unZ+cTsvxkNlBewRu8QA
fXz3mxhbcpIRZNBFUnTC4ZoI6sbsPpL+nBtkNbjUtsx0weIBySZPlYIAMKnqRGyx
08qFLnV0UO6y0JI2FWZuEviLVQFY0woXagQuZiWbL0qTSWEKahkXJzVM0cTjPYL0
hT15MHxciv0eRJnaHVFff18QaNNamL3NIP8BlL6A1ksPQ0dZwOAF2IkwpMIrDirn
gXgjeeibrHKRBAG3s5wpqAizGnG7Xj4+Egbapf0CQl1fc7+mbJ3r/CkufUhYZBMt
LLtOpzc4Va7ZXaOCYztfBdiV1KGAP7O/sj/n7EIYqd5uDTREcEN1fYEo3G9Zb9V5
eEuU3b7YUgOZVEeHgva8p9YMjI2KHvYKrsT5O1PxFrvSGprUsurqLm/eJo1nlYdT
yoDXvdhmOTKYhcA0ywhjFcwsd4YZtBAZx2as69g/Y9I0yUR1K83s6ETJIarUyEx8
rYoR1Pvvm1+fnQNF2yydIXrHs6xDzMw92kFsBUDLtSDI1OhloDB81U3F/yP8w+6e
YgJDx75EVVCc8lN18VLiI3Cs/KPAnlqDK309RnMkYxXRxuvYo3pgcooHMj+A66ql
ORqVHOaQ+aczp0PWwalYQiM5Ju5djyfWU000+GiSb8fymjB8C2TuJGf4l1uRhIfh
tqJjwr1quBRjOL1JfJKSRbVsoDJCuvBTuAxkJA0wnJVhELhGO8katnE1bDbFMtIr
XIdQWCg+k9evkb5jZs8a980PWe4gXyhxPOSeQpHQH9CveaWwssKkY37jqGAldx72
nHrs9VwTxOS76NkgSw6wSchoWzkCxOwucgMU0RDAZ/BRud93qHawl0UIwNzuzrak
ZrLPx6VvY38Muu2xH7Ir4j9or+rU80jp8uD7YyJ+Y0E41maMT9JH9+qBeAPh91gv
k4b31Ba+KHh9diuBAHZWFk75N81QbPnJ8lcSZ/qyMVW9uBNl8JyX+9ZiL6UXNCVr
Wln30/1Fmis2evV8PmY18A+MwPMP2f4bu76icW6zafGkU/MaTslCy7NsDuRl+Xfi
1UpuTVyLgug6xKlsK/wmUVeBrrvyiNSJyO25Ry12aiLsrX9Z4Y9Q9csF76zLxJeK
9fIOEoLDtzwTln/ShcNY0tui4RcUAwSCYzpJ2RNBZPRnAZfIFzZhawOTbVb2/6FI
ePptfWpvBtvHbbPRwOvp7mYMfqyI8QVAFFsn8ewhmcb/ybEwQRd4Q09De2jiKWQk
BSPEO34WdGtrvvexfrM/Pp9G4qgRMETDZ8F/8mAOpDEMVZFFCMo30c5MinwrdoNp
QOo+siegHj/hzd8iZA2a2b91Jc0O3ME/kydD86/QhrGXDLx6OKWSjfhVzQYktwEW
tjwRJCr61kvXMUDZlV55A1BEFiI/jX4jf3bIjLXNSX3TCjXSS3fQ1JhT1cXcFh+W
57OxD5wYn4gRWmt1D7awzlEDajepOMusNL/hbaC2P1OB2cc3yk9vrcbl4DHFT57I
lXFydMD9MDysNP8WNfg11rBxfgvNw3Xn+eNX9HpAQQUAVTQdJmS8gUxn9Hbiqtk1
+PIYxDzUmnS8kNrurCNiUSjQxHvGAj3lJNRRRnttnMqzrOdAWx8zjCcWECgLpbuk
+l0WdyGhBC+DmgNLVHY3UFIUet5cutttqY+oDCkC4HTyZ6BtzmzewA5fChCiFdlJ
FnQLssFnk5d9yIO2w+018a3Wx7y/QNGWivNfgCn1BbN+6CQUeX8IMi9vTQSKFjBA
kpcUmSX/I+vlSZf/YxpX6WCjL8nlNJvI9hcT7zDzQ7NvFdla8AXx8rzigKi2QylQ
+HkYlnHWiWN04ybkM7/96/f72SP2ZkzZsR824tq1VmBFosMK+TqfM7BAqiFuSmgo
pv/NfrmyNfXPJEfkP1Ek824n6IicRAhANFroTO6p3Uewzdws21Q9SnXLUgK0JyWa
jFqrngTwEfkm5Qqrv16dU6JMTiEglsYUwlQsa0bcKAaLnkoczfMP5zo30u6J+k48
Nsvj/W8P4np7r38bPcw/5ArADYUGsTNqZZ84tUqtxuFmVBT8MKDcrT3Mrkpf2B9r
cLCpeSaJyv3ps17Az1lLK6H5DtDr0/dXSCQo0FlMGcmcqQbC5dyZ9xwdoOX1gy/M
VhZZiGJbkI9U7nQRUYpsxBLY73uWg/qyNlc/dnalCxC6J+05owZmlUBKfnQCmqvX
9y1soKmedTpYB4oXCTsfLUGlEWAvORL1/qqf2n7scA/l2RRJ9p1JxY3pLqJtnASl
GlNsPgm88v4Y150UrSZhXOTA3qayJGyq+t7cpjgY8YI92WjZzJA7LZZkjgtM4ZdL
5Wr9yVsu1Yj1vaeuVYC7WbO2XDwkuW7NOA33fHbYAVC4/zBvA20B066YDH3PKlM/
8XqR2gscnsTRNN13+Jv/y8VKv/HWEUgK0XXTuFC0jG/yBoyt/BEzfRBAbXpNsgRC
TfSFgAbzx636IRgciZwDqBeW4eQVAEuvam7rLojjUAcw11JnS9iZDm37U22wMZJr
xnWlMC1gGv6E7z1TC9+dvMPCgBK52U8q4/DgYqPXJG8EdIHIc9ewh6UmGJYoaV4g
T5OO+INsT2hFWRU3qvCk2nMg2uI3pWLN8nIkcE7tbPzKbK8KbWZmBLWH46NLGKVL
8VFQjsBPyFAJv2c4APx4+Q9v/ZQEJZCeACto0vPFlR1d6eMUDBfBBi9waFSOdEFD
H+8dM3Wg7srGVHda41cSFrOEtcADINEJSAjSUK9OniaCJpEA9tQ92UnwjswtnOIO
nPe3SJky5L13sgnc7gKPlKNBxDvA8OdaId8iFfS4M9iH1e36a0IGfg3n0/GC9YN2
Wlv/fH3rRXsKXrDzf8D81lhmMiWCcETMlSZPxZ8NGa2UrkEXeUT39niLhrAyIZ9U
Hiafzx4LlrRgN3+QsKStXbbeO4DIL+HZvxblgnRhJj/KF9LflzX6IDVB8uymd9MA
1dBU3vsoZX1r+m4zK347uxTcovW/ZtYv999R+Vqm7J5AUD4J+0iVo6T1p+cxEbto
utLe42SkEaukzAp1tGdidXL4ZY1bC5EzVrrX6uYVWH4Z+9K0zV/WisWIDzKlCc30
ehxMDsVEvQ97Ab0iqYUCdtF+Y6xpW1yx4u6zkrUzUoD458ajNk7VzvguKdJHl/1O
7qSnDAc01boiVSGMgkWUMVV1FNXejtDIenQy/yOQQ3L564pgiQRMdG3WumjNrCqG
sKr4eaUVGM1/3ysN31v7J7rfzUgDS6J5wtYqj9C6388UjSpXA4PdFCuckGktFY44
Y19BJJfrVa+f+HD62mplQFUPYdxSJkuq69NYJeZc51Mv6DZqyhtVnDFZt+13SyYH
IXMrQ/097guia3qwzh1sQ0HTYPJOo+LevXtts9oSyU8kWZq1ykmyCFH2BeMXJMFj
3lqPfYtTuVTnuGViQQ5G2qL/VtztZ2bQ1XBZKKlDyoVB+y6egYfu32gSIoIDWATf
tJiYU+J8l+q34e2uad6eU0ZxmKO/mVaSiqJIx1/lBNk/NxMPDGZAGhKpTuG6gKFj
lCK006tJs7o7TLC39AD1EdKL2CbRUTh9lxztr88p4OyaKyxPqq9f+tHWVACZu2lI
SiboboC2xwd2brvq3Q4HGpFP2TigQqRXYZeBxsgIvUGZ5AcipTiHQcGU7D0NaELH
BLwrJlvd6m67IKcFUyQUozZ+o8mdm+vbLpSWCS7mbvGJFvq2p1mD7IOhG7SF1V+a
CM1BeSuSGwkHwn3ups00Re8RIObJ2GxONf0PZEML3a91Umpk5PmjWRg1qRLHDb46
7WhGVZr4rr+H8mjjr1pbiR7Cey/L5w85Yp+McP6Pga07PlIMpdhSwDRSk84qIv1P
s6qHNxUEYUtuRRZrv8fSW1EdbffzCrmwf5gJ4U/d7X8KGCJIwBAmXYDDc6R7cYvV
c8IqlPwJ+O8pcGB5n1thv3yULeOL1IFX/MnJ/bRMDt/ZoeNH7s3Ce7Fc8PH8SZ/k
xOwjpb46AufWRlld3yQMSGTA2SQlupyOPLS1W3junC6O1mFCuxirwpun7JkByYGH
SmaRDRnrNtiLtFaefW4cucN/j5aIoLgkKn9NJAqIHj7pSeFyGksd0ztvw0wNP0aW
aEdXRk5klGwNnUiCfu+L007F35HLeelUzMG/Z5o+WQfnx1270VqDqGz1noS8nA2o
kBdoOQJpjTxEBLWUYl36/uGucUEUtSkyDJS0Vj8nmybHqrm7ts51bE5LOjioyNJP
JA2Rm9BCEhXWOP2LFheJikahXPYOy+3/RjD+DMIQVqmB7WOgSorauV7htPHt5dxR
MAiMmnO+ehBrOYwoskJu1INAN7ygSvf9R5TY7+IbJzYdZ35fFBh1icnivIQrlxBC
64yPDJFr2yirirf7fipBmFs5YZUxLnvJff6Xmvsu5IbGp956tlKf4z/E4X+Np9fX
XQWN1JSVk7O1pKDDKrdch1VXgbmBwFlkC/ghgEXE98hc+cDUbm9ieNUW6NsZHA+6
CwrEYTnmZi2x1mL7yw98Q5rwMB/bwW04Ksk+IA9enhJsfDsrXM3uiVxOmUly8BRq
Jl2CnJnoBnKqw4Mrm7VnD/vlcqRbcvWKLFx+z0T0edfeORf6kP2IyKHjudicgNyB
2H6supH2+q3yAcYk5PznXTuLQaLcpbc6s7JQIdlAIYErs6H03HeBTvJQ/FwiWW/D
KBREu40t0qH6fu3LBAa31ObhvydEw51OpYS+CaBlFxO81/ExIK0DGceR/RJQDroC
yqWA7vNMICLGwqiKwxgmlRJCCQ+km05Zh8C9FGlWc/EKVEHAa7FfOPxL8nG/7c1c
B8VVjJBg8ylSPxjDtWb9IqjymLSeSNJgBvl9ECV3KPS3BVYGnm4Jr1VfsJsQDdTJ
weiboJjxLbyk7z8CLhMf/pgQOJGl9OCTuHwcVlGMqif6t+WoWJMDXOICQTWZYa3d
koIAhkTQhC1XW6qP5xMMWGiCKA5gVYPGRNEu+cigg0POZ+yBUpTEvToS2cyKLaXX
ZZPe1cQcGKfhlP/1qULb8SF1gZRc5dc/0RyVTT1nJ8ajt0o9OSc7A6PZkLErxo8F
1YFMcjn1iwV3/lUYCZs+MSNfcXmJjNUKnfj70vtzog1cBdUWG6KoLG9rU+p5UEma
mzjTxSVaGgYhlkhKio2MIvzA9uHDbLdUj3Zodp63F8CK88PiNjzLjuTJP1De8um7
UO84MDYLZfXF0ZOf0J5WVRDzMQzXNDti/E8swd51xxdV0dpcZ+KvfQ0LEwh9MIup
4VbEa/U060YKnieTiry9BOEqzTwMKfKjvrxJeupzwIZjGMbVPxEg52LNZvlQpz0y
vU1RfNNiDqzx0AGX37MSUlcjM4XdyS3ha1ROaH4/IiqmJiwdZpqn+DzG2KPVZWHI
k323pm2Ld5Y/nTGGp2cxbpN7Gf9fHajnyZojzA/iS317NAYHANR9ldH/TeG5q7/y
XXUllWOoV3box/L8ZPPSuGC74M7Wrjl/gsI0ud/x84MDBSANksCo2TVkulE/4hIS
Lh7R8O+5IMRDWWc76HQS34+ScEZDl+TineNCIB/V/lfNFMC9PXzvLwQsKDODtxpq
rfFhXpDPLuhREqAoDlT2HyOFIOr2AbPG5Vm77Ls8Ss1iwkyXhze4vP3+8+Y8lpSR
gJ1rv5+BaJtM6Z6XXqWMvVrQUXtDWA1ZL+S1QpM47E+/z/BY06TiDQb/gp8rvgps
Ji5vwvC5dYSCF1EJ+8hqKWr6UiVzHAocx6IyVVqY50MuqWLA6mA6heBzBcfsRH7Y
qjxjlV0pknWnVQ+KEWQCfT9Drz7nQqv2TC/MtVbt9Kx8Fqi1Ic+0vIwjVa4Xcbp/
PUFkwU0CPB9mWkEo4Pff/858yStWsP1ZWj6S94GSumEvQ/DtBMKVBSquu91LbV1F
dRqzozCsLnfbf+TcDp+qwh+nfHLQXNjRvH2eK80YmLDbs2Kz5kIaLJUz8q5n46as
XabBN6ExQERGvkwmuJvMtxbDykSsmHt4vh4EN9H4LrJBBiah4J0yYTwsYkDiW6Z5
Flw2Fl72H86kRZxDc4ItMAxJViXs2f6wz0VGQ0DBkD+UbO9k/psF2LVJhYzclZYm
PRls2o6FZTLXStt4UV7Q2HazYRdO4m+muL/dykKt2NnYLg1P9FTrVDkAF4lM/hiD
83wlXyeq30b0K3mrJ8DoPQ3Gy5xyD1eTr4880ZV8m9iMixukVMsYVR+sJ8Le95UU
aQBcixin5MMwQMIuAOV4cqJau95VA8JSg/Sk0kqTRh09hXhlTDJCKgDK9YirSt+0
L/mdZTu2R7exewt00rSwI/JCkbGvqJK2kUOAeNE2E6zE3ob/LvGqSVf5xLXEzehU
EcRXvGv44pDmWDwHXxaHxaH6KXyRWufP6iduSYmL6qNRq5OOALWEtwjzGFYOHxse
boCAoWZK2npJ4zDV9DlrZzTGdBkdoG8by6APA+3s9XvzaPzQfDWT1HkzDelW6FpU
bYgt5fxeMfQN1jduA7AcJdcttlAf/Y6AIvCz7MeFqEUl1TiiYU80nS1xmp3MLDGS
zkTlBMpm/C2+dplr6vFp+wU1T2GjV3RLDoK57gRHBxWL/AdUStSdHHnNCfvG8qlS
CxR3Z/+LVCXnw3Ewi8ASBfOooT9dR0cRFOAVTqOnvkeoYjPkVRMk3xMARRQ4N8Tf
57z4CeGrjt5IVKMpqVmHvScfJXKsAgve0yJFllFsE5BcLp6ag1mSvrsmwOVPQWWF
pRIrzn4pSRFFoanZTedBDGbpPHpwk9bq0KBE4l2YMx5xXoGbtVWG3cJdYRaEet7n
2cq4cIMo3LPLgtSQM6jFWsS1CxpmsKKtw2l0wVG8cU0ATmeifwaoeu328UvvNj5Z
0JmZqf78RF/mtvlYW3c+ZYM4UtbO/4UvG3XMX+G+qXMH8Urhkc6sjKTVUxWSi3Lq
JVCd7xA1eF5UoLmEjIhOYBKxn8bhEmTRXHsHl9EJncj1p5NiSrwg/Vxt7KH1yIiM
cIN59I1ndVm0KfjW5TAVqxIFvC5c4Gmjer96bOaiZ9yv79fwlmBMfg+OjBX5qDvr
iKGgmHTG8a+jfRqztRZ+fqZaGUk6EyT3vcF3/shmKUTG6UrrZPZva6xFxSSU1Uzs
/OHKraCY/We8VFzFW8wciCAFkblakVjYFXRlY/fRUTd0p6Veg9GW/O4i5VCU7fCo
0W66howYKYfYcez6JfPsKtLzjy+NeK0ydV3q1J+/szW7c8d8F9qj4vsyFScNymx1
VQNaymNbsa4hdIrO53fcU5a8rtJkFC1l9Sk4eT2V/9s7IG6MhwClGJj7BGKukg3U
Jr8Uz4kzbDp7+MKu81avuB/iixzfmuMII9SoARLd9Kv8j1Sjxqd6oz4NpJcbfmEa
Gu2Y22Ltz9jX7BfJK62mAX1TfEDrC6tgnK5ET/TnLMRY+mRh9pNVmjlIR6YIudd3
Hcz8ex3Xcevk4BIjfBRsHMFqMhV/RZUK1qWxwmLEYYywpHGj46zv4Tl9A4p4D23g
c8w2U6vAeOT5W1rTfEMJXqJ7304xLGbqnDQIFOTHA0k+x9qkLq8VscodU8XvyQ9f
12uPz+y3/3weUhPfkfm0qrRcrHIGJHFLIjpYGf2cNCRiYZvRcpBNF1aXRj+viZPj
vIq3lW+N74oIh/XArTjP7ZWqhuf+GvbISA/yjtfFHeJtzYq34LroZXf2vf7Sb9AQ
mANHm30YKdkJePk7E/naqErvSf1yLkxLFMA2Z40ckWHo5V3t6+cbJal9IpT3mdgH
Pqx6vRfCJOCZ50N1NpBTYFhrYHzcC1iL/RXN5fKr7zf8EjZYoC2BmTDd8W11F77P
0ss3dDRlP8sdGh5jeH13YRKPRey6FCPjRdmYRSGbzpHPZvQofBabtQ8ATsKSBuAI
kB4OEvR54SDA8XwvDAnGikxytCeVxiaZDA9bHI5XVUEANk61IiEozFrBl2lxYsfl
aY1kY2LcmLbfu7YOGnvp3bBsr033Rp6KpowtXbL4y/Kdfn/UOp8Hvu31/+g0x2Ka
tVr1/SuNZitsDVr2aV2pkattjyFDV0m4qHXj2PgSYQ/EqjSaOEw+pGEmWpe6KI2v
kAHDiLIFFb4z9HK+vIvoza9TMxZ53b0L5bSyGvtqm2OfgMtT9TCOUpMmMdcRnxp3
7EBi8DsLXFXdyW93xMHCwkY+EEWrGvw3NSz1BBOoTabMNnzd3J5YQAajKcG7YS6m
am4nfy32+Cp0JlVTMQoD7IpZdbiKfHIPrf3WHpaAQnPWTncMBL0DIOepmhCXT+lI
i53IF50Tbi0QpS98v4WTyfR4se4+MGL7DTQLFt61Dfa/PjfjFVacVPt39CalUl/f
f1r/iV/Ae+k+M491gKp3SnWxiiG41KI0IyFnL/l8+eO7ztputcUBciAzLEhM9APa
9c9G2o6r2cTvxNNwjqjADxfLM6tohEeKUJ1sSGIa8MKZTnLkobIJE78Vq0BKPzYI
TMeTt9Lil8ghuZwaIv4HqDEJR70s58Eq+hhjir43CdE/Hm6fEDZnWsJaDsLdWPK0
Vr+CEt5o79rnioCDRTP3BhBwWNoTS9d7N7T5I+lpgJop7/h5SyB5GiM9ygmF8xYg
A/hWzRv5E3V4r5FRF2gIGMp/Ba341zaPmo1s3AefkvYEJPGAW5VJoDMGXnYViZQc
1Qi+HPYH6AlfJqivTuPTYN3pouhLDai15UWT5uCAiohSrFLzrSix1i5itCHEBJz0
2TC19QNrB/CeGDoILOnUe4kNvGzHNP9iAIfUO56ct/RkukG1j/rv/9V5TXrHqByT
uwgHh14zeAGE9ojGPiE0sbb6HsBTu+Ypskl0BH3ERCscvpI5E9BqqDyC5G6fPfEu
OH+AH8GiF357l7t0JfugaIZYLotEBvbbvCFnEi23p+GPtvZjRlZSlN+Z7gAUGAVD
vuDstI/vdMHDS2i9+G0W+9AkYf21M7tgmKpN4gxY0k7Wlf99U0987JtpZq6EDwgp
xBBSZ1REFAbfPNzDGoejxNjlE4XXCvFpfiK+AE7sFESuh3IEZg4eea2Cl6u4atv3
42ISBPA6NWjrta0uyo4pRwQNibTywN2Ewv2mQh8D88jnEB5tArLDIhlqJeZFg71a
06OlNmJbpeTdD5PaT0672zdijKC5fWQXybH7swb1S33GA9DDUjr79Cm+wXuietqH
0rNpqHnlz+M6+jyEmdUeczSgxoqP+Tfknza0DN6Zk5w7dLEbzYsP04l0JSezXpyD
TymcqwOHit1Ao46F2zYjVdOAMkQ3iY1d8A15sqi8Ma/LtFKxWu1qnxYet8rbzZZu
+NPhprTZ2XxgU/mT0iTBPufIdjSREKrF5RSkby3rzCNpUEtXBW1Fg29FM5/C3xWn
oW9iLx8ujWxpqTAJzIP86PTfbPM7z1ngHtTbInsngb7Jx4ua9x8T9YGjlaChFgTd
jhYs7lI0kGAu0kcqk4FcCzH8akVU785P9zPb8DRdrSo4JbDOee8gpqHzLKVxyvtu
joSW7H9qMbPAwr1IbmWUiOIKOSSTrwqyufsnWPsgNpHFKY8JgsutMRzHC/xjDq7k
ZyMGA2QRh3OvWE9QuV7SrYkswziSkmpyAVfcKt85UmBeCg6LywFvJ5642IH2lLhx
iexUsY/n/Hi2urh5bJwf1fMjqPCZQi1iOT09FjisZkAHbnEPc7heujoQ1WUS5HhB
SCy8w2BAaDWmAGeOlN6gcqjusSYjO4i7irWp5eVc06biL/dMTb3Vzkxvd5zxbuT3
y2Q+8MNeKpBnxqTcANEjjduhRyWHDlPbh9EcnE+7YWmBmwITkrA/hrSq1iB4O3br
dboicbBEeFtdDhIzY6qvU3yfgz39pSDDwZBeMja3GzynRuW0zG0Yp8eeX8wEBaiT
kto26BC7Gy2S9DEmSZtEuE7sGlDACs4yKd039ATrBdb3D+FUnALtm8vOQi4tV+tb
y7PLFLp9uqQ5x1ta6ztF8qcTHahF8mZ0YReeXBAZ+MX6XPmPBlb15DipL6dIlDLo
GpAv0+74LoghQM7rdDpLaGzqXj6fhhUraiPT+Kn+76WV6CyTQyMXomDhKXGpUhRA
f0z5bF7J8xv/ulAoMWU4DMYABWQH8FqXm0ygbX47FfKj68JON9F12IMq7HkH9lpt
0x617OU9IjFKed3Kmi0wF9zx4tnXLL3gfwnpHms/9/OR0ugdswS6MMfkPay98pkA
rK0D+Oh+2aDdHp6nrjE1mozKi1qgjiIc4YHkRv1dk3K0mFfPoWlRPLmljSz1hmzd
NeKYJ00yp4Jx0bBs8o+smU97bMLLg+m9P06rC0/NBZtiwQdyyW7y51XDpX9oysOD
osCCDymKkx78Z210h6FYDLy3mT/6MQrOVYryOlR36diJaNRZA4oBbO9C90scCRfY
yohnn6Ao6kbAzPChIlETCoo5apygg9fExJ0E0/oMNG+8K+sI3sSfBLCyTeWHf6ir
0USpkS2X1CNgPXY9g/3nJSuSEiEma2x86IcHa87MZGDluj89WSDXJKV13lYmSP1d
e/L+Quotc4ikqN4qC07PjVxmCR6omKjNT2tYMl0oheJ5KOf9A9gXiiMBeTkJe7qs
CzS4aI5R53Az9uo05vjqBxKtN0oyyQbUHbn+AJBsEUnm1Oxyhh309/sny5C4zE9O
COvjUIxIGqCU2ZXSadRoaLAzu7hkE3SMaX05Rny+PUfc6eWEFh46t5Khn4L4TuiS
o2LI0ENNcjx5d87knQT+hoM3kOL9dhWglzGPcn3HGdcCyvBvgP5/LkcgDd8Ty4gs
bmrLiiOr//i6kyG58300uHaxRPSEvpC64hpf8FBrnv5nF0OJZQLRy1tSxQAzXKSR
isRdu6PCT9mJ8r3U3oVEAEeae9DFoBCLWS/ItB07hJYcgFLb+p9j3zp7KG0DruIr
immo9LiHvvl4TDBRAWVCTEgNENo6P4mHR7LTzgARQk0cwfKJY/VwpVuZ9yfFVwEH
zUtDXttLk0rwmRunMJrVY+7t8A9PQ/4Gufkeldf5SEXqt4jNvDxFXbz8AW6kwOcE
q2mzKzQkU1+95vsHbhtMJWl0jYPCNOeTXdXSpdBxqEQ6xiGw3M7AqCtiy+FC1ww8
1CXws81YF+7/BWaS8r+9rsgiTNtA28Nrv5iXpYVvZ5/5M+BpNvX9p/oAH80UnuPQ
DttROBaZQ53LAygpQG4MSyOigRUFqxjuXNXhP1WLtOKLgceZDOVGDcR3j01Vimhz
MMeVjEjFXDcJwzFfsEW7RfE5frGg1971KQUbIlzyWzs0V/8UeXcO70pZmbhJ7Xrk
fHTnVcLCuX7ndAAzfIqtHWREk6JyLdnP8PHfoyq08qMiHhmTsrU9OBWHQqHG1V6I
WCeX3Tc9+fW8hICCXPe8QwaWOgQBIJsZ+YRuXFwSTELsajd+Az+qWh3nQ5WGBTSh
j16GtCpR2xM6Td1Pb7RgRDRcbcjkItsFmqQ3pJfzn6RqPLgKmTLtQBbGwD4NZgXh
MA3uzpJFHaHLGiQi3rV8N6/14vvcMWhaulwcofNzDaunQ8ErY38f4Q2MUZSXBw28
Myf23/Tv/6OEdyPacCzzz4yeWHXlFK2T0VgLVb4GY6w05Qf3aFY+3Mpt+qKJkuOO
ELasSrA2ah/Xahq7oX6UeeAzMBX1XA8t64N3vrM8piifvm+2+51iKvOkNBVo6ofh
wFw+0uZ+eGCHaQgWDUEMCw7vqt+gMdBxPrKMoZ3Hra9m7wYSPlG0BGjmxRgBDoGI
06eNsvxJC7AgbKeLlGJG16pGDwKQ6DmAN3alWSL8ko61FU+/pZoDGOZOFEhKiVN6
HK5oLHIZnusNRYkSYtDUzN3LyznDpwaAmf9AWXvd1OW2KwJwYE1Pm9SoaWnLTe3Q
iAavlbuVT0UuNtWEst/mnnGkVH5cqiKP8X4UUmcijO4TKKqPnduZKdyWTosiJRKb
YkVB945UgOpoiHSfVBq2NZev2s/UF1sdY14ZdQLCUjfV5ZqLvEUBlhLDBu9cBGHg
/NOOLh3fPKQoQEshTxXLPJYFlOJfsWugSjZhhW2h+2+CtM5wGTEo0BhQ54ohzi4N
1lj6fmQMxDdthPvm/0ulnDVhkCaWa09n1D8j807Yj3b3O7IJaP2IOTVOseYPrDOg
u5ydIScQRnCeFuSFaN770smYKH5akAubTVTr0m7DGTmrqZUTHqGuGiM7gWD9JcqR
Yyd5ZHPiJmy6QtbmShuowHZe3vKBeWBuSXdtxzKMOiBVqqcoywam+dCrfiPiwD7z
a3t/WnJYymJkIjjcq3pkhiflh4XnYtafk7O44YjjwdsVT8XwhYobsgotoIzcrKSZ
b6mV8UsVyU2F+HAYYj6MdGaGiWGKEIOmsAE582+QOjRLX7MBYeNb962R20zD4LgS
IwBTo3SwENPbNskzgKW3Y+Pahwx65C9VxdEz95F8EDXc5ayUbrlI3MqPTHbXMT5n
DA4YOPMosS08uT+3qUF9NCR1NBuBKORV/rIikU0YX1NMzpG1j6PtrHcfB5k4mdGx
QH/mnutrhVPoeKOMspAlW89Q/OvrfZnD/jkEVGCY83LHyCeq1Mm4c2K8rY4j+2xS
bJvxwzCbubevuTaJLzV47MRwq5hdzCvMAbccrcExCfApogoZ2u8NJZlL+o+zuA3R
pSJB9QCBO/cUGvaG/R2G+XAr8sifcTedlzKCnaxIpEfG5YDalutJVbUTuQW5f0xd
6BULCWRY7S7YJOWLO5e3A94u44ZErvyyxQr1xDW7B12koex/+RfvcCiOgcvKQDCC
jDNhQt/Mbbwai14SzuC1/WIJU4kSnHLUapg6PYawcnPCiya0nJWgptZfD671su9D
zO8LLTxN6HyV2GKY2lwA9WlWgD84z7GxRuvCzDhclvk8u2oY5QR57B85mlA3da4t
RgYaVC8ydNfMihObckxqx4InrVkAHtIDxjnetepGM+jUHnavlIYS27u27c7PfgXB
GWMLnL4Ju9d69ktB39GxQc2+IRUVI0Kvk4jTdhZ4sEEnJgnM1iW3jXhZGmlGeoC2
yQmpSTJbRrQFN/lvMktS4fiNMgWkgv9OpLfg8cPF+0lXETiKUE3GuyTgqV+qH5QY
+GQcnVQnyQNyacx8DSeKoyMy/Zr285AV2lg/4K+FJ3yUDDno6Y2tsivFjTskRe42
h7G5bEug068hr23OOx7s3aGs92sa+x5akbc9hCDjlbBS6Bx20nfIBUtbmnYUfZWe
eedmGJ+kewYpLjfgaqgEFZ02pPDzk2/hSEXJWU/NqNpFN37+VuE0QlWWiYn3NHdx
b+nw4azHS0/DD6NpM1w0skGbyr7zb+M3TLOPWndzlIeuaJJRZQD0D9oc0cGy1Pby
OnAUZQtCqbNyZu9S4NYTEvmZme5DGtCh806pkztiY/jmTxUaXV9G2iUtKOcbVIFl
nnHocczlmm1FEN4GhJXhb1IX5ZXMeB6L6qHU/gXwYumJV5BArDNmm4T4hky2/p6R
x8aYrgu+cuosS2HA7+9Xc34P0A1Q0oP8+jRMOTJjFVUHmXG+6wp2Y9/Ml5ZnPFAl
oKqn3qHKrNhWghQIkGpW0OpLy/LXJIRtBsm0kVtZwZpSaUc9qIQ79UEXZ9gKMhma
oVcQ1nmRp9yopvkQKA86o1QBqfT6CDjLGuI8xtzrZIqyZ8seBqRzyTxzcLvmn3Ad
j49fFbG5zeld9pXB4No8f/D7xG7g26oIA8RfvmVFcCrHUe5+cLYhb81ZJdo+LEeM
cQD2S6bZN5HWiCfaVBEEsH4FQGIQvrm2CXYCGMWGTxYnkRs8wtEiDtVaDiBdPvMQ
3EYworXuDijHpb5BxbELmbBTXUNVIqGFKOHxe02CFQobXi5OPk2BlUb1torGRU4c
ZCWTqUdCgLAMKphWjPcl3sgzhyF6Z4BKEfSkrHa85MMCVfR5MuqekOWF0jHQxrvm
WXOThL10otrTnhnPsQkpHG/IyBYjv+gKtsMiMvDParVz3G3IqV9M00U+F8tGzqAN
mGk4Xbtqs+jpn+hetlDim798mnmfNHs7dHXd32Gqm76RQSyrpFYnJVtYCGHZyXF4
9es07WyuUmAckrXhKNFVoFbWdEdXAf3RAdiOGhZhVv22AoZANyuuqpjc5VfHRUzH
eFLv/oEvvjMJjaimgfK+/ydzEq8lRSJSOyvF08RTO56Zeg32xZSUc/EXq2r6+QR7
k2R766ZVAJzoCybEJYUJcRBrlQ7KMzTG28QDJzxpR8SIH26ofRcOgCYz3fXEBuwb
IAGnVjtNwvnL+S8w/VtCD/J25GC0KbScc6lewnD+DpitzalyDAil7T+qLwnd84TO
InZy2LO9a0xcLZAQZ9RjIY7nofcnrwp7v2UyPfUSik1ftp74rnSC7d7DjmD3jK64
dHIUTTqmKDuhM61tqOdQ66kfgzUu2uHAm4OCrK/xy8SbuhitMPW32CFpoA2SUxh0
tB+fPeEKQxmYi93fSyVHfmGXoonYFX422f5ztMK3xbmHqxCskqo5TJhxBJkW1LSq
tO5LO2V8/4f3WyswFW39PZYqj12+BBEslh8TxHvDNcdpfEUVhPYbFyLd5r1tXmbf
yrnc0pcZCyuHw0l8IcjMs9L3AMoK7hotFIxH2y81Mymz5kp1maDgSeXv9FzT5nuu
zlmNVSy7A2WDJmksS2zlzNs7EiK/P4Li4KuGL+2RdR7taTntIelbzaYTLQ7+lAwr
nZn20ZFqsDpHKthjTR0Ma2IKHa8n8lxI1PiDk1bpTfVE3EB0dNQnEgYWSGdKF57S
QY7IYyAUpeJvNyk5dGP4DVDSipSHT+XoPacrEyFtvhhZGA+sPV31HCNcmc1IoLHO
9+COyCvCejoo6tSIqGfqnYN74Ttf+eup6Rkt9zSUk7q+RiU/1f4oP67yMWcsCHmY
bQcoXniGtL87f7UfWrzCPkZc54mOtOxi7iHqBvt82MMCirTHpMPTsgG4Q0N+KFmp
yJZcM4SKQaHmzeNLZx/qmBXcQDiomd8eBpEwbQXOtokw8szYkozTOK0xnj5bRMni
c0kVvXyklYyeDeqhUFsHyYsj0dFWNMIBDlpY5DeS+aUacTaTNqVkQonTtTx+kIIv
jY1pD8FpYaVQGeqZPcGDdGiOko46WB6IbYAUe8lk4WTyi8Wwx/DeCfHcCzbEZG0N
/VYljgkAHSi5ZMStwiwN2y2UQfAFje+Ac0SSVf+Izuc=
`protect END_PROTECTED