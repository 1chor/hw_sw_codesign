-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RqOQBW/vqUNIoarUpq876FSM8sKGMDvPHoJjMDHX5+uj1mXi5KV1IztZFj2k0QyVI6oKFDvEi+he
XsWDc1CnwDCiYtFHkwzm588HXuVmrovXwo1jrpwDZ24X6rDGmABMJO+qFXxmKARpjifjQ4SQFwrn
L2nIWd73CBhIKiWPYkQsOX2ljxiTDNcjtC4VZKHLgwc3ZCyvTPDup7nArdspbrwg9qTqpt2R7S8/
0ERiweDg6EofvCWF9bYId0yfHHfxAUiW+76PSTm6R8MrTwRSvwaNsoXt9Yao+wuo4mPwBIOs8Vph
fwJPC5ZZHfVrjFnL/I6h9TC2tFBId8bL0/D+/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9808)
`protect data_block
Cxck5hemoj1zyeJ/nMm7nwTDSf3gAOHS5BAiALS60EeeDOXJ/lCk1GP/IeqdhkgTZy2I0NwUB+zO
rrgNmuxffxt0brwUouJKD70ldzn6jXUPGI79o/7Hp02uh8chnPtGRxVpgsKwV6HR2GblRmfqdSJr
0EKftqTlckK/EZmN/y2iWLXObAFgzJfy6pDRnOt9Xn1mUy1FQYwqowVqI06ZIvI59OPlwvymsz0b
kDrNoI/5Vg/Mwc8UGHBY7h89gVV3ebrWXIImZH3GNBY+1YXIZsXE33le67vy//6cAu90H6bdnDAV
FBNXLQj/qinJ0l6F7YKdimogOdDucVzAf5fSlSpB0JdlMNm/45msgsAfut3jqaSOsrKpUxguaL2h
qiD3YZm40MD77XFrYapmhP7cgn2Uc71VTfDPGqGA/4fP28PvVvuzrAvzPiTVGCcZXMjBsxpV8oNg
lcDboZLp3PaUbcbWjjbEaB2DzDlSs6yd7rwGIYFtOAHSfRRoAchiq0SJoA1ZvFgkIRSbuPpowkb+
c3jLYSeIiExkvE8Zsm3/PTgeNDawQYUibu7jzFSGxd0HpPfF97VrSrXsrC/TNfQabmdiz1zw2JRk
ZEn9tvTP6YCg/8yQqkl8br3TWTiqJj2+qTdttRkYy0P29/6o1sxWxV1G+tMVkDaCUtITekRYqVMk
fLM+aMDJKLC9sy3WjPAFPYJ1V2+BBWfBqLPW4KMffoz8+++8RtJX7bGFEUcM2Bc42Cn/asQ3HqQD
FBFejEIPmLpJ/aVEkI0o1xhqEQNG1X0y8XtAk3Z58mdvY6DRW9XeN6RJZZpLk1D/FbHXVDOH9i8p
U9S+fZgHf13tTCubCKBkoRB7h4crELNMIdrbeIwvlY9PsyrGa70wMJgUeHYpWY0wHsb7FA9iVY36
QlcyQJp+KYL7HzXb14L8vdWt2DCWxxjzH3bJvodwPjAHTGzc6KjCylKI1gwNOq34Uzl00UTz88Jo
LsuECPTqMGJmLiefUrW+kXKlykrMxq/LZCPcHAa5Ej3WEBSRRe7ubgX6Pq6ZypGR6utSAhzTCT9A
r5+oQO0lvW0ybXx09l5CAVvRH1IywQUN53NjnIxAKDxwfnLqDP5RYQjAlyvF1O4fBHyKBBF6nvgs
Sqd+DDmCUWU1qRBGjuKiGN3SOwWqjLLVcfr1XUGv2VjoIcHqgWRYZKeGsYAyHtuG9/j2bruPRRiz
8hsPb8aa5VrRfnklbChF51aG27Fvvh8dH8JVWKYDdhCJl77PzNAzSmuL6BavEYHlctdHUMmglRqk
cvcjY6pjI5eTj/6m/lnF3bB0GtTs1hC4lNAq/KtCIyW/tAiyWyKXGBWeV9vgEW1GMgsdBcrISyPB
SrD0qx4woPi8NOdMsoGr9WRW0pFOVKUjQmGvqmDUyPg61rsm/FcUFnMfzdKEkk+dBObYY3sOn7Ac
Q+YvyyO7qLAuuuKKSPMdxZIZ6FMHCZGdumfHhro08dcW7GqxvrJZzX7L74rf48JoJxNKObdFo8EY
ejwA2TiNJc5wC5o8ec2mbYB3+yV27PR/fKHknOqohMVi4rasIepPFIE0R71bR9rjz7+wl64dyFx0
/d34d1K4CnnTncVEk/DI/8B8dw6OWVvmISMar+ufIV+qly8eQFK8B1i7RuB0gx59Uw9WQ828rWlT
qEMCxKUwU3Bkwl+i6xLhwvL+G3D0YAQgXbBEuMOVhOkP9Gm+/WjYbydrPJG98YcyK9tCXtaCdq16
Y1YUdMfU1Nr8MMoxLdtbqGU9aUrxFiuVQlZpItVVF0iKPs10I6P9gGyiauAzaWQu9yzFHehjImax
7q7pfJPrwFLDPyKVt8mcwZMUYU8qcLoLwss05VZ658ZPSBgZYSOy0x7mLeoBitXngXhkjpKXiDre
sRMI59eP5qWTLADAby1fWaoeVlbFv/PZbFW6iEjpfoG4CQNHiNkkXtlxK9EReIAw9M7O7ivXTqM0
QXlrq61FgFeo8FFu0Ohe4Y/z5HEh4r4hs/C5PCKSjLlLQoFXttqA8Gxoufgq71Gbw7QOdy6oPmUe
TAf39mSdEXKg9nRAL9tjHB8sXwLP1XLCJ0/FL3DYxPjcNJ1zf6MBdf2mvWvj0yLAv/GK6KPjPwPt
QmDntO+0siPmbWf/lBt/jNsnBh6gLgYa289YndkVKWqK1ntNloF4k3eyxiVAn2dmmofHTrHaBRn+
xAKCnDDhFy218CunfgiUfQC3g5pqWL3HSIhE3Kzt9iDFdM7rueFxWHosMWNbHXev4XPElDgA4IWy
2uPx69yhUDjIIlQEi5e9Hzk5vPXQzraLzirEFiIsY12jvF9PJmqloVg9kllbiplFHV47xavzg1i1
l4qR1Ong7gFUD3tddj0UoOUiHl1Vx3AUikOl/R8qg7WwinAErbEBTQHip0N7Whx7XLvLlO67jxAz
0vx3TxUoqmTd+YXw1q67FR05ZS3DPE9+DXQ/SW5zeM2XyeGwKxnVSKug8+j3ynv8iuR2zPcU8+vm
QjktYF6HuO2udA8LrTXj971TAjdhb8ay2gZ0RE/lywxpnWml8rGRYnEN5JelgNUPUkGypwS1/pHs
HNActGWg+Bc6f2xKOedk7s8yrcjgrwGHB+SvhYu8sHOHo8fccw8X8PIbBf+mtjj4PW2OHSTQrkaO
sHLqsnIP/gv2HpHZi58YXCpJsu9zo+sMg2YyOY4jX2uzS0RSJypgzDci+y4BK2nUaff/I5mZfALf
hJmaYxUoqyXPtRj+XlO83DZUUWl7Nwl37P+IQyQEeMY3BQxOps7zlzuCg8pBi5n4gscJoiYzogn2
2qgimur0xYJfXnsy75P0+M7nBV1VuBCKzUZL63hy0kj6CbGwKEFLl7y5errt0JQZ+PEKOuST75sf
qXokanvMlT7Cu3uzkE48TnGcH5Qih7UDAcpI2o7WPPbqloup1LQLOdOL3Rfx/0x37eS0T9JIgNUp
Zo2hU+FrVvQ4czdftMaHcV9A6VX0cidf3X8slspMtYcBHuEJnVun1BHfFiyMUJ3Djsyws3lqDZC0
aNf9WD0VsC52kVc3uIx6LqBvLnMCh5TvD1PWNxyRud1ABMEmws9mQ+PpmJDo8LZ3GJUsof46KG+N
3Wk2DZhf6/y0m/ZE1+Q+ok6KvOGnnYv+VwuZbDtDgiW/o5Sm9mkOVaQ9+dPP0bAUQUS3qw9j09qh
UaS6huHF17E+0MzfHpMlPscJ+KhjeSDOJ/7iWulcVxTKRa2BkMU9v564lrT8xYpsyaa1D2HUrHuC
faNmLlsToCNiHXwkXPYVbklC5/l9j5+09VNwE+52Krglv1nlQXQqnKzHyuZL7JQ7FoGhTZfrzKqu
HyW4R5P1Wf/sLerSAXp/oChSM+Qjy5nuZScYTHL3MoA6xexiXzVyc7n+60HIssqKhKL71UShpks4
Gzu2cXIQh47/mWRwc2t2BvbqlExHGlV36C2dooh7DuDEcAuuCruPMojO1bPeADiYzes/4qr2zifu
GOgcFmWKqt1k2b1d3XczjL8A80vnN0NUn+tCvvC/ZJk7/zFJjfRs6MJqKu/SCcwayoVq0n9IpxYF
Dik+IPmpgkobKGsr6aOeJE0RNUXVPHtFFiBZbJ1QZPMV20YsyNZmenj5FjK2Or3jTW0Er6kVNBc4
93thW51HzNApKvfG7GpyXJVl3XsAZVXrVkfSOA/NfxMAizI4jmYNBDpoNUF2feYGC3rj22PfKP6e
1YC1c4bbB1eX+okvy7n8VIcPn6qkpB53/bs9lCEIa4Nz1gAHS9zJrCfBqwaClLULdmRv6oqZGVwa
oIaxly6gfwCABtTDAEVIkOa5RD7XJy5lVfWaU8rrcL2Ix6hwmQYA8jYmzFYWoQuM5jqhaOHghqoY
mRrKx7vFO91oBRM0B4U4U3SUjaxC0p2Rdr/oXMw4Pm9TvDr9hsMRGqOU8sheLSwW6R14IX8BI/43
J6g5PP9In0CqZBU3WxM6u2vW/eWai14oZHaDf2zkIJBIWJTlhzXQG1f7Unp934nZsqtYxkaXbIZ3
0vgofw5H4Oj9LevzzOydfTTNc0z5vYBJnnfSy7KAo/IU4n6UH1d0JW5I+HLdLVs8xJyXt+g+37jj
cEM5w9UMqCaTPGi9mpqjo+dHi/8pFHqMkxQ5ZDRtRqJ0eRsewIQ2o6g9ldwU/EbmVuJ2sKjXRzl8
Uh5+27INWLY/WNwEyCaMCGXrfLH8yeva15yB5VRC4ZvwESH+dgJaANBs+CuiKLFDSGN2ONkXj8EF
aqh/kI48DDgBt3TRd9+OSHHNORiB1LZcwJXDHDUtpP5I2Zp3ZslElD/RK+mtYQyCnp4TX5tsApLj
9yNIi5lvuJ9DhVddYt1K42TsnbLbrH89JskNIpbhQRGiomLYzrc17P36w8dDG3t/OJ9m5+agMeEp
FfHZ4Cx1Z0PQrlm7AbvcPuDcT8LSwJJoSrtIyPe8Zs1QyUWVEJbftVvQnrMqkToz23q4sU7tIbLW
HEpVj4Zsj0Ag55rVnksp1abNdrW7dJSO6R7q1heYHSX312Utw4ZY636zqtRk288zdvc9fnmZtlRi
UemxZd+mndZwolEsOh3fN8YHGgE5C97n9XciJr8Zq7yzuAPfRCSfsBD/X/hZj1dkmG6+g+31z4PD
5bKTFuNajmln3O7ptQGYUwZwrYVLp/eXurDbmIuWblk4Fhb+S2Grx/DhAnNA40atXg5frHiAdL/u
uZ59VUWrcStVNZRQTk/aom2X2hGDjkGsdj35n4600zTnBFXo8AupjkDNgZkuToqEiPWwlGxrJ5sq
kpXQcnNZTnB7ZObDlGAMhtu/MEMIWYulQ+kVs0avJL1QpGcLGHS6b//sJ4QDX6TXu5l8s7yduizU
MBaSMLX567P9icXwOv3YvsKeHP9LOXE+We2q4Kr7GsE7lyPfQN77M68YatGLA3OW2cbMSYIRIRT2
0UCYNRERe2aGpPlhh/k4JBsJ3zDf3zh9svXKD5eSB5GUMCzmMZgtlRkpuP+/Gg0MRl5OvEwW9P8s
1Gt1N+4YSLyO5ZctJd7hQzaL8VWpzIqy0oluwiUqfnjYTRf5S6PX6q1AxLDkW4Pe3CPiHlLTGfHc
FlpPR1A1+auZC9Y7nChhXhuaTv4Esax2dbvk3T4/jwWKfXPSvWOQifLOoijFXIAckuehZoZYRrHQ
WQkt2GSZiSi/hIPXJ2tjwu1Pxbq5G/jTTpsiUyd1mo0RF3KcMN3pYwyXPyQFWiyn/9qCZcMES7Er
pDwfXINeUbrOnCxJ9BCTyRmuYKspXC31ooaQkqt7yFNr4QirymVagzHOXobocc2AOZEuFcWiW7Cu
GzaolcMISezmdRixowezZ1Ch4wUq8b5N/4teCqC2X4yQznJwy+f1kuAD+s+8NqnpBsXz9KKpTk61
mG2dRMmzFADEtjhwbb43QBKVhcSiJfPSfJ4vJzTLWLVUz+RCQPeokwyTPj3mtQOobzjXakdxqL0T
MFkc3W5yQd53xTObUe2eX/WZQjrCH7FiApwteYaMToJ/2e2zUhOynH4l70rJoxtFapiMfnrJd3SE
ayGM3zkupGuWv2ilxXE5SPdO1G5MbetwkNtNiZuBOobp0AP+L79EGOHHnA8Iu4aEhnleOMyAyUQT
oEdU70/W8a9uifYi04HNMwYEz8+vZk/LnLcvJlRRuDEQYPZWd0H1A8tAnO+XU1s5XJgVY3GHlzbS
oCYoRiJ4VD5juyalSTtxZusN5PkTlDsvFyEvbtgHvxtjrltAiteznEpOtLmltN/QkmOX8sQvlyOu
/AW0x06pNdSguJ/JBqK/zV5g4MTjp+VKHdwNqYqY/CZY1dairCOQKOwJEIuJov4lay0os6DX1KT3
9CvPvr96ylmbHQ7/D8ANg7bInySejvYlfNFLoEMDBvKOM91iNxeLdToXb4inD5lHUhDcLg1GriiW
TQ8tWV/YS5+3ggTUQdmvTSFaCLeOY2pcren6Qq7GU7VyyUXcE5HM1oM3Ix7vkZ2Rna/le8bW3sIz
R/fE1Y2dFkNYZA+zwrar1bBBRXTIQoHTiEy9UIMsClLRRk97lMPiWsTssJBfVySWIFnD0QIlf8Qy
8wJM0Jwm7ttXpEKII6/B4vEgEB3z82HdizC1TDuoy4ATg03tIM13/09VYF2cl6BZXbc1yjUuOoHD
QTsGwSotb08f4xxp03NP5Mb2mPbuZqa0tx/dMOiWon+rGo7orMbyFSHTcZ3MX80mTuFxW7QiQCki
lUmjIna1X/5vG4K4fiXvVbI8Ky8SmZ2lPcHPA7AoUUR8EmlXp3U4zQ+cF87qefNFVOo32EpcqO/l
YyGf/NoIHovv3XWj5VREO9MAI2frgWNuNbam1h0UMoVkBWUZwcQiZ7nEW/czwNJO7cQY+6eJ/efm
QQydfOXj/xDIiW+7n12y5IYHFH/zo+suKOS3v9e8ARAEJvJSNgs86VNa9+98bSYbzglLT4I7HeyY
d+teWsuxaNRefQl2bhSqLJQGSIULH+lP53EWNOQjRYkSLaiyv6ShADgqXhSyB37Xxw1JhbPV/5nb
NB9+3KUeXhNnfW78saxJ0mpI2Ueipqm00+Au53GkFxCuAaF1DEgvBAK8Tq52NaRWw02TI96GQUdr
210yrHCY0VGUFReXQwh95XaLb7CdC6V1FBIlxMag5EoVCteMlg8CezMOR/laN2okqb8ReOh6XZ88
K7c6NOT/KC1VWreM27mzHopj8tLgEk6IU8/y3qz4SBA6LWiyUI5zrNl9xuTGps26BBvPaHFLGLKx
/4NPISgl9JMMASYa+xdB+NyeYiGWDXb5gOnzyBf/RKghhcj8LTZaFewtLzbhPWbPSwoLvW/f3un6
7SaWdHMWPyTBEe3fjTKYBzuP6EI8uHScr9uZ1XfZJIOr/0Wj5HUH/nCZzhZ508tkLMsYX7Rf2T3P
DoT0mAc/ZcVH5n+OFuEE8qd5aEIolaKRjRztNcPD8lAV92uxl6QvqA7jlCzAAHwHyeX/vlAm5Hkz
FK3/HAWyB12K8R5U2jXn0nlogNrnG98k9NEQRMW/x218SVthtw+TFTkkIL0ZBQn3tmOWskrh/v+V
VX87xT+4ZSabvIAU9oILCakSrUYkXlmc0sfK1kktvJeglycgnasfm69gNZRG6Z6+TrFi7jO5mwkC
hphLPkPZubP22c0PfGWLSDJYVu+QsKYja5HdUW6FoGO+oBnpUmRCpjJU7AltptpeUW6QjoHT3oX5
EiHf1L+O0Q4XKTZDQUoKO1hPV7bV3NSd6pHupHbIn1hZIzxTykBlcE6QLxvMcBFok7xuuE+1L8XG
E9QT6wkD608S/dFRkKgvDqfAGUXl6Y4R9kBEfPbtDMQSxjtkwZmszIOkzyFakT2tROQPGC51NVan
qbIQ/0fXot+jeNxaUt+yLKiI0CoXYIOuMTwMsK9vnqJcSkriEdHKd45I0MkdWB2ZxxqvokkhLc/U
wi2MQVs80mrx1tIHNYVFWSmJtwtNkkPr0Sw493IZNXIbRPlRzx7eiDq9pYrUDh/vcbOIDXfOuIfF
SMimSyiq7vASB1aj5tqpmg6ZBOOZ1z0nhEGpL9+uFMX72knpS0NPtzbDBIhyVaafZBETGttKV8JM
U8RmA/Z1VBv4jHIGGwJScxabA49W3BZr4yRnDnrZSEFYP9r8Q2lDTDZAcBPVj3+pHMfeW02A4kS2
vZPqcW53gvV64+wfhGnXMCTe3T6aPFCA2lt67Zcc5+bwi1rV+YyOkgGVmkjaFz5uXZR1VMGIue5J
5XtE+gfVbYU/X5j15m2trJInEFaTOypxpvhrl6OM4O9idxU+sI2f+W1TQV4whGj4+qL3fNzaKNMe
i/uYAX6onhhVwBszLCKn8tixXzqhaeHqaX1kRxozVE39o3fcgOjYprqupGU7oVbFMSP2LMIHD7/f
XTY0WYNy//6+XJLzOkszAzR1HUXlrUR/IlMpdHpJlAxD4YEslxiE63g4ug/Z2fdT4lImWWZhn+5V
tsf+T4aLlAZmJIBgtTrNpa5wEUmE+9OR1SXQmFglHCJCYIgYDSHLrbDNhwdeDyY5vMnnOQC3Bu7z
kGvf8q7FYvKDvLRtEwTkSJqjGafB7myW+/ihgenOa3lS2W0z4qlAn6vS90G6Ip1n/MJLY9EI+rtx
/n2/+5XIfperJK5aP8oIc0Ppr/GJaG7etQ1hjbfTyMu7UOMTv0uIi/asmc4oGc9CFnPVb5O+3+CG
R+D5H1cmGrPSj/+IHyKuoIbZSB9WLmhRNpu5CA4EKXVKIwprhDlI6jnezPLDyB4c3PVUWGzDiW5E
G+Rwpei4cMX9NUjVy8IEGx8ctQzkg6jEf4BM2CuRZATwX22Sm8OJmAMGkVeGgu6d2UK/v7p/1HsB
KjIGi4q0UxUcc7PteFSxNSKrZa9xjorD4EfygcyjryRK6t6vMHUhWGyE7U+AFSSgUas6W+d1epjt
dEqTeKjFbgMe4CsDrp7YGFYEpVXGdzDZVszk6Z8yVz0FuKWiCCdpPAzb1eUwGfZ9wlvODM47s458
yPqAo5EKzCoKJXJD04dVbl/2eQZ14N9vaMRipkzbRbjN5IkIpJbC2l3I0+Y/RFPDHF1QUuiFt3Ry
4D64rKw1xXzrQBvu8M2O0WASxL2DnzqnrT8n31nMVWOrbeZ2hnxnGWiKSaYZvF1ci9lOQhiF52aJ
uJ1+y2pZ4yzEIFeSxGyHC/Dn8jpnYCHn84NAukIbaqFKEBHpkAap8CH2dFxqqCe8iXpturVw6d3J
XM2wuHve9kt0+2S2BR8M4eUXcgVoK50TRWbJJam+xBJKieSBICM7zBSyrfnEut/i0iRxyznTh0vs
tWiKm6kWNSMSMkHIf5yvVU3K8DyMzNwcK8U7kz/TjggYFazPlZZR1NTthPhjrHmvDS+UVsRoUGAt
NhyGK350N/IO6eaYQUTOBxwW364TPclKYf34TZw20cb3e9gUOV1w/vXGhG629a77RolKBYDVtFah
zJAdugbQHOn/ny8PPFyIiaCEEE+oToW5TgWQcHmES/qma1PyHhoh5HHhyQBAKBLKNVqSsZ0cYHEY
NgH8LZ82mV1dSvJcjsswT/kfsl9q20nr0Bie5QbOtsziso0kLwPvVNTT6LAyw/o7sRcv0BoiBtFd
uIGfTgGU/4BLk9mV746Rz+tTieDTkDVlwBBZPS16Tzb2CDCSw8Enaaym91Kz5upCZFn33TwbgP6a
WHgrb8o9NgPrrw3+MA7Ta3Q+9HUx8sBv4f4CqGYZ40Q9IASQ4/UauQh+0BJR4QjxCE1ALE1wHc4C
WxWtxhtTyNBAqQrnOQ5eGOZAda8O4E9HJAZ3VaC0ExuE0H36s1pSl1iDxaptYf9hULU+KoBJ6Xx/
XGqR6xfr23OKwfzVoaOqV65tX8FQ8yOAGmK7o+RnUAJpPBa/HbS55I2lX/sXJSvWgHiOc0d770jS
CAKXTQmJaFPoOaJHV9Y1hwOmtHPhrwtpB5vqLmuNdxyu05Ue7DwkuRd5qc3thqvU1neV44ldUR3l
zPysr+sV8OdXdM8XY/4TBkN8tO/JMIFeLEC1YMoWG/6SRNtJytNuCB5DbMHONOJA4DUXw3SIft6S
3xjitpfBB1XmQPHjJPwJgvmHRdMWY4ceocL4a+uLhhtjcjIVL/mCoxtVbydZhM24W6lQQPwgfgpj
b40MgBnYufWH0fZ7tAYK5oI3xmNUIuE5lSmgl/6QbUrvQmvj7U2xmbPUDeUlbN331V/OpY/cxztZ
ktR8rG2oENoP+4YFwdecoJFa/6I7WtSwKakB7z/JLYgJJNM/kOXJ82H626BB+BVtBd1s9bRFDnUu
pfuJWNIicsSoCtzX55CAlb9NSdgUth5QqFmgTFyJnLhuaX7ALfN7LGeA61hYySyjQzr3B2YDSVHq
JRIbcZqw6Q7UUyFMamnB4VVZe8CBFT20aLM4zGacD2a7zV5wjSqUc0wh9veEugl/6VRjQkpnG+42
gS0/GHrcJrLAzx+ISTHNt8PQ0yRtTIS0tIlbufXULw3WBjg4f59SOlWXSAsTj5LWk8Hkf1tOiv4Q
/J3G2fuadsh0cNvJD0V99tVRCZx5GR8ZtD/I+f66XcsGyO6krLHx2s9I3CjqD8KnJzm6r2lEZFU+
+iFC6ylHEzZDRfGKZEXm4A40QqknRdhdkT3yhVRfYGzAdVuDVk81a4oebkOhsq2xu9J3tRCYZ06c
siyvgjATOcM1nRz1MtUnp/H8VNafKWP7cEZVRWSzdfTUckTt/USCgu2JPrj7e29AOhdmvSv+1JBD
TX0Sx/CEpHAXPMhvYo9w7AAHI+FqCyV0Vj3QltK8et79zMlsrYEu93Wmtld3SvztWOGz002u3G3P
8GHhAoDF2rbjl9qWMbSMLlGF0jQ4RPRBAd7AE7WC8spRJwzO5PHu0S0L5AwrpmoauXsLpPbW+D13
fZ3yblvMvsbicLc7xxP5dQCAOh6O9+8gFrdedKRighx1GtsmbMMKgmVNhVV7XB4aEC99MtGU0RXZ
XrK19nPQd445nSBwQqqK+Z1A2hRPM/kzox2nWmnpBfDkhI7SJfxeLEJlJZeshsFegQbzU8wMs51B
mrM+IbWjmpQyp9bswkahDaeMbNmeD/Lk2Yhd2tV8lxuPyqzp1UZqXhrQTAR7Hp/lh4pGbshEe2gB
Eog8Zo4MN6v6VEQPoWYyBtQiZIskTQm8Yq8SEF7AkgGAFYX6pEyY94y1NXrE9gKOnR6NiZIe/Zxy
4ddt4YOYEhqbry18qlw6b1gJyk9KOs7+a9B7JCFL7yfXSsrNqHB8cOqW6jSUphMituWV/chJEOTk
8D7arn+jHBjLxJqOapu7prK4P8UOmQxvEwjcyrCS4xHDlNryP9buBngV2nJBDvaIZgHr9dXwAX89
EhkfC4amPaR4R+2rbo8Uol0cmGc2uJB87OFfWC4DKNa8EpOtR1+BIwOY+rUNqkUpueku9HCYrhIW
yyZb2M8Qdxgrp6SRj1hKHy+vxe1wQu4CZPpJBuEWCPJW2er4tHYWiLoh2jyQzGXzKeQy4cUhQXWr
+kzhHpjnOGnF7/cFG4x3Dj7IzOR3XJjdRTm7fLsHJ4186/o6cMr+/HIk0uggraJNOCZnN0UOaeUv
KAPfp0eA0prc3C/0HEZxJaVgdS1NwmwrjAPYd4+n4XUGCHpRhsSK9jS01fEYzF1BgbN8pYqK4DxU
pGO6+/YXjwEIFWWP2nefEHlqmcIq8Hn0Ff2/FiRORPa6YjN3R7Xo73yNBnb4DS1Qa+XQ+WHRZHeC
kW1oiovmesTeSM8Dpposuk+h47d5Hrr6U7wDKd2PZaiivYuCMfuJRGtfLpDOBNUwX3dBjw31sdP4
lBwtBZvcA45gUQ8PN36Ne+/ElTx2qLgw/c5DHWuW638ohXgc88JoIW/VnaCK1iZp2Tn6pZhqvQV/
aN1SiwmfYY0NlAh5dcV2B2dtiq+ToNEJGom9wzzHJLI0kGE8GgVknhHibO1qF2qTPjRORF1meC1S
tbH+brSqkx7kLPLtw61yNHncDFuvykcEUnGBC2EdE4a7aoFvlkzGIwd78+JHgi9Pxwy85sWeSqxD
G/iWdXbffzuhrZMj86/Wvbl4Me9O3T/pip02Y2OpPKu/HrZ9s0vjtX9AJuigYJJ8r//fgbkW8RWk
ULwdC/glBDfzH65uPLWBBvfS1onMh4Gv3ZLx9EVIo/GrvGT4ID+z1bjsJuWMM6cdWs0XxpsmC6Jq
4XP97y7YV7R3i11rJlk9fP5I1lSc5PTNbrhED3kKgAIos5JZV2HXHwQlxQWl9IpmRzd+/H7d87Cp
bwZ1v7g2+5C/uiwZaiYEbWDylN6F17Cdo8k6HuVZCOjn1QZJ7PiTbhoq+1a0NDPLScb1ElCBFBgC
87SzpFVox8X5Tg3uNs1Ycmet4M6S51SmiBPbDD7NoSRXDZM43zAJrtCyT2jTs7/CTfMQp8bys+wS
4eBTgzfdG7hA/BUcl0f2QInLVnIFsYmX7247w0m5UcECYyQmjWoCt5Tb7iTyxWqD3d/qa11i5iPe
O9xE7Lch9shSjbmTzXbgpecCaJkKDsV7sEJL2U+HngAnkrReyySOLEOkTiiBH/yYvo0L7jtrVyjP
CplCJbxLsMhY3KVNmGFP4GCJ46cqbBCUWPANMy3WqwSJtf2sF747jEtMqvxCaANU1+BrkhMdcTPg
Kg3xAa667gP6IsMob7N+dOmE0C5zKktxUuQ++y4mw41YjOzZTVKDzxq8gghJW7Wg00e3mW2wYqUS
xK0gNFI3HqIa2XVBKHBpRhJgm2rBlltqB6J+9ka9QEXZu6+YXmTWDa9XycKKMpOwebKPL8QDMCRJ
yvB6tUbAPuUsDptyC7IPYO+4loZbEYkq3KG11bR+qx2aQFblxhQS4gTBEu2T4AujQkZmU59ojtpw
LH3yhZTs47yio00jFKOP4t/Fr8AYfiWmiUdqc5FNlI8Chet21aIKRC6wsR/OQfdk6yzzcCv6cZPA
PgxnMb2c2yK0na5ZZ9V3CPIQZN8+w+Hx89l8AeKt4f+RgCIaMJnzEg1MgrGd4Co9YTbnPGoP4NV2
Q+4PyVtEbiPSgO/4zkKl06WZZvKTrXy6DthnpfU1MISG/eetXSU41/GKKrt/cy3KhZRV+5d89kKP
LJRZIUXdtoJuromQdwqTj98y9CpXZeFuuakNUsYaRYCGXmY4zZbdamGjkW7fr620dfg12uyPL6pS
QIW03gOChZvt8pQNUW1tMnHp83xz+R+b3dZ9WqY1IILJJclI2umJFtlqICN0DCqB5dfq9lQIZEl1
kdEP7rR9uio8oGyj51+L0bM/N3orJP09DHVD1pol6Zd/r2NiMyGidl05n08tTmjxCVmo4EUyI8VB
tNeiyhCNrCe7tj1bFNm6XSH4r0/QGCKZ4h+r/5bENNJIpiAmXzNajJVYpMCZTyvUiU/FOlqOeNDF
vveLgS+tP87wGL6AT+gGHItVhgnrjOmQrMdaCf/t2AItsasstEt48LocmG+ZnNJ8TzkLtlBLTyhQ
Q/NVqdRHNPaEGbdD2pztLgG9EoHHaz638H8xbC+PWhyjYLNFesWPVjjlw28ktk4sSCoCiBm8wdLR
M3toOw==
`protect end_protected
