-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2YA7kOVJ5Z410HYMsLMOtIKHo88g2nL5EB6qACuMny7UkqCF6xWiz2UApg9E+cKQ
sL26nVvc4/U3dWpz0/8fe4LTZG6VFRdjPcIDV3Ni1/68lVCChlSWV4DMVRk7hW3A
PcjuxYyHqlUUhSZVGMoBxiuHCZGu+BjWbbtVKbrnfJU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10320)
`protect data_block
8Bnw2CjcHsdDYLD+5bzjm5m1vM193LJwPVQeTzpMdXMJIlBpU2MpaobzCLMBV8wy
NEPrSvpglGfvoe7+4lroQyeh/e6yhZb0xfxiFWLUh4/36CE9La6dj8lCpWQ6tK4A
4BliFTVh2fuq5/+kV33T1uyx58ksTMuSUY5fn3TH5ry3oxbai2CL3hmoxVy+o5X7
OhksmaY1OrzeFy5bOT9AG34E8n+rG2np9OOCvLuiZmmsn4Fb+Mvlts0MIP4pSM1n
5TNqGKhgryKbI2PbtInpRDP55g5Mb+BFkPZBh1EgADM5EW9a0Iv/KCwYQ6Js2obv
WQDPWysE/t0eAWRYSvJzqhQTLJ7Odc+DAQjmE1Xy3F2UTrl5x1jJZG8VaJVG0vcz
MI8yDKLh6M7MGLnJYIn/u1zXfWwQYXCA8xEzfrTMgJJ5Nd+Ql+lAVWLfrDEHhBfD
1Ium+67LuBI24Ju72ijxfOC2QiQ6wjIaiI26EUVV0JsXv8RuTdnguMZOacru2RqY
Y/kr7bJCm6qRvUd6J2W3vp27w0Wlgi0HidySS4HlQibg1LTRgs3NEtVevfh6xTG7
T9GDHF3ritCIvDJ4elpHij11cwjbxmyjUfp5PfEgftjHIuy9NGRjB7SckwUFR7cp
R1ddnxS9qUeCkyMaFAT5ciymWAhsX1GUnCtqORGpuH4Q/PdbT6lXIuHyB3c/g2N/
bcX8IVeOwziksj5Qp9FS1qMDnlECPl5s3Zd5aKm5NJ8Rl5vUeuRgXZ3tCiYC7cND
bZEAj00bQ6pwlyyxGjHEXkp+Qf5SrsFgsKALNo33rrmUqGpbVVZ5DFxRPNH58iEy
xJTRcIBWf+XGkAF/ecwhoLm8yV2WytnOdQQmz2e7TTF7v6D9AHrwbc8CN5ysw1X5
QJgxrabRlgZXMgxuufcLzjCcfh5hB3/1e83dR+/rZarpzwEBPpeJSfyKDfBvzRB7
8A1Fzkhameire7Gi4pHBprjh0w3NiHLor4l+8uj0kspHlndYGe0E4onjk2HGOoj8
YkdbzzdbvZgiYfdj8n42dG2cRE3OJbCWiG8XPZ6JeNGVQ5oEfs5FDOwAJcsYIa5p
MjH9bYIHnh3BJwRJ/mP3OGYvu6UkfNRW1nOTVExdqNZ99hvhfKCf9yTreyaKh4f6
Re8PjO4qztp/drSD3l3RBug51GN2kMm7qYufUILD6OO4E+KgeE0MptS/3qJ/9ULG
D75UjMuKNP4a6xkD7SbcU2PiGEsoipjcIyQMqS2HEOvKd/Aw2FhHDu/kym2zWgsw
f6LD3iXarYSiLlCJbZi1I0NIq2tt59xesQ3OeD4jHwtrlym/0aI/mi1i3nrSde0K
XJ3f0h5Xb1wxQ1IH1GQ++LYEeWZAplDtXmyxkMf5maUS3NAB/WbE3lrID1ZX9Gdd
rDe/UWXjxy2mizcs0Q1HvetFfppCs04Z8DJ9jAI2WOV8ozn/oPSBfA/r1NEQNXGf
1GE1BqAylRiUXTBIY0+W8Kemx1jOs5/Xycaaady6/Qe/hr/d4KBGRTA719BxeTU/
CMQ8+SJUbDahTimD9sEBfTbLbF+a5/MxBM4lfH9XpzDG+1rTNTNSycZoL15OGUMl
JwkNuXnKlGA0e3dAfc4l2Egh2xCN6VYCBCoITP6GtSgzegT3fplXi5rgaK8JdVut
KFoxPwFXnUeabaZv6cWLM/b9sFjQsZGF20mrkmkd4Xmz8B+EhgQHREqko/mRTDDe
Ay2L40Nd0GzuDeHJau94vUifYzWYI0v4cVbnfpzQLrK27HTfL6Iz5n/JfyPdVDwZ
Q8rAU8xSLuPjYJ4/jA0TYewvu/2kysyortgLO4uDW/Wrl+KbCzFWi116VZQdOm5j
X+YC6+oACFTveVF7XVsyV1zrEvj2tfVUQhh9TTitp/ojNoS6DrGP9KDuq/BxlgHi
toqPhLFjh0HHuACYLZxVZeox37xse0Wo6IGpfDPGNzyxlOz1ZZd+IpDvJPtAHJtX
8QX1w/XN+vBdSw3rT4QtyF4YHSK9QTftrmfyKguzC5zj00Mq2veodGBWIefPnbqt
WjquI/gAhoypoUKlbXu5vGUf/NFzj7iJCgWlYLe1xEIsRScA4p0R2JPOUZOVRr4B
aKSYO/0YJI2Le12tnAYASi4dBLZGReyuQFn96EfnwVq2tHzIt1vw33C/vUyqyDEL
1jc3/IUt3OTHnU8dHEuylbSnua/PosNCXmVFYwori1qBM79YKQYn0NgHzGr+33yQ
PeTUqyNfNufkDO71p83InJlx1fIATWt5CdZWIsuKGc/3l5xhp1BD0E4h9/p+yLbo
ILkORuKVm7GeG7QEwGOsoU7ZTR/Ak0Y0z4SswXtWj3aIseOCXQjcHt/GTGPWwRBd
wn5LzL9up2oAMHwe5fxOLFHZFIa4RFtfru0Jx2FRPc55BbevZZsyx6RVcBLRVxqJ
++Kkm+2YplqvAmDTg87pmRaImxOozCXdQo8QZCk3k00V3a1mpeCIuzqKmYR6p1OT
4qomGU8YvuNFoQKcJeXgrpb7XqJI5+C1OUxmD+74OXoEAEKx7XoC2Dbrrs0g8b/S
ZAer3yx94ML53Wiog5/oX27WM+c4+U4lEtRPBNyTJbx7q4v5xUAt4XLe2t4uar+p
5QfkyIEa57cLlmFwv2a2PlYQW8mHNYyOmQfxRwtFAV8YsJlWMPzXWLra8J4fMcaS
oIXQQKzzR62xN9ErpaAKPCt0XNpVc5EvqVcIUitaofwUJ4hMtrcimqkpq332Xu2q
Eg1+bG0VFNvMrscSBmWmuH1T9du0PfaA5Q3KxKta7RSYYdGhigpOiJ58sX/XQECj
17AZfqifn9s+TVhbcg4gNFmCW6ynjsPt2g5rkWeaPSHcEMnNT68uU9G4kLSDmfH3
XgAuxz7G0CBgCTAKrm/8zn6xdLavmWhg33x6ldG+Zl4F+oCcRUcJnY1f7cjOxfiO
6I/uj3/ROI5kbihLJuPyoq7rl/Y9UBR/JT3kuIZSPbFQ2mcC9pP4yh/1FeoKOz+w
ptrjkxN/wlB4p6oX0FmvwNWS9bno+meRRhNn1NdLKm7uNbPtmVYml8jatj3iBxgT
ILHV/XuaUF7XG/R3JhML8X4yZIZJ8pMV4WHD/0nNncMtDtDo6ggD3alx+bI6GoHV
GCHamgsRg8vEQtTEJi9/Co4UEWAcQgevfrifO0wrS2hZKBUdz+X80LtJS2KcXTrn
J9hvPHkD5umMOi2dQIA8dlxsZgcJGNFZDywjF20FPiKAKABUAR6VV0ujvnSVEMu3
cejHWldbPd8QqjQxJYnhKqnLe94bWnwQTHpevtAZkc8oeh9NeOawjZ8/Mw3UTadd
V+TSTE0rB4piEW5wyD8LE+D0QCkGnw2ckVXpP5BrxYZHEER4sWyjCfzgTDVtNvyK
X70kjeCFCHeo0DEqyxXhmZz25AtgH1YR4jTFPCDWQB3u3gej0BWZS4/GHPwIOBXm
0D/ycWovENtaYq8eVk8VWzs5ruDI8fhLqbLuNw1K43ODgacHvU4ju43GMWJfW2Kk
ZwcKF31XD9c47GThUj2O8t2caTnNhVxKNqfm7mVhJZqUEAe7cISpga6tuc8PXgAJ
hSAAdpfxtNSINlhn7z20HScwm6obtvOZEydC0CHgKrCIkdA9D2j09B2BN1FvRkZ7
dfMW8/wFSiUE4kyqQqJHLL5IgaDy/tPEfXToEveZyUVZZeoy4wZlavfqkgx5hwa/
I4BRT3iJvWV9w1C39H4yaoU40instmfllUk9Zwv7Jb+xVNIveNCIubH5dhWvg+Yq
6vfqaMz5ISEl1QVLV7bkmPkR2iGiaSYQSaOa0G2Uv8AGwNWKakMqoih/+upJp+v5
f1vnycAgAUu1IAYLTTN1k4ZNjuQBcD4X7pySI60tzeda7WIvIXBn9UgXwsgdck+o
2TBJuQqY2kJ0l9TIVkttn5AZ/Zyk43NtrBB3uE3oderYOULpw46zTkxMWZxCyIc9
wht3iON6LkZVLchOaSFQbKE4QPrKiVntnZMk991SDlDmBrnbPJ8YzVOb29SAeBLi
46gAjYBelyThaYiMKIHPxiVkaX+O2OB//saWuTUwoYV3WO5NrEvVKtfkGNm05gRs
9Luvqgnz1rK0LwIOq19CpPzQ4wqNV18KflCIaYn92hoe4jwRXx8FzP1UKNUWNw0l
2qiFGakoo9wPT3FN+k0AyfaUKwDlR8AmRluvrBkk0wl975B0sFpMGDBoV8layoBa
JZK2B+AjROMq2DSuLbAmR8+AR8RR5KhtcxgPW/PK6Fb3goNeO/fQzEZAivA8x5+o
d0UOg7STgEuWQLgtdguKiZodyVIhN/okp6a41ErLyFGiFS/Z6aJP8S1G7+mYUJLb
qdXgYT9QqZm02hhXM+SKdaBQMDck3fWsZZioQCaZRekWFa+EAULMYFgoYdxAvxag
YtUQa5UBFjoP+ivoJ2CiyXT9rljDJuWThaV5N1BoORoXQg3c1kqpYeaeJuTl9Ovi
aj/gIAHlKNid+6kMf3VbIeaQEsUbf9rN3nh2+wepjKOEI/GszzH/gxjVHsBGyx+E
/c6eCIndSbBThLCy9Li3MMfBJXTVc1FN/Kh7gNXRZC4y71EuG1Ik9QjqZMCSpmZv
9DAgIlsEcHx7ZRtjnfs4sVKaKJLlR6iaKVxTBkrxcbIUcRKmF11bqo4WxswpEDge
s3lt7fuOpOiuMwJD1BC3ZD3PEAXm7WqNd4gEbhOZO3eSW+/AmnD8MJy5JwQm9dop
hnGDb8jTZZmaPuIcwPWbJc4tqctbIdYvl9Napn8VtDzg18HQdexF7BWJhQJqQY/j
XjunwBO4XA5/xDV+bDHv6+o7LI6lo0Wm+dhouKbvG4qDrsJmIhbPc7Le5kTdGw4s
yqWR9MJZxCE92+f876kZ+0maaVTEw7HXq3/HcVdDR/usjTLjcnaqAncqWsVy2l0N
Ms11BNTnZJvhnDTnTgNJ+Avcupe1tlN704zyZcNTFcR0+6/3jgUd4aXl/Cn42ZqY
7nbaMZmdzMAzePCvrp2mOiOvIJH4Tba2IRWjSZ9SOfuEaYOb0XtR5tMuelG0Vg2q
x025tpwdQrwIm1MTZGhUZXpbLr+b+hv2nrggMihsfdKf8xpD0iTRqFQkCsW6AxiF
5bF+pn2KxwWF8jtJI3g2/jxN/ghcPmtx2tNjgCRIfmzS4xRWJM4w4RirIpx4rgHb
1o3ztR9V/XOKVpDZzbMNdgvc2GfrNCZYc92pbmGdVpEStGcufDhVuZs/xoW27Sal
/dfOTuASWfwNaIkCHan7uRaCsn424KwkWxntcqTePtE+7t5qSk7fQ9K2oE0UkH4F
qreGMy4MYnN3ntnhPrSrkVk3G6r55VFP/zrvFGUpUm/LL1r7p61lNIl3SWnXBxDU
jR9xdSp3mEokhuch6YFZhEge6Shaa9cw35P90vAKJ6hFafx2kSwxjoM6NO1NH8rD
E2zsgguga1EUoivDZ7l74SRYemWHIFSozKg0x7s6yVLWgcbEIY7vXbwytkpNRgVH
QqlaLIuZ6P6CtHpFAUf3ZLA01VY1zQqCN135G14ZgKCpMpDIMVegD1Z4tmo2LcXn
ytwv2+JoPyG9cKqOALz8q8PN98thK8aANwqFe/+ou452LEVQCoVygpRmCW9vLRSQ
KKyAnpJAs0Lm5OdZoPEErzaXLCF32YrI9yCKgR88uiai9DHX9Cid8KPYiP3qRRHj
GZJvsYcwRNKAmurMk940e5pVrX6DvAsyXgSXZbNY7SuYqo3wX6nSOfBPmjoYvHng
G8iyw87FwFuEoC1JrZ04T5EeDqVc87NG/kju0bWTUrZ6L2fU9A1EMZZtmXe6S4NQ
U4RcXmTCSDkjCvwW1OF8boxTgg6n5XNxdfMXtdxV22Xk9VzssLwSm4pfWt0szu5a
aKOewzgeqJhGKUw+9pZJhODhiC2Ft/kUbt0fmmViC48mItCN/XrAcGBWDdK5LCgq
K7494gJkkATRLvn/YYqMPImoQSp62bR7bjTkyHWPeyI+JdvTsP3XD7RtRho3vKmz
AnnlADt1VJt05TldvkRz1LKcUaBU/Ijlcg/UPy2+NxknBQostpZm0H8H3XkgjMOJ
FJKE1EM4dydErZeQaZ9FaMXISAWDw3TTdFiiMjm2Qel5Z8+0vn3JYA1lkgsOnwDx
CRoiF4NdfX2A9uG1j4EQWGkdhPf1Yt+d0E+uEFNE1ukVC0RHI7kdx3WKg69+mWd2
ZhSrUZLFSXZSGqufTx2cvBf2pA647ITIBmDdmsW2seZhF+qogcFoJBvD0/dDxC/8
ihGmlUDrCWEQfhyIW5kZMiJn+XeofUhLp8EbnBsKzEx+2CptOY8VAMd8geAcVR2c
Kn3tavQXI6W0QzD9jk2DQkgwKtXJng60fFKKIIQ7S+iJl35CdiNBOOJx8MIL4y/N
49sO+FzC7kjhoM0ab3zpD1xO6D8oCxYolw414PoVvz2KKDYCnbFLBhbn57DK8IdL
/Xs3U38InD1a57PhE5SW9fscVZhjpINoivGF/VQoWUzxlAABvhIt41saq/lbfLEn
mPcL/swnXXKncaWXaIdFIRRI8vzyJGN9ciRk/FGnDXooYVlrnKLvbh1J0qE5fToC
gJUCWfhNsD9r853Rx9UH0rR+WJh8Xx4WJiXfl1VXq+BhEEoHqGvWJ+Q3XWnpIO+m
v+71YPLJB5j05B6ReZHcvISTP6iP7y71piSTtq50/OFIaAcoFDhKjx0MW/pRVfya
pNsAleae9MPk0B6aQTEDjMO6tqS+gJxh0v+fRqxUJhfMMVWOkEZLF8oWc5XB3IT1
UQdhQx8oBsch+FXyYFULo+Tb1mvMJyTOcLSB0KBJzo10ohThmajqg+EzxUsQVG4B
uo67OzhRrfrlbfgBUgXYaegs1OgG0IYlYBHg34juekQZ+hGVp0tNI/e2sBihc5MW
K9fXQdc/5499ubCOZsxakct6YzKWUyE+m6b+gNsHZpIGVFy8NPGSlim0cEXOWjHm
q7fSSHF+PKeTSbakDjGErTP4kNdJbM2GvIOQlD/6pEzJDcWrwm37xIRExm0eJYOZ
5uE6n3gG7rb0Ptkb51L1Y2XBHlr6vtGxWtUgQwV3KQVg//kMhdk+buiNDQdjrWXT
oiud7Eidu8tjdwPxXXnKuFlWIFZEm9uDYPU+pkiLNuyUY9Xu60xMoBZGJx/3T8/g
sHmywrQvQGbJKdnujqvcdfp9078ik2WbhgJ+EaqwbfrOJxOsghH8+BgeaVXyo0K1
zUB4NupojiUdlprFs3WfuvHyl3ldcDV/MkAIDlEjrzWhFGZnPVCVHkOptniAZcEk
G0pjb5pt310TuUXPQtX5UV2fliy7yYcYwYwIgGEQhVLvRyL4ltLWzH8z+lEJsiuK
j0UT/ZRjBlGTOVu5LtHiRnIogZOUq5P8MGZWTSbAlF7EAaC+EDK2DUaOGSX6RSzf
b7Th9m0qTnryc9IChP+0OD4vnBAUp2uZGZnbhMiksdypKhbDPITnI39/LiJO8bBd
Q1szP04UNm1t90MfdaPnKT+XoH+AYjoHryHKMIBi38MVSvGf1O4rUpbE+WaQBj/P
W3gf4GQPsLvkFMe9zvIOubgE6QFS6OgwuS/3atlfVyIbvlynokpaFkx/Il8EeNLu
py9q0xqGU0y7U/aS1/A+BymbgjeVjdU1MYoOkvRYe9cm1c4L8zrHWyFuPj5LoQes
Onf/hLB0Q2tKVWGaRsgMa2KupipWU9hikCKm3rWKWBv8MDz5OTJYdYh0aQCXtcOw
HvZZK3GsqktSbAiAS8DbMcAGBJsvcckRf5C3p+ivJpD4rqSyaf6E++wON80q6cRx
rW31mX18j0ecvMQBdk9Ya0w/EzrdNRjBhpFoTRlhrapzenVgoesib9M7lYoLvxrG
Z1G4yEsZp9cJ43rquh+oNlPD1S133EqIHGMBQIn8i5/nl282/QP/1m4aDW6hIMvz
IIZlCVCXb5TR1w/JqTWxjnWbi8MJOAStnjd5mJo3THyep2VZdpQoR24rAuKNA9jZ
qGqpy936mCLDShI9td2lL+WS9qVok8M8DLGD6p38u9bjCVW9DfVIZegRdENj3yeM
YkgmaHs3rp0ZnVS+ohJQ6b5MNKLoshQ5a6Ohg2D8ORb5/y/Zf3HR1AVSdFZdfdxS
eW8H6GiaqzQfXz9hCr6bhLUe0Xx9bTATZx4KWX0V7z8pqbIHi/bN99XNAigDn0Hd
EmpxdY8af2pnQUPmv0j9uRXXgWll/7l9IHHFDkuoiWRxs0A1TuuBoW2dqcO/NdZs
LOR3sbdXdzWSvs2IUVZGzdkfNISF+2RaOvQP544RETSmnhQokGomoi403JCJQmqC
yu/HGkZJ3dq3yw5lCGLng0ebjhwsXUm9+JsirnTbvE5QjROUWCEqVfofw1vvM8oz
BNPIXb/VyTdAS1yJzB7YBF/jpaT3NmuUd1D4Eg+Fy/Evo9L9DzU6ibjsIa0ublYK
2OAbrDxAZWOPMj/hHxQnuN7xIoOTdrvvzdKzEf7cBfQgcdbep4VgFY9LwAmjVL4V
stUq0nHFaCJcUMV3BDDD3SvtaZzpqOiw71Y3aRsOwrutGgPoVrzEW+Cd8U1knLiU
AZpI/ea13gbeCgVxBrM9/WyLZhixdeWtx/ofnzD4ofDMad7ba04bgdXFc1LPwmQC
XhnmEQdYpi7RtPz7tcWzK/f+DSc0tbQ3oqKH2bEKYGL0TCpYPHrDZjvM5gXV9s2I
MzA7YMxLFZoJJzLgUUAI0qXl5AqP1wQGEtKFhCxsmnc45aVM3XjkRuHMT1Ojygim
ZfG5EshwCWd6jq9M1Z8imBYjN0kVj9a+6FWWxQydJp1dPDQ2AqRqtKVakXZM6pKw
ad4LQyzO8GCKAztw/sfdBhacLh/Iey+cnDrPX7NFFGXakZGaj+47spKi6SiDst8C
XxaFZvr/bw3Rh44fBZ1cRK5PncK2Cc+wTTT2BvWh3tlzquWasaEdOMKnFN40VBHf
4kzF2/qoeBZ6CsHnxDDJNSU4y0u5QQ7ZdeSMcBXig1xBdJeik/YHHIoSfVHLVTco
wNV3/PF01HUSh6FyF17a1RQkkYlJfqqqgy9ah6p9I/UXbn4qPu76Up5Bv3T2G9V6
tpvE9Jaic+37q3WSyfRhfwvzQsH2jTUC1NZ6sNscSbekjEelHLYsM8pM7jkIHaV0
qZznueFhdNQdyzmWVctQFpq4LCbYYGJhxJJL/lh9IUQFtIeRHKuSIb/zalSuKwYG
hAamTCFTERravHk5aszbvdZygT9+6DYSUgYJNHqS2qo2JiD4lGZVSEfRteB6SEbm
1A/EqlhuqSVM7hYvjZZ8ViShBCku6o2xzpJ1CJcBGJ/XU0AVFhmah0PmoJmWu5sc
VpnHhe6cG9ywSM8EjOGV7IhQ4SmINfiod2jRS8teTRK1pKjNT4aaH5Ugma3TTiMy
qI0OQHvE/5pQaynrldIU5yrykGdpuBVTsZ9oRfTT2KvOAIhkAVsEfGUxeIG8DPc+
I2iCEyhtR9YwOaQMiJhtgwjL9k+yBB+Ie0iILmMrvakMixSh4z94grIPB6x26LO1
odma7DaI0E4JBHixIPmTIQR8m4GOgzz7Wac3J57x1xDwDaN7j27CVRtR7IPtRNzY
Rvv8Rgs3FfpcIttRL9+/dGlaRqA8Qx0yrK71Vv1ATECujjVDn9kOGWWzySBfOUZS
eHDzfi/AyXoesN2ARHPvnktWjSQUtL93u9Hfw5JU8zv7ob8TClz72h3MEOY+lXoI
ZrS2Lv8mAYfF68WLF81u8U65qx9Bf5i5CdUcagHPyx/YgmAbKbSHyehuKyuMRs5W
/LEU4tHH4SMm4GgBanOegstppTE+/H0JjLatwW3CeghGQFdrXePs5g6VwH64YAs6
HN/Uoykvayfe8twR5Xer3omBVfFt/pxzwKtrThSQMJt48tug2O3EXfLxF/BwbkWj
k8EPDVN2v3hY65gno2pXuNzootLPJyXw95IgTdjk41mi0p8KrZ9D4toZosXGuhgL
gJUc/vUCXhV7U2hKg2Eyt2lKUYsAfUqwoYGkfYhu6vfj+pO4U7KO0iS3KAhxWNuX
Zhw5WWT11CSVARLmTEY6utf09vJ/J9kLoaLUhSNZdB1mMv9CKgWMMimo3LP472eQ
jb93i0NG+bae3cddqGmEOUJdzLo+QYGt4I1oguVR374DrSxa30+lPIslSPp19QnK
HAiCvTi4iqPqLUJ81eIZlADaFTQmIb3lQNBb12tCkWrSVBB70AJBgFbq8M8lvXdM
/hbBKbIYfj59h0e6/tyE36Rg5InUEa6jycKyFFY0oZF0+o8t+dSoi6mzmRq+KnqN
1jie4kDQqMVaUrR68obqFupRIrOpVTxSidYmiUhpWK1CwPKNb+mr5JGS3/n1afI0
2eCxKNPshysfaTLGeKNAjdO8swGa9IAuPb9AnaPWancywo70etQhlaIQVOP0YaNU
ZcbLVSJ+xAoVJQoWGOde+xKEhkyObFUOyM4ZD8N/234TxTfhHCrRpMn0RPrIxqtj
HLyRdL3RYb/VltKQ7dKttxUgkwn9Ls76RXgYlrRIZV4adxUHWz0Ha1Jv0/ExpDmj
zx8o9o1uhprSA0V7GhJmLmILr9MfIuMyzWeV7CUqX3n9U6US9pyXs0gdIv/MuBS0
9xXEu4fZU7hJw1t66MaSCrUrazUygfYOmUkrClKMngyQXj4fFC553xgeXt1R6paj
z1LbrQmoT7EZF+4nI6e0RCdhKmyMRvBjrmXHOyUlpL/QBTR5EHBe45WKKbUJAnjf
5jot3eeABoKa8kPE3WJzunG5Kd+SKrjHiM4AedBIIpBxfEzGskKLuW7vVbypvxvZ
VzZKsuUqC06oRjo1U/J2G4nw43SgjPYhJFeCD2TTod56eeLKeV/wit+SNzV3/ZhU
UyoCP1Lcli0Ak8NQUrKwN6JP4OxnTl2uV1dZzht2gWD6WChMZs7rVVutlIZ2XZ8U
AJYCEYZg/36V29AUyIWP1im1OoIAia0mtZpUwgrmwb9YPclo3Ob7cBj/DbYTngeT
OcoZqcFueHclbK8Sroy0PbNqrmiSNPSPm9qX8kYz6Ub+S/Om50IuZAdev12csj0v
3W9DiJ/4OjXuo2t/X0Mb1wBulvMN67I9q7eKGp7zwpwyPYS5dD9MEMpwD9V/RGId
AldB6R+p9J95w7mMyc3Vp/RpF2vxyOZTs4X13gMoUtG5kuDbrXtaveXbHWb1wPw1
WlB38noaLS3+QGWU31JUdH+PhUhaGVN9hGDOjDsa8icX2GPuBS1dy07SULSNGMSd
YvNXhErRaeVVXsC0SotR30vpXfA+g0OwqlHO72E02J1Qeu0smZNcITWOUxP+7eTj
X+awP6NxRWlPU+9zme3DNhSz15pgMWiUig/is0YIl6qDsRMC3RQQlIUoPdfJMJLZ
XyMM4II/hlTlrFGnDBiYsfUOv8W8ONdQw/NV6f2UfZMyjqDXeSw/UFWICX7pssUQ
1aIkB/ukKwgBEnInImNzNbJz0Af57+Hov37l5rWoXS2j7eTafOfIyOXl6xj9ILG0
ZWOufYCxLyTYFHOqytNZmy/Y7h4mzjmey5s2nbmD4FBBBkqhMcgtBgmVHWawlPYV
i2StJodFnNW2NJdlTeQh0nFvJcgpZiNDfpY4FmkslFuhTMRz7bwuJNWUxFdmEtWj
mhdGDTcXlKRLgKNfmpfFSNTy3p2YD5e49T3MLb7Uoiekth9iLVLQcL1Xhslv2BMc
0zvYG02knR0wnyN2+rY2wUdvORYASpT5JrvayZcVhUg4brBZRS91Ai/OaKnW/Ud7
kIrc3YU9wrVZN7JI9FZjqt4dHdhmEXJocemjzbLAYznbz7RzAuGw/aNDb2kEtFLn
drn/+IafKUm3IPed+fym37bvRej/mmjMonHPJHrpRmVfA1M86f7j5q22cBzAaDzT
LMoOL5BIlXKHRVHHcRBouOKvkq3qtHs2el9HG62ABWfu65E1VMj2yR5KVDhd03CU
1E92I80WBTbJMENQWLKzbjSBCJWIOD4zUA3Ga+luEvtHJiUn7tMIIqzA6PU9gi4v
9cPI2JjEopiwYZnFX2ckkFhfwfCBzXZZfwmcgKFiy8Iqv2PrcdIEdJzmJQNP6U56
sP4IBGcGAROhiq5A9pHMPwimtjVsmJiMUEk2cAo79Y2VeqgcjtC2z2DCSYjdGjUQ
hZC/GejGGgb97RGJGD/LQsz2uiwNlQmDijKQTF11qs9wPTiq4N2vl086B0KqZv2P
7fqVimkU0+enLq8ZkLqY9qrbwrbsOsbTk3TYgMzeZRoFehdcsqJV0YOvUicK38Ss
kXdS1djiJ1bQ51azuDwoiaXWvYAqMFZluEBs2ZjNyF+ZSovYlSTeOnxMt2qUQ3et
NX8O+uYEvHRmLgbQA1s2Clfjr02kHJvXAyElBlxICylMbNtxoxdkPa2hrAWd5XL8
fC942mphNpaQap0843naA45Ta6K4iwQijwK3nGBnkpBXEfqNKdKFcpnSE2x3codB
AYBiLhFpea2MTPR0K3oAWriswtZ9QVFhBnNxNJ8z6Zx6xqxck5I3jhtHsovs7ytP
ztvN00KPwtiMYw71NSo4r49XhlAWRXT3pAXVMdQK6Q+ZvlznvoeIZpzIWAVjdwkn
tnN1WA0gEubjm6gn81GgFlbkXnK3dqAC2W5daH5F7b+yEqc8KPgmyrBbIa3ewEhP
mdq8e313ZUD3voIVd2b+t5wSNThtIwELWK+H4eAxHkXXitDaza367qrUonNajaAp
eGJJwTReaAQ6Hp+TEz5XMht3R6+epU64H9G8BzOJUfFjHK/ZzXSjO1ePB6MsfByI
8OuVLSwzgsOZehwovpZEUsiXulxD11SkT0pAqf8T8/Yc+KFtJjTu/tNMV17DIZIw
qLyAZibqdNFmI8KXy3aDcIP1SLpIno6Rbze+seiNpg15h9Od36zV2QBRT53pBWBr
o6vG9q3dXy78AqdvtYZvDL9PXAmf32d9P6crSFY38nSRqh6Z3deiSJy4WIVLa9YO
lUUOqqDe6npgDs1Whd96hW0aSzCLN76tq52DA/O8cd0daIonE2ie82hudU3WYn9U
7f/zuZYY3wwmGWlVtTg924vDD0oKr1IezVSVzyei7CgrIe6hICmSd86WNlMChujS
6IL6W4Qc/xaQynTtasth2WN+bNdATPOEuqQ3OQoqxxY3ZSJxvoYWHFmpcg8beTJZ
/dLmzLy2BUrQJBJIClGNy/T9igRXabxgPwcy56QGKVE4Hr7H/fR1zBBibNvYPqoG
AW8/Z6I1+ljwnSmQOlLP+cyoANvNHAOhX1QjZg7QE58RwgLeXGBJzUww/HYiB53I
TW2RrB/xAatEKkhp6HVeKptlRVSVwyHI13pAWNGciISueTaMgJG0L3epLyrtuY5L
5CYHOpInwhHrAVo4DsfzP6r+KkE0kli9K5bnwub/79SeNt9s6Oh5mpGgQ25cNYbl
vBVQO4wCYK5ZdddzSyO0hBCOuWeectSL67dUJYjUYbQ4HWaV/jbNhn4hnyXM/XiY
jSDZYPQ8rHFbvcm5dYs3Lm1Oh4QWPy/XHt2dstk+1lTrLz+KE9cAcaIzxQ5snSlJ
fIwUaHAujbHxnbp3FSbHUl9x6jirNkcnoLQNj8XXr5qEK/5SWGsRCl7sBw3Ksxg0
5GU3eq2iC1b6i/Mg3F3U2uQ/LOK+gu8E2aUfVqboTaZVcA+fuj4o9eifWFksNDYz
XVidpLUw3qIufa0YXabedC7VTqslXi7Q6TgeCHKHb3VM8IUhnYCvV3/5CDSJv+le
`protect end_protected
