-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
NLLFxKrQwW0GMafAsRFbrv5+ykClVOQhjsOZTOoosqRBnK2ZOnbREYwhyHJAi8Xw
/TDhJceutFap0IOGMQErqrZiK3Yg6kk56fiTHOir/tyfQMguK/2c54g16i+9K6yn
KgUbHj6CJVTNtq9XX1EVOkOsf84Vj2dJO7Lf5z+7Lkg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10496)
`protect data_block
RX4lPeu80XF8FoWrc3nZeVRDaUxvuDUlzZUJe4miOsuC1hL+5GbnCQOoazLXW0vI
lGczJBhlz51Z6CN1L46XgOeupL9BNe078aClH4i76UrZx7RQoqUTa0BtrSVmCgeE
vC/k4oAoXvxxrjUKj/d6Nn7S9TWhcmYnDJCwgujOa8QHI0k8UDqHnqoXBBB7OVsy
k/P45BSfLagcT1eYM4WRG1POypPMXXJss1CZY42uR6XtGLSR0tQEQXV1S7QGzL3g
Wokgo+sCjf9rNzJ29B4F6F8Hls3jEWre1EXWO16xQnXO9ocey0jGBP6HbFBkm0dp
S167FrrBYmaMNFLRDBNnxS/cg74upbQh751iixBiiPXbJ+A4ykFPOzysnaSwHKya
gX4QbfWp9mTXW/bET9LUZHFBFJhxrUzQ4WUNJq3V2Tv+46ap0EDVQ2zZEZhn0plo
h34pmn+r2cc8CXd7LIiPuBuFO/rSJjNO9IlJSK02cD4LBmaOT2CHaURF8ENBYZIe
1MAnV/F2//Yo66ESKwLadkPb4BogqP6bbXfwopfPeUlgh2CboxzU1FQhQfkDkkHQ
4ucxXNsSXW3FjHJ6x6Yn1lGsbJUeopKaf8iQ3hRrGezfobDYiF2TloMkAgxU8FQG
lMFhKkKLma+WSv76/u2/WyJA7SUeTeUFEgbTp8tlkNdUzhtYXx0gIsRVyVIO+hEf
s6rjW4jkZrxUGFzHVpBxReDX2JMsxD7zs/kW8eBWgHkqyJp+U7Dq/wMWxo1fBAk+
PB/RUWUoqxj3gEBGIxDTSkmJaS5Zc6C+8IYTjsh00bF7aWT2ukXd7YzQKynmzpk0
8VC7aYE9O7//tDwAhrhxXgwIFCj778sDIQYyXlMDk9MBlR4wzli4hgRdrTfGg3DE
pgKIHTIOFwUrhQiZ4QZ77S0/LA7UfvRZxARIyC2+b6NUalvIw8nCNTE6iIEEaeoo
5Xt/Ucc1RYprk2M6QEfGHUrArMfOhPbUljg8m4oX37H8v1wxmrluImr/COkbkKs8
aRGCxSTsYR+8l3iL9N51fYFL0nCKlaKSQaOcaHLa/4tjHbNqwD7N+gjluVe617X3
qA7drLlYVtyYgPp3wbSSdvm0iT3jIJv6Q5Y2zsnGWM8T2dlIBlGwUiC1nOSQiNdz
+bXjU0Kkae2sc3xIjNnn1CMc4r4YCPNx6i2nhuY7qPWj0BXJE4ydoU3A4vCH6PkO
lS8teLzkC0/4dYhzCqdRJvJfdncm+gHyDK8TdG+eEal5+1NLoF71Rfom/oO1niY0
twAsrnOcJTqqNwpYTQihGTRJTZOW7JyiIhfw3ETlUw1aKszt7k30/C0XCrN4HpoS
qqZzf4dzA8+FwidtsfOTH0KZVE/QPAF05g4NcjoDj1PbBQBJTTGxpDTNTH/4rauC
oSjL/zH9P1O0rToq0/2hW9g3Hl2z+onUsVP4hl54eYARfPkMmB2NT+O5GafW9uR/
GazV6EY+khFaMeNjkovJrNemXF7dvRPMp/RVf9IKXtQ4/axIFd3WtmKIcaNxzQ9f
/Uqq/K3R7weIZ7inBC5TuzYAgpzuNKWN9UGR+jhByKYGfieACHljlFA0bKxKDptI
z81gVLUDLiDRMdq0cQy4v1N/tzGlAbcfJDMhYWzs2p3AOHod92hfThHDYiiVpnHH
eoiLVj5RJBZTj2Gtvy/nQkN+bBjl4Qlrm2B/LGqoUewn5IFXwpxr2Im9Xt/jDxCg
grwh60Cwr0V69IZ6cQb0pVpxy/RLePqxFXSZ4jBylQMo9S0qJkZfuMr5H0U/kDUE
Y5aAJIV4ek+aChd8LhdqcQbt0a+XFieZcPuBowTLt4Judz4OlbR5pOyZydwRwiL+
JmBZBJNFychUC3Dr1VOX94h9Rt+zyxxt+CHEQSav+a0tcxHmyU/906c26Em2aqKY
DNJ0EvdKBIPECzThcy9EVBIaAOwTL/XqIfVSFFrGrxIWofxYGr6cjBu8cZtcgLBk
BxPFhnUdTphCJopuOf7QQ05tUCQ3hXv4TXf0hX+kNwo9unuWDf9ShmZzrF+ywMFi
6FtjO5Nfu0ACAwu53u3fLjOuiH3wFp1qrd9IWf0fn27+o4gcazrYCMS/SNvNgKBU
DEaj2C+TxfwSkw67dZ0xbi7QrJSinOIWBbYAIVDRdtTXlAhJodohaEE+cYv+vA3q
3Hu68sR9Vk/Osu9kNAW8KRI2pkTDPmyzjj8xLSwLq0sPUycV0h9VTwLlB8uh0PWw
If2WfFvK93laSj1rpt82WAC3a932vgGYIeV6M7BFCLXt6HQujrxS/2hZ+z8k0hRL
2naGb9avQ+z3wLaVbs70RcLyKSLWjvmnXGV7zkdqfbXFVqWvxtvhDf97FHOXhqlQ
sFFrHpv9V9xgjWBesHBFo9durYQKMmHJ7Ai3Ok/dFu97AMPcyKCud0b0bnQdZ4B4
k5KUPDciCkVYva2HU1n0xiF850+ar6bZnZgWmF13dF6cLnVNrHVHLT4XFg33fb8q
ZsZiQOi7JK8G1BM9YSgYSlG6eYJNT/IkYjbmXD7IAVl7ViC81z5Y+EW97qi2MgPI
6aGvOzwjW5lDtvQAzLdRHnqo5bXbvq7I3e/Z0OERhs0FOQPiUV2VFuU0HpROubYZ
tRDaABKFfFffcEpiHON9619ojwkUsOZ9fweseejaEYsKxLzQB2B2+XL3EUyHzrri
XET86nduUv1QdfBhtJVRS13DPBdzCInw/LRz+YUu62BTIVdK/03aGkr6GcovB7dB
RNbj0GyHkjnXwBoLPRR8/e9dtOIUNpO1OA28UVurZeMdAAHRXZK10YHBxfO6bwt5
5ztM5IsIBWACIA5vin6OdR7w6vwnVkn/eC1uLjZ4Hpn8OMrRsf7zSxL8PaBTSAM2
Hg+mJElJxS44TVXrmDi+Ar0lP5hGrDCDWDrLthyc3VbDLi9vlJwfu2fiBQXToT7f
wdhGN1CF0uWrcU0UF31iJNq1Keo8crS8TNSRMVBCskdGj2tDbz34djGCK5mRp4nX
G3QoM5y3R9EZORPk80ucvF2T8T6n8jqKz/6G4brAhXPizkiLmqJ/D287WalUi7IE
hOeLdAf/NrYcXatv+xYGgufLU1gXIiDN64MgBgp23hJJwG0kO4Wtd38mKd3x/87H
Msut3bMRp1warU6hNvUXACHa6GL24muD8jnQ75XZ5M1Mt/LeJd7niJE2UbkTBphJ
RXtMktGdyDfB/Kt2d4QKv98ajVhL1vLsheEu7NbpaawJgvBIEy6ohANn26lBBKZ9
b6xDrmF7H4gMu+CLq2zohqjkIPR54/8kphpjXt4fpt84Gz+JPOw4NvtXGI52vSqF
JlpKbI2NhrbqTvvSo5PAm4MnHzUmYgNLs5hBaOCgQyXQjS2Q6LxzKixrbw5AJ1RZ
AbhMlUiOsUUEfPI2yx71XnsDZKv/JAcEo6mrYVPToJUldd6qzTpuV7Ob23ZYHTt0
SNsORaTMfiV6qFxGUz4QGcOaKxEr0pa6h7IWo+HG17lAh36mqmGgEHhQ2TDcVrLz
sp5G65tCcRk5iMJIR+ckUHOPcidkv8z4MrX5btsMbEqWIRmwJhZPvEZ3yrAhOKon
xe56VqN8RjHRgDq/UTY5o+58KD8q39O57KKodi+Tq4jaL7IzXbfYYBF4WOVnxrlM
tnJSi1vi4bjYhwrgVutU6ij+r3bunlkpeuTAAY9WzU23BYSdqkPiy3P8C6RaWthq
VSbLNlpyiclOJAuZm9GPL9xb53lk6yDpiEJSVdxxHWwoMYbugknxxVz43DZT/SO8
odUpEoXKCpDmL461quNnZoBxiJKbTOcdoPbkdBU+CGs+v1jPo+n77qLWBGKr50Tc
92qz+sVQQTR86w8AOiBTm6Ul1L3apiXw5zHQEJ/osDTAIgjDJ35T5GRAj44Pzj5b
dSBXMnfrAvBgA+gO7VBno0cLOUlMMkYxqVRvcARA+hA+cn5/OzH5ZJkcOdsuWWIv
0GtK1i9NMb5+mTo8h0b8tZ1lDE8eMfztVmrhYZ08plCRgQ82BZMARdEDdyS3r279
shS5kGygXqHjL1+xO9hQsvhY9apTWy/5eCm6K1G5gLYsNxaPm0bHNlCUr0ZOxVQo
lzUiWXFTUm/3y0r98WfBel9rPyWRt9dNfJfkEP91sOrgr2rdAKTHXj1G+ayfPWZl
ejCiJzK8DveglAjh4b/ziser9vyr1m2px0Z71q5LxYW/4d6EgDHEGkW36W6oIjEk
javmgj1+Xpf0Fyh0K4gC2osUzWI/zAU8DKOt2VbICxpJc25cdEboRk8dn+/kuwP/
JkARy69VRyKQuyypWHuUUqDRBMzhqlbNwSMAgGgRjgzmaD1KhQ5U9EMxhOoaA1TM
68aDRgOhx1FcdSUplVhbwvwR2IVBfR8Ff/sp1kJh7sj+RIALCvbHJ9tdmMcL42sJ
PQCNlJWZPABpSdkQtg0tALCb+cWheZH2xR/6p2T3UsWfPjRzmYW5P3mQYKE7jf65
fTIzSipgSG6CTICQHA6GTMpH86AQVFaBc5vCqbQ8fgUp7ETZ3OdEH6kVx8vB14ox
DbbnaL1Ai1o9yDx0dNNkXDDjjZRtJndQ1DI0A4KxbWOqWpYP3GwjtvxbNVh5d8Vb
sSogCX1+wA6WPw1Ncux9fQXdtdhY4wLUA487XgqT/WtZMjbTyVajtnDp2+nXJh2a
4S1gsAMUVqPp4cssqhzR9ghhTcYykVS9l8OZBlgZWTQ6BXqGoHUcJEVnyhJxfYyz
NQOqFiM8jKDgE8A1vodbn9kS5h7Stsmazsyt2jEi/iHjDBuyZGVkvcKdFa/43oSL
OKb4ViRFHTi8KdRWE8GqKuuWeIphwhDG27lhREwmUB2V35oWxBWJi6B5gxmWHN9L
AjA04LbpgxG42GsfOKiIMtQKNZ9NxYf+Q2CpRqhVYPaE9Qr0mQfOMrhaA/tN1yLk
BEYtESIq3A4GRwVQjXmGLcy8Bmc64hCznJsI/YlbweeuoAOag7ar4zc27b0jTy1Z
MF3jUdbNTjylEoWwdMjnSwaAbhQq4OzIU7rASoZBcvIYm4p6r+tlVcpQ5JaE8rUf
CCoonIk6mw29IagXh1MFkXF+ZqoqGbvmteRta71BQ4Ufrap3FqcPfDjiVwLbDNos
z2qlETry0HLT4NMDAzYivTpMGJBRMa+Ocx8svUbdCjAaI8KxkxJR155RA/KiDjlV
6Y5yCXwB1MXuJVOYz433O9nw/9hR0UDtGDdpfsjC8InUHTqcXmJIj3gZDscjRexk
UzQw9vcEd27pxiEjz4VUyYsEnEE1NzS1YyyTdDfKG5rnktB5OsR6tIvTtUsklY9K
htyB2fGErc2aAZgZaobrVtZRxCwEjZ8Kk5oYfkMrZgxN9iLusTJ8gBbVcsp0w59Q
GR/iW4cvIlZCVBnFvktLYjBwf+HqYjjv65hGrdjO+oZ/vpwombzkowpMpTO2s6sO
ECXs3FNDKHa9/SNjlXyVU6xhKXSpKmbu/aTgqoziTRgeeDMKk/dpvpS+2HK5NYfI
xijhm4WjWRvOe1lJSvxEiQKTu+H8BL+tsAYx/dqHOJ+gXjepF5fi2eHm+j3do0e/
RgdWKmaRInt02doymVgzmbChXOZg3J13zZNN/Cu8Q/LoyyE2d47dSbUwgoqS4geo
X2DoAzmXsysVB+mD3Rh1ItcdbTzMMhK30joTbSbxvD7eu1jlrf4wnZ29wTM6Toog
T2M6cnDibc0C2fb+QH21f2KYSC5CrDAw66Zfa4RfoejfnfH35dkXTmvsMtbpiJn+
wBnuqGOSX4YFmARTvwiXNXf0hDR550tCHb14nDKi/6A1wWwzrHXAtyfB5yN4s94J
Ea5yi/GSiBuC3ruuX0bdt6pqF8tn/TW792pfHv04usaDtHsXhws8nRgnupbs6xq3
3csvCDmLLk119un3QsxFTRu7PQbsVdiGDKKEnbRFRxqxT6nqUwGboItIIs3UITIT
hzYM/6N2AH0lH4dHWyMRX3En+Ibj/k7DzdXYNs9ev1/s1u4bVbwCRejHHwo3Ioaf
Q4+LfEbJbSV9MaJFiQJRiOP6ztWJxnJT9mPPBaHREgShGp5T016tRaI9foKGYu5F
MlbAV2hQouxZlynHgS/qAA7N0fZDsgvynfTuEO6NoAVWTHDTQAB9PomEUVQDOWd9
X6tRrXNHVwdS0QcddCwBDtQP8DaLtUQAnXIoFYZYNXr7htlXl3Y6QxggGe7vfztC
jnR+HZij1nAW5Vd7tkH1ZfNZL9w7e8Z8KFwEZSE/qIyncj4Yd8M+iEF1cUWmMYws
a/HsiAL3b9Euu9wYxa6A3LMq8oz+Hc022PYNR50YcTtHK/gz20IdOTpS3x04se52
u3oUOowA7UX+5WyV4jy2PyvQ21m6xs6oLOtIYXYXpYVL+qZsxZ/Otg7abh0Vcdtw
/nYE/3VfKKIw/W+W0oV7EOemrUvcbmIYOfivvnqGUzl/BGaUWWp5nB3vr4tVoa++
NynhG50gsc9TCDKRGsDOl4B3xSDDP2Awphmm3QP6hPrjVY7Iy9UmYyKl4cvl7x1J
uqAG2/jf/qBHbFQ7bW2iwuZIwV3JB5zp/eEFZrkj1OlvsEcLgh1N4YOfR+w8IYtg
qnqk1vrDypGw/QQwCn1fWoxU4lo//eRzpmXPVQPmZwApbfpxEzuM659VE/SKkQ7i
z81syoeO9D+e+I37JjmfiGgc81zHnGAnDr62vK4y82agQbcErE/SajchLbMmGCfL
Ra6/Lo9S7+VVrKf06BOZCNmACiuvR/npPwwiayCjqLSYRU/mWdPZNCoDMpoc48YD
9BsGFYiqPkqi3qReYHvBxdkhr04a8V9l22wHoAiecM3Fxtm69M3AwlZhs1an/3t+
rjm8MgjiQuvq/CMnqATtT82YfMXepG5hLRE2w0rtMzHkd5l3p9Q3UkPBNGWh3kSa
Fn9IlJo1MygDYMNc0bb+UzW646CXcCKQvEBj4eZs1x1EZaWrWkEOIns981FG9Cb8
5mYOOFB/7dgtFtGeTaVvFLxFCXHXDNRuhJ4NcRDoA/6EU6ss3Ae9aNfFosy4bnSP
7zpz5vsjBVXS8FahCGWYUk1x5IVEKF7i9AiHinQ4lb1L9nPXMnzIUMU6/Z9l6DBd
zt69yR5214P7HklJi4jxfc5iHJESWqiZ5dnncVFIhMzJT6FavnLzS+TTJ/lTjXcQ
ftQA/J9fRSNCt5g+beQvG1JlXw2h7ztVW1EFov3i0FAul7JoTTQqO+Qs68BbRzIl
8y0cf9agR5gsd+lsnp20wXGlwL4vO68NvJku9SxTiYw/l50ekFCDnzB3I2Szsuqi
8QpUmZ/wP8PmNPp1hoO5Xw+B7n28LiIEV/kPlHn22c3Wjbk41D77ixehnNyRTo1U
lqoohFsK9ZYDRvDZZXdlIZ1HVl9fgwG5DfPKqxdYb+ldeAzet/ez2N1nYMMmdK+j
m36Xpkl1bFC3mVstjNyDaPmnEQPqHd/GzuZu5ceoOxLsiGJBGBPOzwnnjsUySDPO
lg1dhyMSgQaCQi4Hn2BXxHTlVHInFDiMTfB1/pLq8sKzN3MZkkf3V6ccmEQeW2GC
9GfpHVm7zLaYuTOjr080mR9R3+4TR0YB+/xAtgTTm6VvT6Pdd/QIDdKORel5TL7p
sk680JbvK284AT4kvMYa6jACS0SpP2jK55p3IJCwKU8McJWhD/mM8JCqSBnPPyK7
6YJXWUwPescCc/jf2O+3vW5Lhf0524ENw8BN2SqHxQP8jRpVeIhZDvT2X9Dv0CSG
zC+bz7Ga9GO7oALq+ANyETu0m+wK19K0qJ2aCVkVIdUV9BmlUg4vXggykkeXzXbf
VXSMmlXiwXjItoVbrT1IV1lZV/pK0jguc+5rPl8qy/nLCDURidAvBdbEQ3z/Nyft
H4EkOoEXL2BWDA6l5wGKg95WMHdKbVCjg0JxMhf7HXihueJgIVMchXpBrpvvCNrB
5CiTT/o0maatqz+7sUMQi7uwZMrxAMRHjR73gQ7zEn34fopBcq/ZaXHEembLgorK
k5dNvFTsUepLCo9KaZyt+JErHwuwMTnB206kUIXojNrPLJAdC7vjfrouFNBIx2tu
VU7a7PQKWmcgij5nICiwtOQ/YeaRU8ZBTMiSDfJ0p/GU+ZbPLSTinNcYjM91OYYJ
zYoOTKSNjRl4pc8teA0LOQpBPph+Y49oEC54pOdODodQhwvKqK1reM//nHR3utPG
YiEta56T97UV3pVdtXfAhyh6zkewa5oBCclJF4fjRl3UNwfXOmI2Y6f4MsI8WSpA
5KSE68LV7DWfWVF3LH5dPQqVD2SF6qYjr3NwltA7u4liFLt9gSBDPT8X1FLt4leR
LFahIlD6B/Q8ElvDOfL5++spQsj7Q7K78EG2hpSWkAZLwbskSHNU09fGmUS3LTHZ
8SfphKTngfepXHhXzrdv8E8yUC/8DTmS/0BtG/W1nwLfdgWESXcBzNUJBrWdCAlC
VwQSVyL6xLOTCqU1IhEH/Q8QbaP1eKdIJ62sK4VhoDmQCaP+VuH1orLsp33ls4nO
rHzNmkuZDFjG2h200YnY1ORTO/Va1rJlp0ZCP9S5glV3hZlJNINsxYJXEdMRLO3D
Fhm3rtmgml1f1IiZMIKOROOakUkab1ge6U5penzwqgFsyWVz8lgL59pY4laJEi1w
x/HH9HwP5PVTP+qpwOzHZ6ZxlIOhqM+/JkEKwJjEp4QNKCo8DecZhj11QHkp5cd7
Ufha+Krp4YFxFBIZ7Dhx4ZuQouoMZdIAvQqH7cv/iWtMX6FSmsoZK8Ljzeyg2kw9
ryzW3GzgYhtg7Ib3AFsCGsLEx2S8oJGOlfA+u00lW5RqlVWoXnHpPqmwhc0x3ySP
tBUeH0at5usdIweWqnDPIKc3B0StYIQZ9hSgRxzolAbilUP+zuaoTsszTQLWY/Wi
eVXj2TM6lpaFWwOlYsVipfbzlQigLo8PzC5n2/eaT6/F7pHUwH703r394adx1XxA
pYmc2Tiw9oQEL4ivABlcaQeB1YpBsSikFyB4/lgK2o+msTjtw2B1QpDj3/Lg0E85
FCb+JjTbHGxL+u20PGTaKI6TZRcQBbDuSj0YHQ3DsoCGrp/f9dRgmfaEPSwfAPkE
QxrCscmuIvixLzrTTRC7ReBGxc7i7/X/KtQS0uyul2detwKtgCp2qX0IW6jfJDtw
U2GYgwuR5RP/fFp0j3pcchPmovg6Egup5omHUYRhc1AdFVgqrxDy1Gipj76EeAJr
FQFH8b7yJ9Kxrsi29j3u3KgJaDDFCrXTVY7h1JDDfPqlrZyF0waRXeKJbdnoKWiU
oN7Ao3qwaKumhs9jhAT8ovYidD6/m210Ge6wQaxyNT/tw/UPzrlNYNZ0GwP4XwIW
BQt7LFdft3saYH0idS1QbElMm0b2fYUv+ij0jQKsYjAHKJarWs4s6IB7lEjJ92xU
aR/apE/MTdRBlsG+7/PQrBOng6EtXaLFDEMmFT96Z22aWkPEZfLmRDpFbwUhsDUA
2qyQVpiII54g7ytaTNZRCuSkZLd7QqAUBqzkib2H/XV0L2uCE/52EKwIuuIIausS
z8Op+qfSGfZXbXQOH1l9TRQH9iMJJnaivACJhPR2692M0F0lEVX6zdTGn6g2/Z37
8nUrglrtcitv6Q2Gi6a/bF/PKISWBjl89CvMlKx69V6Nk9NTh7IQ0ELMfO4j8TtJ
1JwHqv2b2Lj05E63q05HUQZlin4DU/PZyF0rS6fPSzZOObB2QaNWIm5rTV3xrv4j
UeR7LcvYL31VhNW28s9alF4Qxe6L3Anb9NyplHB1E14BtT+8B6ZvBkTdhSr+rYZd
VND7wTBVeuT7gb2mk+aCwUrWlvQpoEZJ5fQ+Uk5Ro3p7c5dyKFISEbNMJUQgVo2C
2FKUydLJVYvhNUYSz+AlgYz4m9ZTpzhu12GF/3bjClEAz5RwuccxRVaWCwCo+4P9
RFSGzoSILF0uvC48FlbBtkwuqLFtXKmYgTlkt7qO7F7+gtRiz5vJozh3K4UuCmyE
SoWm6CX1xlVXk6bTJVtcHFz9vEN8A7+/w/Nz1DIs9R+ndW17mXh6neJQfTeMD+v0
xFE/TTtodXCb3NcOADjlmufciUVFoV1tLjziFMoukRM/JZuF+StWyXJ+UiAGo3j0
G4QUWFNLnFM91C+oKKYn5kYpYKk4kOLpVDvgeol9qyrCo/AylMOY2Yd9a8Mo//H6
mPloMtD5UMMWfQcW+49cUD0ouK8k02M6h0+tFYrtVkg9ofqau3Ja2ceUaKR75iUY
ASVOdGf5YeLQ2uD4z/USjtKHJVDm8/EZKhUTDJGRUDwpm1z/mnFs5QWNMqBQH1Yi
CwPNckQ+fjU0DDDfeBtlzM4rmPJUXRwYa3ddpnKeBVP4cMMIFzFvMGiB7+BS0UlK
XJ82PCN759kgeiOubuxgMK7nDIG8H13g2N6M7EOv7Vya4OCUBHieLZ9FDEC/GLpv
CW+uQB2w+9xKWNtuOiDioqO1ZBsmKqRwFww0zScbs8izKo3om9SnQKWe5lZLwpav
QAFkzHfLjkQoyJlqYNJfn42uNgWDUUskk6sUa/3Y8I4vQgWFPrsBxcRxf3J+l9rZ
rlhO19p8WcmJMUqVuuVDs0DGma6ynGEdLgJuxtDYgI/w3Vhd73MBcugCJFwW1Rno
nAs0LGjKZnGEW7FiLvqLj0E7SaQ/y9B8nks4FfoqJMKDMfQ3aZNCnJq9TdWo8eom
PbEG/QehKaWL43ndoykjtHWQKJk93i3N6zg7esI1Mte/2JNFO7iRTGgzgVHZkm/4
XseHCzqnK8z2az+QoflRz7NlgWIMbXUdpezkGwjhSYWRtzbHmFdm7kTntP5GZeI9
01aGNbO73A2iAcBqNwIBbcg/LfOWYdsC4gA8joohchY6KAZQeB+rYwH+QGe73FS1
uOaNE0FJekZc1jm36++nDnb3cweyDPJ79AS4MHYruS385XxlXq2fK7D9vrcakY2l
Z8XTUT18aESSjNuAysgyPCzAwZc3zBCY5sF+F/skGDt3OFYi8DOkWMFfrxUzJxxJ
DAD1+DTbWHynxi8sJFLpQPmPSW8Di0vlPLVZvQ59iqU7AZNGRdyhyojozCQMeVRO
l0UE3yGG95jtJdpCQkNQN2rSAcjd8FP42DAMecmj5UFzMU1B1kVTxmlOrIqrtejh
tx8XRQHXDdh1r2X2LYX69cTZKWCfDvNWTL/bqGovkK5LB5TKk17mjB9PfcNf6oGG
BpIDuuVsD612AO1DcKtT+b31mEIkZNDmNZorbezrnpWLvViXrIOI9aKlZYZ3GSB+
3X5dtkAKjVLNQOOplrbXc7bKd7RzWu74I3REb6NxZ7aaz2Y3F3//LkmLKE9TfO8J
0d/gz9RgfNLJ8eVonbl9I8pzOnRy7bWkvNUghgox9FDLOFLVPN8cmu7cGxOSpCde
rX0posD0VeQfN10GLUVfU9wkEzpye2hbXbQtKEKxAt4c4U3OYXYU0nZbteF3Wc6A
SVwfn9RGB0tqCD7a4QJwghsVuhq3jco9EYXpYxRG367ZKu2p4fii91LRz/zeUfoj
yC7635mrsZHj3MwBJeZgag8Uie3Is61eai9jOGd7JLrSxJR6nRG2ybgJsHz4us9H
u1FbAjbEf8Z2IZfTAkBU/tj8AxEHuvbpZGoNZLDHhBWOc5PyM5PVaKJ+eJiLmqAY
UFL8/LAQeNIWSLCGNuKRSCQ+xh17A2PczArU4duZRahsAkQu0u4fmdF3gYzlGGMZ
9qfceRmf8Vj6y5NXhzjil1nDBh3QFRjh09W1QGPuz3FlQNPiYLDVhCbhGG8q/qBE
jt/b2fABLLzuSeueXp/Ldj6PvGEnDAdXZAV5nnsneribmTHhltBfaIUm9qhswWnx
fTr4I9XdvzEShGS5efT909aPqon8klGoFYS/sdbrx9f0pSRLDKjV0j2hNQwSRjgd
nkgmuNyEO1XcVeNwBOUFaZVwFs14PulANyRKFFBuI7xUvpqUKI1kPNCrG7VyIqRB
MXuIREjjHhGUbwSpWdxbYfJtD8Nm8uAfVRQUwvZwRvMKxfIiO1YJsglGKg/4DeGY
fzSYSGQcM+6ymznTDU/MDF3sMd8+HYMrJKTce1icFtueNoxv8+rHM0rQT0iPMHOo
G9+Y/NsYfcKVrfAOEQlvuadNqUd+m2AFipMRlvGxJHvoslm2q7TCHHSTJHdYpNx/
7F0WA21xZ7ZvObw5CeOIDp/2TYHi3XluEyP+/ir2bqhTTXkl8p58mEaJuqLM5P89
++B4eG1Q8g5uM09qq0MRCjemxxi5ZvkjBVkQmsnDUmzClUVC0LrVCA7gbpUvmuoW
PqTak7BCoQk3uwy//9zAzqV/+7xA5vK9/x/d68nz2jueEhQkUZMoB5WqUwfrjguu
07hBaDIdJD3M3c+f4PnL8WXhQONX6W8JR8asq1fm3DsnQAx2DAobtKTQfAy3jJ9x
9ZTTg9ZWDtIjgXxtg/rEHj6QDG7h3teh/0JvkGx0FEr9Fq9OCOkQY1j8+eWo4P5b
dXbpr7OujBHlXSkPBeb/xTNzKLusE/8SJwALdudRGgF4fonmeWHlOGr8GGyjHOYF
a98VtYGjaZDchgEC00SliExsApDMgEurdJyKDxTgz4rx883Q09caLkegizFnpHLA
zLqmlTgOTu3yJE7O5FSMFaTPZ4dfpE9Mno+wlV33CDcG2BpvYF3aMRIFBGWn91Kl
F7isr1KmNl7iju8DkMO1BdBsu9YZK3XaJPBvthEJlFRi+7CJtzX/L8eRXDdfBb6g
WqqdIUY8Qv7tscQANnj/nZM7e02RQXabQ+bROFG9mpfDBa36/YcS9UtDAjIOIP0e
v3bXDfBTkn3YKzU/a/llo6wN/fJg6G/5Yc3Wwpdu0tomyLVsVYfn5C81SoFyebdj
Q3U0IlM/TZczlo3c6zhrGtThzlSZnuPCkJsoy+vzzo6KwxyONtFFpDlm6r+zEC4Q
0cohsj0u2xjAm1/c0dtgVy18HNNDJB/QOGT2UeVElH2LD5CUGzNRPOYlY24gCMGP
/JzInkJiFQ/yMA8cSNhmMcwJp+Uk6ycXhGQczv/AM3C1r3Ipr9IWHEnOnr36+IWF
OKFKzyAe6lvBDhQxUeXhrr8PMl1PQ4aLX7DUdOKZ32gVZL9o0RIV2j4y6kZPndlW
PkxtpdG1YVIAKy1uf08FQd9Vwoxp7eVZ0OtKZCJeCmzVWp5j+6RZq+KY79jD+3KA
57v+a233Km0gqxkOd8NZb+8Xw+eZp7ndLzekw34v02T6+vs7xVjp9Qh0+gYwv/RS
I04FE2+sc4s+QNamjNA/03R67pPGaen2MakLTUYjgC7po60zZoRjfzVNyNGaH2QC
NAPBghyTDuwlA2AW/U4j5KOHNg0URDiVLjSFslfWY82prLTST2LYxKBybB9yo5gR
fBzbh5IfPowelNu+wgdGuQHAb/BNko4lLHGTEveVXHJO9DASfe1Sd+ck0zp0aWa8
NSCnTuKIDvIoKsZPatkPqz+uJHB1KcW+mxkXcw8GfK7I7hwQ5U/rsPbtR3UwvjwH
9zPZ/LwGLLu2hMMvj+OjgonO8YcRMoSbsncr+e6a4dbpgSFxHwGJsFhzKDZPZw08
AhYQtFO4gVr2N3vI2Ox903zaEnftuhhhZBLGmWzxqzW5fzF7rYeNQ3kS3k5mG3S6
g8T/wBzR/4zjdQnorFLJ7gGCZ4vx1KLImqnG/9VNcnVL049anOkszQvRfS0AtFEN
2yI/6ZL1/xm6LjX4KO4Zdhxyue1r0uvCePIbEq9OkBHVJJv9aJXTDsJiOlT6F0M3
Louglb6i71mY5+FsTlaQ3trKT+kSlnKD3xV5vMWpunyMh66EKs7IynLXzdvvyHfJ
TQzvYKqWsyi4jJ6wfC9Aaj1DxHeyPUXJxcikoFfMXyr2vbFHaGoFNKmdoFBiO/Dk
ClGrOTn7IiMl4RIo8SbNzXLDeLQtNgkUW+Me12pkrnAPWuvFtvYxXHSRxkN93syw
erwE2SAwVnvoJz0kpFsqX9wa209E9LwDWKqeZ/7gz6c=
`protect end_protected
