-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ewr0EH/GTs/gztfFDh2eE74prrxcY+qLmgZSqk0aHczepZk7H2yByL2o/HAyqvk062Tb7nL2QsOY
GpdyfsnongcFjpVUzn3ydkecE9ExwwNIj86+7MxT/caoaBIYep9HYt9G++LNhpLNTAPQNXE5Ru9C
wPWcrVv2jIChUU7KlrMSY7tx84lT1i7nAmQSTvM7vhWPny+/wgdzzvSGomHulQaC3P5OnQ3ob8mZ
zWPjHS8wfMX6X+JedRT6lc9DuN2LOFodTamxxmZM60fxQowdnLqAKZSIO1VdB+aOcOddxYxSJ76T
iJU37pArtxcJTOkm0r4F16Mik/Lxpg6YjAJSaw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 34416)
`protect data_block
tCryFBXOLrDF3j+h3213cLIEM1Icx3tAXJHbRMxp2ipNujofgmXq96YZWeRrA0vdzIN/99iMZzIH
j8LlZXLmLCR02CQGNGrRS6QSizMryEZOHq9mpFUFy+KC2k0t53TCQkPlHPzE5t4SzxW0rxfI5tQM
9sqvNaZWxSNOY6iZzMgdaUl51bhubQENtPDtuWiODl1jTUFdt+PpQRUY3Fwk9sLcNgI4hjd7vvOD
7N5EvwdszA8zW6NTqaiRxzjs255jotCKzUuXRZN11+QvqxvYwHGPDwAWpOXlEaUQsirqE9yFD0N9
S3xYFbraWzMVj0KH/gbkD6EVEmSty+Ugl42BjfSaGTFREtdrOzxn1SRr6+a+qIwx+IXHfKgZ6SIA
g1LQumZCfuuU+BnsdBFd+Erg8T8cpJwNcJmFw2d84L0dkHXZI3FnE56ZL6q9PKxJVX0+BtYG/+ts
yqAOuGEV4p2oV1sLCDrStVcEcNKJ0KTehJKwv+4a3ukaoUYi5Z29STC4ds7ttKbOTxbogsBgWOaB
t5WSxxt7wzGoReXweH2D9t74k2uLg3WZ9p/8Djx+XyFPURHt7Jz/Go9mwL/mLuM+Ya5mZ6KwEMQ5
d0zDXVuXs0KkRVZP7nAu4eiRBNh6QwYGRpfRqceUbmr8Z3WQ/0a3wwADKNb545mouhnewfu3FNNs
qxcAxsFHighzk5nuT+knPYqWdRsQtEqjKLPqbeR5hbwffF7AtPhTiUUONLEb6mtUX4kpr5gL9qqn
SL4ZomUntOvNUKtt8RlqblxaxBHCeGTFSyeBVDRzGMd3kuzS55kNqAPehM4ZlFYQ7mcbLMmU0XjV
dIN6hZN0XcEFq4gkjvzKnTcv6sdQmEF6KnyLf5FuGR7R8OTYFOLj0ftfO//k6LSVyvN/vmu+8hKW
d7brloYpUV8LT9TYycGD13+8sP3hvphM+ZPAovOionbp1J6q/+15IapLmM/bKmJIjxGU/2zLpIg2
WeOdub3X5Rw3+LsIROv3fpJWFjOi2QyqMoYSI+X8NTFgCkbi1qXbrUSNTfnvRdNeYY1oZL3Egjc0
1e3QxuN5zGTuie1pUuKTRAfDVwDrw6NhunUvf48jOoK84uAr8UudHRWjaEMPHDgTmVsA/uzxBUSZ
MLCHDqjU2cR9HGomJPU6eR/fv89N+VxUeW78uQrWuUNBhMv3GA7kJOVZu6kNkTeTyP3QF9zWSb3C
NIIZxFmMy2cP7/SrhTmpk1AeZglTt/Rm+kfk6t4HIQRaR1xclb/1cNXBtPlkCz1iTtEnUmgbKqbO
yEFeZo68fhTZ+y8n1D9ViKF1hRA7s0O76wemql1++pD3yMyYroGjnh2iXdApY3xQMeNDi6PFLqaH
WMo26z1AJvZItvlxQb5PR0k6CZ3frEcKXi6dmHyPqHpTh/mvyUzwjxWNcPzmbEPXb342A+yKLeCf
6JJbRkgCcWtwaOJDlSQLjyOo5NPXFkyWjgVf9s01las01N+Co1apmBVZiDDXNce+UMzLSeHS5Utn
15GcMUiI6L35sKPnssKAWL1kG5UOMOkg5lq+LYyR2u5C+kig4LPvN/IU74Epll98KakOiPnUjWba
GGem6XmfO9Y3aP476alHvz/nihO/e13/67ruzBHwIa8LP9cAkSQTrbUgvr3lAluNqW/etBpR+z1I
CUQzmqO8MdxYRuOkBnVwiQ7j4OjIFsyxWG/I3+HYjdCG53T74pW10jBcbPX1MkxuS1ZgVK7umO7J
8ZXLy9+ZBAlbMVr05l6Ebc5aFrFx1G6Hw0HyeRJ5NUk/B3hKkOIckyToltqk50NKmTsiFU3EiDDM
AVy5KqHa64UMMAJaDhAj24DYoJMZqsYNjQF39/7h9Q7sXhEZHE98XZyG9XIaaMZFEw6gdZobxSdG
fKvWoWuV05u1f6fBLrHwjP11Qtvhv5YIXxxTIe/cIq+Vo9nAA7R2QpuJHdRjSuDdfSaSRsWtaOdU
Mmid7ZyK9dGxSTYv4evfyC254e3NZSl1LKrrAEkXVG+YkckZvjZZIPQH82i/+GjVWdIxS7vGhvTi
U+wQC/HpYXcE2nd0Ys/MjGA8+Lem0fBzBO6mlz3nJQP9glCSfNWqgYNLGazBWzLLgZjZyFQHcP2c
DsryhnqclhLdqGLwXXKusEW6GFBLY28F5CGExyNU63WgtN8/Soi4aBWWYJgiicuGNyclGoLcyDfu
KEtRb0Fi6Y4+Q4KWCmtSmhgiCrTa87/5LpgmLX9eX13yAKbHXCz/X4xkpbvvmo4lzWwzWR9CDyU9
0/OdlS7Utr0V+3K+A3TTyOA27coW+I2jDD5/+uQ/dzFCeF+qwrh2ldZxfwn/rZfnjvh6Xewt2gG3
QluOYHlEDsN4RdiG6CNK+pLvG5Yno1VpeQ2wKljj3DounsiOjEXrQe96yhrDEieNhoYENTRFtiT6
rTaIAAAYwQpQRzHZyrpNdpKUXN3iXCDFQjjVpr1eG9TtP+8zor6cOwE4UtxlYf3WCt9qO/7A7RED
kE1LyP8QxmPcCa1cp24oUDrjdJfx+ZZfriz9OiHB1BVVLX+PUDbL5LXTxhU3ON1HVXxv2ltdhTTp
9D1sWYDIqFmflEt/vFARf4CgBT7RTsFiv2SOL5zhcFdxOhRrQzUksJSjzoQSWk2pJQzTuHrTB/oM
PTKRQViwnhEFygeQDt36wYHwKnxSkPdfuwKpvxTWcPJeHBkN7QdRO6IKbaIqaZje4o3HOLGKNEOQ
WATpphsmfn6SfkhNeh3TbqMuhkZhnUi1NnXeY5Btc56ASmWvsir5S5ajZYsyvbVWA5XnIi3WwFqb
ulihfNPWT3xri56kbZ7Z28GKzxUvugcC+rlF3cGe+KhguARgT7BQR12dyKu9uAtrf/iUAIkr+9EG
VdAkysGRNRQoz6rVpSUqtR/rRQ2uh96tgXZn7uRjOd4wItjEKw+MJB5Hj1P5n7ETubYR/kCBWqAy
HXKAj4+215HKKKa/9qM4mCzGgMVqhNMzaivd6fMJCbTBiB2rlaYsuVS+VoD+YnShmnlKkXKSQUAQ
vCEKDYsjB2auMs7uX32XVjaiIWLitNVuz26VHQVVTb1+39cNuCE8q53G1Vd4Sz6N5uZfvZarONOB
/DO33FpMCgZKOE71PhrpfIDeL+JVTzMthlGsWqf/jchoBpzJvrffjHKArxAwEQlRlThX1GAoAOKc
skeb0XvN8cUEAhEKsLur1L/dj8wc6Q4lPxzq3NiE3inJ9aoTk5AG1QNoFzkwCayoQydg74yq7YxN
47zJ6AK4bjQmOsiIfibxT8HwjQ0S0Q6XXP1tILexj6GFUf3HBaWogTXK2kCmMp8PjE7cMzld3nOh
/Ycn/eJkTweb9bamz7m7FfQE15oGaxnptmAZw5JT0moF622SbseJlqzNQm2fXJYBfO2FTgCNyVpn
Jm3HTLxfXxOGc9Ay8WqtJucWzi0CJoZ8qhi6RwCqQlwMaB2gsSCdcOwUizlb/GuLsyeX9I/IJwsI
us6MZ69xGLyXg1HrhL0Pxtr2rIaV8KqZv7SzHyClhPNRTohZN0LrJdwSsrUowVKgr5ya1VkAP0yv
Yq8cngQg6NbNlirRaxZFmEaqs8pdOc+/hRvxOJTVT+KRYjuM2MmfSijHNWJqljU3lp66ZEL898W8
h8hW/0WvAtjwUAL38AkNzY6FCm3hcNXQNnq16lmRFk48uGSUSqDURr7nUnuIafIUpYwXA/0cvcFI
X3JcuR08y8JDXnEfi4x4H3bACDfvfb1SbkK5oZit0udq06mzurGmEGtYUTDsfXXzzLlhPvmHqbOa
qfDeO4vYmy9AIOXTXvZOkblucz3L4OhgzL+CRi+3bKX/06+WexSvRkRkcp4LDiT+CYbk0iZlkSv9
S++jCW6KIabJnJUXi2v+BU6OjwxJklPIvYs1ydwntRuagHbLi+x3eZ/14rgED1Jv1PZ18T25m0bW
ka9oEUXSyK04YsvfXmwSnECV5EP2N9Ay993lx/jZPUjPeh7DjoaN3VxgKeR6UU9Xorjuf3xU34Xs
SV7wURs61AcKZGg+w3n//74kI6l1+y1C+iTr5LDb4nyygLp/+QX7l+Px5Y/uIHPLt4TCGpW4A21M
9NdoD9XSHSJX6//3eA2B5TpAxMl7rulddVsnTgnED11dKujGbNBC9ry/pXaZXTD9RaVpeNvQ8+o0
Y2Rh4KvYuQrrS+nAh9nfMElmOqjaUoU5DQOSilHoAEaMY1jvAXEaR9qK0WTQRqwgJ/Luj7SAOvfJ
nFQHVQ8m3l4BIkMnAPMJ/+ZUUGd9uhc0h1lWvuZy3Soj5pqQZXJ1uw6aGuoARFJhcje5/Ftr+cdp
B8983BdL6eazBRQ19EkBU+/nfNjs5hZswYG1XvrXwBo6EZvVKom2GBhiaYIKescmDA8nn6pytUez
Cz/Of4kszTFKDdIzxnbjDt5uyBTEgzP8fyQ1A87E4MYaqupSWrNepMpBnz65ngji6suR6qsknZfL
brYlRIePjp2PA9d0OyENRRYZHBkVvuvKX8xuBBDZ+gsw8I0b0C0VvhPfuiwfkurZfW/q0h73DGdV
AY5R1EpzWjKCSd1KCCJtS0OBVn4akHimeBn0bd+ZpCx/iucHSVwSPzCkSvMhSvncurocgyO23w0V
tUlnz9NXHCE2A7b4rmp/n/xy6GPVVVPrZpY6WvclfgbSoxaynkxH0nLEYc3NyuYERyguU8SURRSu
yiBGoKb0rZZZ7XHacSq9Yu++F4XFgTpxa7S7vjPnpjdGZ+k3G6k0YlYEApwpxTdN5jmwV/mddZ2w
TU82TqhPd1hcOoolrWI3Fliyu5hX/F03KwXjMDQ7UC4oFLgh9U+EHAxIOjlVeDQZ9yPdETiDPYwM
VJoXLqnAhS/lOBJBelLlDliisqOQxrujI3G87Js9eYCWRIwdxGWzPP9mJjHuTkNEFs03pKcVryCz
9GnVtk6ZnK40lXJguzr5fLqVgJL3LK3GjSRKw5Dj2Vt9ggU+hD4xIkpR9ANJruR160ncJntSdQuQ
JDQuRZ77wUGx+D+WkKWNwgT5pbNW8N52lr0Qv8U7NH8EyXuTsQALKXtczyUuNxRJAUE2MzTE5IFU
h8QUSwdFpPSloiwxFK1dSByODYMsXrNuVjUk2QK/IKyhqXIAnSl6p1RzzbI9XetWCJRx3I8xn7N4
dpJP6lNGzzxhRpcP2GF95OkWCtxoWrJ7ScJZjYn0QYdq4V4lTSIIwj9LRPGv4hm8r/QRQ+clZ0TK
oz/WkeZmh2pcwT9con9wAj/S9hgdHxVHr4n7A1H+g27ZJRvsaSuGctrACru96gJT68IzORz/HAJX
AEkq3SyEl1TUvmS3g+SwIBA5aFI/OnvvFH9rVg6+tH9LT3WuXRu6FPVTGUurLCkYXhDi824tznLf
lvk++8uv5s0iDwXAPe5JxxjVYFkZwrTGs6r64kB21oZdAPp7APIoWU8fZMK9KEi5XxqE5DX74HJO
ePptoNuY6tIed8AcpQGQf6wJtAVZLSnV2nm87BBjkx0TeWWUyeTlTTidwMsySr+rk9G6TCvuzG/i
YOg6rFiEcnmzSVUjrgv1+f4C/oQltimz77uMdqROFfV1b7vx3bQNsal/cWevtg/qAorjO/w6hWQv
dnOfnJ5PKJ0qqX7esMhyPrrPtkTad9v+0YOTibeA1SZIy/XLeIxxFqwxVzI8PyfArHngZssyQaH6
poonUWYtUT0CTtXEsi1OGt5yECxK7oAEReja/KGz29uaruwH+loNK9HJuJpxRDCseVY2fW/4jUCA
I/z3KNt+5GMLLSFZlD7YnH/RTpSvypR/v9spl706L0vUXz5OV3YIkB8YrIh3RjPKDfHvzUaPYfcj
oKrdIkyf/JPzwztCpZCPziaJPPPvuR+GYEvt41rlKonc5txduLASJf7xnGwFYTu6mcqUAYJ/Oh5c
JKRy3WHT21GqCSVOuFNogW5pcnpeBY/SNMI8TuFQHPOuxl2C6nC6p7BjRAh4cXWuQWNOad7huca8
hY9AlUPTRSIKiFuzXHe8WKj/ULLoHGmYo+30N4xc+ALh4mJB4AOiSa/h6/j6OQYeacZ+cgEK6fA4
dgQaFNzDrVuAndi467N0mDE1rY+3RoHWhjxH4vszHxqCipcaYZpIwoRu3WJWgqEXRoxHFYBCeDdC
LZSBnyu50DccTSZdUTQiVFoCcUgtSQWxiVsfBnf9mMpB+bQGKDB9cPFwMS66bMsncKf37I3tVvdS
uEm4q9sT/JaMZ1iSlfVU4gUBw+ZafBamFr2Z/iyOolJTqgKQrcI5cH+gigGq1L3ZVFnL8lUCuyf8
rmV2UVVDgGHUSWvuknydZCU7WIRSEXTQLTu9qzXGMLGKXu5cccTB0dmpallv0nbeeUSUt5STr7pA
DyZYUB22RWyDJcs42Klf0UN0LmgS10QIw+eUbWNRsOL2DqVmZdoMwTnwESofSwTwdnYdY89gp5AG
cyCoYQCA7jlofgLNogDz87fyNOZUrkIwZ6CixFbGUQm5RNtOlsa3a44BO2BeztfzttR4FeB03ig2
JheIB7cyjmYMs6C5/6nrdcIWJnE5dWI9UeaD7ouybfibRgAyIdb612Gd0v3zAST5bzYjN878LXnh
+r6l1oDpb93OgxPN2b984IW2sla0Fenv7GY3gdCJaSoIe7gGiWRn6EFCguvybb3uIk4yvJTL+2TI
SgUWCPFozfH/KuifafbQm2iU+02Fps2KWOec0czy+bvlVfMh0k7wZoujKGADWI0cLtMxd0HdNuQj
+LbJDMxEP7JQIXv2ZpdxWRvOO/svWTWwK4g5XXcdEGINkW59w1eUZDVHjO+SMKkzUZa0zaxw7kf8
xCe3ph7cx8ZjiEEQS3ZFs0R574BeheB7hTNujMlPXq5zBHB7CwsgXtiEbzf8/ltBClbpnl5alvCu
t5TCU48gvL/1XD7IESQbfQwXYBJ9Z6TCKnvTH3lpORamoNhoCtcrrrgBJFTFZfW24s2B/xwEesJg
hwlkvbvmCfpdNoMXLMkGUsn8fzsBDBdMmzEbkm7XZ7mLhZypGo4ikDtWNYsvsF08htGAUTaDD03d
JemmjbGtEu+3QGhcMQYHZ5nRyA3E5gig4ycV05Zkg8uD4pdCyeYO6xUeeHT8kVpp5xsQQjwBK+4H
6/NfjyyztkHgtv2ohw4oWS9vxHr2WyTLp5LfdScZQRsdsMXKhVJLFLgtYkC/13NlDZM99egw8s32
Z1esmJfzIjQgt8iiji7iieCPTTWbcndQMT89wNL4NDB0kjNtK0iEDRlVogQAexAB8M2pw/+Fsc2T
x+WMIKtxmc5w8I4jSzDKmrcQp2fu8vL8VbDxoYfm1B9TsN3HPFKzuxtTI+vi011R0CdgyOidpYZf
JzJB6RU3UnB3C/Ws4eIzk0tG15JddNqXDLJGyX0arhOM8OlKm50KqLHTcKtVOVMak5VUST0UGXBC
1SshtqeFo2SRlP6KCXG+W9BRg1G3qkrLnLs0cLwmQbgKVOrzf2Hy0IQatlLx64BjSQI+LFsAxU0q
DwiMHtc/inXH9kUDRiw6Tfu6M08xozb0cGzZYEE7VT2dHj7WSni64PhJrOsO+RcC3/Cd0jRRMiXK
adyQWZREXfrMWpKHsrxeaPh4bBmpqZTDaMdSh5AEQxkgxHUW0RrmLkPNunlKPTjkjqI/pB4PcW19
X4QiOYWEdVBstHH8VXEokuvoaWjYQnmZBSBAkrLXrZuzM9d9Yowc4P5XGILB9UWZBxoh8EWuTMG0
1o62qHO73sEUIDbgq5RP8cRuThfT1MyxL7GUg9Cim7/mZYAdWvsXjDHujG0zXxoA/LkMKi/hFH/r
pJXep2mAAA3Ar4TuO4BIS149vsUdTUlWFgH8a2w+L3JYuO7+Xrw4OP4+AMaQdSLaT5SoGXNfEDeG
mksAShz5KD2CBetbz/C+PIto0dI7n2T9j5QhmfTx1RZzugrL+GPKlNvju+qBSk6fHBcmdX28lPLs
3x1B7xbiCBZN/7lzwiFz/c20zvY2SFUa6Q3PTbO7eVA1Vf2AclDmg6pfqT9R1lV2JUGFdyX6zR9O
K37tBKN6JvaDnbKyf86FCoWySTXD0n6snlyyboUQXlD/VAVHACXAUO6bV5ZlfRyuPW4Swv4ZuzYd
RHxV9nEMjcejKfqqV9oIz6oRK8rOYC/XiiO8CwrCYCAR0yqr16P+exduha5/CHcYV32szrPzmiyG
+HJRIlK1ezZPZCbxThIA2e1rZW26D/S+Z/fqcRFAnAshgnFXLsETqv+yPQkh5FQ/BR+rKyy32Qtv
STPbKiklzyOSdpktdTUxQN85MOmOk++bol/SaGvoLrUGjnTiajvZ2B76bPSwyvXL75rJB4nVzraw
rWRPyyt+fXiW17HuoEYVvNsbo1cTfnAkuH8LqD/a02lxQ9ddwm9n9bJqgElosmITmHwlNXtfE79s
3BWWMBHrbbfgQIfdMJFQ87in6Z9xmoO6yLu2SQzVkxA44oCmNTj7f/hyBRxblUzehZIuBN0ou2pW
mzXDjmsyqSmut+S/3JLtMnx4YNeCakcfbbX8R45ox6n3ITunHkBtQlJkO5ZocMlmbXRzHqcaJrQB
DiHiSwJObn9tQRfYmrThllY8a8243A2CTQoe2p1/zmCBgpbGQBNk/hDeYxY6VcF29RetXPIXcBg1
KZD/ElryhesIxQTl4+f68Ofm5twxaNRiD3/s9CGlBGcN3gUrCJTa9qzmXY254KpHJtTIHZZot1hz
6Ep6bPpv+iIoI/ntp2QO3nySfIUwpTVlrUdWbcwdV1IZgJ9/Vl/bkWG2yidrE+UZOc4w4QyXuokw
pfjrfWEz9EocPzkPxIOlnESVeHfF4vB+MIMbF3qLGMPiEzWxIZZbBMCMWtKIFpsL5TT4V9FBlko5
LY+6RMufVj9uZj9peyCTGSVa0GW6sspMKz7aZfNALF/CqVZM8RkIeRI3rbnrkZQd2zfV/EeRpwvZ
spdWLh/qrn4a7eoahTfymD1N3sk0dPbnF77hF4+kWqZSh60vzdnKmJotddBAE9TlZXVD/acz2Vzh
njKA2LEy5G0CXHtPz5lLxKFrB9HfJvAf/J6eJDqb5Z8kwvwnXshkpYsjaIdmZg6maRC0KyM4sP+4
4HbOB0mhO0prBsyJh7Xkpv5SOETrNIc+fUTwjaQWrcY1nimoxua7h0/d3OZOXNNRKURD9WLfm5MF
/c6QKsgPtPlKOGYwmpaXUPhkv0UfdZPUPdJj0o28uP1vtePkcSNKpT1my8mzP3xZ5YHTynLAQYhx
SCtgn4cLE1s7rbtW/LqACFIveNAOIIpAb4BCyt0lDbM9ADqvNvdw3en6/fvNAhATN36BAuGuiaZ/
SgmLA5lSwVJGl1As1no4gVJF5Ia4SVGCdNiwe2C89iSuGOMmyVxJa4aBTzs6T2AJlfdDw79EL3Dn
s2A7oBLOZkehxKUTzScCXVpURwsbmLM3Pu3E41XPVGCH1QX8gvdOYvgWqysUPy9LEeKnZRbWkEoa
6vQtPyFSu0PecQcfoxoRngVpN1wQeZVRuKSc5A8NzP+277mSesLTkwGAUTaoP/UTtDvgzxuYVCFQ
GVM1TUYxROhvuLxQTo8mHJPxz/qBbOGWsJqYHNhEdY35PV7fcNWCgFeKRafYa5CPDxSQhYJaPPlb
SjRd0XzE2FkivP5x7gQLskChjlN3QBOVfjnDCaPbiZJECghwZU1rRlsO84mITx/xPQcZx0LyfUzR
FT02gHxla2hzsie57MLdL1bf1prTak+IIiPZDeRE4251WDtKe7TZ5svddKvbZhD6uK+VzA6AstL5
iXPWUxquiX216SxE+jbgZUfSxMdkE2tA0Hf5TP3CgHxtrasVIiC/95zGcXefXCzaTgZa1YG22kvm
VMUhB4mrv5YdG47AXkOqRDUlNcj2cJ8Mx+0nKyQ/E7VlxqMe463rfAhNwvaaF1BRkkjir0R7LodU
1ybSV8jLrmnnDg5oD/48TLWP8rM+lcTmpOnayag+Rdek6c9ZGqPOre/IXCudokzLEBOcMrcYEZjT
QMRgVqBxAu0UtXRLBSnrbkWT9Dsej6RfZ1yVp4jkJeqgWOfvi3Mssds1GEHR5yLkHzRmF5zX6Wv2
1kz9MXCG0NJTBoXKf2QP0YBi7y/SWAJYmanSNX/oAwqP0SfjPnLfXS4FfnsaWA0RQ5oFoTDna4pu
v8grOX8NHZC9bkkTI5VOnhRH98nb6jVXPrB5XmMifUGvMnZONH0wwCtz2ob60JTLs5miGxYSVxAM
kxiNqUCd6Z/McS3+EIdVyT2ZdBklSuT3YM8nwU7Egf+6mS2aNq/uAZzuwQHdSrK00vwnKIdlLfOh
y/qeH7uCf2gvg3hYPt7HQC6pUo+a3pw1IaBq2QCneNixchX1fyRThgHVoQyH7I+YmQwvpekgNAAm
KQEsG8CEg/GHXzXtLl1lBAap9gG0PSici0TgiYMMLtsyB1HTapD5YZi8jmdYr6kqYo9ugUMbzQlL
1T3tnTn8k0mICQyKuI0mjsdS+xRGRgiHWOIaeqLN6xKTogdAYWg124ZdJ0vq0yWMvtpe4PF9SeVt
s345iai0OG2tMLiyT+pjsWegj2XSXZULvlQ5jZXZ/iQUukjUZMaCwsbEjxgvyD3xFE/sfy5JonI0
Ay2Z97Vj5qfDLZQxcXZunfuWy1bHaGsFCbkbUsczhVDvQTJMZ9wIy6C2JiVsMBO7CHnJqEz/trBp
I96cHfIomUK7xHjOK2t9LMUBl7WUw4UZev/B6xOeH7RRjwTsxNP7JNDn91pPuRdfsCspSWVVmmTQ
IoE6KWXveKKRoO5cOglSZqIOLYt+h7NvNdxDuCsV3d9rLfE4VKDN5Zb29KXCUPThjSYTnTs+j1mT
8Mr7uno7AtsKFIVae4k5HSj8XaH1gF0IprH0zIJbzS4yyTX09aMPHb/O/bmlTodNcAL90ieGxrjo
3LkB12Dla8TxS0tjgk+At6L9GidfZwdYpFaC8AyRfMZ3NYyJ8vYEyJV4MUkehz1xPDK83Qe+GFVd
OCGHjm9X3rPLm6ykqN9npbiGzAPzkaZLp24n/5y/AtjRVDm74yJbzhwRFzSG+tEWzOiB9UJrnqLl
yxRBsgiMv5XvugxNyMy8O9j4D7baRTi9KI8Oq8Aa5skxrp8H255tKcDdTJk0goAq2znApREgDbPw
BUsb5xfRokpZfc9g/0KYsPVNp3u4sTDF64HoKdfO8gGDKpT2T8bMDzw7LOxjo6qmaC8uvScmPaJM
vSI2cmp3zKHOtpbnR2irll1m+sURry5PL0s52VUWry41Bl9deIzmhnONLA5MBT53KNzrff9FTLjq
tqssGzeXw5yxff/6YRyyjQ778TlmDMxhzkdSgARezujZTh13q9nQxom4Ti4MLyaDxrRVjR6EqOqa
Mr5sBnOhr7lqEPvvu9nIm5mxXQHs8KNUNCGF5kzG60uB564TBLXYH9Mn/IeNuitzCf1extpO1pBG
3ZmO1AZJ3d3C61aOCbX9JIJ84AteHg+5xrGaPAVCSlbfh3dafF0gXfaSYcqHo9+6s2uIJbz0Uycv
1J8TPBDLyxBaYgEYFW7N9r2dZZYuN3w5LWz4/zP8JZpG1aXBIolvcxstWwqlkLmrjr6F9tSJ4FlR
9eDm6mmTJ976nl7RL1UUUn3jebqb+pioZLe1gq13Mh6sROUH7F9698egk9b0hzjKHiQ4YM3oY8c/
V35z0xOarEcXc2dSYralPA8Z8mbdRiSYZM/nAr3VlX+Gh1GEu0EKnl6FwlaKalAZszJ3QTEwEA87
AB3aag2yqJOlTNbdIpE77V472ED7A3dlkHDc+m3WTSxdVzv045+zcvJyy5Ta6Y6wXDYoJORBza4S
4pbFp6F5kL++zB2OHu3KgqSm56RvmBvAiaxSzvRWOfwD4t7S8MhjRpwUIaF2bPrjJ66T8M7bg22l
82PI9Hkv01F5oE6prI/kmtrs5E9EtJoufjGpF9/Naywv8qSImSNoxUpSvPTDCXeRiqKFepbM6Dv0
PPZZt+YB+IebLKvj5xwcB7U09srPHbnQgKJkr+9FLJ6fnaHKZG12dciziuWs3rtZtL3ypQKnkyFN
5hVJ6RR6AIYmnkimBhW4EjPZDGMuZ/nrJsOBMHM1fT/u2qzG5MRbcfsgtC4Zn+11RN/ke3MbrK8E
g1P10w+ctxUUpwVJkqJMwMk7lqLudUsDrV/bw6JLQ/UKn3iSqvCYkXmOgRihXVG0EpZVo3srcBh7
9fxAnbcB0R7b6L8899hQ/UFazXcQbjxMd8fw3oYH8euDWZfv5DmSCjiemrU5Q932i+qXbDegGNuS
8YriaeMl6eIQUrk6Pcg3dqwhwJI8Vkg7w2+/PQCBnMD03CffjQRvrU6fusZDdeYgMYWHU0kyJHiC
VU6kvNAGYZoRVBfprfvPX9VUnf4jDKJE1F82M8Mjb301kzVMuu7uLjkrTUzsWSSOXLmFbuon0s3F
yjGZk67D6Nt+eRI2QtE3a5fWly8NLu3yEx1Im8OeE0sadUXLKTOBFhDNku7hXw+19xzj3T9W+ddZ
Lnbq6WkNY5UzIp5haBDGPx61zjDBA78brobjZkdne8JYpBwghMTPvCZFqWQB3xXVbEEaYJEP9zZh
9NvGW/oCj3cuQvPdfH9snm63EJ3i8wrFYb1ZtMax+gMQCVuXt3TxKVzlP7ICMBVGHYbFcSIJQG7i
XaQg7kRwgnrrTvtve2INPAJbMaAMA0IxBsWDfID8FhCsvUtN31ofOQGW7VvnbDVUVS45RJCyU7Xk
0QX8QsMOm+pCdWhd5JiBGO4KT65RGkhX8AzMXBLNRfPf42LHhzTm04iM89dlqbgbwjndK9O6tjz6
8XT9SVSOWlzfivr7qQwnqL/j5Po4LULR1bopW0MUIhL1xeIRKBr3LCTB4AlnDCuS09SAN5R2W1yQ
qMOwL3DfZ2sMhRejp+vOZzTZCs44I8OcJ7sFLqhT7cysfpi2RhaGu1PmiEiO30TcjsQrjvF0gAP+
KeYBQ9IU2gHmKaozPgFQZNWma3k9lTdzO2BKgHYckRXIqWJ71GoRv/mNki5W0tQm2w1DXz4QJqGB
8iY3YTKHgwXpq2yhUjCgkij+DK2Xj3vlPSnGVwMtEI2DOi7aYJTd9PjNqdFfG+EzvfgvQzr4sMqx
sQCAM7/+20zygjv+f7JT2RN3J0fmIFcttU+YibXRUYVXMDsQoFUNtpAfL/kcxt7NXjdAqX0jbZ/W
JvIb/PLtYcAiYKz6S+vvNjdUsUh47ra2tqH8EPPrPj0ZVq2Gvp4DFamoz5X1ZZs5MYLom8EH/58h
w1bTW5DrDLMYODFWYVZqvH05xE84hyzf0IreJN4mjEcpvw++iQzZq1joX4CdPwvXZnN3U289v+Kh
7NG/1P+f9h3e1fvXn/nBEZ8LRXFYF60NJUJz5CLqQzXLDAcm1BbskCUDbB9QvnEWqQW2G4JDtZYq
qXle+naR64zewkh9UZMHSC49NK/+A98VekjvqsEKwZ/2wyHPnGcVzfzO8vGj1ecdm5jwmIJO7+Up
Hvhq84mUEUIrTx2HXQNPXkVWzfl04C5jvzhh5otAmpJlY8ZuUmmLO3mBnhIWx5v9PBoQq6AjHBjB
3GdS66fpzpRi9qvHpG0EGNYdhxnEjLtl0oU+JzsZ5uDS7T6y1krsUQLCl7G+Och1iSHT12xMyj+e
NuGwng/92TO+n+LKa4/D3DjjZgEbFgf/ZG+wcDf716CSuPNykxXGDSOYIbjImW8vlQvZ3Ol/bJiZ
N7Q+q6Va7ZEJ4bcPVOBqTT10mPA6yWcHR171IG/9S4iEY4fpnKHwFVO/c8cRAudecQSIFa6Dj8nh
SKuPZiByx9NsxjE5+k9ljFL79RC39mQrX4rK+GUekzW4OF4DhPL9BG+PoioqR4tdWucCy1jG+EOY
6N/UiL9QDy4NCyOjCNNLqZv9+zef/ADd788n6dkVE6NqLBwXPaHK0Z5SJbqRtKvmDLKkG8je1YZZ
s98AkcL8HN5V0zIV6v+8JBaPSsJQMpDIo1lLTnnIWO/xgSitD0kMqgjENHzDwRpOb+xzQCUTIJQQ
gaZsNxzx/pvbfYXUONtW85OxSzsGnJeuuzJ/5oQE5QMImTxlb5hYB6XCNm16X8l4hh47Pa3Es+VS
032ePUN/VWfmX3hLEZqaPRf9H5izpB7KcWoVweXvnnQgc6zlmt7AeUEJysYyGiSK8CqXaSdi6tsc
Yf/B5IZEJS/Llgekdf2NlBTmzwUNVWngWj+AOKZ+Jagyp4HbrW5Y7oRX0el1RUggJPpdixccn1y/
syoLCy91DtnbtOHV0BjrSkP611n90G6tTynzdZuG4Z2YdvFMxCcE7A3T4kMWpwo/H3Lebvj3fnwF
3jB7i4fkDI9SPcQzZYcuq00Opvnm+TIgkMmWlCGHFTAanwaUd37b4DhgqmgO1wZUC3Ebu47biOOG
TQhKxrJNwVUU5yToJvs6QY+skFgm0xiDtIPNlc2lrSlBx8ztBW/T3+UIOmxakJTWb+FEWUsVzRzM
T0M625gh7rDIGlCARmChf1mfKKSzgn72KBdCDLsO2oSKClCAhhmUD5psHcdQYFHVYEmBmJXI02Fy
8TELt0umNyDrg7QrEO/1cDTN3DFMlIr6d0fy0u7zXe4GD5FJVY95NX02wOPtlu8lD780Tzn5iN3r
SSj2fl0G4YgQqQ41Xm6jOOXMVpiVaYJqvnQE76WtW8Yn1YoY1HaVyziVdU9Oj3PY64cVC6P4Q8sP
+AxGEPgo3bUHTF4F6XY81/cOYdG9+xoZ/l2rO+vF/oru6PZ+Wft07JdUwy2tZ/oDMkKdohi1i8xp
uAYtIqMafDLJ/xc8WNmVzxhj3BElYJgf1us/JIRtKQ8S2uyV4QdyVtAEgM1i+Cpr0TEkgFzl85Si
NyQ5U4xhI5dcJDFJJZoNVvNseU7X9VEst8lANjT6Y4UuJsenbIVyl9I3jbicyOeCsQNR1LBpG0us
O33gBd7vbXJ6gQoCD4UAi3tvj2sa9UcUaJ0z5dOuZN1E7tC5Zy4553xfLIIJFQ/hSUXB9GAafhq1
75cYwDs8S6x2AJRjA5lMAsdZkITrvjWlAvBHCxW5GRA+z14OD6rH9QWQ1d8dtJlpMEROdAihMGeW
HhFJsV7RP+G8r1BgFumuv6ZzfjZbx+3Tb3ViRKIGqBTEaGdHJceDGFgcec9RdNHWcOBX+hzk1AE4
K9s7U35WQVUSm529r6qxA6tpeHtKHEadmUoMO/8tc4BF84ZQ5DpIYbb/2EZwn5fGXJJWNCBsfyD2
essp5U94aFPIo2bFL52yliFT3RB8Vtk1Ps5I3TS2YipheCrpEe8gy82Z9YYV8jHlzKFsUUZXeouK
Uf8WWDELCSprSL/OWPOzf4/Je7iibeDJkcPGjfNGQkmGJ6uQvKCvssZHTLy5DebQ2PK3norGV4Rp
45x5So2rOfss0p5+mJtYImzjULufkM49c7zG+8uQ3OccGhXrd13K57HPRX903cxIgYjLQtaBaUj9
7OCfKHheLuAUhVEyW7Tz1VOUvZHF3DOF8HTGgGHuwK7NE6JssqbGpPUwnsPkX+MiBJwWZE1IaQAF
WK/US6bxW8/mwvzF+UTCXSwmwvN7aIKFeQ3Dqf72uhVcQGO9oosfEuBKEOOFq1tU0VJy6wVkBw09
66l9HlpzMkRZeNnMkOhRBSrVfpaFSl0IXXHagzI72Y1+jgs33EWeMpgD5uy1eQFXGYBE9kGIWm9a
M8qiHg1bJySzVNHvprU47Hznu2lfx+Rm/6hbL04tNG8Y6v0UDk56GjzLQfvgS5FWAfAzBEoQ8mK5
QG8QiPNYueDEIMMnFtvRoNBvRu/Nwo62QHrC81rHYYW4wmL5qVCsiu0vknfwWMeVs6gCSkGMOKhV
WM90qksKyKAVEJDgFUN+vpUMIMR1IyxzLI3NoJnHw/6OW6qhGJf/nfrz0iTmL4j0LBPnGyiuKgUP
AKZ1Pvkg7UW/+rTZXp4RLj/ZRxxU+Gtd2iSWBuqqKkZB0EDakoKCp+0yibCN6jZpsk98Vi72hxCT
xFnalIBxeGeauMDXANiuhrb7b1e4wj/Rj7Va602MlxbLylkDD6WL9V0DfLF6iCpPqfzacAMIPuLO
TfRkpBaRsLis3Yfig4/VDvm/KolGBtM2A2BcjwkqCRrkmRR8DJUvl/hshfFRtzv0fpJkMi02XrEY
dG+CbY6ygxo4w35fmtCJIoksE9G2wCIxwuuKsdN2CrgBEZNQj3+DUNqmCaLDTY7zS27t9xcZl8Ny
RhrdT/LjhSuWLPc35b6toDihFlJfAiEpUywXbit7HqfKTM/oNvWmH9zBHgrRXLtLsbJPfJItxMJ5
TSzb+i+eNXnxH6SHCYL0famWpXAcfGTozbGN260+GsCoNaE6ouKr7fYBM+0otRSMt5+DM5ZMzKq4
mJvOAan2e2TbzQlm72g+9m11RxWu77j3+jhiI2LPv95hsjbLH8VZLDkPEQoEbq0sfs6zoQOBTYiI
waTy2yDGIdvSOr7aa8sq5W0ltEHKPwgVGtqMLm0IGTkBAPx4Se14MRxj2dEmwRVyOHBGuEK2ACfc
Iu71MAb7V9H9Pv0RP/4VsIU0me4DBPZyBybnMwEnnvpWvP17BEWbKAvi4KgDXXsP2VhCErP/2qyF
Iz51KPpOlmCxm43+FuTN29LvfNWNguXmDXucXcv1dVOGW+C7/8dviJ57Y9vwQNatBt5ko8r1eIno
bnvKZ6zpZQKc78wOMGjXMCuEscMWjzpt0yJQ9in46xDVGODcO6JpIb0eCnlvDR7I2m/I1N/FdWqp
4BXKcEcvry3LwEtOx6kzuTMb6g0IN1XOskB8k3NHf5LUZBk2yUXeYw5xH5gAH+WImiOhwTgluIxG
8E0SEm3L/ABzbDlRJqcGY1BIYiOwISVxF9dpFro/FTkuYpb+gpyQ3dsR8Ql6KBCgJuFIddEbiQdV
o19LJ1Zkd8fidxyRoJB63OPcdBArslPPeAJRylNBCnixGBtnz9gAiCIzpmsEnGew2LSgPpZFjjfF
8dHphLew0NZad5h8EnMgkvf3L5h0z4cesVOZg/TzNjO19ZlxXiGwZDUR6sy6+CQGAbo62UuDpCNU
+sIt8ESZCfqiZkq/J0YFV7RmgAKGiHwIHv+wrk37SQIXfv70RGLXYvbC7hl99saPElfknPCvwJXk
2g/lbXWv54WT2UHu/YuOMW7yMVeDRQdPm7YBCVKHYNtouRXTyiHFQHdZM3NDGfnuDnK444Qp9xkL
iRHVF7tTO38LoPoxc3eSvNIBHnOdFMUMih+6s4kQfQ3SAc95qJZ9IXGV/ztExLL9oiK1JP+rX53S
mE/mpxhWT0kkMDbJmFuES9JFeRs9B0hjxpOPIGHYv+m97XHlBW6Jgg9fBvbfm1Fs27UP090F5qZB
T+/BY9xMKdN9KAj7IDwbXST/iGhJAAHye2m9rAX7hn4ByNKKJUAbvLRiLfZfFGChbC2afu2Cfdja
3blrPH2mH2OOD3VHnRZfggbg8TRVcwhY2XCEjfuT8FWaQUs7fuaL7S+yYMVNiZ5lb+evMdl06oT7
QnNB0QcKzADBqLYazY8aUismmCq1/+wpYU8Jtp25v69LoYYLp5F5bcs/D4AplGKfnXqWfQ69imLQ
n5UdjXbI9nyvm7fK9Ks/le0mjS0z6NQMvZZmCyg24Utm8m4C3vGSzzXryjj8HhMSJufoC7/fFXeO
Mu0wXq1ocVlQQh7GdH1WJjI4x4vVTRPxYzVZLfGKa0sg4won+rwM+EY1PkgLUPdgMlzlaAqqvlJl
cNwspzAtHL4ImT4kA4Z8JM4/d5SijOJeQlggi06yIg984bO5DpNPB+Te779s+p6YjxDQz63+S7tf
+kIymY2qkdWwCmsgETjAxLNZwdtl+2ic2vZon9g2i9lhTp4G9pRFjeUvn5zBg74b7vFXtOPQuqQf
5BNXH88+KMrAHcOSLXXiJ36OqKneVg0tjB/jUoM7seIks9OUN/f+CQeAJda8Wue+BlftE1hgvv0h
pZxrCuoJSAisCWhHz1594Q7xHpuCJcv08t/VIS+XOQztJ+PUQCxcARRBrKPIv3j7aNjItUv3A2KG
PqI8WLpMLEmDtuZ0+XxurhRSE2k9e8XGTmpgXN67TQcqJB3p5d4d/ZGfG8rmNtO+jVh7YQvvZuZs
mS/Z+YlMXHWBj13uzlHa3m0fPwafcYQErUzezDj6mgq66bYw5gcGgDb7mT/DftNekIVycrinNnxR
3CL1kSO865OYnmhfkPkQkgQBQG7vPoxldohyFxfBp88/Nsi7uDpmiqHSW8SfFfUwZFq2tzKMrQLE
EUcH7WZ1HRNgjdmglfWlSEHw9B+KyQDg+JBldqckTzxp0LekWnZymENgkGA46epy6M3mLVS4agQB
5PHIhlJfk3cPZjciaO90ylPytaQwQBcqGU4BiUT+Xaewx8XmWYmfnwKylpnhxswV/Jj0boYyCXIT
wrBJCYiGGmL7B+IB2YWblFA3cr/WmuR35XJpPNe6/cqE3LiBWl05DV1omeM2jl+VTrXtewVJvMY9
vNWRr2BOZn0Oah6iI1I4P8gzk5I9CBe94YWZH2vo12Vwi1twqhzZduilaw0lAtajK7OTAvb6obMa
pGOytdY1hZXGKRWBlFSR/5bQTtFOdfAP3huAwcpaSWxARnmmFNdmWjODZsAqfc1B9jGrqp8FDjdv
admRxJ8Q/X+FcBKBh0Gksi7R+dUInfPyqBJrg5hBbJh5oilFtptGOtrNIfTp9WIcBheWeniJqTqq
9dt6q8DwaSE9cGGOTDpTx0Iaikth+3VDBHgmPRoSAgV2QEprR0w9jvIE5AgYWUkqwoWBp1OkYan5
yNMzn7iIbowp5EhsUQbXm5oD74voDEoag7nKpeelWG/7/i1oCLkm61zZWyc3IcxMz0jLUce2/dJM
kP04Z2RQ2lzgqR8Iyaowd1RK08/JCY5v3cunWZdpZvDjXl4h6HzxbqaGVlDfXhm3oZisblbGm5Sp
PJaGuFLmyOaLuuU61cOvwQRGgqa5XWl7dN2GPGY+g+k9HE6+mh/GtDEd7Yv/dAr3K43QQuHbszNR
HtydLzHwCmZimuSmGqqUpX+ZEdtbjMTYX/an7VegZNY8fkB/m150IFOu2Soxg+Zu+B5iF4JzB+SC
dDsImJbUaqgQkikgi5msZZ6EFJcp4OH/nZb7DQ7hdih4/WvksIEn7Fz2Jq1U02Z6FHG+FOkU41rm
5npcu8XVE1W8EQYacHLBJnbiObvoa+AxW5eC4H77OuJ8QrK3vhwhH7OccVpxG7kvF2e0KYappG/p
ghh8DJRR0CWwhlOc3BvB0cfrCXl1a7tGI7v3JhH8SA07ZhTnn34O2xkMIaaehlRAvloVldasDYSb
7fRPRmpYqbFuLt5Twfjc6FR1g/lkpyb6VubMFYGutzQ2rEmBNR4hDHWn27Pt+GiG90fwg57niwl4
8Jrd/WA9AG1BQ2mbRyUvwbsln8O/a/2OaEipsNeEGiqKO8cEWdVuT90X03phUvDmV3HUtszAfpnM
DPGJDZnNjLfyrkuVI+2Ggk4FEGGPCoAK/BHm9JmQ0IKo/KTjK5PHtHNTVhTMEDOmVRjY5ZdeX6SE
UgJtHT6kU/2ou2U0nXgcuHbbY9eBbe+fKAlUKmBGGvjY9Kq95dI+eys7U+0VHsIf7uVyk7TrB7Nc
bzQDxz+gJI5FDb3F6Dz0ESrDV4HM6FYgI7Y39JAM3eSUTNCFm/p8MTxnHw49/BB0gXMtkOm8OUe2
pYMsLq4NQTX4f6PvjQxCqCoWJ5yVSvaUWMaZgtyeEsPuHRj7wmi8K+NnMqR9xWhjitPJPFZWwzD8
+SFvyMF1PaArLIrYGW1hnQZq2U2H5yQlpXY01pGA3je75KtFRNbQmY6naE41uohJsGViWVqyPvfo
/OiRY+2WPiJpwnbafgdGeuNwTJ5rSIEjNnhzajfM88MtRqMBo+hYVhL1R9ulwso7OVsPVYjNRVEB
7aEojnP5TaA95+3HUiFcT+Dw1z34JBN5cejCN8GruAUIrqNd296sA1lnIXZnNd63LTkLAJQ3ftC6
xA7aX7oPalpzpVqlcbccrPYyuXziALeQ3w9LOTKZytWP19syRvjjef+RYE3oblhiRn/EwXhF49Qs
lVKpWQivFry1ILXwbrT50qOvyPu8RzQzDAjRavR0vQ0iFv3FC5Dn1ZQIjlvtiKrWZvsKo5ldtQ2m
tCzYJ0q8KdztwU2HeM5VjnnN+ey5MO+QFFdHuU4j85ZG9aXHR9RquZjgeWin426r3wp5J5d/95ju
n2rgr7D3yMSfzK201FWmELeQTEagsitvRCrcnn1Mi8vzkiihWtBiZ3GdrgYyk0Z1uCCSxnMNn5mX
kX2nZ3LxyBYJnJ9ywjj5HrKV4onajFGTuTn4lxEG0pcBXBM97cy5/ZIJDLWQVns5dw+zUTiRTQeW
E6bCTfHNOtsl6//6JZZOQUS+fpI88eUlEk4oVffKaF7UVoyCsNjqzDuG4kL+Y1iWXhY01jyPi6uv
eOpiHsoSEOAdU5f41sN7L0PZsZQN6hVNRkhNulM5OBefchBZIwc92gY1KLVVPQxgb/dwucE9SPOe
PoOgPWfQgs4Q+/UQuMFL2UqMlgKOLfmFVmFyjgabd0yrFEPE27e37qYtiIyKFPMgGCkSh7Bq4moW
v2oZLOpufK97FCL6xksyhJ8FrlQIpUQE3pRR2t6ml2nI91Gasc65kYsQkX6At39aqrMq7ldTA7ou
i4LHf/qfPFt0b87NG2fGCKP2gREnD1airRQfQcYXifuVtkUkTgIyBYV7F6XeRgZCLyTz5Bx1osXX
5UbZOrsdfqz05aA/C8aWVeXm0TXd4iQV613gBM/eM50lL9LOorjDACHapsgsOVGK+ZXQJ3ZKUG+D
KNrBYQSKMhj+8/PW4T6co5/Xo0OnikgOKjFD3PXbaHVYOq3Fn2u7ObT/FL+jBdTVq8PyOLiieGrr
BbQnruJ5wu4p8weMQ2+njGjguUJ8+e0sCyfXv/iLN3qEPuNWgDox5wOFJVwfZ0CJidFTT8LxGNWj
Ud1MWsAhW7OKwNNrCvKoUM3zCj9VQfZT5zmVWOYADJ4ezy4QClN69C7c2gqSSjJuzOE3ej/neAIS
Ez6ePRC+f2PItJwLHFVu7MdBGfnULO6C7q7erMq4IazAMa/uy7iboH+MQmZ8/rjnbBng07oT/id0
Nc52CMAdUN7NEqRCR/GQxmnr6jk5w3U2EDYIJfvmeR0I+TKg1uQ7bdeOo9tVcMRGINFUDIJ89nW8
7i7/Fxyxu4wQjNOij9QRWQGjctmAkc+dB/wIHuYV53dhnXativk6A8Q/oUx1a5UOvb2KZC0//vKY
tCn29Sqwy26uy+eQeyIzCDZ7NEVPLEBEN1u6pfqym4CnPZGamj1d77JnBLaKiX32lL0LNsut8Uja
eC0I+EwTf5L5kHOuc3c7PpT3HrHrMN/qu4MlRLzVNf4ucsBD96XisDV9edW4zaCAG0brMYHyRonN
9Me0Agy2KQu8TlLSJvmR/33+z1xYAkT8jEaHEo3zBdrLoBfXyVcetl0rtK/J+L24dm/exaUq0p4y
TJfAUagTIKlvp5x+A5jQHJZuQzHRrI24MjkCC5mR/0kNw3UdpldY4AkMEL90owZE2g4bJnHhkIWQ
D99bY17fXWQVr1laQk+3yYBCLAKW2C5JTBCJXG/2ISdXsds2j3WobUTTH+Ix59n9ZmtuC6nIUV/c
fzeyzFWOyETivXxPZrAb4LSeXRKRHhfSJSlHDDyFU383OQ9FQfGkZJxEyU+XMqB0tNvgjJZJGIvw
63YH1x9PNBQ03Ds/t8Q1xE8SArrxUGluZAm8Qi4cz9Pdj9jAhyUZ4DDPeTPBm/59RJNag93Owch3
kig+ge3UJrzNvc9BOtVs8IOr8FIsxEl1WaL7+ewBEie2vdQUWtxZgTxk3KVYN3YWITgByfbRDCQb
4y7/JwE/ggItAvQfuFHEDNkHvEdMwGVppRDGARraVYs19lzsVuyo+LBt/d+cH6mfE5yqNaENC22k
WlysbXDMqeygg4lFCYGUjuSPPKm+u4ST25YtTSxsO78pcK1E0m4z0GUjt2l+HqDw/GnhHyOV9vmA
mAi7MEPbZxpmmb212K8Z2NyLW6bVyZITgetKZ8iCUPnUbSfXdugMeMrkDDk8DscX478mw+F6zG8c
V8TlWecLBcSUZSn1SWNH8xh/wu04TKFoaAOJWwEgnQ6ME3Z3VTv5wOy5Aa3k/GfXeYRyKnX/DqnN
+Jh3CYId5My+MljsqP9xe73i2T370eeXfYuvotV5gxC/Q32Izqxkcw02DxZHN0UyXgBByRyJLL6B
GfMIlS+4mb7diRypotjN1VlfSZK3FZEHfdXsJhhwkQZ/RAgaW+07HUxeaA2Ca9lY1iSS+0ptb6AU
JK3ETQIaYlu+29gPxyVnZ0bMe8XrJojiuOltgeuljyW1OKPJwPvAret41C3PatSKGkRAiu3suoT/
IHMBkXJw5kRHhJ6xfkgtCKLe5j06rTQXsE0UeMzbHkdUnsn8E4k7oAqaTER7dPVozzkd9e7w0w64
eecMigCxeR3zccB8pWMBlmVYUgj0+YF2gyP0+cMFheLFx1Hf+MVMZcmcDZe3d9kDXhk/dksXnCfj
Je0bHzHMN0ItGoKl04Q4GvjhcWloztyI2mljijIn5oja3tzAGWyw+HidcigqU179ZKVZPFdYVN87
zUb0XT8nHjMzkb2t+V+WdMcz9yuXLNzmCw5iYpIiHyY6fBa/uy/eFzKZjy4xKVWTMLzEx7LB8j+g
TmHJ9QPqlBbKNFD7AcckgDdcGbIfgJD6hVxtSjpJuaMMuhYjqDKMzN2DtvNoZDBNXMWrxzW09Q5y
+8m8+0I18z8uG04B1eFDHadl0bjODLQo5hSLZ98Ze1wGlNl1gvxXgSqEk1LpGlZmBQtHgukByDMe
4I/q11jIY/V+qbRjxEtqeb3QLX6EotvfOAZ8VmSVHzqTKdpG9aEg+JWQS/BVhS0xJiimhLvIlun5
XRpDFdXgJfN6LVmZ5QZDlLeJ3QzTeiZK2fiaiZ6zpiwPM+zWM0kIicvjoxukGOdY2RJojByXxlaF
m9qgTE4Jqh8lV3LTemtnh0/kifCVSvpnZiGn5eON8fljw7ceOB/Llr6N1izJit9ayFkHbT1Gz9sj
6fwk7fzhH9puhN21XGwaSGVT68/62vzoMWkgWRFrLi3k4mWDr25ZGCgCvZ49goCylclOqw6Jn7se
1rFyWlzfp4g4+uE/3Q2oBAaVJF3TX4VzaqrVJsMALbp7KBep0aE9RIp4XFHPre/12XAL4Dl3uP1Z
iP/zAp+QpFbvOe6ID7HiqnHTPo64zUlmrUaJ/x1zo12gzo6HbsG4lDV+huVP1yMq3Yn3HRRGTFqB
sSW3oR8XuQtczB4wp/YBKRDYd9nyakeuj37JMXXjqktEz3pSB/Q1cy6nLMNHy/yCU4zFLmqXmIq8
pJGcKywn611SHbNs8dlfqjv1Kg1HQr6Ns/H0cR+VkPYpUK01SyXM3GNyLS+S+pZaDPDvk48/fLSR
S7upqvbEVyXCAvu1T3CDHbV/bYKi0J6MgROm9EzjTnCzskfKy+lCODmNundgVRVZqb0wHYrAoE1x
Aar/MwnAoTS+pzQxZc0BYoCUbxpUR9yFxS6WqpCFQOrJwaTc7yefzcE+zyohUFGGKUUZ5SFmM0UW
pj/BwIU61zhy3QxC2SavaH6BLzg8GfboB18UMnm0PyPftE0EEc/9EXWT1snqRrvCN8R048NwBrJR
lfGH0dHsOT36T19yIXEelzRqIj6bpGh28KAPLr2/x+HmHcNYs7MWx7J9d851B2u+nrNxwceTe00b
QgqDk6CYXllVe58o3D8Fd9jP2TvzallOSgZjA36s+5VauvvNzLcGyFAtCh+4bfTEpDmmxPCjejTD
EejCwt0bmq0lxGhq+1iJCVlO4s65EBPCP9YH563NmiWygVomaBHkcI0FcWOcul7dI9o6QAlYYba8
fbDIHL1HWDPeuLTb4V8n9u4MBA4g06OIGrXjamvfTHG7RfxBsAa/Hc9JtopMv+dpT3GrUB9wLyMW
lEzQPK5+4uf6CR+i7xbQFhdVux9tU2qPHtj1Zj31cTSuJBE6BzOeDp0sOyzn0nldKrMPXwDCis9+
nk8I0d34a5R4IRUEaVatePgk5hv7y0etSTzF7GQAH0sjJM1j3oQSwgp7jl9A7dWHtsNdIr0vv5q3
hhUmlSnZkkw+lUR8Ff9WbcXg4ClbPgt5UX6XExxJJilDo7HtzpFYhAJkf9Orlh8UPeNmtQffFjb+
K936Z4c8jdN0bys967FKFdBaQrzKpBFDBXLBH0+XcYUgICwCgrYDAsKW9G1xD3eHB9Nqltravof7
s7cNnXkyDZ0bo/yuz/AEPL1Bmgjt8qjXomSJgAq1PzkMHrMQeMd7kAHjVZkKPGogeSzEKhA/RgFY
FSfiJpP6E3cVW53tV/gKa57qoD5QtVTa2GKdeiB9/A0MbpuTqhf9m0d0EkFjSd51L5WYN8NMV+1J
cKFaBHPWYkqNb+NuoVaHGYOXv+QYbhUVu12wXGGrDzzxQhgMGtoVD/ZBs9TgBx9gxqsX7LG1lYqR
IooHd1sVNRkxAnjbfCJwPrZgsq9dXwFO4yf3qcSeHXkSy+l5QdZfmRV64YZvl1YiMgBIzXzltQEP
pwqVeMke513hxVGfVueAO9lk1NGkG6hnjfW71SHAQMeDoUNGeT4Uw1TV2okAvWU0uadkoIZ+73nO
w/MmAgvRJvjf8LsRXyHdnF1U5lxUry1tP8ikVSlVLnG93bAD/LoBNedDlb1K8/1zwWDzKwn8/S/3
gjrgfmCopYIBO4RlkFH9NvaUsVM5YCIIGLsHkrpMZRjvSPIuo/WMBq+IO71YUbY/s41cN2LzsDhM
ECIdyaehNVZfkY3TGPSneDxpg4LLy2vVz85hNohAoWx3Pv3KuqIpzZ8rk88IEc8ZXObODZ5vtokH
VWSxqFsUJYeZniiCT9aUjJCxCHzn9fsDEVdyrdtzSUR7tGLKkVlSiBXoPfQUqjtJHL4Czoz+kQbn
s+K/GRGNAqFvhgEFfsVuXgl3i/hVgTA+akqJ6qIiVMf7f0v/dSGjiGlqh9r6CCvtDASPTkkMiaiy
HlRCOW0KX87HRCNNMj2o7t7bdjFBgesMZKmlxRIktq8DmD8lX3VtrGBU1G+qZPogwVBxxIELaPOy
tM5ZVD2YMUIrxVvbiqpCk2y40R4Y46yiniXMAjcNA4pHnjg3AJc53EJoah4YjzedUdy8sjzd4ipw
3Lmj0UNvmgpRej7d7n+xcQDQur8kjKJ8CywyPo16in13tp4/zaGg1mxxMYKrFBnmWQXmuy30VHSS
mxX/+7xqSJtor35aW29hsjrR7DlkAbGeI/SbQAC5OEWR9Ym15yl60yUeEidq+uVpx+085TAWIVy9
HF8NOI9gP4+vDs4KYQ73K5atfRKL9bo+OIiSwPLv4lmQk0Q/7T2Pkx/Z91uG1c4EfxVCs/g4sRgd
roEcrwGP1yrHy4w7yq9VLc1AHqG8IBAYmwjZa/nCZbo/gz2vzJw8xXXIjSijFTnTn4pC7P3cgt/Y
94UxOK6v6D8GM+gP7iJI9HKnwH15OSLQ2QE1GfTfNY8/Lw3gEKmfhZCfRc8oUFdFyf9vC27KPWaP
cRXetxQdGXlUZdoc8EnNznTZCsCWM9/O5UNiXmA/8S0/Om/AN5LN2L+a1VElQoDJzavUDmoX/4Ua
QFtjfcFnH4kGQ3VKmTR6iz7qCE5mmE6zoxy1vO2DnN1gVtjmmp3r72Nvwm9WUWqGcteaDq56oI8Y
jfNUkm/RovN5Gy4+pAxUWnMoVY+B18hyo7uV4HpMlJIRwAqn9BhyrFqmp5CMDA1c82QozL3iSrtf
SirRHRBllV93iAB7bwnRACVm/SUTTT8bP/NC17qExlMu0njF57+ofSit2K//a9ht8QbJ3lio8Cfd
EM8KRH/v+dFTK+84Cak+47V+idDEk0jJbiyXuc2dnLcl7ktCtxrCWxedjePGdLLSZncGKPp2yEm5
M3CESr0n/gxXn/Ce1NL1cuUt0hO6by99DoPxOqvL/X6uY79YSoipuMaJnpouT0FVox/IiRWxKiGz
SrPLmBMsA0cKPg96iiVfK06s922gEjIrDzD/yiYXpx/Z/W03xpbuLsdLUZsot34DHTcZP9BNmpAr
Jcjd/c1jKu6XJOtVTCekKS7g34aGLjEksBKx+FGAhCKqBae+cnrD1fozDgq78zoRBytrOoU5e8eD
YYx8zjTGIAhtPXioxYo2hdq778GuZS1i+0+LChKDYHgfXmHTgbCgIlikzcsbe1RaEIUhp6n6gqnN
6Erd/lYVEqeuK/7fcmwF4dxuzQRaz3lw8ezPC8OuU/tm9s4wuVCyIt/FMpZzlOYwQabRUTes266a
HoHX/xkk4U4KcC+lZpwn3YmXsP+UmeUGT3cyb620V4eA2Le6eZ7ySRX6RBfByg8gy55XVa3L3SP/
UR0YbKuFVfv4bdKXl+acqsfA0EEHAQIrc1myYJ98D7HH4z6rK/a4E1KCqDqLFGIu51/e3/OeUlJC
vR1EYdB14x8K0lxNxPxBF6EDQCcd8pZlpFSYK46eHzqcKug/WI6b19B2dIxPIqNK6ig2ruGOzZBS
CRAWLksuyBlHw4q8PHyz0qohjdvsoeNjgIIpCGniuIuLTu0+L+4pXcs1O4UI/7pBU/DGcayhrhPY
X2iNSGslKEAyqFwCwJQ9LhJz0YM4y4/SVU2lrn7rd7yXoc6QEKbsrfTES3DuNAjvh2RM2W0c97A8
4NJgVJOt4MLLhYgLwN0tRTWbBrQc41pinX7pxnSjrKVADQ5Fn/o2GdKa7e5qoMisLGRvZNAFGBq6
EYt1u2JmlEpuplgoH/Ae9dGRO09BjUwFA4IB5TbWRKc1LLNaxa+awpsF9fWfkwycTdzzmhDuChcK
JA02bZ7G6MCklPgAUwwvMvzD8J+ekm01fkK+AM770fSubbK9RzKl2Yls66/KpaZUzFelgpBbyC7k
GfeNdeeE8hD4W+GUVlrwjvbb2CeWhnarXJQ52xvncYTe92q0bBbb7C8YC38YX3gBYE5L1f5YnEkt
ht2Bg8i6AstKjcPeWKLLVPpzOLRwEd7y1KAHSHcKydyfxXvgg8aqZjMXcIV7iOFzRck/1C9dpaVE
pnVqOubAH9Voq4iHm/KOfc2o24R5ZgsEFwoMGF+E96Om6ZPMy0v4dII9BqC2o5X+FOXiuEuhc5A9
vSlP5jsIA5wxB4nYYO1Atnv2IQDJII8Hx/96w0EY7XgBwVFvdZtVzhR2mjGIQC8MtFGiHJBkh597
U2fLaJBfLXHM+oBhGm1Ydxo4Qi1zZk/L/pZ7qM38gP+/PxDeqVaV2OEMD82n2c39wEGIYlDgGb3y
h2ucZ1a/dLW5YFT4aK4koIg3tBo7efvex2AQyKrZbKDUpxUwLWwgAIMoMuq0CSFoFucxuaHADYHG
64b5RzH+q4Q+OCIKoloK6K/Amth4WoTF0JonLDzZPx1z+BTPi+u5kmgLg2b8iLne3PmzoE1LEsbM
eiwn9Ek4/P5Lqd8qPYdODXajyKbIVDAimqi4wABDYpZA5yvsVdXZt80aT5LbQVQfwOKFyYKzXz9C
66gP974SqoOnM1A4lq5pWIA4J7trv0I09sSYCx172LAkqaYSsMNCwSO1837ZY2h2+s9DHdeKQql5
8JT6GLL1KEBVsvaXCx6knX2ll/pFuy1VGX5AJU7F2uBqMWKtApQYzUnsr1TtpbQbec1qFZJyKMJY
GS5ojHBNS+JyqakTsUVX92HNTF3Gmj3KA9pC7WOjGFIcfT86XhEP9w7BU5rEdS9TMQoG/IoeN9/b
TT4MEp0kREoJtB5vD5R7nY0koHSEDmb9BqlCahBc7nHz2ypdlJ5CuEqAF+VeOIvMGv1bg1VGzmox
RDVAgU6+ormtCot5lor2X/JqmynSiGZAKz/SxPP/TQzjkeElxxpSWwylkfAoO7Xs/7D0HQkMA2pU
Sl1wNuDPWtBNefVhL/WUbWlqod9uBtWxk0MADGv58Kf/uJGdSqTDpdwtfHz+48jUrp4mou+sIuMd
nYeYrvAk9b16AMRiHCgADRSgJyKZ0zsrTznha2nMh++JLhcHq4gkNfV9M0q6T4jD/P0dUJWLyeVa
9a5PwqA2No13PPk8y9EdWhJQXI4Aest9so8Yf4/vXg0INnRxH8kSC/fbrDRi1aow21xC3889i9kW
k4y4r7xzuYzNrjL4n3wHk4eDfR1gqMTx3N81bSva96ToM/BP9kUD8HN+F3TWIhDE+XkqDRyvUN5u
+ahuR9df9mhVLq9YGhYsWOlbwQ28sceSdFvbw6SQdTifx0n6pnoh97K9Ep1BWj+zZmnxag+LezpF
yCUc4jgnSD3xcrFBVBTgbe4Fszhv9rgoBfhdhygTiQYoblWKvfgcvt61H00AcZfnYpve/CALfD2m
gy5dquFmbzo+4O/CYmXetweBsA/fYQYJoMILsvmqNkHcfeBfaEXStQvz8GQEpfbjdtr1RkYDeqWT
O2XBxxzvHSzqL7VJO2oHhSFhXvhIAoO/TUcluK/ZcSWRkCeMh+quZ86ZAWthPv4n8W7eR6ePE8LI
EPlOiNYZP19YiXJR+QSbCvMdzksHPDtErD/Ln0YWv5Us3vfzoYgEY7v1RkrujOc34jWuKpDbmQj9
uN/d9cNnglmIp/gYCP4CKyixME+JsoMykY57e0hvxKwhrp9X1C5dDVO3f3A2OoS08zH6553yaQUP
EM0HC78Gz0hbG1sLXWBa/pmREyJGxYLoYR0zKzm0l0yduUiTZvlFFXOfcWAzhRSVA4wW6wTmM1bD
HaXdfEHtXNQ135NNPTRgxP+qNNOAx94B3kZ40BwqrG8vc/W0CaaIQktgaYMDHXmY2Ufx2mQqZ3Eg
kThK82gExvLPHyO8YziyQQc75tDkjaymUAjU1NpRWaNUdOT2uz5xiBNpbOMPkiF2KH1xCSbWFRLp
F5impHy9pOmJNZl+EC5f9Ff3v0hzJMuZtXlH05Oe5ZJMmFXMxtD/6wcWvA2fwewbmX1GrgDy2ouN
LerQ+a8/40dkcSf3J1UTfw9SZ2A+gkqsDTnZSFwlBzmKxrqykcFSq0Iis0YCM9hQH4cYfZ1URfk9
21/nhFBNY9Ev1f5JXsc8q4dSeoV5YpILtTD6S6TwBg+GCStGXytDh6HxAHxX1U0LKYwPRnENb/v2
0SNLEkD7Tm2jmRrOwgct01kBzHGuDVbq1bfLtYZ/URoF2RoF+T7uMhzHFgP6EQu+W0g5XPsWa97T
LgJsg46ZakW9b5PxdLtCGkwt8FcD6tgT1ZW6e4L1ynssN+xaJE7Rhya4WR406cQL/Kmuck+zXIaL
RzeC1pOnvOGrr/PxaokR3ETDXV4ADSUsGO2+bvqGN9gScKEDnzsohTwUbFYDaND4g3uHtLZXmzrW
5SYiCLb3iQ6A1Lul8Da4nAR86mkhNByh3Z32OBq2BLsl2h5QkfnXLhCizJhhsnTMqkNbxn8GiTG1
aL2wsFWd0qIGff7DplV+mMobhBfxPnAsD9k2zoxLQjmUTqealxhXvImTPM863wBXDY990I/1GhMX
MSKLy4GXJnwbaUS7xeGYX3RNCjjHNAuxWllMrbmZUEygDHImSRCIPlCF+DC/UxYeR6tm2PcEfog2
tcFxABI8qMMpwsCwkj0D51BEAJaNlUOzKzm7fIyWNHlWerAVpMySkJMV+n8n0pxqAOHWL9sji8V1
ZTUIwN+cialidQQPfkE3iLzHmAF10wuPas5C1EIxiYSBfkJMFTnxvVLzL4TbEVOgCFn0aWXLVoL1
rDYF8OhG3lwO/6JxPbL7RYB2nmshRqy5T+AftJHax3uIzFglikkXEjW2d87rM5gjL7zymWVns17u
THOtjEYP2n22mMK8LMQ4fMY+fVaDYYt11dpJa3cXgLZdHMyfd4P33I80EkJOT/5/Zf6FKS3C1jIg
mlIWz5alXkjnz9Y6Y7raWSOWXeI3F9X9ES5byXaEDM9woSJ/wQ8PrjG7ANN5bnCtFL9HNgPkmeHA
Q4QFJbMBytL5q/LPyjpl/rjh1koDq74R57kr2HmWC1JVeCoASPe3Y6CRTY7B6SAQJg80iQ5uTixK
312F1jra4hYR4IeRPDE1Vv3ch7IICH78NFy5cs2Ct/DfAmOHRX3NKpC7YiIgKU7pVkXl0L4TG2ip
MoL5cYjz6FQX5ye0LuPiSbKZx1K5Y6/nlFBgr7OCpXecp1SHA8WWwUjLZfeCQAVT1wy3PMfrKywF
GpZYaDuyh0sSyDecwLBFUND84iL9GvDElNWbvFzMWfpkAuTTDGMyGRmlW8WIBSLbrEDsV5GZjN4j
pSI3eKiRrgFFifd7ojLlyp3OeSFpcQj6/eV3EnO42BnC9R9ub2pm7P/upyyL0OUIdfYSmEB845dm
9c9U7lXNhxvoyMp/1KuWUMR6c5eqtW7dXB0QnlhB3k540+fWg0NwKdpfwfPfC9BXG99DIUCsa+kr
3EXgGaXAE0OW6alfaI6tm1rBvkjRHBI4SvkPvw3GmzIzYF7MrGCNxQoIOvVzuVU6gPCxyF7p8D2X
vd09JyizTd2bUJVPaE3LaejDmxYq5gs32DUSdE3Xy5osqVHBRTKR2fBT79Jo98TFtW+9BixABMRW
KeXszJWX8ufyT39fOVX4G3YcGFLR+FA9FYGsI5vA6B4yFNMuSp4iAXxf52weZ7N8FJXIH2ARCRYv
PzSQ5Oh3zFNMkXpeBlGBdkPvuZ8h4e07pKNUGcsAbC1XRv+6p7Nsy8zTH7A198OD4BJQkPh0oAwv
p+oPW6TjcDWIElLqFLyYUp66L8A1kyPI/PiDxTWPfllVgWRPRm8UPgScVnNJfJ1iN39q2vT+giuF
Jv4DJLInUd7tbE/Nura4MMSKVPeYffpprAf33uvb+AqLXsmsGeNDJOWohj9qCdWodxxP7hS+kJ86
pDwbVibrwt6VGxMCg/MDjkyci9fLYl/xTVPl5pYSW+3/FvMNEfHHDTZTvgYurgj7NYgHWx+d8j6A
ddbUXaRspkIORO21/dOBSkDi1yoS8Y+wJes6ZVeeuPZNLW06mY0lNZrvdihawlWpQjhsEu7HfveT
nHAtRycNK8wSAfYyaM7vG+FmyQ0AnED3SnIMCmjkNyxvx9iHq+ybVup//k0zLeFYiWfpqlQQyJXE
8kLamV5jMhsGLHuWckox1kvpArajL/5vm79ZCmv7MXxshu6py+413CM1GsGRnjCLddRhj1iiNgmb
UjfHFECw6HiSHXgbWh9Akv5KOcwKAYh6D9uAdkWk+cE+3T/ZrScZEaXfRGl+eXgnh2l7QmKrRTr4
iv09eJl9MSuOtinykkEGtIsTUZpEzogaDD69BRQxQmO9KGhKuhGY2SbK59PP9khUYrOG1T93uG66
77m+5+IXI+SEv3SgPkQjA/nDJRC7GbPVND/ib6ZhhW4POCL0ekiiMfaUI5Blju4Dl0cwQsMcUZXB
1xHiPhxwUGoLxF00VL+VNad9CJ9rrvveZXzhrSAi13Zw8JKIkFdqA0o981nEgqjVAsK6Ms7ZsNBi
tPklmdqlmIYfdY7EM7N7g8VWXJG9AyAFk7WlgNwvF0vojldX0wxK2FJvaGSdnjdOdEHIqs4VCNE5
QwCtk/bFEGA62fdYrVupJIRUEtcqZ8Xz3CzNTWtqYjxRmqxB3cKCCVn+uCj7wlU4moYmQ0w2WlDx
mN1w+nv8G0NIAqKTI8sW8WePNyYYe1bVsQOGhLxqDALkSpBLrQxwO8yCi1A88Eb7bbxGdmbkJ4C9
L58VVmzSCCIs83eFN0yJwnW/dSXjtqXQhtlyJKea6GHoa51/tRSqw4r1aFGdOqiv7VWzWRv2xR69
Bmhrg8g/ExjO5b2IqfIbX+KFbri76XfUgopndx4d65/fOKMmf22O8vQNEwuuGgaLak6lpFYlWUsX
iTNlAtDFe8slmNtI/s7wUOWkpotI6KGBrYAcTXCi/jnS586AV9xgGdBgNLEz73xPIybNs8Rf+GNw
yE2M8NrLjWkPWLBfLHVX8xrKH3t9scr4EcQ+Pt/pIgdzBXtmpavybvBkHebkVzfp9WHw78Ac4DLd
vQL5Rfc4zU/EtNxeIV7MhgVuniS0kutUm2kNNHLit1l1ls6osPp8BHGdzVIla/ECYYYta3H6SHf/
XS/Q5RNoBkTIu4DxJYQLO8VVyKX9BD25IjsfIL+uhI4B2G7Ip9lFj1PNkvw8eXr5H3fNLMnvyVdZ
zPl8C7778ZefdOp6ICZIsrRQMHNkbOWOnW/jHATdTxKzOBCEsWe+XgutWjAJetbjWOJdpZqpxyyJ
mKJkQrQEOzkDSOTWbsQqyvlvYV+UzIEOkYtSBOWMJMBGydZz+U5m7doAYKYdhBPJyBfCS2jAxYfw
4Obl/TRiHNax1dD86jDSa0XwULX5SYdALsYPqlnHY9sDwPBRXucUyPManYaha7NLdvBBBHfiIErr
UQxRu22TE5PmEc5+PWV5XblcWQZup73r4mDHaDxEB0Kv1+3kled1VCPNL/lCU23JrJUNaKGFRKES
fiuJr9wV3hgmliB0aJjgQs4A7kbvx1LXk85nZ4wCd5MU7TFzyxRsW/N9fWSY+/yuMhieqvD9jeBg
RW++nMPAPQB97xLm0QdvMwcWlGBKnEWKo82YcQvBDO23yeWS40VckQsQeq7TZVYqnkV+lM4XdeA/
iHVmbAlRURZtXMPyeR70eaJX4qgL/HUwDpUu3O7BuFdikHSaofIuxn0L6jgULUtWGSRkNC9MEAlD
7Ghqu3sflshKvEFIpVQKEHZbdbk+JSMgGGi/pVRufB/gzVMwp2/DUBk8DGBOmw9ldeRtjVMsmTB3
IHgwbp5jIMrAwbiGxnxtsIWxAleLJ9FYBv5I7o3CpCXM8sIfsa2HolWerDnWcEcZV4q1HECCqHQ9
EE5ieEqNZxgBxd+EMWhc6bNbGCwaGdeBcFBOJ9EpJn1YD0+14n0LPOD5Mnam/5REYolSmHJKTGa2
4NVzrmWek22wIIv6LJPnANxenmuv76wqW3ddvdQfUO+UygpbP03nvSXgi+FMrSgKaNhcTcnBUn/M
xUMmKg2s3OEf22QlhmJkws2z4PXE0oP2bIwtVOd7lEGNElEwkVxrX+SiWINMPHiu98/rvHfWvLJc
duH5A1zSfYsAc5xj9tGQMKJ2UCUDMI6xXbPLlOuk37/s/7Xeb11zArV5gUVl4RcGjx2iEPnwRwKV
ulMEJ/DK91FpsvuKbV8tFKgDuP0CazmBoCPS+RuSvAA5QZvG7MA7e6DceqdqYJ1XNy6E1eL67URG
M9rVOkcB//gPCH2zdVXHYzaZrdtY9JRY+r1vJDfXgjSuxLuQKjBoS+YJN/Lm5KlR6ChGFA1mxGZD
sZocWi3uACClY5EyPjyBnRKxp1kIcjrKbYxL1skBp3uR1PZucJ3RnSTjj40M6pm6BId3z25zp3/t
KmMaGqe1teI1GoVqUmKworItICB9CYruEhWnnkdpl7Zd2ZxzdO/TNwOCbzIMkzYsO4gc7GeqT2GK
Pn59SepUhBvIrjMSbWsAIAs+LRzg2wCpJUSVmUQ8V4LrCdv9qYygwg8cT6l/kZyRYtOQQYKPvg8c
NetVsRmVux74JxWuxZ3duI+Zh5FWocbthRvueVDkQC/WjtjmfIMCrnTMjXKnCNeL6ABY9WHFGYlM
LH3B4updmitN5Gg7ao9jykvfpayQjEvvFjWFUMFfPP8uxfxz7kJjl0jl3XnDiHidBV1kIF3VFVIl
JvGbLtjINZU1IF0xQpiRqE+7LAVYYDhj5SBReNegbEhBjVb6C7brLfCLB6Cd8EsrqVCnxoIz8VKL
VIfZz7RUDo8P2HNaFwPuSkDxdo7QaFjhi36tLQ0DM6uiubeGmP9gHpJttN0vPsM7dvvbX3LkYIH9
u90DODwnCM4lNbJzBDK/Nag+ghEFaexFJGyxTf94pRCZirq4x2kAQtALFQpT4rEJTZmjJKAT530O
xLYNfbV9azu/eRnW5s1lBIbkSE7W81giZli4asvrrS3KKrUAcJ2bT4rlKKO0pyTu9H1p3xXMlFtb
L+IZTPITzYlg+TRue7F1UDUWMX5P3NwgNoRCgUdgQxKVO+SyrmZVEP3Gxr1SkdCfsNKNvNg8owQ7
Y0gYYHc15OsfsRPXInZKCtk5OHX9zFsaz9ZQ1/V/oMiCibn3dYuX2dmU/SE74extvzb7OlyVA7AY
YrxPY9qFePRPxYDg446f4Yrj87P5ZeuxwQcs5SBOCRqeYl93MvfzRkC4wmVkx5gpSrBd3MHtN0S5
cEUPGaUIW3+w153x/1nFpjSZXubo0gwPAyyRo3xq4u1qF+Rp4k6SAW3HYtgh6NMTZLMwcrXGwwef
SDia/sLGgzlQqO6IwUVnQlJ3mYJTTavXYQnti7I1Dab2EHmQ6C0UjE5LlS/8jMSePGXg2N+yvgHv
RhvS4PXvObn8J7OlcBZXw3YBwNy5+9AoS23u/LehZ0jISoK2/9GqJPoLIkOTXBstbPxqqZWmKSJj
A/DbiHDVx7pOVqQAw4vij83jRjr1zmNgJ2bGurgH/jHjPNA1QLG5ey0bSA1lE2LsIUK04vJUSFs+
/s9zUHDLbzL48STua+JbTES5uvayv+mdrHvgm7xWvY2IrT8eKk/OiIBQJ9xMJw3pv3i9uG//CeWz
gSU8MA+mJVAtZM5wERMFaD3x++Yqc9Id2UTi4ZyQb0Cq4X2KgWUV+dyHTRYbxEZGNSyvozArQSMu
ZBiUz6Mmb88tZrqFdXGpcgiayZBHkM9ndbtsvIR39yl0xLGPObPHH4IGfRkBBIfCLY23XSSVynXa
62uFc7b+bitr37hG3nXlte19/uNn1TYUcb2t9uMmM+gF6tETNxZifD7ATcy8lhewVolc8b77swhQ
AKoYIszuvtT/WROwOzpLXrlvfQaQvai2dHLhGDIv76mk4hYNSVtS6pYWPWJt5WQF32vjR1lwJhAd
rFJFPmSBplS82m+Eh9bM04UnLVmmreNo8BEVibVA60k2nkVbcsjIYMr/6tznNn9zJWNbN1J+8jVl
/E4KnpngzaW5GQkUcrdglVaP/bOZMlmUS0Sawkr490SwZvY5c2MvxHWvfeJ2qhzt94lS01zMEGAR
pk3bDxiyi/aYigJkl2AsMh1hhwSaNjYGfkC3+APpsLWcTsjC+yf0GyhC6347ElIkcKMhJm/TGNl/
s+N0cHDT8d3Aq1o68I5Pn/yeUZW5twhJMlNkrnMplTIsuwfom9DA1LdCI96Z4H9yOY2tbRNNdmzD
fCzdt1QPq2lIW+6eTJLt9vQZirNiDX//tQEAz5jwJB2VEA4hyAm+dzJTzg9dOOv9mcDF545HLGFa
/wXm7Ij9SSKOg/bg/5zuOJJQIlNolQs332n+j2NpIx3I7tpaKtzrOR+K1Okj9ZpnRC71mZ+xrXvy
ZqjPbW7suk+GuIYm0VhhlBwCjUOFlx+lv+Bwa+bKYDD79eoLPZ1GyKXPSElBvI+aDKqnoeD1baWQ
CiDX9AXbMhdPKskVzdmnOQ7sFn1X+rn//CrJwwpkGq1WwSaxkLJ8bdCz6yJP0E4Sys+TTxXKp7fK
hO3gqvUtiOs1//5fI8QJVwSAXScvh+79cYeNKw4Qi19H/zblV/nu3g77+dD6dlM2jqKEO5NhHDpU
9zP4GF7KL85NimzP4YdOLWLeFnAaN+JaMABKifi2nQM/MLu/TnkPS+fbyqZIxMkeC3u+C0IWsUvL
lkQuIbxx6b/1t+xkTq/MpQ5QSRbOdL05B3wVdr33MVGdMgp0wEMOdKzxSwX1XmsE+3JzahTCBBD3
TqUZshB89vmiFOt7XdfXNNkUJny+JKyDdOhUcI5Xg4MUnGoE7OlxczwtGlePLxDd2JeGQSK8oKXO
G+G/D9e/OwmCVp5PICcyk4resEnPqbOnpbfPBb4YMfrlnnYGdnzTpOAI1Cm/jJXjDjQOajd3UgN5
uTvVKxkyZfp1oj1lqwHJ/ZVHMmOHqzZDyG23mKTAcLQMedkMmjHtOpVlvp7+FXWTMiIuE0V1Eyjo
zRmS+mZa11Lw1ONnseK7jCJGdLdjOR/vhFoBsYw1gtEPzCo3WCpDemak07zcNIAs5k7zpOAfuAkd
0WCD/x9RXv1m50oTzU+JvSJk/eNjXE8ZGtqNmoLX8TmzS68hFAiYpWZ7M7XOcxLljxWA4S2a3lTw
TgHG17oJiV38pudrJ++HhhusKkTl/esVddZ9LoQ6h66WD45BZa758XUe3E84zqaCycR+vvNXSirC
mBSq9Q58XL29NDljjw9cGwsofYnrgBX+GPR2VqWYEgyblJ5r9urks27kxkpS+VJrkv/TJXGlaXSQ
rjqduEF9x2kwI2DebmKp/DRXcWbM/We4upiDCnZnszskp9nv2nsYMXAmPMhrlZ+4XFfj9FYjBuWU
ljZzxOXe5g23FZDM32qO28eLw/riI0/YxdJAOoC2Hpjnt5KOfB7QnPhNb298y6q9aqrDRazHrQWn
7Ti7kYDhxGG0ZEOJFNbUFMXSTgeHoSar+KjBxRrvQH3RQW+uIJYSLt6cyALRz11+kJS3mSNRf54e
T6GTDw57WonMHXdMtNr3Z4syXYjf2r7orWalIcT+OjWXtCvs7/8OIM5Yp12dgcDpH0Ew6JW3g8XD
BHFRqyLNWSGBMUaSLFwRutpb/8R5mKm0VZjU1BjfTSvdDaiA9rcKIhkX75RtIc6lsNqwVRBOYMg0
RLGK1e/ipyTEifwf1MPnYRfd2BWtKMjt43f9n5sfQW4mkiwBIUrxOCAzKO6c1ZWTZTiYLUs06ojZ
UMkjTRIP3wt3flaFQFqCM8FVfJnqBmVSrA6FWmy/46DS9xeMbVqwrysBcDPVua5a4QXj/bBMdhCD
AV86jR6nKIIVnHLZFTnJL2OR8xTTBvHa4D8kYbQBd2OU+MPmSXYB/b9QdyfZjHpvHsTE8zZ5ooz/
6DKCFO+z9fp1gDyMd1Q3taW2oDzDZMw47w1k+19seZ/SKmfoa2bcOGkigaSmg664NaIwPRXBjf85
wnZXjUM5Kq9IPO1a08SMx7IGJF4N7evBy/ddQonl5bxmtSpcaL0MwNZNPYQyubWCpmJ4khkKRT8q
OpdQzf1GnHUVRqHHoOUc+vsDLTJd3TFv4bNjQTBMLAF0RkB+lPy4j65wxMMLqvMTxHpTDxxsh2/L
fOXTeFKWhX/gnB1O/XEavUNb4DkKek94h+QGiuQFSm9g70zBLZJ3ni+iwrYjvhY1EX7pA3MsFJwk
LvtifBIaTwKkU2rwSnLjpU18hNmsZXxLZHX8UMTe1SeV2+kHDZo8kn7OMBiYZwwTlUxy8B0Hu1JV
rs0WLpNct8tBpPZNcvHE2OB8W2EKZAs4FIPNekXGXQixMlEHGvtgW79PdFYzv9EXGvY/O5T0MsjG
Hev1Yq2r9Tt0ij+eEHHRrjrwvJpijtURC5DCBkHTEqIhAhMRagxeoyul20gxPJlKPZRwinpaB9Mv
vEl/3SlDy2reR8FYZVFiKLfj6GleVHPR5pqpzMOhi8AJXT9lipTJ4f4QhU/4gu9Y37jXrMHYblwz
dw+nq8zN/i/TvDTcHfjTYRNXPYh8Z3CvrWd41zt9Hfhiir6luN85qYQ2FVBoTssHwsUHL6xYNOgY
pZv84uNKv4LrPMPUCvkEFp4DG8EoXhK6TpgnlDT+C7bMvR8f63sou8A45qwatHq+CTuuq7KswzDs
PKTb+NfwBhqa43M1SOiRkRX8DmEGYoU6T0QegEQIDtGTGo1gQwbjexnDFSHFKuv4lTrEvSYBYn27
sLGH9iEassOQvNnpqM5uQ0aXLBIdcZyD4QlTDN3gFup2lHKxLzaBQlvnWQPa+8TemoEWx74YsRKp
F5RB/6IFnNgR+QFB0J4DkkzO92xd/oZ2MS4vh1QAed/CvEV3I0whSFXUrRdgRDcav3bWNwSdiyGc
iZTaqgtELIZMYnMqg5o8B8KnfPNSA3S0uh+yhbSyRG/5owXY9gi2tODdmrwMvOJ7nA5Z1Dt19gZQ
Xwvu4HRbp41KedCELZrPDuv36VsxzwWPEULyT45RvLR7T510amoqqOaXpZDHg7k2yH5cbVGIYME0
LfQLKSkdThW6jAOD1BQQAa3v32JckSPuKKHQR0z4danKxL8BnYld82+srXCBlishgIAViebddZl3
LX1IDd/bw6UcTJoNZSM61SjcnPmhZzXGMUEvgc3HlLiJDNCnCwuQ5OySUWMKVvHo+VSA71TV39ba
NErXdNLKMQIQuSszfbdA6alTXZLic7rx3G/GjZN1fYiUR0FPyQ1Q5cmL1/P+1pTEkahki6AJHCyd
OLn21qAZToYdQZJUfYJZBmv2SmYjnPeEfzuUkKpDGriaaRpMV3Uv2w/j8mu2pvvWqM5w75h+TTJt
i2qRxcumnLF4FyaF+cIRBlc2DjuX+bfol8zx7otSG9E/VbHTiNbNSpcZuEB6cxp8w6eP0VjWTRuj
whOGiHY57Yq2juP3Z3r0xkQRoJCGZiWO6wKIeSO9eH2uXnNwfjUFtuC7FvwWnjQf/zdRg3a+ACsD
YkrO0V50UTNNL3vTbvoXL0hLAFOjNRKD+dIb5UyxQ9ilzZDlXm3hIJyCPYFEqQeNQghqT1z2k0wK
X9+PEHaZEordYFm34E3LMMOC1+fCPu9jjc/vuQPSv5W3MQq4CS1TdX/feRVjVNETaF/zN9nC2UO/
9IyrBm/YHWgN1VvoJ0zrF4ys1TVr4JHtt+B21Vjb39RhUhbl3aJBE24Pifs1MojmS3DnbtFmH/3X
0VPM+Xcwz9U4fA8oRxirj9sjI+U01Sw4iPQUc839nvi38nv3SQlTFC5x45+4yVj6IgwzcSUtzQTQ
xCXshsSv+8FkJxOBTEtqyzR45G52bJhX/rIueE1ZI9LG6VOlzLwgth8Su3Q9RQL0HQnST033v5Ai
u68fGPKE0haBWnJBDlmiadCEh35S6o2CJidLawSpxMZkj/kmJ/zOS5eBX+e7ACXGp0DPVGiIWKQG
0Gm5gaXL3MCqLf+zE3rlGeJdC+rdQIYwnF8mmXM5/tFh1eAZcLmcNMthrHqtKgq20/fxwSsR/3Se
SYPNoki3OsE/Ho+nKj0IxsmibxuYAihjfoxLzkU91Aiyq6lQ+Bm1UxEhJpNPnLs137NSrS65wIso
bhjFO1z3sMmIYsiuzFXLohxgTFNrYDrk6fM6vIq5Z3a0RRkdyU5/ovNEEuWD5U9ZGwotzmCpEeLp
jsCqaEDATmZKlDY3xEvjL+obrx7bg6FwOy7crs671jiZQXfGNsvCUFwBBXpja1x5RxSbu1uL92Vr
LS1eL7xWBqAh99f+bxsI9UDb2tH22Or92tE+9Rfw8eN/z+1wJpHP7T3eVSFqleJrY7WEV6iHFrKF
KP6MxaIHvn3gEVoOqN2Cq/xviaDxaW+JWFKxeqE/JLpGfznE4emgsSlP9xCAeSzBlkqBm1fRK8iX
CcqGXHTfs47U1Qt4oxMs00CgNkBI02ySoBFuGArN9Ks/7WP9KhiXWaLlxb14tnALpH8OgaJmvCch
KiiDtuq9/0ZlxapIpsNTM/dw8XUVTgrDxcL7vAz6iRANROQ7+tDGjlpBbiK/jzE2wTtS1VZbUMZR
dFmGFnhzzVXlozHI/jT3RGtS7PksWAkkkuF/fXSZFYVathcjaTadRq+x7DZURalKdPUg8oXlp/sj
LrEvKPFdTz5pIU8e5wyUeXM7h8NnIqXHEjgeXiyLqu2oMBSJ0C3NBhEMEranu0zYgwlLNR1roJzr
6Wg0FLkNeemT/AIdiDcECG7Jn+FMhw/3NbERSKyhhqri0diYdl5OGF1sFYOJgz4EM7IRO9LzUR43
655MmwAob0Nj8Agc4KL+dLhE/rJuwqCWsuoCc6tZkCQTNqoDtHaPmdFtlMaYRDUnU4zzCobc23f/
mT7GYx5SbGY5+oi8d2QeUiQzSxSAJ2QMSOgGiqPzQDUUQezmKppOkdZ5swKN640d6k6RaPCXl+GR
ZIXUBy0VgJmhxgMljsBJkqLmekvnL7hebLfIgoE27XCDMAluieLgD25UOHX/KbfMHH68t5vytczX
lSpMM2syL4/zP+EDq3lUMQn1JkBNFYe6VX8J+/ndBymKl2rmly3A/T/Ua5E2rKwQpzJQJFuZ4xqn
JD+CsV+vcrrIuJMx6J2o3ZCxIeYp9afb5BCKs9K/wjgjL2fDETnWHbO96brt4f99RxzyIqwUv7/V
IxMYSlK2qlRjRgEMlMc+lsw0qSKDKA0COk8clfryRvrzMKQr9BHNbnLq/zrQRGQiOySZmaKGcCr5
BVWAtqWsMPKVZKzs3+RU/0G0XlrmrdefSuzQm9mg4fstxNSZR39WZBPEAEF8hcv9BoZ9ptO1ON5+
hkhVW7FjJ8cZnmlkk1YiTYWF6Tzl7/uwBSyH1IkBsUFIVv7QrXJ5ofBMzZmp2oE8N+ztrGQsxZjQ
5JVoWefKb2zJ0uAns84wx7djogcHEOk2SKY64xNNK6DPW9Kc68NkicGihg6o3pb5oehNPxoJ2aNm
mFqYCB7vfBrwO/Vc0SwKFOcduKgvk4qgaJdTm6AejTrftN42vc8jxiD6NF1pPjcp86B5KKrW5Sa4
+9tg/V4qsN4LNa7dirQgvAY12QFI+5SjVcZLL7rPLw18nKHbnz2TrGz929P01DB24Py66PM6oBhE
ey/FwS6V/xXqFYyfBUeud8+zokxGQ/wvurfdb+kB4/svrJT8C0Yf8rZwkPrULMKk5CesW+1qYheL
N3kCOm0R8Bg4vnlX2BpqrE5ZMHbMXldg1uYk9D/QsWW2hkM+W3FVq5d2uBLKizh0scsSIkHTcrNI
eN09PHzX32k+wmOMRNDprjRCoWcFwufkNj3grM8a2wrSJfekwbGYIIL/J2fh1pMUzXJO55xkqbXO
vgdeGLwmdTuKYQTqev10DkGxaNx7ic4J7sP8XYcsXJtCW+YeFBYRFEki5f8GiJ3oKu5pE8xWLKEB
ZKxe3W+BsNlMfQK/YYlDsTrBP7aGRM6z+rWMlPRfJJj0x6otGVlQFGa2ALm/iDpSGWNzTCne0ozL
NhEYXzCBGozz5PUPWXXtWHgWEbjFYDhn6uPzH0haf7ycXUTKWOSG8mz1GZ8NcinWAqDBA7sZhRip
Cx62Kxy6QS2rhOI0mi7HaM51oS969uefU9U49+Te3gIlh3pvUHd/h6Hh6fvKjNcx+tWRUGlPJXFn
5ltF3h+l0UYQdq3Y7P9fDxzhmGAbT0zVVmEVONAqRCYspSE0W4wX8UEhaAVlExhWuPU5byW82Mmm
Sq+cW7XlgNS+O7P4uTVwJLaq6OQWV0NV2QuvkAj2hGbOXpds7bR5u25chC50h+OyNFRS7PmPeWzE
Js0pMUS7kecREWRigI7Xis22tt6CkT8jgKjQxsHLjxnRanRhFSO4OlxHwxmVLGeEQ/WaNXXJ7bbi
uohVeQ0SWfL5ERSOOjRm5x/G6QnSNC6w0kgXvRoiZVJyIGwN3TBriBW8ZS/icoMAIcWFA7E0WF5I
Mama5bsRAgJeL6ZwR9Fgt+YLwhOAn4ecPb3rBeXARMzqktioYhE9K088WyhX092HiVsNY5VW08Rt
raF3UXSlI8fCt/RZNSLefDtr0cmLu4Q+ssN375uZ52e5MwrOnogM+OWPwlMtQsUAssGkEIXxwHQo
fuNayJb6Gu9YRRpKDt0FRZnqAJMG0bC94PHiYCTzxV+P8Ift8G4meJ0tDh/6nR4ER7AlIy8xWFYt
9kpPDQhBhbohiuooHfsMSAfBOmwKB++rLxsN4CX21nzt0Sx8BKLnVD6NfNYO5vuynjcNGvXXVCox
ZgeNg1ylsfeA1U/zFFu7tWqND99KO0Yk1DCMlwd2EKRfv4KAqda65EWHTybaep52o5DceFjaw5BE
iRvtOvknzp4pQ+wLtjyFUbi91RA/20SJds+eYIwUZzZjcNoWvz6V8bldB/rYm6OSJrOVh88Wp+m3
lb+DPD3MlB3R2uiP7OeynNRqL6PyrOTkAZj7I9WF9/nMeUvKWvjbIDfU3R/VfhTfP6X895mn2glS
WEZxXIc/BnMImz7CmqSMsFB/pwcOUDfBYw3jxeRuC/NrEu1TTDiuYICrKcFxKOU6miYC5/jx01Pw
OXSXX6fIRSi5+RDbPko0ce+Us4HXLZ/qVl5pJly8KRKuErqbhcV/fOwzFO4JwtuKhmjW/GHvd3eu
gx2V4tfMk06IhQwDUHv7B+nkB92IURFgVpVr5DRDYl1QZIJG4KNsR+XK4hYT6gppcCx25HgOIlwG
7tJpnJ3K4cnSCmMoeDJYKhEEe6cxpA/ZWm7BxJofAvxwiv6+w2IX+DnU4bhc/DEj3SFCYwAZs8m5
rpvt4FTwz2yZQThJqvePuvbG6EAePQUuTbp27Q3QVBwOr9NW3yG3tNlM4TmAqBCcEsIlh0cx2BlP
0MTq6YQqP18KFA5W2zw10aaJKywaYtvIXccczC/TEhk9YI8/hQA2kI32xcREyLd3SL/YiiLySSxI
ynA3H5V2L/e7wphsOVddKFVCizZWsCe0dKpX39XQDbAzucbWk1o4i7oRKDlJDSEAT0wOjIAQoK7z
Iqq9+gdftirAie6RzKPKO+yyPzSNBPAGv8MVp0LxVN2T2km/lYucJvzNiEFirCaYq+Fd5wPPI7vT
bTopW3rp/zG0Ui6r3Gj+KnvPpYDw1UW64ARws+TD/zpc54EHvItIZGA2mvQs2jmjNV7YreZCwjBN
buOKkmOLi+7p3OO8/1CoF4LSfM9sZeqJ+TVHPgPnfs1Ig+o8e28kcpCBdffCzhCO3E4kvhL0xPkr
jQQxdVIC1/t36Q/4r8R+dgbyWbET7wm+KSHCxBXMSWf77UxqI3HX6Y8Z+hdOFVThz7drkT1QgS+Z
yjHblXGhOtxL88AZm86qCS1sZgnof4Pf7KFl55SKSbtZXAvOpb5Fxp9CnRA6KED9cGqbYaAUJEdM
oiOC+slKZWgqmsTygii4iVvFK5Mur8Yrq1Sf1Lb7yD7SjoAMw/+IyXjxGqcysbAERD3sPJGhY7cA
NVnrcZ1hjKZbcTeVI6gnzV19sto+i0jhiH1xX1mLsWFaBdBLhlyd8jzePCnDcD4fCO0blkDbwaDH
5apGg2YjbzKjRUF5Dddel6lXqOAqblA/fyPCXnvDwB+jj5nWMzzFpu3jz2AisAsaE4UqKJ9jl4mc
dnO3sVf5eXHK4/4GFJxytYgjqWKjjX/wMJEHtfIj8iSMEcsDl0pHVziA8qDeAHon6+/d5BZr5oRw
+U9Bz3u3d8d2BrklF3Rkq1o4N2Avu+/A8Jb+6WN+jwwHzBVtldnBcb40JzEMT58sPUSGJE8kTapf
Ac/XMU6LPbiT+t4x0yV6RnvUNPdv7XoSAQfw5nlHRLV4OTpWg3wflGl5q+RKxrAeVjypaRN9kysl
bE3kkOniLFmnqwTNn17O/usNjpNc60fMnuqxLfbm+a8dLjUrVYZNQB5A4ju++QgxZdGbmDHAfIgV
bCBCPrFJNWUWlUEK4EdYzHy3dEagOZI2mL+B2kg0d6Tz+xeVBGUueaWrLGGFe5AXDpWGXQGTtams
o3ks/M4XryDclQbR4uDZu+aTp2YIS8AWtDBqhb3lbL61513fmVWDUkn1zJ+HvkDTC+fSjtBB9uIE
NyUl3gUhTz4ZA5AV3IiCpGVxfh+8S/Q/mQnOetSnndfFAoVpQUcp2MrG/B6HIT32j0gEfOgQxDUg
AtJMPH7PTS5CLBJDRkH21OL1OJn6p2Ydry2+4Mwh18t1PMJ9uyy4mUtvfedyyGiqLOxfdklsHlS/
hyR7q29+wIhGue8UBSzFjNnZ1BVIxVaFomrGaLS10grg82uuqrkY2oxxQvvjPe63XmaVrbbqvVKA
y/IJfQrGYymQfU0vPZyDbby31HwZflsnCo2it5TDJYVlyZrpewgkT/ngFwVGcprGI/tWLoaX7Zvn
uOarDdIzc2o++t4Rqg3XQUuPn02/VUc0V8DJDThVxd7Eng9D1IO7G+AyG1n3yUm2W4lznyBdFWg0
FfVytvJ2v50hI+VdMPXLjfzzc/83F1ZPJUlCaCVTBsfYLsvwy1D+ZZ7cNqyWUJWocSXbS+caqEaq
iMeko1QH2CkaB5WKhYgDA2MmA2XiDkQ+IuiaBUQr0gazQ1Xkdk1zKu69MlifPBPP6NzWr/N2I+zi
M3d7+wHTMbu7Gi4RnkhnZHqaxe0mUrOLkN1qQkbfPgJD/RuT0g2zBO4N33WOmZnSjlEDt9qL8kqS
AJIeQ6EKJCvoPFhgkiNd/98NM7n7Q1f/wrfz0XQZSrXmVlMGEpHlwNjznLykFvupBY6GFShua2Tn
WhGzBkJ/473+OxdASIFjop5abGvocsnSorNOV+A5t4h/14A/5UgiBZ5DnBapx4bnSTh1OCn6VQPH
2x/8JHO504OaYPL2JzZBJW8SqcvEFQt1oed2YFQBqWxsZr6dud8+S1wstNBEmHaejZarECMMdP9V
wJzcroAf9/OpxT7YqjeSNWk0oxMhFihJxkNZtrJFxdvR29j51fWvBLGDlLdbw19xBaQ7KEriJ201
rO4V8Inbbe/OhfsoTCq+Z51JZGyrszshjGpHT3qKZr+gUlQIgQSzBWWrPlO9X7vzEhQrUpz8MSZh
gBRDIVddP8DBIr8ulE+EGYhkhOmOr7uefpOwM4ar0E/It4uLllp7X2SWO3Pjqff+CzOk+PZ1IPKk
gUe6eyaedio4z/AentSkG20ZI/alg/xey4WRw2I5F9qvV6ZfwgeWytfb3cqjkANpCobUclnq64rR
u4FQgW0xiiM44zk7yPV9tJzbTjzIHs9M5ZcyVy+8k5NRAKGc+dnwUhlx/JAJ0IEIC7bsJN4/vrbu
0KRUR28v1TVExfQN57SOuwDH8tJyya1qEaf0I2c49iLv71ofiUSORcwksL2zFz6ctX9CXu3OlWoP
DR8FmKPnLq2C8QKxaT+RUxBw5lCUaX+tjLSfMkqYrs4+/3GjJOuUeL705t0dGpTC3lV2e6JNV9Ie
PQ63R/XNxLZKsHAHWDAsqhmt0qGwoHAA3oovq+pR6t2dI3/rD5jGBsebVA4+3iqPSGvkJWKPvr5W
bray6mWGsaxd4rApRQapQ67An4erwkLWsOXMfdt4ZPwubfU9dkhw/287oL1UXWMo4v7d4px0ytD2
DNy9lJTuCD8+LGhXx0zwIWWnB/gvrVzQRQUk+TFEe0MSvRbh/SozwwgYv1LJ3TZbzAVFwnNNwkP0
FBLCKMlRCnl0IKkveGz8cRAIYpTkBy45ktKIKKe4/LB7LKEwLZYOz46w+C2v8ggOvXNS7iJkqvAW
wk33yz2J5cTW9hZzyW+vRrMZ2E2bzOIFS0qZ4OyCK4V2ya+heQf+R1ljv11Z4tfLQJTIXcC08sUM
BgV0TxTWVP0Jucsv+/itBWglr6OOvkcsmyHa3hcgsYdaqOR1dj5NhrPz/RuNDXrrXY4TsStT1F27
0v97WpWq04QyErJQgrAJv0f3sna8x4EcbMoTVYyaiQcJXoXfbTolLY9BJYEwWDgbq6sheSkl0owM
dR5KJr37v/Ef+NDRTE59ERfg4QwJwyax1BVJVOkyMDZviFb4oXi3piY9pq+6DvK27ZjVhK0p01ru
g6pQ03NfkwoDbm/Izyo/BdGofnC5jbLNgEqg2lGRUUHFBRH79Bk7vVPvoEZ5dXhiGaW06bhlbgDy
ETu9OfrkuD1U30OpgtzZtG5IvNIKO8FwUPhtnW05bMgg1D7al0BaZfj4INjJpsNFuked282eRxzs
PZ4nbV7wEJ2xHJneG3nBf8SHE+4urrEeTALCRsMgPrihhHAQSTCsooLqImNM
`protect end_protected
