-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
eYTytPTdOxAsPKhx7vmma7NO69AJc824UtMW9rpjzP32l7sAortYwgLP0pWLzIu0
qFmfqIiIjyjOKufE0WWC3swuGeAd8QuWDObxheko2QcCezj4JaMDdO2ENrwhhrqf
njXo3GcU2LQF/JIQQbdx/RiAFC8T1tTcvHZKtHF+U6uV3vMnWL5egA==
--pragma protect end_key_block
--pragma protect digest_block
NfWadBHLJJPi0rCSwUsn8zV/5Cw=
--pragma protect end_digest_block
--pragma protect data_block
kc87f+D5B5Bsr91Ql5ELHrB0wYF38g8p9Cbvvb0jZBQ9azhXHgRK2MGGsD3gjf+h
6cShdO+ApPawckS6zobenRnqSaLagyPf4DF7suMUsgeaWOgEehPM1MRss/rEqgw0
+G4b35FD2wY6Yh9faBKpuE2POffqspIlc5aUqfJNyZV8yrw4mg9quAfQ2JMHYb8E
lBWU6KDLNeSztYmkqrBx9zuijaXTW0QCjvWpirrFslZRVFNG5Gs8LynT/CoiXOP9
RSL+oRPv8csH4b11nP2BAUTFnwgRJHuGObRC5Lt8KXEk9R1Uxe3qE4j6jsfsseH2
PA44xUbxJg6KmgU/rhdujKaGidgm7I1eWhAAxMGoeMmoNaorAzgzu590BZys4dIa
IWsEhK/RrmPVx6b9mG+NsF5CGU7snAjlF3/LN08hkAqgSy48ykHnqPd01ewFallv
/1h7zSae2Peyt7hwTZXoWRQioXgNsdoI8QMOajpAaDRxaYzw7TCKwBd6DOdHKoKA
BrR+4GFG4sF/mhxfFFMNYGsXRwN60GEEFiIYLqAhL3UU4tGHgiBXwJjO7gnqKF1Q
uv78WNQAsI6jE0O32XkSbKSvDGFJ9suNJ1y6kBh5lsNMm+R1ax4BB7uTGlWHa9Rp
UEK8ETflgRjto6yKrlN0yCoitDjpcI0Jg2uV0sG1vxKqUj1O5EzbSCJj3Tf4IZwj
Raou+3b+xH2NEIS2ZCukrqp/vnEuk8ViiA7MGMJmv8OjA4noHur7L0LP2KL6hBzq
tMEeulq4zt+e+uvClPMKCtujXgbhQUKIui9jFIjKYvkTIzsoU1wA75Fj74wvQlDj
xNJ3W6+vm2DTAwWAa8NTj85PNXHIXYFnF5o1vd4Ka3kOWFFPjQJAx47vIjmRw5GU
ZUqLXAq5fe3wzBZFOiHeixkJQf1eCAPV2eq1HQk87/RCCGjDmCR/tUpYpSI2UtJX
vLrwuC2WRkbx1awUbwnWXt/lWyw4YwvPAdVMYJF3NkyC6NBWxa+jYQ+YNb94MOaF
1FOsAOpI2Z6rKXVHfrILu8sDSgBRdZB9tEccUYkpvWEtDFI/+Q5j3hdhts5X6EHS
sqTKa8L5QpVPuyH1wf+GL8JfY55p+tEYHE9SrYj0VOvHLUVBF/+EekSonqBwOkPg
Rht9kPrSCwikRPbON5vJRGDbiSgfV7ymlwzrSHvMFp1wyXk7oUjRmjPXCPkdfZfB
XsiB1QvwFE3hEapOou8NYYDMXGWaVL+uDQl1yK6r+X4kwE/qrJ5LGoP/T/Tzgqn8
pta7ehX0mdFiMMA9HkGOomcMp9qJPZF8xToNVfWx7WoZe1K6g3aJCFPiB32w6BBa
pUivg6pIog7LBdLqOIYnTNvhG3HvTFFw3BSyhBxIX616qGMQmxQ2vF4QhBIRcEP8
5iiXDs5l1L/+DURQHUBtNmN2cy7Mi5cstiyCG92P/uJh8l0kGLB2hAkqcWzThg9y
bYuy6dN6X90txph7ofwW37pcCUTC6lesom3kUpk5Xhzyo2Q8qFSeJNKDdbgmEdNA
BOqBZryhbhKnJGQgtQE3HQw1HkCu2kR8qNI6c/qFCoplpKwgFCC6gwKHetBgtalA
5e3ssv/nZywKx6kMe/0QshruuahgQM/bIzJSIJx8NtD/qrRN3VTsDv61KsKBeIlR
/2SDtchDsMgnCEaeW0qJPji8HLz4fjwzzqX1nQxZ3DJdEhQHAPsgq9N5ZIKX3Wbr
7beUL7IXZmFmBzMCnioITkNY/9RoM4YwC4Ep34JXiYxaKC76iDLqC5z7idxQu7Aa
i3GdS8CWNw3tzbCszc7zYhifRyke25DIFLmRiVKuAnb11hvntNTsPF86zuXMHqEY
yYjiuop3QlVHlvlbZ9eIV/7PqHFxTX4KQmRC2urwUrQZkF40AB9xlbPePWK8gTiJ
BfO3dFqg4k2KvmuPRv8Gco4+20mrkqNEXhhqyUhcm/xirr9GE/Cg/4tfvy1CSSUI
gWzS3Od872BGaKAdsxnxt9c7gOQkpv40wCdffQV4qAXCVZWp3GcVJTnJ390FotMX
gGuJ9+/zEyLyVvKwcdy39SaorSnURiyyr+mYjvYrDsmJfgcC8tdpRqQL3E+uy4SR
10MDBtC0PwaJhOH/E0o2l+V1g4aAmy5ISJCR797jFbkOMOtStpi0NsTSu2Sj3CPY
SdbFKGgmUBI1wMrsUn9VdDhXuzCccH3/bAmsGMfN2D2/otwMfBhdbGW21BnKAU/i
ncmO6jd4X9ItVsPHcJU52uf45Z69SUbKa6ABpcweXbBCy7lFPP+vAf7GS+n2P/Ln
YYgm/1cNxQZRiMK5u1jr7OBKZMm1jz2ek7NMppoU5VOSmRnyIGdv7nMyAO2X6Cyy
NvaNI3GH3+oT3x2SkKkzMNjfbIcAoHwNS0Sedi3MpdbhtF6iBGY07y0XA4zOXx3Y
fmB+UjWtEs8v+O8vsKSapIsTsYIk3Y529Jzbojp8Id42T5IIUmKmTLW9/wPw3qDr
2nKDLQ9uEVlSsQq9hTQ88lzo01/UVHhCD61ncTrVYD/y19RXAGdyAS8i4VJWM4C2
1Km9o3/+/vezTCM4PzwA8QXJy4Y1rJmQlDsKeJWrtJ5kkPy/b/KU9cQT2d02jYrA
26/nkPNLquDLDqWckIWP55RmDryv1XhEEr/3w44fCuqgP8BDEW34wX8mttOuJtoW
t+A32tz7KqGgsH4OErU3R7enuZXHZBukNgVWyOMe2vXHbnPktcRe+Y+9TjK2xFXZ
hPVy7tNm99FcpwILGoEbf9oJsvAJINTG+C1sfIIjej5Y/MmibMubbOewv8jZEkmV
76n1rvnDtBED4kcfrgmanbXK5I+q+wd6LKYRVwBLLMhvC532hZ2xdMSjb47l+OmT
HoQnXMw16CgnsXKEihdFzSbL3z87wWraDFnVejlWgFxWqbbCyvLnCUEjyYn52w3N
3BFGS9+i0ldMFUSmnYEjiOvpwCdP2NKXzatf9vtA1k5+JY327Xbic/gKLijhE6jA
u36TW+zkvlvKgXxv6VDgQvnIQkuWdAREn6L5jMc18Z4iD8RLaNo+b/c0WYuTsUFV
x5sHHTS++qdFux40lcwxBb9VA55dZL3ctb/01V+lg93a/i557v95aFDMgwy/WZDo
Gois4YwzoNRrkWgXHA5Ksoo30/M7drp3pTsJ4/hmWuDTsRdF86pc87B78p++wdv+
I5wPkw9IIUepsfZb4khpS/EBukzPTmUJrLzCe+m1XP6hwGeR8ezjDLoDYM1fM0Ud
ySJdhmy1nSRg0Mgoa6Vy+F9vXo+YnowE2z47RcqQcFthNE5b86230RvJH8IcjFUv
I9UZ6aKorYFTzkzd2GXYu2MwWaXj/L21GQrDrx5zchdk4c0jsHU7boo+w6mBltN+
DkiKRR+zHnIq6BpZ8JDKWaCLVKZRb6CzYpTo2Vk+P7l/bGZY9MgkslLSogXuXIaJ
HVfl3lPUQnK8EobT3NeFXz3vPyGy8VL/UYfZfDU2hNsJ+OUPZVmrzAT8uEqVN0sA
OOKhfnhFfZyeqhHqL24SZyGegWl5RvycmCGSsvAFDguGr7i2wiWcLgZdngkiUWX2
kTG2XydbsZ4oonwdlx1MmB3LU4KsyTmqP1pvzzXfyjpMxXB5OSItj1RCvFMeh70g
+4rzIRVeSF21jChkUBOCNUKbl75ymKQi10AAyFxyNIDc6llr0FWdE7K63MDSt9yM
hf8scHT5vzEfbEV3zkeX+djx5TeACudY9Lg3K9ZeJC/fX/8dAlZK54Ou2/PhvlAb
lZzu6VxfPSzAihO7mCPekrXaIVcMnwJtkGu9Yf35ZOlq5r80/XrpgV8hTWENfuMP
RzwTIYlfxf2fJFCWXIrUARl/aKELRLrnKi89EGkc7r8t7bgQdQb+ZXY1kHirkR1T
qDpMJD1jex9+sbi1QYxcRArYoVSzlqATafHl8SR8N/bm//mcdcg6oktcpRTCGYt1
pfvCgPsRctYnU/mDNCNlON8gCTl0yMGev+JB30UzIvZs9N4yvFHVRkEKdEmM5OSW
56mbdZKQC4RqdwM0iDoPf5zewK+3fP9Mjbe0F/AHbzdB0VI1+nfzQgshw1klOvQt
IdLvgL9POiSuD06yupAzUlL4C0h0/FSXb3+xZhg3ntoLfkkRH0nGKxq8I0wykYLu
wbrZPRvALGEIGOrXk6fojEvSjFHSCrQSG3vTmbCma4yxwnIhetq64W95AR4c1KoC
ouIUpplAAHXTAItEvZr+2c7Y781zr7xti72Y+BjIi5EG6vOTidAYOMegg3cRqXPF
WcYQLQ3tHeFMN3QLebVxAZzdtr9FysFLhqM3qmUWdNSbft/zaTd+nQJ5Q/S4cfKA
lzZ7SheNklcKbmn3gDYKTUEVi4ZQOqikO9B5m1JteI+T1oJVemVzvdtOwUIcTnPQ
2RYdtOizB7/zyOlC2a3Rjldd7YxM1L6QvfO0Qn/ZiZUiFtWyAmvQuNvOr9BYgL8r
1G87nYd1FiqAfHEwYPWQR643wMYtLGVzLUWbog7W2qs7xeahKlzRuIoP4XM69gyz
rLcjU2z9i43wAPIhGoWPcxyEsQCkRxfoepm6rpOykto3S5z+k+aNLFnwri5botxj
YAFCNr8qr816p5Z3RddSO4KCJj2yl45Rx9EUtJj3+OVR0/z98GKXwBTuhu8gdzTi
Fq7JKBhbSRgrg7g/wrPVrTKbjfcgUn1KqLUgtQtZTFQlvxdOCW3dEi9EvdeSWgfD
L5qQETgjdI/lGNXqQ4/tDG4DMWlF79rgobKhcphUXGL1d/2OruNWpVZI2QmAMcyV
2gqDo7ODq8vopmJzoc60R5zi6gWJr9zv4rSYXjJDf/igXYYTkfb2xBvcYWVIapCy
pefOjj/3NQClVVbwtn8MqP8/5LbVAuH3ni2nCxUBFbgsy1UXv5h97T46IM5H5L7R
igjXgN5kNhA7e9NfVLV43J62sY75fRgQ4FAVvitOdd/pQAeHvvX7VdD+bWfTxxcH
MQ1+hhnf+ogc7bOJWtne6CeJQYQ+INqjZIQ1h/dAGB7wfMtprSSMHPG/RitHC1CN
mZFRiyZjsU/Vqat0DuY41yELqbllPLvmbD+14GKinLxdqt+6BTXu+DpVEO2NIldG
IcIdOaHXJjsTStXhWkAqhrTSLk4JUnnh0EAqtVHnovOqwId4fOdi3kEEPErIfDVN
HgYTJy8MWnf6d6735qsW0SIKvhfsb7+ZYRJM3AAYfouQ2nVh63g2aaEP4jyM3TBr
G/rkosnbpHH8GekNe1Sou6p2JuyTa1+M1ojuPLm6pfeks4HSLul98ZHc/Pgia74U
kJoRZXfXH0AZmczaIP6FwGQRm4gxoM2JxdHtt28lqmdWOdtDTVA6aNTDVU3V9RVh
1p0yueX41wbv02ztWQruN7BbA5NFf7gifdgZ1RoA8IWG1uIk/QARD4Btgc5aybpH
x3QGpmVpEUIHN5SfJ/zNia3xfYP9nytZVT5CLPEl6Q3x19CY0KmpTwgtk7sxRO5l
OfIErnoDF+Q1tLhUOzwl4pDRBMfZ7/RRFGslU7k7rgYAjX+PLTxpfRuptcBngk+I
R2uoGQCBn3EJe2IixhjeItwNBtLB0VrWAIiR1mDMa0/SSco+fUFKmTN5cz1QrGi2
iDyzU49l/PbTDMFvuSgC5K8SGHt3FcEzUyJPrOu7MvPugZYHzGpU6BD3amedYiL4
TvlcpxmnZmoQs7OvLW912SGMWSClEWJ+SJKfx3wu5kb7avEbE7Xpw2XlNGtzEluC
TogvFA8rcYjBg96YW5LWKLjG59dsYQp80qSvl9fE31iqmAKWjTx4ZhD7DVG/Y+3Y
xOc1aZhSGGKpLaBidgPtjmxCIN/iDoMH1hK1dThJHsLJfKoS8B0PTdwOrtLDXH0E
ZDYDPBDChrFoceQb6BsigaxYAtr9hnnFdiOtXi7VqEmAc4Iimmf0MCFSUFlNvifV
nzOmSUosN5vQf8QdyEH+xjDGcctuStYyTt1C+WX4cmkWkxngcTQ+L2p0aqLRu46L
UNHtKz0vdVBEEW8qXBq6DWBLnb7yXoAgUSAxOl1+1IFUJf8awsPcd7gPuQ1jnavF
7q8Ye9jPMVWCa3N0ws7HHJ8Zp1QFSoTKs/+FdGXriFDs+SGeq9yYNUyGvZ277G0o
x3EUJK/D6kPOYlSxR8CX6+ohwKUXclTOeSUJrwVmboQOrQ1oazEJJ3oQmL98jpr8
FHOwTlJfIoQ+slap+8947QjwtfklKeSJOFr/h6Etn1OVekFZ/tyjD2KhERjclsAD
aiLmH9ZePdaxY9Sd0+Vr+5rmmfvyqYKI039Eq53N9Nj8sfaADWECJIxfWSDL6+G6
rc5HGIqinD97iAeH7KyC0p3WO8PpeWHBPDOgwxQpF6n2VfVciU+VY0F9u+Gvot7y
0fX3C4cKjoOhLdQMy//DSpolypV+zdNEUXAEF3GeDPZz9yEMasgYTYWH/MNbZRni
ReJuERqNhbu7zhNwaL7HS9GUJef8Y3JPAR1+67qwMIxXYyS64d3jo3x9jwvekxin
NBXuakAKw4uM4Nqw3sAIyQocTNdW5DrJijywhQQikPWy741wIAfqAEVsQyjNb0v4
jWuaRN+vZ1zdCnnxNek5wX3whPrpWX5+v4Hyid+qr/R3JFudUtC+gDJttXspCbOW
pq9CaViDzyS5s/Z8eF7brT9Ngc50Fk941Be8eoSrZHg57hxAI8O63zAw6AEfYvzL
uy6PuUySX+73NKkYCC08eREJpAR6eMjIeE3gWge57QdOYQtb2l/8vWDVVPdhm1BK
8taRhcmCBpN6fUG+dzJythbDiltORyXd6tZ67tTDL/ZrX6xlVS6j1fgyajg6Cmej
qsT5qRvEzNOkHKVnOt9wZlQKeyu0CutI6IBQkhTrCOMKqohza84lRIOfo7TtHApu
keTJmNIe2omF++JHW4/nN8khdpBMscttJ4A2vatPAjrHneqqtDIY+mFf2MT1/6Qu
au4T/d6iqHyRJEt9yiZNeiAq0uBT4kINmdwLnJcgsi9A7+VuY73/3DNv0JcZArHA
xOKNvvJyBchhksMeNXe9IMqZg596y6ymvX0Vjsb5ZgA3mAHuT9kXe121lP+NKOHa
XZjbOVH4pZplqafGERyWafqb6nyR1HT3esSme/BJjq0NoY8XY/9e3aLXJasjKXvL
17hxLquB2wQekl3tH0mI0gk8F+ZvN0BzrdwGY23HKolWW6pCmEJ4swMCYqB9eGW7
zQPXUeV4y/OyF+Va/3Jrl4XbQ92nGi4G208shEraTjPj3YGTyNVjM+7kWyBty5iP
d/OGq8YU1vX0FJfowpaNkHtpThU3zXK239biDvGMnHUPZIs7UiSuCouV+/U292a+
YK7Jy0riUEJ787UC+B61z6Rh7s6Fm82Inb+W85tcJ545MetaC+d544ywXoigMeFk
nrknSiQpR6T4ZoJHMLu3tlYX8WO92sT2hWzKoJcm++G6E3/Sb2G+REzbTzSA6EIj
OsGaMxUZCbQaxWOjfQU11/j/YephXfGk6kcq8k9w4qOwCvEc6UqqeaSSH/YRKOVe
ej2uX53f/X1YCLMAnBJGFf+32Alg91N4IQjsYRFeMJPSW0xib+BenNvj+9GLy2g/
wT/7TpPaVqgxNp8e1y9um4/fqKDQU/j9ewhnmuhXXnH4WXtuZlb1hFJP1WtZYHCc
BWRUj+GhCkVhSCNLReE8QX9b4Ra75FoP6piAKkmEdavo3WtpRUMj8nODqOmvaP6X
m6ENo18R1WzahgYoUHBkG+dtDIu7u1IV+LzC2ZhND2VNEH+8qaNMj6XZ53uRyP6Y
u1X57beRvPiZzSwnIv6PAdodrI1tlp6WkeXHrWR8PMQOUmao3+CGN5HmEWJLIJ+Z
6FO9JJTYBdE+PxWnIvgWYvYbMTNblqUqoJjh6rjyV2mynNKrveSkARHiYIquqUIC
+gC7LMZWyDEZdD+gy/ZWC99qgNUNuevNPMhYW+MsBTKTD5nKoyxnXvGek2JmoE/R
JuRbaeIGZdPpQcwglMsEZG4boCboh4eT3lQKDd2ISq8zt2QFDWFLGVY66F4+rY+5
bg3kv5d37js+2+HEUaOaLYliTIoYTKHKiiTRv91cF8dmvwlm4NBJGXCy7sp7HNDJ
cT6gYpSbvxehXe4OtFwqRrMSBNLXOLSXuFr9oZJK4BCQO4s3TQU+n6z57cRCnkDs
Kgq7AKmb1H0z79NGXZjBsI9edH87iya4dJHXMR4OIygJuf+L4b+Ful6EXjxztIsL
Jg50Gy1X36lp5a+FoS38mNoyLqL3JgWxAjGDAe9Xx28qb60MfYzGTQAoCWElg8/U
q2ouf7alBuqdqEjvO4ONOtb+A0lhRWnMLuDq4IamU1y3ZYxky+/+J/bh6K3Rr8Rg
DrySNCrYeoiufobBKV3wutDbszGctDydr0GSpycgKtub1Iy6Wb6F/SE4jSLQy1oY
cDglGqCuXBLb64A+ltTqkZhAUim8DiAr6+CJA2yeJ0BKiWNDigzJ54GhWPA59DNh
mNxOWe257dXTO0AWCRwZOucksYxcSpc88ekKSpkpnDEWmsSoNigW/Ggbb5QhVnrm
AmDaHBdESGzsplbHFZ0UHcQaZePbGQQ8/9z4t9mtP29zCod//73SWpsLPIG4CW4E
SGGRnXJQpc693I94eyea+spdhl09uja/u+3GKZABeCKy1rx0gYqtUkhpsRWoh4dw
bjw+xro851Fp1J3Ucxq7jEUhUet4Yf5VGTf1Lq0yETo9BdV4wCr1kSQyXQqhSm5Y
qFlqrgVCxBJRC0Ia6PtDj9DUQt8DlGbrYIt2h5+KocTZFR6U18elwNgTtDGk++g9
rWd9yE4YB/EHU4ucmZY9re+g+1TENuz2J5VngsXnkOSwfPZQZTJDzX9TC0ULGrSX
RGXMl8zWhYN3qaQDEvNV30KBigDXpMeJ2fTBq7vAZPes2t7K6TEFG/REoCbIHKpb
0KTBqqYD5e5ey8JABrtmSDZou71hNcVLUCY2ylMRa5xrQ7L5omiBVfICFP+l85Fj
i0ueqKQu/EW607YmkQOHHk5ri2I+uexynnjdi5EIC01aSzXf+admera69g4XpWZG
eqpKeZvf01I31+PDxzDYueVWcaHpRJiI508v6lilY5XCrzXy32q928pVIymNGHek
Isz9CpAUVbnVyMLpmRgQT3/Yzg05OdXE9Dtq4xD5y8XHDDpxt0cUUJDD66mPWOrP
78/hrDdHgQq306DwrsHRET7TV8uiuqLOEPb00MBD09fG3X+H7RSp5VJMWHJu8Wh5
3K4J14wG0IYD/6ZS2pPuUlLlGmTUduxZU8+508fDzRlIO1YubJuDdMbTxArA/O/p
tsbOm1If9bFFmtIi7Sv7vn73LPOj6ud/936tT5bRRoJwXdGQ6KQtDGFv0MZ+o+34
EhNMnx2raCcVm+WjuneLtNQWoCIvIML5+nAbnilM9p5d8ydQNzrHMPrMEHFLoR1K
fCQZjvsoeTr3Sg3Yha348N9JjzPfWDtqF5zugAOvvGnQMLvPjb0cyTAtQ92gxMQw
DJmJb3US22fg5uM+nB5tst8KkqLb+1Bd0V01IBaxONr7FXR9tB7Nc3fp3fen6zPP
36rebmKo4hrvuOd3Ap9wKJwfxp9XdhVGF+y6ZdyTWOECQ//IcZ/BlatCsIOz6/fE
T5new5KVdBdvYrDCduu6tT2Y2OEHe2pI/0IaiEDex70KaTBmY7IxYeaTyPwkPyEs
wBFbDoDItWdkUdn+tbWUAbk6Pu7ZASyirwL7E3tqE/AfApz3AKmUSDUAAEe9ARXK
uvfRpyGeTQWZ36WjNPG5yGB4x3MuuuIJrOnwdS7d4//tqirYde9t04jeuOlvihXp
cI0MGcxMSo4lFXdxRaiMxvDdQ9sD7MDo7hWXW/fCYbzKXMrwWFASrsGe4mIqo0y3
7dwMLZ5xQCL8MYmsMQYd5w5ooJDneqFfxTDkKJuUAlW7Q0ywofJgA5wd4xncP1mg
OSOrdjbOEEsT0IH8XFXnabR1bW5t04oUrg4ue5RdeBnwKgzxAWo3TTd3G2SfNhvW
Mfcc/SebeaPcWafHL0SPVDDHSiuXg/HVGvH98p/s6oa0DVP5kmG5OEMemdJx90hg
T8OXJPiR7nbGzzjjJGTffkSodTQY9US6S5yfu34uk9QG84WF4H+HnZ+XQF8yrzYh
+GGDz6d597qL0XuGxCy8B16yfmds8e1XINcRxnJuXswvR37G4LrbrSiGpArDswjf
8fbsg9hA0g1gNVS5GTLR24fHEGw/OiIP4XoIJnHvIN3EoXMpsgCUqJ4fOMJ+wom3
pDpcEVK93zQoSphvgoSkWNAXobqP/6tu1qZtMmOANav/ufhkhoX150XZ9jE2v4Ak
nD7Xh/DPCCQjdKzj9/SwPGeF7Y7GpfUqPgbJ83t9XFrQVBug7TJfM+YQhP8U30gR
7UkjPBkm64V42OfJa3gH+Z2SaUDbDRcJJKR+YFUnAqdfLytow40G+PQdrADmfXuN
CgHetEbawHey6BaQq2O9npAAiMcbpSvIp0C9jyI2Rbu50E5aISj+q2MIhfPOcKWL
QGNx0ko3eCzFYsm3b4vwOP2q7cvi4qm1MXc2hgZXjU6nYOCzwaUyOQ5bIpNMmdhK
OjlFmyCVelxSazxNk1zh0SBmW5NSAg95U5YojxYyQ5x46tYRVK4EzciKJO2Vt8Ey
jiG7cBIhNTuSAjeWK0ymlL30zLOvgWlfcCvolGiWv8UbkzjXLLsR2ljY2dW+FJT0
gBs4up3zVKmyTUqbkBZqtnxE4riS8XUX1o3NCmfCMAZsGWMihIFaRKulvSfJPfrP
h5twFzoN65dZtE/uEcDT1MymWLmwcWah6ZTE8dIXJeVrjjcF4qDFXHNUw0ZdGyuG
gBvoQfiQngYRPa1Q1aOJ72uOKqaRJCCKgvnDiBuEZZ9g1iwDgNLQiUHTIVTz15yp
RrP12I7bvfTHiFt5HNE9bNB3UQXw8gvLG7aLXA5yl6OcT7AqlUxNGU/w/VOJIv24
IBFFCADn1kDulwr+IW+Ks2eVBgD0pB7Le2awleXSIAlwvKQg8Q/kxdu5ht4Lp1Oz
15M6oIT/IPy6LFLzzLud3sJJKJX+OGlgj/3AS62IXI2J+yC5E3d5nmeRtWDHfsG+
V6juB5vxQtR3q8GGHlMeSN2auF/X0IGn07hzVnk64nO/64ZwLsQQrzEp1fjtW5+d
tsarFkv/7f1WocSd5FP94vgxZsnXypO+6e6317v/5QGv6surjd3Z8T2sEiwHQ2fQ
Kogd8RI6VDMclZWJne4Iwdcqf9CDBVc8th5esWSTRaParF6oE9ek5m2q/YSqJSDQ
GS32c+2jtUETIplB63gnvipZaAGL1gCHvT/APbkUaRVvPbhh/YzhHoz1BP61Evaj
Vf4wV2BcRZ8ayuM3XOBcwTEQ7kiqJlcUIJT/IZrtW+M=
--pragma protect end_data_block
--pragma protect digest_block
5+a+3VM6Qte0MFHZYzf7R918aWg=
--pragma protect end_digest_block
--pragma protect end_protected
