-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
hjyxfhoE5paR56ZQrblYQNxARmZuMvzZ+RRlRM5MwC+oPPzw4+trEDcjTdZbDolv
keHDKNXkgsZdBd3uEQCcXB6uiUbdhh10o5hg6GE5iG0hegFe1EeisjwW8/0efJlQ
V4yEuf48ZwGc6G8Mwq4KERuDWG4yXxjFvmEB7jRd3E2YzI4oWUYoxA==
--pragma protect end_key_block
--pragma protect digest_block
86syHlB1eLsFfDWkG57IHAyRK2w=
--pragma protect end_digest_block
--pragma protect data_block
UmFGwHraunQ/f9JHn2q8cbUgcQuaRXrKnCxbJm6naT6gzNswDgy8ptM6M2SmkNfa
G7Z9/dUO8gOmL+7gflCyS5XQtJpvmpqnH3MBl9BOFqgQJIep2MxWnQc6y37PYADX
ltxPLmwJ1pIrugq6oAYicJ5mLkmMHPmBd/PrQl7bJR6a/mMiX5R7IndNF35NDn2x
El00eKcdqRSqcqoOClL2ifMWbc1q/RQaAJuKzWIwzN5wp5jGCsiNwTeo57DbFNk/
Ac5exoOXAJBupmHGb9cH8JknBIRNY1uVRryj0mqhps6qX7l0cTvPpqMiKiMif9js
NQiThfnIOEN5RIwfs8Pq5gQYt0/AN2B1vNH2EeZIOjv8uz7EC0cM7KV9D0k+8ZU1
pHiGZY0X0ky6bQx87uUWoWA+WQiU+4zhg93oU4iQ/0L4Xch7MQVhX+DrlPXxYAgz
ILAgEGAt4g32q/gJ3lQyCyHsIfAv177NTLLBk8aL4hU2dG17gBknNePqv5EAdk/2
eP1tvK7bNPf47mFLwNr9xWYgvPei6t0RKaGKfUYomG3xO1rW3dnJ76lHW6M6gjB2
/w56lSt8blMHUTlx0kRDJa006fIhLjcEViOIBRWv41DoHULXg8GBrUMjwq6tmLps
CwrUmV5KqZ6/o+ZLLEU1M6gmGs4D4YyvrmJ23ZFygG7tBfbVVmzsIGpzsfBxggxu
nA2zfsYozoi9PBKejM5mih5Ss4uDl3xOD45z86p6F+kC7+nhUUICl9GL+05WCKSg
6j/5zrucXgoEeSDbMTiPYRFuEd+QuNm9EIwqsxf5cHlLP4sfvrvJMWAjIhDk2K4U
9/NJ7FW3DKxNHrE4fXboqd6UZjnpRkhJjVFv4VcFuTsNZwTgPaK0nANTxh9mB0zR
1mff9KS9uS5Lg+PdW2er89qrgWkUPtp8TagyU1iAk/mZdSQGzLcgpSOS8gLeMoWf
M3zgnZw/LnXjeAO0p7toH7mAn/WPbfr+9Cogd1fl4TZg+EEevPuQ5BHlgrSrBCWL
vrvk+t+4Uo0vzOfsG0QiixshVoCqWJoVdyd+IawN2SbYzgAiE/Oj3d8CjSvkGeqV
wjJ5Y39WkpipGmZ/3e2KdTJGJT5tdmxusJWWAKt6AGgOucKRLmWDtqxr3IU2S2ni
WDXgQ6mzJiBJAYskQ6MMoW0KNn22WM94kf2pIbZdK0+JNi24ENucLPyphzdb285C
4qlVNRlxWkbqpN2vtLbBM/LGXKvYfCMLwQHlMj/Iby923dSF2ylefQK1e1RAm3d6
O6tPGBBvQSaXAHFNxf6tpVdKk4G+IYh7K1f2UHTKMjz24tNLBJEGcQRNJr7k4aw/
Z6C98IlGbMj+71d778lg0Amo9xCkoM+SQZYdKTUA7i7hicNu/O17Mlhq+YRW6McR
H5fzHiDsGk2MwjglfKI0yUEm6pOSWD8Az/a4BCYiZJjx5sr+4oMdZk/x/JvZ1fMk
ckI/DPqqV1vTusJkAoAb+lPKbNDcTY0l4zv04FgUXaFhT63rkPhAlRvKXrV/Dztc
J0vX/Df3ChZdE88SuQsNouQZhzK2jpErRTofTbVzSqWCahNikPGRnCb3YdNKtSOw
O/OfpikgyQuBRrvRYtsMbE3nLQ42QSn3ol4xvgpaXT6kWKRYbosJVqZ1KQ/JybYo
CVaHUxY5wT35xtNrBzVv1RGZvzFftRhahHA/urRdDHLZwKIh1RDSSJeZVlsDPvVG
50rFsE/T1wKv71ze5ZB7tN76NNSd8jNPzQuq8a7aFEeQEqgRwFF+6FQpeJWeesVK
wILQXIwgCmwhgG+2ZA0MGFZP+czeDun99aXtwXHzVI/pvaEzHr3JUigDA+fhjPCI
3hcKe00pKIYo1Ex0bo13bVV80AAXjgrcjqfVC62O4zjoFTF7bA2xvVyKXtjqGRX7
PLUQayTYamT6fw4QDaDPdBEgBoVRge0FFWc93h+QPcEWfSt/gidJfgeJjUTsLglE
pmxYnjP5/68ZnO9zfnq1Dqxn0gqmWIocQ/KYvbdITqXXSckqw6TZ0opuOmxoNXIJ
AUnPQAOA9DDgnnksOe0Z1wpxHJlAXOobIk1/4RI30ol5j9G7tdcsFtQiyTpYgtXd
QoNH5XpqM6yaz0WurqOk8dpbrnbTC43xVPEvUt2EiiD2dTfhSb2L/6DdI4hCB5YM
VLeAXZD7iMTpC8O5bjpZiWstdRxGe++fA87blEMbYZVMTjYLZqZ4AFg+rWHOJmyZ
eB4ZVycSETuKNmgvgzaj6cav8+P/1EceWtGQ4YNjxgXlNI8Eqka4KzpOLIHgtgPK
ywLUP/65g5aTp6He1KNaCaNYGFo9cAEY8ZfnSf6uCIoltsOarq5qYGTUdTHIYr/d
lOVzrm6T2hbwk+6ZxzwSfHjNiE6xPh5Q72YN/7DjhLKScD5onUmyCPAzWnHayJDI
HrYGB3AUnsKUl823uS9OAcRT9852mY2NIUdWlKC6Qi7OH5nBf7dKqxnCox0eXGYq
NEX2q41g6ldkly40NZpxw8rYVUsfDQjiHgGQ70KnX9nV33Xi4Gi+o0jzflb2GFP/
m6NeUCKouPuroV1wtv3DiYYrc0wFKlxIIA6/MWHcO7tW58+xwZkzZ62frfv2ZBjv
N6o4cN4GttsxTFz61y9H4kSpAIlo/r2VGCsRFDaDeRc3lUS0Txx9gXVlEnQ5d+KF
C/hkTW7alBscD0diExJsUIyBnVmuuS3AwGSOsLFUS/9EJU5Q0oA3sUZEvv64vD/F
z7Hz1Wau5BLsafsAURV2INw0J9OeG1WpzpAx8fqUHN811LfqmD2Sux0KGkNKU4Bp
zq7NK1zOPnvy+ee9UVQG5HlxcMPKyWZpu+5C/3IiPTHBZdycVSTfa9se48X8AMM7
E33IXQtRpIIaogNsB5ZEhYYwUFfOztJV0l1kqXOWxLq+BsKqrDgYyFw9/GsX2B1t
DCNIaOiYK6PotKvAoGlgthaWz7BH5zDY/CwHfLoyEf/sn+8S6Zg3TcdeQViqI/UK
T1OgkHlwxVPtOwRzb90+Og3OiErB/WNNciNAoByYfyCHREBGDPOtceD+Umf8ibWJ
xTfejf2wlPZL7zRNO88KHO3oATMnOsH5qezilPP9a1UsVIRSj1+vupodUpjScrls
xjgxFnAbH63xit6mlnoLFrRYs84bf4nesOq3bo/P5CyiqhXH3z5ACET6ww/+Mfgt
+TUFqubrerXs2ReMd/V+EAbbSq0zBQGIXkmSnBW8aRiKvOJXqWWhABdDs+nYQssx
GGOU9YDJKGMlchEu51Rj+cvkVd0hyk4AYxPSXm6+uvZMoA72wX4T29S5jnJINWxw
Dxu+Wy/jj/94WP5tU72ZSgXbXePIKyO6yx6YlPiWR22cnz4OTlBdwMNIk1rmmb6w
V1wDm0Cv/LxUaBcClkmLJqaEPMV3eNNYL8KlXmkpiU+VZR7Mv+7FBqLs2ufY2fPe
xyDHXVjLvb3kIc0g7eYjf6vIXHQQMsUkXBb/rNiFQ9ODbnvWb/mE3HGcTqWEd9ff
raQee0avIig44BGT8ta5Mh/fG77rTUpSVRiCpAdLq7r/2I91OYnLjmm0iqFhlwMj
XS6xfueO4uiW2ZPhcxqWCDZ0QDONlcQ8Y+O6g/E38WED/h6sEDP8Wu9KXP5YzvN1
6jto3jau1k2G2DdIvrVKWaWbQUmdEgJ8ayRyfA9rfJDoPejTAbzmquqbKKRAEoBm
eba9ScSyMab/hgeC/0uaciAyAyFb3oFvqPpB+486IN8cSZY3w59SkYgTJKLso6oj
fGkY87+WdpKEqCfL1OeEjMkp3+P7t/YVsh2a5Fn3illpbhxvo+QwjIoemuvhIIR6
y89DZe8tsTKs3yAZ5nw3yOXRnir1kNOpmDujlW0Q+zCy5ZY89Alf8xYV3ULmrWgl
yN/OkAE3WbIFI9K0hqM9ITKjiWXDE6DXovFWu6jgmW9j74WQG4FJnJY2dUrjCgFc
iPWfpoWX7HCDR61gYEiYypdbrtbpZtqJSuowcmBQ5dfOcDQPQFS6HVaHXOVfqhgn
uNbr+R5RIxFQvC+MB1umn+H1VgSCq8LYc/wutE3y2piMTIoud/w+QB9774ohAmKL
EIVJZ65TcWhqzNAUjsGMTjgZnX+jBcUZUugELjNBmOQYzbPKGAhyyl9TEu8XMTe1
41R9TM7ulxZaukfiSk06arl0nyo7tzBONo7A5V5+F717V3nAAWSmqDtST8KD6VSV
TCDCksJOU5FJ9VhgWujj0eAf5Rhb8cNoFexVoodDoFY3wObKc4959MmRjUalmReo
m+na2qlOVDMbmwH2iCBa5jS2BW83b9xddAhbLZHiAstPlLF4ra8vQCyNG8bSxlVE
ZnIIxBXPIYVLKaU40ACBWhOkNlw0OUmcGCW5bsIfQXuvl6VM4+Jy8ge+1+dWYnAJ
FNPXqVIEUj3I0PbZRVEb547FW2Kp81CkRkboEQslVxZ6R9cER+czlqmINRmhbctQ
ugB5clIE4im5fL6av53dF8BbLrlzSJU0FkopfnBSGVcZlKItH+eI+Ko2ER3iNWbY
ov72tNQwE90+VCGHNln+8lorVpB4jpT7JtSx+AApN37yXiTUdku+uBKK4bpAJN4U
UWI+cfSrIRmdj66oY1Cvliu2qAnxdpQ2kbSyfNvQfNzCWLOoUb0/hcR9dPC74qmw
X33JuJPgHgNjcMYKolXuXWdq9VVvX8nG5x7sY2HpT4+BZAOE6YILFx99IrBZbakI
rdlCsjatAqnXk5ZscPqlcVu2nI1FaRB4EH8z2kzRc28cPkYojazdY1cPILlMiWFO
88YDeCUW2BiG4HZKj3Btu7iQy0kON2bNWH3osQN443EEfQA2p3OLi65R4VEC+k9s
I+LTRk9BOgV/dfVJUnyeaCrHUcDGa4jlGwQXeF5TNGv3YhpVZp3nx6zkFlHhAizu
leTaA2KROEmNIs64P6yT36M2MZvn+N7/i3G++oU6cZIthUJ+2XlIJlGbQE6iV9tC
XZg/XGO9T4GB9/Int6uaGu64HY8w/rbeZS/1p2u5mnUTDYpET8rTYH70z2vbO68E
idQlX6xV7velBgRuwLcwshY9sD8ktEzHy05gPHujP4L5GtjuuDnsk3MoPh/lujZL
f2ZUb4SgRR7Q1BpBR1kIHBydC+IHduqBkOk1G0XlV1IutDAaedLeyn3iOUM18IfS
GqWSGRsfO8pWfM9A4lF7mhDPiFzjbEFhRFaw6cIjvmQkIjN7lTe9K86OvM+6mlQ4
qdV/MPgnm9nw5KrBRduYph2a0YTSQnMxt7bA0JQ5/pljncdox7/0m8bmGxI5kE7v
Ci5swM4a6jXJYbB/S9ch+hff2MWldUcrct5uftdoItBKwg4/tv2yoJijHxFlL+sP
iEnWOpMoSQ6asqOltsMbqITlPkJlyt5DWlMgYo+zvptpaGCcc8+jHEYGpOhoutLV
tq5R4Nk52KkjFEdWcgbtAyx45NsDNDImGNTQgIS8lQkoFG/2L22s1BuxXcHfItGM
kMpXMgfxMl9QkKaO0u1dlPCA2EXu8dozVGlpRdAUJKtzsjTekPhlcau6QhxUTigz
W6jok5DlQR6jEGKyDHS2p+eGEmX4STwfdekRn/gzqpHA+kylknHJ91BabFbwKxk4
7lksZfekWt0PIEDk4oosD1+GLUzX2inYZwJsB93NvP22mabyJFQPt0uK7Nf9jo1r
9QTvJk5MEPh//ifq+3gwHrCgLWHBOaLqD1V5ckX1JPnzDEG5vuMfoQ4BbT7ADB2l
+hV70FffrVfehmUjDP7O72f0vwYfNbaf1aH+pOaDqvVkyx14LVKAq0FBTfcv6ZHc
y+5XzmDDAxKxc6hrZtSAM5N9waHJaFOsBS+JiTbtMLuEHaf70ulop0IRruIvO4cL
j26umFyuLiY4cMaDDwDtNXbdqEzEMGn0hx5S5s3KLGphB2V5w0fENu81YTeTpeCJ
QTGJApmUiGluvd1ppEDtFXjzoekk0l4VARKTtmShFZEfBDkNhBSoCPY62gv7dN34
/cohwnihpHr4D5JutPbTf8jaTpJFpFd7IXoJtNy5C7M6KB6y4fLTFezGviXkwzQ4
xh5E/CdwOI8g6cizJOHpydFPQeyJaehthX1eErnRBsIWE5TUZiSN5kbEeYJqhQxR
Rdb7GM1/w2yoruf+I+65VpWf/nE9lPCREURDa9uZdeQYD8fl6AQkoQisPJh0nNSi
N/8AsEeLpgOiVQW2FU5jYvrBbwvizrHx9ONSFlcJuwzwldw6JZwcev9qzauLbrv7
f7aHM7cUj/fsB4T03muVodNQu62xYwNwMEDWmBiR6V79LG3TKo8jA+06tdkLSx4k
cFsgzsB7NcAxyDBkOIcHLik7nE/isVPbyXHvmtzNwwcYM2R7hmEQROLf4lOulw1J
P4aLKLA4qJkMQSCGT5IsGxsWsgd9j76MfDrOV3/k58qI4Xy417z1WQ6wOQBSLt5X
/GuAUW0usmx/moDQTwU/e78Kg254Fr7czOUW+oqXnqXuE1M6jesXdzxih/a0Ej4Q
vHBy3WwW9E1GopquZhroVNEOCaprj9zdjIVqWBnjhdJahQHpCHA3IcC1QjkRQg2H
bMZi24bzz80yMxUH5pCJcMpzdCN8NZY95zi6n//zLkJp+gUQRj8PE2fhFKCqlDID
ETCk2jzBnK5hH2aCnnfGC4YLjxulHlv7xhScchnteBYZf4mYt9VwmVKVsKk8GNBZ
zsKdU+hCxR8aYfPGJg0+W6RDnPkiJbDvBDlX3AHlXmCqNprHq+GBeVMyevXUO/X/
adPczZTmkuB9UtlnFcwspazPRevweA6luxsiJlzLMTLpCQxqvh1U26lnZz/unZwA
Qf/WRZEC42akxUw/IXW94vmoszg+cROFLO1AnCQq+kULJ3+fgMp8OKmAsrHn2bxx
HSH8DLNpB1msrnxlQGf//5TUmEd8y7OBaz7brk+lnzmfOWBrv/IkecPf5Usp8Ill
k5PHxVpA5sgVdT9d4ZTfcWEr4Y65Wm4OBtMhIhPt61psjQp7LFftaau6B2S+eXfW
pnNznKzFrySQQIOqDGwwp1O+LoJZbwrfEjQkNpLEhRdoVoVNqpesEcG43utQkYEd
+yeCD9KWIDYFea0enRYluOG4A1PDo+VlnaOZIww6Ad31MUZnIIuohTgF6EkrVxcr
uIw5jJpVmapooBFrAJgc+4euMVw2rUeGM1676ba1YvW2ckmQW7NHzVQVx7A7KA2P
owOClxL9g1kdwAEzCAr4DhzSuuSFf0NQ7IMIu7uZL+KK/M/DUflT+lLtU9/+Yyfw
7P3I+MkLzhlADWBXXKp6Ei/HFQCpyCR5UdqNObZuZeRpaMx1dUXlG3H5e/TSkO6l
4Bj5xNzZYchvA52zmHLabYMVlZydu5xcRdYRy+dO6MpsGK5PynQkusAEFp5nWmhB
Hs1NFYdBE0lDbvQLAr5vkLNPjmhw32F//C2+4vFisbwFN78Fo+oABKKXDVK7cLdz
ALW63aImqn48oBHRDEub2rKRJw7Hq6hhxxNQ5Jli9f+fsaP6xi2FJJR52TE7Q2cb
HW5PBKEXb9mFJWXu/Bs34FzHiT1ozupXtT55TDDX+SNvYMGhzp1RiMiaIxf3NhPY
tDf8SctcoJOoLbtS0taiSn3uTO57CeZxAcInheSIUytRmpdRiBuFlbvS+EHNNw4I
GBjluQcCwhkxtAOHxBDUeBQM7ftDpYuuv3sbtflethsW5Zm/I3KFqUECw9I5vEYk
QXG/ze6ObKRcFbcGeoyi1Tx0zOC1/B6ay67dkM/5sakNRpn6R06zpQQ51K64tpQ8
WsLYKvBohKZgpwK2ulkWmNzg1osDzLK4XZH4Dj+WeRjmB4crYk8Esl+KjPehM/Kb
mseG0Kcqa4WE+CSXyA/n6i7YItbq2sQNYMYC7dSaKp3LzwfxL+jKq2vUBVhRLlLH
xejFxkL4SJBiGuUPJDzxbagSG1x3qxPGoBC6jKfVtTJUtECQWsGLGAqktDQ5Gfpz
wJsETvUnWwrct0MpqKNI9/UKpXgmrgItgUJLHw+Nu7P9gTmD/n4krpuxzw451N9a
ZCiCbRjhFBjCA5iIWd3KNwKcrMT+kPZMkiQftcyfKNnGnUJv2S7vGlTuEsSqrRAR
lvccjqgv4Hg/yVbZyCFDjdb1jJaK4RIW906Kloy6xLE231v/Fsk14778nKVHbL/e
Wfq+GnHwAzkePoAEo+jjwDrWKmfduj+I6ruhDRrtdnONcdhhC/jmwCaMcmV2/2n6
jp3Opkd5nGuv/k6kWGr+h5yKJsc0y70866ZBl9Mi+BQWoz1DJTdcCQJwebXbKTu2
WaTO+N8iHkZjB+IV/fseF1HqiX7p4k07DkmN3J/XJQKm1Y+3+zkkUgVJb2rgpJrx
VhH6K+2kLZt7Uo60qYV+yccggPZLvuot5gnFp2+s8H/9SnZNzqKks85X6Af/XKIB
GXnFd/Lk233U9uzxwnhO83hRp22OwtfKifj6qmmxIWy/7WV6842TULrlWgeY8LHk
nGds2Jipj3IjdAtC+Pne5wMpswsq4DsxKugify+ME8yZcs2qMA9SjfkmKegeIYZd
2uPmVgWNeXl6Mnigut0zHuPHC+4Y9aOlaf7FrhdAZE5Z72FnCovNWeW/VfxwR2vN
StLydZGEyPB8rlAndQkrwLeDWKTDb7Lq6g4AaDnHOMkj2PvqTvpeWLyAUHyIty/y
S6iuLUCWdB+sho+R4n4ABP0grgCBGR1G7LbzwNWI/KTsaSz3Xc7N/FNPvFrvyNQL
N9a8RSb9pW7IvKOQVs2fFbSpdlaJvxJakN/m/q+XtwkqaFn0wC26XspsepgQnH9V
v0x0ZTPCD1EQV7DS4GOLtcn5H2YZMGKj4JtHfOVZgazGKNRGbLLIh8UQBcT6w5TP
D6ibE3GLofiU2tTAOVpPjRz7Vhk0C5zwoy4PfZnvAnPmDdIrJFMNv87/rzp7d53L
Z+ymB7GTIIfiobYjxsE1hyaYXNamf6AMrdgqz0kFjxKGqrVjpNSFkt3usH7vExpa
H8tLzLVgXKkBiUDC0boIt5sttPse90CE5S6QOeHkjAZLuzP578fYxceNC++C15+9
ESLQKJ5joe45iYAhLo/NHofMR/ti2nTgc8nAHhsLVg6wEV6FVRIuZiHzbbZmSTjX
PP0kt/kdbdhCjIexjqaQWERhREX+RaTwsZkTJKIrqDLIKeXpVnSPkqGfEHYxA55J
6cD33QcGc6iXwVQvPYVuRaP3GWWmFNLGwzFu9S41ylxJUR3C4RvB18c+p9sqEtFI
zqlBqlfITXBLQzeAvq86Jo4nhfOaUQPedk5DzeTUbr8FkB1QLHgB7yfIsxeMHWQQ
xs4eyB4YFWkwfHvlzjEAHNvXowwQriybmY4Ink/skZz98DQf1ysCKBIHvCAkXLk2
otYktkNEGpIRtYgbNjI53Mo981Uv5R/UclsBLzjpufNNpA1rMx+LUBAl7H4FNVXC
8WPw0OSeWY4R6gTLPxRJ2cCXuIGcZgf2TF6nLJW7J92/mYUpUT6rJe4XTnXbYjGi
s+rmjhe6HdNFRrm3M0p7Ak0mbY48zEIMs3djkVEcqdxVupanCNH9x3AKxBGnYw75
R0Hf5Ov17PfVc/Y6XAd2U9sVClW7AQfujRmTvs5wME/mZbBfbfSXOj3LGqLYR0jO
s9+M5GYTOdPGctnhOt30bcP+U0IFpb0dNahvEa6u1aLzIFermM2fO4hgClS75U4S
+2V5lllr+qFJwApkppCU3b9QzpHiVX+XSe6iWEzNVQEKP2luPu7g97bp39GEpF8F
yE0ymHlob6MBvo0og3R8/BhEa6dNGV08wwHZ4LX1vCPEKY4oY+tLvVI0Q89iFKmU
AKPNVRB3EpNsDPcjSltXdvjcZ6CG89qMRGdLM/wu4bH3C+bqt2x3YFSxdtJCF0c9
8VLF7xQ5+EP90hZ/2IyMqd8J3kiQPENggKAhVZdlQRCze62lNvyACWaEz/H12Mo4
u8X+lfxLDjTVbc3MPYJgoACZbptt8w0CUNJXOSIZSlouc7MsFdce9D4uV5GURbvB
friZ5+sGr2c7tKfC5Gn8N1oKRfE2tVsJplumuw+1f5d4Lh3C+RWqVu/zPJxA9XTv
+ZUI2Bpyt4mmkrSYZwABJntoznLyQXWGXKbtQYjME88/hcQJljmrCcyHAZoK0+Jw
IdPc94liVwnt7u9CUdO539Q6R3yDv2ovTs1Jg9jYqhPyW1oBPZhzp53ouocszvXM
DnCkH4rnQ23Ptg/BWkCJ1fXrGB8kgLHsG+VyH0gDv1ddMtiBxqF0A8gbAiYPvp25
cpTtfGyyJ5pcnqbewz01nxTkAKASgI9AUGuC4t7FeMh5nmTAgMcoXDizJWFp+dlS
zH2buMWSCBlkWGSvMWUCm5WSV4h1tMV0qnIsnnCFpFB4YViVmcQsdSNgI20KPDSs
HnJp07zQzxj2Bh6IdjAlzSpkfZgdog3LJ3/JGrc9awh3PALM+Wmy4nUJsvfEPbTg
LVcZQ+0/UeSyWfArKzhuYa311qUXk5QaoLWurqTA/h4mXDhkavzrXJS7oxPz3SJm
A8D9dCl/QTG2qVwIiSNkMlHW1yN+zM48P2w8mpTx9sexMVWK6KFewHHoi+XvrXw5
fwUo+sS9RqrcT0FYcY1pK1LJ+583IOQato39vHULso+K0Q/c0kJPqEienRe+QuLh
qG9bMm+p3QddDOxOqR2A4Cl822y6jYBxbQiqcmNmRpZdLrydTjuW5kr3yjl0mqam
HMU0gjNqE248YPPD2M2A8pQ02iWy6l4gGcJb5UkYNn8MnYnMQLbO/5rlnpOXUat/
+GCIyMhkkcZxGnwscVfpH793N/se0FQr7OeTqZrT+xUrZUjw4y8BlvbYz/d0axNf
I12u09vdiAS5d8gAkznGaEJbj17DWw6siTrB0U2EMT3cP4FcxxqXed8AUzodfRvt
5wbVjK3+wtq3cXYIwgQP88lRhoMHGP0ItWl/tCBZyeFQezMcT39kNBHKTlnu4Lee
WgRuEY+utgrlt6Ygq5IQOgOrHoqnemkDJ1HK33/AiCNRBaCeVeE/TjKMyX1GpcvG
MVUW0qfREf2GcFYpotaCmsz8oleeO4Rb4MbKZztsaex3/AuyxXKOSjccSSN+3mdP
Yi2uy/inwb7pbcVtutkL4xONgJf3u1JyF6TAkjgfpBmiBjI3VI8NiVf0GyARJjDC
2YLGwsrgibfpHECtTgQPhgE2anb4ji0NxMTpBM3S0+D0zOOq6nTMRzsRxk75yZrb
+PS4o4dKhyZX9aGE7gx/a6hNXcRFxfVZBKS0zJAYnOOv+yFLmjmfgRdEt930XNus
99i/Z3iuy/9qWq2bbn0xv4wNBGNYzwOPfizeIXkv1Vv5wD0fhiZXhElnLZKReKdq
qyzN++9CWlE6j503YxqqBLP+eJFdwcsMtUqCVE4G9MCHlL20qV4gUV+a9tMNr4Nk
1AN6H/gDLbEXZ8y8C1GAuZ3QM8ml+OmqIGqKCHRCQKbcFz5FNGmiO9HdWFuwmsug
zI3pM1bizpaLzY+uHznIONTN5EHDZwxGNP5NugyotpsixQ+lxcFbSCzkdFkrrjmT
Voo0L2d6HV2ETqVd4UDSszYzlT8YdfPUtKC7gwG5t6CmMR28tgFwxVX5QgzFE9SP
H1UmiptzHvvRsl7/GYcrWAOiKF5UhrS3EYTOfEj1vnKHmEIIHfTL+vaH9SJfTszS
a75dUNqhLSETf49DqIen5AW3m6O3MHczR5IBjJ0TIr16aRI/KZrG1ydZuZJvaAnj
E0r6RRGOY1PpIX02N766Qm76kXpLm0ASqg2a4y60OyiF4esDlhZX/gwaC5K4/SWw
6JV+Xi103iSluHKnrhHcOLsXDeLexQSE0xA3cFdLFTfu51wRjsFlZQvWke/tI5TR
Iv6sqcXo/5sX4LAmFX+zfW1axIZa/ba2G90Fe9Zi7YSFnUuclexfsBygXy39T8jD
APi22N9qDYpwA47wBq5XFvN7gaDvny8QHY2dxSbcHhFX2gYWkKcBGno2/D1f2B9P
yeSNuxxbwNWWEHPo0Dq4ZdkZGQUKVmMFm6rtXXTSfS+HSGGjT/vQQg6RhwO0X97k
anC+MpL0ywvxyi06+yz5KZNbnyQ/cg0dBjq2PFh8vyZ07CGE08HGPYwoGcuvuvLu
1Q9AASPxZ0ClPp+qydoZkV040wjLBvshmVWkCO9aJOaIcDfu7eRRIo9anSHjtfl2
+Z8Jdi/iyJe2zpsIvv7K3228ksnWh1bJo7HKPgCgcvhC6kOB+DBS3FNTBGRit88K
sF5P3rXvm6D7FluIj8ZFLLBUV/wz6e/RDYSroY/gBMANBa2Kj17YMYmLraf9VaJh
/A2UyhMXN+wcJ2g8dTjrG8IXiUf545cIRKjhbbANtMbMlUHPx04pZHT9zpKl6QWD
1aqYLcPuhcvUk9q7+0x2NqvNSW0uZNKI/SQNyHoVpyxOCj7LDyLuHVBgaZeLe8D+
w2BL1Kkrs81WF6unq5C7SdZTSp2K99HbMVE1CZIaiHJ0VvO+0nLNl63FAS0VHdIG
yKm34x8JBVfYkUFIKFMGfctVe00pnPD6Hlmrp4s0eF8OuNzty0WnANLV8IepA69q
8MwLlGpNTz1T3eWo+sGx0a/s71IeZNbVLkFtCvSW+4Iy18ATrA057hHb3lww5BGA
4hWhrtT+crurTGgHTyl+mfd3RBTBR9Ke2wd9joZ5gTWomEj9w+UaYftuSRwf88yM
zLxHM1l9Wtja/BS9+NVRdQ0ZRrrjZA/VpRkJhNkESHVEEMBBYxyaChdLJYzDjZgb
m+Pf7mCvWG6P+rwnQR9n2ZMb6yyxBApMOSRfrAqBCpbJz3EvosFwRpKad2tdT6t4
qNU0V3ZEpdD4YHEZE8nf0cIbfdoa56EsIrfMTChtZIwX+dLzFWs2Aoq3Hay4/Er4
djDP56Zcw6+fTZlNxNW7haF+gfkUKwy4oNpItiPyditR/NiBiyQo6k0WvmGKFeO9
Gx+XdvAUrcina2EL7hR1Z9ZgCwWN9QUvsNayE4j+WWO/bpCXoD7R9ZINMjPIINyN
00JXPwk1gA9CuZhttcbKnSa8Vu9vypDM5uFcPIeGpufhv0nzKPgwxRPyKHZLwQHp
ogffL+rsi35N6/AcKfYoxKkooSVvixf2L0AAan4VHSrNppCHXsl4aqp9yAn+xc+H
4b+x8HpcfJI0aoGiHsbUpjA5I49lkH+pm6gCcCjqwv3GZc9+IohHPEtTs8RxCh5j
pMtONajzHaHKLtw9gM6ekOEpHnkYz6mTOl6CsQWR9I9rTEds4z0wwMHcoMCMdkk3
O09Q+ZNOV2srv/bgwdedQVDPI7GcuHusk0uY2arkAbTZcBLVwiyO1Uie8XbMhLG7
bsvLF7UFpSZJOvqXHtJHtR0Mim43E+ZXIRguH2h/vu7wpFeohVsCW21eyRJkwsJl
vg9M21FLcKyB+jevRbGwRCJw5W+3ZOqfoVRbxgE6FWeQZHrj+T2G+N2VNI52T/41
d3tPxEhHqmvSw39Jon0KXxsTGwynYQfQaaNKiPnT/9cD+jKpN2RS3858I3TPxqBg
8SgAacBF4nAQ86xO05iXuhYt246dbh4v+G7jRMjAqn/bGLQSSYW37fYT5den3PJS
EbHUDA+6TafC9CJu6WGul3XNCVrXjIIiu+Alr7hOI3d0KgquXSs9WT46m+1uqm6V
jXHCN3Gzhb5HpTH6uiPAhEEW2C6+Itj5UTe8thPOgBQx4DW4uIhFPcAllFmsp6cl
hcEFMeFKsma2ySLWc4uyMMKj6MRy9y2mWT7VVg2G8tsWgEfcCOKVKcd3o3HNK8KO
r8dToe0l2WV299l9svWadPqtYzGxTK55z6wguV9eVezXHhLb7pt5ofxJsIPG/BWe
FoGBOcif4C+LiM+vHXNdRICEK5RyZfptOmiB0q2aHrxClwK/R8uqK3KPdUZg1dA+
hEx3WLuDQZ4qQ77y5E1Z7H1LtI06O2AGsr9s+ouqpx84/KaX9+WPkroKIK2JhOZX
s21u1sfT0AV/TMmM6kKIwGekRdUGFriHMkqc4YhWf/1Ki64Ea/VkkRA1jgWSQ93o
ekHM8ZJ0nZsPYIG502GOYGEOwiHU79Ez+NrT0xpvP8AnMYcvoqkxPUJrKLS1U4Rh
W3JmwnnSsUIkXqiPSxYZad4RffiIFU9J4a+kPXhXP2OGNkVdlUoPNPWl4cvGuzLX
aUqkYnZSmlGFKi+JagGM05jSTWC58+ywaa5krPLyKpH3PJfveURekAAD+d+QuxVD
9oGHXRSFnAPTUe89ZQvXAVXlOMU531aPmcoKtz8BNi0D1NjEE8PSolYHdxvc4Z2J
5eLAPgR9WYQGtV7uX9lQ/m/SPrmk+3I8a72nvWQAyBhykVuQC90C9XWhIz8fP36F
8GbFO8fu3uYxXfgZU6+Tq4CqwxCfLaiEe2JstK02byRUj9YVI7/p5xk2UhYBAJ+Z
2lds/3NP4sOJow1m27GvxaX0yzR/h6CPTjhRDG3rfA4jMhbhAUXEoIhaGBEvELSr
dZ7ElSMTJshPeglbvQWzBo/JNckHZ8zWBXw6e5rv0/rkj2rJHahjmfPwVeuPDoxn
mwWbcKwY+HfhLwPSgz8kEmubYuIOlh77/5UQJ1FLaeLb7XEG7+YRgZiI9Xc6d6YN
IZc3LPWM0vgR5/7JQTC9TQ+gga5tDQ4k2iJI69W00pmzbrZwMRl/laA65UIEyJ3T
XJGUgdSQMP4lj5jvmr3LAV/C7HFW3/3wTjyrLxvbP40MxQ/vyv6sDYVlymjBZyPE
ESQL12nMaJ+9suCydPZ5/qJ2rRprc5mO6cNfuAEuMo6/KQjPwPEi+Zx30zZ2MqEI
kFDYgmG/YLl9yvlhLo2pRcGB5cxiQ81+h/qWmDv5JEp4t5qsjReINdkqWkifCFzQ
vqlLzIZn2YeN5l7ZF6Dvq5gkqQD5KLHNPO5lsflCWuBb9vB5CJe8g7JDzAZtqAqP
4+7GFfkJjhbsD4Uum2cjSoF3OylBT8uEyADocPnkyjhikBC09Fy5/Sa3BrUKRjBZ
l4C9p4d6nBxVnlRC6MsNhC7gHlGQvCrjHyjOuALdpqW3b7elrpmps4lWpG/7rmjn
Dq//GaVAbp+nuR7bg0gWl6vp8/za2gcpsTx1CYdmapz1d4/LFG+nH/dHdB9UjCDM
3mDr0unrAPru5y1CZ45aEnedIWGoLH5Ne/9Ziqu9nMufSdDJg7TFu/ZhvCm5VI+n
qqLFkoFoue8u3d8VCTZU06Kv0xjF9kpHyKRAmfOAagQpP8qfytN8699cup2jy2zb
9s3RLW/kk+cv8ZWpM7xO4dYksQnC2zcB1NLQBhb/YknA/CDX2HGC2/U2VnY/XbYL
+75d/XcIDnO+pca8NMDLuK4SYWfp/2QUWEFeDd8i0zdnvjnCTdUpZQx/RQSh0thA
VfndBZtQXuGTQJSxPaBSHTVB/UkjKbcy9TnKfB2sig5Y8kcAdL3qK5Dhjw22Mk7Q
WdNAkNZrfRUhIXsjU4N9rDO3mRAO9Zcku590Sza/WROEeIXs9gxt05XxIg/PhCTW
9fF6omQUz8bCpB+i4yF9q+5sAdAeycxdVuB0LRJNf+cSZ6bko33v09x0CSOvr6NZ
nEoKXi4NCfBynPCaNAiQT9vULvN8A5Ysh/SQsRwIME9EXJw+Rkp8PMtd1CplfMF6
L1df/ft0seF6kz03FDWPx++MRcdZrpmSz7j3PwZBm0EPXk4LderWkKpiEKthCLwG
Vbkngd9//YN82JOvtEyA5uA5xH7f/SniI7qj5E0fGgH2l2ti22wwF7X4xgMpi4rw
9MQgYBn77L1Bu5vS6qKV60hNgG7yqjA/pWN6tI/nqbJjFwmUNCCwY8dx7mB0Mh+c
/ljAdZtF2olpBDZfBYoBGSci7vOiHAiUeHw4gDDjEK8g4I77kZusA4pej2MWnMFg
mA68Jd4c49DImeFNNNzYyZD8GH4Ka4qcZuKVOESoZkWFfv0VG2OYHJ4XI4tOVh/5
jsLcZ353w1UzGWxg4x9gIupkfycYbuNIpCWX4alWlrsm8eMMgFkCUnGD408rApIm
nh3rlNiLH7MRhUa0Skj4ZAzneBK2JQVmidcjHxaiUPhUByttIUuaQBwKrP8thmR5
7MFUzibGP1A2KtBEr1aJvm8yoTdVamAezfWnKzqpeG08AAMQ17q7Gh0WqKo/MvBZ
+iMhgQ2/brYMp89hbgXigeOsVTP/uGa+cDYG6tBaM++zYvJHBTC6QPQ4326tgJxu
WBsEoScXnsbrHyIi34UynBIGJ0SfVy86gI5CH9yUWBzAAfQHE1JdCB4Wm+yj5zsF
Q/Du/FkZHZge0AhLUYtL7pA1Kg4Op/kMi64FKlEcAKJTLv9LEREbcvrGYAEhhEgJ
dboYNyDXZVWnVpsIRO8c2M+u5zpbl7w14BTqYW4E1fjcb7zDc15Z6VnncPW5HP8t
cIRahW90QRirwSzrXbqWnJL0yto1HVKAcpyNGp4pEmPHnNwUCuYtSRFHbBe9IEln
gwrbcf+axu/rO+cFOTuEkO+wN9caE5/v4p0nDnOJE5uMyWuu+OlKxPaQDVzlBOEL
fvIF123toJgU4A1Uxlog+lZbvv3D9QdeVsmwsN73eXLYMvGTLo7jIYSP54+cBotf
za4rCZIsGMjjdpsL98Xmi7XRDnOQn0Nb+GgyJ4S3asYrVkZCQIAserPaKKSwAQSY
OHBfrDu/QX3wPftlYyWmtfB4z3qEudySsMgxRFCwvKBmo54DDs76zFAjml+Yw57l
fD2QXKgiLzwP1FNmgmD32j4e6Hwy3b3zK3H7pcFLVEJlYxcDa7x2QUxi8xOgGDbi
KihbyOhZFBnCZwRbKNOX34Mdces1rKTP8KnH2rE2jnHIEKjrOoWklaMIEOcHJ+tc
EV1+F8XE56J6Mk3UgLSSxhBHTfBg5rdGlJzNDGNVUD2t2mwdWFK1kZCpDS2ck4Yu
FEQ2ag4Tpwt4KCTqIh2Gz9TDtD67eIViXK7TOt7Im82QbH3MSQvR/r/VF3VsIs5b
KyV24c7fn7vnmdEtD6rd/4QY8gxNw00JxgcQwiSq/q+NOs+K5WNpfE1csIT92Ccv
TytnXBU8Lyec3doXZBdR3eljIHDbT4iETZ/1HmGb8UuXY2v0TToA7iLwyF1K0byK
x9n0YL2ZEZtz6r+nTHkoWYc/3+fvc91YmMmNW9j/rUSuTWExIQARjIc5aLS8eXgy
4glqfiODNdgIdFocDwaH3vPKaz3vH51Aq4N2SPe1xbbpQ2IMf2YPkc0s5hvqNPtn
00obEJYFgdzDijI7jd1ehjbXgKz7TYZiHuMFk018QAo/n18NxiQYhN3961mZZ9kP
9eGI0PquHk7VNmY4AVia7SDM9zecpvU6lx4RFIak6ECr2O2TrOhlSNijWxGJjHeI
OeLGOB7T8kVaL2SMmcYp1wsszqrYQONmTLZ3nBZT5blGIeNBojCVAoUg7S5kmqAx
BVmyAUb0gBZEuJb5LNoQ09YW00mYgfadFIOXGxQlFfI1p8a50WR2QDFcEJSd/HFo
CoK6V6dq+ANS/hEYngAdhbsWKmIdiGqsl24hw0BebVo910Eb8NKQQrT6MFJa8TBD
fcyKCgWTzCB4vPrFLE1muN2aR0YfI88t4J5SpjNFik16TwUf8m3yPN9MDZcMqMJY
T7ZpIG3HPMw+5JZfHyAdmDmngdVQjTNYyKPuCqWHyfVaKlwU98h56xjBz71imzhE
Twpd/4ZTjxdh1hX5s3lJxGmTuFAW00EIAkl1R0Cz6Bt0kPORFgV+6KrEVtLOyfnv
839PkZIf6E919/ChswCyXRv7myNhJBa08ImzZ+fjFJB+q2s9dxna5XAAMAHqVX6P
s+h9YLQU5IaZDQrKyqA0Fes1rZdk5fHjwSlP75LAOrY6V36aXJs2a0SIxoiYyyfS
jU5EnGeBvgts8IEgkyL1CRiMDoolR4UIXkUzCcY4EH8jG0zxUlK8vS6BV1pNcWqN
OxDEettsycLe8Fni6NrEjrP3gORNa57dUuCglXHZkGvLyhyD9atlfaWPQOpG6IWW
Z6CfUmYb5H44ojnzV4n0saIaQAh/TuVTu2S7bmVw334cDC4hYC2dalQcPIFx576w
FL9xySWf8AUYluBOWKvP5Tz50cKjANa9yTfE1NP680ZTeo8KPMVROJUHihFxhdpw
ODofKfc64l7Ko5yfwXPVK0zKIRlxvXMkxMtMiFn2TeXOLA3QPcbmwBpYVOfSmS9D
8yfv1GvRQ3/mcwRq1zC1Q6OSv1wJ0UOpi8ZJa9mOJgv+n0gJCPAXakUz1nPqcUQD
4oqpBPWnoG24ekz77qZOwI1plgwhSoD6SphewV93KiCCdJDbqbvh/BlJRJ1QX+k7
jaed4O/RkajmlydhWD5lPPQGr1F7XC06go5oaeVocf8WxfoZEKh/K4lXFa+iqiW4
z36cMYnprajSq82Dbz8VFQC1KA/TzDsI4q30rahjOrBXxXkiCtzdv7FZ037rhuWY
xk5l2kUvkd+dIpoKcxvvrsdzb3ZsDANbL90p/uyhQHDsuo39bkY91cQf62xb2QlM
+r46MLg8PPG2IXUSkleCJiJlkDVcPStcco81VhT3NCRg5/peh3sGqDNSWL39QQlo
lLSQVsiOtlzLd9IkT0BJIfml2qa+8P6aSeA6kk56xDJKJpawY3ymBMWv/T7vV3xz
I5XBsvr8rW2aGGJLkW3R+QjIy5OJj5KzU31Fqoj/HqGUUNHeturUuJo8ClLO2MRH
OyllFo69zAJIS5YuvcKtKqsWgiyA8VeTjjC4EfSRktLgojOhmNHNk0mflt/u93Ki
sE8J/eookd4iwP+RwjuyFm3PbnkdIPZ2i450KasHJ/uJx/lIQkbxT9DkbHe1SCO1
DiRsyKNWBmfiG62GCQJTnXrdlDLbGKOIamuAaVVKXdfEx7PgSe/sIKRIPisZAVmK
IFeiisUBadq7BJUjcxJOuhs4LnUKKy6KXZ3O9IwRcRb1WVM4gcHb0rgPEdNLY60k
FfyqjwZTAJla2cY5y6J0S8OQ+hkSGcJVBNMDCsWvbYtW+fuujN+0qe20phfcbSAO
LC8rZkwbcxLyQVTpxJD4i1zBKQ2NaDOB1EwTIZyA9fp3yCiSWHsxI62LW637avkl
GbXgTjHeVrlKWTO6a3ggjf1AMbbeUsB3rodqXRHNSjHUIH6G5Rh/jlFMRh7Yu+0C
OQVQr66L2fkCCGk6jkJnC0YsO1dDp+3E2zB+bE5u55rbaALV7ZHo2KadoIzm8VQz
VUQBc0ygOXMtvyt76XJSKv0cA8xsHY0MlvAFjZVHVwSAwmXD6fsK8dHwJUA0eyo9
Wuceh7g5LfYhCnclqKti28IrJw1BSlTE34tQ4twqaLhoEkYk82yPZgkvWmmmJNYw
LiFo2pUK2nKrbaY6ANvaZpB/00ib6SQqednm2N4+Iu8FnKomELEnXqNE9DojFOWP
FNFhD/fwSTfEvr11uIfFKdTEeHDGcUfD9M9JkB5MgT2X738p4MM1mfChxg0qZUt0
vmRqaahKYmZWMnw1v2oMOM31YQyL+bmQSmmBN4jmMLnvN6iohDMIeygWdxOvGt0E
Oy/CREG5UaXcP9Qrd7206UMeNOFhlk11hPd6h4wP17n+83MuYmOXdo9iZbhkvL20
YY0CDbzoyKoDMl+9eML17QwBwP6j+uWQPBymEj4x5lqfBuxl6C1cm4tRioqIPwV2
JJS5LsfT6TBKiewgs/HEP4zA0veNdVwoCwTRtIG5JZZPwpWAPess8G1atZXjafqI
hin3k+XZLhKrj26WhRevSC4ftMeuoMd447t/8LoMoTvyEpFsPdi75Jj1Hfjzz6Fb
hViaRhA0aVyFQCqAhyGMUfUmckyPBae/VrEnFN2Xuuu8TfyIXaMLTe87jItz4XFN
dmzB0aqohF/1eexKoRtGrqgcObyVyC5jtusCSippoKstECY+g3PqJzK3sYAtaRlc
oMcpajWYO50X9+g30JizdJChmTfAtVrVvAZQOuNGfhCQCNvC+bcP7p4gE/Uf752f
zoZMH9PWHLsyv+Zlj9W+bCRRv9L79okeC8Oxmn7z8RhMO/SpW2g0qA8EOM0c4R3S
beJlq/Ji5BDe88KmPfZ1pQppF1MyqQ9jADYbl6lhX/JRtwp0Ia2g2fnh7KRNJm+6
GQnWTFDV0nd7KBgvMzDDjUJqGxA4lIwGJUn42KugWna/rlXfYH8Uwik4grOpiN7H
ckN408fsupxgZV8MUoV2XREsqJimBFNt64gjzP/jf0/7RUYIgDmlZp41L+Wgothh
Mh+0G3PsbaYl8nrAW+9En4jaBK6tf9jcmd0Hca7XRGLBzqvfpt4bfkuXrVCH1Vzx
dY54qPR+MK9D/2mu5CXSYuA9aMMrA0FELCN9isBCjjnONvxKHIblqHQjxxrwe8zN
lhkeq/b7RBD8BKyx+nhQYvGbzTuoYpw2/Zwafo94a9cy8eoEQ/IeK06Uv4BfjBnz
qH33yedNLlwPzGGV/jL3g3bKPxZlQjs25tUaiFOS/NfTdsUpHSfHN3UY+7yGzyhM
fCTc1VilLcO3pzAC8m7VF6Oa0DpkyAyk02rey5NfPmcE+Z3wATt4I/3Lv8LI6VVB
aQpD9dEEv6EtW17RSThppuKXgxUAXAqlxLHWD/kknjp5Gy1nHZLpCNQPLDvGgCPq
rExcZShlP+X7mtRoHv6D6JQC/7Fe2HzgN7aQMtsehD0u8Yu0fmbEiVLMzYx6zmsC
PAZafnC9uqZr2qwkUUIy0x63RHGZQqoN++2bLT+SgR2PnDmzvjfAESoVQN81B0YG
3ZWwLqn5XtB2iS59U+ys84ArgzlRMh9cfgVw+zpdfTFW/pHZVfAy/zXZ7xTfq9g2
XsUoCQokTjurj98zbZcHPiP8B6t3waK1C1j1VSlHrFi89DCsduZdLtI3c+DsiStp
oPX8jZ4B306XpuYkiIPzFoo+xcax1GSdBgun476a/OyRdblsVydwqAG8bVspXhcg
v1IbY32c+ty8GxfadjR6/sC0N3bxzYAsD6I6sbaYUz8PNNk5eJ62AwWeQ3+ohN7O
KLPbdkDDyjvZtTWws8RXRjHtFu8TURfqgSfnMPLHoW26ero7y4FTz9HyFALKlTT4
ZHnPtPtgkOQW5XPTQcwTqLbQvcES2IyNL2VMNSMREmEbufcOAeAnSmRxnOMxlmtd
ZVzaDy778+Y/geR+ZIiqJF+NjkK+CBKDJDZQoHMi3fyORIABNrzb6fMextKMCxE0
7mAre6d7a3nOUzZTkRmEtuu2FGeYArvtlIg7ThKUm+ObmXOGUWzcl+IM3fCWddDg
AB4MR+MuVDdVTeYfswUPIwQT2CK36l4zCvYwyYi2APwQYmlZaPr5QbdWuOz4N+Gb
1jHYEp0OM9r0SF4sUboIHUuuCAwSZZX/k61dOe8pXfw0yKraCVY3SFoo3hE55gP0
DpKYc95eHh1FuyoqFwu4O/UgtkFc/boOtlmT+voi/y3rpRjrd3NHhmjnG1EQJvQv
N9f+OG8MIKaVsS0ufWZNfT4wVDv8i664kRtgSwe1UnyPb6+7zB941F+bxWITXNGD
zW4REi7pz5t0p9nt2rHogrPt/2QilVS9ciUodYZwHslYIU8VGWdNI5w6WWyHe2jc
Rb0lYO3rrB+qU/dIphwmW4V6ehz/Hv2dXQGygyNOrXb709d62yI9JtBja+NsC/I0
qPll0jDJ6RhXrU312aUi+RJRU7C0mELNYP40cXWRH2Lr7+f8tjBNXrgATQVsWqOO
JgtbrzxGqe8xOSb0yEMhG5eEzJd2q1xL+tuRulpcmwA2vWfq1GRqyJTK+zqZmApm
Tbw4RuQM6RmfWFQZrDvndE0tewW5CC1f0tr0k6ctCiyqFU5F/TMdmyRC/f9TQXb5
q4ahPUpfieGinJSJrwH9fjktFS/qGH9O5EhdL7UUNLDeBEOG/MxuH22coyFmh1IP
IOpD2kCF+JQrEE+0xUvQUGyOJ3r2G6U+Hf53Qrm2mj3+N3U9fYRuj9wXN72CzVhz
0LiVyr9maxvACaxpDRet079vI2yeed1qWUV2qZsyd8piiaIAASFO8Hb3syf/MiAJ
8qL+yDQGolaJ+QCYlC9X4scU72ODVo98swhXI4Ltmrs3YniXuyYpPLAZOWFr+F8b
VvKNEEj+j3sdyxzZHuCsrzRsPsYLQYI9XgGMIypLLneGAjQOGcDLOveYxbjvYIf1
qrEQFFD/Ekz8vByyQYMGMxz3P6So7Ywer8YweBJNEMfKYwLG9OsiqSUuFY1a7dhG
Z42Q4D4Wd3yNTSqeHVBJIHqNknOgsPC/5j7ygST1U2soP74jA46Qb+KVnc9qQqC/
3M259NLRbCYrscI9ocrBqMrmDEYrc1wqQxe8Mj3+W41T8SS2niUaaZLSLzXUpedV
rVXj38z3cFF7nPvQRbL5c/rltwyo8edtBvBYkRYVF2KgrISvaZwTPHnI1mY8YT/q
FNrw8iBlPLl4sS2hJNkRBUDYC4SK2nFt8nEfICEvfRe+kC2mCEic81doj/j0thbV
hofAvDVGucVDKos6K+0gPf4hndnsVDrRC39mtQUhyq5x3ux2oDzP5on3LxUALiWb
NbWDCDdwzlVQYSWx1TeCoAQwABiUzcr6Wynab4IXFGZmktdTMfwNaMuKtKZsC+w4
mgR+3Yb4AYgwu5STmH1NPuDX+WdZyU0SFaQBYeW2naO/Lxg9z9nJRLvyYdkDDfxR
yfpXAP31N04k4TEySq62vzUvXAAEVk/uxF7JcanHmS731y35famA6NfenCYsq9zv
+FKKjGUhEIDjZOocFmZ48Gayll6W9CNWUkbF934sLTuEFbHljTtadh0pMPDpX8v3
Lf129Q0QdWniZVz3xPmrhWe0WyOfTyFzsji5l1fdjg7aG9NfW04q2eqqCfPEEqRb
6cL6Kdx2a+be62Jeniz0qrx+7moe6eWBzhgcGHY3N4k317UaSnBeY3hGAyXs71cn
Gu/pSk4m+/BAEg3ONp2aEggxJi9kkq++Ls2OwwaAx59wH5z+JBdA88ZGbw9KvrpQ
v8xb5cnBk7FUISUfEw+Z3FNLQTJjc8dB2ap8k/e6ygH94lkX0+d7pb1i3T07JXsJ
3FC7DWTAol0z2MlD3gFdiXvvasl2y5x7Qri9dlGoBmeQABHVfc46HC3/NoH4z78m
LeGRZgYBAs+vf6ERbMgLMNenePPOebzcD08vr2BMaG5ToKGN2CbJBYkDPJZWXu8w
gfWlfsBb2Fggl6MXhHg1rN3fgGHkmSDH/YgOS32CdMpsUn0zeP6D3zqIA2ZY7aiL
aIiwXkoVKdEzjZGTe9wPY594jhUxh7tjBIFm1nfPyjeu4a2ybOkp0lSc7+CdA6sd
n4DrGvW+bj3+sevh5Qr/PwSBrCEWa92qGKcAMU1E+aEYZAB1TAAOT4i7axqA8oqy
tXMnkRxm5PB3sHfRyYJ+pozG2pmNNVzbLpjHaioHPoSyWmQ2VoReUe+GADkm8XdW
ZJMeTu8iJqDlk6vxRjQnYMJnhDYRPc5khJO7bWFW8eqmeF/YP8vX/DuO18Js3IYO
B1J4AgUH/MRUF+sb+vKVKGITFGEB00zNBQJ6WKk1FC5aRoh2hg/WrW42LvSpos8r
xfGOVd1l83vAvO7MB1AfaAOj0mY0lC1b2hPQgVaVlI/5Drcu8sZ9ywURLAfxVizK
FbjEA8DDEwTeL454UHl4lFXVBZq9BCA+7AsBcB3tRkZkpHva2PHJTzHtMsduFQ7o
P8xBdp/7fQSJWOkqmKyKmZMEjO3Diuupjhf/zeaaolBDkFMBKks00Y5zoj0dCcNy
5kseHOmzhbfq+6VYARuhBSpaSyiwft1S+rXenlwWZyexn7xrnrENOqaXC7BTemaj
gXxubCIPSb13FQia7aArPeYkfrhBK/W88znMhwNrPoEeYc4rJtugJEv/SkPhTBao
vjHQ7o/EnHDJel1XAmBUAAqZDgHbj9EW/q9lrD5FBSYQDf8AEHDtgDE/P104DJkE
7U818ecak0XgMdLMY6J3vvVg/5I5tALkE+tEsMOTScZA7jxPxx+GL8J2SqCCYaRL
I9+nNGRlo99GH/hHKUUQdpYXLMI2NNdv3B8s4qu83ZHsmNSg6WMAMYtKxTgf5wTS
n2Y1mQ439JpwngBnmxxZz7Rt6oregSOaqJo5ujsc6XX21b5m1HS/uEivpvP/pIT/
7NF/0Abyi8lObnkC5EEStCL9nbdg6/IH0mL5REWgio95rnurZZbRVZuUxDXjhUWs
qHU25IacyOfj6lj8eL2qL0s+m5JgPdfr5saq1h5H/Zu/xHFTderhJdHEhu8l4/i3
fyyAIuken19uNHuOTqG3hroDQOmA7dJQYPNAGKuxBkOXqt85oytymtnKqH577Y4L
L/ndWPQreiigkHnNM/otA/Y3H8ftlX4O3jd9olEIvRZQCTXy3nTN6cvczyCqYiQ0
yEdQvOJtuJxaLmOAwYmhqlw1GlrwuxM9d569FTJIM/DUfw/YuwmlM+/w+Jox/cM7
xcV8eJ1xSkByPH+ohHP21m7UI10RNQTWHxyanDMc/Bp5AP8j4K3PDdl3yNfW2gHX
q5LhDaBM3TljCHVJk/KVC5q6I4rpYEhwEYfN0QmJwsfZl0PTY+EPfKGDWyiFkLQi
0Rc+X6OlHbQorKPOYv6Dv/hTXzcapBKEfh9/VBypLJskBZf8co8RxLNZk+ZLd43Q
hvTwPxcKHrF+T41teKNYTuNq7ZxxyPP1ONm1xUusXRT9yBqSmnSebrZfgIBGCiKI
mpSilQahvuXT7yP1pxvXuaABzjci13iibRp+hZz2KcTlXGbYfppR/FSTbIysnu0x
y7g53LyAlDAibRLrpvu7tCZwi8LhkvQruEkG4i0K6Esy/cIFiviWyjbG619Rr7xR
YxDqYNAY10LF23unHLoNYO/wR00SM2CuvdbZDTXpz4b+O5bGm4MnYk8Oafw1aknP
eRnkXFQYiGlGfMZx+2L9dN68wbDxOnOvzEHTlcbrLXYJAfkq81QMck32muVJpnzk
+LpE8FteJp2Jel9t81mkAupLbCH1ju1f9YedJtjeEhfAbzlIqTkvUnMQMdMiNHSS
k6X/5qFdDd6+V5evgbwdGlK6Yi3rrg7hmQ+shlqgW4/ZgQTHqTQ/KJA+g1LEef64
GapTUOh6kL0uEVagW4X4ZA125CIbb/MGcPNuNJoDZ9uayZ09rud/9sxZzC4V65F2
nblWPM3sA4oKslAICuLSlW0vt5f8cjdg2fBF1iqwDISFT77xOuNNDSTiojz6FzPF
OGHr9C1/t3U5QXtrqTdqOvRLTCGjVRdGwAwgrfGcA68yB0HNNcEF04Jq20XAHEZO
AXgNN5OToK6gFpI7N0F4cBGdKWLlYz7QCR8Z1QVrNyIg8byvtd2HsOi6vVx65mg6
0pszl9c9fkk8ItHRnFgnT5tThquJcSCeXPL2HhkQCBZ4eypGyDURo9Om1wSOf8Cm
GRm9OBg2RU7s0/dErfxN1pAA3I1Nna1LiZrnR8CoKLQKq77XearH4JGZvQJ2mnt/
qWh4OksOsFhEZHGTJiL8+O7uEkSCPW9m7JvzigOji5bFvzNpeM+BLlp8Y1sd71dD
Bp7qN4tOjjNTJFruHzuAHS5F0In8661WPAasRKN3YFNk31Jyq6GZDa0z/aVjVFR4
dEmgTZO3IodqtjXVz+i7T+GU5TddFSHzbD81YoR6J37KwIEU/0+R2oa7/ypbakEK
PHah3DLiTzsG9O+PNrw/cb0hhtVBBgj0q4jQZjdcT6s6TMATw8b9+VOkdNBcZvXB
lLIajTRjglwx/vMOXeTxyLCoEYWHdO27FnkK/ZRUrmpXQwAW3eQVtfxtOuiwT+O8
hRAMjVhjNTRBUXqJOc9DL3ABoa8yBjpZf75xpxyKGhKJAJAbNYILmlc7FLU3VyTK
BzxOB+gJaI+iQFh7B2boIyzO42AmgThhBNS3RYRZaxS/59JY6S4nHdd1ZqisufpJ
KuVHeuFBjXh66hj9hCzGVnQ9PesWOiWfeQBH8JYki2adxSrne/rTzcqJKlY3yq1E
7GmnTUU6jKw28Ku1YWMtvAPUHVI7EGUjQjOgbn/B28r1SrJVIQUKK2NLCMpotdaF
leHHrCcVzFdA3wKN/jmJDP2cbyD5ksT/vaEA8KjaIJ9fT6XJjgpq6mYl2OY8J+PP
8mdDqjfLvmw4Ql74owuhaLXytpvsVs7vZ1RGjMsbk/xkUhBGACkLT1/MGN0zJ8w1
jfcWNw1BiweCjdfrMH9kEhy7a84jCbEYNZtm8cA2T0nzGz3vSUrvkEGjVbEzJGYl
vOU9yLupVg90oTXBAKlGOYrh3vnGnYb5nurdKBW09l60LqB/lY/09nNuf58Rru/G
ZDlSuhr5tQa16lMX/2E+O77nqS0GPJgPWmikGqjHh3jJbyxm7m10n+guUr6QPxDV
I5g/0Hx+YGz2R6iFnVJlTkjD/SmwGkuSYm/WYSCgt1ErPS49YyshyDssMvvsQni2
Wslh8GOC1HnEnDdImF1+1Eue7BgvXwOKii5w0GBkFG2QBDjo0nN1u1RQ8ElU5fb0
LclhJqLA4KN3hVLYL78qUm3FToHZkGtSB+l7r7M0sidx3mss9joKyw7edLj2Yjil
XBUU5YbDMZ7AdPxBcF3hQkZZPHbzRuPmvrAySJ6ioXX9eILb4YyZBOV1DbSTs12p
aGlICpo2qo10BAySKjyZBIRLFDfT5Up0N5UlhmsPyp+0jGezTDN/pPDsh8u71vEc
SGtalKKQz+wR3Sxt48FqCDwldVORP7jn6wGcoEZmer7W7Su0+PIZSgVbbqAObKDT
bSs6l50dLZxclAceeT254cPxCAd/X9WqOnlZyBcSTRA736qfHYtL5HS81a1A37wX
u4BmU4PDuchfMjC68E669YByTllRMDPi45Vv1e+98gR//AqzCYHRHTc4ozIc96cu
kcPwFElztK65c8XVCjZBqwNE28MLRq65UUBgMgujNjDZo8VxphEFZK0vYb4mhP/v
LNplFNzUy+UveTonUfxNbTJBP/DPsWbyYaOJ1wC2N7oqnJb78q+zSkEjPgWpXYuh
2Q9BMAmnpr+/tGxDh941QpdCdQfsRC1CwUGqcXxtW+Io58KG43wRIY+MduA9smvh
N29ccsbeC1l0dTrdgodFbtXBHd18vZ1Gvh2ElvYUd+kQHMZDX9uPc9GMu/UVgBk4
0a+deRM4RnoygfsWhFPsR1pK24GE7qY8+Zd67d38Ax1sbX77e2cKrGGS7Sq0PbXF
HFs3xjqDHGEqcDslK4oJ6iFTkl9cV59qc+cHFPsJSGmRFx+se8cRm3M6GVwhq4aF
th7lxqXQGKn1x0InKmLfx+QvGwD41mgwIWLzyzu/fPEVzw4tESY+Kr7j8UMlWC/D
/reihNg0oo+xSnQk/CcBKlg/VaDOQbcx1bYYj1adg1tczUMMwJVTTFTfh95mst9+
KCGreo/7P4yRbSQmNY3xj235KpqRGUbwdS9nhD1i4nyUnvqkBi0GBZSmw32xIF3h
I1jWyTV2AcNXt2hDnqh0P/qQiQUfMx6YjPf7425MqGaPk+28cTEx7OBC1nhSdpwA
XtztRF0cLdhVq5ncsXD/CJRSa0KevzyqD4S1Q7OxgHPZrlaOr8rXWZtPx1D/rZdM
i/lEfb7WzqwAXNImR6AWR+40aPa3IRYKwWMsHDCV6bLXBU97eOnrNi7bJfjkrhhD
RQf/U+6T8guXkTgl+yCpqazGby0fqUgZJZVD51T1X3pwZsFuOoK3+kIoYrfPzF8B
bfWI1deJcrRsaoR2EWTD69kDVqCz2hoaiNsXlXW6+FoOXI/m8ySM9Pzfo+eJp/Cp
3kZkybmDiAjCgeIBXSR/e0KHYmUGdQvLTR8BCDGZT5052DM2gqc1DUWJZVuCWK2M
mm0t9zoZQqtI3YSfPmgQx7e8yyFw6ip7Pgg136kr97eihipmcbaFTYTZHxV37lf/
iJJTd1fHOnQHFchtT0SZ4IgLQfMkgtlvCY0yAQpkh3PFx8zg686+Rph4UYTAcnC/
cX9Wmtphlb9kBAw924q6fy4F63jf35tX/cgwT/1Q0E6Pvb+tcB/wSsSSkstiXk8R
IvHl1tqtUeGqYNw69U3RpEZ1XT4ALFKRHQbKjMEv6z53k6ffaYrUXwXznknGZKgh
jHi6pLIS5OJIy0KvmjbUyYS8h5wk82H4ya7mdo/wTEV2j7n13mE9NMdJgFJjtPnu
2Ritp2IRw0OxZsAcSRe2yJ8I5DYQmYt1p5Ks2Q4kcdub3WpjHeXVqGMZ9GTx8NnE
RnRQz1x7itCA6Iqhl9GW+ghyXaQLr6g2NgPca/KxvV8SvKHbtyjHy+WmmVZQGePK
eySekO/z0N+HG3sRny7VoDx3Z4xhASMseSX7ZEIUatShubZOSr/90pnhw0pg95AA
ib7vBnT5+wv3Hjw22cCSmS0+6b4hwshZdF95xUKTgQCzmPIZxtEVq15NVeiFWcep
RVDIzR9QcQNu1UCXUB6Fg+Y6GOveEJWFu0PaVxCbmLhRcwh3VPAUOVqFheN80CTY
Yk2bCyQ6wNTlactjH5+hr+Pjk7Td1j2WlVGZZPz5RFi5Z+GgIwP467iYfGkFx2Pz
vqXCDXOZWLiijgRsBb7+dJNawyNrZRiRWuL/scbu/c+oY8TRH7Tq6qNt42MyuDRZ
XzWAJtGqGKvC9jDB6MGeYyycsrQhjSn8Wkw6GLXjO34Oi6sL5g+4GYrCbaDPBjB0
FtpAYVFDucZ7oI2CHHZZYUOmej2zKR1YhMMUeCrF0i4nGERaqfbUXHObkxEoT9eG
BQ40YF5vIu6p0qxeKsBymnEnrOCNHXbib4mDKujj1LJWg+hiCUt73HzXu40cjDZb
WiijU70NJen9abf1Kf83tV/WCxbzlpnBsSGLCPkAy7wwBEGHe4pevL+y+MRAzB8P
zOwJLQJf9tnWTjSFRrLG1ZqMjAY2ee2WLvOG6+uVYq6unaieoDCLWVUfaYviuiZU
ZOK/4rcmTTr9+MXUJ+sl2AKMmCOAQCj4Z4Ba61Qo2YgyZ92KQGjNwR/bZI+ddZbs
ZdMzDrYF8T9mBQc9p9jCtS5x4OOKYuhst2/1Np6y9rOXWgEBLkaa1fdzOW0ZX0l8
QWlaIv7rygRnZ84Eqd8TC5mMzqcDY7mZiEBGRExX24YKKNao27ckLxGqonbb96lR
gB6TrDG4sWQZXXwkRoQiOsUT9gB04vfAfFf1ryBOnEd7ppNFV4PJ2W3/tLQhC65z
adzHWAXCUKFrf8dPBosLkKlB+Hm8gR1HYnLCjgRJLSBwz7RWHxm2wPnHVZd6W8Oh
H3KQG9Osp84orEJsOvYXTeMNgaM5VOq+VO0B88G67ZPRUsmyHMhe9zGbLPFy9HwP
15cbZNvsnRx6Fy6XYvFCxq4uz6FrJ2G8BrTaGi23sihvHWKttBj3QinhGKYyAUo6
Prict05kCiLnEaIeTyj/sOKbiZlwnwU3Dd6K81apK9tMfwH5g9xN+Qbr6OL5Sy2I
NZRJi5sch91BfzIJTy237HFyg9zM9Ux3y68+3spBuGCkY5VJDciCsvB6SK/V9AgK
M2EmDB+JNjwf3MeeDvPpVlm6mMxW3X1VcstE9uuJzDO5bAThUfcDMDycLNh9fc8e
hYAMRKNTNWKLcvkVg3NDF+zGIS6AF7RqxyKZmUwVtpi2YibFt8QLLR5t0IYpruWb
RcQcfUx7H2YtVvEU/ZrD0T4wWhdSsNe9JB+JtQp+jbV6X851XZkVNHNw02F0Gh1b
nGqn4WMOFbYoZlRJaW5UXXZKUTZz/1Baw4rIb7FYZiu6Ocpz9usE3K8fvQLk+2/I
cV8LB0trFqCveMdg+k/VO9ez0I1W5qqUDz3yYOIlCdbeZYgQZV9XKydFVMo4kXX0
OGk1XGbvZQneonb85TbFFLbNP2uN/Kf9fj1GLfbQbOTdEpNdekZ6DUr2Xksm/lhk
RlS3jqiX1F19VJ1V7JGF5WXV5A3W7iVcx1nDe4/4VlH0XfFFYPIkuItBNstHCcoz
Z854Q3O/yugjCTDgG0x2FISBqFBiOEshJYxDW4w4jek5A8hMU7aQZIO0BW/pgXqD
sG8QXctw/W9QkjM+5PF5DRhxwwNl8T+OrFMz/L4mkVtGeMXQ5wj9oCXRgkTblXNU
GatW64rxW7AN7QZZJZBbdZYvfV6Umzn7YYbEnOesBbOxs14C/Z5Hyduepq9N3mCe
ONrkMfT+1BgXZx8NkpRn5MuN6wN4+rj3XHwLsyAZN/36qJYp9qWQ2el/cigVJxcR
cdra5pGxz88g64eOOSSOmAv5Q5ge/eSrUS+1+yHOdlDKJZYpslQFbFDP2RnyFEXi
6JxBpDX+sxSFijcM93GHrRgP5U//4bXWZvf1tF+hlFZEjOzuiVVcEQX0Nfhy3SYr
OasGg1ijJ3aF1r+ddGpJw4C1lNujbqBsdDZorjVHFSw05MfWQjbfzrHS0wm5H9tc
wtYkdOsD64DhS9jWjlhm5DUn9ShysmIUX2eiTD3+2JvAk7q3ECSkaGejNEPR2410
5/l7DYXHlD/mpf+bOTvTXQK/yJ/IQ/U4ZzDx8StTW8ZoJMcL7atXqcTBn+SMz4O4
c6U58NTgFQoL1VtKVJX4bOg390wPnCK+bZT9Ry5lEG4u+gua2efiJjeKCqyxUOym
yS3TKQjtTwPAoKvtZ5OTMuK106tZo8fx7dN3aBSvQxtzRYJgi9ugA8O4C4Batj8A
GcmAIW0OkH2tmjxaBKoW+9RJ0xreYUHqHKHHPLKUY6HrjITQUGT/kTMyHnVkhgjx
P2+hfFjfZY0dV0g5GaTSunh9ibH0i+ZgTWXyc6JBb1CuB165GJQWzpClhIh67WXZ
5Gm8yb+HYScewSF15OUaO5LVwYZVm0hWq3swJU4GVoWdImLhkRs3XvS3/sQwerzn
oz09kkcTlBtwT3i8W9DLvi1CIN7Svj4u2BeJJLKXIeojyYIjym8+kKfbEnxlLo1l
/EgEB5KjACDsebYNQx+SMwqN6bujhA08ywkXXtxWDmeSsvyh5zgoQ91zvSBdg0xV
X8KCxw3Gj2FWJyATt01L4HQCxv6ghiSskhwp0R+FGFEE377Z1BFMwBOEepfWivdB
DqC4+oFbXtCdDhdES5JTszmdNZ8533mEX+0x1A9hJb8LOpIViPbW/tsKWepWFY9K
FXrPMPdkZ67421uWO56zpGL7cOMymumJP0SoH9NeKkNZkOgAVBen+Q9AXw83jW6N
6/lL8Vn4+5QI/kn3xZti4S51Y2426WWqQV4gtflTrZ+DYmf+VZWG4CaGlBQwU3h9
gFpZc+KajAj9fRnPpqfFmaywRrEQe616j5GIWFTEAt2EzF46i6wdy6pLmMLf6VeQ
MzoC9R5ZTd7W8gY2Dn9Sj9pCsfYXIRLsDCOPXRGfg0Hmv+7m7maviS65Ig2qhVRn
5nnftmGggndh2Be63aHiBk6vXKt4zf6gm/VxyvQhdeGHYkq3+XV2CC/s99UOdw6g
giNpDcag7uldrtosDm2TyVwMXwPVoB+mzWHVw6wqTihZIXt63/8O2c3OeOThwxUH
AMO6G+IxOYp6qBevOkBwxUOMn8x7xu6h//C5RD6zVvjS3Vs++HINq6bKm6nvTYHF
+mek4FRB70EJt2IKR2uwCQ54FnvdXlNuUYB5x1BQ84263mqwka9PUYia/9Wy5jas
NsvDZcbGhFsHDaPgqrzj33m91/tp/XfTY8nK3ea5KZlQR3WnkiQV8v4vXsp9QWyq
dsLh7QARBop3Rx8hxvISQK0VNNxRszm50k5hxfSt+f/f/FRySclrhP+M8Wqo+bWd
wwU6582SqTZjozs2PGl8j1sAN86u3jlk6pPe3feVbmYkyjcdlFJO9YB+zkEk5kAt
SoQJsnDmFQZ6eIbEJJqJUIkrNmJf9mI5UMFMdWsrNUd4mwQ4UGB4dl3VdXjaemq7
uy79gV9WGEfFNAoVndW56lUm/hFSg1Q+Fo7DZomCTGFgc4Oke/M9iWGKp6cCPuh+
jx4Os2DeMLM6rxANs1MA39idNfINhX1hk/ibGXpgZAXfc3cXzHup2dizC/5ITeUD
sxkOqRn5aeTl2Y5qeKf6gHIYG0ritflEuiPnzaOULYkiUsILl/9Ntd2uS45Z0b50
3/aD1y0Fu2MWvBM4sAjLwEnOeDpfokfs9N/EYd6wWkLHvy8ms1tJVCYKORAejWtT
vv3rJ6BYJ6RBQG19RtQCg+w4mtmoxMP0rmDw5DHw4PcBLlsaW0bLiavmES8NfX9e
WHi2+KT+mnwDyfMf/ZMSblBsIeLYu8fSDIZlhNFWG2KiLGKfifJNyEDIqKjN5amO
4GRo/sW09RNT/n28q+QxkEq/7TIHSEiBoZ5rRXGLpiDu/7MpgdRDoPkWOIfARdfS
OGOG9dYt2YGOsh3l0z+LKMs8719YLnNSs0mmVt0vowq4rDi7AYfggg0PgAYTjOf/
Y2kPZw3xbroW6zwkf+vbor+ZJEMLrUj8OYvBa4FLbJ32FlbmhiY4K0bIVRO03iQq
lKijdbvjYCh30ofE777pikGxkI9gTUyBWJoZBWxOIaujvcWGzT+O0s709jrxcUie
Is8Bw1piicV6+CqMVSpcI73NZRNjgjZGfRpR72/ecOfvkm9OEu0kSyH60LEB189o
9zJApuKljKYrva3wNn0JYlcC3e24snciRFcFoW1qvhFaT/30yDg+snpVapDHaY4g
M0sulkVF5WAEEdsf/anOp4c5zr5hMEXLMRnkCNXv6C1d0RNmRmaTacC/X6ohdT6m
TNTnXrgzAv9RpT7irWb+xeTrhpOX7SrOQQmdWTULlITczjwsOj1f4n9sCW2Juyh2
JEMRkcGPot2Wh/uMW0+aU44GZHG0IpP4F+rcB1DhNH/q3IpgF3lxSZ9Wt3fnKCs4
obmKGaagl3caF8wrFMRALIE+qC53ofYj3BrZ68BmrDkvuq8XVLSFdjZTw2cA7iph
P80UDbXFb6KYqCzv9pIF3FFL/nY7YGK0Zsjhh64OVPqtiqProKfwwC0XhUHWtlGz
gRGodYwmuP7hcUeLAJUv3su8na9Eb5POv9f6sZbFj3VHUKT0Vi8TwVLAJ53MO2/A
+qUousb7hlT9vNbb/2JFUXxFDnInSL95Iie8LhbYHlRdnCRnUfx5ErSvOYLcY5U9
dsd7uPXQCy47psiR10pNcl+4ekLKI5oGpq/8Zky3ULj02u7xrkvP/5vJWmW5Zpbt
sNKr+i50R9N886ayIXJVkpoCkSjTmMfpq33FPY/gAwfMoCRBwHwLbYooA1bxh9nA
4jmNwsEtt6gZfB99edRfCGR4/m+jWUVAcffPFShZgTR25VdpKy1CNfPK+hAR1kop
pmEfQFFRobFc5Mj5w9raBZ+Qy+95O8nd7cpSg58IIQHkkvvvhHHFp2eyB7/vofTU
jw/ku+b7tigLBgzBM3UNhkKyiqbIDFyfUwM/fmiy3ZbWPu799+MmSTcRPEUe6JxK
PgjheR/wSo8wzSkgTLDFjaA3fMlhSUsBQqLXtXv+eeZqZOnxTnsyH0Zwgfcs6LJw
ojOc/Juci/WKrhytPAxuo+bWmFnr6DzjgyZTPMpgiOpa7sTNOaDyI58Nz2yyEnx3
erD+vAdvuPfznmzT0fj4D1pY5YDYMAazar+YADFyOkA5YD+GMqWOeXVc34lrSDOP
fq0uhbFccMB4aPZl/parAM+CM24heKB0MPca+a8CZD+u/fZonuM+7juiuHuiv6l3
qNGnOetl0l3/ihJI+VwZD3A7YQIRlMnCdEMqotvlbvAUkOwgLpslrH0xcSpRVbsG
gqE8sd8Xk+x1UTYkz1oW+HBHCORh+d8FLyBp/9+j7cPi8tnQqCGBnMiH9pBGgtV3
dy1piPPPYU4Q2hfwOncf29JoL8t+tlz9sWClQS4yaaXLI29p8dmikxadr8slNu7L
JPxB2RuS2pUPkPKpvvmDSjxLdjatGED2yrm8lDBoPnifPblDJkl+fXG+X5JbyHml
obwrYcNyrl65cBXtXhZBrEK/6348PS3ULnOyxSoG+9PUJYd3bT6VK+um+Cewl69W
QEkibAaWP8EewalQ+Gto4Q4Ev/lPqlBHzeklb2Dm2zXux+sbG/us+qXpPIKP2RcH
1ztaKPFhwNxek4lliTDtkm/zr9PeZ2HCiU1NaqXZDlv0afG7GoJ9dpAVNp57S1cx
Dh1GgA5PYPllZFWqUqUljZcgm7aDTPE9LQ+XsEVd0qfiM1eO3elaI6q4LfrTAF4r
FDG3y2N9ZEVY4LQ+rytTgeIyaq+3xZ3oSpRkuLAa4IrcTLJqbHmRLzTClIXYwyNs
OVI2vCySjt1kp4dnz/OS3mcEDjwzJ3WeelUiyajZUnzl6yjU9FRNkFhXB6JwXqgr
EF7vSLydweVnXieFkOgM5LKm8vHt5dI5KnJGzEruKZsZrv3Pln+TmT/jrVWQCugz
NZDElAYbr5lH5rzxCxgk+cgHjtHRAEP/2+yBXT/S+c1v1hv+C5OQAB3B1dtukAZj
lmparJDU3QqEZyNQaaNuIV6hg0l4Ojb6VDVEPQELj/zt+7xMFhVZPYW9dQ2YfAZ7
ju8+AGyerhsrB7qlJG6blP5FuimH5b3uljbEZwr/TATXYqvz+mTcA/pliv5tWs01
4HeMhYRE0YfLNRviUw6/XeppeGGQSGlFWNU1FfnbkSbDIqPmqEJ9BkLLMrqNKtIB
MDM45ZngqfFb+HvKrS8n1x5fRfj+14+rsFlrvB1DkdjK6sswbD4QVKBHTMVyVhpM
EDJ2G7mEZI+NsAxpSc6SDjnBwsK2QPbRw63rLwfh/irUZfaBoxDigNBsOtdx+MWF
cbd+AF55tjirani8p/nY53ZFqvMv/h1+UhbDiBU8XYzp1c9VP1vEfc8oFpptN5Rc
BKelqHzfBg15WNh9DL20c6/s7LhkGWZZRUMalcVFsE108vvFdlQIgkvY4hnsn07l
mF3GmtbQVpIDFfpU/VBFCH7LJ2P2Xm8sarPfKGyfMv+7SxDzyS07vXr48OxM9dpn
NAcJ2/jaSClI6DkcNZxVw8dXgH+kLmUH637XsUblzMHLpWOD1Y5SBEW6Pq57DlEC
kPJSW3oQI3nDMwVjaA6ggHN8uqEjr0NVOshgVZganWXaH9S8JVe0Ni3ffISn1qEs
AQFirWfXGaLcyI1xg/IGEhq7kAhWV4K4hUZf2i0cGfjdJ14BtCxHP4Z4n25Pcbck
6+BQ4i/AZpYTlo/9yEZC+VXFQZbu+K+ZOfZMzoyWE8fghR3v7ELwCtL2dGQggERm
HEGRMZtw/DhqHT4TfV8hdQGVloIYkVQojHr0+G+Axl6mcDUfRJmO7xfqTU3ai1aj
LeV585ytGhqasX6lhzr8SEg0mnjiIe8tKhUxf3/J/5zJIwiOY3k33tpU71SAyt9f
XIaUc1QgL/bB1KirSJd8/40tSyi1D8PLTRxyVbrFW15+jScaRWpufT4xbm1viH8b
2BvN+z6/4K5NwnLpeHKKPyAvGlK2mokGxEzeeeRWL8ui5Tc6KnfBUIL8ODTO/0dd
j8L0xoP6CK3V0dG2Pcs5rP5SqjXBkrDf4YIDpu43GlLpwt7mgN20+S+m4bx0jPKD
Kl53O86cln1royjRHeVZr/xS22uEFI2WwzChWtnh581Zmmpc8MeJjMiMSuOZ66Oy
VjzMiHGnwTOFfRKe9YDzXM9zJk4sbZdY8IxTgSJfQHXmxrKhN1c3VPIBuAMAMk7S
5UwZSC6XlooY2Xf0y73nAhHtVjOxNKyXz+WYtQb7/jhTMCCBHs9L+Q/NBvxRSkE9
khkdx4HJQ1fk76MThi7CijdaQT4yeCgC6ntJDfuPaK52XUX5dxyVeflOE/Xuf0ML
sXNaDC2IL26rDup1KujwwflLLMd+Almf4lnvYLmgAeu0Jj9iWCBIg4N4fuegdMcH
cyKnw8FbxDcQXJZuN2RQyDgD2Uo+bfiFzzMFFi/DdNHzmA/OHK0ENhpVAZ69gWH4
WX75p19egbjBNuQX3olPTDwdteFBuio1Sabr18QEMe+EO441++Me94waPhn8QM+2
c8CzeWRjyYiO/CnRnvRV1rllTyS9aocqJIhkwC7KYmGLyqWip7nWcgl8GGFQSV+k
uOFWXrzlTW8G/b4Ff7u2crqxzXokSG1S5qDJTGIJ8as4J4ux+eLdVivuQ2OmKoAs
faiAK1QZSa2ghehBpqY2lIG8vRytmnUsPI3g+XR4y9t39dr8MECCE0AqGlZceH0M
LWoVUd8syvmlazGfjJwDHnecN2WT+Z9gSLq0rHVCWVOZ17ktDVAzsbFNiClXfx4/
a6XNwhhP8TQ2JDkljUoLMrV8gcuaO3rkLLPBSpUqSznAdjuzNQOsBT5Svj9CjvTH
E3PZaBsit7MS+dSsE1UfC8c79tWF2lB/PQnQA93igc/Jd6g+3qQCfZrJ4/pXj2lh
P3XZlCoPQ/SdsjZ1SRzaa5/CksnGLhSANRLu0TE+cX12gpBGeIomuBnAuN/x+Niv
7D5bCfXbPVOJwxNpNih1EMYQtsb7GlAz3EGLQaZjmPyep/pxCstlOTxtqcu0CuCX
OSBnStAhdD25o5BXxwT7T4d2Ez8pFn5boefoiLp4Y83AZCllph+ihqNaudowpmM0
WhQWkZyQXppGCFYVGlzClNaXk4Pkg0HokjUUZH8AvR2djF+vbNnBhzo6GQ5v6EbA
TbxWKQ0LzCcrrZ8OWO0UoIQqZrpg1KF+Q6YyO5cBBq37a9+gDGfnmX0016T6bil7
vHL8Tm7D/faqaGcLsc9P1J/CVWcJRQlagJGQs3AWTvFHAZBnplMaPwVqrUqr9LPB
Hb/8dei8rORQUqq2EKmXb3JPPXbYhXKfYhYggTEW5sHB9DIqTS/PWDJN0Oy7CEwK
RRo7PpUUcF9xeLy68wX37/20Bw2yCQNLTX947fKQX7wqbiCX+ro8JIYxC2P4nUg5
SRau9WWtazeOcov5N7Jz/gBomw9VAhhPSeKRirsWHMrFXYQpPBXvN+OsWDYpSI6h
t0RWocOqwUAxxC3X4gThFoUTKOIOiTtDYCa/025rG3Jv19t2Y5ahnjipEmJA8bIa
WubUN1YevpziuXKcAn29vgi/Nf+ON9d4EVaPIPNYXx+3GpQJMWat+KVu/wTHxmkR
sy5sztI0wvSMb/TVpHoSpExtCZEVHUnZpmNoL0T2lzK/mVuB9frW3JijYjX7bioM
MGdvcfO3TsuNWwOR6tUim0ImjsHpsvxgK5iHMM8XMe6VuGicTS5J5ZcrHfMN607o
n8PgY4DDs9xQynJQJd+HWzy7qELWcANu6IOXLCoRJ7pw7/uRI6AMXiYzcirs2spH
MMjJcvMDVlLnZJKBoD08lClmPFpJGAbEYoe5zDlzkbz8pnK0T9qXZo9APNek/12q
tHm0eyuxFeC+ADnKqlBVzCxWq+R8dzfE3Jq/v3AJhNIbn1GgETAJICU8Bt6ED6uw
DD/lWVHd7BdpgA/HQ5vFAYZuNijlOx4zHQwZ39wwV3pBf15kR13857Y+QbrLex11
TSNsmTFJliElfYEtlVR29v5LfL02OWA0EA/KaCTUHFIlwqg7VxmIquslqKHB0ebp
B++Uvn2iJ8YGVRM2M5gvf4EVflCBEiDzWO06qox9OboCG0iHzBUH2vNK61GuodTh
2YpZc+kubxvMcyrcBtMQETTGSpNqMZpZZK3HLN5E01wBWfZRcdGs5nqNr8EljFi/
/kvTjPArM5f2I7w+dKr1GIxio91KDM01R/u7OQ2Vqea0AHMOp3DvsIQv0helfIOY
UvunJyY678VyUjrM0u6d/7/Z1z0gzy5qIowaBZIGr6/EpDGOn30L0cXTJM0p2/UC
zJ3FCZYDJZnrBmeT9BMQIxakC3v/Z6cHsirCg+Xxmpzfdt6+GcqEG38wkxJ93eeA
+63j+NkFtFTWzfRvgeymVN09DXf0k6/DdOkarqZ9fIZ9rLyvglMqz2YlaUE1gJFi
/9Q3evP3JK9yL256UmB0E/easWrKWe98nO02ClrvtQnIAwYN0CJjrexS9/cG0CG9
CK8qBZzyxvti838pnaQha1NKMkjaXiW2siuu9jU7jSDiJDyHzkt3plo3/yRdDyjR
G65g0yDqMBfowlI1oTtSl5ojeHG2v4deDUnaR+xc/0Vu57g98AxSZcwbLptYPtil
b0g3D5fgpvQ67TrHw7K/+OXxiEtToICB0Xyh37g0qE7ljyfd4ZTNlLg75reWh3kN
kAHl6z9Jz2eVfWv9AdkMo7+3fcva4Lzt1MmEbsL4AzAvbS/2doRqb3bVwf5Zwvkl
vKQERSg59F043wGPVxI0b6cUQD1uWEyyOvvrxOLz5o6zrxUI6Q5BBLQEJk0iOGAU
mmyYZLnPGfp8iOHM5hzzuOFZE999G4xVJAnF1llqcqoWf7n/RYtG5YVlqz4dhGWT
8SNSmCzrLsaCSDuwC4CD5EpEt1fcysBN7UpOSD0ztFqyrb3pUkMLAI/W864iOvY/
VIVn7GonfVyXni4fpg5IMBVo8JuKlTxfjg/UIYv1y882yBS176CAANDRRFNkw5xC
/By3shm1CsjR/aEICysJN22LC4GODkKp4hDv/kLSt3VpCzTEKDmGYEfdlXXe++PA
jjBqJq4JBTkahEigtHNMk9O+LUqhrMptuIu4ivFNcUJvJ++/qmqEESaS8GY6anr8
NSKvGqwTha6cUWbh44ogG95GuhO2B7a9Yz0Gyw8dyTmH0ZfR6srwh2ktXLLHdVZk
Lhplw1yKSS2H6jdAd9onurWxjfkhaOTrfPQvRlmoihI7REWXoEU8mnZ/OuHu80IX
a1iCMsBCnNyCHTOHH0HTrD232MeDsQfMvuwZJ8m5NhPXVKhtHDq5oxt7rJjh+zkn
WSej7uWlruMECxQmrqqMip0ttvgX8xONw0de9QzgqkediQHFzbYxON9C6UdszmRK
Wx24nLTylHDnig8kD16APRW1nTBhkV4gyAxwXm/Nkg8mjUZpoC83oer6G3k3Cohy
Cl3vKPVeW3OeCUIMH9aKyWQMj9h7oEY82WbA0DP5QEI2yDZ1n8Rv1SEuf1CfdRNn
I9eZUczSWUPEYhiaaMoSAaqrE78sH4p9QFjaLKDvrxIv7dp/0+12C+oJZLOAPo0v
R6xOHjQceyyk75f05seGnEWex21bXwpJKkS5L64Zk+bf3D5pih34rTGrZBYFn2+P
SvWlEkCIuQV7NlCvkfMPlN509JNtketk9Ov1YV9BQlbALLliU48TKvR8CUGROHHP
x/n5UM1wyTJVK5VYQF8NiQVDeuV9bHQUl+e0Ltx9bWI3wE2vnm4/GY45ZmWTzy0+
nxrwCXHY4B//0RGrCMCKqL3F93YrNbBhDqAMZBjTRjYlcvkZrJn1+y9qICj8/gGp
+CoyAnezEc30bZFZ0rg4s1YjNdQm3JMgjQcoD/6XL9q9CGGpPI9A4mv6LEoG1YU0
kQMFc+BNP7vMpY3gg2GoSPOVY0zm1xD3MlNVAcvZgoQwaVG0cKAe8oF9qOxwpAPB
E0Uku35ziYSezjKCMEA1P3/cqLCPyYLpK8Wg16i6jDn9F+WjGK5Mh5Wvcn+uUjsu
3Yzl5+V9fA+qb/d6VpzguBN0rCUGlnKwVAbGLXWJUA5Uwq73v/08/aLGSo+Ogi/M
D+Y8tCW4l2vqbGtldZYLSaR1N7gxfgJ4oe+0gm+Wk5Sixzz8zzjQO4I5mFhT3LQD
mWuWvHnHOTR13dfw73TqYzucI9kUKNjSK/AV5ByPPZY2TlbkTcm8E9uxVbrL5CM0
CqAaObHit6Xx/Xc/11TjyHvIHigPbp5koLZFwqNmjz8Avldemkb59dSPjxmcEdhN
NJ6Wjof22w+Jr4VH2ibSb7eUsMdoK6cIwmWDZecbcc0JKzkJOQb4Dg5PcrbKzK54
pK77MPXExsFrk++MnXt+1WS4EN4O1IF6b2nSlozt5qSLUVsptT+4IYVsl+bkPvQA
AZkkPSINis3cU9GZ6vsN9j0Er8n3cZL9Dir8a4EI6USTfV2JVe05WbkRwX6PGFGz
p4+tgThNGSTG8hTy5iNFwxTZEaPqw8vbSkoMI1f2BiqZ7g2yYdauXQm8J84QP8H4
2ucVDVxIzNb6+6hwlK0/vTFvRxGuAhB042zxWjYtgoagCxrgNFTZfyRJNZZVZYoT
4UpcpqeRIgotCrjulkJcYkFgGaOCn18NJhBM/0T3VojB+Ta95u5/GFVg1WvIylAH
ubxb16V11hAxxPOgmJgOJ0/t7b0X5iUbVO6PEwXrFKU00KpLhAFeior/OQWTabak
WyPuA7oT39qDhw9QnhrprysG8Ilk0vK08SmCpQNf4wCzVG6UmXuhdKbZzZxH+7sK
R3hcD8UfuIK1oaMpH85d/wFLhFaE9njTRL3b14tSbl7b/Yo8g9cVCMC9AAfX9inV
M04vf3CtE7daZ9r6XYg8YGxRwdd307b3rCckqNOtEiEIZR2wsA2+vN6vEPKCI6NG
S0odqAiORNGS1G0kEcJFowyPFFIYK5tcevQTCl6ZKu73fqKG3G0OYcq9jKyI4KRv
ELc/dMrpxJRZjn5Wz3QYPbHidbl8hK2rRPNUOr4pXka24tWZjKhG99gIxAvZ6FJg
+T48GRuMsh4u+dLV9/ciQ52IWruR96T9j/7+uexGwFub2TPJCchm4J+ZwXesEQHZ
vckCbqL+b8b/bRTCwAILRzQeeXw80fxAi9kBJtbzjWSu1Em8gY5LFnAbE4G1jc8O
Ay4ydZe94rMjjlHhXsX+w2LuFFyCDsIzRWKUyRD8JeOz4lROuQrA7ojBl/QKCDoz
2No7qmSNfLaicIvXE/S53SVUbIVIg8h/97peIa0QcFDOamT2s3ZWC1aLnCUAfyIA
N1hFdgzWLj+C0bsICT+5O0ZI2z4XtTQOvCPRBE/mohxoS2qb2atpFeDypqa6wjV3
Ym1T75MJTTUO0hNh0PAKx+PRszsLo/eH22rDLgxtGo8lnTpzqc54nQoQMwayGa90
OQXhgI/eNX5QcmmnMnT/xcK7rUohM4hMTT73BpnMQf6aeOeRRC8/Us2iPboJXKTX
PNvMvuR1ToORwESmHJ00HUr/3brqudrSR2mlJHaKrLNk0UN2JBWSQGv2DAWTQ2I5
kQBMKlevY7hyaeZ4KpbFhvF/VsejFmrG6u6k/8Plmu6kX03vZNZTboWIMsdZTZdl
6ooiacUl5XUb+yL8LGXR3f/bEPhPya5fkvMR+NFAHJ5VIVDjt0bbT6Vyam/DBt3a
Vvt4cEQflcSwIhFjSCbcdmaI7Xpdd9niAEyR8OgdPiQBqAykLo/2Pq/B2NsRznRs
usHFUDCL4va21sqqlyfSS/9tErHPdlx0MLaHErj+mjeP7mBVDKL+DEFwVDHgswJM
7cg7kiWVBkEFa6GcdPqtcA6oiZ+dORHuPsxZlIEqKhW+/aDx5sDkgS1BAfeaIhcv
8NWAAnuIfFHEyUWXf9HLQl4Fy3D3go8KMX0P38q6gtXaGnrH6JT9scufI5SCCwqy
GEfkjf8XYMCMzLwHOx4v9wBdfeS6ujtLag4pyN/LUiD7J4/xqAzYLQMleP3f/IUC
lLnClyL1Yi/imIef1WPzK9QVlrJ3tthaslIEDcN960z2wbEabX6BRW/EWZU0pw5k
nCfdGHVqR8j7jehdlCrvtWDn0oeY+U3vyPXIq0ZVPFw+ZQ5XffAxp2nFurcZGVBN
uGZHPAEONMRA5imrQCQRQGVzgBZ4We1OoIicXCdNpppuFyFdWFpAZfAqJH4EBNAt
d5WcWbuEmsdDq/zwfUJr838zwJgjWavsP22FreERLJzFHdWVYSzHtXJPq4qHghhB
cOs/suSHJwVMjnbM+rj9JYsKzqLBC1a9hw5FGWZPKGTteUlbL1tsYfB59WBMbxhH
QvXVn83qTv/rs5qOFf9Z7DC7o8d6WRsx7kIJ5yXQh1odeZVsUgj20OPBRyXw+/vI
YScNZwh53hpixrIsO6qKnXZzlWuwaqwnfNm1jWeZJ2yjf8mWWV6AbrwFOfpvFuxm
9LoBZeERRFFr9+1B1ZuiGShP8H+U1U17wQe+J42MQOJT9ooNp9PUBrHDWqnRvLob
EEdVr5SeYcApUw/vyOF4flnuP+78KltVFA2QA3nxPpGqeP14sKL2bwpsm91ghfnM
otdH1B8shODtJpVf2c0W+gbkJ4Otmjo5Yz4LdAqZnk79oQRV36DuK5thAHM9pDbO
/jqFGAqybDplYUxahMpJ1pGL5BtfY0RsYIVIAh8bR9BsuOAEGLDEyzqR0/tWiLe/
zzMqK8V+iXJkeTKquRg7VXoIU6VTtyYK5EFUVQletsWQOd457/Q9wdG4LT0lPFx0
S9Sud+qJIBPNvmJ4Da0+PnuRTSzvToAyTrsrTIZddbP1JKl6TrUSk8cJEdQvghrj
hFKFNuuOiDCu3VKNMoTWvTZibRU9k82xdvvVYFT/S3ULV6cxMCZWv/7APMadZ2bM
aTuPOz63pzZdW/2R2KE4bDrQAa584yHzAcDjLMntxRS7wX6GIqutQoKxK3vhfnGD
YtJWzJrl3rLnrPT2nu5/9XfhAK2rAzaFO1IA1UMt/zp5OhOsX4cUkSPKlHCsxQTA
SQtZ9zHSU7VC21yAlWh1in8uaOOW7yGD3qBLw047juiigRl2zpQHtBlrN6vvbixj
GdkAMrWeh1GT0k1I3olKfqqpU2K+Dl0viKJih5s9UpYCcOmg09a09XMlAXRtRrPe
iuJZLMMuH7l96ZQHxUVRNhYR0rAhxrxjOctoVPWQ8LW2Jj4UIEt1gDDw0jWBWNWZ
icy5n7svHDNcQzr6uvtuNz4JfJ2dszIBPHFarURWnj9knPU8KBwPUcpzkHHYPXVn
w/sKtEspzbWVd+xp7ZLQdCbY1CaM3CcIzCIyjIfwqUPtVN3WlZPsRgKLUxJyvNMt
648wd8fbKSxnVQE6TqRaoQKcarJkYAwdEyzRgWw4FvTi+QvquFG7c3YAcYyKu+KL
b6A4MgSeir9moH0euq1qteJer7DgnofqarK9j8z4TIO6yP3nhDMnN0ObZz6rnBxq
aMwb+vLtxdsUWtfIDOsoLN1I22SeN7hpQ/TAOo1AZ1jE4yw6SH6m0r+eP1+tKl59
EmIfT9fpUTKokC5eZcJUMpyVTTOkygV0fRuT95R1YoEq7uUopibHuf+wzCu54yi1
Yf0e18ddSAWnxfGSgbbod69NuTYRQYDb2VSnqxi+Enwu5XhS83Y3UWhDyzTfBC6c
TNdBBVK6Ni28jCIr31Zbx/ICtnP2yPul0P8UngCrIs/Txm9u82c5WwYyKwpbg3+w
wSLLtu34npI46P25YS8+6MG6+VxQBoj/ZxlDKwHPOtFL3qBaRSNkKjCMNOI9CiE3
4IOPa10okxGLo4M+3O35Fs23PMSNQhZ5aoqUGsQ2VG9hUGYwiHTaGjwoQuw8Yu0n
Uw6dOpRpWOoy39eUYcFMLmQrNTqKR1ZaySyA5xsG5oLvIS+z9+Zy/vz77nxIddl6
k5B6SDbiJIRntvWnySKvDDEFSOfOgyh0PtXs200rlHZ6fXK0oHbmNlMnrYHrsCgT
C9DVhfQ2EVOhx+QaPxP9bZ+eYDIeaF7uV3zNHFlK+G8aA9ov+TKu50qtdtSLlWiz
cmWRrkPkfDImQEkOVb4HtmAi3rQEYfHYNCDKjocA7KqKu26M0dV2wpOaMSei6ME1
lbtZAbOJHMSPWEEn7IhX2f1wAoBs4pp9glAHSq/DoM7HM1wuXsGm90o570JZGRBh
e9PpWBZ3mobIaCGyxpDIszemgTrBbLfviC4k4bGigDR+Tas5RLgTsXDq3ErByxCR
nSzsciH41wgTXyFRpf5yjE8vNcg8ZuHdPE0KE9nLyBIe0GLIB/zOkn3MJWAjW29B
SE/IfrBLLuhS00Adqdg4TVzUINySMhNpWYwmfUPH9ooYIVnJO0feEUlArWAcFxtn
EW22lgTa3ChpNWztlRQblpHLxYAW4QeTDt/xQ6/baE2I3ZNsRzGvb8jp7RI8/Neu
V8Z3q+/JBUjpLuUKQ5rVrK7/6sbkTuIWgsDdZhuQkG0FlJteVuUySVI6joQxDuzl
QWugS3yy0uiN5GPsSkk/Kj7GjkjROXkQQ39eFN/C+6sgTQ0H4XRWCdCrYvyQRBrY
+zvT3OgNKRNUG/xVVJMBs4BvIWy1bOwZVWlmOQ3d77rwi3yk8yuNRKhouk4/o96P
dIRudvagyX+iBE2TTrm7KQkgQbOKqGO+MkUEw4FLx5zYr4g7sJQD6dIsSWLkHthN
+V4bxU9TWSZolWqhRBYDeLewleo4YfrbTUwh8g6DS1AsM6xTBZC2AsEwPlEe71B6
YNmFWa/kVEshHHjlYvclyfC6LuKkv7tDiSSxo3v6JApEAFD3uuTXO1pCu2iBHBN/
JF0uwIscGCSdq/u1Rs/W3zaukUETq/Al1Yj7+cMq0xhUtKnvlCFIPfuTqyukenYn
3vjF+JoLU+PI04vzF8nQ5u7C1ZgvMAocg31yWGHVrWZcC4nM3Bj6f7xwtTmWtUjZ
9QyPXdq8d+uCRNN3WIaaRkZATUD6upxX9x4shor7CgjspcWGaolNrSLBGeQM6+Lc
avhMiTvNjVBPeMsYugI3z75YnN47rqWUW4YtFiQmjzWNpj2APyDU2M6TmT61jHLz
NShgS0+LpjvFvjBExTrnrfP8dUJ8unw2uwYnnUF2ieg5/Mr5cUxyIUF5/+b8fFOK
W9baanCiuodKhyF98Q2k8ZP6db5c5NLW/RE19clBVnE2CaxDapUg2PRYhhbKIfeP
3FCjFJCOgesYbsj9ldX0sEgn8Xn62KeWE20mHE1mF4vlNU7MzbsdlQPhPEVbzD3L
S0MEpYpVN4cLTLsfxXUgJ4Rfmovtt8xR37z4ZDWMm6fQ1WlqWUUZPJDGcoBQIJc0
G6nvsiEfbabX38vlYMAtIy539A6opcpQgfma+ieFcWiZCfdCcpMsPAtu7trXWHPw
CqJnrsPl8KwLqX/fZBv0WVLXUva2U31eCbGDX69fSLaiBnGuO5KopUhQ4BPDwmf6
Y+PtY21KN3/M4zW8dmL3N3dcKj+WEe0e+MEeB2Jt8895aW06ZiFHoidJd4bK1aWF
uvICjqSITvu+/gMALcRM27UsRd9u2NvP8Cdw8tSmpA3mt7jDc7PyKbUXw08zSml/
EisUX3FyH7jq34G/Fs6mBMF7yYrOxIAeTQPuGU3O0saKoEZiGcAWf4OyAt9wqGJw
zyEdO121xA/EZvGDLEQssuoTwwoYR1ExBAlsWFK05EaVLKjZ6p5WzarXgHJGkB4U
eDyb06+npjYqiKbe6xRJbBN23QQYYsqL4TezejyACsdY7aXbgp40q5aSmxyHWnLZ
3vOrzNew/hxNOw6R0Dz+SMqg9ZXqUjCjWHIYCJZJjBaEGbAzIny1L018Jiy5gRo3
fx3l5npqVEpwMpGrpkrCBxkCODuCLgYx2rLHwNWl6ZrVT3lqiLf6cUNC9RSJvmWG
xorcbaFhZOtkKgbYQpP/Ri5OJcmCPN3hl9wzMaVpj488xj9WuvWSIUthkzscFrrT
pG9kv3E9bqxu2lWIaioUx9oK4FhloO79i/8yjpL6+BSIxapQzMRtislRTq3CXm83
yFi9Ar14EHki4PZweoQcH8c7PG+3rxJ+/w7fYDY9FFejRVQdOW8LPyL80UxXjvhM
aGeqkjwX7VpkoSIai+hEfn55OkKK3lVADsx+DqCKDsJl8ajpqCInlPnVbN1Z453+
D2h0a+TCeeFX9Kmq8+UnrFbifqaaWI1b64MmsjVw1ONFXycVKB8Q8AyEQqLdrVBD
1M7YfN3+jrVgXYhD5xqMT58myk8SgJqt73CMdPTSL4k9Ni2LK+zvJKGkwEdMMZHK
SIc8EtGo9Gys6Kay2Y1SHcd3yyIWbKtHgVW6fC0+YtyeSr+sDR2FEGSj9HbIiWsW
5EsWQZtqUvEzCmFN1AxI2JcXpdmnKvhM4FRZyFuu8Ok+QH6upblTb4kcjl3IiVOk
NNZxWvRlnSu1oYAdpltKFhg4T7c4pEReSqidt2vz4aqyS4v+YbCU2mi/1hE0Lo07
eC7Y/Z+Bv5t9J54RoIwBbfLLCdUcfkjCwWxyGluvSfrfgHwda25vtXFMe/Gkwpjk
2WkIQunkVeGG+C5NsRcP8Y8Mv5pvWgS7ioo6DwF6EV8ZW+4oHvIdj57c7crZfhUE
wkaTk7CwH6cTcS1yT0cEpZwXLqTKdUi0kbfwr2N88hUb5v0jEgoMDgjBUCX3VQiz
twGaC+65HE34u1gRjNyFxjEBVfnfU/0y9Zrf0mRr5HCJ/whtAtF+A/3vN9MdyBRV
gNOZDqm24qUiC/+zLxC4KzKeRtCwVjG0XUGf02zdpBS+Hd2BjMv3+DunT9o/xqiX
aeskBRtx7lkm/Ho7TK+FnOv5gp4Ednp4mPK8IyNlct67Am2kF4rL9ubmYHwcutaw
NYINrJQTrE+GiSHpKoyLILz0OlgHTmnMAxnN0bRH9CKJZhYHpwYSqwlfNh5ZtZfJ
9X/8HtZXiy3FKZ5bOWI36/Q/LV5Op4VFgOdoGNnP8+/zk4+pFCdwXUVsNXz2RX4Z
RJ+vpDsxqIbPfe8EZGvq0BIWONdOvbZBSEP/1JJ/Nu7JOKOuKsJLZW8E34Zxjey6
7VLrmKDj2YVtNixr1Iw/y8zh5wiaxzxzWPYVRLU4HggiVdJRKtU0rd7ayfjnaQNE
6jsvCjfXkdHjkZ6e1BA/oiDw7zpco+/I2WuUMQXF6PX3TR02/OlbMkQbbPrHQfjX
3jCKA1GjkB0Iifl/ueERCZOTbsZ4IAQKjUrqDAvXJdP5YXKu6/RH3JwpeN4NXvzt
Rvm/sItyQJl3A5JMSB90bA7G0r0BQigpcW1JGj6r7qJib6laUAqstJDM+Den5GI0
YV4GwNTPdraYH/oWKiGBFuSRE57vulVzZpg6njM9C3d5Osr+KF5rgj7+PpuvUyxK
xdR6KZK0eB5locaM88IpGHKfxDFJr6OE2v7xu1EclBiFVno2DeAeZgmyrQD6E4LW
csusEp3XgappXImk1x82vTNJkH1zRj+aWPjHkOe5K/8GcZhmdhkO8WnnyaS6YzFI
180FSdz1/SE2lva2eiVR2RjOe1RM67Gn9u4yR/DLTslWCUPGBukp9ThHvNHYRmw6
Vxl3LZznh8+TQwP4kYTBfTC8rCxvU0rJv11z0BfcIXhGtUyIpCcqwxjNy6orr49+
EmLA0AzMG6D+Ug3oBR3+ScGSWU//hv/1bz/e0fLJqtXwUrmsOHxgFvEksJKoWKno
ngIw3jBX3MF6nco9G9nfYa4JB1Oeg7AnccsKM1iTLbWeBjGmYL2jys0OD5hs6+tG
Tm+xJjMnXYiW+gOv8Fqo/GYX9blMWpoF9QHIPUR8IIn9Yl5HWMOEz9x/pxVw1+j1
gYwqR2fKKm4xW4PEz/QNAa+VbgJeRbcwsW6NtE6cYKd3ePbzJO+CV646dQkbkWGV
sOVJvJXXw6uQvCVnYmc+cfRFUdaceIjSXeHzuCmJHMiI/i0udgWw0BiZfSTcEzWW
K8drwWiFaXMSApABi5nnl3n6BVJ6DgDXaXqsvP3ze80ftS7qmaJ+5BifflOWHVri
ts9AqBx7VTFKzdJN02oYbANup/ooIpqb2wXKsNhwImEyQf36evEKtvSOV1+Ka1aP
bZUmMA+Sh4YfX7MUmyxYJ67moXfOlsCamCPbaZ7ZzHjkkxxGyuz+v3QZfYaMiBdb
5jKmi9TFi2LI0kJ8n+R+VMmM7GblHd9DVGsI7PUT2puiXHVbzCqpKLKXqfc43dxC
Ln63yzZTPkFveqqbEJJDnIjSyPHPJbeHtJJzqyQeCFjgr6qtQz86cY3wggp7kET1
+pUqXh2aQ/82APpez2Apufcj4J7HUTYFhw6AI4NOJYh7Gln9lX9imV5UBcJ0/ScU
+7jMF1FJqv/eawR4PwkzQUH79X0sIRd6RpI78q/UqfCb26EM3KwcuiOs3gBN9q9W
cl69/Wy2Z7UmXNmGhQoez1OJbKjssN6vWjkx5Y+Nq5YY/dN1hRF7XJgcxJBApRfN
zJLgwLqRcInH3vZSZsDb/cqCykP4bv95SIz4jhsBvkUx/RlXnIOQA+7iXuRUnzhv
gZGiDwrl/WVOa83khTGOuFunXkBqTJw3BOB9IFJOWHqz+gUqiWGi5Ama23MnyKjx
Ly18I1h/m6IIJ6d2ky5jzYTqLs7ZcmWSNsboTbHkdWVCIcAVupgIE5iqw6EkJXHe
mDm5u5n+FpFDKvwnZcklFyqmKP/rmQ4JfUA19RRMqxRvO04Fn8BBdVIL+VCi6IBJ
F2bskiqewYS5IOzqTPljCJDJEQdqJ3NP2cZUhaCWdjpiudBeb6uTRXd4udjtus4s
b0uEQbNtNwpFkEA+mdIX6IhpGpOf1qQ9V5GVTnhaDeUtcR1RNLNbg6qVxFKcoaWs
3u69ljBJXMgxmvX8wjjpJ3CW8X7qxkG0ezxUrRHVOqT3O6RZd2E+INIn8u1stWPq
44f/RZFkcTeZy6OUjoK67FCPp7ER2a7oixzMB2mWBaqqB5P0yfO64f1VwL18a86y
eSqPhuf0/7hHkaE1mo0tlUNNmQSSMMziASavmrqkajufzp617En3bnl36oZzmSlw
J//Gj0SCCZKiMri8tN7JIWtPwkyvT2PZaMaeCcjyuTD6wioMXJ6EmzF1QxWPfm2F
E6dpqPa3qpPiJFoXi8rXfOHKyieB6IkFbR/OM1R+4IzFwAZ0HRLc9Sy3htnf1QnF
umgqCsaJreH4UO8IUdpIjwmzJ0ZFoc9V+HmiafkudKn4WBLcIUjh9UvI9PXrP9zs
DKOiL6JpwaVauspm7m9DChKHrXDGLyp0q9IOXsyVTVVyaH9/A+fgi7rdGdeugbO/
/4p1QYCC0HWwDcGpIvl4nIWUE0hATw3LH8S72DL+hv4eQSP71P+00A2GTCbOoqBg
N8oSEBjmUDN76HhiVfnkPsBUpAd0KEePEqkLPmaA6wMH6GHtuyAAm7dInuCehiaq
V9tqyYwDXGB0McS8w7eXx8uhg121vOhHf1t4v8IRJ108cm/TdLlkcSx67f32KZGi
H62B7yEuHF0OTA146OU6Jj8UYzpKojnuzFIaY8KZ7kx7Jp16F/tyyKiCwfngapdP
s/lgUvb8l3emMjMdvSTU/dkW0yQJjNocyXXZR9kDdyfm+wDBp7VtsNqvYoUhTJHX
KDfvZOqceusYdoGuDjl+4EsFQHDiT6F2as0YSjcdwjNSiPCmGe1OxEnPzPcy9pLd
lfCtFCFSJYmiqpW2bxZvMf0cLove71zlix/DH55ZlZMIJoB8xxbYNRkEPweba7wq
9YxR6v4uJGN2kxFSeVUT9b5XZ5to2Tbzhd6T71DKM4hELCAxed4UcoqdvQUTb7dx
4tCgS6WqbMG2KOwojmZK7ye+DN2ZcSuwGPxwtW8oq9VFI/AvnRZrF9qLC4ZLmYmM
RCBdhvwzC/PuNDGo0rsgGljpdIe+asSEg5+etDnn15m8Xgom1iL0YKOTqt/RQrEh
1RgGDGPRVkdYioUOmaOXgXfQe3XaDIfJZabmtKODBOSkNuWmO2XHSj8szSa2wJp9
VYGPICeJwIOkUOnG6QgaGTqDC4aICrIpII9n4zG8dw6Sxl8LK3iYNON0dCY54rfS
nN32wkDBv6EehOyXE+WHX6wxM6ZPTk1HYx0uDBLw1AYr8TaTj3zDs0Hcmv436bTj
9dnSf8hgrX8zfzqnLA8UivN3jJbQZx4OAJzjKCNAKiQZYYIRqQqSfPfD11edDkFy
8fnlsTK9DXM/8DndVucNjheCLRrct0zSEHTTnlpTbiiIwn7ucqP7KdzuEK6QI8WV
QpGV5+Eg2d6Rj5ZPbZPHQXLf3n34gP/v+oqI5Wf6OQrepeaFpN37EEcX97pl/7O+
W9pqU0EJfSl3QGi+1DRbY+0weskFUzGRL9K9aoNyx9VblKRklXIxDSi+5TojEc9e
lvyyLTsb1WLF+Lfa2V4D1rXG4wCaEhHbxMpZylPVQ8JaE6m0/t4vS0Hfy79Trfvy
XXuK2Lx+vNwXAym4q5vrCgvEAoBC+JK7D8tu6/MTYWqGeZrNJQaIRJbIhFduGJfh
9/P9Kfqjjh0C1jCow6+R2DmoehfFDJ2B7KgFKjYWOmAYDDZE94lYgcJMiMkqe2l0
Tae1D49Odlzz3Nt46pz6eXPV6HxMTHMLbAy2yoUirA+KCcCK4Imiij7YqTvDN8eS
r0OZoC6jpIkthYa2NRAMy+97tnIcVO5UGbPbCrk4OqqJrGFE7fF5t4z8QiegaRhB
9Qj8L79opvDT/n/Ee7C9k4fwhCMjE5o3Q6E9v34dWtUl0icIMaT5Nm6G4crgr2+1
bocInNv+zr7wZqAV/3YzYGSbKJe9vzK7xHMjv0dYoXR0U/fWQ58fz+l7zt8AP8kp
95ewdr0eg28q1JpBjZxwfBLlO56hIOSnakYqxhzXVmvaAfLzUZbZWxDeXBcOHUjs
Nq5b2rlYxkX8SU4V4nYUYBVNrnZBZB8NCFW5oWpc+LyaYLxSJHWpdOGa4z6Gs+ab
PSZ+IY+azKf6H31GVNZD1oTJeNp1Tn9HWD3ugPQcUa7jbmJLwYatkbuHQxmCHogT
lMz4DnNS4nCbtuUTERTcEx95J9x4Vqxm7N7x/QpKC0c9QnCTIK0qpcyXiVADDRHW
pOM7j3wgMvZ03TyrPquWFRpSfUZ6Qre2++y9nBTF+Xz79yzzb+y0mOljxezh5DXw
Vz1BxPz+K/s4oioPY6scErvdHV7TlROTYpFSr0qMUgDkDX2rUEUSsf29qzhxRGnY
KHXtKJMWkK/50zv+IQOz4oIgGSCXE7sqi/19rcHUn2tLzzfprbKwbWf+POsu7EAK
DoY9TuGdhPdS1SbU6y39kMH7SCg8OjAiOXzLQAUgDxo/QNbBTs6oEskL+4qOlmT5
/vMNOidSqc5aMxCQ45wf/d4nKo94KwfGHUHaWZROu/0u8UQ6wxDA7hJLuMgis4Ct
dl13DjAasEcaZ+1sDM1gZKbvqfX2TIwKw45HweGwjGzdmlI/y5m3xK7vyCst1f1i
gOxdC3GW19D30yF05ZZHBDSm1e6RhCtZVSQJuuUZ8Ard8r4Odi973tELWUYQVPvg
zNdtp/7J3Qg9pY21hdXaZThpA8bS9qmpSrZNLBcv7oEYU+X4g6aMBgujtEJT5jZM
pKqY0hhHZRenUQA/GvBRhotVfitSWm/YZ6/FT6V6tDs614LpA7GDJ+fQFqVADo5p
CRu2ElWrJDPCfPEih5GEFwNY13I2qOsTQanoFjRPtNTf6qX3K1fDzaw+2LQ4OiUW
3FDSy2p4oCYxhOzDOBbvF9wX0+RgvySLFG4GM6oExTMTeHqFawZh4iNNJmGRJ6+t
4Yu7d6PeWSCGU6Rn/yKFC1GOKxgTzd7c14zBGaYLfoa6nPT5fgmi3ugEv06plmRZ
YX2gHZ1N+pGT3P1b1DaY96X/afeAfLDdGZVQhflZGdsbZppSqAIVaI0NSXG2YTny
bweRfg+AYqQiE4mq5BEFYB8ywYVWDZh19i7+IJgJQJXFP3OXZ8H13Y+7SVXhTDl9
VlaCrPtNifNviBywStigNBByAAmoSDn22EAdKghlTQQsQGO4HS5J384VajNL27OR
GFvoIKOrNllTeIzu9bnL7T4HiUb8gyBdeGNZaU3bCMhccmJp7bSdneY1/CvVXmhG
7BvhEemJjJmvPEdO49YhY4bqVArjm/DwDvlSeVdeoywxObx4oK8TWm4c/ILoJEwS
PPD4JfoY4P9LZtjmWKwl1JlylAzEiRdZ3bUt3WI0m2M3RevABi9ifxwVpLA07R/N
Y13/2Bwj91cD2BhsOrXSh7kERUFbEr9VoZ6F+c9kk5wuuGWeHfOVSvEkUPoLkGMO
3eHlC+oSqdg2jraCrYJuhIt3nxpvNqB6P07JYeBPqyOvhel9VEayMx2SVpIpo2jg
LYtJpTKZWevp0wJ7fvouX4IeMSNrowsTVo98jLDmTSJtJebxFeOZQkiIVLgLcTGJ
5tgrpZTI4Xs4Y5KRESS9vOMktM/oTFo0cdIUg+kv09nrKzsnupP2R0zAcVfDRfZq
c9D6dYx2jZbRW/R3FwrEgF2VirpW3pqG/v3AV5aUsXbaGqjyccRTqghmVr4oijuy
C39wkkD/y1uPNGExHy4kOuv1Ooe9aYGu41TKjkaRF1u7ByIQfnFUmaKtTzCIht1e
Wzsy4KW9i2sdNk07vtxj9xtOMjV++aNaY6jFwBcx7OccxBaTF3y5r/H8WojWu2c6
Q+glfWDghFeNKJa6e9FWhH/d0PY9rYdrcNrQXa7uMXluBXBWTfUbQTDe5T8Q+/vd
4Xwc71iClBMCbked3aQn8GglW4fatRY4pEgXj7i8h9GFMYWz7eG85EI5yzQm2FOJ
33v8QxdeVy0jp0Z2rMgkT7nHD6LttTXAVF9Qb72M78i5FpKSiNr9mg8he7M7xO5U
DvX9dqgiAetmuVCTcff6FQZEuQVHP51jpqwcdUC32vrzZqzHOIx/XoyahDOqDiuq
N2lFtVeLtNDskvggK15nMcjTTpplifA0E2hPLMjBHmadrI85TmeJeD5K1WzF7/OL
b9J3sfxfQwLOMLbvXI4f2LpU3TE5kWftiqbiDurhNWQHayiProM9H4uVmlJbYQA2
+hPjJyv1RSWAg15jgGafJZB/+iewyCQLykpcFXCblfIL5ADT3WFOSB8gqhcVs4zA
d9JgWLCmDJJZLwJ0okzNLFDXvbg/F99KlgQV07WiWxbH7QDcGlR9DFu/qmIHJ5ji
vszOWwh2JTOaaFpqSvh1Cp33WBPotrQ9WTbZ+Jke1Ohz0AxBbQrQjGhR7VPYXwHq
yxVTMducTkc7KHBk1uTNCMbPIDy4Ua/fwLzyFpoQev5lqC+HNBTu8tTNdCA/JbUe
E/eZpKSypailK87L1WHVu4CIQsqbWY1JRwdiKqMeEHlatx7OnRQKEGZi5+mmHQiw
ABrPJl9qGNrKSeB3Vvzj5moYh4A9PzoqIFWbWDT8fSe1J0g6pBvLD5MqiXJvd1zM
Mb5BfBWdZSCWO0bxxvCjU1odM+bqOuHwRltMaXSI6L134SPB66cPsu4+t6uecfXa
PD2jAU31fx2xXscQi/QyDMfNpD6UrjUiuskkDAf8plxut7lfCtw3q1rhGanpGBh8
LqKbZsDvYZ6S889g+OtpBX/AO7dhqm7mj3+jjKtClfu72JjeVziZW6nHjl2Hm56D
mLEHqO/FLIcfhhdyNhzzZnC0RZy92pQcj0RXWIKabZ33MzvSfjH/cmH1HKXq2HNT
XT2M8kzlgua0EB6NLEAGuTvCPC1TfJlfCAiuMXKWe60AWDf3nEJ+qjPs7H9FHZsr
itMRruyDpIunMbyG6KwsdOpQniHppwzcgQ3rU8jnRICz+WkasSoxUz60BijgbSIC
/WI4xJfLFN778OUlgn0EzLe4c900jrYIxHr7ro7lLW8Ipm/aZh/svheySgJ5lpcA
hCaNWS/tBbE6YIdm/ucZex+Mws/DWYyA8YSqVrs3w/aBgVGnZA9C8mnHuxvDAz65
Pj5AMsHCUDmJrn7fKVkEokL9rV+oN/vCbsjDfuE/rRfeuee/AWRaOO+0G678eS+8
8wCWI+PLVdO98vPFeQRQ/1JtvBXNkpAQ3cuP8wUkNdLYUQwdMPnnjyNpPBt66K9G
lU3BjJFykvBiylcn986BEESc7qhoNjpAmBmss7QT3Vd+JxgU3lN5zaSu7qTDoQ3I
4ue1AwT2yBnmn9owjW79lUqsIOLzYAoo0H6hOaHaNTdz9Ltwwfrmn2qxsrAn/DjR
TnpE6qfQQbdiF1hNWpf3rZDRLFj09U4iYDI+I+63IAB+OfnFOPb0i5jX9PTfZND4
xpVh43ZNYc84W3sZ+JfK3/zEarHvHpDna+OL4nVKS88qutXOBBTD21P6AfRfuPZh
k50GY2WhXjLwhBb2xl8MGQiHAcxUL0lJncGcRK17KlfiGjgJTGhPG+ErnTQklpm5
99vkaxfgv4lRNVkMMF+7fWAkrvFCxCyDlr9EiwRbDnxyp8q23ijvxlCyDraJUiKx
/zUVAswY+gPwiet8WaduXT5RuofmzUX5pOHohAc6yxUvITNm1ZnYb/jxbo1Kwqnm
P+EEV8WM3hx9R8ZloILDv003z8V133LGs3eVxTzrmIkibrEdyikzbeVkLPYKQVRv
CbyBtBACPpH/F1/hKMOm6F4LFrkiD3eNl4sJPJg7Qz5WalrBT0pldPCyXQxgSULM
g/qXdBZBhWKWjosqW0pSdtVoJgFljdXYnBMF3Op8jT3vbos2gpilWTDjw6xBlkk+
NkKFo4ISxl3lUrYWcMIJ/qag999Wjmko//1s9xa54QRTZuhCrLkJ2yRzfDURcQao
86OMWJc6R1A3Vf6pvG2e/NWM0N0D/baYLmc0b9HxUk/uKyRGqaANYiPzWwifoYoF
cfjXt9IEI2V6wIC9Uaxn/l3XMJ3IjiAB4OWxW880+U17BcIgy1DnrJR+BVeooQgT
VXk40MLhbOpOFmqJrbYoraZmCJgFHwQeRqKQRCGySKcnvtwFbdx5YaNiQbF3CSkz
nGuo/Ky1Bq4DQZNEEVWZ8l53L5PUDc0Ydo2/Ew8BkENf5aebhHsTOz9NpaGL4CHy
Wbqcb1I9zTTpoSgWeaUTGRfLjsWhVE8OpoRmY1dUL8K8EGxYMFxZBna/te3pkkV4
Qgl9lTi/0EODzF8nwJ8LQ5dZpIGwEKS33YmOJio0jqC6d1jO2m+cGQNK5axqhRlA
iZ4zJaxPE445xREvMlAEHQ92gB8oJi02eh7P0U/rQUSZZObBECn0f2lWPpwYcltw
RWeBC0oLBgq7LAdL1Bq9hlmV/sRBSVWfxbdLHDg54LmxzbRhNtKRjzxi0FVugFPb
8JYZnAv3CjyA+5xnIqtIbvpkXHdnkUHPqUCrZInDpTX0XqpId2/buinLasCx7cc6
6oB6oib5h4RSfxaqsxIv8weTg4BjU2b3ZphTSBbhFteqj/Uujsi3MtpUDkoM/k+h
lp4tst77MRva88bkxpp2uIIbNX2zZdQA9T7VSZqNOtahLL+vR7n0cpaibqRsE39r
4JV9sJHgVCpSOpyj1ukRA2JCOl/ifK4B2vl25BWnPUmzR/rdekwVtQFy8hTI72Pk
xlxYFnD8nWxaJQRRYIB76LxhWvUhKm46eFHPpc0fDJL4fRInAaOoBIYYIWIZV3S1
ithIcGVTd5iyG97RRN4RPFX2BVYmFRzwTK3MKmSd9aMlGDz0heEkaAv1/mUs+iWp
5tT1WcC1tZ+GlI0+Bx8obizUrl/tHRhN1SxDAExUH30tf84Wm7WoViba/Vb+TgfH
8RXpjRExxCvzxznJVHpl0WkGbrPWs///WNJ80z9uDrfoCLE7MryHSvMckWQCiw+q
HJBzQOtYRQhUPDlANRSGD1obW7BFrgAG5nhdslnisu9HPSR03c1SX1J5W2OULtvX
uMj+z/dxzOZ4mPZCATnCBG1ZWVbCjL9pecDJycuSqaKJP3lEHMOHNeT+IPEomTX4
CmSNZf++0/b7pQVTDOgl9MSRsfeBcIt1+YZdd49B1oYwv+LL/+8Er1Vh0W5EdLgl
ILZAcQeuaRJkIKL3i7wOAByCKuRfgLOjZpJQSJt0AqrVG+i1N8wUt1Trp3dDz1wS
DhbvYGVuYcNMah2Rn8vZKGHtpik7gsSLbvyF+48EnkGX00bijMOA9dWg7HRCUzDp
i8w7AKmiWFtqbPDRUkUFHhAPr2LJ+/to2KKMXTeUJs0rl5UPzkPNf5Qh4ApxhNxH
2Ns1voBOcJuaFIWrQDBLCgEO0u+4Z4FbIUL5KtSJQiD4apZ5wIY7DqulPhidaU7f
4moeH42BiFdNGrOHwMcSuQ2II69fR/qA4THSCzGQ9GcD7kRH+7mUB36fFI8d7gZA
0buQdARRAd4Y1o0VVy/BcWTyhUwJrirIeXWSqVdOViF3QxXNKTpESIysHwtUYrGx
zfwH67zkPJN+hPVj3RxbdpRZejF+HMHgoQ2KpCVVhlN9hfG9FuIbaxjcToogSjdH
QquPC2CWOuOYlof9r0VSsQWfGr3icJ5F+X7y8IiaXt6539WTR65VfYEdcwLRADJm
7ltdbzHrsCdxpIyaIhxSTphP0Ry1I0bG7Xk8H4k8MIbqKPpWOVAOADT/7PlcxeUs
pflBek+t6Z50AThDoPJyWeXl3X6g9BGtMEN1O3144Rff7JpSJTpoplFD7IOUMY2M
tFt5TFG+8tQt5Dvt8LkipyxRqeUT25iSPAgZI0yByTYTMtgzLYzUTwUzJUy0qn8i
Qp4o6F7iqKOHiJBegO+0XI/3khfRL56QnKznOUdFJX3PMITFkzeiaNCU8L6tyQvR
A9XV5qOXIL3LLNNTMzGQuNArUjf2qAQ/AnMDgJK3FSDsh8BmHqm+yvpUBEiCxyfA
ooimLgAO71fbdVvz23L1P5hL0HWpb7SAKPUmP1yik3LBLAnmXbbMTVdgRrpMJOQX
TwUTMJ7E6XQa8i7+aC13I0GGhEJ4JP03lkOwQl90Ty/47CEs2lg3iFVwUnVamzza
S9PN8A3YeKm7C8XqI8UsGk+jsQoYk3BtOF8jaQ8Kdb5x+AMjeu+D/CjL5Qjf4ugd
8qgup6hlOn5lO7fK9oymY43O/NlhJEe2CLaFNpUhT+DdGynxf/rNKas0C2533KWz
7Pu7RjSq2M15/U37ERPl2JgJdZXCSsvBT0uoE0BOFuBUMvpWC+slkTMbM+IPErN1
jkJx/6R7gGhmxQbrdzVMiy6/5lxtg2g7/+Qc6iT1SOJ2dtW/Rn9OBAyPpFRtJZIJ
862j6LA6hD3Ni8GGiixJ3Fx1mr0zk6xK+yaeieSAccElkJ9NpFxqpeF0pc8801Mc
+uD4KCLhkfjuMuDIwpoVsM3/847VLdfc0QOAs1KYOJDRxcCmCzeOABn01n5dQGQ1
lJZ2QiiViz4faUcyaYaMadLju2Ijy7yHRoON5rSXYWnd2DZdr7J81gK2iktdQVTb
NoX8px9FitNzZ+CavJ8pLxjUACj6TC5Q4arvnx4dsQwBohOKtnwZ43lJwwMdCDNg
/pvQi1yU8yx1+9V4+MD/DQ53ms9xpJtaM9tbrd0Tf0Vsni5xn2j1ezGvvSGc7YTt
e8zvKSV61kA6oqlOfVSQfs4E3dJ4ZxnERNN7YNYoFyNeIH7he6IUy4EX1kzh5Md1
f1WYVaeaCwCcBUW9lZX31GbGOxvhaUcbC6ZGTq0XnMKwbYbZkx+9y1VavCDFz2Kb
alYgoH1CGMEyJvkNWn8LqmNwwRd35+XYS4zewGG3k2t0Eao4XWsRbOnnAjlbxWZz
kFqunNb8cCDP6wbWe2FiNsQ4O3TYrq6QnfSztCkOILInc5kDUMTVZZW9/aX4RbtH
ckDUF7l3t7+l7dy5X3YCDEpE8YwHNP8a+IXn0OxIMsi8kNQ8k0k+17xp/v+TZog3
9NPaVOHb9M+Y3ZybQ2kpp2BtuTkja2/oNLME6Lv76ejfS9Xq99UbP5mC/7psZUrl
uJMnwVhIzbdvbprv1aRsyzi0XbVDfb3klO0FFLeVio/ogRkFqAezpHz0x4/GeL43
ObBgfVitMcL4OmnparjrnRIUgHWL4Iv/kFb9FiPSR0DUAhs5JqDcrtqO1coruiGS
r5dG3K06uF4eFsGHVcLUzWOs7GPG71cXP6le8beQ88aup8xzurSPTHqkoNO/32O7
zhGpnOvRx8UfCA25xXn7nvHF6bDeyfSVxHbN7ZEp/fwa50xTW4slrS/gbomQb3Mx
4X96uECo9+RgbnI1R4z+gPELr3TwAdfGcz4PsoC5CiqyHmgtCIhuxLIe2Nnl1cCX
3FS96fd+J45R8ppo16ddzmiCaFoKDt1E8Nw3OHNET1JBASOv8KQUeFbXzG0wn8cM
dyUetOSgFukmbyEUtKWfJWkHKYX1iFG/iVCyBHJBZpKjK0RXPuSiyJ2YMksj5zwe
fm0vlyv9MnO9uEw+2y0rttD78/15wJObrGfjDL8HdO8zI/LtDZaAz6I4yp6csU47
ANpYamQBHE5Lplk7TTp4f+iqgoZTiSnv288uvyKVG/WqnZRRi4hwyqYxXGD88yz3
Fp9goiXGqpCIVhyjCYzObcVpJb/E5grexG79EDuAJ8uePGjLL7Ei141E/idcYcnJ
cr8AVFI1lzVir5AShfGKCNGt29LsWTpuWCKUA+aBQME9cM0VjITftZjHkEhhnXDt
tfasO+HwJZhXwpZk8tjzzCKaPZdY6G5S+i75w48YHeMB29xQVR1BAHpH8axbppPv
iimYRPtRNpdHbl1IzP6OEqKE2A0eC3o8LIEs09LN3xb6/4VYw7Qx6bDzHRkvJISj
sGHcj8XBU1kvYyKahOHAX/hatQ+URlhz3dY+ZKGJcVUjxQCh9egjb/cuNQgAhOP0
zcOvgrjAP8nLsSiYwIAu/IaKXOSZs1IJIihYBuyedHQyvu/0Q86EfAWqPUVJLFQB
m4nvnX5v8AmT0V8KBCc088XwGW7Gx3rjZ6ZtBBeWRRKm+9BpQ2pShbBBaFBnu5pf
vFeDoG06mv9QLfFmPxL82OxKHHs452Vv9Eaq6IOFO4xpKg8YrmObgnm9MfwT8j1Y
jT6VKlvh0suZVCe87EwARKBQEjXOYZXrPN4BFK67MCWr3o9fvS5GFVGkKcNF2CC7
0EiZ39yqHdapQHhKHXxZf9IR5l/243bQeqxVULQk4wtzdwAUqCPH8JUotgC1WuaM
olZimqkNQoqZnzbMDD549tOm4fbnu6Vzb3q1eYp5jw70yhQcHym7bsY+FLqf3CTZ
n6yhw1TjM0t/LPGoqlZrv0qjz88WNafNAzdUZEhpJ2uEDEUkI0h3TOM1hX3g0aMH
rj2+T2WAgfYuZJ38H4GVQLl8LgPRikFi9ngYrqfl8/XiwGQb5oAOnVfd9mV1g88F
UDBEyNkwzBJF3gszJiIotWK99IrTPvB8XVGJ3oBv++6Br8k/ebTblneslTvD8JIJ
TdXJuQLpGJqmalQdfB/uwqWWfKH6cPNzYrWpsDRaNPLMMjI1b9qmLrgC65xiO+qg
M8nb2BuIDko1/pKykHHNbDd73CVSJWQhObaTCJhRKneI/zmOGM0GW2deAO/Myjv4
toSly4wBKKyLnCoWWQ1P4Da2kBY8NQKARlW84v5VQhkTl2cHIhVhI6pGksWbvgOA
1gGR5KT2ZsKYZw60J0dP8UFKfjczQdiD3hADA0RtyKcrQg4PTYohWhr3FN2E02gs
OPejI7zN85ra4Kt1AYK+X0DP1978txD5wwvlzlcmDEm1gGGZomY/e5SRHkM6uYNB
AQ682Eeisx3NDI57MPr9ans68fOFRmAd2ETejOuHbuzjpNXGIUVlDw9ooGy7LkdT
6DxNCgZIQTGJWcWnv+JghfjBo0mEapx3o6vSqMKjiSEeVvTlkEre6ZDv0+qz+hy+
T5WhWezoLqlUrFCco40NDYFzXv1wgdtplWs1SAK52rL2NJ/M+mNUDIE9Uo+lSWHH
IjSwQ3Bf0HmWQWfeHDnk3kiuGe18bnByn3VhlixJQFwElpzbREAyxRHWKCCnxZq0
YUaj7iprRCx7Tb2D75b8RFf3RL/07zrZ0IyMG7SuI7t3yyVUNBm11QHl9KjRTeZy
02Vdw0aQjps96pPfOKztbFf9Tv/v5PpFW/ccBIfFYmZ7CkojnfksrvdXV3yF1COG
DZng0gQSl/f/niXjYnd1kKYl5ujFp0UYORXhaIa3u8M8xwo9qt4n65cpxpFmWgsx
kcMDKEfZdZoMFCjMC15hInjeVvqk9g1QUkEpWGyumPBeWfXL5F0glRqqwxL/HTXq
MDYfw3J7hqcFsPV14xp4HZbU4STPQucsr7HSJQqHX1d6DpW80DX7lgmNsGsvupGx
/yWWFAs4p4novMeW3FG5tt3Y4hyFZVMyu3Ha8wM7TgU1EnFJgaZ76kSGVLG8HfrV
k3T2aCscIqpqKtSTzm9p1uo/GvC8iIwD+ve/SphDQen706R2Qd0tZZtyQUG4u1Tr
1BiXYQZUXXyHv+lLLMTOjFmlA4s3xqP8lFSOp5A2ag2zK7uBkiVAzB1WGRrlnQJA
5bIs/t4roEbEcYXM6gjVybOvu+L3KXf6Q5EVbPYo+NR6ZkJsrR1tWb/ibC5MyXWZ
D7UGNXevynFy9sC7clyvbz/7cBdzbkK3HmmXVsIiVcolI+4Z9VM4w+5rIRwcp/KP
i+5QpDGvOxuGcqc2sTfQifYmRO8a62XY9piBy2RaZbQJ0PkJZGFbrxnR+uuqwM6W
N6vQ3Dp/YZllLU4e72eL6byFgbDPtob0v6LrLFr1MbOOphaX9pJF3dQt6yQqi9nH
sVPAuFLNojVdSOp3bbaOV6tNtbuvg9+3Lpi6yXa1GtCbcSUdmXasXjp94WAo3Yc4
DtvgOMC7vg03pwbN1w/VCvxTSyN4OKLDRmb3FHbXCnpm7FFFcgV3iqa22kzs691y
gO5JLhbBRJey5u2ytLkRuuLL8EmbSDwpltNeixUl7dkXzL6DlI3LA2OqQtJw3ZwN
VGkg1GgFsaBilVaXytIKQ9OHV5ND7eR2n4oI+2Qybu70tTIRZ/Ng8VgzwwZz3PUu
/gFJ8Yg/jtxaf+g98W2WrjaIwGSfbGSQKUu58izIcxIKz255/IkvtQJZjXvAb4b3
0H99MDLXzuPzfKO7zU1Zl5/wlxGw+l++f0iL0ocPfz+dTC38J9d5vDjkB6Kb2Uyz
rp6KP7qEhG/qAw/KkUt7nEEJenmL01CFG8xFPc2mXUolGBcnTY1o6NF0TICYQ/mX
F0TLXZkjM5MYEvWQb7xCqNYk3EeRCBgjKa6hy2TJYu8CEN3m7Xz855FQ3DXotgIT
9R3KoxGoJvvfTrZvJTA3OQgEfj9Dz/VxO5w08FsMbYxYrB63quS2287GM2WThRca
subb7JGUTxzranK+IVgfZdOca/rNvlIqzh4f2DJVilKdYloM/7jyUH2cHfil0axe
PLsDtJrqGJvlEiLawcoYQtbxiZisPqzvA9zge1QwyyolWJDA0lZSH5Fg4UlORx/Z
L7EzaAcgH66F7kjF6QrEjh8E8tQndjXGPGvqghgOtU3GdWsWI3VV8bxP7gyi3YbM
NtikpoCmXNn/xAY97XKh45vpV7k+MT7feJ78S60fcFUW/kOUByh8bq2wygrXJea3
N6QneTuTIbRvu20JrLIof0YGyod+6iZ22fkaskBZK1cjRpXFym8wK7NfKHQHo7Hx
kzJbNbRpECl9434gyH4sxlZ6ZJLtgvp42NOP1gaEna9rUZ94Yir2cCHF45NZBldP
Oz5eCDgoY7OX6N8tlO46x++/JAxzWKUxbP9ZpQ0IagzzzNRKc7PnkHL2wA54tvtV
arVmjdsUfRN7Z6ovVB5py+wOC1fc+mECNsLryP7WtmnapW0d53/9ceRwhdOw6Js9
xM9EUVdQ9N6fR6WNeKowdKkz/W2tXtRhAqizB4nP7CUnkCl3pQcZxeFDf9z81/Xy
yhUB31WAWWGFRyt/P06A7RXZ34o77Bha2P3SJEoEpqOhyU0e/YkNMHJJOx+L4RIv
5FcLR99mi5zU4lTe/kT5LZu7L48g0Uz7tmKvZ8Z7WkcWJk4usvUhLi3KZIRv4mvk
vnsy8ebBWwPd3ZdH3hmqxSXLLydhXZz9gqu9j/WuWlAkdYPe1G40Dh3fBfWky/tA
Uh20BcHxwSjmYxLU9hwpJljqwDnM8LPtE4qXQ5G2TP0NuCVlz7TYxxd4f6W12YlF
oApaQpj2GjMwf2KEiuM8XMxdbR3IXd+zppzWL5qtFwHmIhg9SMu1Qo5kI0Nk09lT
OsViaLaKrsV5ZKvPvvA4r73VM78PSn9P4YKKAtUjEGj1eQA7DeHEq28BKS+KEJkK
l27y8aBVBnLe550/K/L4pv7LzJJgtt2suxZ8QUcC5kCW+ZSfzKVw+SnUU6JBxWoZ
gxS9sbC58ucBgCFX2S7aaQBwo5GM3bZ2NB4dYy0sxHwz0GlWG2ODthk+WPxsybNa
o1xOImLX0b8haR9kCY3re7+OOHbcBRzZxevhupdo6tC3wPgdKVS3m0EqRwZM0DZk
JUIMMKx/zkySpPtQLhfI0wOHPIOk4X0bFa5Psh6pBVmz9ZFX4IMvlD8iVevG8Tna
pNmRbAQ7e1dSUdPNRiNVITW3uvM9yjfxVR/ju25Gh/KOeye7CTk1jJ2xNRPrXVx3
gDDsxnUnogOMs6KfQxRlFCoO6easUoBRqCmtz3kV/gmq8jlLX3EZZNI31PvTfEbQ
bwc1aMrMMvieUVluZFbpyM5xeRAWo9vMX9e926KWNxru62pXy3t+Qq9bAxc89Dko
GYY3uT41cKGH7aN3hBnl9BOlUO51XH52v8ZDgA+VqiNB2xhGJOfK0ZXjrrmlICLA
NVz+uOkiTFAwCb/Ut0ldeAWe/gXYBv+B3PmI6FEONmxHD4F/PJhtJgk3O6B7NHTS
1J9woG25MQrLv1gH+s5JeZ5U3cQsqS5dJoMzWyC77gC9767hOkiOaBaIzEIzjFJu
Cmf2n8iO4exQvDI70xhSGqb7mshryX/nS77KNvJm2dOgWF/gUS/qUVEmQ5dOYWOu
cvyUtDN/0ZnhCq0z/jnRQqW7k0JC+VZahwcrLzwOLKZqmFo8ZAxn+fG0YPfEBG+o
ugwzGEmgx7rBuL/ASJbigE2zQIlthTDhyn8d5u16XBGtpLyY8ZamnLnqotfxX9+D
+2tJBc6b1rby0I66BkXwVEsmaV29tWtltThp6nRGJaSE5U0bFwWJms4dvdmin74c
sQ6Ouu/s4FibzWa02cFXsq5oSGuEerHsNPghh4YcE0ZisyUULFJeyM0vWGLQnclZ
HSP+e3MCymB6pQ4eOQUqJU+Wu7XRmq7fqVhv5peY1s7nu7hskTzs9C2pawvj72XM
gqOWM0StTPkHn1cEC7AWLpzQry49+3Vf5E7BqSdU4aIEqZgCMY1NPJqNaPdbR/hV
6lLRLgmorbsDGGibgh1f2bAVk0Y74GWqeyjb4xQE7DRRLe4T7JwyegGTlbKei9SD
VzBB1j+OQBWMJ0IobIb2wDw71zK44Xb58q6SlT5+WYmu4TjV6xwrOR2jpDWSc1qK
mc1A4A1V3pViE0qgN7T/U2iXGJPysEJAbcAHbIiEmAvQwgO3ALL5ZJ1AM8c65O1n
f+frla07PJK34ltrGOUSpA1iyvFDzLzHT7F5E4sg5+6jSVKpvwtIIJ5IymGYi58B
EUTc6h39JFeD06xsCw0MqVUQNpW3BmhGGbv3davng53w/4yS1KP3KTK08GX3IDJg
fzwCkw2T966KHjocUDvrJmWeEvwiws7O5wduuuVvg8DKtBofDXZNYrCD0RPRTimD
I+u9M2IMe/d7V1hqbCcZTNo7jXptPVa2+il1F8f/xhTo/nAPMLa9QJaqezIs+AeJ
NYUykSxbHjke0G22OwDrwR+mFWLStIODX2rInm+zulXbfQYT3GKQ7bpqhBtRJb4s
91AYt3rfKsOciV8wt/pHJ/uDP+2OKTDm1Ci4BQWpo8NtPNBAm0rWLm8S1m2SEEsj
YNYQ2YtZYQemwlDa7bFO50cISAQSzvyqLe+z8gm7SNsaOuq4Fr3UOyL4U5iEsTyO
3cINvfBEdEfpW5OaB4sLF4141C7CH9TXAXQcwMvOQadGwqNa1X5/9W2txX/kK8sh
z3pOMgkhmacMxQHwS04OwELsrY3nztK+5ycwh00RWUIwn8Bmn8NF1jYQBIIyOJPg
FxstxU5CHrMna+taUYlznQQ9X2MUpTvm0y325qdGAEc7hqlL62JSJkE5O4ZIpi7c
34/iloO4ATb0Z/sYJApkTfD+x6DGpr4HU/WoPbvWe7bNZavVb6pKvDB/vCEaCg43
BoZrRKUgZV+pQK+YhZ59LseEkidJxVHxEHNp+YxCaA2XbAx+ECKr9LGDzVX0M7ns
jTQfVsMs4fyd65mK8j92tVZV7CRzSFW5N2PNdiDhXwEcsOhHkGx3alzmVSlpafi8
XqBMz357EcdPZU07QJxk4whvVJpv+CbVGWnA1UfU8qMxKGNmj1nyHrneUCdkBRiU
Q++Q46H0u9WNgWYE1mDJQMtodRKApVym7idVd6T5dr3Tmh/hJ2nCaw0WU2GoOJOD
hNzGCPduiLfCT8gr+queWsQJiWKWrxP6/Z/AblJgP0NtcfXi7N84wDdcRflSY+m3
Tf8JrtI0pEV3NUZpLk7O9q7QTuB0Ejy8KeUbpwYFChI27WQB+Fm5L1aY7wY8zpsd
8pcJ0QVR6yK5uy65W8+bwA0n7CSrPBwU3JgbbICrZGFNT5N2O/LX+kr6iM5qoUV8
is/bDdiSehb9x5Ov8jWRp5GiyQ80XEv/xxscbwcSr80tc8dbrcz9YyLNBmsozx95
/yKmLBeYE/tvaoyEzGuCPOfj4dvWix0Z7llpA1l3DmlGrzYji5bY+Vnsui5IKUwA
lRwMiyVoZsLIM3+mI9klTmSskdSG8TuuZkidZETGKdv+VFydiJIt54fxyL+i+zn7
Md/z9+8GaxKIiJmajnKdJyCmgm5Z/Hf7s1qESKFIk0b4bG+C1bgCug7fcCrWU8eN
FT7S47ho29FrY68eOlPGdd/hwtwM38UOqdtHOYJd6JGbmE/A9sixTtj4LD0onLkk
tcAgM2iZ3L+6zBpPUpqaEI74bqRvfXWXPxuKBmD0Fpp3gJBCZ5PyMqZLRoTyTrbt
LtYTkwk6s/9XlICfuCvQMyphsaGi3aQkixlqD67rZoeWt0s5kfvf9Wc0xaPDj8QQ
7WR4dlhzjZgxhxZftJutpQDLDNgtFMt1+Gsa6fRPPlmftUk3jRTtNJW88xzsqtzd
/PLzV+W4h46b6mf4Uv/whPZsN9UOM3p0eQN0H6f8xt3Az7d5i1kUNnZSbMujl1KR
JDST5wsszZg6jBftOA3Oip3ugzOd+kHTFCDH9Q/Aj0UQjYU8xzfJK4WYCDYPLmBR
ErqP5AulTPWMhWboPp0dSdzhqME/CHPmHX7ZHFlJWkQPtOoviun41wLHhBaXOoby
+BK5TgZtiLTKV/bgF03bqKcRPOAoR9FSy++VA79V4xAuSBxyvouDDNR3hQVwX6hn
PIAlNxFfnD98TBbhI0tlzXeAjJnJrSywV8HVL22Zhb/l8nJ2ew+w8sOQ0C2QDXNi
H4h24zzrf1Wv8IK/DdbwLxj7cZ5JCq3SmOQb0RfQmvxXVSM0DygTJeEXdwTcG+GQ
+Ptji58eWm22EetHwwLHEbQ+9zKB+hCCTVvbgE5/zGyug9m+6oCdbB5kuJJb5oz7
ueuHRwhy8EG1IKgn3t4ec5VQ908MyQEpB2Y0hZ6xEhRnsSVWNAzJUL3E2pRygVFn
ag2RercJllOBwOANtZ0IR5JFm0z5ExYaeawSYaHx9NmJ+lR4YkiLzKwR8dFVg8Hm
Os2Sy1eLOeQWZuQ6dRDD3JlDT84aa5d1TO2sARkqcXAvC8eaeaMWMKndugvWoBw8
JcXEnaniPXDMPVSTpTnT5YOwAHwiAW9aI1P86AChKAY6X7QTFMPdtU9EOd3Eal7K
9GN2HbFyVljtCU876GoJ1GaSyMv4f/ddy6TVdS1rMjiCT+KPIRzU1kzD3k4C1lIN
/17OCdwnOmgiv+2tAHaQJMaczojSBLsQ5E2hey+2Bm8BOmTw65ezzPxgYCFY+Veo
xmppAgbD3kUZiZU0c7o4sfELg+qXcRydn5WKaj9ltmUtr2PKzP8SJNbuQihpHXuL
uEPSrvd8eun29806+cshETrBbBSI2KwhP8aRIzHMqOBQ1QvdKcMUls8pNRPhETHz
KCkTkKWMM7C+nG6Gn7fD6PjEFC26qId5qfIzMEqgGJ/1g22HPZknTCcpTvDnOKNK
QjGjdDynCQ12kYdbKFzjmQSg+QI/JjhGUtfMlPqdsmZu2z0IICk2qdV7KjN8AWQW
Mir/ZjfaxJ0qWaX/Kri+PpnxvLqIl2tq8W0P1lS5NSmXQQeaCVlorWfZbG7S9vCC
CAD5QVwMQbRg9fp60omTlpxE0sFcqkuBhoChpryx5uBbiXS9CN0CA0R24QJ6wDrP
Cv1JjV2axX74NWdHKlxoOzVjFQ3z+DL9ZUK+qBJltz2Qm+fbZt6gsRHWWFLSzMf7
kkGevwVVaEck5RyblzZLo5ZdjV128lMue4wq0ssCvUGucjnPN2bfqNyUqnXdRMn6
56zo2D4xxoc3xCcXlwEX6Ztla7iIB2Ej2US1t2LMUJPwwRNosycnDumlkBeoXhzS
mbYrO9vKl3zFdsErVsWuIyvl+2S21TiR+rELoO6HWDlXjkYWgKiDPygcr5cEUd6t
zNg8smbkMwQYS4ljefqwx8YLaErjuBXNECG8mvS2BJkxs7ucvsZSA6SAdia8O1TB
wQWGSc+xhFHGsITUNJVN6d2E1Pj+B9qPoVSR+dm4AoVsodxfyh8or0vw4G4q4UoU
ApPvSwI9g7URZUc7F3odWOZBNOBpVo3gBc18W1EtavEPXckZKhYiytakdGl/sCdO
Lxhuj6lB+Q9/oTzQRAObfNybGxmV47OJxBtCt9dyBW/3kYPymSoFhIN4DyQ0m8er
siHG5LkWfr1vLNMz36Q3QxebrQ/mt23ezNuuJqALy2JgrTFpOTbdtcoowjlXDDHY
nuy7c7x0CFA1tP1oQGPcc5O0XJ6eLaXzlLGbVKng2TCUaySgypCZeplk1tMgFKL5
cMbyytJWxHhrz+0H8AE/4yAI9X19CCkYLsgbrZar1MRHChfCM5TQoY+WO7SylJKJ
qnKgSEJmEQQmQKEpXLziVDRWwaPIuWen0Yh3nrPz1qphLNYRa2n4SlvU3MegqUZ2
S5QECxNO+GR7VgDaHHrw6q6R9x3zy91FojTxakfim96xlCyFH7WC/JrWdMjD0DCL
jMo3aE6bGMKquDxH42f8I76+NeOblCPudGGZXNZLyWaop9fObBLuVygk5h/AyTp5
TGCILxd11ZFzcK1sEoD6x1uW2GHDCFe8EihfmFWYKFGsl1Ee8LU1iRvA10Ky+nRV
IbLM1qaw4qRATQfsZgGSs8MilEqAZnbAbhd1SEtjguyezM4RwDPSxo5q6p2U4UTK
EWbR4fDaaZKmUEPeWDopArwagK8PoantkThomTsoyNUnSURKhUQGjkac4ZVqJIF0
q4+D63DBtmk2qbCsTyPeQVT5uJjfo0DzkkmKrpma4f40pSX4r+2tQWBcnwyNSoGQ
XrxemT2pR/ik/PJGZAUK1eq7CZSqTbgOfpEfPrbsANeINP9rYQOOLenIxY/yCciQ
a2Mo2R/UgEpZvDN5ioMOHs/+RfRidDMdKAsqBsuydkIDM4k63OY3x2/pJNWU9REM
mF2NdSMs/CDMQ/rZtKwOii4xjvkvc3txTL2Y0hAfSMuvqpcDqrmONFlcSPXQFDd4
VVzzYQCCeo3HN4Np+kb6fDy06Hgm31NwD5Ek7HfxqoEyVHtIcaE8PA+cW9XLqIlL
9BmW+oCITp/UdJ0MYK2idIjxhafTVqIAUFm/oqLhSCT7lf640Bn9K02sBX25sHin
fF1RneOAZ2gA853us6uu6lBmuIV4D/bC1Iav/ipOmd4GCHZHZsaCpUeXHGbqddve
MgK3XZWLL98pRfKJEHIDXNxIDII91CMfjzVbq9FyH8i8vZ45PTsdy92yDKsYFmjE
Yo+mbaGFReceFBw/tpkyE/3YM4Bi5Oxg6ghdwhDMlyCiTfHRCRP1UTuGar+Sj15J
5rqo2UsoTsX+e4nGP8e8EDs0rekauZBrFiJ3AAqEM8nrfUTiTJ4U1I6YxYO2W3Np
UC9bEQLLVM8GD60lwVECbUuZm/EwebtysiK/wlyhP/oyyCPsrkZbgvSwVCFQOxpl
6WQXwjTe0OSlLkeO0nw+fu4DJm5g8R2oqESOReqg/8++VRteHJ22yoDIiXMU44yU
nF7+QoJG7BfPZgX7G+Um3er2TJT9bhEBar8wG7e2mk3qt7NfA9j+/OCBm6MgpQ9Q
ADzpiOqAeZ7gqI+ospGGH9gG96uoVhEgY67UOKqTrsot3RHcJil8uXsgm57vziIH
2gGa4dHqdCy6FRonWus0IamyYLZGhKbcoK28wgo7d6o3DDhCISVgF5Cl3oF88kWy
YQNjU/+/Ekv8t0tAM1RZM0ZBo+3VJ34alr+LV8B1JzPR3hUf9s7ilWjPdS7pKR1E
jB2R/iYErjk0PnzsSz/3oJhRjbpK8GAAjul5urOpco7mcwR5o2DvbsgvLe790VKw
VWc/QzStkuxABJTceGjm5pAAlqC7a+Bmj1fIMyTAtGZYe8tiB/F4jTpIjqGxIOSF
NtERmy9LUe3ozm5Gd2Bm4iBjV1xeUbuc6kSZkOXEymBrLY7HxMVieQE5BflzFeu3
zgg7/Nmm86UyjvOXYGAdCpd0WSubvk038KhoNNvtHv/xYxpgcvFCvLCEAiPqZ6vx
lWKOZrB6pobHVN4TBsiFTy/YnYfrEJfEW+c9MyyFl1FbOxB/2+ie65SaaWC9cp1C
9x/h9+aaYGE4N+pQ1hD6jsGvv+x9NQ+iv4GedXy3AHaFc7rcXLoYoZR48R/zW3OH
ARbp4arQdfHKdd9UUl+RvCznX/e5hp1yGaYQAYdX5RNwy9ATi/u+3hnRUyiKiYzt
NIRH53vXdDtlUrlpNZ5RcHYBbJ/Vqufg14bFl4Svmc2aCRv5y4+qMOmZQGnYin9n
V493FGjVTlyWZceYKF3cIkzmpOziIhjApPPnkX45xBoLAJpnJukL/QEQiCjvFLl/
l4THKCtKOXmL9Ayz4F8Jj6NiQplXJ+pQXh7P7GvfQmp49z06DW9xRC4BbkRcKRGh
uXeHkbnULGexj7d0rdKJ4RbM38DVve6YQyP6wnJl8FCy/eK/jOI+quGBvgnzRJjc
+6WuXBH8tz7wNbJy6CSIAAveNPJlsG4i9AlQgLlktNaHKLeeiGl6d058HnCfKjWv
6h6LvILjWwjC7W0fnXF1akJj7GSLdsJKcnsiaQ6t7Y5qxA4LHTc3cyDLps0oSAtU
KNUyEYT2qHJn1dpcYoC/mV49giT/nlwdXznQFeUiQbkRXi9kT+NBILhzJNMePBMV
rO6zlC0g1SWtlnMXl/FFgo6FD+pSZjaKv5e97qVWTQaLI8Qo8G/Z0ULbvcZuqU10
aZ+Kk4SwswZ5wotH7qo6NW5w7td6Cx5YXz8R622Ym5eD7Wok6PLzmoOSnr40rA7r
a4To+HzZ6jF7vLrxdLTTrNr7z5T28jOgJm+00Se9s7F5YmpupZBZtoqGbHxgTGjb
jjElnVk1WWkeYZQQp/BERBKDUKLDaN1ifxtPHfVDuQAL6jU/wGGaVbbEQDG7rgby
GMycSa6HP+WsX/efAa1RH3LQf7gdCEUxSHsivaFfLywkbH3a6HBap7NRKWu0H61O
Q/s5wKE0dko1NlLyg6KCPuwRHoytJmoC3lMG9VFiBPnFWvxuJx6BOiM5swwtzeHy
B3rXcc7c8icVO8u2pqA2zocwCARpLVs6Szia21jMNjqTWFlvb8LVNDLAxOyFgkGM
wcp7AAiZxmlhm7pJXJRoG4iWeemx8dVtAuS8O21d0h4WdVXpudrVPyZfeXoQguec
aALbbW8QaziUWO+KCN+krLTM37WM/64AnxN9SrU0aaEqSoxFrhxDLJsG+Gga086Y
TXHO5GINaHul5E63E+uXNHQgfpDAtGpqR9DIJCZ3uRS5C9NhgWTkbx0RQQOhVNIh
AKlZZFnUzEIxgqf0UGakpvot5YJKUFPWwWt/lxXj5QX01URcQAfeAl/UbiSqFCpN
h5wFaq2CqAfRcLzXwIdIS34iqAvOF0NKqa7Ecwz3x3Jz4kzvT1jhRWhTbN9BrIbm
eFTBTXRxEL3gg+3j8BunvXs9uAs38d3D13MnOQPG0BRRlzpp9Y0SzkoNxWFe2gQb
YqSv0nHQpNPVSGo5tMP2J4zOSQzWqmTI5rATBv2F820vRtn3/h4AEyDBHe752Cay
I4AK5SpRXT5dmxOX2JNLxtgFYya3PF0HrwdUHL573Y+zMR+QAUq1VnLKiB4R/sv4
AowWwrhKrw8uYbYKw8VFUP4EyOpbDjZWyw8tVzz1+8AfBlQ0b97+Pvjd829DN6mc
uHUq40+oAw3wSD+n4Mc0owc67Tq2Iti5nvLd5nwlAK7VykogPOUQ3F526PuSoifQ
gp79hQBlaG8+1AGqN805Q9i4bzSF0FwPH73QZ+KzbFWzTdb2LorfwyQz1WjqEtOS
i6vNvDyvDA3Nebh1ZsVeNUpWiBvpsS0FADw9HylUwc3mUqvs9mq5Hf5ps5qOhWd6
BG+wmJEXXFXyAVnw2+mS/m6RvgvI0S1V+nZ6tZ1K3SSjF8ScAbW2tqrW+D5ONACK
m3XXZLXzmLOG6KwNiU6VdNIDsMRY3DL8jLQkPtbU2wHsRrNlS5GvqbTOaoQVdY/S
WY1JE9v+T7za8T2MlXhwYm1LAW9Zmruqx8gU+7TfFdkSzGlI4GPOxFRdt6u5+VV5
K3IJR5UBm2zDjf9Dvc8VJPKb2OdB0bDjEBOWj1/+sZr2Oo0xlKUKJTpYijuwl0SS
67ke1aHOVn0SoTJfCgJWjc8CTUQfX6JZC7DZSjUWAJ3LA5gyu3WL3x0KhELPYhee
wogdGSi2QQblEundEbUXy9sINbtyy0ROwd1U3PuFSdLOi1NT7wPk0/uA90UT2pwD
gzeoSJoWKOnNIea2f2Qr8QMhSaCFrEM+09BjyNaO2MLxOqkYgqhKhKbEfBmg89ju
AIM1eO2v5vB2pfvCck8NFTuT62gq2vmBTN2NW6jGZcn7qqpUhs6k7bsB5ejN3ky5
0CfE6Ft7/w+ie8VR8t0q+32LAkjGNmhdO0vTNdKkPHt6dph0/NssOrSTA++F5xaQ
WTRNwWbmctbuOKcSIr+OxEXINgnurPyFz4mzbok5duXipZMSd7+Jfp7sTK17G8qP
QtrUA15Uk9D/hLfCh2/y7OLjAqNbTf7q8pF0IJGlLk7PLBwv6ffK0UirSMW+1BYl
tuvAXoTDrhTuh23v7slR2AVaPVejKlwqlEUc4JkNfpi7ZZJUmfOj+S4e5rR875ZT
+Kr9TfpLeHN29KFq2ethTytHDAyXe6ge8soMiQAIVDEDnTHcVfvRXC8fqcv9rYNx
B2QZY8dJix4h28jEDzPB2irpPpmEx8FrVtmWAQGO94428dh9MvpDZozZ7y7rO62h
qY25HG1UTrN+ph4N1o2s7KKmr6ojij9DoEhrKJwck/53oWkvIMYAG/DoBlO9SyXQ
A3apFA1l6zBU+ppgZRIjonJIjlaMlMtWYnyHWZGZSexJgsGPc1aFTjh+7FqTydQC
wrNLGZdl8j+U/dMEIvDNddd0Rv2AcWOVQZcJsgkxlmGIJN6I5mo8zQIfwXjwdV4E
GG4HnMxW/F1A5x/Mm6caXbVTvJHCpcOfJH+pdTS/JkmLx2nhxNKOhtBl/WBVK2tQ
1gcs63dz1xUxSTBJe+AB1kIMb7NO5EFz2CVOa72EOWn1xqdM1IpNfffwQI6cwthu
SbzuiAFAHp+i4asp1BdTm4D78hNWL0/wL8WTgnUfnfei+E4aycHMTQxPQ5EU+2UX
7C9x9u9UmlJcCn0RhcbH8pN7jS1GATgwqfdRJBvHerwH1qFLRI1wMrvh8pyAF+H0
82hKsIJejCBWrzqQRuFh3F68q2MQqO2BjFemcfH5sKXEtfNP7iNCwyLMnyJoQoTF
Vwoi4G9bqmmvi+axAogG893NwIYtjokEPK7NU6ZnL3VeNJ2niVJ/44A8ucwkI5xQ
2aDY2ozJsl5Vbly3/jAqppEfRMxHb9SkVZcN7qD9ou0pL8RQjHljqlX0tDjvT8aU
cyrJnqr9Dx6JKKKp5Q010XZ9pDKufmCeJaAyYZzDWb+U51VXMC8y7X63xIF3+O+8
DEr9fwSmQ7t7HDjwGbiybk4OGZDWILRxWbvfi6Om6CSvEH2jpz4mLq0jmNfYa/vW
Nsas0e3PxGSvwaV0m+5DUGkUlQHdlexubgfESrbXe2/9OeZ4n/pods1Ql1GWDEoX
zvNb423MqWp8oDfBZt6LHEyXCg6LpG8yUD1En0DaV+cH3ylI3JptJe1EfxDvxCfz
klQf6Qy9nlR/u9PC5MRjJrV2ZzcHDKANEmC7R2uRKMQfkIJ+VzK3CkQTRRtUvVVp
PMV40kJyH+tEf926QhlSPV3it1a5jnjBjQqnHO+TA8RPOK42fpyZLxbW5LnC47bT
P1IeBvW+OxcwITyfHIbFcU8ryzPicBEzAjjSnzRiuFZI6kE05FqnRUzUj2bksKbO
7sVBbtBsGMAjagHxxR0HSy8W0/ede26GwFeVZduGCJZbSqovWjvRc+el2A9gHJR6
dNOyB8pOE+RteCbdywMPxMAcs4+7O20G/wILf6BwXFh9/irQqx3Fpq2sr/eLp4sZ
7PcM59dkDgnJeM8SMD0eyQM1QA4Q+y3RZR8vy9Gf+r9XBeiqsFFtBxyFKfmWq+AN
dcbLUrr8VYU0DBafjSvKMjgbV9b9SWkpNCWb5WOhxFVb2sD3JhC0rXeNVbAu6RHV
RDxJxOzLJU1vOQ3S05llgkYmfD6zcwhDbvWU5QfpkhnBHlzSwkFuh8Mw615/naIi
6+EjeH4uVvDQJQRijzGmc8wnIO0xxnO5zx1rF6q3CQQxPoZlVgmo7s8UCMC7xeEp
NgRLAgz0O18cqwir/k+zrjD6W0+oOun1TB1cBq5I7S1ociwJtoW2SVJR4yFpwJ5m
gV5ehSJDdsvXnCXm6QLpQ2M0jq7Mrdp9NFW8Z21Z9n0LZ9sZGJtwhFOeDRHCjJnS
xE4T3iEkCjKFQjqvdR1NPqb6kByn92vzgJdfSdnSyLTen8lE+tsO0ja4cR11SA4L
YHqgumpoXWSPj09jiiN7kRQQjWp1Dvj9I+hDzh2QTxjiaTX5XypvAz3cZL8DQyKO
eq71SAfK+BS210U0fMRldW+yC3YJ9RUKDek3++r8bH+gWC6kcnBr549iNCILef4m
JIhpDIVeklHZ7/yDaUqXZyBuNPf9VgPClZCWP0TiUN02VD1EUHaTfY7xwumVTQw9
btBhigseIAHxIB+9YpaxtcB7IzoVYF3/JpwF71el1Rc920K63WP0UGfesmu53Xo0
JSMTy5ay6xo3oNO8h3qgNQF8Qgsg7y3nbELCg7I39v6AMxEMwnbZ08XczcFBU7Ko
/d33Pt7UAC5i5OjqdqPo7tqIja/cAgK0zS7OA12xpe5Jiv9wQV+9Qjk6jAJwrSkO
vHvHV6jTiUqSdpnU8cziuxmrPN7uSFos2qpJvTsnrJltuBAmu7bmQv3cC5cWJxiC
xiKoX7rFP4dr5d0YuYGTdhBLqNyqIP3pO0Udyi/1yKwIF6DDvV7o+sKI9+ielyyS
hPUmT9/ld6faRmnS+rru5oI9D9YSulnIG3NUvfOushEXhEGVjo4jZzGqZIKUWbbW
E5nCV75ofZHWnDaFwhi4UOEWHhmysK40QbJuJGGvjoYNCxvkMeIFLruLXPXoK/50
aemN6HP5c2zOXKL+MouGIaXXZTSF9kiNx3zhzGybXug74VIqwqLODDbAxm7UMsjI
s+1ehdLLcvz/HTiVoNpt9ftmDsK9DD5wQbVV4MyAsHH0Tk0pmgI21FUWT9Vb+eNo
Mk29Gag1J2sKmCTpHRj4MxWolVaw3GjPHwt6jIS+vFfjJdjkRrzyPeXxGVM0/b9Z
LA9/uXmIl5N7wxIgnH7pKo2btAST9KMtNSsrZda1tL+3v+DuUlpb+zIEEXen956L
FhtKeDxBvQ/Cy0AlmszDeuECF2ERphlfhwrzYfdFYT9L8oRRIWh7zcpOpEpZDnqS
sxlHEd7Uur3TXntghLyU3vXHTUg4V6kueMnwRAA4Ar7pYymVXBNpn7dqWwmnUkJ0
clilSaaw2E1N9jF6CLO3FU8bBtpfCQ7qLyQ24JdBaDqpVJkfMWiA4wZAAlH5z3lZ
aXAyREV6Y6w5QvWpOZ4eWT+EqOuGRn3qWpFO/F9mJpn/q6MKteQXtSLB0DR8a+tR
Ux6e5z7CQN5wd0qifFuCr3l0llU4fedlQac+emARdxZLtZXRQsmIowasx/NqJwG+
y7UIgO6+hqp1Zgl5KUKfh/V9It/dhZNM7aSt8ywz5v2FSDFK9tRTCGUcvT8RDx6l
o38Ai3KEFg7KSq4xvMrnzJaHSx2qCCQrLMOdLbF9egkB0bdXl3jXLUnDlIc0hXPS
GvkKWs5PjXcSS2gMkuqIjkfgmdKb9NwBRFF5GuIUS63Nh/FPJ3UnqhykyycUXBYJ
RRLkdA0+cge1Z45HpJJko3l9dXcNeSjJshTUah4Dp4jTNwJqLQFGh1vrPR99Yu3v
lEqi3Hm8vjM831xd6JQRCeuYBN8U4aceq+gf86+luHMD4RUbtO9bKFOHG3mr+02o
spdHjOYEWZVUeurwoQB/J24+heKmonW4xUhzTpPtz7cyPy6C+ow8H/GE9vie1xYE
qa1WagArej5I3WEZc9SRdJDF/lNMqe0ngWfJzdKLzhESEi2seTo4iAdH8maDrDel
v5JgUsk4yb6GjiuE1tTCpEFuIWk3vMYlZ3dUsgo2QgNMIcWW2zO1xGpFWWUPjfAc
A6ERxFFIEEiRm5I0s4saxL452vceuaXUciDvyWYZpSfFpLfKJkyFlDAGADWj5DY0
R3L36Bfrmxyzbr3w0uCIyfsHJChzLdbEpir/KMPxEbULQ5s95WKT/MHIYycblItT
sqnGcGIkI5HgQjf3z+q49AtBW9BtvxqC2Y8/7ey0QU4Q9xYHWqjzD0p1eAiLgkyE
B/0ajo6FDWlrwVsDNQ0COStBIH8v4U8mgzKyQB6zqUNPXT7JNOOI4n0boB+GiKVT
GigWc4mdGi6ao3gUDVWaBTn75jTtdK19oRDFMpEgTsN49vwUbcLNgcmFEKIlQ3R5
LZF0dW5NfmbehQbdYG0voqJ583AjkQ2/CgNv74wD60FhK+5r0iyHv5NKjn4geZa9
r+6U7kCPOtg6MSva7MMY//SP78TPlB7Z7U6LQuUqdOwpA82oI/89KA2atDNOzq7n
rZoW/rYnslNAODB5EJfsQHUJn5TZL+m1JXoWCNv+dmScJ/azpG79TgTXvy2ed106
+W+wiGjaGui+8EeVl9AjgCDRRBupgzRPACjfBQLF34Lvlxfzyb9rD7tzC5LQbd8e
GXf4QMU4gUdC8O1vZTeK6gU2d3tRl8jFFIopirMn5BEqmWtJvv4TcAVNOWF9XaGG
tDxOJYuUyKFZUf51Sgbw1iS3qoXwuL2OiAjCiAHE2QmHXgyOSIdIEIxt4GdGMVLF
fWMfSBs+WBVJ1v932VTz0giwELfG3lPyYEltUPoVTEDXkAe9AsaLPvNq5957spo1
vyq1UmOX6Og86cyAMC7BU47LYewSWp1Nvu50rKzpZYMjtnrSvR/dzJuinj0Gxqyq
zY2JwbtkhmXsalm/UB/88QPMOOdg5noY1gmgheMJ4BiCgpNmvQfI8U1Web//srD8
fKsXX2yRv2evt5bjWboW9WgALtbj2TcsTq15SdHa4RkD4JWhafrh2FBqQwR9w/kS
O5BHmjmO3J8bv4ty+MO9gU7/Gazox4tKPAPYORHMIOONqoau9skL0GT/3dZw7xNO
665FYSKVCOV6XeW8XM7xs/0rfc7G+YRjWiJKYdtugfkqv3JeoO6KF8Mp7k0OhSD5
efTAfb67xxO3ky3nQ+VSM37F8MFBRK0JYelkE9pOB2SgxHEIZGEOPp27WX/EhxIr
+vD/fnWlre5wC/XwtOymEHymKO6SaMomekbffRuFbDv00TcSeqFo4MI9jWgd60G/
+JSXIofjTVfLSM1hoHJTrI8KMl5ga3szt28oYkP/80dlds8CcouEeo+Jovyy63xy
BCHoSmCdpFZIYAjKnAs4zXRfIzoPWP1twuBOsCNwENXBKlKVLUd/Uk5rSgRcuuO+
fEM6NZmSgfS1Fe1ADm9gDEjQOvVPIGRD61djkFkCdmUy+R2vN/sbBRGLE0afyYWM
dWRNpHbnpFQoofbU1L5uUy5skctu0hD/QErco2XkqBD5TuhpEw+NXJ8eRcWN1bj+
3zWNWTgqKEmhcqM/rjRmnjuYs+6FkCohAYv8CeL/OGJAe4BfD8TrMv6VqIbfj20a
EfFIEVmGf8DkhLzwrih+TkXg0+kykG8RaVvjwu8iVIB0v0mBxDbnUKcrJM1xGnq1
IlpnakdQkOnh/hFkEO8iJMjlWIN/UvZ4KfRwJxgW4TvQtB2TZPACEIId5BhTrodI
2vC82L37ruxO6qpxg47DuKxBJDJyHicF8efIQe3HIdZQqxzEsZVhbLzhoaePCdWX
k0ORFs22kms3KX8kvM3uRVtoau5n1iduG9Ah0gmvJdwBu+MXJYDKxnfFFrQOjQuA
/rtQ5KeUXZ5PN/wyEuQ06IGa9r+Hp65PAe7Vvg0xzjmxLgG4571WkwzacEwsMkyb
OOJXOKGB6+hmVhvM7GMfzgCOikJEyzogqs8qEc+uk+vtKYM8+ZrKwUjdytUtvdur
G4C7gn6WowkQg6PJtE61J7hplTELjs+pURRHwxBfQhUvA9ytaRVUTgP7WgYja08G
RP8Xjo+BeQkjsaxxd1qj9x6OmEJ/iLZfcLcn7uW2rNwbr6ZizgQyORleXZL9HTYl
70iT9NV5d1VhWKZIUPBFhRNAj6n9FqrH0A233FcgspofQdErr0WVL+0D+60Cyr5V
O4T/A6hSPbR7X9juOVgpnmEeq+0GsyFo8Xf48uzCn72tC/0mFQWN+2jhWE3q8NVP
CqgTaTksFWYDOmSgHrj+9h2An2DdhoqDMcHhUaeUyUf9OYPztKJjqcz1Z6QIeYrs
x6o6uZEyTVRS/a0Vz8od561FfttF/CJYrXeFXAZo1vYq9qlye72qnfF0urOmxDet
aIuSwCxKbihTCuCigOychPXKnHSXCx9cbbqS1G+vzEsbtYThUULt1Q1E0gb95Vg7
BQNUIc8dfv+Ccq/OpPz14jc4gxZm+ENfp11EORfPUrg3FJR79eOmgnMWtPHX2BWn
CCCGPbyFyH4od9Q6d+lQsR0sfXuyA1FhA4rR3FqnoGDIs4cnJC2i1GshFME9BqlC
4kJt4KR3zd/ZlEBexOFWQW0WCc0gG6Y3ibHQLMMgimGYRjIDPSV+GYrZg+jB64nl
Amgvzhfyua0Ga9Vdin/E/VfHMyZnFauy4Jn7TQK3w7p/qTU+gMqynHeHGjGgB9U/
CuD70d1WHHufrMu7wluaW6GlQAXmEZHq4tEjsPiodY2Yvzkwt3y3FXwLxL234hd2
1erx9FHonS6mi9akrQIpaujp5bdnVhMyLITFUSSZGPhN2QkvWLP6nkX1TvdmT4B2
OZ6SfFDhLiV4GOxVqR6NGfnSOFVg70FZkqY5wLs5sFZt17CT1pOTlh98sEoEpDoI
htBSBBxl70yzWHhX0+HtmbQihJCFqeZvKFvq28KwocUsufDsP5vt/s7r7HnnGe/B
kZFZUpmhOb1uQVCj7+KcqZ9VB57jkRXHJWJb2GsE+oF1YRovZzcYa+tasY00jPwe
piJZbcBtJotl7ztQzYuMtn7wkIIWAIk/0VpYTkaPrgfVsOmIimUmvJ4a8SWNOCX+
PKUE5WiuNdyM5xGJe2IvLpW8azAFOPL07iVqfWK3Hdk4aO0q7ZsavH2uimg85BzT
KcWTuRnhVA3JYPDp4H15xel3YRs2W8SV2BIx40SpyqK4xtUJEWaQimKzPWVOfvIC
+0uk/xLx7CxNcpt3LmpZy+lTpMMH5tRMTKJF71psV7Jt6Fc+3NqCEbpSAZXQxPGS
1z/0eNaqJvwQnQjrWyxjQC9BgaKaxdtnMqYkvCPao/qk+xLweXKyO7Kn/e9ufnU6
FWspmSNjT6PcjKh/QRQq/7SPuLUtAZhk3WhD3OZ7BnyqRBe23159z7r/nQ2lka4j
Hp4X4KSyA1Y4TGg+iaKHxPHPeVyQd1MqBJ+4Osbu11UJmKyo7iENO7UsJ8dI5Ou/
XHdfn4os6MZ7Db6T9YYjAdSXPMIJnzauTLDwBbbIzr1bCChzMKGKwlYhPwU/0akc
Y8n1AE678b8qEBG4xj7tw5vlXqCePPr69vTnmUlqHoBI2Ymx2UCHZJVBIN6R7v9Q
PW9RvCPLtS/NR2b87EcxwDP2IwfAYLiHdM7LCY1oQJhX3wSHRJZoS8pcWBCRfg6y
7H/9CWlX1fTwvqLuXG18bEYM9BlS30HJrqYYTl8mw6PncNVLytFYTWoFJzKYGpnq
FY05z5XGAJ7AdwApWLLqeWSsxSA62xwYOR7IozMWXpp7zJUYFuCF2Iwe/Q1m9eip
g6BzaAh3G29rpoHHC0n1SyAnYKSC309KNCJqta58CSkwKORPELWdAceMF3a+RJ5V
Fbj+6b6eBnde0ICdm6XO59auDsUhXf2S/LVeiCdmF+9F3/BVxjXeWM050ptlDYBB
rZkCAT5mdlgsvGhJzeYgr7NHgvW0LVr8OsUtOjzmUSP8Sx4enDhGFB/jV1clI2pW
m0OS30kgsFFhyh8ziSogv4ISqTZzDgZh2MvAi858OP8Cu3stYMMZWaWomM3sBYUD
rXaO9s5hNyXfXXSsJJ5DscI2G8PIZW1qS6ZRgY9VhIFthM4T1WNOlK+2rFm+S0+7
P+0bs6kOq5AEm1yu1a5QH7I//JDFtI0UIPSYU0DgbuO003HpnNYtgUw8rIuvsHpU
4VMHhefW0ak/GtxHH7qNFFuM8qPo3XvFa1VZAG6Btpb4+chwLncwmeudCCnliMa0
oQYEDrAWMLorH4GpXQxSPdk0uqEv2t6lqtSHELUA0N4W4n+eRy2tMa7T2GQmTumR
7wm2nFrN67FwMYM5xnAEYavvN/B5TvmzoYF2IVaWPe5bwsk1+kbOWNGMKcNZ2gMi
TmK9ylP5GO3VGwUJEQIJgAw/Aakb3yYVsp8rABdXMB634t9mVscmIoX2er8zn4xJ
NVh1cI2rxiQZgggdiP86xnmQImLyObxo6wywSzLvrMKcm0ohOevZmpd3mWe1eGEa
TEAmPidTkVN00JMEFJJHU4sMQMaxpZNVvgOIXpbXt5ya3RNkL7/kyBckOJQN2nfL
copBWHOVA3ARAF3Ci4DnJlMwyMkKPQQCxtDvycGqm9EJbqv1lF6MhGbybHghU+Tr
uVXPPac3/+1QYPwI9M6IpMYobqJEITpG1NGIXic0UrlphblOVAAPNROmjFEdaylp
L88OJySaYWECDQqlK3igBCfYhDrK7m4lvZX01rlwowZkV0oaZ3N/zT5Cpks9bk5p
vRVfZTj3PE0hyHB0Qi2fPFdlD+tidoeGTAXNEoTWncETE6/S5jJ04QN4eakS4A0X
MIlc6efSJYrbUB3f9zUmj7iijHn3MbgvLM/Xt2eUJtelNhQ5mNkVIoJ/7seiPuH+
aLUs97ftGTEIzthLRqC6AR8NEiXEHzmFaRIB4/XJbmXC9FoMo6rPxsl/uDpHIDNe
nznxzidNbR8mrn6Cfmp30R80iXbjQGo/ZUIa42is4e62L1MOgND8HPh5Mq6nm0RR
FhiCEpr2G3xJwr3991HIBxbG2NePyDKWSDkHP8LTJxqTBjA/C79aVr8HiJXfZVFU
97EcCaePOpF152xXDByvfNLXkOXSuh8XE49RixIkQVewcgThIrZq+d8bPFbBq/1O
vYd4+GxZIH/qw9woaGZhqhHpq1qX1JrAWTaQ48AE8fix/NAKzn6Xp9U31BJPSKoY
2PmiwaP/JosPTRclk58cw2V1EfPEFpFBFkWnjbj+i7EELg/fIbz01jQkObqGrWGe
O34nfnxZ44SQTZderqJcQGDh34G6uLI2iTV3S1YqdZdPfLu58Zri009PttJxMz56
Mq2Hn8kHkqLVrhv/uz5izP6GxUlnNrB8+a+65MzwYEjHK74gL5VOqzDIEhAy9YA0
XS8aEsGvZjGCRI/jbh8l+ktjyW4MFOQI3tabx4B5ojZ6++h0FBvGSdU5BOyNDMJf
gcuTh+OU2I3f5dloXEFr/KZYfov9SSlZ16qpj44dgOdmKyy4uJ1XKXSOUsVZXMi8
DN/anHHLQ5lGtkXYDx4MwvhKPpypUT8JTUCX4vs8eBA13upw80rpiXzpWhWPjG3t
xzasP0uRYcconalNAi1uTJbOQD5iPNLXLM5Upioy90HsSNRe4WoDJurAgl7biSkq
tPEvRxAhDEfa52SQabOkGsENOJ+pleCsY0XcRkkgp+or0lgPLaq+QLvAEMn6Y9ND
KYl9GPkDxmmrOzxv5RmAq5UtIzke4d9xIViSJlux/5QFVPHKv124wjOKumMzPV6r
sho0FOHlnkzsQ9qf3OwhEaXhooeFiWyFPOvkmX+yfJ98xNjWZi8jFPcsuSzbI6HY
GAvwnRycltmd0ugO9wDYNdTOy35dQ+a3j/wfHryN5GPYbyCfqv5vMHOp9fVVpm3V
vclaBQttVEJQnWsPNM6el8i3geyvIejyLHJZLflouYK7CrRb0xAOdbdTiZKeJ2P6
276eWFrhwnIZuN+VsEdhqz2XpOCy9bTbZlPbccn3fYNUgNZ2JoOfqP2Qp8zB2qsQ
LUTXuV7Nb/6dt9vBhPIqBaqP/XFUnH3weZTvpP2QuVxQSbu3EUlspUbRU3Ea/ijm
0SuQc4RZh+iwFPxSu79AYGNgiGdCb1LrMLE/UJS3+PCQl52CVKbfkgmdN7mgeP/D
RVaROKFef4Gb89YPNXZnUewfjL7KyjQJ6l7jE3MXhgS4HMUFpmCGrkCLWC8g2vQn
g38iM0e1eUpTczkIiR53dNguZXl1VmH5DN1P8qOVpD0caP2EaDGvhm5hRA3F0Nqx
u+rmTiowx54pgPeyBsdQb297VIUF4lN8ziYqJx9+ZA/AA/ZZJ13JNDNN3S1GB37/
d+ExmGPdEp3oxFb7T4r3D6IyyWGwsq0g1Qm/0DzuJX/GbORSLNarV5QDhrTwDP3G
7gHRgunsya45f/7V0FgfiqMU3vVJfFT9PjkdYpJ9eexxLJUPf4VMaluUx/IPTc1G
0Y3HWXpksZp0J4PSYIJJ6GBgfi6zN/OztZCCldsqBBUTMvsAqKZOjuCu992PVXv3
dxeZsGhR6A5DRgQRLz1lJA/fDj38IZqZPjNz0nV1AgmBjpHnZIw/ODVf7HRZkF27
aaa4eqA5LsRHmrrxdaRU5PYl8oOSmDaZjjWXEB0WChIjXfJ6pR4dW3ACdqwUoR0W
eWApZau7ueSp+5bXEY/xea9t+RZ8JV52Sun15JzHFnUzT2W2FvrmM8sTD7SzDLU+
o3MrQlc00PnlzHbH7PEOSaLWaf2pcF73aXDNUMiQEIRBgztaO3ju+spEPr1bnRGV
jwhsWM1ixA+5cO7LBkO+5rVv/F4dTcgF4uH17sUSIfkmu5s4SqQ7NCTiFbEAeHCh
aevOFMTAXc7xpM2qniiIexA/qRMtPt7/JWHeh8D92DIbAU1hQH2AMbP1kb1XTivd
i3N/I6NFTRrDZWjdO0ZyXkJY9EONmaxLRjKYTUm+OogkfT0yGbHy97lj0LMBPZVZ
4b9V7qqRUxYGSjc866ZVE5BGah376pN/E5gPnAKlQ5MK3/CROoQdecfXoPsblhma
rCW27kcsaT0hgLZPO95KvijDeYNmMawfJz15B4AfbI80Sz0eHOjkFjtzJy032ZBc
00VBhbbj51VcdHdKKoLfW46WPQt31SA4T7yqKObKprCMK8NjSJlVfGJCNMQJbvba
OzTkNPS6xJeMXFWIMRyqmpthe5jFW+757ye4v8go5v8NhVeSVO9rBeZC9GRMeq8t
LISfu97i4pZWpqo751T7aWOHDDxqFCtK3x2ywTupSB0xzrSGvEHKjQadJcSXENrn
zVZyq01rq/LgBhdSEykfp6fgfnyvLvVWI5P8vawZpbs+0FwJiSU0kS7NdWN37wYt
tITTw+VTJEPtqcGIlipYR5N4nNh4hBlKHFNN9Lef7fzNiO3Na8RAhlejPNhd0aFX
979ndDgpHObnnA2yxZnOWkq8iM10aHFL9+vfWriAhuAdcDnoL14HCvnmphWULcXE
orJHE6s+oVz0hoob3DsjY3RJsJ9X9H9tLJvux3qEzpo5/zymDs6tq4vmKQAfLo5J
w8KtoLe6DufotyvvRwOt43Om5C8pQv+tMfK4XNyflfqp6JnrAdR8RKXuwPJCEL9d
gQ46QXAejpo7DrBZP1mFu2sAHiiqsJYC6+LFLmr/taTaKmYxLS0xclzexHvF8oiG
rcs+8rIehCwlOJs8JrBZdUwiM4xVGhcUl4dcdcz2wQTqN0hsl62ffj0JG6VedklM
Mg6zgDDss9PrpRsmX1Zg39D6tKxGb5GNRhHGQRHKRlmb8eBDWKQ9gQwL+3FXmDwF
D5Nq2PgRvShN34PRI2ePpiLi3sFUyS4e6Tc0s1dhvhwcG8hpkJEsqYGtWufIdufl
yuO9rTlQfSYMA7DVhfqzCQOrYgQh2XBXaLezKjitZhzGANw4WbJbmjq8t8Hbk36X
JMv0FGurNznL79MDObehfiq5vdar97G8HxsghvW1QsglZPxzuKw2KWc052UE8oLD
bP4MCXfiGlLjN87lVURXp0cEyB/jE3u5JQih66vuk91EEQ+ilmHxNnKKPH7JNTsM
nOGOTLWJwMD1VAwxnCbv/9x1JUh0eYYxcYituW7UNyP48xsERcIBwhhfv/iWaBSO
pWJDlLJ9skdasgdEXhuSxF9ndW09ywEzCknYYUkTZowsU6yD8FnD39/kl9llZchE
l4C84ebxms+qRo1Im0UISCAYhmByxw1+1ukvEQjQ76XZJdJ4ua7RzdZvf3NE2ccH
swG9mZ2UO3ekEh8E8PTRx1jLEKPTmN70yrNLy66b0eh5x1wcEkufrapGJ43Q94yj
a4Lgqt2+efGmEBpH/45VMp47iWMabmN2P6h4lt6sCddoivRTZseTY6ptX+fMUZIs
+7XC/ApnVL07908cP/L8p+ipstB008xyBXeWz6a1ywIOE8cG2s6Tl9olu/XT0068
7VS6JdveLx+MMEX+Y+P1JxLB79lVX4e/mBhko87k4ZuKyciGZSYQmW/jg/bHx/QG
eLrRGWXKZiHcEGFhWgTiH99X9ScGwNfHDClKFTlMsbEcyi/dujxoa6fF1umY90j3
pMhsmAKo5IC8+IkVNhrc7Epg5pHFcrZDYZcC5dFXeNF3bws4xsRhAD1I4laAjgk1
PQVWpOJ3C+4r7zKdYEBv72LMQSuUoHgHYx0DDcaRJKnxSQKraaLe7I7kz1fNs5YA
ldsDSUTKuAk2i17gq9WfAiXFkyfUhgsw9WztCtNJpMoI4Vx43/WPSjj3kXQV8PhJ
jB7KmVgFe4jNTHYWAUS5fHgsn7dsRLIILdYQMLz6eeQIEJRFMri1oPvbal14zWAo
udzJg+6GA24Yr26dfxCUn3VoF3bPAq5wfDwG0djNwcEqEQ/delqVGmfoQwnY1mGe
caAnt4uyWoq7ZQ8psX0bs4HMfwU7kdo82vzGtLBUXlZeyOJJohBydz4PoG6rGrha
GlymdFIi0incjvz1bUF31zoJC6qSpTuhND42znuW1e4PzYKJPnVNFz5UeaeWDc/m
dTpVs2UL5MvyHFVAPsBmmYl7qzjwNP9D6Rx2X6oxmMA1oKmouvOsyeipBJx11kTI
Arq+dQFgAO5QHjY3dTrUgMwOZj0I2dgCeXciTB3hepLUYN0E5M1EpAxH2u6qO9MS
Rqg1JBoYFn0gS00BcyQSs4fmBCIox4YQ6YMuJXtc8czf9w9AFKvWr7fiMkBiW/wZ
sYpLHLZaTOS4XE0x4ZahRPbzfAZC7ngrSxxAUo3H7FSHrAzkjeAUBGJ2ybwM09dB
XBMvLutrSmc/eG+s5Lzk2hNTuL+7SGamWQzlPDYZLKYj8zFLvlErk+54d4QzNoK9
nXKPdN+ocmLIomwqenrWuEcNSqBDFFaa4aghbTJH66q3Ajcy/XuvqBUf6Blceotn
UaNtPVaNXLu0LgnUx/4NrsaitfArLIUXrrWKyNAWLuqpFzZdcEDDqinBUcCsU9nk
MN4qa3aBNT/9Xmb28IymkTTdG3MDDtCDMKkx5k6TydINpfyyQrXsi1uXO2inxX9j
5Mm2e8sMvff8n5fFcntTzdO7am3eJBxxTdxLyW4FdIITLm9z3PAhT51fY8oHwBqo
I2sdsME1zKAwa9mvn9gTrYlzxgGjszUVu9KjzfxORWUqw/oFsq+pO3+Od5+M2283
KONnTltIzEaL+c9DvkcdZU4PA2IUczb49CR14UwyqINsW72xqJJ2xaJ+JbrDhenw
s6fd+WvrsvFdR6ixdQ3xfWkkmKnc7QFqYVnPAVtcvRplmtsZVlEJEsSXalrQrj9J
hRi/mEhhI+AdGN2asMd6vWsFSLuI49Uez/+Wn/wbFFxh2r4tNNADaHC9ugQwXTvY
BSZCAPQHBkpc3HNZxNJ67uOyCgu0zo9NHXo9To8iRIczTDvYxU+Kv5ccfrGevOvp
2hOKU+1MCU/FLkwETAKib0zz2wQEMMaxJchFg+0t4DvA72a7JnU60G/Ld7rRtNqD
XBeRuq7rcWazB6LWe1Zeg3omZWmbL/hF3SNBurmgPhBQCxi5/4elRqRxNZ2mtGZ4
tVX6336jcv5p+6SdQMXWqTG/ixzOB4xKXa08czp7bRX1/tgGHfH7IPctg61daYhD
yVXa3JIO0bMBx2hb6WW4Ri1ez3bpGx/RO9LN9Q4EXnOFwzVUv8lNiM5Ep1RZTiQN
EIWim0MoN+zikCjj8MYAYosiXP37cZLHVYbSisUEXGGIaL1wJsXXlIWx33i+4iD8
k260HlVHYts6nMrOtdNkZ2Ao7bf362Z9r+1/0uMbYh/1VcFLGfG4NyrMrvwHIGbU
7KE2TQQvJLlCjvbD4sI0qmplmc81exRB4t5JDYPN8wwoY03bjvtY1HTocwID/vPk
JP++qmEAMwYVc9R7HwbtOjEmorR5jt7+AHOZUckiRI0/iFqDztuRQEQF5JoQwuL0
S7Jc1+a7kgjPDCdg4RYnRZ5d2yIRv9k/xsY49/fehTk3SG4lz7XB29j1Sw9iThGJ
x5F8Tt50WZS+OlPQhjLcpbitMkJBsMc0uQa+Az8J3cxhIh1H41yz6WlM0K24GW9p
CzxFL/YVtQYEH0uwCbNZuCHIP8dNEjv57fImk5584HOEhzgDdLegOtHCGG1QGfYp
Dx3qcwHRVU2CGB1P2qcEGu2sxj4U5TNBzkcTL33jhnuk/sYsDaaU6qaVvl+sFtQj
DKH6s915GZOQhEOdsfFm/ROJoAy5kw2IYRpE38MfVq6EFHDYL8wQ+xbWLBVmm2BC
XDRsA3SCzAKcnwCQEEvA7XaYwJX/tztETu+1k9pzkTWXcd1J7Xeo6ONUQwBsxyu4
MkGvBbFwdD7QYJY09UGFoXohTcIWioOkIABxYUeUWRkeYdQiY76ICvTICCxnBzB9
sTaDteLvTiOKLAja/p/Cn2g5Kiqc/w4jcZvZ8oEfc0V9d+wXaU8NFkTJg+rDh3NI
XD4Wo1asmdTXycMiLvk5WCM95ZmKrGlnM8MqEyCtaXzyJXawuxea/2DEUAZB5O8n
aH8IRKjeoQPPVMTz1RF6+sh0nnLOCkUApRSXSLJhvrC+gKDLGkbAvjWwhu7oXAqC
WtNAf6dWZ/TFrrW2s7EkugmKPsFKc5vCGGxTWBrrgqFKk1PelOQfk5rxW/iKUnkQ
iQt6pws+Zd/V43uP5hXBW/zpp6nfhqcfeE7WisY/uVDAcFyCWF6t7OTV1qv+LnEW
mPYA3Zs9/yuKbobkgo3mHy8q83eN+mJu+CTBPHMyiIrWcfLBnAnM86tQmg2WfEDn
gdIzT2ys/K5mnOKNn7p4LlliBWEQa7DD3kB13655PwZhMzmX0rp15CWbE5vg9kuE
snUzR3PKl9SAl2mWomezehgrL23IYdbpPU600DpL0DrOe/DnkKD5a3gNm4hyEbKX
rTX98ZNo/KZGFsjvcNexYrcBCdUg04oLiS1xHdTZzNq1y4hK+6Zpewk2Tp6c4tEQ
IVf0jS19C7FQ2uP9xcOsbYywHhvTue4HLrGg6izbM6MzJcTaJ9IHkeC9nH9agLDb
rHbiGVXHwKMw7cgxSpbBWHmRb4B9Euuu0GXl1w2xqbi1jGu8NBI3LhdJAohvgnLl
e1H6h137IVuwJqTutrmEpyS/SmF+07T8mqapWa0tXVZlBG4/8ClswSOZybV5JHm5
eAuVeWBUO2htDWJRld4A9CDBGnG8s3MfP0BsN/ERTDim0IP2Z/za26s/MoygY0Xz
3cM4pxggbqpE8AOL9GhYg/jWam+Zwsjmv+OmLeSQ3Kov6H377DiXZsMnq4juM/Yz
AYRRHFTdREhQTQwMKEGrhXr4h1rQZJQ1+scWx1RfEzwqrWBNOvuukmXr7bAkr18O
nxZS1OiWSvPSUPwlt4GEeaPpeUd9jiuwcklPVBnKm4ZEYNgD0DkshqI35WLg2WG9
fx2hglDUtTOkq9IBrAmtbtRSOlAtJOeVI4MKMGvKhEejuXXHHu2rb5E/VHocLJGA
CIzzge3HYtyHc3aM+YPj8avz+h1XZgxeeafVFw9aCBayKG24R1UxaQWAS3CamG6L
ZhHhTHeXRiBZmtH23IJB/FGUrIHNPrZGQ0zTbUYMY9SsNFoZUSDY7i1lRy8W93R4
reDHArS66+9vxQUXe3CviW+fITss6MjDmqm7c8bx5OorHG21aS2lZKTzakE0fpVe
xcv6iZ8KGqGOT5naPTaN3UH0VNv+n9fOMQPEOu0shGNgaN6B8Iw2EuB+MrP5FjKc
QSSNjAqRs8QplbFl44t5H92rFoAZIReOqh3iqkL9F0+XFwcIPPnWtbHjl3zeCoXo
pscukGqVxxYzaugHhHubXTsAfCjYdJXxfIbjruByv69zQ6JnGK+tVibyqW7wBz+y
dFcify3btA2w8zLbEIc45wkn3vXy0z7lyoJm6cjXgzLJVDcWPwqSbBHNqJSqWf+l
KbyULPKeT4VUH92YiInYgNhwCeYFBb1GsEHjCB/4DCd199aQKmgg+qcCwLjESRMq
ovs/D165XH5NoxMBTasWLB+Tqy94VCyE3yA4u2D4MS079bqOeQNCdzC6OgDLvJnZ
Emwr8RsHeH0RlKI/CUTicc5XDf7ScxVqCEaaRPr5CBV234XASxm6VHMMxUMLmJJW
vofaV24LrFE+canvhfIdZXk8b5UMk4E09d4d17awvkIY7q1fzZyxYMUmiwqkbUxG
M/D6jzXWdz+fl2ee83KOFBg16eLg0E7/64ypeN5sxiN8eblo9VmWrvq5fRScxbKO
SsWWq2/HtPPf9z9BXSkXcF8BbHvvfvrxbD85jf3K1Kj72vzDh0kVRbvoMaI6s/UH
L99qdD7OBl2MzQRgKR+B3NS3LQc+eJ5VLdIk4bqy2dUDqZp28gc1NkfSlXMPAPoC
R6+cD31EBqf2aEHiGXoWfdzWlNeFLR3iNlMBOWAHhLkw5ZTHwf0C7ZknbLhwoBIX
HZlKJWT2Uh3EwAEEAeEir6LgFhUgwQNv+pDzxssNt/Yb6q4Xg44qeEQRcLZ1Hx0I
n9x744SHNhV+hDsZMTL4FhH9FRs5QW05NdkpBX73fCJwD/nkuo55beSAMC8ILygq
F3pKHHg32DoalCmHCRNFDE4Nefbz7MKWswzg7ExhzMUEkGKUC2bYfC17PQ4LGm5g
2Tq42P7A4fkmwDaUnplWOYNKOf3ho0fEGlDr/ZNAdTeK8FyXgY27Ex+7UpHeG8Mi
vBjrhY7i+Ac5lWLEOOF8ByqrQh/xSwvCPktDwN4Ked2akL32pW/2gINtX0/6dTKU
jfzBGzzdmN23RQXICCOBSCTTReIj1Krq0hUhpWONjb3qLAJZf8EUUV2u76r66cs0
S6rKRn7gkK+4cAMjSnFmqA+LbVZ4SMq1P/9aZFDARv9z4lUuZXCmv1x+hEljHLhk
tC3pjC1OHMct8E5uw1+3gsYUkpuOcfDIr93ET6AWWL06adZrq+U4KnzVaiE14SxT
9p1wHHhMVDLfjWygsIaOptRsjVXw7AisK7fMivU66xxbzVvXzuVVBnXax6e9Lw8l
g0CdpSizPSN6owhgLVVNTgIJisuPRAu577JgKJf4AmS+p0LAh98yJWY8RhHeuRlh
tnZmswMVen4ytwpaRTXL04hpr77YNPIdUlKlPeE3fejWhG0VR0tep8N+wioUnh6n
O2p2pCkvXq0JU6v0uhKqZRwNjvunf8J1IjhgVXfUnFM+1asUvlFxSXx1f4Om7ck7
8pwl+jiY/DoWcbzMVxXeLoLcBbAVHK/MWLHsasuwXQad98Fw1CGvTNkBttCYQBUO
WjOYiXMCR0fguLzp8w1FJuuC+C36/eBLc2S6GBb36A7CAzyVjjLIN5dIimzkG3K1
djES39FHbrLb6U7u/bjG6jxH2f6FF+hM1BNjNxOy7QyxoQ3IszT+ZAeTQBzV1xuh
ZsuEZuAAknbN9zj4gI8DgjfgTwtqTsvuOiCLTVq/6QXICvEVnA8myIw6Ez9t9a+T
TZTZD9RNwo05CFysShWDLdmxwajaoKmO/9I+49/lr7ZQQ3asK6FQ3bb/00TuhTHA
XTXeFij8nCSu4899ssZIZMGATe+qiKyWr80mr9kqu93eWCdjmyLiTdAYb8oBk3wb
v5wDmmRjmFuZWCeEoJ96ooDcioln/nAhfaafA8ykW37hDPhtN0TdT+4Ce7pWa2nM
CdwvixIKx3L6LNWsUuLp6AI0dQT508hQAx81iWqXg/cSWZxzjW6BbHfrTLCitz56
TjU0+hyRJvRaCQx68OUMx4mDPfImeaZpZxLdCpbNhtd1RY4Oe2BsHA31ZDC8Lt1E
NGjDSDklcstvMwcl7TenfLCzYCz49qvvv0p2dhLTs8v8S+rz+V5B+ZoMrcWtyUiq
jeDP9keM8z/f/2H6aeym8/hG5xUc6XoBDqRuqpQqqdW2E6KLg/uZwVzvGKSOzLdT
HpmleHTqOT8X3CtyETKoZJUI4kCajAFQfUPXQB41pkftGaoOgpr6pA5Y2OxCiI03
OQrBPZo/nS184D6uB412BXylpKCNdg9vBOFAhCtlMuse1Ez2pqqYwPDtZUvhKFdW
FbNujCXQPypKWpcm1WJ7tn9uWA+UZLyRUE63YordQqbRBOc1SoNY9sDV4MEyOOQY
8any5X7RFI4ncB0sSGIuqXVtaEJ/Z7Qlmu4lt5NLruGTacu2UuGJZWjVZ5ZhAmuk
QVv624izudTar+IYbangn9Z1y0xz05JsyBiZtK5oBPPssNcRUCDGucykpGV7wg7T
dKAwGK7stsF3+0WWkzGyKiTGiRMvYLaQsqUoorpZEByakCkVBXeSTrdV50iM93vC
5OimASxn/AbamwUZKYMj/7XLHGleJ8xXk58klOiv9Dns+bzJuVCkCtuHwZCGVPha
MbcluohCm/BO67mB5MyOW+HiP/rlC9kMAOQ0/16zof1aj7An2llB7XBDvtdMGlw3
2M/luwNUQT2EvX8kyNxORlYv/fC4FR3QpFumJb3uNqBJWlB7EgK5Qwu5cOJxJmwT
PO0kZcnu7K5GAd+mNe2opFjXzr2OokiNrmowQ9qSZOaNXeMPdzgDyi/ltAEagYHw
xKy8js8FBlttDrMc5/5ieW1elqOGRAapylM9bDUlLxFSlARfV1yhmuQjGN0j0KKr
U/qPJVxMShdSl47ybGipgzQOXtrtfRVW1dtAs4D8GapR8S9gDuUI/cE2ldVERZ7c
geloeU3YHQXaj/Je0IDD5NfmJiDbpAvyKSWeMyipL3+vVBYA7u3zqvDLBzg/DI5c
ztFXG/k2cwzoEeTjTiBgykVlAqlQ8eF0Y36HTP9VoNK17JvGzT0Lf6Xu7OmuUv89
sJjFP2duzbRcE0KLjlLVUL444VYrb4OcJlX4uoHeSZaAkw0WU3vQ17zFW2Z5/dNA
xicYjJ6bZ1AsWpPu3oxZ3HO9ukQPTyxz5OSSdOBNI3TXA/Y7y5F/u8E+EaqFoWvL
JVXLSWxCtb4ubNAFPAwsno1N1KB5rnrcoXTkJwy09KVsv7EvNKNzmQ5+8AErak8m
H6F0GJCpOqoE8Hm3nVcws4d5ZFYHQ/AasVZU2xQyhjwUcks3C+pvinVx4lBM8GMG
UrOC2LBsWBOhvsPTRPmdobiTjcUkcSKG44CRtDjQwbWI++O/5ABG7p4jQJWhEcU6
VWHbPG0/yZTd74xvOjSrZpdyHUXgsy2xb7p87V4Z30sW47MdPeMoQJmbvJbqnROd
kXcHe6bkQ7wXkKa9lfhz6oZADBxc/4qQyyJyu5HgVtdNzBVwaXPdeXr+6++Ad7NY
OjjNs7NeJu9u/JFy4UiV/or4bGLKrSQD+ZK3k6ndkZyDEjPO4SzKIv2ZJB1huX5A
rPpmc7mpqpwjYLzAgS482MYRf+IBbdnb9K3FGO/JVeNiLzWpFWkfW9uI77EdVmJz
iR3KWKTw4O93Zp1ji2pgpVLnhzVdruZFgxHd625xepE5rASrl/HsP41vEZIRY0ZR
uaAfOpFflnSEOCTTSbpPiuKpIa2hgUnEw1UdnXDa2ckqpuSTCb3gM/IXSZbZmLnN
AuaRUKzTyHC+A8YTYcn59onehrA+761U3mXk36hTkN9Q6fXR8XWc/zbtk9+LrWyI
ZUwxQsaxqwVgT+H5X9rXVC5UUItkJlMonRxU1RQ7tGxp4WvzyXeBzhkAlzWX5Wsp
tgTFXciZhalddSpjCnOZAevO35sdZUeBOPa/ualu5bUS41SWnpf3wfKdkH5qsgG1
/XrIjunTc9TneZL7tWe4cb2B9EtwZIXIAlZAMnI1Yr6G5wiQUU+K00sSWJHuGmwa
vT6BzTyEE+nobGMzcgXd1TqCTVqhLh6+VqbB7639Vp/k9C9yG39kw6iw5WGrwo6x
IxC72vHiXo5+bPOEDJ98g109Q1p/61rj2OS+eubEmBHqFzTpA/C9jOSRaK5ujzTC
1RQEhkP4wmYmZqX9qLAk5P2P5vNm1EjX7LWG0ls3CBz2czw2PLyWESBgtj7Q7iYi
+Rr+F52GC8F5OibFvdu4QoPI2WvSGisbDk9uxy/h6BsOjMUBjSv4gUblesjlKC5K
dBjsrXx6DpzX9DN2s2TUySkTxuRVahjYqZzLLvTq9rhQc+3p/x74Fj/tjo1+Zjdj
A1yUTpW4PEFK2/ZjDXvkntL7Dn3hvLIUrAiXdAFyBtWAFt2RvqCG7t6ps/mABUFC
v+c1thKJWKGeEyVc+pzr2GUljT67G1IHEO7e23BBNXVxbBAzsNLE8jHtqbHojSy/
CNXZMzFWs6yVdlacfHQTHUQVCt0Beg6l4HeBuwQXiJWdFzPVIJbsJDdZ60NbaSYS
14B4SYR+0/hyCrIVvJxF4lXb9g5NXutpCP60rgnqjxpyHqNtocR2pbpYIcW0QBxB
6GHcGEXeKPjwFZxNvSh2pJoARBD4R87azKpoc1Ka21V8/OO0HLSThxgSFTFud4WW
vzjb9n6SIAiEKK93k/OWYhvxE8XEUNvXBc7QdsIiUfolsMaU1GQOBYMbPG/JaayT
Fcjub1X1W4yFK5r/UDgFekJ+cBCsau28DZaTMxpkzZFzsxPomH9uHmNezzzI0UE9
XnmKvqwH8m8pB/w2459BeZyJ7U7Z40+7PyWhncvoEwKkewkBd8EEblDh76j/JQ5c
XS0snw7i9iApTE9HN/NW8pA8Eu7rPXfa+UpW8RSehDIKvAFYY1eVFPOobsuBAFUQ
VmS224h+2JMXGGJfvcIsAbq0XWFB5+/wM1Uw87oik3huBmd4J8EUio0sXfBkDZqu
lvBtJEtjExHt7Djds7QqAW+LWj/5muLqpGfH67uEBdQAlDrdmtMv7EnXwE5V9TB9
GqWoqZmSet3U7GN+sHghsfWn8LwAcnxdy7rjaHdzUaK9fsUa4PPqYIGTQxlwkXIf
LqzGewI84KaX8n7lxpTArCxlDgnebw/Ebi1Uwm2ROj0qY8uWKh1CozTBWauRkC/C
HyzW55tg1kDgKiPxEw2T23/ix0auLac/TVN2H5Y2UcLigW6SkpqXrLsxj3PNkng1
+tSok7LQIoLFIGXIOrqG4uYKZW3DHO6MAnPI3Bgvt4JTcG3qsb/P5dYnnqNxxLgc
TZnhcMCk43foQdCmPmPgC96EXwmGTVcA3gvhDbX/ANTCjpFM9+IC9JwYiBNTw+aC
y4LkrqQMowmyHBLW10fIvGZS9VZ5JzgFdm2IcoDofdVqn+zU98rrkcBtr7021Pyp
Zpn3Qp2026zh5Fcqkje02/nTFQXUsXi/gkOWlHSdY7dqzjvJefhIkN/uuGdhK7Pl
NexskWoYW6ERuEv5dD2B2Bi+dhO6bygxXVEt5fQZKNLpFQBqkwMuqXhZaBA99Vqd
VwChJA4KE2m867CG9TkekY6uUcAyiUSFX/qFM4l0jL/vGjdZtm+Abmbmf1JuHKUq
Er1BCXj8SwOcJMg3m2sIC5KyIl5OBc72CJWTjovkBHxlTGQyGohBA0k70bzPwc4O
YQm1VSzmMG0p6XoGQSnzYmAPBsGLmaMw2rwrNii8e+aCjmMCoq/sheSrslbcSLJq
daMboO3aQ08Jd192YdtOJOw78z+lyM5pIF5zhDwqmnBQrvglbxM1ID+E+K7531SC
+J7tzuowNBQu+Bl4Iqh9tV4/42mPNQSPSx1R0NC3Wbf8d8OAdm7rIaKr1+Iv/DQe
y7Tt6SdXk8wn9+O17O5JGs9wRymHybU8O73tcLce2ibhfUiB6zv81ETkwtgyFWCB
OWalMB+R6ZiVgxA2NBkEDQBQA5A34Ries+qiwvXaMaujFjHl9ikr5kpog/ptkV72
/u5e7EijE320/hQ09W/kwL7n8yYqUuEG8VNtZSENd0UyB0nLjQWOgGqdvKwsdQx/
oO0A/N961W4ShgjVKReVQnjSWdFe8oUK9weBvQdrTid+KR+nmJSSozDUCnaoZ0S0
mqb4ildOH77zBRAZfnFyz3948dRH5YwIDMXuEUW/1wS6ZJ5nsquxJiY5raHZBfxk
7uQfmAEjrpVFgxyBvEjML33krJUoGOY0wGp3zZ3163bsfZ/+hPmXYvUBZr7u3VaV
XJgEmOVNB2nfM3gi+Jl9QzFFgY9xNpxGDhE935QRzVyiXUCRDkbMyOYg+QL7ebKz
A8sRanoQvlvS7qdI63ojP5r/hIvd6qsJcsx1y7QmgmhslxojTs6wsbacV3wpkgNT
EOUvFMXqmKkGVE/SWG8MxYbkDMXvOQkgNfGZepmt1jhwi1agpEmhPeo3ltwI6o+h
isHSosaTxTN4OnDXuvgm6fZ8MCSvV6rj+GKRlqzm06xRwDIFgDMNdiV8pO+ehCWP
iky9smD8HpU9JmqR8Sxb/8ZfE51hIGm12XSVBbdJnLGn0/XLxOZtArv+DBXkPAO8
52TbO94ZMni4buz5rW0rEXsriBH7zVwPFRP1q+mpjrh6lrHYFlLdOzSjxHcFngk3
XeokMnGcbQcivbu6aa/gMimU16qinguBsycTCQiPR0HrH/AmGqYhQFkF4x36sda/
+o9qP7nzZlVFecbJ30Se2I2rxPexwnaq3KOLWfDAYNKJkm5LFxC6Z1fr70lTTVWd
qw4fS5L0lEI9N045nUIA9FTXlGUTikfeTdqFWsX3+N4kLL5vPMXiELZeYquMo5xO
7CupRjF4ofBGJwJA47Ujf0xNIcWsIopXT5q6RnBoJcLCiRHsK3M0TlWtXGxY0Gfd
V+wIpzRbkj8DcJy3sZHyYh/uK5dyxSDIPa7ZsMftfuNLB++S+XhTqM8SLBXeXkQw
S8cqNbjrHMPxxe5oOt77LHhKvl7l44ZIJuFMbI8e2qun1bDtkRXGxnoIArY4VHmX
/xn0viFy5Ge1LmhOHnqNVsF62Kh3YSYRqLyWmaKlFZV2m1z7opkmSLHznUhU/iGL
FRkkBjZ3duA6mHIQL1jhEXZTsZflvowAVRFo5DG4mysp8Lx5Ul7/cgmnC4QdbTHZ
xIocYhsQIF4L5iAlJfmFAWQPKO7GDZLVEDm1nrDxnlwDOOKN1OSYJfpTyAVEyd2+
WMzQg16Bt78n5BwBYXDCPczIOjHq/t4n40kDjNbWY3zeKlzj41kh74Gwi+lPwOFV
kvQTziLV+cyltw4CRz6ePv0iMzB3+vfcUrZL5udGINz+BIgxt2bbFJmP9PLx3NwG
mJTeSbA/u9mGqJZm/dSWHULXT5IALvJWWHjArqA96rsRofSp///rmxKlmAXWROzp
ZvEfqORJmpWcTEF0CSvGWyQyt/t93GbSRZCAMREaZGZYEhJYqB80LFwkLEbBrLta
q4h6nWrBZnp2nOIOQstmH0OI44LPPvBPFWa4wQWjKASsHRm07R8mBpcYarbCZVcZ
Fc/W+/WhPq0Uti7SL6+ege8Mbagr5bZeFq4gwx901+RIeYv9RwEITKpm18VqdjBI
yhrEXziReNNboL4cu20TPTOM4AL3NP8sDfydLDUFD9dMlhkl7C5Y9Ng7gXuoz1eR
rhcv2CR1muqX1eq+Bg4iF+Ys10AI0BqXydzO5xyN7HiysxBdOcyavTzfIX5jiWnx
43bVmKDhq/tXmxcCBITcFM/p1QG0TKH1kVRpD4TBA94jPY1ENbOd/Uqwx10D/0na
Xr9g/sEjk2sV7ZCmMQGADMZN/ZL/gDmzsCmDxY61eHAPhNq2Ym8eIbm+AjqCWw0v
b/jUXJnb4MoIy+RlEoY7wal5O1zbnkiHwiWwBlpgC/ODVMVBuMktkn0JivqeHiih
Wl4+puqd8uREoMeBSW1LN1NudK82nDHZBv9Wv50+BWoEcauxcWabDKaL7gPABg+T
i6ftQB0LC/P10OtYLoyj+M00CNJkVbSaRExukQSCMgBpWwaPKFJDZIDNlLIOFcuK
V5yXdhYBps0IYgX+2Wla2duLIVfwtaVNPvUtxUTxbLbBGrJl6muKUkr7aovX3kUU
5XypE+JDKEHw6AZCdtk88em1wskSYeiCra5xsos10efoK+S5HaBZMVPhhNnHZGCx
sv+d3sx8BisfuTjzrcqZXPPm+UMRCzZxB6BW13Zx6seWmurLHzqzF5B9glYevtbX
GPFOxrxmNE3jFk4cidlKSa5jE65oQMtMulFRr79LSr/FTiFCDOpGaaWYGx9x1RVk
jGRXzXusGs3ya5TgfuHtuA0YmoRuayrOig3rKIXk9ZvpPsQ0DClHD47EGhsahnu/
TdzHvkf+41SYltYh2JWuns0S9BezyPss8kX/DXSfNaIcKCAbsevpA+0mggH2OONH
dl35+3lgzgkEOwVIZljFEsgEQw9HO2nrQvIa5UUfu6uRWX5080ARc1cQhG+pHBHm
DPnMTl+TZR4jtZ1p1GB07tvWrsD9O4zzKbuIfWXIz4+Pu2/kjVYjwEsMvipRAKq+
AFP6em0gopHHIp6QI81RkIyuFnaAUgQCAYqkDVqHRJsIaZv6vmIFjzluMRHpwiTR
vpyfXqJbmXxDggmNmsh315n7VriXsGP3UqxKTNqEPQYuFSbc8Ljx+v3PobvJun5A
t7dlSEleplRK1CW0vxay3mJeEfxMFOXbUt/kYoCmg2XBaNpBYsyFOn+H+pBEhAZb
tNWS2GssSmYuTt40dE8YEZOC524x0i4d0bd0RryGX/kbSNmWkGEH8s+OP1j+UDBH
GcbUmFIgq8IIF1MHyvNwuvwHbDe9EFBEes6Nk326IkmCY/ZaqDgnXS/1K/MUloaZ
1wtgpCAk3jF8QfYiKLNZcNi8ka/t17uVZfRvITG65Qej5GPaN39nTU0xjOnFVN5W
DqLq7ATAG7cuVEAmFvEkyC2hN21kwBlyoNkLnjo9VEdGcwb5w76859wPzLDWOA5L
dfdxhPhjNHrPMx9ewDa22XK5cijJEkUlNA9EYgTVw+noGy43rIJZLxsxf71zfc2/
frrX6Ua+H1FUBWi5iIHgy1BlbA29q8Ls5zGo6gzGtTJY4dyYmqB4B5yAeDlj0Eka
K8172OYk7mNinm7paMyvUs8IpG3M5geTRLJhD75lEpLGgaRACJL4rRqbpdRWFXFz
zCTAKh6xQGQh/SGqZnykewSzROAAUHpjQDrnp7YERIHX4Hl/ze9gpLvcGbyC9vSZ
F5IcLFUXCOgivrCzc4cKaNxmOZxL1eEfK7EeNkYTGte3pv0YkHmCVqHK0cAoyvy/
CwKTJaGLksFn0OdYR2LdYg93FMUT3DFuFp45b3MTuB/iGHuZ3qdkedRZftnoJyYV
760FUEnLng/k4vLyJFDwcFgIgxzMTdOp12jbWJ0bbby29esM4ak41OHOAgDUc4b1
xZUeSr9nRy2VQcLks9SYuTkSF5EGyCvvcAdcLeP27CDoVEh8tdGsoznCKUXIMB00
6AG6OuOdsSOzIfpN0AkL8uu0NLn7zz/GpYDykriFdaUIXR/SUcBQdd/fUSV26jtG
dyi2zXx7MXXbGlx1sfXKhJTtW60RivJ9ZIy4x6oCf/C34W/OcngpOOvGIrgY7VYH
OpZkcdqj7kaRhEQIKR2ncwsj4LLwWR23jhFY1ZnOjgR2gW/u8zY4FtYMbCco6f6q
tlhVs+fNNO3LU8xWJsajYIadDDin9ZzaLYxg94Tbj0VkRm2vU01yiNZcgjMfk2XT
HfrWwAgY9LajqzqhwVjc5i2vv1wnSbXW3yUvYebrnx/ubXvZa4wie3fIHzUILBOs
AaWuw2cw9XKvG0STxR9RrINFlMakoiu2C+JKsvOvxn+9YK2xqKohdGxflFiPBzDV
VY11sYqInfUKsVwpc2HSTJL09eXg3d1pfy1XYFxUXkEoet4VjppBHVWN0YmtVqgv
/iQZ3KktLHuM3ZtF9inWxnjLSOsmhmiu9M5tH3eX3Mqx2PQ+QgORyyUAXU9TtG/G
wBj/jW9iVpK1EfJydNZpP6sf211M1BZGS9xfHedkQt6Oln3x/0e8HyExMLRGSIo9
jUlM/XOujlXJHha7sow5eVYGT5IqRmGXZN04eF/QPJ2rQX2fIOw7UGRhv7cUkbRa
MNsJDK7c/9OnpjTjVBCRsJdE4bDAihX5ZcBjGREfw5fQ5+j5GwbB5Jee7xyGL/Qw
COQzulidFUvONyc5G9RpeM/5pkFtJ8fuXwNgHk+LJg+qfMlK9QrxFH+Ze4GPdfKc
GcB5etlkMJwIc/NnPEz/UJVqBypQowFQkgcOu8p759Az0orW7JMUrZCfw/EswdjV
mio4/Tdx1PMIEymCYlrSWxs9fxiSga5vADo7x10yoNrcQgjxfCV3602DTTGh2vz6
up8PCbcVxgXIcNbV4BJ9YwsSzMNSht6gdK6Kcvk03JFEbu/RuGJzwdSs5x4Ne6CP
CmqOmJLXG1A0ivs1cSw4UXJXIFv1dpyVTLQ8KdoUe5na2y/UFlDRCQfnt4ZnDFFk
yjLPxV4EazFHKPwbTLl5QXNKLOHupuO4mKdX7B3xOHqO3rE5fGsr4K+P2cI2sONU
p5EGnavVOMDF3Vk6sZlkf9nAVY0xYXFORPbDLQObVUfgOfZtUfL0R8M/C5aA3FrC
sLwx87edIy3MN+3h7lOPR+inFWDH5Zi0AaEuP0fdnV2Yy6TP9YGpkc0WMjyCxRbk
MK6FvoIIxxM+Gjg2NrSgbMOm5dRbBu+N4d9jLpHfJlBY7IzliKwUpaYTbd6p0Rdo
4/dPFDWx44++gZreza20eMFQX8WKD3tD+kK23kY/fQV0p6lkbl2nrSmsUGP2fHw1
BPCJ92J8DV34fb36oiHz0hAzzOySEjH2WJrWh0pRgt9aaR84WwpuZ1z1RduXVzIk
6JzkEQURr1gxVr5qn5cqMZtq9d/UXVznnZSwZqDFaLWX09XHQExDOaLY42+TltNh
5SbBM4lI5z6T5+Ir02/X1gUxLL94xAHo/7+F4EI4kWGj5FQBuBs8LUHTZpjPhAFS
W/WfoVayFCvLRzhkxhojtABjopbsMda/cAw0Weh1db9l5wm35447QT9nHKVu2B9c
kgfJkiiH2iEJD5CDjKSBKia34qypfElA1ejcJOjdPwu7A27iJTTUWA7pUJUmZyib
cpu5eHwyc3B0SZ7w4hFiRlPSgNI9tHoO5jz+3vcZtlK7HNFHUkv5vmw8HY288RkH
dDevRRkT4qHlrGA2/yutuUMna0l1ULUTsfzKyhZIPu4j+QZkyys738N1W4QRXamD
YANKQZab2vLEwWkAK0qpGN14g91gHDLAvn6SSCtEIYl98yjGmXqEkicdbGB8+aKz
hi7MF7x2y6xpsJ1leADnDbpqCXI9n4//hG34jUqosSpnjIfTpJ5cqxd7fg8lM5Vt
0d1pQ49bT6gmMHExIDqnVquI0J0bZqaILY5ql562hJXXkoQN9Asp7QY2KuU9RIwA
EJ8fSBzAV6tLi8Af2/5GZQjNYW9k25HvTsSs+zEo111x8oF7QcGA0fk3rxLs9sOe
cZPHmJZpANlpv2FC5a0dxVoEHwdcvKzuXwR+hA89mFIXoYgffrtqMXc6nj62uV02
aG1yUPYBz7no3Z/STJ3PV1TFrUHBmdS4WCVCQZqejWqOM5t+hUJCiNq/B7pyoWbs
0g89xDH2vTNxAgzUqY0s/Sgv3PfDpL563nHula59ea6IZMN8g8sEpxX7AUO3BYpA
9p6XsLljuY0FbGPFJ/GZ4o132vzMXFQkoy/FxrUEIwIcO8Zko52EFVEynrthuOX9
w3DtdC5ll+mBy/z/mdTR2cpTAjIcJm5cAQXxzjcVtUYHlv+TWjtD4Vg9APRTHGHB
sFUMps8sMgC5G5lQFnXafKUppY+vol1ZfT4l61cj81/fBORkiZzKsp0uq8aVeRN0
gOZ1lnG7U4OFgvmN3KtbqBgkJqS88dRsoCLMw1xaqTTMu1EwMm0JpW+FldVXLGZB
zdQHLIaEndczhCzC74G50BVS07ndSZ1T9q+LKg4SUDn+Zp2JAwHtUbOJvkSmfSoM
EPReg2hHuJMmP5+4xjLVZoO2wcbPNUOo+Sw5Vmq89q5P0WI8ZFIkFxzHK118UdLH
+D82sB99KFuoqSsOdpyko6nJRhEiOjPc8DNXFjuBh8QYU6eknSRdcVeG6hzfmYaZ
0/5TWqBSSjb1Tat+fQ4Bv/hpS/8CD8vMq14GdxL/IfB3pLVn0Uy2ON+JwO27btil
aAERI+26ySBCHoumGb7X8a5Vcx8KlZx7+LAsUbDWtVc89d7LvBtT0mdnLPLwU2gx
6nCfRcSZi5Xqe6+T8HqCKu0LcgncfLFqZOwJmhyoALlPBelLEsSL6GeMbIWy0+Eo
zwgTo0kGRQCTcinA7+gp+iiJ5ztZA1nnCVhT0jgF2ESypX4HA66jnlouWm5Etz6j
F8CTM6QzRCXDB3BJhRRXzYvOE9GfAJSHAJUEDu2USwsS2hVahyfgfm315ajKDfPV
rQvs8WIA3jMdTdkv05fiWEfls8VJTG1H+xzyZ5DRkRHlc8YmWveb5fYdwa7X4hOy
8RW/rq9Hb7leH+XwLm1vo3czUgCwZwsgU7DPufjovrWtKGENV/Ph6BkFhJ/Y0UOF
IXp+13utatKQTnzZHLnlS+AZXVZVVKGNoz26v+OHFdBKwiF1YoEdDgmvERkgrasK
Uqu4w23oQyph1pQYjAKz6YLKqL2PhZtnG6XNCedFS0QY9A+Vq66fj59RXrE78GkK
VPBj8Qx3P71cV8S7kJbbCDPhOmOySToWlHOZfbmaaV0xjkrQcCK4nLhzz3BK6vqG
3BawdtyKlCQFEh/VlqbFhMmZohx8jMBn/QKB7nFQ8Epq1Xnf7AKErFJ6T3IgFX/c
am5Uxjzak1djyz1TDFdy61Ag2FnrF44dnCBKPdzHSIjjB8WJGvQue3YngTR2gtLW
BFe2EfaCNsencZyx8uoshCyJySOxge93UYFpe5CVccoBChiEvSNKlOyxG23NcN5J
SaMr+jY0mVY9mgLNksdVJCOosDkwhNceWGh6q9NtcS8XAtApRmc6RSbHncbzpJHy
yJi8/v2wfzkQHcgJYR22MQ+dEI/D4Zw7ios0VoPxgHrZPw845L6AAx+egEZWI7cP
eDue/vEtAp+pxZ08jgntZXpfBL1GhVZZeqjbbWXtkCEMdDKGZnsdMYVmH35d3eif
e+e7wY/u6mNg2bc39J84+c7ZhkdiXSVkPKJVL9sbhR8k2jRwx87PTzguPZgJYrKu
vIXhXL+yLR5S41Zz87d/Z6kx3NwZnUkORyWEf/aeVhmpjxMxgKVSJmGf5SnhHOEk
jIug02zIGhmgaLKg3n6dJ/i7yCGH+cpYHGXFY3pSoSh2bJtLqPbFxC/wFqKKJPSu
4vKqXC6R3jYw2IYI59t6gf5S9GQyQjfCJDliih0VU9tZjB5g2y4JSTNNPiqLyCY1
6KcyfHtB2KewqrFHIQ/UThVVnZKXa9PXbCF/jpIlaZhsv4ApYTZ68Z27odOKpVqJ
pb0Kvf4braCL9CuzoWYAM250LWgI7psFg/N64l8nJhj7fLW/BM4/FH52wGwwhznb
udJfXBYks3DhNt3sOWSsRimgwCJXfnmvPgJNhJI4jXiH59pCMj6E+u9YzAt7xcsN
Od7GUuc2dhUrNnPmksKUrlz+0YmvYjXvoc+HDyi7SjYd8PV08TzRyxNZkEj7ZNzp
6tjE3YcaspS2liGOLJli8ZuoKj/j5M9hbCiFx1HHzB9wtpMTZSij2lqofNJOMSLW
6XrK5sN+J/0SMn9iZSG8qkycux9mp0Glfmh63UUy9VaL0e3oWI4xoWGrN1hbufDh
wzEl0ac9Jf3xqQH0P22s4Pgv7vnkepOFHx/N0qFPOO2rI5vLBzHHMNjX64Fw95vV
9hLo60/hXM9z56bOK3nHSSfsx+KlxTq+HHALIhFB8oXUrydEycNQkNZuwmqpNwxX
b6L5xhmI6owz5kVZt/aI42cxU8PK/EHnsIgdaE2tQS6PVmjS2zME0Pamjorxfryb
7gv/0TvfQTOciH5HW+7/KQiHw8NMJcjeGMFPOOYdc5Pwn3ptHusmiXMlBlKOgEea
TV0mC40eh031alfPgj4qc5zSYx0wiSkMoP6EEVsWDtESwoM9r/ktZM36ABaad+QC
nj5czSJPI2ryo2SRzHMZv9FACEh6aGxo5CKhWFceFQYz+hYOiUSBJBvTl3S2Ju6Z
lRqowW5Y+DNG0SSd+7D60fbwC7WcG15379DAVJPRfbi/1osMBv4043W6qz+hgaZj
su8QonLJKtZojRVGbtiU2VeSwzmTH7qDCrOOhwn41ey/3ilGVaDBKlCClvjWQv7P
0/n9kIxC+YWOXVzkSSYJ9P/dQhw0shPgpDaySjHNQsoKSt+zsFYwWo9GthyCfieI
CsNszcwQDdzpTTYglSu9orSHxGmGxQwfpw/+HW48mzadkW/SF+efxvIFNUrtpdWl
76j6x9Bx8vcnrf9/nrDvQ42saz0D3Tf2jN6D+HDdhxbpHmrHhcXgcDcX0V3FlrAU
mh9V3woj1Md3yLkSNnPRm+MuWFiiHMeKQZnxX/njR35vlpqIVtix8aNzkhsovgkq
jnsZFpXhfGHZTZTKbfvcuixX5iZSKdZiluW1ODU1SqwEneUsN7bNvJhbQJo6KNUC
4aWC8/cb/yq4s+rDN1zPZwUuJRxk64B6U69FjA8W2otA5M2qRqFZ73GFCM4CK+NN
5+JGkw1lWwIVZygtjI0nk+tyoJlWKvAQ2suPBcujdMin/7obrNb6pza24BkFE5LY
IFKqBYXqywT9k+6BL2Xkwtq7f8F2iAy+vBMYjC5eD/PhSrYCei8/8vBk+XI+DXUI
haboWYb2HjH2fkjUe/GkwwFtimi6AHjU96XJ6qD05+GXb0YBHkvd3/vd13CavCo9
fSzBFFZtRP4RCAnIl0do8ZCc6JXOWwbGg7OYXdtajEYx7biUOK85qSo9THk170VX
7i+S4W/EFqBWB9VGcmjQO0uCdzH9/OnaKAq2SLEp8actbK7TNCKhI+Ii34J/WK2G
WOe43L7xFAH7Hr4cHd4kjjjMR9JxUfDJblhY1+bge2mAy8K1xiRVENjjfLSxV3VQ
8y8065BgfS1Lj7dFAIhvwyo6ZS71keWX6DbwSxyR8WDNThKJeFonZohJEJmaFNMy
u675xHwmoS7jrVH2RIN581zFlxiRBNDnphTaw2JvpINYgTHl5gA7BaxmtncOCoGE
x1g1jA0c6u+OrsuMttM2EN1DRAXjWHbfTNEiiIeozBw8lcWJEotyCr5hRdn4iMf1
faVjctve2ztxAwNqs8GQVPVZqhxRZDq4r3l0myKVmb9/LpDHCbn/OItA9g8M2KLX
ybivRWRGV7H6ppjpQDJVBioWtTSTJrr314PgdZYmTvZARKjlUrN7tJESbnUgDdm+
1UC4l5hNrx0Ci7UNr+K73Y5ZVPVzI6BEe8RH3OtFDu9UoyRrxit8XiGN0UG/AwWD
7NgDa55/Ay6DfOPR3WN0S4iNDh5nQI49KB9Rui+QuXDgve+kqj1N0IdwgWDHBMhL
e9jTJYXFHDfSe95Sfa2hPmVAE/OkDxYnn57Isu/m6IhaF8MLmcu8/YwrLFE/jahc
jyZrb5fQeDc0P8LhRQSoeNlpSB51X2t1y1mBfiYSZCIJ0eUY/V214eMq/nOQZUgD
ahCG7IqUJBAoqeGY+Y+cl/onlWoAiBCQXzyac3Pyy0lLTLpJ5gW4h7GlKthRCvhS
e5bPD4C3POn2CbctRDfLpThFdl5n9B+wZ+R2A1HC7Hqu1WkNekucvkF9X3fq+Qxe
OyckwBTl/n3XDTHBsIRJgUAeUf2FFw4hyBQ22nIkaiB3/8EgU/vsWbw1sqsflZWt
lw06NAlqYGKiRQTIq2xj+LhwbIuOqUdIe3jWl/9sxLS3xo9wd1KzPTqWzIMsuYny
YepFFyR0w7PbcAEzmHbgHBSYUZYiMfN4emN8GTY9eE5UyOztPhjpdu2PuU9eURdw
oOt5GdyaOWrNNeaTAG4TLxHn+isWv7BAVmAlumGn8ZUhzUvCgSDYP038epxc7nnP
ZJ3jb1ztR1HwkK3T3zvi9FhhsgpWXrGtX+6XEWLwnvAqqF2TleL+VsFb1i5y+kxk
CRt0XX1J5I41jV7AvC1PMJHu351Ur9Bu4x99i+f37ufzoLxpMC0pUpT46uCkJgFO
NK3Yzp4a8OlByQdhrUgr38tE4rqYZBt2mhyN6wigqMCqijBoU1tQ2oifXswDbHLw
j/CsvedAKpHH1wP4CopTJViIpf1IrRR95hzIb3GaNlv6+ydjDnFeSuQWSHfbzyKN
WYfdrJroZ6wKAs/9zOeLU49NTtt3bYYCMRF14sUmF/zFd81tawfUi3HKBq+R+TX0
wZXt0TdsPp3EvmTMDQkyUQwoEegkspMTlZDbPscbRckNGjnyU80upZ2qtPTgrzGu
5twxVUytFQ7kUW95zG4K59DhhK+8ECe6JiYDfip3CcrXZ/l3tLWebpV3xN56rMPW
kiLNVxSkTgmCxlQX4JNbc3on9SGQdcLISSGUy29K8r1rWKmC5YTPAey3l4fzgr0V
oytMubOpd7FWrqcRa2NAUy1dwQEOGUIdWFzAHxm2KFQ6ESBa+5aj1khYqS/VfrSD
r7Fe3FOXHIPzFcHMPM7KK1Hku53zY3hR5tWE3iHu/cee8yY+4SqmpD8KVtsWti0z
fUtZhMGHBiPQtIz+J2+tgH1tiBG/xiwWGrXkstGgqK7Ik+dHKaIGXomxB60x1/Ck
WqpSfwbCOdYEs4vDSrR/9ZIC/E+gxE2A5+BYQTio5bdrLWKxmSJs+NPNDlBdQ3zK
zkLzgctI/LHllxB5J66zh06H1g/SwBN1KVGHvLtsuBuFpYzD6h3wk31l8xAjS1zU
vDnAWsfqbTTlEt8fIbzyQuaAnVxcIX/36tX/i1etNZzDessr07g7n/JAaqomNkE3
mKS9uEUBEZSxLlxsKItUTe6SzWAtcd+AJ4EE6x5OsKJj+mfum3heiH4/AwZ8UnGS
5YNeZHjVaZfQf8giOX2jLh9OP+7YX7LLYYDqf4c3zAOmmw/CH0BCsHLJsJY1qI4x
nqRYo8ZisVpGaPgb8SQT4OBA1I5uP529vvTcp94GnTRMP0qzdZOfNyg9PhESwf7R
9QGDjJGZGZBkupAX7PnuEAWJxt97TRB+0zw+G1/LNtjZov3FKslTD7/LA3br4XNt
wIxr9V1X4fMUtjwmGVDwwH4eUvz8O3VL41eK0PoLVmY2hldcAICHLM8xBx4Jtqqc
KsTBY5khucdlivt3ANh3fml9eJ0mYHbVG6r1KDyQm7u4l/U2bH6kw4tn75xa77UJ
wGb2zm8DLRE+yH04L8qWbYi7tnZw9xWeJYg84ryFDk5IGx7kEkCXGRhpxXltieKk
2i+aa6vGiY18UtTSgYfeJK5rakjvd5UfOfvCjolMT6ApU+w4KewMFDf+yU2UB5rm
qR7QWevQe6A5HykItyNiEu/WykrdmnaVqBftWY/Zk8PoMYFuIO1iQ8o5J6/aUgB1
+7Dr65j9JqiS741VbSQmbCNeqMyhSj3Oo0uJVATjRbpjYPS4niD5V+jHXVqqN27T
XZbgZomIm7WLfxGEnI+tUzIGd4D5eJkQFLayMz4Qu2DUK+uVH3hxquw5kT5o6nBr
VahR1Adf9Expx5SmeLPJkFYgqUl5qUw3m+SBnOGL1D8DezLWzPsTQuEhmzkmqeFk
mJnsXeumPeqqy65OiW/8OqyoygHFUyhQQ6s/kRcyYgDrkavJeUvp1JsarmVZ+qaO
TRSLoZdPghuTkRaQ/f+baOAx8Y70gON+e0Yjx6Pz9f9UaMSBK5gj0JciPSXwBXly
kCKNUCUyewKlQxcXqmTnklzHOcOj7LAe/sFKxsyBcVwWAECKFvjaR3sSTHHXe8e4
EwkOlwYQB0M6NYnOv1Brwg1AFh/PKB1h4QNzpSjsRMOXwX27Ge3ydJB0CXztSZeg
LxnRubJFX18bQ3OQWMKdeZLKEFBauysxULLv2fqzIV1h9ZTgFTS72XHl8LEU8a7C
HOLNoBz2cvRFdmKjkXWLjcFW7u82Tv/bomZZZjeyUiwqJtxTasJc+mg71BNZe+3c
ylhFXOvgOVyy+aruDOQMKcxLQ/1pi7oWsbnxvNv4Q7X2hBfj/3e1kSF9x7F11Bq/
HljcsnCV4B9TV/jo+GUo/pb7ojHz1nLxBuGBfiq2GWMOqQHFxNY6NFfV/A5QSLYi
P62yjrmmlVXNqMQ+vKqqvFO3QEDFdbQg3lIc6zngdpW+BuTSi9tQkF+e5bQGTqD3
po4vyb7WPeA6acs7U8fAdfm8CwvSDLiPpKpeSLiQR6UJMt5IKOZLQGm6sev96Xhb
QidWvXwnM5qCHIO4rCE35UhR4i1kgs9BTd4opoF1XKvPtjYhrLEU52pqHY5RfyZ2
wKwmNd6uk02ZyVVH+WSG5ibkczHR002MLT+fXwdfR9R/6zI3j7PvYiqYfh4eIq6/
Y62LV86DTwK69vsdfNwvhw1HKEgmBrPtoY7senxHM6Z90QM8Y+D011D0W6RIy972
hnGr/Wnh//RxxBwChFOVhCVA+cVnSfT/KFFQVLjkFycKzFv3TGtkBZSsxpSwxcL3
rQZ3ntcE5IErzQDuEPOzw0QWNJqAz44eQG1p49s8/F0+VqYuhf9dUwhxhpFQYD4l
odZQraV1RzAH8r9WXZT26SEPL4KjSo2nUC+jwmhDMpKrILWTiuUtlpxeA7tmFMVu
Te29tBWzWN2omgwW8oQzC6l1BYtb1ELtDAF04yTaKu8i9hmCuSB3bVyqnMZZisKU
b8IapaKCV2p39h6T+hkHbUnhyOJNdaimG/lLeyEYxYhVkNB5ONe6aKeTBK8fhfdy
3L/HkY+eHxavNmoLdgV2arK9cY9ouqfYup2K7kz5lzS77qtdzVDQHrb0aowwOdk5
mVv7KYwFS3tlRVMuZlREIrKtpsqA0MDnprIKxlQz09RiZcadsBzwM9gfYFU0LSwj
H+5fENzek6WqrsSzwPg0qADSBozw4tDLOYFMPcnYsolskHZlq4cEq+SBihQwWqFu
Od/PE+s1b2MLoWEv+SAO1JOwFSN9RNhY7nCojWoO/nH8az9vVA/r3mJpBMbxQ5Zh
aFH00q28jHU7UJ7FvjfNJLXnNPWyAPtfUTBpeHmsbtVlFhkPFdLx2IgAVSwhvQCF
hbEhcmBs1BKG9VKE+a7yA8cKCDU7pBUprVNdd6lb3hPYPxlhs481//XbNUdbDo/1
n9Iog0wstb1FFbQEbMKo90bIXmb6izjFWqeUIUTNkdAnFeZX8SvlEAa/UxW9z1NN
PUEE5tIBWtQ+Zn+L7F+nM8FlLby9hzoonDuGju+zYFhoW664t7+iQOe+gCvw/gvG
k6pQUv+qC67YondWRXWAgMx5BxRszZt0TbKm5QUti/VEwcfZzDa+rygJzmLQDb2x
h18QrQRiUBG6pVj8dYVpd8RN0eJX7EDeh7OOZXaQ98q0CJENIef+Pj3QpxEJjTrT
kfdWvVV4lSQGoxZHiGNbJ45qfMneYdGhOrELf7fPOntDpDi1QDRZmKo/W9eiPzm3
DSvTA0zpvvkE9mm+CldlYhESSf+IHtr+F8kPs4oYhNrhNkdH+HyGx4ff2YWVBb+9
2zImv4OeFDALp5p2MXJXfaUm6IX6L2Ov7I9edNf/n+wbkhR+LHXAJGhHkJ2uWMvl
ldzza8e2TD3yhNu85FKQbI4KhmxBh4zGwOCgAPymWbdrO+0ISrfMBD2lklUbmd9d
ee4x98Ojp488hBgLjySrfu/UOyusRTkghIfw7hG6kcyP9sguL36rhMiIVU2WgQ6a
6dVOIxVaMal5HExMoFzy/onkomFCX5LWlki26nQQFhL8pK/eWmqLfgt8LYUc6PJP
o7IFKjzGERpCXw8xKjU7mm33/KEFqsZY20SZATSwdMXmDYw0N3oSFQNJ5EAckli4
M0EVm+5jMA4XEV1V4xdC2zLa5JHeIk2g5Y46ewuLy+bw8VNjb2IhKIdYjca0wjiO
6cErL5U3KqNuG1NBaOzk22m6UNyiyEYKZudkOTbz506v0ylvVb96Pk3s2/+ODUZ3

--pragma protect end_data_block
--pragma protect digest_block
s5ucqUS9BO8kuZ1ugAJdeRv0PkI=
--pragma protect end_digest_block
--pragma protect end_protected
