-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gmK0If1+Ew1yFg91B0UkBWMTGsYwbI0wDIjBh1Xi60AaaI9IwCaSSpKQPi0HwzhL
lK/V4CpyNvDczVpuaLfJTxLQ0jt+rskDODv9NgADrhpEMQlw2bmOWthcLsloHspD
GcSWw3JtuJi1zVZkOSXI+ZFHX/Ng4S4xv1lL4IFTnW0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 116307)

`protect DATA_BLOCK
NQq+MH+sibpASXD7jxV84FqL4qJ1+SmELAfDQIN/cp0Ke2ivdi4uU8RFbgDTOa4I
nIaSHaqiLxV4UN2x9qDnZoaVJDMGeq9fQlLWmJHMt+ZY3D75AEdkm/eJgV9GCSFT
MOiQ29IBeavufAXCmWtWiGO1hzfTF48DXiaNfG+vRzuATI+F7cxOYpd9ES4/JXvI
Dslg0w2e65qZLX+HPkwpurqFuUU9N97n4ifHuZH0VrYndtKHMesdMahASys7zd9g
BdRzIO6lsfnpQEU+FDMM4LK1pt7emWjVLBSFATHGXvFd9v5uPYW5jzZ7rIgeopEX
scYT3pOPIcCgo22bmooFGTTZMa9VlZc3DA86TRY8KwdXhZHYLGS/QKA1Ju4+jxrG
LJwIRCdtKhnzozTQUDWuwt9XcospZFWgS/iQRkJMRt/YYioSc3qFay3CX9/2Gp5s
XBOrfXr63ByNl9fRK3P9prnZsfct+wwyWh1nYow1sR2RkzHlZ5ePPb//Qw0XYrC0
lyYQBdbprpSxFPEr4YymnsuwajdtqkGyXjCuyC/iMYM7ZxpJf8Hqjp5Oj4F62Tzd
xTzmJ2QV8Enmc8+wTtFXOGt1J0OnG3xDw2zCB98TiWn1Qv1J/XmoW4RbNgf9uL/q
GkbBgtdgt5cdk2pnbTfld9uZTdGWDM/RQFJ9OVEn+dip6mBvu2e4r89Ng95p7DNX
57AQdeGwnnJR5i1EZbKEsnIPxB3p+QOpO4piXyLQZ1HHred9+dOSVAwimB5MWnmO
I2HAmlssZmNlHyzL3lsz3OmVzWEaVEVSQV9PiBHwPQDuPCwBukQfACnCVxNq/UQh
RTAdpuLcRgyVJ9tpEyq4awdwWw5NpfkfEpw2DL2Nyg+XvO2iQZlYRqZ53SwChR7S
VYEw13I6Tg5HQCy4hCqIIbuTTXTpPkLByBZTcBQAyV2Da6B7vpjmgngYeHLxzEot
1FcfFb5RF87xNTEm6+NzzhFQPRG7d20iPeN2DWWMCWkc2l4oiYpjCoC+f4ynd7Oa
p+TjQQdQ3UJMqsUyRUAGUXuJyALBKLnmKwyzbA9JblT/mI2zsY9rn4pzXO2uvsVt
wlm39qrDomRve6374sncdUAwcgn0NIoOzA2WWT9Uk3EhQZJ/86Jg9moeLDmoF2JM
bbs5/wvLsRm1HU/uh6lrMRfhHZGX+7Ew+3puKxKc7AH60VPiRgP0wI+9giduxgQC
iw45MB+s21tR60w6Ri7DTZBmFBi0B/jkBfv5sS874l6IffoK0k7Sm1JZYSy8RURl
owTpsYy3UYeMenkenE5hltpVKzJkQ7za8gz2tEqoirOzJrO8zI3PYHcMx4FBee0y
cY6LlNvNjPTdjmVX4whsIlcWM5saBlBdY6XmtrMQIP/QS7GLXuBR243u9hgLGKfn
7XprSPu8s0JLn89PLmx+Hn74mLTkLf2XfFskxWaKfCuZpXqPfmGoxyUVFjxkhDCg
9I8Ty9rsZprhooVb8yn1tWgUl8ny/w/VInNE37U1uWf3soxLP1/vfEWgJ3kjPVrb
SXXyGA8s6vbp5/V7vfgdgp8YWI/wF8OFnWz/fMXYGn4ULaK8hh/TkBBfHtDrlnqa
8JZJwAkhg70CH9FGO7jtqJSovWEhY6riGAb+iJ7XlthdrP+Oo/hSYfkWqFUGRzFA
AQJu7RL1aIDDOS2hAowpWgN6q3KFCjXcABEj5cUNK6pjG6dIcETaPYsVcHTZybau
xBlwjbzpuo8w9vnacKBQvxZwyi1xnPPkIlDnXQOXiTp/XCkEGZsveky3wsdZaj0g
/95Fk4WqSrqm5Bwy0NVbLA/KOQwEcUiI25SuXm2QffAhdbuabQXTZJizqzoQIIv0
ZwM0uEFqVUobK2E3741pFrZjnWhTEHCBedZCCq4J/b8LozvvKniOlu57sGLEfh9k
gj8fLvaUCQe1w0knbEVh0HYWsXizNyq6eurFQIDdySK/al4LajlrOEDS0Zkpj+jc
v2nXsjNPxPZjKj6wLDMXUpdNobgXSN+k347v30A0kKSlGx3nQZ4OCCPNJtYRYKrN
+Vl2Ct7EOJXgOOSBZxUo5yJzPjyvuEyvE93x8oAUvOdNRMw3tIAL1H0pOjoNNQyW
7/1vfgMFV4yRDlzxa74GSkckBxGHwgNclpplkWScToTKQIxDhCrZ9kAxYGg3S4x2
by06OaoVbpd4W1dypW7GF971Mob1cnnZGwj1524joeA0Zvsfc84kS3CpMEv/xCCP
3en8zhl8cjLJdUs7H3N9eCzVE8Dqg57G778WTHAVW1kdCD4kc3qweEajxLq9RI6T
hwpMleZjYFR283fH8iM+iBDzT/7rAfHk1Es0sPJqmJCGms/KJesfS/xHpkZH55RA
IP0TgEco5YdQ1vAB2BIvhwvlB1L7ecLwDoRWuh5fbCf5gTpJEKqvOK/tRtYXYqCg
KLWVJvaVIfvP5Rs9ObRvQfRyODNEVSOsv2DJfcSoeS0cxP6rUNhp8lU2iTuOx0AZ
G+3qoWRyNhmCEJ8qf7ndzLwlo49QbN++jj/FyHT+qr6CJIP809GNPA+H8ga5naXm
3ArKuzRV0ciGzEsxZG6ZIYSeLl+kF3ma9TnQ7hDI9xZDFDHIt7APtJWCi+tECnnF
N8XUPOmKj6wqiPdjlQhekrwakvYJygzCAudVkN7MLOhQYWI1s/xqQVr72Tg7EpaT
i3H3ZwVG7TaedUnOoJroqBTwQLVsNaYfJE8FbQ/PsjWd6Fh5hoxm5y/UP73bbK8L
5lldAJHvW7G62k6Kinc6K+6e7/NiIg/f9cgy6q/hrIAxz+u2NPtj7sFInuBbXQva
RwhW2PMWiSrormJPXW5J0gTReso6zRPydVEDUn5mROHR0QAhmEflsAc3z/q6iEkH
XAG7XuxnxWWmySW3Df3LnMGoaNEzBdYlpnVjpD3WiJ2vIetovsg2WM6X7NmT/0T1
ZF4HwNmgDToGiEC2RiS7sW5/s6wxnk6Arf8G4vmigJlaCOyzOngY+9zSTWwYqdye
nqVQXk9j7XtL5rz2fb5/a83SP9gi09SKZfQVXdQezomNUJrlO/s8aihen6fuKWmz
12RvAnVJsb6rfds+gCkpNDwncAHnqn44hPrGmsnksI5fxHavLSibNmCYNtardBos
AKW65t/Lxf8db34Ekoe59GZwWcc/B1CB1vO/LdO1kvzrlnyeNae5ffXRgjldzzTc
bU6o+NnPGdkP0WLRzgqG0XCOcbN42cwl2Za3LGb+jXwRR6hbDWGCj+Li462wVEAj
rINsi8sl2lPt/7M9Z/Ia7jrZzOxp2BoH/pFElTFve24lMb9XMlZyqP5iC2feAtYN
2v/vyJm/lJajd/6xQQMBn0Hgjvufas1j9B9bu0UmhVuiKIktAoGUjIrO+UdoyAqL
IAydfhTmfSGGTft8wSKy1gmigarBcojwz8qFcwiW5Ksc8jeBxXVAFfhKTj9gLxNS
YVirrfe07D5WWLgMq4+7i8IRG4jY2DuefuJGz19iMjg/T1JCGqi56n7FuBzvQjmb
uIx64K0/8nPvMvEHVd92WYmcPTQeItghagysuBq/c51Mi/xDmQuQzTeOzN2xK1NI
ZJXfg9uMmw9MX2+qrcaQdXrSXfCpOlXPfQ696HQI6JgtLNxeSYYlaSb5No2BNT5d
+BCCmYZk+03svoeWWhWOletgjFBtPuWj5xCMrrD1u4zVzqIbUaGNjcJY+bOZMI2y
uxskPVGtC+nU8z0AddQdYwlk32Fhab6/9H4Gove54NjGVQlUMRzIIlyfF5YcB+ET
LfZQ03j+ITeOa8uoNXSj7aY0d3YsOPvBt1LqyXvxq+1ImjTCIpG/LhrFAYH2pO1v
wHwcOIWQ03g65qmZNXfYju9WVpjudkZVz3/pn4VNu9U/ZlP1AxzEQeGqxxBO6nEo
j9SBKuzsaEl9/EV6viH583QmpFGYGjn7r9FLDvrm9pwxUbJUch8HM3feAZLwg5N4
XZD9qNDWxYmVehhsn4xzt2scu7on04iEU535VkwTo9NupgZ/2XzNRQ2CphKWQpOz
prIJbMlxkIbHrHtonT4/9BNPuxASGc5UMRqEiky5oLUeAKhFXOo9Pv1LsXwpzYgt
265Yh/YNdZ64u/zGTb4Vr5lRDldaFcc9ydjnJrM7EoaiM+IekwxvuO0Ru84+k3BM
qls8gmL/sOvt/AOiXBAXUfgqUhw3Bn3BvvkCiXEqVn6t01U38GTAwqCquLT6H4ES
jlUxo1XrtSIHsv/EIlCSZNndcGXz3GuuzcvHL5sJAybM2BTYR2nqfiUZORDhoayu
t7MKU+4LoFD68K8ddZJrbxneODrDdev7EyAghjKPwa1u1ba5Nu70VaUuBqVcvNoz
UXVe9QCKtga8UZGwqiw1gDmijyplKR04kE0QF0JvzaO81MChuuBO3XmwxLPtFPqk
HFjMWTQw4iBwbZ3OVzVyzR59uV1+X6vcwZFv4JgEx0rSZK//qNZKF7hJMGGersaZ
Lvh1BxNzlmUPxrvEftaoz6zgZgjHaqNMjTz97msfnP76bLP2S0/QP+zXYp+Skn4o
LBXCmORvdv/i5MNqQkycqfFDZwZDJRvrLSR/JyiutsPyygpQoI8pkGnuG+eNDA/u
hQ3kQeur7ab5Icuw9gGUnsdsg0kVUusHK7X4wjrJM2hi/HwwarToH37u6g8WoVBT
94Lixd5M9vP2dNNM7SEjHnsinrRznP2TPtdNCqnwR6cVOsNxPv1iaZ4Iiv9JBJJQ
HZ7wbNvvGOTO+51YwtHST3m0znPt81Ox3RSN9e9D91O3os+4OplA/6rk9gJVYuv+
YYJapgZlrx6v/x/oJspbK63n9drcHSpNgKr+uQtqbg5xxgKU6Y32MaWkdmzQ6KB3
XDhpYyebZ2xgOYM6P7LKu1h96V1yWhP94the+SzBipVxjdBaZbK7PK/bfR8JxOfw
7WW3jDMlAk6F4lbogeDcN65qMXnAPI/GXqBjmVWVBmnD1h9J+KtdEn91Eda/HLyv
OREozrAphPSyNL+4ed+B2NweFBBFSFjDo6+QWCkFiC47e//+RN6t+Pdi2L4GcWJI
LnjWqrZBeii3CQG/hy/38jQl6Lb2ksoWzKzuVUnQhWEf6hMf8ep8JAbwkaCYDlHL
IijF00H3+eXJXRwLCWg/NptloUeR+nQoxjAWcVPwsQ+wKQWUOnrry1UiHiq3MkDr
rg1CqOPuX04qAjXv/s1HMyDxq5Oi1dy23HMZlSYB31pSZf/88jmJKrAuEVKkeL38
ZjFgUoRcLsoLg5JcO60K96AOkAA8oAufHsdb0tOe4ap/GF5ApWFt0noOet55Kr4Q
fs7VYCRFtfgT9cwWVXatL4l4fUk0SayAY+f8+WtH+M844m4o2mLpM2dDNfyL0BNX
IY3KVjTIxjOgaK9TqP88KKlMbJ88DAW2Pm/W6zGxl4APZf8HKHlQwoVfKwolBkLH
6zexP6vgrRCivK6rtQrlf64nHGUVpx+ERY4qN+ZgfSzUpQcyvnU2MU4e/fUpTZA2
/Hta2frodDLY6O+GtxyF6XHEJrqTNcg9iajwQ+0I+yhRbhHrttf4CAPB7d36yugL
epeydkh6I+MSziSTtEqrlwY2sUclyGZiXGg2IP+cAssEnxwEegTdGv6CGix4R961
iIKzAQPI0rkE5F0Fw+5/JX51QfRPHO/H9IzhaB88R2f5IF5E5XtmfVCxRdwjtArP
kp/bRxp6kThLOH4fOnhjZFVcRt4L/rch6muRDTs8wbXhFywZH745nPveqRoP/LwB
mkcLGmWGdldK/NozzjCcRnUgcUrk21q5baenILXXCEC84QNwM+gkNbKiikg2HNV1
4KXyVM/qJ0B9OrSbNTWYw0n2Gn3InLxmede2DORspgReglLwliGqgKCkaGsIM0Xz
iYvLzVfbvDLY/I+tHJQufcd2RH+/SNZ6J24FXcip966LKg4oyYEofwKhg5/e6y7z
9dP0Mrrh8D9zQ++S/f4fbnDxr1h0q2i4BEzboSyT5XlXZ3+tBb+UgsI+7ahgYZ74
Uty9fPtBoeKEkEnnes1Vuvn11NJON+/4RgVUH3y4yaXYsQtjPaac9pw2kYbqwxxm
mjX3Q+wmPZQnRJzHHygCfdC2i0bIoWpb7Jcm1Ubp2vU1V3Y0a1xPRQlU02CBu42V
okZPcpAVuUQyv9wD/ihevzySJwseTnht4UPDmjS09vPmNvUUQ4lKuWFLZmr7IKMh
lZlS9gtoAILYS3DqmHG+ef5dpvVaH2TqxKna+tG+UIjnJbKrUa/GRttPe+QvuXtC
2I88Sb4GYyGlJDj7L9kADdcDwdZsxnoEhEp2CkTGtoz73bboU/91mNknBiE8Vx1s
NzC1I813vhrkTU/tvVxmWx14YKRokk7X590zwevK5GdQyFaQdSdliXyR0U1umBU4
vsixqg98WCU2MkiKmgVxPD2S0AvC7mRXTMnPBwbj52rCJjGr6slwAm+YKcWQhs6M
pUyvJIoJjB0e2pDtaBNmPyiJDK7BKCDjS+Fy+PMR3jjKGaA2HLFIt6vjAv+Mt+gY
6u8olTzplhDMjYpPApg+wpo3ITdNasMYktPWPUymyfNt/p99pdidRWU5cpwMGReq
+iziWAYgWEC/c689IX+YhS4IjzGAfwjFasxStzIp/INhG30ejKNg8CQmBwGScg7x
VKyQAev1M4OVql1yN2l6cyxhz2QLTASJvPQRGRZTqBr3h6d0QAHyI3csomyG/bcy
8TPaBjfvsDmJHduPY4cISNjoTwaq336H3Y+T6zE1vFaDHgVl5YyU+YWKs91FR7a+
+pq6CI8TWXXjTxxgBjJdRRTbdFNotGoqyTqHMZk6xVcBrovp46GP7VlKhC2lXezS
LpDWHgThI0QUAgwRqQBbxeMH9Mf+H5mhZF77/ugn502L8nfyicmq3+0ebsHaJGQ7
Q1zhIfMDkMZpMy3iUId7yWmPXrkxGKH3I0Y6TajJ+pAcD7T7Mm5OTkVa+tFaa7OB
ThIZzKqiylXptkDGGwoR5Cou2f65ll2KI+FA3aEWQx294VY7r8sWQx4FxrfmIEJt
jfajP/e6rYqlczAR2jlkpb1IhSTjbeWbeBBzNbXHuBvFEZDIWFkh4gZGLhGCc3IP
oDJF2Fo6YE6ZpcIcirSM1YSAGQrkVV00JyFIbBeH0xno0MpQSVhIT3joSNjcbPT9
6x/dH4/mkpl/52azMVBDxaNnhpbw4jgFZ8tlOXdlmeORqCO7Ca3k6hVkjWJnG9QC
1dpwQuTYiNefHXL12SnimH6d1umAAUxZj8UHjqPjR+/Dl4ZpKDapZJdZYZsVHdkQ
+HgBHLNT2kPtK4E4ZlGQSiEp3jjb2eS+z/dBLuXx/m56k6WyN+26KKBxIqDF7b/H
gEgrP1KAbwa4ohj9IsZjVu76e4i+zNKUWshQg10ki2Fd/KmIZOxrTG1gnf7Ul3R2
SRKcND6y3+rZ32HwzZe4lM/Qrn/DvdKhhAA0q2O4RvG/QnikptwfIH36Ig9Z4OTw
vSLqFprNa7qAkUBy0gJ1v74PS98+QNoTHCVayDKy46njt5XuPAa4xFW06QJT66bu
dkAOz75UIOCMMxvjCVtLXtuHnpop7t19Y6oucvvcMncJnYDH1F49999N6Z1TQHIq
ruSky6H42cUrbwiZliWnfDrNtmkBscmhzUNrG/WrmXez0OiwrZA9RYqcuIUCJX3Z
F68/kD0bf1WGlU1M2IgHtd1hFY821+GV2u57Ap4HqJcxwKtOh+3ogy6ZFbBDNuX+
JSEzJREN2wuNvX/ZQ2wuGGZRRQH5reuhxjt/X67JAGs9KBeHp+96HUDW2MnWapST
ZB7fctk+v2Kkf+dX5sbYfGsNZA0+k/8jrBtO5N1vXn9UDVsv8dSN+OYG+t4/6sln
9+2bjkhtAnnxCVZ871TAIl52cmEbECnVbkc3cdYp3G4hbsiT8e3EeXiWv5ZTEg7T
XmdVq+PP9Or2735K/B3z2ZPt2oHAKoEquCmSvmg2Zc9KqhzEHxnLjAe9oCLvhnwJ
Fz8Mww6CGCjRbsEOFVKt601AnKpzHLWi3K/hIDCC6PuxtrOsFdHFU8oL26rytCMi
cDHk/ZOfM2sV0Q5WMz3cpvPeeIEzsF/DtqK/NEejNF4BeetWZxOYKCy+2zTq1YZQ
lYwOD2tL4XOezOdgiphbBTv7BDATBkEShMdkkHS36j9n44zgFl95Ra2eTDQq4+uB
ZTYmuIsKX5SLYxDczlG+jH6TNHS17ODpUTEZI6PVfF6vDd4Qq76/e+Mfw6pYFCO2
VBMYs9MAv4Cl8gpvj8DixE0OdTbhfuBPPrieJwOcCmTu2IwKm+DuTOQLN2xqso8g
is6n2cEYPWzqSVRI//JISncmCdZqfoQwbX0NwVuXiaDbdtk4jUFFuFM/N+sxzYwy
pxOBVhCgHPD2ta5JCzoN87c1GHtzPyfeCt86BG9A9jZRNZkcyJOAEythxo12gWBD
CJvCCuHS7Oub+Q/s7/BJ47gzWzoMrPfEnfAbGW9iNkcL0idiSTW93aXbWsbNtp/9
cTF5z3J2zgwnJIMmCktwU4sSoJWQ0k6Yd61D1o9cT9SNMNb2DDviBHksBmgzdfzy
4mMOYa4Aux1UxDR1O9PU3b+Ll0EbPaKTFHLxN0MlvF12ZatOQkjfLtU0jkH4GArz
ADQ6vhaBbaAABuOO8fKfHKemXIeSPRF2qtuNRVCe+vDmZZQqrFCOjos6knOqAt7g
EWbRq882Jt++1Ma4p3SOFhGgTJHEvlUcr2Dwxa5MV9LWmG3386M7OY5ie7b4rFnf
yRmDHHJYveFXdffCllQsdGciNBPQVFU/JwdW/aIFv1mXBxH7PyqyfNhFv1Z+G9Bx
HINrzAIyTCAwLJ3oSNqTmsoJx5KGtkJHVX6Byw64re5M4c1xM1j5k3IqOkeiMB6p
mG9M03U5Soq6mmJq5jrWhyzFmqJLEV+ix5ZdIzSR5D9VFXWJlYhyUM/FK6VP7PbR
cDXJYBVTU17tUg1CSj5pos3imczVhpEEGudCIrctYg31ik7Zqfv5IUZliDzyBXzm
joUSFosnVXbm/1jeR6FdFyXREVCr4jxwpbB7++IA0CM1GShhW2fu6kUugrMYGqOu
RwX33d+ZIGYDfmv9pUC0RCrpqCk6Fu7ZuUo8CwsKmMlYxByg48WiI+cqO5WWcaNy
Zr3f2bZ6aRsIJQlTlPCyGPselU04Hx4qmTznMHCizCWsBdlpi6hfWFOKEjE2xgGs
9+DW2XBNAamDUC4fMFkMsi7ISgwQ2ML5XFowRfoUsC11/iSjPLQIqVWONkpDfnXg
bbJYCK/EdIqDPgVgcBRwVH+yDGO+2qWZsLoKdvvuvEwRpj3TYPljtrcQFGfk3GpE
kKbsLCmfDJXGkPL6FU1ctxL9XTFdZXiGD6JaHWHMBHk+JHxIa8RyU3yffATQ+iCG
B7C0O+M9dzG+rN6c35EABN1/9Q4dmEcxrVN3WybTke9LRbjZUe6QwMXXHOlVgtGH
fgXxwaOUQ5aUgX5CL2WYvRZsh9ut1VOIpbO5Eqf1RryTNJsXztQvBOrhAuz9aah8
y1C9BT8pzuV0tZW+Lri/we3Il7p/fk4HW8FL0SjhHB+BzGkK+ARE4YQMIdAosxsz
Vh6f/09y0TvXi/anu75m0Yid1l94Axe2aP7B1jhCBttFmJW/6A1XniGol2G3hgEi
toN/XYBuToAWv2Kv14lHd1LQgxnQkxWBKJoDa45dfAWeHRtufWT0Ob+mpDz1RjQm
InY7OGjK0qIPZ4Z/zTRmZv+dI8xH40iIRw1ox/z/waHrKsz8UZI4fhpTDRpn54QN
0R/Xm2ie5zyi2+tHD8LC8jTYoMhDiFZ0WNThQYHCgMQnUEALpmfi9hRiSEzDrtrA
HJgsgBNslMH/57G10PLS4BhcDtv34rG601NfBQZdfZlNFzmY6At3WN9BHPzxzaSB
8eedmHrZYYNzYilJvv0RYRJNiR3u3rUPTX0Y2MWxAnVDCaG9x4+RnazJW1czN/g/
2EyjDu0Kq4akYRhCpo34sPMe3JYi8kDzlDqbDVwt9J021NfgU0lrujmZRRJiXy0V
HClKEFJNlhR7pg0TqYTgpc4OHz08TWUcJhjusaxUK9hSVWCpvU9GtnqDgb6UWeF2
S0H3TTcY0CidbNrQJw5Z7aI5gkZw7/bToq487MqUi5i6JGEoOvCeUkD8fpZcvJJN
4TvK2u1ktqe3eAue9AkKVuzXrifzaD/uOhwoRMv0G8eEEC0gyirpcZZ30/l6QuuZ
bSv5Ww+019okFasaz6sNg8253w6M+GGLNh/PYojfPbQJdaEzAU4FnJ+/rai7vywi
9od+X0EtWhgELzcrrCMlkee/00g4L0N70J1gT2L1QbFs7W7XZC0XC/GTer2Q6IUJ
hUBDCOqowVr+p9MSBKueuJOlFJ1pvkZwa6n14PicMDcsW9RI1AJQOLMis4ohyNJd
jNPK9qgZNsSHyqIPVC//qVAHKxDb+na1wnJgaHteP5nXQVUxzQA6iJptrRtd2tGP
Ee3xKNHC1SMoo2mrbhJzDwfMtmPJWKWtI5vL8Ekg23P/cLefPvBkmIb6sPtu2qus
5vyI8455KcLd6rJsnV7kwuhy62ZkAtWiCnLou2OpM9JSFQ586yjsJG7ersvt2bVL
BUp3DjJO1UugCnrm88WhI2btCJb+DQe5QfPjhBGuyxxQqcYJjz1uv1TtFOuhlpaZ
eRGZoMQ2/UirxWBHvL/0DQOUHrvGJOdU0FPF8TGAoT9OBezBfkGQUVMXYqEmPXKw
s4O4PFjeBLie1hYLAgzubSzY/j/rPg7VcfS2CHvk8zCAmIArdOCMSlVVUFConaxF
3yUqKRzdMEBVBzIlvuE6Bs/FC7ph9XlFBIKuuEfGAk31j2Gd9lgYe5ujq8Ses9D3
f8VcbCqdykZzSJSMwIKhO2uqLcN7nrM/VH0TPi9715r6TmzJgUAyuRH56J7y1X6E
qrIC2R3YH6U5SUFr8zBfBQJ0xZqs82t+DCq7rsMyu+B/orPXGpmS1IVuiNTp/hjx
OL8w9DjLOM0wirdY+VcqvwR4jj9nAVSe1T3zpcnkrBRzEiEGTDY+U6ctghCEQkL9
Z1qwGrrp0VGzL4drbvu6Nqs7mXjdKxJVbsA2hD6glw6ASy1kM4YUje3NjSjCriB+
zJvBy9hPSCMuKHTpmAgNW5dpublgUtew5Q/H6vL+ARmKgY7sYLoXB/glz4Umve5x
+Tgz/eCb6mZcMdeCPlVgZEvXM5hGLuzf52Z+Wa9Q+SvOYnm4VugV5eTZgmsWj52g
/Gn2Od4u51WcYTMwMPghVU6Q4mvsDDu51SDHNn7rc9VnulX9Cv/jGdF01XjqmJXe
2isF6QK90s4cpVnYoEl9XNk5MRpSmIEx3J1zC5ObC9phaC3brsAQvxY3MIN+kPi+
cZLmWGv2aNWRlxDJ1zQEnOQeAokMle3Arn7PhzNUPwJ/YV9TPsK921ui0inhMqCG
XKrhpSLLs7DliLudDYYduzotSRBMjswFqOu+s05L0x6ZMRHok1O9KBSKOngClvGv
7C/R0Q1aiJpzez5cGw0V+9pjWD6dvzAQQZwRlLq3kyuRc4YMBon6nr13CxSStf5c
760hXi+tpRqNZ7pZRUurSxR5kc9GqCtZsDXOKRQ7B3CbfZ7wcNDAkzB8y1Zotny7
WkDxac1hDd0C9SABYBbMgwyjwI6mEtbBXxZwMrdKb+wvKfuVPzpxE/lkuPYWKA5Z
2osS+MfIn5YQ7LE2ChO+yI2V3Twj+GhW74faBy1qVST9syf58tx3UpOo+lwulaqC
H6q5Jn/bd1HfapQ77DFouGdHSS3oG9edeaU9G+UX325KtldjX3Yu9rD3Q8A8Tx5M
VJ697iz2zI3f0jDCD0bX+iG6PyAgzrNXqdIJQR2UjnZ+mVSl0WgZbFpT3f6SlTm4
itJnEAFSpG3NhcuNCH+FaPrK8xpricQSV57RgXcJa3j2veWlVvMB78uDptTNZx9G
Fg7HxRkyZnybuK38wBdhUvBYfbaq98OT7ALlG5WuqZd1r0+WHiIeCjN6FOj9z+fA
wmCcrHIfRjan5SlMYMYwmT3CbLKBhsu7eK10gRNBdFdumwUvv7utt8dv8J7kgz5E
2z+p9Lsr18z9QtiX9feYpJRe4astsze8mfOA3I85MBjO3QDnPUayXEkZTOCC3fnI
W25nI7igdQK2d+j1OKeVGBlNHsfXER8JyHWht2jsARrAhDv+HxV+v9clclsAjMq5
poUXHh0OMj4V6paeIgQqJKIFAoEK5PaIB+YkJtAyJ/G3RxbCIMcO0FSm+hvvCuV+
eE5MjRNPekFyxe6CJiPBX7OpA/ORaeLkQtYCnyBMiepSpquUOHmdEX98c7yQSP17
29CgIDJWfrjVHiCS9IWfyKeew+yylxpqKjGq8IVH/xgEDIYPRoQTnlxvgZapfZKm
z+VCmrHhygniloBaI7hhtFyAaqsBeHYBBLhzzpxL9YWmHtq6PXN77otdUDn67lKM
Ftv/fg9VO+o7U4NYz3xB76lYNQf/b1FsvpsJi1Qak7q5lm1FT8qWD7+GrmGWPeer
K8AkUXaIKKNDB7BrfAOnew3ifkR5HrFxL5qRPaWkbX/SE+XnXRF3iyYMn4Tl3pjd
iW8b04sKzcSa/SfCk4fqE4i/IlI63/xt/v0vPm1yoMNfGdSBFXC+OiLHnXpLlOGf
PO++BQs9JEWRvbJxfWxQJKx09ZcyAYUWboQI7KiMc7KuJKDGyFTFxDdI5xxsiM9n
g8oH1qmyt+uIeg8yaykQ5GQrz41hVOg6gFKD8f8BEj2cCCQm0x39N16xNaCNiDV1
cjYjg7AT4QXmDpaHqpeqgHGDzE5NsN7R2SjnaU59Kgogf4qMDwesVpEWmg74saVV
qk0MXGsQf5pCPV2MtP3e8Ex4noqevnUfkzcGpDnbxEgJmUXc49qdJryx8DBB0RD4
0lPCI3yt/hmh8lsvpN93j7zOeps5OWinIaRmPBeO4P8Hu/9EG1kr0p3IwHq9OEoM
K1Ubng0PkJsltRaIcCUrnEaHpRGbam1mUpbgjyFuXbIV3Ieskj6/LxuSmF5AHh0J
fRhu7zn3Q8zueQEqCww2UuHzzFm3E46KD34X/Z5xkmFTFa6C5KGlHi/c+GraUgd0
m8miW2RqpbIFrxcKRQMSyp3jE5pyROTmytd1ikKbNxnzZFBGS830HR0PeOEIaiqw
8emjruWrit6UmulC+M8fLES490ygFd+YVCD+SN9kyO8TkYu58W+vvxa6Q8R2S+ts
ufnkHL2A/RzTLmI9f3JwNlwpTmEpgfoAAVC3JvFYPCgmIbP+22+KGPMgUNvQ5isP
A0bpOsx5gdPuuv2MtUTBKXVi2+9wpWI2467BMaDRa0jQ06sEiTZBtGEWbBgT9rf7
cr9ICvEyszDgN7XhJNZLvqUbPQ/15Oqpw7eVwVBO+NutSOE/bP0+zRX3aF/pKe1w
CU+VyNG5Ori9FlpCh3rtVcXEQCChkkLZFQrwChAhXGMOkVcB1c3RTS+X/rBOvY2I
QnX2JczU53rdzvd0hwdZ2lqW+L15is1EbDVczel3ob0wItrCzgFgxfDndNR9WACS
Jqajyc5GMkqBzKqtNAyBYKY9bXySjo8eo7P000/2gIpLbuWJNNQkmuSg5EbqDeuV
OdDvhme4lYZJakXpGzbXo5uxBtLHVZnKy/t0s8+DxUu014P8Xqs8BTcjQeRWv6Hx
FN9BBmvs98BYmc3YSBaImByqKW645NaJ0rFW8z3VTuDI/zglXp6hu+oaA46QtNTW
/c9THb78PYwdPRlsvJ95uo2ErMFLaAEmXg6qTqU+1+T4Yv2++pno9Gmee4cv68Ip
1ORODKghQyMd8ngQci06nUtd2b4l0/1FZ3KxaWzGC7G7kpyD3Z7jFhxA33H53GT3
nIz78rrdXfa/pGwxmTRZUbVFCVgsPHtGgMWjTXmUHhuWjzIeNFQ7IV2fGiF8nPpT
aSh11qYUTDclsyj/dOhIoSucv6nb7gE5iBIvezdYKb7qqAs7CwE6FeMZtiHRMRiY
PORiZinffXDkQ2z41H1wYRl1cayNtYvywgEt+SGfVi8eHaY90Xnk1OO7/9c6ZU9K
gBnCewNZGftCr02wg5I8aKNCfE+WtNdkIAEJ9wDNOFKid+Vnh7op5Lz1HwPYnzQ2
kRQWr5GU7KnhNPawlxQmCdBXIKO4o6DZkafNZpbmyOWn5dGL3bQG7fZgyxwRLXdl
nF4ufxZEpWcSDShjd65jCPttxpzktgFlOjwimhNUqFrEQz53qGcV2GoTnpqbmWqR
PvLChPNmINhZpbKS7c699bCfGUOwdZqIHxdw8llPgZyKc10HZhI4H7B8gFa3XH0X
CAUbO2KHd90G1oZbg3NwSrQwI6p9XscDQW8Gzbj8Dc5v9q0x0nse4T1HP0ar+kDd
QIeNTfcPanjmT8Ipuade47S7Jhq6iQmB9Ra4U0Jka5V8uFCRPB1zb/ZmkoASsWB6
q9/gcCiIrxIYaxKJE6CZG/9Fro6EOLkEReA6uUMFjErU7phNNijRG2UMYAsitwIE
hw5KlzDsVdEy77CD4F4anmMojxU9m1V4mBZrPv7CQhb/zEFFkXY+lFSbxk+fpinH
SpTHROyrOhWTx+fd+WRNk9z+BmpYztSDH60W6Ghghr9+pcF94BLrJHho8ECYkB2e
qmJAUvvxFiCxAdjcDJCQGptBm8zvInzAAVexca5lsJOkRvjpmkQ9asknTh+C07T9
Su056TgPTgyBxXtEqI1yXc7tAIblzYX5oeMvaWZ4UF/16vGXgSiyx/4PJIRDD2XJ
491fwZ8zImcsKsKzOcr3Hlz3lSdDojk+Zgvd1wbhVwmSCsZZIDVd3NlhLUa8XECB
fKsVkOnQ6e2op1nLsiUmfw0CCoG47BsT6fUJxuG0BovC0OjOMZaBTwHAddBZO9Z1
UtG2YG2/q7ujJ8ysNxK5gThFY967tWqVeKcjIPzwuSSr4STsYCF4eYa+lvBICFnU
RKDVjkyRO8O+KCgUaIRTydQcFIJTSGkGxW51HO93rjhBMWKt24YlaEkk2J02Oewm
AreJeKYJc69TqXQa3DCoUynlB1URQRdjpdaJ+bGmapd/YZjFYD9Ea8PHoETeGvus
J0PxgJUOFGEr9R7pUaU0wgf3mj4dCV1OH9JNj98Tfj+cg01Tkh4fDh96FZcEIyP7
dgxNHRgAgTi3s8NZqjdS3r1EFZXwycDfMxRN0qdGETjpX6Boqg+OitxHXsf/nCLD
cDLOHDUWirrPg1iYWNzGaxiGs2dkjzPSGNrm8XpjPVZ/h4M0829nIO4/0gD+RXHn
qUdHSPz4tGFkfLcn35s11m3yk4tWKLN4GquuL2l24G4KWWk3l1RBgsR6oB9K3+5h
cWdP3gRiYOlK+my3JsYXlMJbDsvT/tIp+HoXSp/0HUMqELAWoqQl3ZWHN4QH9V+4
g+Vuq1ArYr6Mr7mIWxTy05DfQJbCp801nLt/AHQHX+sfsZYIUSyZt/0KGgB4B0Lt
uVLH9nk50YHnQgmywmaz4GDLLVrECFTTwWcM8gmAC6UF4pk9W3Ia4lb71naOz25T
zgmLSvobQEOHVgVDV+nhXpaRJFkM6J2oO/hwYy0ZZ2WJgt7rWpE6pfqwvXNwUj1M
GXrKL+C0mGAgwyDPwNOlJ+99NLjn3TTTA7sb0unkus1H+W10x1k4XKOG1O/zGegL
8mIXq+7na1d18mkGrak9HpmuJXFeSLozUpBUIhZNQCds1mLKNELDtop48Ljp6YWZ
ey7Q1Uhkxs5Vm/OJuylNZ/P3dkFYKlS0aDGspFdoEfeCLBwjJFSqBWZaqRlfFgdu
VaAzdZA4GaavQsdCNUADfI1X5pS4mCJH9qwXe9NohpmuaTz6EQSr+IjuGLuqM6Qz
j5TwLjiBcPM2m7+KGdochiNZca+sH97aDGKK9SJuiskcmk4hJfL4rz7gd1Rred1k
MwtrSpFo64aoo9omBD/igTDrHJiDik5iUzWE219NMQgNeVsHhS7pzgHnInfw7auI
TjR2o2v8f1eOY8kGqrUEMlyh7ZcIVT1SsNo46jAMXzoq7Mf43bTNPUenw4Iq5yxT
fYDt/+SJpO+XT0dw/4NjkrwD9OeIYJnwDfdA899ZBZFQECuGr8u2WxfYgMM8Yva7
wXAXPvS7++o6Iud/R6nn5LxqW2LQrQF8jq3JDqWhNR//Cfy059O9TzLlC+cKjaQf
1N+2PW9DN/mrwbCmYu9YQWaezO0Daw+RJu00b02Hj+IS0FDwnuWZ/MSldM4BTDGf
MjRfoiMjcakoTtwjK8i0TK+hWxGoB8ot1iLFa2cpkiCRbgMsRFpzZmB2sFaOmiQa
2R9om3KrByp3xLXVUJsRFXBEBGprRSPT3rK2E6IakPcbdlbHIW0ro1A3/0IFTvfo
Ub4SRz1HLhiXZCBrP5c81JKPDeNzPUnENFX2o3t9Vf8Q8kXBIRClOjyzMibW0E+5
j7Fb0vPjTGn/CME8JyARXcd3e0flRKOsEaoBLZOQIw9nAaorzNzdA+ZB0+e2U1kj
qN4mxAYgSjPUH6GmIv3vETVgBJWAIPR54RCI87OVZyfduYZSNDX+mB1L2+pTlDsd
1Ludz1YNuegUzwS2QWD9vpCJWMRJTvyrkVnUVEiw4df9+p53Fm0EVBXetntlPewf
PM9YRFfBsMW6zQY2OqXDDGGIpWm9rRXw1IAWjuRQF0An5QvOEM2pQleWA9mBjYGb
WUGPTo5Plg+sW20dpIiYsbUYr7sUioU57cWOz7NwcXJlPcbIf3GURiAaz4vrWWL6
p+S6c0SuO7HZWwaXtUr4oK63DlKoIBRg7V06gKsjckjjzoHBwJ+USSkfGndcdNxX
qzMQw1Py++jtvLHH+m9RclqJCw1+U2x48yb7bFV+EP+QL5IHL7fMpecE7swMt+6u
Cc/ktUbFjbZSvGyIJxVvinc8hJWZw9D0rJoRLmMBkmTg1eHuuUhcTrh1EmSjD4xd
oV7TOMsfI1MjulwXUpUy+vgfuDanKPKq1uOjgUsP53XWrYEFSyhqFq4WDleLriVh
AFxJIgmf9JYZ4cka62epEXN6TfqYMv7k+62WvPrtzBAMUuCbAnWIlAAWqvOnBwhi
fPWebWL88jcj+/vOmLOPDW+/NblgzVMUe/GFkgwcIYKi30iLNBqfeWLlZ7Fo10ni
MjXf2oOZj0ocEXJUF0LsGSFOgnukY3BQgNKhRAik6XsOY1Q4Jt0yE+UBch29OVyY
eie07b1qUvLg0GyD3SyKWpwnLwOY6tsu3yvJZkO8VNuIR+Lf3Zh8l54p7IiKoeMg
fjdH6P1EWSyePVFbwWj0jfaw6eM6SE2R2MzSNJmY2ogWi+lH1cBxJ5mKcPqVLwWV
6So8REQVIy7u0ypg3Efelo0HxJjSBmGiPUDyHPk9Kt9yfWJM2d9h1t0wqOQuxM+u
2ZHFGIeF7u0V6UiqQqFeDr1WzMCHHewQl2Y2XmNRqOXigE/4+p1FKLKOcqC7fxVK
3EdRFnHPlow4+6DSMGxdBluWEAp4aX69lAYQKCLrlJJ1fjfZZhlkSSzjnnZ40HEb
LX82bILg4FixzRnvYqxu78nhP1RhYDHQnvcRa+leZjvW0Ncix1G2lsorQ6t21s2o
FRuNxeYeg//4ew76RFMdjD5g4a3bjvUbgvLWCiYS+Fnl5l/ayhBy7bDzyjp78Jdh
cjXwctC5RsQii5ASLqPkLU55jkw+sBTyZnZhTIkS59tVwIx33iHWORsOts0J17g1
jaXrebGs28NbPtjJf/lDzVkNsHfIaxcfx240H+YQ80i0xSxk6hsWkZMoR9nKKhyL
lBkz8CaH/nDqyiHVkaOnXlfAnjIwCe0ah6ts12qpFmSRZaQ4oAIPmdVpyhaZMvKG
7VFoCVthfQ53DRWux702dl+gtUjzvj4enzhrUz0RZR8ETmTYWEB+BLXat+OnnoN3
r1CYkRQHSU0OKmB53VIDsNoHvu096O3hzLlK/wPnfWk08KQM/HeIg7fYu6KDiWtj
uBIIQk0WcQk1yGy22yd1PW9IjV/g5a1I+QmyyFZYGw74uVCGu5XryfKo1U5e7ClQ
Iw2L4IrPPd5rnKhvpvO9vdBfCduYDuiY1JyN9IiwzfY4L6vMhMM9LKLMxN1jGMNo
BN5v6FDHmp5aA+RUUjjxoX35nY+tb8CZ/mUbhBfv5CbA44nRr8z6dvvuicXYtPf5
VaoBy5P/V935RjMJg87gjHotBrK8vKFfS0QTDFW1J0Ysi+3xYkATuhWRu6HHNqVH
P34s4tL3t86/c9MNVylNH6x7DoXy462PlODhtIoJACT8XEM4qbPK71FIza093Wnz
P3h6r0296nfy/2cLPg5Et5QUk2vNzaBe+zgSRN2H9yz8cCpQmI4xCvSHhGvRxiVU
LoxpIzOLuQWtTRh+4sApDTP2UWlDKSxVMC+UtUrGhi+SZGojpSgeewFVg704hsMz
VWK7dB+oVSvFaaCoreILqpyrhRRQrHwOW571Wea+r0EDbsAobg4XZ1Z5RLTonsAR
ILo0sZp3n+oJSaGQKPryL8RNd85NExIDObxJyNzJFRUsYJSMma+x/angXYfLaU8L
SIkzu0OytE9VCdS0yolW127pv3H1KSnfTPcJqYTmiS3kJ6QT+s2N0MmXSsNkMSnR
1WZqRGat4MWq4V1/pNqnoeVzgb+sDeiL7gGiRspmK/dUNQK3MYOtWieqAF1TmLN+
mYcNypLpBCt+8VZr76/FMiRb5RQkIL9VH43u+J3kB1e5uowBAvO7JUbObfThRzcX
K6RSYEjP0cJpW/ocB4e0fG09+j4qkYz5jPyhDb684Ou+x1IUw34tdUW2x42d+x6X
Tna8eNmV36ouUTpKlnuH46OdDvhXUB4iA11KoLvdOOAJwsX+waFV3U8drZ1ru5lo
MDqgAiwBdFmwz513CI4O/8V+8vqfJr1/3wbl1aP2uDBuGS2T/ljjJusPnxwOMKFf
oputKBuCgPBQZs7sBoghojJzhO2l5gj9HOsFHS9edQ+PRVgf3GyEQ/5QQ8v5QEkN
022kpHOVZ556dqub8q57TMt/w5tVZS1Xaw8cchjh4jlegTbFrLFHFFdrPHC3yM6J
7kNt28en8r3LVDSQ0oKiScsdjZKpOkT4ELcrLGAVeaStC/Zs/6hMIJx6p8WjNH45
/52XN+woQNnMs2MugmQW2kNk/KlWD1pjEKQBTgWRcwgUFMrqGIpwImSYWkvxfed5
9ngQUHOLFvGf71w7fh8JaL3IBUtR4aIC3kF7JbtdI2XDHWy5O/78xiDtPTVsgbmv
inrR1rZuFXCCFkG20/IfH+SA6jnt/dI9jpmctBEOyj3hpYX2AWk6EJrW2xDxDJ0f
Yl1zHAlRaQZOIbh7RuxoPSZ2Tn+x3NzA9My4eGQKcrZv9b8fzxQBe83g4V15n5KV
/lH5k8AngFAz29KNPEVVlO0LtIr4KiGz7vAyTyc4uFNVTdxfuUQ6eArHsvmbD4zd
1G5uhKp/Ubv8SFqP7/JlSjqWUNU0n2ficNROo9lLCuEhiK4RS9WBgehIKjaYY/Qh
4zGjGdHUIfjaIdw+l+TtMZAY/QLC8w/w/UlcKgfDClGBKin8TAOyIbhXou58hhPQ
VdYw69KKWLIQFfPtS0qCXZRlcmV3cRMFYF8h1xJQJS0vaip9e5RfCLOmRgXBuOmk
vwq4Q0Q86uaHIpiSay6vqKsPn1m9xBpY3yQOocMYPnz4S7FIDCJHl8H5dyPIBmB7
j4sxhcF8N07OlFn6x7CdPhMVF1Crj0ZlKz1LtGQjRcAjRjx+HU59b1z9dRGoyjYi
FDYIJVdycQuWKac6UztSN4JC4kex/nDuY8WVaF11tfCIWBnYeHESEx8ZpEw6ZXoG
Q0cqOHfJ0FmVkBaSf0Hpjol670+d/Y8SAJuRmJQzOwVuOhoG9B2tt/mhXQ9yqJni
E+ZYLTmLYgPhSJtxk3uYXyZsULWiKYvH8MhhSoLHzPHI3lq2kEfbI3p7NXbtm2Y7
Rd7NO6MC+bt4Pi8b8NQrMqdq7hwNUtaJqpdvVA90lB/Byi65duvY4ORK2IzwqOhK
w69rB8kCvac3iCceXxL1wTeCn2AkoNsKEKA3hOFL4RBnFXUK3894GDKjCSd3/2+C
/meKURGljtEQKIns5pOJRO3Q+vqAxomujgwjzfRp+zOJWTycawJzy+ZSKmyKnNcz
LRCowqkNojWbvbm7g3uKdeaooD3+TZBU5S9KDi6Tr8579TOPfxv24JR6iqeG9omg
OpFftxU4wE4pkHAr8V6XpLiB+ef66rbW8hzejbZ+xYmI0pa/E0j6MxTI1a4rSPa3
ZL1COZDtn6zXZbT9SOPW8Zad7TfPZ4TRFxER4BOXikpOszp7AYbXW/r7sobqHVIi
Vs8q2n44XLikAZYYZ/VkgmVFRmv//FYq9/4P1G35pYznGycrACcYtG7zf9wczf7Z
P4h6OXEko7ae+YGz1NUo2J4wwTxNYoo+XHFcs2BDug89YbFURTYNMMzyVs30nyz3
A/2HqAtWi4TBR1Uh7IsuQsViCg7/Qn1DQcKRC3r5Y8XQYP7EVCLL0pChl4O9s77m
SizGyXfgzmB2khapUgWsRczh7vwlruTUEE4EtiIpQzdpKtsoEWi9IDAWxMAA7p8N
OW7KBn4iVlPn5v2f1aGp2m/PiYQWu3Q4PApS5Gu+TjSJo9qSaXfEzXUKyyOUxJQf
RX2yoX+PF8EZdXI0Sfpr0rMpwgzBDNDYxKgtxVUCjrMjFJAhcvPPD6qFDZTrFwxJ
S1qWLKDENlEUd8JPsXNpi+fqwF4cZRB2KVTHz5jXcaODMfNaiyh37y2u4C1VO0bN
vPSfAEmRNdlPeIf0BHJjiaTcb7p+zp0V5BTd1UIqvU5dVOtANZ3gNBHgeX94FgIs
WplCx6iUfTaPqxTRJyR43aEHuoa7C9upElpdSF7C5Y9BkqkXSTaN2NRREoumOApj
PT7NmhHw9mBaVLsAFgYFCUaiDDADC/3KtBkQVnhD9FEbTBoOJB0T9jir4sN8j5jH
q8qunskro/f8S4sPkzAkTVstpjHUIwslzQiSPxdCrKQAJZgon4mHc/OkO5wb6lFT
PgUNSihcD4aAk9E+r1kuIQN/tBBGfi4GzsHtic4+QmuMAcXmo4GsNef8mCVb6ExR
zZYB4IXNZx8aB0wjRlkOifV053ytdZ/umUESCE7mJDWrgXu6+YuwFvzd3jBGWIqX
llD4lqt+flTUVFBNUeyEvzKbOMpjD3RvxWw+N4tzWoGktjXYs2LjFc+pHQ7Tkjqe
xu+uLtlwrR2CdqFxCI5P3YQyk1nzJDczlCIDHSdYBL2a2SQOgedceR9SGmTPAAQy
IeX+ssTxZ7/e08tAGf0r30Fv0/LX3wF+8o6KaTCCKGoKu60Y3bulEpbFXJUzzHf8
Yi5ZC9odjn7BKsJ9DVLT0Cr82EfsTRsYPUmDeuJ/qNLazjt0arx94Jwi6Oj2G6Nz
EFhSHZ8SGt/YCHqjPC9tW05IoS5i05S5Zcs7StWugmr+A27/82evXT2Vvv0+F4Lp
ctqpdPS9Zw51sIxfgTCqXYSDmxQKPHlv1G3UVX5mDZ3gdxhle48e21aLFwGyXPc5
M3waIKjUaNysZGu34w8u90lGX6gb5cJFj7dmSjFLRYXkmj5+MBUQT6B/PRjdjuI2
qnxySTzMt/Q+tk7DatIdZV6BX7o34JU6ofGu2fh5OyF89AqUZjVtVqJx6COlEPyR
MUZESdPUNYFifL5pjnSIlfpvq5tgZ1MrIujaSz8Kb9+tx3+pgOjFwio+TrO820Hn
P0XH6m5VTFNCm7wSfNN3MHKRP3cM8WuMvv8lVY0kuQTI++/ZxKZetqQe0HkjisBd
zRfQkQ2YqloNEF14nkf+5PrFe/J0f8jNM+DHxuEqqbcb4jCdiz2Am8lPT47VFcVY
E7N+/qjklagatkbY2+D/ijUtl+/hkwlBS6NI9U8NhXjvt9DD4YPRmK78OELZlKk1
lAK6lKdm4ZFhe08qYUljTSMxxEB5jG5EZBMzP6agnKUHwNEYLmdpjdimCu15bvYH
MactqVJ6BDqS6Nr4+coIZNPXt6ObhR5itV/kFXoFMnj8Gn0vJD4g6Wi2KfVsLvQJ
PDBqlcTD67Fslr6PeZADe7sySwr1n5gdNh6UOkdK2FjGH//bYZZK8I4xEj/JTe+G
orZRzESwlVUfkLioJ9UXyrAB++IEI0SLcz9Z7/0XQAmqI/WERZVPSDxJo7WCKJ72
3NQbkV9DTd4bA6cJDTPlgfYZ19rKbnL438Oht/Z2fQYi0FmHTOW2CKFEvhh/sUzR
r8mvCiJo8gCmBH+JyH9OQySPDUqa/zbBWX8IrFHQt+POwP7FucJBhbz7GfXjuOe8
PprNInEzavQ04QIWjHh4t/iTdl4EDlQkm8ta7SqRuxj72je7QRUcL/M4cRVD9aLy
jQp9Ya2c3FQBJRr9N7K/y2xnZcMGWwgph1ev3rugX5ldW3/23Bgqsdu8Y/ZweUHV
PBnX2ycXBE0VT5JLGY53/Ja6Eiv6uMgC+aNgwlFbgZJkf9DfsxVgW7+0x1gaecEs
Qzr7oQU+uV4WVuwUnRLfllN0QXBr2Lfl+St2yH5GKcYawyGHX1zqK+hi+6n2n+cH
jreANFS2HaSeDVGrI5TzPXbxesy5OUAjhQ/M+FOu+5vF4kujc1oHquq1atMuIIy4
lkvThgQt1IVAJRHwTj9LrMBiYNHLW+p7KejxQydZU7IT9Ym+Djr4BDLA7S4aSqWj
/Hh7Q0n0KaVC1SazEJyaxscWrNUiXVwfZyNN6ivglsKe7m4YBHFx/gyXJZbAUGNE
CFOOPle5gkcOuH143jP0ktNUFKWTeVtSvDSWPzs3SUtZp82Gkz//headLz5fKkuK
mFyGyKS3Ig/oQdn6th0KqG6KrrMiBmCx+Nt2NioCQVDbAL1T+GEJ1Nsmz9It7G5k
GXpcfHlmB5fqp0A2KAfJQxaUaE+GHRInt3xlAGkkg9nADuSReJw2DXvLNPEr9O6H
oZvG1QUWROViZx8/Ahvs4ubDf4m0UfdqpJoAcW5gPqcEW/EPqHc4g+OTXjMwlKyz
VrGcJSplYel92Uk0CaakLn4qMRC2U/tfPjuf91LZuYTtMhJpFMw/Fx1ruP/5SEdt
ncjxWZ8C9xx520DkMf65eYQsV/iBFcSooobIET3dYCBOLuQTHAGMtT5/KLs7Vsw/
vwThxE3ulN/0LbC6Km3Tj8CDuzWjhwv39+L9jB48VGJJDF6hGLAGTnofnqTlkjwP
EpxaH8J5BZ1DOSEYyf61he/GbUaOAUE7n4YFU7zXqVDB7MwEz8/cwSWoP2WSsOUu
8y9kaBQ+m7IUdF5VWqg9pL1Gw0E2DHp1W5anqOlzzxIasWBBttBb+RHfRpD0EEVM
IonSu4FU7akao/0cwYleEt8CJzxKHkA3NmAXT0gSAinsjJAs16ac6PHIf+O6hFSz
CxD5gVqV7+bzOhtOEF2gGlOqMduXjuwX8FhK5lsdGrWiVq7NDVDWInJtV1XFGNtU
fsMDUsjZf9vQGbpDRIroAkhEjNIkIx7TImyuorv2FXPgF23WmAX2T19Zs2Mm0qgS
dEHhDbMdKOQz28gZ8LqZR+XXuw5DUYK320G4lX77RAU0rcKXw40qxlGIn3X5ihWG
D2mz/f4lCzI/MgXZKKjTlkwZWjU0VdAYZRRKE0r1Txp867VtriOJpLMKCXwy7O8x
XY6u/8KNxaPjaEIuY0Eg0i91rDKfzWF1C7RnkhpAKOJcMTyv9OL1tmHBA5Gt+4Cf
Fh47VoqePrOfgrGT1LWbpSXqxrCEP0jwbWytxstQBTrbdLlD5M1DeeaOWyYPTN3i
9wrEe5qScO/k5XO9c/5AfyQAffuveGHzNbki03+WR/pjucIMdgFmRmQyxGnFsa0s
/WmlqdSTfGuQ5dFxWMw0pnHTVvmzx+JsusuNw4UjkBaZ4YWb/7AeVd7kGTDj8/qo
lKCI9CSyyjEKj2/la0C7R2yO93g+iDFew4glvtTYQW2GTAOU0S9rjrEogV2DWvbd
nzYKi6XLT/qjjU/pE/jDq0pfMfj8fMl5SQ/gy+zueaoauQfZqBxRTMgs/k6f4SGp
aRwAZfJo1wUZBFwVxTB+mzLhC6RFZbK8h5XmTOwpnBoAG1bVadumQX+AUfWoYKiW
eRss8Jbpr8cyhuW61bppitL31y2qCrQel9Xkr46XFewpk9nOFVWQ0uazXzqed9R2
gpXh+Xpydgx4Hy2Dqm5VKQrT2386pJRjKPYGULo3yL3nAK9oql+hag+rl6b0+Lvs
0zlSs45hoJeKp2B0W915g8X9j9B300Zn64cl1/rSY7huqYj6UQKme6iKITT12kr0
he7IHYSwD2c1ZpwfZup8BvPuZprzn9gaJcm91HJ0KB/wibAbF/5MRf8DKqC5c9P3
XA7lVO/8wBf204QS6jVNT0slq46gIkn7iKClhSNm8GG13icM2APa48RAwlcL6IAt
SmFsZOOCzJS8CHxuW/tpSo9FaSnWeb/c8scHhX59uOnt5gD6S+bV4QKfdkHvnbtt
3QJWCqQmt/Q9crHuhOGNr8r3/zay5sIpPZFZm+k3CTP/Av/naLIme+uhtO70vpq9
qS0Qd43jdK15xRIjVYJI1NknKwbA8+w2cWu4d3VYQl/qSWt2JAu2OQYFLibO/N8p
eI677eWTYJaX7ihPiBnoHZAo5D1gy0hjwTfSljUEiZKsycsCKn+hRFcYzsDjwrPq
uWtyjCxAXJmLnjJU1TZSjle/vvQbVm+lT5hqb1WARahpwXB5FEPeKYhlgC8FBqLq
BaLfdFaXy3GsyNoiZaNsbPte12HBI4JawX4NI1zcB7RjU5nIlFi9ZN+kCxVO/Xpv
jbvfkG3g9INiRPd1uBhaBZ5K+6PazWxXOeMOmiuaM1hqk1wRA7veG9fzpBSkUJML
9qD7hVfZTaGTe5T9bz5oZ1uFqDGMvjcaUlMFzOQDH/cCBqPMmSkQ1fRZ9KaMDvFy
EFyzi+uHlseTZDkSU0DSbnFGzUfHRYttew4c3Cf4l2ASSPfNXFnPrm0Z6NMb1He4
cU/K2ELws6rt2vZiqqjRDfysIR5rUI/Hrn2ojQ+uZc28fIrUe/70EVKvpoc+m4EH
5YysORHK+Wvj8LlqXRyiC3QoVucrfCM7bfUzYNbFMYvk4tM6KnuM3uN64Ej4H4vS
YvQP6qZv0IdJP1og5izKAyaU2e1RSMTltuQlnOYxFUcwsMqlD7tPgkaIyLiFSP3L
YugH3fw+wX06qYOBvTZ22ONBlyb/hQ6/rzR8r04SI8SiVqYnk9QwVwaGd+iLi8JV
doOfMHv/hlfEux8SpvjXbHSxKq7Br7Kdkdf5bi0R1mnAg9tHW9737DumZYjCAn9V
b+jTBTF19xsJOK99+T5dPLAG7qLVtM3f0mo0vLGO9P8dTUoKSg5ujhtNMDIoCRsV
Pk71tKg0xtF1UvyQS47MEmFr+YmKl4AOHQIJXHrwUDAtAwgFSIem0f27KmhzLwoR
NIgxdDosAkxPF1iN4wU9kTjJgLCRHDH/EKR4/CCAxU0EK6nKq+YWMzKnmsHCHOgC
urXCFecxBfDVV0wtHNY6jqvGn+GSsp8AuPEIY1LNhoNJqYDRQv078ou0tYTXVcrs
w4YP3nfIhdOEvnlY4xhQJHZKau3IjN6znxguKM4HqVdf9ztO5VwhvohxNgqalmkB
MLdMs90aW3bfP6zCkjrkJgNNRzXMCtayTuvTIWGaxMo6b7Y4QnHfroe8S4ENUhHG
f4jI7dN5jNxe/olzbuoKc+0XM/U81zBA9VdF707KVjPwidYpz1BswwEB5F1ZxwnJ
2rtHtH5JXr0iMzGF/YoYTAbO6EXCyNhADcKr+kLjSg8RAvAMVwVHd6tu/SujHPa1
WktwDYiKxpI65Q7JOAqXN/TYXcra5XJltDXhObW+NQSHe6WBR+quVCdeLswpZF0f
CZp6REqlZVh0LCxgjJOv3mKDfix4SlpEFXIGnOKrnkMPIyIKQanuGceH8Jf61SIP
2X+8ipzNMUdDt6eWRc+w0uKNJYtvDNbMNtiXDTIBB4s73i47yXH6Ti5GnbUP2Xjn
q1Li/BHGW90/Vavb60jlfC3Xa2NVvdkCWEnAw8Vr8/YLevUuwkvYum8fGCRcpjqE
wwTf1nQdMIN/45KzF2SS35HVTSSkV6mbw8qrSKef5T4N8zzuGZsSwAJNM1Y/AtgK
IHRzjM5n9nibO0NOI7JSsIXgvywOKYsPhfcBoZHnplEzaLyCWUFEnCIcUUI9RIjJ
Hh5RmSExtIROwIczRM94Rz8yW9J6ARUJtGv9HpvHhDqiNXKWUOqpzjr8pZBXoCAD
0okN130gdnVHKfT6b9McTOIdty3Kpa5hjiTpGA3e1EBemvoD9qNe/DM7Xw2jPox+
xY4YwGiFn+F9I/r+sSHzFGWO6QOxAZvwHP0JR1+RjrQgs/j0lJQDNhbbrryMgMM+
Mf70FVha4GNtiamPCYFqv4Lrdt/yIPJ5gM0ofaIfwBaOK1yEPgs4hEQN2aLbvzfh
107YiQzr7/s5Oasc1rjgw41Bt5DKIQNo+4GxzZe1cDIrXo15jeYLCwFHuBdR/MAy
NVq8/8m4t0NhJTNPIr7B3r2GtVc2kDrW1w3k+IITx2WBHpWr0OT3sG7qm8cqRNPU
p2FWBK4F77KFRl6yEDRBLeRVpz854+a2eqtRmAcOrdUXg5/UgeL5qFbnVFcEwQFw
rUjVFy0OK4deTfg1V+IutStibibndqDMdBYd9xMrhw/pSF/dOrTryl1P8n7ESNVJ
rqOommgZme2YFA7AKhSLnLSvblrBodNHL1TtAsICeHXkxodjiFgDIhpncZADIbbi
2CoG6oLrF/BLCCfA+iuvInyG+wNpP6xAVnfveH61wUV9+wSKRZ5wF5ZwSgGkXRdc
0+I8aVgKjacDOZfo8OC/W+6qKYO1wgBkTsNs2uXOWVyP8mVOvEqrodtpxBSFH4QC
ZeNtvDuLbOHgD7tjU1Jbz9JEXWcbWfewd8fKOSwNmJYldO3t8iF7BvrOKT5L7fGP
M384jxEGdljOxQG4VV6j9+4DYiSBHgT/p8yMMHew+lqTyMl0CaX3npzHZV0mpcx+
j0pqVSYqmOp9eb4/ECJa/OfD0eWgIJr5iMf+HvKoAdyDjP70AdFCID37hoWDz0pr
JfvsSE8sqSO3cZsC3Rcit8fARouD2M6eQ0cN8A6qXjyDxK6alQDAlqJHn9iaXYEN
t1Kvm/aNmVj9yRCXbZauiEkRD2c/PK+blb/dsexvM93MbBh/GoJu/3zEmTiqAvpR
McHBB6/vld7I6GrzQTqJLUtBFlh/MPQmVQysUtlG48iT2Lai0aX3PZe/p9dWpouw
uJhdR+kc7BI6wJ29VjquGckvm7ir1hXpkpKdtB8lOvCLYwYIA20jDXT3Qebqfol0
jmpTciKX0X0G85R8kPG/+Glq0y2vahitMRpgOSd8+OczBffRunl7D/ig6fOfOqyB
oMLEPClqFpsjIExOavQfqz+291cbRXBcwcIBWvyGbjsmgNE3wl7MfE7xNbYHdpdc
nQxQ9Yi0KSJusJfZZ6yCC/P/H7P0oGLV+tGa50/3J0x+oGCK1d3bJCQ3kkvQPyDD
XmQHNB6PeAJkQYtQDQfjppeBtY4sZqil/X1yp7aPp+I+SzWznNovwbbZuW0HYAed
v0I2qdSTMfHGcfO2UshDHDIIbsjTi/vNt0bS0/gEkOsmmtG5J96KP5xZ7ZldhTlq
ta9+glrlkpJTnfc53r2pqhfynB1SKYbgyf7TZTY0oY62n6hO38rpOHts2O7Z48oj
eOExzTz8Pk6IkEQIpIrgJQ3uVLh9Xf8PCTSzRymMZiCBT7pwS9WTMIox8b1bv0MF
q9MvE7kAt5kjyU8wcVOuiraPls3CxQ/FKMJQ2AmsgmHnVuo4c9VIVswJS6ddMzqJ
q5h+QC3zXhkmAxDue2s3Co0vXjNMzEO6uC32mZ8f72RWsrrzlxMGujAwwvYW38ya
ji2ewCy82AkNepr7Ntt8NW/LJP2J70o4z673AcOuCvbnguu+ALZQI2CgFFf/vjIm
ElMBG1208V7H1ooQINQsYi2bkxiD9DvbrBPttMOmjIlr47ySOzAus4/iBN/u1pOU
QLozsTN1SS4KViKhxkzP6knPs/6P/aOwIz5oRQGaDmFYW6L1EJeBYbxpK6iVZMXx
tBGsauJugeofXi0IYWcMZGB7rBv1Ai8C2fkxvAnXszBB/guJ3V8u8qD8CKQPuVLB
UsDSWJw8PoWzZr8kHEnMvtSw19J3qp1QyxoW9CSpWJV1bDMHL8jLbCQboNqRzfXT
oszwPQDa7cKYdqoVpY9Su2Js/JwLF51Rv+xzftlemA9vBqqqqxnL89JjHLBhoU1V
85QaiJYCPSbVqlWxy57xw24K1QbVkQOsMuFtaccgrgsGSy0ZjTms+a5O4xH2wpGA
tRvh53RxarCORGOoxW931oFTQ6/Owp96+PCPVVi66gY6jHKnoR9PrhFuBJUfSzqb
SSiB7qa24bSiaqRh+9Ie2a2wOpUsFYn++d1f+ZUoC51WAApqwSHBHOd0tCGOmm8h
Y6PqRb8je3pQazfCWD1kLs6Uekm6FMOW+VUgXwY0MuJASNH5EsAqjY6VaRlAOU+B
89g9caYslclfNQ+v0Al4xOVhKHQxoSQcmaJL6IaiV9KeQrBqJnLTm7NhXErvZCEz
O5OynsvNOAR9PdQNRlNCNDgBii5PI/yj7HHT6Z7ZqGR74ZglOVr6JZGotFbJ8Wac
apKiaEAO1O4mSSyJLohPL6e5OBkDiOFRCJ3ixGTlPnUw7hPFZU7ii47T09wLNUKs
btmil6bhkSY05q5AxICkNkHSk4+din15259Ry6KLrYP+unydAc7zJqCGMpRY8KVw
cSaGFzY+InAgEqydzD7HZQKD9PEcKM7/yXOWmu7mUzOT/P7j30hJLwR7mAd/Goq7
ZFFAz6Nq4VepfupYYTVdkVkYpclj2lTPyL4booUMMgiZJ/YeTSUEuvSxDp/sxshs
i//9UyiIll9SF9DCzofiPsuGH/iCf8eWPwMCm5jS+RBFO8YzxcnETfYvaMb2/hWk
SMcJbA1bZQy4DjOWWtiZPASl2zjA+vhFHtilrKVccOMFQATACVPtODxvAwYuFqRJ
d3SSlNaaRc1l79eNaKHaDk8rOoJx37FpBDVSel0ZJKTVjO/D8gjjxP9dWUe3F3vb
+1BoITkGRZ6IqfL3etv8Ne/VlNl0Nn9NS4CFh21wwhLm77ZXy7Lt3ifQ2tshOgO+
RGImcUE8HkdHMx01VC6OKos4frktUUhSvLXS3rcNGeMxHB3FZu1ijSAxnzgn1kiN
YkdIIBzm2YvJc8otYEqZHLyAEsPSyVtItKh0ht09baSI5yzV9uBaInDIbLjzCuTc
jfluGyDr+FbShMQDrr6NaZnzclNaST/FRPM9EkCyIGJiTUTElO4cD1I+7MsFfbL4
kk4iTQ10LtTjl0Oxw+FJDpsHyRvmnvUmWM2n7dfUjZRUZ5A6mhiRiXtyx1CLznZe
ArmyyuhkZr04A9Sh4IBoiLZSyYDBwyts4zYJXyk4clpvy7GIWEn338Czi6JLhkke
YJHTbTQ/qM3whq8eIW0iiAyq8EaY2l6QXyq9ozCNhGGGIBYM0On6M0KZR1eZxG+w
OBh/rrzXvIIGly4X65pkiXBvJXygOlImC4V65rDQg0bUEAxA3OXRGogZ05RDRCBp
HqvKJFNv5O8hYuFCT4SDGSBR6SHQoLTYbLXTfkOo5pX0j40GMuukRIIPGdVa7Emb
X0vRA/vbjmCI2K22D4kuvyktCi4Sd1NMVZbJ6xc9HkOMuGw1QAzfmBgF4g1hDQzH
6PdVXGXR1kTge/m2MWcyXTLhkgTDo5ZXeBnaLwioBNj/y6/aJAVm8ZboIcda7yZ+
LIGr/9e63NNuySVumPAz+p+q3APzDpH9Uz8IglSwwTaNb5yta/SBEDU1W222gnem
Uh1+QYswGYVaXNuindUwPVwK6gNHx+jIW/Id3cHsmeK+KqzSiNg8elw3xzadX+gG
8Te7B+nEKQqqF8fU9qy9+sVn2J6+PMjveL+AfNIhJvBt6JVk4MFhqHs/I0l+QbVx
SAzrtfKggmY94jbOGg98derWM9+0ajTN/1aB2+C3cLgrLmspX/PkrXaTySKQ/cod
nDVG+2zzcPxJ0qNiaqzTPeRvt9urrniUzh7sxxdRJlwfLSUUKbxadjACH4Pmaxc8
XuRTdxP9bgJGX8MOoBMilVlSB1VESdrFD5To2lvzG+rsyv3WEvndmaePLImjgkP0
lO4ODcsAOatHh/y81aaC//nt96dfHDNWj96q4toJ5GZBM6oD2f1i1qWf9CAZAaGq
kR74OfCHYAmvYsBi9JTRV7DSHxw4cBI6Ipua9MoQ/ut16V5hZiYWj15iI++4z3YF
2v1n1cPV/n0tPcdt5eD1LxDVG0BZzfii42im3LsFsWW6dYsFhSt5nGPdVmxfoVJq
8H8STkmCCjykl97AXZv83winX5wrcpaSy8qRZ55qXJvnh/gFle0cQ6/Z8Y4tD5HD
JOHtSkmf08xV9OwuSC94NoH6zIaCPwaJ+tMi5ADBksWFajdDQPDWhEpPgkvgeWxW
dnQpFuz6QOWD6E0jwACYkxCAcQn5kJYkHLMaHhIS1dXNOhLgtLehyZz1SaBCLgjW
ZVgnsb6IfOENvFaE92Dzsg5RemT8OhmXDs/yvV6EdIcSh8O2doWtcV4VOSjLBZbT
tNEbnOtz3IAnsrETVu1C3PEvbvkFTgaLnkqeZzPMzfp7q+S3g8oaQBF/KZsx3IIj
F4fmvsK8yj4LKsiSMrRxvrqbLvepSZY4JYrkw/p+0WvhWc7AzV2R6Fo71VWnyFwK
6bhQUApU53/0By4TphyNIKhUnZHqdv+1y95mHFr9S7HgHDIdf+esF7M78corC0BS
MlLkpVfwunN9YGuJOiH6piVHEr4VYXGuAzU34sAL2KPaidfUUKHe0XQU7TnMiNMN
+Ms6CB7VTvLQQ+nlTJzLqHyzBJgdhMex6BZKH9YZUxRvemWE7/RRDsZgJqbcOKAn
NAFZYlukUT7a0UfzVSno9BhqTvJdyGB3Ylwr76bEOaNA+2x0BSUf14zsOx3Sagxk
8EJ/A4LcToR+R9uisg0ddpAzkpU5p0TwPBqkbCugVO4pWMwRGNtHVZq1nkIl8JV/
iVN76NHZAhQqtCdh1lJ+P6Ap1U/9RUix+oYh9RJ5//nvEbfp2GrnfA1i53RXWEhh
7dFqYSiVQLu7RfWHChW5wrQY8cgoz+SgzanA9EYa5ENqpnw+cL4vUqQokrocdCsi
jNcTC30WF1Bt2iaRFTtez4y0D5OtNZmOh7lzjtT63pkiLGoeUSllSmHTUxMhepPN
msiuYNq2YpxZfJA+2NK/fO3t8XC8746FYT3LsLvo4IDq4kxrioHyN+tMr9KqhWvr
JAC0GpOiR/LKG+C/f58j3WR34t/qYG2gm8IVWUoiQkrncx6RqKyHbvLUs+4kW/i7
QenXogXPgxmum0K0SkDrAifi3bV8oRPUTnGERpGXHsLHVeN55W3i4JZp77L+9qzg
HAU5/ZrA3tkyC3TGZ6XVh12tqHAs2YCYq6nPaDq5Q/thnSbX7BsI+TsIKuFSGtVg
00FPcdPguvU1Qw02PGCxNb9Uxs8sN0pZ4OOPgxPusAwcjAK6qFwngF7CswfMlhdM
9Q1jB6Xrf59PPpNx9H2HRBuZCoQrwDe38Pwfc9HID9u+1M+Kj+u57WnmDCOMZPy+
rZxf/+hgz/X5S3fggPefn3Xk0txhLkAmpSAxmQllUlJ5DtGEoA7S67wdvhKWdhuF
M1MLbrn+9UKZcrUr688W0orD3jShgMCEdU4LpeZoXBuvoeZU+T50t5RSVGBj27dT
R2zcI/KR7fFAcBmWWDFyIy+GShC6M1hR0Dm//Lf8ejpicg5t2YVeSoMjkcBCTiIm
pTp8Jn2Z6FxwSKxWYuC2dqXi+5mEpEm8iyrFyGpuXnG9hnWdWqqLT1JkHHPe0XmK
JpM3/8/YxH3QZ3hH4onD6bzdr8TR85ifHLD1IW5/GRvrRIVVbOQ+vzIojXspLIc8
kjYzxrTgn+8Yq2J3PhPMV0nY8niOttGxKxGHHtqeLlKQHiWEFdqO9I6ecavqcZg5
BxGCp+YrM/lXrPaGy++fvP1x1oLEsLecDKVVP1hik5jjJl+FTXzT4iL63FwAPUsk
Xd9SswOc0P+VUhLxrai/82mFEimHdg4KFg5GPHOKNy2YP7YQBsXz5rP+h2/zrzOc
muyR3ZjIWCuWxue4DTxow6AeqDMOOjK6oLX+d1Aj3pfewPZ5suAjsAkomTFT7g5j
H8GdLwqs65aPP5ejbSzLeAXptGYDHUFfTIItQGfvhpbQo+WuzhBv4GqLNBRJiyx+
lOY3Fg8jQzK5AT1rKuVosCIL4Z8M6bg8erDjBdCSJmh/WarRK44Wh/HmNVGsS0+p
34btt6dZ8jDiyZaX1RYEJqRT6ljV3cmdrtnDj9wR8mZ8c2O6eNrLavLTKsQVIOne
CNqPL+6Wf3mZug/yrxLd9V7NV5o5/YYP3lrhObVf0KhcNdK1HDBtteK8mjbi+liV
nk8MuFKc3ijzjfypWlvYgkurb7fSRJqq9spVg0MhTaOiq88Ey5z2z5q9EQsc7iAq
z4dzTYL51VWguG1G0abOLOElAj8PABuMBR0tHt0lqQ1yI40BROoaQswmqa5XYFbK
Z5kVuGoqjSemnRhyACqYipMPEULUkfyYg73uuS/PLGhALvCHURtNYkvn8NIv0pRl
F7pYIPRz5yfquXPcm/2uqsG3TIZGk8bN/WOrRQ2cV0z7llpHzDegHPpmPbSyDgqy
+1CDZW1GwCyaJ5R9XWM3zcYjKMnsQ2k5Vqwdd+P5+HsfSmeNRHN1UYIoToGkpxg5
m3K2xU7SwP+vaxhWRjJu0eTkuIBqyF8lx2wO7qBBjXFZMJtzjMmfsWwg44PcC8cF
Og3JYhzyfSY/+V85QSUaEYIrZ1bnmrA7XU1e1In0+jLmYzGcTqXS4M8VxAFIrzvN
J0Sz3IYkePYAt41HXUcBnNqkKA36XwXc7/iGLXQhPYlkHi04wOQChhqhwzB29FsU
CNvlKejHSVJMKhImH91cimRxfHScrGb6hCl6ShEf+4PNlX5sbMN19XFZhSVhIMjo
RYO0v+iyKBshGltn4fsa0DdZCH8Eo9uhYScGCorlm3rBk83NQ+wGY92RWjK+78xM
fUtm9VjOzyVj8TuTYqNQ6C2y4zfTwhhZlHwJ4mOcpc1Agwxn9Kzd/F0Xf5SY/DXm
OBSWrzqvq8e1ccku8l9810Yyht/0C+DuMhc5lxY7wGJzlh1ycZLeLBJm7LcBMpRO
k0xRQ0cr5SOMm3MbD004ja4Bbyzu+OJVcZ2SDfmdlom636MYgNBnYHjhz+MUtDwq
us+VWtAfgyko7IhMSvFAotlY2ABnz+0Liu+/WWS0W4jdwrwcPeYwylSIhD10X9PB
+pynoB6Okd6yw/zcI3Nbttx2Py2iE8XegBuGahMpzmTDO3LbO41bRn1hY8TU4u4N
OO6xKmSdn6junnTWkVK8F06qFcXC1C4vl5BIeVPXecYVPfdeIPAehxRGOyW8hxry
xw9E7dXu8YacmDDe+cWvTMO8bpQhdaygM2W7ghG6kuq6CEaX2BudAsJ3KFz9Qzb/
Lh9BB5GIVlQ7Ph1/A9X0+TEGWlKeheKsKFhxQNtnw3sk5fLmKhZH39jMGpFDUOAp
/ijobGZG+8n2TZTTaAFkSc9smbpRqikv2Kum87nFVnSWiASt6VojAKphgv9ZW8t8
hlZ9roPNpJUJRVEiXp2X2wcY4rSF5rWrXizC2fXBthfV8/ISeqfXDXGThpAUxicL
x7ik6fA443oEwOyX+IOEoeAmArcqqtWdM1tXsKxEz4yJj+2+R/au182+nYonJkaO
I6yPHaDsigeoyxf9LZzWm+lry/ljJb6d0Vky7NnpoIuZNd05+X5mWvzkv/gpKaCm
KithrDj8R+nra3y2RS6Alk60fQQ+r1amNfBH+UwvAhUWwJda40wHDrW0NRzZU9ty
X3j1HMGa4G28UOgUg9dsEEdtQ9otGPT69Zo0Qp9dS3xw2xdc9/rvigatSdXC54Nx
mp3UTs5FBISVb8Br3cXn1tIEicfRQcGQmNWM+39rzl8L6f3GhZHR+qffxTwUebg3
591XECZ9tZn1q460iteZLonN3Hmhc6hWtNt5gOPRJZHQtC63y8R47V7VWj7X9M2t
OCKB1l55Uitr3qAHt7rQdjB5FmFVhT3v0IBwDpdwt240XWgP+6PUR0XRZVjv7Mid
ODAM/4Nz0FO98OE5P8EDfxzIMR+gf6V8oEJaSoWL38wNoDxbJV9r/+pYghvryBIj
MLQMOoHc20R4BuoDieiOv7ROOWhkA1uLuF2MYLXecFC4SyUbnQtcL14nQcvm1UZ2
9IljNufYur4XTMEt5wSRRUHShxLI3PGeKkonTeVO3btoCZR/ufZWb9RCdf8ZJ/Vi
hhWZfpGEPO5T2+Q+m7F5NfILassaS9CqFWdFWyv9o21EM96NZoGEAAHyZbzOKHjg
a49rLgN9KUTTZHrQkeWQA4BtLOgRqozQlyoqijt5/OifX5H5YpcyAJlTS79g3L/T
uk0lB2Ns0FM3+6YY9FQmhoHmpufqDBf1hQEBeBeOVSv7D0YL5ME/r3JEMqZyEb6D
0Y40pcw4LtkvsNkmKrKMnddQS50Db1m6WlJgI7/PRXlrMz/Fkm/I+t9UoELjBQ5X
+p4WIgiPVwOWs/AON+rBjq8BrNAd8c4QL18DEwnnBhefltR4Yjhb7JFzZY1p45mQ
fd5rrMez0gMRUW0vDWNO9/+AYpTZvTv4eQcKJcIHYY8gBy0iMC8UONYnFgJZRXQe
+Toi19XqJtti7y2bIPo95Qfo91yeJkYzHz+c2V5FLshkJ+oB3BC5w6gw+od3mS6h
QPaZyNoVGOwxUKfwRt4f3u+U2BZLOgxJ74ean/k/ZsAExEPBcSbIu41ra+Xu85yZ
OlaGdCUYqwu0leyTv3wT3b+XtdsCD4Iu5Zlr+/tRQDvbkoh286A6jRcBHfrRWIbY
aqX7wTLEIlbjsCM4ZrmYcYFfQ8teYIj+0EessTsPLwEIWAuWtTzdhsmiCKAZXfGU
Sne+zhLME9q8jrGFaiXE3KlK3Bn9MlPLBlbR76+G4zkd1RE85oIWmP/tCzgki6jV
s+/wmfgEWMpQBQwc6ynjAOWN8sYXZ2h/rkmh6YGG8FwNMOtKa4lSG8X2Ut1NFuW8
lXGd+rPTiAXwWgW+ewWANpGJrOIuVDz6vpa2L7KdoYarJbXC/tsBPCM9cJWuaS7Y
Nz+5l/PPZN8QvfFnNBkSKsp6qvfCnE/6rTwwoWYjXkuReGXEhDQd2VASVj3zbusO
mA6luajp0fSZHLdvnhu7JuRIKaZH2FK4ETp9n0gXb16NXbgrv1R1A+MwygmxCIbr
I38y85zNQKJEPClnUUg2F5kEbTDDafm/VfVRr6NuOYH/3wweTeSaMX+7QQHSCyeU
mcWxTN/Eq5Nd0ii0VKcPRBqQ2XyAy2iRGdlUtdyw+WOSCdiSmLSzKASruQ0AbkiU
c5Xd8MCiRSX9mH5xFk8PYqw4F94mWxEvNpU6raVnFq8vAMxWvPMsr0lzCxtt77at
I5Uh3rTpTElkVL5mtyKKsHw6loRqKwqKg0UwVqET8aIiRJmZlyBLdAAPEvtg8pTI
tL6UhlQYMwtoAvulRclY/hbjXeK6ZBYtPDC65GyIRTWoAMfkIMe0hO3QwOvAd7/g
5QJHD/XgMNPq5jaVnJyK0iuyqDdl8VYze1v2Az+urev4jLMLHnw6Qo8RexkP9AdF
Jiv8urYJTVu7zOrLhW7iQ+Eg++Ddz8zPgFyJxxFF8GDH2tIJX0A5AVX7A3XCz9wf
J1qXW74n2+3iOPaRDbm0C2Km1anJWGhscMqa6CmBREPDSIVddKtOWMahsVa66rIo
T9G48TGy6nbdolfSU8tL4Kj1d7cFHXcKZSqC9yei0wNTfeMuqLnmOaP0Q7pXlbcD
6hM2eD67cuxuCtkXrOM00F0PBy2QQpVCxgcccFV+PBY91YIaVsCyinHK5lF7TwIk
ajOUTvSGsOWG0hS5mnaPqmvTexKEdLhehF8zpZiHgaTZVgINlGP6tdCuOU24Pfx5
SPXfaSyPjD++WRc/+CQYK0Rh3tqczThyd7Fy1JSPj8ZQCJsOXw8ngujpNSiLJLbH
LsQu4zsKLGKJ7UuY3g5QiS+ptkDl/aiIO3X7I5x3JfSO5ERzlTWNXVilVjq8e18I
e9r2WxDudNB1F8JxjmJbM+QoHF+Q/PI3UGAJ2WztOdsnsrSVHqDhNAzBQM6zvszk
RRi7g1Sf3lR5sW5ojDXgNsfB36H2wFvUzR3C8+aZxttByXNnL/kv1hs3qGKSQEZj
mOO6lhAICfpbH8NxBBE2rG1fYkoZllD9cohjQLB/6zwsBMa1G96eT3ugAnN8HUkh
yFsMHT4RjQHSkDt3ATizlX/Te7FO+WiMRlhv63/azRwohYMSUa30Pzw4XZBxf2pg
nUZHmA3IfnpZLuYcAxKFzwkHkTehk4POXdLD+1f4VI9ofXCtYrUTpVbgOge8lTZX
zSqq9Ie+pXWn5El98UOznI8D4BgfD0AuIg5nKJ0FemWbz1mYOQd2VDcFBdLay/3q
QSx2zgdd3ubZHepslI/cK2CAo+yHJgsdSSuG3JkkoPyBKCoCnQFzO0UvxGg+t1c6
N/0Z9J00Y5YvlLoSrHsNaWE8Ivtstuq77lsdQpoIoUp82Do1IhGGwpxRLaG0R4Z8
d1SSHenw5RVWoPAJ+hJ8ltTj/aKbWC45y9fXvHXrGewo49NXbK8uFA6U4izPP3t0
UzeI3uUA6/UZBFw3I0Regrz5K5MkPNbtIUzkzdZ7NxDjBb+AOPQS+xQ5SI+C8qO4
sB6wWsXsPE07C2ibHbjnHicK3Ghy40INCnMnxhDuZ8mYZsz2moeL1NUnhOnRcb2/
vavOeWk3Av3zd2CU+RdakGZPZdiiK0gtFHinqk1gAyXyzYpx3T+BGNLdukegBsJ1
8zReJVRtqoo8pGbi5tOTWd0M7B2k0V0Rx/feOqwlmvWMC2PRPvv37FeZmwUI3uWn
TJiD0RwGaV6hb34xueyyK410gOObd74vZHLw6ez8IScNapgNlsHb92bu7MwYUQou
+6TBeZ3j8wGlNSGaIbCtfJ0cpxEZQC8YwfxfE2aOZeTmMLRWuvT8Xy7jQ/RGjL+6
QpQvh6UysMSEgFOfCtjW4JfCnoZD/WtXWgzLPLs7JVeNkbIDYAmQqh7SRUUPB984
VAWq99EbhVSf7Mo557fpm5tXg9vBklDmtYLyd6COdLHf6KIUx35l/RA6zMpJgi8x
48mASiThTf+JDHfaRa3dXQmR7ZcwsF5V5LCcDiuJlTmcLufGB/+g++9JRGMqUuRy
ANXgYlv8o8DGDRHPiFoAHSbM74HwkeL9JQerXS9TGZt+8FMifnOR2qc3+7WdYj/2
dknPaPYypJ04xs7hyNwFsOcbVWEnREaMJh96glPJ3je5lKyADZMwzlEEINErpu2s
C0JbKzmI1FuAr+wxUwBAhDGsR8ta54GfhkHfWRbjBXyEXt0cllrAh9BwCrRbgRmN
ZtJbKvS869+CloHdpgpUpT43JzKc8TCu/nBMoVGmv8V/GY5xKQy1S8WwsUM+nfLs
KxfI2l19PkF/39rMYSS/dYRLU4aFFWHWX6X+uFnytRO61sYOBBM3ABzATVqRD2v8
MLDmRkrmyWB2Nk1mQ3nWX8DjAwbdbI1VjkYFYCmNELjmIKXaY86XlvMHGjZ8VUPb
d46tCdNo4e8BnOEBLthiKAsRzCXKeo1Udv854NsSkMaDpTWGU0F7ykyCAC5ZlMkB
GMj42LXW3Xf8u+h8bmYTheFk+dDBM3vTtwZiuvR6xYlI+Ubu1EOBKZkrMHjUt3ys
WtthLMbVRfm4tseWv80viO6nqvybWopksWF3JG1PnbZvfnLooaKrd/59q9Ze62t2
cEFDjXAgDexaYpqp7Mbi4GnTlnj62RhKEj5ziU3EcBhdlBWHBQ1rNociw4xvvkUw
pIBB6NfsYCotlllgyMwvB01QUOsGDJuPOyxnjgJ2OaPEi+Xc0n3dkw7zjNdWR1bQ
1La9b/DUsIPK6YPcj43SCkzanhmIysu7N7PGCiGrTYsUPejZkFNdgy07U0n3HPIP
eWlqR7PzY4GMZ+LiA0pBYFQr3Xb0dMslwLILQiCIO01Q/8FTO3jwo+vpVDUhikcS
yevhMjw8W6yJ3J7Wrhp+fHPn0GUBnBgRsNDB/+4t2n0kecfmG1beFXAxkc0VfAb4
cIBkXT4dLOu69NBHF47O0CQz7zS0zDZHSmK7xm7sSNrgQS4pXoDLlo2vjx8Th63W
l7KXmaI0HWfNmM2yyYurtLyT83ulTZAvtkLr7yYu3qVyUV62/tKm++3Z/KBsbMFd
k5sGA+N27iJ1W3mRqX4fRswUF4ONKgsD9ggfIE9ge9f0rsDZqI6pHB7OkzP0yGnv
xhNRWgw2Km5Q0qM3Dwzy/Gg2zSnBPtRdJf4NeUdFxXGw6r0VBIExqBqzeLgRER1u
QZ5C+mNMORfxAklLioKUoY9jrTE288nVR3uHZqznDauSNibykawjUgcEGKF1PFqu
7HEY8VOtWtGblivJzkeLO4Ge6CRfbGgeSUXfeliyEfEeJc6/sea+nU9FBOXpKUDM
2zIlIMhR9Bjcqbg1q7eg8PQcapKDcnYeHluuOxlJ3Ehh5f6alX9kW3M9MbsU8b6L
E60mq+JQk4JflYgp/GhAWspKoj/2/6A/u3MVpr4DvRGfIMFhCelwwPcgGaeXD6q6
6ozVNIRYw4xHNLaP/uwEWyFD9Bvgj8lSDRP0/x7USprtkqpu9hB757C+vFjenkcv
iYLYl0ADXaTTgccKrxeOIEmR2aCAvaFYCvCdiUONWPZt8ffsDeSDfwfx+1nQUQa/
mSg2PjnUQpGXMM6QAifCrsUfmpjk92M19VOgk5Nh0UPnOzaKKSdPmGd5G1JomtGz
h+apY3sBc6kuTe1czeBa1MS/UBGHTDr0BMkT/1te3TMp+2Y5lFlxAwQQOmYE1h8d
y4AabtFWkIsZx8heBIe0GFW/N0Bnh3Qp9pdhDsXrF5ggbxbXyEJJeWpc0DfQrLNe
CSQ1Yw11delS5gzAXnO7Je+I1ejiZphLHU79ehJSiur70ebn4EN2qKoxTYL0l6ZT
DYp3aDF3hGgwPjnd1z7gQGgbvP+7pEPcH3R/UAkXpVR9FNcgkehH+sYlRI0wCzow
nReHZfipnopHnx2VZ7CbMp0Pk+V0i/8t7RsJ6dA09rdr+2NvOgbc5K2Y73dnFHS2
IF3sKe/eIt5p89sVcAP7+yxv6q4IYLATG9bHKaA0F65SN8z+O9FoQ3IlV4whe0JZ
pb2r3CEfBdcWK7RcdP9hO6AFmAoDa0007ErPBSyI1L+57EpI5B6Vh0v267QQ+1Ab
CbjkeZ7TDEQ5Llo/F3dkipyJSHofqhzKt4LN6tuwCSv5JCcLpbJ7Ea56LCqU6cW9
b8qNmzK2EkIX1bp1EJrKehu8wcHRs0ZZkkOuHHcXtOrcR6YV7UopYRIc01/TaB95
IWytW8twuG0IT8TGfDyQX1i4qpLhtLjjUt6Kk0g0vopzrxB0F/QtpecvUAMwbT4W
B+bFd8Mk8lPwZth66zVbTr8EmzNaaEeYoDV2YWok2/XQhc69d9O2dpEWIPnMCfRK
JVOHE2WBHL4j5aRmZKzjDmyGv3s59PNHr46f4gjZ6vbKkllTDRSDda9N7+5480fv
nEH/j0+X9kp6fcDASc92v9TIaKm7RBFMXetnayxogMngBjq9AIQP6lDEJDYN9bWW
5AwJ6i04fUpLL+VtMRMMJRFAaEn87FWKalralmz2I6xpjpBQ6tz2iFoQ3XroJHnp
g/8segfYHt7CxJlEAx8NgFuRxO7E5oRnxzh0ft0ayZAkD0rE5RTqDZEWDv/jhMQf
mJMUeIS1Lpp1LOrwHjaOWxcFPL6mlBAcGEUOn29yI4v8S0xnMuAY/eTBY6SLv0ve
Viuwrzta+4uVYu0eQucn0dQxn44VT4EdskWDGIPuNcrJdarcR8uGz+W/6MzT8Rwv
H3II8r9ud79XI7fFiXz4y1TZ1VCdVgQr7V6K5lp0NnvmA/tU/N+PgvTAitRJbRzB
MxJYHMz96hnqLnNq2Q1MmnedXLCB5u/QRVwgSQMmg2fTleTsk7f95FE3Mvw/UiCc
k6BVL5Rj2uKLGPIRl/ntfkUBOgxv9GUIp26zV9eNSjO5jMTjR8VDAkuWBaisWx5j
zg9e1RQ56UuHXyruQ698dx1qB/rBE2bkQG2hUsr3e1Yda1giqtDsxesJJY2y871s
kvpXcdiVwHapESkcg3QhUhgZODokxwKbllBh3tsVupiPS4Y00C43N79s4syRP4HM
M7Ee5n+0Xe24k6TzO09ZE+b3i5NDtO5CnmrAYJS43dOlyz7aGmBPfociTz2uoTdI
0IINXgAa1WDuat99Rnc/UQBQAZP5Q9Pfg6KS42q2i1Q4i+Z08wQeOP8dNoZs/PTx
Vy6TdE6Hre7d3tsOtMlceOqcsLaahmRlCZCozni0onl9FuRbjr76e0jknN4e3U2m
yBGxcxKjgTJZiU3ZQG8Y36Zr3v8xnURTPtCcRiiVUYC6noGVb+y2i6IECJcLp/mD
bD3EwJudcg4eBIsAT7H8iVdknnixYJHENXokZXQJtSsw58Q5Wv6Q5lw6013dnZb7
BX3POdbA74KADPWsMpKWkVFbFbXwfYmeEJxKR35XsbYXE3pxfeL3XIxwLw0oJqi2
ekPV1CUR3z+6qitZPZyA82rbATBQb5E0CNB7rAzkQVuypoW8xT2CbwwuBNiun26t
sAwSIgGRNRES18l+LtiJgpCqKBJ6SsKmtwtLypgYZXiY9D9gRwwKMvJhtsH7EwWD
4Znuvb+QKFswF1EsA7W4/1b0BJnbo4xaHGwWOgsigeeaBBLOO/dXU5TCw1cYiQRC
KzS1024WEtgSgXeQYBtv547vFtI7koiz2FsnYYPowdLyhWMuIA5OdbTnVCXi3vUY
yjbdFASARzl8pklvBTuj+yVPLzrPkNVX1ZUrCseO72bQ3A02sFzzFHOWFSTmQ/N2
VoaIPhMhEw5S9H4+dTH99XIrttXNC5Xb2qBPQXBHZ4CVrqQuYeCWWrYAAToCwfZa
4RGin7ApqIE2BUETsWN0q/WzZm0vIOIgvRq+jMsHP3d4brEab0z6Ms0LHEDaZCNA
FhbJnHfXg/gSeoF6TpFxhrRY0Wr2tFrkDprsozQQxat8v9ojyoUGA8SRH64+tdGE
iIjlWvo2ZTe8DgVOComOqtMTpV5YyftQL1k0A2G8kM4rylsXI06l1nyQr29b0emq
yXCR4yq44e0/2BR1PN2H+uEDyCsmYe59NPvl3qSiEqpV6KWrJ8RPZNo0q3DWse3i
gNYUPH3SgBW/8ztcuNwnj9ENeHNmbqyleAT2YpLSL6+IuD8YDyM4pnec155QeYBf
lU0QeDhCxGKRtpE/uTquTMPtKuoZD91o3dPwo/m/b7wJp2NdK7Q+4XM+6nAxASav
FixS+rjUK9r3eUuXGsN/mN4AlxLWgnDro3kG8TGEByZqbMImyopiBMCo4YP0KtI0
dz43dwL4v8V4f65JYD/2GtO/ChQIinwzXgysIAM8SsMoz166q8R3e8cyC/HiRge2
LIgIKBaQ70Ehh1vNVSqK0b2av8HVLX8lq0crkdgazvQ4MW2WqXuO5UoAsNRsNcKl
/YWQ/ErbG613zkKexUSU4f9reY7r0l8yz6pR1gw+npGpnN0ybGcrWhGr3xwOHUuZ
we7MSlKLhRx170Q9w1t8kEKsbeVDUrFNgC9gDa6fymIAuJUsBLpfjaORVNTQAUlD
7kp009YvnnmCC9Hb1TzzrzteTMsAgvrvH69IVY9PKN5/ewKD+8oErALLKr4c7pQk
P3Xzwn0fS4a+0fsIDf0dEykxTAsk5CYPlNGuz5BRgHSTjjeNJOL4lrBYjsbRbcQi
J1cTSgRw6hfbHVgXOiOJgTNS4FT39QFVOQh7MlMIG1hwUVBH+VuskZ9PXb1sV5bA
uy8UlJnqbu16cdLN13XsVej1D8lU3U21lqd0MKDnwzCkUt4nE8An4J35Iw0QCARI
avmD1WedfxYCYgyjzGXQmhaGj6+BGuLif2yHTy5FGGE/Qzi1vKtHk6pjxKfCHT9U
TRpNjHeW2bNeHHvfhEabICwcf2SwzdgXsF2vjcMpB+cWNPrXj4PUGu/CU4P8dRru
pTplEKcjYO56+b+aGDbIND8ODqinF2lresh2g5zBSNkVvsNqIraHgl8O82loPacJ
YaTNBH9wVD4oRPbWSayYQ+P2TXdjJgu/worTt8FzeM+VarDmCp83BxYHL4npAeU3
UdLdbnjIw4e2R4KgIB/t6cKled8hrYgvED+Xt5mFCjsWCZcvvtgVE4sv1CG/e7N0
cbWNNVez6Q+czebavG89yPsMRi6uRu6rTXWvME88AArJqUKk3SP3FqMxF8kHOcve
zgIilmPGUBt2H9bkh680c+x8nebLb8NUKtczikW+jndaxN53oEiUY0JcgV79vJuu
aPd4QXw4Bn4ClpZNikjYlkpxf18LHp6mbdsQiOYTKZmqHJ5/1R/vC+griVe2YLC7
Fn+D45TB7sowSeXQemxzn+JJASVkHUb7ndAh7anA2CZ8QRUiPTEhPHVkyWElHVgJ
/oQSfx4CGMdn14o8J0NRTnh5hKlcl/Wil9nU+XYS06l8T4Rg2gV6+S33t1PoPf/v
mO3mdlG7VK9v1P/ZhKbn9BAJO9lKm6Ldy26nNJMZm/lkXSrTmeCfiVV4/NS3Z8wd
ORu7VfBeJ+S4nsH95dAlCYWE96nZRdQKZE6DbqTUHcON/TlSzhKM2/2nYcTJTAuk
an2gRJFNGFMAxQcV2k2tUHmtpM2BGykLtIARCN5c2KBP8XzxSX32t5mcUY5Q5trP
mBqA3lBHhXqFyUPSgRxuJygslAK++t1U7ZIdJ9P9DnGIS0hX02D4zlpqQ6RrXwDA
twSGyVvcjQSWGMpNKyuIzLPi67thMy1roSBBnSNP/nMG46p2qZQtcV5cxvN6fPK5
vhMYc4Dwj9CacIlYvFGQCAYv7HElTLa/z1rdkZfcM/R6r/w3sCD0jG3RT0cBFzlp
/nXey/OnY33qBbkMFONawbt+edOwOtP9KpXk+48Wp8b7EDG8POCm9030YHh7F0JL
XgS3iSY9hnh5pldw5F0FAWKcbBfUIK9pFJfPhoPoHO2NXuhI5+oHEHCdTsEKfPsk
P977WaoyJStUc7vmii4r/5JalrOoigDysuRZOWKka23zl5i7H8RQJ2ooEnLgHi9O
cLA1IVOht/wsuYxLdFsV3x9d32O/A27HwDVxouLsJKyOtpWh46XIAjIqhhuYyuyN
AzMwpe/tgxm5niigbeokJAgk0NU6wOVHEpMcWit4jbxFGlJBMT2wPfuNMOcdTBbL
okAz4qBGA19x7WeqqgOQlUqaG/8vXjlO7CCt2gk1rlkCsbsUoNJlUxShoQPHYcLI
P7gLaY6ux8rJfTrOSZeh3ChGwlw2fU8OXH0WWIrj1jpJwHR/77Vb/fGkj7tiNmbU
B0vdonShpPpjSaFmmr1euqQB/Y4trbohgdYe7QpMC8oOUmC0YucfGDTGqTYbqAhX
cAlgC176KB5uSYLN3Za7ZSQT61jJoYpivsbgDdNWW9KhbqUXXSMStLOyfFCQ6/Jg
GV5NFxHZzWtzQdqyyhCBmphnje/SKdCJrcS+IfMrEOcDpomm3UM2kdBlfSBLemLB
laQwt9YFpskd895x0FCAF+sE5Ab9jq3ZSjQrkrRXcpjZ7f5ZBWWSE6bad4+P5kjh
Du4X81wt06CPwQsGNeqygmFAQxKblCsWGGGjbZpX29MTU5H5T1MXuGXqOr04aH2h
OksCGiNQHD1ACmE9Z6rToU3EOJ8ckEoVOKr8msb0Cg7+kzJrIz0lYzYdYSEvD9wi
LDVLDZl/Ci6tin23/Oni6zCigYPL+Vvr6+1PAKhSqeGedj6bNouqi6u2/X4gvTcg
6O7Xle0C6n/1qhRCQT3hnmwz28s0gZjG9/pD2LEQiqZ4S3xt+913gBsuHftWG8fy
7yos14ofMY8OYJTVXuRorFp2//fSpYhiFLrBP6C8nnnagcmr27IbTwfHpyNKtRNy
eJmEEowwBQE5OpvQH/9XjL+Ojpaym6KSf+AJri7yKMq1yPG5pnWGt2mz44e2LKzz
byEg+Z65sAlvURAb70Ylpg2uYcT9mD9L3G57J+dD/Zzk/1cr0ZqXL7TYh5i83Ukb
GzoZwrh4+B5gwKJj8U6QDO+1HeJc5AbfedUVTK9n6BoTuinP/31nGQ2A6vwQQKRS
HNure7d4JTWO8DLw6PP16+vX2pyB3Uko9gH66uhukmaIfdIQ3cpPdLX2Pw+qoWZQ
b0/Tz7D3CdHuJSpJFDm2AUGaNqxZG+qbc6L3oceGxHx/hoHFmRiW9fNj/GP8Vv3y
JUy4J+F5Cec5ikI7JqOM9lbx9QNQ1NHk6yc3Re2Ej9Cyl+qhXS2MuEf1rtqVtuNW
iKYkCl3xZ9X1gF7yww0LLn2X8PuoG4Ci5lZqBFbjN21xTzmK/xwfUmQ3rs4vOtJg
r0cq4z3fMS8ZG/Rwd0R8SWAJOFlqOXaJDG3bxBTLDQqieZK/53sLUlO4rCN2gjcF
3h3ovqxJfwUfC1wdgCaylwRVlibsXaFBFF7NIJvXTl6Uw0QzFa8COVVf4wR54jQU
V6MKlnkFNxPpXV8XGXilfNttS1C4FS/+JHi1JfDwMNe6cN8t1nfRvnbU9m8qkpO9
onzfRtKOSCtNdGJx56P//aWT6wpMUtliyfpsn4G7Wu0x2th7MraB5TsMqYJXw+w5
S7xvwzR/9Ldmc18SlUAZCUbK2fKx0CvCObhH7/+wmImW4WzAwFtxJjE6RKHB8XbS
nSSzIMkhzNVDMWfXLQU/xcy/EpanSjYSx+vK6NTDjiKEYr/9LYFTYaD15uipjD4Z
r4rFjDyWnsq+T8qI7KJnR7liLaWzocAIbB/7u60gD4mdgSIN+q5+yC0Su2CfOs2K
kh1S/1yLMT7d5nz6IAkRQds50Lu/hLe0mjUKg2Wju2Gbdxb7zh8AeY6CqIv2951P
koE021FbxB1cTZDCWGmxkRBlfUptHBhveKrQbnWp9HmYMfPhtqxW95fMnVvcuqFX
NTOPFEqPvyDgphF0rq31U9KaPn8x0g1L/IFYDx5EuOYLLF7+J3D1PkYv/IOHHlws
jvTdFpRi1zXbUxO2ovg70BoHCxb5QWG2M3h/xCCY3mn25C0dpNS1LpC7cFvbgUfd
2bSqP6uU0sJ+8xGEruu6S2AVGx8v2dd8ye1Yd4AgBixspSciGIzSCej8EJLBvlGP
XMxUtmeUnSZxN0o0eDGKtGFkdLboLPFiwXwPy234w5buR0kCHwe5dNzCT2lkww6F
KLMCb0i/uaC5LDav3Mdeln1JpSz5/uMsR5oeT6rHlSb51psIBxLWRKnQjxLIlE/8
2gTo6BGz/n54reVV88CVSmnP8w4Jdl4w5Qof7rlS1tUEW+roCmpa6+7HgKVHVQJW
y2aSkErypM1FQ99EQIW23BlwUb4yZopgznFJbdNWyLPE/j6Pizikss+ZWbsWtN/J
/PwulWMLe9W8Dw0+zsblF68ADjq+yZI905AX2YQlSWtbn7PdPn5YLBAvkkqvOQcY
84TnACM42VBvZl7u2U72PZt1i+ooXDpn/JLdn6fq9j0OVAtxyZ4GFc6BtQ2AXj4O
81FzPVWsom84hk2BDfRSL6unEtKGCfAaU4HzXGUzSJheqdL7UCLV9iaEVyz+4rZo
Nd4qoKvkhbs2JQGGfFjfKur95aeUDcgsi20KRh1/nmPDu7PjEo9ulzm6TcHkPsQG
J0lvrlSYsOEGz5r8S3a1cMu8hXBUI5LwBCt+v7Dj6+8rpb0gXOo7oifU3olwKb+6
g9czGjxmNIoi+jr9rMlW5WlKXApBAxkjvwBQnRHBECO2M1leR2yRsPknKx855ZcO
glvKxZ0fr31QIx+//9Ts1E4sNoYpUsKjSeLThWEbEkfgUFNyIply1oTz3aOjcn69
70diRb1bT2zZVIbeJ++sYQcGMN8bciiOxkbJ/HT0n2HS1MHM0ctcyadXyhO8ULFR
MphRMbkPwOoTDpx8kb42kpeNwNzI4aKRwAH1jJke7/37ugavS7NH8Hw4Jg/bxVvG
opEAf5v/JNA11+nn4IWU7B8G2wyivogBij/Ezmq+6VIRRmd7+kf+wAKMs/YNmK7M
ge0N5nVkmCqV4bISfie4MVY0AL3rwJlR4NqH6nfKPxDS57Dsx8Ghc9wynQf0il+/
pu5hZ3m6N8CKf81U20CGAtg0jKIfvA+5YVopxncsi6YhcOvyRk4mN/hjTj+70dUn
mNi/2QfMn9m38TP5ci5ms9OHu+jFg19d4yUo+4NtmnSwqtNplmzBTgvYfJiF49N8
JHKegtrEfpESVHZnQgJLBjkPK+uudwX9ohWpdO/5SZJDhxbjMTXKxqy+A275wtdB
MCVSbswTYZGtaQywYaMsguCX3LgH0Hgqv4J+Per7WRmTUTmWYX1X0VcJUfb8d/Y1
ULJmcDWe2I8br4UPXLeXaWX9CgO6cj+fBo9fQ1apOzZYIK/JoUxKIxS8HqqHszgu
BQr0rjCUEZaHyURNu5TBgZX91ZHUa3X0mqqvEASx8UJHl4QNbgrLW7WwnZxXtSHp
r0PL24lI//4ZiXJp5qQSQ2GjdoZm4vIrqLXAva76oH6hq1eFChKcz9SqXwC6+906
v2bKVxsEpQqf2OgGwjc/JP4c599lpZ5g1bo6T2k28w5Bq6kOcLdHbYg/v3R03LpX
PibR4RaQdFa07siPgfDPiw8RtHzq7hAfDqDv/HYM/Hh6D5BQJnOpe7aYm10E6lrb
Hr9vfqykSU5T3flA4V+uEOB/P8+pgDddmGsMMkhe9t6nCINVAkNL/qusvAkyY2iS
Q/pgdGujkjRmC25qKe582pyd3j0Z5GDPkLQ02TnRJWlwBiXgv68C7UNh62muK4Sr
rTiSoR/WND6F0ObynsXzi2SeICJ46kHBEU1LVl/PkFmyuaX6sxaosN5fyOjOCyN/
YN2QSeMJC5e/mCM3PhHyneAVxMyx1Tq4leGprKAUSiVGNge6Pzb1Zu7iNxzDRkrD
N5riYXFMDoODMNTAOR/AjEKg//u5OyRrobc7144pAi/H9hn4LYujRinZA4+XGDXD
VFY2fxS6Uw8HQ6oFnLrgRNRHElXRZ6Qtoble2GrpJ3XT3xdK0Do9n45svLK9xWo/
Ck0R7pjMiI6fXhVmghWCfi+gcmSdU6avFB2KYRpDWinlvkcCii6/oV4O1dPboKJW
077z2XMV89f7bS9uJaXM/sbdTAeCB1VAQBlRhWcugCV1iXTunYjOFklXTw4lCKom
Oz46RnkJjptkvOBBEo9Mvagvf5S2NmgEpLPtXm79kp5RsPXEB1GefEefiB4h1qkX
p0104wlIz24FvNuDEDri4og+F8A04HMf4P9xD390jv9aXHlTjsVO6eNoTrjCQJFj
izGz7hkH/XDYicQKEw2kT+4rRYDCS6hPyJgyMt8ziqm8g9aBG9MvvIoC9DJLzvtW
vZJX6uKd9My4zr41ndqgIsOEW5a1TtY4Z7eZ5u3ksg1aMqrouPh5c8dL2VHHYrOC
pkRQ80iKM9CfW7IqModTkqADJlnAi/9va3fcni8E72W+ahbq5Me/T//1QjkUamjo
giX68DBHOGmCrJb9tCAuC8vFTUAheJKA37KI9aJha1En1eN28sSPB9V+v+8kgZ4A
GfElWIX78SlcPXcIl54dv+ux5vJb6I6EtMjhUrNpE6xlvZ1zf13ymk2ZOul7VAf+
+/SwJa1L/WtWFznf1tzHhIRieiE1Ak+AOP074z7/F+H7f/JJL4/ZLqXgsORdKk4H
n1J9tWkjFCUcnVXuOfO1zSbWR9ZF9xP6+qGwG+G+4b0frREARcEkNfseVMwoObF8
VYzZ6qtsWCDAlcZtl1mDs2ZzodX5vj/1sRSIlUsl7CEyg4idMFc8M667hnXQpzOb
pQa90ScUBQatx8u8v5p4yNnjelXcpzyZgwGP6K1vUD/BCWS/F1Qwt4MvXwb2jJaL
TFBGFnk5WjZkO8db7gX+1gNoQano8chUuZCAuVw9Dd6yLCSptxF2atJqiuAxDAKj
SB+oYiB6bOieTOWq3qKhqoLoMXlfWi6lw66UmcXNN+5I+sewgXpyqF/PQICPY3Am
BXYiitQgGtna63w9w78yFNiq6NkyB4dmnm/e2avqnYuD4c9cgiIoBa3sgSJYgzMe
UCEOmEdy1w7Y61MeMtwpvlC4V5swwVrcuqJ/z5W3lBMJoEyqxl+dvrxZwwPDVTa8
BA7UObDJX1QD5JWfAcjzM84+W2jfWvYW0yILdLMb23vF9eKZSFGYTV+w1jwzBA+g
EHEbEssqTyXZuEXU9J/1ceBra83GpdFqb3dCt79bar2oVYH1dvWOVo6kx+AVruth
p3UwtNuAqUB+fdmnxpZ/RJJPJWYTfsvP3CobVqnkuAe8Ty68c+Ib2vXQe9W4+y8a
MwQUO4RnzZwbvsesGzgIhSBetWFfH24a81uPz7oK6qBpoyew1eDPhHPQ8pCqfys8
q0pnaRrEgeoGC7qXeOs407EDk/MdfrcLcNEDMusQhMb6hkZuqKY+JLdgyzxdfKyZ
lKOT8t8CEtQQh2JIJdY0suj/xhMhmYprasDv89FPt/Gngudr2O7D8aHcXNAm6hlm
v1eH/rnlDczSRhP/rvtDfylT1FPeBlEuVk3s/eE/HGIt1GqnrgUU/c4rVhmeJcXm
6rysbrmyMPT9H6/eq5h0C0qfMsFhxJxQZW/Q3KNRNbJN1Ap0KtJOHLmeTSrtzhHk
xSvHecaYPInz38+tyVPXcZGfagSKbLLqnQDk+3Ub4/FfLYmArmQm1Crjlmg8OERI
cE3RIR3vvPML4lwVqO3cQ3AOT3tqQFu8Qkbr0FIcBY0t4vU1faNnNXM2k3j68xWJ
Z0duyOymmRFEzhKi/lsnQUpSDWlhzjbsSDOnbSNAGeeGfBU6qH3dqsAZRCSNu4U9
gYGb/Ui5GnAlm1mCT0xXqPolh01EgK6UwB4CvI/L7vJxa3Lxy2lo/D/3ron/ln58
1hEhp1QXd3cY0/tEfI7+azQaVYuihpTGlCE4FayFDgvNoB6J9IZ9AjN87nSYH1aR
bOSpz7LpWnEnNFQALTxpofJxR7aHnM+Z3wpNaD6xjQlXwz4YD5w/WKpO9rvDAQy5
mUpAdJmEFeupcbwE41B3vhkWAhef3okC3uvpdRRcPntiLLEdzJ34J0Vgv80rOKOR
7h234K5na235x2R6KtWsVM0Svcl1hgDMQODDle7f47UeD3s2mRGZR4MI5gHl7yYW
GLkQUGVO2Q5q2Hvy6t2N6/eW4ruJPFS4QDywNM9/vb8PYLTQWTGW9t9l3/RChTfd
sc4Tc+WsnXHueoOXFO+Pw/8md0CKWlCBOslBjIEK7xgMjo30nNthqeYVbTu2brHG
zJKw9t+fZILIyRE544tkZnafxXsOYVl5lGdpqwYNJI+0RysqeWXQwHCBoM2BTUux
/Q+TbrpyEOnWY5dVBVWLqsTYSedy+jkkRTW2CFwFFmC+S50Th7A72tLTUIs/XmR4
c7sBMKyWsfDv5H28BZifPPDJHHpsUAORDR8hkrSmq9iTJGnVBTJ1BLepgov54qWo
mEqTtMK1lzYER7gJAV0oy3VLZKdbzJ0baTOjkf24q4wbodb8jKHudxzfZpK50AuC
yOpQV5HuxTczm8JqmA6XnwAg/yqAG2brYtAJCnVClf/QFloS//R7Ay/KcfkkEac3
2RTTIpQRxBvnLQrqTBaUbN+4XtMSStj3VZ0kqwDBxN28fF34KBcJEsDEakv7w0ie
t0VjSrQyL+T2TcylCulnlAHf9jyn8OqobY7s0o2Ktoej1I2BxkBSksjfMy1SNile
Eom7jST5w5KHByAFAFMIghZmWvvs3xze2saTEtDLK0pdeJ3K5Zi2kiE14rMS4SxL
rwzRf1N5by2x0nuqxx1xMLaG7/KiEeWC+HmA2D65jDT8qzbOrdJ86SFtIZ6xzP5+
sHBDnvSeR9vs/GZVOfeb3nAHXXF+fx9P3TekIai5GFMUAapY+3+t5KWnRietiwa+
PJNMuBXP6MwjbP4N3PNg8XCY256EIHXlcGGzK6CN9H/Odi5+yGk/WFEs6szNz9S8
FWY8WjWpyLnDz/y9N8hQN+XXcYr+xU5UOWZ4cD8gkjlPyOFtDXRz3vhbbbDuqu5x
+y5gqnVLeKrBhkeQ9Lb+kzRO+FYRKk/jhJC2pn29/6icmZqJSv91zim/vLM46bJQ
L5ur0CriKHllgZ49kPfCFh93Rvj9NkR3fzUOf1R/HnujUcoGwJ8PnglFsbJKAEUX
gabwsnMMa6e4kcIIdDY8VU+cy3iGsusfE6utt7UnAdfd6CSA0oEiRwbDdd2pnpW/
8My7PgURus3DJTgeOphnfc5ozFsTm43+pXMIy6pHm5FnM5VTL93hxRwTZHSd2NBa
q6oPZHLxzVJIgkoP6LvZs9INdscn64bl2i784njhS9Z4JPOdmDZjSH1/IibvW6v2
e76UtcfSUZDQ7lLko+FkvglMr3Xn/XaREOx5usNVlsy+CeXul4QCpzdJ6faz5XV+
g5g0qt0939lMZg6rcggvaPU6+OslN3/ZViDoD3kvB45cvmwSVKFbpWqwQw+7MaVz
2niYKpKAKS2997a/JmA6HguGyTbK+PyrABjAeL/cdQFs37zzl/FIRNxsiBl9MwU9
KMUw0508kdjO6J/7Mbjq9QP+wE9Vh8F71b0CpximEkv+KJfHDeE0hd6ErNzHdLPG
XrFIUXSoLxgu3mm7HiqOW1ZjQr9DB5S0CRggLR6iZWNkzX5xGjLtiUvYsY68jdOb
1JXFzKZIViNJ6WoioWhDrPHHvlKYU8quxvaIXrIuJfGV87iogdOja3y6zk+MZLOa
ieEx3N2g8XRw+NfCQCbyk0G2SfpInrsa3hYtfYGrrKDkM0lAsIrT3h+PB8y4d4Rp
vYEepnppVc3yRPpWibkVuvV4SZ+VjimXCMuIXdYPrwv6lAnTV8SKLMh4FiXJe2rn
QYekTjLQSpw8m8OiG/nsh18ABdltriPLuljH9N8dk5x1JHbiXe1SsFiZOzDhVOko
0v+12Gj2x1L6GuyRrBZropC78ddr9KrEe4C7n4J4L2qyB0dj+5764Bv8Cq65fY2Q
kUE0GUJSuqtNYrWGVdUHk3mi9PrzTd8Z/Cq/ovZstkuj5Woz+fJbXbdp2NAzQywo
0wAFnsg0emTv8++w+JLLKDYHb9Q2jf8T/NCHwTFHlD6o2J3q+C+ZWLUKdBaoMALW
N8/iwa6KC/kDwCGOB+gGwdQBj1DbEz72obJx3u2vu+uTkaUOCbDVcwy6ijtnrn6u
3YuZVvW1j/tO3oud6Nf/IQOpoY6LUYHJ4++bNPxjDTeaTNFRjdQ+GwWt5HMkw7sT
NAupMK7srlyyYBAVWNoNnCj5wGh2+D8oKDuTPcDf+kJuPU4Ulk9kH/ncupRXBK5W
BIQpD7vxp1zrd0iGAEANy/NkBhvsgVJsiPymsLW5wdZIAY+GTRSG5FhSegkZyf4H
rzGIhWZcqCDFDkODtc/w4giZMNVGJpFRHoJ0ygrn6yZc/I81j5qAl+VDbuRWa3QM
TSX5f9mTyRQbm8UOhy8+Xes7zR2hvcCUa9eis60bYRxbMwI8O83qHviNP3Lw9Ssn
/l65uCsSqMC3vq45BWo6tht7iGlrqEqbatBSJDYtUyM+ngBvOZxrkISDbs4xA1Kx
7HRZ38UtcBEZUnvtQMJhjjVqCBhPajW7v9MDHBP+LdPsxQYupxZnNKHIzqJcd2De
G0bcYEWw2beKTB/f/imB0Wb8mAAvuU8ehuZxAE1O/+P1R4EAo0N7uRorF/QlDzcO
r/YFJ0+DpGCtoIKt6533avpguzZtbi754CXTTXGHjWRmLwXrrlUhIrJX7V4mil5r
wigU0pls7mT2zQbhW0KrBt9ozm37/TXRNYtrzobj3/1BOwyrynIqxCvWPB2HhZX8
T1WB8zkh9AkuCVqXwway/54CoyFmM741EooWwhw02Pm9+a+78Dp4TN1J/skKUsBm
7yP8SmiEL5OIvFbzU7/ztodMSDXHb8+HMgSf7M24ab1dr66JpcDm99upPR8nSain
ExUOlMQq5wrprX/9qq3Irg07yCyFlAsO89/a56Pz0Qd1LM5OSp+rTVzqb1wRjeYd
KB3/iHM3ru4zgD2enn8UuErPn7uWQ35M8qzrJahFW3HRTpwqfN8Loyt3+0RJFgdd
CjFwOiq7JuiPlNenkL7oGr03JbTFEAMs2kHbTx+JAeBxrUs5wwWVLz0KYEB5RjC5
zwxkAas+UPCF2x4mAF5embqlQk6HFQGm51roCDaWRhY8daEPhjjEjybKJxpZSu0h
7kZkBXWL/O1OeyhNPXI/GeoiCQIw6snzlW1IPLq533MI4ZHFEo0A1S8PVbk5+jSP
tSb11mTRBG8REGcFUaX9YE2dx264KmLO9XvxlC7a8CnXBaICOJo8kkfN45WFNQF/
keZGnrMagyrdKq63KmmxYRCyrUCVa70t4/h1uA9eiQ5oHe5xySZYlZ6YkhxU5GFx
PcLKLlkytWHJRvp8ID//cuxtBmFxIR8KID9T06DPIcKOxk3Iz6GZ9KTq5yXc8rCz
MIgIdGqeqCCfuwFj9bKgQFMweNcLUGsW+yac31CmKwNN9DtB8DUh5e748w0VialT
5LhBPjwkiEMf7iZM46BLrTevF1I6NrR7V5hmE2IhNtYr5VuvxhltpxoBhlj0W2b/
Dkaj1Pk/choTGm7/AuSM3Xwp/MVjqJkdJ/JqfythIHHpAsLTe+8CpTBGN1JxLkXm
2viy0OEroPzfNAuZ8iqMMRfkv7psHHOx0JUk4tYCW0x9+xcMu6b5vvIR8qTGX70W
ub6gwlY4JIHhFjB5RwaIdgWE8HuyounQncE5pHH2Jtt7aNi0EMz/raaxWuiCkHDE
tXrcRQP2ymH9xEkFm6wY9gTmdQRkAkUfV87MiyzmSrptfS4GtZLu85TC+GivmXzL
ZTViKtddeaWjOyeZxkOa38N50N/rwkhCvi031JPHOueYvNI7cz9gAL426gp3KdhR
EJsVSK6Aijm2NcpKswJbYs/QCEW6iH+utJbPgfAgxb2VTXa91Ern2XIqN71fGUv+
qAdIE/DDcIV6KInDzmUZ8XzNR3bW7w2VKns6IcwyKRob5fFd+4oEgSQAySh51MbY
Pq6Cl6zs4uExnNp1KUUYwxR+LvTjzxXHheWER/LCwb0kRF0Eb4KlzMfGpkniO6Ol
jKKwXUPVGwlfSXqKUXTnDc8RLnMVcK5Jy0EQDUvekzZeR0+6IVVoL4e1VCenV/Yn
Z5rdqgB+BbsJyMPqpU9AlNgpjADFgu6/zW72BYO4V7czoRc6diCpQRSryuUBYc5g
mL39hmE4w9x8BIbWyt+EIWfvl3uUB5XzZxePsDtaOlO2MK/YzP+si7YvEMbxsnTq
yNmmwXX6P3yaqjNjH/ZZ0O5r2IFp/BMrE0XUy7Ok2WiiBS+sTXPIpde95+XkIv1J
RMFKx4iztip9wfvGt3y2obfkhIn1hq4WusKBl+wxkCxaRyktSvZcOynLlRCotUz4
QY8SWUOGldigXkOfa5nq5ynP3K+1hcLSi7eqZapVxWyuv4KGUbyvr5MVJ7FwdpfR
BcEzRddJRfWrs3+c38ecfiEsCjiQRnLRTz1zRV88f1qTB0pD59pioLYx/xAnAex1
MzNuksmYTg4mSSQ9GCBDu4dXeh5+eAcL7YheQhWv2GgE98yDbqCL67infW6LL3KP
TIZg2YoCAK4M3HfqmbzDDnIWhAZWkxLdN7PGIfh2YSVdWKt7FeQGmqd0sdDDE8Z7
5VFIMNm60O1eCbnQRKkcbpPBRzC55gbbk9RuSe96HuHpvWjx19JvBUgaL4LBR8ZY
ieI+ORH7eL9jWWbyLtd812yO/3CvVpykoSXSlLIjv8RnzK8YVK50/wis8+/AeWFU
6//HXdu7YsIhCkY/lOZC23C7K4e+F9+k+Cn6pPIUYJYT22NWolYLdxfGkjJxbPnC
xoK7v3DINB5iofD3lSWv2Z3MUqJZIGCJQ3SDqFG+nTzAvPLn01dX0UikC0Y2QPAH
0PHHrFDMpNBo9xiSX52oU3P8Ole03Hz7DwCkxR4Mx7Q/1v3wIe7L02BnHbk+sBf5
bEpS/szRzUTEqdunzJid6PozUuNdsqoK88/LBbXEWdqXmiOqwS3K9qgdjcWGZkV2
qP/wUGWluLQFy8UxsOosyB2tHbRc07yD25wMSEozGrigP2REqSZPOLJjt0X2t9WC
jAlMEvm8nIG0vbqSfXHsn7hyHgKocOkhUkPggRNADG3/woACouFXMN/tTK9F+Ba/
AZm8JPz2w0w5KpPizE6Qgs7E0Flkcfgc2YQBMsyFvVyYvTggVkTIxw/ZKdD7Dgr8
9KpVMr1Te21bk+KZAx09NmGkL7MqM/CZ45UkG01XkPiaO4azXKGOgelM5LCzpqpz
LFtt2FRDMz5k6RuxneJnkuGezsOCb/u2DKsYc6yILKFBrjztUFP0hOt7mY6+El6S
eIGCNE5qLVLXZWQJSQCV628B8eDps2vY/6/n5cqAgc2BJLFlnIFOPEJqX9s6JN0P
yawQPZNDuN/8DpTvdbPwoOIRX1etiW0rbeyIazVEEqUZiadS2b9bD+jCLbyOtrRw
o2iF+HIgJ7kmT90Fm+ySyG8w1U7ta8JrkHSKgLtaGVUzWmepn4Z3VQazPZE5McT2
PkbxhmyZoyNHbiQM13588bGpR/nh93z6sTUqqxfLGgM8x+6D6YqcLdjmX87p7G0V
xMC4uIfCEihlaDqwR0VvSATBrSUVtXsn5vBxJJ8st4/FoBHYmxknVJGjsIC/+wz2
AHtd2i0X6yUJH3OQkq56n2h4VDmsaIo44NjvH05uBjRfIEvoDg/TdK0cBv8vx5CH
JcqkUqXIipYRzTiQEu5kHqqeLlw+OkNjnxH0EE/eABHmw1jf+Ie+rLsfJ/IWwGgH
TfXwE2IGlyomtf45cdfr+9OVBVussP45PmB5GYHIXPqWsEIJr1QwQPNhnu3IqUnf
8oA1H/VC0v7rvn2YVfrvQxpvODxifwoJj+axFn3OKMKSMG7oWo91tkzcUdzyJ2oj
PWRbAxJMS+JO9krUTSoVea/sl2/P/CBWVkKRikroKlrx9WqSSQZOTetrYsAXkb7P
cPk44ILWknV+PQLOMhe0SXI0hLU83a2CKKpJ9suUHW7TPI4mCLLpt/MF4eLCkvNE
zR31+jFISVBQup4yiPqqEqnXgRPmfThHIO1b7HYaA7eHwS3yB/Rmzbg6FLRN3j87
OWHdRcUUWYfxnPK0S0vTkHX34eMUc/hdfA1sBgkguexdMS6yg54+VEUYSOz4wZ9+
+bNrFU1p0cDD4SvUV/W24Fbq26EWTXxUZ5/SxrQGT0n9jTaWhJh9ujL1sawqXKle
eFUhfm3Pxlqppw1TmCucxMtaaDk4bUPvk+88jStxd6MbcHmt3h7fuWfnTyl/CNqM
1ski7b1I81ulh25c/+3n3Qmvjyy1eNkSXJ2qgWdskoRGvxOLQm5ZVhcWmyD6kzgF
q9t/rO0O/SylCHbKraD08SK4bUq8r8Qw4Pw7c/1RspZLOZ1EVB2tWKbUF5pNJBMS
qQlzhbO/yQfseTAPsFsCd/x1WBcDI5lCp/KrgKiRQTuB2o9RwWjcYXV6NyDYlUyO
Rqs3mf1ExLqhGnwBCIuhEPj5yd/Br01ytHBIbE/xge9fDLBrVROhlvC/UeCXBIxw
6ZeQlpelSnzgBZZLUKHd938O9BWWTfCcz0kegXTkqy84WJ9tb2YCCZRojp5TMB5d
kkDG/SZd7/517UUQcEtzRHxvQABphC7iyxTkTE7WQ647tm5XCNGga3dDoGvIu9Yx
9qfsi+CapOrarmfGZ9zzh+q/jJjNichqLtAtaTlYNMsonlGI8E0NdLmcPFbpgEEd
dcQAaTsDlgIBGcows77Zb45MES55ZmQHRrlvi7a3e38az0o9Y3gZBR32Ds+IXWp3
lRrh4jDRxFz8TmCTzFRM8Y0gySRUO2aAwCcJmLUD2CARlfBooV/MzACcowZALa+x
eBuDxhRU2GR5a+pPNYYXlmHgoa/dfIo3sG3gfc3yguk5j2qitMPM5odWUjuqfnUj
IR2ChUpKU64JG01p9GuC6qbMXgLXPxg5nAsuKEo7WEmMs7V48zcFGxBYSx+6DLy3
uTjpbwV9i++tNQVYTJTIIoPOlG2hw00K9q8vemW4LlvHWNeV+mPL7KSaiAduARam
TsMCSlOye43NUhRSfyvfc0CK+tYLGGKHSKsJnqZIU+QHujNKFhf81ZnSpEfP+/I4
2uDcKlxd1eF2kQ22qyt5aaAKJq2DhKNVziYgzf8XSc5MNHhTD+9d9iE672OogPGM
NFX7RmmYvMomCAbU1DnBjBBMndZJqEHglJ1Cg8yJDZjq0+yuruIvk93YwVsox/zP
iTPKUPi0UAd9C1dheZ2Nu/w/ir+7q7LDI0g9GvuVy6zYA9ad7Rx9IJC3W+3W6SxJ
WRnEOen7CWX4P52LvxGPrugDm4Xzu/eSU3PLkPybkjyiwde2DNwG3EPww4MyZQ+n
QzOwAuWlQJYtT7QhcgrETrLERr1AOc7lJMgNIk4jiNbdCZrzLGIGNctVKW3RC6uW
NyzZlPCYuDq9rtZEajvfXtg7rnOHHdFFcgOT+fzdJIoiE0gpyIVdtaTpAVkwvBFZ
O0SvwYKcb8JFvaQ/z6bV/Y9NzPp1THMIpCVcP6AgDT+DOMC8A5xEsxPVb3hEO2In
/akQyn3GNQX5N8oSOl9ZCOKZawVJ8a+O9BrqIL4bpQyF7AXkQN2zgp2MfVQRxhAJ
KZGS8myf18liyD2aMr+fcJmK6JqSXBtN77EbvodabOPgy7O4/1mGLHZ6lAHc8uGF
1DPMaXDyHwJ/uFWqqF1MD8bH5WKdh8XsRFpgwIXgZ/R84hM8oqx+qXzDcYoz+afP
2oGmhFb26h12EWY3cq7WQ1hRxcxkIviJEoZMD/y2Luj5Wa6YVkf+v4Q6hYU3ZB9S
0tz7/TKZW6Djb2wNnoryO/7RXw3Iu01+XSJ2DWHprILDA6S7MNIZ7OqJL1WGnM9y
ZM0L/FKMW0l1WI0KynPBEFO/ZFW90eCh3GfgJyLkusFRIX63B8BCqXLC0ARHmcGz
rJeFtoA0gWiINmAVX1YrGkwLiPtochl6wqiC6UWBcKojaFLvKwWtjNrpCLZ/ZsYd
CuSBteLOOWECGrTdSjWVpUHpQafRQ9gnzOtdqMnd4nub2fEMMmeuiwUbra/m33Mp
KloCLiMRDPycBUag18W/MbwYt/tMMgHC03DwBvqgPcXg0+gsfGgT7xkv7kPDFVWR
wMT55mhIRgogvApRfuQO9rOXIg4a+eNaAXgGXfZ5SK9kXoJcEc0bVpVRrkb1AoVt
JKBtiPU/J7dyugO3p/Pl650ZE3FAm2UIb9/TcoD5R/qO5RnJfAqi/DCFbb64Eaau
XyfvAyTU7Aku+AlUdoZQCfs0NVkqELepm34e5IALOSP65rDm8S2CsE6gc82hkXh4
h9a0dtQ0CYwz7dgUcIjCa8LbuQ7giwTRjJEEDnNloADlqg9oqmcpvWVwYQxkHOWn
zrI9kIegK4R3SrRuPoma2kspiVL3V13XR0GFrssYotd0BfD5JE0VpuPz1r5T7J0Z
Bj1Ucn+stakGf+bU1cJWvCWDlQXoyYeuER1DL3BavX9GkYymNG3QF7cOIFmEqjWF
GaWpo7Mtjx6IpaqD6KtfVevZT+L5AjFEXxORSnx+MHk4PzRLxat2t9YvHc41QI5i
Zgpf0Fh9ZeBTpk8qVIYcx83FARlsDum218PAhmgnbNhalC5OoHxEurfKZm1uNkrd
Y9rLZTGD5W7/NSgpOCA6I0aCLIfqJNypRZ9ro1CyD+i+x9aUACTgnnhLnFlXd6rL
mbJ+B76pxiF/VTMIA3SrqOm7ZFY70mR2SwNSri+3uuAmUVKNK/+MRn1CseJ/xiY4
h+V8oMohNo17WiZfw8p26i5Y07ZnCnBO3o/jMo/HOpsudGcxPzJg0wA8XAYDAtGJ
IQA+MKoQCzn4Z/iZ1WFmbqnS0tR4k4I4IKZVZfmNMryCr4MI9E9t/w62oKnhikv0
k3GUVSI4sXO8/S8qU4ILkb6XjjhbvVJ2MDLb8ioQrxuAyBGgYLhV3f039GoVPi11
pbgaPxiS0KE2jvAKy29wNZY3JTmuBpxyNNnZmyEDjOJrEymb6xd4Tvun3vvhAkCg
5qNA8UYnNBqM+PAKxvdEQ1GF/8YSq+mcb/Jdw39QxA/dznMGgcJMBIPfQm7fxZYB
xI3pqsW/vrkhpWdI2nJWg0WcT+DEp0YpztYdxinPYfI1j8MjCxIOl/lydIIqKzaF
YXS43MDqMaFlMxp9v6GByZNbgWDUMjB7TSvwiYaYBIg452nrYYwgyXbEK5yGjNLF
Y9fJANKUtsa/7BO+eZQ3guvr5QxAn2EcU478TnN+5WKHKPYKeGmi2j0DvC/JX+51
0Fz3/P9aocfFZ04EMHgPj4hG7V79ATuD8DG5YY9San35lw69eSDnwIt9KYEh8NyD
RUzPoNhN1USd0e+q9hyx5LMGj0RapNJfceD4QFEkSSuzFOaW6F8TGgAJGF2i0BHS
zmvNsoJ5TauOtofcpe2yDMWymkagzYZJk6U++tUqWatgN/4RZ1PAMekbaQDKZAu3
oOdUnnbFCuRe3r1lzTclWDNZf33clUY77F5FKHuuMI4251wBtM89AawngaZ9KRXE
6E2bfxh7v4aH8bGKrlUOLwPwCP1jBPgbKV1w+BPgjO7H2WLWDs9Dnk+iaG+yQNEw
nXAx/jw0ZDe9J07Yd0032d8+NbwiA1RYsKgYIt81dWH313pxWL8B96gBQyxk9RVJ
5U+6GTx30oKNw8eIKTYhso73jgzyP2oUw3hTt/d/k1JNk8qEnlfKnTBXPaKoOpmb
lKgVzfPhgtgVtfy0hxugX16iFr1ZyBq6Ama33XBxw26AmQQSN4M0LK4Lxc8YB9aV
4yBZmK17xKkmBtlxtsMx40YHqOj+sFgE5dfIWfc7rJTZSPjR6BE5+FTXWox6QgMu
qOeuE6RqufsGYPqolXuzAQ2/3tyyIXcvL+6UB8kMfjB0DZw0R1Bz3azUcHa0xD9k
oWcnnrB73rlKBdvfpmp/JpopSmG1KuhbLIHlA8yL2Fy5Fkdczpz6CyDqgt92/T07
w0oMzGcnO+0Mzoi4IthcadpqYtQVVoZwVBbXh9nVcdiM6X0R/utXlJcmbUg/Lo35
L490Xa2DdOBCtDjF9oBTrHUOX+mfNV/FyQfRkG3GXSaAeG6/KEa1nzQCAc7mLgdy
/6w8MR5S2q5CI+8oIV/fYVpJefDgPo6/gmc8M4zne+x2+TQmSfsID7g8EWAFrC9V
9sTcI2ISmuMiCtPlr3rcILkEJM7S4ZkLCs7zz0jpx8zMTZ8nc7374Fvs3ClH8SXx
BgTtvcHcBrBSWz7F9t6MUmZlBULzhXZulpmX5PMt9MIU26OYDCwBNtjwr3WYO6Dh
cf5lfCYzPJCZxmGyueH7TNFsyqy+kcfMfaFLL5sa+eP87kkUgX/VbS5iKZ2uYLZZ
eeRoNpyw/uW8udtw7tarMR5wDnDFhnsk0ZXQVVx/7P82dqcGN+9K8le0wMA509UK
f05uxznlGwTuEbVqp/yjbyN3bLhsZYVK3Fq3i+9etyyk6Tr0ugOwTIh8EapN9M5K
lp4GHS3MhZqnz2N5Sc3wD89LfW6Asu+pAc2ruaVdtbHXI5Qj7fZtcSqWVkRu6OMU
BdtfjnI0SvjTTbP6YJFCuUXX8POF5w6xqSJN8vkYPjsJQdYUVHpK85JeWesISdmW
NK2lHUDcCLKTfxsiP/NIgpt9v3XbghTztyWTsyTjsY2K/9DnmSXty+1GwpZ4nCUy
4f0c34JpYWFb05Hg/AVOnK4+jaWWZlR6P2x2yTw0VUYlgL/DmNFOmSJtZNXBFf5d
dMqM2yS2fn64n99x2gSbi/fQefL/J2eIiuJbkeImQX/fz58gm+ot9BikySShph0L
Po0DnjY5/a2h/aZ4mr3K6WXO9W3BjasYjkuw7chbhTF/cx9A6cPgjDFUjssv8/Kq
sL4dNKMFeVPQ4f0hR6LU9cRTLKsSxQOFrHkHXLxtXWyHpm0JwUu6lYdzU35V19dE
IZdy/aRsqiqn98e1ZgzqtF+C7BLbu+YZEVxe8cGb7KE3AaB3iA0TgDnwuggrDe1t
s2w9WaJTPy+jMlxxFp/kotcHTS/eMMV4KlCMSklSlTcCOVY4gVCr1zthFkVivWUc
MkXu6/jZvDJHo56OXQhv9CzPvaRBcOh7ZA8/uueRmrBlsZV7K6WBfUSMSe+Zsu3S
hQnlRIqMRugNqexsdL6SUL7o1QE9811Ev4CSrUswvGCEWAPefFOy5md4Ig9JkwuV
lhkDYLlCYBQNLP9Oz7XqM23LxK1O6Zp3otsNddBossgCQa1aGtNosuhkrZf+uMrB
C31r3gmzzCnYr2Nv/ZuNMGhRgOYKsfl30vBHx/U8Z4D48anjM5EVOBDwfCO9N79A
RgfIbt1UMGpzwHurlxlp8tTidZAm6UXZO9+EkBhNT7bcLhsbgRCswizCb3/6u/9F
9jpKJkf5Xkt2tZkV709CfZxXI/Y1QL4BuFr8ZQUsqhkSIBfBbRFKlRIkZhubu3vB
WJId6G4bD6JT2Wnvy8FDH0dX8T8aMe3lS6FUBiKyyLTvUIGSiZ1PCBKmlwXkDfxd
lUEkLczBZvjz1SIdmHUvRUyl/D2wIpXK574Rr3jMzan5RYIQQLBduLdfArNLkw8E
lAcq7lHxeiQAUwmhAH4DuDODjZmstljhEIrT+IkEFMpP9H3lTJh2grGu9Zshxtbh
ZraoM4ibJWYhrLkBnTXXfZr/FDO8GmTnAK5QoTV8y32xmcZm0HuDJu3Jq2rrE+J9
JKLtx0ewEZRLOqt/uhA5QyZ0tZEp990b+Rl95+vy29Igl8giwSFhuurxvv28RUQy
9UDTjhQyp08djJ2ksf/wHkQKH3g6GfSICbgDNA28y/yvKMvwtrsw1aFjxgKSq1gr
ZlUuQdBfOtnyCh8aO3uT+7f519aprfuEri88SSmgra5oMnHFXdqBbRuG67CvQA4M
ctvHlZhaGnCQZYF0v52+K7/JunW+OQbvHdSDk69c97ncv3eQulxc3xSWL4+ktzvF
rlKB4bgs6vUtbupCLC3DoYkCjdSs+1fs/apgaSuddcv2NoYAsqpJKHU9hE6LopuX
ZxMwefCmVDxaPupmNwuFI3qtmAsNIcrlb6DCFW1YchBfRDbELkTzTCITQUSNMLtt
UJ+b4GMeR99BbkuulSOYI11i94GPEZJHDQkW7OkyjfELug79f+cg19DLtswJ96EV
vvipM1XJjgXZ1IxGIGoK+JbxH96kPwOgR5undFXigB2QWwnEHvZk+poSSGkxbyA6
CkK7H0FEEx385U7Ent3zsWtRKAqmPYvyzyJmMBAze3apjhsqQQdiuCRlC0totE+R
DNw1Iim41fjUH7MCi84auI4t0Tn8FaEtDOmP5ClauQj5sPcTs9PCaizuHmZk6IQR
OJSJEh6gXEUADQGci/8BblkpwfzvxDzzrgPoZqhYxoyF4r3hFy64ljEtXB94zXll
VkmVT1GwuRCYCk/vBuN+4xGuIHIQ9F1d7C4SDHwwg51k8KP6XovBx9FDdi+81RSP
Qal6+oC72hIhoaGh1y0aMjlc0YeXs95Yx69txJpeVh9gGriSPwh0B3Bu5jf9P7e/
i3+e7qmzygHplEzozbc7TXLzUGhgIDtJDsQvSIpzvTJYSWl6f3zGdSVnyZkmbImI
UgfN6be2ll48cCrqKg//UpUEKHW18ts+FLKkg6QQa083joizTQneTSinaXaAF6uP
40W20NPqH9pxthQZnscjItykfyszllfzaOPJjC7MGFD3AHWw5UfYW2+qUOZPf2Hd
snkQW39xu5tDjA50LkwJw/33n5lAmxULZknJe8h7eyMQ+R68iiRFupL8yXRSgfTW
CQVRGyGeacqSNaO8IWWMwsW2KoGp/gUGzJ1kkTfgkI1MuqNTgrPvnDOJALsYKj19
2pbCHkjWxEwJ+BpgpdxWmAOqryKGQBZNLGExwl2YknLsUWQa/8IWMIhVAzNFslRG
/MyoaGosQMTlR5bZVAAPq0YlrOAhmmumsKmYd3GZQfq6deAnP4ZMdtJwpGvLNjNP
MgC+lCJyroa4ETMKIYi6wWVl8CcSGoYQQTrs13lCEVLM2CoOzZdskUz+c5J2Rl0V
RsQZzZObt3eEaFDTTI1BZ50aFB9ebe3McZnjNnfirsCSFPVlhclV26LEoEO1pbeB
QtErMeODtTUOK4KOeIDDQ8vBY/bDBonh6AQw5kfC376GpI9o2b/wO9GUZGUCz9An
DUP22YkAvb4Yy2ARnhFkpQjlNmZEXOLXrW6mnYMwUuVhkRnEMUkwQIaI3tkrN3ge
vTe66ec2jyo+/MpFeHrRYn9+UJsmzZ5VfVoX7zM0igJKkeumIofC70DVAb9auKrg
wmnz0sOPoCPkHbARztcEQIlhN+BmMUNaX77/5FLX6coLggg59ygPaUM1260P4Uo5
v4Zn1TnT9qX/VeyvCt1CKsKr/XhoI+blbWGNcdWpCtgcf9lolDiW8kKP24TzFzGk
hQzloruoq2ikGwXJ0uie0SIkTvEy/fXg9gAeBMc5Gym2252006Q+pRB4i1kMHSD6
SZJL1TG9X6CV8NFXi3x+tEBA5sMOFJYWWyAKY1XVPRBmjgYIOrsGromtLueBDrLK
eVBBIBvQjSJYtG5xI4oiGza3zccs6aUpRB9w9QrO0fVWZRBaCibSLprvJePOpAWK
+rLnFyrBbSAOU1Y/84onWimVluSpOBQkYkQcsQKqwP4NVAupAhlQsOB4Ib4h0O8M
bI6dxEnPPmTxz7P3GwiOktKS3jEoxKvGpC/eBLg3Uy10TGfcEc+kqOWvtMgTbOqv
B9DKBo9EtAX7R0+AiD/CmeUvz6IJC50PC9kVs98tNAaKC3XbphkfB4/wDmo5ckfw
hb9GcgSQ5e47127Lhpu+nx1rKkmaGn+4x2Nf9KuQX6Bc9/yV24cyw2DUHpQT/qtj
vZIAb/XTAzxTHk5DZyu79/8UxJiChWIZH6Qd0T9K9qeYEkbv0AXqwENqpxNwYbxO
93LsMt+IM3GRAHrG7FhiR8S4i5XnemDrglK79Deii6/VnBjjv5tLA5lJe7y+l8+G
VlOeZ45EiQHFgK8KEQiPdBG4Vm4g7x2+tYmwQgR6D5w9vaQiXlwdYdk2uR7LUsDe
WuOZGGVxLl0gQR2kBIplkJtMK9HA9kFLYKAyDgk1jOEHGU7Boxub1Uqyd8x/GABU
PsSf92e43h4dwSkrlmK039h3cFptb6KTZQkZz1kEaC4HOq8dVIVPgiD1xboQ1nW9
f9Hjx9N8btZ8G7qf9xf82C4s5MEj1uJR/6x62ggPw6uoEswu8K5EP60atAWgj9E3
uOh3e0NLV6HsbqgOSbHj6ty3sYVuSLS68RYfKe12+yNfErML+qcA2S3Dd1IoOFOG
Pe3BzVawkd/7nUr55dcypvNzQUJ5bZYgDEX4L1vdpg7XroZotD4nX3hfouIh3/KX
zkruEAIJydC3B+/t/LB6zODDFujsz9kgSbohhOyQwNpGQKxH7SAvhYWCzG/JmQke
zwfswyN4dwWrUw4g7gnCqqkyRmQ2JQC8cul7FQG2IXNdyJqyTCviekbZU2TSE5K7
CteHpjwhyQ1lHhkRQbKR+yzvz6kxCsid5+KLl6uAuDl0vspLSx4okkm0LtVyh/4N
ac5RHDlwILI2b9pLM5NI4bQVr4flUDEJXRd7koq9m5N4wdkvKwwKSCEbtVTahx+E
0EuiqD2t2HFzcSXzgFhdveYYR2bS8MYoEpuzuoj5APtRPcTMoeLp5xx941IuwIqI
bdZlu+zk/mbOfc0w0wHOdSijz4V7VyEttnBbAo2TwHJnDVjfjzXbgcXRnC13SehF
KpoyRiuKu2VOpQQIhPhzxqY8sYTCPqHKJUUwu4Cpvk7aWkuyUTpOkUSR5y0Og9Xr
VeFp/iE6uKjPUL/Y7WHM6zbPTHJ8otSfOleICSRQ0BokdYqoLOR+pW4cA2LAkBV6
Ejq4dz6DBAZMrYMFAKEFskWm91RX7MxBWIiDuMjzs++s4kA1UoNkS0bRytflSp/D
BAlYDuRUgg6fJmSCQ9RPqU7NlcqvyQ4Ll8/2TxPkL+qPYiC1JbFC/db15rfFfu9d
AXrMnyCC8EZBQUY2oW+pacFXD1eYmv//ip1bfw3XAem9MahP2qZ3czbXrV99Tqtu
JbH4mkiOMVZxaY1wA/XhXHrlcEP2gwotcTlp150fUi8g2Vz2Fg5uZ/hQx1WvY2YI
xC/QFhU6YliVi6+usgok4j9RXo553rTj6RZm0jYNuDDDk9Fhw0fHylN1HW6GbVxr
P7g4FUFUK2xuk8owJz7x2pK1oUV/aUqX9iaK+6Gac6SSCpShJuF7oWfDpAMlFxVT
mbrNN6bH+M/1/2J0l2ryJUa3hw+8danUNx9XazXgrX84Tv6pQ7e6NL/0jD4QNM7I
fNy3IeWmHzCEyQ2Ph9ZKDIguzJ5tHhEvsiVME8cZsTycc3kBLH4C2iuBEmExg7wH
TUyRLKPMWWF/QoBe7DF9ymZYiQmlihNN9seacZzZ2P5xn06GURk6xvsGD6/zPKwp
+G7eZVxvqRVSb3lhTJhk2ZS/mPcYuGdm5bej5sDXSe6D7VynevLSoU7TxoIx5ydY
3V9ZD6Sp2n30vSSDivnzlTyCV8lN25VvRHGIZbDMIPTzSIYr7ILhd3UhaZ1KCTXK
LHBep1nJ2yYmUIfWZMXK2W03BMsnK2G8LBxgxsXnbzHMrWbVMV8oza2acAMAFUD8
dMGmTP+lQ4I4+S2a2eIOvnWykIqZLAF2p/7gfLvt0pbC2K02f6DV0Iqi0YHHI8dS
9o9JckG5Hd2awyf5Zz+ubT+0hRTuEtisdHoWnv5Di7U9uv8jBjKMFPqfFU2xXkwD
KVnNX5LvzK+7eavIbJ18BpJUzBAhP/d9ehFCyizwxpCAezzYwTTTPy7umdQGPfFo
yh2jty0hsnGkGZb2rX0wVu9/tGRncUBwfIex2TUwyGRdGjyzD58uBTGuD13iJIDj
I5rc1FI4KotNtQsJxm3c10CO4OvD2xntAEIvkNOeUwiMCPhHKDnOqoAvbApE2AeW
F7MtmfmRd2Zv/smvkZfHu/ccD09DKacCez1guyc39ARiQyovDZtsScHdVjBbWzcH
LHQUeYXoVHPhdDP4cnB28jw/J6E189tPoEOvQZv/TgcVBI/xVlUX3F1NAYC3GwLi
yJoGnEpY1KA+p92FtSoLTrxeW6a2xgo6AamppDX9GQuEtj2Ja9KVwgXpJu5t2Hij
X8EUXyg52NGQ+EN0Jw3qFU7mGjL+Dzqfl2onZhx3yuWykCioikOvkKvM91RDwyzI
uy3ESfjGGZ/f6+VY4NnJL7P8NLHUwxCRt6h65ZH8Ch4uhl0o319oqmKmH8Fctqme
rpgysbJexBIHsTLjm2A0av4XBD1PkvBljWi2rAUbAdn73ysnaCYvY4/faB2QJZ6O
J8xvLTYosb2aFCZ3oUT6NUhonGhd0c5RrKGLhS+CRE/eoTviZElsoZndEuayCYov
8ef0LYBHDAgQ3ARzP4NuYmqSha7JkLBLS6ABSA1Ou86Ud/Kk96esDwuPqThO61xY
1ZjjWKgr9CUVYEN8nBqhxJx5L0DsveIxY1eJedYfZFjxqcstTlz3ACiYpFyhJJNO
k73KnAUWSbXx/uEymTsrSnqiuuVIM8FM9/YtVmHKuSWBYEqVDbpf2eq5NRt4Ug/w
YaxRHKaold/1KC3q9a41pwDj7R+GVmhKtr4KKHd+fdtTf83AxEl+1RC5Q08CDQqj
PxhSsB0K3L23ZmfQ76/zuskXQCHRLlulHbiyZqnHXKWuqtTqGksM9dTPMGBoyJ1u
oC9OFGQBwqVxU+89GaSxVsmIBoHe/J87DK6xAPWksqvFBnmAhs+6BN/b6YKx4G2f
thdlnD4QVvMhvZXtMjLij33MU3MK3MVP2MyWN6b8+OFa1i13mo9UWxIcUPUCn0dl
DI5w722PS254dVWP69MCov4oLj6wBxSWbPq62YhVYmjhJLhdpDN8n5lFzgeKVIv0
BfXGhOvwuFSYwfOiKVphCDmkWzrBkIHnXhh0MN+bKKnpDHgW/dc9jswAiiqoG98M
qHATO1aVOCc0k630X74EmAiv972S0pFu8Y6aasiBH7Wb8Uc/U25eFyhHA+Ubr+ff
hUqS3ukj/IBwGFv82hYTf4PjqEQpzGrIh9F79YHsnMrwDKdQ5pmdOqGS/Oh3/iYb
HX9AgQ6ZrBXdEc1z3RBkI4t1ZbsgbrjxzjOsRxYGrrsVreb76fsR0WcU+8dAvTsy
XTBlFaQgqd+L+IZVUopRKLjub/8JM4E+Q41tgh/UpU5xJrZDadhFh8/WPmqEY0X+
dPAeeWrHe9j7Te5mn8fSW6GhcRLSTPMuFpS99U1g3eBrfCtZRGoEWscLL16bJzwC
0XEyoXurL+aJz4c1HsywkRVnZ5Nda0CwBrKt+x3qEjK2TG/Uio1XJwAYXT5gjV8n
WlRO1eH8yWMA+8YflMNiYD8AbOCLj8A86i/YI208GeYzh/VGiPA2bZ7YZr/vO5zB
1yv0Gbj8Dijhv1G6bxygKk9NL2GZjX/UCn5Hb1hRHTWMpS4wcbmaR3+qIx1etoe8
lPXuHKNXuZ6fQN8axMZQea5XKFL63fusIKSOXqCSQt0W1CVn+jECEBeqSFBBJ3aS
wJopxuOipDFLhMUBXxL2OOQUj3eGii1btxhxzNxvgU/ocWDypRBYnQHDnSklf1Go
MCpglXt0WjH5sqmOmb07w6smTeEAONN3Lm3RU63dd9N//wFBooEQ1I7lAlllhChQ
5K5DNIHuyaoyQrk6yQ1hHnJMDrdCurH6lEWjcszvzWQrk2W8SesUrl8ieHN1CGFd
g768FmpCkLU/9wG58NHwAdp8zrojHnap9KXJX8yyolbQVYE3z0zC7pgz08BlmUxQ
+ZUoQe3yFjGT6T5LyAPnDXW3KSheENoGR3ihL1C8okJytUfQeS3V1010FiE66Dsn
1Gn8I2fIYjuSmcK1UHlZhUTv1Ru8E1K/3byF7JIKgPNqxrwlS+U/KMDJ60y7fEw/
yefdV5hzVz4q2gcFvp2GoT0q2wrMzS6VrhOplNtiOTA5YB5k8VkR33bYfK+HmbJz
WUMA/obqN0N0K0Du5/n0dXzRb9V1UvvktHfkZJ+pngOrikzt3ojH11b6jCr4bx1y
HDHHwmCBbckVl1eSGAibKP10/Aq/4Yl5M3wyv23aDh/2KDSmaKr52JH6Rnsu8bmo
eRmRNWpJUreB1krWxvF9HGEN3S0uKQ1y6b9QVzREYw+fosUDVQC8UCYTbMZ5Og7X
uG7mTHwtjIGMi3FVjF53N43LUVl0dR7Wb+iaGpy4QJjvwjYxByGUMki1FBJNNQoR
2vNUj/sRu0r+MwRQYavbER/H4Lc3PNh4W1+RBHoxjHMhnJjcLgky6aPh6kucj0gr
71XSkaflgFzMFWD9JvSQIZZv9imlyM6arQg8XUY7+nWmq92LSCEsCcq97bVdf7u9
RGesZeBOfSZGqYRuPXVqFf+iKDW6O1LnP7nfqifTUrncoLk8l7d8lQCdncnToYfo
+YNGt1tqXtkQYoEj6OvLbggltk7TKg7rryVJ5M2tQg1TpnzRuymwbqO94Xo7J6x9
fkmVI6C7HOILxIy9S1oTJ48WU6+zdiv2xwlNLRLR+S/ajIyLeZT4aaI2b6fZutI9
QRpYKLA5t4bGA9lWIeTFjqwxmjUuvsmfA4GtLXau8im/SXG2kGMd9WbdIxw8w0AR
OHNMI/Ls9mQmLVLAwgAqMxpQWu+2KiCbZfnSisM5P0vwgX/jfKwLMxI0rokxmMRm
8KPIRRdURqshAJwk2UmLIWrIwJgWdv0uGdo7gggjgiGXJbuzW3CDtf543hsOjFl2
IXQi+2VNvSEmUYtR09PWqQN1a/eVlWfEchEPtbPHCgTPEoBkVhaYXbBVz+eIiwiT
J9h6CEst2oMwKTttecs4YG+4SicIIGm+YrkuyPyt86AdWCEi2RLZr1G/eyRTbX1g
AFxNN29kve1juuqk03le6513+iD9dkxJxFMHDQdfWPtkBIAz6tfGGGAjVPD5Soac
GcZlSYUQVPXD5XFQgLrt3B8fdozvm2VOl/VqmX8OPOlCKIp/jrsflniFmX4gGMvZ
hWa0WXm+WeagJR5zOE+x4xGh1KU1ZAqsK7YYibpdQMYLEOmiKU5g3GbE1KBqOEe7
S8iT90TgigbD6ehCXvyblgwcWEuplK+f1bJSm1OEp0iTNm9LiMNnZ2atyrwmfxLS
j4b3fA02Khwx0sJ1ZXMX6IOUwm+c+dR8D+0z7phr0zbHifZVYyRSRuBDUHycA5Hp
ACJy+ZfwqcL9KXoF74O5b48mqKyHD2SFeV1Wt71pxzF2t2JXluuCr9p+/Wi27Ylp
NFhoT+9qbBCz8ljari4uNyBl33XxPwnnoidB03+WWBchkeI8V3TAjTIJ7I+XL82F
yUH8ywXnukcrRtOjeMz81+aWuE6eFLYAZCpFl6zgialnjYkbpOv0phjxkecuNmRa
i8hJbs2uxAuw79C2eC3NTCBk3UvyFz0ZHjef4qUERbhTuH0KPFJOP/MUW1z8UeMF
Xlk+9Kmqr4U4+U6fPFHrcNkt+Aw+KfQIkA2RxWknznMTkP3vgXrgvhneB1tGD7gB
Tr3rwZ9Vvv4yKNM7dlm5R67QS9cwA1SsJLtBswzilfXNN5oMnpKpEsdHms3q9/yp
qXSMhJ3hp9JUAq6B4NmVXC2v4Ws/2WxewplB/cJtpXYbkgefH62yCY78LIVgUoei
SXUO0WFl7Xv+Xe2ROcEf00qwpKye4sR3Q4aRypNSI1YuPl2Cn2+fgcjmuiR5WXX8
el+1cvxcO+fMliWyEy3oIkOaEylgH+MYpM8B/ALDqnso1Oc7PgR1g7RlFa6txcOZ
8igISqvCS4dzVM/0rpMw/9TWSYw4Ztn5vv9TzU1j14x+DyQbJktsUPo58oQu1ONN
4fB1aQDfv8dS4QuKAEBZOExp6262Zh9PTWQTuPo7ostIYZSDwG9G/5Gv8UKiwAsH
2pH+K6XT8juF5dO/Vo8Ak2A6GIwbfOLvLy6XrB7ic3klyvTqgr8sValg9spWrteC
uqeHJKuk1pu0i26jE7BpSjKL4nz3aO0mMKjCKGlOGGQ3wWs3J9dN+ujrOVHEY+tw
tkyOkzwcKuwpy/eghP83boMITwLoNdmueWJiMgZ7K6n1viSUL2IzBl/MiNXSt9xV
SV0c0nzFOpfGs9kUtNMNsWMxFt24crUv5PDciRihYWn+TadLBIMp0qILRjv1DQiT
M0IbbnlQRBOhWXY2I6V26bEk2HTWo9XLn0R6/a5KTK8ly9eRiR6U15o+FN4HWJkv
SpHwcoZ1ZMCxRHLnr3NUchfVgtWl2aqNRPA0XOdI8t2PJagczYkWEJ+T6CSqAja/
+tp5Q0lHPN1lK2FZf1yJaTAXr0DEOAfQqpDIebj0m72KgZZvQWUQSHWq0jythePM
+1IBWL78S0q6Qd7G32KyWGZuoH3CIbQ1Xmnnzn/4Zi705YlCV6C6TeTIZ3z/nA4g
AD8KvpqLrzSwEvztzuMu+r6BxAh6leF61O189i4aNQPjPJhLx06kXJUxaiTu01/i
1+VOjWXZ9JvSeDZis9Cw892TrkcXRKXUmaCjDsgplpKrkZMSzXUsOqjutctKY66h
zkT2mVNTgBfxykSFmaGHwaqZ/mqlaQqpZVgzHTUi415HV0/bOjLhwu63NB/RGua9
BffKjbJ5dwQf76EV9xVm/4HLfrQ0sqkBCNHKu2Fuypr+/oBLd1gCjAMKEe1f8mbd
WJyfP+XvXZdkdxtGobSV0vQ8wg9lHTG3vgySOatFwAgpIEtM7HV5XKzLU3SNgCi4
jA1AKuHmZs46YF0Ta7XyhjDPGoPFumZKvBEqMGhlG1ZfwryT6ZZMFq1fTACaYlVJ
7Eo4R0GCnpBldO7Fby8+tD+sY78/ti0fNBCouuRgOo++5CAVVLyGxJV8Gk44H6D7
Dqkqacj1nylR9QEWDOsFY57DZsNIKf7URGFZWAXhq3zYTVoVHVGLnluGipjgWDBs
5Ijt4X7YeV2kymI+WCYqd69G9+WTpV+mbFPtLvYdMCX4EQ7aQWk85jieIW07rFJv
t/l1AvoYHvVfvPwD+U0ernpKmCL0U0eAOhbH00W6KUbkNarSb1EtMCSAYVIdyJ88
NTgjzYTJtlFYm3TAfMx/bTJEwVAugBCCZP8URmvpKyV6rOsYx90hY/PHyC42QYgk
W+d9vTpshSG75loIpquKmpljQcxEUlTy80JE0JhULdLSOaS4djeAtZcaprmxLF9L
6Q4jhW8oMd/kVlRpf2CushAhDwoxHPt8HetJoQ9CbpX92cHA1v959OsjfPj4IbsJ
ABPnOCU+Tvr/17zm8FijqlVdukFL74EqZqZmyVDRevqDgX7c0frumNO2WFBOPHKE
aoQcuvxBYnV6kGpsxzRWoMYkCJ6Kytzw/I8hfr+9IlBqkaT5EXpylufbTHCKFDaV
XOzWdcpMtnlNc2WohhWL/dS6brrSKyb8N/9vQ1dfQv8CZKKW/dAMw6XPewvBUUEJ
xKKwJwEys5wP4PzATQjCQdrIzeelrzdAol81f+gTKKQupofldwx3/RVMR+HKmsT+
osnbzxfr+JJOULFLWdg8f9n/U2mk4NCtzvZqycVFircMe6f6T/aF/NdkWSK9uyUw
Hu03Qts6dKTBEdPM3brY5tPYr4NX8DaUds5rcmZ4oTiSaNhBVT3XcywAZSsywKty
2Qlx8XyrvpLD9zIATTGasDv0ZFeb53PC576RfQM7uc1SZUHoipujVzkwfpiOLLqD
aEbbq/EsCikvh+4dD1NHBAUPEVHWLEmSp4a1vXH/SvhTylkO1pWt7jiwG2cRVEPs
i3+H7zwueR7uGNd2WCDCtFKmeeQsAyhPAcmzOv8hFrCZtRDf9nPEdP3zx5Wtqoq7
qc+iaZDVszg2cwkhmF8sSt4016KqA4ywQ9Htl5dou8OJtDCAhHC19Ehil3uG9ATV
U8JQnEXd4SN8ANsovPuinLDO+fKEkHeEPNrGR8XhdG7lALw5HEq7evn0KLVeKL9W
7fcpUNpEfDKVifoo5urVEDJwL7EaMcyWEeg+PA4zXS+mNFeOGeERV6+KnEIBcBee
OEe99fNUWeotUmfZbpnJ6sSe0OElgNXvxIoygYDkRWNEHLcuAUEAEgU3FwIx1acZ
8HHnKRvW5qrSzM+fcjxrLanq/dmvBWm+YsZ83CG50rmWEqxiLTvyy1jv6uV/oC2s
dQ++qrJvEkj+PzB+IgA/3PPdkME9q5Hkw6eJZgzm5ltG6w9EL69QCd1rzqY55aEi
NVn6m3Kw9oBhmZ5vNlxhvy0BIyIRx7QADlwHTybrtlKr+caIQxK85ckjyPLTb9mO
L5Iv1yr5Kh3LFfVXV5JX50k+a7vHl8mTPkdDo0D2fCVptvZsqB5Tjs6eMBeuUFkp
/VcnIY6RsLBgtXyeHnci5Wfg0ZmupFdsEVmTHiZNK50C0GApr7NuoRL0CwRIkGQ4
IoUJ9YHT2Cv4EqhZWre0NjNB3t0B+BUhimK4bM39q7yza6yGhJlpCVI8pHx7cXQl
/0n5QKuxtLDjwJ7unD6BsrtrUDZT4efsjjRVDoKo/uqOScF2gtibtCM2N984iURO
r3Yt2Qaf5qpaNaUu+UhPwdU9pc793Gg5l46+ToXdBd8Lq9YQfes8k59FUgQN536E
ttK5B0AytyUjuFAYqOfwWhgB0NbsRXT2SucpgRbrw1quTM4JrY9zv2pUYwYktirK
rGUxdq8wKBx2lcwLfaSaW/oJFq7ZecMzF3UN1mOWKXhDMkO8iibV0THfEV8dG+ln
PjqIJA8zvo0nCC6qxR2s2Xh2DRRCBHd8GKunDelHscBNeahHLPyPlfnQ3vFwrdM1
jCuNMmsEgbUW44Led9BpVG2StolVVXJnwmJAO5adWRi2jFMnrO62r/hfYiHMw+g0
hilTc6EM+oGEiu+h4qEFGFtrc3jmMLY2ieZ3JVkFpwMwDk7yQ6HOAVASwFb6Cc5x
PnSasEfyfK3twjE3v5mKtBetje0QSlQk35ZYzIzbmQE5izXnbGXMGsr0BrvbIo9V
RqceLg/zn1HCbHii+vbhOPiutr39dn2+ig/YHYWJzEekPGyP7fDww+GQkfz7ubYr
NXwY3Pw5zYSMGj/NFjVICYWdeLGpSUrXYY1ux41V+BVa1MrtvqLmkvIArEukrgWA
y7sasIIx9PM2z31C7uoubE8M7ShyXUfTJCUoxardkyU/wFDEqUbRoLlyj0vPkDmz
ef3jG4NqLVbfyZy1l4+OMbOReY4qXQUEJzSzh0bDJG4/43MUnTUj7AcMbMt0IAwS
m2HJNQE2CK5aFc1P7hA6KrvXBL2o8FvoM/BbZR0NFJ9nWtONEAaM+i99TFrYxO82
POUGterF+mph9kCPRTVd401oA+XDZlAniX4iUb8DhqnUMtTrtbxsf6odMaI7SQ8n
h3Px2VaA5iV0/1GAuWrAP5Jrgbp5PE1hOOXQL0Qk26sfACExYt9+tqim6XknIuDh
qjc5ttt/B0mz97S2vDi2rVvsVtNTWlvr6tbMRZrIQY8Hx/9jIhTNzNGK4Ha4w3rA
YPWgW8cb3VO1eJBNPDS5lwXbcGl35SIV9/ld81rRRSY1k9H2dV6zn5YN5MixStup
LDP8d77LNZpUb/fW2P80vE8iB6nmam/4vyt9hqVFElxFJ12E1KB7iV8IzfsnKpXd
o1zqkrk0B4klzmp2ppFVMD4G7HMwYK/TdzWZkM/c7ztiWdvQgC/mnkHMju15f0xe
xTTFfC8qRapwudzqLhZVFeayIzZ5GdW84hmMj/scvbl/DxW4AIBpzMN27SgUF/Wt
u2AbCHn/LBxwkitKCjeo3RP5/kwp/MgyBPhS7/pr1cmHowacJodyvItZ3kn/x/7/
Cvf79QQChoG2qxu3+hXBDXm0KBNq5fuLpN3g8Z0AesIGgqsJoNHmD/PrgiHKa5pt
R8Dk6PrhK0uqXuKQ7J4pec3EOCj8Tt4bZrYm9IqFoCCZ+9qvLN3anQA6l8xbBA7C
aNYEM5aA3bhRXfr7PTe5W9QbpwwELcTAInjDSX7XamAeZTdnvquIio3Vz5PXg40F
dhgzxJ4hZchMdw7AOzfFTPYCB9EdkPn1933L9x49K36QxANJ+ayAJ6CpjW8cZ3RH
Yn/v0My4pcXBqqgDUClgBmGfqYPlQQ/XHzuTDG5bQTVu5Gx9ev3AzLcfUDMJVrHq
BMj2rEhRtW5Fiv9ad5qA4RSxftJKHAFwt+Gv5rmRCo95tOzykdW7SSVDMys7NBzR
D7886/zkwaWNJhIgVht2/QqRSBxRyyC15SdNIAa3w5eXUEBTN3Q64Ep424HO3Q35
KEdImXaTzjWtBqIDDvgbYYjlWONZrrIYAxDq6pnsuHIuLLb8nDBfhejCxj4wPDJr
c3AqdRGX5+KcxStB0Ujnu3TNGXseicyaFJHqn4s/4BN7VnDFJl5eiQPqgIVOLNt6
6AIp/S57wxQcuoB7A3kHmJ3ndO+3WGcblt9dgBB6nCVVk7k21NVp2Tw+tVMuFwQ3
gQKMCoOAMhL4/yZvXcIXzhO57hO1sGyoiqqXaOe2lm2jR9Jr9pEPOiBNl7WVzwOZ
KAEGjZliCcr+ZGovO2QDAtAQUJtm/cHwWkFkDqTKlcEHqpRNsO89bHSnTjdyD9AW
s+wLJh3yvxUhlBOcm5bg+91+QtwWtpXD3vLd1Ln4G7gntXC0Q9rBAPD1ODoYY9Zd
kr64BZTudCude07ijmAKklD1G5gwu4+9uhOQRQBE46OExOgaDvfztNG/W1oO/Iru
DmI7GZ+IqfhfRBgLJ6ubN2UScxt8auMKBVKEvcT3yP/RtwqHfK4T+JSZZawmTo5M
Vj17Q3zdeuw8pxUsdCuEeyr50UWsxRJLfw7j2WAuiuEC97rSCeuDjRpRVsiYJs1m
4KKYsUNr9ZjEWM3/tiPvPUJbpGOm2pS+FAuSHhZFT4VecHp3JrD40kGCvdi8irxD
naKPq5MdZk+LtHhWPkVDr+3AbSTE4kzjlvqFVAEQmk+Hg24ghwkpuxLECqLm7G3C
b2iAx9Ai9CndVzWp+YS8y2oWmOqUj6Q+V95fFuGh6xSrJmyxwOT2A43ZIui2/NrP
1MNelScxA4gFmpDPz7aqCVxQjFCmFDPrtxLAy968zaJXn0qJTaY9DkwAftxmFkTj
lLT//M4LQ4LjTqR/LJK/et6v6+ky5sXoRc2D7FLnuhxWDS3+Jjyw/Xgt5gqLML2F
XWKWtLhzpMgBKSoZq40wySA8JgXt3sfIFc0b2hE1A5tcaOQNMmMudGIwXgLTkCzf
Jj+HUTVYep6Vc/Sk5T0XMJXCqCiSszRUm49I/19LQyWUW176q76+QrLBcILFlheV
bpwKHkXekb8i29jWxfWrpPQBcqJGajDfN6Ipe3fcGhVw7hFKUZusYbGu6/SderVX
NpLgzc9bOLQyDNh7Y16Wi/ocLf5CF/QTX2VL9XvrrcFwmStYz1qgTIWSnVu2NnKX
DrJI4av9fwJCYHTpwG50/Bcd7SNZKxBShKxhY+myR7y62PEGbwD7svmL3pZ1VTSt
Xyfme+qesJKktLfBXZQ9YzOd56/BXvza3NSjCjJffO1aooqm0FWEruk96xy+3HAr
6tD4wymeBCTqTSqLZHM3zB5Am+yjKbMZ+Vpo9guJ48of9yNlNIiCClDqo8yC0fDS
VRK+/d83dR+IP3GJDm5CQXxX69YbFOXegSrUoESNSOISryWS38CgRjNEkrfbskFM
jeRVMJAmKxfh2cpJzwAWmhvkWNSUpztU7nMhkNH6EpxW3sj0/yc/Xr1UD3RTPZ77
pnnnUpMp9sGjWWCR0iXttoleYjty1E340OHbIa/zmM4Q/VjZg2QhCR/rPYNWpWIn
dypisZEahwYsjyRZqVKt8fccdKBWKar7MP8tFzcj7Qq1jMTXPfBUDwtAk+WYRr7w
Mh+QSHo0WxIKzMT/ELO/UVdXrp8/Sf4OojJoio8DQeH4fcpGfPZJmsdMAs090/SF
IcpjtbXP1TkwYqoioE06Rv2KYbQ1dvECjma3U6ZY/pZ3i/LS/SivmPpSweecHxX0
XOL4Y30DAf2q3Bl0M+MZ0XTCc+jHwYV3Ec2NOkAuzQz3XjNsjq2o+xavqqY2k3oj
dfne6nQbxDVgWIm6cx0iNBEyr8PGmlJKyMZAPMFv9WMs28lfmLr6PTBg+yWxQnRD
UpQ3wst2gAkgXaqnighyzO23O3vQNfcY7DSZ0wb/RQHXOfVIEiwrrZFVqw7KWd5d
Ygzqisac4h5PQ8fKqNYb9hKkLChXixKsuMuWhaO1KlLHVVpxSpr5LcLi/MNT9xb/
VhtLQcB+ezHGWtbu2Ejf08GXryfpjFQJD2ygypRPVIEbO7e+OJ7N1zfXqUH+Av89
M6PVxx7lALUNTSQciPbv9ZPXyn5V92wtznwkGTRPEiEDh3E1t9ZjAT6X+attturX
P/5pLfW9SJXx0o95HctqrTqHxjPyaP+WJZZCmYv6GZ9g7WH4BmxoFtDRGL3rYLcs
VWBypl3X7hMOJ3BVV7i7+rns8CKbBeKNlw5CGqrX38ZQXe4swCQUwBv8/VCCMk/8
e952lNgeVo75IaEf9kDKTOHMGGgxdILmszhaFYdiPrJ6qMzNQR98K36M3J8aRZfJ
fgn/wj33NVZfQ75/ABhRezEqm3d6wXcaCRdTALZ6i271HaJ6tncN7AJVDgfikMvn
fAui5XR7a7nFI1FjiRjywDDXaZWrPqUMQlykSHjMPHZUEIE1ftdiZ1uGAmPHrUS/
OoQ6p5JS4G9H2xKHJPrYCzhYYbAye/gpnLYbfiGKgR5S3WOqFSRT3aPfdZlNVMfU
fhDP6InsdIbmUHhbZ6KMjwUDT/mIBqSLZov+E3QAEXbWnoE6lo4rRUQKX2lM/yja
ILdTz32qEITTRl2kTAITvo67LUbMEFK4CFiRzutr5zqwRb56T8UQRzTlUHB3yQiq
+wkwoU9CDB3ALGD+T0+SuyW+TBFuqBjV6FBot1yABb7RbBaDFYXFT9aYA07vRISv
T6bFYgroevfS7Enxxgmxy7274qP/caDYN89e5uzi1YpKVr2n9qtQ+JPYdDGC94I6
8087SCIrevSFHEYOS3GoVD364jwrNO/GQZXrsDEO3Qzg17pmyzOo36vkye9q4RlY
e8byirmlYTzZvUWHU6zN3kgcyk8jHOItEKfoWylQ6w/KaxEk3NU0U/TG13xK+DXL
O3hIF03Ezu2yH9psni/YFkOdJTwUvL0xizNbEEfBVABFJIkj2M5KB0taHdvYm6sx
7nZ3cOH37JFljuI6ZGVZY/oZtVfUwH5U04uCTCINKQFumznOtEq8fkP3Dx0++/MD
JFnGAnVhRh7+WGPhcaCVPoZHVIhraS/WgAf8iEYrITSPrsFDPHNTVYAgtPHXLNCP
TaL7VB3VkvxbyGtZYgB7+4KME4ogQaXsIXSCJaUHeG76liDmFqatstymL+flqpTn
D+DTyCTErRMm4fIAYEh3bIGAl5caRBnAYSMOQDQDyAFhKBr8mj8ajT4WZ1OeU/Xj
HcDoRYrJ3mx3QuRfXFoJdv2rbE2jmRbN7FE7MwLZf79S2KhAU0KXVoQFbrrePJCe
hr4MN4GraVC+UJludT0aVjh/GkJkZKBvKRnHbhor9IzDGTOkElwkDhWPbBayCLxx
Ynl7fEbtv5SIHiCke5x+b1q9hnYmxgUf8yqXJXxQcEUPqp4Dtfbb6Fqqu9Ut5nLF
Lz7qgV0s0c9kUhC7dfaZkBkz+/FM2/7h8/8tZH6wnKtXbTwKOKw864YINjbUIOQN
PKjurfC+jUe7vfbSqzsA3+0HPJmQ5Hbx/Rg6PCQaa3XrW2nDyXvkXbljWgGbcxMK
L74N8rq/Yg1M9m15tbDg5NjPZTMvYJq/msk8iRIg+n9DIpoCV5DdTFNHJZPEOun+
sLiSz0MYzsAusey4xEG9Qlkvi6PxFcXPB+ytvhiuX8PdBK+XPXo0E3S2InmsONcK
mlfPzGGGvgZrqXRABowOK/eg6qhgnw5ZBpMAsGHClEw0hVC24p/xhuHhTvmX/lh3
UnR4YnmGErt6ikA8lMdTsOfg0Mzp/E6pQ2WdMKhB37/kmIoa3yOtYAM9PTkJHtgg
US9pKVeUvBARTNvga+NJhzP3I9WkSkSNB0dyEY9cttNNTYg8gRUTeQfuYT6tBy7D
PtMMHgS+m5F86co2QtMKhqIWaC4/8kcjRGzobHr6Cg3icHm7XhzU0s9kTQaBMzyK
cepu7EB3XHnEupRAMTs7iPU64ocbKapfxmMGKhJn+CyxNQZhjsoykGuc2mqD9bY8
9VLTVWw26t+LXkGYXdBd3q+5sGoVXziKYofG0jKTbbEJ/VZrv54VoU6q2Vio/coh
rvoVUe38XE3Wrn2kiGpf5p7Op/LFtHzMS1Bvj82BDuzyZjJ3G2fo7yUSSFQgnUJw
Bvz8jgonOEVdI86Dx97DTE4g2GpDG5Y/uXiq4ho5O45RvrkIwp1e9By1n9fPiQdr
anHnx6fAv1cyZfp8wyn8N+77zmyNUuSipUrk8lVbQyOmMHqm2oTkpRnUGDGFm2BO
tMQzV0YNYA0SBPA3TriwETyg0y/rrObu8RB3nHrvAv17WL9Rxg8zaBN7B7EvD0kP
kCPQxDkbQq9NSA3Cewl3aPxCcm+PiIKd1fyZ9cIdkia1V/uUO+5YQdoray7szr1L
yh6EaqWj3OnFWJrtlDafpf5QXWMDk1YukV/Rq3/g7wEjSryJ4OVq7HDI/VZaYwVb
XltTkUU1gANY/jL/kAwm6HHTwkPzbEpUatDiAh4YsyvZbPR7ph53kYbHES7PezSw
jmdpRZvNntU1rkJHuMxiq0pa3hVglnjVcvi9D+CU5G4rXQEJOmQxFAHzi0Gz8N0T
1HezUunCekSj3kNcJKc9ex0IHbwwmdLj2XRShqlql9SSvYmgEsx7eqw6/UcPhEoi
ul/58JZIwMLLWiU3wbBO0KI03TuPFnlU1Nrh+a4vsjnbYpNge1PCr1y77Pv45YIz
Ikrcq/S/NdfkLO4djfkHGmKdwOGLAFFRsKcHfLBLaryLu/n1f+mBD/SAyYRlUSpw
zhK86fWPH/wmenvZe1BU93SrOaHGnlDuNVwtQUHyGvxtF2GNFOr3XdYAm1gNolUw
gN3DJ/q8qXBGUN8mWjW1CU8+tm9NmwGEP94FGCRi63SuqoCDCKkJxzHbDsZULfos
R4qtzYgrHQ/7bvhEZ0/zMkrv9I4PbdQK7hFXkeH84SpAaoID5i6ZBgCokmjJdmR6
ZI9N6BBVTy1k68CMf/8AOEyWl9ormnAvSjKxF9nHj4eLXojH8DkCSvNwQ/3fMspx
24DdVJ9XxEdzIus6QJd/aQCcNxi1BpOipv07MgQQThQPKDovoN5CYgpYKyqy2+T2
qjkJfnMScDRfZ+joaYiHDblnHD5NI2n7psSKuviYfu8owaCR+fxU5yeQMGkycIl5
tc3g6GmrSwTAxW0k9JG2cwSGJt62W7Y4zqnSOagZTGqumYqtBz7YlDwor8GGN0ap
br7aPoAe31V1UCa/Ol2tlEinr8SniCZwYbQoVLFeaj/AE8pq6WrfzFR16N9myOvn
S/i4Tw1eEsL5hYdHteoWSaJnAgnKgaYoNq/u0QvSHjk514gBwIX2A3wZr6E5G6rq
xWasC/fWQWZjoxMHfUB3z72XVd6P9Iv5MRu6AKf8IaxM6LwlLQuJuImMzax00O5G
z+IMmV1n9u43ofcgt4a86yJ0Q1536D1+5wHHpmo9SaSrzOoJQFj7Rsd1KJj9R7Vg
182zPw6vpaHKrDUPVpfWdyvAWrJ4NXI4T1p1LY5V2cvgQPqFcUXc/mRrOG1iqXJ7
ltQzQa4voh7HpGTbNj3h2OmXoZyZie0A0i6wNxHrvSAb1Ak4GIo2GhFkJesbAt20
SjNtJ24oad31M0kxm+0nmUaIBvQL7PENKbBRpGwoJaIAxFULLRy+1Q182MYe792N
y8gQuRVGPVZjWpFZSROdGUjuTcuufPgMwkCbG877mTeRvQz23o9iJnqe+scP+mrX
LYT6emrE5LMwxWN1BJuowg9n0BYZwjClO6ChWfcBUkrnLblWej9TdOE5yYhbqoAC
+Nd1tLbFE2OMfErxj9jwavPfNdc0ZYXb7cPGQPTmAbfbr0pC4tTRc8G9Z+zKXTrM
qMTsStVqjhQQtcKoGoaeeTgSQrmX+fvewrFyAlfGJfsbFECh8M+KoNLJhxbkQOaD
lys4qjiTgYCS2C08rPg261fKvGdyiFuTrWlThqQ3I0gpZo3LMxvB/pO/V3Sj+6kj
ynMD9b0qzU6WwLpRkey09PVVurefLgGHGHUAnDPiCauvlaTrbcPZqH0QhtIWh9ry
YjfdxTgfW/stwZutNsvhR6MEuMIYUWEcazvhWMi5sv8GmlSE/azmIikKLApOGSOI
nKsmq4zdDB9LrrdmignieF9MBQ7NNJ4LQBgHgim6ayCzdEgCoze2XAsQu/Xf+PHM
J31wBfDtdz8hyX4S6Fnbwn6WsfD/NK4we1XjUff37Wds4QiKqmBTmlWNECJMv3dl
KJUMTIA4mYjfWg6nPqI0QpO9pDo7i9PJ1byIfZV30ivsytwp2F4QRU9A0k6m+P15
p3EMir2kyyevapGmf01HqTfY/swy4lBKMb1VCljwcuo8yPJ/B4Jd5d8aU0o19XCf
zV00+3mVs5JT9/Z/goy6Cbk/h6LalFms9uEJLOaLgQlUrkJBhDpj/Ryt4qEuVwl9
OyNe3L1YXfE7g93aCITopOk3HJxQmEp/fqv0oFVu4InIudoO0IK21YDmprZnNoS2
UjRvRX92nS3VuFCTIX0QLJ/XCUsbX4YOZsc6o2VWSX9ZDWn1Gti7JNFXirFkXncJ
WyOMHHGMevtTdmPEzfTVl1zlVtemkwyEdutPiUBJQ4jequJSK4rdMQvkEd3QwYEg
xPTbJ7MwLL3lymKw8r0qiJJWLufyItZXohQpjvYK3WCCsximSfDWnk0hKQPFU79k
vXZFV4Gj6H4wmsZ0e8HDFQbC40EcX22WPSJfG+oWh2D4ee0hQCQ885846bcOrdgT
WqQ/vz3x95K9AtSZZyrFFIFPp8AOmaqQeHzphA2rDstYVSeI5fQb6kZp6LfHxjIh
sICfRBIAikgCfvq6VvPIehv5ozjw8vctkIVpftP2Gfa+gZfJYC8SYjszfFfPIBKW
vm41dQPYVhE/DfyM9UGZGoX67DR50BeKZOKALNYQHt/fWylBMpRChoKNNzAXww+U
2LaAMgMDhEto/EEUyxiFsFOXfl0WuSMpL9twcOIbSX/GrpE/d9ht3mRun0jaT3IR
01XHmMLAdVz8493MZs6FidZaNQPihmiyQl4dFDOO/eCs85HB0efAeUJgBHxzv0S+
fFEw/LC0yoKRezXKC2/pbBwFtqq4kyAcA6uFG0KvFd1bCsiQGIxP8jhi6c3n12br
o+ARyM2s6Ko2wr94fky42sW+TPSqQLiOg3ghr3tl+f4sT3zeXjZQIE/je/AL9Ilz
jfTG0bXIdyuHXyxomVcVmaSWZPaXQroT7+B2JWnL6Ipi7o02hHtOhbm93xaQWr/F
I53cQGJK2DamRTQqWHUgC0MCC/qHOxTeRDTSf2Vtu3FjMLBTmtX/x/zD6o4WQQeI
CLC6XjUmi74C0Ofdkh8uO4NyEd3lwEJCHZCEwPVMkZSsiY06Sa422irZSPA6vFbz
A9WnhmMZFAtJCdfc3pGvo/nkeP96Ty2lu2xqpbI8rF3K8c8jW8T1enJlazb9o8ka
HB4pqE3HnOBrhXsyAaXczlUoi84cWZmadzQsUMCqXqioKC2b9Gw9PQmhAuAYvwyO
68U4kjqHypOa/t+n5ciS4SmbkblWhkn6wZuyPM7yXIRXJPYgKNuPG0y3ZWae5CAi
4BLQ1Jub4N50YgtUg0Goq3QG4AMhhA63oVo/n7pLy7gGwudOqBah3piEB5e+WKzR
LDv2675a9KmtMq0OlFnhcrhF3TLdTL3IC4Vo3urgwHKiiG3UXINPglY+y45NH2zT
zEBqIvHaEY2hjLB6ZSfCqZa6bOzaxN0V0aE2OnKorFo8h2joRapTCF2RrGoBY+B9
qJ++GdIa8FHc/mPI7Q1MLhAdVr4/AKJUZyu6GfUyLEa/KivSXebB6CoWoUa6JiKx
T2dpCrh8IXKDgeim2HKYItQrkmy2UOkfcdFus5AyUG/vxopp7OqoaqIeKw8TbE+Z
15I1epDIM6fv3I7hyuUd9DKLH2Akde5k2z5qo1bCImDnekcPW1GCCQouAwpCA2W1
WPfEsnyQCUK2GI5FEh8QIN1MknYVzucDgcCjYSREhz7oitxYtv1naart8ToM+uk0
ASiNLzPS7IbA0sCb9XZVNqTKZiioSTOjPrfba5b91h88myacaxStuxsDuF6jUWco
tBYI2O7V+OTwZoq3Y937Zz9DKGBRwbHB+6QEEid2pyQlbZN6yhpW8W/RpHkK/dsR
vlayDXuKzflDKuRP1cbochAW2Hkr4cXOnyo+zPkVZGjwbm2DcqFXnzMN1VWGzxr8
3nKJ3NKgDXWcCOts0t7rIjm9Ch9lm83bJXY969rLuPxqd0lGBFkUXKoXGs6xWVA/
9PdDJfsanQDjt2Lke+19lVl8Izwu6b6mdpAqMXbTtuFAVUk9GPareoK6g5pc6BQj
mt/eUORisGKnyV9LZXj86f29Y/nxrsJSp2al223CoQFkXVtZZW+wrmqQm+IoZ/91
XUBd6fh73Jf39O7yROV1GCZOYm7QEYfSEUt8dD06ZAOXVM59o+oQ5NppG/efx2fH
HmtpRnHCDiz0myP51qnEXtjA2o2atbOS3pnzlSmC61+xM1UGsDeVbuYqVdYSEM0F
NSeolpyVaRL4k9NbyUBrPtiwX1lw7oMSc/NGvtEDyD5bjehb7xOZ/lX54rycyl6i
2ko1mOp+bgFRfqCmAHw9bO03Uc4QFNrPAI7RoMCZfoM8LjLklYzcfMJi543Ij8OH
7IFGI71durnaGXqu5TBl6j5NLXRITnQtQ8UffG+77BfwrwGUl58xex2hF3KwewTA
e6qtU1HlUzcKrNJnF98j4ba/gT+Bm1vROq08HaOSQ8USZKgn0lm0Nnir37//wLeW
tKUBEJ4tB0t3rImDlrgqU/a3pXI0muulS1P7diFyAH6uVVdWn7ivZFTn5bm6n7bu
bU6rpZ/ulCMNSwKq0jkGSd49WqHoWDh05Dsx2wexTHfc9XfoQnxewz9EtqzdwWI7
yrMkmdmsk1cyFrDFJTG3Ai6P7hQLUQe5yxq8/A4Rj4s0uRtXcy17hBfNxJNlNxS7
32leJpYqIrukkOQ5uk7+AI0uytkLb7K7BzPUbDw1a3zTyfEYxWo8K54ABPX7GGzl
Koxx4PBc0OocswVwr/NVnJKCBETAMPFSNW3qfxPRyEZJQ+H3pPZBjbhYQrz//MTb
KkTWPcTDa8HoL5vcidHT9F4U9B8EXy44xx2zd7v2Qm0pECaXbVtDgEq0Yzlw+9IZ
btXTRDhHWzAPPVJlDxFP5yDUHinvBgLWSOHLjBciPkP+PMfWQr/hBEo0Q4iqAklP
GQ84vH22Q5Bdn7xViRRmkMG5NKF59ClKOrME26OFrLUa+iw8xWC2uc3iHiokLpSe
DsBY7vPs3eH760qrafJ7KLM1NUi3BG+WCKbZhlh4XaoKdHb7NcNxPmUxCC/Q2mF1
gUlmKVz/ZuDJ/RzkNPFI4GXbypC9sHIZnDSTy8szF8+v1SGmCLGEzZQNEHwvqBPc
h5DEe9K7lzXRr6zKrGHBI/KnRUtuGRgY8F6SopMfiql4LTsGi+CXebMLLvVBcn+A
V+BE2sfMhw3LqEfNEDYoJ7Lx31YYtOVk2ydg2VRZc2YCfnE7xiQc9D+f9C0gXgMs
Cknjc7HztjOrns1NxwB/1lpuWByUwpb3WoYIM9LjwUXa+MxrzOgFD7poW4Is9bNb
nBaXkNqzwk8IYJ2HhWVY3R//DukYWljX/n2DSvBW9GUQSx9XIyF7JGmj7QUaKDer
8J3J3EQeGeSbQkWUuW/c1rJJya/Bw6i5jK85eNzQk9w7Yc1gPu/jSwiLTuJzq7bG
sonhOYq5PEMC74nQRlEqP85uHW89aAY1ZnDSFgXw7TDV6wA2eAB1etoUidqwQi8x
MFN5c5qVbwVQkEmx6UviOlOBr4gewbEZOI2RF+LTqOrihE/SFFsLpQZZh7K2Bm4g
THKZLM0gohSFDPVRqO/YBmJPWHUECB/YWvpECxwPXUtt2L6RP47V9iWihGtmDz19
iOKcuTH3moeh4TCYZstq/3hISTtGcy5qjL14kRABO/iLoBVA4Ts4P2okZASHXWPt
W7wipz65fmC/3ZrE7iwJajjAKupkCJ5289qYFyfxalLfP7y3chOAWBxXki9tCxRP
CnSNfIbsamZAjKyn1hlWiUYYz5RcBshurxAXY0fwLUPXkZF3+hyBkQ0htoW/n4JL
tGnr3g9rmbsfAspPOA58VbM3GFdonV3CEl55V5miSy0hG68SU4DyToGFWFn46cky
tGmljKDPP3YoqsLXj9GVRFySa93EHBaTP0ZWeS5EKW08Uzv0M76DYQI4W8GUZ627
ksyto9+ExCkXKA82yu4I9tpRFF1KWJTJZ1T1SvGMZkkkZch4JZFr3I0yazSuhmYa
3bqbhuG2hsUJdw3kCCmgnwpfiECUbIecXL6ZrZ4cSkXPk5TS/TgkJhWhPN28Vx3B
mlfDSYTvdYgYCQ4PVMr+d/jUyFVYriJNoRGvJkNQBgOid0qXhd87evKqD38JjgXN
nCAhgjHUDcxc7M3AISuI7z70U4PawwWJS2tkgp3zuzyZyjCo16BAo9gtllW2H5It
D2iqmSHDN8Y6+djLKEoM989LzbgMR/tR8XS+cZIYwdYcSYSz6/s9+DJG/7DAyAVe
wP0xmr3xOrIPyuV0j62UurnraIb05lq7FANkf7gBsgLzk9NuI259407G532zINwW
rCTqWzVgV++PjH+6/du2MVz1XdQWsm6ZjCHE4Dg/kWUpVA8w0k9AU6UXtFqYo8YG
cskW3mI3Iz2mS5WdVOBJ4iNeaqLj0WyoNT0pPjv2pFxJsjeIiS3KdcPJQpSbmlxe
HU6nOC8m/FT/QeFE4L+yW9SSvgwoyTX+vLM5QXObZWuJIKAdDiOS3G4gE4VpwvAE
p4mhwHlj8bdZPbuyJaQOTkaUQGI/BB+bP/8ed35qYMk/SZoM8GdjC8GCr4F/r4Xp
mNI8U1F9uxjQeBG6PG5OvDkwEJEB6RkN4CDokxTgegUFcjdOYo786QSGeEaAc9KX
K2VsBTpjuhBWDy0WRz57j87jW39gp3KeR6D95h9+yJ1909orPCLeWQJzhMBQuuPf
Bz4yDfCI5eFDsD3FbQX1j5WCbQCgwgF1AIl3oJDQRXfkabdcJxE92YhZ4NCQr0LC
qJXfeiZOtm9cV4iUti5O7hwF2G/81oQDTTnV77e15FVBX8rZW6zuo1502Wz3yZby
4dIjNWLu2kkgjrGyHX4BoY4+BB/5i1gbOuTHFngXU6BPCCxbPyqPbqJsUQeotIqw
xtVxRmf6AIIvzhR/L7qs47YBOnmtH3k0A3tE6b9vEdncnxKvilfDTTD6jtq3LBQd
aMVSY7zyLSWvH/QW4lo00YK1OGWftztWJgI+Oub3lgq3M6+URC+FQD23vc/o6pAU
kVNne2vJCYQl5oRbjpQIL+ZokqKr/qqmhQm2KF1+0XTEhQ7T4xTDaEoozP3s44mx
OCw7uWPiuDPsZEpxLwiOA+CUx/I3iepbJ6hW+N/84twlhJF9w4Ch6jbmjdRTY3xr
kT/BNmXRqh4zYleaZQZhXBXByOhlgqa4pN/iu2cPFAIZk2mkoLC7Ac7y01stEr2T
Z1SpglVGGxj9QklSjwP1xy2IM9eDPKf22P8lwiPqkC7CwEIEwKLj35g1LgUi3wOt
bA/Opk679G+dU+uQ/9Tqsoge+iAcdHf4QaGfpqbJ9snEBvUOy40u7PTnAvvUL86B
5lqi6Vso1ZimqXoyRjzxwMHzitG6QXGoFcYsfppLhCOzUl9E/dOn9+Nc7JbCA3uj
kqYd1pSmu+MpNd+ewfy4UUYQSAhKeRFlt//sBQW+xnYj4RJr2WZd9nTjjdWkmOe/
euIdy75rY0JR5/qRcQoUBKCGdXEleYNEJzd4WnV7ZvyhssFZWiPFQFCPH+SYTUmV
UsSc+S26LCFW2URpNITrIL0Gh2tSrRqI6ZqWYpuc8T8QDAKrth8WWx0YwZ7IAe9z
x+Woj/MbKIyY0lVlQ4M9CdgN/uYvdCyAWfjgHZssSHVz6rBDFOKKtKonZEyDJ/iG
HaRcD/tXgSUOngvzk/2PU4t11UgsOtMxYjXsoD1sza29WbaNRqw1tDoIC4KBsR50
kdIUKSxxTkCqIp3WQMHeUrRr+Wl67OM8AgN3Fc/doEQFwS97mLYhdj3mL0HZ1Jw+
7xw9yTONd1YMfYFZ8jKaAtzp0b26X76+Ct4hvPZ/aL/FyiHUlUBnVQWoA/hdds1l
BltMn1fDNT46FhUcEUu0SrTxGlUo32LFXp29AAi6SbppSWtn1dCS71kK978YIrIw
wT5AKUwSTz42dyK33fiuPlADxDvgeM+FTbBhCEmizpHzXrA7avUz5YqYKA0aw6gN
Lmp/nml2UfXByzwqO5EXB7EDenVGft0/vKMdkgf6TDbO3Aft4pNPbhrX2M/qnyu6
bpMTwO3oBeSw5BpC+WaVCukiY9BLYQk7YDtZI50Pf2LugNRQfRraH6xLivvPKOm+
zlbzt16YvVTWfDoXZxqQZFNc4ryO4wuo0RgwJ+lGM1sv37h9r2AJx/OQT1yi9mnJ
lSCeHyvj40Vsfc+7A3Ua2Wjb5V+7Ldx1GOOBT2z5jxKNUbL3sQVDAYswROt2ZO6v
Y6R07o7NWJIThF9lMU9GWHaS+dZux21HV3im+/eZC9+PycbXK8VjWf+XNm+1eYLS
hgCB6QvPigusG9L4MI+aEILhgBRbhRzaVQFI52Mn8kNJOU5TMALIAoPaL5oNzS/k
94xAYCZJ3VB/JVvVvHiC2tLRrxT8wrKFrnQUsEjzaycEQ0sFJrl6id+2Lz9Plii7
pKcpbxPgDq7Q2uRFMIqGl1xRw66+s7D8rLQVOdFFa5hUDyLVWVT+slLxD3op36k/
z0Tfk5Cy2727q97hAH+Iu6rgjn1n+CyVyk3xHbrzCWNyEqWEwG9ATPfK0zGxTOHw
1N+A0D6L9NIv+bDyvcZiu/B5gqiORKaxsD+W1OW3UumdM4kDi9k6DEIZ317eU2zv
IDthmzed2aoG9CFzCaJU0RIQTZdrDPvuln2KAsKBqU9ygDm7+/qWmI+ODdJLLeIP
xTvcjNfWdtdArOwrTDSwVfLJKmSWADwrPtO4poomt9M2s83MfJLbY7oBn3Z/0pBQ
ygBRawDVwWVbfpNztqV+9+qQvosS3GPv3/tcD2I6VBfyQ400DzSJ+4IvXfa/v9wg
eoMMXsAC93hWQk8HQIFbHuH8TohRuRl01kpv89HnSB4v4ygctaKa3khPjSbLaYBl
kVV4g3dTmG5BzWiLLJtq5Aava5GMGVM7Ox1jB79m368w8tXsj1Pl9pqW2u7aMzeT
FF7zYE8tbuvvkBXp19yBCmewd2/n5JvqUai4hpmdB8EA2tB1otS7owv/CLoWo7I0
JMu6CturlsbIPye1YDa83e6gbWwo65hK0mIfkzFh/ND8eV99oot3uL5jwE9qB3+q
9BTuJ0wmD5KdWM41velYBX2Isiv5YPW32TzWPtb+VgFJfWgxn6wbwae6Rq2juHq8
oI3oW2JrQqK8c9UIGi+f37EnfAP5z9gnvPMKNajr2oAglEzhzGO72HG/IYZqBgnb
v4/rgNaRJu+fVSI2Y0ykPyf7VXJxp+BTCtZz8a9S23l5NRWC+OyvwMYrZI+w3Esr
AnaKb9MdXtFcWSE+U0xDQ8DyYT95N41QJKl9wR9ZNTBFQJuauGywe1ykcsBreZU+
5ZWCQjpiy9KourOjhzQGmsiAaZyyWYD8yt1K4FLRa5JvkYUZ+GJ80KDxkVl0ipid
EtIsZxSXgyOSV2XElpSeJEAZ/+eYTz74O3Sbrmy/3jCzsj3w6pQtjRDg9x/Vpvim
m4FJ1fjjhSoB/I+9b8n8VZU7lBQO5d+prkuaJqCWjzO3gjCTtRGa6S7ZDqr77EdD
y++FCywVAQSwq+pWWvTesnGTJxq0lPcDfR/AZVwWvLK4Cm6eUG1UyYWP732KXSjb
I4iXoalqLY1GkaOU/0eoHETeVP9HGYMIJeB4lsJv2wbirW/FUlNDAynKq9ikPDD2
jJQ8QnIUWOvWzU9VkyN5A8Epv6Me8UgHFD0gouwF/Z5tANnXhtJ/A6Vf6oGPld8V
D4zGtBP1befurOPW5aHJqlwP8L5l3njDhgmTuyrPX5kpHGbORjluDhAdESnXbgqk
OMwkfwIxEp+iHYNABwkd+UsnsA6QpOMieRneCHYqwL6JUfB5sPOSjaq8qosXXJ8+
hQHcoh7BW+wUqxoxULcnMh6xJNE6bNvjQe3BNtNiX81b6iN9qnMYYzRgVJSiwvxH
FwbDt6DUIWDDlHyYes5YzCiUOeMtPsPRot3F29I6QWGE5PF8fykGdGSY4dRZM7zQ
ck1SvxJNTSqUW2dRfT7VIfeBZuBWqdlUyRX6lUUFeblZ12igYTkIaFzwEwyQz03m
qxgggDlFGfC+0iE1iHDVcu1JTM7MPAD1YwCcmMmKCyWH9za/WaUTjSAWA6XUbn6O
36T0a0SdlP0Xk/BZw+p0RJZe9oY3ZGYuEDmZtjYCZdKY09u/EEv0OS3ypIb1p2Lg
2WSKHI5YTmCOHmjmg03T0D5SNiV4m9PFQN83G21yZshIQvhXWVoBHMpWzrotTtFQ
FLIZ2URv0IHUP/chco9A2M2uO/W7xofFLazpMB6vLv5wwjJ0tMfxccxJPabMn4+3
2EE5F8TjJA0ZBYFhXRSWoGEmyIaP3ffqBtOgBjKIS+xa5xzwlCN3B7iSzMXq6RD8
B+CscmKEyyM+6pU+gczYC5weVgbWps+2tFXo8i3+bDwuUiNGU8I1q+26xMN+zWYy
a43BrpOP1XLy+VXFrV9EJF9Tpp7FQhgUOsHzUscFoWGoBnulJlUNz1A6CRyMnzAp
fv/mD2V3uWwFmGBQ0ZSJLv9dDWm+z2a5nofX2uDgHG3buP7to3Ngk5t9iFFJ6cNF
9pfXZtwUFRQDSVjk08RiikCuQbaIKqFrny34DRgZo+pmKBnjOS05y62LVk3cFVmz
VLlGL0TUIwOljf+Gxn77knQp3HHTUsMRcq1Fia5UtRRvdhDv5EazaM5hueV28Rkd
P1DqkTMK7H7zoFvlvZfYuhhmHFOK1xRUorqwoA/+JURXLg86hft9ncz0NHC3+cWM
4pDn1Rtyih4jPNMPwPimgufG1fB1ECJEbfbEHOniVkhWNz0ubS/YthL1jfSrEfCK
JEv9IGzovPCxliflt08C6Ri+IjOT4aPpX+n/zWl25p5PRlEMuu0Gd7f999ra9SNm
29za8wNVVyDvEJsSs3ogl7cU4PvNjTFdU/OVAEJqW2I0yGg+neX10CB57QIzyUKa
ZoBfalZLKM3iKCD6nrsfgKyCwbw3FXUsePIDJfvjSgqPcYsnHLKrIEllmkzqGv68
6h+lxF75AHN25QV7zUg53j0btGbZr+0mPQ5RAFatUB1BqGHfFT05OBEOc6EuOwy6
5PgoD5ycnv2wIIHAX25CnSWJEgOUvOIY+utDCsR384puYteFZwFz5Jgv6Bfu1niU
FhDo8MR3wzz75J2SYEuCw/VcnPGwI6Q87oEbtQHiIDscJT3DwjSOO+6jvWvRfYAF
DHcFUrQCnHf8ISss0FRtNC5b4vWJXAPpfZ2We0diS4hgHUM+lwAOqXLFIvcWw7WO
xZ8zzrQ4ywhZ+qab8qJrlUsUYsG8uYysIg+GTLTIiTarK3bbVY6qsqn0rPuVhWeR
F9qzVSmHvCco+JB73kyODjg+UZN9TDevVBMcLvdgoZ84WTR8mBympAftC3fklF+Y
sAEH/RLylYpJx61yY3l306Dl9yX+1qQ54OpLJ2NvrzcY+SQePz4OZDFNBugNjdZY
hz+zgklXEBYH/+TikLoNQ1kDRoqzAHrsDEIN75FbtAxi7rdoc08V2LACssRj6l6t
iu07Yx45t0v6TmFYbBAIMomLonwJcnXQ/WWTrRuZb65c1iVcXFoknG8yJdmry0vY
vNUZhv79p7gwvdAQFO6BZqGMaWJ+IVUredSYECozd+A/pc2tWEjzX/MLls1MkDRN
/6tiiTJIDnGPcQY5kARC0PqIcTykRWJZIz2vT4KiR+vTil8A9SJBAu9JeqN78cVp
KWlFAyF8twNv0+y5MQ/VMJ8bPHgyj6vv3sz2BWlyH9GzV8LPIuuwXyRXbKl3WWfS
EJRAhFHrdbjNTnp4V3Jl5s0j9pwKEwzJ2dICCtMf+xw9uDDxr1vGINEfEbjAB6RZ
2BCG3i76zLZiSFBDpNNBtXwWT5vX89UwjNwHaqNHSpxGB554j2383bRY6cDS9UHw
4aNFGSsUpubFCRDdkU36nPusle2InpT9Xu2xfisLa70YZ5R2F6CJ26oJGe52+B4s
t0EQdogBmpbbDXOlLlcoKg212sKDRCUtTIglAWiefbMx77xA0nmXoYMwyF8rc5Ny
Dydy0x1VCiqlbYnLeTEIhOBxtAJcqEQXJUjhaKuyPQaZevuFu/v4xcNGle8msBAH
mIrOH2oHwZB7joa9Rg2BfdmYGCA4laclKDGg/odXispAcG2CrDTot4ZruGieB/+r
TuyjmxsWzJr8qUO6fxVkJYXNB31fcMUBHomjYotKcslsm/L1/6ayHmICYRfu9g07
Q8DlPRh9/Ec+aEz4J6/DvF8uExh28dTyOMaqkUn/54oq9KEYr0DZ1ADEB3kA5N/i
xDNnrM1VDzTP6yLRwVUvVOLuwXPQBpUp96SiNyILhDCkRoE7IX7GxUHomPNUjs4l
gGS25DIFp/YmcRE1aX5j0Epj8HpNv08a0psKjd8sl4hoRY3miXtxPoMqQnuOtToC
0xFm7f40iwU7Zr9VKHXTtMAM8+h8VAQV08QGv4qDI32lSLxGQgRzyYlrVPoHqA0o
+fIB7EPLASG6lVXUh7vr/p3ZFaXcmHJrasa9cHwYZnk2DkmuIHwqpCXNgUXHfiGz
gbuL1tMIHSfBV/oaLfQtUW2GOeiG786hsqf5r/icI95nGm8WFIyaCRmzNUf/p2SH
uzKhPLuv/OnCjwGvfmmABsckj1rqftHizXhHzMXEMbfCtNGA/8HOHpOvL/sOKAGf
jgBz8zjJhxoVyXfffBRhsOM6gXQfaSc60xRoQweiPwjeNUr6VCIr07rcJb41XP/a
5wsG76iWoGClBadvnFT2Pv0JMsvhOj0XkjvHDloXRrsshbKRGaFHP3SPlP9lPCHr
WcVvNCK9YsRBLvzX9F5l8VRSZ1YlWMmppanI9XQGPwp36ri2Je5AmUcquoPbYB7j
mVwIQncBi8yn2IAs9vvfxBIv3AO09a/FaMdQJxzUbPH6r6k078IzuuqMFJuQt2fG
gI5dOtMaSG7M3EGe9Y7fQ2MLwn5g1rsQHhDsv3AuF6w2jKPJOeQge3uh65L7z2U5
jFdCLmS4kLVrtRdns5MWVgyJVBE/tHYWa+k/g0NGdSBu7RhkwQkd2ry/+mVrkAuW
IpbIuwzyy5HX33vYgYGXWe29c0oCfINqKdon7h8SrEQkCW/9FBbffKbhzw+ZOp/i
aNfhVlufm2MsIWC0lcFyctcb+Q+HwbUIPke2eaRxgGDATU+VmYQ6Tam0frpmp2Tw
/rwMaocT64tqw6o/lyT5GG4zh1wkWJfSyzAw+WHATWADjXuUMg+7F+/1q99KTLGw
porMel6e6nknK/Ws9xQOwNjnEWfvWU1f06fakApO7Y4vSH4Q2+wgi1mBIguGnrnn
6e+fjmV+wecek2+BHXY4BHvvt+0meqwxIA9x5KcizbGMBiB69nSoNss/LPwoztP5
05kqYqIMpCtSRol2U98jYbfyCAzeUyGBxleiXjLtalxLuWx5s4/tnSOjwiAYfLHY
Ji/B5ObFmBHMgux9JOrrTf99k5aX5U0GUPDF4cD6MflI+9a1S256E1fEW5PvsZgN
C/883QZ9dyl/XDTSPu8xfBRaxqJNMW26oorJSVE5ussRsjFZuxMUnnkgzMOVmAsS
2NdEXY+N1ohj/RW0pJvW99AnmRQrzVYi/gT13OPuOC8noYVxc/QjGoKECre3HxUP
cVRGMmIrtt3IYRNG8+0DPNJM5w+WfwsitSiVhZAju5WUOTwz0+l5o4z2rfNRNoPu
Is5ryR8E3CdaPLMEgiScWhBHGp8ZOAtVnqgelRvw/ex1vlXcUbFFyaG0NPKrdG/e
uXO/XYu3IcFWbK+uBm6bvsTMo3KJmRGorbM5KBXtyg15MQBEo7F5X41vMjyS2CsX
tvbLNnbXDST1YIQtUGZ0+AaGRAJi4TCHEfMaQJLy3upnQ6aO1jVVISpgT0SrjDOv
eibJElffxHcNN+xJ/wSjTz2SOnSRsm30tuA7KefkUPX4a2vbg7gdtPGoS9I2lVRU
nx16UOCRTbm+HAv5fDeP2Rs5t+byK++rnr40ISs1qIRD6SezeiHEWjty51/ixt+s
m+Ro0Br7sPlpQAjZI15DnEmezbpzCSJMnuZRDM7Grk1C+EYGo28ZXyr4W4s7Uwu+
JgzVtoHLSJcWn+v7ri6RRrASy/oHurc9oUP+3SxJN+XZ3z6RWGPUQ6fU8vOUcEJB
AEfBTa26KnbL++p+SvYjn0Esq5OeOBCw88C9gBe0QbhyEG79hS/LrYSd29ZTakEo
dNBRJJ3yCPh5BKqgufROF2zI5KaUSJhGi+4GeM85LqN7RwauUOcbN64xl5GtC9Hc
RaBazqkfvx2imn2upPR8ojMZH3C39S5L5Ci8tmtXtXZC0l3h3+M6lSKrmXmwrc/V
KgWTJjDVP0FOxrHU3rMOHd6t8x6R1tI/ynBlNOJ0baUiE/Euxiw9O37S9HtO8Jo/
jif1cW8vfEyXI9XaCgjEHVV10hRaNtvO+CPYxkerpm6ns0y8uzplsme2EX3CJ9iw
KLCc0DAYOLEbiIT/o9KDy7BXsGkCrvT6h/MERBXqxzQgRhhFDGQvhK4FvhVbX0lm
5M9GCf9UwzjwnrhQkL9eMSu03UNtjibEB9yNzy/Reu2I4CDxNRPRwQNJEa9cM0Oo
g7ZXoeuFkEw6uPnhsNm1h/t0dzYTj7u/iHF4wxyJQdlcAX+P12r58Pt2DtpFTHEx
VatOK7JcY1icM4raEYLx5s9v8tfsiUrl+LqK8/nu5Yz/WFmjhUDW/VZntPuIus46
pHW27L1MYAsqeiPzfALrg8I13XUsYjBmqQTp1PNaItfVJ2wzl3iwlrhP4lYZ9iue
0jzD7/ICShUYlVAkds3Z/g+XNaW3DwIQi9NnVVCYeixeRYKkOLiFsOT5qOJKvAUM
oGZSjP8BVrpwxBnp5+/6bv9rFmWRhhd5rxsQAc5p3YQ3dgjFv3lGWewY9i/YWglh
Uod4urxgJwa/PTfNZGTZqyUwTrWe0IzAFDgfnstuxqt4zYPl0wmYdWg8ORR4ses6
ScCU0lFmMsU3OqW+7qXpUdmTpMfGS5mZiLlS24Z4EBAYUzJfgG5Wjvipx5cr1dd8
b1MSuKx4IktJ8oecozud82FBYXSIdVENlgDdR8H5tYtpSgJuxkX09qbnOa/Nesac
h0PSi4JZsj4lVQbzbk4U7Cid1QCL0OytIQOhStz15daZt6zragYn0lvxrGfmTOdW
dmkPzPZ/im1tPCS/lVNLAL372eAD8AyMKZg6Qnbi1pY179x9g7TPg7ynwH25bmly
03LqkNR4cyG86BIL1UHgKkAwfT9AXxJ+76R22UzaMxzlh1DyDIb5UC8rNPLfumg7
CmwZ+8Ozl8Vs3xJyCQ1IQTaj2o7NFdYXHZ0SF34txyK0mjNJRH5+16YNTrYzV2N4
MtqgqoUUFLjFNB8Fwy8Lnvd7Q1cFn9fBS6URlEOPPdOS/Uayce4oOTNHQU+IDhrB
vlS5XbYobLZeRgq8vV2ChG/lLfk309ktvuEAQpHA+mxLOHpiHT3clALBxYdIk0FQ
BpS24cyA5keycza5+sVAm/y5ft+9aL7ojQhEwg9z/LK4FHfz1ql4cTljPGsQHBkY
wn7FKtcHb7TN0kRUq6kACuXbqWFCPgZnf8MkyzJhla+C63B4MANyw7w7G/gX5mOv
nG+e5qGkdlDNc4CS97G70Zg1+g1NNIrO5GLKVfMezYx6WfHzJVR4mgtaIa/G4/CY
lDyk+4R+XXq05J1ODFkH9iGGbluS5qyK5y8xm8Y7cFToN81EABEfRZ2tZF1oPVh9
NMon5RVy0kN/jpJ+fH8yVzIn490+ombhVqb1bCeLm+BdggU8uwOK5TOJ2ALebXv8
xc2WMPmm688DAQZTl0kA+4jF9bzjnDkwYT/l5pCwBuDiM2hdBC15MxEDc+iI8cZ7
Y+EF8T+G6tBuljowiuzo3YL0tCPtOXBYc5/TV+K946w5lo4YEBM1HQbfQTUhbCq+
qEz7v7Kl9agDX86gz2ELnMFFv3PE5GF2eRlpDFkbZLDogyEBdIXrQFvhgXf6hR/m
n0GijIdshgW4CP0iDs3V1V1Ji5/kv/nVcQWLh37S1yKKISNlNjaYt3I4+/+pz1b8
bp3iWCtBctIgn0avN5J8ovWSoR2WIh+XEmKjLSWU7JJP3M8i0gpC7rec3sckbteE
/6JrMsmrS9x9vz0qzNmDa9tdLOUX3pf1hxu/Yec6uxQ0x7HnhMznfUxPZphPZuKT
irY51hp4Z4TjKrBRkrLrq+4tvNwFYfOdAApAoepZ3yYqIA4rhw0EBcRBPApInqt+
ZSLeUp5oWmK2aHFMxAld3fIPHO80yCi0ERyyqf3ympo+nYu7e6qUYUj2vT0C32oL
ks6XHa3hmpN0QFJ33Js7+UyTN8AIc6Ml6Uk6JgYnGbZ/ZjSzv8H4iXS7F/YSDpkH
DWPJ8jeG9OY92cv8blPMgTiYaahHE44ND99vVx4H9nQCEYXClYjDuBiPpgbVE52o
09gAkfKQYBgRO9VXoCA0Lqv6catzqzdiSUaC1qyo7AKzVNMAW7P/Xbg/qJI/5dr+
ACxCwYO7OvHis9QVhJkxCVhUiK7AGRgm8xXCHjeS8LzG1IRMZCZlimYruOJ3ZKS7
UbFhAVsbzqs+ZaNjwWxLIlioEP+06ddzuEefR1TrgMuqd+KuXkrow1CVtiFZa3FL
IUaXqByI0+pxuRMu0dVSMB2maIWJ/BudrwmQckNj0/1RxXjB9VsG9Ly6TZP8i13U
/q3GvKNT/JqP7JRwOIebqp3sBmMZAbMPQjj2KTmSmZrdtLiPJGbVMF5UlYc7uLFo
CifhvJHyj/CPM+cw+tlXy2SC5a7PGTx1coIlIa4itU9NTReQqD9ZFDgXSVQS231b
3oYJO8+sfwkTvsLT5wrwzyVAYe+xWZFi0ZJ22KGUtmKlEOV6Py8HCSdyRSbFij60
/PfmSNsoGX0OLJccI+Xu07MEivP4qDWy87WI7pHGXYbNV5Z+Nw499hMD19Eg6w8r
Pta6Ur9Ty5aCN4IEMd5rTj+ypL7Ew04bKhT/L77njHgF7/+XAfLGoWbe5M+SxpeM
l4GOxMlqe8aB6/QT9KzmP59TESd+KaKLDr30su04xpMn3m6qS0FdtoGB6leti5x2
yUtdVwddl8VzjIxddM1chKQ43wZt9zJluzwc8TISBZXVhBX12MNFweafCSGrW2KJ
AQwCw208snFmsqNLC8za1NkBcupJUntCFGaDF+UuJtlPQ564f0fiWgF/ByS2hJQ9
A/G7Gh/QcJnbZdn9nhh8HZ5Mgbu1BnYme8+71lVU3QNiPV4Fxyem5rb6/ISptGbe
LdDouYHMJPyOSvdPhwef98/tFbZVRefCfAnyOLf6iaeY7NqkEX4NtgE6GaLt33fa
HYrW6k/gLTLbmI99707PZTeGyY+Ctf9BR+0e+NmGTA6cv3AFf9A+t5TnGDe1G49T
lnnczbjsHWGtCd14soFytjuGjyVzx+n4nPEgTRFyvcK9i9Qk/LQT1lS2OUxHlR+A
uybegIiG2Qfu7cfu5fWF4QEPRpHU31bVS/+xCLsm6Bv8OM1FWE8C1cL7txYqQti1
y1YNI3C7ZeZ7Egkg3EG3pm8RG5JOVT9GASuAZz9ArZ3wCT5+TyEUpVg8TVuuQviY
P5dX7hpVZ3UZs7hX3mhi8aMGGGhIERHBOqy3cIh3uklnb6QMlFMtZhYc1sIvjkR7
WLXuRC1d2dIRCVv6gMns9o6x9tWuP3UqRPFLIDZ3yx5/dNGJT6cuqUvPScF/tHNo
vW8pAUsXQTerE6B6cquz3y+7tdXTMALYXhw17gz2cd8lBI2D82zyxw3iNLXkJHnQ
HHqABCikWLTVaJiCIy27uwT7z9T0MDWMzhlqk7xYJ3LmFZzbKagdbxmAQXokRFgJ
9NjbjruELh1Rwgb7s02LokKg8glSFlnnrirPBghNb7vYWJmvujopcxe37tfRMowo
p5qh3Kzu4y3MrLbMomfm3a2PsgYCt/ZHelxdOs5Hd+rv+j9cG0FgMZfAYzL8qhV5
8iaknTCdaytlO1fr25VhUHNb7yP9AMoxy8sQy7aPz8tcACJHf1Krc2B5VD5TD/yG
ILr9BYAXc+MGsEb91Jh053oQ8K7vbHNU1O//dMG47GRusK2cwfSkufYv7I93Bb2F
V2pNN1Q1x10dLWWHBk952b2IwhIlMa+zKBxV5oaoAah9Nv0JHwvMh8UHxlJKWZZw
nuU2yG7MyhTxISsnOyHapPrJKZUIRUccEGvP+lTnOe9jRtHcpRv8Z2fID7TDg6J6
4fGDtvUbK7M7b0YND5jyWJKXThP0aRD+k/HQv5seRBjxGOhygeZwhIgTanpA4u9y
cA0OBHSSmdVI1AnxWH4R1RJYSkI3pufWz2b+TjIz8pNqCX/UZL5vbYt5FDfY94jo
ioaUB4Oqe1T8M93gORknhvnovpn2Eah2fl7+M4YQqoTm7gagI7CS0QAEya6enoty
NhbWgBU5w2hKABDGlRSk7IYuvoKKdVhKLrGI2NebcvaRs7eyLAaGo2xE61bUH3ki
xPfs+chRw7yF1kDL7gp16Z1b1JCuKNB2MR92sGhH+9IjGNhhcuQpyzW7dWQcZ5kl
hlHPJ10bGIROtDfPtmBfHL8wyMCxZ8V86TfH9LlFlGMJ+vSd4V1KBZWoxm7+WKrG
wtiYXtX6vf61qa4o6cas2PmlBhSRHXvd5tLLTdVx3zbuYBMDSfbvsJvmMxWu4fra
BlIj6smAdTKlnS87nIwjN410G9Xru1boNF9TSO7j6y6aQYdd5hAbHsdMTsuskaOW
GHw09L7ops3uxRmkXh9duZael4mrsSeRcTN3gXKPqNm0IFVVztu1cpqdjChw+4KB
x1TC88fELvhTQ77wkHhkqdZYZDjlb7n+VFx+rIiw8qSk/ldvQPrmvl2hrF+Pt1Iw
CTtCH27Bv0C+tKJOSduKkYjdafUgWQzc9Pk3+DOu5oQSjtL8eFzx9dOokrw5R/a6
J3Sb/6gAiMixHnbLdwFRfKCwGAlhOEVfr+FQBQrNdW12FNlcHs32rgCgIbuK/pJF
Bjc9g0jejpEhlBmXwUt7lCrURS4QXJZM7Bl2E9pcOW52FmFqJ8Yhm77HP4Qq9RLR
SkMQmB2obcOv2rxqrZSSh+7PdG1dOr6ELXf8Nb1wGltDbKdYbJj9hA+1JbXzh0WX
4mhnprR8IlmvJi9VnpLmgA8oavdQusJQeUFhNoSe4Y+LlF3kYqGeHzLov1uwjswL
Xivt+3PMVg4uEANUpFjaaf8JqXt0ZjUMo02c+GhvKNf/NWrkJiNWMUy/LYdSWq/K
8crRZy6hT5fdAWQhlVIJge4tyx7i0oqSrT8Mn83F2Np7U6H4QpK3P8wxNBvzPIa/
xqtSDpYdgK4BgReXVzj76+WRr70bhRFahsIpKNZ70umNjcHI6JsCsWukQXW7Wzvt
d7cxsPsnzz1RU9sj77lelbg0fpd0KfX8Rr0XCytPYp/BqgFmOI/VndaPAXRSAhOn
lV5B6tj7cU8XferTezpVm50b+lqFTy0ZVVteTiJTsl7082UM9ovoiU3In1wR16ay
X6SGtc25GnZg6UH3ToYOjoY4JqIOtlQyVpKpfjujrwBrznMLHcP2VoZFh0aaakNA
zaL13NucN7Kskj/M6PggVllbshTZ+/rVSIquEUi1/X8yHoWCOnwQNIi4G8Gfs0iU
QIe6LxNguhKcpr66Z0lg7KiP/3TAG3k56EJ6YHbd8Ph2PiyN4lhX/iqMcstyczdJ
kHHhjuzMoNxE/TQAsiv6O95ZOYyC751fxPw6AqtuqSbeATCmXphaWEyEHbPzGG4/
w38nQorl9sYgL5BN2e565fWQ6JVFx3Q/DSLpGk4xqffW+nQt0gRunx0qWfF9pUSg
kPT/FiqUjTJpzI8doDbu423hFWmYDAqQukID+FVScO1H0NrhWXGZ+NAaCTe5iRSp
R/5pZljsnG4lfFpbR9NtheqLKLAH9D9Kxs85XsMQp+a5VwieY6fZs88eQYSg1lMh
puZH2uIOrWhNsvKykmED4X7vMmMggiDl1uPBuxA1xKQvSaAkVPe5vCwGYO84JkPP
CrRqbl14bHxUGe6539nmMyKimJw0EnHdMIyyhW+mD5UOZFREMVWoBlqbt+/bA9B7
vYrnuptMhw5xHmFTwb4uPCMIy3hr2dbFrsqc3eAHZndsNluC0X53qXQaZekz+ubA
LxmzmIBb0FHueu21Yj2gcAGN1YzdnMtIyce8g8PNGl4xxQnLo04dC8rqhzU0/sSI
jggiDRRnl1erKHylAq1/5BnIldSvcIPh1ZN9bRHIbG2lkW4ZiNX7cuGld534j8HW
ncn7ARVp2LH3cvwaTo3HrjzjZ1nhJ5iOaGJrhojHeh1t8p5V/fMYaoPAaEk2VmB5
BgXTrHh6Nc+NSFRofq6NTOUCKLQTcMWFY9hOqnyTKwrG5J5weG6LvZloXbi+DaSI
LiZdH0jT5JRlzdqb0vQyY5TfgYDibsNo5IjZUD5Y2thJoq2H+c/KxqaokSr/HQi/
9XL4IU+VWzOg1yuGzL1X285H3NrS5gyDioe/Hn2lLluJFsD3NLNppB+B/RO1cg5p
en46/NGOYGbg4UQhS4cHCkKmvSXKVg05O6FrLK0wZ6/e4CPWWfOYywF2nrlpaFIX
cp4Wgvet+eGiE3JtcyMQ9BVrSQVKMxewlfKoJiXhjRLIiNCs16DEcYW9de2uAvKG
u1MBxFSx06AQ2mizSa3QOo+sNU++9IM2UCLPiNFmsgbQ7U+G1CzvDc7p70TEluTo
K71c0x/46Bh0s8eu8mnCxBRAEJxshm2L3AZVAGm8ejTWId2I5AKBKz1W1ciR2iSR
91QpCej52I1eLBzNF8QFwOtF8XMtuaqIhcy7lTYE2JScM5aO3OCfwKaI8NfjPlIZ
6zvhw1iI8RwG75RoEw7J0lFNohvlNekZQnUp9qitDkBkWtmM8IWw4o1EGmxAK8f7
0GDvI6brMrVMp7S3qIFS/RPthK06pVkOTtP7cF+fXv/6rAVCn8b1ETc/jzf4a7NU
n6zY5jnreZQntnfqzNVzIXn81myaE6S/iWql+FsHYT/x1F0lnrcGQVKKtwkW8xr4
06NCEMlpy8XF6geZxCkV4lL+zUWSDcoQbEn52qu5ODInqHkklllVL8bZ1SoXl4sX
opk02tzMt0LOw/eN28zUroIUmFkp5UI9iE03E/07etxEUMlZIxl9H97DHwBuIMx7
egiIjinVTph4/J4eC1uvR1cOSbGMctLKtN/fTG4wWSOue3gT4in3B8B/4SJSFrYS
QhL4VJIgTC6vRlBFruH6DkzsNzHdIwJbNykRDBySw2udSafmM7qiH28LraYvzVcD
R7gPCAGgbyOjPmqvy/0PARR1mAwQADIo2tdJc0ihm4Zwq3FEhDfYTNEphMtIfC4L
BBXqO9pAiqgFDGf6R9ZjYUbR4/yvoWe/eC3prZHMQ6ULJO0nmGbK0DPUvEPtMxqs
jCmU1o50+izkcgvvIEUpk2GpyqGzMlkz/mh5+VnJnVBV14g/l2bph8fwbwiOet5Q
Kz2WnTewhxhE0uIEPHaMQSv1xC+VM+tzLVr5YyrNxetnjOhDCPlGsWVk6woiDa/R
6jhQYtu6YlIiphj91qRSTEuBTgtgrSMLFYzGVpftA0cpw8ZB054+yHYxnWiiujrr
hJJyiQcLY/cY8GtqU1ID0iREehY/Kn17G1YeGdi7SYvf2cHYxnU0vE4TGivzYmPJ
HXiGTpLTxw9E5VoTQwtpvJAZY7IYviRYFVT0rU+tO6PeV04iynxVy3jTeWDSQow0
bRN0ZmbDLiurIRpoyorTCbVXqRAQ8rKM1uTRRibQrJ/kpe/ot6f4nR+gGUlq+sgT
Z3kU3pg0611/iCSkikqWQYZuTYmY2t3OZSkl6psnWx1q0lgLTd47/znTUYCSzJkS
a4UriCrPx2dLskL01jDdwWMEda6fi9tcbBj9ZzDKlAIpqe450YjUxkpa+QzU/myW
Rz3EAZHdO4CSn13J4wzHO0DVZKpnE2M55hW/F/CRsyqye1JVGTTLE4Yr0fNaKaOO
pk257HahSK4YhO4aLe0alYP+wNk49xzQA6SJQuTqiJB9g/pkPZ7G5XKUxWS3PNg2
0e/d0jxIu4COielGyqVqJ6MN0DoYh62VT5hXC37400A/pYTdUGtVXY30Yrn2otKk
l3BsR2snGitP10W/jeEw+NWsMlxJ18JCVtfAmLwE9OYALUzJ0Nuq6wQC57skrqcc
7XPAZCs5C8NgavqYemmvOCws1+JOH9QsYs1siPwcr0tzpA5XozYlUF0TV/zhZZXb
sKp1zJlIlLWtdorlTOrS1KjluxzeROdbedsg9kMeYtTFM2r31kRrY5VGqrnX1BHW
45tW9tVUkRwp5oLbGIiCCwE37tH6XlvZPSJmplSwNjgaJm2VMdZ4jM70ovfY+QAU
DkTgnAkdq5cPWdMgo4IublORXvlQujHPjl/xFSykQ0pUHB8y9X9isV4Sq8d32aA8
DjjYhqzqGSP8dxD7jxSoJ6N49DCR2IGS+/qUT0cpn4zsVXWG5l9fdjfxA7QvDLQG
yDCjr61lQ/SoDSeXL1rgj5WQe08HvoVF4uZaZhzq643Nfl+J0BtQajabkniUl/pE
SBl2L0WszfSW+hN48KZ9uXAWlYNuk+faQihMrTMdrFO6uXN0DRZFikvEolY36w4N
i3Gn8RLLxL9bFJWRaWtwKGLuhGST2qozKUkqL9zcKTYdgvq3DMovY3CmhqobyCwi
mM1311z+sNjQPysYzG1DTDoToC0YdkHYiAQ1OkEKcVnuFw3ClXPA0uFOvIWE6A9D
RhDnCCfj5pBQZ8luZrnIAcS37wMkOyt0tF+B9rlrAZIJXkSemYNJ1TAvQi2D+vG0
38+wS7OrQh+D+LaU/R9HIP/kwq0LE/hCbs7A7aE4YadNkZZd+Wc6XoRzhnEbtfQm
2Ah/LqhLco8FVNdcKc+EPAhN+ZhDRnMzAgsPG0DIQyMJgY/K5DzHjE06Puhd+2xh
IdE0TXAVdS0KP2TKkfznRs2SiX8dvSPw9lHQV/36C94miv4YN4vt9WlQjOk8ac1M
x/HprH0kSdPy/tRMiiLEfvEQNbPxaWDBl0gWDQGKkyvgBlE2ISfepbnJP3F9U/we
HWTfHo5s21asqkJ2UjxTK46RRflN1/2WgOhDnMk3Yyll1Zwgl/S/UH50BCSiZgAN
l4DQ1mIp5UcXkXcAYDQf2fTxjDpW6bKAijTP/Vx/rRhX2/d+BztDvmlDS/ANAjQd
Hj2xsiVpqDevbFRTjtMBEY8HJ0/x6LVtlU4G4gIXImTWS5c0LXzLzniA8G9KNIq9
oKAFx2ILHoz8Boe5SUye2jhVWx5g2c0sGjjartkEJlIQkDvdNHY/93AC+vtGfevL
n2AYonADZ8mDQRgnFmSyU/nIlrebGMX2y5l10l5moQhB+H4YtaTuoHKrzIxK5kyx
P2TeXn0QREKNVAwtQSSqzKR1KG/9uPqujR4Da4WmPxdiGqPHFIV5KnAo4ZAbCgj+
40Ko7TZg5oFeOMA0lNdxRl6oR+8usk0RuWRYf8689Xub8O3u9+lMKDpCUMONdCOF
JBj0AjkgRCMuY65CedeNvfKxJG49Jlgn1QzwU5UOxgP+g7b+ab6XNrEzcMki4gUC
gPfxNeCrPgAJQwcfS3zSlg0Wswg3G24T089406d9UOj3Zv7N59/F06wTBLwZwkW8
rRT68Q5Ft4u9BljIF50vgNd1EO6uKNNAKeOWJQ/I0tud6/D9V2Vw7uvdsH1GJrwd
xHmlM0vT1ZBusCfL1mMGm/1SfLttYF2Sdn7hJiHyryIrYVKnwHytWMjILitmY9bX
2DOx7F5AQ/vr2rN2XBAbb0u0i1/vkSKqj9H380aJES9ylhkTiXkP1aVActL/+dsU
ioKDEzr8W1L9Q90aA3qVhUJ6wOJaOdChh/w+G2sR3m9LiDa4rP2hyRU+s8kDu9C9
sJbvcTj14K/Uv3V38w6F0TAZ+7vz09L3cg7WOh9BEET3qvElQRV3g4EpJA279vK1
Lrm493Jripy3vxSVWNXD9o3fj1vBZlCE+L6mulYkTpGvF5pf7a/fHJrxvXU9TZOg
5iGUVzpK3J+0ET9W9BqrMK2FU/FEUupAKmBPuvUSbJBvXtJYiGtL0GST3VikCwm/
y8RAYQZfGtxtxTQRiZ3SeJ7fqMrkY6r+yKByyNSmoTn1oyxQGgpqGn3UZJxb59Ie
7aAGXK6MG+JkF1h4ixMjh/GfYHBlcbaQctaH7DGUr/QOFCR1fxwZxTg8fLXmLlSg
aRaCezBOwOMPUGnhd73JCA4zgB+msa48MiUFqPV8GlU9B4+RLl8QbEymZbmjDYjy
78x+xfC1no2CsNJ4djjsy2DjihIQ88KbWGtS0unSr+0b6RUVZo05PJaTqP9gcOYX
k595ufZfNfBVaEdP/QfJfZ/e4KATfTGYV+5jDD0mRr0Ef5Qv1toBoFFRpuQr3b5g
AOC3YWZ2YYEjmpgg8uO46icnyyO8eea47thQV0FtGg7rRMmoQ7DPiHVIbjiy7NHT
b9mTEMFGKWPKqaA9IDlWfvIkirr6w1eNWWGFWCpPgLkycQLrWGBtGEbqncKeDzB9
QGWuIk21kSVcIASJDXcr7mx/cmL4iWtIV5febPLXXya2aoVKJMTWZI37fn5Xrohp
B2phd1QEXiCtZd4tr5XM9EE9o/52XlkT8/FtWM7yBhv1XKdyzhCZAPl1l8JfEHch
n1lCnfWwIgIK+CuN2deBUJxQAdEhOwkcDP3GEJaQnfla+yKW0ZwP9PqYNw/DGu/C
qRpxKDHqnf8TVd2pPAgeiHkPZvUmDXDbFz6gtoJ2kZXjvUYBpLY2y3BnwNOf5e08
qId8aNujjmpGGjtUELHpTlOnfP6+LONJjcnCTe5au8jEOndnMaZCChHfaNxuFds+
rpbNZxKEghXbQxC/1gjANxnxw8b7MA8ZzhRnNL3XmKRFKsdNbwJxwmCu5rTi80dN
758oHedvRTPeyTpH+vSKBEQmt9Mu1Kdfna5j3F7lvGhfIUDFLLqh9I+Dz9yB6YSV
0LyLh6QxMRFQr1HGupFCB8q+0d1TiyGnQQKNPHzQcEeb4W4O/o/s+dFbNsrUIT+L
Frp8p/7h8z0HhSXQ5txhlVirtknCemkHsortyWL9sZ9mliBQ2NIcHOforA8/FBv0
wb9IadYsv6+ha0gbGLwMMMarNmKzN1vWuyErrNi2XP37aRkUtu+GMMXN9LyNp/4n
AbKyPYNvDDy5SAm6OdgrRK2auzW+JoXtREWh6ccKHXxupKjB/Tjv08Xd5TZqehWj
Ypd/KIYLlRzXG9sYjMxgRFybgSxa7xELlBLbGvQ2cSPTGr7usfuRIz9DXEZQmBnN
HlRlyA8xTBxV39yNU26UNRyA1clblNYRZ6qeVkRoi5F5LqQhKdrUV3tnRBnSySnE
g6Cj1/bNaWYdx2N2Z+NS4985yjpinR8FOtYBQs8SHbV0tZvAzaiWNDla05lGjMO5
SLOOiW2ajhpZ8oPKN+d08XB2nGTo46+kEvDK1OJn3IosPeL/H+wUu+dPjpKs1yE+
Qt1Omk2/Gt5ofLzfeChimwouC84kbFyy3QCTGIIATlZIZegVuWxh9xV6JEc3p2HE
Gg2FSh8hUp3tjr+qpQSBDXH60Hf5/u3chHYhvnhR3UxELl0z2gMmCoWryDAMqX4Z
LoUGyQ5H/RMbkmdx1fd570sRGmTurXcS1cvy5p1FKHglGYP9BBqix2trLKm8gdLr
Z4Uw1p4bzab4U+orZGjDMlAnUzGjmqjzY/aomPmdjfMqqVRQLJpPN31YOyb7Y/3k
hwOthpcceiqEuOqt0JqTuMWxMDwuef6kpI5K0odXRhoHRBMlfuuaj3pOYlzLzBri
YNIgbrJuJ0DGb+StCGXQElNk4S1eGhNef8Y4Hi6L+WhtkhHss+Sbf69PwBotd0Wn
QVj2ou5mzclCV1yDjXYdxEU1oxz/Oh8/55E2i9e7Ty6mv1whikmiCdXrQ5e+wtRl
vIKbUFpjLCslDUPY209Qh/qVWtyj1LYMLnkq3LUYz2BsiU0KWvwx9jcpnGl8CD2w
JrF+CUhqIrrclMoE1a7OTTKhIgTxWyjqhK2qaodY5ljMZcrzreMzEb+ha0hKQPlx
62IdQal/hhrnD7My9mimZRcjfBECCpsQdtgKjfP5CXnydtqhforK7SmsfPeX/se7
K/VyF/uHGVreKiiQqW5VSYe38Lo1KNXCEQ5IN42dcA73M60rrLQgCbYXgTxaG4AV
s7Zb03ERDU29Qii3yoKcnof9YvzFctOdhsN6pSErqZB2rOZ6OTlD5WjaFhLqzCtL
IU/z8eID+rTIZPOoxXrX7Z0f91j83pHB1uMoaRFcJk7js2LhZQ4zzqW0+VYsLyM5
wNUy+NfCJXBaaFUx/3+BL2h+EaBh8bz4IHDh4AWEKZ+9YrNaBlxvumu96n6Vo8AJ
VrsGwZvyUPljU1mAUSgs0OIAazOH62N3svGqp56Q77WgX6CzC6J6U2EPZgcRPeA5
cknpbIvumrpDReeGT0Okbc54RQR6wHU1zxi4oHQz/i5uNa6RtNDVdtST1i04jBhu
eFRmSl341ss6Z3cmK/hoCAe4Tre277XqGHzVMi7Z4xcpVXD4EFZr6yWKHW62pPQe
NopHw1VOCIcwz526wIg+Yzg0RwraBIZKE8YTrvKR0AYee2dw2PEcfR7VsvHrGbxg
cvFFLqmDmxPodl8xfEBR3lIsYyu4VbkTCqR9O2aG2tvDfdjp7MUIc2skJVihpZm7
eARw+vbR61jxdWkZCNbXdThumcfYVx0XVHiwrZGrFU+32dASL0c3gMrIe13lIKhQ
CSMWHEkI2wKIA0BOGFyQh0fdK2sxgN8EYAozW6hxvTYfO5ao8rrROUpez5qiKFyX
NSUfLqe4H4R1uYXHynT4g9pzekT09OsCFNFyhKDWOPrg/r1ZMWKDnnx0jt5FBogy
eGBLN93oDln8ZkczV4N8wi8HWoYjY7+wUglF0XzIIdyIv0+U71GOekU5ZACU/q8d
nRAhBBwcwoZMXVwAlNEBA3pz6E27mWORzonDCW9eZJa9FfjnUlSyVLQWNWp2hocr
crdqbALw8HMHjQ3zHmGEH1PaOS2r//c9zSnxTz/kuJNDaCJ49lbT7yW44veMrE71
uIx1xzWZbM+zVeKAFgYIJdmFCNEdNNAwfdWx7Cwx5l0NYmEo5jq+GPmVzFtgyHUX
3v9bBud55LQjG80vBKa8aFw2B4cJdMMllt/j5CyjB1xnhcFbOBfQLCySfDnNJRO7
t4m6H/sOV8bhlWlMvSwktSkx6Zgl24cBCrgvnRswhwh0f/JXekw0qdAxdIwhqOQs
LWI/FdbP1ka0j/0rjja4P/8TQWZiIq8zehA6sOjZepdGOzuE7PwO5AdKqIiMoMW0
DN24ZqqCUTmaELHV3cK06mlsJemUE6nxoEkEqJ79GIzZevM9oMTHvlW374QTYTrp
Yz1KgLC3OqLSreTztP3YptaohPkxWbQAs0+5lgFGISQrHoUotGXMniEAns9ECjnE
73ubTJQ4Rsqp6VNyt1aB7uUdVu5ssonNgtxg3dUhymPSHV30cDvProo4EP3kvHQE
+Eg9cOKT+5/GTSOluxNiRvQXYa89VlSB5UcUNt4LfbTwPhlRRCKjW+JOK7mcKneE
C+ZK6EZjq3nrVTJ1P2YzNeOqt102GxVAZ5zzXUEnMq21fUdGGW65g3t2b1CMXXp2
+H5nx3ssWcs3k6juQ9k3+AlRLS2GjLqQnpQgDdWDX/Gy7UMfQn9VdHUaMcLvo9tL
T+h0L90wHs3h/uG5eqGAffU/1/pnBIY6jGD/qeWNTLCQ/1KEx4dFL7VDeppQyV4v
HVTbHpd3H8UBXjyTfqJ76rkxfpUcqnxf+Sr4bEFGuD+rrFV2SgXJaVy2AADOgIsU
tk8YGTIO79+WoT1GRNOr9JzDVvtk8uaIBDSPxWxP4p9yfRoBX8xxVWJlhVsc506f
LLjifa2+Dg2FCVkOjCsT0JSlAoFCO22pn9AYCrVAWtSCv9Amxe30kWiqRRuawtzK
LcDYKYtsm1YCN67YlEiKterf2kwa5vhQTqv9lOZXdN5yaC/HKexC3RqMtIqNXaSJ
LbzUApC+cl660NoEzpx7MeRvXO9TfSN/gm76VG63kTAXdJF2UR5Tn+OgHYI8f/uI
PDtWXarhvwEc09PYQDTgTkgrLg6tSRCWeTHZbWsnUXdGsRuUjNRWgw+wfClboQEm
6+0OndAeJPCdVctEtzNwwYYl3wO1cWdClo366fYNRdr9lECsPwuWSbR2ZuxrbVnj
xwe73jO3sdiXYwIU/y+qUh2erir9/+1tx2MBqGxdmmhrRnGII8CczyyadAn0OVL2
z5GGAlJ0kilfeZcJvb2rFFQGVQxSdbAgHZGWlGNM1Ogmux17CMRyvKyKsvQiPSQo
4QGGvShUJuEN/VyY/y1mjCi3oCLEas/aK8k2CZlbvOJzaVADLh2QR2d6tRIZhSjf
RFaoyKB345R+nY4wDGunXwBk4pMbZ4fP24ClTRwsGWD4OR0QQSZn8yEoT5RovHTI
X2eLrlLN49lDUT1Mr6uL4SIZ581gExINkSrE8mEA8jRb8CiBqdVn9BNpEit6eM20
bPyLb9fIkxLZ6F+Ory+6nG0ni01LzAhNI1cL3RQezRxHuPzHWoi/GuqIdzLujkk8
YGFi+Pyj3Z4jrMewMX40u1rK9Zvj+68k/vLu09RStRVu3D3PR8Ycid8Y2cocu+hh
vP2qkFH4zklmBwaS9Q8Xn/v+tEomsdkW3kZZwFDiU5Gb0Fpn5QssAzn3Nqtu7Npj
tj7rNA2dlktF/6JTy6EuecjwFpR0ZTQgID/nwZVEo1leIeW8JTDhkv4kR6zYDY1l
qE/DAeVr2WVPIVn93ZDvN/jLmoaE2tkVcauuhKPFFuR9lEJmbuc7KdFWqsLAJ+uX
/idOzBILOAYpBFmZ3llrTDcwAD8ZRreSZy0Cu/n8trmWZBgzy5tNX69Ja4DscMUD
QZ+u8u7mVAwusUIYRFjUbP9CrhzhcGqyjFuurTB56WpPvHLnCz1lIrdw/FU4ZTsg
u0van8bZv90FQtw/z/klXQ16q2u25BgzTEMoVh//BslYCGK6FfF0/xFVf7o1CAoW
gSiny3y0s8V06q5R6GoBw75ufPYQTXgj7isCqnVfnM/NeC+sZF+K9j8s3+yqm9X5
MYLuy0QHbIErpoTPsDkDuKse32rzkytY19btiq97PaHhczdPQlpa+RF83GLRXFtK
REeSyIGAcKpkpTuqhVAHJ+BAJv9k8BY35F5knDvI8lQpbNkjzPoLynj80eDd1x3r
5p7H7D6qQveEaWUpd9pFJ2h0kCS8GKxHQ8aPHL1wEthjSpgCGBAGObwlDNtVIm5u
cPU1wdlaXojA5qFYhowRTWnNE0Vp/NiAjQRnD884TpSNikNnUy8BaUCSvBSL5P02
pb74jUX8Lm8Gki8Zg0mNNXYTqxWuW7gdbzvUSbJGCV0r6eFgP4fcA+TivD+wwxri
Jcb3LDoAEbO4NA9WyGbw/OWcdiKFGpp7ZwRWgJfJLsZILVmr+dkL2x4yrVlyoLMe
I7Gty3/pqHn0w0T4I0kTw+9fwvpUjLhwL7qjNZwOy+HUQLjR4M/769GswwSdPILW
mDth/Ko1ICAsVtL6zOLagv8gBp1DN13uwLejad7dWgCzTw4I51CyHPM5YZp3Bwle
6P/VKeURhd52Zv1B4I+bnRcSrKIHQzUgSDZPTbN5a3GQm1bQMy3cRCUdW+0/rzOP
ypVKR0fF5LVA6bJwQfLySrv19xhmvuvMFhy7HtoovkjUUuqlapxdNKxBW+KfYlGd
v4oIexmVcH2woKxXZzWcpHeBuZ/ReOlNa09KEqKISZjM+/zfXLucdkvCgkHl2/3y
Jif1Ex5oonVyTlCLCAwrgx9rP9DuyNVBuvqWwQ4+txQBvYNfz+/yk1eKcoEwh2HR
PrQV0I9lQoukzUhX0l3SIYbRAGfk/aRmBTZlo2DRR2MYJfKHP+hKOyw3WMci78BN
F39k4f7cnYNSiWNjX5zL1nj+mY+a35fwZcBh2sDJejm3qZ+fCuVNvAUbYIr6nRB/
fPTM1gc/q+35ED42xOo9qWPtJKvfT7Rue3YuVqEtp5xjkmaSR9dDs0w4ci5qt4G/
ralKR6FWJoVCurf3ZnshF45XaD8aoFdTkLF+ev39/hl+WVoGuc8kEDZglfSqG2Kg
kcE47luepRpII2h9qf/8+377D5/y0owwnTWi+NdZ3ecrUZ4TN5NHq6FrkJYGAybZ
GjdaUG9p1BAFsmHw8sVB+8VowI+4LPmGMpey6OU7QMdqL7SOTP6vYqsntbeMh5o1
tR1wtVOlw8j5AXD3y7iCThLJ1jPSoLkD/byblRWFo8AN+NNUFPhCYlyiWOhE4i0/
FqFkQAsqy3Fk0h4D5Qouyl+VNoWB2sSBd+impdRPWQPAYDUwGfMrpP1javWTAUoa
0X1bDQOaB0Wj81oXgOf7FUaGfq4SxQ0eAinFxZGN9RKhXvP2c8hSAaHfBnOhou/Q
JkNJW489kyXf0/aUaHnWDFYOIj8p1fjikGV0VaiwkC89lm9v2YyFQpjmwVtwZ5Q0
ICeSQOtJwhHiloNsMhuH/AW95+bNnYu+JVj76x5A+xjofKWbw2N+tfHlryW6W9xR
PuehGLMYJzeRSfDmYoQZxFhtryj9uhiZlaxjebmmkkQBE5utkI6TXfghPNLXrume
91g8qq2Z+eBK0RueMKDm90+gk5ul/W+/f5mpUq6DfyUfwOZ5Go0fKPg8En5+54aE
MpoNAtu0xyU5LGJmZL2Aw22xB/543EgtPL32T10u0gbbpfRbHWvnxbLLcgB7cMG9
x2Ig1hzn7DpUNwQncBvJlhuVBL2dANeMh9RsBgmJNgRroQHbAV3A5fdcv+KvCzfw
8Fyhbkcjsc//1a5MGCPL1QHz+aqdfZKxFGanIhoGzjZV9n8/4tTPiPGUiidqTeHg
ZdUtGscEf+wXr6kOGQJcIPbkdQTTgMNybuYgWOxeTuq/8BSChhFMBMncVOjYhm/W
NniShR6puVQngrdoDNoDWHjQVFlYtrp4IlOK7jjqGtrYikQtD3Yh9t55TMfe+Cnw
4rJOKMiS/QifUab+z8vPO0d1TQuTRvNfTAGEbB/InCVnEoQ9ipzeR0/bctLVBSQH
bUalSpMCS79NHIT/ZggJ0ZWW75uHtUMvHrjUTYyhYK/+Z54EfiAme6ZF6wG0WArg
F6Kdvj+LKf+TjIoeZic7tuzdmzdXoWuhTOXcdKz70EPH54GIDqQqnrtQfwDXZuWT
I/2I3bFzLNCIK+H2MRoueBS/eUzQzhmhu8yJ8AF9nJcxvh1see0MPOfsSDwUOrUq
3zde5balMwpQkIUi3JFF48xoNZHKcnsBZlmg0f2Na64gi0orn8UGaHLsSm8W7g3v
nlL3cKNHj0C0WOjs9O2cHr5aGzJ4onnjmXe4emIfNfbEMXCbafQYl5TsDRfUZDvF
wWXUlyKdoxQ/uy0WeSdATiPgoP9lkwW0lBPoZ5bY4+ZjB9h7eMzWr+gBBLUpOoJQ
nXc+JRPLKCE05Xdhnwp+kSEnohH2iSigVEQUWmV+pAPiTxtMFsOKC3v0d75w3nfS
8vAAF1VZvuRz0J4v2pF+sk94/Z2SowPwqieMmWV0COyITgE4NQE01Mp+UPWeaFTn
ZBZGpgpgSz2zyrMB4OUooxxVK4fcZ09Fkwn/zzq/AXLPnDdNDUbnY2iSPqgef2Nj
0NrDYTqAqLGUHDpKIbe3LrS1kj055nAjpzSb/U8MrqsQoyDmb59HDs7SJtcE1JBR
rsiMkLlmTRhneCgMxxlweGEpc/WQaMXbI27ARdIpqQovHC3BSM+EVPWitN0oQ9/C
zMvZmOCtKgoO098nrvyh21I56Hz0rjT84OC8QPZELeJwOcUdQDoAe16VxFrxk0Sz
1Fh0j5zA/+REqukw1M0XhxSNgMb6PaE23QL3bxzy6oFYwE878ibBRF47KEUcBpah
vu7Ql4NVTRCO+XgxhGnpEGVr8zAUaKZE+yBPIXeZ0Pbg1dJF5dlyGH9PnvQBautj
l+Vv/vqv2diHNwYsyFIgK1bxd89R1q3KMhRJ+29ta7yc0/cN0dbHZq2uMl81ikXB
SIxZfqISKUfCre1x43u0UKijs2DY1gxKlmUr718jt6WGOJPxQCZRFXHDbz0hzzrs
F4wxR9BVU/X8rvKl7B8LMnd9/kUW0E0POw6tXPUAqVxcJqAJwShHTOEYeWo0ek66
R1ZMxB8mQqh3ZZcUw8XvRF5qBT2Dy3lhoaD5IujICNAXBpKf6If+2+XTYSgpek8R
Z9BcKoLUisGl3ZfxCGvUtMsvsPduhNchKPyiLSI7NCTWXTv9+9mdhfXV/NvkcgK/
v9ed0qfHDbl9s7ZE54vJ4ga6PaU5D9q8oOIpGTebupMsRJZgSLK5XpLlK23MdZut
tVu4Kh2tAXqAGw/CgX5SArgDKI+4DeKfq+17ZvQ0mlltdzXg+0ne080KU/qKg/ZM
mdFckVCZc8Mdf7Qz5Nn2px9k08CBvDGLue+8dwT6GhMJcmiVoLJj5MDGxqvjL3sD
UdvcxdtwW5wUHqdIOC+oaGvl2R+5vgVoreZTIB4h8cHnomi/owdI3wmiCMpVpRF9
NqGgT3QOHc/8SqNQZkquR5AixPWcok61bZ0AcNBgAoR9c27aIfy7VztXsJuBeUfy
vSTGS51FND3L6Re6SO/tgBZmNd0ac9bpE8RWY2t6KWEelXOKgaZ7JOXo1Slnw+3p
1iUbdi6SNBkxwppr2JynZdHaMKOf/4rSB1ml10A6/UC0d+zYtE1tFExtf7OAWsXw
WCp6K/YYc3AychtjEexwj6oIZrH+psw+azhk/iv7hQu5A8hvS3TsvfH0zEdwzd3e
SmcaTH1GGwL9KbwZ9YWo+d/77Z7v2JK/CK4vxx1SqLIQLyFIcJtLdjRA1QpR7GO7
Fl6PFyKCA3la8bd0t2c/AkkHsjmmo+zu9m23UyEbQvY9/n/IQrSV8FYnExFuVDj/
HgbysVSmCxq7p7RgHqOXw34pdmUog/jp88fwSvQnfuYv7DkXVR1CIfAAMkGA5x03
acwF9P6bqgVvKOt5faJD/S8rbfZhMf71Q+7bpoy5ATGwWczwZO828Zym6O8VGR5a
8sNjioHosZWTB4mavJPJ3jy7v+7N5ZuwQh00BrA2/tWmmrOfNRpZyq9oR6S08rGu
Voywx6wE9HXIg+Js6b5/ayaphYwE+njmgBgGD6wkog7q/ft7UEM3b3t9P2PTgQNn
dgwi8qhstE9Kvbb5jKSInrhuyGivKbp0S+gObLl5AGm3KhZDO/nYVDw72ZZ0dsTC
fJCDMGOlPnLA29OnPezOlkVFfykkoPVkSGmZnR1/SqK9CUbs9pLl+f5QY8RJ8t+I
9YvWSpRE98olZfa704KRLPauWX9C9KGQmOs3I3psXJlsi/L+Kpg78KFRoX9jTmva
k4HpXHYnu6XUN94G0fEgO1eoYvk3yVMvrAM7G26c7iQlQT2OeDkqnXQi1+CJIkms
p+Js+xSi/FHqKmjbE+r1cJc4uUJZZqXx+CdEeoP/5p2BU30itIpekcuj+sBvS+Kj
tKrF/Xr/oMHaa+YYG5GPk6N1tgvWdjOWR6907gvKbALcaVbs5D4w3ci0K4VkwgRd
gIBmArrXbA9DjxKRrmQc6z6BxAlsyoriYvniF8Eh0JOUudBq8uTD9DBUxjGTBSyH
S3EOJVeS/SdeiPvchvjMqEJGzkAPaiRl5r1gLqg/LdwHUXF7GnXnrGVuVuiQdrW3
Rsm0XQRQVTvu6CI2+2sQD9G+drSDq9+oByEqHF6t2HrZ22ixeDavKnl4BzKsFRnw
buSm/1an5SBoKyGJfgCncp0PintP+LULqpaUXuK1BK97NJarDv92YCtlEKRfTVKq
9d7uuU7y0qJLsHpwhyqRlB11qm14QCu9YNGmVJcsgApGx70WsdodTFOvZuQA/dvE
RaHz+Xz2Ij3HoItn0uofqy8sxPsCk0+J9bpl9GTjqAGv5mz7lbA2mW4qYnMcq3oe
2ToDRdnegCWYW/34cFdn1VJzzQhJYafE48pnZGqboHI6p+GJgs9lfFUtYsKmtiXC
tUfnUaccULbizh+fvHZgfZKGq5L4FPSCkTtT5TfZydBsZc2zEOvFWPjjdxkVlTAx
onplfOCVQVM4HhU8lgZk8nIRvibpTix10rSrMyZDuJ5Yd/m5ZBkhl9jGyaz4LM2J
+yZV74rqz94EAQOevz7u4epViYOKyMroTS6Sprzvc6Sxtt61yGQFA16N2Yg2uzgC
qUoVzTa5SLtqW9HCdbHIplqXl6G93MmSZ9Vg/pP9sK0XQ72Ef8vmWGyhgIQQy0bL
qa0GPlMGz6sixo17INEL4CaEjZWQ+N0ijz8aTrIwjbPJrJdAHJZJfIv249rpO9ep
BIx5ZjpKxHm6ncWJBCGcO4ODyGKZGytl8WgXIOPABJg/by88VCSgX1wg9QUvo6Oi
OMayLyzctUxPTxuPvkQMXrzIMGBvEiekvLNLudTxoWBBlKHF1vyqslhQ/qybzD9c
ubByGOXhIbZdpGQykCms1l2gGhH7sLm8F6TmDhF3c0ZFttYOpCNJVzIPs++O+76Y
mettY3EUWIxFwP3v1gBAJkNWNFOR3ryS45zeqJ4+bNDTJwwM0Fsuyfmx+i8t5RcI
v0JwTtYut2TqphF3qqWdIanGMwR7loiTPTzTtmgUVs2euYsojI8UBPouCV8B+OsB
eMfyfpcmyBeX8Z68cQFZ/taTl0cGAKpy5MOTlLi9Mu/kTc2Wk1rnpa+9lqEk4C7y
CEe9MJ34MAL60D2R1iT9CcuPoqOKT/ImU89JbWV5m69017P6BurCEwJmqtIpEJDN
/8Dvc2KeWu3OLuiboR8Klzkr3w08bBEzaDSUfAHCiELUztm0DbQvug6uxJxTQddM
Fcz5Kjdv7u1lOTx/sJzIZwBv37Z4lblsgBzlaunGAet3fk0t5qZWzh3BmN10YJff
LGBIf4GBcCqrbEuq5U+YQ/MXH5P4kkrxrfuo2AK3M7NsNNh+sAIcSrUyRZ5vGQN9
79uyYMbOv7XoUrsEidXZBTCWosdqsr5YLmzk1iFQbuZzz3OtKQTK+NQ38QyJyPCM
V6EDr13DPDpwS5xfk/ChoIAwULBOTZPOUegbyGk1ACSE5oucjG8YA9Az/AwI4Nvf
k5ieJr33lpiMuc+NwkHwct5LMDCQCpgZ1NCWmjosZ684Pn5+mO9lzHvYr1p+7txL
sXF5lpQeibpzZCivDJfS7cH+KrtQyA/clp1Z9gUl2eFwXdbzRxUvxyx24y540vHI
9dNveaIYVC5qlLejHyAx8p76xYI0l49d3B+eLHR7jBQ/qxyJhY6aBF52Yn1ssa2P
gLMGkS9Tewcsv1dJdtG235rWdG8Y3fkgOLu3uGAF3DwCeVjB3Vq4/oKVzgJawl0v
aqE65VxnRAmvGu+r8US9g9mYChiG4x6BxAoRDoyRgcuo4pbVlizy50rjuYi9Wrkg
diy6bl1pV9lUtOIeh+dw1DikcUHtZz+hN7u68MZVaSP4X93rWde8e9Na18MKDfe5
zWbPMn7vi63YMSsVSQWtarWz6Um0JkpoVfGNQultD8p1Ms9kYgOWYqvCx8iEkXIG
mHyFFr5ju76+VT6DRkAuB47sag6b5al4bw5senjQs+1PqXrRyqUICpPl2h7lW8qf
n+Zci3F3zZNo/UcMTtu/D5BYfGhg/ylAaaUczKGiSOuT8uFUcp9ADMAovkkkk8t8
WK624+pRo0CpAbkGpXNLnRdScPn2xgNQaVQHUAFh9+0AkoIxr57XVw//T4FlHEiX
QLflk4t0R8BtMBIxwxDVQfOVsVNNI0kVmJP7qgCDmYm+LiiWAsolrx0L05U7TiUn
xFctrSn5Ak2J7JDrbJhY68sz/42ow4YIMAH6oSOLdkfuez+RohWS+4OCBosw1CgP
nXQB7+0MKlSmgIQQAOt1viAP3gYo/UNWWEVxHwCjGd+Hp1BXEolPZpb/GIT5sJ68
L4KCZDaPMiw87rOG3fI3C7WgvzmN4+IZw/8aQ9cU65qhzPWe2ko/ZTeyCOOwKGVd
kbBumcwuj4/Bd8/hCTR+ZwZyLcyqOX1tU9X08/+C251FVZgXXWV+//A43KQIMysU
M2ex8e2FEbEolcDGO7barvMlXIcdxnGLrLLy2PbfxiEgUQXhwWj/5FL75WXmALPD
mqgTnoJbLPn3127PXgVkBzuZSniNKkxAT3caMOZDaEK7lxAID8y5hOzEc7NsoJSu
MeiockR1qgGsc/go+smzHXei8RKhoEb77nmqYofvyg9s6LJhlni0GBzOP3+mvyEv
5fXhZCRqcvoHE4USJAh8n/5Yugb6x2qdaqb/FeyoA9ek5BMTUlv8+tZuk0hu2MRn
HMbGQ/Xzu0Iyo3NdRTk2X2xTkJt/5PzRK5nAUjN9dZbaToHIJ9HkDBkSaX8QWcMz
1TfDSwyESMjauQWSG8RFJxbwunwp/GA5iPEwrpt1euvAORe62BuCnhcWhAXLG8hY
NcAwFugb57LE5Gycmb6tTNK9YkzwgH+LGb8ZMSDxePKdeW5DBKbGCfeKjhW5pm+T
JandCAeK3+ZloILd20ShjPKUCXyv1IvuQCI0+Qa34AuDrhWthK6lS09A1KNV00GI
FcBXimR/xIdjkXouKEISeEvnc+4UMc86HStjRCm/f/spynnS00CFYVOZ81uvtiuK
LYU2gxooqAyGfgl1rxmt3tCxAO/tLuYg/ZMeFJEUu2uSWvNoII4VFlJkCg6MUFzk
LhUKI/28PapdbSxsUy2Mb7QMRmo++u3Omg7ErHWf7gkpRhG/61tZKO3S9yebXiO9
3Lilerq+nygMcOFaOls7B3V+fH549yiuNZU4qKfK4ZqR9Bmy78xZ4ByMSDdGozJM
GRPlmadmFc3EhAMbyTLCMRLE4Y8zm6S5NdibaKBWvGK1IZ6YSsVuqKk4HAG+7DLL
zFBXLsQN+WBCPj+Pp2DQVl+R8Cesw323RuRcd+VmHIxNpoqQYqYnahMEFm69aN3G
aZf6P7Lx7qvUc9Q2Cqd9pzqpZVQdqSmlwsJ0zb5HEH7BmULDuziCycawF1qOjGA3
eTaOoQyqvagiR3UQg/1ro/4LNPiKF+WpnF+2U65XJil06ftUvtV32MRgc0srH0yO
gAqpd1ymwuNb9fObpWhFfRorlvzvwmy/gH14brUnHDSBWd1vEi0CSc1HmeYipGv5
bpsImB8z0AQ8i/ZouJ9jbg6hgTvVxaYPq9YzTJVeXnZfOcNOH6FdFpkCla15b+4k
owRVEHQLd1Vhkjx9v5KGZKUDCYrEN1rtCDMKuqa49DImQPtnOha1NB1qUOgvOfHa
Ny4ZaNfZj23bdTuK9vtq8pE9IJEgGh/aeoYp9/F2blPSBNsLKJcbfSDsg+D0tMwL
vUe4wPJtOxp9OP8pdeAUSxehVl+XKX1Zb/FGfC0GbBqV3wGsOB1hWUSmKnpjlZsF
Dtd6feREqkmU03D+Cd42cAxFvGTFruVe9JgMFXgcBg3i1+vLfQMQ8NAwYB5LUv29
fNhYMJyuSuVNhViFwGExwbQUfn4CAsGypk+k6TX9Fu3aMHut4E2sino1/UsKFaAZ
mvs7/0ivHF9j1uC0F5vPBbBlfSkBSYl/zv/4Ag6A5bUtg4G8vvjg9ak6L8sjRAXI
9CXJA5ro298nGXa/Xin06lH141fHby6WKE3BQdlE8foZ8o6doLKNuvJg5QAbDSFW
y8j/exGvEJ/PjaAKC62LVCXyPTC6c+eXclaJI7PUBdcv1sTKkl1iPFxCkZ52Z7NL
Iw4Jxq+PKFYwQdiLyIlwL8vvILiAgUrv/ghqvIpEZLYZHkXl2aryOqJ3qlNJnX+M
Iqn1lYJkHYhlMFnl67zos/eeuHk7I9Iu0MNCAATqCHDed+zBe7IOEhtGZDcnX4io
DAm9kgoMrEmjJLwRTkebF7yFMLkpV9Zh+lRKfM7wJVuRwnModIkrE60F9Psah/VD
VTXPyp0KHfYgPtss3ED6QVmggyJO1VbqV9YCKoB0PNu0AmSL7FUZuX791fn/CAdr
YSYyVMbXLzjdsWR0cNHA4DV0JhWqV73MTbpQJ2IO2QZ6JMLA3fW8VctrU2Dy4RWG
v3QeIcVwymwx2vmVNbxXH4+xgW5Yl/CApmn9XbU8+IBqWgvHk2w3HsvhIbkVgauU
xizMoYbXWaSrSaxfulo8ZbsFZj/dA7sfIOF7PsWrkNVKyMbW21S6CAnQbqLesxE7
NWiWzt/YrilrRHWvzUrKkn5iZX9dIx5xEOlYi1iujfLsCIcA2A9pcu4O4pTnrFbS
VJ8cmqEg3bbk19EmgDDiGOQaKq6qEH/xqqLZebTF6lbNSOHaRe5wq0r+/ACsb4kv
PYbxPums616NW4TmA8yOS/umBc9CHzY+14gw6lCjBZMy/AT9EtGbt4BPKzm1QdYK
k1sTkGjGnIOv4aFCbOno8iGrTO8GRZZ/Zpyed9v4WBNxAjpBtEFaI2AMksjzv1Uv
4B0DrdmaLrv5Y5Y3JFkVwMh6q9Re0wHR70OWYe9q3jHTLXWqKbGR+gGve2mIZ9I0
tpRsmuQX+4E/DU6IdzhQH1pV+k+ZSoC8mZxqFiMBEovqM085Wj05d42owlJ/syH8
6No2kM/apFfno9YR8EGp1cLkIPNTJ5zdsbosClpUzXFLDHqRQt8vCbWWOIaD8dAI
W1LDoncIyQuV9s9VpJwlZpGRoi8BOA89aS7po+YHCcWx82H4jTEiGYrCsEBRs/Ra
gXV0TkjYQYrAec6p5X59yk/9cZjZ/tTSaHYhneUd7HvB+bdIXErBsh1IidAnCV7U
FfhozTtm8uc7XbmJpMJ14ryqpbP9mhb/R8ltB1A6BFkzlErfxlZBV0ZEzVo3mUA4
kW3xfnhelNcyrm78jSne4Q3P7EODnRM0Yp8DluuU+k0orVzTgY/9PoqolrVDExco
U348M0r2AUW9jK2Hvg3hgtqhAqBl+Y5E4Zq8oidA1h0qw8Ih9a5RaVmygS35t3FB
DEQZ/DFrEVxreO3FOIXCj3uczjwPa3Fy+8MViyzsLw5aZyV1A9rx8BVTDO9x6Idf
ISnGmXuaHcREv6YdKACw46SqMaxLwyEBz4NFBawfxFC9z7qK7JXdL54D5aZ7RwJo
bZO3dA20A6/gMhLuxQdGwp2uzWmk3o3gx6FrdZVNp9Nm9Q8weSMTTqV/u95cbVQ7
peb+Ini8Le+a1t+gtbk1lVQsnOEjX7Fs6xXtkztne5CZHRhqVzspZvK6sboW0J5T
Mfpd5sEsbav7S4dzB4hxg/hY4EakaO23if9RRU2aenBfn5WtoBdrgZMCFG+f7ICr
1IVO6ippNsAGwCpBsAsY7U8rJFmIJQbUho2qz5SDkAxFnRWr1Q+zoVkfteScKggs
iEddjZ0yv6T/nd7Upr0/jnc4yDPi1rFTBRmtqby5ioHIlTM4aqUmz4AxwWKnhET2
dDnT/0F4Z9+k7GatAEEXAq6V+ivZo0xLQ8UMqmqOQgw924MufO+JPW1T9iJDGTFw
MLHWJMEyG9haqIGYt/gOC4xQQdWMzumRe082Ekr89nI8L8itdOd6LUOnelrKtQAQ
LN/nnf6eZBIaiTzeEcF4xrzpxgYiVPKGTIJrRxi3vsOoyn4dX+9JHhHnbpVUZPGP
EofR48044AHeaV1aXapeyzwXto1rbyBvsWWYlrOhioHa2RtipuunvQUNnU4mQrQE
bvaPK+Wv1PCECnzoGWqSEnc0QGTaiRfFcGUjh0g7sMtQeV3kdzvNjPd1Dsw5IESC
T8Xqb86wS4f2FEmImCXYAu9yt7ojvAlvgARlMA9zXWSF/Kn6fNxOL1EXA+xT6hkn
xPJFGfR5S9FbQ0sLuIaSrANsHxGcoQYnee/2lToOI1OiJVcBiRuLajuuKgqJemNb
XBLBxdpQLw3cb+hCM6h0oALlXz7REiQe4m3s8axjwOrpmFKkR6oxrPbDvV3t1cb1
VYxgXX+rYmv6sOaBnHuz8CXCT9Ky39JXmiqqVqw8T0t4BHGbwnDp/QOBl/AoP9lh
TYfbv9Pl0nB/Ajof+3ffy2BAg0m3TcDwAS5r4+RlBN8UzDWyfGFaY2mLJcCnhczI
EH+j99QGjZv4QXLlRyqJvak9A7mtKFmmNauQtV+kse1ICTXJiHB4AAatGMxv/QCO
GBq1Uc7yajxduINGERnE+wQh4Yy6muyz6Bo6GPbpjng50woZyFhXcg3QQNHaVnkY
mPwIsAQcd5D1RUQul9mHtEO7oyr5fhrDDI8/NGOoMiycD35+Qqp56NkWlMY7Z1b0
KuhaQwUdS65eOtRvYFISBQyqoPZbdpCFbq72hb9LoTyg1oOSoYnePajMiHIdweCM
ppbvH3bdeY8q8fiK3mLwNqrMyheloaZ3DEb0xJPviAW/oY2TNoLvXUjQLox0zYp+
8vcq45hhURY9qB8Xi3eLWEEsL27tBA6bZECgEzsP9ovEU20Aqzi/2ypj0VzuF5ty
enN+OOUfKGAE9bS7ET2D/TJyQ7PM/TGgL8rmd+QxZdazb6aXVQhBzt9xg7lg8W37
nTMUp/woOSg2+gOCBvaxj8PNbQXXuX9IEJxLRduLc52Fr4x0kv47XrFJjCaK01D3
e5sJwI88WhB68uAA9mj5XG54lGqqk78mWdgTwbK9865k+Jos8IgKChNIG2/b3yti
tNRO3mc66f3usKTI+9l4D4eeeEh7zNQNKPJB5Mo5oBjST4onutjO0xshx4SOTcS/
5TE42MQ7yOSxNdKWQyQ4nzeZd3IcuPjzCZTXvoIKScKpj2bPYF/KGQFBpkwUqAxp
PhMl80O1sN3h2yGZUjZN5KVjdwQmk4N6RmpO/H3oqjTKA9AmkPBK/ILA+8K4y6o7
SDOazRdmyZSoKIfh/5wODslBZheE+tOFwuxwvZr8SCtLZOyMyTfHfZ21Cjl8P/Ij
kI5B6ELeo5ZxTeQdFK/PW8+xtGZsCxL5k5DP6pZq7TSWS+LP7EotGFGwxGo9c6eb
cbc1Q+Wc6g1FQEfL+1a9oDboq4Ajir/BMl7GCfYVPQpRooLpS4wkeF5r/G/MoknD
xAsNcNGq9DsrKH1BkzWrfjQ4oZtahNJHyWT3t4q++TGytUboBT35t8jHCmVXbIxD
oXDzUYh/EEBxYnzCVv6RIGRiBTawJvCbayL6ndQtTfJHB92nD+FQLK8bBYKlSUV/
T8VZ20WGucm8LEtO37dedPhMU3JBaezlptvSp6ny6JwUp57oYzJKnuCBKb/Zaxn0
Az0JzZBPjzqwQV+oaobsUc6Gc7GptEpkn80UYXToC04DpR1zmnLc8HCeNZy4KE43
ARE+ngHfF8cOPOcnTDAIUQNS4dSHbzpYM+36hYkCDxdlZEdexNE4VdMSKDwHUNAB
L8C3Ns0YcW/FuRFZJT20iz4mXbWUXy3+WMpOCA2Dt+CNBRbLGqqGinpw8DHtdmUJ
/OuPFgGNox8lpTtv3Z6o1LugnaUR/sd79mnDtZojJR8wfALg/W56BqDh6OFMOacC
gyz3EGK1FKnX9SNGxCkzy7QkWShbf23eWXzANWsl6XhPVQrzqNQ/QI2WuP009RGK
jizZ8JZpIdNZ6byOLANG9zjB0nZ0qnKa08VsE4v3bIXWWWoklJoJlOxhkpV9/V+n
/ja/dOL6GhHg4kMwKiULpxSuLU2h7RmYciEdXbARGX99jAr8SXgVfkPaxX+56HCy
FuGbgQKhKzc3t7LdbzBx4xdLSDqO8FsXdirxIT6CJIutWIUTets32G89+6rGZx3g
ExOijaQL44F4qsIZlnDmYjul3T8gjMYEXRsyBON23ui+rhT643654tsozIYD1KSl
YT7Bjs5OyjZhaajYFr5vwyG5D8yqP/H60NAx+7YAJV8JiBhfvG9nEca6pXSwlH3P
aYjV/f9+yI2Izz8ZH/oGmA/JvbjOCY2sE0o4PBMFFXl7so7jrWGNp8IaEnH2TOuw
g0LkLG17JBIZAmRYZ6SFm+4dJhkvpMoTYH6XMpLBXwZ+t3KzKAsIOap/UfubnyVZ
ijPGzzcvBc6a5jilwSwG3VAhMr63n/OCc8CkTKyeTaa8aBpULapZXo4iEtYQ1HEL
j3BX0D50eaqAEg9xljhIasu0UpJPEqQCZfaKYmiXgHOLgLawx0p+oRxVJsJHnPGb
gRzOjhi16vYZV9UXrShWD88oGuSe+iat1OOcljNPMQjk8M/Cedxgpjb7iTRB/FLe
ZlUfMukSITOlytEGy1iB5ddyVGTgm8+BlOYUQ7lihJUAXj2r0nMalppwXPz/dQ00
sw+KzsUabVpcUvfwHr/Hd7O6v4YA0dBqJs5KAogbl7uCmLza+qSbm3a0MxhuD1mB
zozwOzlJoJaGbksA0oS2hi0tZW1nDiLvMOgNg2yRwq0ENJrtJLEKm6lKuHFnWb3P
fT4r5hatjy2793DSiNgLlCRk9PtKqHAhraxN/UGNdlCYQFC2trm9v46LB5TfIukA
38EWvpr+gknoLBPp71ojloQ/ueVeAn53X+dpcuKjOKyY5UxW1XvnmgUlZ7NBRpou
pAv25nnKgE/AP7LHnf6kOgSzLNbkNN0uyjYdVnX1dGY/Y+AZYDlXQTxAdeIVkGLp
7FP4LrLlaL2KbfjhUasyt1S/9LlPZhP12sR6gKnpOS9FQmc/6s5wngf9YW+5V+JS
WBt3EL9SCBsoYV92nNL2FmtQJVLwDmZIAJmy3tnKdKYIq8eOEC5V/z7auGex4b0K
UR6t0LET+iIP5g5VXXLuco4+1KcBw3ONcs3rwhJzDxo0eCNj7WgF9jAtdh7E7yHj
EcTFPNEuPXObvl4oumL3/RTXeODbdFk1a9o4snAqxz56ARUpraf8OLC5esYb+x4R
bShknrsvr+yfqwJsZBldmMFVNKcmNQ11IhHPxC8dRA4rksG8TgoFnqb5uosQ/0KK
Dl3i+W71YhyqlquBp5SDyH2PAkpmgqEiBMH7eeRZSnQhLKo/sHs8bYWOZPpqu6WR
B+A1KLvK5OZumq1msog8W3qsZJBDON4hc1XrOBB16mQqHPvCbDWJftSRqTwa4m6s
44tQeiUe6AkfuEszPwDsV8yPR127GUYMIXaWZQiE+t23K8bem/oxRvMcZR+TCc6M
Hr4MdoFr800fdK2GUvpDKPS6ZWZJgmhRCPqHPiCFmUqJOPEJtOaeIAktJUWk6Qv0
pIsRQtFhJp2hiNy8s+spMjzIRSN/a1MvrnrzEn4vjyyJ2QHpQWY8geG6MMBwB21B
HZCdGKMN1O/lMwYzeHfnZIjUgHWfR4QY1IU/Aw4QQmsNxZOayTtobU4e0HlMLxbA
o/wIu86f/QyuH+WT2lP9eq9fOErYkCycE/KJvSOLR0J7+eq0oGqGuLIgd94J8YIr
zAh5+u7IX//kuP5A+1jAABK5AHZo/b4mEsbKhThEW+IeVcFB53TPzd+gR2JhqGyq
pVFiG8rXxsZ8fZDtdcPU52aWBI3FCTaKbHA6b9JShYDu73NuoepkXZViHe55zzcK
GMsK6XK1JA2QtPlT5uMqbbXId94QRWOYhRggg/EGhFC8ZNZmSpaRnbm6JNSov1Jf
H47lCAfk6CtAFd0Km8CzcPdMD3VF8tClswnKgLLNIiL4ewBAgm6LrUJSUB+KF/dh
hZ5CIJDkfwaqG+A+b5Y9YXImzdMnxt3BVfJkLUDb2PfMlR0PhrfLfv12zUPobcM5
11ZKRlBT1k8tGRw7uWEhtkCGIW1vYEmdhxFC7nJTvJytx5QPx0Mjy/wIJmaiLJVj
RXKQGqIQmQfJQ97wDcGrtwxOv74itzTSmrD22k7xRZtijVLxXWCmzqYqDfZ7ZbQD
L7bjLIjOi+lXzEDHp68kMnBtbFMA1gWOgbvczVGnXDUbx940/5vpDc9BCNxIahGG
n+8rarLVAHNWGA730GvQZB88rSM9H9kObOut+i0zRdfzpLtBsXB5Iwv5Asvn7v/l
2V5e6FRJG0lqZ5cGDl7IwlM9MNtmjZLEwhAVNH4JHlQ2tBGFaJiFdWO92777X+X8
xjvqW4KjauxgPyMmWpoTVkbhwFvf5uBEC0chC0Ilqp15FMALoWpP9TYK8F0tcNaQ
awlVpVdEvlWbXtGxpqLriHMraF69M4E6H+T7tZRp6IQ7TNzvvn274z4S3RgKB4BB
a+6Xdvejau2YuYky+ZG90gJDBc9iqZEq/Ip1Qr+8FiA2joP/YMEoMQjxTzRLSSXP
KWyT1TnupigmrX6Pym4926wJsFGQetFeRS5rvct/gtmeN4SrB3Mp/Ya9ydrDX7R1
FggZn9dLBoM7m5iAeiorEa95GMF4mj9T9aYRygXVIxMmBUTtmfoj1b4jVyG5heMk
byPtSAmTzbB9r8O6N+0OQIeOfXhbt3/g5h/m53zJEZg+9JrDm8Rilcr3xMA8VVrE
Jbqvp9Yg2lfrfIo0nOgoUg9hQEtIrQim7ZJPFXH9WC3S3O1MntMf1piG/rWperN5
y+pKcL3VfBD2CncFAJKUvyqVsU4e9CdMyueM1QD1Vh+ZJdxwRM+ns5BmRcEx4OdZ
UB0hA40k5YwJwcl611RGa2EshqZxXPQCumwy6wLNa4mQE9ST3kGlT4+O1nRmm9tS
mTh+eChfjkKB5ldwZBz/JGyEUbMNCECuM8KsG8OSbPChX2FNrHsfqLmav2mfSnHk
lbmvyJmZ9TXkQ97JK2ktsRQnqU9wbEDZcbaFrjwoYZmltbX9OlQ2UvFVWL2uCEIl
5cQkrcCTtWtPLsAl4/TdCPzBO/+X489TCwB5SYPwHgrle/uISF7THep+795rJILu
uLdt2TUbdUXIR6zX5O5tSHtb4jL5QukAkUXzUvy5jvHyyssQC33Er4j6C1PI+4C5
+wdo2XKhU4OpGNp85KjfFfe6PAoHll9QbwtYphr1ykTBgZxbt5nrYBgG0jcuT/9Z
G8N3uVKhidLnmnyVYIENn0qj8sGDhusHXNCgn0vWUDPunKRLifMmdUjtpdFmkLPJ
2JiHLMwV0C/1EkIN+/FNx+6Fnmi1E1/jIgq8StgLi9zNyCSFuinExAunxzJlC8yn
CEUhzvJqASAK5MOlATpvogIlDPpiJg+IqwGRXJcfdO3tNSskjcv/wt9GPM/QaVkf
EVyaXr83n+Eaz/GV+odHrnYdZfZPFCKFSY44NINjbPKxY3rQ+BOd7/VPHalJ6cMH
yZJvfpduSNSpWINZWrvctusUHITQSPXKVCnDvy/sE9RnoZzDZWcWJQElbyl0Wf2Y
jORPZn9tDigCDGH/2eSoAJsufbtQFANmuMK9ln1FM5qOu3+CEd8sJ6y/K6R2TOL/
pdP66mPcL7EM2RdwTjl0I+IJdEerI27KFoJ/4Sbjf6YvHBSWIgFL8CHQHYpYDZrQ
NwmBbU+KmuuvOoUneWJh5qOXoVEs53vB6jxuLZZmtObzmHJTrW7YilEct1r4+Wwq
Ze4x+IzdOMjICwTH5lGN/baPb1L51iDidjHAVTzs84YtPS8CKHQcbjJ823wad3ON
MDZgtB0BJuRwy2MdlL7VJd6LuZyYJBK3pxGCcEOxMDiFPkwyTEcf6lPcqTmKgab+
OwAPIF5TrnNmULdzbLW1/91rfOesc7NkaVUixK4ZIparBVhgqypyhWxhgge48GMJ
TKY1AJ3wTDbgzTi0KroLq7rKj2cPqO6j7ZEs3W8LPGcTmzHByVTXIvihvSaEtVoq
pJ8Rh55M4FGZmR4zp8RQcMKrs5BZ5shJIT/Uw5o4uJYIslovrAI2yjc7MJnKNMnT
MHvgw+FTl+KQjhwKGeyODMdpJqQrhdg7llF0kD5Zk7/vpw1S+/+kYPLaehwaF5QP
yEiH+W7GV49GbOF+QfOM5797+3mXLPHDahnnPDdJ3vnWo6c6CRlr5teryI/n9bGa
tUmcBwIA8tp0T9phSoCeILFhP8+NHi3EGpkg+K2pU3LJHQSCbYuoYqNCqy7AnX1b
GnBrr/+awOHSmG9hD0ghWXeZpxJU8/5NHbzs/FfAWPX8arDia3YXyTgx2tx08RWg
JRhPkrF4hW3PmKhdWSXmi0gFngCKxct/qDI53aM8cX5bK8X8lQ5QXmeNfE0cutQS
g22SRTUvHkkuyZ03WWYMtrxnHVVFE/5N5SL6GDxXFvtv+n9nr0OMSqtulW6cjcOH
IJ4wqJCoEbdNgQ+I6HZtcf+AAFa43oU33s9df5rDir65FD88cGviNZgAYgEgxZCx
5LMioT19/jqa5b6crzXaPbaU5gXuIe9F8QGRI2bA6ODeo0f0l6WpMgvE0RddlxiP
w3/w6mBEZUIOUJJwSyGvXDK1mHP2jE9oO+LQRERIuJHtqmC9va4c8VlsLsSDlf45
Azf68FQlJYdYEASqZ6u4SRlVhgUKZhiNYh1z3RPNxXvjWlU0eT75OpLS6dRVnmRu
2uqfR2nhOEubeko3HO1VU20WQvU/YSOtj5vnHZS8dqtbiCTboG3vm+GEoZiYDTKT
U2rXWrkmjndhwoSeZ8iMAjBQxAJ028jZbQaCxA0DIywz+JnBqy9KOoG7gFHlCALE
PGKDe16/1R4Yzei255Ur7wcNfClM53pfNgz6/apwwHEQRO61Y9iZ4dk/DIZhXr9N
aRaQzGFwioVkLMDwgXcorq+NZiQFynUdNbPn2Xnb9DeW5THvpwoqVhgDdqV5jUzm
r5V/qjWUqu0moQp3Gj5B59FV6w/DXnYRN6+vFQ+DP2OJ5n/qpd1l/pOm4salJILf
W+A+XQkhjDDzcmWENAOF2tkvp2bCa2P6F5O+l619a++/9ErTWcU7hHdiG9/xo4fw
yr5NOMnKitcheKEbK2xjdeNAkaQWcG4XVGA2lYWuXqfU+ekTX7k8sjegT6+jg/ny
gzpB3EuPRzKoK/jnX7UUe1UT+7AYJqUfnNg96FCQVKxRt/ZurFuuDOff5IQL+fMi
r8gOUMVtuF3khft0TgciTy7vsCGyQkJHZL3am4s9Tmeb77yHXlkJPOEPBl49S8yZ
zRm8vykawDm7erWWVl+0hMNsRuiiezj+dukMcpuPVkNm8EpzcgxVGuavwsUHQOjV
bXyh61GWKcQ3nJQmwyH2FzzfANIcsXqCtNLwSPOxTdwlGoNzUUsKKPdOseTtX8BE
KGWqfq/I2LIh1emP8NRzrMyET5dv4kcVvfBLyO7j/oku/kTV5SHVYVUXRKzSmS8G
Xl6uB833fyWmJWG10nZwq+oPAQAGYQTejvL8tKh/oA/JJ3R6SRWNGyJLkX1/ThfU
K5nYs0GlUNF05nRDXlDbYxClwQhnOFHJJEHcHj34WXZRUJXJUy8s/otcsEHev2MJ
u3Wa0trGRop/F8OVJf4dbVkTGN01xq+vt9fvI0MJfYS/KDEXIja3OWyvTVyRjXq9
P6rdciVl1FDT8NN7HC2/USi9wJHYev9x+Ags5KnCremwDBc4hY/ZA2a/ceyfjqND
38J/thrzZwjYyZsgHJJSIQB1qISwgC+7HZ9F/1OtLGylXRzYV07vzZen1Po7dxJM
jJMb5plEkei4dXtMAbHCSFXr8gWFEWu0NFvmPSI6ipdO7X/ARt4yk/1S2WV9I5aq
3xo7WApVYWUCI6g3PKOqRW1GD9DfzdUA1IMPeyQhfSqO9PU56QB7+VbKWP4maSR9
GGknuGIkMY8Krwucv92t9emId99iTIjaBTH2YRBowSuGiEFaYWQMUl0ZZNW512v6
z/FXT6R/0FIdXHQjbcyYF+EhpAhGwIupWjZ2U/dteBeKwQyinJzBP4qqrzQVc26W
PfARTXvtkGr5wEvhdk437tj+m04fUxuqLglCuk7NYezgl3Dw2iJsTF+HX0+zXP41
WIWWx0/GkHiRLoZgyXXJT3jZs/tjiUXdO1JJQuKDEmUXIdJ2l5ee7Zt2e8ECSSnc
eNnqlC2cJUZngEJUYetXFIEeNmeIeI22DnHpHQeEmSnxygwcGsEu+B+3AEtZTSW7
egH4Ib+0l3a81uwhK/lRKywDLcfvmliwHQLQee1peAh62BIBYrPD7MAMnWDzKuxa
gt2DDKAe+np3eyvC2TfX4uAPVNVx3E5EF3xv2+bHTjYuG1/G0ydrf1R4R9HyAqx1
J8LuGVGZZ0ibJQjgXZaOOFK1UJNMD+Wb6F+kucoGN8nK00x6DJzq7/VRoliDJhI3
m24Zh+4o8V0JhhgZ645/J+xpbqX9Y6PbtUP8El67q1YAd2dmp8B5Vk6+1gw4dCwN
YnZ7BcfgoBwLq9hkipzhd1on1L35nnYUhSLB/jrsoJ2tkAMl91IHOGaZJVpqDbG1
w4A8ZPRdrxjPMxJPGiIg9yV3idzVCIS3RPtp7lUG8x13JbgWfogiN2lB6iWMKlcB
JMZ3xvAt4OKiCKT4CK97iqGVromw/zitiNGbz1dbDOoTjPtcz7B4+sPgZxz7zeIf
X584ZP24EMrWcsTuiN1BAuwFoFIqQx6rmWe0MpYXU1hIPoDkota410S0C6QlMw/N
n9KJvhm1a0OcpsY3UbXp8GF25s66u9qiMdiFbsvKrehFTJ7HN5TTevVCLwFkGyf3
zioOHV8yxJ1rW3K66rGI2fiDTbN6sQeyW1u+SIfa+qbtuUqUOZ2eXOyVNjjcmgeL
6zD2yTNsMo+jnaUwUH5+zOqZ9v2iGFvnK+c4HvO5YmzeZc/gVPYiXCZOyF9Es0Z6
kZ+kZGq6SnBpW7BekMoSuP8k0HSZNpPD/V56tVL9N7VMWQO2ALyKu9XV9LKEwqHC
zU6AkpwVnW/2ky0w0ZZCA2LTSw0Gt6ZY/TrHPPbMU3u+e2PH1xyLRWEN4YJ7FP1P
Su31EWKgA2NV+J06gzifE5Wl9GEIznTHNs81x+D5pyl4XWD4VJiMmcc35sCaV4Kx
dfIQrSgxDYh5GTZzhLYivGowfaORponzSXMKY4C3yNr44qULoHQvq+FGf5e2f046
ayjNtH5w6g8ZQtJSSppInOm/zIUI/6qqXL4J1wZYqxZ3wCxMlq2WoNQAB+4IYa3z
4/3PR3X1b7fNqLzKBIuSnvwf9FHfy6y0HYhzsEZc/6um2JE3QoeXjByvOXHSmrCS
5TKrY9yZ/4htyZgqY38qd1LtUOUjnV6Y4nNC5vzmLcL+vIy+0DEihapONX0KF4Kz
YFZ2y6vU/dbmmZQiAv3ZQUjYLlmXb6XRUAhntrgnizTkbNPlW09R+71+WbQ/4RD7
gKfOZqf7dVgFSkb9VFpZk/Aej5/+RRZmZXnY1xjcx1h0XPCh/+indHwqQufQ23va
Wtf7Mla5XIqAch3eQ8FZZxKndLOUB2ZzyV0Juur4NqxqwqIg0lhxRbj6Zpv630UI
5T1Ck73Tb4JOer5hBULHCMiV7t0/L0x8TswG9SLKeUuSI6ILISjf60/nH8R3NxQ1
gNQcSJ5PeFYoVTV5hGFXhjThHTvvPafuJ/m1SQWOuikGsso+ax/G0iZLGL1KPK47
u7TdrIYEE/bMPCBDwV7lUNLr2J/4yt1tgCFJf1A7CNDPGce1CrpmgQj4YsUyAry9
vvIAxYC5B1sA9IfRKDYOT2gfh+iWmoc2HqdS8d3bOmWseeg3iM2G+cRcJDyEN1+m
+p3OnQ8PfjQkjbrhKYGSF62Qj+0S7rfBtgTnQgzx6qHDy9DhsRuTA+l69zEpTwh0
sYd5rRleuR1sGXc6yDc8L2CrmzIG4GdKrLoi7BuhuJ22qwnpYELNU+87hcG0zQ/G
BlM3nBP2+UT0v6AxBYwfn5DYdDQshMybhJ9yNEoD6YL54hi+I884n/EPcg804oqU
AdFR2N+SqJU8RE7cOXEIYb+H4RabjMVtFlg1TgcX6sLRrfp1mbNS8Fhgw57txIgM
KbNq7Up/pqCTp6DpwpaGmgxImMdmXL8PSWygwsUoU+FsxqgScOwKBApeWcVJglpV
8GjVKVa5Iwb5gcH7DCjBy0F2SpcJ7te79v3oQJrk2Roh5D9DG79PjZi5Q+jTxxmk
k3mO88UVipD2e571ZYBRw5AuBj8IDx+mMRljR/rfVpborUcpgRIb+fJ4nswRk1aQ
ZTr7mkY0316I3sp/Tt6bkRI2mS4PKh20DPOOPQ2CJHS+nO52JlDgpblDQGHU423f
ZUQEwA941hm4giY/L8R3g475UvLRdc/r035h54/q2qR2ssowLcziYXmPupdCI7JG
rRei2L4daDseXDCBbvQzlm6r1MSShA5owbxNBmOAu70/9cuhtiKh1UFJrtrxJo7/
LJBOyll4wfuXs4qVgY1rUfLzntTuWx0PkTGHG2/rR1YLn9ETdf3i+CTwVN8FKJbx
B8oeQrKr7sSK6vNvh+yu+KYN6LtH4G5RhdE9dpR2R2/PJOEgufnvoZW8z9DpWijV
dv/VaWrDpAiaKNBGJeat8ZprBeF6O4jV9x1YW8kbjSzLBUBid7V5acoFAlkfiCmk
oF7jdycnUHTEUv3eQjkDQe7jacNOsSf7GZmzp8kfScRz2L9AYYGVRMeyLCLM5DDB
7o3FKQYL+9VlJW0oHy2dZhRDM1/4Fm1vbLDBMK3O8uc6EfcvNNmIMmVEhlnmFQaZ
0fuGzIYdHx8juK58ckDce5so7q1Q01hFoYTcnuLJUK2A6FixSqcXTF8WEOwDIbCj
QnDHJ9NWZw+sr0lpIxNu7ttLnPjihuIgdlDsF2dE/69TLvZSIaJT/r+tWrvo/QSs
5Qc0tTVYA+Ea2XmIH+PVodObkx8tJkw8AYwzcBDdDBn0r2BNoNGxbofPbAStimxg
VK9mPcdMC8CQyxgBi3LFHgon7iEhQtrvezUcLzATIMTjvn9QiZGHbrUiwDIVfIaM
0lBG1VNO5vaBbPMQd6lwKrZXkKf3H3p/L5A5myTcRWf7J74O6GFM8X0zj3ATALQR
97l5q4LBfL19xwG8v+oMlR9R9SI+CYN0zRoPofFZeIXGKoxssiQ3zlEgCm0HqDzI
DvWq2YGQWZex09VmiNmMaxcZqFUSKyRIOQWVHz5+pIEwUvK7pDSKSp8eg+VoHo1k
hnOGbapKFhtAM9DHWC8uEsaSeV/QAwtxnrWN6L3wdQeH2CpmGjOMRdQffeH7MkWj
Gh6ISnNrYRK5ahcYP0VWVvrEM3aRL/eiUymzN7RAoTeIKCXIrGGs3i+jr0YnH7WC
va8b1eRIF9YrRI6NkZeyPTLQzFXzm7H+LbFCr7fpZZThgYu8dF+ALO9CCwiwwcGZ
LLrAReEf/nP6HVlEcwdVH/ujIb6pWJbE8/GwpRTBYEVXj8s822Aby3OSCrlVL+8x
E7x9I5bVo5kKikQ7/0+ncQTuqp17cUzDNGLa0IyWRaTvHo0249YcafRVzMxsKT9L
ho3RgFRq1JcMDjdKSbmi5Qtk8xIrqg0A1Py+Q5AijjaK7HgDld51W4tzxNUT6UzP
r9L1oVTF1t+AD9D1w1OOYHF/3diareCHGjIIHdB0FYVs3jog9K8QMpMqsgs9G/SB
nOs1MKsJ5QO3jNDh4AP16QcVG+C7mvADN9NF1lRNoVXuOBnW1p/YDWLUm833Vv+f
30vbQtMIpkP1EhFrhyczND57LHNor0MB7OiQaPSAmrXrjb7jpukKpyy+H/HyVRcQ
/BaczStp5yo5VgmvVPItJc/E1Xk1lkXM1jaJE1yRg7WkOHhKq2HzOWhJ9prRT0Fx
hw5SdHEzw/xan80aFh8UotCpNegPZhUz5eZPVsY/PRzwfgzEo7m7ygGARI35KmkN
gXUWYDIly6RVEYh09mzEEXgnpsLDTkZc9UZBJ9iaMhDCZQObgqV+vGUHp5NCQQyA
uBvSX1h5QbYhmmOgCR2w+KUhFsx8wTozjsQVUfp7WSCM/6h857g2QHG+XVFffzBM
mFKzAyOV5A+90hSQ4G2Q160zbtQgWtTAJOhlRmsLeNWO87my1ENTy5DCJOFEVIIS
2L3jsad4WWHRy0cUliZrtRjduHH15w9S4ZRHiqZnXevK9X81eXaiivQD2qZlGVDn
MIY8bl1gM/mHTtFJRQhcuTw5EycUf9z/AQD+39Wn12H3XemQonJucNQrBdHQKQp8
QYqNIpaZKTiSey8WfpeHoKY6bcsmswVzx3YxInpkcJmgSnznt0UHW50ZCTQ/xbX6
WlUD2K8z7BxtacxEs+d1ZnOlpTzC7Xyrwl+OQDZE8kqQ40cdeltzHgsrFfseRffF
IZbUHo0SCvJFaVmce1efrWy72iQBOcppTybCurWPccnk1Sv5QwaFq0n1tmUj2/Rd
FR3SadqQ6Mc9XRyHHRiGxDQg3GA2dW284RHTY9/0E1NmG/Q6U+4ZU0KWnyCIFzdd
rxu1AHT3zLUGObwO5d01WJo+IvMa00crORNVi/VYiWWjR6JgYmHZmTj1TbcoXpkh
34TnwKqQNZkxdpiwKgXZwuAsbw6+KiIYJ6m0W13xA7IWHJ6lAu1nMkNtIC+p1r0n
djeQPdcmLOAo5h4IerXa6o/E+Qxo7hmYGhdEZ2qp7BLqYd7dauJwtjNY72Q+1jAG
8HXkRFxTpR7tf6bokvW8xBIhiwo0NnNE4NkM1gYT03pg8IWPYzacEwc/2325gDH+
idYM4RLoiKC3wICNrY5bV/0JeRCDk/0gpO0UoOI54xwv6E7sI459xhVLNLKHEApx
MPUklo7MfZT1IgGn49eJWspLq80oQSh6d3+dNg/kM9KLtJR447oSZ2XUfN7dSYL/
OB4RDprmtfuEwa5mgXzTLcfFYtRDUhJZtEZZsPlDJYWVA0i6oxYTgksTrleKpLk9
+vWiDRrweP+lzHRPwUfEokcyAqJRYCNe6VU/4DJLrYF11z5z2S6Y2ENBXJc3x5cH
Cfci9P4oqEeC8dgMtDoHRVx+2pfeIECj0dbuQWaqjWmEhYjZc3DXjQ7RS+UPjadY
WpOq3UQ6tyIiooALZm2A6Yrx1lwOSmd3vQ4aiohrSltgy32I680kIe1lfJ8Ehxc1
Rkn4R4XQ82V7a9tyxychig5LxPdHeZqazWs5mEWK+1yghus5SEN71GSJqtYeJhrn
MMnFVLFuNfjnpr4Guka/LWKNYOfM8PLSGT4dRfjztQeVwq6dpMv8HMLra05FBdCz
HRZ+DQSRM6/v3/hbNuhywUM6e7kU+3DK0rTBCBeBLEI0NO4qg/xGXO7heNyrpMbE
4CNNYm6CPMXUWOFh2k7rYoFNyHcYWYPwKTJb2cGXtiFfDpFlsBW/tJlma90PbOKz
zhqwBvypKDvcUecX1iAMe3CT2jZp0KANps7YxM/KOu4wQb2z2qruDpk/tyxs0x+9
QmDq6tUgCiiqaDOG4SLy5D4zk2Na55mJ5QBn6nH6ufGbqBZIJ+VVlMyJEiVR1p4J
MzSLDfVufCIRZd5Z7ChQS/UVzvtu1kJ0Q9BuHBE2MIPPqmDWDTfluOR7WjMeqvi2
fpNIGLsg/tUiVGCbpBMoLgYIpKypRq0hzP4ljkxOVu9/u9Nr8Qnqv9QYx1jlvk7T
CHCsmhPLYIR87MLS2JmlDXnUTP1c0f45CJNUzkfd/VuSgCfWkcFPlQXgvXHfdhgp
pKS6NeFHT5JbKDs4NxM7Ug55glXXvPA3wIK0A0Tca+vX60XhP07a2mWf5j+8mOoG
1KtItL56t5xGRecBzhg1fcypKgqVWNCkZWnfoFf6qREf96JatcigRJ2vujV85w0x
CfF+7iBrt7UXsPCkt01WepUAW6faCDCm4P1N93n7mLU+teZIyNOy3Z6wl7uD0hDd
cIor0ipySNjEMwFOAYN+y6Yp9FvX56hdsMqw/EhDjAclkaNe50b1okPrLHeoYbZj
+NlKyI1L6YByTUBdC4rWcszvcVRfTQ0FWtx2tvZ3TTM9olbh3tmvZhxpF3ouQxqM
8dgwhh3Khst29NT0v3XsHE1eb3GVoxqRaJLTrpbB4pKQiBGO5AlwWxDkYgpK/8E1
PLKb9wDcsMbTpkuoVZiO7hdkkkRhKxnnGhWYeTLFRyZEFl0TPwcXQyiBXASLswOl
zqwhqxEUZ88sOXPY25vJ12Nc/4bEgsH5HSAj1lJvYsjynf+slNPVIVIxJydqfW0Q
FJruH3YumaUbQsaiuQcAAg5U2yUUzYTXSGqWbR7rclZxafq6MB5TGLeM3nDcgKcP
9xVsIiXIJdVnzIMblpzwjh1BeMrrk1BAtSZ97sRzpiqzFsnZ63GFYYQlQHn+RCDI
sPMLYPZ0zr8jaZo6soI/2MetFBeauaSUAJuRqY4HiYPxnqhDiehjk7TzP/fqgBjz
h69MH6A3ROAKg+hGSLviXE+oEqYJiuFvybvH56/IS/LoSM7Fna02zsCQezo/mAse
axOxx+vla4c83eJc8/Jd1X7nOYS/4+2B/uY9Otoz7DlgQYPJMMekULAmhvO5/Ubg
vTgI+iGuTAG8wGpTJqWBdYpluETWVeWmtkh21F0hjNljkiaKY93Y/w4r12jvFnna
nT/l42wm0fQrf4gphWN+qU8BAiLTj11znCE2zKqwmY52QhEdoeqXb3ftB59fGfsp
Yny6m/s57ihuDeHO/fHYLnTGbQGDd+v4IkaT5XcRz9n0Mf0CInatsvBZCGUzewHL
HSzAd8cmwV6mpiiEzv2ZlDukH/0K91B+39sATkYEfpGPS/EN44BvCiXeGeI+l5+c
cEYy6dWv25RX2C/65XAW0kf+JWq/SunBRb4xIPyJSO5RxBsyK9PCpfLXdUACrTlE
W+FjIeAZi54egZxoUEvXoZp7Y0p4jOxlsJO/xyAchUR/3/mKNrhg1jEWBqOCGFVh
sF1vbfOQRFoN/23U0tDyxF1G1Ozggh94QUoMdOurotpKY4sF3lIJMDPnvayjHzo5
UphRYWPsbr97eP8N3KowMp2Iel+5Q8ehVbocE64tw/lm27kjLODYua07pKV108Hi
Mb+lBsjoz5Q6W7iY1zICyVC3xbXxvn0oMsy9f872a7KZOX9vUr+n45+EbjQFgWiM
q/Yt/tzWdh5dbO09OFOb/LDM9vGoNZsBKJi9BoH5LmBrtRUp+4FNhEqQBpf6mcqI
H+MQZ3C6ov92qQVT3I7oYjFRkyr3uFrg9ZapAT+0vgdUP0Ml9zto8DPYQ4J6GZ8t
txdW60S6Ttl9QBck+2IuC8fR1JmfJk1+XWVgJun8eeIv0pmLOh+oFtw5BbSJoWv5
fOnpplXjiX2gCPq405fvDhXFccWO5eNILwtS3agR9C0IygHaWK3mLtUHIwsi3bPC
r5SeY7tCEENTsV9Cm7iNsvqiwCxlchnVUGFYiZ7QFQUuxGGcfwJKeygC9G7RxNJ0
LFceewgCn8YnGGBgsknygkGlpbsMEw5KrrO0Lgk662Nvg/iMENdzYxlyeKuU0EGq
JYLK7BVJFDdHF+Ck8kGaZf24FYuOGA8N/URHCLRaHxVpyUH6ccPmWIyGdW794hgb
lj8+lq0gO1sTLva3hemWfcpuX6L8MrEGqq/RDxz6duY8/YsxuDJLHsZ6tXm1E5/x
T564RRCpRsGZK73Tu3mYN0ZOc7RMEMgu70SLbNGOEIA5b0TCdQFhBT2xCIqRvkQo
4PxmbRHlnoTkZYm1NpVj2V6psiwDTqFVmN7/gQf/rDfZkIWUh0sZfjSUuhKJWOs1
XqPGJ5D6U38tzk8W3H96ABzhGf2d/POOF0QkqnQMm0nETEzGUsEYOopoLR5tGQ7m
f4e7P9a257FXVEeBngAvzAyq7XFheMoqC3pVO+D7C28YeRuEebLK2zsBM29H/6MO
KWMZ/Lbbh0pz9oHAj1OW0Y7vGXbQCd/GEvAZ9kjz46HXW1Yh7HsaC1rqzEVGjRP4
DivpYThr57A0PT/INitYe4ykgYGzR8Iog6S+3CTCpfop3/vDcRw8XlRG6znN1Mhe
MWB4Wms2TARwAcTSW7wSsFEykSE1fjKTAva6WD5BgSV2TUgh2pYNnOGfgoyXwusS
leKnQVubtrmU5Hi197LVLG0GmI0lh+8aWubDGP7c/+QcqqG8To+knjt30RkMpk0y
PeGautaRo5Pww2n4gFQ6wPbrOBSq0TK148CMk58YeNBECAs6ciJbs5S2f4gHXzgb
zr3A5RnioONEztGa/bHnUJB8y4iuRLzj6ByXEFXSp6hPmTTNJSzlkNch0D2ree6p
z7HYRVQ9xeELPkIXBIU2rMoUkhmz5yzIcZgB0U1QMiIbV5gwur/aE3vUg4mbgCJb
TXvMiMAY/C5xXxe8Y6PBeEaUqfh6rvcWGppg8llQYZ3e+4Q6mUdW9lJOcaHp9zPR
ZgkUXW6C3ErqkegwRmFoimcff7CdowhrV41ha0hUmGWpSlcsLEOm3ByqAJ74u8hG
N310gNefopB02fNDJrz3cghhqWRgHZrcHTl3qHbhJzL28svnTFoG33MLdN+ODINX
xufPhUeE/LCCt+pbRLAFY7DUm6a/TUtJeXP2q+IjTi3+FbQanL13NoCM5jYFZr1C
49mtyEaw3F9AZ6kZOdYapk+MqUqv9i4BcSiphKMBmf7OeOVRCXMJgANk+frId1vO
gzmjf4T/uHbrbiWkvjzZ8MbLvXho1+SKuzLAo2YZ+D0fdn5kRJibdBCFwkke1NA6
ygMc0UJ9zeMBEmnpFuHHP7pg2YnJLWgO7wk+YW55JH+COLJZp4La6hll368Cyj1g
a0WC97vCLCIw5X9aCvTDKxhAhRbZvQeHqPYQc0BLsXW/i06GXvCFVSFGay8CfuE8
8hSjgdGGmv7pX9foIhOTcHK3BoX8A4Us+IeaeO0a66VYslXK9q4qIVd0DeYEi/eH
eJcnOgl7yEEmzbVPAh0M8onKrqp942If6ELXCSxndkwYhh0uv83EHZaZ6t6/WvAR
g61PbB+4b/CXqh9xCPNN+aXuscToIcVHJS+8rmFNl3UMvz1IXONWnLwqUkOhImwY
0VIDKwasufAjO4B4ELx4GrBw2y47yrjVcrnRV5cLhfJT+MRqchWVPeTLzdFcNua+
VX5AOa0nibG3WELl+y0l3hZ/ieRwnA17hv4Fhi7+9hYSgjl62yS7qPHDDxlwTd6k
2tw3MjqrDDXGmu21uCps73Gv5gN803ZdZNqJccwuo2W0LJc7a5mZpzpM/GGAJ0Pg
Xv+9QieevFseYnrCo0Pt/4DPXE9fFNoPyLGY6G5HKbkh7f5iZObNLksbwSrbHF01
bmlnsnK4m/QpviHZVFOoNx4nmbTES0koiDrYmYDafJVq55A+RIwnG6YvsAMveABF
T+A7ehMDM/5vBywo2ifQE3EB+u3J4zwhk7n/NWQg02JjSTbdBKOwy5QHZVbxRpOg
jEPYwUWaCrkZVeoHJv6B0mcZgEKvyhuaARoxptCKfIwHIDaVGnPw6Ggcu8yRGSxR
nw+KyyvzZVkzdkiWu1nRwj2W2A635d7bbYBZXwC6hd23XARf6pi1GEA0AUUAedCy
3VARrN9/r1uSUe8LdjRsByTeXJIbiXy2Zs/UPkLfiUt/z8OP/sgcbxpGKSjKt3jl
QlHUO89vFl4kwmp5rC1WTQCcAWfGmRs89HDvFxGsrskdszyb4YQQHXSPz7hfGXNQ
5fCLhxuunwGySqvlfc8zdsKYiGQYiQZVBsMxa2bIGwLiRLrChcD6Sk16gadkt1us
vHHOue2APWxCQc8lOZefkQkweW/YZnhXVEobs+BovT3lZVhPmrJn0tE1iKOrix3i
VNMfScNnYv2+jfiW2TlwP+tlhpdkhFxnjov+2HxAf9Itg8iRRROr63T43YG7GAZr
osoJT1vSYv5FMnO6aeMY3PSB3nmyjFre4fkgfv8tEUMPufEDgdNQ2+RapMgnn6h9
beKHBYCHIOKg7aPkTLI6MgoiK9ExF1EzQwNAamUVTnt8TFFL9UGgMxQoLvNTgc96
nilW+t2ysTj+WbUeh/v4FRrmkJni1ixxTcXfEg+171TwO2BT/ImEyZpYMi1ydv5f
/6Rd4rkxWdU2iHBOBWXsw0LpGzTDFG9v9Vr/N9iQGhAdA9qvLYcae3MMrIShPe2V
9bT3Bc0PRphEUcf2YrAzoAUwNLIVpraIQY7ocEnFQVyVPd8QsTMkvGAy1j0g1u8G
ekOlPcrcJsggSznz6KjjPI2Eo8Wzvu3RXssZEB8uYmM8W6EZA8X9rlKOBJp4d4il
ENSbL3g4Q709+6dO18rG6BXbLmQjuBWX2GZeKXQFTU+/3eYEA3xzL7EbI5w/BWE0
3SV2bVCVvyRcar8+uE+fndfSY7IkSK+C3ezXkvf3DCFzVxVi2JRNKjOMmZ9deqI+
9ITswPSSiqvY6NRncb+6xPKRoXHG2pvb4/Y/VEvmmDel8h6kOKKBaF7nieywbqmZ
nDeYYcO7joLYgCHQJ7TbeizJ0TO6F9VgQG7GELYjakYhcMc6vaOYY5uUKbAEvqUY
lb0nMad+yKuaq12jVrxfVuKaw5ppSpaPelmdq+WnY7v/S0hxA9eYGEAzYgOYW9n1
HkWZzM0iLWu9Rc1hzLTDbWTj9fM5gi9W1+wnpc69qjit479R637dc21CFqzdBd0s
u9M70RLBsulraKJmafLnA0sBP9bPArZnlhSvzQf2pTse/WFbQ2065OCAkL+Wnt5I
BaX2z3/FWdhAXBul+OK5imD2jtObaAx1X2EDeCTXsiOaYjK5dE8JW414f/Sl/lNG
PyZrUIK6dffW77pTLCk8ia8aPSQxgNpbvaFIWflUdhK/iE0mUZttWTJ7mARaKrKo
xSupyl5x24Hf1/l0Hhoqq2u7GLzwU/HqFnfI/YXlijl8RQfv9t1MRk7QN4xtswSW
33nqxiKXxXKonet3A8l+EkkIy4wVQtSRdgVaAxfb8KGcZgjvxXGXeBVq5W8NHWNS
mtHewmr3XTZvV73XNmZqDFqB94pTBrFjjeoHRBcpmUkoUBjjAl7F3L+fzuB9Y0qE
+rCY7faToZnRUT6mQBFqlwk3AdcWbqr7AG1pd3sB7JYr34FmVIsaF/xVg//iXeCK
TvanTrZB8MRo4J5h5ym16t3M5l+A0mJntdYVFsCwxCJQMdzfWT2bnvSCg5+O+57l
vmDwv4aMQ6Di084fMdvyfxUlOsR2q6sswe8O6XLZy1AbcAxsKo+VHvR78vmP7rgg
ZRtUqQlwFm+HKgQCBiBXNUgHEgK9dNov+M/A2hNYZlXMclciTnY/vsMo2Cke0fn5
9Iop1PoEe+TMrazPluw7wJwsPSOIN1/sS6i137uUXPr2huxOG8hbqDW2XK5mCVRK
mrG3IM23yUhq1ydrhazXzfFieqoDVr6YFOSojCcZvWppjt1rJyU1dt3gFPWT/mp/
BzGARcEBs3rIMx9zQ6aXGbsPvn1pGjUzD7q+qC6Ip5S7cfzXNE27wUl1vDIjIzUy
RNK24jMOsdBti7eViB+jjcJUzEsmyq698k939tA5zCgCeMRPRPAlQyVsBjNmGx4n
A+CxA4tMIKG1/fzGe0khSpauStgr+HXyFAT9VQQ7nEYQLTcmN+O5WOr5SIg4hS6c
Q9KkJ7RxeQHs6cw/iPcZrJvMe7jrnWMssjoVUve35C0KgoFFlsv+e/DQVLv2KFMj
OSNqseDW9IvHbjt8WczToPd+uF6S/+FKL2XUC7ALqfgUpGSvIguuqHvL9DOBJ6JV
eD7WhatHQ2Iu0om78ux0ai2ZahcAH4YkLqpNF9hKAh9jp7eZg+80tk78LkCa5Dwx
DKVhlyAANKp31xR085qs2yLjUSpTvpwrjqacWRK91C3ofhVXQc3THfzWAeeKAE0C
wL5Zj4vaeqpZWFv8rk52jIRGu8IY9lZKrY42WPNlk4TuWgW/rAbogdMUczieDpH5
RtWfmD+e0aYeLW4WhEs53YyAOQ+puaYMbAMmzffkWFrzrmYVDUOZK76+fBX5BMJS
kX7Do8dlFFiOtxeCGkpHhSXRjX4abXV3Jv7u/44unjUDfeGPRixag+/+463BuiOo
RAM1E8O1xGRVVgHTQ2HyyeclgMbGuqNuckV7jDPJkYjDMIhs3NGdBWzkE8wmzVpU
XfXjVN2syxp0uYV99F2wwre6Jkp0jkC5GLcB+auePXVsGy4eNB1kukv3a8O4EVtB
ouVi7f0v6ygQ/jm5kX1X4WJNWJjdBkl5RyzKhuurSn4Tlgtp8eVzUVr+8Zj9xZA6
iLWRkfdun7tNWeBPumy5sNvuQbcbgmp7X2TwQYgh5hzpdc5XRux3XpzzeJHtz8t/
+9IoSdeFIgqJvznOy83Yu9xDEFidSyFkNwCZDd616J9L9NpuDTJOLMAw3BKg4N8I
2tsbQ4nBsB0oGzbYGhFWaGxMJjbsR+fOC2lKXGL7WqpQY82W7TpthO4I9B/Tkj0Y
bRj6y6xh9QHxpD6JwCHYVsz1bH8sX9bC8DhVb5DsMEvwVkqIODZADbMKO++qKjBB
n9F+cqfEwpTTD/Ku7kOR0SOyxfNCPVN7H/Strm4D37vm4nsoboeH5K2udxl5qnJ6
6koFZ94KYxXs9x2Igt5PJhs3dRkdeDY/zm+SxHlARNOslwOvBjfdKC4MPW1+54H9
KBvHEK32hf4sN4HMnS199kEBR4zkSOhkx8LUEGcOV9dU998VOJJY44BLaKUNTYb/
uuYEWt/bpZCmCEPsbfwcCNQNYPPOX1yHeCEGaUBcjDbOqiAb24MNwYuzQgC+CgXF
5fDNzHUU7/D0WIP6H1PhBeyqB8dFl5xJCI5GkWv/WnTDaigT2r+BXjk8htLtiHN5
A2VEvCUuCXWeognX1W5w+UuCPHPGF75XISFUL3uDfgG0Ut/jtJwEiEt20Iul/RMS
urKSTUkwyyIqC1F7onMle4sTQNtLakKDN5ZpFROBPJnJrrPX8FDX5X5kdWBwieqU
Q23PrgbTmejw6b1k0nhWXPpVjV+Twx79b7mUiRjFiFZarCmdws5UN2/CPAe1FGge
zrFyVO5a2pt9YI2Kh0Dpgt41d6yAnxTfb/TnW4T+z0Y9YdvccfOPfUAv4kelSam3
7hAjdmDXWjhnmB/VKHezL/chYqiRaO/oGHxCIWtarIIvBlLXyWrU47BphLtIOB3P
ZGXMpYIG7Ru9n+OQz9rnkVVuyRI2aMxLsUc6pa6zXueI75Im7/UMFmEdvZ9s2oYg
iUzARooJVltZWxBwVmZCkjSE9OwPbW89ZT+oOb8AMS5BUCdPVatte8WNOY7WJgxh
TviVeJkbcKCgCm8Aw534McaiGUbQ9/bCKJ/NYexq8wgS7vFVS71oTc3nM4smrQu8
kE9Ft3PEd95usZKEaeWkxOTPqmOgqS2JNcztSbuejvVMVMH5P/i6zxu4ueOPYGHl
Vepjd4M9Fgn4CbeX3JXz6UUGViM6c297l4tcqep57/nad+RVeKzu4rQyxc8Z6d+U
Rx5GQo8GFiaKU/qahqPacMODVxy4maC7NClsNut54tYNt4zigKp2NS7gY5uZ9Vxl
qqZ+WHOvPjz+E8osK+r5qnC2el7e0ZaGjHI1mEI0fQws4Q+G/MsV4TVQKSKXO63g
es57R0QCscp32kImkSIoW0qi3nOcW59LHeAJkv7QmnfCxKXZV8G4z1tPOIENaqKZ
bakSTMCDVmWYOzKbJWwCmT/rdVMiuXT/EiB69DWjic9zB5T2Gwln+PxibpMkyMp0
3IFPi8PXY7phbLLUI+5Lr/nqZdoUymqvvYThxx2ydcAhFC7Gs5nMAi0Dty7g8LPm
M3fVYPfgXPtn6grrMj5Y/77LwxYfibDZqJnn+fCPDRHkD2u4b6c/OQ+3YHyW2Ht6
WvGuHdQNsJWzXKke1eeWlQxQYhS8KIN7F3+f3TSZHTi6EaweHMYZ5LtM6vhP/ETG
pGi+Vz1QECbKp6xTU6Dd6vRI1SbIu1BAHuowsSkw+f9MKQnfhgav0CxFYt2d/jwW
hCbn163hX8NQVGafZR+1L2AYAChlCVdb6OGj+YINYj6aiXFo22kZOoGH8/6PX1hI
NAe5V9PCnCIXnGQY7SXoZtCzq2znDdJuyEYtO2FH+82uUc/t+nQsmvVFJLsqZdzl
ONhhmCXlHWezY2i005i/TJxC8eI2JxTRAlPO+cCDzY+V/Kr8glkKicbv4H0UA+ny
STcqOZyHo11tXw8ZhUGr6xWqkIH9hBCm3Z6RMd0AhTATCK+GDUBCPCL/olE40q56
jyKTrOsf1h+Ti6XeEh1/Co+3yFvwqaJXUB5Q6QwR7L0P3stmEhD3pAwweMqm6tVp
2sembxqNX7J2Ty6AE6WZZpEdKXDkSiWLiHBSUGoQ7U95FeRkdstSvIW9nz5GVXLt
4yQSR8yYIELS4xG0et1JiegBS1fce4iOmuc5pOrFNoD7nGbDt6BdTgHIFPWyHzgg
Zx+DSJl7HJ4RmI7ugQy9pZ4oGefb8YJUeAbem9p+Dk9JAXpA8v2XFOFxBZ2uU6uV
rcZLGluyKuYQKhQw012/CYAXcyPnqypSSTRq58ZlAyOe3JgAA5HylQ7iCmzdrPwn
C/GlB6Lrqg/RexKib0Oete+slR44NzJQuoe0NS5YhV/Gu1TmbnYryfNwRsgtC5bp
6tpyf9mnlI3npTB86QgPoRFAwrVPwTC1hrKuT3WEy1TD19KdXtiRrfy0lLMy+2/j
xVH2Za1BRARPWsxMGzxyuRr1sqbD3as54ef9hBQMRE15L0CwCaGu5lgKYOaw+wTA
WBbnSxpcDvSsAct9U/THnB5AsXudTRq3kJLOObTRCONjT/EgA662A1IpUGdjCukm
YHZb9PNrHj11hUTMfal8o+Hn2ZVmWEBhUmQmrq6MU5EI1cgzgcF0cEgIMsTkyXq2
XO0eNJeUGIuGNQyXm5DhNfM5xL7o/AobBAlEK3foEamGsAgyrDOGq4SjRiSc/w+H
BU0BJdaFFdmzmFcTWTlzuWWlkpUo/4Rf1KJncEy+N/HV8hTfgYmk6EjhVfS5Vk9i
9G69W74gSNB0skJeIYAqotqa1GiRGu+zld29F1MsA7coLmfXgS5n2W7UGbm4yemp
p3s/js4h3vnt8f0A+Ke3HfWVJ9lzznhMkh6oyzdBNayCXVIgc4Sn9jxeOTunBQjK
DmPGAVgu6JegyFYkUZacY+AbtyxVwQsIWTdhHWuyu1nH9BC7DcToADAiOiojOkrW
LuCgmM7Lzy5valxAEn7s8o5h9etIxjFMzVd0/ykDOH4nZHrqXYxkpVOrCLn9PmFg
05IrPbFu++nyIfAWPX924Rxe2s96T9pb/OlQQpeUe6GfzsYpipfeFjqnHZYEqco+
LRtd4DfTvhkAf0SuLXzguEXcEx5xIHeGrdlZ85liOk1JmG1lkqkUwQzAIPYNh6Jm
7Lzx1h2iF2mareaKrMNjXCpGw31rAoGYAi3CSeh1L8daQTpLosOaktxdf+vqbtR6
temdcTPD6b4jWJLeVsxMn1Zhv3sGrAyOJ7o7FtSxR7TWxX4ynxCXiMh88EQOppiT
tmITunphgLvJa2nzI6g1z0HPCW/IDBfRWNuFfeJXRv6cXgFyVv7uzr3YPUSwoY1C
1I4eThK2fl37va0W1olgF/zWS43REeopKCBSyehZA8bELMIX3UuRSFwVtQy91cin
jwryuDQ2XFt3yx5VjuXzJ7IowP1/p4IP6jgTX2czAqo937Et08ZcwQx5Cl9+xf8s
HvGfRUsJCfJ62P1drVd4OiqyTAEZM2gFOBKgJhKlQvQMqFoA8cnNTeR1ECqAh6BJ
DgrZzSRJZdeGka9GhmRQZYD7E1uLIck6FqoYHLkpOZw6wdLB0R359bZRSyuf/ix+
ujf2G7XlciiN8NMSYU9uFe+Hteghq/Wf1UTLUzlWV8aqjtRxxHkDU9r1wJAD4n11
H4zqwJXiGWeefhr5VC4imXJpfLG2RNozXZwPtQbqhtCTKGw6pT/P8CVAdiKtQmna
q2ETu6IOCdFvYKKfq7NDYbjGLhxptAduKjHLg9qy6HSbX29C/zvGkmD8NGqjry6b
sgDQ390TnqIqwEQbJ+QGzFt5OW19d/YvvNDGubtamaYYvH7Uy14K9dHlLL9Gd+59
zn9ebY0zi+6rosZOky3m7oWJ2hNEyRv5zv/Qfkb4rcpF1lfyiYoeUZNYPqV8QtyH
6FZ9+x3oe9Zg0SZTaL03NtLVXVS5nff8GvoH/7AReDUIurf53lNodJpKfsdjYWdw
A+sxsRUxg4RN6Rg6j39B6aiyUFImR5xnwqCcYBH141bMg1d4L09lFV2MywBIkzay
xsqKpl0n7xvuQKSuFWWTiKzwzn44huciwu2RO8GjnUphLoKGjNZ8ycIUWjKqTv63
6ppMiBFAnNoh7BQxoy0SeMpMgaXA4VWxhzDbek1o2nWgUmFNlsPVujlE4UXREO54
P6qJjtb+QTjB2coxlyvccCueu5Mt+5AiyrdKa+azOiVx/N9m+X2XdmEUmSwT6Plj
Wj/OB9IGWj0tUZVowmy2PTmwAfv41DgMQOCj9kXr0lRoawlIz2/n+jdO9exRuyCM
5lzyFkQZGkLYMJUb+xA8IFJQwDkVsEfVgKKxUP4bUv5fe1lIpaWnweZr/pIVdRGd
qUT8xWj4FNWGe2DesKIAfZm0skKopR3y+Fckk8byRlRme1DPB80QnuC94ydqQEeg
ARday2PCVr0KCkeIpwOUGtDtJ2W7WaU8Wjb1yiNXvanIUygo8X5M7EIUA1f9sgkV
+sNQyMQPd00v3XhmcRnVDg9eOTkYhzjP8vo8CTRqZCtaN6T/2ER5NHAoUkercVSp
jrOO/4UVk7p1mAlDSLeKXX5/QVDgGK5qRrxXJavCRauP+9mh94Tho//lPjnXSznx
RE60bySVbOwczWY+yVt73RzUIVtIxcTdm55WvMFQXyHosZKurWbtvcbtQfjUOoR8
sQjb9WHEQeOg/+8vwFVA62Dv/0eIXhgScHkNXe+HUt5Z8KBKIJ31aZnsstYNmVmH
uLoJD/5Jjqcbptwm7ddSTdxvQ6ng18OsHccLfI39pkZ3mfSLpinsEQ4GvloM0EVK
ndIWktx9VItXjXtkyeU7pkJ9Ok9rjWLX9lZX3gemN5vVloOpMuWnQwOJu6hmrfxn
9enT2H+enjW1+3QobNOPJoxKfa+eouG16aQ24fzzpkQuNhjnQJwIAuhN054oRqZS
7xX6i/fvIXQC2qVcEQU6pq2gdKjZA/TC9tdmgvmzZ5l0umW+yedSh9tVJJEf4PvB
ToqiNCrS9J57hJ0LD6TNbahil4FsgYzB9d+U5p3VJSPThL55ySlF8qmooO6r3YzZ
MbJ6ECEzVrwoh36/ZkWjfmSrt9ZOBmU9DhILYnmLxfDMBZDEUH7DTLBQU4h80TBR
wcft1MoDBZYRzqGltMNg3icHYi2nSZOxWU+2/5Q4JQueFtlT6cdbsIx2gher8ijj
eJOig1brck/Mns4ZTfziG8BTvdWBMdswLbC1e/u2U1S8DgFrAf64uQ0pbK3Heba4
QwM8otC8wSYH9BHSlh8hLVswADRToy37ASlg4bF/MeMF8j2BPn8GZFxkMggkvDC3
IVXneiDcuoNiEIFY3YjpygohLI6SxiArHbeQLbGshl0yaOCsXjEszh6HPtu7cRx9
f4IZIqatPvWF0BSKA7Y7FFykcbiVw4LbgkKSZ+Chp8LMl9vRaKIy/SjACWT36wfS
decregeK2ppc3vslStamOOYJl2Ce/1UKA4/E8VDjAbOXLFtPVFX3ameEsEPPowWw
3y55Tbin/qFvZsPEZIJZLtCUGtPwkiT93QhK5+V9DfmogCcbJ8kKfxU7BB9iZmpP
z0VPwB5Max5hM8aDGqt7nu5oTvjevb0OW9icSDtmtdzdLjpFJzdQVFeDF4wf32hO
rpSSx53494QfHuP+VRPUeqd5FpYQHahprSlRgCnq72akFXzAvaJ+eG0Rf4VMGUDs
68HKGFGD0qSCmzLvLDx9Nz7qc3dXlMIS5n+lc1vji4lmio5Ow6tBQMXTCTxrmxBX
GdCepRKLMkTmnBPXgk7EbBXCfbJ2L3KHmuEGBs1uvSAk6upWQAkwVV0PkVGe/LjH
+5ueRqoR7+opUvCLmiZrC0wauXDOUuOlt0hkjRTlqR6RkycH1mYxPntlm/fv5ClN
lSsbcxSCDImQ0NxLv8muuaCyCzzV98QMTbr6K6GqfdkeuwLElDqolhWyKDvaRdz3
Nx2hiWjFL6oFSZa9rAnz8JHBR8aKmt+WY4bsAzsHxCCXpkmVylTDhobvhsitjUq8
q8UjC+TmclWc9nyImfdLS4MlbonkGl5Ss2CCnIAQ9T2OZvp4pEmX8sdjmX7wSWH3
r4IPQ3BEeBy0PWZDEoPMfG54+ivzLbNIeMlwYYVBv5ZzFEPg6sEm8a5RvsJHQC2V
8Cnz5rhHz7nIMbcFWz20ECE5qMJ51TWlMsrxaQjzbbloft0m5+D70IfcUHdQIDKe
166mJWumRwXw20US0azAgDXBcLhbDnvzjSzIfB6nMRV+5TP6UcNrfpKowOWBbDni
C7CnU1hf+wH1m9Lzcicr1Gj46nW1NJ5aTZAdyzMXVCChK3K4OeKp0xzjE3qaSyR6
yv/GYBkStD3ilDHTRSYwFFXZd1/xFNaqoadOZ+LaVMKiwFTNaQ3E2geyhAqOalc8
LgjsV7t8SpFeM4PPRVpn4iyVncEbSx54e7S+KXasi5tLreKYrvg9kUQwu9KABV2f
QvgHw8jm5w9Ooj9EJqY+nmtyyJB2NhN8V0VVtz49k5ksZ2wiDZyRKhlSU/lMIJUA
xr/KPQr0jqxq/Hm2q4vbUxvZ90sGOJIQ9Ju3PdiNfPZe0EQPd4Jpc2HJ1Y3eeTQG
MXKbdwsn/W0Df2T0/OurLALpzlst+ojuWfByqL3tte00n42A+J8HD8kizB2HQfKD
h5B2LX5GKGuTKyZtTtlOz1ILGMSrJ7ZIu78v/kqTFnlWHeEbNa3b89tRkhk3avi6
ov740Dc+DHroRxQFxsyl22yVpyy1teoNQRFtj1/vlIDCteR6aTT4K9QA4Cy+Bq4l
VBHM/TVH/1LFlm2DIPey7UqoUmhrtWGOECAosIlNlpAcXUoC9W/v83GTB95+GWL9
XRjvpK2HccXZAt6LlYJ7cEMRjMeiFcRSd6atqkKezvtyXYZo9M2hoKhjMbotCq7C
Kum8t8RmWAap/Yq2+mz0kbBo14B8dIkJukEDk8/M6tboIAZSgLydqXTNtsFAE/jI
YN3VH617ObRI6qIZpqNa31YEUDYwaDiH1ARr9b/n8jFP1tw80UQjkGQjXGM9eRiv
LWCri2wfPRxNDUJhjk70tDAjL3i9GQef4+ZoFX9pI7RI6tw1LGjwTvctgOuODZqP
cyERUUKaVIb0pnDf+pXO5+DkgMi2QXB/YcT7irS4yTTgDi28n5cnWCiG4oc7s709
SGqwHkOmn2UZCBwx0VKoZjqT0jsR3RE0jfm9fgX6Kp9yNz5l6PWQgOKRrvjR/iK+
MhA94I6AvqzfNFRE55G15BP+8w551KvzBlBU7fP27nYhgxjX6+G5UFrzRceid2uG
bCKQ+1bDCHdw6WbQhyC3K0e16AjISwrotTZP0wr6IrD5JCe1rJvCuzAFaajytanr
gZouT2fOBC/KRjtOBs/HCLZUuw9aUgpRj7lRqP2O2x4zziP0qcjWsiwprGMDDeSG
hmL4EJNQa43UDEDUj97OUt0WRLfOadOMuoZoz+aBdUQtyCCLm69hL/1q1BdfsCy/
flyGF+fLexnKIiGDOS3oUVgbB6HAFXpHgm2I0FAnSzgy1Qnz6mGhBT/3l0PISeFi
1Zyftv7CEecrw/BNKFtAEXL0FbAgq4OZextINbipPm/IfGxKNS4CiEdPY0xTQ0Q4
SMs21a94DXMeZSBKEaYMsbDB0lfNnwlkxNiaIzbsNFMevONy4eMJN77z1eqmo7XT
P+xI1Qbqg48W7wV1dh+xyW7dyZAHiCeiS/GyOTCLByf6aFEwVVXvbWM14RJt6vp8
/+cJ1nEYUajudokjIT4ErA/DepINb7URPkcUsq3/YMsBlLjqlIsjduWQyZtApRtH
uMICJyjDhl9UemQDPJnKdpzflS4oOskpJAzc0JbXV2uKeYFcyUFcJYU72BJteHwU
pit21MW+MbeL7xbGx4EI9uQ0ZjEXPZwIYRPn93NX6A2B2Da6zzsUWlaSttGQAgHl
4KpIWbsIMMuKlOEf9cAqgmXa6XImimbWpGvpVNF3ynxQL8ysWWu+taMd9uZdpMJq
7fO3qGb9IFopViT0/tsd4dWQvq33OnKTCjhh7B3wbkYOt6riZc/kIGTyqml3hB8V
xAb49leU7OMTdLV6cvNzyP6X3KJWvzR4e8mEAFoz6p98OPi/l3Vy+mZQNZRbp5Po
lagkIMQyp8qHubUbiVBa1i0lk7XwQ82juzAsJdvGD0XniDwFxQnVD5/R3LwPntmt
KASFgdu6dN/J5gjZlL7GAvocCpvIy1aTC1aVTyxSF2FZnIjJQq7SXM5WLNK4a3wT
iOtBaTwnoGHyCRbf6ZUM76SOAFTbJ/Q0WK6n5jVvURj4A0/MotBcd8A/ogu9VdIh
0Uupmw9EON4/aA0rETf4uDiXBRW5Q0he7ApSmopLts9cIEnDZIHToupwygnu2nQl
q6mfH6WQzqVRA9b5LmPA3pxnHTtAnlSdktBGFLxPETbWTYEXI6j+luXu4vurKZEv
5vSVgcmN8DpsNq71ZRmkxFegIyoLYcXvkq/95dDU2j5xInZez66pE9tFpt9Kmv5/
8qsiPZ/NYQ3tviXVfkM5aXwjtbgpe3+K6yPLFkirO5i8NyS5S+8pO74WHBqGLcna
y5isw7t01BauDN5B4JUq47x95D0MzQ8pTk1SDze8+Jvv79JG4Xi8ftC4apFuxnPI
QvwB0ZcIrnNQadOxI6fRh5PiBdh9niKfj5Di960HCLslwZKCcFWGCv/X/tBDIIfA
wwdwRCT1wXbbDYnbbXKG/slZlVXLdpFrTPEs+iU48dTg+uRtVnX3bPyWh+roKcsp
LPonwUBrKqXKuMsMMyUPW7xa30tUfnyDUhGoUhK85EWBok+8SS8Kfl5e8AsNeG73
CEUoBnPsoHwO4zHOFxG+0GVqkmASAH6VqvCtr3CsRWxU8KdPzpP5K1KBU+IGFROb
L/CkntjQxZJmgh8CpVojXWc6zu3sY/0bjShaMxhfBHGeZ5Xd7xqoqFyHYxv38ukk
z/McHz2nM76fBZjs6Wioi80ADjjlhRHxFWR4ceErsCRwtb/BzGCGCz8uITQmOo7g
rC0qJpJ6vXSP07U/pokk2ynNjcc4T9CEZDyxJyTZz4asCnRO5n+fYbcdiZkyiLcL
aribWUuDiQBBqOjCovTIB4d4usrd0mhG0m+4jW8C2kRU3g+hA/Ky2en3v5VuiD6k
vKw2/KWhjt+HUrHWkYMWR3K62Ua+nrJfk2RTJBWMJ5pr/h7Z11j+RTFqQPebIVlk
eQJoNwwZPlw1hsO6+wbFh5DRhXT35jUcpyWxzzvepvnD3IDKfXtA140kzI5+yCsF
2BVZR0PNXYxtwjhHEMWUe+vRSNa3zNIjdhV5UkLEhuaEBJwjGV9duL68+uVB19it
K2yBdvk83F5/nLOKxtxwqCMTbnM2GwvQ/X+rdGEhocKQyzut1Gv+XGUC600HrCQD
upPYsJ8CAkql1qwq1IyVzfl4FT92Jmp7Bd4xewuLU69DpgkyFbfptOV1sCkXSExW
MHS+QbgBkOdpBAFnh18x7ZNVEKPQsFTcMXi22FaD70RxKfqlch730rJvEKP3Piqi
CQd13jlYU5SMG/wpjwZcZs9cfa6KdhOFcAztGQKYIPSTRNmgY8ddFOgRGmmBaF4R
eAkmEvO1qy3Xv1HyYVZBEJ6pTkmReU9K3R2QnFhBt1w9Ch6nu2JOOIlcmjLx3asj
1/jm7mF6dB0UrO50eO5cE1Ia/G6K6O/vZO5hJ3MOFf+AykB6gU0f74gsBpu254dw
tD4yH8mbk/EsMg8Uyl/I8UTxtY3IPeIpeaBqEh/3itq6Ue2P35GJaNKA5A3p/dRr
6LCpDFHOQAeGd2Cb8YlkzJyhOJM3DiAw/uI7wnV+e5wlWb8q+uN+tzinadPshZkT
FCrTgteRhwY+RGaZs0wGyTB5RAfaRd+dyB3NNXax1c4cEdLTtodUlRI7FKgGbpuR
uYkIulA/8imzT12rkPfUQoZ9o5im73lGgMYMPXVvSVPFtsKbMnOxUzHd8Etp60AW
D6pFY6TmJpCUvNv4n3kG+Uboh2nkJcpBnCcK/peqBVtrefoLcDrnKEQxdRcBmapu
yGI0kd487LRPmFivtw1dIuBvQEFY/ORpcMUaIJUW/IFY/qUK90BLo+3MfSCLvmzF
7P0QpHyISdOjLXa44ouYVCFB5ZfgQPyNF9A5y9xSVjcXr203aJKuHB7wl9kuQT6p
qHumRxu06XwTaOYm4/L+gKLCFOvb1Guaiy37VzqXVBTfEkikrsuv8InJdqs/g4h1
3ae221eT5WM8p6YKZfSztNYq6atHQOFLSHbTgQ0UALHuM+dEz3No8cXdzHxLG4UD
KE84VfPE42TS1hAr3EOUg100RrDAOmDlH/NAYGlcVXBq9jZuVdcp0jv5Q/OM0FQ7
+Y+u5Ip0VAG9YuDhIvCkm16P7XV5hbspQXlXyWscbiQ0zSU+I6zPdoTlqi56UMGl
XI3Nu+svCnkCcz2wZutbuSSTmKADRqB86H37KidTCJXIbWZn8aBLYc46HbCQOr3R
Ul/l4AMcFnKxCYsXGHEvpOJ8XqiUifHilufWb0OCyPBR4i7LUUPw0c0Jr8jzdOBj
Q23skY8PdVJwbHxIjF2aGnzXeIUD0hF4dGmHc+5JLPq3kpZLGqSCN4cvL7vK9E6v
6D6r9GTMfXiaAKd5k5fywMy9pJEYbyLrV2kQCSsyScPuotR7UIS28aG+DyPQlHqQ
ZUXdv18tlbhjo6SDC83TND79YbLssrLZgzyZCxz+3ZjwDD+7N67M7bGu2BouFFhl
afSaBRINsZmKV8SrQ2E3FTch6blbwmIp6fEWNKlMWOBh8lYghWJGyhAFHzSGrJkj
GdjjBVkzPtISXspUIWxxcu9fm97aRw1fiwvmO9VnS2WX9aem+i8HqB/9zShPX7pY
qM8/2e96PTOJsgLPAoqfotQoZAsEHyd0/P3ZNwN6oQL2iWwlzwgdl8VfQNAP6bH5
EU2mgAAeKzqDqkGjMjQr5RO1OyBbm+Dm8TO+wAIEC/XaYszwkByxl9pcZk14UiQj
T8T2IDV1+1Spz1tI6bmPQ1yvERTLsgc1sPW+xThsmGsR8P3e4NIYRnGTG9YfEl/n
xuXIHrwn2Pmjdx0TqUp8YfaFgj0uPouFWCkKf3ViRzakiqXti1pGYEAx6pomDHiT
JI7ftU8dIfRe9Na5sxdmMI5PfIFzXC/AUlN7JD8OtXt5EIAXVfz73nXcVKK55iH/
KMqOBcRDAc1wyDsISLOU0CyF0prtLwr9FzmFK76KHy2f2QS+M59rhvytbVMyx3jU
PniVJ6f+7KVVJNEC30LgHhYwO9jNtcVONTy5biHC8cPpozMhFJ0WcP/XwEgGLE6a
4cOl0m/XA/FLN3uWA3PfXr6/ZjV+bJTBZ9yQmWUTlN3TUDIE9vaLLTZfPWWctyrY
lqWBuYf94seoJ2itgBl5UvM3/FgEUqTMGRpSFZu+IFS4hAn076MtKwDpzoNsJMZm
IBB8BI3iEI85YZ5iBIAmVGtUNqkkl1de3Oo0CS3y8ChKwRQFXnoxLQU2bknde5pJ
kRXbi8ChDGQwy/Sztp7GCwI5aYNVI8mw2r9Ov3t14bhw+cCgRAmnAEb/8xRKjrK9
dVqJbsAJ/bTlebKF9bHzJRduFqFGlPStYE8hvOHBDGmSRczgpZ4D9r75hZIIlP8c
Us58rzppcxz7Wx9xr4O+qijwnXdbQfKJvugkLclO9f49UHGjdvxkgMd5X2aKmuyF
pK7MkeTRNQ6MVQXD3CzHSBRtfSdrpfyn+Kj2WbE27jpd9cpsKxQ4u8RfDnL4Tv+a
tpdQLZ1vWnN5NnvhWV7g5QEhd+ReWeI6RY88tJYpaGgSOm2n6X6GPauaAen9UKqE
N+M+gJ87vFEsR4Ljx7qFDUEaH+/TzT/hwbUJSaXFbVPLahxIpOfKF96aMSLkSzgh
Sb4cxhkbc1Z1zqkAUIUX3BItz/dseForVYbEEa/kKUkQzB58A+OAhitE0v/2Tuyn
przQf9etWwrNqTFWLZovfUVT3ToqoU8uDuSkvhYvdlLLZAO6wCZqrbiNmMb4abLB
C7hcj+I3e3HHYLZEdbrw4epiBCC5iUl+UtOSzxEwZ52d9xiWbMc9bA7lkNjrXzsX
dgSB1Sny05GeG8NFHKfmQ+0FYSFvAxNYOAeZ+9BgAPPykxfxfP9xPpLA/zdgYYo3
LGGH42RL0YIZIxkRgic0ivQe812hTAb3W4OKvVj1RP0hxObXUm0+OoNp8mluxuz0
GUeWR4SLvSCYpx3xWzW0ok31D+bIN86emEb/MoKnwKpQNyCv1qOdobkjXbuiH09d
46iujXexqY5z4KSG84mKS4hDqnQcdVqdtTzXCoZ0LyQU9Kw4Y1DYuoMP/n6AcVoS
5DSrQGCxivA1OV2rpWShZCv2T5us4a+2wvccIED8I1g92ZRYlhHjXtwcYJqZ2hdr
pMwVPzZFNSRUXxyBX/K1jNkUKx+uQiF1dIBGHv4LrEMT6/hBXXIZqhxTC2oBKdhN
dgiTQ+pS/d9LcnnEIWDgsYc5j0WYPcrblyGeDGEfeRCFfxTYL45xJWgtqBc5tPbZ
f60rxnxXNR2FVwYZRv2O0UYs2VQxLXtaFrsIBaJFwaaRP9JJHB4picW23D+Z/uwL
AwlrW1M/EQHWkwUXTU5pZlckvFp0qbG8d2SLPShe20ZfgOcKLgiZaz/qkFyFZ+5K
BRSSxqoRQvfMEXLopbesdseBh31qLO5TPoN25DjWsn2jsKWysOlNyEYbcsKJgub/
F6SH8kAjjn31CSQsuvMWCwM+dXMWVj/CouIvCm0SB0a5T9m5/yMflKJMjgpwjKoK
ap4T7DcMUWbBltHzIRrKD4/4I97PiKPdByl5Utpc+ddVPe70Wm/BjiI9p2G7qt0B
oWQJkMI5VTTSgsX+A6cYzsONal+0YuD9rCWTcQFwGhymc2jtto+F0nOBeiNaX85p
YK9eZRiaOMKYZmebDMT3Y6dlE8eTTO5Hb3mpcIFyAoDKKix9qpRAQgB6qiTy/UX2
YJ76wRAUuL4QlRlcBHgc2P+XSrEyMC3UUnQYjrIhcFJX0Gx3xDYrKc17R3s0iL/m
1/BhSUS4lgILFl6iUkstEkKZTUBl3h7Uk4DbCkx7tuXcbsSd39Kr9CIgd4+v0gQC
deEjodQI7q1xjrjNQMmvylTHqU0eJJlqtPu1h/6SOESIJMLo46T8ROuor1PtDipv
TotaJjzfGeOVSwqHYCi9WtfFhT9XH0hr/FCbhi08spRng7y7wxJLzenYz7lWakVx
+vqfns7uTqTDDJDFzIaZdC1Or1319TX1KYI369Q4bnF1SVtGSMrTd6SboiJoRt+q
rRjbQ0if3k6/fSJTb+UO1j6mKpq2rFSeCKTBuLIhdjRGzgaSHq9od8glBMjwgwg+
+wPSdOxWfpma77qCQ2JW+tJHn5+wFver2PmFwFW9oSuUDHjBgbFMZpCYD6GI80b7
MjOmUKppFWAEyco1rACnd7r6xIdwPGNyOsoMEyYLeqji4Gw7e/Bw5FQ40mkxY9fE
Oc4wdakypJprdy2F9nwc1R6FdIyl6RIIkGdmU4cdKWYQ48YPipRHOaRUsATqMX1q
FTme8vwBRib59L0xNBEHjWjn3l6lf94/IhLU58aH3SiTz6Edn2SO8WLT+RdRSSnd
w368N4JGVoKN523ww0qTMzDPmXmr0UatGET2tWkp1BNLuI6CSRBCQjMy5gtGVnjx
1wViXFizrpWneDGmna5UYmlosuRdKAsebwMVxisoJovpS2+PTu0VusL7JHZBRx6P
f/ZMmKTAZsJaFYLbkO98j85jQwXYxCd07wI2JnLapHyxU8lokJSvCt7Psz9xckNw
fBhi5WOG74My96inEeI9yeLYRIEVMXfWaByxipXMrktT1wrwRhf77xmL07IB4ftP
qDgbqFd02RDokii4HI8aoYkuJuHHTQmBe75vsAGtG5BUJ+Now48OxCKLYhoHwfRc
HPnjLkGU2Xd+zChoAk6THS6nfrVclfJars3KyvDi2zAeHXSwXG/GB7Y4dbW2FKwu
YTK/AOVHm84Zewp9+WroX2sQfTAvyMQdgl1/w93H40OLTehgsrOoUMc1oODXQLN3
MS3Fcsu/GAbrZGL4s7m6FNaCcDd23SBZwG8iQlbtrqbM3y0xnUeyCfu22iTmBUIu
UAo62OC4EExXScQBmktAtQUhNKQYtokYVVgmbb440TTyR8I9jIj3suJqMrr0LbiJ
Ztg0aEJmW8SJ5RvxPoG6iMkjxYp9PgUW9+oSa4M1QmlO1wZRPmWJw14PMQmRiT81
GGuw3ATRS+uaNV96THcDHLgZERwV49thAyUaYzEMiwb0Xf/6UGr+FK0QmlyWRUCm
9YcXN8+kVPEfaYT+gHk9B2B8tYyU4g2HFLnZ3828dyvjuiWKkBl3wbDVfPT5R9TT
CusDfZhHxgzsZo/iM2lMfW/f0+0Hi02g55nwGvrnGkSVZxKtgGtVUKfaoRggP52z
988WBVsJTh+nJ91V788rL5MOQxJYNwBlDodwvz1hqCRQsIcbyg4GZRPYKjFIyOec
U/U+tDInR5Wmj7aY/uC/T2zcBtuJY3OHfBz8Pll3vxT6z2lBtql+rkzSUc/w3f65
SQstpNYHEKXf0Ip/oD9CO41WqZGXZOWISCeb3LvmFWigCq6e9qlgAMT4rdgQIhO5
ZRnysLVJ2jifIV6P8Oa8OCRcg0WUr0WNv/2OooMtU4qolrJpbNU+y4dTeflKWMbq
W3wHZxff6jutAnrSYG6jILovqeTxPkvZEXkcXyQQ4ZQlzvSCn1slb0XwYfdWyxJj
O7l7PJ+SyFfOeyoinKc7hNSZUpSObpZpGqPDP93h1DpXqoVC2MVpq2Kv41Z/hIbA
g4h+B5jEsoRf8UjPnvNB6XXvHy+Ha0dP1ZYtyfUd6rfjpjMgOxLVOfuuJUup+Mdn
Y4Ln914k7mp/rJT5eS4AB4qze3bScorf2/yY83AX8qYRGR0sws4JPiSnAmWJx8nS
bwgaR9B0gT9J7+FjcrzHiLisJxXr0oqEALCv7mOYzNkMxNc+cm5Qd/ZysWouDyYl
yrT1kkxraPYEGNXSOD4xF2HPGT7QIFW+Q7QasU111W90A+9oCBeT4m46D5uJQkkg
X2g9kFgFl1usJVlEqqAaP9CZZESuRpDA8H0pevgZC/DE7EDri6maC/bj3Ss9vaDM
nZY0jaMZc64k3KFpEYQ1IvpKsdMphx6O/uOozOtwA+YlEc1BfO4kgurG0iiKJdUS
fcFwriVMC/NnxnjLOZL5AT74bNvUOTcp2Xkp5KieAj5ZTeasUM93tZCM6fS8rgZv
YGU0n0G00Er1XK4ZJ55jluZOTMrqWYQpy3UkDDKypnlHFzWYYFos+6P45tTLLf+P
nCDPXGmbxTcNBwO/Grw5avsmTIVAPM+cgiYA2tKbZt22wr9OJz5UtrHuYHiNWok/
04H7+2n7h2kkHSLxt1sizxviqPPto3aqmZbf+TTzYgX7Tn4YfkFY4BxymnImRdkI
fE2Qld8y70uOSaeRwmSBxcQ0E7FA39EucYjMD3M7IKOyg5Sioj++VCk/CVKCytkj
Q2mnOxhVJKFEdXKioE4aZX8uB0naLnZrPKF7FX5eIapPlwvkHHg8n1oNWGY6/4qO
t0bqkvnaQKk2axQyd7+P1Bvf3N+lUmNZmzzM8TzbHKyRZLjWeRCMYfcSONoDPf5B
iNl5IrE3DnF+Qi4R5aJCcnIeqx9J7a23572YWIHN0GJp0L3V0JYy8pD3jiXmwMvz
q3iTJfhGTqF03KCvAtC3yRRdiPvSmAoJjWjXcNTqAWek4Q31Z97vsCj5mXV9HIPS
VKwLQF4MDGuu+nSfdxONOLqWkrzCNfaShToZqjUdBiAY4BfVhibUSsoVlAiFQ7++
UQBR5i/CLiKDQMhCNxkEgLm8HcsQT/wC0DVohxuXABf5MGmIJDtjebUJgJIrLvEa
UBa1LSwIW9QiKI5tXm+lnfdAy9Y94nmje2c7yTyjhM87eV3oExnfj/ZXj1VGcs0E
jlAWmy8v8x0o7XPj7yYYXhARyDNm+AgTqFfsJoyzT8mSrXzUksUqJ4T27CJC12jT
aTm1HLzg6NaanTmAn4TW6hZrJ2xsnwZPTbk767/AFflB2gIsBXKrf8/AzGKpf89V
QzJVaOXRBHiTXN5SqcJEDvF7namJTCHqpLeRDIv3x5MCyopODG0frhQeQfj7V640
JxChQEY2QH0zivyM4c+1jAWAUByq1alCk+NROEFTdUvSF4AwCHefTIdLAyB2wuRz
iPKX8pxPyO48F4MvgTKVaeVVTzIYdXULhYz5DGWbtVtN5GZ3bLfPOw0LPvWJt0Wb
dheP5Eleszgli0E855iqow+LG0xZxL2v8x/WZnfxaEQtEUcRjxDr3t/fB0aV2CMw
J6/AoCdzCY3u1J4wIjgRpj1uJO0Xx0rV9in7x5uMPLqucCj97dxEw/qKjXy8GKQf
ArgMooxqkPVuhBKMdX7CXHdQ7RVj8NaWQ1lk2Blo4EAYDW6m1VtKwpFqJA/DEHZA
9J0j+9Y95yUDSvRPoRDUh7JICz8plS/nvPXyiqDUYid2Ud7USOowxeUGOSvQIztM
oSJgpOVizxq1Pdyp9AO3Y5sxR5EPGmBXIkJIuDfdFM9ZDbVMD/iBAMrt/CXvWcrW
+aVqfA6xh56zvC1sWrFuyyrE4S38QQr4B3M8kIGBaDlTu0esTIAy+7FOTlJaeq2x
sfKjxLALGik87ExWd/uG8xS90+rVU77aXq5cgnFXLEuL+ji9kQhxvMkm8uvcuPR+
qPYKK4qwp4YrAYkN0+CfyDlfFLlQwjCDozmpdvSG0/31kwGtpSpTirCi6EyO4Sjm
0gZ+ufXOWSsxqLBo0lbJ4fF5e5N8jPV35U2RGZ2/vs7DtnFUAklulidjVZKz2wKi
ln4g0Lw3UT8BCZYTKooqMy9N9o0Vi6b1oRtX9uYOaAAszhQ9KdV8Iq/2Om9e/GTb
mdsHpFVd+x9O6R5lYtg5l66+UBOA5V+BcnOmHwe4kP0ACRQWKLUOI08XthKbsKtX
VIRUI+2k4sP7qG2ql2AR19w3H6S6RihNTMGWwvhrbY9JJt9ThPO7xBwncFK/Sx4a
OB0JdwTXDDHARVg8WSHzaWAmncr7dOh5L7ZpNCSHGXA=
`protect END_PROTECTED