-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Lf9EmA9CB3m4iakzAR2KJw117YjYZgtmzi/jzyJpbovbsZ2uIPtxh8cSLaiQVBGPanlyl3WkP6OM
U6b47+BFTsaG1nyy3NvkvSjxaIXE1tI/2k+8i184RaUtOfvtLu2ax/ZpBtC4qPAVTsc/MVDtKlir
J2jNZ/2upvm2B6vhjyOn4s6Df1V7k16Zrd0AOkAr/BtoplsoHCdbExVgbJoKbVDV/II7HD/FgZuo
lu933fftgYoMen+Y5A1REQuoXNvzYbbKdD5fnVdXWJuJaokTq3WrwSIEiTKZGsJdcF62bWOf1MRF
5p5M04QBJL80pz32qtx3UWcMTL/ZxmBQiDMgMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 116336)
`protect data_block
DMRWlphwEyFQv3PadizfnkYOu24yKHXJbofNZrZbJyqn2ZQyY/dI2HvCOAo4NFEtibH58Da34qe4
It+Az9o+rnJ9shzPXN5LrgsJyFXiyklTH+nfpAp0QTltblSEB2p/hAnJAbPxsjp1McoxhxZxQnqF
9WzzaIfKIDeFEWy1sdcHeUOX4K49AJUt9ndM9c8LCXdWKs0M7p1nbUz13VWBi8JzgT6dcvzvRRS3
lL9eEhD/lxH/bqX0L1uXzyrj/oBMBl5EmJgW/H8V6XWaHnWTGy1+xwiKACngqbqZgUGUvDWsvslC
MqK0Ani969Q+VtLkqQpLWULAJqKjX2Uo4AqkUtmm0JGCxcp5ZOFVP8XNHWB33pHZuQg+4mazNITL
5biNpS5p2GdH96qufJJIlB0KT/1Qp8Nh0Y24ndnW6ppNGgQkj2qzxXRAJ3fpeoq5r+rViNPWTt01
v39E8VnYuxsUrX8eRjekQpuUlCGrRLan9Y4LGhG+Q2AisG2ohr4F9xaRDQ1mgkhWR9wzlL65bXH5
E1eGkNNkpHwMlUiA/Smaqyr2Epe/og59+17wbDfAdNJTZ4kzZHiFCdqCkURl5ic/48bzx6Iazv2i
xV3c5kcPP+AJeuWf7Vjj20zAXKnNJFr6JAkfRBfhyfVkZqIQZsnh8ScjvyRVhs3qvRgzePim3Hfo
8pbocF9CKW4pLutTBEdAa7ppt8DLWmRwaBY6/IAiYUnF8a7KZiDRjTfldu69jBk/r3VifZSLKmWU
E2W46Khk1NX/DAvyRmXI8FdCJnJXPduW2AfdpmxtnKJzgug2SyqNV3+euSuNlrR7HSxU+zFktBwG
b3RvK6uqVCF1P9XMAcEJieTr3aTtGidy7Rhya8llc8/nAibbswZs/2J4rxcS6WV2py/ItmqWC3bx
uy2K3u+aww6LU/rqqCwszVn/V+cdtGtdm7b2XUGXtorTpLuKJ9ryQuu8qsJybOb2UlTGHLRDmTB7
dUwadpEXs4B+f2aaBdhwo6KG4pPSuHAufjRadUkUAM3KVb79m6lx7eiVa4cVRRCaGNDVfuMYCjzc
FoTIbmRUcARJBFuffiFaQ7SyXIBW+kZTdQqJOWxseb+2YOw5HkcUhPS11Bayoesg0PR+uKH5fiM/
jbzoUSGcer3A4L1tQ10/WgqVna7679++lNetnTy+2B8+GAMesum5PyV6Irkt4iKoscbb1AD2rcSx
TZPClKVZKEfDDGHPEOPp7abT/4eTwgoEEhMS3R4q3VZKD457145FPwa9JwKig/AL8GM+YUUBxL91
tSCoL3gGrtCg3r6OtLIeB9vbMze8apBugUTmML9pcdg5KwkvswDKxUAwSZ7HfohKlXU8DtWpGxUl
CC3EOqCP+hKK4vTFUwLBGVKEzP9GT+f9xCqVS5zAFQr+V2hTnp+hQgR/YXIM76EHZQl6gqrHzXIm
DYJTGVMqi7CTThswdR6kg4PVCg9/CCV4PSPgGjy66AzmTlY7eobgy+la8KThDaQyWLjj4kc2p441
xzxO6ncwAO9rrl6LSD1nWQAKZekmkK0Mto+otfCv8wkoKhR1SPDoPs6tEPbxJP7N81iZC4lq5dzC
BuZHVSkoVrN3dnkYv31jI6bdFPkqGRNeMi997eHBBoQRhIlGRXt607Cd46lTfy1L/y1UDwxerXB7
N3QdWOB2ViaejM8BaLLzvCJaOBf3ChcVpDGXxl1LHHAc9KU/wSMxr8uBgjw5ogwoleavMxylZ7bX
jkEk4uiLVDNtViT3hf+JnKlTHa7bh/rgeb9RHJES3NVCaREOzoMM0ee4opS0bEpqyORwVuRxZRpA
DsevuEEt/0sx6+IlzObIY2zKqauvcRUVBOGL0If3UEbtjAY1JuxNW/Mfp6AEXDIL67VDaruj+CJn
J4w219viP1g5XGKf+0NSDVQIF4GNKirVDP+hF3t4lJ13u6dFtAHQsKf94Uqzn5ov6sKM3jjW/Edl
PCHm6OnbswH91HDhyU1iyC/tknAemlgiu5YeH8xoCMv7ykZ0Xn0F9OZ/AA7Yz9H2rwyt8sVa0bGY
1pMA0bqU70GpRGMQVfr92RBekCzwk8RmPMS3WJtOe26uJc7FhOWUWMDeiGG0SRlEcHVTqiymexsS
2OT3TpQn/uhw9Tu5n4wvtgeSFrik6Mtpf8vt8pIVnfH3PtarsLw55buuksI3iIyOdevRek0ddoaT
WJ4pD34TimUXv2OQgunqEfl6FTO8mCNXKw+s/4fxqiNcodcG4LNamWBQMW9yE/H/aSEyIJHXLcxY
P/BoGteBYdHA63h1R4t+Z1ZqZVfFdD7JHm1LZPKkSzoHmd28N5CKuhKrmMHbgPvNqSq0R28E51iw
78BBxk1T50l71zwuXWHgwh2ZCBZm8d2HU3Sa9tewZln6oXrK6Sgj7SAmYYAEq0kKRAWJ6ZErESBQ
e1soeBHZjxMWyMrXWsUf8tFSAxg3L3mD7zAaW6ctK681Qa6P55fksoaYlLrJXtjlgmjdhc6Ip4dU
YKCyDHH/zXIcuIp2gBWsl85CshX7bpWou+YaH0iFP2tFNxXWtmeSP7WnMisuGnZlecSMskSKz8dS
/4+weh10Q1n0rNH+FcAZz2PZSJxKPr3VKGjO5FJBH5BBGpk9wP+yTu6W3dmV41RA6s56YCbNmK/u
kh9VAJN8J1vst/zRblSxobrX/ZIvS56Cx5RWKZywqXqP5CjKjVxGaOjliV07wPnDrsH21oO1/b6/
o4kqQx92C9lAUxJ8tZMpiuj2MLzclViK+ZM8PHrS2LEvuIWQeq8AUhOA13ddg3R3ia1mdN59hTSS
e+AZqPS3nrzVxIeUtYt7C+eJ8wxiD+U8zk6MGCio3upefhjKiHbIK90ihvm4laIwPr8T0QmoAWKE
WoWs4WG07sBm1ASzW5ynS3bNrVpakwHmfZF+/PFQb0zzUPeyAh6DUCI5vjBVHgw0ypA9Xktxtp77
ejDvqh0vDW18Vx8ZPLmvPFUtF54eUC4dOStwzQilAe2XqRUCanMbSETBlWAfPy/dKIuOoLICELfD
fcAMY0gZ4Je7uAwqE6HrefOsOoHYwkEhyFnYdvHhuGpQW08ssYqhxaAoZj49PGDAx9QCyzK+zLzb
8m/08Oa5w8LqKQw96GIpmEBXe73iuysrEiDdKNAdfKKWcub7hFiqQRnucNUs0MQzoybGLVbI/scr
zbHFZkpB/28vaMbtaUh+L0ZMXYSB+Nn7kcgnFny+dJFIeh2KozGIKnNKV4zAB1sc6FubihyaLjnE
JvKwoxmDYT4NfLuvSI/O1Cs3R+jKulFm1n3f0ohCytmhhm2krLPbxgIldBTx19XbaIKH5gg6xtqv
Yw9ZD7GWZMhMFOUW6XjHD2o1T2QTc5KQiwFeO71WyVv0j/0fWYlETpExwZZp/1N4gTPxOqsSSQJy
3LiuPADTiKwLaO2QHBgT9aMzdp54YAc9nTUygcKLlfa2CmoTZK8a5SGwHOyIyljTlL381i4jUnk6
3tUJnUyKA5i8Sj6GcTF0BMz898lqqxYd2A5yE/anrQCjUR46qLbVF4ZgSxtxb2h7JKVHUujLshw/
qAWj2nzCtjGxNq3b2dSsxK5own2b/SBSffxicNglA29rjdjecccth6t7vS3vmaaDXim+jDtv7ung
N6NTZSjtBrcmpLHk2F/DFFO8RaIHvSgmvd3GGGOyeZIP/w++Ij2J3knEU5pkfSmev3nUgmTSm42F
z7111d8JJF/wuO8UWwiWDb4xVujOcsd5uW/yZiaD8hxx2t8KIcMR3S/ATZ+n6ess/I6kgr09MJW5
GDqQ4FamgyiU9wxCU6OOzYTvKT3fJiURuOaqSsPWGR4y5qd7i1IZ/J7/Q6DOGHkYc1V5fG0EgeVq
jBBAc3q2Q0gQeqA2R+xDmgRUr6ZwtErl8rYy4BtE5suN0rEvgJcPHhRSIVpGvYlg1+cvCjCwkMXP
6fg13L1hm4BMcKNan5QF4PIcNI/FeIJhwDccN5SClVulQsiJxMD1PRMy3zAiUG2POx5ODtuLqYld
D4iVyXTSwrSgPRUEiN2PTOlwN/FJpziCj9VlybcmIv4oGtwhWCJ0wSadSpUJgCNV/oh/RKEqAMuD
owkkZMI12A80txRdZf00tOyPnxl+6kfAvMiU5bqbBYBdbbym6Yji549AV2bmQUNgqITDIksaIABP
Rg2aDqhxH7l615SECUk2tMm63OND2mcGVne4xrud7BjkSyaa7Zu97jjTM867wYxafFgzXbAIdZ2D
s4vlX9w1jE5f5ZjnGpAawW53VquhG3LjDZUKRJErWWBXVVCvfrgvTKLVLUsXxWo4XvT1ITfDEb4P
6GLnhk9m0GDihGOLxOy0m+G3xwdK622jD/LcGThUoNwr9+WIA15JTb5PjJr51gUA5CN3c3k38cE5
11C3PEjw8Oq2zsIY0x5BScp4PTw6RFP+h24KRCIvsveKZc4xcq+zyihbpvMtFsSHjmMfgXZCArYg
mnPUjkP9iXgOUy0PAGyyx2tqgS6k1Bs19eIOVDk/mMGCQocLD+MuZsrqcDsjSgDYBqT9IEBGzeNH
sj4WCsQWVaGPwRVpOpFp+loS4LQ2otfEQRHEk7i53zpkvehjyVdC3RD6vixq38Wqdnv99kLdYpyZ
TAPT/MzDdizWTeF5mgI5/VxSQ9RV9wOfzs2wF9CQaHuw8OHvqgTQmj+dNt+yhJFUuYRhr4nVe+Hc
Xwicx2Q8OYhwalNgH4RJnhwCxd9NFP/Xc8w5POCbHtU9LMHuO4DbIsVIMQFG/VwZtj3BnixIYSVZ
yqid2vHN+sBVPAkhuUNQs5s/ehW0XVYo0Cvd63SMANsd70Hr35ST67atroDuTNGTUPL3VHSdnkvd
U2cBv6o/vCSwhocBAwKIS0ENCcnhwYa03DXE5bDuZs0vd/DI5Qi8OrmPS3V6WSMK60S5N7pDwIlU
5lPgKv6nQsVQ0ZemZHrzgdt1Urd875JbVvWa60SVnMsXO4K1lgWF/DCIJT5qmPpmGCzoIast51M7
XKnjV732w9/eXRsrsENN9SCe1CZWizASafFtVEn1tcLyy7+4+f7Y3RLlyP5iHIKAqhT2lOmzEq30
CH9PG7uGUuAWJ6GOHjzA180yWowm19aAftEzuoiZieq68RzpANwS2Ue4CtyzqJCFIwQZrjxNxinf
VhdtL7D8yHuBHVa80HMsttX/woeY5ibOeAvCOD+w5qWjcKTOD5rqJqyKkVgt+OeNsl4Y7yI4caTc
WZ7rSkfiHv6yo3SESZxyjlclL1hm5YOcD946zji29/Eii/aUBLu3j7wRNdPoclMjbO+3OrZ92sWt
IW4KxHYWbJ2dB8ZXWZBj4KYfO8YVcEq1GdxyJ7JygeAcpTtjUjaH+C5z9iLEwFTbETfVnuyn/nuj
xxkJGk0lKRX8ZQ91Wy7fVickiPe0H3bNcodY34sUKDMphxmfiEQWvJWq19oeb0cOeLGFatTjjYjF
xX64vHX8AbSTobn8CuRrIODZ/m78E8030ihP9fgD2RDLHYxwEZ2rjXbobf2mGqvSuTHGeKed3VBe
mmPAsAiD81ORBhZ+gOcW4K/gZojTwxOa2PjeBW3yUp62kTC5Rh5gOWraMdgivaczLscMTDV441bH
ezt0XtPiBtK8psSv9z/rK6q89NVwISAiGlxNp6L6p0z9HvGg0VDmLa5wKPNTmzoyNwJRdWbYZpzF
Ce3s2TaQsTp++aNGIxpMRCY85Afv7DFKNtySWshXArM7xLv9hQHBXrfz6vBM+1P4CuPnjF75+Z6s
Xdvbg2EI8TaT6kaiMbCxQZD3O/9Z1IRo+x1uSsv2Sk0ogIdbZf+2U1Y+c/9HKhKDvQdLkG8jr2sE
mjJoHxWPbMoYiCi+uYqiAKonCXlryX4DlZt3VCIukYHDhgApkDe4bHA4hEpmyM95b1ublImAi2vK
MF3eCQr+p53JMfBf1wbUcFGDWDB86UnGZXC5kHOBg+DzF+hsYTc/Iped7JzIijrqzQLnYJP+eOMS
2lKd7WtG6z9GhOogov9Vr5Mpp/VVJX+PTK3w5mhnooaEV1pXVz/yN2hB9+4ulA8jSLqzK5oMKot5
LlxNVBblqSAakIOc5TEAkujjOoWNA0jiIp9F5yoVQkWpcG7MGzGIW+IlZAf69YnY13PiUKYoIzDT
tCrxVaJFwg60dxK3vX3fSnzCzLRo/aYFZXu+Qci2L82Y4Qvk+eW3ycPzpaqQFVMHI+w810PPXn1y
5FmRsguJ8x9DSEVikC+n+hAbsw/T1iStSDXtd8DihzwqMXQbrzg2vC/yTXvlbLEbOPsTUqeWiaeg
Y6M24NnUHpzynf9QPuhxEsrk10AO5VgIoinETD87mP7CSL58E3kByrHzxc9Rerp4lo1E76oTQsQa
sygKxHVmVSQZVG9+dmu2WuF582N6J+1JNQe5dKEXZnXzigMTC/+Qdu4P0Vb6Bx/GaOJH+5SWMJLB
pkkj971x40qjK3hiG2gW6+vjSlFEFFwxeq5KFCKqBZl5TGxv3g/1tawY8IVEsbfloRPqOBjH//lI
l3uylDyjHEY6PVewgwcKLy8ZqNPPVVyMOfrFHvBZdhk0C+ifBOZIV3jOpccLaT8OxKFoBr6Qgwk4
kSS0D80Ox65rnHbF+BNppNtmHw6ytTfyJXA2nvrTai1BcdaQohAsvYo2YO2L1aAE6qVV3FuwXvEN
0et89wmUOilx0pJCOaEyvDAhBVZCd1e6R3YIKSnDMABlRoM40wFcx3TPN0/mvcenPbOcPjSHcq7f
8vh8Fu3t9EVCu1CuI6zGgDB2wP7v/ZlvJ2lIF6vGoDoFU1XFABfNZ4+T5Xeiw7UKJfjw8iGEzgrF
bnLwHMjiy9oqiV7RjraiJooE1L8ODAba2POt3IivVeTC7uYlSBNHHg0Fo5C5eaBB2dVRBWhMYq2y
8x6ybGp1FbfXm8Ip3HCxY9OTy+tUIRhHZpla5a+wGh0oNhICtGnm5Ep70XnbonL7YuoHAO9RUrxr
QTyxbgdMDARJBsbBdZjUN2UoRPn2UiMlCm69crFZSKMIAd9fPqRqe3TNfKz/TGMTtkiSY9mc1u57
M6hHPzQv4jbO6oKtKQxlDID/C25+MocNKit5hVi/x/kjJ6VRkpPJsDzX6T4uyLQi6X3jFoQiam13
OeswbzI8x7mUdjMso1w173OsHOVl/j6Tr1BWzOrm61s7qi63TdZGzI/bHoiLBQWvPOyvoiEbRCpl
jd2dbwmS/m513ik9ctFDfXG9CEN9GOHmjp1+L5PyTFqqIt0qMlOv107t/ARxXTyVGyx13pDiGvH8
dLdizGX9PFwr/NrfeF1r+5eWe0ZlVMKoDLf5oP6SWh1kPiKiI//XQGEO5Pk+SjTikdp+/ojealnm
KG1NhcnCPm/TDMm6HYW2zceX3A83CJCffWhoxyxn8dFWRxz1jqIme+F2v6Nb5kLXe+fSiYv/pvvS
HM1h0Rov68tkd7m2t4CVOZ0YhnArh5NvwWbUebkjhnsPZwBEIEmGvhk2DhZtW4zWc0zxtFI6sgum
dLeIxcaFElM7nYHFtT/DV8SBe7vN/ulqfL2WODqBlq/DIMs0DaANEXvd4Ad/SmFGCfRs6bYBE7DA
TelfUEPl+D89HuqCTd1dWsrqFzjSgOlqc5CkQLeiJQyLaD5j6d1mBf+toodMr1u1gnroUJgz00Ir
S17tTjetv2aq0H/LvE6dXSAGBZUeTHE+2lRfFu9H5L10rzWRqQ2cxREowKMyT8N0iz7wPaKgH+bQ
pPaMIssWkuus5wMc+2Z+US5gfRAYk9fsMK9ZJR5EUt6adgU9y2Vv9n5w9LBTc6rKbElVXCdMBdyt
lAJ7Msdvit7lMuMfOqYRlybef4aRM41m3w4wj7x0AhFF1AKJjPRiApU1SusRm4BkWU+nKsDpDBbF
jR1EmiAswzjSGo5GIEOUDnFWCUHC6M19oY9goxHK+X+5L33ZQV/kWpsaegEVNUJ9xldmvxrTKm7i
fNh3Bwcv8wWdXA4moFrBmfc85XE7bjFXJxRo+mvJkV/5PMOoUYmu6/3PF0yjOWcaDxc5mzpKxgtA
JJUd0x6AtttgxQJzf2EXR6n/nj+aky8Qk5S1GOM3p4cPHbeCo7HiN1ihss68P+WPvW3glOGIpWXG
t/8CVQ19v+VD1NfEvutwIK8ikNHWM4BZXUIqu5TTH+bzXoLIzxier3mPrzSvV77/e2DYOgXRUHnb
9XMDR9ylzOFAxrCAwjniSLm8vKVmnXHxBx1J5aV7zWpxb1suFVBxQxZJ5jZS6aqRyB4Cx3zAtZo1
g+wFxB2FVf9EmlS/rAve9Nytpz04CwgJ2R02m9VIE7Tt6iWYBG9n90v2Es2MtbBbzm3orUgCr74Y
iAIl4/d3/2aAQuOIJzkcWr+mHfqa6ormvWEUIeFusBQu8Rz4OZ7CD/c/59rzPXzZVmVj+K81mOGh
vRchxVnFvTXJQHnLP5IMZUtBVfDDETx6zJohmTc4gaRiueoZG8Ui9fWctFsBjXUB8CA7XVz99UVs
xGtdoFS58HAhFolLs4fNxW/MhgTK5xQJuy/d/d84UUBUoSuV2EN+teejX2XApPIkeDp3icRTcShS
9nlRZOfeWY3P0s9Kp6wDfyHwdQ0xDhptuJfj3siq07ctjwuqzCyVftOEewv7sFHBGo1XPo5HamXC
b3lNsS5hIwz6pz+7Kri4WvKLWjRS1uPDdSArW8yoABVqg/mV49MLm5Z+N4RmPdOq3qZCULWjTC+e
CkMAcBwhY8xtWSzFYiFfcmAjqf6vO1wk1I1d5bzNOK4on1CDdrpxM+g6YjFD2URD0nJpSrEcniUk
k3xN2KFC/JlfsvEBxRe58kkWG6HdfCfgS9tZmnrkg7lb912zYLU8pDDdfdZjKaVe5NlrgocC82BZ
VIkDMJWtJJLoYk3RmtoekreHHkN3/9Us5gDif4jVjq8FaAnpACcWOgeqnWrgO6zIdmGDfBqUty9s
OQ2Xid6dHsGlCHiAmUK9x0iBqXunyjz9CufnLb81GlilB256PWS7mCC4B6DSuAXRdV3bedzgmKp9
x7QbDURUJ91TdrmAfkqjFF54ms15FpqhpP77dY0WSCVh5WsqAQlrol4YKrQPwyvcKnJ5+qxSOXLQ
fVNAnGz7Ug574Qgu//t0ac821N1ep8e+/u7Y49WCWhdLzHalP4qcm0Qth+4TJ07GaJW9hm/a1fVs
5C6cYpfKV5Vbggaxb419rjC62CUkIjWDuIWNI9pn8MXFWs0et8tZkwZI82HmjYZwH5jdDeGcHybt
5w8qIKEVCDC0v+KegPm2oakt2jZ9R2TWHXiOD1RbcA/OVwVNTxyAJDNebxBJzwE6K+WnqOlNdzWF
7Xd2tA3rj6obpMmf6u71VohWx69j9xNVNAH0ZbtGOrT2q06RIYS3uo0GPmEReyqy0ei0D6Yhp6Oq
E9HLg5CSMH8KJCVK8ZUQCi7yUbSjuznE6JifVckYGqAa+hEeV9Ex6jagCPFRKUmRcGAAbZ97+qwS
dKX1Sz31YyOQEXp/u+fD2IlS9ilZz37801b4kFgx087rerMTTB21oJAr95/gEmd7i3O211JjxZ4/
tR55X1zynFyFu+IbGAhGtNXlGTaBxgXNdFcmGXxu7Yu7UKTXWRZn/ROFY4upKGthvWPQY/ON62bk
WCGmlLykJET4pYvd4XutXXnFkMMI+juoFab0F3IUaTVJqYS3q99fvvSHKI+i/weH3wLjBcMnGSWm
VC5KcDqVfz5IBmnFwulOHZJYIMcFqTMrUBuUljfq/K9VQwyHvwx+h6TiMTbuyLkOeb6bguaME4Wp
RaCUFzxAhsN8xMnQKjDDeHSRIDNtDeDEZA12BCEY3TZxTdlkcnxiX8rFNGN3PXWf/O168fkhVbq6
VKXfKYfvM8OY85UBkpa2ejdNZiDNskE6iGI3JxCPeXRz5NPRAoO7dWO9M08fc/Wl17eVG+02ysIh
Me2T4Dk/YPFr/1VaOYkRkdQ6NOjG+b40dEgfnCP/+L+8m8eh3Lg5o/7Wk8Fq4gJg42BmDb+Vdtr0
SWksvysDetR6HyskYoE7WmFcD920RoOlEG3bmv7QYSeTA1qN6xoMMb0lXRlFFqD5XWQbGwBCLxyl
8sVgWU5w4RLect1D90zECNZoSiMN15hIkVx/CFqKDZ82ypwE4ux21bbunu9pFCv7grG/d628W2aY
i2cnFP5v34PURGYOH8BTFH5wX/xm2ZP95QE93hYXhUI+b6OL93h5cMvhmDzx33XuZNQ/3RVqvlEH
0DDyN8y5Mu9fGnH3cfw5g+Ze/RoY5ZZojrt91neC68au9/mrPBfmJGFFc4WBnbnMmVQUryWbYmV3
+PIgBVbOtpQLryvzRvS7MbVqTKFAC5NI/VF4GGx4hr06mdQ/LKtVGTiYGQT19/pJRc/ieVV8RPWJ
ySqOqgQ7YENetnscVUB3mQxWkBD7vglOCatLZgXVxplybKH66RrrVn7ps8HUFGoUvVIaYjwh/I4J
LFWomd3cS+LNuMc6Nb+bUQSgcUSGmzDRbkZzVd6h10Wx+BRbIJxawTyYe0fGd2OYqcJf9KfG8jTR
88zTSzKcg4iVVsj9HMqMFJgvO4wj+EfXQ3sh0sRjejxoUgcExShIEYjKFYBQGhmwx25cif+bSC7V
vV3NqUs3N71ubCVSGV8JOzaUg+SIiBBTIqUIc9EaBxJbaKSAYipMHYYXLiOjqqZmX+eCRSSydpqC
a4YgXGlZANdY4294bjhp5lvYiZFDEobkN3RBMUxzc6cDGr3uD8Bl8D4EZMCJayt6cCcfcX7337kT
ezXQOIPXINCJJ0jD1hC6Gv2RQdZo1Cq3W7WaguRo0dL474/YD4XwFCO+AaxPg+teIvQarRhDSe1X
yW7/+QokC/69YQUKxv3QvvP+RZS5dKpo4F2W6MzE8IIUpO653qyyvEa53gUxb1VqQpXHRz/aNTuj
R89+xJ0Y8aWQtAvldionxavUQ7q5fbAw0U8ETLcrJYMgOvGJVgzPsjC/dGOcwY6H3jXBg/793IWd
UHyVC/kzUXN35zmMOxxc2w+TnCmD0dGQn1AClypixhOvmzr/ov7BhUM/JvUe/sf5zYPbsdz2nfzv
zF/fjhKhLIr5GcD637sx0lcM3QFX3Vs+7QcEttM40QpiF2HvE+GC7xTyGlWA4X2SYZ/AiHVtqb1s
hc1EJf4ke9A6GoptS4ZEPJS1ulTLi532k++HLWis8GcmgEltxXwXKMieIhFXvgNKEfZclL33bB5h
y2eW294nHJ6pVSHLWQCsJx3ECE/4QXvW3sNbALcZPFbm6i9xmSLBmlkEsb5/Oh8GgXPS6jGzjXy9
Qasjo/bmzi9I/q3WR7T7oNupIQovJqE/KMEWHJNaQoxmDY1jzrifnvnmV+s0oexUiDlAVssGIRPe
EbM2YQu9lJduuvHwj0gWsIlsOgagw81PWeDYIajqV8UZuyhmTswA8nnxFueJw0gloLM0XAdsbgG8
PfAkxezP3m1Cpticop3s2ESG0lpucsHN4UZ10pO73l6tHKV03pRqczBYa8k+mT57MpqLWMq+68Ho
fMQAwZ+Xw2CM099woLhLXgJRmHmnuWUrx5l2ZtDy+2qTDkSzJHoOf04LqtrAFc/pzbqMDnYcfzud
xBPCRCrBaSg78885ZfDXLyoi9DF3dgL1nqMSX0BMpTbPBUCOfPdRQTsdStgqHzX/Td4tHNNMFQPF
iRaQcLk84LYKdR/80dpkFhCvTc4pKEcCmGtrS6mLVPxFtXK4InaXgTHe1vKDTOYE7t1ZPn81M3Sy
h7vqHelzeuFw/Bzny40//FqGcjNzvNp3bBMXMAJg6Q9tGkyvoIBZfVrON6kg6nrAtS71zueR7dB3
06fpixHW/cy6w4XEh1KvTKKzbLS4mBtPQc9H3t9kWs/0ZbrhFVmBV/4aNVR5N8YY1YCsVVdf9JFn
S8EAeQvc+hriSon4kUXrqZzNYJWHxhLmrXuCfV/RmP1gYj/3soQkv1uugZVAOnXvz7UmYZ18sFQK
vzMdeVesMT83e/HNvcFnbXVlT8Uxl9/7e0FqLYwyP5/0c7Sfj5gOj8OUwGnHr90fuu52+nSJOWs/
QvXnyNht3nghbmcGSIOIc0XOIylOcx2uS56TvjXydzsFaSrfp9e0/wglsFY/rPrmEjYyRw/OicVK
zDO9mGA81/e8+psG2U3MuoCbTD4AAUE1tAaymxX8Qb1vX8bREj9kYF4bJlepunlSY/cZqByouOk8
o2u+gPY63MPU7RIrZBDWS1yecRcwthxkiXuwVpdvNvFZO6vtXi7mkJqtDSvlYv24y/TyLQG4mcvz
VfHH7fUfIgFcGra8ew2r3QH8c7bjQKcNy1mTUxPknJodRezEMEBpSxV/X4oI8UUHgDsFsJVl7MO/
xibAJKezZbgT6/evXAXeXZjdYmHXwYk6jW6tp/d7eqJbi3aLnDRrxOCBTfJdnNZMaKA6oWQPgdHR
cFxMBfW3J4GFq8dUGipAJ6N+Sl1up7dn5Rdop2PKP8wUvZmBhH/p9vQIQAaTFPPKNV+10sUHl73l
T7qCDp4jWEc9Ho1YaPEceTKueYxCgOEUULcyqI7j0Tc7018TguiQv+LXAyjQzCBMqldqogH4iq2b
fcPU48vtrtiwtNvDWi75zA25Gb/kOVB9tqtqeburlS1kqahRMjonTo7WVn8MaEeY5sZzmz7MsO55
cZY1PHpoXEB9QdK+Ylwz6gx8wAEDM4Vf3PNTEHWKYmgSer+llOF6em2pZkck8YRJYg6f90SMzF9w
f5ojLqYoVfKVguwjZMdkIHawUYC4eJHRgUgpqlygy0zlS6FVwEYdDTIUmvBW68aP/VypQ+rbBg2e
ODTBMjmIRJ2pl8A/V7CEoHw+yN9x3WCumDsDrwqdAH5WlQWRQegmSatSpFYzloBm2slA2/9CSEXv
48z+CHMJ3tQUWqKH5MltpPZrFWfJ36T4qrUOS5q3vjOrf7tp44e+YV4lIkl5wVL2IlwRnfqzz5ZP
k/l6OkbdRjtdevTw1wcC5NKC3DZIMZo1BpCvwfgN+T6h46tKUgP3ndqVWlez+z6NiuWD6luqk9eQ
66nIkSlrz19zD5tE6J89hZ+fuUWqO2ly7sufpSVxoqhEDLgMaOOao4X9pamUSi/9A35FJWclMRrJ
cfequnSofWM4UTGmkhWuAUdHB/QwOW8Fvveo0QXloxtD011UmqiylYkInhStLfQ1e7HDCyQPJGe7
OHF8JXGh9TKgxLO3wpnkgAoKn1gY6MEubf9ANUYhI9vKIuvvLLS7rWmFxuAgia1XBswsdotLuIuH
wtG4Dkbs1rpG81fqnn/DlhPEnPm15KGB+4YM2fPZbG3BvRGmLaFi+3d2SBykHiBwdU+d10jubqfo
5bJ+lTHMCWZ/1GCxai2uaC1Djxn6hJIdLoMHh1liex28XQXPbT7qxLZxRgo/wBFW8eHnhTViIUwA
WS+5ZN99Uv6yZBHa8nlMv8PAKxKsaiwN2G66LxMs0oMcDZWd47IgoibXSS3ukPUB8T4P5pvjJ3lU
Rm1JjNla1ZHTlDfx9loe8U6LfVujZibMK7QxqhnkO8PVsB0ZvHHUFvTT8H0BirfaBYcTWm7QxyTi
VnguGeJ0ZR0QBnR24XlgGwkSHswjHEyI4u4Oq0BRPjBHXbJb6I9zSbL0xh+U35w/FDZL85GvRLGj
yr8p0J9zwDl7uO5DxJmbdVYVvAyYn53Ak6JKlmYhrErHeeZ1u0bxEuieIiNEFjlQJ8u8qMHtmbqo
BS512rPKPuJIAuC47jTD5jdbLb6tK/+BgdNYnM1Djea9CWdTtd9ToB9XX6BuFqPV16K2OYq+l+0P
48kaIYPrHrbr77eWamg5CZVAS3/6NmskteiNf/JFv1BG1OmUD69Q80pdmCHjjyQQNlTurcmHlg4J
zFslyK/4tycJ0cJ7FwmwERE6zB3T4Awr9TMjC5wMfkHmiwArFuB0m9y7PeKKyQhSSooM89FIgo8p
XeVdv8oC/1X8Z6LFzvbFckwLnhxGFLnHl3CCO/4MJVxWZru2hXjNh2tNWsAsGDNpwIjqZhBRVEPs
7UP9JBVqnINFitClQbs3F9vawYbsvWtw+3KeCrd6YcVnHB4dEAuCiFOTuESaVwix6LnVl900GQTc
CTbF1rVBmOr4ovIeS/CYaVvF2lk8RsmV9v/n3m1shF7TVQhBWYDgeJqV4OJ/IlmQj5+bmCH/zSan
DEgxFz1tDwgcU5715HrSPpQFCBah9JjLSTSiT1tkgHHaMYKfGNgLBv896d7qS+DdgHPtWlngOtS+
Snvh4jMjAABmP/D/iTF+rHuWO0Z9u0jiFqNpFzgfSuWtUnSpb2WKZCNccbM1d358gPuihkmjmPgj
ocDa/tsH6hfHvy/RTkBj6DKaYxOA8GDQp+kjzGkxj30kVKarPrR5GGxmkzO3zIX2xyBBRey+Bi/Z
0NMl7oxDAQmw4XOBlwUUCYYRasl9/FTjvdwbyzfLZ0BMfyec58QMGvEa2w+C0yxutmaV7gceOBti
QvAATyxOT9bZhqi0reAyb7rmvGwuMallSThsGLkLzVsjM8iGbjP5aJTS7RJhIG8yabRyfsblAepp
FbUf28a++h6uRJL0YFkjHBo/MjKLl5FlClC0169di0Uc+K1xkEWy936ozaiPcISIoXvPc1vgvwqM
neO0HaD/7zgwVwMW73YW4elVK5TjZRdhSsQ6idYPF/M23vQCiN9HwDmxyzR3rnhqk175DApGiJ8y
IoLyWNkfn1HbBvXonwE/12oM/NZtDQMXwizmn41yUWF7Utm7EU6mh9meuVi5J1IW0wNrJ7njvuHq
vaebhVBuS1aU50oS7rHc+ZoJb7aeCgjLeg7h0m9ZFYZNjaythR3WEd9UMyMfF9fjGDCSt6kepKRa
XWhVmMM40AJMRXKHYfXE6gmdwoy6VlCDqWaFkeq9mWj3CzzfgUxfATqSyqeItQan1fQ/nZX/znrs
2Lb/7CZDT2hPWbqIffGITNPu2HPT9D78G1zBSx7TJIcGmdkj8UkC4LAda3i1KXFN1/LxT4pLKKzH
oGah+NiADMxARrMNH4y5D5u6X1+lwuFzmnw1KAt+ptOWb2tkgdAmlDZH+J9O/fLpfJ3eGG/tK5M1
JbW9CkobCoM1L6cbhmDJxBXV1rCRCSEc0eqJSzpM4J48zn/ZwFKUduKs1A1TR+yfjmutXHWqiK5C
4XRTtWKm59V7NLhirkJU8z9eSNUT2UU39W5a5eT0qGKSTTfj1Sac1m8jV1UIef//NMmikmO2ssU1
l1u8YMmfq1pAF/OrZXapGPZPnL5X7aE6l3b+4dA/AhIUxUtQSGACJtRBtGad3xNfIfnOjer5Zjb5
Bi32bXeM4TAscPtXgx88QFphKeApslBCQAXG6vZ5uoL+Nx2JBseZq5N84zEQ5O4rMZR63Wf2cgen
HmZDlrcocAoOd4pMedWao3/O2c34ptB72ZS+5gKxwOa8zmns6EhV4CcSN5aygsCVBCDuQiUyA1q5
lmvl6dJDlu1VnIN0nA2bJ5vS600b25mYdRUCHwunOs/MaULtWZb8lK338RzYt17bohz/njGDbr68
niVM0Gw2v7CnZD+aFG8HHeLRgDomHswmVz5MNTd9YSR4jsoxZZExqNe1mXU9wBv1c7VYJdLB+cxQ
0bPHIbQ9BGY+QONj2URe4M1NSN9C2DV7eUhS9yc6IWUFsrCGOrfWohJOqL2bDDEZovCHkR87TENu
ghprjsFsveT/sx6UdwETIE8wTiAv7VnxAUdFiCELl9ACoTIbozcJwoaXI9LAWjrxZY8jkU6QpVOS
k6H+DWm1oAGZrPt+TQLkL9dnv9Zz4ESN+5H11zi1+RvAXYOvXG4QEyyzrj7xlK+2cLBWeEdkALhw
0e93cWTBTb93ruGyW7IpFKkMXtfgd/bagrlH0sCw12gofNa/BHfauGu7uQwT7iWasjCLhdBuVavt
evlnbZozUQvmx0bfO7j+7/luORT3OQ7uRycyc8BlXSfSM8jzHlDk+AREW6OXI0mg5m0uSktlDKr6
YNevujqdfZKPMyGaBDeTeulStgEGUylzwdLqYENI8saBZQ/G9ZbPU2QQsbtycL+Djzs+X7lo+pg0
uMsxezej1wLNlA6FzCFIfmUiclDk9n0oOAcymn90enDPvpgR7THwaFYqtTg72+HufWkqF7HQNfLC
rkzU4mADKH2CfnbYQynW8tzX1A72mgeHoSQC97EvwXQRsCS0DI2rYL0uzL18qDnOL4m30Lf3nt+y
M7tBaLvfOSWqy1EspWkFLfd/riZkLMK36m7yNZN4ilAIWfESoo5fQ5oQoGgN1egqAqKLhy4Ysn5a
/d01sVB2djMWrlN/Dhtlfy7USVf7ODPTYDPuTtQiANAGwxrn9m0lY/OKtHywh3V1o8VRf5tnGZQ2
KLMlyMjgm0bQYre1FY6u5S0ZNdcaFiI/NPgxxMPiv/3TmVNjAuzkb1K4QEfKcgQIN9UPHHpbj3On
kXwGDLAqFjpMWFjQU5W1HimIrJMwRfbY4ww5onHVc0Ej+6jKtAK7czLbmf1Yhqjp4G8Q5wtoWFo/
weNFvajTyqtKCDdmVe/nk9yjvz70PjAPl9pq4N/bnnL7dJIpkkaDedWNFiwLnYinuEujpb/qiI+d
E4Uo6+M3gfDNpSKFfAs8XNW99B/FvM66MlJas2nIxl3mr99b/9tYmbJHIwLV4G8nIc8z9sZ3kNLz
HW5+2Zj8NuaW09OBnAgMajIOfn2eu0y8Q065vN8f2FBC0pjb6mM5EUtfiyu9NoLR4iDoql2qhS4o
2+y9WlOiFf/TCJ4+wl8/r8DvzMJlothhOrIyaMLUH9iLkrXdPa8Ys4QXByLmjuoOBpMddBZWMiap
I+vKRnYri7f2QR2muroCL3WXVSWkKnw9Z3qokhOuPg1bSwSMjsw+8QD5LbLElkqT1YhYm25Ek+/d
8Lm0M+9BK/ek5k6Hk0pCS1MAT2UMiSAthrmfov5IcubJCDK1K0XeecfJfMZHuukwKobh2XOFm0tq
EUxFKDndxV+J53T268X6FNQP3DsHvLDIWUz3aQlI3eitCe5jcg/Q9O86rWkE0K1eyvFgT+hhRRmj
YzDnM5Ng0PdOHMPKAKrpcnBV7KrsZPkx4pm0kZm2YBnu2/rEGVnR5KCiE9P/RUnByP6U2c/7i0O9
N3eSB7HRB8S+vCd+iORBrqa95Mp8+1w+ZF93twKu4qf7iSWGn8CzWanhcTxkpEQ2kSt/SdjTWT4c
L3AP0cquZ2uId/30L5pVYNlQQQO1mUi5AD3QHemVm8WGtyU78YJnYOmUMkSGtlxMWpB6ihGojQf9
5AX/ucmktPolM9g/IJGiqX7RYa3nTKuxzl1Gtu3UuYDTft2P7lUIPSzST4SgiASeHlZSdBb/IlLv
Z7rKv4h4ZZRWZ8u09yWm85hhxCpOSKo2ZQmR1jlrFhnXfqvp1XBx2cSp4IkiJoYe5zMRSVOfTccP
L8aj2+Z/Wmrlwqw1kA/BhA0DCf8PAyX+BcUvYe+nj6Q7OUcf3mJdjvY2v6O4F8xsyy1kFPEdAyWU
6FTbfb6HJRiiuLTblbqnEU9jSnljPZkp4BkrTy3Vg26ivFTRkqQWcgRyaHCXXfABlAsaXbuXcWXV
pKXi0YLK3nUidiVqMxeD/Du8wQZo1VJTNNhw611wkNmvGtXz2dN7RSr9lQ0KA/O/u0UGi9m29xKw
LMVU0T/NjZJQPJShyNHwfhrOJ6BCiqyJaIyNkQEm9yNPFnTRt3t9179tD7KOSys2LhRH8jVBv7b2
7G9Nd+MOJmhlKC4YCpt04ZGPciAvkwTUWQDfAGB1DuC32IcdrRN15Qhn/9IvDXsZNGmJzlh7rfZs
21W3PlwH5j96qAjFS628UnXSNV3DXuX+2/oH0BVktKG3b6sFmwjr4CkKHtG85HYZ4hXQnTo11j2a
fqMbZCFaPyUXTs0QnCtHQb4PckYQB5dTGaIvPwpGDUkddfcHFnsCw/P21EaJ6FzevL0k0GseDZtS
Q3NxM0xLYnYVSfVnREbVdrFJn5XiEhJXb7/hDIhU89xxu58JnqUvuDBCyChKs35GH2lxlWWXkaB/
1kMaiOhgohhI+eP95HfeMBhn/JxzmVJ7k3E4lVFvd/vs7mO3BX4aHBqpJAgvt9AFh6+0cE6RmzS9
qDIp3Fr+mAESNMbB4cKxUDghfkQWbDM5+WMqI4eledllO4M/ubu3IKoxTUJvrTyF8DXz8PRamrGX
JJV0S1YsPCr1sfhGSHfUp9RNzzhUHVHWADdsKrjCycGbyYeglnPy411eDX6ME8KTDXK5sMBdcrOA
E5W55ofXV8Jvh2BkJLD+UPEzD2sj5GBp3Szd+NdcaQaoy3XLBVSQdieT7nCq0lHTqQfOiijG4dvC
7wKsCj4LWEK8MgvvRQGkCdQkpJY1emMwm4lsdatNzDDu/gbVKojqVKB6LFLwrXCpjjnt3atClZOF
VnXsKOGdymZVRzlLjD++vyYw7u57q+cACK/8Qyp9FbSVqDjLNk1ThfDY9fGnzdcQi3B0kh6JSRaV
+qKDZo3DxbeRm1XqljlfrS1vidPk68tioM06WC3GlW/1P64coO4JA2aNExEUbZt9gKiR8ZTUzkki
m1Du1CBqc9GrslomyTszJooQA3kIhK76h8cC+cv7rf2sNGt17X9Kbb14XJV7tlV/0IeLyvLPmEJN
RByYuhe8o8VwDZagAFaCpcYPGHWF3FQ+kVw0PQ95Kpnr9TpWOzpAX9mJf9XACg8tkA8wT9XofG6h
ed5ch0u+jKgqemwU+8n60ZVbBbrvwVFjQSWrPU55NPQhAGfT/N4f5SRyC2yBWJH/1eN/bFjoU3Xd
CcbM+jBaIysa4S9bYFAYYpPzP7a8wEW8ndGSeSy53y6XWSia20B5Ja8GT7XiLyCXv+NUkHhNv0A4
59TLxt41nFpQT7w42bxjVzroMRUQi6aZEjzsu7QN30U4Sjd6+6ZX4yM3qmdrJqq7ouh9R/+KC0Ri
0QlOMYQw7rfYjipKtanQTgUbYDncZd3CD7ePpCghbEKPDwvM6mHLw0Nb/Tu+UKuzBo6uHJr4wdqj
b/gEAmq9pEPISSkQ54k4jDa6NqpXNeJQsESn5XTKkyJB7+NznxT38ZV6AOusATnT7ZRh7f/iSRFr
vUA2FUEFblHV2C9U71IT6Z6pvFXBOuHhwEzEt0OKa5P8lbN5k0Uswjl6iwjAWjxrWNwy8eASZI9B
adXWtPcvqmsSX5T6v4iAv1QkNdjh8CJJ2VZjEBd+r0JjrLcYu0Z9wwmblYBi0LS3U/INLrxJypla
nI0A/2mTDywg2dgzrvs1wKYr/3YXfX9edAUWC5aqjTsCxq0alCgdfZ6kFAuYY2aQFvQpx6gZQNBn
9PuQx7HTkNAbcvXcqyGqtXuVFaA1yufCjVT5WG7e+uxESd6UPJ38C22aF95r8ZkygN3PqIrkKTRW
lEBnZa7jEuOxD+38RHtAiSGDyRlUWPOPZhTNaBjWFzz2bHbyUwdxcvEc6LX2Z2ue5Tj+XM92FkvJ
1my56NpENGKosmSQr8JYkwjhJtesZV4hna5b5yycmaB3XBysAPkEl9vxJYtM8x8CDY+2vXHaD8CQ
gSs4Xn25o574Mp2zIX2Mw9/0YcsM1D3emO6z1/XdyET0k05SpIMEF0XuuHPkqiDKyYpvFL864n5R
BjuJdEDlKcmRvOUN44zRL8HHcR1m9rI6Kp8C9Nwv4Cy8Yx/Dg4NrgVFnweGmPf2vUzE5cnphRsoo
LhqzMUs0L/KYWsJR9P7hXpSBsl3o/hOSdEYWTQqyVS70htPlSht52J9gJmLTR9cExc4Va3rFrJmq
IBpVXt0bCWEOfvVqV4U/bmnFSAIr3hekUewwne8UOjkX23AlJ78ojrHeSrcLtduMFg1eqAG1iiAL
ich2khejJ4nhHBCoOxSUy2MiNF9sBGDPLivC+JdZhZv6begNs3OQ7UbLL/L1UY2opLDDuIQN6O1g
z6VdSkhS9QsBNxpo3ogxGr/MTeXxkvE91ihC1/7an0kl7PTJ2wTNv/ZKdWXlbGIqNJUyr2AwPyDS
uiS/RgfIGFJFHahsF4G7uUkMwnNhgtp5oMveKn/jEgLNh+lY9ME4pggAqoBuCGL2lPwqzvyWDzqd
VNcu2HQyis8L0NM8F1jniUda/139jzTNyDcGrPjS0LQ5VMcLyEy5o8hCJBSdpgycZdGizySJw3xS
NKgTWWBRzEUM7Qc4wcdcQdgdZE6Vjj3YzMOvCko8rY/Vo3x4g4nkqzfbRCaE8Hv0v1zdpVwLvg3n
8dsywishgUqRIbSn1lhyg9h9+2fbp5uZg115CydQGA9pJLAx2EbGjbpPIE6QcjZ/DMkdEPxcY4z8
x1/m075AdtRiNBdYqBF0TX/q0Sn8gmAt3Asl3+syvbPfNBUwOG6hqaJUmjRtU8ySDjzHFYSrSapu
VIn+I2bCaqn27r5/OGnb+9Sxg5yA1Bi4qYd0vM6vKlgrgMrEdwzWUeirH4ySAPJxK17WpPkY96Bg
2M0kgV/GomfOQxQNVF1aCj8e0gxMvoruudxysO4ZxiYNfyaPhHhcdzfmjgnH7N9BHLPDpC139y9V
JF4NQ5EqZpkY99JZif4KnKPp/UJYlLcMWWMtlHdb81mPdAdWwevyxBprD6V2aWIZWVPmC+pRNmd7
SrwcCytNtUJ4l8ghxiBpqlHIqcpWIqIslyYREx7lJfPvFo+eFgem+NRg9pXO0PkjSqP1o8v5h7rx
7CcXRMjYobNudp8RUqRZ2ZJyhXfBovECcbaxltRIMbiQPcS59C2gFJefw5SKeLW7srk1TqoRgLdo
Yldky0lv0gXo2hmE0+t7WwbNcRXQhEbUjOmY4w5vNxDlaqnk2IfUPU2kDe9NiRd0BQ0Iqoh/9K7/
FVgfU+nWmZQR9oTmKsxShA3FxM2Zp3Jr/sj2FXsHjCzhp460gGttfOHohisXcynztif98Uj27ivD
jjzzxZQBpnRNIbRY36p1PF/LHEP8BNQYeEOmMc6ntzODWSL1CaAz4kyPbrnOAPhlLGESZMKpUm2j
BbBBkOpcSN0b5sPaAdsfNeBjVRcZTGHQxH236kSfSMl53CW53JBuFpCTA28YaE3t0BZ5lTjiwQO0
xwYDH26V0FJYg7S/oMXLXNnlCWi/+izkEhu3G1MUjQdR/Q2ecAHbEETU4PkaCYiOks8CXPvTjqLw
GbCGVpFhLghK9xtJP9tLCjvk34/RGxmCZX6VMPdPm2PTbXAtXOa1Q1h4Vmyh10g2R1CVBEV0xafO
n2yeuAKFtuKVRMigzBNyi2Y5kKqyVIeaz9y3UxnccxZLnk3YBKGdToXt0qBynNL32CK9Vbqe2Jpo
lOwy5DvlU7/SZhENuJGOsnJSgRj1Oo1T2qEhUzMFsu58D6rmOzp60iyYr/on4FOpasJqOok+7OV3
5szrP0LuT4iF0qca+bPqmCnqF3/G/EZNZ78u7NspBinINz0putj9JHl9TBUvm4OStdJIV1fq/Yju
Fv5CG6xC2GoHkibyAfTnlF5ZSIuL4I6otgjDnjqkAKrNghHCBFE6CClUyfD9FXsoPC7UZToegbc6
3qKyKUkBBzvo+hCl8kMUOGkaG+RYSad/KaehxTvlMaFfUsmVtc87DRMQyOo7sfW6oE2FTOEnYXwL
s6MyLsGbbpA2B0sUggoyaoNC08pMuZxiY/aCO0efyTDdNzfIfEkthU2eoBy1DTrrZ6PS6ckL1pYT
fAx8IGCipPdzJtZIqmVMhZY0iMABYncXhyLj80zNWLXhEYE6ZJ2Rw8DboPlWIgGCWMerwc+iHARI
hZS7u+IVydgRBdOmyBucfJKclhTbw9r5Bpy+uqHoJ5xtmtKTXFiJZEgAT9Fic8XOPbLFYgQUzqn3
gFZ9tM/pkFQGGfUzC0kldfjhGqhg32vvwZl+8Y+fVaB7oZJW428eE363v7YVN6XX2Rffd7WWaYaH
xhkIBrdAZjT9sazTRV2cdDMZnjfZr2XYAUNUE49g42prjtInPGNmRQLZKPbPzuQIZ/rkdUSZ4G8R
ynb5kVso09OsdHc4BjLj1BQY7WusOEWCd4NNoy20nfBP+g4Bn8E7rqss1dInX/JHKT/r0UOEkOwz
HYUC3EjodESkes7LIBLaJEeIc5hFXjEcyCCYxwRRxv2GVGEsNxSVqojd1sS+aRNodHCJtkgjfZEo
QnpJIn8s+8JYEUvWEHke57BU1fydvZw1K5zjpLCm7je11m4Zl5SAdvWA6muSrymGifgI1RGxUGkc
Maky3iST/yFQfCSb9G9Oz8URzDrs5X/spHSHucDTzxDXFkZkUu4yVhFyI15Q9BF5uJYY9Yti/jsM
xtmrpZbNXKfRmKbA+IzFVNRmc20BLyYvQ/OtLClf4LmHQml4FlfuPYU9E0R3gyhhtqV1K1JnSbQg
DZg8L+HnfswZ6i8Huq/PL0aUOhiMXPDh3q4QyWCAeRaYZnFOjgN1vYE8DZNbkq4MgmzmRVCRsjdn
nXsoEFbjMnFy8lqNUeOA8UnJVlyD7+10uyGJDSa9iSj35bjys7l9eXlMA3wubZcVRuTA6/7JCx9j
dy+YYj4rjaAQ6sMnRO65xgg7nKO7QZT2sLGNlxmZtyskfwUF2Ay2iBN2RahmJAGsnZhTKCtAWWDC
e4NyK/3B330xDY+p9eljS7UdyDVkAJdTIwvqMA7miMAk+JJf9g6kSbTd8RWU1JNWeRV/u4D5Z1gD
BYc2tE2SFYoSmymIFOaFXJXFhaeAxdRq3Wsduk3zWczuxHIQnT7HNMP9N57QdqjJktPfqYid2504
llsFtm3BC5jdEaQiG3PQwm1w4+mKzHBicHan2jLLn5c65AF/VrIgCPGxW97Mo7EWaHVQNalHoAoL
wy4yXyDJH0AW7/F9ScypdwqubexaP9xYGHneg2er8J/d8R67TRaYMHuLqK3C1vF6rnzStfA7WdTq
QnFUEr1Nbk/7zVQbxJRFlMin8IT2qQPXhMmBEA63r4k0FpcZZs+OO/eR+lQSGmIQPBU5o2c14H/g
6ZI5kedeleMGkbydlo4gkHA/4CKtdPc2h9cpt94T9x3eFsm36l7tAEP8+d//lI43L7symIEWMw2o
nHQnAZd9r6pbZgD6AzXHWUs0BS91QccLZYEl2DTWtsc9HHjsT2fyhcDlzKOmeIrmqCzsThrjLoUX
Ti7yDW4LrPC29IXGwsHPS7j0Blu3ZpgZtsL0Cg38nrE4elRsE0pka+CjJwOvzsbWy50waLUh7EK5
r0J9tX2HIrHDes7p1+OOYJeRZuv1LK9OjrxlN0Z6zFBOEtP1wJWizv+HudbeTidd7Agwacg61ae5
Qzw3s99wdbZ5CRSXw2GWouoX+YHA03BaeNjiL5pnvd7axhPPQkO/YsRzoAW6Ja1V6cGkh/KZ9ADM
NYvc3ruhtxEEkFSE+mUM30mfB2nM8sc8yvzGqbSiQiCFIMJVnAN3Y9Umw10Jjt0eA8wdWtnwjq/z
TmAhe72eodony33IogSriUY3VThwOD4LmkJC4i47fCeVfR1/80AQck5maVGD2qFIx5YeMpUPWi0N
WdJKVI6l4aZX5xdesJGIb8ZgLvsdIcXRa4LggCIKijdTwLXuj66UkZolrykVDGpZBQPcpvP1tVXv
p2M1saNcwrvx/tSyix0eLaCmaTgZl+JQqD6LPmeiroV8ST4s3QGSHfVnW7V7+yIl/xcYFC/nipEQ
gRu3yTa4pQ6POz/V06RoBwXE+SYDriTrL1lNWVM4sG8U4yChpKx58i2X/OrDJCugbNbMpX2f9QJ8
oMYgOXN7c44ar3Rj07L8fyJn4aDX9GGWA+vwF5eQ9iuLvdY5uJ2K27su/d14kfxyspdhYEzb6n9e
mp6673PjI2eWdtb9Okx2LERO3wJLA6UZM0O+bPq1d9B1C3t45YA2S87FYmEuD2JEqAUBkec/wNFo
9sp7jRVerSG078bwK9zCALxSBx5uHwle2uXVDbwxmUvkqtzA76b2TdsOAsx7RcoqfT88lciWP1n6
AcYx7JLkwVci8S8kSJ8aB6uGp1AlsPr39GipXOWQiJGjGymPpu2/uU7QofdnG3ljbKaw2OjCsWNl
nXCSJkYC/SNuXl2M5O/bc7LtXdRLNjRdKV3M5LfLXjn8rUXSyKnR21+422hUHJv0H6ne79gbpnM3
TB4PMBZM9lLBdqT31wMUfpfDkWqJPdjE8n/eIZpf/VImAeIoq7a3BRXbuSM/J6kODxZyFfy44dYb
X880M5p5eH9wF96UVbtrAcQAr45uZ9pbCDD3uwHIDx7QtZ7XjnvyopZ3il0Ej1Dle09t70GBqlY7
1UggWlGfez47OTVIFXL2Pe5YgisDmmy+kug2YG8Xbvv3QCHWOSezTIcnkajnGmnAinJ8wnHo9zPc
1wUc6QVZ9aS5dumvODsyj2QfmUEacfY5zOps/BbF23Y1KdujVryFEcMuUasL8+IN8R/w+7WkF0v0
5skALHYal2cODZZNNQN8vX9LZVnVYbB3oFA+iM9GLiGZ0j1AUFHZ8zJZ6ZNT/u72E2w7HD3Drf5u
5IsGFNqeXNdJVsMYS1VSp9AKFzENyZPOQyKVnvT+yIodFh7xYllQkLjwgGp5fRMrun9C6mRTWuA2
Hdmnijp+VQLHHJBOVjVIUCKDcG0YxPyRyW8jymqNHILTmtuiETgJ6MPGqn/yssCiA7rz+7Hfdhmv
s8zPRqe1MXXsTQGlyAhSCsGVdzG92+AjpFUL7Az8DKUGBkwk0UveNTkMp51HqH4BurEr3KmB0UFn
FLEooUHCL5wC8lWVrX1k0Ks237kaEMjBMN9UayCHrnvw/UrEXj8zvHtV621v+LPKBBV9IKlSC6xL
okGblnBHXQRSDwsZuzXqtcQFlF13fniG794yQoD6/BlAcVRy+i5wPMcDOVTJrewuP5xK/3Kocr1q
/doaAHa/mdVr6lCQlpIv8l8nks2U28hHZy/UAkY/TACmie3hWWkYx1TBVGv85yq8ritfxUDJnORB
WEPJQxioNlO637WiByfYvoqsI8Vm2U4dPRfrE2U/hg4lGdt0zUbp/5fmn5/6MhEaRkcyG20gCRDs
kSWEsb0N+j/yNB+9sH0atCuSytjywM9Zq8HpfkDfsZPGDxtYA+iiu9tiacxfLwqRdNoZimjawrOa
qczQR+UyQmjD+OM0nvyMh53SOZls0G/FP996O0KQE4TEK7XP/GOMicQpeJFrZ22q+VdEVabpeOeO
OG11SN4GNC31ES1NVYsrqtEn7R3805dFfENRoW/gAWBTBEDteiiO8/v0snS869de8Pi28dBbZiDC
0Fqoi1ksc6H1XIOXtK5jOtof3PwCQHlqE0bzwanrNaZTQzz9rCy6e6Mr2Hqcg9FqKak1oUaQNXVs
Mhhr8IA/ebNyQb6+4Dd4Gqwm2V8dNLLFzI3qNuJZcF/iAfEciOMpxu8gEDAFWtU9J8m6zeC2X6FW
xqaU/dpzsDnCxFzoEXnQOm8OFjqTVGzYyH0sBhdz4efCMweT4DX1PhI5mVSMEjOiYmX0FurNJI40
4DLurQdItHN0Ezzjy4ks8AG2qfI9UhrFwqmJTst/5dz+FLqKJYddjOILy3YKwSVO0OoNyY4D7oTO
K0ZqtOvoSGs4MRjOP9HGhwdMGdSl5YiDkaxg4F6yErOoNdDtfCgirtu5JUMnQ/6tnaJP+5Q8RyGK
3VrP47lLxAoW6r78Da6WfgBKx9/kdpWL3tAq3hGRh3cPY8d7C80j8XgPBGnsPm2ZidOH7mtqkKPl
8EfG09/0Tkg0KUBzL8UAkJlnTziPiJSfKf0rHIOk6OoUcJp3fLIFEqopdsbIaQ0HEokaVhtZ7woY
ouH8/kNiL2gPkRQ7hF0+H5Mme5JElzidWTXc99qF+Go3dYhUZnnOJyxAYZxkDziOC7SkURCYMcyO
oxD2HlxjVOsjm64XWzczc7wysRD2QfJfLaMkdtVI3LlroYHFjnK2gZt7Nd04lsC7JLim/sITONRr
z2TtQpN7Tp0uDcnTDQowf6eomwJeVJ1QtcQPddyPLNEuo7hXLWcV8HnKekvPxtXPANSNJZCvYPJD
2RhjiwLQw5vAETdEng03/iOBAPww3BSjeKJBS8y/tl6XPAy2ojAk+7R0MoxhQlGHFyyBBTfeFlne
JBsXLfXve6rixG355mkawhezaUAiY/MP7uWibLrleGtxiT1baPqlfolR0hqhLehE5NWlAA4BS0al
LTgJD+gZ/mtMBasXD4iG+rcq9zi4qNvuDfrzg0s3wBLuI6cGrzNQyP+rjkFAA7KbKUZ6B4fnNMBw
Polx1oe+7kfHK//xdYEnBany3uk90uZ1IJcElcbobCg8idRF5pvRR3grmYfYpuVxnloww80BlXXb
7s83XM0H/qmelipIjEVrp4Z1Lv5hAvEJ87fXY4JQ53tJqCWKxs4SjF88E28vQ+oHatWXX9emduCM
joUC9JEZVStYXjhz+KRaz3ffSJMRRVXV3GpYvd/gB/yza4UKLkyHtjqpdloe6uywRtkcHtQxS/Ya
0sVyjSO7nSXmMmzOQs6StHNJXSYyVPcWWceNJFViE8hTJp7rTMSnTLnovpLpkll4K4D47PEXTdWo
A2blGdj87V5QEVRuUvjznj7nv2U1DknIS45cSwGx2sbtd+o0/ezPaKpIc13dT/WQ3rtTc2pYgESD
SNbE1qbfiiyX8RPiWAc1fIHu1kFc5T/TjAi7tHc7fV94pI9FekcJ0PvezAbPheALo+hB5dhKqZ/K
pevuV9MkU7LILcf669kBtF5OFsWsw1BxtI8VkN3Gj6pHqrDqOn/Do+WA/ekucAi8YIyyrzZfKbiE
ypwn0NaQhXa4GC5vwAOWZLOmqpytt4eFicfqaOU+KLPeSl+C9I0MaqJmn0VBhdAUpGv8L5h+qNx/
FOLt0HXKkvVqCsW9rXBTcJWwuuXpNUgeoqDCbywLVaUNTkZWRAZaxUDj86CJMWyI+X7vMhsZPllv
e0oGGUNwVvL2lNLYciOTqGXNWD0/GENf/kxBSIsjf9Vc7+GTQ4t/rq1/aj2DKWous8G+xu2ugjIc
O8pHQPc9C09WQc2LQrn2xbuNBSzILNZV2ggG5ZKeYTVW04jKgc9BQwWWU1ICDdH4q8Nx3uNbDVze
9iXT81J4iMaMDWb59hNQkJ43ERPwaCXIzUrLaESV7U0i9pYliOVb07eAtUyH+Agrw1akCzH2jmfa
1uj246lPPF8C1iAuekOYpsslGdVMvdN0ap/7vp+GtpSxQuTtV37i06ci9utJv2UpHlt7P9V7mWTC
B2p4y218VNReNYmkFxrbYUiNvL00vvjFgCaROMGZGDskgJ80q0/zLGhe3wfTjEJPEeS5IFoDC9wJ
jaECQDenXGc+jn8TbdYHYyBxiWJItzfPOgrtw0gUy3Cxs+SiI7KUbWG4HbgerxNnKPnhOtBOWaJJ
3auGW01bPYQ2yB65NkukNjKxvD3WXl5HEBiZrw1bMkbrARec7hxASholjRcGw2mWWseoEJX9Jk6I
29aTAE0tadD4vEJg/o3tSiVzBCnze4B/plnPpfq/m8bzbO399VjNg79eyc+IexsFo+1ZItwaxOSq
4b9iL1JYbQLyFMfJE+0wSz/I4bdR2bXYpo/Jdse2KxjyDPoT8tE4q50gLagpfwpnVw8+26VVFTUI
4Gtw6YWv1H1GfXCW7jVuKHXTQ3+qXtH8u66TcRNmwI7w/FnbUYJTdbGWNYLNt6la8WDbFQ6G/gQR
YE4UWRpULSjeBQZK7I/dzlvMdmKQiGYFyAHDBSni9Jic24LZBu3ORvU3FLKylQ189ixzizjozqVo
rL0Tm8jUpNQ63l+ZbEMu8itck3T5ASR4qNvWMYSr+Zg2SMHlS28za9ezP4IPNFerBsvUr/rYFwKy
IvgdVgOhnTaQvvs07pXGdnq0WZYcVD4deLSBDloym2MP7HAao32jQ7zUmphV5pfodOcO3PUibYG9
NLJWpdOpBgJ70YSpMPj9Z+CGOHuYCuE4MRLQsuazbZ8kuP8qaBidjNSsqy9qbisepCyoQr5VWfgO
yPzI3mlEsGaoTW0dyYlwyMs6GclI0fedNXshwG18a0Lmr071Z3f9NPrJYkzND0Fku8FVgTO0yfO7
bn5VNkMX+WqPFkcUQXOkzXYGBOLEhsRXxN4Ee9JoHhTa7J/O6elUf8hy0Mt/ZalEZfDS1CzGNED5
GQKCL4BqDY4HGoKZ4eqwXJEXMuFaartEWF2DYVGMC9iyspmQL1pA8es2+vGtA0D/0gCoUj0yx7r1
MJ0vhmJgm5AULyu/zx4/qZgrUayr5HCDapu+kdSgYeyXUHXmq0UOWT5yqrh/wHuI01IiFYYPdPfP
9c0f2M+ttaFteD3fQ0HrPFf5qQmRUUPTIE/XiHMYUIyyBlr4tULMVF+MFoI/75obhudUi08oH5Lr
JvhyV6yBJ/2uV2t0OL5NuoX+IAbTyDbIlRuNHU5QLnBjdita4opbM461o0u0McKidsCY3eGjCz43
oXXE5cSCQkFTyiW37gyeZGuIf9MNzyVbffkrhI4kxtc9DCCLOVqW8fOTDUM4R6GI5mzNAfLFMpfC
RJZ0H84/8oKindC7rkkvqtJ7wRitru30fv0NVzmmVM57ktdxeoWpIPJU1kc5WdqEashWwBod6Vtp
szhYHUR/cNT8rr/T2O3CXBxb9w+KIo7dLP7TnlY3PziBGZulUM3riCyTdAYVwQOzc01lJAjzeAfz
ODObYTToHzl+0QXBbzaMmw8Xm9eA35g2XvX6MqzjAprFWAW/LBnuiNNKkAUm3DQR9s+x9cFQ8Pf0
y24NVMu0SFg8knggA6aHAWiUrK2o4Yk4PytLq2xNJvNbe6sJhH95Er2YGrqfcf2POCZS5cgX16Gn
QIlnkuhbGHDxgNslJQqldGwa9k2C8zuDXm/Mp12CyXlcpltMx4qQDEu75+w0U6gQUeIAAH/HNSiI
3PEerWKOsRy2PeKlbQZTkthPc68kWTvUyQoa/gD5HNc2RSWeu1uHB3Zpy7YhNto8YX/ui4Lu1OsK
IJiEYP3n1Fq94+A8mzpQ6IOs7spWTWTOLQucgIkyO+Uc2EgNS+cQu2foMUvQNEnswVBK/q+NWp9d
dhCvc3PQHeItDcK6VCauoyInAxJz1sSPieaclpOmcth5cv+otXXgVWOcedmT5wIfCIJWUMRhaQaj
6tV7JRQ2WylLRP9R4Pt/1WHo8e5lIYrtYZQ5wBHrjmP/TUEJ4NtNJCIz1daFe7H/D/XaC3fb36Yf
FjXbl6VfSEevF2ljToBvCKTZhywjROeUnVDkSQzYfvwDVkpxP8TM+paREcCLeJUF1371imNdM2b5
l1+jGhF13n8k9r2ZO35JDquT5PPT6c+LXL/pQ5LKkEKVgyE/Wv/yehabeitF6w7SQOjyFFtg3wnH
nbEar9zA84LmMJdSwgKxXGIKzMjSIaZx6A/WxijOhk37PyA7lQ5z8LGj75klM+T8hftTg5EmrNhW
SZgzLOtBSQwLq7UVdb5mHqNFc8oNfZzorM8c5nsJUe5F4Ko2iPkaGAwXAMzRY51Xx38AOw1t+K7j
GPKci8FkkiMW+X9HtolT++XEKIQUhgi/k58xvCcbqge1e5aeypPainPpKwlUmn16gTGV+vCg0eqM
7+7uHFvwFAuZEpoYSZ/0V6oO0xN6dIUHN96YQNHpv6uCGZJbV7Jc4LMsWVGj1B7QmmtGtvhprHYU
59zDn3lOW1ZzFbI0aM+CuZ0nZpbUrVwwYOGiDaO8w3QcsovPLa+jh1BIQc7BN5mtqatUunt2+y2N
iQWkuWihs34VUR0Acn2JKAszmIrFaFJiTevZteFneNabH2+/RrBDrqqZeVLyQ4wFA0Y73PCWSyeU
cfUvcIi3dIRe5rUdH1Im5lKWrTFrPun7e2sj9u3Db7/dEm2Q8T3AIDTMxQvhamyU6q9q4SnQnXvM
G86GBvMPeBD0kOXDcIeUYpQM91oeN+ZeF6oOwPDU0yaCU77wzpDxEV3fFb0Sq467QVoKw2GhDD/b
nIh0wrcUs9jbJBs0iYTfBPSajANHRi46q+6OGCXrgimslrM7nCTcimWU6jyYPf9hpaKlVMqahBdZ
CtcJPjOrKnticr1n8eHHy/bKrL9ggILlD2CJu+zqEBJJrwHnZvSQ0/TfDcjeG0h7CgLHmoTzrhCr
5+xTq5kR/R2lcjCR2+ffHkqQT05oZGDHC/VEBSmV9QtPMb25NBK5ESnk+RUvsbGtQLHLwR1S1XjK
DCm6PM5gcMHq0WIxQlrytpOJVg2AjQBGS7599QlbtBk969ptWrCi/7SD2ZTBIdNrIY1XQdlPwPIQ
Nm6so+PBPSxekHB4aaiV3ZW+misgERFyjdS3yItlb28k/xDTmjvkmJN7iErVG6pgfo5YGIANBxLk
GEplLQaF8igvwcHb1didZ1GBXDy3T5mWA/brhAn/siIFpWeI3AAAv5J+fLcmvTaT4TOlisYLE+ji
SGYBJkx5Wlc9b9W+KZYKp4EJSTja+ZbPqLneOIlqiE2aRBulwIfMj2H1ZYt7lRDPDKDzGkjLEWNH
EcwDPh6N3dAfq687dMV+kyB4UY97iGg5FO4ufmg7hJqHvT7IVQiKASSV5aFKzvWsGPD4fprCvJ31
KvnK/7ZDv0OthuY9RdREVrdg6XSiHpOW+CV+5TG44xUaKo5ntSP5B5yqOECnSEzAtxOifNZrDoKA
M98OBAQFoXjKhcPodQt+Sxw5K4obA0HGP8LmSdeko/XJEoadCVCXWNTyHgsfzSwqaWJXu4CpPIBD
mZ0zmD9YrN3XPzRJ9xlCqWsVB6n8XNuLvpUx4acUXjRwCsr0KUjwLSnF3ykN027Og1Y0u3Lr4gFE
Oll94nKA6HA3BVfIW9vFfHuN0jeIJB6D4zSWE+4s8MVvUQmpobBWPlGPouSzFCxk/qsH6jkdUD9v
nFzgfO2chhQ2SNR21i3MrKVAHAhmoji4pXzeRvqKFSmFq0Vcs4Z7XBlRJjI290/CQS6+iYP/+eqA
5ZI+2YNwLRsN1KkljiBz/zvAAXm+/QrkU6Fqn7fDQeSIIGrLcUx77Wt1LIMbIOf2F5dZ2AE3DZ5q
B58yBmI+SmxC+TaF3DYAfY0lIED7h2toHVo/3XdmxEYj3JETVXFRuo4tMxjeFha8zFPiPlQ5ztH5
a0SvsFVSHiPgPi+Orb3wNNCXZwc6Mr0ybJuW9O2lWfTVCWPGY8T1iFenJ1hmeiYGUDqWb1Q/Sfeg
EC1W9mngBLqcDCTtlcfSgnRk2avX5oNhHrujIdVXolD3XN37SuB40HsFcQ5W4RkbDgp9AAYv44wa
6IEctPEti9NaAazbSIjnRawXAhAxStkzoqtqu3IStBW1De4nIG4SL3ot26x5UwmX+f+qV3/IJvcx
hrarnV+1C/oK7vWA1zq3SEnFTYNjWXjCvKLRrbTvH6fS52y0CQY6lcvMediDkWjxL5ypdVzfTw0Z
eqYnWElxuanEv7iLNhI8cngs8HK5pf9zLVrx3AuRJ1LiTcFEqCqLzoeEx70tOle5WHoJAMhWhrSg
GYd4HFhikgOEp0HG53PUmJfpit96h37vJlel6blmkP8DibllhyszXqRzTDQ3Mk8kegeSBYTKfxqf
l7tDbDowXmOG0p3rdFdKBQ7swSXmOdpNzKH/gauDbR88APggjpBD9kIn6bBSiHT8bFsd8ui0BM9P
u3sP19wY5r9u4tXOtRZH16aFdIZBkfUwHGgFMUGHPpuXSbuz9TVUokWsM/Jh/ui6YEJxfJEXkl+k
iR5EAExTeiL36tF7Lhjrn2V8fOCaE/W0mF7uY+A0xOJEPn5zuoMIZ3JTb6wKypJqz1mjV107yeZe
1+85FTmG0MeyHKSvemFBVC7cyJWwCtCN+0JSYGPeoUCMOUr3e7Vvei0Q88xHx1gA/yGE+wacUzie
wr47ZjdG4TJ5j/qFDbwqpYLOXJyvM+yDe8zNJ7i9TDCVXlmUATyQeSVCg1QAeI8oTiRwOm9t+ABK
lWdQXKX6U+gYPtNeih6tjftnZQbr8VEVHrkajuy1i6WtvIjiQOD59+hSMG1K+5474b+7Go76h76T
8F9ScGMqZuxBHA/3XbzwPmm9FNuQqflmZHWC847T2jnK3oJ8luzY2Q/n3gcP4wt2QNJu8t2ELpSD
ZJyAXyhHtBkoJ5L2CwFV1TgxoMFfco5k/sVAfLZAARmzLHys2d5qmxE+ORKXe4d4Tx2VlNC7TYHS
jw5+i9DbrAUfUWn17BjyuJQacgf9zatXKb7SWjtoCngWlSlCAsTtR1UIqtPUJI+LV7ceiGzvUnKF
iWZi57REOWr2icMsHKXGs3mDZPB6teZl/+GQAaMDe6nwudhpF71YNGwPzDLU7rY+7Pa8XDjmZePB
iCUHMKu0e81UvE+1ndhNnpJ+WrFQCQVHxJ4MnxRWnhUKY+EYuGC6gyxjKjoCw/Hp3oMxNPw8Kx0R
tCJyhjZwejRKWm60ISJEtopDHx1p6WcJjlVgWa/erVK5KDKpb0phLaXxy2aiBcD8VDmaWQ3jL8pc
8j3PrMDXRGPK+6uP8t8eAAL/ftmpJjH7rOWn+pPUP/58IFbov3oUs6TWribzXEUlrq1Lc9QRQA1K
AQ2cWtnNHIPPdEoeExaz7JGVZfqOltQR58HLsVnPgESB2tyMLtaJpyYzpcmh2oj3/MC/Z1EDSKeX
lpTp6W0Pj88gKkpPPUHZbx0CxfwifeHZhSxJTI3Vw78c6JSoe2/4qfAsVn9Yni7hpC8JVCnh8ZT0
m5elrRb5mml+rrRJyf1lhzYIrdvmwZyT5wdtBjHopL39NReo+Vi2XbRB4RdG2mEftsM1ifvBQw2Q
ZDm/gls5cDnWJBilSmqsU6srTXWVaABsR3HroO6HQ5SAuhIlIF5E4YaJhdruDEiC/G9iZqqrT4Vl
aibfgg/eow3OX4hlPoeaEHtcNloeFnvT//EknYmAJwopSLtPn32xC4Ar2FpKwMZgXo2wKW3wywEq
hKsbHfOaURc4yooTtS7iUMd9u4ZLBm3ZcGZwxA8TnhkvU3lEzX0Y2VB3OAeBqLjNqfArUYKQWG/U
wd71kE08/QBz0+oeMLN9def557q7TgejYcxDOPJXnZkhsI3yaunZ/yoYnLbgG/vJbLHdqL+0oudb
A/qbyXcvknj/fw6FRHGPUM+84ruMhpvMcYcxAhnL9embTNKk0jy021o4mnmNRsb//kiNlKXULvXo
lyzHeaebtA1/ARCDKoeptHfqUy0hKW2Ula+QnsU0Te9wy0H8v4QZqimpLBp6pd39IDV/+ffHDKJH
h+NVJ2Os/R8q0ONCu5JTODHC6i6Kg+DLBfvVg+PbHQM6Ung2dHqas9ob7+z9cNyI+HkTCaV011Pq
WH1FznwpWHWestHL1/Gf2AlT/1hUDiER/zQccoIvjLPu1dugGBj97qXB8ZU2fJI7at70aRf0Dj4a
oQf/1BJe6r2CsqZnykJoKbuNnJWuJU+/F4nT11q1tAcWNAG843BizH5cpzx+FQlJ2ZEmOwjXuqIQ
wTYQZz3FSxicmlilBYWLrgI2iyG6jnFaCfKyEMw7y8CZSyABx/ZgMxyT9tiToMM8VPdBf2da7iN2
Kd6PSjva7RaPRsloa4IW9YsSQ9Rx6dqSFgxfmLKRbnjTk8ZHejEEwugqHvTAqIw5Iu6J+JyzJtRx
ZJgbq1Sw8iH7wQ1DLscCulON5qOQhJNmVgzHoDxwLGItOncEsRIbhjnHW0aj3Q8rgEzNhd+4ur8F
zsMCaG7XdBnIXD1KtWSt9jkBSmYLZGpK7k0EG3pKpzGtEtwZBK6FBaeWENOtzBzi/o8rGdKE62pT
j7c+dSk+j5updMMdfcearT0ysn3tbAKS2v1+rhzSXWE4HVc0KpCFHxklIBuVayqH2c42x2o98llO
qRXwyAih87aCpDRHlRixhtQhIXoSCGe27NN4rNdQA4YUhxuQgsvyL7rer6HUlfPhvOn3ljFJP6zH
FJOHvtWsFlEOXh/MKtRocm7J6l5SQPj7/v8WniX7g8CHkhmwRKc0ULGnIl2cyzTIdhyPVTXyrTz3
Mc1SUBvIfcwkyY4ucN5HwnAe40bauPPTj3BoeLnhLedgw8Mn5lu2M54iQrrQGzaxgGCjuctD1ak0
jQBh/igOwvYVdQzxQ1W1dBJI8UP+Fz7k/AVDQEOQLKNa2bS4xq0N0G6BXmfh+aUPZBPw6fO+rjTt
WFJ6c1S7ZuBJABjzqNVBqbZ5Nk8m1L/7qgcy16hlou8HmlfnJ8fkEzcb8A6KbpVSoxjM6KnGRHPT
bEIbUNJZpX53czwe61BvkVnHQdVo3G+z09CwK1JsVKVkRIqZrs2tudavDNfRhCjRggHSKXu55sJg
9fLalICRZgsFfhB/hOSPW14GhLlgUdBRAfbth7II69PD6dxjdZKbkYe43jO4mBuhDI9Y/w8xYq3A
vysNgWDro/JJGYjn0+ryN18ss+dZkHyQmI+cSxBMtl6ZxqJROJuCzF+sknMf5LC9ZVb1DZyGduQb
G7cg5/zONJE4MJCYkAnQl735fltg1+WSuLOFchJDKg4kAGpqec1OqgFm+C0VRpTa5wMdO7Wiicx5
kxPkBigev+yIbGq2mwRFfgYjIZQnruUwELjY8BO2XoV04Yre5us2PXOX6Rx6vkn7yQo0oQiGxrI9
tZkuRWah56Xig8lHcbGvTfm1qT1O8i3KdnENITp1cwCflXU80JLicR2mVD65SfBefetZN2KElvIv
Se3DsnhdkEHyoNZzujYFKKgjB35AcXMUvcmwVSAGXmSzvVgOpR2LZrOxG3VWxTOlIs7W7+wrBhgC
xFpcnOjOBqenqH8bA/Ss7czU+lqrvWBKOOfpy4ctueS3aGH0hOYjcQH9RHtfmeYO3vxVaAZh8FNh
iA06noQ3IyLJ+QHDRPCCeZzqnVh9jygxsWPOzKpLbNDGBeWmKqzTt9m8gQX1FOrK/hPWyxXBXAlX
hyQSV0T2eB6LkorSNbM22nFMPUlnu5ZT7awLnzSYa4sTPg31djygkLXvKVvsM55h3GiHvErhaGqA
+ExjN4D4ec6yZgmqHy0Tm9OCqXV6N7kpd+N3X068MEH1z2vC7v2YE/BiFiAsWQVBTJGvYvpfpirP
Xv04lw7h805pJxO128POHK2yy1FIJsmaeBSsOE1tkRlxEVDAJLgPshsVHRHv75lgcoSv2KQrmITm
Oklg0k0E94TH36UinYAl6c/tisIh6SPwP8TaJPt8buGf0Q9g1hepuGbyI3BmdP88b7GV5Xyv+w7K
iio/wQqtYT3lIT4bc68KylGKxYRaCqV2LCUsSAZc1K1Owh8BQlGy8oUOSpNXZOjvpCrM3rxD+OM7
OvPSOZgvrtmvlujYpfrwGkkz7fjqlvy9kqL/VSwVwsfwUCOJS/HE7y19s9sGfshzb66h5xoPO2S1
w2/DT/R0jbCnspFqnn6ysDgAotyuGWFe+i6MhkLEhIfsTC1YZFO8+mmDI7VF2kXkbHkbcs9HxEES
RZEjELZ7rXgyNnCPiZJrkyxFoV+kngmxYi5PlTMHi98fUXvMhDtFu+h8XD8FKsZYzuxmSNi6Sv93
GF9Kn86rsTD7Re61PBnSOkGtzVzu8mTCFFyeG/U4ZO6FbijH1l3kvHzwIdWDkfodynIfX/qGVNVI
mKBjHpyx2VM9ivldZNWeJKCV8yc79mhnx205l7PSCWB1TDiY2qJhJXm5VqYXmR6i4x/QzsOBT+Qf
eVANEiZRJfqxUUMKBUbVvuyQ424lASw5fhv2+OKRrgGEytVxPMEw4tdPFRX897+uRJR4ch5clgSH
oWBZ3+yH+qeSZgis91shHBWhmmSgoOpC1IvNNqvb6hSSu/2VaklfKnMP4PaITZ64CRkRsKDMBlbl
wap64DpeQW6HWtXOFTL7+lUyXqyuiYuQWYlIH4MJ/kUPAisdPiuCPKVxyos/+RHgaaBqISNSnNaJ
cWuLNIqjdY33lp15wxU0T8sjJ+Op858Q9NteMlhowQLF7ALWxbJQIS/7CpnTHy7bTSFD5KttY/Xa
LFYVvokivjwaHlQpfn4NsT9qfW5pvX02F2BN7DzwcZW0zJwwFn3FuYyj6XGP+iX5URsje4seA4UQ
poSAz+xgH8xaTPTDinSGdHu6YFCgDVpRpof6t6rBrNn7+12eL95o01SiundLLVF3XrLCHMFm9VAq
pgJRRQ+dUVjJGZzcjqZEzA52lcRFnbAgj6Mj7kg2Uoc8IpHEQxSCb3FpgwELJecJsJDQAHPBR1YQ
k7dhpxUrI3mFjMJ60TZyyRp2dJTFDEgxPlZXQxOOyPIAmBosX9dFQGFXn8K4YSJEw5P3hjdgSeHO
hLyPl/nEH3mGYZ3rS9uhRk3+L4f638XRvffCOvMep4EcPnuIkUQvTBoZG3vtwgJPxXb3m8Ho+hms
7BlFbNzOVm+l6L1lou+NLHTfB0i8ptvj8fMpcCFawdlyKwKsOh18N7EdUZsJNYgghn5lIjpCUCk5
T89RialLkOuMkmA0Xoql4B5QUQsbwWyD6nZFuT3IGgIxjNqmo2cW8wmj/Wg7tJHbZIFY+ufLHjBP
hotmFB8XXy2kDi3IQFMUYWZJJ7HDvkFH2D6w3VeU5ffKenK/WdYHQQPrM9t7vkbiSa83zjG7p5ZH
1xVDxZI2owSKG1ZUvZFOTbkKZlyhd+uHQzbjb8w3hdmix/w8nLTZPf5nN7+EzDOSvJBFB7BoVGNI
p+wE/AYNLiC/IRWVNqo0bfMKLth+X8uWnDanacL5VU9f7LBpmSOYHGwzy4/4jzsmj0StRc/jWeK+
VjTfQ3EKqiD8Vq4n5hxa+qVoDGm9GRYL1EZspo8VC1jCF0I/uMzbUDDWwAD1whEtelz/uLv2FYsl
NHBM6sbOXt1/QHHOXlITzS3ZZDk6WY3SJEbIWkZlqeR8U623eNwqo2Y8fVKP6g/Yg9spbQ9MP4yC
Ql5IxCeqTpBLyQ4wZOAjMM24u7g1wWgnuxHmtczfaZ/B3YeEd3DwGkwlDqU4/cUEIiZf2/kcxViL
m25hZ2rPJc1Od3FuFCz7QbaBFHZEiOurYkZ2l7vBSV64XMVwAGGz5ep2VDTlFszUqKjG8rcANnQ8
jtRsuf5hZMKIJn8+r7MVuZcLp8aWiSbaB6tybsDYqLZIxw/dHQsm+e4DxU3PGvq+78pU+SbpKWk/
c/II29zB4/SoCYAKDGs0WBDgGT0V81piyaKHvQPdkJ/FYdLTYbBU45iHxw2XDpRL3disT8MAGsZj
MInO7UUVzdl6VcpdUsBOTzTBafeHgFBbm03szer+Q6bBZYimRi2wqisXazHCyGv/6PUQMYvunOvt
cCoxjr7SeQB/hcjvnf7s6L39SVl2oZnkZ5OJk/9B79407vAwVSFzuqG+mLaebbH8RpuioCEjVdB/
3ge3B9GOiHL7KoLbrPsR/YqQ3iUrEQo2tMUypOAcvBsSfJc+IL4m+ejGV0Iql6pRMA//AiEhyuWQ
Jn0g4AD03+lEtqAvmBf50tMD9Ak/KPMsNKkHMW8fpRe+i6BYfYK490TYkhXR2dz5tAOj/I+hCez7
JWSmUrG/ix5/iVJN4cQzAc5XYTwh0HOE98CGEjN6e7Oyk+WMN8txKzkCBAYEvD1BUkXmGSJuhvzs
U+EnqJnw80WwS1KyuCHaWjv4JBYVajsXK9ZZ3sh2yrBgzxVfdZLqaYhbukoeQ400zd9fyljPvNhD
hJnaiwqLJuDdhdKzB7V5borxh90l/8LsNKzQdPUIx7Ua+xMUkndR423p/jBoVbLq2DcgBo9aq8QC
N8uiIDlGresFBmnfm/QVBV9kyfeP9Mq/R1wJGUiOHk26ERAJINfkP2fcmZU00zaCfYaQTKzw+Iyh
0CPXOp9JvYPKYP7y8oVzhg+BAFY2Wzd31rOeZQxN0xb2S8Wyi+cOXMWD+E8PQ9p45T++Imcbz89x
CiTlw4LH6VaFct0pdxij3vWpxxwIUtYoKcgB3sUUAsA22C1QmK2DSGazeLpv5D8crbIqOY9Kwp7a
oxRFtfi/mr1k2pIADMFGM5X5ObQ/RMU/Lg8M+jU2WN4UXn4OhIuxnJy9ca07Wha+rvccAdYiYoCF
o3g6OAyOl76fMirDdTKEGuwlayLzUstXd+wjSvVAr78kDkHFp3NSJVWaNP45e6iz+G1C9eFrZBN+
bDxhfRGV4RJpk41VLAGkO5YN9qKew5rwJgMjDTmyELhz/HDkRh2QKq/8MiFbVhPdbks8kpOJ0ea0
owiWSoOLSerQxxUO1Y5j930RpoXN+Noj74wN4N1qYRCkeKEM+exfaH3RLPGdC7nmIDMYML4XjXWu
JN0cPd9WTUj/HzZOglq0GLplTb5hDfuUzstvUDlCPazUFZByPlG49Tt/Gpk4+si9ta4POcLSWFQz
U3hDt5kxlNouFv+vrU+F5mi8d8aZqr+S274vUE2cGer5VfnvCesxmPakx36RWcmmOCWb+uVgpPvr
5uz0H1siPxeCvtJBF7ZLYs3qyF3GC3vQJLPJFTpIUWtUXW+ck+Q1DFHQKUxNmVJqZ6qajYxojQuQ
yXou1vwTcox6zXVyTcTuV9kz2ALRe3tl/iqi/hNO3KQnz6EPtuAVZDkk7t3q7ylAkuoQuNX+PcYN
nkrc13nj97AQsD67r6SsJp+ivE7F51JifVPJnWKqR7dsjQY8O46Z9xevTxALSzT9CwUU1i0eD7+1
ohiCcv2GjmX74j7JrjbbtAZKVKpv9IQSSvGiLDPcbg2eUNTlZbMsuxIScrVS8ad7VTaQdBtGF5jF
zGLJCI2teHK9PTXf55KlqQFBQkgSyFB8o8g9qK9HdDeDQlUUPyNIg/CmLK0bj9czVoRqjDnboHvw
K4zwRCa6SzY8zSQ9Me6CE9Txgdeq0GYNxrJ6SQMR5uu8xLrLnvNYcjcpDOYjInD5Mogp1D9LtK7Q
EQomXB5CsfSotyzxs2TYNeco8rQKOQKEFthUTqHXeL4gLUWGoTJIkJn4hPZR2jLiUmORBtVGWt/U
dCV9EPi2R10nHgLdLVWP12Y/RC8zNjsVoshfQ8WMJrIXRUkN5SpLFe5PAOuOXzDdmpgV4kxQgsO1
c0KzkvXVHmPnRxdiZKrKKSP3ELrgQfmcYI7y0Q2cwPfJTMC/7z/kl4OyNlYeiZ7OXsVzudE4GqVd
4cJnM1e9POV2mJH4GVZtxO3e/xRL7+yQJ6Wnk3TMkl8mW/mkRd1mm53wi/e4rPhga2ByHl2NrvGd
LWiVxKQZBYEymDsa28HbS6PzitukDlIH9m88xFBFARne93JBa3AB4/2b0tX/QhNRxSnRcNYJxO2J
f77rMr7YA0n1cV0kvxU0Mqs+EKCOIUVM8S8wvJIV+tbwfHDv5ZN+BQJJWLHoC9E89SIm2EadQJvA
XRPrjVHExsxpp+OTlqckPkgqytIP83gA2t4ggrTjwNJzBsPt0jEZq7dOZ+Mn4t+vj2Uc3yU48JB0
Dnc0/B3h+UJ3UIhyph84dbJlIa4nNTUEPtwDB4Y9D6tM4bGGO34MH65mqlA6uzg/cprATSzvP8Hu
OHVSlBpQL9lazLrOmX6/7ny/LxYphhB9fNzQcoD1Qmwt/T8t8F1iVb/lw2wM5iwJq0g6JtVlcAzQ
tRFOKosiQqQeGGtsJu+Cv1xM8ujCVWNliO+CulG2RoyUo/EK4pii7zVKhoZ7+y5BwHKCxtWZraOL
CTcyyWsjKdFDkxMNgHCKRXM9wQAbWVe/kobgHbKRXFxh+bijAogRJ9rhpQEZhXOqtAIRjNsM56p7
KOnvtN6ub7sNY4k1TaekNWqHiFMHBsM0KY5bAYMO2xAAIQfvndZU7K/TYq0LBN5OEpbdqYuHLfYk
zqKraxv92xZURdmVgV5ijLqXLt1pCusaEtBULZMyn6n4aBkTpLx28Pwe5YFdZFs8UTsm14LQx1cF
gHbB5bCagf090anjmdll+4yPBinYwV7JbtzPunXFJydJAQEf5L/1q70j2hsn6Csa1ZoEsBHv/dT4
6TvuJAAds/4mXSrv+CZxIeROLPacJo2mpWRLgsx1JcEgKt1IAjUytIFgL8xAWkvE2uI5CiORTRru
Z33PuGXEtoJFUeNsD94K5VhBgdSnIwdGxCLU/lKmIqOHJqqrXojTQWsVLlfoQN5q6RgMXaOHnqaF
C/zuTiWXzyVfgCpXhRgXdcjodESGbzjdr5wMcuc5nslbOHZ8vpi5unZPJUI/HAc2I6se1LttQSxJ
P7PSkETWD/T1guBYY3yWy0unOQhRi4pZZsormYOLg/piZF8tVRo4NhtyggSfXLcexCYhwO2ZkgMu
2K95AUgJxBy1j3SY6p6eoqRoYqDRMzTIABHsSP+obpcMjhFXBDeEb8Y8gNQDCaDvlx2BCLOkAkDV
huuB5WxO8VKMAu4E7161u2daz5fIxj2tCk1UF3JSpdQ4mQy5w/IsX7BYjQHiRD7RQozh+Sm43Lhx
Fm2qAYUdlTSdUdyY9G0POSOzQaUlervWgij4ODkCYk3AL01rjQ4hYPuh4Y5Z00EzDvS2vnTZBUs8
L9bGcNH+LBAg13f6P2yB/SiO5wYyYNepAmkjMZ9xaGRs5aSvFDA1GSh85Yl5fsUCTlXDVJn+sM0j
pse/PXATWboBIeh4MC9LgPBNhmEWiJ97n6Oe60vY6mnBTIKmZvB9TwtJRfxbHYBuy9dCkEMm30G9
XNhx0dzU+UTK79QYklFxcxslyN/qF/SOhg+XU7Ei4zeZP4X2c/dC+wvPp1RcCrtDDwCyZOi7b5v1
OT6uxVNqjY+fsLvuJ1NLbTsWbF5yMruFIMBAqzsepe2TUmKdC9R5IU48dt3Qnzu4vUwrnHkIx9nZ
q3/AYlQ190HSdvxLLnxh8SiePCOvGBuqBZd1Zt6jJlgkBuwwsTZoo1UMAY76ZiN75dqlyseaiIY1
gq7+n1euBGqKFvSFLLiQGkQZcTu0svLlPVmc5lP6QPGJKI7DZOrYODcH1QSlFMY2blGQ4R6lIA/I
1zt6493ajNhR2K5+wSO6jABP5tzuD+JF/wFTCmEAlqYHpIDZWGPj66q/wwyq5/s/WHYY2ObpgVqr
rnPhgcCd9tI9Bc67PlemeiEuOE0YZ2fLc32mJ9nXFJrjoHnf+Wk2u23NEgWwR/QJAZCIEz7rr8ma
K2XUElhbyJDHJ0toKhj8jp6ymZriG213i9kZwsvl602eJNe+/NYL7QDwE8XzxnL6/WOOE8URHg+g
KhHjnxxNXtvYhpk15xiQao2WGAWzUkrMwfnk6Cu86FYPdGvnx6sL71xhQV1Zc3KvopwPGD4ndHKy
iAtgRj5wl7I7vTra10Tu1MSsvN5cBp680EnqQ9fOnTH35P7Yff21QDFSIZ9Mjpe5EaMxYkOYllIe
7R1T5q6vjMzo1hdRUCSM8bOGMlXCgycZEldLl2jUmE93qH+x1HLsS/poizG5Uu2n+tDbXU8G8Qcv
sUOJvkobDm9O6i37XqWgTp8Wj+Dy/5jmDeqRC7AH3OT4xz+JcS8xoT5wSbyZPeJ+T0ryEBpzh6MW
UB2PfIwvk5cMBbt/axk7lAmkBdSY5T9I2S6smkkeSnNxaT98Lq5cxctgTIvv8xX+o0eGp0LyM08b
MvHbT1Vn9X8iiB/I5BgDpGbAJkypcKekAIONOtCFaYl03f7Au+wMlWCoK6hxKLY0LkftnEEgQgc3
asfqxJ45PLjWmbCNMHrntHKBFdSSw0eF0ThxPqkEp9961nu9JSJZIdk9/PG0W09nG9cXf6MJ7My+
t52Y+kNIkloKJ17UJlKPw4KXOflOtlHIVFaGqFOd6x7trnMKmQy7FzmL7qh96ws08G8BdQeYDLOO
TmOFYAM5vP5qFrBot/ipP1yitRRfwQ+z03qky9agawITYlue7ob0KzCKwWkhjiewaU7vGZYLyNVV
F8UyqIBYG9qKo7tH3mTsjY1KFD6vjBobFOFZqsf2IcQ10G+9cm/LdEFD1PixvqWEwkDJrZQoa4Uk
7vyCzeX5bbCLOp74f/xMe9uosvoUObbK6UaiwAkCQEklV9LhXQd+yYknQuVEMiZMPFPP39wIuar8
B+5WThZAhEisovWiFCSkOZ9aA05cOh6YS1liTtDNIDIoC2FBPjqPrTfaxbqI8HgsCeCzQy4wTsFr
W707ZJK6DbnHoDX+/FznLrq+TTX/ibwlor2zjvbZqdcEiN7bsCK66gFeK/eeUNGOM7KqHL1+nhnq
plYBQYzVkB9k1Wm/GPVcIrnea5CskL0w2alYdWjdp7RN8SyoGhudaT5NMHvBdU2r1YPjEBWwr5t1
TVf0UGpc4NCQjFyqk3mDgyzC5GWYN3WpzQC8vTLBM8gS8LABZ03W0eOTIhycPLZH9A876VRVA3Dv
yiQmmrYlfqaZ0hfNYHNA73mw4qSygIIKvMrQCePHewZGo884/dNtaNQ7AUSjnOoQeZLo2shZvJSz
Z/YIlKyja9T1Bk/rPJtWI3U/R1C/F3ozDM9Sg9aYhgyhP/IuADTj5S/xRtpGu9qSryFxs2Q25mqt
GmWv4tZw1jcYMONIsR/1qtwD9TSN3mW1sbKWwY3y0XmElZ5X4fys0ZPmWx+XeyAxcXNayHDaihGL
sooaWVrNRaGUTeaMjRbHBT1L7E14U5jositKMud+nOD1b5tGzAMaX2A3DwD2DD9tITi5bhg52btF
09VZZFKLvLXe+bNtIoWVzPZwk/7VCV6mcYT35OJ459RjaKU0Ah/U9NUJiKVI2OMVSnrxsRvA9nyC
QU0LZ3FLPmQYdMsR1yIjRdzvmewP/2BhyYln8IPZzAF2OqsitIOp6j7vEIFJuk6moXvSogcgrkVN
vaCuLhcgBU8pW9zeNS/ie9X1NBvhOZFHXaTtaWrhCIQbuIVy7YdnNXsSWWJujF8YYDBpbsWpjTHv
Q3w/STXKiBxV6aIZBVYlvlN9o/VV05g3kPe3K8b2b7KfkhzfqFPJLjEG1fwB0iZ1b5RLq/vEbc2F
A+W5TEy+V5gU+T7beYC6sOY7goO5/i04v7Ju1dSjBdgfKZcCcYKsB3JDFFje5yEjUEPdWHjk06io
UOJeHSH6UpZIJ9J6ZRgmKNKmFtuJlh7RQ0Szd2yjTC3goujkCjyOXI1PsCi5jBxAxbYnN53TtJ4Q
XDqKt9ujCx6do4vZqZAfSzpXleavdz6fAo/h349r/IIw8lmZI9vGsEqHrJpPNJjFY2lk+JtREkwE
GgpMx1aXtCbHqNHFQVRUihD8tWWdgPb0bhtKiDtHxnI6Ndvnd38uhH8QMWaYbnrfZpYuIFc7RmXf
EYHYVQlMuJ99wWzmrJQZlcCly28H4vXWtSvfUyFnS25pwzGYT+jIAxbYABSQEyeEI+pMk8cmTWBT
pQMSufJGI/Vq2DrzGM4d2Z8mRpeYvek1KTHeR1fV9ZquGePYGeUt7VPbbC4A3Qi3UY7iKJKGVx1d
G/YBFcC7O7c2xPTbjaSenaJiuOmwioX5m20eMMY7J2FroCwqIeuEUBUwFzJ/qeRCoW2rkh5Eu+aC
AT1f77f0sXhKg1zjl2QmY1JGHieOzfAVQbq7kjpe1UsQsJ3m45BlFpU4X1kK0r/cvfFkqHViauWE
mspS7xguqE4R0ZjU4200YxKptjRFRD6egoyLmAJG15uWsiNTq8IwZPaPKLcIxiLvPF/NiyHTm4+C
SVjLvit2fwwxBk8DXfk2kEeaGcXpXpAxFPo6uNMr/8TX/Zf58Or7tE8RSSIAiTVyYUatRBK06eDn
+9NSY7B0jm3VifNyk9QFWFFuiJEKFI53bKYVYB3NM3Kvc3SMWC8gHLD1WK0ZnFeo0K+6mS25t9Q6
+2csgd5zZp2TRyTPm6GzChRSXRQfRyh60e+HuejzhfOw7DUQWY5/8Z3f/6ScgAAXFfeOxIoQgMPZ
52oXRthdIuziCBItY6obzZOfRPZJG2XoKA7pxeXY+8uyvB04AmuJFYuB0fXWiBG0FRwwzTMf4L+r
HEZbshVQkeEP/CwPV4h8K97EpZYYFwJVDgXzP4NkxmK/NkkAynkBNJH8xjbAL6Zq11UVyj3u0tYx
8kLrtOd5O1TLjsNitLBRoDlfj9yLDJ41ideO4T9FzIvcv/pJrLpHF36KqCtapSQecG/OYtQ7DYJh
lR+gVnBfgwbyQnUutPCoHZi3MJ4sgohve0hQlzpTGPETxuQsRJHiOBE0FL0Ko9LP3pBuTaoep3VI
z0s9q6PJV/l4wP0KdTQeLdzpDXGw9QV5LC0d/onXVpfaNKu2kK6885JGCukbBhhqUY58X3RTDWal
+PYLLTppMfSct+Ji+nWXDeNdza15sOjw8FLxa484Z6aL8AVyEhS2eco0dxs+7P8yksCb5H7+QhPI
WnujAXp6DjRGRV566xitX/pYyq443e+2Uzv/r/Y5aYgyWWCb8hZMpmPN3G33hRo3DAnYwczspAU6
bWKp9jYU29KIaeJTRXRdil3Q0eCUvjFYghDLvcLKMKeaMuQQXzeOxgfavYIHsjl624k933ZPbluB
mKMrj8bEGb8++t4p36Wz5XULT28+8I0YHbykDkJUUoJSSDQ7vPCiJdaQ7xi6qv4KL0DYk1U1lwNQ
8nrZ+ISz4kNxLdOabe3iE11ecq2wkC5CZbsof4MoMwQQbpuTWUKIiF3/N401oKpWibUyimLfFo+x
B1mZk8z7D77qVwOrgljDAFsXR4SSuHBSKLew6qaGgSUlU6HXojCZc9fu6Xy+gmRg+sWNMxe5jsWX
QWqRIodl7xy31AtBzx+B70j/ALv/C3ZnkWh6KNo9KINu9hOrdLeLuVvEk2bRhuG+7ybug4eaIf+l
A//SkFKePsdurhsBHqGywVCIq0YSX/zFjVEN7lvPx9KgVd6i7VT8PIL7TVxcKFAgk9qWjI3Bewh7
gh+Snou1WwkELmq+AVXWRJNfBdDHi09Y0HhRTErswdMiamHVPm+sgXtqXk0WmEKROH7fVjT2zTTo
1irKP6DCFMPXGjt5H+6u5ohmoYVCoU/cr5R+chmJaS7qY12DGSCMKSFKw04W8fOUWQ1fnZqgTuFc
E1ZoqVy/Q5z7eq4GLrBEgrWv+vJnppEgr5gXRnBt2KQXA1BT8Thz0OWjNC88LBZ8vS1jRoM5qxuz
iP0D5O93VX0FCCvAsEuoCqKu7G5XlfgbAU3Joz4n3kxYVGIVbqglyY0ALWQ5IdDsS75zpo62T+U4
gFIHTk187SjLUwAAUcBmiZI0AR/9GR6Dd/u4JaYUCH3CHwxtVIDM73M4YAM85tXrEDVujpTCZwut
JL8NzDIJ1W7cMz+/qsjEY7BnAxLBMRack0Z9ZXZMc5URlrig+Fs4s6+Dqbr05PJfdWxhzgUodWyu
X8BvT/YiZQtFkHH7ZT0Iq1o5F3RS1jZKNJrRA+jQlv+UvIlBfu0/paAZXf4HqzXHfxmeIW0yvRu9
BvyePbWQcAf1OtqMM5QlQhy1so/NSrJwlgkVp5qYn2fki9qcQCM1I1uEZOJmVD1jPpAhtqJVJ3dt
sayzA/E3Y96MSrEKb8+YOG1aHBeuiLbyquMZTDQhdVxsSzFX8Qh6OPxt1DWOfi4Ezo+uQCUrbx2m
Bmn+ISUHwL6U3vvBlWgIQ2kvvghsx8hSjXuGke4TNSRPpihEPQLBL9v/wOi6EO5fhf04GG9w7zlz
SGoHcJDrip3lhQ9hDB6OXDkNyTkkglfk5HHDMcfleI7cT0zwS07maP8uoMsOshVLR3bNxK0JduQR
me/4xdGhDv6lLyCumoGSs8aSh4V7BmfgjDlMdQyq1fdtxsSDdcX3VvavInmUEinFS4HNmxzxKvkW
aVdh27f3nbFGbr153Auc60GVOncUGtcVZACgQRYZR0AHgJiIw5yP+C9SEkjBY6kODdfpsgBPOU0e
tctQq5QA1JtmH1dNLq/taC/dXHy3EZvGVR0FH18Uqn14Y4Mi7qx/SKS7+UghtJd+XRAi+g3Cduk7
TNA3sT9Ob2MRnfPsRyLuYcJdGMUD4y1huIEUZt/jvMMahYevoPXC/w0Sbi6hkhMyav2ZGo+JfRp0
uFWsIp5XQtD4w2Rx5zJuDcLvUivEg3qNftEScx76I5vSLC4nxW/+avDOdm/k6iMSIN3XhAS9kd1w
9BaB+QeyWZmxAtiovEOg6/s9L+cfxpLhBRLXUUQQ5yq7oH7MaO53lOkH1fbAygk04j6FL8NwBLcO
R+7iBbR8gl6g6Xk5lBF33PnVOnU/wOl164NhOpbncfMITeqIXzdV2N/b0SRhegj6ZCzxgWLBPsQd
sSExcX8UXL6BSrj4MmlMugL/lrS6NhFmTuoSoN82AgDIPlDKcfOPfjmYoAfCIltr/urQ996f1ybx
aoi4r/hOQ51rLR+X91xjlK1KWgKU3R59qmAG2S74Ce0ClgEuF9zV/XYLgW5Z3wV0lGbYZD7OOO8C
N4VHJfNIejKG/JCQeIPcnwJZ5eiHVXsLLcL3dKibYpWEKpAqqdjLntaeUrZklYg7xRI0IzSXeit8
zsh1qPtW9DTx3aoAnLt6mmZMw83bGkaw+1ophz31vrPGuFkB10ccc16fFYNXH1bXNPL0YC8cClHI
268rvXXYWWAPkFVJCYwUrZQyaeOtUF5ayPGU4djB+jdDdnH3QO9f4fFm6EOd3JcD6tc1ATk2ICmZ
p1y5lsbxSwmIW7noFrQE3Eo/Q2E0ovc+udx0dNegu1C52RMb6DceUSP2ay1uURvxkDyZbHTRyxAE
WknN66BuA/+UQy0kVCbGPamZKrQ+rS/DfY1YBO/AjZPYiadOUyKuTzf79zgkIneYT+AzrtVXgmHH
WwJCg57OHwBckqDAe5nhCj/BgRCOHUcM2V1GG08WYPwOfZgs01LfaXpsjjtnVrDwz3F543iS60zw
WU+d6fJ5t58rkFwaTslCkTxJ2GnUtZheTpBsGHQZSgPh5tUSWR21ESOnqmH+B+OnbARM9rAhIE4j
RAgkXRBFUohzl0P8V3UrxnWbLB954cWNHqB9oGB+/08/4n0UIzOE3TMowJfclJQc9dHi3dW1j2V3
EEj1ti3/A5CgeTj0PZ0Ne1L/yCPfnmvQqz5oj3KiILWTnR5rxLU3oxCN/zpTxZp2Ic0Kz/aMcaDN
/azYjPu9CiDXhceDayLXX7tnKZIj5TN/sNP3w0qBxQSL9rBIW10gYTJwM/5eNeRvpC0PWKXkiDh4
pmMPgc690VlMiZKGqRRz6fnZx7CZc6EEfCbziDCZhu4W4cUcpGJ7Qo54U0ghcMxKIlJFQ40XcYUq
I6FzX9MlSyc6IRA20PrUf2HQpGRyVlC8U6sxxXGwxKTuCKhHPxbTY+cONYHlvKPF8RZym7vFHzrm
8/imGpLv986P3X9hb+ilWLrrHhYm8Z1I+TE7yMt4yIX2tksOjVmvgfS+o8FYJjY+Tx9l2jVcCRxp
Ibd5c06RUTFgD8cQxUx+S9K23Fl/zBde/wOAyjGaCsQ2QagU866qcANn6M+grzuUWi4DWXzoZH9E
NFJIUqwvuDLu45wmggFHwipW229ETOb2AxQNgMyLuNvMbp5LGrozagJcm1eaq35rhllGzCsvD0Tu
tUGPdy4+bM8BY3oY7C2dlPDGnVCt3uz4zVudn2nOCS2uxs8HJYqtaWGunzeHMUNuMwAK7LH8Tv7T
ID8Ji3lyHQABZmqVPiZ51pG5V03WPjO6RmEwT/M0HaCUMudfxnySSkXfFupl7DAWboCo/KJIuAKJ
c2hXeoxyhglzO3dmlTis4FGtvtPcyiCyYwtqCoXcqmh+kQpEjZIFs2v0DPYXF4e35i6FgwzOTyJf
T6B+dF4VssPFr1QNGEOc+arbLClcCw+cv534T4cMN7Vw0GUZRdWJkPgDZye1n7B4fEGPsanLDExm
JN6HVwkAnArcVEmiVcRz7VfjJntZBcM5bXcL4Mp6GG0AUpG3kMfE59lR3V9cy1c4ujTArDGttJOW
lLP7yz4uFVsY+x7OvaieaO0N2h+74haB/yqifwXXY0XYgNT8Ns/CJtJVoQf+15TBs4WfG+m+H+NP
MPOoHomcS2BPELwMmzAXT1d6nOctWOF2FIlyQmqHR5CaDxm5P7I7rKgP8+PeopJHq5cHLjtOsCKv
ftousKbEbl/5ytS28vgoRd/7YXwyD38ZL8mfwXmRHNSWHEm3DPVeQBCwC1MO8uNWn4RgEjqKb1jA
EyWZfY1TNsi/L7bD0ua5pY3DfbHybjqXLArvpr48wyPLwcbn8xl2vGInqOd4n8odqDPET75bxayS
LgXtxWLHzPkwDRcViqJ7pfCdk8NipFY0gfOtHMnp/ytHDYrRACin4fpkhMDQ/ONXwhCOy2mz4f4b
Qr7bvDDy9txhBWICIJLOtiE47iH5AkffW83IbxhdgISbNJHNADGKE4Xic45A//ZzY9Fgl476OBnQ
f1yk/JLmiN+Upsk8mNzxcoDppnuOqrShtBieS8qHvk/thYztwTKazh+llvTKPOUpxxoGWgQQH0dG
wKoqbj4n/NbPHoKi6nEGoAIdJ57+35roLxBQ3abS73HJjXD4tsxPjYEqIPD4L3Lys04DqaH8rFo6
sx16C5Q32L0CdB5rkhNE5kZ97tiNnEcodLTsvg9Ww3qhkRJT2PK5vPXXULaS8AynxJSKBhD5bnOe
/zbZRp350XhUbdA6L+nbWK7jyXu4K9m3rYxFAfyI1B830W855IFEC4kHE8bF2Mq2fVLaZbmbURJl
sMHQMD+/l6jaA++dXIpeBYrmP19hDTkMrZC/KsOS2jrzsSf+bVAMET1rlssroBgT1baWT3hD3whp
3qQfaaccMKdcCzpI+1XlJhInAICrjm3v8EULZ2H9yocBB8yqU5/U8+3E2yBBJEirGdJm2Cz1bfZ7
nBaunGuRrPbbOn2vTU/ET12W/hx7GA07wbZG8q9olMmWzNhm9Z2iRj4OQ5bwQEEthu5ZxGZcYjgX
SxovMMB7mAuKpS6MGwfm32sTIEAnwAvhBOuH6zUtoOSDLwCPdBi6mMQoykI4q8KpXK8SogW78fDd
6tBqYzoFSJYuuxejC2rdedKfIniIrv2HAXX2jswGNboiPGPH/anbMjdzwF1XSaZdOm8xalmLhLTI
QXUtrUJm8V4vHSnmBKyB3gFdutaalWBnEXh8FtC7EIoOsFEXMYx4iN+qEVjnjDFOy5Uio9GY3mi0
lTptH9RKJib4d1I0/aqxFMv2XChKE+k3aSvvkdBbTXYLICoDwMQbIWLhAoLNxLLQhuJRlacl3fPc
u8oXnZAoF13yVujWe1EA1OcnqfbyZjQAPZCbwTYy0Bdyd86AOO7DUgsZnetCxlTlacwVsFasJVLs
dkZK0XhopbQEig0DMc7hdcR/fPHF3WJlF/HA8UiCgdXQdqK4X/j+w9iCxaWlkjOKsaUhbUyB5CS+
rfcv7/aUWy99PvylYRYEJ0rdmzAFv7TEGzzF3Lmf2zaxqiTlfhASk2U6nTzzYIcdAI90VhOFdGr3
J0wVlm5kedED0FkZo1wj/npKSonz3XsrF3QbYLDSEwoEJrqNUtlsaiaq2Ha1hkLSYdlzNor4n7GO
Iwu3QdyoKn6ah+ek7z6Jikq0IWygiocoeJ1YR6FeJ0bcBRzB16OgfwsbXJ+mdl4CsZRYZbkZwKW8
D4/YMGFR6Xj1rMlx61WcKPTdtDFDiIq9eKYaFN7yif3HFdfv2WhWEKgKU2qk7ncmA9gk+eYlH+us
yqNtAbHVJ+LOvX0OwSzl8TFbLo+RA7KHLYSK894Oq7eI9WI3sZ47iTiuQ6Sg+nSxduICZJb6Kepb
zj+B8vJp0o/0ItUuhayFgSsnUX4akBx/h3PfFV9Qy3XITOw9Kigl+NG/S4FAV0zOeS8d12HF1l7s
/HzkRq82EoKmiZGi4IrREsoBdKL9bqM2RHsMHIGoAKMu5cwgIP8xiZhWOC/KRRVcnzhVCglLoCMO
P7SqcLDelS9tpo+iwAHYTEXaTFTH7WB6wZqOyQSe2sSlUmNQIfZP1WVGcg8Nur+oroQgfzF8wlG9
fTF7b6EM/I8dqPH9t6apDkcVe0G/811Ne4JvXTcRLkxrnLBsvI3RmUoFMwLC/TEUTN/Nkyl3XDni
VK3mhgPOrmVVd58GMiSE4OtqQr0GLpm1acdFnQvT6sAyaewOfJd1uPWdu1VltCJivD4JvbY11zBS
MhmHkPwsPsQzoEt6KmUwmGWmWz6tWIt1C87U04CD1sOnlION4EEsMkZnGBwHJGsYAPgXHsv/ejXg
Ubk04iEUbi4E/J5AvFQvgR4gIpSnBBbbLZX5CROhqo2E3jegz2BIajsYHbj/51CNrFLJQHCDXY1N
lW9ZvSIxyjrzvj0dtCw+Yk2nKanfUB6nWl7HfYlzyP/gyQ9n6bSSEQDiGjLjO1WZY4sM6uwYzQmz
7DAcBbHjomyOAZsMp+M/CoTYnW0gN4taonnz7CqHkdVKq2iem5UYqSwTlnzttnHKEb+KyNP2B2R3
qpZ5sWyLWxzJoP4zdZTsOqSFNDLZ484ig3uSPa+4IOGmbchBm3EpNZ5o7KyJg1pokOryWvTXPyms
05UvunhKnGswJmmJtFauAgz/gAPNO29/GkqmVSxP6P0LBZtVJ9FRgJRfJWz5sGgcEqUt8wXtKP77
rIfUjFlhg0NtagIZSQzWr48O0zAWmOfN2LryYWQWFclKZukQuPRzEpiW7MfaZ6+jgtAMmjXiznKo
sHbepF0Mwe419EMJzOWfrY911PMjWQsQVL3EQm055Agbs/5iWdJaHGwqPIWRFxYflrRgKKZLhDE1
+o5vm+uxvDlxYcgkq/jKpxBssp1GK9BDsrQjI9caLR2rJk48MCqIBR7txJ10nQeswykW7nDnS8OU
5jCeOQPxM0mho72VHuPt8iOIHQeWXm4hFLVcWuymCO7iK3zIg7v0RsKpX3Ig9vcgEtKVxz/wk9f0
bIVVffJDEiNxODAY4ZRLxT1j4BC6jCVk31ne619Jd0xQswFia1u77l3V9DjrDveHAXvNh0Y95Tsz
oJCOupfBTxQWm28tIlyiHJS/O/SwP4AkLxtQUpqggw1f3pc6iF+HlIosim7fGKYu76jHk/SxsL3Z
UAmMOC+/x0xv0XEnIOyrVVk6vOCUS67khGDSdCXI5Z/AM/VgcAG/nAL1sbKUNKJk9Q4vjhuGa1aE
ZjXKAg4vmwyoQvSr2z0e+2f29lbzMv0j+Y12wNMpUPVumENq+U8yKIjcNec64Qbt54OpI/jvJs/j
QQPJ1SCRtfDX6Dbf/BHV7e4TylqJFYxyAj8XfK5/vAMVEHgwwB7GKgLFpoTz9fAQSYzvwfDISHib
IB+U4Z+OXZ+e8xm1a0LAqpZ2zIfxDObwxT+/0lGKdWBAOP5XuZTO8jMQdvmd6jKn4HCKdKk0r4kc
6NlR50uXgI58d4Gcj8D/iJF8OehgKvM1QGPMa6puKpGJb9ptWOLqA2joz/F3TZeaYK99pDigvZJY
ZL9AQx4B+Wy2r2/7/EilmJwH2c00VdBg2+1esia/uYNoDDEmnSqFNRl1Ub8qNf/AnhzzMoyrlLKD
7R3nkY/afUu8aPCJR6OA4xNLvTOQK4T8wurDOWRa0DhUYSbC6wIKHPfKT+Tjl8rpg1y9bea7Ic9e
cpj2guad6/JiLQizDbUHOv0cFz5Z8FqYzwPMFeRDIFsie9DUto6ujx/3LeGy1dXvbLdVgrV+4O3p
7wEZuzXe0HLHJS6BatToDMoTCLpy6qCd8eb4jB5dBNXATKvXdTKOFkVMxqL5jNa0i6wTuGpli8zB
MYiA8aY3Tuhbhueh+J5qHA3ZJbTz7BEIqFVN+tLghR5/qXBr5UUf4tpNMFC43r9CrvQJI7+r2mKm
2ulMtcPzcTGERjRRCDIqKyD9NqisNpEWNEPWtWczFr8SJyEBGuqOpuOQ+q75pTpN+O8ABvtTyht2
VdwkffWH6+BGQPqBbPP4r1yf0Rff4wE08+XXjVeRNberoU6ArdJagCHt2fCou4yGipGTvhaIBoCq
ANyQDiRD+2v/XSkhDisDI2/0mSeAYUijtuLD0D3/lCcWS8wn/B+8Ki0qEm1IL8W9BOI/zIXWdipK
aXl8IKC1Gm6mqRkeXc8dhgNx/XVQwZG3gR2mkvaoIq9vsqtEHto/bsRBibbvktPHl4+e1MmxLXNv
uo3WMS2sJTmDjblzBoJXFi75f5rWjIi9m5G08SEZV+SBj8pN79OS/m5Fi/4itF4Iav0PQxjJMJ0h
vdX0BNw3/HzJBEAGAQca1qsD2iKPAPqVCrVsN7K88vAjXkHuvT4SiD+A9i4F33ZGcA/30ycOPX4U
eJ4NVLKHnwbw/BZvH8+xQyh1uh7zt8K62gMm3Fb90FWbneUWpqP9Cse+4nSRnzXJHtxkPKR7X9N7
PGmHk1v+FzvTCoi8v8pSxcS0tsNH9gx8VjaSdNraatRkwWEuw4OxSK9PvZ24cPdrgAsp2SA0Yhkv
cCAEyx8C4bbU1/yzePG7zsPvKry4q33b0qcecvJf3D3PNC9M7TVd+hCC/75Uo0R2g1JxWiXyiudr
68iy9YC7N7mqRxm6v+Ki5TqYwKJSJlq8Ty7F/09Mno7RgMoRF2sRQ4Yn0Wa2DHfYu5Ua98SZWeC9
/c1V6pFL32Iby1ErZKAtyun+q23z3r8Hi2xFpPApsxn7CuWVGFKKTvAZ6SrJLLIGEDrKWcpA1R5D
IGHvCvckrvXZGt9cjT+06nBVBZEuV4O+FsBTwr/0MtFwi78utPewyPogwXS0FbOO5N/xIMOndUf1
5wteuOEsIygQcpPgtwNz49RmcCnNLMpdK6k4zt5NLjJJTIGvrNBOhYwmZ0REWuDb1+lv8dySR/7C
aEqaxkAR8e7crp24HI96cJ+v1FnWHSS0+5Aj0UGX8yaGQfk5ZWFxE9Dah0+WZmzQ4k4/o7JSnMWk
DbpQ7ludy+EEwNL0lYCan/owCxAaatsEDte3ZwYeLasCJRVIIZT/IbwVvqkcn65glEjOdvz3yfUy
KLSJJJL2fRWg4D0uslcBHCWV2K5wkpqjS16S6yyjA/UxvrWOS4VynV9aUIYXZhKtp9Qb53QDaXiY
ETT5nZds/KuDdlOg3OIipG52FDFSOFHRBSbno41OQzD41+rt+8dx8InxBEIcEqDs4JKOTK7S3hZx
F5llGvbR0RMq6XP9OIcrqzsh9Jra8KrpY+Y0dqw432xCT6/akfKZPcSWdwaqSQhBqLQmJ8QJ6UGt
UYFkNjf96UVc3teO/sJaZpp7ShL7wTzETheh+oBeizDSuIMSK6CArqVfzbE0KfDZ/zKAE4C1v4GK
H/RNx9BMHGumWASEgT34QucWM1l3eSeD5t+KDJnw7RiuDd0lxS29e15dQfrFFgKV4P/xLEGGjvNV
O7ytfL+HuXnzJDkyLAJ5oifIXQach7SuRmNLGQ/CbqhZ8flXw2mqYAQ6u4KlFXbTT02nihjOidtT
zhhRc/hAN8HPKwxa54EdHUPuwl19AYvsiDlj7s1zwYhSyZUK/1H3XHfsf3VxSxCbziVaN2zMQTpV
3dgh/rRrxMxghbmr+zd5coz36cCt9lPyU1/sQOuK/FJgg/+fTeq57rDfL2hwrnbtwyxoAVmnrvaK
tUh23c/uaCk79fXFOc7k3l7N7kIguWCko/TDKv/8nKeEuFWXUk6lYNI9Nj06CgK4XndxUZVMgQ4r
B0mPUeqvapFO+jghKwoQMiQ1LuuapW7e45Y5QOIRZ5+94lD0iv8K5UCU+NUUMY9/281HjkqpHesK
Nkgl1SGHJxBby3r6PLMPT43FRW0K3wpCMdDbrcT8OKdrWYYU+4rgbtHUEL4tqXs65VAWtLvMeamO
wCbLQCwkGgf8+uLBXMNsZH/AYBp7sPg9nHlY9MZrO1PmOsE42oB2qZIC0UcGQex7uxtt1fLCUexn
yuTlaL/fPZAsOgghCjmUvhvrs+mWYtb2fIMnv70huLca8QZbb84LH57bHjKLTn+AehzZAESjioBl
irXqyeYlvG50k4HuCtA/GgnCzGjZ0ccJ183cjiRKBgJp2LtW9F05qRB2rvji3rblFdmFzbLNnzv8
AsiN84Yn2oYoZch1OHoaVdE42aytkN/KoniJogM9RnWiKdJOJU6CHq3xL1GViaqjMuTuHRbmBfuS
waA9My6XCdWUEHvBYPvTn1qRILWfsD0cyPDMJfOyOu2WqI7p9kJ4q4xE2e0s35Wuky1kLKoOK1Yf
aYtswd4PUQ6tlT6LHUvUQW7pm+Beu0/V6z0d/jQHMe4VsSCbEM/phJtRgpbg+cRImCkOG/NMlxZg
Y8t2eNMLXEP1n2jJl2ku6l+gB9v/SEBu/Cm1z4GoGOmCqoq59NjhaYuzJRqI887gO4YIQbr5AZWX
RYp3RfShFRP/V/R/qy3VQbbSHpUfZ2iaSv0soA2NVZrMphIZC9S3vmiHIA/OUk3hh7OePwFyiKdf
b3aJoyojkZpGo7CIgoP7WcUWL4H6br8n6x2fxkVoCNSdLeDubCe1hnnBlsJgyDZwlt8e63IEupL4
62/LekRUZ/A99tkwQhac3/Vm5Wu2PgTi5mFn9dSUDV2re75rE2pf4oMpqGJ8Xh2HOyMHC7grc5OH
YHoSk3uiwIja5IJtrprBWicZ1Kd100JhqaWRWzG5c/NwRbZzgMZdoCT+bWVBpziYcM3B1kSz6IHi
uA8UDVrd5xfd3IBEgnTAWKvq/mnlNG2XdouVYoO7ZZkEmd+25zmWBWV1YgeNElNNPlA6LbidWhej
SkxQKCGrA2+OddJZV0uCJzARaCKqZ9hdM92TmTTMyh/F+woX6VUfJ9JDhc5Xn8UC7TN0mum1wSXx
bnPfY6GjBPQYgUftO+BgiY+j4GUoWtgs55R2hrhB+R7xRDH7Aah9EWkLG1uk5zsxgGi9l6E3b1fN
PdOBTc1YknMXt6nMYwO4QV/tKAAhsdaXmByLustsElrdp+6mgHkMORhlqbDdgSaHq4BKc7JQ5zT9
g0XNovaBLP914qWCszGRObW47ZE5wOIBTSpN4U/Z15JwPNwSvtELztnX/gOjhmNowJGmT5yMdyjZ
E2rZlcPAwZ+3FU6Y5HjGmFTVnGFNA7mk9UwDakpNzbQtB1Fm7QOp+5m+JKVinx0sx7hB+S/MYN/a
Qmxfc5IBmqY0B6yfbODwaQeyGCRvJS16B2/TOvVDYgqC9dmFcK91PTNjlmxb/5wAwHx2E+ZLvj6M
ZOG+kvCEnNIXJ8DWBjRhng7CsH41DHF8v1pPohpRtEqi5QvCBt/5GiWC1o8+jwMKhqKK1fGVkSJ3
eUuB4YX9S08XtlP+7jZH/LurOdE901anw7updoc5qXBalKuml4DDcSGk5JqxjvdKuKOQ9vUeXH7E
tjXuUxU3XkZF55O4QeS6Go/eW0LsJ6dMhAQJpm6UOXSbmsqeeqScMOJxe/A39X/mteY0e5CV5wC8
+YIIPfsmaxuPJ+R1gj69mv4YHm3HMnhmUqD/kAC8rbjGidoBXGLmeeHs12fwDE/O8lnvvePMfbpN
XC2mHrJkADfjkt2MJXRJd1QiKjLcL0ocMZM6ceh3xeNdVfgwL0zFoAWpSDIA/fDOS6a4h6O+7mdN
cgDVr0oZa8YOLkYGzNQ2FRCSwpfkVhVKIaElmbDnjK1GNb9niwmMLklAVlMDn/otqYkjXM+qVTFh
mm9HU1GrZnsd5zROF/Zq5vVFafCeMWoBgnl8+89drfqdQOTKSFYNnGBawA/x02W2wbDKjS/h51jI
Sj1DxyCAUj0Ix8G9JbU4uBXd4j9TW/bmBtmucIi81aCEbpmG4lArZU+KqBZ3oodxbUR13XIvObJf
krRI6sP6ODQcUgWLsIwWu66vRDh34KBZ++B9syGGZPr+hLLnOfVu674WXf+E06uCqC4St01a2dXP
CktmzUYdRc1P7pnj0ZhK6SeKLHZA2qE25DxvF1yQ5RdPGu1Dg8TSYXU+vtQSuq115Cr1vWJdfoz7
Vec9ITMxldtd6dy6r8JEIrILeSExIDGEWfQVPEjsJVtFOvOPB6KwrsriQAdoPRtMVedxYNftI0S4
8LmZsLJKPCx25WfoiraQ0cXqCCJuya3T5E2a8EYVWipP8AsuyyIXGACWwfqSk/K2p/0eqUTq+QhW
68gaBV0mnyfIO5LpigYlKiXPe1V7CLB0TJ4+cTCepZFBrn68y6NoMEliYqPByF/Z/Fv/UDjFL1lu
ykSCqWRevMfjMJ6NwJdyiD/5UKBNndLayMy/lsDLr4H2HZ7X1SFb5NsvH03E5PB1Z8K63h2szqn6
98Qr15O+EHl9BSBtOWCKvy9ZAVZ6oThPWjgv3j3POtnShZcqEB3KhJpCQLGvtdb2oVQEStuGDBoN
M4B7dbGqStOPzCuRAbaPOSwLIkXm5kZHsyFQPXcSMvfmDHAeOUW9/4CYA0P0Z2QiQo2OhRvzYTjN
p09kLwj0iKW5D9YcAn5DBJue0PKgaBVZtcAHGMkHiw490U9b+u7/DMzQ3z28IKqbMnpRWyr+hoYd
RaHDlVMB60r9OjE3yqqun1p04nyAwZKJrtiJfO5bp+nXZQWLhT9cVEgcDLiCBoPaSGO1mg3He7bp
BLfkgyliVAIc7fVvNKwAFSZ8ejz13s1623P4KhNJTQ2uYOYCrX0HQNkBKzq2BoF6ErZ4oGp9KA2c
+aqLN7Gl3bX3Nki/BUd5wGMyPyNJ+x1L+PqDiqPg5Xm21IcObgJc1ZRGJowp49W0CwBd+zfvAtXJ
k4uvtdoME/u5zBU26lMQIo3i59+k8kKIP9mo3pjKK4wSYdP/Es1XmNjQaXBU0k63tVktCQ0Ncpev
JoSFcwb+Uc8LXP9xNmdMSnF3LmxiYTIueaIvwFJGbikjwF6+B3+GepyiCGGraPicnPMyZvgR1UbN
cQJmvDCS0Cm8ytVgyGp1A+U6qyawDlQGSYCbdP8gpDgsD8as+DZ4Jaw5LayMgyojrYNlyA+ohSjR
MsTmq2mvzRD52fw6dgwVb9K+lWwHr6hwqYTitpyo9HY27bwWkmKs3HKa0BMLTdfEPjn3/jg5OzKr
7j/w3pt/KBSeLVpChiG26YB7EfJx1x1yhwmPX+gK9bsywUjSHp7RxjBJg/x2zcEP0YHHyXaEOgGL
FKoWwArpfwNefTU0vqgmMPtbYl5R5yLMyUjPs6P5s9IH6kLanWAvZgZjMPSvZTq5THUOr98nYW/5
Pb9CK/UPQrgN6fR/uAWE+r/a77P0mPkWmltnm59WAbyeIiZ/uMG9Mcf/hNCEiClZ5VKrgroAg+//
vG2x5yDDWm45o2xpc/jpLJBEb0BLbh6pILF+wCHRNQrxys5V+MNMKdeRlCVufZcyOH9cSSMGKwV+
WLAzpvG06hmNVeWFtZS+/8gFle6hjAsogjwSG0cdbLVwpIV8cFscaSsEDR1F2gQuuD6z7iBancTL
6pkXRz6OlD7xrm+dh351FD5nwRuId3cIlkYxbs7AW0nLbNBEaYLjjHKXkPKP5MflPv5ibu8IKbvW
NJ5h7p3O6t3B/vUXL1mpvFyC6nlqSbWrl63296cs/O84IBpDATszsHTzxEOKlHWmhGCpw8NVRdoY
+7G+o1TkDXPFHJGuXOStg8iDlJwlgB9JWGfwmCpPJ5rn7pUfaWD2CXTzkJRQTLALRgxgIpnjuKcc
b7/X7J1lnSeJrVhGpnd9cSwD7RLICqO5QcEtfQbvCvZ9iKRPihNB1XjZs45JyIUWpimDJdog14JC
rkIMWqJgebstE5YzgknNyl4Z1qgDK91xXWi9VH7tboDs74CVtpcLxe82BJgvMctqUodhUdiJbVvZ
fQa40Z/JbT7GFJfAU9AidmLemdNPuTaK98LCXx/NeVQ/qdcPkNAp+aUy6MnR0qDs5TFNmlqc7Mej
pylV6lEFSuQGuVDUOdJ/fF/Wd2YRNOnPFtYpJVzPwjz1eni5sacd5+Yzjm3gn676bLMwBUbUVtfg
uJaigpXF/nh3R6J00KNyVWIdVlv4Q2cZ/PIhOrrOIpS97iFWZKJirp5vFQheoozYDFDIb1XWV5NH
zXTDTaoE6ZsUjWMK8C1SAzLZZj60RFQRhUv2+LEeiuzsiLgdcQxUqOk+zH4ZXBLUZ7xuFSuTrEtg
CbDADhPxJ9zOso2HqFa750t5RF/LtNvlKOZdoY08oDtUsUyEiL0e85RdjsQ3ZdmxJoEFBDioxNY1
fUttHhrUN3E/1dPnhW66slqWPA+XiKAMKlwYwaTdVKg7WofReQ1Y+aPMX4E6OWPRF5k6mFe+SejA
t5IH52sW0TD7FP0JqsnRegmleQhTqhYxnnkk6AQbWag0jubZpQQ/FU4rGQa6yCNx4PLLIF+lQ24j
l/p4uP4FDfgzfBdPmso34GLIayk88fhyh1/cfUU4qzhCVTrhadACsLpx5lS51RNJaTZd8f80MQSY
kr7t2kkLZSEoRAj3Y57qnjQzeDMBbv7JytmuCquBZ/oDc2FFsZhtm+F0qq9vweihCq0yCkte17yH
W+cmE+fnHoCs6gl76APzVH/J96zD2mysL/SAgFZYaZ+9XejjXvYQSk3ZRxJ+BUUH5ii9FFMfwc2H
pIzNrFtxZj7o9vxELOB9SvXRn6jt/IZkffgo3cPkVw8tdIJoK+GfEYbUcwSFAkF3gX3EqWDzHYeL
DD3oh6YVh7ZErkU6Lyw47jypkE1bmfMxDDN+IihO4grT+3Z0fMgAU+T3j/VTr6IRjOY5j36sQ2rv
rA322c2tAc9LpaRvsZRoz0QSqAyTYDYRq5+j4n1zQwM4Mrj2WjHi//ioY9Fk2iY/mqllRQdNRCd5
IMEscxONW4ueSbF+VTwDk1M7PR74n598rFtBH/6h2i5/lUP86tXpasCVuZLyQkCaj2CE5z/43JnZ
TqzTJU4LLRd1BcuZpBe7VTi3qsnUgFQyF29plM/xkSYnj78eaU1OTx2lHDewq92VGGoKgbh/2Ghy
w6FAd8HnhjQvQbPhsNQM5mDle0AQAF5RNJ0KiFwOpksrkuDO/vW168lzXbQiBYCMkHBZRfQWHQm5
a6H70hAtHtmc8jxHPLn4iPHwF85zhfFkGOzxZaf0fRaSctrPAj9JBta+FBdabmZDEk+L5tgs20ao
IL1Lzt/u7/mRzAQFjHTvEH/yOzSfl5JurLSRjwsYEkZxP2s7g0/o+ME1ssrQ5P/l82u6qtxli2zj
WAhFer/mxJkVQo2kj7peNTvshgBc5I5ibxlAqoafnYm6K++fnvpY1HEANwK26vi4nBjssvo160+R
PL+hT7EiSmn+ib0MQQ+oAPHxZ7cYbSrf7FyX/bgJQ4KTDkmgeLjqdOjBGQDLJzw+YH3fj+4zBFgs
kk1isxfen5dvP3HM5cFXxd9O0876GRhlZuMglFxvd80znWFNoeEnP1QFX+Y2oD+FNBlFfRNQX4vb
PA4Dz6euDGgx4Mft4MEk1aOo80isCAzxbatensV0elKny5j3JKH0FojePRoxNUPyq3gs0VT6TzC3
fta5L0KOZHKt6sYvTz8QXFSmfWTi29qX01u/kitw3iUUK8F9yg4UmDkfg699rQm6wnM4nq1UVin9
rGOi3xXiQ+3qNQoVjN98uIlExRH8W6IWB8G99069md/t1cEjGwpmq22j5lk79x4IiXTNR8XOrUDJ
uvu7UXNA3nw5gy28N4PoeEZNcGl/pNpr16I78J4MSJn1i46M0TUBPklibkU7L6pz3R03RPaQLWAY
wi4D2KFrKGD1h74vkHtLn2oZ39/Rz+GY7lijDNmKON15VVi0DUOAeTJdMQh9+dpSLfcgOxCvrf2X
XoXF04GH/yMDqPg5E4prW+zZrATxiQi4NSsH05YPYg3n0LJMIAPDrRG+vvlHcfAa24wsqKxMerDt
HsO61a3NGV1JZM9AsiViWFlIr2nfv8Sdpw9GOFjzk3W4fk2zUpm/KhdNPDmSecyAbk70AJPxrt0A
ahNA4vs9IJ+RSTvXXHZiFuCh/IaDpMGVHmvzWlEivduvI1CEDPV7w6MwAGhTaFfN1p4YTeK997+k
jo/ebT5PTLz2TWMn0lG+BnAgSX+vUXVG27BX4w+3lMopZnV9ZMM37PFTGXlAk2HTsVtqjbCLMBoA
HUiAh/1sIq4deCq8uygrNrsqQ7xnmyITPcAhkrGccdGLimy6Q8LymkCz6xqMKcjDiS82BSXv5DIz
psP21zZNtxhZwEYlgyyZZ0xIO7fZIgnfdj9HQIxVXD8a1UMQXj/z7VrPq3LOuZFhD7qsmsYgC50g
cucFcw7vuy3Q7yvrHjLAnZWEzMafAPaSe5LvrolarTK5LxgVxUPYWQX16sibGFZlnaZz6NbTJV7Y
lsFeFh6ifyKOYOqIyiat4BUUeIHA1P749NiBzd9M96CMx7QSx8Mwq+7OF0OYhk9dlCUi9zptK1ze
/G7hdyK0BqW2mTpTOMpz80QLTCA9B3z6pVSjjtnHAA4OCTqxymPTp/wpNkGyv5D+/qPiSNAAICBj
JMbeuP2bzKvNRNeBlLwjGGx6U5lPTFj64SJyE91qGEcnv9me6UDtBzqXmQjexxm7NCRFbOSte5zA
+kmztpVf5711nOjM0g1W6Oay1BYnKAkx+jceqpV9ZNrX31MEKBx5HbsskdM1xsnIB09CaQx3+dx+
ebZth3zMS6nYhUhJTknKDvM2NzQW+uGpSExnHdPLhbkxCLc2zSKZNCLlv82c7t3cwhcBjRPBHLNw
7QvXf1tbTFsmmfTtwAsziwAOubSrisGfkAg40cYo0IY9z6NeGloEXp07nBFRM9LJXYaiKFDhbVLa
0PwCBqh0Li4P4uJf//AGx+JhIzlc7zwJB7O7N+3AmA7h9+W6ZWjHDEzTElaOBBvQhwHJPSZA8EkE
4aBjpSJayr496qp5OsYH3PvWyP4EtdGUiBIBkyCiF6jK30zidIKCGvOlQPy5IR+QxfiRF0z0XjhQ
+GiykE/zErvQgbQuetU1lOEQVJpAy1E4y+rMxeBJjP3fHjrXSibjUJ9l7a7gAL+UwttJXL+U1XSP
cPiUfwUBQw7gAERijddLwJGqiJfoZlyQWWvOm9ytMmbU+rQSIIYaZyNwfN7+b/bbGYeCNNuE27Vr
jSy0wq/GwljDpcqenkM5ERxNf3HYeIAl6/CWf4VJGjicHprSlcULWKc8zfjg5GZQchKKW+JxfIXQ
T6X7bRkNY9o2sZ4xAzFGGculG+4j6rZJkKYiQm7CmHrKSbkJbdi0QBPKABlM55hMkHev06vq3w7t
4inJNOLhlBIJNRcr9MlS3BXgM+k3OYkvgzDNvMx4EAPMN5vBq1WZDIPyJ6Hn8KB6zW0DD8WQyyJ6
FEyPyo7ZnD4hTjJVXkpmLSBC1TlqTdiv7a+/TI9T/MOx6BbI4PSfWF+nMjlqkAxB/II/4D5riauP
sL7F+9SYiASBSuSPHJIaM66WAeq50H0CigZU1H1X/uc63uLomvz+1xORiQyHX66v9i8P/wswiroq
8+2KxBglTSeEJOIiuzKVKT+QL3t/vhd5OhMdpTGI2O3X0pby1OKM8HaElcvnmP0dBk45CSxYQbEm
JJG5TK1846L1rIgi7aVVXcTvIQld8PTA6kDARRUPl32skr10p2VrNtRbuLtcHL5fpI9PbRJRQZOE
sCrkbC8ozuSdGGQgOYFygcedgNkrMVkTLsdlRQFGYXPX9S8ZnSThAIUU3Q5eoB3Dxmqq1/TQogu4
tFNSMym5z2mGqjntZH5nXE5hprNJttPDyC8zixi9y9Pmva4r7ujfDoPoZj+HWOxYWbGhBr/kA1Uu
wOssZL0uJHb/DgECPRC/1jxqm9Ko6IiSUDHqqAYdsesS8nXSnAxovDMCDpm2nbZc+wVUBlpb3Rlt
BxonC49BX0UjE7nl3830ylkgAOUvp6lHJm3zLj+308PHoqB2CzuKaVxA0C2IwpeolyU6YT9vJel2
bXTseWMCAvGFaUgycKiCzk6spcQiNJbrjtgEznZcW3lXDyRldn9YlNt13o73Z/9Nv6AQuSH9wQG2
8cL1K0g0W8bf0w2PiL5NtvajqajSzGCNF5qqKGsv1TnUhBcLESYkZeN+bFH9RHmm2c8f2AqevisZ
Mio+I6bBZR/+Sx8xiVx3Ok21x3C/LYcSQWjCHlzzfLtIAQzCRv1LtpV9qHrsuvkq8KsVJsNKOSSD
U8SYrvusDAXDReUal/URrJtQYCUIRKZO8EXF1wAW6i4ux7x7GAjWhXNTPI98sYo7TUt4qGzImRAe
Lo1fmdzarXAHdB7dlCCzCRmDImMduODdesWiCRhwbfMZT9bEnIhJvFb5eFM6jRH5+mJMXB+krKTn
ohY6NFbeVxf5bqadQWflufZmCy71hv6LujcuFznYb9v5FCoyhSP1eAb6/HDVbXS0olbiDgqGGcJY
aKyGEFlHD0FibtkGzlI41eaHSfXd/mTYSigMA4WCZGZ12DkJD7OvQsXNWy6aMugdvD+hm4a0fEyx
caqeApjKE5DBitgPeorrOsSqSxcw9PJbldDGHCT4JJHCpKpmjWZkWSLpTy9U9NlJMxko9zULXJqz
3XH406DWsSksvyrR7Q+gtPOH5G5ceV9oR3iiQ3Ls3pM2Smr+lk+fSxJftDahcZ56wghL1FYL0kw7
j+/ub25A2UC5+AzvpzKpEPvQPebCauUUn2bX1JwAOoxJ682LVDsSLU8mL23eWo6fEi6cH+MqC83S
Q/Bf9tFEbJRfV9gGmiWUr2wgfdtU/CIMwESGllNjxUJvEtwavmGxRrLHI83wSHHGTf3rLRLk4tIz
ZWT2cnHtPAGgKgbQWZiecWx2/EAQUC43vylmYcCH0W+xeSBcrRZHXJqFVPmhVLjGl0AvnZhDCdor
P/ullR58tu8UpNOjxnGLFg6gXPVrbRhbsCJUagRjGnNYasIF98R+gjJkFUlm4Ixl/3s8eog/151l
/ak69dCOfc346mQhpyN82t62Vpzk3h0KteIQYz+ZQxi2Fb8/c3RjXEi/diRsJ25hdNYdSTtKn8gW
A9IoQbQX50UCo9g3Iuojn5leDVJCNXFJ8dbC722cs6ShCe58rExh5Dj5wUvtAm9prwnJt6YmAfT9
+aAIR0AjA+jWJbKpGH7z5s8CNNMLJriyGcIR75j9p3ZAG38NHlCHg/7qhxjwbkUq0SKp0fANm2m4
eDIDh96905O0Ok5nqbJ61Pa5yflBX0YhYsfFuYGFsOYcVXCAPB+47i6C4+y8jjl0xyk41643jDQB
j3GGzmP6dUy5r8wPMJJIyi9E/4dOLKpY7IuPmQ3mw+CfjmBZWu4RZ4MNmevDO8AiTjvbpOR3JM7H
k71rERe7NIZBja6ie2fGCFlXhHY8rzUI3ieLbAlKe0diIq+HVi9tnMsJ385Kmxt8m/qP+OtssRjr
H++IahN6IqjB7DgAuiiLvYyf4udJ94xFyBgr9Yn2HpogDNp3CIJ81ztp+GAkPOcTqg6Bt4DTWNi0
fvYDLrhkv6kn8O2VSAQelPEo/M62ylhqn6ihbxkBRyzo7Ed00iGbLdOJBx+hFvZlp/v+w54Z/G/T
hn5O/Vv2QpYBI6qOEbzIcbt7pNCxlZ9XtoHrvmxVLes4/Q1QVXuZSZxjmC6hKd6hswH5v/Mld4Eh
gUltdwHkSNm6oLIjCFYtv4kTMs9+Pe3T6tiHvq1lrvRJ5G8Eo3JmoT8PLAHsQu2H/BmqZa70+/Zz
NtG5U9n3aomVWJ2LhM8PVXhVTZf6GMAoPInHOSOkiuQuDedsGzqj1L05WzScw9fvc+nIphfg9wfm
V1JnzdA+gXvYZMYxO5TmwQoFH7w4gYjcFuw73oXWyJzGO+2uDUad8eyrWOkWQsTqgA6coyWeOYX6
ffcns5CTu1DbGcXbXiUWYM43WNmENZ/esJeG75czj3Ji0Tr5FS/vqXYPn9RUI1qWhsoaqLmn7QSU
1ZVxpPsRLEaT5tZojM88UfZupsbWMvpT0+3W7UgFAlzx3jiIVfsZEaGuSWA7Ck1SyjM4AgTqOYXd
U0m53CLb94iEz2stkPaW0SnBLkyh+LDegrVOH6jZZQEJ3LA+cD+QcT+z8b4A6PPUo21sVrz7/gj/
6paRsjTZvFO1L1kE0Cxzp32oYsDji82F9r3ZM+vLvc0NkQ4KWUF5zdiyyODK3txwSS3/QeEGXVz+
BbmA5GfF1vgcNkt4uY7i8ptZY/+ZZdAFgrinllDt8di51fNC5/fZZhS8a1lR6dDFA0Y8tDG7XGB/
IywCSZUI/Tjn6/T556MfF06R1ajNzUIbPaKjxSEEGlT6UuvfxlyXZk022epjGh52tn1V1UzhnGZT
L4+cefDd0v4YYvydpkpMa4TV2EHA4ga3mx/8AzUp6YEOtpDSkwwoN/Iy1+P6/drDR/ZgZpWtfI4F
iGyaz8UK/aTwSH1Swh3OIbaGRWzDPqEGZ/yuaexokMfcW444hbtQdqBKiOoQir1H4AnNre9Y6KB0
8nxJBDkkwGII1+AHr/ut5PH7D/XyDjgzZ3EsVPt7PQmC5eiiQde9ZltzHzNcorVJvsoWGK5ckH+a
TK3homjTDy27yiFGKYp39L+ku3k/BJ2Q1nOMLaqf5c0WlGijz9hBCA2fJvrcFcsXZFpcOV+k3wER
EWiBm+CJsmHOE29VOHgwzbT2OM1NpjSzfX8zSqPzyWoeD1uOJh2YqBnQYTj2b3x+o+PC6QT4/nTj
Yp65Iz5nQRUO2jPbDrWSpoV1W43JB/wFV0UhxrwN+VB2kfKzqSJDhJzej7LlwuD5eThdH9yAHMFs
q2kcgw0syi6LIXTWaaRtjxISbFePdw1ell080FdF9veg3ysGxEeA1rgIJsYzG3HzZ3p23gHdSGRD
aNB/I96OWrKgXJ2PNkpXc3hQ+uZR8iCMYCs4Mv9mt+IhADV7FoL2gztI8RSKMtjqy4tOLhGItXE4
p6pht61hGGwOSojQyxzkGx0i5OSm1iQvPGcl1IF9Y5cqvkTbtDbWhHmpJ+wNqCoxAUdCGq26Fwpt
3meya4Ju1ManFN5ri/sfJUVKbCHDEGqVMW8zIdK6QQkk/ESFPyaUA9lOVGcEFVxPHhfBHeknLf3k
C1qibjiNiHBXc5mWiRy9r5M98jKe+WFC4d7UKwFI3UI9Q1jv4KII9DsLH64ch4IZ02m4n8qiQTof
0Xnhh4mwFWyYcUlbLRAUarNwfl0cOgKxt8tdCyEtr9MTUK/OaFf9fuz5CX2nNh3s8dcCdzOxS0wM
W7klcFBFSpXpdMIzj5/76j5ZIBsFdXxe2js6vySwMd8lrNmW5d45m/iZtiaD94dByDuwUxD70TfB
oFNYXD1IooneMGQSLqFKjQnJneE3euYV0lrGpoayQpeD+gWK43XN8brBpdeB4Ne7v9TKfEaKTK9q
+ASrEjllAWV2Rsitbi6kGyphGXtv+JxR7gbJZscc0vTMHQc/IM3N4UApKnEZuNfsTkPeVlM08EPG
+RCqmfKiaBmWsqUqYY4A0VBkgjH/szrhgzokrfBgyrQK6rSF9UfJ0QYDvpafr8VqIC5Dr/m9kWpN
hZmja0wQ70x8xnPMDVc6Ct7fXI2JgUWJ1tHEuxzVBQVASAYP2u4+Gi006oPGiw55XijVjBbv8pto
lL5kKiAfSypf6HovdmsvQQStSG46IAXXIcrKlSBxXGY0rJDw/1E/SvH8fdUO+h9kzyQx9076PGYK
64fuQ0XtC//r/y2SsBqPdvKlzr27Are4k5nIM3ykRyBd28Y+Q7ibUV7sJB6U2g8Kb7TEinSvtGNO
LQ5RiEjCRSWzHOGeGT/ij+BrmB2Lce/Ty6vEhtSxtcA+tDKCFfXMLyWwOFdKveJU3GyFc9/NTL0h
WRomHt+rh9NG8ygNtVjPAxYDsDj7rgZXdZzSWD0kJLoJwH7vKNN04Pmj+XWQ0ym9mDjXWm9l7rTf
0gxZQ5T20bEFw/JGBi773oNK/oyiblMC9dFsq+N9hSBpZeH84f0WdOweU/C41Nb+EkqECb5NExnL
y7rkVyuy/9JnhdAH5fNhEGT707zTSMLK2ArEzppucQTBw8PA+CrHFbnouWut3ZVNK7eCZoCW+srY
eRkpDiZ7YyIfh16vJWutaQRYd9/ew8m5d7rq93I6cKG54hfdUAmRgGUN4vs6iIqFC5uRuYLBkHRt
iXM5C25i0mybeECFsNw+Mm0CchutMTSt5bMIVVZxzVTa8HJ81XF+t6Z/e4Bc2uVKJpHRUDnNOJAf
e6AoA4Ec9Z5VVruuBYDQC8FNdy1o182+lWGZLwWakEaSZDvSTh38r6eGGZD/W8Hzqywt7AFRSjS2
Ew4K4fBhFVqUWlDw3gOSmj4pExT5i/l3dxwgw4QnF6fY7q0zm3FW8alBgnmR4QINBiK/aEgOHzcY
r7yPtvqJgN/JqHyl70PbmDC5B8Q5Zfk+GS30X7c1nHalJnVVDHO7hh7HPsQ7MRDz/IHM2N9b0Lsu
aqLa5r4BjGE1IE2WukuC/gY6oNiFczFeGB+a95ymAvdLJEKel0DtKxaboiSW6BqGvL6dW1JQle3y
VzzlIpEM9wLTzN722zg1Z+aKlHfEcaLf62e4/RLn5woMFkk9YyDNlvlfZDuQsJFgoHtRPQ7v0CxN
Qozyw5MNdkaaRM2S88bovri7fJ/ZnVh3/ZUDa6cK0xP61nloHoIxKW5xj67uGfuBya9cgQrsy3ud
IcO3jgpHIcKZJNHghgdtPxZG9XFJNP16N1a8a42ClUrFWdNhGeK5oUbkfNDBDKpcCwPTWJLW+WO3
C/OqtFY9hq0XL+pqIm8ypD8I2USv+1xBCcY8XvmWUtcjZHaAAkXLLfMsKwM1YsljvWrTVduFm5ji
/GXKXJMWoG+oUYhGzwQq+ZkIIB2UaXyeyuLfvcvD31/3cPefMBEUkTIE+XaQCqT46DB9y11/eVpt
Tl0jRaa1mudQQWFNWadQB51oOdBotPWcQkb6l7BPMUn2wx9DNcQ6zRtxnON6H1i/3M7DRApGM+pc
OHfcbI8TIUnhH/lYGvZFk1ChCmOhGOVs8+NEAh/9Q4bWgmxXXWoRIBXt3nAPkpbdbCOdEepmAPAI
tXoHRbvacpWy/WB/syGb0iajAZ7eF3rWITsGElByfMR/oWGd7WNnwrW29Tz0+yGmBHOrLGds5ZOS
6dCGIQpiVfFDezqalf1UBAfg8D1wQZb4uOGS9pl3I4WtIIZMfIElId7ukwv+x+VorIzB5PrnBq1A
WsMc5xmid5nC1EiYSfpO97pYLIYXiXiVx0KpFCtG+qVfU3vZwcr8wMq+lHpgnJaPMpWFNwZ8Xvym
e5cIO82cwhEoKEGRLzswF5xDVTOETbuDeX1lQZvu4PTcBP6QbkyB4F+3Bb9woxCNJi2oeWSI4FRM
7B0nd97xYYgwnu1AKbKoQIfh4IZUlTTGhGK9zQ2hlBsBDYBuJ2yi3yBV5i4ceSOqL1iJ4o6a6XUc
jnEamgSsXTNmGD1lBamBm9ek+pTI4M8In+vU2cNvlfukpaOqsZIfs2VU1esBprjdrCUkBTa0AmoY
STJPUSU+sJQpGLrfSeQLTWT1LuKCvU9D29Szb8uLfU9bT3pQN3llsx3l12CfoPf/oWadMPRgaHZ7
zUd8+mCBVTTeTmPSwH8gphiuFDGmH1TOmTGpIJkTXUPCiDIXJg09ZSe3XZ78tOFhFNFjUuJh1Qiv
OwQQ3+oHWwhWc/qXf6KwnfPEkpYYLYiK9Fh9DbgY0ElD0/1VFReuPEOsj5AHxtfFhQNCXTofVVCF
a2wYyh8e8No47Y5+N1nUhiAttw8/y1S8FdSPHJrmfasHMlJcm148cZFh1o3s+FaaCcUOrajNEBIc
ohkexLUecj27fR3ArS4Xmyi3pcJWMQWecHKmcVPjH2l3iHXpsSZw3pflH/BD7eyUD2sGe/+6sn92
B9Oecxo+N5Ks6JJ/8jNWDzhy9V0LPNrqvRNdpRwgoiWdjebSgfp4vKHr9wHkhpBwcLGPLmIEm4Ag
TbLTgy9alTMONYcquFOT0oExcace7GIg6t5RsjYwSuyFuG7PS0ADYzAlf34kIZT9kR/Jh62857Ls
e4m/PC3aOqGaOpRujejfIpE5CQi09Uax6AU3YfeQem5s0d1hC7zfya2xyOwXvnzCGQB2DLQQA8dC
oj4Fl66fBkpiD5Id1EfJwASJ8ctvzUkzo/+KgLVHsl2a3JgE1rmT4j45/ADKNPfks9VJ6k9f6udX
CS46alVJSYq9Vz5OWo3ooivxKONz+bBd7/suI4YQitR3OVM62gk/mTw5orKRm+g5CWeKZYH4fjYO
9OsZU8p5/8PfhNPntPAvWbyc726ft//2BM0pbDT0S8Mh6yUToReSVOiEyHPVVU2Sfz6p4Hnko3OB
GXJrxkWxmL9Uym3tUbV1ndStIFTxsJJ4oK6S2gD8D0Ah0ZmDQ+B/mS0Nk4vqOnd1GniSftyZsYAr
65zlPYSMUoULiM7v0K0D7qwj1ZyRMVE/7cP3W+ohEQhCBE3dC3drwUPpiM3aeQAoo/RmtBV6+REk
n2DPQVHtJkOHfaqS3EhcGfQOVMpnUNVlecYAlQWavopCOUpdxfBG+i6z6EEVu2bQMA3BiaGczInY
G6RVhGg3vRTsyqRfiFVkOQcRbo9fJ52yWrg2THTr7F/0zToT61yXSwrZkALOSzF1qIhdbNjB62+u
5VrEI2r5svEPeeDELBzUYPEr2vETGQHgigtbegW/5YHhEMIiL7aU2Xb9+MMv39AAlTk/tqXPVu1s
Aqt49vA9yUNZ3qa8IJPqMBhz6d/WOC/oD4+dQZf02mVAy5vP5Kxt1mVEe68LlYajjm0QCSaHTX0r
dusTq3HfPrs1IwhXG7uTueVmV/Zv32vTLJZ+zOSvHF6OJly4uwAQ+rQM/43yw/71Xrrid0aS8Yc+
+D/0O/eTU7i7jPg45UzYn8pTML4N6PyA757ugmNBKFS1TpQ8luYTFtW1R6d5ZIK6sLSTx5aZz4/c
qxJwCEoY+sg30epE+fRDZ+no4mT/sLjavEwlkdRuP4gfpdJ7/rc2A8T7ZMXIAc6jN06BqQQwqxo6
iojUFYs5dJYRkV8zt0HwN1pFZ4TN0Rcphduy44SrTLaaC7441cks+4KyVbbO9gHlA1bHo38XJ/vu
2LGK+DR5cGDH59pk0R21s67JvgtbvHyE0we9XJRWyv9eKZr7w+jbRq+tng4f0ogPDhhNjN/xlsKu
0u7bzsHaqDsSa2lc/zhGvp7+DDAeJWcHbdORkUxQBJgtOW6SaVIhVtBvpdn3gx6H0sjb7vw12yI6
WFF1KPmAHb8d+JJszg8xRizNdkSK2hTYj8sMvYJQVuBl6Xmw9kGnKfitnR/6ICzUYslbDHpBhhXb
MoZW9F9Kipe3B7Sc3Bi2gx7LcXMWR6d15gQLKyN58tz2E/mgH2PYbPVP7ydjoRwWQCMiQrwk8fa5
Hsjzlm5uiTWSI+6oBsaXfqXOVLW1WOAUE2o37d7BYMQoSw2itCgrFOPP6tS7c/fIsT1u2fZYDJnF
scLQqT5SgHsaQHhyuwJE4aOOCNYJ5PFqCPSWpXMeUI5f+Fgshe+GVudOPxrG4osIBvZgt4JNANK9
L0TMaGa2fsMpkMN9l7m0xKz4gtMTz30YovLLSNQyIZyktWLTbkOik8si+y8dxMVbfBJkWHft0dTn
O2EZ/3ZCzpvvB0QA+tp1/3op1j1xu7x2Xx+T48J8YMBC/dgLQQ+50Ua1X0C7JsPSvRbB+/thr2Qp
7Q0md1ilqzy+bJ8z1mtylypKzx6JN7DanTORkpsCCLvZr2W1sxHLmZ94WKHS4igUvl16yCuGQiLE
e+E2d7nNgHs6RRffJdlxugUdyk7vvCO9nSRBGG2dVBhovkzCapUljGIXscu+UZuuoDhXgLtOa1Wl
8ZTpmRl77t6m0mPr9kmzFQjBME3kTGWL/nS2XUBVwoS98Bo1GLtbf6wYZKLJ18JSMzZjT6MCqzaM
oz6cMBHW0UlbG0ekDHlr6H/irQxAnWn/6RsrPhUiaAJZC3XZ/BDAsQoP/+yX3RzQGHM5opyiEdwm
9lPzEAXt+okzjJ6IKe/uqjuiR9iDd3Vs0Cr14G3T4E5xPbck/v6JVC/nXWWuTeSdeMYhkTcWhjKV
V6SZT8PlqZK5ZXmRorwuaiLez0Fs0hpACpLc+onMxdB8AbjnST09lBOUCUm7yHF3YwjUXyP7V4iz
XT/FQHEYFUkJIp/czKnbJ19TiMKrg6DYS0ES0FVTb9xpUQ22KIOH7uNsUAGvoc32zcMB9CXz3gLp
9xnYlBlxZpxzHuDaNi5q+JhZqWDKGX65lAftApffchTo5e9wNQKP1D9aognNwKmtKIEmUmRHHaE4
O519Sa4ksluFTI+WqeTkXKzCVNt6m50fJMjoi/eCKpF++YW+gwoWeoc7BKLi2R0WC7pTB2hOTeTp
WWpXHpYx8eqkgs456dwzBZXIrZCio/taMeQ88oAoX2eFA2dNfWbkuVnhoyWNdvfrvu/xPZGMIHzm
3yMV1hzMqMw9rmmdOGFIUGPNmeQ55MT+U1nNerS3+WXnjM5rwWiulp518AAn4jMC9EYlCryVTXR4
0Vu+HDXLeX9M2iD7FB8WFxNgpnfry3MS4y9701wRF+c2z/WdfKEPpPYWI1Euxaa4h9trNNhDAKHY
wh02aQ5/nMqRp7/7V9C9QzynZ4wZwcY35NISNPWdUCaZX4n8Fsi6c+7zy93xMre8egVuCigdGMv9
vTEjFNce8/tFnI1L0xScR2lHD4eIuzeULO6nIw6gER17/N/sXrnk9B8I8luMnq+mqHNHg11xHUSI
ouwZobihx5J5/yb9k2hHR4dEayBBLiJYgdd9fmSSOWL6hw+gt/cy6kNc2xek1oRGKzRbuAOxGZCM
1lOVoLNR/aifTmkN0Z+IxdvsPZryNi/h4/xLulmk3fvurXSMUJ6O6ZAt1/v3TnwUWlC4ODpYDY6n
dYEPi6cnZZP2kzhEGF67SboTScjEPLr8TmOWdOZv9O/YZB0iejplMP4CENp8asoHRCzwyu98BeO4
zbIlCbdg2nnZeSj7CjZa/8CZwLQxo//l4pRsoO1YrsRaT0x2LnaKwJilbPw5e6RgCZP2IVuibF6K
2c9to2BLYNewwwL8hqJobbO+dxcngBdd7QlCxEc2+LJDUNdt6hHx9/bUYE5ES6x/JUfwoC//VZzo
PlNnSQaqQqJl1U44pvSqT4jQDx2WuAdnw2ZqYdbtMSOtVuTOdZmRAPnRT4lCEB0REIaRSHaforWy
rRBLev7jU+ymjNd37gjv73YgDy7e48aE7KckqnWIVLcDiBBEzKYSpzoi/fmerKHChV2IXhcsYJYe
p/4go2gpZe7p9nuUzx7a/twIuca69V2LBpBcmNxbXKfKzuwoiTzQ5zEmQZXZM++xM59fAjxKFl9K
e6IJjR/Nk18n1fNGPxeQlmpjbuQo7tuwrur6Cph0T1MOlWwYdvlVAq/MfXgVthMgrg2I8j/Je/JD
8u0voiHEfSMyPmvAPn/29Cnr2AXMesiTqtlE44+SI3EdCnmD7rMN/gdUJ3gRQSKrAhisUodtOtfC
K23eEEeigEHRKK3G6SBpq2pxHdUP8fMh0xv61KqVKiRsAZI4urB3iIHgdTMaipfTNPcY0NhlOZay
UuFqdNyzc9HeR7lpQQluXCKBX9aL4EBt0ucnxSc9j8wKGhvKTE51cgFbH2SsHsozwMshJpPCdTme
NQRNhcVioWZsBsRWGen2k+/C+vOu3+4B6OFATcpwqBGcDnYL3mMdfHW8xCbUcp7Vk4Yw9oJw8NNW
6GhIgjH8FhEieb2JoXDL3mc++dcPPat4u5RZm/awJNL9WoirYIUv+CRwbiXzyOAhQuKl094PiCZU
r1mhZdYywCU8rliBw3i84GBgBJxLEc1H8Rdcy6zJlAQ6TuljzJsqFq6jRZQNCFjQC7LP8QFDTYFD
bUUSNyzzO2dXksOnY/E61b6U/xdzmqdT+wPyjXrQgvN8MvQ9F5cNlCkzHPY17LKEOBPsaUHd/oTP
gu05K6OPl+1aL8cyPjg9LqDTOrvJ7NB8kx63kk0gapX1VWoctqijwgZcunu2Q+yAPtCc4OKHFLPl
8fKgIQj77atiyFrgvIDrSNHRtHtuxioZ56JHE3a8UAoNeZ+t2vS8RefAQSlDCmSgsjh2RXjVEsRe
gsmCGYlkM+OOVyCEYFhD57wu5kVnWgidub4Kc6FQgOS6VIYgxElRRSPeBdsMruKX6xw0TAl4X+x5
4qLlwC8OBn03e7gKwgB5l0ueY3S2NjmoV7joDtiYUB4t+zf69KipeKOIDhQpfGimNOdyPcY85ZK9
5WX4NJuopXzq9Jn7rH9rzZLDmfaSuUUXw+qO99C0yuqEkJ3j8m2Y/a035zCGk8OCKokMU0/IsZmS
F/h5tR/eArBBCeq2hRdiQFPkyMaApNOu/2YBLGSic2/38RsoOqhuEHeo1JQZaTAu4H47/SFQWivo
xnjLR58QVX6NHrOOMPfIw03Psojhfj0cBHdXtGlHAW1KDUC8GOP8sqHQlduIryAIa6hZ9SnHf4a7
w4YfAqhBobBcZtbYeKX25NF1XynL6AKtfmYkVZs1xNquCx+ZnmyYcDDAK1MIPXiW3PAVqT0DihFt
CJj0GyswKkeNHH2mzMBKKcxFjHgTtGjS869GglUcVY23nqqqcIQX2A1c/FyGcTcRVxO8Xjrq4AQX
QCYocx5idensdnn3FP/LrQ/3MNPuN2O01Kb5hfQMv1evPc05HGrGUcQ5dTfjdXkgV10H2K5KwrrP
FZ6X4vlGmhIdUefrokTBTkPi7ZiC1unWKShktZzxAJZ7591IHjIqqSHA78fyMyWAkj3KVZzBmJ2v
tSyeGNQaHWSD2TmyM0hVLk4YC762AFMXOYUmnO0NzE9m1CoO49RpGlUbS9oUzUU6VbgSDVBW9cSM
/+KqfJqIXK3GguOJBytjeuyZiH1pYSAdOaM3E4Ham4L4QNJFm8EonjoSglKKi2Ljl9sSKuPdLE3Z
ptbeyR0VJjHXLWz7+AYVsZXl1gba/I/WEPobzhiXzJj0LmxaFrzXGupFga35lDIN2ZQEI/nzB7OB
qEhAR1XtgtqaZSvnGSS4pNE3/gm2cawSW++BniFGIKriYGuqKqfE1odj47thrfNwJgG66CsAb0e7
s7rajzGuye2NI7nnCwH4jXcT381YjdDQlwY6h08xKr8AQHnlp4L2jPIHOdXxvbeQ4+MCbW9v4CPH
kqYWPzwZsreGvW43M1vW6TtyVwesMAOZVaM6LNZVIMZGapqVOywNLMxVgpXAMTmTHiY7lGNAUlu4
nUu7ZgLaZTXw4fvhUkjBbAyzpPlPgYjwyf24DhUtZCRD6X7vImil46KOK7D0HdcWkh+McrRnrFLE
KyFKJWZ+dVJKLI6UMRT1JidbJ0bOc+xJ7Tg7TTzcIf9r7CAD9NE6ND3VxuqN9G9PqIlE4gRI+lu3
XR0sr9UKDmmg4y0JTr9INB2oTOe035+x9B2YAKl3Oivk3nQhlZgUaf503CHbUytd5QkJ7Ixsfhky
NNG4ddlhMgtS8+jEpnJklFRos605NfCR2Aw6YQmmM0txVhQYYeyWSemCmsVwqTLIbJ0v+JEWnOzK
plcSaPYlay7auoNGWI9UT2S2gHV6IT7A1q8HrNuu73Bk5cJfNcycgrWUKPdyRaApxp7i8M0/sqgb
PfSlaf0U6ctN5FNTuEqqdkVzaoE+qvESNlmz77orR4YHuY9ySXohBMoJHE6xdr4JNPaD7R1pyjGd
XPyRAxjHyZonJmHP0sZvuD34zRDK5l2QvLTDyXOFUoL6yyT/U9PsXaKgOwKOwogkQEqXGa5OBOxG
4rkTJVb7TP8XWtvfYq24M7y4aMsI7+zH45HFTXewvTlQbrmlF4tYuoZeb1bDKOWvjq8Fh4k2BtCi
iZxA0POAn8YNH35WzQsr8oRkE5EyGesaW0a8DQXOvbBp49o9hMhAZ86Q/vwBfSeNEaTKsoHckVWj
qgEBx/zXNCJNQTTXQkbW9rL0TdqPii2bqmCaUkT5z6dcv859ZDSP+LlcRXftXzfF7MVTAV+ZlFrB
jMMhBLqLQguiU0dleD2lAK9VxlYZ6ttJIRQ6d/xhwP+0PENVPRGE91wHDVgDcouDew46DQG7+Oh/
ViSU5dLfC3sji1sWy9mc3lG8/Xjd5Kmzt+3wN2mqKItCixA+BmnT36qt31bkcxzvLZs+S5A0IvyY
h1qNWbj2t8PK2rN5da+3P8xXdCzg2hPkypPexSYHPWOOaaxmYjX90bha3N+4ZfZT88v2y0rYZO/r
ajFyUIHBqRSZICHWzu6Hl8JKSbAT5CV+XhAwzMc6fwefndSgIEDMQu7JLcCx8XHUiKKgIZBLBbrc
/KJnN9QPuEps138DP52FjKvfTZqaZp1+QoYsh0IVdCw9IZEZqOI/vvicZiSP4AFGN/dwdNJEYOdX
jKS62q5gCmAtOnqNA8nHInHb6xi/Y/BLvRDYRhLHUKJD0xxYRPVmnqm7zYnJjn/vTqFPHOCi2Axs
Ko+9rI5m5iaeJhcnRGl+HGoo9kjbGPp5ss3X023fND5JEMM22Eu+j9GTfMC0lpOyEeIFef2DK3z5
gl6Wx7zzBcN5/9oIiTmmD7lxqZ0/exicxS16oi432ikgWyC3cO0YPRBpXHjE3BIqlGwu1PJtAqub
NNtfrCwXdxWb/Yvh08F70SpzrATP3fh3lWaNwx80KBSoGP6rzlph/XA8pbnCG5UDaTCXrU2v7+Pi
mPK1SqSstxzJtVOaA0lHYf7rvZUd5vM7KYDAJ/YKavIxIIH3tt9uLioW/hSOQR3rQb1KgyfxSRO4
drRindk0VTeGC3nXFJxFK7wzopVqLo1m6R439MprdMsmwf3wWCGA4cebBUw5rXmv/UFuonMZEuoV
xjiORp4Opv2TDjPmWH6tO9vbwmAwSqk4cCBafidRC5GBn6rK5DICSsVay5/LzJdqdYUoUsjb4vVc
2UNWeSPQrISTZ166dvmme++FyvNEfpEJmqFtYMHQfM04/YNs1LzqZxxqbV/LoN0Y+fKGjYLGb8Mj
3hhthcpdvikWwhvVPwuUZG84RZNPfJLfrpF84XPAtLeSgw9tndKJwkAf/2DzSrMbfn0B77ZUTv4+
hVg96x7HobwY1QigFrxKai6QX7LJct4WGEV9LT6+w62lSUxxyfyXn+Bo63Oe0Vh96SisXKKiAx//
VhABRFsuAkUujD7rzqYKZa+vch1xTe4M5BPqobn07q8fCDBmlbCb8kaMgpsL+Jp947ghh3yy+1Zw
jhu1Qr7/PIgjgI4Za49LJYFrvDTpii6Tx4wYUfhFfK/Iqd01vtgWDKaVD6TWj5v7Lt/hbT6NC0ft
IbWwTOTvrKDOvNUmdJXHMA6ArPNBYoBbOukZjSf+QexVLesDM1BkG+6esnWPhPfNE5pboy2aq4cz
dARqMrKvIyV7sREKdNNIKCbEpmFgIB6F/hLOe1Z9T8Ose/WGENxL+FWuTFVvjD93PeCGBX9SBc4J
A0+1CnVlR1lRqyaUCJcBEg4Qfmq05PdN5F17rEFHwpJdgrX73B7ZBV0o1dBZbl8RDkcthpfhRKYz
6NyldUIDgtxiIIrRPWCqXSeVNCoGnNf9YJ3UcvbdwKFu0u4e5OL3cyKsCwWWzF8zTwTxhCkuDEaq
3ly3UZvApw04G2cOEX6D1X3GteG+lonUU4oBqS2/vMcPvbWwZEKLNhT9P04m2hmhRRLAyCoUKvA7
jbhRkzXO2Uk3vsUhdWHCsulxaHJLUm57wUFLSs604i/NmYLz3kBBThaRAx9/Z+JbYHbkm8qEr8f0
cKB9nxUvDUT6uYJQ5pKq2hsVHbPeqfwlQreHlHekISjqGCeF3LljZZF9QoIc1H+WJFThWd+xRa0p
zyjk2Yd6/nqwmZwYk8gw/44BnKuRGpUou8LWZDbgzFHm6zmZ6sBx4Dnuqm/BAULI2CJ6CvIklfWG
8RAlbvBvZmBiFfPzybBa4qHqA5XqKqf9E/kC87A6ZkWQG27NFGdrkRBCxK99ozybBUSy5b+Jdkvj
02CFQiqssy1EhQdzJHAzDQLan/dZHjQvUjCl+NgYCRodGgkh1rE6n+YK/+Z+0DWF16BoKuFGxHs9
Rk3PstWO/QqRmc4RjiuvwuPdUlIm9p//exzjliAjij3tqh7M/MdxUfBqlUNgKs98SpnP78QPDWxF
5vubuWAABdPifU+I/ePckaY5iqEMw32u6c60Yr6/AqhG0ny7BtEYxQsofkX1jBglGi0gf3dfVdRU
6+eRWVZLOiiloLPZddoZyxewbrC9QJwRzuRP71g36dRELbe5dTnIGdQ0Q9iKEB6Vbyuyr75yhNSn
Yk11oST/gdB3WRnABNnY9x88lmRbiXOXxAu3PZDKApx8uua0ZJcjlbRCHqK2qRLV4uPyf0CEXYID
JVo4CRVE0Rir1nkGGYozkL+Ix3YGs/etbRHJ3RAV3qwg22/thfmFR7vSlzl8ruQP5mkSGFaughss
+ZlV4mgLRQorDOhZUJcb9khoJoqfJaSQnA40EYYTzmYy0DIfp8M5oqddN8LegCc84+iXvZO0Hbhe
ofEIgyC0Boiw6mh31b5P/FuMJkLdCRY1ed+faWBuDfDjUIH1MVxNWULgCLG83/NjkuIwLlsTdkmz
QYQ8r6loBI4sUnKxTiXsNsdfQ8lVLd/13wYfTBR69P2XkRZDJS/ylJ9avkzObFH+NuMFpRuZX2KE
C/wRSemmtqIH3qVCXAhy63Q3/mMYKlmzSEQ7EuHlfCmtOVuqghctDBuF86yQxpGALw2/bdrNr4hd
NSLOaAnVx28TJMoLsQqegh32DL6UgFtl75yvKHgbtO+ssdOwMQW3ajuEOfn9hqBw1v2avVk8dLCZ
rnX71XVBZTYYziwCZ9vYeL2YA9dJl+d1T3A4O+QY+hFOHsUo5m5r9e+bM8/spypaXfjS8VyvL+NN
dV5NGPP75iujpLRz3dV46a4V3jnJhjEFfEB4j1OS76nW7y12A/YYWgGza1d1HEmzlyn/ZkKBmaPM
jKxA6Rbz+cTFFnhon7IdKgDewJuZl0naawRZOmS9wbgrTQSSiiZNpVbW+LBXX20p48AepwxFEI5o
12KWsfvB//riRKxca6AgHeg8fgTRAqyQW4ThF0kloOIoNvpP60zG487BgHOnsSxBTroahNKHb88l
sAr+fPJlFEwmMdzxSpJWlIVrsu9I9ye6xCkiekyz+TZh0pjUDkN2/HHvU1fR9PCp2mnVtTpfegQ7
Hml4zv+nzdKMpIDem+gJJWAWAknD8Ru25tFO3epYYON4HwGzndelkc1MIoIrP9/baiDZlwvKD8Ne
Lv5XemO6SZZCbgrOPLpKJhustrO74yUnasuTgCcSnyI/UB7iZFc/jqi1WzgzqCcXBiSZ4Z+Int5r
lvwWj9nn34AP0YiQGVzPBvEpbfmrVrTd+702i8nehy6JTvbO2qmk499d4jKAfcDurov50b4oYxOh
17tQ1UAraJKSeRsBlvlqkwYi9M61SIEy8MBagt1hVA4NLp9ekC4+MzAaMtDgdMZapVAP462mM3jt
jMqweDwRxndqZQXmdRKikeCcjbS5xBUdzQYhSP2w04z4QwT+Bmx7wHHhuOkfVe1FUgrNgFuI8jsy
Lis+jpcMalLHfRsCFgkhMnzUIApwU8LX6shlZ0czpS/R2HF+my1nkKntbbBn+tAMG3q8qD/KH+Gf
seaKqKGXUsCXynQcwBPj7wf3YMclQ7aWK/3iKFWo1qy7X5/7VIVRSXGWCkvV+WyQRl53uXghXn0h
O/nitgWOpdPaJ0LuzYqE+wemd3yicxByePiLM+eL3c8BnML13GGvp8JHhh00iBXhz2kREQlZaKVo
NPrv7F3EMPRD00qG3BFGRmuAgDNWKR9UAdsUG+G3u7EDsE1PMcBglaZQeM33gzEhKU3OALOmao8I
TChj/KymtgBQmS7qiF1LCEX1OHD1f7D/dXfZLvXD+SVtF8EHi1CFMA56YmhO1Qqdg8Qf6ixyFRPE
k/CyBK3NTHOJOekCELUU9Hd7xEAmVd69HfpzRYRG09SIWh1lang/WvBMMdL3UpNyoj5la9h3qR4j
FjhEjn3TAP+Xde5z95dF5LtMc3u9CBvCjWCMkyUvhaFK+8GmpMNKgylqaIOYYIpc5dP1Jv1CqgDJ
pxBGNAlZawupMfUsyJ9w8xFUeeW2K6vSHPN7jnJLt2OXU78UrOXh8PdHHaNwSeemcPTTRATn1DNy
66zd7FDIzxXlqybS49KL2QONqlMYaM9o05sGrStVILFZ1q4KPJPiwbMI6QIspczrxZCnDrBYeqpD
kOgHcn14ljV7dpgO/dzdE8ewmHKbxYK2tMeeIt6rA86TxtyVXTGO6uXWmqfnBUiiIOLR2ocVwAVz
PKB5FxSaO4vKZrruh9puqKttOeNSXtZxDmSdncWoRxN+ZBjtmS2CAyrm3cYXJbInND6YnaJYQP7H
OC/hJ0Fh9UKlgIuVSq5Zw6U+hi7fhhrqv3Jq+lJWb+kIAA3+6n04yekguQZo4gJO8rsYYKD9nKWY
rQBVfWCKmdB16NotyjO1ziRUQCLi40MAUBE7nUihBkv2OMOnCCM8ToPzLGhdXqGqDZEnrdwtmUBx
Hw+i+xb4vNB/ksElgX5LveGBf8nhrvNQAeh3ssSqjbqykRned5OA96BnyiJiKJZe+zDv8RPvYlYn
wuaR1nhhdkqt9MYyqxgVHKR8Tb78DQihibBN0TzkybVCpvOLG2FsF57gfsqQxgA0wVP/JTJxf8Qd
1a1lCVoePn3eTzQaWoCdScQlqt6BbFv887maHIGMom7L6gez9j1cXQBTK434/u6BRfhsixyJrQO9
P6VOf+ILlXS5d14eWND3m+X1d/jF+iPMY+w/7PYse5PgUNtiFcBMY32BiyLK2LsWPWxx/OyltJBC
9nENlID/hC+0tr5c6EsgkVlVYAmFe9dMV+E96nvhN4iWf46EflptFxWdtsbLtR5w359Hw6nooMMm
lH/aRlgrtvSey/c8BXZEBXOK3L+FZpSoRRxosMBkx/9PTPdn4CIC/y3xI+gt/xbSYw/WOUtUUvsK
mMNm/RObB5pDhZs/3oOSFKB9xkUyA6fp/0nysunaAqiWSM2xzhIG3Fp7exu20AVi8flJYcyTVs0p
LriKUq+aBnzq0OBJIn/S6EvLexV1pVurLYXfv/sV4EnNWbnG8Y5VchWGDXrt/LWiR1dJHYHE+nDZ
2AL2FRzoY7DPCoizbOtbdsfhl0VoZ+nJUPP6aJXPKLtDY1EpQantSYORS4cVNhom8JX+2ZomwUyN
r/Q5sbaQaBSSYn2A8G+fGGWHlsJekqo9q7kjfM+7PWcRsIoMw3b3c1dVHDxTY9VA3k4J9dzNwRyR
SwMYlDBe81zQ6Gk4sVvPfaGAcRUqkudPguIs1LuUumgCtt/x+z3hpAeMK9t/i2AbV4YIU4h/+B7I
STt3GnRSJDJQ0APRYu7jERPLBXwwizoQXMb/mH7z3nwpx2AmAaA2ReeftryazlR9zGmuJOCIvWNr
hfA0SsmNcfzrtUhdKQYT1CosXF6QCBeveqv9VG1J9T3cOVjJ+t7lGkyiT8Ckx0nBFGR4QJwTmuqg
axN8FSVL28+AxYo1ro9fOyf/15sKB/Dw/AADk/S9JBtrZxbWMN2m0B0B7Zzj2r4lFmUxz7Ay0cTC
I9KBCYrBDrjpPZREo6iiLSioBcl45W6COUaS73Zy9VeP6tElaDOOrwdrCxuH8e7Zny94mvUMF+M5
rbsaB7l0o4/cRkhAFYom/B6+6ThGDuHsapz0sTzbHrV7D/Vt7JOcvf2tD9GrowBquYO5qRFKS3ju
/xbQviHcd5ooGuOwPhXitG74lC1CPU1IR3ltaTz1E5h2P/nvft8YlZjDoVPlws+36zOOrN5KeDk2
9+w7pjYMvfY3uXWax8roQlArzYYryP9U5K5F2p1Z3f3IR1DD11AGR1lirAtypSigFUJ+b+cXjQT8
LVS1tf99h06I2mGE9ELyq17cVpb5F6ZHqIhqcybsrgWLR8yrmaoHyiAdcZYzXHb27qo9g0l+rqcw
XvNp26oFhYiWd4hMYy/vx9WX8htSqg/S1QndybfAQoMjZ70Mg7M8nRj0bZM7KOHcWlNHy74hdVRh
uMo+TiUfqoPEXYZREv3Ayvi91xTWrYEE5LGhVxSSd4qmoIUr7U+x6NiYNLFYauVIGvb7v5iNr4Ra
+s6teA2mH5fMzk8PnQTsF7rSJ+7eM1mcxhSbUQVx1O5l20yA4WC0AHTgDTzAc9BGO85Dk7LlOlAm
Wb8Z214TlNJowR7a1jOiFPPgsZurOM3MJ27r0IveMyEGKH37sQuqWc4K95KYEOaeaWqo0puZG4Nh
q3zgtJSpt5ptgIN6K/Hc2QeBAxwtuHFE2HIIsOXKXr/xUI6pcD11pkmFcnh47GMtmnxHdTsCPLWp
wnna4wijpeN8F2OT6kwQeTYjXsrY88FXccodlx3Kig5bLNNQG97bKRBXiQXt5bZEpoJ6cIde487+
NjaVXLxQP5JoxbnuSrUFlzg4/6lIsUgKAUXIUOYPZAbPFbIhrhIA3+L2SsLpbn+9jAgQuBloNs9m
V637zLfcT/R6yYyPbbqxF3KqBhEdY84+9ZorkwgXL/ulHCtqFA2UDnLKKf5RSKu8/Qu7OgtSjDOx
st5iIeDYKkBzX+uQZ6WOEC3bNrW81A/kDcBV+D6quX3KQl+gpNYXuZBWYZLyAiBIFH1YihQwTe24
0N9GzAloWxJV3NVyeTOFOPi6JyUX3GTiEq6W+WcEapEJEJhtbqtZjSvOQTPeMqQc8FjGgZN2/Jrc
Gq+zDvy5a2y7pT6bncGqfzv+HSbn7rO2/3DV2osIYhDKE0GG5lttJlsHXBc4Xsn14kKDN7X2bw8R
qjzF+1AjeKLd5hVilPWWE9OaVkA/OztofRxTqRdBpBB5NtIEYhjBzIDVzs43WLLCtTIlCVepuraR
jPQuxc/fU4nmA0/dvtOPvLkQJBqDyvfpU3gU1yJT9EqEB3++MfjUrv/fkk5lyb9l1Qf/wofuoFHo
LzJJUsAbemiR9rDvAUGfRy5Jd4RBaqFnCDYmQmIxSXALH77koE5zli7bJtUDgbM8W1WgFaI/kppD
TiWzAO31Ud0g1icTzxb3LHbv7eOzLxAQ1EkcVKfGi0WT1K5ex5U0E9WOO/NAEVjc5XTqa4gN+OZQ
ixs8V2W+CpykE1C5ACJ9n1o3d5DFMDG0P2lyfwVssQ3XMd2VRQijGJmpx8bmtCzlFD2vecYEqT4z
YpVGOhiLGPAKGVfwKxsCjq9IViUdmDvOoYXfB526hQJuaPJeHUFdqdq8QmNv17L3i/fC0y7j6tu+
cTAeOrXwFUEzy/ilvnIr/zpIaThvfEOhJQrk5kiYuyH5hpq6Up0vI1RW9o4L9H7xon7g3rHp49Ae
lCvbH7sHYMunxk6UNS+gag7hTLtK8Q3v6nWNzxRgA52h2HeytWfu1ObPsSIDOHmozBXmbOg5HPaT
24QocLc9e59W/he7x2HedJWUIHCji4l7xPv7L84U1iIhi3tLComLDhFdIDpRiXGYMjn4XAgYB8vG
joZ93wpPribKzEjqI1gGxMVX+R652aiUwIc5RBTCahakRmejz+ybZvxZdh4HgemPDWqB1gO3kta7
euHjTa0DipOG7pCSMAU8hA34ASxuFyKEVb+ueoNmP8p6Q0sv6KeQag3S3DlIHNJuPqSShxSsVmjI
9lQWzwICydNZ+iD66PY3exU7eYdcsBmDgq0FaMlwG2JmEFAdvYM9wnd5VP7fd6xtoO+hsprA3hct
MomqQpSQbLSmzufysQ79kAYE9LbmStTAZWJ0A4khgwv4huFjcosckA415uTpmx/R1nKktE3LLbaY
oynh8VF82hQXomKAoFVI9sKKL4YrEvpFsKedAiv8ayUokG8dMeIHBtMmkJsSLwyv7Us0TsdpAptz
AUDIEY7S4AGVtCH7ZnD6tLSpFfl+gWg5qPA5IuLCv9QORpOfpncGMxkZeJM7W7a5T2FBnqyq6zwQ
9m1moxxdnnHKheM4Z+PkJXS6XO6ZXdplzJEHZ7R1D9eido4eVf5F801r12mFR6mdYv1DcgyT0/72
5lqtOQxJRJJDbChRFdiMbfLDjIOL0t99UwCx2JPC9mtuq95A/OOGT6YC+/yCyjv36oWLhgXRIIlF
kJxcYzwaqglqHQ9I8n0X3rqUPyIzRcSst5RuH9ir8klqvM2sLUoSnwaADGBq+ca9eQ6h6Yb5oVrj
+b2cN8ZI+egb39F+yDI7KO98kqr6IPmch42xsZtHtfEbhFHhqc6n3T3o7LvovOb8ppSqmZVaXTAn
3IuxKiOxGcKYRSyRS05CS+E7aurjuS3g9rw/hfr1VxvPOspbT6j9o4JniaENdXnK4AclaSUREied
dFiH59U78KxLKWkQC3EV2lkG16XZdUVZueyyxbYcdMwg4wMWeH4RO9vEN9/UOrNKMZcE9XtdLAhm
1P4qNsQ5zbH2G0AR44xDfhjLH9nS7QY3GiAaA8XsIIlFkv/FulNwsDqx7HewsdtnHLTulkIMlHaI
MUwpqP3HjEGNz2p5U4XmKjadJewbnml8RIR3NdEEa/QSSfSNuBYx0HPih08x68egIRGo3/zEHJPp
Jr98ARtIXHmw1zd2i7WgEpH/0iQFNGNE+Im1cdIr7bUrBjTBXazZELcJG1GhOoPXNWw0+sLPx+jy
OHYrJ+yyrNuj9FzZhwwGI8uR9Od0WKlPZ7lsSg0nyoYy56y6m20sE/L6TJjEQv+RcNgZfQUSpcFs
fdubhxrb14bqp/PiWZlraIPZZV4otowpE+Vmdxv7CLBhnmP34dEo2j0L4Dr/dL11UZj92t2s7eWp
9ddUjUe+4IXS9VElepjAGo5WhkBWrqU0ETvCl2zsd9BAAz3RNRFLxaHPpzumvKpJz9bb8xDfgmHx
5cnAj2SWVZwxdX+ir+jp7XInZhmy/sO1vQrY1IMACg231G4fDG/VlxS4jJ8QwxuvKCE3M5gHDrfz
XusNETf1GAwhH2XpvRUGnMvIJMcEdKOwxm6cngdLdXsST3mUO3eH9Gh00SjrlNcloWAZMasuLzNm
VZGHBOf9Ip+CXP+pjM8o6MyVVPdPfo6RDr9f4BhoodpctvGUTvgWWE6HilcxKCRKcr6HOeY0qdTp
rLDZcgw4xnJMhXyMTHdY0pgudEzkhJR1L0Pjf957j6eDQj5ePtpn3UgqrUzmr+fUJnVc7gO69dBD
tvC96IhRutN0p33Gqz1xub+quyXu9Cx1ImgJhAs4xUcmvuHq6osN4dsDKqPBpY3A2T2K6xTOQ0V+
tRzx5PSQjFfzywvFszZZz1y8v+rlqIvKhU5ZnQKZdXQtGMC2gcEx8SpvT097Fw4Xfr4FTGG0m+/J
OcKgGj4R2N7R52G6rOUnt9V4xL85y0uCvKmgqwsS/Euhhn75TBGNDPiHUI3fa1Pq1nU2hO1mbylb
Ral8ydHKaZCdHxXuVBFG+ToflypQCqVhWF9flxYIKg1mSm23/j5Y4YKPDRm420nN+Ne2T2lrDW8m
i5f8A3q2ppJRCH0pmbruBUzBjTGTMukh+290S7Wk+QYTpI2JYpmMSVuhfyaKGfvfbic+vxOxq2RP
C68eXTgeAqEfzl0xdP+ALhmF0aRkK5VTCp73TmKLQEpEALpzCpIrEPxhUsF8MjBnLttkahIwijeh
9CsvRTA9Y7wtH/OBq+lh1tziQFsZkfSj6mgYxBc1DudjY4nKnswab04ZxYscVdoaq+0CjeILLvop
hAhv3Riilnsh1zGEU4+o9m2ufNZTBXOQVLJmAMIAWsWRhgzLxM1XQz3KRtSaHggz1WOm3NhpPExz
YaKyTp23kKOsKJgiM9OE5BvIMZ/gOz9jCl70WHYiRq7RbyXIpVJfSFKl/NgRI2rpMdgVEiFX9LmU
aBqpkHBHcmzqN+mPwRfH1wk10Dw52e09DsL0yEP1WDibPsNtFbNuGaIOuwSiGInMtnV8QxuzEc2Z
jkCyGwTT8sx825chRe1rvxZkwvbYXHsBPVNKrfT80vR7T1xns2e00rTOlrpUpxlpq8Rxki/TNlQ8
EHTjZyzo3iKEiuRchcqUOTcXL/qZagzJW4oj3yLcPu/1JE7Fcw48D6ZN8jY9hFCgn7zTKRBmeASq
U00CcZrMU8aJhXVHRvT/kmPWhI+9Ii+fV6qI47ULyu0TCt0/GM/D/dt/xggRkwvIohqGg5cBCkjS
FIs9ucd5eY0oGLWnXVBBpLKCm/ywlwdX2GtHPMG/m8f/vhJB9+705d8m0IXi37a9qtPjbOt921Zs
m93W9LUiUO6P/obTTaXf4tkvi5HRUy+ZX5fhtQo5XRwCG5ez3asuJRLe3fPbdTUfyR/SnHxQYHqr
bgDYqBFDdt3Uvdw6iPzkmGwCcp9mhE2QCzxrKF+4STYFsep3xrqgjH18waWywZmGoBoJdz3FE7nZ
xUTrwJDroQXMZNfMoGPcCs2jL9C38V3pnbL5FNbNgx3ptmFKbMcEudbDUSvHGd38433BEtCPTgEZ
JMXQB5WE/mW+DVmqPsVfGZRR3KO1o5xLvK4O4tsR4lTNyxaSh4gw2+ReZQi9EqQIfMvGBcC4+G9Q
rV2y16ygJaO+wOunUvr/OU7fo62N+CpNtWTL3nHhiPcd1SuLprwePelqmV1WmvKHjeWqio/NDqHN
+v+FrrjjWoAAZSPLFCC9WFSFFnj0ZKo0kR7wpE6GJv61+vlf/cIo3hYnH7UAMe6Ph/AKuDYd7Ara
Fqi+0Iz6Dii1sdn7Rzn3RsGXvy3PVo41RZ6rWnT+sL5CZ4MqCKEbudQyxz2cR+bISIGZ15lv7YIs
VMKaq+llMdSHzbVT8iRwxeLHDmtwPhwODjWGb4/FAfC+AnESz2Eub5wSO2YF1Quq565AT4li8IXD
9fZekh2CUOfKrQIdA2krac8YRZG/Qj7G7uaG9OW3fGLnaDRm14I3lT6WQOBWNUv6IJhCVzKT5RRs
nnzPEzuz9nWw581wnPoB72HgyjZc08n0OSg6/NUtb/CWS5/Vw7+qF3CbGBtUyIQla6Yhxc7iaE8R
R/Vvx3blVi3U3lq3zcAThoP1gPCygHZqcYEWo+4s9q18Jp28EpFUXYDHWGtocPbUbo/kUaVIrNUv
5dHYq2mlohuzvLldy71rFYse7ruiCnpkGKdokXrz/wnpL2FiZxuca5qWAojm/dpFTmKE8eWch/ox
/K906ALZVJuEj7cj5NkJoiH+ye7nkw9DMrbqY5CjLczJNApmpK05XEwY5bdA4ShStDFQPRk0zMwo
vpy48r0Dp9tPtq4ZpYAn0+Igovjg82SefkVLSQntEWhZJkYJk2I7z+dFtLZkW8vL0p/gnmV/qtk4
TCbexzTFoN7asaD4iBQeekUJZs1dgyFAa0JBXvFD7SIEPFJ6UTAQ9xDlSS7jq3w6o7X9CG3BaU6u
bJHUylRY6GTFT852WK4M2q4Xiht3zT73jo11RFqH3HPTscRAeTjJicjWcS3KlYPM8AcW+hEdA6Bp
cf0LHzRnNdcQsFAiyA7StZ+KM/9lzZABVTXcOwl0aqo2hanSbxWVMkZNDNZuQS2cKQ3qBSOdKLHn
fJLe+9fyGi5F3BW622J6EtqLy21oYABd9+LiqlUB5mygkZ7r7nIVOGYopH6Zb+U5s62CiVlEDbKV
mBtx6H0PnRmQcnP8jNvhDXQrCW+eQxKdjnd5v+6yZHruDKvnDCAX1g9O0CrTGsYohq7IdBK2pogl
HZxEVwBPa3M4u6S3KaSHdN3H1/9zESvG6u7aUHggAUBnIYeY9G1uI8VebZqawalNIbaEIWecn8OP
EFM2zmdu4AS1K0P4e/LwM4o3uvbiLJknbcp1JEph/AlLQcJp1KcrX7WlVPQ1OSa5NWfcTSmOKNrE
WALWie8PrqO5vptoBqkyk36NogHM3YTsYnhN8/3guf3iC43t7zb3HEWn4xZBDCzkmzGmlrrA+BwP
Kg/WHfkkAkviDnuQEqkIUQaVNp8rKi5rBH/ac9PfoCHeJTvIsNsKCjAlTZkjjIopcpFhBKST3oEC
qLfQc1KyYEbtZhRlxutct/d4AFnMjpB4LAulRtzQzg0xYDPoZ51ky+0KEvuNEGTztd+BclyU9zQU
sDra7QiA24cXCOkSs94gh1Eu59DDZ7k+iNg/HrrM09X0z9GkgefrckEq68I/H7+dRuAunzlPlfNC
cVTK1pk/4NiTK874EPD+p8ex1YHv1EnkDeIuWc+khWxJYQXepwzntWTN0sMj1uwilGaLwlqibGQV
uWnvAVTZv03ltacM0NhG7uI2vA7pYk+vmEyrnpREz1psHkD4/epXNgiryh9EJ/QG0zAyJ0EE7PBY
HM0StpLOBludPVC5/CJHhY8OqFA5BDnW8fRlF3GH5nLBhbe2/c8Ea9C2dCIg59iw7NqsiTFMVcGd
XZjEqpw1VnMuWnRbvF95qAFMJRgLbtUB4u0aXecwRFhtqNH9gvlyjY6t9xAkmxbMScDUVMWfDIJ6
XTr8P4A9V2HyCB8jKEsi0h+wFxWxn9aFomkHRBF5XJ6bifMqkudj79pZXPrF8RFNNIXSZ6rqU+BB
2ESZr7yfQV5h00xJ5EqMk3NOTEmrgJRXOzJiIFUoYJ7m+VBz5rGy9PUvZb8c60GJnbJLOmtcOgAs
2hk8jpvMxxpOA71pDGiCAg7He/I2uUDeH+3aykQhNrzdWlqb4+RCfVs1gIWJoloOQVNa7BM4ohAg
Fl+VGTSn/OVcdqN1SSJPhgtp9RkujHp9eYUp4Wc4zMQZuqBJ80a33Y4EJ4gifT831vTrNJDZjotn
8b1YYJebBpOOTU+rUsS7Iy1Ig36ROYOkjiAZefoNzqnpF24F9995bChbp/L23WmDO6A847MmYb5u
xBpbj+aGNkX82EaWXrGASgGp/80FoODcBXlE7c0P6e3Mhb8LxF3WGt7z2PfIrUcwEffwfvniQUWW
ieOClTslQhYS+E4ItzckB164Qro4hUSceIPjB+ON+bZpxMdB7S6uoidwOz48PUDSFtCn9ckTPtD3
waft0tNPboFrf+CLy+o+UBxPI6WN6cUvzPSft7t4fmOD7SKNusCSbaloE2dX7eKBNiXb+qxHBZjs
d7xNqvcS7tdWY5szXomvc1Ap6iBnQmDZeBpTkMKz1pBbAYx5O+C1m6Yznv08WQaykWGucnFCR59w
KFs2yBn0WTU3f2IHBqg77HSB805CtX2O1wtaO6SQgpbxIlPkl2VQNiLpKjn4IvVqvmOWcnIVqh9T
PTyndl1WHPYB3wF32JX0Mn06mPF3rVsNQiAC4yVcjEaiLOevC+5gdFtsl3ChymMdiCxzS666PE9s
GVZfX4JTXlhftAE3VRTM0dkHiWJvTu7LFfRReP1v751Wq0PT0HV3qvwKJVFrzupCOPcYfADjG5tn
qvzysiASK0YRTIGhHoEeNzwO/EluSKRTnQFuMUOVh5UKizvy3DcgWiSukgztmz9RlyjnG/1k74eB
HjklzR/M8fx0J4VOc9LhhNrioYlqI5ElywnYVuVKn9WagB88AY0KliewFe6fLCh10b/0v8x7ksML
t5g/C+HuM+1iK99bAbITt8iTw+kT6VPeLO991M98nqkuMGtoWe0JNjM+nZs8GLQApJoo251QBU7Z
cSOTzbvBahxtYTY6C9U9rE6U9D4RLhENyN7x3WTts1bLq18wJwKiaJujLpNnKnWnswMKgqyH9HYD
O5AyiWXfRvZVi6Pqyto1uX7Y6IHLTdQhKjym7KCHh9GOMqGwfT6ll4qVHQ9/wpk8zBbSTNX58XgX
qhHxZUbd21ZWHPbEVkfGxjo4ieQwy8Tcyg6c+jJVkliIaM44oipfvsUArY+WdMYZwChLNpOxzlXe
DUspaXj3LQdd1vVlTQxE35+53vmOKMV51A7ZA72X/vdrkg69p+soQymqsInIjcm73ZZApJBwCzI5
y7n9G5gq28EwpcX1ae7lI3ZJti63kkQvF0sXle8dA8SglwDy5oSIj0RIL8GxwYJ25T+Rwz85oMe1
CpO3PnEuwTNBAzjPg1lEHfUhSe5WcHR9/tDr6kPnPn7RtCdYFOT4pq4lq/RozObJh/h9VMbJ/bZG
jsexjXWpEls1Nn5wT3FxqK0UjBWIV04xeyMmPOzRb0RLhRdKXaCu2aTHSeCx+op25SruikPfR9WV
E1cccaAFPHTJu4UA0FFoTVCpiomyVY9QQ8lb5bo3k/IT308+NEeMMmv12VmBN0/gjUTUY+2sC9ug
WPEFAOGbyTBzMbvPSyOVLMq5HG/FpykexI0CK4tsnFHn3vb54uO5sZib2TYwRaRLcRYDYTsUn5gG
nxt9IZtyNNv4kT/MreZb+lzcak6HVi92sQqBN+N1oYELAs1Zab44IBBAb8DchRaQ/nvhuxZ9/4Hf
ngybV0eSU/m6uERT1159QG1doS9BmJyaxckUkXe43pPwKGKjqy16FMWZbl+XxC/ELcwQecgnRDmK
xYuyQ9FCSQ3GBeUZa2Pjk7Y9pfefCyQLpkaqG/we6lGHrNnDz/prcHTKAFEqr2WHsUd0YvLCHUpS
1BRWolUdUayaxziJx3YQVBk7CcUQM4ZirD5jKGfoEUUTgFu2WuCveoMVZXh871xbmsVFkvgOa7jW
j/b1Ijky4WZr/YByXEF+8g8RuDvDF1Q0JfPJfpMePfO8vWCT3LklEeIs2t/HlJxMAyKj/2in1KsY
FnMisMZ95XyzJY1F+9U3iTkQFTATR2CNFnvlX26/NVGQDZDui4muz64RwCIc7wtD6IcTkIzH6LXn
9h3sBWY5SuABJWPtb+/nMKbtwIzcPVRv8UIWNlXySEdOm2rSGvHltvP5mcik6jknK/D5VfxH874l
Yf1pSXU/dm092vyLcnobKCYrwCxgkm54Y7jq5rXUW2rMaPPyFqR98FoEy4rE36nMGnZWvky/R8P3
74LWwbJeGYqr7h4nbAD+xEw03T7hq8vDCyFseB0HepdlQDdGuW3sSNGFyX+KD2luwEg28HtxlcAU
DjAdtDEa+gZ/aMwxfTHIbbqAzn0RX9ZqS+W2p6itojJIurYmiH04OjnqssgDOqJXtNoYrD7pPzCm
BxHcVak8wVcaVWSuQq93c33dgeXw8QcNVGEuKUdxFMqXkVj9cY5wgk7chhT9vjKK0H8n/L7P7k/I
nGybzPHHaXc1z7pT02+GQBNexPqGx9WhKW1r/Vb+t1pGgD732uvnRJBiZJ75zJ7Gvl5biNWvakHn
rnzuUxK6f0DQADputj0FgPX7giOSe4dvx/lh9UwxDISqZpGDokI7quMJOBVwvfmIdYAPUalhbszH
KFFuGsAvRJvfKV1IRU/icTv8Aelq1+glcEhVCsTYhTNhgjlImYYrisWLRQPTTFJCxC4RR+6o+OF8
HdDeOdnh2LVkQVl7DUqXLBZas/0yoN79PdWkjQ62JQINoUSn9QjwpOVOOObIIHWySlFBMI7U7yIA
IU2crcJmFYm7H2OUadpwvzTSj5MLkpk9+r/5zwAKuD+KxkwYTd6Oxp9uM2v/n6hX2mPF3GzlAwgD
MPu2vttzRh3fpS/WAWFJZ2vQI9Sl8cnCqhDDgfl85AZqwah+Fnl26DwSB5ymwoqtin1t1c4d1ICW
iA3WdZOFR2zrSCnavLIHCN1vVCUjjOjoUU7pAfJBMhu4q99+CvJ2K8XcFb6FlKkpzKz/TL0wKfE/
3Y+rLKWESU7+iy1Cs5MTYaI8Jgw3O5Tdx2HUzKivqd/OXd+g1wL0CbWA6CWileZObnGjvNWZPZbg
SDnq8aI9c2Iqp4xtAT1bC46OzrAGVePtvh28WK9RpwH8LV4KgpfU8buYRcKNbptv+L/RBokMPgNX
QkFUYUCco+wgDtW01o5YQj4gaiqimF3SSsLzrZbQtwA2dG8cWugW08nd3rDNp0zGoMLNgwcwV70Y
ZmmHNMZXbDTTgU6iPIuSswDEk6ov2+Q+/hN3f5ArfBWHr1CzrW1nXLZn8sA8voVtVyn5Z+Z5OvDy
NypBbOFAAffEht9vfeiGWMo5zQ3Xs9R3u0qrHFoe+j+IaVTm7K+zmU9Eg6Q05kUP09WzK+C1RFl4
tLZP8ea0EZEnz9Y5objMLJUFdJmB2z0cpSdu5pjlRdKDeg/1t0V3WS71opxrtOtgxWv0Pn9eYjgK
B5zlwn+3V2Pby/TUB7KR+Ue5wXmclpUY/YLPaiwBGOP15Jw2B8GBN8o53vWjU+QiubkMZPaeZV0M
6s32QrWBjlJ/CcPchawaa96Kcs0ow8Cy9gBHrDAEKJWsJYfAJNobaSriqXVIVl+/GFxYyb/BoweD
lk3yOFRAToXMt5gKVJBLSjPPcIxh/LwkEE7EA9OuWplyLvxX3e4hVWbYFnKb0ERRtKFbNg8k+OTm
bjJ2q/tfrBwVPLRu9AL6X0HITF2elcyNXEthrXtBio6miOlrucfoLNMsTDtRpWPkzF+fAwmcoszt
YYHQxkEuqzQdyQa87G6oaIx/cx8xXSbb84EI7v2NTPXWmBDlTqtyHkLjAmXCVSaHIMLOUqRawUVH
DoR7XqrbaREpmUkUA2JF/pMsw4GP+oBuWuYw+zS7QEjMm6Bwe2XW1Is8RsemPAeLjQeIGj4XE1O/
5QWTUIKFOwgWCWCvpk2kBu9V/FZGd9iNLbGeEiInUN4UL2Y+imOFzDZvOqZQZx2uw41R8dwVTQ8u
0VISQXbt9VThuBSFA8CtYwEYubPzxA0b6F0mwlbXU8WhoqFvFHv8ML4b7q2D9W7H8rtTagmgVput
plfpTqfDiNd21+AJ8+NtkD54Q2+MREHi6BqpI9cSmMmpH5a1vmAgcUKv13wYPdlJufyVYF2dkraH
Mz/4pgxsXqEyMn7bA47HFk2jxRgmIrOo2e93YYY5LtKBIeKhygE9H/Qs3rBQZXDIelhVtvs3H+8S
P8ybHRhmulKfaeENX7jabytv+PrMOs+e1oLDaAYSqya3zrWW3+vvCVbhIkpm2JtWU2GJMKty1Yvm
Rx1/8tC1LmDfYCFn9xtMYc3+5PUrOcmXySnVCT1bh+beAKMMD1OdMSPj3PfZESBqKDF4ulGY/k14
wI9s9TiKZSjf1Q2x0PNrahfClJX0yDYqY8tiPM1Z/HbOc7X/qirccSbv5Zrb/XkVRBHSt8Na4/Gs
MdU7A1S3XlS/r03vTQpsnZxGbVA1WhqHxGVfNbYM7HmXu42oCAnAE0uH8FRVlqCaXRfZXo+sTxlZ
aNyo8HcIXatg0zZQa0vVh3yZNvEbrV5g6pakk6PbovL8TqgoZsTHQ00lfVW6Tjhly87AD6/TULK4
16MH8EgYyha7H/CQhS74fr5u5IR51x9r0KW91kcJnI2uXnnTtTmjUyjR1opBa1QeL6+GYes0kOEn
+xAD93XnB+jrmYTO8anQa/uUo5F0WQpaXy36EgDxizSgHutWuictP4tcsHfdUzoMmSLKpipx+pC8
Yz8mUPN4b4O2DoIgeVwtu/IOg2BgguIxTQawoc3FCSc/Z81nQHrtHHe4/r1WtGgI28J+4cTbjHwh
ZooDnJjWsqVsnwWhG251Zggt/vr51/Uh0REANwnQ1G8E2TSRL8fpOCDbPtQA+b87ozc3fzDK7T8l
og2qZWWQmTeIEZ5h+ONXnaCDFe83z52nFUvA7qGA7bh6k9UNKvEkGH5LDjfU4HZyTqVY3xR5Pwj8
CH6fyx+wWrR9536YO07vTJZNqXeS06xrIZNajkIHrPHlCmcrTD11FNxbQuFEcehZM2is4ORsy5nZ
m9bijhFlGgkjS2m17P+U8qFL5XJZTsLWNNBlwddYvDAN7ITGpjVfhWn2ngOmJofeMn2ijFBk3MDH
5R4nkiPctmJJ8HpxAy4IKowhak6Pxvmpy2ZdZ1JIE3kd5O7ph3mJwWRVavBrsxNp3uJ/to2Mt8Fo
w1ZVKmtK/UKJHz992AyDyrkdR1eRNYQ5Cg2gGIWZy7dmOCc0aSmXnzUEz8xGso9Okgyt7goU7YRa
DchU5kcfFI2lxWrMfQ6oSs6nxa34QFZFHpAtItoREO6jbahKsT77L9BVCFnheHbb+xYxMxOWScMY
AwiHIV+LKdhJIqg0Aw57EKHQoKmbJe6aCnpxTYA+DV79THor+K5ZzAPR1vwmHj/T80QJpxpxjd/x
4/+hvbjn1qXahq7QH1/ch2HQ1R3+HY1BlF1+mJmAyuKSKVMUxMM2WAet86B+X9ciC4S4lYA8W6ND
E6QVqll2JRrTrWKbxtL1rm8/nc4Gc79Io4rgrv8HswDc+1rrzKqtbFjyO2rhxI9CqGuDSJvezcNB
13DHaWlBWX6440u2t3e2zau1ruM1JfbyMlLaFxWZTX267pDbjPoFnsj340/OGlCZsNhym2e30EDr
PIIlHiA8E6yhV95CjycdZW4/80puUSCh0zRfsQW8krUaDCXheVtNczehIWDX3+ihzX5OdZvzTo87
+/s6wO0pME9rtVDIkiJ++9W6W/pogSo9jcoNoyqt2lxYKWIC0Z7SQu45Wh5+bKanOujuZ+qe8fEz
eRZGMFceWqQ+9P+jesYaPOTLPQVeMOkrQDbAGlMQkcbsBXzG8+mCaLkTJbyid7NY2udvYbVPU9sr
bZEyRnNxJvjDP4Lqzg9b6RfXhdjUeA/lm6NTl+105LyF4Mv/gg/ZusvD2I9jBNeFh7u0tVpfvDAt
v4S0pODPWs+GxQpTVhFSw/JZDmBfwrgP8YRJRJxSlUSUko0NY3m4Bys1wM4KT6hxAKx4uLRVbeub
+Ii08psiAa8G40mwHDroKGr3ZiAVL2r/7nMdleHd73511dwuthyNIN+y0P79cVL7cGvbNKXS2bqy
XZGQk7p1lXgg94DXmpDYqfyCzvN5s4dG/LZr64WkDbsz0C8wrRC6X/9jQ/8ztWET1F0w4R4x2Jow
7qKlmETkPT+T50pFe3/VRVqZL46bCyLGx5nyeSXntXCdx2HJ6Wf36uVD9chN8E1RjHFjeORDXw2e
KHM6/bgbzyfu0Kizn5R+gl2T2VKktF6L6pKxraQtzam3cF6OALEav5xxpzG0GZLaDefM4XpssvwU
tgfdAdAxXYcFqJcPiyNj5UF7lU4V9Xtq8VS0dn1mJRRh8IMH5VRalX0fJkSieq8sed5ND2180iRT
EQsN9j9AD4uRU6uu2ZG8knQyB5rRsyZQRXwewLyR4mch+H/RT56LhMIN7C70Lj4gwe0lY2znFCpd
SMcgLlL7rPQBynmgklh3tg5fUE6VH1Hz31pCVzf7aI/jXyZhhXEraHGOAdeSGwuZlF7cRSGYfgS1
Cy8YOpieFnKpDA1oEUzHPW7MaTeuP+DDRt6XIDFHBz2vVO8M3OZZ//g8Iy9/HBzjxvW4GlHzdY4R
PwYBL3t1NGPlPGZRHjDMwbYdigcQVPuRdL8Dl4Yef0wehgWLPmg3p5wt1WNBEgTVBTTTsgItGiz6
FBTYCpJqqxwcd6jN+FlmbrYOPZN0gsxyQK7bwkRDM3PdVzdLOkZ3ePotep5zMiTUBOYODkdX0Bcd
jHOs3cgl5RQ/G2gqprTJTc/xZ5HsZaO3+z6UMPwZspDZ2+CcFC74Dx8YfUBGsFDXsXuOIQXoJS6G
s4zjRCEJ+Uu73uUMOO43cTFFUBqnEBUq8wzHkSb2h+9CuvrdDQSc+cPQZ7HFr06kp5TZPWmHg+wY
choSkoA2gy58oj5byDeJXmZ+4NJ4bbZzHhIZq6ZgZoMGFq6nrIppdXDRC5hLZMTVLAiv/rEFJkeD
dMJBF8BGDU9x+iJ9pTXZdpDOcmJr6FauSZ5PZ1kXyXz235cpnabfkYxfKBTMD1IiHXeHp0fX8PRP
a1x3oqHpm1zuvee8v/3KVDQUvGDMf8EhhApHq/6+fGcWaaYSY8SeaOasGVqP/vIC6EhEK6tbqp6m
H69chaqIpKFqYdbvOXIrCNF2yDmacEALbah8XmZFGeAXavhJ8hTy8qEBUxUfdHAEc4bYEYNx2ooc
LuJLGW4lc1sat1Vrxu5xln1aDqkJdPyKeJoYYAr4rzKXDlBEYqnnReAXgb+nX4s/RPaQPLguJmME
oidn6CxawMrKX4ZYsuyZ76g9rvMgaCEgR4ILIo1DSXVR0ACGt/VAuvCQ7oB4PSbM8P9uH6n6xThe
rBEYt2kM5WFqX1P2Gx2al9Ksp0AHrn9foza9pxzg41WwjczjnLjY8cUvIFtqihRGLbVxPZ5cH1mZ
Z+aiKpKbiuz1icosYb0efukl2xGUXby33dxeQ8M0HeWiBOw8pPJJjBRmy/cVZDvNZ1ZmYQQQ4cZw
ID1x39P/4JEhp2ZsOJnPhoHvV4FqiqFnEMB2ftSjHYoxwY4uNEDqMf3Wp67AS73N7zHKDwrEibei
+4UcmmBvLv7FJ5l7EcSDui/waam9bza6h2JmfFp5gwHy4T4izY2ZJh/DvMaUEwZ24iQcexNAaEyP
MkXtYd4bGtkDmXnn5MU43PSFMMiTYIxOxk6xhso1gPXucuxV2ml0mH17CprneMwU4GRJ2JIQixS8
KrF7orZToN6dbWLqM//05irLShJLtL4iMd135IND7iio5srieJErKtVfeysIIZtQAjJqCf/WOcwK
L+ixh3q5AUKgyx6M4HVpVeRZu/peLbfo/poEbOnt4ERM4GjaeKnS1qCp/BFNgj9gAxB23gLha1ux
OHQsX0ZMyNGTn9hchKskXPuDUDI/ajhi1AdfJWzWVfTQ5tELz3riNXvusuPSbPoFse0oavINpDBj
nGLa+csY7ClXSvJhAfOw5vnVEGKWuy/nei0bf7rwqMe2wrviRjEXNUJ+zbF8GrMXbQaoDnPH8SF7
AdXcpvWjqj4DE5pJVv7scr9iljUGg97+oHLvZrtvIDA4PEGfjjjQP5TQZYqrc60RVGYgsex75r68
qqP4w0of2CIwEhqAZp4qJ7W61ZKa+mk2uepWcukXms7vPjQfOqnyA+aJLQYMXo2Icn7kxbbiA1d4
X87F8PH0i7oVlhmYVcD0ymJzxQI2XsfilNO39BWvf+SRQzDf0wdtu96DMm2cGQa/8noeoypw1c9g
ekBzSj4BXSNoX8SPX0unyQ9RlZFt2VhzDU0mWA1m4TEYtUZw6mrt++4991sYO9SaeqjR51SzuU90
SEhouamhTWO/B8Rp/ZIngSkh7OSNZhX2KZ9wTO6dOIu3pGb9y29c/CLkfg99e9hNytzYPCn7BGr7
7vaBtQIwK6SV31lLJHMfh/p0ApPJ57MwMuqHd6Oqkx/FjxySjX76hQYnYYA9H/OeUeCvlyEJiQZV
mcxntjygLCRbOIGOVWTB5Tiy9jTAlQGlEbtxYDM/kWoT/2dM+p0fCqPChGQjo39r4wpknOj9j9zH
qKbakGrVG8T47aF7DaVMENaLbmRcSSWZPdnaJhfTeS9FliX9m6BapFkfkvl1fzchQBqKP4LOAEPP
OatG1X5E3SeLTZQrsmVRp6zrYf2AoN2jakNmFw9n3gRjuG0sjD1e7eTaiQ5ByEFnipwL32G2imYJ
oD1aaujfrwNI2gpYkP4RNZp2KD7oQfeeHbm+Mq8YwM+OEQzFljX6YYv7GT9bQi1q/iRDUv94RY4F
rMh/NJsKmXgtjo4eS8M7ie2HZX4ES/gFqAsDv6I4ob/63Gi412NXZbzecXW3bc9NjUVPYV+k3Ga3
4Q3sLyK758IEKV2uXNVFuSiX6aXBwdUAUDHflEO/Jm1A3JA1fAlk3+N677yevk3SE+shT9fuvLRo
8e37ZUHN28lTXrfwvIgasr3aM6sVx7cw3cZhqi82SC+mxj+1n/J+gJehlk1HA3+dFSilCVhYixsa
pBec0ZHHucwkkkpU2UZR9XUU5vS1sADwfF5ZkLWrbQC3965I9A476DbU///OEVF4HSUjreuyOBTY
MBRFjWOt7Man4rubOGmhxa4KwOoGyshNEepihKieT1B+PgucGJGb29GrvvcAVHlLQjqMBFgi6Hz5
fjtWHhCp6JlYRrQMIQgAF3x0Hupse7J5/v/quZ7BRRifQ/fGawj0It1NZIqM4wLZBQ0D1rdUiQLs
Xkzf4JRGJgf5WosnuDKyb5bqe1FBkBgoa+oX9QwtqP9MHA4lZoiLF2jc0P5UdU0Ft2kSEzYfSmHF
wBT7acQQP7pkHHH5ZcCS/A6UXOJVMcLwlB7Mdjjtv21wa9lmCWdWtLMEjqNcFrEhA5VKMNzqmrM4
x5y0u+yZKyifYnkfFY/pQXsnyZgNL7+66qkwK5X+N9ybSsmXVVgYBXhnPtXyyAN3E1hIhY6vi6Rz
5byXXF64yNLd3NneFpYRNO5/4mkB60onJXCYcogEOsoZkEHZ23yw4mP9MWnySfLsiJVuBDcPyarz
6gn94UnS0qP5dGlggZLDiqCoS/N5QLGwYeT3tCryjKrXK3yjSp9fxXrneI1y+ZOqwKznRcg332xh
gyxavbyM1gVV8JlVdxynQrllHxtW6Gqvmvri6W/GowcPYs9MdByKJhnDBi3iiDD/HGdOOUyWfsbM
UXuK6UHZeIflSNZlTsn3mTTJt7Ul0sUYW6LZT9/BD35krwEnaU+2jZLElJDkBLVwF0J4EmOfX2s8
etE1SVwVRWr6arP6ILhYFNfPWs/LAiRWUsunpHI8BAXS54pVIYpzTBwEHpylsA6PmO3QJWwMUvrb
6pazsfOqK6K3um7HQQuXuTh302qwIvH6b89FfLSLueqCiA+d/59za8/M0Xed+Xo5H/vOSep7qzow
ZRGRmgzT7XbQkYSQ4r+5GPsVHO6pBR5mqL19MiDn969B7RL+upjJYc6kPCLwRMsXz+lU4EaDaxoI
7poPxys3bkb7UUiCcDaiHQgHnRhzAeEw0/a0jS6rjZZRw2knnBDRsSBN2F4PZTwciPfuP4wrC3kZ
M+JOQ2igVG7JA1a+aWxKxbQ/iF2nVdbg6y2KwJCPuyrVKfIPqthx59j3+x+/y5FPG5hDG75a86YW
UBaiPSPFHgNAUUxk0+3G0sbF+w9Su+Ysqe03PO8uC6HqLd3KZDYRPKgiSndqBQ5YxG3XoKWGKjtB
bKrWtIfhPZohTMPO+dSnD2oTZoDGgG1u4gvODj+H3+fSodkJMg5UpyDA0W3ct7QH0ycfOXlTYgmi
Ox38ai9vYkQYaqHJzAToJNNZnAaGKBHyiZe886eFl9GaVqf74T98yQj6xZ4tR0lAi6qLb1v5INpE
GSPFF+hRWK3ORFXKw6E6NCiQddxz5GKyLlKTTry2k8sE7nJTSEoSxg8zTMtqoxQqMyo3Kf2Azl6g
5a9L00IVdjNdP3Lq+GTuvljxgr3xsll/n+uSJBrTG+AzJ719aPYOWZlGTilyTtftCu4ZauBLMLU+
GUDK+xM1MzNRlm7x24uJj6JQkWp9efvvqBKyxP5XawqfWCbxZncKi/9EthraOV9LT7sdWXVH2Yd8
/JEqonhSfN8qiZRN43cDaeMRpKFXG3YTSfvYBDMhmFkB+xoqTlLcwxJxjEERD1tcHuDZtsk2KpIh
6PU0YZ/4iaghjRMTBeSBpg8eNnYw9ptSw9quBrafd1PdNvQ1vD+Td5hMMBEGIYqW7V2I+I2HVx8N
Mbtz83AD2MoMjs3eFXpjWBCjxVssEMGqHy+74GPN2UwvYk7P79rggzczMFZkjaYw3T1P/b01jl+/
bo7svQ/R3bCo5jRPKkN+RT5PVxikMvDKgeYkm2zNTQ9joYbeAaXUVoBgEHCevVQM/l4xo2pktwZJ
5B63GXSAs/hu8gnShXGu5eUjk9wTYvG+mnYtmEyK7XsCDZgA5ea6MQLsVwhXiJYtfz6/R8BJVQXj
Z0jtt6UFNyq5eSWRYMntkgAi0rT5Ag5EF/BStEfFoj98uYJ0pASsmlOM2/wcmk20w8BgImgDbf4T
JONNfEoidxJhAaXZhieehhUrvx9zNLXcPoxUQHmrhxjX/w6YQGLB8cit3iED5oxByOx1I8BvlhtZ
yzKpDtmdvyt+SWsHjXM4HsAEvYGxqjp3S7WURbci7j0D7cg2P7PnIeHoq6RU1T7+iFXqAH1/4Hzm
IDqqer0sDWz3FlGefi3OsnsDxXY2wbsgRnBTi3PQEdL2SBhjOdX5FoCnJEjhuy/TFFpAutHxo1Ii
zGJC/MV/T5Muz5xZmTH55WAiCIhy0nt0qJzfN2JmFnS89chCM4FXEPVAWP/DM4pmKl2yA2RhqVSJ
m/HKx8FC1lUzCjZRAZeIxns7eBD7xmGW2lgVd1oY7RTOgqkCaQuCdzpUuTeS5heYzgRVuVQQWsL6
Oiy+5jXSRfn2DPBNzHEBhRPOSTexotPAW6Wv/1JKe4ZCgg8idLtVK6/329G8uVhMBfe86lNOEUlr
HTQBXxmcuy1YlVSSoaFD9zynl6/8vLNR3vT+oEodIIWrTNIt5bIKwuH9GGZTD3gWZYdoeq5p8ATA
NONeSkD+rQ22uWZgIEYc3UhAXhoUkD7WH3XbIXAaZUCefNrOFPndpBVKZPvcJLCzMjoxHbBBoKs9
gXW5z619zMStcdpVhKG0Jsqp62mMYrg8ZBow+TyfkzteslgNp4Ru2N9tlks+w5lbx19W2NZBeb+s
aqhch49rm5gTvSs2tDlcrEuSuylr5CPRLxZOuORjuA1prgbNb8ra4EWmAm37+hDomWf+iNAfPImY
2Ikd0o7NM2Ev+njd/kDCXvlF+LN6UxNWg1GQWurkfbK8PyOrW5DOYEy1HlZ7pareqBzJllzrcp1u
9vcbIii9mMznfragOWJzEzfky5ExP3zjhvOExvfJh/ZES3CR/91eaDlbQCvLTJg92Rrrdk9xczrj
wiRnp+UkZaldTgaQFroQ8baYC1wYR+yIbfNhv4Nfe3AsghJBhLYkFI5Fj9r5C1jDpxMrhAYPGxS+
bEj57skA3qilNy/3TrScSzrYwjhGCcTCBtYi/PD6Ny8YLOkZQbhzuf35Hd4ntc0CwTb9Lh1OKH23
fFNVJuzMtP+VmTggbivd4aSdqzDvPLSkEjuTxi4K6KR6cWGmQbfioh7rA6TV70ekeV6po3ZyzeVT
OPdQQ+IhU9D0COY3XcbkmPUX2wqpJqd9RoZd+SwqCH3Y8UVIAM6li7zRBdKkZ1LRwCW8oA+S4cMp
Z+zn6kDVdq0fUionpGTV+zRFUvw7Yb5NnpgCS5dNvrDq86sPrBYYs/1w9BRq1kmTszO96WrjHhH/
TbuSGE97aHtenc4gn2caEqu/sxIVc6HeupdC+/l2Zra3GqoSCoYTzDSO9pqVrd9cI7ouqMqUVDOV
Lb244ICM79KroEQjLfK3W+RmH7nrOq+WsysBEehF8mDVmJNVwMshMI7bY4JDVZNIsco0PnnlD+bX
KffG3xqtu6VkUJBTfxy+ptuYPg1Ddg0hPTofaZht1t1kR1BlJ6iGd1cGTu1NqfLpSltrWLWXOELB
b4dRz/U5jwy2ijHsDnDluhe2emw8YKS5YyNkZJuv7zlnJZQSi1eoMhUuw3Ti2j6/HX8/PJF6nN2e
4EASYZi1i/y/8HUgMQxagy3anSnMAS5ZbwiI139/06Axpu5RMV8fY/vxcx1v0tLfuPMvEmAjs9oT
dRaycSkKLTRFsTDGGIKu2bSrNF/z7g8rFD8LRr68zxa1gajFYw09e1hZv3AOMpnfClkiZXWr1cic
Khw4sxhhfpruXO2tIIXfu1WjJo0LchxWlJ3C4e7+JvzRKFiJ2zopX4oNCjtxiiHNQ/+m6u7LfxOo
hkGfwYRfLvux5VrKhuU97qQiVIrfedzXr7IxmoQTNul/hXINQr81MPjc5wK1bav3JdI/gWG8zH8E
OqcwDkIAGvR2JsFb4tpiy/tJm6z705kEnzpcXjSsv1tHH67hLwXdgXjpVOZfMUcRg/9z6qDm+dV7
DyXVIbJunSugw6ElkjCJTG1j9hLTjhoNOyY8KeIZveMvqKgHBqXLbSVEtATJTKdS+yP+WOFD3PGQ
Ublsp1h6pA5qjdYTmvyPI1TXrjSIuwV1VKIF2jap00BLScsAdnGxGf2Mbxb4t5Ie7SxwOEdf1HrB
Qa59yiFSVX/AgfQMRJu6YRV5bkvjT+BjGHB/gr754nogGOlKvpggQzUcf+4Ifb1aaosk2DFOfD9F
HZeEiSu58iVizTzfeByH5DiAeiSdIvLm4hU8MyT6pduDhZrCbdLflRSKHOVwEhodXzCYUD8+DedX
Cj4fLs7wFgXYPcK3PWrIoobWHZFVNmRcgxcEDoM8U+XZNsqYgmt2ouOsFjXadhINje1Q9sCIJQJ9
hN4ETXBO3qvMTxA7F8kaLaSXgsSUCybMz4kmuXLXO6eSnPqpK8m4iH0NaKi1ddS6PhRRgQLWrze+
5amYfVpYrI9X9iL+5F6yq1ePq1ZEvg4xI8+aj2jJTzwsC0V+fUKhOEoIOFR8xqkOSrpULwGWu7Po
KAFdeCL5fViDw5FslWVczNzl2R0gJWNjWqTA6HkG9e+BgXeBSwi6KJWLg5Zsur/4JXiLzYY7LezW
ajUQFTIId5hgpRQTDzCvkkltxr2EUAMGW12FEvBUwpCHqAmVHUZqUIG4E5l8JbLX1N861eCEddef
mbJ4gaJQ3QCdUwvwclgaidmCYNBYrwQZ1LaOuPs1tamF8j/1ria49BMp00vp+JsU8RxEhHfCoV2q
WgrhMoz1doSGmhnyFEHkYYCpi2WCoJNa0bxVZ4n9Z7SbNWOY0TpHkOXZ7js/gymivUTZQmCX9qQ3
H/1KNAjwbenf1mKHHOhE+cwu/fx7pU9MkUEx2gMspeGF1ZuUgNyraTSfHw8bBznqwEIl4KAZxnyU
UeBnwZrX3lqfFplb5LJJVFFbB8tdRaYyhviNndUu/ku/FWYOKcIlmDvTLaCJehuFoP0jlOD9F4+w
fBlVZERo1Hmae8kdN4MrQuJjShDT4FY5FaQ55L+7HmbG2CwJuZm4WgLdtIyammnMG205o0WIrLyf
kyALAbe44tj76R+vzkprW0iF49EM9omH6i1QmGa8O8x4xbiV2+v/YiK0hrtY8143K/tGhRo16X+L
9mSWHVqE77Jvl41dOeOVj8neztwDbCx/o4uEs8AzSQCgeLG1ATskDAr9yqiv0Vcl4c9RXLyts+Jg
jyx8qID7U09t7tTzl+0jumqVzX/k9hy4L+6Je1UnFyU28PW12V19yS3ls0gBFRPNh6pu3dng2WLF
DiTVzvBM69xi6FafAUEuI6+gHrKo3O4D/SfasYg7kfXyHysVsMzCgp/IyQtSL56YE+k7jaBcABWO
SX+H/p7Ic4ESeUqRTpPHzB6XKIaxm05na67xx0IOwNOEwAH3+iXXAlwo+O4zuMNq4qRtng7ZhmEa
A9QoEY2HFNrlhIkuAfzjEi9Rs460t/7E/dw6F0xi6D2ohWPxnKPK8rHcTu9h+8fohL/g9NcuUaQ7
MRMV+aE+NA3n7yeUrisyseTQHJ6xjiT8/PeqsMod8MQoikSfugNIJ4oSJyz6JAFl3rlDzUx8OzYN
D8U+OoPG+UE8OldRkdK+5BSZF0TsS6/cDiV8DQ1fxVi4R5ZuUTRj5BV5bzfQVHXys8BYHTt4lQ1N
dbBJyseEK490sYnHZx2k0LMUK/KmD2xUxXPt1mTPDvDUWxCAjqS8yLdJ+GXAyZ3vwa5dBhApMFZ+
CpvGQ//uYRsci6YcuYcQo7LDtbDM4iN8BgEnLth6QlUuKoWuEkgQ3/0MN0Pi0c2itPEPYDZrkcWz
r4enB1wYC7KvTywzyYrBYbl6N3Vuvb2f6rMyZhp/NIxLtkwCP4NU35aF/AaG96Tk+1gsbMQ3WSiw
NfytPgMG4yvlIs9I+Jp06e0vSC0fREyZ6aQnZ0ltAK7Aw1NIyqXue15VSxv09kwZRB+HZFbSN2gM
fF6o+MBF8p4zDRocQKFf6K+P4Jvs8O0nEFQtBFqXyip04SYLMoe4/J9NHXyvypzx9933mqfWBmCs
avap3yqAJZtPxgneqXKFdbaklgtv9Fg/59QAEFMovy2YH4ZclwlRQcN17+3NLFAanAPGx6fxPjOc
2RAN8+vM97TEdp+ttZ9R88CM6siTS8w7uBR+JurRko227MflO6S48m20QXx9V1sY+0zDyUPG/9BN
PRjotmT+SXX9kvcxqVCu+RCXoeWVXXF64ekYRaR5fn/ve9d6OZtk4UNzXmgb8+8HBBGG2UXufRo6
Wm8vKct3H0iGhvG31ixqa4ZXxkyMTzGMvmrLbNn7MMis30rKCcsYBUuxt31h58F8T4ouK0idEfXq
jb9cvFsgESsgVqhLW7Y2AZqTZmGJzNzz+zb1gsw7C5M4f6CwND2em01EcECIbxBo9bLSybOO/AYB
EBko8roNeQeYa8XjRCL+yuQ576m+DDA0O2vDq2sWXmsU9P4rF5HVvIntPqmZz8b3ZUIPVeg3sWI/
YRlmTHTO3jQEikRS6Neg1iBeN05qMt9Qa0Pv8dWzsG780ftBCjx/2FsH7mt0qW6Gn02ymMAHlBu0
VKxvz2e5Vf1VKGJuOmw+0zSz9nyleOMvJMkh3PFsRWR9p6HhZtgpu31fwOLGdQ2lzsdl0Q/sY39C
Cqz7DIcTCtrsjp+XISuuwRS/J+SbK/5PkdaTpXUiugj5AeUVh6XwWavSOzmVNzJxqUqVyffAV67h
bUj7nGDnWx73MiBrPcfaqq5ql/9pHca3y6NmksCckvbCRKSzcbk9IWsIAYFn9nMAHFRJ5m7v/fhn
AkS9tU01s5BmZ6kGLv2bJ414LjFmLI0NQU7bg4d6tj5SyF7sWBhcLHOov8SZiAtCa35YIZKkL4Ci
J6jidQ2ikdx6bPii6HldqcY4acIod+dT4yp3gfRBaG9cQcig0GRW46TA75CRZ7TA85g3Jkpo1TVC
myjwxbcqMxo4b3QKMyzQplxajQq9A/YJ/rV+KVttBH6OrAnlXvXOyYNy20FBhnyKpJ1/VaUybf8p
M6ed5s+9mwmI0qWVr0l/Xkf0qY74WuyRwpiEqATNwVkL+cTSHMxVQ9sKVZMEEPUCb/9XdEnKT3v+
Zar4o23ikQuEnb3p3mZh7Sxdk9er5h+fs+r98feMRk3eAF7eZoj1XJV0qo48/awqg20Cj0I38UV1
cTGihfnNo7IjMRanrovQiEg6gYNOfNIjo0Gmc279ecS+Uo1e9wWwMqJq6U5A/SlQAbPQmZyVY03C
Vj4hxnBjhxPzGihZCIYsgttVdRE98XDghkebbzzCStPQwWk/WH1OY3Sw7PrvKTOPHC8eCiJCqWHe
jtOqXQOO1WryvPfT1lFhURhk9+ByKbqR9MHXlIREpwWQ80EcBBVRAOyQr2E+Zuqp5O0M3caORhwX
yPpEghd+y85P8AI4jIlM3lPnbetk0DMQd4SBbedXuDS8KbgqknHNr1K9iO6tOuGI6qZeHzcmgf2Y
6tWWdJggxVXfZEHceCuVPW4ItK0sY8dB2JNeTD1zucOt8z3n7LvJIt+XhON9e/GBsRRgen/y/kU6
sOjnMqtjVUEY/AhEsO8FLGRToW7FnYVyGKzMDdiYI468oBWbp/78U6gGblMkz+mJ3rRzpFRMVqRE
FK6Xb//9c+Q458LeiTo2NLbCJyFdge6d7i1PcYyxT+wWCTTYNk72G01Ds4cXUA/LgMnRYK4cIyYE
/7IISAek6+b2L4ivxKu7HDlhe9v8nBygoaHBB4CCWAwQSCoQusG+OAUCzQv6FIVKQYjLsxDWCXLR
ti0VuDm5WEWMQ+ORaF74kZ0Jm1qRFF2Uxx/WBeCQGA+cAmY1Z8sIOsNmrptvKq6wANzuYG0e3O27
ZI9D8YnugLk2q0Ij73rdrwWNiecBX/PBj9LvLAmeX5Gdehp/dn3qRgKD//37JdMzqPxy/S1gXIiC
RqPysCN7JDpRe0V7crRsKfP1FEAxPVGOPRQYixQrzlHSUbqx2gzf6kGgcK5A5YJxSUWn+3VvQGpw
zfzxz+fmrKUY/nkZRU6czIjRuVuKN6AmZ9rjvuPni9NRDI6N4qt2sFK1uIvTmpLnDVPZ2xBG9GuE
5qORGLJiH7i+TLZHX/EexvbiN+nrAPIwjxYMSBZS1xgxLIPEgrT55pwgh7BH3M1+6owXWSCgfIQ7
MollHifqI7CiEQNVkqL92C9kBTxX2CRUS4DX6rrJfwgavFazhkamb63k5zAS49uY/aMuqWeF8fVj
z+zCFEGQ0SGmS/N/q0DezNQd3qZwnwvOE7ZzGFVBmN2dLlVNx7Zzibnk0Yjj3cC8MDxqz6SvwsHR
7wdnwP5cjs3WZoYbghPhUUsnQGxTRZM6Bl/5mMHgS9p4dj2IfGJc8DrwpN6zjoF11G1utk6w9Pca
4LDTI+01wlyRPVa8mKDBA7p1bNH5ntt4EOeVF9dklQCdXg97lpz1ej3W179HlfbFg3Mes39IXU1W
Bgsvggmldxu+38q2feSITas2QpySukNuHDTHeEdxBjJpxcjbnAqsaSVACoWRTjsLmg2appYIXNMc
fQM9QK3oDgp6uFz2RvnVe8GJhwGhMAHzcAph4PPp/FG8JFcpc5llxR+TQbbCgkGRD7qA5/0WL8Jo
djPPb1RG9pIYgGKOxPkxi+9sdLvQf/JDdRn/4OZwXlYn1Sv/gcey2mO/5wubA9JpxbaD5VHhDzmx
HhHAyLx09aiycV8+FnlpMfudItASYbHT55zIUKV+zdfP07kTTD43sS+59a0yGBpnrG5CcmTIGb85
vsqa53Qe4JIBOB/WbcORbWHQnZx8P77rK7bYecmKEHSD1zKdmA8qCEcIR1tHHwCs4afEPq7Txvvs
TCXsVQlEL0hKzZx3Rqkv67Eub6V6ELqLrWnPUKQJjcR7kiZOFygvr79jir5IhOBKFdeZdN2+08NM
lSE8uxuxOj8920/dWycERzdP/95JJeXrjfnegi/HZ5XTtrwuaXowaymla2CtrdA14NkGFHipOuRE
2IpnQsnmJde19u7vqhMY7oc6jhtxDXvBI3mEpox1EU4TAH3C4RFpP0UvnL3Vis+8Hwmp+dG/CHRT
CPy7zSS4YlQZmnnztIu7ZSYTamXn2lUarKzE7WpOmLwN288f1K1RCdshy9iQK/pppVHG39yDsDZO
gpKIdaXHsyoTXUJhefZCz0//hygAu0BJEY6V4aobN3QJsOg2YK1YF5g2ZfyBb7KU9ZpS9clsqAsl
D8j/8PpX/LaTZJFIKBZ5ho4euqZ4LfK+57GaAqK5AXQSdHafPsAucuGGm/h5j+tCYsCI+7XBs3xQ
g6EDJ1RfIFeNjeCwxtnlZsSxo5sgEz3ERkK5qKSQxndyF5cmMc/FSYSap7HrjROvd3oe5/trImrv
dJLZCQreiSFtUgBpDhklAi8RSr45uBNzJtjQY2giLEa2fDMwyEX+9aFbsW1iyY9YuJTvwU93yVBf
Ennj1mwqOHRfHwpgvnoegJbOluRO9hgNDCisUNZYGbv8ke/wVmI48vsxj77iWSrw8+RKwwPBXYKW
DuAqi6hALYGyB/RYn9NyuxxNKmJYmJUPRd2tAMUlxaP3VjIMK39C80RRmG47zrrn5BTasmJ3HP25
97F5TNuGxanezmA/k1oJXrpbZ/JEV0lIsntUpTXhNupFNLM3imvXyvg+t4Inj6mG/iMtOUVX5zeJ
WCBykKTjL068XfvW4QiSgrKbzLDrn0xXrRYEbXBvWJLg4IKiwRf3iX8QBH4fQO2t9ZB6DD3X2ohv
Tdy30g1J945vh/IjE7Ft8oFwedrTxfxaDwN7T7kCWwneManIvvekOQAVgH0y+coMXOdTzdtskv1C
nKOHqAWb7ICOnNu+a76wk/iNE3DO7jMQeOi0GDLHHQQ1KgvaNODnsOkgFroJpZtNhUTNinop9Xpv
EDdRxQE7CBme6GgMTjoZdjDnRoRdIySX1+tMApK+ridCXNM1jtTMTYI0Nzzef6JnIdEWvEnC7oS3
cbup+ElrSCbq1B6/eR9EN55qOX9urcp7oRjARJDi1q1MTcEgeh9wOXLCmLq1VQUMIgg3bKVuK1mq
QHXK99JMQf1JYRVnsNNMsVWc0u6cNju3AZpLIePJYLNNAKPrLL3MO7yeHdozJISdJtPOkO//Ast/
3kwrUXub9N+JaWuFkBqCiesljIBSGQun/Cqi+BV58POoGbRYThn9m/7pGcgEK/gGNsLU+YuiHNxQ
ZOYWrBhDxXMV/M/4YIcWFQr1+KV21Ot6MjecssOZyuglGoOhnwDbPB8pbejtSuBQU9gkfPjoCswb
oFHU/xMX0WLIpnUgmX1tYV/YNdGsTpYRyZ3CZfbCLD+UFL84o9uT9HxKWHKIo51yqlqhrFNvjhu3
CoPI22NQB3fXR3qjsPAzDorems61hFnBX5kgRMZ1K8ATc51oI7qMk1GwLMyaPym/jNNLS4GO4n+Y
U5HEbSg9ZoUbXp3jq29ECL8zoW7fYSr0jJgvyZtxMm0Z49K6lLYSM6sdQmOWvG1l9d3J90EqzJdZ
JacBOMJP6TTuPTEru/WM9WSpBv1fNAUt0rMOPTgMF15rOSw6gmrHjSALod/k4m2B0tPaNXqRdPvg
JnnJA3+ATlQ9G/+DNss3OQSPhs3+P73vh6Hr2azScl5/DbzlL4TOGnmqi5tgy1m8PWVYgmPtCbXg
lbwt1O+cqwH/H4PhI8pVSsQTofwu6LUOg3p6BBxch33bspxoRqUtpwszXyUetHNqcWiHwhnfdeqa
LTZRNXhhcPDdm0Ty190q4Wp28SNAETQQLwPtubP6vbjfe3tjRYJOcFKzatMX0gdDnK6KKUG0a8bP
7WdRlNs3bRLnqFBNbL8aKcNcXDI1igih8apOsuY6wnAwEZqRwc+d+/46cNCymrrzd/uQUAiOa+tG
QsfRCPPUcMshivXTPYl7yoEqygY0cTGS4Wb2A6ZsOX46MzPxkzUY0seW0ayQpk088SNVCmiDtZ3g
9Mnkz/pfX15P5nYxaOK2gtnOdRk1Vwsr1s3nsb8Boie8YsGPcYcnmQF/BCWU6A9o1i491c3stkAV
UrbE6blpB52KBRza0uFxMEygM1KbZtIqISPGMauC0MsBxBeR0NcVkcYIifdpeQCPiZ/exZtaxIFY
5jrKx/wncXw9HVK/Tfvka5noTsWZpjRA8tpEHYN+NHhAvLJktZgo7IZIO7ru4nT3JVQsOn9f6Gw4
GfCdkQxV9vUcpjBASsFWL7Rmp8X1o3EBVXYt8WdbHdFYBZh7IlLvDiPy5JHIZf1DMw6mek5cKnJy
7GgYq81LIHL5QCrppE0QKPdN9aODupckty5hRgi7aNSm7nlFlXqvnyR342O9NxDNBubPYHO36ohd
wDpV6jecP9SSR2vfT/4vaPdMIlSQ180kJNv9NMzorzObO+fe9I+iyQDuNFKYBRqLjkgQFMN1bWMp
JA9Eb0qlMMUkUOmHUYWEanwqUQ8tpGVf7WXi3/3eVs0W+x4AOK9oWMDX/VYwSFaNEA/joLvz0MPA
+6oT92kgymgOkjDIqWe8R/QgsQG6JHAe7iU3V7/W8A69tud1+wdK39zgrgHRmK/CapVV3ItvSbRk
RI+YLlnGVgJDO2pZzoElDaJRAjjbfNzkK9hg4sJj66h4YajJuvb1jjeC62puCc47n4cOUmV/cxuq
9ujtP8/NAcLjZhL+9EnmW0Qv1f1wV9c11Whqq1RfMNMmtMZ8Zb7S40CfV1918a9guDf9d9anz3fT
WSCUgfuZK8MKPxfVhRJZE60DaI1U3mHo09FF7qU6uljSgGPr2hX8NsyeSC3vNoC9zdtw/qDGTNzl
R6CXT/QgNV/VbyMke4oxuT7lC+hMg4EDCugFa9pKSbqeKevIt5trU6ZQP2VqUCUXI8apskIPOrjQ
VV8KoereLXMgpTZaXFGbgJhiwgqZ4PfJTQujlG/sRA8Vl2JzEwuPDme4PzbIBFs13y+xsd72EtlY
G+MHVSifi7ymGxXYJhZ8WyysW4i/JS5D7R/cNZ27dBIn6eLND5JWIRMS6VZn3loWPmRFzWy4OmZk
odPMIY3F8we/LsIy7VuMxFPpOyef2IUG9+dH6GZ1+Aw1lfh76h9sdrUbS5kjUNX4xgLrVqoQpIFY
XNPt7qt8e89nsDnULvAhr01LHOF14lvz7Yt7JS2i26iHaCZ51+TwkJ/oVacrA3Kl4L1PaLcYD452
PYikqPzzpCHn14Rt9uarZER4vLGluiVbIjr1n6fa3iF7Z/ProjWkYq8PG9QdY5Og4z+ATSNCtTue
gewDIQJ1TuksNyna0K6QpFUB6JHy87m9Xqg3wb2eZqtMURj+uEek/Z4vujHwoJ95r+Bf1bqQaR6i
5uOK8iKLeF4uX9Ko2zczDjMP69Z6xNY8GF/TyCjI7xlEkcvfQ/DpVDUqrtdtlqGCxYrY35gFm2ZJ
U9/8zApWkwCXstc6IOGqwHCyITFEkqVczHUZ6Hagf8wq96xXilcicZrwyw4Olr6KbyvNCpmmqdtt
ig5tfS7XOnz7SEsBytTeqK5xk5VzAFefsxtKrfejcxWI2KRCModQEfKVV+n7MH2qNPogxUePcuhM
iRpDyG1+3RQNBJzqe1hMhWdjbw7tamj+4OI8QV9RUPhrjnBSzQsvsaqzrI8HVmBz06Us5y6GB2bq
vSnJVAtCbNgjps8phqPXoIT76bLmFIxEwfWtZlVCjYQBljsVjoC5loX7eqXDSrqfIP9rR0ztMC21
P6eMvfDBMNO5f8Pjk4w7L7vPsuer+DK++sd24VaDQieXvxm7LiKJrcyo+5JZ5LhhZZbvxgzd/sri
NEoA0kzmCQ3RFe2EPbOqb8WMQKm+OnFe1QdoVTvcowUxb+t3Fg/VlrJjJvdvqNVX1dUUgzHgT13e
R3irPpOKa/8YlNkOk85GG0eI/pjhaxUBiOtYk9H5Gl1WrQMN52DZfioMmLFE71IrDQD3+N60EJeF
Dg+ArsZ0zZC8x0RPXRt5AcUn8nTAxNutDeZNrvAFr/jQU2TiNnNN68laAV2pR6/uqEPf/NlLhEgh
Pei6/wOKvDyscJ31ghQ1DM4iwbyMW8RCJ9hdMyzbN2+d4n2tzvRZZ+tbCXY90XMKbZS6YJ9JrXvF
ax1fj8O43Dy0nYA+ZGsL+DZI4Y8rwR+gq0J5euyJC29ZBm1dgQ56Jpy4Y/89SNsWPqR5ykjSu+ea
OBAvMKdZBKpSrI6pisYV/gN4Y4ENfTV1kAniUGybBWJYMBQXZRX6p7hsz0UckTiZpoan91LjVyv4
PbbgJwJXUwOSNAVALp2XzxTynIhFdWMp/PvhSlRTZ/Vv3uXFcud8iLPiD8tlAx2rRZLyKgMaP/cB
xxWhhmz7UQKA1w7TaFclHzT8qs1j4WXyEdNx3gbOdjsWllmEs8Pa/8nWlLmPcAqkUbbAr4pG1urR
bdKQiOkBmppMQaYeH9LCjrEn5H66rhxJJJ1w+qs1tWhmiKhmyPCbRguKmdtqLa8i45PhXv8Gig0D
B22MH5gTAgM4jQRGk7oarkjmL5j4EHY6y00noN1ahLUV9z8L4jyA475iFriRVpsK2vtpU4P7yJd9
Cvnt960uaPhda9y4i+rl4w/N/XE+w6nCpoY31s9bSajrxP2HC9z6rnKY4AK0vYUs945hBxGoTJS3
W7X/HPsLhCB5H4FdCOMp5rptkIXEpPSMiqxyOds7FgvMrEoH2JdwfPYJqvfsGG4vUxuo6kTL6kKL
cjFRDgPSKLZY8OGKMy8xK0RL7Y1zZ3Nl85ku9vN6L2LYRTCCp36RYylcfgwidZuJUgZ8vzqBfHJi
Vmkhu3aBuzUj597VICo+/G7F3O91AvPRJtJqoPF/+C2FMTwqK8pr2yJueWEVT10e2Xzg0On3m9K2
Fzk9rmOpW00SuMot60OO9iYf7RZCBukVNwS1ujoPAnPqj6FvNQ+QSQh+HdObR2tXIh7ZHpCRpf5N
hYP6YdxZPpxEOEzHWrSEZ0gcCjvbfcagXWrJyrv60wCwSbvVvXj7NF84tuGwSVizYMRxeStdSN0u
rRL/ryQ8PFkFh06WtbTQfKwcDKp/vjtg3p3b2FNkvF4fadDumq2uHM4YAV7IgTbT4cMJPCL3wxbi
60q9r7zngrCjqkLSpKOKiphyiO++nYiAIDyMStC1tlGmiJPAiAhcV1ExhjINOydvq2BqDAFIAKVD
d++d+68/0tEU8VBmiebopYP6CFGYGBC1ZXJaSI8stchZGRyxAOidaURUP0mK1BMSczrUgx2leHw4
NsWs+NZeG01eDAUTNnY23ChgnjE2eIeG8diyS3AyCe1+8D8WykVeWU/tuXynEiYCxds+gPhVgbpV
Y0IOBdesdC3t5bDQnOfFtBlgPIz+z7tKLxR7oCrBZtUhpeQXQcfb7UoDjj0xTvMRr/IW4qkvGuYQ
/UfUvZwOuiqK8woP3y4LfMSR4XLLnqu7Yn0VqwDqyq5ckvoYi5wHDJTAoZF5tvgq/yeozvOA73Pt
wkDUfiNH3hKrdmRjNKHYIYrZr+Wlgs0wECyNv3Zk9NFfdlrmbOsgKTcKZnV3LPO4Vv9UXDihhhrT
+T4nApaQuVzPpCbaYcSwCEz0YyHy3U8jxUBmxz1hSPrVcJelFTIsZ71cXV37hOtw1qIa5Tvmb9eQ
DsfBOlet8XRRkukYqzOvTPTAaKON5AyNm13FeLf75exUHl/iA6IarjmthXDkPnulIQCfzaO9Z3OA
TH8j5/pibb/N2eO6lEgZtmInxdKiv9KkVuZE9CM0c9FCmhdSSoZJteqT+xp5SbDf9lB+4o/zx7b7
Ro1WqtKxdy8R1Vt8VJ9wtDzkacu/uMGlZ65FTGZtbA6jccWRrsopaazrbzDtdzzyJvfjuhjh2Ai2
5kZWuTJSddvATzOLoG9770qvIZaigJkzq2TzqMdbOTjqfI8fz3YiqLdrq4kaMI5hwa5QmkYXvkOl
aW5bl6uJByaTO097nw2ojyF2d5FvEd8WGYC4PKgewkLVOMZGJVOb/rA8z7idUvI1mr3k3j+Koy/j
zm0jHQxLOkZGA+TGbv6gxUSaIn04h/U26EyI9w4cjNegOCt3U04kxEGuGmjdP9RH1JxpNBXFlIJh
fxdFlpiWWTrS3/QZKql0/84ItKs7gcf3d/LXA31yq/5Nkz+oTdckjF3qdqJWFktMCmIo02VoRBeg
3wUGJuNifCtLOTv+xB8mUasmq0sCWI5fZmWW3DOvbs31WNZol0kF7BzqBaqYXtSJ+DAEYZGbOEw9
SrxwwrPv88E+rNhLxFX3kYuB28T6pFvEJPt17kzfucUBPNm934J/124JpOT5R+CEVysBIk4HBCad
RI12M0BSsbsBj8x1C1oziqgU6WatJUqll/bwZZ3iW5gfHRiBPSEfInUz09OGecjcAqUc4/jtLTrN
nNQflt+ntMsWvhbNf0QfD1OW5Vp9+geKhzQbdr3BEaDYkKKXm+97GylLg94L/J9VCYv+j7JbDkgU
Nl0ETw8sRp7xLP/h3FgMyKQbc7wFcIco3S6f9VtpS+pQZ/0OBOff7g+X/Bj4Qvw9ZghJctAe3EQc
CSUfq+zfiDc3oCchQb1BDKfp9gDQDhgvsh6qP9gs7O3mJXl3809D6p6aCvdbbtCe7ibpdwT64+1d
z8eILJayYRjDfmJjUtOgrCfDnj/E6KnObPKLQ6u6zDzCFxuMwlrwABPTkpnJy8OFU93xoB6KbQk2
5Ejz/goiIw6gIo3B0lZhzmdf2aOwFbX4c6e0361TPhDKNmj9OkfHx5jInDqjERWaYM8Lc95WG6AG
Uue2srQt5U6yWd3TH2Ub6DDW1IvlqJKXf/dYvCq2GB/JN4A+O558xyeo3i8lf8eE+XyK9Pf71kxe
ZDMnOUEEnqh1xZ4VaPbuy8YWtiEV2EEn2J5UhK/H+BvgeZYYL7nYziN+CYq3yHk96CYp7rqQEAzq
b8P4rzmYHNX0GebIPIboz/fNlY7PFeHXsievjN0HAGrV7RzNj4WB7y7CvspE3MBNfPO8sZfa3F2V
PJ+kg8ytHCCXg97KlvAwwkfcmz49cKjBF2Q6DKxowDOstD7T6H+ixSTUCWfu9EqQUesiAtn6poWU
9LDjvDfPW77PmxwQcXIjSo0f0jeziP3dRSkthbo8x3+RO9qj1l1T3fDXT3w/vFvUT/gm7yR7GCXq
gwxo5toHSI4CHYOMZBIVUS651ZHIK7GXdVSEyOtc4NaCbiMW0uNjNsksznMKzYUVy6blFvZ+OjPo
v9jOeGqpfM4pzFYVCvrwyLxJIqw8mkTpdDfX58//67KI8Rj7vodIYB8S5hxx62lCHKLm4C6CG5Lg
jrI1tGusje/BwK7nd0MZ+Zcy6eK7z2X7WaEjsENQXvcTzqOoavxAnm3TAv0F+5vpY+CKCAMbfQpN
uGu52RjjUns7geiu3jyuGXRvBnYBC6sFFewccCoQ+pnPH5MrpTG1gmWZG50K1pBoX8yOHnYPdmHy
htzaUNCbc2kQ8XTS80zI8MyaLNHGxmn2gR3f9vyHgx5Mzb52xjmrlKoE307ZcNNSNKHsnw6ZJ/aS
HMa8X9DJ/feVrSgUXI0g+GCd89kiFMBCxqir2oFCzoplgPOMIN39Wa4dWBVy9b7obVet0njglSAy
77B36aYJZo8Ps/vlRRPrVbegMlRFzAwOH+sbfeIrel1VGNMnSarOT0WRSwwBJxlf00RmZ/zVhvRf
PlQ3Leunia6T2suv3gb6ehI6NecJ4rM2vmHAriNuyMmu+EDF2ge7MMPWPZYkxVA3lz0HOtTFyOWl
gHgnpz8Mwdy5VWc1W32M+tnaVxAwFbzpCLgxWGCN3te+REXZZbUtccWmA1U/6YSwUZWpaH1XXPY0
NmwXWbrV7d8tXW+uvW3rJ9u9soTyqYq3i9tDlaUERVGQxcTPkDH6QZ0/x3W4dhDXefK13540JIwS
GM5rMsHRX7V+f+Chb0TeSMJl6RJntoXTFsnkugOJYf0smO6TpD+oE6A3Grozqf0T0klbbaidZPm7
6MpUrm35csg5IBplhQGZg6OdLI+cfpP1DhQvUF08U+x5iIFW9PKFyZw/tDS8l1geNEL2L7sBwyGZ
dIp3m5e40CYo4AXl9rDWuJ7NYY9m/cTbsK2Oa5HWPBsODqlib2CEwbyfrfqZoXxANdyjJMhYlWN6
ZfmJzMB+ryivgqunKUUB01CS5ztKVxOe6oQSw81o509Y/nIt75Yb94GdQK0EDypaybdg8feqzqWh
7j3OM3nSrK1OgMzafiUWshbotPGLvbIYL/CTrnGiPMJvyPCUXhCaIrdPHwIy5lxyaGAHvb8dLtGf
R2UO3mPT6+7LyVOUb1g4/GFIs+p47mgber4dFsMWtLV6TuiLTsRsKGFqdIxaN4m+zaEy/Vp98i0f
fpcBuOzd5wiYkzbJEh7VTA95iDlNc8LdsfG49R3sT6Xml1bUuG6Xbc4Ixy2mKF/pPY6aE/iNNPBi
+KcXSKJ2z1bS2eYoMhm+8UVvfnU/h2NDsTOxQ3LPzvSKMRnBN/lzdYrBY5RThwpKUykKJ88BLG2F
/A5gb6+M4mqjFR2pQ4n+9k2GiloR2Qx09qTOT2kjw/ZanIJ1QEUPN5oYdz4E9/mB0Zkyrie14q6o
Gfai/dK8te6r7t5ZJ8YoF8j3LM0kP0wXifOJ09onlgQMtgCctWL5UXngeo+m0av2aKavExkleVgr
GnwTknH//ei5VSKszyuW6YczFUaCoTuB4F0wxey15ofmxjZnDU6Fuo1jmDcTo7bZfX0FoNbXOf+8
mGTB71rkQFYmwahHopPetM/fniODOTlHeqMA+xcrxYxoukTAcKMnE3HA0CCI50PI7yrXzpWrXLdY
rx40ZN3wlmZLVczg5/B1N3I3lxsX8ZYAnK0Qhn7pJbJWunVPOJfYVjdoDdAle0k+eONJD+PkcZ06
D/IbcUdY/GGkWYffPd4tvs2ePNL5ZAn6FoUPUm4QryIy925TsXGGial+ejrcIUspgkN6EsCIBwYW
v2N2qiC56mfdaDoSCNewQVAZL7VE74E61oyZfRXK9MGvbC3L5AJGRfZwlxmnqe12X9D/0x2if1OP
ZsGPsTx2m5XNuyCv/0GR4Nn1uhTcKVNLEqKVpCpSzeoewqTCXM1lHpJDkrE7udyBdR1IVvrUe7OT
sBL34H1+ZYQ0h1Vjk8WCj2PzwKAJCtu2dNrVJezWcBl3ZGRPzoC4c9xBKViZ9TeqbUdUdFfpzHrh
WzMmUqQESm+1wAEHwh/yM6wRbU+c/qBN37B2hnDbdO57+YOOCZ/dfgH4NbwIUWLc0hNUPtSaNM1Y
9ufW0SkPFZ2h4S/Vh48uhy9kIoQmqbSE53I4UDBr4tdWMCYtvR75WF0frZXuVa4KVWIcB/RUBhIR
+OU6nBAmrSq/Fkj/Cb7qu6Fs5Am47obu/r+xsRLuZrDLjyskyetP2d9eUgQTiNH9ZjeyAt3tgdFq
+I84y5TzejxiVob54uUqGZaaZsWXE+pGxavMUxEkAoFLHreOH7v9yk1pl5h0q2EsFwgxau/SCTqW
r7HiqRxwL6wflAiZPXEcyalZ2ru6zRLjCee/JtneBmJHjIiDOrWJoUZoxaKCFdac7WroD/uOvE3g
38E6oXVvmakuqyYVJOkR8mTGW4XINg+DW23vouVDRhFlcc4nYsa+JwOUTqo+tSN9ueHrWC9oXKac
EWpv/A7SxHOmTsGwQlpxhMmtNnlXcuESmRCPEy3AFTd6i/6R6EJWcbdMVcZBOMe5PhVhfYrFsHCh
/W/h/o5kKqPeUljayMTuTicH/3APyQc0SuD44L8H7Xbr+S/e1SHmH5s50zLuECyH56Z9DCi5QTEH
f9NJ4b5HVIgMF/I1Kc6sOkt0tq7ytjE55Ml5Er9fPntNiRFzx496YZMYIJJdeXfmg2NkMBrqgRwj
7U1axgIWuDIeoM0yoC9XYTS3MEXsSC0RU+yolRSztHeFSjVdMn7qf+iDcBHdm2Rq9Zk17R6QDGT3
OMSAsyx/QcfuaSKm0p/Syr9jqqtVZPtsHiR3TLkT2f5RQ8v/ivkeD6385lpXv9QT/k/vapcCStI5
y+jVGzjhwpbnZ2o6sp8fnk/cYcsJrmpKZbN7ojzAXu6ROaA0c//TPcCEHFlgiKWEmDuERyRlANxN
MJ7T9veDY68sSFkQneqJqRxl0AKbgY4WBCKlxbxzkMNBu4HeQqfqJy7qzju6GcijUYWOMSLdv3SK
t1b2klyMydOIdIVSOrQwp7C02G7K0cVrj0NsWGOMLD7+3Xy+/8Gc7Lc72h5AwX3JJQmTXD4rozlr
DbIyNUMA687fM5sssFgEma1HNyPNLknbHGTAmZRWlAkCfNDMdP8SAASZJ4bpMMGChMWpCYyS5Xfc
t3WyU/mueuyMK/wJyp0sI0DU2qOPIcO/R7YWLOv6u2PvpveyAy2pTDcAjCzZZ9dyGNM9FeLq6aKT
/2ziG/Qj4YjTC9YO2/4Ggi3UGQqyO1py3OvokMyMvRg2X7BFnw60SKSJts7ADMJ6pf6N2fw9jk8D
HZ0YwPy0lxzM7Mp7lzugaR5cA+uLy0c+J+lKxhI+omK62k3MuGuSqLe68T0s5NvFhO8jZ4rTog7O
PSPLWIYahBtZ+XnV+CBCPcwlxALOP3NVNm6DYzOtXKzeTlJGdupjyofIlO4IdjqxuCADMshhnVLh
ldTCi9gnKBNldPOHGBcJsI0+3K/9VbHdYq3BROJ2xdHHGsm4IiIjFnTSEocZPchnWxZQ9Hui7pE8
ZOBlA1eEZp8qzT1jV+eozafayD8vrWE5TZm5FJKXbiOFqDfOxQWTv9R50JL/1oFEhCU3saCYD0WP
tu4vuwguExnslJAdnC+MDYJUP+cLR67jkrSInXEDj4Y9jcpkTglCTaljqmvy7rn35K7INpSRnwc9
pV7C1d1xLPbWoFPqYNv9MQLY+VvbmzegEdxS73Y7H4//B96YzFMuIIpxsPpQG0zoyrLpbBOLNbE7
9swUIQ1Pv+Z/ruGoxEnxso/dT73Gk06L1E7bDhZlhoXZ7WWPhq1mnsCjCygRDcnJQV0JlmHlSUhk
R54XWXcMYZcdRW+N/PMyaGI69oNtGcT8JrlpQiv+w6DrYA04EjzPSYNoKnx1nfzZr8K13ZWAb02r
eyLiJdd+ki54AN3wzLJ9tNNVih6V75SG8zmKaaoDgszf3U5PRD0a7EbeJdWD2LZyxDs0Gt6DPHzS
eBFnQficsVK7kH+P1eGipG5QZ/SmqHnIrcL9Uj4HV+SJd5mskjU97ZoxGSYLd3ykpAufNMqS0cGh
D358rbaNf0oiwFs8lG5BEgKm5UaojDDujxKsaQG0vJS5SgELtxg8yl8FuP42hz1uoe+yw/S4ynpm
MSQnxBcPyS0T201yL83pukYq9FeTqSz2uA8XDzfevc16J70QMoRFDTo0NxDL5UtcPs2IwYJna+EC
t5nSBr5MGPZQOvFTyMZItfVK1+cez3BaZiHZbr9Hfs4/as5iqXfMkFVp42FK4+RZ8aQFXneYW9oM
ayTDVd7tv3lYLgsI+mIDevT3JBZrr8EO165E4zKl/s/sx0MZtRtNDlW80StS7J1cdzdN9zAZuV5L
fLl5hGLuFhffH6OH0jN/zulcr5zl+9e3HZTxnSHlereezvOyK7xzHl8t4MZUxDa4lgxNoAGqXROM
84IEaBeYCPytwZzfj4gIMarBdXrt6+jpap+OLB9Bjun8CCbKkpXMp7K1fMoppECzMF0XKhorn9Cl
lAauNsXK+TigLUnYN0pfdYefybVFS3wBb32EI6eFwsKAF3HmN8er7yyq5bqnqC5Sk3/z0Ybdp2OH
bNg8rlEcFhLpG/teHJgE7P8Iv858bQ0wV5mILYQyYbgpYF9knAy/p7TWQOBhA359IFJPVGTNIV4U
tAQH73W66ovYzSkemMY5NKpPJHAawgCFOHdjgM4WwaMWwje0paXsI1d97Et7yLeTKJSTZdXvJjo3
nAdTFiDQzc7Ea49SNU2eIamOqv2zzoYEgEguLIcxiaJPSV49r4/JzPNZd4t0us1rRkf9838aHYpP
0CHaXtpjmOnhD8zpE5D1cR0rxmdHQWrDqBzadmUeTw716pdsgaK4sIgE1wuFS5XZtXpKZsFJjDbv
B2T72i9JLQMUShWvW8BGxe30/Y9GFHQJNfU2Mg0JcilcYSEI/U4QPKLOghkBQPFCVIiiEJzjjJQ0
sxB1ZBiblFhLOkfF+zbCIwfZBKIM61zHX/w+It5H0BSax9r5cJPNHBExTT1Ai2/Rsw6MTnhd2X1r
5J9A7BU7Rrf3QVLJo29HVHRUMTcDwUdIJiqBEVv7pQu1sWmY4EfI5CKJrjcWWBeaUY6IeHTWAb9A
zADuv3+B0skD+f8rP2l1rHSOXo62cb+2bIvdlG2MPyC35edQZvigxo2JNm3dkjg59boOSxPenrMU
W+C64iNz8F3ZdrFI2nmJ7atUtfIoSIZgfXTey9eTdbXDI1B/eU1HlxCFzcoMPaZQSUDYj4SrnfD+
U8VANFXiVdwg1ywLTL3k0ZVek4bB30eu8O8hyhW+p6osohxMxuqSbdNjrwFzyWOOZRI/P6DZpO+5
P2KEHK7Jl09yNoKMU43j+upiN+qOWm2ew2mZHKhVBeU9pFkEvCZo3okpA5MMMVzJ0hduaq4z9RAq
kEuucyOV6+tPBsd/rl3TqynNdxhv2p5qOOqJX80VktUfTMZNt5Tl2ddfRXvtXOGPHg1yU79TERSr
5KJeAw4nYL1kyoxH/sMtFEqyzDvXKhNHd4hPRt+ShwqFmhrWI4/8EUIvTRRS/gBM0YoB67IMRZuS
N7OD33CsPRwIfqBcgWxaAF2vDQKgPHKLYGLsmBseOdQC0PZT46yhYInGuClLHyFfgh70o+YQxxzA
bEbI7PyOGsRBvt9SR99cBzeFvDhxwwqEv1h2yyGNJbprp6B7+Vd8TYUW9Z2Th3zo9iAzksw7Fds4
SfLWBLxro56rL7PBHI+2mfKzjLykA8lItuZBoOmlgH1uZtZ/IplMXoYEa37ohaxHt0Sc+4dGPSEz
NkyXPv1Rr3DPn7GBGVMqAyq4wuoWVaWn5JegOVaewKj8Kcguq8b+9tKj3dLLFZPTL1RaOAM8AE5a
XtuIsgrb2pO4ZUk20VuFjST0nD6toi+NiYnsnC3gg0z0meHomogsJMAjBCszXuxe720+oHkKuLAE
iJVp0VXWFTNB6WgBWrgHOhAlYBt7e56QVAq/ImWcA+T0EMvQHO2QSMqsCMZ8QgS8+5PTX1J1ZkLd
4gdJKD7/5LqblwQB/TPVCYrd27wZNlYaE63J6IuYj2OCGHOoM+kYHbX8jxqTE9gu8aOfQSzDYnT4
9c/vaxuf67uXEuPG10XcLinvkcaJcc5lBr77UkkdQH1cx8WKcuaFST0Jo8f7MyK/4ULJswcxJFm4
ae8hS8p89KBbb7TaHN8EYdZZHxsFwCiNhOcSpq88NVoJER+shgrqbzIQUNiO8Obuw2ym+E2vTk/t
47PO4xo38C399zVtW4enbHhVJ96XDhbBWPOmFSSfkp8wgvajnk9NmISD1yL9v05v+dR6IOY2e5bh
2IroHlK9FKke5SC+gbqR+9bL0Kj/PuHimVWBjozjAdaih3PUPAAkSs7deAlAjBTcD1bpigprLwER
CC0cYc5CNkPEGW+9E+IuCJuYcNpo5tpbpnzSq8jse3kEPdxUeZvlzUGLkcPXoYZ7mgBRml0XqlMw
LyxjhYVIDyWtYZtXgPUZQcdNnM6Rpf3dZz2rI1iCKSejG6Q/onZ9lorQ2l1H/ATMoy/z7GRFWspj
daURZkxBY6J8fCmZgULbOb+Zi3PxH6yuV65PqQpR4arhM58PLHvpnyOPxzkvHz8r744JwRMuSgjN
tNTairCRAiigepmKVoA8uNqQb1GwD3T458U+TmYye+UUywcc8TWKkr6f4Yg5bpgWxaeBO3ypIcac
Yed5frkHCy8ye1opqYQCjPFzcHa2sIjB7js0dN/fwMXrchvWnXxxUNMRwQ0ZP9gA0OMob7TX5gqK
fxnRAMavVjqzMCYn5fCpYpmjE5rG1GvxQ7OjRUEIIVSmrGQ9Lavzqe0zYyIFlwMEuVNu4gHRrYur
7GoUzDnyHQFv7IOmQ/ZU7aEVoh08QNDwCApFbkUD6u3IVy2EHMmym+nHjIMVbddF9vdcVTe/zKAB
WvLeU9pxUuXRJnuh6iXqOL++eHrHAJ5c8+3xD3tUq/wqeTM15Abf9Bgk1nBc4x7gZJwr693pe+pO
bpP6S7byIkiq2ZBVB30jdUZ1pR9ahM7jI/SNJahmxRALiXPyYI1PKiQFxr7U7w1gdA4rPZ6L0kzl
3S6giX03v4GUZSEThEgtMjanIEyDykJUg0dhYHA6jTcm3/qYaMvupInI86VuBG0kMOB9EVFkjBU4
dFl6J8oMQsonb3DHTNRfH1nbM5didgH0jVN3i3m3rFfv83wtcxarOtM4LJ1PP/L1NLgpxScj/NIF
ySnLBQthGyBN5ksNIncVLBA8OAEQXo8rE7wqmfcoMEKFnQ4mTB/gg4A6WbBR3aU+Im8X/yOvmOim
9lhG90YwlWIyCQHInecO0clC5+bP+cB/PMuKtizKzbJLzgGw9iYWvI1C6VCcrvIG6XtroAFPhs0b
O+OTlmd2WB4ufgS2MAfkR4BkhFlroM2gyDWBbRzoM9pV8Bvh7q5Vj5VT2+oKANPjYIxlMffRcs7h
EnSZVyiup0TCd9zD1xJip0KyedlUpAJzTiA7Xp18jozHo3KUd7inteibL2HHaAWE9+5SrBdsmOgt
LbKP1XwU7t1I8FS2OZhJdlqASjMuuNEb857zhX4Ex49ffRF1kDZOeXVFY1ZFtzXWZvAxE+VfLYFz
kOq5o1pFqusCQxFBhSpPsOkrdQMbuVASzFLFCrkbWbHUduSw+gURXs0u05JGpuCH+67heNWZ17s6
euGaN8W/zOx6cCy7PjbARzEvozLQSOztz9psbtiIPUSesrXGK7gXk9BeB7LQEL+ylDfgaR/UxVuB
Jp/NlbBF5faYexcZ9qxhSBteXAkoBmsAANWu1p0IxRUHrHa4l8dGCU27iSqqGsqGocn1POOJ+KJd
pPYN388VAYH1NId6y4w50Z7cB4HQFFxEak95ARKZ+1F4PISuhiNjBKybRIkNxldGMBsc7z3B2AkX
hKJPdGFunKCmtWCblxsQADXyqvXob4H4XUYw+JqL0O5muoyxILLbDjs/Y/vNfaPeL9cdfOr2SKat
PtTmnxfhgCZXUQjR8gu+hGW8fSZ0hDwtndoG1vLtzNP5qvUR6uDdEUTz8gdn+pwF6jzT/MhzgZgE
XxGjkDj+CfU98ZWgNbtBknuf2TzTNsgg3yt8CbEFRR/UsNzrh+EgLS7n0zeXBXwQAieyTjMYxh2w
KiblRp+LhLZYeweBW+WavkTK+YVKzcuWehI1uedE0LGeIMkb28XJ7KGRxckyjObWKSP8rxbB5/0I
6Woe3JQOnogL1jzAPrkecBkurrRMI6F05jg4akLM4b6uuMAQpJczzd2mPJ2W8SBkElDGEcAtOoRH
g1ycvAdesnFGxSgi34ygMlbMCBGDzBePISIgpcP83ZRLCYXs3Xy4m0wQgWLQ/9BlsvIYee8XnJTZ
GVWRB/oWxvC9gIqeqw6C55l73q1lYc4MYo7p3unLPBG5TOqYlXVkBtsNAjORJ5Y2yngBF0PBZz2p
5x6mvDjWPCyOd8pVTQh+ULs/wCqSucIm+jB/1D8LY+2j3KC5K5ONPIlJzRj63IqanGCbwYl6vhr9
/Y91iAz8WS6YeHOqMtx9mICkvHVphPpRdH6cU2IAFOmxgpjEINU7AYLrUS4SXrQTepAkn9HsWGHN
241rDrk8sr3n8sgHVBSbw6LsMaacBHtTNCA4txzAFZbjWh0kECl7ifwF/cYOcf/e4iwAAzJpS1eh
zfjIMRPT9VlScUk1Mq2fgCPYfAWmfCPjnayCUDUUCwDpwsPHhQKO/hpr02oycNgeTlgqfjVb0jQQ
fyrCazl2ybSU32hZCreSeWJ72tHkfnSgZqtX6u88QJ7IvfwP0AeEn2i0P2QszeGpJoBysIfsx75Y
RA16L1MMBsgYVILu3d3fkpwxgA7uj0crMWEnoX9YM9JZ9wWNqAgH4k7FSE1XiWKIOTKd60TnlsZk
rvswPbv9+lU4wrqTR0fgooxwlGZ3n2oLyN3d9lilu8bzS5hrbjfxjLQqnM0XJ52ycPcg+N2M92E3
o0OCjXm0goXyEzkLig3dqDC+eG92aOFErly0U7ATLT9acnBd8RnSH5fM0iv9vRqWgq2dyNivzeye
nlEml1x9m7+vaD5v44/fGxW4CKCd7P1FICYGIlRWe2SwT426RiABv9TcA+Sl1gkUISW13sKt4Amt
XaG2532bWFjaMoSHCfN7786VjwCkHs0nALQGakVVgpY4K2e/EaKpYa2eLAOqEPyQep+Ev03j/uCp
OcOsQq5htvYhct5hMWd/YgC8BMiQ20ANkeXEcuyl5YS2ppL7gFtzWR4jo1uHSM6+Sl7jq5jzmyuR
b/4wmcZxRYHVk5QeEL+8t1JqvVvh1COF1To9A0+myYjP5R19htELmQ467H7DfaQmVEr+BnHkqCZF
iaM6w0l0kXJ2lULKIO4bTMbO/jXhddXxflbcJM2h1IERetLpSM/yedL5zTWYl1OjpIPd+1ACeJhU
El/67CfgoHA3NaJLSOOjit+/Ve89i32xbesOnnfwaelW90Xl5vIeWXeYL2LITOclrj//7i140pBa
EiIO9xALJjpQlCVHopgfxeqYVfsNL3Kc26WenEvYaC9GGfmE4Z3z26Sxf/R+tQoE5txu01MYQUzh
vW8jakYhZM3RYH7xQDjJLvhta7475CpMCWIULGhnbs5ZIq7GBzQArVY20LCqZwjSpmUyQLjcETbT
+0+zW6/fNKodqgNicxN9PFizhC1eXEq6cj7iSPj6Uce9WSl4L9hgDcCWmJBf+GypfpOPyrYv+NDQ
XEBV2qqW58fh0kEAc+fZy1vFRKqLbxv9CNJlc1yYjkEGYR++7uF935z89fC8Qz4DM3O6k/K/sQOQ
FLfh3NEJDLHmrumg9MBUkcSN4zuEyjhnsf7Cv0MJSUivCEXKB68Hungble1z928EBXXi+A69yHd0
7umGb1XPUMXQDqITWB7wNvrc29ZbqmvgQk+AVat87WFju9pEXDBVGA50vhAjrfYJY1sQzXC7Nn4W
3jy+hUgihw6uaK9fF+WfDwWkHASbNWFO42EMkSra4G6FXoS0wIz1kfSOrUWZc3zLxaTxjXUR5cn6
e0vFLSh5B/9yXVtMSaF5Z65AbGzMO0Is72mCYxzfNqyotWekJKbv7G0n8BKKKPcJ3aK746R+HyCW
6pnjplNvL2VOofXAgu378i6U3FA1ayEjSrY8fga2TFdkZXbAvHbZ+ArmeOVSQbyMGX9fIIcPdi7I
J3HtLMOvbC9RjSUYiR108cGhhNW7UP7UqtpdprZ1jMogJo6PjY1N7CBqn/9TqH55+jn8Ufk7mo6l
5LNPLvYkJygR+zEQrFV0DgSr1C4AGPPBnO8D0Ooqo1Cjyq8BK4luRSezNs4sHU4CXkcAZWLipfm5
eN26OC8pDu8/xzwc/8lFmcVYW5tUBHkbXKk7F7eT+/oBwK6lJ1sxu9avCq9cbwCry091Ltevm2mI
pZ80TLH660jUyasyr8Aiu6oMuQMraveYx0NN1y9UmNXYiw2ug6LTVQCZ7xKtHJ2u28t4lRVvBIyf
R8D9JqJs1oBaqLNbP8HBZvyKDSC7IRfggxqOPlj8jS+XOTeZ0FIi6Suf8uJDDGYWp7d304LZmcr6
QvysbodgjqkqYoqsvCSXnHOV7Y66gyShiCrpKpeG59vepQnEAWUPGQsdlaZRmUo6SGOJ1A59XmOh
ZJpVMHqTd8PB7Fn7spHNGSEqc3KCHOwlJjNuwJw1Ofb3pDaV+kps2t1NjRtoZJ4n8iaD6rpp1AqI
axOZr5qMJZLgnxt7mphU3iRcSrY91aKSmccMgewNPznVRa254YCZNDJx8PDlwFRMF5yt2CJgkOlH
o23A/nIxrvi9xHdoVQWGawkszLABB+eEdrTWA4X1fsCc+gCcdll2n574838zcTKlL5VxDsOAYEZx
jON7TVGdjAkOv6ZdugB7T5Goc8pkBcIQJgPBT/7OYzAAU0UxVVTa05SK3REK8hzDh0YFl9N/SwiH
rL9c4UeHHW2Fli23F5ys1TnwH2jinfmfYlCRMq4q4AaMMEgVpSD64HVXybZwNQATCFpGclY/eizQ
0R6yZAiseaRabjs5HeJ6tK41TSk9iJHts+vTaFISTxcX8g+Fm/fpLQBJ939FS1Hugfk2gD48w0Jj
Z2g2+e0tm2mD/0oNCB4A0Nz7tdkb5mSNaSn/83DQ22chRxLe0p5VKyviv+k96ZViTVLidNuQ7dJf
YjYLpp2VaqIw2WQAtu83iicdOb/iFQPE8gsrDehL6VdWALhrBA46Dc30nzFDWzv3HNKzZT3c6bOj
3hqu5hPiUN8gDTzkHmZx4aiT0jub2GgLN3MEZQzg3rxrcv9dHscN/DkzMkM9ck+ZlF5JdF6bRFgn
TTMssPeDSaECtfOyS4ba/HkU+ykmhoS2CL0JLqaiQEuArf2XFLqLXY8rFMIMK2b29f80zIHxgBd8
XybwnSjLFWk55x1IUqXDYdqZ+CoY9QbV/o9a+nivazmGkvK6QwhLb7hEn5a9SoyOx0Y/I4Ts6qko
faU2c9+foSgaiETSmNcFW1pfOKFhOYyVB4IBajfK0JPyWRuq3iT3RuoT3uR3LAcHnUG8unoMim7Q
Csx+8Cdy+uMg+H5GLVOk4a0aFcNSpzwiVMUaE/CW86jNFs2UNSvmxa8WyNSJqIBihdFueI4IjgXM
Dv7fIJB+75mPMnPafLAHsNO5aNZX3kAj9f9PSyBd9I2spbztySez5LPbSFuw9bERZlenNr2Al6Bc
EU366CljBAZGYDA00Ohzpv4olZg1I/iSgipypT/goQLKrKh8l5QCc3U0UePTs9Ak8qEqN2BuUncR
IsBT+oujr80Lqz7iSWkNRxlWtrW3RSdFmt0H8v+MxmKVoRSBt6/VVERlOhTlpL15FFnMXqdXigiw
8QEmQdj34M9B4D5NYEW8SsV9JukBHyo4Um1jnZfxjt0WGXA9LHPZ+IxQL5p/3ogou/10hEMPdib1
jFMPrqIdvVOpHiKgqzNWN7pKpVF9RWqFiAT/FTNB3D/Mgom5nEod8RQkztNYaGROQUSg0g0M+QX/
m10S5BcXSWHd0eli/9f/1iu27/Bv/UDU+B9r3ElnU7CGZOwKaJb22KzckhL+iKiHLTW3dBtT4+Wc
nDN/FGDf3rX/50HqssDNtSRe/3BwJWSTNMtd0Pexl+iqFeptSp9wo5itufu7+0nlGUbu75w/OIPm
/hbdiZWDAMG0a8RKFWzhtPhWDj520TEj5Izc9J/k9ECv4JM7n1UCQfNWDzTSbvh0cOQ2ZKWo+SH3
x8utMLvcFD5oKY6bSqYC0r14XKZwqKsDZ5ux2f4PXTXeXwsA0r2LVq7evm3/kEk5ZDhm4lQq+MRB
4t7XYq5TMgQm5vZjQevAGNY64KFIblQRBEKoXUtny+0w+O3sYLqVfDKo92zEbTGBuSBZIHSDYjvV
gGAPtR6wdjae+u/QysCkLmt0HS7cDpqtGTHdXoUA7HB51giLemaOxqgaTcO3UByHp9h9RiXbYiRD
PRWE7tdqhwlu7SSLmP8bANWlUkM8XfKW+/yNomDSUsJzde2YutAE+1GhSsxu7OxK84N6yZSSGPUO
Yemf8pkdGdUnw2dUVUJ452yuMfBDQNiNr8nwpyDsdQW+B+AgnSPFw4QEA92iOSp/+Qu9TxCWOJiW
oAanbRIOoHLKJqaNzWlorPJftRKWklocZSpcBaBLtvXSPChSYPXdrHb4b7mDUSmdYMvpcCIuhS8K
B2kBVgynFQZRLjlXEMj0NkMWINWIveZtvl5Vwkpa5EWF+tF7jXVbsTRfdBzNQqSRFzxdu//F+ZXN
nML48LNbNah5J5iqojCjohsD77RMaJo19vd5HEnvkk1WlWiIF6yk+IJFv8IMeRVVRwdA7pDI03+i
uGqkfQn8NVPGXnq7GJJD0dmUoVS5wwUQ4B6mFjuh25QOQ88sdoxpaQMMZPfTevNWEQIG9guUKxyo
ifBP4e7nv5fp1HNgK7GH9TfbOL33PudFEKkaVPqhuL89D8Fllaz8YcL1j1tkSQOR0WP53jxAWUXK
wiavVA81HhP4tqRqH4mIMHT1eyXo2HS8R6qcit4PqMdXwfnRc9taZBd9DEdRxoHX57MGqvsOt3kp
2aSEuhwENXZGw0oX2a8OmTKrdlPKMktNfb42XFfoKB4qTTDCqRh7rgVUnJLNQQlFQUheABlR219n
S7AIRaDWbUahgYiO7PAA+drslnAVJzSh3wsA9K+fF2wPNMUtdJNe120YnDzw3Tlllx51bYyE/sHP
Sb9GfwHBa3n+d4vwXawnvbGPSRZdD6SA69cqKdHhnpxrwfcKkHKFA++quZ8PJo/RVl2BEIFSE1Xz
2VN9lW2vya6Ukko3KgJuXHoHBq7k6vVfDJ024VDowPZBqiqv4IOchpGatlLXsrpL1DC8uV0wsfGI
GOIGSaJz79DW8GOiEFM9QBJPdHjMEGvWKEKSNyXa+b/ADMDQav+N2nV2FxE0GmSTA2DeKZleaodY
7839BsHcc2hQ0G8CHmwUFICZL3lBNgWitCo1YkalchFGqnvxiwIkerrvJkCTU6yPbydiS0oixFwT
Ywu7GWwGD/vECSrRBuy4po5wVDRhVTtl1N5JjIaRiNfYVxcn8jLD+4a5J9Cq5SodzhSxhzu0Jwpo
XtfVnUGCaXlVlR+tp1fYZqTDgsv0dBdGw6GF/PQ7MkQTX3mw0uZWfbSF4pGAI6bljFLF/o98RNbf
DysgVg/cNh4gHMlyg1td445Ie1x2FEpWfXvkzgJ1yHipedem2S/O4zZ4zgeS2oLxDKjmVEcF4JGC
0yBXQvuXQ5yqjaTSUnEVjUTx4F8F4QH7odwrOd4W0UNQLcPIGNzPwK08e7NktAYnmmMRYC/IGN4X
vA5C3DeuUlG3Tovx5hDu6s95MTdgO+R4Jc5FMtnylZDWxteFrsjW/+w4GXGxHX1zm/a4AI8NsM0d
87rnQjEAXY/jahKfOFJLpxukQ5L6WdIWO8RQvcSi9u0OlAH+EjP4XZ95Dwc6AfRBTkjScxo1xB0Y
84waF7D1WOX/D9c2RG1COF9wEUx4a0LEXOTP8bBzANpJcq29nkqB0KddIyXWzhcNyJJLFYOZ2DtZ
2tb5Wp2q2/9aXwPYHg2q7xdV6YyOhNoAa7QSRbl9q1c3g/n2nKkZ+tcRn0dqm35Dpy1K390rl1Cj
tk8ViSWiP5NBBhUXYvOB1AvNlkDs/yVqc4j1SRA7O8MVaSstGEoGk8Ha4kIuZLo64Czjb+DVOkhF
JXeffjUrjnqK5SYn7lwJGu5TgAbMsQqUyR+dW4MP2qB99hT5JKIccFKo1nRkIzAD7cPx4giTQ8ig
tbDDnoqBcDmt7p5CiG10JB0OWSrNebDBjhZY8tvmOabFtBD3FyZBlA6wK77+rJTvgWjoaGSSnLQd
rT3B3Fou9/0t6qNmTwkTiV8MVhI+NKkH+AW6R5mEPh3G6TR2R4a+UNeW65phqLiBPtFoSz5E98N7
oF+GzsyDV1QsZtYjpYA1yPzfBU4CitmrRh8j3kKG8AFRhckGHLgkv6tJ/RftyAMOAa6VNK7cv8lc
kY6bw7K4cdZhrwmlse9HC/YpuNSn8CQA7aimcNXZvjzkXC2/SpHsYK3HCbmC3nV6OhUXmB/Tjev5
aOUTJPygTn6uYOw5I3GiOO5WpdNjTnrFjWKlShtoG2ye9llgibMgwXaxin8vjKuEOrKdzvggfixI
39bxQCP0Aqi1lgfvzEnGGnS/8MbkF/jVZlmhzXEsCIqMXwilUXrhKwGFu4Mirw0bjFEpA4f82T/t
i2saOeUhzDyKgu5GH07gyMJcWsrghMe8uNSW/DnOpNvmPNy5OVd5oMKvLaY0MzswueQXm05tHzFh
hCaNXCn1U5QDeO+AibIFvVn+SFid5dpEamMD0YrYLtAF70WvobNIkxy1XIKlDxU3qzxZ3rTNgScG
DYiwXPINvhBnzjBc3bwKjy453HuWzUQeLyKAkPLjTT25WrKoR+8xWrGjXRcmXgt9lxiqqlyYVPn2
jP4j0ajoKDeljBG8GLu+a17XsNqG/kESmA/V6cN98aZ5NvXs7HmGwktqFkly9sMFP/IQKhHhjm1r
3b+WAKgDjINRjzUZS40wnbNeDwmKX93CLepioc+YvgqpnB4UZX0HT773UYy7FFNa5UCrGnEisdFx
F76vMuGfCdpppb3AxviSy5Tb9VR+w54PRc2YWxpNCEPjsaIdclqI7GYnsxtTI9z7Wllng08llRS4
H0yJDpgz1LbymKADxHod22eF2Bk/1gNAXTY/54Q6pRrNOiXqqmtTovdYbN/H8SKfa1hP0uExseZX
z31B1pF8i3vTdKpvFsCpl1hC/O8kfYaYWTXbSW2iO3zae4W4HBqiBNMQxQxmdv+qk9Bi+S1bm7fn
bajqpk8UGGmwtxAiyAUw1pvWjTjZoBQTK0vu7l8D3G1ScZDneptYHjB7QggKBXAoQk36Ia6kUF+b
xCJjJpHAWudvUWYNGhkYjmt2RXDsJU6+ZqsIhmNomdcN6SMSwRPBQ9hZGScqg/Z/PB/2dPwONwU9
x6OehEUaFJ09Kuou+Q3/vgyzdaoK4ea/AGXWlrgi6DSz2dG0KvSFjJGhjx6SK1Mo5xicplcTdPq/
86lNt6nyV5ZgBuWsryuIxwNlYNwhnUwCwBGn9ClCdxkwwwGlFhMWpjWlBnNSUIMSTk322XmiJJ98
42BI3EI6vJ2VC73xnpFFCY5aKu0UtxGl5TXy7DfuYC5halQmcM64OZzT7lMcYuJf+EBSwJ954HbO
otv81c03cBH2fKLoH3zgF5hjZMKsQ906MKBE3S9Mi+z2nU1qInAEOCT81REUDON/2tEWE0cpAX16
EMcA1iY/ozjc2nhPLUAAG+u3QUBSz2QTZDOHfIKOw3OxGZGv4Rr8D2anVE/ZAFjW9ydthtT7MBxO
q9OlsF8heqGLfCiXe5j5U1/+RRUEM75Cbwoj8hRn83NoW5GZ0H6HmxjEXVkYqexCnB9hg3YDC6/0
a52I6aa8B7ziZOv2f5+DfIcjmsUzTwERoscNgFrjjXhNegJjHRbNz+tU27RRRaFDhRJQO1Mi2tpW
y1ZIeznSKCpu8RfvTjzmwdEwU8HkZg0XvEA1K6fBcy5gOiWqa6ivw2jFJjPC+1mmA8ucguNXOLLT
zMnV2FMQhw3qPh6Cxu6UH9ELrnSmsIK8sR33iD/5hC2JOn9pIB1iNPoJHjKIs3jBxyhaiKSjbX7K
9x/3BaKA0NSvtwI68fS2pct53qSw3VvxLVa6AZnVp1vKvZCRNIP1nXRFOSjnC8X7cSANTiUMFu31
6PDQQlAeBs0Qwd3+82pU2haiZMHN015ppEpGr1LtBsKumBIvB3XI1W6qFDbQL7q2shuhK5GTYxn/
98Ccs/RCooD0cLRN5D8+mMuOydPz01HVuxX6lnqhykHx563tuBJs3LZIPgGTsj9uVNIHRJET9up0
XGLDBiCF/yhqUjjaF/oF2kkRGj3cbjMfd9VZnlEgttAaW7S2x9EeU2SQ3kcI/JpfQ3sywH/UR+x7
xC0bebIePyF7vlMU2upqpBICGk6wmX4NqER4ggNhxY66RKLSGwGkjrw+JoXOlIG8PGcOAWqr4kPH
55V2YP+DaUg+6moWx1xkRGqGthyOvbZ2DjsYYI75hQiza6gLR/FSxV8cuRj+ZZ8ZO0KIGWruOrTq
vynEHJqpLWPdlanoYiFeHx3fa7c9F5UskjQo9nnMpF3/Z/2GFUfq7fPcBMcNT6b4nVVhVH+nLng+
O+qE20xKr64Qvqiauk4R9PMdHM6EJ/SwUzWVMQX0Vn2jfhwoesHS/ilqighgVzJUqCBAe6FGli9E
GeFvHadMszwxHfwcy0ViNQxNc4S8wDNJd/p2ZihjroND8Qm9vUKlPua5kdF5liebZfHgfnxpbhBL
EyOp1DHL0CVpqmRAcuBGjGOT8AZjDhn15qqDJRZsLNbxXj+jfVKvJdnzlyLMnlY6JIhrLJM+n1PZ
SmElHWskSzBGYsALv+C6fEUqPTwFZ94XgY9yCIX8cu7C7X9M95yoX4nxIUS4/jEQU5HKmQ6Nhu6A
xxbY7vJtjkEI+iL/lqUlBmGxLNJyDa5vSYkM6Qt6nWWylaHpJuVWLhJBuDYAZXGI8iY/JPwIFfAt
TC2h+Yloz5L5fBwLRUcmpm3NzGqcNCClJyi/aEIdgatOKXO2AFn1gBS82qtvpc0jsggG4Q0U+9pj
eQTLWZEAVsLaydKaVgM08qUCjnZPyhKQtsQZc3UzgO/Tex2wZn0vyB/9CIjv7/XhXuUHAPBHixXB
8Hb67+VH5t+3v27GvG0RsGD6j7vIj+Lc21PrRb8M9OLhx17RRC1k/qK84CDoJvWzG2g5qroZ4yz4
UBLqu/xCR8eAqmvktD0i+5mBTknQNaNLv74svm76djP03RqtEYi1gUmBaiQwYEH8+YO5Ub/qG8Pi
xJ0Q0oGGP6kxlVPmqsqGsXhD/akP1ZOWd0Omxcg3+1rjUsd2L7y7KdoRjBxh68Lt6m/xuYjg7/dz
n5WPesqOMeqfpoKUg6/qHSB6ZJ+QOVnCmSpGvjXM9CSLaqtxh2fSR5a8nWbasfXh/nI125S1oXYO
V4nSipTx5LjLDV6CV3V7lTm6eV9rbUb2LCdcjwAqCBqGDu3huVHTx+e0odCvlkkl2ZHQhqYFK3Pu
hGznNQqRX0xmxuMtYhX/4SDaMPqy+W6pQ2EtIZ0Z+pQc1Fz36H9zH/xPRaI14Hgra98Vqs6Q5Wf5
DqUkmwymhYJGiBRiIcVFpHF5ScnSb6r3QvvXokK6SbnbldmvoxGfeSbYa3IT/gUkyp2uobqYybf1
R25ZNyMYlX5w4TALmf+ePKOMFLd+aBcCLwfzySoFuhBuFbPFmOH3XD4N4ZVwTY+7xlEevWN3AzJQ
RBKmJgi4eGdmIe7fBuX7VSzQlvbhOuY5ezQW1kkZ/t4XrjO7mCTmUp6RreWHKTy9fgZLgpuPeRKV
zVY3m8pu5y2wvldyltryhfxNhVaxBD7Qm7NRXQXzaUT4MU+aWXRKhPVrjHOu172cfgs8J0JfiONV
Ibo113WmLLhbC1/n3wqwhKDBAwP6YyFkIavhGKGpT8Sf3XbeGyl421Xz61KpMj6QUwk7hLT5By1v
+MtA5QLd3uvEWd67ToVrotq6k8GYe+wRJQbirm/hsfIgIMi4CMpJ7HyBiQ5zl5C0Sd9WZy2mTO/G
nC+nHWp8o+CISvj6FOYQs+NJ1qBZwc5JrPYrdnZTvhKp8HtExlnzhxfDqUgzzDHXlfIWjnuisGaW
5aRQ/BDzHFpPZcZhJu2JRv7UgOGk+b4FIqKyYGmZj1qgn3O0OZejU1EaKpCO/2DGI7ChN+/j43vE
hlX+4LkxFUtAOnrbZMsTP6sMNTcUcx+v3rhL6Qve5pWgNOHJbrPfKnm+Lpn97j9TBmeqjOr2dHv6
rqf1WCWxiOokHzgs3GsElS1svEU7gUHQ2goLoKwdSwkeLZ40MQXS3QslYgfqhGIZn5n4u3AozVK4
sSIsoxlj2oKsMXbdFernHsq94awlO8f4B27MLJ87Ag+ttLYsv8vCJDDYID9QHn/f6CXu67nnG/34
E9LZehl+DvJOxVZ8vAKEQfPMHJzhP6KFcR065Ryzaz8Gh2wBZrTX61m2AZOZIVs8sjFJqamCNiyz
OMEdFOJr802SNEBtGDgfT00LKOXUahMGW3S5FMxewaQr+WtEv0AgQACMmxR2QsgR/GkZv7L737nr
ojc5PY1rLyAHS2debuWpY28ow2hVpEeyx0HehZUGXv7tegxALXqWp2hHIhkA9SgGluvS/zzHt14A
biN6c5AuHAM6EcmiDrC6UQ1Mjl4RscwCF7C+ZQ06oIfIpaQEKKyncmX/BxH1DcwHTNX7aZ6jxi7O
BfxZ6A58A/1EmVz8vg0koe/933I9zKIj3YWnUqIV78eun111cBIKObiQdKkyAz7Rgc0eHiiLMqNd
xhkFl4XmdTyUW2TPUAF1q2SEZpalwtKIQdF1qJkZc7/FxLFsvJpbphJpXwu2iIj48OLcp2/l0YkM
7sprfEafW9dTPPtWDPb6Zq4U0A7aRUxnk7j9S9/aFYIzEkG08KGgmL6ZVQyesIHdadO2unhDWmqf
ONGKJwDKECXFgKL1V2gDdTWvMhwu6ERFLrEPk87DiDYXjVCX8GXeow/xRKFMTepD32U1Cac6wwoV
BccPqnODwXRKSsFPujJ1FOHk9GjyD65fpyCpdIkrknJbvSHnJHlJAXKQdvT1pUbMT9kSrW9ZyKHn
S+Fgmbpo3JT5RRkJUwhqYc5bbbw+MnBGvjwPROJ5iHt0bXZ3G28eIGnOgW5jJssIhiyty82qla51
f13iKYd0SbIpPyvptip5WXMYucUjBIC3DSbr0riAVPR96uOBb5K4bsoxZS6fae3b+l7JfzrkaQx4
45E2xqnfkEtzK/nZ7m2jXCEg3x63ZiNbE/+fuFPMfY+/lzECt6LlBQ3kFCcCbaLmCqNdhMyNXpZg
En4AF0vxJWoU404RX/pnK7bwEPH2xn5Lj+mPwIh7KsYJY0TkaKY3M4yeRQPWH67hbKxYTlyMulR7
YenCq4zxn4t1L9sR9aomTVmYslrUHdt7ryGHyC7n79nLdAoMMypxAJ+buqMO3AuY0+KXXepn3v+b
aE7UP+jK5CJhnLJDj985G3e0A1hNUmArDxGpdDmYxQ6nvq90y8AOqlh4VqnV/pjwdTMei1jOgE9F
I9gR1hULROm4HgZNI3R9znDMa7gs5i6ha5n2KjR+tJgCpudNnm3G3IGvCnXTspRyuOg2GbmhWAxU
S/PcquF6Sf6/5wK8yajr6uenFHAxua+eUnhMR1tAImA3QF9tCteceabuyJq2ZztsV19zYImScBHp
4mX96zr9M6oy9cxkqXKZovi28iGHh3KUJPWWqMcTUARJw9RhPvI82z9IZVDzAFyJ+9NeGXgJZlPb
ZAxMtDKZh4gn1E+noFLnX7kEM85Pxokq5W01bUg1hOcJmD4arzO1pCon4UPGolVXDQ5ZuNr/Mdv3
nqUM5P4r/viDHf7/TtM84vsbdveGNBX8qhFMlvgbqFCI6q1Qvrq6aQ5SrZd7T67a0cehhPwIh/q4
mGrvDFFZ0980QWB6BjECNhHt0GgHclev1cGFSAiodGktaazooo4FeGbkdwz/8TlosVQTkPOwApOf
L3IY9UkhnkryHMpHQF/OsQREBvV7iHvoR4Q8ZrwbKVBdk5hpmT9OLfArgrS99ND0RtjNBzq3KZgH
h0ipl2h6ZqMrGn5RdGoN/9m5msN1p54vcFpFkz/JsHAmskelxaDIU6IR5rygzqnjDimHMkqpFqB5
58aVFep9lUY4Pn/F3gGGpdPRjvdmYhagsNUMZ68DQgrREGFF4m09vkEkGE90cP0MHGFfv8ZFs+K5
uKS0akVbr0v2huRSjCg9IxUosRzpJr4eu5KN5z6yiltV7i/tM9cKO7k8eGbDjPsU6yPl/SjOqYLl
AjkqWGoT46h5m7YmjAHrU9NbgzV41MacLvSQGie9HCUEGxO9jdnXrZEIn9WUYL21nH5D2lAILW6J
LtCzjkCww2PHpchaTIORdkB6bkM2WfIZCxvuZzdB7fh+GF1iGp0rKB1PizyeSArBKA0MogAzRjt+
0GKQYakWV6pAzkcXxVnbkc+kb7h4kTvz28sSEEBwroDUpTzfJuPXNjn6EJ//i8w63kPQ+WGQEBHK
KNGy4t8zClxRnjEPdhupyPE3UX0YFWBsNRJBjLNmhJpOgK7lOdS1xOsRFjmhUoUkBsv/FfqEF6l4
pXAbfmaz8NnySzv+fg6QZHT7yLJJk46ffSU1LBSaF6H7BkbHFHP4LWwpWgKA+32623zsNFEqWxPx
AqYWoL0NwqL7xJloR7ph8TxvX44JufBnYVO2btp6u/l+yvNi7I/Y9e52Luuh86Ma7QIEJaWj0nJe
UcEwa9bU3fMRe24fNGn+NPFT4bVO7ylqRmGFdLtN+McRdb8ue8T7Nq7paX6LNKJx2SYHZfgnVflB
ALuh+7YbmLpAVu/VJVidhDrbWOLR1zwf1LikwxPrDLnt5VIncVKb7+QXQmxMfTOwBYpSQbbuYKGb
Gd8g+AMT+Bf6UzVnHN/qO3mmQy1eO1OaoIbJesMnyigQSRfI7cs+GkpFOtGTbenk1KDegwOMiWqN
AzVFfouO1POSZHEOP+zUaImVgTG/E9QXKtFXTTvcJ4dPF4HEiMN2b32k86RSpiDr9YApXNRrIwH8
6XJkB2Wc3HnubwzFhFeuV9fjWJFTsIH0/t7jot678Yl6H903ABBVdIHUZ28WpDcHruhchds96SIN
udsaOz1OPHdKEC9RuKhZb8OP26haHpsljywQZq9wlz0ZoZil9vl5NTn991Tf/e5KsVVCrQ6R9yCQ
6wAZtEr87HzByJorHCi2SitbcDKNY77X39iTGlKbdKBJSYWDUnqF2OxvTfuPIqq34hGABDHARaC4
ut7ICn6NrQohjyRs/8HvvaCHP5pd2SFFHPZE+PuTfF9HwTSGdfRCF9z6WPsmbuz1E9sA4TSWLOFB
nV++TA5ZmmXHDlyCW79oM8A0ZB4KuTzn6XrVO33/dhf8SPYLndwzdfd7RuVIUsciGHA3xMAgp7W0
ofP7XLl49FkTVjZ6XOZKOhCx2oJO18cINfinVoyJmui6G/lNxWrQZJikG3Qv4v3clNIQfksK1MIJ
rkoNOiO/4QLJPmTykO81eItj+1FN7iySXoQE/WM7tBJOIywBLdxXPDzIvzIolAcquIMAaecwkeLv
7orQWywt9Cu1mEtU4CvsBZS6AN6BzIlQfYebSf4+IKaZ/VmXlW31xPUt/0etZdbyGBr9dl4YFDEO
5Aos5GNjU5qeSkP5Ejg1tGNnRlwOC3BZHOyD02xXeCGL1RAfmG8AbKFB2cmIdmgYv/QJABgSAqts
rvCprPGOnza+V8vFW1aGkElHQKvD+OMzWIR5lX8kchlKoDBeikiujgfNEG8F+kJksFB1qbOVJ2QY
hEmkl+bD7AT6vLgFo4oPpRuBJjWJoUNoS3AiBM4YHC+96H1Zxwy1DNsRN6nZyQUCHElF1xz4zzJj
yem660JK1qZCghHmAy1FBebCWpYqlOHNNRymaTENUlLRAlxzkadWdNxstWMwb4gyzOEYT2xxo/8h
AEC0YEPUTxJJFPsjQARqxFPGLzoxHzJk/YzbuYOwdvxIIVF2DQyFr/18EMU5vNHGWH2cr0w3Gpun
5XBsuzXeKeNH1xNwKhQbKSN0PwqIPyaMam892TXcrmioapd1FUa7NJkbjTp59zTRgjdXVlh7YpIu
Al9V7x7OT9HFoqJlXaxt+08V63WfFBnGCkPr6/RPPkij7JLoxPLrWgwV9wRU5aZP13dFqXYzda6d
7W27phXtLRRnzlRQgHUkJqR/fV1V1dIp5Z3khfto0hfBrydI7WCAGAbNiUmdLFcilnI/USvN0wni
Kbs9wjOGmZ6az5NaxjL2t80E7afeGyn5Qy6XVgZg3TJtzcsb46/WdIUvaGB9QxzdAZsEbbVmYH3G
yLwXaQwS8u84lADIlwivO/ELQJTbYjtKTybYn4rcJ96roDJIdYcCxu3pFIT2mnVer+Il94XbeoJA
F//C1IthOdT/Hcas7K/l2wGXPSDdIAN+/gldlpfuEDRh/YC/P3UODXV8TukqnwCNNZ2O2Pc/r2oo
a/9PgCp2KzzdnM+FvkYKW00BkPOl75jkxvsmze6a01z8y7lUX+jmyWzxax1OdfV9kDfuhv8Khewm
hQvfEdTNTi24WZdOBload9sU9HcxG4nwV+xXsVk/IFwp8ksgrfIOggdAKGxR6qssESGFVwGobNcT
ECVzVdThf6F3mSxrTB+Drb26iLjbPPmzcppbXFiHfo2L0Td6uwE4lTCMhoJr8XBGU7YJcv5VVc6f
xZv5OcUzzgnYOz3MucoYq6RLgd2VT5bvXhQ/JcTCkMxpREpyRDD5TeTM3f1eBFQ3gPAtZpQyiX1j
aClNooNUeOfv6u6NQ4UJeLyxDtgeNA6MviNqTPk1gt/r3Yc0FGnRhaSW0Lh/quL81hPSTkzdRswg
/o7w0jipkL2CYKsR+aqhn919GLPxcM5+r38gP039W5b9NeggyngIUl7PK5O5nzXN7xOh0Vqbeloh
EQrIO/sIJnEkaRlk9nDwTZG8nOpVZo2gpz6jQ7iHgAQIVvIcvZrScs2/VUpZGbQo4BMfPtlYxAzW
tAF4PmefUe+zWRGhBUgo9UWiaiWuOj5udyLcJMTL8jiWqDNZZ9rMoHT3nxChdj+xy+FxOB9Swzqd
tYW30ZDeAxgQlvUp/ydM6mK09MSJmvNVX/ubk3LLs2bixkMP3mPtmwdqOv3ZAI7Gtej+kK4elj8P
v7gtdunCB/OnO0CWgP5oHdjoYLHw8s1IU9+49ZjQXnprCA3X3mHhqnp3bfBVWPEullovUrzLTLO8
vWHOKmNe6Tu9c4tOj1o29VFyIqDA7/QQuN6qJoVySt4/TKGrxrbaiu9e4m2hlLCJKbn2uhblRqaG
ntkilwoYO6jQs/D4f69oZJXk+rPdBrSxIwYULy1mlfUoIFPS6BDDAE8M2NrG4JFBDU4p8qMYVCia
gcAoHbrO4zOH8kxxJ3BWB42olR+HVX8A1zpMVPsuRK1e4x9DTLCS9qMpnPNL7++ABaJ7tFfrT5rw
+66zCkvSy2Mtxud6WPhmpEBitVgn3VLr+/FFrPFAAKYcbGKjXKbUS3VhGz3+VUbFbaaeIwi3T57U
o4cCfXJ/dQ8NAzwGjVNJfvw5TgzEvgFXlNvlEIEfDGpIGjXy+xHBTI1ezvGng7HGpYwTqEPbknn9
kj1lLVrIT6yYsTSuYEylpRVK9NQLkOFm2EDLCdTTtLL+uhcZ2lEvuG85BWh6H8USoz9y5hUgXjV5
M7HZypcAaxUQbeJLdjkeyXXTQ0NC1fAqCvBnnv+gSOsrGc/oG5w93vEh5UqIcVKTymZoWMGZn+xz
lai1q9pe/q5ALOExdHerQ6noMV27A9BrjvhwSTrEOO/Wsc6a4953HD5bBeVDFCmXx1xKDZIMdEef
x5X3wlG16wY+3zhJlw6+C/7qp5ar5GRuK19FHG+7dDVKA6zqj9jClL671J846ShX+GJ5ThOrCCh6
9ZRTrp73B82Q7JckxjEvJjKJnj7Wvoulbm1voh4FDLWHi+anjZYNi5G6s0l8h17qE23YQRs9TkJm
TJZPhriihpwXL2rGVMBJDce+Tibpn0idy6R3OnaGwO5DZCwmyi1iIKgWlSHbXdOPUo4fJUmGMqva
2ybt1I9RjswPVi67jY61CciwtUewaJ4DuDY8dft4XKuDIMwCR8DYp4qoZf7oHvomB9ZYh3DUBzdH
LEAQiEgNcCq43Q6zMFTLKCPURLOuE64pE6PzGkOV+QqUmL9hUNxZc0MFel+xL8m5jY/9DtpCR5c3
P/AA3xUnTQchft+JssQqWdU6972t46neDqVmVHQtFVvxDb4VNl6DnZJ9xPTXBPt+9EWsJUrBDeNK
vKevjbwdNX4YvDD0PHI/IBTmokm7Zqkqm11iOnQyqccNTJosHAtPRfgl2AZAZ6NGdb8XiXYrN0Cd
pyuh+Nfkr+86UXHMaie7ccTt4iFa0+r0hO4hg7/YOsQPkPO6UL2kzC8Q26uImL2GChYQ1fGzh0lM
/5OgeGiV9F1G5cIygeL36vdwZdbSEOpwjf6MgpmOC1Lo1hChpPUrYQZgfAE4Zb9SBs7t5v7nLG6e
/YB1pf1sPFMK3+sw07wl8GP4EHfJVCgEMOcSVrO8fpt/lHw8KgxwTAz/RTRI+SARCC8d6b+sx9kx
YutUTSQCAHKZMoQrmKvba2BkE41kh25sP9eMZC6JhA4a36Gl456b9IgpFqWqcZ2JW6y1Q7q15hsV
ZSUwpCzoMqmzXmHW0Nx54Ndvh3iPYS+oZLTXwaeSCtIy6qhrb8bVVKNjZzPrRhQ2sc/At4oRmSm7
QU4EjR0wF3naALE7ZyRfcmFJCPiZGjO9MIfuCg7c4VshjGvaW+T+FdZlw0RL1sEVxQbvnN4PJQjG
qmZd1H2a75bbvwOOCp+QkOiFaHFqB7Tnl60Gwht2gyh3xsPNkKQU7x9q9lycOkpQta5+J78IGPbH
xq8TrF2cO2l0uzRwXEJ0QoxSjCu45KCjSpAl9NDz33yGq8TUWWYrlELJwaC1mPtMQbPIsos1z4fB
Z6tVJEeBZu4V792LGW64IH9sYYMNeYcTcSDK5VJhXC25sWPUXd2WgatvmrdWl6EhHkVbGo1zqcFg
LzJNAZSGpUWXQAft86SOgOGXkXiAM7vX7MZ2vyw8I8uvB7lxuboRjhbk3Pc4NYwVdfGhO/bqjC+t
IH9zZON8OoRBpX7xHNp/kftk5wUbdN7OMtPWvw2VQZaj3dFY58DM7SU8SFSD2wHpd6qIKmGostQk
Wcj0YB04lI1W3tEapTNh0yl1ZbDMarhA2fsr+39uY0K2jotPQBfwBsq6Jlgo72ThP7cUTL6JCtoR
WNfAUfA2iBQiL93km23IFvEHaNypOorVbX33X542B5qS5rH+CNJv2IJZfL7mZNx955ATpqhT7511
zLIK4pG4Hy6/mr1iBVlWqEqq0X/8tkurIQxKtDiXIFmUHqx9nKdZdxdHobJHh8yziRcrCTjsBtsH
n9ryaw3OQ/BjXjpBnNTY2GuI5V53iempZrxGIkzqXRZ5TWnyLRb3X66bfm8LRDJLgwofwdyhohZu
3dQ616Csu7MKnv+LmAwvRjnMBkY2xCAtxra8ENWKW6RG1C5W3rwn3Oo475jsVTE3x4CWgdeQYk6N
LeHCOoh7pTaSRT7DDqv6XANs/St/LeTuWFpDODZhO/IAW6eGk6jV8wzrLgl0WmHOu2ykRph5W4N2
/2qMPFbpxVLaXMlvbku3UxYqw1nsVdwLom3bWpKGvZRJBx+CoFWp4mtj54XUVwGpQLCyii8x/gsq
/YoWLmJXN+hiNsr1bYmDcNtsdhVilMbMD5y/CQZQVLnyX6/zAESt+AKKxILG/26GP+qMaxvWOcCu
Wju0S/qreMHPYO7Ts/ZP0QpDqCbjYsfQpDhdTHpRHWphYBKqN84BZthOfsr9olCHwregXNUmv9QI
A8C0g0+VL0d3z10gKh0sAq/JuyYyhRZleHpLU2d6JThB75wuq+zhhFIA+8njNHoT5sbRk3fnraFO
j2n5bhitLSYylKOc80ll+6CVJuGipSnSTkztJMVaJ0Y5Fgz2RBYEXgjSWdGc648wDH8ZSEG7QNtE
Oi+/qaSDF2ULOtYcTGEpt5fSODhsgoSyD0OiQFc7LBXGEYgXN2rqq/A3zkv9mmHD5LwovGfS8E7q
URGoQ36wwW35wVQj9NzBV8e7thydjspaxdpgVjAi3DPHMfHXrxFlMFs0NmjrNVWg2V87KENw6KvG
xVuoYnK0dHgb1sH13+wKlyP6Y/UoKT34lyO+iTgL4KbHvkdp3uqumQy1j7+urbyin357WPuyvPr8
dP2drJC8xII1TBkB/XvPDJ/lmjMrwwDhMt0RBZ6HPYxr6e0TdW/9b1bubk1FE70MHsrFdBTL7xWK
5RKUDNz4PFyS5nd+F9f59KeHFXJXR+ASMknrzQwJldN/RqGAeW/3F27WpGys2sJf/WEunsRdb8lM
5c6aTWywrQtwVJs6ch2cHtowvlsKuMcdgQgYEh/CXU/WDEkhJx1RzmBhURdBzB/20JZMt3CCdGlj
pxlaEqB5Lr+LVeV0vg2jbCLa5UD09W3oTeRPAB7ZCaqRnths2JWLmOmHjMxEIeovjZ09NyUjHLvY
2fTEBqlIgyTv6Zm0AukfxZSC4/cjHj+tReI2RtBoalHyeNd1A7f7AfH3lXcgUDAAicuGSygTYw39
shQZ+GA+8YUrOiWCGEm1rPyY41S0oejnkvwM9fX4xzPOO/Mf2TSAl5oGLjgA2RfFUCXyM4KTyuqk
x9YI296K64vZnJSqLoRTWkcyHP13JrOKYfwAVCLThjUBygq8yCD2Pnv69dIZfmU3juCCExSebDrX
fkFRyTA8gT4FDgxnu49IQfqNox8OvVk8gn32yvFxh1XOKlgGZe/5uBY/R9Q5q5Zch4FsZsUtq7C+
IEmTYMdGLNASkkz4i+6NrNs7CbxKaywfGzIt46X529utvSBavIFDW8iS5FRV4dGQ4EIhAKlH2gEF
tkluWA+SWY+AZ4r80OJL44CPi0C/p/cBpa/oDBnHT223SKAIDjjs4U2yHoOo5P+myQOax9ClRcgf
H4AlmEQLB0idVSLxRq00eJq660otKVdw4pGMN4t2m8CiK9ng8NHFGBd3fQUYeDXRqfCKsg2K1mc5
7tbzRa+ZbF90HSWsxfxwcORdVfKE449dklNTvtg66Py9V7PZYR/8J/I5CTig7Phdxjlo1dwvSMer
FYJEt4TQ8kifiaZ6cRvo9yxVhKP5ZiWNBniUW8EbngONrdzdMCEtIdFM/j1OyBOJNQpzBw4oyMRm
Q2bIwxbuo9zNFvbU194jvPRgO85D9o2/3kVsCBOr+JTZ79AhQszuyDvmgmdujBf/mC7IMeyrBo2g
3TF41Cd8+/zZ91AK+KUloFG65rhivKXVYzhDyz9AKlT+k6jYt9ZTPOWfcL1HD2sJSsNhgk3L5ufU
j9WyXwE3P3+bUold+juLcFcyG91/2mON3OwXC5w9uTBHJSouIO3H90z+M1ri/ec5GFFJQAsU68+R
rWhOOkhmdKPxIYItBGlgt9oLoKoz3pCYIP5f18NysJfADGyXolu8nQRXVezzPf2J/MKqhvyYAzP3
K51jIU6HAutGmN7+1Q+18MULwP49TFlAUz1wS1CSIHoiKX07oHdqx/kKlidMb7y9gwrhtk1PUK9L
7q2r5zD/fJAtePSov/lzXYqC1ppjmtdipSzxF7XIKJYbHcoT6Pv7zDV8HRzdkLODuftB51XIMeeL
6fmndUgHFebdcrWwF8NOlDn5+QNqGEtFHnb7LMWM5K6Z1DLI3j6/rwmYFNfS9PtlzH6LUGNDQXaO
jBocpJAjDOW9XLq6HzL9pgrPnjoLRGBD94E071f0oWhYUjllY0lvApIXwPEuE03Etcl8UcjmuewM
lItix3myfJTAiUp3w8K23tnsVj3V3pGMk0ZbxI7paWZpya7MvwqRUXenAdJVPktNNH7aj28aXQpE
Ah7dHOrn1o5OQfFc8UW1n6BFchMhBmqBr/adrHVyoL2WMVTOeSyzYC6bSDSoorTcpsItRzET2IE7
S1EClR3VY0Cy+jUw5NdhOz5FUNMEky3DtX638sUv0KcJleRvPGzGBFWcXWHJ9Wfdsg42SwZwIPPK
dr1oJqDhatxBHPJzeRgLFJE1DMDBjOzfg3SovzizqmpLQLZRmqH5GBf5DbhPbRBnWuqv6WNNp+6U
2VZuwI96WULqr9D/UPQh9yIdIEXhliOwyfHCQU1pfh/oql3V02XJRNK2XNY0qDFqfR4r8N5Bv5yj
WSZK/vfUnLfaS9L8S3e1VXMmp6qlMlg4wr8nOm5y/ugq3sxlkKYkAG3ySm+LB/RA/LdAT3GMfSXc
RuOHaadZr0ilXvaiDHCr2j8IyjFz1yGGQoEwYIbX8ZFMPvbSEW1jlvRBJ3Lt2tokae1V6++dvXnm
R51IOfWCWBWYr7u8vCEDMzhcLtb0UmIzpLJS/AFrt05+9REJmXnX5MzqrG2XMgCLG0D3FT+SIA7e
Zn3t42gM6Mit4jCnrzlubalSvZE1bBY05d98QOHv1m9OM5zSfagG4q3hd8eDF35VB0yvID4PgOwe
2gobBwWHF30Rq/3eTdS6/Zn963tNsXPArWtiEq+jTaqqdu7eF1Dtc0t7QvjaWnRA9ctxBNKw1xqj
EJOat9DX4QPoCG42aYPBWBkcAtlmaH07+VrxGsHRKkZKgV4QkUsYHKXT0nQ14+8fUGVf/HansDLp
B2xyTFR/45oppsnp51PPfN0SMb4GWLfrZf+tSxVdNqUQQ4pqCXzTN3JMxkZZkwNTjMYGLEYmNxwr
cB0owz0K/54goeCrVew5xgdWwLQjXDjl2GrFVAqgN9kRKAkdcipkSadKMPnU6COJQmqoNyXvzHNo
gt15ZZHddgvpd5mM+obqE94Fyv/9Jv5z9GD33ddx3B1Bbd/yvzNORDwm35mMKWGuhbLz/mCACwBv
t5lq7bffT5I4N+CTAoADr7mNeQwD6n4bAuMIQyO5yAuYiaPcsAdiXklfw2mTTfJ7gqNVENv6O1DU
qoT+JsEgVw+NNRS9Gj+/7U1sGPwacqs48bHqXXNJrUqANgqsg6D9blPq9xNd7ETDr/2OkCut1Pk3
/Ya6pp2AkHoyoTmmmhxELSN9gr1L3TLcl7+Y6v1ZO5dWzPFQz5q7n1ESo2u67FG+YF8VyGUiVUVD
xpPE1j0LGRDFcYq9+DK4ldItwd+v+pckd6WtqNXuUXkF2smH6Kr+nNid+bmTOKToXqqkwYHHhxcw
SJqKCSaQlxYG4/uO6gY+GyCFbQ4CWV74+c3Kz9D/IEUmhwEfTpsXGy2Ht2NqODOqVt1Zeq7W4Ffa
7ZVVl+P6grrzkY2FSPQ7gw3XIuq3HIihb9W/7CuEA6vSGEjHyPDNcaxmuVw04z4sQP+gUAbFroKV
o3Dvtn8BONGnWmYGp2zw6lxSILLZFaxOikwl4EvHhptLlc0KmIfqrFj5I04rzIoXVyAU3x+8p92X
O1VtNsPCXo69S55s5x06oGySJuoaWokmOilaVETE0fNTduzKjAXBYsBw1ly4QbWlR671qELyAsYR
aoMNro4R74XLCUpIlc73gVvWwk0cB9+X2q6p9wueKmA0t02NCJSnSOOFwEDW9dN604bxbRNGjDgb
6ZQWyEEGn0z1ctQyQf+g81/3DF5SW+rBeWumN72HjP7Kkwp4dJDsOwsYmYKZyj3+XKCMmDuHf6oY
wvOXv21WBDXmuMBjkeYHciJOCNnGotg2qk99zO+OSa8FWdRXqdQas5ISvHoADDKgDMXx2ryUuXxh
zjdVVl5CO1zilM+fln9H6yQNCn0MqipHbjrBJ50rlK9Y/JgILhBJ8JjPB9Z4w6YIeHase4+1ahc9
iiynTHswNGymsNFzSjairFlJ2nf+I5sRphKBVPY6zxKwJZ9bgY5KwirvkBtxTxlAq5r5wk9XYp/n
9MJZRuxv0KHcbBEYMtzeW5CYyUpplzCiLCANHMt0OfdYBt+FlsvgPQf6HAHc9YbthifUzL5Zcm1B
2/HdDK4gpw9FIFGT+8Af2v37hbOuxQgxH160w+wCZJ9WX7FsiyRYbjqdBn/2+6QhQjRxKWSaGNNo
dFyRBlNIvjOdtRn8IJMlPFLm7CbFyCb7Q0LjXeKY1S99d+UXMIVGRNIDziLUEzbYcJrOxvbvZ7aS
Nm0qUXosp19Yuc78U7dLenm43wK+m71uh1a4l0p5pIaS7QApzAFeBhxeeudaKc7rcVsBrF/TihgH
yR42CvOk+jXVfk3nCKpYwaYmOEGesgun2XL45yVArOVoiwHLx0CW/calSein/vCOKUDmJAAIMH1D
umtyDPx3WjjCN9ZLgAEi0C8Y35IM9p6wiEsowOKc0e+uN07Ab1KpKbB54SUCsrrN57fo/s+AVCcI
s2iysBPj7rN0Jg8I15bNaQPrZuMeKpVoNKYTMja85xf/4YCmpeLzoxBdjC53H8zE2s0yFYMBhKex
RPERru9g/IDmBFWU3DZVSzRiuLLG3guiU4fUchlgJot4Oo0PPIdP4OiQsjB/FaX481k2JXoyy1JP
+TFrsTCAQzDlmLlgQdUn1M8FwpBKebTkFqTnZi93go+AOeTGQ4g1Vt++Wx2gL/o6wL+L6mzIMZkI
1NGdN/qd92t002Pp1M2o/eiW7kdMNXW03Xp88AIlgZ+mbkghPkPiCJa2Db0/elHiSeaahGy08L1D
6A4D//WQTEa85rK4noccbuR1Jy2Tee4r1DmnXzNF8mzZ70GuE89N+S+oB7dy/BsdCBj60UDWqhQY
2CfooUctBkOodqXLa0sqqq382cwOH++SqIYkAsn+kH1c6MtHvW+pDU/BHVPrVx4OJJQEgqaYbHnb
OOerb12nhl91fihyX3gpZWaad2C6cXDBb6PVRsh9fJR8K6GrBTj2dYxCfS8dZBUUBe0m7cQdVs+c
OWcdq8YOAaAZK0jE8KBCudeS6ncVQAlBjEiTp17pt4JRRs1u2r+p9pzvJIJmILtWq4t9eFBqKJ3Y
cRehSdOwc45EB5S6xHKLeh30YuMTrQVSKfAh7Giys4CO/DSCXYCIKW4v39eXTzDRmNt5eDu44pWF
ubY1meQEK7HLq7BSEUYBBPZWCDPbUko2L6jBBDlkFXjBlDxSF95v4683Vpkojxcvm5skN2rry4NC
D76j8C2HYsWHZuxAPNFiWUBr1DUSFOrfviqoKSuR0tmOxjfcRZZBa2nCsg72PEK1qQM9hNEJYD93
RTkLDIs3f/INp7R4jcdtmNdWCzPBDxFlJzzdNMs7S4WX+tg911iWHtKCJF8BlhQpOPOVhNnQ4HLD
rHARkf/+bn6LDAXP5L2poSaCZ/mw3kfzTYMFH/4PZtrFrRzBESC11bE9454iYjb9iQI1Cq8xbxW4
TXlSfLV+JmMne/6434JDC+7P2nhJBUyy5i2KECdAai2qBN0tH3yf1OPh5s2vAjFOQljK6Xw1ugMb
t8bfVe4OWisVC95dqtPTiMidp+dG0uyxHZDbjh/axirAfgJoFlURduhUZ2haLyCGHZsI40sz3Wmd
6cAhsBZ/qGA+4xs2CDRSdjGnxnO+HiHf+dQyMnQbWBtdvurVUVfs9UNE8iJ3aeDSynQYv0hfOClN
GahYKeTaJHhUVjFeplKDjabVp5tnpf7L2IJirlpZhSRZNIRd59A9vap0gHLYVa5gH/Ke27U3EYGN
g3FDBDZwMq4UJo5zxnuZTnVxOovgVihXCFFEIppik3O/4ptElAu1PcsH8PMFTblrIUYAa5dkIQcs
DQXYsZg5xX9hXFtHDJaEb6TPntP0PBacOF7/m6HvhvfF6jAfGXmoeQo7ffc1rQmgNBdAgIOi8dtT
9iq+FwnTx/Wk7NiW2u3KXrlZuHuDfXKj7KBjVPUG+3o6X1F0R/2Yj7BMDE0FV31+XQfQkW92KmYc
wQ1K9Nlu6EY7VUzq8/WuyHFSXWXB/yXFIl55/bzx0HN1Z3z4FDFtDgYRV+mMdBEwjyghW3iDDAKj
WE5K9xjVPJYfDLGGm/ix7Yji6YN2mMFVM3TcjdQhapmmToaECDpbpP2ah9Q8qkM3Z3a38fRewYoj
HmVCqT5kyeZkEz+evC2KmnVX/jRC0avdlTiwSY/OArvlk4099RpqxKBdIU0f9bTXkC8FH3LjNYF+
D88ZIi8sKUwyk2ib0t9qguk1Auw9thpFYqaMz6eNVm4NvsmNSazxnBvHd+fOixDRWto5j7CnEhsR
TWb1YWru5LmfX1T4GlHaQO1234xJOfmjR8WK9NES5OA1faf/TLCtUdfkGKdMtRRkw33s6Q848gdk
uIgTXMFXgyF3Ralg240XpiLbBqKZw0zX/2VOKaP2gwlrkASUL/5HaYfK2O8wOJr/CzDPRph+2Ekd
sXY5zezkKiAAXvz5ntD6uXnDrZst/U1H324A2lYMgzMX0khDhntoq3y5he2FdJNLLxwEd2iHX1GQ
NIOvBcZxyfgiT5+MttrKBd9EwcYu6swwg1Krk1QFfYfjJFaeO5KYNL1y0a465HHtQwP5ZC6XV/gY
4xh3lpbaKsHEHOPa+7hoog0xZsEpRyuOcVa1/ySdy3rSC+Flp57bQ6a701i5Dq4DfICVlRlve9YF
LZVBrmGdDvSQfafIlyKx1bMTMvawQsKjfUPu1reRcVM6qHBMXlAwTqQ8aAoAZ4pSpGmDRAhTLRnM
o4aU7hJRPz7qx7zomnUS0TnTkYPm9a37Cj8YnE1n8alBfKL/x/fqkV6eSb7HYcAtJj4MPUnNU3lw
vATZSUcuEuXiafeIDcfAsn+bnVg4Bku0SH6kNUFdE2dzp6olLsjdTJieAHQbrz2zIeFS2uL6vYgg
VdZGX0S50MgJFwaQ27AsKLCI+t8clf4cqC9qcEss7TJZvVblmT2wIp7Ds/MxTavVNDh3/d5WM0MU
IEEDKHDfkTFugm5JvRh+JaokPGPn17AYJcNsmvAF3Qm0sw5kQ9dTTJ5haY3+GDmMb0FuqvnUKJ/E
xLymxy/qkv/JGd89EY5x68zyywIpPu4VQe+waQk40B1bkpwP9+7B0F8hmmNVPcc7Rj+L5DDsUlfy
g6aYSp2qbxGwmD3rhryE3ZR3IkejtY7g5sKZbzGNzDttCWxBU+3FuiKgerVcb5D9rfEpieZ6XOn8
wOHL/LSFbFViBUIWT2XYbYaaKJUuw1wCuQGd9zyj8lZEWZFbrxkPv+tgpRvnaBofl3apP4ugI20R
7GKMDmjz+umQpt1OjkERQCWMdxz/jl6+RDVcIKO50cce/s9o/3XJ9BXhZsTxnb5VzawAFP9VzEVP
pTE2AlPl8KPjB2thEDv5/UaBA+BjoVNgXYkv2vMhP0pjKUFU9ugwHPRl20jP4nhBRn8PlAdTjvN6
qETFzzDvornwaoesjEqS/eHM9+DKWTX4RrxNSWY3xdV+FtK2AeMPDYkSFD4Ao7hCB2twhSd3MtEe
o5ITUiULiPBwqzGmVitQCgr/VB/HOZbcBr3urPgzORaK9Kx74m3urb3u4J2V1nIwRoeY7bWfMwqC
/NW7/BOiZtzc3HQu95SxhY2Lx+uWNrsl750sPhgirysZd9GTtUnDjr99h8jD3+2U5ZPvBDSngiCV
A6YERhiIX5PLGAgoKaERXvyeF/KlmkNTyYArpiz8F/8M4IYFYSUsINFvimkBYvA7/3ZcoF5+bJAU
4q9xCjiJ6v0sQ8ngVW4gHsZN0ODwPKKVMGlrahOGl3rzHUoijk2zP+c8Bstm/yS46RSk0tLm0AtH
GbSTh4WnPhdZNVCFxrWq0Ce1RyfvozJd10H/ypdmwtA55DKTYWGyzETbuQeCb+j/2esR3HE7TDI3
bvNHv4Cn9DRA2MgsFaK5vSuyOx8oo2slh1SgpsaLg9ZtxutHl8IPKu0++fFWcnjploit4oocILmw
A4GuDK9GlUKyou1eYCiKQIcuB1Sf14Lw/KNJ3pYg3bTx0OAQubcvH5705ghMOoNwUnI4mLP6jV5U
nhW+SiJru/OXyLfii4w6ZrRfR+6hEIwD2eHbF1Liu2dweVht3USn/2kDIvHzx/U3b2LPe/6Nvcid
v0wRYoG2m1KG2er40dpzL/cenVVjkm7aZqDv6tYqQ1Gc5171dKJkzs+h2/3Pkt4m3zdaRY2A0nNW
hV4Z4YXDj2R2LMynUooTa3IafV017I4bDBowLHdrjJ8J3Sc2W3knfvCDH7g7HknDm5xa/KqN+1bp
NXS9R01Xtcj53O7v2F4F0/8HRdFR0Y7JzJJpBo8Tj0jGTPIk9VLR0K8KDaMY2UDEFc1nQOwWagVj
AFVqquLtfITtP/88MzHhotvCgqFDkB2qUnqbk+FeTY9Rdl+GniGyeP9IA7sS/l2NtakruOzhTPzz
QE83lBoxF8BELrdJKkJAdQzVChBDg27GZHQX0NdLQ4RPKi4QE7FOfX7SbyvB98cPcFzYDcRckRgk
YFlmjhxUVAGcytSx9yidey9ix6NAB5OIGCPp1yjCYlC39q6DP3DmCvnQKiAQhQaVIGwnYqRb7cq5
BHwzK2nxqYmnw+1uEopbj0v/CCuU/aNCIcAxABMq2DOrz3QZjKe0PQTEveW0HlmOymsf9fc+7tEH
v7OP3KJjrmn5gZS88Z6MgMsh9RurYeGnXVHxdQFG25HqzbAHUvwLsfPVzEEJ3Xm/7WKdFrg8SvZH
WvP7n9znuiFwb96DHCAo4AI/Jf7TlSdISz+x46pr30LFF90bjLKsr1Qi/pjVgBhvcDVfxT0/LABv
ql5WNvT+0USg/eipn4s9KwBFf1owVONpWvubzfPzDfuXJadd5uLjJU6Xhvl6QL3llOGS0EXOdwX3
wUFDkVyFFZ3zg2FR4FQkKfzCYxwvxDvJTUsYDGxHQU9F98wkkhS+cmx5Y4H6vpNr0lAkPfeZ+KIL
+S8ZhTF1LmaAytYVX+gi0VO46aSPYNxdHsGZCfa46Yx5cSm6jkaZZ0kA09Un8ocoA53bUX8e/vdF
1Oo2WKQFIxAQtIAZGIYyVk9PRnPtgOSwac+vWIwqv/mKVY151pTiteLrdmTN5We3tBq6/gGFdd9y
+FqZexB9VCetCMkWh+xV+JVl3ZXR7lXcJ8dExrRwtxSPmEQqWa28EpU/ARoFfGAmo8zO+MD7OiWf
F8LbFn9/PnbcQr4K8zd83TNbdAmAblgr+wkKZQyiXJzEJ7yxljXffbMPqvEpEWGvo3Sk+qT3wPMf
HwXIyGb+RjC9bcQgbZ4GgqnPUIkUpKt+yvnhNrrvpwiTnYp1Bg9NMNQWV923HV33ESzfzfmpEacw
8oLE+7KTtyL0KqMMRUJlJ6tBm0ER+HT/5R2XMTr3X/jL8MbeM3DP9BHCZSWQnLxA+P/lNaMOv5fw
bSfCmRdrQPrNg3OR5pKRlCbzB3jVfjUFEuIL8SQuM+0gXN4akCim048Db5s17klSjDFI78NxGjv8
eNCSp3/FtUeYN/fFJx+e6qrpD7URvIarHJRpHVkGEB8h5JsMQUJ8iaQE6mxc2vEgOLqHn9qcYsmt
vlf+e/QM3n0l+98/GGgOyL74ofjiMoAWiczo13Wn+iYmxvPM0Q8Ejrh0cumrR4ytQlT3RlYOFSnF
5IRtxwVhZfxuMl0JIKtdMOBFpsJ8IP3R5/niGtoyIpkB8/e2BkM67btzDt48aoG8jCKiPeA3YMJL
jCgBChN3COktvW4i68pSjUL2fj+xeXlwDYtf6kpvqoxrQQ72zbq05kuL7/JSl15QLdV6fkikLVGy
KCvAR6ZEOy5PH/3GwvFDsV5BYPbAW/xuty5+3aRVmHrwwH+Fax+VR5iLcvBmprx3KPeGaKQEB5Rc
zReNu9hNDjZ9q3g6QTx2W6GXS18PZJYwZKxuzNyz4uM2DC9MWXewaOW6tTsUNIJyyxtSRw8UNgII
nY3Wlxu/uTqy+nUlZBlob6UyuiemuAKwHzuq9y2zFBOAuG2+0nfNce6hG5o8kLCuMwsvEkmuSogG
oYqVbeGP5KjxFbj6Dice7GfVbfPIbHQ6GCmeNTydRVwvdx1JIaTW3DpwfxxYqSR+LECk1ruT3trC
tHf6PpsSWZB4LGhyTpXgSDYuHnSXvIkohGMH5WI+EfLrlBwFkQscKni7z1QU7dphcDIQwcFxAMWH
/407VziEkEntfQpUOPrabD1yLL/NeOMc0cd8Uz6wgXFdDVf9Mp3q+MdlTBWPrnt5xyQjpV0lSrTJ
3fF/zb+4yi8vzxqURD2zc6TFpITD0DSlK+KP1FPBGxZ17V+3o+HETfuccv16YewT0hTsSuFUmlP7
fG35DIOU+y8TPMn7FlZAxgR62L1BYJR5PYyHTXa2NFjZk3Z8SLkmm/ZiKJjtd1shiR98eCPSxlTT
HZW8ndT6YReQCx4CgQs1SM7QEyHtOASq3wMDzSATVVYZoFz33YeG8A+j+BNz89yuDrgVA77HREqn
pOza8qCTHTxCskcKn9CFktbEMD8bsX5bLNhhMMd1JfqhdmLFS7mMM9U5PvP2rnNnGp86yTSF8E0Y
vdMPrrCjrQ4Uaw1yLi4TU4euFzklKOFpuZO5g6VruJfioRcNRT0GuxhqQxhYFbU1lP/Pn6SCAjYK
5o2IXmxMLOUQ1oObS/8EhJQGfacBgqxniyfyrQtxfq7dqq+bq+G/acU9zKHUU3JUNQT1KSo/Jt1e
s9Zl0mhs5wE0DOJr2Jsa61Ituz7yD/guLd5S7yob8fA+PEG8LwWyaNLrNQ5IKXVPUrlgukfa+gCi
7MshiUmGeIojTBTyXgPTxxAU0arBubXXCRVdxoGjVuHCFp4b9fCj38RP/5C26oohSkt8TaL9kKo/
RrpePbyAJUJBnFyxtXA7cjawTIuVlFvVnmZ2ka2kx/Ei5OneIirvm4dc7+GOOBbYI/69nwlqdqs7
6NSe9umKYFZ8SRFLwvaFT54rCNwsZZmXmTH+mhTjXe0ssbvpy1ob+/3VqEXbfmT5Kg42vv2s1xOp
z0Bedu7GAAHBKKG8AuKPHX5BOki/rFpKYiGyWTi8oCCTv3a0np10J65DVzNQ5YrRwzZ6+qdf1hhC
OtXMRFZU0F+8DzzHONJSdUVWAFEuucIrZbC+P1drbV/8ta9w5kOZh04O5+N5P9P2NWP04vJRDfVV
j5kQOezRHnxptjwoFJDo/2Gl7I4qE4kggdpnTDX4n4oCfshsw6pPGsupZvsRDhAw0UTJwkG2/d05
HzLZRhXlBG+ENvdoWIHnjT7XN9yausr68CjV+36AtXfl10Khxa1/a9vu4Dhm6ne+3Qjrd9ihVLEp
uKVXlucY3aiALqLVcMHjsrjIySZ+6bLqSFAHfyje8ebmocBsn4/9I+Awacp88gI+5/wUxuoTN4L5
y1InSU5GiVRn3saFcwo9czmMyor5MI2ezVZ67/JZvRKpPj0eB8Ge+rAf2yiLMy9L76CX7+E67Tew
tuPEdH/c9ir6PYmHmf3dwpJKDVoZt5oXdocogfsyvtr1gUNr0qoPKA+wiamazeIu24E6gB7FHoND
EgJfSoknCnv15whyeUihUvp3csCKDzRcpYRdE6PDwJPg2c6E4n42YkjxVE1Iv8gaAYDfMvuHW7Mt
FJucK5fofBba99rwex40G43eoAoOCc3rGPmnF7RLlG1jjs+YAYnDe6svlzZWxlCb5jKlB4nrkm9i
RgJQXRuGR8cSzSRUCaDlbSkU+YZF3bDLuzpirBqxKvgU86JtT3YbFg3r/kujYm4nmD6rtSD0Urn2
4lNJTwa7OAOZ72p6J4DxFayD+Oi8tZZu00q6YTjt6ZHmulaPGpP0HAO6EHR3G+71tw5YVtHH2LCU
n9rgwglyB8Y+cdbASxytHsZNaD2O9uEq+O0OaczPoYfUZZHEMX0nBjhxe1icoFgYwnIpupuBQ0bh
qAGMyVqJcTdKtOnHbKowAHVPwsLF8l13KQpl15andFkaiKG2vEacf4gClPn+00UltcmC7uHlBAJ0
CbUfYPxJkWl8Tr/WjdvFXVoivJoLQfbM9NksvlNFrcrOq4pHxAWWmlD5MBhgnR1UEbjAsM0WR9YG
AgmvXcf+NKjTUg14PCiE3NpPRcmKCX0jsHaOYoO35EDQ0iDeUyRin1ZDhRqOLUXpyAfwty3ukWN9
PdUnl0Wkd0NX0AWL6q2FaTTn0We7FMGzbUm5ELMiVfgebw6s98tjs6PeuloA9lGpY+n/AixuCMuX
Wwr3hwvuO/PBd0WtZAWTlojh0QLyCUIKr6R+BSYx+BnzyXsv3km0k4pvryEo7Kknzx6bcVs8fE/w
zWvuDMyZzBUZYl+eYGK0pjURTSwJ0PUs2JZJOdM0eWk3odlZyp9He/dnrWCiGjn8kKDYo0y7x2cU
rfmWgZrmGRl3JaxJGvXWj2z9EaSpjjxXVqpq9zY/fATiA9CLPE4m3RtsA5cpNYsAmdsm9gTWyK2t
aQAG7K3ohbB8AMRJMjnJUPO4hEwJhETBmgV9FLrUC/JnxElG0UzZZYfCR9Qtu/CZjBGl/fZp751L
7/z4xuwD9j6QlriMNT6FLFJ318HYxZO1yTIsFCdZN5/SWBGq8Q6H5aDLZal2aIRAaZkkil6lFsiX
uAj9Jgj88sLNPzH3Q9yNJjfDynLugB+Jm/qAzCPX+HMusjVDQv7Ivcezg8zmDqyFCUBte9jpizGv
N699bYRYYfhIXsv6iJ+PwkaveXAUzcIeYaLUf25HruNOdSAW+yOHTz43uqYeeYOBpTa7lsg2PQPh
gNmOh5eRKVahQjsNbS2ijBesaWG3JOk+cUVgAMyrz+r+bV3rVVBd7twYh24MexKDzC+0f0hrsNBK
v/bWRQ7cL7HhUXeBfExotFuXYr0YYHnXAD2O0iZUlncutMJRohdYqUHpKawZU5lyO6XPO53Xd91r
OebxKIRKw8uzADGELkR71prIhbA0O6hnKb05TxwI6GovFCwH/eM5o2CknF7/OMhPGEOxD/3ArQMb
6dCfHc2royeDBcu5wm7/a4bDj1/Aq7itpsch5QYw1fIdnWP3NNTCLQk1CtWpn/EwemLRSfznm4Aa
IsjO1VcwDVM+TXnameRHag74Muybhv3QgIzNztAM1EoxBLpetPjzJ2DFbgygCkvGweAUtIn8QwBT
hfb1Qy0ZiiS+6SNvazho3NL/6ffTuCyal5wz/XklAdzwoQwSp0dDBtsQckhWOuAOEYjiV0+5itOE
tZTkxMUEEzXpsIVmh0Opv4Ey+tGUXxQNubrzfkzn/XrCaI4xNZex7SPR8bx9lEdM13M00UHRAUR0
ejeE1plhAaZtl0j7iZWgxMcvIppOucD+FONTGYlGdMy/rnJFxbRunwN/EhbEqF6gcl+OjWmyagtC
QqRO8enNnDHkoQCnXIl0YQadhV/TqEbMkx/qBricNcyVNHdPORAJ01r9xzSybzuNVohft6Gg+8wv
uKlj+BSXwlDKZmm8pfzeIjru94Wx5SvgZ1UkBoNcrYeWPO4Q5dP69cJ+deKuhiRh4SiF2NyJSo8l
mhgCuqJBGqLHSF60ilWhPq2YaMb/PZ4bgWT/d0jFjBoo4Qn1gymZVCnmT4n+gkfqP7VcH1gTKH4W
fC7qBqgAK6pyq/4ui+dNTX0k7wss770yS4TVbUJ2qliFuJHpzOdZJ++LNwZJg9mrMJ4gbFwUFgiz
p7bc4/W2sUM9q6LVL+ANbMiD+rDu1Zy2OndcEGkY4fA36uEbUWMdmOC2l4Ou5VRC5L1DunOaKTE4
sWPLFoIbabpom4m+gPI7d4meRhgWnKR+86V4JFuDD/VfN0Y6OEuUguSLccUfW1XaUnE1HIMhJshq
1F1H+w/wQCkEFO+lRm6qknf4PKKR+1mTKfQckOLTMrF97PA/kwK9PtPCkZhjMkPB/6he6KN0KFeh
9lBoB+0PlXLwVvUkYhdRA3c8tuWNbYwSpBLIEir+7ps2rBtekAWVEE06eCIpBOVldTtZJyyfdc9f
Ltp7DE6+ZN3WMH0vj/Z2fCjbnIL6lWqfF0nf4Rl4jFa+8xfq7Z7ws2GzFBiE+4Nn5tzJzKaBeegV
nHYDA7dRX8i6c6cJ6yqEbd0PtRw4UkVLhxd0b0T5jHyEUQocn9ek6YTJjrm/+PQrwrGtEYFWmZFu
Q6fjGkRqxo/zOio08G3+ub3wXSy3x3wG3PsotAzF0/ENW0cY7Fn/jPQG4B9nvvFu2Q7Dbly6498D
4hH0yfEPk4En70Rq9MQwpq90JR1KPLxnBiM/mXVW2F6PNwNHYLNxlEhzzVrmY/O//qCBgQo94eom
nuPDVZ4T1ehyJt79NKi58VZSZAxMvE8/UkCAp9gjAFmDYcZknjTHtPFJuKAsQ0wtHQeVTDTSo4zr
NSiga08Ybz2p90DzEEcvi7QnTDel7wbKbEqUvstTULBbfvS28PGmChW79ux9OQP8hP9si+C9GuyN
0hN2WjT9pHa4YZFpS5ntUoUw442FXxayCyUg3BS/H/q0HAhKAInwqNDRFIXzTf6q3qKGdzYbjtPY
fKM9VD46mXgJEUku7pxWmhMmPYUX7k/ULm8nWMiaeoq4Qvu/lmUCY9b/hRBKAipDxxaDbiHp/IfV
MzFJL3mxlTbqzZc2Wz6JYZ44eoji2WmbWbwPTkjhJEHTrZqYbjVjwu6t7yxwDO5ftaKl1Ag8ZFt8
5lwi3Ko77Xr406t97LJ1wNBUUMEpWOlmZ1cRU5qaL3rVRX2JUtOg+Qb97HuK0qrrPrPQY1hBHb/I
KPEzqwxAz02XdZTlMcdtb31k84awazbqSZy87ImXJFiTgGQZKnQhZpL1f4DvcDPi0Wpau7Mttpe/
Wrt4BqZE3OP/pW+1m36jJ/ICCzTmqVtfj/unTuMraUAHfwRLPu1wxxYWOF4blhfkyqiDisJ8UWas
O+dVIFH40l1wJtLjjx0I6r4UY0rhUflyuTcU5EpA+Q4QuLawPIgQRriWSqgkJ8MeFWu0H6YHcZBa
8UnwwOSoL9keCgYG2pjNcIPZRWqPvTETOkiHjTX/XOq52S56ypnh44KNyXYVmGtS2Bzs1uv5z2ap
RQNqO/2g+CpOBW52LO8JSnLvgO755wtOBkBxgokKB2WDAOH/W2txRZvPmKFbRGrjHdtwdTmK7n1s
iGbZPv96zFJlrSUNze1DGrskpQArhYl2gXvayYx2qpOwokUjWFiGMI5XRLsCr/4ZJcsZEsO6x/LL
HJVIsM/qKf5iACXGP1uTedb80javh8YX/coAU/3uO09W5OoW33mRowQ7ELrdJWQBT0tXkD0DHu6v
192JSUp0tyo2BmQusr3h0hNnUkZ0NZLDQ3bBELVVbFeYqzI5U/lB4NQbhnhg9hO5BmtFwNbFZGF4
Bmr5oQqDsS05ES3fZpA3BE4CkJVo4P9nlO2jU+nJLjYlcPuik833VNu1JAHSMvVMsh6tMNSHAF76
3nvI5KTVdtphRAuOy+7jdHw4ydg2+7Iwxp+3rFeb3ObuPzUmpj0UmrkO4rh2d9rBcxgYNUYMpVX9
G2K6VyOI6nq/YBEkAdG1/dTPQVXAqAsve2MvJTcAhbg47Wsdyhmk5ryEOEyvOfG9WONo/zWiOWbV
hiHHDkW6x/jBwKaCChpGbY3FpF7JDre/k6maQPVN5wFrBQG7VXR494DTBs+pa4Bk0hqG/2aSM0fx
cg1WKQUjJPnxejEv/4zr6d6ns8dT3RJiuYwa4sft4ADnPXRSvEj99OcQ1CvWK8yerOzI+sSh9USc
PWjJAUjWJSMzYwzJmeInpsagRgm9knBwyYK6Wd4kwv/vhCgDULjN32SH8dQoKmoTfEc9tRFH3+Hi
bXULKwdJBkvqpRlq6Hzm0Aw+p+4ncX5EGP7LalrFiIu58vZT5BRhAi70xioKA03nCXRGpKOlwMdk
F9CV5BGb1hSwc3clmJGYezS67pNYPN4vTckLnce1VkhUWtTd3HpDQBzY+cAGFXRpmLjbVahiT3uS
m96RjI+i6MQgxmCt52BK/8uh3D0XhfLpMh1JjDCUCYshOs0jDth/X7u4J075dd9rOQVGvzOYq7yu
xEwCn0mJmzcxgVFaiE75qxmEOucKKyeIUE/GaDmf0wDXcJF71dotO+0ErH7E1Q+LMUepyZm3BQyS
cWSKZ234cb8spAMw96uEWQx46HJyDEPJtrJQen7YWoB01xGdNVCnCc0oQgp6QifHsXWz/Bl7TiV7
7auCGXxGpFWOV+stTi6A1Sz5GdeYAsKewwR6giQLb5PnC5ey4apGIFi/3INK7KP4yzoMuDFkd6zK
MKaEj0YgK+wEMGtYC5DXny86JutTnQTwYXN7G0tJHEMqZAWZrZhHyxVW03vsq/j4VrA1gMx8Nfuf
x6Bk+akOOADdlroMkHQ99JIjwJoOpit2tIJmTbUuekuoF7XTuOok9WeldULw1DiTMNUqv0NPHfj5
BcUUH6YjoUfHqyC6v8IJyvKqS5Xzu0kP4GFhR7Yx0poa18KM9JqxMIU6toglHVF6poqE+ATXpNuA
dGGBiomB4IB5zbLKjT3Wl2FeyE5KCBjMwFw5FMI8NyZ0mO0/p9sCfaUM6XYut+muZv1dMeG/EeCP
Aych4V/b3LYS1sZVUDK+ZVRe3CocR9BUucZ6OKQwvSTjyXPxZVvBFE7v1OpDmynxRkoe/9tEq05j
QRJrZ7PGNAKox+RUdlslKIshVWVHfu4OaPaK1uvPxZLQhhlucMVIaBmoru8kCN0duM04gvJUqdaO
F5oXmcSfNmXIj5S1z36S+pvsJjj+AHlWlpmsePO/BuKiLQfc+P8j0aFTVA/w7WGthWGEM/5hwcVK
/hEoPn/C6qjyiCG5QRhFiD4lHTL8HK8E54a9a+NtN6Gh7vby8xMYsFwFRZgQEGuDnMYyGf1/OwBA
uPGX3qauIHxv4XuKjJbko+t69k0GyyCO5EyMHUr1aASY/dgLypKw86jc0SOnW5DGkDmugIReSG16
5+gFablRyuBd+D07u6VW97PXbrGrMEAaXFdhKze9Iu+xK/zwieXfr3iKaFhm9uyy1df3/AAuPopm
8z6pdaHhvg1SHYIThK5b/DdbAakYw54gTTx47xWXu3yC+BzbEP6mPd5h9lrQK8ni2sfBHVZ9z3md
ie22pF3FuKA3qzBjYCQFk7ejlpTgHpnrmJlp5OtLbxA3QJGnwLiWo5POQgJWc1yYU1eHmwPkxA0=
`protect end_protected
