-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
3HGJiJDkDOVmgEPUCUUt6E7lb3r3BLUujWCEoUVqN9+rxHkAUg42/tQK4vl4VaB0
yfCnqq8BT+CZrW5AtDQNB+Qas/4GLa5TiB0UXJwhUR+fh820FhyB1lMbprvzoTlm
uor1xfoBPLpbMPoBWGr6mD7joSWlZODOe3SxpO9vyO8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 29760)
`protect data_block
zJVtzpUnor8FqJIdT0tLYvQuRwlOB26RJdAXQpuQhKEdG+aGgdRbSbThbx0uPlCq
p2Q1o9eE96KBaE82oIxOMGrgSnwDcIbGZIuOkprnD/IesHY0FYFKkr3ns+n4PZ/j
9qmeaDZihvIkUzkOdOalpXaVimZKHPj4VuXY/IEnTLmKa6W1Et+cC+XXpL/9z92B
t6nNAPl260HZ38fN4cNENQ7bs2xpEvOxsoupr6MXh/M7FEdxWyYEq6oLbN3rxDXX
Pk4CFozW0t0uILuXL66eFmpsslFsv67NkE5qHUeMbEH2vCE3KGBUuxA4yaQtKur0
MXGTPsWsi+5Tk0gS6nZeAe4eyrAYuicuR+eOAYXkd/VPGfrewrhBiK1XTWNNQzlx
5D2fSGWkwLxe4VMPboXO1HTmzGcRbSXQIjjM5NRYtITu59UK5zHslcKfQs5GUMou
xVTIEDVooHNHG+0uiULq93JLZQy6z6dI/SE82qpkYHFxLrayVKT50CZOUkfhIKEJ
SlUviRNZ1Ndln9l4irbjbf85hMA4aHM+nX+l9gV1k6mGUsYT+Qdh4p6TO/T46wGF
ME3AzFvc+7jHLV60rTDffi0X+E09fMyM9oe9PMCzZYlJPgiweTrlNXsiW+ztHzOR
Dm209ETijYYBtABCEFMLE6bxDKV/FvoQF8SrqyDYpvU0vU0bR8Jus1TxRDFDHyqV
D3h9Eb36sCN5romnD5VHtSSj2evnIjh0LtLji+1/629MTCax0oHmWccRzFoLav8N
h6PlSPw0AipqUcz5GoJBwtovudUPx+qqeAqONZ6toJMHwq+VJK//IXq0R/hoWLJR
xMW0SWdB+tc8i5WrawP8EO+rtDsfxIS0NJciUijEx+jFj+vT+pd586lBBIjtOwSe
6rShhJ4zYHXlNJftgjholDNtvUZ2wEu9eSQfXWUsL0qbLBCIHHusmCQdGLVXCn8t
q0UhbWLLAWie1+6QIdmTshJIt9mAB+UOEfcJucA4LZj1Y/ce/gGLgqh9eDXeM1ti
QRi4DTDkj1FI59gipZZF5BCDMIs6zuKPb3xgt54iMUbxeNDK2yXnNxHSga6T8Ya1
a5r89RwPs+qkM8Cdipf4wHoqByaS899RDcqY/xf9sl3b6F1csn5CefNLBlkAoDTB
paGkryUqkJXnGhmjCX1iogJyS2gHD5aPHfpSIMw8fM6wGhBRnHn5h3KkkqyO2Y5u
cBpZnaZiUWUKFepvzskq1lXSFEGHaklo/0x4Rbgl9icS2x+qOoix/OEjlDP/0+zB
cMEK/OLujEk9cyxHNBO4aJitMrPB6+RwIHXwSU8SRp3mjSmdbxQ3Ma7Fv5InhINh
sMBWDUkn5w1DoJnT1QEQl8AKxgaNof+jMtW7Mm++1JU1rC20rI9pI33EX3ip2hf9
YiegJwKLLa8MCXDEog7/gD3g3u4E0KAp7WRRYpYeDcDzfnVxfZXWR0VMPKlFmkzK
jxF0t356YQLPLIeIe8Z4e2ZUn7c7M8c5peTqiPlEE9S/ctI3cFHFqWmX6WxFYIgL
x+0K6Tg2S5SwtAYqF8AHFh2bd0R1rlcohFMH4zAiiaT9eLQL3f3LVvSYXxy5YZqs
Hw3He5YDjLWNhj0Rc3ChWb2AXqXyp6lThFDCKYNUvSPq7rMZ1n45MjpwmDCwx2df
NMXdcuPC8ujgGX2nM1xLzHS721ro5hJ3yTJfJ+R6ApBe1SHJBtXhGOEscvgYyv/T
+yezc7u2rxkINMKkeL38PgA6hRS3CtWBlJTwpLG4d7e374KMpcTV1fTZoMeLGx6x
lOg624+4qeCjvm7zPaH2oe70HrhKe71LqQ/Erv/H0ZibWVwgcYn8+LEnfbH3hZgo
o25TnJrsbyRM/r9mlgDi6Pnrfbgv1SCV0h0kY9CmNFP+OfsmlzXzre4q4L12Ckpf
LcN0iFAX1hauhX8gMZOaNP393tMwxAYFmvTdza6dYtdAwXdK8lmxZBWwfYTVRhr2
9lpP86+mn7U51UnGmgoUC9buKZuyFtaAkGzh2FFZtaIAs0ilEnpxDWl5uzS/7K0S
xhbYVgXt/UP+6fzhK9F/m/y3a/XJyNhQV9X9sOnfii+F0ucKjrcHTti6hvzhzwjK
8M1SlUMiq3mbtC3faAuxvGBpESGnK3fjO/37UNrK5T4MFyG5xl2/7eEPVZUBf+J1
BXL0nLyvc2DY6HmWaEv+jFLxUM/0eSKh4s0yFzmQXtoT/CsgImHDy0FCBgggtVob
68JAX4j1eREMM+k/Q+7F6BbUqmB9uYOeXsdLQc+zi3ZS0qpWArieKWiIdW1nSNaV
+SeIY9oTf/9Q+2GDXUAGlSJuFfvmIB8wd62LHPx14FA7Tqpu8PZjrAytbPrt6wUT
yRUaNobLW8yMv9bKHck3J+C2tYIyYMt9rrxWd2pT0YC5wbqCP3soRTvxCFOlhXTN
WpLHCHiEL24No4kYgrrVmzDmpGTxDb2XiEifRssQwmgkOs3C38cdnyfLTLdscTGK
Sr7T0coPjQVje9GqfvDAkA4nEm3Yt+nT0WjbGdRM2vA4Ptqz7NuG/2ElRhYR3dD+
Xy/gnUkfPxVJfFrUQhOmGQsUqieiLPPf8nqLeW9GLoMGHny3Fy9Ht7GcJYRTc2/o
elB2ZGBqoBPvuA31uHjvCAtYEBvnuRe4M40Q+xXey3cYrYfJSX7kwCn3rAO4QWFN
QAZxvUAY+keyYAP0bVgMo33mQbRgYKBcKSTK5jn6JHGWKz1X5LzT6cxemCjIKb3D
vBh4Kuc52YhMORC0d2J+LBIgdpAggB/xQfJ7dYFfQ3Sy1hui+vNXBA1kVQIJit/b
a+GOoP0nSGY4qcjyKnp97P0u4tH5qt5DRknbxC25t/nzWBDd1c6b8LMFk50A/vp2
fzbyQ+J1LWuHEY4f8GkOPb6K11YNQlyJPE6xPR4rR7Z2JGOPsM0wlqyndM4jVHdG
dPItKZTJcm5OBi7MiXX5ZWGEchuFWioki72XHqzVKcftTJrMPKsYGQsz452W56CC
kzZ/b20rSfgsHfpB1adaLntRmDQ+a/5L2nYA4fUIEwYUnjfS09oGxCpvZD1mtOq0
PTd3mutokvKGtmjxvUsmqcpftDyp/A2gvQtqwJ6c9y90xN64vVUFOVFYc4UJ1qkT
7lODeriRy26E1TJoqFGZpXW3zCZKdXh464Hfo/t6Dp4lCfJbVH66cGeNsG/DgPKf
ZpFw1Eznc2tQrrAsDZP9NLt1R3OqLZfG2bw3w6dZHctF57HLXye9t9HqsbRvoDSF
qx+KIdN6xv9HSdSDOLbu+oGLYGlc/ASv+TNarFTxVgucSvSICLz3pdCES2KWWGPp
E4psY9Ut8ZlDbslJKm/0drJEkwV90RKdkDaY/xIE+4RUd8gHg2ZsKeba+Mf4ZYnv
4FRaWD/DohF9BhPSDOFXoGm4hYdGANlRQoki7Tu2C/8fpgcDUulNf0CJeL120rHh
ns7yYP0hEuv4AIrs3/UsnmGn11RVJuVIwlXdC357fqlRFj9288ISpDGyG3Pwn6c9
d0xDi8SmRk1PLePDHrI08RSJeN+Ooth6XUx6sq440t+Nktk7vfG+LZFIIBJjbDMu
kK5OEFgROQuDK6wbTB3WATJHEVGkmJeDI+x9PR0mm8IAhqGnjjFSJqzkQ9irC/bT
8QlvIGG8qukWPme7YHi2dhVwoxRdk+bDf/x5yjvmVFsOqsgOlC+/pbJKd2p3NDpN
bFFy1qChHlZu1jQCAM8BzfBantnOXNedra5RRJVRUvazarKAY9gwyJCjohSoc2hX
JP6J7QBd8gq9VZuFvmTSEV2S68CXQtbK6oAm2OGsu0+udjFIcSxkq7yPIexBTdeK
VKczErFvJCPSAPJwaXWAfkNiZDRZMHFsX5cpCTy35XBjDqLig+Jf/WE1H+xkAaWB
TOLbogl7b97XHPPkXsGU/MKozR24Tw3/9GWBWkaTifmyGTm11ypDIwclTM4+bSFV
I9yryWUXrs78Ava3m6Oy8KwLWTUr+aPUDrUESUjgJ/nk0eNqBOGhYehJmLxeyLtk
7eGGpnkkM5tOp7hBSD4hod/DRNpqXHf47ASZWf3W0UsRwayn4OJV/8aO4mOnwThj
9o0ZNYvnW6BAyoQELE44ipWlfSoj+Mf/I4wntd1/yYGyW10cLB48/tRGG8Zk78We
NSrVFAISfEpjECDNsNyCrCXWiYl2z+QNmVQ1pEiwMwJgQeuFekCvUnjco1ry4LMf
ZXGK8el145dUjlTJED3+zdJJ+soMG3yBRfkSuDQVrRvRXD4Y69by0otveBq8L/Sq
LMv0UoG2yJg6uU4Ln1rV32Dp/ooWgMTiLoRp3uCTdDPn9WOWRDyKKyQ5UXVSYdES
rjAUOhLXJn7NwNl7v/dYCgJeGYpjoqxldGD7SJJNhhN5Ewwcz5C38rBVaV/ykegR
JdfeqjZzHotrpk7tpXonQODSjDXPOX+bim6enM4vA1jbeB0MmLIBjp7nIQtT/1Sc
oqp5JYOpzyEo9F94K/pZgWZSurYRjXjQD6QpSXva6sXAPqFunEeoFTv9+fdrY815
L2QWKxyV/Lj9Ml1vWqz4PomKl5MgqbcOALebRyDlVx4DoJ391dD4N2wG28RVUrpZ
ayu+UkahyF5W+yp40DjgWQGPH6U49Sxo6lFlV5Xm/EfjbKSHO2HLYzZnQn9QXzkj
UKJeVfDIEyX+Eolj0B1mOpg4pZ0f8TR3ciCqh+zrsrPD863eD3i5DKBVdniD8Ogz
/rBTT+2RjH3pcsesJ8ylcFowt3qEeiuQT8tcdWVeVIA7ajv87tLL2xfomvIbBloe
V3j5gMehnvaX85K2aKly3d9SYrCq08rMricYHPTovuYw+oWsDuxjuSmSUk6+i9Ur
oPvuA1OqpF9ldrpH1lwcwpKP57fHswr0uL0wKKpdjiTfQvaKh4PO3XvF46XdRi+3
B3Tu9Zc38YQ1RIYHEYxY1bW3720gBEDRXS08/TK55zvnPX9vZf8VTAi9ZL8A+ZXU
mYs+eHjQER8h85DLfuP3u2I/JSUAD+BnHOe4D2dBdWl868NDd+VrSCZfboRsC7c2
VC7ffj5zJ/36/pFhiya6OIj+NlKdgJGJYmHEzYuEyWu6MWtnUM+3N4ANvApHBwSH
k43bkFmTUMeu4bEl1yIAwVNxicImbDdhfxkjjh8xq+l+hthAoIT1S+6/yhANXxvg
PWGcPlf050+Y9YULa6u4HDdGAFxYz3ce8jDEOxILzZJ1G5aoTRETEt1OMmvEYIyR
I+MGOZOnnNsLChYAq6WdF+SPYcG/38PQlFehVtLZCDeF6cypQMmLHIxPmHj4Fkp0
Noqxyb2UB9YAFfqWfFwog8lGmctmA+HaEvXXTDIFEJ813BEir3Cl6zzTCfGouuCJ
rRC27GUyPwedk/VBf5k6GOm+NyvtPrus5QnfZFz1R4Ve8RdcdfbWVjowi7hxXFOg
ZJIoN8SiilGNV+C9pnaWL51pnxGpxnC0ujJfiChVVhgM46JhAx/GwQ1Yasu5Budc
hSnsaYte16BARqnQWOtL8BoeXhbyTcbcex8C9SvCro1o8EDgMo+yBj1BhQmnZjYD
azFdY4Nrxjjs7NDmD8SpmGDpRMESxgMah5Z9QvgjOcrAc6GdNGVhmrcrtTHmxQcI
FyfQi9rSJXbGayqA4spndGIb455Uh8Yi+B237upS2uBPKAlUjEnifwFH+sd7+47i
SnFu+6+cUYLynTtBp5zn3sk8ozEC901DzXwmip97tosFe/CwQQ3g7nbgU9xLiIcl
7uVBMoRfOxntrV7TLJWBRA/FWb5RSejdpgUw5Ul123mKNobpX0CNNxIoHQlDRn/9
q9GcCAwZU4DdYFLIIum5cCuQMo8sy1a8sXHmnBchWUhMUk6srhbJgsvkHhRqC2pp
nRton5JxGDhBKys65iR6lPuvcejtLDz7ToQTSMepzvxDMH5QXH4nW9c4mQfcSxH8
lTnB7kj3lmhZSnyaC8RN4yKMg0+CjIJVxyxFpCTvgIQFM+s81RvI79C4/+5sx8JQ
S0YrdPmI5d5okr4sXa9oOj5Cpgp+qzPJoKussHZJ130Ii8i8s+7ITX16Se0YgVck
MVcl0wx3ZKdEfhJ8tR+ThjYt0fsb+Aq1x+DedvATwMmAIPUI0W9aoLqS2aBj32CT
jxJTJBJ8BDgd8udMJDcH/Hh8FT0ZTQt/mx4UNYKyd9Go7COripIGdo9nV8zm5lpS
Tlj4J1MsviTn5HigcFHL7gKbzT6S9myXmHUPdgEvuKTQRxt89XtMDQaUjf+2+CY4
ojM2WGB616k6kyRd0SOfhvsIEfzoqoPw+LtCpTe9OzZsRw0LFRbhotRyRKGJK4MA
+w/7magbOBzy8XrbRii9lvo1qX3Ae3MNPwLT5XNTkZ1R8UF527ROEmUs0LY8iv1G
Uj6etBr4JjmBY8a1tk3t+KkbKwmZIQztcN8rpY2/5s2DGcPZaCSwjwAz3sXY7V2g
qlay79t+kUUmnURBG9aat8lL/Vm7PoCAwiSLFicj7O3vyh48dfJzNzNXZUBin++E
n49YadKQo1zbtCLxY676uoIbB8XiY1HNFZp35BhV6XkLTBBup08cZXqnMZEGBGN0
dNsMIaZYz04ArDKKngOkb8ry13c4IY4lgqcFybNvq+1MA92J8+Hwgd48sBiIGrSh
+B0JrIgjOQpxINNJ40HAcKs5mlo6f/naouzupIcbnsa5YpIusURzXJTB4AHWAi0K
AigSKhjR+3gHxHDbGNJcV2uwXNKA6GR/GSkpj1HSptgNcKmKjmMvkxMFmxiA7K0w
RRFwEoeRn9IjE1TeD08Po9bEhiMIgRcAVNrk3s/m6fk0TTgOlknOkUmQQNQNJaEY
qDt/gvPrwbzTQq9hAx7JQCnINwSUQrt/DV/6TK6Kafkc84a/Y/L8mz90u0PoP4dN
2WSqQpaQEWFXgOfB9yprBvkopM4sTe74wRFgL+PNwMpOrzHbtAT9ozjK9LlZijVX
mRJO92sS4Od1m6V8sP5xGC5R4pZ4wmm5yFjdnieduFBtoW/8zoumNR5veaX+Ad7g
QeWLeUsPVqoTTvMlv3WPr1pYt5T/k4VVRKchvz44tQjkzZJrKIUzo3OBnazu0s3d
ccn3BHfmMzOlOxS43330WWkHk5AaWqa9OwUMHYRwgBSnH6UcqzMsMwXq0pn+aGsf
O0SNykzInVVtVP3kSLCARBGIKJxXoJ1WsZ7g6OJrt5k+3tkRzlZMekCWO/VooE54
NdZzm+YI1Wuy1z7mj/q/Mx3JLY+bcdHV2NxhjxkRZlwa/lM/BsvmayhlIUqooYCa
zb6BVYGa3c4CQ4ZHx4tinH5BuU9XlhyEdgYrcJ3v38tVK0ql2KdH+8BUel9cyEb2
MiUY1bv7RUH/0foG81DSKOikfYQ/YVyZ4/k42CIqnuhkn5xp1cebO1OuWM3TW5mv
inmTIquY/Ckw5wKEAFKnUsg2b0d+U6hRBu0eOoRh4KwU73kpxQJZIGh+yNAa3k8h
sw7r7M747ZL8VaK24A+fy0P8dKMiQIn+JtfWqWgaCakZpcChpZJpf1IgfMVOCHJF
Rx1BiYpk7Tr1Ijgg68NA3TB5zuSgSDXddBloeue7xesFo1I58oVtAtVAsjiSDxYQ
b8ywkg/Nr1DV8c/QuEF6K6rxi3F8f6niV/0OcphEUxjPpUZoP62/xrwphi9TijAO
mFPokgylo2t0mf0FhwYmtrnJ3CpNQxj+NBxxYHR+GCDXmKdvlBmpvwXkAvQWP8su
pjO+yfsKXq3ufOYyQBvnxHChDyWU0VC+xxWZL1i18n/A9UfrM0JdXNvzhsaxLBL/
30Gy2v9x/j7feHsoG5Rpxen+GDc1glcKv55jndvVGQ8gFZ6/NUS4sEfon3dcp6z/
1os9miv11fGxbQ9m9E58zE8KXq1tS5orih9F249BY3a1kdn5ar7PLXH7v6DqIYFM
TaOUvo40ShEDzTmXKN0WMn50rPEL8g7K8954w9I0YOOpTeC8vUrfvF4rgDhPpU/b
Uuf5HfozIkPoGdx9DyQp/pcVI4NVkvuI+d8Kz18uihxbCJa56UrpyIofSPOJcu6x
qj7hPuzf5lmHw0Q80wI+egtQY021DeY9SfUYSKO4YSwTqZRleHWRKb+2xbI00TMo
OwYpUU1kiSG52Tj+1VeUTzOMesNXi8LF50ouEeKEEnbCTUkNDTO/m5kO1y/AGND1
cK03wVIKwqPX7+cAuULaA9hXp8IG6D4P8AAUQjvGUMZesDrMzk9cbjYWQGFEQzQO
5kphuw3LFMwfC5EgL4oztxh0kdqurt2lJ/+QAe37aahC5fNDpJVfJetzbdyb3aw8
tm6MftxDdgFFQoepywo4m0me/YB65UgYxk2UQF1P7cFTA1oEyc3U6BOaqqCb2EjT
Lnbuzv4rrBb0dFaK2+AndUtWp4F17MJ489DCyVJ/RXFmbIDQje/IP2P3W9Mgs6Ic
WQdqsj+7TBwLGmq6QemFuGvTuJZpfK+B7figPWm7ztgaexHuQ7gLs6PnMHzeBC/B
u704+7GNMFU/yQvVYye2yMhQDZarjCnuTOvshihisGtw2OHl7tywfTXQTFbfyBeJ
zeMSd37wabH5zjDBeuVrADYeXSwMK6fd7yBeEdOkRuFjdYxTsTE0bDPKBfLVutHT
wNeuCw9zFxrGdchmJ6Gg2eaT8gZ6e90a3qL7MjQOuouvIDYUodEJdP4a48qm14D2
hMtxvMHbf33Gsx1R8ZCc0cZW9IOzTNEkC5N2VcaXOTlCYj00lfSDW4+vtB+MTif3
xSJC6EEpfpCnhqhG/P9f9SzUcoa01jae65CuGqvSYgX7oXWS3NzqNhXt9/hErEIT
EUifDJ1KsnRgVpMqAUalrTpL+h/PwQMGtPrPvxrKYn45AkKE85DXOKC+wlajjn6X
iA04Dq78Yw20q7csvWlZYKpGl1EYPahFx2asaFij+hi8LevVUxsj8g3B01aSo/PE
r81bOqZ6R9AeTDo286LUziVXXabeQbQsYclsi5GF5Q0XZBLOm6AWpLrpvR5siyJT
cz9mKU9NSHK9p1j7c85aQTDQkY/0xiIaFyvzA5daD+drKvL3cZugAP5GnO+8BfSV
Gpvt+HihgTLaq9kaP2NalacTZhEJcZ0FfEUDU+Vz60jj+BvNDiSh1WhpwAqsPrNj
3R3br8r4Yi7Kh02f8BTrsm3OHZkZ9wNj2hf4blDQF6wfDZ9Gs9gSyr0BtYof36Qt
mbkBkNxKgaJ9N3tfpihfwXc57tQxN2SmoNWEBAQhKFbjmwfdar/aXkEG+6tOzGrv
eBfx5bcqN2+Bsl5mkqZywCY0QYGG65z17MiPuuyolpNEdvxs5W6+eda85ZEjhfOl
kHeHhCK2ctka3wsfICNFL57oDS+QQi84X1sCBfQQd1F+omy85z0Ibkii045tmoHP
9z29IahhqiM8gMDPxfzNxiDfLFvV6dnxTKmGFyZfi+u2GRPETc3oy4md33GnQ56I
bV4W/bZ1dwEMcfdFgEAZyzhxb0LS5lPUD+PbiJR6U3QIz4LA6ZsQMGvo8JxUnyh+
lHOQcVXzc53ci9+5j5wp6IGdAliQ/7TEe6c7PGQLIJTXmVoJD0eP8X7TDtYD6p41
0jTwe93jw1LusDps4ZZWx1gZYd24bWk0VmAfSpJl2wRHI6uCiHi3+iHD/yKgxw4j
hrLo0topvn5VJPug1xdG6BcDQnXBLL877UoLmDTbh+ted03IICEBi+u6Q3pcDcSe
Zd677nQtWuuAU2EeVtRPAJSsE/RKvotagRv+nk8FTg192KYX7mPDoa4O3mNr+po5
ksKsJEssBQl6Qxu/M526z6CveTUeHMM5ChaIWXT4pdGmd2gl0DQ4LATTHvnulgm+
NS91x6ZYK3PSw0dFH/rGfskM2Apek5B5FCJhl/rYRV0HB8lZf7ZniYvoMaiPpmxH
Uygm0+aSO+9gKcMLP7Rik6gK2lLyzMxef/0F4TdVbjYXtgC0h//CyWc0gDvS3s17
mDrArkPF8LljrZmfatZ3dDQauw13LXAAz1X3Ytf1TCbh3kA4kThEQLC43WtQXlSJ
azK80gHhanojPeZk42Ud/YcHHHS0mYzbBHS7gMFVCj+StIXl3uVFzFu0lnCuXLry
2CTuktha5h6L54no2XlTCU0/u6YvQ4rZJdXUzmbngTAEw0/1lhieqY1QHXkHNFla
lJErFtR3DviwGLJnXW5gRsQsQDDgqbBODs8XAbpyKl9Bw9v1h/wkVL3txRrf/74B
ARHzJUdvRw0A2hpN9wkR9VyZZBS+dsAb5RPKmtQOOboo8ghEy+wciu5zSRmp7ZMZ
EfdMSWUNUIi2BdO9DboqJlGyILROprCe4M/Cx0tShhM8S8eE4yWsGTVV5Yq2adjm
V4RG8s4xBZTvnJw2RBMW+0pnxg8LADbo4E4Qr4408y3ZRVcyXF9rKXTG+Qf7M5T+
KowlrK7UZfJasM/q7THP2Edfd6KEsoNqyCieEYJZuN9+XKlIqAcI8CcNZKjgWyQA
zQqTU0ApaqhHBMdWpkmNDBUWXzUAr49vkn8rAPmZxUqbQYhXQ1URg0KVajlDzBRP
7Yer93BWxFiIEkGdQxaDBZUmtgpElIt/YGRFL9Yrgiz/gVDb25NFc2VhH7AXvFn3
BMVVplihr2Xk8o1RmTEMkEFn3iTdfdGVyaV1ytbyfXF1RBIlv2e8OpxDZvKBrH06
x3NOGseneM0tkaA5woCOKR0STjxsvoQ2Lrjt/uAh/kI0wGm7bERrXzVepgiavnYx
PnO1AQt61dXd58pTnRAbUkOwnzjMzhQOew1mZSnTrreMOY8trBa4PDDsKw75f2ny
H4bCuu+pEKciKfcOOnFohfEkt/s1/nFqL5ZNDGXqHmgUpUzY1ejzbLoxWYbo1ml/
izrQMhCVK3YD3BkWGPALqPG12eOvzZP5IbvES15nZtVL1F6XVGAtXWA335WzVTWe
MWI/m5Ie/nRcnMhOoWLqBANRllyd8jbHQyIbRbX40moeMAI2R4ibTr9q2QJl5uJ8
5JfaQOZWofwYq+25iqol4Oh47T+6l/YIx96nEd5buby+DskckKGcOden3uVWhp1U
mGVI7UR2/5H6Gwni9NW9OCh6/kCKkyuTFl9o2zu8OMYO7S3qAOr4ira+QVORHV9J
UwRIk8VkPd4jY3sYHuXIz/MfcxcH0os77FLxLiFsXg0ppwVygezNSduupm4P5Ylu
ZSr1m8w4hxaRKnhC/vy0FxH1FjDo0EN9L+E22OmhJSxDmDMv8JYYIoCOPFK+uqsk
5Du5t9qSAjrdYsexjyVee0bQAOxL6OyGLSB0SP7VsHyA5ibvt2j5tZ8vy/ccf4U/
dAX5ARN4ahkGFeKZ/q/EnOHo4o4/czKkg4JF7rqyowD3zfZ04uHHrpAVcHGTePVp
o/BhTPEK+04GoFCryjum4+aKpMvZ5ljyr+QejX4Qc2jTz6/6fxTO8HQ4nH/orYuO
i/4MBUqpId+mEDocdBosAvnxA9il6e3ge2l7U1Qadolson46T2uh31+rJKO5XFAu
KoYFrF746WFwPfRDXgoR5XyniLA6nMS1RjxpZMHyna9Qu9aBnt7EXBUdg9KYaXP6
mb+nnlVaVNz9anqyDiZKWmR/SBM8CmVEx0Y3BL6hWN7VUTdgnbUHkYKM8K6YlNV4
VxH3RRPVL0adVfzpEmk2hJdQsz9x/te/45T9t2f2TCWAQ0djR6MYrLrUXAfbh9F1
vhP9X0JaVmOK43NiMPYI4MK/l08Kl5PWs0P9CuuMgroZjP7Svs0BEu3K9jEYwCEF
bcMGg+q2Md1Hcg0vBTgH7I8eDeyqjH8E3EOZ4qFB6OnXVv/D8amKCQv027e904Ft
7zvJGolSVT4bvuqvvHFnH609pJttBc/5TPpgWQ6qkXd1uadiDxxu4rbLNXPMhoq6
kJhCVQEhT96RJjKXL5eztP/7nQZefctvK7Dzb3+2EAQXvN35h/KwB1MOhmgugDAA
Q6aFxiQ4/8ZKkS64lPz73hJTZu3ItklxjLu97GRFncuhya3kQ61P6fnEzSu8FlNG
gSaF3DQIgzUPEkzrHleyGWYUyQsiEiOYKYQrL8qp7zOinasSGAtdjCZJ/9+47Sha
C+T9grNIoozKpVbg/vbC+5sdMDal16WURheXrMu65hPEBuTqiDs0M+Av8OL2Bxpr
WIhsvbOMgXBVlXKIgfR8iYXFpcWT7f5YJSOO+JMLA/Bo3UELiTC1rL/DSJPt1Qy2
01dF4Q3uiRf5+Ygllm5tY4OBiE2NXrVorMFxEKiAs3AbYb9M7voJ+2OQ+50xywTb
gCYH95XmdGn8BZdgxLWardYwHIUko8z6Dor75ijyd2MCpk97ny5wj4iNavG7eyas
C/Y5w2Oo8wTQGLrfxflIh0lRzKOs4Tfp9oLiCYNh1w+w7NuyhDCMjqZwZR+OPcLl
BRS4iNjN1kdPIAReo8sbzz6hcYa5vbh+h7Q+J0tf5pEeciHXnjAq6ymr1F1itZJ0
GLGWFGOTpxibhhYeVxbx3mXLQ4YfcXwwtKQw9dksRq/fBMaD+wjhzamSq93C3ksM
jSYHu6SMZ/FRWzHgWQ78dBkNixjm3J9wiCP+OJeHKxwW0bxd7EFCkCjhZmLSJ68B
T41cX/s0YCq3YORQ0CDSEFoEKLFpKm+GT7TGbSJ7JK9QKcCkbMsWrMgV7GftTJMd
tYuGSra2p2nnUjYhhltLjAfqKZ0c1byj7c24gphDRR6CbQECI3PRKu5C4U+P3jQO
IvORTYQ+tIUkVS7czl5uP0q1QJAJw8FHWUQ7r9NKCbQ8FD/vpguLec3ieWOTzuCJ
atkyc6D2VmIpRKRF+PMUsIPg6Acoy/5F99+r2oxxgPKhifnNQ3cJmcc0UDcFMURv
YfVbpgGXlaj6xBVmHZx+WFboT02iJv+i93vHNUYzZpxFJBvJcR3Dc8TwDSlYAyQH
vyFUEVzK5TofORXa9aa95Jl/vwgJdh04wIfSB6GKBXS6ZMZRu3sWhvY5xFTMsE5e
5dYAElMToapelB0BWCobjaXzv8MpEAAyNFum3MXRIL0MeKmof4PEAyC1e2FM2LYr
Dlq6mZr2gOPjA42V7zJbQl/8W1WM367NFAiL2XJ6hzOzevv4PDXl8o2Hwrb3kcv7
Q8DOPEHFe9jCvlJTZYTrAZpFYVAl7FB/Gwc4Gdo8A0nK72b+h5HHpTu4tIkmLakZ
mzY1iypnm5KI5p3QDP7M3JlbVBJpnh04dEzN1WusStbOkakILFtX0S4wWH6zq6wm
2zvdkmIM9lKNJkWQpDX12s1KpPhBUJNzAM5OAJ6+em/6h3ONp6eKxv4euHV8dlYq
vDMDz97h6seBkI+M/lCNe/rmRUGB/vGfM/bO3v08MHpDbYQTaK6nXcjw3r5+TCLo
R5XoETr7uM7qf7+QjRPVEC1D0xOzc67pSpXIpKxVXmPg+2+Um5VyFwfd34h05dUL
1qb8+Batu/lAR7JZ0egERQAmfSi5GeQpz7R64tauYTclM+etyN2al6dTtAIv4usw
EVtDiRicD8I+ycJ9ejDyMVmw3x+ieJ1EQ10HHIqkFbtvYabQSN6cN2dw96FQLTJU
Mlg5+kjpV4BuEchJGQb19Ny0mhkCXMUJnAcNK1So1XCLiMKiccZKd/Qy/FgVNfZh
OrIKBfCc5J6L+qyAqEQnNk9fwTwkAquVc6wjkCL/VREtiosrowl17YJzkfRA5/Ky
hAtsR44FcE5mm6UHOhPG4iCWH2YOKUvXU5kqCxBO3Y6Eg0CzaZHn6mPJiLD9sLSA
yI/6BgCF9I/j1btzSw+w/qZoWd6NmQYBpyMXu3GgYhjdEzNbRCOZe2vPvT0r6y5o
tANtxdvqPxMfh4SaWWh0FQ5JR7Tzf1X3+3Fi6NgTmQsQC5msRly+TnMeS7IVWRje
iTUFVnpiL9VwL2GUMlwjORN33MJSrhzMkIqbUuvlRNJZYpV4AKJ+G16Q7OmVTUcQ
qZeIzZieRh6UTpwbi/Fxz9Dx+CC8PWeqGEqCmX3vbptZJ3cUQeUqlBWlRko4vfs/
QN8DWKXbkLRF8bhYaZMVXSmz7VGssoMHKcwwlctZ17kpaVr0I69wQd7g8pjoYotf
o/MAm2VwzQR8Lyo1EM0V2VJcL+llmgUEvVJEnMmetvADOe09AKm8UxumfkOx72qM
LIWFkOKk582osoIemdUVwhkumvke7QYryWBniXC7LiyDLBUk94SyryaLu4jB5OMg
Qar5jpYBD1EQBGahVgpK1GdkMPzed+RTpbZLXCAlvRPyGuhXbhipZJLMxSelROhi
2I8vmUl/NKWZe4uijWc5sVyYWtOB5xWugKU1ARy23YucMCtt5SGB2nsFvf+El+Sp
eVftVKB98imAmHKsCypAmv1OPD8HO+6GWqk76UMAkxH8O8WGJUelgUKKZphBleuG
T2ziT0bmIiWWqOrDG+TDFAwIHew7mLvaGSjZhPNpRtCEBW1iE7gqXHfAr6Ixgv1K
5k61bkmt1KKoOF7SDTYhbddYsqGS6ZQtNGx/2Pk9u/4nqlAhxhnlZW+XhF1t2Y2J
AUqqHg51HP+fUyw3ynSw/xewPGMrMMqHEd05GXDWGQTaTPJmdQUec9lIFCX1hwoJ
Ar3pQq7AqZifqERaJNVj/krpGIygaybyxyeCY1Ui4yStIu5eJ54d6Ldm60es5QIp
vMXpMlgB9nbKcnrWewjtBBy/13ea2knt3VkhBAs2Hrg2p41ALw+5ceIkrNEK1DmS
h02Vtp5nrzJ2ze6iRT2F0QTBUcarfX0p4IYruNL0rvpOoMGnsIENjczGcBU/MlI7
dO1o1EmE1aDXgYRWJgafoR1Qvt+RSBssu95CP6uAI60f4ZbXTSHVZk3QZoHBG0aC
Yhw9byMnVDCSqQg3MExqlky1LiZXyoVmn0P2xFkxqbOyKEs57BYhXDbxK2PqOjYK
p/r/EIWcq2K4Lp4IDpkGgc3rJffzI8ShkRbMAGzRLw+vCERwmzbOvZQFVWNd0/46
t9VgoioSGYR7LHcZXj4hypO6o/Lr3Di7DPc+VRAUORJumbVBgE0rb5+FtEdaKTvD
K68G5G599eTqWhBhxG/cqsyOT4D5iCZ5LgPQQ/5KDgwFsoSBbFsW/VVVt/mwH18R
f5Wf8JORJEnSmUiGzO/ZFnaU6R7+KZ9T2xWGFRD8H1LZ/T7l0b01lB/09Unt5A90
PUTNuEGw9oqkj+UC9CwBs3bL0uCFw4nvruTQBdB1+4kj9qd5kKJ60M6PANEZU7pu
uwt7dj7DREmfMYtlSNhDcx+S7T0BfGi1oWK+E6OrBIw06tofeYQPSnYRJthtenSf
d6RkRaZm6adi/n+lqeNfQZrEmH5nTsJrfNHZa9BVBmK5q4QrZEJHVdvuaTrmkFMN
KFcs82sSXglUsutKFLSLE386YAFwdLfagi2aPOzvrLgy1DOnRhStb8xV90sImvZn
WQi5smHqnU0tkePawiIJkozJOPu6FheWk0JsPSEEnzQu4794tE52Z2s5JRzM9Gr+
kXYhvf6kH1mNosh9kSirIuPb5alNGLiQNqiJJbvFqzxZT5o3GLukb2R9CEOb9XP/
Tj80bn2y+tNPvEmplDGrA+VQXa/syBnHmKx2zI+kukbHGZHa2AkT+YhcNKk1yb3t
EzXP41PkpZCCpN3HtFw3LkPtZSJNKEnZRMPN9slK+vw95zvUOPe8Ns40tWsXToJN
iBnTYnbiAEXoHXUrUDmc935jD6hqCXa1HgjzNj67+FpBtFtfoFZjSoF95X6UqjTK
YHpHHz+50QWHX08/3iOkSUxxzoi0W9aTnWTCXz5FmwWdQnvazuOuy1L56FHOG19T
wkdC6MA2RRD71yXwbmDN04BIPbuW5tnGxbjLa9k5n83jKxnBo/Iyws+XQTtS9/D5
yPQGFrtQtgm8Cx1lQ//rYumkagGbAcBfQIqrZX1/Zlujrn9J0ayOJDTVt6rLFOT5
QovHX9BBs8UYJXkIIE5cS7MmcDzQtL6R+6QcSpwq2AcHBERReml9+4MzTZDLdxuW
7HRO619jIJqaFXoxUMJ+PFsp4delLwjuvKSHHzwfNCyQtiOyeAU0KsCMwbA9i2dW
yNPvtPYrGIiePVUSd/xLkGVXhIHzDuCOfJuKvh2sBNJuNOGipzN7bTMlMIr3UGhr
OwezlFb0Xg6WvZ3ljKv7e6nIDOr14qnsklFdAfsEeStxDz1Fb39rwdhA4/NcKzEn
GbDJQZtpHRM9L8JXrEQSTiZ5E37Fmk44216vLaJRkX2pRMDP8iaIeJJ5wfvIgpfG
vDgKHIkgd+qyxJf+E1CQvldu450+BtRzhK1kVxR1jLfZYMEe4PgiMm3ZocD4zB1G
Q120w8veB7og9ZhbAO2Tttiu1H7V2o4lm8aWoKk84FIl8OOQvZK/agp1K/f48ljj
3u8cJFfBzP7MLW751Fr9yU8uHVbGlm5WAtHoAv8ZBA5VpK6dWWxiAAabJ15MJCC9
s0kBff6tSqq/a06zY6TtiEhoe3zPB8PB+g3MlNL/tXVCwH/OJHjbqelK4xxRK0tz
xwntEtwhaCbh+5aX4sZZPhD1kpp7p8B5+Aco6HUVZijEXhUJXCRCvFbnK9uro6yS
icrKgpsvzZW9KBOV8JY9RJJnjRpbv8F4onOFRdWDen8x6Cewvy+FNEHP19016V1V
7QL3Nhr8IwxvJS3kRplMzQgihgSNo3KC8sjlYmvLAKL2rjjLM8564hZbiss54hXl
J05gcg0i6i1rfHur715CX2qkthtY6151S3tUFu9HFeqA7za1mQbaw8Qg1/sCiSdw
pAa0VMckz0OE8Qhg+561Imk4YSzpNL0n6BraSSW6OFu4zJg3TxJkKiBGA9KRZMxT
eruq22Sym8Ko1H4XN80N1XEFBqS8adq8BXI0WQrH7IsF3utqGnz0Q2XGvXi+4Glm
o/YkM7NZPG0tkHF4ISD6c2WKis2XrSZ3y/6lLYaFS9pzgdbbB4QJ4lNCgxu0Yj1P
n0Yu0nikKdqlIN63Wke47CrDKrtzHetlqKvpPujSLtvvRriVe44BpJaP6vp3XljF
Q2PkT61t0g2GRH7hicmbALrceAgVmlMD4VpMZIS+zspCJuBBGu5vzAGR9UbgcIQN
//RHxZcVYV/CWKKeOFjRdc/LvXjU0FgA7S8XRb01On8r6j3oT2sZ4OploHjBtc8p
ioKHkk24bfTV8Ii9OnSyXpZmGc9MNOS7lGvlegIl6N0k+1qpr07UaOg+Bhdj06r9
+egmtCIZMTKHFaGPdCVJvtCgZWpC2cSlwjAj32kx6FcXbOZj7jj3cTSDRhdeYJDM
ML56ST5U2w4iTJcg/QG1EcJiGBoBMzUWnYid+p0YrtNvzpVg30GijHua0Z27sL5l
GLbJ/hEva0nN31CeIPFLsZNKO/Yegf+3shViMQuMJ4CvFhXf+cWBjQ/EUBWec6Ry
IhF3XnZdxjCM2aqqQPjWSeeQy+qnXrTqb4tNhLu+hADax0GBH7drsMZ6x3ji+XBz
TfERuBWCv76xF9y+yp3tMecHgGIkFUJdXoHNfuwSph8kk26RV4rMed7oyp2UufI0
ejxHbrjWRy8fGhOVzjDSoDjm/3WP7Ac7jvjC/4S6V+UC/WGRQSf53FJqZx3FIdzJ
xC+ZxOAbMubisA8VgBYesrYzhtNx+J6PncDXbisYFqEXKl5Fa8OPurBQWrsHU28R
jBg7kFe4FgGcNBlbo3qiOiy+3EanfJFnOJcQjOQlCh20/PICxVYtIvf0T4znY2/D
6OgzLv0X3ixKetBiyDtKSieUVUyw0A3H/tzxepgo5rVRdxGm1y24TD9xpdW6L2TZ
1eUvt56OK+1ZMERUSHnc0pJaCKzpIznw+3SKjcqSiiukbiVh5UXaFXRAtyDvO8Wn
8xlB13PJ38lSbryfdtSuA7uE2/WACM5iLjFnTpzWpoZyLMIAnRWCtLPHYnl9wBJ7
kDVzDQ61DH1ACNShxiOVWwLYMVDhQvyMNGjF6qlfG5hDE7dMblfNaha+eT10SL3p
kxRjwfnUKrOo/T2hi+kz6hdZIAU7J0tqrS158liqvdBex5p5VrYMGn2spK/CqTJS
AnLc/kJR9HBM8Jj0s+dsi6MTS3v8Y+S18CaLEpLob6J4LHxp8zTlKEklVx4C+CNe
MdOAjEG9KU+NSBgB4Uq09OWgUkBxgnmLSyfidFKqwlO+9WBgp1JUsamLvfOy4Ifv
3DU92EzjnH6rm4d28Pfb5ned5V900BNto/0uunCpvqXNy+XV+yCwbSEnSv0DcOne
pJDW/ZXhLI1srZ7IM26H0xwGaMpeEnurAthZ5x4uNU/0IEmuz2uPuLcKUpf4PAds
MGwB+AO1Sm3bv2g3EQCQ3IAdm5ArouV3qXOVCavA4/akBGgNrFY43RXwgkGGIWGt
uqE/jQVucV/BViQNqOcYo65jGhoANWoIkQteVl8/mKpQRQ5qy1bdbq0nZAOTrXSC
1ZpNs3KNTDuNlYuEPxszDOtwU1G42b8By+1H0yLHwGouFkF8BR2VxRYsjUvGfWNg
+H6lQFtVKTIGNZGsfhtwaCy/j2Bz6EHH9spEkfRpxYwrztlRR/tyKBEJf7NTjkfk
Gokty7NgRje57Yq29tcWImHQSSBpb30VNne9Y7KO3wmmaKqNjnabvSAdSs0FWpLm
8Cj5ZuxuPy2pIxLIyO+mL3BUZWJ1RdVKDGv6OwxCdcOmksc7btTWO4Nzeg131ODi
4ymZlWZXiw98IgSUPGQ+UfXXQLwSfLEU6G5wSf3Gl0n4OUz5IrsWzYeWeo5dSEZ5
rpQw0JNRk/xKSKpQgHh5+T0py9bsKqem+XTH6hX8agyhWt1d9XV0v3x5mJfQZoxb
XhXe11wXvq+qBO2tCITxrGAOEqSsByLGYjizkYydXBkxiXKYTjWu2swgdM9CWt3E
VoTBG7pI+VajhilGJPmvTjQwqQebI3mTQ3Z9xHkhL/5Wn6LkhO3E5cVXQ0K0V/Vq
NBkqyt0Yq/78jw928wRv3GqGZFbriVvYurHdUQU96TVs2MxfMuG2ToRtX+bjv9T8
0muZuSOT0Isj9oWWRC3WcH6juYYtGsXF5f1RSz/Twx9AF7tAW0ozqJLp+CP+dNmg
0T3M9FBF6QDt6NFr/DZR4Z9IYF00rZagjpjnbx89x94wTsFmkf2JMCl8hHHvXuHO
3Vu08BsI9hnUGQSmx2WeaVpAkQCB9+7ytGRKb+3AEP/jLK02RjGzQeqJrmEtXEMo
PPvHPrY6LjlUae7l5ll5sjupQTxDD1Q/t/featk2dLcDXVUF01VJ25zyKPxDf4PE
6wmUFqijQ8jUzJxYrULO68pLcyxWVIWiTWIB4gwx65sn7MWm+18NqZQnyGSbEUd4
s0unanvi/PQCVowNu2NeFSbm2CpAB04OGHWN/PYa7GSkpHdU/SCInlUugAwockU3
ugaqGI/R6XIlCBi5EUPi2hTjJMPZlXGdo4s513rzcGKSVTkOfcJYMGAQkqWzRcL4
vWFE/pR+0eU5ENTjhjb1XQpWpWhleaQ8B/ZudUS585t7a0/ds5ord/ZSK+vVplG6
jJHNFmwsEGNaO5RAZvMptSy4y+6FADDCIzLKqKJWgZyNEdtzXPtto8iY8fd9Wlc9
E+hsJxnZZYhUTUbAd8XqSN/GEa2Ohxxek8eijNE/ShHD9ds17NXbow3UlQxliVvq
Ham5ibMKYRzjpG4QOaBYm9IZVf0XmYqqEzW9y211bSPtxFPIIu7+d9ck7g3ZK2+T
YEB/5TohEGmSjHpqto7yA0kho9oMIAcy5RmkOH8F86f1QjI/i9O+1+rcxuZUuQc4
ewZ48Kg6JwHaZi+1PU56n8dOVssUgq+RopMYhAUZzKjAGhYG+9mlQ9GdAwpjXFNi
doIpeAJQaPjwnyO0pIpukECPKrorbYIoh/jSQlOMbs48uV5ayPji0v3ZMqtWhCAy
IscbR5Y52XxSoGX4r4HB8fDgBSx0ZZ1Yp9r4veL9bwFbHrI40rVNr/+HxGHfofom
/qcZzfLJm+ceK6s7jjbziMNpAGA1Z9DeEd1zzWyuddKhv45gbw6+IDrTQ5ND7c0W
ZvvgJYhYEoFmYTqsXCAutls9ld6GroOJynFpVIzFDJQWJnsuxjpfQ6nFhRFvSmRI
fO0FgYi6jx8ZxiOH9rXJ+MlvxcMCXMDEU0+BkKBcezrxWHs1pmen9VKI14+NjU/l
dXDvq/oXyw3xivLrotIPIR4AIeXgE2FgY9QN144F9odWot/+ij68jt9JwQsu6HFX
Q2ibgD2m9kRBWGdsacgS7aOrqJ1JWmYZ2D8Ci3RLJS+TWSf6KHTL5Oy/0I2/6DyM
mGGprBHMpNxHFjdHHcKlx92rQ7qXXAMAaMwlbHhOC8S+Qh/Hup9DDnYe/LfFY7Qk
7v4h0LWd4+zrKPTVypIWQRyjncMqXRUvIzZkHbawh6ruwokM+tBhnXX0auHbkJoE
Xk23q37dW1e2kdFgCidu+zeNK9NDJjI+swF1rcKaqGBF3eKQylYAaIxFujtIf4cD
bIT045bNmeXw0IwkFTGSA/hdzR8OAMis85XI3Ot9qNyI3atLL15sgSvc/r1y0K4Y
U9uUsP9EwkU0u39+lvJ6tUuw1Iw7Nqy0k6KRl+GxxsCCZWrTNFofI1w8Ovg9W/KE
Y7neYYiBKyQJYItyzeVimuoKeKIeTkmUTgczul7pX9bByoEheI4CmcV9BO2dMNS8
nM446oSTlXm15w+L1d2ZhssImcQgUx9APKJTPDS3HVd5uCO7mdJXE2TH/fr3cL3W
pbUjDheUOa5hMK8FEX5CDb9uBmpKMrHDvOWeolSM+VlA3WENL0ARz7ASFlH73Gfk
GPQTQ7hPgUqbyDlUeSfKsdePKfwWAsCzk77UqoH6bkMy/MJIeohqDdgEHCSEmO/q
OwozTe0+lMK7YERnwgiUeMN1iZD2FnFjlLVpKMi5tFkIbZaUnNwmbeyBwo3HsJUR
lgbU6wXQb5xtirfcP71vP2OviA2h9GQmekRSvXaer0Y441v7wKWZHHkmKoWJSy1L
MLSdOppdvtG/vNmZZ9MSsl5IT3WsVZpmafs0yHtq4wY3rm+8k9HbnMP5nwMzoQRJ
v4UBkRxdh7BUHPBvva5OBLcEjJ26G6TNB3v1wGwp22rYZUcXO9Ka93tQ969fJYKH
tA+ivzZzNvZL3IvBE35bnl4LLYNMW1M/qPqig1PWGg/xrxCpPJx13AJdKpEJIewC
1f6YOraAVxkjzGKKsd6b4xtRAUF9asbX6h0XyZxh5qu2pG7wpstEgUOdc+JtE8tq
x/nE+W5GUZn+NExGI/i+/I5Uq27nXFsWdsm4ChzQBIyL33zRuF2ImDu8Hi9hbVHW
1jZ5iS86jb4H5fOIXVcRPlANARSWBtO7mo3a3ArhQr9+T0RQ5Mndz5wYKWUtuPHu
uRuHn6OEFZlhrHZjB0cBDdCB6iRM7ya3tIRvTi7NaZDpcgHynEsizO4+9hjjzB05
UfLVJVJAsttQxWngNSYz3SZM8DksCz5G32XPz8+nS8OMRJ8AEQ5N3ScZ/HUshRMm
kHm746O+ozUW6+jSDAAOLWo9qLGXqJ1BEGjKJl42Yzk+G82TeR6UTVKaY1c41I+o
DQSHMByvdDb8+Rlj1ghrTw45WIhDkKPPbx5ZaUwQUBrsnEbxBwqeDPOWQi7m2P0p
qmRWf2hdlU4a6ZLIT7XY43aC4j+qIUkoxLjb19U81lINAmIUGhj4ffvt00tDfSlV
zwAaw1BkfOCJW8Gt7A5tVfycRgZCBR3aJiwDbIjL6SOLWMVaVAxjQBWqOAr4JusF
XXRHy99gQdm4SEY5EQosCWuIdNrNj7BSstwNNL4dZUjJh1jurQ4P5GMPRYL21XHU
cypVz8+wWdag27T/vZa2EsIBNrsmqcN1wQojBxbWKgh7YUNgHEp7mlzKedqy4tHG
vFc46LtnHHGrANm9nfRNkL7b3fRy2c0RwXNI+E7THF/F9L91PxGz9d8wuH8dmK0o
x09MjycqwwKAwvZ51E58fF6cayV2trSWLsreB2GyS/5HdOcGCxHaSekOXb5ecpvX
2P7l/R+FJVOYNu1cScbyL6gfY4t3BAAeRHxOHvhjM+XyxiZ34GqX2dG/XB2/A0p4
1PEjReZghjUZTsQvblpQ8u89ZYUJIuZt5+pfuN+YxQT5W1o11dzdEWxlJDofXX+I
NyHQnUz3pw54PLsBHVNZtL4XoIQ/kVJo8NsF84M5k/7kGm/ej+vodftdwp7rM8Nf
QAsHkyTHsjvNpFiqtUoreFhUPLY7Tn/z6bGE8VWy1uBVdVLOsy9hfV/ViYoDB63n
yynlKHWYjL4ehiJpcNiFyz9Q0IiIf0/bVhmYIoeamnVVBj5O2DQlLMUOwOBOv1hU
8YWm55bG2Mt7JhilQgm5nKk6gCH5BuFVQD7IoiRVDS1hUscWK7CukG78YQyu09xy
Xm4NQ2UsKR+tod2KNUFujfGFhGdhfdPKTx14uPvs7mRIEOenQKom1Gk9vwQ0BJkN
XIns2WKcN/Bf6iUnIS/RJKZp7xYBMbEFgwR05DnYFTzHAopeEJIkb8EIjfJEbGxe
SHDVqQ64PIlj29oxaYnw/6abIWN4Lsa3v0dL+u338cV02Y/qL6dtMUwDyGE187ru
qu0w7275C23+MbXcVFCDw0831Jqvn1NyeRODnP6sRNVwvV4uAI08IrVqQG038uNg
Luy51+7erFvjpcqCMzSVl3hb1LcKMIplG7h1uNWCKsdUnm9KGjlo661RrPflmCAj
NOINSZlbfvHRp/3lACuzQlczvt0AknV7VMEg91rnNvhXurUX2vHz9yn6xU0frfLA
JbiKMpXHjZWbyixweZo4URAYX6LQ6yx4iZholGIfIR6J38YB9pMxHgcIkCey4CDO
sGrsJn98HTP+SxWC+h+PWr496TevEvuMrNecYNjyxezo5dMcp1SLnSprmnMJfMBL
L+qBoOLnyjKagNCpCiP6hkLxhzuqW3LjUJ+uwr3Qblb3gfIr+/pY6G+vek9AqJRr
SpUj1nODEY10kDH4d+ExUy8X61pf2Io86FxYWR50HySbys9in2goSsPybrAQEubH
IXpFHtq1HGfxmyYMlcPHe98gEaNMgVDsXjG+y7IsouOFhNjkxe+3N9Gp0jxFBMyN
JL7QqhqdbLgXwX/0HbGVZwiWW4qTHbF+u07nSBfByxkgvqM38PwSeMojsIjN8U0s
Gy4ZZvqpacFh0SmmfFLiGrlw3v4/AqF99/NRdjP9+NG6hCAT2IQ2RwnIoWl/TXSV
3eQtzecopMnJHjYjgemGaRcwvxJrGCAbnDOUAs0dUhxmja/+f1geA76KdoRFdlcW
dWCOYyoml3Rwv7vNp/zdPMfvPW1Odn7ky0OLBRMPhGf62tZR31/+TG3epA9usJ1D
9AdbqWN8Fbsz6vKFJqu4sBP2BTqoskk0FE8cyCy1vCLmCpupMoswXl8XJOS0D2jL
AarbqVPkGO70aVzMs4ok5zTVIhmfNys64Ruo+TrzP6cW6cs633D0gg44cq5+4Uxo
gNmPbW1ZhDCi+kYqgQGdt4eSUgoegNPPcJxvVm/er9fPYKMmtjdQbITY3m7UU3Dj
DvRTRsXjpTBfzh7ZZO5o6cQKMFFEya4OkOkQazHYKN8yHZclLXNJWCr043hlTF5P
LEq+8hahaEp/wcfiRcx5Puqzqevz7NG4IE3Ery/FMxAenKOlqRsK17qIuk1mF3d5
kVXycGh3jROde0OhLk6LkNwL5gLvB6yIFc8eUQd6p2FA/K2kg8lIG2ABrq8x6XiX
D7W8yE39wjKud8R2KSHbVyqwEUiTvVF0P9wkVKbUdiXUVt2+RPx+RFkb3SzTaFpP
R0+ORUKJDvTqjdX1TCMPkgkpNk33B9mEZJDxbXDj9TzK3XyhR9/CsycbqFpVyyYo
f97C21UPOmdRNFmK5qdEziaT1Ibh4m/7BZXZwKsxklGTOQw4Cqpz1ak3F5bDJD8k
PSchs5JOqoA00mNnAfcn1IudaN24QnAAE8519H0Rl1erfYfXh98Ty3HoDyLcRYzA
HnLwW8OdVcOVzgejpIvvtODN9lSPv0ZjkAt/jLI3CevPYCWbemBYwdtF05jcF+2d
uSV4D0wIFB+1Fbttnm0q3lw8SDXzkW/GME5oqeook6/aPx0tJscEQ3DJwAll1Djz
p5iMwam7t74cD6Dgk6ogfbUdHtM2wz7v3NHJ3qWFE/Uf/aHTUcbHMeZ+/NBPeNWr
qWEFljafaqzGD0zcMbGpFY0VLujiqS3Te9lDDSB0keXPBWySLsyQkZDXgNwZGoMk
jT0rpvwPfUgLAKStTon8ldHDfGo7TbAHt6oAHa/Y47gp3jH5Pqd9zgtGw7bm4o2e
7XA7qGa+vPR+qAnGrTIlKguKe9hR4mdj/IF5cpvHi3VnITHXuOlf8gNuyt0LHDHY
MLZS+MevRpXXXmJB3zhCI/CLa+odRntrz8qyxa141eR9lp57BErWnPk5ZKcbuKKH
BO45jfvKgmg6k4o5ciIqdEmliVQOVVI5hEtreJ2AlkTiyD4xmF8uPUQf9+etinTQ
gaQfGkUBp6IBN9+/lbdaXeri7vUdKmSrE/c6xfsmKRiXovMkPPwB2eQiWWPrAX9M
3eqzFP1FoKsypgwRY+vuybfNsHoKJKvFXNCVunv1vF8jbzPtSRtXVFPAYN9ikbbk
W6kBteenjgJ1Gy9770oJ7U0SlDaFcp3Ew/O4ljPHW/9XPjDbDk9J2YfrMIV3G4J0
wh5bhK8oM+yZulM+PKvNoRoXRPFb4IjfsAGpvXUAhX7wUd4hswtViQhCnshqFGm1
s5Qp1pVlueLUQVxSr9GfsAw61QWVHgFNWfTk6oh75zDkUO+G8Ct0/YFg73YmXcTB
AKg3FaFcZL3M745mU8gjOPq+nYB6KuZ8uZcfeJi0vjxXqlzw6JJs68+GU0qBo85m
NU2tKf4QBayVhdsCE8bruJ//GlRxwVvvxB1QZeGuLI9QiDhbGdRycsVyeIXlKeos
FQx1GtbsIgR776chZifSLSj/s8dDo7HARh9+4+Jh/6+ftWfvm11VF4SUukAC1OXc
vbthSEJvSBVQhdxjHq1+7WkdtAwRzyMn2wC5bZnNXzHjRYHzkRSgHThx06v9IBPb
E+gGnUWZikOsTkm611zck8W9NizObS+gqntCGGZVDYcWMKoV4Upx3H2MtKnqvFdA
KKgG1WzVh2/lifMJ+mk2jrjJAVp2WMNO3ULAvtLp3mFo7uQ8pyOKJ+YVL2Jgw7v0
nrpCRqMUMkn9hSmwNBWH7dzf3yX/1Hcow6boAWKPQEpLZy0Ro8CtQZ6ohmi7EniY
yyuKlSp8Omw2zHFdAAuUQ7zFEf71ltwRbFjnNJd2rsdR4d1UagNuoBOa6GwZouI+
DLmg+RNjn1yWTYgsuBc6J2K+24N6Q8dXq8loKXQhe78qKAoYZnlaFRYv0x64fknL
Aw+OPtVvaQBmp36pt3vgNhdnPyKy8UCXSEpP5ajLF71UyrHZzYOThJs0yAkVCPte
CyeS9T1/TcJBYwQ5nGFDLDdcsmXIj/aYxrmU4IpAroqU7MFnnXuCC6HkdOholWuo
gCijdZMOd4AVkcqLCDPVvyyZ6FF6JYiS2VeJlynL1mnJnlHVaCl7PPYw+jZKWZFQ
coWjC4Du7yBH+LHBcZjDJG89+Lln7YJTDGOanlSnM0KTrHgd7fYD1CdRSTawJE86
WLsTzGzg1YncR96AZgwM4qptBnkFDQlTobzR2yayzAtCPK/q3I8SzDSxDdayPng7
2UrzHOyRiRT1/HUK5n80nDuV74KfoSzjQTO46t9h39i2qd74khsLzxCJNO6Hmwd6
1x9XVyxtPPDBQiOOfMCiumaRHCByJlXGNUfQ9XS1HpfUlygs6OCRoncu1erkMgdg
wytqgcD3/w3xGH7DFDQTfQorU93XRibCzsy1xZGeHg2pwgIi/o4quYu8/kQl4sDc
FQzSrdRFbjfl2JjJq+DOtJZ7/tynyI1fo00flA8N4Snt1mQrzU325N05JSXaB7Wp
T5Iwnr/yMUvBcav/RS7nEMMdkECPpzUMyT1FKlLM9dXXiECMakLDnvBwLQtnxsBy
0OGQXQe8SJtHUFos88yaP9OoacVXhptfR9oeWw3iGd/FEABXRR/4JgVdHGgWCLm4
Z23BcxKcGwkzsEMWS+T+2h4SvTxOKo/NKxJqSsyibJ86u5TyI8S085fbhqGIBvjz
Hm3PbczPgyZvMayESRsHr9OvJE7FMt+vvMbt6TyGjMIE002jwVXmwF/PfOdl9thJ
syD6y1rRWSCJQAV0C+gITsMLWf6QS5yjM3OJb4y45ACSzusHfLGPM8l9dUUjjAH4
saj+aPTG7p1aLrSsuf5AGnyqjvdIDSUV8sztVPFsouWyICQgNnLiTAjlfzLIF//4
OKtEQjbzEDiaCxrGVYuALK4/oGKLqIfyCiLKqRqhIiW6bnLk4Lj+DZpDtd3inWH4
ErCnOX+jZ+MvzlNQ3la1PxpW0E/qLZ0HoDEvlgbDerZjnR1vvB4D6tEWgZbzR0ti
1yE/2vzR9JHmrfg1SsBdZONEyZemu7Ps3AYKs3hLxbuiACBDKuwhgc4XzFy1kkcr
pWvUcvHDdHi69RwdmViBiDuqp0G/tdxJZvQanIdW0ujOH3WO94FVd+KnNO7IqTTS
yTutibjNF0DoHhK3pqILLreHCgWaJ0UunYIH/KiGFTcH21Z6jCk9GdgVFQmZlj/8
g5tbSxYlWVe6zfLBsPiTKlYcbeNK0u+ftfhrO42CLrU4VhhIZHpUFNN2TuLwuGLe
225nLDPUYelVfKqLaf2sNBezstbOdG/+DaXRLZIBCZ9hCndknv5a3LTO26HI/5xP
DwtMoqvGN+wevTxyLXGhpQw3LEDRhuTtYs2xJh1czjRTo48e/IIKjWMH57+w4INB
DhT46CIWcI/ruoQli1WZOsHtiPN7REj+PkysCI9nvClb7tBknPI4QZXqmQrcr4iM
XFWU8Sy7R+RK8b5lW1Un2/MRxxEhUmx/NlsXPer2CjMvzntB/Iu/PZvMVupd5rBy
YZEsvfX/Go3dVWpwKbx8UuttQwrgi1Lj2jh/Y++foEv1T/oY+l2UtC4LgjOjt39M
wSeyztLzElO63es6/Qu4IPPtRed4sBCPp5VSKPMHBUxWGGcNfVlvlKGgiQN/sCn2
Z8J+iqf7ypejr10v6RnvO3ptf/q+yOYBHVfmPu5823i3taienEg60pt2sfFND3ug
arGQnh/4u0KJVJk0wvsYE2ZMMuHJ0slvV//cxIOGJMSN9sZQ54aKF5Lq8bcOYWPf
922NihUC+oXn/pL5ahKW/M7V3yDSzUf8J8Gl1PO0r/i/81ZmNtwiFmxlZkTMpn/w
BpG8H1pJ69/OuTBE8eq3MoH/49d+h/HcLkpNORIuc6pdvsyjkJg0W64BlNDRoaEg
qgZJXwnhBPOKwflT5GPI/QjFfS9vm54tnOzWts2SnUYoMrQJgjpq8gm80Uf15kGN
5d6odo32FeGiFMYUoTAc1kh846IFzK5irR/8pzwm//3HjmRrZVdeo3kGT6CnOT+W
RLDj3BDFbjiGI4R9m5bJ07JNVwP9EH0UlxTTdbDplIIh9cPU9hjQynqxzgeG2zMp
IWFZIz6Yx5tHOb0jmYReLVc6WCBGy3m5wPynuGIWfGkbm9sjfxwlfDxVZstl1FWC
3hvd1pvFT3ujeZYXf1lLAYg+Wo+roLumlV9iu5BVUk/ATGbRwlbUPBSLMcB8GuDE
RT7vncQu84gyPst8UIw/y8NipM+eGNGeTCkPN3t7/URF1l8WxUOTvyXqYBZdp2yg
OMN1Qv940wYv35mfHg8ad+umem29fM9tmmWTHrtY1R9U37x9g0e1ofp+oFCKNwIM
B3C9Vic/Xu0CFJ3qvYVn+MX2YtEr0loXB2Gny1MgUtRh9p/yt51XJ/MQsICYA18a
pftUtjMcsGdCVt3uX2AqRdplngButYlAO4PTk6pLVAIcSEmiwPd/CB9s3dR++s9+
XjwPX+iRDkvVy9aI3o7i9jmOr9n79AnjP2VVyDRAs39wciUHZjBhydMGRXMXWR7a
3wm7gMr3G42kNvYbIB9V34T1HNc49/0qsgURYbCq8ffsuPtsQqw6GrQeOA6zwgIR
Dlw78lJxVpeGCGfzqRdCCzLpFiLgHA8RavfipYGqA7+OTSZrrjvzjigj4LQ9qGO1
xX7xScQSHM7GwMG/loFoS4of94ILJrmgGCqBKi/4skm7Xj4c8XJvUPdDRpmIzCR4
ydAje9Mi86EtwzhfsUuRi9xSESOsK+dLgiApjMLQ8CvV0ytqKbqk5ttAmeHjUKW6
D48zP4Sp2WDyldM/0VzrH2YwKthiOuu1aqEeYtQMIm+nlS9VMccQ5rwNnqFbteim
pUUmq7a6rwkl4XCQ1EgaNoPpa7J/xBmWTl1szBhlfoPWBx0C9is/om+Q21AnabFV
8laG02jTg0QmU1+v84U2KCsp4mTGvQNazoAEB8uEtQg3iQrds9v9sIvqKoSaKEXb
6573EktWepbMSODZyvqaQ3yu7VIK6DqCo/ssztnbuJS8LWDdXKZeqDwupylioFO6
FlgcI+94qMl6QgJbEtlQEX8sbHwN+DaK//d1eXHKFNQhIPbL909wNmbaSUWrNneK
MJt8y9rKI9Rsc1We2eHRzo9//0i8sBqy1Wm8O+Pux7dao+yYhmtrnehMLiY6EbhK
xn8WjGlMsBO5IQBns+4qpnAhMd5QhaNhgcIWf4KPVg2+/fME55QA4NP3etG3KgQS
IWJ211BBkaAKaTqKePwEwA34ZJ7ucFg7fbUtKMXBNmUGVokV2DRJZk4zuhfhqU/6
+pIGd8sLbsQIbcPQtSHBH7pN7JmMpD3H1+KDHLtl4iEYK4J++84U033vuJVLktDv
jDT0K3eHOe3GYAWRvyKeeL3pb2dsLxYahi/kAdbr8wrzd99KarwOv8F5CHc3M0z3
c3kmhXWvrdrtFdhAnbwpI/jHlQkCV0F+tscKpUYa1Pzuxh0Z8fZl+YN/w5lCqsz6
hPoW1yHSqGkTsWYMBLWaBNHtclA4vKCBxoeuu7X3RhFNEnEkBH/bQeddN21+BIwF
mY//qgS3Xnvq/pdi42NG4old386UuG2Kf7fRXbHUB2MQfOIx70jONK2nomOV2ATL
c1jWt+HE1Irk4ymQ4Epc6250Jtq+Jlp0Ji1FHtQej85zNpNq93y/rF06Bqv3Qwfy
Qq8NIA3grCHqPVaQ3EL9sULyvAcBOIppfs6dLrmPESS2beHa0gE6JWc0OJfl66KV
JUg6gUiVYVS+/yJSqsIltaNLGFE4Xu8/UCvbGePeLXRq4VYbVbo9IqWlRLmT1XRB
+WcJQH3If8Y1YVdTV2ZsS4bf0fqGpAqdqjc0POHLp8RCNueP3eLdkVfaOBu5KIXb
l0kxANcB3bT2DAO3nLLiqOM5+8rctgpKEByBWDogUsMCKansblAb6bxH7KhXWNnr
7PGpxz/MRp6Y8l2NAuvU01KxAhJ7Lmfx5ZrcsVIwLNFDOTMUR4ztY7FhWGTpBKdT
o6vRgYd02xVvC13JSfClo5lBg9L9xeGCfu6w7uvwhQzv/jMzqhiKUZfXc5z93lgb
yBZ5TtgRFFOomLNnp41mLTqMhP/hAVWI/rB2S96yBmEpy/u2hS0MBEhaRyk4ygCL
1pHeu8BQ97T2/43gILtwtM0bGevWIaoAFtO/VjMTP1nq/tLipy8BluTof8+NF2nI
KUofjcZkfv3r7PQjs1NUyZso8yYCFVEwKBe0S38FwPjvypseur6hzaX8pFcgZVQr
LRsj+0MG0l+oeKU0GZ6eD1LAefbz4OEf1gi2YzmAp+hZJhysUZFzBzUQngJ4JZwp
eETKNoOCGQZPhxXHxbxvaybgKtCNs8eggMeM83RTiEaRp2UE+CA8bfW/u9LUE4ni
1QkoErZHtLX1Co2oMQ9AsGdiX77DU/zMMcENTtmeoNFLCB6zKg/GZ4s8mMr7G2vC
D4hRnNn2MTyuLYzmSvgEAdbYud0LoCTlx+OqilAoleBv1MwG6/IkRbqhZqiuRRUO
IrGvEasCCQPG6OMUvRsI0DZiBUb35czoxAyOrclB1CqNnUmwSGANZnkwwyP+xlUQ
bvVkiLQ2i3cMSBZ+GPTngkfNUgZn2jmq4jSnv3hDUGaI79W0rWJCa8Q8HrLI0QIs
dQpXrTaKySxRAzJ2XL3XqO+J1QjLIiF1OxX8haopZkN7cdBlslEypxHkAD2Fcn0c
OiDQFKp1vWxuBzqQMmsiU85UQohkq2blVYTQvyUb5Tk2N4hAF+gNKkJkrRZOouAK
/I9ZQPGVVwpebn5cZAs1GKEHzxFbHqCudbouJIMKfTSBFCfT1FbijAbnU7gFVF9i
F4OD7hG2wdJ6UzoCsI+dg/EfwHxNK/w8wO5s0AR3EBqXlv9KFzx7kFFVNkVtrIWp
OwNdERa9Bje311H0VMra72ze3ttjfFjFfFBAsp+brWJzggI7cFxd0d+qL9oZT+zG
96daTUM9ChjuxO2Mzq6ptsKdIAafg2hFrurxH9dwkE0tK0fZZXBdK+EeVnMAS2w8
YYHZKpSGchlrAJZLfa+mmYxg1FPp9cxtvTGcKw9C6RPpCeV0rzwn2AfUyTBEGqIW
v7AQt7fEW3Vl3IzsOx7tNDSwjuwasUHGtfdOSlhnCrGBCcNM22i0eN4/Ce3+zqMR
vDZJooINVpt2w248Pq5iA2xE1fi+tLLrTRBJjuA5g1kmrCecZfmBKQicH6/d4slT
FYetqcy76rLfoHkifVE65jhJcQsejgVKXj6VDHh1GtY0smcrqWXVG/Hg/iO+5FqH
mN/tBClo4B0wEm2H2grkRM39tcfUo014JWQUm/dmDD4bUgElrfZwU063lWLVyfrW
Im+Mrats3i1EJsE2riSjLTR93MSbr4J5LAy+g1b/caT3L1BYPnA1NQvy/jWA/dpW
dvs+3zyI1cgHKM6q2uiuOwo3SFNluIklFHn659GrdkO8gJEagLMoh2jPWjiiR1tT
itMsHJv6zvJ5TzdYU/zJuEvabcxsUYPnHMBA+hCwr35txmKX5kItdZtsYoAVVxYW
iQNxVWepv59GFuKFbu+tMpNra/Xd0dNhWWDXNiSPFSoWpRMEvPGbnIz1lct8CMV1
dr4UpmDK3YeIcBR9FYAMTtAzSMa+rbLn19QKMYTzQ2WKD1xeb57zDgFGhlUWGi2+
yhL2wW+D90I3voVyyeABJe6PJutLOcOq6aIYsuiJzS2DKTi8ckgJcLE/X3OL1aJT
qFkPwGM6Q9gHSjiJG+7TZweypecZm2fAmVQf1JdFmHagvB8//01W37un4VVtZ1a7
ViREOunYds4F9jCrlBRiWqMAiIfkGm6pry2x/u4rLhchP0ezZuNs72/z3K5fmV6g
fYoQHJ4vKKfN4dUOHxAoAMolPw7Knxn0SLalaq9qXFXaqPwtUmOIZTGVJcObzssX
bmjky1S6IkpsjI4jLFO5n0RV2tBtSJO5A9W2fpyBo6sOtqem0Q4Ui8B23/5G/1en
YYFWvkFIlruxTnzh7kaZ2LXfADMdJHfi1yPT6z4Tw1KGpxPLdRX2IQlUUQB8R2cZ
8zUXGYTXaDOUiGKJdnJxcYMkazVlUJWKggnv07XHYVT6YIRzh6HdF8eJRa1XczRX
qBlH9PoUYUu85Vcdajfi/uFr9nwRuUVG4X3KYyzgWnv6xFScmG5CV4DdheafKWn9
CT5z+OVHbRKqpO9yJtqLYcTTr9UhZiZLUPRNnZ6z3OBhq7H7BrmQXRjF47OHNZsE
sErhhl3AJQFD0FioTMdq7qvco7rQYNx3L8W6kAp2AAnxxMTGP/otdYoygwticOtI
UU8jGdyW2wQ6yJarnij9inU90ftjYJXkyD9c62igwbcGl7/NGOO+RbSxCepTa3Vx
Q/fqTrdaF9on0Xlk+ZrNLoEMBwM5GWgYjgccR+YDWD+nXwqjaONS21dx6xdh0M/V
tb388s9Na8KBq/PPnyyJ7DvkNotTHKXdKzQsVEvB0rCkd+w/jvomqP/DtSSoRsi9
pd4cOo+9xp2NaKc1No+G9WC5aadGPtEh47xB/HuTwzydJMhNpZ8fWjwd7VqXGrEZ
DPRfXwjdjBBx26JeEc1GZtc5fOgQUJPo16fGERIYy5zVWzSsiFtCqb/hUQ4zcbLM
7+j+BnCLixisLJyghstBxJo6jkxHr29gzpbGTIR41wYPt9QX/AhR8j0sxlgCl61y
9hb8cyTyQCklmmSII96rsYZIRHqMrBxUQiyMaBnXGaJkLu9V4Ie8ljS8KnLslSXm
8AWqmoWJTCSZssX6/wBZw5KF3Rng1aXU7xoRcNDb1wtYj5JH8plPTJKJN0c43I6S
2n+BqUMv5m51RjHM+Ng1hrUSvVRle1JJsby5HgFhAgD9lCowfqO9bQaVqy08jqhG
PDNUhUrqy+UcgU44zqhAYvitg+ETkndp+M+Pv80OGpTpIPBYJ0V5pGD/Gj6NHAux
dgvZvlmn03dfrTT4f8ecUjNjOe/o2epDqgP1x91LRsreSjFzTYXdHOzQHBVAQuSB
zd7ZJ+kuu+9A3KF0+zYvBrY+paudJ/lJk/Q/FpFnDkUA/xpunrg5m9BC+TpNtjqJ
4/eccoqICp9UVTRGcEvql3HIZXpPaQOiErNRXsx6/lgMCV/kQoxJT6Bz66iIqyRk
+SNAEI+qIA7n7fqv4zY7K/SkMAu22B1cNwY1AdxKTESbe3Sn0iQpTswPXNWinm1Q
lzsetW2ny7qkotpSb1tnUQSLNoNrtSu8p/yJEBqV7eFxjnY2yB2Si7g1rkpp+9Sy
vG2oa3FM2Tgm5KGfOPBzPZMGR25Ph8vGajhEEuUc7BPuytkpd6KAA4AxC5kdTaC5
a/AMUNAL2GswZXVUIbp9JgBMl2Dqxtl5xhFBKSFGHBvv4VhewikBA6+3hZD1Kv0i
WKBMIfmBeqDcUZR1jNm16QtzEYgmcL3y6tVD5yisLyUov5or3EaVjUoTiW9fRpnR
3mmKV4dZyxbE+MV5Y0AAk2ylHLjYiGAHIBfxKqV/BRAoEn+niJU4U68J9lb5VWrL
ShsbzKWt6Ay2eHF7g6We6Y4GUlG77acCUA6BxeHIwiaRdHBTA23tlupnHD5PYhZs
MZPURitRJGqITbtbbwpYUxQ9QNpXBLxEcBPhj8uANdX2g4IgPYcL/7Q9MSpbvkbe
EkhXiFbk9t8LT0N8f1kawowSjCQI4ekEx5UT4qYZTw40xw9Mho5MvjcQ9Zfd0mBC
46M1MKavJzL76qznIHz4qcDV69QhufibRhCVRQTvVzKMS17J4OjqsCwDhYCiAr9B
UYADnlQkldrLg9FGwPEbJ0r0KFa+O6AzsRlTDRJwCko+bKj2NIoPhCRXxA9+AdHE
QXs27WRoRgyGTnNd8njunPNtlPVxqYc8ymzk+MljHkj/ko1uLOUyO6FDPSF5Ho47
Pn+VK3eNaBb7bQQduwkSc4fZKyZ2AjNT6gqO5lm8Tn7sJ3qK3m8KvFqT0eM0lRl9
CkRLCNVrkCX8T6DxtF+NshvoA6UpqKZDVBkpp5ZhACssMWzZresuV1QGQ2onIWMH
M7k2L6A2hQUamKJzJr8HeIMP8ieI59/ZmItS2xvKgZyg4+uUmzHWDWGxdMbZSMt9
IRKRgxcsaGBTgo/rCJexPMNoQziIqHTLHQY42tIL6A1MWqIIzs++2ZAdOdGYIFad
v0bMTW2PTXDnLqbrNmnyzVYG1FPtGgxwInkaijIEtaj+CCNmsp1Sdd99RKUrS64y
czpCVd+X4EqZJ9nuArjuvgsJXVCiM7Gi7PBNeQUYsWtPLN93SuRMNcViiknHvgsp
gqiVLikbW6J6ca3YBnofZnTb5TZDIToH0dZ5NI3d7+MUQVJPqKF8f0yuJ3iBDn2R
9qUBsBg5DnW5Fd1nPfTvizfijb1N3hesJRHpq/hsfVcvM7iFm+Kf/cr9JUUpGHZe
Qovs6PbzTDsA4XH1kCouDi+oMuzdyNgTY6qchYnpMDhGueiToT6t5LUz/SiC/B4y
Jj9NQZEqDTuzAk1org3frT9wXi16ZmqtAj2xoZjzmy5nVLE/wkSuO0k6ya9vU33c
ekXcNtdkybJ7qx2iLeLCJCZzIqdQGa2grEAPFPVTFIEi7s/yum/2txXN3GyDbttr
Z0o6+pNXn668Pe0bY2MDHjxrBHF5kNOoD3JEM7Usr4/pw2DL6OVnWUrhHK3OlYHs
V8AKlMIESQLtCdSLd0liM8Ovu6OcGJgo3DUY3Qcp03HJZJRXkEL4PXjchrvhp0Fm
QptpzXIQ0udGzSM/1I/sDQoqRwbmiIzg7Smc6eCIr5vsQ4Lqr+Xvsdwy1ZbtxRcj
BXxKdpoh5eqou0fcjTrfLWMZtYjuy3NDfhOlSofT7XEw6Dw7GrvOMPFc9rc/y9zv
tAPwPhuKXAWqZ3ytyJsGBA5qYaK2tFwQGzHdoToC0CSG16aimpoPtU6pAl20MM85
h7F60/YMsaoVXaBglAL11c+iqy5RsvMH9WsKyiMaaPfxjeHRvpsETR+hrIvXrYgc
9opOD0qh4qxCE15I5/NkKGkN258EFihvYpvBFg2P+NDBcD6ym7ZCP69l5W8Jc1lT
Ps0k50u6GptrZSOHKEQshzO69okk4KeUDRM+2ek9xp6GnD+stxhWyjaDgqM2i2hI
ZRWotuzDedcAVXVQ9z+SvLC7g8yKEwcDnl53/HKRV8S4NlkG07JZl5ANjBG0PSw1
qB2w5nJB4PK1imuEX8bLL3Oq1nxm07TPqpvazU1zpdaFl+tRdJYJIOhGSK7DVhHj
n4uU6MHNzKWGAY4Owg3BMXOHTnMQmVhIxMu+sH9P4I5MMyxnmz5cmwIs1GT2gAys
QL7NgaIh+JxhQTpFxoGeiAKSuFLz2TSziafOT68s30Zyn9mb8DzFgimAY3LfTOTh
Pk2YpSf/R87m+eKPW9jWo9YQHKmhLmt/QRP6AGL2zBHjLflzp9MlvrqJUyb9IbZ+
xv1Nj9ZjUVYDff0z76CNPpnpwZc/c2++JM2mIhqvNILIbmrd02RhFI3Ew/traWBy
X/KYz2r+jLWxwgGhr3VXopwjJYdF2ntZDbhn0z9C/yhgQvVPLrcFN/tFpwWJ2bCU
R3GEg+fMaED4lLF0GWeNYA7PYpI3IDiLeli+DG1tiUYHT0/dK7ZWmlGUjLojWdi9
+7G2wA5/rrR8zYir+WE/zTKRSc7BmgiwOlMwfUyKjpAe4RToRZfl3IaYykpVIjP2
45LcymH03vF5fwPrs1p/rBhUw00i3QtRtgM6NPuji7+4BsttsEWnYBnmkXgFwccl
ai56pm/Uo2599iGWMGThp/NGyW/bMhGwYpH7fIxCxRDQZ/0pmHEquJpVW3+L7V8N
XHtO+PBqYuKENmaIU4h8snX9cNgq0WnAHNAbxYdGOlnceYduCOCR9WXwUUhre2Fz
KulUHdOsYRGJmuhN5/cSBGoOP+dglGh21Q6S9FlvCkMQv6mkK6A6OUi1hXLhL5pC
NRz0euGtBMWTRA8WCyDEP38P+GuOmvBiTmzYpbqLEbC+8gQ9MyLZVEyMA/zXTmoW
xdbJGJ2ZTZxmR83q51awVh5Qu6M3liJIEJVsglXZMMDqwBm5MGCMaSyIJYsKVU2f
/nMdGsHP9MudaQ6KLwuxKCJFzSfVfqEDSMfXU6li3zNx7rsdc/Q9tZYBoynBQHzS
EDucf0kCt8mgYNXvOKMUZVhz+8HPhafnYcvpQIRBCuD9cX/QQV7p/uVW5yLXd2sG
/n7GHy5LqHlUBWJtlHEOsHKjsLER9LB95TRq0dOV53LH/NZv4dlt1HbNPkCltC2d
Yx6qOaEguestQIjKiqfcQj1OSzjREHyOjuagL+RLajle9tUGQD6PTkugUy4/MDuS
Trl1ZDcm71GM6hkqZScCuaeAez3UAnxtD+rFgvDlIJR0T5Msl6I9Ow2+FmiG16Nz
Fxgczs532SulBKxgk5Bj4xJmVglA42gC6Ba34J4swwXAr6wK0YMXRiBonFyMI3No
sV25aFoGiKk1A4iCRtTjyh3MBF6/hMgoetKzU12wdGLdznz6wBw5pHLRL0q6JTfc
GNajFVckNvB5iI8dSfGoj9ICyXYRZG8PbZv2c4NvfOnQd7pBCrGz/LzgV+y0Ar0u
OC3IAp7fN8ihKDSKBMIKkC7tuMXxzMmqP9Fv3aTnRSD7k3dXUJMB17teDfSPu45+
xIiOSXmu3bpdF7S1tdzTgwjYS0xnxOIfc/z/T+izwWzY1lzALSJEShek3gvzFuKN
oIpgy9WiZ1YPyE66XjcGPDGmDLg+MNeU4LNXkt8udD5lg78aAH0lUr1LlEVvL5uP
V6hWj3BNh+VR5a17P/tRzxUGIFiks/lt4+k2YYODfJ3l3gAS961bK9x60lSVnG6v
G1UOTg9lLGTIL6fPITy93+J1iDMoBhcGaqd3LB+sjT15gsmKCUEnQ+NY1iK1sxdT
msbCY19Liwf362gwigmcQ02FruHGtWBQTWe2WpQYju2Qm9IO8WXm3VvPAJgh0j0c
tR/FnVPlyJ3Dda/mI2VQZBKCWR4LCXbrIkyTX4/5Ns3h3z9fgx+iresqYykISh+v
HfFdyDaSSOympVUiPckA/+OX5kK+aFLeLhYIecVPDnCX7pG33XW8rD9zfUCcgVq3
OAhD5NdGm6eXKzoz8Ys26x/Q23qqtsjFF2RFpCk0z0fadC/YRi3L9Ib4Hylunw71
gmMXjELVYIQFs0u2+n5LiXfQpept8kxE0R8o+2aiGdwbC6uC2Mi8aH3k+fB4txPm
Pm1xcO49AL4Wsp+4KFomMOhVuPakg/vwySnZhBmvikV/w066tHFRcKJRdc1UrDWK
1W4NZZRDL9aqLTG+6ukw5L4fD3bdcgEmDTB8Bk0eXQIKHm22gUCcLdTaEGKw8b9r
Oz8y2sqjWerWplcSgzUn2i+dQkUIqxsyikFWEn3Lf+ADwmOa0MacT9Bp1vjfTTL4
xUMXRO9rDC9NiAqKywiyZ01jcw9swbK4JDV4ca/B82dmsdg5ZLoHyTbtPCj2GJqy
hW3V6EAE1mGnRbFSqV1HrMdx8NVsK7xcfxJVjxRKbY3SJ77h63yZadMP2BDlWjEZ
B0YH7+7fWpgsmzFQjGQ0wO54c2Sr4K6gvc+5YpGfupze+hEv97t2a8uBjQD1gnX2
5Kq0pTkjmdhomnVbUGg19JR4Re83qwCAiM9ZR6l9csGLH3/MUvUzjgaL4r5Fuofd
t2SZIMu/H8rmgXhkB7pG3u14P0LN+nayKXWQ4TCoo1yWrLvucR2giD1ecDujY6kx
2W7vNtFEhErprLVkbmoA7gRXN9cUjLygCviNvxAXwzmUQzDjcEDpW0M9P5JOEU/X
hDCTe3/62TJE49trApYM0hZAf1lAj6EOj8zoYto2BOBR6ZUFNWVrngX+Rv4yAdzh
UUv8N3o7XbRJp7khsvDFSNf0tVR+Yj1UwtSLiDokAniT6C0y5RT+6gU+HvmsmXzS
Bj3xRNmC7TdoZSr3LYB2lfXFmKHCpz2GepK4sNLl5I7iCdfkWOILBp2yOHH/JrnF
eopVyQAo5u/lZjyloFTtEnoy6a3ZiYCS7EhU2vZy2Dola8Ih7B/UmJif1awUMBgv
A6PehuW8Vkikhp3RdoK9Ryz7xJ0FNHjKSq9QZC3Rolb93Mi8VFl8uug0zu1Lzkrg
fWOU3Oj7X2UuIpX9Al/zKl8XHCuArGSrorK6rOJ0TPKwOF5NLw5MlluAXLQrAHcv
uEQ7IQ+gdSx81Y7EPePjLqAQqyAIqcJ8ryuU7wqGqlcwC44ptfKZp1ZwtvuYnKnt
nkuoF7zTwmfWbj/vQVubjhZRHWgd+tt0O3yejnxReXqhAc3mGE5zQTdy/GFmfz4r
Snj+NtmbaNJyN5tCrREJKIjjXs85H3NMLnG6pGmKlYo+GrbPwCEwdvZtDHxDJzKy
OdnoiOI/i1qRTDX4rtWPTFP05a7NUG0Ua/ZJ70ITOWK3B98sQ34pOde94l78BVyn
h49v1ZEvFKLn2sak+Jg6eW+nrbFEC1yafz1cbgTLn5UbuCd4qc3kvhfh50gAGfgQ
D9Ki7FXGBtqjnf2n1eVvZGVMADQwAuVwIW7ShA3rEec81aSO6ZKxJqdV7KOTJ1xu
SvP65MwVfvBx+hFh622F9/SFaUqFPYTfA+ujdI6uTkaQzaCZi+DAklcjm72tNYre
/LEpDW+i3wsQZfUj71YCuIiuQZW0TqiTvg4Tc/MGnqILDZXiaNaG7pPxuScAdzvu
+s73PkY3nyHfV57MDtokBgEqf152bXwRURkRQ+OHrVSnMoFLAbQ0lubz+xtpHrMd
bjkLLpYH5d8DFe9I8mHL7dsD1WjerUbyf8puP5+4gb6HVdc14+bRD38IkKFDLLIB
mPMknIvN6pnS8i00obd3hYLpxoK8JemDzyCG/o3fek5pCMVs4efooSiab011BW5J
FkE6WmaMsxJdNHg8Ik9NS3ObwBzj6Wq8HtizQjgiFmbltTLhkgAVTiqjTuTAJ484
eBmST/9sjLZ5vBcW9bgelYcCLkcwekKW4ZrZhSlDw2bSTV4vJBm+qD1jV3ySL22p
LdQ/Blg848T2buh15YlcH9GvVQ2yIR4RK+VILBNnPLsDHwjeTAVPnAqK6VXzokvC
EurtBFQeFzQWF1cw5caL05zqum+drz+MgPaFOqjL8pGyyFBMdIvgnio/UOm8SBoA
J4MbNNxdIVUfObRW7iU1stNzm3AMTg3LfpNj+hgL/y0g0p7G2xQidcj/0wAQkfH+
jZYrwcdgLO3Q4jBtpPIo6pyNEkp3FOoboLBpHbahysFPPRqivU28F+wAd/CAwUZb
OP4aF4r7I+LsXKxqZUq06eQViTsnjkgM6VJFcsS/3ncVeYLNQaHiqPvs8AsCFG8w
ZDiRsq+WENsSjeZxXryRdX9+P0cfjaRr7LiOCtg1O4zRcDGXmj3qYqpCf05DeuQL
2XE9dzJgDnowKrNrkjetQQMssBJeOofD/aj+afcQsMkIJ9RFQJUJiLsCTd9tcVb9
FC5lUh3pfpewuF6wwZ4hld6QEaBoSPdB+qtbqfSvAwcIQUPbstQujyOuFtJETA7I
zQNHIpdX41NbIfyWds5Ib3bjqwOgbpD/SvC0y7HcscIt0bhtpWocIFC6AX7227Wm
n9hg8Ft+rKA+3GrGLwRrNFP031cCQuUE+Kh7ElzU7bxXdwkSBW9706HzTgaby9Iw
GqzEHM0Do6RTSD2TDPSEiMxqiXaO8btgxxDr6VyMoCa6MFrXIcBtuHuqMJj64nlb
SXIVo+i3CZcifEyuvJ0cTVmAkS2wl3aj6TbvsQkDDRfNBDcFj9bsZIkYps8h6NQ4
cMQJZkmf6Y2oo+zGRjBVZn88hu0th+CgbFh/S/UONzwl2q7MeRLyJzoXQibp2OkU
exsedKTjgvIeNtVVn2nXog+SLbjWHLeIePtomoAdbP9WJ3nyVN1n2lkE4ScsxkFk
S0EX83ybjhsnWMovcNZzEcJ+MS+O9de8PjS5ZdORQYyBYdHgfWKzOIvl2O4ku4aA
r6rZtocpP3P+fKp8gDJ8xmBB6FG+y2nszRiC69f+lxycJCii6sCgTL2TrVLfE+op
z3Qyo/n+oEfi9HjEP3UdNkm/po+lllaql+YXkH3cIQLycdmyTWsLyZI+6KmwRQ7r
i3ApCSCfEKg8IG35Tmcv2UuRgjT1+RXpzN7phrKTeFNXBaJtlZr8lp607QPsJug9
`protect end_protected
