-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
y5X5ZitMnnU6VSn4yTrTKJ091yUBYKdPizJ71Z0GIIDuo3/C5YQkl+aqFjXVwGkUTlDQif+IyiyZ
069fzZ9qSQQ7iJc4ZNtZxhlbkhPPgcWgIQjHELmuvt2sWchMWzE3Rr//MUqJSEtJpeS9Ave3Ss+t
3WVEFHieRfX/UafJAmaD1gsfj0wkADaWedNJ3i96xKtrIev19KnpxxJy4j8vd0x0fr5qbtnchUCY
Rr2WCBj3QXltK1ErBnRo1Kh5xB5vU1mV5fo6Gt5HxX/+h2l0nYx3rhSguOzxkHTV74QXZqm8cVWI
0d0wpsLniBVtuxhkShsZ9Fxwrx8uWUn8Q0zQpQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 34496)
`protect data_block
ot9RAGBm7lpQU5KOlDRZDy01EDSEO1BJr2KFNS5JNu9xd9B9v67Hf4fQ5PSKeMb+WSp/UHcdy8fy
q+pW3rJHU/l7P8FS6CCKFrbJb81THJB/0v+5EQxx9Ne0EkOxHsxMTl4PVTDggp2CbjtYzxvU+MDq
bNfH2wz/Z9d8jBBzcaj5/NY9S5E4ltQKjgUtfBubdHYrC48aeVteBTj0mbNIFD24dGdbvmKGT3dp
CXoYRwy+Aphlb5HAWVv9ixZGYR9xzddNfJhnec82DlgO57i8bXLcHXlwfXTeJgfL5i3gG55FdqZ9
pRkOlDTsLqc4HWAzxcd+qYpRmlAk9vsL1NRTDoUfAXbq4nqFRX+c4Z84c7wnl9N8Nm0xp5UN143x
bPiczfwYyBVkoYiJWciE14dYLGWM9I+SNZy7/QD+3xlv4ok/5FKyaNWOXUY8tMeZ0rTG8RaU4fqv
kMQrXY9VEmYAcPXudrobx5opyZD2qfPxrBnBn3YfVn1zTpfftmdBBAcrcMDmwCMWJsa+hCZnyVPb
UW4/EACzn7MQ5q1eY3bA0yh5dTZEoC9NJsWMxYflVhwv0s1SRkyqHLdfXXS23m6PbAn2Nce4MPHT
YFbRuyi1n0YRWLlwYQdoD0A44xxjBQJSGQh+fP+U6mPUC3U6TP9glmTsBaWWmJP/sWZWau+ilnuL
Y2Ti/aKD6CW0+gMTOAWka2MDMtptDcLvOgLoCkJYcL3iORvUsWy/CTe7I6sJCzNb2FhwDktpuVBx
9/njAXzQipTNuIEjXQxkQO95RrQFJ35X5ZGs7ZKkx/Jmk4LYPjV25nORkx2mdt1fL25mSA64Gc73
mtmdFxd1pxWO1qVGseZAgRlWGrKS1OuyWzGReKZZL1ppZ/b7V1G9zYVFCadzYtyTDGHyQpBuHsg4
7w9uzKpbl3tBHcxfbJuHq3in6UuWlddRSXOTz00Uy8v0aHS5fNqPedQKwC+oc9NtfWPEKt4k6W/e
y2X0U0dwDxxfDNJT3bvPPBFi/cCTlLX/zjfqNyfOX9RjpVqJoq9Iztw/ej1PF59nS3UL9xRyGvka
XFSCu/yFH7LlD7Nb8VEnXJSq1Ps9VohUkQwykEWlY9bjzuDC2RB/VmCSP7BGnZa8A4iunHbAbWhe
1SC02NrG4X8ebmwNwz20XiwN4pSKm2XXiwwFaxhs+dHDF7j0ITxHBbQD6f+8+Q2JEShv3LOGajoD
cJBG8xV+eckc5xPvmYBTJh5yJZw1cXjPmsKaJodObBc7M0BLacSMrvQM/anupxIj2kJ5A204LEKb
sOODEQ6A/yJY/9HTznBejBcMD5IKwBKaAzM77WgZznzRj037U8bjvGEJg10WwJtUov7Uq4cXZGx1
lGc4FJjaC3dZZotetONGDKzQWqPQtx8C1+hWekVC7lYe8IHfwtdYHZCSfOEGyPipZt2w3ts7Lm9Q
stEOdZof59siZwSSmxSsDiIOQQdmfA7WjK9EeAsf7wl3BG059stuq5Zi0/KZU+owpuc2qdNsFRdM
oWDmNOL+NgygiUaSzXZouVweVWAe6SuUsWMQEP8ynLDHF338h+kKXwJ26FGes+2sjlIwIp4eS9ug
MxijltNh2AHMX7iRnxHLjcBuUDpygsj1P7W3whhOB1ODd5fECYuniQohyoAT2gA2pRndARtSGXAQ
EqmSFLWoqSNxcj+P0iSoYlbznTPeWRkmf6o9R7wwexlucBeZWEReX2Z+knbrnYTN5UZ8XAVkbozh
rvIszaufS1E0fAzbyhmDPp2jAYswzdP60lljT6psPKPkov7FQxaBs4tNmBBQLss74KHWwsIVFmds
CmHgeBBy/H1mgO80PoRkfBkbcEPQG4JgPfvp8b2G2hbYKCH8pyC6/hD74WD8ulvDHTwFxTgFZrTV
Q0H4wW2q1eRCFT4iACKqTLidNSlxWYHqsw7EdGQs5bfUkc7y0FF1WNbwUqlj0EYkkXjudethMwfZ
xMMgbJvpxUgZjf+kx2txOx3UgW3LU8sk9MhUP1nw5U58T+uII7AkaZ2EtiLowI3VON8ovKbmnfVy
0pZSuW1fUly9DV+zgH5ISrue3nP3VRcLjXFEnbxngm6JE/RiHwFeQkN24U5s0b6V5RvSly4TfBrd
XtvOh4uhI0jCa/ErL+aACzhVpyNbAZaiO7LCpsVw+QYXSBPD/LviXVaRPL84lqQI+yrk4nhw6TCV
e4UptSIfZjSQYqB4hTu3EOt2YjdZTeT+Y2l771c7A4QZcZc/SanwhPBkb0Zo2jSyEJSJnIV78wez
syneN9jER7GL9x98lL0Foxi/XTeIj+PwKX4PqGpdhUlGDkzjJD7ag4MldeZizjbRsm3Jmh/lXSUC
FcvLtzAOrq8Yfg//TN9QA8O5aRIV0V6Fk2aEjsD2KgDhZZ5akw2JbfHzjk6Qk/nYvn0N9toadxzd
NYD6Y+5sPeOKKWYrJLsmn+iheOn90zvnIa/MkX6xiBQVgFMb2Z0B6V1H9Wp9YWSh+TOwYaEuD+5n
V+20aVS7eTo+g0EhNi2rjGe8t3ijvIokSJfpK3+9+Og5OAVHmOrT1h58zmt8BUQfbnRayveogE1u
YviOmrrvTnxt5WUMv+cPBFjdpn1Uy79FjP+2hZn5O2tKEOHt04YZz7d064S+Po4kcdCezbbDhOJ2
9621hFClABel90EO2BJs+afGCzDZx3g/EZ75jB/HVyziI/UY9+RMrh4uogFrrvGNOVzwdc+kEq2R
9ec5tEpJZshlSFU9EVueA/oFevv1Yvh+DsaCre7z7cqZGjpiSv80x0hjB4xGSPMeAE3Uvn5NitZY
LkiwSezv5BQae/Y9ZLkX30YKkqykGS+lsd0DmB4mQCsSmn+A4//bBGN/EGNTFnP9bl1ArDsAPA1S
+Y0DVZk3VutDbhjYp6NjEW+Haj8D+hvnR52cfGrs7jhxskN1L8mQmbS56qKeJj6EF/4QEuTCXnhg
lQhsC0MiTv3/I6ykitx4iL6sdCSWZ6cny2im0iTxBHKq6gAsamORvNZS0nqJUU6no72B9AQaOd1h
64A9HMHL5SwJR3u224N+eDpicgW3/4kIaMFLZxNbB8UA5j3p+cwsMNu8amGmAX47+Zg3RHpX0F1w
d6S/rKw+kSN0U7D1Xv/nL/wcjPG6tEkwkoyRLNxAhAyWlGi4IwHSIrmMsjYz0jaijARbiKwDPKb7
QzKUMrjJGDNrEdxCbN1TTPI5JX4Q6KMxl+RElvpMShUfXTJmPpyfMkAlVK5UQxXHCpxCXma6R/MP
CFbIsRO/Zo+PqfFV0DN8tdsC1+0oh80wi8Of2RDp8eoMNT1juxA68fefajyBX8z1t813JDShnx+D
FxGPbSm6KMO1qdlsEf7PMxadB/WN6ii1k6RkciTQcp5ldrEc1sSJoAQmiqTNUpXQVyh0U7NHJuhl
P3pB9HTfmqWM1YSdBmnl7jrNPAqigVSp5mRwH6WmZJkHwDfHhCi8qouBE6sw2xFR0tAGECdT5BPE
eoAc0gYmCL6oWjE9cXNRiVs7dG4baSWZ7F4g1Yg2vBY7PgtSrCjO7ggbZh+TZC0Dg+f55j7py6e3
xGKfERmUFaT29uzdGO4yUGQYZmCoMux7JI795WfCk7NHdOw6RU+zu1n0rIA9EJC5wQvWjgR7Yfa5
KHH28GqHUegfS9d+htDD+bU5fRdFXePcxjbQxR8tr1PlS+kVhGQmzifuyh+ECmptEU/pOVe5tirH
5eLda5FE4BwJCtxSH+iYaRqbIOIrZeLIfu3FI03ZLv27wZj2AYvyZ2ThG2g0/+vf5ccaH/nHI/wS
NVqxhszbCo7FCcT6e1GqsYArfi4UQVCyj5qdSClqcj5rCREXhwB2+YI3jdPp98ue7PAX+DaBi4Xu
/v4KIpjWt9ynbUtsLVL2ihczT+0HVK07xYUF79x4YkSgFIpNrBJvDzIKfJBTcE6WXojjwgsJr+MU
it7twO4J9bU4qmcIVHSJZgQ05tHgePyifuq4206sdcntzcIRyUqUP/FFD3cR+TJsBCg/S7dw6jd6
AfFpdFKbqTefBi9yU8He1nb80Cc86gwnJbL2LCFhp7QUlNg9LZh6MwmhRBgI5CqjICcLBU3B30jx
w8M07kiSFNmXNQnEXVEAl/FEOC3KncQvy8f76HZ8nXTOSjKMcO1m8aN4xC9WuhkqQ0Q1Cs8cG5BP
ZVX0ZPf59SsSGEyBAjhp5fhAdOx1EnoeUvdB0rdZrjsno3qZs8FWYTlD9mlmFx5ytQzVIsp7VOHz
uiT+vunxSR625s4towxNOIwgo2L5l59okIGol5Fs0nDbD4hfeb4rYPoMBeYXzjHhZXsfbmxoNs/v
5GRwy3IYVDLr5i7FfUaRthTzY8d5RW1zueH7AcpRgj4mHo0Zcy0Wy5JVhydsOVqpG7DJYhAeKFwq
3iR/8/asOsn4b8bKsY4q27pgHq/R7gvF2K8EHki9RT80F+xh4p9Yr5QCAyNHBxxY2t62+0vmGfg1
F30rwCT03kp2/NPtm9Ud1ZYbWo1MZh/91BSq1WkwUwsKqFVtk/JR4b0B3U7g9gnF5qGN9SBFu8DJ
ItvtP0aFGpOG2ldq4luMylhT2TXqP4aVjaNSBqiYdenjaAAxzTAxSZmm/8gfCUqv7Gy8GLXepT2n
ujrf/wz0uoyHptfdip2l6odzgfeOaMjIeQ1XFls2tJWANLgz76MnlhUw1f1uSlTk86Eb5Pq0+ZYI
tTGPtRRGuMNgww2lqUhKN4jV7ns8B9FevxAxlmonsLvKw/qeXEliybAOEERcBR6i7HLy9x9cs/Dg
Et75XGnLHZQv8DKagajy0xL24lpIalc+MlsE+V9/FGNQH1hnJrPnL3/RBDY7BlT+kOSiZkN+i6z7
n5t8YohC2rmy9YLdf7Vid5m74R4ylzZ2dGO0JhFuXzPCEbdv4kIAoXoXtsclh+FsQ9Gg8/u+uK8f
CZ9O+cnC3AepcSxUnGKIOjwBG1sKGVqpeaVAiMk1d1n5hj1wx79oIzENZH8J1rPNjRVDmZHEnqUs
XVP5cVkIfyH8kUKmdTFdFlnvZfB7xUuRuEY3CVZqI66osIuRxLrr9JZVzTGmPUTMBbpgszwQ5TDY
ndMoZRYlXUYjmnRCasd37fhUZh1D+9pqgJkylOGEVpSZrnLbkvYr/gaBMmcIWIqNcLIxEeVEpjc3
lJxr3TCX6gwfmMdVeNW8SE9F+jz27mKlgwu5elf3uhut4nOqvUVT+NFTB6SPpNBd1F+XwXEjwQ3D
Zsvcb3Hq7yBf2oaqwGbwJm3gnf/UVFGrnWWEfZo8pIB41lRfuZWjDUK7e9epUmTLfItZjLoJST6o
7wVnBdzjihdR5n13AsGPXyfdsaSJGdX14P9KHErCNXiIzzcgt66kToClvQQazFmuimZ3R/XgVbdc
hmRtGg92Md2iNnjs6iR9nqZJznqH7ssq8ubgSZWu4wj6vDo9Fjm7viLd8YkphJ0EmKjQL9VQF8MN
WtJ9TjxuwtdhvYtNCLjnWXGKkWzmL1tLzpmsbMGRMM0xuAj5N0RN2DT457gNf1X76cu0ZmoIp+Rz
x7y0/bqm0VsNTzqXQnTqvLfig/gY4AS1Ovlmi6+RtfidaJBZ8tVN6oxLhJhV6XK1Me78KT/JqOf8
f6A9XPgj0Hu/OuTfjWFV7E2nfvtErNhUACr3GNoivXBEeqnn/MF4KgTSsOlYEa44THP6YcSyVdo3
mBUItZBnFXOpHxcBuLZz5wEyyrxTRJMOJ4rYjGKheThlu7pYC+KUt2CAS9IzUhiBKXBGB/qygXfT
8HEboHvrNs4oIRjbr523mkMnlk6dtbAQImNAv/PdUZ3Ivh3iz625HeTnrRo6yGtD7PCS77YvVCGO
dKZZfnLoCvJFjB2VxYdwainb0pKHzrDZtdpwoh4R8Ej67xEmLao6f48+VOHhg+B2h7M9O6Sv2FHT
4qa6RnHrqdRn0rK8ZRlmkgS45VEfxiEkqSBfEWKSCf8O12QUctpIdwyYjfPSUZBRt0KvW7FkoPk1
DqzFpq/AD3wrO8+BHLilUey5GnFkCnMXLkofEsiKVOsV/9RL73n7FtVvZ0N6e06e59crGE3YOPDZ
1gXEGwr9t/GRpi8WfIi1JnzlRLaMZafBmTOkDaf4PmoIOij///UaYUHNsearUhQrB8VVzfDSog/d
bPDvMxF+wD39DmbU/reFMV4s/R8YG/ccrakI+sEfDD7v3Tn86kyjiEyVOpmVPifVxbjP1ih/s7Zu
wfG6H6ot76hXPvFzJKBNL0nDyKIvxDo/fkzz6GHRdKAjiMlho/IjCYm8YaGX2EahKa8QxKlS9hDK
hssK3YFHxM/IiHBivLsZuNdjZESvGZQsXblamhTNuR8TO2U4rEoFCYyZgdjUAkkfo/rd8Jo/h5S3
rdQhNhprwoqRcB17JKpYTiQIvGr8GAIptew2wCNF1cPbizA5ag+5UWQ+9/6w8/r+AmiHzd5CeHBz
/a/IueOoJfSiyUegistBG+Co2KZz8y1EWzPyviV7D9oDqGe0vEglWuAdPXtCVNUSJ6PJBJo+wZYz
jatlkPxmAcMQT4ZbASBHf76ViDtzt6I8WlKuZPvlmpTfkjKBgUgmMyIvvLE+ISCilkphnbs82akk
dZx7HF7RBOlnjOpiBfQv27gVr/natd0QGADG99DrGDp/ZygGXFH9ThSTVCCoL1IsIxL1PQhtIvQq
kdD6U3/miH+nZvULwaKu6VhQvylVqNoXAbo1F6MkCbySVPjDbFJRUrLATTBAEsTUxDUibD2jPnvV
Hww4xAz7aMGXvNu02YheUcML+us+l8QcXFpz7re5mNe06p5Iovg6oAoIhWX/QjFjJ3cpIxJOANv2
7pe5hs78Z4+De5557/aC7XgkwdY89T0HtCO4rSX5suDcp4+yMlyNZ6ZnS2Ic0siSBDBjiIIGV6hx
cHeaT4/MnO1HYDk1NIwo3ABSuuW+Ebqb8UPw1NFnlsg9rlb33FWlSNZ7MgOmh0xyzN8JEhJiHroP
o/KpnafaU6fB8eWhQQ+eize25a4Y4CLnu5tNGI2uw6e10oyB25XxWfFE8yucXR97FGe5/Hd5xBWw
aAEI9JP7RKBb2qzn/xbmsPvJ9J49Hxt0mMafT67/DB9F5nXbXRXzZ+APscflOj+DOv8K8+QNDifH
p2hC6V4ayPETCCw2jEtpz/3EGquQA/HIWE28p45o9k38+dYAKzYw9bar6q85ThEI27RJJj+oG8hG
+sH9ALRb4SWgMR5ZWP2dfxoFAQB+DjUId6tZ0VM2gIsA6EYNrDCsCMYro0DCJcwPl0TzRgCvoW2g
njW5jMBtJSSLO9JPhvdLeDfiV8Cn0eKPBSUHD018D/hIxHR10yNZGuwAtNGGvRCb4768Kf96pAdT
OsO2DmnQFPh2bwA+5a+nzDqZfN9W+eMqxyxAcjrZoN81iSRF2H7BZc/SZDSThEiY15GB/tj0M6I5
ljyykrHhgArWu1bgyhEsDnZglVsCKby/i/0nxsr67aluplMIu5SI8XrAwgTTooEgesJZ7++o7EJi
aX5Bnm2avr/h7HztDKpti/OL7GAmlHCtitKl9k6HM+sKq4qjlpaE3Z4rGlhMsyCG2BI7w4xywUUm
n3FDm66JCnQ707L78ENsxSSi2Fy8y/3CrgjtuGn8NjxkAtIatAqi89fEQXaUsqic2kPLfhCBiOmK
H+9bW0Iq5LJVjrciJ/7QuV5u8GfaVvuL2tTXTdBKclhFr47jopuzxYLpottBVRN5wdJbn3Q2Ekyp
ylZvM4Mf0fW4niw0sCNAhBnI+Z/FM8/I5ArpxgVCn8KPE4F1qQHLPuHBJ57t8Npzt6StChHlK61l
q4P3L9EoLyeOKbQyAijLRitRD6UMcGoF4KO33cHmIN71K9RyK2m6VCbotXtgs2f4AoYreSjhapBK
SGMyvSA1ihcWkWLtBp2QoJpFbIlplKlP6i38PjdrgNRtSvmzQCEmoGWd1nFeKAl2bWGIp/PQBcMn
yzdEGgqVaCbq1mc8XAWWKkJZTz9KIfIrEfl0vrTrfc/xD+fWqyeEQZ2Y/lcOXfMWHKMSqglcm/T4
BVEVGHRkce7I4o9K+ZGiZmqkIxtVaP5MMUSeghquUn1B03Q3dszYbZwunQ+NyFIf7SlkR6BsGHX7
MseGcFWpPP0WwCGdYDUKDeirKkDIM88/MnnXFoMgrNtVCIhwiVuWtfp7RKqk3XMpEjMdmcPaV6A8
X5H5+2FldLcnOLRJnKlwOMWrXYy94YB2rIVgJg8AuPC2fNZzipd3/dsnA+aD0ZJUcTcAfOEbaJYk
/LNsAMXy0h0H+wfVUHsJJatQft2EY3p4BiJhd4a8psI8ww0Q/FOKFY44Vnzo9mVAH2OI6xTrhKHo
p39bO8R6nT8hfGiDRvm5MjpjCW2vV1rtnKMLkjBIXXMSBrzuchW1UP/vmWQTzVVR0hMQzi9BY9GL
+Lzns5nVrx6P3PQe4VtUpbDn0jgeni8vreIG3by0eBc5rc20Rml5HVm1tDhEO9xnIlrQCcYOcto2
vD+mk4v/aNtQmEspEsf2S91oYLl2ZVnYdmrPHUk4XA2pKmGsnGN8hoD0LjMi69YLOYKIvuJ3OE68
IvHF2+zRFsPDTKii+cWi+2NMTwjP+euyg/5OasJ03zHcuk3cVok6SAC7KTkJAfKhtgA0rmbgHEnL
/wBmW4T7fcEcZz78j9ZCqBfmUobQJhguqSl5veG3wXG/cFQCaqyKOcVfKmJQQj0GSpywbDe9JQKm
S96TJQQm6VY39Zao2naBPlsi9H+s8IGA2Gwl65qQDzqu5pRQOkQ9jTxOJz9HbIA18nPeNCEA6Vps
wO9UfdS8/Oz9r7vKm1T4DCX/sd7af/48rbB6nQVw09U/diBb8538da/ZytmNpcEghSmcltF0B53t
3PbRQZjM9xnvDY+QlDGLxeT5zSB8uJk2CNIev73JYmrgF6f/xLY+Kjffofx0O5x9JtGoQqUPUVjA
PsA14G9M8H0mMZZd9BrLOSQqVGPbcBz8JyH1d8M3iz++xQ+TZIfl2wuRimj3fkN+Z6zzQu23DZla
WDULHu46aiG1wjJIpiPpmbAZFl3On/ZUMafHX244GvzNJoLFyYG7piSSVKOrlniVs9+WuqZEPC9r
mviHuq9Cfga3drxOLY+matefZQNZGCJwzjeYjOIgA1qEx5Intjc9lEojhxcVRgUCqxjHXV/xwRs7
tLwmvZQ36uaB1UhSR0ouwCGvBrDXNCwOO/6luW8X3S/ERsS/c3jWwGkYghli97M6Wfq2/SosAVSI
+JF7MFO4X9SicXfuz5zS8sRAoTgV4+hJh2JIxEKXyEy6dj/67jDyBxNmGVZAIq5W8ntCX2gdRdRh
D7v2vaT0yOpQv247d332qomVRx35WjvrlHqqap7b2PohuJNeEQMceBVNB4fOLUcu7XOWzu5zmx6j
L8Ug/aqhP0XdemUtBjJ2cz4NmkmgAH8RR0/VZKImgcuoo3DtNNNYtA8o4fXOBcxEXE16PYSJjqfn
cwQLzvg3s50MEDGvE8/bs7VOJtuC/cnZwAHzvro73Gvk7T9fBz2FrBNk+z3Q8+5JjFmixbwDPsWH
Ml8MX/c5klyAitBPyC0vAPT2TMp6oDwBv4necFQRlSMrbFEZbox3Td4Dv7t7zAipyengMjrpgGjP
/uNJViZNmiJxk0g4CSEN3dyO7wJHWLhuR67TMpvhBVW628j/v3sSNsw3/8g73j/PYN4vJWO3yNR4
CuqyhUKn9gwtPlbiGk0+irlkz+5pC1nsInk7GTx0EHqpqWwVVq6wGk4GucoPi4ej77NMbnD9euFM
Tl5aOhI9F19eVi3ehF/OFbrABajg4+G3u8uDAzDdZvT8Zy+ZjJytBLZG0uY0stbYtlcix2OQpJTM
F+5cyxyrO5NlTq0Ja7f6klCkgXhv20mtakClkZn0wLgWWSQIDYY/GZE8NWivTI78g/UNupnNshdl
aeYhY/5H1K4B9gI+5eI4fodgVrh0bPK7woGgOAH+ou03COH5e4vw/H+jhsRhkq0Rxx87ayIZYpKD
gyxmqHX/vyjGeLgUo8ooAUpV2SfyGZ91VjyxlSpilGT6jYvRd+A2thHjBHQR8Se8ahdeLa3SCpnu
sBMQJ4tPc+XFBJ4bqIgA9qRDdbhlNtCo1chb3WJ/Xq8GmdI1/U2F/fsjRs3YciKD+gRHpU1KM9KQ
W6ferQAd+cyC9QtVgEgxY6IUUYnjSpLPvgaJIGoo1DsbZYktBWa6c/0RyxfD9nqsclol/w+DSDjE
R/m5YoBQyqUrPURBRebvr8PT0N9wdxa+NAYRVzXFsXKbMB1t4Wjs1tfaXQ8NUjpQKNXD2MtEkcHy
CAwSJdRA/2ApBqNmxyCYZNGW6sl99bnLtU+FNlfQXzbKmWj/InFE+IKd2x5m933V7114D4W85swt
vnXQW4Heh6Byt1RfPfah0sD2AfOnKORnT3DmWk82MUoDh7z1PN/+F69bvPvVqpCtF5dtrp/pQcWY
f3TyKigGKz/9RbbXHk8y4OIECyrrI3QQ0FOt32aaSCQQYKBc39nvWgiKApUlhrjXWYoqe5Kg0zFY
zD8cM0mkpQHroaPZ+R6klc/8fFPLY36iuF6zKLRS9CFswwAJEQk7151mUNk4cBSI503+BCi1+MeO
XXvRvdkgZWTDgVwLo9S1RY1184gsBJsfNsI3GTWotpGHGyw9Y/qp4hinX2ABwcr1vL3TTJHAd8iJ
z1l5aSlvk76+xqyxy3LApOD26GWzdPmFmReGt//Spf2EpciGwQ1domnSsbisgzAl9JwBBEyI0b/I
yw33OpO6AysXo9sD9b+K5gWGRzOJ46czjKgC2WOIU1ESHgnzS/wyGz9fFmyjCpocXJfremH6rJ82
nBuD4O7Mf70xR/miovpHQOwvrdOGbiK2vlYjNRNG0Q+Sx+4ZG05DP2l4dN6XS2BU2vCUzUwO0Hbp
0YC3dHgb8ecwcXIqryc+RtBZOnClK+8PL35ro+T1nydHSq2oIJnlTWI6d/e8YKcPRW1aCzX3r439
lxmBqWUldHgErVt5DSyRV699yMjaeXO4d4YPXYo8dyFwBCo+ZB3YXt3UPtbDo7jBzAdlrrz2uN76
bFHqItPf1iJQvQ0Ucy2VU70iG9cBYN45zJMufBCGE6BtXCarEBbfg8dEqSZAoYGVw0LxkSaowsFo
WWFfcqVVDz8ZdrhgCsxn/v7Oi5c1F2HqCD07ChvdO3ZozHU5HHz4VnLVJIExZ812GbDaCT4tRpmG
D0OwmsZP2mU1w+TdvEncJp+oWlx2ZFU5D6+jvSR2YLMeO9ukstFDhMWDd6crtOhl9Dm7/QbqiNSq
kaGD3sqTApMcU+HbAimZsGkP0DF8GRf6Rx6iuvRQtiwwvM+i68mjEMg/pfx7YRH0cVkccfBkR1IY
kYt4u6x5zRgspq7m+Qrokt4Mmd2dyQ0UNjwESUYAbbcrjuNSD2OONL5sEri6TEte1efkQ8kY6kK1
kpgBjPC+a/mmxtxahc5G0yhrraxMKP9lEI44CMp0hV4FYydMTbpGjq74lTN+agqQC0XAkP7MUvkp
CjVkMfe7up9dNE6qTkS1q9HOealMXQWvMS32sNMnphfo2eY2nTTyVZaQd0iUa/hpTLwJ6PAJjSge
AZluUS7IMCq8hPLHxhIavroS53pPmMwOlljHMirAAPtcQawMgdIS7w25mgZY2zV8LvDKNms0qoBC
u0V9PCPTVYGedpCmajCIC9IDcryvwOPOlZzrm5o7tXPCyRIpYNk/a4QvYdJDQ2ZrdBIjFnHGK0v2
htBGhAJObTZuHnfip+tqTPeNG+sdZkW7wJ0FxpHVB2nnbTu9OKmoh1+XllGFjzYYS7CA4edO6xGc
xxP3CnmXlTeElwa9zH6TXZEg27f9cxLzXN7j7+L6bQyq4fi6qHWkQ4Qe5aBfitPuFoxFv7sQ83k5
r3Roh408ZoXEyEA9REciGaYd2zlVWvawW2YgtpmHxChmk35HtvIxK2oGlWMfYB+PQqe5SasToQuP
I/W4kYvOJb13oQUlKm9HAszCfxgkmaVHDj4zqqfl5R9N0bdf0yH/OxCoxUQOQpWgS9XJyoKufdIu
G9BM2YdGlsvWxVpI70D3cvkprBvJvQWiVxVwhGO9GNzXuY2IAOJqgduPzjbWxGhRtSI1mO6zlc9G
7UKrtnvFR4Y2752rSYp41GCaC2ZPUuZhapc81VoO8M3LEw8wDl0L8JeoRL+tEv4bsVlwE7GvpEH+
1cnzTprc561mM5HQF2kruozCdw1og0R5XCkwPet3RtrNSA2FC8w8oAC4u4cK77VKJbzGrqDZ8wos
RemgrE1EycUtojLTPQiKTlNsnnAZHHUOPZ7j/aRfUbl74i1NydWd4yCrDc2WmIdTAVRA3xTZXnkx
hhiSxNztAUcnOOgSO3oJE2kwRSv6s4JC49cJ2qwmFRPAjwmNKloFHzE1bfdTBR6O3LLDiJo2gcSS
s2HpoRMxJZwxyIsXIbDK6iNpQnaZrixQTUQJYPuu9eVGD80MH0w1MV7IVxTu8W28GbsP8ccYu/hg
g3aRq5Fm1DoXPhAev4uknx7HlzzGmGhR1gdGJlm+PxulC8La/V8TzNFxBwAT37QR0yY5gBDPN+9R
On/7b1CEYR78zernOQeZri+is3b0Ao/2c9eVXJn3yOpQsf8ZbRYhBXIi05iyc87QvsbaDLN9Zvr2
NVCjWQN07w46WPsjtHII7zdS7BZ5ZVEheiuZm2bZvoGbb+wXedSctiB1X7Qob50gOql0T6xEzFBT
n1rAyQW15ZpWIBsafV20BhPgwEgcbHnb0yRfimDzKIW/M7olHA5kw1BP5Ge151g8grEASRtsyC9R
A3R+IQQ2DS1CHzi3K0FHkIbqZSZtvTu6tjBI3hJf+F17mfX2f3ZBtbO6qn6r6awvpJ7sfDdMdO88
4hVTIdA+OpoTQOkXfGD457NueE7REyzrqdgz15kDf/Gkf0iAGe1ZdJx1IdsNRqPFRYxbtZmTmE7i
1nnSN9iLUCabCW0reotc43rwQ+ittonoSE81DXz4NkEQnndSuM1qB9GuCPYQcyedqBxaehLS4lhy
ajWJyNZASDBZfBzN9wEgZuYcI2YOb4Jb18BWf+COxNhcxFUKRUGsVIQDfveEuThzCTHg91C0Zg/b
CLBaHtrKbe4ha2NQuttU0cKvQkfUi8Dd3Y9BUDdiZDwEXIDieft2o0D8sgW9Kwx4szz7OXQLSNj5
x1KL8tTggu/ZCsSx1vls7vy0D3TqoVb2xNx20eYNCQiq31mh0At84GSVUdJL1yPQO4VpjfD94Cit
2HGssjSZz3YvPInG8kj/0Q/w6blGs+6tYVkFCrYYGmJ4b4LEXRKj4b2TYqkGlwmpZJxsF6MwF+P2
Mhyly6iUKe8anY9WnTXrK51DThOih2mvvfSHgEWyMIMEMWNHmGsmqYLt04sRCTQGx/w0dOwEJi6z
UquS6WQ7X8QtLSwEpd0R/nDMmSEhJHjGEc7Gm4XjAZJmeWnkp57AMU2fQ3WRYWNBgiLXHQ02flI4
txWsGGxWLr/Eq0+9UbUk3z5svTvTVSXWdVkLpREYhxVtXGppx6iKhoX4JmDQQQ+hcvnnZ5231fAh
z9hXO+B4nLbDx3D2ACSspz/zgsMwb4ZzQYpHWex1uU+7sOm+cYsmsHa/ofT8ji+DHxAlSbDIHVMr
gi6Uyq4kmqGCaLgz46gcHaW46LCMCInWMyVDFMvnBWgMcG/PizsdIExlMGr4vpMRweLV8H53pAG5
nKH+KkqIf2xjPwmwDmg3XLLSHnpZHQGeZIDs1soBmGdNXpHprCEhHWOEqoxZt3d99DExaEP//PRW
R/VLohULClFKqnb8QjgjCVJO8xY7j1H6wj82gHhf2jWzmdc7YnfdBqnkquVcJ5QKMz6Jtd97c7ii
H/KWfSmyvBaKwgfF2d9rDUu3JuII1fTqnyzCSafB55cD9wkqjH8km8we7CQAc5kSW2s6508OnS3R
/feMAwSF3t4CvCSGtTBzmpBZIFyQx25q+qrYyq+JYSi8nBsivmrAi/wkectbZ42RG0NmYRPIKVsO
tjocNAej+yy/2W7pAdNj7JGYM7rz85aKyh/yN0KBNF+WuShrpxIJaj8J40UViaCkHYHpvn7tPzJP
CknLKHva3TRyqpDpWbBiBcha/rOzQ7jZ+Srg2udaC/ACXun8hKgy8NVcIoLSMpasE2KB60d6feLn
oVDrhIRIjKblb16A3s+XG1PF5TZK5mQ1Scx2pA2ldHHPxXsaqFiUwDhqO4XyqwofmY89xpNRIMgB
aiDtFHY8gmTK6i2PLEZ6g/AhnrJQZH4OGpiYsrSQPbUN91kJg/LZtdGq1i3eFPOjNzJv521+W6DJ
IDXjkncaW3r1TZ4NPN3uzX85dVyDcMjx22g8VO7tNspIwvQTXhnP3Q8ZAKufveLMVqpvl+X46zIy
TLSjNYM2efc6pbfb/hjth+EtPnXic/tRxUqVuHWebVwhTTUd239lk7YlKHxWVBh+Y3Dxz3YfNYID
i2778WO9BxH4XBcu2s+45SQL3qDE10Kn+OC20ztwa3Moebm1vCq7WCDZ5/gAxleIvGYaP1beVyfs
l56Q48XTMsv6PWahyFUFuqBIPmqhxToLc2Uhv93Ev+NFJrFxUD8HprA6yg5RT4Bu7ioxn7IfbJGs
MxqmC6wc/s6cw3SiM95D95TVnkfwRqBvm/pvgV4l5aAoEnZKqB0qTeedT538sLBBeTkoUcZXy6+T
tbbbLe3uPvZBbGy41OFpStEfcJjim6X8DI9MEqKwVozFP+YYihvXtUVmftxBFZTahMnaAMab7Ahj
cUb5s2gIb3U5DzmoYB4wKMqvELF3aUNurRGHX6lay1wOsA7ogkSFHAULih6bePKpDRU4kyOMesIY
w0L8V4y/48iO+lW9cSE/O6FYdL0T4CIECICN6O1rxEh2k4pS+idmp1xGra0/z1as4gl4sjHT4cgi
OwRnTZUnImPmtHPrQ2JFbNynJUAAYCs3tdJ4bdO1Q+OSL7/tLcKNmAh87TE3I5b+cKztkAobOcCT
YFGLgl1iYkyzYPIds/Fn1DHuNaFnYJ0atwnZwmdV9xs9BWE9DU4TbfzVQT4X2TWG6n2Ba1K3ioyk
noEgBcacH/spP96jMNID2PgH3S0+GTR0b+7F6Ss8pR39EY3Rq+/WFleXY7B8rCmgST1NFSdWPn2q
yDBANpwvpEc8tAQW/bLeQ8wPwdXYBO48IMVHPyKX5ZrKzPef4aCQ7npiqllD+rt7GonLMhgA2Aq5
edUDzgjkKnf8/WMM64LC0HclEMZwWC52PqawEl8QgE21oU53ePhvlc7IQFccGB90dZJXx1R2XYkc
BQYPpRulB6t9/cnV9os11eA1BI7jQ2XCWEO/adGPzBva/FCA3Qhrnk7XqvLzkB82225kipJuo0G0
0WsUxD4Ov/s6f0z+eMH2dnnjKFRqdXBIbskrNZo8fSItVU723t9cUMGd1f3lVtFYmPQexfLoPn9H
qGTTGPZXWooO/msCcL3SviuuixCmq/Aeal66Xf4Hdzcwh5wEcmA8cxnTOqSeC+cxURiBtEMskSPn
N9EfeqdnZOLwjjCExemYwU3d27toH0V3k637p8Q+fEMSw0I71+govFNx7n0YX7BmWwEo+diZLAfe
GUs6vj81dnoq/5xLTJ/rY9/F6skMFrxLjJttXHNyz9VfEJMda/TTUnhZ4srwy77dy5EGefHCbg0C
PYQfrizTnYQ4YCu6cRYYx/5ZdQQoUToMk4kAWaVEomL2TuwaYU95h6gYNF7rI6lOH7/uQPApD/IP
pLdJMi/ArAdxd23Gcj7rMWhih43Ux6H7EYJYWKH3NCw6n6ST+7m8cpMHr5TKoWEJIMc1QLLbWkvd
qp5+lDRcAPIqsicG9Ql6Y1wSnQMCP+291JHSG0KMxosQcNYqdXRd6Z8qFgaAtd8KyTDHGKwICoj/
GROy74giJRSqQ0jS0a6tmKOT7zbt1Ti+xQGPOk5nj7pCwQDxGaDSj+m5f68w1ayeLPcEsaMCA9s6
0hH8jpu0hn8LNMjd9nHKdZQB/+1w51hevF5p1wjFO334je5C26skdNWpv8PaKooKftdVbIqxHHoE
Sqs91irhH8/krhEVdAMBfNko9U31mXiQKaL5TJjBLQg/jrPDLrVNJu3Fmooo+eBgauTir4yQRvun
X+RaYxZGSklZH6eTYwSsDgGtrFIhzb65avWsbNQjl8DcrheWPME5IBuZa6AA1e4o7yawFvCR/rG8
x0aZyc7r6n49IbJDE23VQAL76XzMU5gTN7M2FiGpw0xuJqgu1SikJBQ8GnWvUw4FBKcPFin9eJpb
xtkh5ZICniwUMvOYX/E4H0k95uUkP9iIdzvVwElT6tCLqlSYKrdt4eNrOuvcr8l6Q0IhKsgSpobE
tzpvzBZ5Tp+dGjXM8k6+OxfNDm2NDvSTvvlNVpL5cTeoKgn8edX5XniQD67pqoysSl6E+06bn2XU
V1KMq4tyKTCuLSgyOM/bXo8ke5qat1ZOGjvtew8z9SIaURbEGBpuG4BqFDZRpC9FJAy4ndOfJM0G
mJt5y+zKPwXz/g96hoHXi5BpFHxr0zMHaKd2INoysRj9SLtZtwp4NkcSHYhLRGR7eBiFF71b2T6z
J42sfBKvwY24sTP8pNoXQEb2n/10PIVobg6DdGvqG5qCE1kY1Vl/La5UFjbeuN0RWrH70N17UR+a
5MI54WQFiPTPXnFncWQP2u/x4K9fXvRZAU+sYXZ41DP7r3Exul83P0/tIWstFi91vaOjgKt0hek6
fN+hEsMN+OdQoTdZSnAfbs/DPn/SgEhex8XJv3J4ADCjMzMRzaTp6Th5Y9j+flC1e+sk/6k39Mil
uS72B/U6CDcdqGvt0P7nPF/gygzsxeNeyKrLKXd4MMVOVddSD/rWoFCg8UzgYo044t3EcP9Ijwpo
7ftVOe8VJsUaC+275/4jeNdgWFR58RxyGUuKppV2L2RjniDZ6S8S4LJlWFKsx2kGTUnRzDBeYs8W
K/CLVGiwXPHsTMKXy1M14XHVqIIVhAgkKUVv9TVCDqCeh6tdI51JXnE3h2H5Ur0AdZpLfHd6n+5H
jUyyXd3NMTx2d6lxOthZRxmDsCgcxJaNsnp8STG4bT/iNhjz0GU++WDylnnWMEtH/lLLUphB2/x0
o1iituHThuwRgWUFM06kxXYzl8FNuYgMB+3To0szp/sTV/HhnNBIoBzPVJ2yNHUh1eskDXr53ttw
OQQ+T7b7qXwxzbm2CR0ea2sQ/9QEiwNhrwSygeywo02gRPkzoSRv/vMjpzOdpyypuixSI8k75f20
yS+N7fdtveIker02CC+AjOuDX+xviEunikkwcNb+QJv38P4w7xRBP/Yd8D3GcVn2HXaze1URoj/P
SNGJ8PzLXIL+yMm3EAT7DKcqdrWxVkulcbm/DoCuZqw/P0EyoM0/kXs9Ud8QgTXuK92xAGhi4wja
o0gyXJ+j8M0Cgpz1Jlj1Gut2r5FiXYfj+okEj8TR8/tMbnMtIG3ocymfGS9rBoVkAVEpGkuPV1jn
tbepWL2byhd8T4U3VN2HKp7Z6X0wN/38dst8poNxDMlW+WEKjOH7ae+gFDenZkWgudj691hhm/lD
fKdS4bl+GDu9yXTCXckFfwES2Iyu/7kc9md/qe2cEG7BJEM2sQLAY4/Uqrr2FZKg6/vpBHBqN3sF
uvPHdGErFWILJLsXfZvno5LY9M8DSJGKJrVT0qG0xQj7Vyh4JRjeQ6Mgm9AgZylGiOKh3DqpJMVC
o83/xgCxBMGuMjH0dTRb773P4OsOxsDKcTWb7Z1rhDe6WDndZ6N5I3d4C/agCdI6ocsWTWISDdwH
GqPsHtwkCz2tHxAIkj//2DJ4FgAYIM1/3bOCszA7x4ROylzEvz6Bz/HZHVmz2OpeZVXKCOAIc8AE
+5SDX11Dp5Hx43IQ9vGaUmB00Kr62rc0f3YiD29yBLfdxGgieeXizIG1aKNzr5MDv5lDIs7KiCr8
OWsSPySBVk00zgrAxHA2B4SMlVg5/Ni21+L9r519397Wa2+nXu5/vk3t/cfHQ8NrSVIpwlu803iD
dSjeYiFXFtLXuRnUCMcRPYEcyE8Br7GuGB25tbC4DqY4N6txPeI9tSKQel9YBwos2sKwg1zUHdYS
FJr0emjLw+Ke5VoKqggptVLX1ZA5cb6vYQbCYkCJd+TeIxoS2G9+3QI/HYvuOxnuDoR9SD3rKQxG
8PFvrHGZvjLnRJNKmYDcEIKSmyTnr2TD4aDscPqZmxFrNVrl+YkTDHS0CSAFTy58Tx7SXDidaaAk
FQ77bn2ZWlezcvG/orDybdBzIUHVh16CfkKxGPhhiVxGDS3QPB1UKyVEJfqibqdDE3EOz6ox53Up
fz3H5DeDEbJNZjP9LHaohlhY76KP6EvWwHwtThfFrFGcoIGl2su+hxJabfrZ2puofAfhGoxmApsy
9Vrt86UnlH2rRo32znnGW2OC5LpBwknbMn9U+6qe4t1jFwf9h3LXM6xQT7Hf6fi7tqTNg07tzLcw
r8GWQSOmjH8RPm3727GkrgVYp5P2057J+QwzeEIK8Lon9LBcY8W5YqobMAEG7M5Vnvd/iYacBhpR
Yu9vQq9jbVZRMZmlbXC/GpTUMYZHMTFROTRZQwzPssZmM3LnwqutALnkThTTr9FKMqFnOgWpEO3/
KN5RvljWDArwzPrD3qza7ZfLKDhcYK9K/i8z1IjWYDMvLaOrNexLKgxf06bI2hcBHBz1wMsd5A5h
4PIVm5kxRLHd/u7a/34vdbvKXNths5kLkF92yMRUhxqjK6db1D0MYecUmb+EklPVslHwcXy0d0qE
vIo1qA5tQoFjvqcKJxS0lMc6N5cqoNnBUaX+TRt5833HZXArHsB68jWe8SmyvjGClpYIIuJUrybo
pwtYAlpScuIrhX0pligpwHRPiGp2xfhoJufynw0L3W3JfXLf5gib+ADjTIRycefhLS/ur5HkcOMK
/dcjofEO26YorRQHX8btqaeF9t/hmWvU9sev1hI7/R/F3A4EvWLndwENaLNf9HyyUqnS7aRJ/74u
iyJE63rZsG2oszkeaSiHLOF1DpgArcbr1DEcwwc1/0uXIQirtUMOIEzfI4ukoSTnSlxT2kcU3vB6
rlVl5dV8ld2TqH1TNUSq2hHfs9domdS/FyWSZa2++LeW91TF6r7dZHCMrCH9qJd1vzK4idwYNf3Y
N3/jmuFxUj4blE84RHZuHIDN1biNgHG2yJVIIM0SVfPRXEwXs0Eut1EorKvPDv8gLWRi/J344DCL
JmwVkh6HnEXlrYAr/n1Ez3nHgkuqvLyvzoMbZxvOKBtDCw7MT2lDZ5rS2r6Drdm3psQRaDmwsiyj
SPLdl1rZJP0s/Yec7Yx194GCVElLu2Qs+Fd67t0Tp8n1xgVKp0DBgg4ZaT8WpmLWsZ4oF6+QrXMg
YpO78A7Mqqa6KxqLyrDzXw7QbTKK8JfmGSPQwJjX7I+Y46cYb6niw3sMMXpeoQb8QDjm98lR7FEf
FEJ//fqklYdyZ/JhLYwxoitxd1XoueNJ+mQoNboXr+nHcZ3SrRTyJdn45p9M63fdm4Y9vEMZd7VP
PV8nmCZcZv+50Q8OPFx8j/3w4+OzScVHOBH5IY1zn5TktrWK/KzbZOjWvTcxvCzq7xdfyRsK5+db
Dhvwvz9vrVKOOZQIs6pTeW81M5+FKB1VfLmHRZaLMsZ0K2kp33PYF11l3ZWmOVUT4fHDpxX9CfVb
1ibnmjadQdrd/NaPYCUAOApnvAikmGtTUYLhzB+fMnvpNTZPSncYo8w1337UgvsWZL+oKASOQZ+V
/KZ/fyxNaKCEZvQDdrUWoxEHMWRTNUg8dnPwfwW9XxDpSECOpR6ZKQSJ2Kj+B2PeyQLVotzys7GL
35pN8dokxucs/jYwWg30LJ8yt8IjkbrX+kVv/bkjGzoVk0hnWwpHqOQsbR6NRj0l2WEJ+g+6yire
26UvPhy84Kif/XFPGCZ6XgUXV7hzW1vce7n91zgYe511QBiVWHY66Ec0JXFiUIWnzbTLBvDO2egq
Fu4ubTc7YZUw6+AxLANrDz/9vNZN0NFhjfZt+XjYRD6hbpXRF6VX3F6N91iI39+5vwpWe701cd4o
0z9azN1keTkoAZtpOduo7B1L3sbmPVlabbVkhq7xBLQz+CW4/AMW5+9FTBRozn2vBX3hcA+LP8C7
HwXkWpur+FXWyoJJOixBO+OoXmwauf9W+NeMCGH/qzV/qoBPgf07Q7dGs4dW9+mxhLJTJIlxZjzt
IVKzd5p89cBxIZ7yLT6Aoix7ESTRQDiPRF0xSd2xmIYOWaSFIm5grBVopiXjvCMQySmppvUc5hvO
TigfP97zFNNmPHdeLxcYj/1gwB2FSvO5z+L+mWDPD4dvlGD7og/nTaRJMkpH5WwE0IgZaLzOqxH8
CVyLFEoah2OtBBEPoIm0cbkj/xc+AaPPtZsr/52aWw9PwmqYaULe48v/9GP1umAJzx7oUXxtdfKE
wU3HeZp3oIwDgqhq5ObSVQj7sSh4mvxJtt/gJQRa+kfTNKCE6OtRxCpHRcrcG3xB2rlq5T2O2HV3
TvjyF1ZOLEwY4+eIAqLEqk5B1oORanCQZLZiCny/nxVOOEHxEs72eyeUdIFx2Dypa/VmcvLYCiIa
fleBt3RkOPaiduT2uHwmS5kLVYFOMcX6071QvhThjePNjqhHUyQvzDReV2MEB885E0JqiU05l0fE
plauYYMlCv1r/WPgz9jucQmPWseY8H+DXyt8aJm7Ka+S/7exOBmnorKgszLhddS57lHnDPUK0K6j
dUmxEL3EKkcHu83+ITfuRGFsafs2rxXxLHXIIY2IWH4t6x4ET7GpmpQrcLlsJ6brdgGcV61wHDLK
SqZzwkMHzSagDJQy+GWfasxMlxSFw4d0Idq2XY2Qf877iyeoqRzZpTqW3E7BXpUCbVKsOoYy4/Pa
SFCNPyU/ErmvHyfPMGgHXEusK1JfZh8hTwigORGWDwSDv+4aA+x+jQm7XTkLTvZH4MifceQOXmel
ORkpkkwrKfo7zeHQcZ0mX1cSoWeX2fD+0Yp3kRxqUJXK9iC0z4+i39RICUbCFHZizBcWsk8WhJiV
V5rFYbdRVcZ1kx99QgSrbUAfPSAv4yFcJmXOwiPEHBn2PXrsy+3meCnb/uE5W5ACJlRQTissFCiy
urOzL30AMhnN/fDiXRVRnxDSffv9hwhqLavGyqKhSBmBgtcG0RpLBnW5OALIoP0OhcknlIXBdHwq
0DyDtWpc9QBZKJI3j0WBpHgkEXMtvuw82AjlI2UGREZdAScuh888zQgeyFPosrFIGBh+cd/vEm12
K4+Z+c5VxINgQIUakcSmMwIhHCNh3ApwT4mWGuoG/Nh364cXQKyj688CspM0vpPJAouty0Z5teW8
jBAOIKl58wZLWAw5ZmidC1k2H26GspCgi+4CDRI5/1Q5AedX5VLeRVj1U+JZDRqfMQgWPuor02/0
o8ft2qhemAj50sYmO/2bYbEr+OkIxhaCm7KdBBsjMncY2qRcL+bAf8bgOfh/PxmoGPcVibw88zp4
yqfmSmcGdrpdBmGqORQ1iDNPcfya2F1N0Jh3An+XaLBXatBXgo1c2TmQzzRCbZAvMESOBwV1vzIX
WI2XDMgmBaIOsFEzPr6ra7FmNAAfQAk7B5QSdhg4iyr3AUjn072pgDeRTSgQSCRFSjd1DMsuDukH
fyMVS7zwrroOV0ukDeEpUhmpkO29fyZIfTRFFAlcQ5/95BZwhukFN4lSj287El9vrY7yCxSAv2d+
4ms7ORhuPCWVgnLc+jyGn21uKb3iXtfGauXI834VmPFW2Tt9hTALVkZH5fMAC63Dx8SORu5muW95
2+gxci1SwB1/iCSlN9NmkgVZMSAfWCgDG6oYKmOB5AM1z2HW+BfT74cVWjxfPvIEq8LFep+jdywu
sQCSo83y/8Gicf3RdTSHzy+E5MbTZyv9XJdJKoLVOMNgKfAlzrlOpz5OKVnu7WjUe1A84zbcgOgW
9aIUiPgBYdFgSypoK5eCHB0b8O4kZKQO8XeMBKR29uVdMjRHgUuc8tYbRdQdm9UMMLvZOgSVF9Ev
ShYsRwQ3q40Yd8sbsnXm44GxoGte6+5wzFWyRfQiSTsRtuGq8uXh8Ndivpr49O2bONJZup7Yrqnn
7BExYhatlxrVa5w6Mfq++jngQo28+dpdGBAy7qlVT0XdEp72xp3PBN5BdNvQXvP8hR4QbINbiWNr
DGFVyV2qFiRwudp5OmAo/cyca4D48Ktfvu6A8ttDZsjBm466vcvj+leINh3qGK/0OvrhV43tvtcB
T8gbufSZtR67LYdnTyUfSehnW5FfUd52BARPUwBgvlDPa43g3TygfGphdb4nBNO0EV/tgpY8qXy4
uZOdD9VGgFkjzaI/m9miLt5K/iAfUhCi4SeoHH8dI4l02mIfdKF9wOtBuM+lqmw7dTjqu5ao6lnE
rD18KgmZUnb1rUjYpirLaHdZEB6LQ27WVuhx1mQrVQfDt+KmMLJW+/CVIUl8lKG0ZcahPjdx6LEL
ObVFxXLxVV+dIVmtYOfUCmHGBvqPHQwsqs8HD+IgflE3ljtQD09agYjN2W78/xX/wiUI+QateKv6
1VxittPgNnH0P7E8lEjiSt5tuLn7ZwAs9j7oAfkAYwGhILvHXCfgkifLBxPXMNHE+CXHar7l+dvS
sPuziRsxA+21N1OEWqH59PS1cCUZy1+kPqmDK9hyL6LgnZ599YYc8EOoxMU6sw6RDctbrSxdylQr
C7XFaAKdkkDQueKQh6/eiAQZsk9cjd17np6bbpooGz6RlXfVlgQXk9dRzBwOzZBP+lv68mfG16QD
ivW5Xi03Klwt23XibZQehnRYwXDQ0IhC3OYSbJ98WspHKiV0qDtD7sXg+5XuLOfoaJE9yX8LY0wx
OxpCIlMySzMnSCQ/kJY2TaALWGRrWMmTMWoBBRE2s7QSJrdJeTS6iG3Q6iMLyFit3OKT70FgBmmn
Vc3K0eTFleq/YYhC+1CFKiadzZBRw7AC1n8C5mVfHHrd9bTVfLlzftcn3PNLfl9lsT9BhxViOQzR
rPEICmQjptA1QQRbMM9wivKZHubLT+WaLXXpCxI8rziedTzBpmnKuiXm6qbXrHqLF68ShgptCVwo
5hfqTtGMWWwbwvFXztInHg9RhDCsSG5qXrrLoIgdFJmas5nWUOGEbrJkxGoZOvQNgzNIzTTBHRfq
eEtHPfr7/x9gbpR0rYlCEvL9rOniL9q6RUMA5VSKe5uLjSxfnGtnzp2bSeFKIVWnGJRydgBvMhji
FUEngU9DaHE+NW1vzCw9k0o7KyO7amcNbV2lCumUSrCN3DbDMCWPMil/myFJlh9l/FZ9ieG28pys
L7loeO8wOm65ndFM4gybU89INwvku1uAhVZq+sWmR+fOksDF8SkW78u23bJyr8Wm6XZDJROwKlKm
wf7990qkMrL+wqiZvFj6vSTaMnrKoIuih37Du4wpaMSgvKo/n4OSuQelpMdYh3BVE9BYo4MOmVOu
cUzHGku0HRbpJa//R/XOO2wCZJeaolIGSiWIvZm4ykpnnJ03oF1rCrSC1OXWptqAIaKyhllB2Ijo
rDiOPAhpVjiuSaJJBIrxhE00STvHvPZBZDn7O17oQPSb+otdFiGMpN467ypX4qtWfaPIatNro6F1
dT573sKPOfNfmcgU6csbSERblTQKCBa2pDUmhQAeRMImvTQ+cv03vrAdD6PKFWaKWiMiOzWa7xaO
ul3Klu1JPP0PkGADOrQHHzTw5iepkwVgnoswRKorUG63VRdrupI1QRB70ZGibmavI+M1u/CtRFs6
zN55tVWzhBuySkLrOIip+dsCpK/C8kcROAS0F1pIpqWFfg/aNiiNw7h1Eqjuz9iyx712+t6KxEyo
dhnFKnzjpEHq+psmK/dVG3voySeb0yYPaon685CaiBzHZWuKr7uZrVPzOZXlX3aqxOWrLrlPt/ng
kIwNXbGBkXadIiLM5RDa81xF4e3eZ3AL5BlfIMSIhqk8OcsrzgT019Gi7ycfrWKMrP/idOYNCyVp
R40pTvgvJuZf24O/iCEqVLlcdHXiej8bk4Mdc+1PsZmZ7i8URBuBfYXhGKWcUvQUwMFe/jAPAtma
UXDORljou6+PuRLbwGK+6/0QmBVz+7PDE/OS1+fIV6QvNQG3CI8try/UGEKTZdc7rQiedK2azoqr
jPw6YD5Jb6H4AKXuu/fpzcTHym4Lxaj3h0jXCmKWGEF1T5X7Bdvl0b+DIlTjPEHfPnc1RtSSZNTf
zXb4Bfj5Y+GOtWRHAXZQ5Ft2ZOKKuO/pqhv3z12wXxI1qQDAQcVOqhYZq6nMmwLd4o6uybyAPbtU
bQw+BwalB6CEM3JuEYUdUD8yDWzEXpMmjjZwBajE30dyuVyHyWv4aWB8BHb4Pl7snpF3fSTg5Vsv
B80XBD4TOT1XhxP3Avz6zLVQDxAltJIXtlkGSn9Y/dw8CvapzQaxLNyR3nPA3wNwdp1mY6bu4+T9
S38M9VihATwwleOZ0cUzEC16ZDUQTyIl8Wgcv3uoFf725VUeTLa/bLlVUcuKt9O0lWkWzGksbCTA
Na6ZnOy7lpgBWkfSpFkAhYDT+5mVmxsH1Am/zScKw13MMeSjfXDkGT1eP8KVFkfPEbkT8tCBuKJk
AKDexY4dO8eRO6p5SCOwKlSDkEZs0xXI337FCjpkpn4hSdhhVVfwOh/LSMVAOm3yM3ADDMqLQ8H2
9HRv7J87uubiwdo0eAKKfzwtXq4roKRErP1IRZTOtl5yCBOXuAxOlv975pYqNNvni8xwW7a9vxDh
rTz+y3ikle5Zw3RkPbAIkbw1v1nmXSgTWzsUDvjo1h+I6NC8aMmt7kkKy99TmWATI4/X6Zzy6nfI
CLjG5FzjyFz7WGwMW7e6RAkw5KHbQmu1jhKUP4oXdOr+Y6LT6fSkAbthCCNJkLEz+3PjP/OsDzKW
yUVuEpHxp4tyNlwzIfvfv/iCsTzV+VXtogyQqzykbUrb4jkzxRHlOMEFFq/XZ3Oacx3h8l2NpnM6
qpELveB6OUSbyzZChGoWr8lEHr/qRNOsQSHctwJpk4D7P+qxtvcsV+jqNih24VBcIhWOscV0Iir7
WQI9AzN5788b2uV0HJKamGDAfIfdDRSdVJTDBIy51/j3TuU8s/XFLPsXN8pevnbDCjyXnq3Umw/6
mKXy6otbbYlMIBp2Ahs0OoQ43C5CJmBwlMVHw6/yUFsFdftQeeTLOKm30+1UuADlq6f+OB1czUI4
LkSGoLx9QA2jY5oSMSRdzCN26tdAMV2L1WiOL05xhu4NBOzlmo9fX3u+8a9urVTSr1Rd9JIk0PRL
I7UDthFFZbNVd5lNgf7PyqJpf5mf2gyExC8GY46i5CgM29pxr00FqKn35I0j1NArKKU1sv4PFO+u
RHYxp16eXHGh2EJwFfb2a+RQ82d0QJBrNxTR/LWRCfvXZj/NnoNBWFBptgsqbwxXZhoqusi61yhP
diEP0RK7Cg9deeL5FtAiGP3ni3bkunKeGEhF199k0OyCJnN6UrxfbTTZy8OR0D4scoXm6YoNa6m3
eMWtMKc0a0iPgNKuQwOsmTCWpPaTg1Hs3YgIakfFvu+UuGL5Euw12iSFm4UVHk8h43VAGkbxELvS
rbDoAwPw6CgtMtao7famJCroW9Po3f0he8U5drJJkUNEXv9b+p4/YtWrN/VUHhopGA1w/1s1BZ+h
lYt0gZ6US0Bx9aOnHU5CN6xWrlKh66OBN9csv1+qQiT6asYnxGnECwIyiivrDWhQBCxGFSGhxatN
XLnXsL3KcSSiAsqp9WDmaaR3n1CA9s1VheZKzKUxbZ3brcMJL5jBlWrfxwSeak1SSj63MwsscOfk
inBfhZmipl7o6JZXyHmkh3l3qchZrP/MHpeFfLT61s0Y2Iw907HspFWrq17tnXEKfNmvcLmiLIUt
eD8lcnrcWnBjv4zk8grWucsDRUVJ5zxDuovWU+dMF6feq2S99OBie0PoKpK2s8pN/b1WrIhdBRnd
UvyPdzn0/if2Qthw/ZYKqM+OQWja71F4h9ncBgw6yqv7WNozaX5Lv/1IyWCoG67qPBfQhAMkjOY6
S6XrFfHwej0cGSJRT9DBIqxVqPmhtSg+wJ59DoofEyopcmCxBZGD6HNhT6hlvHUHPuDxvKcoW09f
wtsaBfHC8RpHxh17KUY87u4Gma2GDJ2ywihn0NTYFr7OKzKt/HNM+FeeY1Xgcb862HX6ykDZhTK6
eNamRahvgXFpWU3GzQn+8OIkO1AVnN4+dD8YxTS1P4tMEKkbAyWtef3oDWkse0uRT7rh5J9dy0B0
d2YofMYoHpr7JFPPyM8Msjadf3RUC03WuQKs9/aUSPb1iKhuBoS+yaUXKpQJ0bHRvSuod042Ewzi
9iKDcRkgl061khtJnzwKwAoS5HhQqPMy0mb8DQqzeWRYdBqX1g2e6TkhYstB7O8BrFXp6yl/iLZn
1NeaFn86wf3jkOVwp2j8m46zHJypzphBLZUpRGEkwpuEx6e1wHUaHASLlsz+9CAn9v6Xc531tnZ+
KOn1BwbZ+kPGKwAGiJfcnH01Hk6JgV64t8Z9Y0sgEGsWZpwgaVBZ3eQ2h8ZRGHS346V9uUGu9wUT
Ntk4EC128Q9MJa/F5pti73ZXRXs3FFYgqCpywL9VCoyQUtjkFaiyjikKNN8yHXdrMl1YXbijZRs+
CXnyS0wQVUzzzZqKkoSIwQyuHUuX/oMTlxtHUPNvU1HqIplxE5DrkaXa2yQKOmtrNi/1N+Pyia5L
ihBtxplY3F8QofrxOoYNtqBRrPNmg33gFVo1NqibB0LR5MszeXVh6+vTNYUiVSQNbq/T6b08NVef
bzGwZKuBwlrIy1pYxVuUMx6v4RS9b+VnFPNSOkVQZTOIXKCSj+sadluAg4RJUSPfDN9CGi4BC7IU
hPsCYfc+dIFsglT1hsu2UmCipydRWALWWnjNE7syglmcEqy9CL0+Zp1h8IcUUHF0p4vhEc2KbGVG
CpmdbLeq4BQsUqFO0BPXDBXOgujcXf6kwzEcNlRgoK115yhz1QZ7rJC0UJTpfp5Pdlq+XiMqhiEE
lolUkx9YxS5uBeboI4nl+oTcjDR2fxRXCH00CV8SwmNCcGE66mOzEQPwIHPNPp/D7fMIP8K4NceS
4wygp+POowp/mXSNNbmq+uiLQnzSLDjVn/v+gl5/U9932BwwIlaz6TjAtwSfmwsGUOza/YaysfST
NkboGL76r79TSx8hDUDiQLfHc3AIIpt6T04wUGuyR6hdmF5NT6L+cWadn8kGqCuomoOt5CbDutMV
8fFe4buFvTgcE76+qo1StJI99fjElytkBEQ8sDTrVPi3yiF2xaZ0D5KIuBp5/teMwq8U52dhCw8P
cEI74d8glFg+cB6IftR3+VOpHuwGWL50CFrAZyPCSmsCQ2BBRzgCgpxJEtT5IS/MBl0X12esY92l
qX4hd0BQGd0oEW4GLTR1pDI4BlS7DhKpEKMgb6zYOC8CG7x8KFxjw4SJ2LO/3Kv6TLPIUZWyBJ83
S91m9B0Pr1bD0GTLc93WjMQJLEcqu/NQk4t+Mtxlsd1B/NZPocHmIANlXXMvgsFDWa/RBa8Y8gvw
pQ0fxqH5m3eSnhfRlBcbAakptuFzSEp/QUzJ4hod+KTnaQUyTuAXA6Kuxh4D8MgHs13OqkXoTk7/
mcB8/WZcC6YHXjREulAC6ZFhFiZy6gG4fuqVkzcvpaNqRMiJgE6si2ggsPdj6UBMKy1MZSYipIpA
k2kjNTntfJdrXikYHghuIkDekB1CmZkDUlFH1v9ekqdtwHi25NGTBBRYI334FAZ31vdcFoKHbqxn
kBPhML1oQS2WGITxbId2qsmwTkPs0FI5hgBcXjBk49RBBm5KqzKIO9pJQpFKoxgICWV2aD8gf8ll
0xVrzdqVhrfc7/8q+ayqBgIpNIYJpAXw6AXSMEp3Gyp35pJWfvMqgpE+J23Y54o5SN1Uc2MXPc1d
gaEy/0yE4ozS1ZIH2/ujM8dab0tmJ0Vw+HCA/OHVURnNpOxKZAoPtf789FFMlIxr1uzrKAhDyP/5
geB57kxXuNSfjLzmeNYPhtYTRZ+BFRm6AamlEcAsTkaLZqJnX732loh3kzD1R8cD8pOedJwGgyqs
nn+fEmaw6QVPyG+6VIgjMRJZ8QMSvdZqHW+Gg0pn+jWoYnlqapHQcvTXrX1RpyvfaLGqIJLR9Hj+
czowa+l1mg/R/Dome3kTTHMbTZ5CNEj+e6gGJZpcmO98Xfx64qouSAMOKWqazCKmh1LNH51Q6wPl
AxIXiHXvgVcAassOUyQkPDJ3zz/QcHx4PD8CUSY9HzU5y6rRtHhysqFD/x14zkigLJMR4MxC3THT
HuXR3xuPrEK+97J3LF9fJ6oxEU9MAAqPhMOQIq6b0anR3AyHVFBs0B304jZ/7Jtea0FaorTkMc6G
BaP5F3tDHUAAiHjkcywqPkBMSU23Xlabi27vcwXrFHVzu4IpzyPEA8wvKEU7055R3O6vJK22NhUK
YuWt1Pf2H6sCaWWeiKw1v7/0I8P7d1dnF1nlXERKgZRXlie/eKAAuuFGW8REVHCPLzTSGyOQ6F6C
+F07VxMJSwJ8RG2G41s5752/Y8+tkZwH0hkOJ7SYqehIGkFOnNxd2FcizarFWEvkwGsex0L40Z1k
PQLcOSwLWAHp/UuJ1fU+5BL6mGU56KLgowpDvIgbYmoSD2p62GHdaMZnuRLb9MaCVlz+9Kw2N+lA
cSnqwFdNpiYEyQf/XMyiDKwAk9r/AmHyep50sQnwjsFIhbgkmwgx/5Fu6ZonaY7vcWbPuGTN86O1
PbDwGL021+6SSEjeJ1AsUJogwXSF9Fnvyl5HCarsETT6KNov1Oru8nOymOaGKEOyq8rxX/GZ+Mzm
HFEyLYcvQpt7E5C92jYsYQ8xnAjibBVuWPKcTXX7GS7oBW4WOFAAoft6xiFudQX/FkRBl8QjbQSO
L8lQvK5upr6uG9VWnnCHkQorRY03tfOaNualjELayWfr32w/jLLpZcAkedKwSVWouK/WiLIRPHQ2
fX+GhuGqi+xcIK90uvwmIIZfOzmYiUrA4fa/kj28S5LsGF0IJVCXsJH206sLERKU4hOPs4YkGAzJ
fFUnKkVB2AsWZPq8/Jycjg7rJsJIMfo6MhIh9G6gU8UMQtFpWtTDNXyGhjIvkD4w4zdLIhHUoAVh
dE5jO6nnUnwwpu41b9dv6p/I2jIHghEfiez+mLfDyE6PGIIEtLzsTwgj3aBl6eaFnYxGVk/IcJX8
t+NAEz5TubsqRjXFkjgaWlg5cUJIS17OOypqsKVMnxj56/C3y+PlIhKaGwl1rUHsUrmlMNU3yIgt
2odwsAufdH9i8R+NKrbNmV7x9MOJxZEDRRoFW/0N6iIUvC+yDQxHTuyk2U/adVY77vbC3/jqlb1P
pdux43mtVy3RK4D5Og28OpNGTDQCtMqbbzdcEfmNwSmM4ZZLlyqPGE+UV9TWTyR6TiR0FnQKPIWM
HXs5FY4baCZCDzJ/szFcFEDjQqd/pFtMeNMFXtcVGLtZhXB3JKFwZ44+qtAHelfAryYhATHYWFyE
R220QwPGS7ypHZ7+yJUYfJF2cQzr0fQT3SywL1sqw2PqkDcDlbKRkJcz4CBloR3YRP6kJjCZIWXB
vbbVK8SkXJRAC9Qf0OiP4XmUK8R2CiPNMXR4nSgd1n0CZL1i7hs77VNvTEBRRhnxwoF6kaufAYwY
V07ejJHwQ4/i9gBFyPU1UnIrDXnkSYplz72pwPcuGl/LptIRta/FRGM591pK8Sf06xCqyQ/S0LRg
4h6Y/vdMevmuHBdPp3n+h/fE5FJ/qhEq2kronaIH1rAn6Q+lNRfXEBH2qVYVaS7qO6E7cut8QeFc
jS5yw2z2WV5YGcGSX3kRsbrvoWF1mBA8sgcY7oW9U7EHXK0UQYmOc2cU8/a9WebwL8oDA0ydRE0M
bwR2TsJs/84eiGQQJMgGd3UvdAcczM8lIchjGXHGfoGP5tXcOA2ukVoU2ZFAUkC8jP6fytxiyvEH
aUi8Pi0kcxUB/M2nQHcEMpuk1emIcQmTwmAGAsklyOCQg/G+ER1JTN4mClbaiD+K62XuhgNKeYVP
H7skdMo6tgf1pT++mw1yDm7z/a/BagAjjUMlws1kEYRjqWqESwynpIi40aV8JYPIPruDqXZA193r
/JARrF/go2UKcB1gixVgq87qiwIS+mV6I324graxKmlkD5n1JSSvP//M+eoRln4cCXhx6aU1cPUx
YViSWBrb1r6MXrCCzL25ozwsRy9lXZILATn9xk8nLGMIj4sANfTEZqUOAxoMZgyZG0IDawOSZW4V
7reHGEvR1OuAP5cO9BsbkJfyyCOL+BlCTeeFjcW9HChmi3MLjM+Luhx7HRUnP1+cNhcE+BxqyXZw
jTrak7eCF7CEuz0lPCqLBymu5eez/ai27K7ywgbjc+xHgsdsprYjB7pl6Ls/DWkh6s8tltnJS7bf
3qgzKR92Qs0N+5MBFCAfbGwvuVwloaKCKhCjtNMrpxNnSZ8TW9O09DfNgQoc3E4SnqCVDXV22nDU
sb9xrawDHtboGT7zAPvuCNPfcef/X2sH1WFSDFTPMI1Rlq7ky3HjQtsGwrai9Jq91dAA0IkOT3Ni
C4yaoZGoicDBv/lVQlny4d9vo4TvHcitUYA9tNzi5q1VsOyzPUk7e67dybBaIL75LA8NAXqprU3t
+puOW4kt8Nph4KjRZBJvy/tt6VskuLeuBFpS0ZHKAa7zSuaV/e6XQDKH57tmUJFKXflu4fIoSnfW
6OYGjrY5F4DRzmHp9CfTBiy7GU0dzXrxJ2vRmGXUpA6b6us8FEt9gnF0VaU3jDMyoWDB4sRSgPnl
hHdPfk/5eW084hZWgLwT0Wr5hYLSUGdpghTBOOCydFyAbesgjoTRkTHVVCQhBIznwFAlB2IReHJR
q1XEFf6VEykzJjHMc3J3mDEuaugr9aFHtayMcZxOiGR3jm+sOr+VNDIN7xWGVImY7CNUeMl7PtG6
9HMOTaOWwyXSeHO5uFUeqBY/JNE1zoUiHmmylVXLx8OQJbIH2MWgqA55UBKZ8T0OrAWvmdhgHf+/
bFE0Z+b1jGHwlHPsjrxp5HArmPYXshPdeQ7ySCo8oIFmOzfrPvNbQeq1OrPa4zwPVc+RntyTIApG
Kca0QT6vO4w4/7MO2ajW7vFXLWJDxCH4S0fY7O0TN8CcP32zPyhrqwfprB0bSYdUmWdXnpU+Jzl8
iKiQUVuC0HHjx4brl9KWRUsIabQFK54C4vvq/AhapyfplGfrZ3KL0iKeWgrNUHW5TpY+eCYuw/4b
XxvFJRdkQT3AfRad+ebQlP903VW4eJB9wYkce2VsU8FHaInBEcnMkcpypW7vXVcpArhbdgjvkOLv
yfw9HFqvST4QiZlR8IlWd1+i8doVt9ttu4upZ5IUBUl+6S0uLUIRTM8SO5+zD0N+JjCzTvMcL3PQ
MrpBD1IF26kJa05GGIJy1nNLLjXUsFdyurOm7KXx6LCkSdo7Ain8Lk5nK2ucqp64dlt3McujYOcR
/WgLyPnD762cIVXZb1BUFIvGtBtNmITEZOxGDhWbBme3T25O3h3OU1J0yRmbSDffAIYLuUpYi3Lt
2HsfIRLjjc3z9a7WziEPjzijhkHLUZz1Z9SxhwI2KDfkFI9agGJszuuPjcInsyfXNqSM0oPf5PvY
hk4By4C1TFvqRg+9cEmh/sMnt5zx/vLlbm/pwJUB/A0aXp0Vg7vG7wtGZSpWOJ8E2qAwEpME+qOT
/qAJk3VGdQqONMgHtri/WhhaHAf2gXtuY3QF72+/8hx2e3gJLF4dfbfeEdqgqoTM/SungwHteGam
/3VkG8lD5ImmJsdrLXkMRYIpQrBXJlmvOOe0n0KXzaWR148B+YUKbJwpkiuITEA+xuilZtC3srLs
G5UiHl+kIIabIjR4ajVw8bo6odOMSjuqiFCrIa3m6Y7Qfd9JyqkhN/UJBWqWsNhvCEz+e3Jqp4O0
/lijWth7XR2LW7dfUtxINzxP1GJsmmqiXgwL7iqLJL2X4mm/G6USSKXxD3lKx3XCOrqgH4TxM0SA
nQ3u/iq9ApHJ6IcyY7KLgeepoWBxJLYUEY+CrZfe//mqNGWzINP+cqrGpzv/aVOIwYwkvi/xq6b/
u7FPnSKejOud7nWfus/CCfeO/QyHIptdciAncbioTK71Z8UJc6JTZvTZn57jItBN/JeadJ8vxpkr
r5E0l6D/ntaAaKz0jyugZSRUsNMNXyJYLktYTcHgkh3DGBjFv5kVpgVV4DVoquMIFKVLt5S9d3Kh
Ok7KiZGhKTU9YwRK2BulbMd4lxocJIssFMKzLoG35SwWdKlX8cGYl6GhwVyAZDQrcfDEHghAIzcM
7EObgw4TCqYqqTcluV44BW2IoPEPMU0xkIuvWFQ/nf8dqVWRZOLpH9TZksjSN9AOGOPT1g0qPies
ukYN1vJ2PtFM/tIuUCHmYja92ElfGkXlqw8e3a79Y/Bhf64JHiJHVwOckxRxMDNzyoyo+jxww0JD
9qBDoODz8JQWbopNInSAMMcF8fg9yUEvcLjHyGIPgYYKMSNOIkhJd4SaviTEdTxTACkwGfzzhBgj
7BQBqEAmX9tuF3YtFfuqPXdQ9deklrYcx609GQ377x1vAC1y3hjnGpHw852mhBMbd4qxVVhDBEpz
g3f37X8TjRYViAksuJGESf1rqw0UCUkOD+2i5CVGqgXMMVouf1Lwk9hVR0AqdWKMi16zp7DhNw6n
rT/NP2uyMz/Av09Cg6wA0yhcqb3+mH0tuwpuulKr8eW9doGvd19k7xu2EheVFmIj2IWm6TLQk/bb
mH4GwChnWu0Oij1lEF/IJmfZULMzlnYvy53GMNHxIjggHmKrirSl/Q/FmGC82mAcHtvGxF5yEaHO
Z8dsCJL4pfeimlr0sBNX4KaiSoUV/pj/1FORBfWWecHT1miwGhr51fbx4GAvtC2ALOI8GHBMLgaG
jJdnkLFb1IHL3v9CepujQLbnoO35IvSbUduBaZuVGWVjk+cPKm/hNAr1d2z4Mv67m8+18HXrhmFZ
fhjTA1epkNbw4+YscPIiI+Ow1sJyiin6w2x/wE9QkgWBZaLhGN66qeBXi4PfzjeKZXMhUIzcZxhg
+Hf7VqPSE8nodDLvKiCNtFvKqIM3qKRHG6Tr25lYsEvG/jQ+gFX0ELGWWwydhG5JbXmProcLUBo/
vkwOZHzRr0AxdvswjbcuouCvRRZnwf04XqxlQWx3RySO1Mr7nyBRdmNoQYDOLVDZfElD8ShuPR/4
y+TApWLkyY9bg34G33CkxSGi2uzi5OKVF1JqTFGXLxOY4WWVt6GaHQ+lakhw8+9LEy/vCcRZY7/J
iYksfCY1h5Izb+ctMHuXhcaVdm7Y+1wRKs+wuUAxi4AKuWhsmrdeGHdA3BRDcz7E1lFGU+nlDQVC
oZAiJ2V+oXpkbs/fioJQBdbvb8m3fmUmf/1eNK5oxpxy1z+TTYI6kzvEOqN+8yJI8p/gOhiRIdbY
Or7lrCMwepQ1G5O15+bL9fbR5HjA/9RPXwx5/Qf89k7CsAiKsZ55bYQ5sxf8BbKidft6OIirn0Tw
SsO95Pb2sr5JnjsyibsHks4W5fAS7oqtDJ/StxstdDMI721g9+LXsgtJPWutnnXQgdikUI8zuXXu
1wenJcLe492wso3ordCtT4M/s5D8uiM56g5abnXLtHLd9Ghv8aDF1Bn0s2JhB/rhZKqsa1FpDaFW
/J3T0uw2y9as6d9tzmtlmOtLQEJefC1r01TqOynPRKUUwls9p9ONplMhXYmNRQM+F5P8pLfFUwtk
68nvT5lB9Iov/F2twaKSyieEO4Z7NJYChH8m6/LOopxv8ubIiHYw6FbjMsqYZBkMH2l2K2ZghBfl
n23XrvpIdDxUGVr+eOdMZe593H6GEpU6NHZ7kRWFjBZiD95mE7hbY+VAX2hWBMpyKT0SKUFmP2Ya
QTHQA/ltETdwBMeFm+9iph4sxAihUJnaBOg/9Yk77iiov3Q7GOPHeChgbThqx3hKztP52Pvi3STg
/gFree32RYa96kqXb6idzkDLlhushvMHS0YOxI6sg/NiElphrzVDNF0sxi2KZPRP2r2Ii8Rt9Zfk
SUS8LV/L0aOAX9SKP+nwFMWM7gXQsra50yXrWEocwKtfREEL3iWHod/xk6DaXUigwjiBQ90PrJEj
2Xwso01irSXZ21aFFDR/6AZ4Rs0x4ctkqpE9DustwF4vSBbrQdNWs/LjsUmjwsnMduTv/30z0d6x
11C9PMGK0efAVtEPajvIt7q21UOeJUL++hmuU6YJfvUhRQARmpApVFnilzzgB+/f3mAOjg6ZUVLK
K8LO0RMhauVDRTpT73jmqOsN8mS1QETTikGXe9Utg+H3UEwaNLF8Gk+HBVp47WhqHtquNkP3S0hd
Jrxq+mTFK09ZXE/adkBt9jFoVtxzKiWYXTFZlc9grY+62gq3RNet8nxXFlY3y2zobZvKJDCIFR+2
5RIbFTaTEDVSg8kNrnUfjnZoHWnXO2KHBTxwf/bcdaK7x+cbmh6QE5MJ1LUjtwvfxRAU3oV6i3/U
WqGba+EdpIH5xoM2WJ0FqNeSrBKl+IOYoxBEBRpxpn+ukXRArCmAHEFXOR1tGRLEYo3He8EHtIGx
Tf5rXwWxIv3xjSab4iBjRcu2HBd/jCB5xelLyYz8PXwKhVnSA5nh2M9stagxE0UU3s0Ff56EW7mf
ptWe944eyQ8VKsB/kVlJu/F8eU3lnwvcukGba9MDAwKO5dlM7spfbZtIW53a8kvChZQ2WvVbitYI
QcZkZzW6ra93CiX7gg4ijvIo+uk/4Xa2/kkw/x/HTOvyMl4/5fSXszqa9IeTDi4Cfm+B5o3PCQfk
1P5Z810i39GqjRVmMkvDjlvbYD5+yBXBDE5nkLDzJTwSZt5T1BSD6KGe5gWK6gqQCOl1g87pw5DT
KUX7oYZw0Yz4FOcDxBXWDcl9788xSpqm9NCPb8nApC2tNa6w4kJvDl0U6hQJVloTjevVFssZCcoD
S9t/fMokHJQuMTocHgZhnohTh+gAtelxWOvLNGft7VYlGpdgtLWr//bzbinLwsQ8o87jSVmIdEQH
Ik6DL5AxwacDggUUaVL9zSQGoOEFIfr2BMb6lOGOHgga5+3IzbH/w2r6YxXREcCjvW4zu44wGLNu
vtzPQGJ7hEGfKudXttEbm787Ak+F3Xrs52lfLC5FTSDobD0v9Dmxl6AcazyMha/4BxTlSyOV4fKH
9dDMonTrfHESgZgUH9KLCsm1e8NPHcJ45UxhyJrErM5NPHgWLFQ2TXQuILKRl1fABc5dW6aO8u37
OSq9D0e8/Cn3BP8cHV6ob6vDzeATkYC+SZZhJ+xUYrxIfwZ/PouVe6o9w5t4I4J+xHbbSSA79a/+
aWnE+MR4VfhN2hB7YTJ2RYgUHMmgrLOUWrgpderOQO0VFxFpQLdgtxmdsy6seB6D7QWcZJQ+h0kY
rjZOZQcvEzTOgQGxW/BBIyDljoRTT0ApaZgesoYcDvQoQvo24IKFOAudQUplPg9m7MjMgXZ0SiAs
2+0CVq695IEckDEmxIVJgJ1E5wbq+9sicQiheQR83xTk0vFarDsx2uJUda7mTLtBCFnwVZpuPmwQ
Ua08GyDLaf45naujWU7lhjfmAsYDzghUvYG7v1SuMUsKUfU27CetADTSQp+0lrYnXc4ejSApqII0
2q3WdJKOsbFqUezeTA3OyRnh60vf8def9yndlZIPwtdgSJqlXvNvs3C9quwAHhaXuin4m01zRsi6
iTPHztdPI50lymm2JQl2ydQ9W+8pOVeV+Ciai9M3QzRI2iQwu0eExGu/OcunN2YHNgJvjEZbHKdR
WLsiuxKIMb/d+52dA0hSzMVFha3HMF9QBSA9dxEjfuOPFxY4XyXCv2GgokFjhKXHGxi1pOxgV12X
DGAFFDe7BuNc04ytXbQWx+Gf60v2ggAn/IPkJfnWTLwiYAsjBdLvuG8TT6QY42c9dSVK/+TXHRA+
CY2aTvkRzr3JXv00MVMssAZEUqU5toLsFdnfOcnUUrE7ZqcyMbBB5j+rOisduVVuqIqRnT1fGQDu
MF2I1nm3UDBp0tDj0mpGUHviIC+F/cc76LXOHiK/+OEInHdnMMYhRkDYdvV2wFeZ/N4VaKOejhTL
rpDzKeGrOg5aB8Cls9MaSwWzbgc6ONig6C/1VaSw7F3VmWSrUODwNGbhRBc86KQVWmVvRrPqtzrd
T7dd/exAEw9nnY0v1Y87I4fMZj7yVeby4rPYHqaW21ZBamNANqHGGNBDpt3BNOf5ssnf5+iXs9Qh
c8O+G7PAQFCkruJeYhSgiBryH9nyAvtvYJ+wNSpOeWlH6sTK5VhimUUcVLg2cC+MceIA6nR4MUoD
pnNjSxY7ItygghI/HRg4BVYET2aGWsw1gMo3t5ekJ7rEskHkhzFqE57fY2M9GyntMFMFazDIdT3c
iDhuzNnT8ZV1HJrdbRMNE9k6jNgf9SMJaAvvB+hT+VLb6lwJrCY2FUu+3Sk0++Ul+HHzwjqjL/w5
WocLjarEoT52AoffiRea8dX8Cw1baZ7WCMVl1a21f6LRARjECGerq8yYNstumN7+PfqaLu8WzcPq
3DLS2h4OFQZl8oID2sg+BGyGGYSoUAAdh1bcP8AoE91ljrjBlIHWqnbb+7G01fM91rQX7tWksC72
T6syttbuqoVWF4tBlPdLYYp0rExP3h6x+eliIgDwWS3sB4psvwljQWi8JqF0gkhjTAqy7odex/ND
r0S28f1pvvu5SS2zhg1jL/FdjsfHrHiLKOV4lMedQcnvnnMcXdrRU8Bnsn3uQCsH6Hrm+KHbzdYi
RImf5y7tEMsonBDkBZ7Ye15jT8+ZAEBgRyFKFbuqPMIw7jzVd5Xzq5nQnKD4TKbzwkLv59OeBXAI
MpIlAal5P1SbHkoOWUZh5Kn5g1+Tc1TWpBtMRO3TWjOEq4tiEYbealyM/N0OlxRz2t4NXMc+O6T/
bMLeR1HTyOsaPh+owiWi3AJWRGXKepcndMdw1Nxd20dJ5+WthqAhicJj7vWYoWqGF9GuAYqAdoTm
Fk+QWqfWkI1GS4UNhWc5mP4jk/kmH/+nmL6LPwcFIiC6id8yu0P+ixBpuW5I/jO07CkIZPZguY97
Ycvg4dAEd+fIJNs1TShlfp1IdMKj9ZjdmpVMgnk72KL74Cz8mlfXnx4t05SMNzC6abhByhCaBvSd
nb3Ru60LjZ81QxdthseZqS6GdHTWnjHZxJlcbiuiRNUAsQuhDPLsaaQZHy2PIFb4knpQSV9chHc8
/ztIhDia83I+4Y9cUhCz2MDsWDHrpNx0uH21nUm7DzH9cRqcaUMcLIGgojkPn30avrszMH1jmP37
hk8DmiVMu824eXJsZUgCLNJb2F7jaFSt0SCPREyaxX4Z68NdsDzCUTfurLURUsvY5E1AqZVVig7Y
WQXfo4zzPwctgzFl8Rl6FGygQxUCRdNQRCPVf5elzahrNJS2x0fKVxEeqIDrocVIt/O4GkdcVn04
St99ixK+dNYlvj4KuIaTNYDh7Tf7n2M+/PWHDjmYvNLKsvoKo+/LVBdgvTOZVJLZdm52UtcQbvCH
klkCTyyqZsbdNgti6R8/l0r+kBz1ZDNHdu9dxp6p6QL/CD4kyLHHnVLBxJ+h3yDtlr4vL9MzmBcE
vrRqKP3ngoL9DZ98/8L8s3u1RzsqyOXnGiM5UNYygpmD1N45RlD0N8tYLH1pYKA08dTkZRAoebs+
VDUXRAji0lbbg6VSyLL6uGVvtKyuSE62DQL2prF46KFk6cvz8TWG4m4GdbbpnE3riwey10t9erMg
h+nzCOW0ABQeHuUwDVF1i8EwPPE5nb4GbFmNehT9zQrMYYq3iGUEW6uDdMLdWOMYH+3tD4oYK7aZ
rEUb/AEqbGrqDRnkWyW+ZyJpZWNloZxHGsCzTPtCpSe6cjEeu4+WX1bdd9NtyWF9gS0dqL0OzfLG
EoOcKjoU7fLjzIue1ycoAkkkTn+rsnsfly/FdDT3nKyaL/orb9F6wTQY4tKA5Yl9X21rgE3v8M7k
oBi9TBLuH7xaur0TwfCRjSGsWzwgydEUx3MOzLcCcCRNPIHxy7r4Qxoeg9lKJX0UyGAy6y/uGxod
vPm40fDZp0pt8VAluMMHEyVksWkujRCA88EXo82zTyut+MJCcCejXffSR3KpQnZ0e1k2HJLdOGdn
uTyvVM2giJZrt8GlYE6xVpjMNl95qHbt4f0H4DcIXU2i6tIsesPCFhvPJghby2/KlxqhJWoxFtLm
sigchUFRDpyawmME94jqizi3Vv8nqqZASWXdUSgVeGSD9IPRLnbCRbaXwbQsLkXulBLRqv4JTSeM
uD7nqN39fPpPKxtKVYYKfD0CWUOXtqUUJh530ZPsLiyapmICz1WA4ikOx5LzYGrfpz7New6pyRUU
Q0WA24uisuj3LU9B559+rTwpudPWSMqnSlo1scOabi1Sm9yOFdTRjhsmE95FEQqzIIRxPknQ5kHg
iQeJBm++zUeyZ5o8bfzJZGuqFNpCOGAsjAaqjVLQ/9WurqLPV523Cde6G1OyJ+/elqyfArVU+3LW
BTLcFn9aOn2ycb+FVMpFEZPKolJg3zr1aQiGp/C2++jEw2xKzBHq+P44xEiTPdXB6ZUu00jvvGnn
4AMcUYyJpkpObJ3KqxKoMZrskVyWr6VNh5VIHbVYIKXOr/KAuiimjw7Dtw8UK7GgmVX9H7pp+huI
0M+UjNLYosCfVVlS4rR628P4xxRhOGmwFW/0XuFgqlQE4/o5JTiAIT8RZtLh3Sm1Qjqo/lRMq6AV
7v+QHKeakLTXqnxn2V0lSzuY4pQjidTQ3AHSPmNHZ6XKlnDC/mbfXlUVS210mnhlpUlEA58TSdJw
eWL8QmBhfWhrGZnvYFcpAtpaiznKm/TCwu6vWNgh9UIHcXzIiXN6YkbjkPkgDDSKkze9Y2mJ3wJe
cu0WHXIRSHB7/GPp3YfErtxL6N05P0ioVwZJkd4OzusVYvAAdRYjoFmi8df15HkCx97oGMFbHagq
RuR4dn2WmrwODK6Y/XSxnHReT04ee6VR/5bfmOlVXjLoXKX0RTDYZVn13SqUUkCK4B9TrF7YB/Gx
BfgTkspWuIoeJrRzb2hqvj+EG9VLHzbYesnjSxzSFO270WJH9OetmRrC89AgsKtMMrZyn5wHX5sh
uiJJvScFQ1yFS2wdZ9VHFyxhAq0F2AP00aOL/fjZuR3B85NP5zl+ALvInzYGaqKZNjG5inNvh9CG
XRoNYW+WsCLL8QJrx3CMZh8BbG/8+a5B8rltk2EEtadWI96ejaarQ/xukBmmJCEdKzk2aeaKB0ju
LPUipfnunsMdteY9tXhe8OSAYiUy+ObM2/Cd+T0yYbMIJpKZODyICH3C9anCbGvIZdUhi+aDPwG7
q335vG9EvMOfTDG0xFH611HhGEQL4KpL99kX7F0F/Cc5PU3bMRXoMpsh59MirePx9B4c9WKJhQfk
WWGJhsG3/NH+ZFAvk0IDwPxUW+rbV4deXXmNQh/8a94obmeC3uufmyySOwgjihkSw0P4p9pUoV4J
DhHPmKUsDGw2fohd9QSj0OcUfesfuSTGOLvqvbc/MWmRX/QTbqLahgrmpWV1CPc8k6WqISqPUNk5
gZTGTmAohYO77XcAjK7A3aBAKl/MTqPMBtlol5Qo2WvoGrGIEokXYoLyzdp3EJYRyVUBx+fVsH7R
3yu+/N/6CvCUtKdykpD/lu40y60+x4rGk4l4JFZ2q/H+3Co9HIXpCT9jtZowI1Nzm+LjvzahmIDf
TeDspYCrjZIYDVjOQiidioxjBt+eUkCo1lgAefOGvQZ3PcIxMX3tDqUifYTsdq6cyXoneVztG3fO
GvHMaOGU4RZrrCLW7ceRZqG5odhqk6vWg8dM12oCaVTCVtSTZvG26yZtdtiCvE6UDpjaviCNOaYg
EzDhwcJxMEcRomJtQyy2q4EQjyJwvktREcmLSJCL4tYvSevTJwmr5ONDcK6QgloI+SRplumDoBU9
nvw19aU5i7enlsE9MkwYKTLIc1AFkOckH8/JHApNDmjwck2JEWdQbT1OQy5zxkeaE4iL6y6s+lMm
ayoxI2AOzJwhyEOQPpKdoSjIa7AEC4BzMqqz81ujOId93sRRCXXKeb8LNaWv8xmB2RjUW6VLJQsD
EQrcuoetq4LQwNdALBLgBkFVHRu0gYObTTXMkVgTOCabMdUeUJybthchfuvzVpehMx3k5wkr7bs4
hWkC6duksXbB3YH+64K+PfmSj3Hkw3ieA/h2y0gEm6gyq/pWTR+wKWHqwpsD+Hj+BDjBTkheC1/f
1GxLLAlFhSOvyUKYEwQa9IxYsPiZ9NreJF7z/ki+57avedSog8LnII4fSlPc9bNobL48wBUg9LLv
9vjM9SwsMTcOfFp9sBTkN+bsEMHcBE6Gyh9iuPOmK559d88f9N3h8KMEHh0dp8/qLvy0Ctt5lzQC
ZeM1gqjJYM9mRA9MloNd4vHmBkSs5ZX2COBDQqFBlv095LDQ6phyGLZ1wKkrf52O1r5PgI3yDjeT
0cnltO/GFb0fDzU0UU6944U/BeWSk4z9FV3VGjVVU7OlvhZzXTYGoTjAl1HfkktqtHmEd1XqVbTT
cg6u6p7NAs/iJ0U9eTK/8LROPYzmETS5DZ5ZWhnGF90vKM1V9+NfSnzfG7DZF9sg5QIU/2VIyYPa
CWjc5AZaCcepy4gMAcL60yu8QJYvg7bZMbAyf5nA2nJqsgKjDlhJ8Hj2MT2xiep/zrJFA2Yg21a8
dGejiIjGqIVuCdrDPx4VBqTMc/ALw6o/1y3ty9Yy0vcBN4+8lK7CJ15BAdwB3bYBVnRhI68wmobO
+73gpsO3Ahrn//eQzQgrVdNi3tOPxLByv5HUDjZqWd0/Pa40x0yDG/coP5iZMmY+Byw7CDmabaCn
BLgZkGXlVzChlcJkP4/xSM9mNLWYafyfcIk7RCDtgrIzYPoLnT9rDBlNsP9EDXZQrxnDXjvlIwLb
chmbTfvU27MfBOdUXmKPQsyH00JwvfBO9UeTKBprmXpNXqzJH/enUyLJ91jl/I5vvKRbgGjAPUCH
VEJyp/p+ZtQHBGVTnCIuPI1JmXUVayCgKEoiXpJ7MP9uiN8nLUxcxXJ1GEIlem0UTq/zeicm9Gjn
cs+ojeYbMqUvE4tSrnnQo4NqVeR9W9UmavaDpZmvEVV3S7kikB3Ci7QsFj7Pm/Bk8x54l/IJP/0D
gacFPqkfQt8eLsPSBEUnw392lSAqfYwsEiMypq8Yj9L4nkxHPMx4szG7mQARgveszb8MkAC6pjeh
pkOIg9lJ/kLmY58/yE6mIuXtKTXwBgm6ygeysnbzoNeBVFz+JFy3wOye6pn4QpcggxwcP0YrqegV
zJnMslAZNg1BNmvSDU3ObIoIYYDEfKTBSFHWqduLlcPMbNHqaEQp/r/nGYKqcXdyNswtVSVj7xwA
W4pCWKZnZxBeMSHASunLYqRq8Wfv3Jl+Ryzkt9IxTfx6ujWJ45vq8c63elfRFJvemlW6rJYimpr+
A6ji3eLp2esURT0dMtk2oaNS5sNeto/Fi3kS22Ra/vf56T4JgABtAdKeLGiaMOWwQck1gbrFVos9
G9JQoMmcewkAfufouy1Wq4XbDcYgc8x0QTqBDsbAfpVdQ0U/ZJCJY5c0HI7ZMNiRvOVoRxmmthvK
BQkQJcIhdp9ry5rz5jKpVR1vnKuccAXGZkAmp3hH0l/SDjShzwgeqCovBaC/b0qmunyws81t7N6D
Jx/bSVIyiOTN4hu5Jd7C+dnQAyor+4YRqweMvf/Lje9LRIzBWRxOiT/wgnBHLbXkGzJFy7u/V4WN
xAA0ABqH67Z+X5uNuYXry7GP5/n5mtcQLlOcP2ppJosW1kB5X/xsyoEp5rxCJ0MqS9tN9g1Aj0id
Pm0VwEAJxPlkN/tR6u+kuxqanULcrcRlGEUJbKOeTr6vbnz8SHTPeumIQCVNh+SsGs/IxUjuZLl5
0+XbyR+xvlCc2ALJR8efCSKmArZYAsssvjm+cRxTQZpc/PhnuRQ8XsuSOHAIcuZ+Xv9pKcwzw0UP
IACXtWKWN+9wlZZgPslPm4OTxf7VlUF/8CiR4e371uFcsuYv66hnLaxFP7NnFGIFbj5SU9n2VF+N
w9wlOhK0rXwggUs+tSTfoIydG1aOImFHftiTqNljeA9QwXpBKmk+JNLBNQ7sGY7oPycWJVbCJK1a
Dzl20PMZquONTAJF9Fmja8Jl9nXa0d1IhOffJxuDbGwzOdyobeDmXyccyC1tyFkmZfGIjB6JPhFO
/KCbSk19g9rKw1rLIqGm5FdN8KfZSsTrYWM8WFcY2kOaDza+ZJ7NV/TrAEseShczc4VDX+Vikm4x
qQI0EHkPol6f9QkiihFT6TaMCYOwaEz6VZp7XWOrnDJhK+lzbuNByHIH5kj5YjmaEp6b609L8nb+
zjgR5Zomy1NBsc3BOiZiQzOW93WvYU2rv4J8u3EenCLOL+iGPzTnghQLA0L8b4rTnjW5DTaQBQt/
1IVWs3E70Z//NcqdExd+UOA6DyMeRImbtNr2viyr6Ir9ZTvXf5BqkM+nJLHtZk2fYgRYq66eGC0c
5mOzhZdRS5QuFkarXjRMGC8KHnlFAGgtBo/TGA69BuBsW+0pNGO6C9lUUj90xvOSWhFmC5p8yYIQ
UncJsurLdkFFkJlGLWQ0tTbbH8tRxpi95nx+wTcQv8r45ywXfen/9/loDUfc9OT08XBeYx7z7kFh
U2g0KRBdX8ENnR84w8013plKOF0LMFpkiQHCv9qiA9W0m3U6AY0MrUyS+5swealXTQc5CinSXZ/b
TsaWkblsGcuHMdjH3J2RVn6389BFwBlifIUU47YLIznyzDss29vXgq2Os1MWo6osSGL9rvY8WeeM
/RhDzgyphIPj8iXZ3TtfTp4sGLzEbyUC2cnixDmiEd/d67yZ9cglBCWaKgDUTp1lZj2IJZbjVpLY
2YYKk1ZF863mmIy8cvRuua7TCDZ53ALr6nJsmkvLr0ggqSFXapGBHIzPfzHKD4n8IIsl8W9BZ6Bl
KO5Mmcpo8ICxoJ2vgmnSXj0H8TU7YpyxGe3gCtJJORZ+w4ocwew3KQFu2xXPULJE42nuS8GQSTG5
G8V6uKG4c8GOlg6T5ImKt4kLAR0QWV0U+f1DYKJsWqhSteKd4U+lQj0xWuC90i8YfSGuMwAl+5PH
HYsgwQxHcK2TbNJg4cQdB09VYwodd9E3gkfUGgTGWRefsB2uEKI28/vHEP7GnjQDn8/Vz9V+FhyN
/YemWdcBklf9uiDCVVaeTtKNFFrViW1G0jy5YAvffg+f8B5h4X/VG78oqSHFKLrcUzwlA1uwC9pM
/tJS4veRFXDqyh2GrkKzOcAFmV0TWT+YnY8Soc026p9c7zjQb3U4gi85q5rBiIhJHUbvq5KHmCfg
z8xTG7CUEiZD0ZhyVCstHKCGbYjwSvAavsZdYZNpwRcweobSRzt5Qpf6JVe7gK9ka9ItpP+Sdq6a
LlXBoLwoZMx8ZuMUxERIYLvlMbOBlHpzyek2gaxoUpeJmXBpAutuBE8kZu3qeKv7OfYJJAwsQLn/
eWhshdZWhTjpHkTzvyjQFCjlt2VxrvBN28tjI1Kx/9rVTaaC7lIB0uoOUW6I3wtEPrrOTVm8rhr8
m67FJo+GTsOcaX3MtNOmS/dNySpaCOu3uAWXtm1y8DMmez8lK/UegVu8DMsJ2KFsEsIQf0EAIkRW
839A0bAvgadyaK3b65KVPVF6tWIEJXcJStPYHPuiFspKTuM3azmTcgRFevbETlDTbb9VVpoMuA2B
ITBV9ok9n8ZpzMxe+Rx/2dJAPncpKhME96dRCwrgNeXo2eyDNaGy0V04RzfCbEPziho4ffzea5pJ
nWVA5aq9A7A6UyRJ/vawooH12buv/wFJECdRlYJFOeOAa8KAcm5HebU510GsM7kTWrajH2YtFN+/
TOaA7qR47C2hAdL8CioR9X/dxvqQ5iUj3H2Z8+m/TQlv43M40folqXHZyoJl7M/FiNQNCOkVc1kM
hjb9mcB2QgbB4t3EJMEteOBliTQu7Y5mLiPhtN7GSS1bwMyv3iJOQLbqvosnDA4AN9VUPvvPGdCY
yhaO8dzXdV3BEVAyrn0mf0c67kwM8q/RZq4WClsVKSLB1HnAg6SNyjKm3/BcHOjR13l+toNDXkHh
hQAMWbwXXlNFNb9KhSznGuRqaj5smJ+fIpYVj1u1TBFK2rG5wfagUjub1EPxXfOxRdGcaA4r9WDs
KDc0JuF/l9cwIfAABGvEmQ9uhtJqXpK8ZSJy18SzTTIo6CiDiSVP5Wq0IPon4lSCQSqAqXDUa2Ei
/jMybs6caYBq67PKqlGf4BtRuYM2WPMLiXadxZVvSNOK45YJuSY1QSgO3DIFRsd8g+5p+JVf9GWK
e6n30aZrIsYXK/UKs8jT8FXgRoI7S/bJc1lMBWOjBiz5ixIgXfxtdNuGBqzNb5jW9jBcW2Bv5Hc1
4F0wrRnDIP/MpAaDtjVo+rTtXbVJOoaljPJ+H/lObIlhcGVhkcDx3XVCc1+vZQWQh6lokSjAhkY/
MuCHNqsi4Npxo2mEdxPqfu+dYAiS3KN4WavNgk/FRuiKKnFe0uhBHQKRh34kNuEBwKPLKD/ogyiN
ZlwzNDcevn4CuuQ2+oc5Brz4RvRfspLVbGcPgGRttGpEBY8eBB8evlZlCM8LUsOQu12YWFxQ4Yxu
Xi+/AJHjBDyvthpsWJ+yNPcSBrZWiXvQVcoWRDIvbI4GDuPfQYetiPKfptJ6HyN8lZFbYMKLxHzg
T0muz87rWkWQjR+hafkxiQRLc1QEx+MAvasyvZLFrk3ChgwuY04w2GTJPIKYUG6cmohTE990H7EB
nmZkRR17/v4ls57T+Y09fSYzZcZGVVimct7pOhhXfbBQfowperZug/8XrqsBtSK8ZiPQ+KroYk8b
c9VSl2qGQBWQeH0rM5P08arkK/nIdiLhAPWElAEvMOqaRDcXnO7BPe9d6wcLXDvJNG+UdI6WuFEq
k3X/tS4yqjVkmevwAhKNcwR3jNprvUfXfilRbwW1SmOCh4jG2OA4+fGVXqaSMHB0o/InSEYk0dM8
WgMlPUNGDv+5jv1kUDxroQaO1bsRwmw5UDyL9+VVKDeZXIcSdcz6pD7GF7e8Z08UemDUlUdmNke6
Kbj+kSTkU+4fJtLayZQz968u6bzk3y2S4+bHepTaEIQY/xVMV3ZenZNgriA6BrGyQolM3SiKMrdh
GPReJB6sS/SFauMPS/LHP+25rPAEZVYoxmLyKJBjYrr79kujhtHAXLeHoZcm49hBii+A/3UXWq3a
zqBzrUfaK19/CrP4ehLpvu8wdRePL03DDcpUwiAN2DBKuUSL+WefpQ5o7U2ZIn5MuW9vW9pktLOG
diARc65EgaIb392bgKnlagOu9K12/uEgN1KwvDdQb5xVRx275T1jr8mj3t5irzW80LTgzUNrjxHF
l0MK/Q4OM7aIzH86pTbuDzbLnVAa9PFKeXn2cnqf7Um+C4tIE92lzWkrtN818QLHGHfOfT4acym8
SJFLs/G3r0cwiD1/nEarSoxR22uPfPo/EUwCdnjRgLJa+wN9vS4KaO3hI9EqD1bXR8Ioeumvk+oI
QnV43Tycul52GabBocOL8sQftCMOHDdZAfzAQHULVuEHzchJq24KIHo0vuFL757va/wfRyfkwfxT
bFFWdwceVCrHcMi6cOrTLX9nB/JXtUV556fZnMdeMb5dtjY5jGnD0d85lsxKtU4NbTODlUONhn1s
tKfHP+vhs9BaguX94P/L+vmgtgy/zntfoeKXETRdc6EeYse3YOpBoc2o3Di8rLd3RAP1YGsbwq6O
agInNwmf4eyBGGA=
`protect end_protected
