-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
9EVjwMOgRc/9jfeH/eFDt3Zre8tBBs/3/G7EgKWQ0EkQHZ93Kz4tyLNURcdDOPfa
xmcCmViYlDRvTzoIYBTHgmo3Rb4cljIK3tqWxduYFp47tUzQQN9ZB5rK6gkgEm2B
UhUb6PyuG4d3V7BB0cYzFnXgef3TkuIK9Msp+v6rjWVxu/GRlLOu5w==
--pragma protect end_key_block
--pragma protect digest_block
jDBMr33YafvaLRry86u4twj2sTU=
--pragma protect end_digest_block
--pragma protect data_block
NMeFZyCBRl0otHlwAFGuvh5bJkTjm3ESrIf3OHgTWBm5YzskNE9xad97qZZnexfe
b44dVkiSQoHf4p4jZ4LT7jmnQOL/1isV/usa29EKshGiJPNpKhz5hFnW0HdpTijO
kk5miM97Q9OIzaTpVzoFg4FeBdFY9Xw5ujjfbgiqvmHOrTrwEHTdzf3k6qyeSCm8
Xd9T1Eq/TWNw9YgaqutE4rXkNPpzxNh3yw6y9jqj9WJ+SwHiFe2455xyOS9g+fdf
Gd/FTye/I8/tu9igYgudee5pe+lKXfHygQKr4v671lA5D43i7XWBnEsrbJ/CSEHA
JhROXGHJYl/TY9R6mOjOso9w5RCzebYZbnxwizur9mtR7hp5/jB77g7gEaqiCzJZ
PMTw4SG7DJ5I3kJjljmf4H8s9eZO1MMlQ6KU8rAqaljLRZqhzt7aO5z9ObVSTgSe
2vJz62Dhu2468ylZMpvHP6mDwCV40tt9SPMn2pIyuFBFPM0eh6xUehzupMEngpiq
76Q/tjG7OsJS1WiAoJgI1rhMRIrY8h8KljEhFciiym8QJCEw6LO+eOTkz6asrpf7
sDEyvCNC6JETInDWJQvOf539YJVZiNgXwhZYXyb0kl6IsR+4rTNX0yd4gBTPI4h5
0cbZCSXcVyTljm9+jfHZ7h0bf+1zO9lOWnnTDis8UwsV42MuVj9dRSF3wzitgoUl
scT0pXkRWcJ1o8AZNfvytXxlcD/YTHw+Twdj1I//2GgmR1Ber+3x3qdF5a0BJAX4
hlm9zzQTAPcNShxBSfQTkNqZmizlm7iZqE4gFnaaMZNQ2SWS+rzbXVRI1UUlt5jg
lBGQ63CX7Pu84M5K7ZXxeDDlRZWsfpKT2SHSW89g7mEYJ+mXsz1yQZZ1+WdMulc3
QPwzqfYYSUD6qiNQHRMxErqi7LsEQ433NTSiIZy4xGNjlwbvrSC6EWT0Kr0mhz/s
XvdoVic7EzI+IuqBurIOB0/90vpDwVlNyvDo2xgJ8Nx4Ar9DsFaGP/AwWPJztWCd
ju+vZfm456G+8aZPVBLMi7wIGS8t4U9Tm7OSAjdphklqNONGTwyMF7R30Gx83Lhr
qu2fOJ7Ri1gF+NGARBPXelysnzO+Tdh1sCLqBHfidN+ElkoJl9LA7mBjji7XMISx
220DVjhRW88Syq7AZMgvGls/hLym07MvUV8pUniP0JRZTifKPwpIktHJkyWfFWs7
tJRdYxETZy2oykH51L39Wc0iCGBZ3gG1FRanSJr5gvqhZMUVos1PGyOEHS9U86DB
ZMYKr1/j0E+p7ea/zY1GjAR7OKJBZILznmkMrDjUYDIR9QI7GgTvMprH7Cf6RIIk
fsFMNZeGiUcVls802AT+kJ5aN3slvWEo3+SyvaOQ4/W7155XYq0aoaaTRIc5KAUd
HYOPXwY94a6hkPBgUaCZj4ut2vika6fM0VHR8hV3u++nUjCc4ADCHm/EHJ94JgUh
gJgbpQALvyHApNDiKZuiuMyZMQae57286Ai0hodFpK7l5zbTKEubh47vZICV0DtY
DB88icX+na55XcdjkaFOLNUXyUsvmu/OEQEmPpR/+0FlYufeheKn88jWesmCTqut
Z9rOAVzyzgjFdSC9Md4bWL+O23q92xLpa1WkkgLSLNEUq3FjBg+Liq/SH1zsUrn0
nO3D9InhVmSPQSXRkOEUoVJ+BsuC/SANl00zcYOspzNYz4CEof4mrp53fCP+v9a+
nPSNVbO7fHTJxqhlybiwIYd9tIeoD43TYJG1mWkEXylZdB9aNpo0RNHp0eSUczAJ
ZXoS8ChO5OK5/mx/nmthxpFF9/3SLzMP1x5WR/degbQDktbiVffYekUzvSi3n4gh
+9S48pMJ4r2807RKubSeMKC2VJ+Qqy8lH4DyRhIlt1vY41TXF6BQwg7wE6GPy5+Q
LT/An0ci5eNB3PtHBxnlOvKCTOywwQtDz9Up7Q7B4s4mPwf2OAjZrIw+ovptCeGj
me2r/kLTSZ1k9s7BRCddVCtV4ZYJ4AtYLlbwP0ENtoOgPuqgAPkMyfsLapc/5jKv
1Aj4m1YmQiIXks4TUXc82ISDJEcO4fBSPXc4X4BxRlHlSXHWVJ5zCajJtW/lcIlt
TRnuifyCSokmSaF4+CEusSycfd2R5ACUwfDzTOeHerxrEIoLiNUTZS3ULl6uVgxK
Eegy/0nc0YXieCiVCJX9ydVnnKOiuVh72E0ly8LhTyhlNIjC7h49SlhO607VaNz6
psIZtXOx/04JnxgZhFvrSci/aHiPnt+G9Xc7gi51GV3M2sWJTEKk9Avi2uXb42Cg
Zt+Y7u50wjhc++YoqvkSI6WcCgkYZO/I2VlZ9i82YzWRggORRtMULWPvT98hf8Ye
JrxYGVCVdGXz4MtqekR0flwMclCHyH1166kGi+Kf0VsAj31U799/9LeXhnpq/R1j
SlWDE46piyMkyepeXQDn+j/BvP1qTfOyUkEMlzU+TrQm5bM4Fnak4b42a2e/vOCn
hiFEpzmVQ6Fhw1rxDWHxbrpVXOQTU0V73qR8AbBUsBN0EWGZn+tqTEiZHXNERx+t
tFIIcqOJueo/8wnqUnJ0KTHep8fG/WwcHiaWHiqnxkcGbj19PtuA0LLP/dDN5Cz9
vQfp9cb1JwWYEq62ardeCjPih3oHrRJm73oBfxrz2Nqq4eBS3nm8K5qHcD7IQ8W3
Jv1JDpd2vZ6ryYwu1KSD07KvY5uNPb3Qh/BCgVLcpYb+wEG4rRimxjQlmMKFMlbb
1d/K6dhU9bqXiaAvOqVLtNY1zfcjamtYCDRXC86SuC68KufaJdkC63DFB+S/3Qn5
zzXpEodKvtOtB4KjGer97J2l2ZnxFPksuetZVCcwedgsIjpAN4YAdmhFB4AAloKI
0ONqX7U6YF+P57pWjt7UoPDumhcECq/ZFEXMWjXPwO2BRnbH2KcRZ8X/x8M/kL4y
6bTphCYxpsq98P7tsvqBMpM8KFHM5KAeMidwSb8aLIoEntFA0x66jWxAlIE0oAq0
X70DxEuOIbzG7hgGEnNU8Gtiz7xZDC0iP/OSVex8ZRzI+cIZ/IC7Cjvt85JLzGNW
peuXFc29nnZacuzKNBK3ZXTnsEIoKcqZXe0Qk4h8ZHsYBo20aI7fhbeQe27B1sx6
Z6m9DpV/cNjgN1HPETIWqbsXxyNfGzsEbiejPD9kwRA7VGULoM1xF82p2BwZI1ZT
oZnE1Q+PPEKowABmMYLPRshk0mhgrVlDD1zcbDN6mtXmCRzn19enIUqusVmU/+JI
1wAJUqHTk6G8TqZqTTBh22stYustPJnplVySELiBypvFeE6i6y7JcuNLYWZlLGBV
avnYwDmNHZ++PCkTZEUEvcSUw2hlPSl4YzKbSrYI+OHLnpNVgWcvWo4QvnQb/VBq
OeePjyx1AoG5KZRHw1+uW5vNJfhZtBksGRuEOwhYEkHeOPo9Je9/LIUL3vKd3WY1
8JoMUxrE7XsBtKOAwoFCLvf+CWACCdMoYgDZ1YVD5IqKjhAbCQT0Eqj1ZHM+zWlB
+sRIMzw56HlrxThVhB8AUIGrF1cK9+gavibKcEImhNKEc/iUW/hRpS2GTgmJvZYc
4MypEpDFCMj2rD6aVmBKxRTfxz5maHjsvUUeV4/nGEatPc5PdlvqlTps8x98DMZl
gQpcRF01SDGkwkNgqxFefQcJAbfET0P0YDST42JPuwcyNdnysvL3GIGnclUod9gy
w3EEUflqgyVn7fSJmWrrglhZpLX5mMOhBeZTL4MmoNxNV0yyIj3KeMaWRWTPAMfc
YUxp/QLAWFFvcWGGwM/y7D8UBqmbic1mYqP4WXuCWkTqFKpd5wgGfOOx/Hep69Gv
zK+qJUnpUs19P3bz3eAqdnFwbZA6eaTFdFoEaoZTAkZNK6SfV/fW9hRLTHpQ2AnE
39UNizWF2iTVLHdENsUy9/r6sR5I5+5Uy5uWAOG1OWlXUjhXmPKKuPd6dNZVA/XA
X2xs2FAvVIPDwOpyR6+KKXG4nJsuJOLgBFk/CeyTq2BvU7+Cpbkg9ggFd34rEa6v
H2P5M+DQsPJfKg2HUMw4a+s7IPLAtQh7BJkwRGLlFyx4utjESJTnkMsa1opYncAn
91XRhCv5C2eP9mBm7BtmNiYCsrEVaa+6uhMw7hhjsFJWerFlhuuJEAZjBJKaZwG4
oOLq9E8RMJiwQlYTUfzxRvPUxhou1zjUEJOAIOX1b0+j4J6Ih1MWAGmGcNNBQX9B
sB8+WwCTID62XAMThrHlv0noTuNFyFtVpS+Bu05rAZ6rVhgnB2XDVBDCC+iovKGK
4FS6Khw5KPHJEyLWxWXVUmUfut6NuDazmKUegv2vF33YicwShi8r2rsDW1JQDZQn
XQW3rELYM5aGtbcUiUr5g1fTTMHA6nPmqEHrXB2XZsDN3e5k70ChwpP7k/o30Mt5
fWMNn8bP9Qa/nlgkfa5SQlQGk0+rPQnVRrK+JjY+hl/IGt6VJR/dKoUY7ds/9mWA
H5d5dvrsXAuuZrbwjrRvWZ1CB3f2CidYqSux0v2Ck5PVEmWOkUq5daXr00hl/O2z
5jA3fnGLlre/ZsqX3Sp+miUzEYDTsWl0Xuiy0m48V3ln7uMrjfKrSt7gQbtKTgkf
pnxOQJp+ZlJ+0+/9+V2RiLnZ01msE2lnnO4fZi49K7Jh8BUBP9b8N7yk4VoJ4o7K
CHIBrZii0EKPdhaLuNCPjHqfu62lPtNCwfSxJ7RtiA7fS4BP7INA7Cn1sML9vrIk
exGHwhHcnHlvYb8WwT0/sfgBrmH9IvmXLadqmN+8EcwDY/IrXOciFTKAKLEYsuOB
zpqWtVO9GQ8NVTD/ELP3OmJ9Uf3R+XGlyfXtInJWWfDBfSVSj9OYpEWQUPLFUpfh
RxA/iOR68FGcAtKKwP4XUkalOkwMbcBrWQk00iPjRMmjFwYbpRv4tnma304TspSd
XjvEzuh4U0gwhhZHBswDpFIKypT2XeWnkmJJZOvRhpcQYZIpb7+NqevQThjxhF27
yMM9DjiEPy/dVFY+WqSVLlFCAzMLa66LSY/I2xgJnXq+hQQNbfDQawyjroAftftw
fIMmBKtRe/Ioy0xuxhFYel74Ivx4nabZzgylFPO4vVNdvXa0M4s1qcGOLcB6O/R1
mGYWtdA/PQoR91ujhD8luRiwx+Dkjp4OoceQ5oRebVg1n5ZOUoS0SxHFdXb4ihIh
JVgb987yC56rFJUvawqrTiOkESrHnh/osvdJYdN3uhJTXxR3xD4fBQUaACj2bSlQ
T212dmWIqBIyjo+x0MJ8ILNjV5HpE6+XZ05cxKUfNDlh5KnThEcbQ/uyu5bsDHN9
oW/594L38ivPgYnUs1kAyh66JeOCWpGJ2T9fM4BsEWiEbDmdtzOvpyrc2scMAmco
UUTCkbqxjreXYGzDvcdd6WenCGOitM1yUj0O0qh2R7tz0PyGJCSnAwCbcRKqD60f
aAcfLI/AZly9+v82OzrGfT2kg0Pwm+dLhD1Nbav425RayhL8QPYsGgS8czQ5nhEs
fntVuvBbKIxpkgwkH4H56JOTeJwbp3tZ+Q2BnD5gfbMxVfQAgdPC0bI7SYB3zLQI
syZqaj3Qb6zRQRMH9FAZDgJNQcJxDH4rt5ZNHNKTyEpqaQmoLel9xJJbS7K823kk
zZEgdD4bdDxEJSY3AOmFQqsHTahZOkTgBpOI2BiJjUKGbjECMG6zfkY52e0v0K8P
/1pqgen3BgWlQeSmnOH3SO0iS4MGYlK2EftDPlfFlcduTn7ANosbkEUUNX9ymzxi
spzf3M86SL4aklhWz7S5YW2BQfpuaPqlaR8TMUWxdfdBoPzdTghW1+OPwvhBacNv
t5wR7J9xoaRmm92fNOmsc2NJ90hpnmtpqFaev4Tk/UJhIImdtxHxr9kGfeiCZm73
Eti45NxF+OgSuXN64aYw/XCBP5K2FYlIJ5fcY+ZZgI4AlibZexHMxJTi6q4fA6JO
SyBh2x+oxS4ihtBoilwp/M+2JQgeri2+mIsYDp8+6ztUsk3/KOTez0QlYsVcIE+C
8aG0rgpt8A38xvYgXGi3HI952PQOfmb36be4aiFc8vBQK0A19II58ilccLDGMu0b
h1esyoy/X9WNYjUe1SGTcgFUfelRVfPU/Vwj9vbp1FxSW+0+Gxh/gHjWdbCiYIKo
gXcqhlMQ1bzoj4/Ofq597GckMG9T+/ThC7E8pQRrkZIpmC2ukNr/TEla3H69VaY+
0bfx8Ubz3uMJvDPIJwqfX0nL9AgTJ+5nhc8LfVGLWgwsLNtJh5jalke7u+fY3YfV
FnJC4eFYZAInFAodfPNULbZ9GaY8Sh4mpTizSa81deCyEUj4hX7F6RxQfC18Q0Ha
ADLKr5x6liG2SlbST+TJ9msbMWFh3q3iSo1+s9evC+O4ZKiMApTXTW6xjwm7hi0a
qR5Env/Ac1xO1EfTFj36vnTiAcVMbNHqYb6DRum+r90a0D2kkdCkiT0y36HkNCT/
ndwgf9N5p/myv/1VBMESs0ZUT9PONze6aqedUoBNmd5FeEOfAZO77gXpaoZUublW
PGlPs5FfRcge5hiBaO484o7lfkLxguq2AVKU615LPpiuqr0toFOYFXyk3t5nO3Xz
v2gPQOoAebiuahZUYD5g66gTsCrgXSDn7IULlcKbQWRVJfsh51spevqOXeORznE+
Zx6LqxnKlchMREY/uuGk/7HIH6IIeth6CMqSZPHMuMV1Q2veQC/Pi6o8tiB9VfZ5
FEJqgAnZNVQ4McrrPRmbeuz/RuZR42UIXWQtPwBfy7eHCJ9SnVIt2RrAFs26I2U5
pBRxTuAi09T4BUigBcqxGNFrlN8R8G3NBPmsJPCf0eAaAOka3Y31cldIwTRjgOZ7
m/c/kSEAWgEWFzvqhL9/NpkmGlixsqsWKW4pwcFaRERTjgWEpoJt6UzIeZeprlG3
V4dO7b8JAjgDWRw+zhP9CRqlPWThzCFYvXioRfipS7JyWdexIzTQqPE2sEBXimtE
4aBX5F7CSdCeDfgyEwCdanmsirxnm8lCzCZZUq5XUM8Mm4fjv6HT1cMY2H1tFr7+
8k4nE+jqJgonKU+BJX2Yl5KLLCteYb8W6X5f2Bjq5HVhfjtZ/T30UxEd9Ji7tuc4
fK1m97LpofcrBUi1Z+d6095DAYRGWcyNkTsns3TlwNsodIgT9mPP+W4EzfALdbJV
cyVUQhG3HZsbp+jrqlZlnk+nJB97gh9POJkMS0TPzC83QEl4XXT8kA3ntQWulg7M
1eOUx+JNr+tGXTSMQcb0Z4lOyY/fbMJh+4NRWhL+4aeLdgaxWwosbbjAkdNJElBo
QTCmhQvXB+2fW5tBmSP/drQiKFiQJER6z2rDB3lkDgzqMqXxWKqiOJBgpIcy/sE9
xg/7In9D5rkWoaW4gY0ps2vC6pC6F3j978MBTIL9k7TZvW3nhAwJxvS+58dVp3cL
IKDe16v0/EjyYWdiLkjkjRA33AQKK9r64DnSt7y60VOfSE9CcOBl/SKuNu67GMMG
TNCltBlYHYJkC/Fi6mRPR4h3KLU77GLRwX27PKO1fjfhSisU+ya+TCjiyURDvGiS
JUVRDi4hWcb/1NH4u/7QRyk3Gik3Op47aPLNrGcDmg5ZvlXppMPFrg1La5pSdRTg
KEMCvVIoK4vBw+bMEIuGmI6jVid3SFVXsmnTzomQwvPjkJrETuogJoYHi5o2UJN+
g3Y6bC7xWs1EhHTjF+Rlsr/GQxEpz4d2uXTwGcLPg7N1mq4isWBMZ3qD2QSyqDiZ
HQJNQxnjxBNKhfXM1S4H64235d9Q4V6vQiLa1ax+j02imuoH+IH99+uRl0InBmYX
ynzViTC/y6IBOWoNfxn7bM2J9OwHCVgZSuk8spOLvBAXcPX0Q1gXFbRIrQGUEU9z
SFgnckyax0JGkknts6iAvZe1KRDsep7phN+pPJx+/KM/ALIk9cmD/KcjVhuWEFSq
ZQVf6Sjd/KN24Njm8DTiTS739+DvasAgMoyK+LOiu/XooUOAtB+hTvEM/AD4XQcR
8l8l+ZYkRHDZ/lotMNiSMhEvyBPLdQdwIZFzvmN3J22EK+QnNx3Lj2/0PE93GSSU
ROQQLs9GhVJI2q7UizpbBJuNdNvkXoFKb9wcN2+uaMupMN0SrQCMuhprNdx75VJ0
4tAS/CBMFrjc7/fE8FLsyNhkgpLUImAaris6P+9Ym8ZZ1EdUeO5hCMCgPzir/hUc
+aqC2sHV8QLwwXNVFRh87zrfQNeTgXpin5ws+wvJyrjk0l3bCuDrYcXu2Ogs5K0X
O04Qg7gBroNP38i3r2Ii+zzFj84TrBJp+80lc39BIP01vmd2JHQb9LOchWLPB8DF
o5r3gB/sSbGW4TBA5EI5g2X5D9ji5pEjvZhWIU176GQuOQEH6f4chzOB3bh6zNBy
WCl77vppiPBcln1RZMwMlAjNno29DWHPp9uEVWoy0zWVTEh1JLiEwOTvaBaGxPyh
+muGxtmH4oOEPCQwMq9IzhPhx5+5VtRWxAAptuIBHYlhCnzDAsINPn73OSYfqPC+
Gh0NqvKQyvsSLJFL4L79HZIRwXCs954qTI+58NKKsrcw1QOPO4lO4dWSYPovwJFc
Pm/HDLylpWoAjwqkpFw3gR+RZyL/bpHnXOchLj1m+5Qu9+WwDn8Y9PTnadG1sNB1
rRVhNrzO6kxBKtFrV9JeqXJULPQnV0nrdwYr4TUDbYb4WJhqaeNr+FXglBMgk8kE
UlduCEQtgG6qnxcWz/0oxbBDyG/cGWu+RSk+7cSA1Btvtw1hXNc86ws93uj8mEqr
es1AedA1zojqvTbqWhsJLNxjHQwwoXvU7hMa4nWjk75ZFPPWP26H/bWNQiwZ3bIH
Z+mvSz/F3g369FjqhKD/9MG+jVHhO+ELGW5vNnygjyH/ReQLWXpqwOasdQFVFHgd
Sxi7JMEOJU+BNP/h1wEIAJvb0Nf1DuKWnKU0GKBPxMmlB+vCandA5Le+krb3yXc4
jbI/zmrd+oqx5dK1zNAsSweTpVoFiF1lxjSuXCvRENnD5S6xlf4l/qmu6FzMTvtQ
dtEM9fi/LZijQasudlAHPybJYFWd0c0DihHvPEnhavyEtfQbup3ADuf4OKOTK6aN
OqDK/j2x/gL0GmQ84hyza2X1gcw78gO0VN5HhHJ/SYc305Qx1uKQpzlMpw/jlxAJ
Fdj9Y3IQKzua7WPDPIiG9e7vb5xxGeuaxftZ4SIIkv2S3OTs6uS+lvGJoe6iDQG7
FOwqNMm98ufqFVFri0eWQXIAVUhuS6YwmBHYvLeXpofLl91/Jbv78ndcGMvenX/2
eAds3D7p7SCJhDKutU57dddiXg6e7Ftk7y4aiFUnxt6yfinVN3UOujOshfBAVRov
lKT9mc4PEWAOooRwvy+6dT1MzHt5J+u9RAVGYQSWzhP9ENpTZJAiYDM6j+ki0hNW
Gi09Ut4TgRHvMxeukFeQl4Zut0WrF+wnm2zFXTjfqfUl7+8w2oDtGGwDBn9Z3wlq
iqsXpG/vYY7vmKPUCJRdRNqzg8vE9Xk8SeZvIqW07lAiB7LhW426aXjLigY/tDGD
pKuJi4wyOZ6uEKimJqJ/yV5Bba2LwGnb4ctVLnLj7IaAjUVm6eY4CvMFzSUg99eT
p+KXYAmbZpU297ISqIx6RFtnv58f+XGmJeguSDuK3Ec20UlomqzJIgGX8n0hThKM
dfAD3e6U34SHgznd4sVqVGQFgknCVYsw3Xyk0MQBlzL2HMFvrwzpQc+C1vZ0FPG8
xPvn6qurU3Fs3COporwvGQ+mx1xtMg1RM68YZ5I0vCUNc7+buDac/tIEdO6fsqHH
p+nmmcvjHygcfVjEZ+x74HreWefpwr/OszWbT9zoSMFBsKy76Qw/75B67zBapXUZ
AUkPjDD9z0zjVNQHqtV3S8DmNKDLnMP7INVOHot7kIQZArKGGSskFMZ4xKMjUvet
hJCLu7Udj5Y/2zbLPx5ThnH9Ac6GIDwfpn9ajeXIjzfIeoGyOkBliY9MYxRCrw43
hWosNFlmZYqQFwCjS+EKPdLfar/CiUnjqikyVw7VLLDOgs2mUa6+kp5FjeSnls4X
2KZ075jBM08GsYQiS3WuO37F0Lksj3mfwrrgWITp85Na5xwObNahrt/X2UZgI2DL
U95FdDM467q7iPmcCDJdHC19P8d3iXW7mfvN+rkFbh6BlfghZnEo0itO6KRwbZyk
q+UtS0JEoBxUAA53EGqgHazOxhtSqIznOWaTuwujiZK8uunEqRV3FWINWjtV8wML
yHXHsNBuzRoLOeDuPvR2WTqHhaaUhBHdXWf7GysUHfPLULC0p1NYlu48jpzZd8CM
E46k95BvIRS9fJc/LJIocpbyH03UhPmIZcEQFUyXEilZaDEi3X8GKcV4wTHN9qBg

--pragma protect end_data_block
--pragma protect digest_block
BYdLtgHQYU9uvSXY6dhZus3qR4g=
--pragma protect end_digest_block
--pragma protect end_protected
