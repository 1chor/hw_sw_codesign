-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
VYvyHplEySw9EXBTYmZFwe4wKAf6/KgEq12HU0gMSAHdiVOXwVMZIp8+S7DV7CLE
cYKlDyLvpKZi8/WINsfyYbd3827Z2GWX4Ow7V1WX1wdX9svpYsckJOkyJOu4Lzeb
DKNyA0i913HwpYrIgUlHsfe40dIbRON1Th5nib/AAfU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 26360)

`protect DATA_BLOCK
lV7LyUb5PxI2m7K3Ygq0rfdVBHdrFqecWgxW2Q+DP7ZGWxLz7Rmlf9m4ek08gt87
VuwbF1pETSTH/sx7j13Yhb4WNjWHtPmPsaExgnUFVsEvdtE3vvMpYq+JgpLrRe2m
7gP0ZIBrpYYhh0Hyg3lOxdM3jLS7YONWyc5QipRMxJXfcGW7U0sBoeeB3ifObOvm
YewOmWhOrHAQb3FIAJqp8s9B2fZZB7Ru9AHZxhyLApyzVbH4NJCqggZGLo5L1yzB
iWwTjaSk/4lXuDtS+uZbwBBil7hWQgKLePDIhVb6vUcsNk9O2pP4AXUGnCrM1ntS
Aqv/9iS1QhV26i+HmLz6datwohQ7oKC55hGMtAAuxwD1mTpldwfQceI2wt4pnSMG
1iFCAKdfpJLqbuwYMCxNR6+HoQHEzaVEVOxs1unjqKBL4aoz/W8QrNBbxmmBMYh/
dyH++J7reB8Tr9dXPevPA+AIuQ8gGc7nmwHtD8G1uLH3wiyO3x4g6PLMJHfHilnk
aMbWXxTY4Y+gZ+smKErGKJSbcVCi0Nb5j+4qEVNvCRAHIPcKC08aQo+PrchFJ0rb
P6OrBfQ64nWkDm1zeinkFnLsBlP1lRlOCrR5gY6OzKT91iy7gYzAVZ5rSF3E7WrL
D2lKxT+m3LsyEiaZwx7p/OqVesFrOZcIR+ftrp7SQhuTGbWzHZk+I75OAVwyC7bx
HwqDWfxbfmdxr26eXcGSaGcLTDEoRdiTt4zzL2hiBpDCidPBn8pNsYlTR6DuKDls
Zv0vvVcPJGl/bjyDMU01E8fcZZpD7V4bOeoPwOFPp4DeOGp5dIfhYSX5yMCLpgGi
YJoNxOJo6HmJmliNtDbBFn5CTnPALkH0fJUEkCT7WdLo2RTNDMxCeU2xWxupXn8A
D1v4fizM5z5Ndb77gqfxBtuveFoinr5ddNDg0NUckPSxQThpUJk0FcWSyPlhRkjb
rrzJkAvbu+CX+g396qJclC9TQQ5URPi6GuTh7QXMvWZrurz/Oal0SnS5r7GOgWct
URP6UC5giEQS4Dv4Vk25Xf7sUApwHAyxx2tc3raor4IXyckXhzOdMCSKKai+pjiM
8cIoKa/b5BGqVMTaCO5JL5knb/s65hR3/2YN3bwDekQAF1uVkuK5615k3Eujmanx
qx5LzMbY7HH1s3wOhqW2SDHzDkokmWq1BC2O4cJLvg7+NWdUgnGcdmSA0WGjsVkf
oNiTjJNX6Ze/mVwcgAr+ahLoimrxCFUjvof5Gg8a16c1uwjWEfJ28IZ6aayPAmJV
gpFxYC7AyW1ONmwzQfhSOWc6UAjiWvLMtNB0Fy9tNNuDjhScFdjwyluzYXm0/iMP
cxl0eniW+oyE0s8AFRj6yxBUkq0uRcHfMIrHO+udtLuW1cECNbSUuRqgZ2JdQbZd
tZ6hv0yUyj861sV64IFcWQrKz1HMYS0MPOBxvI8RXwuLUYSRJ66hQTrmT8NTbpQK
zr37Pdrh1sgEqQ7hVE8a41EEz4heERT1Fub1IxcunTScMkT1DVzXUjI9rc/qh622
DaRgZaFqR2jQYRl2UOKMT67OZMx8QW8u4vuFMkaW9yagTMAthxeMJq49vuARBXIh
NVbxwUxsKdvbZusDS0ZpNXCK+QR+HtXWC3yvs6nye7reBYEax1Of/P0yrdkRjUW5
r6mOgXI1hI0D42B6yvI4TLPiRwrPwEUAcOqu4FrLRQXiczC/9RrSjROBZfzmNRrr
/PzO/XdOUv6fE86m2FeiMgIzMJst9H8zNaGfi4M7xKR9/4C2SqmUqtOrZt3aAyuE
spjo407n2atzTmgwDNS+z+SOFe6V24U48RP8KICE3ypdwzzBYWXR3gAI/TQhnPyB
4GYOjjAKD9wUPeT/c4gdvdmDYQbs1sX5pE3HjrZJ75lIw8yoOQ9ZT0wD2568PwNh
8eehKOpY7XqRpDnQCGG8barQKVQ+2go0CYXyQ6ek1EHOc5t1VD4Zapjyk50KDmbn
P2nGE3lD5aTnPb7VZw7OAYxrKFkefxZwNBTJ09FAlgIVV/pRyk/CBDvlzn6n9uFU
2EPtf6om65W3CZQghk40VTXwYl4MD5iUuodafxlfGrFSLvqJrvwN0vjf6nWjDwCd
loHu9gyRQYEjdK+UyjvawEg3XAMdExrElHJHf+E4Kfzt/mopn8ipY7jY357YAXVd
aF2LhKE4m1UxSCusWJNEMMLVyjH0jT8vHmHfk+eiD2r5VHk6oQTw1YRR+YhG1F7z
uC62IxTJp92OdnUQv6K2ji8HUN4kXNY64i7Fv4BWjZSMEJasqwSs1PZmBfyc9MAS
sS8+h3VwSrQF5IUtKelw2YseJF2MlN+vTId2NXsA//yWz2Xzmmx+NCK2O7XRvw9m
PNB6DO6I0YmV36jlJJeUnJzGvK8XfrRoWPffNrtFLfPQMi7sZgnjsusTEEOeq8Zt
CFfJiWLmrWa9Zab7l2yD8nem8u74Lu4d9HbI2s5ov61Htm9HSbBPuVJRHoAbJZWe
E/yG6NAAjXt/nB8Tjn1Cs/ImOPtFmAFbiDUOrzNvPf3x2E4ujKYWgqz48x7Ye8T6
AuPjLKsovRuPTXkHlKxRxDlXFcPUM8gggyMgvAB6iOL2E8HL7tjrxEXffHjNCh29
ufAerYkvzzQ7h0e7c1S4GVCHxsJFKSg16u/PBi7hNXo167qWrb1T98hGn33nOZWA
OWLFwoE6aN0Pw48vmQp1r0ZHK030mrCSdj99IZLYWCqtyB3NzJzCf+CQ9heM5t1w
AET3BreXa93cCj0TT12H7IfzDEl9BMDpS2WKyrN6oeVRvQnfEMhyR7f+rMB+d4qe
czlguguKsGdtZwStt1lIfuslwUHEtO72fen0CV40zfY/qVwtyRuRKXT1siVMpPvS
Eqh16t+EY4YsUFUL6EswN+DarQgvLTjwVCiaFEy6oIuDmaYyGZhJI5rVhxCSwFz/
KXvoOz2QrwjEM12QPq6Tes7Lddu37bcBjHXVUBTQGrpNRE7gNb0CMvRV8FddNHk+
e90gatPtQR66YCAxUvhOBVOIx5PsyhXoZ/P8EBtTx63rcNpZT9MpWhgtvbDTGLW+
XJ7dypBEbwdYPPztLWmEeccutTv9+4tI9487PdxPuSbM8RyIADVWCN8/94a4kJdI
JV+847ognfrEZotj1Zq4ULKs07sK3E6xBG/CacRDTIAwOLmvpCG+r+8kvuA7v/r/
tYPWs6wjyV0/ineOPyetYQTypfMwngpuB4orm7vOqN+t+mC80zrmM6wIwz85wWWf
B1BY5LRyMp52Y5Mwbbt8+LKrNP2XmiFbuwpPZ5ERKgoKot44QXppl0GLshrBRR3U
M5FbtEi9W5DSyXUHJYwkZCACkzOO6JO8UR7X4IGo0QSBOsHTnDOMO8FO2hnNXrJo
JCJxnfxD/29FO7JVLb/cEoq2bjOKBXqSnnEBdAVl/WkuLMEmBsH6o68by2McwIUv
+vitmrujIVwmk88GKJBZaE3AVmANRrb/Prp2a0ETvjk2UClC6ru/GRnU8IHJJnaW
4imre1zbVG3XKG2/utVyAk7K5CgiIc1FmjXF+LL0By03w+SrDnRaz/aRgLuB39sr
hc1hb01qnN3Nwl7iWcMBijugVTYoL5y1mdEZ6wY5cI9nYGrpW8teGdO2ZsYnSAoE
95fmWV/CTr8TaiZMDI01K7KK4l0YKlWezKhapV3MFpUzFqGefy6IcjyYMGMKtFrZ
LU6JWDlxE/GrsT/bhHKrfWHjaHwUYEM7R+AH4Fqj/FtjD7Pk+JgwX4edH7k8TOod
LXbzeYLlkljThceI/y/rS1U2KEX7SMMq1pPV/kZSEFF1acrnlh7FkwfUbpnJSdbU
fGm54uXa8CXxHQVBS16lrdAO+iCMwu8CjxtInNrmFBsmeTVwVI6QDht/cD2fgsJE
1fjVMm0bQsryPg1VMeBuHToqp7XawU0SinGxesVEyJ9s+AZDhvknX3HyA47C+4N+
cDCnlJCv3RuuBNDTT/8O2khj4aTP0D2u+U88lDRT//QZ/nn+YHCPpBrb+U7OghZM
SXqGszJOpjSnW9wnjOM5It1nrK9lQ5Wu0f0v0jRfbGR/3446zUnqYjHDDzJpiyl/
z900yLrVv+IqNO/nMav3AZxz2bEiGvlo4K0H4Sy5oYmdbjGqrJiso9JTiNYoz6Fk
bTCTcpSSNpeTWl8LQLQJUtqB7t3LdjoXB1GciNYjLeAeZPKSTGMAwXdx4I848ofq
1CQEFYT/G3sd1wDURD1recpPS0EK1ljNyPXHAPmP3SV2bHkJunRKHzz1fPyKpwO9
VOtcqsHkPMU4C8NUWbXC8nbRo3zhhd6sotCq0au6e0+TPqrscoQRfyjKUl0vMdmT
43mKzo4JL52JTT1DDGJosWtaHCZU7ph2KwrQCgucma9ItfYeDkYm54q1ATtEmv5V
/kww6KPzwfoiOoCwCjTt5tlwWVqUJjk+/C3sgUtvimZpzgWSGBsK6s+C2N/NioW/
4366afVw4a5HsUJZzgk6AqOvm0RWaMXmjES5EZNOfK3EwoU/7cHosmuXd5L1WGC8
ch4kXGB/qs6oSqsehWjdb8nFNYB3XpIGds/61ucOqAX59Fy3kvnjEWeRh9Nn90Cq
ccBiThvEuT6MFqLylaKIKGlQrh4Jr31H1zlpdqdLZT/vof6lZwzCsYI2tFFqx0Fe
PfJYp74P5TzE26ObM3hCZc861iiwFaht72L8TytSuK8MaAbWPPJATxOW2mCEw+4c
qKXDY5PQnSeNz8RcpGvzZ5usnjKL4UqcvMnXvtt3/kY0yXyxhoh3ghetHau4bxxf
oPSqwpVcbAQ5loQo0yNcc/jc+vaaszpumE4kaFa1sGRQD+aPSVZNs4wjsJUy/vuV
g3dk57iiHIUu9qt2Q191hvHOt/9VYXzcrjsvF1+hQR4YBlZW+R07ijmpw0xkFu6l
yBFv0AIcCsnAAffTbhWViAhPNBGFO6G4hvc5Dw0UrzB3euIlXM4H7LEMRRmdZw2Y
NY6BchF6ViHuF1QzJ+ogYy12YKe8NmUjDQJnJYea/Y1GFhHGmipDGcGt8Hxh10DH
0HMAcCs9U0iw5C33RYr8xjyV6et+/3Jnn7zp/9bPnQwFWDkU9kNRrTJyNQ884CnN
VvPrLGTXo+78zAS1ESEMZrTOvH1Wc/Sah0xFBcAcrs7nTA62JcRNoB7a0tC17k7s
E5NuIih7BFGFdY2oMFygxlkrLhLAZBPUWOA4d6dRxh2TCqbw9HHkm5RIPw+rQBdg
SDu39qcZWCQ6Erdli0cFeQVETM/K4JjV+YRv/DBbi0+ix+xN+GwOw+tAWw4GWy37
l533nA/63HhPRakki5jDRpcAKBxQqWuHn7JOF2V7xcC1agrSOBZJLW6PltfbL2Vl
+mhCYPj3ZFtjQ27+ffQ7nhS584SHD64+nizav3LCdvZm0/hH+NGCm07V+iAuV7vd
IxEb79IEvaX5yWQfJ1ja5DPhibY47/XOtLgpwgfN7vvwS1kbJAshs8PfMN068r0Z
GnZVq+eM2G+TgH8pN3OjaE7iv4kYyEGLnyhWgO+QiMMdye8CmsiSq1iLQ5NnJNDi
zgSqFlW/uaaq9UcIAaSJCMgKdBUkmNKmSCBzGkzXFMj6JY6hYFZrXVGvublDwhX8
CTtzrM8nt2sIitX9mjgXBeC6siwcSkmg03EO7ntVU9gti5yiAU2au2MEnQ2ZL9Pu
KvmVglmPmJYu0jd3oTZ7z+uhws1p1GrU1Hbg2jvRhazJjVruTZ+2esz/xk9CK54F
i4g7sh5E6wqpaa0+oqrWQBeiLc+cQ/XL0QzYUXh4qgvxII6DvcOv9FK028orAiZm
CgXKi9R126SMyz6iC4Ckzl7gdN8VHZpGKwgMXAwZ1ThKH/A2d4kezNfqu5WNZDPB
jx3sLmBR874vsF/PDYVI910z+trDtRAcYoKvoWtQrCH3j0VoZ6o0+LvqoAiNVVM5
lkpYjt8x17Df2Rf+dgVg3Lne16lB7I19YjulgW3bBvykKDy7QkKyD23LYmLp2oza
WFUXd5utUy3HfjfWs6pkqMJmSGFZ+csgK+XIxSaV+spjGiBgaGe3mwm8m8sNxCXY
zCDCCkKnQ4gPXevxUcxEyB0Xdu0btVoXafcXQ9gsS4PureM5C54nn+tf8XuBBAyq
oEJwaycKa+hYsQRQCf5WKRbN/3br/e7/qFyfNopgoe9DMlDLWldC4KT8OOJHjJ6h
o3xyR9PZJ0rkMeYjWCr8z+JWaRvx3t4kIJJ36dfl880GZTvdPYp8BfmDnTVgrvEd
R03A8xXLtJre7fjKv1DXjKxbDg9hwKQ4ArzPSR+IQqb7OrwZGyHGBQiT7Hqw9Q8u
oiAiX8nuzc62R8SBJIlgw/SaP06qhbjOggehGzPjFcPKufCiTae/pnJ6Y/e6QzWv
AGAXYJwEbOQguwgyIWxbP9U8AovfG1FHgZUxgOrl3spoU/27sN3Kv2LCOspAB0ml
gtx2WV51nBFuv6fsdyglpW53Oh+TvgF97Jn5csfPrHMePj+vxpNI5iIJmbLcz1wk
e1gBIfSyvfKxwulzs6QwP1hn6dhtiCikoeounfjFRrNuxUTWVoC83LSeb9C/a7Eo
V7NFbn28PcGq19EZZdJcQpG4xct82yN8MuQrQA0MpcmX2sWKtt0Vjh95ajDMXD5z
WJtouS4VmwnimCj9vXR2rO1tjhg1Px0yJVLM6r4+AiUnTykp4yi2EwELxoErQo/H
/Y5zVdU7Zc8sIvOY8zuKji7eo9pg3+H6RJX5HgQcXdJzs9/5SYFxaFvj3EWgeUDk
NoQ+/JgXCI7sApG0a+2TJxRafVkJnNkBTWpIK+bKU/aIPBpq6HJ2yuxQOhPae4t4
+1wt/cd1WR1lyXUrZZ7roAKK6efFdbd3kMPSf895G87JsS0ha0ztfutw4p29yXgi
FJDLG+XLlMXdY8xTuMxvT3XodQisvW0in8KRREeOsPtVzMEY4WNZm0WAU7Y5X9gc
8Xx7aPLUXC2zcAXnQ3b5EeBI9R7gM9VAt/fkdMKHqk9WK6DkSlypx0ay7yPFUPFR
I9yiOViiACuWsIe3gQAAR/GObVhIIgg3meWKv4siIpAPTccwGuORzlrNgsPApLZj
XdCrfzoBOUd0h7FOOUfyB83z2++1bo5sSlC/8Vs9PXx9MF9APMVpdisoA1GXZoSv
r5Vmz2hjky40gFsJtnAQ7n/nCcyXS3ab48bcniBv0oFg1wHRKsTEAB52L2q3BOFX
36kB0nfoLvxaD8K58YArYkwbnHH2/GaxbNDo6z+AK3SKpo+CqsCJj4oXZyGv5fBo
p6W8PEv+5cQwXm68HfQx0I0cj58fygWNfvW9I9eC86NbrzGNX4HQg4dj8ymHGFzj
lMHKfOfxcOVoPWQvdtEwCrxMBwsT5087plFjO8rMvFvD4Y2feSYdL6IFwxXTmZ2u
aP89/H6E3mlnt7kfdzaWlFg7fIYL+Pu/OWtWWuZ3EryRG9u8CQ3vf3OWB1r3USik
r+5WwkAYu19MqPEokMke4tV1KHeOss2QlwuW1uFTC36Rqy+yZYQ36zhvX3oardT1
p2fW87xaJlLrdZt9iNiAzfHEuQ+1GM5ljfYbywoJGlctmGm7JqvVDR94iDh8X1op
teYx2NbY1Jd7gXVv9h50fZkJLtjS37G8pFzDUijYKiJSMbJmEDKsGpdKeXxsCB8w
V3LOyNvKEphFOfkVsfJWAwnlnWvkkpK7sMdjSKucGrraVsGT4cPhdQxCGetmT2Vb
zrC0ljuZPYQkuLvr4rPdMXNoll6HVbDevbxMw/Ug6ZXzZuswsBckQHoyA8hzkNzA
SgOi+c3b9u09cq+eaS7GM4D3EzYJ0CEUnlJAeqaYQ5YW20vuymTP7s0DAI6li95L
upZ0s6ezSpjOVHoNe85bFkrZk8xVdsJpyp/ULxNr7CHEUZsWBtkwOFkV0I9mFP7a
i3PWgwuWgqXCJ6tu0ECnS6WlsxmkLlLpWo7CK8KuJvWG3ASTokzbcv013pzJsGEg
S5R2yK+JFwEpiPLxGQsUXb19r8cx5NO7cxqBf0uwcgBlcfEm9YFn6B/PuVcTDtNZ
VRZ6g+VG9X+b+XMOIRXHg6DjpUrcnRsMiU+kcnn9eSu7JPPN0omKnOhSyuR/Sgw5
kErWOXyo4bfqkCHhUaf2j2j6VHkNghFN7D2BrST1W7PyiG3ECom0pj3bf7vZH+ou
tID9SNavR0mrmRxukaJzHbs63ypPkoYd7C7DcFD4WJ+3NbM5fgPPJH4AZEp1moYG
H0NiEFukQ4JCeEsVdddMwTSIJtaT69PHJVeCM2rU7L67WeTUur4i4uuhhL8zdAts
HlCB7mPLPBeMGy1/wyWlTRjXk2ipogmv9/U0uVMVxEGixMVKRT3hRYPJcW4t5DH5
acTadc60hv3PH4waRJBYkdFiDYWFzAuCMBDSfIjkKIPjRlae6KYcvn6t3E7fVuWa
CbWfN8+lcFlUzrVbx+YhpmyPWwSIROYZrHBFuv3C4devZkIMBh/KjfJbzoQaTK9Q
SPAIM4w1b00CoANNAjRZGEbfjCp7uSxYKtYb1b5aKzlthMOvBaxT6lowYOZwBCeN
oV1C4+zpPX8bp/oPdeVIr4f1YX+4bwX4gSJk6D74TdR7eGFU8TsmL+Arpxl3ecKs
NoHUmJW8TSiOth9mazc55hm//tJuEdQ7uZ8ltTqn+uP5AXl1VdigaRknnQBCMFHA
umnKcHUyl/EBkWsNXhe2gs2ROC7i8Tj3kSDHMbx02QmNdG/ZFuAnUdd9fjGV1Qlp
kbVxVbXokXlKVL1eu0E/ibaToXqFU5R9LxaKIHJPnaTGNFLc0Go8aMMwYB4fwOFD
CAQtCmvSCjc3sP4l/R0l2K1h7ZE9ej81XBMCffR/3WLiRhwc2XzNzxit7ZBDheFS
a0n29ul8no6tH7VkvhahbG0zkwysJWf26rqk7QqzqXOX0JPtyIkjR47sRabXXEKk
jC3wxNazhNPM9/vPnPcSyrES8XRZioNNLgD+I81rQTbimUVx0ucjYlnpp3JNfBre
8mnNRc+RHnGtrHGE512k+io9f0kRHOx7SWHBEMZNvigwGY42SQGVioh8Xr18I1sr
JWdrFE2oBB+QosT2SGQUTKdsorddhQfFhoMShr8ALtfaPmiNdpxpLvXb+1Q/sXz1
/qzy+VbzUlDpQyGFlK6S0W9e/xdjZ7BiVkQXKzjaADSjUK8rud9GBfUp5nTbXGCJ
i3Z8y8Kx8VkYeN6s96YT/OXs7CiSKh4zNfkXkbhvpNS5z1fNT6tipGINbXfFQtG4
AVqTdkCpELbGophl3wF5D7SdwZMV2sQvf6enILKTKUbZVmFuJNkv8LXuHvAXRdBc
0JHBStAQJBOfNaxJipMhr/Pk3O/2MReemSXIor4czkTUo8WCNbvib2UpDPPIC7qB
o1TNNwTocKQg+EeMZDohgSV5tY2t8MeJuYFm9Ud2DXft0D3Y9cWLnbrAW4oQKO0U
Sa44V7CqMC+dK4R4oBw6Mke5kcB+atCVknGmuB+UAVff4oXMR7/j+vzdtEWpvwO+
2eaVuJ3Ew7/tsVKQak45Jp9EvoF3Ayzy1H7OIf9sNTqq04+g2rD1qnyFNob/qUwP
UINw4vkkaDoLA4RMArDi6Zcfoxi1yAOd5m6K6R3HZ+Sx2DfvdojB9TH1xw0knTof
YR++4FnCLZ1xKTlS9JA8aya+eUJSMPlNs7cB12ZS5vCbQCr5STCu1HSl0HUoH+IE
LIQHnVWOrkr2bYY6VeAz9mZ6bVHU53VbN+KmNbLyXJo6hb8PMZClVUXpdsQXveZP
+rTZFkjSbH/4BmZYzT8aBVvn625RMD69doA+vpMYxsxxRdH/v20ithgDho5SvVMC
LzF/ritIUYWNZtgjIQI67+zrCrAa+Unh85t0ONaS1mADK5FwjENs5toNcAeMq3z3
aqU6ftSnpaJ/5OIibspS4n/hT6qR3jXrLxM5kjZaZ+rImJ3nMmZ1s1N00UO3SKCI
D7AICuziu++Px+gsvp12XvP2ULwmmuSad2UnorFap0go0Izd/9SRMtlphpqtiQiL
ZC9Pgp42DO1tuI16fTZ9fWrOqKqXIv7hg/kCp6OnUJFkiYxPGaPC5c62FnEzF8I/
aSWBSDXwGju8KtKmY950NoyPXC5QnQNsPLkq75zn7EdhoGCZ+W57MjFZijatJzty
fuBsma33naOVUk/1d2LaFtc1OKRlGYuVVtq3WMjB2PVtVrUY0bbHyYEDaAegc0AR
DNs0l/4lfe6nm/m0VZxL0EI0fgmGdSDbgC7TmVN6iCDIvjK/TfQBuvMBaz/tEWUO
UBmeGF0w0TyL/OkOIA4gPDYT804TQAFmw9df/0CYYCDkzdRMv8DQV8rmfhexcNmA
A/r3o8Y4m+Ewx9h3hHqJkirGroEz28lc4AGArarOwBZIHGiJKfdkxCfvC8K6YRSX
wB8NiwX8PAJhYfm1xYyJPIx3DYPTk/BIrWFtT1vSL1qi23VHY0A6MwpA6F63+oKS
spksNkAD5aDWZ8OmW3aw+8dC3uU/vyJ1UoAvEmQVsWfcpVHVL7UVoA3X7zaqHm9e
K6IMRFcm/NJJ58l37AKp/csAT6p5XTr+F4RRaHUD9UtSJsqvGwaUBGtcyCBFM3pO
HCAyK3r99Z8gNkagmf7BEDw/8UYmYCmJvAHRpCenWZniczlQDMbtET7qWbLamge9
s55dCpvDNnZVEsq8da0b2h00AepoRGDcgaFT+9ast4zMUyjJ6wG6n+HXOjanXljd
XUbzWrqvvQ/FFe2nQd+RhEPfRxV0lRc50xFMsazQXY4W393bTsy4u6ZZ3TAKCVGF
IFY+PTpqTeLFfedpRahd8RhO5jZ6quBRF9mt1hl3sQam0g1m60lgaufLDs9PH5fw
GllrChPaCp0+zfrfL15d2wBeDZSiPUya6f6Hq6k4ssax8TGM9fKWieoS3QF8Dbai
6jIPJYazHOjzokCChHPUDG9EWgWIOl7BKISaN2KezQe3C5iK//2akRirJzzaAfOT
oVxnbGP4CEg/E+nEqUTnU3yUKDM+qu4sNTfNBoQwlLgnJiRXMhXfCrjOA5ZIsuLj
IEDxJnkoONfbntcaxClymyhQ7QLppbLz/NtIHaMzToAnyRqGYXtNix79zi4J5b6n
5Ydox84oYjvSCU6t4UIXOt98/bJ+Mpfc+cf0i8w1AeoCnKwbZhRZzJbyNLoMcZGL
Rx8sGwntli89YW/qD1unPL5R+3Yr7eKp+l8BijoT65DIjILrBrwVi788bSkQq5P+
xsTwhPlEPo68j0EqkQLR4Ewm75WY/eDGne3vTw9n/qPvsrjhfngTOIxoafAOo+Kw
ULLrfOHZDCgdlv0vpnVXsrcvn0RgK6oL1Gucaelf9l7Z53UxBRFK4yrASk4w/DoQ
WPhIxdXLos5MICFPVUqtDa6I4L3FeaXrdLz961kdRfsWtLRGqxSO+bVz2/l7zy47
2ms+XdQaVnZG9xyo0ulwYkr6fKIPSft36FoyX6w2mnNjOIeejsz6UyOX4zw7B6A4
SuN8zTMrlsO+8TVxJPKkkgDu89wzvKCMTTS3Ocjlzr97YdJExZgGTELSI0GZj4W+
QI3UYZlHDwBe3ibsMDiGkZeqxota3nsZgE+sERWfCxDqGTYG3YlzOC2L0CaLH1ng
icOV02la6AA/g6VC7aW3jyf91sCApGhEgniNDZfhpJNumv8juyn4aY8dg8HnPqMc
0eCnkXRNgGJ+r/4bG+okVBsjhnwYYnM0q8yJ0X94OFaDXRzSEheGwchXU4wtGa/+
WsTfuaXXiDUXGftnXl0LdjMIUYFJHJs+iVowWS/8nu0Hv4XbauiGDYu6hbxglqyj
JaY8uPISNefbym6ZcvVXxmK/hbtGIjZywyR0NJKyXt1wEgGTuJG+lU7dBqOXjXLe
OB2NSw79BmtvyKH1t1sm1u63vPuiae+VF+cHf70B0OWj3R/4JUwQw3jgaDSDAkRa
poW8fP5iH72F/VT2LRP+XUk6BSEzzqR7tPPy6XUJRWCkwm/i2jTqnECqA0Wn7ueJ
cjLfUCyBaNmebQb5DIEK/RWf0R6eQOcvqFvLE/VKA6HT5vM8ykmj2cl/9yBFQGx6
RKoFI1nDs3numalKhFEfRBe75ryBRkx/Hg7xxu3K5mm8lqYenXqvoByDqalQUVdd
XqvhJOXu+csPsKge8rUvXejJDvtixvsjMsG6zSMpiL48/HR2FJTb2kwdOmbEPntx
O5IN2XhvdwcGVlnYuzibWi73M1S1A70lyfw0rPOzsCwzMmXjbfqKEeAnNr8God4v
nEIWxRgynwYkZh5fDM6DzFtoY02TMUjvuNZfIT2MsUfBHfugqJxuW+jcFCB7Uj9h
C3Mt2jlliHnDt0Y5P5KaC3utWGxIuQAzqtaZ2aX/YOQqR6XU42np6ouOTQWNovR+
Tx6iVe98j8gAef7zJJ79ZOYo5cNmyGtz76D0Mj3uiLUinRNtSK+xTSAnkvBSIIf5
pXMwkNgUK7skUAVn7v0ZmbFGaLtvtQEfQyr0eAbA4KGAtP1O7mvJ0kvUMQlDGsU8
EKYrwGxb2toQCFjID3KQa+1r/GwGz9Cg8u0g4lj0Ns0fNxZsOVplUPm7ekukMKSO
W/W+MPt0ElpMMUmABn4nhEsqxKrRHD7+4iLt0gj/IBJq545DOtY3zVPJO42FTBRJ
vBr7LLzIchjcSwwIBx5/whERx1LsqvzybmIQVlwwDQR4OON/yDa3QCnJYUwHGlhH
/uFeupOMEHgaUBLkxbBR3hAJulu7IlUf3FCgsPxucWmn5KTDfLFyPTmXbWQF4LDl
FL7v5oQEekNUuxiux/KQKafp3hxsdrjNgbI0dr8eAtYT5HKuIZJ/g37z6JMyogoY
UU5yyRD/ZjHqFIZJRcw3rsNIHpalFPrioeVUbVWUcc5k8hZvA78r03a0SKuRDuUO
oAAJrmunWHh9nt48odA/YVq+Ij/ZZvAbqQJMP16/sV/wHc9U10s2cCEXV/0eRqNt
ANkC6p5WRAquGqXV+pa4SPFKBSIZShn1oeIjiHDLSB4gJOLdp6IGdurTj52Ua4zd
bFMfqPhFcVz6fnjiCe4/2FqyG8259PR8Jx2ol1jNkmQVi+6d+fDaThgpHEue3PR6
2AXdCqU+dhcrPUOD44oN+srBf7gQfI5ghElU5mRV7U3mvuEVrSlFRFhFgSghnGrk
uglgcJyrkfcmYo+d0Alld8zAiGWMOr2C1Mna755iC6wARfOtv9Lpk1rxaMNHbor+
fpXpgXkLtVHIrWjEjDAHETEXns1iq1ezocJvPsWquFrpNggu7AepwE0ADgh9+2ey
QqlL9jjdoOyHahq0Lc3jJrefhR/S5MgJbseV/TzDGZOR3vq4AIMU7oiVTorTUcc3
+bfwoKfm+RmjU8ctWUuZcCzp6S1uhg+2/S/c70YvzjY8DPi9Ci9aAKJ7ovI3lC7v
IqeL5HF1DVTsVlegnxuSeS+tEmRhXkFCRfyMlgFgWzsCGLTZRVEWxiXY3zrqTteK
lUou6NCEPONTsxOPj2OekJ0pcdg8fupbEVxk/jTdHlNSKHmqCSmHrS5GRuhFxTZh
ysqMS+Bs7lh94O+fl+gvKiL82OCwcrcIH8gcoKuxYrxh/vH9Bg+m7p7JO+av/Ihy
zcPe4dPZcKM7iPACvQaw1sEcLOmFhpmTfl2o0nfJU3gZ4ZAWa73LQZJcdqoUPURf
kQRVaCpAnJJNt+GrypAc8jvSa3AdXNbph/rTgfD9id+lZRhhs9m57wCczTA+ORJW
ho/GKXRF7cipJO8No/h7TAYOn0U1T0De98BMfylaJNoEqYRHfZ5DbvQJZ5B7SjSS
IP8bXDP+Aixw/cRaD4fMhnBAPwY334+RMlVJIc42d2EJ0uvmzCvKqGD7zqHpF/rF
OjkcpKcVeJVoxKLwECfL2qPUVzG3NAdiwk+SjrxnS/Ki3wXNO9egH8p8pV+MRU2J
IFAcrWiG7t9M+QXcAFB1852uuqgXbPYXw35H5m5UriBhrpXECnj6kvijARiPjXDx
n9IGQ38S+RzwmJ5kachYN7YS7T3H+zWqk2TjOIrF4SBgMToE1UaakCqCpoKPw2/v
GR1gUCB483XaJOkqaIaHun2d8ybNhWJxON5DtNilrFGpHwS9MsG0k2DEEzRx8Eal
qiJG5Dkmc8RMzUF2JCe5sZH7ROlMqJ3lZAQeE7JHBvKC4hcTryePjY/Ga7Mgu50O
EionwKJCUpw1QWlrnKuewZ2Ioy3q+ZLThnBrmfESuJuWoO8FqJMLX2c5i1f1lgi3
hh7gZ5QZXYdD71hTZuNC7k27suCF57ZKJ2YgGK3u6F+wimJ8IqBD2Fzbw3XtKMZQ
A1lUV1M0WjLVTFnwXyryLRupqWKFZcKhO3U/pK8Pxvh2GN9xX8CKhZKVZgeQ8Hpr
HOi2MwYv98UCqoFTOnRVkjVg6MBkpfFBESLdcDMJbJqVxEBlXBO5UFlF4UD6mZ37
BLg13Ak2w1xmDBjpOqaO+g3YP3o8wJUzr1MdWgnG1qt/MEGZao2Wol1vfpmfd/uS
pUu5XfPnC8tyWp33LvIEtPxqDbzjTdiMOJvD6vnXWec2MCm9LSvEWMdWKRjtTX7w
l6i4R7qguPoWJmE5Li7taHXwgSrauQWrU/UWfKtkbzFnMgRfwJBGe7ZURaXbefli
0JT30PW4lAu/hyVbiXquuabvasflUB2HsK6yYqIDFmvUgiHLj3QjOowCg26KwviP
EoZH9IC5EymFYGnNHZ6gANrSASIhyfrekyF0PKNC/W/8stDRbz/NVcYK2j7PX9lg
pgws/REpQlRw5KLAFTjpgcKyhew27hV9RdBrDPBnk6Jg4BtLo/7ZrvfnbB0fCUHb
A1wn5RoSulW0Lzzq5PGQiI4N0lhDxMmC68LfjCcG5vD70Qa6EW3WIcEf3loCCplM
PHHb21H/bfKEcvLzNAYYDhWEJLdQi5FsDMlgiFYtR7S8Q8j+wxk+hmJtnX3A7NFR
NVDOFTijHyReGsiAMyVJX4NBQhfn2u+wXTKRopocfyYeWc8xZjJq8+bGf1vi7KbU
o4DKaI3htZ4nT/UoMD2l4FFo+X/ohyOMv09kuRR3HLbVq4RzeF5XS9UxBgjyP2GG
WGr78Ws0GSM4VyWc5JspkMIxdv9S5F79eXaRZZlAB4oFjoWBBbKFc1ZKX+BHfbYb
GMI/CIH0q5aPQSD6lXE5PT1SR3ipusZ/bgPslfGmJ8G6WywxBUJMla65rDKPC4Dw
mu0QzYl+WcP4Pvc9/OwRVKmuDnOy2jcm0aQlLULi6Iky0AhMBLgp5d2dU/WP+gnP
rt00QzMFDuHsS1kBoxvA3/x+ZpXOEx3yBeSywuj/T2OlJ3s56VhFkhujVGGay2Sl
5RfOg5fc7K1/c+KbqBRU26meULmkZZq3qlelAYd1mVdVaTye7uR1kLFUrnmM5ZZ2
95B2T3edRn0rvvsjBtq1YMf/N/3kz2q0QFxwkmkTm9ogX/m18YLklDnHRB9FxJPx
GWZ7r5exCsVJB8qqq3CEgEXF3tZzgEy07MC6Jm9hXVcA4dRV65AKHk+a+ogf882x
mKXG5//nG/Zi0WlSKcQerepRrcd5U+puJ2i8WrdyL8qWF6mSlbkeBGGCMdk7GxoJ
8AuY9OCFzzXRLlBUiHtI0Wy5RkG26DnjBVej5RjKB9ww6sJv3J/0Q1BTMAhParts
hEuJfuwVK/wnE/MecOO8BrzNlz7G0hBDfavFyE7foWKDCfAHwQzK44LhGCORk0O3
vl3AGPguZRWVN0fN9LaDd8FZ5YnlT4dXmIbLEhrnhThIBrMNFhdHM+Iz1AGjehrO
b5RPC3zGywGPDwfyK2igunPlmBzLQkfq5MAs3rz95pAxP4MFgJoXXZCR1d/8ZNoM
R9wHzf04/jGfRwdErD4+83I8hzyFiYfrES/sMnJd3QFQH3atLQ0dqGCurxQEdoM9
S5hp8FxEmkTrsNUUOSFrEnz7f4krNiuztfgwMT3DNShfdmfB6EsgY01N2Oq3fkiu
nxbU7RdHvqeR0WDvT844/1pungbiuVz6Gkj60wABmLXiR4AnLqAS7X84MxoG6PyU
mxoIBuQhN/0BCcf4IoSSS9Gn3Fs3P1z8gDJjtS0GkvMOgH7SSkYbKFtUXJthMwW8
H5ooX7Fi0EOkXw27tPhKeJhfIRHL4t6GXcdRNRkrBtYeGRLbVYPpkKDGEeUzf7YD
VvjuujAeNx6FS1WAOx866Q8PZ7kBy09xpSEvM91WebOVk52PbpZxf42wmNz4Ncur
B967cll6ooHQPbGIUntJ7Nl4ZuEhftqUV5LUEI0QbFqXzZ1sHpE8hLEeY9Zow+nu
SoMQOmC1cWAj4fkRZYdsuPATQT+BVse4yAe6v2zier3WpO+ZbVtIAc9xdQE06kPx
xRzGIdgwnMsV/GKzIuMbyVL3rf41Okqv5PjNceDSLoRhPJna2nPV0k50wdFMV5SB
F1afpNyUSPeK6fJ6Ixmjdz5rSV37zoEl+gFvNgu9/y4Vz0cWpf08BCMYhI/rkrGz
/dL9ZOeShVDfazdjGCO4SVI5Ldipo0yap5d/ETcdYt3yzj7M+K6tXbp1dDxR7z5f
OhehlQPo0Iffi8qvYIvEZ80jH5l+ZyVoyNpoIH+/KDs5TxClvArOvuSp6jeT1Hww
8Ft4GXvHDhJEobqhAouuPBc2xPWG3/cglCDYWz8vyz+sIvV32245HjGIDjdwafMf
BXsEDPIoA8+Irsj/AmwQfqYlpR1U2XCbH8o9by146jQC5VSlUmslmRQl5D9/1ZYi
e1aJNBDYHJ+piF3MuyvoXL03DVeyKqb/sGLpvEd5SK5GCF5sZkmZoLbJ1XhqKQAY
CIYZqf9DLnTagVLA3dvux7jC3/Yj2We3H4htElmmsTEhJpZPlIH80dzg4QZmox2W
HwqeINcr83mYzxtBRZJNyJGw978aBHEv1bA9z9xN6etTabLkIvtRueVXtNlyveVL
DJrvEjyUPYBMj20bbPKo5zhX7/4FAcax+7qfnrwvK3qefH7sYWgHQiTHqcWzog8O
dzNzK7FR4TW7AEFsgz0LLgP38vlx5DY6jzuU7tR9BsXTgN36nwNW4DQYWFvVDnlu
38rO3yWzrhY448fCAl50uighK4WXcCRTQKIhTLyuMmvtzou1XOxqpBDMP9iaV6jR
j2iSJkH4qXG+l4VGqfvPxb12xl5HMPjQKMOfzaAEKg1g496DMV3WNVss4NhEeGF8
l7Ow7vgFdZeGMCIrGuIK/d78jPuLPgW08ieUcxpMndkbWb9xIVFnHgubVmGYbC5g
6KpV9hzlIVhKpDcSTq24qahkGIpVQ1pIBkMelfNfOiM5tZJJGTH8GVbqfGjFOby7
ufuUYFPzl+aOri4mOygcALEPyHTN/MFZe9uFqzawjEcXfAvw0DcdTLRz6WhUyI4P
75r5KbFFTVG36JdqRZG7Mo3bA8aSxjl+QJVvKU/fvZJ1x1Uv3cPyN5MdfAA/B2LC
7f1GilRuK9PY4x/+Os50d49eM02+vrw965LHJPdwuqLUtlTCGhZJhBgKfRr8+CsE
Ua0Pvp90HiGC+pn3q44pCYIsToIHsnMiAlS6lCHLX4sDv7ScjMFRHLxqW5cJ+FyE
z4bvPdAYGAJ5lF637hJ6JDJgjmZbnIvgXeCscqh1jsJaBOv2oJxp9toWAgBG+y+1
DBxf7gA7J0jroPrFvMIkJvLhS2IQcMyYN0yfrFNfr07LshyogzVGv/HFY8tTxhZ0
LLutzlsYuzAaaH+RUzoK1df3FCL9TJ12x38hDBCFz7dAOCZCZ87jq/VQ775+Idsa
gmhn4r8DubNxGUDpDWJMSIXAdcynebwcRAU/DadNc7bJgeWhIQ4yMp9yZxhuPyud
yPrafsPXg3cIh2jxCg5gjwaDQj95hAc2eCdXlBbuOOTUV/Fdu3lTsA/LLzxvOnF9
6Mqv4DWCfvFO5RUW+vGtTXCLqXfvk2zPdprE96lvSvISaO+2SqTY7J4pCf/LbweD
lPLfAABtZD1WxcsimFIJdGadwosL/Zf5Z+xZbPABkJz2NyerQ6HpTzwYLEq45xU2
RE7TWVjqucoOhoPsKYxlMuPopOZkV7GiRfbZhSUlm6esw2sqymZ1fF1gWokCdiap
IDSd1YUVUhJxuQZoWCl/Z9lq4auivbJDH17IhR0iEYDnMyU7qbnkGXAO6dEYJSbi
i3+Bwa+OGvSuOt38EOfk7Vzup6xhCogwE2fkmfYiwGF97oP80hBeU2AVARv6MMOq
ttfU8CVuO9c0t61ekTER1kPqrYsrcykeyYo3wsuTBw/DLSNEAeOZeNRxe/MPTlG4
zAb+0X3npFERBvwVyJychlVcNsKZW/ZfOH1PvY9DA2LXDvT416P2TER06KWtf/qY
g6OezRXHLPJ3lJtslfNzG68DW25RZTRoI2huTylIO//cbZIxSJIvTv3BqhqitH1J
tzDW0qy6uSFvUOHwKExaPc1d7EaI5z+7Qa8QRhbaHV/J6i/WMI2WaI4Y96T1/+Zp
vtcqtxu/jxtbZaPd7hhK+tFN9zAFVTiRmt07Glu2I6MthVIB8bgHq4MjYnXALMSP
7lkjYyRDW3EtZJp+argQNcLSw5y5PflB1WTPHnyhEgVTlcGtgpqLesk7DXwPKcTV
JtQVhX4oFdsytDHmwYdXfGOT9j65O7fgU2UFY1vdM1Fn0FtLcc8t7N2Fze5b+Nlf
P6MWmYtGV8use1vCAdlbnTqt/6uB4/EefSlBC9cOvHjy76XouYoUvaUNy/dFppO1
oqbcpvJDpocEDXR7VR72ROOgyh3Q/xDfw9Kqvz+LPfraUyr3yqMPndkZc/q4WFn8
6a1EMvTuR+BO3NWo1KW1BZktPINCDAC16mAEyLkTQZAcKfbXQUQzCxuc33Nm+Pk7
GyibzEmG1oUhfIW5pNF4g1pykO+EGYBa6Aiu8GvjgPG2D707f7Cg8x/WEAcgZDmU
dQuUj7jmW2oPsEO9HZEUYVS+KjRlymlvtZ7hPAJyDLzi2AYW4foXXs+/b4Tl9pSS
2j0ka9XOdaM3cGf7o2Dk9NDrudWTWDv/RRGjjS/lubO+I2OtEYuHOA2VvRG8VfoM
iLTmf3fXm4KaC0Dn0VEbe8xjMfpJO2keJsocohsedJAKbWEfHe7WcxBENschtXQ5
5RR1Yg7H2cOTAyaVshdYZg/aAsoIauPM/5BAwXdqHQE9F7gUzZ7jndVIb7Dw/+ER
sbBBv9X+iUxStIO54GgURnchPfAooXTmi/I+dcOlDQHuPGWQLjrLRDncd66zOPbK
THwA3vixSQYT7XnrLPGE0uM9V2AM5Nrh1uOg8cnmVaQ0C33MQJlZIto/k+ZLcoDa
gsIyTQ0b3McKbdo9C9u2x4lx78JMOgqh+9REVvdj0Ns1FKOzeAeqXPFLycOIbRny
hlno7zldiKQBLdNx9Ok8Hf7whPBxG5S27MUv7NlQLNk3OsvPMjdAoAQkM4iOqqyv
jhzsiqSkKZmCD4xx6BIHi5CUCBEAV8KltpP8Sbk+MmXJPl902RmbhXnuTvAznvNj
RW0ZrA3VmuZADXi9uj9omUN1U3x3cUHrYqPPPXAHHgrLOIxkdK6EhNrH3N4qyhlv
0G6y7UEcwsMuUHnz3CGrnZR6brfOv0yoqCNWSJzAG8naIYf2lywfv2iXUExtxwEm
D9CZvMR5/0J5L7rrz18APZI/xQUDn/YRrpHQtUNxayCQl6fHiLt7ODWdxT4qUuXi
zll6drj5+AlX3cgFPaqCP/Dc8oCWavvJOs9xXN1iAXWn9aaBkgi2cnuhJJYbxoaI
Jx3LC4EWqINGbTOuCntsTJv+ycTLpDMEKdFfQFmsQ1UNdfQVcaL1hltrKO2xFZIz
fD5GbaGjuYDY6dcU1hNxMAtJdkNqwpyzIahE97opfsN0g11XHRlwDiJstDFpd/ba
vSLlftmiwJwLBTHpsAoBO4oqgd88xWN5zdMmNUDazzCaAMFf9g6TEjxyUZgDrdaU
b04NVJklbrwN2fBklqfzpTFkgiQTuBFtrMC5pvvwM34vY58FXIWh99XHOcCdGuc/
B7g83vUs836x/vy3fAvVn+dKv8Bu3AT0OkhQpJ37FFslXf/Bgz3yD27Z2K+kkk8b
QWl3OJyQdOYcKCwRsruY1K+z4C4Hy/7azsE293GHQ5TWo0SL44eSbLVRq4nuAQCf
a5Y0vgB6Jq+QsyCpIOeHlqchuvfGvyK87jFNEr5SOOtaFUts2V0rlIkC+8u7uliY
/F4kglmK/tIOtYLFRq1SfQGLG1RT9EQprdHBS9am7rwpyoyhZ4wuCkDTKeHSNVsb
Yx/ZZ+35cfvvGoT7QVF6l25K6L5iCjk5lA+xubBCKmfNDVFsVUtSUeMyTa/N9zot
aKKyrdbM0TdCM0xeGBW72RZ5R0g0C3j4+hdFAlH4Il9hcNBYZDxAlF69dNUnVCYi
L+1JYXeqWPyPTHSG5s6BYiv/yTtuWc1cqR7AtEyzDdSxweurEgC6O/GvYaCFilN/
YbSBnSKm2k7j3SeLyK7sXzfY8Sss1W8nlavRq2gnAr3dPpX/AM/lWshOuIMTqOsO
Y82+CmKEEsvzGdi7uVZqIzZeXWQUxUOpw2b5v6NvUtygGypYDKBI76t5hcTDz60D
nZe/pvr6lcb1LMyk2HupBx9uTxea3FWwXlCydgmXi8QpOrfWkMwkVNegQbyF76W6
JHYuloSDfeq4Nsb8LS6iPhH176O9vSd2J8qlqauWjp91vMZbezvYJrQ3pX+PBhQS
saOCpqLSf95wYWj6R0UgnX+qCk+JtN+0H94EaFifwLFIfgsSJtutVgBX6Wgu2Q57
ImEwx9Y7Kd1+LRfRjrT4DITEutqgTr9AlWY8Yv68jnoYJpaTK0bvtq8MtK9asHEt
0ynFEiyKee6Ja9qeQsg5+DBEyrxT+kK3Eekd69rUChWLCKgXBiY8A7Z6m8xJWSuO
FHLfDlQIZNADYKt89WfVzppP1X++WoKR4a6JPCosicfEQobtptx3InuVP0pyGVse
3kmgHYh8JkqRbd3Tdcb2VM8XA766mcKcrkHYzx7AnYnrlMKnRxpE8SWhHBMMfLKR
cbveaHHhOWUz0oHDB3XdXUwUSEMUTHOHGkfviyVnQWYt7fzZ6WQC5udUyLYZGK4v
sJvPV8GqRQxHNNvQdE2vDZwB3ABofTLdI5V19KTdILcTvggg+iOO4YEgIFS4sBGJ
srjOjsysHBEssmJHbSkpe0ARV42lbvbvGopfFKWP+5xwrbgVjxXT+n+GIyG92bbU
W+R9R6Uj607OOXjk8si6uJE1Zm1e0naFZWzF3AhUB99+aqScXLE9nDAWpE2odLXR
imVw5ddCAiu1WsSS4aY7XkuXS7LhuYF4tYdlus8z6hjmXvEQpUI9Ml+NaGnGO0ht
LDfGvX7ayqx/2asbQNCn4U6Ikt+mu6Pfwohzztk0zHALRSMFiEEau1vjKZw/sTVU
eZmGZkCEaGbZfps4PdzmZ86DfCgiLHAvZwMepl65s4KDnPpOcAGpxhRV+gbb7ZeJ
vGgbF3jwNLbYexDGQFm9OWsmWDISrfXoD6Qal/K6q/fCTAb/xTjkFgNFIsZVgWYl
NaoHsuDY+AYEHx+26cTz2dQyuaEz/prQOPgz41vw0TbYWg7o+2Q7H7r1Wpoxyl5X
Bs6/4UcjLkbJbNOHh0rHf+SUDLICIJIAQxWz6h0YVMU5mlt9AnyPJxAsLp+FZEg+
2rVRBYAtDQllwJxH4hX4rJcz7pgujdAMGcS3j0/5xns7N30to/Hr7IZHJ0asmu71
bmHHTjtqylwhy2U/j7scTWP9Q9k54AMfXrWY9z5doVQtS+wrADq4U61ETZ+WG29x
462EI9x55f0+l19F+vljcHu9KnmJOnBUCN+TSPCRi5UQ2GEnZHwKV6MuXs58hbog
a+rRd7OjEbvKrkzj56U3qveZ643mH0z73Mja1TKmf8wRtCtW9/Bcp2DSiOBCnJhy
h4wdEfr8XfiIsL6oNyDNKk7IOkd1a9Z6kWVSiaAaAHB99wqxkpPB+JBJ1VPTjRQ9
0SZIjx32dbQ8YknmMxTVH9y5CGI64MRD5F0qLebxgC1ZbOYet/f7dadD/3nw4EXh
dBN7rKlNz5Gc392uGPOOleBE6mCWFcP1qXeTT5tz4tCjX3Nz2I4MRUN0hejpUdw7
R8GObG/5z1soZFgd5UfqWkYcc1BxRgYp/I1oaRFzgV4x1EXII6ZEMjg18hbm3bvi
m0KACnHO6cmKlmaoQ6MB6pLbKSQ/uxvFABfLeR5jaDnY4PSC6vdIEY2mTdHQ2+Xl
awQvPuQ3R2LN7gDoecrww1HBNipR13jGfKK9uiHY58KqzotqqCk4uVPa2du8NULz
p0qoR4rl8hGMTTSgdxXE0OKkJaxh4hfMj3e1oSw8zva9wizJxxbPB3pTLIA4gW35
m0XzSup2ClYkf1A29EwYmwSZ1zrQpskOBXx1PVYElNKdYph0scRmCtxroBUHDjv+
Yk8n2vilETSKger56L6f2iS1U70ntTzboD/AY9pj+y4NtgRwdMWRDZMtuXG3/n8H
5g+BF3upIVdFKrxF0glof3yVvb8kAoOEr38/d6BHZbny99UWoCjAIl8CJsqGBCa9
IwHJ1BI5YCnuKRVHGXroo8Op9qATBIf9ZI0mAxKxqf6Yn50QCFLSEdKzC9FAr92q
kjm2bjnzgqctln76bsAYMHtv3gXqQWQjVEVle4o+Ho2pDHXNmt7oVrIA4RU2/0hM
v6blydSN/gyJLdvPdpzxWxcJWAPay2d99SHFfLlOkkvMyezlQB87kp6lGsj3GZp6
TR+tgBkEaG820KvimXViYpKrpPojZmGrw/OGBooLg3mu2LwPCwOwH+rUVZwzu/Uf
kklIvqfi7gpMe1OfVSldyZi13wuKrpHSiAtlzAtHYve2NTwaHBi2L6PH5iJDjpuY
YvSIBa5+9JP+WeZZYzmGA5cfpZo3wv3ZyLXPRYynszor9RvjsZw3BcKFhRzwdLxl
kRIpDUb7MJ5x5G8mZZwOlJraGESEWrL39GfFc+YJspZ17f3tBICcMGxJlDsGpV1S
qMgr1a3zBhcIH02WNIBsmhv8UmoDIrHwGWmJg7LTcEuA7OeA1Jfx1Yyp6C4B0M9d
Yx6siOFVpjPuVYaeS2+rUz5okrV7new3OI14soSSiw9BwiBjSCyFQRzNLu3pCeLs
wzoLwveuWDXCTOwHuvheysr1TQK/t46wk0F62VHdyxpyVJGA1n/DRvGLcdkSPUuQ
VgOcvueLmDwWU4c9mocY3Jviirf/IxkPmx/RxKxOMHxZtKaLTTfxxOFcVabw9ihm
B1uResgXjP07CPLFjMHN+06/qOusHhnKj+1oyY6BTZ2xwcxupCCZ4eRsNUYiy/HK
8nu9TmzWgH/JfWFh3DEj0hYQPI1e8+ZCc3Om6j+0P4/fW3mXob7HWS+39s3/oI1H
LAJcJDO2OuATLqhoY2hBbLE+24ot7UxvjJZ9baYDb7zow+edawd90JsIb0Lv1Bu5
2bK5S9P2jjmxMbyYyEKTaQvc/m51nI7Rkr7z9uWJ7Z8qB43NqGilrop53ko/QjPT
hYwfbRnyLxNUxZKTC6Ibgamg/WH6/WfyKa6+KqduOgDJ9kpWLfN1rCs9Z6YHw+as
5HIAKytS8HuG9rHC2iYjFLEd63m955T0ZghEF/FMCrC0wawq0iIDkgx2PgygmeDI
eN3nfn1Xr/nVCVGGB6mCpBQ5OW1uAaJ6z5JBCr4pAWaqMpeJTfJ6LXzEEPRUMGaa
FBA85fZ2YX48r3tOZAmeTqW9J9UsthfsGDZJczyYteE6GY98+5ljbg6q0oo4Vte/
Dr/Cy/pDrr6VyIEiEoHGoS2nCGXDlixF70wNbrCBKAZAUcQIYalJPQS3XIyt39bZ
KvFRP7WZYyvuKCtla0GtaD5HpLN57PXgkFA4J6eXo18k02NRocvOoEjwoVfJzxXi
2o+auvu9RJNIFXWdduQ6PVjB+F0kcSbq+jiufMkBhSkOXiAEBrdfLRz9dZa7S9ue
a2MRkuS9GMpH3MtM2RjPvskQlPw6GC76Y1ZJhaPqwb5DcJHX38wAUx8QfYEYwF23
lut/rSNLd8w/wXIdLrnWfl69G/Zz4BouZF3/DaeneNdzqRloMZP5egJgy9ixSsGL
1s1m+OLtTtvXt+nqYXpsTIEYKtikV9+jMt0XvQwhN1ydPKlntBQgg8lgTymWPNxR
vHOA6IWB8E1cBzOhPH32Le0JEVEFC3IgfsM7JlPwRbcUDP6eDiFcd05j/uwerXSA
OGRJ4wRuwRJ1mUhnqClK1PA4YI9mq4OGZGit0OfJltBvasKGuj/uXkeULP6wt/Eo
I+Rb5SM6vLczS7iDIUyMvqRFq/5/Fm7rI2RErZckK2FmWWtlBaF4AAFvtDBVsjSM
Bc5g7JarAL6sH2rpEukwT4LpTgm5Ud05CKsIPNhW2nAzTzfGcKOnufnNuUXB+s/r
y9CPqk90uVg5eUZ6HXZHTVewf4ysexNdP8i6XrgHCsDhAAQDdykga33bxFIjYWKb
9COFMgL9UDR+L5d4Eb6ffvHo2cO90kGYD8xumKtnFkbHwPK+xVfYh9K55Nqi+Fig
2fxJ0S/Co5io8hGRREj2+IxDCw2ON7uVpx75wapZWjmvrfNzsykcoO2fsgwLgPPV
qWPKrUHgQhgyOp0jyhUaO+m5Cwsnw3PlQYVDEDTBN2pO97Q9YjyxkcEnV+pawAbJ
YqEoirX/0XkKwrcZVn2iyD08KTt9gUUklAQH5C/+zzgMXAkAzOGEbTiTUpKtvjdN
Wsehgg7OdkEBHFwl3hP0aD9TtHflJx5V9zJMTOlJMGL5KxrtRju7/BSDq0pk4VPl
cwcymq0VtEn27TbuzOxxncKsPFbmKbSdUTyOmXkOpodjPFWRkbk1rTNHLQ+ihDhP
f0QpxK9heIYwweMoTmxWiUjXN247kB1slodvTL+qw/j3xPKlgiWZgp9UfsDSAn8w
RJh7NlUkxjjyev4QvCsrjk5N1OgJ7qYyKiIZnKAHnbnqqZo8I99pdn4yRXagBxX7
SbXa/RmWRb/uE+yLZh1+PhVb+5w1YdfCpEzurRmyjBHh4w5wi0gG35JSEw+HO9Ji
Gzg6FvtvfVP9h5cfBrMYOIsb+h8eodnM20vV95J146+q2H58al3TUnOGy6JDBQdz
8ZsQ+VdFoXQwQa0Vb/o/mRPH4ytIEFEEMQyOaMY3gxZ4zN19lNoEvuQkp56k0yGM
xnkALdJ0opqf9WpXYK/3z8dO3zczA7IlFfEWyoGKRu5YWAd/Z5+uX7zM0RL05/RV
/NJOa6IT5QYj85vgBdEZsx2JqWMcKGm/hH8dLaYzUMEpKP5JvngSl375CdZpnxp9
yQ8ZfXLniJ5V9DllgxYs4CcOJUXykvkACAmSIQG7U9Z9YvJxA9n2au1tjmHF47u/
1UqFOrDqoPeTkcYDRE4kP1DXGCwqLirr8NyUxg1DPBM+tQ9FfKCxlcPBADu9LScO
0hNdDICKvHS8XTlvyYFMJD77rmzvgsXzLfDaqLzF111cf+CrbSpu4gR/zquW+rRe
Go57ievRp4hRORk3umG5kL/4hi4YbdvjlIIZmYAziQi1zyQ0Q9U3K0AGm/3zwk/0
zWIVKstXT1nEn4YsM3wvsqrnHySkGPDfxWrXIsMS3z0CJnfhUBm3cXZWPnUYTHU2
EDvAp04fxfMa+ZUSOQJajtU4MwX1ezuuZ7V2o6kXShkzr4LsrNdzEFFFiqPQ+E3j
1a/3Z2wb6vpLta4Ezd2ttRa5ABXwSwXFIqdcSnDkNyHrOmJinTL+dDVk6ODDJXml
i2B5XttH8Y4WOPq6wB6Ik2SZ1jzMir+/sC8AGXdSPL3hsttjuHIzhcMb/dx4ClID
7cULJZaBKJsQVnP0IGjpnic5AXcP+7CBT3oB2lbDXuSGObjrZJM065wpiwlKUUX2
eVrYIgVYjRFXHLs1MImJVjNiHFlg1nehhdXZiknpGXJgS3WtPkrwOJfpFPSB9xph
/wOo6AKmK2JwAbYP6TcOnweAlKHdpySLMAbNjhZV8iOuOzYcctxeyG4og8KeGBEv
PyQciNOvNorkr5cyBJYNfAkwY7Eg2jC7LZrtqO7an4aryn6Xf9C540qMHlStia6R
kne++nR3HyNUTI9v4MdzA758Rpb60LKlxxCj22HdQBvVO0NJiwYmXiTd+MrINniF
uJzj+iZiiT29DJ/YhLcm3NcC+aAdZnUtH5O7q6UTPsH6531us0Jw5iqE6DewMSQ0
mZHirbfQ3i5YnCUfcWJSXvME5sqprWXNWOmQhOCyK0+8iEX+ffuFackf1cYmX9RF
LiSjbL7rq+/JFy8E4OBSRGe+7aqZcNG5u+5hPPuCnu3+GwO8hQ+sVH41Vc8qIeFQ
gktFt24W7yHhaxba5XtR7tA8elJ0RySmtYk0VjREx2E8lc9glxsvPov5utIK6BM5
RI+3u232STJXcSCa2sfkyFoULs4R3dl0Ij42N1QezHHL1gW3yY9FWGzrFzTX4llz
+eBXejEtXhHATVtRd0SJ9mg9ZFWs53Lw2IdNig+CwCPwUUbFRuH3q015m1iVAojl
1SSnro9SgpF+6vYkSgsNyNvu3HC2G/+xbnBgzlt7AdT7nWUU4lF7H4C3EpWZNpK9
fL2m3zDlXlzghZ61UxKvuWzDvhzYW0OLnPqq12vVHRp52ymse6Hc4Or1R5h9jb8n
QUjDuIUYcjsQ8Ay/0Fkr19KPRgW8IP2o7zOx3yukvDaWANGPybYaT3BcHuFOBVlz
x4XQc+eaX7IL9u3Mk6OwzC7q2yz6FPhjyMySXjxKEfvffOm6vfCuv5EfIEtnXUqD
SucRzqZkSkJM/QPPRXvnb0CyTGa1jU5HyMLb0v2qJUzN/cBFuJw7mL/KG0tnmlKA
pGDNn1S7vGj9B78yX/QOWyWxOwXfE+FjV5rCsa1HlFQOUvOiEhwx321of7tf9XpW
3bhapfg9pxsnLQ/nJ4oFug6kYp66W0s1XMVyOwKv2FW2z6WBfibThyBtmCAaO26O
46C9GZBr4Lk1Hia4tyiFLRPVvjZmtGxOAEOUBcX3elLoVLVI9x4f9ek2v0GZVwco
olfVirGYKoJCNIzfLLqjffLHDjvTbMJ7fmx2nGDKA2f5D6SF0RxJ0rIxDuSh0oNr
mFoI929IJ/UOJVqWTDVFqkvfTdRQ0KOyURkxoBiKiX8kWXxjsyhHmHEoVUIJ4B5t
LSLuI3sCmfxqdO0bKR+Zfpe4RUncl5nMowg2hLfPw+rBxgV7QlIQ21Z8Yl8RYAHz
xsAWF+VhlGlYDyAoZhhZ0g71fcmP56gsWY2A3QhO5aMe3cZKWguHISWFdj/7URqu
QSaElJakT4sZYps3csQuXUybo/O/wAio9ZJZA1OisDTGCOdQXBBFHGnbYZb3K2pk
2jFExGWuZ5zz29UP/oCp78PTUGEAbU+T+rtDU9szPi97QoTCyHgLlFiyxG5nEkzt
n2MWpw09U5HPS8In90qpJQyBuyKy04AeJ8nnuwUriQ31W0RiEtUL9AzxSm9ODWuR
Cs4Rg3AZuFKIxHIVFRv/UX3bqKbsadH6Fua++ujBnviy45Jbe8X9/M+NSzQlDvb+
e3CGDUibOwEGw0Q/gxqnb/ZtqNwjMD3zVPOY4HkMjXMI9EiAW9pFpEiMQoSwFpcr
5qf2V2jiR9e9N1aYruWs2YuDXTx/AalxgsPP+VX9tSkBBFBAGR2wn9FGDimewLX6
Fw6Oq5ahUUq6u/u5hIPBnAXsG5ZbjbGeoztLQI3RzSGxpqPH+JgETYLQpBhgdBZT
jdtAgXuk2zYeU1u1mJD++M6HtV6P+oPXzfG7OM+kNc/5a0NPDg8TinR/vlz4ALU3
hFwWiXqGt5WqPEMDylIwW3fy7JslYBHcb6EwJc/rI/bUYz8o3m6NKGrhSUz1povt
V+NXZBnjmsKGtYLE4PUhNzHupNsYHsekp7EdeAYvEFbT1Qgd1j3sxGV632oG1Ko6
/7jg6h0Id+bzpETjrLD355j/LNz7AsCwNJgMmk1YJGPZfDTzp4mT1Bc74n42nusO
gTTL/qdhgFxnC4lqK+ESJx/ze91cHLDOHUf/oWL6z0vLnANxTjgh4GVOuHFBl6s9
0cMvnErsrCUMZg/hhbW5UMpP7EIKTRLAjoHYuVVKJG6m7TH566ToZU1FMh1o3xPp
yRYI9belsUrX2NZZFN2n1P1umIqLXX8wbxRoPdUReW0WfctrcBjjjiHJir7zs0uR
Memu0B47VyvxJkTawqdd2gD4rPLjsgRLRXQ8NmMNpqBD+WTGhrqdzmBHjrMWDtr9
E1H4/3CtllfSf8aUP900QlB0IFOiCrualTdSH0jXp8ER/eBCtD+OoIIV04nJa5Nr
BdKWs2/Huthl5PWUPxH//tSAIOKsRHe6YxAFoNzgOxxCs3cAtZnqLODS+MqGcbm5
RGtB29ZnTxsYCVs2vW2/T7y5tNBenboWwbUN8c7iEqOI07A3VP7etr/ZsFRqpaLK
j+zBmI23pEPgsazzRe4SIpkceTZs9vMRL9A9vYuPJsDO4icm1Cvq1INJbV6m3APm
TE33pfuI8uysgRqTxGPrIQEbKrd71qE97ogmw5ps2l7N1OzKlzrqNOp0kFsvuU5S
aGDvtu/FkDbNgOD70JMvvEXwyIq9Dk6cCMkUl7HesbWg6aDryoAscLDP5G9XzE2H
wokGByO1LKb/Y5oGidJroWdCxu8y3YCNrhcsAPJw/MBPQUjRRXE+/hzGJrMLMXL3
WOqf+cOkXuxbi8EOwB1zDSMsN7ekmYzBgKtCZnj/qE2cs/0mfYhk+22CDKm86bWx
wnzQPEDwWKAKfmVDvjj58/MoBjw5Oaxd+wpvaFgxzx2SzbxNeN18q/S5qlffF3vB
u3sW+brWo6KzOBFJg6ZUIyDVPiLHVWwlTmLP1R62AgzuFqD6t4+VPKeH0esXZLPu
pzm6iA3uiw/myMFhEjkMzIeWQY42bG/Km9QfhPK3xuCKRtJebLE2QwBjC6R54pdJ
FSgHVbo8tvN12RZ/CGQkzX3djCVwNdl1+vI2cpaMAzbIlAx7VomJFM0nwoIzatNS
3F3fnHMs2cMbAOBMEpqTE67MCWex6HOKKJLaMlISXuYMQs+em4XBlsOI9JQNbayK
6J0zTewFTPGGk/3UGAbmZwuwylDoLLNcu1JrMs6NeWyREUkS3BEXL5mf6kWbCsIg
eat1C0Gc7RNS4DSvfO0cN0u+CX8Rh++CdcwJ+tz0sDGslun9APO/GmTgPYCWhqG0
4g7ZPWIAssBNRvc5QgTPQQk3q3OOKVuO4ofDB7VnV43LkHfav+PvrxhW7LRUzIm8
/dAs4jlcnAsOCYPcfuBQr+y/zZCbso98U5n6yYVwR4Nch5mbQpjxPV2DuC6S5Anh
mSyL/yGWrB4CDtHUwB34Zj/sPBFgSBPex8DHY/we/5JdpGiw9hhHh3GfZ1DVEmgm
Emv7vWiKpZunWJ+wbo35BuY46FBJjTD8m4WZFmjhHKSK3sje5ItGlgyGuo4YxSw/
cDYNoGplirI2bg83La9/Dh30qreetz7/mVm9raRsitHLt/Q0BoyQ3IV6u7XpdYFg
BlTmmptzoffuncdL8gxa/zZDxOSFqbgAOFP3+wBrEoVOmankIh+qKMNRQQuWvIH2
jZygJxz1wpCJpmuYhm9CYs1AuXkVnL94mQtpRTZ+On73K9MU5cn0NUldJHbVBmMt
aekUxDyCKmoFYuYo2QTCFCwdM8bfzE7GUKN2pdY9uGk+BGZi2NzM5jifQwJuOZPZ
kA1ZDpDcYdR4Hu+Sx/6w6qUDQd2Cbj1hV0OrHK/E65vq9y0Ko96uf2jr5IQlnxqr
sO8j3H6fNsKmIz0kIrVifUgvYvY2HHS/k66rVFyIAOGNCPtjwLoucu4cOMfy+Bwl
m4NKoA/53eeHDgU4DgSzc/Ecfdm2s/yqM1xgTrRHF7rvHENvCvp9wQw7oAZaKX31
xpz+t9l/9RQoOLw+g9yz0JSF0dfUlq4LCaFQr7F4H3TyDYACii1ASyobkW1lCUOM
RVg6jvgHXiFulAhhZeIPbvZca7yvNBi/nlSSFn16xvus6F6TCOFDWXkl4Plccgrf
Sx/V5kYBIeoEyKs+cAsyf6OF9unX0OkO3+EUwaReoP6H1j4a77D2e6sBaF2Jb7V7
LoeIES2nzw3+BiI5udUDKOVjpdH2Yc24Xx16lAa+8M4aoEt4ukHM5pyDixV+C1ih
syMMYOQEuElb5DUebOhmLLomdpIHazpuNqcfZoiNPC/T/K4MCbEDL6J4MpB/+RFa
OXQk4UWiDhZRM2wMp0fXQ8JjRuTa4RSbwpcyseW16vqHGyxLfHlIQU4PlGcVsrAY
kiOeGBqHyIfEvoyPzhh/j5qJ8Wurk+3oqilCOlebhLyfn5jvHzi0N79ugKSZ+p/H
EhJTdqvZ8QVG12I8pW/QIDE+uxDgYy9L2e8/HvdxrAbJgyUS3sUBaBAo6yRXhFlQ
abJkJe0/R8qGHk1ZA3PJPwRJkzQFM2TejIjxbEfc4NAgLGsc14tl+7paWTabpTaT
6jfvvzerFHu1deQVAJdjeriDA/4yM7j5cZCJdwCRiAqnQLaTRf3iMfNEF8tPmhFg
N+i/d9D6dI5PbMuGdy79wOqZXNqMslriofPiuxAN8xLhEKZKwSZmbp7ypOhSrEdG
wjDTFq/rHYL29ShUVYkX60K20PUNgTabzvDmfETTTk27ySWA63ra7VTrDhynq/JD
mIvDjElvioM+4tucStnuS7K9EucJJnKGSpKc6RSJSs3hHlRwpK6AWGx2O55RQjJl
BsOtP2KNcqG6hfvTx0KXYDRZWzDvpYpYkDowshKDFIO79ziq9Ka7sKCYGpea0Fea
T15RqAs8m6pMlWsiCFSsoikibYVohTcmsxz5Ca6BMGedn+HWHfso+aiYCQwDtoB1
BiSXJ3upNrBOf9OHLzb76VhMUq5ZPh9Gr+ZjqVtF/g3F7mXvWr2/pbv4e9mIAXdz
n3kJkCa09kI2Y8UlHCUNUihOfOYvdfJXoT/BMPHBjrmtZpPc9uoviJ0wMWc1kmNL
IQNRvPn3SRxd8cDKCN36Lis9WnDqJsbmilT4561hwFRsfat+wodw/JPcTneCn4xL
cC2fnH3P34UZ4h6aOq89NbScYiKIs62gwx+qYTu7vH1qzauZ1Wpbwwh3ySqa19aj
g2Uxd29kqUpnO+xpSJS0BZWXhJRYxrhzB2k2YwaVa+hP7j1acDKEJyW1YbosX0ud
Vl5sw/798/7ZA2F6cHl0h1jXT8ifo1shUNVnBiJg+sX8IotzTGYe4AYt5C0MVbkk
xW4X3Ink2eFJoEi7awg+ebnGb1lP10FoCckKwc4YiOGIn3Jg0b3LuLlEU3qcspYJ
lFndD0+clo2qGl4XNOK8v5L4QA6dLy7ZZ1D0uRz39YGIk83J8EYBKUDB5WzcaLc0
ERMwuAjrxSpLnx+OHy6V0MF+Che4Sio6AXjqSYgKEBT1VI+GgO9SNxwck0yAa0X5
CDteFHDGoVbyA2vCf1IY6TN3FhvuH/ZZtxGFmkzOLr9gIG8I6NnRRFwtJhdJXOcg
MCXlwSlfDMTmdbp3DyjLeKz/9/+m0wQbxxxKAmsucP3waHh4rmZFgEaQAP52l637
OY3gtHeOSQRNpUYY7PbWrex4htEvVDc1GQwygCbh0M/GSQnLHkX/koNFGxCSKwGU
aqWq6KktlCNfla4cG5pnyUGQpyM+SRR4J7E63UyXgw7fVOzlvAjKtsNiAyJzK+Mh
aU9Cob33WGwaDcjgDEy9fcS+AkSl75bA1sVwLC+HSFlSwvdfFBrLM0u/HdBC1ie4
wnLAmfymiJ/felWashHRgpxHmiKwvWD3rYvkCaBC5d2SA8BJ84ju9vUg1zJkiMvB
6iACtD8ZBYyBXwRV5ykaQuomoCEi8znedYlC/CDm9DX1XZPx+tS9hyKEDr7UI6zA
yWs0P0ZeY+d5lYdLrvqSzaV50yKDW0KgsnVobRyqMPE6228Fc5o9Z1KBCQQKYe3w
pVSUNy0zuqCj7uhCZLVnskqWaPe/j78OA8fKAXAPYeMmCxggCw2RDlY5KnwhGW2L
fYoq3k8DrNVjhIaBO6WzjYTdu8BfhsBMzIc0cstRHXw03Cw8tjwjs+FPfzsQy/VT
LH/3P8nxtWYE8j5zB9pmqNCSh7JfJAohstFUNso+83lsCobuyY+d/JQhlKD8yK7W
ceWTbjfG1eg+KIJYSK+cB7shXxhGgfMdJxRws8d/C/udxF0ZyQwtk/14YlplBKmP
o3fmqC0aU8FaGL7F/UrLGPHn7TbyZIJnqQdqN9ro33V6z+6thqii5S014a6c05Ir
UfHT6ZKfrZJLnqS7Xxymi5gY0lLk4Z6EsuGhRVwZJFi5t6baERp18hkYos2DAldR
W6G+CneYt+16JJ9ohqAnU8kOanuN5otidGivyc9h7i6/3g2yRCwGGBL3wsJIdATP
S3e/N0ps/XaiL4xOjjIb4jvKTvmDQCPfJAI80TRzjpvRPrEnkJJs1cIeqrBorQPA
X5xnZniKh0BcWaYmzHFQQdRyRRVuHp85bH/caK6LgSuF+q2GQdANZQpOfyT3P7qB
M+4BVGkEiR4gjGTSvoH5us6oIOUJdY73/N1tmGwuLckuBm0QHK0d6BH/JBMVH/xQ
M4Ns2bRkL6J8WzF4XhVgV5j9lC0CNyY8eke6Q9Ec+sFNpxjaGAmzHRfyxByPjYGt
xlqhzCakgrWwYQqlQq8aSJqlDYd+AOPhcJWBjQPrHJSikq8ARcY2WrYT5b3MRGtB
h+pj22VNYX8SdpHIei3mVEAOIHLU+K4JektuXUxXLWixSaJgVWZjGlX+JZUvsnQZ
XlBLuTUvfMnWwxvUnRkd9Un2XcwejWf7Rbzlg0ysteWCE+NwxYNjISiNgWKuEu4P
ih52gtTd1yTilswwPSZAKVbjrdRdiC6a94l2/7Lo6HukYZAaWaiU7UHYt/k1cUy3
cISBeFZFXpK4kfBSbHUM3jnqdUsYZAXkZZLoqePutgPnwUkkDITyN/dMi0rJVJj4
CnF5GsBsKaQxtfGbEVXjMsSDiOm7b6AEkr8MIMe0z72YRmisC3vb1I9EA3HuNGEy
vP172m8Mapn7pAesMDJOjZGGCBNkfGE7Ul9japrwxvbKGjX18Qezmx9ApMonLKYA
abhDR4ym6b1QusEbXj8pRpT5sCKJdPzJjXXJJ/B5fKcLJjW+eI0cCireCEG/epui
GPsTrSXzM5PmeQaykAeqXf3iPl4KqvTNazh16bgW7E2Uv1pJ2njfP1KCpMxTJOGy
kabCG5ml9oteWX/Nk3gwSjZlpuTXxNM7kHDwe3EnddCVISVgndVC5I7aXfNeAvs7
GA2DSvd71HQt5dodBfZcIuFh/PLGtThjn6d7src0fxAPIFYeFyu7Sl1X0+LXWYk0
6EbDQm9DBui4LlCsFNyKiSS1AiENybuT3xdPyMOHt6HUERc6YEwI5mz1H7Vnyi96
Qa6wIGvQQfji8qRZO7h29Ab2nVVRjHRNEHuoyi1Ny2byXgPrcnvhfYJ/RHbqxxy8
i6csT2LdpESSNcJG14xw1Fj2UCLqCbooyGQmAyJ9ws35Nc3c1k+yfa1OzYcpc6dl
ur4IrYllZbJBYTRf906z4lLb/CW55kkLPBsbIu8tEbOYopagI04OotsQkColqXhb
gZC/aw2D0syiRRxf+JGaqIEcHW0lSz0GCxoZDebKMKCvRKG993LVXGofVSud5rbY
AVGy2lsA/AMlIBnqOfWT5v1lmz6CNZsocMW9SGWH96lOHxpqOu9IhACTL+rcy5g3
mOiMIFoWa1zQokLBMpYkKeRVo7UCGg0dbReiWgfpDTOwbOLmJggenaMpfHBEoudr
ZE9xjGyRBWIVpWVw3fOWWTPx9bPfrTSUBDCftc4bQWq41QSubkYGFIcHXFf71gAQ
msp+TKEFagChRQMEkU6JdaPPXgCKUcOw6b256DxTbptqUYeexF4aYLzBjigVSo3T
a8WJK2P1J4VLz1DCwzSRLLAnppP3jOZECqgxlwFjQaXJ1FGwdZhQ0dP/0XhuXhIf
y/DD0NnYaTH0w7h8mNBc5gN3jjrGTJiApVwU2ZNScUFZW+iz4XF/d7/XjhBVnppk
ExzAQ6/2cvFPFHiEzjm3NhtlwPrZ9Wh3avoLOsFrnBANBdoiRINrnxWtoxlyn8lR
KLH/LLnPzB5KtXusSx1L2S+rCxl8gHshTJnCrSa/Ir6rYXorV387tKdxnXRIWeZR
c3byZdNuKLdJwr0ywX5tYSuvxCh3uJ68PqJgx5qmb/IcIfFIM+b6mbXjB8lOxWX8
35KHeLnCLqrXjCY+7VIVRy3ZYhgQ7dDlJLiRplkFxWMNkkViSsdLiWTJeg68ENpz
6m/d/NTLPt69WNc04rECWvuw6vfUxtslQBUWgF+dmvO+RYteE+TYFkNHoZFaEKya
QTCkWyUhV8ECxYmWW9Zljv4DKiUKZcZvfjMRZLvGGN9MHvZEPV40KEoKtQIr4WzP
ZawvdXLfc3S0/6Z1Cunrpm70a5zg7pSMTXvJxX80CSmvaSXSeU4MkSnmtKS4E3wq
0RcAACNxOfPS8YmWvjjtZbzT6jlxickgLIt2euv8J3DFJ4gv1K4jZMZHoGY2AlvD
qa6+MZHFg3h5xQ/oHrchh3bhWBn4Nx/W/dN84q8md9hKqj3BgXf56VFDgE8DirZ2
vPEm7iBulOQR7TRRbjcswri5vcXA2hIq1RLaJoECDV1/iAlGCc3jrLql+INIFje9
DDskn0dxr2Q4xS3lgqDr61EReI8P3d8xnS8+4+P313X0EMkkldlK1yVB29mYaEs1
sb5xvwg6KCLJzAQprxW6q4Gw63nKOWgRMSp9QN0BbM/2t+kFiUC5TvGM1dnrpFaz
6tveFSmX1W+z0xxkXKP6frTftpBtYtBCWGBIAAeWNqz8YFXtS4YY6m2cRLqlXxiY
o1rnzOZ6CKDCwtFg5QNmgZz2/8NDCdMB0ZgA4s/AiFp3UIrGsczTB516YtUWldJ7
8x1cix/eZCGUV+BXd1eepJqFLU06Vm7VdgsP5HBj6TDM/kXUv1/zQMduoglzSJYy
O/2VZpTFskFoOUYr5Sc10JZhhn7I0749d+BrkNd2ZXMc28DK030d9lA3cC93Vaqp
8bnsCNvxNRBfpdC0scHyp+u56qsEi5bz2Ey3ewvbvek=
`protect END_PROTECTED