-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Vvt7XZYPckCu+VTmsQpp55C9H/AEZhouHVhWsf5B8ZND4GmdVkHziv8k7oXxpKkn
NI/tr0Ys7jkJk/vi0aVcQAUFPBoDFjYma7jUaa+qskSAM20h15fTYYiKlME9mSYx
3hETW5VsH0iAl//VaNzn7W/34HbNbngWP7hSu4AVkUg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9180)

`protect DATA_BLOCK
02mFd/NsAZxTnbiiAWn2WGzSbb7cmYq4Y4vC6qT3QQabxfVN73baFJeQs6YC1gSY
eLO0NloO6USe61zQany0xd6XQgp1Ydtk7GyGVnEbCobsWsEY3t8vG5oHrXJXlfWf
4WES3c8y6do12e1+J93yIk1i3vU1MKo3zDRYKyvsaZgHh0gtiNHX3pd3TX8Mzy01
VcIutAgrjgJu2HBbPpi7iB0fKmWyfAjshZPdfY2ZSxkleycBPK6wIwwh0SzKiSN5
uhURbwDUws7pCiB0b6hoH/YrcVj/YwjVxmOaVVSTGGk1uQQeetqhFeaxTlrbeS3c
ClThGEcXjjKKzvLDd5y/chmDfJ1rqChD3wjSsvVq7JvxyLkrc20K+KP5RyMN6LUK
7grHM/RMIIb23hfXK3EJ0aHNXhsQjZZvf16m60bmJXvV0wB3NnaGKl2ejc1o02GD
+u+Ik3sCnDKJB+ZTuxxo/xYtW5x55OH05+vLqgYPQRRWunlcOsCKAHfpf9nR2Pom
pZMQsm612HlVnq9KHRUN0wtTgVBazkkUzxhiP05AYaGcqeBI88/kVsoDxC6lfjpq
Jpxou3z0Kgsu5aZ9R5MiNh9eDBJah2QNlAU976iWCoO/rJFv65182otGrEaPIZph
JJKTQbv4IIeGhdVE6jjqo92EuyqgJoSMU+JKb9RBLkjY3NsRkwH2RyuTvRBniHp1
rCgwKksi/bgwITExpKjj3t4WpkJTaozWYha9wg0mMTzk6Yq4oC+H7ON+fRa5kxiE
5mPtggNgx1SNpzcvA65WKXdC0Purb76Y/9adJyxE1fad+m/SIpvh65LsRFNuT+Sn
3SFRfOxZ9D48bCaIGEa9XSD2HVYHuXRV+P9/JzwRboJQrDM9cJGTsIBozEzspemj
04uUTtRIBOr2xTyiNWD7EfUbNQz4MpdRyJk8dMcFWp0oOtOgCWn3Me6pWqI2XQGU
goxdj4h3pTBKXamK8ZyzoAq2NsKPJL5WazrwCZHp3m1qoVQxfqBiyqIA8+yTAiOv
i88CM491SX5swUUDjH1wBSarT8yto74TvQcTzBNgXiLv5wbiVGqwwpDg8OYTFmeU
0XV78JbKs2edmC96zpm7XN7CPst7CUhYhD0MuqhnkUvCQmf58xgvBZuLpSIqVECF
gOyS8+cw1ktprpyYFPvnLs3DTqaQAHjy2xBPYDnbk878kejBLIByuVTg4/pmqgXC
N5c/xFZST2msaWY4mzDDIkUFwhnxjVCiewzLSoZ3oa2bLf1S30gg8tEJphcCSFTa
wpSW8cAb9U5CgCf6rj94CtKFkU2Owwp7BTuDAw9gv9sy604DWSRTwxlkzb26fZUZ
wKW6b5qKWkfpHifBWyiPp2LNCXKcxOu5Rr3b/yhyQHSl0O+wSGXAxe18tPPSg/GP
umd+PTL5pBg0cbb7tfyGzvILhBBBCWFG5x/lrafAvqE3B3kaA/8ZWAcze+oHmOkz
W66GJxtVvFdVp4bJW3JEiSZfwa+e7qrudlwrVVH2L6NBiLPmbEh+jTbzPA1kz9Ms
ASWnti0NtnKI/tubsiBix4f21ZcTA/Q3p2rVvKB9oOP0M022Iyt6v13JXgACKiPS
kajaPjPhdUFOz8EPjpv1sxPYV9dr6qEUNj55+Qdgr7WdsPe/KGL3RGTUqUKB2VWw
mxD5brSh/9H2NeAaGc7yVa/dtN+y4JwyLeRuXo9U0kEfDOw+GcrZbPGXEuoaSz03
9A2aBm4r42phZQJd9jM9Sm9+0+9nbPiID8gttM0yCfhyDsc/JOV9RfklFoP7iefF
OZirtDDgG2+126FRvRkvERpeEWqLVT/JXBHjs3ruwuUgDleODGrCTtzNDGc8H4WW
AaXOUrcGEkvTJc+Z5hMPimNhNNhge88m8JFGGx2cVsZzj9BWRJEh9kmZEeOZz/5D
bVMvMidD7YaEIi4FmWgFgyywVrim0OIVCIrHfDH8iCvcIbZT4kiQv0k784BB5REy
FIQvKSn/6Ho1MS6WDqfdtEyQwNkTIngVs1fA9umNuwxWGn+XZ+VYv4ijUpubhKbt
Kue4K9GgkNTk8apYQwHIB6sE00nJ22qZkttEm2IkyzXmzQHeTGgoEqEjFpqM9goZ
VJrbzMrT7f3/9DTq8dNu+UN/GRwBXMw2PasNPzNSIyesVs+AZsDJ9ynYQ5LBvVy6
TsvIofpeZS2Jn5aNfGbkX77Pq1mYFTAtImHcPHXllAEdpANVlXJwQvd3gUaFrTwf
alHoYm7GtbzzBf4I67/DTaHVrbmKdkXDJ5S0qflbl0z/j6uZcZAgLzqQMd4T1lMw
IWlDdC0JjrBx9T9qRGijfzdWdGDv2sWNp4F1R/3Y8aGbOcBxns1lTtsAXEA/ct8q
LEN5XFqAHut6nIroYXkuokxoGw6vkm/hTw5SvrV3DlJFDN3JLPXfFUPxNDx3/9BL
sMI7YQnuOdcGFLwNUjGhx0amwNqC0cnnW2DnYBQBDJX+d2327iYuniPw/ezAD5cS
/wElAI2cI4l3hbg7VytaK2gkY62kyepL5b+c3KeAYH+Wl2hIEw5vaT9yJZuhs73j
H7s/IWKqB7Jdg1dVCfLAdmrYwkaY6sTF284JKtEi+rbpk/kIP02SHC4m5KoI+BCu
C6qoGTHW5g3uZn/AcT5M5GXabldRxR+TODFxraY3i4OrU6r4Vtbi0ZwFw2cFVKc3
TUYKkYbJHjpeUjxszfrKT/6vZfuXPjPUpmKhJu+3igzlDxtyh7A2ehwF5etn/hFA
sUbpo5wx1HCmcl6MlCq46ccRoMLiUw9oK/Jhny13KvaGhaBKZ8gPKk4nTRRsLVnN
0Yl+QSCqouHB6LXd/JfivdHBa4s/OcMQbme+EzewHPk3Ehx4Hvka/m+5gcmdGAYe
hvPnEqAjtAh7zbiBhgpm9/m5C71RjyxyN53l8RYuqvV0F6dyTVMJdpMRU4BiUom/
8XEWsyMxTfGZHesHcI3q0kMLdtCpHeSZwCYh8QJnWUCH/dJoNNG85kdXq1d6sZiK
2x/vNx9MTqzmEWMyBmMU84kWHgpwkpAuyynkE7QCkaHVgSh0+gCKZx0Ad+/RGgYF
/21p97yJtvzZIrQXA6qqbKg3Yy2APWiY87XaxxEvGjBJOtR2Iqp3Q9MWaD+kDZMJ
/JFHzdFGV4ZrhhmP6wfenldXNFHSeF3YEm5zsztqBuGZzwCco3CDf8zQgv70AwRs
vOrZly0n/FJutt6pWZi+yi+mYrR73oGiq59/RL2l6iJwTZLzcy8IKkLodkGK4sJD
WlHkp5r6gy3ICyY1rBKvjQwnfB6B4CyvYTAmtVy/+vgpPEXe2asgcpbIeSzXVXpp
P5flZVRfvJvfN7E+J5C9YaAT/BHxqWL/b6Rp7xECz9mQgbGFzwgcHu9TYcATV0mO
R2hl+3bkeB0WwMZT7k0d5JVvUOZ6ablmBLJpPRwI/DnqaXCan0bPdlqE5U/1ldJR
6RG0DBoXcRlBa0ya/XR/pU3X9UkuWknmimausUZOy1XVQbp3MU4+HcZfPoSbfzfM
IJzRHUUKIDmQYF7ELIzbAOvEqxs4hC/E4LADc7QAOzzkPLVxvBkY80YKKMG8wfVS
/OwL1qZvNhuwqPVHndYSOyadBIGumQRGMlRO6V8f51+EnA7HBmxWStc/212+Gvrw
wyVjPwY6UiezY/zlOgzT8oLwyNG4/ia2gKTx7AsTb1/s16ijllbYmmgpeQcYUaFT
XhwY+HGDPr+TWCpLxNC9tUDw8zn62YVNTyxP2RC3pkvM8d7Y6D2qMaURp0sqVZZC
nMV753naxHH8duq30Neo2cv79tp++q2B1LwBqvmDVodlhY0NC+ieqEldD4KYGJcn
vev62TzGaPgwqFNBCBPVTLc4BShrgXmNed8wVJhWKhjFA8flwA7AlReDIaRR3UBf
XnofufHnmH/JwpuatNzs3FlnFlIX7iAULhfQF0lWGjGly6A9BcgDvRmr48opscbb
bNkI0mNS6zG+cyLtOdyokI3blAyzqgq1P0BsC7346nckNkV9kMBSROUXCRLaWyn6
lueWQm9VxPOePIoYF9Fd8FrqNfukP6tmNVy9af+jMemubE5LYqTCTzyWY7qvHkZY
Nv3lbwZH1ZxCG2RU5AT2I/4riRDzQXtMdsw4Xsp/vqbOu3VcsDCaiOux0YOs2Cok
QE9WamweGpvE7H1bnlWaDGe7Af9/PePRl82QpWYNhL4736dQsIYxEdpWieGvRyZ8
8tKm8D0u3NcGJrUFYPG4x+YzEWOwB2miDx6HIq7LnRpxmUhpOYb4CQ0xkFz1oStg
wk2NRt4Xn+GrCqAj8oKJZa0YfTIU5zYc3GrcNXLlawW9qASREr5JhOQwY+l6/f1T
SP7IQG0v3ZMXNbzcAJLEILtimpI8LdKvEf2Fnqlmatwfc4/pcQvaMfITJoOoAKIw
hZbiryv/7R5kQMPuIomcQMI3tog5dpwFfuQDuh1LgLA4UtfEcGbF+NXbutdLL+Gy
EbIw4nY9BtWbGsiXzyNq4MEQFcTNmJ/mjVoGCgirXV8Y4CpUvVauQRhReZ+CtxGw
VZUDDUkghXVjLPGiw1iHQTlGJZUlgOuMJ++XyPMiINYfDYFsu9rqaekurH2akZoS
ZZgMA9GzxCUds6RauPAifw8//ZOYgrWEKcdNEu5k86pbXcqp+KHqL6Sur3ijueYm
3lmRjtcQ9diY/V4KHwJvQd4stNLgD+Pm+ot5hNW4ripJmcNOJ5bQF0OmBvtLgPab
QPaJMbHjCCsePoVskX+muAotvw2C7GlJJxvLBD7ZmSNoMcLMMI9asuNQFM57dubH
m63eA85n1lbeEsOGrsvhI9JV64b4WMqRDR5bUcimBJlVu4Ivm6J3VPEu79MtrAQQ
uNiy+OEXSM/Kv+QJcIIAtRy2IQaEl1qE4eHl0/0Wx5Djm5xYT5+VFkRmXh9IssPq
ECsWOxuA5CEUT+N2VE52yalq934IDVIHBtJ/6I/+G6DwXCzNmlBeVb/Sg/citOgE
NjUEtzepNCSus4pZM0sm+cYvr/tm7IGS7qMSQX40Pk5vGb/2Tb3Mjpxy0bR1Bq8K
SaPJ+h23+RlsrMFppbImkLXgZLhA1AD+LZMzhT4tH4n5gvYzu2f4EzHRc9El+YpU
VJPw9xrSyFe98IyTmlBxuWRL2YlkkL6sEU4S2+iRCaa3qh6a+ZAiZtP2FCfZi8We
0oVoXyAX2OlO44az6JFqsnZ4mWnVBuSYJttAQ0g/v67FMyAmm250HFhFmiM8SZO4
Eqv8SofR+poz1g7RBd8VC0MRbBU2JiInsVJVvB4FgAIOmKSn7CTGmcXPaUdPUg4m
5rBjoTeE2cN5A7mkvgX24/xv7nB94GV17A6TtPi7gIftd3pABi6hZP4qY8y6ow+r
uVdDLx0anAdlwMWU5gNz+8u5XkO5G51ytoANwRVHcEntUrNCRyonWzT/ImRF+0jw
L7mOgx8cwG8dx9qPPgZ8PjU8O5l8Ewt70dSZkJrBmVupmaobDOA2JcD5NJRlWDE2
ZK7rZ+1x5UXepysaXALwtPRCJg2ITzjkULTiMcnR+o8pYfe8lUqYbA0GHFOiLBgI
grzpEm3loWttSs1r7kmag2EFRyUtnJaL78fMYMe9UaYi3u4B8bmjUWc5ObDXe1y7
6gfcPpj9O43zkNIbbowMVbZ1EvcyAPifv5CEdSo7OYxAXhB1wCuN+5Aq1AKsn0YB
d4GuA8i7PJ4ubF6xfSssTWRJ33LFspPwLp2PlTpbtS+pbVeS1g+hH7UbVesHU4B/
x89qu32gUkfCYFpIkUtv0i5z6rALMWVH13LesFFjcqH/31KhCQwvDThzxGhWY/6B
+ksGvVN9NXZmeeNKlfptNW1a8sbBa5I3Jpl2W9ltamKeAh/NR3+JeRkMRUMs+oqj
PP21ruiH/3+2AeI8Uu75/8ZRyxzCMO6NcQKNVZSRV3xk9GMci2OCGbSiqd/5sJuM
THVuwbO7zBJVu+05jDsLB8Ol2Ssd3rMrD9s6WNvg4OIG5ihPdB9tg/e1Xk73WLZK
u+Wx2nT+klRMy1pJPfQxvfxSe2B0gbmBnoIoY4fk5Kf2j0p/PzKNAtW7MwEsTVsy
h6mjsFHnMNKG/uwOPgg/o1JBDvP0HSvcaebPiHoHOzMc5Zd7SAMhJCs7/b73G2sl
ilCep1oCae45SwMC4+mDxWBzS711agA2bL2wSTCAF3hwTAerSOg/ZCenvePXbx6c
7PlxkaxbaBFQQ1xzaGdvP2AyAUx572bqcUDXG9zi+Li8EvrcDRlh6yOFM8roRXoi
B+OninM7kiHKolvFu7JxFWf0ZYs6fVwT81uIBz9/PfuZThCeqQYFEUL4AgqMA/Qa
LmfpGvormpb7R29irXk4OSxG0MfIBJVY8FqxX9QbaK9CP7chGaPylDihLpQxQkmR
p7LFWtHlInNFLDUEGmFdLbO+C1j1wlVtQ+n7xAGRDS+cPrRWLZmI6Sqqw20UK9vg
pjPSXE9W70JtlB/UoL7dff5Ngj2dQ4/XMTaVyq7qiwFAr3sifMgEwXumy3z17+M9
TK4sX6h/ESGANAd4u42w7mIwZWLfnfh5cu7lkmINNC9/qm6W3LQD4hqkY2Low1vz
xSKKBYlL4Y/toni6a8SU0r8SsSSa5rKJPyowtJhFydcxLPOVXA7ArC63QIPyX4H+
/RsJ75qSJ/W8wZliowLjI99qss82XMAfFf6auWEBYlQIdK8KmLzEmRWehVcYuFtm
gqzldXXCS1llN1RamgBh+9xmui99wdY6zLyofLUeWHvDfP18JulsI/pdUAO3m++c
Dc58l4BXYrs/pbTPqeNxFu8Sn9ibH94Z/yNTeIX/9GsIeTKhnxAmqDWrd56bffW+
5L0W1M0MuakmWOqaZMRnKpqzX0W9E8T6N+8/yZS9ILb6+YIjF8eUVPmzlRaC9YpU
cOZVYhivwKCP7aSeB3ShophloHeqpE93TVA0Ad/hLpkt3KcJzQ9INjmXxL/fuq54
vfUGIZkjquxXd6GyDfM8HECToxlZNt0zhwzXyYXvgFw2X9vrtpiqA3gyb82syXDU
h5mLtSNOQQDHQ/Fi3dEqmluL2jgJSyiY1BY5Hu43S5E5ErrnLkjJNCzOk0wQ72jN
adf9o6a/rltfRsdT+O+I6tVFJ+7Tn3w03VOzigCMXxk2eYLNYiS3gZK2WSJMxmAS
xBSreBU7MWhbEIu1TX0mr0KEQKoeE7RXGiNCdrwsaPUpgX+Tbl+sXYx98pfPWUPN
9ksDAeUSKUDDAl9yGkB+9e/1zguekdxhfhi+lo6gCW6b+H1AKaoiBy7Gtvj9lPPP
sniMIOe27pQP61mHZtwxa/HmSFenGgTUIBI8h1WYpoy/EJxrZLESUMWYFB7sZ8B5
84z2sHaG92VoVehlyiO1TN7UOEwmy0RRI8bIQfdYwEt4+BIKsljRkEYv/IecHBr4
yBFYcOjYgC4cLpRO6gSZP8+BsPX7hyrbOOpUYTZTHAb9dMYhqPWtaAgZSe/3mMYU
9yWlBT02ZLFhRlJbcBMItIEv79FC6xmnfT/o0pqYnLdJhdqeEAPKjFHgHaV4d3FO
h1yp85hWaajbmidNPPxKRbsNKNMUv1TX2dWGK72y0UNZevCTnNwVkRcF00ic6Edq
ncTei5/oWZFJSSflKr8OJTxHpR9zMpgQ7kyUuKqiuydG867ERfV07dHb4XVTsFkM
3pytVSl7G5g0OC118khGzYAMCgV/D8wV8kalH4FvCHjaHBrAe2HUwcfPftYvZ8ad
bBR9r5bSZHgCxlIVmpp6iz+/byKbyU3s5TLFSuLORkJxQ145L96L9yXcPkUIWQZ2
guz4wzDGjs2rlCZJ81xn3bqtbtdx1Bsa11tkb570d5EzHJ6SclYhQP9WDkxbjgsr
0Z7Oy2tkEZQ9AtJrxILMBo76o0mqCNYstPA3e0nemh10l75SAJgGGGmN9h9HHO9N
3+k6EvboXGkb6ZgdQcDO5VEHug3G+uzUd7CTnom3DGu9AQuXFnfhxzkb7VzWN/+o
v+5Dwyilh61kWkdyUNZ+e+vUM059aAQ6gQ/L18OCsLeJ9Ugt1t8BCquze2Aggbjf
QlFzk730FwUHDS0BA3PwpODBn3hOcZU7vSTrIcfFq4sAue2pkwzonuPPcMWjqEp1
bifQ+Azu1nG0/cSWZy3l1hucXiWCkN9Oo9FwgNWym8/JbqQn1vGv+B6PKfIUIN56
CdExYZFNapMgSnoP18taer8SroyUQSr69IwP2+RUMjcMK+WPFX9gZ86fLb9q8oyv
6JISfKxZDHHvV2YvS0JnxCsLEf/trI4qv3MCpd9XJeKQcnbFszDHJ/q3wDY94W2+
24HKyU/6rGxISF5lodIJtSTod5d+ASDeLS5c4ukmyOV1DmZhvhHIAOLooq2Hkxin
xr4NvvIsMijsnteb3nn7smdd9mleGU+G5aMSL6ukU7qerdOQtLDdGu/Ww+ovHfbj
63s4FZuTA6dFBsEsIxNSEegoF6W53KqjoooenjzL0TbbDp95EqH93d3+gTof56bA
g/dy2g1WgwhwgpI50fXdRFqRT2JSgp6kFK/XHv7RigxEu61qdvq25reE1L0/aRtZ
2ugw0cg7iGngtLjGj3jWFtRzZUPlCGb6y5YkXbHvuCiUzyo5ynLODF/XnzNrxaOM
delCIyvfVgfSf/9FcoIQ4hRcAOhfDZhk+RtqF+rvRM3KGLs2xziJ+9yCPSHG6nmf
AaMIw81ib5TSA+CVxMuSX26CYMkhO7meOruA30UanBxUaUvFCqDndU8FLMuDDkyY
f31wNMSW3iQsn1JxcKDHo1XIPJW20OTpOrAnYh8MVjJ3n7Ya36xa9UABvYJ7Pn1I
oHSUkoWFD4pQe06tMUC8S+3TKsc4qcymtn6fsHDlsXHc+zkj+U5C/ZETA7HW828W
kQGwjuyCIHyLdZMYYvbDdTYdDiXvuMCJSbB5rfcmLrLcqR/IJc+7cu2a0Ra89xBd
pAEUaCRl2sqU+QM9+yPCzK6EBiSqZPlw8+GQ3PslJdfp05LP6eZQFQtDKVsUfVf9
vRjG7p5Wiql2RX7Kg46EPtniQXri+P/IZMVj/f47im3746f2/nLwCU3OBy/Hs72F
BGPaXnuSoBfSL5+fwfOzGLuxIF8I8a+aqCB2jXbVLkkZR9V0PFYJFvSuQh+6yRDh
aeAkpFNP+ElBuy1OGA6bVtxncG8SaMiCI6eKTdMfSjOMwLVvUk+eYXY6u6oKCzzI
AaxmbM1jbyey8+GrX4KbpT/MtKirhRS/HOuyqpsSPZOA6+y+a+2y9Kp8z49CbhHj
JFSwyKtk/raKrj4Zupi/YEP9gAnBHQECUDg+/5F/0uodgaNmhCCE3pn7xHAmP9rK
i/N2aqSbqhVz4oWx4fO0b45F9nIVBvqKCrAkXS0+B6RsuboykOfWkkhovk2VAheG
zpBliyivtQrXINBYXCyUBDuG5C7ghtDBYEIqTeZ/mKELZ4AKKoDMKY82FNp84NSF
1GGbuy7ls7hk3HC1boEkCfzqgbk3V+WFWlh5cD6eC8LypyneHqU3nMu+mNXXREcz
cecV+q2kac06D1HgxTcn6d6oyBEuUACJXSJif65x9XgwuBXr6JWmfy+21VngPrKs
9hSDJ1WKgJ0StNntFrB69i4eognPXYZQS81GdM330i9vxtc84SyR++Cuv/yzB7Re
S18+vBkCIzl0oBXKGSr4PD+x6BwE8uSxbKuSAp2DtNGX88xRElgxzHd0m3IlZ2uZ
o/bXnVEVjRlqS/odAWI6jkY8WicLHaV+TONEyswle+o7isusRJmx1wqTyo8s1yK2
HGlaDgwOCZDPbuKPVIaf+2oILqNXPVwh/Sk8GpgTMcyjaRZtQ6ZCnFJwi4udMaHe
YFIrtD6AX018Hp13ZXt4Pi5vumNs6+wgDu8U8t2FtfbWLOoIYmqelTDTv+gQtEGT
K2V6adtpdgRryT6x+FCcYE4Tddfq/Gwl8rzTuzExGXGxUr+5+SayWc81EvNn2kYt
fqvpLZsiF69WJ5apzI5/9nLyar7uObu8NVnfAvfQ9w1UkSNNGQaiVi/2W3Toz8qq
0nGq1idd6v5Dm5rvruGJy69yKxfQNM+PP6OaSVvfPKiju8KTmpZfseuOM7gQ0r9M
JXfPrGAi+/ISb8towtdSead3JV4RgG6tJe43XUw8elLvQa062CZvPH7WgwfSYZGL
TL1R82rBRAwf7vhQWW1+ehneCZO82mymKOqp61vRxzEtbKa1wXhsvJCGVZsWnZwR
F02SkplI69tsnKy1DKNmbnoaTtFNTvTFPJZfrl7MKPYRDWyBFtCXfrDHaVLzhbX+
/TuxZBWdlB9XCHzfoYY9T+lDXzqzbU1QoElHBbqTeYh+OVMO/eiFw+4UVe08Rys0
XNy3Y8RScPQtAMocw8uksbCyy+jHBopIVUasAfezEDegJM3LtMGAKovT6SyQ2N2p
vszdrSuHFrmWRMRSsxSKPFmN1TWxqSRO71ptqYK4Hf2fkLIjT2VsbFISESjfxk6Z
49xcUGRpGWOpJ0GZ5SglFrN0zLSeYPVKJwO23xKyp9xNO3BErbGOYE/lb6UGf7wE
Fw338Zb02yzWnGek4vKhd0y6wzl01X/0+EpmduC7XI1fAn2/Esb44gJffPrV7j8Q
2tzLEp8JC9D2YDEPuMHJWKiHTLDS1hKDDCp7TVK4VMrPJg9SLt9SztzkBR7fX+cN
b73oxtY/D6S/eFfFBghg6WiORpsjaDWvB6hDR6+g2cN8PCESbg12CGgL3Y1R+C6+
nIQlYx1ytjaPDr/Bn7GOIANUHbp740S/ey2yScGEoHZjZTfCegftkFA2mX80b8mQ
jZEcfG2oICtmddpGkX9aVVWgW2ERrEBIAqUirz61S1B+wji01ok90wbRJqU8/mCz
RlIGcc1PpE7Uj/MzzSz0BpSQmnUdyuxZRa/Sn28FHK1V9u5WF/YooLlDrirlPpBQ
lswHxLZEno/l+3AZDOwI6CKCCB0XObXVd9Lj2X8U5CkWx/QHQVsOjAscL1zg4Guz
js2HgA07etzVpM0Bs0VhbqRDVwUwJe/2Js5yqO1pwS+fLmt72No3B0KPQpyjMAtM
dqqejCQQCAkDs2PzheqXvfJiVfuJWktH1uP3U4xPGbCuA5PZCM7hV7XsSl4IIbPz
rELisjYKnschXaJSQHlvg9YZs/hxewbysc4loApry38K8dwDPaZR6PBalq9zdv5o
hXzjsbf+lEvcOl2D45O+IcWlJa1nkqO1xW8hgf9QBVa5vf8ZChIThxvAlSh4BSPY
bIAy2r5517daLkmiXvkjDaym95TmS9BVS4JEvRo91ozwdbskRxwkd2vY283xxYb3
Qowe/cHBu0RmCHxmDrkjMAdXtUOdAqrt73QUgvrKc6jITtkZuBZ8AACc0ops38St
AI7xURffgnJRMs5R3n/n0GLffcdJ9YlZVXY0qrx2Y20ZYkSzIyOl4WJYGc1UwRHg
7jRmal1IM23dPo394X4EdFIhNKLxMk+5nijBTfjHxZq8CjQJXT203uIBcpBEK3vS
vXNdhSNtb/15SwhhOhWeJQEYuL22gvYo5PvYfaauC2UvbTN+8l57iPLVJEJWzizA
O7vuXmckY3599UldDJAaKTyi1mwxLD7QDzY75suETns9D9vG1S07T1pqBH0h7ycX
eoYdl9CeCEtcC+wZML9f9LaXCgEfvNWfWr8CegoJfrRFGdoMasOqDno+ST46VlvT
0G+1/6yKiaI69PTK2zpp3Mm1ATZxsbuAzG9EzcdC+rDIoVTojb9RZL2xPgcZ/itX
BFbMwHoDBoMtkQ2t6S21TWl2iuvumUVHvqIgZEfqMCFJlXwElcQeUO+Ny+9A9Al/
JPo+NvEY0bp8cLNb5MoPvmCY8qfycCrHEAgfIprSW7LfbOP5AYTVkzNPtoOe/ORH
NzuFj49a1nuyqcdHYFtq0Tia55ad0gwRvRlGihJh93u8UzuYURj8dR3jHne3JjFo
VWhW7ovNEyDQopcfrahOhjHxxyOYAUQay38P1/m9Gfe9Gzd8PrKK+PnS7oUtc7n7
zuKVTswNDzNAQR6vLhKMvnL/rxB6tT3qb+EQXLUCQqJjsHhNXB4pRIaj3acqOW0/
pf9vpgGIWN0fzlP7uckDJqRtvBd1Vo4wQS/7LvRrL7VgolrZAk0N0P0HQx7fjHxm
Fj4gPL6bdqzdygSHtImt0ragi8OGn15NUdRAPcJRfv/+8/XxA37W8ZeUujwPecWd
c5JkudsgJ6tRRNUuFRY6EH8tpFDThubu/psi0ELBu6A=
`protect END_PROTECTED