-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
NNxGcc3o9b5EUiNN0cMrf/cHWLiV50FcAhBO16AhYl4NULmV8W7ZR49FXC96p6DD
2GFwGBz8Kk5S6TVsNcoXPM3DtWFts9t0CZQDpt0a2Kz33VnZr5wTUfnJZstY+0qt
nsOmyylXtsPigZI/0h/yYTUvoCMLRe/G3z6OEO3U9klfp/wVuo2hig==
--pragma protect end_key_block
--pragma protect digest_block
669wGBgPPj+Mkjjawl6Yho3PNgE=
--pragma protect end_digest_block
--pragma protect data_block
A30WnQ2Yg073FTmo34iAAW2gKqQXb19Xw7RATOsD0djGQNco+M2+zDxoIBQVVc5O
qiT9nwBOkrDqYzvr3k2m9Stywzh9jQ7NaUHTDmSGvbGgRxaA09Ee0Z8ntkUPpZr4
nMRNwBXS0qplpH33W5aPjWmkSW2jD1MdozKDW7cbT9te5X3F7T9Hl1J9b71x3wzx
7kVMLJyM3bQSXrO7g0o72lwYd6bR2KfaUuMBnkWeHAlBCR+RekqCx9WwZJqkmK23
WQUbWhgyXdBeOfJOYseaOekvUC5DL6m7p4v2zNbQ8ZWiG9zTdZqfNngC+rT4G30v
DNlkS/Bq1Sz9BTZYzXEzoIAQ60krH6+ijDCnNu7Xj++OUdYq5NY1WRVwn2gpl1UD
qPI0JQ4KjnIDpogfvpztRUHX3Ji4BW5wq9jsebrX0wAaFLcMVrFwIZNRilZS3KUL
2ZxqKYjYZbBamsiwxRxfDjCYMO79gcdz6C/qwlQ+ehJQdEE+RJtMqihLW0Au5GVj
AcApJVd9sbI6hqy3wR+GneOZimYJNf5cz9WW3O9p/JTm/HXvUd5A+p+Jdo1W4Nma
rduQK7bLDSa0BFUsf6FWEhTUpS0J+Hvlxz8Ry5pkzrF3VwwtZYW+goHevwUYA55N
7uoOOkvTFR4hQBMJXSpGt3e0IWu/aRtw5aMf9FalKi7Zw0AERANWYGH1OWhFFqSu
coNOsCUdIcJ+hy6Fq26ebTohQH8gJx0/V9LTnAXllkYWIoFEmdu1MhJwa+iZiQmx
u/3iOJbX3vb5SLhtXdDExXx35qvjJCQYndrFRKz/VrObOqkYNX4fdAsEUpMZ/JmG
25/srFmmJV02knb+gEH6SlaTzsuYlLDN56XmuhJUWHTdDYqwr7Z8+bKJsMQDITq9
Tiq2BxqNCslQb4NgHRPhHGYAk86gHK0PUCs7EfOQapuik1j889c+tn1hQNxEtlVJ
Sdj6vZ5TEpYtJoq/Snuc3BLNZWdjzBxxf+sCme6x/t12bdgckeR+apgpRl/HEhw2
kPrnTbNlHCbvCcjPB3W4STiuN9uWYiTEuw+QLbdaHt7fyAnkGlKHZw4dwJqNdzrA
adX12g8Tw9JJXvy7sqVslZiN9MdjPmApdX5g3xdCi6Ssj4TZhvEyZVQrvIHt4P8S
092B6hR4fY/okq7oruoTBOWstH1GXHmPNZqrbSvctMEkovuLtlIgBdqDyPDs+bMC
J6fqbcEF3hShR10//ukxrb6bTlvMriOiM20KoltoxoQg2BjBGWl0WjS1LskZIfSA
WuFTBS+Dhbk/O7dcRBYLPfIkNT1b3BkS4k9Yz0pELmZIG/AeVxbjcEmBdJEy0/ax
Jtb7pSZGvPmjgXTqOor3MiYR/5UvBMB8K0sfWIJkzvtvdDZAPHbFNVj+hq5cm0Zh
MH2Um5VJVXlOHBCS7mAh9N3k56xMjLWT9tY6CCTeEYyhhLJzdBAKf2QYUBCEwmRZ
RZ1tX7o92K7T3fGcJ+aALsbNxjq39QKaXh1B9oUmNBK9tO/5MuWljGojeN3RWg8X
fTr72eFDAiaOfVhEUmJU9gFlx3P/2g092TOxpmkKSvhznTMg9NDjeDIENVZp77cc
Z1mHNnJA3ZvE7oqDE1wuwLIPSjAywu9brSJpIuE5mTaO95d1LpStagFJsKt+UhVo
q6z6MAIjZ45hL5aYjBSJR51ZJ5tuSVRiq7IM4Ki8S7F5kCABM13NWlZgUYo+DCIw
ZYJGLz0YJX0ilJQQLKQQBJFa6pFEkQfahBUS/wiWdAztmjNcWATbYAak+N7nLCyw
2vMUqwMY+CtfIwo/GZmnkIwbPqz+tz0ioS+D6dKsWZ4KKl81Zbvwra/fAC6viNgR
mlpAmOXIRmUzTq0luvf2CfNYSlCzkgV2rS2uoucwCQiNiSWoDGToi88bCqa+tZpY
AArcR8NUMRxwDys6/recGJFR6PmtI7QxuMZVjkPc/J3txBEfDN7oNbU8tRwUZCDN
29wTZjMlD54ZX2yH70ieM9phFFGrtWJXEYt/85tEg9OqpRgRk1Ky9BO0RsUTjPNY
5o7nTvGhNBpOe/L/vkV/leWi6AFxluj5ImTjU7LkSecvNpmHunxEGG4/ixXyjeML
DyxxGQIinyj6r/LJI1tiRZ92sj5heYUZ9vV8uAyExOAdrVq97lSc0kp8IK25SL+9
errY0zH7H8eqbr/5RArDzaXSbkRgV2GkTN37njolnyJPTFejNsQawt7/UE9dtz71
yTrhfvzX29KhMitYNSMrvmeWwjQezCV/ZDN0tNqnup4mnqXUlXTR9D6omCayPULR
XZI63KKXG+vv/KOwQcbrIhDVOf++s3JitZJzJNa5fnMMvlc/PmN19O9W4xL/am/S
WUDnNMiZPUMNl4Y1EhS14YO2uMC7KXazRXf9fOuB6fMSfyAwI+HpBOFyro0/X/8l
ngzd7KWUcokRctoMMcvIKm2ww7TJygCnKTkcKvBKad/xBC+IqHFLRc1dlMnb1ih7
6QBNKGNAEiJdFQJdpr/TdiFK6QYAT6bChtKa2+B2zlL7W2+DJAuN3Qh5QSJZWccN
tno3Yp1FA3cqBwK3Av4Jg/wAA0kOyfj1ZcO4lv26D6m7yMYDrtV0vo5oLGqFur+F
dpq67uurSP+nrL2cL0OEbq6+n7+SdSy8ldWvlRX39EwiEGtyIym1KL8xbWmlF9fu
lS+K2dxv0CcrzKLxMk37pSu1IfUZSQEnzqz94vipSi8Uj3i6+CSleiRFhcdkrJ8m
GnTkXnHJGD2beOB7CN+srUT2v6wAAenyL6a33vFF7NIQ4awaXyHktaIb37UiksD8
oEmPZSMJ00QyeIH2xdEKtBcUY0Sf5q5vL01uCPBO2fTJxGYda36nDiadJi/H2PdE
7IY07FrpOYaDNqjNlwD/Gcfab1zinfvehdeaR3bkI/q0HQbcIWEjPUexqrZnjKqW
KkUxMjmHOFJZOPaIeqsjgb5xKiP1IK3jYlTIRNwpmX6cGFRBCMjk7CIEIep8xBOC
yC/bJoItJldcPtTX4WaBbZ2VYn3djLLs7LkBINx7EI0gLcqI2LxwFcYcojBs/m0W
nsosyQC1/61lg6ipHsX1a/4tSt8YJccVe4ILAPACOc6MX2tTCyOm8UVKtWqoTwLG
FED9pZXay3dihRa5YK1FU/yiqqisVQHH0E1KJcG2E8kkn4tgPuQovDzerXO3eLx0
M2s49gM3q3xACqx3iuFnkmjuLQttO7DD9Z3FtQ6/bJH5i9eXq9NwhZ6o4cX8B0cu
T/HWd7Rm+rK+Ww3XdFSd8hJANrflUZXLKeSEdzDH3gh4ewU+TgpM9a+rstEWP9Kq
BQEzn9qU2NspKTVi9mJ1JNjbCunJZjGTJuxR81/TjvC//0A5xxF6PGSJX9igZBuq
2Kx0L9DynM20cBJLc66bpKot0t73wKJg5tlWzGkwWBePh0DhbdNs8IgjqpmXHOb7
ZaW7R8C0/n0DM9EJ6i6hg6c1E/SEB9yRgENsPzJSNB0KLD0GTdnxqQXfb9zXPgoE
Qv/yil8APBo/nosZywP0pFbOZ2VsJwzsmFEN7ci52Uxg7y6C7s0+de5b9aO3EGpj
MtNFqyvzn/JMB82SuL5sAXiCkBNj6RvuP5kcG4ueZyTsQ9eAgew7KT+RtCvGtiFX
TgFCdxnO1S/ThK9j2J3fCZ0APvSv8xNZ05YXJQpDBFeNJVrrO/WCQn2C2L/gf1/q
xlAevoYH5nxWh6STgIh9lOuATh0vnJEm/+TDgGLP1yMfM19RxXIHkPP16tK5jBU4
R6pImnl4DpOLuurl4xI7YzqqUGUVdTk/XvZ/2q99srXxAfi/b7t36PSOqCCcl1VA
5hSVGGvWY3YZqLzxz2mdlOS0duqzDuQXpfHW3Fs3NMn94DMtYYZb+sZRTysOr7b1
WWPrj3XG6ckwdoz8TrNHOkqLPqqcBDg0dQAOUQQvMJ7qR1ioKtfz+vovJshN5Q0k
530PjQrelJO5W8qEW4nQdhgjpjpWsxkIhpe3+1X2Kn4YKkmhv3MSWitkNd3mOWUf
K7/ybaQYUf0aW5Mfw8RaFY1oc3l3liVwKWqmq6Uy9+jyE3MKUwzyWpm4NcFwRLcv
LkuEiAh98aa+SJaSizt7HA3e+7+KoXth3084Zo4OS79zBN2PDKlr+N9bSj7TPXFR
WyI/jteFWYpSWlq92LelM5AlPQISJAgn9E1oofxCD3c7LextzqqsEolx8slRjumK
AHG39/KTSXbntKp9X0YfgXkq5Ei3Y78Gqke/MFkhUV1dTQfAT9dty41lRkahncBm
F41tRV8S8fNwcqzgkzyXH4cpzc2QpX4Yf86kdPaxxLIgls8vKjVi65bPCcFY2Ga0
EDBDUNrBnlU7BIgVaoiKpYX/po4VsIJ01lL/D8pcmYFmYFL5SmBq0GVTVkeEg+mG
41lXLkHHcDnpR0267y3IJkY8nokUOX1xv7IXm617/KjbxDW/iOv+WsO2yrmWWqNb
q9pGGtB0HmFK1DDnbIMv30UfdI7z8XrKCo6raCtmLpl64ktO/LYrYFCeRHgXZmYT
HLqGIFb1Kkc0pVTEdiHVSMURKuc+3R8lg726202aV8vjAxaSN0XTPmGjn9qOgKhh
BR2wR7vwP0TMuIqZq8quH+BMVC8u9x0vJE+h+RhLVX2/jfbZ64TUCsXZfYdDBcFp
/b65W79vpOcukkQB2WHTkv7LL+VnNTkm3goNGV5U0HmfG1zv6zV5tH8xHgdgdXS7
a/vuu8cspTt1vIH8id615Sub4FNxaArRudf6PJF5Haxi0MFym/+RFQk2svtfpdCZ
xs9OGRH2UfJEIPB6wo6l6syQ71eAsr2f+unf8N8IR9uCdjkU1DhX1ZaIjgf2J5qI
vl/uVxCoI6oWb86/wIIFw+sc48AnfLTdfn28U+oTcPX5l561rFFMMT1f3zHAuv0Z
d2ym+dXh25Lav2luuP68C5cLj1+fbNMRO4I7JNjc1/KeBwXIUgrl67tNATXqMwE5
bNQAEQ0/zHcn4gKenDz7IW42AAEszLIIiyFRA/68BqNpWzpGEHIEgO0RIiee/L+b
VuaogT/mqEv7d7/YsFHlquE9V6nvzltvNF+3UeA81v9wMvhKOmZZJXhcrqU4XHPL
uxDmj/jjBZR/kcWtTrUoOSOjCr2WOvUIpsfJb8Q5ByBKHhqvf1DeHbO68LfCi7a6
Ow9azbBy/7p2JhpA9s+LwO2yCHFmNj5ZTPZpOp8XRyQHwUnsUEHi3+FCGCSyUDzY
6MHmL83e04zjOkZcFbHHIQ53c6+MJ9JcHlpp0Pb3dJkbWN9lbo8Zf65yf1b9qTbI
wX0fEswQUuizadgYkT+x/sLiINcDTVvMD/GQ8y224Xn5+dDaJHO2Z/KWHqmM4Bn6
a5gvVs7bTk40O4cc0ZuV6MZOwKADWsJXvpC4oh9tTAOfQptUIKoC9B6JpQBoKocf
/uBy55MqZHtuzODlUYOChGYpnebk9ITwmiAU0XvNHmSOOzh9yGcNRqhRiu/jvKva
V/CGZGP7OgMoiOWXUR7ZJMHzxSSmxsL7KNhKkaivYzgIiQHzzLl21Ztiwikqi8ZI
MWZGgVUdIx6SdOogC2kGelmCz22HePM6YrF/UkPomZ+U/CmaS1sr6PzTN29/SsF9
HDmiSkmYcMtkzo/u9cFyj/6zBBLMO+KMfwB4ev60TN6dSZaCOaF+Xjr9ZujTH11e
25wgzUwzVO7zCKQCEsxO1JOfyYYFKUF8k4zAvJn5c8yoIixgFAXRtoNWYF6FS9wQ
Z202sJp8FBoqPtQeSckLLLlwIysgWbUDxbMfkmGpcb9dC9xuatjs3yhxQbX63Ill
+kOkpEj0TzZVLjFggQlAMCyQR5/WXTsRGy5ZCwb9Hv19MxlR40UUCulCq/QoLC4F
G+P8dWcijex/+ncjceAxa5J90lFCiGfago6vfWZE3V+Sp0+glhrr17HGLBkz9xRa
aXopXl7qVY78tM7I2GIfs9TKQCh+SuKcskqk8Qspapur0L5zQa+SH1C0UVQYZ1ps
44Bj1eRcO7alDkNYDLln7+cUztNp4QJ27h7tT65XUaCt1iw0ZrvQZrcNAHap6wLk
PyXyLVew/NtSW8iNESVZDy4Lky3RgGlNiK49YvcP85/fn/IiBKIfPmxLsR+b273r
bg27cY0g9R7EVmLcr/jSw61DX+NAbGTPrZujm2Cg4e7n1gfrKztXXRDvai21ZVjc
FxhTOmgjCJrT/JdSdrSrx5zt+rR5Z4B4w7Icn5FI6AIcfCVxrKQ1Ijx88AWG+R3/
KMcBqKXXPnAYywOH6rGsXuvzwv7B/ZxVgAZX0thaimVSiiIyKl5l2skWdwOxu/V8
4cp8Zl3+86CtqcSrjzo3RYBDIkgNBY5r+d4yIMZvG6yU8/+T0JwmeXq8RE2HO9Sr
5gVA/8asT7/eAGu9GsU3n8NbKkiDY971s6dG6GUgTKXFwvYbZpkyv1B8VO/wNg1j
1qgl6QDb1cZ2HIDuUEZ0I0CauTtXLJNhs4aQAm3eLid/lkLoinTC3+ffAuKQt97x
RqAFEbWrqARR/0wJ8BRX3PidJGvcKhDPm/Ixf2zlhRY14KENvtXbcCsiZBjxDZ3w
U4bidG6ADZrBngm1C+ckvUjuitQBJ4RaHoApZ/nwqX1pbH4FLnQnkWP5nYe+I1kY
Ty5aXeKN9dRHNdDPmKkCgfEsfBpcZ7pyZ3Bjjqq99YpHeTogV+QF3FPXIe8D+qW1
Mi90BKfw7UUO0+H9Vuljb33CiwsOLOqBeJ1BsZDP7pOP868c8zeqFb2tIycUriSo
y9jgk/48zvBSE0wzkXh2FY+YckgT3aBooE2xWLlpa4OD2gTEH9C7JvVjqhgGskFD
CjmVEufitFl7C5HD/T4eVmi6MafVllLU5osahLRO0PpOHTea9C2AKdybps/i5pa3
roBcLYOVyb/FrmniyiC8jU3UTpr+QW4Gxn0oluy5N/KjHeVZnrDNvdUKGq0VjSWz
0Xjy4MeCjdzXndTDPVewLYw0WgungcfaL2OhV6KEf+eq9zDpzY2l/kBjrJTvXzey
holV5eeDaPriOZ3cwh/hT9Ve9/fO/cydy+mqo6v8ap1HT5Ei+ZDheIR8/tQh/7Bf
WvSWJuCvIQi5uTQC71K5CgmiUtnbXmKNbxY3zz+nnsj6XDtFjTGpQkKlYiVSEbI2
ATWJyD/QOQcCz9AQHNv6G5sjehkGy2IPJljGgCPDWuz88VeTsn9ZQ7hP+eTd4zSH
V2GikHVBJ2OIQtcQ7EaxvCzZTXN7yJ54nXYPD/QfbfVvLzJXxQ4TKtphAIcHdXjf
OVPXfctwKyc6ZhymmA8V2jWoC5VMzODPpAqZNTPYhJbYrLRTfuGC/75LsBrylIhA
h2Q3q54sln7qwEDfcix07+KD9auw9zqHejBajYv709QjmEYe7ocRb2jfPnRFvVfC
86TarLXHRXYQJOFcnRtbO87daA9m+ktBpUaaRNlKMc7/KU/bnGv7utjK3gNTPphz
2mY31ZLH2qM5kRPd2HQe5uygfOugoYU7lcD4kAd3+930H4x1PtaSJd9JXch0Ug6L
utO/CXYfBUj9QlXcgCLbBx9ToIFkhDVrhFCDQLAM+hUMCrkQMu2p0O9YU5QTFZva
x1HPC/4w7LFRYjHGimAJ6yXUL/HtAKQLfpUSgraiIWrJS3WyAT8KDnKY5oQcJf72
BO4eIF7V86XSg2jlGfsYSXAtw1tGuPwKr5kfgRmW+HT91gccOe4x9uuWWXl9fQGr
7AXZtGVLEzRCDCO/mYcq9Lv+lxUn5L/+CS4Ox7RgesMAH07gXSDskU+Zb6VT8GeW
POUOB4wakTk+CLFnP8OsUUvxWu2xaLtqOqXY/g2zA2rtPrAmSVOcACM3FnhTn21G
sw3oeN+BsDPsDSB18ZGk1VVpJM1dMJWj8x/XWbyiF5vfjsx3XSMu1PjJefzsKdv0
IKP6UJNrONa6fkwh/z30H10nOU5oeyR+dmgZyUXZeqGkKVqNAkZVnXQsXcPBuG4O
akLKQ/uOSmYcGYwzyWN9XNWpgZZ49E3MXDGHKgZ6DToUPxEYcv4ff2YR9HsY+q8B
hlpXp4oAsr7i3aNoN2wB7a0hVSJgdesRlk+lT87Y2x9J+QTpnFkyA+7jFfgqnkAy
pTIWpt6ygChV2ng0RlJ4UtIYvq3M+iFsfflpUkG33cV6hQyNBY773eK9OUgxB9+a
HSgJFlR9UjbjuJGoh9de2jJHiuKQE+zMI7bpf99zQLgXF7F2Y2byMpcoOrbWnDy+
Pt3ta5gpcQZ7bK8kicm1c46y0BS85rCjxV279iXaClalCS6K3yJUaTMxQEoF6PUr
hkkyMuXNPIx0BKwuFhqHZNOe+rZq3T3vK0XP7LYX2fjC/3fbIlKsrINzCFJmzfFa
nYGtTg5P4zM24NTCcXUYBe+OsnmAlTeFsocXnNc1m6wREmlMaAQDkO7kYNIm9PRF
Ecs1TsY9OeGnQS3lZMl7cgPrDB2dWSDW6ewVlmhW3BbQSTxllQsMG/K+YvD7qJTy
5dkWVwHKH1daILxcLY5FceR4Z1HXWYmgxSxE8tj1TXQtd9fMX52YZvJL9ISS4ycw
MxFxV66ivedRDQgvJ6nJlZQ2pru6PEJpEvocpjc0eYMVM67/oHn9vsHKHEGc8Al4
HwGaqlgowkT4b2W58oalUBaHQGsiliFLt2ItwjbPh1/TOHcYqgPIGvUZTChIi7PJ
X35gLDgGXEpyjgRUYHgkPEqXobiXCuo3CnglyynoTeOEAC/KAlwpcGiGdDUqLJOU
GOocFQ0DchkBsmqpaQcnxvLIVHQhnWF10rf3Dndl/qWSG/Lvc1iaMkZG5yRWU6GA
Fwpn9Q2TUKw/bCpQZAF+cUNYNUopdDaUsUf0X44v8C2wCGrGJXpWdvb4Hegbr1GX
6dRPhbX6qlMK+23bGsz/BVQbtJ0gt2Z8BJALMsZ1g6qNdkuQW/HV/eivtw91KA+a
hHlrzN8HDEr+0Ysms3XujC/sdRRao6Md0FAsLmSos67JnaM/JW85StL6iUkz05ec
dYeqj6NFpgBaEY4UPSwyo78B+J+ANOMAzPNFUVx9DYyuxDql7jfUajcGykcxYPVv
hCnp9tF3ZLvOIPU20AWzsA34R9Mmv7rG4vpPjTGCUzIL1ento5tqtQC4Fkqrd94f
N3VaTpqRiVYKjWAWlRwzI7a+FpquzyZ74zTalj+XFCQwH71J3QSix+K/SfwUVRN2
cj4Cq7kVjEDlfT87wPH/B7fib/8IyBYbFis9c1O/SL80Rn7JV23QE1izS1XZBKlx
hEAO3CKIaUdQ04QBF7+1060FAduBdEULy13Pk9pmRNvsaabunlnvgonFWF2yBNCq
7pUw6YD0yM0QlhQlysc8uEDkgsXd9l/3GA63ttg8z9VAdP/QbV0b0YTHZg4wiNY0
Q41dE5lShLauHz7YRETa5oeK3MC+wsJiP5j5w9s7XQbduWYsJYoABr0f5wcNF0Eq
U3CjOmMQeuSU4TQ8oDLJrXudAum7gW75rqP3gtXtxh0O/pAfm3Q55YkKquI1udE+
tE4CxN81r+QeLIJUjPz3737g3J8b/dtavzOZYp0zp7SfvkVe0D0RIZpU9lghLZLD
0omJ0879ktwjb6ewJpJgwwnhhFPwGBjs6Nq32Mi92T0dRAdYcouDX5a/djg3VR9U
pMpLZ+DV94/HRa1wzvDUHXQbT+WOV6Ge+a4EfM8nQgrX2KUZxcc6TVYet94/Utbm
BI3U38TxhpfanrokK8XEKXdRsF0LtMexvXruyddmpgFa0XQ9w4M44AKtVI9j75eO
VaPELJ0RRKbzPbaGS6THZXuYCj7ZieWXUJLflAzsZCLyHWxJ2uXCqvc5IwzuefV9
WBzI/phl5jksDOMsyGYnIpztqp1TL+IgvsR5H4kNDou28j1mu3rDNt013SDYOyj3
zkKxx5Tvy/HJ6Z6phm9cE+X02EL5O2Dg8+5pV5A+KYJFfHlCvJbUdgPw17l3MfFI
Ghyu93vZu8K5c4VYY4QcM2PEoH3xHMr//Z5MRggDkNOveqSSlwtsf5OLsJ+VWHyT
p+/kwkOImN52syvOPz17EX+JimAB1j8m8fB/RQGJB58d2TvQGt9zgOHdhNpMHtRW
x15J1iH6ExJOJpyfhaRRQ7d9zvgUA4BORd+q1P585ZNqbOyvDD93JQ5h1x/YmJlP
GQ5Q0F+SeVc/RALI11ksuAkuWsYmf9J6gJege9w2IH0h1FpTReN/yy6e+Sj73uX0
8dfjAPNuMdHldsiWQJEt+atLIqGbOCQlDAaVEClyCjATuNqZxzS8dgGC8MReU4ka
UTGzSDwyCoeGShd264Pr9D7isuYUyr13RhFm4zbOsUbfEbgkbo/jcQ/rm2A3sVQ6
myjOdlDIl8GjgOWoer9ttW+RlRrDGPvLzpff7pd4Ff31gnNHteruAXo3LboFTnF/
UBUMYTx7cSQXds1SbtaUgjgbVA6HJgngetzjClEvtoTWyonWRTBGdxWsXLvvSwJc
e8x5ASz/+aWbCjstt+ZHKwaZbpC4fTrktwGe0VCgaqUypwC5359pjiZlZ9qo5TMb
vSWiyEFguWpEumgqV6yWoHr+3xYx9kW9A4tK363EDwZT2Usq3FUWfzbJ41Evz6P0
8yFsmfTBustiEV5LfqzKTxVbqZPN0+KmccVrB5yOunMyy7hsehFVflgrJ8JVy2B0
lwZwyUiyVWh2PHqW84c6EYwMxaTKva5gy9Wk0jvqTDf9Ck65K/GpIVMfxFLBGjgr
v2/HVTAHEddcodtxtaI/b7KqSj53RmoZbGLWQDZ/xvVBlswEK7PJkt+xaovccAaw
G6jsxFXaM+YEm1DJKnacbWyx0/iSfh+NoIJA7Kj8e7T5cuVzxnJwm7+zSrRSnpih
bRdh/iFhh4Utmy9J5lpu1HxNf4CXb2+Bfp8FhJR6OW/efleu9x6ag0c6avNS2wTu
W/tCx/w1o16BqqnJNrAQIG3ambB8n5Ib1m4RQRDxXUe0wmcpYFCzcQ0JyF3bdYzj
IFwEQ7bvABqyZAWe6KtPoAik4MwSM5SMKDx1ybmxBx8+96XmcQWm+8rBtbPOd84A
ExKMbidfgjY+N0g+kiy8rIhaZ7TkghIJc/SGegnvLi5MNrxv33hQn7ynbz6o2I49
D7qDMarc1OPZn2Gu1kIBkY7/LBo6f0cy4mcHS4b7RfjCcVsJPr4Q2AJOCRTNjSlM
LTmHvLjSx73tRFgLvypjccdDIcgUi8EbIcahvyWA6YjBLJ5z1MuJihXWr2FhOTSq
4ZBld0n9tBjTHqUUkUoHPOM+J3YxrWVH59Zpgjoa2Ix3ABxx/O2MqVOqrKMlfPO9
Kxb/iljqnGLsD4BKsR4snG4aQIbvMn1nolQo8Mw8nI9NLPe8hnUOS2KOoIK6wpJu
z3Evhyi5if1pVb6AZqMyDQ5m5w2b446oZiMLvdx3Ap2dMpfK3+X3j4Zhj1NiurAB
nCJDmkQSyh7GcYVWLe3MrkNva0aC+Bat7noWHyGdksfpaT1jjNOaLd+GqlYaQMHY
Ir34PaXcudfSG5mxciN+oHvRahcgjCRzcpNwRYx0Dv+A7HqW020V7zpt9OviB5ba
UXg4qMh7hlC1/mJNca8pk6zgTtmxVz8vX6bKkWqzKt+kdBtNH7qzBD0zFzKhphFf
Rw0yjWRJpZx80+NHg81DR6ZA9pNtOim+zMM565mPW9ORnr43EZA4MQQKa2v9CKGa
R5KcaLBKmm6TQ6PFUTh555663eQ+vQ19nrjtQmIBFMI7HWMiCr06uj8HXS2JkRmW
r54mNnJZ+QcP5wbe+RMZHh0yTisfYu0rCsTUTrNot2/LvTlTxZQuurkDgd7BMU32
dB0W0QJCnHLULraY4v1P/aHYWELwY2IK/sO4tSxc1mHnNajKm885u0K7TfOBM3Ga
H/ehHXvJL9B+exWvaHdvefoEn5sNwsiqikr+EkrXIBYdCDvHdow+Gg9odw4gdWkn
MlwwE4zJTzwzrtNSKP02WIANmvecC2zm87TUZxB5v72DmYAhFCU79jjyuMeuND1p
K2CjtV5uAun4FZ3wfmRM+idUVJFnBdst0we/oukfffk9b6JuRQqZwASVbLdi5CJm
1S6EvRkTPiJxsKPUp+eQbijDEBuAyV0TMWzjW8ISJuY46TVqM6Cs5k0/culSowUQ
75b+OcMVSlGipQD+vG6kN53/gKjpr/Sooy+zdxWSO01j7RdOBZSTooCfp8NfJpN+
bMwd9VGu9WaGbAU43TOW5S3BAeaLVty/zJatM613Kk2pJPIMakn8Fh4HXxjJPwPM
K/Ax59sLrdMq1muLVBY1L5w8nXKhyqkyTxbrfPC812iwYm+6ms5DY8Ci8MZsY7m2
5ptW5ygnjgCPAFvuu6p1MTHA0imkXuCG7+eVJC3uBkq9Gh4QVcHXx1NWGBRXmTvW
wxRgsg3+6Ud3uWwAzULx52Lqu0+0kZfRwLVvCXKW4JM+Oky5PbhJ+Cpbzsi4ON9a
KgJjQsuQvaZg2byToHPJMDhHyDKrZGyWjiss6I5rDMv522g/EtaKHxkzlmDIH0MB
aW78oGfisXdvV474MJaPz7MnZcYLhWFQn99pcawtIBWlhtL/F4q1PaBk5teJBTro
C4iZs7pBdzjjzc5Z87jR7xJagJIKwQRAx7EK0nj0rgQfjQR12nH9mx/riYz3MOiN
8ekHlyasOHbxDW7P7RALVTfX8oFYRBRWfJp7/eAh9phFTrAEKGEVTcqUYUZRsVVp
ZruqcHeN1s2izFtEcW3CeFAEZkw/LX5omqsilFsFU8+bDRklN/qg609zrqSvueMT
5yxhRX1VPgfIsYl4drcrhXr2FyWaPQ4glIeN+GTBB5QpwqXOnp0r8RKkZaQs2Rpb
evVoFgV+mWA0SJXIKlYpU6PwzXnosukGiTlpD1bh8qP9el5j9t/kJg8dfB6NMf/M
aNWqjMar3Rq8taZB+LOXyohiWsttdoRqRXZAGvjnqjGU91hXYXa5Os7h5/d/rd3B
aD98woFHoP4jBKjihp6sFvLaF7A5g8HgU4QnJtAWXDMaQmvDLflvh61DJxrneBHs
edpELpLXlxYN5xueXLIkGAGT/D6MiPCvHMu8TJnU+NiH75UtR16W18D6uBSUlO+m
JwEIAh65r2kS3Z32P9aOjMY3/DyGqXPdpeQIW7rDjoilzLd7L6DnRshih3E4zFy8
wykYOJtAlE6VFbmDup313GHjZwQTHXX5qTzx23I+YeTpVBkb7zje1DyftH84u6jP
W3tnumz9MmC4suwskS7yRNxlSeTzcve5IUF90b52t1f13AklClJfXto9RDhx6Ydr
N5cs/7dWdUQMf4REMUskdCu1m1Eatwrx008avWaMvCHHqa1UOYffuNEzUJZ/Dpot
LUilMryCHp985Gy+xVSYyMMYSWpT2M/mKxdG2fW16V7IC0E0BfH3IfoeMBcI/8WQ
+aZLiWDwCRIQAmesaUDooGMU6aUuHo6MjIouH+i+feSvcNW7cOckyMF972gJ7Tim
bPp5niUiuyfhjHg2JXaAYmCO9RSC4/3wQZOZszdmfJCt6rgAPVMEhAgeBm9ubngW
X1NxxkJHGHRG+2h2qtq8yACgiwrfGb1suOHp1pCrv7QQHggqv2pqiN6rjLtrubEO
8JuQ8hm9jN9ZD4NXzVGvrQS+iC+Zoq8WYpy2CVFjBJYlnFUjOKilhz0OMHB6d9HP
1zfwU/weDfhMyq+U8UGQ+A9KGihbJbihGT2mnoW9E247UecenMhmC0XIbPdV5yif
7PrUE1e6E+3QTGGC9QY/n2cw+3QDU786vfe5k15RSEs3F9mwMimzAyRL+tYUEBw8
dEalTG3wZPwmtAWz1g2aPiOn/4F2RoCnl75pJUWjzQsmVsForwNgDSJPJjGNOT1y
UBNKGNURVRfLN5m+RPcNWq6ogPAnmxTO8WI+BWTrzdCcxwEsq4urjAQ/K6mJjiMY
qLuUIeo2mHg7VVcwLKb1dUb4yCUTiog27qMBdt6sJGZENpk1rhEt+0cZsR99USKC
1+enQ/UfSn7H031JwnLMtq3oTc27mHAj32SGpjrGQCT3kwdBcAvw/7/VeKgP4zkC
lFUeBXH50II9dZnwSsL2pOVByuQW+O2tMuneu5tmoscZf8AZCcwNApYYcK1shT5M
MmVMHlYX7OaManvCMyO2uXOw8zLf/GphgcFNDHfRBZrMMhXGmkCOeFSL0jpvdE4m
XJFbURBWClRyFFex3KOFjPCHWjlpgJRs6mjAZYDXI0jeUJyhxmRmVh8+7+UUVBLG
Y2EtAiMjYaiV0MKVWTjX8cgJ2eFdZvpm9TxViMHiCpyP7gkSV75rbdNJLjb/Misn
mmGhX6N1Yah80p15n5mF4t4KER3FNE7oL2yXK01HhZQJB8rgkFwpc/dE51a2WoGd
Tc2m78RiaWtxyKIk80aQiVRCpkaOq3o4G9yvRR+Ox7mFRAu9uSgDYqya4nROb+Ni
qU0Xby/QbqpBKKMVWwseJz15U3U6Ev0I2ZA+6mM70B7KRgCghrvBYD5rYEn+COUU
dgqz+9pdeXIixRzmT4IK3o0qz+zUfWhzR0SG6NdTIFctI4q0T3YGgBV8IO4fkHFK
/ictiWCAJlRM8JMcv1nk0CODQQW5Y6iRchkHKFTxXEAmZHTDlq9lvVPBB43HA0VG
IwIF/6YR2E3GVqzCC3ZtE8VUDnHfkjYW/shcB64X2O69jhsqYPagzW21WLQlZ998
ZDolYN8eF9n+bI/kspB0N1Zl6OM5Itedkuep82F7H7hHiVnrnajecT1jtSzyFHeL
vpM5X7CVmBaEojJ1OBlD1gbal6iBY7uUENZvPCHPPu9x/hSUpDi+argioXx3AGU0
WDmpE4rc4QiVrX5B/7CFdRLiAUj8310YgiicZQx+odksgeKQIFfKUiFbxe1HEp4k
bze4Md6IYrwpwMtXJjIqhlyzj+wdOL9If5pfrOKDzIdGgWmFnkGrBxWoIqlvQ0yE
uZd4hVXQi97gSxs/cJepptKYCaBWvuryXXODuB/PK6ESXvFjuY42OZtin0Kr5Ze2
Siin0XApBKfsnzpqg8ZmYdtEzDt7XI72aRz5M4xJq1AMwqO2GyOGdjCugB+tV4ke
3/vcf5KbKgIu1sJz8yclXhScK2pSHbG7rW4cV9dDRQ1VdSRU4ulwd2hfBBWEyoJu
ECRk/z/cJNu5Je8KMukxhokB8TwRrC3zJHQ7dT6M0kx9CH6XqEy7kkVrhj8TOHNH
2w5fe8V1vebKMPM9Rn4oxy2h3f4wahjjwleb6TBFfZvku7BrWcLgndVnLFhkJPeq
R6sH0v7z6ysZZPZ2UZz9+GSB8HqTsf9MbGjKqc2m3pX32DQtE58BJ+RzROOwA+4D
I4EMpdY6lCQbq7TJMr0O7Kn4hsGK3jXSExc4rjVBo2kS2fOgkhzDVXNrFAcCOB/2
faV9UWsCycNHD39u8bbJtJ59yr5+vK7vpucUJTIBg/63m0dkM0wOc5jbC7oyiFQ/
NYyON4MtncOInPljh80ipvd1z0TyEbfMF1diOKddTZmM1AWw+XWcWNHAn39F6CAh
2y5bMObqOkN0pfGxHRuY1nH2UUjzhhhEua1Z9dYL94PPg7q1c9lzpLV0HjzhZMDH
O3mb18jZLclVabIzBtEOuyyMCtZjrdRqBPbGt67IW9KzgRUKdPTSjtGwW6z1/Q75
atPcrKYiO28ZOksnC6pNfCINRHT9252pthIV7WCXCgDTG9Utb5GNw82dw5UPY/IM
T7oTpcgbjER/Pb5EW9RNdrFsi8bclr0RTRdu8amNyC84IxBnRuqv+XkfirJ2qjtX
38QLyHUiyBq+k2TsHY0YbysW53ykB648vzrO18RONRMdZsTZ5imSsA17NAJCWEV4
39VRxgvosBxquLoZIy9loJ0YrBmS+LQhk5XMrtIT+xXUDTiof+9cm7lAZwetYO/F
mi/GHIQZ2qBYnBjufIwucGEXSkzJcj37ZQPZD2fCPpd4OEc51h3OXP+cXXBQkMGa
sKmVxeJaBkHyAIL+dEu++1wzvT9IEJNle9vO3J8PAeM56BifqfxZj7TVqS6QhXBE
wuZM1O0pvCb0X68rKpUAhckRXr0qmHLU4Qa2XQ9He4aUv4QkfNGfpQJ67VfkD0Xq
J5DEKXsTR2JN5rRmRxZC21C3ce5CKVLS7QjVAGI2vnsvfRDnNLhm8UeLBMRqRY8t
A664k0OmovrVDAGwmpSOlaJTq8ZJLCBlItL5lK86yb2DT13OQpND9mVL2qTvdxuT
BH8uvM8qjxOJVYPQ8GXv7nuvawLrqfuexgSAgf17QsROBy318+q5DilAPd/ig8Ov
csHEhTJ0/XuLhAIjqInPigDhC9dpLlD1rw3NdlKzgNBEhan4o85wES37MAgBo4/o
SFhnCd1WBcnFiXU0AznLHXfhYXQuhEaCR5NlyYQ92MlQmLHFcB9h5Bo4eu7I2FU5
/Nhq6i17V6WIEtc+p6wd9dKfPapD8D0IvwiqZbGviGr2C/UUefexRNnbq7l7TMWj
Kbe5CJc45GskeYtaNSI8AYVy/VQAKumtNhzihWzGXDV2GKpcKipDw0ej4nJzmrVV
mqveAGplqUIF0Yx8L06xIkWUREZW/5Ln8sRb+M5b5S4Vd+Co94AffrBjF88M+jYS
Xlx31b/iSRRBxo2OnNOuPJH7bysfnSEbAUFJdc4/ZGn9OEbd8G5VDw29CHmCRz+q
qaAQF+nl5mcTbeXgSAhymHaLMqWICc20O1Vt5D2ccLcYf8pa+z2AqTm8b0fQupxL
KVK3NTt0WP3/Ln7oQwpsb8D4DeaVZbHvlsFDvYX4RhAcbT5NdKtUfRoWxTGYcT8v
6gmuDHn8ZnddXZjftf6hz9TEvARqj1sbsD4UWTFb7qc6WFAM7QqfHjOXgatWhPhe
xwS1oqN6KBHNh0kuTB/YNHp3XdpgfZ/n00YAMHjmvbK1/hfAqOfb9OenJKJk1WkT
PHczN0JCCdSi0j2vvOjRUS2bfK9gDcZ3WAnvrM1DyBI+rLfOUxvA9nLMR2G3Xzhj
vAxYR2UiPeIiN46kS+51t3WFqVOsGefbqEl0UvyVYcBYv4wqsFhjK/GliLNYPym3
kfemx91PwvKu6M/DOszhNU0qzO6ckzkMRLpebCD3VRETrKLuqq7RfoMWBe8+Ms2A
J1gYmuyM8vXLT/z0cdMsvRa/vXTN42K2DXxR4LbrY4kCarZ1+8DsSP6RBBB4QviP
eYedG1VyNFV5GnjaFN0+xi/+LsRgrUNKEi5A4uQxSgVzbWNPni3asYiyeUDTNGwD
TmhWgbM8meGxcHnrJ1GveldTeclXzEFHHg3LPpDm+Y2A+oHpbkyUiUQk09HE+m0B
UrBdbQ+FjDxOu44JsNjLYFtyfCEqJUBiO69IBOZ+NPWasVedjGDVywXMZeVZPhUw
rxXUai427SkeOA7tkPRcVjVZ1fnEnaSO0FUrkQ7M4b85MqRObAP/1cg+0jGgFevW
eMPwmPkIHNiiCxr3e1m+8vTqE3a0IqOX9lVLPI34WBqsrsZDB7VgabZHCiDmwFHJ
4TimQbs5CO60xgdr1rxgmw/yiFE+MvOPQFh+uX9HrqnZVXomw8fj9XLlvZDgEe9w
jXNg6uF5jv3P7RtBMnDer0asqtJdqZGQ06m/3NKOFKmXcCNFn6WNtbI6FpPXx8UX
B6L0/z9ILvFoa/MYkY/xsbvGkLFOipM53jbklweSfpCVqu1nkUtrXvPH6g5i8SQz
GAj9PQhC7Yjr1kv6IGhQxnyVrhiZ+nWwiRYnsSrYthJL5rkneHWqXcf2iVvBUlMZ
6DmmH1Ep0Myxr7vOHAayAiV+r2h5xfUzO4UKfcufKEA4KyQAy2wqeF8C1aSmanj2
LLowhAXg9SyQ49Hxcrz+Fm0ViLzACvwnyKZmjCyWBNSYD2k8pk5sVYsDIoZAA5N/
7LEH6mNz752IKz19saHhM4aQUBHrMzLrxVuJ4aS5Ze1cNN632/N/L+3xFN3nl35i
hwQNCHfigEqkB1HRyKXGjurbVkmhsIz4LExN2hn7zwRgwRamwrmvLb4Ti4X8p2GU
gGYEZeI1HSzMWs8Dl+UcRZq1VqPfc0BahveiODzCstc30KPDsRUAX/U9qdrlMLzX
YdL4W7X6EyqEcvdN9LiiyqOjALKZjIOeuVP8vQQ39x1xKfgw5n7kCVUlYzvn2GcI
ZQiq51FJHbXm/RUkYl19XT6FYD1uSScAPXt1oRQc1xPx2NotHC9aTvdAtyG+8D/e
68VmGY3ToAP8am8j5ndmFTAD4ZIHCdZ7CZai2+r3DxX2c9e2m1VwYCTYTlUGLTvt
G6qjvAuVmp8NqSepQpYIL7q13/Lu/fSU7vHTkArPwriTDhupmhK6PXZww267cuy2
HHrz+oDQH9zFbbtftw6SLFAhrYIfNiMHHtCPSoX+2kib8PLTZK2bZ6SQTGnCBnrt
VljWF6rpVQZCRnmTi9+5l7fERYleRCK1Lzp9o4y7DiXesuPgVHg6dKuCEla9cj8g
66U53dNLzUVxdJyC0bMgsOdkuc7dkmIF6+uqsNljodgYJt+QUQW3gOUz42eU6Orx
st05DVF1YxCbRwUvi46WkVXDi8O4ZeIZ/n4Hsxb58mqX7CQmOA5LHQ8K+4yryTxs
iMWRvOz0ZMn5q6Vj5G8uQsbWGU86yWV9SV/ufUongORyRC0nChYToeWEQU8zjh/U
ue6giqTXFUw6+RcL51HUGmj0SwcNBZTpkzFu9vNyZbSwDjBxHhAWkSTCmSsiaNIy
4nw9xe7SaNhaoiADTaKmWIg2yxu4M/k2CLsAxQ8p6f42dNmp9iCdEL2365YED4yN
Cw1M5RrK0zHDLypCOXWfXmmqHHWgA0wTIe+EDymcwQPq2hnXFIpCi2StdW8sGbI3
q3xR8NgJFtdkM3LUo9w9gz9AUKy6FdcqCj9LPuMRMjj6W0Lq/TlPfVwWv5TnL8W7
N8lcCIQKb48k1Zyu93aGiosXtQSCcUfEaqEnR+8eVOduy/noR0WMgWAVDkzLJY00
1zmE3EL6NHGs6jUZfgra9q/Nbu5i2j+jbS+/DL8KDFaPv0Gj59SONWO/5AeGs0X/
tHvL/U3Sk37TubGZuc5zh543+M9Fa1x9yjefypwcDWB5ICyrlHJRjWiLTJ5cUTnB
dVc9JE7GRXGY4xWEZYI7urINXu8mELeSZOpa2YCFLZqqkUQs/Y0CPgdWIrYX0Z0V
WaYYu4s4Q4g5zw5jY6lNv1to6xuovr/psAAKve7pGCgxlaH0W3RkO2LnySkPvNIG
RVelFZ23KD36APxqhKHREuxFLp2FP7ghE1Ln/+WSdw+7SFyxcjaXp+za1fwBqebQ
UXVtmu5Koeoxbd56/LaLPd3CRm6u2Wqykpt6UgD/EzrtqKT9UAipkBdUO+on3s+6
h7x+MjrSWQlA0iKhYXOax+7aBRDxtEr4RxL1hEVbv5Sispgc8Y65vNNYDqaRXZyA
lufEbS53ZN+FNMPi5YJQWt1TJX0dzB13a2Zu7OrotsEaC7R+JYUcEAdm/p8q2wgI
QAIsFnvkvyLgCozQOK3Iu4U7vGWlPCxyWwEXdjJGlrrxRe0BzvtmESQxh/8ubrvD
zdbe8p4JjHVxebYJN3P0SyAdqoPwEPoHh7lQvLyJkMzJQooWPoEbXPnfMUepF037
LoKB8R6E1duwh5wrrANkdn+FhHTOphyR67DUdC2wYEFMXTDpaPJ/t7+wuAq+cQWT
TCMuI1Th4wl8eiuG7wXUxQuwpqV1o6b9XCTFZFS/K9dQ3DgXRlTwwbQsmAq2xYUv
mF/m3jFb+W6PDkMKEkM8oWr420ZoamlhLTeCZCAMHTO2IObKFnPo6zTWuxzj9dW4
zgYsJ7nU7zHKlkKVcd/BTvOQ6SGH4fO9bwnAhjgSOsPV+xhFPlF9rOKgv5jtsWep
g3elvwjZQkOeqVoHZ70+nJPCetEY5VMJfp03QQsN4nzbugZ5rU51f/cYfikvMLll
oYXhnqL1mZWPG9Y0yLuvOs86pnEkjMJtZU8vBmUL4BBR2GTSW53G3LAfCG1wSA7G
WYLz3odPdR5UR3ddWPK4TRpLcrzpRZohRyFa+1AXD/L8Yc2D2fenCp5SrUNbE3Rj
KoWZzf2mJpYV4JeMY6Fm++bUXCOd4gncM7UyfgCpYk0ObRwMgHYvWh/kwMB9LCNY
f49Fa0QTBr/jDUX7HSd0BfjFnIG6ZUefd9Wh5+ZXuu4UeIeIZatW2I9+dsQth5Pc
e3WcG98Z7Z1wpjLQK8iRQXb0Uy/pIj0UDSPuydCzkdBnRSjgvX30qcf8Ix34s2DI
A9ptJLUIDmRlg04CI2oXd0EENb/H8Kip+inX5JGVkw6L9FGYwRiWT9XttYG8H/6+
hXpTjEs0NFDH6V/bHnHjdlSZ1c3sG/xuh4xcqf1C5sBHkLc3a+bf1tAAm9PEISDe
w+IvvpB6GcaHcS7fJNs0ZmzAkx9fZMOs2X0E7qba0FInAenbCMLAKSkwTSCIoxo3
GnwDa0BmZXJjE06mEthDsxLurvYIs5VnrslTJNcynB/q3EfqOT7dc6cb5nkRX9XY
uYOy8oiVHTM9mxrgi7s5M34TfWTVB5ktOVSr/vZojcrn+13xyajM+svI7p0ky5IP
KbeQzleP4iZtH2vp4hKDHfdMg9A77lzzGIiTnixap7qzkR2a3/S6afibAjCQxzWq
dqzSr24ZUwnrWAQfNaygOVSYJJRzhoS5bmuuU4jo++jfo5kkcp4lBp/aGfRabtET
kNaW0dDpV+qrEtl8dx0wBfDvHR7jeQ2P5jx53dQjIisP5kar48k3RINH2vBlruPs
cu4MPdH6PpNbO5C3xwnzpK4HQVL+emNcb437nZvZaN7e95rVIXLxmrsUpzNDJ6lK
tOHf6tNZjxc6LAZGD6N9Zf2kFHwkc0A31v+4oVuDPgRhikwcK4znGhRRxwU/S9Hr
rIw/C6WxwFZUhtr2mehZVbV5MCs8ewnzXkNdQC+EXTenxh8XYvIJ/lIAqDzMO58E
sb8kahaOl/djGfEyZMeI1HHc4aFTqRMk06I4yf0xQIVRxeGXggfXBm82WT4bTQOb
VPPSZ+9qhBVB/0zYuJvp4LRMB0k0pJQ+rSuY8s0/RHTTz18/y3gcI/m1v+JpmK6D
t5Ik0Oacq2D1rG5nIJY9j+cPLXvaMBi7bxUjpefbPKbCblWEkEX3wl1prgtCUu26
lhSa2X9+0u6Bk73npwlhjOMmvQsx5l/qDEMDJGhSFXTUReNj/Q91KakXfqMH0NW0
RLl0W7V87/45659jF5Bkj5fUGMmMyPGU3V1C2EUv3NqC02WW/RUklasI5HDPs7XR
hWSaCw9n2Egjh2w5dApbFym0Xe8rwCzbyMskrx7H4kMLdhMRoC0F7yuNVaQ+GU5h
bHQysE5jc+Vg54StP+EOLCMJdOEtzvaU88q2H+zTjmk7oXfe+4PEeqlPTO6DUCfN
2Qy5hW/esIRWMMvda+ulEekp4JDFJrPGOf7I3fryxUMSNOxOEmMkT7/p7cfaVn0b
ClIyX8yLzBnLoZ0rOtKvn9KwHELPolVt+sst2xSE478ANyik5uSAHWmV9PZIID2f
gwZOw9A4HAkel1yE51kWRJ0lhitUQ+RBIT3jNtKqxt6EJ0Uwodff/I4UCVQo4h3c
kJQbV1Qof2g/hIl8+9hb/68ieNZOR+nuA+WZAIFYNBf3NU9gtMC+ZA/4M9HMlk97
CGX7XraI72Gfw7BAHTIh7oaV/PCC0nKdHSQqGE12AJ/8nTxQMVAXr7OB5koxKmaX
I6IoJFIOh0Lcx7OZcsmTAFfG9Eji0hC4eSJr5xcXAP4/feo7BMRvofJcC+RiMMYZ
suROmhDf8H4C56dMe3PFs9cZQzs4S+YxbxPpfdLxLZJmzTq2NOboJzO8pBSy2kCW
mRIXQKwcdmRiImC109lT7G27TJHsNCIItyZOAmAf9jaGIBisIPr9mv/zWu7IQ5qa
GSrf4UstdDSSpPMs9zDsPfRIio+6K91LlRzB8OZh24BnZ/+uZLTfZKr3HtwKYEbm
2fuVfeWU6OXya+NU1XOAxq0FmFw1CB+GSBW3ADsYLdHlEpAivzNoGDa3M7X+vzw4
JShU2FdEeXl2FOo659nKxPoQVPqY7JSoCPbuKPsaPyCalESIfgb/3HYD/BodEiB2
RTYx3HyO8/9kbeEcs5v9Y+JTioyPv2BfzqTyu3U0s7TjWYcgjGhcx5LvVzpvvXQm
pyE7GeE/QoogqFpaMI2GvpF32BA1NBGFs2TOjyXfyUgQl/q9dJkeKItoMWQnVFEK
dE1j00SLR72mqWSmJPLHpCvqsS9pD5pqInkWDj1sbn5M49T/KcGl6y2eoZ5Ue7+h
eiI4TjgumO4zlHh4zkla2XEi9+1P7ppoFpR96EsiEpqy0x1UAvfUxGFTYJK30mxE
29LigZceCY8sz3NFqD6nff0h2jrpBsDRTDX7rKNysh9JAconk998uW5/2HOEir5s
3vgF0ARJySrYQP3AhL5LbDeGDiwQrcf/wcDv0uMhaEFhCFCIdP6zMWcz+ah4cPxY
8Hp/4a1pSr65aFOQKFbehd2fu5+KokjsuXAjqNvfRXsZq8/oOpRcQFHi5YzELc6w
8ggHRARBdm7Ow1bGDBFs47RZsV6m/qZt/CaHvGVacQG/3KW6+0EHISdzxpMuYEAr
7ed6hER4lAjYZRKjfIIzswe3reQOkrSLoDR0PlnmSL9TN8gCF2B4CeeaOamMomnE
TKrbgSVzSQXgSn4qeLtcXBeiWS4idKBzYm6ZNBl/tgEfjy4YWlY3srwDg+7HKNFH
OfQY6w0a+7ILOfqaSxr6hbQ7Ip3j/bNkfSsWm0saeWBFQPJwgm9czUIIeWObeZl3
UOsfkWrOVTtPmnZjPaqQcbJidRrnnra6Hw//2D/kTiiZ9bPBElAcQr8Qr4eTB6Ub
Al4hEeib35s/rIdbWp6zDDYYR61QG6ypGCcC6Tw64SzNji18y7ufNj5fRthk0xCH
SmQfvP5PJ92iskWfmIDQWwtnyoKi04XdFUVvrXqPCWVDU2Ixpo6DapGnKh9rUMlk
OpWYAG/bFb6dcOxjJ16dc4QNV3mMz7Z1EMEbdiQP2z7KHSZH6fXU7AJ0npdT8dvE
anCfjLujWlvf8fPNJ3gDpKBYoVQnX9GG7Wedfqfj0eYwlqi2KpetoroVGEyaOCQI
nJXFjR7XJDA8bT8ALNTExczXkg21VCQ3EMR5BTqX6O9k16jbmi9HZC2wLlrMh+V0
EHux2M2AT5Lvm53juwlKhCi69haCMxzwyIhc/OsDJkZ0JPxALVrRTGRqvy8PTPgK
dm0GNhxUr5cOhfTaJ5muWfvNyY2eLvQUBAnYZ7fhayB8hnDG7x7nRh+0fWi1RsM0
zn1nf4AbZvwM5RJnLpOKs7sUUyjk086t5ewmo1hJzfu7IUAjC2F6hlEH3O2APuzn
qKdDodGgWgwB9Y8rF5ysvD8F0LPP/XoDloLP4/c6CDZfYP0lnBM+HXOlcAr6ZX4B
5lS0PcZrh1qYckzUEa4q66gjDFdXl8Dn+1QelIfpPFl0GuVB2JPlAUz5tJwt9E2x
2u4kha/Ok+YZcr5u+MHvV0xoMTFdgYPfslZXaRjwePuZ0ZHwpqzeg8uWymW3EeE2
a1++VIU5PaFQt+D/Nq+pZLby/CRXqgj4e1bhCGYu2mfaXiTk59cZRVei+fHcs+h1
Z5/hHmuo3SU6JXCpIBZaFtFKm1jj/ueHWdtKVFAkAvGPHBF7nCvsRDudBNTV5aEV
Fe/Ra8awH6bAgi+jjMwpNyWoFejfNyVj2d7NyP6C6vuLOUEY7fpKLpQJ3qb/KDqb
zrqCaJT1BoARhapIzuaK8EzaoXgTT7P8jYc/+MdqSXSPg74Z+gaelAOokGcIaweZ
rijbIYewgWQsyLKvqk3bCxWcN5tCyJ4Z7jgdQtXHGeY3Jfwx2Lp6lzjEz0LC2iwg
E7vXGeaUQ0eXlezoX4NM7GV24d2YSIa4snbZXLWp19+4drv9605KoJExmZHVM2RR
Mo9Rdu9n1BuqfSxRLfWWTJX+rdVSR+lY9cpgK6a/LSzQPcNFC9etEvwN/MONNEHP
aWygV29OQNvlTRfI64NWu+LMYNIithUfykorYxUJwpJWq7f3XVfUMw0USVUPry5B
L5NVsBRfaIMPPAQEJaACYXTmT6Y95rN7Lvm86sV7GhdDah8QieH75mt2O3iEdyt2
pfGZB3UGaDtNacqtoCizPGi+A+YCsspRfvVherzqotl8ii/07ZxAtYgpvY5VEaoU
Kd9sCWLBHSgs4hz2FMDp9b+Mj8E7kwm/saN3v1Lhj7oJEzUA5g1urNbLALP3usjr
k8v9ZDQ062kHKFCr6JLVLleJv17xVo+KhNR8B9TCHvyMVh4TDJAz437xPwgzSVFv
Mm2QkJRXoz3rvu1wAti3FIRCsgzmwW73Qq5N5HluGLELbYspx13H3Qhd1ZsMyjo+
D2h3KSa2ai0W3PFp0Am6Trm/4Gdsjy5bTbQCyIB3h+ogvfoWgymhEgTe52OUwIkd
fWFK5L3ivBhaahRx3V+UnNI5cd5O4hANGv9Hm8nf+K6HCDKdhY7XTAWXOOAztTbj
ccQv27itYy0PpwlQ+dlFu77IyuDZ1d00xf+RhkWUdraLYQv7Whb5ZeW76/IWb8AY
nBbJtNc6bqz3jSw7FUdPdjXY5Jz5gKqoRGVQiuDCnwt9AxcdEQ3AW6vJx3d5ygdb
PMF8VF/yZBGBqSh9cSl4n7pIlRS6iQ5qwjDvkqpOm534A7uAqvzBeDV5lU+qOHcb
GfG16oTKRk7iHrlrVJUXsFPe6iKWBzvFKT0ftdA+8/e4zx21OoXyoDPQVV/0c8Uh
nURMVREgrDHHMvULYgJiNoYgJex4eUvvbNGKA1tsp2eG992avWomOEXcPPZmNhMr
SrI3crBStZ5vT3916ubXBDy9IBQtcYTopUH5P+3VQ5NrVpZrtkfAmKoL4LLhwecO
jKvV3nJQm8UkLzbz2gkppaTuqy2SWDlk95Hh/FkD6UoshssLfq51ad58ihGSs5BO
gatgyzjnvvC2LZnMtqAvGkItEM7yOB9ii0w7j7kDHesLGASWrYcWMYJr4f7eIIKi
AV1dGzaCYu5Dtd+DEVzvIx3iqGaKUCd5HvxbZiGzlSX1WUxImPtSeUOcadXak8Bf
FHIvHD2hUSedQima1xblMAQ5n+fDz+kVbJK0UIxFoZEYMMoVjjzsHuq4j1s9f3r9
umwlH1CrvxMoa09iJ2jz3BPw3PEoMtkakOPRwS7yN+8/mSkpI0hOdLkpo51qapcs
TNiKwYv5/pWpUQ3DkSj0Uk/tzk3frT4wkF79k+Yvpvtdz6UzfWidLSz96tC32B05
4GrlMSH4NfoY0zM0ANQ3RHJTVU0EYXYEryD8jPq/pxn+1Rp88lIEiEwmpsiCGESK
MBTb5UwT/TG1OsZkSZu+yskz0gdPZrQkGQe/6PZ+L9DjKKWitEPHFkTGfXcNOo3S
tI8zV0K1QYhX1sITJTr/3Kw2xaqFTsCW0Lf5NttBw6kooFwYG2oVrZ0NwcnQRpY5
7KeuPysi6UXgLgtL6m/+3inKE9vIkN84kKYF2I9MO92O9uGrqzUKXyEd3ANYAfz+
Xa1mKpAhsZ5li/dRrkOry2PMgZBiBAUFAOG4hcbSNK+xSqeSdi5LPJJAJdNMJSgG
O7TL4wxaigtQ7an1Vjw4RdXW7zFoMIIhByT1QVkwO5gmS+3LTdvAF/EERC+yHmlc
wUt9EJWx8vgKFP0TR3Jp5XEh9Ft3SRymsiHXNovgoLr+vNN82gMphkMlcBM6oMpu
HtmmXR+uvQz+tGqTBUOoZX/ZDTqZqn208QEcZ0g/3WFl106AGqfLd9ujPGRke0T4
O3H9kl/GhvGHiezcY/sgjsPtv/z1ryOWzusc55U+5fu12kKHFWjfyLZozL9D4he7
b+JGojyTEFrAHGvt5+kAo87wKx7rA0+7W7YbIvC7oDnXSTJepU4wbg5q0cu9Zx2Y
zzr0uATPZe1LnlSzvtePChMf0auwZAeMDnEs9xJKr9qULJU75eZR+OQJYmQF7qYa
3GiINNBzx2DvZ/ZTIc8bYIefeE5wLdS1YOd6HxPTmMAnbwkgoQJn/5DYDO/XYoyT
vwwS8/42ncKm+ZYpx1T5+Nk5liHokuNPAO0ntIHZ/GCY72LzYjsl6KHlvoyv998t
eYNbimX0/e4eUbA0lwBqGEkYvOp0zuR1kNcN+60XlLNF/Jy3kt+oITV2imdfgV+6
kFMJjCBdCWCg1y4rXl1d8RC/5cpNoeTu5oEGDaqbR2qgaqTfra0jMm8Hns12ZOFx
E/QMXY8jIjEnvPbkStilkmB9I7BccSwyJUKNHEnLbSn31DGCojikaXOOOvGdeaBS
Xe+CWdmnLXlWhumHswA2BaB0NLB9bMNfkK0zdNoIFGtUl3OUP0KdA9s6cxz4FyjU
n04oaZB/7lOLtbQj0p/xSuTq8BXEBj+5knWQLK7SCCOOGZNJvItatxXlRsgLbqlb
x9aW34NLlfHKusJQQ9BrEfkpzCxRVxsSbyMnM4pFdgwzRxLXH9Q4r58nQ8XWoOJj
qXy/JHoxELO/Sv5rnq++lDp6HEv+ILb8Mgv7+wgzkYMZQjLjWsysf6PBw0XblG33
Tmi3ywG9GmUCXLKFfMfr25gbTn/2aN8cU00l+yVWvD0d6MVeQXi+QTsernMi15h1
7OwNt2l54ss11hhNWShE0PVJe12YW5cj6WyitbxZwbAOvyivMumSTylmHqBK4hSh
S1XHxjlcGFvHdMyr7fuV7GH/zsT3/hlr+DyelgCujOoW5PgKEYE2+APizoSQS3k8
76jopJbWPNi4Ip2tfbsLc0ZX1IZ6BC/0LVj2+fl25FfspSHUu4RSeiLQIdFDmDGm
uLNMLgMqyKDz2obM04yQhTZlzsP8nf3VWhJxbcMtHMa1CifRfbJxPmhJWqsaKvES
kRDT3spcJ8uSC2fviPxsgMkeEYMVBdZxbssfDJ2LUiuVbJeF6Ddy3f/07tWmSvyq
BtLG7vLhFa+C1yVuc/tjuu1QN/uHaArQ9f7A9Jf5vf5vj745HOua7a1khpzi0ypY
E8qebg7XN4Z43zg+AytBfUjDWjNkZ9D6L9LaecdVRfRNMv18lUAHP8rVlNy//U+/
UO5fifi/so+6Z/UB+hs1cPFOs9joqswOVFs4h1KK4dh+DHNPahF9IZZXJUwLd6lJ
QKREGfLX/GHZZKveTv1hYFkMWIj8kZqcgtdabk2623/jA84Eq5XCM39Uvj61L24R
g8r2BavcTkCu/3RjgyysKa7pEoePUpw3Dgf2ZS4I+fsGU2kLLSMuGp8SVDSwaxk+
cU9MWY12wbADYRoGFG/n0AAl/GJPbFkVO92ZejrgVW005EsYgCaEU84tRYVmlDlB
x3SZ9/caELCTZSvyl6kuPXWYkBIecAFdRjvkH0BqlyP/BthPadepSMi/ZW7l0SXF
VPJqElSPu6Z18DHGYtvRlpBNkXmv2XXt6Yl5WexqMn9T0cILssjzjTEEfAymmA1Q
cPOCbtCmTe+jiA3OCeEfOdX/5mCyRPlVYDNgnsb10DKsWXVEYqMukEerm0VYxq//
+6yuohOni50WD+fDb2BbSZFUSjo4x2RDASbenVAEWkrqoHdysLNhL1E+qcYVzovj
SzzokAv0YAuurtSNd0Dv7Ez8RXtLemblEumjfRunAfV5wfM3r29uw3g3VM43FY/9
uEx74vRzAsbVadrEaOkeiRD9DGAhMIIRVp1uu5RjnI/tPWxyjeAHt1QRi0wzdB2M
y2uYMklajwj+liMft2ny5QFCTQheMqiivVqK60pLFig5omduc6AK5iH6eX31TWri
lNFCgh2C/czCpYlz8NLrrAgfACe+9oc+tLPydgwHZ7n36bJWsxHNnqot4qtfL924
xvQTmk510mWwCFtyJTwZK8kpg8ugilBuIedaD3uT3Q/DSzac1IRkXQK7xS0/d3DJ
YBVJ15W4QGRHnwLWOew1WYIV92IFb2j29jy62ulzmRX3NpYhVvGEmkDL+vlJdTTP
hFrTqe9D2PCF0LEk2KJy8FF4vvuDsz0rjlNhRSZ0i4WgLFDj3efasUCNqMUjCfe5
PNT5dwtBeRXt/ase5671y6Hwb79gGq5Uccglskj1cQSLczbuFMoXkhv+5BY0+EXq
GYkBc4F6byAwyZSkG9YR9JzLlRTgqP7tqTZipnNihJhYzwojsHENxPurELRkZF77
IGFSmKGYFd5e3tz60R+VHi+Aww4ayA1kvqPIOOTrDDCmiXlIkHszrccV62XHWWxl
JD4cPvTGofsVmA6UsBJyvTyjn/HqKZyPl1PHN/BNX035ubIAKFtZX3RJOuoGb8WL
bPWxloOzurdc5ojMzWiZA3iQMjWv706yjIZcVeaVvBbNZHzhwLNXSsNO0x9nUlPV
1xM3ivQPMoFA76L0Q+79YOJujmhC5OIjeocS9i4+tVWrB+C+0oqukWyQpUYVdaTG
SgjGLiByfRvPKSCTmX5T42K+0hJYLjmFWDnx0Iw3kF6KM0ZIXNef16EpbKpJjpvv
Q135AXrNiSI2OglrUDF3q9truhM9zMHko4TmN2k1oHLVidcXVIhoAjLVOnec8M61
v1fZCUhfYNkvgbrMD1zZMTlXzi9pZDeOew9opEFp0wYKFRGjsSPufB2kkA6FFBf4
vkKAK6G4RXpWk7w0Nf6cEK1TBFQgSR+J74QntWgX53n9ap6gbBOELKCG2AhCMMrL
2wl24isvHgVfJWFmwHGHphugLr8VHFfKkRxUdxcrEpMYiRlIgu5LxuUmYaJOfp7u
HJ4Y+ge0WxGZ2/7zumEH26DcFSSVZ5UGOugHBvg07sx3AmoA21l6MaL2F8ICV1pP
bBj0qndZ1/r04P8+y10BOm6e88wvPXuXd4bKQRigyca0x6jljoRtxuJviDFv8dmw
TttUEQDuYKRHbMMaG01I2n3eBUy18KTDyo2dKDTfYX0IfR2DphzQAQFHsEt1XVZ4
EyQKXZGXIRoKt8rnp8A4aRSVTIa8DNL90Gi88GZdbJ1zsLGJ6iOmOc3XFn/Q2rq0
aNlPdw3ZS0du/82mdzpGx45d3lNhZs8jaFYsUAiBEiSJ2uZeYxkFX64hEamUx6tV
e3ZKjHsg/O2FDEpQ6ZhsoqfYH6F75IyYfzNgK3Z7R5FCGOdr87KwOMGMAX1IyIYS
O4cBFkFxdiiZgNGpgVcYzHN/+NLcLZjMbjFK+LzzutAHiyccVpk71/AVgo5XODSb
nOGToIUk/cyavYU4FHHDiVYJ0S+UEuV2hT+MlZIpVyBa55swPSSXqbi7+OKcliDV
Gv/IEjax6y4cq8zTTGIEq6qbSx9BLsb8uSgb2TUe06u7hIj7APM+WYz9Fc3VKL97
bHAvPheOjbJDRX26US2AI5ZldDyUl5vOpq46TBwkxnfXdaDb/wmjMROPbM0v1ggp
2tSxwh4/cu4QK2YChm8h/5bl0PQNOa+K6ae1kdqiqi0B/+4Vo3K7szqHl1v9fu+O
l55Fa1Ku3dxUeUBN6PBdFbqr0mDLBHWspdPAidCE5i0Gj9S0GXnB0OPj9Ct6+I1r
32xdF8WESjjjSZlcSh/k96EgPNhPR6tRdsgvvbpiAZq1Pzrdvftr+hknnv7lOtuq
CyJ/spcLz++0sYPrk/KnemlS9DtV9FEqkILFIQiBy/U6+f9IREuQMRi6y2gQjQMn
TFly0gEnhhGCx7p24yg8CHZu3EFkjvpBALhFKqMUSo2gCYYV4kg1SBpbXyczpLKJ
r2Yh4iCcO+WgIGrQ2by4wuX7/aDLbZxtsurxL7ptT3npb/g9pINzqshQwIh1wuRr
+X6lEmI0tZuF1d/FIABxczCaL4WAHRy/vTEv8+CFFDDEECxtoFC2ixR84xQGAQYJ
3MDbC89K6jk0PAzPfb0ereQkdI2YDwUKL1faT/d/ntEWqxWo4QS4hYhmaJLRAYwX
4/us+2rM1d55Xz2Vil/7IWfyFqLIJIm8OG4yfYw02jE31ZAqESpuk9ZC+EOdIxlA
5ioWsxG7mhqb6w3ops/+dgOeq89lOv/JxbnUqf5orfHCovg3uRroPMIsEPC4tKyR
fuI/9FX8UKyEvyk6H+SobdVYdQ5bP/Sed1Zy3GxNYfi64D/ulLi9pTAYLTtwZou+
JvgKhmUqbUqpCer+FT6hcbwgECKtPROwGgVH5YJWACa5GiE26M0BILVy3xr4WeQ8
4qrlnCUXlpK3cRjm2EROgcOEjhdEOaqzmCuJVfPesM9fzFY+8xd3CKu8KZni8MmC
TqOoJ8rY3hAFzJPEnRqRKRikOv0cSIiw5hSqvbWZZa/j5ZlngIZCEAePOFkkIvpI
QAv99trvzqnW+EKuy5NwaLtR8rZKHnO0ngSFErAETErBJAdjAUX16FpXdtblLhaU
nJpOZ+8weqxs4ucOveN8RZREhmfXFPOLF5cCfL7I5P/n5H8HEAC9yHS+AZnx8CDT
AX9xuzy4wT4cqEqB0AP7BGx1UVEhzJRKSnRcVLy/TMyhjc82joooUv8TtPOKQr0k
u6l/4rwHnr96gKi/mLueIxjAskrrKQKO80y7+Gpv+rdcMRoS+dPV+8d+b0DwxWWb
fDEA1xy9NhDk3njLoef0088O1UIWLvCgDXpTGC7XGTAR6TgzaaW3p65VDzOqqJm4
L54zwnrIjLoAMWgw7WWm/r2R8tQzRQ+FXfCHo7ZuR5yUNwoF9g1SDIOqxAVJWtt3
KMlDGU6omcjZ9kQqOsNYQ6+MTtXiA8wwwHb41Z/r2mpevHK+eL0CnDHKJ4MjWzVz
tPsT2U01fUBU2jl01WaMaiH3eXm7tgGFxyAUj3makKieQAxFzGGDOYgbSxc5zf/b
Ate81BJjT/VaSUv0fs4b+poxW3sKV80E/zuPhCnfjZ5V3qGn6dGeE8oAflwN3wA5
7rtEkGyGsjP+0q7w+p3f1c99LM4uQr9du4qbtsCbRv4zH1UPIygOqX814z8kcjuv
ADA6jRqDgVVrlzzC61o8+tBUIQRwvwNFCoWEY3i5mIXGijdkawTSgwqwn5mlH4H0
uQaR8J/L/xulcm/fSTA65yOZNhsFQoczencIu4aN88gPMBvj+sbXEXJbzjditfXk
cYDJtstQljdyRI4Va34UqO384oGrHl1e9BXhrDAj9uukrjEa1Dop1C3QW2fzAo1f
28W86C61oLfg0kIJ3WpvxRA80MjDdMURC5rUT8Nlya4wsK0jWQJepBJVIYtJWAFO
C5oNMBrUhhoUUqAJsVZST40L6QkEvY8ihsMZV0284xvzP/7GohPON8gTg6Q275e2
z5NwzAjb7zLBFng2BANBxPZ1LFu9lmGLu6vCwNAhsUrwUK/POHGP7s0UFipxlPL0
fPp2LwNO6lg4YSJ5zgm+lR3XGDUrIxFpEvmQwP/D6BCF0FZY/KEZP3sIf4YIASfk
ENVNMHLT7L/q8ssDr2vjePL7aHiv4HNKrARtaRKAT61G61GEa0duCrEtDio4fD4v
3c+GzOqfc0FH67tXXES16Lw2qv1988NHIicOZ2uOdVRcQuAuTkd+ZGGO36fh+Heu
NfM2gvVxGFy9PUuO4PPH8/wer9YJp4RDd8jfR6NBmSnI2UnqokZiHufsU9G4PKWf
zc5Y+O+bOC730+faSn7vjskQIakUSUUgcEGNlYopN+NpBI+Jl+yDhN6iadP3PgsO
IxpVTta3FUSqeR5unmugw1SpzF/lJKoeslJIte3wbaXibGRkvo0gCpR3q5TM+5ML
uLObAxpHwL/1vle7sJbAQzK2/Pma1XjLWHdEtpjSXoODSNGreargXB/KIVobaqWn
oytuDtGtpgcS91vXYLBRb6ojngD0wJoI4kAogQFOtILVBqnS45vOCqsbumM6pc8v
YVQXfi5Y4nMia1PdL0D1MixXUh+fSajG6NQCc0M7ijwpW2nd5ahSHLxsNOPMdzu4
CcnntlQwGD+yNKEJKQtvqgy24lw1J7eBcpAPn0SPABF5f+199AMGr9XvBzWmCWbS
LB2NxlqzI3JXFh100e4qX+HBCwDBdlOyhxmHhfFHk9zUnmkN0+/BGjk25pWVul+3
/vwGRspudPfEgHA9XUvX0oKZl+tDWS0ARyxmEa4vP60bQ5nmDXje0n/jF6RMhnK5
ESOc6XzKVMVrXqP/lepvnVnA68KM1G2MrJz+m+eXwgl3/WV2znoo3+yZqYgPyejC
SaieU4Xq3QprmkH68d+vxxm3lCsCI1IT25W5LhsX+5dIuxojIRzF+KGpFQqGVR6A
B8V5c0dmA0kecZg3wp91Bj0tgUmasNTZEkNqEEq45n9EF5v5DlAsajnJfN16zVeo
vHudOsxWaVyZOpCtwRcDwiVGjS2ekvScy3vIy6us8CpV5iEuYuS4U+BdNnJ4MMk8
N86RpMzdPXfIK0KjuQlVbc2lMwxmUzzHpDSHId2jqNPMh0CDikL1zdiK1LFSv9Xu
0qbEmvRl+VY9jWCP/ZzHQa+EDcHMK2yncHvyYUnMd6kh25oGxfaUa+HEVOUENKP9
fQUgbbkJu+NkcU5AAeO4SKNahflYYArLVvsTfm+RqJaeZ41/zHjGL8TdGPUtnW/9
VDe7j93izZeuOzPPEI/X8b7hnU0ToYXfRXqVxYOswdJP28RAjgI7bPvkrBj7dxnX
WGS6X59is3TlybAaQCXTr68ZGAS8FrgvIzh86Z/B0nGyStxDWk0trC1rRku834pK
lX2gcBglqeNfQBMd5moQ2tLZqpmpjFbNXHktXyGbQvWbOo90qhCH702sY9l4iUS7
ko0fgMQidgVyLlWoNomnzN9L0cVYn+y9aTv0NV24CurBVs94gGOuYWPINoxTvlA9
Sy3v+djRBs/88cf/GiCwsqEl1bRywuRSMK3U/JJIo8oFc6ccCF9D2wu9mLSJOahy
oVDqFkwyk0iQ/tt9d1Vgw/Ak0vY56A/dzARZgbosXFygW+GQmV+Mc6f++z9ZsvY6
k3qLaVwPuE8Inu4Q/6I15iQObS7aSxPCE0ZE+ljQz3G/lkfrVNThjq6O9g4qdy/3
6KwKUIcSlyWDXYmCwXYlQMV4LuxLZVvsWgpNRO0dYHVoyQo6aFOmpiDsapbdWQug
YEG2D4lGBPlgTRnyEw2g0esT/COIq1plJEIwkgdo/2z4q8fsfhKvkiM1wi/GMM5N
phWAyNKYkKSE1Mfc1DR4WxkFWKF8D8sBHSlwZ32gM2ZTupn1r5YDd9EcxRId7LPB
6ckSdeLUvVTCceRddYyNF77qtR+jinLbHXrZOFswuvwIzkLuxjMyjW7rPDBE7DYp
iUOiyY45g45Ep95CSm0YByo1jVLFpXS4ShuvXOGFC9DwGAjyc/57ctcMQ+KXKFN4
DOW2AZ+TM2PWcAkRatnMKoIxC0iJUW0E/4KDiKs0/96QmN2+NvY7cYkL/6YLWtlT
ahQt7Hcbkfm1upko50DgOOanLxAFZ7TztI9RpA/m0LlwNFeqoMfyevjT8G+Ek1Sa
Fa+x45PXgO+IWyeMRc1DoO9YQ//ti4OsGFz9WYZwxs/2sm/t/PY77GbkRpPV2TfR
LijAIsXqf3m6X97aurawC40bGwguf3sBSBy6dZ2YEQktM61eMIReNtvn+wrTB1iG
BJjUSgEFuGAUWk8mL4ODWN972WspOIoB6Ih8D72jng8JHCbdmkBPxvl/Kjgnqxc8
l4j0X5Erf9qHD5C7b5CilZRn5ioOwGbQWHuFTf+mn7tZnytwrDyeVERp7GypsvQu
1NijvDlkSdXi7gz+g6mjk1gM46hkWpyyeMCYFmCWEuHIDvkUOFj2CyYiHGGCVR3Q
hiU4g26BEnEzp7Adn03lXdBLQ0UX8tnB6gXmaPatXFpZ0MYaokfq8anAd7IywCCa
fwspkopegKok3nPXkqcEW+xjAbxkr9Zq+RO7H1mC6q4TOsDu9rBlWwVboiQ8kCJw
MwYg2FwDk2/Ui6dvafdWU/eftOTAyEOoONd2DrA+cH61dpJw5Z7gKEZMbxD/Kq02
FXa8DBYNf7d+c9WjCVUnVfkjTXc2ODm51vR81BTSio3ZyJVJ9zVEutk3Oag06dZA
DR5U9B4611yCKCONQMBwroqsJFfVnFn2AZUHDV5s32iFpX3pv+zFsMvwyeT+Pcap
o8nRcON9CPbuif3kbBIy8GIJ6S4Fba5XkF47+Xt0CsR2jFHKGhjzuQWrbDieGr9e
A9lws2vMJX1IhCzl0NAJw82DH7uGOU7nBUIiFghCkNm42kKF5uTiYiVYcJop1e2k
oG8y9rI1uuju9WArr5G5te6QGtp9J4RXi8/BsKhYhKFNu6328mRhj8sFhPzuk0N9
Fak+tJeEnyzXq3DtRLe4TnGp2I0l5ImfLRs2uhfEN3Fnq92HCWSndg9Pwjv8tC5J
FXEThYZ9crbCLJEQwMBwUgXkavom37gnroXRxEBKNfVjUeeN72oF7P0iCm1gDUcT
YyYDduyYKfGAUj6i/02losflB9t0CUA3AIK3bPGi8UvXW7sgRGOtY+nf/dp2BMVY
UbO6sV5OVqwgR3TjHbGAvuBc01LuNXF/IWKfqwxQReZnctwQjNwNXIfdqre5RJbG
speeqgragVRs9yxI3EBfN2M7MSNVe9KLeZzZocwDXp+SrTZ7AjzrHTGLMRw6PXyQ
CridisgCJTeLO3e1SvfQ74TplBUBEncMAQVfPUHe6MOlY5RWB4Rz+lNBmIF5F09y
a8S3Dxgrr2oAQOFYK1/QNuYSXXhfwtZG5JFlnxWm5o/y4Zw1BMDCo2T3uOXdvsN1
M//EIYdckpvzS4lk0Nx3olh9Efdo2GrppEwYkBRQSNZVHR3c4B54ym+1sgGGPHWX
IrmHoy6JvjoD/6P8N1ZvsRh8ZOoODEiDNl/Mc0r/WanILLjC2/RAFro0tI7pWBjb
etd7g0F2hfUCHiySIr/LT/ov1YOBzZG9JOnAMEcDSqvCw8HHuE6MeKGPbrGGsMpw
aINuTKch2kGABgc5bjqCN++ebE/kescZqIUbqhyXwpCtTnAfaY3aS0cXGQI5NGC5
M36gsN3Uw6+Vve5Pb2PfSbabMwC+wblBndIdIdEhdDDSXcy4aAmdDMjlPcQzaOQH
OOg/sgna18iPMHjXGIr/NOP0hMqT4W93fihTYtX1nGLVbmXJpVk/8Bdto9KsvXeT
+euTxHREh1dYHm1X3lRv3tyKjZSFqxAO1JOAzzWcdx71vr3je/Q6WUncZuoIv/pN
xQIGRGZkvDEGud+OOqaa8Hv0YCEh9ovuvtNH6NGPHH/DAGatJy2DppL9X44n+9Ls
pwh+GAGmWp+mUPbpuC64AXTszbpESjRtjDNWAAXWNEbSJKU3oc2ClQ5japEg+9T2
ED60gUsBgZEQbnYXZk0b5pBw6JWjmt1xSYjTpey81PSwQOJD3Pog37+afvzyV/80
08Cta75LHX2SGqxlD+QCIeCrTIQWO4YZcZmNKlUjP2RbZR01zX2Jg4EOI/YQspUu
imR9KXfuSerod50lkKiosyE2DgaYTup71b/W/COidOFliMA1Uk5kdyYsQU+y7w1J
kdje2ofcQ3EnhN5PM1W83hpxxKvr6yYa8M7VPly1Mw4IsaQWUkjSbMu5jhWHgnsM
S28ho8yg0+btA0SXf3zqFZFc4y/pzcIluc3sKTeFPSzGsBzX+/OE+MNov7XFDbMw
QGbsqLr4NWmqjq+skHn+VeJsLO4tlFS/zB04MkU3Kmdjq6krwa0un4oLzg0ba4Zo
Tq7WZjht/7Nj/rVk0jqfi+QPGafsuSGUkWRQCI1H13G7p+lGvdZvxes99MW1Zzs0
d/xnciq1do3pBjUek+En+aruiBgLVrWnEi+51A/zHqRHcZbVRJveMmthmZ8kUkLP
zpafs7/wMq4ktM1ayjWvhhlxzlQMLdM+HFdsGOCglJ9XoMM+Dhaz0Z2Be81+NGMD
PO5pUhiy/mdJDwFFpXBSUsQpu/y84BidFUFGbWkVwyNjdt+M7QK1KbY/U2BFerZO
wDl6EOkFL0K5dB+nSDecQsKkiu946bpEgbptiGREnkjTOrwQ45g2xLA2OMiU0Pro
NLavFra10yqlCSWrfTf0+gA47C/xfGSffysHOofjeWyPu4NXf5oHQmx9PaPmalaj
4DDWMXFrP3VRs+kCCscZbB9VFbtr9r22Kx9QyZpHoK44y9GSfC8RYNnmHEK0ZilE
jbCSpxZXlV2qrE4C139MwDPhVTOjL6ihyXsWOa9ibdniL/bWeG6g/OiTky0UThCG
scE1CVtT/w181VgtgnlXS+R3p885kTJ2jpvIqQ9LSik9xF8jAstqmLunL6QD9I/c
C8pnzYkmX1oCAT5EKlkRnf9OV+3Loocc1mCk8Q7eB/TeC6pNP1u0TJEEVrEkbpaN
zQmB8e9wN1m/Vv2gyPhWd/kGE4ZTgGhvS2gvpKAgG6Z/Sq6MMkid4CX5ykkiddNe
NSS7A8yDaZ8/6ijz3bsitwFdhbRFvp0hdLz9qJA/rF/66YvX9+qAnxnGoP36Gki0
j9gwGSU3L6MPyTvenPCril1uX2tCHYbcDLcAKj0cy1cBFn3dmm4+nS20N/KFZ1uZ
krQCq2qIcQ1F0l1AkBClaL4iIvu9hf9ieNewo/FQP/+VcZ0/DaAYCKI09QPg4T0B
cPXaDXtiE8jBZ2sqK0HHk1xSlgpA/qmGOsH4cwLNINRRBsKhxLxwITPhkS0t0JIP
4NGmpfQQp9VQ+6Kv0GlKjNXFk1ichBQgdnFs2XNfsVySWIm/II5JFCENMrA5herZ
qAEn9C4zWiImpJd45dpr4OfWyQlYu4F+Gj5msWeNkWb24yRIBmTNDmYyg+jn0gXC
Bhy0GLW4cqkFItMfTmP+kfd8Hjkqt46qn9eIc5CJnVaLCQ9iKPH4ems3WJMYFwEx
od9R4X/LY1GGOMyqy+SC2E2FZD1lNN7HSrq5nJUZC6V7082zFxkZiUFNsskVgR22
jUkkaWUPrvHHjMcUf21WnYatRxCMgiHhiR7clDJ5L6a/8hGujLvYlBSvxAtzwNLJ
pxkI9RFybxOqRbIWss9ROz0LzoY5VCg+LA05vLrBYm2N5Fc7ALCfhUNxMCsgLFG+
4X8JhYYBLV+T8kW3ZCjIq3Zx5ANlsNHrMbbie1Sc6xzyHxtSdBQ6ZlgCmPP6Y8La
iMJPNtGNKqT+3nqQXJMZo8xKIdnKbFtdVrTJDHxx+j9eLYr4IM2uFGWFENrgUAal
nXTg4CU1w/gtZaEQvYeRJ08AlDIv16XpYnasE2E137O7evdFmUt6hZUR/5pIBH1y
1eE63G/2wKBHOJkyVNAVKZIArFbCbAC/QPmCflT1DUpEIfNqs4YA4LMMIIOiB6pC
BGhFhewjjgxL/KVvNuigQ/KunbalLOz80z6CtJVO4a41Z1KzRA+ieh1WzjWSqJ8a
kUzYPbOFcr1CWefCur6A7hnzv6POs+Z4XX32Em94p5rCOd+6uYZSBqPgQObdDWGN
k/hmt8ejMr6ktoFfcnp9WNF8fr9NnjPrnvvd0RpoAFsCuzY1AJDQdgfp1jWokJjf
5npdXAASNY70U/tuWRgN92JnaDtuWkg3hpbY9OsBZGrg7FlMgtH3DM70EExCtF1i
h3L/MJbqUn/P8QhxmwNgJBu78V7YkhS7VcKQ59XHXsxgu1b0KulwEWOqaL+DNbi1
0FCwQsRHX2h/57yTBduyY2Hm98E8lD1s8mkgCpCafU+fPbt2FRZN/J5j76slagQA
TBnCwg6wlRptdE8cJEFy6rD8FQi/HqObLTzxMg2/N4eR3j4lpk7su6bKRb8Ajolq
XpYCfhGn382vzppOwaCYVzQ7dSPy9DRouG/7K2LLcOX6DTMZKgtXy+PUS0HdtjGB
t9XN0mISrJ6EFqQ33/tQABIki4ubpgsaIK+kRExI9OO6DJvE6g2xicTzSYP89sOu
DsXaPTq/SWDj3RygT/ez9STkDs+OBeyVN2ZrWHA58v7Os1F0VtbPS4A0Tlackw3e
gwB3ScyKNaGRdQmzncjpG8ID4Jj6MK40nKEnKJECgrZJBTl5mf4/AsbZ0wfDIzet
NG7UCS0jK9GOLKfmNPGehMTtXrWz+pHNv9o8h31nJn6lKoaC3wEm3JUBo4ZFpZhD
Qd1RpeqoyKEsK61uE/ZpyTlKsSk/0V0kfG0a022JIoO1LP04Lf5b9ILFCRTBTRz1
CW2NDRXmQzGUEQkJspVTjNEL3FfngJVqjStuzVOzCx53SzCMfTcoBDnB9+izvHyV
UqoUbkOrL99eCDOAPnxFSlfDHnfKi82PWoLbQgG/pb15TkFb/JkmPL/Z2G1it5GW
oVZOWGaSsyIQOn3tJwdvVvM2hSSWqhA59wGAfIVL0x4MUldWMv0UrZCt5hfgteWV
6t0Tgtnbt5OC6I4rYzo6+xjH9sqDBp+xvveocM8T8B6waIqZOr8HGV7rWby5MVis
s3G8FUis7mtZyqYEDNDUgc8Z1j739P4z5N1gLg8jC0x+79wUdGPO3csrecEGa3SV
Hnz8tnIVKVjnS4kTMyKrG3xysvBWtRQkfXnOxhIAqk/ORIIu1ZkRuXR2qteCKBcs
IpFCHvtY6c0mcqsmGzR0JctkawcTXzeTNAQn1G9l1CT9MQGxV8IlZahCDE/MfoyP
jV+Vw7SLBJyigwxOaExJQmW6C5LIXxLHskrurqMEDdKFEHBf7OVKfe8lprDZRgNo
/be1NBIg6fSQoBIhvI0Thedoqi3JjkSfTezn/A+4cVEHdSd0pGdOfSQlGOHHx5UN
YqPMkHk/Z1YSvquniNMkKiaC2D6WTb+k96v+lxPl4DP/o/wWsdFL5R38/gAiTbQD
evzVX1OIt+3E/+rnZzDEq9n17CO1naoTStOJifRmlZ11ST9uU9xtDuIwfcL58Rv3
CTAGBME49ZfNVlW7n9l+zUVBgAYjH+ckljF2qVdtimGqwVCvgHVZaLY/PCxFbz7Q
rTM8FDm3wJKzmoJCYQed9b262+VbI4m0gNbXxVjuBmkRFbBhsbByGnFV9iPo5tAI
f1cyUoimK/WzRcU/bETKdZTF/0yZcit2Wkbk3LdH1y5O6jekUTy6JSI4pVCOsEqz
H9ixHX5h8t2jjXLnf9U35l7fRTckB+l8jK2Yd0t/DRI0nBh+uE+ku+XcDyhRB/r3
Wzg+C+0VsUIgSgWECWmqHhG05iVDElbUIbWgaN4TJkXFYNgiWfD0wFJXSTG/tnYJ
4+iBF+g/M4X8voc5I8sBwjvKLKvjlFX5Bo6ka/HvfQsAna8dmTkOojTqotxt+iNq
IRWv9PGcdeQCkSQixftzGMRMXIuIz7In1rhKzhRtAUJmdXaVCPqAYNauv94Audcx
6/2zLk/oyMq7VgaUK1Uk0lALvFxKfaBrKW1L30Yk+ikgt/CvU8abrC0X86+hcxSt
WYxllthuUitzNMqwmMC4Y7o4mI3a5VlYNpqfBC7JJj2Aa8hnb9osU/565oKj3XPi
4qYzqE7sOfHrBv1TZnQK4Tx5aAMAG9gRw5xm2pj51a7jumRmJIS49O+XLyB3K42V
ZTVQOXANzbFPB2eWnpm8flooNxpUoPMahN2q8LZHFsaKLiMNcJbntHrdJP8VZm4d
v9qyn8KIB9SuacRsWR29TB7LY0wpfB7HVM6I+vZ3L+jmlbuTaxCIhwbgvLXZsSb+
sTelQRNbVdVERdhE2CEkDqeZ56WY76o8qd2b1P5H7/F2qBwzXLALSrM/uYsYkbVJ
jkUIwFFHJvVoTRqoEsxUM97i79BPi3Q4FrTdbaqMGX1wM3BBprjY8WVkuiPKqtis
Cd4K9W+gF6Eq2lx9xY6ZUTeO1BQSd2tZH3YJes/pziv3+79Vi+jpekhIgpaAGIsh
Fon0SlwS9r4XI1aREzGpRWB8y7fY6t+f4g8nOj/6HBM1G5cKulPY7u70/4oDjp4Q
eynOuI9sBHYX7UTmnhROBywvuXe6W0J9vw+o+PAbB8nFJIClbEKhNDUOttmOvHUY
ePKuYf9okqlIGFg3O+OAvTPEzKSBuK+5o/YVI54dlDTuPdsGMrxDmy2RQSP9MMoS
vG/59+A1hU6jgDQn1sIYpJvTYWwrKzUEEOyQruuuCWf23r7znVbwqIKlr9Q/MQkl
assxkxBhbW7Y33JySTWsXnA7FfluO1dkhYKxBij1lhmCCzcHqKVfQUWy5njUZjEi
rUJU8S1+EmjH/7IbIcghQuOMisvXJRlYJnGkjqfdBHC2uLY0ZAketnumoUW2C7dr
MpVQUgEY9aslwj+mAZrr771go2sRMeOiNTHMQ3NgjkCGa2OrSDFZUWi4pTt46RBx
HjfJXN7q72liCR0ZyNp71IR7FJuiMDuSFoITH3BPoE/JGmFzGqRtcHO8K8jH/tex
MYrXTA+H2OKp8VIwQ3qBl5UtWE/a2cADxJrdufn1IIIPXbvrtC9QXaAJWitzafM7
049m2ItAgoSnQ8WtQoE7Llui2uOxohERgHPqqdXhv4P1aTwruLdujPHlzgfBtmCF
Q97lTYp56l1svLh8ePbyO1fhUNVUVb8jZyWfZwafviJPLQ1NBW4qVJ+KCIdvTLmK
p1RG08am4hw7ugGkDQpsNXDQRPRic4k/tzUfpaoh3CXC6Cggppr9yi7pAsKUjVcN
dDiWIRvo/ApclxmaBZBmPRawh9NBTsiFsvYSXjtdj/qkhQq2a4aJ2m6mB06x6rSL
K+qTIsuwPB6qzagfnYtKU+LZBBqf0KRymsakEu2FUS4NTADcqrLU/UFlMClKeiva
GU+AtL3HuG5UbdHeo1IaFkzIusxX7si5ajEtphHeW8keYIiXFAqMs9bTLfUVFGjn
JAhA69lcmxY5/GbavAQ4UaJfOZct5hGNzHZk+nEaS6Xzd3Gl4hVfL5WHxuPGoyA1
gJGpDB4a5CR2/ck6ZUS0gJoJ0TQhcWuHOE0UizVeQz8x8vuJghuF9osB59jtrUoG
gf7A3UeVpYJyx1srfXt5i8ceHm1waN/HqX5rQ8ASFwXXrI1jho4Xa52IdPmvUS7g
LlXDq0c7L20hFqvns3dBiRgJQgLB7Sja/71D81WkOgP3DnUmYCo/+WbONMi7x0y8
/n6mlbSRYrYvWqF9G8RjRSZ6eZdVh3N/vJAk/1M5I8AKuI8SDsa0/cdBppN3N/cy
fdS5pZa2LlnuroKapTCQmqGyT8iDtq7k+7d4u4h+/dEZGHAZF0eooozdH3+1J2nv
wLyAiz8b5h7hkFtt6d47pDaUlx5Z+uzPnvIKxpxedHJ3Ds1X2uEswExejgGDKgWN
pAW/lFrtQjaZhzsTYZwtWQAtsKHXd3LSFtys+StPD/V2Bvu9D2PLosUy0SKal6Rt
lOMlitvWOlhji7Vjjo4q7v6pRFB7PCP7ac7qBFXPm2pv54G67FIoBlCYfFOhe4jj
uirNhxkCUX3Em3BidsCUhpE6bFi6KTKAGsjKcaw87RVQfPRUmcAkvEyW3tk9/QlV
3+8ptZpsjcVFnZsh/AAAfY7zDgpUrOSqtBQ0quVOugFCTAoi14+pVah4bydC2/ft
a1P3b0d56XTDjzHPeSh15UZFf3kxgpOEEzoOmdVrH02uSjjrlzCEackTKpg3RLGL
Rt9PhnTT/LFJhGgxaL5QYP6IA9q5sFMPCWTJs53llXAxThd5TAIlNKCIBnqXaHkl
zNY0HFIqJVSM1JOj8MbgP3raTfgkRALPKafQQcNitMlc/An/lYmHXSFXSvT/kslQ
hObWaoDfi9gpNcsBBELMRsBitohf53e3gnaziF6l95VUL6iWMKeGyXGfT5VChBDK
VVoIozc2hl+Mbf9HTqf6tevjNILnTE6xsJ+EeqNgGFfCNkjw1Vr1sDIysebZYqWZ
TNIVwbvrNiJRS1h4HpwKX5tO6PB/SXDngC7hMu5jys0jedpERQcrW8Fb14/70Qnp
HqpTKDAx9pmVOxRKZDfCLWeg9VrszmlyPxGl94msGvnzfJxrGMmgHv5p5zWoDozt
O4IpD5THxQgPELHvZwDIlWm42xyrTB3d44hcNzQCbqjs7InlxBPmSAw+mC512j8A
QZ2+mWfgWtcbdd31ZPtelz1E6sEAAuzVHHHLnJRh6p+ymRLMYyEtu79RQWJ8Asa0
cmK3FnGMZY/cxyAH/9pwPdN6czBfLQpb/jt/UiCRPCW5V85koBMlG3SnREn4lhFk
+eaiUSvTttscMkrdLuEhLW68j2C+W8o2FSHIPNvm+rYzs7rYuijZA27Mo/g+T3SG
Vb+5LvTUlmIWb7yXVOCAgmZbNjPuhzZytwdaVk/yUBUtZYFEbWwt99F7XJ/efbUp
FF76OWHhN0T2pzZ51cr2JEBkY5uPhLWJdrz2TVwj44KwUaMK54P2tdG7fSryIi/0
CMxLVpfggCNi5xsoZkoZdS9IFvCEk9Bk7hD/DZTBxZhSq4VyIxztJ+cfcUW4xO54
yHrjxAz1zVqhlmmDaAaSTQ1/N6zHmdO6eVE8nQxA99Hu0UQzxgg9btX82GPVTSFi
xEfq50M7qtvdz4lNXLt0eBN32S8nrDRHwZiJJQ7GVBLisU9ZhPp8jMK1cbixxPMP
SOi3ohkRy1S+Z0pmUufXqPQopgMj9H27JonKcamf+e6gbrPxw4/3NlsnJsoNg5Hp
AmgqG3v0emVYODD1F3Q1ZEUaqKpqf8gW1y3fSuPpxt/XHLD2TSlvKuh2vrewQofi
pPo0sjHD9CGxvl7hTXEZKLMBUuJIqC1OUC7C9cJTccoEO+gHjzSTRMbQWKNR6HQE
HEQGIrfr6DSvVjP/fyjPtDuOVfCs39MfNGYvec7SyDerLsnFOcO6WAuS02c/uNvr
tD7p0OGVRmE4MPan28TjxaszUNxO7YpSBwlwhmiZBSV5oc3br1V55YFYV9f9SetI
3HPU6ksdS03OxhQFfAu77XYCRIzr0LQkieVqFlYg4UoVEiC/kIO9gUDAT4FbUNZf
CPle9KONDeB15G5ZPoqHbQLyGO2/S+KTEt60tpmRe4Fl0LNZ15Fdv38mHHqrOvHy
wos4zUZ/mT0upUtX5k8NB9DWvrUL3Z1W46Xk0bkNenKNgm9oH3EsyscaZDIqBnpM
XUJgdAmJ8WgmBkfHqtAN2PDVcqrUHsFG9FNGpw0jRxNj1Gk6gNm5XaPWgRkzQCXb
NTjpdWCAwzwGJUHmvfXAW9qmwko3c5kvMT5S0EmCdEwByVLeJrBBmUC4FQ30iUMv
pYz5HAob/gHRy9lrB9Pl5JL6+jIp1KJnlrws3LQPlLgNQDPLWlJqcsmEyBAmA1bd
UdXp0IqUL/MkwkZrCpswrnW7BM5DuRZJRRRAclQu0A4uzfPSh5mjtc275Zg8Du7w
DPiRolk4C2cdPk8LiWxx4KA1sRzjPcq2jq7wWVdwbqj9F6WpgdsLfWw6WTLoqAon
jnXhwtKYx5rv5lXKiwF3AqPt4mpUXKn+uJ7ytobXGYCeX8Wjtu+qk38MY44wihRk
hu6R9rlVO5PMGfdmYqTVRdlnOvg/bOXumWfQECKVbyIoL7m39QOgj0JclJpxPUcE
h64G3PFTVcSMU4JGI0lZrhy+lBlu2vy3288FB/26HuUcnAuBNr4nc6nwxs81j5ho
Dkn9HxgNdhr4gEs8H77R7N1IVDn53rxptxoZjj3hlJ5WfCjgjER7eiqYHDHiwKSC
WRL7+hrE7UfaFPguMkNjicOYYEr7ueiPYIFuOfktXJAAV73i48DqwDSe1cEODxZ3
0L3UC2blmV1LsGwPvetpdXj4wesyJ9CG4VWFf8OLfXhnzoMQKvIOlVZXIYVev146
ChnSXEkObAFO2PEGWES3pv3ztw+Ze/sQo1sH8GPrgtLTFbqBYih8F3sGXAInADbY
KS28BH5OgCcuwOTaXjleirKXch/3Vf2jUYqk2AimfROboYx7GrAjXJp6fAXWps2o
/hMiVHytubECXuCnLF9Xv7KFouK12rxUtiK+uwt8yi6jcf+4umA6kzskoMydnpKE
GZwmXwhVbq+4ZzlNE0LsH//7WDCLzHwMOJ/dkgpT6Qum2CIyp/icb7BxVsgPd6Q+
iriRGptdjw0xdNgnq9wLJpMhCTYewaegPJHYKomz9UvEilArGvYkhxzX6CiLcdjZ
6dol81yN479+7crZA+OcGdepmkVjOjRzyak13j9JUKdF+yzqlghwD842vsARqFy/
Q3QheN06r1SMnsZMNl2InhFbzGnfAL01JJni9MfFUwU746OVw11PKXDDYfxxLeZ6
Ygc+VwHnGA8C8+NPe9XevYg4vyPtexoOOO2+KVK5C8U81bLAffRCCV5KGRB3KvcO
Wyu1xT/TrGE0Xli65sEZowabB47jDlG/YlONexvAsDYYoYQ0OzbGIuwpu08GvGvA
P2K5FSaVbej0MdbtPj+hUNKrICj5G+2DtLYEjDv7ovTHcrIQkzpbqXd/5L6V6CHM
LCbeIhTLKUW3mUgo36G0c2I5Qg2ktnVGM34eXNg3DeH8xmqN8wRy6hZNTxwSwjPy
jjkI66glb0K3DXA7ZMB+OZrQyoLS+czVtdvNcbPWox0+CuFrkKTQg/qfMJUyc9wr
fTRs46iBkVpeRiQCDrWUqgCbNsp5wsBDs4rGXo8QcHD2VZ2187vd9qp1/EhxX2JS
V9gUVKjUGG4ZKGBuOSNFoOR5IpmsIsyS5ajH9Biee0aHt1S+08Ay3gBaWt0mKF/r
dWqk3Y4eL3BiApsdthUX9VsSf29MWH1DcudsCibAUupJHf4Nr1vJhO2vLwe2qpgb
twIJ+kSpP0X627zp7A79wKssdTOgyebLGGh6wuBEcxqxHvMdQjftDSPdgC4jcr+2
pF09kBwS3Gd1+oAHMZkB9HhOjAcduy6QvffUaxw5mxWTCgme3TLxVHKKdt0QlGVl
Fs/ll12Z6bQ5MJHXz32z41LL7qbLtABvOeHH9T4NhSCSkjBxFEV7/JrlhTssJPa0
hrdk6fVgR7T409bmqg389d1L2zUvRTq5pKuBFXX47UTsX+pPixMN9j2U/9nIKQKP
Xo209+aKZGYjN248ZxmZFaHgc4mN+cGEwRKc7qQAGrSrKXaTAdMWKh7aKLJPo06b
GzSX2h8dYpiU9pMRatUYkEe4HCV8/np1tV/1Hqsm7JH/k9gbv//lLg6adfVg/Z6x
gHuNWYbzoHMj31YEBSFV3pTC244dstZLjlk3ZgbrdNKi8bJUsjnimNeMUqUgVpq6
+DcPUYMzst4pq3CrGUQow3VSCqT1O16guUcq7Phvyfu6IBgkN8ZOPhHeoqsQoSOa
JH68k8U9PCVK35PSic3ebfp0Ey8Rj25Oy9O9TVo4z9hGFJaIvMZ17cloVjEYWIIa
wI9CMdKPOZl4vS0PP4Y6R/ngQpGgjBXN2hs/jBOG1V4BPOdLVPRFoHrVMBwDohvq
weHjUG9rCEvRTJxrYTbD1F6PWBokhF7xctCYpp3UXHS651790AR/Rh4lui+zxZqb
NxQqLSm+ciSs148L48AX/5QKUDoz+eJs2CLYCleW03nkosnfaA35GZSXh5gOckPe
WFoBDqm+btoYSJHMasoBkv/chydg61ON5LBCPzxWJeq60cQn1gR5Y6sz/yZKBBIt
xuZZMk18oZbk1KgELWmXB8ELvThiNBFC4FgcpIPb16gUfPJNLxcmoM3CvzDkt+aN
YLU1IEB5UtbmCBvq+mefewDjeCbo+HV3y+l607Id863NnADhI2KwBAITOejgLugw
nDvO5B2L0tpY1M3aoIjtFdK+tNEz3sVnnWm6oDFWw+oV2GkkeES2j1YneD4TOFzI
QM+U6IE8U60X3oYpeHL5aFreRTUz6ujkQGOsbpubeXt0ML2JfIn833Hyz3Y5fBKQ
8Gp33u4fI1jDUEFPzRFVjYPPVeIAYBY7HDNr/L3F512lsMPRczDOsh/GUKm3m6JZ
MGUqz1ypNamia44hcHCoLLuMKDfP9CvXDqhAGX4WjvrNIxcOX6om1MpHFfixJ471
NSUbezPCWHxOSwEiQzIU1/EMhTv2fycj8gSbzlqkGq+AWlD30N0LRIwMWcG3pE9W
xtU9SE5wGE73twIhiQSXfa6zov2HPwyCUc3SMjABieRTzc5H/qGIh30s7v8IOM8x
+5D2Abisbp1f+xDPVerLr94UszYoUAiKPyfETQPlnt+QM2zxJdv+tsuhYwpjCUb4
AjMWVr2BeHEruQrY+nBIl/+hzyqAWG5GYmLdlOA2OYoUoQghMUcqVHcMUX43fIVr
gAOJ6yQG2QxX1ZzpVdGAjtQAixDMORYu8nkwhmWq6+ia7Uu0st488cdJiHfPqOe6
J2+2Eet/A1rNbneBP6n0erpF2444AfU/R5eotv7CxvYjUjZRde7DDjSzrH3Vurvu
KfaWgFTI/vkIeEiBisKgZocD/aHx21Ho6QFhmkI4NhzfO+L4Mf6ORCG6wdPNMRs9
6YwQto79tGmy9NSz6hu1PrihFOyAaxl66IkBSUzbrNumMLHJO3WEtpN7zoesPFIt
fy6OFn//8DacqZeI/aNiQBtpyDnOUx+rlWfdJkt7pS9Cvfr1Uf41CcgFhL1JOnTS
11YlMR4UZnYEN3QvVmrrnntzodbBHhO6HhQOlMpMR4DLVQJFEKIXWbQM/YSyu5qW
vdc+jnRLKIcbLxaSRhzOhdFOwT+0raqjtN5ZxQsYzC/rhkxYVq7+wYAgPdUkZIhB
PpnC2vIVOp9xg+JGLagaKtQaF9X2ElM1gelar/9Ef2q67zvoRzAg81bRBFJojXUl
S7xijwcPQUsiRcWgIP/3QqXqW3XUqbvHkwlEKnQTOfAD8WSN+Ny7X3okfxzRpCo5
SshtfP77yc/UfkjGzVY6mliAkG0MSp0T+0s31KcSRUM0x9Ez+tK0/N1e9DeshdcY
731VTV/dU2DWMF1PlZ78uJzYL3XPdcq/tek2wt94NCnlpS+czuY9RwNsgLj2NSsC
cKFw3J06hEw7wagDeI26PK/ISK1o61VR8T4gWHOzbgDNUZdRAR8NhsBq1I3E/2sV
hwG+/Q7CPcXmz/vzcB+WOjdCOaa4RfwTIDvG74hd/+eUBdV5msuPVTn9L1VJHaiK
H105/u73eCBSZjW0DwQqjMU4RKElfd0jCAHi8ZyMfreHlW0IASQI4dx/IVFKZ3M+
zepus0xvT9ZBy0e+2u6Sw4IVcIqeOyrTY7ZXjpxyq//3vDB85h68/XSX6g4vrp74
+Zu9emcvfsT3DulU+TUYFCFVtazMskI96aHoHn38tC/iZdHRtNwqTDCKlSFbnuIk
BkuH9D77JJIES32+tZx9DzqVVmtHI04GD4VCC9PhNKWkE5P0BNu5BSdz3xpn/DhH
FJkFNbdpulWZIyGhZ77eMp/n3kYK9NFImsQSUDHwzS60N6VOmjeMR3FFMrjowSeu
aXwO0zVQAT1uA1u+1kCNdOHFFT3P0T2tt87abl2PCvxRKKuvfVb56Hc/F/YyWVoP
HgIKHng9zItT7OhE7fErfJbkxOnKMUFjbSeVGL/XYgWZYVe+dhMgnlC5n8IqB5n+
yYIUeG3iLWOUhUBanWYzKK3T4/1yj+2dmGfAae7ovlM2m0I5xxX4RncCuiyHRUXR
npWFDOCY8ellrOKtsN5CBE4NqOD50Z8IIyxEdpg5VkpNUjC2Ay2DGBrHLvAlcwGD
WtCCQaRzDeCIeqv11konR7fDLQukvTcgT7uDuc3KiH1xze3xG6sCzaLbZcQz5jvw
J+SQF/5GbIpuzOHzoZfK3naGVyZuuNKMyWYeYP/c0hHcnbUhVKyhn3vBtxzc8+KZ
j06Jph4KNHHRbUSnDLhm7Xo8lCm6r9RZeak0AqtDWXT+VOnUeVnXHBnzZBTc9ZyU
HExr/IR9H9N4dcc6UXNU/nEpB4fJrXWHNpRzS1+XFGoplIKfdZGhSo8J8grK4xuX
PmjTSnvvfj8jOgkZmnuFzoMDlaLsdBqFBsr90/7D/jvQIA/33zRUJMHfdjrDnVk7
skIxocabJmxEu/X9AzfodCIOIbvjUjY6zAye/KT4dVlSgrYnahU+qZf9+eKuBAbe
iftfFVZ7eAKIQN1+S0+rGL5origcDGlEpBzxlASajs4PAKavzgZUzVFkuqEpg6iw
p5FMFxk5Ej+uLVCCR2adRtOx4soisP6S58n0Uo/LgVxXybvhWR9bL64BJJYbzRvI
5BzCdmzc8Rude/1fjiQH0D4IDbcLWmLEKZebNN6KvZp4qckIxjg+2IzeThY2AieT
GVlNTF1ETKkH9QEs1cqWIXnhUmUCKPSFYM+igIEexqVPJXSsuJqvL95ixMKEiO53
ig2tN+GU+9ofAhU/pf7W9+on3n3evyWaIg5nlxnSzT3dK72h8hKV9S3u+4e+3EWq
IvOXkfo+6y8E2dPzIHpWKNH5MmYwJFMDyrzWmlOXjkF+k1kWLoS6DtrAu1PxIXsp
OiL7Nntkx4RlL3Txaal5idy6W3XtPRDKr27fSODvcTe0CTy09qUfkg9OJ4Y/Jwib
qg4PMPCsF8o49aNsYbsHhuNAKVk6NDlQ8iZP0uxwurEC7MCtouFQX8pz41c1FVM2
AVdulD1YK4qwABepYeltFz4dtp4E9kqLhuK7LO/Wsp62FTso6dyEkG3HCOsKwHsF
WQ4+8OqzA0w7rGr4+Ftrg7I8t1/17jez3/D52dsz87uYqnZaLDCvAXFMqW3k282y
Ve9E/3/i7JOOpDszofttv0Sb/PhSgTpT3JKlMXyfQMTzx3ftGOxH7q75EwCsquUK
ISIt4pkBS/H3LvabihWt7D84fGIMIrVxXP4pXSXnnAX6JUE+1M+dFNRtFNv9Q8bS
CPLIobKTkZaPV+NSKaubBsuRVHySuYfxhAuAUIrSoexDpuah3VLaiUdyE9GELsMv
XyX3tYj9kQyZhTLXIyDGHbdg3oALBPmDSeLwqsasa2z3RttkLP9J1PS5OquePm0/
eB8COJmYjAvV2fxNSYoKd6w1Jb2p/J1eNozD3Guzx064RujdUtBczepAHNwc7of6
QipNiMhieOaET6VTQUbsZXNndCVSoRxuZTHepA2mKKGH2Mm4hzAYQd5nm8Gy1h5m
pODCljHFHTtb/bcee88LEw9yxBqfLadhPS1f927hq0RuYlSAikqRy92iQdBaTzMs
0HGc9pGDpEtatkUQjCt6SN/fIjs35x8mkJT/IF6NH8c/uiuF655MrSgwSGF5cdhp
s08CF61oQyLwErY5sEE/jBnCtExx6KDkQA61UD792ICaz9aUTI8tMVzHdJ0TEwNY
47Xwofqa32cJP2TpYhhELQUxmZr+yNQ5VJPTywclnTmxjf/mQtLVPF80550KSm5G
QpIHunavpWhIIhFsLg/jSQ16HgLrXlmNqYOtPMGaLw/6VXMf5p7ezZl6rtbwT2sL
iV9j2D9meBA5yc97WY0u/Q/8GdOFb03ELw5d5Y4Oez2QXoXzAO65VPOrN9PZ/DKC
Fz62+nrvQkewXeTjWthPTXVDXwUzNYH9SIXzroppCJZ494D3UChT12K7FrklnoOI
pJoX4HbIFIU9+5ap3kAmByOnERfdCuCf0ZuyTd1lgjaFxsr+Ia3BhBSQ9Iyjbohs
Q6jmpGxBKpCtni9QsdEUxOJCn0N4jMFO/A3sNni3x9rlgaZ4ywAnqBd5PFC4vdUH
A7QaYWM7/KBTbLQiqvuG9xl6exZMxjbJrptS/aKUwPJq1GwAK2KWqtwmR5C0kpiv
lPw4ktl7wIxK88te4P0oCXXUiECkEbaVkyARybmBQ8wfjwjjMh3dbDcOvzzChSvI
/JW3niTD+oTknoQ3a8Mbo/LmYZ1bkhJ0n5HDV8zfmuB6lUAwM0pn7yfVK5yvZIoh
654hsmxDvGV9qVkMW1hT72pMdkTJWq0gVV+Z2Tv6uz6sIqvJY6R0n4p396Z2iV4f
ORoUVe2YgEK29ZRSAXyJsrOpEfZr34WkFZkhwlQJPyjhYPYVIF1GbR/65XCbNKXr
izWw8GKjZDOElselD7DXF6DJTLbFIMBeB/K8lbJoHSo35BZ4FNiubcieCeaQiZDF
FaT75qcxb9SaxuJlm24+QsdNY+wAmb0gyD8Ofkv+WXgX4s9ng2iGbSiNpiE27nha
322dU/NW82zKHco09JXR3h4AIhkobS1rBylV+UMYxGBOSSLB/yLGzTz+OxjP2Zut
0VDNi3+mSxiagzxoFSNTgbdN+/MRnN4XR5Ul2DN8WpUdaD1kHI//SjOi229VsIVh
WN1tKYBXZfo/cwDbCPPQsnG7JMJ8ATEzzIoOrsnI9wIzIMJ+nwuj87Y4X/PWEogX
eLukDfPMrJreYlllLI8c6ZNqWUQ6CVUmQURqlWTcgtWr/eHS/w1P2oN2quhAQVbI
Mos/AMunRwZe4E5bJZKj1Z5/K+8DF9SUEqkN0dh8oKgz7UdeTd1wsohuBpHvqgT6
p2lItHA7XPfGVtF3uIEEWWaMm8hp7vwrpgcLTqOGXMtZT8uw4qC7wV1ONZtxnnOa
/7ywR3tKAWHqQAZ+fjNQeTIXdZU8aegIM0ZF8CViXG6AC6P4HQTw5+edMoeZdPiy
Mlcx0gGP7xrno+uR+TrgNfopx4dC9I+aWIwoYPOaRjp6L/pDCuTqMJh9kbhIIKuz
IAWoWZMdABnopyuxtMbd5eyKv+doA97yeaMPn0WdWVZSH7FhCS25PajtQMk8iQEY
zsme06ltbw9btgvvhuoicimTlkWkAHqMgfeXAFZxS3S7A1ns/El13/TZGuwmCpp4
53sGf5C0vO1Bi5RobUFlc5wFUL4rbf4c5NXmmUGyOxQr8H5lENpcxzyqJfI0Edpr
3QJocPtNtJxsYQ7ZTHxpod6bxqNMWwY06V++dQvTs8ZFfKw/FQZf4Ujy1OX/a+gW
pZenJAoVELN5VfPutSEA5RwfIoHImdX702IvSSdjYVwRSIChG6SJ2aBMkbyGL2Oq
u+J+IgO/1HroSM04pgQHozi48lXuGJaNEbnVw8ROgVpdv7bxE2dkRnbZvttrCsKu
QixWkheTe6Jc7nUrDWHOAiyJU5WWGYcdM745bHedoaphEifz2N7nQctiuATIEphP
E41q9CVQl3zqlpwjRANBnoCnM2Gk85Mto5vIOVt/mQ9TO18U+fF+D3h1lnMidsFf
m8OQoXMINO0qcU1me4EwKgE0Iez6zH90aEAvbUL6V3ZviOqv8rq62Z/zdfR8XVa6
NGxVhqBYSmJjBnpKJkTwmhmHUJkJLSETalC1BmNCmFfNJwn9LxLmuVNkyyXPcweD
E3UV4uCBO9GlhpoimZbm079hE8kbWxVOTFHp2eazwyiHfSyJTjpMbxAdNZwMSGKi
GBWxQxCjn6eqV/CVKL+Kn5o/YLmgeppUFuikI5gU0mTcbDju4Mrd4hJKtAAkuM39
rEJs5+qaLq8r1RJz1GSyBPZZMzE0TiVH+k0RNs4cBr4QmCfI5FotLlZ4FfDrtG8v
T5zpn9jhhk7fedFTqg2oiAaua4Wkd1ywx57FdOcJG5nyZtPimZFsW50sPRemcBRV
p1qGs9nzjBWh+h8QXwCm3wkSz2l8OJuY5dvvhfVxPRjboz4fgIqmy5XmrwUIQJGO
QmZEs9Fgl39s6Aoh/BT4GSIGL/Kt+vnZoYucMRDVAtmx5l2mfyNmhad7H8R7kS7U
bZSwu78bqknOdy5PJc0PM6ZG6kRPROuJXE9KC1e6mOak2p/nx+g0xWfbz00cSDK4
BG9eWJtJL0/WoC9PM4m2DmOEGiDz9i00g5BQo7xps+E1eA0VAHtDKruEH5RqM/7n
MiyBUZKy0IG0/jSvARFWwg35BEjmNqi+tAlDyyTB2+inzzzL3tx0lWfJtqmH3al1
PZtkMdtPJOM380arR3dkjdqCXE0P+nYBABolhruSxUgpGDtH9YYdpAJ/ilRY7qzT
cFM01oEmIxo3oeTOfDr57KbjQp+QZG0YTWR360uvLZ2/V+D1mYP8PrRQqAbyrTwH
Mf4OJk2ya2zuBNk8uhnGW1OH48CGeUsiM1/PokSjzqbNEXCxOwxGpwHlj1wPL1cF
eZSbk3Bbc5erEUFNk7yGLta54bSEyCZXwGOXPgD/kHMfCVIcUIKjHaUlRfNXScj7
UBaZsvXEsSTRXz+MDPGdNkcIpCZRd7oZuR0aJNRMCnERZL1DvoCenTVRHqJMpXZ8
U4u/WAsD6YIup8g75IZUaO6WDEYc7oTNV6nkv0PNbtmp/gb539itRNgiHGjUDzEm
Eb7Cg+JtOR7cqwOMft9j9zFsqxOs54wd2CQnwNl5Ze29y4YlXgBqv82Ykf352Zi1
R85sriYCVgOdwoBbILffxYXfZMmAYuCY9tcOhScGKycKVJwY5EOVWdt7CFogLKNt
+mlRCrjzryBe/5KC3gjyxeFxq+Q3JeAJED1Tb9wBw3QpTEZF2RgeSscZVRil36zP
sW3LNrUNpIdHKM5ssEqQP3Ng5kYtvqM/JJGo4P4Osi6YPnVAqmnlnnbnD9iyLsmc
WgxlnEIT26/PgNdOsW3Fzstsq351Qp8N05FltmY1qL1bYo3AYdDseojt6ZxW2Z6J
MWDMv2I5GRcX+Ovm+D03V81Ah4u5qT6Ha+5MTJjDsRi5hTHmJeHmYMAIACmR27iJ
SqrQHDNL8UNR42JL0tSvT96YxenB5bBHMwpe0okrEMnra/EfgeA8pdZYTSkFAbGl
6vIY8GDUFghfqid4dk/Bl73BpLUJdvHs5ilM1VH4k8khcJwR+kvhtKjaVf13e4II
OGSpI8NLl+QCyJV8cJiIqPxkCITVByKmEJrIhUGgMr1AZYoWMUU50r8wOOhV+XTx
cU3cfTp1EAA/g6Zu9Ue+OsDNedXFCdhXduA9amnbKbpTMcpSO/NsMqtHLQOk1+d8
YRTLUJ1Q9IYt9whV3aLI/y9aNdzI7hBifX0CgrCgfU5A0yjhu//68lcupFupgIfj
xuibgU3Adm00wOkRs8a5hlV/h0EmMKw6dSjHboCD9HOsWTq++0qVsjBi5WNOZVmt
GaaDUlkByvW7+LnhBmoSpAKlrcy92AxujBaxX5AY0s3zQyYUKOnni2H+DhHDnBhF
9dim2okHwvWxp2gx5Hr/mg2phihjPJdY5md7LBlJ8nfeHQ0N31tYIH/WPTiKENju
pb6RFNCAPtSpg1SUGFk/vEMa99oEEjWAQSs/YvpWHUxpFB9n9nb0CWEQ2jq6NpDX
74WIH9wsxwKONEbioUXjwwwpsmQyUCxGQfXuj2aCkJBce67EeN9R/GJiFxu2dQ2C
j2MEc5VebjZ7fYtmxPU7viMs/YVn88n6JH9wGzHdhsUnn5Zj72i3+EGjs2cvBM8R
Ou15EN7Ja4Os8ayDeLky5nP3AyTTE1q2lns3mxQe0+Bxm5ce1uDBoBF7uR1cmRJ3
uUdBXT57uZ1ljD+hSQ4YIAFza3IXt/Fmxc7b+5vSwv21ke6UNj6v5UA363uaJDSZ
JvIHgvYyn1WMwg289vbrR3uSm1p+D19lErgl/FnJb6HIYnQt8/q7T0r5zpo7/U1v
+sfmrNLERC+3TNE3Em7t1by/Fs+OVpteSRCvttniYk10rYvPbXm9wJdzNe/YAeCI
3xu4uDeojjCBzUcbko14Ytg0oRlNixlUlEZgR12Ycfrk4y1Nu91kHx/OptnNYV0T
Hb+zxZT2qgNGoZsJlff6NYTKjeSvrDrWucFLY3PsqA/pDmg//hZkhVXyOo/78G0I
Oo84XhmOFYgmgtaVA90wBRqrBVBhQrQ6vp2nNTqCkyzJgBd5XH3Gy0Ph3eriNTPo
LcOkBt6lHJVgJZvGfhJVbEF2LVnNAHOk1UG093gtrnH0YwnDBjLKo1FkBIJrbPsf
C+X1hTa5jVqwJrBSmfXLa2E1YjkKUtCxE/roDE+GeQKMYFWq3f5gZ6b1AeOQyUqn
17YKu+1Ck1eRimwAi51/aEoHEIFTPmVfi6OZtK5KSQv9qPXTsD3PmD/bJihj3nub
J5G38bF29wDbX++lFZ+/NWYBm7zN51/bNXT2jUK5lN56XHzabeRZn9pw/JMvZKtZ
U1EW13tSoow0PMdOtN+yjd5SoZ91tE+d8PVXW6p+iJTTmnrWYyE16H027YVT1ifx
FWPE7KgZfv8pYUCOkR/P7sAzqFSJT1I5aWOEZ9xAn0AIRv+c1JUKzg19eHhoc8Eq
i52bBW5kM4MUzHKGKR1zBp6O+EO0GSWbXL3mu+B15W5anK/0LOj29OqYxfArLOXn
E0sFaICMqmSiA8nZCI1Xou1iD04a3PFVKlB9QFNvfJw/mxRGRctZ8NNCnS1QhsaU
ier2Q8beJxl7GcwGXoEaDnU1xxuJFF5TxKIZhjD5nRWdHbuY/cjPXB6u15qYZRCT
zyRuO+pytye0PIF4/Z+lxCR5MhjUePAYZcxL0/tnH6pv9IrfkFODBezN71qKZxbv
I5NXn6jgARAjLSW7U32omms91M2IlqmqPcaElR/Ydrv5s9RhAc4uSDE75utB00tv
AO2i4Uo2C4Xa5flQl83df7noXzNYjmv3Efj8SiikE7sRlBrWtCDkLuToQZ1qwItw
ySUX8oObWf5K9R3UPm0KvRzTi7Hchu/CYLW1IiD+YiF5Tumb8do7HLcGJCoOrRW6
V7t97994t3vUPhEc9CQlvxrXyNSFZsgXdgcV58Y2FDJn38b8M9E25W7n9Px43uSl
lpZ6PRPk2XfSm+W+jDH3RmSkF/h4fgez4Akw5HdPR1hUOafSVPP67MMYZHZajn+y
RyejlqBtRmkqHo+hYfOkHwlIC6RXsI5zv8+myRn27X94PgPCR9zwzSWb1FD+k7dH
LpGcEykZcMur+OdeMfOSO8BsnOxczmv2UbKsdyG34GbvF/V2B6lpW5Y9yzxi5YK1
asuTcUXF3EbhDLw/e+F4FXhD0R2QDy2/wzcUpURrUoql+8cW47vCZtFnam6fzwuX
3sSlWZ79OECFCjYzcoH5pNvDNWiRTUOdTLgILRZ/yFDx+95wUQPs1J18gOx/jrpT
k5tqr7KwTWp2bkyydxf0mlpFfOaDPreQnAqfw9qelG6h4jjdoPNmvlWlR5grLt0e
c8dgLHlCwoIr80xHmqgdfDUcDCvR2e0hIV5MPdQEb8Jkma6oqR17x0xxDsPwOuSI
lOaJNv3aHwGjam1nY0LqgRdySzS9Dw1COxpIrPWlWUot1nYBV0Zpi8YuoHpjS7Mx
NCZInxN+he+H7rBRNjok4nKzVw8X9CxrKRCK+b5K6S9Fq50VpWVFMo0RP7LMR8R2
dAZOqsBObre7jX6kqfJe1y8RXuIt4P60fN4O8eRveRYpYjyCV13jHiJda65cz0qd
0/kZB+xUTy2LzUr8B7rnIZZkODBfYeaavEZ0BhLgdz6vXVs9fRUafZuRoKp9ReAk
3NuQ1zO8s4gP6P+qGiLke7drxTpP12Ltw4BjamxkxrkkFdHutfxjD8vL7XjMnMVs
FnUb/EGN1W2Dqm/HiJWiJb1X/RCZZaRgwslkgJXvjiVNiy+//1ByOYS+Ecet4W7r
GXXdDY6rKXOeRwvyQSzlG87OqKnu2xWr9cCuQ8kt5DpQ+4XJ4huBK/taqSS539qX
qQphk3/vJzxYa7K+/FAbNsSZjp6YBc4fl6vqxW/xdMRJM7vug7ilZzM4ClYC6Yih
YZJn5cIBdvFEru3OcYovGmqPEWrkdOckwICaNtdx1FWRyTMMYNSRGpF+VmK9c0ff
znpLsO2EgEqc09DlosX6Oy8RyzsIvI0b8O7rJ4wuvGtrZ1qkfd0n1XW7yI2dNKRx
sfuhJkEOrA3Es0ktuZnjhGfRNh42J9Ev1pf3zq3I/zZ7rOw8xwRRgJn7YTU8Vk/A
iWcl0U5G8LfsKckJMadaDU6/H6tROICIUwO9ACboAGVYTeMydzZQYkbmlrl1AbZl
tTbRKspQI38hkjlA4lHNR86mYnf8Aifx4lXNra/vg2MLSV2z8wdU8LsrHqYkSu9/
FKDZiBrnCDtB4/DukQsr7vKaIcLF/30skLHbnZReT2EqZOx0MqJbX4KfCPtwjBG8
uMayPoXCm9jHG3tRzy6myqRH/iHyRL/QJlebO+hzEUZOQ8hEedBjg1DD/klrc4Dd
msjJgniQ6xvTmFQ128zpafGzSPogrlYbz3hAWq6jaVaizNKjht7jH5rmGMOIGM7Y
6/2INqu7D9/JqiVntrrHxDmZFp4PqSAEWi8egX1bTKbDd8enrP4S5O+MgnvRCjuR
AJWNxD9wl7cY7cWByI46NO+4WDW1xD8nRK4DcqrwdgT9c2DPaaxGzMqaLwYVlgsB
lt14SZ3ZLyBY710cXd1LDAtUArousGAVWS4Ml2Zcit25+vJSBH0lRvw7ix/KkxWq
Q/DeAy/qscpEEnUuXcXSdu1V8mf/AiaP4L18HV0/kJulxwSaZvH55f5MtH4zwVls
JnABSW2NDdEtDMiXrXv5Y368g3uwkrAuMX9vB011OZInReaVRC9MO+/z51i7GLgx
7irUpDxKMdhBr1dqfxsDJT9x3w59wF+3eIFDaeALfCa5v2+trzVZDtV3GRE/zY3c
vw13efC4MgHQJEFjBuUEXClz6phxKEPnRGwIM1ZL6xx2PbYtcK5fMBUejwFUY+mv
YYjomlulC/AIKbtNeMg9emJLsOJtSRnrwWJyzYthWnrfsDXhk+hWu6RMvLMXSnM6
HYTA8ye04QeVmv5/2/jK+LMaTSwRqFq7kEj6njYKOvMITMGSM6JUWVn4k9bqvOFm
+62hT0btmpGfmhzoZVwywfnBbTN4X5Ido76gL5uXLGSY2sHtb6oITE1R1gIpBKzh
6mXuZBfMEm54dvkZbDIBF7zsaVsw0Q6fqSX5yj+ujiDhIiS+yqiwnFVN+OgcJJ8t
7wal5a8TSZWeWSkSf9oKCvEHfW7RU/z19ojix17MWm6rDT34BsonZKDApxE+19Cb
A5dhY27gDdOaGV71Kj4TyYMD1rSUqzX75Q4Ll8muQwWVM8w2QKbTVLk+ZwCpUU1y
2KIs6GvefTxvO1Cj75h6Y7WMTDM3osMA2JQseQFeqSQoeweSYZzlHID018iDvUfd
vI1VUqLo3UaX9laxOdzeBX6FRx9pkdPgmBlAu4x2WKOMVhNBgtfAw9gzlZYhJVC6
8so+bUZakzrdL3FlGJhlbtuqWwNaMsFgAmjBF6hM63vg4cxfwEQvnUoFsJd/qTcR
C3bA/3XZszDKfOHput9MWwY187AtgDvdA7v6RR6os15bQ1UXGzGPbG2PShu961KH
AWXNsrY3rQzyD16pWnr2dL9enCNxIkyUSiHlVVFYDgIRZGcWEomHZ5Lv140KCOgE
KEzB2NUgAiVcKiGblKs/jE3yOoTrvYSkcH0MwQHZ2jt5bzjFtmOOnRp/nBjkejRr
RzQXzcjwrTf/6dHtnrbjOPhZOUJaP42GTfcR7wyuGei7aXcRbKLOVree+eO9QLav
rTfSTW8JUspJEZwBLakhetLT7MlDgoRooAPFUU/KUe+nVArliGcvF0jqYk0S5MML
fv3Wxf+fNHmAIPI5pDAttNxhIpzqmAHte1OcW0uvXs8+RNG+bPkkG85dFHOOawWS
75gDc1izGagpP7JGdxbPS4JquRsiaq5mRt8j3L1lwgyTgZnEk4Vu4DvTLjYET7PL
28Hy4s30yaQ7NQ2FwWGXHzM56RRq/7GfLjNopFvxReseSXjJLhX2/xqq2QYPKFQH
rfo+JkG7Z5050mWCPdnYs5pSbK50ceItraBvnniBKlCLwv0+jBV/Xu7JLynD+cI1
6qF+/JGH78GI2vZW4B6JQVyvsF5sNU0F2Rr1j1bNF3roJndSn8AMpzSsqtZUcnFr
eBvQHQFFM6dSDFWN6QhbPguQLuPFv4AfcX5RBBLGQKoM4o0MJuwzRVCAdnoUyW3+
iMsIFy90cNTHMjhxzMPYZaDOgYSM6m8LLtxbKEqjtow/GZRVFpFyNfw2jmpmyqt/
lxQa17v3btugZXnIhf/qU9vJ7O8BVraMiHPHwTATVOgBCS38vjCls/2L5NkpMEQr
ThIXnC4+RnzdIm3ysMBvgRscLk1s4N7irnEHvF2pYpCLiAu6IJ2+8SAk8m3t8kim
v4pKwGaBpNpB3CQ+OSo6viaDwNFmlTFsEYZZEs9Sj8HX2V7r2kJeoEKgZu6CTaIA
4rynLLr14Qzpq5Koxkkt1yGXtqSWS9ej50Bcfor7X/RqA7L+afRYvF6VtVcAS5xI
YmtT434ViOUibPDuy3qhlmf3pMm2FVolqWySWwqCL/TlhuysXhhT9I2ylY1pE9uZ
I9qMwni3+FF+8J/JHOy6phMYmvfwbBOdWy7mLshzndFb022Kbe2Tj+IabjcDuYFi
9MOiVggXzYiitv0mL4JUhAJsTNdVvoWrjM4G0aSZDl00AX+oE2CWJsftb8lhVroz
9ungDHeUWOpzicMVwX2EQ5FZBSF5j3zh7Cz+O/UOb+8s1322ifiscDKiFPrAtECs
pCyCRq3M/AYRuagrELrx61Jlsd0XXnCriH0/VM8Sf6o0Tm/zEG0IQbXwBpQoJ+TT
My1xuDYOv3rUB/CBIgeS2kU0jRJrIjPpEtpqovrpS2UZJzejS1ZXqxVo3ZvV4wk+
cPua5412VjETTrCYDpk5FlT0Htr4UONgTV4k/anp8P0yWG1YhBsXHt6kFvQTC/vD
QcCQRr90dDn6j4LnPluZFLFU0Z+MdmB0aUKmK+C3kpbG2hnz8z7Rmg+hotFHw8Y8
QnP1fNiaYPGiDdhqtlTFCI+8W3F2QNZJ1VnKc5EV7sZUzgXBEfcQr+VQNJnxMxtT
j5wj7pDHR/TmC915Dt55MSwzWvMovBG+jlhpPlnc3YsZinZFnNZdnWi7SzP87OF8
KLhpjj218rNU34f+nI+BUuUU2FPqCgXGkLCmOROojyEm54lTPMvkL4hd3sjLu2xT
ZXPBrAAfvozDddgL5+4wJL+3ht5B22wnIhjmyLiScgdorHZUDFBpdGBaTWPvETw5
yUmMfJG3NMgHmNGERXa/is/E2bPTwe4tRdlxjJB7ArDIlnLKSlVQ7KRyEbeXzxAt
3DXcEvTI/RE9KWLDCaidogl4riBuRAKjJU8Jpu1Lbdgbn0ggUI81P8wV1GNJ0Iop
DxIjKsr/Uq6AoSOsDJxWI7efK7Dk9ZUU/bbRkg1J6D9VrGwSgJ5WlhWU9cI/zF5q
Nf5GDvrbsaVmoconEblOelFxtzf2Eo52n6ZG8yM6JXU2F9gyAk+FwFJOrrTVFrb8
Fg8bD/cH4Tx6Z4oL0YayHx5iC/3WOG7GDRtYV6sq9j/II9qubaD5GWT2bmj66IGu
nY6P5MwaTaVP35EzqU7mWhTU2MK/acB5nwGU6U5nhEZQqUbHhPsQyC+rBvA9wdXa
gUF5hj4yTeoQ7O6q8xCdriwBYt29xUi3pFwRq7gTiIZvOZXvnxvd063pF3bP6vFt
rvfW659iZXuVTViuky4O3yEBqhq7H1CepTKsxYukpg83SyISLWCz0vw29yAbdX2N
VGnYstbHJQWqqnSJlPpnpNAhiSZmT6yCspLG6PF1fpPioarAEdmodgDKOs9+Bxio
cI6CWdhyNTdU3Aw0Hok+0Qnw9+Lg5087NbQsxBJgDLos6HLEKu7HfYmnDGJ/HuAT
Tezao0mGgb5gL/Aja7mBM9EJLLQohxPEFypMbLB7HOm0IMNLLshOK9ycp3HZJsuP
omv5MV5rFJB7bS+lx898Ysl7858CS1gb46JywkNlZi8f/aXUAxhpkKDqgyhZ45Ig
mrbu7LmjBNop1snmGhPZpUy8thd7mLCH/qmiieLEM+Le1N0gU7ADAB6RUNxcA7OJ
SbzP/Qtl77Z9r7Xu1cIhgVrAY7wDBi8th0kOtBhqBZU3W0kC1E6f1+C3eDHt1VMS
kJcBUdA7zsHppDUJcPXVo2sqo3w/cL+J44tBhAcVQBY2j2vJusZC+umCE1vhRkKd
plKldcX/dC8h+xYyynpISBSa6QaxUsXrXZZTDeDi+kGGp2uuevn8rHT9jO2aPNHO
fRgENJDjqDVoKCcRgNTz2cCDcPca16OrWmcVGQ4x8cKF1VOoyALIHAiyS1Xu4iPN
/PRajefXsTUayi3ii8n8C1+IJaK880w1VEBwI2MzBUHmjDp2dlODRQKO1jSazA+J
a+GQmKSK7PCj0ZjGXE8ursY6DDzRGg3CVT6T0eeIsApu0z7tYPt7pd9TxLhlnNCh
HiW7eIQJ/kDpkCOh5cMb2IITLHt0dBS62xEGNgELXgyY/NZpZ9/8mJBH3ZzKTWVu
/Cc8L31Q4CwSVLX1CPxIWsqQw1tCkGVjf3gmax+6G+N+w706agc+s4/UL8HxHWhi
uUTsvDnXvqaOYetvCbFjEuobrObmHkWKbzDIGMntYpq+hN6wBboqXIIdom23MxKk
mwF5ImFNqXbdK260Vkm/qkKzJozJn0s2GfSfo4W/euGwo4oB9UhXkXmprDEQSvWC
vBkmd7X534xoK/AWQ0jWz6BQuqB0POZZGnPPjZKSHUbTZe/WKMTlFs4ZPn0BJf56
ybaorzWnjXxeDuzHJRcBYRWXh9r0svi0l9xsJuOowYJ9ae0mVHyvZMoDNw76KH00
K9/lCO12fvtDY4FE2PwZOJv2WoAc8S4rFCAgu3hRFLA5se1oa5y6R9w1QSYVA3L1
ALgGcn3AJO/RKS7bN0pm0BE29XlPEsn0OjbFRnB0Kv0jFNdkChe0Pf6Ho2WxO7U7
kGFTOwDDpqRUl3aoKAu+Fe5A9OGZhXPTNxtNOXzUbQXXsxSjo+03wg8jlYmIJWBG
NN9/vZZjCBD8BryIIyCpDGqU3JoQJhlPHy0F8dHZbvPd/2q50dA5RhienypvKQzi
IlN4Z7qeWdt9n45qEyYdmyhd+xXwNRH6ylxciuXRmBazLyn0ODIH2hVlnGANzEVp
k5sXX2X3moybMd79vB4w0IEj/VRZbnVJyzY5kzhtRJij+M4QbT4YZKAq1x7+1VYw
6yvEL5TU5pKCUd2eFksL31uieR4X0mofHOqv7+cl0ejU0U+QPRyKfXqrITHLB1uE
qLyNAyezriAKPel8qzI0uC+jb9Tp2oCmiWp7XyJfCF4Cr6iT6xXSPDp55OwWC7Z+
MYWdcSL9wDjSzFqOSOeLIPXkw/JAy+pbI9K3Bh2mBZXLR7O4JwKHeucyUPsSoFU7
zaoqp105bn2OEVaFyDKeP88vnzghioJpvF0WYECytHvo/lySjVM2/Jvro8rsdip5
tSNAs5fo+EsEFAKnpVxno1djQq7va2oP2nxiudWO9O0e2NUE/auJ09ojlj0S5W62
mzqXLpXZ06jYGS8tVRVtPwQ37g62ipLdlEGZ4+zK+nSK/dOnXM59i4hpZPUj3T3q
OjCGMbdV8htVi3Tst5p0NIj5ZEyqiFJrvQxJL17A1dTo+xHTLOFPJRwZvrKlJGsr
FWvSlqvHpM+/xzlRR4gVp1TkvCIqR1TXzGhfVjHejL4Yzx/72tuuL2+OE0bpaNvs
zaCUZQNqdA5XB3eyFvHoOatRA5XC+y+2W1OCBjjvS8up5lvDXe2M04d2Az118RWn
RoNCcYKHFdQENtH8U1q+Gpx356K0MQoieTPN8LNYFgo7+1DjLhH0bfaYqkSGplR7
mjDrLrw0xs/4kKgf8LMQPcq2Uy++RPcoqvJsnExXeioA30syUUAWYe+Y0ucxxTWc
4dYrc/ArNfFrq6IGey2zdBqn8q9brCODP6uaplA6FAX7gVhU+pxw4N1+rPyb3G1u
qpJNfx/E+tUp0pay5d+b9qr2eHWae3NAakmBq7kSz7k90sddJZyGoos/YZ+0CBw1
4h1FtlAJwsVyP7SXwVaTvDJxirdjp/B0uZqbr9ipPuqLck/TB2lfzYFLbi9y3F15
gmD3oYME2kGfzsbzbokbSQlKDK+HfA5qpso+1R6YKR9uaNtBr/UFVIWJVPfz3Hgx
tF6q+V1FqdTLf/9h7N2lrYogwVBhouDxlQLrp6AgMDSvJKSRvWLQ85P3aNRw+1K3
TXvq3YIRsfpwebrHdiOzvV0TAoZhSdC1iIQUuT3L124wcuM9dig5VSfFe7JNVGH4
NPJ8wAPmuos6giX1oJQHGnBDTCo/f5nqnjLkzJlrg6kN99SkXHq8lKqz7qC8U+Xj
YvPa80J5uEQCTKSurQxsC/WZ4LeXhQScD43uRdTLcDFJagoyjcs3yRb9UDyrkVSL
eRnUrqq9EWMMIqMZ6D4yUAZrVjSUBrWnha2QX3TbdYY+NrJmmyk9n+tUrOXxyD6G
7VPs0zziJxRfBaiJADY2mVPmJcFOzriBr0M0eqktgwPf1OIHtrJ79T2yFcJMzhc+
lgF3aEVIdu7ymGsXeD6kqAKl7LwvPWUXhThOyNa+sYyfLvcwOglxaQwUsse/+KcE
c6Q/S+3j357lKrGUyqm1N+OYcq5j9LhW1WKN0t8IDGkS29bBy7ykCef2vnypNV/v
rzTtD4izMZvbL6bzeZPA5cuTNjV9Boxu/97wYq4NaXKn0+cJ1wznSoqOzcEebTHq
YuK1NKtaPTmyI/VyBA7eb3C2vfOdoM5DRngR5c4aP9O6p0Csic6OlcOA5h74Q/8O
566p37K4HgRIfuIpoW9BU6P+W1je0K70OlLplNw2K9vawCUj8fIWA6EJBZgsNBiQ
dH4m9MHIvrKU0dO/K7zjSR1Ohf2T02WJhC+2W4P7qUh+NaZ2J0r8emFmhBMKcJKS
GhmAe0XyYBu5KCVyBk/07j66/VnFGogV44LchEPRzhQ66+0zUkMjtCPBSWaj/ViE
5um7zzRZpcKai9F9A7FfLJNdyr/LOZ9vfgVuRLoGht4AXgPAsUyChpT6s4Fih2bW
kTZO49JZ21S8PKlZvkAbvlVTAj/HGSylM51Dznh3Wi1Ga9UshJNXEVy8JM8NRMcD
KQjchIxmdEkgcGGsw0LsYlQRxbPeXwHKv3p7InvxDShDDLG+k+aVwF33pMOMikxh
ufap0AuQ6/jslQ6QDkrEW/57jdlwiZ146yuxtdHsPXa1Eqtz0WMzCDOgD4kG+aPJ
ghaBGM1ZobFADPX18GrOiuc0q9j6XYnf4nsVvOVQ9BUPQMGlRRu8hd71UofcbkGA
iqW6Lwb/6RWGAIMM0FdcNqo4cb+jLheMt3v1JVvGO5iJLa/zhKRvXk1wGaaG5r1I
xnWTorQ2m9Xi++Wr5yHKjZa+bZckjGiwMBU44vmj9+kCevbX9IEKoMnNMA5KjRM1
7BTizo7Cn/+Q3+OR3XlDYbPdzQV0xTI4csuUgqILuDhssmcxbW4LoQKbvs+NGCxt
FK+Rm4AUmd76FvoMJNdnNJtrbm4thRloPvSsVbCiha0JXZYHP0MDLktl5PTkrWL2
irO+yNdBu0PwNND/Gfz2ms7p2saxh1bhtYeFd6RxV/rRAiKIrFfc1S5Kxw//1aI/
LeX+YB2l/6wK6zJ665VPFBmSD6A42oTWnbSdu5lixr43TfqUltwCZceJzUZA9B+j
5XvhR/fLypwp23+naRe0DJxn7nqVi491em3PKnwGKQUN3d9CeRzeyk8gZhnxol5O
uMI0CrtX8BQaXCEHKL/A4F8yeELlsY/HK2ImHX8YalxzFJZv86ehElsh3b9JN/q4
CjTrOK3PcLGC5+9bRIooxiot1sKBOpmNtPnSUI5AHyO9LmrmnCiiaUbhaM9KM4B0
+/QgmfiEFBRIbyoi/rf4tq5BKBcE1dOywYKmpSWZOhYh7T/I3W5d+0DezVyWlGA/
oYt7S13RRyNRGIjxsGccrzvE7valWpriZMy4OuZB720FHtQfAaK/zV+Lfum0mxRV
PLiNVdSBGA2muiaAYUqvJjFMf5FQI7Z5kgOBCbL9am5gMZNDhB7/erIMBxRL1oKl
nvsbdwwf+y6AOyzX77kSRgFPeNY1e0bx6iMgxxnCS05ZXD1pT2sW9+9QJBpgEhVy
kWGlh0oZ5A1QDsp7sOndvZTmyPuGaa3DeYzyPYLL7elReCpBNqK8FK5dwzXZNQsM
VLWIxfNQTCEs6awqVS/ju8JCfbtMJIaFeHxk80xJeBt0wL3OBSgNJZIbEWtCMIFa
T/+FgWHUPLDxqlaQttrYZixNvfwwS8ahLaKTbXXKOoPX7gdzT23cnihgqXPlVymE
nceoLvp6uXn05WAs2YmkDBrLSiacJX5J38e4L8IWU9pCZPNOgqfqFUn1KToTHHbO
S4u0HuhWFeTnLbp42iGAg6hfYrJ/ZgVwVcvnjygYsJ/UgFfuuAVWD9TpsatJxi5x
04kqwMSfUR918mdN9noHnbwc6XKlASB3pwswhToI71YDE7rSc5vdhVlKIvXK+wBM
FBL1xCc/9BLwqdAQucjWkwJMhp3qulvhS43vC0nKnLd9AXDKerxJIq5K26qU47Jn
b7Q36hFRXzvoWrRH7NX+Gpq23SdhJObiGxnpQYuz7/ePts0IGIlRBYpGRMf3H62c
JqxZlMwx45BrNdJG/A6Z9uj7v42/9wY42JlESlThTNPUsQqhHiQOXz+OGtg8lZFL
6CZghEmM9N15veDMAWSkoNQUhX6o+8b9tsdi+ynUTEuFQq4t7QeSbj+n7AZ3tznC
P7UODbfFFtdXSaYyN5W3TCvMI9nqP3WtYWgqTuWItte2yaMVCWfBps3chpeoujaf
e0sKf7lKY/a+wBMy8Rqm9ohKuJJ8+59zQ1P8assLjAUfP9j19WsGxFGIfK9im9b5
sYTzmOTbdzU8InfiA9uEogiifSV5t37dESy+JlzahLC5aFzEc3ANEasK3RVToJwu
9ZZ4zP30k8C1vleb0CiizIJkFnrxFc8N1fimN+OLqLk9YVIVWWuF7zPWYm3rUKVl
DdJ/pLHLtMJXuYMuZk58/YIPLV5VsmQivugUSSbnhQfQTamAuYNk+9Lgh9nsO+aO
PR+ck+f7CEDGf3TssJIx7f5i8STn+36sLvHfeN2ACg8woY2ZjTBlZ1r0cuBIPRgh
Z9rTqyiAllsFt8CuHmpkp0JVa+RsYB6O6qyljRuC3wMrv8CukDX28395AkMfnfW1
2eF8FI0u4DB1SLyDlzgLd7362z4moRD8ObEKKVKjq8q39qrezK2QfegHLijhKcX/
PQcqfJKcwn5PANJx06q1StBpruhgRWx0HLtpDBGdw+j1hSb4jhEA3oKyQOabG94a
tB+tHfOuochOyZ6JKN7qeFcaMcaG20BY2C9LBiyj2LB1xHZM8QIJIZXt/mdDsDBE
Oq/SsPWB1SujICGzIymForvq7mn2GdzxSxQjlaS8Iiuj2kccPFJLPhRSdLnDWZh9
Ma331IfIzWBsnN42YcDMj6pI5Le1Ec07lhLHXQT/9fvMhkBKRVipnMQu6QIzWiL0
TeZX8+sG71OguVTAIQ0Ur7DS8UvJZiTjQUnT5e77sdww1faadQvf3x/3SCpeCwQz
3y6T4pf3tT1SMjNB9VOkxOKpmy58flyJ3Kdsv0Xau6xOWMsBvNKHhgyqOH8FwLdz
nAnGPzwzxxdy8SezPu1L/0TdHBuvPFbe+sS07PxAkVLSg2HcrDt+z3TNBtwqdEAc
VCvq7HreKWNkeCiAl0+0bEe0KViv8OLjweE5NlGBqzulrdL8li3VFsQe/nCssuPF
LYjrNayOco7pr3puxCKTzSjuQbOy634Xk0Xi5OOpyltJ0F4qANfwKhqO2GI6ZMt6
B5VPevZD8dA8FJLuVmwRmrNklge26jNBA/VVlhrkYYfrrQQLSQjjCSclM2J2nk7i
QoIi+7Nny3xeEm0H7VhWADLaLLidzbr2gsR1Buxyh2u+47TcW0VafkpuC6LsmO6E
iK26O3CX3p0yG9cVIXflLgCCrNscGYp+c/JlzACwfGaNWfCpDt30r+l0NDzfPIa9
LjLCy1Y6h4Bh7tiTXuqiSw4IhzaCCCXtqC4Tbwfd6H23a8qfrbxd1WtYIqYSXYNb
s6kxA32IJ+A6R0hM+YazaXBcM919/zOGwt4FCdutWQAJJhH1X272u7Nd3zjqqI1d
C63ou7ojymYGJA22Rc+HwqOvUVi8I3F5lqw4Y7yTm+BRPCz+MFS/1kXtq8UYVjX1
Mi9Bcs71NR46llvaFEpEw/7L1WTWEbtfdfGDhK/my65GYQnvLjXLAeqmBrbkUlEo
/wV7A/dWlJl0PTuN4Ek8aGN5JadLoKp85N9k1EvdYHqicRLJkO+G71P53zb6sbzH
EfhvrM8MCBzEG+Dc3da6Ie5Defgd3fgOjNxFVQvMMNAluGhjqXTl4w7x53Y6oz4V
iuE7OzorwxuMhhL7bM+aoqD+820t/pGnojLxTMLKQzTR/P06JRKD6+dzYkBJxrT8
pRPYl2XTproEqdrSk3rv6b69zoBHpOfHD2D1HRCQ/grNjuTwiClaiWpiTk6QeQKw
MhUdvM8wzfH26Q3AESB782Sszm1qtkE/mPqwE/ESxeAIGFe4VHb0ItIUAIoTYGH2
X26J0/7q8ZumlbbUKcyuTRmTQ/AtZufB6TLUXQvLH1vKq5S0a0aks90VMHjpIbXB
G+zVaAA/mOwsEfb13PfPp9uDUUGF+1BzLPyqPR1Sn9hfWQC9iLyC9X863CNDDviH
Di+E9x+jnlqANs0hr0C+HXHL+qMhyM/F42ri9LHF//+Gvpf/Ca2KxvuTWcnCR5Jd
Tsqgcc4N+YUzWr6fbLaaV+BemNkf4ik98r8t8z1qPMR/a72POEHXWuS1gO1a6LPw
O1qVVsYXvbFuU4QfyhhAlsA6NqFljHNZgv4Y4NUpf8uudg4y0TikgX1m0CUhZb7j
iimEY0D7HMxRQXZJfqjJE5OC+ykvLDQCFeThLknd2W0ZZjk084An3UWpPLtjhsNw
5daYSY0RSLritfgJxLLBSPMaR1tIbbReZjJZLu/fJw+bVxsg3VN1UxBIQpFintub
+jY5aLDGg9uZHL0+ew2c8PoRucsld7OuJKLQ6s1JnMZ4tYuEVGkukZAjUDU+3eL8
DJzGNGx0Dm8T43av4NwRK3/nvD3mJKwelZGFCd/+Uv2vSYdZ0HK2IFctq7PuqUHN
t5G4q+pn0Fa76nz2qxZPQqFbiVuYt0uAUVfUEr9z5AnKqJuf6S5nB/JR8cnLjpiW
LLQKpIvqn7uiPtX42jgd/2BW/AX9QeZwtsMXEGjJGet9ePHwTV89mJQcPsQlx9bD
m097iyOlWM+cFBFU1egoFnkGdVuOfCq3+O7pnvwftybiqU0Nx/FajjRrUPp1sXZd
O+1fTXyQThM5R+BtJgKtec++B3uaRMkUdfyeZF/2DsHjAJ7c+fEg2aGkrX0wTzlL
Vk4NIBnmBAvufrsNhIbrS1RjDsWiu60wFPjslv2Qfpnz447g5zioQoGvoJbDsbpt
4GW0+yJRYciL5u7ngQ0cI6EGFLzkE9eaJ6NXlv/6rlWtsnd6Qc268kj+aK1yw1hN
ID8fFU/r3Flg8zXxBicoZ38iFAQ+1Rtb6vE6T8c+LFGvtdZLtl5TWS5bwCasrdxZ
ZXQW0NtrviTXc6gmhsBQ8vVA7nEWtqD6WzvzcQARpnZ4nTPkdPevaWpFI3KEX6s9
gmX3197qOkwGAJtOgk4o48bWywKxh3G32inNVyyfS8YEY04YPyzImowhZ4vxnDA4
hesZW8WAUKN+JrR7nM+pAC5Q8OZN3CAXv+E0XwaqK5hk3xa3Y1HhJBXdI83JjNSF
qCXBhQBilTKoORWHVBN2AnH7gbT1s11hCl9oPxyKcf3boOQqBBRl3g6Z//CGKN1N
PkieGiZP1C0bgMMKusN76HGzEbRYFnYbHynherSR25wNMceYk3PpiGSTqbYtLehZ
qH9t3e1u0joL1OVEW8UidbNXwdUB80Yby5aB42I7QAH/xlXfJezUgS01KzSFz50j
4FKVhU15ti2HsrerUBXzAL2JKfW280A4UnS+GG8wUtt+YfKstGwlUsH9OtjTnEta
u4p6hRZtRY2cV41XpO6BGS+WkLP69z+Va43ZnXLWP9wsBA6L41pzhIpWA9P11WDb
STX5Hi4hMgF0J8b9pnTvoofe6qlx1KSPyaBCCPCLWJ7/h7+8pDnCOEK0GZQzeWqs
8k8/3NmIwoWe5sOMi433pmN8Fgsj98/I1gmOURJEYWmSI+OPA54qcaCKBGMitq9F
qZs6ZCewYbR5QaPaAyHndbdGnKu15137OFPJIzs/agoJfPCoprJB4vaY2wMpteDH
ZPiCuZ9sKvYDDob9DP1OaauNC7LFd43LgnnA98iTR9sDk2dE2kAT64flgOVFqNIo
7iUhOUcN0XC3PMWI41wRzUBtPFBXb+DzrR9C/C0AfJT/0XTpVialhmL26qBReyob
ZOlftE7O3ZVn7sj4+9UOAg2GEv83zJ2lxlnx8mogg7PyKlSKcbNx4gsOPSgMLxUw
KljDIo5fcPc4fQRhY/gUOCEyD95W87cMEkZxRAJAXfMWLBlLGjLdbT6CChKVrfMH
eCFT4ipQWaVD/Eq5AqVowxyHwezcGiXeTxhnV4iADDpyTH5p5tztBdOr0ohD6/5g
fwZsJht3h+GDn58kpCQyAwlBEsOv2WOdVpkKvKPQ6N6dCGfRYwemw08XSeVrXWjs
vZBm1Pat71boXK8I15WvefNLqL8aqL4uVxiRrIxBBVDvUdYvhWLg+p6zC5Mji6jF
maJZrq20xlS3Xb/CSG6/sWuYNOqdcWiPCJBk5+j+DUp47alX3RPkNsC1lKFDxf8y
6bRDzKHjHRkf3dt/RuOcj/weqAiNDz5Yue6X1YSNLrvhm9CQLmjwf92Te0OY5Tx4
BhdZh3qKgELdYrjwsgompJ7sYRk9gpo2SfG2A+2mQrLOECV0U5Hh8bFjAsX3QNuu
Guv4pTruzV0rP+K6oR7QP72b9noVesQEEOQrFRgo00up0PURacTo4i7Lv1+c8trE
e/gpZTGGA6Fh/mQ9i3D8RfpCoJ2lZiB5byIw4X5Y1HmwxOctz3T8fsL+BBARcyIA
86tKZVVFTlOG0WpAuSjk1t997Wg8AmZBQY97in3ey3rf/xPEA7o/DlGHPneOOLLs
a25+ajNZn+H6sN6Uk+VfnRABrGx7ybEzBUvMa66Z+er2sDw/+q276hyXdGtErYQH
vW3wCDu6rWKrpTt1udLbofe95nZdQEvpgYDEkAZrAICjXeYm5PK+lNnGFk63IR/Z
hoecHFnhBdAwDe62Fzx71Whdym2jXXe6qDz6pgW6iIQP/eDTRQ2h2aur50XD35cI
HP0HsKIPvl6W2nV7Kpth314eKt5oTz7ZcnNKpwExEiL2U2V5zRMwbv0zM0RCX20h
x98VP8KUh/YVY/grKs++OpeZnyyKJtoiq/iHDwGc6fIuF0VUDL04ThXvfH1mOBZM
ZaC9yIWE2Iu3sj7anS5YSsw2CmKsLzSUBqjhAprYP9yJ9U+WMyC/jFBVT2uZyzM5
jk+OoZgx+ke0V46uY6V/ueDmT1y6RKrfZprtpphXZkNiiXB7SEXNqdonX4pWK29e
BLkA+etVzUiHegfKShyRw79POyzKhr7E5WbNNN6hYfYHj/Af3i0a0NVKRTwGBwkc
JRsYEkK2P8gKwh4liCKk8Fl7af4pRVtEY92V7gkTLQ3Xxk8r0uhKeXmKM/14jLpl
LnRLoTbOnlQd7zsDjWTLX1ok5Om4fbF8MCMKj/JQZxgX0Pv7VBMKneBOqgM+Zx+4
DPjJkwBY3mv+9ctpdInhTsoGcfQYn+RdXZwt5FBal0Mo3WvmzP/EuQVq/ljsM7S7
2Buys0eWr2WsPPUk7di/R+ux7N4pBwLj+H10JaDZeCluTYBR0w1WH+Dst9jvuFUQ
QbdAcRpVH7hQFWCgou6iGFr55cNHnTrC0PBrrO6D4o+0E1TCxpXMAsQFc+6gMplJ
GAQXdb8TbzbqOpyHQ7PexKa5XMr2PPerskLxWsBlOynOrDMR4Wr9udXXtzTKOrdy
dj61INE5/SpYQCZUTS/ex+oxfkqEdVjV0bXdvjM75m/eafSoTpFxh9EQ8IetyBj+
dY0iFXEcj4AGD5qLDP8s1JTGYoXVH8JC6usL/YbtVpzoano5JrLzYr3pjKt8/kEH
mp8Eqn3NWsMT9W10brUp7QrUwr8HiN0ASPO1bzf51VrsVHaJAWXtAWwaJ09B69cu
UeBtRR3vgMXt+eFakVDXj8hLYHJ3TuHUxHNLduE90inWT750zHV8nPraql09axSl
H7YvW0cTGvHdgtihnaxjIX6ruVZ7AyvTzmF8D24xYlC8dGuT+6fWl18wFwLkkr9H
aPy3KBkyjGrIwoiPD9kWugfGypt8b7gSiScdyoQ6tXp0PQ5NXXeXvWNhfsEaD7JP
cVS7VL1U8W9kekUfiGI4DtpyeF7Hgpder6a3UtccaK89mvOS0wRBnj1r7d03tnVx
2RKUYsWa5VD2mbBoLzCSXqDXOBS9fljTccjSMdXY0fkS3PQ51Wx6wjNz8fzwWl/X
sNUuPbEghQ/9d8lwkpPQo+Qk/IysetpxJP3Bf/dv9kLMT9os5y6I4d1Wvsn1GPc6
X2919vWAxT2c9k4+iYS1x/w/ZtpydeSBGOof3YAGpEYNPMX4ccGxvTPBIngKmVY5
Yrp03+gVtgjobVZZvlmOfK/S7C51zDY/r6aKruZanoRKkSqL3tx6jCWBEGnFSDq9
ttb5mMKmeZf/oLPl1bIsHTX+6pN8CCW3jhLpnv3kjmrcXsOqPnTZHmI63cJ2jL+J
1+ZO2ta25Qpc9pRbZiA0GBdmKNE1c2ZG/12Gs0nI491WI7wmeJliImbSIAkeIWCf
oD0Gt8wIGrHzHUN7vwvdrMIyeIg+Si2SEngRx2Kc77cl596HjDA2QR4FvIrhhmqy
9L0XrOoMRajmkslpOvSD10g/VyZXhR+HXMnnzAxSeMckWv0x3knCQZuxapzTuWxG
4OHC6deASNBFqKoI+Pvhb3LGAvxPxVrcGxLRSyS4YKv7FAH0Dm8i9yW0ubZlX8FY
lFicvicB4+zGhVs9YSuIqWzAJHd1pIpBr8jkZjgn8JUyENoWmLVC7dUjbMyxU1hI
TDsro7PduDoBBNELK0vEuOmUUsLn8D+rfJ5X1QVbwLKE1ZQG74KuBFh7vntXK6RW
oO3vLl/N4Bv5jySHDTlTtEBIdgpNqUuQCwe2PZmOsbbKHOG1GFF6EVVYBP2wV1js
BPNeFpLFmqoltg0JxX30HVVaSV4HNva6JTtyIvsFBcox11jVylPzHwBuPRM06u50
B/ZRMX3EN1zwOfOJ0Gz/dxmE4TT8aargFk5gYbBdDLH8RN44Rrs+v2YhcdV9GAW8
BQgs7sF6cpR/n/AJCKrLdB3sJg0WJ/6n3GVfw3rt7kj3AAmzl+RJFgD1OKzNge1l
PGtsYjlykRkwmVYCj924VIWbDo8qijzeOiMfWab82hR0Dx4P0mqxTH9wy6swZrQn
Xc5aNkilAYfzxxcPRV2r7bmPHia5vR6y0a/bllDwZNIcbV5xFLsWxAgMf7HuF7Z1
5IntT0f+Wqj/Pz05ILhYhDUgtLbWf6XyDIZeG80oXV4u5Kuz3aWEkjY8mJzU7cXU
FAzXCS1ffSlIdmLg+J4UtScOiZDxPH9tBENiE/g6wMsOSeSbxHHPRT/vaVWbCuoT
TK88vIuZcAlyptZ1Z1e/OJY9aTPIdbJqByoQE2z9w5liwLNBSSt2jS3BvoUuP/w6
yd5zqQouNKbGIa1ZgoOWvKu8OdHKDWfNbptCtNFgIX94GVAyNn+0sA3U+uFy2R9J
G4ribriWJR05uBmA5mJAgXGRNNB1HYkxCNDExf0+SS9c5GBpNtorOBocGM5Z24gf
3gHzHb4sM22iSID/LjqWHjFpXxYdrBkrS4ve2VFyWV8H+cAOSUxP/Bf8ZkDiY1mK
84QXEFBuUu/zocPM7TcP88qs22iW7AEogYYfetvxFT3+jBRJFtADyTu343gaVG6N
23gVm0Ckd1Qm5VDJcMkxRdrGrfImtbcbL6Lg2NgR1Spk6UR0wgoKc0k9zKEop3/B
YokXxK2X2zqQQoDQ8zQ15c32qzjYP7cUy+H9Ga9DaFUdnyJ5rQTjZeKrnGbwVv6g
qVbzlqUCIVu0qUrMPDlZUQ/SZ+iv5uWTrs5a2aI4TmcKDp4PrtpYisvKXHQfimQY
JnQ/ZJBU/eQBTRQAYZM9cOIWu5kZiLzdb7vrnJh7BsUD1lrVBp7nfiFD5UX0r90x
gSfj+kZp7M056Y0a4qfdQqzWy96HlDDbrLR0uQDLZb1TG4nx4PfLx9QsFneehS5z
1mrXTtOZS1bKiVOtrCFj/GKHT9IzS48e3a3Lxt4MGkMA9N0AmG6pBaN6PFe2LPQa
jFKON23h68PV7CttAVJ7+X+7h8TItNPElCktIO/oXX29ToVQW1ZQev7XzBjkF1fm
iyxht7AbYL7WcGJAOBrt5oq3DK9xIQWrjEqoDfzt9d8B1BrleBurkXfZUFZuYkEM
2eyixSli+sDwfIt3phvAhWV1QNQyAS2UtfZjMDN8LgMfaEOLDyKIrH1+Bx7qFhrB
puBfsh3qTYdfD05OmiuRvqucmrIkG4allTXBY1Ik9l7bQ/3wd4JowlluQXL+ojj6
EISIBO6OeKqSoSSha4Xq3QbierrMctUb+ZfJPmZ/ZQnYgy1Jo417Xr0UetQLgG/H
TADssKLZkwHfSkUeOEhnUdCMAuh0UMkKm3dkutoL+/WqUWTsvDNB2mQQRqa2RdMN
muqbswp/UJnDFb57jCcW241bgWDO4BsOD7apBjxT3VvvdvbqBvSzmBRRYXuVZURM
03taXbR1Sr8qMAlh/YhimmVScj6OoTjgMrJ0PwlA7uUalvE5X+f0ZrOViq4sjT2y
z/axbLO797jhj3DER2vFfScBh6NFV0NdN6aQawSIMj3Ej4gRHb5yFCv+vZCOAPaX
4RK72zYubaCtO82J9iKyfDIPCN7DniMqfSZACaaYdDR5MjL1LPT0a/vhdfOuvMDU
Q7828TERdGpHHdIX47IDoz5tK/t3LdIV9IXa2eB98aWI1yPncXtcpntlq6Gvn46Y
nV/Re3oqCU2j8ZzleGaXzywat+NMQhW/hVAQ5rq5IPg79HsugI4lHhKJmsEp6s4s
DKrp14wggYc8N5BZ6ffYkYbIiNO7eaSgHYZifOgC/lMEy55zjOx06Cb21Iy4oOzN
AMhf3hS/mq6+qdDj0vHVIDcf8fqjxsbRXR9GlEVvTvHDfhg8BfABA6tLLEbDcRN0
8Q+6oTfX2oXb6aMfAKvFPhZevr3Sw7YKoUpqcCeNIlrGKhPj0nEYNOAc7Amvskcx
Jh8irERP524GW47AEmqkz4FngqwJhHYHABwoe8+4oN0bke/Q6oFLcpv2A98H5Sq5
roNp87nUUU2uT3xYjSQ7Fhkl34Utq4Z+UYchzvqO3Z8mvIITmGzXG/Klvubpb1rB
eIzICiPbIpzfUWtrK7AOyRiciiQuhlqIYp6JNDfLsT5YsPkMch+cymg36zHgVHYs
oWM84n+bAP0QViLeXFTPQ8rrj/cjngpdza+CmfMSJsC9SHBc7z1j2bJfoqv9j5mT
zAhfzGCVuvO4m/w7iNo1oHHqZBsf7bIijyUf1uLmvxW41CrLpLKDlOWr3fjTWKPI
5Iz9xN20ZruRuMnrT0j0wRNg9ofLvXLDlqyqatGQ59mtjtGC6DY6NFDom9L1NpGz
U1g8jWYqSCox3mJURNQKp3ai07dvngFfXmT+bjNdgyQ4cSJk5HBpkgbb60xZILIa
YLr/LqQl4mNE1XWxHKIJHa8Zr3rJDKQB4/IeUtiWRXBflaAf1LpGRdaie+8VXkXS
/l8XcN8egZDuwgky0Wmfzz1G7qFHJXczEdsFWDKzKnjvI/HeQWuHXtW9/2V4reu3
+LwGMlfrj/9sPm65YU0OQj4xMSt+hOPDW74J0BlJSmGvEjhmZKhl73ZsywmacwIM
mOuZMnyY2RTd8OCoYOJRFCOfd7rZgQ/l1llX+BuKWUXuS18oRaC+z9NDAiEQ4qa0
OtCeRf58WqbZpiTXzpq3LtRTFHGypPi64cQ1d+/m1SQkMVvDKjGTKMN12C8GtpNI
yU+dMlE7OVFQHN7bXhlFOfYZKP12IELc0RAhkAbMRTKXVuH0QtcLiLvlxklGTeZl
B93J4LNY4Xs+Jx6vO7O4AITo3OENzzE9Zf0ahTrR+Bzo6oCXAtrnuaoRbeAEWK2L
jrPvHj0C5zpITPc+8zvQ2BAiyhb9OTbRvu603PcT4RnnjJ0xJoBlGgbqyZYqZbK5
7ELTQyE1AaZX7ik3kxEt0mFhpkyHIzBCgtF6+GDg4O3kCAg22to39eVTzNoxaxFR
gJpgvtRu79kfIawngytgWWdFP4lTA7Spim7rdxv2jDfNkRVF6+J17EMuNRWGM3dd
Z+fuQQNDCYgn7Hb9bq74shodtoNkd4eF+pyPEn3wOUDzcurafArhzRykAzp5dH9N
PyeqR5v3oj+ZEE8r+RhhEzgz6ZOUSIvD2BYgizDvuB+TkDL51CbO2QM6VHTj/tle
5baO8nGNSs8cEFbZ9P/OZVKMOzcvjT8n3IfNoRhOwyDbpoF+GWYpTwDZYgKo0C9J
BxWlH2ZzfBnsivCH44RWBJgX6e0sPTv7u7fOBTWfQtIyByC3OczTzMKjK2lIXcc4
i8AsOQAwVHrF8kmxuYwBGCZ0izpOJklib3btWaH9wxVG8dbTCs489Im71KnPCljI
ONcOt0wGkMBtyqCL6t2OyXBSlqFIajmPC+N2UJCq8/GW0PHnTOMsXRcpgeD2Mce7
5J5S2bnGteU2/aIOz6raY+uUT9toNn9cuoL7Z/wEvaOWFfrKDtzVJE8rmMVdVOGW
ndoKQS+d0o0HRHY+9NBuBZLTTKCs+R3UkICYm3k6lm6c89bJmBqThzzINTZdiL+D
SaZ+cZ/+dXg2Bl9fyIUlaAL0JbTlUFNdpG+g68ZAAwCbuzGiAuiUE0TBrpJ4j3dU
lJCsj2HzMHa9inYKukfEA+Xrukwm1fkBbEkGNB3EO+mwVNCYisvCcyUcEwUwrefc
t7CFT6moTamRpdk+njBRKPkuOZQbRFwCxluiQgzYIzv1wDZfM3S+kQL1x5pY+5l7
ssT/dMYkaWK1I+w1cSqVLiVPkqc/gaAPB9T8NzHLXbDkJMdJMcqfNGoOeIbib4z5
tC/sp+v4hRtBSwfNzGZxzJEU7jN1OxbRvf1q7P9e8lONwOmltMJQXhP9Z/Fi2Rm0
Vjad3/v4W5yqCPFbpL+s7higfAPVckQrFGvQ5jCzhd9XJbagbS9MAZets73NDoYz
A0zu/ijcQbFjXCRqvjCiRUwSs6OEEW7aa6SPEJzbAq4Wn75kErdUlD4MBfQlCtvN
71775wKkWTtzexekyJne1NtBxNBPehtSSJiomiPhTxub1s5tanhIjL23ROk7wnNF
WXGp9//zki+eMi7x9lAC2E3B90NnfgxRD0WYgsvjDH/WUleUaNfqA2A9IDa9eJLt
gm6wZhgeEoM56sCetNosVXjAFVXMe6SV5vnNPX86zMvWBQrswFoN/EoQeoOg70Rz
1lqU7mqw6sCGPfDYIDw+VHypczJqo+1C0BDKSC21lAgJCHZNX4MofF41R9/jWHIw
wK4UokaPItlrRgnoCOMbeZInZqxkZcRF8srtALnsNyFee0JHgFuyV27xYwOHnqo1
dQRURHnZJyd3lpvsYEqI802AYqWyzjFuv4TaUBRZyK56davaBlMM3PyQPS9WDJIj
IsHlIlu8mGV9xVzD6TX7qqlJTKafI8PENLwGxQ9ylKXYFBWvEvkTadzeEh6aGP/N
VQtshpDd1cXELYvyLcHe2QqGxdm7J5Rf8SEQuLFsU/x+2seSKJ/zhCRdglff8cTO
JajmeWvsVhsGAPaHFbqbD+kcF6c1dEOBkGYXmGrwEpW5H0PLwVr6Lo4Ou5axpi62
MJqN37lNj/ZXfDtZY9O3QJe6KpqYFHFI6BwmV0tjWHYdY1jdOdrWEQ+NaNSlZLxQ
y+YGK7lDR4A9gJu4MB6XDJ77S1dHEifK5e0voa2gGEdEmoVuTTgZBpDLt/Djqm9K
Zv3P34igmN/rF5I1Q6LN8kqkMX2eBHLOorR1x68n2/rtzwcRwUcTx2yYx5sZNI8M
TELDa2IxPz+h0dGTDaTLXugw4kGQLvw2+Xdw0oRfFgE49D6R3E+pABc98rqMsKwG
UJS75uhqX5gnyhrMIv93g+p95NQbsagVT4fSYP0sb4KLV+YNRfpymDzsyfMvUxje
DxkVwp9I1OFebb0mwGgetimkiQDR+iThPPcCDn5JDQhjIxhz6kUM8jjzR1Tk14+V
JvyYmR5krmbLiJ4VG/7D2kAhiTJ8odaRsQAREDydRayXKP344VkoYJeYKORxbYMT
MZBdUE8/qQkuNak3znoYio5XIxPVACJCyEmSigWrjOokyz9nA7nX2eNsidKoOXK+
dJDGHLBKpH/5eHESD7IuelbC2DyXa7TByYI+WQt6DtEqSeAj1FXdJhUVQddq+I2H
/Maad5BTzO09AN6ecGVmx+xC13ZdzNZTxBv5mnxl2aKGR8xPWoqDGg+n03/nXGRt
QDMzfyjBJKX9fkUn8kFdH7vm3mPvHFg6v50GcpbCQIBWyPSX9G5ErGIcL6O2v2yw
bgfHa0WpkXNtqWN5y5hMxlp2GeM0koeV+1ZKuR1BkWJBHwvCmu9TSW2AlDldj6eR
Ckng0TIePGQdfjWYnsciBV8sjX90/k1w933xCvJtL/6lFOtwQK52tcpwndlHb0+p
jslefe7zk4NY7lxlk5FiBndbCBHeCj1tabkOOn94fbpn+wfbwaNjPW4IQ+WFg5Ox
vSbAgMLwHfEU5L92AFfP9nzuoN62oo+uDOXYRSb8OrvuQ8N3sVtKcEJ5RlU98gnn
UuJU/uzbG6/ewN+GPFNcfZLVlAL2zbtkU1aSmuoco3nN1SXoDGYbsmdYwmn7d9x7
fjKY4YQI8bUkAa9S2Dxt2sw4HDrcfwpIJ5rCYuUsLbF7wJVqXa9O/v6vcLJX24pN
Je7hg9yMMa1xhxyD4AcZHZcfUv8hhUZD4AQz63innI5KvKGUMPCCIktWU+jJ94G/
RQ4eaJZ9vnxatAh88aigArP4IPOwbA4Jdd2bFzOyP/kJueyQ7Q9JS4ET501Ju+1G
O3fAWSIdeQNJvncduSgTv5Zx2NzrYKSJDBBJZycld/IJWZsss3vvbLoDdLdq++7/
lDc/mxVoJlh/5bSCjOiDlAHlZs+Tyo8UxzjbvHNbV8ptdhZaJ8Y41WlJ4nfIMwVp
6mMn4xCCZHJg2eazWnoT4KYvAz2w4TqM8D5gBxqE0bJQnSdZ+wucYeWR+64kVLzo
qjo7aUua+/0D5bnYEkIzhRmEuQwlCMXxQqxWsOSbgvsd/S38dNqniHuOqsxmwCCk
QsZqKwHYs6lQEBsWDLFNoneDlGN8MnsZg5Vn+dr38yaML3/N/3bQ/pZ1fS0M96HZ
KEui3NSJmd4ITHjTVOTgJJZ6AbsC2rpOvttGlTsuEdgtJ2pmAqqcqD5/G4fUcVB7
pH6hMCzOuKiz3Ehd3NfhFlggtnzD4UdPclk+9LCpUX84/B2ES4g+c9Sn0AghNs7m
90oZY2Tw2drbP/Bjqa7AmvoLmhIWkVor/Lhe3EezUHnKh191kDfnEwNtl4RMosls
b6hr/Y4HmI9wxDI9usBjxtz4KukoOprlsJqS/T65Uv+jI1p7Qj98916KNeD3reHu
fWyi6m8nO0hBYlA+Du4xup/8THtY17dU8Ppv1GEQN5p0rhx6dF/MMl24ZyVB2QkO
sJXXlNNyLwoBaOL4qV+z638aPpnQbuhjHfXsGpQFRPK/FXX3l1xBX//O1ypc54yy
lDCz50OVZ/0tq2jXcYPgTElXMyKjhsjoylMxi5s2+Nu3Swna5bnt6siBhObGhL+m
DdJlRroYgSxvWKjeOxD6LCLPquY0mPzEoq4uSHUk7xuY5ZoBdDfYIDRjd45Me6UK
Ci/6AtOayzY3SywSgvq6T2koDjAJ8Qu2uvZvW6JWGqLempMzi8Lh9Ol3QLI/8j1m
vz7yZ+dKra3bqe9EQlKG+ES4ayGxBhMOxWjXLD4InD5DwIgdymLNnLJugKJkL1Ut
877EAqWyiU64HPGQZZ0NXlxarflKe0vM4Fehrz3byNrCcBy1ZwvT5Zt5Uo6mklR7
NJoCJHvsGebxYT1VZ5lSbaaL1rIdiwJq52QGoErOQIEy4uYwxCIr9tmlvqB1MnYy
5KVSiV3cttJw9CqG8pgr1Pb5xUbNu6Ud9pciuBIVuRpNNKGkOwjF7Yz83606s6zb
jKQuqhX07Xlv8BRQowXQ0Uhma3nFP9ciIPFxnORSEWg5Qo+6BanfpEjOQEG++TzD
tkXO2G7cNCMUgFlAIODWoh3lYdWnU2Llyhv21iws4olvkpvuXIPSeD6QZQLfJMR6
p38A9BNLBSL0mp+or8MtskTJaQxlk5X8jV+pbAv6dVCYv5HujZRb4/+Ms+ZMS6zc
B3jCSQgIM/FLlrIYAJhv38ZkxJWj2irBrk9rzPq0kq1cJqK7q4ZhTg16ZZ39SCJD
bpuFULwgjgwUf+VCrYZuvKizUaDWIHh8Cb8QbmWWh1yLJXGJ545+oLzGbLbRUeCh
7BUse4mSHsFoHLL17X/Jxv05l7qwn7hTFDM/t9mZTHxIUC4UCSyDjNcEE0hwNSGE
Qjjew26y0hK9JWVT1WG/aQ8+V7JRwTfsGKOyx5TPzdAltnWn8ATVQPmZPCq30Y4h
qIWJVxGp3Ie+Z5t0BZx6JnviKtMOvp87ZhtOudxRQuh01wXPd4q7qW7NgCWxaj+3
WiTj1y1DPGAuYrX0ZMqJ0rRelDHWFt4mxUd/IgWPrKiocrJqWRdfMKtLMcXVqB3c
XUfubXbNz6rICk19jcJNy1phuL7sltRLSxWVlkxwwrXCcoi/kO9QzTtGGeytNCnI
hzNacTmInTlau5GL7ikpM8+hdFVM/PiM9ItXOsw9RlHAb4eoELvORKXK566yw6X4
Xnoz6oknXTZ2jVulq2PR5pOW/+0ms5VkeEJSGA2GEMj8AHABlIn9sVKSU/pCc1XQ
hgIbNmjqR2uri+wzvr/qMeCHi3BPrMb/MM4me4xnEd7mPoyWeYmlAo+OaNAq0BpA
3MS7RKUhySS1QHZkXFcdLQvQnHL4SU7tBt+UUb9BRc29rHiM+Rgf4VtEpWCa5vlI
EFXHVPurLCHbWG0L4y3E/w37DiTIYoDUU6BcdBmzxjfJvIh0JrAWJnz3RPoK820O
BaTmeJ4i4dSExXCc9l8gpiIYMNJamxbiVrPphNbLdegPfGJdS1cb007FarKY/Lzg
zbQKRT93l5rcW40zJ6d2awPsDFam67yJIUYFJWZUlCjsUYomcsz/aH1LKTCj5CTo
/XTRq3Re+tDB/YcxWOBjEg3Bo4wO8x/AvbiB2HYpjDFmaSGCWcE5EwCAbhX8Lrxn
IfFq3x6qLkx7inCzUfcnWXCHN234eppvzuWEjvOuNRXouEE8K82XTTcd1mrJLNhg
bTV7Rle2xA9tOy5syeRajXFibCGtMPqpXBbLlxP/i+/xXr2kpamkjCsKcdu/CloL
RinPqu7v+5okGc2PulwYqHlam+FNngMMfCQd0KHl8xBOeddfEvETff32YoI3y3iL
MhrhVgqhFcf8jFthOg957LT65ctOeeJWx5feh1CvT2B6LFKXo91XI9QkHmbbQtfm
S5eJVm+LLx3Wdlmlu2jX+RFnKUUjq4hS+72z3fU2fYJ0bdQfFZLDn3dOWkjv32+M
pv7rky8ej1bPyD+Hy5xPKOkOf8SwJdZdHJzFrHNRtUKIBBpNakaSxNVwlsxlrodl
h3lKG+Y54qrdllIxZns4oHjNSVpuFM4O8RDOND0PWVP4s3O4O+gKrHlQ6nb7KcgU
DZppkBUTAFevXaN0T33zk57NTVEPNvxJS9F5vsh9CDmjhQ6t9PoguznGUS7iscy3
ONSe6voRHlM21eP1eHLpCTysy4zhzYsppr2GTypMiGj8H052z/5Z6GdW1oweb76y
Sygb9NAG7u0p1RlHspkmELkfejJZzMraOFGG+pZybPT3lc5Cr0DXjS5wir2CDFAG
jF9Mg88Qzuv6k6TIU6uOu6x/LpvqLbCmL4MzPJPS7x/8116chiAFmotAmv7NO1yT
AKRZxI+INsp73Ccr3Af/OuudUtsd/bfIpuq5k86UbFy3x7T3JmIbcIVPLgIcX2VA
GRvSZNgsgSKdpKFIm+uInZswMU41dYiVLt6Y0op4g72EfSIMeJBKy/itoj4IXnaj
Bj3qwgCvHyra7lcglPDjrtdBjNISbVLqfQjlZR6abiaFrieJExa5z1WeqtqJsNE0
bcPmlfllnTBtT2y2Zdcgmlq+/ZNzsdVRW1CuidREzRgdiMewmEcNPHse+trp7wYP
+o6Bs/pP1FpR+/jAlLq5GPPxLsHsHLTbw8IXtB1BV3sSddUMjx5K/DrTHi452dtT
caR/tUELNoOdEW6vgif0IX05wE3mamEdUgyEn2RH2Vrhz03TQqHO8M+acgJ9QMUA
ynSU55uS+rAa3ufKR0gNvoW4Rp5YEJzPmNnoNP9Hx5zxSQA6lds0I3W7FQ9JrTs0
w/2sCFbW013wiTTuI8Mu+nvyZT02t/KnKUAvypEIfKAOjQ1d28laBj4ci9+lZeIw
vG+Uie01y12PvApQwdqjaBlgVLxorpj+D3o2UcGN51MbXnD/zmkwRTaxD745M110
Q6W5uD+uZctIdFS6ce4o+fyl3SYrPYb9MOFuXUMSQu8+eWrY31hx5lUprfVg5jxO
oy78YxxUnrlZlfU0QvrNQOMSpxUHNAmhK+y2YIyQRmjx4U75lcfdauicQ1iPe1om
ZVuncPkwy/VDp0szDK2GYp2ihPzLB7CDapbu4hwk/3AiH0smBtHDvnbxnhoqnsid
cQuZN6+BA1Hk++XNxpwv7yeQXXXN30WdqAyIB6+8/f2OPgLTuiwEj9qu3IyHRUVd
NUOPwHi46uFaGGF8iCftce7rwCVuF+xBs8RC9qfjkRfan/GSDlThlsLqiyNscj/y
sv4eMvDVZL1AFL6uHN0MFLGUtNB4n6t/zRkPH70ns+etN6yqt6HIrkDvaz89p28I
Lgb9GeBg1vZcC5RCmJo2E1Ma/EiIhOYZJihqX8d4bSh+bY9NzTaIqIXrf8T3vpwm
ihntZgszwKXR7kree/ADWTs9FPe0XDMc174HwPQCWZuzn5MJxNBt/0oXLkgofFlA
vhtN5a7D1voIWMzZtRA4prkQoFMzwe2vqog3cZebi6CbSyHOYmBmf5E6U8k7EgVK
m0fkA70BUbBsgX88ybzaCXRZH4mzA1vEP2srBd/Dg6qt1itvTJ7QPC8MFF7m0jWU
veRE4ShWiqu7KOxWe/CSSerSURhRGwMMYICTLjHWEjRj3HKdjW56Ta2OgKXyF4QD
dgkMWsh9hW3ffarVGPIAb3+LU+dnsDpdMxs2y9R1UyNICAm5lx72y7V2+1m6/d46
sG9cgM/ws6GJmwxY2YOiG3N8Wcu7FuiPaAQ+qNesb0EX3S9qRTOZIptyhUM9/dn3
fBCme0YK+SfGPBmkVAUU4dnUbg+GoVaUIpy22lL1WNWxyv+a5TORr53huImLe5Do
+jSGaSjNrx8ZAUw6WB6abFOZtWkOBPVWaUO4RP+eQbDrELY4sr09j2PJ3kQcbGe4
OwPGtq9F/HNHyHAZm1rhmET27GrCZKqmJiKGoa59XyvYmgfjDPejQysx0ogTuE4R
Q8tu/5afVSxPE/Kg3mDDU6sC5Sb8Jf1eOxy2yP8KWlqjwn2Y/+MD16VoWKUH6UpU
FePBWznFhrfQxRNyTQNIAoxK2N2iHWq91wPIIuS7XD8H4S4TqrL8SZNIQW8vKqnZ
RkD/TZa7dmqKzvro8uCR6gkiytET5ZeLsJ71dLk1vkbHsdV5nl8L/ZB+W3vUH9VR
o6mI43j0nrH8lmo3i1JZDk/Xx8269UAuYxDkKLZ/rxUsAwSIWOGKNbkRRewgh738
vuZha8CN35c093pIaRfULgt5R8uNYVPO+QZ8NVsESCcmGnk3Ibct62bewK8nHX5w
dBXzVXterTW6S03N/e9ievmUiVYQ7xMgoSDcEb37/yvXOzP7rFCxe0j1lUaW6l7u
ecGyJXJdYzk2RfSj+0S/n8qj9iwg+ldt28ajDkZ91IDscQZ4kT9SMiqBtzb78CDo
Q4WgQus8fep3/hQpd2TuxnMmQPlk9oqpfZjTXu/rVTnekJmvIGCoWgUIMBBF12HV
Y9kSxqb67oXZBYI27ggRqdwnpmsCVTlXnTzSbQQcysWlUidlehfOmQAnYgE5FKLC
w3Ryv7Z5wKSBe3p3JhSES/hcIyZZorHUr7u2j0NRs3mPFdqwVycv7/BamE6EmgJh
0Uet6G9YKeD/KwDExc4UcmN1nuaXZQ+ZqSjm6/d/DicNkKzJNLHMqU3nRP4GZPWU
20Veuycw+9L8TQSdP4dl9F1jdS92weAbkB8O9gX7fmCyXKPF15jbgO1j4iuxgsar
hSul+ZUC6W6aFYJ/dJWKF7UC/ccDhnPLZFzm3TnZphyPIxX0+cXTDIWso4EwngNd
0gD0ModLF1VFJCqcJz6KYXH+rRe64vdlLBECwushSt3AohYAlXDgDJ1a+RUXILBI
Jfsy8i3t3a6k2CmXfyQeCCN9j+TthwlswA6lUv4bGvkdZ2gDslhO3zjs7RRC0A4E
13ans2JrmcCB9wiqrEFhz+da+M6fUDtsprWFzB1vQnZHABVRog/Ugxc6OlmMvvcd
UfEaWwDVn/0VsSJxA8CwI51qsqD9zHKr07Q62AIn2v1mu0JrMkyMLpL2Pjzy+GWQ
oUmX46A5BeUssmOrCOtbooYsUMoJ2wHCAmbtc7SOGLe4pqwcxJpGk2BZ9Q+x8pM2
LZsO+2Ud94gtRfBwzYncT1rGSwP0CQyq87jcwZvX0XGnPFc54XxAUpf5LB9nF718
O6dOsygBJn9oBqPsCP+Fa396yOq5TAch/xFtoE7ggVOgGmOtOcCtyjEpsKEUxovR
CZO14ilGK04kkTkuNtCFPZSNSJxEL7nbmc7qRLPQ+Ui9mswZwXKvQQuSVztr2LVX
DhzJCgtnkVakNeuM30XecvsH8B9Pzd3Y/FbKEi33ZiZjtN0+cvPc4CpUgG18JZQc
tY+xOqKk45IHqMJAsuLB1QwDnrf8hjP2zG11K2Rn6edL+L7OUs/odA2MGzayls+N
DfWZoQGG0dpKNnezY2lNBYtHxH9a9Jz74T24lPaEETEKq/f4JVuknUBXWyX6cAb5
tBbsXGB0hMAvzBmY1AXdGdcURAOyGT3JJCXKdXyc+VHSKqr1QXcE6JC4thDrxAS9
S3y38DAlcqn8nBqtLCBTSdZ7O9wgt2eublq5RAQJ/bZ0unnuaG348MxFqcS0994N
NV/cmRePxGVzsKd88RYmQEYYvrPSLiJ/Lkbr4RxL5HjH/nq8oE6cj8OCP5Etn6E2
RhujEmr9HVRmIJQyjmY6EySlYhflc2cvBFoQ/0r5OXaVOPe0c7v7qhL1oViHkgDb
yvkmNs/Mhoe/5Z1Qg64CtqhcD1ucKdgl/MMAuE/ViNjvkI0gWl2YT/eMqbYx0wYG
d+i+FjnREoRLyyoT4i8XLALTP7+MzsVH7qRMsqUYcwYF15ijThf+eKIrs2+mF65s
vm99o7E+JGVspHVotcjL5tnz9A/AXH7Szb3WwXt1izjDQzs3fG7izRbfxT/Dpejk
5ojo11LGcbzqewGbkpfy+1RyTviKdQNXZvXo8dqRNtMF79WiMOsQ0AaFYhlJGes5
+xZT1SCGl8jUY8HWZjLCmPwUClYOMoen7STjYHooJ1rXIaJHNeqcDgjrzuntwNkA
+e4+pk8Tyo9GjoknnFegUsZTONKHCyJgB6d2Qdl1xzsHKlUT3M9FGUMpU0JphrH5
B3Twtp3CiiysJt2EsrGik8uNHgdlhubwGucTKpl/ZC+0/oX2mIdVhxe5d8MQR5FX
SwhhmJ544FMJyad0PjqOZGp78QM6Vkg+imZjMaL8pL4n5zm+vC9k5VzrAiaoPp58
iXSI701hvNkbYSxFbPsSQa0iwQbe7dGc7biLnlLYQJPiZTOgjHIp/b3dmIvijyYH
pKAU6uddKd5AdD/Pbrq2PWSmg8YMLX43J0NZVha4ugjQCBnNssiOBj9fmZyrCywK
4JK2t2dLNfvulHoRGk7bLTCUiINV3Mi2mHVfciMOoibQdGck6PTsvIT/dYqk3W9X
bAiG6Ul05S2+VjNtQIzVqG3ZER21aYoN1+0uRnFPJxz24/B+nhNbEjYmcgzNR1vd
oNjwoISx8m1ZmM82ypcpr4+ZhBna4yqORdQbMtYt46Se2SefN8DCU4/LuAncGBU7
gHWasfOxrjzjMp2gcLbZseeck4ZlqCnWROmRUx2pOqDPfdb3QiyHZk55j6I5QAj7
s1caoCAmxMcLtGREaM20WSgxWtXKpv5ARNcd53UYMEB+/nTzgNYkbwPLnDQfz0Qm
eevba7WQuYjJTliSY3eeJfU6uuefhnfGyDkMO/W6Ja1SbOYj8C7NV6xjPlQieWWd
vhbuFnlH5UHmFtNjY1d0xJ75Vh7WwcegEgfbtHRdARrKtqfEUhXUWv+JORrzzVt7
UUM3dd3NA+d79bkUBavLHkSO1ioGuNS926DJyZB4cy01YG3oqWAvqRN97AlAa9KP
mJwl/wu5NktshxWvQGclwk9+Ez3qCtjP7BkEOw0vHWBKxy+u68f7F+vV9vGN/ypM
rMmT8phTiS0sNtPXUde7k788NvukVRLiYqfOF463miIx/Yh+6nOfE2LWwZ+NCae2
9nLljOirEdQ/EfJyWaWwdQYzTST1El6Xv9cXPhNMCvF9vENg8EIHw+ZgFYJFGOf3
7IrTfX1B7+iTtu4YfiECdaEwan6boRzcEzSn9zB8g6L9vel25dbyCRolOMf+EJMu
7ILxeXVGYwqB9MDHGI7oNlgBcA2GY+1mTmcKduqxhs799OowUCY8UjYOBlizhaJs
aVEwdGSabRwrgZcWAX9+xx8reegN8WZVJYBloRc8IH8vcvSRdjQTQM375ipuhhxM
vAZmAG8tGrsV9jb/70CtxuuNNMJ7Zan0ps+1LtHzMv4HD1DZsRGK6vD24Y8rjyqr
vU9AFYtetjHMXL4Zz/dM0dH7MUKfZBoOXttRZuO0YAJOnIZxmrZ3NPRByGvZkrLJ
fo8AQSxLbFRGK7foZB+fKvHcmCBRFRydLN/PIit3Y3O4r6zu+oE1m3trp6Ydyb4p
vj9bYoTtejR1Bu61UvtySfaj4DWjnC5Jl7LSfVy0mJwW2gjTwX0LSTu8eJ6LOax8
qfQO2qKv+gaJbz8dNX5J9rVNYY86svf9Px9FXX8zc+NyrNVXeiMl6iv4tVw1wGAX
W7zIccQPtdYNihWNKmYpQQ9CzNytjivaJtR5A4nhvS2+M1lpohmRgTzY0GDk3fGY
jqNFrx0BCOo47mhvL+06nwh9KsAosQ2hfAfW/otR8G4TFUA0NPzHng/pk5yXWVrM
lTFpEVqFmKRDOt2V73whcebOygI/e0nrbMSn7gAlwiDub15ZL0y4VlfxAFsDftuK
OLmvLvCw0CvjEsS+eO1wOCtCEwkk2Q6T1BkwnShlSCIzypHsCzLjeEbGkOYJ/cX2
LrbjXhwx2R2nrWaBX+0ttAaL930L7kXlaFdh8iQxmVO1Ha1DirLnVzw3wsNHY/Dp
QqxWWe3aEWViW6O3kdjwIjBGX4ue0+D81Vd5gM3Acsicqx6DqgDeH1rYGE+2cVJJ
TeDb8aqhMUQZmXywZIzE5Gi+wGcmhcaHIn2kK8207Gb+fzaDGV48dgT/XnWEj/59
NytYhBSw0g/qBlawM1PrRp8PVzX8q+goCcltNog8Y3V1MEmN3/4Z0s10BkTRHnrd
u3cKhv28x4kDqpwzYVPxVqd6RZsHoTaszENkjddzj05SYcDEpQqoTM8n8NFqvQ8b
I1I/W7fNrhAV+Tymozg73K4LAe7yjuYym2NAxs/QP1K8cWwFpEAdeltB2MMefU2a
r21WmHMPW5t6sFjL8moHU1pSO2snwSNWmCyUhym9c1XzL+o4rYwacr4BQ9I70y8w
VlZsuH3vL2KIKWMD08Mnb07eIy/KeeQH4JSQBLdyV3btuLMUpN2T61Hn8dV6gawW
aUPk64WNX/8IAk9Sxs8oxNu3CugBOHLd24P5Ns4aOAxCPHkmoYN2BMNZigz6JpBy
8KVxIaxvd884hKE+T6gXlCBCKE6lBfEcYsecX85SLfOAXRqdh6VIvayBAfMRDl0l
OVwZVo57iGqc/OZbpOCdCFKIUhhQQcMpCXy8nI3w+KohjqbWZmGh1kA/aAeinpi/
45Zb9bGqcqDUTlHFANO/YB1L1ZiAiNaYK9ofE827DlseJJdFVVppCcZF02Y5F0+L
Jau3p0h3njIutG9k3qP/fS4OgTCzvqpUjKZEC0W6bLszZxboFq1l9qOfHI7Zd2QA
+DUViGPB2uoDXS/f15CNg2FUd8CSf6lNpBEZBBYnzZqzhGJizyBsQROFGOTfjRdu
1mm8hoDadsVDC9m6t6u/GALApSRA3d76ZfwNrChf1PDiyAax7r8s+Zqh9HyboJ1S
U/MMnG7+8IugYn9c/QkFrEYArGHVOq8PdpGo3J7+5OlKVVmxT/81UW6YlAvA4jE4
lfoJhgXxTHee4RKlex0Kg4JqM7BmWWVrVliydNOw4dfOyD7s99RtjJ1fobPYWbdk
e2dS0bitY0Yq/N8MGhGVTMKFuEPvy+XekhXRo7mtaftWElD/4GD+/mbByBJ5ueX3
Di1EWM4OFnuyX102brUu/38TTkcY0JEDxnsL4Djs8atQLNclOqYYqfkhvsr6LAhe
n/BC6EsW/LTMymhl25voVRx/4qUjj1D0c3RiRsgL1ylVeX/WXhS/3yURz9odxUeE
1msJsQqFZsSdNbh3gXQI0aCwx54l6t9WIbNo7Zhne8sBNwz/Mgg7wZa/+y39jrRf
CBsF4wybu1s1o+hfFGuyaVzMP7AdXbcfrw70EJ0VlmilP1CqeRC1gVnsuZFNxUWu
hncwb+esQjI/dZOp0DIbiRQ/t9bliFik/OfqxfdHKYSjrvYDbiw54uPz9cnfkWhM
LMU2qcIfg6DmJRxWNB0niVL88rf0u1rVIrKwp6HqHCY3livVGONrU3Gh21QNojRV
tF1oLJKm6Y3+jJoRAvn2PZ9JleAKVesr+mxSGDb2uWNbRf84MiRuDyikXWSsRmLB
lOLpFiWO7PzIe6+7pq/D5rpRtfadS9cDmB229EuzbYbOk2Fs1sOXkYhiUVG1aIQG
jbrAsrvgu0kLY4qPx+DQKgCNFpwV4B4YFq04o7pSDzTz8Li5J2Igjafbfh7Udsxq
Q1te6sSn9khA2wT30ogvjyIYtRwnxiIAHuk+n4HmU8FhzVIS6IF0XtA6r5QbM7rT
CSWE8GpKzvH97DTFcHIh8eoc6KoHjS9lWgNxvUtupXtTRGWEqim/m/PGDtuJTHTb
jZQzSO5D8YbK1LlVExA0WEdU4mLZ1M8ibjuNVS71zqHWh4BEFq/8rNirRgcnOUz6
CPg6p5FpcFXE8zLq+Hs2BtywKHTNIBaY416w0/J6XH7wbq6OUX/30j8zg4E04byM
fBtPjNz3qi+Em3UNvwaaYrsgCAUl10fLLPdKyyW/NcjdCTysi1E5UPSQU9qDtDEc
LxPsmgZZOtXYpDp3R4s9Nr188I9HEQ/xf6JL0D9qqFT/MuCI6tUJNB/93NW4nQdR
1FHCyPDMkLlVUZGuwba93ISJy7xmHCPtykGPlH0knu0dSrvTYr5ggB+blUa8v3X4
E+Tol1u1Rv6khtFlZ3Jio42qIj5xfDfodx8qDSff7xsiLUko5HdGCXh+QxxuZjzX
Tq0euzgOmSI22E8xMBoJY+2M6OD0O1EFGTO0ZrdYlD140x3SoLG/qE8IaMvohOqo
b1iNK3P9pQgLHHT+c0bBpNgSKWwq5PlzuYlh1BIhr88neDHMW/eNrg2Tvw6O/VXo
Qvr8/pyCSihjObzSWj0L/3Hb8C6NlNcuxb7fDHy480g2/8/7grcK8e6HqLIbyZNN
e4smjWMQh2XPDj3kQaqlS/raofEn+rpJsMwS4whV0K8NYquTS+LraXtkfKBJqopm
TsKHg1mHZhfl2Wu1Bv8obpZsqzdlBNlWsMkA5QjQ+5Q/Et5WYgiFnCtGCJaVsyAq
aCHqQW0lY1yxYeiCrl7eOCUyg8wLoLiPJOBvqqgbYXPn/qLH3H8bHwBDvlbaJQJh
eBN0gOLWJLU5g8imzecuY7IyAKb9do2uJsTyuJKX1B54KJDSA24XdWiIwc+y9mLt
RoNdXTo1N7JtSeiMJo4dc3GbIK/xV5Nev9wTHiv4pQ6Qxbt2se25JAqW2myGVe0q
/QE6PX0icWoTp8Ev/MNDhZEvPkCWpRn7n9I7oBGVAFl4679kD+PDIkISUn5YKj/F
AitgfXyZGi/rpl2vjZ61uuy7SizrJS3FNHDJEBaHENC23rb/1QpgaWKFnPwdhPJ2
nGdaVyg0VVZGEQBe33/c1NVx2YaERg+GK2UspZQnUPqnoONd+/GhwbhEahE7qtja
g97TjRCt272CnxY/8NJDQ5pALuIubFHjsXoNTEmpTSaw5lShqo3kUDk7wj+1KAT6
v2MqyEuoIhmEybzSTWz23mdXoO1MofhxNZgVLT8G6Y/YjrpNBZ0055a0eRpZMQLN
0+K1JheceOR0x4otFZXwVyOR8Lo+m2noRF85dwGVfxeMblBZ7M/EEio4J/PnAaD0
QA9bGFHefQIUgY/fOPzylL+os9fSa2dj96YB27XdULaqnokHxDjW1Np4JNFPBMJt
BmCp2xYNPhwhu1s8NeMLcoxyG8BTVWcV8ilhe6RvIDS9igQ5t9vR0D0aN2p5+snI
o9IVFHkK/GAJlkTUolXh9GyREjORjr2jSBtRGI2e5mPUmzBFAUlIR+4+/mVh1eEk
lwbZr+BamJDngoMgOZtXtS0fR1sr4hjnoP/uQuw3hD5JytPYvEyi7mMWiuZgBO5V
lmYx9w9ERfQ2YqhgfX4OD9iwUwQAAJjyncj+80Yf3WcMKm4kd6gVsPN87m4IIdUb
ptWjHnajTsnzyyUWswfvhbEyLj+7h9cioRxcMqcplYP+mR4GkDj4wcTkr3AHVt7w
VjNzcXKxdzVifoBNm5SYIfv2AUN9cfCMYfvgEvXlebNvtG5qfQ+H/+5wqK5oXNdl
bq+fNuvipepG71hE2RESb6F+9s/twGLBDIVYGvNSCeyCS6iAZTkAC/4+pDJShSYd
OnvCYyLf7jWwdjPuGd3PUGaCUP0Ko1jW2+Hc/+h+DkLjmJxu6nnC5S9eAvvGAbay
JwkVxeESt+0XbL9eP9p0+gUrzqOaRbSjeEtXv3BjKoSgZkCzuqstuiszIt0xy43K
qxC59J9Z6oS8Ij8IdmRzGY21G+HuV5n83KFHnYjwO4FaPYoW0Rcqxf1NIAGjkXXo
owaaxNlo2mgeFrCmzvGklWYz1uRakK1ztQrnVEtpsu9QB91JWGu9Ytgwq2hIfHaz
CgOd1oOFr93P44a+9XEEG5qsdEzZustuohy9wQxN4IoCRwov2CqR9byW/EEuoC7u
VVi5bqAO23RfbVeOVQe5FHsZeWxyMrJGvW6Thz32gMaZsHl2Cny/QtlfbwTaEfT8
724IOWJTAPUmVnoFdXkhJU56BWb7mLDO4RbFeZRoIwmIfzEMaiEwDE/boiLX1teG
DMJCUlGXEk15D94htuZJSGh1soaWveONsfUfqhdgFmT7zmMeuK8ETCBDlf0Nejcz
Wjl4AJ4g9cfXdcmZ2UXcGfBuJbY2fJ/6OUCYHec5hBpLKoiq52r7XP/e1Z7pMMdv
jEbQ5gjR1nVG/17opWVRSM5U47WkvMGvIcj3Dar1T5KHc4UImb4C+Zxc1ytwzfpa
QsU6/0Suh1KUNViLW0a/l+XAOPcCMzj1XjEnn7Oe7bVSp1Cvqqm0yCTXlpAUHj89
e5sLVwhuRiGKlxKrP+gDHPc47woQyTk5yx8pYxJAVU7+Pqj2jSFFtRPJns6k4cNR
zgRu6pqakcPiCYQIuX4htCw+61TCTRWayxDenvVTjVVEgijSUCYqDrHUTBm+iAvw
WXD57An1OusUZxWBp0Qi+VCp8FP85u2F2AC0edgQ0RH8FCkDo6FGDL4h+jI8YAYp
Pl0Mz/q4aNvC7Gc/cAZk1wluC9JgiQ9PyAJ2++z356qPHdSulw2BEEqBSa0hvS4O
9yvmutW7n5hcx8Cxnn/1C4cohgq533fmGKTwPvtIaV4brtYLyARgBzCAmejoBiKe
3SigqL5eMsB89PkQglwYttiBGWkz3xj/+VOH3/xLpYYPREwevKMNAc2qgBA/K36J
Q/ZEe5qQ4Mv5H4G2vnT5/hMifJQ+7vYdlwnAYklQ507nEOfblPJUspK9fnoXQuvC
NP2C/fd2jZuPRWZMqXn3MSHZPbieJKV88Jfj69cuR5j5iyrqo80S20hqv0xGmAt7
EYpLahi/34YJ0kTUz1GsoyONbyW0K6NdEcVZY6lYtUSDhRT2l5G4rthKuDehRLBj
oe5WeO2D+FyVe/on4VDFeJOO+wqbXX6zgX1+UX6MdD6lcSaHXOeR1jJT3EgOizAp
gsoJVzosAm6ihNa8lRnKufYEBfLvtPhkLAwVhfvJqgFj/eX0gcTMzhdw+tCRY8BC
mkG5bFAzr/4q7M/zU+Y1JMOfJsV0xYOxEzs7dqJKLg8elH2qwI4O9HupylP1zbPR
/TBeIse51rXprVnjhSrx93Uwjs2lhKMG4rv8RDHamFH2M6fm3IcJovG6rHiWaC9Q
lFXFqj6L0+lkTJpWeiWEBNts7JeAmS8AwIjXYkRjw1iY9d1snN5H9vjgZQPnjxfD
Jq7wxjTewvOfPFf3bk/J/jdJD6xOJ1EIiJxkJHxB8PXAFxLl3sPLItsxi3k51+u0
6BPAfwXVPS+6pWP/n8ZdDgNgbQZOFNhrz2kEb5yN4oU3h3TD8N1sQlRF03SOJsHO
j0ewE6wBo3Xf+eAtxctVIMVJAdPYs2+JweKrWJZ/kFIwZq2Rfp/6BN4cgErQvv5q
w3F+K2jEVeejiLw1WeGvEwzjDuIVl+c5TN7Fc5ZggFKRDI0FhOSeSQnZ21bV/txe
TEgmuEAzqGy+im9X4/PYQNW+7ByjP9N3rFVLOxy4wWWU+xKl+R5v65rs6cL1KnPh
mVu3+36s/CRhovWCoP5lQHud/lxKAfhtLLHPCBEw6s6ki2yyexsX1KO/sI0H1KRO
FimQA+EPpMmsP6OlOQ5YAQaT78wdNy8kthbqIwoAY80FPh5jKIcOxMJABspEzdNC
dG2o9U8TvSIH6b3febT6dBFWU0DPvWnnfSqi+HnDoddfoNjeZZqLp2DKmTMBR7xt
UmND7X+zGnDa3L1U1FTpT4nFZlOrMUELx7suz7VdNK5YKZpaqHNQBw1u98vTHlEp
rXHHQV7qsizg+SVcM34FPAr7OeF6SVFoXcdsiqfIO3iaSwewfbAMdTCR27itAo70
6zMCkCqsNejGsP4kzZAmJq5poxzX/DUCDW9lIJyly2DIKJ0gX6mlf2w2aZNeBxqV
+Cqv/ES0DDvXS9VNnmpBbqxtlZC0JhoaR6Ocnr5RijTqBOkgknlBOeCccypZqosv
AafP9kA/y/dPzKTw2l6HP0/rk0fV7yY3SXHsUl9bezMn6u4u+rO/jXVc8ly1hbCi
w1pzbIHHyM3Sym641Z9UJ7Jhl2SqLkFUZGuu78XlXzHP448yVCDXN+DeARtmCyxQ
5tgKL804f5lqI7cDozrND5Fez3XQPh7CoAhJAFhHOjij5r0fYhQ3Jd4CzBY/gaia
6pzIkt9KmxcklHfiiDv2GDxmufnOk208feXw2nejtDbp6gGwVeQ8zMIpMzZypMIR
k2Mu0N0ItkN1Gi67kCHQMrKf3Z+ct7zNUa0vMrY5ETRJv6bTZRAv/4NQJdIZbAcx
pWvDzVV+0Lwrp6k6/hna3/auxChH/Td5XRks0x7+4hfho2AUYLpkHmYcRJA4gc3d
Mmd6w+qzT+hm1sXvwhtveiwS6c08nAuRVpujTMjHr6WExn4MUUryRJ158ibdSzTc
cF1j++dxwF4qc4FlmwvQlLd4FAXOhctGSS4mGe75BbekCiXNhgaLjUp/v0tquy3z
zdwFNSWdeA8ctnFxtufDqKMwvzMCiQL28IYQ56GG1KAzlqt8JQRsz2S/JKwYAFBI
3l7JoREOlXP3aiJtpC0UcnAVIdPUJmX5lc2SAN43xtJ7sVbApQq3aiD2ME4cpm9z
+vIr36r6UN2mrIPcs+ubyctB+HFZu9NzeQN6KLIIlW+gboFP1t0J/CrF7gKu126Q
8LNxoC/0znSdhUSqzicIVaGzT2DI0VCaGJrXEwI1Sr30cuIjYqlsfRYQbe0aAixB
akizdA4TxkLKY7mbZfpPy5gABJ5PIBhT6sAE56TNA+sVem20NPWQTlVyKhSQPzh/
H7QiacRR/u//6khmu/rPDYa91uwz0wGRL+P7ww75BOvkA9l6CpEn8aphGfFVvYbd
EbYAAuSPeHYegaioMlKG/p3RrCfj+J4H/b0AKBHAjXrObXaGZ/5Ljd+yZQfm4sOk
jxbnSzXFQa1tWpDSk0cCWv0VK0ft/1+I5UpIA4Dler8LZkTENCwp6ZLC+XeHBUXh
69GmGxh6lpvw3f6BUKAJjrx2Z7INkptJhSvVKxavigTOl2USstNIga3iny/rkfIP
JvQd1WZuplhkFLJA+WhgWwWp39znBIC8wbF4Xt/4EX0uDUa1qOci3sk/Kk0n7kCj
42CI+Rsl1X5p2Iz0Mjxvpn1qSUCDVkPONV1Ts+saCU2fKUtGJTYjDrb7jYkKiGVo
MFEHUIz8m0K3ilB/zaH5EtZ+1TFM2u8jHgL0k/1HucM9JZvdN7dTUcNAt6aKePRd
E1/b4DGIwyldy5sopk3B1HuZ63M4Sm3Q20Qm5tUQoVpk30rGtb8jQWIQD7o0088U
4drV1XZ+mzAVNE/ib14CRotCnFxupMmPQ21+wTNrvovTLzHftCV2yaw7Ecn/xref
gKNsAV2hvS5IYLEjFeg2mzp5/uJgBrhb5GzfpN/re7PTekjk4jduYIX3F+H+3kbP
WgfW+siZdAeX3QsmHufIKTSQqnid/Dw6gu7owK9TP1PL0h/+Ktmpj4P6Nqm9iFXA
xFJiac8v/04I9l1RDHJclF2mrgiqhMw3Ull0EBj48zTimFEBKf6flqufzInsoMxd
1e2K/VfTIVJJBvG7Ws4dp9PVpOTi4P66pyqjlbbHhwwrcO1uB9wT5AcaH6A5WCul
B+UJBScSakk9gcSz3IAzRN252L+rZCUFisSeLlK1UhU7TBgqhWXiiH8YpINEnieJ
pkWsEDQmWQpww49mQRchh3Xhimbd+hqCTA8d1qGewSH3sncedjOJvBXPMywVdmfR
oUqQXXA3LAuJ8FBXeq6BHYMA89B48pWyMaqZmvPEYrrXmxO7gkvvzfq2528Y9emB
vQyKPc0sMRyaPa6HblC+kUAt1ZSS+ZG7YO+k7dPI7Pb9M9TYmcn7pDAOSnbTlReA
qRHL2xhGIkRVoRTVEWO3qJwotfKM2ZkxSBvpqteGzJzTuwygpWrIRdT1ow1+velT
fQhzkEQZcWwNQ2mM5CR7ZcqOqqX/tVZ8i/WNKIKTX5VSjKakDRNdAstZtjqAduAT
tCWTarjkQNECNztm6nkDtQzlVJ3yv4WJrvXRLrqJPRT3kbygsSsTCjh1+hLK2/xL
f+0rz0k8XCSBXxJKQOeFrRIRChM+gICsOnYXgdUkr5DEnwCy4i/m7uREynRlkMzw
Tb4guao/z4115fnnE8DD/YPMwW2ugrdnK/k7IM5UbQMZcSFAUUVvKCWkRcYA+Hry
h762Tq9REFDgOf0NbQGvkIS2ouCVv01Q/M0YOy2naka6s6GWTauQPyee5kSEweZ+
PlHmtOie1Thl5rLeGBg8z8JAyYNbEYRS7sVlRGhejFrjAiWZhW97MelzOY03TfOb
Z7CyKfb8OWrQj9PoZlFQa2txw8qTzMdKDFvqPaJZdkxrzU1hUNWHD65KDOjzsIIT
lbUCcgcjEMjSyywP0qzMUJ0Kdix27Ljvs0IlVusCnlhZnUOZ7QqSbSs9feElwZeh
zM9zWEqnjw+1K2jU2ScdwfxboNojGZ+ZuPL8nzxEoTw4bnI/obnqKAEuURQ53xnz
X/iNmLeEXVIuM9aYJ3eIfndwE4itIz9OYOxMgcKNWjLFrnXu6jzs0lPj8U17ypp7
xw//1r6zGKQ3eFnlbfFS5278wSn6Fhts9p9lINaPSgWhzyEpesqXGZaMw05D0sxU
XmCZVP0m0KjrBTqbNL+7mLb+59qD7QItWLXSJVHiHM3q07AFo6r8RdJ1qQROnt0Y
oWxkvxGFUn5SZy7hyXZujwsI86UF8pCL25K9kKdWRblWm3H23NIIoPEJQdM8BDG/
YVAQg4Uw6ncwi2krpxKO+MVJb82AE5YJGRzWsdPdOE08aMHn8QGgUs2ij+PB4TYP
GDbfGManeV4FQ+p9b4kKgfrWkHSIZIrNPQV8x6GizzEDI4gj7Pg7+22t6D1yn4Gq
PXi57xF5ln4UjpqbpbijejrtitrwunHOiSFurKUFq1owdWvzJpkE24bTK5hL1cmY
/6KRyiaFi8Dznwiit3TAY5WCu7dLaRRAbMH0wNI0KQw4H9leOlgFTMjog7Z4Ki27
XcxlG1N+slYUhvOVqK3tEmfO7lkmvFtjX7ECcSITTO2Tpx8OwxJvNDAuQ57E7RK1
xWtp6MkRyCvGLM/KyLiMcvqDSL8nhSagkN0BIAiDW6kCsKSA3Y7sUOd9fP4Ct2mI
6D02JSV8H0bZY2taJyZvi3BwRFRih8zUNKxhCGUNdfVLPJlmpee8+03JTHnMXZVr
muTho0gYeLCJ38W29SIldZGctp1aMwo0tfOhWKY8yM4an4kDU7r9Sbporbz5Kdot
AZVd+vB9RWsQEVJ91FrOvhjrjGiDCpqo2rhgkt34r8vmFMOKyFkvA0mYsZwI6Sh8
BFx8cpiSLFJg29g9yzYE/Svyp5xfJ5rmPOb/NHjKtz2jd6GAPyB5K0nrbypC145q
bX3s96A36npQ8AqkijKLWC8D8A4hXZ8Vi4b07m8Lpubh/wnYizi5+v1RQwo2UtdD
NepSja7awTIz7iKI8fpFGTVj1MiF9QfPEqvGJmNbDjDQVAy58WuyRbGLxiYusf2j
CSam4hBwaf9iak08oIg4YMXS3FmjWgoVG2sDxzbVB9kdc95FMmFa7nNuM3FojIAs
DFrK0m9/PCY4QF9z0RRJHsqwJhe3gj/UHiwancac37p3eism+9R1eR02S24Rambp
Ht1/cjsqprKgTN50yUnN0cAAhD0VVOYo68/k66Ho1Df1lCG/ANYv5nSqinAR11kD
Epkvjyd6w6SmBVsXDan7AlQ5cPsB2CTCM41WnMj28WHNn4mo4Wsj5HQvoujd9e7Q
7U9NZbtH/5MNHKcJwaoIcW8k7LnOcB87RzWoWgTqyEgJTV1Xf/mJ0oyjKqcVvOiv
rscgKeqLIOEY/VXNW3qcxyo0gP8ay6V5e6Y/H5ZLIGdpWZfR0jNzvh6nDU390YVR
9p1rAjbNQ4eOU9Tc0I2RVaVxtuZO5LeWXgKSOjJuHSfrKRXhOC29HlQO9g1WeJSo
5xBK2pyRKPQm9P3UracVx3u1cgRjhtwlG8yAcdQhfvjpQVCi/tdKULkmKzizSXVy
TB7qi0I2eUVA7aWnhC88q6A6e1N2/rGQ2k5tp7koEPzwj4N7NkjvYCECnEHoIngp
hgLcB8ykPQA8N6psfug9pjvDulYQriM4HHJHr9iV9RYlPwN7d4kEqwb6ml/noy+j
1I9NCIHJ8/wgWU7rqvF32lRPDcGMEPAY8w75xphDj3/D3cJZxuthMIw86yk708vJ
jOJLZct3aA8tCfDT5CTMCLQGxCHds7SZJGZZyNCuB/ylBZ3+BrQ2UwZRwNy7poqd
8+BfM1XjkzQNrtE+L3sMwaqkw7rNBk2AG6POPQKu8UPcPUhG4dKMdaif6d9yv0Qn
F4Bg6mGvCeTvX8Weiw1s2OIcycO91DT+FLEywijG57QWLzbZd2bXn2/leqGmWdjc
HcSOl8Z303Kua7z3Z0AYa8yDbF4GSx7YUcQyRO2FhoOGRIhn8eYiZ+TCr9gTfPlR
z5UxMa1hZWxkoaIcuJME/Uj54J6T0HGKZfsve74DYqvQ7LjSZHi3zb5hQ2VoOj5N
VcYwSK2gPsEp4ZpZVX5D9/SLENhKCr+QQCRtJ8anN020KUqxLBJAcJ0NsFckpl0h
eD+Ur9cA7lIWu1SnuNIW8lKtR4S0D0gNIB95J0+CTNG8jcS8mwNQWS32LKlBMgiW
oioT0WD+2CZl4+Kf3MgqOnQ90eHFM4fdWsxydPXNvEwOX5JAXcH64gWPJyMIPQa2
UcUM3smqS0eJWzj3rNiuYcQBO/sRXAww0F4X+M64YtY2Mj8Lirmy0X0jV38ZqFfO
tKMe8BOkJj6jz0/JQHMqafiOioiMAzZIGU+vTTtQKLCZwsWVL4OitD1ze4kUnz6O
0X2f+Ha8P4Q4wDaOQJV6fhWJdzVvrm1eBjflqlHiK8dtt1Abno110qTBvnPB3PS2
VZLxOFYG/G2CUdZIY+eCj2LOz/t/pHduHUaEFeYFD6dw4hbQFa9wybd5DdCaZ4JS
YS+uuTEg9h5GP667cRVmEAqRnkJasOQE11sfIio9LsSW79XpNPg+xirnhJcCaoHr
k1NZ50SA7VHFcZ4Xd0IwNDO0MR44e6CxOIcxiP5mdgwwKdWTK3etz753YpYIM886
l/xovb3taTaZqf46dLPy9jhMmNQc2wHaHPg8Lb2ljJjYn7XSosjLHC4aIyheSLD5
lA8/A5RDv6fgFi+ZB0HHvqeNz+BYFH7r3KkxZN+MfgSxX+9XFH5mT13jDWVTYghR
uPv+IWIAvq8wmAsiKtIoHXVttKSwZO5MxjRdX4pAqnS5lbEJBIXX1OmyarQs4rwF
zhFNpR30rr0IBDdfx1gQEP9CcF7xF/u34gd+5SC8sTRranTgpdW6sbgAUYqDUFHp
+QAznBKC6owFaAv68hpCcYciIzZxpcL/8qZKUd5zpkVZol74pKiEJSyngBsQ3WIe
uCWAp0PJLbbeh28NWwgmwUn10b0ExuYf6nFlyihVDXrKpL5eKhQxFkqP3dBntgA8
4qqKKZ0hKEUdHZapW65+O+VYPne9vK3EnlBSTXZRtoOL1P3CJ9/nZq2TqavnbB/G
xcNmq/c1A8z1ohsH+WV860EFIyPIedyRJj9oHWEzhvoDQMnG0/voREmsEtRB6YeH
/r1sZqygcyAgyIKcT48IVqeE0F4Sg1TrzhLp7sj7L8ml/s0LVRDw5gWp9T+8yePh
/ZvHphYRNftjP+vjVkb4h9qEOOz0WqVLL2Zw/BAIdWT3RQqAmfp5RHrjcooj35/h
dsuLKEu92SaSsnGG2uyRl9y1bDf2vd3LNbSZNsCLOxCqLO7k+PQCm1yDv6msJHhx
xdxAw8tavjVEJcf0RDrRynmlrs17e0oH36NkEi8IoJ+ge3gNfC7X0FQGfcCQWMNX
+aUmJ5/ZylB+jnxIOeBTsOEahcWSRh+mMsC7wuHwggPoBwtOWKp3kJPJLBps9jq9
L0vEw0eHGHAd833TurxMBOss/AtXgPAPTZ4jR31b3FCuiFvNmz0ViYv2rKU+yN+n
qL4IZza4BiTZa7PjwTArzXcZ9tibgdWwcFmcBHpaiLiUtH5jMtmMxyhjc2+n63NR
MyAEj98R3q9wWuvSjCV84/Z+OBKrahx3TZgqnBVAo1SZcjbdXTx3DU4EzroE03eo
ZBt/oY2yO7T5mNe1YDyT1YvuxjV4wGXquVZ/tQu2M5umg6qHkjfHbLcJ/mF9Cu9Y
UnUYHDeHzbuxdNKSXyI3zjbBQyzHrGeVe3ica5bABUcXJpilmdjNe6kYQ2vZwaWZ
kCMQqnN3Wg3Nhur9R8BvOYpnovV5DFqbVqYuvrieDoPTWVINvkAj5qFC7iQ7LZhm
hqqi6YaJgihm50TLpT5sEpza+zUvyi66x3EDLeElwZF9nWiynvNua4PBn/o5bEt8
11QVv9zSAc9ud61R/x0kS5SmuP6gLgt/TYyV5bTpPxzuvsVTy25FOtMAbogxfrer
5/2tJEV7upxIKuJXCh95hwwypGNM+iZ4RGdnzNOBEdz1/6thvGM4pkfo/+qh6xrJ
GRh4mqPlMiJe8HxDvPU5HoXjSBJBAcUYI9yIjk0c6kbcF0KzuvugImHbxVh9kP0P
r7RQRGWG3mQNbIOxAmZ1AoTuEogIMxNzyIXkMbPBtY9nVmTGJSEOHUMow8e1+x65
4ssUBGrJ+M+cft8jjGZw9c6z6gBWNX1cZV3FySFv8336xnRsoRZICleASQRk3Cy+
hI8RWhEfcMqmToc5676kH5rO3iN7wyVLDZYzw4POtBDxbhAnAWNPfC7qeV61r3Uk
JMo00SxdRDYDYw8T/DUpG5GY20ldlISKvOzCikgvEOn6qLR3adJTluOLjt2+Ke4m
HHliAGFet0H+LGDGK8Ns5F1dqeCkzzoi8DtY81ZCbCPJt7nRVp7FvnGcoyPHVSQg
auTeDwY4n8nrLwMyq+Tu7QFSWEig/yUUQKSnbdzCrf1x+a5KtIjG+r8/XNEKKpM6
uueKespTkIoXKCvh9CvPZxudmD5NXTXcoB+EMHWjSGNPrv+18YvQx4tfZnHr2dqf
CQ5le/kWg4O89qGwl7pvQhg+qQOWZ+HrE4unr6h5ukwnX5aO2xQeGsXzSgbTtc+V
SpAgov22geRkWUGGvOa/awd8U4hBcBmIHYEUI5/aCMSFpnWG7tyEfOAyWacwNnf5
xjOmFs9BvZX6T/hwfAqHBu8x7BmzvLnP1QSHeq70ozdyl0OQ6copRtRVIwG9zBLn
w57V0tD6H1LU/m3QE0UaA3TVXEACKvnHlt07prMRGVX9ENdP9AyamtQah1uSMH15
+9G/DAmxCyC0j3vNGzYQdkGQZ+0ryKbH4v/RrFqyqdrh6K1tggfS3PE2V31+65hS
duDIoyfyRXQKltmq4K0VRPyeYTSRvuSmL994jWDE5B5530TjqsNoToeplzmPBccw
UuatTQeg5YvaywkeV8YS0XYOyqQZYKpDJ9pJzCfcK9wXofhItoghEuObLmcYevMN
3+3qcGaARmQZ4PwhUfX9HxmeKsxlj2XC8adPugoOavfZyjXcpALt6qVlpMu1Ush2
M/2/SKhRXiKhGwkBGAq967KhbLYD+wQE8VrTZBuT4StV34NAaROwNmO11lkXI9cH
FEQ0c5ZkpXZ6rHzlePqb1xq77HkD6C52YV4JRQXx7HjapAKsPjNS+qpqllE18Gby
wUeSJI/BV06o6bl21klNmOxBjMp3qhzg2GnRv7hMNgarKhcj/UQSA7HKtxfdZLSJ
gN8vK00Z3bjwj7DVU8U0qixpsTpExhS1m1v2lHHXtJlYAQ8kvX9FzW2Ld8sGfyiD
9K8AfcgC9RYlrpAisVgZRidNVgGA0BLf17doPXlZL/4nZgJYwAHyfAME3gU8hHoZ
fgzWdE8ArtyVNt43j1ygFGJiXea0ni6Lp1+/DeJh6FSSyJpTu3cS61lPWjJm9M9w
EGOQ4v4PvWbCvtPZnxYbiS3o4alrBaEhOvKhc2MRLUlVn6WA+mDD9bFcWzVtgijQ
4ArfpaR/r6VPfTvrAIqUYP5nT1078V8UOakrwgsnWhRSgkJk1bNQWTd+tZkuvipc
J0WvVIqFYznda3eS+SKaN6oyfCFg6usmfwKaJUHrB0gpjTcb9AI066V+j7VgCDid
iAoowG2Cdxp703lrXVj5AmGEKyngZG8C6QIKnIznC2zABhdcwpkMRtFJ7x3qdDYa
CgwC6qSe4HWJLFaIKzebUhzLHzgRrNGlq22XmXVFxozGxJUitmhxBDRQAlbjJXoy
jNVVVH/GFD4NAHlWcgWjS1NeQGAgIkDD5v6vqAwZz3TxeA1ty8uzVw2YoMfYWzVZ
txn9Lh/nAR+3CVAY1l6N5W/1gAgAbg+sbL7MubJxbWJaxW7eQCLO3a+5gCDLXT0H
pNFTE1nW+VD+EpRRaDbLn3HmXG0T1DxAzEDFyw2FGwN9qlaMP3mj6Tqd448FR+c1
okSmaLGQst3R4EEPK9hjABOo8IXeNxKHUSJWycW5J7FV/ZvKZmoQF6eJg+bkpjtQ
EAM4tu7XGTOjPVpDtoprcATG69uylfCR83Xk25BtI0XCRrnozpcXOXft0zOvyy67
8rtC7cqzdHxgdUwkGIu57VSHvCvID1WyUUC/jyNLWHGhE2WTqVfBMNRTipNK/j4X
8pAwBJMDnEuTwj3q7lwhHRha3uY7/s7hoZKdzZVh9TbUoN2YzbzgIGI0/GdDYwgW
PYG1+v19JA2TpbwUDkvSTqMURG3F8iWzC3TDKgb3UXP9nfbfuJshADhBSrzUrSGx
m0vgDE0ccKMdq/vVCk+dMJzdM6lOZ2fLzwqzMLmQ3pjWQcppuQA+vm6VZS0eT8T5
E9okbN58Zm49VQl0EI+PLP2tegTFnoUWOUvDym44Z0PuGMgYs6LkdYWqJz/uqqcu
8hXSzevTu+fmFy+gyQOYh047R1HiCLipYWwD+SnxKteJR1zYtu6UMrvK/Gqyrjuj
DBc3GRKClhp1K6duCDyeYE/du5QoUYGPzRfK5Bz9tOzwJcQvJD9eNok8uEOkuL5k
daMT0X7i8d/pso0DMuiVBpTjHN+6GKrvhSJsJpT1NLL7SDCOBhpQxCR/80EtP0BB
NzVB4HogeumS36X9QFg0U8ABKp9mqnwCTXLPkNWCmrA1amlUVHgD20zlZ2qq4tYB
RX16rMvdaY5tLGcHN5CR92byEcM2TBr7TK+gO10wr461Vt1/nQulzjkmHOQar29p
EiyMYB+v5SizwSbhIUIgAPLlbvPmPrRkXefkJZHIq6jRfdAgfhuk25fE2Wyokiq0
ql1It+l99lzOqBYsGAhzUlnHX0SHtf8MSmmE6Tmq9+ACLA3SOvCbuKcj8UNvcFdu
YIthLEl8ld1rptW+n2NHYIPRp0YzCXCXgs/fsBwtsnusRAf1yNiugvcCrdgvcgM/
XgYSyLA9lILjJlYP3v2S37GrdzaAC+97oSxUSPbFb0SCHrxqOLEuWmLZ75Srf+o6
LCQK01ak9hDf9nUM9cN6MherN/u4RjmMXffvH/bmGLiB/SUEfNNpNM/TfJheua9I
9Cs1OLnLyvz7gLrJzxx2SWOKWaYCDrQJQUtus03WEAQAubSau3es5Z0LOJmuvler
8UM1QpF/FdH20jvLfyCPSB16vzLruw1SxojUNb31JZMwyiEA1HyWCne+FOI5+tbf
Hw1I5dCxKfmGRZJWzohOWtniT/ZGGN/oiUrX2XHUC/qFHnqRd4V3smyc/Qs6uzA2
nIiXWRq1m0yA040PtyYUfWcOovwzue6YZ6f21NXFhE88fWAM/eO9plKOXq2204Wl
+m3jf0k48/2THRWSB+usR4msy3+/xvp+41y/f7QDG3D7jGGVwCi0EyD5HbLEFIle
0euFqxPJfcrJPdpEOEegG88MUN+Rq0BZjec/FDOAfK1PWSC3Z+FqJyjfVXDD0AQw
CtynZFqG7UOVkhnLh1ddQMyEPtzSy6rRQGEBkJ519V5TVYtNimccFEfD3OMHL7gf
5WFHdOaO05rb2L39DJ1wH575vkHx2AHBmaKUp0vt1u54qxNyAL8dCsGvWfPSYwDu
puhkVFhpNlFLP9iHxSJNDUxp49x8WC5+RbSCeu9NLT+kL1aolVRUQAI6+5VGhZgO
gvNqmviXebrwFjO8QqlDdV+t/CvkE5x5vgmoFMM088XcoLxwVQUJxD1O5MnQEDjV
+T3Ack5ByZd0QKZoMybYMMsuABPIIm/c35Ej72zEW5L40uEGJFCDG1IElCEF7avz
ivD6TkYKbj1pvNw6b/jVIrtdZfJZ7opniIgQLTGE87kafruQ71uaS+8r+xEucwht
WETPIpVlJ5xR10aN4kxX2CgyV+ozoWeujSHjluo7WPRtqyS+BmvXv7S+sYvDiaG2
C5FJz/vah9u0J+kDChEL3Vkz3Ikzi1Ybh+O6sNQNSapUrgU+2oy4lECCrccnhu+Y
jVxJzAKpvoVZRRbZuimE+V2MHdpXyOlAsF74k2QcYGAtVEsV+nuW8Ft+32J4VkqS
4eAxgWZUa2dqRS0fQUPeZQ64hbVOroH7b/3Baqpm7taqrvlzR0Wyilnc1JXdxjNY
3QVEiLkgKtZLUXodMB7OdfPxSwSGcec3FkojB5ZAhrXkOc6oT4bEqFMZ327OWJOZ
nhha2QtydFW2qCvbOCrNqnZ09s8dxk/jdA+tjMVP2bqWedtsnTaHaffYYQcwFwE+
m7kdm216PGT4jLVFFJmj7BKy71K04NrXuM5qa9ly06iP0ET05PtxeI7aQPVRorK7
dS6RQsMyP0y947GICBu6jlQoAUFeXDvknr8QgGd7aHSaW6mRUCmeFYjOe6wlnkgg
9JlvI7drx+Xybvpp5EoKdSLJdnVUsUA12U+zxpWJJCnZLZpg2xCGRfUsJEdHtvba
znI81od4YpqWxkdwnDNtUYuOtd6+u3P5L68VRpPhgcTOIeYevTRM0CX3kd/d3inH
XUTDtEaGJPYwnl2S+jJjOGHMThZeT4IKD7bwUm8l+F+9QMdxHAUctbseCcie2q6G
Em/doej3j6QRbBFufWYVqDdIBbJvz67IjhpWu/7/MxYuO85OfbeYNpeiifX9QS0V
hCKrzXtTHKZ5IKfNoE1MrQ3dbt74DWDoQZ/CABr2BGUkEfcY776StVttisT7M+Zd
xXJDVLNippL+Jde25hDNvrEaiswLj4MjKbt1ospOd4V06CsBi1nCxo2C0W7aPOw/
kvNh3RIJg7RX9ZCnqSI0VEwvpXHzD4eUc/+5/32wIcMApAImjYb2SGIa+6ZwO1F4
aY4oA1s5it2xlwT/SBZmO8iiNwrD4xwtq/hr6KjV+XWVtTHMlgpWh4CrO/QvEi6K
zfu42S35z6xF6hAmd2HX3aoF5dLnhyF7v8v1UNfiq5mHet66wUXCvvJob+HV1JNz
KbIK8cC9jbYfWImk69+l+ZKy+XKQP8xe2kccM3wvlYl5ziFpB08+s09zICKyuMK6
LZmuZIKGzNKFWOmWvszd+PYK8RdSb5QtKmwmRuuKYL8a1iG5QTep9AzL/cp2hdWM
kNveljyoSAeN0r400TShQKLeAlSJrpsNoc49C7vquxL1NcIEcfsdFHcxOpv5nd7d
8bptXrgFF6mM8NOZUKO+SLwTDEJ85/NG01WfyUeElCW62jovumf9yOLO10DqWN/+
BSmdutCtZZZYxY3tYI9h7BviWUQodL0xfyZvxQT7SK5+VhEFQMuUz/pTK0rr96U1
0txBV3aVhYRvfoHYqpvuejQ2KOcRWFwWoEbgWhUqlbn+UHMy9jqpcIr7SZK4M2xD
BRp4xfOe1ZR39OzFtoaK11qYPj6ZLmVaNPAWNnPHnWjp8toUk+hdXLgkf+tKON/6
iPMI+EbrmLC0BX0h4yMvIeS3Jp6BtQ4k5VaCjJrCfNQ+i3qKDfpPsm3fp142Fsrj
Stl8DVrWaea5Svj4MuAZG9pNY0ieBHTqdwy/S5dkIvTvTdqX6DjvwYvVn4VVxty7
Kffg2kqwDYEZ5FCd9ZElYGJN+a7PpGtAfUtWPLwq7lx5rYV/M30ax4Ne8Ke5NZp1
/UgPifOQ1faOgG4fiI+BqK7erK1gubn06BGgOfP3HgPtXm33SORQTC9nz9CwbvcQ
GTKfIxFpYADDP4bZlHc0tno+W6r2EuJdDZlDTgjc+RbHdffHybNQQ6G/2al7+Emx
9xiLn3L2xBL/DB0s13hYEjVc2VFbqAb+nECyMmhTdacoN+dT3l9Eg3pefH1WkN6Y
hO9pNvoph//SoFJXPjeaLDt5Rdf7Lwm45hdBfDCIbImQ0otn+yBaA+SBYJhveFbN
2RFOo79FdcEl/xeZ2RHSJyt5GIHyjoU8AhZxgPRDQyzv+JikmFT+S+5RuWXYLH/z
2NUJ7vfkcSQgGsoQb/Lv8NuaOE5JOoZ6HQtTfS29MFUQQCAt63oz0sGMiGsAJu/8
1GkB4E2H2+fl4d6uG8oyV/Z4YF457rnonyq98/Z1KX/JMTIuKiW5zOBv92Cj0qrt
K67sx2J5sEVZuQFN3phU4nlL0PNs/gU8atPTOAdUl3+/4RM2JKEaOgJuWAiGu7kV
K8C/hRVOkqua4f8YKDTzSlcjqTjoQDCjl0HTe5o9GiHaczqRT7oLtYfjPNOuzAeh
xvV6lFqNlJAAVRNQkZzENFghgxsb5JMLcGz0YWw4riQ2WjzzqNEYeoDTAnvElnDy
BnX3mfHsHLQKKFxsinBWgytZlsV9vwwyNuUJMI2LxVqcQ+tBRUNio6A2t+cv0Tz4
xfy2HMGYQaK0+8GJ2YwASKQlwkdO0WrG9/eNNRT39lNgZKPO7vrhGZBNCQIp7Kby
UoKb2E2z4T+R6V1t+LN8wPO39W92Zii9bkIYnnP3Ec5Y1vwwLxbiiOyJclA5BUU7
odW6DDyaaadXJq1ZWh8LkWVB5XCkp+P84YAN22yqCM6wEluLOga03hWe8eZYA25m
ELX+xqC7QcDJgjUGTvz9YPEE92T65CLxQILFWEZm4knqawZRpEsx7064BIq2nf66
Ku5OkUJKMnFL/iw8+HxeCYqjpTIN5FTjq2+ST+rz6NaF71zxOsmD0+WancIBXlhX
0/WaX3DovyUqxMNCB12Pwm1grdwMV3akOrTVd4xQQF8YJOEwUdHm2G6UzBxsUrJo
R6Xeyaw5ALgC2ayYb34qctq+cOGMENXoG4utrXIpYS35+p+VTLaIzDDgxab904QH
G0R5KjmFKTpxeMmJTdxXIYDLaRI6gUmeID8xRz5gqum8FowL1uq93bYpEUEpzzOa
9/kB+9BiGvKpHtKusAJXgxf7vc2FZkTdi00CBNCeQeinFKpz/Gt1q0/+f1/+FsN9
PEyCKC/EjG/4Y34CI6u1Wf8y+aNUb9XBHtcJd8oDIIelhDMWgwrrLk0HuKdRpI75
6teMWZiCtUQMqhlV3y+Be/tg/9wDRjJ1f5GyEyh724uvciWNNXhnVv/ydDoGXXQR
O9HHasS8TOlEL23MzMDIl06oXti65tDsjSxTJRMIWErqnnIrx8wNyoUaLp6QY3Ph
YSQzfIggq6VBjimJLj5nh05852vD4zzBkm8VETdRLP1OtfVSCXICrnnpQ4qMH+QF
ckWHJeXrGpjwzc4OvseeurVC82O2+UQqs9cp1abz1Kfb6HG6bNgNzOR2ZUPYx5Th
vX0sMLbhf5byT0Thu15RHwl5+z+7olOPtQLgEGJyMOcDKfh4VG5iVKh8ud/jCeaB
gKzLSx6bQK7leO/hGbKJ/WKj4ZNdFr6M6ltd4UYdvKRStc3ieyhueq37Z4k16I6w
DA3hMKUGIqbIgrBoODBHjkb+JkAmjcFf1ditoFYQeEFPEYpRB2WgnnkbXCbIWFHR
q0ugSgQ3MwMgd9LSMJDyP8lf84pGyKRTGIZJRvj7Xyz3NnXvGC64sikTBAhDw24S
qmrjIW2MiOh1nhxbiJYZKinoXCRo+auqNbVdK+vi2FqFzEyRZsh6Yw5+zk9IA+7I
hYw8RDYibWA/QpNOEJyMMepRidgOHagtFIeS5ftQb5lhZistR05ByYHaR5NaYpsV
gSsiys8NMq+3Qn5RZYJXeaZ6ldyiBYyZ51kmsqJKod+WJBPd3zdVIU5E1YbRSqNH
UGjZ/8ilxKqfJf/pyl+ZFHjSC5AewHkrzRyUV7OMtEmGQ+NhRBfUm5FsqQm/fwke
EVa98q6zNPbY27xS4f5aw4rATkNKvc4JSOpyfTejiz4hMuuJw6r4KuejSAT6FStK
BkfuzMcTfwswi3XpOCP1tG/wX8wmVfSD6nc5onbhsUvkKdJO1JDpVNi3fZlbNec9
mnJirsG4FB88R+pNTtF1sWH+4SnRdT68J+yzeDkeEGE2at14aaYgiPhRaYVvSUFt
KXj1eVCWq0tOOivAhz0OctbGCyrc4OAyMFSeFNvIIKa0WBEem5ueVWGkWWudOzvz
JvWw08WAWr48Ue0xQgbwKrpmYJdYYLMT/mKeevV9LXGXMmtu0J0fe+1aL35iQ5IJ
z7CbJhRq0NVZMs2ZDDNYf3PJDwXazu3MltjXbFoEfa/3dM0qlBP01gfIffLX4xxC
dhr24heMmcYS+FMcVOYT9BMo4o/vnBIzpj4J6klDb0uEq8KjaCv46EmIZ5BBJheQ
MJuGxgtE4PISKtNQQ5M4yP44VRrGZu5gi5MnaSFYSldim/3pwtpy2r8UN/fgFuZp
NbnQPWq6HLDDuAmhS9MJfrWU/r8T1rbydBhT5okNZxIqBhY5LV6e+E0nrQ1RKLm6
br6dooOQopKTAhszdpcxOBA9vx5rG+UkD2qR9r3ZOjyHdNHRxw/YSyt+KBWyBH++
puqVrn8thQpu8uDIbu+bi2zFu0Y9wqM06FZlqGZ7zYIIEI78W2feCfaYprEOSgB6
kjr6V1p6nVg+faTg8+gEPvQKUL4Hj6yChg1bKcv5qpz+5ryfHltpHTZ25D1ZkDNX
aTehA2naT2Qw30tYQAJQQtgnV8Yy/azwFKNLfyfRmJB1NNX2TCsULbBPlGxebKLb
aJ9suEMr2eFk/b88gplBcSt8iovGKsKcHH/rfnk0lSmpxMqOz+0eCefb+hKaKeOj
EMOLU+ktEc+rTm0jURDYf67O25WLA2yvjFiyDyOYNvThDP/L4HAcsJcQ3xOTLkcp
gCmVq0sE+f8WQaxgD4nCPWgnr51Irt2goxvXQ+Pscrahi7FYQG493n8Eo0X5EgaL
Ues0qaa3nVlqabez/aVFehEyrdDNZNmHxM61tkescCzZKcGb5gbpVISCPRBDQIFp
cynY/FQuB4J/1j+Dh/HfqiZKfPu9lhCVMSDq9cTzJ/BN8rox4DDviNwFIYwQp32i
h1ujAX38bW7pRCs0hPclO0Mv/dr+PEikmUDFeMd5eUKp30/cbj88hta93iPVgWgQ
e301XngzHqkdqMgYtEf3CwNauU7zW/JRUF2WB3P7pdI8dU3MQ0AnNBljhMA/Q1h0
/giwo4uZRDKP7zV7Q5/RCSYHWRqJkolVbLwX/oliCdTGWhO2SZM0OXA8n5oCBzrp
1MSbayjvMhAuwXGym/GZcG2DgSv0Rqo8j4FdfZF7iJQwgiXhLbTThK/EMBvrEwsC
fdmJ4/+/JsIkESUiRiNGwtdppYSkp6VIIfh5VsO+c4IcNJu1dI6qsVZs5gBq070X
/TVsGS+YajRF3H0haN5DhCJcxwu5w8YLqfId5P40UeFhbHPIym/368LdcoXZ3GrU
bV8uz7ZGN/AQJoet5Ef10LbRF0ohB7hJqBGmanCzh020cwJszc41rXFQBTzEC5rd
WfdqlmfAo1TSWTAuqEomC/iJ6VdXJ9eGGpMdzVowjj9xK8L22B0u9Rsw8LcKPhJa
cTrQU7kUvQicsKCUxga5a6WrR2ZAi/tEbIBgLZp/sKNgyEB+ZsJrZiP4Ha25WAlu
uKhYDN7+y2autOd6g3FgaCXuj/gsPWZiAazV2AlyHEfnfwKl7XZSm93dnSsmQ8ga
lk047TA4AACKB7HYBFfLH1rFmmjn4usOWPKdC6WagTmDBO6dcJ26HbCOIwDHitF4
3bRuu822baga3MunpJarzLSfo2jNHSM6hrB1MUL1pLD2LWIMG8zMz62bvf6jOCs7
Qxop2dtlYTHPscpvC7U2otgvtvcMe1rWg0rFrIkZXmziXEkgsis5bLRM4941WHAC
yC/aUKAnMPJI82NBljR23i8FmsD5YHW7RFuUBVRysrZBMKAo3wz2GtTpGaht+oiN
2D3JTFAE8SJ6CQ6dLMUqO8IyZIPWisvrbc5VYMTf0idqT3Y3rFZj9CpWo99C81+A
XOwdyhLabPvZAh+D5AZV83fT84d1KWweqUIieC/93hi/gpPNBl7HYd3xfB/s9dA5
FLYVMEzEZFzwDstx0cbuoHpo2aNuFzP1l41GDmFWvWQxYoRFDQZI/aHWU8n3kxO3
pr1DGx0VsGWFfoydM6xwV8gxbXhAyOYd+286S1/TmBpwJLY348h013xqUcxZGhWE
885CM/PBA0JFW9WMO9lG++dLHCTNNmpT27g4p4usvrOtvjC0MucETXMzwUZoCBjA
n7mLBjsJMULHiw9sKBc83wsmyfqkkQRZXjmMnZf2p/KrUNmk1B3tFJUmXETwy4Kr
a77YaaT8APecpqaY9cTCkhG/TRhHzsXF3mzQmaeccCz6MAyH/ipmM+wfkUjJ1WQZ
qdx5kRcWet/oyFLtGXA42bZtFFNfGLd2IN9AKV9pDfOIyDHm7dbbrxAc/rPo2blC
p1Mo+ZLAB88Nyl6bCjECsKr9r9/CtEbxX/rH+FCaCQru7hRf/IxYCl9kW1OJ0xO9
6aXHmodNfR1dLi1g4PudxegIs8NOw3uX3oc5pddi209rBx7ryGh98gJ2hlYvG8GN
JLvYvE7V8pUjiKe8aBu6T7Kq6iu9kWuq4n4ipf7IBADYvJCkoIMtbQX15SjRa63b
a4L1oAhEyvfXyfddOzlxsHimlFueQiEA9DIw01Oru2kX09EG84XhZ+ImAmAKw9vH
klXjeN3rfBrzO8k7lVRuxLX16sD/y3GVt1ftioEc6BvTUiK+bwMWswMER+tcUt3/
h10M8nISKZ/ldv860LulJM06tVHVuJwMNaF/eqwZkw7XkHwbu/VRrgyg0bwi2MLs
wriGqJGXmv4XWrPgPhjMbAnsT2yn/7E/pgBj+MM0QmFOSNB2l4red30an/gfkt7E
f4bBpkSpnKP2qNos5gX/MgL6Wt7Qilqi3ZVVeYJ8m8G82cqqZH3CCbm5Ly7IOU38
aUPH3ac9r42TM9zHmPcNUJz8QBrTyNFWzAAZEMMtcPq37T3vZLLZyBA60l6kFJlR
4KXUAemoX4Jy7yB4CTdejs2wj0kuV3PsL0j2GglxhqQCL0SRa/gDmCaNQ6Yk5YH4
p8NsGL781hlTXtXj+cVC4VAxpcwsz1cyN26kmH0Sp9OdETcllFeUNnytcNLkiPkV
Hj2za4pg8Y2fmoF0CYr3PBJu1uGUYCZ9pfMouX1x3n0A2lN6XmL/+CoP7oMU75Go
VvEYZ8uZoC/O/VQeaue/1ZaYy+jlVhf0fxRQP4YZromRhz+39o6tpBBnOmSHmvHL
f8B2QwWUQcKENgm7RkLnHfTCZcfeN40c8XVEuKW+w724RpkWYLMUuX6Os9IjfiBE
8mdWQEqvApNSn9SAs00B4dwf2ViGmhG0EsdsER04huUnfnSVb1pdmNJS4ngRogVm
Z3C7gIPiHpKCuepqmehF7FtfaYczqpyRZOEo2vqtiGN0EupVw1b3fnAmzYPr7wUp
2hFROR5w8IT2eTDYq4W0rMFiNTXhiV77MwPvIzVhnGdQ2T23wfFeh5B+eDiYfdxN
1WW6ypmAw7KrHzUXTIVF2g89Ro4mX2/6WC8CLpTQcypwhALC2hvBQSsoAjvsORI0
KyaLSMbJTfp/xriESsQYMtZWxNm8zDQUKY6og3zJ0cx3XJvDhSPf4iTldHb0jvgh
5BHgtID30T7GhHCBfVsGT9Jv7KahlM6WYPvtH3n3IACOXGEE6NYAFmZ7H/bqcKBh
DBkiDlwDEhuuw9jUX1qJ8I4QgCpcKVgBD5cFqUHWSEXI9eMq5chITB4DvtBsEQ30
UYCBXIp8rJzpv8RwEZfqEfwX8JVAQxTwEkXUE0x84z0h96skr1w2Py71scFCTBNT
hgN9okjh908p8hoC8U6tJywmGRLZb2bndiZDFKVC8Oz98x05RfwbAchApKbxSg+p
aTwDseCAfXqa4V/3tSK68LFmgdoDi5smia6dBW0qlbr4PZM2Coo7BzMJgPxCL9Ek
Zv98b2cWt0vHhsl/Nx9DtbPEcPxZj5Rq9qJFjE7HNLn8L7hgiOeFBD7sNCSGotBt
BZZryBtFgoMG7R9Mmi+wTa2paJh7K6y5nNb+KaeaftxPaB7TuNEtWuGieEmcAT1F
8sKHrulYxqgCmUWpj7gbW1bL/fXtxVcLmxtkLCNAdn9VD8ViehNkOh3ruaU4dh1d
XNCQSMFPDyodyaBHHn6dpwvKx62ywH2PdPGzFNWj5cjcaGi+eyXNjpy2qfTiQsWZ
BTH8qZ5ePQoVRf/pAFfRDj7AMLwxCQYpNqkBSti47sozgb1/K6YmI8fV2hp/AInh
8UNL/uQ9RdpLYynAmyw4vNQfLhQISAojcIXytAVTDBhnN2CXpFqXbZizzkzIeVPS
BMkfOcjXcBnYACfWHfefLUf+uDjeK2V8Sd+eW74oe/Sy4aCpbgU9hQ+4XIGKDqZ2
wlxSDrk8Zzl5zv3szZh3+LXcxZyqSXU0JMvz4BTjei/+aKdYDpwF7k0BNVKUkQj6
V7PcTWq2v7+NOVToefUINkn9QAaWAJSVw2M8luEBlXKVtxEZnijFv6iB1r2awGMU
QNYjz/iC/s3jlsryzl7BN/HmRMJ9ydKm92JgE7VJFyg3GiYwV80u4iwrNOaD6/vB
Vx5bgux+FWF15tsOIjY/0WmsbP4qqnaDxGJcDLNIQ4iqAKDx1NJC++/++aRzk+iP
2f+lDoEYpycJn+RZ7pWrQFo1/ayrVdKoKpETTC3wQJEAf1tRmFFHSPgcj/2K5aqJ
9PJUCx/8kicDkf0HE+O0vzsWtrUl06z4UMMucElHoQ4IRaLL1tU6DjZSXqubykzP
BNEkqkfu5poZS4SGhM/hm9tuN0rtiysRZFFTBRJWsLkiDx+0t0CiFP/YZ4zrHSiy
8yepwB3U+SkSL/+6kzDhkwOtZoqP8OtmHCXk9gS+Ds2ellalRMpziEeFNNEJAEdh
X9LSfNuUumdBTBr4Z8O6/6JiPvcrM9HFgLdAJhM2ZSVP0SJlcKE2YV3wXfetyvUj
ZZoRmoQBKp3iBZsvMJytnhXGs4NyovrrTTcljsUdY/E4DK18su+oINEaxoitEWuf
yXxoRrEBXk5cHt5sh7T12wQTO8L0sPCIPeLs6GTVBxhE3jCOGbfYy9iF9H5kZ6r+
qMdso+klX9Usnp8id87GFXs0PUSuq779ASfIEMPAE/39xbrHt2FbZ9O0mvU8E74o
60PieOMuD7oRaSywyabEbztExEKOkYr+jyv5lgU55k3gztvn4SqGmzbWa9dlIJrs
jasBKZCniLCVO+H6G4u7G014G5Yd5bWovqGYKgnxUKJMq1lxaoJz9RS9u1HPByNn
vHXtYNsvlAAzkt0dLa6UdyrUZOYnUUAIZ88FGtK3QGqSJ5rk4X7fEgsyUjCU3bmF
uf77LrMuN9EMv2Ko8mTUuSq4hWcw8kiB6lUJ3bRzWaakbAOBrRtJmQWbHA+HFq4N
q+vAYZ/uVRMrVxz3E3Ev+ohHzaDd0j4XLF4a43jJscXwLDiyFEUTYV45Xr/mL/NE
gVlB7xW0EtzImxlrGGM0kSymvC4ofJgfaf82NbI1l/czG4l6HDmaD/l38yii96MD
CLkgCvhU2wcMkUXa01B6ZFX5PVQxEI7hQCQoCCxPfJRmlqsWSsSe6o7PGar5D2bb
lOFUemyc+j0XdZo3n1tYU6/rbOSa1C75z2ytpOluJLUHhj0G6yJ/lUoPiPInZuzH
1V4l9r0kVxnctlrbGQ+I94kLI0GQAbVrbFAkZrHqKif4QJSxUmwVfTSqTb2GWH4b
SFnSmHp1/xOoeSb6V7B/x/b9EEF6eitBpC8TEugQDJ0f0vIxU+mhYd8/qdm/K0yj
kQzxWjixaQleALClRN/mwConHQw6M/qolfuTMDBsz/K1EkL6tE4ohRTS5MHBo8A+
7t8PBSD7SQClpc20Om/z75NBNBamMW91nG+XWPO9Ix4HZy8g59kLU1Mp7ksYW7Xi
IgKBqsRSkvguYVQwQhxh8xW4ojo3lQibsFnMLTnKCx5gW8Ef01fu+0NCZV1Ffiym
plFgQ82BI1bOaL7P99sSf1K3uaL7WaPzoC6E5OHpTBRk0pratK+ijvRutNubO0OH
dZbh7o2owyrQ6YbwkfAseRW/PzM5jBMfYxhEhKQuUvLrIoNZw5tJS2a8vIwix49X
tEXVhO8W58h62K0/nHBIlAys4EQ2AnSknLTLtx31DL5+/0rGiokrKthbohv0mjre
E45M2SS+thZ/fhsNgreC6vU2B3vvQ/zIr6mo9ao5ov2+ZcOe4ILq9T3m+Z/OHDYE
4DvtptdUcCjNR58KcNFEHgdkJygkt8BT0Ff+VA7Wl12QqXb1p2veUMCtimGXIpur
zlB2sr1ovwc8oMqYOnWkS/BWtH6y5XtYoyr5fchKwhx5RydnpuuDZ+1504PS2Bec
UONdUhwzcAEz5iKzKKZiab1sLDzTW/kt5NeW16cmw2pXt0Uuug+zeRZNEyFETUfn
HRGlDJEMmnQyLAmGGlZwEZJZCwBIjdYeczBoU+V3cAsNd1cqLJ9IsWzfxA1Yrzwe
8eogv2Yp14VN1tWs3JWoWiBwPNdIRVJ/XBn51gL4ADIUSbPcJUseyZosKGQkp6aG
PdbcZ7NnVRq0siRwsqctKoaP+/SXqF+VlfwliXI17DUcMon/jO/biTBz7UDNRrIB
Q7z0FlMVtwrc67YsO8I+16/E7al8C+D5GYtfDGT5rrl9h+ssClcFxrIWkSASCI4R
W9blSQ113hBs5xKwZYu90BCKY1VIC3NfJe419tM7RcJgzFmP3V92i9tthV5n/5nY
HeOwvfFzL6HLOaoMQkPWkgOfKBAkO+7n0FAuxaS+TyoZtdObKtcf19oYqRnzBLIv
FWiLXDPJJsJfkfXlyB1gotIn34I8ezt6T6erQDBKO8mIJ1oOAJwsclmxCy0gVhuQ
FlMvTrHIiif+IlibCQ8JjFcgOV/vnG7vlCDWvCG2xgCviRlw8m9Ej6MLlIKoICmO
0CV8ev/jKqjN+Yv0mYohPhatvCHCMthX1WC9zJ+H+lOSIEb+SMxDCyaZLJH35xs8
w4HYfJV3tw/GDP8yVsEjm7MqSqZq7r2fh9ooyyBXN1wy2dVPLHlFyeVdUlmMCcRO
D/h1uN07y0RzGTNRqHF6Q5Wby9x6qjUmKviCJ1afMOT0jgsZsrpTgF2RSEJUSOwA
m052InCBRY3Rbl0BoWETQP46lSe40w+53jc1F4Dd3B507Z8YVE/kNfT9i4Ihgxev
20KgOIWtFXlqGl8Y+2M8wHpo60zawXmXWzRfOnRBkKFks1C1TYCZnJj5pV+kfPYS
Fql+FwgbeccyGE03kEDl0EAFAy6MXZBmKhfjwMxaV1H1QUOVKoVJWkdjWP9sMPQE
tjKaGlx0CueowE2/FZnqq4EDBVI1cHgSV8JG1rbnS95+8eAel7IPg2d7kt2aOI0i
iGO4NzVzFxIwCb6Vqy/JLoBm6G39CmCuH4GZy12tRbhtjiUkJA3Nvb11mgFpIkTi
YKL4nBAqda5Oi3YtGbkMtFphThIDIXCQdm3AWw+DJbaWBFTCAeSFiG0JC+SFuVXS
u5UX/rRQWYEntV+MBg7u8Q==
--pragma protect end_data_block
--pragma protect digest_block
w+PFO/aXAV5atbUcFMFA5tqxxlU=
--pragma protect end_digest_block
--pragma protect end_protected
