-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
I9FS8OBjYA3NKk+2Qaoeq6gZMhYqBamIqQ3pjJoAmYZjHztDmjj/FLvd339n1Iqs
o0GbDtqy3zeVqtsgE9OZx4/V0gM63PyAyIZ1BC41s4nhQAm7k3n9gVnJQ+4JSPaL
NQvM2Kuyh72w29SVekY0JRhWIxrj655azTTU0KjnIbVJQ1OkUVfInw==
--pragma protect end_key_block
--pragma protect digest_block
Vb6QJx/lo1PvBuYQCXC3tLkfz+M=
--pragma protect end_digest_block
--pragma protect data_block
AyevtyrHTvaLl3OGaYxMWEs5OVtugtokH6jsFDNXwJotKiNKVx7eRWnsNjhI7Ydr
0G665cequM2Y0tV07o5FVHS8IjEy0PjSZNZw7NqMbbwlImzYTYLtuUELkui415HQ
luzel7kJzdXV6GciLp/YNK6R5E3Fr2IkrLVg3t634KKIF1i4eBcxV+/DnlJ0qOmL
CNQvKkL2S9WAh3op8q/hHsqfRNLTO6cAXGENtbAl/ExvDVx4huUw+p9ZTdyz3ATr
vP9KRjfv/OReherGS2rJV86lP/fK6xNzhRCS4cYNMEBJNV1WTndur0QCO1+PKqu1
/LEEHYD5sCnXRcjbB1G5LTuMYViinRZ3l9e9+nOEkJjlIKzTiN465o5TPzeAMwhJ
sS6AyOgD1SK4oDk4BIRLyxyZFW+EmtNc7qQdeJCTXsOA6J3ylkmY3TJNS+FbvITt
Xypj8cTPTkY9GEZBLdPwV/MICY/XW1UlmZOOZPgpyMiXqbQ9wOjmMvPF/NMERJQg
rfIGZmH1NJYlQgXrwYJdvP/PxWHNx7HyUAM0QGZsj8uQ2LEenoAlB/IMJxkvXiK2
HWAG6QzV4mdgvCV0TNdBLr21MW5EiyixATvuoqb+uTF5U+2Z7XsJBPAWLc7sh8mu
+TNaJ1jr0Vz3j6+FtpuTQSt0lmjuQHZcSEkiwFEMyqNvnXdeKkhH6/lK8PONMx3U
UjPsbkW5+XhP6RRRXyn5UnAuDzFGKPkxVLFaBhiJPE4Ti6ufmilFqW8AEYGFvEXs
rIukX2OQrHdY2nIqgNCvkfQMymwWQxyjGLOdAJYFvuvpoG2L/zP4RdwfVThmjCKs
UGZccqDTmFExkmQwAFNPyP6lKxBU82k8S02R8skgklJJJpHeF/EPnhfeuevie4VX
CeAeInmI7ug/VCTvVOVNXEi3V6sqym6PPx8JVDxvqDZHiT+X363GzFrOIXJMGVhZ
xirF+UjuP9ONMLNCuaAIzbHerx/uy7fhgamX858WdH73nmydn4P2u7ThksVcO7fY
XSfxpiUThNu5rBvK5cV694SnHk7fLvNjGssuqlOCKSBUd8DjeroI4f5f338lRpUz
cIwT3bOfot3kPTFdp4hfT3u50I0/0oMkGeBgIyx3WxxOt2CBVmkBwxwz7/3Dmkfy
J9HR9588bC8q4S++V8ap3PwuEb9mRRO3+skAhMbtpoKy/zI1xVSCip4N/o5w6dbn
4hMV90MDDCQiTikUMjRyOcGqVDxK/IJFCrBSAhkdxoQH0nkdTQsam2WJTG+Xvwfo
S3a2JQ0U+orSdPGJiNQudsZ8o8W3XlU9ZWO1nClhLgpuqPmEK9usxR/q5kXIrHws
8Ja6y0/m3+hjadFuVb8GXyxZe46QPWOpK3w8h5lP9Yq0sooA9birBfdmMsVQdy8l
h7ls2AUoXehNZEYINrvrJPGEiYg59tYa4Ij8ovn9SvwdujwAHQT6Y91iR8EvzI3f
fDBGymuTj0ciJuUuGWnl0DOAmKHPL5v8KYTFvmBCUpYgJ/QU95Ddx/O91QruGJwu
df5xZhTyQyVVcUEWNeC6thl3rrC1l8lhTwdd79zBmKGnvKbD+lpeJ3dWCLUFNu8b
Zg39IkozsL5XjHfMMvx6Zs1xXi8GiPpzu0iI5TC9lAG22t1y+uK208uwsjJYh8i+
YhjJuB4cWJlE0sz1fZ1qsTmYdOrGmiNuBJ4oO6624M8EbarrLCNk534f6OKReg5S
bfPZSzCiTzBTLfp40X7/rSCSbPW7sZKkhixPhHnG9VqKrVfXRBWhhdJbrIl+0sc+
D66vftw1NkJ58p0BoDV5DBeTEuHx2/q+lotUefJi8few23AW4P6ewZI9lkHzXXtI
3trWvMMGGIFYXWMSBJCLl+waBcyTqlvh0N3QcgaQpNoTfxxKivEA+XjZo4IsiCzb
xe06q/R/XTgTAMzMc3wI/t/PtOYehMxcE8PwAWtumxfJnYanHXAbc0RT8R6HMC/R
8b0j6QOx5nu6c/h5VNx0EZW2uYC0oACnZVxzWC38optR/PGP436ILeq4bm91kW8O
Lh4oyqG6SM2pr+mgmO3l7bV+lzWxMs0ePzcf8d09Ptm9ojUdHwpnTKH2c0/SThtB
SFwdob9tWEtbuu3z8UixtRut9WZsZjB3vS8JNxM+F2k5+YfkKTakaedkMm9fk0HW
MN1TFDp/en77HT+bSqeyUzqkhSmfQLSyxbUZ0UONveJ3y3Sg4Xl+gykYhCp0swA9
qcjJzBMejY/y73crVBO4bLLznLmrIMjoIN1blDSUC+oGEKokTT4zNmaHEdm/JhGC
tRkCm79+xQcUWQ8Vj8Sf0EAIg5PwRwCPwOZja49vm6XvxQYX98hRKFPZ1jV5k+Pk
GM14P+lx1vmXHNVLZXvP2184iDu+FXGjt4ks/5YdDCmt+/RY958C3YUAaif+K2kH
/Zhenu5LtuqEdOmVG7IkuTvGP0yjQv11nAUlPXerzn27tmpgjwqBdZaaTbARbzMe
Cy11kbKz4fouNSu8sHGyBSIXoGZYgYqZfAgIZVMGcEWpRLJ6gkxpQNX0946DXPK6
UPNo32Kr4YZtM0glvcAT9XAwnX/SYQxrWdtx7oy4hSVO0BmWtr0agWN4Fkd8J7CA
dr7OUARMpalzvMtfhribTiSiv6+qOZHcQGnTJlabLiH76Utw2Lq8g1B+NKhJjeXt
oO2JkwbUrIaIYbB8Vj33cOv+IjoSBG95ob/bhbHM0KPro23+We2dkLTEwflVz7vT
iYHwVqHPv92OdtudNASsSWD0BDp28rVt9ZvGjmy8SzdY90gd29QRYHwWmaHQprg9
c/pAucGeQH/7zL1NwNHvjYwJUC/ceWwC247wwfAyAPZJcKAdJX+kxj3+K5nEOQD8
u6/HwdTzZJFfBnDym705EkhiiuXtkbq8/0MEh76IjHqLQ9J8Dsx33KllAr31BPci
A4L8rYDvDoS3zmoIms3MWKhk3aVKL62YpkoDLNIN3LHgjfKBJVeTV208QGwXD2Wl
Fy9tlnZv6s0uNjRX+Mn+2zqilgp5TTNX/kL+1N3jJrEJzow+sy9vXnPTRlTwRK1w
ePhQYAwK/A4g9g8Fk1dshPyEMLxCq/Qk/L8mmgAF4JmqCsV9kMm5yT2KqMbD+vY6
4SOYjMe6deyWyuJufb1txzbJIixb7XyAiQz1kZjdJI8rwukXBKcJ747CAne+MN0E
VLrPayaOJ8AzsxAG1186hQMRjsFCC05jfhh/pZbLRbTO2lAGgWrBmSqNcnW1TGSA
lvv48u7J8QkX5a7+2y8T5nmsB2n95ZMjYlmm6jBLhdExIou2hChjvKK3j5xJwyhR
/yvVc+gt/YnsLLJvySRuQwBRMKb76hD2EEldcCg73VgDfPKu6JimdimUq3SL5h4y
e8qQAuiHPzbBuE4P4oGZAOelR+8IjSfSZvtrySIanICZQ8v16yLFoFSpWDAJitd1
gDQhH87gVWQ2u6mmI9cCOgxxhQqxgpB13z8JtZ1rRjTUL+XmgDb/3JZ+oamn8wdg
mqhCqFtbNOy//si117/vHOXwUygf/9Nij5C/snWB/e6jKnd4V8cgXDdurglE7ew1
PLWDLMAbcyVL5IYuLSaa3yXbAH54k8aNdKzyBhcYSBa1r7Mw9THRQMrNzgNhMaws
qKpWDS+umz17/TyK+jGPYyRu+2C4ny2K1c1tRPRWsbG7Zptj62IOXuasl7GNR31X
mWrq31l4TgtUSa2069ZKeu2g7MEbYxeJKib7ttiTlBOkBJlEeasCvZI2w1D91igp
4C/fXY9oXEl4xzZ8mSVKwDBx3DKojFQOdQHQSjQUm+feq2bphtyZIM0vZGLSQGer
6eAjkMxe9/UDQX+3qND/zaXUz8w38N1ZtgvuRXJ2YR1Gn6qRxUNVXBkc9/uZYaB9
uXrZDwOXrYsgwtl0IJR3f0l+0b+NfA2vG0sObzy3gVPgZ1eJKypqHkamkTpqF5nr
NpcsDyzKCKtD7CT5L/akHPmS2Bm6HX4wGmolKJWGEd6L81JNS5nfJNK+HFJQ3lh2
ojn5I4NVmnR4tq235Nc0YMaHbNASyvumAmigOU5TP1yJYIpKI8OixYQjCsLrtWOR
P4RjAz9q661AmXQfeKehYezYwNtEC0JiSAWbxLwyOkkDaiNJ9zHvRW+szSjeKETK
oQkOFKKxCUfm86ltHqwcFbG7WCA3FToEhEMttSnIofJohlzbJw/PcdhLfcTzZ+Xp
Pizt0Gi7/uiX+TWAK1UQw5po7RbO7GwLhjPk48LvcgFWdOtf3Sj/x+UeEVi8LEw2
mRREdToYvfHYnCcYV+0+1QcNQ0o+/Sq5OzMYgeEaN+1K7Tq+iDK+cbf2h3GfKAa5
fB+GAlIV+GWt0YY+cJ9G1mLgS/Cm8zh024IOeE5KlAF4UloYf3//yU9cBffK3H3E
auVL+yNat0SqiPZqemftVBwgmRszm+mIj8lQOuXTBHZJ0P1DQpp+S0VXHjALP7jy
gi4RmfJ0CRfomKNsh3j8hovWXl5UVku6v+4dwo90hqgzmgaaiA48b2JoSenJ629K
f3u9z07pkwXx3Mhg7gDLtNRhAejK8+Na5ssuNXvy+p0WLY01dRab5PiPJJdGY4MJ
DGK6sJcgYnNAapyXnwF6jdUYLVwEu6KpiP6QXBx9wPHxshIHXAmiJKIhHqx36t66
BG0d7pn7AaPfX+KcErc9HrfnNBV1OQ5VLjQfoDmcO/2Ps1ee7FCY4WuIN8DnlsUn
AY/J+LiXxMtgi2nzdZWOCt4z76XiEPe7/rf0GCHBOKxatrIGtnVpmF9jvmAsTRQt
YYx+odRO6tD4rrxTBjA/PIkSs7MjDo1NZC5mV4vFUDwF6c4idUFbggQqAx9QngFz
oYJounjozV+/cqU1KL5elYDxxzoEn2eUNFXTggQ+GimP3TMyD+/29yirmXGGj6/A
qCVXXaBbGLdNnZ33qMplyWk8nKHIUA/egjxOWPASJ8uyq9+j4KU7i7AzDtB29awB
E9X6WlEdgigt4tClA6Sji/M/lgwCHwORtaHQ4RqhFNrLq52JZ+rsH6Zy8raskr9G
uY03Kbxi5HwdzogQVfD3UBxDDBkgu0EV3pREb0pkSYs2gZS4jmP/mgT787XugNue
MBslsPLRaJBrA2/yahG+bMi0jv501NKDifj2HVmNhFwCADCyGPFrJfuyCZB51LdS
CfYct7UCHvBPkeS3Zssp4OSDxolmFbmokAxBKlTlzejt6Ryg4ushRdBkENrba55y
aG5AshyDTAZiCoc+/AlcyZMg+CAVWpGXGmPVyc+SWKFlaG+i0SfLMg9IQTs6iBY/
zXcomKw8REVUH/VQW4uNoBQcBhFyoTYukZ2GUxaRowPdn6t9fSwqNh/HfGj97O2N
fWLxpYxp51xD7uhOQeEd8to3o1rXzWEY49vMXPUUscxdzc9N19TzEmJWBOT7kf92
Zyh18J2XtFvMqyL0LuiskvIrYH1bZB3ww9VGV97yX2P5qA8sRrlzXur2UhfCaHeQ
cp+/Dr7Z1srFI/A4oGcbj6CzRkMrvWuxVbxxZVN76nxEMN1eMxs6QpaeiPNYbGGw
trBxm+j12kJr9WKC8qnUadzsE0UCYjAHwSAiX5UV2Hy35rIVHmQmJ9WEX/qUAbVY
D8VQog748rQCtbrZgYF2pUwL5qPUGF+vnO0Cj51vUN/eyP0g3TE6x9FQ36Da+37x
j/ohymMBe8dqyxLSf93NM4hhxlnnsWLE8figMQf1NV351D54BKpDIgMeFb/Mpi1q
Or+0zaPLArnbrwZp+XfMfOsFkgVwzS5vk1y90Tlg21rQRzeu2utiZgDs6Ne6mYGS
EsWFQC/t/ouQTgS9eHqVFSfm5xw+LyrELC2suLruo4O6NA2d4cuiL1GzLhUxdGzn
kKgazOc18b8YjpdGX2BVls1E0uubioFrP08rU7LMGmzKbtQDlhYiDOQ+PyGRG8aq
Z+YTrVxQ5nIYQkaeCt6DtyEqxAt1BgDqjSGqOBfaewQMcq4IZC3aQzEZ1Hla2IbV
Rms/WtJTaHmqHX78x88hlT2VXjAF848fhOI23ojAE9Fip1XqtSdL57nRvklOUk5M
cyfEccZNqGnvdvCS4so9uolm9RNo/GD/RcIeoiISBRa65e4FvboVmBYdPx9co72C
U4E+86kcUqdAdquCzd7HGGLfdYbAeW2XXv1mmuIVjWFUvGOH12+04Q+2I00dPmOH
65poW5bLtPqn8Gy42JtBkQ0Sx/MFXC3u9a8cTkuOR175u5eKx6+ZZi3sgDqDg4dW
iH8TRqLtMd0CLuAUO8lpAbZmpG8xJRiv/U7igmpeWQTmfrKMYH2OGeDCJn7RZmQ0
o35ilJYT+jDRXXDZhxSCcdFwxTNtZui6F6OUXBFD/3M=
--pragma protect end_data_block
--pragma protect digest_block
p9iiOv60Jl7glZvLE+fqC+vizn0=
--pragma protect end_digest_block
--pragma protect end_protected
