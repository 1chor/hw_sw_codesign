-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
VCKho/Rx/sZ+vaaY3U9eW0WgXnevUES7vLmOwkm2kUwamPFE7cVUwDS8a9yrAH9z
LI9Du8JuR85aXDRDKCUTOcM71aBE29b2Qy7OtX7VRUhl7J4v5QH4rZtkovsiDc1/
f9CTsMMeGmcl5+JhXGhYKUIfIvQXlpUfO+EEAaw9Uec=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 49775)

`protect DATA_BLOCK
8GwZ0yzWpd7Ev6r5BdrY4SCfKQLWIrzYzzHQ9qTghG5geG62ZO+3LwoeCX++cjVV
4BbE6p/ZUrJSSbvdlQwGA6ZyFp/mzg75wokNgvT0LtEn5o0MbWxZroSYe19Ek3cE
0EAYZqcPR3MQbNTnsOk4fDE2NDQ+rDuRV4VkZ2rk/sBpTaQW+n9zHTVv80gbcQOb
Q1Hf2QYPdgz1QSlhWezeNqvlv4Z9gCPwigE4Uc0TVAtFUBC2iXDn2EYR/3EXDWMy
3Q+KhkhLVMpeKAOrTL5aqRdWCBY6OolO2e9ZCE/tk3qXL/c8pFnm+Ay2eQ3Cdtgj
8Zv2JtihXjqREkSqIakrehSC1lnQ7VTGt72vRDYe35G3tdkVFg+iZmp3C2URM9ww
zjDn4zy1mTWgeVbjgXrX796D0ghZ/8molvUwXEwTgamhH+WXBXTbI426YZIiQlaR
NM4q39eRyNT2t6rYZ4U0xXGRnI19Fqs8a7fmrlWWTJFcU6I0E3D0OCDDf7FjpGHc
0uO0SfeiG3exb+gug1fAXQm5hE3Mqzd0pzAX/xTx/um/SsUb4Fvw5styieVc+imB
oahfQp3KAWcGNf3QcTlJCZlWOAr8sr63z3Jt5Q2Nj0vg1a99ZurtC1at0cS6ecLP
OhsoHaXq0CMKjTdFzLDj6bv2kX5Zux6G9FT6maHhNCmbYZhc+hWGRn1seXr1fsOP
hjklgKieUl4kGpj7sY3CaTV3jChxmP5mBYhXQJVClpNkN3VkH26jiIjJKzPwiwMP
4JoG5Cd2uw4VRReakw4JjAnJjYVJhKgESfavPZQD4BZEYa0DBXbwbNjh7e8W6rEU
XqZ/8LJjyf0PB9n/sxUFN61pMkDgC5nM4TiXAmDXLM9J/ado7wYgnbaKt08cf5GG
U/jGet0EFv3PZ+x65gWo8pr2vlfDfuU+5Ve3mDJHQKX6z4qT6a6j7mSGPXXtVwM4
RDTQw4n3F6NitGV+eP/vLdDu5I6PkhkldGi/1xSZoyrcsDx6y9EbOa/2PJepbnEk
n+yBOGVMPmmoAVD5IsB1LOgqhkv1kMNpgAQ7CCISNUwxndNaWQv6YtqB2vPw1f5z
QOibE9yZY1JBgTX7dtAeqjMr0ZG0mNFO0D6/eoE+TKDJ1hwfszFdeutgNigqMyfB
rse87AClvy6DdG+s5L0nvUIbMT+Utn3u3Y/17aRl0euwbGYqXgbTMoxH9Ivzbbtn
asbd7cB/1C8H0tc6Ht9qPDeTICrtN60pdWBPDKI+KU2rvRg5s0RJ3vPGhk73Qd16
wRLjqQ3ibYstgoFFk3AWNXqKi3cFCmIwJrkozn1HJSKhxidm1JvkFRHEF0289DD8
ZPVgqgfWG9E6/lGLYvBPKjDu/o8jvYVJYLxveGRDRk0l7a9luhRWoY89qv1+dn37
sEH/BqFswvg8Ebpavu9B9Kd3aRBHtfI2dJBmII7Qt9Kia8aOInnkLN/udQUJIZ6C
GkckCDcPorAnfwkjZWPkrW+Q1w4kHnwx0a9znFr0iHo5eLPjEFROlVNGvu0+/Uql
U/O+5Yl/GYHnZWyUj+3XwzllDBgx3WOvLb5LCJrK8w/dlRPltNOkjEwdh0cLFfZq
/WP7ZgkwZrYDB/v3plpi5TgI9xDFNtUZqT9RV/XjLCjgRJp0zu5sK2LC0RatvCIX
ukW0HIaP0chn4SLJMXLF8BHB34DLFFgvBL+dRFeOZjoA7GmDULv2wFSUXBgCMWjs
3TTnlFWvo3mk50gEEZzC+dE1Vma4bJXwktmLCqrzyl7Tysy5UfTOd+0zIq4GrGS6
gryInQFoynvul/7fVosl6vRV3h8HoQx66Js283o676bP4xg4OdcEiBX7uBLxy6rp
X0t3MLnj/C8VPGS/EhfSqMwlxWyJBSE7DwS8uObprl6WvjPoA8DtakpluK3xMTyQ
A1I7OoblKJzo7qOwsVnzUToE87bVKA1pn5BTYmTMGQf8YQLON9JpR9N33e7zHSfK
EtvRw3UjrhFkuEhuFSZY+5e6UlyCn5DdfX+vyj+tW7sGbsuLLuOAvOiohIPDCIVy
JWe/9OOJ4XidEzCjFuA4yNPnlxIQYUUvfodwuIEgIymOKzn80HbD3l7mTNO/m9at
C/EwKj105rLZgffuh7ADcxzA/tZxwDMK0KZbxHiV+6b0wSYQd6XjKacsqimEL65t
YeAm5iDigU7PpaIbhUp1fF9XkVtWpXX4UwT38+tnWJER6iL/R1eCE3YIGbu0HV8J
BI4jcK1Lpv/0MllEFLyl8t6/LqYcrStDMO/HUe7TCCMp1AnZb5q5NeBhBTXtm2CB
ycafMlt3KFROa8DMjxJQe8s3CDGjFGzGt4bIuYHDYM+usswA3E4WpegTcF0XkZrB
Oy51uPy08jd2695ycVe1xuOSAHTEixxADZnncvqBV6LX99pLQbfIXT+T+BRKzT4x
8ZC0EsWPlHK4PnWbxlw84UuQuYFPZSn7vosfmeXJOqxXTMs09v6jv63aufwHYxM8
dLO/rfX/yu1uzH/h6gT6oD4daTxAJmiqNDFJiZketbQpcwyA+0UfnMYf1jkUbHeu
if8tN2jURz4YFODn9gso2jQ55Hxqnsg3RK/EFtli+ZO1v/UXATm98WofGnw22Rli
5DEYHSd0ygmRYrIGFNAUevORSXDuWyL3MmlnlpxKHX1/dT2Yi0iHeH3hBBcGpTCt
vhzG2yahYkxkr22BuKx69a+vgbmGSwsCXEyqb/QIIWDQQxbKwRJnEDms2nD5fRDX
+LkS9HX5kv52t1xvf+CE4jTw3WWRRQflvfOVnejbj+FA8eRyYyAZ9aW8PNcl4IU6
hCZPVOavhAG1RISbgV4sfjug+n+R897y3pYwKiCkG6QuTKsBTck1q7UPeaC3ayL4
7mvyIIMe2QtiogbH8C3ErVNbRbgQU6xGs7EImVqcKsKSvIzJB8qQSjYdlMXwSsRM
MR4TSaIFsMeAyQrU8AR/ySgMwlPVK7MYtbHK9H6VjaalsXgIuXrAQCqkaCRYIIT/
P+z/jJPBJ6v5MOf/yM7LZLRNpYFtWF/T5VcgBY7vkmlPEABoRx809/Ws3esmztIf
l9msctJ0JplZ0rMvKJvri7FFwLvB+DDWr/8HnXdj4W1b4WDTEv4ZC1kecjhhrBIM
ojQbUOd58bnjI1Qb3KB12j0OWcKHb9Co02+fUO8bYZhkWUX4D5M68rqEoE//q81y
2ynAMCT6Fb23WR2xqwDY6ZZWeVVKgPgHnWqF8qB5S3dhj7HD86Yyk3Q4lJSyWOXZ
uXqpCkFAm36AtQIq+wi2OK1qpp8XJxPoLxjKTUgwiSStpAI5Lr54midiOzrAoHgf
ed49LR4/M1H2j5sUAPBfvkj2BkATKw7GPJ7sQOvjAplFmBumeKz5D+Y9pUkhA5zI
JQ9dDQegjWcrsrwStPLWnD1mOhHv5FSXFEp9FyK/bQAIhQk50CzfuPRTrS8BBluH
dX4lxaNDxp9OVy0+ECUhYKxJXeXOzl1JAAAGrssxVkOskys+KR2MUI0mmMt3Eaqq
JTm6+YicxkHXAUvjtYm8c6dkAvM8ItQKDL5HL0WPhggWUgS0YTwoLv9xx36JZSa6
Kpet7lBOWBWLpqbtkZeHVG/UEdDKE4AW+2HtLt0AwJzziajd5cw3ntZFRy4GzDn6
hUGCKP2FlOmd6HZ8Jt7qrVqxaZKXJgMZXLUuk0mlP4B7JKsFraC3noXOWy9U4KOp
U/Hbb60uYRPfl7gk1qXwJTzs2i0BWDspJ+GVaj1VnFCGsiI0D9iLIP7A2wP7mv52
ba/XOc7VJE+jTf8q48Y1YpQfgoyaMHaTIbAnX4wcrAQWqDwo4WY1Z3gojngsxyhr
v8To5NSEZDG/x+CHAs5ugHolRgGeyXCuj9s5Amu+8SwUjOBEUmn4poWrkYhePY05
W4y4Y8V19MqlFp11pvu/6aHJCVjTmhXN46YFma1DnItLNxZxdU/TCXulZed0gzHX
OwdRx9wg54oKQC3nRsxI+YQmz6VDda9NGHFG/UmxmBcWMmL8jL0qcOqVKWT/fO8W
4dWE0hM3X4NwHzifZqltHRn+DFepfEjCwY4QVcvmGOhsLgjGaIqkc+lLYAlSNpw2
3efWilnUD3DSkdVkeKLa/akLahsdijWLo+b71Pqcah23QDToCkP00/vwPbXB3GOB
kTXPmJuQMmQq1eFvDmFPfLOtbv8Ep3xryagVI4DJdZbzBxK62RWibND/0q6CMQmr
FVaFLI8I7yFNHdRQq6LpK/FVXYuQVLDGWmP32HfI3FfH89sLyC+U3AcU1pFX4Rtf
dnuDhh/faNhN3w/G/Ce6qNBrGvmZCCqJQUNcfsg7pIlJ6G/AAi0PCBw/pW68mz0h
36FHKjSEKicDzb9ju2wl2bsj1fqQXxOexWqEDpajTlH5HCdeYwqbnLB0HXhcvUke
i71wDGSuoVlk2ZBHGmV3caHWUnVmdFr/LmbjfybSPgi0HPLYv2Gp8nkFqRkxUiXt
fS/R+FsMdUzZTPy2WJcmt3DDwVU1+zyuSOt+uKqBzgKuE1/+pvGJ+sYzjRgDHRTi
o49EWvyoJ9g8R2t4Ouq5kVosUzyg1sJkMPWi1txSt2M3/HrONhaxrba4wAvddSJt
u/CtI29pMC5wV4Jp+ZlgjmLM8gNc4W2xsF/MuL0R/lYz2DMcHUEAkMqq7qW2CmiG
giAJFmjlxKOBpwxqrLb0XE9f4P9T4yKleiMNJCfC+ZBdZmVScKyI3wPTrKMXTL/A
pTE/BUR04NurA07CjTW6qCYCE9vqYy0QTudT/648a0IDDM3ro5HXJib9AcXe+H1z
NfdyygH/9Kk6iXQfMdDEP8z50XBPq1ZShzd0XmpNfKnV+4cJ87CJqgZTrj2YwDsd
9WKnNYyUg66ijl6s1FrkTQaT8aKlvT3PTQ14hEs6nQC4TIYgCbf8V4CjjOZOQh4H
ktZfsJprGLtAncIcbJQ47vcEwRctjpDM0KdJW8pNJWKP0o/DgJLIwn5RuInPL00J
zlu69OhLou0zu8w9QYAQxWJVoX7+A3xy8dLQnQ25xyT/IAske0OYsmTQfTV9W/mU
JpPMuXIDQi9NSWWSTkuBCC5G3wGiovR6/3H48IFXfVClJByJQPmKk9ODcQdDRYBC
Kh7ixfqDyYTBlkvJ7VnBdYpzxDGdMBn9RMY0I0Pdjb/qlwhNnO9rGt2vYvJpd15Y
5FsMfjeXUmto6Fj078YEA2TmDtJgyjdKjoAORyvjCH3+CJrI1if0Y3mZaXop/cT3
VQ7MT/g78NZEFN9oQx0Poaok4LpSFxlWFgt5BgfvbnfASj/y9nrFj5tCn6+ToQqZ
jQokWDcuhoyWjJ9/W9z9yL8oLAd7VpmUd0LqE8c6JjitDVfs/qsJSheUrTbDAoPY
M/lw4+Ve+vy6PktIxY57uG+pl02yDTByLbCE1i+9U6akpQ2ejbYcRNHiyGWay/nw
qXEz2DvVBx6yK4YPL+cAJaMDelsJCWGOkIliq0QKRwNdPbVr3pKUktvWHMvEGeWP
hnxknSmnr3sp848WLXcQpppB/EVQN0d1jEBYpceztsp1UiUMxuL1b2MxNJNDjr15
lwAVQXS2Pm7MCDvAm1UsM4vVPp7Nx6L4WsmQMW6BSbGcOPmywZcTRjA0HJ1x62az
nVyFGdn1Nev3pKG0nSK1fe+gfEPg3sFkqMFnoEQTMCPoA7T7teY75oExBbaift3A
aq0hEish47tJuyLsqPxoEaASoMDtKexc+PrgY7HhIwRdQd0DegJQlYGvqj2zPSd/
T9AWt/WIVO+U44X59r6jNSTZ9hlCnkmakvHXNZpS6+S+MdNAC++whmfqQ6F0pBPJ
T/QLyG8A6Yq4GWPUbuhIqSMv9YNOoAblnuFpiAeH3XQPRF+tnS5nswu6dzuHKvLI
vzswLcqUDra1HDwqVstEWNWY6x4UFdVTW0QWz3OXloafhSjlcLB43jahOkxOT8ut
D05DQXcvzHn0PJzAsiSlfSklOyJvImUe7km6MyJRym25FnGeNB7lj0P3UwvMdEsT
VNBnYH83yR4XrDBuWHTtFcGZW4XCvIgfRNN6yqWaiCi+FzThrj0oKja6VJHIzjNg
nbC8pUZdnqdz78Rao+bozbtKqUEG3a+Nycni11ufeGdOZHgqZzhq9ks9pj20joM1
I/sg5COaEQVB/2Xy9PwITg9WKR4lrv3hVnEOXMzA3Sf4BvQQCNPb6iGECERX5oeF
zj+cMpG2ygG21/IFcoVCzs97NABfq6thwAdZIs70ikv/OjjuHLaO2YniNH8L+axX
/aVH+81b7WiTKVzbZfSvoY+TDFoGOOnsDASHpazIEYaJCi7inqgKpuVOLeRdRNhv
OPT/BxeScj2cMbZconIJbbUQbMjgXcTC/pzAbaTiUYIgtxZI7E6qDBcpI4RTovJx
vXbtopEmNJkwX/6esHhQJx3rFjauFF4HxZgqjsxSlk7irfZ5cWQHJwvZ1JDmhv4M
PGuooiOK2+jy7EBGQrb75US9arka0988anGh1vESMbVRdV07vCnqJjP94JMpjLSF
g2aOTNrx4eMXZA1nMJNcgsqwXmcw4ufV3wiz4MwQ45ioofWV1cQWEsfTuUryGe/V
MutNkveNcZAvTIz0RoRpFta+OO79wdMMrtEsrJznnWtYON0nQdxW/ZCzLJFL63VX
afkMzQ5kPN+C+im34xvJaeurj8hupt34KBRkWLRmZHjPvyYh9XiN5iBInXDdytis
i7NfVr4Y/gNqt+NFWC8hKENz5Fk4ByJ8gQMB/FMgziEdP1QPRfMrpj/KxV2V+uzj
DLuFq2rhKlReFlYCdFZfOktzM+PNE0r1XMaAKRwl3AkNRK0ksovMss4ZfkE6/guO
KrMZVQ3DnQaXQH+1gZjxU6+lcKPzt4MM6tz3VEeS2jVEr4pC+DfXcoFM3QSfmCTb
PR2rbhu36NmZBnDzc1hRyEjFZOs1ldRDeazQDpg/f/gJfb3sJeaMTVFX8bFkokns
xBdTHflkg4JB3wMVNoN4VFQPdxePQ9CQ11hhTsvdTgHkOHb0+hCPRza/qKS1tJ7K
1jHetEzKCdA+fzBCQ4g43lr937N/ZonGuvWIwhwYBPFwXS1lL85b9lMnnKTL0s7k
Lo+F4t9bOVD/dlQ/iWEs0p79zsAENe9+QTMHD1Zo/CXzLXMGwzsJ28Mo+xsN4ZFA
x0MtRy8pwiltoMwGfZ4IDcPABvzzs7HZtBClrd8yrsNEPXJX6bs5H8lMjrIWK4KJ
TFfjnSSdGJfMAJemfyi8B0hdN3AzepWDsl0ZluCluJBN+B9O5aqpEuiAM0K2MpJD
snyYf4QBiXtteq4TaMZZUKnFTIIXWVLuzVqdjK/IDZRK8A9lTE0d45hp/tmY8bY+
4OQ8ksNEsx/LWktvsH18Xop0TQKrRb5YmsD/sLaailqQpsCncb7JgeWlHdRY2/Hw
bD3Hj65blgJw+P9csw/mQzsXBMzWFn3Qotp4CAp6dm0udepRX5SORf0xK61gdnnq
XgEUs1/L1YIq0ZTHtvBJTZF+ZFdCpxRpek4Vh+Id604B1N+erUyipEJ33HboVJdw
oijgKazt9IdCduVBG9G6fIRtcblcBCOmT15IhojV1Xd3WHDVuV2Nc4/KZg8XkdMH
MJjo+ryWuIr5oVaFPwNrPTDKNLCeflW6Ay3Bsj6Wv5bGObPxDL784b+cN/wcJTp7
y3WZYqmb96Bu2LO4gKn7381RY45GiBuZkNo/waYigFsJm7JpL4gcBvfLGk2Db+XE
TuMy/9fEsaLodKf1Fe25cOjBAXG4x/MNfUKXeE81FMweY/yz+5VqzP15aAeyb8pR
UnAEGLidq8PoIEMShXWrF1R40A7JIEmNS+YX9y0vuFMWA0S1HETCKNGj9xSAkm+9
Y8+Fqy41VvKUUudJCxs5M4yj4xp8SF3UoUKNyztC0m0UARNf6NJ7/4HzhhUd0yZ+
E+i3HXZaq6i+TOYT7t2w9mvY1ccJNEFlK15I5R/WdhLZm0bBn/jOYDs5T04cExpN
bXiGVw2psvu6KY0NjQHFnMScSs7t5lRR1GSES/VpkjHtvcLhs31k7dgUhP91uctg
Ro9f+26EkiebjJkKNW3aiKmA6PNOFD87q2+Oegi3pI0/e8o8oBUXOFJe8RmFeISc
itOme+pPbNheb807U5GxKFp7rR7L4pCVsRwlPS7FZMZFB4FbbyVo8IPPmEdS849M
8WhsFrHyBMHLghGIc+AzRvyytvVsOVMfQdwwT1JL8YkvyWhlMt5IPLaclFS+NkUb
l9ig+1KlAfv7o0JDAkArpXOgLW7RAj24Uc8DTPFh0+2+N6T2vuruutrcdaOr2QFf
G1VGC6jP1yOD/mDHv3MV3JgYMLUx0aAVnAt92royeUX7KzS1lKWrR4uJKVSSbKkw
gb53lu2vkmsf0gt+ORoDEyYmY88ACCzp/g37WDGNvwo/rnETNk5n2EbFYVvjtplX
UO/gdj7wUVcZN7vWoBuBrGeTwek01rXwVbtj/cH03n1CmIentNwjyVohY+PMvyf7
G0eCxWCx3dVLulp/Qa7H6OsYMY/npK6FhWAHHZauxOibkVIs0ooR7l1xATtpw/MQ
AwrtRCVZrwwTQ71fuyaYgwGXGFvQKt6/mGhZ4Lk3dTQEhhC9ZLBHn3Iz7JMn+Moy
Z17sNQnlxkqlj3aI6DlxieiXD/zyeMsQJDAtAK1XslOVzia0ZpgFOE4lDZwotiPm
CJ8jHnPJlEkNmosy2w5U4YtQUs+BHKUka4AUV1HM6VHmPKaiCD3F2ZDawLhVwc3B
Bsus6IE/OE0VVwAknqtrotH8Y0K/sR2j78smZXd3880uM19FErczIQ09mfs8hp9W
ToqIsQQBdEUwAImXUh6N2Np0ouUZNfFSfmW7rnAvjZ2VAcK+j9AHADhAgptvZrWM
7/+7SKXnm8BUSsSW0ViKUEsx6hEztTvwPa9UxCFqOsGFEd80Gsa+Toyo1QloIS8z
tskveXmH5o/e3hDQznJNrm7VmB21Vt0BxfsIdNyqE1RQhVvpDJ5hDddyKRtp88DL
5UAOIDJCdEcWF2aIIBqC/U8sr5sinyDz1eP6llV3oP0Fg8vRXyKq98D8CBAXEgBF
Im9LnlFPQDY5HdBOlDpVWot2Vdj6kgu9EZ+OmxhNmNaJ1Ti3OP1E5eI58xpCrySa
gImP1NzcEJ32Hj5JynGKRtrnjhBdzcGbpewVxiCqgg6MCDwb12pbskN3Yd/wMx83
7LUbXpXtuDmksodtplxBJVBIv3V5J7QIYrfk3Cld2hu++XgQUhPaZH7pX+Zlq/Cm
Uzl53e4CMDEhKHgWbGiTTHylP0iVivvTrWXgDyu0lNcsjVBc9EHKVaHP/aBJYDXy
BCJjstdZO34exZRmFb8GRDzZ+CuqQfET/tkPwLN26FQP2yV896h+jtr8NuujUv3K
6DHEWRgNNXJ48I7ImSXCI6CwVlAXnnCpa0YjR++QTx0O+Wu2CQMeQ4BwxKmtGwfZ
8A4ahtSgfYcdnlwV89i3PEZu48qjilaB2z78X9brZK9Cu3bxPRPd+x0IB1EXqLCu
a2zOEhIu+jIqnK252oY65Yx9uJzEbVmCa90lIPqiTl0LVV4Pdk2nGYg9DVU/h1g/
lENep2wa5yva+1W7BV8FirZcDchjY5V6IhV9+5r3fX2LyZj5OXEE/RTYM9SmCiVg
eLo9qQSjk4LiWgO8alg3h4vv3Q4GHmGxgJiyZFVEanAx1KtVQga1CfYLO5ZtvB7S
znH+yauCiFLDYENoVk9wWlUoQx9O5KCHVe2aE/C0KprMYToFFlMWASgt2e3ieAzS
XRWTBAkcw99M0f9U3mI9Bz9nayPnCqUCcRdV7Q21sACXz1JykPckk0h1yjue9ZE7
+Vl+qkSjI7qxjKgaicKFpPcwD+YnR3qopOrHfajmSKZTKcHqToR4+/JeBVqhJGfY
uI0uVDL2l8mRsLbO9ak6BC6ArXP+MBszwxlR46ZwP5EJ9udWHsq8FGHLwbwCZT+i
LtIvmCbMLJIv/YDP50nwIIT81Tq3/YB9tEb5kXyAlQ4wzLl7LDucgjdap+AFbw6O
9GMBlsi5Ey8HiZj41JWL21SvggcjfEJqskLg6Qe7Vq5b1ymRR4/BYrM3JOqkIrZl
GPSpLXF1kQC6wlI1WIlaQz1NtWbqMigJm3HTRTdRNx7xElvZKdSInjwKxw3XS7KS
1oCCxzdg/S9SujvwxE7o/sO4oimcLea5XNhNPkZChKrz7NWZsd4DdViEXczj0MtD
itwo0IC25NAu1PJcpN6KQYfaZartyv3tC1ax+0t+yrevq/12LiEUVtcbxcVxuHsJ
KJlvu4H9cFHt7WAlyJeDpJvZnvpu8vgKeCUxKhNY55mRSVKsfsdJoABKf0dz1cdB
G25LKDYZHAY8JNvBYd4AMatHnAMznyd3zOIvsVxLT29TPEGXStyFYcPnuOntsu43
SDF+MPu/5Gr10HnjHGlwFj4GoPOZUFuxz+aloqkmZ2e1+WP+2mcwlunaiA98vuRC
rnMaF30FDMKSUuIAQBVyMMIOY3OHFNbkomihrpO9k/J7X9nCAimTXL937q3Mkg1P
v8g0EId5fASmOZh8YX9MnPyfz2cA3o8BVkRoKA7InThF8IelD4IShjS2CTYY6O26
dHMGzpqPjSk9bOgJGwcLXGttYX9kyZ7ocuizSO0olsL1IvgeLymMoJZaSZivUGhK
RcSpTwyTtRf5rWMwK2kRDPQQ0MAHeUmBjf36nKcmna6zBtWpd2uWLtZm3CZtAuzj
+NFjpm2DPajjN0+bom2yw+uim8NMuksiZ8m85/oHB4ddtp78tVLWXJWVTLaOxOnJ
w2LHS+BYkMpDtu/BXwea5gz+qlEZrDw8Kl0Bq8cTHYaGLvQMFvPk3Q2YLn88s3dZ
PsyHvJsu2QOPbzW1h4MzF5tP++8+Bi6eFU16I17rG27X6V58SVe68PrKWTTLctH9
TXd0gUG/bSaZwIa48jl3GjUIGcaK7R0YSlb60FIiq97p3UtKLhjghaHYe/qWYbg5
eCprO1jbqhiDTLN/2Vlpaur7LTGic4WI9V43m541Kz+m/Bxjoc8/hFKwMywJX5/U
XIdHN+F3B25OPX4lfQ1HmcbUQ3Pda++nZe3zj6dTZtEhA/GIhSUZwegavKVexF1O
l2uCBNaFL42T+jq0QiGhb09KPDOJIUYSjulWN9vUQN+qGW1LCdQcBOajtYCac1bd
G6gQpPJm3z2+O+F5Kb0WAmD7hIQ4LdcbjHYixlTMUrwUBQm0Wp3+AhWcSlOIakNp
C/zskL3eZJmn4F9RbziFIsf+ieS1YCkIF0O4/4lKMUD5MB8PDiDWaF8MYmAhEq0w
7SSbskC4RIjeQOAuGxqEhOhdeiqBeT9hc4hbEXJ1SV5Go45z9bYiy8f0127P6Rse
xBforo1SqrfjMAR6rniITREuYONCNjVQ4ZgpG+J820st4KfsqTKwnnrVPuF+dKUF
TpSjT3L2y+mzGpqHSQAT888OkQFbaozcdvGGmfb2A9UOGzqHKioyOIMrUrmvJXGN
ZBcxn21u3LU1hfSSYUQ3wSQHsnx3zQU9fEiP2cZmH8a9aGrNalat56kq/jWHAujF
RGpOFzwssot7In9+UPJaOaXfoUNb47VxWCeCEQf70zbiLjTcbldmHQr3sCPTNwRc
nF8mH/cj3eftrsbLaeCTdI+eg53yr4g0zXGom26qC6v//6nqcC/h2xYc/7l8u4/v
xiVGCFc6AL9MKYt42mxLL2M0tPJaOm7oBXA83cEhTbwaLSMuhhx2HO4FywlYi2h1
aFFOYUYKKQ5I5ataYwPZm3ftp4t++i/T2E3ZqfM5yTU0C4zbltZKq9aNLK9WVem9
iopWvItKWetNTSTLJvgIGlm4eOmthVCZcFGWw6wzndP0JYGFBaBaFa1YElCjz6q/
W6xwP/6AHp3GzGJGlxRiilydqShrjEYPNhwf4YqPofk5Du6VJHUQ2JKwWW640747
91+lwQdpoeaLqJONp2F/HHme+Y0izaooJ2JiqoyMEJDUxjIxVqDddMqDbGVja0SQ
MzhS+jXawD5doo5ObkOAuRjel/dJuigHRYI7+DbOWcw+5cjYlDT4zV5d5G5kTLmG
sSkjFg/Dz2yQFtW6O5LJ6s4qRn+KR3/D8m76yWEQc2Vn05IZWRD4c+tyTJNJyFzf
kVr8yUxm+2JcYHOZjm2i56dolEPmmlNzsXh7ygncJNuLaqdQtVuEurYHPlD+S34u
6fNBeYmwd3y6JNJ3D2HTmXCf04y2q1EThKq/yAI4NxgBUnutctkhHmWeLpZz14kE
kGaCW85DnmIH5+grveQWeTn6X+gwzibzLecW/6w3AZ3ghAmWwy5b0t0SJyiN9GTi
mFiO8ASWgxRp0mvST7qynVj68k8rCmzVkSvPj1dgMJXXQgw8iqAxMiDnbRuy2w1Y
mu9B5pIuoakDdMmpkT2emAagh1Se4GxJfvOYwqtaQFugehpI2IwPdkANGABciZRM
RkG9z9QxVI1tdQb6bvjJNw0cTjWkPPRMzCpTbAsrFzGAeaf+t+776B1QYa7JRHEf
h7viLDbo5fxCHnfD/AzzgXIlSghUpu7kUH/0dpe8Ro6eEL3jz7765e2y5aHyjb0k
dbgaAXPLIn7JJTm9Ge3pmIklVRt8qJhhCxfbfDq2ydXVM87AsTevJ0IXYOWQSvvz
XFaAwSTcwJqQ7RUaNmbQTEEr+eFaO+I3J0tk9AGhhWaXgqup8sm4Aq7d6fQOdVQb
rA+25Vic8iHvm1Ln62jBsyMpq3jB2p9bMkh6KOquQ0z6KfX9cQ5jpgakyVQXkKis
nP8K/8oGnoOcP56EtvdJgtwhTuo0MvLPMYqDIwxswHOZ6v8PfcRvirWzWNm/cBB4
OuroioDUp6/g0At1+AtnNVfsMLK8YCWkj3DsR4+fI1GlkYAprW3EpTSWBFwfd9mz
xXBw8aqwfmwrKDtamz4884jWDcr1JvoNF+LqY0XKmoW1JlZrGNGKUriLO9nRBJ6Z
0O7Yfc3yaoKutKp8/vzzOZzFsBTKbRKbg61HXIm1C6qMbjO5uBIKnCCjwNCqWGtV
RLXFGlbM0baWnaZe4oxptN+U/ppayS8BxliUJI4Bru3VNIYaHAkOuSsEhbalUfj3
PBSW9Zm2CrzHpAjXQm+QjnoZBkI56ZUEKqpZ6KByOo61hRcybKkpbHwNGNYXwPCa
U30+vFZ57Td/OQFQSoaifzQMzl0c5Ps6y11Rc2ZPWAiHg49OCF+ZreplAEdsAQJ/
kuFE5zzB3/TwhqAcf/LoghiuysVPwxg8G0tUiewKdLJeEPucnHIkw2X1lgOsFG9/
kFnxUGyurHRANrCfKCyduhoizqVn/bcJCbn0B6uUf32iCr9Tf3KQ1Sy0V5AlSDgm
4cb8uv4XGh5EZqlow25flltKscB3/Ds4k+sc7vcsdisdicEaf1FAbkBfPSSLmM3v
VsoLbOmFUggUrZfw/QqhafMgkfAFzHBDlDtuWS6uqL+in3ZqZgTdiNQG9Frr92oW
wjXRxfVwxY+44Lm4A4vx5Vn0tb4Ltbj4avU84w6GDShjeGQURtRt83DzsmKgyY2f
vYG0oJ60rSbbCI+/idTK1SiG3E3V8OX2BD+cmUAkA/OCP8TViV5e78PHtsf2vr5H
MAMRxL3FuwohPoKsd9JyaP5yQBv0fZO/yxHIcd/2hqHonh25Bhsp9Ti9RYvDyHrn
GyHDndTSGnFubuF0A7X3PdDY63DdSEQkHzpdWn1y0ui+xwLMH2Dk9JslR69bpgpK
FKDiDeViKv6+NiYMKRcCrzPgLlpuDG4nRgwgr06l9oXpuvAL2rjsjBaEHIR+8IgS
RWJnlMk295911DJr+KzsLSYtz6nXiaDiwZ7UpaIONDfKz84bSmozYJGsFMVyaECl
r17Uq8y7b7DPtps32n42bI5r4DBvAS1Xkche10QAmwS6jCiuTjT0rVI6vzbHJatd
wsv5LSC+cUeQyWg05W9jwpCC7A0FnXH85JrBo3rfUjkIxKPJoG3Q+dbwD+2YBx51
E3YZROlP0dvnUz4gOhXAGU1GdEOJUOEpwZtv14AM3O1tcowwLd1EGpL2JF441Az3
NJBeWusGl7s9CloWjCAYbIA530DDdXGd2rX5+kgEAxBIUV6MCgGYOW5Pr8FZq5AY
d6dj5KpL26d56TW20/7n/cB+TqhRNQo1eBxW0as9lWMJQjHlFeVObRNJhqBBnfTs
REg8dIQbYjqI9IXqb2FjaYqulM96uoW0Hz4G5rCRh0UoiPn57+z243uQVzleDSpf
XGIaP273U84t+lBULKBWemOFOcWD3RiFJrfH9TGjmE2p69rdM3vTefr7+oowi5gy
hO+ZBqKmg50hsQDdjD9XSyVJiOEowUif5sZekp2DLt6t0Y/KFFmS6M2PU2GJDltG
jco7VdoKty2g4Rn5DAJB1x6XqHst3+eSSYwxBtPXIltbYViNAREcqYXtZzaOymtF
NBR2g8vhUQnHoC2ER5iKibjzE+e3znobOca/HYzn9fUQcqwVCEbp3WI14vI5+sPT
ehxd3MOBflVreMOhbAl1G5nVIqbK9XAEyRSiiyisGxgW9AoV/IObjSY0lIIvI24z
L0Q84VfHmtbOx1grStRXgVXDGLmBCc7VR1AFxH93SRl+nuT0MUgn9b2WYGM1dT4b
hAj9C6EbkL8yqQe3uDW19USfePWS+6S9SlNiL1XRIeVfd30sMwxXtMPpCAeRKNcy
m536AdgG1/NECXpHqDcj/LAUsER3uHQSr4oUSYATKHXdfuHjl3og/ccFUN/gvOG9
kSbr6u3YS41mgq7V0F2b4N9Moouhrom+fCJXBDH9ocjFnt6pI0t0mwMHn4EjQcCS
d9AVFWpA/HF8ZKI5KO1STPCBWO1x+1LGchdcfLmye2pShULendSOctJ83IZfgIys
Ibdm9Lk1HqT9osHQE1kDcrwvaPvrZdCrVWtN5cr4gyD/FhpLV2prRvsjbjSUGHvY
4Fzmt+QydrlVvhT+nnav+RtA+yZ50mRve2FEkHPbUbEsoB2s0s6jQHAa6J30ueFY
lK7M6+tCDMs4d7QwJRiKuJFWAW7ClTllR1swv/qjdf0p2AvULQCtEqKpo+0M5WJU
8sV5Odw5NaRBGi7612wdvpTGSDjcPIMR2CU4Qn/g+0nq1RsGQBHuMfRo4WVgU6zZ
hvbgw45BV4RuE/QjfE0NFxIvPaqdvFcJOFxNhli7oEVBZ5zGq6RPbgM9LSDVvoHU
/Ll5cwtetZFmq3x3afahHYZYyafkfxlOcwh9GUcU8eMYGxTMYUtkoYF+kf+o3CXQ
WrtytgLhGlt9TW2O0RPoGaO/oHStJB8QPQYChTMKQAN3msdPh4ivOXU0FkYTfb+m
G2wvAwfG3psKAyccpzq4oeKgg3bU80ZMhsBS8Psv8xYJdwZ/0suD6K6Iig9YYUO7
QykY0b8X5oEZU6QxrV4xuOWxDat2FLeu0InmMQVwW4RQ772Le4NPlaHohk2kM56Z
plye3aPNZnUudVGwAO+iWW2Xzd9er79NHxzevfFJixcba8++0tUOVAMiJdjR3FXk
CtitC+/djWbX3mf3SiGh1lRn38nFsZLW7vXQ5O0kubq67lYv1PUjJMyBbXh5et8g
mwgLypZlqo7NSQtAiSLFC327v1HSdXVggyFRcaOQh+5Vug+fXtQZkMhw4hdEwOX2
34JzKyMqK8bpuZJ6VjTZpMhP/BMGz4RAPYX8x5C4vAl+fDzpqp/PCU4EjbpNoohb
+HCxCOV0c+Um7TDDOGexCP+is6gsJ3+N1LDGJ25VpxuL/+B6HwK/0cXUXxHds5l1
WtOueZyFsRaZPMsto3gBirbrRxfvr8ADJSkvd0KQVHfq8GLxycEGPH6CRTythyFX
sXs9af9wlUa7LbkNYmNuvkLNECI+yrjx7GYgA7RJ8SgDtgQ9A+E9VyN4txf6lpnX
SjhGb1CvWlz7VkEAe0H4CalSumDzRTMyoGQpDHF4sst4mMK9awzSWiRLLry9uQvH
MIFcMekuSFu8LrkArC/OB4Rzk8KCrBxCpxDz6CllnVBNrNsli3VaGbrh/msh3sqt
7BpertmAAMpGAaUITwVNqnCQD9/7kFAoe3nvGNBwgvZ3bUxESum4LOaRpkEY7SLb
NDTPCS85MOGleqvPfRS8IDvQpAkLBxhXSkNBtxJMh1HL7EQ4M8tHHYbSNkyze5zw
DjmWyh8MJk2IAFM4zXH8Fyg1nv39wFoqxDJCStbjEcyRtUJkNCo1qz1T5ZEB9dY/
Yjw+aC7mpzgNI8Q/HO24PZHKVjxD6D28/N23aXKfwN0HPODlbSafiPFOKhW8hHXL
H1z4qA0WvmawfEA1us9EbInlrbv7rPnmu4EflXR7lTPj3+URO5dzjZUviNH2L/7R
57OVSCxkQvQlQBXft60LOmVJq5ek5oJcfyMrIBHpUaBI+z8OMppiVX6U+0WXgqHB
cjNzaYleQ2FS6O/9tYg39EvIhi+mhsTSE3sHJLBa+ChNhaZ8qFJoYo07azQ7q1a+
UHdYRXppoWYfefWUkG5p5tGFpUEs+laytCz+KB/QTRXKXVKbLYdotEg3Zee+wBQ/
WG1oDBCsNm8ed7Qdw9CfTiZ9kgq/yZY0S6cPFt8baFLXFgPGMdSgZk1G0YdA8cTQ
XSDhdvDBu5RY7Gnp3I/wMOEifo2nkr7ILdEjFu6HwotAtvjvydy8iACS3n4YbG+r
5ApbVLUmT0cxk0L2EpcVVpN2mga6+Q72yAcV8mmaK4358F0BZgsvkfSggRq8mXov
zkapJxf35d0JfsRxJ8CBfQYRAdFUuD9jMz0+ZqWG4s2gnkixH3XSH3E8w7/JBsJ7
2r7NCHIylvfHyCh56a6kYmfikHkBeRXcEedQNosthWMGMCR4OOpV42MZBbdy/YM/
w+D/GX0xcZhKTwo9bg68gHD+f9Km71yb3mSfHno6plkN2xsr5P1wv4UnSoggLUM3
y7PceU7vEt0Mgtgk0+p+hdxSJXzU6Fq2Z6HumXw9dYpHnFb+K9FppmyOyrREnwdI
6A2f5aD45jhBK1XV0L1nmfn4TkPVHQn94dA+ySIKKL6Z8q10yhsKGk6x5DPg0bhh
fgMQbhxA3XYuJCPWrvJ5NCQ2gysAHJQ05EPKzNbmR0XjDYpr/Y1YVz2dJ7icDmQF
deknU0ySxKyU1Cbj4LJUjv2CfMUotaSXqbFEDyi/2b6NHSUzD9LiVfqQfeBlEIuT
McjFjBG2N+Dz7VvW5kBDBJQEgi9Mrvu3qtGVa4RWMGlwZ5BqYBm/uL9zaLXqyk51
X3oi3FDj2zjcPhuHsTKRPXTpz0UCXkAkdaHb33jtah4Pbsm7aml6otTtEJ8BPNRH
rnePnR6bPW3pE/I1IIvPH0bwfbcd33k/5Uc8pnIF+v5lfScvmm3DSLUp5nlStj6U
Z0kSDESsDoA1C6ZmpyggHmoWkzoaJwRgWaf4/nmyc/qxPy5aB+9UVkGv3D2HLhs8
hcs3RE82qfjKumRikQeWERcZqHJXvTEkN8K4ffVyNjZEbq+AuQ8DvV0RqbqFuS0X
cbZ3GAaTE51AMxgXSYeUFzs9LeBcpQipF950QGF0wbqfZmPscNr2XEwARtwZCrWr
LUm3XP8/zqvwdiBulaVrA9E50uunxGqKBn1Fbz/ICnoGI/tSAQw2M5QSadRme06M
ovmrcPMxLoOPx2KTXAYeBq6gtQjJKv38DvZp0hzK7C6GTmo6LeuVeMxuGS1iZdOy
fF/QZLZdzOr1Z/16jcTVXnOGKpne//IUddvGbkXYyIdT5b6E/8zG/j19+ZksvQ3r
WCxV6j4qOWMAgR9wZ3PLd8UbfI/sXClGDleKBVdBfXLJWtoML/48nCACSEeUlgEO
tiSg6xmXE6tt3zxHjOaXndc0nMH+ZsSec8QNgki4WAk45pMEw4nHx4i4Dmhn0QkC
zUnORyqWyj+5TnyM073YXfWKVdplKkzJennMOyPObjvE0JaWy0+4nW9CADDY+0ej
8IpfcE0R9pWllQVVbSexqYZ6xr+aZzuLyrIvA8TTmf5wWKQGMJ3FLEUpxGijAChy
WOKGuSehUZi9ODpwdoEKG4ZBtqJ0xBqe0pVarQlzGjeqIX/Ondqw9XDeuyKsmccC
NuNXuQGMYHDViQ69l+tAbnaE5PJkTsRmfm/kpLcL4Ecsn2Nk0m2eldHu919GE96F
bCy2frkBXGUCoOSTwHyN+tlSuXB/awAXJKnIwq5f5hheuuqHqNArUZo9tUau/jBi
1TbM0xw8Ml13QQTfpo6Bnsw/9ZNlJ9/Qsh/SBeK7lxTjTVA2A5nprnbnQk81U8EG
afJZf6wOZaHkVULchaGSF660Wl+pBv7qMwjIE4HRMUsrdAH/zRkGkpSJflrgj1LE
eU5R06Q3LRFL8b3CpZRsEsIHuYc734HWoFZloPWZNJJxeyhHwwm1C0rjWz/fbxtk
8Kf5TXpOXJkVUV54qWqlWNx3qC6gmaLUxwkmHCyxrDXuAX3T//tj9Od+y+OGooap
TsyuQmezBjExde+f5PDkoa50/cE4tRWaS1R3rBSSk6kMmSCc6kBmrbMRDtFo9HLs
qCITXnf5T01kEDpAcTYrcC10mDkLCKaxDgOfuEn7JKQqXS+65aaW+3jefxpa5083
/Z0k+XMCeHvjE349dmrFQZfBSDRq/l/QSfqaTfJtsBE2FERi8Sm0c3/oXwH6aHYJ
n54MaaYV6xePRx3POak3H+Subxn+tlCDcuV3lX+e5hsolRsO8v1HUDEPQYXrVoQl
u6XsFE0EOyCL1yWU9l+E5bsSR53/kCSC7+74NMmWMadLzy7Pv7i8/LMVLsw34Rca
R79kawyowmZ4h1XzG9D5AaiQvyrKSq9GVceLZvWYlnDcGqbVKFU+HKAAEAQLDou1
ILwd63SlKfBMl2kYWhSn8anFIvnwUywtjpp1A3gg10LpiaILeyu6heZmjdG1sWG0
MLX9dEyD7HmIvjU4/jpPJbVrlJuZWoM2cjealng7UfPYYYOwQQ8o8GvfsoZEZsy6
sESePJ/CbP9UbB9YTlJSfwPEqNP4PVAUogBobaimClRuCuJGoSWmaS82eCwFGLOR
mOBdLKSmU7B+zr6OVNHyHwrigOVWeP77WiXA4Ypn8Sen2GOcsYt0ATnnZ14e5o6A
OaVoho33kL9JSD/l61W6QDw2lg9qQ90qTjXw1GeES1JQWaVXpCenxC9CBQhL3Y+H
tLEc6e4uyuu2DQtpxaHgIezTcNhSMvP6f84uJMQghncyPlAmYChg5RY6kejit+LR
f4FH9eKqQCb99LL3gT4isD6ZlhVV7bXxFLWSf5ab5/furCNkbKNxbQvWAuf1plhh
nR29gmVevXIZW1eSpnmXug6Jwbby/G4n5qltcK56PH7Prph9b1OZLpArqwuvz6jv
ZLwdTK+EyYj2a6LjDw0C8Y7N+/k9pZGCjV2GyMTwG65vfGwWKkI2BzTtENYkt3gO
g/lqUhAFRIPs1RDyHG2gsT2OwSlKFClGPNjXRYiOom0ESpaHM3//YsBMMfGsIEXl
bX5k4hbBR8Fvx5FZpkXb4crNfU6PMauj//ztnBhnmaLNpM9aRP57uZD1yAc/8FSW
G6W4qgNTbrk96Mz/aE0L2czkvNEY70L16ouXJJuuzTScQmpoTlDtRjF5mCk3UEdu
hA4VelkYxJjgfY/OgGaXlfqjqRb3ZiROuUEdzaXUi/yvDBYXYNcR5HWxxJsFtT/K
Kgr+X+Sb0cnuJkTYX75jC/DVVfbMu20rzSi50th0GRYNuoK6RUd2rY7RmreuegeF
rm9/Gr/z0z6mR0ouzKiNJ+EUePFe20c+7VrZYGmyzta82VX2sxDiJ5VBV9sx0tbo
qj0YgzYPYT9BYl14aXQshZdpqaL/IqE/BikXnASQSKusm5jWhEFIoVe3Hwn0kYo1
r8U9hb4qrm9yvzqjEDLcD9AhYK1dLcR70MW/7t8Ve+hX+yAvi+LEa9y32nyXY5OY
1RGj83AOW5Scb18TDo58JKWu9CD3suy7SYdtyHGyIJ6JPlOi01i6G4/iXA4PoV6I
2KyUFoNyw0unFGxWlKoikwG1ZtJwZhsDBpygv0x1I5pwE9SxDYVFQvuobvpXet2Q
dqDbuXW8Hj6Oyp0/pzTarnxLANzKuGK+XV5DMKktXyNAo2bj+z3ZETtsIH7st3j5
T16EBcoN530WND0oQ4Pq7AKS65PUNB6OYahR1GInRfARiOgiXLn7U7nU1IdMLND8
rd5MT0HTCKKTlWK8zSYO6lh2dIJjB2I0wfPgHMceuCnjgcgyr/CrFd0rWQhmKu1o
WBXx8l2tiLN0AK7Ny4JLaElsUHEbUhCmnleoTL19+mGhCxhxTLY1/W5bTlbE0wER
QyIcp0GfcYzNsW/+XFDhutQ2o5I/W+SaAdrE9tlwXV+ZIVmAvIKuiyFq1h/5xOvz
AoxR4UKwW4FTLGE6woVuzNavs7tVSmHEk1drQkOcAFsrVM09/k2ZJgXhXfPytEUc
nznvyLS7QFkYe1VwZOMZRVPdtX3DFk4dk4YeGGl0oChTOff/Wllzp5Ibd1VMRdAY
Oh6vz7Z6K5fuS9KCqw43ZDZTdg5j8LOg0RdadH5LLoKRD9sse1zKOLXVKo610giB
nQs6XRuG/+/nmxtMCEyKOj2n+IIbkSYSQYF7LzBfld/9R8FSbQfLHr4PO0yqFLDY
4FvQyLdvnSaPjWdFF2bh+zVMUvu2KQ5okhqy+baWzmrf8GLvvhA+Y8Ee0+SHtGbC
6PRaFWMNY12B9XxLmNfff8txVy8aYLfkSzayvuG6afTzM/bfTIMI2xgUGpBx5Yit
30ic1n6kKbiqcdEQnxFhwTsZSZ5czXt33IOomKdgHHT5CKNybdMAN70U7gj8ClOs
aAQaHAJx27e1lMdY6tAvXA3n/RfC2TjvoMqvr36V2yVc82aei3oSv6+ujTTf8XFw
1QesWh2fykA50wsleAm6TuQIWdsO0XOsVXWaF7DlyX0rHovtZK4k2kEW/6sD2lzX
3j2nGMtlReLqkdd7Xl44Re9/r+KetDWi39WCFJLQTtIMyqcRENzNGziRrWwbkpkx
o+gCNWfawQMo8bj3Ms7PtwMp5WhU8CoCusmwPXMVAF6yE2P8WKGoqlHBw5oSef17
SJzyuGOkv+ijx/WTy30LXIV3zxZeQfUVcHk8xM3ezo80UTQ0pvYxpMEbjyYSUUR/
q+r66bLFEPK0xd/A6TYrIJf0l40YyOTWk8YCPK9A+a6LFciO1najtfqgf51QxKgJ
GEDRUV603X+gOqXIF1hpYoneYhf3Y+IFo/y0C5k2bRogNero+LuS4S5tOhT+OZX5
wdfIAta5YuqWH8zNAjPFFo8+/u076S0JGsRjEWg3T13f1TftT+SIuBkSbRoNy+Lp
xooAaBahCHzv0aAEowz6UC5EeKG0CwfJzVsoWNSsTmXCPW9oIvFA96yLkvjQZpZx
W0vQOcv0KEs9um4Gonmu4IEKippN0GWInC1ScejjmeKo/mzIZ0XwDM0MEiAsWLT2
99Zcbcl+2MxH/TIOPwDKtOKMSxDEpdHE8bgg8pWwb48z+k8Vi8/2EWVyiS05XoGM
MDtIz4YF2FV9QGu+2/tUR1NygQqCya5k5rZV9fd/mHGmEMDMZVagSB2Hl7D6/Brz
h9Z91AJGj+707mfb677T53tWU6elTKmBDQfatEeq+c/sLx8oRgRRiFmj0F/IDc1R
p5kxjs8rQ7dMBxATxqmWmKtYZmP3qecVX8m1j5mPljfv5tBPIR9+q2kL1c6YHrn4
jgP50yucx6pSRZU0z8oal5lD7h3kwZcdwhvGNwrczTF+kqCRKqu9ppa74jbyaNpW
/lLhsNP3TMaz2vmzmOhYnKbTQMbYXe5C71jvlVxAdyTiBjpAIo8PaLTwpW6IXmxO
q7ZZXFd/osRdci79m02dOJjedU7Jt/gukHjLGok+1ll8VmH0P4CBU69VpKqzV+IJ
rOXVvTMXM0dyPWbyg2kEs9psttBdgPXrejM+fDKaZIAOSfFqgs+Vwo6a3ZNx+Pvc
S3nYiTv+BYlxsq1L17kfIOpuCmHJOX8bduHDbtZvQoA2X4nWBbNyLJ9S/lNwZeJa
UKGI9ttjYTHwT9Ck/QFgMemnrel5t9kmV6aNF4iffQiDFAwDao5KhDUST4CJNgOg
AgLsjGaVJnXk7rFIEu1kw0je/XNGiHTk8WFqrBzBtgJounUvX6D17N8160POhHRq
rlk36392aI7ZAmJb0WqZiYUBbEZbn6JnKiwBb68qeWN/VMW8Gt5ZmO56+d6M7t+B
zgTwfvYIxksFzShUN/59hczrOS/QY5ub9GDi7tAt/Gn1gxz92wxjQyMjSZ0c6luG
oB2qRlZ5wxo1g8VuRrnICSq87Q66E1JyQWVj7kObX2ZlJUgZEs2H9NKeC94xEtGY
zhKMNqlLJ49ZiEefd0DJ/zebnaUF2tWOEREh4s5UkyBEvQ5izFykOOao4PX/wVoa
tpgJwp6KXnK/CJP8dGAfCg4VyPtrEU5Lo3kb1ug5UH05PRm7uOR3UUVLNAN7vsXz
venI/iGKn5ErVwu7M3SxNP1Dui/7iBfc2NIUjppF3enHPbbpJIBeP60BqePSAGSx
K6jh5c76b17BxSKAtCcVYZybCzdWTQzmGS/n+bCyHCayhh9eJCwULgjrorzY4/i0
bihnVnJIKX3b9awsf3ehDSTFOisYn4oOS7/KOf0lGqdHgqc80H6jT8+X/ldv3XUF
zaabRIfen5rEGPCuCQT/1m0o3PXKdqw9caSByAPtGb1kv1U1HzoUt2wpz4vxYBL+
IjdjHSFY4nA7P+piXxK8cV77H1aYyNAfG8qdqCJRKkkF2TUpLXIBibhhQS9G1+MX
6aPfiURO/b+CUDM2zu1IHlK+ackr1B+Eey8auy3DHqLN31neTtDtRKF7pcg+NB+i
Qv8kKa5mov8m/PUrh0NYpBLEVyQIMlzMuMhySpl7D9VoUn9Q0uC5VbvR7xxe+sxS
1iwgKBUgoh0CujfVURwwBLmOPH0fMj3gbuYrhZUOV7HqbZp8T8q0DYNyRLj4vRKm
7qDqPfO53f6/CFmTZC1BLDAk1Bhtoq1eE2jC69zu+baNgHq2/a8OFkrhmD/mbbxt
kjcxkw6EDJ+943Qz/+AgnoQlLT/vfYS7wHCz1n/b8LMB3pFx0bBB90hg6i4TGkJ2
8k/du0EkuPOyROBMHBjFsNvXqoN34tvSyHFhdBEyBstuveh+8sfNkRUXiibq6Z46
IwiJKptLE2ohDZqjEv8UtNrB6Q0iYnRb1SD62R8BtDD9o0M20mNSmQP5vi4PFodR
UszwSaQHcaklIAOMDMegOSlCwE8vxyF9GkZa93nspxpr78WGfNBLPme8KUVQuUXM
o8msqvEx1xLIIu5JLQtfGoikqvsTTXrO2DmhignPzFtVpkrxvq5HPhZhTxvw0n8u
8ZoqIs6l7XMXGSgn3HmlRBzwQztWmIIzE3vw/x4Vl6LT7UJsd4YVFZeeP/H+x48c
rrxuPn8/COacECQUjdIfDP0SxWhlb5x6vW+GG3/nuSMacEXI/hjjS7sLm0n1Q4u6
xu/+hbW0mfpR7akMz0bn2v1IpQSSg3SzBOeXrMXh5L0Uwvzvpo/E/6H2mtXYy60P
xjIbR7rn3N3mwTCYqrgXVnmNhHPw/lJGc5mTMwynxEE5NkPxUf07pPWxKY4LpHY+
UyVWi8Hi9I12OlyhY19QUGOTlaZ+LGBQa2GBVS5L2SH9CILrV/tELNWblR6IhhYB
VLMjGySjxs41qE8EHzdV3ztf3DdwDk84+OpB8qo5DISccNBExSoQimMWE/NXAEd+
5bZMJyfoMrPUrqDYbE2weW9659Xlsed8oblvuwqyX6KTlDXFoTaKlJoedwBR0JV9
UaX7RqBh4uPSYqOQA7lTbl70LQUrYw0XU1h2LR8ij437vTAzu227DudJZx+rWAmU
D6o93mL6CxyeTBs06tEyXZApjiHDAjQ9razyQie91OOB6JRjoZeS7Y1+sfZEwBis
0sHS4IFYhnhxwo0mKOJELy/lLjdSYpRgvXAECpL3hyf+7jazC8VJVsJguri8YBXP
+5gISUkP8u3VkEWEbaCttXj1WVQNduJT16dD3OON6JhEySRmVa/sq5IMmzxew66n
0Ej5ReBTF/UIafoqc4Cz6Wps2Kp1r0xn/3n+UYbwwD8olUY5IKKgrdoYpHS/r+xp
sCu+izw1K8DEoUsdBZUvjFxKVaoiwrsFoid+tOab7if/cFG77ZFiL+OXuUkBQuV1
JNPw3J9ef0hktIdaWELPLmKM0H5q5P+mF8GzaHW3Z1ls8upOFjoHG2oBdYr2sY1s
uBmVZUXIFP8VWDbg5g6nQDI+ekKiuzWkRjC+IabCHYKDl9yeZxUqwNqEOw2WkUhF
LIbkMMrU8SwEb6B7Oi6Db2hO5Sd8uCxCT+X+fPK+KTaOL+KfwhRXe2khmYSo2bOP
slaacXd5T7uKveNPNrGUnUmp6F/nlR6RfzAkVS46HtlEB7I8CAAAf0gsc/xzrvzG
diZM9XXUC/w0hDrLYPnvSDQoLn/XI+AikUgh2KAdk2STi8zaPOhd4ayLYV7jmsix
DKr6ZrBgPatp3302trSR8KddWodtvPddZqoQsv25iATU6VOJ+t19o1sGOuaqZNHp
ntkRtY2SRBeERE1i9RCER94zreov+HRmj9/QmYgrL+FoxKhTY5c1F9KsuZM2RjDY
Rk88/4zRxSlGFtKAzg89w/lZ5deKYRvFWlm3GeyBPacy+dpChwjIfe8YB5ZyaA79
gAQ8fGSibY2N/Kdhzn93qi49XEcnHMw/baKOehM1aMe+0WNigupFGAGErOYlS6BJ
EF1uLDM3RQMnn0G18GbKvzr/9GLVOCE6Fr0pzmxmv/9GVZKoor+M2DWqxeg3tD0l
/tQmSqfL/jYbyMPuNo2a1AtRc2uVEwSFMmJnh/LG57n3YM2mlYdut1pcGswOTtdy
qtB0GioIhf2G+oKLVpP29AnLNZr7rJlKWnl0BaVbOoFx4Zuul/B/5Ib6JaVY5+FZ
vwuRzztViIwZLFzH2fmyKRSnYR2Q/VNfrcqrYpHya+VThlPQrcwVnPc8QYZvuAXM
3eJfIsIzZvFfbhfLz7FL7nIdm2Z3H3SWRZlUWVeG1rdgSpbBvgC5KtOaVIFdCT/2
LQd1fN8wOril/53i/rxDoYU51HUhxvNbUEjt8UtN1Ow863WVWrYHo+hVI+2GBtFp
4zHBRXWya0GRKq4GTpuaFrr24hbh1oGMmhTK56hrL/9jJNSe3ce6fXCkJcjnHy1J
8cbp0E12tbsx0zeTn8DG7Kwus9xZDgebtVu5gVJrtxZ3hwaDnIcagYiJxywXHZvl
sgor4rsXtEsU0BiNm4l10Wtjvj2UP29N3/RrzFap8Tjd2StAcccNSrc26OI9L/tg
gy4su0dFedaD50y/AnpWfqP8VHbRVWG/IB/FbUBqA/YX3JkHi3BDSYi9iWLXtf3/
B0lEkP8bag9pKDtVcVsVARJhFhUVuIG/vMnGJGlt9gr2VaPCzM/mi0wsK6naDUPw
ujJDdckNFc3xWqiZRltAVWsYIszA/0QIgMV3qzhqezO/IGUUKc2/RX/78OJT7WOl
hh8rZ1II1alxjaFWx9CjRxhHATEEabrTwkmo1VJr8noa8Bex3EodNS3735Jd/yPU
FLwygHgpolYGIugRvdfFZplf7LVjQN7D/9SyFabeXYx9PoE3RU3a18z5asR9dpy/
GBZF+O2EOXnYyEaOz4kW+Wl1KMlvAZO7ctI/H5yFPoxmZfd1oxztoGo6Y2LKW1ob
m+82ilVMce+9eI3+3GOCNpoALoIbS8Ruu+uyMpPXabBdWM8MmH1rK8v58g8FQ7ZO
G+J6GL08VQXFxYoJesfRJkWYJgmaZWRTSKWOouxGBuhDUYm55heWD4ez/H9GFpFa
VSPEin2pnfdKn/V0tz9t9LNzJLzV4+/hngBdGDAV4dzreHMdeahFrr1gmrnPGf5U
C69pmW9nWgO0SvgyP7ISbWWCC9jyYhgFphKHjAdxk0SWUXED4QDOz2D5TOMl39hA
X9GhCyj2ftDOWp7DaGf4qPtq5WuL/O2pG3lm8/I/puVX/00158UbaFldiEbxOY1n
MLMRGW2rIy+wxPc1UKJZ5nHFR7FEMZTT6/pODmsf2TCH7BE6zZKNZFVibHYiiwwf
Qq8kaqZzrkxx3STOONljJ3L4FBjROjbXJBgEPswVGrgBFNG5Jswc5iujWySgQNhF
b5j21ijrbyR+bC1bq/gewkRwjM8deGHdaMYNDQBB7makE/ZtkWgafMGXWBBPuGXA
xA9cHbUgHk5nUnqvlxzHykTZr59AREYnPssxuaYZ+hmCanwZ2cQZFvicIvnA4CvX
bQzyUiUwL25HO48qWwlvROK8PHoPIWCBEjJFOWzgqPM2KfLHH0dRx2JeH6hHHHpi
B5+F/7Q4H6BHQ83QysPp1gGO1ZDKuCI/eyfo4Q6ztVc1PoHiIOoQq0iMA52eeBMe
+enRQU+367CCsDp9mMPBzm2vs8XXc8RrokOBudin4Cmo4yvedRe3DiCxlugkO3KJ
0YAgnHawJUoXlYrsJhqMfaD3+kT5bJ1TglyTkjpiRhZFHXCi0nqksvUT/cyI2tp9
WxAB3fwZalrLOALPv6OsnIE+3Ts5D/u615dt0MhMPGFfnAs0yAoqZnLJdwwvjdZI
iQpCiJqS5RaNUj8RKBEB1VYp1vLxqV1ox95SODNUMR8SXf32xgwY3XR9HH6pMtnW
tFPPKpMKsd9R1kLqCnfPMHDlAziv+Y2Iy827MCz8NL2accCDCoeda6HWcEZVaUnj
OVqYtHmDenYIaOTGisfX4yq8lFqRCQAQ2Jj2TgeAQ/3/dLW91s8xWhMOzcQT+Lfx
Wi1lKx0UrjdUFm/r1f3pCAYZ2w/IMBmBnnZmHfNJ6hzvZwJppmufkDKQvgaEy8V1
sKshouhXIJXSS1GuAmpb6s+wT26Y1yzwK14tuLelpEqrxFFb8pusH675Tsw0yz6c
DSt5DcfJCZucSE/DfVa0zAJSsGFiY1hWkrdkCE+SWqEf+4n5bfQvYK3wmOnPoMOH
r/ViabtdyPZgRTnzXOMmaAZpPHcAXEnvnpGK519uF1tDnVxWWSeylKbidoY6dPKK
EGh/mc59O6R7BO7K+/qqNGUMuAjR5zcbv5MPveSvZ94K/ymbVkHNJ5UcWRfXeSFa
vuHgqcJ0H2yYHuGUDEn1XjMfP57o1C7VFyozNtyqZw1m6j591qb3V3o5pTO+tPaa
FKvTIGQEJ3SjYRXIgVciw3BHxChFWIllGWnowLXt+h/DMA0vJH+laRIKUoGa877l
Df+uEuSaUNFCMwoIaaOQd9oChWBAgNRboQiRNtkhSX8AFIIMH+RavhDSSb6wkLB+
KWqfwsWDLRkKjaslzS9kxlqkZ834Lrkq92s/eOUCRPk1+GmL1jb8wLnZR2W8+H9g
NplbZHe99W0u8kLnKFk0EckCRhD1S1OPKLf++CwYrGRndS4ei+qti3WgskxQI2fO
y5hqJXjRkCD7tpnHx1F0m7FZR8bs+eSfek+p6pRvts+jzgfl6zfaHmu7kEFU6IDq
eyi47Ld//iR2rvJSrkJne87YnUr7D/5dyj53T7eY37pY4abQc3n8MhZ2HsoJRmEv
9HVmnbJkx7JcIoYwKkh4TDi1sdSl4pAJ56AdJ7WltIOOWBngN+DqH+62jdbJy5Lq
kt+QxrDkR4g9YzGUusbxbLf1I4VIGJ0PAuypZrBLt/CJyI0BO8KfER9oLVe5VgDJ
sbVCAz5yOv5y7t+k+34GlIwQFWeFnBUuj1c28yKCWNgIGPC6zrXYy0tHfJwmMsMh
icKFCP3h6E66ITkmRfzmxs3d4q1HPOzIGMjsEJDwb19T5ofCMmQllO6gQ5m4d95z
TfEvhgElMwQaW7xYrIxskHDzkym9YZn5WDDWXHE9+C2MEp69X0FYPKOWE/fgMgUq
plqkzHkrFSmLrkM3YvkILdvMQ9TSz5n/iNY0NICLY2w7NaMK56tQ5YUopoohoGgA
6ShvQ0QBZwEp7pe6CQG0u6ItTKjC3nBZwd71It+ecanc5W6YV/QpMnEeqzvm5+OR
szzRPixEVEJGzhEIhjzEUqZQS3//hfeLGPTIBniA7FFs0bypUjcjDeCruiWtcz0q
xtlFnRt5MI7AeHxdlYz6X1n4cyoACxU4rRJFMlARy/oz3J9Y67Urko6YPR662ki1
EKCbe5PcXQD7wHMnvkHf1b/XrUC5ADiem7jIdZr8rVvMBt1tXhV8aCMF24ki0mNa
AJ0NW4mBvJuXDK7hgLATxBc64grd5q4YZ/HAjiodxAgQbVt0MD7UkwZjInDHB+w8
U+8urWFO3kXzbd2AJ3sw6wJDF+YRPGu4E1Iwz95lFv7ry+46tu4wwNUDSwNYY5JX
qUol0DxuRfh6um3EZhzJVRJuz7DHqoQp25Yr8Xpf3KHixdh4GiH/uBjMBG88a4lz
UNuuVMH25gnRYjcNSg4nQccE6eWAB5nxDx6KxTJQGZD1L2o2a3WEascDaCmgXg6d
bmSHYyadaMc4L5U+MQvCDVq7f8GhG2bpL4PIcnwzijb5QuLuqWilKIvCyc/e4y5m
93X/U2U/59kuRd+2NDkT1IYd0MD4vubmOu3Mh/vSB2a+RN+WJRP5W86zt80af+hU
EqwPn/JKSSQp8kK8tjTmhEoCtsWTZMmgE4cG7RThbTeTipMry6y1YqVqqbi8L+ez
F678l2y4U4tQBIwaU//0adQVx8oBl9dqNjXxnQtDHayKaksw5ij/IyahfJ8lve9C
6JJyIOKm4HwqnbRWC5goaIbduTjXf0nGrotvGa6VWTL1xsExXlxPnrV1rj4o++G+
033fyUetNrzRTAVjFFev/CRwm6F9idpE6MC8fx8YlpOpTvCETdhlnb6LeYZCy5A3
eVvk5daFWEGGshxAGbzUis1llGgGV+/ct4+LFCd2c1metOPnV8a+CiCF2gIpzz3Q
8JijKljT7jiR0DGBOFY+RfKvzWjdi0HvmFSToIp7yQdWHDgTwt7ScfJqs30pk2bZ
ATa+CMeLyGoNG3KBdSt5QHMSrA98E++jgChHEAgVFe0fOMB39cHXCMe94v3F8WFP
W0kTDZuU27ID6lrDi6OVZkhPfjWoU6uWBEdwy3YeKZHiABdr8WR7h+MGLj2lDW7G
VYSkn/DArKKG5o5/qCbNMlYG7endw83+LkFW9ERIHn79qh8b15oHcfPrKEXEwfRf
AH34Ku1ibR8TXB2JwjNhuOcXhs2GLrY1I89XV5PCmZNqOuld+s6o7ESXMjh0fZNh
sw8hY5fQoVnZpsAfe1Pv1H5ATUTvA97G5Kq6EAVvebNTYgEvE958UmcRqAsARXZY
1f+SKatVIquu/RdKTISWdjapjsryBTJvmcPcbYG0n4nNYDJ68SN+9xAJ8mg6uH6N
BGSx36WqFretMbm4TqkqhaDuG7jF7oF8iZhVJHHAVUeNspe1Wr87z6yyH2cwtEN1
9G8KQyjV0M9xaF2S6Yn5EMf0+IcQOL93t6YoxGmSLa8MwD1CP3KUTYzcK/T+17je
jBVG4Y3eGvYFZCUK0vPgDVjqmM6QqZsMh7Skoui+IPGbI7roMwLN84P5NvB9GHYH
/QHEXvHLCHQT4a4Fr1Ae0tXSwtCs/JfAg1g2f/PJOB8KzgDOTVCXL9KUYtsJG1wY
UNHyRd2vciiyRSSt1hZdfZ4waTEvPVilDjKkCjypMfBOP/S6qCIMBsWBl8b21sw3
5vvbGa/3zCnknyySUeRbpRfosAKDDc5n/mQe2haF/4oeJuaX9s/ecIFocwZbru68
3ok7sPDLZER0ynxYKfil17B34jIlDw8asKOqGdFP6ahCqwnWzLPAJHDc5P04rDUz
VejJq6BH7BQCm1USZSH2Yi+Q7Q8noLms3DRt17nhP8n+8ARgIi399MxA5oF9PJPB
yCZb+Z0qlcNoQ01WsYc2K2Wc4ZNQkWmvZEhzOptaerjMrpEmvAnefwiLPFXryKEZ
Cnl41+2egeLXhjPXbG9Oqrx9lhKNM7szgMWIF6qqVMR582d7cNN97t/IgdRyhjc5
xCW1/cKF1wuN1jXKlCSteS2d3/UM7DikjQaz5H/H9NX0uIqp4SyeU8Gz7/puc3Pv
7zUdCTmAyfJAY28bmd0rzVXaIaZWsPGr8ga5mhLj+Uu1/z+8vMWdiTaCAsUL+er6
kFhegdT3qCrIyvL0gYR/hhJCZ380h9onf5mye1Rf03iF+13jxBEZdlLzCrhLHaSI
R0X+Qsya4RDayYs5O/XIMXzCW7AiBD9o9wxbi8Q2JQo4gwsVdQkKDljHI4CjSzLY
+pcLtGqmM/RMQlhkhROk792DFfwlYHQXqAALystH83bjx9Vm6MpeGYNzD2a8K9Mt
tEswC3LBS3g7yJv6LHefLyLvmZnRoV0ljNXCY4dJ8yat6hrwKkHO+8xKfXQ315Hd
6mu00zxePAqF4QbwsKIWJ35Hypm+lI34DVeRLKYXYGSc5an39VS8aAE22qPIwvox
Sh8+CVY0U4bf6aUn1gwZh9z+SWHx6zkVqzfC/eM+2gtbc/HihT40bsoz8B6E7Y6q
al9LnQ+M3WaH2AL5rIUawLu/VHEsJHJ6+kILR4lq+XBrAdeN5gM+bgQmFJ0wEJ/M
P83JJlaxNIiJgWtXg3WUdpa1zE4DFjBxqn8fdDtsJBYmoxguuAD3vVp2TL/0TNxS
P9uCxcTAI2Agfu8Xu0D2oL+Poy238ZnIW7Ke6ctxW3KAj1vjHMijlvyGQ2+V0IxA
M2nfvUBDHLW/esOFS5OCeC3B8jsp1Mmov11dkBEVs4np528fJrLxhstrS8e1KAB6
dTLlhKTLCu7g6RKVzjyh8IbGU19lgH1sXUeHcpbvnIl97FjdOvfkUOQLVABONoLn
UkdhMPAopay48B6WnZQtw0LI/O13X0XXg91zV9KCqoF8p9aP8ZwUHZ3s9cwOyi9Z
VoMf/6JiK+oLzTbF0hC2PPcL54wV3XkbdfCkvTEym27Qtt2V6aLvz0zwxz567EnV
r/CrEwnt8JYXKl/9hXGSz/WcBDm4A0IHgTup5WkSPmjKmuSfzoz9YrIiL+W8OYaR
9GEQthb3QvvHfBtMXGWkxvd5+jJVUF28DgouC2iOGBDaAL4RWC8RdMRaeNl9mutP
yaGgpLNAT1WQQ68RnBlbtQihwESDIFc725zOp+jPjnPCkfJCatHX4ZLADFnqTVi+
t3FE4Ff4S+QK3yAssUkNG4wAjf8YEGmqcj9rJvxolWHZdW8eLjevCNew9816eyZu
YeXkdsYZDU1TnfLOb0SHQ/+vwf/8AXuL78d3+07SeAeQimXGae8nX7zY34aR39xW
FN2OhGaUZnGD9rFie6fg4HVm/x6gR1pDPC7l5bmD9cpHOT/pats+QNnoI5Sch5pA
DPUuTfD0HrmmQTMwcC2lPiBWWnvOTnVfKceltaOOc5JAgsswJ/Zs0sMLAmtnGoU4
Q9DG7DA+aO0WMgN9nO6vuUTaPQtN2JMNS7jcREv3EsIbhjWmedsmTqB/WlZmnmhB
TkWVgAwSKZhN+1buOUU22dU66R+EgtVQUe4dFQsEGIRkABta0FXZgZbSHBo4qvjP
lmsUzko4MIPb950OkReYUuq3DT6NrWfX9e+Qj8ff4/eaas1KSFt89Q7i73KONC9Q
1g+sH7pnDm4NsCEriks9qyavxzZvHdmD8H6OG+tPwaQcC0bpwIt0qiax7EmBk44f
/aNCprrohP2890+WbehAPAqqdp6jA/J+QMROwXaVTKRNDSKy3bYpiPKf30dghxrA
/dSMniExd1xaK3Oo84GfySb1gHdBY7x6wCRk2Dlqn3sDhj/FUVPs9g4Uh+niWRcC
zgaAsykXr3VHQDNDPIinLEB0gXikG8FtE9O731DcwFc9rfwGDPnCkaTJ0LNvxqtk
54QVzkSpinT2RYJQx2eSEnyyhlONAPOzeymPdXVvfNCG7pr/7yZ8kx7Ma4sdh7Wv
h/wMteIZSqXjf5e5eOQL3pnJMx122524qoUaFSdEa7baF8bVzmWfjZxL+Jg9OIJA
08aQ2z680Xaw2SN7d83JsPHNDqJCvQA8mVLncnObOy3ZNzWwNnhbkNOVb0KrWNke
yeIYngucbOgf9oTAPM5YPtA2CpuMRh1+FQm6gq08LVdNbrJGw7Yhppj9sLPhCWH3
orLC3Fh+vGznFbSYfI7/VLtC6NUW1NW3qjvfRAmgYszY5Xl0BZxOS9xqLrq834bz
X5ZuVMzoE89bmEJ7cFKI8MyTAlDePL0Ma8bG/Zw1LKHTN+FdOlMoAslU/i0qNvMt
UXXQ+gOL7Uu/vkXyRF/bwdzp9uje+ILfUd2ugI7qKnIm/eWKTBYTF1aTfgDojdW0
PZUt9E79jHUpSvUIJB7+L2uSYWZeXnEAO3R6Y6hh4n/gnKUESzuX0Dp+ziWoKtzd
rmtpUpeBMsqhq8fNbVBCGk5lNlTMNGGGDvgrDXEK671auW4pmPpJag+DqbgM7r0P
rjL9ZRvUQ0ZESqeq6HiOLNwKfdu6tm9yceY20rerYztzyD5cmrbyLXonpnq9sldK
9kcN32NPw1dHRWRvS4fyCb617GmAPb3IiH7PhWWxQ0Q5cr1Q+jmNTC5PWOCmCNsg
ubxmUHwbagmMzaDGrtZg8afeypW6EVA5hkkHwzZr+4d/qkpOM7AQ4X2DudUKM7JY
Kn2RNDSUXxB9fgLLlD/GFsKqGhB4NUnsX5WMrQ29xygjbhLwDCNahBXp5FpQ1o7z
FsVLj3ioYWIK+YUX5NZTQTVXeR2zHUsnkXb+BUjmTRhlb+vdAOATYCStPpMdYSCH
Bdh42SY02vQS14x71FrxoOoaa8SFGgNdZ8TRmMv7mwbZ4LfNq3DaefLREihKqoN7
Uov8OTA3gNRg8SvIG0OKPhJkaj1PQy8wvAeVRaFAeuoSASiAskd19d0iXHaAxKVz
KHuTpnAY0UspH02nL0JFo6Rd5j3wcS0slbCJMwC/grnhQz1hPWqyVqY/2Gp3c+tL
V+Tuw8NA6dwHfpqpttPHBnUan2hGhQiyZMZYKgggomlki9Fx01pZyCF/iPD0YOov
Gg42mTvxHYE1O/B5tiNVsBwu6pHOfUG+mnASFfEP2S30nNWF0bOvn+c7Mf6GyATR
DU/j9YAJbKFLnanszl9vwj2h6rB4cP3LEbejCdItfHXIth6YYHxrLbZsz6WovuL9
oDQ06xKiUANnc1qBIB0egm/sP98k1YOaHJHQW3VF8enOtHGHg3xfTZg6jhNphIBE
FFimAJm3mOSxlCZgsChQTiNTIL+Epwl1XuBXtEMD7c5txnllTp6X22pFkm3AZjuf
IJsS5zgfTjumlgoaIJdwpSeC6SVAomt5Tj3heuSytpUwalgWtE/ioH5nDdWkkS1W
MTwfapbzbawgUQEorW7bEOmi4tlSFXmN8KOkKRq88ItRIPP7H6cAdXi6Lb8Gj8xa
eUCaFEm9PjaeJqoypEwbEs2fEIiFGS/jwvQpU+hxoDJEUFXgRagz+cEeGJDsK2+G
c0EZNUFww+Dh+f7M1Zchma0tz+feACuYo+C0FzkO9VD1Myc/XIrYRqstG6cqKC8t
WTsQgIM7S/O/s2/2DHgX46m6bn/cXPoTsGOovSpJWkp6ZUw/Xmd1h/vqVXkkqjvP
7nO08RlsNCuxb7wEGxGkCU/WFM61GQkVvR/I6k8ev/I9bnfgWqS2lbdQtOiixa++
XtcZUxxWHr49YzCUBm5yuZUAkvFybUsa/Pdp3eOJbfn9g55JybtRxMLt8hnoTLl6
hDVQVtkRs3KwSZwTkqzlOejqcnMkd6TjzchbEJVyKLkFANCONA0j9YilGwe+JHvh
BTK2HJxgT63U68RPd3R5pr6s1SqxG4+nm+SzOX5DXEqEvae7od6apGNRkmyaaTkf
2IIzkh+XdbMk1LNij95IoN0uoLIPzvCjSczUwrYtGV0uGFmWuG4FT2m5/3qh3Coq
9cgDTADjn76B3mhBkDVfxbXeXUEPkRN3Vq66uH+LsHR29PFoxcEFtbBynjF+vxzZ
Fr9WIJHYCf+sVr0eOLCDU5Jp1UxbSJXjyrMYhcTEfu+ApAlLYrI4odoha1RUyClX
BuYuC4EcbC4DMLPlZVrQdSrpTOj3dYIek5GTK0nu9wLSfuloLY04B7GBAZUfm6t/
KNxX5V/UM9l7qNXWohbzXiWgEpcSQDXNaXooJr7cDa+Uu6O8WzBY0M/M9MBBtos2
UDnZ4kVnk2C7JPCSb2qh/qRhVNt7y51BRaKzNethA2clRc460vZlh/aEFPx+PcHx
PDuzMUvw3mveIK8bGfUApD37GuDw7vxygs6tL4uMs9cOLkoJlkslzD1o6Hcqx72G
zCzdhLsyijtUrPktwiGJ5PCMzLYey1pQUSZpIu8F9YMeJtDSzGzm5RCORB38aLsy
0jEHLGkaaNREBYSq/u2Q9FxJaFCWcEz4grmL5UUOytYz76MijXq5d0y8Z2a0rDLb
zhBoVXHYsHh1kHFPEbcb6udLBO3VkgQc3W111CD4qXXR7eznHxZXBGDd7nd8xrWX
FrZa+2+XDJ69R6nJ4ExT36LHrQtwyx5cAdA0BtpGM7rHwCvsfpQAlkVW+sSW339O
ZWmpSjUEReNEpf1hQOmMWhGqqKYlb+yMMtgVW2N4XmdC466sM6Igp4h+C6WHnLVH
kDMlrx5QgP/jVETALbWwLx3cyYkbHhPCYuwap4yOalheLusVcobRLNCHnmnJRgf7
FIeVNuj8H8Ksb5G48tUYJBRRZf/DnnEIGGA9NitYrID7KZWucw03ILLT2XYypSPj
1OAvubULeV3G4SKVIsJAx1Ur5K8rO6dScRkde1Bv2ibPpFhlAORJzC9YiukXT5WD
Foa1ItEYRqdagO0ZITpar2yakxFPdXtYl5U5/vva7AiSt2VuDDbA88KIL0WguOWI
W6DQgUb5oQMVqnFEfkohS3tz3obzNGi8jn67fcxStZhhb/NF7mVqDw8eZ8eBrd6A
HQOmpKc/u8TLr+HZBQqcZ2GhXSIBL+23bvQ/dqloZaFb9ebl6UMIX7WW4F7UOXLK
1bXhiVc1HMwdXHgy9p6FbgeRMfPeC3lExZrt4tFLmGeLGZtmraMUHJjjp/YXYMX2
e0LwZc/Voeo9Ah2JJvnfVP8AGr+nNmxpbTKoTQrWsdLC72OE7kz5F2BBWlbKl/91
d9Edrg8f+LkpuyxSfkYju05pCxsUIRqNXDQLD0sJDgjgXRAVcRFO0tylTddMiSf4
XTxqglPQ2/JMIsVplTGLJIN9bWbUyErjiyEDdTFVfyEMusIHvTn8MM1Qdxrf0Gdz
R0B0iCGLS15QZr7Cz6+oUagZjMiJRcjtk137zDl3FSfJ6CTLrOnE6ogz5Q804UX+
+BvXxtdP3tqA1pBT5ZSrhvkgIHij/9kA9Wv52GIPuudzI2HugCNFcN1s8oUvPn0q
Fs+vd9L5Yfur93USYjD6oJSPKNgie+MzVkMpWaz8mX2hjfgpXZK6O5UVmKgQADGB
LFVia4c0FMblDu/mTK7j58RLZOehc/tTsdnL6M7NGYB/sRtXCAIDVPrGofuBn2tb
vypyBKTWJGDX8riB+dabWKvtHwRtL1sbCxApzAunAIl4w4j7iYGwN2Q1E7Y9Kl/Y
RpY62mZr60/Oihd0w7t51/aG1o+i7muWaCN1qYeMYAQoKfV0WVeE3pB23ox6Oanx
ciWOypjnwGDXT5HEXBq1WCuYL37wODDM3Usd7pCR31hmpU2yQlkrMozPM3Dl3rch
Kr0HXyG7yJPVNW2g8uc8P1xGHYx5vOuTioLPTR8AJgEXAZJ/kSZwQT6oYMPCqcx/
Bo+WT2c5mw0Ey5wvTS+t9WAMiC7m7zQEU5E08gLAKMDQCn4ZN9ZPPqBofF4F55Nc
mgl90RR0P9ymYak1X3AebIlja5nwMuhKs1ab7p/62oAkSAG9HyTA7X6iuDJV0sUG
dvhgNbW6bkKVRr1r6HvmBoUgwHmEn59+YyBYsrlBOHr+DUEeQmYatMT+elV46QBO
XYREDLCTk3v3vvz3xhlKfZgZdxrSmOMFCZOo+GXibzV0ObfyQyXEmfmMJMDdDL3k
kMi2SSFDn7TnQcRAOdwylXQl4wIdQLyzBT33iuqtFAAmqZUrWBm7m9t5swsGZP14
fm47/vAKqPT8Iu/+iwzUYhPTRQdyeJplNTjCWU4pYjM7ulF7UNCrQErdiW1zEkp7
AYntt2EO8QbShSCfrJYMWv4ukaoEFSxKrVZ66C4QAInpSjGgVJ3zBU1PPFWVQOW4
dicr3jvftiG0mqMtBeIrPXN+JdpjtlFgAZcHpaKaif8wjSRvkL02Zv/LBUTw2yHL
xEcMgqc7C6cdZBBneooWyInO+X70DjBQr4LQQzRaAIF7n7UXlyfaNEHl96vDxbrf
d0Pd8Ggqzs12cw7aena2+iCk/Ab2733C1ekmHFL/zFsxhtn7WFd8pfmGVlfn563L
8WaGR52CndE+b39AnUCWi0481Mmi9dwRn9GJf2MrSpdx83oQgIuU/XjmZVXs3Hmd
JCRy+fVcUzGOlOE/4pXpjWG9t/myv2a1EEjTVxHtn4PtaSoRjsEtYreapf02461T
0dqce8zGBUQy7RTThy8sDcCn6TJKIpCL6rw9OI+BAxLAwOuyaVX1xFKLjrMVWI+M
txsg5qbwMbvuehPI/G5D96Skty8aqQA1aQJzcUwM3xrSNciXlaL5pysi2QyNliLm
77QAc2XkDJLojAD92S9fKJKD2leFyaCzpl5/6aQ/YROS1svtDDAD137rEsHBEBsz
9d2W0ZYhBqZ2+M/AH6r0Q5z/DUIIDZ7s49qVRnprTJos9YbgkyXscUpVzq8QNtSD
bHnL5OcdvxtUAAuBeJ/ER6m2BLBrxY9gzScx52PsjcDICay6loZhJl57p2Pwh6/N
8RCQDgkGUzzgpfHNZpwSBXU5spoWnsy7owVBxyBsM8BQq9BZR8prI/dBRiTjIdZb
dqrIgLj4I2CzNYXDba8rITYRNkLAaRh2KdnrTGEnTTwcZUxLZV72STTmPYcThycU
W179tKDJ+/0fcB54Ke9XS3UNltj0ib1cCFGbiW11kGE9iHG2JJ/FzcqFooC58Rik
hACLCu6MxE3VFm3NJklpSaScfp6EjktjeGC8YpDyS5F4EIiOAvzy8az8eG8NYDSw
8MKwnbmefyEiaL3GEbYxghjOylicXIIF2MdBLvqMQNYVkjz2Uns0uqHZaOReseO4
Sz1e5NbKRT3nN2LYvr+Dfs5VSHO5R7Fa9WsxbGalx0FK+CMcpoMnYfRclvLou23I
fmipsWgkaKzpgyGnaVav5bY8dTqTZmCqH3lpdbAGH29LrJ0g32wmfRYy/Yd8ZlRS
565hEH3FFuHOse3FLfIg7+fBs9RGmadOIJ5fRVyMGY5tDBmeL8ntO/JmLwfoxnUW
CJdOEc/+fjtYZvRCwY980aAs/oKLOd7dkpv1+FO0pwYCt14A+Tl7sqZbVLXqKl4T
aGWggI2FbbWQrGFacpy0K7olJ8r3TvZjaWc3qaWrwWMUukUxSB5fgEaKMpxpI84i
XSf9+4CF8ROG3WO4goGukbca1r1hWz4CMuN9kx1Jcozf9zZ3TgU44PN6TOC+CeG2
cgGraqU17XVT6cKOz65hnL0Hkuc91sszfsmTtRZkzZLmj1TkXc7wCyl1SjINmdts
DqPAs72V7XlxA/Se1lbTvLfCAfdUtAdQ2tfZSTRm0Be4ZXkFCbg8B6BfWIpibHe8
W9/yO4qtS2lJVmf5L8JfohBoGHY/ggowKoRzmwmzPWuG3p1EzeEi7s/4r3vfMzkX
e1DEcKu6PtaAkCP+Mnwn3d8weLVfr4RHzKtc6uup7CxHVJegdmE0xYInFWjWoa19
lMDO9g7ymtY1XIEGTkJZRNVpWwluUhML42SchLjM5Qrw2vdNR6XCIN2KlFL0Z6dn
AwLMqgxtrDhvkboYr0TVCjJeHzq0q8TYsKDC9KApAqddPmzpiKsh1Faj4F/KSpgn
ksMZqjPeXNFr+VHV8vfyLqNNdKtKXRGJT87e02/1whV1hgZlspZfBCdtpHNIqhFU
NX/bCVqPLGWov0SelPJgD/ch2i4HoPWPliQ2DSKA/a2mU55kWvVbER45NKzgKNAv
KcBWXHi7WF9O5qUL2DpC/2k3slNX+e+wW2JYndLzDuiJRFcQISMwcgGIlPTMd1gk
VQbw0tC+K8kjkA4N039rCWEX1KqpWSlXkEX2y7FUu5/4dn6tZvROcZg0zzmjosyl
k5KzPxZqFim3t5dqKM6MgKkNaWVhQ6n6ZfqTB15rSOaM/FiXeZvffhdTOfWEl57j
hU9IWPjY3PjXIxfVe+IRq5VYn+NMUlhjkzgXVtqykaO2Ur0WqJpaZIBJ9X8xh8sJ
bKKK1E9ENlIg0/pVFbyp6KasaGP8+YTvsgDNzbMwgINW6rZ4YCW1HF2+AecKUQMT
HNpMIizjJAQbB9VTXPT//yIm/g2fNk29OvOknxE4VIv2boLT12LNP0GrTLmNDP69
5VbgtlhPjsgGbFXIksTfqii4tYqqMpLgTe0D2Ys/0L/nepltIzsmdcOH8NaSf4Wb
/0C+hQkey32SleM0UQzB11gAy1YAuy6Gz6ZsR9VLvMxvk5a36rDQmNfJ+1BUOhRi
ZtVNktH2gm0FHBn7cATJ8UU0qaOWWqMpk+15z/ow4lUOY4uqK5RQhw8SSgcLJMdR
3D9UPG5ijRbN2uR77nAEKlLqdNpHRgyUQO9UeczyRCR+MAWGkMyfyA2GSfeCBFqs
CkkE/+A3ocBiASKFJ4Aqx362zhqP28XWEcafDeOjqW84rfP7o9yNL7Gbv9c6Xcoa
U14ZGUpG2oV/8V1bKv+w3Cb33RfHleWrfZ6Zyhag4KNWw0oGQZUrI7s5UU5QcRxi
GzhuZfs7QglNrUmPb5uxphJS2+Xv5aq5sTt837AOVi58nl1Unw95DDoOuJFcZwk5
NwLNxkKfqqslFX1dWUua/fTkSzJKX4PXv2Y1NgId7N8ctVnSNObWPeN/2k2ZjD1n
FNVSARKmeBg4OwscPK0gkuY6XtnwHhy7I0OP2+51K1vK8JR21EBX4j4Mu6TIPgMz
OKSZFmYemowCPA1pEO9KIBTum5EznNy8rbPlyoKIyKj4HIAo/cIUZkmPyYIAUWJm
WpWNUS4ERmna01Lemh58/sJ9nsq7DMuK874EmQWjixjY0wt9xenDo2FX/c8gTXOp
XQAM0+IEMplqSbZYOl/EI+QsI6nQSgU3ih3+WBrMxCsiiufpTT4CtTJKjK3uzBcF
MCjj9LUJnAca1npci2TUH2BJ56Wt2fc494OZ6DbB9onS5o4rZl2BzG/2Gx8E2OoF
+4C69aDQTg2+9EAkCBc3b4bQy9vEYpfOYJPy/j1Z5WJko+4bcnilwNbJmhubXCk8
nSEmVsgvH0fqRVlBx1nDJAq8nBraLsOnHJqAm25cjuKrbcy3r4/lb/ge6seoGjCb
xUOJN7YqwcJx6G/RhzcC/70H29iDtmiiBe93lsfAJ74kr6FsRmCxSMPb9gbLxi7S
0L4Jf1GmFaWzZ+5E8xBK9jpnI2C23Bwwi/FxXJzsbh2yie2gaRJWIRno847Beb8/
f/1Zh94wx56t2Ra63L43teBUzRPAo4j/UIbtZUoBuO+fbCyd2r/WtPS7QL8Nmf8b
LCUb+iYjLXgtg1o96iHwlGSBBTOYpvxH/b7RcCd7el4OyrkccHUG7sDGy/yaiP9L
OUb1fgOLnQIEB5we7iOZcKm92zkpxkMGomTT6x6aoQmhHdcZ1XkHEs6Pzxaj/jCm
TcW9qByzqX/wSFW+ylws6HlV6EenUs2VxvpPCBcJGAhPQ7nEGzkmErtacA814lxO
m5CCAYRKcrbhG+ddHlUIZ9ITy82xPMl6QZt4HxLfjJULvRzoJ9OTVbqN4puczplR
z6fyrleTBto751/uJKnDgh30qmyMmTd3gMRoqBWtFJA62eJycFePhfwwZJtPaazD
6z9YzTJOB+xdz3X3M7NegPCwy/PW+68EsT+NcCFBH8TJOla8EUU4ajrNNB5r28gb
KcAaS7yugBO5BIHx7/nZg8k6WrzNforgmdG9DAkSWv7EYk5ChcuXD43wIn1fW1kd
ceOICgAaz1aWOrXdg36S0kgcnKFU+6/ec+D/kt0y7IbO5FTUajw3IiRuNFajQvs6
bPR+j8kDdiWZFz7xP0F4tymkYd8IVvBNW5phvClkB3+OWRbsesGMX69j3k9sv1Yq
LJ35hqV9plI5hMAJuzqnhPb9/+zBDsbi+qdGIXiTyMqHMOhlhewAUBd683cFoeVb
tySJo8+azs/820U/MaJ5daJqffOJWUj8uLehg5Z4jE/w/To/jxuMRIlj9kxi+Na4
piQUlWEpcAys0JfbOWtF3BA0Eeb8MhOkW8oow9h0FyseoV+C2D4BauY3oHctG0Fz
ByS6ogsdGLMbCxRf2Zorz4J7q+xDzPCs/1B1rewfc0Gm1wLx0ElKxPTf3Ag0a0un
q6JfUDZNIkqfaKTl/pJS0mDdHZkh53ODSYddMxU0lmtrAWxyHn2gQCI5Ojx9IjyM
C15B3OCj+KDyrIvMHBZCE6J5kiSJ7f5d+I51D271tJRHQpgXiRbCXnwpbd9CgfVB
4OQul0k60Y46QuqIjN6dqdDg7K1V92HsLGDJdgfJU0cK1unmzOQxOjQjsxy7YoTc
22n2r/mqwfB2RdcjUtM9wRwHy0TuHm2jIrhh+X880wdwR0RDT8MSjY0hHNQQoFFR
RHEG+UDd4vje52bkPxMNhop61XeZqhGy1hVVlDLwknsSL+AjoNjLW/x8k3CkNlH8
ixmFfjo41KU+So8zjPV1ZyCcDOvZMSicRmhwjAwarHmoJAAJl2r7Z4e/ytF+Tzcu
wdwRBwgU+aZJcneepTpZ0/kYj001+SX8W1ILyDEyq37+343REnb5pbR9Ramhvw8E
4f7D2CB1ruLnC5CZlnUQVULBuf/oH5DGD2kdoq0LgAyeOAg86dDQZK2gfH5NUeSn
QIg2nEUpfmpxyubwX4Q12xt9UCamSQwKZ/ZohASrUVcwJdPl75B7T1ioGNEIO9IR
9SBp4fvm51FF2PJsvz2CS4DvVjmO8HaPbKcjRPPy7c6sX39tFvvNtwE4EjDgBcOm
5uepiifIr5XDeVu8n9dcBtr5nMC3n/xzYjEz80RGMjjCTpbd5KKe5Z3wPgg69Rpv
BLDXXY6p78wCpQSbEL5iMBLYptNtIbmQgHZkN9H0qU2CdHJn+Y7h84/nVzHRrm4Q
Hm2i97Q/Q2pDTYwjLUu2x2BeK2oIduWcRPC/JbW3lhI9trgYxHbCFBJmF0XkfH+L
PgIzT73n1tDV3QJpjE7G0PymSOGv8W7z2r6Hits/UalVF+mlFOt9Gm1Y1Ko8GOvU
HiIAxzYN+F0htwY28RHYQExoKFysf9l2oXIRXjwssyH/pVdvLSuwtarV/BUtX9B5
n4O0OU3aGMl2baJ0P341uyjabOXoltODRh9RmyrjgNSoWb/mvuOkW8HDXyUE2Hqv
ZRbvMicT4Wjbdo64Hh5xlBc288P9Tj6MuEZN/ZTLp3ztG5V8+D8hqXYcQotSW7zf
HSRTDCuxmZSX4Qwl+EDDimcZxKmvl5021vJa+f5GmGzIuwbR6OPLSGzYVJZCQldJ
MfUsOheXKOAMgQjzt89Jq3QxVVTz2nnTkuiniHfAqwPxksBgvH9tf5Mw9ATStZcE
jSbJ964VVcB8RK93AA8e74P9sCaXO7Gjmwbw98WvaifFraneQSh9FIWF97JnatoY
MUB1covwbAU5DSnYBrhOa68iuBMEjeGkdL4NrKIZvCjQLIa2cLzJWvhpJ24rTQqv
EOE1oAEOeUmsw5YT8LHMvOHslRG55y7ahGdEJHQ/WfquM3XDR+Nfj0Db6p0TAm2S
WLTQaiDV/xNcuP/4Ongd/DYW7BnrjRRCDfKaeXi409BcBU1A6iRYkZC9A1DWpj83
svSTjcfPQA3sTPmyjZT/0HUxg0hrGBsXKvWjeFtwvEPm002OSs9+gMJ7Z9OMygRO
XKg9ReATdjuv0IW0QMrSjYqqBiC+Cf0jWZWaNs8xonWSIxPryJBRhSw1jpSJJ1Kx
C4BNDJGm4bni+nsNpNW8TSrxIKcsApYk8QUPu0H0wkwJ5YoZP3DEdobNDvfEV2nD
FcLOtn5j+LULITDat6Xh2EnMEBua6X+o94sTIrCRINxDjMiytgI4B4K/I1nzr1RM
tBF7nmOYy6ALWFpwZKvaliuLH7F5mYXky/AvtEbi7pt09jR5U69UFFxiTfSSI8Rz
A1JNrXr+6+WbIYwkY6bvnAnWVw+uNihUMgdC/zBRtouiIjFAxE3MyvXpRnr4TsBz
VgLljk/g66Rse5+y+YXODOUuO1iJpXXLhOwt5mP/uiW3leyyaWwb6LXFNuGXAuKP
SB8eDqXrP6eubeK9HDgtMm2ioKbyeIOah7m/YUJ5GrR+bb5O/s59bITPuBevVmwY
4+TwS0NC6bc7b3oXI/A4YG+R6e0MJm3TpVp03SO2y2a80Xuc0zwgV4U8CrH7pFDN
VO4bl9xOuGB7zfIM1KqAZpesU/HfSu4Mq3HDu+vQjTAGsUVI1fnzpk5ezBbb+aUw
zmnvQhKjiobcD7WqUz98doppC/ebVuhxUa/ghRb9/6MKkLPZljy2Cs+5auy5Ld2b
WpdcDjggjh3gm+h6mnjs66gFNyU6EjQVmR9gM8bN9N5RPHta2eJxRLOyhskE/Fm4
QNVF27bl/Nbal9K6IqSkc3pVYDdOOtFhImq1dlomp9ox8kHMk17DmDwcNNKc0bs9
V0cnGd2QnugRTGDCq6EUuM1oPCnSmS7bzDcy/BnhL3c0n7X50ccHmjn4QL4uLVuJ
R7RJ5D9gCvrYgn4utO9wXabkl/PJs5BmBE3rQTm4I42IgcIlA6K1ojWyQggkMTiv
rtHYcvCeWUrbFOt5+/ElP7rfXjLupycfuCzqXs4DntuvtLJ3IDlsRLh1naXZ3qlh
CPlibkXkLDCDHzIG28cAbUo5ekmZcS5CBgtVIXFMKGM3UYwafmgW1KeUly3nyt3W
LyI/4xB4ODlbsqop3JEQTpje0xuwPObQZrU/Pc1AhYEF8J3qDfdqiHp4IFF19iYh
7wtF7nnDEyzW47T+VscBpIuuM2UuKj2lmCJ6+aB2k7SwU43SYogArHZbUvVR/uvE
0YbAh3SqZdm1jokcT6E5RAEpMPKDxEXluj9ddtuFm6OZecdU3GkxL/foxyxoY/RU
Ur7uxujT7bVExKAUm+1yjH6IlABYJqtRYhzptbnoEP3etCzZkE4PSxb/RSzOSLbM
CHc1CKBzsdc/8bh9EDt9TjM+xkMDxbDeZk2AezUSFvoykFH+cE1G2BrnHT4QR/Ki
kwqm5Vh5MqXl5IGNSAYevKhTODG7MX9tnS0ntCy3kzRqXFvn/VPSLhLYOH2xOSJQ
IfIw51hDGzsKADZ2bUckcMJQDY7Fnt/JT5iKPGvOxLPnWRndV+lU1BSmhfdSKvH9
JS6hzG/dVyi0YplPdMRnDrBLTEheZhnMxqaacWEOvYtiBSvuOPEg2FV5VAytPdmh
WmbPw+ZhEFYrQprEU/0xjQmFwryfr3EmPtoA8WHxknF+sshBuXuuD3ovae7DtOcO
pVaAB5nPbjn7GE9U4SmrN08yZTIG0GwFslU7Y1xF045OmedEMoJDA0f3ULcD2Ywd
uIXWJeyKiY+7ODVsRMv3VpIQ1dAQOtFfLax0QX5KQ0TvFa0tNy7K+daP4NtBDCU2
Rqai3v2vMiNjdpNDh/vS3T0prN15k9JX0jaVFOypUSEALZBu5zLKEentNBl9GaB7
3kgBOKwACFP5BX8wjvQs3BIpIrb8efE7KdKaV23WSP7BHPlupRAX8rhU1A/qGCYz
FAsMnb7whm411oQccuuog+McVZVQ2PcqxBAn/1PDPLRhZJMBy2QdGDI3P33KVl4V
o4CxUu71t/+f+zB/oGAbeJzSzNApqiWP0rw80Gx7xduIQJYKP2C5qDQeK/+alfsv
W2ZNkrWelBXuUsQM53xoA+BMRGIrm8aDsEl9nmF3FqT4Kf/QsibIzbiaD8SFHIip
3tAfnCbDfPr0EnNHB7Ezm0bOiyb/wonkhbuDEL3Yqk+i9BYbWsGTXj6Ldhd5mJB0
eGPwxfNHLIibz2pfUj2CdYMpb72xKv4Ia5froAIdp6uv44M0qnF6RD4qSFARkYQM
NIoujJQX+PGnRHUXbzRNB0RkV8qL4l0emRLv9wHSS0xvY4iCTzBE5hv2pVtJb7Pc
pnmwRHBfqmtY1cUxbDfXcAqXLEzRFwl2//XKorXSXYxuQuvwBb567mgWbyl5FiUT
g75lbkndGQua/9JxgBTFWMWHFFcO48MCtOrwU5vMfxq65vmGMP9Dl9+DWOGjs6XF
BsDV7WkAXatkU+0gMCFtRKjt7TxMw3dJ8ZKGJ/B8g5gxWNpdQTrnRPAhgxR3bOAl
eDzzTZmOhrXnV0+ZBP8nnQ3NswhryN9pfOlLEtJt8C1VnyMiT0n6aNGZL+ZXHF7w
2K4uMvcozija9EAO1pkUwTHYjuF3YeASRITZd0/zxAQBR+FwHgeJA2q1OEEmnBxp
m1DmYcnYbVoUMKZRq/Fo1aTJxTSu24MlS8ZMHQdbq36/vHEyF257Su3veAoebMOF
z6npNfJYuSWQZVYlHZSpwDDP9RrpMI2v/Fc4d15rM2JdJjhcc0MkLqgF9vshbAZT
8rJd4+TBLQdzNPdaE0LMdMZhFLdcBa0Xti8Mwf/qp3De0AxR5ZELMMYQYJso53Ig
LAPgk5AV4WfKCRh+AQ2S59Wrey2kJdhVHNDM35Ws4b+YvmLjhmIrE7iuR5TnwY6h
XCBWhWzjeZcCzwdkWwXAeG9Kojo8vH32pPFj0eoKAclF+zErIBEa5nA427KHPdpV
pYdDhigCcfTYncHcVcV4511p+P5i15B03XQSUNRcyf3gIYk2wWZlt2f9eI7QhPHI
kg0RwzyULKBpgsY4Um3UAE07HNZtbDgXW0GAoWMo/q/gnFtIpEkZCnEg9ZpmovXX
/mAnhpjQG7JZTD2+v/14J9JSSIbjC+Z6VW5aaf6XId3s1CEjDxE5W6MNigNFB24S
+7UjEzCZP6z0ujruAOwiYkq+QBbs7SoZoeRgpeLxb0j/UGqwIjh4YnrwzbFcdpNx
IkdwoW4gNkSI1eCZC69ZErLHrZy5bLoab/a5XHZq4xDamcfOcAlKWT/6/6eDeWnl
FjkIh7l/o1sYBlJJaNOP1N68Yn9I/QPdISlohvJD8Wuo44XZeHAcuSksNJsCjXNR
NZeV2z6/bmcE5zClXzxfgS2E7IPS9rKuX27mTtJZku+rxJNNkgnE0MIhybtXzuBC
whVfKC/3ueLIlEnW6mByJEiCeDQtoNXCt29sD/6gCYyOm27+Ybpyx5yRPozgbPFz
qeJ4Ofi9pawCkiRi+WJ0Q9LLdgdEyV2p4/r/qnycSFjR3zqZGTjLy1PTqbUGi83B
DM6pHMY64nJuXqolUN3yJNV6Kb+nWX8ORU8Vl0xnmuAkLxLhDpNrSwylAkOWvW6w
RUxT36gMcSVnpirp7H7lOIliaNQDZxkCXuGf5UsAo8yq+lBJldU15hkUWaMYF9PK
JlYilWmfLtq/dqtwCjoEMF2OVch/LDq1aQ2vfJAlephMx+yjBE7+Wt0IiyGeLtsj
cM3Q44EhApR77++CEpVxw3wo7xB4xC9MkQEk/yPaSbPZnCKF/Jn8sC5ykD1BJeFX
4t3DfdHP/Mq/834GqD82Kj9mq6K8hckc5GHLHaJTRIytRwZUOu+/CbO/hBrx02bg
Xh4Q0qRCwZNEnTTFBbwsItbb1rPzFUjNB9qmtqtBVog9LqR/PiwzvkuX/TDrRFyP
unsuZNPJ/mOqnyEH3Kq3m30AtJCdCwVQnM9ht/5+WlWhzFz3bZXYNlrlWs8cU5AF
1qcMtmOlgKihxfzKmCQMJmkXH1wZclfpcQKkL49VDm0jp0AlpL4p/Nn/JXJC99SZ
7aM6q1x2gg54PEOZYQb1jZKzanOkiZiP6QpsJP3LbuFW20J02DHXz1Yf0r0Kg0Ox
36sGcv5+zU3pd0O0f6R2KTdxF15m6/eQaHniZmlS4thx/I+ufh5RZzbohB80QJc0
8/APuVkwZKDxlmRoXB6oVek0X30rHFJaWZW985kyDGRLSbL4Rzz6vcEPL6L7UOEL
f82ahzGg5iakI39CFNLaSaXWx0Mb0S3oOT2MxVnz1luEDdBXKEix28jqOq8K9CrW
hNLrvXuO0m6f3v1CKdzvEsqBCjXA34/CAdzET4hdfm4bnEZnowA+HUjKWjGGXs45
B0ZxOJv39b1VV2zQhYfoPLlUcxTlkoOjgvRwdqGV01F7O+aGkIM2G80RrDJeoWGx
wOLgt1IE9JfsHdfQszhQ4b52xH28DX+lkXcfggP1ISRsF5mRe+sMKXWthFzNwxaQ
07+tDVCpph60HJ+tscvdEiXQqHqzYaHPshcG5+x4TW0Xpz6nJ/izFwNR4axhpAFv
SM0SAO4kMQ8I1nA2yy3jXOijY1hd5rPFADJNDXmYCWlsJEqLqW6GpU+UxzjjnvT+
r2xl5tVjLzJXJKGHUth6Rf+dC/YW7AwJUVTLFdUndvdSknCso4OdnlvXfKoqUBLn
1WXi8Iq6J8wY7stxiwf1GUQ6SscI6Z00t/w9gfKOMeO40f4oxq84tGwLARLi0YVa
BdOWW514Ba6kQbubc0hmeEG9w+64GTc9+R4bMaUmtfjpEVqzlYZPq0v/VdLtbbrN
dQYLlRI6QXWDS/L2/iyFIbwWc/cqEt+plegJM3SW1M/fVT+v0jB/NJ9J9xkDF26r
EhhLhn4CKAUhhZouC6b3mrajDAQRmmwTa/beCl/7d2yI4eXPcr5OOyxLkYhM5pYe
a2VVXeC7cKIAjAAFz958K5WyC5Om13mZBBwo7GpvXRILJ+hNoeCnFEYsG4Ovo+5S
8Xp+sQ6XWuC/bohZhdGgL3U6G3yU+EfggaB9KH3LmG/ZqZJlVZ3hBIuLhfETiHCK
qIpXI52YBhIqm0zNnu77iTL7jhPkhV1uQOD1VPm3TGNEnPbAywppBesLQjECAZ1j
RoDm4pHSZ2UM91FDWR+KP5y8jpsXWFwifzrcAQqZpMfFy7sS/ijXhzbd8Mdw+vwA
BpTDRJkOQciEn5wnLa03llCpGfOmX9G7UvG9CZMZ8FCvDVDnxXMtevKfsJpJymIm
uNpQETMR83gdEInQ0YF/bmCVRuQYTUlvc+XdRtgJUX3CtiSOA3Q49FwV4Cjw0SzF
d2zuK2d1cQWv/EWl0OhLe43ywvT8cUrzKpmurm8gzzVthnTAEAnfoRi3yyBZUz8D
U6zhGBgA/ApTnKM/t8KxcWCeD4gqZJNi9rIZ9Iy6OfN8SIASQXk51Ze56XmF2doY
3B8rZuckVKvud+GoCLbQXiy4B1Qj+obtLY+YYDt4iilB/7xzs2KBlbgTgHtAnCZx
ofVN8x2WwR6R73pjnavrXTO2iwvsGgO9RtVFgsWYrSaDv1bYZrmCE4JePGUeTBNU
pBkR51BV+WodfeW24qfIUT/ArjCxSovvuWzHnV7adCvs/6U12MaFisZWInKgGorD
ZGj7BkM8pVD6mXYkdkI1mjCeRstd6LmTruV/mjdOgir/46/okQTJAkOBpoF0pTtX
xC01Xezu87LMbm3sqHeAlsuejhH8hwncdP/Roityf12tPmm6GZ8XFT01OAawVi1h
ZTy8TnhD6fnZANlBMoQcoRlYwPlLcodsEOx0wCY/o6Se1ZcFDXnuhXy6a2I4z2z/
/y9fxSf1CtrTNzQoSDoKEeu3ENqQBkTGetz8K1F1LY533Hiiel3cP5mFSaqSlmNX
SXGNgwpc60E1uUetF5UGPdZcSwGAapn+7px7Pjoua5SgJ9UdIiNYydG0gb8AtqOi
mmaghY0VTgPDtygM6OBJ1QTopS37oRSVHMcihkb+hk+CdIf+NGLc6obNud+X1H27
DKu1e23PiAX0LWTMX+u+tB84XxqGGemDkVLHhgqZ/1Z8q1/GnD0nbPLcxUophG0A
gZ3EIF3TgG/XQ/u9oHTvpEmSk7BDqDASZQvYzH7itcyG2CkuVEsX3aepSLx/IQ0i
tLunOOeT3uLx8BPZ2ptZIamS4dm9MnedcME3Ct/qj38ApBKPIGFfffYtdAbGYW45
mJ9w4yitcaP76HpB+zxbyzGGbIApuqCYIaI6KbLD39CpVf6jPnpPpi0GCHnSMYo2
3iK9fOz+N6VRjrLPtTTmHmMzScKC4qsD2gRyy5LZA63F18XfI1pDbOd//3DdxGnR
oSHxU3ADmnWoioFLmd73aCYKOuyiuRTMEzzJE3jnbQ1knj2a2p4sCVilz+NdpWl8
De2iT6hlpVqfzhgO/jB0MuaMkEF7I+wQl4xW+IhGMQc/tSb8Pi2Fkn6Q0QFs3mZW
4cPAa1XNl1x4nPt/MUts0NLfXd86EnkHZPeSrOAz7b3YXvn6rIj9H2NhyEMFbCOE
b34/5G0UG5l87v6czSyUOlTvo+z/xh+prGBUh49tAk1PLLIitxHr6iT667P0KVwf
qMudovJ97FOk0el/AYohb6xgx6I3DXjRYdM7I5WWU2Ikd5HOid0r0Duewk3qi7NP
iY2YwBPcwl3TGyrlpB3o0KaAlYa7cexuCmKG/e+0uw45wrTEUlBT5lFCueFDSHgk
dBLCJlZ4MBzoLrwQ0e42oGwLV7y+I3Df41+kzVQeCOTgw2adBd9f//MX1gLwduwt
FWqd2J7gpMXGIJ3YkDBxGXx3INkkYpX4+RReMVepGQp8/MEPVKZR50Lj5y+TJkDk
1Fbp28McvIAoPsJV7RAxGpThM8ygPoyrVuzGSCBcrxkbx2Yak7zgwyldpJcMK/V6
SE3fIzEHUiYOAMLiiyUprC+uzo7iZ4aunmVBd5V0COVPRMN2ytTLiO4oA6sdsnQZ
v6P3D4xMRVa3Nc4zX2uLIj67eVQhEdkCNICqlUMuW/bCf+HTxH5Y/Vdt8xgKrDhu
SGExAUhikWdbkgJ8uIrp7gxHZCIoF22T8VjSILN8dCzCAYAI9v0taonwm5xmqb54
UJxhLOJPysbjAEOmbomTX6O30JclMbriA4/LMeVqZzv8CgshKlCRivnaemedAD52
c6abhAe9NbHzwslmzPqBHweEu3fytHYSqAfYvrZi3RdvKYuleEtB/7F19sFNWqym
isZU++oascg5bl60kzdKKF+cHSMnfnY0bwbT4rNoWwN93xzuW1fjoim+V4GHr5qd
ZSmtQWeU7fYXol9USP1r7LCO/Ng9fhvSnNtV2B1yF68/1+CJ4UZLWskQ0BqPhP8W
Dj8iDB3h1rRkV4YV7DJpPkyc0NnKAVOxVODzCsMeC8eiGtNvY08ZPSG1a2GM+vdB
VnNiLxjEsixguxi8pVUzd4ya6kZynVfENKO1e1QT5BPGPU6uF4IR4ak8iEjGhEKd
T8BEuhwGzM15d42BqpXboQniex44zXFAuyk6Thqs/nrkpQDlb5quLUJCZZsgUPsD
1eRuhNapKBNXXtEQb+VzF+rFa9emMPwK/S1jqu3ZDUW902rzMQ9RbfpOsAF/e5+k
CDvAwzTdMS3HiEToAkx4bwA1ezeFhnAKZ6q6IEzdFhlAhYOWGZ5vzxmVxmP8kA1G
HWNVp9+pZpLEBxbbPR5RXGPCOXt8sSn1hUKv5DuLkYM5CHo9mxz1HBBVqOe57U6O
xXh8QutOpk3ajHz3pTepbrYICLtmPVRAImkH0Yjs9ukHAL+TGRlmJaMDA03v1JRZ
U/OCzO20/l7PHFz/y54v4jxfVw3gdEkbz0fjKMIGujncHIvth22D6ZRXAbHlG771
+4IpBehq9m0ncTAycy2zwgCoID3AF7k0xTl+UqtUxBnK7bZNegm5qWlPc/P/3uVm
3QCa35sCcROslTqTo/QqOdILW+xWY8ZdmztdNtyHYT+skzJv3HNWEdryoEVTeyjr
CpSGREiGu1AqEVDSwuGV9Co+XEQslIASod4Lxu4HjnluAZ9MkNUnZgvgViUa+f8q
RGkGFR8norlx0Ss6KQJHPq+bbmkXesm/9SVAT2lO/BW1kWJSD0765OzWavCVvKe5
oJ3IPSTu7qCEmQGcAPO7m2DzOxTsiyfdfBLjkCnoylm5F3BtZSNZL1z5kj+6sfZZ
eRWo1gL3v0fme90D+85AfK2Fycq0DTkOdLNte1k5YE7b9JVRiqChBisjSY0FwP7H
N+nJrrQUxadwK2G+moVkvJ5DrI1tcQ0qkEnRG1rWe4xVoIDygCCxz3tkYSKu1IHh
rRYp2uc4NUkkEMnqJSeCvngx1cONg6LFMJG1dmEHvdTWdxxvrqHxvAxHe//3sw0y
LX7afQyb3feXxt5byv3meUg6+lo/aHVm/bCg84gkZSUUglFDl2hE7dGcPH5lmZdP
wyM8yWlYCBvdB0wQP8pj8ZvLaZbnz585Ej+ycYHiTRiKjOv/n/T9ZApKmZPV3WSS
JU1X4jIduLtuGxNIjyg6vurWtHsZImhWn3PhGe6aeu5SHl2LssR+c7u6paNIhHLf
93qsPFDHXdexWJoRTZdjLS8iZreXaNwZWTJiZbxD0gfTCAYyz+K1rFhmTzRLQx28
1qjNlj1D9E5wBgfL7HRxQxv9DoAm1m81tNhpCjE3XjFPAJT6njH3BWskoXWUZTbV
usD8/DEBlvE7Gl4XlqRuSGYwnNeY5mFo8kH18puFhPn/h3yA+m24Sr74gOe4ZGmP
2dwcvg9VaFISbnqT2/0ZT0zJJXOSi/qmGnlE2ugsGBG354UpcKWinNJBDcDExpNg
RbKD5XzD0r6n0D6T25MZB8QO6DPjrCL6owzmwoM6j+tBd9y3BrrHnHi7DkAce1Tj
PHobCi1stgKe6/akZ8bjD99FrHTbQVuThyRmj2RyusFjbuifBrgYC4PzYgCtrCEP
eDjokhnajRqbhd7boanMeZWMpBGiOMBMddTlIOOqSYmq3lWVnowD2CWmsO5k/DSr
sbXKHNxvjQRTjkyjCi6cCSTF/2ku53l30SW26PTSZaRVKvN6S3LNLsCjiOIFx2iP
yfbNnxUVEvMVMXTB090PF7UXLNGnqcPQDOI+EAJPWN3kTilVHLK2OU1Vjn1jAn07
ioWcX9bPBQe/oc1jttxFEQfbgXkctKqGlZ68kB/but126APyB56p/VAyFFIwWzYO
T6fypz5uCYvROkjYrGIEF3kUiWxG68vQ9hWYFCGJJ2RmSKlNBkDAxwyqLc17wx00
qjRYjLHVax1rimFbbR6YwwDJSQXq4R5qobExdcIIUbADtOZyh4CgvDoqowj8MjSZ
bE4ybkaaOpvNA1zbmhrkKdXziuOWq3+XXuRBxEx8Ac+O/1LaOeFc6rjbhG9oVhr/
dl8r3a7yc9DWwBulqoQCjrHxIo0GAWLOBbcOqXSsTBupP5cvA/JrRHNBHK24SRC6
B1Nu8z4rJ63m9vLWReF5yiRWLJ1jg4Z4gxJu/NNut347CWUFtQHfoT5TO/VM6B8q
mK/dcylQMXwTGxmZTdyec11sHbmVhsxBMAoECx07OmcsEpf1twaELXw1iG/WljpL
S0uPDGiCPDywec6g9wnEDeBDQxiy5lFDaNy3nr38VYnbFUBtzct1Ik7OGWQReVjr
KrumP8HdqRxt+mdw5vGC5BH/QlrPauRv8pt9gPGOkPqo1venLDnPgY/qT7BFHV/n
EixUut4ehzE0YwwmCbxGJ8OH8ERfWRcb3CyFLEQ4SYVVjXAybDhmYrWzQ+Qp5JD7
1fcVe/qjMoJRNUwpbCVmhPjlWu/RxmGcRcKi/1Z9J6JGjxCrNRApfV0RKe0ZnFJ5
MEQjL4y0WGoz5J18jliE0RJXg71LKcVt2wDn80yVdx5AGK7SGVhSE7VEl8PIzjAR
pVIPbvs6487Bx/qcowHDmRycTEfWbjLluYdG3u4tW+As7bWxwdvVEoELma6UxSzO
PQykS/7vwTFdFB2YfK/+KvyTmaK2JesPm3qp+QofLvQNM5/jF4+84sRUEH42cSvj
k9Dl2t1slSq9JlHWjfC3b0efIk3nXQEyLGriJHbYi0dPHw7AD2xOp7KcbL8e4IXS
GOewILiho5mNQ10hUVIf0yzcS/NEw3+nCEiN7YD9LtRPt/bRS3Df6AnwlUDk04kj
p/HwbjJ46xjocq+bRZIlaRfVWgBffkBwsAZt8/kDitpBTm0a3oiZfGDcuPwgWwqE
IWbLQAv//gR3NZnDMRAcnX1ge2jUcn0uPoBh3dd8XatKqVblXJysBFnFVTzdRmbQ
V3QXd/JT6h1/WfN5V2wstpf1D8wJ7ZOqoUv3WyduZ9cvU7aY7t53BnfprxjtG/HG
HUpnH0uCSADEmLC1FcIPSLuP4WG093jonneLQYKVNuCNQb/AwunP2cRvLZZcGmoc
gvr9mEmnsOpf0Eg3HBu4Kmgt7WBR40O9UHAqOKB3f44XUMLAfDr3DtnZNcm/SSC9
ZrKj8RgUaOpZaaCAkNSgJIAAYAtZvtNOIFqjERI52keckANzg3XCOkUfAe4corRg
6wQPjEUldbLYFO+dCYoBIOv/J/8GtuEc5fI29YERRH4X5/ardZCume6VqJTZ+yZk
DBbHvyDN6gwCA355+0a7olj1nvAf7MOUmT1JjRH2PFo6yB8ob6xAAcNw+2YiuV0c
kq0Js+JPVkEKQfMwfM3WQedy6bQeZ/DpBxkcqvpeOg55cJBMzDmrw17xDO0iCPt7
IwFdDNbxj8XCV6QwpZPjwgzMyFwIsrk+j6uqBKNtFLGmFcg/zIJ0xwG8P42lxlQv
3MoHRlZGQQUvrihxdmi/Yrkvae6j7x9jYv8RKxkCSlI2+632CMaayFzbwf/+K1bF
UPpPUhIL+tbvDqw20Wbb425eybDbG/nzvTXK+XdtcLGUdjxZiN1Eq0ABmi2X+DNj
mSJ5alde2YkUGDkwofNFlXAaRQb0+ZUpQvntRPnZpQA+6Z4JQFR9G73NOELPRXsZ
cKJoyA6gQpkTDqNh3sBryPA6QZzbEO8pentuDY81Nislmpupc7JEAo41slHXIymw
qZ9BQ3Dn5zakcDUXpLIPkaemQcbJUfPKZy76vTB/m62I8fY2caCPcszG5IX4nLhU
Uh97malJmVmR8QSgKIPQNwhmst7f8WjxsWocVREwqnt7va7FHgc3usJIYpeVKX+c
tYalPKDSMkntGGzfgqAyYl9d6ubx970vcM1btDhOu/b06T95CKsV1rmOl8fgsWX4
9HCntVaJIlDleguZsGycJmAOAYd78+uUs26wXrAmgVpaLSItfPEa95lFjYTTQyb/
GbzBmy6tj6GVy7/3yRoBSGhMSkbwWPPxcSNUPq3OP6MgAjy+Kngodv0poC6+ApGO
5kqw0HPHMk3YH42KEf3TKp8Z3tXv83rnMwiYvi/kB8ujvSCaOcRele5b2NV9S7XT
9obFnp+u1mciDX8XyfDqF3zg+Suiq+QFWbU0mSARh5pw0EXHPJdLi1Bgo1w784qD
kR15I1fXv+LQvZg9I7RvxZvmGPZhcLoM/Ur3OfFp7em7Gk1z7eav3pvHvRkSBpcN
9jKtUdME2PWG8w6WemFDNVQFEtCZNm2j1NbX8sT+YAvg8fUvMSaac0+9lgXug43E
N++CJCzw8uxCOHQUUlIXtlKRjedigOGvP+KtLEEtagaRyXG8K3qAucc6rIztbu9d
nAFb8rYaR0aIKABj686DqlvEMZU0abjgVmhZey74+PuZ/d2SCdablNr4NGYDKWwr
xxWIIRURQRhUXGHwX6kMvbN592GE8TtEjiqlSgCfRrIaiYBRHi1Rk3xuOJZ25jNQ
EJZ/ioqyicWiN+M3+cqge4DZoramTg42jI+TBMUMDQlFiPruzR59Nr9eNU4m3Oi+
yWJgFP8AgLsDVHAzQ22EFDfNdz7J+jpWZ6C8PDcFwPZG+PfWb423R2jA1NZv+d64
ozuQ0j8cDQYQionX3xbIlUa2EEjX553VJwONJFEp7iTE+NxNwGZcGUYlsIAn96Nc
vhCEEFaBQPVUtAVkrlDfANX7li7u8MWqZL7ljwPaEmxE7lvxoDBaxdZFccX7KHVN
N9hKf11wHrDuQaVnZb506goiDtlZOBkbHf1D4NjSITHt8eM7SchGDkbeD8yBphCY
QE52IXvEr0t1rfoTWHR0eyUzs86AETfg7g7WEMoSnyCNbdL3nTjoFjYZFsEi3Jo4
OA6NNZldbxoeHvhZHZcNY/hCjwQWRoIEZr+Ecd8tZiKWPsT1hZoEH7Z4iiZiO6GE
fIfxxV6zMT4RJXOrYMLFX5gIsmx9jdpa95byElfCmkfIhbkslC+nEYohMVyILiJR
G9LX/VRh0iyRjvMpq0fruyQ+bWpLj3aLBnQx7+f1stlER4uAg4pZc6YxvttcL84b
EKoA97pn8LUGitn0fT871XQNzOxEj13i4QQE823N1o8M33FGfokteDWmFT+nNC2n
QZHVVAPbqgEfOCYlRqqfI1nBiMubAc8oVc2NOkdc/9n91q9CGAYkZC1VhMWsDwJR
Cajnng15Nrma7LhgS0Z0nDCNBNhAVVWOAD2mRwKydg8XEzIpv1ESoGkDccE7JtfQ
nvfNPBNRLEaDNdoP7Nh8Q+4t7MGklCAxWETOA61cuGOGTd+Uc9iQfqlyti5Ay2eJ
8+ImVSqFGsNTOp/bPILJ3lGnFWDWsGHi9J5wjhqnE6ZU00c4FowBRBD6w+JY2Y8X
4F2Y1o6vji/Ogq9UhYQ2rnrkiFq39ACQRx98jQ/0deH/TlvrLzRuBR4TJsLU06L4
Nopp6hDNMgZ0bhJkPSsyEWwU+ASQpXdFjVRy4UBQEKphI/gw2f4lZpy6tg/UxyRb
sWm0KILW9ZkxMv3jLLkodhrLLQCSrQXJVVpsPpD89c8sAucwIsKNxw9YYY8C5ezo
Or/GaBIxYuQcjSlS/wnObeQIiNbzXPuQ9cVK/j6yUPmwm3xxUCAzJxrMx+gIj3kf
JJeBFaF25sgjJocPPYnN5mD/g5vNx0TeJGcD8MWRG2eQIbSPY6tOzbpaTEjUQAVH
0KYIvq0jDm4UMEuqFiJ+tap1JsBIIQQL/XIoZ9E4m6jmKq4JegklwNp47FFOk+H1
pDWqd2shlujW8n6gl0QlKQH3H77HefJ6etwvN/mP83ml5LoTFXj9RRsRZLLX9gJd
OZuNEUiUF/lse7GZLoHtu4EEPq95X93i42/aQqCC5lzG/eizK2fVb2myXTvjHVqw
j92hqEzPL8T/JPVqT6MLb10QR6Z0eNQ+Fae7YyNQ2Yq5Uz8nZuWaFmAqt0qQrqxZ
rvAolvOAaESCLjgMrFSs2GGA5aFP8K98FJsloo1hK4Aa8vLBEhMtPVKogZ9wkSvw
IBzAAFl39fSAWpENSXtxKwcIiIM2KVUi/vIe0qoneRobec4nAvBc7KSMAfNw0but
xtqkMDbl51cYxiRkGGQPKGv0ogfkpdv0NlgDW2PfExl+ZGRD1QXh/vQylOI0OHBR
NaPPiHV1QinIOg8UgKKTcpmGUV0QfWe9RK75CwoGQvHwjP1qaZ1dEEqzjXmMt5UH
43Y1ApDW5CieaM424oGSYecDc2kUDEM6SziMLcarxzLin2gambfZi1nXWwjL8ocB
2/ccQC9XjDiYma6ZcjDAC6yz5ZGBeJAfI/SCSdpiJT/rCkrjuq8vNWqZgPZK82OT
OJMdH/haZVO1rcsyJRzYG+UExsXhAjtqoB2hQJEHEXRMa12W7HqgcBn+SvyHCbut
6QHcs4hSV+4VUbKRvv2gz90SNnqnINFcdXWJh0JVjk4GBgowELmJEKP/gs9KjZRs
a4EBj/ygF3XZ4r7gc97JgE/FyiEiGQVRax6fwvMR1OctxRc9/wD3iUiuTLDYrFb5
jQhN6xo7lSCIFvETF8CQfR/K1Ct+7RVglg/0RMHBh6N/Z0yX5BQthfhgW54prBPM
BKKvfvEHDIU62Ouwn595Rx+qh7df8D09Pb9Nz+48vD5i233E3fxexl11rFXCwxCw
L4AhiyYb3NO/P17Ib/7WxT8DZ/d6o9tCQT1LbeYQIb5f62Qbv6X2lLB+v2WIguFF
pp3LVpU/4Sm/z7EqZPmItQFsBnLjijGAy8EmK7vfCNQg1mccXp3K4rTlJNWtjieZ
4VsZOSlXAiJ7VLdYgklMa6WomVK5oItEVM2hnGtDfn0eGncr8C778ZWvHK3Plh2G
OAau16GwW5Rii9dhKbZ55KowAjiFbA//w9c8CZ4JcCRyLPRRkOPerL95mgkjTcxL
rSIuJUSQHGLeb7KrYFtiui0dagVG1i3Dakr23DiFnz7g3Jqa34g2oFWUNc+aQ6Fk
uldcqLt4zhRiyOtsdaYJ+cUS2R003movBtQZyymtxiCiRmXRg1uUplueQv6RgeQn
UCgYqMeIS2X5dPI/XxIyaAlqzfUtnz26ho/0JtWErXwYqL+dh9LczTCJrjEOV+g5
cf3y833FfdpY8bip3y75lu7l6nbJPk0kT7cPvcJrC+ZBgmCWWSh+6Qp9GhG/+Gs/
/QDXS7Zs0LmeoktRzFm3YpI/Ee1IakF4nrV7o0iZ8iQ2cKVoLheevnMOW1c5TUQW
KeLviLyCYfVEpQuOVDulWfa0x1YUfGiB42G11a+GF/56xzjDKmtA6MlN3UHK5ekX
wlLGG8Dl0ohD0rZ7v2kGk4kW64crvA9znN5yrXzD3jPq1w0gkAgN0InnZXVQsTM7
047CTzyCS7lc3WFL/VBedHC3nKtdPBXjLvWU684gZFF3Ql+2YJlyVxriBJkS4yKM
2uoZuC2k0mioFt95Uw7n5bkynbh5yMbOH/27Ng393orlsigdpVx3L3tSY51Vzfgi
D2e0liMu0/W+VwlzrXu/m2FRXxaZlGD4D8bpQG1mLO/2yWPDlGtnoPkoc6rtatbn
aJkzDXHhuOoKYM9EFt5dp84riwQnlInKFjqKPUQx8Vhwz+hx433USupHya4CuO0j
lINJiQQeHwc5nhk+O0PNQJrt28GgUAeS3YTirCSWYfAyuMw38PRi9FYJaWVQYLZy
Si1DFV5EmBsQvI47hNDzFALi/TPzpF8TmQRPiqVQ2A9WulOQs88j5ceyVT/tjR+g
rx1OWdbfrhgPxoLxMfrOuIKPB68FHD5C8I5WmnMn3hDAko3u3oCemWzDsEx1O91U
G3wBI4aoOth5QCyd5K1UOyaYB1bS2AcZiw9DHMC3QorE6+tbK95CegDhtk5fqteS
WguXZur6qoCQZy+TSzImpPJJg3gHGKWWY3a3u9SDIXcSqVJTsL1uNdQq8KqCpdJW
NxBXToxk2K6+URcZLw4f6rWYZ1YU1NX6QBbIpfThBfcIMpzm+jzaPQSJPDogpRiY
sCgAQ3Q9Kmv5RZfWZ6vKBUNyTqDcod5x+dyULYjJwG7ieVEcnbAAL5b8HcjSNpbE
aF4UVnAQdrPkCvXe3jEOiMOP+b6weVle7piyNDnUBqVHOWDWjMoN+WmqOrieLxGX
DRDHMedBINFgpCAImdEfgVwPl2sqbCA3ZixAcEIOGAsg+bu3hjAJg3hHss1tQi25
VSLMLa44F8NeHyQU/dGuf7x+Fc2zvDPHVqmIzfZUFAuJkQTwpPiGXeCm+aHt1xn5
hSh0UfcNat3AsPjuSrbzavHI2527uPPxcHyenYX2VKkmGKlEsmFI/3EcP8+NkhUF
5mhIpQbjWlLGDFZzmUSeADG6niGJ4aKquzK2wM3/SnirK5QH/pTxRXe/geEAPLq0
eMUho6GLhJN6RpRXyjioZj1+kxedSWEQE9V4FMgEbGuVxtC+kpkj6Z0ldhm41HGC
ryTEej5qSJzePEPweREr1Qqa6/DpGfmTz+qgbAGlIbvCLFUqHQZYoe26MlBl5JuL
a1ZJzjcigqaLQt6Kvwo9ZuimZXCxnW6RF360VGCtH1GtDidLhozdgkLjdQi/IVOa
Bpyd1ID3GsOr2d9T0zNe3Uy8VtruoLys4pN2ebG4/5zS7V+pRRoFNQ7tA97Pk1bN
A7lWDZT6BumlBJ2DtMD9OMJMaNVc2U93inJAPDdjeOT+grWcdVThCnYI0UarOlZd
aUXoWxvUlXQaGynqQ2e+4WJYvHzGQ8CdwOO+1iVVFW7XWnG7tdBZZ/awBu+Tk45F
hhAHRYETSsDV+UFYi/FTxoJ1UJDklEDtTWYi2Z4+ge23BQRvP4aY9kG+RCHpAuSb
qtPtD6KTh9Mmf4BaYZTDuURSl8Pgh7zynGbIIwg/D9RDzHobVj8etlQ4Wlrb+Btt
uPARdjBj7BZK111gifFFvJ0h3VIm+B3km7RG96NzWKii81UwIr7jETuNeBMTTA/J
5hYaXPbEBGMZqUUc3FeBYAuFj73SV3NmJYOeLwO/eZHFVnISatiqmoXO1sImGgSA
U5bMNGxxbb/O/STrh1vgDAWDEzv/EaZFWLQhDb7KMo2x+Q6+60fdX7p/2k98z6GZ
VqnECwgCwjz1OJ4B2IaQ5C0mYwech1eHgFMRrOIVd6IpXP9iaSvXogQgWJEE/NR3
Z91KGxINfDgrFbR82Neopiiw+SBqDnpn6UabsCq+P1bmJw2G5squr/N4IyPXULNK
QLLw3S8gAsil667lILzKCufbfuom0ooRW+DtMN8Tc8LXnMgWIaLlInrSCkVyVAK6
RNtajaitTSZiCYEqJNzUBZIjmtibwTF7QowY+V6UbC28O9AvFGsFNjt6d46HQQnF
CjwTB3nxy72+yrB8oMD5YMNq5BySd8ozBkEtEalaOqatFQsCyYcUAE/Yomlis9Na
zFKYslDfBUvVCrQEmlYwWeSFo3PQVewZfgxSz5vC7jab8Hrs/5b2P6szQ5izgPS+
NHoYEZlYTtIdBg7HMbHA4Uw9RNKxEEfgXq40iqc47mLZU89geECwucb7gLmjwvcr
RcRcpOp7XLAJiQiCVqm1jcXDmGz3g3oXJsE2xQCMLsw/QmyxQlm0DuTcXYOBLTA2
rUtCxT2ARhxPfRxBOTdDhTMBc1yk2aGc5cWbo8wLj3CPjiPljSKjLiKdyC4OhSmh
zsdLQD3sZEBM0/R4TRBbpXkpIONdkJzddsHjg9dJzyQV5XaOZUsIfguREMpuJpFU
c1C2HaUnwdypUSoGR/KodhjLPhywHXRlRcbABUzvY5AL8KvIDJuANUhXnchSQTNh
vPOgDIIfNc1Ki/Gi8qByYaUzcR1xJeT1/iugdiGC+xMr1ddyWTOp1ysbvtwloBGx
AC1ugBGOh38xUZTKsyPr9I/NKK97+VH46EUDGmMH5b9QEC5otLy0ImD8cUfLgY+n
GDxGu05kCVPuI4PhNgopbmUjYkWk4wNbyaFLDW5+rK86Ot7ska2NQA+5LN+aeF+G
zTpIHHJrQ7VeFCyucVjhuHq5TP/dgfwYgmGz6NNsu+XBW+bsJi2vgrSTukumkGgn
BfIfKoL6GcGEnIvrApO09fBtL/4k2tXJ6gYPlnXJzPXlEQS6tc7KAFbxtkLC9crb
Qm0Z3Lk8zWaDg+x4axt+51TcvsjsjhWSSNP2lkJvNwRSwyP+62i8x/EfQ8k2Ic62
BCMqrwkuYg3jCCDSf37Iy7enQ/OzQLP38a5uBGse4YGZ5qSdpF4Zd5VBIaq9Zm1n
0KB/sRRzyoICswhxP/ngNbbKHsEzLUdtjq6jMiY8YrVwJZ7U7ub09cRyu04XXna0
1cQ3Zv4BCd+GAAV1tamD0g7ri4uYK0yRVAiDtBw739pldnDtFxyd5gm+Nc01WyAx
V5E2NZSBnPw2oBrvAPO98ps/dBqpUKwSPAj2Qqvc5W3bT9WhFY9mbpS+6xBQK+6E
Xa0BgjIBEImYKrMCBzHGbVb80zCdvfud9ecAI0lAC1g1U2k2ujUVOUzxpHxc4pkV
NBQ3Kq8wT1iblporwJw433pR1sn27YqmdUkadWJR7EH4+FXIVk+JHPF8Sbv2VPT8
yEzhZCRxiqPttwmffeMv6dotu+LvOBlIm+4b/f8GzD5RJ7IIWKDzk63mGTuKwa4x
RDocpDIE52WnnoBznxjvgpWbu1SNKCKfIgCAJ4Xbzo4W/JgbV97g9mHRCVagHR/X
2oze+fFy8sShoU2VqSQExNSOpv87u3lBhr5Ujap2CrEwdotdw/mbDs5ASLCS70nS
4/h85aTwISrKbYhbAmVkpV3c6tjIE6vlZ9wOF+zJh5HA7QyZ9WNkfWlMIuUgemRA
B3ICCUb6A8nT6aIjUZvbWiY7vthOgAC0JI2ljH942ZbSvQq4NnWFeQLtH3GyAzCY
+drM/PMuc2Cuxfh2yBewUJRNrtAEfCl8i+elSEA18ZBcK54ffLiFcr0sOAXFUGBA
BADumHWgCw18rPHiJnJ/tEsWu8nM8bTDd9NtXgvQct7fMzQcAJSOw1rGvFxrKuBt
sFiqp6b3s6Usknav/6MIGhyHHKdChqCP7on9w6jrJtAzEbFD3wrKkssTIyrhk6pp
RBom7U/de1orRoyo/wDklSLyOJXN7P6BnPONmQ80BOW5z+v5zSv/feSHi5xCNZoQ
PXD0RrPAsQrTWcKgME7gUNEjycM8kA6JmUx+OefqEuLx73C4R1oIiYcGa0sgODX0
DrOwU+iRVAiQJpsfXOtWvO63217ZM4ndAGy5UgDWaNIAlXzMUdzlPNGUqH3T28vj
396mKw4vHykaa6CkFrxt13XKUtYzngFf+f1pn+KqEz8wtsTVyK4MTto0y4InYBTQ
gK/vMg+coTwhqQjBEWMWxFpiwFiKx1SMldxTlsx7xHmqMhbWhtEUMpebiwMzFftC
Y1XIExF3l/fsTCn+kxx+kouzWxBFwMYGTbVpU3GCOoF1a6lB679HeGIvlyB+SX6t
fHrrEcO5jhKsOYcrjW2g/M6ZZ9+9ZUb6Z2st7gRnX/02oEk/lgMdgSMmialFE03M
aCzIhKYK6uTX7i9kmV/9qLiHKKRJFoKXu1JSaUPAA9SMIxBV0J629ivhX9fNI4AR
AMHh9ljoUadEhHoQi0bEi5b8OyeVawOHxEc/SqdEcP2yyp1x6jZuCUdXf2k6uFnS
xsLc0ouTie0ob6Y2hLwxMBiXW+mE3ooH2xQ8ZdxFAJ+XnhUCDxObv06fphh/LqRC
8zHzXwgpU2UDwBkvPEwokDacdzVI4WAudIoyZsxXrLDIpzYFBgtuHNIarxsliEeQ
XrvFbSIOjyRlOMmxaKigsCiDR0ysBc24uo+ezO4ltsQ0lLLYxzIt4i914NdmoRoX
9ouDziIOfSu9hO/C1YOK3UiOtVLSpBI2tlr51zXycWvHA9JYuD2vmM1wcd3oUAkc
XQq320WRdU22jHzLTdb70D9Ii/Dkze6Ja7PlilgUqwBQU7TpCfuKkYqKROYAZCDE
ijUotO+bt3RmardpGcGpJshkVSb2C1IZ9EvAauCCzO2bza9KszjHhLZtMHq2EPMi
LzTWuIDsofqarI5c1/yky6hfeg+oUpZl9mi4KGwVvk3RMZO/7s9ceMSMVyrhW5gF
8tFEaxGgIjoxUZNrk6/ZNVOgIHml6UAyX2EZCuouP0LPJWhomlurSrXOiAGaG5Mu
TQZzw+2l7cBE2meiFxPJMursA25heWXjIth77VC5mf284fkLhq5tkM13JndNJAcc
/BqPBfoOf8Ue51OAengOD92bFFr9TyeI75MoRD93Jr7JvbRDUa8j+1ij3nSNtkvE
RJox0G89MErrnBUYXit4bqdVd4GPOGT0V8uAzRAWdln4QUaLl6i7g8uWN9UheNLe
7RpzWiqyo/hPUIoIYdhK1Y2exXSUpWA4+mT61cKKWZObcKGs4erQ08wGUsM8I0/Q
bKCgHZWihNT3JDBpDi5/l+iHCfzFj0xOjtW9V5QwE9j4zRlLGqZeNVl8lcqObr6u
+5DovreH7cqGIuIHOPIgEE76J171h8Lgtg+7M0mKM+5hwrfanQadbeFkgV6arV7i
tS5Lh/wzGJTYY/PZoPSn29yC5eFUt1h3yTN5S3rhGhP0cPQOopxsze652RG58I/x
AiLNWrpf3NFVDjd78Q0Rlyw93/fVMmUKGfUgmb9fuekWQ1J9CQxReqXvu9Yh3DkW
alD8TxEgdCIUCLR44441Ocwy2ji2hB5v6BIMY1uB3Z6kmJuidvyFVAwgQ7/rWUKm
q01qqIjD0ZJXjUdoTPqSsLTnkRZyETkx2GzpPR2Otzie/7ZpoLRdCZvAcFqP7igX
xqXhdxqmVio24x86OOrVqXrzIUekxStZk8lDpjtBMzAvqqeUY60GY3D+Uv7xDIM4
sGLOseHH+jUh4nGcxmh5MrBcubGfkOmSE0DU9TwXmvFNjsKxaVthdLFBxIrjZOTa
9EcYV5vAo1XTn2mdBUPoCIIXYp6uNfC/S+7XG83zCMrwrh0ngRhkIMVPD4WzuYyq
wW2O31qB1UIJ9A7fQ5wUtn5Z7XawqIMEtahmM8BIu+hGafcn8af+ShzlXPg2ISWU
VgnB3bCPrgnHo39ES4foTWQE+cMnfWS1XRaaHyRBDtDjzRPuXIn5+ytO3Ah83Ztl
xLnFuvqQYsXDxziAAtWx2FoQ7cz1JiN6o6TlITMycTkypM1Xk8h0BpCpT+LAF+L0
jWeINBoAY5Ha4ErHod9n9ddTRbMHN2X8e18z+Va1uCut5xrJWDzE6pQSjMrVTs4t
VwhHQYxvd+bAjdenFRcwgY6BcRngX5DIGSef5SsFikJhFsB+ISoKwPCYZknZL9AB
CrhyfaPzhxNX5M/UfTI2UZBonDe4w5DvRFp5UjV2lUaF6E7TjADaaMyjtqYx1TUw
DVwavbqoaczVa2HwDS9m4xv9m7dGK4OzXke7ENz/cLwdwvqXgLvEid3G6YB2ivxN
V5QikXWANn7+WuKrcgsfvy/Ydy2yFeLHEh6xGFNi8URc8bgYD5eyasp1NArLcc6o
H9VRSjepYCIRekeMX0u8kaUGMwbZKhQhtEHpYBml3ZPEYYG3FfUpDMcsNsRpK0D0
pkSPUIFX5IIHIdDmFQKJg1P/0OA1VTZf3d41QlulUd4pN/JbdPPygxwJ60ptkWij
b2CkLmAFDLMflpf9M1sJSAQLIA4yNHEyrcQASecWgozD9iRv2MF6eHE2KOZcrJkj
EflVT0OTMmqfTXOb5FA2tWKHvULbw/ew0gCUhbcosUIj8Pllb+13bFyW5CU3chMh
dAXysOF91F0t701m5nozg5AGORtx4/LqeGxdQwy+JtSp8Tz12frNgtRzRu/jdtZF
lg/WpYV+r/Gf173dYFSm0KFk+DAe0IQMuRmnDH4UHGyiFclrnbVOUluZ4K2nkYkL
itXndjGrcAJh42PhPUfwOQ8Cg8ptrrJhrbEmCLFFRsNzQeFV4Fw6G/vFGrVBlH6M
s0QvZtBtBbfSymMrLbdJhaWV1fguyz6D/udFCE+bB/w287DY8C/IAhZXE6/mLHV1
KE/smiNFobzkv1QWJL8ZE4J5LQ8g0IdQVearB7sAc/aFJ8+MoukhRJS8dtctSPOH
foNSsuJAyx4hmGEbGc4+f7hSbHcJuVeWIeW8e6RJpYWgx/ZkcbRaZAKFrSsLwB6L
QWvsCDartY5tJ00my+Af1InMEZOjqbZ09mBD2gtLUS7b552M7ZFaG1tVVeXwNEkh
kJKtKSb975yR0AmB07F8FNkVMDuP3bfVXCuuvzxXOvYmMF7slCAIgQ1kVIJJ7Gi3
5X1XIqP5gie+kBw2PXhSYmvT6QWe53b0kfgOv2ddnRRg+GAN0zAUgL0PrAO/fAGX
vrzHXkQv7LVhDQdMd1e5FD/R3A1Vriw4FMxff9iWMZpVYka8e/0DYmLcDPmjnWkk
+mzWjiAbBcOmDZtt3guNVG9tZIW0Del9YT4MpjrcgMlbMUzWWR7c1pKTHyB4kowC
i6dT5wbOoKd2x37aGgG3whXKGXfCHByD/j9eEjb0J5egPVfBkTRFzhNCJ0miw9qY
tjaUwbVfI0VGENYicXzvSE2StfjN1qv3iTPTDZaAsjTFN8ZlWTltr9T4hwgOMM9Z
s3a97SN4ue59oJgMhNkArvYuzoCRX6vl5XEH/pRqbNq0/PDEeyt989nytNzpSYuK
ECzjaPY1lOTFIHDkd4ZOQVqKHQvF0WZEMHsCl9dp2o+4Do6yl+nmAfOUwP4mV2g3
IMCgbvxAUTRGIN/K4MEsYuqQ6WxB9KV/jN29Lg1tLwQlXuZWOooM4hOwQaKblD0h
3dMR5uA9EoHh59g3MWkhhFUcLMmGjuPC+ymE9P6feF2GR6PpJrEOc4sxQKH/i/Da
kA3NKRjsygPx7EZ8NND7vBQ/iGsImbgnL3MnkwuW55wWcGbXcd960QhizXUlFUNv
EgdADSgqqRjbLkrzAt/SeJoyWu6jgON03Vy7ep73qCEPyepydXZaloRIkiNHq6Wl
Yia2jrpwUIr/+Lr5530wDx0z7orWQmK5/gvm8L3rji/PTGu152zRYB0PM9X67aax
+MiolCoO9yrkIqlU/kTotSdtHtw1KKMoP4cDer+r5AmRXzFOl721hBEM8Od0E8l3
q8SUEZkKmLl9+NJMFgLLITlifLf5Sz2eHrxvtOJEgJlUBRQukLH/LOUFJUkedANp
/X5S2NEFgiKN1yR3gE6n3nDlN34+vy5/yFrWB5lXvlO3FNZMBxxznuNGzuqE/MpC
jpoYPGjliSz7MlxxnDk2ZgJfy3wftJF3uraHGz6jFXoXN1F/69K2ddyIdIWjVfpt
4wqA3IWXYODZ7+miRVHKuo+UYbYCuoZMK0HQVARQvpjRVLJrHOYFY7urkHMBI9CK
uK2sZlLSbbT7WENBaw/7A7LJf+UhzkG7a5E9Dn3wqoasYDk+IoXXSCSX3peB52sT
oqQ80B5Qdv4fx3ZLabDDdUXk+M6afQW17RlDLp+Mjaj6mRB6dHrABVQVmBi+doAF
Fd99H8A8dAofwNUccx9hUm3qNiPozlsxk9+T5yKcfuUZfG6k0uy3m3uLWObcmlGd
dGQEapafmv+KS6FpWjqeqJaCkBQE08XOPBJGkVscnEg9wCM9TrBY2C42v25rt/F1
w735HZ2iHqldWH5yweGXDwbUkM/GobNLen7CeqJ9UB39o0HvkDNHsYWoLZWStv3c
k0EhAjY0cOQyJzwhzsm7qE0LR49aHZ6iL7WBXCoOrYdSk4BITIgFZjaopKEdQF87
zPaLEx4xY/NqmaQ9kO9mLJl7Y1wW/J1f3cfpHEvp2IkDCr2CXuo9vtiBCOxSHO32
PRu6U6gmUYihCtGni1pUnzrST59wsVMnYXBOV3S3QKhxCrx4w4ZEl6/GpFB2vga4
f0FP+aev4I7wE4F1QP5O2rkqaaQyjF00l7gf0eoG5tc8raAlXuimGTrReMAVFN2i
SmWAAW12gS8/J9QJ70949vJb8lavTcJNoWkoEWW+njIS3ipKu7TU9HWazPuHK3N+
7AfoBTrGM25KT9vnB9KRYhN9P0iOBeNYbyIdVMVtC5CbBrsUuCOlCDLdmhg1AKE6
7AAcK5qnOPgvv//zuD80l0KsBWtTyyLT9K4j+fkr8/8rDuXhxtwwMATx5/4zHuys
KGeyX73AcO3UldK3iRQIX0hz8+oigLsT3GcvMD/prcv31TkDMdKhxeyQgpUxUyIH
6VWEh65Q0LTjuFwDLFwuFNN/qjnNQLXOwqJDolSt5CVJPepaItxviNBShdvxXypu
lQrGOBGV8PRWhBNMr/wU7QXc5Z0EEKHtRPBbiF1ZEOqW8wYO+tvf2LjCQaHX3ntj
oHd6CNNkRm8biUsEG4Nq+POeLLpdrIsRXWewM69Bu0cF4az/Sap+PLQwV/9Qtu+q
Ye3hGVO010JRoYoxsi7z8G/xNpanI4Fbq67t4ok87vtQDisHxXIer8i3i0piJO+0
umTGlmDtBg20Xcp9mS0pLmb2bqN/WOWvdDemTZP8OTxEQKUy4YggEe9F9C//WVzK
WIjOgP1IygNkPO/YQH+IDBqXJl+Ppm60kZlQ0Z7rWHDp3YNUaZN+FOmraaZHXrJL
mN0r2AJVNfIerGVn8yHKwrm8LargjaACgpED+OH78n5/e1bqWP0W0jNrmm737uLP
C+C4u+vqKvrfYY5CEKrvRrf7aotPDYRKcLb7kR3u1wgskt5RysjGGyXRMQ1JIvrB
wuWPpw1MK3HTWNoXuO0Dap/HeV1R9mvsuRdkXldivqUkdB8nQNewFCKV5NGLxWGp
R/GXbB0KsB7RveQhpM+CBjwNU4weDg04+jjG9DM4WGlaHAJsh9nXefpj4g/AdGOQ
4jae3xL3j2fcBdWZtyhHGbOQN5/SEsfFKm9/5qZkdZ8QfV3vvrUZX0qqcK1w6Nki
DWSinAIBgNKK3HET3Pc/Tcx7MFAVLlFLMcZo/Eg8QkrLoJsuVD6BfGqoJdan+GlM
MdZihVZ2Chkrb+qRAn8gf7KsmOqDmKY3bRe1zzxlUbJEtY03nlBLhicN10LgTCWF
y5ZDyC6pQGeuxic6gUvVEA==
`protect END_PROTECTED