-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
LzkezjcPL7JoE3cvOODSyRn6LDaWfl+RhHeX/qov9Ac5JOxg6eii54F7ho7dHgsd
8dqw9aBDIqH3OlgQnTyrq2b/1/pU9zG3SfkrqXo4dHk34/EzqCmlbAfTway779Ut
HmX+auuPHWkTI/A8MGlYkIGUdqiJ5L27tirjREMEFVo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24384)
`protect data_block
rre7b/vynPZh3gtfaf1u4HEwUpUg2h7rrcL0i1GhpD39b+PXkO1l2oihx0klfvUK
fJAYuKsIzpP1wsOnkKvE44K6HeDvm8oaKQz2s39zKFoVLqmpzt05TsvuRPZsSlyw
NohyGtGn/WVbRl8FGsVwrRLDEdpt3/FuEs2z87EfhQ5FUXunmwrBvFjXWm3Az7Il
7UfS0eyUwD4aQsq4fAKTFhyJIqhqKdfToFlgV7dUdebvDgoeopTlt4ExAfFGVeTM
VlelG+u1luCJMXuZ9dX9IKnTD4gSHpFp0IeQgoeMBUDHX00UJqnbarW7VrPGosII
Dj6yDGin47Fnfk9q8zv3cSJE/H9Jdzd0bBIev2tfTNYvx5fsylViPij9H8gP+6tS
+mcqRCTYUnUXU616q6K4giEr7cWjsIkzm8C/C6n8r2QeksImlhx8zVtBZlxU+BGn
GOoQFUgNp3bwuQJiUx5dts1hbK1C0Zj+DrMYGe3eooR7Wg5vXijzhNeh+vVFfbxG
iwXYkdYgm57t77Qz3CsMl4lDKM29W7t0HcadWzU36ErX5+Q3lDRbQdKMwEV6DqZ2
qSS7Q6w1kwsbIdfAteoE620p+1nvZlRrsnpf3ZI3gom0GAOHXqpGLdaUoublIiCE
2z1JenxfRDnpkC+3/vi68mrWNomdmySOWPdA6Uw2h55J5WyubDBDF2mSj+43gh2n
/AIv/3tOslaXDs67J+7t4vEwZnBngs5B/f6+BEkIdXMPBDexCKTVotoGcdtdK5Dw
GFu3w2XJ8OybyMlTjblPRYEn86OVTFzKREzdR44767f3l3Qif1FdUp76I0bcE4za
zw5If+Y0s93h8Tv30c2GZETdEtt71pWPQBk9tsABAbtbfauUJ/oHRQzba5ArR8Oq
B3YoanpfDMzosHVoGxBEdC3L888+7Fjs75veBw3fzchwZjPOPrAcFmkv9Pl0Cqtv
SFw1meqNrQLknyTyxiDldah97pm0JCpbhz8eMInxk1VqFLP3PxlAiM1cOZpgGuiD
FD2ZmpjDh5mjQs7sYWurY0s5HiQeFgO0yUbw6sE564HW4Dte5gksHxIG3BzAd189
V3NjsyCMz5J1R1jsRzaeXT3Bq1W6m0jQvimB18HB+a7rI/Dfijl6z3r4CSe5bANp
bgY9w/Jz3F7Qe44T653p6rFedit1K8gZo7W/6AqBcY347wnjVBZyubzQULAJ7m50
kXwNAFn5B/8zu3Be5ZwmkF7dxaL7bvi8of5ZD0ZsN6g2AyIxyOdQuCfVWd6/Nx8u
gp+/CsLunwyEc7lLXe3j1uE65IX91xncPoCSNZf/yRQps/EUjQtWecqidZk1ZNq1
LuMgeJNvVNjYGbpvLk4hZT+P3/DqgWey3uvlYZvUz+nz2MowcJb8/u+fkZBtIGOm
NP1Id+9aOat4cBu28sxXD7kOXgbPuMq96inqy92JnFIpsDHb2yogvPTkkqgHiu3F
Nw3xA+lyieedmWdjJLcEiMYjx8GozACh96toqPPO5t1mk86uLzIEO0JHVipLEjPL
G1Ui5vtN2AIL2JNfvfVrfN67zfSFeYU/KrLRzQRF8NC5c58WDWS2T+6o6Rw5aNxR
70HEGLfqcmi28frrSKzz76QKdN/UKhkWu03fDhU10hEHvBTcm35k1LryqWJXqO5z
ra+k8QKEs4HAemU2yo4r6nihUQdwQ2AseqPV1CYJqV9+IyJgLtI+96gPxC+JdDJY
2rV+faR93C4ClVQGO8pYtayNoF3q2W/Laxd020Z6smEzY8RJ9YiRJyB88ga/v9fr
qRo68gSGZdAoGmvRH655aInA6CR1InF9RVGHrxTZ60DwP93HYyAHgFk1uDLaDYfv
7iq+5xabvIj2S7aMChgzK+HO7ZLlo/Fwm7g+9IWQQRoyLybvLNSUJUFOwCLtqEou
PTcNTIp1QxbnbH9B/+/YsparH1S/+UzB1LqHjL6D5PZf+dClYnCsg39xDTu1NXNy
zwaF4wW2ko/lZNh5P9pC0axRUgM10i/jHEPw8tga/YDAjqTtcYKIE690b2KqDCB9
1QWSqlHxXOmJ3EPVjLsTYzMLNdjp2R8mhz/+0wxn6qb6q9o4s6qyFMgjKsoB7nXC
jjV1A9FDdm035+6X0G/CWG1AE047DjC2ktKGibDY+36C8BZqJZyi4+Qw6Gb5I+My
TbYihikueX2pZkJNVh8c05i6mMAlbb7Az4qJqPbAMweD212bKlxLst8f/gFM+O94
u9YiYwv1/i2bzasB9O6Kc1NiPNH3aHfctqySTJktA4giZ16Y9bw5oPSnJqoN4fMS
WCTu9v6vcTSNkoJ5xsJ1TiKZ2wlH0PCew/iBn1p1jXqW7E7uVRfJAANBz4U1X0Wb
jtVY3IH9RuZipt9TGzCXebMxYwn1V6WyzS/aNuBf3tf8HdxwOG80+OqEJd6WASvJ
RWoK4oRH701z4epLPhTv2Q0xO4YdfqpFVVj3YjRdmDKVWQJblTt92jKFSADoW9BX
2RDICvLlJAce+jdG77jMZ0DPe5L34il1PogN3Y2VeJwAt7+aOQdyFEpV606WLMUX
8uSSrbOWobbkST3568vIhx3zGEzvGg22I1rl/e4N+6VbgEnJ3/XXAMM2CCJnt//x
3S0khMXoKrjJR7M/wuTJa1vcpUgFeff7Qu+Ge7BQaftsQgV4io5LhOtbtnEtbw+j
z2NTqYftQR5bnYwO1BSz6uQBoKHVYZK8yJzbH7vGHyfWe6KJuBkZemB727TvCtDl
Wjmlh/mhhKvyuNwBoBbwMF+Laq6hMywGnMoYrBwNkJ4IKp2+9AWlTvBl5wSTq6Qf
9HPdDUxicQ76aAhUa3uFXjRysWq8kxmSmHtdqG8nH/ZTgNJPWeLLNS4Ig+76QxZ+
4xenWDzNVAveU33xWtPm48kEsvVbZTWdAuG8N+gQ5fa6DcmNKXCBgoDEvSGAnNyN
6pXRzDMkaLKbr5a7FXnwgvjx4aeeRNom/dWPp4wnxVVGSF22b39HsUnq6HtSIvxs
yfcCApVYxDKCorIYH3xKyzoUjIk7fyW8gHQjRfyDVGxp8Ho39jV1SwV57XPBdV1S
l8fAzqr/Fri0By6Q8ecbS5M4HRpYQHHPSnKwp0sWRHk/82ZA8a9nSAoE18HfDj6X
q81yzP0kELOaqaajM2iP3wPGphgZvvOV+B4jauEhjYOSmHaz4G8kfDm/iioMwxq2
7Xd8HBV0o22Cd9RIPDB/qsNcK7R+0X5OkIV2vWXq04MKWpTQ2yPOo5JgxneXhGdn
DQ9tVmFvKqNSZFHNqzbwTwP85a6G8gNP558GpbBhG15A1PcH9pOfnxi6WQA0wDQS
LLVWYkF9StIG94Zr+ObuW8b9j85yZUjYzzEz7WOuk/Txg7OiEdR7vXgItuhFSf2G
oNbWrxd73wFccg7at12LwtANgwuDHffmiMPnIrIvXtVHvemhOHG66yYXE/SUguB3
JvJuGouC+O/B9wcI1zPvvMPqWdoOpo+giSvTQNbP1ULr7FGCb789VqWEmeibqXmp
tv5yitYBNy7qm+PC2sXFIopzp4fRWO1fns3cuhrbR01u7RBMbwP0mPZeIKSkhKCI
SYz6F7/FRWCWNFjTxLavgWBG48gvO6TYgl4m8c3vE4bIK2saTVYKrPeQxvD3PjFy
pfWPXsFSmQCydHd9jt2KreSlRMYmkJAg8Mn3YshVfJ690p+QgJehHgSyr+07B0sH
WK0noLDonq1cNgwnXcJbHPIXQ9zNSj7kpArlevvIQY92W2LSNWSlUWODwa8ihp0G
H5rGoGGaYfOSG9qUxqd0s8tKa4Pbtk9LfgybXbzEyYQ0Vd8VDgbK1wnG2EtkK2Fg
q5y4m21rj6XFI6blZeNviTuQlHlJwyp/3d3o5yWEtvQv5mBOWFJMLKKnBynr6I3A
JzUrQ93N6sto9FhorQ+1/sy7NUf42J8/hLBXYy3+3LIA0mgPlKi8wY+9lsm/PfmF
6nqtn8WvoJ2VV27kbW789GA5nhFsPTFSACUPBumv8woORHdn0QTLsVj3n9B7rb9H
/xMnF2/I0qYwWT/2RwbHLfW+rQBhnmmqmQpO8xtl3HChsMjT8GdNXZLJIWZSwfvf
6pQwtGMWeIyTJlzkKGXR3aj3YLdgzn/vx8aQ2TBg8YYftxGKh/va2epvdCgJV1PC
eaIiyJ+LRc+9fzPgwVg0QtXXwq4PUuYKk7qrgqp+q1fan8xRZ2uWj8P8Fhm5ycXY
BdWC79nsn0C4aPSbgeJMAGOaNxaaJsVRnynlAqxZGpynFo/pKx9OVkeF8h9u/p0S
MuZuztJFXcEzA51uYMmJcnKL/PQXfkRHSaGptmrxQPC25CBkGUBuONe2rHcxTmPK
LAM+51N08FrZ50Vk5eY+7ZRjarqzc3nL9VgxGK8VzTbEx2/CHYDuIO+VKl52o5i7
LL65XPjIQHZpMXzA40KHQwqlvfR4Qfhx78Ayjo8TPVhn3MlnxEyvoWXY4WKC8DN2
2jSulXQ3nUvlZyMwfuQN1Pp07/NOp+pNnHD9SyhCfdYk1bVtfKfjQ0SjL6wa6tbC
HLEA5Sjr/iE5aCB60eAq1oSEGdWVKoW6GlBMcPEBdwjGmexFZU8lcEtgYEz5glOI
sfe9TVulEcrjFCx+PohGBfIz3rOszbzJDXOfdbTOzee2OihLXqecFT5KS/67VNaI
sAZtrlU6N8huTUyIkRWYvkbv8D5B17812892N6aYAM0FBwjgxxaUUvZ/9Oeuao8j
ZLSzYaiOph/NHsSY6XhIJSgWiS9eecbeGZgphI/5tMVhXfpgyJ9y0GrnQWgfct6s
OpInl1LSXZq9F1R9W+/9RU66olheyd3Vvv8H/vZfeyyP+OjUtGNTQhan6lHQuOFX
6JsQXFvqYUtynl+wsqGoYFBPDMqxLMe9i80EaKhAIVb15qOI12wncwGWgIZbPhBM
fPm+e6HehuyaO2A/5qfO/veK5apPS4ANXEDIh471jTSsIgHTdIj60+D0Z03gt6hi
jV7LLiTpz0m1sbHaDBEXfq/whVXqOaQ2ixLGO3kTzdnGr9kghAmtgTWioVwjdQlk
aZSCpJk29aU3PvdjMgX4HOAe2EpzocdjlWGgd4X70wB2CenhnDd2Kl1bYXFVdEne
ahjhASN6omw0F/me0NKhkDAMW9mrJBD+cJgW5uNGYnbiOsEQ6XJdaN7GxcXO9C72
TSa8Q4KkGS5EHutgjZX/WhN60d/IJOQwisZEEjOaLH66Ll2oA8ldKSwdfpM/OeYH
RPR9ctPPynYFywTyT7/h5jsmTu/HR0VjHjWvhIbVTpL7GDk9kw3Sv2GzYhMrSALX
vICtQEgkOeKCWdkCMP6iEti2YLdEwUhF+KDfLhO0l+dEnkaalWcscx/EaLx/JsAo
aCBPidYvQoYvgNJajzNFBBpv2Y9DegrWrrXG/bOpxGbkZ/La1WEnMtqXfNZ2L0n/
jkiM9Uz4Gct4fSKcMK3ThTeaiV5PZZT28htcQursDNx2BOqLB9DX2I3jkvNXHlI7
DwTMxsGF2ROKgSkiC7PBHjf9yPSX8YHl9h4jf4AlgGkzQajvewSmYZtyA6Yb8T3z
dknQElo/vy0p6QuSoXZp45Ct5X4MW2alqqylO2Lasg7qWWfMAX91zuaa4PjIehue
2m6rk+LgGYzd8RjAcD8CwMI8Qg/PFj0ph4LE9bSRpBVw8l2Uhi+wtt2t4Jln9EPo
GQeAtPTE6B69luuS/vGiBowNyIO+1QEwJmph6E9QoZU9ffbLMsoOzvclO4QWd0Tl
AEd/LQlI0B0u/1aSvcbsjJWlrgJA1as5wxxXWzhqnIV/ooLXREbE1fXIAhiqID8V
DOzGP1U7qc5dh7/6iizRO4gBIGghBBQ6n76DObZTyhERQvSlXEhF9qEzp/loon8S
lOvY1iHQf5D6BbJGFUglaS//5tdmXtrNK0ixjf3EuvAUisogJFJ42vTmUPk29Wad
8+NXomVim5sIBA8UNUXQftG9k0MmIOrqOiKONyxxYQTQJVU+uKIWr7baIX4lbZUG
YcTyst6v5iQPiSF+TRs0xZN/sJ2ImlfzuKtjOb+tBOUKeNyzvGFPv3Br6ecxNBzh
t/Eq5d/I1cKea+XVXMj3MZ1vd26Ajc0P/m6MXCEenF6ITi39lZqW+eREZjGaf/mL
YRbkEkvOKv6olTZcBqz99ueeRUQ4x1BzNkv0Lg3qlZVjsFAs4KB4jncZCW8V4Ckx
lSL8tdTi7NUeJkDMg2w1Z4MQ+TBbsUhNuT/2U3fvGmehY1cYWaZsVXBHnXopn1U1
xb27a0xUFVVDY4W7j+F/OCPDrok8QFRY9hjEnnB6RnfSqSbkAqGrieGJyvwS6pZP
GdG5UeMSh4HPt2CW2avZZe6WenIlxR6JYFBrxjD/eR8jphsdhTgFoFw6+V12G9Xo
/N/O9MUS8hKCc4FEjRP4IdIs+/qoeJjn8BDfOa/gYO6CUcPHOoPI7HN/+4KIgtnY
gc/qI1qpSnSBaA7Q1ld+9Sism2i6eSmGxW6PR9J/X/5H1kPtyVRNhiGZRwKfz+fi
LtDoStib7tY9nuvdH5uMTzk0e+7NoRGwS2klj1mUvG7lJpntUzFznrwyC+gad+SN
+xLmvBaIjEHkRiViiVG+YEK908ibaqSjsppNforCmYNlnsBeziXKUFUoBlFfn79Q
+toGUWm8X4eXyZ+6mpKpyvX+nkx0SiUAJuB3UZF+stgp7BR7n2K2f1sJnRdVxGLc
rkjac6HcjICguSE4mAGsP2/q/DDAuXnsrqZkJ2fna4XYzGzA56Wg3bozJqJ/8MFf
de/yd+OO8pstaeuFBjThZfdzeYdpRHZtdgdzd2H+XcVL6xfpOoxXQpNjhdJ2Ri9v
OawrqXf9FjtjDrgnU00UG52GzmZE28FD9RDxu++onOsynUljAawWysYl4zEYh3BZ
4ccCqgRXelRSf6ND7IXlPcYLmp6CyBkZJ8250UA11h7+lt14ncvQU1GJV7S8KEZn
OLXqXU+HeIFEG/WiCpGZBzaJnRdmcyY/rqWBY1fZy9S8UkMiC3xUbK/MKGugpflL
UeBnFmGu/OkYGVfvC5HiI9XJ65Vw+LZp//ftyOsZCD0+MelOBa49E6cxHGAurJW3
KtZFCa7/4cMA3/zLOfELtqHBgUryzZo5sPJlKopGRJsL8gwIxvfY5mvLllPHaUgl
OaZiGQiqa9Wxc17x3woDw0uC63RQj2XuKKVhWaJdH0ZRkxpYykSKUHy/Hj1j5/g1
ewC0x88L+xaeziSZy6y3V9WEA7PZTiVaax+7AgjxncaQM0ykxo/07D+Xv9IQqy+v
9AHj3W/vBaQnDT4COcaK4C3r2uV1MORVzDoF9IN/vG+zkUWdng5BkqOjMRAwRW3t
ffRxrkmWqANx7hBSh3duK9IHJ6CESz9EOE3M4lVtRlEOGIuJDM47bD6bVvz5zjZe
lE5hQqkx8EaIbVwf2ugSyF15rwi9eFcDysYNrLq+cDw7TjhsStsCB5fuvlxnZQml
bAnTqP3whoWUlJUX0dBhiga1ScT4fhuND+1afPHXoxIi+HSVIoWA9/8+pmHv2u4a
9StMB7sVCwQctBWpSBtRCIAiGi0hJ3grsDHL1prsOHuFhw2bTJVEoE1sMm32f7fN
uIJzenTqqQ1FGOnMX5ARAVcfzvwGw/Ogue9guIlC3RIPocKHaCLr3Etf20wtJAI7
diO+u9nw6wUm/8olk1QqS3oBMBuPAG9JAPGhtlCmsRPDFy5PZDNM44yj4G2Z91EH
Buu3ryHDy5I3HpTsVaNcmZKKkuMIpT26VdHaql3VO5tNk50XcdziMZhnvlnhSZwY
Pv3JWhc2EL0DW3aCNSYmvbcW89B2ahSgsGTyQEsgWfCKj8Xq3ILOAiy2NLuWElyK
XyABWnC6/WSjlMhvro++hExAzu2OR1H7gXDetYSOpUKqMahPH56g4ZofX2hIwAW5
cfzxGroYbhItLSSLyTqANvHAB5SSvtxD4lvMoKMfWz+Q2bMjjGN1v2arXy3PMrE6
WqERi30adsO+nYcIgEYAzPFulBKqucRFbvDi1MWkjBehIoJRHjKRGedXkzlcq2a6
/bji3EbS0Grfl/7U0DBVsP7vTJyqaPGNl9IVNUZdWqr3cuYuSCQFp5mqCXNRAYJU
jodUKakFWfkZsl5Eg507d9y7MghrF5SDHHOqsrUIRRGhrKIG9B2srMX1vl/XxYmK
7a8SQCIpienyQkdD7DWTGQSnCrYl61x81i+gm+xf5XbB6vT/LTw1xZRh5M7fvTP6
97pnXFWcgGBwfsoW+1Wvyu8VIizcdfzsUgM0fYgkOgoc1FIbX2NnVrKLTw/lOL/H
LHX55OOP/hHcPmUULci1gjuDM9iKvy3Qk+Q6SEbmyGVR/kXO4huPz596NfO4m18y
5wr0INh6K9VeCXdhGp/MyagFLDJyWmQQDIrK4OoezLhvx0q2vB/JBy233chAe/91
3aux0bAAO4hyyRHI5pN5HNr3eiM+thgsZWyQ/5xtennGqNUBJO5jTe5Pg1uZh7hj
c7mUqhR2H7iTRs2L/0kf8rz7KfF5h0iX+pQmplN9ngACv3MMLpGuJfCIz7BbOPNI
CRefwRo02nangvgxM+jMAHt6/mk1LH6dl1cywg0y67ZKjTNHKCaYijtUip+iT92T
vZbaMw+wRDxzQsU4ULji58rT79F5F9BWNzBzjsptuudj6z/Ecn6JHcCHtjpYl90r
3C4EKIXP8yIxdCLPP6Q+OkLrbnj2d1gQ+IePZViaghQ4l4DR62IJaj5oVwFMrPke
ekxLE5jPdPBv0VWkuZnMRzoYZhgRQlj0oSDP9a2uyoFN+Wjfo94wsw2WZx6vY5T0
VMDH8GDOZMavFh0vyiJKu2gj5/wNca+Uw2BPfFQPNbarvzu5YemN5utyCdIu0JVD
UtJ3mdgkjTNERImIDXnJF+rwMYRcSmNBOIXxRCKyLz+dDuwLCmMlMmYk3T4pA1X6
ltyGfXNNHVlgR/fl2vk0UyuruXG9Wxf8xrWOww43BReeRBJL3I1GvKYjlOrYUoEw
TOjrnv8PaqYoOd8fZ6fghrL7W6QWECdzsFx2GwzYkISqoCXAxX4AsldmIT79FgNL
rtNlchJkjdEhrPo2hTe//3ih672GZqFEy6fVvh9GQsMSrh76wFs5Ij2kmhg9G/D0
yVQ2STRzsXkXgMaF4LezDcurplQ5VujYf1PJ0vrTk0799rc0QS9o6pkoHAmSxT2Z
U5pbn3YdKhum4v3/Pv/fpG2f4u3sA6Jy9E/7m5g0BXFep5ioc3p+dlbm9okOZNcg
BvY8T4U/y7+AFNeX8QC3cW+1ytfBl4DH6Cgt64uWZ6EY3Y8bW9ct6PDJXs9JePhj
H7LiY8jzHTHlJeMj6OgnMb8difUG0FgQ3L39WchJVcOcxpNqPOxY3ngco27b1IXQ
RaSmFcSa5L7l118mEnA0ppFUMQJjVL0SFZvvM3seJFfaTH5ZMg7LYYfggwqfi9np
H+yk9L2J6JUUquwWrHouIOJdtE2xIuJDIW2iHmxVylX19ku8Gofnv94rVsRTBl7T
i0aeB06ywP6WlZsj5u4pSObW2dJkXS2B+PLv+nD1yg/AmwBbVlmDZImcfY7ODGoN
pvK/VDY9j+e2JD7qLZ9Bya6RvylF3mBvu+PbcK7fugxfGmrxyLxDv3cowGBfRhTP
HfsgbV6Bx8k5UqS1JnfID3PV755sA11CY6Ugwm4m2u4aENA3uUM0xzhCwpwd52/v
6LfxsK3EDUOdUR+c8qbFhvO5TcSS5DxEDS14UxLqlCr/eGmj5A6Yu06FUgiieCED
tpNu8xDaEFeT8oo0KrPMCU2odeoGtf63HqRCZV95xImQ5thsUf6noYgAPoyLX4qH
tQ+Hr0BvCubQOjAEOxK0TfKJl5KxFNf3i90QJWVxb17nJynNT5Xd2LYXXoWXrn0x
nEE/SU9oSSnxT+6jbeTQ0ZTCcuBLrCvBsDTzTF98r248fbDQlu8b1+r7A/uAfJK0
ZbN2SZwqp3milEJaRKb+vUu5VSLMZTph4D38TItkpCLvbMQTv/ynj5umlqY5qes5
aiyo3Jtnnegzx54UgXqdRhYsDGi3jTA+RmWMCQ1P5CD0w1jipxkyLexZgvUsb1DS
4p6nTfMexE3umRWLD2G4Zl0d8ZGKrerjzTcR7RTx1o0qXWnEkrY12PNSUDmnKEh1
T+R3bxVmOOAcMEUW1dF0MxYu7wzK/enk4aEt15aX+XJIQsj5W9zO2tAZzEsh53i2
gWAeEn2o8vjM88D/OIGKTDVK3FH4b9exDvXg1zbD4hLUr/oJGXmwKbPEfKUOY6ho
5sfJd0vEbImyF1MyVzlTVusP1S+m5Q5/1BfklNKHGdggrcG8GTNUSJPGrgVnljI/
TWDfsLMKZ+iO13yB7ML+I3WNiPZoHCuBTeyybkdl2ogvn3uqqCfTWuTslZwp0IsN
u580vyse2XydSgER9bcMkIQBlfwilJJpBo/Nvgd1RXqoK1YNBT/nbiDcSkKb4PQL
ISczNT64aFBAp/irMEyUl8TZ/VWxC3peMLaV83PfvxOH8eEFUI2N2fSWP3eVatXZ
UXlHJn9RhVymUmELmrgCBMzpK53q0FHBJxissibSw6byOtdaT/P5WkIBLtxDBGYG
3DvaGCNMiLuoCKQNWRpnqaO6dT3hSCsod1xx2Bg+yrFxJFgrs+ZPRdMVRTalAn8o
0XxKhxhv+xyQvK4zpmBitEQPUvatGow+1RnlPcXs201sW9vgy5BpT6H9KM+eJhlQ
nLZH67XSpYlLaJJ3OWkjC8ch3AeSKlxuVEHFANQj8Jr2jJSoQ2JS8X1zu7CisQ2o
JhUmj3bhpPQH4bd5IrhB8a6dcMUlWjiHysdYxP89ueNql+dp5BODuNdkI29l/bFb
ywrG9PzVhXi3AeKnigj+mutUZbd0k+p6WiXrGohtN4HR5CtEeeqcNYrIPaFGsm5B
M4EZJCkRzKEsK2fjk+jKCNZe90+6hQsWe7ZbFz2FleQqYtKQ7zXUHGr/dVYjubhp
w4qY7XPHGTR0G/oCMQXW/8P8ZTelFxftAfFB2wpXQ/+g/z4MIyzXYQfJZ3tRxrmH
hHyblDe9Il3lPhUP8O/9jaC5XFqOO7FEue9tDiPubsMdhm93rqlOyOVX6AQWfUql
1wqEPmtG8a3Gc5ZztPhjGSRwlrYsOuMG2VMeUaA3EdCJdDjkZf0max4zwGZXn0TS
D+5ZYHAGYVUunA4MHPr7e1oMMlr+NGceIrsGuoPU7rzeXXh8U35wQlBo+zwSJpcM
mVBEXYwAqrUWXWwHA/GVBz58JjqbcMP2NREYfQWUJkKytGDHf9VWJYCL0jNB4Qbl
1Q9iO5HpHjE4xYiQZTD0RpOnBVLPgjVlkfyj1zJFhWyV/GMbk4KLzRIT0HKpKMlZ
BhXFLKDUtLuRoc2/xoncQlk4Q+YngEELNmhUg+8ANCkL17jyKB52v/jph0bOJM49
nZcd4kxmD24OUCHD3iZ+9NcYLtdST9bpcsrQaPeaKctmFKlqbTXQyg2Sk6SW+abj
lsl7QLLxLzxV4MksZPexjlZQP8OFQOVdI+m8NVCtUtdLjsou7OPWPIVkOYCWTEFm
zLb4J3u4DQA+vnWODohxIKO2hHEM43GkCxfzwhNbJPhEnnzhz+ZwYYELAunO3c8t
2cIJaIwaF6pC0p/kDbrZ1WqJ8/qrZ0Wdg32h49tBCr8cZNGjZ1bCSrYg2jreOmQ7
Xql8su+oXNxNF8FV/Vja47Im9n0vxripH72KSsHu81JPQLgvFzaNaKu4pZ8kxSyw
GOd13th9vlo7c166CNPX02q1JPQOrLFOEIQKeiobmWVaptUKhyvkVrqX1BXFWoza
f03QCyPqCSQGZ2fKEdcFGnoZQ/XFp73LgkNuVi4a4w+/JdV/qetKQIdkwJVAJMS4
9e2FitrscAwlrcfP1tbkxWvUF3FfAVVTeHDxztPLPxABotw22e0Yq/hSDb08scIm
ZZbdN9iiS3VP/ZFbHxEYkEbrnzdP25OwNvNvSPQAVSA6fJyGzt6hy0E+nwD/0lEM
mFcVFeydHTeoou5zKq7f4nRWV3Tnt63FcwlFlo/LjwwHm8YsbXT2adM/sbXG+nvh
0Bc4lYNzIlqCVRqr686FY92GZ4OOApVM6nRGZWWdr+51H5CdYEKMExvcvDpBgP9v
/uob21bbijEe6AlMgmAjlP1svVMcicsn82Fw8fqvRKpmrkil3CVHfp9RtuiVquu5
Ozmq/+Xf8LqyOMkx2gak+QiIn6SE0il0nyBEREDQVix0wzNkV/3smoyUT3DKeliJ
aEaacRIuMYbyKW1nnV4U9FSEZ76NAivmmGvmWHV3u605rVg8b2MQ+nLEQKptgTJE
wFc6AMF/2ichgEv1j9etQ9swno6fveRKsKzwbsUE+iIduK5/nrSlAXRfjyC2ekxe
VvITjSarnslpVT2DIW5Vc/y1vbWR08DDEvZbIwj93b+AebS0O2a3eTdIUnGcL8lR
LRa+wsF6IuIRYQXbFfOTuZNvvUu58PdfEzUBQl1t5DxZe2uk14Q7nkvaBzUMQhYg
6hkZ/YUecs1mJIO4aI2frTrZ1vkyuoNKwRkiLIgvj0MfHiRbrriGKt9ianwPbnBh
ie7u28VGkeAod55QItCgGIvKlRrNTEDSlBcFSfQctaKYLRVZN8PxPrfcdN56ijOJ
FhIE1HfLwTqe44ZloUUzpna+8wO2hvfe0AQnRI8IMNLLIPleRD7Q+HAF4GAWWFql
0rVDItMsQ03aZ0vj0vWoCSbNSLc/YTPVmZSdZCoqP79XIe5RFh5v1ArwxLLnmtH8
wDEBHCTao38+1nvubUmMK/yc1/rUgoNpap9xEjJMEoDyrZ3IMD/pW+3LZ9gdp6HE
uE0jHQqbtnjU7u5au8vSWOZt/g0pC8tObyVwi6JTGS2oUTwhAUjvqOA71cfOddk0
2xlgUZuXsK5hOSJwbnMgQb7OrRRd6b4hNkqkEBd72MCsOd0G8ovl2d3ahCuRU+NT
5KEu7nwoawnQ1S6/c4sfVKSavSG86K2p0Z5YZKC7mZY/aCtxzIItnRnZxFyCXeFa
Ayzq9lHWWvvKz0Y69V8Xwd/5XSmXytNNrvroFWpZ6LfHJMlLveeOkrcQyvPRtcQo
HruAO5VDw9Aljgso4kGo9e3K+XGHp7+2BU115BoORab8WzUspRW6a91gJQZLnB9N
diw1bfXR7iYAcJ4EH/g1dBzEk7hvF7iXTLQTbfh2DQ+olParnyG1J5JI4E4VWZIb
39b9TUqJgmIe7hfTTkCZznhULk/i4EEINDWjhotFX0YLDoCOynN8XwD9ROFEOTKe
TRpS8RwqOjT5OF7/YBrqpK7m7DEAsdzSEDCRrJWHk7Fbc49zO25KEle4M576ODVJ
XJsOM4rTLCx1xHo40m86BHpk9tT/nXXHtFgeTxFMwkWXAsWqSXFwp6s0raHlGKvU
eqA6n0htYUO9aLOuWzvQIAgZYcg1ika1hu57wYvC5+Du3eI5JSS/CnG1d/kGu0G8
IbYtTHZJXXJegZmjgkr8/lzNb5xUtcAEF4Ljlo0wmL18lyw47J31CMPZRAjbocrA
2ukWGkbVEps2TrIJ1cLO19MiJMPG+IPs2i5ABUnpjs7OWad05yCZ8Y9XggSVSO30
+NIXHkvFLpcGvoPVe5VEhekfy549LnaBDDJjAx6TzeWJEIq5LRC9m0IBpFthrf4c
uC/0zzrieTANxC9XstEml9TWBBqq9jG5+rrs8UthnSde+dzSA0JMOXcHfJb05OaE
dPrk9sJHmaUYeqaDKoJ19LMApsQOTsyUKzMBs4+nCSz8kEono8zW6V9++s0KC2aY
dfZ/NtGmD2Q8m6MFZrapyBdWK2IlrwgFP1NaWqeHBhtXxfo60TJvNAw3v37HDXGN
xRNzr31HKAgYyNkdG2UHVsWQYRK3iHpqu7sMy9LxcaLG8t6e4VuxbfbirGi3TAd+
k/Q5apPQ/y7wRHJuLovhCjW0cNOXSF9aSlq0SH5HzF8kzX4rRvhTv/nLpKxwr4dK
tDKTv42ssz6WmnIq6M2qkeyxSnH2GOuuB+ul1oTf+ijfXJJiRmrpaM4wE63ouuHa
0Sp+IYopj3b6s4DYCzIZEn5lumpnPZsNuePz9ZF4slzIh9SzPs8zoLcp3lwzztIU
KVlCG4rXmPzd+qY64NAa3fUN/wE5g+Hfwv9rGOfVc6M9piWOGk7HWxQeviqSFZ7b
hhCwLx/zi+FHnFGVz7FCLLG0P6AakSXvvliESe87By7eoQf/zcaju2tP3xxCscvg
MarlZEn+K9RbC6gaEuf58ZBInXDggBlp3saZWkrrlU92U6Kxq+H2KkM3lo4yCRZP
9I3l/1nPyhZ/2HyPZmBOliPT76D0ImzkkGMBo5A7jMw6m2I581JrAe9+tFS+y7uD
tFK+CkpwfWymdvWuUospDoIwlMdcWpD1ePSY9gd+ncwmezplEawpX+VOQRmlFigS
2qHIH5iSlb15kIhkp/h0lWRnzJmvpJT9RHJjrl0CYc9ExwSBmTL2ZQsibQpBZoy6
aziY5rlySB9Y4pk9WKEtLh5jQurRbKvfy7LyqWjELLs1o/8a0W6NLis6HSnk0q82
nr49Ys7K4/HJqiwLLG25jUG674lk4JGTWDqXBwKAM6fGgBoX595xfTOILtZI5ysP
gF2TPAKSFi7I2ikA9HT4KcrjoLArcBzFapg0c+7mvcjCfWCxwMdaEhYA4mJemWGy
JDtSKzwr7npN/xcxjV5QYBnHOTuRGeVFxdGNLhYlTw4HsAobmv6c3f6WGoXH2ejw
xileQG2t0kEdEB+4bkWY01l8dnJzNiu1ZrlSkfasU2GnorvqNuZMfi2pW9JTLx/O
9UDifzKrPO7d4oViUtpP7I5Owir/qSoO/AwLqJa2wxTex01GDL1L8bbH9tbBT8uB
4zV0H+frhi5D5uUXpwRv5isPqeqdLbwA3uVXtwSpTx1Hh3UMzo9+h//M5ARJcm46
kwcxzK0neX971yxreFGQLQO0NpPtYeDJVuBgzahHcT6e0pm1iE2u20qYVb86fx7K
ZiZ4EW62cIaCli3BD0oxUrVSofRWgM6AfWesMmWN48sJD9/aS5WTq62Y2hvq+xLJ
JlFMqoMMNkW4ahzU0ww20fJMVu3FIokMTFxF7+RTpIwNQVpFN/9Bzp4gKVw4PNOr
UsyZ+L/kWha1Ct56ooY4MYTzhDEN8rA+8AmkwXe5NwgbKMuRt/Puk3F7u9OrTubv
KuEY8j3PiwB4IEK4qr8p3w1TslnQugs3ZlC6Zdj0T0lJN9gsREloxzGUrXUYSgef
g1aHjnT+esvVGTppYURsGwri0ExKjiqdPQEgpjcaxvYOt3mC4B2iGQR0+8AJfal/
Av8019vUwMkaD1Su8Zg4nEJ8hNXfnZuyBL8MxnVpUCRz2IeGVgSLbcWdyoH1t+aH
5RJMJntK1z0X55FKdM6qOtQqJl51sTTGk6GcKZO9TiCrOUPEM6wuXd0rH+9FPSta
eM2a4dcEUx9X5xU2NLStoTKsgMDjH5ZXYpMf+wpqwTgf74DuQULnvEieLAnU9sjC
P2aD+djMIz6BrI+GMHr0WQQqlpC2xoFYS+9XAiK7jH8AkDEsVNWpRlTiJAdnu5A9
O+6MyGdV10ArfnUsC3cU4AweoXP/Dgdm9Ics+zBfZXFSoNg8cD43QIUH6+N6/gAS
3DbN3fS5tO1PaKIirvg3MSmv3vZcAjk4klif2hDrz2aW+/8o/+fBNOCcPR6Ijzi+
V4iJPabqq36FPrc/9M+tu7Fe9NFt2XeYHwo1fo64+o6QJKKY0ZMCI96WQSr31zM+
fnfNpWnEag/V+Q2FThu6yQ0tWUdfaPrIJIIIp1OZhzqBLbD0D2Uu15CN3EPj2aR3
Vy/ZdpnLAnghX5JYLl7LBSxDOcNYVtVlgloAXBtL9wPLBYm8Eiw0C6/O/FBMtxbz
KeyeAaJBkd5DlDYAOcyr2IezI7oEjJLTeFHJzWh+/km1x7nwj7mCCKo+R+RYHvgO
cAIBfeCJZ7fiCFAHK8giN/ot+b2KvMHJn6Vt0k1YnT4ZeOvDs00FHok6uKbqOtvQ
+5FzvoK8rhytXQ9OIcW8d3FUvYWTpn6SSNbpdHICSfGoWUno9952jG0nNQ3gUKmR
8AivgbnmAC8xKJQPsY5YikkSOCPXCFhx2k9eIo+rw0SC6v9Ojv93cIVIhyk39elW
k+9LcX6dV5k8+DhMocbgmBgPFCVtHRWM//ihx0JIy0nfNZLgJY60y467EEengXlU
DPWjxRI6LmxsdlCjBIEF2EzPGy1MkP2xjFe0C8BddNgk2qe1W3+aNPUn8XQxErQM
MRyrPTaUVyrrJWITKwwpgaXXHItE2hcP+NcPiDuwWwr5exx6tkIiUUi7feg/bII+
eq8FzWdORa+YozNNWc9EAj+r5kk1sQP9VpdUxhNOg//wxwsvPcf9JINkzI9BrC1p
FyoTIOelP2ains2TeixxuR5VQ9cINP0Ghdnp+iHFfHZJVNadntY1ncriRE2441mc
x9qJjATB6uWc2jHGK60WkdD8cWObNy54S+qYoBPjhoy0zGDwChS9FhGvj+kejrM5
SNB8OJyWvrmBHqswtKTOLOdUzmVM+F/R+tkpVijJKpvtYdtPuXq4kIGD7qgBBNxy
yAITF6bre+cZ7Z/SJ9XHSiQflTLzYzvC0RgY8VtGah0LhYrBNIpXoaLEHdZ9qOZu
aUJZE1SU4Ocq6NupvjrnFfwBfBmvvmsWfam4sTms/bEBwtGtqZPVojC4P4zrr36l
1FeVkrd2k3FG8jeytH7ecAh53LFRfgYQvBaJVTwnUwLt4Lvk5Dmuah6kBv3ldHML
+FOEg9fVG3G4jA8ojShzcbiQ6xRjETjzpYv+OapPjHeMGDOxpQTTxTfeuEPPOEc3
VoEYltTTIfpdLdgG4axKdYZMMm1pQ2BQFYerkMxa/F+k4uCLA18G7b6vmfUTAAqC
TiwAG1fFOLVXqvfkqBYlSpurMgwG5qGHjSNSYV+Apt5i5leyPDMqt4/XLieTlKSh
kNT5VUb4lwxMHrqfOMDcTQUcjCCgyvzf74pk4rrfpmBqQogmSa4focSqukuYxmaS
UO4yTFNSKD5yf5HNXtLkOcm7XUCAqtIHwlpdWvEHIIng6gEZAqIOGmaTBe/csTML
sQEcjbZH7Hsx4bAFWEbx/1Sm+P6phca9l+q6fpVTUqvwA49rr3nyhMK684zliSG9
HL8qthaJyNjX7c02A2/v80KLi/vVGvER7icsoJ8KVcDd8eNEvg7zoSrqm4Z04mr+
aEnZSiQ4mnPkij0zyIttJmw6uwzvpl1+00riO9GnIXx1mYhaSu4DMHWvG4B9U5EI
v4tDPAw6789mkwihHQiQKdnQvpxp39+Brlum9kRG/fgIQvXamJj0yyQ6jOs8eXeZ
/NgzEkkXDLMw6dANKqAwrkos2PwAAuZYJw+k1VKAFUd86uuAQcBhquIR3mwYc59R
pt30c/DGVjXgi/cvXd2akRm0v2guIpjd3bBPl6lFPoW8qXQkzDH+FzdtsisHylOi
DFEDNVo5OXUGvWYquLAQpOPymQVKqXlVB16U5CFfPMUseXXb8sXDAGebnG1kubAe
tMryxdBpmgU5wyM+tfvaV0gPVm6urt2VRZDTrlVRZA3LVS5I1EdUI2EQ6qhMr7Xp
SfyUMw1Q046EFAaGNfTcDLreZKaOOfLo+wagnadtOWz5XvBYRNv2RU31vAwsbiF7
zbEzQKQA6f6b+qRLGLwpR6uB8tw8rLgtaXUoscq0OfCENhaioig6G3UiIo+eCxmM
LxeVOcDp0s/FxAOxrdrxEnC3HFuAJl35536WIGD/A2Fk+XOiQB16aY3pIWm/YHuz
8IrCFkK3fjPpJ8aIHj7OQtgJfuaLRmXoYd7zgsGSpfgVanF3mksBOWg7xt7BTXJz
+wLQ2wLgef3FOJAR9vtF6czzZzNJwrArPiYVcZSK8JIkGKXFKycjRiZ/VPPAOeVP
s6bTwJwStvXblPCcE8VZCNVui8Gx6jn+l/wViZsT+4PIUK3TcIBx3UCMdtgSvmhz
rLqrgu6W1BCDW5+DXg6HTzJPFKRBDi4REUafdiVZGqrd9QZWfPweGj85SEr0FeUk
dj1YNdxKN9WdqByLy6Bvu4iTLo7WAeHBPf2M+fRwzZfi6+yYD4+qgl1f37t1LN5a
rG5frtTtOBFprG+t8BRwx9mwzXcSMniWpfAIM2MpdBZ3yNsXP2plZdy3uqeswMS6
Kny/pKD/X94SSPR1ir4ODMNuM6QzUiQDedNTFILdyzY2ooVbC2lL08Ukb9rdE/hv
qS9qUSs6SidGdaS8cuV+SG0w3vAz3ona7t4k4D5aTljvZwly0x9fOzd2rWKz8mft
GTFEm2HXZadNf0Stilkiwm92PIawztrlPE43VgO599HOAxDDhRWJTOr1R93pRIYt
/TuOY9XSx7pRs7Y60vOC//SPsfCkYgIxNIqyM2MTWtnUJ0kxdd7QHv87xYyBv4oQ
1+6GzJB+hViqVOTqLc0UEQiMQt0rz0lq8TmDJzl8/v2wJGXtE/qAEzGytLVfgKrt
6L2/l1sohs7q51tIg8j9zsTefWrHTMyXYpCdSnxEil9DYshFQNc/CSGVpsYhqXTG
1rqbNtc5RxoqzaJJjkPznegSHd5tXJ5b4ZdREmWfWnBQLykLVvpr25rA7YSDiZiY
jIgKPe3oB+OnBaNcIceOzbQXFjgwIMbUcQgoQSyJGYMaSSeZGJuMbYKbegPIEqcW
q6BXuHZXN5LtrnEN8NI//eFhwc8w67VuAlhKrztWJWIiA/RunsKmvsCR9GQedFnK
qUYho4VNI/cN3b7VkZc6tfbiJbpjd6jMBqhBBih1SjksRv6h6HxGhO0X/yfcpBwG
P0O70cG3wreEXirmXAq10oXy27WFfbGhx5hTydTTJgoSIo+UMD0buYPsimuH0h1B
n+eOxzJhZvsYOHZgA3K20Vk2SidTDKycSgv1KI5YKeOhI513oNtG+XAteTseHrR2
okLH7lWjZ631pTzXhuJqVYylF2Xj9X5vcC+1GHVfmtqDP62DGs2ZWDHaCC7qh94q
kCChxhEXenbwwrOrbFRKCLc+dJBbYZ8iZ9dreD/bTC7nkUx3nXOKj/suymCf9smy
KxPELy/AXsci7IXNgyW4ldornJROTLzeEaz3EnJFEdQ4OBxbpsnNh4qvSyJcp+tO
OyTEEwEHw8fPjAtcHip+gCMXBzNpysQk+3ex3/nRz/C/nK9W6n5wlkCsJrz8cEby
Pallx7EH57JIfL0MoSn3eNWvUdAO7KqEofOejRezKdWxpAEdSc0B0pmkDz3khfKh
ldbdv9rPVtiZyrQbSzE6h1pRWQfYkY3sUg8boHxn/xmYD4IUDgYJYsfCY1FC+WaU
LQAL0WFGtxQzPZgElogiVFQ9vkILd1hzUMKk1b7G5R708abBB+NJpCfg7TrKe4E/
hby7fpRn3mSQ5sG9qthkKTIGbeFJcuKuOyh1QIYPRbutKMhdLMbS33Rq+kWQLe8r
pViwPKMC6ls0BMzS9WJ1JuwalzeKMbQjSi0fLYkwKj+2mk4XRovQijc1yx6Adp0t
0KTP8TwyeVE+EtSlYCjHRzlTbVeuOyRVB7g2mz16NUgrv3ICKKPj5TtZHO8YmzTM
MsFutO/Cwkyjv+ThPbcFhhmWjYfEOflmYEvcddTqnabRY1jtVjWbXzZtegwY1dMF
eKpEptFNnaDnr+2/yxe4Ykvtwx+s6mm2UPzgmxI0GAbA3D/TI8KGxSQAUQf25qSu
v52afx/55y0hWQqW1V+559FUMG0UKAlDPWDxCx5el86GQneQVG4Gm/UDNcdd8m1q
xcX5nAFYrN7clwsHTZkLw6bIJCJjQOmEomQqyFp2qLfUNa/8OgN5WlqBrm3VnJPW
K/zfrKlTUDgEPwdmqpdw+lcakdDQ2dMQ4aA1KdOXBZ/hjrhPgajr4zj8KoGuQUeU
OarmtR55s/G6gY5lnBa4e9w3kiE+3NQp+5ug3JsXslffmKg8gYn5Rmz8UHnYTWaq
xk69jGBn3EhcGNGbAIulRAVve8GSgA/9StU3GZuLiGFwid9rnwY0oyMya5i2vEFE
tl3n5SZUdI+QxrPRRuv/a9gF2F10mZh744V4VPj1gMOLA10EOJTszmJknf09zDVo
p12b4abSaB0JViwvVlvjmdbTl8W/i5zWYBdqCyxnjDuRQxwNgOPYyuPK8MO23tFV
xQ+VxpNrNh088itw/5ZNs2EddFvUPwcwogErKPBj6O6sGUpjbi8brpD0FD2yfvCI
Yg9DX2w6pw+TM35rmQlNbiE1INyRG0uCWy6E3Fq0pGnKwDxRYCwMzA2+dkkms93L
PgLdp+D1MxuVF6it8MvNvmSjZcfAP4inncvEczmnnk94KvU3NfrCwmvWP9kbDN8g
m9BvJ0zI7ZwfXLZrL2zkC5Mb1tt/IunUeJaPtJL7MuVXpRJTjAGnau+1sbGst6tf
k5iTYFQo9M0qeOSU+dkLSwKiRLXUS+9IkWlynM14lYc9hGVW3mxspn8R75H4jxRV
yY9/bPd7ptSYE50GmYLHWbR5366T9SUXp6R569lEHqqO9TuykydylIJExCqnwlXN
SZd0zrvHWBDX/wEHGgV9r86p22CwQUMzOLDoM6clCb/okoLLxm0OdGKfVW3rUXws
D9qcLYfAs9AyoGVxBDBiQRtwLnxXMGbfLeZgDsKNJoXaPOqRkWO/qtAGxmvmMU38
vlSfI2h23hIweZB3xvPcnXq1jpt4ZVAvdqUbI+A4UVhP5WoUu86b2HJGfVS24DKL
JFJ+zbMl8FP+tVpSU6YoQoYN9/j9FvM0oSjpaSuAjY2rKpuFKCaGHYfL2JzXsXg3
uUppyZy6tx4X4V440LR4hX6Zp7lFd26YUN38hJU2oxuJ3sZrvCi4jXSrNzYqDY1E
F7Ld8ixYDn7ZJit3tYMrAueuLFDn6QwoTnXkNeUdSSBHmG2VbsE6T6Grg1YE7Qu/
1CUC36iH7QAIq4dWJztGB1TI8MjRiSkPseKGNzc8OnZGSQFHZXYwsJlaRfH1lFxZ
UC7sLDN6X3EvkWr1E3gOvknyadJ+/STWfYTeiWaQBfbqC6KtVhmRcanGH9EEEUHC
5l+2HLdRCdt6g2i/zLdyuybtxOjaT36EHClx5DrJhLSQBCT03JjM501KGqKryYs5
VIgIp28382UZPlisdNlHTJ6d03jqjYG6Wx6vLR7eQTNGh2WlrlI+8LWA7YyIs2IK
6xZR90ndYQXeG0F0jLOAfQeyKJ6llPJUWvifFNC+IWfVA0j+WNNrQu4Nw5u8uEdT
9zPqrJHsYX3Yr69cb15I5zNCcgMkJC9vPi3Nh7TONxR7Hw7tImbZnVn4LPIlY6XN
/aEPHFbo+cl2EGsVFRqMWvArP2N24YfPhzhKlL0I/IJyOHDsoP4ku1aQDzyyu4Gz
AgVUUUSU2VAFXEP8wwoqKcXsD55beqYJ8XFfHpgL9ahlLUvIWsDzDsuNsS+XLOq3
lXnsz29uHoyiAdF8smdPBAINfJXVgx3CpcXe18Hmz6VNTFGPz6hntIOI6kebBeoW
nQa23RyAT2g2DaFaiymp2F97rIiE5ggsMtRFQC0DL68rMYxypvuJRYVc4BbD0j2X
5jqqTHsyJYyoKcrLNZjT+ngXYBny2jO7XAGnRVkv5H+oafRM+iPPUxbxOUNtafje
MJB6kNER+2jEKAujm7dDhKGufOzAGmI5pqNQsaDXXq79ySkRy1W6gSS6Vc7o/F9X
FmXjvvMlJNwOv4ctpI/BcaywWMDquKBTLe4j0QxfRu42LE4f+wvB/i5XwgByqTHY
jEmXzmVyxQWnkuP94QeTrgv9PnP81CyUt7XdsIGfC0FZ33lGWRo9UHPd9ZYSodAZ
x4QtcAC7oi0oV27nB1WgtdPXk4Nowg7oNTwf63ba6Qb3quh9743+3wfQIz7yMDKG
TIt/NYfMT1ur3UKBa7wOpyyi5JM5LS1GzrMFxmrslE7h3hdCnvBLENj8pU7i4u3M
thAZL5LzMgNeG8M0k8hw7U2MfbN59aQxLDk06RTDIHxDCFgu5hlTEtHN9FX2I+sm
go27ceqXhOXeGSKGfCXnh6Qy3EM20hnT5Jy7+eT6qKAPwDs+WZrkwUQme3JFm+6c
RHzRaXvq3aIw++C8TlFqm20IdVj7Cin1vPULONm2rrFB8ooKZkrb4zk4x0sUQwx7
s6I3ekxBgZxW5haQrk4V82WZFvaxvKS7FajzraB6vuYha9MP5iQejjtrkibf4e+l
/9lLc0QhW/ewk1/TpyyBSlPwGB/txm9Vx+7mxSJlm9RrSGjUo0CWhbput6ZDHZwv
jqLpgQ2/E0ZJPyvX9s62RLQPtkLnJzmugQxH0fTKUfwCh5Tvb42iXwj4MPWkmdxZ
Nfwwo6iOkep5XNjlatP+cDm1+r2HEvxlR4sUirDNJABHtcRlP88huV5lmZBP20wC
0zrsjIBM5u9G+zdcwI/AW+C8A1MeX0nPHkg6kjmnG7Dq+VDjdh5bg7QR/ZPi0rfR
tlnI/v2+Jo9GZM3t+C9i/eXpWO92TJP2Guk/XeVWYYqtifC7K1eFX/pJHRzUWzr1
Bk6mVfD0VqFspEVfCqkSe/+lcFRFHesvMZ+e1TcW0RlrITs248mqBSzvQbQP5VMl
K9Rm+ijOoghEFAkKWxsKsFEVA+kuUdoMihxSDT4/8+3I7SsHLjdHZ+ua33NMZhL+
BkFRyFChoBg2Zc5lHPhXCG+6+X2VkA+SphnFUG04bOBpErD4cHIephaX6wYgRu3d
QCqvE4834+GmVTOOyEH+1XeROx6jbgwo4IfxqgN+y78Y6C89YeIGBzl9Y5q5rAVb
BOCfrsaBY3XdH/X8UCIbryEJd9KlN74N3eSQ2O+txQaFFFmWKdPns8t/zfAI6hrx
GB1KibNMdc3kEZIQn4aHX79C3XuJ+b6FV8JqyWOCeYjuvC5CJaP22oPEkhfFSrAk
RqlsFXTnXu25u/g7eVp/qPnTm0nVPfXYrakoJtUN39fYdBaMl48dzcBaJ31cvX69
z96XcHMAKHfe0EMTAM9how5/9xEN2Ip3q4iG/HE6oOK5jUbc7dlE4dwL4K9NVtLU
q2Yipxd2f4hsAQt2Nq2O7KQ2jopWaR1tGRLn631jJONMRZXztH6QYL1prjfxWefZ
ARhOb4sgm+96/h+FIzXnGqqcV8S6csj+6C3Wq0+lS6qbK27lT6IAmprT8Pf+l5Fp
7lifW3ma71e5/94NsCR86FJAJs5jt3ZC78jz6aVvSqf7eGitHLyqUUEqe1bYC5ST
50RvjLhda+f0eFsa+sX8R6ZLWLQiWmewKed/eXBxHRoP34Ml2+FZEArsqZeaAb3u
YwuUsxj7YJTJJ3sx6LEfgOuAgWu++Gacma2clPGv3Uu1APNFXTwuUG/5ffReC5RX
0YwLLfMg6/b46dWRv+dqJX+q+G1Q6mDCRBYQQoUn6vi47gXAGSP85YqE3J/uMXGU
qcHe57uJrSnwAj+xjMQKczCpdl9bpdeXHlw36x0iht+RCFJnNSBIGL9gKDxAt/yV
p1Xbf0wfytjphLBHqCefSDXxhEsUKRrFCN+VHu425t+094+L0Sf8TkUDElRVpVW3
8sniGUe+OmZXqPLjC9eSwUzuPAIB2iCIRGTPZ4ITaEGlFpdUVUkdHuGF42xhLOxr
GVoF9OgVkpk/dFU0/u97J0mu7qewcB2XOIjrK5O1lMdZ0fTU9Q6ldD973DCX5+2a
PRo6y+EuUwF+76gDXSqj8P52vgt/ML8eT6d74mAXC6gqPS4Inwy8ZrbWuaIKKiBr
byHg07HTvLcJEB7eXdTcyLgyD3QkG8jsMcU4PJt31ld3Tvho8vTAK2PfiS5BnuKh
ngrtDjn7PmQBk+61KG5MkWYp2kqYlknp3i/l69Tf7kacneD0f0yK3Wulr8JB4qBc
wGEreymDxoMZ8D885zVwj13A9a+coU2vmvDzz2rv/lzYAAcRlsDYRQB/iCTqVOWY
s+sz3P+b037UY01whWLp/Qw7ZqZ0M8+yrteDTF56Qyar4PlbnekwdwpzFbTX4H8I
eEBwPtSS5gF15P2ZUM1Ev6EW9ufXJA1XidbYkMObUvEUEKeYBZnb0NVirZF4LEEV
LaLYUC3QTMQK4Xk66SBxjaqs0IhomsOS5FXbnSZaYhNr8mZghwaF8nZbWqgBCzgn
OaYbNHDiMdFfi/S7wSt1r//SdONWJOUnORsbjJIPESrzCQUNmLH8IqaortND24p1
jeHIsbTvVibKHYeHfCHZ2jCVkj235s7m9xm94iMCszLSdMuDr4rDDl19YfnHY4i0
O0saVBVZeKr0mjQmdrtmHjQ7bz0t2ziZ6Nfg6vWtnUkZrjJEDYjXwzFo3CbkP8Xq
1F1v3sgnyIbyIW7X5x4X7WFEcuz+AotyWAfqq+AkU60FT/HAN5x48XdBU9xxnOYc
tn86FkBYMkhbLWH8wiY1BshBbNTMyTjCQi/g1aXsLwh7zeqoWjDhmLGZKwtISKjk
asUmhHksNYglBzd/YLIXBOO/OH8FAKrYd4G8TrT9xQgprPML+xRSW5YiOlxLvzJ3
xPtREOvtMgj2WZL4aeYxjB6RfdvU2LOMWdXktaLM9g0cTU1AgFGFI/qamR+9u122
SqFXX2ZNdHDN2PRj7NG5VhosPkR0mwF41gjK9BEBnm0Ob0dsT4j0jN2zUDO3LtgC
JrnCILZRXzJkupC5YE0/ElIe1+tvjM7UmsGeUDK6jSQ6GRwQdHTIRDshD9+GtL6L
1EXjTmbUs/CJyMaQFzt450M5wORl+Ys1Bqw2OPhtqKju2qE8w6TFxeqNKay1nYfA
H/ScqC77p0XwDJ0yYvB2OAMTCy3/kYkQqrpVxMtdKxyMK/Q67QFvw4118J6RaEWz
sVWPGMWIxFY4rdCqzBQ173dVA6RH/phGKv5PI9Kk7RGBjAh8L04LaLCs4/iltlMH
TiBoPGWQ5kGt2JkGhrekvYRh0IoTC2JkLNr8H/rCvPcOM7I0AI1z02kz9hfK0cAq
8BoavJIx1C0Zp3rh6y1MVVWZPJv2uHNsT+C6RXsgCVFTAy8IfzAwSfLTgDNAmSSJ
bxr/Ggh7eYwRUiClKVILqUUm5o5GaQtOgUlaZbtACyAumZXEsM+OG5WGaIEbkpSd
2tS5Pco0bITaz79fg9TU0Rvf9QeiHx3VBGgLKaqY8/nMqYi37VFZ8GFDrYLopiv5
48VMafHrdJFpjaAWjznz9KTpkcoC1bswO/JQeLHTCafAt5cwD6G8+24qDAurg3MF
4uYHwMex/4tApSXiH6HtilJylCWG/kIHWASJ3tCzudVIQQlefCOoHohGns+POneK
UOEPe/orPX5coG1V8ah6rjtjH42r8OYAJaX/CO6gBANA3lybmBNnoASkHoPE3pVn
1SGUBwcySpv7jFhn/BXXBvykYxcr+lqhIufLcnH0DVf7pwYe4+6WotVD5sMmxR82
5sQMk2Do9v/xCcIDFJa36W9+ds5mQd7BnBi+UksPmH0i3g5Iq37SXrFZXavzZ0dS
wJ2lbEO4/+5lgiIx7Ql/toORYFhSzkzuDY5uvLYptTUpFITF6icMA+M8f9vzOzIl
Ux+/NTrdelIp0MXlh9mBUoFONO3ciHFaag2zB7+mjn8RAi426bZzsFks/AOxEApo
fWA6kuHMCp6qGuZcZNf+rbfJd0ad+/a15rVLW9JSZ8OawTk61O9DqYWkiKxiSf1V
r8VyJW2hMPmi8FmsPYiygeg1+SwdyNH1GFDrE0lXuVkgsd90Vpqh8aEXcy17dOqt
PJ+qzwAFoXlXXOtaB/5hWzaVtzRh2jbEVOiDYpuCpwdjb3oxjxY3qBHfHH4tBQJy
m0QhqNQsP9VmflPFYRynRABHmmGPeLgMuPEmUXU20c6VxV8D5p+GPKswVTNkaRnO
tMsIYNeSpYVvyNn0fl1WHbj+bNrwrcwETiCW92zOPOHJoGfNNsG5uJCWzOSpKdKO
sWmwcpZPZS/UiPVYn3Uow1bLe6MGmGT7ul/plq0FrOIw6WwfRj62fUcWndkYfA+v
LQR+bL4Aumorj0Li1vrj5nQUZQY7RxmjOjTsAC3Ck2QJuQkuSgrv5b9QxfYMKhLV
5528w0aYhkirFC9TeA3ehsCVt7WK+YbG+ZUOlUc2/78YiKZftslZlk6INwNmXn66
mfh2pQG7BKlDUvvzrC4LX5w/JucAGry34DKNtgZyZm4HQY+TTxfkS0Qr4eVT9GWF
neXp+ZN5nWHGzYI7nJyk7aYcHKeMvHoS2ZSJ4ae0GWs6KqZ9sFR/rwAO8Ov412SV
bNiCBBtvLzEMtQdV9CmYmwROr8IyE0g7hiCcP7ng/Uc7a7HVO6pPGmxNz8pcsaPm
93UDOVlx0Dzm4kCxvQjdo+f9sjUW2AXj4UHn78Y8QHJXHbwmcd3TFgJx0LQZc72A
f+9iF2oHfOxZMgPQLeE8pWBgAgEQsBIb2swhhqdT1iZNQeuSCm0FzoTmPPurf5a9
JhmAMYf6gKa2tNk2fgVbTGUTQ//SheZcg7286/dP3CZkCHx4hi7WrxhyG5u+MwMc
dhefm+vd/s7ZcTf+G9cnnx77+3lb4Lpj4ewXh42qPnd5hxP1vT7hmqlsuMsug+8C
EWj1YEv2gYQ0dpNdPn2bNeak14jUsuUgM2hn+HsZH1p6qKWN6vqKDQvNZifTEudP
MF9whXyvejUrvskDh0oC79qiEzUnLucsyrmbu33ynhhmNqxVeRuzg9OId+v2OO08
5gIkuyANtRcsi7Jx7Lccur4JYVVYNof1vtElCU+zpC49mbrPiuHJVVsv2gyolQkl
LIhQrVMR4VlT2eyT4W8iIXPolaYotwlOT6jwqcPOPCxILzrnNjA/Vg3r5lm3R8Q6
39CYTYISa7Zryhp3auvJGPQPQUcWgC3SO//9vanTQAhN+4uwLo+4Qfq67RR7wbgs
AYRH9TfulCBnDWCopKJyYHcmidzQPtJ6r9OlFLPgM/jIScyOkMU1WdAKexPCVcQ9
DxdaizBxgGBwrqXGcdQDf5WcSpjI9HboghI/kFlmJcZhnNorswamdSIybrtrz/uK
TLN5fVtYvpsntiqfqH7Z+TRIHrl1xcKy9jxG4FU6Tdw2TPfpUoHUAGoGT/VPy/HU
lmRzTLbINrEaj59g7NHQivA8RIsfbmqAkgh6EDGl6RTSDFUD0Vs+aPnhw5pEsd0e
7d9kLmZy3HsDixxKTqFDRbsvAkTxr57fLlIlRN8JkgvaasqqcSWOI6N/Fo2V7+T/
i6h14dTVVUE3RXM+MkJkhlbbBpSWoim2KFFN/OeZT5UXlX6Hx+9rf5lj4NXPfge8
aHNkNx7+zFRxbC7k/jxhHmiiFuPaBMfB+WHvvVvo3WUIWYzFr177XoNpxi+0wxGA
MrBYOrIGohbgCCvdcjtmztqCEZHKsXHiOn2x2J0gdKdmmEGeHRYOUMs3GHxSrkIa
A07KgYerSNgGhuo6DVXYBUXBcR7Z9eUCU1ohU2QRPps4/srRYv5fktImn+VMnyVf
TpCTppQ9MeHqwkSdXVYPFh2xGidWQzcsD2ON9I/4ZvhvS7IfO5Ehm5mUwPUqW4CB
1IDjLuZ0rlQjmN8iLcja1aRLdVW8cX5I3Hf1divDE39SuPkg5uAkeedpxabKCyLc
Gbu1yBKDDN5lp72yoVDFE3DnXiND6zdk9Zw+5oeFJ6P5FRwyZKuveOr8NpXdgTRl
q+scePbmBm69IDu10IpGRE8RO4Iu3yjQdSfPrz3mdhEPslX5V5UZpYGcOS4fzbUM
iLhrlpf3gVZodPOGecBPnxgCOEDfZeqFmKSwwgk6xbuhpBuYhq9CwUEO/9R+VfEb
HfuldevGBvcltHGQQfg19bbglfegzo5SM6OsAq53Xsn9tx4/J9fskB+FTZeRzpu3
5xnxmgqAX45K6YsM4WEbux2rqdkgF/DbfasNSIgNKRB+74dlpfijmRkOTINkrn7f
+ny65OxN1wxip+e+KUkroJpv93wzMy/ZWqNi3XBHxM2kr6CNP06qogVYQZtgymBO
K0z2AVUhUktG+iyFYptopY9b/h42+FtsmcW5u06xM6G2K4kVeXPeGarvniR4/FS7
t9M41vGzXVOpynnozWwsfhTVpYg0ohmuuYFpkOheX+8lAGgH2U2AJdlOWRxCFisv
kLg5taaygogziNuSUzrD3oRCdHxrFXUNkzHwLFoRX8uYX3p8jQnkxio2k0YUHFh2
IURKF+l8GwpAQFPe8Rv36flMkyvKbtoiqk5nNIc5kxq/ywvJ96gnvoX5Rrjhge3f
/91F4cI9PFHAZvNUzyLoPMqpcmRonEDAoS7w4jAgbx+JHyaobyE+/W6bcWHOI9FZ
RqPVz0HBxi9eV//2uWh8YaDhi1AvLAJgKCKLMBOaQ1de+u+PQKGYxs5wTQNtoLlq
HLDw40TtLzXuXgcTko0qZhFf9ndtHP0DQIGn+9ZBWYcN4E2PPmsI9o87EnhM7QZo
IzB2Zdn4IGOnwdK8E8aVwTuY2qqHx3jOsz3lTxESs0w3Fq7SDiEugHk3S1zfXFNm
DUbhKU18SrsH025GySgF88xUEnknQtbUdFZlXIYMYgHDOIb5cYIsbgNgljgWLQ1I
N5Gu7oDMjhzvxNQj73Ydx+NVPIkhFbIHG5FiX0pEgiZs/G0FTCGZOMQh/nZ19Tij
HWiLgCIlTtij9RhV0/RNMxZAH1O5iNlaN01AlEsGxAKOAR8eFOXM+9ZCzsEKwpnk
tkZQhlAz1s0ERjBEQ3CmQIZ9WUx1FGXv/VZ7FkfkXRgZk5O/x1XnwdphiW/PzGqs
KwMdHpNrXBJ9tmy+vxYmGAQSdMvjhyWLnD7aS+YEFEZxuF91cw/WWLrFEMWU8PWi
bO7F5nGcv0YS9YL2kcgc39Sc41qe1DENqrZW5CakvL5iCspAetrfE4MspdTiSWRH
qi+a2jpkqNs6b4tS5SCeOBBULgGgCM1UpNKLaqeazUWlB61uZgmD3slpGxQSu9TF
9Q16LsPzpK7ouLQQ3hxQfI0QrHg/mi5/TaBEjUEfEBvZv4MoZVxWYsEaBnaoO8vA
O1+1QHrndO9wcuGGhSJH9tBFKUv2KH7979AIiupfjM+e5LIoDP+V0ubZGW6dDyJG
NWnpL4IZoNxEsASm9zGlh62o+nlDvqXHIIIBp4ZVRNWaZ7nAAtjctXvXafAuMwce
RSrUWJnzP5eSK/GiED3Ium0UaTVnuFn52qax2MsDiw0ecFEYxUz3kxap2EbeCVcZ
0vyysN6+yT3RC5ujNTVeQ2RUS29a3j5AZ8JKLLTL+VPR67vh1XHjqFmf/NgX+dKD
BZ5pgSzUCcCpoSfEMRL+O23xn1csFszbRvYZ67MQQPAfnGW/0D5rhhN1jTTg4O33
NHwFHfJkVut5J0KzGXauoM8pmi1FUtfgp/KL8lGb1Nl8iVTX7GIGc55mJQfs77B+
kxoSkUbSlEPPIMgnyII4c64NWdBS+nmOzi4ipFjBM7yT2nddLwPOntBec2AMdWpC
C7O8Wy1bUheJcGElG/rsuZAMdjLjDSO74fAj83X812LZN8D+qxnUGiHhvLWoEmVk
5ECijEWU4Hfm7SzY47wUAN4YlbBjTAwxJ38A9//QfTPFQUxthKIeEiVF5NnZs/8D
19JkqlH+GUwupddj6zqfNJkNYn4wYz6Q0of+2EvJO8DqKKvwJ579hY9i1Qcot2J0
Jt0Wl9rGukcjquoVzmd69Pg39rQA+PbJ/zQ5NWluiiDqP6WlWQPJhiSlhRWcjD00
Z7fK3KyFsa/AcoV4AXOiAr1hK62aS/aSG/w8CY9aGy7/Ktz8nUmcQm/gm22QD+o+
g2jrriZ9qU/nE1CL7U9vNc5JjmGOmZv4GaEC2woFMjbqX8N1zlJhvAVcY6qI4m/x
KTaia0OPag7Q2BT5oKtSDJXLrlJozdiwptFItr/HmgP0ewmm7fDMoWDpDw0H+jdp
BTKnTdV562PzGHxixpW8lFE7PHxXBvP5KQkHm5TOcY5+SL6UE5IAiFBcBSqRlk4x
lrZW4YnjnrvS0z72SQuzk7QBoyxzYawLTvAA3Ty9vo/iiImAkA39V8jTWMXA326S
pw9jzV13sQFaTImgUM4zKgRygnnMIk0hLB1xN6d2A8nx3p5D7/vkkpxKKwOV/TeR
U4fY2SaNhrzF7WE0ZKfR9BkKq5dM+FoyK240dAPxb1BMmMeQ+IReehFE30Csr+KX
G35uUmbLIEv3pNnBj0noGFEvmklj0koBUcfq1EhtFxW8XEEjJhEvOBcqMtN0SM/1
VuwHeMGoIxHsHuEds2oVvQsKGxPji1CFZBpMteW2+EimATOw+8gI/+fI//EAngH4
saJbmphkn7I+4FVIxBIjO8clhMbLJs6rzIw78r4VmPSQAe4pybK1/C7WrlVzRXCA
pYHLFPHxGgn3yvzKIdzPF8B+0QCHCn604Fev88pNfKXni65WVUZkKQiooRN6UFrc
72DiwplwihSWIarSWeKt8bJuwGjwK6anWVffw0bNfb4Pp4EKgVTZ3/3Qf+XT24vq
1lx2kzkcF/4I7vGY8kuTnu0mKWQxZrHlOvyj5SKdrOC7X1uiRsdI28FjY5LVf/AK
FO8/Ayi/OU7BS/RRbzK9ZMML13BFYs8oBcfyfhn8K7qUXGyM8KdOIiMXBNWlKps1
r3PuKFYPQxovw/3EM9MZkpNAgPZDhoK4KYYhE+HGHWtPTjVlpu8rx+lKrB5w3CQN
58MoeUckDFd6PI+U6iEasGbMjknQC+lNkcY0ACv/UEAuK9/LocErSRC/BeRBHuk3
DMbuc3vPj5+566w9Tj6bnwoU3I8YA3KomxKo9mZNOthA9+nuQg1H9y0R2TLCAgwM
n783VGx1ccigwlBYdrvZAicZlSSVC+Nj0WfOyHxtFsH8vOKED+Xozv7UnY60dcGH
4poz08l6N0lgTYvvKZSqr1VF6Uy+fml9hjhcYnRZHz3A0jJjCJ1aO+vCrTaIkjrQ
b6O8a6MvjB+RmAbJS28qEvHqf6Kbq1pfFv2yDVeY6OHLhhoYRQf7Dgn3DJtPTAkI
esJACgU4C79gjrV5pQ4Ouc5xm5WfwpSebfhSAcxT9xVk+yDx2g73Le2oiukPKb4s
bhBCXTh1M1ACwwzSypJLCCBnyu02pWhSTG1QbZ1GzGEazadNejRRxTxb3MrvAuQR
c6cLO3Mc1ki9dxlw5VrvPcumAqGNQGtJM55wvXyU8yfaSiEbVhraDliBiSLj1B07
tnqMcMy8fV/oDJzcaUYdZQmO7mmAKWe9W7Qpz8HriYmW2/c6yOEjKNwiVU/XSfAW
l8kx+k4WJK56O989uOfntcHCtRf4jRpNe4uSN9dF9Tn5LMUtlLRACoU0Kg64L8C2
q3EkOUQsO+k1DtQ3WwvfyKovlQF/RwUXT81fA0OHQK9P+qdqi5gAdII76TbyY1mp
kuTbCGy+KAtK+07Nh389r9fe3Snb2JbdhAk7suZVcRMM+Y4u2J9hVG/nJ7w+StNt
oNJRcBjSeEKJRpFk2craCOFSMEtYq0L7G1scK7XORAA8/gNoCn2/WJNbpJopRj0e
SM4KSq2OT1PNcvQfwM3RFg5Q99HyzrbCFEIEY3aANhgtJ7wOsM7Odkd2EkV4Vx1d
ckYfQkXCYu48OgTcuhSPOH8xcxQbFC58ViijLqQ8FJ20Cek7qJtED4FWYRNk8xL+
hCQqWHPpUVebu4ClFmAGbJQ4DMZBqFFy5TqEMxp3khNpl+Q76Rx3NzuYARh+4Sbo
sTC8zdJF47m7YOFEJPa0rYTHlSt9NS5RJqB6hXmr63KLrQJpxA5OvGbcBOmer3Z4
usYorGxVOrqbSfIJK8tnjgMObBQG0uDd5AielVIUZOJYXWdAmakdGphe+b9khe4d
iKowotEfVnrFsiSKx7N4HCagQ3ado1/96uP4Q4sktfMiPj5sinDHvnJ/bsYNO7L0
eSPvNy+2C7RX8+DUdlD0HjyUTfk/3GpIwm6L5iCNJT+prA67gtYPRrBDfi2DY8qe
t9C9x1ONSKSRXoc6ft0kk5/VW4P3IuRcdRbp71HLC7wB4+kq3ioAQqE7viZ7H+Y+
LweEUk6HVj5kYHk4wFeEUR+dBoIP8gHHrPET5iBevfUeKwA8DrKe5z6aPPu44ANt
9ELfDPEgJvvIyuvZHyZ37W3fNPyuN7Z+vFFwTyXj9jxGFLWbyEjo5yotEdlYbxIX
K/BcL1wJ8jCYi9w1y9o7Od/UnFM2PlkVj5uHqShqikUP3hPrRF522gZunCdQcIxU
IdcSbg+WsJoD3RlKHgpIJjBHLK8vitQArelfCjOlmo9assEay+cyrPJr9PqbaA23
3WytFa3uk71HvezDcLyDZXqvMKk/3KnGJM7sKAxQAW1HfouUhN+F0C8PXCgJGjwc
XXNzJ9YJQn9ykXuKB0nwksFpSwVIvT2eCWab1sAvn2Ov/2VUoQOxJoCROfsGtjQR
BVg6QJWFngFTarbCdId6DZMv7S1j3k6GOkgXI4H8SqthiNSnwj/NS3zy6CfPCij0
`protect end_protected
