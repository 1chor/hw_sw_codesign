-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Kwu/3h66zHVwiRiuHQtWDEfmu0Qi47GKT2h8jmrf/1cYX2VJTrkVcFw29UPrbiUHTml7VfrZ0p7z
bFXdt9OPTheFfSi5bVMUSG3Hv1hlxuvxzqdk/J/lDCX8gGlf1il4PR5ddzI47/xfqRrSY2Hq3uOs
ZS+K2HDHjkfEM+ViUr5INmQY1w3tXpfxSscUeJCPMQiCFfKDB9+GiuVfVDIJsR/0SgxbZ2daT4kz
fNDF+ixC7O8umoxlWWuu1uNAzTH9XFR7fZ0UlxCbST875doHLhZETQFN1xbbIN3NU7jMJfij8h1b
fNZpU8aAxiDwIhCgBAqhajTSiuUgkX43HFyFHg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9408)
`protect data_block
LfrMFqywHroov2fgu6rk8ToBokxvpslkNA0eG9r27fnwRO0YnKLkHrA1IdekcELcdMV5JIydr8or
0Fb4oVj834Y4NsCPnebjXZ57NMiinCV6stUhPhdtrMMI6Oo//sS5GxcsPAlguPl+MyAc0XyDXlic
E5H0Do7u1VxpKqCMEPFGHsdE/itCZy7AKwIVxiaWwhwC2IaCx3vWpSVGeXXFDg+jdD65Pobb5rUi
WOPej0mbKhOnNiZ7m4Rzmh90SglWZd3bv0PxN+wgNq5NRajNQHaMXp7XHFjw/psncCzSqOl5F2L3
tPo+GhNekN+a049Knr/0Tia1ab3XIkiZr+jb9zVr/iEWDgUYo6YNv+xLBnlkQYX59/7JnRxV2x3x
J2RdHYiVMxxUBXmOuMqHMog70wPgZ0FKRph4hseKR/xSCZpQpil5CAhxgmIInWxfctHc2JBbIK8R
0whOufJ0LFIpkoDg4+HuXu9JSYBNDyiLM54OBO2wUvBfgrkr435F4DiMyuARGguRtD55TECZ9v2f
FFlMXl6CuB1Ct+AMCmb46xjt99vl3R5saNR8UbY3dq9B+LfkCvo5ik1YFZ6SyCFnM4Mlx2lWzOpD
YALpjvodef2nuzsQpJU9gdGeU8Gh0X3TgYmu9fv++509UrE3wVqBxTOUWvboIuoit4hmOVw6uqEB
zKfnbbCqUbE2N0L26bqhWgCin0KuQt3l/GOsCjHwNa0hF/s5qTHSbTfov/ktEGFDL4knT8bs8jK1
Bv0AVLwM0v2byBEyH4DnA1Cq9zmrjwmeNhIHGEQ54O3JooxmlsNKREMhwYai4YqQMWPVN9n8zBMD
wQqEhydaJU7TQkZ2Rqa336WD7a4Z7PYYpInPHIBnVucrMdaUn7AaXZcG9Nrjj29Jt7s0E0gDNTf8
MKcoiWjVdyKbwFnzKUJ7q82VIE11O6IeWb02IPmxeehRSHehwVzYKT47PQPqpvxfk0dVeCpWblSS
Hxmcqr8asVXriiBsDUcSIEfWAmTwWK3iPmhx/OxEMGIDtNt4HdKNdhI+EZ+CwqIx03waavnVHpD1
04vbZGpEymPbn9AjcfexNyifCNhqbM3TzZ8M3V81BtDMIuLsqfk7Z2H4+5+eZpxVb7+cM3AIwaNF
9PDIm0b7/nIOfQJu99w5tHwR+VuK9HCKXGd5VBYtNNx9a3DOCxchrcUkVw7QkRn/OoyX9QK5IYKt
dMArx/h8AqBdfHwc0Xwgo1cffVLybW6yqEoLBGsv0DRsvA17XlTdOoD2lkA/5ndJ51doJgR5b8HQ
PUajctR+2OOUaVaA5WdfDA9Tas2W8M0pYXP9vgbraPrGDO3vkqmmSUd8NgZjMcZuW0pfIXm4uBzO
WsUSLxi3ebMRDMQj6B4fkD3iAemQ+fU9ftV/IvJAbUDjg4PLMGsknE4ewoBN6e966s+pIzEocsXl
Lz3WLDfMKjBQKKpxS5za1Y8Kn3CSJi9wLniGMMvxDADm/fEALykVN/W7wv2jPn4YSR30R6x9lIcA
MFjwV1OlZ80iN7szFL0FKfw9bOfJ8FFPKPU4G52Dnnv5ClqLk5sD5MSgaSR4RaBmUVxClALS/G1i
Qs+gQdtq7cOJHilDUEp3176T/koYV8SnOowVVwBWpYLZBMP2mpsBdPBFFOVL60B4kbnEjy3sGyR0
9tD8hjs2b5SeAnNykrvU+il1eqTRastBQyyAl/bvKPp/aAfszTz6sXJqfeT0NjFyT/v0n7dS15z9
uCD9Q9ynU5xvgTNFzYteAXHQ1pAwig8zbwsnHwbbTpls6JZzjdpkQC+GblRrA1NkiSmdyuRV5NYk
Iju7TVWa6f/4sInZHWz/qSAP2DJ0Me+43K9gzvLTrU6XumkI9h6MgXCJMbfZO1EV4ZS0TnjwBkvP
2tmzSamARe6YtBs+0z9OsXdYYDxVCIOiUVuDuydTJHQlUoMKWaRL6VuItp27z3u70spfjay23rFv
6RvYrg7/C3HzfkRnWqglj3ZZBdwAKy+MAa5bVcc1NlfF0CxjP5bXNTf+R0aAsbEXHnwZNENOLtAe
pPp6qboB6uku1nDV8PVgfbzo5Z6kVMXhj1Ih9jH9zuNz+YHPUbMWl7euzbXp36VyhWkdNyr1ZNcs
ziuHiZX154ZvUnaOK3qWbaYOQKP1nl8l8uXbMv9DUr95LL+ChB123+tMrD1OmCT5RHDUk7fQ617N
c1ldQNtQy3wTurp9pdD7zGpUeNreikKfCUE5QLRF50TmLNbu5zsIz8Qd1hKgyT2ZK2z+J44rMRzW
EBupYFfFCR8U99U4bu5yzxC1jCqa+ETCFMIcf1zad2EPn+W7sDNz1C5kfzlHKlfAAQcqARP90VjM
4iHTTCje/xgUbAXzC1J9akJd0azhuOMhMSo7RwR1snFfXpzqTUakUYliuDCqdEUCi4tacq8WYD57
GN4NCAwTNoQSIjiHfA8lcNxRX09wnu+b4Jn4TV7tHtb/sIxqi2RMijWeTv2gUsU/D9ybDUwW+fjV
9rcgbLq8Q25W24YyykKPXGemIt791lNWIggR2TTDgN18OptQmcRpnLwgHBUSaCr9+q32xP5fqq9p
wDx0YDvPYN3t9PraCiFYy0S0mRZwXaNIT5XxE+fYhB0AWY/3du0WZ1qBKRNrfbTZlnQ4hqKWvhhR
r0En5Vw/7+y+TL09yTbJK++keYPbyiU6WcDqHSnUQXYsX5bJ9f1+Gmgo7YcUA6p2cH0k2C24+hXl
Saf6cJv2ui9I3aPX/Zfc6relbJR1Dz4CmdIV8QHdrtn2AnWVCkwTrH0D9sILBFGuQTBdj+H8w+uu
AvbPcRJc9e1q5Y41gEkWKCphojYIdrSnT6rAb/z7dr8V6AojxX9FWO0t9hcRyI7QJ7QqJWkEY9Tl
O5f9ti1lAWyG3Xo2zlgdiWQFoPuwCUyUAKdNs23cfAa/cM5CdSgKkrkAkEfwvF97BmRyLmKA+X2x
kLQHPoud54VTd/x9fziSD5DmwktjtaUELy70cuuVUMI3C93gjSnmcNHdxgm/KOwGQMwGWNaI+ROX
HYf1JNMtBeUsBvQfY6XY/pdTcFjET8OLch2LyQSTAt/hE4G7ZjenDrr9HRn3Ns2p7gfUyjztY8Wl
7Nvi98dA5j/jCYTxGYcNHGr9vtsa2evskWJq3nkSoEEPB2RHZcTKV+BorT3l7N8msrt35dN8COSE
yEd5rAoFK0LqMpgUM9vRjkO3YrbOoOs/TuUDOeKlfrHqHJi3eOH7eHEmKcFF9UQVxYYvhsIq0lQp
RcaYLcLCwe1vhGonXhopLxLW7kCbJYPQ8fIMYD/sFxB1ni2H12u+4V0DjDM/X4QTzGUkdcDyrKRr
lVJ1zCXCzuUl+MetwYM8+h46IVgtbrGXh02CwdLMhmN/Tsf/fl2wel4HMK2kW/dCDAIpaYcutsBK
kkOliGU6VZLqMCstS2KmOdWPioiHsQlIWKizKKlb4pkE6lXqP1uHM7BNKdOalF1s96uWQxew3s3t
IG2wHD0xWIf6kkDYYArJpb7I5esrFTrWtqrpGJFsjwV5+UUswE7Umh2WFMmIdDll0zfbNKssZLwu
2kg3CFl/vkLPgqV7dOtqKDcFpRsXd0PmEEGY0x47NEZ28n+jrAOw8L3g7CzRJ2H7yu8tMsV+9ev8
x5ZpMBdsyhUKWVFi3JkaMWU9VwE5c49/zl03COTkgbrVkCoI7X7RN3BvfEucRAly5VbiYytrAY1o
9rHOlHk1kUEbvwOhuIdkpxQ4DhkmLJ6i6H++ptcw6C2VAXQfiyV5Hu/qSXoKW6yLruxhpLkTo78F
ao8/j1Ygh/Dl8JjSvz3aYKVHbMfO1torJE+8GdE+HcR/OOB9KUIOTAqIRYHKOXybRr2aZZ3ZL80a
+AMunhaJ366UPavmqp5a78UdZmXXPkKJyuuUMNUb/JyLm3pUatXK8tnoTGH8pReGs2UGk0lEtbBx
LRiAMz5weymSJWnGdljeWWEoOvQdUOb9zhvUMO0ACINYrcv1N11Iv4RjTlKz1LGGGBmZamf/vb+k
g63TxOY5l03G/9k3aS20C9OyhkQ9I6bTKjiUH9FOMLHpDXW/cAnakgiK7T841peAkDG2OXKekhvJ
ZE80WCFRncdxPN+X5yGlvJtHukAIQxBK2JYcZHoJFUA8UZfI/qSVx9gO6GUh9W8zzdO4BWCHinfD
2HUTNvM4+zMnyHzRCDUx8U9HMR54hVz2ERtt9cIfQz2I5w8NQhY/AdTUB0xyl+vIlI21GlINjBQP
pCcvreMeBMlFdi2tJHyYKAGp+gSJY8asfbnbSzYY8lUJkFjFcwrfYTmRvFMc+65190sl6lJ+tjmr
VfiNlr4ICrGYK81WxO53xTQGSvLotWkEk8oGsGDoqrhzXcptSdHulCDVrJjPNnDRw+PFKjiCdZqJ
uYWlRCwMxxFxnY6wiryqMVqO2izYYRuS29bUZrOSaV8UKboXvZJqzCTWcCCSwP4c4oBNlB9ts9KT
bBzs69jexty21kUyzjJSL2hAs6SApUN+6kbYnVQQYC2HzrOS7GAxab8RZ6UD8LG9rBkvQ7Vh9S58
zivYviKTJNI3OMg+mHkRr4lkGQDLYSW8dHWGhHhdT8VMB2KYjeJtT8iqO/K74SCzZAHt8wXd8FL2
SiDMIc3LMpaRnUGULoerD/ryMfd3laImtSM95PMsqeutLl2kl3MO8UH0fluajYWvSVpAtO20bILy
m/TH9kUfIsddeD0UK5P5bhK4x8XVjRzLsMZUI0pyEwHpsywFt4/JavNXhgf6Fc2xhFAkuVfyAL4E
VcYgo23W0z0MTDqI7fxOuE+6pR8B2Vx5mZKdWFmsOHP5Us2wp+KOYRLGTsap8gnTG8lKMi5Q6Hf/
uZg3BGPR8T94G0MsnLrZq5oSR0Wv0hqO4GRbE3NpWxkP7aCyHH4KFNbdTZvvGEw+EJZtbovs0uwK
YQtHrsyGSWgosXCRoMI/11weLiycG44TIpqxJtYk+OAg9FnxJIe06TBFDNDJWfVNtkuW524ZPxRv
CPt2X+EQM18EL2uaFxOMM5JX4Z1KYHm6QQP6bx6EJJe447URYkK456X6NXkcJ/lfYt3jyXAwH915
3HroMO7gY2HxT6SoXZX7qLuYGu7iic//Q+a/vanDYhI/xL5UJ5N3XTItelmwqTS98m9zq9ElJTgc
TJk31mHFlaBhvsOjU/n6Y7YTHh9jjkj1N80HLNsFHC0+O63OaA2sBaBrPMplVEjwbn1Bi+A3UJti
Ki1LppWzKGDBj9Q7YWH0MsuuyZlhOC9bHzxyu7dXCzplibQh6t54Nl1W5T8+mp6+NDLMnazv0i4F
2Ffj4xbaR6L4856Zhk/3zkgpIlJOMueufSp0J6JkAwv0vqUiKucyG3nYobo5Ec8A3x6C0/xIRWnZ
ABKm7AlKeaTP81xo5fNWp+jcAJkjav2/V1HdwuyuihgmdTplx0txiMwkQ3FNqvWPg22jTENVvoUT
so/fldphlS3LelCvlZoW+Tm3dYLHaTW6rouS5b4Jy5MScz0gYWW1eyLVXWkyrfHeMCnIy3s1Jsrl
i7zKUJBDqooAofQTdBSIc685tF6ifrir1OFfZkpmmKVotz9BH9r6n1ZmgnCR/4Rg0jZEzC6ej5qX
50CwBKtmoM4ggqNIeaOGyiIERk3gV/IsuZ7qu05cngkMB93UtWjKThNK/tBRDTQ1RPw386LXdvqA
y+c7SIeyY9uXrqum6JM3LrjHJ3/E5+33nII+671oI7SNUI4ChhGRnsy+BpbKu9HkWC1qZDSWBd0x
/nc+DS4NNayK37wsUCk0arjJlcgbu+LmFyjCfx+/ZP1aWokMnobDhYdAb+E0L85KWuZoyv5gL+5W
U90XoyILoUnaHiBdlHSXjcn8xM9exWOd+JEdrFHxzu/1ejQ3M3cJxM72OEffCXUkMJnM95q23QUF
cN+PIRqqead5lbcX9JuWZ1pzY43RufYK+Kzxt+UfhTNuysEg1MMIySoPcEQLhigWE967XrKUraZE
tUyzGdOiWtrNHni1G3CXxBiqQ2bbHrboe1CzLAUo82E1jyaPTgsMmiRLdnFPspyW8ZbeMe7HJZDe
Dndw650/zkIagXOWQQqzWWpAlGxDcD2rXfVgRORg38fFHKyGxbBgEKfz5XzVevrINwESHGZz+jSl
UTlSjgJmLq0ZkyGeCuZWzftnG5wmuDo98G4x54Cfuzen2hea1MEby6oLwgx0U82+H19Ie2BkXNAr
9DN15yTNwFMHczxJjkpCEsBG+SpqwQL5o1roC71M917GRcscJEKBM5RPpzDQRh2ejbOfbuMaNi1d
D8+Vyhl0R3Sz2bC74O21E/A2xBUxsgjFaQDrnffVJjkFwqA0Zg//jgcNAC8Ljqg7kTUtio9OVJDC
D+QSkliEkY86kKakUA9Pt7ehBEc8JL2RqryZ1ucuJuGf2KFdWsoSbRcmFfXsHy3IZ2sSx7drb8vg
MGlmoOO10QiPsF9WQ16MYyz/P6/y6MoPKM3JeMA3uVGJMnQf4Fsz76aLaAjvhxUQFw6zI0m8CAo1
oqKLLI+D2Av1ly7D84DGbQLdbPY+DbHrihzfq0/Z4+DwbXpQKtnihPoBy3bIe5va5fmF2zfQTOSp
yPK3pSfLO+ngOVGJr4kph9mpTljGNRQvQtye79y7cUg+mlTcgVAOI0MhJ3l3h7PB58XutJApGcrX
/2gHoWmkJYY9WcqBv977cgZvnM8SMbFMOzdkSAU/ZIihOcnw4L/xg3QTo+Y4bnnDHctr/eBaxjKO
ngHZ0C86NvLmshOL5PrZNk6Q2pOxQVk2NVpHE5XT8LEhAzBBgyz4mvJw0fROwLHM84v8TEeQ4XQb
kOlDO0tv/qE4H5dy4xttpnvm1kwgBrjtJ4UVfAKUdgFKnWIjPUn2TmAedt9Ur7nfRTOgMv+uNdJv
tPhxfXD9B8bVbllF1SFUBHv9op8JFN+B9maBq09WCVgdYzfmX2KmF4nGGIoky4Eaqkhj87VG2hVx
GF5d5tWZaam5sJmQA5J6ppCQaAGRd6okxZIf9DxHEwfu1yjqZWVklplhOYgiTbPbpMGorO3NIA2Z
5JAQSnEQSKOr1ubFd0UXx0J+CsgS92Nv0Qu0LSkSiPQKkj+Q6KoWzDkUhwqKy92Ng9gzPl6Opb50
/JkV4tJ/GTX+uVvMYQeWZpSslvc7dNPf4ta1FE1SteJg771cI3HfoVI2q+4rh3tVjlnwVjPzmmr+
qBKK/ou45DxHWhvpTX/xeIHhswL+oWT3LWfpjraDgpCRZPvGBLzZnhq9Kn6B/TMMqoCoZLTHUHec
i5OM0NLZJlcXN8iFb/LiD8UT5SsNENz3QuJoTm7F0vqwl+Tb5wp4uKmox+VArsemSdaSHfBxsWB3
uJ9akj2TqRCZmXyOpsU21KDe0+HKD2x6azWctBCm+akdmdF1GdgDQFH5OtC6zY5+xtq/O/1ZOWGu
yQR90s8Mlw/dVt4PL6PEvMkgdWUIwpkTFv+FemvI68SEDiv6V1D2hlAiThijwD5LgUtXEGyFqe7q
uJpeASN7SOib5VG1uBsxAeCdfo6DCfc4yzveG7gdRfYT0MG7uC2yK9oONpV6w3BAJIaCI/LjwbZC
XuxVhYuTXNWDIhZKz8X/MEqMxPoWcfC5TY6Qa+e+8TQL+FZvOqgZuDybZRLmbLznvMNIS9AVDky3
hW/JfLbgn9ZePIMML57JBn8P3xL6fHYZZx9poj9EAp764RUfGvyVABzMKYo4L7LLrfYkXecnO7td
9I25Fp/ze5Ux4DcrzLDkpNwBokZoBi09FFNB8rbtl026F2Fq1W3kqZDqHPhLxCARGKwY+p+OUMev
8hIRS4/cjGQ8Ferv0Qqg5O0xYW63tUyC6FaSbfy21AJJ5bNirOvC+qeex7KT21v9Gie+kUjR/rpI
qu0R4xAaHB2n0tp8bCln25BeOsKDbgI8HzgGWj6WmbomvtyIu+BqKsd/XDfOUtesGi6s0GXUop/D
ChTisjVZ9EbBEVk7iGa+E83Kk2VIRJaGSc49HB6QB6Ph+ubKUTmvvJNxQnNOhcA9qbfZZR3Nbedu
mTseU2rCPUj+vjctmZMi7v4xGfzBarLRS6HQsvNRBM7rUxNKmqSuwlnoRmwiTDVPIdAL34zAsbLy
MzQTI1P0VkxczxP5kj5SpEjayNBBSF5Y1xSeBOwgysJ6aQW6D7evsEfcGnG401iFE60wlXLVscEK
p/bEISnB+ewlO5LNkbkpFkllduf4gms3TfPcqsCgXqtN8Flm/hDaf2n3GTr11Pbz9ngM7qjMub2v
Cnpz5NC5vZCo2gXO2WNifJb+B9Hw77aAK8iGSf8M0HDsyAhoh10et8YYhx9uXNnmVTy5tbWpNr9y
qnRuo/C+f1FehHSRClQ5vCrzfwH4Jm0kbzZVuoN95tgwZh1ICGiK7CEEk0I1p9k/cM5okVdozWpV
r4EOxeY/AiQ38I8ph6c3phTwV+jx+9VR7+09JabQf/WJMyZmYZ7hIAUDjVfRFuVX+kbaU9PyENFp
I3wPpvDEAo9jy4rFWaW31pGJXf3mFbCSRC5b6c8rEuPGG2JOfSVGMObjOwVoJhQV8EjmUM1h4x1D
++SaNcUJYETNNHFyiFgEKcWWCO8mBsat9UuBMilQCPVytG8fdTbTuYhTBbhJuMO2HI9EC0FlfqP8
kel4etyf+nlVTGCxO75+29eHm+R9+2m2FgS5itguh/DUmsa63dretLQZ1SzXvlpDlntJvWKjOfdA
kYjCEqYcoAdX7JD3aG4bLnZiswQ74lNnlv7CXVfZ9s9JxOg5/YtvgzooK1DBlmWrH2wVSgVOY0xA
WB63dcjcDBlFQj5Hrf+17o/SKmnrpPdtvE6OmhYxSTkjDRRkEcZ763MUZZyUS2r1BEdtlDBjRb09
0VH54CUfvnKO/73FFWO60vMbyhGUtv04d/Q3cUFfTHC5BJ0qPY/N0fQB6tKDVZFCyRkwuMHu/OzU
MNfINjXdj5NbzFw0GsE0IFaPwKPvyakND/qDozauDsQWZegNZBDCv3Xa3KMzpCRqdKbROKtTiX7o
Y8jHwA63HgVPKuadWkxtLnGvaRz0YEBvBZWfRD73bsTonWICd3ZOekLqeiiYQ/vphb1WXNtAt3mH
35IMWsTfixjYHj+pH/ThItn18lAoI/f8ctagRySZOVYA/RjquA81KZeZLd/t5pufTqthmsmt4oMv
XTQvwfxcJCCgriOIQkDfQdikWhsm4PVu4cDrowe0V5y+jHHz6nMX+JgMS+kis4+i7bYtzx518lr5
4rkpBPoGckyboMd6Au6yKQD9Y9FZkPURkDrIycxXpCrQpjXpPpKzMRSuI1+bn2mPP0eF9hgSGOit
fIxECiy72TJdplBLMozxCJYwESNhdyUKAbNDzMUqYqmyP0TQozSv1sYukQq+o/Brr9gRJrHmaPqC
RKtRZ6QXgZyZPmHDdxmTcoepgfdJq9U5m57RBMjyzi8iwxcUqmvMLZElBirWGmjHT+qzWdWM3bw2
r7LFq1l9jrCov0tHMuxYyJW9ykRA2sHH23sEwde0L4xaCMKAd9cjs/826iYpO7BbdW5E7+8ccS2f
HXj4h1Pw7K3/bl7GilBvz1lqBltYRKui6W4gJdZ55v2MxYimtTJoe5/YI98pvQgNH7NR9OeNjPwu
pyTrLUJIIbZf8IlgbSqFKSWEBsxja0QgGR0hlYPvWghroMWA25AHC1slRfmRJo5Hnyf2kSRG5lsE
y9Dykkgwd+c8McSSArxfTNqGNdS9xRLTaCBGoiVn0TyZDVh2/pkvN5NoS73jiVlbLpzR1USk74Ig
v9T0LKKgw0Pxnw6buj/72ByV2MNEEdpohJFU3cPc0a4dg4AlXKmDFfMklbr+JFrlN/2+FugmfkiW
EHIWmgzqwl/cFV1rl7PNy29nSXNiSbfewtfYPV7E/laGUBrgW47x1jpUK3Z2tH/xJLQgkhWwUA+1
glGfuNq8GoYBCP5VciivYh1AE35fU2zUVWen1J6j4J6+DkTuahcrga01HmKZTGp3bfLqfn/ZxalT
+NteHEfScos1eh4S6FyLps4aB/XQevnRq3oPNqK1VqJrxmBxELq/FfkrTOe8G9CpDjx0Pl2NTwmE
HbdMEI9awybUk+4TuwpHc69Olj7SVMPa44XbFv97rXGazJ/QgT4tA8mEm2ndakSAHiwqz9+lLMtK
D5dDCRhqEDGzjufqcE461HkNo1TK7Pn96g+8MONtBM6fXoLHJNPBfoHUEf7EBFQeNRvZbnQvrW3L
pypLwsq6o49DiR/KLg3U2x4bydMKbRaCmh/511tL0OlaqKrDfkcupGGuruA5HL5OIhn63z79Oqk+
R9zSg9BFWIVARsoBkeTBJNtE+tBDHWgGu0SlPqiKiwlwz9Y0uQhK4vh7y62oGRa4coHXmIKGCe7m
3LVDlEUkiO0OpqtexXkkHJKlgwjaegl3hVL8ssonLQgJzyw3zwV64kh8urzLDqKNHP8YyIjDNTRv
Wredw77cLDpV4AJXC75LkKYT69EkC6Yxp/ot2aQLuMIykGZwRGDwa65lx7FPSoUkoq9TtkORNphm
/SbEwysRUnsitl7mN5wSZuOnzzPfJ0ICzVYNLrjbbCOsopsT7XdPjEbOap3rDF9HjubpFneZZzR3
/+N6/HodjKtkuIIYqzXk05SDJ9wgJMKwIXPjJ6N7h6uNeDMvRe59/Ly/AU5RpmIUNNKDlHON6lTb
k+fFVykaAEiRKuXDu0LUGZh9sW/6qR0spHLjjL48QXkut1/7x3R5agLfo6+Ybkwc7z/gia2uL+L2
0KpPRuXZR81Udw39MJ4xA8xevlw86itmrGoZvnIIv5qN9JE95Mhxj0C8uyXaDLSJjcY7kJt0wqsd
QNQvhgOiKO6Palklah7kAhiL10jPt+7HaFvWfVWPqgLo2whFdJ9wkZ/s95/8SSQrKvFLAaSQgxfY
dVXOrcOWXC/Hvk+llnQFhWUEGgd7p/mculI7jpwWEBuuhM+78Nj2BDzsK/wqlQrOn4l5FjGOgh1G
SuVbZ3Ahadbph+0nj163aan4SAEHeGvgqDrv0e79ytp0ZWHMNqpol5rfv1WlSZJQiM/Fs9AzWgIc
PR3CudnABrjk4UUb3jBTE8D5EyBONNVc8uFbC4U5rrVR6ZRo5T4pR2jGfNsN5WFcu9NPNuHD0bid
blxBaiOb9h/2sStMvAmuLuh0D7Aj3ImmBgEJXfx+zko03BXHmLaGb1B/Mqln5sLCcOqWOR5c2gAO
yYSmsPNQN0YejvPpJuQmuTCkd8+dJIY8bhlWLQIvfe8YwTZu9QP5nQ8yShM/EDAmikEZHAidPy9C
2c7DwrTgjlAOqklJT1tLTJYKcL7A3Mfem1iQHhlryAVSR8XkR6XaTJjHmNAQ48yvC1krmey3lA2o
KbvaoGN/bVwW90dDQaBPv5hOE3a5fhf2irga4mSTv08WwI7aUCiuCXtVdZyVpB239ic+RAlFz26r
TKZ4VmyXmKG9nTpGB38cKuuDcrWuUk9og4YEHJ5RBQrkP+kfR46ke2ck0NqKbBIQos3pRpabF65c
2uQbnh7c8mRY1KHcnFIM/5TeYjGWhR21ciwuHh/PU7B2d1QEF5L9dJ0ZAQqU01KzJNA/TILgk3K9
vt3Xliva1a0GdV5o83TVn/Ro39WipLuWIXKtBBg9jAPu1maZGz4OhAAwxvcaPFBR3bFzQ0arxSRJ
e5qYuECpmSc0c/nNh7i5zOgD9PyMVDCoWC4g65fqcc2VtdeNLLOvcPeg/OfufOgRxgoURzR6vTcV
nkEtirDCv80rfY28amYpqveVuNBQIf4mrxjnXjb7Z2G9KAWmbWypUJiUkbdO8E8bLFf9Z9/4VeDJ
Kbbs95Vgqmoi0Lt4xPI+j/eH5Jv8Dq1YGeZ+AB0MqfprWXQiXi2s/aNqMV4Y3yyKzzgHqGG3gW+M
MNRPPjHJ/kKK8ii2P96BtVYShO8i196NKo9OXe96cZ7YVkhO1YZjCu1ROJFsm/XHxSgyfRS9IgYV
1evfg1Pwc1kSaagG42A+Wcgm11XzJeOhIvUshOnQYfwVZLRjwXhwgBfKh6a/u3f7lAWfwadKxoTR
Fage2G0dHxYwmH7jq6NX2lE7YJ5+LP4j0dZyQMpKEhr5sWKPKWQXB/rEF/shC0BanOVTZOUhQkq4
K0PaIuE7HJWMGXuPfdpGlGEYJpmYH/ihMr62nSqvtu3B2ErWcR7JnJkNj+roMm8+wPwMd12ad+kW
57NuQtGIpKimMyZi0sYpTxQLc/bag/TuaFoRofoIKTuleRyMpg1gMUG5rHYsVIcWF6k/TAp4A9Rj
oui17oogTR0V36KS8qiDdEEkJKbxfIJF+Foqc/dPNcOry3Cvy3zGrVpdI7n1ddrghQdm1PKVStJh
6mNSZlr9HT1k9tb5nkZsFYSr6NjcMXbaB8xtJzEA1s+moG57/qgRnNkiBmqwzjlWYcEuhGMEV1e9
YoNsLEg91GezvsT4KLma/J0Ez9s4r8YHXqIFXKmW6C5FOFjWf4w12eb/CJn5VLzrIHxlgDlh6fs4
VtSQ
`protect end_protected
