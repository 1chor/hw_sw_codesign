-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gNQxWyjjzfubepPg+rzML0o33EAeEs37wcGCzP/XNWZd4lJhFiJyDszUdAa/hQDnZARLUVOHRS68
PfBWw4xrGVrI+dIxyAOdn59wQcuqsEAaIPUD9qgq+o95RUlkzP8ZRdgVXfoZUG6nYHAofJRIeKci
VmH3NzIvMCMng/9LeS9xbb6WbwL0LdmiAxk2urgqMiyWPhmTzVR/bpFcvhVLZwprNzer6Qr1GeeS
PlYcbqUjJ3r1XDyCe3I44GWd3Dt5rnYPabEYWLaRPMnxrJBQedt2fMhwM13mtTTibgryn5mC7EjR
RQa1FJznEO1JH1Cu61H/GUJl8JoO1n0ApV82yw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5120)
`protect data_block
JBZzNZ82L4jwuD/4SUKinx0tekWgHiSpBH3RQbFewjgfHZOZEMLB4T4ydZXDIoD7Yo4Nxes5JopB
FqXcf8SvD/LJoklxIUBfaZacZ1Xle4K3gcmOlpq3dhrMaJrJDKaSIfXIyODixfWKr3jS/GEGTGLK
qG0rASWS093+M0cZ4F4bxGP+PIZJaEdLTI/FfxgSFrNlKUeJCf908ci6xXrsIvjnlPnU2HHFSii9
Hmb+ZySVIPRq8M+yIk5SQcghTo7HzCQj2drUtNHemW4PVHE5JIpQKkWAcZi1rEAXw26fIlR26VNP
g660h0edpYxjq2/5TsOL1RzbAb2KHFPB2D4Lh0rG24DARIgRGfz5QiGVuoiLUwt4J61iW7+X/Fc2
/kAKi86lKVMNr8WOiiuSzcQfM/MQHY6ZkIXaZs1JnCpPDCMy1TtjBWmrZKjU++HTyIFpTUGxUaTE
/+DBuh/lgLF//sR4frLIEpE7C5yXOiy7w3NCofExJty7MtI4OiZNaSFTEaTYCsnccKrj2vebnw2v
3E0m9tLQuDJzttbGpUlyiWIx0YkSm2I3r6L4JLCOS1huL4PUCe0j/GipB9F5POhR+CHslz4eapcy
i3YJW23tX7x2yS42PbnolJlvdOqGDDXNLj+iSzhedWIMZYQUZCrNcFQ7V0rQKdDwws4IDL/bfrF7
G2BV/Ta5JPoY6yzPw6CXD5Bfsq6RLKlHcUKg5AU7Ds96mts2pUCNxuuPTc6U8yyaqAsctrWFNT9G
+3gv32EKaE6SG2bl79D/+QEj40WXPgUmpiibU7/WePSO04njZhs1Qj0+N6zDrci2PjA5WWJVsNDS
BCaAMrHP4JwtgChCEqVulJ5t7asvLSi5A3cOdbd3urbKVvVH3zB22LiRLgt1kdDyxpt5PLYktwKJ
AmmKjOdhpQSB0WW5poHlqi0p+/Xo9USmzagUgy/od7VEA8LRh45acsB5gGb7m3NtJQ65o+kcLKcK
orA//RRCHaWCQR8y46WoC8jLM/c6L0j3vL/XpDHgBv129Ta3wLiuV9+F1hrLKSeEX65JoHd0YIkL
+1yUnrn6ZXSEHY0BUgZH3k4CqOj3G8hHy9vij/lCDrQ1Ta7I6ALsSalKo+g3sxGLyNrn4hv/sisY
eWedInWBNMOHO0fr8Mx2IklabmhiIfC08GndhCR4HxUrhy39H5y+cFr2WEPxVNsQJwjagjUbaOvL
smsh5BZWClwN49CYU5PMiUWeuw5hLlj4SzbYqY6i+Tsh3NKZIPLEKHW1dv5UPyXMXA0gHHLELXQS
rQlmqwB2uOXrQEMnetoXUqOty0rqP32umxnLhuKPGqnlYq5FRRocK8szL3S5q5ey+fkSsi1wdsZV
J/C9xue0uv8vSJrUchhhmFxdksydO5DN0AM8+ra94oaBk1tdWeMreSg2rWJpOPggFQxo+qusn9bi
aZaElcwS2YDlPcUkOY2YQHZOzqRWsTziVbeQFmI3an8I809AOjF1X0+1nbXBl5yaBn9slaA0SBK6
MlOEWT0pI98NCyDU0DP1iJP+Y4H1G94XvdBPQ7nZTs6ypVwTItgMPbJ4iG5rQgUFaED2tC5BDije
g1ImAHq+GpfUJhasJ820jrQgCQVQEzbB1JS/3g5BZ/YErQ7TE65TG/q3Lm/tx42yBmTTAH3NfnPc
/KIZ3VRK2RqJX3eks0sC3PoBHyVPhdkWH4qz9Y+aqm/rGIhVUWaICxhOpGZSvceaooHPoi2ztBZn
D+j9qT8emhZR4XQMzU+R/EBdl41xIjXGi2j+g7nsXcqp0YdP/bkhQiUVzgXi90aRNqMMaf8Itqb+
x309b9mynprpysEiqZB5n01NDJVjZHCcynN/bE2v6B5+9sK/IRMroCjI1Kg3YCgLY3AF2pnuKMji
YAxkF4P7ba18RArTfVFBJDSFaPqayVx/f4wI6l5VUfa4rLnPnmZ3Cl1myi/TfST4x592BCZGfTFK
c7BQ/BTKA3oFW9ay35auTe97AE+A4gzhtC5c79vH7UguNi/TAoMBtHRVluEU0kTZSp3eFG7FPsUn
wOqk7jzbo7uiYrBzODoMSCWSzak+oeHwk1jkbDjBXoU92mjnIUEma85X0ia4FPgllkn+fkFNkRgC
sH9j17MrRN/FxyKjoSu+C9t/clpp5xzd+dAte5rQAspCJ8ccbRHQwtpB/BhZ3ZXoE3Ld01SzDpQO
pFCXvLvTc5qVqiGHCrUBeQ34C1ryh2Am2SZLx/CF07PNZQ/kNGlxuBZZtTSeopiJzKawc+0rDjGZ
XPXd4sLf8KGFobGL+AZSf1EX8VusK6YwtEJfSP/nAoJCZxdrxfHhil7MMeviQ2M4XSLsMSr8+NZS
r8V2UPG4Fn1FiiZ14aTfFUDiVC4YmFr6PHkFJqbJ0fRUOs82aSskx0+kk9gL2BXLlt66wDQv/t8o
8McHUBN+HLpbO3M1FdxCVCJgJnLhD6gLQtRG/R1eVXlqOUI8nIm4SERE537hZC1yzjbE17dyiC0h
aYpqLU/DyvTY3O8X4hzg9NyjRcgayKIHR1UQP0cTAPVNgcTncL9vKEli4+c50IGtKuD3BwgtU5q2
ffKc0jp5AJLqzG5WHMDj7IXvtG1isQngriqGuePmD6++Rdwx503nW7J57j2DLnwxlYrGSnJ27jcn
tIF+4++ZKLllBc7nwCwUvd75dEhMOWsF1nSTGnaB2oqmDy/fbI2lNvPYCuveC/YiLuRKfxmRF97V
evdEMxqLu2QdPXVJgg6/A77OYE8YViDQaTQYckHpn8Q28nhsZulnQE7ggbA8vJoHtnUMMwjPYwZE
f5rhfnmTZF8tEmFFL1KcD2QVuECuX9DQZWuoVFg42J0zNDh4J+NF0NWbQuDo2MbHubuX4MF0En1C
wBxNulMv1M4fP723UeooOGlRLMHheGIwdbymqZ834RIbK9FTqGHZHsWDdgCDt1JtY/tXaqB4fRcj
pnuRzMt30ZxQ/C+h3ujLCd/eUn6QSEW3yR+x6dTlSQlFZJ09AIObSgvDFzA3vGv4eV5qBX2BL0uR
pPw0rPtX/Dgut4bP4JgDOoFZUihyEfOLkPYpUCWvWOPw31QCabRN5AlcEckKlaG7wi+S409H3Qc1
gH6LUZxHKj12LWApNuM2zAapG70dSRFoJW7PwlhZumIfbSudR6DwxO/AM84iILCG/gB2+2L/K6+m
VPQIQ3s1n5kmEBU6xXVbZlIGxzg0AuyxBJem5B/EIAeRidQ0YhBDfHtINYHtI0DYzlPjxEEuu137
t7KLVvqXsGg37NUAQUJULuQ0RzgZq3BLRNRYbfNpVMMmuO1LrmpxaxoI0RQ54+esUpFTedZoF3oD
bceIcLsrj/H4o7PfkoHtZqZBd84bItaA4/4FsM9nwULZIWej3KdylZbUBOOGkAPzuNoK8pyVMfsH
cNz67kIMFP9n3iZqTKra8PIlyzpCHaBcF/28eMtk3luZFKiLgt5tLz31ZTxzAQU7RMJLCOTXsK5G
S5w60ECYRiRDZvlvojA5qhH6WNWtjMCCq6TzmSa1sGgtxLcrJJ8quG96OG/NXJ4yG6UMKbN2ywDe
L/d+QoD5ECczNkVhOkD5+Ss4d8DUoXZGcDRqRRQqcvFq1BYTByRWDT5RAwAYLOlVYvuZr94Jk6vW
p6I+p386T+X1Dgze27lamovIj/Oiv/ew/IYjo9h+vKESLN2FNH59rRkRvAgA90L4jzayVEpuNjh+
aJ56+47ldwqriaTqhc9do/Ra//hhR87C3mqE/E98BmVTZBJI/RH4lRr5aRxen+5jMUwkK2PHAC3b
mZBgkLmQiFJy1gdB1qZ1Ch0Wh9kOIUb5soMJOXNecY+TCMO07aYerTqpC3puOnhw0DW8njGdwRpE
+L1Yaskx2QweGd0q0uLhZPlG5UZQtddKkza+l8Jgfjn0K6sddPNybr23eBtb6hmlywHk2vOkoAAc
KW3rCdymxKDp8slT4/EN83rZe2gCiBGoxbrb2Nt//idr+ZLNyAQUJPIWBxM2BqOXPzOsS+TErTgM
RbdydFD7Nh+RysME/8375g9o69q17gmvWhRhJoEGpevRHXyGQolM1R5QhDJnGMt6r80lbiGBUi6v
t3lQvllj/th6xxpGnER5odr8iyKVamcRtRzsOiwCJiNMD0q1URIbfHMky+lJPeXQzxVvrdKeNfDC
y2HJ+IRY2PczFIjeOmsKpmgHw6bvtAzE8IzJdyZSkSKTvvJ0SlkHwVKpg2VoslpFCYJLnLkZyd5N
HMMzXqlD8fbcATrqARoFs7efzkShxeqA/qkEEwRIvgOwqiClwaOUxJg9c0eTlM9LxyayUR2ShWs4
3NWgXSe4cu3Ln9bS3zVCfN3f9b4OClOH1EvngaS8bom6mb3yG3o1VIaEG9kDCfRE6wTech7vwhUC
dex0jiZyfVtfhqaxIC8eXaJPSZq2BbU5Ogx59zRimh73bc5T2Q0l/Vg1qimPHOB948nKbWQlU1E0
cCEd/dDIYuS8Ht9BJ1+PO9IdNjbR6pMmRNSXJ9Bm0BY5/0+PCVLlAYqArEVapdGWWpWIASg0RMtM
oWY4Zr0rwNMKuyt5HH8kB+4JuDttBsMkn6hYLxGZ/RVCshQ1CzH4d938OtX2GTrp2fHWrK9owpVy
eq6efKmGkdufER+kDizDRSvZrxUJLpmHNgxW0xNeKR/pkkhWj73U47KmWYuZD69Ctavj3JkR93Ww
LiNNGA3nbORy5pwD6s8sbJsQH5+TKyo/2BzLhoMCvTutaEeNJU6AVVSsDTMztXdUho5/SVQ5GcJE
PORfsLELlfDM+U8cSjUV7pICQEtSPZBTNuh/isAIbt57NWUWdCCavzuQGy+N76Nmty/ed83WoMQA
DfmosELQvQrji2KA4ueE8a9mW78Xp4DawKYG+CEGK5jOHCcx3PL/TNfdMoCYjkaWuquHyIk3odtS
bnu6YytzPbOlxnd2LdT3Mc+XffEEQ9We3WazsvnyyCpBQ0I83bMvY0qfP2/XNzlJP7qsTuu2Q0c6
ggyMR4Y54ePJu/UMHkoIRbo5qHAYwPffgZA9rC1o9anAKg+jsr1VJmyYDFelMcZiXT7v1WkOgtjT
KB/sUx5BUB6UMYQwPyuOYPihfWOydoaMaz7BLrBT1zaAA5B8YrH5cfG/E6WgA/FVgjVJFyT4taBh
LdSrt5/6qQqKhfqcWxlbCxyoQZcZJcwLIgHs3fLB96FSXE3fxaSZAgXqjc9oJIW9pQQ0DfWCsAsE
w2AYxO29s/6CZSrpwP4jUF1oBv9G7Tvlmybb7PTAUVFCVjjN0Zj+eC0nJ1tGsTRTcp2NGDl0GpgF
YwLDhhXJ2izOVHLrlXjrnaKPle8Gr6eAdZivl0CcHU8UznSkpkfaiGLbxeEN9c7AjKSq2+jxn5t0
xs6eYzfabvARjgdlOBh2pHZY9ZjeLdR2CGmMc8sNBW95vkUin8GVLnOhBsVdSkrW/ruMkLf3mwD7
f60am9Qg11jwWkouQL3N28eO86CEK7StNTP/MynPHiB2VN9Yvn3vt+GEjllvkbGZQUHBiHdLHI/r
fNxTDzPx6D/+GP8nNOPXCwvlYxxb4pRHB2C+aBLIX6dOKkSGMnhILQeuaQgip8CM4QRKTYtt/bsP
j/CmevzHxTcQLxWBgidq5ucWJIxVrjcaPXKwtdmyavnR/BGOncRlE8FwVWsRNlsrs+Q99XQfuXS+
l9BCqhAnBtjDcG1eaz4Qmni+DUlHDBWNOmQo9y+HSniuk5Oq3Nd7G6AKkSLop5Ohzg3ms707V6UJ
K9ZHhxxo3P79wwAc+EvbLdI7K6TlA/E20YeRHJfQ/ykhqK70U4x+W4rORffQLDP9tGAbLOoSTsLh
QmzzPOt1f4jskcPlx7Q/tX5AMFa+OgGjOK3rqGln+nxdVSK2zWqj1wM5VKq9QZaq3pUOABogHm/5
wJjme3ircbfJ3iSrGSu8qS4+5yxLaz1RGxyyzL/dYkY8cKVDubo7gKg+m1zhzwfKK0Oi4IySMdUh
TUKF84hJF3INAzoQhEqe3jiFY5NPPLll19Ry0wTOFSM/HbvXlQwlTMzeY0YL9NCKOvcreVvbbT77
9SHputRASEWjb4kxNpv32FHtmoXSvmuuW/fbQZcgodvXlhkVe9ncPERGtrgmAExHq6lSUVt5k862
otuysaiv8zH698+MVVN1puDm8P+S3920UY2/7x2D4TOCT20a7oANC+pXopM1Ddk9MMoFj4lOaeD3
cqrBxO8pgijgWpDAebFL1xlI9rECpte95P4NNmpDJoQWdnfaBg0vCwsH4iy2cLzlu8zIhhX4w0hS
BnwWZ2/+d/k4yb8NJTnV0ftfkmg/+2ZFi/9qIol9nHk74HoeBehh762VFb1+wkr9qAVHBIOlzNID
wd7eZh4Ycrkx9UbIWQgUh404HBWpOm6kO/YEFUKFa+FZJjHh/0q7GqbENqlCOTXp0raasfa8lM1v
70vXf45/7lEryVf2kkfOX9KZcY9g3+OTZCiA+Px/M3unMSDIdj/XwmX/0OUt6y4vZr9cJywxW2So
PG2XRpwQkIrdmVqpGtFK8aY30a1wbBjKxArneZKrR+M8waW85By06FE2Y/88dbtDx4oMiH+BGfHf
z6+LuZys1rG4hDLeWP5dBea4q5TkqZGsgVc11n/QJ2mCV96shNclxg7tw5UjsTV31Hq7UuxjXGlB
414uLQVwjjOLT5CZRLTuIEiJb7fpe6lZhYSeC5sD2pBMyNJpAhGVVsjOAaBQhrY60fRCvcCZD/Qg
82ozdPH3EFaNl/Euf9FgPxMjjJUQSoWh8/SCkRyAXnR9qGqBVbO++PsU9WYkd40=
`protect end_protected
