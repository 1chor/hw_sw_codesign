-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ofcWM8WgsUkL7Hg5+PUOFI29qEyk5w3TVjxcuYkxtystmD/xzWYy/ob8YTmZu79I
QyNbXiPNFULH0tQCRKV4Jf/nBawkHio5Zu6GgZC2Sk/qU62DYvxNQxsY8/BJ67q3
4j3ixKu4GJSNsI1checwNEMGlf4AnD8G3dz1dwyacQA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11971)

`protect DATA_BLOCK
dQsayPbRlcXE/bCENAZGMYf1fREDu+Xacf4ltxkUh4X0XBlxxH6U+d5HOdt1R1kc
sTcxjpZ2I5F4R8rzfJoucDETnqBZBGBNShTf/ijnux3BmU0It6FS7748GojFuh2z
LXu79yakcv7xu7jCMRDL6N58XgRaGRhmfW2+7DMTNj4WufRK/SsYpWRq/OrhWVJB
vVYkC6t048o9Pq2M+z85Od250T55qb720E433/bEETLwrnav1eEXXsMlwFrT8IoF
OwlHZnAJsU7abVtiOfjIr58/R2ku01u0hRIm8jIDP3l4+l/3ySscyXI1ZI/n9iUo
DMQqQBSNwRQRaQe50MQXUIuk5lbGHSFO4Aeu4aAcdJPIQ8OWnXranHghmsP2q5vT
98Fvhv51Ac8q5v5vklbbQiprpO/Jn8OPowV3ldh+jNLqHL/bMLbNCDq1Ujti6YnB
TTCNgTOaqIr+LHPdbfaDs11btwTsFvadriuHouV8hvm2dbv09+t5NH+jmJrJ7iFP
Wf7l+SUGPmbUCF/LWN+yWDtOHWi4XV/+isSR75P2S6HQYjVdHLd6TAsvFFeNB42j
vKb/ZgZbsG/ZfgQsULGfJsp91gQFpJzJgINLEaJbccA+2aohaNKVfTvzIsLDYzpY
toBj2pN7xQRsi0Jc/Wanb/fN5t1U4zg8vvgQqWiSm1+jY1f+LSUG35LDlv7OUwxK
p3PkTT27b+94/jZo98lLFlMfCSlpdoPe8joR9eyDqs6HG0mC/zusBd76C2n0p4Xs
atoqCLIVFQKFH6imyzAY78nyQ11FEJykGbfJbi40Xcwr9mBaq8XSZozFgM1PxVYH
IGXMtoXCHyJbxCgivFI4L78VIwUQ4EvAr/Wp3l6aqrhD5xvtY5jgiCIrGjuqUolg
u0dBN326c0CCuNNMYOeBACsCtugqemddg4e6Qpzv6hytsbTjfDoNEEtfslRzN7/d
k6M51I7kBvnJ0kodQpQGqk4bSkDalo9HNbmC89XftfE66zQFCqUMTyxi6Xbk1rA3
oXsdN7QWy1DFNRWA2sVEeGqZ5LM7/FKl0Ac2UEGf/wS1qNLN0KYC42lRc9RqBY0u
i7muCkSMG9hTwER7NDM7AEyQqUmdajMdZiBAFLbFFtbPw/xXh8eW6+zbXaP/J87Y
sDVv4KlHht3mh+Vt3QLdeaVbix53TSJmWsXNnam6+lfwFIPPNmmoxOIxwXpXpYRy
+yBbsYaJCcv0Jfp+H2JnubYwLaL8W3FoTJ7j2sTBUBI1I2BKtpbaIF8xvbxkN7p+
VzSE91zJIDi+bJHMwZ4W+ww8K/OzIghneXXC4yQDtyQokf2eQ2zzN8pkn2euQ7LG
BOx0g4mlIMWEQgvHNCIgwZQio9cKOjSRpFRDZklFl5Vw5xukKgwC5ClU76+blZe5
Lq6pFHPK+eUZ13AWvBLTzp+FLltZxVvlusNebyVSR8iXDD3Ac/vJWV+92t8raIsA
TLZTaD4WHP/4RcanU4LGn1DbikaA5lyg2Ewj9oHEvuAQYRUfz/4AAUPPGR9UKJao
EX7sFOiK2p4ZvGINZzItpBtgMzfwx+wpjlzCd+vMX+JXAdHthRBS8I6jOcxDA112
iuFSsobGRqEY993f3YSAxy0Colj9YEXh5myrlYyNEjaxmSYp5oRQGoRJXe9dSgHE
XkghvkknPct4k50BM68oX8GDd1GaCQ3/jursOdfeMLNdXfrJ5YiO7OZd1nZa/2eP
6cIDXdFQ1PW5HrbON0bTSETFOdOPwkrJ+YrzV2eoPT9Qj6F3Tbi9BF5W04MSPE3j
plu6YRejT/a6lhqVY7y7hLBW6NUQS/BR1NKpzhj/7sZhTfBVLtSk4dCBRiZOtsNQ
L3vQ3W7KyQhsXFaJJNVmgu5eZlXYqnKFWPuQCfh3dunQUProEWNXYz4/c8G9m0aU
ldPu+xJYVX06Xwj785Ja63isUYyiJ96w6dVUtaPRjyDys6Z+20FAvNVF7vmO5oLj
5OJiEUxO0GvsDMfW9PPCbLkygcETJq121NcGkN9UPP+WxeZFD0QYA8RykcuP9OIO
nMlt99ZXt2YF5woc7pGoecJEEr+5y0D6GjBcCl8x0oELz/AtjvI9KJqpqlA8YK4S
2pFSRl3YP3uzebbv3yWkyxG9VD2ynBE54PNIvYAVOf2svkIShR1pLHng3m2IUM4P
fofbQ73PB/U2a9jgaoaCxdR/iazl1/1UMEEq1V4jRLGoT3KJqGPDLyIEE8kEWmAx
/mHi1B7VbAbaQX2ahVdBgvEedJDYjdvhjLjzpWllJFlwPcueMuOXOLgHGU3X8Xgd
wmv87k72OlJDiZO9CFl/KhFXVuq2GZG74q9j8UFe6VUpueu6puXmRj1//qvdRE59
ErTLuJ8n0L3BJUSeEsRPTuB1x+/ukHCT7E6Kt4d+yi6/RNX190tqJ6n9jRWIhbE3
XOF2hOjgffgHyBoAX8Jo3PzxTFbVetv5b6sm5QtygG5lYpTOzrRS6p10p/bV9/GO
zscAyr3ah4Aj0V+9AOCF6bDur8pz3HP+kHNpV2kLyHRoK3F0pGR+QOvzTKXyYfGT
H8VL4t2KkABhOpfJxJzRoMj0ldWUV67YtxQDJp+aU48+x5pWrAI/cwsQc8qYa42H
rgJfOXP/lCPdl9FKPGMKd4mPedD07t7F9POVDCYFmylpULIhHCAMGCIr2Rf+6l4l
308328POPJul9tx9Araq2fkiZ10rVS63O1qf0tyvCevIxI+V8/6Wkj9klL3IreqQ
EhTfu32rHL27fatRROv9UiNVWSm78pTSBmBFRWJja3rOyDNheVKGoWmPf7r2FAaf
mnvLOwq/JEhtEZRn6D4iAIQNMogUou0XdHPcvXvgoJenvCh3SLETiujfZVPwWIoJ
RJ3MKnk84kJSxQBpUYXqXdSLRi8ZBYJrie9HtDsZ8uxFMBJGrbyDym3pjv51y4/v
Qxz8SbZ3P6Z70Zue5kVx2bM7FGjqJnbZS0s9ra1KeevcGgEU4KfRcQieo4OGqBUj
N3xSXb+HH04vbdOlOg3OrP6Q5nMQAofGc/pep/0gml+mSlgKBWfJiBwnBZfeloGg
2FrgE3KbOlv8qt0kWZEYGAPofv+C5Xa4GKSUAUDyjqEK0sU0gUK6kBW3myHPOv0G
KveNcWOEU10OrMVVgUq8kXDcswmdENpqHgEC8Tfu2PVVWP4ViWi/ogmwMgg0Ab28
y+7PFPSQxhj5Kbx4ni5G8VKgvQQ92OQA8W8gsWriPBG7CZKFPQJDxcyeZ/WBgjfj
jcoQ0H222ytqKCtAzN/X/8nQE5xiH89alKBSb5SL3ldReLCebklwTdOMgrOX5gj9
DblFjh0RelcOByOLyaJ2wRceecL2kia3t0nx4Okikxorw4E5WLf2r3KW927f3XTx
qgMO/mF/febIC6V9+49/9rI5vfljJ2wY3s2PYrGprAMcByC+rdp2L9puK8nb9pPy
I1Qiv5RaZbrdLdlhFUeIizR9tHMfxPZD19DL+gQBxuqatlN1bgkRsmpTXY/NP59F
8J1EBwzKOYb5uj58xasTSXODbv/yA3CIXvhTCHtbyj4UcaXPnu/M7WE9NOkFPaYZ
Wv0rJzD6XGOTc+T5pOy1I2bLJ7dnM+HUwgvDn6fzzXtjGuJACO42VcOL4OmM0139
QcCF6JW0SloyFavbooD+Cy3t/lQHj/bSH4446cc570x+/uAtT4vDQS5NTNi6+ZeQ
rd5RebDYJTeuR6fuaUB+0ecwOVxChn3lvYSdqnMGbL+v0yuiFrOZXk1gVOqUJz0e
kAKConTb12gOk6M8MfiW+V8UjegB3GSwpNWsW2aY5uF2NJ/3W7UsiBTa4xeSZo0V
e8/AYBusaSMufZeEul3fk82P4UD+sbklGEAD9qpAxzIVtL4iovj3ZS4kfaPo7hCY
vOPHn5xZwruEuUVGfufESbopWpCBG3HUvkTmewYGuVfbyS+52PvC1DP0AYy+Mpnk
WjwMajCDsOm9wy+oO+bW7F32JGavz6OSp7loSzERflCj5uJFSoVKs0cam1kViAsg
Aqk7mlVWXB6tY/dRobinbpSC22XPw9WNdv6fMigJAWAeBEIrUfvfdjPVzlPv+SOY
jPiegIMzc+hDXZAeaSSMSs959XlQoDekvIduEswD91aDLo+37Ymo/b0/kt772pCq
7T94eFLnjTouwdccw0ctVVAng78SW84igZumouNNwG3cBzBL99xliVlmO/v2IW1R
qak+RIMlEUcA1rCi3NixZLsCG8FGxu68DlIPU7P0KXS5e3TIoUS+HYL3Wm4+byd8
H0rWUMGS5Klj1dTZnZbmccxI+ThtcpXSOl3AnKWj0Zpjq4XNaP9jYd5DpfkNJpka
ARxqcafan5X1requfGA0pZgBFIk/gF8Z8QhHvB+FbtPLQDu7uQwtVa8ZBOwci+4w
YVNVOw7Ua3kGZzHVl8Cmyxw9OpYM/75q9UMJdpWSqC+sE88mjz7NkmcT8sFsvyjs
csM5SqPpAkMTgDHyl+EibI2l5CKGd7QkSfyrBYR1wlPcdLSG4jeVFFmqw2kd61pK
l6PJ5WgzX2fmfRrDo2P1hGzaRINwkMXfETjIe4Qw0ENxylNVMHdr7+eVbS2wH+7E
6Q4rgXSPQpp9scPAYdLybfwk1J6hpb7tfFbxBE64JZQg6hktEWQJ17nhdXKIRe0D
zFpKwrhr7GfJvj2/kIgzuFCLbs2Fbbw4t+EObu5oBoDmgmhZIG0r3AjpHawnfmW9
aYnMaZotM/YH2u6dqVDvSsqHWIvbr7MppTP0hQ1HC1h9mKniswyNiNcwW2z66a+Q
aWntPoNSDS+tzxT2kFPXETF8exOZutp61FzLx/nP2tKj4m7IYik9W2Oam+8k8ZmK
qwFOr5RcxE/fdzm1pjBRmiQX2MZQIbsvU9iGjdBeKdtlFmZls1tdzHnKgLcLopDX
9eZFK+Lbf16b8njcypra7+xEthMiJv8hsWw3AcVp0aeEN/PgQ3l4elHOPtkB/1k6
xUv04VEfOVyMGmhs6N8aVr64thQuXx5bng90wIQ4tmxzK9zDj3+oGMTd0kb2KyGX
XtdoNs54FxNRCjtJXgxdlpWRUndIH7EoWgF4aSlurHmNgRLQyydy4F0LV3z0j7hQ
DWUYGtxabOtqOaUZOO4lXUOZQTLEovAg3L3ajzq2e0vmDWhmnCD1T5sRa+J8t/yK
snLLv3T9UIHxPZwzhLrOFWwJ3/Ob7nnWJLzfDNNYwRGi0tbYejqLfM5/QVcai2I1
1ZC5bREZZZf2MgGWpGRij/YjWaPgfXKQPr15lp9UKgyt2Huk0Q+LEuKuU7JdcUdZ
qEQW7PvzHXX2/C1nyn4kBcjEo/exlLlM9MNJFYD7BJIbCFq6GJNXNWWz7cRXeVL4
+dNyNcgpVSgAaKtGmpmuD3omGq5JCrB9hi6KGMvcjNeNTWMJfJUi/VAM5d8dH+ct
WBFzGStCbm6/WklKbfnSkFSKexhVponVKG7gd9kmz60oivnQ+vU/A+ZBXPyoYRKz
GvOFsOfgy27XBhOcIDN0kEIi1AxSm+GGqz7bFtr1vaVrq6ap7KYfqBT2bGcD6+R9
4o2RyoHQndJ8XJ9gvwTXsyrdlw0d5jTEKl5FVX66BPpYxlRcqYMpgaFnzEfAeAM+
9Ys34CioEx94WJSrg/PP6qACHXtiNeoU+te2V+iNYjpfUiJyF63qp0LzxuiJPgGu
/Wsh72+h12zc4rcIJkN5qgGlFq5a24wbhA7WQUWkeR6SpDz/nfyBnonYm4sS5qJn
0/gMBJketVCkFeLB1ZBddvAE49R7HXZE/YchqueKaV/p1+VU4XsL262XHHhiJCdM
qQojuaYDACz9v1GK6FQPP6zEP+q1tesgmqAbK9h5VMfou4uFi1+KG7gpsHQKyPpU
yIFNYKZRgY9ZF3PfUt20Rc16Tzdn2TRJZhHxFzDZhSGhu1Ok6bDhK12zBVehL08+
+xIPIrC/EeleGtuygR2FhGpyvwjjhtCQaCa9Re9ZBoMQntIg+toRcu51NyNuFmSA
7BzgB/+y+lBS+CsGqWf99yPMdn+8erSZi+hVSRypg5cxn/MaA9YNCR/4MvczEYLC
w/85JHYDMzBnsvbx1GdUWLdH2R5qfLPL5IImQHtZehROulBcz07RcZ1BzzVAjYYt
ptb6kZzetyvipS5OjdWti0jW3kb+5hJy/MmpZCzdyz5TBfOJ9oJoCiUJkcA4voAf
Ul36XcJkHSdJ94n6s4iLrovoShIO1xKSAbSAZjLxdtkfc8aeAaCu8Zoyi8TPPX7W
alXe9vnCGvZuI0/JCEJgKh2gE9SvdbTXCuNose7iirh2V06MQZrou4Qvzwg60d+a
I6Ima5OY1xtoDJMMFdG9tDYpEKkDiYDVgzFAbb0PJjlPBKgMqrFvZTdEqufSUoj2
swVLcSRBJ1jDDZqvpun60Zp4ury+JUgTkdNzJrxRxUp2FK5KptQKj6kMkjQmD/Mg
49BQuOnX+IKCBiqvDMsZwdPOgj0c2yz23wR3p0JIWi9qS6jOau5MGr5kOUDDIv1V
evMVCoZHO1zSMxvHe5ZCV9S1e/Q4PI57gI7LTOMtqKcCs+/Xp6cu/mlVTlMAR4Ne
BEc8pNccG+VkBouNRcO0p/BVvAEJGMtJH+XRoPTTHOmMUKBmcHIgIUvpXyPb/ChJ
vD7C3w68+lmPC58L2s/RbJcTgfjqpVVWPEABePI/vLkhklUxNC+rcFLBciSHCFEs
p4h9KotAJfxAf3Z1LtImy/5m4DK7f7s5bR0XX6pI+yOhkl62bg5NWiHm3c68X/Gq
Ms6l7d7t3YQmJGgDnZ4PlBPC2nOifkzMON85LqY2uTZ5I7DSLbCY7kXbaJLluOKf
UNePCoVPz94f6hiIxPOFrQszPz5gTpj3Uo/DFAZ6v0l/0IsNdABUZ+ndBQPaYCQG
I+eyQNEHlgi0fnqe5JBvbX04R6zANfJr6me/kOz7hr9QRc/BVrclGTbuQvXMDNzO
z/zyzVvVJ151haA2j/gfgtRrwoQ59datlbeNfvsBpy2ViAuNVwnw0Ldx+NHbptfw
ygvPuJGQir90MZhVv3c3X7nUn/5uhhxwXVxPsbVFmJ4SClW1WHBOPbHyGUJBs8x8
Nu69P2Vvl0MhSG+Y0FfNpJ4tVX2bW6OZPhHL+6qa+LFd9TClXQYjQOE979KrsRqp
VEJ7Xq1PA2CnNpTUJ0y0wOjnz3PEg7hMzVqxp94ddewjWhCdQn8cSruEindpVI/J
fqNivWlqD/NwvtsmNyjUinJ0nLhqdtYkDt9d1GIEXpHcdYWIGkGDEqTv550ACEgE
sQ7HScoCV9SANMjR0q/auTJAuSINgLSqSufnhyN+sM6uYMs/WX2osjozKV/Q9C49
tq6hk12x5dDvapkuAEWMP2iovD5XdJPge6EwSknxcxHGeulCXJREBrZwstjQTib/
qP8vQ3w5bB4WwU/JHIxquhpSGdNfDG9nYLv7co5Fhg1Q6MN1JbflfAY6T9yRTzuF
9/Aw5bC/GRb+CgAC1kIHZEejF7cY9JEoSgiHiEl9+9d2YQm1OhNtjdreA8LzaMMU
8go/t6eJbi15f2DlAykJMfsovKUcpnBfpyh+w65KeyfmO+9/uQQjWS1q2smbTTox
HxpkkQdcwPmp062dMIhSRBovjn6jzMdD/G+GyvzYQl+uP1tbJxG/Z4X6Migdz77j
Z6it6vg7pHewUHhc5lYmMVjqnFd2RigE9h2+skYz4wLb8ENzgdDXlX79OrFZ9coF
2RcD+z/KiRDXRnyTcbXBX3nhuFRXwNPz/Cn/9W5j3UuOe7+vLaI1HowuXoKHwwve
8fqV0NeTKY52m6fkF4V+qZ8AsPKVmjQxWGXJYOnS0sQZjUmx8MncYBO7Lcl3kvYS
EbuVUG0Js8hDRmPx0ZK3OzAG+iJZ2/6wIfVpyUHwjkgvXkLZ44eZ1E8FT4ULktsb
11URV/5SBxFTQPg0UHOFo6uK2WyUM2MOWLdjI81WqqS/gTovqoPnpH5jTJbvMqd4
RgzSe60XJuDDinru6/MjtobUR9gAHWuMZMvl2EjNid7OpQdY0iTVSWZlDjJMs7Nu
o4ML7YL8Qx+d7tb1cjeC8INUvH2DCW9QFUAvWL6g3BstDLnRQj2DoRXD8tc/nDG8
FHyCOOCQ/zkSznGPdlEA8JDip22RcG6Z/EU5sN+nUZNr2VsrPWZysjWkM7EnULPe
wkL6I0rxEyNXaUBI7QB6FGm6vYvozlceb8mUzOwB6CXhentDcNUooL9fHUqgFXz1
+fhhE560tAZFJGgQxdk+obZ8hQpbW09G8LeNaEHiHwy90JbkWRPFT1PgbUf5DSK/
kKllyaUOdNtv13qlUv8E1r5GmZX5cDjAc8M5ykBg9eJYABaAdZKFJvQ0wVaRpl78
2JF1HvuBDMx0jMWADCkS9Y2b6Hth8IZwIAmV+seXRBR1UhPZd6BGCNVHM47HOFt/
q+TGVfgLYC0wfaFJ4Tx05avIJLdL/mXu5bFiwTuOr0KfGZC8GBurYYiIIx3mNO7n
hGmNlhCngtbyGPxXaBUCcT/q81R8H4yWKhQ9u+tAl5v+2kE8p1aj27Qy14QY7658
X2kU6id9wL2YplvHFyS22i5tli3fMbCDwsMfa3+RAXm3FPZ1EZ13KLIf35o44F0u
UDo5kD4VLQTOkbGNi1IPdV2BOL4JyUjll6ZJppOLp7QZam4g4Br6Dk3l4ulV7Y76
SBcbULRNZ5HDp/c1oBz5C/J7bH/muV85fc1degJYMW85PofFMLc6BC8t2frn9pgv
jRAE2jn4PcDv8RvwzXSw8j1Qgmdc4kxG/WvxLk7a1d3jmKa7bmfp0ptgIm+Uww1o
J/2NxhaPsOxoxMkCFUyWWbPX//Wv/Qw9/BK9QiY79mqwqMIbM4g63TL3iFXILY5I
K+iNC6THDCNL1twiSxyz6ms512wdGQCnWPYPh/eqnQ8U2pU8Sp/xakzYlkA5rHhP
BEwtZDs+HBzBCFBhYdQkMKnSjpjVxRHWIfYBSnpONpZctZpnwXFtcfuNFbIam9je
X63m1LUfh1C0OD9SX5q9IZDVrp/QpKekHt1bVd9i6YURT+VqCSRyI4ZIWLkirzhf
vGXwl9f++jwCeb9f6icyhB07dtVZIQlQvk8tDhc0hMDxec/KmA3Yto72wyA263x5
+z/I8S/XDyZLM+R7ISPqkQagkhLyxL4K81wdB5b6qoAbnC4f/NO3M+6VMI8/N4/n
TgwXLPFZ2elfxpiK7sHcY9iAeWd3Mtzk6p5DoleD9HDkHTUGTfHbNlpYkBfydRac
47QQUtetgUY82hM/kZaCWzK2y1lCuX8hSbEFocoFvCXBHblEwpnG68tPAGlakvHv
dIoTUVbbGCQf2vVhP8Gbx6lLN5PPsMJhu+Ey9eZjFJJObm1vzjCny+yj7hWPpa2v
iss8NXnCB2w4x7M8TNFmw6Aeaq2lr3V/8/p7947w2kKkAzhK8CxF9L8x6FaBLVXX
oFQif2wN+o8GfghGWzKbjiw4Ww8B2pcltt8dGdHEE56BVRY/YqVGS2H2vY2wzYhI
paEIZIjaPKTkRqoKmq06Tb/FobtrHqxoDJfVm1lPHKG5kWflVrShHCxK6ucX6NHR
W8Qg2y7IcWP/JtrVuepldnBiFfa4pjl/QSG0/wtdVrTUrEWPUCj6SLvfbYlDvuSF
qTvJaGdufH4l/jaCL9KerRVwF56TPJMEbMMZYui4ngBzhN6lSgyUnCdmNWtaDtsf
36lkP/siBsMNgDdOEamAP2/EJNXfyQD7SAlPJ5BtftLvmewTo9Dpj5P1JFPfgbWb
viMw62+pyi+3UIcMpu4QyjKeQDtMQsjiXsJfRPzHHt2aMbZxR2lvIE+YuMknYF9h
u3PmefMLZgzli1wf4C238SuK4zz5UYg0KfR7bUYemgMzB7JPGT0SuUoFh1xPBacw
sVl1pGaqrK/nDU21Iik/7X9xXRZr22Ny1AZCP0isLvB99xLYlEIlW+jUShV/ffxh
+jak42Augx5UfH9AcbhEYjhMOLkrc4B8fE5lw9+zWwM0w4EkAVAj/6naBqxQJSRQ
006h8SOGbP1adbw+k2ZQMwA+q/N9O8sY5XOHpZvkiHWfCJZGeThcVxnI6QFVq82o
PSJ7lUGAuOAgCRBe1nGuLE2+IGAcpTMG3/cu8o9fLHMrR4PuMu5UuGu4uNTYaK6S
BL0ibKx46bEKXUBGefWEb7kTU2tXf+uf5GHbVdjUKpO87lGd2fFp3caxtWMWnFkU
hhfTf8tYVIaiANU/wpLXU/ExdttG+3b7TpZOwWM2wDFOSTD2oBSJlR6lknFAwmQ9
G4Ryhqwfgfy41GJsISRAPkm8gzf0kcYE4iz+uQX/GWjZZiq9JyDkzAr9OqZZ46kd
c+K4InyNYmpYdoAuTjcVooMRSsGX+vD/itJ6df7AsjUGm781byNruwuIBPfTMGJ9
cq4U82wkxIKqZUK0Wbl+RKhR4WDdJkMJYX877uW3pmSrUgT8oyY+MgOTaZA+Jv+/
3R4LPYZjUAC7HuQnq9js/OmaKbNsewCMP0w3YLr3Kk3N5e1TuAPtQUqiMLWsvmg2
H7419rugRwze6xOUR1rEf8YM6zMl3ZG7JjoN20e6Zso6vaj6DDrctnRedqTS+/pc
FwKA6Z59LPkofSEzB06ohY4EeUliF0kvxZ4pyN15/uzCUo3Ogw2awbfz1yb7Uc+B
bk3zbNC5ypRBTbhviRQaSSgxH9j6wiwIbZZcka7ps4zcMWOAA5T11g8VteHkdEBg
OMc6tAejZ3cpca623uI58ikwlEP5jcSSO83Be9un4Sdimda9xhBhG78yMkMrbkqt
tPOL9z71AuyDM8kuQshvLgydsYgRbOI6n0y4F+ehK3j3IeOmFBrquwbh6rgSPf/U
QlS+6Ad3NJGlGKywdEsCxTP7tplq8ZwQw02Bz+TlYeqFec16r1nCJtf+JwoMwzJy
oFwz465qyvMeLq6mQqda7OvrtjP7nZ3nrkrrS78pQAVzDDtV9lRBTUe5uXYpW6/q
cGlyfbVxieIPE4UesQn2nj7VPAOxiHMYbwPoDCP2CHHabdLPrEZdJNvNQLVBcMQC
U5Pe0mygS/7jeR9LXD7lcXtvXbktw9h0FVotvsHoIYabuHJvvqljoNNYzgCYtbLt
ZSEsoyqccPPX7KxOa8im7sLwx4vjnO/I977ZLWntZiLcFOfxIhDt/sppbS8UN8zh
a1ZWXrX/Zzd1qX7gOfxXDRFtcxjT2bnyWYYIBDxPQRA6vtescDmo4d6cdl+FQSFH
vUYiJ0qkbwSFLl0tWVfHaSpSy7WejGl1lbamDbNTOg/eWzH/jHHMyvv6n/5VPlpF
qe44i590fZyerp2m7n4aWEzMk2P8nF1dg6ssIZn0UMMTAjwxbInJ3xKgT65oaHPg
Ci3JoFVPXhl5SsVjjlLM9iSI5jC/3XuyPmEXWsjweL0gcC8hdcZME+BjFc05V6ky
GJr82BDv0Kiv9yXJ6/mXsLGFKbceT5yJn3p8jOTxX47V+/DiywbT27t+ziBE2KcR
0T7fsKZJIjueL/5E+b1NIg7qrkg+xyQ5T2z5MY0PDdsO+zXJ8CCCDKew8RyU9hU6
neGBZZlExxdZXLLou6q0On2FC66cTlABaGU5nzfRRqsm1Xz8h+qoDwbJ8YLhSrgy
Jo4Czxd6eTEkIcJianmMGqBJHBaV2BgCYcagylAfdDUZIXUHQdLASiHcv0Y9e1zD
c/vpGGHW1C1boODqKXgAzR+HfIDlAoFZZYXtuPCtQJDl9WYFVDSF9CgSBRLxFrgg
DohOqCae6f0QXxzO7NqRGQtX/EV07sIdH/dGYbtqb3yFOo4fLlhL5vxEIL81BJPK
a2PWvpNi/zHNeoeacOEatnsp0syvSlkwEf5uR5zdK05vyJTjV0l9W+xnGgFuEug3
waGjAryx3HCiOt1JdKEeTF4tNME0NElAcTplbh/1wh2OH1ExiPTn+7GkVyTz8VJZ
HSvPVo3YUy/y0YOblrrM53XKhM40yo+sR87wdyw7prqRJXrW+Wu5la9Gm5ZrjztZ
uI7vABKBfyYAuGZeHYMGLgZmN7Js572pxT0P15zzgfygJVGE6uVgj+nfipXhgsLh
K6BVGaRJKIQjvdwuwGtwf2+yLqQm8hkPopGy/axKK3AxLzzjbhcpk9CHuwKWZAZF
ecsAIaJiYTJdVawypDkbsSnpsyExjJ9vElg2P2kUQc39tk91SuULIujFnkq4zf1o
WXWRZQzWALS8RCqGx+Hra56R7qvnXogVv4z43qyU+KPk1H6cMF1BOeou2EmBE3i6
a26Lk4rYSp2q3avfd8WE+MYm6ozgebBNwkUCs2hRAFKPcI2rKjxiB730fo9f9d9+
Xg9kVNASu3MooB5wHNy1P9cdZw5CPI1ocfJG7ngZBgHp/+UyMD9Te/PoqroVRXPU
ZIh6kDoutr2r0yr+ZeGFQyVauwXbowhXhWdrZUJ12jE+7g8Kd5SdoAnOK7eeSoJD
UDwiJAlSxBA+Mvv5rSwJZgSox2dJ8Yq6pFAbTwl0HC6vcuyx6H9FZ1/3cl72CjXc
4l4fDeRNwhgR9cZTnO4sJW+RVa4AQS12JAcTUsZqArCN5ys0FfrqmbfRBOaQ2p6C
yOTf2cofoM4ypqWZv9kd3v2owo4fFYdGk8DfL+Cy2pOwfIZbi658V96CkNAXckCU
SjWSgnI+CEXKOEj2BTGj/lbd3+CjuDgYNnaCVeQFD0ais6lHbgBmpzxTCvVcfP40
EHjRxrOf2d3FqxQY+BiDX1K5o3dJqYlUmSsGGhRw65gwiexxvNUceKPRmE9XeX6o
6PYaJnMsLRb1nFreoVDgimyvvnByi0Gew5tDzLrY8pNHsP8Zuj8Aqj7jaGJO+6NP
0XCHRau/qlj2ZwDlq5DjhX/idLbxtDc+HjiGbvWvS8CvvvTsqG+ve3sDn68kdhD9
z+n9/B5vz8QKYt+VpC1hcJ2urQipDNv/pnYMi/z8SEhBU6BqY5xjeTtYlUvzGUS7
m29e1HjJjAg5j1v0BRm6/1pfXVjz9vXYNXxjv9Sno9JjoWEjaoZPhxJqqbc+93e5
ofLg1jaj44GqIt4f+PHXHQl9VSvOxAJH3RWuEtuW+3B8w/UPZZtVi8thCtW6aNeZ
g1dlx0xicHybWQE0ul7fSjEdsv+qiyvl8H1Djx+KxUEm/9Sb3mG74Ekcq5L0m3An
VRGRMF1Et3cWOiw5/jFx2eMnnM3O7/FKTv7MaUOPwqMYQZbZ+8in264QMddD422L
AG4xTTvPC2KLB+SK2PhQMzcr+3oAUBdmIrLyiGMeP+u10C1O9k7dUjl9rygJDYiy
fH/Rgmq+p0TrUw6VZFEmDSwF5+BA4wI7MhMAvSeFL6NqDCtmjU6d+H1Kuk37ggVa
quLYpRnkVH0vCn5sKNUrgYKpG2oNyUoe1bX/74oz4tjIyugzvzGg78Hbh+kPP5wN
upNv/b4cfiW94sCrIbCsuTap4003QuoWAv8ZT6+hkmr+aSsdAef1HJdC5f7r//B2
KCJFHVtOhzPU66/Ar5mZEfNY80kZw1WShosW0/uO/v+zROo/Ov5UhioyxUSJjbw6
M77bQxmOL6jY3XaY9poD7NjWmCASr/wkjrI1TG6cN0hiqiVep63gsVI+lbod9YWv
yJpQgMn90eXwYRt7nrHsRYoUt6EbTk29GTq6gh2ywgj/8Cj/w09ob4ksUjlHgzBf
F0oxhX4p7gMZMHqxcrraLN+oVweaSNywxXbwfx/iYX5nom2AlndJzOX+r4dCsR5Z
2wa6u7qPC5TB0ienBFkA9a6uIFWFo4Pw20qXFLOVW0+ITO72K/9IcHWXqyIhG8c0
V9KZI5U69HPLn9ipGVKm5EzojHOL9c9hVVNIQ7onoSc4qwyLEU57gQRmqPEQgyD2
H+jb+SPuabWGpepMTOavPUebInrwsma1elynjMfsw5FeLOJMxlBxBMXzr2/w21bF
N4ljCVpyItN6m1jDQ3OHyUEnPZfF1KZgJaqokyGcpGItVA15hCt9neY4rzqLQorq
OG0ph69GQPi4RWArz9FIcG7o5yYwW36DOjfT5mnFNP7ekSy5fG9D/mSI4Cnl+pLm
0x+Quo13wndKm+xcx/pQ6cfqWboEk5PbRBE2s0YPvLCT01fQCUArIuN9DbZ0gjzq
kXa+MRrmc1/8xKC8FOU2ZB75rBkAW8ib8OZwYZvhXAQ6mLUGPe8Grac9aXvSLzMp
WrL1HcL+i57ooYAEqyQ6Mpceuj/DxRasLNssz5ngWjf4bVjSEEimqLYQgj/xTPY/
OVFgItww01eJABrF9WplP5wMGD+1hJ/XhaqYBiKRkm+LzHRsuAohFxLyILRwXm3X
EGbeNX2n8JB/h4Gi4ZTuKrohWVSQBUqeMF6TttxlUn0PRzyKz5jsFQbUSllls3Z9
hMjgagZ8ORNiUZuUKxX18hIUs6s9P25sKCvXKjSEeb3NTfEeaAbmLKkmN45kLBVS
jw3v5tv0O9v8uNgcJDPaUdEnPKDa9Y+STini0jzSRS/+wiSALNxgL3duOIBFqzFT
MDxuJeLXUSZrgJfJyjY81ywoy1XbVCgNGNcA2zU1xS05OSWlCcYszbi3ZdJ7n4rw
41otXTpLVcEEH4h44XZR38pKFKNZLROSVkT0wS9zp50RIkeQ6tkYl0v5hxY/Dadn
Az/3qzCyGE8u5UExs5lOxdI7Tq0gwfsCqTJMswhItEuvIQgICZqJzXafz2JvGNHS
jRk78++wPcKFQYlwFSd+GVPw1lXuZDLMzK/vBY4LHi43hM1WIbbK3Qk/k/jKOEOE
0emWEILEJpdU3iZ68kbRwl3p6GYjtbtCkRDcNohBbIyv+3nExRE/ya3qrmPW+AhA
Kl5GLt5Tzg9i/D8b1soFQ3nXk0++1Gik9+oEdwbE90mbhUfCLLJ26Fmd9TD5MhGD
WL+rR7Uk74zRpWsp7YRTMSi1UNK6fVGYvHqbGEKYPGZAfHu1vfJWNirUuv853Pfb
g2PybJyneQ4TNPlaNSNDJjSpzqYvtOfmYX1AgKU1oB6Tp+GRbOkOo5moTRUH09y+
oTqPijj3ffTFhcwOB3bLPy74Vl1RduNB22X0GPRAp5FgHOaUnZdEkM9jX3ECvjnQ
+dRubSLHn2KSrnnl/CK6nGb3FBOoWWtUxRc00ovVYAN4A8V8IMrZaWs7uCVY4/Q6
if917HhsiRdXoPvRTOKw+RPPtqE2+A/uTDP+R9xqeJCj2W0pGIt/EYbndIQw57N2
3GmcX8KCLcyj1BrepbMCVd+U/HKIjQ76cK911UBVCvGPVHHhwSbzLDTM2BW3yxRn
eGXmafnrgUe5T5npzLbF5uvbFF1taOL5qeCo0z/mWXYvvqyfbU7FRwsqO3TYZwEC
nET3VI+QuZndyNSfwukxAjl3y94T9/mLQIaWXRd4rbidoAvSux4RPNRjy31q0cRY
qPGL6JjaD7RUa9VqZePk6ezY3QxX7xxyVPS6bMyizuRA4AM2PWZgcAcsQY5ON1nL
vyPZxk40uPALwZiw+aGKsA3dA4CSz97LsDdQwoqgq+tWgPvbER3r+EdU9u0u0Gd7
EDz4uhB0f/HKFCgeVPjWBNURw1E4gfkA3Qa0+1zKjiFZuiHB8JtOhGNV+Ex1NIc1
zRZKwjUCblHG2U5kFvy/7OU41hPLiAOu68cPvwQPRhcKZbkw8snIAUb9lFGrSEQe
iWIHKVmuhD/YHJMx486grR1sBD+/YD7A85+Fn7V9A7vMQLSiJHO88cTr5HDDJSxj
V/K9hCluzmKdl67oyXtj6fReGf2sTH3UOpNHLqE+muf357e0jWBzoG3VWIYQ8B/J
SB6YfbKLS3pRIB8yDrvYZtMLOOptzF0PA+Ei/RWrawl/83qdLwLYFDcTR8otQN9H
g9J/48REnQCNtlPjMRUqd5FoTcwY4wjVlQ+oiE8tq4NxMYlkkKuNOxdG324dP00t
YbbnA6L52qIb0g+wkr1VziknzHnQzbOR0savYkWFhfUYP4pnUBU/twrdMd+naIl0
`protect END_PROTECTED