-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gvuFW5WYeDcyF+07mfjZzGZsS1Jx+J3zr6uAp1Petl9usRxrH3pQdkDrAedAD7LM/NNFwQU5VFF6
AuMCVKVEUT/DczgRYbjIePYb7M9YmUvAmtUQEArWiedbPNu9ufWAPy8T6AR/FBcA7Z1RXVkjDlQM
m4VRJ6GB1TVvGA4N+qGkjhwWCMKDgzb2BmX7mT3Z8VWC7npTVC/d2HA72irAkArX6ryB//8r9uei
TWyS7TCCtWzmW/eVWn58sG1zHCbZit/qUsTHd1hrbiuMZDCatjJqyc9JzdfvNp6/t7lGoL3GoulD
ehtRw1hGf6VE6E7PXyUw/xODFldDUIQfTk73PA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 98352)
`protect data_block
d0ukRLwfZFq98Lp3ijZ+9yeUNMttIOQ4kR0+ZUnRfP4i787tx2X1TJVIxQpETRq1l7LvgJUmQ6Ij
g1SgSxebp/hZbpDyXMr34YixEyvjHoxZPfkTACH7RcjIOLB/fGHL0Q23raS5Srx5ZURpAtPFl7hW
nqtbhTBOLKaCzdelUWw9I+zTG+pSR4c3U5L/4vAmdeXsAoikGa/s87as+TSyhxRkBFHA/iTdpogg
GYoWIqyzaI7kskQaYOxknWk2dif8Uo7Ubc3FOy8ei+QXsYYuMdNQpZ9nnBbtKxyBJqXNyWC1Q1Rd
xR/1vCh8ze9px7Nqa9SzvlCf8f/DNBll5d6pJ8H7aB/PheUSKWaJ94i8JLeiuqlNWYHFShtRZPZR
TCaF/O58Zsz+/YXJ2rDglCD4LrZYTypEbPyFWwls8UvkRHM7do8lQMbRhNYF+OkB/yc96iIonZWx
FnNrXufBj8LEnIlgfA2b6PBUKSUJNRcTn/NYNbPN0v6JL4ah+ltNWb1MqwZEJIkxaXE4M9GxB0DN
l0IgdGOEH+9zmfzuBZkCg/Z+gXVuvkPAXtWHnXHc4tSmrfwcTIVeMjO+SmQjR1MhITorNm+K05Y+
62cwfIAA8m4eEeLXvqgcmXs45J8ZGaR7ZoIIis3ETJuVV6gWYrhOfjbqorYTHf47q+q+Xen/nuyG
FeIYzfPWSXkSN8XzN5ggYiHk46qyu0AS5Kla0FQZk0+z3zRGH7jPNGFVtfckbseuwP79d/YFZ9Qv
2xhZkR502zPXlx6gyrkhWqcB8rEmauSYlMQ7ZSjux3q7M2m8G2WcZOTBqkD5AjzVXMcD/H5WxT0d
IrQjFWH7bdHQdttyzt0iqMgp2YWi1bTNfq7a48KT4ge1DZXET5/6Z45c9tgNpCPZc0WavEGo8NlP
PgaxxCNgaa1TH3PEfyUmmWw6jQ+3i2ESII6m4g98wKXHJe5a78SW504nfD9OOoPCJMyC37mU/gU6
ewzOWNoEZGbLJRBzAjwDjXEswyXnHNKt6DFRFHBSAUBtbYQJcpXLRPkc0gLdzP8B9230igelOHGo
Q4pL5hNw6Zea3GM7uoqpgagIAIEcHirpcht1JZwNXW30//UPeHTE4WlT48EScz6wDBkWoJxOcGN9
BNxGodHugM8t8tUjbSiJuJaJQ9R0yclJxHbZGiibOvQn7UIpGMVPo4Fl6G3HOH7Nd6Gq/a76AZTP
vPIbUaf+xAVt2Q/PuYyUN4jTP+YdX3MOawYE8O2zSoewgBY0dHvRe4TvXa37o9WB9AqW1U2HBPSC
rROjQvIf6mL/AS+ZeK7BfaM3Prar+SDlPhivDSfXYHObp9Bt6lMGNpq0YhVc7P7Ac0LBwTqYQTIu
PMcmfE/0w2uX2ZfJ0eHclYoOEWNxbeRjZ49C+8+7UC/3d4JmPzvqmLkHE1mJWyIbAUCvVVbiRd7O
oEQBKTgud9YbfuZYalP4GxRywoyGh6tTVUGHUj5l+BU+66UjtVtAPdUfM9plee6OtDuT4CZT8Xjv
m9/gPXrx2FmMeXpN2zkgvct9MYZOqruDfPShEYqY1iLtR0WREh3ZFTctZTvxD/yq2iYgIeMMtJ7O
I87C2pueP9V4E2uyGGLNpBdqu8XFPLCHNTzeVLCejmOZDny/0BiRw/0FCZGpH4SMqzMJqERC6tFc
lcwtn8n9sYK2Hn3vKiHdnds6YBrtjXSGw9PgUCv3YkQnH8sJNPpa2QP7kOF8AVVMk71c1QlUnTGd
3jp8zPRmO+I5dQUE8hCJKBXzkp0pyfXfu1lnnhqpUWzikj/mkyOfvsf3gW2BFlDoGY4ItewsuTCh
lU6CR3x4dtBXtPWqHgxufKdu+t2ErNdd/cxzpiFk0VylDXbqv7BG7h1cJfRFbZVPAn6eqmFWe906
IvQyra7/Ih6GWB3DsQAHleB195P7Igw2+YYS2WVyf4EyyrffYr4M1uYBEso8dtUsTykvyP4EYFUT
8kOrx7OIGkpXpZn9LrMTlb8Jn8WhxoxiR3jrodgSroctomnAHjzm/timrzYBi4fX3RzehkvNT5ic
O4FwYXdYszRib6SHfblMUrak/h+1NC9kTVnVG8SQrAwq9mgsiHg7w7wWISIIBYUY4FUyq80ObQds
V/HqxT0Lpe8SIy+XrfZ2fpXcnM7o9lKpnwJ6EtShnTRPD7Iz7uoJZ2Kx7D3qdbg5GFnKk3+x2BPr
n+qcR+B4kz4pfaHInDPpK/lg0xBXxyG/iDgQ6riPRqPtm0k5aaTnFE6Autz27rvuI9avas4HV7v/
mpiaW1AW8WEB1PEkQuQzlnI5eXvTX2tD5VGIp55dwuxo8XoUOhpHVgzFYDXtqy37QRJp5Zuypsqa
wE0IxXe8jl1wqP7LHG0bRl4crOm773hrXup2m+qVo+J1IqqqLQbS7RwnKOKIMOQPB46ACOg5GdsT
lTv5mz30VUCKf9/X6/m1ltk0TzaeNoAW/zeV6Pbodte1RGDet8jjW98PoafaH2dgOekZbict5G22
NQ1HSNt1U0+qo+vbmwGNlJZGo6TRqPpp/cbLQIx7uk1CZI+HQxJ1uH5rWqBbYYu+0y5ytsjMGjsj
/d1LGejdptQqo88K+HkR7RuWTLuqT4nBmPsz6sPjAosoor+jJHKQPayvd6FA74HcFqCCTBx/epK1
Lc6eEUbRqe2grpEJoh6B0xx1YUa3g90fp5yQba9fcZGMWln+b2gB8mb2ZSMxr0YxkRsoqwdqn6WX
E7MVAzMp8ql1b6K78f1BVhA6UwL3dod/XZWR+yxOGrejSMOx1GX/9uAinEkivM30ISVM/I3IYl8M
Il+zQaNZ/4naoDx6ctt30RmVV50yjr6yM2BCIvvYwR875AGYYI3+FUgtfncqj3yUMyHjNlVdH4UX
9Et1EAKomylRKGuDjIAWB4BrkGeBIaQl8o82ngiNxz+Um3EVwSxyMEPK/WK57KQf3UdC1Y77EShp
2UexxL8ZNM4axLlk/p5pF7+6kH91xf3IEkqo1Xvdz1NpD8kxzUGtUwUEnXNNJhhOkBqySSGlzcPX
RJ/T7E1z+E9YE91KaEcIO6n68PoUNjnn2CCwkB4kiRV9W3F+xOIeXRXnov3Jq0U3O9UzmWiQd2QI
Okvl60zk+EUKGxeNiiICG3/3+4AjjS1JuCja9clun54aA32u0+uxRno+67UYmcew8/hQxUaOt32F
EHIq8vG5+P22yaepr8/xNZg26Jmeo02nxiLnV/3Zb/MRa0PgdtaG/Lm7YoTrZSlTyHGk/pPkizfg
pnbp23IKMZQSG+x8g3nYGeapKaJZqAOpmaT/H1MjjrIX3Ts0Yru5QFp9Vrhf7X0BP4JKR3fbCi+p
JovhWg5i5IXkkvHgvmAblohRvnCHp33zGh72FeHR1SuJW6U7RBWvpE/89Oc/2BK7ofajEsy//pKC
ixseMG9eVhm+APyJKM2da+maeJPoyOYolZgUOGMWznkccZ7jDVb/cf1N8gIQORmOpeftzocmw94e
jDP9hk8m/xZGuDvFKL0j/UnIl8vvx4JuLEb25FM5LP5AOpTDmDuLNnbQbL6d0HfWijVtN8KuyvWx
ej5XtL6Ju+Nr7nf3Kr1lQC7DyvToW44otRAcf8IbwZBK0cfOlSc0f3lxSzMAowZ4W+pchthn2JkX
8upiNyrzb1lzNGYdsmEKg2YY5WzTv+w1OzBWT2rS1RsvVDfu/XktfSXhYIASfcWrDzT3HcfBVxO4
cKWWvEoGuUpNzAWebzBFVFfvzKpq8N3UgR3qBtr4/uJiEiwVaMssD1JvkCY10OJGG1cZNQ16zAqG
h0xvp0gnMsKsaHke3s2roRZje9HD5JlvZmjzMiuwuT1naNDuV3ZEbalZGSZeHZlc4MgampsRy9OG
SH14IR+zcIkYROHm+H1cwXPvxbLXeq4xz3F8qdoollWZzuQ7SV7QBcUwKqvMEgve6T4v+dgQXLL/
lMbjoTNJus5B8ON5y4lqDRwg/7Awj25Ou+iTaRjGyBtKFpA/RIT8JuwTUpcm8lFpmQR/PsPe0dTj
OCS0yy89S1SBKOscyodfoU0yXd9wOzDIB22/Au8i5azguBsz5rD0I/WVFLNGncDMdOkmH7h/ne7Y
c3JAP2RQ3lhlRG9CNyrBjpqO4sUBMSpg4JAE3YbjyDlyIdw0hNgRunaTzREmyy1RlwB9kukweVWI
swIM2troNAM8ti7RYe04e395PWMuBkAGlg+TmY7d+CI8SKoKerC2zswMRpqjfQqg5K082BuVTFgL
54mqEmhmIQQz70+k1J33iytRsXQb65i5/V3qBYj81HV201ppCRr7wMoV4tLK1v3vWw0yJntG+VwQ
Uqp3YtGPDMHkayaCleRLYc8AptNbAH254UtjsOm7C4CtaCa2Lv+4ywQ9wFQIvkTycBwRwhAJMWME
nVEMGSR74cpQO8ksT3ttjjv/fKsfhBLisYfuS5EsZ2D4HpmmaMnFXpyp5hTpe1uiOQ2RdQNjxGSD
zkBqei6rEWMVrsZUfiHEdTP8B6rtGo4bu4v/TAuyWDAIpYrVz6nt3GArc+CD9zpa05kjCCB9dwdp
lOWa6e8fJt9i+G+Twl00bpf8Z4hR9/GZpL4S3T/kv3S7L9oOBAN/AP8AaZytqEE4U5fslesXawvH
DvXGIcgk0T7alg6U79UWp6afZaB/2o5+qwAPDkVyknYJs9twbKJhFDWhbkRlXG+06+YvCMte0Mde
Qv3/x+8hUARG4dOHv6zuHLPL117b2XqVAF0AGnd8qi0a71bp6d6Yd6y0knj4y0ESu22YAZoEE+Id
wXR0wgadnI3RL79jRfjtc9Kslpb6VJTu5Y6ll4fImXFA7JV6qkoeR7JSt+PsKtWBz2FAX3vpBo98
VU4MoAqRdjXahqhB75VceOQTOWl/42eraLXsp45YR0pPxkRicNUr7no6BmdjRI+v2A+NeStVSWyF
NMwtGn6FCqKoJOqNAO5pFymTO4FtygZTm3FVGEvnvr7J/KtjKfRU2jAB9T3NU5dpTgcCQWMHjSJ9
Ii2QcnGpmnypFNzirRoPhejRVKtdd7TyfD8UoDo4d6qVgNN7DWmFl7yj3Cgk8juEB3MYGOalmJQ4
51aU6GrNtHM4AkX2i/e8O0GoqWQUjk4aIu5sCxHX77OlZdUWUkGZqjDs+RmH9aVZcgvjNNXLoFHo
1IDsjCBHxnx8LF68j5Jpsei3mjQOqQYn9SGtcQyteyQia30ULMqSLmnK2Ci/9XiflhZHxu9QdH8s
+nU6pUh/9IEGMlPYxSd/vEThtKwkuJIq+QBU7L/Sm040KTWivKsXe+ZrBq6yp2QFRMQ0J0DGYD0w
/67pz+vO0DC96D6wFWuuIA99dKCU8Qd1NSv8w1N6Oifi3kGTlMw5sKHiOtw3dLxS+O73LrJrCkaC
Ip4YgZiKdC1QsRJz4V5LacHwzrJV3OgmVLx03aOhJJOg9KCv0GlB7sXKLFwjkTm81RLCdmCzzuhN
xXMwtb1aLKgc3F7D8+LfnYp225S8CVMr4Yho8cGN2/U7nJgVZ5BzBut1haeccJygmft+HsrjWsgX
NV5+ofLPGrvQfIpflFeeAiMhFzXIOeAeEgpyNk2MmOt3si5ubZ+LunYUu8IRs20JNVn//CwlP16B
yfccldznngD4MGyb1RTbZ+7LA8Ina8prR1vCuArfI8z0BJ70/wXMQNT/nN/BI2MkhDRZ+pQxE1th
hyek9i+4vcg0RKDlDmo1efcOO66y25AwUinaY3Gnw28tUmTE2rt/igHfRn/VoKZRAxo8dy1d6piQ
DS4B41qCi6k7wDFYEp1rY639s/kDxlSTn25kYQRTwvVG/t52tyKWHsJ2erD4ZKodxDHlmMpc4CzX
f+VMe7Ot5GFvoAGFeoxnJUn4NdlZBOGlNXMHZoyn5aXZXevpTp6EBojVDluLNz/xilyYLet3HQIj
yIKJ6vObcRhtexWm3c4qW4vWbfFiuYB5X1QdadMorfpfv7jnFzNcyFw06ZUQQKtIIwgCjgmVbZtI
j9hES+K/ZeICOyvZWb8Dztd9ON3/xwJn26tO+aXps0gZN1KEbZTRkMh0GQg1ZhSBEMNxD+LSsSFx
79ARJQC3BGuSH/0dhpcIEQtubHxalXUdu01xwD0YuvR6VpuWcOvUcbabdKbg8lzavHBK37ZxEWlK
6tV33MWAhVB43TtWGYnJ93FkSdqeah9OIaFZycus8CFjSAlLppBC2Pki96JC6DETpK/Y54x65H7g
66bfFsqFRzfqtQBVtIjsyPcu+FHojV42iz4Iutf7HnJY4Z0+f1Gao3eJBWaUR+VGZSFhF48uXWtw
5hW0y+H0oRIc645+3S4GbunERqseAiRdDe9Ls57az4Tx84GgRu9GxPto8AtBVUnPR/1Rwe7HV0WG
Gl7M8DIhW3lSpWxgM+Qmhe7I+IAT7D48EAHBoWd7qdEUZxwkrx3kdNoSuV9lgacVTvlTLewKImA4
24OAS/tyqc6FXlBYoJqyXbvX6f3N9HqCQFuVNbQl+UDaeGrVjN9LuNtf7ujy/K9RyKJKKqVyKpqZ
aB/ore+xzmpddhHCJvD3itlseXBVGY8Qrjo2duzhLXBjIlY603NXaYLJkP/8NT0RjcbUnL8l85qn
DskwdiQn2JTqFW1VbRRRT+caQrngswUynRVbJUhoZDWGUALg3XuRoKoywWWXw4Z4RzYFiyxmzt2n
5LDMfnRaotMBTO6mPa6RrKJ/YMHXulnxtf6DfnVi5NsCCMXZAqp6mcSmaEaO6NjP9Xf4NTczu/Jf
vJjzsBN+9jYbZUSh1E74mTc+1UWgy+pGYUaSp3Xs6ixLxbJ2OpBOf20AdjQkjKugef6S60OtkOBP
fP8pTy0F/HdX5TYTL20gRYV4gRecROFdBNoxMb3jyFm2H9W6ZmUWilq28iN+52jplQRyhgmN50LA
nluJkJafF5fPs2RohM1ZjzsVWR7z24cFl7/YBAV3BVr1wWR6c6Bq7g4mdanck6M2McSa0DcpbrsJ
Hl/BL78XFJbS8Q/zDVzpKlPGE7pAeOdNa8CisP3K2yUYJYF7q8k9sOg/KrXCoxWnTQDYdFHLyFLl
2OoHwx49EE4m4WaJMDJGknbKTXctO43R2qi2OY1mF62cl2CuqyQo2CL6t+74NEaXB9VWT/uaOp1f
Rff5NbI13GMaQeDJc10b0w2fmib5M94g+5wiw4MqgpajA2pb4GRy1xxB4qFj0ZzyYvWsN79gQDeE
QHlMmHCewSW5TXMNboI8/EroCyHApdHELst0g1Qdj/Gu3YLCv6yTPuhaC4VUY9VFGLF+5OnCBuHO
qVA8+cGk/2HwhTUqw+X8dsaXuasd3DemtutNajcJRuJwJiR9ExlcipuJlx5itI54RqOanWHePrQQ
E6Nk+mrQaz9fpGflk36j/r6nuXrwKC9ZnQPZTyHM4LigI1qhx0c8YWHsnhClj3w2++4XIkR4PKXF
zpoDxbJpjgs/U/h35jrrpGOJcv2eTzjQoEB81onqmyV/Wwy5W5U5Zw4NVBoG9KNahcTQXvlS/M0I
WN1WE0SEp5bVWdoiqCxiKAA2J0eVfNtwFN3WhqPnT1FyCgFmylS1xoTq6MzLvNXS50nfi5NCLkd/
5f1C9ofhstZKYLWZep73Z8PfLA83SUOTHxmrSsV8bWPHVI4dkb6pjyhEDQpmvw/P+U1bFgyMMkDm
CHyGpfVs+CHbMI+DWHT0FMMnA71N+nSt1ebzCoYZ5Llmfs6gc60a7zj6JtSegH3qUFvNuRIrdpPu
8b+m3xRk1PsCORK88UHx9M52esujr+gVamieSHT3T9/j1gus2L1sIpMgKBjhw9D9J24apk0IwvtT
Gtpmme5cHCLtJhEoA2qtUhAUKibiH47RLC1aKU/FpC7Ls2rOlyqbJyitIoaNHe41a/6SFv9sh75k
hAxqEofIKzcFY0+WiOb2mN9yV1L7j05bZPDIpztKfAZ3OJuquRFBFTsVILqT1pk1KZYGco3cjZkY
GZub2VFEQ7U8F/0XXEV65EpgwLBsWejZBA9457X4cmAjg1TaUR0Rayh3aSyPXNUY9+slaPGoOYSn
V2NEUjYlI8B6efP9WbzfiHsOPsFrL97Dl8bLVWMq3fWjSaaFIffE8qz08KSEi5QQslQPwA9NiIZo
O4o/3eG8jwRNpfXcYs2jyASy9+/VwZtcU4u8ZBwq7tFexvi1I/syGc9QjImtRe1w/vBSF9ikYiSZ
/kv8iAK23ioI1NbliD8gnve1auio1ASEw8s01uDEdBDvB7eCQUd8Wrsb2z4UaOp4YTjPrxJRLfZQ
r9oNiu1srWrhrRkPuL2V484jcbCIa6E8rpNffKky2TxengNY4wTbGAhqaTwNuw+4topLLhdeW61S
MkVQksPqi4WxJxfaIEfH9ezv8s5fKaioFd2+oMbNNfGQy54mjpq+os4RxkARPAiubfFVBJJ1u305
wfCYJuxpB6GcZ8h5NQE6De3S4XcTdcYr9R/JH+SiERaJk2EwQWCze57ZX4Xy0/XWAIhfJYkBWbhr
nUYkAxEB2sCnRN+WC/RxjTZF05D6+zP5wXBNABi5uryGzmsoHLF1DQwk8yDJwlXBZ0rW0hwkuQsH
3cuGwvembK6LtilQPmSpEprQ1hAdoWxnDaAr9l+TQxBEI2fUGvFhyMNCCaiBRKbCIpXfIOYieQ2Q
smx5fhLWp/hdFX23txLQtFJvQJBSG9C6RhZ0fCOsfMLo5dmUQYgpBfxxg94884qbSvrZZCqtFOoo
YPtmVTgeBpMu/KRTCaKx5Xgc5cR+uPohVPyg4FXV+oHpwwoo62Njq4LyLZiLxx8Gs4CVxXPBk/kS
GVo5yyQy4juCOupp6pXcSvjsJ2F7ABsWRvnL+uKmgOsZtHR+2wkXM1hX3ML+YZO+TjKoPpB+6VK9
utQZTvtrVv5FniYqtjee6nI/CYdYDMj4XXgaLcx2DegTIXoi3451HQzQHpS4atGvOhNbRRadn274
TxL4U6MSSDoRLZw32RKjtkb+qkA3zyjYkzNu5WRTLADA9DU8S4oOUHULSFbGywoMx/ACwbLLc4Wc
9qr9P0AEbZdTPtIlDV8CtEWd1Ng+XYPOWSy6ELo41jLzkk7yqIjxTFMoEP75IjfF7qSOwoDAelCX
ywUOBO9+yw16DuPW+/V/VCTgvc35xfP4XHPj3c2v00MR5gIeO7sPmb7LZhtcVGZDGnil24gcBrRc
ktEkCaXmsgygwQdg5N3Zws+kX+JedeIRnCaYI89T3cUsagw8dEI2u1LTJVjVzzgtXW+fejJgleZe
J4fE2lB5jt2fRTczquGvnyVRDo3NmQzlS+jf4gV/lQiFJQ3+kSNfSDvGe82Jad8fCqvNclfyp1X/
zaQr8p0CwePUk/b5+uEswHk3fVGrySBUPdWQFvEtK26NnzziOr87VyZfMZDEIpPfwlwKgq2SdK3/
PT2+U8yW79vRBzbYC91ykP5FMk5LtHYMoL3PPinS8vvwQqTbSA4qj88Imt+jOFniExlWMBgcUEHS
cv92t4Tl2WPsvVS4T8351h46qEvHYaQEcsFhSVQisvQ4+0JMqMce9WAjETeihhNUjKHlZcpB/NwQ
WU/hBbqq4r1Md3Uvp/eB9lY/vI89RN5udyHE28g4hqgJmsrJ3PwKT82IuokVxWN8z3rNo3hlCh0p
cKLLimQjipHhl+5nP07owj0iGbeTGAzXVmn3Mrqj07Src6Q4onu/K4isJL8yNIF5CGKquA5pwsT6
/2lAYBsNk3Ta5rDMoMb+KBDaF8H6NOKpIT3ftzsftyPNNWZMV7rfHZNm50KC4zkDsbOGe+XSPjaX
92oybi1aBcI78YCI97CagjFPwHnXmTuotQe5b9Ih5ev7K9CK/t4TVvjLNe+pGkR3qRML7GkpvPIq
sFw7LaxzRvdAPQbdwWcEY1LP/V9gWkuHuzQQiHkCpYty51iHwJlEmphr5AnTDCOtw95zqKhQauac
vGlWGV+jnWK2/SGryQKVu848HNX09hycrHOkD74dUY7PTwTML/Tvl17O7Mohbq3+Acda9m7AwrAj
ujz1EI6objLx9B/rEDkRpltN6yPpME8aIooGfme1Zxoez46JqejUda7OoX9GbuyPuiw1qxC1Iq9j
K4jILZEsFWmI2Gi7WRgcj0HfvV0Mo5hZkRnRO1jESBaUGLLm00HDdTpgKchdOOuBj+Xst5+nYxeF
IKwAGUqFM+FQPUlGt0dLjITUxILPhDx8iCJtbeQms+zxH2cMe03oz6PbVC2msiBs1Vazz5g3BWRk
dDdW/2kC9t+b+3VqqSn8GZxDa9N7bq0PPKW28SKpZASh9aQnOBSmCQPcSzQkpK2rWsKG5iqD6K92
YN7qU0EsMSJScQCuPHa55vmWMA8VakusJwz9SrHBurk1+oMi6qgobY4WMpw6822rWGP7h2c1zUmJ
J4Imx2VvPqU05fTMgEAsR7DLEScafk6CFy8zdI94D7MqfOumZJq2fTLImCOOyrqy1yv6MU2kIDed
7tNAoUUHKc603SXf8/XoxPvK8a3JZpN87rt+7pMBFMiTMZvFhsiz7y1zjPjelU+WbvJcai5Q8fps
fHAclRLkjzl3CnM+3IqTl9gCNcwG95YPALdL8T6U/3NCMsl15DtJTFbnqZBBlR1Q1BUezbFqnXQf
Lzqov2I/EPbUW8nX0pwkEtBsivOwEIKkxdmRh5SfEC1rYtdurmjJoAmjtbiWgqOt7iINHEULX5iX
x9UMoOYdF+s/ZG4WXBsyxyOrX2FgO7/xTzuO0c/sXcKi/Veq9N5GRy55H/9QrhrzrTiJMTeCPKbf
KUbplSCbU8cPWplettJ5iHKrlqFi7iAaPQDimmNHXT/FlgXe5sm++oYbGeMIF8fb6MuRYEU7BYOg
s/n+Rq7hntcu2gr35mcvd6IJOa6bMkcGF5caRuToqc5f0JKhOUrEaY4tKhCqpzWRVD7CEHu7fXjB
wjkU4RWB/aWAcjMhoe5HEZBOUFuCgLFp6ON1HmDChh25u2a5CSjo4BlW6S/c3Q/IfN4IO0cQFsqP
1A4L8UF/30wKikO6WF47v1tDXnO4fcDXHt3T5NGAoWd2EEHICxCDafQu/cR7XfWHL0edaJXQJMFW
jkgy780swmLdIilSoHf4qx4U/sTdnpnZTWnc8K6xTj0GH5oJVWF3/9luzeT8EvcSMQYvWrTJ0XIj
Q3/TGvIOk6jR2LEjsIl+aC0O9ys6gxfXHfRMn4bmRAdEdPuMvMm5tQ66AnQdPRwwx62upfj9u0qc
LzsAc27NnCCyGwVP19x+98BfTN41TQK54GeOaW/FNFJxl6DdjdAzWTadTmbofWv7GqUT4ewa7/ey
0SuwA9PotToehvSuKzIv5M93wwXh5YgbyCyJOWELDvIiMKpdiYphgrxdyDGHEL2LvHaJ+WPmLEQe
KDdjW3eAezpGWNRMJFWUeJuWzoVWiJ6xrx/+8DAV3sVE0WMjCSv6r1Rt+VY5cgw56b6RUe17LHXv
etTDa5QcJgN/XIWu1+tfxKodA+WsdOu8wB2MdN7fYkFGlIiRyM6e51O2NiY1XxVoAEaTEo0zniO5
B7EDZQNriXr/hAYOjECLByRznj2Wauw9Ouo/M/FNRSauDuUy1J9Sh1I313/hCmypA2FsgZRsahkA
ylimK4enVS+GFfkFcIwMaZkRQwA/PVOsiNaZXk9s9kSLUIsIyyxUJd4jqZebOySOA4wct7J0fSiy
ChUIBZzfjVI3N8ppVkGeWwku9j9ArvFRVKKrVUjHd6ieOHZAAhEdsNrxUwt7X4/QlWMdksfkuBSu
vfhcdWhHk9/VdO83DdhDoBD7YZ7V+JecuPG6oL8pD0noC+gu+aXYSQij1QPxhHYaWbt2ClI+dFQy
BednTiObAC/wHLCEEW2h7Py9o5SDj8u1RYFUzaMuBrzZJIqJi5XtZu5ReCl0jJ69PNNJFro+um5/
5hGWqGYnNu4bX2R9dlKkULDime/FDCJAtuBiEdCUL/WXgNQve+JHGZCs+07kBnV6PA0COC2nwRdc
x0Rh9sRXlE8whR/UJvsiO2gwvEYgT+c4LUmm7XKMRWw9h9eSZUHksiSIVIGjaWejFDBFCrW3daju
YKtYIZhZUMMDZexFpMIFToJipKASOVzFr/LPrjlmLFLTMHLfpSwxvpDzryXOS1OyDKWxXM1MhHuO
dVg3Sk2/Yg8MpusyUiRmgsOSgsSY9NtcnuMKPpmkkr2ddN/E9lj9dvvDYkXCZiqxOht+AUMUEqeK
0w8Fvt6GokCuuxpii8dysSbj7uC66H8bW8M+PtfFGcsG9SZgsBkcTpOamZzX9zJDQ1KpKlHGoo4f
3hRrxdMz3SnjWS0iuUH3airYHSSlOl4cEQ6508VT/96xneGunqz5fzrlxU/X0b7nMQqExrsQkKyJ
YDBSVh/uB/hkxLUGW+ISWTtSTAbFLnAfU+NiAMWuJIZIzemss2/sajrpwaPTe1md/nr1ORvIDFFH
3wOa5a5OP9KC4hD+fi7fx9Cjy3YJj9GV+vDtAOL+cphDJ0H0xAkcNim8oJpKV+F4Xx2J1PLZnZfN
l9sP8HkYFs6RnXVlYF3TnqPAgvot5gG3+qWN2QdMyvsgNRmyPdPcxSjjat+zlyH9WdI/cd3jTmzY
9+s3pFjwnVKvDAlg3JkaXx9cr331E7RtoVVAlrojmKips4mgRFOc6OY0gGoB1yX4l27YtWAVTsLB
pzu+RuPxqDizy9GQsXZnFB+p+x61uBc4Sq8aeWAeqOtFDfZDWfqp9wMOvFE4R76e3v9aXVSciRqN
0xbKrQ2xWp37jlj5WXCagrLKX57f533ibIie4AgGoMvsUJTXJt5U6Id71jF+HyUIctjtfKIkONeG
TrH3kOtLiSjW7TVWLR4tBNsXgGsBvu19esX5O7Y/eZcX8SNfFp+zd4TxyVnQ1vt17StzLvslPXLV
pohmmlhFO/QIT2u7eea5fFzf2Vn0Kyiu/Js1/Q0XIpaYT59h60amyaTelVor0lgQ0z2cNh5NpxAm
NpgZsRXYi8dYXvdTQjnrANHsHvIGVxS3RqSGmzpYSouzZilPT4BotMz9iHcf0GZTUTtVnIqHulBU
IZs+5c9G09CAJ70XSYmYY17UPyUzuFO7DQSe2NKqYixFJSgu+n6VyA337KLlA13ict6svl+lv2Qo
MKAOJ+7080tylSs8efJPrtwIpBpArxjwXvLZXYWFKN+90R0CVP1q5dNSV5lWHefYtpBRWzTDYJu3
ocuki7tN5vyBIeMbT0Nj8hiWdWTylyqlHUVUu+ur2pzolh4lvb5Ay6kWL9UgOlUeuuN5dsqRQv8Q
nYy406sb32oRKHQqstnEYhb4Fg5H76cocdCIgDiUrIBqyU3Um5UaO70SoIRgR8X0VZXAWMWV2qMX
kn9wsVYuNn2HgG1D8ihMcIio/If4xlRCLRGWdPRYVBDaq8EhivyklXYNOP1ukszEkmOmIv/QCXwI
5wkrGdEroK3OuRZV3IoMPSkWSyTPD4mxz1TIcj1p/7scBuvKeBFE0GGjN9a5rzoYk42h2eEmVtfr
TktfJgnKlq5kfA7LcCDXEpOECso3ZOdeuwBOBZ0KGGTS4pb3bKdTrDVwoo49Q54IkuwmQuO5ABmS
x5ycKSXy52ehoEiLLHlfTwCPyy7X1RRvgtZ36ib+bi8kEI8/1Wo1kjRISUq88X7g9lbbPLH8p6aO
Nq0lEbxSdp7v1eUn1WygTU4JeOeltplTOhIV0ryU8VwY2Ne7ufWdHsWcE+QIUapPVd00zWoHKm4f
lOXsIO1ABKM0BvmQHuaokJ/U0ta6r0P5ulwyH734Xn1OArV86Q9jkOryvGry87bCnzDEk/TvQ7Du
xL29MRO5mu4ZzYjDWufhvsAymzhMAmFyOwHMEql/0DnRIrchBIoEh6+awbzGDoFn+b2Hvid8zPBv
qmPYvj74MI9iRwg+rvQt9+n4GjZnDmLjUISMPMyOe+r4vlbeKE2uPd0F84YP7c9xNe75/BuD5CPp
4lcvvUuaz5nGVlHhRPyW0Pzuk53xCDpFg5XOQeifUrotrmhSM71avIMLL6fXZMG6mGXZre5VYqdH
oR4RhHhSUdqUFpZ+B8dJIrDN4fgnnsZOPUSXC9sXMZB75BPiWNCzD+vF6/AncWrOtsmsNdmmh4lA
Li35N87kIa9JaPhZq0w3/0CxhswxUCPzarbZOvptFgK1eLSNY5/dqitHQ1MIyPUYJT7LxEvPPRJp
DfZnAilxdx9gZvL3iADhMno9CHYZOYd19H4dM8/QiHr3WFND4mWY4vSJwtUXe6EB1QLWVaeI4f0I
hO54BSP4CdL4Vx/dSImAPn5X0pTNq1ueBCoOURfxYPj5ILXVGmzFe7PD4ENAfLy8DlUC/amoQr3y
4yHXEPqBAReOXDEeCeVPjYu7iCJ6zCkIv/Sq4XIbBY/pn8QQ03rtbx5NjCimalhlP9LSMrpp/IwF
hqPZJWDoWYAo9nFNjd7V3xywHqzQa0ijLSDyBPLCPxQPj6zUHhMP2AYPL4YUqxBsuHO6D//5ly1B
cAgJOMCxYc9p6X9JnI4qJKt4wpHjvWqVpjJLKFgSYYc3FsfnFwdj0B0sAGCj7rEAdTocPwAYQXSj
mwWtA89RSdU/BS1Ik858dwq1aamY6JvmAonCT9UcIPoWt3ZgvL+9LYgvnPHMVoy0Wq11Kmw3P2e5
Br6LVzFsnqWgOeAALqUeyvDew698gmqDnPqkAjvb1qrLtr0YrbJDmq9l++YaasayZedYK8O2AiQa
rN9cAEmuOBXx/69JrYBbMmQ7BUnWib/7S3rtAt7HhNHdI4PDGNE6GJrtZVJnj8+xXUP+2aHTeJwC
WtQ0DRQQiZfBeU8Va2TbVjtUbjhxjmuNPhP2Z4BYGRBqcxadJIbImPupSoOk3s4SHlQhCJtsjvXS
N1vQwxGRzlZ+QtW8yV8IBX/2YDp6+sJnQ+ewClnO9XKWRYQxGkBv0ajJ3bAys5wcb5W/ocGWbA7u
sOfgTclGZqEjekPV46agbtOybEBf8P8WVfmw6ufSNPIoA/8DnVZHzzt9R+TmBRy1N6GwVQHLD4zm
DhU4LTHG4WAahqBgaNkMW2NFTYkKYqA9HRjJvG3sKeYM/Nkeo/MGUjp7lS/lYpFEIVPhxyiGGDhu
17RwhwJW/Qcn6bO4p8brDwb9fYSX2g9qZbq4M0GA9uYr5N0NBDP3DUMydaJPnDsOIZNYQAtcSHCT
pmxS9uGkKDPCSq/8aax7iA5cHwArlsEpFXUTzThqR+x/tVM7wni743Anuf+W4EF0fIFHGk0sx9OR
k3ZKdoBAczAcuIGx27xdOGaDls/Dpfxks1bLGxPHONCEhDmPafatyMHs68TVnQ4Psu67AqV/Cgq6
tUy9yUaanZlH26Dzt6q01FBJ46wHkvRMcyu5/Cz3XYftcawhtjDDpjsXqcKee3J5ttU2MUPYtrCl
hcp1oEmLAnSLPIwm+9m/ft+WRiUBoAcGFY9w8XLlGPTgS4laTQbz1afzEQ69zBQYxgzO6b26/DRr
WBJyiZ847jqbdUD6MAm53UksTeC4MSsizoplhvp1iJauY9ivYe25FUfTI6IuenSnd+y4kBErzaih
opJGRvkP5LLXNB0x///hTG9mMByVIMHn12ci2UykBHlqL2Fyf6asyC4N6GGHfI3nRGZ/GlaWqSX5
X4RzGr/tZSGkz+zDlqkYZCP/YNSEHbLj3HrYkOOtKr+dnlmtT2eMbmJvAwyIqXNWLE+yNRvbwLzU
d1go9YegWd/ibYzakxYgywxtw19gKrtVZMIRKxWsz8skhSfTOInCDVsLqTGwi6AzTPRbZ6cGgmgV
s7tT8XTsqyHXF7GyZOJDgGBbWSRNPkGefmBH3ihItiGorHDEf1tdpGWlM1KR2O/e4k8f8OuJDYme
RfssbI6JhgWDN/47ShXBBCFzIZRVA1lc47aqkzAsNiXl6u/qIHx3X+5tahXmtrOF8CD5QatyeiP6
qJexA19GyPFbyb3bR+Ried4sLm9CuWIRkfqAPir7ajWaSdf4Yu4TFXjmfmUnaqaWQE986wOq8ac+
h16FoYIKZHNkUAXFgiGXX4v8n6QJ1wxGK/grdR08SubsAL3DxtmdDfvXv+GvzKOcbYsg2tv2NajL
itBe89dIGrYrJUPFrrzDJZ+j7WqnkdMcDEvQAicUX6AO60R5KdCcgkwZSWMKU8R53QHPB6cCYsDl
s1CGnvucNqPjTmnc02cIVLbDAms6qT+V0dTn/EZsVK6ZgSsTAcU6o6YwxUDKSbL08B5i4L5LKsMd
BTeOGVhM808g0sOb/Ipoq7CTN8ZAWeq4OSDlnesYPEJHiRLwMyxMSZxyWCY2ULdFOfuAPl4BSzBQ
qxyjKOOpSDD/6ocPWNHhbFBRpnrvfYTuzAslXaE5PaiGPIgwuwl8hQHotCax+qkADWPZ9+VujMkC
veHqV+1qLNFJyWKzpm4WYjnFBfTIkaaShVl8VIutmdFHNwx2zCtVQR9jshzuBZj6AOfibK7cItBe
8IKZQMDHFWm+9UjULBQCDy3p0ojYz7v8AjFmDCuXd629E2TQES/O2HC1+cTshvl3OS0Xk+Uf086J
yz0wTFh+bCSTw1S+kmEA85WvlFKfPbCy1X9Ft6ylCzX1FE9gO5OoSTHM0jAMpd8WUb7SsTXsaVuH
tmN1x2SRrUpDJ7PJaPKN8L60MjE2Opc/TKMKb2QM4DhcGGLmVC9730zrG+ALFmSooCbGhj/zfRAT
wXdegvwGb4ll2trf3KOdloTWJJGaWZ5rqDIwuepvY7/iIjrEutXI6A6E4K12cTsD69zO7t0F7PKm
NNNGsBqs/6ZzVNgaFCiHBASId1t29aEi/x3SuR85NuhieEHZefe46PCVs1ml2D9cX+S4wPrHvuen
VPpXCyja7RGsry3/zL8bp5ZyGzUUytLcWO7jQtZ2jfKqI7Qm6MCEgPF0uPOjaBiAgo8lsh5Janoa
qRBqBvJ3wfiuB/ydjp9HgRKvxsoFd2apwPTGnAMfzVLNCgwOHew0/NcPHN1XGYfJdaVzSZhWpDKj
3s0Q5e2Y0oj4nKkK1R+Rhb6qYHVKbjvBFAth9Jj7zK2nb6l4KUJcc2gyHP12HbXFrQc40AzaGhwy
MsbhOgpvYpfncAV7jwBFSMUFVgmBCRFfJFREdtP06PYsJP8Neh0BoLuSfGd6EpcwjQVCR8DqdCWl
mZ2BHaZSPdFpptJGWVx2PFJiXRkGDxwxeIhXRRk041wVVYJ4MPNMpJFue6vyUuKb37ISPqBqmHD9
SlFTKhai08CiwAFKsa0DhiKS+w+Cjt9Re2fKAkWvR8oFSTHRHmfWYNI0pAYRpCHJLB7CQouvWHH9
AIVrk/mWSGKlfTMIDdt4g6Tveg+2CvCCgYjTAgQrLm7AbGaBJWOFvgm+z67HoGaiWD01QUuSjDXz
gq5w82GyVdJ3GWc1kAVkIMnyg4xCQ5Ag0u4oXgN6s06MwMw/2KXdRNlaznKfE8zy1SY3a6oQvSal
Bw2sAuXLtutT3A7WdjzoBr2gCJrJTVOh/UAcSzkwSrXJJrNXJcUFdUlPOdaktDqzZYPadgulwusu
6V3MnTzI0QfZ/6H4enrJms8eIjs7dIPF6r0seP7CTOQn4iUi8NbcBcHsm3IK0JCFBnH6lq9YL+bc
H7xfVlh1yRn5ZjnkSAeS6K7tGT8JuLQJc+LkLonzsXrnrAgDPeVYAncSiV2mAs8O9hEVYAGKik2P
cFVR1fEfp7GbAMOHm28/oEI5p9NHDBVv0r17GE7trTSyJTzfJZg3uCRqtzcBHNladngvRA5wQFQv
czctvqnevr47qQPbL8BOkt1+M8SHTrYraULTn1APJpFH03LL64X60feuKuQWzgphS++gsrJynk6G
OxcwSWoM5gg19ikgMIUquyglvZQWNJSua/x/OSe/VWq9wCSOxk3JSypLdMFSN7HeQtHuY7MP9pbR
f+U+9YPn8f113VobVBqTgAbcJfzVmsteH1DmXRZDNH21Tze3km/MI4vcCMN7aonf7UUzXzZbkGUe
Np7JqXUuWI+J279T2z5k35LhwTFC/aBPYpHxuM+HtglQvLTes4s3COASV1EczmfRQDsvvzco6uWE
o1HLQsw3sIK1krBNEOhVVEO2BO7ffU8dc4SXXSxJLgCt6e9gF9/tFe0kzsJbB/wT62zqn1kk0HbJ
KKzQD/mDzcR+8C+EY7dRQlD2JUI6IlfkDq+0pURDoXEOOqzLP0ayyhAF3/XPuA1OtrrX2onJDjaf
D9NDKcUfd4qReORDlO2qbFdlrpORItS0/IGZTtAaSWzDOJdN1/VjqVZsdqhx+4wXth3RHtqyPC9u
hh5RpJ/6qJc/eota2s1rHZYGWpV2UpjHo/xKsTI23TBUzx8sgZGjDUivodZ3b+ORTEnll0Dw6Q3p
xlAqAUg4aTVotUsD4lBH5z505SjgLL8gSznb6xEhcDC+fkPlQB+FKL/EPTysp+g921aH5/y6LkXV
TRG1NfJP2rpL0H0NVu2UH5uh3H05pdxHzhFvtIY/S8BH9df2g9fNYAL+lOPKP+i00ZvkvkO+J7Et
lUtpcssm27+d+qQvZ0GzuTjTJ753A/GptAAvzXS7zbHiRpTMj8sfIWnUdb0AtH95jM1dHjwHnegd
HwhS5EvsB41U28hby+j//ML2GPse6YK6lUDrZHWVZISIjJAlCk/ZPHwqnFnKTsmwDbJUml8dUlfF
gqdP721WZiwGJ9H0Sa3UTYGf9RxeXEKE6zT28kWmiMUvZsI4gugekzxsBKl3tSg2aXV3LR/u93nr
edreUnRQ0GKgn4p+B/Ld4CdC97C+8TVb8aQP7oZ9BXgZuYj7hi1BvwWV2XDnuqCiAWL/OXvNCYoL
k/QoNl4vPYUjSUkU/Rz8JyNiceM/U95EtJ+5SKl6yyESqRyNJs2/hG8g5FX2LAe0ZvB96z+DA/En
SpzeZdEQHw5byXHURUxEvuIs5XNARCo6TKti+FEkW4fGPMEonQAnNajAWrOAjsC6sehqXG/zH2fj
rCmR/oz6KHrsjZyHDwuAUkJ6Kkt8C/hL2ddhbEk+qcbZW/oVWOOk1lbXbUnkn9QS/WnnCocxo5I3
6jYR3MhE5WVkTyUCylBgOH+sOZBSzEI/fz0rGDnxvnSG4P59RTpZyxmPsKBPDuxwVkzYkyRm9JuB
GXF3qPAcCuPhrj76/ZS9gYAOETo4g7bEfJTkzPoa/hc8ytPUfY/6lpcC0HQYjHFwLjYwtZtZCrLP
Dwzw2KKDSLUBwcN6+vf8vhlKzYHkaabrVcg8nmsr2iz3Rr9XXNtUi2z8oKi4I4EcflSE8mESHA5o
BccdGfN/MR47Eh/mCZ/pbCeXXxS3RWfBJmeEWHcI6BZXH5VM1s7hh2e8wfuDh+GI5VH7a+UOtXGz
oK2s5oc4gpvGJd9oOirjh3Q1fYxS6xuabeUbGAGwM8QnM51Ho8RIwIo7bxYoCCdWQXFYVVYAMLdU
2QIblWtefSqv4ywKwSIJfBj6HOX2A5a99CoIRn1CDzNOzEaTNId05YX28Hooln8blmiIQaWMfBkL
zQQaVR3r4oYDOS/2/XbV7oDrvi78WnicpzV7Ow3LemRkUqeCsRhyP0OZp082Y0V01rBdctwUAx81
wBVS5vK2xfHAIFg0n6eRNJxcA5GxNVQJtd86Hbt0cibNYO6t7+PioML+gCKCkY41WR7aEu6AzKSv
nI+xq3gGNSIZ2gPtKWz5sG+Ow13YBq9pqz8KDmQKezOArl8rqxVazMMmzfDCeuLZK7gTQtu6/omI
IUvakvBGtVs7EC/aAMrn6ufejrspZE8SaHIjpSYUWvFVOSWNCXQjpWi8NwH+Bn04AHgBVVMyxJYr
5xzIe1WHduQCTL1HFXQ/5wKcXcNOiwX+Tw/eL01zFS7pOxCDW1pMJtfkj+GbNAQhl0Et9dqnpm4W
Syz16K0mN8AKcyIGIVu6dJngDBjMxYuW7pxEhB/gbetu4WLYNVKAwK4ax2DNS/Vh9E5DTu2VI3z+
PIPGb3GgfizCP0uF1LtJfIQ4ycbHL3XId1xhh4PksB0/WiKre96HPd0Cf1MkiOPWxQjmrCTEUdDL
q5jkc2DBNauxsIW7jptrBGn5/USZhveSn2+aN7lXjwFGMSERPxXyBjZtSmIdS5ayJkJuaxJKHru4
RGVWFoeESf8MSXJUJxwk/MsKrGXBFZn9vdfq72wxuc+Zk9olTYdjk8fx8IzXRIm+q5FvAQAh9t7B
sss4XvUCYXi15YnidFC01A2aeUU3Z1Vn3Zaa+XE3lD+mxTFBeaWsLbJOp8a6OnOF3U/SuiugsTnA
+bUF9UUR45/XhnsHtVG34hLSiHns7EUFaM37ZF3FNgUq1hmwkTfyTsoDXfx/wYkwztfn8v3nrfje
TVi65mmZDVW6TPE2AjgFXZ3LhO6xfysNa3h3ilMDB7hy8F4KbNmOVuJ3VTdL8yLYHKOc8uHZekDW
f0EFve58ZEHvAxO8DiY5jRQB1xduqp7ZGqYjllqA0lafJVlnqbub1KsL8j1Q+AAOlkYKWxtd+MWU
xr58zF0IMY6dUbQC+cpD/mPWvKM2IEiCOgF+QNX7GELNzCtJPCTeTgsvJYsejX2f4dAz70BfjjZB
/e3LJgXdGjh+cHg5SPYmsfj+ykPZPCaVrLvs4WDhkyHhSwcKGswBPkJxHBc6fcPS1a4EIDqVh5IG
LTaJ3kf4M01unEpWGC+FhZKaZMbzZLRlso80HnEqn8Sm0KsuV8bDN0rkpNATwo2RX4f6pk8M+gdZ
qumyunf+HIEf5tqwmfzW3GHhmHly6mzvDvEscp5DZsj7Q8Nz0p/5A60qFSZ69tToORoLuDt0d7S5
IYj572dQBo/91sMujlfwlt+lAvUln5+bbxTTcG+bFcKcpNmAHKvL1y3NBM3sdGewVI3xGbebAn9i
YF1IPFOMeguNNjEJtm7Gr9yp/UHX4o+/i+prLvgOM/P+ehCa4t8e4ItBridU++A/EMs/0MxJ/dDY
EDHwixTf841/rqz7njLzKAWBc2pPZLt+Wjbd7HAquG+hBhpSSJRDZ2txW1BhRUtC1mvo8tK8Ifr7
H9Wd03eFSRteQ62SLmsjfEFjduyoRSCNq742Nx998eeptUUnf4L/uGM4vkyG5e/bMviYl5qIfJQU
XxS0mQrzl93PEtg58taj4cV1QfMTJUy+0cwJ1LFvdhggi6SElqpnWeWEjTBpTKy7BIPpsOmyC+q8
pEyCfVwys4QWHZ49vauhaoVN0RxuTJBTPdIi/BH1hUttVK65SbfoxiX5vblnWPG7wV1zgvomZnev
Gya0XjU7P1oHtg6xUu5KsWCoYtp8NMsgSXs+62LlkZBSvfvo3K9mtZENFGZYk2msgz2Kc7K2tDTw
RuL0z9JHyNm0FSVQ5WYE3HUqcYNC+JJR094Ia8/1yAgCeDpuyB2sKZ+UKc6XB5Yt//O3Ubo7aVY3
xh2Rk7GMpumQORDgjIdlmCGBc1gQhNKng8KE8nOf7rGfoKU7ey4RhmmVY00uzK6uE8ryQNrauDh6
s9iM4g2PIbioKvHj0+z4Hf2ZsCtEkbiLecsjhVfXGo+qm/JOXYJLstpR5/pSE1dN/IVZlyqfna18
JqQJlVMvdSgJ8/JNQkpAd4ndJgnlVYgHCpGV3JKXSAvDrCFxyWFCTyvTZ352imTxqTslFxrI7oOW
3PlCCj5VMrdwAVlZpxnCfK0qCDFEOhVxIaDubLhJbF7NclX0C4Y8qNM/geBatGAZ3kQgRpHorH3j
ydxuJsUbeCPnZCoIV6KetJVrjQynXeF7FlVv0CYqUtnTElQg2ifJn0TIt3WKYXPhRQYpONHslnlH
gVtZO5MkhyjshgqNKcfkn2QokXOWmO5AsKpu7ePf4mU0VABXYq3XciHt8mSHjjKacChtrsT/qJEI
LNQZ5Hnnw4ak1E31GkFp6VEZevKGZzb5Lps8YCXJROZv9bAXuFFEz0mDzqyAse/FcO+JxFoFZMcZ
QH1Vigr/WIqbOxmTVY/m4qc3CgFjvC2g+QKZb6Li6FSSo2d8ztLenqW1aTvbHYMJXQyQpk2KfkdL
Wltb+sBAxtJ7TQKKa+NJ7oESrv1dYLLIX9ETykPe1FaRk5rhMnB2lX0PX0E9q1oXzWPe7Ch5gdXu
7vzOFLao08X7Lt6JJ3lq2fxR/vcCqXGsPqjCrX/zRNLJmOTr23AHD6Pqg0wl6tRh2KTZP++2QxAT
nN9lwznEnb7mwKQ3FC1fknEyRdkhqNMPJq4RUTCVMw+kqYrdoYqEExH8O6OqSBGIw6zjcjyEw9hu
k0wikhdDi6gDwBUjtnH7HyqBgY/NgJFN+czXdYqVXPXNNxjqgMvH8uJgJb3MMdtyhMmvUqMGS6xQ
+8q9H3sp0TWRfD988SkYcEBoXZtQDb3nbegAVkZN82nPTv6EtGceiDS+xk9YizKAaQZKgdzzLxjL
tRgGQaZOgAQMmkIJco/leyrd+6Xg0OGXFkroxkmPNxd5oZTbgSyhzHbJa3dFtZveQRwNs5jE9ZK2
MOGfNFlHV3VC98H35R2aipPPYZLxRA0L2kx0ImhXwYN+PLtCmoEeEQAZzczcdn3mUjq5PvXkcchg
6qfxlMy4pV1rBWk6H5fWQ8ydNVK/kJ/JzVyQM4lXbRdcSKz8YvdT7QrrTdLmmqZCKyGrqTi75/3M
PbHm+OwgIE1R8k7Yifm2MzM1gi+w9y1sZAnRz9rlkrI8QqVHT9kxGfczru2OfZdqCwYYD9ZUuIFh
ybkbtQtywwYT9EP/B96IA1ePD53sFP3en30VrpOwtQeMbuJ748piWSJCPj3+Utd/Le0vs/6wdpCy
Vhrkzkc35HrvNgOerf4Xm8+Lf4/f+9cRK+WW9ec/d45tqQdmwLC+5dm2W+mDSiMNBzpS3oo0g13h
83dP8SFiFNFG9whDTTTIc7qPgHzPhe/sfs4hw+s+JiTlrVvcCQhnak7kbCybTThLFHVbFeqiuIqR
7mEJnbNNts5SpF0XBZZddRLAPCRvA0ityUwgAERLttQdGDdD+lb2nNAOCAGIL3u9QYXFs5nLR193
ueQgCiNBNHLJM0XKq7Jsg5SoXawANvZLV9w8XKMOlluSG96q/ofU88rQyRYsjLHr1hnfz9EcT6pM
KVGTUfutFgLOAN6jltzOCpzi0UZzAP/Zle0DFhoBAMbikB4Z/PPbFdDViKF4txQMlXToWW2fhelh
4GIrhgD20hFs4DWWn7/8cdOzz4mZ8tiOAIF4IdydCiOpb7/I1yIfHmVIUTq2LC4H1FB3C7p3Ay59
qFT/92c9w0lWdWs1TbY99rbtYdlCewVw+NgIOyxhq5SDwBYFzXJQYyXtxPZS3y3b7v4Wt4FYkpK7
TVjeFfbCF9+UUcsAusqxCaGd1xQOkK4HpUcOaNocx2/jPdsorPxzdMWv8dcGMSfLzyiYcJT2cl+I
qJG/LQjwq28nRkIP6haWWgUu6tKTJudC645RDPUyxIk3shEj84JB0503sjG+1wwq1E4leWf5Wtd7
FcDcwXWMwmvoBch1SLdpGVysl2yWhNELW/vN8UQ66eVd5MMFy4Ykoh7AL5TMKkeEeyFXuagQIj4V
/oq19mNtk9/vHvjU3Q1uYG9c937U7TsEkK1MW+/0eK9UG5b7IbdnnjQ/JrsX/WLRIujewDkk1JcT
b98qrVRo4KV/tU5bMJb6oFsjBqnI6XnG3QGaLl6Yy7Db9Aec2QMgQzLCRBynN5aRP5wffTQCcBTZ
LP3i8NqtPZwL9+xOE1iOZbhfwHdnPiedb8IOwrOJTx3JzDw8xtQ2wM/HC12dE2BXqziNcpwoIVHi
cnjp8XE9R1d01FcgulLQMAIUyHpJ/XOUwRzzH5BKF/thRNQLvjSIxduqm+a3Uwye2NyfQs3zS46C
zzH6r2tJDMCgbuE+rsI8v7ksW7SxjNpTf9DNnoeRRL2Njbt6gsLdRy++yOi2Q5tSlZkofamFeyio
XnA9X5TZz6ksStmtNMN8L4g60Bhz3FF9L/xXna1fAuq14elW8vfNGBwbTouP7wLBP+1lFPDuZu3k
FTzTpJR6jE+xudObvGoG/RTLaaQVi6MCeOMg0TwstOenGgH5NdT9n7b/adL890T/rd0s9AufAH+x
uUJ+ecyvSJKGYzUSLPqqTNzQGybzH+FjGNFDzVRQPJogsdONyVn0auXohDOoF//CqejyH/S7lv4D
0K50KBn7g8R+8yG/jAyknMg4Asmmb08JZkZr9W+SZl7CYxqhoTr2mr6hJyCYr/TiTfa3pkg6IPRv
mvk2aTeumAjTV4yqeyQceey55VW4zmq0Ni2keDWvEr+HsFVk9orOY26VjbbLpgrWMDDbXnQ2A37T
g/L/TnYM9NrAd9gcze+jQUfQyUUUjblcL+T90CeidcJWBzid0VqVZRtUjAxJdEhxLc+S+dICyF8G
8rUqqzMVDjyz4OmblBYukVi+pF0xU09/uFv5dL/i7wIM8JQ/OsIWxp1SXbDfEjCSm2DJhzechAVm
qIi198SRipTUguCoXSMYCjM+pfVEArzwTYTcPoXKFqpsPJtuqs8At5NWyONi80GjLl07GTiodkG8
2E2iOlgVclqwoUasVB7WcQ+YaGude/JeygyF/jRvwEyvuuRGG9+5OlUIA9GnKB/AWn+e5ACeoR2i
MGyVyeWbCbE/g8HNI4XuaspniR7IRApids3klod2dy369qcEquWJ1qrWpc+NIv3NG9/OY7bhmSRC
98di/EDXfp5Pm0QvHwlKlrbFpvVYqI14ZCFlGl69iHkYrFkhGFAChZVZofzRwlQVB0C4DbbakeFU
j0w2dhQsou1/SQFK991sWkpwdD/wJyNstK5+uwC7+z6TxDEDeor7OMkTcWWu043SmK6kmqtonkrk
f8r3CmeBWIYS3Ak5YkEZobRdyVI4NV70/LBpSWqxeVL8sDk6//vm+5h5pwdFQ2VazRSKvDP1OlSn
Med+VMmd7NdtNQ9Ku7DZEsPw2zTTjRa5p9heYN2uNw5Whjk/C80fXs+9FSyXg3WHS4RDyqHMYFBe
8dv2lJDzXgMSPeYBHf0dcXgOLvY5tzu7CI4SH1RIlVQfeC6bVq//Y8GQu8kn3g3D9ZvNVa3rSBe4
2ykuUQ/obvtSDTiMqhb29dvfm5Nw67eCyzyXpeNwla9MLinZPFSGWFeExnskxlOgebAcPQ7t7nUI
ZNa8V7iz2BAb5M5CdACV8hdixD+kgdrzTskunDzMf7xrY8fvx6ujUHpGkjrQxnvVswrkPYLbBX6R
w3EQzGLN2Cpm6E4m73f9ibUTgbEICNoU72kJ0t9benYXO8Hpeuq40MLku+9QQDuKvRlR3iRXubZx
QLVYMCmAOzDkS2z5orkbMadQNnotQx7zVzj4LpR55/nGXBF7Y5HpYeV7wOgolqcBzyZgJU7VEl91
+iNdpRyl3InACJRyeMZuDE+R0iFBOfKzI8qHMVJSg45jMPfqhniZVYvxHrGv7nGuHzc7i0IZIrWO
9zbCfjMmc5FNxwhX7MBE6yfJVhNCwdNzORjG/ZqUpUZPtMREpNLRhcwDLhZ7ZQgXK5P5OK+YevD+
nIe66bZu+QzvquP1L0YdgY7PgAqSYJiFbE+eRkxaDo7N2nTbpPb+0SSQFX3Plg1OnAoxp+8noMAV
vmvjjSR85pkvgsFSn0/wdET3FZNmFZHSjhod+Um/DxPZzXexiaYxlrua1wtazmC6pFD1PUp9M0JW
EWI68CbMdiAsGB0lU1NWCb/VsSuV15O7Y5rGBOAeFkOkpX2vn3npd2yWXoH/G2DfEVRcwOoyX//x
I/4ehSpOJWKjl1guDRjMAOi9Itrr/YpYQ9vzbVsgPMcfP3uaDEQQ67Ec8jySeHJL+5r6LuKN/b0Z
CjccpDV03XMT8lm4r42gU29EuI13UXXRML40uPEHNxsDmaq0BWrZpRvkfTh3Ejy0EfjboDeliKas
9ZRkwEcby0pFCAz62Gaobboaz8t87Z6zYIhJaD3/5hYJnxTVQqNovkXfHfU+cZQ/fe2Eit9YJY1r
WiGmgS0bOMajgxhD3uZl5puCoBrA9TqOZMNWwjZgm/g5TGygnQ66HeW8O8ao3AoVejQoTgwIenJD
A9YOLYDuuAnb5iBRpy6YerOyKFcem4dg2Cyo6WQbG2vSS9S7w+9ncXscbeqVLnWiZAsT9XiW2X15
VKh2yOc3zrPqwW6RcJvTZY/dA1RKEIPzsO4rS8gu5NThi9+5uNUMZrBZ2xAGsOw92XYCMpvty0eo
9GJCvaRBUs7wHcOpKsT3n3YbjZWCK3riCImw4UGu3G44XprjXKZzM3vY9kPwOny8C2zFJrXFFx+A
9eTPTGHSiV9hgbfD9n8FOoOp02uYPBEbljRc3HcEhsXMSCutWimrEppMpk80paDyoXmOT2gYWHyQ
MFBoL2Fvtp/H+1B12JZlpyAIuq0LeyDGVcHyT0+EY7dlDnK2snYY6sbg7OPuROZu/R8ATogL6as6
U2SSpv0rk0/WgQDE6zXL8Pm3aS/zMuCP5sIFJx5agng8b9uOCHEQ6rxxoIbfv4xQAofhG2E6A/Ke
u20+1Bz+VJ24k+FUc2wEZwPz57P3LZRG0S/pjp6a/+pEu3zWf1Y6OwU5W8vhCmlcPaHn1iOIBkpa
BhchpugyVomyLbcYHeHYXNuZeO0+MFVOS6qfcrYHHyamUKcUEAIqIe1GBJBiZNw0kn3mu+NU4M9I
uzfTYy+8/yKhq84TmX3qPqW26XRXXYsHDw/p0BLo+IBYCd0fR82RjMOSQc02N8BVIdJIRBQP5jGB
0K+2jpr+4DmQNGd624YI3HboLoGepLTAnHiglnCcySeFuR9MCHo6DYvVyLyBA9umcpCagmqXLBCw
cMuS2v26B6Ogd8pdm6qh672lvgaBcMNV8k4Bj+cxgUUNDW/MsT4QGjpZi9vevujDpU+Fanut53Vz
KGXTWA9p0pxqZysx/qLYU/PT0I6G3o3VkSR0F6rzr69k1G3tPIF4pTTzRBA9ybHSnIjqIMizcgdw
afDdeuDtcxyPY9LTPfb+yOKs2jMdW5FhRGmtnJo+BYEFGLV+D4UPbxCyfbyXqAIKhkqK6+xNvJD1
g0BsBWlhq8zTBCA/dTumMhscnigNw3HO4w4X/eZZsN0hLFDH4y9Y5WKzLZHHxVErCFYbPNZQnyON
Tk7TRwZhKbJjxMPSEWqJ8A7UqWTaH68Nh/gSYY2Fe/3dGeMNBwuOMD2Zr634LWihkA9NtE0N5p5S
0Qln33lsdLwGPZimX3x2ArAigx9gx6e3KXvQ7UlhbqJQz1gG+XpkuLm74MAgveETOnZEL59WXPTB
g19m7ncjFYu3hfolhCclEzvskmGq6qhyRrOdGrkwHtWGH0C6XB6TVXUW6MN9SE5vVgzGJkH1MFHU
bjSLGfaxwBbwWeU3/go6ci1TLo7YtfmQnORM72Ab6vKwdVp8EXTBc21TuhDK+27dbiCdGtIanqKV
tIcSoukdlEB37HsQJ41EplOSuVjQfj9UMjRFGZi9NDSYzpX5if7S4cEkDpcb9F2Ve5FpJGghx8Gp
WZmNsr6fUYRx+OshzyOWIvsy+VLXwCyeeVKfqPYCY60dBXyuD6e/sMjqDPT+0LyHb4Fsnyvb/bLw
HtQUxU5r8MBThsY7kq/012gIoi1h+6gj8sordhBKdpyU4ats7O4lWqS4/SmrjmlkYyBiHHT/dDQq
N/Ah04mdtyx2oa9uA8yrGb7Pg7s0+/D9cUGuA+ds+2uXEhy1uvUdTph4uqlLO17YJYqEf6saw5Rw
2ccAAGyb5juhyV4aY21Bi8hOkTJ+isPEqpzSjMRoo8co6BATKrNOw/d/QTw2XdunCPY18ZBK9TRb
RXmrm8KUznGEAUwhcXZaIlGF9l71FZmpCTAOvdNy3XUTZDf4wzBUZy2Zt/SStpJsJYhRmMVYO6Xz
F7w6rzLLZQ8ZeDaF4t4mq0bD5Y29Wbnm+O4HqaqVlhO9JN0t75Envx85F8sExxPjhVTjb4gXrO8m
077azybBgy21aFTpjIipujz4/nY6FLdVidbjMGYwb9jXZeGC0uozZhd4kjnKj1LLhoHrE/Q6C/Np
2UwbIADQIoyQgTSGbf9RvlJXmImbM7Ra9SW3xVbDxz0J+aKUskLmqVbrCiKldh1YpGRjH8sTMbus
sE7lKTkRFfojmjyrCq1WmjmnPApi+MojGskeq259Cw2RckzVWoJTkjFG0WRjFjau2n14C4RqQXYd
wj744xfZ9Xngutcrq/nn9gfciasCpf8ZD6W5Wi478fJeTO21TgijteSi8x3r9onJK5wIRjIw2vWW
PJ78A0XVNcLOSONpaSg1zCkmkMcAZqqqDw3NB6OlBsVJ0fqVoEfXUG1kMFQ+4jHiDLHoeFHB1qjT
5H0L+TGxsd5rx5ixcDwh96Zxl1RQPzbIBcDgPfL61cxMex3kUnVdlxulp2qP8B84e13+x1j3VNZN
50G3x0GGW/u0C97vrnYZkch4MdPpzNCJGJCZ8dl/43w/GxAo/KdqISRwPbvj6Wcpx7hwnJwVWt7D
PSpg65DLCrBOjguoVRFbPUhk2+Id5l7+dw+aTDP0WMnXjcjOadVOnzUsFLdDs8SwEUyaQK+s8v9v
OeFgA2eqr1A3/u1LU7KEqb78/xhwSoq8YJM3cY0aVKVaxJODDQ/wYRNMTGfeI6aaL6r8fUroUl91
sKkjnns85zVy9gn9542WZ64WaMeopSHrHMrIJfgr6wGzh/Fh3ZeJaKSrh/0qpvmzCTBXNQcW+AjX
HYDcsdQypH45w/U7lEjTrHkkUAbIW5eUkiOJzjcUbZgYBbFxIjdoD/6zKAVqYnNDnGKX/+kkNh90
aRM+yBYoqDY1WcaPRgAjGOHL6PxS9txrV6blF4Z5a5LELLkYzhL85xNjfgKTNacro12HEyohgYm7
vBpZAra0zNNCWbSCkmo8NOwnhqIUdEFh29WWjjlNJzCU4GSZk1PkjxfWHrMu3BQNCzd6rA+gkNhu
YHF4nM3YN91oARddW7pqEVtSyinnznzA5K+1/Ajj/Jdu+1iLIgpCTZ3Yh2jEGP1BrNcog7u4SCz3
vMH30k/lPnhVHQefTdmLUY5XWE3BJiXGwImU0V7Fegcslb3984cm4jgXRaxFm3/XdErJfZ+uHSTg
hyStbbe7cfjLwU0Iz/Bws6ufKPvrv50Lhn5a3WWTMUi0FV7emzAAMBNriqcq8GKimKLLHPvghMDd
xJ1RRSFYP/9JdziJ6/FLkHHCRHDEKSflvFJo3SROwRDUAJwc8EPDgA2K8XJA4UX8jL/wHtydLQBp
iVhVfN1R7Hkwfq6DKi3AwsmpPCKRhv3Mv91f4dYBI+Z+UJWO+arecPd5l1+Om0h04ah2Ra82TXx3
o4+WPUDzvFXOuj4ZJqizQ7oNBAx5GfxIeje4Xe6cODGpPbFIohaigL+X1A6E8v8gnrScvIwXOS2m
uPg6qvhENGaYPyoaT2qAr5n73xl6C6qtaf4+CW/uaZdOPdKk5SPqmsryrmwLA/+X1yEsQKaJHPWY
oYEBbCQeOcHgBzXePdZW561zyNHoeD55Z2ojWWozmcrafxj2OsgxoTSO0Wjhce1miX88v4sM4dnq
1aAfejr3N3RTmCrMWaom5/0yER1OIaPyEgXwlro0Uxr99kra4xGve5VuFHDYMUpf4yAcE30r3dzo
7VaDUfnBJ5X/miCdzpuXsqJ8yR63Y/8tIc/sQ8/L9ncD+iejSltGth8Uyk1ymTXPs3NbP9Cq05uB
cAjF77aOxlU8hUKaWYVwXhKDixT1byM7Q5c6CZ+pdw+DJmVCBBveWQMrQIKKtO3ThuqAy04LF8KM
vUczshCSBV35zJmTDhqRgkoeaARJgG+valyi5dVExo7IiohkG/Cgfjzm75EZIvDPyvMioQ6eeWuK
c/Tib7CxkyBIqH57iCzPACQjVv5CA5agwoLb/njhWNLvBAGLhgu+5/aJMHWi0wQx0RfmVCFsdu+S
EM691eX4wZwF3Lmv4iDaTbpSsde6CTRPc0R6mFkI6gNgMOhjQWP1DH4SKaVlMmDdkhaaBaAuHjzV
dzYGhBpYVqAVTsceW8vJMSGdfSsD7WIv0MpTx5P7zYrdHgCYVmJi+mrova+HYpxgf663K0ya1+8+
XHNTF9r4l+nxsCgmgu0+jgnU96RZi3TJZHscz7Xo4c/XACRle3wW6E2H7TyWFXwPhiyoeD/mtZ18
KVbQed2p5vbMW5FjJFZTHqv7XPIkRJYppA51pBoMqQM3Ed+grR33B2mT+S5CL956SriJ++++5wYC
lkh6oaHRUDM8f1wXfRlsdSI1afUW/Q18mfLfE4ufxSpIMMl4ygihXwydaQGDBZofOsjp0PgIjcV6
kgbTNg7DxVjdXBHMgm8h/32Vc+N4OvmJUgOFTyZS+gNRT9xlaJjA+EfSbgGd1xjjB/pd85uuIS9B
1Bifes9GrM5gdIwW07RKYPCRcfkR/PpKlcOTnjBkiyORhgGletm26+UYKg/HVCSShgA4Ut9pLDNU
xw8o5fgKEJongmWi0jCDTGMyt93ej044TLwpGkiXFxzgQnhlvZ/7rC94dUOuccUi84lgmub+h9vF
OOk/GxgWxkcD+RZJ4EW7eYmqmg+hG7fKdzdZ4hbxqSDjLYJ9crveWq0eKuh+rBkcODOtvFHbudBl
bDYz9xK/XgxwFazsdehP8dxsWFDboOdJRIKHosw9QTEnLlhB//kaiDkskqAo1gxJafEUmLHNKsoc
EqqxbZX+PqGnxYoQ2DSh4OwE2umHz99QmH8t1hmc50QLd+di1X7FGvay7TK9UEl7ia8lUHHdJDHI
tYCRDSSL47CH7ZttqY1juZNFjqB604JWeYHkgL1cP9sD2wjl32DGnIKbxrpppA3Mz6dtKOzj82Rm
PvG2ngoBgGt2aF8C+KOyO1+Qt4UTi8UewonxMTzc6tCpC/VA1KZsz7PUjpNeXOIgTWUsi1JyIld6
0ygFyc3rV0bzl/R/le13UwUY/R0yx2K8aMjN8Fr3kF9u6jC/EYnpkDLDztVSSm4bAqE/oVrNPGLZ
ylQyKUJVLOmiVScNwd2sXrPDTi40DqUKpOibkQWGgYT1v5VP0w8pfDiY80gPow9uYEE6cT1XltBQ
POha/1lySnZszS2JDeU7YHi7kbU7ncHcdwOuY7lck3FNNbFb57ss8rvQT4osAVrbF4Pg9VL38hVQ
dQbi26G7W/qOS9/UPCric85l+b8ZzMnodV5e3Vc2diNIraIsGp6AZltRCKmZhO/ZYfiUUkrbUoDJ
fm6I1zTuBlXgIzrWMrS1jjdoP7xte5/slBYTO2ak2Drp11MtRtjNxVJI08reO17yUsEsuCwl8fN9
nBkv9Vm1M/1SqYLpV/Pmc/o29i6glSZKdxANIa2h3xwUrvhH7x+/n+mr31yjNmbbvME7v9D2C8Pi
sbTW49Ap2NjILk3oCgN4bnDBB5beIb55qEnzh1Be2xr0uLEgZlLJz08yOqzJ+R/J+wPTPvF5JYDh
0aMKlQNoBGTu+hHMSby4limom3YQCVyGH9AOtao6ixaXd0nQb6VZUvqS0Zc7VwiTwvJkwoFaEWaZ
7kd9ASnrbJWT/+frHdu0yb+i3mS1k48R+vMtDee3N3aBd0ITgwRBYe2QxMstWDy6ewlwrSh3XEBK
5gd6dHbkwURbgdPtNvRErDZeKMsQaV37tV1N4qyvVsmnLMzzRcUKOuu8yEMiTTfb5NdThY+41UNO
PGKdxWMf18j5E7BHM3gcYC7BYpYTZoOY5/c5W5ruXJd6xjETEDLhtrCZw4W05illQ9lkA31LFmKX
5vcKC09QW1a/KAdMJwQipa5I5E0KSb8nsG9TV6Fea2DxjPFo81KJ0qame0myb7oHEvj9XxE2E/6I
h9ygofznBQxwzllfJHiKQ3l/qH6pUD8Hm/q9JD5q1LLMLQ09uoGB8vLyb18vwm9F3egQIm297uvv
3U6jySyqXhfW8agoZYlUcMJNh3UBzI57qsU3NaC9NRWTB6izxQYtQmKzfh4LcGj7lrD1g4jL5a3e
54wO5Uk2Lpm8rq3Oh6Q0F4+yE/Qq2HzCliHQ1uoL3FVzGt3EOMdoEXU2UEPoCbLc8yYuCBxXg+em
Dnmgou5TAedsSnupLtqzC0FmiXcu3Iq65GP9SXiOWCDDxv/0CuYZ6b0YnR9AXXOvRBGO2LmBDwMt
H6na+vpk6eoWqjpL79bBh+VoAcwHbP5zSirRWLw8PiA08/3wJf9Ytx6BRn3GpfOZxzP7qBEU4OzF
e1seyRr6Ftr+d1SZkQx9LKweH0zrV0UTMbK0a67c6vNzvFUiCE8j2ZPS4860Ztt0QsMuWcSSazQ3
KcdpEaWYCitNoI55P9l9nAHPklzYVRaql9EtKr7kCJonTLNCXyLfP9S215mewdVu8VUQkr29+NCp
GyC4N0HkzesubYh5kIRd60Dyf3cp7daytzgFpGzG/Xjni1HvmAHQT4Ohj4QnfZ3sh5y/U6sk32Fe
hxig4AYXnumtOJa4oaSnZu6iEekBA8U/SZboehetOhW8hzwMCdB8wiU+k9/t9dk5H57T0q9soRpj
aVPeRNklfoP+Mikq4AxqAcc/1RURqjDw07P7BmWsPY6zpLcIu+mx6/X0es93wPhWBtdvDZcGzh+M
vtbPnfapevSV5cEiMMPVfxSrj8Mee9AbwlnXiaeSzAui3PktN1nmB99SFQ6BFFwc1EuDG/VCQO35
llplyEYyc/KTSY58sxV/MkbZH7IBXCsJEZ90V2O78EbPl7OV+Ij5DQ8bzX0OHztjx9avuEplnO+K
HZrIOmh+7yuOCsr6SAxgz3j26Mbdk5MvbQKZCwiDfEdpzsW08txAJCezbGSEDkLOe2szDxEISuka
2BpVUCcgcNxHKGvMX7RhC8E3vpyVbTcm8VRHzjvOSOa0mG6oA807L6eIHLAeS0E1b6dLOF5L3AFb
TF3TcTjLms9Fnt3uRc77co4fbYoA6OuBe81G94AFD2qnF2oy1OYY828cztXr4+q9SU/XuOuugxdv
KYuR99nVpcxQ7f43qOfoLAzUrrzm0e0rDs7mK9jRRmySYL2eBYwmIOuJ1JpzhWRZb8AyYmt3B+xw
paE0ACGqFTitUaYCumm5c3KcqHtSOoJiC9B2Xkhag7W1XwSX/Q0HaByiZsY+PJYcjFgsLNaHksUh
HuTu93UQLzUWSwlPLYWR/tSgkCMeJppc4Z5kalp0VCB52buiBzEUCCPZ1HqDqH+RMq7WssMBnkmI
fgz7X2Zt/TcPPKisV3dURlPkV0ntPH/lAIhqAyP9vTf3MWD+7NXohOoQxXwUuEupxqbmVWjVZwGk
gOU87V5YMcvN80wfysBT5oEhu7gty7w2mSXSQ1iheFzf17TLjXc54JplJ7hFjn2yV2BgdRK3/wCJ
kEmroY/DkRcUkco+bn0pymRImkw7Szr8j3A8kE/JkWMu72eqJ9AAsVgIte/HI3jkvCCy1XaLse8i
D3RoVzrlwYN81RNpsxrIzcBbbV8dIIZ5QtqW7W0ShELMEBGMDq5eQDjYvWoFgpXo9b+OkSqwVL+W
jHKqFatxK4Eg2PyT/MJLfrcmbVjx9K3iHpLElNVDy70lG/8cx9UMSY2ah27utgV4zTqL0ULAoKfc
LjfOtaILgqHGX4tY8QyDStGZfpOPytojvVQ08ysE/RZ0ol5EZEE54JppZO0Kh/DpK6RMyMb6BDIM
KwL/Z9zNNA4C0CmlEnc5AIiQNsTotsfJOMLMgc51/TRZfcYj+nYtgwyxDBxWScMomFPnsZvd/cUw
FKJL6ED/skVaqk6HWmQVxW4y7etTUw42Xi1DhUvuQLPvFPs1e4h4d0NyUwdIgdeskfhfXpJnvi5y
IZ7Qk9ES0dw1Axv/+F/0KXUg7v8MB4qfM23UzwXf5yxnXEaTafVHdLKDEu8oe4h1bjT2UYkgviCx
lbC8lMdg2d3SaqaC9Twh8JAvQ1DY75YRv/s7WMI3IYeRnzArvg+gt2X4/Qct5MW3tbEyYKMImNLj
v8hUvIFT8zdRIhw1HVqrL+WiQ3CGUCDKhk+ob8CvN6pelzYEWBp6vd/kdP+0eV+tyEE4W97xHTOx
1iwiR4b1lsv9tJ0X64JvrjrdoDGS2nITEDZkbKlULu6DNpjEIn6pWC/8JwmZgoUTNLU5nFoexFRf
3cealm8IH1pEaZgSw5XQSwHsKZvIYl8eol7+qCTf+bjj4L6smgH7synrPHX/tzAOGmyHLJaIoaON
i9UvrSh+3uTl/5wcvyf9Db1N1jVPALp7rpC2Y0eIEek23TiEVxqxH/ZDar7x7NPutj++RnucP0FQ
4axo0EQXqX8mjkwpSEV64mYEUS5vDb5IHMAg+LAh14NTw9DIySK6M+ttilvMDaX20CX8Eg/rCJva
5bqlgvBpi8yw4Gi0NAW4ElV0VLD6+WjrmfNLw2vXpT4S+UAr8RmtyBpqtBT/eTjGlYkbnLBH1x58
YSIoz4hh+RaME3l3fY+hEyj4dJQEg8CFvZw3Ejz5Dwaw3IP1GOokrkPCg5QZ4IKdaEWK8jTh1Mjp
Mqc4QiYwCc0KkIr4ptHf/6xM58Hhs8lNmHrkxk24sSOHGZ1Y+Bb0jyinmKMOl5gyvZGGDuIEUkxh
omRyN00BNealHgV7K8f7InjtEizFoyOA5ygbSX8FHJSnfQtRsLVrMQejcCUp+AdqmFYPQ4hymUiY
hOs654/7ooH3dl+r17Fa/wISZhYOdtPcf9U+dY/ALpZYLYlTZrpPTmRSKAoRNIEgVHHHGOIkyPWt
9GnrSlyc3dZ0I5HSxENAVmEzLmO6bqccvcyWI0XVaiXGade718b/btKeNvHL7z86HZdR7xp6tBhy
zDzHhK1xLRePVv/2102SSNqL8BPxQ1JCNrrjniagPMNgOSwREXkPdb/X/vzglpHQg4RHUeG6fXTy
j++NMrlrRWyFAGC5lm2zFtkB0YvvChBbsRd+vd8w2b/E/PVCgPWpsM/Lp2897m2KsoJEbICeaVOC
D6r5Vm99XYso9SGD2wzrfN37UWmlPUramyLKLg1JQ5HRYLmyk9qNLmMBHScwMz4k3yZNsQcHfVye
88Lqeg6Zl71MFuKY4Ke2P4EloJE9ePsSiI+Gw0pStztmM1aleAB4CON60EBtW1cL9M0zLkhdc29M
WAJHQfMdfuXhnirhYMYDNNaSlloJAn/lgjWvLn9WNn5hcpCpVpm37kBzwF1ABLl6cW/JPoTs2utT
YzQTVyW9J/bMw7N1yMja1VB7jO2QjOLJMt5WGs7GNqFmCf6EPCmBx1esKlaqW3cIqLGHmqiDoLx8
y7liEvOUXxRn/JBoFK8/iSyRCWVBbUXABvITm1Opw9pa4LeocFF0mNbOhsDdZ5On1Gzf6hTAF3Rh
F8VBYjnJwR+2d9Zrf+BJgOEP2oST/ubIilFLGz79U4xLld1IY6ehdkiqd0hSogHHxfk3CQ5+Yonc
vsiMGg7lAZ9g9RU6G3cZEGHmoONsKOdDVFJtHr1voBvMmw3frXBk1HizTjAxqWEnEqh8Nsjj2hvS
urK4Bs66eSv6c0OaPlFiOcxRmjN7sIiJosFgnzP9Yv1BJXAtZYFb22NwUmVk9flhW68GeZG8MlWt
NeFsFIAP7HPyuEaAmnYOPJX3BOimo6hIZ6BXLO6rql8hYyxNctVYFw5rqOZV9R47xV0TuDDy6N1k
OBJo+aRCp+Bfk23ZEfr+5yAohVcFeXYio0kWPWJfqH/ZOoz9Ymd5qPyoLoCLhJUT/HxeRn4rFqYZ
+cI1fGmfbUOvCOfIUYRsblZWwa9WkZ2YQM/brXkgAQliGbHBcX/NYzzVvP/M/Kyzd5WWg+6x8mb+
6B8AnxlzoZFwSfoSLEmDcEO36GRrG5bs/L7bimePdkkFylIuuzt9bgE1wbHIS6qsLzQ5dIN0X09M
88+Ip0RvNQBB2+okqdSV+JJNPy32eYVKO+SirJT0eio31bbA3c0At3CHkyhwVFvnQNohTgly33vO
cD3NBB/3h6gMHJnrFuXqviwsOjwpRilLJ0yRH2A39EUCQMFWk3Qrqm0rnQ0OaZ3D80KhskmwNB40
jIAQsd0FnO+Fe5ceZKYItB9TMi9sY7clj+WmIu0E3h8t4WGRLhmnchqxZguQSAJAczS+ukiLsK3E
Sv2Gncb16v9atTlWcXIPfWVSJplhgZMTWp6tm7lGfmkAtPzq9NrtAUsNwnBNyf/6/52yp3bhqVRX
2tQ+SoVoLcBSyOgRhUv8oVaglMF9bbehwucOtp19gWMDTHiqKw2q2I5YD8THFcMnzJ5eurLdvjZT
BPt9wJMLDBcE4m6B3Qj3Ai8R6zf0A1NxP0jWBNnPtWFPSN6mE/f+oqaar/0rLCbQ6W185zO0CRcg
CbB/fEewAuOQFV7XfknlTIRpc7dyLymMYqqxPxPdjVvNbWWTUDtAnootImmuv/XlS6tq2puH0vGO
LHcSnz6gCBoVMyU6BJ/bUYsqZjmehT85g0dMaH8GZ6YbDiHRntS+pt3P0yW5ZcLO2MO3ezgh+zNS
wHMW9Z5Jbw2O341r+2Qiwvl+weCXlGHLCBBMJ2343dW2eWUXRUKLuTNv64O5oURNCviqv0kHGexm
a1kw2YtplEjEEvvRQVwaflVdJqZQ+tEFS3wNA25ueIpLCzrm8jTQH5dqzg/GQxzvLnm/H2pf2DRS
9t/wymxtg5/AzfMkNJRU19922fs+dCC+21PyFwUFYv+ccLgT3JQXljpe5ExHBVI/bQHXZOb+w8tg
Oxrg7DcVEG3W4mK5Itn/hzbXDtgIlWHXpeK2TxlUxv4uWmdaoJyECQTCoRZhjDiNyUqdvFl7FNk2
68Y2CqGl1KPei9p197hTSi/GiMkS9X69oNzx9URyjuvV7k0kFynomyw80J9ey4LskzvpsyTavIdX
fDQuPssvz0Zc434Usq65VZPAWbN/2cGXnFK47dGYT6AxUndLiHxmJPh9K5/3jaGIVMqAEjuIZoY9
cNQZap9pxtm5ZlxkRINUl1n2hqF3cf9QBVKrHFHTB8tD0mrLqVqhvFQ2TPnfv/BUZU+SkF7OP1I9
W3eH1JJxFHk9u/BuEm/Ko/xmcAHbIDKz4TwOxi/SuSrwALH3xCd+QqvrU8rK2wlfWlSdzwaSCvAY
Ti/Hgbe72nGK/qNRcXrutsI2o9AY/npQg30abttuYNELC3PNYaa1ybke3QBDyvSqrmPbdJ32pZC8
DhzflwBrTN7RxWpjo/XPOX/GBJX21G1YKUWQP1gkWgqqJJYEQu+2P3JRc4Bwi8Ee8faXA/4CNfJ8
WMvwa9oox0wL5QwRT6Dhu8jq9z6lmR5RctARK/ZudGJ3DcEv+cwiaXK1iPEUYCFe7L7RrFbEYmID
Y1AAwwnIqyaf7dv21QKQVU4hTmKbSOzOH+5llQdr2vb0HNhUsxTWWSMiVM13I9ugySuQNoOdTZmK
UfaZxpU8zin5KrOjDBaGUgILFnvih0q31XYXqEcA7cI6tCOabCXx0TfJ7tJxIHdYvfGnNOSd8rAG
27P8+CN8mVcCv1ad0mN8jl5DFx8ZZaredkUeQC6BBKY9BL9W6GbCMt7uewioG8oWJsyWWUPDLRbs
nJKK+Yo5rb0cL75xAtBY/UksMxU5gnN5qiv6jcuzUZlY1y0KROasIJ/Q14nDyGXmg9QnewPSqJRG
+tydIBBmaaloDpdNF7wxZQhkucrBGJfF4mE88j4Ge0XfVmvfnwcxLE+zb4cyT6EajuT0Cis3WqrC
z8WJb1e271x63F6rvWwFLt+s4y7vYWGPwR7HmtPq+3zbOPpsE5ps+14Gr3jtTQSIfUE2W7fdFeyr
gYoVENLU3eOufMI6ZRcSJxLftB4Yl+MKHwvPi+RNto9KJCI79F89d136eBI74woWhrywaXwQIvnC
A26iObYhFiMTkNSyR3F/IVTIquiD6TXtaunDr+r/f5IY30kMUoOaBU8gMzfelb+LkSlay11X+fe5
+aZ4hLRq1RR4aH+4xVdnbkQc1H4agZ2evlZq9Ulwm5gS0OEqvWoz8exI9cxAqPZyvkR1u84L9BCV
wwK1qMesj00CDAdIf6Opbp8iNNqyOhCfT5CcmEuf3clYJa8sumX1awkTHwqKgmcVEkwpjWbhbpcb
fDfvhtO8EbsNrVCKaPU+EzZPO8yq1QwL/LAcyuRipCWrpQblYnYGCrGXP5RiTZYt1OyA/dqFFvJd
48k7P/6/KNYOMn4uiCIZ+J7cOy+BUDjhe0hqu2CQzTb8yUR0UtZ8BRSsXojvCaRBJEFOId1vbbH4
s1Hygw9BPt/7nZQ1NwdjxuNuFhzV/d5ST2iVLwUidLEkiS1FDC/fG0iaPSnrKekRFMp8phS2hD6j
9xPvJmVZ77ZzwF12N4QTOt6RDajhqDj4jVXm5427AkAyskD50Mif1+BvB3jy91tUYZzz1wcadsIb
7ywynVZCpeeK7ErtGpAUs8QshLX2OxPd/IZWrXAKmZVnC+WBz1+jp7mxbLO+9LG19g5P/Rb9HqZf
0TkSglnTCnbKNiqRkgNZrNsPA5gZkPCQqVaWaN9IMAHtMWz6CTIcp53vLp9VRKJ5eJKoZ7wXhB2g
qQY8f5HkadLO+Pe3McEOFjsCpv9fIkdUIhbbeYuEqc7LxoaOFMHlTh2BJ8hVQaDOflRsftpekfTt
aMZOsJMJf5b5cB1d2z8ZfGyQQuwzuX/8GzvBswJ4LjRTBg28ZOYjayy8vKtqOfWaeL7lrroZ72u0
q3lV/5+a/j0FlfCUlBWv+rIX6VRb6BuOZj8Y1NtrPUuoWkcRVFirXOS6ZPF+P6jBquzUPvfwHH+w
8tmWQsQaorO0WE38MW2rQYedJQH9KySpY0PLrdpArZP1LrTwg0yFPhkJj9IJVwBjPDFyq0Vr+5T2
ODH9ESlyTWMP0HQ3JJP6DE+1WZlzx+tnU9FcbSWHRvqTkck0dd8vTHemkHN1mH2so5w9lRzifx3K
HchJrHpekNcB0ftwk/nFaq+21ZLkHR6CG96/o50zBnfy4V2BRBvn76Z4dZUdvuCjUFBvEVyVh3s8
itOjvDfGyIhQX/xcGwP5t1shXKNbz0bGC27tUm5mjHac3E1QiahYekWu6RzO029xjssKFw/98UT4
O204YslisKPbb0qUmjS32ekcBWICleRlNWB4o0O5iSJ6LSpIl6VLSodfNIWQXVomJ4kUuVkIGq/X
KpGEKik/eC5Yvav1cCZ/Qo6mPkZ47TgZ++tbwQgWix3FLPM5UqFRGafUqexRDqjiF93EMiH6VBSN
tt/wvgHGAY+cf2QMo0aQsD84vOTmw4dglwXZ+p5XhMPZevYuUFAjtGNtyzJMIyOFQbSQeR3r8uP8
0oD5yjcBqccd600euVQ/LmktKnd0Xlj4yEbOTV3DJeZMClRP/LFu0MvZi/ikmC9j/BZsxI+CWur7
OWyaCpZTUzpFEevtmhNKEiKWv/pIVg9y9p0hBaGuEFH4PNQRkCve2S9L4wwXqy6lzdEEsG5DEiOf
AQ/b+OZRgFuCOrB+1ctEaBcMLCa977IFtHvuR/uXk6c6yiYmOthw7IeQWpLUL/iT92r4zT51x0HX
c86JOZLbsAO2wculU2tSgk1lMc+HM7b8raMYluPn95TJSfrqNzTnSTaEVnssOnFxcK/fitNL1GDD
o9cP5mdypsWeAhoDD2rUWtZgPjjR3NKCDc/3X7TEBPZgi3ZZfYJZjXW0mOBxNnezN04fQ1w/GzGT
cC3RJ7FnFMk1A3ueZy1xz/r4BW3uyh1TaMSpWfQGaUEU2k0YU/AFp092EiyFhRSI4i6ew8XYL7L3
j2VBvWArboDHBf7XT294qUxw45YVEMaiw+Joh7QV9JZ9tfLoz4wHPOJHyg+hrfA1NPXFbQULNgLD
w5rb0w3tpRfL9LHRC2goNm5vAv01wQSRJYBZtKSDzfPAiSIG7pjO0JYHH1pEi9shPyHOZv3i5Y8J
SbPztysVH1xolh7tNWD7P6Q9Yf8mLsXajr/MBPiwznEKJyau9rMGbjMsRYqEhXiHg8ZgTC9ZLN/V
BOJZTEyrtT+Y6zpB3B5dct5ahGMklz0nti9kqbojTJotFg8D4UOi+4GqKR8jyHk3CeeFKkPc1Low
DoXxktaCHW6VLdLtG64ndediMKyaPiuEgjxTMH0QExGSbcFYE/fJjVkSJjXhK7oR3GcGQI/3HvjC
3ELhkzm4CjnHRJULzgRoq7jw0XLtURLaEb+mssTd7DyIeqc2u4DCST507m1/JAk9XlM2bkB8qLRk
QL25Scj4oGeasHH8GdpTJxV+/LXD/wSUf4mDBc5TxrLBTTmwT1rhXgx/rvT/bpf3A8oFugDgse5w
7tOLq8foANqWS+3lcIAihabYoDGH+hzFtR8PfeN9XCPpazRX3v0EsNwqIpqXs6PhfiJVkSFiS+GX
EvuLX46BvsUw/f3qUCqAuLCPWbgy1iURsFNPvW2Za+2wgeazBmlxvCoiLjWd+dAfpW847YisWgiz
9PIJuJzZSIqGeKcZSN6KAJzKQkrnya+iWAYP7iO7YXpyDzPLj/fEIP2SGgyAZqIFIhZR7IfNfSS7
QkEan0uBxQF7l/SSbiRZOWWTgOWxnw3RUnEeqR51kuI2W0qh1mapjI+diSUNI8xxxzjUvBqTUscx
+LujUomRNNxoOj5h+L7+rytYjmrI35QyQzS6lIXdRm1rgo0Oyjj9uq0byfro9i8MXQ51laoN5YvF
QW9elQudFt9XabZV4MsXUz9T+gnQ4F4r4+j0CiB9Q8y4hRLBJYLFMctvzoidytNaU11B3HPqQRq2
27tAH2mnh3oT/O0ZJ3aXapT32wmFxzh858w2y+qNBvsLy0ljAThdRQELgyJaY389vUMBFAqM+B83
SIeH+qGo2SVUctZgzeNCog0jG3Z6iSV8wbSxCYcRM8lRvKckbsPJPwjUaLfEX1Emiriof/dqL1He
m790c4jjx2z3tT4+gtchSQRzTSC0MWR/D2xqpI5TgD5OBRAodJxZBdjz+SbZ0W9qvwosI3RPecGk
EOQr9GUZg8STryBsiS40bnuC4hw4JIuBxjboB70IBWyIvyjSHnKuPHnkSEYKGbzpqO793eYy7rl/
AeOPUj367ZNnOS9PiQAEgDYE4LXrZTu/ZcVj7lLR/loUElGjiGTCdt4dGu8hdTIhp67TNKH+6GVR
1InUkEEODGckpyXz4rdBMwy8NfRoaSSNmOwqFw3bmtlAAO0A1LU3sXe4bjzqrXHYIBuR2BhiiObk
JY6jfigQSYJ6lBXYuJkXZqFoNdxX7+bbA0NgcElOyPxGpl9KAviK+ITSb89/D4xWn1iZlcs9NFBw
kK2g8l1VaLNzpW9UwVN50mX0ITs+HSi8xvk5ng7FQXr58XOCh+lEdD1YMbO8a6aHYt3p2CXngAQw
WNG3G54R2LEMQX9JMGxyFYuuZFSTydoDKhj5D8VDa+IzUSGV01KzsSGA7yd0bBFWVuotqvzfCCWR
CAYZIH0BTIwwHuZfF3BDMPlNBHpcIpUS7aNjL8bD0uJ8x/NKdKwxoGUIYvfkJPVTdWvjDbssN+9j
uhWk/n1fEmfSHlVRfBXKkW/8E7ImwMF2sQX1u2Bi3evni4+Mawk/p0dmu2PPhJ0/g9sChYaCud9n
rP2sls28A6JEphrKTPmSusqmUCEMPF9EYaJdhysFJ+em6VUAI1fFD9i9YQsKshgthsFxhPFIUkcw
cTC+Zi5k/SNFbYm3/ymkyxghq1+L8J+vCVrMqTz3FxPa8hDVBKL6bDXcJSRh4zdxOiiwdoDEfrLT
vYGf52sOgt9w3ZgA7wTaYD6wXghEC4AiryrBRLNTc/T2+hSUgZtWsbbzmF0INgF5RISUSiFZfzMX
IzCPM3zbletILTO3cnt2OsSmk43YVD/qBIn3834zAbnelAltzYd3bolTaqsn99tTzaSA1PjeTvKw
gzZqookgY2rDhCc81G/0o9Kso7miXN3G3z6ZKw+qcieT1srwtDNx3f7WHC2JdinKHplFWCuPgo2c
xVyKHSFmjwwy7ZF5929s9MLtpgFqSaI/VR3/J/BYahj88CYz8pJCM61eiAwLZgNpiYqxVkR2jeON
jJEwbkhDVc928cyW67t3crnYxdv6E/5RZVL8isemZkagnK2Ngyz0rAxyE8JqNcRw4CCPLmO/6qP8
szKqLtxQYPhPjcYLqehAqjCKMLLLJtnCzLA4Yrr63c7sttYKRyjkH2eEQo9qQGAube5tKLBKN0mM
+ASlPIdrC+4jGXPgs+wLZbQHZQpqbdYWYlRGapXyl7J5JD424Fz71q7Z8MCuZlS/b9s8b7mfXAn4
vCfRf8j/H1Wvju+lUAjXa4a1efNrlci9lBcBW9y/PQ/4uZdh43n1sNhFuCeLZB8FHffrNEgU82w5
tbNBcJJPm6i4xp3/c02inuCaZ+rf2Z8B1RQGb+0NzbY/fNUjXtjsjMIdLc9RSAoT8/IcLIa0kukt
g5O/YPH3YksINu6EvJc0/mBelUsoNEV4SmCdbfbSWZFutVTgpyJIa+z8a/OZBYMwWCRwGLk67X4F
4S4fmmJjf6SThh+vRawyne97N7kmSFmqn/yak6PlCoe1vO5R5UC+2HugL/8m2r7wT6o7QnPfxW86
YLifDONYj3a7MnHlBRdsJkIp2ZcOmXo+EZbKulZ3gOYu/9HySWu+GuZIxsUy46Mj8tHDQhh4x6xW
cXf5YIMOzlQN4k5merlzqOeOOa9NVmxKlA4miVjkbmeDs3rKY46twg+W43eG0raZiX6j2sboTaf9
1JEZ/YZwGD44FQWYD287AYtUufbcMeaDLH2DK/fyANPNN8Lvqarel/G0CsFVPaOhG1SZuh/1f9oZ
66pKpkFEq0RuIl0DArj5vtMXukEUM3SOTyHQyH3KtubS3vtE6aDdSoAedZgrJOmc7ofM9jxOFB+x
wagqGWoJs0vvkTE4W8BmnwvCca+yT8IV1KNcWHTL7m8WtrYLjQCzO6gx/oI6HwmBKTTyNC6knyKb
pS7HmezY4cVV6wbcma+f2mqeShUecazOKZZu746a+MxzGPbWWgaD7beFc+gW5vOz/qKmXISblFai
UhaxasIcc7Go/ZgYnCvcTp5bCnT+wPxj1Rmo5bOpo7BIWG5OhLAZzLq11WlBXiykUL6MxKmKbE3C
JqY+87o8tXqCvlIzaRIuZ9t3mYt+oModUQ3GnT0ymsMrh4YHhW3XahW4NH66TchT7GMLN6xo6iTh
ebWNesZzW6HpNleBPqhLTr9ZpSEsmx4SNt6iq8R6/6b8aTsuPp4+5sGrFHObGqKuErXYMAN9MPor
C5SBLrg5mAXnV63GnfhN6mof24diipStHwKmNk+rHoH88vwvcHWiqtnmENDFu5yHs3mEUQB5e7PV
6foaaCvwWCleeV/ELnyjiaBD1Lq7FI0euXxhOGXR7ylZLnYDMp8fhGMAU7zVQra2F+hvyF6TPO0Z
csjWlGSe+l0EGRZsT2PHp4+m4cFXaMbWfYWzvFJHRpnslE5HippfJ1J1IiHIP7/x7alkjuKNvLuU
1wFPrT4hKkBe/TOloeUuqphydyGglNxqXY0tNw7h/g5k3fGJqxiWxc/jR1SBO+pYfv5YBeOFCwgC
c+sFu7gx/1BE63xknZAtN7+OQbPBHB0NZ5xZmQn/bbLTNBRT27C423evGv9QQKwgzcqPNQ4knAGH
vfcRp1Tb223VWDgz800NLZjcvbPPA8kg1PczP3mVWYpk59g4Np5KzcS4aCYu+tDcBD7wHK9H0ATp
G0wMy1AY4w7OzwA85yhFxnirwnU1R/PcHn4qjsmSG33eZeD/yy6Gm9v7o2dyg78fJ47v8dS0KRG8
yEhOa29Vh9A5FubQ6TcJrpEQ0sE63KrtLBeIxjq2OEtN8b3d/FfZwbTKIMi0ARSxRmEbroFLqeRn
OdP+tcIoeLeNf+a80CZo+MtNorclhVYVhC1kBBRaA4HOYE2eaePkEgkCutHv4TQErO3ssN9uBEqg
biZKeOhW6SRSTuvnhON29nLEAZPzF4uMrV2VVhwRpg7xEr3r89JVH1kJsREP+VfL6bAxpZkCmDJO
IYtT9mcK8gSYngIQ4PIkuckvjz0/XAHoL0rHm6YkRdQh9aRzCFekm+hOKbDmx2Lo/NlzQcbWDNon
k4vNimV6afe88+RLfPyhlhRRNlEgDBCXq69KLHK63FLrkdAPPKVZYHve1GniG5snu6YHvEI0tX9s
8P4JI2KOyPFUMj+8r/F54in6y7iE24zt6MVZpgP176Rf7EmQwssYmAgkyxRrLdjfWpfAjZks+dqT
Ywro+fcxjQm4s7z4SxFMoDKRLE5EzYdhm2zFZAsjQcbl6NjBIqR7PE02OJQtQYdOt5pqrCvr/I1Z
Sg4yJ79Puj3nbz+kqdqfR1SdBdza7eDDkUp59CmISceDcXfde5xmdCaij0+SF+uAfyM7hfwbQ2fY
vSkoXDMpXba0k7h+NXiPkApTJaCWtT/B9zssNy9tB3jQJIm6jERCI53IF1LU/6tKFsjysi720ct4
DD93pLHuf1q/fW/Uc2WYcoyrd6ciJ6ZY7wBG1Jig2Djo9KHi00zChMJm+9NrR/jbrpNjh3m7SozV
u5DKaM6F4vy9dLfUGRoPvv/fiU8BTTcrOhcTrjkDLlunYRUTshl2UPbIKcaSd+YQWAeayNkUX4ZR
6iIVS5sH+szegN+sWT3N3CiI8Rwc/rz0/9e3CD9b9GauOWG0O93g+++BBUvMghl48NWd4Q5cciQo
gpYuB8mmecJfx0Z7lHsNF1cLgVtD5QXc+gumJpvkzWBpLaPJ5ts4JZ66YaTw6NVoLWr/fChdUIWk
mEF4DtLs2fLs41VS9I88P/gQTrzkhO+9Yn5Em/dlc/JGhCR1gbDCHwRsvZwh9CHkof1lGXsBvtFr
6gmhfsb8/hoMWezCcTIXJzkCMf45c6QRYCcWHIFmmT094bS3ZR8BERAinjoX1soJfUU7iZT+4xUC
4uGTHguQo+L6qIq7O18N9ssl/vk2tHgc96fOgpXZ53ngxYaezpvi52WUMb8oHdiJPAKBR3mwpb44
5NVgemc2Nbhwf/UUe4DJE73s8Tv0U9ikp9sbLViUJho8bxN8HH9xRMUGUDm0VCudpJe7GOD268gy
m2hyqiiZcaNr2q6OIlzmqbsQMfFlKJX+eFJtMDwHTSi4728y+X4ZG7BUVdZH8TMKJUXxs2AABiRM
DtKX973O0OFQmPT2rzZhxqphKM+ERbdHLABdszq35CWFO25j8Y2Kvkqp410BiQOHVaTUPmlQNkCc
1xORfL3P6RUGKFDgliVuG1plmneMvSw9xmc3JudWEgxEGRy3DDYT9jnu1gfaJiUfCJ++ycr0Bt8n
B2rBxRmmuqJ9vYhOJgCaDXTKk4M7kkvnZFF2qBOXtox+8SNBhIDB1Or/Y3G5GMkiF6uMkkVzNbVt
9nW2XWThj26UOCotPLpMrQKe0C4B8RhZesIACEtvHu5UNYfCjWuM7tZxhFJeAasZJYoRGnEt672J
xYM5+Ta5J7bDR+AvAurf+yAaZkbTM0pfyuf5YRcIIFvYbBTauaTlMMCMP//n76mtExKgqFHP5rZB
PrkOUqPYSoVGPpA0S5nkqkeled6SgxZbBbWIXf52PhMTD8a74NIMOqCPBgdakqWhqNHY7y5qln3E
oSNzjfQsjTItj1vc3cu8vB2eaLlAx42TgCehRl/l0uEB3bqVfI4i7pefRlPHw+HaNzmRocn8X+Uc
Og2oeMMOTSv6+KbR+NTLJqc1buDa5J4YrtUlO6GejHvtiF6FeaswLGE5W2bTacdswI8b0DQKbgIT
T5HTN3RJIp0uBwCcCa0cFITpamhin6/PcHEWqy0zbXlfiEvbHVpANQQUa85M52RygiiO5Nyf3cGM
jhRHPhreC7hvjATk+ySKZ6msIVm7GqjsnPNaDfcMpTchYedYZMfWYD1BYz0DUpYe6Ow3U+uAAu5C
ogKnD1gwlX1Wkgtjra7r3MNfoVTMX5oEM/gGCaNWNgFVGeNiQ63kf55uMSUXISEvxepVI5UoPGF3
gH6I2nkh8sR4Y+sgV8N/NQOoQrzTpOqzdQDLZpv/kUn+VR+kzg0ze94cTGGxEw88tmZy8C2kUD+b
nrJHqrJAFw6LNPvxOCr2LxCok67eukfgbqehwGRd/FinNK/JD0XF9UEytX7Y0FUu2XglMDyS7iMe
GwYeziO8Q0Ie39fQ2g2k41XLP9DgvgVCEkN6MNP0i3YyNRkMNxv/P9ylgMT8AFVINNigq/ebieY3
MCNm+7NUl3DQTKf/cFvfR5lStCV6McVqAbaMEl59/zgdrRA0KfciPlAxoHxjcHzADj9pt2FksjIc
O8iiJBi35l/x6Bq2IhDcoTs30rxyw16MZX/U98WmdN0UJWKXc3w+jGc3IGUzceEVr72Nv5PJFrY0
nTPf63aZ2kPwLwCbleDu/cB6Wr5XgQxPkTtF/sXAmLBkmJ/usvjjYspfxELSxtWUfQp34Bcu2f2+
74JvIcsRu5U5cm+5+cUEORGfn0eUgjdodeLzre4zwoFqfMmOEIBLg+8+bXG24ZUKGwFuvN0AfB4c
BbkwnmFdm9f/bRFZAhaZv6lRCEK6R0Ins0TuUEFritGBoyn6GCYAvyBlQk/AejIGiCDszP8nrv1R
fsHHCUiLh1TM5r7+5nzBL1arZhT3hqeYP/tj08d5CAaIFFYwhuxf5Ee3WELwbU2iL5eqSNE6X0Rp
KdHybD9oSrVg3eoo7Qap241t1YXTmz8dBruFnMjRss0LOv6gmnL/ajwgYkn1ETeRxMRCNi53ubF8
RwOMl0AgGXdLPYGr5oqXEKtfJ6qzRT2TFRjNqODbrpCusWxDzAewnaRPVmY1w1Mb+1Rxspcn44U/
EgWABIpCZwYSRiJWEdQfsZEGSrFcNY6t1ybtWqShFM+APuHTxT8ZcGM3yFWU3ts/KgHHBHohE/ca
cpLQr8fcQao1fU8k+Pve5OPqVZwfVgMtFfsLolGYzLtOOeLVyhtbUVloRNC1tpe4lKBNGQrBTOy5
TGjVsLlHFYPqRjGyn6z7LCeHZJeoB3cfX/AIGLf8sD618FXPhMeP33FfcRlVU3rlBJSNDbY50506
WQjAyBM2iGVxD9tspsGaKAmKxwZJe62xGvGxR77/2VUelu/CkWQHTLbJodSRbBea7xIPwNDKJkc3
vGZxe2fU91VCPpAZJb5ezzxllrRe2/EDYH/4abHv0QATo4YBIC0yyL8yl9+HNFT5ZkAzkwaRjRLr
nmFh6A764DTCkUmG2lWaEvGuuY8zOCuppadaRnWrpPcInP66h/Zkdw50iLI5HhqEJ9kOJpTLA+zF
5F92L6QVb0qUhBh8yTkFWb83zvtVCIGfli5I/SmAXa+DXnbpJhWptrFCokD+o7TJp8W/KLZOk9Q+
k3aeJ4t0HuH3LhrzRWRkfG0dhi9BouV4tZ8uqYVdEcQmCsX0PdH8ZP+LwjAQAsv/J42n/b6Vw9VP
vg8Q83/MtCUNndiwDToRy4sMJF1iJJDkaTkXv9Oc6WLBIlqOjSaCm9beFHHum0ceoMPzU9MkWBbd
prxkbwx1lx52p1lNXSZpF9NKOfc72tWqoz18rYINUsedf7Vmnl1Tdu/Gk9jH7sIaxR51IUPrdqOR
jO56OwYeKAwq/3rXjuMMiI9FPACDJEShJJfDqOFVnjWUTQwJ5H6EXNG3f96MY9HdWhNeGnXRa3hd
euJVQy2pIL5YzYObjf9oxH2wZFL1TtRZi2VACF/qhqfz777KuOtHLZuXGnciGQqObEPemN0MkA5j
R1wjbJAhRZA3w2is5rLQClM48ynYG9GpHDS9z5PQLS/nroQxCiZyNoXfKRvuQ5Ij3L768bywspft
7MqHvb/3B23SvlZbAHEqme4UQgGsPJwzenDcvpMLzUI6QrUQKlJONQMiN6NTW0xvmLTow5vDxJ0q
9GV/e2bmO1TWo/ApMKGvBPu29uf1YOSgrfswwqT+Y406aCbKi9PaXB6E+m8O/RHdKa3xIsS0BQIM
ny6GQnRLezABCK/2QRbffcnhjVb5iPlRAkds+HqncNqC6FrniSP2fjGtvkZI+LezIY/b6AL0KS4j
Zpghk0ZuSboO44qHljCZWks8jAuCRt0UWkYv4/lwOfllTLGYUeD/XU2XhaxtCGM6zUCiks6fWK32
TjCfLvDTSZOAv+aTgG2X1uA3c6953THc0RgQd3CnnkPwN4mxz02Sq8rkooUiDF2CQpC/0FK6hHBz
pd4YRnivk2k7t/hEK26gNLCOJ97AzceqcdbxCfCK0KD3dNCRB1IqpYCJJPR4czaQCa5ahocvo6NQ
ka3sRjP54lStwP2inHreD/hMSWtorQrE08NSAbFOv65ygUi4g2ezzUWH012EKniD8BTjQGszMb3n
+BjjEkUmoWNVEEQ2ISbCRhc6dUnDyOmyTULicsb2UcAl851nuHDkZn4m9v2ol4AiekWZaNweTb1e
3620CwHGnQvxbMC5JuVlh4ZovUKndMfEfou8z3g2bJJR+3LS7H/CaqK2+QIrogF56QCDLlOa5K4z
JoLyquqdxwnLlWvsTUnNLb/M7fxHRtatKsEsTYAvhZ+8SWb9zD+EWHbtUpv/kFGhXVk5RFnsZZUM
NZyA7GspWCSm1SsKPlP0kX7lHUmz23aN8jJ9+7XVIxTCX9gqU/w2CB7F48r7bjBUnGp1AvXTGAcu
SVXWob/oCXQlEtby66/gnxeNOpG3LMfFeue9JWUjAlNONc4M9eHzV8fiBIo53ZGAr9iILYwSqhSx
DYAAgctZ6rHpul+S+ecPqMOF9JUrDz8UxUaCW2A9/Izt8idT0uimzgg9g17s30mTfp5SQnXsEipq
lEV2gAoR5EtTdYOUQrIf8NDquKobu/mQaXRzL7YW507Yq0PAzm9Xo32CRrGr3u847trykB3qJKFu
4eps/qCOJDIgfFnajHar1azMz6I6SYzv8ypSdmMAIPwjpa+MlnvuTsWM7ka0Dj5Nlo6/oj2O/IWJ
pgRYEv1w3lBqLbDzsxJuVrXvhMTGSvUmEIszwO97Lkcezbg6JW4LTORmjGdEhXgZm31HEXE3tcUP
mu1Wcv83nvd+yrT1SSWSOkqizHyU9hAKsgFlPQV+QD7MvS+sNhcOmMMM+Lhoz1L81ZUbqI+5kWG8
SHIhCzMRnwCMbf9O2q6fA8N8l73OQdlxmSwv7g+ru0yHPF3xPHUssQZgcC7Xi3lA44xCf80Gx+gS
Ibdsq32z1gyQvmsE496jjFJP+pm6phFPo9hGw7g0Kp0FR9Pmkj9DLtkzVEB2ie2BaRZPeVcCg9Sw
4anFgfWXU8yXG7VxEsmP59/Qz6yeHgEbWJwwVbgLuT+1pmmvbbRng4+NGr8Y8usSqVeTZO5J4iKk
sVz7fUDrwq0lZwFWfsp/lyYjopP/hSG+JrqlEj1gmwE4Gsv467fhZJwjvaMQRwzfkDiPrr0IUKP4
sBIEQRlLmS3qEFViPlYDRZfrHE/KaG+w2olBkiWvI9OcqjsB4EZDqXW2tHSB/A6KcW74g+lRuRc8
nBgyJoIAbx+Ca237wTPwR+XHtrQ2iXIqpS1hVHQkqAAajbYlCMQAG9yWZCvoEVYruXRd9o7UM/l/
gfwdIg0DOnExyrQnhBuHE08MNYbAZVtavC6z7hJSjKv6juoZL4kFZlLO7UgHMnk2YITNSy/Jx4Cb
xbdQpINa2PjrY4fTVWXHk/S3E6C8gxwZw38CMSONxLrNPt5dXaIliMxIok3qJqTJJxLLi4ePqGL+
+YjlloBrjQAqi9yoQZ8VtSYri2OeZ/BssGijtD5kcj5lWPqaZulHJf9wXOe7BfBCKGnzHvJrqgEX
C9IWLE+DXiczsJ0WEpxYmMwZRhHX/QE8XqBFy1CqB6zzkcMGvbYj6iao1yQf9PTlvFmTkXhmUSfr
+J6CGr0fJukRA6W4aH2qFImyjeUKGj+ll3ZKVT6mLhFmdyC+vmilAAgH0ZGFANSdkU986JhQ8JXF
sXzPuplMXkA7RzXi0EYH17kJoGye+Rh0ZgVzi1fhyZLwWsUU4nSjAoUPzKEOh1tgRasvMP6lYJOp
UYfbxpL/s7a/+6krIXIxqIKjZUaq1ZeyAekvjNbAMjms2QWWzVzjDZ+ZIpYLgEtJnGKQfGM03zOB
sHvdNAZCNkGCBcLfB6+Jn+Uyri0HlwVyCBL6wmkt99aJIg70j5o0IxfRxvH0c70JI4pQl8eDK1wW
+o5dlt/OhWItfvYV/2BwJ8QKvhMzsGQ2uxRziZd6UzwbYEBj/3g/7Ync4DCQEgKSxJACDH6gxG0M
jKe5I8sHz0SDewcb5gm+NS50P9P1TqJtxDQNpHG8tNhvN11dc59v9d6z+PUxMMzF8K27b7gRgoG0
bEhroAtlcRxzTaiFEEVW2Yai+tAnSLoiorv4/5BhYuISaoqcINbkFwRMsLzBbpDKUDdQlxspfCVS
OpVnAMK4cKcmHzNx/hgXoXEnovpU6fq8sQ1noWq0I6LwTYPjORV3TimHRLczOsclyqT1gJ0gj0kW
HQ8P6bxI4WHOB989Pimb8AITR6rQcv33s6JfUxAdVeAKgtMStVKGyyZ9yvJYmq4GluP51g6joaOJ
8kskyMUSoBQlJV4KnfLri+g6KjoFY88U9iH60Z2hR6s3a99oUT0rM4k+XwLoNSb7fNIl/DBNj1RJ
/yCjowwMSzGXg/WLGhDfJilQnSkbiTeB6lKy1D0pYA5MfXuaTrO2QBd7FMYPkdpXqAItQnEDEBfW
IT4jyLpDUOEqDFFy+TEOoQths8rwNp4/KRthBw700NWKyE2MPvfcFWIXcBvHCUcDH4kWrpb2zuhb
6jgXSF21EnEIe8cOTZdq6DODmXpV/CBAurDgBevMELz1YyvbRMCTIWngl6Ndfg/+sm2TV471QZKk
iWZrChrxjdSuEyb4T5zAzshvX64jQcYxK+fc+lGEeGLi0fPnFQM0UMQel/ozpoRMbYt/vvKAcNhf
UM8xH5iObklSk3uXfTI2B8gnK+aZ8jpGwwdZ1wyB8vRu/cSixkZnKtCL8wscCyCs2ABdJ91rz6Vq
bEjMbERvcEVud2OasU9jJLJ+/V35l87n/ABMvkTdAmaVKZYVgoISD02mqHXHne9oR8VqCsLJvJN/
rWv9AxyKvJTQLLugPAeKNRF8dpTBszgAX/n5d6I2NpEAUkPTsDSJGRT52fNvJvtJMfiUAuY7eKzr
2gdgyTB5StokQ7Sx5znGZFlfcs3EYADS/9cvFgAx0XVgahU8UyO5kq6vLlr9cvkW7tD3zMB7c/51
YTqmz40dZ9YNoUpWIChe5D566u55HjWv1zKidd/UJJOYSmk0kr/Mv6geXcBLy+Tnmz4aQaZbFf1m
D1zZ4dAb3qg+7SYm1RrDmm7E3Dofjtep2UvMILpH5GGtOC2JT/dzjfYMOCKVdXMg5lIkXdAZPMqn
lpsRdY/wNv1SeE51LEefSLa4/cNO+0kP8ylzRb4wzvHZ1j6Vtxq+KGZYk9zt4U3H9t0wsykUyFkG
5CfZA14biRbJPIzI1oo3DEO7ZcuxDbl3rmxbNr9b4PzpD+86T1cMfdYhoRTyTibTiogqGD3/Sa+g
SXFp3n+qey1nRpKkKRG2iQJimFo+xbl7n13i8YMWSCc/aQ/2Ten8Pp7ybOXEKZ2L4UNh2qssFpcf
JQWXLPJ4IrKrDDBkLcKORH1RARVwk1HaowFIt6Nnw1mu8BxVXbftX/IAskxlIC7a2zWteMyowisD
cYB365U9BrAInFmq9ugJlGCJv430gA89IsOCqDkrbrwhl3zEAH1KSaQ4apLSqC6nMQx08MVfpwPe
kfYCo2OuU8VvmuORmX1wfmK7Ijzaf9F4EmhUl/EdAg3jgnV8uFmHOIqmMSyousRSUR9dxN9NqRMg
N3YLHTZq5U3MGpFhoClZuhjc/MGQxyHc8QThc82K7RxToENRxNn95tzj1PeonnEu54Na5vk5zAy1
Pr0ob65OT79o9yrnIWX+gPRRADHRKBYnQ6XlNCAdG8BddXjfpCqK+ij0zwyR2mktERxdFQg/tr+H
ZvKm2cObv6ug4+2bj38nvAXUtGQ+Dm85nz3fdQWB/v2MPGX7l16Py0AxOlyITCmbrSoX6328ks2x
NCc5ikxLokSwcDZILGx8TPyUA16n0rFaYBDcHTrHPYohkgROf5IaKjm/n8AA8bbsewLpISBZj7YX
j5uBew9Ybi7uNkXx+LQ5MfDVQ+XDviYp0ooWvjDW97+KWBiuSwhXVpF/478eawwhDUoSw2TSLJyZ
xn+Y1GS4/hRKtpFv4x3nGflg5D7smA557y9zr+O7v1n/co6zTOxfExKnfy8H26SkD5+myVhbYJw9
Xi/HqxW08ybTEI8XU3S5iaAkut+Kz1QxL5hwYMYN2Ptm/MWhMVSDSxsu4nctyhGQ30j2LxEubnLx
E+kczp9RllkzGznoe2Gd57rmltoDD792E2q4VWRHua7K1j7TJCiKYBK1OOLn3dxRBLaUcXPnoIxV
Wj3hPor3Y/dL/ZZgwOBkgAlYDlOkuCe/f3zimBlPFBEw94Q5g83j6NRoFZfw6piAOxqr9bPdg9h7
fNbG6pyxqgx1mVZMzavHpoT3lPJY+1UmeVUf4OXSGWK+Yt2FN/DTEBN23+ECwfHYB01uMxeAzlge
vfYekOjj23RSkOPIWHcRGRPa8eM6HmTGFATyslEidNYyyUzUIzpPIwQTaiHSp1Ge3hpHPpftqd8Q
Rx/TCOR+i70BkuTTNKO0KP0hSwJTb55haqtnLo+A1FXdouE53e+898t/1fL2KWuRPJsQ3d4Woa2R
6KggPX8UpP3AkEtrmqGTYW1JYdD+TdGQwmDD792MciCyoS8m8r3GLdGiHIB6fAcZ6fzAU1oyGHHT
VHEMH9yeQaqZEPQ3jmPiouzFMzu7++NQ2tioFNfxNS7CFjstslbj67ot2EzhZaQFYhaagdCBZIJR
HTqnaAL7lc4Eoo28UA283HDcH1ZbCwK2qqjnMn8crSnWfXw0BoZTYRo9Woeslbp9BPaM+Xkz65N9
jO/3v+SmIbOd3pjjMSZpVMiSgbezAdjEdaqWQNsVKwosuDc0A+KdWTKo364rZxrwWPnMckooKROe
udia2UoaZerXqbQP4+hdkGvfsUyYyRxUa3GwRKDr2nldxxM/iWY9yWepzp/ukg688dJzAiu5wT+G
DNlwWZF2hJ/YgZsxnKfnvvqkOfsyytZnWq/Wm8RGhVg5T4oFouTDCGyz9JwBAg5t5lQwifPnyMvY
8mJttfaNN/m1/uyEM+sc2MZrwd0K2VO96WwQamHTM/KyFkZNK+HJEkwtb7fF8etzokrK8ycsHOH9
cb/65OBVZkhj/QtbNAM0xMcHkk2TgrMSzlTfGsASSinQgcK/qT5LUdxY1sKKIUBJD46onv348Kgl
36dNjgmV8Kq0w3RzF5FATbp49epBAA9YzoL70HPbD4AhpUzEOUq2F+FlUNSgi2gTkTYrT/bsjTQI
lK+oWeMJzq5Q8Ktr/RYjfTBITHdA7IUrbhnl2YCMj9mCClFJ+37LPDGaC/2jPz3RA/8adkyrWW/d
QLWixVVyMJWqai/ozue3yS57PZzVFu6dOYXChK/kHY3VRJNEz00TzszUyi/8aT8mo0mtvOh1IZpK
+nlFAcbzoZybAtYX55Quqn/BdbhWkr4pDer3Bx7QA8TKF1o/36BNis0H4m95y+Tc+Pc4Re2b5J3c
YtmubQkrh1sEhOjKIQA2yN5ijasia8dUb0oE6Vf0nEBVnBxjLSHKUeY+ZzRsNPTIJATjmvSYDa4C
10jOgvpwq2ZyqswHnfPEhyEMYiV8IxpVFw5D475BanX3OYi2SUkigt4a88ngfhh8sPhuHOsNybyQ
FbEkCR6Q7OGKS/tJTu8kONpDizx9bse3niRbKArhRm420spOKXdAtMN5GRk0VCXzR3bDzAsjnnct
oui6yKfkxHaidIjn064TUTnj6InNvluYV4UCFWDvw1Zfg1YGXXS7xYKV536CYvg1fEHXM2A5jv1h
uNJt/LuCflC5IQD17Kq3lmPnf22syM/32IYafSow8Bb5+Zxt3RNIq0Sofw5m3SL//2AnoLK1TSGZ
VZQXJzRWkSCSjzTsmmD7h3U0WSYvK5LMq3zav2usQdAbFJH8TFz816YJ7n+osdGpXax8tebenscS
DIv0wU1E2e6a+usrH5e9vs5X8YBo63WEps0S3u/0fQMKY4tqAgfwmIvl3BtlWso/UE8StI80xZ0n
F0RgyUoQsknfEsqLuRhbp2MdwCGrHFo4X6e6TVBncAeByH8H+CwUw8oARH4rpM42zbA89PqGFEgz
IxjbU2fi9CfZRBrmfKSc0SF1A4vlV/wpj8T74HxICkcDjH2QrxPix6Kv+FtrEtpMazp1SrWxqLYG
sI++s9fxgfgx0djufhuDPrMiCUHUNTy6TJ45l7YcQBx9Xv3P0yGqbdWpMQqelVdWtpfAjc3y/bq2
lMjIOvyRzB8tqkPH/o/b0tAnVqpocqcfAviVua58C9HCvvnfdlcDZPTxC8jYmkh0vJB2WdaxKEwB
aRk5jEkmeBsvBK/xPYxUPxecxT7tgOjA3gi3W9cMyc/ZC9Dm95W7EcBXrBsB/dGHVpZjJjSw8WCl
yk90jp0qI9JJ7Cb+gDfLyQAsKwaLo9lnEa49HmKRHznQbJDhh0EYX5KVJJbbJE88BBVMOoo22mqb
hvHA0y1leWnkcRBaHDgz/twjBwyfsJOjftG3UzP9h2c9m00448XYhap8qvu9JQu9oqqy7jC74tGQ
pqMHIbG6NWxl8YeezLbk+WJ/RzVEX/jI+ZXl1NwBDcyzOOWakzA/6Z54oX9h0moDFUx92YBmgzDv
JTHTFEOQmlmEZaAvMwFRvkH5eSWNCZ8iObJ97QJ7XiqKu7W+Si31ga9OLjpsxWles8p+jowX6Qkb
daRmJmwsYYv82G442shUhDkRslQAyka/O3Axn5SG56k1cAjo+MV1GbaM0LcDECRHHQXFUM0SH3Wq
zkvBfRnXl296I16zEaFB8dPrGXQzFwy9sAw5aXrxpMb9IkD5KT/ucDwtoTyorDOWABgr5xE3rQ45
XQRxqxnFxRiTzBTsO8V4CsdFca8ZPIUB28MjI0DvxzrUtBj6xLKV2cGpv+FJnr58rTVf8buhY/V4
tdpj1X6wFmJL1i7W9pPAlJz3bliH50IuGrC0rELxqRmvMfETfZyQ2t1efhq/j1Go8KOLkyvhqT9s
GxNPZBQjrBNS/DXcusy5D6TOzHcVybAJiSjGV0AzpGE7oGiZSkZyuEAG94j3y3GIijJnlvLpXp+p
BneBTDv2p6cPBpcW6BpJILi9d+JRebNPXrojNCMdc2poTlYgHH/kXqmf+iDUlKmRECYjRt83+8SX
lqWqPRlKy93u9Mza5i/pfRp1DCDAOlTYsu4fi498qB3lcLsYyg6KfsMJ57k0U/NIgc3+Zzbop2k1
ozkDuAzR1jrMuUhp8IPLdRB4FxFoYYuSAxo9qFhpyE9SQfG0AbF4LN8j84tvh+ez6IrUfQqvLxKG
Jkk2hWMlyNxqM8NibqVMJH7AoA42CcIuFkJ/vwNC6mvTtPU/kNRIzLjgpS6lJvoNHUR00aSmlSDo
SA/Jz2xLfWn+9AQAgnSpJxW7rjrfezUEx4dQIEgxYLniQD4yrPbNEbBBSlqg0v9O2EoAJM1WvkrM
M/ivc8wRtQjHLX1aRuoQ8zDwvmD4JylkTG6Qhe4Pqr/QvNmu9My8zJ3QlGDPQhBaNCjX5npHi+l4
0qSx7uiXe8xE6f1lfXI146dc7poqDRg3AwYrXNVmZSZel8MT63zofz/7jj/1CgQufwJw0t6lWFDz
2k03/EBuvwqVueRwA28TfAa3Ul95GLXWKuqxKkNYxevYS7q79nDXi3cHm6qJQ81UPjoWgeQx6VN4
VPtCKBi1/mj57GXFypXUJpdcINR+Z5LE/CDNJTd4MUAwiLGYssHJkw0MrGue1pHw+TNOJ2h5Vcyb
0SyomwVjc/qZ1RxNXLYNndOyHYsVX143+Yhxj2Mk/o4Klu2sl+7kfrOADf/ei7zlMRh56tHQuhSI
LZzwv2RkvWp2lNsdHIm3hq2mk0oAlYSFutf5d/T7AvSgox5dYQ+66DgpC1GuZn5zZbM2/cmVDvsB
PzlBwQ5j139hvKCd9diXNV1mF8c5nSP1gJD3oyigJ371vEE4GBU3JqYb7gKSlKs3jEMWxgGUNsRr
ZeOZHZWPIOMSII/2eYINX6m6z7gAIoON4/14IlBt1Z6GdfnBRWne4Vvdyn42Zy7Z4rrJw6w/Q2UO
YonrXmqt50+elSopnvXIxsHZh59UOqkjlxiX9QVej+xOHGAVqmsxfnKwr8S8TCbPRq77AIjgQdBn
N8Cmok7RC7I4ISpJhS5+f28N9RZlxxMg21hZLvdOB3BoqZrK5wTDPw/qEMgbI1ZgWJsMe++ES0NV
mVMcjWCKKFTARFK9hsHLwQK0y6ndTLFrwmAKLNROAnRx+QKu7b5F48uSX+luh/IqJ7cpxHGmEAiG
eQ8wyoJNN8YX3CPSfnczIq9lnKeY2ZkPTNJTAsDirL50nBA5XHVDZT0gvVoetXqCTX6wwNqWM95N
H2b2yKkQ/9D2WeDTu/HgSpvlavgOW+K0f3slnCZEzwMYXiAEAng+2fDTuyoybuDL0OHUG4X7Nvkf
/wbql9ZTYCl/aZek0qrOmmHdrwDZglHszpgD5H/WGoBEW6xkBIBR9cyYi0Llh80FwErVxum34YgS
/uEIvUzuAWSZiS8JRB60XdYnhVcd1dZ/+NQiatSy3M905Z3aXA115iFYFUvlUwJt989R5QPKK5Aa
5U/6ipfATBQVTXXbuAvZMyThWtgSYDG85Vtz/66leM9AyTEBrRWWxZj3uqVhdDGJ96nfWtpXdT02
vHD7aWFpOTOXOWnVDZLwNVYFLRQq963eRnZbMUyvLkpLIwpGhgh23M8itoLmo/7vwzHrWYOTMYkx
/nI+wpw5ai29wV4asc+IggP3QD/kjtWjtiDr+jGiLKC1f30EIeegJp8mYuB9VglVzhu18dF2QmGY
0MJS5HluPNvaMpyIVTSa5wuU8HgiNmlKrvnKhD/I1AzPRjXLVHmngQeAcAfgc18GcLopDLPOecps
qCs/V17hsLgW+B5SDtyecjEzu292dNbG19sbnDCWCFlFcsIFEHaIVNbciSVn1cBWacN7+k0+85dI
z7hPzxD+Iu2b/ftdGNvcjrn0PwnOfX7QCLKLz0zBIXPctVecbTZ+6sJTp1lQF1mNlaDwQFYob7iB
fJB26A8kQdhblhiWbtC3kXwWXnKGus99D6XbNJWQlHcSwCLdMBt0UZzTC/lonaADXridDhOx8YEq
cWkvfGY6L3QsUu1X8r5UfVm5Iw8JETG0qxs37YNATMZ2a0ZAATH+H3PnUZ5E/MQih/jNKpqo0q6Z
ujuydS4MZSSEBDljUdwhqxuXHsLJ/ZSarLCkeN4RUZsskWjENzAuAw0NMK4odznrDrc0qnjVXLAg
TLLLIEa/EH3dFRSn3rnVpVxz/k/WzaVflsSqyFo7qSfldTmf/xU3yfNxL/ylXwDOowiiXxN2LkT3
MsLkgix0gCV8mpAzBx4RT+IY+BZZEWd3SOh/VnF4NJ9jbW/Gdw8Odw5oPRrqwZPeWP4xb/AmLXdP
fVFdjQYrwaSrOoewuayWA7ZRlVyrCBNHcw5831HfzzPzD81HTpDt5DIZ5bsjVjmf4Zs7AuJl+qq6
ZPf8fPkQxtWvpwbYmH3JPIeJcHbyvNSu9uSPAwDdjqLg+EeinB9oy36v3HQxayutPxWMoSIj20MC
RmMRPB5iR4OX13g9SvIv7+1w17g7/KQHcsF5DosA5dBYdbZjLhQeVlD6gCDFkjSl5baHkV+///4G
zjcr4OYcrIO6EX1x3MmCVRRUrJssQyIVpDnS9DJ7xDUf7/5BrowDhKxMJfpJZzNKAyVFYHSPaOOt
offZmCi02cIaY+V437stGCqQBeozS8wEdcGJ5cTbbVqnYNG/PYN82j8l8wSSIlTGtbjd5+XOOiYN
ZaIafwGvc1pXrFcVNO7hpr8GIawFZ6vwo33ONBFEHtfZhX/r4cOjjOw85SsbIUVf9NlTiM2YrEZA
7sed3hu6RFxB52JnkQEN0LMR3mKykkqk7bK9fhzHpFGQoKMKclSkEgQoF7hPD9QfAubwDgLM89gv
H2pbpy3HUHH7nlI4xVFl/KyFbHs4nJCLK4gBodHR6DM1Kg9xMEb/ZVbw8ER6rrv2bB1Nw9E5IORb
akYKntX22BaCpFJ5nAQuR73QHvheMCQuokUSIX//VMFWa3MzILCFIuWHfmVO5KiZaFvySVCGqahP
5PPAphYbvx1COddOWlap9AAZ4YVN7F/Ne3vN6YFqA/9ikPPiQ1obk77plQUi4Uy0vZ9BE9tE33qb
Zu1dCnaXWAqXKmGZhMeu4VW7ykU80oG9x/iLTb9JFBAwF14SScJj4iq/bWGUs5ukoLvt8/Ep/l8R
kM9Jeh0gs27SuPmGj1rxUjFNFnQizmeOWLv60NowwLC/RnDxq2ClTMb0CZgoqwam0oyywkwThfiT
+XmuWBPNMMnwpBV/xV93LoSw5ZdU4oSbu8b2aktWkn+FEfNDYO6pJk71eucfb51a7PBetK6+sLU1
FV44Ufx7I0jkGDtM+rrohHn+Y1M1wmidMLIP/qnyJeunXtNhNSlCa0z94yiKd52evKW5x86N+luu
ghel3+lZjtUIaMPMU/Pnn/iwNt+TGDD66YDlsYf+Xnk+jiERbQmQncJj1v173jjZxL5E4fDheipj
l7/9sWvuPW3oXxXlEqUWODTjsI7BStfhGXZAeTjoM1N6DQ9hQ/mC75lahjpy2xkrrG2xmS5iuFtm
mqzzC8MvsjS3hvtRUEeVJ/m7HfqVq69Z+Z9afckbGv8j7+4PsuGzN7Izv8A8jSFqydNPOA5g3Pgy
33XT8m81U/11eEF4ozs9uWkrVJkGUIjcB6+qdMKXuSVkT0kANBWFGDHBE5EpZ58Ll43qyLM6f/7I
oqN8PECZ8cg/3iGMZ32XTs0UgWsUU1gZmsfRSfim9nUCPzxO7pslgYrdRfF12ZL5wbNlYZQXOad4
ynq+bYCPAVRY6VhaK0f/3A9jVQTGng16BoNMatR0ux/vPnvj56Ndo+o9r5wLaP9wEHbADjBNWhPJ
Uf7ctg4yPwdwUCJXKL8HAo+NwbTmiZdX4Xx+2fo2osHhXVHT/YeQ+WGQ9qJ1LZAde7+eepCCM5Hf
yvqYqNPWhLFoaIVcTRH7cdMpX8Sq3i5LJogsKJ1tEjSL0DgYQNUBdReQHzN04VTVvD4baTkLMn2P
G4p13tpbaNxTS8+qSHZ8WjDlI/QR4fHXZ9S0Q8wLnXAkMEvfkdd2BV347CoWTHg8HTD2UmsAWLi4
Uwu4OPWaKK106wX1icEF3NxlX/8Zsl21H7jDJFteUSaJnze4881lLJ1rlfQXsGDWC8UFNqiWwZ0v
UKNd2LphrWDHycYIeffqob2bnZT7y9Zw4nhI2lwRyZpa4Xi8GSfv4T/d5q+xZINTBOlMIuv2/UhU
ZQKfkOLq25fY/vJyoS3ZiiGItZ0Coa030nhRvT5GQdB/pUVZBcsW4IOtB1Zwi1DHsVBa6xcsT/T+
1eG2DWvF37E5rklJuY54Y8I5CbN6p+7siJuI8K3+eHXejgyC8eAYv3NCTGdZUyM5JWiMeQqA8P0L
+NQQciSVpTOGjEvdfl0FiGI3vHhKE76+x7KFx+e0UGU6PRhVdQQ6n3aSBLhVNG44X46zwOnVcjGA
MnyoNxnBsDD8knoJBGbPfQEpLvfeNMqOEfGQ+ix7QL4I7OpubvrhYko6zllHgqtkZ7K/MB3/MDyl
sWmJ7rwuLyPdnTNUufOxfkcy8AswQV2TnLrecOTRc1cFNchl40g+6ku8CwQoDBaCza4uAtAQv0Ii
7/9PyF8RJUkQdQHpdcJ9I8HpByVbLOHhWQ0Ct1Pi7+XvYRXp0gki1Z1eJYvMOa0q8Jvy+fp1t1/D
GN42fFePS7rYvB1fxUtlXfh+OHWhXTUAI1qJs2xZoVqfOeM9hKWYMcFepspOJPBFicasqucn9m2a
YcBNq0Hjg8rYME+rFxTdcX2YqUumWTCg/9s+DQLMYU7LmfnBezCt6lUc0/16V3rZMgiaaMYoJu+0
W8MIngPQEtZ9sNMzxN1NH3aTUEcsgab7TSS3gfSJaY6vHq6ZSiYYHh/vY91cTeqm1Ul2mQDFRuIu
UWZJDCkBaa4XrtYxuXQtiExO+8lyAs/Yn46Sjlv4h+O5Y6R47hUCHez3H0Fp6SG5RPGtS4RnENMH
8q6rDQ6aFJb7pQEGG4XRDepSBHVlvUyLSsRX1LVMiFnLCAeA9fLy4+BToJusTisbhP1j0mj5oVbw
P3minCm2M3DgcAgyLIevfFdOS8vgRe0qjXGpDsk1gcUAVouzvwU4yUz1GJQlMWyyMqIUANDvWPzA
NpVoQltk41ICg4HIqEpQDJeeSON0xTcMwYqCabfYITawXsuvYPiE1vLglN/VeKWo9Dz1N2TsDVQ8
BdP3In+TwbC1HMibAa/pORjXoOf2U2QNwrLXVyopx5aRrB/KvIVYIlCDP8xygI6IwYCxgvzqzyTa
8I7iB1B7EzZrZwjddtoxfkdTbHeTn3FTdDWM8K00jAkX3f5MhbaF/5ZenkRBaYLxpueD6FaqXGQV
qyzthpUh3hGmUmBHOI8moELVxifRU51p7RUB1OyVzXXKYn1Q26JQ18lt7tjJ5zsyqEyE9dJ3VgZN
fHFqg0EsxGiaQ6KcW6TXRT5KUpBwarFEth5H6QZiM75QqLBHg4S2SjpgrKf76WMfxU7cDjF2MzmT
oOMW5QkqGVEbIFbRMbo6huPRFL5mwIiKj0J06Jxkrm3xYFHS1dqYCJEIgVt80FTGVgSaxp9H/W6o
uhAiSpDbcvw7HFWn1a4Q4E6rIg4obUIk1aNvI3azmnL4AJ0JdvUTL4k+Y5AkqC7X6oLo3GrQ5bYF
01ICwIaXpgm81Su6ekhU9o+1gnjc9CNJXy911pw050zrRNQ9CtTb5KHHM0SRiuB7MLAhuGTlxqr5
93f/OfZmyEnfI3JCS/Vq/xwopFKQHdpiLKVOfvzPM6LZ/vkvHlzEdwHNXgbC0HqDddUJ/KYLZP6u
z7LjSTN7nB5EeR6rAZ+/y6PPRZu9Xsa/liESKWI5il9TBUbUVQQO1solSt0qHrLOD025qzP2oPIo
+nDJDoZseLCjxDuXtWnzTyPHDCI6i/RWQbaJOfvTczIWwhgMAZQrgPUU7DzOnvKtUig2B6bGKKy5
k94qrU1mLgN7Bq77eVocbt/NdbmPnIDoFzNNF1Q0PkOKQnR8LkrqZxfRzvOyMVmBTV8bXYBQKsoL
f1vIClzWrpkjs0BqvFA2OnbB/DTI1XnDLYuMSTsAWxrSCxuF8xTVIAefAqLKHRSDLEuoriMrHqWd
IsRY5p05L1j9OdllBRYuolHZZO3bGNyoO/FAuUQ+dQQTFNkZ1gCcarv15m81UJBbod93NOdW69rF
1PfE9DoTOn23eqEtNlwvTFHpB/G8wrYDGhzgi0LHacoaC31rsem4JU1h/NExRAE6TGGdfPEIdbkk
bwlHySPUG1jLvk4oEAwUIFM+IvF/YqYAKJBv6izvYKISlK7jvzartQ/4aSQhjc4nftoL7gvtjbHW
qA9ESzSvq9DuTzWFx/a+hiytnDuuTrJkavXJIp4RZNW3oEEiDtPZfN07q2DxyhLPypAhYXcRNoMC
cgjCw8zfRiW6a4ahWTQHqVEfpIDdV5T90vJYoOLUCR2A6UFBEw6XJwrdK7vvJp4GCHpZceZnJKKS
5WYnamMzEpSxUMyCvkeSRgXG1LrAakD1RFUPkoF2aryBQ57n78y4gbr2Zt9fnyaYAfLeRR/ZbXd+
g2B1xWxDowiEvqxJ1XQBzkypRaRqTq1x8uSVvHWF/q1wipqRQMZuB8qgH1sDMVSNIVdTA1YY+2Pn
VRc7yG1eVkTaqWmQ3DVtmv/r6XhU1WLhDSMKAUbuWtKtQnPWOFXwt56Lc7enekgbpQlWGhgKJafK
QTx6M/EFtN0Y3UGD1uGZWIaJsSuhKJyEtooHPnnkcXfFD8YH26Ax7EaJDjMKMNBpBO0r71w7iBcW
uQV/94qO5dMpDliud237yHAF4LPFm4HV/X0TTjv1R4an0xqC7lBveTiWmeGFHJzcnWaa2N2tji/L
NRmPDSl5LEGV5vDWTpmKE4wz9ny/4OWmYb2l93rPv1kCgCzSFWMEYcZohq2sX4dPDZcGjYwW9Cuq
PRxsdswEFgpJRY31MXT8c825R+N2fxVdruDA2lMNC+p6w+4WQm9VILR4KafMoh9Iwv3lBtqKyAkZ
17Y4gAjFVRER6GC1runB08Ho369f/3PtiBMIO4JWAEkVCLNKs3wJ3L5E8cgGkp9OHWF/Sliohr2i
wRw1QQZgyN0KfOg66OyB5HchdAV3Afu113sBXQCvS4z8Qo4y1QfvwndpTWV6OK73NK6GI4hBQGEq
c9cvu9X/0yas7O1Ox3JWhtGJvsNwNjGzICFJYpxew1fky3/hiwHI9wlmiGinMdRO3/tr7c2X3IqF
8fVdJj6qAun8qhSG2X5yZMz5xBeOtMYiiifaUeIWNSPnXgtNAC4awDZjI2ZLUxmaz3z1f9e+HV2K
KP9r9xC5fIKiMC8Xq9iS42gP4FyyB6nEHr6k7QPfJaPXydtXOhntiJxtB4yuT18RI2GNLbaDEwH7
koACuHZH0ct1Jzee1CT9hBdu8kWRCUWNDAdGAmUYgSG2fR9HScumk59yTiITDHyNrPyBgXVpjsY/
5FGb7CpuzQPY02YG7R3f2ZJX6Sud9QDDy9OWcCeQIB0js7JVfTAYUGGRKrMKL7teQ1+898GHNU1H
yUhST5LhR4nNC8nF5o30wWqLSPpa4P3R2wRMmXS6ifEhXcUHnH/9hzCM1IM4n6YioJFJ52eM6Ne9
D7CsZ2U2oxZv+hn1mSE2/JeISeNiyKtLCnD3MLkmWlmZPNqVI+J0aA24Y8oHXdMDGbaFSVpTHDm9
ZEw/E3zfTUrUTulmuR6B0alsRuhtgQJmo6hnZ91kMQwiFzhNuLlzvJPcDdKozuIgRwwXBw8AFJIj
+icp/AFVlxDT/lmR0a6KbXA343ybqN/ajT9QEaXcVWnZUC6CFMA4zV7zHQusmfAFhAz7w6A//i4R
IBcuN4+q2ozq5bcEBD0nHmiWO5BO+DFQ3BMfgu/HkcBIb9PekFwpi18yoVU9+Zjz7xYVlDPYSRJU
XqvU3b/tt1zn5+NDIlPRJSOoAznJhLbnKaK73vNGN5LB7YktTiAW0dFU45IpByKWOencN4AtCPUk
rbpFfd2Mc63grL+m1FuIGCIN8ZLbiiP5FM7rKhm6aNZLW/THonvTayB2atd44gSZ/GRk9YgCbOsI
u4npg7ZhiQu13T3QLq6ThIc4pf8NQZ9EYtbBCIwE7qNc4th/HJaMQyg9fI5aIgn3NjR2jjxfYVTP
HyjCzRHIGJs7m/YSdBY/G7qV32y0skOai6L4BG0T/l1wVPoKYg9g0hKvCPnyB7YiqEW35cRz5l9F
BCrXFT0AeE3yBjTZKoyq8V6huxI2MufpgmMDQwpfzXNiHopdUt7zrsa/fZe/bNeAKY38yWw37EPU
JVUC/GmsW3og/kHvhYpxI69eJ8IefKOma5CeihHHHWfKUU9LRu/zGP/dLRYU1JXeIUNkEqnqpkxS
nndI0DhGjX/iaWvaS4M4JUpDmPMMmeLq3qsBx2YYJRhvHQh0NF3F4jTH/J24sDgkwxuhM6KFkAF4
lYe8ZfZuXX8jlIjvwPDZ0v6CJmL42VU9eFeGqX5eGuI7DE7IKWvtQoOBUHOXrffDuw/9ceepwF9h
0RNYVVLqz8GHI76ZVrAg/KlEXv/7ukPlnN/543xF3McsYAWjIRlnGpmcxtTkLHGpLrhy4b58yvfC
v8y/Ah9qQbiBTpoVhX39vpBBqY9XrWX1EC3wS0nAtP07zxyK9tNqBPmAlfhLTCuPFp+xW9G2l83T
cavTnIY99kywEvVV2h/3CzVb9KxH8gz0Az81l+1FBp9Zq+E2VjZDYG+gaR192vnceveLxdo97xCh
plegvfnE/Jib4oy0ITfVEIGhWCmge/OG5qN5Jj7BJKGF62f4++Cl8b1/Fu5zGMX4XhHN8TQtCSfA
eZPjoa/LRNLysVhboR+DCPdpKNCPMnoIYmqR0fBmXGDD6/rbO16qM5MQeAyVo9FiwAvfhavIVflU
WhhlLBe7cOnizA3ATFpWdr88ZayJM0MzUE0WUNTKotZRcR4sgmLC1gtvXjP1jO/iAl5MxgH3gw0A
kKKHAUNsqlxO3+5nOFucLTLn5Cbd5w53FzHWFRcJmi6fDkrtWdrYck4YI3VFzdUjR2dqrXh3y185
qYBLV/uB1EBsswB2vHxU9AeCB+GFytwQOtZAI35VBtiIheAforQAF72eu1ilV+v3Qk9w+GeLQ6LZ
ta7MelcB55TxFSTuXqzboM4uht07Gm9T4T8f0wk+Kl6iDOdc0tkVbzBxcqzsdPTS0FslRdR09157
KQgVHz/TyhwesEFqLhu3VD3+fP8TdSvQlgUxzFxtHCwVXEDy7PfC8aHoErCciV67iGxRgtmCvpxU
GEk5rLeajzC4m7fnzhlNdeRs9oiywOyge4B6e+SnDFeF9/wksx7bSEX73LV3UVPw2c/6hs4nLHIQ
8c6mFTV27xmkoQmBxf1mUx39Kb36YOHj1DodBn/pNLo3kx7lRNtUpmhU3sI1l+to0Ar9GkH+4s6L
DFHLdBE4P2NWluNr5p/CoOiCtSWY6ISAvPgR1bdYH2Oz+VSU9F+bs1qlSpj9oCbnj7WW4GfZmMuX
EGPMEcsKl0cBUYCov0h4sL1QyuPOyheL1Vlx0DTePZezIKmUSjvj+NZhJnGhNHjo8+BfaucpUm+9
tcSuTm+uTT3T15EIVXu/3xKij5mYOmPFHQV6A7pRK6fatfwT/KwljR+liTWmqhvBfw/10T25Y24D
rEaKVA0pWHNbmkujiMM5d22qLRAV4/keRech2Dgdk2sc9y2yrS7+BMqphiaY/peF5Xb6voe7BV5T
rXtCvJGk93pNeF2WC76hK1ZH5hW7xjhGNHebU37z0wAk2QtWGvnEP3wgy7XTW+2rVSThjyWetZU5
gaZ6o/xEGOWTyoBd2gHKHD+EHKkESmMKl43OzkcaKLulwjoNjeb+TnM83oqzYyXA+OCBm3XwOr/7
xnxIOB6ImeGnCN1HgxDk2nl5brtfUHExXC5a4awdrg3DgIgRzkslkms4c519Nek3b4vmRuPbN1sA
MeMNNSKtN1G8Ij02+dSou5i7u8NozX0SlkkVIuqGVnT/Psbv5OT8fCb7Xf7clC3mlFWytp6QyBGa
uLwUMjR7vfvNbGXnReh/xvPQm3S3sZU4hD5uHa9QHig/izKlH+5tFoFgF7Tex/7RCD1LVxskPh92
1s5dmDDtk+59eoKncagSne5pvtzKtp853NSUhdND3LHJ9yyKG1ZzXYZWUexhFm4zSyS57VKfqYc7
/uWCksWkKkcUXYlnfEHal2HjXXTBM/mt/RYOmpH14J02eOScfKGNB1JfdPJqwj0C5YzaFpEnUec/
/ZhpB63yuSf0wuTRQxI172sc6eCRLsF38zcaGZww4PvsTgOiVkFCw5f1L2VFyCRm/xf1/fk23uCX
D0/g3zWPB4UxjAjBtM5xMW89tO3otjPkaxJcY7hb3ZL7rhBBwe2jlgQkJ3GqMl+a6KQU6RzgahYG
MKEIUUDUiIAyaCj1Tz0HGJSrsWy/jkyLXfWbucAMd7mBgegNiwiwXTwXnQLlWNI4EMS7AwqnJJvv
dgsZ8J0S+Ip8mIk8FJ180wCzsC+g6ZxoGNaLH60Pl9H0tmE6+j+hHxML4R6G5U4Xp+rieI9CPWvW
1C2ZXPAdxtl17kqA5rayCiRf9KCHphi0HkyqFytMfZ9hGqpCPHl9WbAYt65hW3F+sTVTP+ChFO1e
PCBOBcSa0V3MB6d1/Cw3coD5YFI5XjiONSCQjn8apB0pHxubIqaMFg5lLtlKAM5W9P1iBEguvGJS
WPCvnXnkBiuVfCqd6qYJC9kdhD7QYTc4SjbDVga5lg9sexykF/nxQyjTNVzg5CaRjSdpkaMffEl6
T1I+qFT4hH+JtgomjJfW6DXRdZLrg42Mz68XkYMfE8i8IfbawA3GNoxNH5AV4q11dZK/cySbNeRT
WkCR7h0HrTousWREwWHH2VXatRC8ccMo9K87vLLgAzZgHBNVgJBT558a5w7PP8yVyHQx0QXqbdty
89d6DilrIV/XV3Z4bFbBQZ+/YiMq4Ns5kvgywigGI2lDZGaTtLTt7ZAD/lqQYilzLb2HkmB3/AFF
V6MYOGwcwTSGbkpE+6sJDT1wvNwGvdJkFalSydexcxIDwTXvWjikPj5m2DV2h2KCTKF3l0Zbm8K0
2584aEg2GeKQpPOD8cKmU0NQ8PKizQqN4f/iDbIiHtKf7T7yCYc6GYcSrZDcPJ0HYUCnim2U0mBA
Zx+2oeiTjSS6h0QuHXWr0XgGneJxTyBTcu35khv35Os6P5MZGewnnAClC9ZVo+0jUhFtUfTksQNx
fq8k9h4xQpq+8xlhGEcRw1oqT/ffvEWUTNmk4Q/wzDzRrZFwLGDTmzjArh6jzZg3o4GupmAu+mhr
iDFyTCrhoCE259gVYuiZ3yvU1Xz/dKyksJPkiceDQlsccbr+Kzhs2ZN8sUOnHr72oYjnoxtjd8IO
Q4/q+yPNFagxcsSFmGxo5MscVjIGeDyn6quY3UcnmmKYtwYddHt6/v3rE9MgR6q5FXHspst4GLZd
O0zIFk3vpwKZfpRC+XCDPmdIYNFwELmwJFLSzX3cbcEZ6l73IcXRuRT3Z/XcpZzTSwBjugtnRmxU
0g0rbgk881CHm+rXV8FgRggZcgLujo61E1dHIXaPXJqTVlUI79NG5VSfCiuISijfjJK6+ccWtoGR
s88MXTJCFCPA0cbq2sRWh/Spl1FjsSo1kJXNE5us/Ce4iFlItkw40smD+4aZamW4VDii3SJ+9PTO
LR/bcbjolZq302Ra0t4NluamDVxgL6Brmsd6bUf7X37BBdjR1T+LIEHuqHZu2jm0niwaNAAoUUPV
O49VEc0Mf0LXvMYqQsLGw2jMUV4D9HbOZ3q8uGfVx9+GiwRxM7jSS3kI3wJ3F15BuQsElReIwBr+
DSx5+ZKUBn3pyA2Ri/UjVlt9d1VjRNdVk5eqhQRn0elEdbrbphhh3kQKgMOe5JIoakdo6sSn6/WX
2+sqghsYmLgUSCSpkkTjUl5zJF0eQd+HQa4F4OdejLxEhOBSLFgZXLJhsxu7HOnpfDLZ2PUjtetz
fsHy7ZRkyIshBIuhbp1pfx5GBfbNeTZTA39FN7X85C2Fbv4AAPooftwIvVo4ma7HPavum0U5EyFd
FAIGEdLLdHKC85VtoL+BjX0UtdkUSZUjbbeh2FNO+rUOHfJNT9nhbQHDi/yUpKtqGsFQ4hm7Sbni
rTiuRWQxLuOo8KRSjFU0AED1QTJOLGi8e/doLj7OYtWTNS47+L8Fcepb4FcKOza88F0nhBltReTN
U11E8swH8ZOtW7EN33FYdTkmMoHPfNw27allz+03/vLV8i4n9caU3Z0QhU9e3cvHb+Hd4iIpQ5XZ
izjMesttiMqfxk4Hf2jwepEQvwqH+tFGB318rfX/ytFX8zodf8gGYEmVtffoGmyGv5vTMUWqgmWA
/Fn7iGu0z4UgbDYC96K9drBh/IBZpaZZvTE6srDSkfII6dgC3Lhbj8W98oKWEcyjmTYzwfI7Mzfo
u4Jpz6XHI08EFwI5QUQ6KRnTSmW1D8czfKhol70vqYVkFE9l92UPsuQkhebH4MAuADdgeNtM0aOf
ouuHHM41PKA+5sd3dxmDfTJJg/9gjej8Lhu6QSETt9lFLNUXN0rG6Gwcbzw3lUXg9noT+x28JMnD
k9jrnLiE2i7UnnoY/41TmxB+RaK4wLeiRIV72DJ3Mn7hYcVDzYU8T2KgXRAsKQClSsvt9IBS7OZD
3jQ0cqj4Q9rqzfhz5LTG+xhQ+uBby6pVNLDwY79bEbwVWovVC2GEDFml9hjar2bqhl/+F7l6KpQM
4B7UL61iXfXDQQoFdnJsGFhpNUcJItMerCEx8A96D2TvBw6RBi5eSKlXcKT6Qi4zUfOQb9Loou9P
8m1w93D0NAsMwWqzBdH1pD4dS5JopkIBEcj+Ig/zS4Rr5krjRTsXv2qbq0R7Kdqx85FSjn1f+yJr
K8Wb4e+vQHpHkJyhk4bNXpWm0ZyXK0r4HQpj+0wOVSkQdftyHJGrhk5P2ccFxfLrNlluAHssxhml
xvZAisXel4jb1MN2eXNdyW1/cRbxtuSnm8T4VSFPcnLvR69zEusckJdpLezxUqxg13nD2JOEEBIq
bX8JVakaX/fdIX0ct+pvbQ5dlClUn/fp02MlHxxmtGC49HKlt/Y30nTN44t/CNCwzVfOIPlMQXkt
L4o65P5w5rkHnBK+jMEEyYAQqVjVZpwFAgpaoobdHxdYClgu1/doq3JPGpMCC/Aa8vqk0xYtk1+C
IQEFJKFo/yCSfp1uNRB8eYJAH2JkVvX42ZymovHpw1i91hZoxtnczPrwPvYmoiJX8JzeHKvkLilq
ssa+YE2vIpw4ezizUHRoZJC/siV+x7CVj8h6C6Wj15BQc86BbupnIuiOBdumCIc3itynjsXOORRJ
0ZB8jmStI9LGTXyZ2hs8yC51t5yo1bi3mJ0EPC7Oawu48mUEpOHKlTEQYcIq6pl7w2AcfOkcUQQO
NFk9PXGi8I+9slfozbOqQkvFmMsGGfoseM9s9gAoJCj7HU1jTKs3aLL5uvuJWx5WlnPbsF345Tiy
PErPlXJU/E92f4U7kuARlL9bLbzv1MxytIAgnINyF6i08yqWlSTQp3lF2qdw3RwLD6TzZF9XSR+b
ztsBkbxeiqlyuRYzAN6uQuJdClZIimspcp1K+V/0ZWefw6RNV/4AJ8+BVaLISvaQsbRXkfcFPkjl
7fTvwrht3FMMaN6+ZFjO5DP3hjpmKgF62al8aLmt1jRwXY0o7q1GDBOKQTrmdRoyrPKs9DxeSnzW
q8KUxobp34wfg3pdrbmpDN+hSLNwZ33QxsrhhcmML32dUEe2mSeW8CQXexaCZD5ZUUDYwNkRMXC8
dIwLTv2R9Ss0sMAgNEK9a2yJSCCGIqT7gkPh/j0D8twJr6V0GPneCQbmutxsnaJvHaxPpgJGEjFA
PUIg+70CZXh4e1J2f2ccR7MLtr00as7fhARwu0tWlGeEUr1OgjVF/IDIvYKljmFwT80iGRo7Mabr
sr/oSwjJBu+Lf+Fg+rcbTMpdb/wVkyIZaB7Pncz5uZp/0ECAan8Ayw403vTh4RmZUyfR5Jle8J3A
C3puGlGPpkiS/nsx/IRa/paECicX5MOdFLTgCwr7GYhPU0EMf9IQ+oBFI/O5pJgrX8grso8RDwyf
Zb53DKW9SPRyzMee6gaQ+IaN8clrAB73B0yq8UGhQi5pDREEFehw0y9qWyN/8fZ4HvxpZfalo1rk
Sp5DsQ6AOv8d0cQltDTwL+VjUjwSL52DkmVmlQXb476wgVbL5mMZBe+0f1YqEcaWsBYfzXAl6Axb
e6ym/ecCQcxMEh2k7HidNPJmdoVAcmv2ulCMNPlBHSCNmgxM4PFJIRkq0f/tFKlgDgXnK/cKw5nx
cw3i3ABvv7L3z2zfzi+NhT+i1d45zvTe1kPv7gdotruYvflglYY6Ij39yAk/1dLtnTHAHPuW5+Wn
IyLDJ5i6zB51rrJSvjVRP5Gv57Xhjspb+IpFaP40T9KRVOhbYH7GGRwgChbm6M0T/WX3ypur3Jtc
ZiVDegyZ7QL9exZcHblNbf3Q6KAGpNVR3aqRBOgLMXEll0nq/u2lSweDMKWYcczI3khy/P4IEJsx
9W+EDKKWqmjQwEtUJisAd4qF6+PCZxg1ESP/ne2Qc2iOYE7MyYUcmC7ooEHHDu0NItB3VXidFWZr
jhCVrY/2P5Jrresz7T1F4H8VVGoObsDr+aHGUuEYOx6xzR0z2LUaH+tBIRXKlrkUeZBshappeY4x
0U2SRPxraabf5HkLqnlnB4Wz9lUMKaBkfAScMXl74tqpBrQS5pGJazUeuuber+va6Xf7EApPpgzf
v4LeZAJ5UBSlrfmhMEFk7Wye5+uGtE7C+U8ajAgFTIvTwR/3H2ri/7zu6PsLZMJQ8PNfhBAg7wQb
MQShAw1oK+eDqqRu0lzIVYYqcF3MWnET43jiohPH7NJKNSp2q+ATpQYPS4Uo5wkGRAFrkHwy14zF
m+O+n9iNtE6x2N5DJQsv0Vdt+nqdZ2m3+wawGUcTVc2Hx2SL3d0zw57ic9Odmwq5IW5dQje+K5d4
kVDRYiGAtDH+tLiZh/mhMOBPC6noFg5pB66SDqjDzlLIrm2Zdhk1+XGSqwlX6RNw9nkaUoMXI2HZ
p4b++uoHESxr1B8RwdpCmutqlxKffFiBGbO2CQe0bMjECHykgrlsNsjA88ZDigI4J6V89OPpn+To
9hgtdCKkEHXKgxZLWUiwjA6UKvxQ2bfvCpL+cXQWuFlOKz2LgdRdJ8NyZtd0z/E4h/wM99lgZTFz
/BqKpmxxtteG5/EqAri74aVaXQRyiTKIr1kTUOlwQEhwU4G/Q13oUUT9990KnfLIkNmPpyd7LYJ1
GnPUmvw1xoXwRxUpY4ID1z6XLdAY99ZO1dLryi6n/GcTz48Ks60MrPyt98Az/SF+ACDlR3OL63iS
Ok0PHB0cBwGNuye/uoLV8vjqzYdA2GVa+YtdFI9Qci4GSlastT2mXJ/98rhNrYdqjsX5Gogbn87T
C9aPQCHTL2j1ubp7YWI/hjaQwq6AsSKrPXwmiI2oAkNcWdIg7mAu/y07L3RZKMqTfUTjKieikhf5
O5pRF1SFj0mytNvKPNIqfdvyG0bE8Sra8/PLs1ToAV68LcUsEvcRxJp2acB4p+31Pm92yV9g04Zg
OAHnkOFFj/c6sFxnVHv4rODekaBn+irgQJEgv8wphuim0b2Ly0izRC4gQivT3nsqyxajkiIa++0U
ULU+SeA46b6jOTM8jgSXngjPqyJ47pzIaCoZmtGb14eq55QrsM7SO+SR0ZfZn1NU5bIL1NiFyVLY
mY9pELW3VtGM9xgNKk9ORkcMSQPxfOaCPo5YOkTIp9GilqR5SoHGrJhkUrtEpKosAUekNFfMz5uW
eeUT9J3UxDoKWsq04DY15x6cmb9n4DnBjKte4Hvyzuq0Kw4hzmnPbBzn2gnZyRLF3DKSHz58TemA
ueXUJ6urzN5rPm55ssJw5u8/rAkan9ys5+xNkqO+h84OLzzw9IR3bo8kmlJO+2uR6taeiJQVP2jV
qK6XLlNUFy2bljBs0oCmno1786cGliSNR9MEBYGC02uaMjiZb/FMuAtS41k5xYzgnqJcQDOpnECJ
Rg0MGa+Ws7NW6Oe8cx+8lH+3VI7yKQ+LPlItFJqKIIHL01i9qqQLIQ9spZUXrN/d5yIAX93mGl8g
pwr7MhdrM1IkyOzCSyujfwN6gks79XdH00yW3UaNyp7kMysWAQyPs4Kyydv4cRhL4/m8ZePxK6pu
or0Ny8nXTHniLzf9YdiQRc+SA39fkBQdA/4Eks127MY8V4r28/BuhbaL5PdEZUL4+m/++H4ZstX+
owl+HB8CxKL+qgjZJ16NnCj73J8+hSWh6mg073QYER/2NB9ZLFbgkeP2rnA+/wUQya1eXStEYA64
2axuSHIjUARLxym+opEhlF9svcYtHbJZGCbd8n8lgrNQjwnUldyLmQsPPSKgYzHwHje41r1aDBMg
WUvvDiB6mvKZ7SgvtJ+IKOzDe1f5yNzx3BAe2mR1TrSXkrBJnJsrUsGEB6wuDH7dYzP6qmwq0NVi
MrA+i7pxuod1ecBsCkHVUrTvGMgxxT4RNreS8Y6/KcyuWC5eCLT6vag9HuTTjqN4JCZ8KiMiVesy
Je82AA/FI6dm42dv0Ju0DKPC4xvMTPPdjcUOJCgYOeFK1DZsa0p5PMPIwNdUR1j7eyVkONEcbs+1
g+rvWBPFmJ8WDs8nuF4ccO6vTYUg24ydbjBs75gJCyS9ABpq2vMw3ggry4K2YaBJVkX+Wd6heT/g
VEm4PTXCXWTyPEvYE5MwkRkasPC9kZ6x4ePXTOOn2SzlGKlI/QzlGQ5llkldbMHZcEaJfWy8wHM5
0R6CSDr+sdCQB4Z57DQcVVbfJsS1m0ibrrKhtUvMhYFA3eoAXtcqiqUJY1G8FqEMqBwuRak40ce2
Urw21HGFyy9EdIPazDdOxTtP4aq/t7hH6gIUYguauNzSX1d/Ir/QQVSi4DgHexxqxPB9cPaAX7v5
0A57Vl0/E7KNFOTxiv+UXAS9mmmm5Ty1y+fimfEM2Ue1+qk+rE4SZZkUmh64JxxUC12uvcLKZYJV
LH+2Un1Uf5hpmhLTMUb1hoUBgHVW89T+Io4lJcaxHNlDMerqCJr5TBtJNM0Sgm7sd4YVM1CqW74c
eOFSdnSJXNpRVHQN1qFkr5Vj4R+2Rqe3aMRb5JJiw7v/NIZMn20li56YDKGWJODxyezOaVQt2sff
+xOjFdVVnmBawFtjIr7BrmyILALBCA/cxEWjeDCFsWM9b4QA+/Ro++B9MqbfoAtVbK8f8YSvEp+k
nCDtfWJVGR2l+smo9FwJgWY06lfmebFbBb7vBp8/sRePa5mbogsNQ7m6UK6a5x0BAwNwgE9ae/Qu
PTgJZd35CUBok6vIIqpVNW26TaWMUh0juwch/576Rrx78bqhmkCT7L8Y+xTKLkZ8Ri8qKVeDdR41
qH8tfQKWlft7GIvjwO+RxW6WjvADkN29VoA7cqRbBNQZiGo75Wy4KTSyIionGZWUYiqIA3XBHbjJ
Qrd1LKr3A+lCYnN+jrmC9VTckOHDwsXo4VKVzIGZgk8M+ING4DLqjyGGpeuvE80FyOYzV8B0U0EV
hM5M1kYjqtOqRMC66byvY6kD4tRqDgcMflJj9P31HTBqqYRnRWy0uaM/KOvngYw7+Zr5Sc7WVXKd
43b6eM3E1fXFpcFMJ+HJOpPAyuQa9LUICC+Eoszcr9y00t/AyJy8+2N+V0u7lR6t17m5GTh1xCGo
90YhhqNTZU2Cdvu1DYvtImDLgMM6n1K+HyWQUwnLmrXm1CuTWk4YrSNIuJlTBkc3uFxLE+AwhIFG
iLPNq8fDLS87JWnAtCEcb7vTbNq/sxtoVCgd7ed1RxRGat3gf8uafbo5wVFOWcbp3SFCqPlyH4V9
t9mkpgSWbI0iEQvyAGdXpFvc8zmOtmFLtfotzzy5n6GXmAGB1J+1NHdezm/ocbQ2XAdqbMI9aKyo
wL4b5ZF2QuCW+BE215pmperWOl0RD2HpFNmvFQRlEgvr4KFa/taOq/ppYcV/kOtGLNXwPDV/BV13
YpPkAQV+e42M+jLSW1B3sOFsq1FwHdwlzUDgZvzw0fYECy1VtdeqJAEBebJRTClPx5ASSbdqZdax
PH0DzsBJT85Rrjjl56NtLF4p43eLA/LvvJqnECwKQoPazlQ063HAOPvYCKvXJ/9r7xWf2sHqKKbg
O0xrExPXcYD9TyTfHT0C93nsIwN8IXw2goDYZPDaTJUWst+D7hOEvCy8E1wcO1Qn604GtEz15R8p
onvzpnYFo3H4viyLDoVb5054qai/vOBQ609StTqUx7qdKObIPIYMipAagLbZjXPGC9zVJXPdEAlr
nkJ9OtO2x+kV0FzMupHNHHsgFz92poU0AYFCxG+GRYzc1zf2yhNF/Bgi2RZZjl+ifKW4VsISKKy1
GUBVnQVtLK6sotev0f7lcVZUKakQK9JEfyOMRiUQ6YU/q2YwJ2Df79PxgYE4oPaBkdE1uKL1aM6b
9IAR4TdqHecPbzfqRZoQsvUtYl/1XnrSwGMXKo79IKn9M4KwbREicyV1OrYq9HTXBeaMYSNjK52y
yEmnLbab4sjeSIFyVJnDSe0dXAZ6sK4OaQ+dgYDdsBIXQHZxXQfuZO89y6OA10Q2tC3z423iOhKC
5JO1nn4jndAY4k3Ks66M0Utyc64hNoJtt1AACHQ7CWK4VLjh092PceUJkTPjhsDWfmmY+tpVTiXg
s+7/IKyakqm33gwGyDcILKYAl4etoVx9ubTuvUTgi5WYSCki9Rs6J1EG6rxUr1bLVa7Atb8Dl3It
a0juwg3e4T8MBTrYyK3g7c0plyESrBS80K/UwXdx4oUki/1BpAMsAIE4U0ZPm5msbA0wV5n5ctv4
4Uo4wWpQZzxqsatg5GjQ1JByXbDTXn/MxX/+F010bcWLsDgIsbrrqyiuMX/ZJPYVFPvORkXIxd1a
8yN0LOuF2krnly4VIxNJ2eodRWS+tWqoTZAlCHFI39uF/V/HhuOz10+SA5aUHLd4pmO3WKl5NXMY
3h4GWs3ALcgi8s4nK46FlIeHcQGN8cg17+p3ZgO32UUyHEu2LAASOU5vSwsLGQDVaqg5rFzud2j9
g6kfEzWT6WIpsVpT5SG9khM9pQwhi33OAB4K/LkDxNANIMzBvGpukuTwliUiXBdRF03QGpMdnYv/
dTcQOuZWvRUHj3eh46Zoi3Knl6kM1PQmlINx2jqtCZ7Nu51G/L2yI+5hB97YgMW8MVq8oTL6E2EJ
miQ3Mc6+IxB7SzlZ4SpAPsac0hZRPC1m+l8xJz/nXggWwvzbPMdrtzIA1r298S3PcT354nN3lQh3
TR8gVJMlXnRxYnw3JQS2EbFNx1ki1aSfVtY/XXdDd62Kyf92uxyqjYRmtmcRChdbmMFWKggIiBqN
W4P2EicEf9JT+R2IpXG83/kIZiCzOxoMGgKI9NpxJUxcBJyRxuJaj7yLKskmVuReHnvYktahBt0f
JrH9Ly5+KCCSOVGhr6UdgsoSXRfuuy+R5tmFyUhBMFqGLroMNudMIbsFGS9S1PCT+ceMJBZoyvyQ
JtNlRqZE8NjoWVafzQgwKRxIa/XK++D4q54+lJnLA/RCMst6DU3HYMYPBGtiozgAVoik+nCecdPN
UvbpOJmPdYf8g6AvsCo34loETB4M0mqq0NFGmPav0jC9Qb9ZZS8eoL8Zq5J8x2Hw4K1onRCBiGhV
ATfSShHXsd5REA6x7fnJvD3pBCnvBfXcmnX3mg8L7e5Ef3Ye3A2JmeJdtW6LOTSgz8sVLokZIJd+
4als8nAlb5juY2Mw54TKCEPYfNtBF3lJ1Z4IO2hKCUY3cIoSp/LzZAdg8OXq0yrkx16u7+xWU2Ur
yP4NhGm+f1pFONvIiSvbFSSPXbFNb92OEF5NX9i1vH4BBwzqidVLtdJJ/52i0x3BtrkOhxfyrMFg
zRduHufdN8rQUXnrhgM3huqlbVXJhXj8fdzoWwZyRNRdvcYqUzz4X20Hr+MNoqTMEMfuac+8aaqw
TGFcgOeFIyUSsBFayB7XyOx1gIh2MX3yLtMI+zs68+FAs2LmEUJoTDLh00u/JyGrf116tvKlnF8M
qjWZv08yzbFvquCrwRVxdVZaoXkgbcmvRt3DQB6Gkh19CsgTDtWLeyu39nscU88Ma5SW8+avFD5k
NZFOEHsEmzh78XhM4aAG2i6gD1F/IB52m4JW4wSgj5T+MIZNrmTcLMxXEThthWY7AVgrooZDS240
lXuOt0a+MHIAojM/1Pb7lmTZUSgAmlw/EkE7DKbAU5jvBg4cpHLsOvkap7lB0uu6qDYCAd31aGmO
998EmUnHOMySLbgUdtNotN7R4erdGHPLGi8NQbnEYU5XtTpwD8oeRd4rHNiDTDHL2kX+diYyllqV
29zQ/FRwCGgqX1oBy91Jm2/diVauQwMN2821m9nDQ71/rzOYSJ6JQskziOy861tXSyzAg85KDG/R
WO4E218fEgefXQKcvL8TKcjKhwpENQ+99jyWv15AzrFU7HfGxZU8OSqJhin8kF2mC9EYpOLJqHcd
QgQtjtb+c2/XKJBMcNzOmElffT9bjWJWBiwzCBg3DB1oygW0gEtxGahk/kNy0sAvevTm0yVFErDD
pSn0JyTrrQyuDNBDuAZP+7NqQZrpjigHKPeLdlHHmAt2qj4sNKeoP3QmFf0X6jEW/JjhQIB6NPjw
etju30Kkr/NsXnv5ZSkuVXVRoxtbGW2wOtmt4BM7e/DSKGA9a8OAPSV17QSfU2KtyOBs+uK612Eb
VzMhRERDzFKvL1gqwmQguet1pj9jNxzxhdbQbaWD9b8AvW9cx93D9rvC1wgi52Brwv26ABGMpe/J
MYMXzzLx5K8vAF5XhXNiNCnrvT9HLTJhy2nBypfFRylj9QAE/b1++FexVjIw2MyGZ4XJL7KPrFNO
uB5qiMDHVSpipHMEZaU888R239v+/Hr9UiqcmCXstLgJ1ukVOiVm8FYH4wS4c6anDAVKscexOqFg
lJuH9RdSmlCNb63+nUOxYJvso9ihmAj4cLIg0mLue5Hg/ylJ9a8mNSOVpNhSwiJrAqeBM/S9PWiv
CE0lB+AnWs21tV22pJADXfZ4NP+1DlsSRQm/oV5cR1sJ09KHp/VSYfvUY4ORtDCvjIxcE3W4i6Pb
kdxw8SwbxrtOkw+zalUIQATPscmPRYbvpWvjxRmIQuyhsJVVYY79YxcRH2H4Zladq8v+6J9cxiaz
oVfMZLnkQP0UItUqFbLcVuVsgFzx3uZAlrDX20Cyjj0VL/0/ms4pjhZ/D7WNWL9zerP89aJWooPS
K13vBs1vRFPcP5S5TLU9nrURUHN1oNodZ2LCaAOD7otQSKjmVOEh18qe4DgxnqgunNajIEsnPJ0H
aAn5w602vRofHw4t6bqpFYcH4V6CTzGi9e6LpilZ1/PtuPNluTNFHJMAvn3a+EEz86QPdTlJ7vKL
eaOoGR7dUGBTpu8zn0fxLB1YLj4ADFN6gFt2G7FayAit8JAst12fFQSZaEgid3gh1pOSCTnaqyXK
UATNERabYcN0JfAdpqr5IJYD3K8a01E+S1h+ZZe+eJH8OkmnMOnXc3pQwWW6UKgD2NqgtRnC/d6x
DQIkvRY0x+T6Y48b5KtZZmLBPet5u8YY8C1e+if35E6rK2kkoIaD+LD5HypcI3tS33E4Y7yI80BV
AqtInaVb8Jjwp3tYCKqqKzYYS+uvSTrNenkY5kJUvQ8eM+AxM1vWG1lYWk7aRqiJqewe7nGI+Ijm
Nj5MDSS8OIJL2aRWxIjujS6jP0K5p3q8rcoiOV+IeR5wSwTfENCeh1HeUTMeHgYi5dd5yHMrwhcP
gNwjCvLQ3rT/RCBySurC5htoosqSBR2/X4t89jEW9FOQfWVhMfUBZA9j+UngvYlbZzr6Azt6LBN5
tFtzm1D+f2vpRhvKcjCQzcSIANNfs+6EVVwO2REfcQtwd5Uw/BonZbShrDvu2xucCeOCzPhFjpUv
tlBonsjbZGjpXICusPs/dMyXkmD34SdoNAvNyUbde3knjJiU/AOVOMXDQKHGWRJ79UvzMnepyJOF
Y8Sb2eXcL7KfCTFDfwm0WiIcUSL7kkj/zBtDF3HuppvEzjGb96dEQpWtdqPQQMXOxyFP5bhkj4An
ah6OEccnIcGzHkXnXv47RhkBsmb2pF19zTF+25eXez96T4QzkCvnIQgCP1I2RdtgcYqaif2kzIJs
EEHhGMuQqXlZAEtQb+bYpJnd+UCi2fEzpA/irC1mBRval8uZVX6KoIrsJkE6CARoGBr43shYGGLA
IjvYmP9XFgcnaw5C9XRYAl/2fQzSv4kUQzZgeaVrii/tVMaf5MYZImCL3foT+JoQDTDa7jCXjHb3
xOcYCzcUdSYx2xU3/yJaCzTpn9rjWpZWXiL9g1rRo93o+v2F10dpd4ufuQwgI02mN45XuN2jBuX7
SC4dFQ1oVJPy2B+rH+56XzaAeM3cmI9rqsGG2pAmyB5I4FoWY/2f7THO5o8aZfny21od146bNA6Q
3cRYp9sw5CuEcgZO/K0Lk62giDVDLidUQtJ976YBSsQXLIVp6EylXWoKlu83GsPcIGWhryeXihUD
JUfhuu4eFazrBqxt1pozrd8rFwP4XqpG2VBoxTMe/x23DQJjqs7fMaQVn3k8LkwgsCs4cFq/Mms9
6IMD3mO63/13CxL0BgQPAWZB2H6WS9+wYJC4lFq5LqFkyZX7GC5tKB5LQo3aW7sqJUnPUSYAi2y0
TvxSapUx2zn2jV9XBhQ6u/JGuhc31wPkxArOTwr6H6lqxW46BrX20JhSVvwvSb0XC2TUZh/sS8Dp
fwR0yw1DWl6scTWg6r7R45Yjp0P8jGrtRN78QgmID9El69JOTvhTQHdTfKma0IQef4qa43q99QEA
hWjowr4cn2Z9L0r+xr/VCevQtl6jJnfwn/Kiv6BCYwMpcVGOmjTCuYEr2vviibXNuzSjmLGkJWvf
/SS/KkpnlwdnWbQ9AvL+uzlmJZRxKwrw3R04/62LTLrZihidceP+cWChtRPQYnQPASIiQbMirWw0
R0xxsvd8y4QwFBEufyJd9/uEJtqR2jPpjnTzwZHUzRaPn7xy94HqzZBXsjS2+9JS/7gDfy3gRTVv
etnhAIWD22HagWeNDugD6dhuFS88tOzEotnSjN5fZN79XEFsG8Fr+r2K2jbiSqWXRJOkjIf3qUDW
5trl+gb84j7dhaki6Q0Xi1kPpzSV4vtWHykBgpzMq2TH39tQ5wfCztp7MU4jUEF32G2O86HSwU7c
OgGUJYo9toJyKzc2vnukRbmfz5D+RmQ9uZ3dw/JbBJwf9EjgQ34SLztik/29ETHnG18Llv6azK7W
HeY2+5L3a2EfES6WDdXhc6Jj+gYdePScIxaSC82SHDZYL0RDGwVNMWlaV6bJZohTv0cEpcuoZ89M
LrUxyczuNauA3mxTEhhlHRtJxc3ZC5981FSv2hPeEvREruFxFGpNyBkvpkkIq0jGaQxupl+TS9oo
tU+6i8GLv1+dcpuPgq6uulK/ECULg3UKxhKCQzvBhikXDLzCs8jGGPXZnEp0OE3dTzOM0Bsoh6CZ
UuWT0NxTyhgFNwRNJxtdwt/phbXDTavQYFlQT5o3P/iigmNrxOoteWT13y22XFy9zHZQJT88bN60
fe++PaPSvnLWuh7+WHMpPfD7Pk0wUisHZ5KvqPyTplBRAjM1Pbe0sr/RsZ5q2yLXhGCWwpufYp60
mochUbVDr403RdEJGMmWENnimIpbP//YNfwSVaSAJt0Az7LmzzoO8mcTSiMhl/1XwQXxqSbemm7c
4DyfH6CLW36GV9V+jkDyw3URr6+5g18LpsSb+7lFCvhlouu9FBJGzygVk9HkIny6UZoxi2i3mdel
IL4InKBbV7QuS7NQ4HPMKRLLxg5qhXWGTaGTQ7hdQnXk7x0OhDGzobXGg+S66yJ4bpPaU2qdt3RN
lw8LXdvz59ZJe1nK8/mr76IL02d4dwxdqZaFm4IsfVHXOpY4v0jIrVnLZnPM+x3QTu3+9SaS7TNh
UjRxGleAp+w622PmFVwrG5/pqzv5PnsiyJKu40rGFgPcgIcpD2323ymrpJ95kz7dWwgX6feBHuPe
jwqhUPwN0r90gVXC4yN/w7mPzvH5Re2FPkABRLYnGRk3mfUH1MpZj0uG1pPkp1sXAgFLoJfknnCo
OYWJSWjPwTC77iGn82wGQUnE+I9+RCAxEzeZW1nTRZVTJEmK9078KnvesVs5eplgmzpHFBM/Bl9Q
u9XdX9zy1cytKHgqEYdyrR7UraoxXQpx+tOlbIZfzcBx4FUhollmteVqpwWh+Rog0wdrchrBFDmS
3/nIuKwtkd0LLKt01tm8BvvzseoouMVdfZ8Gu5CG90Sq2pByKXFtQvmmFDw9pdcFMngiVFc9kFCK
zXWWfJkE5VZZ+SPQHX9a6mSEDPwQ9yZOn6BweSQpz8fPcedsfDTD0lWVQq5XrNfTlKz3SpTzRYEc
KMBW1ccMJUkayfJ8lwQf8ceoYb/yThf81fPxfUT8SiNYdKWP3grNaTUdZ5RB1BexjlSThyghwy6Q
BMTkq0dNmMZ91kxzcadl0OdzF6SKwgv2NySbl/CmYDcox7oPSbOQOkIr09P6Fz+qBPTmsn0dwmNp
/IPmYug3VBgXjojSuagitmR/hXtWoL/42tNc7y1J1kRy4ajSK08JmFQ2veMfJqKazANnX+YDxOz0
8QDC0agjp4VZA6SqXBm14X3SkV/lhswqd3v3L7c0Fyic0fRX4aQzG7dH4NqypuF1NAIkj3MYoa+3
UjzBZsVNGv5+o2wxFkTV9KDyw5B6apRDvsuVon4YVN3FmsbzdDCQiLZmziAMwa2tbSnUfqwtXF0x
THvqjf7kyFEqdHHQIxX1SK3dSSy1j0zTTBwSdrieJCHG9Jm2c5mUTEdU8dkf70x7impNA0THB+f1
HGle2HrJSBQ8T8fLAmKDDt11sJ4e/4mxP9myXyg4fFz2qunHjk8xm/X30A4i+C1EecJYMPx5GkEl
WZjgbBVXQPDegeb2NmtPtmTwkJcmqeZIqfX5xZ+jFYcWd/L5jmXkWbGo6ZY5fExGxDSYxOv18i4f
j3/rU7pMg3hlRSVqcTwVZ0wveQN+hOzwZsf/erv7uDxCy19HhBxYtDfxp7Bh6XPnWxSIijGEL3bH
djgfxxUgTRf1JmG3k834HDh6lohkR367i39J2RF3yeDQXgWDbjbJGgRifU7rX1cHr7EELevZW3ua
93t7oCxPoiyAlV6+dMNBCQDKIO4bVpMYbrgGa9F7i/BhVvr5WXOIkSBa6+MZCe2jGuzjfTO19akM
Ot5AvbxgMZ051X6lxXb0Ma2oRTvvRzB0+CnSEAibMYrYfDurGMfADlUYsNPN73qHnMi+8Ww0A6+X
j853Gb7DjjwF2UDiRBs1jzXTxQ7l1xwiH0e7BC8XSCTyfS9m3UNkcZNyRmCOPjHKy5DkG/R0stfT
/cUKviEAy8U6TneN18o+hEK9+CM/B0y5TYS8qLJiC4nNqKsHoN/b5zkMZ8/X/27CqylYt1rKOwkR
ZIZJxhBBHg+P7ybd/9ow8Rd/71sSW3zj8dlt0bivc5U7zNtHyUJ3iGcIhiUzxe2A3u1W8JmLCKC3
qRpBa29xt0H02X6P9DVhND1AUWSbB8rWTkx8o2it8uuAUmcvJkbnF5Wlz3Bq9MkDhJc2iUcX1QIY
WkbM+tQmHFd66/gPf9BAqUjfCK6DaXWjjXskIQJbUI/LGUPH+Qny7L6bp7CL3GIyd4LX3akb8utK
6szT9/MMhf0A6MhW/sJ4uHzEjpYlzOymPqbtT1n+FDY0nPygrLmlZcV4bZgAAsOpDSKu26ui9gC1
OiyLmgHtixhXrDFh2n8+5Th8r7itPWUaTOf7T2LQgQz6MVCXP5zerEtq8dM5Q5cC0JYj/SpjY+ea
I3jl5SkMEEXYB2WUVl/r746p13PYuH4QlsjbYuBG9pd2+a0smUvF5pRSaiY4rgE+CwLO9VgRjE6N
elkQDx3KLL7xehLf/WNuczuhZ2dCPhQgBe2+JvW21q28c0oppeX1a/K4VdKt0cM45hIv24KR40ap
IGzg058yPTl2QEHBQ86ZI2kVeFbid8Vh8pspF3oa8Gh25xSgDb23oOad0zevwg0rUELO2A8HkTlE
xZGrZbhMdS4L3tsecYjgUH4ZitdcLG6FXcTG4rOm0DYh/HgNkCFS9u6JgO47BuPp9QklLM+Cc1Y+
XeUmbwIp/fYDdTqvYMGnwS1J9Hs/S3CtD+M5dhrs8odqCW7BDuYJ974rZqlqIEpgqtejGxws5ots
fr1LiV8xK7sG7D5iOoEcJQVocXkh78Qt2Q/AqYHoPxWWTH8zonl+00cm8yPplKuD6qqLQCAFe5zo
w+jr3uvHb+VbAdx0OYF5zaCMCKIOSvOES4aK4dhi89MYImsmreQiBimozo8S+YvjI0hr2W+d+1O2
sjbJyJ5iX1ZUhYgzqSu63qIDuYSGh1vDqrwZgp42ifxiwK9VNPdN61WFGm4WLOsXL2dpO74qNo5S
QShaVtsnRQAxZc/+cQjpkBhzGAiv5tFw+oaTcgHesKh64YOX+QiMiZl10ARp6uzjiPQy0HAMXzHt
0+J/Kp8hx0ZsE/hpZduAR4HqJuPx0okkj+R3YXlW7A1vXhaq2iNJ09jFY0DaQxG3/XpPEsWgMTGL
ZXM1Vr02A4NahwiqfPL5ya9d6eG8Yte+Bft1DqRZNiF/kgCNWNuN0WKGcsCtwuwgkOpxbHSqXDHi
Xr0X8bRt+rVUioB7lx/oUg2xu25i2pmopGmEzaK/B08qfbblqijCmqxPu6ayvrSMkgy2N3rjCvFR
gKlMyoisjqcAT6CKHySwdlPZu1Kd5ZUE4msVFiDPnsSV7BUwwzM3AcgMgN9eVZjIDFpkteZL3oZC
cUj1E1KRvBzwg7epjeApLYDT5yUdrgG0jOudbQxdyT7qd6Fie9tcOnX/VW9ie5gaTa1VxUyQYa+P
rR7mHGAFQYomUEkiQEaeMjhIkCBY3usrKylj04hXwfzpgq6UDMhcSNrizIsO/RHMB6TdDx6Iq9GL
U6bneYUGKMd1HxuNWFlTTedJVTJPPZiwCp4yyAsgx+95OiKY+FJ4DjYOFRqsJfwJ1moOS//06Bmr
L+6LssY5LHdljuxwlbxpFeepO4hKEqaMiKFEiv2DeY9ZzBY8SZR29/FuYJhyObdllSJW99zOS8N0
SGYnwOdHXaYHk2t5y8iDDFZFI2/czY4cUAAlo/qT0qIO3Q9j8ykJCVCh3xObu4IBYlBEExjWbm80
z+M9wZDx2FdXwsnIj5LSYoag0v154mFLFzhCiOzABRVFSY4Ds1RqTtwgGbD45c5bhfDbBgAcWU3Z
HeiiWXBLOiCIS2Wgh2MuS8RFcB9kjte1/+yz0iAX/yvucEFxP0/A4mkg8zZSjedtp4ZaTQGds4Dz
UAoWM045MfQfr8vBAzq5vJUS0QgU+HGqZv8xGMILKqgs7pttogYWHTYzvtSOGnfL7UR9zN5D9Chy
WmjV5nJVDpDFUP2FDt/VZv0nSeuX5ZbXF3N4TsLZR6W39GjbMvCc3Xc2uDGwA4ARDt8BEEAN7tC8
CRPtsMHQlxyVvozuCn2Zj5ofkb7D2DSBP5KPCzargfR/ydoNjWM5WYfuo+SFvPCXHK+u1fDKdZjv
z2nAtbf9000YmrO58ytiYvr2c84SbjY4NMncbTLoUfwNYRfbviBIPyk3OC/ozsJN0jOigwNaJS9u
RFT3q4Vr9ITdruStfjZnNAGK+ufP59uF/cnV3TiwIoJW7YWUDez1tYvmwNUqbBv8r+Eu1DbJFIgC
RvhXzwzS19FHGDA+D5NUZ3w0ROeIKrTgy/i7hotR4mROkq6VSfSHcVDrjplPJwdQe3seyddtdEay
F2Qp/8eBur1H01YmyBquIeAc6dptmbHAaERdFwiXp/AVY3/JenETUViwUhbwsQKNoV83u0MT4nXS
3PRzhYNhyCnk2B94O5V1XnexNYlJb6siftSjdC3GYOwPRBsOYk4qomSIDHzfNZKVlrwq6SoAyrw2
OEfj2SJ+wF8KFwttyk90wkbPDxIgKzbY7cqGzgRx8Hl/zGrOGrGZh4xMc96fKntzhfD641JUKN4G
v3pWRlyMGaeEOBqkBSrmK+lAlSrbXKgmL9ANh41hriV8x4iSOlRev0qPFRSMkPHCmI0ICZCxyPD2
mAEVydlahBl9sugWyTcrSjFBYHP+KIi4HETJ4EyiDAvP50sK4kutEVaXi4zjoATEHqXcSCJqmlP+
yYlB79d0HQ7C2+HeI6mXV6SQUkZGQIn/F20Eio7eWlW7CAIiTmxO3/y1lnhqQQZCFxsIpGx/9bTW
BBXXZ5RQWp8sBONN+/7uRfZx5OyQ2dRUw1/CywgaXTH+mZIlJdRJaJ2SgNbZrN/APqTHMseSmyst
Dx6GoSl7AGwBigvgxjRmw3bab0iEHnubOlz1KKux1jY591OyHuZo5oqvOufeYORKKkDDvB07PAxm
QpIzTKSc3rNRPtVrLqssOY+TSoRyJ9PKKHk5a4CwVUaYPtvT/PPBQQ5KzwORc1qMs2RjZLir+SHb
9njS2tSA50pL5CO44fZqDoRKkiUhjAP0FtJbuRzdZLeAECyoombbIXdt4HedVhcR+nKeQ32XWvP9
hr9FZNuh7XBJWc8xT82zD2whfzIVfZZm2k656Ne0aybjvaV4VZJxiIJ/L8rmBYneYIbUeg4Fsz8N
3lXIsIqHuMRDS35j2N5qBAr1snwZixzlN8sbFIi7AxlRiONHy4fUCD7dvvPzxah/3uhFe7UPOlNq
zRa9jeIwpNfVh3b2tmGy0QL4hb73fmLwMf/rXNs0Uv32QGK2A49UEq60s1KOfKMFQf6CkJfMh11F
qDLF+VLiBS2fGqfruNVE9nSMLADR3wXedbvyO8AakWyolNdWb1deU9y4yUwDnSwnpwRxqVaeT3jU
nbNXGIF2+9hSwm59a38YfNUWtww3ydOu1g4rGyG7o2lwxnRCag8aNRjYXo6017eVmfk4BbGas8pP
FScwdrf0F2JYlQAZ0XNNQWYc3WUx3tmVdZQz6Z8hOY0T4XTV0Oci1OprXI93F2tm4Dgr/hmBG6qG
FGrtgM/QDhX5DoJ08BlRzTgYXloCYUqCrVcOE/dSju6Hn9RCjuryB9jOYdZyz6lhQ/DH9b/xq+s5
YzCZMEKrQTB/SoMFf727Vkr0OJDAVhFLEDKAvntb0yCLiF7wH9XoHsDDMnr03bi9hDkmtzY3oVwX
V0GDChQSAsuBmzXv3ilI2TDS8NBvZuw/3cW6EPZhsReDZ9rab7kMcslQhkHars16uz7xayfJvAJ3
tm9moB+TZuUXBbjca/3k4qMvxOXYbFV3clxlX/UF8cKqjb8WR6x/e/WOoOmmNQJ4KxAHM+3pPNkY
3X38ZApnc1jN4cC29LbVpMYf4iuJESJ7Q+dmHIKcLBEac3QfXjCkdiflJmc6VDMsm6hEJ8buOcwS
Mgl031uhJLu2+bTSat+7DWaMB0MRV0JSXw4W0mkhW6dy+DdcaNW1Vdp7ibwDxzuu8p5OJDRymBQK
6vtpuSOdvaasIeM2hmNqyQDmf6MasdZLPkTA5lmkU5DldTG89sDnpYClbUYwgAzFaMCZFHp1LPqZ
R/rH7tXFdt7LhjF5tMHN8E3D/d7kkb29se5T8r3PGiNceoss3VR6z0zNsnFKpXRTT+4S9MLVv4DM
Qjxg/higgk2cWAoufaovdjhEUFohqeAvzPaUu6v0tBGTQbd7rv4BqQuC/PbDtQiDZRJBhFPl5CrF
xtRuQFfQ3clqRTEnj8uhCILLUVCdBaBaNBB4ogx062SNBAFB3pw2r3NDgB+AsSVz0gMlVb0tTcxq
/Yck5afhDoaE3z8xN0ERMJ0YguhTxZgCSztoOZ803rmTmKWLoV+SMWAKOCEL/Lnj13xAzOAjCPzS
Lvrdnj6SX3z47SLJRQX2hfNLzMCWLbaKo2mYjvSJyP2AtPEcbCJHaH9C0crVLyvWtkDynwrKybT4
bAvlyc+yCuwqGOUaM+o5uHwmqEkseXmAhcma+A3npvmld+0LzZkdsTDggs/IiRabx95mZT7v0Qfe
OPL1tp20eNdrCm4tL761nuTmiN2q9l8v9JbozcPw3cd43mMot2Tg6lERlU8XpSIcgMt6xgqHJ7VO
fcBm8TFaTc/X/ONmffXLEnmANlTjMGNnKN5vtANqoKASEc8u66kboNW2MhWbD9xTrhy80Tkk1uRa
lhO9zVdbQxiYWjfeGbOFnnzQjrjZqtgsIsZzIOwlsRYGW+1yFAfjBJY2FxIiJOvP292aa/l7qaZN
61JQgR6kaIUGxuJoRkdmoTllvkEmzw1RDe4bodyrzk11wgpeyyw5VuiKWkKBnNdA6PneWL5NHwxp
4rA0aGnAJld0QUlNCezAJ5S7VjeQSV6lWE6eG7vmbFyT9bzu/6/VFemvUofrH5E21OIxZpROnkZn
YJ8J8Ucr8L4Lxwr8xlrz9jIa6XyzaS5nWxLN+JHgVIid9jmkOgBRIURH8gnVRWCOioVk8GmXboEu
qRCSeDNfCpaPbEVJtjgjavGxkqxyV5o9OqpWlzmwKPaXMCPXS0is9iGd6kGEOf3Qvruo0VksmuBq
tlZKkZCJU4J1KXefMEtSF7ji6b1UXgG4jmCe95yleZfEkRKxfN9P97Xl765Pn4J1v6pgBa/J/Uyl
1L2VZ8AHeGBM+jP+t+6KqbJS/zSyy9DslxgTCzDBV81t5yhJTPdh1FR4f77F7qYIh9gpT9Wo+4fW
HV34+gtZw04KNpkJOAxfkWWvQjkxMJxCD0FkYx5XUnjCeP5MEoY9TiqZSBFl4ldXbdpn2tF91tcl
AuK5g4I1mX6VsbIdHYdTxOegDhIxuJk4eRmJyvP678epKIRPGwtPO4zP0x/X9BAsSC27JAQ3Gl1j
/RWXGfyRywvR1kmAMue8TNPC8v6Rw/19LCAN4rSdX+98laoLKxEeGJJpDJmRR10jSSfKAtOYl/b4
mtZfUYpoV9EIcvdp4RmHY3vxRV0plWn0unmYOpEy5VuWbRoO99kQ6ivHfNgVXoLqhE2fXDpFaHAw
9NBZedLmixtbxTTil5EpyrqSHwUBwpjnuo7klnD6oRKewQGeNqkj7do4MSTzeBgXLZAb5ZFiOX/x
P3s8s/9ObYK2k2OxO3p/8mAd5cRwnj66IHXG3+AEhfUJkWYbm6CqgEZJA4JN/FkzA4ElxcOGzWYt
Gk5WJb/3fLRxrXiLSpBgKnaSKW2UXzbMrUkaqJ6VKTrRfbzy3pR0Pe808AqdR6kFHXKiNaBXB02+
IX79nMjbWriJpJ//c5+M2xotXCGVCUd/MIlH5zVi2R8Y2iUqY8ADcVFOUK/ZQAKAzifHeCTMVFiB
AOeAYZMqEDs4faycLtinOfTHNT9dgqp+g+/FuTNOthcP6B/FNlA+9HeqN5i6ZpvkUdDyD6L0gAIN
gpc3/9cp2+O++k6EB/Z0Y9Pk8Fsie1L8pYHKaZSjSbjiamTh+fnSaOLmpGz6n1jCRkQ2DQhLNVne
2vaO2r6mhT7Vh3ATDF9o+FjwsCvyDtH5qWbr7/TStB3M3fDzsEqY/VnnhkMSftlwQ+wBSuPAylLa
ybhPiTzZWSCWtm9Ly8V4biJRFxtl6gZl0Wpm8KbWicjMtEp06s+KYFRx2c01061xf5iygXmI7TFm
oW4N7wGsC/kM+B7W969iLf+wROth9iTaj5wd6bLzEEpB+eufbixa/A8NIEwavQIE/S4crYNe17JC
0a13X32Kz/Xvbhvh6o/PbG8RerpFhub0Lj/r2HEUV0PJQXYl0vPE8zim4uB95n+XYTdf9IGcaqsw
/L3+D0JRzKrNUx7tg+pjwcX9ojxG6uYXQSXxxxgPv8rFkXJwYTORfFPGd28U8BFY9N+SGysX0mLJ
Ur1yRHkAQfRaKRLiYkw4zWjILeQhrLjAtM9ktcSNjTi5Wxtl1SX3Ky/dP7nZ+f6yO3EIO7X0p5l3
0ousjrNRmx68MlJQBJldVOjlCC6TGqzcE8F8Li7y2tk8ZIbtNMHhGV1tpcmmgcpPpXrArRIclmSq
R2wVkE2qkomkoKc8O++oqleJJOm3QdNNfC51ORSwVBEwZC1qXdFnWLLll7UED+boo5Pk9a6GUtjT
fKlZpTqURkzN18k2yzn9DSgRZXIcHEqAFvMwoCoa/FsHebKF0a2XsC2HpK3IMoBe273BoiKwwspD
4VqDO7zu+HCV4yvaNJNF90oSiR1/h02r5Jx2Sps6ZOuVxvWSpKAr8W8Gf0Mpg0IHCBPGB8KMFhM9
eq4n6QeFu9y9ppQrwLiZlRBbCDZlO/8Ls7oU61tETG8MPxij+mIC5Y+Qfpyihfk5raa4s81UpgvL
pJAx2vm9mH+TEEAL89oznPW19dvEqiVrURkLoxTG4v9pf42Hsy+l74VlFeGakubVrbXLQu67BlfR
wlRD5b+Vh4ubzWDYHdFhzouArnIQM7kfdfj+zSnwB6c3fWVs38fklL5LU3ApXTz9x+dlmtMz1zMf
ED6THRSb3WP1wSh1Lml58YrtXQHdmYwie51Wrog4001c1sLEgwKn5/eWlDREgHsFueSENGxtCg2Q
OmaoKuqCAi0rZ4TgtxzQG38HpYJwucArIK+g2Do+7fPPjBicQEhzPwY1OJDj+Ns7L7+vhNyHPP9B
DACrM5oyXvPE4tKdXZt3YeH1Q6dWmI3mSSreyf7enBo/8CZfdnHUPP+0p/Q7kLc6vzQnUfVkVyFk
hc+yrW8pY8WXA8IAK8dOmNPZtMYUHI52K2SKVv2IsXNKq7RqMlGrgNrHi/8oDaotrS5dU6iP4X8V
WbQkhCQkdpB5p8v8uFBZUlpJL0CJcSLh3CxA8inVRqBvnO8HCdKp+nWl3lLX3s8TssKKMOiAIdZN
UZXC3c6qJB03lyhepb3h4aHO8RPjH9Zpg0OAOf/vrYcQfeHJmgSczmeKXz+pGewT7AIRMR786SVB
frDtumNiBVSkMEizP6OVbAGthY9+Wsm7/4RrFlAZppGx86DGMnTjY2xbDgOq4CdZZONVfpVaRNUW
OKFfvYblE/ZJgfX1yBzd8H6AmZlEp5z1g2uMu6nHyId/Vsixjtv1YjHorqs29QiGKFZwnPpCL5E8
vkAyD0F/+8uiaf5H8ilBjq/FGiIkmHidRuQxDmi2HSiuseoUCz1bdTNl3ZN+iH99wr1l7BiT7025
vW9qhR6ERI/f+XDICgWRRYtpjLGcdwqDSh//0ZliCdKNDC7zCN8qTerzUBnv09hvwFnXfEv0YZD2
w9BpP+Ue5WHiJTY6Buazr1Fnn/C3Vpfi4xfGmryfE05VvcknzxeJYDE1szz8SxvQgOf0gfmxciXa
T/B82yo7bs65Ycsd4VxCnOPRYxTuWNyJ8NtsfIPaSIkKtC/BcAEh9fQXzLiehgvNaaBNmb8+/JNw
Tad+0OCgY/TV7Y6y+v7z3619OmSxUIW3a/PkYkAC+XRyBjBVUP3qh1ZWSGXAKHv7NZlrB7yJY7t4
tuEpybzqJejWrxRGSooK6D1bE6TS15W56NsGpr5J3eMV5bzUhhBVdKWqoKMIWRvlQ27tajKeMCMi
tVTHmtQ1NdYoJOZQ4f5iKqj8sfIAt+5gqSHyKQ7PBxTOieB5YsajzJ7rCDCTGORIiG+rV0ipodoD
NC5UYVztQ9mNdGo3UY7zY2x4yjnEmAgejP24FjvLts7p0IF76EEV5koKJXxn//pSDjuojtoY9vFa
JpqCjvMAJRPOwJXaGr9OHfU89wxgA+Hj5c3Wly6gMUt2tKwAtai0YLQ3GG0jTBOYvoPqEZvmbeqS
WCOYvmHWNnWcmbtzKcCPX9eTNOxxKlguNMMbrGRu9y0M6mRqArcW2Gyfqrq+ysgemkp/ntquH+3b
35y+y/IuSED4Nt8t9de3UTVh1xgu6uqrCVoSYC54COcATmUArp2JujjpfrdnZabCnQiMZykM7IRr
j86Vdfh2NrWm6CfsW/78BelOb++cVejeSPpxgs15UMlAz2kjA0PaJjsYYjdTk+eTodeD6Jcsxtqh
siDnTdI4OJ+XGR9kNI6zaB5DQWjG9CjwVFGKSrQN2SQNsr2SQpR0pzxZ0i+0R0dHN/N686oKN5Ox
cv6m5YU5dbd9v3RZ3HfwNUarMppMbSBDx+0gH3VCPnUkqAiJeSJaODOc1VfBVEgFSAD1TV3v6OvP
F9oN7TkF3lidVLXgZ9ASY/PXLe0cpuEgSthkTz1X4M+Mh4S6Es6mv5+o2DcLOM/R5DMiFtVYExjb
swbnSUyE9e/tJX1P/QN7GkjQkndBxikvgV/ud1MeaYEdSE51A3HVU0r7QrkjY6612mVPClRiNOko
/n85b1smmWI2UiHZIBfefxYZkFqcdk0NU8M73XeRr5pfs/bHulcVAY5/6MClHVUc8KGZUcrWYeqQ
uL5dr4os5kRmFOjPgJd8AGXhuNt/L6ngpsUlOX4+rpYVrESHOIn5IHQW4AhTNP767R+VRwv50chC
3qjp4sqDaynijMLKvmiljbmjqb0tmePMwYkcLiC40THQvDMxNY9zunb2LnBeORlVhEU45UA7QF+0
d2m9ov9VcLrKaLArlkyQc363P8Gfo184AE/yKRsrn09EPHJ3GyfDJrG8cCPXjHDPm2CgEPb6TNC9
DM9piZq3gcAwTo2kyZw9qIDjvfczkL6vEPN6nFjWiB2LNStA24HHqcDKi54sluBFyHJ1gAb2FWUA
vjXe8cCLV0isTQBNwg9ZV7A93vLGjxXYaUOXRYsP7MLVK3UbVK1INSY8xQDkxPZZTE3hNhMmwC9d
/ITsrAwIGxFGOPW8YNCaTTAgZVG0JjcqURqjY4rndJ41C1xvC9mHBEAW7iKZH1deOZn1gl9sHKgM
Re+SKAet5p/ZyV2wDkR3sY2npQugabWOdFZnt+6X3u/ZMOKjVXufxXSR0ShKkPsxXz6YY29V/cfq
Jdh1WbElRgqFkCK0I5ZlpUL/wfwdP9DL2KVZZXYEYDovzVkh7ZeLboaKhac56QLENHeXgZ6MLgT+
lnSPNxCNVX5MJPZX2Rt8lbP7X7q3KGJe8R1SkWDp48roGeVPP68bfjw6RZdGtwheYISpmVU2bafB
UiebrWQKbpeYIdO4OoD/XLP7gFHy0A3e8uO0jhTO9wnMZuBes9d0R3DortQBTg/isYp9P3amEsd7
IHahSSDqLx2ApBWRwCzyebjsYnvrUUZVNWNwjNr2xQRI+tEwTY5LeflC6ieSv4FA9ttWvGTYLEQR
39OhrGAJTlMOUyj80M4oBuu8aUEmIqCtvJEqx/H3r2K3Mv6twRuJvs0VYrCPBtleMsvK+cepzWdk
vVYA/Z4H9nxnGHT1psxVlVU/y3AwhIr0XYdpw2uq1UgBQ1xJKv486eMHMHntDRiHlIYq87bVUbnG
II046as2XsBfQPKMrlX/leRP9Is590HXiTKk3hCKKRXwLJn87iHKuSYL/jWVe2rYtUvN0DToUPal
nxfq0qVGBBiGvLOv1Qlwkh0KTsfFQAeXLI0qSsSuMZx3C9iRoysFxRwtPfNEJoRp3jQjcGCpGuyM
3KZc288Pl0P+hMtBNjNBfwCdAiaQLjTHfwfkVpTufSRT6EezyRVQff1wCq5rFwy8OlFGdKXmVdx4
jwLLsXZnXmQk0j/RpI3EvfGMQm77PKeciUGxPSN4J8t1gKpVqGm5tcbx+ZUezfOH9PGWmHZ32zKd
M3Ax0ldqT8tCeBxeFqDpTgSwEt/BHyz5CIouJTUufUlz39OdaDt7aMGv1L7wmmgvD6tuvtTAw+Iy
2SkwOC9D+b+kmHhZcwt8R67/S+YYTD6WYEjE8aEXPxVuN8QSVRvMqR9HsgukTorzt0e4oEVnKjhh
HBoNljy4TOdIn0gdZKN3JKAFokC5PmGwk/t4KZ3lsIHTMyPt1CVrMEua/57FOHDl2Yz5TqP2NZWm
CNO5ROgiiHn31LiUGuZtspcL+3551N5IxhKmSncdTP3//3VtI1KLG2TivLO+AtPRhVHt/JjesPfl
b9Py4PtxY7FZj0wcJIzNR/KDnmac2Nste/pN3IYzVrl7EgOCpYve/CvYlTRupgbDXUHnM0arJRgn
MpwTaw8+0wXsGtTnU8WtgzBzK5VXXCTpazyhuz2hYifzwoFNdthmFmJ4YrCmmr2CwYRlhWixbrZR
Q0kIrELO1VobxAfhQxVNiSzPjc5/K1wYtpLNCpK0nCgrpYsdFgNHm9/F18gtJ85Bk3xF8IZEPRIY
nkPvLx4C6ayyUh4PhjtQYq5ZUSGIfQbuaOITigrl9atBc/FFyZ75XX5DWvkZ49hJKNsVmrcWoq5M
fv8guduesgdVDWHpGjN3v/ImYBVYQQdBZzRns9cATzED/g18fZNCyBt/QvK5Q21EGePAGRie+594
DDKyW5Nqa/dtOgQTsnGwgy/s67i/T2u0qNqM5UmHm9i+ehDNMnHp4lskwnN9ckbOmSs7PudttyPZ
rB8Nuj3bZFTrqVR8lqjdu8wa6IfMdiH9D+JKHchZUhqjJeswPAD3oMSpwJ6jmzYs/Pt8WadHcYgR
12qSZoL0qqdEwwmFYIQ+6V3DuVrTlAE0570Pk7TeLhjJfD/IO9bfWJcTMToMFOUKWssJZPV1VKVy
dcpTO/jdMLlx4Hv5RRp2BE+6WEQwXsC+J4RLCrdK2oIomZslPtQOG+49s0uW9orCUO8cw0KTlPv4
N89qNRdoj1N/7nj2UiK/PYS/HqkifcuHhpA6OWT6omZ9hrSWpOz8boc0KaCtuf/UafDZWfRvKTdw
l7wd1cDwjRei2dY5blasvI585KwhCqbJ0myCAM26FQ0Pz+4Se2hmeVDoEuAbEfn9UTbTMiQmKLGJ
/pVRa/coVi3smpbV45rEeJje41wNqzrk7VDjUg4as90DVN1yfrBycsco+vk4VbfPmTAZQTG/SwJ6
a8TFPGA4n0b2j+kl6atin8o4LoB6ILBtFi0ab9SdCgOiFEkqynTARnD4eViuuxjCtGLtjEJYNfDV
S5D8wB3aF37CHU6dbXHqi+BFJ4kiz/qJ0F80M+bEsSWOVnQbJG+YqxrKLUq+ZO8Rr6cTUMAdAtaC
CJw5cJPRN5b5H7OjXrQjSs3TayRTmAM8X3OISne4fBeLDcXYrES6fWBT3n+3qcAtnXL3w+s4Aotl
IqK9bxjLHFBa74Xv7/LZNEol7VZJ3O7q0agoYkZueRgfYzUXgwVqipqVYkyDrm/Bzz3EyVGHMg15
MkWoivy/3pwHkfx2PZom7O2QLjEfxPwwqHNDRD0lVrOP26svkdoVD4gBXGY9KluCmt+boyg4iAbW
oj7nWqrH2A57yi1qF2PHtNVOPJll0fmQqc27rSYJpnCBUiCzJI/b4xJjEosENPEZTjflq9VQVn48
v8tEQGFl0o6K4uuBa2xtcSF20wDfSFPBoBc0/KSURpUUIxlvf+1qfQAUpdy2jU/m9vPFpa4IADXj
MGLW9oyb+sqw9BEskIQteYz5xI1QZPIm6+0PM+F2H3UDMy2n+xoJLesMhxu09G7SKrbbEqq/P5Gk
xSoqEZ00nJ24YfOo/PZ9aZAnIBjSRoUlC4jmpfcSNnCtYB2HVCPkcX226lt27MgVOZUxbr6Aybn0
tLqJtLxicCDndNF62WTAf9OSbcQAZoDE5dCBbMzGUR7PpwzT/gaM5twGvcFF2aZhB3c++LBCQBT0
zIHppGsyJFgFz+dwL3BQNI6bZ2g74/qqoRb5Q6X3Ts6tXYBXWVxTnyKCCz/H2ZFnhUCWSMu/Zvgp
OOM8J9kIwIJjwpuE8OsCoyrVD68B+EY/z4I1ecbkQ5RUPsP4qryTf45Jd1Haxs/9MkrjcftqVNU6
krsMhQpzeL20lyf/P9zzM0/FjBuYrICyHCHXLjZQtZPR0uhBcC0GOJ27pyZJHuJCunyNPYG2DydT
V8/SKdqiP+Wp1ctm7ak4n544Tqjj5aQmPbo/SB8MHb7Q02dsr0zVOyzu/We59rxMupkEskm5Cpxs
BVeuXtwfdK6xV/7zavdsRRRzMoIBo9LDQE46seI5ryL2Et3HEJuBp1je5pASg39PhKLbWGxgQ3qz
Q0HpNBkrMMlKSLyfbHHo9dSGdMKkj62WaC7qe934WCZGJaEL+dlKrw4E9XgBwK7l+ruGt/Fxf6bC
BTUeXsuVj4UBBopaO8LVztix5j9kUBwvCbIhqKO29XpG7dvH/9DC3yuV/CYnZ3M2nDbLYGPC9GK1
im5uAklYbNKJK0UtbSf28aYMM+lmczUchiQ8PuMLPSwqGz0fhlgovtXjDyBCl4lFQy0RWxIpZtEx
MQSuRq14CCpPyhcGYdzvTWDhEALyUiTcWnjnsrqvrAT59QnOsHnp8/5OmLc25l0ArvEuhVVqcB+S
cH7tVLmpc6wXkSRzi74b89QyOgF+Ry2KLeBUySOpbkvzjlmUK5ZFQ6BxYYFiKz6JHaFcPbDT9uc4
++t6xnM6lDcYUgkvj4r809PYbX9H3KdktyXVb36L7zIbmnqiCXys7aTOR/uIl/AtisKOzfZ1avVY
Ao74pKvN5yKRSvIq/nkcavtXBt1V4xO9v1LW17Ybl75Pd8oZDsVuV6ju0xop4GEZjMFB3X74ROxc
KLfnGnuVp0xcOWHbiu8wB9iwGYdWI5zkkyLJP+7uGYh9XjknM0n2XdT7dz4bLPT+iq9LULLcpIk/
7g+cIKzpsr1aHcfTgaQPgj4fYAn2TDbIVax8hATAze5VWL4cdyAxLKSpxbwTjCJfoF31exJRpDKf
GxPGF/vtR4fIIdFLGpaIwWduysPbUWB4FVD6myCwK92fxHzl39eiDG1rUsxJMiwLSzHTXhj3hkhs
AH1U0MHsQPtTBoNs31AbgSnqwaNa7Nh6Nr7zGkh/0Z9nc74j5eAklcVgF/jwwcVJsKonjysCGG/X
vez1rjOFGagjZV2BdStBWfteJiKVm0U3ZiUPZqYlIjl6wH5SuL/aGJUoHrpStYZO+R+XKDJdjEfg
F5W3oPEVuAACaGctAYK4uI/TbMgdN9Nl7jJD/ZZpob2ToqHfrotbTeKH1fb1eh4xjeUNLC9u5+pa
EerzrMjIQtilZacf44HgDVpcGYJrYAeeJ6BGbbf9xi2Smtk/pSHh2TtZFL7mS6ofgK2lGGFzmh3M
XW7Qdfo3MBDLNt+mXLE2UZgOh0POH1TuE0mh0SYAQH/Cw0j7S5zPbzA6mQmp1DPsg1ZCo27gukcV
oQC8GGHQvQh36KAVgkizJ1O3xiO5qAcOOPaPA66B0krgHUDWyrMgg0N0fJXDXmO3ie2jKcMlAQsp
wms4nMbMcz0CVsj8SGP36wNhQm+NweAMTg+L+UAwAKXH+w203Ruqufby0rE+niSwVhbVFNgwVm1Z
VT15WGfjT/SAvcRyPqapshHlU/vGHp42lgrPLE9uGIqlGuaKwwTOZNTU5c/FD1uiUBNU2+Q1Jpii
LRZc0j42BJGVQdgHK/L/WxZXyCcSsK7r3OesUPZz/jH0fajHU0ebN74pqFw5prMXc6CZCd2j6913
R0g6IADL3gfky33/IGl8hE8DI9+VCrvkhSBHaZkgVDHMS3njLqwImNSP4yDaBNAurOjjSR4RcY6/
gZjm5csi1DDblNofm9a/Ydc8Ff/Nz1cia9w9vpsx5qA3E89dmBJipdeVATGLZWF7xVMpmwhEHKXZ
rKEs4dtPI/66fRzJGf1tO/qWa/VQwQ7JIqyzFGWGvOa5KvnOQQWhhdUeLX8P3jIG5aKlBh1ACW0I
TGDhXOEGc8QLSl4zWZ2XpGM2WRKUcbu71DzyKgBfBRXYIP25/J+8uE14Fd1vWMjjXjZquyB9FEen
B9MZAlhpbxiUA0PLAl6oG1AgP3EQVVAg6NBd8bxV3wRLlf7KG3fTyHBW4KQt4ZYNopT07LEyHLwp
0xmdQS05+YbgXoKNAUhs6wiJZ/pADNK29SF0l+qBjr+x6F0bfbJ3hMSJoGSVgqC8SyjRr3zJvP7h
eL7XontHM04cahfY0rLlJs2Gqe7p87qxeHWee9l4uOdiCU1XlgixQugKofK9ta0i5A7IrSNV5Rkr
A6F1vzjqqfT2TiPBwwyZQdzqgWL/b0dDib5fDbZhEKkOxr1mn7gMUxD4nBr+ei8SJtZOhokJYqpP
w4CEfdJZ9sADdB4VWb+D6YczYIsqHJ+DuMtly6O5Nn/3HJK8nHV/O8s4aDWEMvPAssgIsSp7wtZz
kcP8iPSWGRLNpocPLRRUtkunP2GCC9+4xRt9N4IL2CFXs4bgCctW1UDCiUI7doRVFsA3/yhiVqH6
7WBM7MBVBGoIcWiOi7NicTVWwdu9sg8hvrA4+plUTrtPNEtze2Zmv2LaTxvFMrSmnFDWScQnTuL/
zw1epLgf3IrQglOt42GlTFBkU4eGPee+cpyTTVTDBNkmLtGQCGKah/Uq9DQ0gpX93MN0gfW4UFc8
mrOBEVG4vOZc1loY9uyw/iVYqW1o7iTX18P0LtNQevrB7Sn0cWZeN6Lkwlpa1iJ0UfsODtCTJA1x
c1odZVcwK9ZgQB5wL9utTupkMQbSVn/x4YaAsC5XZmXUIuDcb5h7TNTKwTE49KrS4XmbpJ42dB4w
sc9gn7kA6uBbwT19op6SONcGixQSTe5C1NyNDmYbJpMH8MXKf1Jc8vEVDANLl0776zVr/BuGTe1P
yEYZVsAHywy2muIHyRFQW30NW7riPwVTU+9+yGdvdBFvBqjEp2KnGMzFLchnRJ8kI3KAAdNP73J2
el4VzS0cxGhu0vZPgO9JM0URXyjTgG8hST5f1spYjO5CzO2Av0vea/dMgk8Dq0qZg24IdWbT23Yx
ryaMc1oFbnsMT1Ir5vwLi5bsn/Lx2UBG8IbJ0LjJeET1Q+9s4Xj9guWx1Nnx6yR5S6ReE965KnMK
aYUREsDWIKT/FeGlXkgM7BeE+w6fgiUtmkK7XQ4ri2IcevfcgcBMAPv2n7MSyfHU9O8Yoy+49PN5
R5zetNdEwnC721pgb6XBwORBSOTcXJDel7qnyl2hDoW6U/moyixwCLioj6Wakm6Q7srQlaHNJ8pl
4uPHm3hJ6xZwBms7ldI0YY+eRlzDaCJzICl9964mD+NEwL14tkQwZNxbDtQKYzUQHZKFf7Axab8L
zvC+G3wmzY3bQ5Aq7s7q9mdu/8lzOLdyhcbRym8/YJaHlcZcBw4UsvoN/3ZcbrS7VZnAg74eZspq
wWBLIIn5mHqLDO4d+Zg/KmMtlh03phvb2oqK5gHO7fkqsMOeTXv7Q+HlGIqJObL0HMObHWxc8NcZ
7GYFVbNZi7dmy1AAXxYqq/nqQkTso6cNAMNx6X/cq5/9jgXvRI5ZULVjjs3QEm2OpX88ujeU9Bzu
1dBH6sjhfIku3xtdfAkdFXlNI62tfqbEBJoBHd8S6hxv5YSVzLSby3fCusSPDmKirXM1iTVE/z2G
l6zaqraMWc44O3p0Bt6o/P//bT3GJ8V4J5LrOm7/vgZvSfdNVWFn2QR8wyvoW18dQ2xP3c7gkjjk
wL/eNAxRBpCDqa6ONhgo+yXiUbopFHidRg1WMYjl5m1eHDJGOuaOKGUPPL4wSwkIrK2odTLEt8X0
cFgYmHbwVX2aBb196Rzvv5iJdBGymyzYyfhCOFzZPbxx1vq108Lbqag5MbdrIshw8o6kntX24HPg
3AWDupHAMgyvXzsWubJA035buYcG6ViJe0hUlFDg9tRviiQ/+hpVoudYZ1OV9mky1P9pNZDflej3
6KeCo9t1XEFDJ2OEPqItg7ZyRDBgQakppDaqH++WPW5awVHCe2e7GHtok7SrhIM5E6ZqmMFQ8VWX
YvNW/nRvugawx+QdcP8R+YGCa9Q0OWUZ/cvKQ92UB2XlaMv8Kl/vvUrebvZMl21RDxDJ8if9tY60
tIsY2PnmGI5Y5t3qSE2dNc0LpQvX69L5SSoDR15w6D1NkAFI46n02GIPHXt+W6PHafjU5sF4MT7r
WcDtSw98J7X7ngcZoxkv4zd/1ZngT7hKN/SkGEwAkEtsDrS1agIz/b8qwr7u6x1G4k6/I1DTO1JM
698OHJA8jsy2idVqr9J/0+DkQmSP1MqbjFjFZBc30SAefv0CAQI8utzvNZL3GH5ACDJ8vYluooGP
40cOIx+IgUyuYlekjoJnaV+bMEzVLDyfUzLgESXkdm38JJXA/YHyNRn5RGDI5E/86+EIUxAUWlsg
MEm6HCJU6XLf0bDaEYNjSM3acs0iEK6BLxClrcDHSckDLC0Z6YqPgx5Hv9Rukdvr23dB990Vj5Ec
tmkXadi+atgtN/zgssUE2XJMjM48RFfCrc7Pjda+nmNRWaDzAyNd/xNABVjDoJu+tXUWxxx//JmZ
cWE9RbQkUN+7DFxSGLVEaTxZNw+l+9ek31PouS+Yj2wUQ0HjPqt7VFOVfinyefqPmkP18Dq01ALK
lfaeT0GFk3MPW1HjiWuq3+z3HMGWinQkyBtQDcN35ZCqNZzyjf6jw/2VXRZWVnm23jk3D29nfrjB
cqxInSYJqL1VIV2Tu9lWehnPGuFy/m8PGN/Nug/rrzW95QbJklYigvb3RABqATHnmLJUiyY8fIrv
fAbEZg6S39yR4jBO2GoGjvlXvNyqvgfzzySS3pvt4diuML3p1XVxQH/QVwgZNFZ9OKc4lUgD4HQ4
8qjm3zUdHn6CQjl6ikWbrIr/dklnBMiuJAkNXmrz1cKlZRKNzH9vCAU1HXSo/giKE1zRgAhgER/Y
Mq/oV1ATvaDIybK7iGOEABSQicbCWRg+QsI+EWbKQkdPYot0NchNUsRrnP7wBh9yyVqUJi5OjtsO
oLujjOi+8FfKfSvwieucvBhsEGqxJsUfuVQsaW2ImsRFKrI/gGqDILZtaaOWoBLo6Rh5P/mf1kK5
v9U9GSgwWc1JrQXI5/wFHozYpBajFtGCFTEYTndK3WSnkottkzy/+P0lOgjvad7RN5jbfdO3NG5b
N/3BxLXULrI7mzlwZnc8mUCp+k/PV0kh2uNIeo901Xw/uc8Wzp5XE94W3udX5gX/GPJEGe9eg0Q7
4NOjdmkI6mJ66nPMdSpz05unJTJcj7W6vIARLx7dDo+TRmrNKk4CRJUU9ogPPRPkrzP/tiEC85zb
tVFvc7FSV1JL58MwdBPLUhcWFHTh8fbv9yRy9/iGc4vgruaoBwLDt1e7yZkE1jUTfmcDStEJUjaH
bP4V3oEe6UDLl+tR+LA3RLIf1zajIwxmHVFdrIPpDe9SrsbXUy+h4WhsW0d3YVdZgT58BmbB8CXw
OsGxfmS/ITseHfsAAaNnu0PI94O7y3Gdi+z+rhsFGREbPIdC515QLiLTr4Ubp6baxhR+WdCLP+30
7JFGhw7dH8j0FMHuKpufhO0tLhWblZBCqe8Dr7IUBXg+9YXClR5ICNbDvFPy8F0h8mYzW8/GbPbC
Y1+lYXs6RdM/RvGpznrEPeweFB4KhrTk+5yIN8UF6rFMf8nGbYxZ86r57qbuc4OwOmRduIfuDY29
B1YObW52UnfVC9hsG2JJPDTC7t2L8zR9uHr2umxEay1YUil0rwFCdVTrkzBayPnMXNNGMRMuxcUr
sFnSq9OiBeQBSOO+Mtsb3Yn+AvCojCraP5M45qBmOC9Z0Dmy2zL6Hyelelp/26/SWRjDEy5FCykn
LBfA8u+8N0YSsnVc06zT7sSbVi7MejRHpoiiNf7fj4MT3CKyx5PjLkWSmlNA8fb1qyDr5yFBGfUm
FKYEyrt3uh7Ee1YbL3FFRwszA4yx2goBzwLofspuiXTH1BalfoLki8jRmVvQImlPPKgY9bzh8LoG
6B8jbNX2HdcXdzSlPfdbLqnr0ZmmzzAuxNRQq9d0ReM769IbPPfrvc29Y8EkXPEpSiHfpjneP7uG
oQ9KABZXSIpXNJRhFXkKKSQ6aRuQNIKLQMibOQrYlfu3QOvOgzDkYSzGdhyKJM2rc6G8jeTL/sO9
KEUjYSYN+XxE6iuZA39r70ASv3qOFL0kKAwnIEfT4vwN7VDcB4GTjkN/KubqkNOCVf/+9A4JAsNB
HlgvJvjUCOsK81Up45b0sKNfowm/iuQoLlCCCPoN+T1tx9WQgQXmjfBm6koO66VKGNPaUKF2sRwa
YSNyrXZsL/cIXvsB0EIs1dYZRTf+lPkBukoN3PEjrgoQ4nw+UJrd6SCuH7sv9p8NYsPf1WHjSVdn
n3WqTFNCoX793xeoD0saGMQDnt4DTRY8YwcXeisFoES0Oo9R+B9KjgytRgbe8omXuB7FqNU1RBJ6
cm2/uJBzs0dRyG6eVa65oC8EiEz2JDWc/a/Lon07TffPPlM49QJzX6wbOcD/A0kgFW8JLttY7NYf
sfG/NlPEhDR0k55TZwxbCl8C43BnLOs1XdMd7Go55I2/O2XeNf/xzJM0cv1QBd8CuMxdN+2/ay1Z
5iI4iUngtX1kR7wIeU0Ol1ol6n5Ma81EDUUiCv5TcvLluEbyXszAB427sMm6QMAkepxJowwgEt03
EBZpJBJlXWrrljwFz2yZQmIcrRJgcIKtit+QpTpbpFR3xKcqUXHE2SoA1L+JfMi7rpyjyhrA4Lzm
NTvWw+8ffO5qsbHoq0GRZ+lKhu/6yin7jgNDBxaW/NHv/f3nNKNIKuCCYhOmvwWgg+P/HQMjOlDu
jjIYzzCSom4pLyNdKvKUUAdsA6mYQWh2CXk6EfgGBB2RPh41mjdvn5B+2/5W7moqypxIikvGf7dm
5FMxiw8DhRIV07R+8UudMIqZORur1l5vwoMP1/7jkKPkoh8qBJsORoMvdOXkdZsVSLB5ybVZAgka
LTXu/BUXg6wA6392mbGCPxU+DNy/Mj700PnXmtutrnnNu4r8DnHPe0zvdD91iV4ATe+5cZtpLWvQ
hfb2e/S568aT9+1DivFYAC6eM6w9KB64X2dbTn9hvAw8WPTQvRuNYoqNNmS2/RiYF1QsAlwjqFO4
aQ5Pjcbk99DM8+Tc1qtwC6SUqiX+TNR/3zzf7QN9FJJuoyqHn838a9tn2bW1ELUX8Sn46btAzidz
xEbP466Gh8FBkuZBMvPrNfr8EDk/gKGT6FRtNaV6npQhaHXvfyHGLLoe/cnmbV0uhDgLAE+ZUpC3
Lg7RECcqwRBmGdk/lROtOdOD3/1BS/y4sBcKCVNQ0IYew0l+lQx60I8D04J/kvf/xSZHCibr8GOi
F62eRnJ5xclf/IONAFJr2jNyGjRnDlc6f8Kpe1JjETjRXTVegqDezLuJY6g/ltWlO68M2WpeFkoe
DUvns5vwFExf199x7u3pRtypbUa0vrBRHDvCVFw9mQ9HA8C8NcA4v7bjp/AUNCsphURm7E/f1tQP
bR3FU6pgQ3uc5WaZMohLZlSqID/sf2CIvSwCRKnwRo4jBO2vbplQQ5fUvumma0nziSxHx2bwfxfD
Re6l5PdEMuLqPcREYCveYCPVi00yK1lwn7VV4UXeshrq/kHvZLDHa6xa97oSRKpWLr7jl9cHaLlf
T5VM9rzu9ktJNL8bG8WjkIVSojan/QW4xUb5PSngVm1iy8T5FnOp+aofsWm6yBW1IFvY18ND3Oox
9ZrB1cLvdKfy+U1D1CLTae8TKuJMM9Afh+YEJc+bm+ru6hWYEs4TXzWSHbxnXLDO+k2Ey4Tt2gy+
E9seEtvIhaaxWDHJt/Ey8v57Wl+4wGn3roRJciW8hGsO5ak4zf4IeY3YeUSFSe7vQAQK89vcDGMj
ICC9Yd2ox66o/bDhuxaWc/koSflcVjPhDYQ3yFKfbmrh9XY7HGYNOqlDzZKjE8/k08wjviTMj7cv
Y1t21dfUcmou/hbgGT1/qmWF3iqQZ1gIGwcm+I7uXtq91+XUdUMYLuRZZIaxKJjvA3twyt4eRkQo
Egaj2BUzWoTqvtOxNq/5DchON7wKvxI+CbP0BVI3fmZkJamHtE05YMCP1eLsWXotSdklr6hL6prM
ujWwwypthxgPTpWgHm/X0We6pmbJ0DptSVgJjK4njl1RN4wkoAS9yfco2P0UpqwUDioT3xi5wqi9
GOYFZ4sjlQ1O9aGZGumXvzJ7WqaYeCQkeixjWNAVPFoqJz0diXury42oGUxU8W+CsNrDiVuMNTuW
Sa+eM6hRQmmxuD6DnhxayM3c62KWhWo8udk6p4ODpX4/hmyPnm9R2sXjEHwaIX7xBQ5ANcLsrZGh
P55cO1Sw1CsTXEJjhxUz3KSl1//MxewKMbat6LnWRbxK01YM+XUzXrLq8pfdVgj2NbRFwYdNEZ7+
3K3tsaQgSz/umkIbQOOTVhnlrcExhRZ2gOopzWqatp5yEJc698czTZFxaaxXbmTrvUhNLyMTsSE0
XIqGsm+uTWGJnHpJxvb8Rdzoqk1Si0TzgFjAdNFK+YiNp/TqHEO5V/B7/tSD7XPSuIfTN6BtK83F
QEnz7mXESF6GO6tKtM20JbMV505wQUM0atn+3AlMmzkHcMTe3Px/lbma8cA3Ux7sWzce2qIKvnMm
1/LskIcBTb73YKSeRa85qIRpVoPVvvyKC25EMVWmm1mDjD5k1UBPOpAoLzvRsr0xZ1c0LsNFz1mY
AChnvHvmnQNg/JfozriugB43vxLycts84dd+ZJvsc+EQSkIhrPip0FscPJvpvVqnR6d0vRqjh30B
SxKKqBd/bOtwBowYkW4uRUesu9OW4Q7oRJip4KQAfa6UTC3B0bGsa4F1ghuHTfDyOTcAYy3i+tn5
3r9VTlpXOkEm2w4VvTjTQtCB0MtUV2rOJrU58nQkRMIQeVTKEx+Wh+N3HbK8odCEP3CwJGhREeKg
42I8CQFreNOUD4mCwF1rpdvkLZFttFNq4k2BgLsZgpIbnt+hHv/8FrjvXZjpXgOfaNRbgg23qpGe
XsKE4uw4RlUrUxym0+iST5nZEREubhVi65Y++UZbS8+NUis7GfUdResAQ+AnSaRu1nl6gu3YR1Cp
jkExtBwJWThwQhueu6nHqwMxRMnFviD/R+z+bttAgrAVoApU0/ILP9lNkCq8X40iE9OPKdM5EX76
9etT1KMHk5myY+n1Cs69OViwInmo1WREsM0pVh7HTnqSJPp5Yil3hNkgpX4gmGqVmgaEUAcpnd7R
h2ulKJbVTtXcw+unRTsVj0HdJryQcorsRj2zLh/R3IlIZ7rD+3WsDsjpyoKzu49jIW8CBuHplOYC
hGxcQjfwuF+JwFh+M+aRuNXmr9wc8W3M0R+UsuGUt6Hl2ZhssSzLHStliFSQCijas0mP2T8NO+fS
p5apwWQGe5VxJKEhML4evdvzIJP/x5ExJ8qyNp+krR0KALv1ZtL/d2V/HnOfDbVSGUQeP5OmHFk0
xFUgRS5HU9pA/QhPGnClyw8RzNKjRhDgnKvmFuSWa+u9vF9BRapjX8bO9FmZRyULz9a/x1dUJr3/
vezBMKxan7VtC0USpX3D+8uM6yWuE3B6WiNw2BNteKc56Lb4w7cctUzcUfVwAMGPQgAhFdlPkDk4
WrzBgLldTE02RLDz1Qpt8iJMEwY1zw8xvdkXeBwiyE7yqmtksIbZt854eW/EKSYtFsEgu+wJo3yS
otMnI5Z0PUeGJk2KUI813Sx14vroCdDUikcNU1pfCLtmWSfImpTsaiFCrOFlcnHR6Oet6zrWGaBy
FIHYhhw96xn58YiEFSHT1l4yz8sfGBCVGJ8uChBidoUwOgOHTqHRvcc0RRmRIPr4PmMLiyii5R/U
MKYTMQBhQjrHLcjPa9o1RAePlbIU+cMn5axpVaDD0OWBDb05qGm0TicaHm3dbcG5CBJ/0voqwsbi
zeFSaFvov95PJf9lgGkodjr1xOCXL9C1Qd2791V5RdFRJC7/zkgi3vXmrTGndl0zq702av8+HL9o
KqppZlfxrKISz+0eW6rJlQtI3UOATXuHXWa8grcNzSN4FE5fdcoWDuW+2FSDyVQXq6U8iym8ZdTa
g6bpUOsMhr0G4ElY3HcNExw/0+GEuwpkjsx/HCX2CDClV5e/wQzIL4sNy00DZ0wVasTrIiPFb30l
48CzwRwHdq63mlCreYrVuWEg3PxmGq2Gy5XrtK7WEYedyJZOy7TFPqjtao75Pn3BrlKV6reHCd0E
+Vv8kzSh4eQC3SS631ydp0L15FySiZoA4R8b1Kpiqqp+vJYK4ZRA2pDkDMabCXjnjdUImK+ODvoQ
90oi4Jvi5pBBwykK3oZKsCPogiUcZyV9kHepaOhFAmzpZBf3ipV7kdDJsIEyr1dOsWwZSi9H//Pn
jzlEtEMKEMrU3DHPnNHm0RFf0FkgEFV/sehqSjyyaTTQKp4eX746hxKt1kI3fS5BWFhIFIDUYfEk
Z4L8JeBMLSjvXXztfaNc87B+qZnBb/hCua3i78CYBLJrcOS9MqQCsIODKgYrtgF8sXLLLB3CaB7j
orfppWcgIHmXXOyZ3EK6gGTfZCNG4Vd+JA51Bez1UrL/g9UZthNsQ3q5/RH2nHfs636liLLeHzuR
p7fjyjJcDP6rrsqkHCJT/vyPRA7AudhGWMNUOEtSW8bSES6jntICsXGbbvI5JGnmAlHLGHVngTam
xhJ3nCq0DU5BMgTmc+2Z86+bOi71VILAkGA4zzkF/cDFpgBShmdNvTepkMpc3YMsyF9tAUbWoXff
Zmdn9pfdREee1CnN7CQS6J8MimMSm+SDqjXVWEDIGH6Gv/PehlYmpTW8xVJ6Td/MB0/PSV4cyG2N
vGwUVXUgHSPwehEIPCQzaMQsPIkToRr3JI2qNiAB3XhPtMWocOBKI7360XZ9GCmtr+LwoZRLFxIr
nk9Q/MVyuGmhub25DRGUeewpRtYAzrQ+fVOFieCPg4x7uBHAiMDonLhA6/gp8zgwvekvOqw8DqWG
VB9NUsJQ+FZ85kZxxwSKUvHZ5khaQcsTb1CYurWoYsxNVe5oiK/aDf4KkirwsG6K4Vin/oeOEVOn
W1glqlao/Ol7NBVTvob8aE27/09LovmMN5chjk9e9yIHvYQjgboLXyEo8A7ZswtB9Wywx9JaxtSX
0d3Jn4AXrVcwNuuSc/Y43Wt6Dt8mZIBzot3DkzKucvGtHjX/wnnUQn1pWGIBmL2+KoGWTwL3ihlt
y+HWJOxdlYvJUfJ/gevF1XmdQLQGILJ54wgCrsM/+Wowi/L6INbgP7NJDpzwXWkHjfdrSpyd9lUB
qDFylWroyfFizbPJoma+N8vuMCX6XA+opbZWjSAz/80XnlzGFz/Tl2/5ROv5tiRvr5L+cQOAyaYo
JDO9WJJ0B+z7niTQ0e3nJ5HBJfNMVEfIbyel982EDQGhAsAv1lfmcE25Kel450z1saqKTPJpZ4nI
nI0J1RD0ubCPE+acanI89mdlc7PPN1z3t5iGzmUwKWizWCxTY7bI3gsJK/Hj5OrgirExw8uB2E3K
+RqKtaGCLHRWkbSjGu3QyazTzSfD95SSEgAeruQTRngF0e/SNvtR4031f4Wfg2U5Wdz8juHnkrrl
Ij1PiW2fLpLgivo9edRgEI/Mq5e+Lw4LUYPVuk+v/TcRJFxc7t+DR4edkUvtMcU2I1zQXPKpEHcA
QATCdunmLLy3F/0nYVpMzCLkyTqKcb6/1CzSim8izsVUrRoZyFZm8GyCjojMxejCi3XVDv0pNXNa
SYMLvMP1rN/vNfadu0McPPSsnDF3mcO/gpJmPmfZ+M/eCu0DRNAmaoIG+LuiJgmb5+6KUH/NzUI1
9/deUHAWO+dLgbZdCsuk0w2AMQZmiudPNhca+V8lDNGMXqloHd898askJldi3Id6AgtEFBi1Qh74
bF4xJm305juaJe/jjczGPWgX8M87fEpEUI0dUGuC15oDQCqwi3xTopwW05Vaxh3Q/Krd9FV3wP8M
hsC8NDAWzxB32E0uaJ4AqNfgcqo996ZMWexpMOci5lLyIM3YVYP8RESraMXs9zi4RABdMCLEc9Is
HA54dtTuMYdj+HHte4N+EczKV6hS0dDNhPo6qNvkWcTM+EcvZlQQrhJdGKM9EO3lwQju+ILYNxrW
NofyOjJCs9cwYFjFwaLQ+8AdC7LeDGi5xqFE6yad4+IFmbK/UQFIqU5Z/i0hRAZcfmT1v8M9A+8N
7gGVg3W/3gCb3+fedH/9j8BM3PNxa09ajKLQjhwA6c3dJ+DBwacuFGFHX8UTGJbBbhLuN+dl7fGy
+aH3cJWXxKS30NZPKf0UC0SrWvTF1zZa1rRt1uOm0AldXrtrIW9MvuSbKQeyOJaYDnoBIlBvyN91
KhIwawskXFx30Vg+WwabknoISD8ea5opDAdPoUSIPlD8M8envFa7vvtAG6gLclvUcYwfvXgVfsLL
kOt2ebL7ChP5QDbH3XR0a3CjmcpUlqLrRl4bcINermEg1L2p62p55TxMyz4ENvG4MtFCCI3jrpOd
/w0/TL0IyPp+Kvy6LTfr7YmWf83gKQz5wXxz2M2+ydk0/fexNVwUc9hAPNeSWpyByBc9ySwwEB2h
tETILu0IVWvcKykQ19v7QGsDFyvAGAgwtu0GMNutjBz6JnWZtW5jYIqpt8XZ5EsEtOrs+f/IgBhQ
/aNM2WXQCgZix3ukdY3sZbsKLV3UwVGlt4iz3DvLvHdEv+5mDijmcEu4gYgHiHLOVRBnwBF91BJg
jtungDpyb27kDoaU0tmdfFManFI9l38VNOFusBTf64gy5wFDok01HpEklNFrn0NfRhSXAuW1XZNI
lcOvTN0wQ2QZibubWP6o6oPoqs2AJgawdiqRIB7YjVM9UGwlVEduPikQWSol5zvW+Y9m+TBsEweD
qkICcNMbsiEEs2Zl2LDhtWswi23muDfWcQ7AhQKVsffgO2hN5+aeV8nO8mA9FDc+1Q1/AU/IHhr5
w9Xo4xTgHk9nfVBxjSjKgiAChS3ehK63ExQ8o3FbBCCjzeaFx/AaTuC30b2fH64ZlfQMPxPRjln9
JKC7nkaOEfCEljaFsAqFAXdQJMvWpW0hnWpURcxWFjfYcRI/iaLerzGgz2jz0OZaTI8h/R5/G0Zk
gPa/wclfvkN867vXZKXhIEIwMXOAxAz1uh2NZC7H8wEqAxf3y9CfP8pi35wUSGXUPJCNBnJ138QY
3SD2/79IHeRRgy4DjszwxKhn0mJ6IDJj+fX6+QI5aELSncwUWYXtmsSjc1dYwNsIQiEoR7LBps76
hGNVAoIEsPS6r3tZmWcgWyCprVs3UyVZG6LN7BVCoT4++X4tmF2kSgsvvMvdqxVYGmZAZnH0hPtx
P3v/PrXgk1wx2DI8DcqOMXu3ETewhWmnLs2ABoiSkaa7HAN4lJTyz9oDu+gG3mHiCL6ShY7RWgxL
tDrWZIG49aK7lMsOG7M3AMz/fwuo0K3Aep/CAdwG9K8YllYTo2EHdMWmXwfSGMvCynq2m6RZ8SKa
MiIJnY75U7xqoQmCMSUTnZyKOIio0/nCEKIvLXFPawklO9KCwbN8GnaEUnbIek526jVYOYLTRSnI
Ql5cMvnvwojmpC2jlF6Aj1LhCq5v3Xadug88NKT4RZCiI2r9m80tWJIPGqIyO+USOYnFf7YC8JAd
jv++r86Z4x46iSQAFJmHRR2LG95Y7omoWbnSDAx8ybEIY6n2euMhdgU0Gjbdb/tzrKbC1eBSOq9b
+RuxNYa+3jEfUuRLYz3FNA/LiA4v0Rm1MsEyhSIs1CBtXeyqYrl+CA+2AOp7MrnSdv4xzQgiK0tM
V9vhpvXSHwuOI0NcUcJICOg2YiiPMelolkSoWnZqFifvXZuRgkgd/gKMOpJlyuzPh4n4jcbFj+xd
vPMsjabplkg7KJM43XE6EvrxA+FMQsPvhTbptnsh7/AnT1bkVkKD5UHA8GcVflyOXHdS5MI9VajI
Z1ETAIxQJA+QoxI0qF/eHVn0JKniv3VFTGbBoOZ288nXbf+3mzk8OJIdIh7VzZ/j9j8pyHMuRs7P
j8PbA1Ymijix5e8oiZOqTXUnOMQpnyT1P6s2ekDpDVWAtwmt8473/4JrFxiU44XaO+Mm6pr0hktK
04OuG6TuI9OJcc0z6y4IDdsp0F1DqqAH/P/KifhJ3NJXWN6xhovpS1wqn36ePDPwm4nWHm3SGmqH
7rKVg6UeFiKbKv490AAwM2mc2zeO6v9PyCjaMVsO6UzBiQvwz4vYdg0upE/5fUU/J31LKEMfECvJ
srv1ge1FOmETuPiUN4J5ASC/4aqk0tBP+p+EDkbWMrJdUjH0cLaPJQfdskgKlp4HNJ4EdNqv9Da7
xhtkCYGIH4fdEmagUiQd+iIr6kMvMz2cgHc8aEzwnmQpfd+tuQ0cGzgb/PHoFehTOqUVIG84gKbU
CPhZwQlBWegszBnscWkl6zjzQcTX/4Li9iO8r2w5D2pu+kzSzec8jutMgwZI+tOjrgA3NLaVJpIp
ZJ5dpLw/rR8Mw0NRwy2HLL5FV56UycdEBuPJmyZ4mYt8AO1sJrXBMx35oloI1Ls4giDJFfBWX9On
yLZpZsY+uukAPlHzwlPsCTuEP9WTX6tcvpJc3lG3DmW91g/8P2C1FFpaPUUUU3q5HCsRAR8M4QVH
ckxqUAOH/jWSWZZo1uNwFIOChq4qSwrwdx+Mf9Z0odJANFD17KG/Pz6bP//kmhySkyAd9CD8jexn
KINn9ll3RUGQw/BuTGCidQIcx2pFrSr6YP8M1Nnrxuf91LT7h2/B/UWbWfjzSYqGzp8QeJrh5jq3
FKgZIfKrbFWMOUXJiZlcqxskimqpMrl5Iw8MYf0IXBq2MQDXU0EaIrWVHxoQTC+smfFbRctQL5Uv
wW2Y/uT5ioSt5iPA0rxkOfJ9P9i+JAzElDaMhZqxZEjgF43T927JcRUA+P80vYTRUs4idwvrygJ6
B7ueDNo/foClRITEq47OgtiFki4Ips8qoWeiMmeDHtR2M0MyFXyY2pbw40l0l33B96q44CeVP35I
5SutVxRiOhP9UuLUiNWNQ4YDQrhLNW1CvYWHAcsrLOeHmojtR/ZCnxHjMpDmC/3tHBEisDVwlkSb
QwCQIwucWqW9fntKwGjn50807vfOhrPNOxNwPOD1fxVmxN3Vu+huXTlf3K3rXfkKBw2S4pEJX6W8
Ut7Juhl8AWzs6EMVMJPkmx2steVrwKgGtlM3EKBAFEyY8KxwIM9NICEMEk47Z/m/rIgixk4TcA0I
7XyGRm0mGeeiXGkjD/Ex8eoh1+L4yn/oHYx2+SYW3RRK63xjvPI8eHs7494aOYS+0AjyhADN89Pn
hz+3Cu2vW1rqVHEQ/b4IoSoM8c191+POrQGbhLxNIRUErkUr7zN1rZdCLSBn7JsQFFRjn8YkdtEy
8JGUxUb66yhj6c6kPB+0f8gu+LCFcz8KBSZu28dCfclqh+tV0ZSJefT/q7ier8/DQ+Gf3od7WJ1B
6s0A4IqUsPC48qUzWiB/6thkiMjeS3gK4laA0GuEpWbS8vD9p7fI2jQ3VZw5c/EiusNc+5YFk7I+
xH76RJciPTBvUowsiXcChovSer6MfE0OWd2/HH5u3CD/Wl5EdxbovEVX+Gj3hSCNzOgbavC00uHV
J6ZHekcSmZ1WA4Nqq6DWvSjwjFNRJwJ2tv72AWjdjQQm+vgZlasHEMCTHyubuS9ktAGsYQ1iQj4K
CvUZpRsXn9zQ3Bw6R/apR8IIx7H0tr9EFTEqyMIQwGP0/lwz7x5nqeCIUNseAxDF11FxfBF5EEk8
KIzEq+SsSshy20Px+XE9MIBMxiQ6OCOtvNakPsLrFyegN1qkPFMfwf55IhdlA2veWXwIabdFq6SN
0u9iSvRDhNsR3XQ7IPt1S8Jsxjm3giulx0V+hI7iYzO1ux3+ayJdM7UBd997mc+UGW2mVKcNYOQa
FbgQMrPKyVsIsCa37xkBpIYArcxW7Us8abNPBFq518Cz3A2biIido70FAervXx6jqncfr+nJx8pv
81DZ0qn1flUkBdpST53efXz/8Qigq0w/DZp9nZQuJwzb6kXaVGcHyko8FcZarWLBIWKi14GH9Ldr
AzvBVOASe9aw9QPfQ89Oql8N5vt8TvEsAQg8/VMXiZSNVNGv4aDHnK2ngQs4WzojygNEv2MiShUf
tQDyn2D4L7Xyde4YIEEm4q7P+B23uw7bAKyxK+dmwGXhoIVif4n2jpHWlOwH8TLH0tyTadmShs+H
+W4xVHZmuQPBXlerqVuE5Oo7zt5+k2KJQIulNJzSP1zSXr8Hopy9p83GFear4P4FYqbzIP+aaaV9
CKIM2IWUBPlwqW5dgS6U95OjvOZ/n4p79c1rBrTg2aRLBbnBwj7zYC3HIk7h30Bl6cIFuoFx0GVP
NLgs+vjIXVQJ4gWOqUYERnkCRI5jaVidHp4dS8rZlJwrL18opRGOrdoqT5xc8ZlTDHJ+RKYwW49k
NLAh1Z+heilfYbGODE/gBqkDpHN3ALPgShhjiBRN+dB0pruy66syBuvJzintyFLvc0ukvz3Z1aYs
OmGHjZlxGBv1NRtalkPvNDPeEGTYVwZBd5f/Cr84pCil/RfsuRLECRxS40BLjeyergdJQ9bF4ima
kEfsFWVXP6O2pGNmK1IKClr+VzRl6A1rE7UmzGZpGp9AcA/k+2v+613rBvnT6vuc/pjTd73eFmZy
7voGd6NTFLoJFmxpvkC4szjb4hpf7odUt82kKStMEiKbGpAs675fHQzYhdsFT91RE+eCrBIzly4N
DQ1wlrm7iw5yPspNC0aR73vqPrQhUziJGAhOXWIDt+S5iUSSofMrUxMhqOhK+3WueVrnJM3vM3lJ
foYIoF7mg8sktpKb1v886RsGYbRXutWgGYRwrlxEAlLVKwtZfQmWGNqz3C30IP3YcT8gVvS+cSL6
a6yE9/KhtxD0Ol6uOUyXgGmJLKqTCJ43XfYRBu7IyEOq3Wk/nAt98i+XfmUPAiFb6AkxcRNPVyyP
96ndXc4rwRlwBLpPWC2ccFfhHpQaCBn/6E/Zbrx3tM6Ar6BIroAKj/ksMb8UuqgMT8yyGd/dtPFD
zcytq3qdKchUWA//JNuEF1VLlE21CLypHVxLnEi8gpyzfEqu2crrtRVQiB6ygO8B8uwty7gEeEfW
uv8NJ6Npq/bjAKX2PXEY1xb9OKtcfa/7QcHzxRzFUFwOTSEwem4IqEN09x1JkxK3WcAu0bRAO65j
Kb9KCslyr8FQNkLE/weADilVqeTHbmRob7YmGMma+iUvV3ukKdr17y4kQnfwhOig1g+PIA/lGBhP
nEg1O/jEorcooKsYBcbJXG2q7izBAEmjO2AP7X/o/65qv0vu7Q9GeA78KkM2/K+M1qlFSFxfOIjw
xjkQLxsNtiEVHifu1ChAzWBa0MUEDz0Vd6P0B4CRFlNYgZktijUf994goAu2eLH7YadJ/21gin3A
5OhvF2twsYNq49brD4bD7sQrw0+Q4i9rl//2Rt3MrvvmTHYqdDJlvqdAv/d6tFpy3SpKwEmfQEtd
XHa+qs0l2nXbq3JFhcuLkOjMYC7qQMW0NyN1gitapwPWF1ZOuEoLKDoXxnvUp5UnkAc0Qgaq+ahW
RTcI4tSY0Ym6v9I86etWTrOb4m4ZsPX+IO54NyxKesj5aDNdWecPcjHscHnqjeHvDX8KiC/kXbz0
n4rSlEo63hmZevsqcEZ/pbTGKUcJeN7LHdNZvxdbfXXzkzfQy3EwYqQKLn6hvZNBotfKBVb8AVJH
QWP8bv7GWw9/gQBGpnno68cgGaawuYO7YGgWHiKRUlq9GwsFkgPCXKJahgc5QJEaBPXSlYIUzvzG
M7koHoJHF94oJRlIGsk7wTfCurtOehEwZWmm9LMokDx0vKMWu8tj4Jd0Qzgyr0RgfQB5JiH5RuMy
DLIxBclOwHId7MlkEp7GawDr1afm3AMB2hRQBrRfqug1tMr8gPIwdPzTSKkOZRCYYCQFLwlObPrA
FL8OhDHohBXp3F5TWwvNWi5RUyUvmXYFr1iP6MWpBtBUnbSKr/35PHkxE+1A+gjlZr8yNTfNmAVM
sAQU7RtKwVOs8i9xgufo2DUJ/1nerl6GBb45UuBtzfSdWrCSCnUiDBnNUxkgmLC/E0PaO4Gv/NoO
ECqmc8LVBIzTvv9DydZWIxgSepBmyYmbKrONMFAPIBp/fyGG5GfdqQKbWOViedouDVet6q0YzEoS
qlEDC2hcBYIDsy1sbo8xpF/nsZUfy8Gbar9e6lAPIdOyT4j04cylaNpnLNTb9TmvIhPQSjjU0QHN
1Q7CAQTsQ/nShi+t2sQ7Yef/NLNindZR8AckAVWzKd2hAaCL0pp+o2vs4dTLpl9P7yq58v6EypIl
m9aF7RmcksL/UEf2kWSbdQIQZxJ0Ax3eQW1q5yyeIFdgAMkJp0QtgE8XHqqHl66KwKDV6nnCOnc7
9ZoN0hJp9Z8/IL4HGU8lRUEZYYtiHg904SYyZ/pnxPRbxM8hNsGEdtKDAbq++bkp/KAJ6WFGgYSN
pql8zS1pZYHZXllWZHhdAk9rq1YJm6JP0UaZeP9YNYjqk9xXUGfQsuhKJk7n3Ajlt6ToF2p9RxpV
jOL2gdOLFRpuKSV+aRNiG25vlt6vuISrS/f7FU/bm7DHF3AbD3u4dBhMKk7VwQXMaR1xv5c11dR+
UTYVNfLUqe5SQ1bGHYsfiQlie3CbRcK4yf+H09D6dxiWcZkvKQIj+MYYNt1uXUvFleV/gA8EwntV
YJr3HcU/69/RE83tS9S+QAszuWrB2EzFQogYQ7WTrNvivPlJQcsF/cENE+fLw0I2fyuiebbt0d9i
JlQPIswkBX9WbJmCLJbkV/0/5JYrVNcDjYJZR09TvGvliGGrPfGdlNNrjzNBduVIP5j5RJopBrs8
WRXXH8iV2VPIYl+MbZfkqd92O45e6eOnyBLT2PagoHjHUx2dKD8GHaFfGtunNg9Z67vYsvIOvLvx
jN5zQGwEq0L7OraB7Gf9VH0MJYi2jzac5wuoIJZ/1ji3JXjAINFHBaIvZzwFsQBm7kldYwKLbGup
24fe34XgWozWCQniqFYQ2majscnyTxonllf+Pl7AxGNosSW0ZemCV8iyOHJnxXhhldbnVa83SZgE
RAX1h83AOoXo5i67lGD+XrFBZyOPKviAr5GWcEkPyjQ88nwoNZ63cxRH5F0oA2EhnJXoLmMz8Wv0
AZnD2I9YyQ7co7wqPlOGMCQS60I3QRn0MYZagLhBZwa6dPilT5pZjMy8ySD81pGGoSHtfbkin6YZ
I1Ji0FyJ1pB0kN5T0PdEg2PKtAB/99XJrK92sOjUtDTBo75RATPtVzYqbAvpFw1nDs6WxhLy4ZHD
zZs4+Q5S5BezYOpuSTWdO2JFFb5p0p9p2EAd7L7CF4KPYREK4pTp50Vwp07uDC31mkkwVmEUmqK7
oKIdGTQ9qohr19UCSxglznCH6SPUkXZAD4S3kfZDVgGYLJ6SyE2pstlXWc3wes4PT43Wh9xBsTVR
sSIUI3DPjrdVUyTjboolYlbGq3B2MsyO9A1LdU40BBZswJC4S5gUt8P3tFmiTAASsWGE7/JubOV6
hfZGPpbTSj64jznfnak6NkTLqMATwbUqQV2hNhIf/L70gZuYbHsmtahX1IcgbRq02uClNayfAw/A
dFa+UFmxt3mRebE2t8uUorqGWKqa/vgh81lvkUw43uP6QSNn8+z2QxzhnUGkCeJcPJ0LCbtCtkoo
xNYptJf7Xk4ljuNsLJrcS+iHRlKdTUut0Vhnic+F2XbhFFc9XZ3m03I6Rm5OQ9hibTGKnezEs6gK
KnR5XKTmxp9xzlT9MyE1jSIZBLntT5lwHYnITH7ayrrJVSAvoaV1I471xPWnpEEhVfBxU+6cKoYv
5G3LOw2atfGNeLEy3xB8sm9tzPr3LpQW78zxlEOAOIn3EE0tggzalplzCJhNMeS6ugxr0DhwD7vr
GRlSqGD4X/al8dwugC1iH65OtzKEics5XeXAIAFRZko6T5BZ8u4QbIkkKkwVbMP+rGnMHILlzgPK
nEUmDeG4/MjetfsgcqIPEEXdupuVGbj4DwpId/lsKwNoUocPwTWU9GHrM7gq9yVjxFm+4XKPurUy
8aKNMB2ezVEnAQ7WZCWTfrFn4RnRrlqbEW1IGQrwHg5ShdFTF9BGMB6TluYL9hfcQvUk+VjXAUz6
0F7XnCkRhH0CjBoViiq7k/WcQbsO/1XzhJcJG/eLO0lAOtzf8jv3mGe9bKdnOE2/e3uP3np5Uwg3
U6npBIkenpTNTo8J8v3tpG7/oBOtIbelPH4lo7GiSqHAHvsHIfNH+YTwEB8ZDaxaocwIyiUfGIyF
joaL3ZQUTPB4cbPDrUbn1l4AF9QRxtNKK9eeL4a+8H6yyCZ9rwEv1BDVzqphqrIPgKkl4795eiQI
jCW3err63EqU48WLeZSbSs+Rp0XgHvsdN6MCudH5mkEB0R+hVSTG1g/TL5V1Brxaje2IJwaE/YyR
5dF2GZOLETYI+tRCjlQqya/uzZHKHtk06W5bNYNPwvY1bZiECAALhGZ/wFQ6q9lZ1cA1WRPvOMN6
FiWUslabfM44Su96N0hW9TrUTZOCG1FUtafinz/o+BeEZGmbZr9M3dLFoY8NupSdu6FWN1wvBkAD
PYUj9Jv/YMDUM7JsrivVUBsX/sGQdcBsmJtyvga1cAFrWZOtv4kwhJlXW2KwLJVm1YDQUAwDcnN0
f96LowMZ2ij/wcCdj3Z8AUL9lGquczum/8w2QnIWKkH1gKTd1DZePZXcSzv1L9mksCDTfyNQGESi
DeMRzFTb0c8WD965ej3p0pEGd9SLHq7sOj9wSG+nVwQVm0nbN9d+MXa/hXuxyJOHEz77uIxRIkHL
lRfAJLHJJHz1JB31kG1w8hgXMz6BXjrHuJbY+R7pbcs6tYi8boQUnSyTxrMXjnQLXEZwbNuijpei
s7CkLaLoUxNh4lsyg/qzhILsP0KJ9RJBEqWAa5wqvA5j07mSNaGRTbiQ6TKovWqJr4d6EZ8VgiKD
QGOARFknMmVa5VPe+vOBnJJjCWfDKJPXW8C9QJzE2Ll3i3+P7tpQ3Ti+yOLCHVMZBgoDm+w/ztJt
zfLLInm3VE6spuXdFQMjNpTHUoE+xGPCBywsH4yHmcPBUWF+zLriLddh85c3MkHGwTDmU/W4MHgI
HRFuRudDh6qoyKfm3+dRmyp7kXcIhzBDczX7rI09oJLw6emgaoOoj3bHlYUXJYbU+taimKG2rG1o
FcUWkmc95tGbiT1Ci12j+5MZK+4ICviF1dMymg3u8CVShqSCe3ciXOMUFGamhOW6ZzZ7xrtU5Elw
DZ2hQ3q+JeDJOQM5h9NAqgWJViXi9GtZSHO7OOtV/8KrlaNKxnubXxO5tTuoBraSko49vCgIcyZG
3ua1GFftIYUA6dnmK9b+Z8eFgvxxSRAHb5PgCKEXz9PX2Wgbl3cf3lwfKLxq/u9I7VorISO0Osbg
l+KsEqHQAyddjaiKs10WB32WcZhpef/PogAIQ9U7qk8l6HHaZt6TCDOo0VONtxdCt+GilNsczf3h
f8G5TqwOYfvzPKki5qK1dBmfab0Lipv73Rv5UQYI4jOzhqmTZVkqgMl5Nu5ODRQBpenHnLR5ah1T
qvquv3i/3wN+C196veovv5FlRFUkn4KxJn373XjuwmaVK8aqG+B5oClig86ta/4/kywVfLL5w5wP
+XQCH9ZAxnUmuxeOcYrd2AMNT1AuDEJsV/wjRPllFn8xpHceLlBQ+E5baeWWS1cq5ONCeAhPo7+R
GygEuYW1qvi5LQ5zUQYArQGRQ4OGVJoXl/xalMjyOpBzX/uMAIIQ35ytaE/mNtq0MpTh900e3IG8
3k6A3iwLeWkhbnY/lwneR/5wkMiYJR0XpzGwDjQjBEAJAtkp3iCozocMfsdG5/2L6dkqOuku8jpS
KtrjjLtSPPQwEx4fGL96rhmhqI0NiiWZ7qvjZm9egblo0LMm4v1BHrnkTQdI9jtAN7fftx/RXoNF
cQwsefDAUFn8duadgLHABAEWLCwal2BcWS/uj0cNKLXOX8bjMxxJyKGDX6cwl+qAHugDcKXY+JYb
E3aPDtOKrdTDokcoMpW3tXXBuJb4vUI6Dpenfsbd5lIFYtk+YKkrYaHQvFXcihnJFC8smVGiB7P/
L2XIaMOhrhCGDonmv94x2wbXL+7A2VLkR67sMRVBPyMAdJmLhd40TpROcw6pNKU3t/1ajFYnSHf9
VzjpSeP0zycDCpzw/tMKBGSJfMody8geGW3pcttkTNvl0sHd/WZuMKe/dtL0ZngI/LT/mHCD0JgN
T+/DlSr4ZMqOn4KU+nJHsBS1qouorogFE7EynHjSzecwaBzgUZjkSt1yIgvC9RpzJcwUdBgEINmm
UAb+rY2ruRRsSLGmtvf/DLkeB/8+L2xGvKkBElZ2o/0e6IuItCkZtTxfYUoThDaT4BAZMc3E8erT
6F1ohPU6Yq3ovCd4/qr1Io7eg7UGWOJIMRj8smBe3r52t5UUd7uIWq89KIc9/r+xHdlOrLEPTHCv
8MtC6tp4znCLocRn4XZvrOzySHQA0EYRISoIvEBsYo1DinRNiE/TpaknRO9nxg1h55Sg1u88Di+3
k4UpG7tni1jWnD6H5diRikBHUmNIqOsB/qa+ldGyziew8dCbK3NQNzVrufDH/o0pDdriU85jUFc4
fTXXByI9CfKr9JBK8JanWnFlzLvJF0lhCYdBVq3tKmJkaFwjK5W787aRSreL4Ma8WzvFwCBq+uKR
cmV7GlT/UOsJoJUxbl5H9UQJzxif1ZizGae+9NgrA+2LiRfLSTqnqKbgKXhIOZ+sS8Gmt130JXk8
s7M+EHHEb8quOB5OM9KOyu/Mwu4T42Jy14jSznOp1qlrzsSsOy6Q5lEVKAFvfbiAf7TBQupoWx4+
oKZi1zGNg1pCN6hdcqdL5r5kFFzibKAkrQKZD4P/9/sizFDL4rlOA2MxGokHY6AkyvxqjazFcUsG
iyHhkbdk98oR1DRhgac8PEou2UnlCbC86GOBxYN3msoqfcXC/bd1nPY2P4izxiwVq0Ea+dydqNDR
Y3qKF6aOUpdJVtfE4EvjmuJugQ67gFkUAktN2hs9HOTotA7DfoMCNMBYIZxoImiXM+JZFbv0xDFf
NzCWDoit4+FVp/ykq86g3AfgvF1stpmU2yb6Ez/bOaemdW/AMMGsnqkhywVG1lxtRGrwkQZS00/s
GdaElv2nx8l9KcxcqBfwnEjU3/seWtwMk0vX33XZ98fl1ImchEl6h5qrCHWpzumhaaQx/NIsYWzP
ALguuapRsshwfd3WzpJIVfBuWQh0KuL9xv3ULWevdHzvpXWJrkxehteH5WvwXknDh28rM6U/rruX
4olF/RJ+i4ByYZEzyqbw63cdvE2Lfe9tGVyr5IMs3xCvvte7kT73Q0gGm1/2+JIuVD1crgQtpcqn
iKPyo1eJc1V9e9KkRGD5Ja21zgrY6YFd992zqiHDnSA/hkBMCTWDX+pVBwqv939QuRb6NhAGdRIQ
BcPgMgffzFwADIo60SEl9VP0DzPc9ReihArnoTX+L5PYBLwmxO8v+rsMLTi6Qkj5IouWUKEnTDUe
kQhw+SUBHHxF4RmHsHDOvJ5fGalS+JzgYB0vVwliK+sU2zWevijnbOAKadzbJ5BuVWdDWkpKIPcw
TdOq0lhXm9XU0SU8L2WpKd9+aUsr9fkjei+bJoT4nITjcMtuEnH+IDlF+3j3bx3o1V3dFu9OPwgs
xGygcq/YSj4s/hgpftHkuG82o4o9kXSfEhi3frn8kMy+TdQS1C3fHU53CYC+Wtlt+Tawju2r1dzm
nTTQvPaBghtzqQqhLu8mA3zbqwb7a6Md47SLzKrRe2WfwTlGiDRlGsQhgPZGp8zxHF0onRI9kBx7
lfrMgODvI/FsyeqVEK3az6cRQlYWtvtL8EUv93wk+/x3wnvGdsztH0SW+cU19hlWgVa05TsL0+Or
Jw8xBuTVE6DFY4KNuw3I8qd628pawRSxB9T1AVa1E8RGp0HZNRLN/awE00JJiNWsGn4KsIVB9nr9
et4DWnnA9t0EMg6ISFsv56wZMiYg4pyB9x27SyVXvDrbVT7D9PS5DJCPFotZDCWYJ6OTuWVyrkB1
5Gyjqu9iqCT6PoKRjRu5TLTFnsR/mOS+bM0RlLHyP0orefuhalBHk4llrfqhHvW2v5KO2Gt1UR/W
Gb4/mYynwZzdxyB+Tgh4LchycSq9zmN35a2SjeH2k+yLhFHG7vy0PCezs9y4auUY+Xvo0N57X3i1
yhyGkef6/5U1Z5qyHkqjuIubgmP9zo7Rj9Qa9owVUsR0l7svtaSOcwMTU5qvu/ch5ysr1M60p4Pi
hTkIEdJkOQ05K5Dt1hj4hctwh3iqvX2oV8edATP5OGzylqWllhybvWZxmhPMjdXvVOYaQh5g3sVJ
OVZ6zM1d94sp3wFjliY5xs2rF8kHKme1WdVCsa/+bq9Ra8UeUX/LNpQYxX1cKWHATPL4HnGhxjDg
/mfHkuSb/U1HsGWjxw++gih89Ed6Rx6e5wibjpmn+2q/Q7XBL/OcEozGGWT9+AjqLsM9T9jio7wZ
8y0riIGrkU+osmZWTywXh6o8Uke2dpeBp/SVs9nbHpAXk+v0t+1pRNzc9F4H7ycR7MokcHDIHkMb
vwQa3GahxJt0z6gzkSYeI+Xvkht/aHzRTUZpjYbZZSSe6jnsMili1O9sLVo3t03qLjPVCzHMgbr2
fXNopIhZ1R/WicBzJEUF7oK4FR8JwpYoydmAND7Y5KtFxDOLWPeYfx2aUhwm9TsTY/Pq4rAMHLzJ
VmGnlB3rS8X1X18aidMNmKFTf756xL4LAQgvtlqrGJvY5l52+3Hgs53kwRL2EAG1xLFMDOrfxPgb
OsNHwSEKXY47BVFATta3aC2UXJPfg3Ablf5t+BZ1VxnECiM0gohC1BPwTkW3b6CZnvVZVk761+dB
6/xA78jiEXdKHCLls8Z9POUlbWhoVqCEyTcHW1oLY3iIsl5/FT+EXbTnrfVu5rZ/abiDDa3vCgAx
hw+QNPFZdmL4+kxs8PoBhzbRmMmHSTPa/jIsw5Swmd5GtP6B7sZ5BacHO6cixz9a9LWFiuADMJ+n
mBnhbP9+VKnYOaq8S3k7DkqdtdYMydMDUGcuWLN4J3fixq1ipvDTNPu+FJ/vKu8IhrAy5r1xFbCD
ve/EIf9dBeKqok1pq0NXIOxF3HWLA36EJFdhloD4oaYmZ/+/KwzImJEmZqpAq7ApGnPLMb20B0Dg
KGxIgCzpqu33/96m9QyaLiqlwDKNTEoU8ETWlxx9WhTwYZNc3NPQkkos/rZC9Hkndo2u1GP+9xba
AuihjUNVdUF5fTPre0Ie9rRCrDyqjPWI0NIll2G45318dWFb8MpPDewkG/4B/RY/9OOV+NRfOFk7
spS1JWQpy4863q5T54sOvEvNch4AwbMS0pmjZTMAUYeOgHUyPy5bTst3AU+u0p7lVrboVVilO3T4
mb1reSZdDfG2mdKS+Jn5b+Q7F6ErN/5pYckPqBIj2C/Y+Z10+Gwnpn1YmWZLeR2edcBoJ6Bg5znm
oK+TURczDujbhtGRSnKihKjFGnEhGit9SoAkSYuRwPTzIameiI0QoKnp6MSP6tmN1URIFvTxT2aR
viIoomFdDmI/XXy3qY9SoFG5xJ4UYnh9/lJP4ASOxiCtAVD8+J7VuvRfNwxl1PtFDVxFxw0et2FR
EzRUy5cw2/N9QUIxZZ7ob4CB0GpL4q9kWA2lITSYJ4prY43SpIqPiDVghYKnz7409+8t/1fGdvLb
5Uvoi9e4xizMdOe8S/8oq5qdPhx0FAr+SDljZDuBo5qSOpTYLiRBSYbeSKaRKW2wiEezwFfOL4VR
dMbBcYMVNCwswbdVEaPO3D8TYx1NO2LcesvItqmmc4g5Hd6N0sr6qKrCcUK8wqr+Czzrp/KV6NSY
urYDIkG7OX80QHmcE5KgitbhFIg5vA8tapDzOEcK1PnX/NZZz4Oq/f0AxVtRVxVd4km3fsUL5TET
TzyxXRl2GQr4SlSBnK2dE6gyIvm8AVjMDUAY96kUUcVqhWf+YEB6l67owj/e3z6VqQFvJlAX3GOm
5pAirsSCtGbQaxmgwtVZjt+lmJOPyToMDRSCpZ7At1VC5Oz8FbW5cdcltOQf6mpHRzc3l8BXort8
V+605MYWfVVX6NgA0+8PrMHwh1QGWtD1BAMb5xY1DBgG1EVVbrgQPlh5Szl1lNeL8kHPxwh/LQL7
v+FXSsCN94i17zBqNq9o6YJrssFw2v+gxcM7o66oGxmSRGta4wmuSq/VkPx+MTmyKDpoPjG54DGR
PhHepOf/J2DQSnoy+QWyUev/L1rNdtzIxfFm6ZwiQJZxrG/pPxwfzfloPz1VKMeRfSImO2seC0Eh
GmQM4suTSUmjhZFxUZ1SrUt2jKLnMv4s7YVM9vJoxQgj3VlB5o6wr3zac3CFJByRQ0rTcoRIzFza
o154qGwBaB5xyHVwIxV2X2eNcCpRz/d9po0YMh585a0e8c3zI0aYcTrMjsA1Hj8pSNF5erDdwIfE
PqMoBLsEKMPhvhJbqFeDpy2N6sxHpromMFIGX5YFxGByd23efTGgt2NZaPeMKhQuCRHmbcG9cBwk
P+vXI93ukxjkiAauRN+D1miNQ1h7LmCU1mLO6wIq3Ea4yYAYVvpCEOmTE3fPjcmniqczjsxEU6xc
r4FK3bSPjz7vUvHNHVraeAfrKGEaYp6ZH/m7LdzUnwiTOZIxYdzdvOs+wxTKTvuoCwkTBGyeI/aa
317ALrwEVTP/oRamTcFQGmtfia5MTzuZud1tCDuhJU07qnrRTBpXjXYn6em1MKym0MM6cUIQHOAx
0JlcvVIMxuH2tO0bPuAWDe9jAXk7wod89Q3wSDlBCbBO10jue+DvVE5U9GGTAsEGfj4kF3zOewX6
/TUKYcn6Y5N3hB7GhPyi+lTkd+MnMfTev1SkEanfNjwMFqjuNU9w9AdO+YKV6c3XWY59lgFkBD90
BP+OMe39+ikzv+bDGmo1rmtMrU4yK1p/dgzvjmsp5+7KTXbk2IXtPkYT2CMgOI62VJ4NU9LGki/0
+xX4n9lYHFfJSHP8N5n3ccLtk4c5vrumUalVUUdO+Q33objZEKRwv2Lw4Fqb6b4hvqVCQyO4ijJu
4McyB3qW78R4Qn2Qiu8rVFSAgXzLrdZydhlK5dFoUDtpZUgsVWH7stNRgSg5GMiY9T4zzIDeFChf
2e8nlqlkph/KLG9PiDBFAtO3fJ2plLAhBlgDZEQ0pkwcVCambHl6K9Id/OlisHhETJKjgGIdAprz
WUJhPNlxBi4H/FkrQHxPKLJVd/kr7cR3STp7SyDNkkiaUOldFp6bJJYvIwXktB9cKLDOOg3fWsyE
PUVwFEQO4ERhDf6i0IpKs0+puyar0ZCtQehicvKDLZNjo+TurfA5XxgstXGxlN70NEu9uWflHl4t
vbv6fj2lwyOHFU8g/nitN3FdjhfAaLGono/+5WlcRNAMrY1/TYVkKfDbNQcMlFVrxITt5wVxq/Ye
Jfzzx3F8XkA9T0oiE/Y3wnJALXRf1k9aVx58mpJO6+tTNwEenOsTFKTYORc3QTyZ6bBelDdlvjCZ
i7qxZpbx92M0M5JIja+ArkmzvTotQH0Gs1gqzkahZkm7nhusFOTCkYld3v1bmmXPB4QPa8Z0Jsln
XyNyxkl/l+W5iNjjZIcn+lzxNBDVEy/xcigmvuUE4uZkuIojUEsoO3a1BwxEC3yVe1eNU+E8rIqy
P26G82yw3rkZh3KTZq7+d8i0eaRNqGQzaeWWZ3heJGrMXm1bfIaGVY+VDWjnFDDCjiRHATt2aa0a
YKBhbJ4j+yXi0eApex/f1AdnLWiqUduhMA+YyGupDE/oCp3ar2EDgXCl+UWhSfdwiufzhQxMFsuD
Ybs+TQugEVo5qIZJBo0IQ1JFaEhBHpiVQbF5222BmmpnG7q/r+QZpdhf+vUTk9NIt9YIqvCTviRE
7mroGP/Q+7pzI3YlGSuFHA2q8sUdk3Jf2pU49OUK3ciLYT9EkglOVkKR3PilzIZo6pePqFS/xo/1
PkBhgZl+riArdN5Q3tB27CaTPIKzfFJKVszAy02q19Edv+B7vPfTuG8RRN4+dI4jRNJ1pB+pe9dE
9xhLmMepVvoQhmaACl5wc0Br6ic4fxKZGEkdSITZnKZFfdB2gK/friKMlxfYCMTEqnk0cbW2Yq4q
PSUXK2oRjsMhPceK3WGDmWLy6xikExtff5sf/hUBCc/sfohd2sKSafD3G71arU3s1evIJ/0Qsvaw
/SgzZpjJkMX5JXs8AlVz30SiWU2WNGa4sHVOGDAJfAgKFvGyhr47/aSPT+sZN8UawAwJEquWe9k0
l1jP+tqKlhU8SrgjUhfn8PiL2tbcMZfaW11TlQsKYHqqZaa2pnSPNBpkd7nRO9O7VK4oNXR9j2ti
482CWpgdzeTuaw8ayJasoX7en+grFSqgkd0xUA7EncLCItQNHUtSnPMDcbSjnmoPIJ5gEJWiT8b9
66Knw7V1NBZgAF7uUMQo4oapx+EmqD/sXixiL9aNqr+N768m/svsyZLFC9wA2JeX7QEqibAvFB+l
ssyY/jVuN6VOgJdEqSUHRcWjltxYtaiMSVmusBVPijqYL2anWj5T69ZFZzN6cveTYn/IcLy+tT2O
RR/jEEAMcXXksvhdAcY6gdS7EoCy5bH9WargZSiiiVKdaCETrtFBZWACDbMp3FaDJ8cFTrevDBYo
6H2esJU+lai5ez/1GkXDDuckucZ23EzeNSzTCLaPJvB292k6Q2YDZExaSeI6Sfxfm4hAn7X/z91Q
MVGgArQp/PwKr81ioAhOuGHPA+YCqhjW9RqIBfR10zyfmbhMNS3TczZOb/1SLSjMGgLXjE1GjQaA
p2wKstVk0C3FG0SiXuuVkiXjh8rZhjdYYoMtOozzehNiMdvs0snPETERJNf3bA09en+pT5xVR/1r
Ulyl+UgPjd13UqHiuRDHx+quy/VJMzMWtq00FaV7crfBcxBuBXTI3k35jUOa0tJZMka0/VNtyu4C
c9S7/hH9su6P3HZhMg+r1wFvt993UPGzCDLwF9Eccw+3UtKu0O2kVMJhk0dzhohAbqTwEPq5Do8L
dMVqW+VszsTiP7+d9deRUaATEasjaLZGv1KYvJz5uSiKmEmEZAfbkGwYHgeu0oMIMFhlyJmIquPH
4CG0zLGtvOhyO+s3CTjVKrEGGQ4H9mL9GIqJm4zmEyfmYXoiUXbqMspT6+LlBUO8pLjvF/P+Z3Y+
eOTE0qFue9Fbg+XXzwtz3m4CP0SwDi0Ywvzu7c/gHgnCuo4sNKoCgQxelQ4iJwrVbneSyTiN8ezE
rKp5ppd11UFRIi8eZ3B+1srLfr92ddYa61I27qi2HS0xAR1O7m46TZ49lIF9LapRLGbWhatFGXNx
Oz/1IRBaPjrB100VwyQpvXbHE4imLdT5AbKhMXCSWR/Jw+EbZLtN4tEcbRUbOegr8+kNQdx1Bnid
NOFqKDgh70u8jx9Gbz28OyFT2CoYmXWUUeQz8uav1L+jdaUVebANFZyDou3V/z9U5AtzeN8F5ZtH
vIGAxwng/aBCD7r3MtsFc1ecx4vZ/GJy9sFksWmnOM6xGsYRccr59RasTiCP0Ert0kyefWbf2/Sy
2+L81ZiIpMB4hty/yQKaYtLXsUYFH63OjUpi61P8fX+z57IgHad2ZDaURwu5Jj8F/ZAIAkbKZ3NU
6F9bSdsrL9IkzUBVIOtmjlDP6jcXn0hjyBWpxzgaTTLFJebPgryE637gVcaApW7ZmQH27Z7QVQqm
himl2vzuUaBie1TSgywZafLg8vgVqCU4i+tgnpd9yE3BA2kE6mSzniCPtMzKqswffgtW1mhb9Aaw
efHw6BpSTUpi9dNz1RPDjR5B4mbiS79n92nq2TOTiN3nv4voi6FZeqKj/KK3cEIG/1JQBAUjAuiI
EE+C9eIYrunCVfFW7Ucr/IzvR5uc4qFdlk8nOqhQRaDd3/oQO+dhG79NO6FYEeyHGD5zwLFKCrGM
ehYTOt0A/eEG1tCevThMcr4cDTOB2xfWnmpLD4k9tDo1t+xMalvJDgCaj7JKoYpLkYyNA+3gq3KB
3qoqHhSkEbKNBP6OhXQmaeALYi2bhcN71nlfQhTL+KVacycM51UESER0Q8LtV5qV1iQt8aPaq9mW
nBIbZ8AlBODH/UzxN7mVpkFZ7GZynleIV/ruuEH2mxPtXDxnut27XFysTkCRP0qi7CiUW4rTzcwI
5Mj1N00BWdZiItqV6HiJmEIbCS+XSvngMqgMtNgsengkmXTO7tlSdyYiQ9UxYrorL9Y9Sapn04Jo
LhZOUA4cXHv6iv0HhXah0e177Jgr+BcdaRLTj7YwiEyj9Q9RTQR4urTK5QtLMO+UJJ0anXZWuV/P
mhri06TvzqEQV5Wzc8IeybOYX5ptOMERl4Tzu1d5hK/arCe7T1ZGeLhJhcTqmLOePCzESXTaiKhR
zq7G+oOGug9g9wTliAJ91ZBCJoV8eGV912xcuy1c2dqVCxqwA9wCzFKCUFeTFv52rRsdYD+/FzCc
AaT8MAIvSbQGRktVx05re5XAk6OlX2bpGOw60JWB/3B2ZJQsyJqOG2m8pUdUBCSVwXFooP/cl9bq
OnsO15Z5T9sjM+qOz8lHMZYqsIOCfWlWxR3V5IuDVrbJ528qAhBRFPh2nMEE2zwuQmr3D7TJLb+M
NYLBXASR2ibsmqwhtl0BO438j+XmJFv1Bspl//E52UPW0yueVdcFGvJbmj/OiKEsBOpnWzKA2LBO
eaKhLLJdusBNrBsKnRaNxd7P1EL8qZyR1jiqIwf615/d1K7F5qU2KbLuqnJIc6iXSCDEYQ3T9EPP
CgVEt1hbEjFGz0Irdpc6ZmquYqrcnkgjdRsH2mJX6+EdT5pLe4HlJhqP7m1+cPmNKEA7sX5lLXWf
wl/0INBdn8Cgb4aOCRpr6K40PjHFMNyuUMQ7YQ3j/MQKt1m9427TCPQI1oFBwzeu1/X+jA4tEy5z
8uRNfYi9bA8yIqrRLE+MZX2fMmA6wssK9Bj86kLVzt1sbAvQlkgrOyT6REziBSNDV/WlsRVxj76z
REToQ2peqBtHtZeE9BcWcC8mQR7qWoYL66PG51d9bgwbtxoZ2P1SKz1rlkSfBVlHXt/LFfLSTutC
m4BxRdNE+ocnLoCw7WyC8kaa7VqYOnIHepIROOgcjWfaRw2Kxj8m4nZg8H3qnxanfyHIK1izgptz
/FqLAExkfdf9BBVI7J1pqoTFthg+Vmt2QHCtgr+YUJpyNgUGMp/+f2A/aEn6MxufEh6FUgPvDBtK
gA+8kfa0IMedP6d56HIH3nTECGZKLFB7n3o+5xX+ydFncMBWQfWSNjwwbdic5gwDhQLc41GSl49z
gZI2Ci3d2RRNVyBGvd8tqoxUnvVhFmDIIVNchKVpJOjBFHan5fRTgDKaUouuGp/Rs/XKtc5DjEJp
vNYryjybWlWX8E2Axy7DVIz100e1vY2hwUsqlwdx7RdEOOMuFeU2ckIWwtsdJODzVW+aiDk5gCT6
gnFqLvy1fT42fowWFsLlRhgMTujj1nrjkHjY1gS68AYeAp82Hwaseu5WKtaY+Bw3W1Q7DB57+l8H
3IuO1LbqxHux8Dk8lrGk5VoWIGXSfPxyEjB0ViBiPbyww4QspWaOjvxnKxTuGeCTTZY1FAjVphNa
LthGGK6fUplbyK2aPLE2mIZPbUUY1DWCoPpg4E8nZcnjnqMkoW2Z4wHaclovH2O3acqto4faVcku
Mf615/ba90v6W4nWd2zirVoY4+lV+yhaPcLlm/n3auXHtNy9rKQx0QCyv2XINBypVSQ2QgzblqhE
LwUrdsX+WNNM7mf76ln1PPSOwav9oYwSbaSzIr56V2T7Ypoq9D/mnqV0sOGwfNYHfjEiy1fv5ptx
Yv2c3gpG3nIv8IIXnu4GS9Xzc4ckEr4nkeXw8t76fdy64NcLNxzPGe1BFtLB37Po0dDvbE2To34t
OOwRDm/CXBE03dASDY0RBxpL3K6RKotjRI+D/uVr4yHqlKWTrMBpLfwv9UFOCBLmviTtdDcztA3z
2YIf0PuS80Qnkiw3/ScOFKevbkJs7Mq5tx9P3UFv7/ZRR91HD//zKYgQsmehL9n2xoVDdaLG9l75
PQrgOEHZhYCXLPyN7hruwl3LQIIxkPHktNZ7p1u/H2gaacr966ZCXFLVhhrTRY0gdfil7B1GQDoi
K2AbOryqSTXz7VRVOqe/AlRcFVC/o0z8zYwYDiQy2Ku+Pt75A/rBjeSi6LINblXWqu1r8NsOZf53
Vd1iAfUsWPEH/6qPuZ/dB0+vhFdilg5X8gT+dN2Bb9q0Hj/8fYEs0KdeiykiXjVVbml22st6S3vT
wdcOdDtUFDwO693s+3/dFTxvuoxrrkXINTIa6+7256c0RXzbLk5Ec8UE056iiNFAc5gM191107pQ
3XpVqwo9wRid6Ry1q9qiod0gPv0R6LUjaHwTlyykTdMiTcus6+/vAx6Pj9zMkJS3scvwIzusovFR
UB8ZCU0THHfwPrFi6LmWjWmLk8LCY+0zAPx/pZaJUO89C/QvlV4ib9Htutb4prKOEoOuhVX9eBh9
AZiPaZb9UTrfHeRW+Oa+lPwxOQMdkL12AhME/AXBmYzFHf9v3Gpx+w6nFo4qelCMDmaNYtTQ22f9
fCwP4ekdG4/0MYj3d7IvvBj4MnzYI20Fcz9YjedqsfWEu0TB/SwOxdPD9EHcFnlw9xRZfz2zsDz4
OxNgY9uCsu91DjrJTRL7I0FA77DDuc2U5GPfhhO3V0b3mS22rHFFnyLj8pV5Z68i1HFMeD/fhppY
sknkPlXKLNktFsencbOTAO/DNH71At2E38paoNVf/YkGA6DHDxxi5tZqMXrfdn0qM1OY87joeyga
sCGti4izz918NDQdCbylsVzrROwKZfG0NfawHIyGYN5zyJSSpMmdpMFpCcmiGxyfTHX2GX0q7Sa0
+BZxSu2bXSCazkq6vTg3+P+TxBbRUA6rG+3FYBOR8qihk4zOxtQNm70NHgikAxGME824nSPZvkDO
zeOlY+fkNGXqHRfijsiINNsvwBbEmNFIPT6RpS03EPohmQ1s6hPNK/kEGx2lMS7nPYGEZ0tMUixK
cDCqL9IHx1FwpvrYpjzdcHme92sDEYli5tY5Xfi2YY640VKR6G0q8Z6Ghoy5mf5LQmCx2tR7+set
V+QV7J3x9B6qjPnryuIKbR8/XBIgih27LSVp3COYzn5aPHpz9bNmtrRIrZhvGXihnds2e7Fd6t4l
La87MjSnLYnnK09pmgkfc7a3JuManQy4apIcQj/V5M1kcyPjBIewF4C+09K/s8vKI+D03vptRG6t
sWHNtnIF4EoRyAn/uwMnBRHsVHFNwABQ29KspdXvwyyTT2HtaOiOqcVfzebKuKW24gu3MRg7yoh5
Akq0anjzCS3cM9AXcwVD6p0miMZMEdX9Sczm8k4++JzOuXZSuTWgngN/qAhCzJs9oHY/BtI+KFo6
Tr2bfKBckE3af3VrgXqNvZkxPbNFmRto+utp78UZQOaamd3RqRbZx8wWE/pRAaGXy8SrDrjrXUx2
EK4CkNLt2CpCIy8OgAz9VOx6Iq8v7Q1pJ05QQmu0TidC1YVoasdgvzj/9msN8kLfIZ8NHYXhGbYy
oXrAJ9ppcIm/wwvYGVjlyvXEwQlGv15gtEzkywhkgyT9YZZ5EGPjz9rAo0PrV3UYHGuiWdtk8Mdv
SldulAM7hVf1r2weAaBQ5/KbBxfNRco/EHQMLyR59JdM1dUCljNeid/LSvbzm/UUcOvVKH2+Vmhl
iqdogn6MMQBFeOp7svpAE+z8qnvkiwP/q6f7amNf8rP3AJxFG5ZIJdBzNHnkUVUUUfm8soQRWDb5
2iSjXccs426SJ9z7lYBJUmWsaS5bxBAZes85MYOGYlAVHwo75zLEfQYJQG79eSCvR78IR3TdZWiY
sTRjqgt8rmLNdPST03Uh6XQVPHSg3kSRYFa8x5TnHK63G54/kgrXeEV18FnErT55nVVzYsmBU6sW
oE+gI4nXNeT15dFrzPhalxYPcXJsiLx7x/9prOCD5FN0Z8tB+mWDXyZQA2aNuTV9vQSm7doZtmwU
A4dDHvuw72AarczKdVyR6AlfjkQKuNAw5Vrghln/DbwL4kRbpHcS4DFVY7O1lUNOuV8haEZGHgvR
HMcPrjQAtsoX9Y9+L3VuuImFvlTs9Qfn1ZBiQEaqVQgIjZ2QsboFgDzVqpRX38ax7EBU18usA1lw
P0sHHjPoZ25w5vMxj81p+tzm7CsluZBxYVdAiPVMd6OYCeCQwoymCgBevj9jqBm3eK2qmpVGn8N6
JySeSGKH+V9BvwDtL6En23ASetgyZ//JL57ttopBAXYb1Rer++T6Z+LBXyifaFYkX6EZkc2/uCR4
2Ot/ww4MiE8rFt1sEYelahsj5ZzSlBZSdZqfh6PqwqgZAGlV2HJY6D3fHWvCePtUSvzzY5kxfoek
U8FPW/K8lUWATvhaU0FaWrdlBNXmBG3ymibxpjxtgivOHz867hVeMkt+mYMH6vaIbSEdaTwKfAGX
dsD+hR0F6mMnZEbHpFt5BxSsH1Fhsm9wTR0i4dzvrPpF+hP6t2bMi5gnsdJEYpGq6oueBELtTpCw
8UYNwHTPjtm4IjO1CsQxuSIKC19+zbEGMym7Pl5rx/crbu8PDJTQWhJzym1XI2J6ikB1H3HFvV9j
By5EUlXG99D8E6blSegEC4yoMb5+ZKmAkKDOVNfkMqW4lUr42L+Va7KLzwdchJPbXdBY+KQ48x2b
+FaCnWzW69yXyDfLFimmu6ujnaLEVZschwA5uD9ycpUge9Ab5s1D3KWifAUhNwbe1s8LK+1G962Y
bz5XUqutveKIWFDt+0iWbCIcqgoZlAirkZtuSsSXIDvFAuG5r6bopnqJL3AWhwgG65U0rEo7ptJy
woRrqMh29U5DhPwaTx9bfa2YyLfG9BfRoH3J48VMEBCV9Hn0kapb0kdsPGF9n0NZH8Qtu33kC9Wb
yXYwXrb4qxUBgBxlWROu3OwUtlaOAyEiq8XGUKRnLlm3hbw4xq9OKbkgd7V5gQkzK4BqONpaMoRW
+TQYYLeCCb12fhx5X1Uv93HJbhiLPAe+IB3NchGLFg77Hwd7RI7YvxDr3zib/arl3nsCENnsqBYv
HRTqSbEDqZmdssDzEdoLQ2SquYGVhpxdnHf4DQ928TgQvD2tBpfhyYl46zaFywoR4ZAiPWdzpJ0B
/4wSywWIBZBM3SPBqw0WyBFiu+v4Ra3vbbAm7fys9/46krk7I3I9gQPtMCo332aFbR4ogSfw7I+L
9TkhS+VjUvdo7SZK55tzh5hf/T9+LTI4TUZxVK2SrAaVce3CK/a/bQ3uOkkAPFObrL9+IXfb8nQN
N/rHL/KDeUqgT1iw6Bv/zH+CAHHJL+Ahxs7+WKTU9gSS2qs5IVbv9ZPd7TRsBSJcKYu5rG/lByqt
/oRsgbBI/LLCmK4W9a7op8E97Ywh3EKBnvm8uWjCfVv7xwv2wJbSNaLFgw3t90M3RbiL5F+d1iZ4
CxwHZ3e/E3ZPNgjiogWQMLIM0FBh+ryrARwaZecv406zqT7Asp2xIOD9NxrNsp8N3OijNgFePlL3
Or+R48tOhwhiCwXZrvFRcOP+XtYsa7sUmE4fTdJpiz46A/GLytGbgH2ZCiV5876H7D2kf5gYNgTz
8gI6C8tS72w7pbU6h67CURxRxmkwuzc6owojyCvnElrTCyrVbenrFS4elie1fZVj9sT4/ul7rRfJ
7PeqhtZ7i9GpHIf+ZQoyAVkwT+Un3HR4LLSmgRZtUiYwcyutSLPu/VqluDelSTHAcPxqgwCXL/p6
bIYNURjsjHu8qCP8cBxsvUi4KaVgRLTU3tRypUDxC6EAC0D4PUrMVMIs7zhCwOIk9G+0mIfJ5qfG
Q5f61LZ+yiykj9/pauRMmTb2nrzCHwjTBHPA1LMz8KJQ+AwmubAmQxr5qsnGJoiEWZ0vk4keQJdC
fiPX8FkCGvfacjh5A8J9bIds2mM3OA832pUH6k1OxW2M4QTIbUAIduU9f6kLJXKIuHQHz3cEVDiF
MB2JLEJ9FycQS5FC8LFDgGXQyKL9RaXBXSg2oTAdvTvU98E38fNn7EmByi4ajK0KS4KK6SkTKuO6
h4KBiVI0X02ovSYvdZ4X0y1hHY1ZfpmNyKyvNzgKFRE2awXJarENnzLYvZmqafmOVpRJ+vOPhiyF
qGfv4whIITM8iV2ZU1fXg5jJ55W00QB1GzvOkRsQpMiKNw3/PrgCYYifdnCD0Tb3ckjevcPZGUJH
AOximgVgGJJceHmapL84mJf08gvvdbZbabD9Ea0PAVrERe9pvYYeY3ZrUolZT3pmJ+RNU7JBXV+g
oDmcjyX1LwMNBCZQDh0QYCz+BqlK71GxC2NP+NbvcZomhkrv8Hbs2/71ulnon6ry1WsPQvvb6g3r
WNVr0l1FeqLyQMReN2ok++U7y0m2FA7O4L/1dHYwflmqzkx4s4jqkhFAfsr4YIwyPdxH/O3CHEqO
ENprCW92ZwHJ01YmiBhTh2XF43ElseqhYIapZjA0fSiH9aCJD9Wi3F0uiEY1umGnQH/uLMFl27XK
uq6MUozuB+FqJmlLIjU69aGzY0390TQe2hx9OH8XDbcW3sRgemjJTd5bsyVwLQLkGzSQHP7dNcZq
TPovCSM0yDiLi5/JIyt8bEOkpvT+8AwzPxJNWfmYyLMcHadkfiqglTabVtODw0GunNIIVyGfwASy
tVCN5mSOLT5jAp9qSq6OcYy7wYlfAn+LdNhfohQjILobEH3akN/68MeMCqMb4QAV/FUzq9ofOLga
kFM0DHnBYQgHotCKxYwHFxJxLEEEVnH0I6ZZHRPFv3mGbhFh5x+6F3gM7j3+xBzn7NqVaH6MUKNh
SEl0enYvgjaRsoSIX50gs0MAEMEx/gDMXhyPqdblQYaBt/MRKd4OnM9aKNOLKA/BWHFPfZjaSmLq
/+X6Zk5MqZFfIgg8ChcAbo485xR4Jt1ulcnEEyijAsw0PfDNgp4LdesWDDnBDF3LHW40Zo4KBcGI
M9oWY1bWqtTYSR5LRTnJ0Q40v8hzejQmrYt1RRiQOWZpLLhEf3x4319bX0RjUeeT6eFcCJyzah0+
f4Y5BtJBJDHmYODQAuiQhssHJu5j1djcOG3HVIGj9zAcTPpfH3zU/WUuvsRmnhrhF1z9YEbT2uPx
fUtR/P82Kp53mE5AdPFjPRzWGkjw1vIhMGfRcFyzIdqG+68cm0cMrtFI8Zf4ssC8YpUOudmmwX7y
Nv8v2L1vtLJFPyAGUEH1PN284jUz42dnGcTO1/xuqkWw33cYllNuU1surIzt/MlfaiEYPa7BCRlj
w24irI27KDFCYXirIullQ551oVFeTgyxEFEnEnpejTBIhUf4UwOYV6XdWc9uzZTFbP5Vx8lpB9KA
C4B0J4BzTFhHXRtBmFjd7lsLMhbCVSvTqUBZkLu1CXnAVpkRob/RnQHRBeSulUOXo/cudTK8FnQ7
sw51nIlEYQg8BKUaDFgU4XISqdtYdZd3Q1QspVvnbllQMOo3Eb3Aoi9PVIEem5CADKcZ+ulX3Z1C
DsJJTdpZzUbXW2EEhc7bibKzmSlUg3OJwDrplrQ4PwjDSM5aDe8QTLrQ/BtQkdET+5hPnO8cOBx5
EZs8IzzMH7sIiHzfC3pJ2Zmc7LpjJxEEP60Ng5MlwG3K69VSUNA9zzrTNtwuH6MRTCOBs/1nZBrc
ryYRWpBX8c6HGoVzNNGqbisG0y7O+dNp9l9/PoTeheN/Yq99S2vkegyuWLGJ+G6wU4ebMOCFb0om
sJ3rSvBS4syVs7irJ4ojxT+wytIf9omGA8rV
`protect end_protected
