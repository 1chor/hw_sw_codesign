-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
WzLxCVv6RFxqiPCl0I2vKp5nP9wwx0Dq1AK9ZcQ2pxhwBNgRRZkEQt4COJuLYszX
SC0SXBJnPmDX8JEHpvr9GdW6zpDjPSePmZkQJJsTAZ9gmyHCMQQHwllMiBGzf+SZ
HFn86afA+ab63Rqwg6TUm4Me3CqRimC8Ipnk6DmmKLUYH/jdvPmxig==
--pragma protect end_key_block
--pragma protect digest_block
eCQ9CCHWdhDnHucdOF8SW9O1C/E=
--pragma protect end_digest_block
--pragma protect data_block
vkNOoXVDY4LnaJ28D06fIyNZ6R6C5zvSUWvRglMNfWRtaKwv5WMSieNMGQkPipNg
6hXAQqinXMTw1UhAiuiO8sG7/nxH7Q+vUDBPlzmNvyxsfluq68537uYy0/3VW/8U
ktet6poVTse3Zc+X6sCdFDA7xQiUGZqfNmxfvl9VCig5KFNAoCpLDaWa0rzbkBwM
/czSGV85srRF3ehIcfFl+9JmXWT7GpRhK7nVOJABiV/B+DSyp3kCiKIZQqFFIHmn
SO1/3+krdYNWvVKNgRlFbtc1wy1M2DLK39WlinG80kJs6A01HHALNDkU1jgkW+8A
b7E/e8V/zJNB3W+3FQbIPGiHAp5F7kvFSeOw57zZFAmhAMqZ4VFfXbs77ZVr/DQC
LBsRteWBkavsaCz5gvBKGLRCaBhBvg16gDzCCTnxgL5juRWGWJDk+YvfxgngjQzu
flIuqE/oIlzl0qFuwQt5gzIQkUVT6355q5zRNDGGPzNm4AcsGUt2QUBL1fHBd8VO
ZNTAaS7uCIQhiE8dS/JDjhDXpSExdgs0tv1SDzmbl+6z7nrSDQ1mBLgR9T5H81JN
LafxCD55zmKEeRxv8M3VWfgXFLjC0naGaoDXr1SVvsGOEk2nS868ppq7ATYTSHwj
uyrNjSY6qt8XAmlvzH53lJjKUnJ83dhBQ9ynCCB7Qdf7Z9Xw/OtSUGDLOrpAybKp
xMkON/gAo+obfvQ5aO3vDcIzmGBaDQmtxNK5pGd5K0HaNU0oTqxMcM1Caa+stHPG
t2Q0fJnivJr7/n35HzEl46CH4wjoz3BMUZLhz/CFKxU48bylOcAoumEpWeR5dGVU
U4X5r00PdfsINwQZUgU80SRruQ+oDuNHUaCDDRb77q6V9Dupas2xNowBYIxkIlkQ
a8BoonWk0ilVPmXcaVSwh4eda1VSQc/SZv/rg85dsMc/O+DIBYneV5U6HMK7U4i8
a6bygaj1GjthiF8BHeAm5Zfr2DtfviufSpz8L82eOnipDJJeqXBdWEWBHwYVFyfS
igK0K88tgZzG+b0Hj3TfmlKqaXxR41FBqvzWbRd9fvOBTU/OArQz1iKjzMoUhpdD
gGC2bAn1haL5f9oQG9lQw/0scitSvVH5/WPYZGkyuv7ZuhR/7fPFxV1EjJ6ncXD5
dBaNoDq8nB/rQefuIDl3b7++He++I9cHJWb9pJzhZ3d7POVg5q8Ntk8wkIABXMxI
crKH0BFRx+p0uTgZtY2AQ2vLY8RdEeBA9Cj6G92DKOy8aTKQ6hUdOy+wGQxGtF7H
I0VFMf6svsAq3voBd7aT7gk/FySwO0smI9cSTffa99YWHHOH8Ae6+JaXoWJWxAnn
JgPRwV2R4SgjdQIwHSWlu23syHMbb4bVbVT8pZ6cILhDyFjIl2qrUDb5RIddotPp
UV1i30FUU6feb1Y+8kNhCbo9rfOobM79SjCblMJoEPiVHzji4OUzwyVXy3dTfFD9
U38F6iaU7egas674FML7CZWtRz32mAWvOdpPni5GQpPP+xZR/RBe2gpq3RbN8EwE
k1z5yTwpqG0obcxv/mlb7sRIsqxmD4BfepakWb4auOUiDlB02vT5qWDOUPaoJptU
evueGYbEei4hhAtQdthF5puXfJZcT2MWvEGEKhXswLYjmoqnERGH3Dpy08Py+KPX
+SYHpgKStify7chCeg54iaYn9ZlIIbZqqNGU0lbKRUFzTvRVh3JfVMxIATo6QlSW
g7u4gmcgEjk7wW/ph6s+WgM7pj5n3ClzzsZNRj5WT4peMB5kb1R9e1VNqgVv6Vrs
Q0vQA4jXPjfS1PBonDzQ+xSBMLnSGPO5bvmAahb5hASOesStIlwZxkYzOIinW2Wk
JWTSl+fpardhnzcR1AE7f095AtpaJyguhak7DI1Uz1HlUGhnBsIZiOTZJtx6uN99
C6dmacesvYipn56WKpVliPR5BBhwzMWy7meQpXLo4+IUyXPfy6NOMQMbB8mGCmRw
nz5tauchgqAGp3fhGRELnMooZmzdk2kQt5euyDMuCYw62YuNr6Lb1rt8YTtifiSI
e8Q8QtCOiEKfN/s4bCGsnN9WhGGZK0gbutjAamxzRIpveLYf/UagKKrdtbEHTz/U
iITiFRxYfX5qRYCVX8/Vih6tuRljDbd0FbngCtXGYIMv7JPYT8vf3evoRE7qrqzo
2pcRlVWxn1x5slN/ItYeK2KHPkWQNOiiTIUZJPBBMfVGyKrLCCUE7vCgT5ydsAwR
Aa5JMLOzxrf8myL/LEa1sZntsn8JG8XAE9qXECgc1rHXULwWy6eD1Y4cMi0S6AMV
NqBlGLlR8ykJGHUAq3gSiza2i/WCOCtmXbLG3eC+ABG9iEptrItixn2B38wVpxTz
0fZCgDt6PhlcmWnam7bpSfu0LWDqpJucsI2r6DUjeNJL44uPXzY53AOZyitBohd1
yw+S4+jIfs7CVyKSgyE7n0s1Mz6RSutPVV5eOsa9+IBr2ghJCTCbEiRTYHfeFI80
ltuEK3dRr4Ac+ePrL3+eACkqXp6QqPmtkEjvBQ0MaBZxW+uvqFZfgUB8wKXy6Z1R
mlxvBWi0gBgMXR96eow4SKlGkOmoLsXlHQZDuhnaDOL9GH0Q1mmnsY2cI8YSeceE
laNM3hFMGJAwnYyfGQDeO3iN8UIqpPu0UsIhvkpts91941UpumHrD7OHJFGHdmPm
CrVhFoHKcY9HD9brYVyqIjIssCS/x5d4VzuK7qS9py1SmvXPYcdipvkheZchPmYz
gwQtxYFLtTIKsP8xa5jNh44W3TzbxzowcozaetDpWR8O8uQixVXEaORJApYtteCu
Or4KOhBaTG02U25HHYxjGg3GBdq/Oo0c8VTK7MNMJjoV4suPIL7LiciafF6PpeZm
k9jXnXJs7ERpKrarRQA0DBQQG2oWaAMpuWvWbuU4h3EsQfW5YNwyPdvM9QuNxyJF
iRzLGC2v+/8PHN/lXWz5q1Xz55pc8XKamWmka8pOPKD6C7WN1wpLQY+enjbVkhkY
p9TTTRoMD7fPTrEgChw8QSJTbdG3XudZZyyDNEtQawxrd3vSUsE4eW53nGM//2B2
xtaw+5lJNqfc9wFWvtD5ivSm1AjUQHY9ueRwxOhQxw2NbvjSRNqYDAR0bcTk8xd5
PThEoSMMzFVTesdKGuFJEYop0fCuRCD2adCOB4jcIitR4TVHoSHWAMUxVCAZX+CB
xMww9hbxP1yod9O02yxWV4PuHKPDEk2AIIq41W/iD3QTDD9pQMoF1MvBVXjvzcm5
KYKTO5dscIXkXO2FBxR/fus3IAbq58h8noin5lFqVPwAFGDhdhqbj2zzkKHWkoSe
22jlJ8HPE9+NZKkjVDVPdW4YmF5lZvE1/GxQXmq2hgBNgFfB62M6EaUwRjRxw/xb
Y2aEwYXQ7X/PUbggHjLYHvfnetkgMrHt4jKwPW0ObQqKuTMBowwRmW6BE4Uw8ekX
h6iG65bD3hmLtEWo4WyYQkZ3CfJz2pIAzGi3BgtyfVIvgY89n6PF6JimL84qDwch
DFF+NZB8HPM8U7oYVunKhfVyQJgZJkp6LxPoZSmAN/5m8AtFm0HzQoL8IV1WwCKE
eIUZhp8ehtcdQwpLy2qPLYtHaCxmFwilwtovqzPac92fG0UOm9lSlI8ZDZQs/RSB
F0IMIBPDMdGZTU+qI2/9G2CFc142YWVCmgQoMcxK3tDAohN/ETeN0nrb5CuzP5D/
mXNEV+64O5nl5WmFRFRxCoCHR+1VejBuRGUA6x1tVaeA4F1sbfsBnWiWpPGiNJcT
dc70LdNK1zDE3zExr65eeHJc/oIWtc9Tk2P8mwi20NcV7EWl1okHhCNHtchLSFOT
B+CN5vuQIgJu7MSjLm3qxgZJSg+zK387uSNwwWpKEhecXnV27l76FmFbTz7B3Jo3
ukgaX+8HYKPAL9DjBdGoslkZtQnKJosaqtwjRBrSau4FBXQFuJ+/esKR9sj+Zokt
eb/r5d0jENCGFFtFXMdPLv1R2Ih5fTXgErPjY1vE3hLxvmOAari+E7Bb+Go/MLRK
/BEillXnTUDOHfAWJifDqbpsS1htRg+gz4NAhOGcVqgvtnwrBr350ZQ5T2qLHX3V
6VPIrMlsP7aUAZsiLMpFNxe4WHGowduQc3YMGJFlo5kucZtmtDgpAF0S2unwjtTQ
xEx34Me3HioCfIpy2SuMM0Qz9HtSX3VmKpaxBsG04H06yxF2H2wm0+16zk+vsxnx
QsR6X9tCiWR9Uo/pIbhxiON/j57rdL4ZbYGlbe6tl+CAVBmOoR6WPk+gdgbejWyP
32j8HcctuzYLEIDU6RK5/lAfj3JunGVVgwHLnustlaC4gOvEqW1BQNeo0tgLAaM+
CaBSRzq/iOXzFXcvcGPVDFdiKYQ4VV9t+NFIs8e6iiQn7w8g35utTu9t6Xao2vGW
3/VhqImv1Q1YmBGNQCAHaIyDeUCOP7vWuz7XBjhqkF+mPchifDW3e3nsy6RyZ+Ac
hWkeGgZItZmJ8Cor+VcSg3rtBFrIWHqw9jqVaBFdssFtALqTiUvl/RZYGj26cQUc
zp8TofIzU6odiiugelRojhEWTCtQGXiMD33mtV8HkivFripbl9qLLbvHEU4G6rsw
fmDN00ZrmQRYf4sXi7mURcG1e6GJX6YySabytMhP0PzgSX/Flg1oOdsqTvRq9uB1
xMuR1iyHVijmyY3/NnWPDNU5jhA4qFKvcq62WjRa5fevo/V4xQJ8ouA5WYYlFTdF
5/febJ7UoXocSCnw3cHA1LKqoIGeI+i/s/AdTdR5O/uh0XPKgfeDDio/ptTlTRvp
u1nR9sZ62MpSvGMIX7GQeK1F5fpJ4cyblUqP23mIkStjkkjs85QJxzC+j9j3DPGh
cJHdIbLO3mI3kftVzUm9hfn+KKcOl9sl8sq1fTgNm9HvyMQTm0USSuacAriu4yIb
hdled0x3XtcuD5ep0Se93YGLc8Ecp5TBnAhANWbpFHd2+/LTl4KrsxYCEQcLm4/4
JaT70kDJ5OmwVAZ9i7V+G9Om5NudhxP5G4od+SG0B8o7AQkvSmv/SsFOQydiREHA
sJFAlil4O7GG9SAli2ld7iE3BPRZRvIr9zQhwxSNswLaPSIO1LSAQuPfBm37tjZr
kZ8mhYNeUV5kgPsI1qs64MKfrFz9pUwteg68ygGTZNWCmcJFd70P3yljxoyA8NH0
EOpT/BeDgDswj4NZinBBu9Ajqy6brpIXb4MfseaEkDFjPI8tdpkEgqfhOZz3MABu
CbZxhpyX6HzwxVmzUb33RzK5ow3o4THcYnQlHOpGgX9GkcY5MQGD4q2JQvaBUj9S
xSoC9/Y5t6SLp6OsSRC0OWuONFvLNN2Rsv4Fvf7VexRBTa/xyQN17FSaoF3W1TnZ
zZlssZdOjUkm8O9N3JMIaaylXJQXcG7Rt27j7xNjROLs4SHuHTjdAezl8N8Vvttv
AqnUSgVqiOJDXgn6J3vty/ZrWKuk6nc7Kq/udOP+3vXC8hJsySSCxnS/Jo2C10rO
udOj3A/KM+wCtOwj7ZixW8HFcYiPwsHWZT4zxfQTkHLUJm2fr2NyukBmjszOIncI
7d6Ta0zXFA8YCGHS9T86lF2OSfqF+a/NOo/XsO2Uc9+y80vudCr3+MNac4D1/WcJ
BA+SXnRCPconlYGGWGfp4NTF2iUhvBvEPsifZXo0YUymmtaNNlDMrPUGMP4BKlof
NQ5WoE91SpmTGTaQznDSeYf4+9Y4OZgUCikGG8ARQo8dlvhxR03jOeL9u/1HLkzb
EyOhpNfr7H7Y3avPB3ZizFqRj5ysqrndykjZc3CwANJXxV5L4XphCLIiBC3VdgiF
Cmvs8Q5jBYjXA9Cj/ViM0YDqDFaW4lG0y7EjxvGb6+hXaKgxZYAlYb6jmy60/07k
vGeAVhUsLwEL6pOKpZmeb3T130W2sqrs0X9GfCqC0vmv2b3j30rcm8eDYwjVEGcx
exy9im2w1OXhsTtb8SFLLFc+szVfzV2gSZgp/OVmf1XkxwqHZz4ySfo9eQD1nU14
cdoXUJVG+qNChH5e0rZGZ+WU0OBmtKwV16jfoz9uFLNogW/iIUJH9Ws/+5uBF5Mq
p/fKI4AzR9LYg/UWM3kdJVYNZ9BIf3wmr/qOAPu6Moga3zQV+pgOq2RmJq71jsKe
BlUo+4/bi44QbfjMtjBmg93yWa0sgn0qd+e996XfglkKfJI44W/5A1MX0nyOjH/A
BWL6KVtTjrGX/dxXkUfqJJLwS1PJ7B1KQimL/3sYh9JioIQxjXmBXnhCz98AdWQ6
WKK6xSJet9lRioigG/3z1bcvQ3YRpuEpk1tCJoPzxFFmxUJ4JofIS7Z2Ao9MUScS
N4lcGsEP+8fuAb7eOFfbSCDPBHbs/jisTlCnhb6Pu4WWvXeyY3mYSArd/w0u7ckl
6mf38LLd1BVHEBx7q83oLfmSzhqRVsUudpsUUgz46zTeJeUIi4RV9OYY3EirmQrn
2ejT+3mE8RzMpXz6zVapVFXt2RM22uxsB37AMWf0qZzcWY4x3PXD6afpAkK+S6uk
01b/WiclNSQIxHf1Zrt0dinNndAB9zxHK9DxDHEGDJXt4AiqBbAAQYv0s+ot9oGE
SXuFv3KVw9gPYdRa2CZiseSMDhy0Ifv4dGzotCxY+k6jm70gaCZHjq/JU3kI4Zlh
LIfI0C/ud7MGC0obLWsjxsgc9ksc3/gG+JbhJ89XNiVEH7GipI/MDV2YRQkUGi23
CCHfM1/eouf7NO9GAHscStxEnNdvL5YX5mZgTeDfTcB7CY23W0Gy2yMfXXtU4/LU
EU+Gpd/VTpRrj5S91XTbUXBw+Qo/E88SU4K+jfKqjKzPQInOl/kFokOUGhcj7saC
LsjhBkBtAINg/c/U8Z/mwSWZMHKF5EH9jJPGLAp93+lu5Vn4EiqLLTmzEFAzzJCu
8nchEqfA+dMPAHSuEha1c7ABQQINP/an+VqU0d0fkaPPR7PNydiIwp5RvhtifdVL
EQgMIwAb+GFIquBAexq9PuR0614+Qx9nFncI+ngaiSy2OmqK5XSojF4r3lh5EQXi
Png5pw0IxSMK6PcMI1aXo4Hv5BZk+QZbonxadpbpVt/cuSuF/CrJyZMrTN1FsCWI
U9OjdOVN7gsi+arO7ASrd88x0iZcPNHV1JKQEBgMWnQDBO3ccWNwJ4AWCce3xKx9
To0GD6glSH11OKW1mrhkF6xwpxAoOyBsCkAPmNN/J3mnWAzRsFCi+0ZJs3yROFWK
C/crymGv/K/tra2Z1SlcXeT5LDaSRs61ND0mvxNMt/O03eWseKACg3hNacHVQMhI
5x9AgeJ+NFF4ceiORq/MkZ/a7ru7s/QvpsmejFTl6Zh1PXlH/hvBY+e0xUTFL5st
EbVXuvytBZrAnmIqqV33HpusovlzNE5hmT8q8XicaCHabOER/Jf59yjoZtrTXvvK
bPslIVafCuYs77XsxsQ7tzJUKKmW9sfduFsZgvCnFRFztCgvI04tnaxm7U9ImCGo
Rb0I8IidWvfWFtHQunIbQpmrHSzoKsq7UAUl4RyQsHXhI4qKDixGJ0SsTU1vmWH0
asPBukT+xcNeUXW+mVeM8m8ExQEIFWAUJGApAjmFyK/+Q2cCAATPQAIXCv34fvdF
R2ZtYXTlYRpOPVuhoj8Zgu+IY7XJtDmF/EDOpD1C8gNteaqpSk/lMUQ+mZx8ika1
Z1CFcYsF/BC1s4eQ9UhAxmJc9UuT+rsQnjg0Wrgp+HciMJAGgG77SHKRYmfmabsg
ongbhE4EuzNSYAk4gmk6atkvgVNtneOVN2OV9R9wLeczxx86J47YncGoOIGb0qAp
4tiLXY/vG4KU8tLPDMHtXsUnGrtd0VeUjLFS+//gYkeBCMhHx/1lHvoyhcyDe1sl
t3PMYYOaSho39DLesv9SAj4NOQgH4tFg8k74EbFjn9CkWtNa1V7p8c6PJPpt0vfp
aC3DWfe9LaiXPy+DogLuJEzVwWqIXStbkotMnPz0Zw9jKiHvyLFERr2g+4Kr1l8r
Mw6kRlqYG5vq0MtIByl3PbqnF+M/RilkVzNe6ux6Z3rOTfX9SA+g1W9V0VzbX/wt
YfI1iq4wUAYPPc/A/4WCsmAAf6z9SNMsJ9LBy8ufiEeCnTogEyYQ43UM/FiGyN9B
JfZ4SukiRD+WvzfNxomk7ZDjrpnikn+Z4YzWM/9zoA9uhmx5bEeIMK/fTEOGp7O+
R5uDhB1SOa1ZVhb6FuFoeGznBneM8XuFAmp6cu4TNWkeDlS1FxkhhqGuxPD905PW
UQIjD92r2RpSxOv/+P+Bx1aoD7Soc11CnKJ0FWkQEGixW9MpV57n1WxP2XjVz2qu
/IscJUixeOoOGKU1FhW2vZr7GzkoePRrkfOJfuIFAK1SF7gwFiLkY/0Xpq2kYJ2/
clrGRTnDF/rQw0hmYu+XdbhFspZ1GLJWCqEaAKUh/z/Yv8wl5kh9+7ykarwTiGrq
QNgKtPzshgAJlrxqc1DctIpcyRc/dqjcyCSWcULiI0k6Rixo+sLiEjMlOiKRX7UD
EKghhXHesOZyLn0oIMF8iN1JpCz3e8hktmCFAuXUvwPOwK98udNYNOCR9IsboOKg
SaTIlYTPPFHyhaaMnkluPii653PLeAocyyShBtW5eRoxjkRQzIZ1K9g1FbAB8Hc2
NeHhYqgFhph36c2jIfPMa9odydOOrTwSLKttPPAYecixBuxK6lTuBlJqaEBrbyg3
8UJ6MpuQjxuw0112zbPdneQrLRPgULWQiTmyS7+hb9UMr3t/RVKrJgDPD7D+e9wn
0q+R1z5QF5WGqPHswFye8zxlRG0NO4DldJt2I9FPY82X5uzB46sTxqgRdaGXJSt/
lOAXwP2a7gDCD68inp2k2g+D3ErDTavt3a6ZEBQ1ZwgwS5u0OgR+nc+eZbiBraJV
HIoU15dEItJHIm13SV6auVwbbyuocXLyNfeuhv6b5w1gHUmxa0YeMBe+xvgzQjOx
O5u/zpzoWjkl+Hs/uoDOL1zdj0odzQ0uJy87R9zayTwkRJErkIiQgYScKANAZw9U
y4JMQPLv5H17FlmlV7Bc7vVJIj6SWtDj5+XnhslX7WvfcwGTjFYE49shbgaSavTv
M+nu0M49tj/NyHh7Pen3H/FP86rQc1OBrHW9W3CEA0pGjhpJA8NmCaytYSstrXlu
3r5kxtAUerH0u2gsi8dPAXQtHmIlDg7RMmWnGwnSpZdBd+tAIOMi9Ek3ti45mtWV
W1zfE6lG3WKVSywz+udMIck0DTY5Nv59JmvM/miOrNl44SRgqR2iHVuiWAhUFQLL
XA/NpeFXdnOGtOo+LgFkFlPEqER+rDflkOtN7WJoygK0fmZt3JD3utA0AVZhzOKo
DI6qqKVvChCppiTU1BO0KSzzRGzKIJzfSBozxJ+rl8PRxabreALfXIBqhabZZtvL
yhQqivKBFooR0Ta8LM0sjPoIo3vew4zDGqaJh+PnVHzt/dYhiH+soTnE9Y+ZQflp
R3GspZ1+3VvUtsZ3KdMCIbDHPhcJY19lyac5sdwZdhsFRkAgNz3WwqbiO4rQ8AsJ
QGz4f5d+VCIJr97q20t4rP3U+BPmjAH3WwyB+4nTsbbm4Kr7tl6awHLhwawxIBgw
yYV//PC0VNS3jvQpfX+5cGKRfNciilHq9XybUbaOkSc91GgZ91TLIkhA4EXymD7R
z3Z2sP2pWL7rGgBj92G5M76M4kqW7EOu4PmWshcndNj235UXeX6gW1ApQnaKewl1
oUBv9tHzx1igujnb/TPGOhjNG0tssIQHUKtEvlN3k1AL04Vuu3JVNNb3/pEP6MRJ
p4DGR/u1MVtpNbhGXh6ept9wll+pqLKid7HDNWYnp23Rb+4DTjGQJ6P//WZ8ftPK
9Qh1eiJXe+FJxsjvrehvy5aOG7TQ6jnJuFiJKsRwoReGUoIYNWbop0DKyErkBzq7
ToU5mrdmuIWdShVE3BTdWJlKAJeu+WfD9CI93teUpRZtYiD+agNWpxCzlfPzBtlr
CPgmAJYERS4QiWtCoQ/R5QN9ykIkldK/hqcTFn635K7Tpm9rsqRuUoMXu96bqE7C
3hfCGaqPsxr4hn3I9F+Dp0QO0Z5/FCZs1L3dg766wgn1fT5ijGR5t7GBheao5A1d
bSv2KOcsricQP4O3GRR7M+NgKySKcYSzY8m5m74OqF5b6TFwpN/DldH1ayEsyIby
dEiLayNhwLUAKSp/HvikiFYS28PzmzMvsGXPfEWKu3Abdvrcw8AoqJuDlbug8aiO
ze7WRBsSgv77iX3JV+Be9DcT68O/leEbUrOdYxD/qJNRYvZRRQfqMn8ixpk5f6HW
aMQhB2f5W2Xz2A7Pol1UxhPg4pJ1eDpjke99B3y1ykRMXh5mCXOMj4L42xm7iXhv
pJ+XuC09uQuQKD4uxj7bc932xwd9nCeOLjVuierrGf9Pn82egHc7mYriaIi5cfBD
ZbO1D380Wc6gaJynQJReP0g0yiDlZyc01PJOGSoT30QJIGVFQgKS+UhKNEI2eQgf
41ELoEMtOv4JNLX0K55toAx58baXy0WJg78cB7AaF2iRBKqaH6PYSQ6Jkwt4KybB
vI4bMriRg/NHskUMQiWlKeguXKyYIqN34Dp1VwVTGI0nelDHDXCpHuj0x10ZFQID
nltyCcGnPgo7Xagxt5fxOWL4Gpa0tsuWqvuW2AMZy7mfVuJ66X5hCnHYctU40FB2
dsohM6LE5LFoaItilQid05HbttNjbVwT103XF2DWEIAUVfAeE2jIr5MfUw59aoWf
gQ5bpR/5fH8dGpBhBEne9AccdULEJ1D4Y4bk/ahoeuUt20ZLlXhJLsmVNPcm2qm9
FoClBxAl5lZ1SOoPu7XJyByJQahm2O4fKgDY+HoUvVlZ7lhtDHnvoOCyMeNl7y4k
Vavns38wRx7tGQS5Qsuozyqzo/Xrp0yPfPlg2//eU3Buxep5jkXOv3e14vU0J+NT
eIYlmud7Mavv79O0e6e6in+115L8uOS39FAIW7MQ/ZAz32h151iloXEO2lZvLvPg
Nzami88W6AYAW9eakuY7dcsGwMIg701zf0CsaQx7nnJRQdc1iC9ZHayUVCRpDyHg
gODyN8wzTjff6Psimdo10DSiOWeoka2gW1xqliZF197FV4ie6YLv1AfHYea6tJ9x
sT590JTUhjwGvpQMIdVmYszE3cm1MrjxkeM/8VEHUSYuF8lKHnf24uKWe8OW+GJi
fYVRfgB2wcqZ79r80eNokV5X28IK55Bz42L7SnjeUs5BeDV85eMaW9n+6QxVH2Lz
oaXFj0eZiIAdOO2FC3hKsxlslUOtVhg2tOEHs86RNSKu9QVGs0iaFbXZo+kbd6iI
Ro+ZYMdSfMjjLOtN/fNIcAvur7ioVaHZXMGHSYZGGGgkK/5NSYH5UKSAUfVxlkls
8qLdpRBT+twST0wIWZyY9XHEIomFEn2qGuhAAKbuy2zfcdylCmjs24ouwCQ1vfRJ
dt90Mf9QCZiuhp4mLJNYt6D309UwlWVO1218OoGxBIcQLig0y6xg9M2d7joVa0eG
UmdrUzWUx9zhZV4M1L19T4Kr+4J6VK9h3MdZJzo4OWV48ylvOJiwo7P2gA1WlgXW
FLenQy/WF6SabyG76D6Cc0BvstTb3TRBeZjf8xsxaViALvSffYvGTlptd68p640m
D165o8hcpCjld3Hnxyv/feMwGoOuuw+gO7Ndq0IdBePhSWhVEMNXic4dwpmTPIIk
pXrg2L/QmAnjorhVpmEHkGSSAf2xKThyXfGEAylX011OmPIhfSy4wm6VxEfK595B
Cmf/ubgZxCWyY3Yre0RMVaEf/AzJ1ntV9+12vAcI8YntkctPprkxtgkKEDT35IEg
XUwP6QtFGV99bSaI2iIwbxerpXvmx49LiT5WS0rR6r70uZ+H51c8xUygmOV2gT68
GCf6YLFbNgYMUm4PgJXcT85BHi1oDUg7tP5Icba3VD3r7hyJf3C3b13hV7Za0xjP
vENA9/Vgv3k451hn6m9sXSHClQlMc0v5LacoZ0nho206yVtVxQfel2lLK+4xLU3D
WT+v0eBafNpZzptu7Wvs+KogxCU1Jqxr9gmgSaUggxDNwvcr1wygtUZyW7AskFgK
URirH10AZRB+JT7ZEUS0VZsDyPPKP0uMYxaAhSLKVMwjx9nttY6vpA2zuYc8dAaZ
HfuLrt32S7C808YlbU/PFrtSglIXjSzQQ6pEtkSOWo25V/qZ77qGQwfrmmDl1M7p
qmVVG0VrdwpY4Edy3z9whiSmcr7FwDvJ5aUYEEGsj9oBpQ7jRpMh5eJPGOCIotFw
BdADu+F8487UODUX4lbuie6IRw8UxMQ45HXgy822m3M2tydk6+OYYZolKvJKmABK
XXEyTBjyL1X3II9R770Vs580sLziNka4PJgBv8ULO1qJmypX3OaZxJ0GWoFrui2C
/oj6+N+Y8vLB/UF76fZ+XkCIaf2XkHeao2Ej+s7onibudgzTNld+3LDqarTAd+nf
7niM0eNX+SszWg68mFpvHg+StpbJRgOGZChGPQu4fH/NPTN7MYGtU3WNkrbB0ZwA
mR0d+b/UYBOzCySTRr2JeV8ZwV8gh7wpYjsBHLAnhu+Om2NMuOV9VUqn5qnkt0cQ
ielhs0J2RLQpOACM8yUJvB8kaaaghQ9SSwYNjzjzxygz3TL5i/QMLzcQvs+cMtEk
o7Ngrn9DqmmW6f4wYgkOUq2MR5uiS3mJoW43PXlJboIxK7PgJVIx9kOgHrMMjESQ
BENWKv4AHTGQ/SjrgXayAwEU3dWe7uIYNatEArjjr+AtZzayHjTuD9nsoJzGCUYf
plotKzWULeBthYX0e+fcba7qR4r22B6ili04a8npJR3iTfoIZrL7p5qo/vF5Ksdx
DwfvAWGW5n3G/cbuQiGI3E9DELOwps58+d0KsoZA1Ll5P5YA07+M3rSt4xEqym3I
fYpt5avsec6tP9Yp/cUAxePfMaiqu6zxZK3RRkmd/5C8tgPUaSRXSX4Ft3vhLvw5
Om+zD7M+gjsavGkGjzibl+33rUaNjmEDtpa/LudEZ/LSq5UpZJcpeb5ehhC8iKbS
52+IYxmv9+HOr9/kOLEKAia95JcDxLIxEqG3ukBURMhHGj1fvnKtyJz7u1AHyzZ/
mBdJMKweOG0RoC8BnjBh0+m3dhZLdAEiiji19g9zynFXvvDWVtaFM5S/Vd6Nqtmm
K5OBrzsEBr/BjIiHEd0FtTnl4m1F/zq5AueACszfqOccvHJqd7YuubV4+OuwaPHb
HiDu1U/T/c2VLn2Gqhp3U0Dj65XkB4voF/sgyfESW6c0HtaK6FiX/1ejMJRi6g95
WlITmZQgK3nIihj4iWZrnPGh9lATlq/+nMcDeAnhX5yYQZdzBnoGcOv7BxW88lbw
wi+sQr2FEcuA9GDbCNftt5LX60TjPkBCamdu600JTPz8m2PrfwAu4/VubL9mtktv
7EjUVtApsVpj5rLRTzv/HLp70fQuVqBHwO/n4DfWhZw42kMiicn7ISmV//sGXuQz
YBzC9aWOn5YuyWIB6fmQBCl8FnvNWSJVKgy6JI0kiixAgzY6obZZzCkBLx0DzVsO
5Bw0vkhNxOr7NIcEry/FiwvDNLIQ02bjSoPOF+ywBhibo8ehCA97/ue1G2jnpBVJ
CicUcpObmOVHnMta1T776xNhdjgCrogUG1Z6aim6zDCbZ763cYtSgsmPO6MUFffs
ClcfReWDDP5dAsOy2sOUnMdW1ac1dxJQzWXL1SgvlFMxvz4kmhCU+InbeMw9CbjO
QTTxOjW8M36TvsZ03cAN/IWT+uXhoMnTen2bNtLtTD18ldwgay2qnR7JRgTgzJmT
nSNozdVxUGiEU0vI6xRgRXnvnE7IY1gPT79zoWpay3VEBLqdhWcRcY4B1hmPd8aK
EAvruv+6PSvVT/NH7ycc3F1nriNhzdQ9YtSWV33zkesJk0D6TtNexzC+rm0ezU10
lhFEXAXMfI1BwT9F5XP9uVKLNfH1ptpuoIEim9GE3L6I5SiUsbRyBBkD2y0R01RR
ofqF/g/BWg0O7egXLf0FUx6QKA1hovyjTlrnB1kDgvllBg453M/5f37mroTKJS6H

--pragma protect end_data_block
--pragma protect digest_block
T3VrALXh6GNZ1pYkF/F8taj03Gk=
--pragma protect end_digest_block
--pragma protect end_protected
