-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
FtbOhCi5jRJtipk2qwtzrGmBEqu96BRT53Y/aU7Gun3TJ8r0P5cC3Hp1fTBOW6dN
dM9YmgNx5oAhGcXzi3+cVZJNY6XQAeldFK6stL3rtJxxS557p44YuFTi3q/MxVfc
rz0kvw+2V++Qj/7OgFfIPLku+QCNKv61Anmly6+30uA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 20784)
`protect data_block
4rOa9X5zWLLND7KNG5ySYVbCuX1Gz6b5DQxVMhLeiJqWmAxkXZ8iSn1WjUlpMlLK
STi3vWStoGqk98urxcwez0If//VJcT62xgufr25z+QLLfx/Z+zHfeik+YKd7KW2D
617lAK5tqiG3eNXqvcPriE9MJbgJzHAao6wIK8iOpC6aPend5ix86gH9t/zVjugW
i1TF1GRIAEiAj1tubFadLA4ojc7Rg7SNyrSsUNxy1HxZ9iP8Z4KVH8gG7hcwaDvi
9aCYMIBK6E5aoU1KgquQvkMg11TU3N4mod6TNtTYVjrhWNlwQvlhYrEXOJVb6yOT
aM+tYaTKvxnDoNXiP6AySt1nGhpVUw3dD3SqK8cYMA+m5Ot7x0KvoYuXKummQsXv
qvQaLsyMlh0bVdXqHCz0c+RH4WSoYKyEe+OgISxzewT0zQ+G4FsHU4Es3WIc3M6u
7GjjZDirye5We8j2Be/8prNEMG627ChNf2XgByM8Dp/W3UwDU6vbVRLAGNImZoSj
1Lqud/ppgUOzqLMqEZFC5QJ7TTcVpLLAVT1vlNR9l0glUgUitjRaP9uKGOyHEsUG
TNOFnqtlxnRmZTmYo5qozfI/3mBonGyh3+mm0NCV/ibV4TbCdPJi28yHEY93SHl7
5n/bLLgo69LcW/RuTIv/vYSuKTyxaYILBE2fjhIEgBjmTwXMHnLF47ZFJk45Jo6O
Y0yioocw67Osp+6BnPE8toA6LMtqjn0zDxTJ3RzSwfL2PBSpAq58W2HrnmuOoloT
aWRJPghn0F05tDehr1xmoN9BmuExkyok2swzEfXklPUKJJzm2SCKTxg2D5sH0b+u
dkaeKuJThWCDRzm+PortXbVTRFBVkIBM821hhSxtli9e4QIO7VCWdrpKET2NZjXv
H+W4dmeaGB0AzcM6wW6eqU4Ask8gptQn4UraszeV/pFZFfM+1+OuzX1Bvy/YL/MU
/l0DPegooC3GvB6YGuWBNSjvXk3GVgw5X+F+SndZiUFolu088z6yINYtp9KAduTr
p6kdCDlXo/ryNYUubiXmRDwnbKUzc6a1mXfTSGU8mGiwf1MZ4j2lJA6KAX2BNz1L
t4TLA7EaDogiuy3MUokvs5P3w99TVGMoyhw4AsDa1hzjZATiCi/Xb3PZVJeWC0wG
WXjYl0UCVtr1YizFLCnFiL2SB+FuoR0iAf/u+OODHGvlkTB/Yds0RtSK1wIL0o3/
wvdeGLkxJrgk3SosoVvrXBaVoJsdY4+JMKtpqgK15x7ZCFYtf+5BBxWm/pKtkIyy
sS9KdZA0oKKJq6zua3rEcZxJWvo3ltjBLyZpNzpC2cQdrD7tGbI62Bexl3s0c+1+
lkUo1sKEgSNCbrKYzks2s2wFhH6NtiFbIW5sbHg4PHoj+aFzJj5FVSHOI2qGBZso
Jq4HGxlA6Ok6SNhf/hCum5OalIT+9vJ06ZC+l2eRAt+L/7MA5ZC6ZE73rSIYajLf
fe7iITVVxLrNIa7at4/35KDIW/Tyg49tcmDgzOZWQNe63rTMIMBi1OzfJZzpmn4p
HKL5eHu1PQMOGlMb18SsoDIQnrbni44x0iy3LykdI62vbPmTpSIj9Fqm+0GqvmFX
DDwzUI0rZEktwhtleU/gimycemN8vaR0qyAnA3I3GtYFtWSKXyjKBDRVcFOJpijl
2CKHOlifqmFw0p33O73X02WAbXd69SCIrJvE03gaOHJupVEbAZ9wxozluaLH5hPj
bpKozSiQ2jnQAlefLofY6NlnbdRfEvqhcK4maxNtkNEc6kJc/fg+a+YLEvL4C5Bx
z7VFitWy51mMqoEN+5SjCzcuvtf1Omh45e/U0swjEwoh8Q7NS2JxRvdnraQ3KWM2
i0hr5UtsL2l2/k9rD63BVuBWMDEStKz7K0PDqHwsocZGX+SgMJp56OfT2ZCmAHsE
89qD6TqMGJZRFU+5fpsrvej/Utp+9Miq79ko2RxrlzVNbO2Rih2clyb5IDQpsyXL
nrJlh5RLO4WE8NYQURVyck54plRV5qzfAnfXdMq4ZUj/5l+e3U+ilpAG9okpg9QF
UVg+h5f0u9PtmE5SR/EV+aZtA/o8Vw4nhwXCjKUIrU9t6Y2YwDwaWTRbFWg4WtnG
+xmIkbFod8quT/giD8b6inBnnR83JRoTkRfu/0DWq/lFOmVA5XQ7zCo8tBWUsSLE
VxKElx2TYZTZNGlDn/xbNOqr7U4gOexjBcifPMVniZKIXqRM5zffqbBA/V6r7QlM
JDUDZNSJg6g9t91WXTCvx7hUeWFRdkvCckWGp8IepWtVunAQNLmSR0qUT6/7uEiY
aC5HGa0C9e+ffNaBotWp6jvqByeUbEyv5l9ntrlPFZHjMhSJ01n0ZxRNU7H8QF7P
KPSgzI896sDS4fMXoSUHHB0rJnLw/aIPLVtu/gGMVjMUA4LzwFRC8tbXZotCjF/T
l607Z7ZTtLrcjbFxKfBbwt2Uja+RFy4Azcgz09SmBC3kc6SMN0TtKyvjViclTmbp
zFvIVZ1IXfy9qd8IH1m57Rsas4kztlM2jQOuBRK+wnRx77T1JSIKJEd9R5Ou3Mph
GbyhLhx113LBb7iFutED08SjsbViyJFxjROkCseOEAuLJ/ZP+f27Y/uXZqzbqyD3
YKxioirJ551SdnEUQjIsf2NQqopbpEvCt/ywY/f6RK+I0xHQCxVyZcvJJ1KdC2bX
jjBM08kiSMSGnOp8mV4PHP25l00smY8241NXAfrtRNKxTMvHV3zf11mmhCFJBQSg
SMEplA8fcfSBNPjXuKoTytWa4WfwdqL49XAAdUY5yyKgl3L1L4L+trIRDNVfc12+
4SLKFy8+x2Q6EUcSGNJHvBVgcBpyo6nJrR6v2tOxmBVKrtmtzsIPWuaXR1ckFZ90
4eBrV5dtUY8ihXgh8loq6/Q73zVZ2xH4L7zcy67nmyfmlhXJCW3wvg63RW0t16Mz
VUm/VF83C9lbZQBpBK3VZiK7a1FNbDgzJ0SC+M4D7MvIaVgQTbpSaou6wyBNz9dK
Tgotp9smpgFQoXdCgMl3YUdmhZnuTPELZZzXK9aPI/OeYz9Exm/bFDa6T4MDZNVf
z3CMA92ZqGByiRFZosxTuhcIiUyD+4IKRHXBIeSm9JpDZCTAuUU1tMjZoyNxS0ss
Vm2I+acahxV/Xg54ayaxUyStcG9ih2WiEKTjVn/OlyMA3hqKgr95DBoa5XG/tAFk
7BFc1JOt5fGyHfzaaOecdljzmlsiA8cCrDK+rDSTsR71chuL3oRjo0k1laeJDehP
FxjrglN8V5lv78MY04CNJ8+YNTSjrXcHWLBAJLo1uXbSMzux0HCN3QULMy6r6MUv
MpvnpuewXzmDZ3UWmN+8d58jw3e3+vJKRjysw4uDWthNaMGvIGZIU/76L9grwkzP
bhM0YuplWr/dyrhKH6i/ABb7+6/CpPNBjNB8mjntH8ijL/G7R5FZAWHpH2OuYs19
xeA+gJDRD92nAykXkLaP+32jhu40c2CtlG2Leey+FQxt0ux5DcPjBpIlhMDDYlJK
MhANazD3LWZXDDi8KcZrYMNJ5BeiyeIZ7eRBqb5PWUbTcD5wEz/9eAfOdANwB+Nc
1TTlGqTX3JvMP65hDypHWTAbUhML39MUPBpn+3JD2dKADRVqxDR0J8lSUB/hpINI
2MH9BDAF1MJmf18i6V2Sdw1RzhdXuhPUBDrV/TXolLvvhvy+CtaEFgknINEShiI6
pAH++SPxH0fm/o2GMWqtdUY3Lb/I8riselNISrOerIPjlXX312w/Ri3pnbzrLktG
tASFweE5+6keNVR9Q5aWO074oxoWrGEz/Cfp7/r3mS5U0fPpUdTruNcITby2kNf9
HBhb4uQrbqEaooyBZzl10YyNDoL3X2rRIX2vR+mvv7UjDd9JDUfR+3pSzt8Yvbwr
eaPq+8CFGSfqHyg8A/usDq+Rrov6eQKZ0/4UlzOm9SBwjRC2OZQKmZ+Y916asEyq
lspgNdzf0TTmotoqo4rzPL5/HDqNvjkKZPvq5vMNtyS96FSe5GMT9IgKOuIzXpps
UWM6gqEW7zp0jWsWtOV5CZOkEwxGJz+BBhn6M1gGja5p8jnpnArYy7eBoWrRyz1T
ACLyJFPKyT59s4eKiL86xG+N4Z3fY/rpGXnYOSc9gsvu1ou0Ex8h8/4VQ1kkI2l0
01t3hdoT6ziQq0RIye3ffsYfIMmC/7m9H08mV1b45da17ZhDvoOPm/oBEs9wx9pZ
JbnhsCvkrZYJu0fb7yDHr8bqsFw7Xxs+oOCRG67iUwMVhBpKFq1tpwWswFv3d3wx
tkSdl9NXlVe7DlJO/IgL6ipTYV+xZzy0OenJq1ZtYRn+eRaKdpIDk53Af9/IM7Sv
6t44wPXcb0wyEgdCE5eMQ59cBVLE7LHbwHWUMN08h4ffyQP1uOiCK2a0ylWD5b7K
BvPK0YISQdKjkWnJ/nTAw/qb4MH01NSKiw+Ow6i1HEcdxLjlEXc5IywYgurA4yap
aRAN09W5tXGsHV4ufe272wI+KGXfgBTaEn9RPQxaViju+jFPO6fA/INC8XJ6Vp2t
PSLvdTP05Hk5NSlyOerfOs5gp5O5sYJAOsDkqA9Q5YxNv/leuo6tkBMIQboS6aXw
D8PPG0Eg0kd3tkXguxLrS5iqqElIphIAmuCf81BZO7aASd8eSvfMxxDXLHBcaDDi
xW528mLcNm0KzNwbjQPjG3dzl5BXtcWYrm66fM9qHY9Measp2jSGieMLWwIavOCA
3mN1tO+9aMsY8zujZUPqWABYC4tY9Pthq+yOuAeWFp5lmKh3bZDhvv2WVfiXkRd9
+hoD1Avfe0TNGnfFEQDQkT8ZjEe69pUIVyZFfV4JWRkv/YZnRF7qdGL19d6FB/7u
H0ajJ83/gdK1i8tiRNB0sMkvojQWz5B91ezOdkRPSffRojtH3BvK46j2UwLXuRfC
dS/WhGrtfv12aHWSbkidXI1ONj+o02yxgszDZfr5UuYjhNV1jgPX2DvUXQF+Oidb
Lm7GWYGcbk1HVCK1J+uj8n0jZRmQMS2aRQMnh3FoULRqiaqoxigrdpFgu6tPI4NR
49huSVnbYj6zDrSO8uThSpFGnnFMXOCTkmOxu1Xsp/UcNW5i2CdYgigLXS8esUWj
919E+ILAI3D9H6Hi40RoUlP9UMFgLxf3PTmXpcPl0/O2a7J5MyvAfpeI8qP+GQYW
aLDCAH0806bGqFS9ITDvv35eSqRb8VwJYEqM9mxouQ9IiupZqo2AyiBGTSkYMZlD
m6riHQYDWASGeocP9Qxq1nik4Gfvykxfngvth9HgutcObYECHHv2w3psn24GwoEB
fbfgZgdXibZzMkLnnRpEHBKrJnxDc0fDIgNhMa5XET9AmVmMyOBIJjETHdXKvi86
Qq9yJ3FNtorV81ssRg/pbBPocUvNwvV1ZyQNIuXFB5BATTt5iq2OX6eBdHnnzjmM
ZbCDg12dt1TAB4KEnoXFncnvS3NJbVetWGB5TSwVYPfLZmoHPm6fCaF4PIM0U2Cb
8pHHDUPhEsQOM595+HKhXjrlscJb29X45GNuHUC15NvYqQeqCB7eF9p1gctyYYnq
wpctFLKlnNAaEhiKKgyVwcxd1seawHAcqflyu8WVIFkRl53bCJrvJ4yNer6JjOI2
YP+6UFUL+s/WX7ClifSiZzTcRTtuWV8gWwJU5XbIrDwjsTlNvqaU4QZS3N/8VEnZ
GlQqpuLGA/sRMINU/x7Guk5C4EFp7FQkB7vAWWRhBUiysNEuudKUfIE6Nh1qmrC4
N2QeBV2NZ+h8bs+8VKme/+1QNW16mHOWsG4d9vst/kPNF9QMM38o97y2kQC7wLOn
hY8QoWUPb3wgVu2Tie46Pvag9MnBNr1bBhMeVR0wgidPMCl9CG92SN46skBq1VGj
3nl/TnJOK2iSHN2Ufi79Z64TXn8QxLa9T83vxl3dCYNCvzvYuZD5mQR8oLkeZdpB
0lHnB8pmr0biAxcxKViDX1Ym/Rfa4KUHtD9PvW9xg1NnuwQc6AIkeB1tzMTQ1ZeR
i6QQeAxegn6WAkuUYzrT99CchXfuAce5fy1Qb0x2OmhSqlN6dHEqpqdSuMPXXN//
ps8ovOetHKejBqmbgeSIGbZp7j6wUcIkAWv7vwOZyzwwbN72V9N8LmeTdbxkKAI6
8pMnFGfN9wqMnU3hOPb3Nnj+FggJmCe/DWniRn+716w8BmWyxyZnPYlJaZf86k87
NtWSMdNsazbiVghguJPTLz8gyWTV6rojUnrwsF7M24lnJ5W62QMMVvejKMUwfYX4
cmvnXteshyAiX30/A/zDI4A8SCr7sv0qU7FtblsZCVhwTUYwItP/qRcZMDBhOSWZ
pPqnjs24ta+uIxHfza7roK7N0+LC8hAc/G5G2E70wV4Nnq+cWYZKPrOD7oSNlufE
syj2t75ULrOdg45y9hX8riVuo3dJ1IV7ObRVCK8PbnTjMPzap3idCFneHfvDklIz
WDQoku2KIC7p9ILkES7E5huYgDCJrfE92dCWfiwrocJb5bZMVGIVMDr53gWxWtM7
JacuSdIQiB2qMbXZyqTDIXEBNaFLeevO4Nj0RTqsLRhI8+5vYmv+5z5SN6m25E8m
tNaTZMkYujUgbtbZEuoVbMaBeE9XaXXvCYNOelSAEtyclgKbi5X6mMHkVOP+IENf
MxoyFrvQPazsfIPAyFryIy7uGw58kVNADBzwz0f4MB5g7XMvxvzmUVhQyf8JNzqr
pZPAjX3QBjQkenQ9mE/ArGi0fQFAjd18j2Ea8U06rvp5QvonQtNOCFKPIromJ2Hf
EeQGEywgwx73L7br5G6+ylWC1lfl5sieXugeb7lyZHOf3cwnzJO9drAMhuVzUIpI
cvwpStnjSOT7RilM3hbnUQUNp1VbPBF2/IKrKPcX+tAJBzhYwQqalFg2cCB7a+G/
KXyIltQg12uO6BjE4TB2SyCf3rfN9My1AwBAKCilz/jG2XOH6ebDD/AjCuISiKAK
W95n6c+dt9H2fIP97xrjC/Voczz5lHX1jSnO1JCGXRswDbycadZxxID5J2kESMQY
03KgV0Kyxk60jyx0ZK0yvPZwK6wnDAwQXRawy90a/pM0L02LMxq2xgKZzGwWnw8O
psS0LD9woG4xmd7KGNUB+tQ05xQRE4Ad0wxw7fSXFjXnip32tHG/5/DgW0P4KqAr
KsGREqFHr3lzVcHwj/R9cJXzIfcBJ9c8P7+9lXnbk3DJEggLUbp2mRG029cYUyRn
FpoBcA0ebfy90wHLUxLT837t9N6GOGX7o+cTt6685epSH3fVzjyt9/DMQlvS4Fk+
vBYrnmSC4qGrWT1qjU3pStUjGQtEwNz36uTkbEOTqJAnE8PAsnIxOKxiarxe2hnX
gB4fP/CnFYRmlowP5XQDiErUtX/SidlbANmKBcI/T5vrP0ts5rQcwRoWSMRD5fQp
vME+n7+aDPpHDM7ubDnwrTtH9dMvMJhUaAM+lLPugogzz5+JebVtUrhRDX1Okyb2
5BWfG8X82H+cXHIVDLyZaifn5m5iDghus2NraxNeDQ/s7T4Gz5rP5QnsfUPG3LGr
+p+41OOsNxGqU0tKxUi1uDWYoUkmMGRYw4/MPDLd3vmIjF3ZhJzmprPt7mpv96qo
tPugHj1AY2Scv6k/4y8BQUMlDCIr0hfzak8e6GTZEVU7HQoZ0/TndcLYUdye82Z1
h5Hxobp2+CS5ck9FvCAsgJFuKQ7FGoLPuTTBF7g75m4vTfyShagxqujtJ3d9owz0
QyCJfuy9YfkdOS4OoyeCiFEKBsUlfP6XmWONeltpavLJgnE9xlQfOFaJASuacq9I
ry0IcBP5eJKhWJanSx1tWad8Z+t6uP36coSCCgD/+jkVo+a6zTzQRKh2UJTphrLv
8a8RBy2PYL6xyZ/16K+ow6K3/M/kv8STuW/M6mBN7+9P7QnFNyJGD+gHedJCF9lK
u6ib/dmCW1kXlEIvKqERjY5J3JUZZQRUu7TTHfWREmm/6c+acU+VPj/T9eEtfahP
38stzgvpk+3MWTUU2x5s6wPpP4R6ZYRONDPbXp6xxpGAhn1NcyDR+f3vQPlfusfF
KvrtP9DOMLSx89fkCZfvFJ6JJE6YmDdNRF7Bqs8NSU4N/OXwQmQGGrsJzOV9UKCJ
QdFFMoXtBcCqGS9SxIEWnXYH3dlUUtwqojQwAMFOtlyDg6uo0asD/jjf49k4/e18
3CKxjMW9fvBb+E9wyO81t0BHSn7N1YOnTeR/83CCULHoPQl/Mp2HDaj3ksj8eSX8
C51e2dUKHUwETew/0yp1ojqyWFQR6YoKL6wSrfQgvlRO0q1fgeKQPsxRYt9JN2Ml
WibPI/LEz4QuXFIKN78b5w9en3Tn+NGL0nbp1/821Vig584Az6t9yAWpD7ogCtF/
rETWz6ja+A5zBAkTg2orpu2VlRfGnCDYVFeFii0v6g/JnaAxxVpHYLmjKvT5ktE9
dM6m5MZhBpbng6URq7aiJmX4dTQn6f9Kup7HrANiodaXzmjVzZBJxLGK+i0ochxd
4wVPM+zg8WjLznuMePyt5aBZcOLgt6xLKipEJpo5FL8gO3WgVQBcCKn/GHFX58cd
aoczcXFnF0XV8NGhLJbZzG6SebJ/a8IMtmAFa9xRIuS3NXNyMMM83PWkUAfNINBu
FB8bKTOXjFN7ajXFhvCOSGPsgE7lnDfQPhMo1abLy6lh9V6CKI7CNJxpLrqxUG0O
+sKzmZvmCNEmz6vESJvZYfHdpJScNOZSZGSq3J0HRSrZ+xaiqkwyw81VxPNPtGzp
zZxqXI09lQLlmuJcuUHsoELDJ9Phd4fL6dCeyoHUnMIfqCFMBb5v6HkBbXpCZZ5x
0/hFkZsX73+P3+to7nYK110JfsTmQovupfZVAe926EMpDy8HR/hR1uC7nKtXjLeF
KUglrgeChYFDUCILvJFEut6GT0GI1R8Lkn9bcAgE/kI8F8q0W1nAKhvF467XuRM3
2hMCZ6Nv/DN6gqxX0L+YG3NQRmT7nqnbvXeo+xCA3arIQOpVgfvIIzrXixPVG4hW
nUF+Bgd1ZOs7qWMPob4v6JX0FBe1uiXXWWr7M7EoCFYQedXZSFN0+NbWElKGipgD
vjW3RyXFiMG8JzaLI4ep1DzWAkyUzcdo1/dScNWqyZJ0eWu76a4pYmc+JEdN6PXk
4g6CkTqvQXWDECcJ3yqsQGMYNMxsR0S+/rWxw1ijgqQAW7EvZdKeZ1i5YajQDHCW
PD3teZ13b9eMQf2x7d+nU6eTT1ErvbJyMvXg+ca+QjkesBlwD+mIcC2UAxeh17wA
bG7/g99JoMflZ6ndJv1mwP74YrBGLENW2sS0BaPtqeqzmx26KbkVgviVi2Bq1YQx
yqlUgcMIKmkJFvw9YipOx7HdWreQAVm5Zk3qqUgesdsBbu1Ayd8oXO5xw8mdIjng
nHhzUJ85i7FtN+05+Ytl3C2V+ifPqqaPdFUg4XJDzfi3Y7XS4GAHfA3MNn86iK3a
GKHzddRrrZeGG5F8Ltg8VtDZi0LqHD+I/QjwX9VgDjsED5i+lAtB1QT5yuQNAA1R
YiyYK+5ur+SOOLb+u0/mkcGCpElrQ/GdNnjsdxfFGEmSjYlDeor1UDC1veha+hHQ
6xyJIEx/OrIZ1lKHMkF8a4SxtTL6I+ETS3m0gpW/NX8PHU7Sl4KkEyuKoqhJ3Dno
YoF5jhv5ZFLrvvsv/QasepRmLMIsPA4UZR33jyPKD7dA614xh1EoR3XHIe7LU38D
5ImQ5dHZDndZ7kfun24UDlLjHE9qLo4EeIutlgInkQdEd4JqXhC+di67vO105Qbj
dkg2ui9QulpFl7QbGO8yPFDIrkSyJ2vOtqheKwQHzvqWH3of+gruDr338YUlBAN9
hAVeLXcgu+MgK7NN1WehD2CXrRF8TKfYVu+2O+YJT9Zh2fgw2HpSpLX7fRs/NNWR
RwVADxTw4CDZ8ER4HJLYH6iraPMMs9G4Z8tz/ECw7N80wxd5k5aysRHgLc9cL1LM
kH9eRl17aMnLCqVVUwMCrIAYWJAag+rifrJ5uHRIbU2Ktxrkrcv+UOBDxNDW5ACV
0AiPymz/cUGvWrIIIFlcbjNfHO1Om4U9SXy6KnSEcNyCOMWqUvPgpeO+NGckDzC/
P/5ClbSrm5j60ATXFbEpnpGCpz0VO8k5iDxo+CTuwr3e0nOyS27/AR9fnH4uvQid
+84NHuou3u5akXrvD+9dgma6Z+lO5No+DLwmZaIM7Rg/ACmqfcsKx+MZf7rg6FX+
KurZR/Xpbj9um8T8A2KDYymm1IpMeIEzsqzwMD+1cZKzEVGoZt/zhdt6oZlhLKfI
R+CyYIsvHE+NCbq+7QHYPCFNYi6+9JYmXXzOyWBNUfulX32w1iZEejoayckj3HVA
/fCOapUuGhK6P5tTxT96quTF/6x+/YgvTwdv5u0iHi6mxehMmaQlw3jCy5QH6cLx
wGSig5tWTvyw58mu7IbgjHcQfKxvrwbcyqTFZF9WOoJeNFBUix2PK6yXw6j9z6uj
ClljBX4hfx9K/csEy4IfLh2vVP7AI/UvaUYxVGVEG+hThpiUzgS0eSZSR20vyqV8
BivSae62/eIwyls4Uh5rJXzA3VXPc8bO0AQ53fQHC8CP1ANbwx1VylWPAxLku6/i
sthPEQKHbsGE8I5Jqwi2XsXEgd47zuUFDvTt3EMfkXbcwapqwSuwOXf1jswwAgpN
uB78BgjGA4+XjSsTqMajBPqgS9Krwu8r7kY/+J1jJhc89A7P1VEftE30iELedndJ
G5XJUb6TMBLUv6zq2ftiGjgW98pz0LNnK3qViAbvvND8g+yHmsZ1ROkoK3GUpTcu
l4RTFN+nOTo6FvciWhr03C4D7WZPTy6uZcGBsxvajsFGqW2PgBFgM58ZWbvSmFtU
kN5CQ+RnPevv9ZI94uAgq5hY0RWPtCOvYONS44yZHuzJbLoJ+rFbLDqA7L+NwQwf
ys+7dZwSISeARqEt7nxqsJ5mBU/vJzNBR8yL+Jt3RS1sIvOMFHvZfWyOXdOiuY0H
fLv239M614wHhyulHynWs7dCIy+1AYUmFTh69myU6sbuFXRQGIXCrBxLNFRhRHK3
b5gA3rFh7SsSKErtG4zVetHstg++aieteRLe4Pnxh4Pl0OgGg3kp+L/MgSCffP6K
vbyfvWmmejP9h65EMkwNaHhudMCEiMCg35ywqnvyNcwXkugA+h36kPmulR0T0EKi
qqULKyFpBnMzX4vY1lGRUt7mZW7QNdW0qqYvipiLPBEQZYmvrH5P4bSBGpNWKM6x
Qk7YYZfwl+SyQ8kjxRTTO94aR813suisj316sfT81BllRSCbssBntxHp5S7Y6AZV
gacmpL2mXZ3Wj4NmrSa0i5++3/DZU3HxzxdCKSmRRgiadRdtGy6t1Wa1kbf0HWeG
/I6tvd3Y56VwLo1CK20tXcQsEejqYLtXJZYsSyK7bpiUXwf726vhmtXkt0YCfhxu
518TtA0I3PwQ7BxXvMNT1Z+i8uRBEsTmv/KZMNltcNW9etUXKNIEpTKmAA2sOvL6
o9Z2QcR2p027IBn6tezL5YWJ/P4Ttsv8SEmYRcY5AAoFecOYh6zoqEDPuaMKNwDC
PHpzKf86nn19uQqN50E7kwlOPr/ggpiROtI+fijEqNrvbXQjGq4x9TWqfHk95yUi
uhrd+BNNqp2xHIM+yoRVu2Gj+pXjMzYKzZPJnUIu0fOvsHnI/iLoURHCvIRaSt7I
4UBz+MpQeB/btShd9HDbNpy6MDnkL0cRmuYrZ3Znqabe+MOVyg6m3orudXjVCHuz
IIFHKOl5dFSkswBcguLbGUNBFeK9Tda5Ma4JVHX/IBuY7jhm4kTZOePR72TeUT7S
+uXXPXOtt4vuA3tRzbwyl8bYp5+up4Kw4UN5yGZgqo1hvJGMg/Do7tf1iLeay0Kh
Sb/EHBCAEm4nTTcmVUThC2r9DrisnikZUK8brr7OG2AQJdXKmlSYsnSgGr09bVx4
5Z9wGdEujLVQa5+SFdz3bh7dUC5uAqgGtYmhhwrDuvxqnjzYK7Q2jraJLXYCmJU+
gZzhArXOzP3eQvWKzIEE9AMGaVRr0idBgauEXYKeSnk4E6++yh9DCsVSHyvOYK96
i/Dv7knYjJ8Xa2hPJfEC2pKD829ewqPL1xfc1OdDLMTN1xS5h93GqiRrM57VW+u3
fVfJEfPjLRJkKQYrPjaCQWwm2zoWDAbrC29k0CKwvrFPDab4MGGqleoQT2w+8I4t
ZY+4Hboi2iAbLc12gwii/I7EHJQJ3fLfFraZbmiY+HPw+DZU2Qv6WEwqu2NfesHo
s5T+51gTyeIyb9/MoKhoixCR0CUwWm7MA086EFmjkU7gOeFFz32vmrJTmpTcw196
l/423VekR+PuL85RrNrCa69HYM3bRQVKVHEATyDkcYOawhigNemGcSLkDcroxX3W
DXmLtMsrlQPpz+r81jOl4tSh1XBHwb8SaqajPLguDsk2FI5XFqPY7xCy7o2uoQRD
dxKUkjG4ViGjo7x0WHidHKLVFygl3XKnXAIarmd+MtuZz+cZQsf+/4MUjGRkGXWo
VHco86upLEiL6lfUYUQrTAeLIGwVg7Xi44G5x5xvA5ma/oaNqHRmn9QHsm30N5oA
47RFdJIXw+HtO9XtFhCcLHOu6jdoI7pMX2o8jFwRwUSErddMMj/BqhlpbxIaiMRS
OhoK3DQberRGYM0Folz4t7czfR5nwFpRdPun/Pvj+FfcTePJ7cxt1NrakbbzXUaP
EpD1jA5Iu+O1k4AKHJreeWDqsrJdgrzVROrizhZiH2RxcGMutUCbTo27Jo/dXGWc
0HeSGNrcOi4IBjC3GB1oWdEtSJAcO/sNe+bveiLZc0MPWRv8wYq3uVCmnNS68W5d
326NDzI/Lds5WemHAPLz4WhLwWv7MsxFUyaWEmRj0ZDL9hMbCmvSHfwcRSx5FkVG
vN/mMmDgEgDod63z0+DsTDQQ0669IJYNYE6YiFIhf3wHzKR5Nk9I7PkmokbZO4/J
uCMuHOuFGnaNraKCiz/DnCdQcRaRRF/j/e8GmF74SQf+J+cxSK54wlcjkeilZd9p
HPFiSS9F2+/Nxgrq4bze3FMvP4jR1LK6z4EuXbl+BWfnXKuYdRcpP4eZGNUU1i3Y
2397b0ZEL/f55vlz8pdAA564ovMOLIdFbV6jS3ucS+0e3tokurLcJzcvrYSHC9qX
GNSJVvQPj39yWJx6DM1419SOt83sMIu56de7f++jxZf8H26kjDy+ZxvF30haMzgh
Ia+m6iUBRCkDhggu4L1XyYOVCxmC8J91IZBRIopgBLx7MEd1XKXW9cyKg5QVGr4a
hck4ta5Be0NkIenzFceja2S2eTxyDuWS+q6g/hxRdXQaBUW3b3s4a0xk72tBMRLv
I4twHez31Y1uPPel8jMhYrhTBaPKaJg1mxfnHtU79DD0/+XDgSi/tIkV772wmhAI
MP2y/nqVgPqF4XFBLKvCKyLttnCn95UFO5c3/249TcCOkP78Tk1Iv03IZu1DGgcq
GNL4mP0I37prySW3kbbj5P7wIPNq9R9oW8EIBeE56E7UrVv2DwgmixyWsyctzL2g
93792DFsjUMKVudBbxf9vOJvHwQ1AXazDh584fPqwTK5ptRU8puBsDCjdVFHt7zv
1SeGt7DsZ7EUjWO9+uU6hiQEYYFVbem2GG1pGMIcAimpQirzB2QlrOaHFuVj/fh4
erBA/wYLxnPQLkge1yUXArS4cQRlhc8/mUXaN5DHR3160uJlVOleRsZiZhinU/AP
5pZmVascXRUAuztfRExEgUpTO7nAvQM1Z3pjzkIQAoKxWPE01woQGAYQ89jTWXFu
hi0rGMT3c/yJKNGorIbussfxZiWfBS+ph3pjtfqu6a/g8D+xnjo+gDivXFQbmGHS
kUXrTWFc00OdB8S5COZIHga7tjc6DLYiDQ8gcmcYlInRJTW2zdykqnRTmA1tTQYU
qJaM3vUYfI99MZfYkzo139fiX9Ft1JT2arhMX3FWTs1EGKsLf2D/anG+N4wX9PZq
tr5+BM65HvoZdLFCsJjBEOScaB2RNJOI7/ORO8CiLhjR2d7fu3n+d34phZKuonlE
EOopN2EE+BV4YvK2VL4NYH0iR8i7HmeMzUhIj0H/RgxMS9SldxQjB5roP+dT2m49
OTGh9FzBpvc9L3+dtw9Z+9hDwUpZtUjfEBfQgvPr+DMyxAx13otH5/RShQ3CX+qC
cQmA9vwvBV7W+WHQYP3BEwuoVBpFDDR84bZm438LeQLghs5VrfLFYbirVa6VpL24
oDaOl3HCTkOXpsdwUi2D+IlNHS2O85z6PZWhZjt+YBQ+ApmH9/LASecGUEnL2cxN
RwFd3sf7BdE9BtzzbnEBqCJ4ZDjb99Mw9pZERSXfrKLDogjH5Vv31Q0Kxgg48/sT
0CKQ+0X9k0G3bBpSeJkeFnmGnvnLa2955V59NXBRw6bizqS2uuN9SQNrbvuVonad
jKyE5+0rlcQPn7Xdi4RCi/mR0kpEC1OxQk47weD+i+wcKXKxnGU4T0WX56B6CaOg
aHM5xt/N/GY1nzuHQY6Rs09low+kwuASjDcBkod2RI/ik1HX9NcW1eOsT4chOXwd
tc3rjSkBUG9rvr5Bhp4NT9kobE4ULiry7CWZZ/KISNbJ5un8CJfKyYcFLwU1aDLx
ZczlU9EjXNqvBUimM+pdoeoqg0/vz3bmmDXXYtzn66TsI5D7wUE6+hWEBOqCNrA+
SN3IC/6HoGZyLV8jqJi0agXXZoPIZqxItugwF05aR7F7zRBcs+3WtDzPUbtOsYNR
JKY59MG+GIShvoXZV4nzzSz11NfGHqYZe1RgkU3GePxS+Hf5lFNg3DMnqbQsJmwv
3QVyffCE0rv/1fe5J2Z2xTQO8buJq//jxEnb8/a7XMXoyT3rsEpGGQ0E587hefsL
CHILcQBaTi0ZFQkE2ALsHcekiGqMtbyZzoF2kb8q/eRjSAvMkw9UdXbFMhdQYpRp
shkX/ClpEYlLzvoTUaQPSMBKP6G9nTfpTicyz3Ww3mIXkIc2F9zUX/oknQR0aHFI
r6f9ex+Bdhp8F7S3OdWjGs6c6jknMdx//UQ3P72cHgBuDaspi5WCFuGyPUyTIS5p
sXMQGKNQr6Cove539du2xWMEcYm9xWV7Wi9OgMecL7rrronfsz8mcWlBdNdgDiwt
RVlezPITnHNikhoNyq8QtGvmFBoEeAqrSlPu+9tpBEnFg7uAaDBdRNC96BH850Ij
YumwIWt6b1e1yLDwQj5S8isx9m5ar4MSgC/oZf+M1cz+NnK347HTAw3BTUESdSLM
i3QFOfkFRU9r7S1yxfWdnXGN1waPnhzSm7PcMEo4EC3vr+ye9D3eeMBJTejZD8oB
uDNMvc2gvaT50b2aaa6Wo1Qv8ar4L44JkUZwVU09Qzj21QQHDuBYMIJ9JMv3gT+L
1QIYE/2ZslJHaI5YfMwO5lBC5tsrpbVoYKdT77wM87OMGcLbx++Z0yfCgvtXkfok
ABBkH/PEq2TOyQ8sUOXE6bwsEJWSYBi81AQ38v2QxF0809hjVgCG2F5o4LQNsZzY
FyqWNm1zoDZfmuAf4BWb8VNx4mneKmImLCoQgBHhpXd/u0j+YVDE6aNc2ZF1YfpU
bFIPFY4HQ2SqQjenTlna5+mJbTkWNK1atci3wsn/+jn1YFk8yiDWh8Ai4xyTUVsa
ZGGFKL04ZmgcSBXSbudKRImoMTYUz6SaMJuvVKk5HDIYIvQpkd2Vr94ARMK4WebO
e55QLa7pCIO4zYIStaEbxIxKIiJA5FYt2ZERrXaG+lYY24dxBFNK51mL13t57AGA
JPqOF2bTGt2g0LpoRlwxKWYuDOrGHI/R27N+w7aTamR+31DkeeE6mW0fHQkWhzG0
Rer4FG4R3w2N2l53hd+5udTgQvMNea74jfhERZkXCoK42UW/ooVmDcOVsDd9Gihj
+cQTHw0c6oRSwUJaVe4gjL28pp2CrsVfTouXsiNs5DhPmLfOOUvMSdFFpwvgKi96
xDj5YvBEFyswxxyEEJjO9bQNjeY5dPPs6zIgP079qCR06yfxFQYHeeMxx1BI5kHa
uJveUyQcQb5f0yHmZ8MP3vvZXoO6sBHbGIxW+hBoj5++025GHN8cyNlg9KiNm4sE
a68Dj1tB4vpYlFgIAUkScEecwbdB5vOWQuLdTHoT3PLew2RiglAjqiJzSgaZENl3
TZuZu+CFqFagXLMwk7kj8xnKtk8VZGhbEaMUY3oefjsnnzbrwsOewhl/4Wx90hU0
HqqI/TOLdB0VAI9j4F1c6Zd2GdMhtSruTgsrSmlTiyqlapF+/FUdTD/AI5EfSmEm
QKitI+oHyw+cTqEeLWsE/0NYIi1kZPg0wUsFuAYymCiIRwU1QDG7Q4d4SpnulncZ
QUuU/5rDXJx+q3nptXoWQp/9KbQrJtSLfDHWvznYxZ0/A15+jQZABqCRN+XSv4ui
HJhwdlsTh0f2Z8R69pBuRdMnuOJWyxbUtKo1me20Xz9RtoTmwuVSXCjkENGADcwa
7MKAWxMJ7kUW4Y7PanYh09Q6oRLfvzspefiKBATssmurY5iOgVREomFuhmSXCWOc
bk4mi9KCwulHr98N/yPf01ZHl95JsJyLWgsHX25hzUZ/jyr5SQWbo1ed1VhWPJeh
VzPdbemqk4ve9vAHahRAWFcgjAyeWSJJGe6QBBzyRdGS+41cfGnr2HRw42jsCgWI
7cNLM0p9whqKkaw52TXz0np6ZlTthJ3m/tIzBqTQJ6gEV1yvMnDZl7lYEawMze1O
SgLO80/m4xhUkd92BNjxmpGmTLp56Z2dq+KbI8duDsdJ/QwmJBrDUAtuqeUmOizJ
BH4YuhWIHUhqgopNmjVPY8nUE+a/aXflNKpq4yH+1azdebu6q2IUoQU7SmLXtjVQ
PX2KFfkAEjDqcENERI0eEgUb7hiln5kSpqyHDUb08mTG/cASFPDwYT/KrxQuHqVp
CcHfN/jrvxWoMH41tRKSryAXSTvyjjCfZHqSH8L8vC3tRCInp4XgytGAKbRfw0E/
qPSwtMqoInPdo827lcLLN63+f4YTg85lUuHBv3aF3JYFI0uWyOwa014fdXa7iYyx
6yBz+/YQZvexQIol2HTflrdVgKgn8d2u4QgXtNc8l9+XCOk1fw1NJB2Ln8nepbZK
8KaIq7nsscrGccjDJtqLRnbvWGXEoCTQfGj3K7s0KZbqtgoGZbV0XtOxFvLy4ktW
ppAag43vq+SZwwhhUHqzqT4RteTRCdgu9AaFmp1ino+zdN+o2s3M2dXgBw6pgYvI
8YBABp/3VsAlmHzdy3eUonhqmbG4PSGtTC24g1vciiyoCN5g7tysLoesBk6QmUUg
9+g2B9mv7K9LRJKDciAe++Z4zLV0ntetQR05HiEEYOriuhk3I15iJl1UFjZHmZZs
glAQ3ISj3UiWnfO9jftMA+eEyFN6Nlp4Mvc1yZGpq4i43BpilGOi7cFHOje4cYEl
ev3GSb/V7Ma4BMTIo+ErxMvN+XNxfQs1F1HnznT1EMmMOJcXNPggSZedsLtE8sAY
OaVWO7+eqHxNpZ2ZgxVI+rguY4RUQFMkeV9r9+2YieTtgNymlYaVP6hxwfOKZ63J
mXfZO+01Td46Z7M0ybAr5OmAZl25KZH1EjYIWxf6jxbzUQgcPM2DFK6H4lp0avQs
t0LCuCwbi2hN+cKkg/IAlAekXmo9mFb06T//ORmuT7fuEXacIuXtZ7Qjw4zBRv5n
eD3NQs+6qohNgCroQ1qrjqjNeAEb11/sgkNX3eheBK6LC9p7FPmcm1mwHwaqtiz7
hU5Kmx9/0khSP/IXqRwZdKdQvPMpwj/TcGtEUrOHPlG/TelZfpdtX7U42oAf2QYL
ws4ZkaYxHPOggFJoyTW//kS73KJqy3H+Uoc3XBDKxlK480Ph0L4TRnOoh5GRrXci
e8yw7cC5Il5yrDDy+UnAy3rY9WahH5E0zXzl1IOsQ5rs7BQU22CoiW2hvOEN+xE4
/3mstUNUfTrWxJ1b4CS/fzNhL5AKwSy3K1BsnJ2sjZ4S1KqyEliR0UDlbpPuWg0H
zdbdoqGxeFcVwBpILYaPDhnUj+2WjWLXCG9kIzOjvmlN+iTD2Qq7pfWaYzcn9HKX
5UhZVJ2bMBh/hDxUrchifdLlkFbBTwTmCfuh0SMKhpxkHfyxFFK4fV5ApfUVUDwj
h6ggUdSmSoQnykOgj0CeQnELgYAcmY//50RnKTHP8RukDUWdJus5Vt2tWlfkc5ed
MHEtKSkg+LPI/H3OvFdi/O9cUY+VUzijOTMLop6gwdkTsr+aUmZnk17z3WEBvdtS
xTugdTwQbOk2QUO6WIoRqfNNsYwQfMHKpFFClsrEYMxoRA8qDr8mbOldJ6DaSpLd
fhAk9cnf09+tV76+IIU/8wS9/KdeP6hnZ1dF6Xr83WuWyvQy5qkBmKqNRF+2gOEx
Mb4iz64Mg0QfpTB7S8uakbVEJMAOIFHDTNM2VNUOtaUDe2oPOg1HUIzVHhN+eQEP
a18f6rHqCyZbKZPbA/kAiNCP6LO5WkqvVyLWdPFx8+nZA1+7DtvI7Ri52WTnAu1B
9f5BAKMinfb/6K/1iSKkHKgDj9YNKfa0nN8UMgRp7Q/djzizemTQXzX2cSnkLZsx
6pzt2EsGt/xwwAHaJuSq7QSotkaiwYGVSGoJ9LF9rRvukunjzw27qW0naulhfSLA
eT2UF+sIsDUFHSnLGQxx5jyPJDhFEwOGacxkFyeCug+1h7LOV7kc8gHMJsLJeb0p
oHMEMZw6C/s+kbdn4Rt8Ac75sB88KSE/1Us4plwuz7Xt2HcGUxbx+yIYiv3ReNTr
BClgmuhhW7xQqcHGL5gPsspO7lu0uL7NasRJlI2/3d1ntoMJ0LVnfRF9+eSKalNk
C3I0hI96r6zdWGpU4SzoUwS7Kmu1vKuYCtbh0QcRrIh86GwrAOGOiwM4qrGOe3zu
gckLwG3bC7sKHIeM7fQKqJSNuI3Ddq0yRZlFPhP+fe+B1T9DkMwDFG8ckJ9DAYjM
PII69pha8sEYz07I/zfVvRtDuJk12znzmCp3+YcRv9BXe9WQcY3MifFGNotL8D/j
LSZ7b7Hrsi/X9pW3KY36uV9EPBKW3Xs7UQYasr0Q6j2+stsFhCfcM3yn7pMSF1WR
Lalrf3b3bn3w7F/ESaYNOJtNd3GFqzygXsSiMKg0RbsMNgHcA5qYl61+JlF4atDH
POJ4LOSCs4dGLHXjNs3iWWTjIfZheyoLMaKdEh0qk5Jgn0rXMfyxJHxqyWhV6Sx0
kOwpmY8oICeXNcl2PlbkQexO55Q+huoJ9t3TVQEVFVeIUeCPcZSLCPE0qVqIUnR0
SAf7YnqJcgyOgtmADWv9/VsRX3GOEbaJDhCTZgTGJ2LXpSU67DqrOk2s5tnQvw+C
HHYBF6RW2lNWdxdA+n/82K0pUTnTrjm20r9W5kaSqluCIz4h3Mdu2xRLrcAQIyXb
D96DkluQgk9BTWC4jwuqO0FnoQlhRa2nNsLTCU4+XHasr4B/JA+7KdP8YfZ90ZWd
5pUd0Y/scLHh1t99fiHUtPeXLT+ZF2ayMogfzZzC9G26LV3hcsSAJGPqh7snSENQ
6H1Ue8DnYUaezImQlE8IzJsL7u8Mjv4TYFIjNkP2NwesRPDttJ/1AsIfKsfXhL9Q
xm56uvoxhQRy+4FDqyX9dqLeivlm33OPoSMunfmwZNFl9swA/NzMfhnsAyrgfokP
jBID6Zhau0hUK3HbmCkMksUYo8crV+UnnfhZWGiW0n99wb7oZOpK1vPBE1Skopjw
cvKDWLzeALK6SRXIbmR+oZqLc6QEnlghn+XGElXn34ojvOelFd1wuPOp+W7zk3q2
4O/HKsEfMcM1hZNA6lOhYtY0iUZ4I2xX1X+Iki7SmGMnUk+IBVkaumZNt761Tma2
YXcFaAs2bYI4gGZIRS9zJtfcSG9kNJwg/RwXWtpFu6AmfmJ76d7KBVVsaFk7TkJh
Y8cVBAInfvh3y44hSpXfFdT0wfM+6uuCNjzb1c6rsSdvZWFmcOOz06ieZrxsOC/w
awfXTVTUrWyrL+uVLOYbMiYPGdMciLY8IsmFxcYfKz5XpoRnBbhWiYbcJIKjcPeS
/jnQZzlDOc8jhYSdianbnV8X88c98u15v994UXwiSuBb+OpnAN4lmaX3WKKcCun4
scr0KCGbnIVT8G6Gtu/RLWfyp+Dt8W54RLbw3+T12Uf4z7TSr9QN2X7Ef6EgbnLR
rAU2OH38neH4fdvQZvlJbVNK2PhO/xH+Ksxe/omulcszX57Ho4RtgSwjE9KeuVAI
1pOc6KYwPMmbiE2LSu+/u11JTSPJEotwbnkaw/Fo6GZjesq4QnFoRce/BYj5yf6S
G5xqQ5y9SZQjaQHkbVew64b1ApYELSlk9g0eWozsFW98XLD0OTvBXBwhBpoOGokR
jBhfDdukcuXZlAyxdOYkBHAGYMDLEBF0LkJ7iYlNujrhd1vOFmRalJ9ZamUtNKjO
vlBvaqtBD4RDz0qFVfS2BqsNNbzbFxERJkU4+CqwJobVQwdUwlh0liTgH2DA71kQ
qMNN2BjRToPUoxjPib+rC2on9fQ8Cmp5/lv3W0Zfsw1yDboiX+TJaoQpYAU4d7oy
/JOeTBT/Cmzq+FvDqKKn6lierJ/eIjmh3NUrTgk+9TFaSpeIMW4vaSg21tAzmg1F
XKBwRMJbZDD9xxzrjKSyd14+v1mXiwkB6EuFrkC3UM7IjZVbIbq2b95XTLys0UwL
amCmFbRziC1FvXiggaG+0qr4CLbspwjMLLp93+kHRzat5/YqYvrZNRs1bkX1L5Dx
m5/aehiYq6Tg+OKHjP8qRR/uT/PtQuuzCVL4OnF+E031xJDes72y5GLcBkTt/ytK
5A3Ifq+ZceaMssb73rdjk9W+asXOY9n6j7e+MiUZEW80okL49GaCZ30vD6Zsqq1W
R2RcMTAgQLLZWt5FlHV6T0oWOvN/pvTHc8+ezgXFbfM3dAmav9mcsPYsVss/Msp6
iEHoU7s4CVhcX0v5/Ugt3/R+JchA3l7B6GP1sb9e66/arVKmwvq3fFvf0Th/QnpD
jEpAIUZEO9m+iaw5SjY6xedMiTBNimC9RRyIOriTtbZKGUHPp7kySCxPEp1uDyWT
KOYbFFdWqTIzC8nGipwt4A656v6e3b3cmsos4aFtHhwr8nQoUUqlCLJtMkxOVZVD
mWw8aZHWLpsgeLRupkazivtf7gGAKDeYa8W3m72ya6b0UTEXAqzP9bRE1TPrZWH1
zaUzerLmPv3bjomW5YtShiDaebsqtSAOr3iQVIlOcTJqaKwha0IA43+LuTmgAO+O
2Iajhp1ZXqbsHgpofyDipMVKVbfZ9CDAdTCDFzR3NlQCQ0w+FoPe0BdPI/dmAzde
jPgx3E6r2cAKerb0T41KQ603ykIDHKiVG4Un9eZyrAMlTB+53loz+0gR6FB6GeoY
lquoZyn4uLhdWDh3PCrfKA0pxCMmIDoE1nBnyTngIReAWLcO2iBgJP5T/r5DzIED
rSqHZJUOWAv691SU5zvRr/wAZWnnlJiwWY7n4mBHPwpRENik9E4wdkdDeJZm99VO
bF/QQKn+ikDOhCILbIpiqyMKhHoMRid4+OAE5bR6phxZUvTF9uWaFweiqdBO8nZt
zpc4DQgBa6fMgahn6VxTEewAlHLnb/7lD+6P1tqQ//VOaMtkVf+om9Z2kNWbUtpZ
Xbevj/Ts5sLctzjmrkDOzOJkM4XKRL7woWtzsxodOezzHoA+cU61pinHUq1vOZ7n
wQLgKXupc6JRb8gR6Elsd6b0LvsXqLwPLBMuPQpqQDJZ7340b6clPbBqKLu4a5uj
74KGar0SsQ6oXu7Y9mRIFuTGILlRa4ck9gj0cXPOYnh+nvzUUlXheADTjjj4Y06I
J4CcxGQR4NLX+s8cVm+UzWV6OkdOLhPvmUGG3K6zT/HfMOANfOtSP7UNdQZx6Zz6
mDrZgEOIIgPoAGc0YghdGD6nrmpO6VY2lq8pQztFlH6t6a0QIqe3Kk6iKiWkofK7
0Trf75oTsqgLAj9XlbAoja6VHmEtIv9pR7OPk0HRY9/5hJEi1k6wtTwRSJhtK+j5
EbyUjQoDINcHxXws7TV60q4txFoAylKV23I+oECKqMCZqUOXj9Jr77LRPn8AW+KN
ybKDNwlQOGiLCuEjbGmutVL1PoOVFTNvf3FzASC2pinS/a2snkBRO9G+g9JGvBXr
0btzTbC1JbxkmhFl5YVv+7EQFqaqyYJ1meoFiHBbj2UnKjBfpoHROfWu8sZfzPD4
JYe+OFAJfDJtVa32MeVn4rv2K8L1O9iK5FBS42w84dDHj6qt8LeI7yXipM2bxIM1
KaFcrVwX3zx10aCnAdDodR1py4WUSTzQxwrex8kodkDNJRnDNWliM4abZMLpSfnX
3rhIWMrqzyUs9RgxJ3vMpqcA4Q6kUFbGJs7GHd1wTols6gl6yK/c2oMFILw6DWBJ
iS8+LkjDFiIOn0PX8No4+QHzhZuzlni5sH0ruaC7ZqdxXVwoCmi7KuQmrk6maABp
/K78UsRP/28bairRi4ggAUucEO8GKssB3F3+WBPIIuWr5kIgz/U9giBnPsWjcOcP
SLddn3d7L5EWdVZ0porwBd5OGSy5E8ynBIFJy3GRiAMJeZa0V0gDzZD8sw65zSP1
QbwxQ8gJ98vUbpFFsP0SW1g+HB54pQR8dOydNZQaofHquEAONsNVlFTtwscenWFT
OW7p/mt+8okY+FDH59/1NMOWCBKwlnoDVr3DFSNpzdIV0IEe9xwcMYJkDvkGSgwz
e5OUzPudDbc7lZR3wk2kO5tahQM3SHX1nAvSn31VAWX/1sHZxCR5iwfwMLoXA5DN
hsfixE6/gcAAgo76UlUmv83Q19CkzBA0DNJVjdmUNmqwai6WHBRC8boUb0+nfhWu
swbO1d6eR3dxQGgZ92D91ytqi1EBPAYuZh8KkEj6n1d2zZvxWkPDwBqk+7Mt+bqn
ntwkqLKRtMLAgFL0uj+MNML+Q+OEFW0wbZu/BDAvVNjYdD8/L5E+LA55xVEOR1Ps
aFaVTZVOF2/6XiURIdzmbeUpQUl3ruwU2nr3XjToilsoFLh10c7D2Ag8KXNKLREB
4lHkzfRe9zC1t2Iko1Jniv6O8WZtPX11Ek5g4WIwqNipbjxOIHokiFoS31xvNUFg
4a6P1Vqvzy+ozOHD29zBlxXjj8s7pggRyVButU95XkoucrVrldiAwVgIuxOpOedh
ksbG7oQPfSeYah8itFbkhomgCm6oXTiNs6SlQUfT66LicRhcoyYqkb2Y6d2/JSx0
rVxuLjwnfD80x2lhfnjP6fVXsqzmWnTYU7eWKxgWzEDP365aJS4NjyzIa7u5DP6w
x8MqZ/KMxkOFEsvLjz9E9N7iIvB/4fIKzVdjmgQzNJHVikP7DfEW9BgvA9dBSlNj
VJTjW++yS9hoBhmWAneLGHdueglnHrnXMdl10Rd5ZjD7cqekq8BE1TAu/d3aCubu
053y4hMjsHfUBXa5DSp0vLRjFVzatXeqzV2dPJkqziRPG3Aw23ynqp5W/hSfscLe
UPr5czcu8LDgk7l1bQFQzpukRlTNQvHciLOJK+f3vZ8L4wzqoS/1GqyUT9SxwawA
nZNTAIy1NMSj+LxWT1DwRRoXXoEyO9JONpYFyoxMUN+JrTaDYUA8gfrP9nGucbtP
gv9mwS98iGwp5ZoSYvVqYmpbEwZ/Dkc+dwqUiA426kA85iGi8ky9qASSBqaSuBEL
ogWMOYMF7MPSqbIk4qcjK3L3JR6ZehfdLfVJHy0N/BlYWipbjwWocPiXxl01zqLq
aUZP5c8Q332KnVcTFh5icRwtE4acMiP2qrMNWbC8vypzvVX7Mh1LElZZfhYZJcPu
NN0PW7gE5kZW5hnhbU4UANJ/D+nOSF6fG52XkNUrGspBBCwZTkoOiSpJhPFrgqTU
L+4xwCGFgkorhbccW00X+xAmRfIF6JTA1ZmczJYqjlreDT4Hs1kvc/PcxzQC+kA2
6Dk4MwiQkslLQwuPNmEUlMu+3QuCoRX04PcFeuaHeUmWmhLZSTi2QbK9AepIqJBK
ffCqbZI+xSv9XQn5vjxTuqyHfcG1cnbvdbuELK4iPtjpy8bskf9tWUk34BtDQJqR
ZzdKg+bnwpU5jFIEORlnXgnjFWF5y/fM3RUngxXnmcW8Zju9vypSCr1OR6XLW+M4
ZDaf7+TORxO62Vnh304mEQMNe0TGgkma2JlGb4EFerL0ECYQU2KaO2Pcp0sMuP+i
Fwj035PMloQj6cCiBv+9n+uj3a1yeDXL4Emok9iZid3ATMIpabHbqNWq4p4TN0fb
TZ9ScFRRje5WGbR1ziGYbhxmLItqNbv3DQq6+wpxULZdP31FC0OiP6JGwxxMayRi
T0BNPBhiN0vC6KiA9g0cNEDocSFMnbLf/HZK2j05d+OMjAVYX5bFKyqX+3SL2a95
let1oh36CSxynep7gfZFkPJVXMu/t5Rf4/ghq9q2xmVgGzYV1PdPRR/5/gHZdybE
IdjpeEqLqNEv0VopXPM7ufwssoPRDKjsqgLShLhTwIcWkAqpvXcTLV9tGO+RjzCQ
OsG3cF/2IV4rVKMuB+JBLFVVZJgpuebkU0rAwpCNI5TmV67ZBc4Gq95nJoDuPMor
BYnK2zXXCVuSKP6AFcrqo57dUrwEmeqTKqybT7eLz/Hxwsy2pQUBLhjsS3YEZa/f
BLFfKKIKqqueLANG9/7UkupCe5hE6PRN4qOzMjSaOebAvVL7f++0bdw8E/FRsZHo
2yzcm+ci+RQDmqXDlpy5RRVv2l3MQypmoU8OzYknBLZA0bzuZ7h6/sT+W1PQCttn
yDoCkE9hGvg5v3Z12yKjTFRJIRcI+DURC8U/tJG7ArJnm29u8zswgJTuUZz4LJxg
SR5cGk2LrI7DPHVLK8tiIRJgY9uKwDYOoebGYTEVDgxswYgS3kg8v2FVtvIkSXTy
XFK/gAgXA0DrIWU5l/jjr9Xe2YvICYyBKTjVNSea2rfIzVh/Dh6voNUPY1FB+Ut9
63aj7rbiKEmpvJheldh1O5659/PdmUN6iVc1IopSAoIa0iKqCTqRYKFc3bRxkU89
OiSmWqk67Abu+CKlW00tr4V+oVNKae+9I7e0/S5LlOTH3ZLd1mZmO89NcyJLN9lW
d3/gFStvbiIxal9bscA/4MxxIk7RysmxF7d+NuYWrL29SXWY9vlTsP36tCJDz/bv
IjJ64jTSoLylkglFrUXe99p/y+O1XE8YqDJ3DUkhvYw8cviZit6vcnAYeP5KBBJ+
kSMXezH6OwYECpsK67pfcYSz5ERqQFG9k00RV9UvHxYVfx51i6+DzrA0klvXdNwR
LkMrIvMWQFESwWsVxk/mdD4M201TNNyE6S5rRZpzhfycxozbUv6xQQwwvisHKmsD
hsVYfCxsdwlNpphnBCMlXjqjY7/SpIzAEPbgQh5ttQ1N0pZESWtzuJfBa3M/EkvI
a+L+XI1zVbrqlmE8cp1uo5DxFGxOqZJSg539F8QsoAF7+4CYlGh+PJtZkb1fF1p6
kJLCMaZ1C4rglgwipaG4Yni5ACWx0Zk9Bj9Su4GRkPLGUrVOR1CtG72jnR5UBE5e
LhVbY8+gG8dTG+ZlMuIRaW6WUrJnxlK5HqNmgdHIg0h39bkbZNIos6NaLHPM9jfW
GGFesBwVFTlvXcJUzPQseMZ+Nomi82fNJO3t/lizgk2J9jfK8fOc/Cyl9n92/gTV
9OvEdpJBqrlInuORCbyeFRdYpk4RC8vH43Pq1GKAECD+sGyMJJoSyzpYPEXvU7Cp
FFA9sB8rCdjiSaAFGHvgEnu7CWehq2AFlmFXth+qkWVcVtZ8Wg2ZLJrSo8jXESz5
iFcu7jddrhPqfAiy81BCRwjk18fCPBCiNQ+iQ93BSDsoo70tA8ZqvDwo2j4nfZjc
axUaLeADTZJibDYu2B+Pa8OMPqiyJrEWDaX95yXM+yIS+2OSkOuA9utBkE9Dh5Bp
+v60pshZMz3Npj7nqAwPAUnWR0FelbT2euXa2fNZRGcZbwuyAXB32EF7WvIba2Q6
msLojCQ4os2UOb2SnsLBHI602E2WZ+koAeAEMPseVj7tNe1zMHgB7T1g+eMoN98t
R2zOrhveaVLKYqmZlAPC4T2w0dvQkup03yIQRk+F1nLKb665m2vHnvuL2LXWhKdv
B+VNY0FspamlN9QcV2/5p8Gdqj+eXfyJrSPwphPQFG+FIbIQZHavbNf+pv0KkzQR
4NrkPN/q7Cn0VPoN87K9ol3amKewHrRvUxfr9LTDeZ9TRlb6AtfaWta1e9mqu4fF
V+xqU932D5RRwxRvvbQcF/Ynz/CuTFxGoUFKNeXPDlLtcg3HIaIt+zEnAxc9MtPV
OMBMwjoW0vqA3nbr2IKQgYZmGBQthExLuOCkVsOCwNtYK/xQHwBy2EPKXD3PUT12
oJOi+/BYNWhv6IF5fHRPPQ+tBxjOGQiErnMh8XlEJkkU5O+xbms4YiKeeZ3KDP6E
6uWfr5nEX+ySCYs5tVhcCzSX3T9n4ZpYr05M7l+O0MMdzkY/JIPi9TCCgDZA2NKB
lvNRaHbdqFIBrY6e1jiM9KxB2ia7rVPqLiwmFT2c3TzvyUOZpzHfgFZ8N5Q+OOik
ZtdG4aBXna3+Xg5ArNbjxye3BmI68R/e8hF/yGHlqO4MKhBonrBACmZLzNBPKVzT
A7rsuFPnT/mZqX3NfNKP2JhOcOVfU3SO+xdRNOyW1Ri/sMRkgX48sspYtbmJl7x4
Lz1+veb8t1RSEIce+efpbasAVJ/cEzSKdkiiXvDIiBqtmj3+MjEaTDkJabrioAs5
MzS80cdByL6zzwd/nB+Nx4lkjhDWeCChmUT2YKffCB+tonOzA/BKROTgHEquIX3i
Nrc58u86TXhzxakkZUNXkKzCo1BWcOl0xh0pJ7ypIQlfdFfKVt1s4k62G3AvmLxs
n5pyra9G7i1lrMf2jpqkdL7g6yd9OgYPZXu3oFAI0HAMdlzuX2QhnDINTVdThCr8
Rrril0RcsVKBr7o/hjuYHVhNe7gfNE7Kb8aeZiVwuPoKzgk0hXQ0JPhdRdhcesVJ
iDJoyQKI24U+NMssuN82fLknviG86u3+0Ooi6y3O9adssjaFpavVte+yQKtl7pih
vh7IKaKGJ66JxbGjm+2zT9KMfRJ3X8fl4wKDt+sVMD+V0oNwPtxzSs27I0lVq2Z7
6Sh7c3NroW1UEYjb56TgbCmMnnyWvSV0DlxxjCUXBlrMi7B6Y6lBXMNm/R6xrZd0
Rz5l8VN265i/zVrHJKPb2RTTt2bMY61aLEzQ8Vf1mivE/mj/35v5MqUzYLFcP2WK
Y8rzsg1zs9v2a9cElvqq/T/iUjZ/zpBoe2weBtfGUKh4deffmS0wHOmfR6zJ11mH
+1saak04YvoQrRJEhMnKjVZBSJZnbYcBz4HmQwBxjHPoNvZnZy3EdEiGSO2LLc9y
0/bbhe+iWO+7DwBIFtdfcf3hz6wLmw/xBP7mJKOV1mhgyjbibY4Rmx6z+3WE0AZe
j4Ex+BxxFys4xWFHEagef0NFkJ2S0nIJmVLuN0f+M5nTGz9Muv7QJKkrtG6OAMPY
gMHp78FPQHKrZ4fVsmOWCo+NioPKJZd4DojWzHMvIXJpSatnYjwu7iul6LENSes8
xRDIucCMiLXRGSJVsSI37ooZ4G0U7acq6mAsSq5RlJTYz9GSbEwl9lK6aGkahnGr
`protect end_protected
