-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QjLWR9H5eV7TLQh2ydTnsDK3iFbqonyZFoJvVry5L4ct2q3xMuZLHY66A6v2fQW8wNdHgWRUodgY
yxUdSlNxWYs464FNPD87snDVCItYrNvsjxXNIb2CoBAupZzENX5OYqKUHDGy+sYcxwqfOrvjXjfi
FHr1MumptVYw9Qq82hRtN/uxQJ9QvPT/w4JXczAr8TahjPFLTNAhrT/b6ENDQLKcJUsphtutvFJ1
hB7RqEYJP/A0K6L6NCKoPB6T3kaQvRCDGKfDImwfPZb1ZaFGYkbyQKEhNU2lvWs5eqPf+1oCbj2k
ZIZFDL8KMKZ/y1Kdvxqge5QLd4B7osvnJkJYRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4560)
`protect data_block
FCObetYJLQNHaiDddVO5Vjfs4Sm5L7yODj4j4aoAlDfVbOhkipjg6zZg4t1C4Gc3ckqxt3igU08z
G98D9hEyq6ybFtpi3Bd2lSSDhcQDQW58lDMmv3f8V5BBX7pqeWMwMYOKgg19+Bgw3vSF/cEUFMJk
np1RzxyDq7qsToh8gHZWSImfuzHKOQHFuvRhuYE3oY0lIuUtgb5Q/OMyYGBX7S+XwmGWk7xFiaFh
aLP/JQ1DAzOg0CgYSJbs7V2flHz/vsL+cbtH4Yt8aKQCe5Jrkgujc7NpBAdU/s23tNYCYIIRq7K5
zdVVEbEwA5UzC13buR2DOlsCE0xM9CoZ5PrvepPudHt5CzAvbX3RsgvWopSryWhQMYTFyyQEbzXS
0UNTfOc5hQGHT0ZMmWWp9ecXGmLf8L56RJAeypkEa0SmnfS6RyLsLzNw08H0B3MEtUdBS5BZd6wJ
zTo5JEtS04zdT1gr2xHokEVHCKNuYsHuAEnnAnImfILc6t2fgcpVLkKSgYNxON4ujGyMZ4S6s4gc
3qyzJ1mnfU2gw7qqt93s4J8InWjWmqzH/R4D470VMMpNrHQ2j354wx32xZwsgv5ObIAU0xFDAp2e
qubVHJrRlOprbieTc+SLX7+0xXQeIVop/5099K2QQU0+HEJ3Jwqaz7K1xybXiMWHNfFsidegP9Kj
amS/ikc0GGsYThdK/MU7l5rfGzEmRpVVns5I+IlIggBFgwKttgxlNajcgErAcBYWUBqwswEPIvka
a+jjdBzBO3fsn+IIwxn4CftQd+2VaoqmZ3+YNRR3IVFag+4NTUcx0j2+tuF1QoBXr70FR4HTvMXF
51/9sI50rRKv/VW0nzdS53OkX3fWO/krzJyDUtytKTTLzLg70OZSMmaCHqmXJOc9yxTYYPFfAVhi
DrEGWjVoeexOfhuf9SrXUeHVXkNyEPNwrDQCOCttSXWMNSg+XIAJuGZP04x1NMH6/OcH24+J4Qg2
BcGroQ8EQ49PGo+AQtT671IASsq4Ft2k7DKKVzs3bdxMVmHbHhLGYTThamh1YWxyV7CoZyZAffPV
jhQ226GDd3/WzO2Ot50tOII3Ypa1l4Pdk9Kiy5JZwwNaRzQ1rfmWYmb5OHcD0v3SZ9oitREdDUsY
FikVFNHohofSqaOEDtAlNrWrZP7E8HlRvlNHy73MhOodDm2DQLb6olEW8Q2O26MBNblzBScu40tz
QjdFG15g4xZ9qzTd+/gJnSbVR2mM7z6hQqQ82sLRQWvlnB/wPGzGsM8fUcuQTnIhpdrAZ4MbpGb+
kiB8u0rTORo3ip92Qgf9e/3z+3lCE9Fa1oxRAWOtuYlU+R4uy5vOtceGS1eKSpNgUJV/3yezsWkI
z0lOidgNQMuZwsgftJ35OKSni07VgbuZEnsWZtCT+7qIcC/wAjkvDYATY3gcUuDbIQTlFy3pr5Kl
nRifuuTcGaoN+bzseQCICo0kYlgellP3ckVL98rkp4S6LQb2KtLWzuLuQotOlhh9Ybm68Taf+1EX
ncHprTcgMYi3oZ/jg1umxp7MgEueTpzE55PoaWSbe63eTeXoE1VT+12wZkz6n5h6/zw+C23Ei/ew
VzAZKKGfoPfQflC2AhZyKD4wlhh4C8o7+Zi+Bn1X5t6Wm+CcCnwIaUjxF5HDRl78+CW9/BIdqhZe
d/KAbV++VdsCw9yIHmMAnrLxEEi8Bqw4FNc6jIBdS0BIkxeHySz/ljws5a8/DNVUwQmMwTW4DGmF
vVn8eyr/ei/XMQNlYdgjZkZcjM8Sonqa5oBAlleg8c70jKz69WT1fY5TMhbQPsjPBaMHalxqKw2i
cINq7zXDpxanBdLas0utNpkkD1zEU6JmVXpp+AVJxsK2fMyE742h+iAJhG51oamDMMBBLr/+UaEx
+dRH5Lb7M69KBLNBsTrmTLojuxqecvhArrb0qu6hYBXj698yh9novv/dVeedlSpq7/v0cZm7IBH3
kRpowyIuLZzO573smlmldz1uFfXwqYPS+yJJEeDYf26kp0AOWd2Wyw3vIPzwuMw2N7nLHBOPPvhv
ZftlBsKBzYMYVNpLZ/oVbkJafF2gm05ImPTgMkGvWZhpeyqvcH5Ujhdu7SuH8sX9H9mDWUEiYohm
YJLmS6Gc+HsUCpB2wYkMvii2pAiEGGgEexe/YDEAOGeBLVWjVSF8tfSa7+dNCMac/ysqMIxmEa0q
4PDP+hJ4Z8wmfefVqu+RAFkzcneT++IAFqGjcFPDu6FZFTACaArbkOKN06CNWyVdwGjPbgjqCdjR
9rlhJaybPaWizKWpIz6urKWb5AXFylvnuam9UHkWOFXY64/0Gvlx0aXEtgaQwaGpcqZb/CCoey1L
rVFhqe/cJZvaKvCemIc4gEki2/9DsoMA5ahQ+WQYWOrwLx6HQyXoC5yLREYJrvpsXECjfwujTmuI
IVOrVmVYLyCDUQo5jiYk66DHQNCNfm3JaHCJlb0teP4gmEa4VvLFg44g77N/sxiwnJscOBFOLSUY
E/R+l8PdLgLBR7s/nkdkPWNrE/2buprZm5uP5qGn56JbQhSF43WtpTzvfafCwe5jjxH1HEy3Bx1s
u2WrHEY43p05qUB+qpnd5jrnVe7cIncysRnkiZMdrXhR7Wr/p//2adVwpslqvV7/daaEHwJUVdOx
QwcKeLh4AFZMfoQYfkaNfyQk7A8XB+H0n91Gs4uLoL608mJM/tgS/uObkpQYDrHDpeZdHDB/jnzr
muzIl/O0fykNvp9yLzVNyJEaKTwNmMS6+1Qzgmmb8rsRY9B7IZPIvbanr7wXaZbsPLB+ylghgWWx
Q/aW852LtG0gyMWIwQdddgY/HWcyPy5F/rJu8RTnAZGNr/G/sI4wSDfy9UIQVhQ/CTiZkhjDdXnS
+HDtkhdlkIgi/mnx8AEdh3BMxvlzdzP9EgHRx1STCGTgMKnknAMXfPy20jFZJdBEiVcBKxraYKOz
f20KhX0nXshbULVI8Wc5tu9jN4CvL2q4vi7Af2FNZqRlYz4AaxlgDoHUF4FIgWW+VbAkJUI/9DQ8
Eh/jE/sNnCkhaQ8UZjLeQEvEweu7YLs/MHFYyYE2/t5x7WJgaTmM9LuZEnEuLbRZwz4ukUhSLjaT
3lxKhioLM7vaBer2oL7ELnbhR1w9l06N8Ktxi2Z3nIIWLXX2YRgQvPuQUw9kqHHekvaXrMYrFHUi
u6kVoDpWiS9LLpomuAPKaM9a3XPJtix7BSMrip6/7/rDg/kJmubDiE+EgqbmwzqnHjJC/y070Xdi
cb0DDHMcTIOczE5zLfIapVPzQYLe2iKeMjchpPOqIM5GFvtzDTSvHuNCtePxw7GzTsX3taMB1ayn
wUuBRYOHXVlagt1vRJ+izJFSYD00SlHCms6ii0bup6NIhD4AY5ap+dMAdVBjIK+boq+DYQxI0YRR
6Jzfl4HL18lpLNWLBlEvFnlLn9+y+sKAKwQrVdWynZ9SoJmHVCiYl0bKmHoRB5J8Y9M18s3Fi6AD
/v8vzNegCIvQJtnAMwyiQzXEMbzUlpt6UIjM3FYnjoSuuewTXZJVKRfRQbwfqcAy6JXj1Y9zz/fo
gxJw9NlT73DgRGuX0Oie/sJNlCaADbzxHQa9r0jsbsw+PpWgPWHILevpLGYP7BJEmFrfJ+7zym3u
ISUhYgt4CxV2Qj3ruI91VPlALh2fXA+6d1TjD5OzHAxzmHxFrgIkQHGglRNfb/FIDs3UwueTubad
ORpYKqLhF23bHloFqEy1owm0nlZTXCUUTyStfgOqFz4h17z1RllaulRsRX3D+tS5JodCVyqxtG/8
cXgmw2rykKjd5HycjS8J7IhNHrHCK/HwQ3e+Psu76v5KPoQWKucHaIGbGK5ZK4NWHZQYZlMvvgIX
uXT4O0Q4kl1KT+0C8roUCaCO7ej4Y8bbqo6qqZF9W7UxpSb5XAgHzEKcnUArluU5h4yejO0crDv+
4mfm4PpjyLWSm6xlfORNfpev3d589J2us949S+Eq7iP+zWPfhZYVj8+0tDqGZSu/o2WHFed3tB1H
Bw4L3Wa90+FMlKEQAoaqLXWMsWnbeDd1DQDlzBkFv5bCEXbI2O6L73GVOrUk+cQbBJTAqBE8t4Wn
CefDrEv6wb9Ml8AK2cyq3pa7qXc4X7UXO2yjK6PKT4gF3DBCZgdUg/k8SW2B9RBLNydTXV0za49l
p9nfgrQsO1quSm1KyRjx/UH9rt2avLq21RRRefAr0bLDd+SvioE618RGXOnZB/WHciovJ6OAMzRo
jHEkz6bkKvX5ytn81VWXUK2AQ1FJyM3xTfmT0O8a1DPaTIBKjehdVthHfTwxnOksWVgu21ivpeaa
if4qeLBGqnEcZr7FFw9ZKj9ldQpzaQSsDEXq6ON1HxX5jX5bELaasIPcazY1wjPX+GM+JNND3EV/
kUzYFUEps49kse3iVhpY1mpMjOVRzvlqV23W+HoNd9yv9rjXJdmoyZymjxE21XiG0zty9sJpAunF
u39dcs1w5e7kgUUfmqz5/2Uv3qLAIdIoJ3BMZUUDzDHhMitm25RpS0A08WiRkKXdIINEbxaFIG39
tJi+UNG9t4Ay0ztvtz3tzWtLQllPeJGvNacgMNZknHMig+HPQAIjCVq3mQpluHs36478lioXzKTC
1zQP7O+aiuwyW6KbgdEyiLPiZLIDz01BHaoNX6qAjnja6TOZBk8Zg0bu6wy/1noJ7jyCvhuzM9dP
ptLhIHTx+xSMteh8/z3ixLz0tbn2QkD4ELAPUtLTrZ8QKIRy5GAGdJ2yRpmbKdi5XN30Essw2CpE
5w6u6XCpywfXV+ellr2vXvyusjnalvPPI7H/st9w2wtgx3gCoE2MrLNDS/K8WI3oboua78IiC/dZ
Mo4Mnl/5tvLybRhgKKZDCOUTqN2SMQhMb7MK7bP04KsfB1abrTwdjE0pifWYoVf+AmtrY6wln2zC
wKdLDjewYpMJtnhXCdKBhnocD5L92ibVqPLdivBjyO+wfJ3YbCy0cC7C1UGYXAz4iniixVzuyPk5
axPjMD9ZBR7zSOOYpTHRLFnYO9gVWeIABlnc/TSDeTeeuN7YR+Z7VXpnlJH8TvAx1j7CzeJKBRFG
P5jW7sCzfQOVHMDmjvHbQ0pI/bsQu3P6m3QgVczy17Z4Z1DtR7j+o8StdtZzzzNutyU5D97+/WkZ
h0b79Q/F2485fHbs/P6ELn34GOui7pj7dvha+HhpPKpRyPkPuFIDzMVoty6NrZDrSfnWijr0k77o
Q/3q+beq7WGGi0dbA3p74BNSgGC+6NMV522hBYGwpI24BMoDbiaCFqzoUsmiQaNM80fb04bprEVz
1hRDapwUteYy7emIeUg3adZfDzDFBCpOb08IF2NxCRFrSexmzTDxcHFuiWgqvB1sowicUU4iU36b
huMv4SaKDgIChPYnuWWidii/l76WRMp66Gi+90Lmy1wB2oEFbZF1lqj1aRUCpVRm/5+lxYijX3YI
btFO5+fdGbP9Y9znuCNxT2s36u6AQ9/hz76SNoZXcOp++776k+OT9I7kc4oidMFVfUXIjTae8zcF
12H+hMT4dGfEYZXnDjUJNIq9BKu4v2bqFH63xlXRbn6ECAPPflcI7DtErlL31nqtGeGnfM+/otJn
fABlZ/si765odsGFhapluH+en+Uvdraf2LXcBfef6h0kwvk76Klb6lJGgb1k8T+MZCCA8pAPgiOB
t3C8pANAH24ClveVvLRfmejnQZEMBvtkOYPTXhui0BhX8M7TrIYo/idGNvpA1Ecs4zwiLhQ7vv0D
affetOFzcR2RcRvLnv50Q78LnOFmhyMIqw8boLx2iMoF+1BVTx1X/U/Wi84fu7DV9TgrZKHTicKG
VUJOtnU3fQhLUrtY6fSg7WXkMazh1KQQCnDGHX9YELNlnIFswn13lK5o33VXiz47eqVbdl9CF+ur
jTET23ADD4iAUl1cTrrwGNFPJ6pIIM1jAfvupXtJgtIbpKMboZrfMYykLU3JABzVvjL69CP2hZjc
PpZMgvoVGhQeaFgQBNvB+CMgvCEBmujcVzZQ4gknCszza9bPFdbSCyYGP+mhlcVs0h3NwPUKfrf8
`protect end_protected
