-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
F8oSMGRSnv6WM3nXbonk5xdpU+YjKtHBgbhkG4zpcSnIPwev3kjXskTTS9jvDW3f
z1KtqUZOLfa4UghQ2hJZitZkbBJQOhGyQzoMTaR60801uj+Pzillff3BOFlSWSQG
O4YTXRXKwgvSEVWMJpua4FPQfigwxu/jMchyrYZCrVU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 2635)

`protect DATA_BLOCK
zRxdpaymTabXlGLS8fgzEYc7Fl0xUaeXjymCcXT1Tn4sBCMV3wKCKiRW6xDQ+z+C
OLMZHNJDt+7yTzPYOsLK2cHwsscSze2B2RggOzeGMiZmgRcv4P6Z4taL+7Sd7AJm
YZ2nZuyNLCngog/Cqo7xKo2Q9/b8deNj515M7s0819/hbQvvFI55rfqeAHcGDgRt
Be97sEstPs3924RpfuQHLkFB6QRwtxmLzLPM1IDQ2AfzyYysNzj7/pKqAZPlUL8p
bZxpy4dFhDSDeiPwVYZL+Sxx1zOERfjfjsZV0eZhZWba4WEOltuiQlLdA0ay2biz
ZepxeB1YatmwZ5DW4mSHSywcHJ+oPZz0Hiw0YATBNvKlkxBS2FWwSe9s7Mv5JVHv
hC6WY9jtVx7UNBCDXR0qM5LW3Y8pM2HikMgAz4ZuGovHkDTHrF8wJts3VwvZ9N3X
NV8QGKK1Je1vDax7PQjgcgKMzIzJNSx6Nkd7w8RlKNGi+3EBwf5AH1qYW1QkEt5A
Q/e0Huoz5iPRM0iirJejjRrZm+6klHbPlLx70NmOPAhYC3EauVQK1BAvr+JHxL4a
I5LcTZa4R4KcgLzJckZIQzwUReteRHJG0VZ8GCUeCcAgtZNW+3lxhaGoHWuLWifQ
k64UyiaELqPF8iFTRT1tF8X67ab74TYgEG8fFqzjpszqMzU+m5cho+/fGEzBVVMy
FTiFLTgBaVjb1NNL6bW1SIzQWVllkOGCR4X66N3uAyeAyvCqhZtV/E16CA3rlXeo
mEPpZ4TmOsdHKTX+cQtePWt/RkZ5+j5S5346wZeu/4NPNRQTh2URF/55rtZIvdO8
6h2OxRub49B2/EBa7WgDTiFHKt5B0IbuMWFFzmFaauPdr64qmxfdrOjWFXdbbQDQ
3l25xNkcD2aDCVnYETsUpsqEujcQbLQ871+Cu/yWM9wUFpQRBZj9YVog01l3vlGP
FTcmQvIu4LiKIMJ0zTwjUwu63ZvTsO3nt+znFuhBz+s82OUAEMlq+Qherh2lcplW
RMayRi6CR6enUXu+bpZ0pVyJ2LDKOyR25ydG3Yck8FNt+1x1Xyl0H+f9HO2pPh8A
keY55089B464HClzZOZ8LQszcXOl37IF1vaRRw/+enlDrZxp1QooA5ey/2eBb2Rt
TYJdsrcEoBi279wPGI9z4vn85qbJ12ZVLO+uAujRcthdtmNlDXY3pSPrJ7Yv+hwx
bfkn4ZAJ4r4nueB2VxklonNOaArazJrIVxzNtYkpdD3apFxeCec6s/shqOqKKgHN
ENLW1gHhqbWGDSLrO3YT8LvaQaNBT5sw2VZb7Bs/R4431srkOP2W5wY4WlVVK8YR
WEGFV86uGwgFQKwlYX8MvB1bf4kku2WrMmhLuTL6zAf49/CKcHvBmRBMgM8SiNBF
Mn/bEZ3DUicL1i2dkiguJLTWDOgTB3lSjMYw3dPSZBo5+R5JeK5AgqE3+82b0uAh
TMP18UPk3mRQEqi1Riey8kXMnEUu1k4QlyivACRjAb1nVTqLZ+e1OQF9D+rQxSC8
TM0yBnXDhtd/LpJ2sNIBcW0nsP6MbeUXeWpsN8jsAyp4JDF/J/RqRMT6rogaRVCb
pBuhZ0oBf2WimOLpIUG/1tZzeSze0fN9/N9Mrjc7I9oiZNLPEo9EzwNXf2hSqg2C
xmLuTeSb3ylBiojvD+9bgxBcqloEnhV/FV764TVki/hlXFOvyB0j60PKsuv586nx
PJ5c5jMK0gEoo+WO/pL6jsHy2HuknJfjKOAFOCp3D8CQUUjokxmGTgA2LkPRWLnP
oY00R1JwDV/eKEwM6KKkJ/QbCcO9uroxPsgvgpYY1vTdtHAGGMNiQlkiTRBIb0tX
k+7JlKqBjs/pdkZh47WRyR3jNwciOOlae0+pa10f3g7O9hy/Jlg0ykJg+1r/loEx
Wvi2LXeWY8+8kTMBpGU79VQkzsd9vZmYeIUF5iZAMqbb7//5fpCnv0a8p22c0DOh
iZLO1LXSdScLE9ZytYdmzSf8wx92dJ+5aUxlLrNJbvLwTIYM+RqQ2NfxE+HWabVA
kf/4KUX62oqS4WzvD+JQHgJj6uvJ9+3YC2/8WgzqaESjFiYtUIOvfy9vXSnp1Eqm
vz3ha1FI2VwgQrzZ11VJ4ihpLanMeRJgDUQjybZ37vkK8iBetg4nC4cP0FDvQqL2
dNBgYmK5+1UWkpwKIdbD7K6HlpCWd/zaE7sBxmjCHiWQBy2slBWC29YOMyUOaGP1
P20AIPsO8R8j0O3JRyNLvFs3aU2HvpfsWoRZMtQL6SZHE/vN1ck69E0nTfHZOpFQ
bsA4qigSC2Byy1RIy1SWr175zHWQFhs/pkm0/bYbgh7JaOBunHQuCnffllRzPVUk
SspvyxH8S4j4G4qmVl4PoO0PQXt+sP0N19LCZt3bkorfdH+V3sbtboje0b3bHCLg
MS9OlktTiPY2voXoSSAQTlZ7fJUIyOiMO9v03CTPBij8xQog9coEgOl08DN70BMZ
0x1JJALZtw8OEcLpU295QIUjIi9CqTe3yolJMZAIUg7tQ2StaPNn8RWdzgWyLdOt
Hf67ll9Lo7g6EpUhKYd4v2/9qpdciHS8PRVNkz/bWQHn3BoD6WpS1Y4VN9kWNC8h
xlgn4WDZ+uFFAbLGdu545AAH9fF/c3Cce2TvtMx3DiuvKHYCX/hl+o9QhB4UHLRY
WDjerGqryw7mkPXwmfzY9fKY+1gGHkDNfrw+YrvozZKffkNs/SELjvAXTav2ckvA
E4JWdAyeshx/wXkN3ofv4RiZu5vuGt6adPIEa6tNwcb5Jbmp7JcF8algRV2zk8KE
DBwTs+wF1GBraijq2rD1LI3YLq2F9YfA5BL8DPM97O6RsM8Wuyi6Gy7hJdvRIqn9
2Nf/tZjda55rJJ9ggwuP8Lrmi7WhsYJmWyZNyVs3ijH3PRq/SUA2CLpVCuPlG5a8
qmcQ1R/oFJ42RagoLymrJERgtNBPzJnW3ooc1pNEkkLS1QTQu/+ybJ/bgv/duvl8
k8ZnD4KGuBiaeVNVsKZDUn8sAY6DuefiWzUn+D5MNPNXWiibIDPVpz8h7OFs+1zS
FaV0KM7JiPSnDydB2rHTj6lyaByNEn/5wPxXlc+tNJbCPm6frFoFgX8xjx2w2fOF
3CYX4JAUW9h+e80pceUI7eo+bNbE+ekxc1TahD0599rzOgY2JW86DviM2GA34tMf
2SZX/HSWDW5kgbg9Lh0QwgUahkPK2m0hjqGnEdPPBYn66+arqvUMSGnomK7BYr2A
iDMhyABAIqv2C1qhTbmY0ZkdvbnsVTBqdgtybOrqglyDVKxOYKcuCtzEVNyiOuwa
K1R6pAKv3lEigEAHh61Db6HsO62tSxDJzM3YqoQnXWfY/ZZ9oJ9t9Z/ahRD9kvU8
oJxhpxuP4jaAUuBNBVOPsffx1MTDBizXBuh5gaZH52u7XNty6xMRj/+H2NzTrFu9
hZOG5/LShh67pIiiQ7EtrXf5E2hDqxhEnO6QGff8NI8ttYQInYXnWyAa1gOar09Q
64VMye3ORjXmZfXpK1Horw==
`protect END_PROTECTED