-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
wWZIQc9Xqk9+yuYouB53wqYNh2FqLSk7AvccsF5fo3WxSkXBnCdhPP4ewvJP4JNk
kzm7fFQFXMRTaRA+i6+lT9vgy59m9kdThMwBwiXm1Q+lXI3aim9QRAq/nieQtXq5
bYwtPCF6MjFvmSnUgeuzrIUNHEhzWn6Oc0ldeH5b63k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5632)
`protect data_block
t3uqM2I4wb7Wh56KjTrMBCuUfuG/CQBPl0VUKOcfjCzen9v9zG5NwibgqSToOWk8
zPZ+jGA9uMrCPpmK1A4S4E/qN33+3yxlnl0I2dPcUintIgrlDuGmKK8KYaohyPIn
vraPcnQ9+YtyXeSxRDiTCSOh2gEyTsLgI1vm1k9EYFnS/B1UgSzA0OPobGJM71Zr
6Yi/H1NI8TPnEEtL4X1Ij0dYfLQKWLGIyY7pu2tHWcYA7lcpV3d8qZnousphWwZB
KLOsB0WgGTHN/1wcU8/DrmSPQ/I+cO372lHggsaCR2V+siwOX3cS/pNw1NQZjyec
58xtVMZYIM654U9kcQPRLC1P0URZCuRq9cL62IOYldJt6Dav7FESSHkcJW83lV/i
31UKwEy2dWTJflD03EVC+dRUt9NyBPPqwdfv6kEDGxea1QP2DdOmUrR+AD7ciu4v
OtwUBzYNlMYLxzuio5mvFx2wO/TBYng9i7iioRL4yNJtdib0De7ugojYR7dQF8y/
akuFLch3cz78dqSfWQJoLQkBDnFk8Uzjqa3FieMN/UPoGKVw3R1CBAbhnqiEs4cv
tFCZNRw1XbJB/SWrvDJkA9kegMkqejVbdRHbt8Nk/ss6Urf5slFds5kENdPu7F23
qXM+KOjZsmtt5YZSzx7WaYSFHRvl1oPyZpWb2pfbjqjq6OzQCB8iC6bB9Iq6pgni
0evMNWzCLAUth1KznxKRTbi06rCd10bvYXxzpt270+rgxajOCO+dr/9pHNvVZDq5
zB1ORqgs9Rq6yoj3mJm8Uf2YwPLFqKU4H7c6M82RkThO/Y+gRKQTgKLxB9g6VOL4
sunxji7bGKCOpfaCwYXYA6xcxafL4UTo3TM0FN4bpd/p9wygSIKr1PmX0Vnn6WIo
axqkwr18QDSH+aNyDOSu7XLjQKR/eSkciny3hgbVoSJCiUHp8t4uFgxOtBShNM28
I2bqqHr+sQlCEPr2T10lbfZ0ayxpCGV+Vu11OF4W6DPWfhBtCAOG+JGg8eBMkDr2
L32/u21fVJiVRCyg+PIlvHuMcC574As7pp29dcLro4pW+mVKZYO/mnr+3mcuAQgS
a/73PjZqGqK+yEBQPw0PpIt/CIftp2f1jEfseVV0nGgg2qsoNU2bcPt5Jn1VCumw
VppwBBxG3SLt+3ck0qDmpnFSYCVtE7/FNRWGH+JXiRJ7y1VDE8zjChxTox+z0nc3
rrVrPzqCSG8ysH7hyh+jBiwXHn/QOtCuGT8S55XEC5eS2DLrWwsO25ZJ84Ou1VMo
K7iW8CdWJHDRdMghdrtBn+P55KtZvipljE3s1S/hKQJ1l1wtYWKknnwCk8cg/Rn3
g0yfwpjygb0cd9RPMaOd0t2NujTMQ57GPGLA/NuSEmCp5/WtI3MebwziqYjkduSy
dfbP43PhSTfGWqG9htqaC+8KQTuv56a5KTtnS3ymwE1OEmFAXe+uMFOxtTt1EL1V
OOXS7w39S92L/CNQQ6daRuSUOyD8TGOYkBCpLOLoU4wXPSZPwJ4AmZmK8cdo4WB3
wmDn9yvDRvCSGk2WSMvwQv2GpFpC2WK2PzyN36D4QnHgC8tLUtaGEW1klb6WfX14
5Wcft+apk/0k9b7dg+teN7/+bYeHF5h/d3lkk7l2bk6fItIOKgwIQwSbhuJOw0uf
21jhMwUzst+1bZlsDBiodsQDRrMDPysh3B4QgUS48XOBzBtEwpTEnyRDPC+GLpqv
vKkLT5UL5LG+DgSN9oG8+WLvZMkXcBgBI5FVpRyX+FlhYPEqZO1Azyh76vVsb0dc
9OUpZ0bDCWp75nYO349p/gYhKFz1MdFMiSFI63saV9CaFJLZS6uhmNzhBYC6eM4q
uaSotMzTifCWJ9tocyTUlWx8yB7lByhXRbBfvg8xUTbpTKUMX2GRtUCAl/7WoiPV
vtoaJtRRGk7Ywrtq8+PatL0+D+mbXff8TbWQgPCOQqL4mUq/+KO5oKQgK+ppjajT
/iv6RekzRI65zebsdun4c4I23bVnDc2gTmX1dQ0vaML2MyF92RTlVpIAYJgUEoOe
Fhs/5E8/9ZDVtVzfT6g5wLn6FneEfQLtK9Hq5V0ByINwJkMQlEIPJsztYVN7a9Di
f15PFL3YAnsuPOAVHgetoX8EM85z257G8KYT77o/yeyr+LNJPk7j6E1eTd5Dc1vB
Wlq+VrtHvTUYzhNSsJaXPfMB1DEbrjm8IHCLhKEvR1dtpzI2I9adMEbwBlDMfSbz
r69HNuG30nxwVukl2Z1saDJBXqRKsYaPf2uUL76kK6WBg7BdqGIhHI5xiQtSWv3y
fJydrIa+95dbfOkPCzg7vfJWcJZ3eMlG3hC00kKTwwADmccMXXdc/1AwNnp6WdIY
oMikWUckUKR8X88JFsX+2eKud5xCqYKrhh2bXQTSG4Bilj0ytZPmdqPvDUXUkbnk
euZzLF0Q6+b2rY7Vtwg60UoginSQCdSc6viMFwbH4/FdMbYGHPy3Sx2Obwml2Z24
vMPpZbBGsmeFnoGmqSEi0oQyK6NwuEM9jidyLI8Rx38xhnH5ZEdK6pE5TwYmHvO0
lkXNtUvqrV4JwiKdMoV5izRgtuD1q/M/Kc54bv15yfWPV/FMbVLVdmc0elgL1BI1
9145Sn7CP4dTE6CDnoMsL8F+iuVYsqRG6DzM8yYe8d32cB2Eu22Ji9/IElLNNXTW
v5zkiD7IEUR/q8xtf6SyCrR6fOpX7MjFBy7IKmGj9HruzoMb5W+uDrLPIpElUPgg
xMltxUjbsJpBXBwknkN0SAUs3xmbpFvf93NQz2C/Z1xqWLm9j9F6773DqIoLs6zf
QCvWNqRPTA/aaVnbY81bBt7YBooG1i9zyWOhmh7yacWT2h/8Fa8M6Qg3Lubp+4Rh
tT0v2YXnHwfcYuXFjYjJ7R6EkOOS6MS44lE8lOma4LyRQSoggR7a0beAi7TFWIue
MbtE9wbzMojU8dvnQSsIyIDgrp+FTDfG2ibXYuXog5nzjCmXqCHlvDinlWI7Ha4w
uYRL0jKSEDVrw07FjqGgNC31WbnwvLOgu7EM5rN821/4Hr2BKL9oCUO1hSZPUhi4
vI2baBcCO2VVFVodbxOmvkEvgig7reuptmX2wqJm1Bj1wABeahDEG69vivlECsfy
ragqZjxumRbsbpFimMHhLytmImSXNkWkEETRUOb8h4OUIj4yfN3Nmf/FX6y9bEG+
SP2uBr7zoVx++DL0AoO7L0HkubV/8dNuZ4g9HdsJkLpMawojuNap+mVPe3fHQ46w
Kg5xhZI9d3H34fwNVI9tXnavVUBWG5ngNt+h1eDURySsf+iDDE3IZeZInkdFRDie
K1CfGS3fspXOtu3WmKhjBfcvZOminUfnJv4V5yAmkjAnVKAxHGwZ/HqiL7howJOs
/vREg74o0jW7ZBItC/6DVH0jAgY0tIX3tungas4m0JLMvPlFG/4gypO4VeuTU1Ye
T3QUPK7L9mubmXxvVBPmH4te8hCqN/8aAk6k7j6H0fEmCu29RO0/p9GhXQHCPUyk
BjVBpQcOv0ZFscRIoK2CVNLsAMkXXHtdMrFAzyAGxhDa5U0BFIf3IGWdur4eU4Vf
U4xR2KB5f93s5f9aY70rZZn9G9zESo4RWFI86ssttmmEsE/3gf4X+VKWLjmkXG9V
rcWVXIHRhEsrlA+q/17L4iy6S/N6cYjo2KAZ5dfbqQ4X1SG2Go3Ks2oTgJA/GEeK
VHWT4hhGgiuAkbBIp0F62qqFl4bFq/K44WIBQRo012E8oRvCDlh/vrbGSAkFcOTW
b6O9vPmjORvUHYJFCp4uzBaJPIqDDTmMn/6C2LmBwcB0n4q2VnEZ+56MijvyLv//
wpw/IvMDG3l5a4J4sH331RuqlTNA8uePi1exjw0f9RcbJE6+2BCZhc8pYcN3uSt+
U2JpvRW2qUWL7ODiUS+ESPFd0WvdQxH03zNqMYeMh9yFTLn6+gpmszyDLFoyIeQx
aLdDHqq0P8IM4ithEadJyXR+xkMXpg8c80bDrwcm6ZS5QWI8fdvhpsxsKiOW6ACF
oRDps/Wd3UBdJlbFrzTm+XptVk6uSDTWS1oaKnmhoqOxLVW+guCMd6qcN99SpktX
xRkfebD0EN0CJx6gjx1mrmKZEXuVvS4OO4PywCC+Muh9vkbdvRz2tO1Wrd01nGew
eUJyy1y2gguFycRMG823pB3vErRgNr77vevQxyj3u47UZQfdFtvxdfaxCsKG8D63
e78i4Dg9dOYI3J9x1q1vvTx+iul8O9NGnIAOkrEjGTQSSNDTG9rcdhQ3YYDyLMbX
kC/ae9/f74uzelOz2j5xNeGpqgWbZI//jsPYIhEVRtnECnk1s/ik6ijMn3fhVpS+
rZDRQVf7UxFXjfeHCLHXz9c4fJNX17shgB9ZmuWdFr7S1CpViTyN/9AF6DCNn43m
bWjENN2rCFSM2teXPxZAAcBvSMJrcLmR3BGbJE+eiItoDtylyE+qPJmngNDtBBjE
/0/qwpdcYq9xxgxzbEF12vPPKaKQiEGt8ou2lrLUF5DkzMuRDvNwKIEwE7gZotDd
HMssi32UV3FGYltRInJwAvx8XJc+fYsZg5u4tXt2gRxcMOTzFGKqgo9xF9Vl6EHk
A2NLar4CDosVvQzR6smHzmop/9qBL/eBeqfnd3Uzo9GV3ya5YRRsGVdvXv5qPn7L
/BY3pLORs1+hCsei56meKxHK7cfCC3ioC74dgu5s3Hmfc7BReg+5Mj/++BhCPtjt
Pl3hdjctKs5dwhUxnI4h0rAI38Mjf0ukqI1MsxDEQPk8wh0+coDXTENE9nRzN3ql
6y3ziskAuOLqA5lCH7P67ZlpYtJI/sNV34TVDR+eIu3s+jShBAsx6Vla9Bjj2HQg
ZdTPYg5jeap+zQsRUnKQbxNYJu0wiLmk2tmFPr5m3oap+1+sR16zyZCa7o2pM7YM
H5EJu7HGuhIIX5Fq+ck43viArr7qyyXw4PRirAjNkeHfmrZvml7ai8czR2KyEL/y
24WQ7SednwJp5Eci1E7yTE3PjYxf/91Ldwo+mnWJCU5gBYqsOj/qndKwTMsGmmy6
p5tLRA74i6FJbc3s3ApoAwaT8gTjK26hvkcmfMjaV5DX0097fCyCymTxHiw2xVll
Q7VTAV3i969iE6DqBN0onOKJBlh29IaEq+WDoqnPAdfYhQqDeuDVpk1joBJi+SNT
1e57lmv9N+dFDJl2OfRyJTyaDRlZ7VEQYmZa6t9e2zwPSXmQYaEPbqIMvjiK0EAz
AcWAjwhZN7AsEzg1avp7XxPbwE8U9wxIvb2rNyYhvDtJ2aZzSk9Ncs2g6mpit+rN
LbIrljTWJCoknz7Tihhl0Hj4nRRJ4Z2I9nF0mE2gYe5/o37vi25h6Tgf5bnYO0lT
pf1O+8Bb5IKFx+NIepPQDmXzdahIQXMYQzVWg8IdgTX1OmGqfPDPvKbltKfRwKXk
UhQgog5W4gZjfvtGlrYzAE+hNXGRLRcd2WpNbQ8sg423P7e4hyopfSzxAEihf78x
oBHeEvN217lT3spCT8yrICO/OfIviip0RUUGEiv4m/886lN4kIvIQzKv3QhAFiMb
qfztnFffgK4mMvy0zcA9lgsj9XGrTYLI3vyLK4r7V+3mWL7hjsVxZLjK/32ARnq0
+F1zaemKr70l2t+Ldka/1vXAgJzEWdq3MS3+M+PRFfsCozJhjIpqItAaxq6uAf/X
SB3NtfpqhX/0ILq1wjk5LcYdGwfITZ3aXkzz7joqIHaTJa8jJ/i1XzSKGSfBEh+H
41cSvtYLkIc5qZezVzBo/qZhtZVBfYlVk4THhpbjiJmhPdLcDr++X0tzBTc40fuh
wX2Wb9PHmaldZswMIcI4K2jQOlJdl/9mX9PUpio5lK5dgNkXkn3Npvm/gMhftU/+
CK1U6yKCJqVYq3uwD1aC1fr6ITh8MD+TSI0ZvRyP6YnnCGkGKotm9tMsLBhso3IZ
IK7neumTsE5yUG+PWyZhBAkmlPgf1zyjIJdhkson7vdaqxuKNo1qHr5xfJuBOBS/
KlPJH6OiNIlpYWXKrJiVCAfkuFx7FwrcFWaUUiXRtOClVCiG1W2zQIPgbmLizNLc
D5+K8BroxC37K0PyzTGb3pqoNXeQjk7dFzay3sbCrvzsNcoh4Wgip/zvKMjxRrW2
4x+DO7aogONYHhn+nlGB9CFS8iFlEzJLYjfPWHch6cUGLWc+nIJh6s9qR97EBGKv
vQ+Hw59GGb3+74GLDEKD1ZQBEdSO76IEe9vf33rIdSTnEzGNBlrwYxMHnBt1M0B7
uVfMgAPxUyF+2RFoRiggM4JC8SUcMd//JIw6ebOSPbU8RPhj6+HXx5nu7LalffiZ
6fP2zhsHPk8yblzBHXZ11t8/GxV/UQCgvWmB53Faf43c5MQABc0Tdn0+HP9CQpy3
Da8+oa1ums7k7JIecRYeaiAXBCJafbH6VEX2iWdfMPFVKTrQxq24IX5m3jsd9+yx
Qla+Fq0TLFE4oSV5LoUrDFyi7N2BQWSyIugPHtsoaGkOEHNW4gYp6ogTZLELRCfu
mSoXEAyae26XPWb0fvbkJK4lMrn1waRfXpoKXkQjEmMLRxptLiiuxdz0zq7cFOAe
5fo1Na98xOumTUintDpBx/xipEr5m9yR7cxQqcuupAmg+05JEk6RTXSgJAjlE5Ot
11D5l8//5mczWYVfRJPb9ZI1Mp+U9Q6n7Eezhr21OcAQodFKLYeNtMNnkdIHuF8I
D3WKzjtX/UNWOoYCHUNSZkDo7eYce4vvkG+p2OXfIwkWCwpHA+VRtLtDEIr4mYZ0
KP/eDdnqskgjDtFuStqUGWRt4KIIqQOB1YKDKmmYTomz6Tzaqs8+hxlkTj+GV3DX
uNY1BFNO+QvIyz6gX8jIv7PT4wUMeZ+nPBTwRMXQJ/Limp0urS5nJpXbxPhPAXna
mAHTYz5Tj998bkEz2mVM+z5xCleBGsYm/G7vKw3gVSBllGkrT/lI0xmOxu+BKNh/
2oldTu4gxc0+udW2yR6N0wlt3b85/fnKeZPN91aOpuNFEzbRcpBJTMyI3Ne2W/jf
mvrC7Y45D04OQz+evWj6ANdJNAAyoL19f8SfcHxCXM7/m2gyTjVq94r5jUgqI+Ia
sHtt+FTRMOTtyCcbIkqvzK7XM2lmq9akiLIErGbb0LnXzbW1LHd6M9fOMmwFgBqD
iVX9wcmVfU+oa/jdTz+allhImalYpnpbvue5w7OTv9iqogM7K5Yi3cQK6v+oleUB
EsHRnbR7YRyv+/Ajn6EBaXVF/XXJwh6jnI82SiPV2K9e8gWDlZmB0IxYj2jU3fw9
A2lq74ZQ3UymiKHZdTPg/Z78VsRVQ2sJZI/Ve08Ryk/Pay8o7zQU/AN1yZ6xcF31
hmNbuznkURJLgC21TiXlBEC+VEGLSwM5mHOSqa4v/pmpRCegJItWgXPb+J6i0WD5
B8H4MP1t3J7BbPYwQmbQWEigsSaiL87zfqWwbzKhqxeMKc/JQoUeGFLVQk8UDW+D
m80nD4okuOizD+V5jiKPaQ==
`protect end_protected
