-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ououH2/TZaOjgh1TNO28cnBiSYo1LCTf+Ql0EINWYvqIN0JrxeSxHTc6zzS/Z4+N
qHhLAzDnvSlJ9fShb/6DDVYkzHuGdh1REzwnEBkOtDEYzCAQBcW0J/hJn9yUQdzo
PgO76A/5W20igL+Uq6TkHSOgZ0rWQuyv6R7Odb+3SNb3/HOTdnm1ug==
--pragma protect end_key_block
--pragma protect digest_block
aOd/Wkr3OhyL3E5YugHqlr2nywE=
--pragma protect end_digest_block
--pragma protect data_block
Zi9pBFwCPEmf4Yws/l4eO+/kpFB+DZR26XXi/5DNq+aKLQJ0rob+cceIx7J/etXj
h3m7775laVWZtYGUuAAtuh0D8cJot4y4iKm8OXdbuHeWGy4TnGAhdHgUlniWdO68
FNy13MDZ17iNALHtzj3jhAVTKzfpXQOhgcxCwxFTCNc20cPyJ4JCbvL6N23CW1vd
EJSLy6md/VGRMt+dICJZyrUtKFbeOqtCQtArvY/cydk26NIxoSpml07IV/msed1N
UJwEEf2ezOIuVwX6e0RO43WvrrjyRznF41qwpbhRvsKaoZj9hbXHBqHtt0W8DA33
1LnCr6eBKuP1utokpnPn6UXzxiIpdlTjgBN+Vwl5N0oZ+7IgrKVTQHM8tQW4ErbV
ED4+dcLx7VYd+Oyh1cpk1Me/xJWkiUtvd9R0m698iVcb0gexzzsNKwhF4LS7O1V8
JnZD6redj3aBA31CPm6pfj8P7MDUZXud8UCXBkuSnu6ZPaa7zygVXLL7FGW93Ddk
5/hZfAXLuxh4fXxvWXRYxVUM3n7GZThMOBNiKMzOifqKsNN/NS9FXbrWrUYa325q
93wuyxI5lp0twFYPZeT0DcSkw3H+DUCM11Du0JfE4ozJrnK6D6i8Z0o/MSJ5yX3x
S/rQDKSXfuIEZT/hqCLiwj3PuLrTfoyFjmtbKfTBxZCO2hXv0hGBEKZd8RjH4anp
FD1WzksjZ/gonLmu+AQSzeYsF+S1KEgGCvsxTeUNgv8i6DgHMAboOi1A6cTFXTez
oz46iPfjGh1I8Sel3UnGl4vRUypfW/oz5/SArprmZFd+Lwr+1keNSuc61GC9krSO
jMTuHKTJ8D1R3KfzqPOvG5e8epeb9206ikWPL/8fjBsb/e7gD6IFXRfqw6KpxySH
bPv2HhvgqL7/FycyeGcwWQyjyv2O1/wvEwN71LfCLwbLyi3qHtPQFLPjdJMRIlRU
63Jj9/5A+c0JB9yZUOqSH74FePUnuxT1/NXqehPyIFYOIoCos7KDWLGSWNgTlCiZ
dmSf6xLO04uxpWeNVWzydKgbBAshlpkaO4LcL2UyjYi9NhfxX0tEeiEpsiMMopbV
XHHPC1JB+0ao2zfdZq9ePPTqb4X1Wv87R7HIKDbGjMsjd+hjtdC7dAZBiRfj1rmr
74lNuhlRfjUIgToxnd6AN+8vdrg90feOpmjQ2frxUr1tWrS4ABgxEA/9v64VcP2R
mwtubWB147+ru3zM7c8HL3BTdqfBS4eRFVYQJDXRnD7d0P7Y76ATsd6Ot6pvxaKW
Jxcc3UVs4jnBTUgW4xvgMpOcGmr89G2cwsxVTLucO+jC+mE3DYSIjMVY7wRHWiMF
DoMuf85lI5GMcO19cqFq47LwL/mTeWyZd4RVOzF/2BmT1MVDPrmbYoDvUjxi2GL8
qnvwFQN8DvQjMKJTwWiUQ51Zog4G2/ZmQNhthYeRJgxt85JT97qLr4HdgmZ6tIWE
vxMWisUhr9PgTJpdTVFLe3PGYNpnffeyEiLDKHBbIfFrVMATGjdAEKYteb/pJy8/
KjRX9Svjz763Yad0wk42JeK+NFkjSFCUOmhWpP0Qw18JOJ6AAScU7BL8FGmbKSr0
jYavfE+st9I/j0D/A/nJZBkX3lEHy2KsMg3YScTRZ3V7maZLsi2f8/K+43GFGcGI
hjlPfLAzmC2iZlRJyCpkp9H6uMAGhMXf9CyFE7nDltMmlQsFGSNRNMdip+/+NvJ1
VBmIXaf3ok6Z09TLyC3/xmGCcARtU/c1x1CMCOIUMV8qCvZ67AKVevxcK5fLhgFl
ivN7uxCFQHape/Pe1OP8WomIREyqtwGVEmcoq/6fQov4ciOCVRpskVlVw3FhnMoi
C86UcjCIcOdNkl7kkkUGoqV8m8v0AJMgwHCp1vOtZxCPepYp0Qgxjjm+MizZw2Cn
Pf44zXLgnVRd+8J19OUXnZL3JjETw/G06bRiLnjBxhoakhvivI9Vhurq6YWFQpiy
1ZXemZkIury9ivGXz7t8rV2Jyw0Q8NqgLhxgioDhZDp1UoDIZz9yRgbCvkRSkzPL
Sruk7LpZLjmNxGjzd064nHHZkIyrtOUXSm8zZF1RE+3Km7BVrd3Av9hBMJeFYJeW
sjewb/7ZvzydowFiObOn67mY8AfvF+M5oRhpjcenWTDRR4b9RgjODyVW4s4t12MD
NLJjuYlGrL/p2zGSE1aJ8snGBhb8ZHj+z6TRxYS0oOgy1XCuEMe9ds539Y+Tqswf
VudCiCiNYTi4KL/nZcCyaazHlnQbRGyeQKgRo6PWUrruYGf6N0bvugVqZXJvXmEX
uBPo8HGJLm12+5JLyry2s8JBSzHjJftY31BkldkjUihg2gm0WNe5kmgGfesVDOwM
BqFRJQ8O/hUoqTiIwdUEL+TIlSs/m7saNam5iaVhFeSfSyzW2dSGNylS0h/5sPI8
JT4NTWBAyUXqRPaMgelEepwIgeT1m9gi0b6eJ9J/QN3RPAXBepn0sLnGkjK6v1ks
F6D+OfKaBynFUMgemOZqC3ogzHFN7yJ6bW4FbXjDxIBa++UyJ7kbh7oHzGu2E/Dg
E20fM0GTmMKlGbaj1TtDk2lY6hGl+8xdSPvga+elHqCztYc0GCh5rrtbysEbnPan
sMtGfBoKE5KtJJGb3wY4BidqaaAvmLPP+uST1MvBQxlVTa1HqFOZo4gbhtDqVH2N
plEx6n+mCQ9l5je5RCTgy7tMbpHUYgdQCSAbDUBtptHlSPsCQOHRUWdsu5qdJRL8
64RPp5OIZrH5XyI/ML1l+sCFH6iVoPdwyvS6Ab38VqmCNnK7SSiE8q/5V/VboYZz
HeBiM7OUewrNVxZTu5Qr78Kv18sk3kFl1FniZ8dmBMWqr3f03/Mhe7J13DZSExc1
eetnfJ+mBgVBYFc+kBvx8d96xjv7XEiuOfofxoNTZcVSa+M0hGgWZ4gQZ4U+L4ei
cH5EsmjZdBm35E/GtzJN3Qxh3EAuD1tk+wA7QuTfomWRluk0Jf57PvQ3Njh67kx/
4L0qHs1WJ+pH3yYecv3STa6GEzM6MTYmGR1I/VzPBBO58EZkcn3jcaCGsZAAWpoI
sld5ttS+pgwhCyemfSLUblMLQz69pnEPHv4u7AIB3R3z1qPQto82HfFaOOJjgxH8
ugy9KW64O7X3kubDSYga//BCHgjtDB8tkSRu01NRgcpASfVCvYBqc3nKF3RgrdH4
/FhuUccbVoWrKjoOAXKj7cmEeqvYM7DrcHE7G7Up/UTsrwn5RaxYLI7Eoj4noUjk
x+wP+ltSGIX0YOuJ8YM+hFTa85Y74afanwQjiE6QAkKbgRxCF2G8Kov4D+7dbsJi
Eif9aubRJIOEAzC1eimExgPmFyXTZ4HYmTDckF+Mfl0N8sPyvqryKWUqzob/WHo0
kHRJc+dOv9cNDI13G8w5fh4mRWAZmkC1LW6Od+1+2pi9wu/BpNfkILRpu+fDLNjw
l4BTSKXI6G7jeDjvfh6Crmb4rJU5HEtLQx30Sg4blj7gbUnbOq8TEEettoFOJ+Fv
9UsubIk+y51RFAb1Uiivyb+46jC/TMIun3+90f3T53Tr2/ETatClMyhyDU9aW7fs
scxQLtFpLcvptkVOQWVHhPz3r5WvFuKOc2/HXMZ9IBy2vUd1+79ZtVUS8/4K/uSz
NYBzfCingZOL1WM3alfuGVFvofaGWrlfRkCIctPb+uAY7x+RhLxX18rac0CDHkgE
nyFM8PCqnN0P8hUhnn/GsK60eOq5k0VBc2qZflZHpzHGW6jdbS4sVdWE+WHEGdgR
XwSWsE+WhJsxw1FKYD4MCl18Ksa/DiEt00miHQg74j93wHHU9LlC131rykC0GoGl
IWq2Je/121aZ8mavOtFpUMxpQjBlcKoFdIA9bXg9tcfu7R12Su7xO66CFJKSXY1A
B1IaXLT6BabpPORlSfTqsHAnjrkFU9+zmY9DqOeTYqGkON1fI3vaUMYxfjwBpQJB
K4XT1cPH8MDCGB5pOpvJIizfPN1QnAWtixCW31NnfFddkQKfSOdg91trk9es/ERx
X6ZAqEBNuVd/6Dsjkv4aoZgb1ukeIq8N5EfR3RwNM5wyOPOvHNrz26HGE2sga81p
48dM7e3Ns2hhyR9gBzkprbjqVC2l7LoSn+dEWMVGWGxEUQQupE04cLYfaHiOQErU
1OvF60MH6mzDCdWreMucl5vS9S1hu/9BwJsNDfl/KL+iGDg+/AR2X6UxtIRJTEWb
lLMj5MgnTVhg7DA44PBquO/726fs5iw4OZZDzipE/gafrPd2SVes1m9uZiJZcMm5
4Kv9hCLEkbMJWPNK1mhiLCCYq0C3SjH0W5idS4pEk2D8cWrufyBVXNvr7ZoRbh9D
JWXxEaIGaAdrot7BnZR7U/9RNZhH9mgQ0gy0mKM3UfeJEvhTxNx6ip6ePkyTpfMp
Vh51PZRMQbEHVJhidaizO/ftkBUBwnHJOBhg8Qcusowd/R3qwKoftsEv9rK11AV3
cs+myhWAUGcM7fgZ31ECYQYXrM/dZ3Nx695qIt+3jeuFaL59PhUJU7ZneEbNjJOQ
w6YzqYyKWEEOOmddDxRecXUpxl6KppNnzKrbIlPBtAGpjlZBGPeNnF7CrdihoZ2u
ebjOdhrVBb1GXqrs/YjMwvfr3coLC1DrhmCYX/6IFBm9wRBLNvij8WUhuH2DtKe/
OwlfUTGJBzpeAAkb9r3fW6xLVxw53jgQZRZiZw1jYbXCJvJ10uExZ46H5W2dykAm
TOjwNaOWiwc8fbf5o230zBXFwgs7XGaSA8NSTzudxRCsQZOI7KVgewqFhxtQHsUh
16ukNkuIFZGY6+2ddp9fg32vsLuLNfHJnRqdseIWRAF9TOvKEIJb+9UOOOtQrPI2
oQ3V0Hiu6YBaYqENSWNiRsa2fFUkx29kpck/OsUCq60Z4wP/7f6QwfsC7gJiLIGA
mvefpAWRzR0xSXeWWi2TC8xQ5dH/xArvCnyOzS2gvDtanL2lfmT0g5EjEYTtMAJ4
0dvQYYa3+fRJPXZtSA8BKnjuygbi+MG69Fs0y4tg6oU4//M8Ksyfew3xvW54YDoS
4kGBz/XlgNTHbW7Z0CbCIPojBQGbN2DchnaYEIWinoeXELSWZAhx3H6zAZnqDYPZ
FL4TDCvG8cdNzzUg56sZmDjjNimtsKdilIXwib1k/1/0RffMhEhrLL8gxTe7hddS
Qc/DGo2QO8417wFAEZ/NAWks1FjDIk2JyIoHE1zlkF1MbKXwfh72D7ACvcdLRchG
9/ESruNel6K5WooECpfSmD4GuW7NQhAeae3vswKZVLy9bRiDNhf+PFBuRwynnx3m
XtHDD8KhlQEAhM6URiBTLqoYAq+VaaM3DMbIydXfjmh7ioWXMF08gVVzWY1Mg4YL
FuOpcKPIcYZpCoHW/kGetPlN0MaRhjXtTuNothLJj9lcbzXyhir2NZ3IdK6tWrcT
8piVxOTKnmoK8BSQqKJi/2peUIcEY9w2VOZ2wgJvpLWvfXcLQYQ/jLnOFLrkEMFq
QYNaegXjUwecbI0rnY/kVVCCEC9jQ4sIxRO+4MV7CKGAFiqrhn5on9kY1DF2TCz6
45qfHuup6FiYoLL2NpEFjhxuOjD1Jkbsjb553bt/Gn6p5pRx1dXoWLswxgjaeRT+
pJMfAKuZg8wG9HdaSjLQSFY8/B/7VWHMGaMUDKgGsmj/crJVwZZyno2ooDyf1f9X
p4WhLdoIaD835zG83yisENk68NTc7GNmuoU8h34xA0S+j6uVFR5rU1ECAGi7SCvk
LzXmQk8oabSpd98ptLaBo/eE2janS4w5yHEo98eNi1mD6u3um2T3M6p4GiWaJ1qG
KIhohfDe/x0iqe/rN5M5S8Sd6MFsCOJE+WPp/8eEex8Isyz4kwUefax7anAqlbYF
36BEk5yqNP7ud9UaLreF7H/mNIx8ZHCEEe08THFLyWI39zUbSPnn2bQGSM3aJC50
PjtQhFji/PWwQ1SwN9fAkisXb/FQvE3PdC2pGMeDvJ+M22dzwWXDZ4BTaHNh3Wgw
MFTMyEZOTBSRhHqWGAJNGDzAL/LfSs+S0tQlP4C+7pfasMSNT6HRzBCcF1Iudc1p
oyqOXQUmrKSF9F3xhLeeo2Ld2eT4ztqi/1CXEVAMuWW6Z9B3hkKoF2Fy2CXvyC2Y
XMvT94i3e7RvgG5UypaFBQvWqqb+4yrrHLqOMqEDkFGzhZMW1pJhxy6WoNn0Ulgk
nmEBs2yUaG3WpP6OYQ9VfzkhhvDkGVdWJeYQa6VwTzZfiV/aKr02GODyS4xBl3aA
yiy5YRO6M68SWUANrDls7J3xaaSJpiIBUo0mT7tg3gXGqLwFeH8eMsKq3MuCJaFo
LBEI30xjhjP5jbC2VeHJtmK4x5W+BAATkkCTB+2Ylh9Ab/D105kfSnDUAw52vCGe
YDGc1PtV8cK6qBHcKGxOhect2zE66pCCT2O6zMrduEDqLU8pANSfa0LKViEmJqgK
VW8tFsQCfttNsyPDL3/hTgA1/xFoub/Ic/sVttfSc41MXm+VKvOiEypFPE8FLm5I
L8TFdv2dUWI+GWPx77a4N+a2L3TYYGflUe/8I+wxise0o392NILvCAeEwL86cVFE
bN3DI+uRgHk6twpR4Q95SFL3ZDWgcRGn72+DjUPMLZNMvGy1iQ49IgSGpJfRRDdb
PFtI27pCs70cBBcaz2Jxm19xCjOCSqyINa2hdo4L9i3nGNudOe+O64vZcy3zvuFG
b33kkvXnXhAYjT5v0eJMxzzgt4u98oNmx1knXlRb7dwi4UDUJZU5hSibWMi4571V
XI7V6MVjGDExkVj8FVvXYlmXxCKiMQKl+HuH15RYIVDRnVcBxKXmXiRN9exIll6L
4A4s/CAEzhHOmhitxGWEkRt7bRlN/7FmfDcCVoKsD5MtDzIpUV0b/X961gN8AWVs
tO1ydO+19lKgqlMlJ0Gj391M5odnuyLfLv90j41k46gCnljgcnxl1EMLX61ylTnk
QHCK1hn/2pkSA4MkKciSqLxyl5g+YMC5+UYVzSAbEfi963bg+7SWz238JeYz1CHY
5DaVGmIqxq1wikgZjqmHUEJ4CgoraafBc4a8knHuMdftE/wKEaq06w4Yy0I99txm
v0gDFGVLo3k2HJnDc+z6YNFia3IPl1dYZJkoZNEbg+Z3TKiSyR4pwWSrjZiLUlO1
+qrFT17lK3lXs3CjIGuKGVZKQQLnI+dpCvMOftcHl4Kv5zhjdnb/7DcKtKYPyCwA
wgGOvVcSM97DcIHrzi6PPJ7B7VhTouIJ5RhXgcFkRKvY1C1L4aRGQWj+nw6Zvik+
Ova4vPiuyQoGhB6lIYT0g10zxOgJxRbdMhq/jnKQ3rfFHCzRUnJla3Dx5564i+rG
/XOPPY0i5YaTmcUCP3iJeU7y9wqs3br6pU6HEhwyx9MYJI8Lof+iUw0/Cm2+MGup
dnOGjyAYWgw8xhQRZ7VglucbWifqHHaHl94oVBC1DGKrQhyGvlV59IQAq+2QS/xO
i6yfNQU96tAaDoQMFsuO9NxOLpVtyG5tDnR7XSusApNfgirJi4w4oNiy3Lzuzo2f
X/6bQOpJepEZkNCKR382rqMkTftyTipjA04374M0qBtj2x8u/uSniFcsFUTMOP4y
s5BolANUvOEXtNDqiESVL0ZBZ0/VGgvlsHYvbpKLtJh3rWhzUK9EPhTOIuPcqM6U
pX4btxrhK1Hk8fnZZF8zKgPbSPYdKOJb/6E2e3o2FCjuhDbqafLK9NTsKDdqqeGu
1s9PZ13raQwNP76tCEZ5iseaywoJ69pMXv9wzUn0Y2apnfhQT/j3S0+QPyONO+Gz
lvCllvPq/yQD46u7e+7oS4JpNAFBMDUHK+bmyiVAt7NEVBhGhtBoCjBsV+dWGTeH
V3gVX11YhbdlkR0QBXMbrkVFq6EeMb9oU6W3wTBjmp/8MQrHGXQIySmP8F89USwI
aLJb3A0g5Jk460dR4kvUT7jSYjQoCa7fxNPQoUcwKLu/8fFrYd5JplmndByLS290
68EfjmVnvwHMbqJdFwMJupF24ej+8pAv64IoZkH5D9OiraIX9wTgSgzJN28FE1ms
EjcZSbvHSmZxB4TbvqvIftUJUrHxtdc7XpBhkpXvvysXo3gCpNigl9ZEaAOmJnoG
OTGcnGLnX7x3HM5c1+lvFN4VmwrAiBK096uaufVfn7Tuzcg+j0tpyfPahc+XQKxi
qB8ibu5nEQcbHW9gSw50d2uT9RL8Ay9q/W3Xpjb8MmvjJXmIAm9RLrDnjXMSk69E
TeT2HMwuaEQep87cZg9My0JdzoOQ50pkZtclcY/OrXYK6wkVU+Uv7bn2DUPJJgOA
z5zD4+0pbm2R79eQmyyOr+CSjmKz7tfPs6VAy/bPHxxcYKMoUW7rfe0GswwkJsGx

--pragma protect end_data_block
--pragma protect digest_block
RxWIIDNieVXT9kZ3/RAylcQimik=
--pragma protect end_digest_block
--pragma protect end_protected
