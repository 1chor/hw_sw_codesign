-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IZEU6Vd968+qbYRW/bYW4jyq1AH7gk4MZYzS8FoyRm+arBeo6VmuQVyJquQewkd2NtgYDUxeAqU3
AJr1qL7DQ0LX0XnVyJ6oezYjhh/dCwfi/0Fxg2xBcLMwiUuikrgD736OS8Uke4Ql7OvUDxci7YSi
oabg+pS/uXm/ynzYS5th69al6hvP3ZhHNLGGp/qS076dt2zNzf/DQLkC4XZDoKYRUZ2xaRqbE7Um
OjFDW8yBqCucsbTHJ0hLlHibrurJ8ZNgEQbzSff0XaUXuxig6p7hmb8+tKNF0tF3cbRs0ADJ6pAU
V010T5aNbwwE1nFOD7csyTfyiaJdzme3WUcbkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 29472)
`protect data_block
UfzyyQY7Fz/GkUleT4l6G8ePfgUQfoblI04aE7XQwTpQ27X3JWXeeulU7M2vJ2lZLfaF+3uTulXB
TkITr3x1rf77Hox573TxBxKzhQdcqdbcsH2hp1nOaWRKXDc+Ckg+TQK63ILWoOXp1yYR291IneUK
LBgZS0xBIqRopujrNcNCkoScyrFtOErAmUE6p9eyP6HQsUlzVT6+dKYNBbT+Q2AYARDOvV2Uta5I
zDsZgeYH1WLe0U7bb9FElFdFxh0z1G73ZAYzrVc2AFc9GXeZBXOdrUL+uIyVclxeR/AX4pNcRGGT
yltZKNMc+q8EX0s/74ZXQPAXSVoWYVyydLt+NC+27d3AniIiR4P5Qe+cVZUwssdrXZnNST4f8GkE
YVFxcLWKFuM8ZGgfRVXLOq9uDjOOAnSEvmElsgh4e+QU5zozFu3xqQh7GOEXNZOPGRoWxPC9xXXL
qiWak9194MSCV2y542IheG2t28RbbvJDr6vJ0AJZ3Hgcmu5fxGMWUmx7245h+6PnknG8EEe45rKG
ScHANAd8dbyYjy4D+pgBS4/VAE279SSpV2T+0JuhLH+WVcWjnSv2qPU/JWA37JVnIHS0TGolEn71
zG0srQNpn5uJbqOrl/2OjzCIJAibYnsKkicllF3qzsz+F3ZRfIQxw6X1k2JwHnXFwDhWsU7ml3w3
CkAocJHkSBe/Pg+n9NN/pXF2MS7UPqMFfwahfNuBac6vQGX+DKCGrc/6/UZRuBF62l/eunw4BZGI
+pm/2Q33E/q0npeHVGg89AuyWHY43IWEGq6zEW2tNPhpm6B86IcWl9pHJr7XmoiUr6dB6wIVn/PW
d/2XZGumH+68e/OwdC/8+doja3OQT+IY+B0KGS+qU6hoadohD7tRw2fbKDv3qmhj7fKiQoWZzxJD
0GpSZvMiQU4JbomnQn8hReX+rPpgqEASDNn3lyRxZyymXujs7/c7yoZUWmDSHNUSJYFprFJeyxpr
inUB6IfC7LqqVl0NvtYJcYKU7wvuYJzqfkDKiqSLOUzmeVutEOkaYDn5tUMJh3Qjop+snl+v30Mg
XLW9xY3AaJWUwACgX9jCBAaLNXTb4y32rzgTNZTxDm4wrgIg2hxcbXwKjG0mjmgtFxygXIGoSzQV
VBhpS9UfHWp9cIFfW5CyxyhU8r20F+1WcKfZ9ynIT/Y7EppxuOdmM5i4dg2dRyuLQvYsb9k2emId
dC9rGqtigMv7fnkcuBGGJDtIOVVZUZF6C9uWyS+DrzhhgXBd/vjBBWJqgdISe+yOjXYKVLSGSCiM
MFF6cvgD/YddI+fLnZeDhe0QD7O3Ut6NS3P3F6xB9pcII/xBCVfTCt9XoMaVf+wk90nNOug8q/Pf
wXg5LYWJl0woODYoVst9/mOF+8bwSU515K7OMqg1Xm6XvcyA37J8je55qPfozeO6/AtWiPaisQzE
tSLfCXs8QWuslhzMxDJtnrKJJUrfrz5nzSbbIZbNwYMzhwek8hEb9E4jI/7nlIIdtW0+N0DR4eTP
bKkrtAt8aC8vKeGFcSxYHJjBo5e4R+7MYWK5WWqwNHHSm+T3z9NKoP3WBLRy3TJp1KNR12nRGqQe
Yz/bnh2GHWUueBpD8B4GkNRKfLnjO3How3IKhTbF5GaOMErrBsTrPnQLpLE7N2kL0K7pFn79IP5i
LRJD0vPaPKK0d1s+xIqgW+e0MrdVxU0PrgBiy2Nnr8CkKL4zEDWsrjBggmv/rfwrE/iaNWKYes4b
dSeL/xi+Cc+Z5D4TrfnMwtXKz1pVc2DVskROqt/n8vESVCvqukmpshx1K5UiP5XpTATPaD3ffVff
IycvhZRAAs2xJ1sqU7Bvz6zvyg5nV0mx/YAHshXPUzMjTxXoITgCQegYlqP9wb/QFhNhKcQdcZx0
1zXySeCM7BM7zz6aoclZHdQ+LnT0AvKZtatlM5C3NUFLzN0mbDKc0tuHqVxYMLk4dtqwfjSFQJgl
vyevLKGPnFUJFoLSBZ6v36DzTFjf+1h/L4w7FFDOHLcPl0/8sbayTqwuMmhhGvpp8cOkbKcfTmmo
HkQp+4M8rg8OHpfx8RwLePqpz8cMliZ4bVqWZ9sLaf3JQWnqTbxjr1a7loQGeizq01qzHB+Q42TB
B0TU/iRQFH/ciA5/8JyxEgYPh8tz8fmq58lBDGRGFWkof51PBHnUTRyVpkDpbeSuFMc/StQhPEWe
eVRB4rfrl1A+Zybc+AOO3DW03CrmVmYAgBucQO3qPCBnxvgT6w6mqqbf/M+iS9q9lAvcq/+o4nTG
okmtbVsJK4pKd23gpLxzv4G2tSAnLJBLtOaqsC2CrxpZ0KXbeK8WcEFaxhYGzREOHtawQFokUBXP
8aYbIaUcU9GwLYmKQdOEaru0IMpXmfZCSJVddJdXqx2vj9PyEIWRvXq0ABF4Le5CE9A11wYC7OkR
4KjheCPKn8ji+aS/9cGKVGH4zSXis/sZS3JyaTUiZldqs2hk7W6rUO5/nK5VRgD0w2SBe0ZQNxLF
gOEHELbW/QoPLFLKeMoFBptwl0doz4lYLTuMnn3KjiTjNO4ZfbQNoRPs57PlSfqOQqat2Qo/UBXv
0bg4wuWGTbNqZrH4xY7Hj5+gKMx6Tu6OxUJZvWGx9IQRDYfuA/BedkqFXRggvOZtv5APrRsh10dT
uhayhJykQT5k13yaT7+koUUdZ5D/xMN3G3c/gZEB0PaWwdUhzthpvXYIlFMGgaK6HY/UOga2nPkp
7Qx/6x4MCofJN31JfVZb5LJxYHUZ5Bt/ExTHkuIxY+4q8nHZSEP4We51VJ7z/StMcyGpzMI61chi
n7aJwPlx1jACyLLiekgngXUOw2ZCQ5iyQ+uByRZJG98CxFYxCn+nwewitrOFb29CXYlHtU08X3Ps
tAQZPzbz3iZMJsOMqXgnaWGVqK9En8vWuF7Tq7c0JRC8DpHNUjEH6YFGlWNsca7c54ez4EoHrQ+C
gLCzMYVHFsPIavlY00kfiAaEys6IM8QLIwH/1UXSer3kBwDB4ICdEYNEkf2PWIpziMkcclTZkI9k
2c6dXiAtlGpPo5Q2C4p049O9Jnpb4AD98NmUJ/oRrNevvSAjzqz+1/C4xi5Prw8FPfLIVMU7Mfx7
Hw6a+noFG5EofA/lzQJNVvyVWm05q5Rc9WZr4TFUo/S1HeqyvMj43Ak2UZiyPQHKaPTVTBHRqOyo
09VmVNO5tXW5TEsNZIzTBZl7MrrYfXW3ue2/Tz3SakkvBsN0wRkbaengQek2U6R/MWxvqmmCYadm
h9XcYS7LMNHJ3XqY5tRfQ0yK3syI7cb2rLGR4+f21WVdhyvahkzSBljbMaoP0BXlsc020iNhQ42D
9RZtYllWOvKoAUTcfqOgouck4ZYcn9EPmqLJqI1IOak9C6UH98o3oIB+jir/j9DqM01k3sty9jQA
q1theB836fu8iTHxiVFyTYSZY5ad7nEWWQOZuB01oQ0IdWOkSka/a8GcqnA2f97cMzacjEakRKMn
IQAhFoFr/qHTRY7Yj/83kWHw4OwCwAIADsz3q+0NQk76KtXQgAycbJrcXQeb43VJBAnUmMwSUMco
X4Brs3b1Jwi4ugrVVevE2IcxDFkvUoJlrpfNewtMsLuhB7zPgO3I0G/Gm17eWvKmY/jtkeuXpb5S
OKbiqH+dBb3bqM9YArCmBiskYJxVVuWvcSbdjzSq0iq+mRMkTNct1pf+2av3/tUvU5IcXCYU27Lt
/RbNwoN30gRrpSKsYcVIqhWLza9TTXud4NAhCGV4sniSGuoAEJT1Cu/uu96P/wcRVQCRY9X/Qrui
/irbkm0XRKLJnjvcXCfy0zaNLBuS9RzATOuQjbKZ33JoGJ9ZOsmY2tItVL6gNeXYuBWphcmy45zg
9YSThosE3DZ65z9WLA7USAQ6+rXwE37QVzEWNFKQV/hRf1peU93ZzdWqMq97/a0ZtkdPofCikN6D
WOlOEQJ+tZ8ISBeEw/EMxZLot54inGsT1DDcrT1fco1tj8o30g6JOitPeScNSyd4C69tdOhM/vKQ
k/EoNa50krtusOQgQSrIogAgNP+oNa0t5JmS0e5Dzvtk8wpU3t6BLsNnbA/AfuLOub2F3KR+UuTs
Nsdw0H4Cw4GqmhxiTb+6stKmnKYmChCPFGp0cukzzKsGmG71pm5x1tExe8w78mS3b5Thfv9ppX3G
eDzQ7lLF6rTlvJJPwm3o3JTgu0Qbs1tYXn5qDOUIOzaePGfqinWUFHoHPEXbiossBDpSmMeySrda
YgviXikRoE8BrjWneLcmOnLsV8dIxk7zp8j8Nur3DeH6VFgYxCCmeYyzfTK1qL0aRh4lx8LFgIfS
GMN+YAakIa4LjlerJ6AL2dlKArZnSPD1WcllnCUH9HXXNbyxEHuJczkaAZnjSCBnN1Z1qavm3O5j
51G6bVIjlL1wiuTelFbQfG5g0qaH/Vq93/MfCuXfodXCyhrchIkPz93cmEWd0MZoHSHRjnEZ/vIv
I+CtiQ9d1fEEzgSTyTbFGoubNIHiYalK4zBDe6qpU32w2JVKjLodccWsgGA/00MJFhZfq9ronApA
VZXteEFlRIX2vwUuyuZEsYClraLEa8Pg57OoTKDQOFapJpo/8bIEVNRuV7YLE5t+O81/tIfdaep0
Tte/YD51lEjTXwDkr9zIz8h7ogEnAbS3F5vNUdaunz5Ut1vBH/T/DPh0jJhjQ93FyUfYuM5ZZQXt
SOeDyTOwIK7wew5Tr9PRGtGFTegQdHmShmjM9cvRjwOoTPSw6WbDcs3l6T7hNkuH0FaSdt3NkTS8
3iW5kZij/fvnlpp/dM/I0IHrSOn4WOUo80mz0nriqi90F9b2i8RueFtCSmCahtWEPYrmzKNoocVH
r00CX0OyCuz4PRYEz8NUYIQt+/vYe+XbE60bz3Q2vOcPNzxz1kRifkNv1ORhN1pshCejXC5Ahvdb
H9/Xjwe9rw0sQDYUZSZfKZCOjz8XjHHFFAdLX3uKwqZc8eKjF6kil/LKYr4h2mpB2p+Otcfl2oyS
DGIm203bEJC1UMsI1nbyG7/v7O/UOFanaV/ylIDtcVmg/P479bNdHQCl5QG1L/chnP7i2WNRmLU2
Fw6Y5gQcy2pX99/NgVpYugFMuCNx0C4YOYpQf+UnViLBSsIjzegKibJ+IZ6Gr2Hl1Tqrvub/c9a5
GQ5FVtr+n+ufcaBlYD/W1efLDxOWAaJDkeJHoaNml6/ndmP6v67vU19iJkBj/sBB5F0PRKFkQYWQ
F1FBhqpzbtfpf0J62YNOKTYWq8LT9Ku70ibBOSceMm6EYf2zM7ZoDis2UwsSLOmtDmE0dfZiqbE+
6Q0Ya6JmI24rT5CD6YiS1FSjDyl4Oo9oUM3ZNYE+MxqIU5uVOHcy6Fe239LnJEJNL1PVn+wo50g1
1IkidlPDS4YfbG5ZJxpBzqU+LlglGMySpdJgk4uT888KkZQrDMb3eMhfZwPtCUPFPhv3YbWt3Lsa
ohuFukP0+5PSHPsHsDLVH7ufiPfeIFRiv6FHyVImxX+w/4QQSZSw6odSwiibJwKePMy1jNvaSRTn
Q/7wmRNheC76NGZULw4bUlck+lofmNuZLfwNzp8xMavF2uVtg5qZ7sQR9YvVZEwY+n60nnHtVhAk
8sYyeg94FSZx//D8wVKbU4FpULt3XBIXHo2cEP/FaB048FBO+xinxK41w4J7A3uk524WetjxPtrL
ziyNznVm1HfkIT92Q9+KaqC6y9e3kHwVkCDgIq0Sq2kvBrYrhs8Oe12K3KCm9ht3ONX0PHq7SBCQ
Xp9xlPSrVIKIzBoioRaf9VK40GPd5THlmQxSoGPH2FlmGHlDUT4b3K5hjOXpg3pFvRAoOR37BZG4
3ThSm2nroMDs+Yuosig3vxsMeJgJCpV0PJbLOA9jPOEFN2t15f88eW5td3jsjGc38LtcxaBBHYAI
VUIM4ojXubNX1EJWJRnhxAucYea6U1glCL7czEJolGbNC1qeBBRR9u0e3k+X4uy/e0e88D2YL8fk
06O57TFP9nazvbnsB5ZI3c2Ih1Ut+kYB0QEF0Z6hC97NFjamb3l2aYGBEG9kHlKdTN6W0oEr4bon
3fFjGguFxfApbkfpXhU8UzmMzY1fVpYwu7P1fRkiNcWBZu8qnf6BsBtEC7duy8iiNLqwsjG715sA
Fm74mHht1C1sRInYsoLh931Vx6fFkDXMiCqKvlNcLcaEAVcAPwMW+oj0/j75l+gLyF62TwZAad6j
ElNGs+k9ANREuDSuqU996MQO2SKtYwUKiyXMxyyirNCz7bN9yuhS2FQS+m20PJ6NuwRIjGEPuVLA
yEIc7FZMQk/eu9uEi5ldlBeI5Nmwe7glXs4/KXIzdC4BsZ9irKCbGo83N/fdIY09yF+vCtYGPCED
m4o62M/U3mSPleYmYpNUB0m6JOreMTMNXXF8TYDSwfIXTPGqHbqrjdT1AlclXxMw4NIMKapmxvEN
DkeqDe8XfBEzPlpTybhBY/zmyF5tQEdAGQVDvMNZCrR9ISBj6+YHf/NkX0aWMatmygO0Z8D7+6e6
B4k2BXkKx5YGIUhVWj6CszqoC7N52SIl88Pi2TFp93OpHVbKdCNWrmjr9aDsHnCcnx3+GP73b6xV
CaJyCUJqgFnSWKKwe8IjxXVpGc2wHwLDFRp0+Lb4BWv1AacFSErQZkxb4ABuixaj0VC7XmVwBg/y
p7xGeexQaQ/tLajXsQZZF0BK2aMRka+TtUDVn8BcSiDUXWhAfA4asJFYl4ddSJdp/sUq3F8YNeAt
aSa3D+yJVKm8R/d+VlTndBYBNjEzu9Dh07CkS7+qJktcfLMZcIdip99/TgFQXlSMsZEg2z2kSy9s
EO9Q4RnQIW229j8bMywEcmBOm9nZm0xWhPs8+hwdX3XyvYvG6aGIWvHLIUdvzL8HYQlRT+GbPzsP
YUyxmH4Gjf01KejAdtkNzKNcbyLpNUbiet7Sw59op2TBSceiLxe0XAzPxX4bl+JIACfsx0uQctQy
1EqGz3weL7lnq+IL01Kkbxwz+URu2ID2n+WK8cP6x0oP5RWqGFw8w9llDlFxS7deBN6UWhiVP6t1
j42L4e0J4wI4Q+5XDOxqzy8oxE4D4yylNgK9T6rNCnCD84o2cHt5IvZexBYcanmQlM0cdJEjWU8l
dRL+7c1GtR5yPsIJwSNIi5aKb8P+ZADT0PdMKbmL+OJMdo77FtK4kW5hhRudEA75stjnh4M8mD1b
yXbvtY/e1Q8kGPMj3/AhsZ7MuHodME9X9OsZVGDGAXvEq3DKOHPQ6vyY/0NyeJlGsVKKlG+sKll/
oh40uewiRTTMWy6HflpdrOLSHSmrDkP3LDhA8fsPmdMuHNU9JL7PPYsG19wHfmboMsNz61zJlcO6
CPQt16jFZLXJQTE0+X0zXkHaTbXAFf3WDLhhP6l8Bukj4MifuSovLB6et9cn79ws46vPQWqle7Jw
eFPgV8k5ArimUbg0Ag+BWSffuArpTjXY3bMm7iQxHt7avJVW1V8y6qHbM1Zow6QBt/qUqH30ZVEz
hNsQIUO4Pg0QoprjybAwJgRlYm6ZDyoZ58znRGf+ZNdPZvEWB3EuNEr3wlH+xtE9WCutpZ0l8XgZ
ZTob7JNwkla8uVWWF1kl3113juHfVEwgCxMIovIr0HU30dhYeuuiP4GiDjIadNvsYkd6xab/H6mj
8PGlZiTIhNvIA0MU5n3xZSp1M3v8Fn1mpuLm+HUezEWcvPK4bmP1ET7gx1YjPjUr2mbRM00NpOQ6
YNERro1E1G5Lkd3gakFtyg3L+U/1L+Z3hx3r2rphZp+TsTiJU7l58fcT0cv5i7B0oN2Bt4OTfHo+
CnXBpPmC1CtBgl3+U2Nl0TS/AA7gdUaZ687LMNJ5rPlsKB5w4Rf6PpFN1/F5pHio/xt8lTYKjRdu
/3/AoMxfVLcMVqPtzKg7Xx8hDDNXY0kCOKXyjYxrq4MRkwpK7/bozPOSYY6m8mJh2Ont/vIgs/hM
3FOyeXlleInTabU7YXda6nSVGtdHpVsmwLr2HyFrrUsCHpeVSJbziYPkq+LIcCyJNS6cXEab3BsM
rDQgqyOjoFkdSDM8frthIijeDHhfu54s7SJiM+nXftWMQpYs9gHfW/rZEfQ3tV72ePpDFKQyH4hT
ojddEd5pNfw7USVD7LjmmdA2C8nrrw/Af35NL2krVflw10zlvJCUt09hVblWhMDyJhbxsSjaYATC
WOCydPVSnCqszr45R+YW6hbkjJDYHft5cogSfOEEhM8EPWyOU7g4j9WYwQOc/fzG5a1zlTQYk59i
H96H3SeVevKi5Cl0Wcnl554hMv/bNlrTZIRgsxW0XG/vwOhRWBr+IO/PpYeITWo8DCmsGU4kuR8B
+JIfAvBsKktDt+IhKdfWkxNco7SnR3pgS+X5zfGizU4W9yzLeCSFuC2wARCvtb4nYzKeJ8gxfPoG
WZA3ZAnG42vRaAw8r0B6mElR1DS3y8r5/2nYQOoaAQXJuDFHd3O5E8vYcSGj5y6yMyRhPcO2Lkd8
BVcN6vAbslKov6VdZDG31h3AzDUk8vUiwku/xGXdvOkfRfymRty8+KQLJpLDGODskyy1c/+YX+Ct
hLbem1MPbfkvLyAgrVwsYcrn/Z62Lp6ioU2xkR0pG5oZcw0P/zJiw9HImrWw0lpCuUVvDswi3ME0
ie0NzplZ2etLwIHwwFOhh0/md1sv7OciJ6kLCayMf2SiiXG+6IusESySRn9XRm8CHIMF697eexic
xFZ5IUAXSEJkaUjd+oSmchkyaKNdG9GkfyGgP/EkChgkA1KDGxxuh9+Kt7TVz8irjnE0CT014Bsk
0l6VGFNiZqICyybxx6tLbhxQPeuRKD6VjyyEoYOlYjYYSAwO5zDgMXi24cGPrhDv1b1cN2rxs3yb
4dmaqS20LvPS4rd6IzU3Rnsy8XAXT3ebVNDqByOePy1UL9NZzc/yC4Pf/Sa4BQFE/I+wSd/6wAbv
wCsArmk9O8ulyj4Oxr5a3VjeMB9TLN055GeZCROaP3LDA7C1MNOkZDKgmf1GtBqgbFCd3b79oBCl
jT8GC/Y/IlV1NbW2N/JDenS/Y+Dlq3q2eGdm92RjyJrfVGagStMcyk0Q0nf1IROKJvtkuumgxW5l
tboYlDVa6b0T2+JrYOyJphR1gp6fuxoO2g4TXrf2jVMKNTJZ8Y5cdgMSnXWAQGgCzcbNOcCpoBbd
TX7NO9hmDet1sLWMyhwVsuE3KitN/REXjN/mGPNOwOdv6DghY0bBT7a4qX3NcMUxA4dY+G6T2BY4
pIj7jxvQCZZ8jgX03sBhRAmFVLYZbmcBsaEQslg8wqc7/q3fDvUHut9QDWu9eVNhPlNm1fSL6fUV
JyrZ4KT5GVDFDEGR1NU5KhGz1zQTb3kVzkz7s0rdLe1RJ462pnXTQXKJHHLtzbu9LEYnLfL//Zc5
GygmGGyOnZZhzWuriRoCdEKrnTQj2pv5IMNn5231gOUGf6gmjqV07cYrDok7DD7I8tm8/u/VxGaX
UdXnEB//cC9zsvMYZiAc4m7duMcpR7rzBVBvJZZTFT5hMsg+4/2RBcMcaUuTkyZql51WZHv5nz0X
EjPDirsIKsGPZJJblE+p3tiFo24QPMuQReB5UV8UdOFCe5nUlacBwmSdHYiLWJHEDdOfHWQU8F33
XDwhU2/fn3LR5kbsTkHdqmui7/4r2jSWB3Irdg5K8gO94PgPNwYu6/V/WOOegLAvsJKY6+5mUAwk
HnZh6JppDRj2Gl0Jq2tNw+2WZ950HPPm7ivTiHe2qGBbdxxjCBLOCW/G9wBDyUn+FibX3txQshg4
UomW5cKNikDEhddZ9xAeeB/cVsJOnAlVRn2BpXx5hF2+rqqXFcXMHrIiwBdPy3XXr7TnQc67EYcG
vlvjssC4apv+R4e1vnzLzLLL/IDCndljrHEISWrncbkAcBMIdBwFBw+yx2py9FW5V6HcYwIVOTER
wcPXAseey7RAPZPSjpAYIyZlWbUIJYx5imLQc5UnAekZuPlCAbHH9BfNdNh7NQSfYjQJJrHHuXEr
6Vhct+XXNVgQ3w/SiLhIdLO+cfuH68QI1P92cdwqEwH6CUz95SZXAuykFpCxgzfotSeWDrd54+db
pQgNBQoG8Wuw9SOr9XyPPw5UFYlthBbtEIzUSmSJw6pkt7ZT/3ye8B6tUeGpkeWRLzl0sRsKEt92
FEHvvVLmHnJ3QoikNEfp96u/EEoBphJJv574XheWnW5HQpw9G/eplv/NxIco0MNEGb6dPVzrOMt9
3Snukw5Pa93r6pDGv0hRXRNjF6BWvgqfNB2RoTUxCwm/RjpXDM/MAeEHGKcB1cmY9g9awWs8Qu1u
Fo1fm2P/hPqBZCrkgg/SaUPWyVOp3fo5HMXDZgvi8fAuvI2m87gAgVFan3Oa2d1ka8Qd5Q4iEXA9
X9Q1JFBhBoHBPG7VW6/urmkROoLzzZpj5Jo1rov9ppafoCl/JizR/FPSyqyAfaTW6Qo5HtWdvrGl
THyTdtJ+8uf6xOKTO7gxVOCtUqSidkVFerGEVKWTyD3fi9bzDrSh2VOhFDYGglVM0z9qoCbD6gQ2
rtlyauuetOw/cJdfqSM/nH0ZC2ZzhD/rJtdZ+EEcannwNZznLDEEvGh3iyNHAtrgxDQNYezrlhL+
5swF7WfjrP2sPw1k5rPnR+bwvAszhRMK7RBRMf1rMakLu0PBWEXSCi/8tN9yojWs0Q9OMvPT5ZUD
DQjogtdv4yD9wuj8t47WWaNwoxuF5Y+cmgSiX5PsZdoffddWJUv+0yJTMZXauIvUpLHHK34OBIYd
mpesDGaHMc5F67H3Ddu2nHJvkxsbBKx+cDxZ4v85KWS9jv7L+mGvshI7flWPEnTI6CAWv9vbN9CS
jW6UmfsetOT5kBevYwamggU/qogaXvILKLKHJl5yyzESQrY2+RwSkYbMbr4y8gA5uVanWA+NoisJ
59Lo2xSGKkEPkKXNbBshKkF62GPo5unsnDYZoQOul86QeGGEQbSvnzyGmh338WDZN6jmSDoQB6GK
EpvhuY04iEOGksWKzOk6adu96RkkczzuSHmWNd4eCra3Z+JWV/3cuI7mc+m9nzIAzxaqkqpyWDV0
ZTBIGZIOqpQEk3aWA1zQKR3zDeZQoAPJt2LlvwgMh74tPZj3wh5+a2pGCMR/DxgWVIlvLz0icpWR
hHtIZZ42wcL23iBw87Tu8E+Mpy4v8svpZO5ax1g+qBwfd2eZmNhh4Bf+mK0Ms79WvxjUjP/HsDS/
igK/aMxZEa8cWLmn7rlsjkEKfakXKXOyj/MO3vnKYcdW8oy+sikTtb5tw40BCM4NUKMxGT/MwkHz
VFpO43bmnRRqPs9WuZRnAIItsIzugaOI/W2ECTHnozsk9xmP3kqPZFtefjhTe7+lSrnHQVqaW36R
6H2DcxeJokBcQIjQoZLqasBnxztHbxyaJ6i2nhGIfW+LHSktx8iad/7AGThbkgfeWsKN3DXLaCR7
CaYT1tBpIdXRIXjh6QqgMBtxqpP+NbL0fE+Ppmkbk02adVd2NOolMIbP5A44/PQ/VL5jV0T4cln9
1hapKbfAZ56NdHHB9U4EpmzwnN5zWji1KvSNDXg/YIe1GBhkmKbpH6eJANCnu8IS82j2KVsU+lBm
G9NV/p4Tl4Mdyz2tREaGnPk1/jeUWnQTSi8c6PExQBrB0XuZf2TavbYu1/WZLnoQZzgn+jWzut3x
wm+AH0MzqUFkQ2jNs0jQfGH86qPaZRZtPfTz3kaC6D6sIvb4Xki4hp22oMn+6DvPwWH7nYQ4OZpk
GuonH6pird1ZllxPI/Iw5gXLKLyhGojQ2fS47v8xsCuMJd5JDn4pnV/LjCk+bZoo3f+6gxgWgDBH
rdSOqMs4SP0bdZWPZKzO3ciWMJdKsDlJy/NXgYWIqhwY+mDZW3tdUjAF83br5zSkThbCz2tdC28q
FoQ0IwpRAj1A9aOOmY67h+qn81Rg62stf6zvIJZfgL/jLk1nwA3rWppi2i/8EfTeTb4E12SFOAQ3
CZml+aYSb5Z9CliyMplaLpk+AGV6rPGAqSyj/T2VvZnLLtf5HlCl9WSidbo1Enm3giDoXPrFZxKA
uXm6xWkIR1Gjr9H4EBmUAz82r8R7Cgcx5qFfJkPFqGIBk1VB/jLeAOKcmM8BaY9fHScwMlnuN8L3
qX9tGbR738MhSJiEwPytiywlkPoFNxWPnCRUP0BkeAlm1Mjd2VhIhUC31NTdlUP6kMZMiHfuL8CK
56GngguhHKJgR49D2SOZMbn+1C8B3YkcQI1rHdea1d1JQpbf6pxfWbY1wFwhJg5J9OUedo7x2pUw
9z8qk1bj2vZOxF6eMgvK5tDkSa/ANTwtg6VZ+jEuQO0vseD4IJT4ZXClbXrZdVP7pRevuqPB2XxV
MyeFZhFu4z6J+DhPDN1CUBlUXdbHoI47jYpGieH1xGSbU1zuqYVPU8bM6z+V+oDQpNSQUwwyxEqg
yYuzt/M0m0bEVqB8U0pXwND9bKzenzSjVdUDRbNt4AMfV2J0YsLpkQuIRhQbnG7LCBvlw4MmJahe
+nxzVyLYwXsgbrDKf8tRcNEtZwbKtuQGT9LsQk/urOi36Ct5WrLvOgICyE1NTd2XbZZwixLQYAsa
L95kQhDkeSZTOZ407Z+xd/C35FWniaCysWBs2ss2qf64+QdJn6vEW/BzqQGzPCmwvfwbk6F0zd1z
cZME785Xcdf+JQBlHrfUecq7juiluuMdrSQcXpnghRR5FT5BkbSL9iL4tlnnnTmJB+xJpcc+yZux
F08QwpxcZNSYAqlgSJgpkmMhOOrfqEol4FCvdi05vD4vRmgAJWN2kCW5UMfuU6Wl/VkXLOU9Yr0k
6SqLB7v3BFWFy5wlRjpAQ+o0v8wdvT+U78mn/9GAwdMD3TMR+z0h+ujns1+X16IHgvBcAi24oFra
TzCONgcCQGtLZz6Cb5bak3sx8HStQwdJxVjW1Ly98Vf7jIhkH2ydrhlrw8MyicA6qZ2L5Rf2RCRD
uAul44H+IW/QqB0STr8xMhm1aINJwRgUQ8MWw6lvfW2t8IgcvqRt4LL4gUPu/SIxvQaq1OXoWj9Z
qnenLzY0rZ0k+3OcMpL6FaXuBdfxGkfM7Jb22tO0pgbJn+Xnb+idKXXWXvQmh1a0fhQxUGu+EtRe
Zr+DZ7tA+65BDfgpNWGh+G7p/4VffMgrJ7kPa04DBP9WF2q4c8uJwE4fLRBNChZNtCPKTfQGGZvh
gPltuRF5twvnt16I12M0c3eNZ/TyyyWI5UJyviwrFGDjFv2hQZxXPkgBKwnMU1ysFJxz1Ke341RA
mOQ34RYpxXPlSZTQg7l+qWiFGLB8mJVEYO4D5uOTLuiKd4mHrPt1t8nCTPyX0Pakk3sNJHwDOam+
KFlrK8gxxzmZbs1cu5FRix1tMs1dQBqXGgOMC2Lhbi35IchkYCzdhxlBBxgh3aeqV5df7dOKlP6E
f9UM0RIciax5qtIQ+fMdWIZoiA+iSGbwVPNvxJ6s3I1b1ydoRmRdrTE3Us/baQ6p12KfZK1/Y1JR
WUZoiS6valGo/mIM7G8LhhqtUuWDPX4NBBI2CTsHtWCaXlW3IcYftROLn6pzYjHQIo5S75/DdimN
f24VinTpB1Pj2focisdFk+1+zHwYaAxRzhmSW9UPE7rIizFRx914waeS4x0ue88M//Pfyvk9im3h
74e0qTp8UQnfT9nHbOpK9arh7c4SMLl5ae7e94hK4T5AioWK/JqDv1+AqS8ywz/1JG0XKVvNovCr
w9mdFc78yftIYZ2qWg0uSOY9CQ7J4h+H1oTTeI3u7o4gKQvY4R9r0xjTLGB+bq4TgC9Ewfv6M38L
Ewqc2YONXc9tme2UtRLHIxuR/OgFnFVk/3yGo/K11EpGTNLXo5s6rECFyJ+H33NdfIamoiS96ux9
QVETDD61SRsG+bzkV5/R/gqSfGhpr6BYKYr9qdfO6iEKg9AJYiWX1V5Vqiyz3BG3zVmMCxP8u3lQ
TCAzWe3vKEXaXK2Bu13bifZ/HgwetmxC8u3+ChMAwDnXZp+Go568DlalQwsEjqATFyKtlqzBzxmq
66FDiU0uwbMGf57sbSi/J0zAGKGwF9iCUTbvyLl9VO0bQGR1J1028jtDM+JETu+2OmriXuB20hI1
L3UjK1E1MyHTPHEoz7nzooKbRNWUhOcYRo53+v79ixoFglC8I5LWrK5PWvuHb7S9wsRDXpGUmwD0
RgXMNp4170dJh4E6tP4Pk6dUqz8DwVWIjSUskG+g/ZXU0FyW+yUGx4E6CTf81FfaAC8sxIl1drXa
TIPaPrKDxlMvtjVHdhICRFLSVaTWjxNTJkD+HNmV4Zt4+xD6i8hHjNnZBItdXXOWocGnZIIz7Ng5
17HVU670PZvc+NVp+iXiELvp23Dxb2jp41pxcM6ter6X2PChaG07Zwh1O1oIVKIn2ox/IUXBg3Yv
9M6amg4G8wCRs9/MYtJV3oY3uxYAw+U+74DEhpZVKKssbcYOine6bs7MyCKA6beWLh+t71a5dnYf
j6LT1U5dpD7xp4R42mU58qmSg5IKBHyv9IEEsZcRN9IkF9Z50DF5Q4/wtX/O9g/qEwYJ/jDZgadR
5p3rWdag92yXgkNiHvaXnBmZFS4TEcUIsZ0BGz4HFdfCHqUXXB4YPACS9l/vIsS6rBiJaOLhkIjP
z8hgdfugF+xc2C4wPXFLNazAoZzrdIP9Y7YOuwlBRMkFUb5eEKpEWeUiQ7pKvI8z5E/zW7EzI/4q
ANwBBaH36GZfvGxRQgNC9OhwkzcIPJE5ZityJLjeEQDccvH2zE6zFhWJsTRbPPXURlHvIW66y92c
6dd7hYDjbDoexc5pAl0BAJH2A8k10NNH3Q74SH8Kn9Xojb8EIA1apOVkM8qWCbfbHCeWoN+LVJim
dRSylUVnZ1xw9JccmX2un6HB10mWPf+Ap7x0nMPQK0xvINBZkGFIdy5XRsfzkefJXBHkV192lGQ1
Ayjts3x2P9f62BFsbZOUVCpRDtmqZs8IgRWYUVCiA5Yotgk+yP1WbA8gGlbunvv95g0BT+5/ZWQ1
qP/SLyrll4IBMSLdzQerOdWfInNuABz7mDr7ID0SEJiWyxn0bKwgzaGpCxXw0JGSTHptOnxeS7cT
JlK3Ab5gDuPsJtZCiw6J98gZk10BF5fu/CqhUY809rcMrL6LT0LZYnxRGRIIvhlr8uOijBp69vJW
Zm4F1zY5nvnnR7uuacQEfjnBGHdrvC5vVPVN3oDC04zRO0+LaCRJMi793LxBRf0iLMl5I/RKqAJl
qns6Jw2vEyd58c9h5pufQ99RgzsMrWumk1kBDxIdBtBxtYpNAv87m3+eHM9vlxSKRQYhThNLTPSH
Fk/m+4MurIftWjOZ8Og7QVYM0TeQ/s0p0YJJMGCX2VZMiGGaplXv1ganl31jadG2gndp4UfM5B3h
1dtSVAOEsV3ozKjTx9qZiSQ9R/zc3QXq6PD8U9U8bvl8md1co/ruJaAeE7cdEHrJJwFhQKdViTwK
q3Ox+vFOdzyvjAqaT2TVW7S5iitXWnSAJFWxrc7aQj1ZKCeOiUT6qPGXM1/IyZygnDMRQNJlmkRu
YstwZ8wYxD1DQ2CAa8OIhJjNekbmlmoOQFUuA5y3X/wLAdqTg93FZKUuOJ239i5+aULzUuYtlqts
nOoEehiEeUPsCDLfxrhKA7CxGlVrl6lStzXBo45rePdSeZoBrbbiMGoRMPQ+BRvkyjIVtJZd6Cad
IZYzVMbjWh1ibq5BI+tLVxT4Da3dMaYPzvHiuyNSrbicElH26Gc1F0iE5iadXp8n/9a+ILXsaR5c
ITJoJaMSNCuwtWLLTHULJcuZqUeE6YoLSstcuIxXubVTxFttPHjq9jOO9Hpn9jqgC9xAz6V6WOiW
FggPPUgjLiufPizw4yfPSiziTUOgVG3Tkqb/ueQOLEBEIQihG8eJ0U+egkmo+0FTVZeTkrGKv0Al
uqLjiw+KygFfLH8A+aFrpBDK/PN8f95rc5gM1p7ITfRNYygwbScii0RVpoCgD1dY7rqeCkA0C95l
f8ssUWsj5peWGFoO8uylG7Y0btivGWVOp0szsp05IU35a+bdqpz+ibdSBhKhui+Y9yuep47lPaMW
zbR+3y26sxpUmGQayuEI179HcD6CrMeCNZKQkznGgX7sreBPVTvMTt32h+e+TwcrVKTWfGzQhaC9
3el4K1M+VUcNuq3ZXekKVWxJTVaThxo9HXY6BSogBt3Z0XlRgrUUOB6/IHErW5hG49sqqA/wWCAp
nC16iwmIFcHXDZqksBQRGqce/7Q0O56axuAItx7PJQ89PDOfRbi/yv1Sl4Na/9PRLsWFhqY4qPAn
Z2kX3gFEyykCeNfc+DtWdE9PTJ/3gr7Q+QChSycC84v+WLOllIVION/BkRBYLAoxtBuUJ0GTUcyw
F7W+mt8HikurN4e9ZOSLKCUcT384AL2ofdRj097CBXXVu3Wt6d7jmVA7p2fXQUnLvLaMp4hcTs2l
hI+FKFMQtrJr7+yjq4Mh3/gBRs96Cd2E9quxdOEpG6dwu3RN2MFmLSMk3AfxIcqN4vTNwK8d318k
N9OkBMmzR63YJ761679AmMp0ArsM5WbAjiOIn0Ci1iUPs9JrcUNiDkrvLxjAE6Exe/VrATGHeyky
TXKxyqIQCQIOe7AGx2+iBO5KYq6bc/WUamC7JXP6Gc1OkQgf76gvjar7uDlfzAPEqA8WJOcP+88h
6R+rzpAAc15TSf+ZC9VOfTanpL+u3oQHE4mu40OsMq8RusE4BOXS5AeSrh2kL++GyPIPs+9yNKeT
MbwVohmREEwLomSarl2fRIdjM1vz0DSd97FyZYIeybBITNeq23qQcUHLw/uKwVR34YbT3G+qFdw6
XS3HjJYh/0NKbdA4kxvnEBDqEo4b7dCUTq5aRtM7Hr6YiKTd0WkkDE686ZzWkz7kurzG+ldIUvXr
7t/n5/3cdVGddDD1/j8yznWQlKK/cQSDlKRj32V4ZA4IoJ6Btrb0XB4KBEZMBBYYfsAt4RDCHxRZ
9j0Vh8Jn8xNIEgUF7e+5wAGwmgbtnRNF/ZsgPgbblwu9y/qHy/synPgdJGj0IwomCEFQZyRg85gG
mul4XzdLHWdEWFW/WV9YrUw324KDHxbd2LC5bBOfstpiFJY+EA6wMgGyXrS3bIwxjnzx1q4oVCbJ
Jro/tGz35g2XOhHY+ZMRka71HZErkVntREWXw2xjBhfYitIMnH/M9UKFHIiFjPjhKICiuHdCcVic
ZIGc4S0b++MNzKVrlZGqFms4KG+VwKaEWdXUSmBAi1HQB6ynPgvIZUirAzggQlZozc+9+9tIJKJL
V34waF1bRWbUS7I9Cvkq3gRKQ609fp/GfhauvxtgEmyiJtSX1yA3nRZtf820GuEwVj94SjcoYJJq
ynX+IBLLkJjJewIo9ShNGcrGBOuyrjzuOFyQ+EM2b4UIklyNOQ3hSIUbvA0zntvaf9r24GqHWOKC
7fmevuNgJt07Ls0397MtTZIkoY2wOhjfCOO4xkfGTWidZHS55ZH7f4TlBgABpqlabIvTjRM5gA5Y
vmrRAB82upDfMiGx/2ZFRy0yT/y3AfI8qDSKTlLM1KVhOHlY4UtUV5yPlVbi/eGW3UsHFr7uU9CN
Om03gO5MK9oyFBlXFvYPLWthpaBIOQanhMZAGX6+72Sxhwk8nL7rABTrMvIIrTbyYBy7WVqfAVzA
ZANhEGa+E1piikUzasuzf7GciPjYhGjhBuRdGYal/7PggQgdlN0orgIC3CvI2rFH+DLwhBrBk6RZ
OtGPf8MTrisYDX8eSmAS41bCDPk0NYTdGo2XmcBD5/lmjWo9F7RTrtZP1Z3+rwtRFAueGaBlP5is
47bYFUvxpn+HntqJZUhMc52EEWRjhEoc1caa7E1hiFlPGGMKEsCAqkF4BhmdY/HIjYjww99mb6pF
HCl4zwvvQzSzozc11rFLCWhjR4tXVGe6tSoWyJvjLk/n08BIZuwRd0Mq6nbkG4PqxJRREYVwEz2V
C4v0rhyAL9fFqJf1TRgXSqiFJkGOCrRbjQei3TFmYTSXuTPAsmSBSdgQKfHlyYp/4XqCbiLYNg2s
qDK9DJibrX8i0jBiNABBtrZdDt7ssE2PwSpJgNjCRrW1WIWJy08v+9n1KLk3CbfBmjeC6KLCzA05
kMClm6p07NM8vnxqdFNNvfbXWKbdIwN7TU2isXRb/5K5Gr2Ekj5r2QYCqSzgv3nz3KbptSzhvpCB
hZf3GwNNU/Pxsex8i2VqORsVMUQVxV8ZYuqGGucfDjH++Yk1X9U9l3HWst7VM6TS91RlE+ALXYjl
ruA7r99SYDwmYkYn0MxVQ0Ak7jt8twti8hfcO+5ixXWN7yXp2yUBY9JOIlpK6/q9u5itqdHuOSqn
qyfSgnA3jTSCJGvS1CDKQw2vwA/4MoSicN60GVV8FLX4N5jrj8lOqBCU0BH2fKgP1ex9ELWl55w/
xN0MZOhhYmUrsnOSdHYFl/qUFaHDO3B+YXAWR6np3Vzl5MDTo/4GXTroVl9kbK9dwB8WtpytEhHv
4aLdUdtFYIdcujkui9DdxZTn/wrPFKyLR3JGO7ZY+a1n0vp2PSgyIB+8vsxZyX8GXAwxYGQDf10M
fwV/tbi7N+XVrPEZokvYT+/S2wiebqpj8CVvfdseDit0VawQwLo6eTYKIReAnOUjoX6+OSIKZsb7
tVEYT5H3QBhLGGGWw0CQIcvAMW3C+k9L/w1xx3L5HnNGny6IZMFDqY1jTk28obU5X5/S760TyA4o
U8SVmMvVGnasOa8UpHO0gfJON1C3rHa1asD8OB8CQkqGrrm7HGiosNEACkZ5p0WEZHn7g9PaS8/K
mcty1viSsAeUnqzGkc51LNnPFFfEXquzf6koODQ9DI+l2IFVmIpApBLRIkrrnx92g/d4AfExolsP
UO0fwSpa4KoRBRqEHRpDIx2E95mp5OXw9HDahbufemHZ+4ZlECL9buZqUZc/KLQjJICybbYq7HZ9
B21vL71WVZe6y3N3krubtC3IaKF0pyLyfy4a318XUP5Fe+iHLgCXFhLb3iW4/6yuwsE2nXW1fLP6
f3bS/3gdpM1dkW2PdwugsOm3hh26IuM/P3ui4YZm77xPWk1ot78JztqduLjxSHMlrN3NJOihuNsn
9W4qx58MPRuWmscX10VJwssPbvFAw51CciG3oThIV8grSnwCRJfn7rG9iIRg/h6NQDQdEdyvsdW/
uKokCqCiQMRpa0eLYEsYDInuNVs6OEmaXPZC2lF9g9xzwyo63CLz5BKwkJm1/3Tb0QxyztYMA6sU
PyH7G43FCOa1Z8Rs94qSPXwQzqwXS7VID7pF2w3AM7Rz1JhAyJ0q+WYM+V6sUpUKZziST/rFkpsi
Hr8AQb7NKkq2Cr8cNFj8aM1QY9X5hp9Vv+khPfNxukYezeQD8oXYK/kdK6/rJSt0n5+02XEoVsFV
UpCE9wR6pV79pHvPjnLIViZo0i6M8l/FcJR+n7UTjmR5fGjEL37hqNxrpueo2RX9CdHnWba2Pgto
8NnXKAwB6cqjbMoWWU8PyXS9xv8TLAVTBBWCZXRd2zQMerlzCvgL6oYCLPGtHSPXeKRxqs8OA7I4
Ts5heRkFBf4nxHDiyoCkLogccLvJXANMVahsLajM+Vgv6MeswBhsCKWHKOiVrY9lQrj9hPoNb68A
GjEdB4mI+hFgg8ZvWG43fjERCjytz29bu2nZigGHJFGHULHShAaLb6lEQSJoWBfIIffeRmMCk2h8
U+gNL6EkWlieR29iA+J21GOojeP0mmzZy6IHaN9Lu6PooC2rpzexmSWC4fAp0+y9+WfR7zu9e3KX
FOAdYqcIC+PN7Iu0mC6dm9twLr0c9PG9HT8QhI/9u8FB79Omy9Zhb+m/R5YKaQQvw3OxRls0tOcP
AWwk66eTGeWiffWj20BAcu56MbftrwlZyeXbcFN8jDmRnTEjceK7VXUD1QpgLKrhe1TBUvo7Sx1i
zuv0FZlPDAX9lr0SY7ZpAR1bgsVfjhX9ldglc8dmKKACgnI334nl9ICmUTHBEFG6bFmWqDiemTSB
kv/Gwy+EZXUNBumqrDCC7pgJ9u0Xbiz8C9615o8Rhy+us+2vTqaxho7DgHA6ukxRgkMq8oz+dPYu
oVDkVpn3WSmTC4mrLKqi/DDvDGDBnimIFEu4D/SellsKJ//qwdqa3QvZvnxG1o5l0EADR2Lt8FV0
cDOqZVyY48TQ/aoIzLK/oFwczvURXooZW6TJnZb2WxtzmBqW3M2T5DJfCisY0zTcUcKeTvYP6Wyt
urf32nAXvrOpZ5QMcR3wdVxinOt1aUUZg/5+D3slQDPELI6kcgjEygcLQsW+7eRfk6n4+Dsjqhiq
MYpy/vQ9E2Mu0Tdg7jQWnPa+U6gbKpUvBjpT8mHFNxgbldqN7KqyU+tSLdndbsO8vRLn6cIQ+SQ+
oBPpGr4ubyHHOart2zZo1h3C7+hAro3aY2PzO8Bz2C7hEuAcAiTjmVS/tbgD7eNILPNM/AXAa1qB
52XHMz71u+wz23v/qdFybxzxHtpXj0vtAhfTPnagP7icIQZPjZMZwj+hyZO5CPo5TFSOT1LPzeai
LkHhpK42wWCDoyCBpkKHgEVvcZ614cAumWSk3B3WEzn1oVUvnHLaiTKrO41cfUuqla8YAuxGTUU+
BCZhagjnTKYNYeD8ekgwt28IP7XKz8aJB6IVyWDqc105t+hb+bzHAEMmevHhQfwwskQLlAX7M1vR
WrtegA9dx14PaqFIppeZuX49xzu0Syr4fnUwQAeoKxBGUAUfLzqyERiDxzC6EygSMLFAkZHIW72p
u8G3oezRgfz56qdaw2UgH5liz1bArSPzOVdIFnABCI5B+vpirVCOesdJMggfmPyYTmpUxKZLBC2x
Dpfu4fDhq4opMmEWFZ08UW9HXNYCNvShin231uQQ3ESYvtsWRORrIwcIOF/6zvhmjV4oaLW6Lf7g
SlOhX23a4BA4a6coeEczTWRZ7lj/GRVIeX+oHbNbZN2mYodlDvPKSZBUOy49w8PaiqLfJgEdC9hA
Bb5Vyzal9lT1aEL75jscSUSN+G0p77A5vFyBSFIjL5KMm4cvpeLiG8Vg+lp0QtfFnCN3/XIKzhfV
oTqmihTN/zb8gqBj9dId+ICkOTORv4k8ha/mwQ733fhx5JkR2oo4OzNQSho+saS4O8l22E9QjFVL
RbR5zMXrQP1BrQNurpEEdQu2/gTH+st05JA+YcFSeaqZ2yKqb33+PjhepaMrLX1WsCBEDn/SXUKk
Brckt6b/N7FGDEC4aUZfb9UPCHaYoSRokTsudtJ2Bg357bdBDYwAiqnSTIqPTAhZfVQUb3YWeOEc
2B0PSJpFKZjcKN2O0bXNa+sT+FgZFKRZRL1v9p1z2dniNPGFGvAsA/Slh1hxmlLbkakG+xzQFy7I
gjyd1yNJZSNNTQh6XFaDHq75nBzVwodod7xpEnpKsH9Rjv4nO07/fz9jcI2YqF/sxUkaQrZJO9iS
HRrKt5VoHyiHGAW1XtDrgFR5dSKwMiWpwSo3ClEZF5DGmhBwB5Tw/uqQRrgsUPJSwBK1qvQOzRuY
yUb7Lcr6dOH+jAmudnn9P65HSdNnXel+/tQh4tQJZ2U3V7Bl7wOC/jcbANz9DioRvPkRTWWDvoCL
rF/6Y7FNoDMP7w84DTHIfoNhwvL3p2sb+BLLS4y1OJd/i19YKZuw/diN3WcHCeBC/aqwXUTDsn/j
M+5Dc4EJOqNC4VuvMX2c6EKWNwCOx5yQoGFLk+lFk3bgQIlaR9K+Pp1XxPnFJ7HI9zTMnehrg0Qq
/kFm6dhROU6beNEdYIF7KpeYyMXeYWrXT7U+aveKBTPa3BiO2ee7Ne8gz2KasvHC5Cee6KEFkohg
WX8eTOkqkKkI8INOlDypa8OdVhYKqC9E45qjIuh5s+TeMmTRNjQXL8Xkpg0jDUjYvJmaZxZ1cxyh
AxE1+rQfxX/GmmmxXOvwegXJaVRTtVg18Lx8hrQJz1IUxBur4nfRsdf3ErtjqyT/vJVGwqi17GbI
A26+SujtZPG1vb8e7pmt0xE+QajMrcqWsPh9zkDztMyORedkBB6t5Pk/16I66SNV/2CoSJ2DRp+V
ljaWeOTyr77QL642RBDjOIsIswhUaUBqWEDw06IO44rysWKAvdFBiE15p1XoEwLTHcQ2mpm+QDus
+/Jf4dMUCi4RTM/JbdUbDJsy5PwwlC3FPXJK0CJAhATFBHIO+mQ+W6/Hxoa9gxUi9DQSZQRzSIhn
j5l2Lr57ZSRzij4RRugXy2Uo4aCNwHTFGHX32qtbPy44akAbONDAsCm9erSHh0WLxP3NqN233rZ0
K9BKm+65cd+7NQj3jooLp/CINEbADXW0Vg61wtrC4kfWduacoKqS2AqOcpglCFkwMITbdZXsqHDh
VvMxpcq1UpWLSjt4g6nX8xV0ak0xuJZaW8yEv0DDBKtslqsc+cFYD/MuqlqlwkkRCk9JhupZtoF3
CC2VFrFt1UjoJSAGIAYFNyIcrPJTa0jQRY66N6sODVvEbJXAxoung0CSkYvFajHX6dyNF+5Bonvf
JtzEVHhZ1ZWk+epXFQe5T29Zp5cTrpRH3Cd3AvdSisOhIjP+8ASeDr4bD+mEHP46tk54xFiU2ZvM
4FS6r44mZL/EMOOFQOlTLrZhyeepYGkJ/yyQkjBcOYXPtDUAT1FPz7+D3Rb0SH1FNo0+iPVST0UH
gPSzzg95WKucbXeANQJ1UeouG4HWjQZNXaNwAMHyIs1osOYMkq8HuYWwJZhl5Sex478JzVHIpk+V
USPh36w8z5wlL9XdYaCU99RlAZuY3g4bm0vnf404cC9KCvDKHWDTXICByeOE/iE0SSCmowvTly45
JFPwbuQyEDUT/AqmGc/frAMyNYC4VZVDLJ2eXxpZJTF51ostC47j1a1tzTID0xctyRky/pDj6Nfs
Z03hYBZQ9ABGFXqUOLSqpYA7tppmPxNcDJc3CUOTUCvr7PNnNd5S2FmL81hZ+CQKBbrgQptWmkcl
Fh4m7PGVtYEfUMUyZelONFKNxnjGoWvXxQ6lgL77/0X2H+4aFWs1orV1lGz9gcC5pZYJ5tkj7M0w
+EK3ujGkk35djs775RDakcQR3jgzAlC2MCpD1avRxGoBwC5vKlEJgGdCffK3ydvls+jOTVQJX35s
j/DNDm6Q0kGTQB81HTfe6pqFsG3fXzF/VqGs4rpQ6KDI16pkf/Xj3/39s5C54elytbB3bj3a6+F2
MYHY0TfHZGncoW+RRk0O0pHcQ2cIgUOhnJJUooyuewiJ4wvf/uD4d0wANRLUAMqsToY070b+xx59
87UPYecawIqK9XW8Du1I62qWeH+x09UWEJ1RCrv34R40ViGzYn82N+NJdxqYM+0CLiqnnyNW/NVd
kTg4PJIf4XvVKUDrsCqyo6LJKKurMYvCDZtp/ynAjLT5AyrGnzoS4vrBrNXRilOQSPhFkUj7aqrV
LpnlEAjI56LA7AOBYoC3IeO4TAOTjkGKrOdW949uAYewj5nG71s8m4O/v9sNy5NjaJtsTeQLd2Lg
1ubTvwiN/eAU0SfBOdCzwGuujMZqEdVJqXeSNCHsTebY91fObQ1Emfiv4xIUdFlWhFsViOjrquAT
hD8J8DCpu79SQY4PLXfz5enAM7VRvrkQjAJVJrEnnT2mkA7vKXipGFrXNyxNG7ecBzqrn3akwNNl
t3jjXXbaMiYt9ItrzJJH6pPP7obxxmNy0Mr8mqISq/lDvfZXILQb4K24vpXs64PgXzqI2+gZWK0Q
pnCdfZYiP2S7hICvfGtPq01tKN58TW3HYq8hks0GvBRbY0pBixQiF9o1wsZJdc0+iTDfRlQxcsXn
AxmOTKR2NJl/2X8+jkyVrk7JtiO9ogKt4O2FEYAbPwkqKN162ThfHxWOHwPG0rPlZfiJTlgxYbvy
+5kEm4hzxZh7otyZIwFJxAd+u4WmdlJpTkVSZQDQp+K1/iZzNpDuIM5JndAdmuVbKBnzBxPHRzO3
PJO0dO2f+DZuulF1nDYX1Q3F/bl2pxaYFWdVCekdAMrE9RagADn8Cguu/m6p80cjn8rsZEx/4H6H
bEUytGD4VU/IiwuxpgPORplC7ztKLODWxaFZeriNVchelOs9HCCRDx6E4O3YtoiUXZpr7LDktbTh
ZwKWQLk0tUoMNEiZDz2UtlhCC/NQKc+4EDEzA56hGSNPYK6tVYuSczNnW7VOALQRKEr0vy4XA4vW
XWbTYCNrTRJd7qI270Bd5LH1IhfS7LMfg9Bp1fpusWucmMyiBPNQ2J6lY7EOp7RJp3z8GDygOkiO
ce4q/gyfoRc3piibLLjoXjv9tzi/yidqwn0FuVL8G6WiQgeHvLLK2WwEgulybJyxtKNQpRlpSneh
hxZxFjYF5sQNktTKJPzaqqAFAWYEr33eiUOAfCeLoqg8T/XEVWfQlhJF9FDoQApMF/5Nk6rFfCC+
o0YGRdL90UVlfID8dFRJEaw4hivX3ssRc8Tx90iBsf2NHduo1qL4RSq7bhvWzhpqjz8wFoPaMCCl
j+pJfqceBZPwEduA/NhtVi7XNptaxbvg82gsQYOnSgpawGBEA3xprmU9cSijugS9zwyvGHOSdYek
9BIPDZFt4Q+p8SSxfipWtmKTumZyI5KbR7e0l+EbaiWuE+MTEnTz5sfeDxQYkldnrVUX6qOIqkwG
Gja0kfJZy7j2ia7PQqD1w4f+4jSZBKSjW6Dw3aHWtP8fDL6gT93bSFkHm6LTJT0adiyRIvuQb9p0
MbfraiI4DLiDN91geuKxy6lhUimLiuRPC0O+MlqAESS7TxH75KiPXA810evmVk5b8wVt0airenw7
aJkxCaZtG2zIwJo0Wr+jkklK/T0PHAUXD4VGL868fLB8BBoVeHI7JsaXkgM20ZitigypogsG+Uv2
FyxDUk+nFBMYXEX42WyfNvf2dw+uCwVPvTBzOT3+amY+LgKbesykQUXkn96nv5oYNcWmbt4Ztw28
GJYi1izcRgYnHROnOJSN8CdInvEWnrkkci6cBRxJwNOTJ4Q2ZybNRhtF8EXXytmzT7woQ2Jm4Nj9
Ni1NB4kZ3xf9c3SsnLtV4GK1B013jEr6F1FkWZ9UK0txox++P7prUU4N6WGrSYiCw4Ld/wosf3R7
M8IzxkeEgPIHiI5hq07cd6AtFOWB9IbojYHpM+IZ2Ub5ZwcbO5X2XQV61uaw2hFNt1uX6Ss6OIPF
zDGCkkGAtwpnOnE4CI8o6XipnFyG9kY7FRVhN8K0WefKMdWgoWI8PtYZhq/TuT0cK55Gv9xsiwqs
89Wg0hBg/P4YlQOSz2YFz7295WVj9MGB3yRrPWMBWROQjFtpPkSL7WDhiXNAgfSWYRiZCgrU6EwJ
HxTw0LaWA5aazY79w5GR03bGENbqfozejMxJqdnDxutxi0d0nfA9zXbxnMQxq89wOeQzpIChXxxV
fmfEMur9DQ++bbQndT1+BH659iH+hbCljMjKLwqGPpPdpv5O8A4iUha78tS985xE2PhWoufaitMw
e2hUBjUstsO2/NyJc2glp1ix/2YXwVI6bB7q4jnwxgmR1Ap3tN2nKjgM6upLq1Ddc5bgmt4hhQ5C
QIB7W7Aoi1W6z/U9MDIb/qKtDP8jglgtnjnaETzCvmp6btZCVcPft4CpPyRQuej6dZNZddimPNG1
v0E2LV8nxPQAuu5+RmnlacMokZNV8pZYMNYr6eudMBytJn8Itfw6REYdGorGSKu7tOfdNVkuiXyF
jj3+7JSL3QQm4AIPEAISVArBAOqUH/N06SLxUtMa92QQ59iZQscJ1T47L1q56Vn0yklJjMVVFueO
juOl5yMfbQRIiLsyiJYP+b2Y40uGIpFAFI5Ti8Yauz/bR32PlpSNKBd7ELEtqgVSeUMv7w+yVQAM
0+795nyPqrIQpis4llgJkgUt4w0xL8VLE0tF9K75+4EkvkyR9fXghNMQzDmqiQ0c94DN5ZNCMvZF
2dxL7WVjJvMtkMOa4e5jHi2PwNudKklpkIFhhtb3T34HXyEDLNBL5UiaXKspYu5F5wgWqt0grkmi
hanjGqTnz5KH1ZzWyETB+2rH18nhdJI23L7tXp10S3h16ejqbErDDp5dkIP0K+j8V2NDETkELXax
cqjdLx77PSfeba9sxZtfcZ2+ULwrlNd0dXaOzsHglOW3vhDghoGso4PQOqfPgFYanLVyQU7BvAkp
tLpXVtFuw6qijH8eU85gwgn18oyU4BVY8DeF2VNtD2Qr3CuyX238oLrDMaaEorJILN3oVJ1rvcF/
3n3yDYQiQuudRI8AAq9VMiYH6uDbeh/21YtK05Xffi7Ro6abSzKwXnX89JqjNwWkbkdX3w24rSmH
G3B/+PC8HqQug/hv6jgaFN/ZEXQJoYntQSpKrcWqunetd9Xeo5sOIYgC2ImbCsNMOZy4YThGKpPV
SNDwLx9yFqf6kdgtbLyo7VrlFr355jRqakyDQnWqw8CIkZPBzDM6GjtXU57My8fIubOd3Vt2N5us
mkyLqCuGC5KSKvgg9fcAvKX12l3CWU5KhCSuU6qDTHT+Q4+o3XMiRKRsw/ZVpQe+hEqR1v28Gb+B
NBlpHWkBV5rImoOU0LO3FgjzXBuFl4H8KYHlpGaXs70agTaWyu4jmWb6dQpABnheDs098lu4KmHu
tbgc6B/41ZfSXEOfYKjI52qRMD/E3uNsSKj8NhBM8Zx7UJ1upifjfoOQISFKG92NPvC9pFqbD9wY
zf197Hc59L6lzYoYHyQw6kff0EGtc89LYTwP293HTnSTowYoQJZrMrWMtSA4xZUREBbMHy4naDwT
iHMIHUbTFPnobdGfGr0nUX4myBVhc4BoGT4LGSwV0wQXjEx2DHXXsxLFl3PTQeCniPeXOIL8hI7i
0W0yGlMRJRXgPAOvby9rrOrNk5kypj5uD+gk6JzKl62SjK0STGeTPWirl7vMCIo25/NiBVe2jx1Y
yYz6P6Hqqwa6SSppsTwiQiA8e8OAVeTyhrem2kPJ/lcrmUtyWryfopyZcV6RUpJawLWBd0xjxbM9
42yJCNcBPkIFRt1VWPmJr4/n5gdEocHtNNzlwYROfegqfRCmoxYm2BVv6WMpPrD7I/gJe3tzPies
/U7ahQ0vZ+4GQFV+e5FqvpbwU88al1EP7bSLT7E8KcIabKY2jU759CcQVvOQxFAV8zIImMISXkND
LdK+vMpMTaA5EBYphRL5O1YUrO7/g3doLB03nR7n1tq+r6yV+yAIT7chtWrSZd7SUPOC6qNBRyGg
vOAaijLJmUQCb0LSgcN4ySAigShOu7oyQtnonJFxSNL6aCdzFsvvUMlN3bUC759QOlBMzfUFIaWs
UMC6cVB6njqUXUzsndlcVo89IKuSnkcjoInSfhGrQnlQ5nPICfmjk2u+oysPDdhCBHQxTvZyWmJS
IHfR0djNU8wQektbE8E0Ol2od4KdXBdhVQtAEx/5EQaohKnLbHZE1Et0opfZR/r2jJIBpXyKWlOA
u4tRO+eK+OTPTerTmR/5j7V067Pzr0WM9vDEO1RqZkaczxeSB3/FCDGesYxJ5D1QWFjdH0/TUu76
DKjItoJSGxG5sY28NeI0HEP+8NypNoL91LfxjfDqllnoPtbqS5RZ3LOZbgF4a3kCtpFAzDTWdMlV
15lrAuetVRA3Q3IpMpAI6Vetj4WmfAZw5C8u2B97VxKHDj3yZTc1B8Tl/tqqRubNzm7XigIZ+4tA
cnfYsT5BuAZLrHg1tx3M2RKVI1lflhNGUfASa8uKLpWM2N+Jtra9IEpEVmy/YeUgZ3/0fIY+KHI4
mYvz88IbslGZPJ6jebgYeApTZKVh5kb5T0C2jsO45qp2Iy/9Z2V/iI9cOgICC+eLKPHo2AGjUb38
7iXmcTM9Ich8KnPnzj4KI9bsM1TdFxaSODnkhoMaVniwB4ATbUlyCwBPAhJSdOb5HdFIB3K/6dDM
mF7fh9pCOZ1Bj+72dFUO8BQAJ28toCNknPOLYk34zM+6IUtgmgdDnhIHEe1KUOoaNhrjf/WFduaD
a2mHDR/p8j1SZYH1PbUfDwqZ3NegAyQn5ArCxzeyEBYq70KQX9TyJLObiadkKKsYX0ExSjXc7zMf
9wSnTGZKg2lHhfXgcOm80EP8A0EStwlUfsaXHNdpauRhmi/ZHAuKS2YuyEJkdxBxOPr/DSimQegF
dMwouOpFsFBuPCr5h0Uj4kSpj05aDnwyPIpX6hbbN0udF1My8BRZxuAC5Qr4NfJUnsl//E2cTBjy
kcNP3wlXuFEwMV02l+x+xy4I8diSoA5BDNjaQU1fzFUe796H4WRb9IFpR/19Web3vT2ft0f7TWOD
yKsmwitbULS+/dUwuL/IEHzJu6JL0N8Nu/GG8MrRIGAmXYVSBcwd/tE1V/54X5D/jZVnpsW2T7nG
vrDFYB1qnfLVhDAyVKqau1o5K/1fjAdiOqUnhPQhhNVYUUOkZ/pEEwk5opRrYmoaXEOUnPB6Bzfb
3il94Eo+lFiO8uvgZT+Ia8wp4trRvIXIEJgwRfV+9uYgoM2cP3KHBxFyQ0IhOxrGnBj5A/qGnJx+
62A8DOyN/dOmnYxqrK8qpdV5thNjNGgVJBp3+xJjEARaK3l6Ee7o7iGcrRoZ6oXlv21FSvwsT2O/
MZVKeaRorNLS9oYJ2aXoU19l95BBhNkCDTgY7JI3AQHDFkmmH3KheEh9TdokYESub4u9yzC3ui1S
D08wDEmKTL4hEPehrf6nJGEJ4sgAOmzs3dn+yV60LKpx2fzbPT7vc4RbNs8zGGlT47Ih6b91xrRh
uL4uezHoZhGsXNvGOe3YnD24aMgROXTqK8hgEwEsKR2HaAIE81vSIH6ufYjDOKrkDCD6Fch11zZV
UUTbciQX1ady2Hgrl/ii+Fs1m26URbbNq6et+QoP8fAloraRabNfLofqdJKBvKj9qAebhnmRsKl0
DkC3Vfir/Tgf36JAa7ejIwAAgtUCNfb544MSP5S39ogqY1SDWkwuzaMwdTcGFx2ocYVkAOCXSgbR
Mns7UbLQA2/Pu1CBLpxBnvjIuRnvOeK9cY9NV8N0prYth8EGABPKYf3lIJeOoFbQOwK+i6xk9D9l
YtovlRv1xvTI/4wtr7oE/mJ38OWBdX2wnVBBuq3gdmip0MhlWaLjauRWKtRLjSgxEz0qUyH70PQu
dcn7QCU5wl6tfjtN2V1yYSTKWUX6HdY+C8X2KObUmrDVwJVVlmmP2/ddDC2em48uJSRRdghcuCdj
arJUf4rLKlgAvP3cbG9/5QZ5TkIMs2mTdIvuKc3/QjJeJgOc/w75J4qHRaITNnITL/Kc2DPaZhga
q738KvQz4FU6pjMjiPUmu6q33Ryo2QC0sYzN4lA0GPeYcQhr18QaAOsE8f3xyVvGt+H+SlPOFUsm
LgAEo9iXckMbuFkB5mQ5f7cjCxFtOsiAiUAMuuj02phoc3AuPJ7BHcQyUiU9dxj1UtQqZkM8HaeN
6G3zecReenRVORhPXXxQhUCK4qzWHD84/8BU2YWnkbiNprx5u9Ef1FotREodWz2nQFbUwiI/Uhgs
wBO8VOyY8/f1IKxZZMASo8WPK3rH/2AhSlBvbWW+oHiFwv4mEfanlIgaO1Igx2t9gULZ95BDY8TM
NNFuAjkv8Ee4fDKPHfQLvhWk2fngIw9L4QcXPLuOSmRJrwkqBV+s6L8cPwhO7BfhtK0vwoa0+ikh
X233iFSiEGBfkWzVmuvmRh+Su/SpF0XL+QJRBarNsU3hl8ugxt3LL8OLvxqdpgUIeUqInbbdIVCN
L89i4FZBRa99fm4/QLTRnbtCUNqfG+IIzyIkvm65cc7CUTLhNnRdIFsXQFGB3bUQbboWFI2Tt/7k
9K2+svV16UBASfo0+X+hdG9SqWaO++zoZNYbjBgB+zgjGPw/vAIr/OvO59z6jNNusungMLOhhYqa
oY+cF0k0/1BVg/VOyTJl5nomZbru17SWCeUCvnKvIbDiwFyK/KM3pcfarpSmwqEOsI67xF9GTRJx
7F5Zfn1Bew4yIl7HViugXyI61OYb7sTv0X9mZ9rBH3sF2KZNJySZFeFosOnYkZ7JRkTyKL6z6UPO
2fMOWDKLyA8DsuWSvYza6DLtCJw4L0EDYcTqKCQKypZOMEEop2TzU0TCS54RgbMzloaliRSE604A
924wYgw6zgdTtTEkMkk81tnugnZrBBihPBNHHQHSI1gla2LO0d6f7+U/xUubHXbjkPfXuLkzxbHA
WOxwOHSKS5yMVHz2XE3V6XCw73gxsAhYzQEdh0akje4L33X3hnum9B+S0YS1TfkX8ca1okKSZ6xb
HaZ6mauqOm8FSdJlIWisPdtXQOnJbyjfY69r3RnIWv6SBr/t0FIVuZ/2QYny6/6h4iEjFfdmfH45
EO5n8v3WgmIrzpbMKE7C8+uvuc52uDUjOA5nH3DcyK92fwSQMJ0INkMjay+RyLyErEnQJCi8T/H0
HZWdEo6Ml6rWVNrG+RKZ9bAAW0idhPOu7f6hKt2ixZ0dv1lOOytPgWqSlD+YFdOulO5nBl79EfL6
WP9vFd4smPoRzUzJSesZLd/95ko6IIgMj4OZEJzvvJYUCcpx87NEGLK6PVnGRqqG8Gt/X9NWwY24
66WaS2ZGqkpmZK0se8ooSHqfk+iJwFRmS6rCjVrbE5ONLF6KeyNzF7+GE02AL8AaMA4AdFQCfQzO
jU4FGbj2l1u8XBr+5l1YUIzggovy0tvdGRHqnQfVG28yozfWsWKrhaoUCrRcP17PGwOwRdLF4jX8
OAeKuqz3KnlXnqAr1DYuFT0G9iPJ8k0JpW6KJdxstfsSXqyFWWMWP5+qfbtnM37ZCEE3ZS53uuAl
/SYPGMrpsCFjmZMAORFp4H6ZC0TvXmT4AzHKsCtBeRlOI8wEpZkXsPAsGsytn0F9HWlGVQ5rTNs1
oLrutDGHfLBBioqRHBs19dDEObDyuyzMUe6iwEn1t6Cd+L685p1QYyrHF5NI2SLFIdqhBcq09UKz
/hpnHa88MxZdeBBOMZxxaZ2qnNSNtj7iuUva5wFHKPwrm5xDEB0RCpF7V6iT9c9Cj71tddnkhlUY
Xng5mwqZ7ABQlAkwQlxEsuYkSbcW61bfJp+3wFonwxwzVUtkFlqcsXIJ+jkxPoEicqDlzH5nUiep
IsNPJZQ0aHF3dJbZ78rZFeqBWkeeAOO3yqAzO6q8K6taBrD4x6Itpg/63E5DgNRWvGCs2k25qavn
+zepzv9wBNdxyM6Fn8kb/bPj5BaJvBl+69PijgCEIWQYMLPnh8/WISQeoCzSP5IutosU4IFGnvER
Tmyxs+KhSd+Nm4DQukrYmlzfUxS5SdNMSbbPnE7f2n4wDrH9bK7PC297+mT5MdOQHd+YIqlrvDtt
nJoSyu5ldOZe4CjWBUF6EZbEbB5nu0HqixGCqY/oZJi+MujeUq3YPIMF29U3nwWyMGPT2BcwCkdT
9sIQsKGp88YnVdMkRBi+2dvACysYfos/pp18NoU7fJT5JQJXsraICTk6jiYToSrGQks32vKE7VOB
3Jnwhi5cLcsfRwyCGZ7J+ku3FZZWDVL+56C6hn3nUGWdIbKdbvJWjG3LeQGEUu8260XSuO6soQQv
lnzvWDu8nkCZQpk5/Mp3lgxDANolShEDNS8vIn/09psOYbGFsrEmQIj8kGJIEPaKdVjI+NiNI7TH
RtjcmHbE6zD3QDkjatj8F1CTWw+HJW35sVEwzIb3MJbk6Cz78ib8z14mWewFEVx9+mw3PXZ3iCbc
YYcnpgNzZemm93afL28i0R5q/0BdwlaxwHS0LMK1ut/cyqDmuspZu9LzZk0UG2oABk9u4Cs0OIzd
M6fJca614uecIzwNjKR7VBWS1Zpl6Ak/qg3ou22j3BrJx16Dg97YxJtyLeis/SqTRTqa3ujdunq5
nF5XMYQkWV4+kQu8hn1kb4MQaQilC7U4T6n2IQQcSw7lKotwHd+sPvk6wYFR5bJEq/QsNPL3h6ip
Jvph8Qr8Gf+yJ67NLE50qgVOIwmfGFE018zhux5UwL9jbMvbSgVg/cePgqtkC3MJK0hqY6P8xftN
y2itv2RDsQ7n//1qN+86R1GQ2olftV4qLUlE9MBhW+ZofT8An2ECHEWZPkNXBpPwWVhT4GOc9qHd
dIeqAy1v8mpYBKMGsUGqZErrA7mEI2FW6y5/pf9hY+EjMMdYaWb+lnRR+VTGTIAeosi2Wkva/JiA
rXf4wkKwlFJHT+IjsftJqs9/DzUjgpvF3Jti7Ad9hHw7euyDg4r+9P/t7Owwh/k19B/NxnM2vLQQ
6nwhtrQmiF/6ofvmpjPWb9luwuZi3sf3M7IorvC8owS7FOOiyQxs2gDsWkVXbi8ZqIUU/5/0+tkB
czFRoVKbLG2i2aHzQ/ITm+dUXZBZXcBsJgHVGBE1ijuEZOQ+Xf/gyIyv0qI47wP5zLGJekh81g7n
RDopxBnF8Bz4kWeRkJkNDK4UrRG1w6fe5UZGMMpIpEyX0sLYqbL664BXCDwk+XjQGqa7u5O1yoiq
GJklQUm01Pn0kPdgvhrHK4SnMgzwH8d3mHO0QQarPPzP7MsTiRFeHWSSFlye/NhgDXubqqo2+hzy
tgx1nPMdkIbfcH8o8p+w98JmsWTleOcGGhO61l8pG/wH/cE2YUZC5JmhIdyvaBdBqSZliPrJYOgB
IFarOM2rY6vjfJASJw1L+pojohCvkEGZp5aKe1RW6epKCpAMSR3cfyB7gR2OpXAoy8B1YafntmhA
eBrdBibopgvKFEKYN2eQgQLH9AcSup+tvJqat9+KUSeZm4HNqvP8UDro+HUzctkODrv3uCCGYQDt
JHNkwA2dXxPwN/W8x1Fu+WxxUmwlqnmePJPkOft/T+j3yQbZzQFr0FtsnXbvL29MfFVE03ZKsG/c
AWuncbi4hufiq68zRfZcHdjK/rFO2HkoI4nzv4aaM1rTxiFbi5dhAYyYwEwgtbP+3P0leKdKKELh
+UH1CHltdPRktwiWUCQSBZ/2/m9PAoQlL+qzqHChS5/SNJ8InhqpNkvcpwYlcaK4A4DWWpdT1/ha
yHhBBzA62vDme3VvTFrsUBOxdiwJUflL/OUW0jLrPDhn/Gs6x4DHHLSiBP4VSrVPmXYg/wHu8H5K
+FpsZruoKtS4v5xWP1KCnftJnWoO2LXtVJ1DoovOnzRVSRZkP8nrvOM61PrG4ZvApWb1QndZ6Tgq
UdqAWl4aVgbtlExfzEI9fQ+ZgDtkF27fBFnJSPhqxIHpF9GIYRq/AijNSOscBF7uAiTN+M0qJqn3
kAhzYysLuqoIvM21XB/ihordcwK6dF8mqUtLUAs7B5RPv7MxNo3AeOpgnjfVusKIogUDehiCQCRW
sQG8YRLJQibGWjzuQga2Gl0Q+EL8+bdo9IRffh6JrRIxvW+3cacLayB4J5IZ7SQN0oX6Xb8mOtbM
92NumrNneomBk15IoRIhtMiYoZOJo5iUzkzH0N04C1FnPwJ5aSXXGP4MoFd1/PT4Ork8ixRAqfBB
gVTX8/SGmKwSdsHloyAqzwLu2hLF6vSn1IBOw3ezobsbZb2JwHqkqTZKvqW0475WjppCd/UaqaUR
49CTdabXgV3mnu1/cYmU0RIXg4EU4GG1+0BgCbQmTxMRyaDzLrBSvaHwfs+R7jc6yk0QU2dLI2xy
MzMNq5CtGycrStG9nOcb/PwhN6scJr9qhvEEsaoYh/ajtv2V25dz+cYduDIP0ztNLuhWpTN5Exfp
HxakpiY7WipI4uPCZREjhfpu+3irgezpSnHC0q7Q1s6VTyVDA1AuDp27eoY5keBFt5KmyeldlzER
Jn0WRF/2MML3KPJahnPLLl1M5IRUmm95LXCFPiwMlK5ySAteDzjLDrjdkN+Snz+te9yRYE9893Ms
V8hs1NnXJLsgseemviLq+PACB330IxyGKIuthi7id6h9+K0oiYBBP4Ymw7MrWvSNsl93Lic7V4dG
fzjI+ghwvJ8r5Eh/ChGsInCjX9Gun/PHT8nUPuBYyFQA3BWwRwXkhZJyOzYD6B7xUxMF0/h4d6Hl
h73mbfGjHPl1AtulsQw5uOaP5/HZsmHXHd9BeAD8i4UPNuttSVSeJ3468Z4SUWJ+E18PjnRKAAmE
rHW8Pq/GIfj1ZaXIF50YtLLKoxfvRtliF3M6E1duGV4oEC+C9nrPjU5lhyujnxD869vDt3Ch+z9l
XaZtNrRMgdo61AKFRzJWziL6ZxNj2OnehuvxtUjOSEgKtIOWjmtv7+g0Go0l1jm9us0TEPLJd+mK
1Hgvzy16F6gwCEoqPoP6/h2xo0oINGUUEcziwkhnwfh1K2K80hz1VhgV9qwcsRhLFbR/akGAk0xh
GoShPL17sfcD+UFmDiw/vjLNnxYjgYfp2L1H34zznQZ+ya7Tp6yVaTXCR+ihOQBwOcSS+P84Pg+A
XxVao/AGK9o7WvvkfXtJRnZphsDRBeDDA07pVnoY/movKfILjNfYmv6ageLcEcb0y0sOIJG5iClC
e/qRQ+6432YUQRDl+zodwENVChI8XJOd2k1wk26AO+GV1OyK7t2w78EtXuu93FqnnSEyApnMeehE
t/+b3T0g3SdrBVnPJUxgetaDNRHnzF3d5itq99Xg+CYB54877RcmvztX0c4gYkFulNwrk+joGOpw
Qu7/g64+kFem0EWl6nQZU9ftsRmS5CrWHpVOy0YswOC2+6FcyTOsIAUfrJEp1812r0Wb5fzntpaO
IxWGBcQP9hs/3wxUBMcphAZEuu8kv6JTbaJLTz1eYx/MxiT3gdEHynG1IJvf3Ak10Z907IuSeK2/
Pl0agGD0pWAwFBofmscJmqv9n0C67nhjvLZOe2kCrpmu5Y+HW2TfYh0sd4xgRAuv3d+4gaINbLOB
PKlGQDyYRHLN62sjUJk19c4cK92gzFCP1YOhGQE5DvYVt7YvKGqfFPX54YbW4rZPqfRGJzCFdixM
dtz0U+w482eD+TJ8bv0kkk3vwPrQiv/XU7m8DuN1iNvT9wzC8usFQrBEKtxVvJjqKkdJ79B+JPdA
2kzuNkWIw7P+6bVgGHq091oDQZ+lRQifDL6aILyR6xtn2sACkb9JHw+UQGapjJeHUJY1z1JgPKCO
ZYgkY09FaQN+MZ8cfdt1rFiQ5DhXbRfDLgJWyD7zPZctHD/7MSHaMHIcXIYxNsdjcgGWhal9nU7/
XlfpzPzo0i/rxGz8K196M7qnbP7OBAe46SvYF3WRNVbR0q20ik1J+bnUrEyfjwTmjHPc9sjEqylc
z7ECPO3ldSkDQ729IDNV58hgTs4PCzZPtVQv6RgfmSD4dN5UOyKW8JaLf7LlDL0ib98b0q04kwTe
qtTAvXlaqgrYcNbrYksMr45wQllRAfecSjs+RgcT8b0sxZZJK3EqzhS0MFNybZtVnj46DzRv4hz7
D71BZnDSMfrZlJVh4+GhxYzaGcSKJOCY4Hu35wHAWrNtVwy3/0wcQYiB9v8SD6wxo1xnlUNqGAfQ
02Ih/2H6PuDZQD7I3j/UA6Uy+CIc8v8Omb48n6zR3x5Fwq6mCP1UWAbyuaV1mcZRIryg7HhJzh1M
hjWKngJPlZe18OZnuDYUfyjxFougGGpAuupEOTe5bVe+glfEl8avtfNfS3mZwtzMmqZdw7mQyk8a
Clg3WwpFuYZi8KhsWBVu3QTSBhfPQE9bCCj60axzXTQvK2g1p/OxMGPBBWs5cXWuBNPUjCHkkQxQ
35Ar7pKQdOejW9CQIL81+bdcRaGnxNuo380f5g0E9Cs16A3wosdrstRME/oiQnkPHykKFllTSr9g
IlVWHepmJcmCtbcQ5+1ClZDaYyeZO8M9lOKRBmOdhUBSzK76E9gcSLSK9hZYgBRmglfaCYn2M+Hh
3Og0ObXDWXL9/SNNzVxEiTjJ6p2b0tzGUhDueEnTZUi8v46gwpeaRT4p7U56l064WT4faH3OkFuW
FS2dr60qAa67NrkfNMZ5CAok73vNGELcryLwMbfhgXKXrUGzEPi7PXnoORkIabL0+VUS9h1u5TLJ
pOOniFb4GEU9NAB9l+zpXCSFKxBrgs21y1Nr7j4nXkiaIoozZebAsc6CjN9/L2HdPc2h0NqMWqXG
EBx3+SwHCpMa54NtmDYWdfykYzpVkJe8xAD3nGcxMqeDQpKYR80iThsNymbtBXfYNPIbE67SJ5Z/
QRT+4phFmKt3/7Kimwn3jQ2QvIv1RTN/pUxlm9Ued7UM3utXIAVDj4POdMzJhcORYgyTVaxFw4gY
JUsIJyGS89pXBYG5sKjhegiSx2DbiWfKXH+MKXjO21vakgOatWW6BaOlJ9jAM2uS1Z0vMenSJUPd
FUNvrLGLf2Y63YMyfZeYJDE/+sTrhiKT9Sas0LeAXHYPChFJp6ODB5D+IWJoG9ZAB8j+yePaFlhn
HQBT4jgJ5PLPqjXW/hYOLY2Vjl+Zg6ncGAiOhMSXrwzHvd2vwPfmd5HeMtqcbkRm+twHZxKLjzXH
PY3R76ifnDXUwku/pLQH/SLox08e7+1LG8LCBEIpQ1BBylzgxSjltjNbefFB8Z+uLLQ/d0TCihAD
5jLzzKgPe/P8CrbNbpos700LoLgq/7099fdlB2aIo+oHP5d0L1NN8LaFjwts0D7JdObQ2DF5vVeM
yN7jN6/5Ry4cON9H4rhNmoeZBrUDDbsg9/FXp+rr1h3/fNwmG9cN3UzZ8NpywCIIO3VWKMr/XMTV
cRY7Z32IxxDv8ifLlXoqV1WiJU1GS+TrqRJUN1qlhNG1hVfZfgOX8ziMw7yK9NpwNvqJDbhPhwLm
dxYXKtshUQn81ms39clsXISqm7SPslV+wGwa0WpPmGp7xaQO21qxYgCDYqU3HyHEgVfHHCAWETF/
dzjnunOJvjIo7Jhrv8gOeZz1slZd/f1MEOZlm9bLhfgB9VwcnAIl0kD0dl5G4KsDoWfTLDd+Vyw9
dM1kyXc3Iu727ux2Sel1DdocAfNBj7VUY0LTFbtmVHbgMSbVt+2aZPbJUJ6j2LFACeJeQSv8A0QG
a+NftsvAQuuAN4vIrE37zQ8342try1QgkuxnjzqPutMVdxbHep40DASwxo2PWlZv0RLViEjGKhFl
v8c2XF8DSCznfRw7Dq5ShdzRzZKZZNZm53uINqDehrubvOTuk6HKiC204FCCwaRo8+Arb64RKj1P
e4GJbmuKE7u0IPFR1SoHPoVUA9kzO0z1cVjrMoT8yfn+II1QLmvrJyw2Adf40QK9FrOTwJL9Xn3B
4Ey0DFbcy+5NR22J37CHtd5Q9XCZfOdZNd9v9RugDI8AIHB4OdYI3AAzVSgtiRDMVFu1XXHZKf0e
PIIFdJl5DS3L44jSWZrJKus0UOLrHmRztHglfpuD4xSbuiULss+0BK7dgTOFEm5VubP89fH+Yxff
se37CKyKaYlwbroF/kCrcp6tjAI0GEgy/Xz8PtLH3qLi9lHPe+arrzrEw2w8e4kPXxZd4O0XMOc8
lBIgVU+iFpdrnbMQx4ae/3rQlNPxrOhTzw41XsAYTtHGcHP4D7sPhTHcjdysBSIWSe+NZygiF7AV
sW//Mf5eXrtN/tgXMkRl6mYCRbfiN228HY/cxUQy/G+/NMvI0++9vXjbh/oYuVVGkjg4CIOMe2LR
4WPfa9pj238Dn5qR5VL4BcyKQggm566zKGHEtvdc2yDqC7CPLhb34qOd57+jublHKJDa52nQ27Ab
/gyYjSmyD9Q4VV5Kg2QoI07usYJNZ82tmlSX1tWRL3GXuvnaopzP2U75/X34Z9vuRu6Xo8zcSIS7
nITRMoxyEsn+y9IS5EN3cnKZYwuNN3zvpaUyMLVA1V61HkbbKy5/a5c61GrT5lBpDgocB33/hAC4
CrDR6WK7xLdfHU3+Ceglv1P+4dfLcLs35Ed1tSX/RgzfqZsxgo2bc7s/qW430dF2pz4VHSTlVdFB
ZEaJ+LQN3fpbQXtZXtPEXMHjlFM1OUaY5hwZkdf1IPNwCLO9H0mex6OEYfVXdzs8NUTH8Zuklxjx
ST0zffY3KOxJaA3Bi+fdE66sXGGGisRY2551+ks/WgOUyCOJCpC+4nxmEWzqYjxpOb0A/fdTIkhY
3/39Gd/S8sVRRgFAeXF/mgB4usCbfgQCEzB64i8h1cQHvFgwitZqtGRKsdowUkdLQRMBMCVrV+gW
ijPxKyyteaHe/4HFqF8v0DomgzZHQ4GTSfQ1KBPUvPh5mJo+WGN/pB8CM0Zx2RNrbn8AQ2e4B47D
11rYOY9fLJQQYgxZyRuCVEoGzyFy0fiLQ8oJ2ceNgarEqvJ/GSWuU8s+tF+1b/ypTy477uUOS0HP
h0KAFHXvJeTy72K6ZP/qMNq7GHCR7nRdN8HZLyeuE6653/jKLamHXU9fAzPZ6WKweoAgJAefJQ8R
HWC6rFgqJjFhu4PNesi3Q8a+6damIKnTjn33dgPi4QGsztPklD21NU8oAr/LCjOkcjQC2L/czPhK
rDWKQJrtpUYvc6qnYlq5TI97r5vPvW6eqjM2iVuGN08/HGPid9SxGwNAGw/6Ha3oN6FUNtfVwqex
WN7CdyWXvFLq+dMXg1Ru1+YrXDQe7ETO2j6zPAoy1MGZzBp6PKBx1Z3y/Di/+sNpYoTbh7TRXdAd
+xZVuqSia+1AYwctVjxQqvDG5OG/vpxaqf1SwFdt2lWvYNsF3aiHrF7G7mFGbOTfZB9dTvLqQ5AZ
EqktyO0RoGoGzoQJr9Z4KLtAsjDSuAgH6nARh1ecirq4CeBsWB9AchgxBrpFBud+3VeAYrHW+TN4
jcOz7qVRiXQHXwylQnMa4U4vTTtQXtRLgVxV//Lt76bu57zWpfi5mHbVk+MgcuO9Ts12Pgm8/E1V
y87P9ppCO3ZP6Sc3IVSOJvX8jRJw0A8dCWfsUsVQqjcH+i9xp5WYlSohmGy0tZg38X64ufao1uVB
oF32MZJu6i99cny8lDnLaB80+ostzQkGIK9sD/7ouEeGxALCkye3ZWceSaEw/u8BxRVEmk8MmxBO
zGqoCRubhUnpQdlW4kiisNfgdZTh7/Y2J9KNph+E+bW4UA5SIr0kRvfyqxr67o03l/zGpjKV01su
WtGMwIV7orNN7TkOZZSEE71rxsC/Mv7hmKnIJ913c3MVl5t2Lw/F8V75fG9H1ty0olOxQxjXB5D8
RQBD/2e76XJrX0L+wbqi0R7tu/Uxi7FauxYqt2lcvuBAbATqAHOjyQiAf1uevEYH380+PKsScQva
vxqd0UvLsfh8DKQHmv9D+2jHIF5G9NOw/gpmO0+HOk7s/+nzvLgKo0bcHS30Xh53i9I+ZVC+/BP0
Ajw9
`protect end_protected
