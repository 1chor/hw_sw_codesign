-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Lj1v1hwszytWAI9BVqnC6BYmltRxLkroU9QKPsnpT6RqfdoDc/kxKPW71dB9rA8XpFBuF7yGmPLJ
0nX5c2+KhjagPiBwlMtyUtCp9iADxJ8FLZaV066WEye5sQNMoKCeg1Kg/aQo6fQOEsA/DIm6fE6d
aIT96s1Q04PoUGV/nG89YcbDfTRgvdASXkd1JRiI4pSc0aGkNNH9hIjC3h7q6IAbbf/6wz+EY60T
afa07truHud7erua4wbRNPFP9pzWqK8y5T6lqJLN8hrUueN7WtYVlSRWWFRkVOhj0L4WR5ZYuEdd
x/357cMf7pRJvKNfMiq4gADmgyNQsHrBF2vIMw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49792)
`protect data_block
wbFeSka7DVNsqDubelxyBwly1/Zt2KxEobjWA3EbdG2mzsyndpB4f3/o+pKz8r99mQGsVkwK1HIR
zsM4Q/IViTywaBFScEaQ5wzKQbGbgSqB4l4ySyJ3voGHJ+11jK0tarhdv4vh9rEXJgppO2tBbwQ/
hb0KHSic/tIsdKRPLlOXtSUrnmhXjp1xNk6KCCntx3du4pbwLEkLjWdlQkQ4eKzyIe3xe4za0u2U
oR0kXyeIGrR124OlpU1YRmA96H709tZDIp59QIWUN80P0e2/Ue4vGOwrnUIHZfrcQ5g8A9mmfbzy
2jqO5foRiEOIBc2A0goqC0sNrzBJGss6tLDiKHBvWKhuwCTW0wEuWwAeV+5M0KnbU4CoNHzyjTX9
x9yp2YgLDRxGRx5jOSc8QdIyCJwYTwvlRU92ce+KFOqBpwOdzBSOojisVu6YgCNRsCcY47BMkT0l
7JcAM/sWno8sfX1zLTVPtJ65eezkZbJHSXQ2k15onbZAC22QdIid1CtZM2IgP9GTId8RlLjRwVR0
bCgMIHfqdSH7Ee4YXLLGevEon4P8WoIqnqshyhHBRtYAUdyNevCRLJUqVTzl0MhcQr+6kWZg8+/l
S9hA82v5hAENNgmigFsaCQyQ/g6741U+fUE7VHkODxeYLQ58HRdsnBBJCPP3ksDz2JhjuD8OqUeK
kCq9qwynTmvEYzG1E7lwfsXvOZkEzLN9QRWB51q5jxwhVNaVON70NPTFAijAKeyP9CexwMjFkEKJ
ntijppJIQfnoVhyrcm/naQ8Y6btH4BJVBk7zI6zlCelITL+9AE9yASMapOlM0dCAYYyCImb1qpy3
odmY9PxD2MicOjGKlQpGe+4YFbhxIBh+G9uEzW7InhSb35hoPrmAr0VuWBoU+nZd050mjj1sRNws
DGPSfC8MGkoqROFF8hq5YSVbRM+4HebXLhOmLaApoZKS2Q/114GUG4IvdeBQ09kX1nVJilu2yRAP
MNzLyZR6E0saKwD+PhMMF/xnGabucJa1fStUDoFHBE+zLr9VPIwBsqYzl8pypzX683/alLj588D2
P1MxdzKOe5hcQ11jXCZu7xWNsKQC49lDmhcqF/s/rjxMczpXmCLk72uPm4A7xhal+08XjLbCsY53
OWVWGNsM2oN90Xq6Kil91oTeHXTQaAIrqORIpkPmwZiNlww0I5H8wp4yISjR/SYuvhYgvR9THfLx
rdzfHWMt4+arHBnupH1C93kd15KOb5JA4f/0dQLUWEPyoG7xb24co08fDGuVJ7zKU4CBFVN0+yNF
iNhsJdcR0R9D9ueSttavTd0LP2HA1Ky82rtklCFyda6UbCKBJ/DxHkdsOhvdJ7oJrpnuf6Uqg+s/
PY3lHIDw/IV0nMQ40w3x+QGCnHox1ABdHRyo7iUWiBZJohREdEboZrWbt+w35KtMBBeguFq+Cquv
tzPM7p/z2lXdQivsp11XqtuMv1D0HlukzqwHhHVknDN5IFP8SwPldRRGHsMjqZSNrjGwcxSwV3ZU
4p6dHPmfDv5NZl5ZNrEQhKF6Nh41BCOsV0p+Oz4kNx1huLm53w33yvoz0PQPDT07zaGtSc1yqaLk
v2nLPOIOGrJ6Y70GUBjjZ2BjsplBvYtqxkxeJSzOIGdzgzUcp0wUfccYwPHeG4Ey+sqxrhsfZg22
1ABToIK2ac+pmEG180o7T5OlO8KXnF6qiMfa6W5fMQ+I9ej0Ky2WuM5E3H30lJlmNW2xrWEneg+s
sWBnJNL9+1m9ATYRyWU+66yInURTCVNMciIUFvd4737+CKZ1hV3Tic3PTxmJu+SXZS5V275qqkcA
Ii39V4ZAos/nTGRc/SDkBdsG0Z4ce9vl9JEu8LPDOyJpBAXNBpx9+gkpc1prwb2QzyYZ+W/kewHZ
RcT0/J5DwJL1q27XNnvjHY2lCa/JBBjY8A0A1h6STwPEOB8qQrl9t56pxwF6Mtb56YMRYFidR/tm
qekVxU66qPAoRVNIwUFLcSsUyE3s4Ryf/niWap2Ud93H1UsiOMIPYptNPLuyKuzkoXIIBhdIwA/p
/ikGeON3JpfeC20zup65mZwqSZ2feIvmkOHFMJmqa0u59gpuqTdLRyrT72kswGVMWXNJnZeqyg8Q
saQjz1llUJUJN3h60PvSsnoeFtWQzIsyUbVZfppnh+v40XC+qWrOTRN2xW31leLjbaH7Xe7w1u0I
BraFeVceYJ/QzcuUsSLbgl+368zx/0dySg3XQ9r5BZqQmTcTjrAYG1SYKFJfL4Tzs7bp3RcZsW27
RsXOqwWm5kAJB/IHi32W+jktoaC9uTKOnCE5/jOK4fTyx94BUVcJLMtEj5uBoCrBoaXtBkMDbK3l
eUfAsXo4uKz/Sso9JcQdVX70DsOdaOyQEWCbUj2Jm+lBEDKNzPu+rn25Z521u4JrGKSOitdimkvF
cEb9jkfX5xr/kJgX4DI56qiEmNnyKLTAaguZfa7tav8hwgNTNFC7yl3a6sK8TFVDRKx/bEM3drRD
q0UUg0H9mQiLhVeRXd7zPmExiYkPWkFZwS2WOhkuetyQ5OXmFeLCHi+X/10ovvQl/Ey7qmzxEyjH
iwLNDIaq4LRSYMyos0DQ3dhz/M5gfYtRXObNbBp3ktYF51Yg9AoMDhDJCUoV443RlWr7S+68pvZm
bwAGs7kU7z7Ni8hOwTBoOYooX6xWdFGYw1tz6kmMG/vQujW6cH0CeGWQMk07LlBMP3qgauoW04Ov
VI6WMrJ7VtJu1ccIhB/i3XulZjJdvfeS8Ik+bfM3bj1vEieuSV2mZwl2jxdpaBlZVq9/O7LTfQbp
r85KC5dQ/jAiZfrkIcpVWAOFgqjxaumcB/qcEhprYs/eTMCMqLz0Axf+PAey50odzyQEdJjqdsvO
YERcwYhBBqyI+lUhjPgcvLqOFVKJBY0rKSWCJPC7hndwJ1B1X/ZflTWdgEQzS38pU1SMWxFaNxrX
VpYDcNUyl32QpHNU9BxB1+3nTmKxgwTA1PuerdJLJ+iCuP1PHG/6HUVi0eu04tLj9Wyx8FX1Bb3a
M/4YcpNkwmy9BEoZHU6k6MuRYQ8lsF03AVz+xiV5bOu7x0sm+NB/Z8+bZ4gs8+8nSWa7p5uDhJDO
GXJIV1SEwBbYHEmPdHQ3bPt+NZMwrGj8jKi89kSL3ob8Gz7wII0dBRYHDKbh+/OFjD96vtR7ZTlZ
LITv5nk+r3Mdz1SCPMkVJDn6e0k6gNu9bPP+AvtJ79coFXuT0EJsJpuCA1s6KO6iU7pSvZh4gEZV
7NEEO2VhcZm2lawB2zJwGb3tXN2j7KosIv4tlv8qfDHljL9IYz3Lh2CYasykZAiHW9/vKnQjpyAg
GMcrC584ufvjJR5evKrFJMs2+n9g9EV5bTtigXxEXonxAldThTbbfEsNjpNXuPiHKpJmDrCP2zBS
Gmi/6xGKvXp2z+21sptuebRz6mWlqJEEESHBPbj/KxoAyse4R6h3NTOmBkxBo2gZYnKDvhVFW5NX
bV1Bsczd7/HbxZCW9I6H6MoHmy6ihqPYOaLf3G4fy6isNVNvLG15svl42v5IsiBKYsBP5gwDW0sK
odRZ99E5unpPYT2ZjYu1j15ROIl7G5OsvUwVOV4kf+m2CcvN39Xof+IfUwOolf54mw9l4zad2K6S
9vZ/2cKQ4KlC65AIFla/96ct7fkfZpPEbxPE6RqJ6sTnYScKhBBJwCPP9ido+K1PPrbAocAeqiu0
NRDNi44jur4WpDkqYb6F3K4RToLoDqimuf8PK6W+qPLg/+FK2JRrT7x+mfnqufZwxETOGO93H8MN
dFE0ccxWG+m70LIxWkX7PsWMdH5b36A6TrvjHqctrwKIbXgAtAObBxEKkiKu9givu16B63jI2oZb
xtJGiEHAUipYYLXSlC3U4Tzy6ZOKXiaVqNY/WQFcKdu/xRNOINJfsw/Vtx2BS4mBZiMqNC44YAcJ
2bz+a5J7dJSwGRGFTJC3TfLRQyoevg2lMBtHRqm31E6Z5BxIMpRoJbiLxSJ5vHbxwicwwlLpJ6HZ
w4YEvXN2eX9bXxjJuz/A828nhdV2z3uclmidAKlFpilnw4g+ZfMVjp6K8ts/AaboiSNnnI5KHaKE
VmEaKPhpV/Cagwlrdoa3QtggznxS03qlmhxlIRczlNB2qClfrGr5FQOdeUE7qptMEow6bVUOimoS
kTIVDCns6QlQ74cjcDuUCIQK6IJ2EaNdV5+eiLv32PWCs1gjrLef51X9scwsls9QjQPslhzZePND
PpZvwWm7dNRzbArONEeEig5yV5HoHE8/oHfrvRZfxPRy7qDxg32Iu+RdDKlxR8KuD67hRMZXWuFd
g1MNAP0eri6XBuwpqMPC75MgwUjmTFATP9aUC6XpltupZ0oYwDaYpThnPMo5xKjt0S1KlzLlgPPp
3Hk2V+ohFDe7Etg+LF88FOYwZO9eTDLNuSaz1J+oYdQjZUBBmZtvcZnae7XtwJm3QwnP9HYFtG8n
0F0G2hp3BuptXvUmJ8X9GlFrP4Oq//Ude/TLfhlxYGJOk74GK1+zFDQ6HtyUMmoiPFwmnEevOsrl
HgjfXYxp7V1IdrHDrsRd6hdhhSehvQBxMo0fhu5QuMK/Akz0vAIrkEi/QXSUCoRVt+Xcac0vCsZ6
FbMS+DLTu/MaK8ruTNvTvkmS0+6t5hO+tMxIyR7Ep7hu26ubzQ28wbe+lFmR2Z4ZK5TN0Qk2eQvB
1rLgqZOYyjOAyVActANTRsEvxqaQSjt8v3DWlUWmLFxdtmuUdFyLQnCw2DZLwiyLp3ibUXf2jLnj
TEfqMTQc1SnoASUBEE+Lty7hsIN0yAgLf3megzWX3JevHXnd6u7VuIoGxUffMzNKimxdLLIx84Xu
hPOVUL8ibltSQl0lu+wPKs2i++NKwxrDYpwCjsvdigSSAiPUMI44FCptixOeYClhbT6LFA9EYf2Y
KclzUjtxncPKIN3sBGpmm3hEQj2WxVckSaWxUU1Hn3GnhyV7b1M9ZAQzQ1wqsWYajHEu/y1S8M32
dCQfrhkoTu9Myy/zqdxI3v1NhQJKTiNaLvHChvx2L7mz/7jbw+EIusxdk7wVuDquYlXKi5DKwMLD
6bFITpMdNM5dJ+iG0ecF4hPHyMWYbdeoFks+EInacoYVnYT7wsZENuvghJE2ppeczJPDB6Xb8zlI
nrD9g1FebaBg5NMPwh1io3gXc6/X9oEtI3go3/azVxZ2NI96WR3ZvgWRpEdBTbT80vOY9tX9zSVh
s/EDIZ0oz1+MQ2O5Wazsa8koLE3V0nBdhl+FcbNMl21zsePrxutBTXwGgAemj2AJBciWoYDC/I2+
Qm3lSWZ1nLtKYANuF/W6gIuPA9+FfLyxwkr4EJBsnZFWBa8u183m4pMc+lBKujB81bVWFWPFpbDL
bLqcTGm71NCs/12bxRvcYyjzZCatkgaT3yDnGwM93T8PWAK1e/eInJa7oD4nDCA7kiwnIMD01C0a
1a6Yc0LWi7hQV3eBG5O+CPBYAtzvOlecuqJj0OOXADTWORrmiLOOLbr6KIajeBNy4r0387DGW6m4
S4uzDyX4gpXHK6OQblBmKfW1dcmgkrb1p2QlCQ+9FOF643vH8ehYxtB65VVDlUf1uWE+aN/XZhRe
yStL2iNTf387Krwh6sNEnSeXU6s3UlMuhMlAIxsSytZSBxCZ3jvgz8qjCJsHO1lbtkRuw8T0y5oC
8YbIwQVe8mKxuFsPt+czuC+9sy7+r1XuJ29ClcTVLLWNtnHwfdgo1qNXEvWhyD1m5fwwcfW6lSWw
pzsupiznKsp0sOqm4bEU+rLv+5YIsWcbTrTzpCSfsg5or5ysUg3FKGNWLgNBUxCABFk/8nWL1ffU
cjF51vWZEb2hRSr/qYd646uwh8/n4Gkkzjn+b+wbeytx1WWZDVJzKtEix/uAacBpnRLpk055kEWC
NsNtITteY5BEXOdB7X2nRPM8hlMUFKp1Vb6r4RX0UALT/1wb28gWJ/kFFsFWi9JKj7KoUzNKfPEr
7FJ+RFIg8xmJ4Uta9lvBJ4W9/rMtfo3khB9b+9imwLkjS5stb+wVyEDWNeuVlmdvgdnVcSlM6LqZ
xH5z8u3xlCVjO474OBYMIG/eX4F9v7WqbYuYSEUG8hSKi4nCHxMEqw/ABVCP67jtiUOlCL/31bNy
was+qWWuyIGydaXYMlLk4htzT2377AChGQTByI1s2ZYD2BJfBEKZapkx7S7iQv/GCCuHgsU/xkL+
2fijFdRE3wi9SJWHfMBteJH0XtK4X9xmuqrU0RyAZrgbY3QhNIn0yienZe/Zunkp0tKiJ8FNf7Gq
pGom2lo82pjLlqY05OLrSJsBTVQIFaFBhfm/z696PuP4BjYkY+BC5YyD8E87uYoR2ZyY2Ep4KNEX
sgFMXzkKhf6AVOwTnb8R+bsHhI0cInG99iGZSFmBCGIpsWw1+czg9Qpp7DIyXd0z3bx26n/3zsBp
IhzgUfWk7eC1rSLeRMIYqFELdbWWLllsiKIJWpSsvFywhBeDa5JLzIDFzmKec/ld5eTXGAE+dYqK
qHk0wnHRlz1U6ifs1chonM5ME731MV+OfcqEk/riYxiq/AxM+usDGd+ej3AF6ZAkq5L2//mi2vyV
h0zmMMPO0+SRbe7cvDPjCkKAehw3mFESG8RP7M3kQvREKJyOAYYzjnVKigUAOgxWRD8L+WdRKb0f
88dJVxTi7bGEnlNrfjAib7evmJ/XX7NRXTjN6WlVJzukw24kuP48zZ5Ts5uNXySxhiez7lthh40I
Qoa4nNRtXLEfyO+OVE4yOX0PmGtBtPGqp5aFyvydKCFB6aLHCOrTXs2rcaYg30cs9IVaX01PqL8f
Am43COclcv90x0lgsyrfNzCI6LHcEjbVyqnVdtlgItW98Be1M4yx9+T1xv+TZwpTsLlExTNwZikd
VL2xtE1ZtBaDtqoW0349LtN3QGLEgfG02KLlDKCC5sGNHUEFtA0VW8pZCQCKK5G2msMq+CdX6HOW
nPzaCFYQK3aQPBUSflqtff4M7DTDehszB6YwhnN/YNTQvk+65bb5cLPRSobd+oXwVapFTjsOzSt4
x2U6fftOX8oSRK+VExQ/BwL8LQwNQLy87ZSDjygPshO2MagALz7+qFHh0E0JGsdz+V3bfRdg4YrH
oxJXzXq3LaDvKX5H6PymkSI1jynRtfiWVAZ7m2eN4Umf1sypDdrlRrRxIfyUeQTHnpzGW26732Qd
1R5LkmMpPvRczMkmB2sCUINSSZyDgWnZUdKgvV1wzn/jT8FtOyTP+DMqqOgtjY7oMO1qy5lmJP58
Z2PuTlzyhlgaq9bACkPX3b19IehhcLP129gEtHOBVDnlgvopVUqAkqxoLvELbd9Lsfbfa6dKJPzY
BTFhMpjRjLWFrMHisQ+D0XgOH5rInvGSso8kS7HfTdNn6W9oMVBA25n6sRHgA+rGOE4cJxLzLw/L
U+TPVyfCMeCXAMughf6TdQNueARe5b/mHtYqqSIB3gr1A7ul6qB9woaQ8pPFVD/CyQ8n+g/NB0xW
Cv3mW93Hkz2MZgYTE1Ezy9NlTUUs7nQ49tmMERQoTElc5QFqD2+2UsJjjsJxF/HBzmN+9OaB4U8w
lpjU5oiZpl8XTsVc/WDrLXOyzERpxQRMHnrQujFuP59x0bp0OF9ARH9p2hi40nixW6SqpLkmaX0d
bvcANtTUH2ECnqlvQZy412iei9H0DGkkM6kun2pLOWp3n/HYP2ymZ9uuANGF3fTjo+G1wz4G4sRE
FqGsWQs49BS8VeEDOlf5r1QisqOfbhCYfWr4JLFBiHPAo3HZMn0jut7t1/dAaRmr8ZPN6/3c0xa9
BKDgVyUSe4XcqLTQvTjeZEXrWHJ8CWd1iOO7zk2i8ef40pSKhQiV1S+2Y7OGYxk9ahhZFzILTFf3
xFbJ0nLwmu5f/Ezm28MYAvWAILaeAiqKYXnLHft87pje3U/KeYYYeWZ3s//XKihobCIcnBrnVnBJ
iFLA8tnNI7XkjNZFbMpKzDb9LJhOipO6zJYUVCOXulHN/wo1RkZ4JyxuTSer1MOlEj067BPANVbF
k1jMbPDo5f8Tmc3y9ZcxR4v+XCwObOghWvP7Gl/a+VAHLFCaUjUMf11yCTYDGzBAhKG3PFDnT5I+
HxZAyyKBFMgvdqCa9PnlOomnXNbOEb+s+t+AZf452QsfLz0pcL/PVQeZR484f2tsPTvscZ0pPSfd
Mnl4z1OGdLj/Hgbv/HsO4AQcm2/Z2yAcjpNUez/6hW+TVRJfhtMwR2es3wP3kyO8El48kde/zyMT
UT7MpNl5X/5RRi+hVMVZgYJ39qiyyROa3obDHTjowo/mpeGeKlVTNFMoREbq4XlbewlzmsLdtSYU
DgBeMh8+sb8O7XEAWd6D91u29QQJXYbLzHF5i6uDe6n9nR8IoGEz0cnGxeAY2KnTsgLgIEZiBHyI
chA8bqS5VPW2bqpfr96ZX16U1/8zkWZmOy24vog0lH+iRRIZtKWFK/94y9OdhWOIvu1mI10yCwFC
JZQJhRR5Io3WrPMYNYdGIGH+JLJwc9huFf7AJt5ovq+wfn7EyZOkQvyWoPrqDvnXDMHIWaFNt3fp
WkUY15hv5RtlFwVoOkBu8OsSJi5Iy9ltsh8eFfAg9GnhzvOxPLbUKzfUjtaORlY/vVbLoktB650M
mqWLTLrDFiJh6UZsLHt3DO4aDjLLmuzz9JLAqmFDuOIehhOBTYIEdcHREWhwInRxo/1djjTpqof+
oCyO3XIe1ODAnXImi26Owl8X/jpeo9vKYr8lQk7sOknFxogGObQJ+VYbSF+OxV6A7BQ27eMV3URD
ix1pi67W2Rl6mbpDnCdFzsmkMSmKK0mU5P3LYndQyQ2dnlRr+2QifBZr4y/lzf4MW8tazIcTwt9E
yzXx9XTFYc+Y9I2StXHJFjgUKqOqGH7bAb4OFRqwU9i/0HsPgnaukF8h6TtufZvlYKd8HjeuugUu
srWjD5rBkvyN5tNjfyceCZz6nqtRS0pW6KyWuVR363/3w9IjlkgBK+vvTHMZWJOnaBv3RIiFp7Cz
a4B7oJNY/DzkMjefolwRH9f2mlYjmGQb/JpQMnlI3Ttwx+D2x5UMVXUinzH0r+HHrq09Ww16FHhR
Xs8Zdh0AH+FFd0JjFzGGaWsvL8erfrwGyk6gPlbnxrvTVKvh/5UzYYr5i/EKxu8JNH2rie1n0A3b
WCf/0rP2BEGMn2l+Ze02sKdDPOjeSUm1RwktwRLN9YlYnRXLfb18HgMqSRJty8XexvOOc8TtiFqj
5ux1c39tYfF5W5w2PF66fKq2IrgcH0x6aoJ6NNkt64O5Sy0PUzivRftXjqpiyRXrIo+csiGJ+bBA
jHSFW1vuMQM6vUSDauCUQxiG5+qa5gxYWgzfshmkuKoqF8RPgeoX652aiR6zuR6BPvvY+HgIkxMo
lCgfE8uUFa7s1gMOW+Lp0bSmmIOxOtzxpQRKhyGw+Ov51EMBWzaZtnb2QZIU52Bj4swCxvzqaNn7
IHojHrJAmZ/mDLdhiHtMklRJTkPXT5NMEwwOlqjwt5CVuOM2TlhuQZmCZl7EokjCXBoGhDoJUa/m
w9AIyAedS82a3o6d82wNhYfbkZphsRVi/xFCCRI2uLGuNYnZ3pcvWUAysi9/eifM5qnLkDiLxkhV
QN9+9zzNSjpYboVBB+98DOkMPpyvW6F3AQPjaxf7alDs8UiIX8PVpBZTkak5MTj0xXGgmS2K7Kry
y1zKhqjxjxmZ3bGP0cjYqylZZ6At5mhx62SiJO02RtLC4OC9DtDUamRXxdxIwRitwdJ9CcRSXRpx
viyEXszUYZaBIsQKF5xsgKXl/G2GWbKtmk20siycBBktp6ufxo1CUrj0wUjGhzN2RtkgkoA4St3o
wgUE+vrxLAKJa8Qgz51dzVkmjp0iqaMbKgnbmjabctveQejavfOhXW23c80yROpAIS1emYd9PJkl
AMj7guRI8n1Vs2TZZIiuzYdSViyRWXQ/FaGQZ6k43MH9bRNKYXXHovQDVdATdtp2m6L0Wmh8pekz
FYiEXtxo9RwB8grg5AYgqKTMpDn+pyLJPQzJKhHLumF2kxG7pebSx2Y6IQQvaoMIJH0s2XmrfasQ
AMLFWaGLquQUoH9GkjbnlOZSFrruUzsTBhBf/eL/PdoMAG7I52vLaOtScRq03UFGB4U+4D4nWZWJ
9EnIg+nxyKJSiy7Zi6fPyW/nhQUFxii2lwX8pEtDILM9vWDWg6lDDmMMjEjNUYQ6Fa5egkV/aYL1
aEKFMw9Od3AQ54OZ9mT/uZvdYFUxAxExBwHAw60DLtkZ4oovP6oCWZyJMpi7DW4BSCF/C02pU9lG
RJtEKehGpE6XbumlCQRArjV1fv3AJ+2eJ/gsnTlqJmbQqi49ImMeJqHqdrrCmgfrozMGAZOSv8XA
0fS9Ym51tYSGupMubzI49zWSlCbcT1mWg5ej1Wk5q7i0m5m3FyomJm2IXesdvKN7TfEcXBKPFeFt
vLs722w0czr6rLz9Dmu+IL6q+ATVzchhTvmItJvwAlIIYNl0CC8w6QpI2a//3IkLiYYL/64muRde
oGleRfRSHgOazwjDZ4gkiXx6/s1QLuqn68xHIGijD/OppuBJjhycs0iRAD57e1gXn4a9XK3xZNrb
w2YGyUKzIuceeI86GNaM9E53KdACffsL+EKQBVM27mbYBl6zKGztZP4nvzLBd7zYM4NlbPEw2PkA
+THu6xE5A9NYk76CKWe+Aje/eaPaTRCaOyvf2Tdsvo2HW5ChyzIN0GapoocnDV2264QqqInd1DQm
yxZlAiFEEmA6dvfIuw2ZUrK4i/DSPd0erhgCG8dP1pY42Nwx0FyxmvdZCg/dNBPRL7+Q++U9h6kI
tjrxh8ZI72dhJ0g/3pJgUVmqp+zDMj8EJnnre460lDtWCU9Nw7aswjs5j5HHNo5u/zG8kiCMo7Nw
roKoL6oPFrKRos+601AwZ1GPBv043wlhjvohwvpUm8a/FUGLX9ICSr6X1UATRSd/s06h/AJWEnN/
T5d7m61imGDeYzj6X/ym79FPwsBh/WWmLb2PJ/BADeatUl6XeUVbOizCRUDihAxKKbA9IQ0QCl7B
DN0TrBwn7o19MG/dj1nSAJcRBleV44tWUHZf+itmW/Q7K0bIPA5fVYfi2R7r0iNdYCWA9/a6DDxb
gIF4PdID70GoxcgLSv9bmefmhNtHqtFDiIRnyJVFVZXu3x9COrHDEVautqUu02lHYiFIPA2/xh+U
eacKw2oEgfPuCd4KyeHFtUlq9GI0uwk/uZFEI5RfjII97RjCTw3H4jP8OGL4d/728dqan/SsbS15
34Fa2X0fDH8QTvScVD3V8CIuXzG9pKpwHLZTmibNa/lhWihEEHP8aJFFiyepwXwUPx4pLTOzlg4S
TaM5n7sEuoQwj6g59x/Wfc01LPfxK+MJVJVdTUVLZSN+xyaSAQt6x/M/iP5MV6nwDSt8hqsmNJW0
sgmXn+HLt7rXdcunVVsKFrCmicPULDsm8fNP+IL4DWyq7ZxFpL0M1N7fVp6Vb138a/6rDPoYY/W3
1KsFhrP+6vQelfIM1XHBqWpVn6CQxTQEcy85nGORQs9QUHe7Sup0UJVwqDKxuxSB9qz6ACsHwvbH
Lau+2OVBYBVFE+Xt6flgFVKCMxwcOUd/mvMsuJqgurN/5GB3cf0ldyJ4J0ACi3CxI/8OiggNcoJe
zPKeQEJ4VmEHMjBCj/O45jgWnqen8PI7ynF2juUCJnuCB8aEn4FfFrHudy55UBdF5fvU8QBdozmQ
KdzJ5sXL2SYJY5QBbSG4mSVT6OFJdjnDxuASZfN3to4D56TX9bx/PaTiMAplQAeALFaeRKNItEZT
uw6zOBJR8nMFfooB6X6eAy+psg3iUcb99njnYBbHbq/+AfbJVYCbvrFTur9tZZboWZrvMGwzi9tP
ZAW5O4ujNWUDhPV/mEMwme9GKylGMyaAqaOk7p7Nkn70mGUgouwP84IFiQIeqh+LqiXMwFRDtM5b
FRRDlpf8PZt6TmVrfhYx3zUcrmCuhMXLwrWjhvK7p78ktrl2AHZGcLlFL3/oadp23BdxqsdPP34u
6JGLosb/hiilNi/4P1fz2hjzq9XryXHKB+lyZRCQ/QGmN6bZ2RY+XoTpNmLeIH5WCgVN8j4KfBol
mbnZQLlN0TfHSkJSEqKSHNlvXdTHEmwadyz6DXNvatx5bpQ7k/7U2Irgtx1qAVfEGIvDVIP+r6jH
6Lge6EikiwEfVyMpM3Xi+NgEXIdvdpgQGCNzSAevegkfiziBJccyB6HS/WYO7ltb6u2HZtbNgmUC
E+8BRkvSaEeHxmT7oZ8ZuYfrVwREhmlGwWXEmW3xZgfySKuOFLYhW5ma0qLbKe/ZPH1fbqyOwUdR
ZaYWbKEQ19U8Use4v0EhqZ4J7a6H4ASizjczBGkl8Cdii07nhivBwXc4Is1joLZKYMqla536lHXh
LUDhUu2/hGgVq7Uv4ri0FMBaEhAliKCTqd1j8FH6VhV8t1YH4b+vxJZB6oD5F+ICgT2+QTjeR4c1
9AcsmSvi22Ht/BkrFPYA6Yq7jsYEhC3xvCNMkhel5iIkkRWPGAcGdLei7wbqVoQoDL0dnzO8ey51
dtB9m24TZrxgF7JuGORQUS/iQr7rKe7EI5X0KRMrieYBjEM9+4R0tik127xvRwzAgia4LVxz7xFx
9TCVZVk4L8Kym8w0kMpBd+keATX7LgDT6Fw8O5EHml2VsBWvaFmWUGUIssFqPSzYNSysY3yV0PIJ
zy4vTSp3/q7xv+xjetIksGyU2w9uIowVGQ8lYDkZe1Iu/OqAj5TMstLKFOEnQaB9gJxAyZ07a+fe
7sbJTJimQqeMQ0nMhIcSdj/u+5+fDIWQ9w3Zx2sQbgFpIsj9PvcluRpd6YRHOpYwLRxOTY9p54fz
Aw38AI5xXuqBAaLrBF3K+22zG0AlOr4bHpF1Z+yfCF28wue704QnYjUfOP31XZAx8y12oKlGPUs8
XL1Gnng5ntFZ/DeZCJrx1Qu2dqQTk54bA5pUkBVyA3H8VWWnn7UDzfLny9U8vcBf3XTZhPB5c8i4
OsiXP0oiSzYi93BPzKTWLkChvd4YVbMEJRGzpwkDUbNSvdGfZW8ST0RLlA/pXk2DgL0JTPuANfgh
Bm8BvMYUDTsE/Z3fWJh4rxqDN12lXTGTS2X/VCS3CNy68G1VbN1/Ah24jwk/WSc71DPuzgiNbg6F
1ios7VPwSCGHTTPLz3v7Jx7S7Drmhen8QUu0LRzIbgZAmgZPGG0SvjwdBcUC87Oh6PBPAnYh9/Ei
aBIP36d2TOzeHqfFxzN37aQi88Yif/aPDN0Z87vSErkBvrmQaXQ88crKpZq/8vs+8zpXtIw6JsEj
OE/PvyWMSa3r/DhIWDsvPkaGtUl9z3M82foEScZJmTw8HhQzOH6AGvZSVmtFEhjmip4cKGnJcr4T
4lbhD3il0JOsgCxtLhyHtTR678nMY6M4/jD5QZZdPymZcLztNPTtWHcYOl4CooetY5RPfoxOjWfH
hL89hDeDSVlukoBxYQzLoLrf+tSyI2myTZIWAipjxNAeXL4hg4Z6ADY6l21X2/DXk/whD5cNVQGr
mVMcR5dAJc1u65SNWKXY6r0MgHhZsTvU7PulXYNR+6ULbvnoAuYBlbwIGmY+X2CscCL82WnNuCFR
yZQ42qKG1KFKPBznj5jaa5Zpk0+XlzQ9x2cFdTAsqHVCgH6X3ybRK0V6u75pqLNILTKzk4M6lyEI
t+0sBJVVkkXjhRYpTDSOA1yJtzzjrGXQxGCB8Yrm86Grner3Nb2LfRe0h7zMYiO5qsucuJjyvhxA
0sTPNSaPmduwYmuom1WifRDXfoz3CgGu6If7ZDm/xfydlJsHT3hwf6+ePHUH+k3OTgQIEwhSJ92O
sXx1DNbqb5ur0QIsrSH7MN387ryhycKfKJVvBA5e8/Zk9rF92VQO8/1jUEvPaPbuKwOf+qEmbuBH
cC2/2Htq9K4u5EX4+2BdjsQsFjvK26xxtiArgR2QeJqUypGYUK42RvaLAgi0egFzXdk9qs2WDECi
IUu1gtuk6unizH8ayGvEgKA6XRqAaS2bUDVaBBSZtwtiNJxn2A76yQHf2k9IslnrXOn5hix2twPd
U1GNtGQvgiO1q368Zc63uJ1WxYoudB07LiUIqk0PmrR3WMRBozMiZYfHt69G9uyuUVINMyPSdgYp
F5k5BZdHbaf8w4rcVCyGl0OyBY/qCebrA5q4NEqPN2nVcNoWp2fOhQF7ju2hX3DoUKUlfuvCc1Yx
XDqGBCZshOoynGDBvk3uZ/9bkXzQhjugl1q+WkUzrbtOq835TXeTjl6PJW0j38Ozw0tAI9Ai3lBH
DNOj3nvpncvXBdyp/hZLaLWOueZVPo4A0ogd99RmpvryOMAww3zWFJ7xMNmmOetuEqPFaAiPDwUT
+XEbMIze0q2J9wyA6FSG5/CAc3oron1vja9LMUtEyaHriU33R756C8fVie6m4WNJJaeIluu1Eg1A
5TQw+bsQ9ers/1mS3oCkM7sAtzLts978i4aoPixJiyRHejYbKX05ixMf/x8QlOrX+BEGDhJrqWfu
u1lmNGOk3xiva8VHIkIUXxLfXwPFmDwpmz2M2N9BsXG2ZnKZSGn1BCPEeeyjYir6WPG7WCGMZnIh
oJa5WCWhpywRrWwTVP5kQ0N/dvC9EjWGZz073HImMRouWX7uvPOoy3iVoS6C6UX7YoIUkurHpy2E
gFLJY5ehHOnYZVxQqDBn6UzRMylBJUx6yc12xNKSrYqCJotLy18CJ68oI3kIExjyFsH+P5rQAKkK
CfvuxuoOV+LsGJkOJ7O5PSfyJZDkKjM1A5ZU6LmYzHhs3xjLLnr911JzxwJLDcWJMzTg2bYKjYj1
MaswCT7YCxL15mPsvYN6wyxjth1SbZbul5+CrPYb4CsS+/3dTqHtpEsdv9Fimy9k96qXgaUm64qW
6sm5zRHMIFc/DfyiXFfZ6OXs2hyqx8EgN1Y0+lB1MR2SaSZyIijKIXLQpzOJkMSh9M5IoJ5C/DzD
7YUKdNM65pDIRGuqvi17RFG60P5fL2NCGq1+7T2Ca/lMo/NlEuL/h6Ryp0Z1+4dGW5gKzzAsOtgj
K6fxiNzYtL/yiSpjsXfLvDj1OE2i1dk3QL4I4l29vU2iJADU5FlExRgTo6pKsboStKIf9/tCgTRZ
R815bra2eeiUPul7Trmn47qwZr6CWXbifprUw5nPrP0nV0ZhEyFUOJd3T9lvVmkvoU7z1CMtlxiJ
9ac3Mm/VekfAhXNExzSvg9qMwlTJBmu7+YZtoPHAy1E5UnZZUnsDrrGL868OKqKRynpCnP66RwZF
kdYCsZ2JA0CCfp9cX0bgBGHDp4c275+tndjRRLraUmPNoQYfyeyCcXvcSi46f84Tp/vVpC35/b8t
wOCY1gDytjQOUah+/Rb14tsQkceh8EbN8BvxNV3Kix+1qcrLWlvoM+uxIw5i7T0x+Zq/jUYf4/Xy
k9tBuaSjhU6xX8LQUX5u82otWEZhuDj+HlLDge3VY8b+on3G9OM7RKRT2X7eE1b88pMlLqFpVJ74
mi7O4/++/Mw7UYn3XhlIPb2bDX+O1koCUNDehcJqTAC6bYVU49/YgN0FphdCDU8ucO+8aKpxC/8n
dwFxEe19M0SX4p1kH1rNjpCrR7b8kdwXV1DXOQlQdUlfIJ2syIV87+t2i8rUpX1tlz3bzdamqqb5
d9YFX5ch4YA8ecJ6Ql324aXNd0MpkP4ZEgzVCseFUTeM+hPHIBGTo5OWVCrmTCQuEcOkg1La3ZZK
HMQWJr84g2bOdXP2BYoawM9dqHvFtqMiibXpr6Qsvb1Ce9CTlq3z8u24A4I99fnmgYIMv/Xu3TQz
kfC1Oe9kkM9bgDx1XZ1kTXYfI4OP+wJMRVApFGCUTJOKueaEwbrqO7Q/B7dpnwdYMYjMwNQvXj7a
osvg1V4dJvco4WNWupeLvNQGjJ58Tw4fe0DVh7Moq1IeaaOmHC+BcsjxaaiIBlSqGp1OgPwaLZEa
a0+sX7+1iS173vmHU0hMUxLJ8yCNc20Cz3I6TGmGDwIFvPVYFq28Ob708myyQEH0Sh32tbmx9I4y
7AZmEQ1BhSwR5a/t8wSJBF0PO4FVkzVyqp+GRY+r8u9KT8MEYlYGsAEerpwgRrXyt9HGB7mqQZFS
AGx6jPt97cKA6MMC3Ni3UR0PRvig4aHO8caTbQrqEaALe5U9mtpFXuyYannawzWiyp8q4ondyMcU
T4E4wS3+7sYI2tBy2dz+NwMk5r5Ei3H18CQg8rrQoLgIS2eHbg6XO6chHMOkRb3CWL1XgrDW2DXb
uCXwezg2+O9x6ELMAIe27GuG/7KyFT6dfZHGc4LLk1KxaG2RhatzJzgP/T2N5OFrsRNCPxFfHQ/l
NvvuU+NsIFBiBZtjmD+H2RpjQbtv8/OmzxjR5bTIpD4VG72avjUGjNDWfFS/i0wsarEjbI93n/FU
tdi9YjD3NAjXdomFHdRiQIshthr8AmjaBJthUwekWrdxTdTyArBnjRCVXMH20lhhqYGr0ehD3luy
xeQ1XqSapVulYIU4KQC7h9N90I2ZbzHFX4tc6H1b84nnPaB880U+yP8PQEVcxhQB9dLL82Cn8i+z
IMy1wyE566zvfHBo/m4WkFPpc2L5zpXnLmE3q36wWAeG5TxbLUshnsKwnvtsi+sMTZ2d7PCouu07
3fFFsRU+EQ4bAnadW0VU93EBKjSyqxEOxiVLrPy+F1DxdaKm4XK2J8DDJ1V3DeU54qD1fZBrypY6
RKtXTxnM+sppZGEH2jBtqMLtr7yjhCWN7ahm5jLQsCX+RvgtFnam+pUOzUEv3PvplY0oxJIJEkgr
3ZRThnzRyj8Qg6JJ9LAJB2/NX9dXLyXbuPt4wFNYTd7OW7RWN4doj8/rjGS16LaQg/nrObuKjEy7
EMXMjJgNRhV5dC1wMd0ZAoYg1fo65Dxti/crUPa7ExfrU8ouVgLTvfPXFT95/fiHJYroU7srVv4N
KJwxcOy8iCjhfFPiTPepoG/yYx3x8I7FmVXVsAYY4tRC2FcocONDl9LetiiImOTxw2ct72zEYzCO
hlzBFgKpSH6FtaU5MMVoXMdtHOgvLcyYkQ/RfTq7QqfKZAH1E3uPbT8cK5JGUnDnerQqI63uPwwK
sjO8CVfGctq431wQ90Mk9DKIcALEMlk+McH6LPn4GDjOep55atiudy8cvCFhbYpv7iM0JeWYgRGa
VDFyxu4mmhvzxpkAQzu4Jaa9DdgIosXvf8VuLh1d6v7EsLbqtnKTKfcgaT024GHxA3Flun8lSOje
yTqhSAabkm3Jxog7mk8slLr03lj2A/fzWgT9UZ57d/yXXcJ/F65wfUNUXICSZ1BeefkWeHFyNFG+
ann/Bqew4GxyEKL1VXZuSpCB/sfooC6azsiAq0uTkEnOOeeZ4fgVyW+iQ3oiNAl7LOSqLCQeyyQl
xLl9khOS5REuzGmTEDPdPqN80RTm0zLPmD2bNxaiT0CXKXlrX6zLYKOvoiRSFSfRXYOrelr+NuOL
qK4poIithT9/ORpoyr3fqhofoJd3yl3JMA7IudlOY6IdIUYP0vTora3Y5KxRY54JHw6HBMbYazz4
bT+UP69i3XNzQ41grZABxMjST4CbBbleipBrVdHWOODq/dswTj6FcTulajmlEDHyEf0rYcdXaqeq
odiJbE/giZJk7TK7x884/7BN4md/r+XaeJPLrIezm8BXa3ricfpCORSlOe0hDKINUQq/eO8hGh7N
goa3ACpsbJFboXrd+HVNc2VbaXh5100I7oOf0IGz1/dQ79zwdXI6EBoCwOeM0JxRbdCfWuxH1x05
UgbPv9JIddRwpHclGZBOix2RFzOdlL5QH9Aon/AkaHwM75Ro7s7DZYTRzQ0R4guTXkRH1S5i22sq
dVoD+XcW1QM1zZ7xX0GB1a29zu3NLHC7Fv118TQ7MdnYTBu8DqFvuio584dklJCKxxiC3M/cr90w
DrLdlLb2CLvtJYeWwnNFZWSreKXiFZmc+8nC+u21D0jlu+MzLVoDaKEsVmFkvGYzbrt/f+x2Ibyn
dPKnL7uys2IZme+xgmANFoqVGYjQSUrHKj4cuU8dS+m8l3Jo+hBKrrz/C91uo+KaBtfJednulcb0
XFIWUlDQ4Me3OmMiTgm/M2/z5FV3NRMlHLjiAXpA0d0/6F/HAFTsu4yvhOFTF8MBOyAQKgg23y8/
65b9Cq7fwvrMDKsKYNUIkeldHrUW/F3RX++vbL4a/2vJxZOVSL8v+794A0aqhGAf5wf4h/ZHtEKG
a0gSWHugdEb4ga6jMeaXbcML3hDtyKQ+tPLMVxi8wkIyYNcQvDdFYumdgr2pl7donyw1MbumNwza
RY7J18l4RKIzxAOkNHi7eilLKLrwDf3oglKMDMPEsVAiKvJJ2f0f/awKoN5+UYPzJyvaGNBxjrir
7iyZ+NZH1PBnnosWFmRJhGiANBn3A0NhrSpWfFXP3pbo9CVxWEjE17IaATg6dU8P6I2PTqXL9too
Uixw0gdKEL8Xl4an62rbMfXUhQlPmjLpUefJV5vpgNEkDiNq8s3ULBApRbw5IQM/Zc1Rg4phaO/9
TUavCtR/iQpOGJ2yQAtvPtYMx4JEO6/Tk1M+vI5mbk1sYRv1OGv7IdELZmv820o9qMBudsnYt3YT
uhjZB+lT2xg6Vumya5RTcSRlRKeIpvhVpZEyTRjnnqUpPyLlVGiXpN2YJ1Xp8aTqUa1OkUIWf3CA
/nBTBtqiSHAyiEPfob3DDH4ipQIvGOUAk3X93G9tcH8iDCpT48ofdj1O430lfT95aFYAqqjzNUhY
LKbU3lmxWW1CoTDmf3p5y/Nt7lJuN50AM2zr00OzWA/2rej4E4xUH3/2HrdITMlgu3d57lbB+uIK
bvotSHIwdO7FES/wCvl/f26NIoQzEf0c9tcRlZUJkxSb0b2YjoKd6FVwvr+PT26IYZFFCVMt++hz
G7y/Mhx/74VP5Yz9tiWyID7AFmj1M3/kD/Clim+lwyeCFstP7XSpEhqZNqhaCLQeklo8hTBoAD6G
CHXwlCphoZ2PecVk7MKlxTn0AjDjKkWQYxc5QkD62hZU1dMlnmvF7jsTOjP46DboPHKEk8wdTL7+
qIuMNDQJeBvBU8d9cHgBzmdvr+nSaUJnBrNZPcJ/7Ho8LmL+Dipc73JJSCGcMjDPAKgWggYf66a8
THA9J0P9yb0mH60y55P83WO2m6eqfRbDYMSvsLHPr/ZRzAoRC+UrU3PfUf1DZydrQNFxrdbdhLPq
QBBNbfP7UcoxRTauclN0Y68sbwNRIWdTADLmoNie8ilM2yAMjT1eQk9q9JjvnJfhDlHDXmm3lxCC
ie2I0laMVM0z6ePmDECmeHJo+2R6XpOyR99FyTdMvWkel+2lvwVZQUJHnvcvbbNaH6eSi/0pTrDV
fdjXdafK3QRwhxUQyMUf/8vX5HQdQtT83ghR9VEzu1HDutiymWincC8DCuatsTZZh4KEFzt9P78S
8GeudDY4JF5aHZKnd4qZ9FiKJnIO9KZTYNH7FQIN8132oGzmv6QNeuV1FdpZAkzdfj1DVT7c8SGs
Ih8BcRdoKr1qVv6rE87Qr5ZB4l00PV8QdTeRSa/PSo/YTks6wbq9owpF0HRGBssWmmZLkgKeTq7W
Bi2RsWHZe/LkZRl7nhnM/T2TQ4QmLHsNlewbZZLFwAgTRVqHD5fAKLwhFJ2fogj8ZKuQRCXJ1HEh
LGIU7wqrZRqHedB5tZtfKfPHNxT+ZkXT5eNggOyMMlLqKyCewo3CW7vX1vz3/9s0lD8qkP0aB3fT
80tXiF9L1fNkskwAaS4YEl54fNZ48CbcDROnazn61Mlss3EcdmjjIrbZd/t434zHiyc1A4rkf+e9
KxhIkhHxp7hJU3frqQrkmCQbEz3Y3CmaZ6i3koGIifKJ46X1uD/91PR2kO8vg+uj22ewXX8HlRXa
tjcdWvLfiF33KfqL202UyQDbWtC2iFHm1r616a0WWFPK/QD6Ugntb0kxfLmJdsCJNQ/8hBTvcAMP
ExDUPItEI4wmNNPwh2dZ5PVAzQ/MhMwFFXX/Ox/gGuGIxVNNZtOTlYX8tfcqZl8W3ZTM3qRC5qXw
6e5nmk+Czp2Jr5V7pXC2EzjCEEmAE5H7PzBrI9A0esAl3SQillvpH5QHkYmAAj4DlCfqGo6JLzK9
53IRW2QK/hKDze5HPxMWJxUcyplK9zn0jvHeDwLANPGV0PQhnFZbpTDh6ctc+0HXQH9FtUUvAxbs
lprgC/JhafxUNYisB20UnAv7B3wtYf3fM3zlpwwv8KMjtbNk/kH6Xp+zb5tEdVWelnC2XewMqHUF
RbLvdmjhq1+INufhknuei7KjbKhaUJ07WdHK8ypviqjTe9Kn4ncIe1LeghhUaH6RdPII8qpWxONI
+5YGWw73Oqr6wFrARjqeMxb1Hh9gvbK05eWSNn8F7c4wcNhWcnLkkZbo+71erzQ5/sOAXbeG5y7K
g0hLiwl3SNtkqCKO1wiNOqtqs7upSayneg41xawq+5MmhfM2K1r8pKufIq/+1QtnW70eojUejrX4
z5bkfZFQ7/UwK+LYtPQHHUwQgpKqBGYCw9MOhGPonlTJRqKbc8zMZ+agNaFohnQZsISjgfKbUn4L
d5bTM70y8nRD9U2awwjc2ndtM10QNalmG9u2H08lobmrWMraKYklYM7cobTX5ATEJXP0M/3mKOVH
wRyFzTDbXc59sOb2hMtSJ1O5NFgE+kl0et+8wL14wrnE3HfWoy+wfPIiBvO9mnKGFHNi6zqULb8z
E5lrC6WSGp7l4Hy9nVYWsW3mDIUr4jIlgbkeEtptr2YTy/H/3Ll1FjHGn9LiCGHO1sjRNf0QMuA8
cV0oWbxbk4u5NLalKicuXnvX1LZizb9kGpWLIGlQkogrNxy2I/iDzKtBmZSk9xmKNM7WbELsDZuC
gECI598c72ISxNvtbWea5lEfLBBGsrECsBkYb6maR8be4V1foBQM1VMixuDMzHMsr3OHIg/L5XjW
zhqbm9hbRv+eo0VYZUaR8b+qi8YnQpKTSx5Z6FYaH3o6CPJWdUxBRKN8+6EsbGdUu5DQe2AqaNuN
LE9UPZee+ylY7tSzn/zm3Od4FDva2k9Qrl6gnu1jeU6ssBv5whCDs7z4rPrSwgsXFEIfsrtoh32I
9ZDhjvnRjknW7ZgSJnp4ejfl0WP6f1wJYU3sP0FxPV7gSx9wl+knG6oF4RqtGEPkbQ2pyvAwMivS
wjl+6631Ts9ZoVGNmo1iA3SZLrqZYeurqgdzco0j2F9FHHum/EEiCxeBNMfi6jHP6vq1B5DQ3YXA
VbLRmlXZBTKv9E9Sym2bj3yr7x8+k4eVYCxQ904XCgIFCzaWn+2wU+IDXWJ/Lt2mecGhmGivKw1f
KQEAEsU4gcJcfkTHNdBfjksfpatRXzUhc5dIctcPq7LE1OK/k6gQzeaB/5bv423RS8PmfVYFxf2e
KpIcArKdRFzkZm5cuGxkPqFCV3Mb8HvsaME60bJrqxsRPh1+7prYMArXfM8S9lJjer8Qz5jCX7KY
E4iki4XJdEqo3c8NjMqoVKLs8mRJfgVaIDrX9wOXuTgn46uVWCE7nZ0bYPe5jvJf56nysembx9/o
6x+PFCVZn9X+3xZA7fW01dpgC9/J3hBm3Ui4UDawNQReYBMlKFz4nz26sgNicGzwRH5uDVI6jVg6
+sD90nkxrOEaPyEeXSiUNHESw2WjxDpZwNxz8RZXYPELgMBbIQeatoQCyuDC2XXpePGCifD635dG
UBcs+qh6RyItraR/dgEe43RQsahNXvZ4NB9ca9/gE/xoJT3DHYfR0l8rP3MEHhLcvWxt8GWBJXWV
5n9DpYP/xqho2TMOgyOL3EDpmL8RgyDxulJ+k3RdwiHjbHRWas456itbsempcz/KvgCBNItPY3rh
ZdP0RaEDliuJoizPwtZRMqjwBszM8vm/JHflcUWNEc6wP5vmNXgHzGvo3Y8nPWl6uh1PoBhjIuPy
3tJv8waxQO3j6F9iJJynON0SlhGW9txiYeK+/6i4+rkHUGn1bmGLDMXhzCpfdNev7p+wZTtJJT24
bJRTyfc5uAX25gSud+T72aFmDsHoMe8nP9BAyiO2OmcVwzZsaGCSMrirvh2243Q4+DwNmEjDPYKV
dc0w0+gAttLu40k1ckbe18uRQtgCp86F8J3OfkdX3OQB2C9Ob7MkgTffX4+qKRpg73TvJ2Nh3CRT
rfKCEpqjNphR7QGwm12feyZTl04+rNSE5p2+8BsYpYKqqYu8hxBpgztqx/6/pSOfDh5LCt/4tmEW
RYBEQOPdKtLYJHiKYVUq52wijwMC/m4swcZOFfdvemkQJPN4M81RkllJEXgDr6aPjXVDr+ObwbNg
yUMc7Ff3VDfS9d358RN6uxuIN9Kj3Zl2GI5D/2g+f45h20Yqck/m6qAp3RK++ZC4oWkO1W4MQP+r
eawXDIBKZCR7Ex3gdYK4XRwRTtGhTpziWXU+n0r+KtjT2m+H/8Y6VaEb6f5Kj11Alt0oo2LmM9wn
0K2C2QgVTHpWFjJt3ZHhxcotB6C9PoNp4QHjRX1s4yi+3RbNqK9a81mzWrZY401imn/itn7xrjuG
VolOdCA3i29cdzYkFWwVnazPPCD2ZfezEKnwa+Rb7tQZHyB54RrxGknAZMcYUhU4V15FVLmeeEcy
RW6Emil7Noy8XKocwGzG1NkWqHgR5p4F1NxiJU6bZ2s/p7lRGVbH8dxmt+Omg/Gy8umYEoe5mjUO
VUgVmS+wqT2tk5JAQXaD2O64SDMBQsfg6JxYVR2lllUjGTO9/eJyGzRmFDDNWqg6ti2aKd42CHfw
BSHgOzyUBcD56dZtqtoXPtffP0icgZjGcyaa353Ga4KK/T8rVjZy4mAbruZcPHyLZfzfs0ktoXQ4
wbI8/bgJqYuwazIhr74dJihRE22VXnmok9DJJmF3CGC9IRtJ+3ZfPqG4QtCrCoBbAnIurjUG0TfM
UrsgWt4Q5X8vfsJso8MXmzePFQNAL6GFyCaV1raGNigjFcq8mNQnKv7tOFZsW9GCd9v0LtzuWyY2
qJ4TGwqip5eLk/J2qAJre3Pcu+J8Osu2Q3FqmeQadng6Flbz1okGUmCbt51a26VU7DrCvDjQU5jx
nfKeW09Wb/nMoN73anCEWwc8uez5INe8QFc5BP7KX1U6d8flQY2T8LICgpkFEQwI31febtdUZPYG
5SL+E+206RoJIoL7dQ+dH5G+8MLgjzPK72El7zAq1d18fia3bDN6r9m7Q4IfJvadq+fRoFQoNAPA
tmBMOSM8+Z7cpWL4P/ffOUJSmbJ2vqzBZ3n4faLUWKAQHhPdXjdxKvcAG07cho8fYu2oF6R5VWFg
O68F1uPMor+/VNW0BysQqM6IYgsuB4LsS39U6WwyY8V0vYA73BmFYG0ypIQjyoPorrvdzKqAT2E4
D+ehzqsbSpkZu8EYXB35TGDcpKoK+JHAPdF6M8dYzfvSFeDJMJN3Z1ao4NIMmxgo7IpuGI2a4l3d
fl3A7vDdp4zOXbRFKyjUB0VL9+BS236tBWJQoagAiDdqJBz7isNRrysYDHAd35n/LVIODodmjCeV
G+mMXqBKiPC0XxCqN3Z1HyvojlbSGpIXM75uwN5f6I0SXQPLMpG2tzVYD+3LnAcESSMgmiOhpatQ
TjREcoVUauGnuTW0h9OL6zXxltGWxhPDm6zFo3d0e9DK9KVnX8CnVruqEGd6MCqbPXYxDSBziOdu
oAAzxrz1Asw/HMKPkeZtg14PQlNafprbHf6kjn2EdBujk+sTHlyT1/+RoC0PlVl+pHKBNCNBnRwu
sXyWlD5NFJ347uHfrhXw0R/tqQEuVM7CdJIi1b7rY7AbazAxtt1ulTWhxhiuB0TXUA920vmcemtD
BDwtYb4oM6yWmimdwzL7FbuI171kgSsfU+AS0b1WPfJkj2ElybNqywJwfzdaBZTLA3Z5jF0nAn8M
2r3CqA9CuqDi2dcelgCpa86dPF9kgDZPaAXFWRgyuGHtqy1108NHcxPwuAbGQMfotmfNpaLGKg5h
7M9EotnFVGgUN+Sfg1TY6471h5JkiwvlFmfKvdA2d8CIoYKPTqx9AeeIr5MEueXlNEgCOQttOk0G
/OIdnR399q4WdSZ+jveYsJkF+rrNDMA2r0JLaSigOISada7NI9nLcqh9r3ZFQ9qpcMetRor3GFFD
mSmlSK88dq3LvTN/9253UNVFFu3Z+0VyfQE3uM0DwcLhGxcMJTbA78yd70e/fXubedwTYV8YB673
5wKeUbZxqviD6RAAy5SDiyjkgiYqHK5JkmEoSvdcOeGX1Xm/1AtNwQLihAPMf86jG7T+Tm/uXMNv
Rl1kRdx1Kg6VLik3Fds7dz/UF0SWHvmHv+vTcjJRNURp6+PnNxMoxxfsR+g+ChRhfTMG0BSTbm69
SIyKqZPnpVnloQwn10rMKikulPlX1gbutAb+hzhjiQ/MGqLJFQvn6ZXAsZr5KltOf2d8XuPgdPv5
BFqqwIi4WTTeULi+yFJLN7uqZ9jOGV91kxlX6hZTSVPxRRDVZ44sACyI5ZlJV1HnPrn47pZszrB1
izKvx5FsUk7ioVls3VKRuumIBu4T0VJzZin4jJix9J5KcUNSydKZv7W3JFfWiconiOUCnmhwMnEu
ZtVvtjkMKrMbxIUcB4LmRX0DLzzMzcjD4C6Zijc8ACiUtnXBDy0quLbNb0b3PwR09eRZ++UTcJe1
RH5fCK3pGB2gaamqg2V+aD90h6vNE3Gz9yygYMTabRe2okbw5vXn5MqeSNRI/kd7DDaye+5e3oxg
a/EzIliYtzuAigJxrVt/A53DrDIH14VXQKNu3W75bN2nHMOfwR9u1YWk4g+xWXkK4/zhIh/fSQsU
WhvetuVTVv3BPQ4DzVYRrA8bKO706in8AkIjy/3bh9rBgrnPH2wCoMlaq0Nq2rYwuukMlYZSnrzT
V/IU1Hv8YP+HCDxdwTXg1SZeT1wEz3OJ+/VeZrAo1AjXhIGzntxtbgRy5flJX0HOLRYIfyRYnIWb
KllabSX8qzwAaf1ROW2BoGd+BoDR1FrmQW3W7YRN226ZLEjlKP8viokXcW3nchkugn4Ny0vTx8KK
E45k6dE+oiREAjfPH0Q9A0w0IkHy1JGOThe8EY6FSxyzN6DDJGk1GC6/nSovvQRSlEFdD4PN6Wx/
SiLXDpp4KZO1YIMQwYaSasVt813LA1BNvfz3dpRfDg7Uc7eeA/sM+dja1Zk1oSws6LsZlWbPABEx
XYNX4Z47ZEu5sK0oxMm1Lb7g3eWX3P2Bt6yklFXNzpjiR2QGhtIrTid/ROHVjr0oxHeYxs+g4Fhc
8HNhnKKMjkbyQYRszhoBhxn+feB5f23Y39SjwW27fZUOovXhmbCt/uOYiZjGVu3R0Q0qioXu+JNR
MneZ3LOKJYalRB04dcjIyxWNc2yJhSNoquRQiUMxL4F97onsgnl6LsBd6XapjF124+I5l7tKBYD3
x0hGS7Pjg2LsLf9e4pH05eIiPL0ww56AaNA/quafZll7sgXDYwOg15Zlm3rZQQDx2EHYl/E6aPiD
9p3Q7F6D/RK6gJ+OL7pvSiwQx+0tEd/mXwTHbCdxZr8IVaNSiFKpk+jhKzsl+LnDEbt9DS5Fdc/y
h3mh2dlF+5Mkz7J6isaen28U44Q7jFiwus7URonzKhHR/Vxdt5mXlRwJXtNQo87ugfaRetin18FB
LNqqTKPuaH4YtjXa0YOpvTlgBLgd0dANb5+PBMZClH/4rrwqQErkOR3sb0UpOO6ljNGwWAJUgORH
3Ovy1bqOtH7Sgr6h1Fv1KQft041T6TN93sarUWMEajztEeV4+LUYbvDPOYHk0sfK41m6psqQQMOh
YnI5KOmlbJn288TCu5utQeeii7UP4LhUmgu3WDVbiyfrude+VB6TJJuVKMMOFY+huLt4V4+SQEyw
sMeeHgdbNZW4JgUIN3+ARg46RotHFRaDLy63M3aAxc7aaslNHsn8EDn7W578HLetd4Tt4yHSXGPP
7UWzifm59CZgoXBqXRMzOTlnKYKh8EL/O+k6Vuqy1HrKluB5wK9DCODO6lxteo6YRXNkxLufqA0o
5FWmttdGPDqUeP3Flve4+BCfJBn0dgIOiCrgFf1Y5Bf4/rJ6s4/0Zilg0GkkBhXzJrRR2ayRetjX
xwWzi91ztjJ4UmFdZPmCjtgp1AoTnm1F7KtGdp+Ivj6PmB4VOseCf9A4W33T4kAHgLetkxpfXsf2
yvC3CibLbFGL4vPvZKoeadLR/ULnEGUF3UoJ5wVxyjZjGNuXWJFbdsghCG5EIHXmCk6d1E69A+P9
Z1b19dhEX2exTU8cAU295foxAMbGZjZWtEgl2XBVHxTn5AsFYahsiyQNljS0nQnXaP85h5WvrBcp
Qddmxe/2MFuIRKp3qjvVl0VPNf0XpAZ+HGu2y2SwPpi6iJ0/HKQEGMQMoxLQP4YAFRXCyCqEMU6i
K0RV2IjrAgSQus+XzMLpex/ElL61jt82lklc7xWXSjhXsAgZbE1tYomA1nOGxOcZ9BQu/EHcjtkE
b0O+mu5kDMpyzBpxezeu/MgVavMYLvU6jWgvIIYu4MuL8IaYaIBvLB6lyIxtc/g32P8b6nAuAWBT
xcm3K4iFYbll2+LcnkDcpf+fvlAHp5vZdn3TRw/FQi6PIR+mQZBFRrnws7YXjcx1YZDi3WSLfdK1
CkbXDKZj1fWxrupr0K7ybe3XuG/QxVPsI+K/7fOKr5ci2GUQ21WVngetVkC/H4ztKQvdFE/zLJy5
VOuPkTsrwGuVfBgCdh8vAcIbYm3oxhdIETulPQOXWUzU/nXdg06/zUbGp7KjTg3LTBUkclnXnj39
SDgK69AaphHw642yx2NFbuONA7CgFUv6C1nH4UFM9mpVIysKkvJZKddZS9VjIwABiLaTvpGX1yPx
2JL0wm1Zrc28r5qEiu5RDJqcHNLzd/u/EDHrTWpq8kNErOJvpvHsKjzt9r9KZla0Kr2PVL3uf0Br
EzLByTh8tFalGM9BPyja9cwa/7USdCszlLs0J5OAxPaKV4pqlXA3SVRkmNJiHl/ToR+LtG5YB1N4
DtsDOlZvdAVnQd/8x9QkNBp6WebPKYspgdt41nmaclIYAt/V4vzcV/2gRxxYmGZR6FgkTdacI9Z3
oJp49JzbTpcYnTGyPaMXuJV7JOhZpLBJYbkxTyPz3lTy4V0CC3+JG+bKX+a6XvksMInC3CdA2Qg2
Xuv3KEbXAH2zbcSGrm5tSQ/cP+A/00HUirhkJR8kfVlcsdC/rgoWipCPvLYAdZcuYYfcGgWQCpBy
ftWN1RGrAYCZJvoAc9RBoUFzky1DHeSNkFnnbqneA1MPmVCCpPtez9+qr/Cj7zfO/39138l/PFOV
SOWAUgCXdGLuDbNtNCYeegvpSmZqvhDheYMqezogRNmf9FKjeCHRaeMZiUnWWIdzEPw3aKMwdhzm
7aBp87c5nh8XLa5DfsplZNa99qZ5Ru2gNwmtEOGHuTeAIl2rQsvHiPIPvtFSRaREO0AqYWOFlo1r
ojrXx6zx+InJKGqltAZBicy63hXqTeiCSQE9OPq12xtEbf7U0J7wXMEWzV/ZenmnPeyM5kTHjZcG
++9ggGs5QSsk6ZwmY/QIJq8vIFUbJDdUswRlepOOnmnIiYjmY8KgGkf2PpVUSBjH6Nux/lM88bgR
RRL39JaqaBD94qRd99Rx68SFasgo0uUUpVAXmtOSLwB//3AHmf23bT4tbkC4LzOu09dHtciYSWwE
8fJ4RFC62P62GSJVM8gmfHtEcY+WRaAPoozUj6cqcpoH00alKx8A8z9gEw6OtVqzXZsUU+ocwKZe
5n7Nw54O2i1kDSTCakGDPfEhJggFdxVxoq1oXtyH60i+RC6iiurH8+gYfpMEfcxOeEsupKhd5oW7
JgQunX2ZUAqD7Sif5/GGV+CSFcrBo7MKhVIkRLGzdkIxdBBFhPGOjECPvkD5sdNeELL2tnP+OGHO
VMXTYXM0AERizaB3Wh0aZ4dQHAbb5Fy5Ha8ypRVNHiERVPTskJj7t4FIyVwvvz+NuQACsjS1L6fM
KqS0PiC8Qh8tikg8BbIlX+IZiSuKhiSRTPe4Nu3n3cwp9jwhaurCExjKKQ0N1/OgX2Fyh/Vpn0+L
mVyFhGMtPt1i++7alnofNLTfbxnd/tFfTqHIx9b2d85QYi3aprxF/Ou5b8BxxAr1zmZMMu7YneA5
j/1DepZ7/+8mhNemQDaSNoZLRgFSI8lP8FYfd/npSkrt0lLAJQK0R8E9Gwewhkqq3THacWSbHv6B
JRrzIY5RCnz61PRPb7OTB2FJW7mWczoYXctfSEvU5ycAD+9NkQT6aL2fKi7sS2PPKY+CFS6LtRpN
vgES7pHucWErT8e5NJOF8pTkMAIGu9y7peKj6eiMphRBAw3/Ru5xkrElkrx6bW6gx8VGbr8H97ig
PGPwaOxqGdHHTH01HKEEZCPrE02jzv/xdhQlVemVOHxuUG195Zjxg/IAp3vpPBAv6xBrQK3n1PD1
tLQ2DP5gB7/taCljHNerbFdraaV22HOF94uKm0ClripxZ2PV65bmhfDfiyo5buy2Geqz4hrCJM++
y5se6VlW399o9B4XFlwKHJE8jyQcEMAB2fkTRQ39oLGPJH9+o2uQ2lMdl6LRFCz8IimITD+cI2sg
QTurFvzbfIk2+dyNJ+kwBtY5GwmgVn4bLBBMvdmGzGCxa3mYcCaccwCg7FhCAUka6+ukP5AXtW8t
dXFd4s7A4NhLCHYk9Q/mHM1gPIJ8qwGxEeSrJN6wKr3OCAAZdm4RFjdfIQ5pAfCMqmjKyWOnX6Ox
r0YVv1Pllf+Qd9kVBZtGzAb6TLUq9NqqHKdfrufvEUZFTVMdvdKMVfZPBjcKyUP3P/Kz7zcqxqZR
Qqf5DjNCjjTIdq1U1m3zV5m/bvsz17PDUFH13agCWRCkCnjxKhsQDAiMTI85DXougNENSdx0QFj5
vo77jOR+/3AiVkqDQ9rmPcUDV1dVOpbPJKX0sfGnQvcXMihExfRR/ZXhVkxKT0Y3vCVlHXFrAUvj
gG5Mgp4krz5og62+1L76HIATOGaBms9pibIViKpbDKJSpjnWw87GCdht1UOtpzvsD9nuWt/Odgg3
VYj8bzyBKiE9+/ZzbZiHmTANgsV3dCRIXyshadqS/tADiwI106FQZqrruGmBqzHcyU12mJtPpiTJ
ahoIyYx5TQoeirjH+VSxK0nTJ0VcnNU5pSBoOyljfXSfJ/O85nxSsyDb2Dd55+jmSTXl/O4MKMne
ZiiyKWTkrXILW08zmCJ3wL8kuTXPwmL0t2Q6aPW8CQGY4KByj+cI6jk6Rqi1jnJXyEj10v7Z6PF0
Q+UuXes3NJxSMmeRTayPTA3OOFoatZVs7BKBtnE28NxyzXeLXA1Rp+fPDaHl4IAyJayD/C03O2dY
RUM+Fdnj+91hi315Qb6xo0+aCvHuwzSzPuFSIFiTvkoLbhQ91vXQMKWDWF3K4qbaR3is345DYupl
J7c8inc20LgI7y9VToExL8pmlzH/sGBzWbh3flR2b/YDFku0dS+ZemFtxgni5ED+rPZVpihos5Fv
jleIZuCfRsMTU1HN7WUV96+CL6b+5826MUTeTYhhvAe0ELQ0q5aF0QSxwlK6RboZrfJFFu9UWiGz
itxDfMg3DWYWXBRs+tinmpsUQP2zfFx9ALmyTPIWXmFpzRzwy7d82TwM3zIn3Wy0/9F+7jP5dMh7
HcY0jBx2mTCt2loHEM/NuEuC+teB64BfikBjxqrtvygVGkt1X1JDFNzeFvgHDRHcoST06XEDLLYE
C/HzpjiBUvg003tyALEGXG/5yA0rR0vpTNSsB1VYbQwtz+HHFwtLfyXR69UlvpzVMVoVF2Zwb1P8
+eiT/8LDgr7YNbVl3mwzxKWhGRISLCYh+9yRSNSFtVptzMurv9+jUyImgkZl0sa2EEXJCdZUs/yf
E3Fn70F75npDckVwrO1iPfFO17WDyBcdhD5RF0CgP+K9guf+y0QCNwta1+/GqZ4Sh4+7IExzcRV2
cRRiHv4izxoDy40h0/sO3N5cEEyp6CT+1M1SfzsKlfprPm/7H96CfLBZm08K0Vmp2dBcTPrFGeJE
5IG7MKg37zqdKKo1Te8sK6PgkAKP+nT17k/qy+j6ao4EswTyopaFGUfvkbZoj8srdhvNcxaKztFg
wDHSRdWtRIHZfxom8IqucIdZ3G8+lGQqitv2lZrC53psP7gj+ywSWYLd4t5dznCkVz+yifD3SQoB
Q+BcAWbXS0PIJpjzPNEuRqgA0Nm+RQLkUWKLziyRJKG2JEkvyoEbf1ZuUiH2j66RMWyMTLLNM67R
HoXNXzG8xTVgr25vba433beHN7h1+KktPDqsYoM/oDUn5mMAEoLfqsXLnhlhHTUPXP3iW93MIV9h
q3uwy0OsPy7sMhzLDBBLL59PKbpJ4j5a7HUzvzKqd8S8+f0AFKyk/Ngeerz5+UNBiIBI/+CiQgdk
4oVHJoInjtIzYTuGSKjqhXHHZ9cyYRCeAV0Bpl6PJYhsRME9I9Th7Nm0VsVe2PsMgB7nt369wkAz
sar0X+/Un9g64LRwzy/IdQOE6anyAVCoNn2x9l+lZIInHJXM9E0VREvDWFtDnDDGjVx76I5eMUk6
Rmx5B9FhaVctsqc3UPHuNBAlgW7fAl//dhpCJvsnbiVV2M4qpk4iWrUaOq7vxxhqKB5ud5cFj5pH
qa1D12sJgsuPiVSWex6cdj2MVFpmjz96hFodzCn7pxpIzQDhHquqRVSXnMibuC1iqf8L+05b/F1W
tcN5SCxBP1UZOn/FMdH5mIENInnDS/8VV3c6ZhWd/a/1B4uAMygDvW16XRDWHit+drmXZJPH4aiM
HPw0/YTn366uCbfUw7kcGePbbrX69S4hG3IWxUyzGORWjSHxMsfkQXgOfTUxIjucjq9pW8ZdBuwP
WiPUkZWerDJQXSzevis2AyWt/4grXsof7ECWL12bDI5kJj0iN/QRjM3ZejmDZkUNshr4mLJ6lkKT
C9AK43/pdwWJuhmagE6kgccnmY0ZDs5sCe59CCQ5KAoEuR9mJC0kbNCN3kp637pB6MXVG5u+LAvX
RUGZ2qHB3laiCOEgvlnulZqqQclCsnAEvrZkogriqPBoOXIJizlN27tF6MP5bu4vp++0F7bymEdh
csxh4s6yIVUALzqe9nUaAVSu18uyQZvad8JjzLY2p5Xq7BaIK7/Z4z/tUk1uI2cXlSEjwt8MQfaT
ypLGGwVX0DwaZnN7727N6T1IbpLLKZBboX4vbmgoSdsww3beluW46irwVoQmKjhhQKodUtXA4x1b
XAKLLoB4e5u+bXlpy2UYBlt1H8Dg6F6fsIO0AIJSR/XuTlKi3WT85E25wxHBCtJ73Zokltj/7FkE
TKqHArRbJIOjZGQR5a+v8GV81h6YcH2R6U4ksR2EZDl6UM9Tw9ANnt87zSK/VKIB0Um1o9+Lollk
tBAAQ3+JeyrQ9g48ySd9B64fgEPUQqTI0AjIkU/CkgVWng6BtyWS3V94GuUfA4/hJb9MdZbs+A4H
57Gejlb7ZcTJQ76pjNLtSETHqd/FQBSmhKpYXcTdh2Uop58KoGnxlPpFyRG3rYBdwN2shDdq2IEf
He3TNPlbiRZTv8Z9JsjKJ6WPZTe29SWdkx0vxvn7/liA86in5/kgceA2AzTJpqTx85U7wrE6ctYI
kZXNQXFyfjifihmP3WbG2wGjZ85H9omtxTC5/0la0kfMFqAHkJS/Aikd7pZJNgj6P4DrwzrvOMMS
95u7/6WmSU94BfE4wOwblLfzCOWxZX6VpCRTbwRdNm//jZ6XLebQ05VKIc7U3gBKcFO2RLlYrRTS
FZY+7ESx64qO5femQJexHsXYwxAhJAW+AXGc5hV6XWR7TodqDOKnMCEmaDaXaD8PV0A11rgr29oP
LnHWc0ECrJKsg3ozoi9o3O6n/dd9bq3H2OmE/PJV7lORKSQ73oq/iRDOo6OedDAfP5nyUq4yCAPl
bGSZbMHBROystOG9m6x0/1WFMLha1Q3lkSDSt/rWqZ6PAsi1le3YgzmM5iEhPooHyxLeHwOU7nL3
DLauvbHzJlcdFqohwasKtbLvCWn5HXck7iKCbnUOCwmRn/k4k8caJ0Et3sw1e/R3U/7kVxJyXrXv
z5Eje2Q3bo8b+KZGYsZz8taUrDZc46oIiGsbXVh9AHBy4/ZSu9bBjzPUrEdpIPm3KRREkcutGt3g
gBVGRjgNn350X4DV9KRyQnZHLQ/EtKE3jYkSMIRdZfCyqkildI+RDW5tRDhUdDEhl1iMoZxoP0Jm
JfJ+BmEyisAv7tATLjjX5N9432wdOL9ZnlcVcvGGKvmLiu63Q4YGqzGLHD7syGchlCCQjgAIhRcT
+QNgLnp2lDLUlvdL5FFmBsUq5TwWdRva7rIrDWAglL4RhprdMqUKFxG128Eb8+6Z1XL05Xrdkk7R
j4pHvlMuHsiltZnNqxxS/J1xZ7a7jbkUcPDpdF7/boHOXmkmSpfgEdjiWTtzz03AAgwbOp3DKinU
eVs7hQq+LdruDu4khn+O41l+TVW4dGuYsMujjiyqIHoYDaHxcALHL/MUaoGYC2CDoNyVxmH0ScFn
f0oLe0FJQGgxcZEVJHQMaeKT/bh98wKMYDNQUahIDURqiYC48PLKht1QDxqm/OMOjhrmceexTf9p
ic+mmQhX8tTL1q4FgczVsnfOolSFko96aqqgLktaigE6oMyM9y4XynF0/BNPP8vGjHhiuw0I6LZm
pMKFfMqD5c0/lYWHXdtutAq4MaRxwJ2y4VAZL7wd0Z3+QyelNX5ZRi6u4cHIDZwph/t/9jDLAx1u
G0N8aDt7u5PQJwiBY+TBKtkEacl69yCERgbCk3hCm2/d3FUhiO1/05EkcZ1+zkkNp+0SuT5DZT7c
C5a/y979G/Kwh6JoIItvvTU15L+bXfUkv3B4LjMfmLbkffUF89D4c9dn5GdXIwZvsz0pnD4FpcJ8
IwSACBwgf7qDN2YIMU2JUzr+krmBQ0y0mZJOBcsRonGhjeKeusjNqBMAyhi9bXMFyvcUemH2m57A
ggd5HyfGkSQYsAdnk0DFIPibxQ8yR3i/ntzgFewKPnnIzIsWp1QN25pYcQlyqtTUUG8IFAiobmPR
MQLArA7quW4Ga76zl1kLRbQVaui4dtR1qWIZjqTjILq0FtuQDj9lyCSjRgIaHcJsUJ/VHFyAIPn6
dM+eikSnCrfUC8S9vSnYVBTbj61OaNSQ3J2FpnjFkwt2QVUE5rorlyPJlX2vkr6owsVcjSzceDlJ
LYoDfxM+LndC+vJkT2SADDcnFoFzjyx/LQrxTzrDu9CHOevOItEj9SWFB3Q0FWu2da1pvIppqLOF
/oGDZ2TwVA9eeW+fs6Ed7KQPDQwwqA2lAu1JA1xFTJ8ggV3Ni17wjyJzXVtb69Zt/gSM3yocsY8W
yYbG2NhJ7NqTT7xp68PaPbVv6bsIxkhmr8czCHLGg8Fafw7KG8+tvPF25uW92OE2LrjYnQj5IHQ0
SQsWkmV74/fEBTrRub2BTeeOe0NPWZJvtZfRuUCTWa+udzuBovT0Hr10vFiIbpVm2Q8y5xejhuCH
Pf46FnrZFtJr+ElMn1kOldrgqxzxXnwYoVeWhMMtq5005N2Y9czZViQJu/wXUzXxw7FsG9dqgNCU
7l2EroPWgtNC2j1JcSbXxN6/G0Cp67fxWhxa76S4NqgqaSwlPX0oUQr847yWwY1/R0bv0psPeD2g
n96W5MQ7XYKdSQOtJ/1E+bW+bDq2rOt6wKYwJzdOPoaqeMLVeMVhZ9a85yFnVQj/sQSID7ncdYY9
iM8EfBPSV+BR2UsgnbG8+EwexEemciVj8oYQhFqQKKk2gLh7d0io3pNUFo4rgRMVx5fFLeAIjCtY
rriGzJoUMxmL6s2kehRmiHG+H+UKxHpJrWuHU25JNEz6/4g5hTy6VTwcrmNHvqu0YaeLfr7Ha3an
IFgcJNXwG6UHTcQVzS+CNmvfVciNxqBovDmx7GAiUQkPNjBQmSHACcS9tdqL7/nz6xYAEGICre1S
cgAxS8Ggenb5L9DiiP46b2zqCmQsVi73ZNDQAxbtBdPfSzN4nD8syK6qKE43wqhLS412mQVmfBsP
+IrMYkpN+SholSghiFOfEeDS353KwlgPvlVeYVsh1bGHsu25wKekd5LzU3S9cJrwDdMPPHRyoDNX
RW+tvmPEYKGFJEmrEqWYV49CE/nUdtjtSe8noY+4RlctTvDgB2lgolFvVAIq1WwnGQT8BQe3Ymil
tnzSfrljY8sXThDQ3GweLPl8A7Kh00m3Uk0xt2FTZ4B2O91kEutFq+Vry1QS+AKieTylQb9d+BpJ
VeXxt7cldP5ADQ3VCoIqKtD8Sr88rV5hjp+VtJFzIfOPT/rdfFNU3nLWrJmgrbeIN/mUmdGdLMhx
DGckRDnmXCU4YvM7YC2Qv0eZo9zRIHfsxK/NfmUfnWV2ZpqLK/e+hQ0/9v+Cd+cHSHB57gsOMshi
6fzboZwLdUdRW+7L10gVOp5vOAdlC7N7UDtctfMjOwEpHNy26pGaih+qlc0hixmOi7igYyHVCgzi
ZN1aVnrbDQNp6z34YOuvOgcqWJwwaNQa53eJ+XeGHDZCODeob7UGLdsjCW98V7AfmyD/5bjZoOoJ
LTry/Ffns/UqeKZUoAuHs9Fcmhe43lJ5sqU02n3TN6jnfb89qeW8jSwslqBDoi/cIER6l+LLTNQ1
SUnsGDx+HL0ioAKXsjqBIsuWg41eS4ifekFP2D1+KdxBrMM5TSzrHdMWzjHDzhHknwEglzQ4uYNr
xgqEfet90WDtbjRusHR3Egm6F9X2cHEUjdnAbybMyajeR9boUcUTiRtnTR3DgeSfSP1yx0OUXuMV
55KtcUq23urgYfxKnCOtxwPXTQCOrSEGLrCn485K+9MmKl+Wm6Bq6bkKIO4cIOUh3ZXUxOwq+dGP
+7Q7Tkp2MPOd5VV+L1f0AwGbbUNKsT+hUe7qdjI9Ksls54LiTL4R3rWsuJj9QEbI83L2MI2DpcMh
l3cT65Vx6++wi9mx+9X1FtdO186S0/v/RG7/WYKHaP1hra6WNhM1Rfzw7WP8g4gjrGSO2XDJG4Px
vmOkP4nUsc0jCHR1ZAifnuSMEoFxHcyvTWBaZB/0ILV7EtEACbmSpiYIwTqz1ZihSN01Azd3T1Q8
yR82/XsK95SdHAWesWJqqdLKQNiScvOG1F13Vv/bLZvlUg16vpOu5yAQUnheLh1xe+n62wq5jB8s
wvzCY4eI3EG5K1gQQ9S8oYrKBfwmL5sa+HyAM44mlM+Q+rUL05RUZLTo1ouoSMvokyrPQk4+8Qkc
sietsmStXsY3xfrEzb/09dlkFIQj2Su0UMS6Noi2ulmHzaG1Iml7rAxWqKhAX2MEZQssxfgTF99k
coDxzBYzQ1zvAx8ud70YkQ78npj7kCefxLNQ6OtfwZVTc0nDqg0Mbh0j4lZAOS6cZeIMrkCKRS7F
+XH4QV9zs6oA8BwTTohPWAYBfNFfloJhWz7Gv5Za5COtDk8IyW3KSJCOcxwlVoOf0ffbN5lnpSUm
SuCtdh5jsXKvMZS41UdCLmAVj1Tirvyh+hBkXVclr41FLfgvETRz38aT3mifV2EzqRxbNLd5qnXC
wHDu/QInt7HaSo0mqzcD8o81C77kEyLYOI8cC810ORy24hef9opCn6YogUO/4H/sRuZsgoYUnxgR
jgtpP/RJyA35g00Gv7uChyXEvABD20r4p7QJLy70fq4yhgx1wcIeyxdqS/uvpzu9QfBK1AEnzpit
Zx+MrTcLk672ss9iv0DCcn835UfUCZ8e1PUbkdVjMsqf//KuKVeuowcQxAZqW/6KHcffzr2w0YyI
hrlLK9N8e8MYxOnp59Ox2bRG6UkJHqsWoOgJAZZ5NfBa5h3WAXV9iXKGsM2lce8Ba8xYaHXl5bVi
x4Fax2M2NuWBDN582SFCN1Mvlkn8w98wr5vhjeqfr9RLjnXFpKrYIgXgljICiCr2bNOJXwOpML7Z
TYjkkrhbU2+CLbtyZ363z3P4L27oJe420hhr60+iR3crkqCnfuJL7qNgTNhWio3q3eM9QxfyH6SH
YPAl6YqMaKIs9Isteu3cuB+XmVkCSTKR3fV+CJ3helDgbi+/x/JfaDFlHn4PRlyJURHpuXftKoDI
TJhjsOxhyfgeuZ+e+3g9XgOgPah/im07xQ5DFYIMAaSNX6qcxyM5D+7AcOExT4h3AwEoNJWPs5/z
XeF9+pzvrw+Uw2m5ZKb3lWzaPuMvUwhmmA8S7bxHSp5/k2WxtqNIDiDEs/uCE7+I01clOJx93RWY
tl6fFYlVZI/JNHHBRg7Rr/+VQ4tc+dyZNI0L8cWBirrCgwp0/mkCuFavlWkYZFMKDOTvKnGGEh4Y
tqK2WqAw8zgX4Fz4s6FxUtXMzqj7L7SeJ8JDia3Iutgbs+sgSwTEjGs38HuaJpEPgWuQxiMwWXPb
dxFiJblR4sZ7W4RssVz+eJUOrHSRoZeZgFWL99A6ppiQGbkvPmBwpcg4jkjyd34BksBxm/pQwQB5
l1KfipIJaXsHPi18wg/Q0DPPvNkY2CHb917f9Az36jE+wqPVz9w9TO+zfR/UDZeTT5Hnllm0h93X
nKRPnf89F9uu4RTk8FS6H9ZwTyz6ohL4Y2LHO2TT4iM7ZP45GRhKDijY54RMm1iPW3JgAFLECwRS
nA/hhfCBE+fT/F/zTwcLiuriFogG9NiACntpb8TO4E7ei34iXvJKwMwYteK3CUCw9SP4OFzn/NVS
0RfOoBT8V43V2jsOaMV/Kcj961Do8fSISUJmD1Eq8/ULhdNil7OmloqNmebZxT/7EgTgM0KXAf7c
545qRlVknHpHSWZxlbL6T1WxhZHgPDNbACCzeXG4+v/H4XpvVnyPgPGLamgE7N0C9s/rdykpYl8j
I3p6rrMTAbv/wQ6QogyhSx2XyRgYZpmrSnDk5CsHTWjgKo1tFVJTUwdu1lOOWjW9Co73iIyQdnzk
5mVkI4w59N6gsA8dPssM/PQngrr7hh48I2nEW9oSXV6gGbi5kHWytWd4g3D02QjLza8SwooWJwhK
x1O/iCpwTyiCAZfUYl9zejY/DLgfm9HpIHWWRPQJRF0j0RDW9Fy2i5ndvlp9lnVEK3n+k4I4sR+p
60q4xCEXknM7vBn8+whJdmCTtXdNMthBPTkZhMCV0wnSSY6mFyH3cmZZMm/vcR3IvHrD7EndTUub
k5oRs9CzqcHuzdefIdAB9nFrLao6MRjSK0dIf9r7XOZdGSfeQccQS+iil3by0d943K2kCj/11Ckb
4Q6BHvBdGk5OLodTM9Wd+/va8K542RIFt2DO8HpELgqkGSPt3KkxARnJ6wGP5wRBajaj5JpWU8Ta
MrXB6RNVbisoSH9HYp1RUYyDcZFzIRUOK6aGqCcgMCKEYGbjnN2HlJBXO21MRA2BcLUAGa0LwF8U
SfEH9j+mDPgteiaIe0AMU5WxYYiiqQ1Kigu55RkmGPbsPUGcdrdTKb2xUEZUGDfyYG/cEKA5JaX9
cwikgN+pmWNfnMkjOcPkxWq7hE5GRkoVkN+5z+k46pKvWa6OosdjI4o+k2mx6r0WXIa/FX+lDI+a
M12Ef+e4rH/I3IWaAoHiYWTEBchJXf5nSCrRMVWjcUSNB7ictWJOVu6qtC4yn5E5vFwg6TEPQNSY
JzeBAAuH7Yu25INaIMJSXT5wsLWfCEFPN+8ampOqYnUs1VOhvtzUCIKPEe9/McPL87ffOfthshBI
o3qaWHK+QiCGgBPR59q/Lf7V9UmQKh3x3wyZsGhtNbvkVyha9hb4b0yNBPyPNUgskY1hRgcQzIRc
hjVAq9j4ZXozYWD2Lyiim/S20pqNQ6yGMD/wwCVXiwvkE8Ucp6l2Vy+LNbrQiBzGS3LNK8GcQ57Q
wz2QYlCWK1RESq9I18vB1YthKt/m2Y5gqEABafB1/PaEMyApazQHUV0ZcGwpj+NPDJI39Cob7lXg
m3rnbjV3fg+jEUOwRlOm25ShfviqTrm7Vi0u0cbsZlvK+DbI/May9U/wxt/sQfax9tYfUESpuUpV
vQBLT/c/nuhW9KuYXss+Z+OD2ipkxOtFBtY2yq35pDNo4l7Fu8jKvYhQGEtTA+5PkNx4eIXXXBnc
A3guTGdiXOBw1Tdlr38QVWWfAIIUxgb60FHUm4SWAoWkrX2EwEkaFDO5tzvbo/KSuYkGgHiHjqur
y7U5lEiht58iQAZkRiwMCXIVQsSAg2xM77uwPs4BYVmoYQBkdWLohD2lU7XnshzundIgz/J8aJDO
vWs07QLLvvYRhkOFztetDDEwQiKdomOOPDzLyb0NR+Ij4ESE7+ZP4ieItT2d8oigCENxLdzkN5nx
yDo0Kn7vOJhgD5uO8k7+1V9W1lbfn2NLJgCx8pytb+x0dnZBlaZGu4HtxE3yqwZumlmAQE5C9MAH
Sd3G7OMHkjVHvYhaKFZf+vTFWh/JveP1unozfPyY8I9+baSCNf6XcRiSTkknkLw/Jr1wxVq16ffr
rhId/PJIy6th8O47DD+81YinfE279DiSVf3yGtrT5eyYrWfbWJAjK0OXTv2uLgUxAnMzDHKnqvbo
ai3448d0anXs7czQYWeXHkq//B8nWVr9TA9ZPenOIlb8vfqO5cYtfZSi68kh+QBWqgImpz4P2yX0
TDfTOj+AAC4k+b6JmZhsGCcOd/AycNRZhf0+GIVsYD7Tbzg/CZdScCYgXn2h16reT1eBhzSQqKzw
qtJRQnvsyCs7gcxGo8xGFJNMgCE4yova4/Bj+Xfirdb83mqIgw87SySGOIn0llDx+i0+72AJyLk8
zclMYhRQ5/4XyBzchvoe+iWM7jTXj4oXsBLqKv9Z1OBtlcB1iMPk0PT5RnV59dmdUarx6j/E1w5v
JIgCC/GN4B50DdBQ64D1rQdky9plI/mCVC8sKdpEa+Ug8a5b7gXMT/E77VnUZOzkvBfPIo/MtiTy
DqcWrZyX5JrnFuhTCQzmV0F/agqur5h+xF9spx/9swAYVBl9H3GCM9HX2lNGMXTRwCxykJOes8H3
5o5BhqBHRiwnc2QcWvC1E0pPFUIbKRdtEtp1wvPKkkBW8rsWjcAwOJjGJ6OeFKfasJeaGUtMTCig
9vVeSWASpiFxJ8aYfFVkefv5oyYgUIOMhhPkaFRbfajGL8kLLUmW26yZIBsifXaXpc/Wgmc+3+i6
fsYfH05UF7D112rkiQhJ+83j3r53yOWKZRdcq8A3sqMIxFULL7NsziLpuggyC1/jWZXcqox+rkIF
oUDPIumxT1VM7mhcz8riVTyoWaIiZx8g213zDvZWntoF81mnIXtIFroD5SR8QIGUJcpfZJ2F0YWW
VKIWX9ni9R0PRiT+h/uMbf9oauxTMRCAO1+NuCfkhPx6YuGL+5vZGR1DbcK9JJNqJiLO3YGbHdtE
kuL9sqoUEs6OTcGupYemYbffwE119ixvV/jJRi+1k7ejvTsKmgA+qJUmY3/YrQgZPEpMNIL6gpsT
ZLePhOb6h+mTNR+YXCOVwPzFZV1L7uRRMRkYnkvtHVdmt1jCw43axzMk/E23N9g+l3JxsKiu/CkR
WrSz90I1cGbx4QDaMRU6AU6oSky5qw/cFzRPj+wAHxzNQ4juaZ7Tg543LV3wduPCbQL+DVw3Pn7N
vEoQFlXBCw2tZeNOHT19WKCtyM2RBd668pdn/B8mqOz3qXMJcCiInQ+uWGyomBtrXCEwLmi6VJuB
aZ9jp8FT5hF3o53ZIncfto+dlstminv52YxPL/J1Ix7HXlPHce5ES89tE74FpN17hN33KzgexodW
0H9BnFeJtEKueUIa74aUZQJYFYqRxNjukizVbBhimfqcmVKZb9ocNfkZu9R2qGwF/W04KgBYyFoz
1Ty8AeXikGUVYrUkqnNLCl1TkdmlgvPaWNP6tbwoJaRg09jDHb3VzGtbpC2+B14zDKiFY5Hm2HVr
k1eFPyXESvwch/lswEYxNu60Ips/B5wOPAlBNOEwDeo27Ctgbl6F965iMgfAmfdvbD0lDv9i6pLW
Q/1i38iM5A8unIFQrr2Y8aV201na8JapNj9tSkis3FBeIJ/mIJqYMSiL0Zqzbhcq4BGJF2XHQ/6b
5rKwwkTDk+V2vYYUV0T3VKYAeMy+TA90QM8KXS5XaEkvzeGXtss/b5Mdfh/sdcH3MQrB7uPm8QHE
7t+e10aA4xFMahLBRSeXgkQPJU+5HVAhPMIv6gKU2tREcVLZ7lB7TxR92Z6eBYIQgXsuBYKu6Yo7
1HnGqyhJ5HsMpkz9jI8aEgJceVk4BWSyJUxjL05Hq2UGAyYcaGlfji4P6er31oWAvEnebodkPC9s
MvY1mPwWlcYrB3sYLxDBSmy8AleMKsPWHGPe9JQOr5TYAqD3mhV4/bM+I7/QYWr5J4DsdtImMOoH
XDfkN9z5lgR8/BlwyN6My59XjkDxAYekQOCDfPq/5d++1bUp5fNO0ZOZiJ4tzHb3C6hNLhHmlg+o
wILwqcnF5MDgcwJ3ba9Y/UX0Df0BboolN5gfg31RftyU6wR41e3DVxLFeeAzFVTFo1g5Q8uEm13x
2GznpectzyIsvdbRx8pXMHGHRTDPLP7dibDUgP1JvE+4AU7+cb3Z7e9qxfp/n8T1w2z8WkAKNdkB
isBidcUDsm1coBtIogYiQVa3XBfMjNdlPtzrbJ60py3Ec2j7BdoKZfqbRojj7DIzjhY7p53v2I+p
XdfEesWlKyN0HRALqMNg+hmfWsqdPI1QVKvgTwK+tH2U3suXMEJxyAUQC0gq1lh4uxjb3i9GPPlA
cGxxMGLAT6ZEFWxsvxRAQ4RdUfJe5/ULBEvZL0Vxm30NpsA8RrE3jK5m+0KY8RSYcmzAsPjqk7eY
fWvZRPzjucRBUEGJ3xiOBp2qDbYHj97CwwYtUTvdIIruy/n0UWxvTPe6sy/f4fh9EGCeT3k+lhPX
Y1fODRp8n6eoGzXsREv2kBE9qw5KA4aZ8yDvAIXNM0gsT0WM1ByHwfTfDazbEejthrBq9YW3Rfua
34k8uhb8T0Ze1CKoCdld2nUXwvQvTBFMmjQ+rxpXyjNvUZ09sqKwQE86CMU8fZ7/+D/W/XxklJ8N
v93JUOMyROfoTHVMiprgN3Bdl8QQeTRBUImoxkfQCJm0s02GcNKGSTj6jg2GKeLzR2DRgY6eWPMW
uUuUqp7XZikrv3gszrmNI4MInWaNFiZ91PP4PF0+fMh91lmEW3atZ3/WxuIZeVpuQAuK4UlaGvSf
FI6eKbEZHnAFg8PZSYKo39PJPT+Wc3+YH0oPCjYFUOs/9FH49TuoJkOFZ/WwBrDHu0MQyGGxxz9J
cloyWrpfiflcr7xTq8IdAe78d1yz6gkWpKNbq4CWCBaQAvy7n9YeDeoQHTWX+wlM2r23NIYiBlXf
vq1vzzZPiPUjB4oF4Buj4VNoVs1IOHBH+jBLZjA18wxxnBctsc6RRbD/Evx3eXJQw+pDP23MuL1L
kV2lwtoR4Zy1pxSh5pJe1XmnzITsGkqPvEk7+QN5CyTdJK/RB45rq4lJFq2fCC7lGagkhY712jxB
G97H2xUjghsDzq0f0i8RpQXB4VbVgcRc5bsBNX+0tBzl1jVWbdOi8YWZlYdiOIU/ybeT1QTyqd96
zltCvFT0Q+crsBuWcZsFK/4Xmo/bhBkXmgzgFOERRgGXQQaugrU5R2H3erZbxZQkllZ8LBSusgRd
IcIJTzyFr9MoxRTXF3GJoELoNmfD7TonnUttEnzhzNbVSO+mic/nz6MrnimQnpTy8vciXX4oKQyx
AbUHjdlGm4staCjXYgwUif7cq49ae9A7h0/1K3nWrcH1Dygyd0E8eflISkPk1tZvASuSQMLlQDR6
av8ZJ2/upLAnd823k29ARiiC/RQgMBl8kwQiiWkVCB8hJABK3ArmrsZsrYgCV+45D1ZYkB8Hij0M
VLqgfz+SuuewBh6hv79DiQPaKrx7xbOoybrrzUb0FpQIHkJdMd07fpf2MtOQcOOyNZQMMjMApvvP
m1YvNa9Yd5SJM9FpInP4d02kw37e/POWhEPkgCa2eGY7/WEK2t+N+LmSAuKiyKQnlc00qjlgI1rY
pme6+KYokAm2OOERuUOEGfB5EaAWVInkAVCzW2gnJEPKXRDJug1dY6nmw0DNPspVU8wT1wzOp0C/
ncAxMlpUQio5IrYBdbRaRwdgUOTfabl4ax7irg1iEEP4nuvpRF973xdAP3j7Ynw6PnmYaR3bfkFT
6PayMtLSBxYnmKwECUxlRs+xFOy9IEWPzeHMqMDDkU9orBTptpnKMzV1JZW6tfw8+cq4eAx9KSSK
mJ0pRm7JR0SaOCWuMTPvOZoDKtAkvrCbDes9SWejiZD/++v+l7CPY6RFscbu/WOg1ILfedPf25VL
BskzNY8SgmGFF8skzq7L2T2t+SI4g7/SnWXbcceLQI8/flCNoWN79J4JPhOiy92nPyFP2ElC+J0S
+mFuIh6Q9ldo/HF3gqozVGTKAy3X0Q0MF90eV1x6rrdaT3srUNcy19aJ9kKEEpyG53iUvEK/cK9s
0suaGAQ8gSxQT6N8IiMY8L4QMocfErOausyIm3tWSK5Lkq0/Tzt3YLFlsOuftbmpWClUyYH2ePjB
4p31BUs8+DyssVejLEYnWB9/C6tnRQYIls4jQsAHJXv+dYRwKQr/84GraCgEkKt+cy3HBc3NW6YW
d6rP61E5XYzchT3eWC880hZKz+02LNaCX2eemFA4O1i2z5TkyBN/ZsUsdmiMTxtwjW7VbhIKGtt0
ooGA4J2C4m4BLLL2qVsyBFpxUBNsp5aeih4J6UKcSRzfQrw2LQ8M8cG1vpif3og8NArGpSia51Ba
Qo7O3OaNeDLsixqVRp6X7KTOQF73Wqer4idyxLOHumqQtXPZ4MmoeZgvKiCX9wUXhkRG2E5yhsBa
ZaNZR4FX+E3Eoa2xthjdUPVBAwN4pJJXCywBit7pCt/AMiUQWNaR31ixzSc/B0C0H6NBXCznRpD0
xra5aLN9t40VYA+5Su+gK7aDHSSjY88xKDLxt2JDcsAIcCMHIoBCq0SOOmNDTtAz9djC4ReAeQbt
uLI6rft1iC7R9MS4BAXuGzSJ2mcO/ZVGbwR+aUrSi+ZVmRbV67WiQ1Mg8a9fMxei9sdoiBcqkvKO
oAbxZTZd5tpS29qhN+9VAROKb6L6RazB+TAHPM/2lOse6BDiebpKbQf9ZLqHCeMiCH7epPMmL5ui
JSVXCZyXZ2+4sC7kweSfJ0epwgwBEZOg7OdAUqID6LvYWOu054kH5/a5COCqE2ShfPmkd0Gj+ljb
oapLRwKWyyNaYZirQWRGlXPgw4HA/NafFeDPHd1ZW74hVTSljBFMr1zxL7CcIFyuIVKzdSZXh6if
CXpgUWyg/3vNadg5U7bhhrlchsr0ISZqE2MMuLEtGBeynxduBKHZOj1frAMx1zXc41+jyDpmiDlh
4wD4jDprlVCwbCBgQDukQSEwObXzvJ77rzrKHH/hoYriQfP+2vcvu2ji1hwY+/6kq97cpH/N/aVP
UE3xAvvBizHS3+UD1hQF4oHRVWq5R7BLIWSAcDkHPgmrotUk9KbazgWapZOo1j5XlMApRiSgrsik
3IgfkLkK0OwpnuNBbqGBsCpDXNPdG3RWwpS2agBd4L4rkdTrVZQ2hjsPnq6hzACDWJZdKIyp8wsS
3e3joYKMWBVuArxAMCS3RJ1QqVnpJenA95KA1cVZoMOL94cqAtRrN5wPp40nGoBlVoznEdRPygrp
AV7O7NLDFHHP1lOTcib557pdrSOYvBSA4354dPlGBkF3lF8LxhMvs8hmpiyqxh8jWHs3yAzRfo7b
1HwXxkJLOzuvq6hYhMfN4AsXtxaQIkHSV2yQxy8+D2WxicTA3A6X7EGCMoY+GzehTah4Q/CB1myt
MG02mnHl0wun6ErRNsBElC/3Gl3DQsZqRzIR1HurS3s9IxNWF8paWjEhOHrNVaVXBPZVPHKEg8/B
jtz+jhGisSJh0UUD0QOipYV7Z4aYT5ey632K3UvFnx+wuN8I1oCjObOTRzgwR+mb1s/EjzVHmkw8
QGAV/qaCp6oxfQZI+SXCCMmr8lR3rybVLIanQSeCfYuvkdVoSVSEqrAJ16QlLUhpB8gvKyi7oRKF
VNOjnfjv4eeJ12dr4WLNrMSN+zoVOoe5m1P1r96cIStXZbFNPBGoCHtW7lgxEvqE+LBjk072O6gO
+3JAAuUmPKHpoGfLIA9ZWnRjCVXgUv8K4AIFXqQ4I2jm0c+zyoaY30+iZaIE+Mo4iaxE27PpwN9X
6KLXVM1UvmBRR2I750IgAXxoyI/mNNyLQId4XyHCz725UesGJ2sRWCtpQ+UFp5x5JkbQ0JtXucOw
SZnAkNvKHujdu5+T5vs/AnI+I6gexWUNnFNDCvAThRvtT1I+mSf7qFmUzRMKRke/V6PJHa3SH1a8
emcyHFUE5/gPo57Ew0dSOz2QNsQMG3m/VR16J4PB2qnDQJwT0cJjoh6bPZdoqW676yw9o5V8rxWL
ujm0PTOxKJmRAqLKuHfSga4luSO6qC3DqR+YNIsX3O4XWlcIDpaEpl18n7h4BzF/28wS967yWJBj
5oyiOtCnpoJerCrCIus9Etx/3zbh2OB8TYkbsqkcdvjeKTWxYUyI/3HRA+iKME3dETVKO7iIpB1k
Rdyamb697vR6btH3yyf71ISeilEYYb7+Ma03Nzm+KWTJu7n5hUrR00M7wkHzeglpZfV1cwGzrUdt
Olcgc7v3hdVkeb/YqwGOwGc2DHcYCQkUnwZatJwfIE/+f+YlTjxw1RjTls8CuovdJ4tGusfsQZ+9
TWQO9EV7TkZn59+90qPT1fmZYnThp7zB/pY58O9naZrz8V/8h4V4aqVd4+35/BgDfKGMQ0fkVqb8
RVA0aKsAJ56P8owfDcqe9eAnNCPm0VgPGzspvn3wkKT2g0R5LYHskzcxrUufw90seYWSPU1Zkd4g
dRnV/mfMuG2kSeK3iJWZMHcnhzFAtUXUHlURZyDBCy3sEANetdzbA0RVxWBlh2lzZzxqdv1efIp9
Xy/VVB+X9qCTSzvDTSa7NpnP7+7RrnRt2M9rOsOIUx4BOWixuz3/qYzfIkduJByJ854FhP0THkHS
oOUrCwH4WBwzHJbMqoWu+Hs/jCR8ACTG7SCwduLqCN6/QzRer8fEs2JbpYSbPupPzipgLcCgLViv
uiBuqqHZZVxsEpvbQHV37GmsDtT5Op3uC13YJTSRZRXdgWFhTFIxyeV0doxlOUgqIlLao4G4HAO/
2zjkbdJDlQq2Mr+6NF5NpYNIRN9swI/UQ89GYReQTY2qrEyscBW1wjFUiDUWWQ0iILhzHY83RnoF
PL3ZSCcShCAVK2e9ngKX96fT8KBTnfHcGBieiyPetRztDrWj0fYZsYJm5nEuDuNRuQ4KXB8bw0rm
jG1Ju3h4fCnfXQu+LZU9re/FhY5VzdoWnP132F4Ia7DXph4lTC7XGo+sIXpQGVCIIrL/NgPvNi9w
vN0Zx81fdT/X9/3Asn+YAU9AybGz98mmZM4sH9Dejrrk7VAbvyHGAdbvJ4vbkR7JDC9xoLQLhQ3v
ljIaij4zCIcSkBksDZYx5z3dBWoryqRZbRm9ZB+Gb+/hP77KddEUGzWxR0nxC6PjjzrdMCVzNVcb
XPvmMniYdrcHN/daiNipPje8do5gwphLfTVJVPuS8ywKMDLdAD0aK8h5aeMAh65FQu6U05Ito7C6
bLhCuxPseeQXxSGfYSHJtiWv+4X3CWd7hN5sKdP9hu76YEqi4aqS3MOfQQMTMO005VIU1cf/gTKT
yhtcnLRZIcj09xcFWj76jmLszEYvEknyD1AymMayNTeEh+tQgDibCh+jWmfGBecoz1Gufdo8nDC0
3XgPVksTiZph0N7fe3D5ftYkf1T14Zb7l9mVjreqnTA+wcOFCb+NFa1uZ30HAqhuCY57DU7M9tnf
/M2p4U0GkdVc0eUCzOG/j3JO6dlJThbSJoDCJ0EqR4ItKVGvqm9e6ZhUvfNF61HtJ0cuEs3Vm3UP
A1IBYxEB2ozECzVqgcKCa85CdnYEj4n7wCsW8OZfaj9ofhkTirdTwGzSKWrArpO6qgsGMgnGz9ak
b2Q78SbnV4ENjLCw2Rrei424UwExlwVAJVLeG8EeFectHW0PCJxUqf3ps+mGpd/lkq8wYoJqHPHd
OuEEKo7DvQQpFmFSTgKzSenEvH8v9892VFiuYDy3MNdifkMm34ceqIK8m/qR2c737e1zxD6gNETi
CB80sy357q2ELYkf1RD6196y776dp4zPRDA0PkodSY1GKeva0iljsmbq/D6Qlk4rxJmDaSMwnGDC
1etsLInuSIFR24gKuDbt1fCbKSZtV7mmUvSmmnzFuD9VYP/yDt96rjDErWkZdLmcVUBpCNoWDRjX
fQWI8uQ0n4hFVOxPaFtxDeMcC8ma1WqZ8AOF6Mipwrz2a+ePip8QhESHgmRYv//q1XTXy8YrRxZr
n5FHdU6fgWYH5tYQ+7kRZeP/Y+ucFx77QIOI+TUFE2y1op5XKTXtLJCWdVGarbCs0GYPpti2uNO3
zn1xRHw5yXTSQF2LJOFxB2dw8dB2wLwEueLpNzT4X4hqNWqG3eJNAndwSUqibtVEiTEZd5BoYdHU
0ukBCWs9dZfLOLsuFyRkYiaypLmU9YwSPjJqte44bLZLWmnSoEPpKHjNd+6G2NfYIqDmJoftjyAs
fYe5LBop1ue3k3iaUk32UH2dJXnQexHWRrUhCW/5YSRz7TV+jdgIh0HJl3f6WexKV/J4hRnfSlkh
dp/AascUW3H2Xz9pfQ8rBB7yfWrHF1ZRR7CyJB3hOY7A0IYjUyTDitoq29oSdrDZrH1924+LCGkl
+ovvE1roiOEeIkRIo8ahhKOlqqPaNNTh/5jl05vh5j0E/2JOSE1emLXtExxhyWxbelanc/TpNXwK
0GUVD/nUenfD4P5erOIHUkeLSmwglfqdJbnWYol+V1zmAa4kNP+tIL4Ao9SguLVq+9YpTCapSSUs
kmm0ZXUZeDeiyjAVIS2cSItH31w2ryOgQZcNOvlQAme0TphFBmsroa2SMklRSOBXS6Z+izsTrMiW
CeGNbfRaws3YKy22iTSp+rqjeY6blZP3XgvYkc/lB5Nl6Vnjp0TeVDWvb3+eQXyvsDT9r8SmZvDx
1a+IGM0lRQ2RjutZOcgatreifLwfAMf6vTyhnMjRKhQ89EQ/v5yBjDdvDZEQUeOQFW2RbqzzjIAi
YNLdZl/bVNMzPgUfGuyGJQcVmKY1Et13REtpY9tolVLLN5Ko+a1SA9SK0ZsCZYfYzNKTYHG/7hmh
kqJJDTEwR6WgMHv8TTlXtU8nESNM3fnWqsjr+QemyMU/6l1uEGNQPjHiUOfYAb2jaQrj4p+LYxvS
Iyr106xL2jOSq0lxXuYZ6JjboW49Ctz06eGyQqD0u4AaGeYaXNtbQZyrEt7V2HgKb6j+WsVLGw4w
cvGum0kihrKYpklx+n6eXher0v8F+CTjs8oCKpRNAoc400iTaDRcDx4BeKWqPCYvmvMWU1Ek1LoO
vH7WtnEnRtaF9BMsm38Awn3KNvig8/vrwzgcz/9WjGZXORhzN1x//IAz+oJe+8fsTyhYz31RE6P7
EigSt7SSTz3IvogB2FWInT8JIY5BwKnDtcLwjafty2nGiONETheY28vD776/wARN/5PNHvfLXwvD
NE0iFkMA9+DkO0F4qHRqCsYjXgPqyXIHxthqzehFlDmQFX+GKEc8corLHJqXnRzK3sWhaA/6qu/R
szT1IL9xq0HdlJ6dbdkVEeorv/VZ5NYd5a9f3wbNd6gTdLrZLVpQnqLts51mPce0kPRpuHgaGG/N
Zm2TCJuGfZMFhtz/e2RMC7eb9AccpYp7DL5vbUZ0pH02dwJ9+qlFQwabTgTCddjnI+z75Fjj7WoX
aXgAwXe107FOFwoS4keucREdkHHTA9izp/H2UK0HU7EqeGa6Dlw9UfemZg32Hyf70OYRtBeugEkt
14PsSFhzigVP61VmReLmP+znOYOzKRc+QVQhSzdek8xawQQWCEy/sxYxMrgqWvdA9hLgl8DQJAJT
5OCEpYWK7b7cfqaMW6kT66SVwBQ9Q5wDhDumSo15hyohwkO4e/V15IHuTrVgceiHGRG7NAa0UOms
i6FWE1RsC0SDgEbL7x6RYAAVEZjxiXuoSZzfnGdLEVxps4DybCw6/wCAKiaPTZRWLxwMCHtWLDRf
T6j1YObKVOWI6LdT5C5K8vZfSFerzBwdziSrhIPDNad46bHLGONSYKcbtavY9ecA9pHF0QjCTIJw
/v4LmHLOnVXdyvTOqHo/XACOOiap3wy8QO/YxNRdEIJblr3DyTX0kdhfrRRSujjjsnHdE5Wpu/Gs
OUiEqgkm3Kg4aLofYTHXFUZuJRYvFDAFMz+B0Rqlx09DdrYuUjaAjFJSBUl3/eoD+1Nwz/VbTlQB
6sDml/bLwLMvmDR6/HSrd9dLTZ9Tj40dVkeU05Ay8UWOMePyaPDxEHJdBHsUoa7tQnOy31kB06qd
2z9nZKmU5QUHy7uXIG8q7zTvMK8CeBDnHwIXrC9k7OT0eTM+7JZPbfNbIcMehHb1ZSkX6WhkLph1
vZs+s1wrre6jyRjg1UJ7x1SOUiWi/AqZt4+8/jk6ppPzQ+1+z5M4D8xQPb4I6OtItlH6UC7WSvwi
6yITde/P0DCaV1HKRV/WVIN8kNIYHF9rTp1gDDqp5uK0vna9Qfl8PfaMdH8Ry2v/zKp75bCbrxdQ
YOVj6yA14jeOimO3DzDd2yVHKtKQ0GdA5Ag7Tm71iNkBOuQ4iSEq64XwoZil8bs8dfYOz6DZn48a
gqf86UDs8+czL/Y8GWHb5TWLMA/Xgln9aKPz4aP5ZQnN3D8uvp/I60TEsIersqzcNPmtkU+JkaZr
22rWvAmVkHM6d+Ku7qItZ3l/iLC6HBSHj+SRpI4nSCAHP7zlB4uS3SEkek5BAZFhbfjcWzzis0x+
MB8FRmjTCxoUeiXAfmAQWYhooJ7kgT97jhUXfLlQnSpw0GDbWWVBIQ8LV6Y1VEzEW6gI5qIyOzoj
6qThWvq3RtuUryaj4Vg9bt87mpHogLLFnuXIIgwdD8Sr5sO+u4LwyeFveC9U3SXcq8MDA1ZAM+cM
MjnjRda/eyCayrMhiK8TSceQsbeOybPe62AUFyQ2ZW8whY9WOzLsiwcL0legP4QqZeOc4UD48CeK
FE3V4vVZvSrHQGQJfwv61CYc6egRWVoB8bWPm0O9qVvg0dx+Rvdu/JZGNLBzkpMxAH5znjDDqNJ5
Bu2xoQlCeZ9pBC5RRPozLWcgsiHJzLokD6cq9CV+JJWoCUIUifiiv+/64L9dg1IxFGcBhoEFOLcB
qDqMG+XzDzDAdxDKVGS/0gIAs1Yzr9Pns84OLbyXeggwgOwyQSfCXMfIKIkBPYxb/nypM/8096mX
VO+VMv13qGqQEAInZt/thEqI3VBfDo+KKuF6MlQTxjvVfn28wdcnCzkorsPHuvNnJkHq9sppDhEM
RM0kMjW3of1yg4oO5DbPqjHbWFbfp4frz1Dst9/1ixkhlaKGhQC53h7162HQfsV347XRHt9qB8rs
1AeAAL5vK+P0bq3rpiak2COHt5G43u/xIyNU1SLs5mKsxngGz6EkBmUXq7Tp6bjyxYz9JQk6uDpl
tPkF8G+s6CPT0OaHnKat+gldL/ABKt371J+4rUWMqxM7OjMucVD+ZnBY1EgnaKHChpuy5EbCzwZk
HLUj89U/Gp+ge2S27ZLp2SODjPhKELmXo2P3pa74HVdylNU7D0hFE7G8JdHDGoDFEVL7rKKWu8cY
C7LmN5VenyTuDOoOwmE5JJh+Jlm3oVvtYZuOrU70wuwNeY3+q2erEG/afnVXtz9EMoLNtgUk4p8u
Y2jWH6iMBiLajZW9zcgHza7VyUEy8qemzPBSYR3XZksUqR3xvHUALBbbd+C78TR1X3qCOm8sVfeE
h4VpKTkVwaEzqXTzHBcqp9OO1AgWDrn8Ila9s97t4Hq1RTn62wfXo57++GWBJmQ/KqoaUAisImO5
8lGMzYcWRp/axF3BSWXEFqfcoJhffXDwzKbMcvRFWrCphJPpxW7UcmhIu89T6cDpo2B/+By70D/E
UrYLqMBnlOkPnc/xHCdi1hz1xCC/QVSvpFGYf+k9NCfx9sMM7cnoToKPr3ctkURmmSxJhGAHmOfk
hqximRU9uyy3xBBMLu+MBA2Uqblmz02oW0dvvc06kHO5v0njyrhdVD1+q8wUxPnEyeg+449QjKRi
9GwyOgCDwCcTlCYDuY+QKoHmen9vMKx6JhcWd3P1Eql5g7DmETxAsxXgH9ZUFGoM0jfQQkrVBq+X
B6Thg7bha1MOFAmzIrVJB2/8EWBaprt4NqjcavjUcYTRASzbAENyou7WQnQXG3Z1GRr6i8URWRIN
Za3BeOQnVDX7OuSF6eJN/uyVtWLxW9hglBoX21UQMPVkG4rPZKvQ2u112llz3YC2TgZPRq7lpO4Z
9tdUGZycrVpBN3Z9Amyws1UbouNHihNOjkRy2HVyTb2ZTg9fvx6y6rCFd2cMqo1iH3DcQEORMw6y
zrtfZAF4PxdceMZLn+5XqzOvmesJS43R5F1rMsR59t1zuQB9MmdaWBCd3GWUdhSwT83wTvTWn/oB
qvZjtmylDK1atzioRXqTrD4ClvlUKEj2ZM9Nmodluuys/CgOFE6N7NytJ1na7mrodJKu1FTGWNq5
q1/ym8nh99khLJtfmiSvuR78nLwWTxF/TaWBl/eRpUKWWD6WILuCRDBAwb+8jbOiSTnkD20xwGeB
BHw0FdCYkHof4Yzz3IJlndNCjoiq+MDORV/UG56vglGPKuHaVdnxZy422cWTyPIJyHWcQZerZ0Nf
/vvvqAkDSkxH+ERj6Xle/imYi5EqAKBZQTZ6/e/oyyE93btzCjduWkGepZ7gJCl94zQucZz1D3sR
X2tsthVvl4YKMNDjPM2FnK6GeCJJ4nKKVMVM2ObyLH+7Ot6WiYAkJe421w00VzWcc8UNTXqJJY76
m6bXri+n34fqYjrfFqxjnNVEl6qunNEpGDc2SzyhCr9ahE9KzEZJfd4b5lHmZNraAmRKnOP32cJJ
iORgfvIaym5wx8Xp1rdGzSLHLFwwcJjlbMqPbMwTiJ9M/tyijX/ndsB56yz2jiG11WxyH/06TK1S
+gvb/eYcu1gQ4WjJoo/JKP9m2NU0609dlhWm2EXaHbxiWBVkc+2hz65c027UPozK1WuF2V4ry4lu
btgBSQW/QqOYyxS84Y7frx94xkKP4ILf1X8uBGVHcs4KFObQUZInMyLSe3sBl9zLbcFIkX4LMsEh
iCdE/iEHVGHHuskdgHNCD6beMEjS3u+OiV60qZ/a8e1RpMIAXa+moWDPC5P5yB7XWGlBzNlAsHdO
+LStyXYyc7LoQRPjfrmmeTCJkswYuvbdKEM72Tx7Tjn1uSSJkgTTCSCPp2+BXOiH177/F+MVN0yO
kPfQVJJ+yB95oLb6KrvqlVT6KBVWbdWvSp16FzSKrCWOD3fWeo/qliXPNRsSsV0558IMup3ktsTP
/cYJ6FWvxMVlteUng/Kjys5CEHbY5E7q4EMozRT/zqKyXQxEGoqNKqIqMx2wpjFvaVWxJV2EiceM
y9bk6tIil5sndSRXp43WKWgtRIzRrJk9UREOxkFiuN8biQa5jty10rlrJQLGgfHvbuYIvDM/5ntw
z4GVUfOldct1nhrQy/HTGPiYaU3mdmHz9VJud8YnzyVB2dwvgjudcHnCdJh0ZbNnwQrdMt5AVHZV
tHGLVK+senb8w2VwJ36ctHWxiNnrQd8ycCLWddoY4yibVJxi5wYwvuG6I4Dh27KuqvaajedWjBD3
ST4dHY+U79izMlfWqeNi6wu5J/hDYEyewrLFoi4SF0wmBMUHAu4hqgJ9IL3VpO9LCzXFloklHZzf
+RvaGozwi9UZtk9ZYbh6lfou1BkZkI5vnPWcyBZazygUnWYAAADdmjNy595Qq3vUmv5caHNMCcj/
jk3ryDyH7weP5noY7cJNj7ceH5l4UWVMyuBCsFkiYldi81qB/qZJTNB53dVICoanzoZ1MVGiOazb
Idvll4HGo6HFhGJe0cPOKQHjvKVvx4npUDm6sasAXezEbm9wFuoZXhX0FHI0/EhiHBs5w+bVuQ3/
Icbno3gvMMq5PnXFivZUbzjWOITemlkijb5qgrVV0uUU6f9zgNJoE6ulvj7YJikoa6A6yE1mRnKM
LORasvwFoJhwsjQtK2Lb97oLA8u+S/B0k+SN24Uizp8oWz0AOFO76s/0P0wrRBsHvcQJAyLF87wZ
XFXDjUIJiUf9JMFv6S8PmQBHBh0JbTYWTxiI44C5vNsfblFn5cFUDIfzCgpj+S76hP3/e+j6gEr5
s6rc5CpfTtROl7NVVfD7LJ83GGWOS82RW+/LqdNoQOsjZLYIgCF/Mp2n0m2iMgnOuUZueweHhcTe
mUOwVK9/ZUUWTHje346F7YfZsCAl/zAmtffZ99f3IYVOkfxwaRbR7JLz8cZvXcRuon39x73hpKhP
8E+A7yk9/JOa9LiaM7B0Wc03VwAWxGmVCFM8stVymlAo8tCLHRvZEE4IfIJ/Jra1iSj0dL6zXFBJ
q+a62S/o4dR0iqj738hXhDlb5FRLei0G7L8KEu/vRqvlimmBcDIUWA60q1BKZ3O6rXcVSJOxHc29
cNwFY4h1wlPY7J6VjzG+hFP7zj13aX3IPccelifNZq42mkuKjtwopRj5wpM+CmcXV+7AXuDF3Oj5
KdNwWZS/YiklvvvVpMp5mWQWf62GMgPQ/JgxKQu84zqeEE71QSaVXuc/hakHbw+RQkgxPEcT2B5j
Tg2B23Uf1pwYfAIHMqjkpA8W+wCoyEMvC1qumqOSVYLRD+FbDrxbiKFgnxxHO/vMrwnSMXjJrJ6l
IABflvx2afFSj6MYYRAPqgXovYJrUTILoRkdRgdSofcD5mUXx7hTvCXQMwyas5uVqZAz9kKRuoTR
lcF8cpKcAVCjIBOlfGoNTdPpxNy094JwpG1rtdFVq+Ks+sEHCiTWGtI6QUQtEge+D1OZ3o3kLMjT
25Ym4hN4j7fcU+qKGq7lgM82fcsdzYH/XiwFhNhjH9ixBTwXLm22j4oeUz9N3vUlKHEzYPU9XXCe
nzl7TXC9Nm62IXM2GePEz3jOcwNH/gnaABf9HsSLK8zDf0DGitMrgf3rFCBFZMAk6RjI8acjTrBR
tUMd+Ed1RANkYtIxpFa5kpC7+jTk3wSbcfO3GggG/dKTGszacusJVxKRoEcA62PFLRLsZjHpu5u1
OlFcvrb02F3QHS9o6SmywOwYszPwYrv7A8Nm481DZ2/apMtEENAXtKnIF6Qgd6esXU7LBNgyXi5g
QQzpvhw2ZAbSq97NX2Ezas1C326cpz0NB5ZGudkIPPqG9e0tQX1aNggCDM2rlfv5XgI20FISy02j
sxTFOH9G5JabP/IMndnUTUQoZ445PuxzavE7Pp3Ey9Rq+fQBZDoJx620QTOczPHYspbvBtXd+P/k
yr8fi8wcpsPiNUrsCCrIzz80+PMk4oAip6yiZR0eWNYhWrF+oJrSo4Q5M+WyLXYIUcr3edYRkTOb
E+15RQWO0aWvUWiDOFd5wlDmnz223YV61pqjo/a21YRfUYItUv69oNrKKMVk1ZbyhTmtvDvYOGxo
4UodT+lQatQ2GNL+XFtUH0d4fmOq6uxFfONXoqO/uLd3P2/2CgsSqU/ueT8OJkMdzIl4yui9wGcN
mLhRmF7AnTxDTrYnGqrOjn7e3cBR2jDMZ7deL/SU2OdaJJkXXpy1Mik+sGhTge2N+mcPvXo+2NF7
mFxPrCBBABRW9a2YJtPuw9u98BnhHc/YP7vYD+PlWFEiGGI1xB9eVv4ZM8ccHQW+xwQ553yi6UXP
J2YA31A57h8CpoAMBksyB60im6raAWoxF03UGQZFqQXFbR58c06KmGik6FszW1FtweX37lJcVrQP
urHx1Pwlszek2Ga+rvZEJU+8grEMgUT+v8q1v8Am1bPuOcmJeb59dPCzrU45SwlDAZWgH7GpbEIB
vPloLpyvgKjD/yUTdz3QJoXzELjqnENOdXepajLm42jQBnaOcXNDwG8dVjxIxRDxKy7ND/H1rDtw
r/97iNtcykbYTHwtU+AfqI0/jTeLSzONjtXH4f/xv17WFEVX9cgZl78kJ8IhYzvobcSRT/cosmGn
85mtcthUAylAHnYbIIbwIKrvHyPLg1iJPxjN3Df8q3btd4KuYWncBPiGIxF74mjkwLXYbdAbRVwG
kvWmTfGtNA2lu3mOzDYQyyk9/UfnBTSszwC2tIGHycu8VqnCF7N7XmcPlfyB6Zc0BQG1qxJ9j3dI
X92nh4E/v6GciTbm/XxLsee6TzXq1j8w3kGUBXwyjTTOEQ9wkwDi7uvERq1lxiwSONuESCYkZoj4
QJyqbL085C3ggUO9IpwnMVYRVr33gCcGOHaMORM5+TWSEgMi4+3j6EiYYw6iop1kQe6BoTdiM94S
zHGLtvh4PR8FSTV9u2VEqQQ2uCKd9aW/mzPPnSGiq5PmvHZt7YGQJgmBonlgZpg1hmYY0tONu/rg
MxN5aOKtXYeRw38HZtV4qNKeu+Sef1WJ3x4gPFcMp1iYVpJrEgbnpQySqJBLA60fno+BWzxuDlaw
CXm2cENSpTshNnyAqIKxYyo03Jix/KqxGXTGPIuk/Ls+q+KosrlSfE/MHwmtpjhEFSvpNLb9UbZH
LsrI25PteAyN3fUnL73/V1zrq9h4TRJt+3CnVBxvd/5QyITjIrU8HK87/2r0Lpad8wxu6bSe4opy
CVGSYS9PKcrz5ZjIGsS+IQqJs+tUf5PhgSgKru03G7opGs0eUfiLUe2LnXvhYXQRCrqRGNnt/1nY
J0J1fB+aEnI7S+A99/5ksfil5ecchwZR0qonBw9W8t7aDGG8pw/9boNqQF/kbAzQ3iNTJGdsSoGs
FLGTdI5fz1T2+HIvkR2emEEX5Gx+i2mnCimwm7oq2MuMCxCKGFb+mn/kY6sbZDRJjx/1pvIIjmCx
67NaFd2cm6CCTjnlUOK8ffMMLI8JGVJNX4HUGYzXxsh4ENsAmQkyzees2rkbzzMaxyGUKDDXsWnZ
FxaGXsap0AP72sWSxOeTY3AkLY19it/9C4uD/OsABiw379pX7+SavpR2y/82saUb2mUeP3F69i/n
DvuCMUoBCSvJBGd7g8F/AYAxWCXqFdxiUMgnYRQb2av4rur2stV4zU02BEGCJNSNxVA6H5BSMAlY
oKN34SIFS6lIt7ekZURou1/ktAr5Shev/GMapVmhM7TUV8dcE9J4zCQ+glEiX72omTIa6SxDLgJT
3QrvCELV1gtKAXtY9WXhmWvu0+9jpESCZfxCQzIiIJfV3v02v++ajtMBokxR/4ITr8b5o1FtrMLv
HZHKu4BJ4ydYpAZNpRlfYvXUn0q2zdgSBqXLscxxIQdKFAHFDoPRqz3OFPqLwGnSxMGjaWlSucLq
c6ghIuGjliky7dHIxH1CaOjNPaHPjU+VImzJ5JmcSC2/zwyfAT77sSLJ0XeDFps9rFvuHQGBdRTx
drcuA71dtkowbDaS6i4IN8GT7Dp5DtiprJ6zw+gijYnpCi6b1dAeY9L56aS40/mrL9UpMb9XkB2i
GTUXBW5d/32ZZQ/RQbIzXR52KHh13U/ZmngtIxQVfRMhF0ycfPLxzd/S+Laz/juyh+wyxHGwAj2t
MsPF/XtqFO12himB+98fLZFJ0ixqm6NEcY9YSFkR+EpG1U5Lx10iqR2KXZpaERbExKb099LcI5tL
gvYps84AwmK0SeEbkbqp1gYcHQ7fZdaVka4H/pd+Fv6QTKjA2q2ibvuJJXp+IpvXpX33EI8CuMf8
iPM35Wv9j3Lba4VgEoVVtWZAY4O0dhC6lv+Kgi5DyeKWCjSdVe8K7cySQor/L5TFRMeLVvpjruBP
t4U3rG4jeejRakdetpYUF1ARnBRE9Ib3vCQQtLooM0XR6HyhRMmu/7Mz8blhn+hU08kFviSC6OOj
yc0NP/LWUWDB5UxfFEqM5gmilNX5U7YVJrlrMR31jg4a1LW2bZCkmQWc5k+78GSZPjo/Ofr4xkRw
HzVRRNEe8ivFYg0yvzG0Cy31MINhnaugecd2jTu+nka4YiiOoYQXNi5QNYtSyH3VqL9ut/BUJssD
taDEyGFhSvZak7s0d8Y6dBFTgnVR90nmBnMBtobnQXmIb0EL3kKcKlocd56noQsn1F1JevIsmIKk
c2XORPkLb/bikhiH8Q68+avOkld4O/KPdSr5EyJ38vzMgaHtHfQofODLanY9knbSVOrgTphE6Dys
+7clwQWyLj4shhUqo/fvmlK9U8W8ZpYxnBCuOqZ4kMej9m77B0NfCTkxItT79h3BMZgxyTGvhdwl
a1ODS8/18zmaEUT0DSOORG5dBvgHs8L9wtV4pOXRyKcOlWRVSjzknrUtGzar1EI2CeSejCiaGg1r
ITzeMM2SFopHN55Pdhn2v+4VFvEx3xs3GIE6Zfll2wTQ5XxAjVm3zhnwva/SH4ub0H1gIQa3heIf
Bg4QukHfn7WhU3cZOiv48ku+B4sEw4Twh357ZD8ExNN2Y29GIpCAQUk0a/2ximWB2SD+jucUwp0c
K8ym19oHqj/pctPUmf0NDNvWRX3GTzJqy89eJzwkGgcaJwRya86RdEizlbnoUAcksMh8zTVmgN1K
sPVngLTV5taePPEdLJBwEcaP4zzXzST/alcguWChocvNmbACteGs7URT3FOK7ocInqlas3PAjWkD
MhDPTkwJb/EU7455+MqtSVG4JjMPGi5MbSBqaPoJVDGNp84jo/0YX9Jqf0NDmf7Un7YyJ1wkxnIt
asMiwNxfU/sqZZoPrNvwyxEMYfJM2ZP3f7cqE1xM0efBXCxMgkCfttGJ2OrI+jEkDoi9k4bwVNzC
Mi3mDEhFWA8PlYdgtvzUfUaqIJrzEUDhuS8bbVuMwYhWM1oybIzPwApQb+HUWKagNgt/3AckBAWD
DJ/s7NrJhAXUCQNPPQcIenOMSfnSB1q9ESY54AP4Sv63C9pSS9GZLpWJqQgi2RXd5dQjBdp5au8x
EW7VHpne8DZQQl4WASO0r+s7WdaVXYSGZBjHJl1AMdrOkjgfjt6G0I07EjuEwCNXSVG3alPPjuFV
BlvllUVEDUTfBqfgQRjwZu6cIDfKAqp2/uqrpkCT0Xi1bfA356+Wh0AmfBFOfI9QNtdi5cEkGSuB
mwuChzhtdQ9AQ8sJJvMzeL/34pmJFCSlZFGkwPTn8U/AxUgcnwtT0MlKNavil1nLxNPay70Ok0uB
9rj7yunOP4uidosC9I4+dB3G2qyeXRTPrwMMJJIi0uxltVktA5IJBIZMN+JXgcGaq7lX1uSOAWCf
lonRnCaOLucXhGolyX06/59O5GhpRKtXuvdlbvHQdzKL4sIs4xyeeoTrGE9LqMfe60VhPjeSPAYR
ruvT17OnOsyWCwTxi3ZK4LzRBid4BteuXw2SD3EB6OkJEOkpRE2hHwEfpVVhPXuBEQt3nj6deqen
WvfYJhL2ONv2aBCeZ80cch4ZmBRXPJYncueVg18KnlCugc85Dty5soTSWu91ax3V2dyXdsyuXK07
Xu+rr0Czu1Rclq+dIK87EahzgSAL3SxclbuNRal2Qv/ha/3oSTgmCBVNMYo8eAIgglO9fu39Ribq
6HFIMIgoNrszHsECnk2bVNsUF4HsfQ85eWQ1gaMNNIP7seJ600lhwS1OI2HJ8Zv8Cj58OG/LVF6/
d3LgpWraOwKcL1xJLhY0Au3p7SuFNWT5fKEUQITBzgUjSOyrH5aoaf7s0Nq6Q3PKL4yudABzbdSL
UgFsUs1hqN5FeImfVmUuOTvoj+qnG0HtyN5IQrasa3ambhU0mzerHFRbop+fkPW7vOYevjvxFX3k
lXk2Bz8gsETHHx297+cujVSv0Qxb6VZSpgVKFbzkPtc4vHSXGbjyHxgCSd67WrV0Lt/LyG/52TXo
k9KwOYSAX8vD8gRsCPouPGquSWWZ2t36xk6x/vckXg4JX6xhUuvfl/8KnEi6XAUOPVQDuWVcqL6J
lCARHuUMHxagH+sg08u/aPwoxTuFSWvWkRoIRF6NtTO8FseKMrSvv6xBrZySVxc8JNIe1Q/ANyi9
GNkshf4PZQJlGvv56TZzHka5ruEI5C/6Iqd4IVke6EYgvAMHU8usKU43DYIk5UbZ5IbKb1hBHgMV
VXT9PszTrIrFk0q6C5e7hNLik0JbtyNZTK6GwA5BBWJJ9eyTqKF8hUMCCSsV2XxwQ3KxnCelG2F+
T4np9F/lcIk/A0pOot9bdZbZDkXd2CtbYESsep7gqrdYdwXxklVXABRSzAbAoXPn0Ipi65KQN+7a
HhPlW5Ku24TcvGe0zcEOUZA19ZQ3Pfk+bfsT6nrv8v4fJbEktp6+wnRlQeXbCiu2dwsGYmS0uaDl
XZQAlZifAzZgwpOH1tLlybVAcUGFquXn5IRL+83qYddnMi6vI8Mf7Xkk6/3VnpwyNWI/cqyd1aLp
YymhZgxPClWt4eBYvCKI3UBy0jEx9GSXymvMS/pjzQgdoL6Ht8eyeeT54uN26xre908HvUimv10J
UO8wXlbuKOqR47hDQs3DvVCRAGK8qgyRDmAN4MsWOSsjHB0EMlvJCAey+opONfEJ2P7vOzJ6mXuU
dE0m84wkPt9RlHwNnuwRdlaKKiXPTg5t0eJ5s3m3q/jYyL2IqnxcOFO/hP+DvxvaJUGx3Fe9fR16
GcIBGxqKgiOzGCyEooE4eLB8eeiELIkPGWF8DTEPSyBu4rAG7KPR2Y1Ph+3/318hW35MjWTAGVUX
KeijIQmeTyNAtpdcFMcR1CR1I1Xfpj2WuwEsAn4SqIj86N0YfVTYHcZkr+qEemgRXbvWQYlIZtjp
hJz7Al5lpRioGaO3L/0mIQzDr6W6i2HXXIGDBy+W5oW07xb0Z2AUaeeGlNiA6ZS7taeJ6eKxnJAC
M79frZ6VlEMoMXRmzMGLtbLpPVWWeCCqOJQM2PBdOaFmEfuv9EIpvlaQjw+CaCHyOLBMgCO9YvRs
fsDGxr+wnYK516tsgdNEfawoGHnCeVIOdNO0rX+sf5MnqtBO2/u/Im7Pmh3G5iszX1nrlV1q9g8h
Hk/7LnPTIFGoy3Q7TIKqcjTnYK9C+0DusXAYh1yuUNN2ttpRa9LJTKIZ9/U/SQeVNK1l7AVJchCD
7FuT29IlxfWRbQOc3cCICTkNfTeSRMoFHBgPqpvnS0QWnOxXDQUGy3liYFa89TcVXxO6Vh/TaVsl
GQ5uX8PD96+iiovbJymD2JWeU2A7rN3TTbbyZob8YA/1TYSjgq4i/08YWBCR0ste5pgLs0aWdzi9
cb4H5h32ix/sSFvgN66sULXC/lXZveDOX/reOK8nbpd9CtGIRHOeCrvvSSHNdUmdoPj22FDn7VSm
yBGkl5WM+fqxyB77kKSozX3NjSQTL0fC5sSln2kOgmaBV/cMxunJqdq29J1D8Mys2bh5fM7lGDCi
0guUtVERB+Jb5U8mMT9UkC6gJ8+1iLXkCbzl0DB0EjuUEHewrv7JwJ6JKk+BRnb4n5YqyCSIKmv6
ZwPLbAuupN+LIH1PoQvmOidrL3S18E3fSQUJn5abvvnvZBn+Zl69W5Uz9Ng/NNroIA0OmEbkx5C6
jhii9wGV6Soq8WJejyIXdOMTG505ASKWCBWZJ78o9MX+PCzfzxpJZqoIpWqcpraS6CjClj1swQaU
cuwlLzNtyIgVceOd43QOOkceVvx25WE1QbEkMPW4YWa2bDC4KwyxHcBTzX1XX72bor79c5ILU+5x
hYOI3+QwfdC/gNDP9y9vTDR9UNOmCLqTGhBlGMjv5ewsENpJiHwPWrzdxdixv96u8UjC6V7WT07M
9DT07Dz0c6GMTeRatHBekjZbsolZujrPWOSckUGtc1zLkgUXJIQRkCR7npHBuE1zmjtkaGIEmDxf
WiTprz9RR5yKOGI8CW7qDcWJNCja1FteuEYAEGT/34lubvsliIN6tMWwmr/nT+ttmtsyhr31wA1g
EK147fr5RiuzPEscT5mR2G+TEPLuoeoCZ+fcLCMPaBPFKrqBKhRWtVn31KzkbZLzFj2fxLND+DTs
ZiTg8TAS3qxfnxoGhQlkuO3j/2fpxozQ/8VXzTIbz10nUS11daKtJoRWHKpRhxY0HOKVY0s1I58W
yFuiOszpzqc7ZhAzZTsmpyDItyL6lMEZauLfU52hynUNxrQefdeW7gWsf63s0/MYIszRlkZv5pAM
NStMDt8SkeQMq37ocgVGxnFHWm/qmIShF+A16bM9nKQfZeq71l3LKHes8x2ymGg1mrZFQtGbHH0G
KHflce0LxH6nyVGP9HMZpnGdRFgoa3/fzEfZJEM/sInMLqAmwrnuFRxwzEJIqJbWTtd6+becZbC6
J36YUa+XiatYuChZjX/gOYUByEfNtVRLVOWDV+BId8Ec3QsYO4vXFneGr2+eJ0gwTX5kPFeRX9/i
1V5A/qFjsQa94+AISrcVrApshmImWiabtJKDl7iyknfn56+MS3fADhbmAK0tkmr0LV5nkWBH0rmI
J+WofbM1rmdtm19Tk7IfXQCR4yrW3ya9r2UDx8W/RzWtzaptgy//K2M6GDxWspaa2bkTZiuHvOWn
MeAoPKz0WcpkLayrhiiCYygDRg9IWezbUxFUcggZYyoYndXUs0UBWHk4IJm+61w5p9PeqekUZEx1
ZMUl/Qi9VH5YgiDoVoIbBzJBdOhF9/LX1+MsZjW1qCkcozWh+DLB8wwpLq0Py4jjyetzM0GazHQR
gFXls1zZAg8pg2XDLbyQtS4sm1Dm9qU8EjPQKY0S8thRRpWB6MSBSZ0H84/ZhEvWSfPr+qmVYbcY
BwqrwjXnZp1RNLC4BySp5e1frFx0CFFXJ+4P4AVAX0pv6TG+iNcO9FzufftB7kO8yhuLOotv97C3
CuTplIYz2BVbfPsFdTFxvnrUUrJSvIchPbqPhTfN1YEx2xyLX7gi2g6sKUVb+NZqTOjLqlKSyLsZ
ra4CUvP0RPhF/Afgw9zckCSrpFg3Yag4DSpVStb6EeOK5F70+yRmeC+Vmd2L98oQL0nHjeoY+XkG
SQwcYi150CSEcmN0V4Z4Pev9aof+TTvTw/Wfolezh4RDOJ7VHpahUP6u5x7gGLqiHrENreQijNs0
I3Z9ZIYC4gfhfZHl8xJqo8rZLcPadEHazQrSBMs7hFnw1nzE6M0koC5ynHf2qj1/42gnzpZZtHd2
o18mpfdCPpvYnj4oC1+4nlWj8EXRePEg8CgeILRXZMrU1eU4L0Jvah8cH5cZDaPo2B7goZDkAT9w
t8XH8gfAFions4qXsbC3WhpaZBr+nz65mtIrpa6se/GAL+qRTfYaJ09gnukaWIS44YoqlwI84E5N
kbJ3SJMnyzX4VH9VOJSafwR725japR5YfeQnHfjuEWuer9lgEpsQSGJa7pHCc/iYva6TO0KqyMn1
bDZiUxDpAapaRrLVLPukRGo6ZlLJyHK2ohX5VsZvT01WpL2uAwyw9XNtyiGffC9l9IiQXhnKqj25
0FCa3yJ0pPwmFkrRJu66UvNSiKSvq0QzRCj5T2LmEhhZP1i25L6yWZ1jNH5H4nYM+ONeXX3zoJBs
3OiCP6qHDU7+uvRRLPose5A+8mh6MJcjSLiE7m+7YkKmrbEVh9uhdqffrwdoavtAMKMafiIzgQpa
2KPLbzYzeQlFWWpdVhWaTnuxx+o5FVEmOvv9ILRiue6oLw1/nn0C++HRYLa0q5XZkhKJu5t2Llfg
kzVt8KRrXLz4rNY2bmnLMm3A9050D23p+Dn88JlE4qgNZTND5A+Xt+SzfnKh6cOQ4hS2BjR6UtpD
FDKAgIZS8mPlIworI4e/Eit7xYCk0Zv3DZcAqcdD/P/y04rL0nzouuCQppJsV8OkhKh7akzE/EHX
tA9vy8ugQttBTjat1MIYeF1yApcUOjlVN41hJhMwkAqIHQ/l/+FlgljCuSSF8y4TkzPaaUOosN/m
8/3qK6O1ZbBNdDS787Ljkk2YGVAmxSoRM26rNLkWv5FixoEWFmKwXD3LDxE53Fki8w9O6e9qDDjp
AP7VrNP1Ffed0czpfICMU2daDD/Bs+gVGOtlT211rdadmaySz+cC7VfYWWfqlqSbqcLdYHttqiW1
Pae6vVr6lnALY4yv//E98Ib1kpPkInodS+WRH768pf+2XbNiRSUGyORVvazE0TFXvRzYuuK5512W
Oe3GTmyAKRqfb0oozqwcpJzp8V899CVHXa7XEJmwsQmAonMU+xtF5bn5TmtFgg+NsTqev4rZ927Z
M224HTqWSh5WbSOn+FpV9bNtRhU6M40SfKLrUDHGsZd1NSzxMMHx+VD62g5Tb28ZK8GzX1ibXRyz
OkH5TM7o0WsS5pPZNXAyx6ynOYShkFh9hArpinrYKC7iVVCnN0uB4M71KYPzfWlNCqRXlPMVBtdE
mKMbUNcX5tn5aFI/8wEQr8R1wvU0x17Re8+dyRqzGCMig46Vv+KRj5S55WlbxYDZhfmLbjZq96f3
uYnAj25pkUxapjinxThTMG32X3XjVtEXjFpWDkBvC8LzrcnmJfO6VUFF4OQMGmrFBsfz0g6q2XzN
XFNYt4xNwJ5OK/bMTN/kwOztuzquPk7/PmtL4N5aNo+XvZPDR2ZuN0RyNYqdBQmMyNU0jwXfQcQy
30cosQw2Eo/VCRJb003RSnyzMs+zWdNkZJoPe0h4/PAd95QWjX8E07vk4LOgAIsBwTYrLwgUH8DU
1kvid4boIaUycPZFP1K+s5oc6r/7lE0Nw2mYiM1px8IF8fHobRS8QIS5Z9fZu73ZvaIlTNwLXCiT
Qaz0QmOIi7xfgQ4kwX1kyY7p5ceM6JNIiJLp8SbFdqyjAHMPec5egnQ4/0ACPAsgyN6IaQiBCtt1
GkexmtG+8KI5CxCDhFhJgEeFNGOGULwCQ9yiXODNLSJl4NRB6sLS57JMSuU3uRvHZH2P4u4TyvK0
YyFtXoXOO5xUbcfyynrxZjj/va25ocbMv7zsF8l8qp6mGVsmf586FKSqyROt+RYtllJvlw7zIPiq
6zIZWXO8NFHtINZxrwtJrcL/UV4anxLMIhqo6WhJi8IX25GwtEBjm4c4RteLxKR/WOQTdpcjzxYj
5dTXMk2R9XFkEsHmeSRGBSzmdt0hbL3LGdcXaw2m8L/ZnYXffymBaiUu8sane5Qr1x/3HjOmWilC
8v0/UfN3d3GxRhnRyue2h6V1Zs14UAqfvK/0xnCNHbj/4fnOe74YBHPy08f3tvLMPVvlnrjSRX7t
Z2sJ88pp7R1PDNV/pJ4uCZ2F4gpLMKXW9XgeILKXwO5842HQzaKRcMKIOJ4JGIDg0EZkz8H2T+KL
8QSTB93jXUwdgy31KUqahG34RqUbUKqjxOHc0+U0e0G7JSEEpUV1BoGLg+qeSuqGmu1Dg43lx1QK
6ngb025ZTyWGwBxU1OcygaC8qq+FV7Jm5+0SpYP3Sl/O+z5mN127IaJoM7Bo1B6g/5POYNYwsZep
TnYa3MY4B3jvNzrwHUv2HnP065pFAMfKt29NyToc6AZqpEUA8CrxUr4/o4fOMl/8cmrXWALbVq3Z
9Uf9FIx46IkhJ+QSi0x0WmV9AEHJlxczy5RrcrhK2KK7bIKwUw737qmnT+Q4BIkO5iu1x5zfXCls
n4q4/LLbCHKfX/cMP2Z0BbFJi4DyMqSUxkS7gvF7fg5kaWNha+nbGK8X/aR40cw0OpdoSskjibyf
lsCMTIQg/xMBs/x/+jVLoDcWzEMVJPwLRy4jirfLkt9IokoutXD3tDdpE9QOekh1o3lWexOWkXq1
GjVHs7fYtcrvsI4Jggk9ygvPCWwNW4hwS0jEuSQq9+e2CLfS3ULmYbRJ9DYoNNoe33iDQs8EXmjg
lWPdf/XqJLPaS3NmrBd/LLhhIXcpyTcdHom48vQbhVqhlHqmTAow0GV+mS4ypsH65BwTTh8LXECm
V570du8GK0wGk7B6VkjkFHkdjDa7TzsD/oRFacCIlqBwoUuD4dnQCfX7pobGpQsAzcdHeVWcedgT
YJlGNC04HxITcGJDK5Goctpx2jFPiQfkDQALZhQbn+W7X9pvWDoDO223W5wfAR/eO/9bH+N4vCUc
RylckJzAmgwaeniAW8exrSNuA8spfaUjDI9K6L8USvA02wvVGl8EY9hzdl5ctr8MaGjwvlNbLrcw
yzVRs37g/hFQznfk1h4kkNF5QK+he5fiGFcD8tLB3cYStLBC5ECtBW5A7g9GwV/MGlaL+WCNyMu4
SuLATJkWnV9CHBUTYkXpMy1MbwXu8s4BOD/+yqjpFq70YJMxHZ8LqaMxGnC+GAQnoQL4G7TT0Vzh
dUwU0pTvdBSLMwwaV6a+OaHBYYqL+/oPY6GqZigMJ/01HRcH9BBOkilp4kEAZx8hP+MnG/rG6KPV
c8aI6gyTIWRw7yltzk2Xd7T9HsQyKgTefyYktIpn7f5CAPzJlxWZlE+XEoeCQ35wNkafbPs4+mgw
c8Hg1npAhKrlDcKe5/3Ws+vnaaITHz/5EsAgWfOmwDxxi0bz5cn6QyGKChoodK4zJD0kqxZFRaHx
oin9oTYWgVkzStimGuEgTK1iC+YKVPSDY0paZ4xqxxQ6jgyqFzmvwyhkchRIfJA9veMAGndBmhLF
Y2sWnLNtA18W6C2xnBii6oq7l/tuu2PplpwBFntm5vJhjbYEX01tLjVteuCECpHBuqnvSzFxXDnI
YuoxG1U5/2lbnxNYLiNLMhYHQeku4oDJRxXAcBM6Dwz7VZF1Rsw8y6LvE7Tj7GyTCjdP04nYE7SJ
poRCi1iBy8mVRwJV6jtJoGRsP8jxn2Gbup3PUwamVXTJethacRtTJ9vzdeJ6hANyU5XUVL8fT/7/
H8CZYteCLE48qvmKTFBt+x8ZKzAzXAmFS8iTNTBqtmK1Ydi1PmLlEaGgDyr2eLo6nVJ3fG/FdunB
kFYt6F6yHv2cg7TWp64kgEhojgqbQDlyImP+S2OqEgRqrwlugF0XbpQceSQabrj+5U55PoGxAd1I
FVGtlgallRg3ofZ+9vStCnYjs/aNDUbt5B21MzGP8zZOxBeVFV3sfD9PKrvIZiefAkI/3vMNh5jB
NjGxm69K63tB0sa64Jb5RwqXCFtkCcWP0KujvQE3NyvnzejOwX/0PzM65yaRaNfOzcqoYTp9iWUN
pFUx4DMSLDv3duONGxl03HjvrGjCFrdkYNGNHdz4UwxQRqNZRp7a6eDXXIxehk3k+u/ahThHZhvF
oTIn7yInP8TEEeSxfDVGElQbMrO92SWjm/X/w+1w6J0NASH1l+VZ+57GHtDxiCxpFTjNn/l5Yw4P
ea7qSk64qGhmA0ptfy9u74gWnuGpK5m/HtkqWNy0RbeMYgagN2FPCRNwzX8mrHxA7vuxHsndP4Wz
KUvgSX4nZrh60dIZsuGPZ8DGV/lBoIJbgyD+o9Cr7KdwiSngJovryJgkHSKyboeGPK2Tlcl9YivC
tPwNM0ZaFY5NxmOlMblZkLtlDY5eUgT4jfxU2XjIDTKhOuQngi4u5bgwWeffQu3emsDEbc3Gwd83
fgaeGo7mCybXkyiPJl9S9XbtuNLqESG5YzR/NQ9oAv6suWXP7O35+7ySOTyP+8NIxxYyptD8d3q9
bWkm4G+HyfqeFylwy8YhxGqTTrraJrT1tceYrO+BO05Uq+wkurbj2HJLMdua0KXncK1GHjTHUukk
6UMPBoXXNztEDx5JxDTX0PCXQbkuEL6oRWhWNfmM3p4OTvVDb58SgPWPOnXHcl1ckLTHTZ0cFfBn
CJhYyUaXe4mql+OlF6NpdX1oVuoYaCDmYzFPai2taKu3fJbJWgXNxsymxF4Vw0tl3YajbnN3BrIZ
xz4cVSZx+W1sSPxY0GKQZkGRJnIIpKO63+zDjYVk9SUqk6nwVRLNRTb8SvYH1nbQQA0+0gGK8N/R
9gZ2UvJtUDV4WguVf7y40qszJ2W0WK32QC+MYKgP3ovMRLmNVoY6wqlD6t4jczd1FXILfT6aRVmh
K9eOcRgNbv0SCIOWHusReUZeLxfl/293cmBOq0ZWsj7I6qHzvDtj6Ky2banirj+6oKN+wtwJZOOx
srudJpEmiz8JFyGoBjxjv/fboz+4DF1rtZ6nYfjeItY78AD4k7DLE5HZWwxQiW8Ibln+XDP2v0En
IINvnxRDWPiMCA3A0pnqHsQ0ipsIabwFQDjTB+E7KA==
`protect end_protected
