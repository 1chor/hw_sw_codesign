-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
la5lNQ6R0DwOeCja7zZpm3Rb/QsYn13tzWn9sdfm1udfZah36rPyHSVEaiY+sRVW
hqelMKHw6H84X2N/Iwi9reIpHJNJbuAHO5LDxdOoUclM/6MufebRq1k/U38Pn+zq
F0Hfg90b07uxrcWDbtpHy29CNOqq6uYVYN7xwO/1duUjlqwpm+0RRQ==
--pragma protect end_key_block
--pragma protect digest_block
wPClxcff+mQUpcEg1rXKSZawqfg=
--pragma protect end_digest_block
--pragma protect data_block
SKbk3ppAYtMKCrMgBOYwtIwfEGjJwaLVDHb3IcIxt4KFv0XiNGfWQJ6M7Hyk4mFz
MuNlF+oNm6BxaHojdBHI7AKmvVVFFGI4KURGW88jDM6JEcO1XsSBkIqPpqKbEjVe
x1+P2Af7BMYIc0Lgoy/nLoPsmfEXSkvFSBfK7tJ/gI0I4wcve04BJNx9ub98j9Ce
9ynJa1OJB4pdW96RIO7sf0dMwYiBlB23bjEHlWteBZpyNGpBRS9ap67I7bnlKVes
2NRfq3IrAwCxsStQrJUmszeC91GpeMZl/wUb9yvh/bN1vlGN/jlw1njwHPP93IM3
XC+AQwQhbDfNihYVuMJkOL5DBT/iGJIlqqCvAUr1ELhKB+VR1/GLIDjyDWZ8iznV
xg5twDMXK2uf6x0LHJ2tBpcwjMDpkBaGnLVXtLWd5kCl9UABml4bZhO8drmyN0oi
T/gtgNQL+sqXF+LXW+nmrp+ir+IWPKwDmhk1rCDoQTzYjb1kp0bUm3JrrijOkLNe
+7/1ggnlvhN0snaNGpX0MgYJMCf41Vt3aMwbf31oFd18z+mjqEU2DC7rEJIM+bPQ
pKwUtLhfCO6nzAKQDMm8u/kz4TwLC/wgk4M2PML+Omz/X8rJK0EW0yNIBu3O1mXv
cOTMMeCVG/brgx9Fc4/J+Gg7xkStjEeck1G1eg7hNOpyZruaqJzCebI+XnwyJwns
Sjwfpiu95O/EbG5eDmHAGELLTs0XxuiM6bKe7SowYznTsIauFEfb63XnyrU0dtvN
jLR7vt9w/UPtY7TX5edIORUMLxWmFPaPywqVDO+ZD1xvqjXcC503+YqsBzeIc1AJ
GLH1w0uQEM7Lf1jT4mdW9qtcqt0650lXO5goVDOhXLOwytI4MIESegLsCovCZMUs
eaaM3THym8NurVfrcYGbpPlpB2VDFoBcTN8IY1eCBDkikcEXmXURfCvWfXNJ8ofu
wYXdBdvzeCBQR9B9dvS9rYz/bv5zpmLjONguKDm6YIe7aSWwNdvxTbCTTySqGAPC
3QnI+aov+6dwNcesHU4TURp+kkMtHwgaKEnXtJZqvNViBP7t4TO/RkW8BOqStKzT
JR0ciP1mb9TA+iBGnD5KcNeLE//NQUtKeomiOXfODQiHNYIh3ADjEN3d9fy1PsGe
soJdquOSeDrzul0SIzgawryGTcf6R9eM6MAZn7rwgN9hW9mkDnxuqeu/dRn7HJCi
5gIcG+h/Ljl2rTCMxeEGSfDXIR/lb/oSO9USF9swFa4/jVWkMogGjCOc7sWqOh3a
jgVRfxO1t6IIEoUKKgNCY29AzCJRJ3te3KyaFHVLRS/Y6jEfuslYjw3KF1jt+Pb0
ssZ8fA0KJYqDbjyt6Mh1ydQZW1RWZHD2raP70aer6wGU+njEcWKfmJz1hz6QU63d
hT6viO7F2VUQ4ROA3ELA2Mqta7Bsk1FtWzk5mhmSsKP+KC9LKq9/SdiYi31gppkh
RasauIWcdlBF1RgtSIAJgcCU9UUZABpkaC+jShK9DIby3UxYG4KRUeN+fBJn7ZKo
Gd/91zdtAcwK3NAeOI0czAU+NPdtYLXW7A06JW6TP2Vp+TfY+vOQcWJi60dXPeAT
NdSSUTrET860wptGJYp+5vTgDFZm5CrRsUBoyuZUnHSq3kp2/4oRZrp2Ktx5BEDd
gZUz8gdHbNq+EyLagOI0vWZqLHtAPPa6VoiSVM95qPfVTbGyJVFyzly4g1DlhDtg
0ar4tJt6CFBJHsGg8vM+O8fvNAr4fXU4z3swNBymiSvh1buUedpjJZiK64DFl2Xi
eILmx4AGceKERkTywYe6S7CTE1F5QUvFn64zIceYlzd1+X9RmE1MU/sw1Drj3R+V
h1QCHuJkMzM0K0cereUV10tzBOD7VfBbZt5vgBeaKCbhW2VH7gVAoGvLh+EXP/Up
FeIK9WCX6q50L0+74RZLQHTindmu4UbIBXDWvjkWjgU9e2USNNHB0ruB3aWrYp1L
CvRzWDUjC9DL9iOmK/9x8kkX1lKWRd93LegMwEKerDkw6R3zL2MGVJIlgA72I7uP
Y3BRjzNaYTzJtWY/Cq5tOMy/DCviWMlmnJ6KTa8rbdg1SXO2q89sThwxj1XvIkLv
kHu+PpcTg7QsY54cv5dMJW+EX3+DIWw8HjHmbpD2ejN04CRyWBtBiSS7PTi8GSsB
fVMVIUCjoyEW72FNTfcrHcOY3YAWGj2x6KsdL7j6TO65sfxhH1/5chOvuzOI25bF
niofsABXGohcQo1eempRKxsnJEvcKzSOOkK7Fb7MlCPTXLciHMZEPt9nZCOFtF5Y
GndJaOFPab0lQx6Zjk65hnZYwb+ffJ42H4rkJwfs1bi9NcskSN806e+4HCFwZtbl
c7g9R2+C2rb7RhtCgKuZMSihu6kwgEz0us0qoyoTjtQkMYOQXmDGGKEL66LJEIFz
5GbVmZnvUr3RL0DySeXDZrefCQmNxOs+/cAwcsI6DV3OH6BGmXUpUYlZwqfjUPko
NATKLRDYvX4f2ZmGrfHLnNbwjj+KwcfK2QDEWmxJaVfiR61fu+VMnJz93gC2umsV
oHlJfAgSfoFd8DVLLUcNb1wYDE9cUHjjlrZpdRLXbe0Q3PveRkbgnccTtibV6qCQ
hM5/DsoFz+Uwe48YG7K9g5463R1NEQ0nrH35zJ5M4Gslw+IUT+6cgG24N4QlKfqj
LFtjjKyxU34HnN1ODdYtXN24tfQUz0x5LACXO8pOxcfhsr3iMRRh3DheaC1WraL9
ysFrv1LIvKw8s3VO4DKM1cNyKg2EB9b0YlvHAKaCu8rf/ddkvmzptXNw7/AoK1vU
j38zWvHilu65ZlnFmsp9q4G63PKWdTdOpi7ShX0YBQPwybOvg/gpMD1sV/XFtKCv
LZHoL6UhvopVwTvHt1VyxqATMc7hYbLkGHL88Itvra/snunJEn+/jnVCctDcwK2T
baKrq6qv6pOJyk7RmRaztgArRqzS5pXccpS5NasGU+XO/fF7A37HAcD0rk86hg6V
PftKPdNxy5p/z5AlLBhRFM9FPKW95h/xg/9+eLJJ4+WM48lz3VIndI/qN1oraRMS
UOPCn18h+SAXHJrZNoY48+NZHETbGrDqrqqL7P/sHptZG0EHe8vqEsG1FKCXjPVf
8yvhVVw66x9myi1RJ6MBfrMbL1ko16swbm/frnUFvagaoEqvvFmiBl/uoMAgSPoX
7vds8VwMEn+gqCcHKRz2e8ry1pxrRH7g33i/xctPmjaLFOvZV1VBhsixSOC90/n2
3vRgfLFnJMkNzFBtvtOxJgwRFTRBxpu2i7GGHd+qZBU/hVMIuNMZ7dpzfQYdr1yT
TOOkPt9W5C0RoPI7GfxrYlgzoYadGXR090rLB75vflurHawzNU5Q4axWRMulycyZ
UkuA11awEibID6kxPp4IWM2j7zBLAVTssYKXQgYux4gBal4DB737YXOxI7+yhYq5
CzxgYMNfZizYga106piZqHb5GuGhT6gApNYsFufGBNhKLzVigvcDLktM3m3L4NsY
uNOkUYDHsLBYGSUQdRK9dmPvRUJbUYmmJd8QwJgH0yk7HG/moYP7cYQt84oRt433
xQt3zgAgzqmlC1ecV6cRB87SO08pJ5tIE9fVGVVWvcgNk+4jHYRxPBibcymQQ9a1
O5CZLOAvSO41pc8Oky/pkafmV+ZWc5kP8Jci1dzSMvKX7GlJA1IYBqBJqunSxhS+
iXuoStp+3MLXCSLxLS1g8kgiRiUa0UJaG1RGgwQpN95H2fvXyKP3OL5yplze8Dtf
qBsrJ+XkuIUTPuAWLaUibZR2A8pE20nGZexWpkmlF3WAZdwe2EuwgMV3IMyMmmsH
x5jmtkeYIbNHU0otBKdeQuxyWVza+jl/+d8yMhTQk1ePaDTgJLYadANSc7zpVIh0
t8bOsYELO1Tc2kf3CGuMAgyRgrWg3CJuGLSl0lZO5kGBTjSEI7CMNDnk/tlfTgW2
Vu1go3AGzqioWJbIwTz1GDYFlb2HSxLjakWAqkoMq+A4P5TiEtGZr7Ub/MHg2IbH
nTgOUsm4ptvzZA6E7eeamgwdj/DXFYGM3aL0sOv4aE8cmWVyCyot/EHaOVJHpToa
Ey4L9D5FthN355mBnPy2NiSnvvGDRlR0AgOP0Jgz1nUyoZfNk61mPhhvGA57cPdt
kRZ2FBlXHhnI/GMnocUXgv8lDjdCR3FyAftp0BcnYiiOZbFNXvxnXtOOVkiHKTJk
P7hhXfBkT3G/N77gaRBtvCDf75GWVH+WeCP+p/AisFORsg2okv1RNwsQiffinrnr
sBbdXgzxhjIdFRksbrgXWs+YgBrK5XmBiaAYSGfoNSKFUW299eDubIbdJMrNM1hH
dBYGTjIxplMtEtkVfxax6/V/KLHhh65vHlc22VR18dJG3M0ce6kQrjKlVXlF3hUL
j5hYmvEgJFhthEZAaOcLAC7nlpYLRxhrVq0jS/AyHFI24yuZjRfSYam4dmJVVthv
2Pr7sI+z80GFvoL/AhiuOv15snKuBNCxghXrbTG5yAZZnUhDNbnjLfCbkAPPeMjT
wCewWT4OwV3GMkF7Lfq4VLwcMKgwgPTcY3mZb0bJfDG9Hr9r2LwQabDB5SS9fH1M
/arVi29ZHNWzZZngNXxbmoFMEOFjM+CI/708o1+AAY0Xq0605DEg/yOzOSyj11fl
b4wmjvuwyaF9Gcv8+yuwM9gff1oi8qBmoZlFr+5uU25ZD63pz8s/Zl0xYDulZ7k6
/sw0qK63ZUOQzXAast76+MmHvPeIhFJaVM7OJslSEM2GUWD8+JGLvAuMh7boea75
ryMOURWMOq7FVrYaoZNY/LleI7duquShPYti/c5pWWLLLmxxriZ2keLIz0zvoD+r
QOzpn1O10NpPLnBG8oBpWrwozp5TUb0y0frgbUmg2Mjzmo2Lp2azMTD7sy93dU0i
VE6H1LfpzO4BZEc0M6BtUXIWAQ+d61KEdi521vBIhNVQM3FXkT7fycLHuCps1ax2
YfUHHpSb2OiOqrAMw9gRRlkEq+lRJVKNiSC/ljVbzZgOehWcIbHxE5KYsxMHrVt9
F02IbkiJSbFs6PFMB7nCEqZ5fsprRKAQz+Ap5Cfhc1MFf00qCrT87JbZ4UihJMsg
M2qLG29XYcgG53kBd8B3rnqZ+HEWxWMKpdP9i4C8cdLPDAlLpX633WS3ZTcFv5+L
I5KCqZL1rErfOln8o3SXf+wvkwCKWiGhhVCjz6B1ceVs5D+F7EcOSIH263kCAL+z
7kxJGAygTl5j5tlu5vZiw0PfO+1jfvh0dYSuuEf/0UWFzZhSckybZP58zMuFwj3L
tBiwrKOk0p5iad2Szdk3x8Q3hvI5Al4vie5J7rqTcHJFKeRTC/v16u0xUw4t604s
hPVlb/RqUfdBhhd0MkTgKlZ+CwPSKJBY3qQwazT1KpJkrSEvHjgi1AN3DQHLMGSX
JAvdBOmr/ddXKW24nIO9m3xZDJT2RvYNu390dYu9Y1J2WQ8RDNugDo1fYysaVBwl
2lFuSofKHs+FQ0cfVzX903CKD108hYJqahSeJlt/A1Q0p2oGLTyZouu2yYa7vdzR
l1aPHDh73J+UTxEroLj0e7JKWS39EaDd/n+DtOdWiWm63dobRujThxQ7/LJMw0/G
c6vQoZZBTfUpfgXQ8z4HyMNPKv2V+j6dVEzaSgFz0gV6YT/9eUMxPjSn9PajAYii
o62ya4o7v0kpPIK4h9Pr2EbuJQ1Tu4LcuplCMNtum9y7HvhbaEWaLRO13lw9S5ON
h29cDCgV9f3JIHsBujM//oRog86UJj0RkHp26MW3HEqeYiIPaswDo+bBk/xqvVnB
V7366IZRZl2hQVlBOXsM86T74ELBea8HRF3eyTo9GJY5ACt8l7/4h3RAlepZ/H5V
1eaRtcmb19XBq8/NnLKEOcn6vzo7nvQ6py3cUztQZHt2NmCngdUml/NVGkoIX6kL
ScpbcF+ZKfr1HOQedWsLYaTNKwwj1O2L1Uix8Uaz2ckVUszhJdrMv7KSdi4p4aJB
lkVN5XZgiirDmlIXAiEidvVW19BL0bWiagKmvQDGIPqQGLJpl/GuUEve5KIXUuS7
gJ0EJaxEC/L2xqir3k7mq39/CHfCezpaqFfqMzlxEBCJ1BP/V8ljCpnt2IZsXFJ7
HKAplmKeriat3eCJ9cuUtcMBQRHGOD2HnoIOyGzpqYucuY8iJu4QzOYlTtVfb9bC
3K1kLYWSiNt2a8SFu3cOlvxMCG6VQwXYHnCRcrLjqY+k9dHCPQgJlV/8X2Q58uZT
0srxFrVr8v/LntxzVuwIYiz9XhpWUlECZgVP4Xt3f+1L7kVsyVTjhPL2JY2N9hSm
iBJqGJDVIBkDV9bxo16k1/+FFWXUybpg0mvea6LB7bPAY1vqkzTc3m20RKH72eqg
AaERpttd2KQ2ZS3x91jSr+xmDgv63XbfY4wdtDSAerolt2fbSgkue/zAqP/4BUAm
RRC7ihMvJVsuSWfmZ8kng5Rq8VjtnGSL4VcEqk/QxcgoUgmaO7tIFgRCrqYf/zwZ
06SMM6VcSxgPmlOGLxNiXdeF5xq0dQQQAaq4X/H/qPVFL930Xg8F4HMWiMx8aWmc
PHn+hzf8SP+XJb0acGfwxb/dT+mOHPvB6ztKdzk9Rcrw9lIBUa0hLJOiAmSJE2yw
ZniQwLohWjjFxyFjmksVNM3Cc+RdHS3bEByD2lXDmR6iLQbedbupIFvafhpj4PbQ
rPORwCK1zw6BgcZQJ4s5X/sbxOgSFvIJMSEhDZOEFuvVAKjo5BaJ7qe4Yuf6mA3C
Rzc80G4lOwS0kt6I7jFBaVHmJzswIymwmBYToQcI3LRc0vR6xr7BNoZ3+3KKK7h1
+8vEFFDoltBTwrj13U1fUPVC2t+bJGbnzzH57TFyn+CJ5NEfxRrtyBCZhd1vu6tw
vVm0V4IgfTTjsngQE3tEfr7elgLmAp5Rg7CHtoTu5HMkC60NhOMUgWbyE/wzPBwD
0bGuyUUeTA6SACxPOW0uvgM+0JdDj2dc9rIhAqzkIJLBcOO1iJNO8Ih0OAW4/+3q
ryeW6is1jN+7FEyuhLIIOOkKnLN/jQ9H/80aOLPNidNmTOS9lscVAhFYqwZlLEKy
TU+JRZKvfIPvDpt2XyewxivZKE7R1XrrxnlenZmkBphT3bddvh6QBG9RrSn8hFq4
v96ImhvzCTTZ4fieZ6IYXGgmYMfFVqoZip+3FmxmRCpM7rRMv30FI1m9MZy7peGj
La+cxupadNJxSizqGjKBexEVghYJbQ2gSx7PKdZVe7RR9twwjhSMowJ2tl3Pqzin
Njz8fV6bgymkK4CPj6Btbroo9nBf/Z0vfJ0hHiucnXFpJ/mfVil289NaYB5XLHOn
7um0g9SWCrNQlQhz8yXGK5V/rCAEnuZVgOg2FBdsu9fP48p8K34WhML70cI3ruQv
onUlLereSxkV4F3agyE6iXP8qaQizB9caGusNBxQt5cFKEruQ6ZWUWuQTWxC5c++
cwS3eJOt+aJOdOn45si7Ah+DFz9xIAxjnbL4z/n/AGN4fEAGp54rW6WrrGNqflO6
dKBRt7skxppJKqETVi2fLBlpbsp00/Pm6bhhLNbMiErNLvsm1dq60CNtZMuHy+zp
9AdG9A23vuAlSffI4yKm7wuUoKNxc4FilQ9wUBIW2T2wmqJ9JpPMhIOn+E78jrfo
zrFQbA0gK//Eol94kY2qtv3a/+zWAvN+qXnQWG8TxMA4VFEWaKKelqzq4j40S50s
eQ0qIUo5V3A2WcuGIMmSgqHsWXVqoEaLSQC/KdidrOgM8H2qWEDgcfRsLztKEJxc
y/kH+ucTtzON/2uQ2TPufEEv2gDOH4nbwC9VlN1QLdrVVv9Gt0lRxcNS7pkHjktQ
geW16Wnd54kvVZWSNY2ndZTOfx0p6fEDuV4i2EOJnTYWBomgyWDpjvC0GU3C6baL
noN+dFNqT4L0Sp+RISI8yHpG5BPCdx2f0kkuTI6SyUi9vFaQ9zKMSnn8sZMMdjId
TTbB6JdQ24odPqv8wmGCtPt8eTk8kCgQRe27Gkdu8XslZKQ9EtrVXy3iNaTzEZ4c
HtsN4H5kwa8vk2NA6hdepaTitu0BYi44yT8Yyx5jGBfYVQw811zD6BovKxfQvJJv
2S7MQ6pKI4oXWiR13zyNWINNj91U0bi54qOeP0WtxNQqJ8poFtCOSP7vmlW+Mfho
rtF9hjpBFEinEDxdAV91mKKRMEqLxsWEhYoUCou+5MMRB91fraasrVA5pcx9zyNX
++A1JiOQsK1KyUJjK44SqlEbDg17aWkMjQNs/1ySf5eTfSvwDZSqqVvd20EbG/fc
TdkKtj5bnJAWWRRdH2nexWkIWduPTonIYu91oKXYFk87ZgXFU60xymYnzP2DP3lm
HEvOPbWI0cNvv7/xhvA8TmKFXwXTM/2RbnlBVYxOGsLX5zevbwoU1J2b6pJwqy4t
rCLthXzIoFudzXf+sDo3EtIC3xnGctjjaCPambej804kCOW1B9ADK2wOhf/xfsci
6PZrd6FFBHQqCF33N22M3w61dYKQJpFPbxt3UwDMoSI20kSFyxSQoQ1XkdzhPL6+
Ekfs7ZMeaZ+5RRnbVJwgKDpe/L59W4CMAkdvs2QKgujLyCXUEzHX4YXnH55ZfTHI
Oaf609Nh65zw63iPDNLt9UogzTEd3rzhX+MCd/jvnhn+CZlWM6Pgy4i+45LVNV0v
VWRKXNmwWHK1AdC8eDlrq13AaIr7woakIFLmU3ahE9yOTLa93MsJjooDxL6VHL7y
V9EsI6DeC1Q94DImtACxs+C70vWR4zHe9HU/VuKwHXHaJo91VKxEGmWBwEaBr74N
84D+eG98NaVTfyrOqHdGXRZqCe8B9lEYmo6v+8jP7t/A8erfraJbwvANaApLfL1c
tWFzJ7V5M0yLm+ipBX5WbMI5vXERsyVCxPPk2Hw9bFJJqbKDBs7d12XUmJe/PTFY
OodlKLZPsZmxC+KNIVUvcy7EMdokrq5wD9x2UHO3gLHmDOAE53wf0vs1qiJrWTzc
J3OGEYMeNX4O6/qpIcVc7Vc1wM56lLfYmjef3yiqQP04Gkk6F/mwBAYydRFPldNm
0u8zT0SmBdptynrJxgpvs5qXnabQ4YC4l0r7S/ayZy2Hw8z7aCnTmHGa3jfPya7D
Rdc05YTSOI21Nyvbh0Zr1wdYLl1DF8/rfsQ4mAdHMF6Ciom3EYzeU8rO6pvDBVQl
N+e5W4dOJ4hEBT9CrcmjmROfW/HZnUBJI7wD3/gti2bbr8vI1222NWmFCYxRGJ+i
IRX9ZuGnqa4TAwhzAvIDPme41SwD8IOiqCKfSsZ8yIgNx28+nkqRyFTdNObKEsMS
OFtLCdbyDypZOhY7wmr3ZkOVnA5y1zN1j8wUgeEzz5hVfsYdKUf9PICjpgmtrjFT
K24vNAJBlSplSSlq7MLYcXq6lsJOyXZ98ugTT2r2qHaKT917jz/nTT//pBn68eoF
2dJuTZgoq+0vF3Q/zt6V1gsPOlXy6OT0C//LpUxVyEi4yEPUuSD9JCMWH0DZdPRM
VGJ85vdvNNJa9wWfcoH0MjhXuVXqdg0ALDnoHLqegKDIMSwTUgr+ErsuTCshuSdC
eJA/pIXY5g0XhYM47zGqjjkY7eYvpz4yDCEoT1K13BLwxPZOAg2tk51gO8DqA0xH
48toEPedkezxPrGpQ/wlZEyVXeb4N9eEkCO51FfiTzGvBooccEUmFrLVq1MCEKW5
Sn+pFJTjOuIQSG1qWqpb89NxMDIsYed0YMN/bRB4Qpdow3M25uHnJOaxDEdS1+MG
q1OUUCmy7btOvI2ZKWlH6U/gKDeyecDEu/oC9lP7TBvPDB4z6NX15qJy2QJiXKRy
yemBPjhZqo5PUrlZInD7UL1TdsD5RHrEzBgm0Xl3aQBKkVkyor0dregV5ikBeuRC
Rz6BGCciLByLNCsVmCE8/AP5rrNFpK7voOo/hVuf3KsCmBHJ9HDooIYxUXxgtq+t
Ry9cPgLmQQIs65x29fH4Xbp1QGx+a5mVbxEXjAQyHjeJjTVvD85ccg6xtarc//7n
9kOnC7VcqIs5auHRazCWwgZ3RiCzNiyaacNSoXzC3P07f8NOa/yvPziTK6hb83TN
0LqkGPmDk6/PLoVnlLsyPLf4ED62OeReLL0Pbu3/906xbVWL7yxBDyh1g5Bw6QkL
6D6zMdHhWlBoMneLgcI4kib/rCPFBvyAh199YlqsYdOufPiu7jQPAcDpjWIje59D
eEI41KOav6wct0bYtsRAm6UFuQRYYb94jVnb17NqNWG0alB6UiALYPGeymw9xQaT
saQcpUptEQMJ+H+J1lLhcIIwRVwNeHbclfs/ZHxBKFf7FWIhefLYr4LvL0M10Ti0
OMKHfAwVzXNwvSeyJ2PFxgfe28N0Kb32jR0I+S0kFuozY+flZg4KVlRF7xM5QXpu
LKaMCjif4Kfl9x8uemXMN4WFrgpDCQz+I6kxbSRb4W+Vlm5X6f5yB80DRQRa6PnO
1/ZxeL1grZTxY+lfY2XL1QIYfMhWIA4xV4li/uLvG2M/52PeLezNfAyFuvQut2Zm
hKOCLYU7Q+qRBkGCSTy23uajH8YFwGQphBWtwGOMtHI5t/WPz5ziCcFeJTrjOBXy
+CAlh1vY/wHvbWEuQQay28Fy5le7xRcoj5/Ke4SCI/4tFjCEoXJTKdCE9wtBitPa
jsSVkzLk/tqJSQ9ZgT01Bu9/gbA7Cb4Ox9bammDssDIxhMON2h/lBHisNJT2Vg/Y
gYqgvGo8x4CaRYHtW7ZXPL5sAFyr53HVUd1CQ68i6zGFPAhKx45P6CRCdYS/z5LS
1ujIrupMQEIcxQBaCgpNmaAQXV6b6wB5S6Gf1dM5yTLv8QCKlQm03aL0AuRJ5jQY
fPpZ4VateBJkCnAWzSo20XRIWmmh5xgzlJEa0ffkdWJHhBIrGOuIRLLvGhI0Li8F
9sXEgCHuL3SfCN7/6e2evZx5H1MiIGTuRdVT+/Q98mSYyVZHkwJQDxI5XuxSrY3P
9iG7gQMP2m0LuVmN0tFf4O1SvHaVfXDjOpV/atCHjDY9X/u/DSA2iDrzQmSJnS0j
yJlsIIQ2jRK0g8mHFy7MBdcHKsLVaI2ZG0kSfTp/jVpZoX/eekWGDYmObzzndIPZ
fiC6cyq1YbcTudNP3yVp++csiQud/U/s+/ij0/teihxd/QwIb9qFRBDi7U0wvmwZ
ZtOidEcWav3U4JwmIYEBvYWFAe4Z9xkqAgb8epkExV6om0FRJgRoYHuCd18CCM+i
knyoC4UPKVwa218zE3j+df+CqGLxuFdmZRatHVJA8yagNb1NLXBsrR60d97b9ISF
p3e+IAMKhfxpo6MNjE5tJGmQ1bD54hhVVG4vwXlbe0Rs5G87avcrP7zS6LuZ3ckM
6a+TqYEwJYtOLlFahn4O+XPfrYWBvQuEJnM2SvTUrGM2Gt5Gq9kfdQXZ+SkufLoh
nrczFwFnVnP/PGDmNUuvx1z/0ahpSjWPRgfXr2KHwGzYhSrBgjeEafwHrU0Gf+nD
whS/9jhQ9kEr0atq6nvc4hZGnjypVZZpmrUv5mkOAEkIOF/faUkkjJbIwftpncoj
Xf8OQ161s7B4OzqSCuTEnXxYv3buZzULhWVD2u0cbh0jcQIzHhV5vtGjXiFN2Uwy
nEzo4qAs7nC/Ys/sCLp6FsIiNLjKwCy98h9CCV4A27PoNiIOddfoslkyrhYNvszO
otsM5fKBZKnpcdL6SoRc/avIFIu8whGZxIIg+TsKJtnYy3gzVJW1AD1VosRzcuHh
lE4To+WT91KFRaOgKhX1KpjBUnf9IL7PnYWq9rmUKILxudPGKpO7y8D7Fz+cgv3c
3A9+t5+BSppSC0a4t1Sc/i4v/Vig/ouykwptssdukf3McyjOvbUxXnZUNsWwE3QW
zmynicHyWYYlRYMyWINtH7a7SvejWZZHTZ941WOvv67gpwchWRh9xSy+uhbeRHS9
t4ZtOzTAWvXWhYjKuZIhRRXobtyX6335jLAXsovfTfFAcyNbpkLgREA10f1EBIx8
B1kNfF8f8BOsphfUvF+jZZ3pGmjbAAY9rXakoEHA7/mpuTFRYcPwkXs2n6eja36v
2kn7tjqotGbS8kGnVXc9d3OHUjcZa10jaLSBLVsqICqQC4AwU2rzjEuVfUcO0GeQ
T3S0uVaN+ZqP73cHKQxjIyn8UKiiDdMfAdHpHuE0aIDE0Shk1VWDZg8omEyQUm3l
kPlbwcvwev/SNzSjlAfcAA+NJrol1uNg6AvvzfRXeY86i3xZDu7WiJJdIhYDGcy6
qQu3nbq8NVFzkojWIrwAl2NYWP1o3uVPdpsCiT5Wy92Dz0WsQhZM4NzLVJLD5cCK
uPRZR5fbHeQ/oCojINPXeyn8L+Tz5flL8R0BMtRxB+MltJumltqRRjXx+pAV/NVw
qArFVJBVzfksLOnxEPDmB9vMlvCOXPd+lMWB+kBOYBEEvkmyAHhYG/Rz8zJ9hlfP
hysxgROgnTAZZUK0qCDqo2l8FOw7xx9c1uwLLFgEEXgQP7Z/fvhJJDuypZK/azVG
lvENh1tC+vuO4pmGS5uZPY2NgM2hM2rudzmJcngZzXi1i9/LfoxK5QfLlCVEY+hA
dQ36iQu0NU6Vx22U/rZ25M8KGn8OuZfW/6lBRySCtyhOhFoUf/iSIJiItpJAChnA
XOs0wRdnorlU0968B1s/7UL/L2q+SOJxPavngUA2n6WEoyoisp40/KrzaTEhQklI
vKwhJbpkcUeOIwPsQZY+wUEH2wPoKQgQ0hyTZFsy4NFPjatj3Rh/lilNc/p6NHal
3MPayPUjju7KldV9LMRAfVcoKUBAQMrUWndIZpEZaZTVq/QiPRWmYtqGqZiRoC7D
iJ7BngrLPjxeY8GDw1vMuL8NC2B9sU7mTgnaejzk+qtAmUrktqrON5cHwuN2pim7
GDMGr+qmqRTT5owMyPS4R9VN+oF+iWNb3ROQSZbrqAZ59qhG85ZppTZbOBPAC0t4
JsgM2Er9V7PE2vTRvlqDPYepb4keTlirKK5k6JstQyUBbPOLcMb3oC0WHbsSyk9Q
sxcyZY5iHNGqaj65hkPAvY7G0r583mkhmCnkQDwg+Jl6CijXh4RdnSWc6w3cOZto
8TOtRC00a0WMgpwTZHrIuBeuzBdbZR6s6MYNYWNnpn7REy8wlQssfKAkDkJykdk2
csq3EmyShzf4yevvIcYCBYAlr7P+ValG/DVqdQaOdzsCZUJsVqu23dhmA642i1Aj
LmLvU0qvBndB+hnDEFQl7sz4+TNm1MbEVjEAFvKI8vo8sCBgWVMKEG4EmZ14H9dI
vzHh9O1jwXceG+7VJcXg8vvDc9Oj52dayDiVk/PN+u94MonENfXMuiAsDoss6nhM
+09t+APe790lzPSR3ujEsWc+mSH1QSZmeROgEMP/fQv5ONbZCqvFjyNJDUmEHSkv
+syElLLLAuuyE7h2EcrRJ3bFZA2tIWyweKxvelLBMmQz8dpvegGGjsO9gAtSBRjV
9nICdy+/UtZaFWBGYnFwYIFouQAvteNw/szixsdOOSbZTmdxqNycyeT5amahH8qJ
JTTcEcxQg22vVueZlYJu2nNj99+Km2G9wZ2uyA46/bQwkc26U9uZVTlDA0RFYEHf
QnP/3OEqpkB+gY6V43qKP41Lm2hLmJhwJfh2+l/+dYELw+PFDDek+yoxozHEgxIv
arCbcrfwjAbvqrlfGC/DltZNz+zjKddnYtU2K1w4qtBNU1gHMJiq9XdMIZeRFMyX
ikhR0PaNVc/9XGQPceHNiJecoz07njQ/AIld7I7X2Qc47JP83p79WrjD35cfGVYh
zWW1niB/GfOOvrnSEJom7Xe2NaBoDWwgzzuSDPuLoVsk07bleQ6SGrfgqHqAA6/I
jQPUcNCqM6b+WS8NUY3Ur2ReKFbWDHA54GtrUtYpCKJwfcnPOKMMAyrp13D0m40F
/6wSfaicOCqk119q1DBRKi23OBa+nfM2Nu0bVt0ssLqmWLVq9WTks1uMVz6GhHj/
SjMmI/vpYVXBIlvuxTHsTsppM91k+U5TPSg7X2Uv8MScvUs8ZdvCktuWMqg5OqB0
KFdu+X7Nl1QecJ9iTcVfw76iVcwkWcShcaiO8R2UYo1OoQSX6h7c1jv4qLr9N35e
c1SWAkUp5KJCj8rBiEF3PePQnJkkGrfa3Yw201hbjuKRcGIzXVAEI+xyPhlb5NUJ
ectImEocWVk5ivM5Wa7iJXeuvjifwZWNXca61nXdZIRWOSiwQAnfpqUTA8aEE5Zl
lDcWgJfP4BBsqXGx8TqEFdZYm4PtquK1Mjq4+sEH5WyqJsrH9mPPZwiuPvfTGK1K
fhQWhSwDoqREjhQvQvYPgcjQFeZL/76/8+ydJIJ3DsPV/qL29R4hS8W8BvHRwY1K
J+qmXokOKMQ3snaZXC/utwA3fer25FBTwtVClAtkkj4cktqVmqljAYvyzkUaQh33
ewvfO8C2Ycn92wIjKaumD2+plkPA01T67SdHq++e4I0GqHCJiY3lt76fWnVBkEhe
AuaZ1B1FUWbACMpIgUdoYE/rOmGzRK89QqxsRRYIxuJeGf+rOQWItRPR3qoF4dHp
ZUFYGOd3lWCK/QiE5o5r2kPlUzmAwTn4sqIMoPmDhaGurAAICocpmJt3qc3K988Q
LExjqDDGnay+KlpifOaM9Gaep3xoF/z4v3LoVRkUOV3MdnNoYyujWoMnwkQjxOGp
oPLfIvghrKVqLR/74lpb78vqxRoBRlwQQTakPDOoWB3jZCb1JR+XuxDbV5sTOxFY
QRxwbOgBonFuusG/Bawn7jF3NB9MFz0P5Hz7N0Phjt97PLQDCnf+QlMqyu7HCBws
HHH9Cm97E23UktxsfmlHY2Zs5Lw5Whi09zLolroShOdPqYr414bNxoUEIcVSmq4s
UcbaBGAu/JmoTEETO4q6o3SKs7o8f116DxXIHyT/HVGXOTOmky4fB4KZcQoVFqkf
FuQ8aV8mnkhdPjhb/pEkj0ZQJ9+jTN2EcFE76HZOiCyK8oyg2FaL6fJl17/WpGQo
5VFcr1OnynusC3OBXWYndHErqu0xP/DGgq7FjbHjFVRX+92T1pikfBDvm7nv0xQC
hdAQubu/zvQsDn8V3S6Hlg5bZZB62PAYehmRpR/6COLQb5Zf6Sf2reeNcF7L7Oab
nWea7ueIPP3naN7rjCA3v2d1Onb7zjGo22hxpDDgGTvenZqqH7g+w14dA9UI3Yt/
PhZsH/NRyq/zZyjdzcjqk4li5NORNZnXqD79/kotOziFSKvohs7fQpDJYl3E+70/
Z2isyBRJhv7vUHv3GNkgl7sMlqVY1ZHEh7KDqzJhZsOuOkoe1c0rVC3LUSTZri/F
YB9W4lFDQ0bFMCFjQIsRxAn76G3gBYBpbfaH3MC8x2GEq5Lxcd++0U/5kLm8lz+X
NukB4WR5zEg0lFIZV9cnyfKKhpgru08KieZp8I6ir0pC55tI7MDtW8ltBkj8uZYc
EAUtHy3Wzdnmxdsb5yuYGxpUBNMfY7vlMQKXJnBxpfaEw75wXlcyYHhCAJ8eaazn
ml4io/b2f0dFeTGX2l+SFSl9dhMZtsPkZ/W0nXO36cGzgEMTL/CsHxu9CxdIvZFL
0RrVFXugH7FdTQmlFQME9j3sLBJldhhXxFel4IFXXNr+0mLMZesBNkhO7JCotudW
87j745fn00sDYo7gJqSo7iyVZ+ESKbxpHY3LWsy83dD4Ca35UuT1R/wCpwhxhs0Q
ypOwvJ6RiDJ+7crvi3250rHH8MJb5+IeELG3YLtDkL3xrQW4dpLFTs/uyNQWZy1C
o9CE53aDjLcJQhWfdKEvRkh6GzjfcIZNL3Yy9ftt9p5rN+vSvWFG/19nyCa+4Pv3
xiVidYas3O1UfFmDdOC6/36fDYsHgyrbOVf/q79ZhAlX3oG3FC4NJDZ1ClDTU8ho
N44gSYdmTnvJ88ty6w9uUburMgdG0ancWeMFReUsdbjHVGsWcCpe9U4vFb26yvaA
tBJ4dG3en8aWrD0i5UwgJ+tTPv08GaF8BzJAQsNeRvUxjINptqIdnpfokuCG0Wi6
MKJifkRx7d4tBSgXdIGRvKGXr9rogRq0u6dDlsh3SL7ktyItlpDZjyeo5IdeyPjj
+sPSnalp58h+p0BR0zO5x6aRDDW/Jgm7xBM305+tWB/9UaVfsH5fmkfTvH7BYn47
MoGFwhYQLGcWIBkU0Pd7bvTPPfYDhF6FqyVfjKw4Uzb7ai23IfinZ5JCIMAs38of
cEBBARusylyd+DxDJLqmOTsxAwCFp6hnhyDckZv2MXwQpjxPtosiltQY1+mb6M79
lxD1zMumYZrfQ9KK8A6UnE5IrAo5aQYeki18NIM7Go8zfPZST9AhRXhX/uREOXQY
ULuCz8UGTMUefc+322IvDuaFH/3MkDVQNeh84RFWJXbTShgZjzaXOS8Qmzt/Tk0E
fXsTFPbOPOmvr0Q0AtbYgWsERsPHXDynOGc9R7fcChNcTLqVDC4DLrA2WfhF0ro0
9lgd+EVB2saFn7ylUVVkgtA8FT3B9LHwlIguHSv1uJgK3lT0cLhQEYxyVFMMjNLS
nqaf7vGZFyKYFqC/JE5wvhhynYyqEDZ1I3LmqgmdmvVcIngTSRDIKDmA3Sm4qMWr
ez7eK7+JFui7EMmDncCJw1HcKDfbRs4lljgOG4I2XI9uZS+HCoRIfsE3VnrLLTD3
4snrkE57sZPG7jDMOS8IDSWTfJapWgTuMv693YSzhdmMhzoOYwHUP5j+Ka3S9Yj4
ThavrspMr0NubxAUxfTSuInLhy65mEtlU0bwxD53sQCBIB+fT+0off/uzKh582kv
ngdJ9X7iYK8In+7+pN+FfbN01myqlUjpzZDhBuTcrRD5RCloSIPnqHXtCEwPE6yj
BQXPiFrcYBA3YsjL+7XQfV2i9GjjGl6hMDuY29kC04SRTgMb7PRL8E0hRHLGDYMv
aO2VyEQ5t0bpPL4p3BMKnfKfpijnLSglXB4xNBVUTpvjPIg4ezToWpFt9CEnXiLz
FrYLIx2E92X75v0A5beP6FyQ0VOeFvZQt71ry4SUr2HKeSt7gkv+iIe3FZfdx8+6
C2g0kSjK36kWeAz6QH6qAfqqNYIUTSl8EC3ZXv0NqS3+SzHs94pCYfunVDnG/K7v
BaXohtFIbcczTSjIOUhSvWLZC6SGwR28qKmv+DQvS/NvBucGPNkcZ9e2dkBh1aJ5
qdrKENc8XMnRpHMJrOzo18rwuYvc9ToOfqhMKqDQnAJEDOUbuHRJ0HfXnA7QdWt4
VLaO+PdZvlHBoeYvvEPBrzD7W7EYsNywlKz0mMch+/dnw6IkHBcrPfoQVVDHAnCQ
k6YhDHKWIEf2ed0U5WgSCUMr2VrDQ+ze7jw85jFJysE9ojIVbIp25W0oCT1zm1Xc
5Q9Z4NYiymuJGjbE4kbbA9TsP86AKrFd7Fd342TEnrZGMxBdnDOCVdKRR8PMxBtx
04EP0j6ctQlvzR81qqq6r4QnKPYcvz5PSFoDR9wcrtt0myYj5fnfbsKYL0OBlJlh
H2hVtCZA5UcEvqyfCPATBB8qoNtWCFeXuj256Qpvs0/apAsfkW79w1boU0HjUBDU
IoVrgGxapantaQsI0DjcTYhYohNctyPwaziGA4U4HWGNb/TwE9W5LrQegu5/oV1J
6rVdESahoXox/Egy1LS9B7MNTw0IrkTPCxVog5D99z1xEjJj8jjpJpDfvsE+nI9p
ORJvqotXFuQEvYaXCWflD2e5npOqg/6azYheGfJyX1xHuDueHMoC77ZW+8cvtkqk
KXgmcTwFnuSlEAqe6QUG40V62g/SVZ1zokanAdLuYvHtbweO84t5NkkMdHKvy512
11nDm0UOmJsy3EwvhNZgibnAyzE028ib+jKIcC5uP7q1yejGlG3Yw2liDf2ScOLC
F48Xlt5+j0Pamk/qs+9cBGGX3x0TYHPOmIUynK6tp/JY/S9aHRTU9bijs22GWWne
UVcY+BAlBEaRX8nhPqgj167drNU0snW7qyZHdwHT+rF9hWvXoRVc3sh7LHx4sXXp
fAppQJsi1X+rb77gCaxtRAf8BucC1VZZwjYmCcnpgvcZZuPmc49mpNXy+JY215Cp
ZPbqkCmXE9rHvOURxbwK+eqCljwUOBJ/63wXtRVd3IVKlLI6w1QqAzsp7awiBhWm
m+6E9KRhjxZRRZ5NOHIKzfkR9uLZlv4/XemFqJ/x1SmIfq4rp76SD78d1Cv9yDKr
3qWXTEDzz/l1Vkk2FSRYWCNHDJzKmCbCCRap69Uc8ZIVThy1q33aAU4bb7JSlHvC
T1k3re4YK5WurwqNk/y75JWId8ShS8Dh0m6ewV1zZvxk2jSowyHaUSTK/HS1OxU3
qcbmNyZ2Qzyk7nNpZOJKhV0/35zQu0uebnyOJOc/mGLpPewnN0OvUPWbmsaEILjN
N8bKvJgTiCQjwXeS2wdzz3BApiumwqT8HOTQnZaDbF5ScCkUY6JncAxPMcgVAQK9
xYUloSW3UX5m9HLjSrzoZuuCejcdWcczIOpbjVsLJH8vd6r1BzzncS1pGfJBqseW
sMgRh2xRLZl23ma81u2/xR78VYn1x2gHrwicEVBn60NHQ0AK5XhFfGKAQe93ZGpQ
ljJ/4lDTuhYTm5/b87cJCgNae+32w2caNqABv4xSxxcU2V2nnT2/7OCvVmEjOp2D
UZQtdSfJg28EWuBNVMA81OADUtLbGgfmt2n6T6+SqvjJdJrO5ESQHsndEmXwDa3q
Ttss1r6634qHdVTteuvhStN7hdpTHr9+FZZtC5oPUhBmVXDCqvqhU2WCfRNMakcT
C1WalP4FPXto62eSJdPAZ/mjCBo6vrVuAvbfaxfcdNTKPYdrSTllzcvYWwEsf5Lj
/FqlH30ZmvqP2ML3kOOI/83xL0LSeqCIWpd7b7SJmO2Hp0PH1lCL/Y/96tJ/ycjp
0jaogUPGDKmHsscxO98YTmKM5ExTdAulpgANC0sBeJUHap3LDKFoxqESZMcQVsHa
BCzKOrMeLtGm/jZCsvT1SXG8fj7lHtcpl5ILP/jGsRlq82QRwCNFSlQFzbGUM7bx
8RRXz98EDdN8lsAJp0Hc+Gi4CNhIAgFKchJ5Mc1qlfo0J7kytYOY6IGWHB6Km9vL
vCTs1y0Vypq3BwUaBUSxjBxuddK0r9qDHZc8U+4oZnMJ1Hj3BtKPNKweaTxC35vR
Dle7svSJFw5xNiC3IRdGQHMiVKIA1VOsfDZhzMhzWaBkgtBvwymTN9yIgAvk2gSJ
9X4pucjAzW+ZcisW1HUUM5xU0bF2uvlhWL3nS0eal2tXRAJldzScRaFH3fQRMQOf
xsw3wLebJQB7hYIGmjbzMG8GDWo1m4Q65S+YR/yc3FxOkbOPFnCd6DyjTOh+AyyJ
vmtmPJPPs/E1VzS26ehSDNhU9igVbkJnvvtjGw/VaTFlO8ewpXDr9ahTdiTs5lsf
YBDK620LOioDBQNzH7JJ6bETS5/k7KaxRfJ7RdIhwCjGvdxPuiaIQLIEbI0LTvgT
AzuAdWIOUdhJ7AYZA/eZGIl4w5zhcXBznIgVU/cLnhUfeiv8MSSuBC7dS5gCmdUY
GdfBJ6lQTRS6sB36ulcOrLDuclPu2iYlgN9xR6clsA3cFYgSe2Hn6uoLLHQXil9H
QxMD0sq1kt6EYAWaT3gjX6phue/gMb7dcZEHsU5BtGTRhA7OvlJU62HJXYuK5Rek
oJ+qdUf3HiL3eAMF6HQNBE9IqUYIGG62rBA5DZinDr/eeH85sy+giGUzJSBEBKSA
Jj6/R/TFGd+Pi6T29DtXGraCgn+AJFYX0HQzpIks+3P66K2YYUzcje+HG6jC35Yk
4+GKbAbh7hgvFjFJRgKLqfKYz/5t3NXkyZIcpAcbkJDZHUqi8bXrFHHDUPE5FXCN
WVZiOHX280cupWqw+yjQnLbzVYc6UycdWHVlHab33UBKTP9bKt3eibRpcj4dDKxs
f1pJXexFifi+jlecCw8d8okxOtcTMpH5JKySGef6gjkw3Vlw0p6l/fKotjnKDZ3D
YSDeLk9IR+A5+6comWjXDXnfWNk+dPUSm5zHuyGHFwPjHc0nMIY4HTjjR758DCU0
kJdJxAnRSeNXFCl0PLzAwpErDD/lr8FREC6a1zNVJ+EXq7toRrO88J+mH4TJnPXh
ehdKGIuRNmJ2G1hZ8sKHL/IyHB9tcKtZlZ5S9zzKJVqB2QYAXeNkvvP6XpBZkk11
mSbmCaT9/eaJ7ZxCX3+rlIGZdKyO5fZrz3e2PmZaOZZa0r1iac6Vi5cFG+su6qEV
6UzFjEV6fKc/mSfjK/m7rxxYn/U0McV4sxlOXBWrLhLTlKVRJ/o0TlnUIFRAs+XD
MqfsmiC0olAsGnyNjHUNq7KolrcodSbN0RcJeLuIN7yLEOITKzetZY0BA40tVkAA
nXgr66Y3Bc0C3OPx6EGhR3H7wOWaf0V8qxkY654sJL5wz1G0eTWEkwA0mZcQ/sKo
SnZ0nikNeJNY5QHhKeipUtpxcwd19G3EPaIL9Qw+redf9XSrfNMEehxg9NnDyhPF
KlbIIzDK9DteaMmgVwlb28jdM6j3uoZDbhzOrzpe6sRPpypA5OW3A3JPvzBM9gLY
GnhGF9/rRzeIgpWRaoRBeTjutTUNBHZlvzY7ELk0IKOxxpyXm/8UGHpvfYgmv9fR
ORC4rE+LZNbFBu4QAXEGlXhpeB6RtMjrfAorsMdUAAEKAWuBG0wlWTqzSzv0E/Qc
eT97zFEqgsYewglYvJs6tAOkmJCTrJlgxLEoKcBCMm+mDguO2OnJQmkCAeeax8gC
ku+8LQskoPwDs2l3rheV1Z7bwdZkLbnegp8+0qBkYC5wrjyFNrjsZrna4CBnv9J7
xfmZ/VHISNBn5FAhjBv/5M6XsigYZIKbvSwCEkzKcCikC7K7SbQiQzoGQKeBFQTt
eadHVjvN9OM3KCnjgjOdUy1FaZUdVFVVJXZzAKR7akX8lyq2U/xwMK354+OkAKoZ
PLUN/bnBMKogfIwqBJMiR1h7oGswbV8rJfyYixHf1YvvDix3ng4fftkMa6EoYxz7
sqtx/HXSnIvut9AuqleBHv6iOcg6HA8j/kPJwspDDaiu4A9lKEFwjr7I52lR5Uk/
94OpxjVhY23yThwZIw4pQ7nNW8fmKsBlDsetEwaTJfH6803e4wzw/wE2qb2qiQD8
MbrvmnyvGCJn+IOtKIjE/ea1zcSVBfR4FRzJ4HTlwSDrw2PASfVUBHVybDNcheMW
hxLR/4ve1i+uRDyvneTTHw/TLM9IRshgHJI/97diaBICvRV4Sf6xSO6Q8a4WqtCu
QqZ2o89yWVMpVqbSqm/e+B6/8UIGLNacoc1IzEhCvRLAbNXFzg+ZhIda1ISfecXC
xATLgy2HRSBfXdjvTGgY6lc+N7YOtHZhwpYsyypNXznGK4N699WaWhk4GAQd9RNq
VT/MrIJklH0G54g1o4g2Q6K9I+mtamuO+hWLp1fR5/4Pc30SsViAu+lieRTLVE6p
1rcW4l0BExRqyYBd0LSZQJEK+NmKL4J2vW1HpBo/Mj45WeUJ6ZDTMorgdRoja49A
G5nrhGhgDLhqUgExaSV7x8KqF1Wyu3H8TP7wSOZL/4EpePymoKaHuopjQBO3QY8U
2L1Gnq5KPfMOuzs8ytLw6MT5oL4dk4N5+FK7DxLF0AEar5v3qAoe13hWUqxswgEm
eMYz0rTci8WnXCIynqQB6VEugvmnZwTnAkQrFrafo1//ViKMZwhg6BcYN16o97NN
p8+qT+iWh4W05AJD/myKNm3HjWES+/wOAqL6KwUc7QdSey9bQQIHKo6J5rO/Yerk
1jVD/0kQR+4HTl/ng4sSF2PsPMyCmVxaGQfyWOvaysnLAtL7FyP8L0StMqBsvBiI
7dK/DDdVMZ6j2HloNNvTbViZTd2PTz8dbgTvZTVusG4EV0qa6amWGiIlfsb4EFKz
ouQdiAclDxg674SmTcVtoMlXBjFbSULwJhoIf/P77bFbPpxlIfp4vly+FH+CtTNo
WwXDvWOaMs8hm5tC9aVoIxM5ua60tQeYiBTbtKmeOJvs5lVCDjBS3zRSiew6WyQK
uywAkY3v5r8wG6NeJRdaFw0wfk5ZzCGvSVxfVhVVWcN1xCVEXiXqhFNIm/bQS8qw
7TsaiicnOq0ODx7/CQl+tltax6PJNRR/U8ZqD66GtlNxf8/EzWGCxWWus5srJXf4
jA8jSrjeorLdn8txcTh+oyKn/UvSoyYs8CUEylhiHwQ4pW/fFvE6y/tKshxGIH7Y
W75g+0ulj4+Khx1ft2HTiM6OjPGnU3xtBhWeXBDSRri2AG/YpVHNKoFAhMlhYfki
xHCIVEpdq5AT+5/kfiZxUiWwTvc67lzLnOCKvpYwnsyloEd53KjDS+pU8WWi83Mi
9Farsio0+ozYpcSDZ380rhpjD2URqohALvTwTrgTWWAb2RukDbNZJeI6A2iXn9tu
380zrAzDIR7LOlCArQj7XcoGNvTxacDI+9lie/B/xxRIAbgLHLYWkPoCxJmXNelf
DDA+1cCOXVXUbPoMiWspE1NXiafKocpyaEW3C0JEG5/IUntzcf0GlyKqLTokeCam
NxPVDbmRoD2TQ2cmyet+C1VMnbYB+0X8qAe5qB3ldF2F15L4T+JDCF8ULAzBxD/a
dGqJ9MSNXa8f4ZOlIAlkCeB/ScbLDC3cQ0fqiRWhTwU5KNhoUEtkKq+xkoyrVGLP
E9N/0XSDxUnM2bi/l1hSv6phHc94uWrCloOXrIa0vd11KgOpPXY44mvfN5sYxQVm
vUkFiqdk+yO2vi/q66ziBL7PQgYeUJKFpfpYdYYhziSv9y5A23Hu+UXL2VmP9hEG
euxcUW/P2eUazKbOEdzTM6O73N+SXLXW/pLjtz60yKqczj1fBw4J6Y0d1DRd6Xvy
z73pRgV9eVVlC5EKF8ZbBuQoC2tm6EBkRfdPxEv3SXaNkTF40aPMgGmN9prkrBYM
MXs7K/jqFl5OyhHgLbqHl23SntGo+nEKniChE2U9OBsexHO27iFIrfyfapw/S3W5
OG9MBPkkRZNiefXY34zzN30pnkcLtp1JE/SIwocnot4RtijyL7S4myfTK5XKgKT5
XnHg0AHaw8Qi/GkfNooF17CFscr1wYpwcWs0gADHhH8E1Hd5A21JovCYusnRp4cA
20Bx1fVQmpwic9ITecn9RHeYemcThzmEj907T0ikF1H8BgRovk2TRAsVtZ2F02ii
zv8RGt0MyJBZGOmpNmbqvLWrT5WnB2Mgiuzh1jt3tvHKMHO9P3Q46ASuWLT9F/rh
gZkGjhdJPETBlBJaLOvRKOk8sYR9P81It4htIz1s+mWI+Y6hqmp0cssKnD5p247y
oU2Wz/qba5Yv5hqEyGUBbkYiOcoutc0d6AKVWnQDH5enonxD5BDla94tqYkpT/w5
Zbm6I0ATQ7ZEZVwgAn/WpFzA+od3QwZ+A22YJ+13CEvSgeOSADuz6PqcMbQrZk0Q
Rl0gJmEJSeoSNPl+p3Ne6hQoCuZ5smYZImntD8DteUHx4n8ivZYMsEQEdWsyg4cN
hIqH52qkQylMv/s+Pgk6C0oIPMUuSsaM1e2vjJ9PXu6oR1dq1Ubs99yzvwB3kR6T
X+iAO3U3xXu63bRxJ7dPD2NQ3LArKfRe1AhY1pykVgCRvS0KCRieFWNJUILX3gVp
ihfj5x/HEtHfAlgXQCixrzIrxWFdSPqT2PJ3mLL/PKHHxqSvy99asEvRM5RIc643
7Y60LHpqH58QvHMCrUPwEmlRdzUzQ//h+FNAPYzMM2AnGw1rIPpooQeac/MUvNAP
ERhJE+iRMuS27OfIEi6MVJK0QtjlkHG4RvchBFqTG2tsjsbVtrWXhFeqRZ7zoqXA
jbGosTUuTiZCT+5EqYiUEzlD0r1vIagqiZaRzv5mENBv5X4IRv/EJ3kEZKFMy2/z
BIj6dPUl2M4w+df/mLOKTYRtDNw/z3h4ZBfhhX6XlcygC8LK1K2Z5rBwoaA/Ep/Z
ONChYQDqjQRpgjXHI8YIaYlYEk84AoUgHCeZa+FKYGQ1o7q2LG3+vH9RaEgxmiYO
osAwn+at2QPO+OYBWONLn56IzynQf9DBoa5K0HdA8ji00WekrHsoPEK0IGFm3cuK
lYoLCm51Iw3qq/vODfrO0vvq9QQ0E1P+gOyz5Ntre3VF08cmMPFsyFJXdr6KiGqT
bvmSB+6tN8IYS5e86NHDHHm7i12GQ2cT5jpdSOSKCp+LEmY2a3iMaFy5tQiHwgff
47L1f22U6voU7/4JsUXeN5Ak/7tS2PH/RIlV+0P11dI3r+rWdDHq7GHV8YVOfHGu
HoDIY6KS8RlVzihvDjxBx9nZvNReoj9sNG5Huxk0kDTULhImbGyVivY/ZhhkSYBq
eE3PdMJFht39QDILJYNsUw+WS7XQ2+WQ/5wkdHDuKuANeNjOy9luOz5CXA1gdpUb
vk7cCd9nZ9XsK+kMbQI9eWcZCrPdiyOttqppmkoLjgpYyaUkNZYOJme/jEi6ED1h
RtZhyiYi/qVQo6dB5vfKOZjSBcFMjbtF/wt9+Fy2efYyu0/k3ZDUBK+LF4R/5siB
h5RCtD51heLKWX+4qjbN9QPkn1f8dTXtg0m6nSp6Eppw/lSlTOLb3ftMVNUEBRsB
pxxvf+lKw706luXYx5ffNs/1G+PprlcosZmlNHSjB8PIy9QMTV1KHgHhWA53i193
t4I9URIoozaN2zcVKZ8Py3Edr6fARQW4xmoc+bY3Lfmzqco5fYcaxav5lACHGRmG
l6KUgkbwVex5UMBQbkUQ8ct/9Zu6fnoKLDAM85sF5LfvKhdxIyKpVtqMQFaL6Jop
sVOC7ktUnrOuJnXb6e8sPmOgHurieHuISnRB4uuMPKdd83WC0/Svh6R9PYnoUWMN
8VCZvtR4NXpQM0eTdlPCChul624q4Wx7d0ZTcC+NK07/T8a/ZC3MqmtsBdmYV0fF
WErbZmfZqeP06Gp1jffPz125qKT5k8O+YIUmkh93E+lkqU2RdVaVYVEKzjQTnH88
Q3cTJhG4Fb17K7sEds59ph7wHfUdaDc1WeOVwBF8+vADns0FXoKyCCKm6Xisph6l
HSCo3d0DekjVHZwvHyeTLwAZhi2v2TM5vIdwolJGjRTcQjJdsHrSdVPYwUFj1GIv
QqobSha2gbi5XOzuMTOLsJ1gxoA5YimoFWQCMnhNWjKICUH2YiOV1ZVevJpfoUEU
s9lHV2pAW/1e0oNWNj9wQzvEtyQpwKGPcP5h05G3y/oE7wj8cmIk8Kk2BFRZoi8k
QPXmgAZkH/LErSOXbd0YtE2yMmOHhaIlS/fIEJGuBebykk3Vh5XluIn6zJ3BY36Q
KPIfB9W1IFx9yKengwm3kmsdKwQlJooc7+4AnA0XqK7i9o0ffU7meC1Y+mAjRhBI
GZgji9H0nOB6BOSv0YySUyYllKK38ag2WQKUZeeFNQ60n/gFwvh8P5IhmcKBHZvt
yVJhxahQ7I7YW2ENTr7bovKhp2llDNJtQamkkfy8z3PmMgCqEGHrpQkVYQ4jFl6k
iM/Bd0dV3lLx5QFnw3IYx1etCqe7o/24cDbtjMGbrd0NJN3GTK2R7TuqkNSshovP
6MJc0yDeX26e38Tn1LQmAbRI8hnzgR74BHok/mPhYOZX4vEr9xCxjBp1Qvw2wTS2
CiGSQv+0t3aAZ6KzwHMS8MlRFRPoMxz2Nyn8RuzArW1OaXpRe6QETIwMc0cT/ywY
N93lH5B4289SjoaIY2fyA25u3DXq9VPitTkeSFnCa4stNs2tSJxyp+Voo0kO/F1M
IX3whIdCx70AmPsI6A8grPg024uLNeiSSdfaECKHXqznE56QuZhKlBeZirxbQGOp
VUDGzBPqzqY+XoNhHFOYfZmEKcqifhsLu16ZDGjzUcwjDrHFpG92moACYIbqaNrQ
F8dqIi+2KO262qp3G144FPojthGgT2xTnAyPy+vOrHa2wQJN0GxmDS7VKvJwqX/Z
wv7C/1+QkvfoP+rm6ccelaNAlxMTCBd6IExi3fY+OApuoLo0XvepBox14x3xhsdp
WzmF7IY3zKO9fLAId+xS1FBbQ/FCtqH7LM9k+tm4+pC9taIYh5xtgHj046NkCR0a
Chzmbx0G9YGtGJgNHysblOKl+DiemT+h/a2XHxPpNNnF8I3nINh/p528f4NnsgQ9
J0RilvS5FAlpHpNAaL/kMed83Oocbttf69VD3+bTgEmnCByve8VEePzFMSccxpUU
CwNzGuZ2g4uS6EbhkGt3SbAhQSvhaY55QFMOWmXVjfv1OzIEkxSJn9aUddPQpHnl
NzN0U7xvuc3si+SCUMuJSJo+DmCSICj6wjPfW0n8KsqIVfSUNMXQMAHrc1v9L9dU
W/GZi8SBdfmhDS3zqv1M4cZlC2lPzmUwo+4y9mNHUfBWBuF92jWekKoLyucLzxhL
NG0H51Gwie6LAuEyb7RnrTwuK9xnUliraW/XvXt1lX6sCdAd+BPhmzY4ZuCjNDC9
8NvwUz+cikiuESmQT3hSqUfTtcAzJMNPb/4XzswZsdS3Ux/L8DziuRyuAf1KeFuJ
GY0Oxk+hJLA6ReLOEwL+xBJlDGYxdG2oBxwm7DymJmoAnpu4dHU/3WJHO/sI+G2C
8osHUHgjhnN4r2q6FX7Xc+elhzUOM3lSBgG9/P0eI+G+pt3uhniaWqtrt7Yz7VbN
pf8x+AURKqekbKf22Wsq+1sufVXGgigoXFYt22wB5w3OX1sfd5Nxdpseae1fJzNH
sjAodP3GZfSk1XuSc0B7LjAucl7f6KZv3asIjeMJDYhSSJkUqKqTvdHO1NiqL81W
+yKgQ0TQrQwkUUn4GGMMZPtKVX+VWdMr9fWzc0Buz8s3swsFyI0bk7uhDzIeHQjo
QpmL20Nyt46csQe4UcAVgMC8edzIHUz88ysnDcedaNuedFwiRSiII2JNOizvkj6a
8AtlZ+GQaa8ts5/WusjI10PpcKPgtnrGulQvzdsfyzyefZDfiJdgAK2KQer6FKrZ
YxIMB4n/2qpbyhElkqOpKnn/XFBWm42Yjf91/pMFeauZ0ozLbF4BoQ5+x1IlhS38
ogNtypykNaC+VbBx3ZqsPFStUZawircFjr6FRBD9pnAkNmDZpvTKKj6KqE88jJeX
WX/GbNu1RU7LkBw5jS4CMeMpdr2f6mv4no5ysQtYddQvamcDDiK7gbpgKYJypJtS
1U28NSmX7EIShDYmy5y387d30O3ZNxnmzL0fCknHVnKKYsfzZLomoMFr/sZtqTls
XRU+6yvYqJU+dEHAvfR49K+pCK0CIFyTF9K+ycnpqv1thsn+PkqBxGrHfM/qwUaL
hamWJB8UZ18ACvFferNeqGSNbHQeZkDGPwhqAXXW1i0Ot8r+ApEw4OKk0gNjMTYU
0kNRINUdGPHyP959ViaeAqkGWl0T+FB+csdqaQ4dhsxZygK82y/tmkrjwwauumyw
fqWwEG+YJwxU/giaLBPZw0t/VjfxrZHm2uROd21bhPvtqvLOEns9tbUPFlqRIi1u
yW/VeJ7f4ouGM3Suxr+0j4kRXuf+suQmNmc0s0TYi3+JMgBh1sbUwJMl0jOlQf7r
oaP+xl7ZTJQwhTKXCZaiVX6Nk7zWxAwr9RY4zTrrDA+astt2AJsNcPJtxrvYKNq6
xi4cLYwdOsCDeD7dQBsoLn1fX69RE2BvLx4/6yz2YxK1Z4q/40DqQEWPd7ZwEls9
35YjZoUHiaapxJTgr5n1lD2DySrQq/wptBIzpIVGZXnv6w1+60Vr52vWspalr/Dq
kXTFJFJ1A+CI/zt68V678xUimMcRMhNW4c8fsiveklf10LRsCKKeOXU6iLBUvzcT
4yYDX16CRqDWnoBs5rMYou5tWlzo6xp0j/Ce7j0VoJDAmcD5OioI8LVEerRv5cub
E1iuSX36mqgO7pHhWGDeEtXGRl6NXwgWG0GcxZkpkESsz86/bF6JM5BRjpNs0AiA
mLWcKCzlVx87/jbL2goM+o6QiFEHgPBn9nfqVnQh24QFwmAvlvPBdbM5gpoSZXCG
+bJqybPT8ZJVzQDZ51CCTLXf4iQxqbFP0BhTo7cqs0HA7FXd21WjxDtUDddbeLpk
PlEvVDnH1/mB4+S2WdqlsMfGWjEQR8+hxbkt2aFG47LCqhehF+a2Vy+qJwwaMplk
aIjov/Ojp3xPOvuzc21cNRRwjc02PTSwbcFoO7qRrGfi+TW4rk5rME2WqIm6gsUH
M6tm2a/wmBcK4f3R10AhJqIGaRY3Qb83ujVHDt0lfHJIu729B4soWmmU597vHdFV
cPEDHeAHN7L9L2aXJHNpCajQ4nhi5jW5eo5lx1V8ruIDyj3u0eiT3k5xw5qiryBD
QMBmFOp7HZib3BkptDQDIJ9XiPc5hws373nMhH40v+wUGCpkYPGR5Z0XpK/Smy4n
5txp9JyWePf1OsYj8c/okO6gC/3jgz4ZWq8Kx4B5wPjp2cfEjpDN4pwZrUmdE2Kg
xA+ZXPHztBciyWVoEgPxiO9DHRa4mR0RM4QeqIdqUxEIdgdfVILfSmM8PsvT4bAc
AjOdgCXnpsl/rzsxO53IN4oWT2+z+ADH0569RLIND97kV1CAGyh9qincQPhx4nCu
cOdz8FQ/j5UBoR4RL19FrOFj8OkdS88jCQ9S+zS2z6ZLugAup3KPKC4yoDVi3wqi
135iPYEeEgb9rN7/ZHFLMAVZIrjMwdRrVsKh95+oZnPH8+jtduh/WqrJ3gPPncFk
UNAJs5eh0yhZrfd7G8jgevdtu9luVP6ZLf6Wi1fG6KlZAC8mx9Vz7H8egD2VVfQx
8JG/5boAr4nd/e7e0OBU5Zh5BddVt4whsE5E1tot0OjiAl+8evzfnFM8vs8vDjNZ
3CndK3d/6a7y8bxMsPM+uzH0UAs5apv+DlofmVZOdx2EoXXl2YKnspgKnEKoFROA
XLgTIwb4IavZth6mgXT/GriI45B3zbNR01NuflLzmiuqFfmiJ0AUV++IiNcF3wWo
86jj7W0RTI5Et+dicAgQGq+4DjhbWLkMA4Fz9p9Z5O2PwVGPATjLVO3Y3y5m73NW
yXoZfyxwHsNkvfWSZTch4K4hs069FTmy3+taUxxv1HkIJNLS753A6vBKtyiZyN70
Ms+8sgF+BaQVGRiNSBUD/qca4dx+7ixVFyH4K6/VW+oa+4+OvJw1beWc63SapA93
xtZR4l/204o+hqJXolpZo6gq7a93w8LCNIoah3VKeIXmzh3ngxmieQIS5AYFC6hc
IqE5fXZNKHZXo1QdJcfe+C0cpWmFjzWZEDpG3jU75DWwZhhAlxxRdhHmF2HgRIFl
fp/0qQC3Sr5u4u5afpBLVlcJR07u4AOuj4hXfZMY+fIGwrblDmnKxhcyYp2R7rap
u5gitcGprc52J/N5wUFT/Vw8MIflUKqlRmcNhbKTn45+eEXmSDJv4vZ1QNiN6HkK
v/8o/LHDaTHZnAHU1cubgPOpWfwiVXWGUn6wccJ/cbyGkaH6nWru2bAsbGTckyd4
Xfu2qQwygDvpByt0XTOAwM0xkcqNp0f+octWNhGfLPpGEqWDX4XlbLFmaqgGi65c
q3AgTtI7+yI60EohPmBefsfTjAtCdm0jv3jIpFclAi+P5MAUxtSSIMiWvaYsEKlZ
pYCFvKA9ang9QslmniR4rFPpt7duuFXo2h1EdZsRPM1Ay7P2w1X53AD36ghV+28S
IIeqJPjhnqjDKr9KhRArpr+6QWvXDm7Ms/Kn6NKNErUaoVZldJRV30NyVjHzzCDc
BECmynZm3Ozms/KXYwmJMlvRC5ONMvW4QSzqpLrTPPQytjTLVQf1OTfBhyBjmqS7
SZE18r6CzsaetWZPdZhCHHPt3mZGw1/AwvD69rYvU2e/sTCcrvZ//IMA2L1Q0zol
ng6YqvXBkv21dEqipDh5OK3gzsALHe3KVvU1b+/IQ4GwmMiJZQAo0Q28hC2Gqb38
YDGQawHdIBemNT6G4zmCrwyLx/XmFhwzzTin+oNv0XRQhQen+8MfQQbaC5IO9+VZ
VE+XnNSEy0jNwOrwUS4qjRcCyVcMwkcteonH/Gwvk65TlYxcGCo7rIF1b0kmg3uu
18jWdzDYkmPH4OyRG973973wI3SUzXnqW/YoVbuw/We+3GQM1eH1os4Y8+HQRedF
xaybLtaseWolFsvj/DFiukTPMi5smwtTfB8XaRASFSwfE3ZvJkhACU2qtluZcYkY
bUeGB5FDS8ouCph8x6qs+udJ8cM2K+iVJ4Y3lX43SfFWQ5oo8BwbPcpda6+gO1cU
0kx0qQ/QoPQ1fZjb17msatw633Zwkg8HoRf1xurobSneOvyWjGebR4Qb8qvXq6MQ
FjFhcsRq2z0G6FHfgNw1+aAREmAiHthcjU6Y7/kly+t7SCoxuhhDA4g5vvl01loU
TTsNTPfAMiZ4jQ1mn7pXWnAVACTJwOaLpSZfhTnsVXFuXMmPsYuKgOfvTkxepkLy
LXmRaD1SejXk05v9E4sBsu3iqjRBTJa1uVjxL8LYxo+7m7ktDPhAzDsZVpLvkPWQ
X9rVP6YnWnme4Q6Ox9JFxZ/fVHU+nRCXcdVQlLxZiRqcsHFwPGRZWe5kYWEan6nt
2+t/CTpV7xnLrXXwHTlcA+2EiyMyaqxjSyFEBdQ76c1S9I7vN882NRbs44T+4kNM
islvG3jlxB5fFINNWimeuRqafm/3nL7fMNVotnMHGZEbfY8m+08cV2YQ3Yf9dkU5
FlV+yZOYehDEm6A2Z7WZwMr0S9Ge0nMx5IkeZULCKMqOUg7Wsf8nwr/3HpdbwJBX
bkCStau3/OppmxdslQchKoxGFIRlxPFh5JbG8sIJAELFUMyTdAk+n5Zi0Rq6VBfX
tfeZw/HHHgD8dJ/IsRNMj4h8uIPyf+txKJfwZs/gaCW1xmgRpCtlePam2b7y8yXz
I5Udoty//BsiSkrqaXUn/aW2zg0CF957bmL2HizFpXEpcKJ12lI0t0QfttuvD6jE
fEuhOlhKrYRTWejeSqL2N9Es2P4lYkeEuYzT0CXn7iXChS+7K9dvOKhbR1aCRsxm
sQgIzvZnkzGi5tP/Rqqr2U4czlQUGwlR8PAqbCs9WGE8RS6fFh1gVEJKazEsXJ7D
DVHtDCLv8u9nzNnqhX5obu7zoUtOxsawNGjPmWbfeWwoSM0FwvcborEoVXI6wj5u
D3QK9uOT5xHq9TUcuW6RIDdvjNsJfJ7GttygG0Ub8g40r43G4x92HWtrfkwOgL/5
RTBUj9dUaDA3ydu4gZmEmiU/tMDWQEgVD5JitkOrGND6l3Bi/nsVzZUy50tTxzPR
lexlKfx+kQV6zDUJsyCa6popxu+KSjPRCkk5nu9n0Keak1qk7fqMFUHCbuVed9BJ
4UoI0rw8WsbEFWgn3WXrWOkCJMOCG/+XTmAEmRig9HzyTvyikNzbsCUjzo7IQXAJ
dcqc28lAgpMd3tV+rR0XhpSTB0aV15D2BJFFKCh+fqMIeFoIuYq8lTzpC5laQWQK
C4up7YzZeUWUuxE38FjBeL5WhP9uZGfmSZQKAzlSnp9w5oXa08Xs83bsiSPZBQt6
DCvf/jJ3wD2uTHPG2DYoweslIOspLJKDjaNWQ2r+2oCyckAvws8YwdSVgeM3qbcf
K3QVpENtWSXBWIJ+jIWJ96L/mlb3MasEovzv//ifTlZQTCfNbbSX0mrnOnWrSKp9
EmRkLdNq57BIkMTdFrtx/+sVlKsjKDZeuRW1qB8uV+f0Y6BT0KCB4bVqYf+z+FYF
9aAqBVxQxwCbH/S9dhxlNflgKj3zCjGUZCq1YT9ICdZjUINsif7kZQSARbGjElws
DjBYjmhmziEJkFjWV7XVsojwvmT6zk7ZRpFLugx6/GxQy048ueUe/ocvaomJ3G5D
mrcb8vhW+cZbk9A7Qfx+VyM9oJ+G7yrUmTpRZ1YuDVAhroHgAmGDKeFxpFEa8nNH
a0dErr4OIdp7a7XOG2yEf5bCmOf0DjqReWQAs6sTDOVSLgPNmj+Onn9EgUaJrOr8
3WaIePwDbShjwLfXkFFAIXx1K8W4uzUpJIFHt/SPzNiQXb8CWbqTmMDpP7q6vI/3
L8QVIJyYNsYjXQxV6iHoqTI5gOgGIGo6rl6W+fI+b1ZY+vpCubC3tyxpRAEYvcXu
5/a0aFyRIpBO94QLobLxXHSwuUsiTyOxAd82i+grmmxqioQGhEqDhr2ssI8EyuQQ
lnzHbmjqR1FBLgrKPkuyQFfNh8cqieg/ltzRl4TYu3uxbFcZhppDvggigE5q620f
/LBiBfKJ0ERxhge6vKfeyztISN3rn+3abmT8JGeAvaB4hIN5J5Rd8KxXt7zg8uiD
zShoMm+qYqoifKj4KgaRD4y0+P9S669pvMdrTM6mjfXk5Q2AjSfREb/l2P8M40XC
DxkkVTc+71Vj5gXzWSyyqbHzXJFcPuxHnxj79nGgcCuhwr+4JIJqnI+HbgTetY6R
gwHPniEG/xaflxspwOLFLhR/iLwew2jCcszyNtXhlQNsKVBiG/J4FJHYdmpIy3YC
hU90ajB4rQVYlmSBp8MPjT2M0Uvlq+f9FeqU3ILDW5Xzd7ZvdTR98/+hjakgeNgk
Zt3/zujyUvId5PMhVfHdnLgzIEPb9cVe+FuI1f+mMbV8oQd14aPszuGN+RSCuyAG
+4LS7as0Nuj3pW+7LsN1yGTvu5mVcw5OZXO03PI9Le5J/sY9OLSfnEetZt23RzeS
zCs3CH9FuIN/hnXsDUSO3Rs0UMifFbB0Bn+1Y+g9+9GuoCLqHu6bhnRBGWl4IKpY
YaLl6fNxiZml5lOwPYUUxX36fjR3JFZ8S9KkmAvdZY+Aj/DQtFaL9rXbJXr/xR9l
sttnCaoBExDYlKgXaXvw5iWIVxvYQGEYQnvl90BG4SK/jrSALBn1W6BstR/5g9qP
UkVFriWIzoO/PQLVjLQY3pN8wXNDiqZUH0/9MOuHaWvRFvulQDsjWVD8qgdGxSlr
uJyaP8y8f9ls7ybdwr7V+IszGOdIJsaG+G5HymT3mZFxeuIr+qidZ/2nHFO3wf4b
vTfcTjairFSOElxUgajNmY/DXNZRkvo5x0znVmkhH65sl5Pks3Z7tSu8HGAdsPdm
t7UUv63HH947qqzmMRi2r3Ru7o+XoFJt9FwPLYa+JlAXE+1snSjNC+8FffY+50cE
VNF6iyDuzeuOatsE0N5L/mePb0NkURCCPl8tVajfeiKkOkteblNSk9Wt1Tm8xiaM
g+nGgi1sUGW81mom+LDPuCY7xU5iBRVWuWl2BaUE/DYRjjDraKyjtitwFmrub9Z2
ZM7nijGtylIQTTHY3VB4vNgXWWwKHOxYVC6aqI6sQEZiuRUv+PkxE5RHONm8p3xW
V8AT2YBD6mwX6xOv6rBGQiVRds2HMDoA9nR/Rt9QOW+IL07nseKFMLnBKu/e7Din
HlrDhiwAz070F3cM2PwcsnMhtm4A58+pHsLUc9jJBooPAQR0jAc/1mxFI9rJEy8p
CM1T/+kfuBvqhb+9q96UTA7A0KgaCyKPwEn7WH9rQQn6gm9aWZCRUfoKsPFv6ah7
bcfnkdiS3rVazLzVigVqRnCc9CRFR+r00VqizHHZjPAp2q9gaGhyehfF05+eYwAm
E6O72pAuohjkFvGk2XCSFqGcp/mSrBAtHzVB+Y/mjRclLvA4Y8PYBBLBdWaBaOK3
mPLO/OsZqC7P3IjkAcUS71QyL2V0fvqOAQTgG7hqNS9iEV+LobaU+qzGuZFZAh4f
1wBaX3IuxVaiz3opiDfXmGBjjH0VAgulTjCxw7cs+4ZNnidDwdbRLsOTSHmdZzqc
HkoENk48+6nnXvGjfNED43m7gLYuzDZzhNvFYR4dJgqUTT7Fp7ohDJ426cPhux0y
a5H3dlKkbUeL5jJzVpp160+KqSx8LoAnPLex5L5Pijat2uj89yzSYME+W+QqSF25
DxGqtPQhKJszqfDS9hy5HXWeRgYg/yOPwU1lqtVO1kCoK0ZFQWSBVx/4K02cOlCe
IPY7px6OFjayoOE7oN4TJrgqV08oGDg63M62VEpcr2iYEwNwyBPV089PJL0Er4dT
XG86JK5gtpxZiN2cXyLadQ01mT6oCljGuYxJ2k7kIY1uAJOOsR5XJPPB0rbrSeGm
4I/xwY/y7u8XXP/nhbgCaN32rNDH/4WSPpuGJTCMe/5E6hq6Uu5LZ5h/z14Hsc+d
ZxArpyvkUh/MHcs1YV82DfY+y0HLaUKldVZezxcQDqyUVMorGtWHtPvYWmP3N/S6
/1AyS/XQy/zDa6RW3UexPAmHXsR2nPvsaD6hlYPOTFwtyQ6maOJNjs30oisdeY21
L6oCQpoo28pURfuaLUWOB4hhEsOjtTSCdbZ6mvx16BqPzM2BuAXmRKjoXs+zML/H
TFakOCxx0W495LZ7+Fe8hF5pHncdU0rYoD8vfIV2Yr1lz90UMC4Bm6dtBzZ03pbW
8IGW3YIpCJzarAnpth2JaXMgcCH1n8k2z7yEnUt06yK+QTA3zx4FSa4rQ2zckxPw
CDtTMnlVa6VbgAuIeXdZE2JYOKWCVrMsP0nRIOPC/CUtnb/7TmaCkEji+SlgT0ag
ZQo7sPC3bmhMbunrV6kwbpUMwmg2LafJvS19J/RB8z2p8z0ErRVD7VxWKRho6XUq
2QzOvsjWvgxEpe6Y73vvkEiJxe3UGDdYuFSd9EDodNyHfQUSIeiB+ARX88pf68HE
N/hmWwzdtiAZVcsbly7Lnkd58Sc4lHvIWJkQunMSuYZtX7gAJ90monZvVlklcrL3
O4XQ+34ahAw4LFcUj01BVoYPzScI8pIK/3DsB6DEcs+lsqh84bY11MIympYOsqrC
g31/gqJNEbQHMPbXjmiCGnQ0xkM/9MWt6/rXb9j+f8J4YQ2Ce0IP+GVZWqLUSnyX
ixGkz/xxK2+brSItilT/DxzZdpOJ/x4rGMX1F5HxChe3veLo51lGOlQB3rZx84hf
kb0nbGIVvKIqdS7QdJv0j2/1LGdHcwS/KdlPO5+vsMNxSWwEbJWuA0iULtcJ01dQ
aJGPVFijM22i+7Czh7QjijfWLymxWTt49oIsYzZfYKo2iXgTR8r+ml4Zj6RxiNvO
26uZFrgGt0/b9TCeWKnzOsQIIX6NsB21SiyxHT3HjUNhFo8BtjK5TN/SPXTTkMTG
AdzAWvI1eNQvaKVA34xX6rhL0t16P93Sj6GelyPDu84JrVRwf8X5bY6y6hVojK/C
OyJWjRrL+B5pMtB9Yj7I3phirFZeK0riwfG8Q/a87qrG0uR7poIVc5Td74mFF+XG
BfWVNoz/1+StgSgZJcxfs7vg3HDzhMsJNibn9h2J2rMBEQLOeEh0sOj8pSoKvlh6
j+v9ZW4kzlSyULMll+Q1+06FKJwBU3pn043Ayk1g3nS3jUUE60qCGRR0Kk2Nm1fn
EheqlAjl4HA95tnV99bD2FtrMJ3lPbKMPIntLm3BlXqU4uo3UJg/kjLeXb74fu0M
Q4P5FbELKYCNpXZbtkRv/4R1dnSJwlahnymEO4Cf8xpK3bWfesBtLxw8kDE1I+tS
XQ11tTUM4/On7NE8/MIeeWpTCbYBvZpL4djMuAvQoGVWxDC/BV+6acUVQStKqCQW
0Bk2d7+cluqoX0TC5vueV5TaG7lOQ/l8pYmSB1SKFMP8uppt+Gc4oDPPDTWLqH77
sW+vyC7UIwsnSxNJP392vwF3w5w09gmAOHi4GPsyuZz+U+faXJPEZTKUZmgGrzhc
uGrgzNimWbofSbIPQFBAsIrc1vYdlS3Uxsg5rIXwP63FM6FGIMpR37sf1mnkAR0o
vYXPrJTOTgnWAlYJPvpay5vBz3ab9dtE8eektZQKrbUs/ilHEfSCciFN08lkJcPi
Do4EhJ47HPb6Dfp6JCp/8zSIcqGSqqvLrpnQx4yy1PLyZeO6xVBy9CeFSNUMEqvV
Q+hTjH94N4ZE/tY8ajKi8hDYljkMGWcB9tz728OknVGlWF5rAtXdwyG5Or9jKyH8
YvSnpFyrqEOpwIheyf9rowPnHjZEsSXtinICnRQydPVwD0qlABRjru0gbs+Bki6m
eJexwCyse/1UmH3BtKxEh9biwSxmX1+CUjEyCG6mV0hkSTo2JrLtfAgPOZ471AY8
z9Rsps+L8gtnUi9QVR82eLHIhLkZeIg0Xd9bwHyWq7DxjTSUvFfZL49Tv1+dJ0oo
I2u+EgXWaZdNcqeZGl0yH+nqI+UmW+Oyp05eu52BoI7Jxks4SwE2vSviEIKXWDWp
ApMm/RsqL7n6izLRJy7ga1ciKJCrLRUk4a8pEIF116mXcyT4FUQq8IB2ccsTsCfU
n5tb6jx8zG2YRVo+xh85Y6rn1ArQzcw9W3clj3r08Sd6lMSArrk7wrbbBgV5afz/
nE5vNpGsq5bPY8FL94MtLCREApsYzPhFg6q+Zigkuup4icUDn+ljtB3No24ir/C7
pkSLGqUSoakzKbsq4MXHqzfAmRx8sYpyC8hpMuMja3mU+wYe4Cdq8pLdHK0ecDld
1I+nmIMfdpHteVuMc2QOyoyQErhs8n7+Q0nIhYakYOg7kXNFSVE5JGF6/V69GIJq
OwG+skYQqTrf5h1zefX1X41D/6fOMPwu8uCKb8PA1zbgtzLYbjrryFpPiN4dxP5G
xghGP3QenBNjjE2TtqKDTzJr+WY75HWvGAh1TcWZAMP+dQbIeIvvhCHGxOBVyuzV
T4LbIByT5Mf5OwxVQ1Kki6K6xTaia9/3fTuUwFc9kBmH+xKTEHj0R9IJ1ajoyuqR
paoGuYWieJ34AtXTZxlSUqNwWSqt5b/tdhOOwN+O0JcCjZLU095bPUhnGrRZtIIV
eNxAOJ2ZkqaLS47dXfCqrSNjZl1nCvhFK7rYVtCNhunSXpv0/t4K7b+lez7dd61C
ggPNfqLZdykfUMeVkFQL8oADgfXxotXPX+/elPSY2g7oKolpmw3678e42Dxded10
JNzVZGEegPWdNg+iv26nx2CTRWvzpwp2NMSW4XyIXXgQVDnJYxXaaWDkdb8LxO5G
a1YGbsk5b3nfaxhijuvdX3GYcWERVgqYN0chLpJkpnz87EmHNLi0xurgQ1INMvPN
pG4Lth8TueNRoFc9ydxtrgnkgQDATSZldv44V37cb1eOKo0TMd/Q+O3MieC4bfhe
1hHloGGYrd8I/HFyVkbjfOXXh5Hvy3v+XFrnvdxi/hVHcDHsrhQ1MoqYk+toaFuT
A6hosBGhXyelQZ2790vBMpyOP7e8i/WuzfIjunX+Qfk2lMTsZC3JrIsDI3fIq0n7
Z8h+/vY4GqLVleYqGrgioaUVXVgXMXHAckyo/XFoQ4duRSojJaV0AJpKntLUlZBM
Y5a2mZ1fjWID+RWvTvNOjAtPqpTd3LaSB4V2x2gStOkzBsGN8TGu1b2BFY1FA1o2
eHbAPCXUT2kmHt920rR3usWbaig5UlpcChuj1diGWTYPZk0ouBeGfP5yxx+Olp0k
rsLu+CODiAa/hnWRe4d070dN6l2G5+VBYtdGR4ldaRSKYjtptjO+FRYLxc+OhQbL
9BupMbiatWKLp1OQX93d3DN8c0RtwsqDvtzbAz1haHVA+DLyu9h2aVq7C20Hd7EP
VA6AZNVvgZWLKAQzzuE6pnPXunjk6KV13K+/m63pcvh4ad4CBOpAtYg1hoBeOo53
ykiktG+E9jueOvBGnN5EjngW8E4opD4YvNZt60rJr8UykZJzGLIcPcrOzsSUmY3n
cqFtClMvATQVrE8nAVEleDsPoUeQRM0ci9BkDW+okgrc79URuZVKwuy7q3YQk5Yl
Labv7EhStquRWTGXLz6TFwaqbhynNJm5L4zYTxonBT0WPGP9NGLD4pa+bqxNWsJx
Y1rnoqxBMc2F2p2JfgqkCVsbcegeaH/2G1hVemscxeKI/Ax6BBqSk3GeJZlFEuPy
UaJ4TUWcCMLGHEi5i2kFOQ5WCUgcwIYUsK9PcGVndbBSNYxqmm7ER/pUAqAynanb
2xx28saXNjw+k74aLu4beuAxkCEvpUkn/FfW7nq1VmNCiSDF51p86hCLF0eEtcn7
jnkbqqAnSOGbQvXHvcvoqCmfnpQviuzZxb8XGCnlsd9xLmiKGd2bTw5suOSNTtUA
zy1iIir4NTW8fjkRbgE2eZyYlQQZFWjliuMdDqNh/XA1tQGp8eP2JV4e88p6KaYK
yMF6cF6ebq8QqOYZCTFO3K8ztguwXDrQK9dTXSHgXBQYChEjPHM7OYwVB8JAkISG
JBo8kR2VAJG58FsY7AGYokL0NITMLzFJLBT7es2QhGH5//0laFAw92CTHVDyqyyp
78jXHsvzpeUfTa2Qpt+EmrNeeWPqTb0k0uaYrEB5kVzNzHJN4tOmRYQhfQd9TzQr
8Rn1z17tuKTMqDJQxsHWYn9xIgjQ67SOS0DtF31m83LsPEqbyuiHqjdOnuWVwm0L
VYZqGJDn7h8l7cJ6yyxb9anUaK2CADmPwQqMcfFUM0XZATWi7GfFW7r2yNg6nPs6
6KwcXz4criR7w0bG9z2fOgel5WnBnd0bazbiGATUosDZhyqFoEOj7ratUSvkAd6R
fzWJrupyjonDnrZQEjZ8rh3AxK9+DNWrAqyvXSoUt553VLsqm90JQkVNWWJW/Zry
PHU2acf4BiBjFwPIeUGE2tcxslsyViIHAjmVIGslAAJH7sMLwCVGYq3kWi5xm35m
T8yQKtl9DNhbzsm72L921U4eTAMiA60/sXBAHac8fmwhFwI6sHqMuUqkXqyVe/I9
+tK6eewKD19VuqwSj3PowcENrHt7QbUFV39gv8rYjCuwwZvUY/Y8/yH1rw/eqpEs
+Q49sDl+Gvm52nnQFoSmuPy4FjfP5drsKuIcNdmEjMDux88WkVbLNyOY4fwT6Onc
LVuGLfip0cLTAvPr7WVZrOOcCUNYfz0tY9kaFFUIWsrpXzLUi/6q2iDdrMa3eMmb
XmSEyjhg36NwDaeKfJ7mBwGSAHKi08sCvE4gzyeHHpGHwzry81fmpdLqeEZuJ6d/
LQw1H4HaqaKad6TTVzVLeVWQSoqIxfWZtJdkqxFTCDYtPIx10LgKnqK7uxDRfyTS
jJgs5Y+KUBjDYde9jpRpV5+l4AvRBg3ybPgjg8Dv2pvfMEbdbMlotzuTP0vBLYzj
SuMDw2rFhg0s+iA5YhwIw/+FOglzMJnFfFoD3M66b12LpjxV+kueVBTOzzUo01qw
soI8pd+wO4VdlKb5MiU56oY2lBNHteQ66G5qzthHz8wLWI6uQyrhc2ElI767rZiF
HHvcJAOLuyc/hwXbvrtzIlwZcXvaKvyBD3an7wwpY0oHqM1MHPJOU1qA0IfQSOoL
jrI7Gf3W5UwAWsO720MWaUUD2j58uhXH7hzSNGPzXg7un08k294OedxJ2DMSaWZq
QJBDEitHZTvFS4X/kkJNf7qEczOqsKt0rixd6KQJwSFYn5yTZRjdQxVxoGI8JUht
c+ZbW8UB7GzUHi4aKA7hybMlRLzIRpsNejLXFSeDfW4nErsG6msy0WQnq4ZeKKIK
CNDkODIoCogp3hH2iEUhdPAGY7YOUcXWrr5vI6TyVIzdqJ/PiYsyOY3WDTcM3FaQ
ngvQ9ZvoBcVqqGcZ8MhpU7ZOW4ARrsddGedI8Xg9fBcr/KKVYWZjnkVVYTgFBiQR
UOXoC8lUwsmsQoTlf0qZTNltbOa5t1/3NDaRuR9XCxvHRTq0mkStMJtMEI+6vriJ
pZxw1K1h8o//L0q8vdeDxYl7KMHss5jgDHhw41qjL1B38JotQULivGa3rNINGCks
fJGjCdsVxX5W8+tqgYdHh55MaQ8I2bCIUkdxx96d/Nk3K4284yoi+EHqNh5sN/ky
4dEz951+9bvB895iWVqjqewQovayMQOjmh1f077S8oWvoQlGCNYFnBgfTOKQdVqn
afICx9ZddaexUk5xt9Ilm3fW/1c5ajl6KRoD+4u7ak6fij5lzwzuFI6pQCblhFQC
ZlG5f5ht8zgRCS4rfxKMKLjvbx7yi6EZMYJa+aABigdn4kyk26TQjl90MdHU0AxG
Lzx9XRhkt+8XRP25Dv13SnhEThVoYfF0Q5IW3Sdl43pjIIpnsHE98KG8rA8WHppJ
dvXILduU3BJOhk8Kzz7rFhGKU6MwOARYQ1zuRJn6XOAx8w9iowLyTVkTzvhk+llK
Ufclely6QEf2I2KMewp1pNuWK0ZZK+PG0uGXeHPEzL9ffL722ZCRsgq3Mud7sxq+
1BIWossepNAY29oumC8sTYiN/AGKOJ2gF+hoq+8fOXj+yj333NdNFSAAH3OtbIc9
0T2lGFxJcn93NgIPb1zLLv2RkjYCZHz3uMJU+iPf/IulcY6oA1M1uAna4YVCrQ//
J4RA9h/DT9VuK+eVVWj3TGo3XPjzHjU+grqX3F18I9f9o4sXHXV2a4jJEUkhrh1b
/Z/3qygtWXwhyModkYZY2PjUDA8sG3ks9SKpUeBBTU1b1vBJGXUmE83YJAcdUplK
XYW3UuN93iI8xvl8iG4dV/EzhZnynPRcDbrMDHkikRkpJiiNQ5YyPqL3Y8R7dxs/
CjgaU8ihJqacHvMngDqLq+0FStLyw73cCNUxvW7ZcFkin6q1+DiJ4wEqM+C/tW7l
KtNCCk2OZSVUo8Ik0lPV8B/xpgDqlrwNwFKUtlV0oS3VODHK9rK6bA/SmDos7moL
m1DKkuI1LCRNwMDUhvF1oZKVRFgv3lpEMACjC6pca8OUVwWbmm/bjJhyAhhvSarE
mzZ7mhEd2F9+r7pEtrBkzh0sA0CCQYAs4qH+HraTYGlo2YVV7TG9scER+CV8NnUq
eQ9nTrS3kdxSXdNbpdRAlW0J1Be9WGiQDYWjkMFf7bCGi6J/BKZTNqNx4aETMyQV
rAql41lCfXPLSF0kfo5PDphCUXL59sSAtzyhOqS8fL/j9ghfIVQe7EHccljSGUPw
6hVaMwpqACx3E5CrhS6FpXWBfzRy/VdJYR+aOjJkAtHPW9L5g6O1g1hYV6xGzRyX
YSSeOAnv8Ba5DfjSPH3ISM4qXQ9YCwdH43wMBEVuGeVTsP23hfz/ojuxsGZIn864
XORC/TfaKWKz+v+EY/mfShxSvGdjIjDiJBQI0+eocInU1MBUf3qoHmMepl+QnPgS
7vsD9JjY8CHsEDemKquJTE1kZunVPU5lfWwLobGPZgsuLnEzHbmzsgvzWQOteT36
vByDJhj8YiJzwtcVzkf2rEkRJRnQ+2q6iBHAtFQoSKMWTVm7LSpFp9Gzps1sK0+y
v/mshtnXNsH8+nmmvhK4beAiLyYb9SPJzCfqokxVAcOwRW/YQSNjeUbHMc+sJN2i
rIxxWf+uxPtmuUzHAGbXkvrtNjsRP0IAN0UeoL1/CpaphNIwLvNlF1EV29b6YNlg
cZqilZ7OW+fDWBC1+wiPiZfi5RFUAwNviDhOz8MqJL8EaB8JBOVJjEISqC+2gVd6
JokAgVddZE6E3Z/D9eUUcIOyEojRYgWBOQN9sPwCM8VoNiHbmIYFpbH1SvfxAjl7
krgy+L+9wPTGqjXrvxtmbSz8GLzkwO2LSNNqdUv1e6Kfz+bYYfe+5ppSqudpTbGY
fIQ8b06N8yNt0dL30+VUPUc4ycQHNch0Kvq/R4iwYJtYp2hMER36cEv3Wh4WoKq0
IDOXlafxORtbViat20I2vAnHwCFlAKvpd4Wo70m+spv6MZ63VBeRKDUPvp62h+4L
R2EUQym+ueDgvedHix0oz3X0UjLxXTNq8CbozHoxEA34qRj8peRcpRXZc8XEzaal
DZmE0Wm2TJ+SP+rXnY0eAyA5NULiGR3FxWRfBUVArLAgNzifCk9w5O5oJ3YtRqmH
oouwwkS7XATtYPSEdt8B5p4uel0au+2OJzLcPg5f02POtjBN5OFEcF89XPCPtJDo
hzCFVkklnFfm+K+VuLJuH43Q6gg/2/c9XHX/qeGQ0+eRr83K0ZTON3jvZFZEmGaf
gnQf7Quo915c12xKZLKazCq4GG1DOWVwkBuwp/JVRDinOC3BWkTU3F59fgOkmrbw
ilPpL5S+Yy5Jyc5kVP5WzR2s1wOGuA99jMxcVMBQ/ijPzwiIN1OhP7glP75j9T0t
BLSFhlZrnb3sy+PVHJr0hlEFP5f75yHrCMp7NX4gpkIxaFbyqWJrmrlSeiVnEm7n
Ss6pqPsCSGJvVKF56YECsvPGxvYr7cYJ8vRv5+yIQEz//Kxv3c3TxNAb9t9lxRaq
s5NBal0ycB02uHz8wJrQ0ZwtyAays8LR0NN0+L16mlUiVTGEySOrElC7WvlojP6Z
PKG1NAyPbbrngNPoJMKwp7/XtHnxOd9FQxhmLrwm3jvYYb/vMi62s7mCpcYqsMZm
z1bj3dq8SK0XU9Jr/W11x5j407NMH/HVoCI2iLlpBPZwKQmUofDnxd6REzhgfw+E
AskxSkzd6iateq0dwBddc0P9v6BTKmpqUAi1xYTFx9ouQmkrutqcC312YK7IlTZD
+OR3gNKG2FYsv4xsY1n2JiR8dQcid0vQN46rOwlyPD7eJaOnfd8mI38FVtUeHFpu
zGuSVT6dFknadlYNvg3AI7KHDF8Nx5CormSLGlpqsppCvAy9XcY1rBZ8qOVmDWq+
y26PxnZiwoefKl15RrJKP/09CW7feTBy86JwxhjGZZPskdQF5qmfwWRe6MGRINkw
SkCZTxkVhnni+KvjpE/2RcvEZ8oQ0rZ+0pcVoL2CDQMPJPJ+oQv41/9hSp4H/xHf
rHjgnQ9LdWESbbLNNhjLjmHwFXGKDRfS1/sFS+F4twONk3jGiNcNtge/TA39dpkn
xGtN2eD5heNXGC+JTAjPkip6mmoOUyHZXsouUuE9LErdQx3xiJOCKF0nJkirFpI8
Tncwk8LlujO+ccNIMtXC3h/YFF06q2pXZzBNs88fWR1Ln0TL5KxBdFFjQrkOqPy9
iEvo3DpnypdL5NCB7MGgVQs/gJBzyEPLhlgWkhbVXMYgmYwQdt4BsMiDzWJwyTAe
ls8D0L+jsQPhVVj7g14MShRsW84y4GRIHQqSIngidfAJ/9pot0PGYisT4IavnVja
QxDNPdgF4Io5cjMZaHULKyqOK6NYGFX5ZH5gK1vXZtw38Dg1R+iBKdbTL9eb8Xoh
dJ1rb2KMAEC46QaOD3Dbx5K8siG+DQi3Q+ED1cBhkS7MdodcXUBxP9Cmk9+aITeF
Z7qP3kvcN5ohaz8sDYuPFu+QQS3sNC9yKILHlVAZPHi0utWYGRWr3JF5764x5wba
PjUUjSVRLmixHuU9WdfGmEPtxOeNX3DNjXYBlp8IXpMVwPcYMpILcYKF/Tr469Wy
Q2uXmRDgkL5BXA5DTrWNQ3gaT7eOhlPo3T1DMwqLINjxyQZwSLm9UT61zmhMkPQE
g9vcknqjwa1YRDBOqFqpV7aEedoxZRAd4Cb3iXT/UCeqaEpUpH9RXM0h0mdxz/Ay
hOTvwEN0OxaXF4Boz4FxP/GQ1BP95odi611hYKj8Ys6/4GcCtB0DCTLObU0rZCv/
TbDGERkEjjRBWRc7J1CO9jV0mQjy3y7SPzZSKh6dVhb/LXjw7513LvuPTt46yt9/
YPBcxFyEY4XcDE5wjbjadR5rD2P0CCZP1aPIXetdT/UHub+fPkEgIQ+ocYjgWyDi
zVEe4LnW7X2syOjF8xAwW/v2hdKcvvm4rUpw6bsq0aEmnsgCyL4aMqxv0ZPYpvso
z+uj8cdJD081m+7gLgidTESyyM7G1qkMLmnwkC/hyetJa3gFVwvwjwiP8PMJaWcc
vanxJbCv+Ts/Hae9GsO+BaNBMLGKY0C5TFA1BUacAKaZd99G0rbSiH+vc40mKKYS
63z3TvtVkJk8n2Z65UoqRS41aYqkbB72iiDZXDPJLiFKEDF2712lVsbT0gUm18ue
q7mWMi8PDr8PflsAB8J2teIdhXJRzjDeqtiZ1SqEkkTHboSZTYNqEczcy0yQvufK
m8DY8srXYolwz1/S+yA96BD3CzLvlqSXxxw9f85JM1pOPK2z2ua+UwSYzI4bjrN4
uu1TRVadAypA4VW8FBdS++/a+orTZqENLFNnZep2rHKla9vusuXC5WuFwSTkyY+X
btHc7arNrMEeOQEhdBppHp7yGW3ce4JPj4ynBVsN64jQ0Go/hAA5K+fCT+AzadVR
twGb0uyy+DY/QtdJZy+2T+GC16HxnUcuc74rnDxd/D1yw9s0BgR8tw8cp8XKlVsO
TF0+jXX4asXC+QXuvFmvjW30hMKKsXlZnqSWXjsqkxZGqz+RgbnOq/5PITtXz2Sa
DW7froJf/hAAzLolgPgM19jFCSJRqD8ZoF83x3c+O537WY1E/hycM6dbiZAeoPbf
FOh6aKtbP/kDX4uPXkKfiAgbwu/vUvp9HMeuZ3cQDUzRHkTiAEqzpmCctAUNO3Ud
Oat2Q6f2QFNHxLGawRf11u7Qd6dnIbrTdwAFuFwOZEE4ZYFhBDxDcOTIHjtb4rAj
is0fQHsRvauo0XJST3OYQLE9MNH6Wc9gTHBMCPAUUZ/9SiFCc7UbNSFWp/mooMXL
AYvjv0eglIV2F8yXsRTnAQ6/bnc1JMWjyDu+rnSgKm/Y7lCuVmhJIeR/bCaeKcDs
UJIAHaT49AQj1tS/smo2/jcrHT3S/IjCq876chOy+3zpBkEIsKr7UpAZihucOizv
dgN6vIcMZzfsDvjSofRDe5Cab1jkhvYeGdcZd17U7MTrhDr0aBj4TVZR767duTpv
Z90Ra3z+4kg3wsS0Q2Ha8logo/+hLXIjumiTYeQislDjzBsrl9N+xnTyovJ+Dxn9
Y0aBa7pHNZ9yT0IcWvsbpDlKHhtcMVr8Z3BnnGNykGbA+q1FpgJJxTQcHe0Hd2H/
BXXPZZVyGCWDcVvgt3OcqaOIFMYvpe3giNfmD5pP2EUgNiT33CzNpmj8W6SQXb0b
5WCwOFdqDrEGRFYVwpgELIPyUW2Tapnt5ayhoTx19Qwr2P7c5b1zCwsgfzfy7J0J
IzHTP8P22UE8pL8FUSZSilI0nnsxidnm3cx/FsLbWTiEQ3MNmZ2JP4Kdvt+5iwbt
gTOeWRcXit4doafVCMJph771VtTS4WvrXXLDNsj4ZdBhCePQemLvdLYwxKaxLrnr
z3NuZVynLQleqhPm9ATjsPkx9FkCjwonMouS2SuJbTw3yfivI/T2Lj9Fxw2Raebq
DEHZ/PmqqJv6znUXEMj+BgHEgQ0qH/SapED/D5dJtlphp+UxeZaTh0p/FdCOvm0D
oxYJ55LXFOrkkH4IPLWbmvN77NP47eG36Okc2FXA9efzBkS4uvuACSjEQ87j2NU6
BLK2SGAbNEkMClwTyGx3ah981f09cthZdgll7xeQbYifOeEfvb9bXdVXxkmzVNkz
U1hkcFlkCkJIPQCGJI9eEkfSj7nJY0DzIIgQBQ7Vh/MjXqMCEgW1lxFZIl6+79YL
+MwPKy9vzngczOxTxnjhxWk364U/S1vM0N/07Wbzy/w+amb6Gz4ge2jZfJ9Zasl1
6pvFEzEoz68Z/OLMMG63gYqvthc2gC+CgaULDsHyQk8pB35QhS2L4eR1LRx90g4Q
rXr3N6bXbqbgHnAFl7YAKbsMgSQ6fZBmKA7HMuGk41k3MSiZamXLUQC2pFIabxJe
lXdhfOhlzl9KKfCLkfIROk607CZ00qn88EAl2ow2zNCbXvMBI7bPYaC3xhffuDG8
DwFSkiFXtgz7Magc3olWNbCkp7A+PP4UtM9SlXZffbwJAAEgUbFWHqbfdRs72pSv
qTGnUANePxD0ug6YXkkKbTEvlKDzscVRxF2DH6bI9FpAtOcyAItUtBbA1lsHk55g
e2IFD9qdIt96srlMA+HKEu5xfZgeVZlYJ72p2Fa3EkJZfSmroXxBit7rf6ptFXe0
3UVn/2u3yyjJ/WKuLlv3cRQEVAaPbk6kvBPavBxXT/DZa2KoYBRpbiIarxj4XqGg
6nsYhaIYJnF2vlGPlq+XBRcwv1DqrRtquAaRr+E5c59chivFr9kGr8tqSuHmxN38
RzhNUg4+ymjcjWGYw4kQ23gUJL+hNNjb3rDwB5v8TRFZtbfzQby975ejtNIfIrFZ
fjcXtQTrH3ZUJ/FY9YMbKaqz4cNIjFR1w5grvV+g2ILGAq/iEmcJ+9B6WDUBSb/N
uNUTQttIOa1OFZUM5BJK5mC/0+5F0Qx3LbRK9W3t8K+mHLKhBR78lxVvkwq6NnRp
dcjgwYC5i+xeF2kA/RcMt4nnrfj32CsE49xfYapu61LA28gwbGr5DzKCDz8rMqHJ
ysq91oI2AdwTx5vBmIQs6541LW4MLFibPmo23Ag5baSNPJSPNbLLsceSPg+yet8j
Nc4X2bkFjtLoGpSDbpbOTA==
--pragma protect end_data_block
--pragma protect digest_block
OAiTJGN92f2Ah81qzIhmoeVv944=
--pragma protect end_digest_block
--pragma protect end_protected
