-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
b/3x6b9AYC9Sav1TKtIKAaH1rpR2Vinpb2Ksc/yOrGJtaLX04q/3UL3r7kYfZMDt7z4FWXbYo6oT
ZPX3irvVIvaZtFf4XFRNs1UiMmiO8P4AsbdKjUBv4O5aVKsX+byRQUrvADIQtWO3YXJAkDQCuyTj
ixQqKnIsB07J+SIEh1tvW0PXEPif/x8J+MJm14TfYnYus6uVSSxZ2+B44ZH9+pNfhONtYXNat+rQ
ZYOZch6q8T0FKF0b+YRq2uSqUQ9w1qECJlGn7Zfwqtr6ej8z7wvMmUySEbUs59NTYuJDvjkLI86p
J4Ac0V3Y4mTbN61/5QGhk2Iz9w6DUkiMCK6D4w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9248)
`protect data_block
HVcsI/qxJCFVQgbl+VMg88Me7JMn6gQ6f7gziamWRzaV67kTfynfrjg5xWL5Yl8OQ/HnHcp05DsN
IFLHrXY4lT6kpKAAhNuLEGjcJ3rjb8IQWM/WTQh24H2sHHCnwtMIW0El6+YtsAyqvfqQUCW+jgL4
VIHaOk3EDGas0Puc81p/oY+RLsjMQM+TkubTDePLSerc0iuYk9HfRPhzAdVx3EllxBpROVot/2+c
KOkItfmLoBOfBnrSmLe1S6PRj9VWdT/1EAHxZQfT0tZ/5rKF78z2xATaCHhXEcbBgpBKQfQz1qSq
ipDIVz7w+CyYzJRpnvFYflH3k3lsfOndPVlt7XPrJ7xf5Wn/tQ8V+NiBoE/J/4Mr9JW9yObbLv5z
iPz6gKr6iAJnniC9ifiw5I7cFIuYDpq5srmKmR1Po8rK9NyR0NwusjKMlunSZ7VdV/IZr/sFzTbg
nJMa08OmACeZU7f44eAMjHMsAbhNyOC8fgthTvA4hd2Lj8yKNfBom3DqkkYDiFCp0CuqzsmL676f
eEpX0NOJKdhmdK1pNGetcov9DcdZR3neTJeBRMEKWWDVkUkZd+uBy7fkuVXjADdzBQ8GgcOkrcqB
meSWEqVARJybAIYugXmjt3Gip5y+AToNDlJogjVJnhGpN0HK7UQl//SqlpyE7voQ2D6l/w7nIY2Z
ZrHZWG5z+cQCA3YsfVQPvOkkVW40Lae4cjcV4fq6EnwpD6J5SkpcBs4UK5MYEceLlWi0FWTIBzuf
7BFRS/Z01JZ6mOzHqczhA40Nan86q4JI5SN0v3MOH0txMz/y5SRQQKVZK/M+FZvRMcpcTg53wRUm
rjqIVJDImO19tb2yy4XaVyMTD8d0r9ggMvHvJ6Ie/fR5UbcUVeTf8Rnz8s6mfzLeNFZlo/ixWe7I
iQd2OfHcfbQeAmR+d+w2y+A1TxH6qEFVKJGNxv5fqcrNgr9uVb/jdIC2p0X/AnDEDnAG6B9LG8pV
ZL8npBcs04BgNe5u5LJaN8OOVUHDNJBLkLqyvmzjVQcRHTp07hvLXyHrdyTceJVU/wM8LzN62VVb
mqNp1feHgC0Fr1C4HixaldR7y9nH5U2Jz3w8rPclD0HPDTpJ+V07asR3OrtOl4Wo7SlxOTD3cMEt
kY2OZQN3YYVQ0rFKJsGX2M5VNSaMKBzVrJ+WzCyBHUmjLOXU34shveFWIQpyE4Mzzce6LON6ylhA
lXGbEt2j/Y0LWYGQP4eFkUeF9fBqOsDnuyBnUB0i0R+RokAg2aFUMCig6qzEygMSiFN1zGBZcNIF
Mtge7Gc14CjGlszKuWYiE9/gP1jm+/LF1BWm+fVtG5IfkYXvrWkkqXb/Yx52qERDREdbGMMTAYLT
McPerobalc5t84yGz8VEAti1Zto2PP+2X+gpRNOWuK2lgRs7dPMknwWpH3u+3nIwMrNwY2Mz9MrK
p++WoS6DeeBQJVhkl3fD8JjijdbSVe6XSyXo+xZsh20YEGHllmXC3rGhDJg/qc3Ouxi4PESH0t0Q
ArL0co+rpc16hOjXc+o7RgViPQgV/rl211WTebpbuM+ubVOZOxHlbCsCgvVGF5IZFbXGPKMbV0m3
aqHqwphTlrgGitVxEfI36zchESLpdpuWuLsk5VmOH2zmxIdjftvISgoghH4rYmYu7UeDBg8J4O7d
2XouuXGFujq0H/vproivHT50D+uykZHM8R2k237IyQKNzZyFh0Umbs0lQklh60Nq/wKOzpzHDrbB
97+nso2hsHIa5VgrAKxOjQyD/coaYK0kZ40XoTAUdk7pV2m7k5hmibF7lOHtkXG84AX8kJscOEIa
fBVrPHdWk8mQygoe3SmFEwsQaRwWgzJ20Qgy/3vZwOkAzqOgdJojfL7z3KUVpokUosM46+CJnuKF
pM9SpxDSLCP7hqJo2OKsUTUODmD/gTKfUl0lK3Fy3VWDx4VEPIqTAJZmQp6tDfm/7HBlI5eZHyqy
vm05FqEv0PBNUREZKuHXXqhnW7SItdB7/P2y5nOPJ4JDOZ1fmzgAK2Ikw7BLNducWJGwzmvt13uP
420hggOVntUgaxWQjKd81+f3ukbBcdX1NtgaoVxOnKCfHocjoYAlIDwo1Aqxks43zuEPsUJQaiWQ
m/mTIzxxWc/RvM4z6U84wwgutO3KE4Z9HNKbzvQGydskB6PS/ecU5B2+wVL6899rAhJSesKjJ+KU
Gx07wmVZZ6akmrUEznmzjsd9sN6Ou9zMREeohJPTGF5e+eOV4eux4pCocV6DRhI3sDKiOe3ZWVGP
cVqcbgNjOYe7dXDjP9et731MooVJb8TXhE8++/0mz/vPOD0MJMLVeViPoz2sNj6p/IwgFcj2Iid0
SUnCmRfbn2PH0DKVhmznWdEZN8pomwqSARCJ5Twoecv8BvzSL9D8MKOavRPywy7YZ0nAjcx7BV5I
snAfBo2G4tXSP6COZqGo58zf9jBmKxGV26i41bwJAUKVGbg8gmEklLpA1QA4taGxQQDMilL5rhIG
TdBt8jLakeqrxF0zv1JcG6qfIEisV0iPAP9wpLQLadm0m2LgbOWibsUWDOY2T95MD19A8dfCU7Nd
80Fkh53+qOAmVmPC2z7Jr4ZwLn881OBK4Ly37f17hIEQKH26P4jZaZU45PobyJgfMMDkQyy3M2rT
KyRc8eQO5f4wglr8Y9T9g1ObyPCgviBZ1PUE8lAsN5pRnXCz6ha0Kw+TfheVTpu9bf9KOxSlz4Pe
OLqFYPKYSsAokGRACZU2/35aOzZHAIJuDzp++Tebd33TbgqMuj6p8nX5iKE0a1vtmpf7iYqBl4d5
NibGSkKKKiqf0SAADhMZANewYgnpNupX8uSeMOdZJmEIM5HQPgjSKthBgXV1adR8h2HNdDPnu+BV
yElXebRKlXv0yhP3Jn8t621CcylPWENzhlaR6/LgpTzkgvbIjlq7AqLWfEjUqO5sEU9F+dRARfRf
lO10cBKN+U7DUxi3uZM+RGSO5gO4n9rKOXs0EoEX+gB9Sw7YHHUO/CxF8lKWgcldtgf8J7LOH+J9
jTyOpSfSHOpwTcNlNnKAJe2C6O3K5ES5td4oxyh0YHMip6rbBB987Fk9pLMebj04WQNCtOaSweSv
hwXVhlz3KMxHEAPVRYY777q0ZVzZtqvm3ehcnR3dTeYVux9vieIfEUP2pPUHZfUOc25BRwvq1rjy
XrNWc2U/t2Ygu86KIzrhAIAz06ztwMKIoxBZUtk81zbIfRwz/iWEhz0Q+rRJWgKbNb+iQQSp8738
HGYi4P91qCr43B1NQOox69xwZO3tGwa3mlC6q7ioghtGwVabO36PcZgdkvm/uDYmnUosLlsoj8f6
cNbvogt1JIqT++VQ9om+nQU3fdC3cwC0OFvtej3bd2VEKEQSMUJPveCCdDHQ2JVwkrrCoQJ1DNI8
H7QkcHBAsXdivBbAXFpCepMzDP+CABGnG55QF5b0mjVnNzc/ZCmqeTbWcFyDbYyL/vpDsw+UyPr6
UGfNkN3mQpOCm09LlpZb+cxvSw6l/U/P2t/DI+j2+ZNcdGRVOCGO1eVaciYx5LwlpZ9lZIqr87oK
blBPrYPBpmqaGlY8ODEX5KCkbTObQ7IDirzggDjLFsGcw20VtZiK8XYxDxofxtywdt9lWN+eCl0T
c+jp29gU+BWAhIMyNYiwVj1h2TCN39oQu19jNTWdaLhcQfuhvg0OckOdRplntw4v0jzpDFploUSn
mM0Kh8zyTy/L8ef7DA9g66dq55MlTJhMR2kahJpwegLnB1rwdaA+2tNwM2x8bTWB8+OCI5FK4Utd
QrbMQ63mpXz4rLuTInZCKt42LO3Ec2+gCRbqeMzGPavc83A6NFrAN4kI7YdVzAsDIptYUpR1kmxR
IXdDC57IWUrEeXYmaoLiRmxKz+xFkP6tGrZ3HlT60x+VL31airQiB4368Lx9QN+WRw/KX/+focnV
rKb23HD19I/Y1/DKaLNhMzhpyJ/wVn7VUAJOyGyJIXXOUBQLPb9Vppw77eckhYiwVP5eY8+scl64
IQgT/TuCjDGDKVPE9yqB3MXe+/T/OZaqqYHrFzeN/bcu/aOYCCFnXGly+fxgTs+lC1XAHnn492O3
kCL/O3kPwDCD/ZoC8G4T7QEht0l/E4sxj4tXoa2de8cKx4BRTvQdW0UwkCkFKpgS52Siju7xI3rS
8wPQgeCUVrZzMAmv1y/giCUwgA8fmPLqhUN8UB1WwM/Dz2TiOWAdlFvlNGCebTQLhMP2RHlVYWRj
YNnwxLyD0monNhdD929uxzcKOcn5VyKzAeTT3lEthZWXm8IW9GGd2PM0NpOAzfo5SCwBcqZaUyI/
Q+qKotNnviNapO8AZxo+W5YgVjY50DKthesAzAS6KofHPZpELlrKoAFq+3zOnEi6bZMv19GIhesx
aqqnS4YEWKDUB8OC58eHuYyXO8muOl/ao1hyf99S/iS7ovtQsPPhrnk1aCry3wSXzrPr5cwab6I5
HJ175L4xzjfhZ1ZAubaLzC2ojyfKPCKqlQo7zzWiBilZjANshT/Sd04JHmq/+Rb1KneuO6tnjvkT
TSyn8izjrM3sg1gEXKJoUma8GybHOF6DKTdOamAPbri3eR0TAqvpRjqj278n5MuhxWnpkQnQx5ps
cgZnlzLNqG+LxiGn1SmpO/bHKbuF2G9FNXOooFLE4vjjmZ3mlCPkgp0EismessbawkWE9vHhzYSY
D1VUl8epDVRDmeoHYLHtYOc6ZCtuOxcs604vVTLmTqLrkbnzqWdwpIYy7sRIFVPVnVdraWhEvnLU
yGRfws5uXHEGqVUdL5+RPU+sE+QjUoC143VoP9xfIWQzOtdfNI3jaapj8Rggkt95js1poJ3juyce
MeVS5FPCJKjAhv2TD0gIpOtqOtdFrWJcWLZGg9IFlcTXMY0OeCsy9jxhLWVsJAQL3B5oeh5yqrXV
LNOhPaIYsvD8NAHSP89CBqqqBaU1yeE6lNvjQKGG6TYwssGgtPGrzEf7w/07Q7/d1nUgjtO61/gy
wSluHVevleq8utO4thsJM6DzmA95mBsBwGX3kMKbXA7PkWjPpCRIE1lSDgv/YnVMXPcIAULWbnKh
jBybapNbo3Mqu4W9HBPIVjIEto3tn1yOWIrBsOZoRgH+UIkKX6EuysAyu5RFWpq+sW2kuL0ehBf1
LmUthXTo3d8w7sLYDqbtUuojj+Bpst0pZzoGtc4rRCp7R2pQhjLrzXXbFMXJvQupY+5WT5zVXX43
1hobJmWjnat/9/wPL1HAnbNZkP95ZTCpOo82KMUE0wL0WsGJgDRize2m/8iE/Rw6pJ7nMw2UT153
GenVvAR6nXT9gdSjYlG4q3NCVDlSwhq89RDP7frZpj5WSQ7GQtvMzLikL756Fkj8h3cEQ6qLflsS
mHTaDzAKUYjY/CFoP3id4Fu9054pSmbwHPZdkjFi7ksw+d1Ut26o9glTIolbarpRnyqvR6YmRjS8
Zx4hBkYS7LDnsNmE+BI/8gh5B/RDX32b0ZoX7qcJs8zuoz12tSJ3Ub/ZgPLP/JyKeyuhMen4FWCB
vDdHf76AIOJHAWnVdPDmmtUtUjAmVd2QYIbqLmh3JZi8xHlUT5qO6UZTb0MG7L4aet6u7ot8f/sO
KGRFh/ZXCwJ8whefFdXWFfBNLXvntnQ0vj6sZUGSD03lbLOx8u64mm07alPvOVGApMWNBhym+ZlJ
3GROb9D7gdIeKJiG/wm32ii4JEw37wBbNWOmQKdEE7RwYKlOXBBUSwin2Ufd4K0XPTCRpP6P5VOV
Ad5jHpILyv8kQc0un9BqCEQwfSOLySpLeFzxD8xuV3t4GVmmBufd8F0rEkRnchvNvWAPLD1nFVoq
nXU5/V4PgzFOTBOhm8cQvL7a08vfvkBedxPrLMj0blcPDbdLp8dciKSIMLm0ts+S79GvtDYofkNq
HvS03Mdg1TUenkz5H1RBgsC+jdb6c9kKctp2e0lil7MXbY4Vx+gaEVFEEBeckNLu8FiG+C983sMf
xS6BxZKFswrLnTmnCcINiGwxi5LdpX8L6l3WHpXe6WfLRfTWh+TiC8Y4wxt1CrEyOOI2V2ikh8mr
Z4JxVxiyvbDHf2OzYtpUiPHcRKo/yGpyZKbsVFIT+4p7nws6e+139eh/hIGZb/BWTiUhwUn1itnT
O3aPLbcqZaCNrb99HLSm5nBk4ECdDHtul8WJhXNqHI4JZz0S6rH8raKtx/cy2jmPqE2OA5MH+knl
Symm+J36vygvOYAyfcS8I+tKAOf6Id1vRaTlU6fq1hxOsZpJnMbfGmbJHEbHPHXF2h3Y3bqSwRnR
UgJQVeHyPuyjdKKX2RyWQNltatdlZxmUrld35+figZkHNbs81fms7K5943nQnCZkxjQpgCSVbqtV
f+8CDGYWt704kaFS7PV0Ah3UHH3heDfRwzzsaoGc0gWRdzeo7k4M8VMU1ogz6wgz1fAma1Y1a1il
KSH/Pgyp7TIUmXwfzUNqyL8nRA4y/KxTOGYEa5Cv5aA2LDEKE2J6Ku1ilyOVa7ybDJHmz6JRX+PM
Pxn+jNB9tGbN1ZKNXnNnUVNcUp0hWsqzyD7rQh4l0DGyRYDqrvRemnfZsao9GDP4t1w9zeec4zxf
+rHx1pmmbQQVHVUtcgqI52t0b8WrT335Pj+jGsGEOrPn0ffK4Eq3Jk1Qt4Xka+uNWAdO2RRMFKQS
mCn57L2sUoCKAe4feXSi1Bg4LF2BACXjUFXAAKgIkNoA/KRf4Xz5MWb1sEsza/ziGOerKfy8DjG4
4FdupXyDrfbeFmkF20aUAvgKR44lVnQFE+QbsPIpKUl78tebbJsPOyKT5Ex/xE0sFcRHL9LQOx7x
a606vtUDZNPoLj68FVecyq1IXAb/4RYXTSMQ5TOp6MvnWCp4GWIu/CPyFYN2uttCEUD+2HeQqF/m
oKvnbEp9rZK7C/tAWyBIhB7sRyoiGTGpo7rienmlal0EY+QYofu0PC/AgEnphbr1kLdhkmsRzVwz
eOmKIp8LL5s0Og2UYBEz5tzt80c1a0Aq/yMfnxG2qBMR8wIJLTZVAb+0QhX+Ynf02TuczQqS2THX
0f9rMuINhUGnmYGQXO8FGaflFGKLFysgrFG0HrePcMo4JGF11CMdw88MybRQleLsH2tHwLo/uwC0
NHbBW8zYWm4S5p8ioMcQ6ZF0vMlVtTQ+y2MIeH38K7ovNX+mgLEVPk9oA4z4lVUKQs997xwAFL8u
ygHKeMZUjEtJw2PO5vAELJdkuLjU1wuIAdKQ9U4H9dKUGGVzV4lxpd0jcHM80YHpnb8tXd72uNt0
t5Htnab37AIHeA78HlO78T8neyxYKL2ucH5DqKsMLLZ2/+uPoRcX8mRFcR/pFeMeSA0ECnPuTiwc
liS1uyPJZHGvvmePqv4vfPqXlZz4qPiiteIQ+JWsu4cDnf3oKE9l1jt6jb/oIVaxsWYGGu8NK49H
4bgTbd5vGJzOrGcG0jH9mUxeOtd8l+uHCQmpbVF1uKT5pOdpJQ6+hXye/cB1ZgKXBBFt1u2uzkdg
d/PnjW5xxYjxARmOaUO4WZwS3lWA0GyD8WkDY6MhIYXAtBuSbATI6OtV2U9e4B63eK3EfErpzJZw
vnabhzsYgYELUHSJK310dBUsYso86LWn64fBSlDq3m/6sosms/eASHOclTmpifYBmwBMoijGZfzm
aEl3QTN4HwznoJveVo7MMT1G4LsnDZWBRCQdXt0WGIP9d2Zc2osHEOVFqX4fXu72izX9Bb8d+NrI
DDTZa6sFbPZWakre+qM4cIfA15NcJa5Vn9FeAYNTH7pt/ETJ3xCCkbMcB81XYi+9TwFP+4n9M/M8
qdi7TVDqOATkLUNjpAWnW5Y428lfY75m5B2Bp9/1LvfOlKqbsVvBTJy8qS1soL4MWSRcKcw+re58
BKqaTYag02NiJ+cwtMOp2iVGYxl0VKHhpibVK1WS0EEDLUUxRawi6Uq1NClz95241JPqJfhpfvZm
zkseMWfMkje8o1f9IRtMEV/M6Tp9mVKyeTzo3u420qAcquzS8DNmvMcSsNBA1h3wkYIruCM/vLo1
48MN1rjgsUng31jCA7zAE85MyOfAwFFAoBaZdoYZpkVmFsLP5O1YT1y2tvn/l5k4CR4cuLePH+qW
1SgtrbRp1+qIOSjmTxFP9kuvLiKVJNbHF5XK910jw0YeuKuYakHllzz2kYdHjobgWN4lykoy9Drd
To/SFd8FXlHkNNLGp9rzAqSnJY4Ojrk3Ox4/RazFwrJFDbJmPnCkFT6m9fsv4J3mh9KDD1XQFFaI
3+MLOmqdRzvb5GnUP3Dq6ByoeJxon+Rr7dwntMt1Q7ZWwIqYzxQf3W3iDyRWdMA+IZCmT77G/pjd
7lJIEY7uQaoBwJABfN+CLwJJBXBIUiLvVnaHaELFby7i1EkLN0wNOO8/cO9Jiv7ZNp3hTmCJNFIg
UQ19Vm45ejukjao+FIWwqpgP8ylhDOjPeSbdd37UksnXfNqB/vd20/RZem1+72AE1IaSXupWmvK7
DCBk8BDApSOIW4O6ozSFk9EYOTuF31NlZCqatL08LE9QBfU2bMa4PwxUnyAD65vPLK52dewr2PcZ
zlCI0fkG/n6Hq94JuL0AwminZdi54ma5gTgoPBq8W8MiQj/SpokTDzYNvk6Y/rZwrui1zyEwjyOq
q7VBE0WNXsQrcyIqvE9ktsmSEB0uHc5T+lxSFSGbkrU+pER7SL6OaT1WymAS9B17IVJrkXjgjDvN
OTdgVoZo5H1eVXaAxsODU/x5R9flBpRC2W7TLbsiad3t1xCI5m4UPmogjzhq63qgwk1uSWGb0YCL
YgB4i5Dx4meJGC9WPhXHuyOfznvOuDLYGRbS3qzsrKEEl8A8o53i6A7CHrxWwO+81Y/AVqViZrl/
hJAxDYammiBQzU1ghiFufuYnAUIWtUEcmDiEFpPDTM49DVmxkAPUtrfF64jKaWFox0BWX/iDiOCl
RmYvEkE/AfeRAPAl0rnSZzyotDbdNOv3MJrtCcl6slEhVUr7BMRvDqiZ7iXZuIO/WiEn62qwFYSo
C6UhLsFUWL6MoHJRgsaFR7qd7ailVvyfRYvrIbCoU3iyI0VyYb/Tv2agWEFQp4OQ+r+64mNh9yG9
KJepfcAV/NUL0e6cCfp0szf/pd7Omw1y2601/j69u+AFV+v0liRbkEGiJHUYQTK/ZlBeL3ocyjch
iaQOejifYJKXcT4VjK+U9EVLFNAFOp2DI/QQZribAS8twywHbBenQr00A7ezWY+NEwL2+4i/eHnj
jxs6o7Ape+cjQi6rcCJLYgS7fv8bCZbWeDqh9cca7iu+JuGuQmJQbjbENyWGyNpcDOTqInOF0Fd4
r5CbwPowOKzzLEVSdELeGWmHGwQFegX+09LTeqLg+mL4hOMwAKcBoM6NFQKP8omlmlHDyd+A3qeM
FeMuR5FPqiCoO8XESHjH+hPkVJFLpVmxYLPAv+weeY8wOwxricpWjCFVavFLeEuu/Am9A6ZCIM4V
vZDkxz2O7ga++8eA05K5CCl0zG7iok+Y/KPRrbMlwxTGWDM2ex33wT2FLgUYZVnyPUotLrQtYSLZ
/3QsfqWNAgtiLsKFZ6mpMseXe4Wfcuc8LwlhUddjdypgXoGgYLnPNalMXOoFW/PG0rrC/4yqdi0q
umIcX/9nvPKHlTs/+8IxxkT91VfxjhryLoif101AlZiwmuurgjQUPbzlYf3epcFre/9GAjWbhGnQ
B/EuRNcO08iob2tdIV5tbY2KiBrNviZlBvmDK5TxN7LqcFuHN9LCIM68hg1CKDHSl0izWskQUDS7
Up0Beu/929+LZx+ePneyYXvhL4TIiK6biu6wQevlEdjUkzzQBYFSaBoxlMlDsZAmpl6EEfnj78uF
LcbhaOHDX5Op/9ezfIzxLfkr8SKiCVvA2F8gk7XyzpoaElBFLNDkKlmpDIYX/Vxcc0mINkW9IQON
/LV9gc3wORYNoJOY/K3DCxSNR6FvEGGu8klU69Et7N1gM4fg8iUTTk4Wj13Ta2hNeQ1TsTtMlceu
l2lweJpSsk9tIAuURnGKm5EbI1dUsOcNZylk5SvoOnVQVSvCc+ta8RcYaz1TkvMbCD3Of2W8SR5z
Uv3riSyGWBeNxcltfNOkeUtCAZu1DL5lBHntajXYWIm1g4CVQmbn8mwCVCV/3fgB03u0euIpy2i4
IEY2cR2CJLwkQmxV0j6i3DWoywSZWDbb38LIlAhgy/qj334UIzFsEWWYvGxovpryrNl8MwZotxby
4CAPjvtSIx1hmy4LcXXVPe0duJPpi0oSV10hd1HgdBROsn8VDjaOkIoGCxax8SZ/jKIfMkmW4jb5
r2FWul0kZ1G9HKjsvIGgTnlTE4saLTuVT5DJ0b4mZHvlx9rXjTIiX8hsobmXvtUhp4S8HBLmEd/V
/roz1gedD1wEF2M3Qkvp0Hp/UUC+62p7vH9HNaNbU4kwlArtxoz4w/K++9ChceV7/kb9wyLpcHIc
8e5kG8UgGcr75nTNIGxDDqA22Z9B5ApALlPBgkeHVtA2R7tzrb85orwrs8a5p5qzQFNGEEElFRUT
0zDUOePU2tdlObOSSZGsheF4UO/wE5EVN3htEhlC3Wr4AW0QDBKWOHn1bbdG37R4FgKTCVjhAqj5
3jLA323dfgsvjtmk8Xok3bn/4NkNUijX5xKcUlGVMQDrmSXQn/iV5XT2ucZOGXGfsH0CLTrdBpo/
TneOj11Xt9ZZhPXiKcvszKFbKKcwle7dUPdmjynFOPW/iFV8hA1ystS2oDW5bWpboRDN1bWPo740
P0P0pfG4DBxhuICrYxLfeYyTLlvfXTXO5J+5OZatAjWi705SXPV1Dh9Wbdi3iZFlg+CB0IHcQ1+E
TC+3SSrW+cJAmCaKURl2QfPotWzUNBIbrjAuxLBrXTJU7S6euRmgL5owMD6NgcRTUBkPGe5NlDE0
3e1CU6coBw8h1/xhEJzSLqtLmBcecJ1J5uOVa7uC1ApC7tL4HlW5ynP6zrj4qJ/5zq5QTUkV8QcI
F2IrRgeAwg/63X88bjqb3o54CQYxUUuAkToIt0mhfNwkXFIPLVjF3+H4eT1cwHEejitwA67h47dh
JRZ/crfpk6f+3N3F+41unu4qm3E5qf8d+EqX1o41RPBy4pEUa9Xfu6ER+xAYFKIYOkhMqeWH5PPP
7N+TFIg/E2JdlcNJfbg/0UtBTPcq2G0cV/r5hOOWgbK6KcpgwL11citwcHvCY7+jblD90K7MFCzY
Dln0Ffee3FG4Nwy/bVN/T+vnxRLpSEYwUKfIBGVkk0GoMf/lF1Krxc+tDQjjHScYNGcZzf+AT4E0
UUOMNfMV6zoy4l1LGJAfdwDe0ayMr7Lf6k2nwkxboqpHRSqzTrGQB+tszpy8ofkXsZAlEOeaozpn
8mpWIkvHf7KtpwfgehlwST1DVCyvwVswWgqoLtJFzZaLvb25bi6OECQvzi8RIN4Qw5XlxLdqr/a1
ONpw34nt3yh3ZzUQ/EjgUxzJellF3rYBPeuMWJTkM6BtTaorpW2clR6ub0dgSVyPWom6B422qAWh
i4StZoeGB/vaV9ZcpoTLsDaoI+ve7Hwh7wnhTqYO4bBBpys1FyFjQvHgih0o8QB6r9FN3wdH1EH4
q6PMsLyJAfHF4AhRM0rbGVo/KZmkTbSBTO3VkhBCPH3dlQXbyiTutxM7JbXTl01Rb8VSawBRyaa0
ym9K4acl3oT5U29K1QZWhzlbLWJ7yTrbTZ7iH7FM13inJuJluUkikEFhmAbY6rmStAwHJYQRHlWP
fcLapXEOMxMTq5cFO+02ypnRsXy3ZqW2mJjdIXiuGIApo2MEpK/9w07t0sqOKiFZHCIH0TDQGA1J
J1WO51uraEL+1Tmj8Rz/pyZS3xB3cdNsw4I+H8KNk74OqRibbuhFVjmkcNHAGvRz6s0wwN8CAEKX
ziuC/B3vvNs6qIxmoXcULPctXhe/uDRRjTePoVtaknl8QasTTh25X049tXvhZPcuwiT2ULA9TKku
VgFf7RvL85h28ax9KNIEkLN5/7fXzeo2kj7IKliW0F9Qto+Tsrxx4O0BVHnHWavic53JyMPG1yOS
oNhwKhx5YMuKLv5di/0Aeh8ZXD44BQEr/yCLpsKqaUEOQrTJy+sOkbbLbbS1Kyfbat47lHNFKJgd
MGTJRN47Imo0CqEyEFkUn0ZvTGL/UJ5h1qPK9jhUr2fzZarsz1E0Ut1Y4sf79Q8+KgWmEE3IoF2m
PS8wYrqmpjZmzhqk9sc+zpJRBOuLAWynyvH8qPKEqltSTCTGGQiWIRk6cTntizfCiAJZD5E5ZUe1
wXPtjVJYDKqczF/K4Fs=
`protect end_protected
