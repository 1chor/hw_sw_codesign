-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
JTsPEkh0E2V2kQ7ArrdTScB1FfDQYflF3htk9qRBx58J9fy6s/34jedHSpt5tAVH
YWhnoZi6dLXPFjXI6EkPrAU/IBBK52s9qjvgy3/6FBGAk+gCp8o4q/a4I0LRifZe
oxnhCdmmpWHp3C+adPMTZMIPin+3j//6FQMmN5Lsz0w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 89280)
`protect data_block
tety4Qi8LNGSwebx0wRSJwJ68O/RhvNdFrpatS7xumnOLvbX2SB579yM267tf4nn
nApGNml6ESlfjYieHYTkhRNlW2AJfHJmd+cxfidmZ0DO5xUDM1Lcn+pdyw1e15UF
hwMn9VgfeBS5NN9+e/MTKt6YL5FsaJFjbnsX2ifQz9b94sx8PstEeMgX/RGYFU09
NOLWN7exZBuX+R4Wlx9hHk+o6v+Aj1NVPfnJQCiHMV/4Tca/qSgwFv8LjBsouWiq
X0EF4WjOWe+VuSGl2elvojDwGrm7i5ZzODBcCvIV30adx1ciVYyI4OPdXRAlVjmd
RFxTrOHqiJAcSQhFvadD2LX8AxZD5clD+ZtCjjaqMdTMNV6ZT4YVmgQblifSwrcd
iTcFxTn9rKbCu8cMzxfhIwMiUL4hn/PVkRJe7gPCqZbXU+cGnpoKy8hbfPf1MiTr
ybPetceiWxEo9iiHSEdzMH1eiwNiu95T0vo7VaNUaUdIZ3bmpSNFts3PqiEZVjPB
ZUESuRHMWfbETm+M4q1OQao0MGHPxzNZA/pSwyrknArcS3nDCCKSt9bg1RLHZo7y
Cg4xPIWa+qnDj87IumGuSCgF4VmcADyoOuVr1D6lOm6hN1Z1dIK3hnogD+cBNKjF
oZmWNgIZ2wxarkB7Mhlnco0M5/zBR36gBty5WA7WkuKAXGstZGB/onG1B8D1WdXC
iUsAwxzYbHC9kWMTF2v0jHKejqg2dxAY0Isnbdpxkdrj/ZRwjN/Wf+vhFBAx+2tC
qbIhIGmQl1b0XKrW4NSr6khI4gsothB2jM0zgcWDk2lz70T05NJy0iwE1R8NUgYi
O2Fz+DUJ/ssupWy1ZzHhUZil6gr44C9+Gg3Lg7Vg4aO05FGHna/fbxuxac0MqG+c
SN2jfOMpJpYA75/3gLG5YSNEhGHFd7k3MQvdkQRbQpmkkNafpv4nQd8zUXzjjwn+
XxPcGM5ixrVMyim6fgrERR6//TGObPwC6wFsjq1hHEkt2taNGn71TP/cQautRYtg
y7M0fN8kDBIw4aH48nbWdGg7tzEG0MIPMNeDOpWt6nf3mMcE3/jfsGk95ziotUZp
J7VX7VyQAOXjzVsVDOzJhhIrlW8rVjqQHr3e9aakIj0o61SzUfehBm+S/c/9p3ro
AWduDwkQOmU/tghVjM0k+Vr03qFx21I4gYKLly8IpgANmbgQL/9j+Wpr+ZmFCbRD
3j/gHG+Khz2enP33FKxfe+jkOv1ZeVl/FKWxWj2L9LzPXxGnBhUOmKDNXV0RWhpO
EWvWwHNu+hoR6SveEBzTJtgPBBsNTPCWSUJiEYKNHSCgsk+9Z1W/m37NZSQJTNSl
9f/L9nKtFPgy3eTBh2ofVuVLchoAbmYoXhMRnDBfjGUOrZH/GlEc34wXtBLQsTT3
is1CgU5HNGxfHpKr8R7WDfJaM6uonIEu2vvYM7N/r73+31hxZE+rwXIT4sGUbCx3
bKSIiUqPg/Dg/uZtkfVM9xDLyOzWGuY2MmYb6kQw2hiOPsq8u6Hyz4SNUbS1jhb/
WHKhc1vq5PMsgTmX98n57XEcQZqxrTLoerL0x3RhV99GZyTRAzDgvTDzkc/PJD3P
QSpbTV6MGMtohHpN8CsIBeLYUYkCDfUCLCg/90/xMKIcRFrkg+riD0EjnPndfZ1P
DTuWyIxfrfhIpAQCPGsmHuvdpBTxD1775kLgB9wq3PW1r99pL81X8eOkES6SBal7
75TEt4u3NPeVWIprMHZQfArvUd9mTdToHoxclanGWS0E4/nvPzVcyPtADc9xweag
V6LeRH0g6VAn0nSdJIz/mbaNsd9N78B/DeTzupM7G5McnyiFKWy+pmIz39ukZP1/
TNClAoxcRfr6ir9mvRNqpKObnL/InbEqVdEai25LOf2hog426eY3jZiQR9snd9wp
uJIGykxB0Uxj5hr/QLSGkoH5DhlqYtrdz53wmRiUnAV5b7L30JDSFrncAoZgcVYa
wp76ywvaqtFaUem1CN+cPDTSTTqnoL3bN+HvKOs/TKXWyZHbcQp37uBvxywKLdz6
qBRqQIW/JZ8vXVhvGJNndHgoqs1mlFdBZpfwSFe0LpSFh1mnJk7LTOO873r8uaT6
LFxdHvMsywuoXo9+SdZmaLJ+LeL/gY1rKZg5fpectp4W31pkmWomwSVNrTOEK5m/
0agTHIFQwbEpRMGGfrnaBRud9tpdZPfshTCIbow3ykSpXatwrP1g4DUmd16WKW4M
oPfqEcRMBDs5aU93kYPq4jVm6Dyl48yxfAEZAl5RfhfRHUs77bFvIGZqwNHYbPrD
q1GZZ3bGYqd3/cducNsghAxZcmHBKarDu3mmMiX/9/9sR0Bx87zPaMqU4c0OmLke
9F0yo8FQcR5dZuRHk3yNbDeHck3CWC4bKUJV+6MxU+O3javhUbq2Zm09HNeAqgF2
e6ZI8Biqr6mz6nAv3/uhrfemv3ROdaiMw0m8ozCCDSgYSu3jFakz2Gy2b4wEoDuY
bcxC+iAG0jVsWt63JIMNPjmUDYZuEE7ZqWeCmrL5xYTMEpBf7Dh0r7g+S6/ZDESV
4VES8fPOWRprQVk5bo/0x1bN0U04PjXzu0xn665QLrqG9+FU2XoUHKc33T0mFfSw
+CXXhaM7tiDoIyrg/uCV9JBg9HVgL+tMcyXSdG8IqljtsuNst50tzjbOr+tCjehY
AxcMUykLayuvZR7a4c/xMQ14yRIrU9wftqBRtXvbXla26ovZ1vWbDV4KS6CC3H3g
CcTME43AJV5O0U/LNTyOIvEVyDabLu7Qlelcq/wSq3oIlLlyuXfAvAfW5TXinR/r
cSbGX7Cxyrl9yClrluxmGj4RgOQNIEtUTisT7iaK05I1bepqQcAbPuk3jgJLulmv
ah1ijQ75rqLlpVqro5a1doru+0Ql16lMuM4QeQV1o4OC8B0NiyqlMgbiGbbnfNds
y3Vx7qzKm6FWEdkPh/B7WvaVB63cv48qHwyuw37g/hOG17NaIJ2jK+6uRU+NMedC
MCaBwd4ZnLQJtZU0EVX2xSH+V6jTVHK8aUDSuvbx/S6gQqfc5Iv4EkipqP793ryh
zMeQrcpemzAz3QsM7ADLA1wxXITOAGWUSzKLm6rh8BQ8jY6qjGOcaxtTbXNL3GyL
RNWzkDnwRLs+wpz7QeW7kzEkwrfICBeMU6EdNDpk/QQpNZgjjRv0iMDzS/j5rZSL
6WwFlOw9tFjT5e6Yd8SkKpNx9fedFY7R6laDC6dMQph9lKBX+P5GQVays8vZaYQ/
uaBlM66xzTDHucFGiQmcNsLQ1AUqDZosDdW2MXgGJEMwH3loiwueiRC1QvE9MFws
Xal2q8BeS67ms3zBJ9iq1AqUNyYA/WFUmOo0vdQMlkd65j7GdoPeVJIMgdiX6aCK
2Td5OG7ElS/MDULhHs7Y89EqCX3KaUL4DR7XX4mJI/xylEIZK04LDXK9CXHuoipU
YXUg27t8leb9qeiRQIho0M51fM/shxVeaaoUQVBcru/51EJvbyRvVn9VfxNX5aOt
kTMp8meR1E9qxe6Q+T7LFKS6EngVX7mA4v5qbE2U9Nf85iGd5+1qzdF9xZMEcCSp
0lS4ci/Af1lQz41zBs+OqmTEzEkLU1q/s3fQ4T9vX6EiK1MMHDCG1+3qnMU1mjO6
sjhJvaa/Me6AnqLmOHV4lzYFZmiOedITvMPTP8U4Lzo7xz/d0/AmF4eCG6TcBj6j
y99GKOKMdX3d1a+B8pm1nnxAIUsNsLz5XpFKH92IUcH6BWlZghMNvcfRs9StSVLd
0VOXxCFfOFKeZxsso0Un2mMFSnbJ4WMmjeNvBvCfc8JKnZvGz8p7EtipdJWSqFN4
3mgj5wZO5hXtuoPdGjfrBBXQFulmPQU28ldNlEdCllJ6WZn6zgu7vEY1GAPHme97
1rXYefg7rSlzkItD0akFc3+X0MBMKhqCksEmJw/BgUjRJuxk6+6nOuV40ObHf61/
pADuVodJTA4vu+vjmoSSVVXuMivn97HA9lDBeFmQwmmftLdwSWrxMn863aDCIZ1Z
fGp1TPyUI+2Lh/wkOdeE+WYeKiEZ8bubYEsDMnUPqgUsemJ53PK7LCbYKGQknzeH
TFYF5iOTyeJzmI3iNDZ0eZqLcPJJQDyMIpKXh7T86+F6wruFEyT5nto9ow010AOI
NxweO2qdcG13WDxsXQqNMpankZ5jV+TYpbhUNqJpc98ci6meYzsi2TU/c6fkbiI2
MpUqRliPM1IZGM5ScYksVowK4nbBk9xphgzEM+/AYopdzgY+O8Pa64PREWx49po+
bMgAvyGbsN4w8vAjJ7BCg02ye7WaesHrqytFi06eMmvBX1TFg9sgWWnWKYHGSfZ6
Br66DpSiC07rRVPainAPBYtcWgwnVu2YVuGBTfHsJ8bsr365bG2wqmgbGuGXmW95
1lpI+D138Wcq1AXxSc04SrG5fvZ1cc0ZeopMpw5LPjkVYF1PY5mW+gdhKzj7dR0V
3Vw8LW2pZrGCK1knCADlKzTY5oPURGkC7CKdp+um5I4BjuWKSLO1PBc8Ji05s6UX
dYlrjGZ8KMezGoupwYR1MAihGOMTKG+w4LZXZDjS5KloxqdiA5N8bA5yYfZ4f3xa
Zts8tbEPelv4kzmAxFnNQCgW1+xEIqcue7VEWw8iVK++JVlgwNNgbpl8nL/DVOAW
qcSZHTFsZRXpjPmtO1QFBCTktIHJoOrCwJV76ZOdJx+goDX/kfRE7EG3RVEbuP5X
pNAMmjTQHAlMPa2Dk9e357QqrocYz7I43MFgTOIEjrjV8t19FRojxpC6W83mrKYN
z/77CSMQprjeHYJe2QzpT2LfvGAdkmJbybd6AUsmggOcW4onSLISvdDPKd27591a
POvk1qLWY+pP8DZIUmwNMPVKez4dpnP+/BRx/bRlLXeRgHnFSyFVSNIBuZO09fF2
AH+caqZTCm+pkB7kgJRrDoh+qbKUzgoUz+KZ9siSXqijOKN4+cHpQ5Th0ROo5HsX
vY3U1O+R2laaBslVGp+Bz7g7DkQLYvW0mbcQtzvGDONARgstpFrcPVI0+v6yPJkM
qPC4qh6KuBfhcmJAlAkmUlp3wKyK9ytB7FBzJudqAxG+ncDmEcwuboxx2UmvBEum
Wp5/OIQMaNhSBwLtGWmjkcuN34+StOcj9E65JT9wwBOlTy/ZQcnSnQAO/gCr9rLm
0fkwBln7WA32/A8MiBhCge2eQ/rzsksvcLRNeKigasNKMSdLVNR2bnlGXwXMuRjG
vLGgsvG4CnYZGTJ3h/JWO0Hmtjem1zoEenwbNcesDW8xNxZQP3XOciS3alLwVkoj
FrDxDAWgt+yHCFIjkQxesJ0Cs1AAUoH/hMRnwgOxNYydoaKMqMcDk6UY3ZTCPxOx
KfTSSbIKf/6PKixhYmODRqY27qvWIklX7U5/P/1XFFEt5GhfJ6pVOfHZRW8cd/ep
S1uCmZpzVm2D4N8w6N9gUbwX2LK4mPrAIJOjxWtA5mEqWBId/la53imjRLzM5kPF
sfoMTGXxxwDZ4PqwgCukjtUeozCmxiE4HukJGsQZIUCVVV8po26lAZpC6zzavbjD
ykUJa+4iAwWo/Vomqfl6Y0xxV84jhwos5Gm4NUryPPXhoAfrmjC8m9orluDiE0m8
NpnuM99PNWNlgY+bQnDy9O0rGtmEs114yY7mp/qf7YNzzTn4iQhH11jWaKoz5EVC
oWzSe8vRmvpuFEMIo1fV3uzlqsGoRj3nh0Yu7INge5btJyzPVb/jvm+j/6EKqDZv
PuWR3rVeparNsigqF5mf6k7oyfKiwM1+u2aW/TvOgneN8lPQHo76NxKrCpIyzrb+
VHkWCC/waWwu397B089+Tquy9qVS/rXfc8uLDPKhhY+fk9t58H/uXey40kYH3pvB
fDC+TWs3Qc2bDyQManvX+4CGr/htXqita0V/w1jcGdAMIrCJ6srRPRlSztCTfMtn
yhuBZwPiFAuRYx8MeGHNrHwADaervsl31KaWdC2yRDaLEZStXI+Z9qUOvnJ+IxtK
MnUMfzCTdzCS90uMHySv3UCDwhCiPES6Oh2ETvBB6h2WJYtriv+0ANamabyWNHKo
K0BiawicoUVkLwp1UkqenctpcNHzAMdHYbbT+8F7ra8yE0Lt9McQ49+kTW0a/MRb
PuR4BfY638gNXKAjFfkXJ+97z2rnhXfexGYszYQQM3Bv7TXY0Gpe2VF5/5ekJXkf
9f+rQgfrCPq6kHG5ivOFBpeVAERdUXLkyd3g3fat/on49TlIYRBXkZmzZH29K1sH
El/i41Pzhzkpag5ABTzxgBRJVR2vHgbQ5j/7kFET1sFe3Ps+xVui9CNFmwsw325u
zhLqK1A4BANNawxbgLLh4+nCqR3RiOD3qG0K8VOd0ixnHJi/txvP9HiOrePJAaX0
3iTUE/Q63VWpwQLRAebmN0RsjqHeb5ZZDm2MbIw0zq6j3ttTbsdoKzZYocthF2Z/
6kQp0ny4gwIStwKeXQo9mRqpV1P4ul7EXBuq1QOijJEG4p3/VaMUhin4ek1Dbxz/
ApUvwQfO+8I7Ltb+x0YGtSVnJ66q3lhDgfJ0cIrHePEXiV4tltP/7LeCLwkOJ64G
IhHrdrqQYeCk2EYmz4EKxkTvnW/zbfBibrgy2U78rPpldhAiRiT3J4ceZ37byov8
Y5XXG0whFfLSKahvKsXjuxAfD/XX1MRFgg0rKlH/kVlQoTcZ+gL9Vp/EGKQQxRu8
5qGQ2uC00/E0otBmlxy0S5b5PWFhCUjcM4Fzt/fXv5XBgu1lS6Byo727oEh/nf7G
EqMvZBdNCLjoV60JIJdA5N7p/uLmpxXIWi5cYvorRLbkMaHLg4PJryV0+8T5cO+y
M+MXMTbQ21yRHcj2u6tvRBPnhqB+rGa+yPxecO72sNYHvQMQhq9FqWqjEtBiwf5Q
NdKQjo2IYRpGUz69aisAwZ+0FXt3XQb+Hxc2V3GfPElCcbM27SoTu/GfJ0/ctWUB
KnN3Upb7T7aqvvnmvwHlO5p/RzNySIXnBVkxKwevWB51NS/tYUznWXRSkNiZBVbz
QRfNnE67ElZz4nWJJ2HS7dLZxKiaqkO/Oq4In+wad4SFgnXwhaMSgYR0Xr75x2iW
TuC9kK00zy9AWd/FbIES8nCQ7WMlfj/GsPC245d4g7f8ctsvib6y+T55Rx9foZg6
SITGd3sfmTvArZ35wxdpxtHfCYyypEVOwSnl4rCDRhkbjJsRjJjb8VJGCg1iNiMb
vVNTW1sbI9KGQiYZZEsbIrtkSNbtRoCabmsIVDH5jDVL54mL3kG7obzXYfrEyKiz
RyCnEcdp+Gv8W1n441rWOZRUBzLneIeZy5Ll1TEjVwGa2TG8GlFhvtuPbmTjUfbI
CqbxaUY0MoRJc93SJxla/vSYTFwFIJWut/blEyMzi9DTFFJmiKHAS8zZyxsnsbRR
0X9+t0EBYSt6e0v2K1ed6fy0Ey7bwdWmxy+oImlgpluPw/xciwNKgS9G5fbHfrMP
cSD3OS5gNL9vA5+HwBLCHGglKRmVvmM9orN9GlxGpmg1LgHLzCRABGt8CsySQbpa
X6PAlen9/KPEYiwAKONpwVRGgDVvuixFE05JG8imYoQHDM7Yu8y0DAJYjJKijKt/
W+jDRtalmjfYdp/2wu3bsbRN1JL+UrV38881Gy6OvdsCW3o8ZhJwvnQAJIBUuhWi
SZy1PP6sXqpk5sXJr7pbpRftcZRdFwVlg8Mp9zJIgfZDE11RoEdQ8X2kfvSfRsZq
gRnSzzaTp8E+jzd9BUMZaSIJOSvFNU+tYUgMGcfNAWHaDNd1I55zpZca1GugtV7F
HZ3ZEbzFrlC2u+PHI1RYI9X599AUS8gdnOtvNIl31AWZLgIMTkAR79IsnpnX5uyL
25HIDs7ZCSiGjkPjBskYQ1/33msFt92dj2Gl7g7MdzbVRLGopoDI+aSCjQcLiFou
gfRFZvpW7KT5BnEbHQETz4fM5ergiwwv3CqX/+kp7X2gXajUEbwfBSA1jI0uL1Ax
U4xzaNMRmNiDT0U3D0MepL0HPnz/2Jdso8xFJ4Ctzs/aj+sRrKlreUATwzyIYFQL
8/X3RoGN1H9qbkRd44+CTrz+vI90LM5kcIqilzkCFGP7t/PVMX8LyriVS5ZXvk2v
kAetLrlfqVtMF3djhVZPhAbwk4MqbPEdIUeE3i/L0IRUDOEl9lZB2dregD7vTjii
O/8o8t7tnlC4bJ5NaExW44R4pAsAA5ZObWtXZ4aOwammEDZgrvbrcOOq/4/BVS31
eUmPiWytKyOo0JwbFKzDekupF8aHCzDKR74LlnmAumz9f+JFqVYtpjrD9MtkzFID
fjFniQkFpIoRzQhT82LPuTqvU+1Nw+dB3lHiaEd21lwT9HzQENHaA7msS6L/0ycT
m73HT8fdYNOwDVdAg3b5Wbjq/sjCbfnHMm9lK0jTOrQT3LtehU1l5ZQCgOaxllqh
r4VvVy1iNUg2+AaFN+yXiugSVGZdOMC6Kaw4lSne6CDNUZks2q06PhL1ueSp7XPt
CfLo4FNwkpe2APoa+kya3zl8Bq62ClFtMt0lUWsB+/nmJzmS2sI0OKgTwzGx3M2t
rjYEW+IrJKs714d5b+KHfBfZWbR6znjNs6UviLcY16S6tppOuRWNXpLIPlOzEVXw
X/aIyP7S/dD3zKa+6YIXMV+o0v3xcRmoFK/1TSB/aR0x/Z0sq7PjXWu3hHnT4Kwg
zXGFXZw+rI5EJGRvyf8RMxKE2N0S4dq86v0YXzNZFZlUdFbxFoA2MMEC++1iOS7T
BBpAoTm9JScRrcwig2naxQSvB0k8AbiPFg4gU0sVtXTkcGUOO/MW8BwGW7rNV8+s
LuAOhlLIsv3H37dBqc6P+PAjsVLinoJ44Hb7Yod0raMtSBkdj8jftn3MfLEzZ9By
yRR4Yzy+Qam32aGcTH9ld+3xVcRZDpxyUGEJZXpkIImK/x+2J06PMgRMhYONUnW3
STrgTfzDXBedVxjHdXBObFJ5ZK51DiB6iDRju6Ur4CHFf1Jp0C0CY3iRnRZab50s
pNgF8AKuuEgAp5CmDeVjefA6v8wfU30SvDTK9FN+6xvuDe22kPpzJtwRZwJaE6Fm
SpjJVPTaL1/Lpht+B5RCm+NNsJFuH9iE1Kab3XmH9uy+kEWTOLL7Ls2Zc7CJoh0Z
VkQx9Q+Ulfy3mQO4W6A3Zu8VYOgM5V9Mp74yUMI1U5qHrctYznrtW9TMIKC6Msov
me7wtS6itdeuf/SCyPZeaSf1N2ZRHGsIhsXAdhnaQJM5zbvPCRqjGcWooz2HIa+7
syUr556xAOwWbH2tjGJEiBcQpqy1Nt8gFlz6RHKVGWB/8t2E0bVCMwj14yiyLEhr
RrDaJVRnW7I1vkmJUXO0m4BTZULkqGyyJ3lyBnNObPOA5H6qXdDsT4OearOf39F1
c9PF1SbRFE9N5k3MhKxkx/1bb95OU0BLjCWZO+TVgE8OoziIYMUIMVrXf4yHtrPm
ML7w6Ji9NLW6zSToiFNzNOayCGsU3PGtIIK+iLOJ4HoGYeqdTTt0LNvMBKvhoL2X
TzYXEMguk0/ozrWOYJMAgHR7W27o02/bWvC+NbPT935zdsmPGIONfl7zOhi67NGh
23EdRKnN4/CA9z6AXEChjitUfI8g2gcCjkIHjfO3xl4OUPgy8DIJqhDCEntyV4ny
3KsZ3YobVqRv9Kwnr45gtLk/EwOnLPSBInpNCeCg0+ew7SsUH5gcn8GxHMWnbyTJ
gSfMiNCZyNCW0c9x+SiNfbwm073Ud2UMQ+qP/OJN07S/XyPWz/OfWa/HRVSG++MS
QUrNa3jsf0FcVrzFsut3P04HXj3vAlUiOZsGKb5IppwJVEzP1dhuAAfEMtYyaeSP
yCs4vUHFRLYFg9tFJ6akK4BmYmtnyF2C7g5mBmBnMZkOFV140FqHBzQ0F36BxGou
lpX2+OQSWVT5cyWt8+NX1Cu/DPMgkJ3oES9OsQrK/f9n1Sj42ErzMLuuK7F3K6D/
EKmdcv/SA6wptk0BC67/9pEgdKh9AAIxtsKjPKT6TMvkYJW5JWiQxoGRmf5HmGuM
WRqgTIVtgEW70OBTujNNJ23HW+j+uEuSgEapAX1nB7uUDiaOPBBJVitsEDbC8Kk2
E3ZWGziAkktYfNDM6Iu5XviOzAqP0MAP0KFm3b6ljj2Eswt6rS1OxM0B8jIUdbvD
FfuQXfwfe0uiJ5fpNvDEXCfikjsmZcISHAUKghs4d+e0Wp6Jr30nDUeSBqZRhaLi
HsHS2+mDwxkLf+zMTA1ZaGMOuYFqiUABKd8MGR0wRIr2RWApLfRaMGXWWQT2I0Ds
/AM2Baksziug2/TaxKf0xU0xOCAydPf+3LCp9gju3yqONKYnbBhb+EwEkwfFm1i8
1TxzBGEX0xk7d6cW1nv13G7eLrlMgp7alh09jl13oxvrG+F6/iLEr4V9yMTiaONa
PdWOF78FyAooccCe2u0O1mzd5RTtLE4JvoT+TeVghll/fTQJhVyiaFzdfBuGFCcB
FXN3OnauNSlORUXSh9gcNVyixEx5V0jplV4jcHi38Uoh5Tap7M4h5mq6biCNkoQb
xDNaDf/fdSVqp/+bzOe/mZZs0iglCtKuj7tKML6wWKfeLo1umZsLbt6H0YpH+Sxi
tBaVlftZek8kEKmhraKsBbDkf7nzc3MDkbGVG2QinByUAuAtYc4CZrD8FC40H049
As2/Y6IC125b7UXoqMoqr8i0bmoIRiqSSUZ5JFsq/jtlssEnjGCtOKOHgeQxHMn7
r80jfGquUV1YS+XwmsFQrAVPIr+RZGViAUsrpSswks95sLVQ0Xput1636chJwHAo
eWx/Ml6JEODuZROikHcSNypE6+uuloet57EpHIeB3wzA3LrrUOBYZE7LKQ5ztIc1
nqLS2K/YWIGFBlM8gYwodNc+SqUwbr3kXtZxMethzC5q44dVTz424RPJ36xjC/Qw
gHNqRWuRN7g1Prv27fRX1shLia7gsr/ZMoL3SWlsDDb/8R3IyPS8iylfewED1bMQ
bu+TCgH5+nir06bFU4v5YubrqVeApNl9JkZkh5s9Pons0FpOceR1gYqcwKirgPjC
ZurEhnPO7FJVsljkFA8PyOiDwCmNaLCuTYpDRMBM8BBVlnoomiB0m9K5DMrZ0kia
0VizIfTatG2ApFrFBRcGZ+FQE8dH6jad8SBcXoAiY1+8BgllfJNFZ2WCk+ADxNlM
VJUPTj2NvbnZN56LtR7uJSfzn22mAS2UtP9Y76BxczQRBaMWLYzYIGMM/BkFNYDR
V87SrDL9xMnGE8Ojn3DTJCMzKJrLN7R07fv9v4jqdI5hu95QwlymW/sAXR+jvMcq
M5Vcuhb+3tcJVtVglGhPc3AJEmqtgLv2TPo7sytPHpW4hsaOg6oMTt+kdRk4XyAO
zB06jd+nzq4+7OP9MZ8JjhKfjms+Y1g35UzIxq+KOKbJYhJi/UB+AQ1CdZCLhQ/k
0rVXTs+QS1YkKK7IRS/plsG8YU5yoUc+dwyTPq0AN1rX2cfAXopW2+Ou7WYE14PK
Amxv5E26klCyGBD65Y64zj6lSiAFrNW2VIF/hmEeXME8HBKq1pWa1Ior2wrMLgNO
L/9ibPpgL/ES8uNOrApgsiYhaG336mjueefvvXzQyE5MHuHivKzaoz39LPge8OKW
LQmDMAFKj7aebKhoHIO3GsLdHOifaRt3rbSnJfHvg2jB5jlUStXTNfPhbUSf0GEr
TFeZ/CTy8iC52/VcryzGeuh6wtvd/LqD3ubyya338Q/pR6BkQ4aaY4AZQOLEyCTs
zY5kbZcamys06xZYQZIAeXxs6sRhcqpXZHGODQHl4r9gy5Vn+uBTDIDZuFEz+Qip
+Yz4H8ZnPd1ME/WkiLTmfOfbPYh96/VdRrVAqdDC7DaFgsZ9G2RkASOL1wQmNvAO
hY0YeQIkpHXCDeqtKkCUzsgKMS4RwgrmiEcHdMcNKjk7/VyE95/VW8N0bKce2vgR
ChD9u/ZSs8Jgw2gezd6Pt9vZOm+xI+7dNuNTJTt1rc5Jz/GQxP4cykFjM1uWyoKn
gkVvVOGAtJA/tTWAJgBmIeiyGm+CI5svEwrhy5uX7ZQqJiD5di7yjci7o4laqdD5
Nz9tVOQtQuZJxA42FTvPDLGNN2o/SMUQceM6AJNxasGEgL+qiXW0wDUGK3g9Npp9
pzQpGMurNHGU9HLpNv+3TjLeq5M9TlbbRC3Z7bWklQOcwWzDAIjmN5RkbVqEG0j6
6yNupyAscjkKqURdd2l5pWoKjuDY70Uau6ESNUuLmoUQfir2CATQviAdV8OsB63c
O5BXGGWS0IVZ94JnF1x2VI3gjFFyRx5QzyRj6ptp2mhCn8UipLL0JMzOGKhr5KOm
+gQv1prjVZ/bPFFUV9HuzWSW33fb2Xuv8cbPdzADvkxWTnbsNJkn86wZsceanm91
0HHOofmrSG1+IsPISQttD720jJO7gpIYfrxEzuh4C9YortFRHqfocNCiyGZkyR8Z
lQnhel4PdmcInqxFoB0qpwOOSy651KqJWUkVbf1QX9mOjtMu+mztY3MbNe+t3PJE
N+JGCnagy1eVpEWe0cDlyADN4lyM9PEYqzGU/ztRUk1ayrwbnuf+kOtuIxMln1W8
qvn8dk56u+9IS02Om3cMRglRrC/ebHpdJVa2I+NDWNPMIBuWfNp+vd9LYRf2ZVQY
uqcYo5dcL1aX64v+bnqRgHoc0lk9UddmqirJPcRzqqWFccEInjzchbO5Ddj9xhsc
hSLdmot6qGftf3COXoYuFUzNgPVwtskMhcE8RZWZqmp7SHblp711Uf304iyVZ5+T
Xx7A54GIMRJZrpUuEfSqXg8JkxcSxQU/0Hr8Bmq4d9j8PydLjvsHDHSY0dm7rAs/
ZhsgynYL8Aj0FPjATg8RN3PjT6Z1RRJFZFcVKCy5U9fqng5VEw0jCUfiG0vnay+K
S4Ag60jVBjUGox/fa9oxaXCowxKQGIg+fnsYjjIWyPBjJKcw381RPl6YkEbX77go
SdIxg9Q4vpPeXeMomklqjFGVIK941nq/VMJAdptE1142QBzjIg8zWfqTXbTlmuI6
qJzxJ8s7ay1XU5+H9o8qNY+Hv7R57D+TfbAI2pdKIJ+VTv/0KfUKAzIx2swmeYnz
U4xViAqlATTjPYvUb/vDN+Tz8Ob5KaqwHkFk65ufS7HnnDBjYPSUxy9l9U/isXhu
XaWaz+vGH2iUhnmOuI1bomQqRMe0SU3fm53wW9RdSYlM67q29cSVSWE9c4JSTjfF
R6GcVovWC5QkOu6KDBlqgyJ1RUKu+Y6HB4ItxRv+2e1j7Z5FqRM7fjpdYl1Xh/b1
+GNIz4HijMnr2MnliwPuU+yCIOAPxFlwNEiyD6f0EQGoRy5yqXnknsowbDH5MC0i
erkj1RAPmCkKdkUVcGFHh4D6iDCRbOGqjxp1rhegiLNqxJkeT78GOyNH5IJ6OLZM
jtWdyYHsFauyUsvw/ydjy9AkSazu2yk85VQ1KzeM8AqEaSU4wtrdwUFtlnu3cM9d
yGm+yB28LzBT4z14Lbr6aD7uQgXDB9cM8xlhcQMOWrS6oUj1UYpSiARIIJUOXg4y
50T+Y5enaDmSxI19eVyzLpBDZtfq3vJT5Is5FujZBMgINIUnBpeegU3HjNATQt2M
eNrj0R66ThXODwGZiCRTGb/EZC/SBMISRwF4M+Kxab1Xm0G4oWnfIpVqkfboXxEF
VIXcXlv300/cNS/fR51rL8pfdW3NhFBndej6kXdUg6BkSlK90xV5/hLhA8ULhBwi
jXrprQRDyJUwTinJV6P3EcPXvTGqCUyoWJBA2fQFHIDZ8IUEu2BVl9prCbka0IvY
efYvJcROxzy1gvRAamISePeG9LH9wlbh2xYN6fbYnXikB8drou/wsqwa1PtLbqMi
O91U/3kTDz/ZhgGYRYthvbcB2/opOFGi/8APq07k/JuNxEkL6shuXzM27LgNSCMo
0yDNLHAhnteChODXPE+y8KSsen7A5XHw80s5bby0wPXs9Yv1wD2ZwlUOx/KfZECc
/c5IdFBZVuTH+2j/1R7x14LykO0odajft00zdHED3EdjKcPNcP2/MzHQvDi0L5eU
N6U7QQGu95tGOvz8XLNBMC5FBPfMxBUJMCHn39AdxtiE7/0Qh8oiloszdIl1efS3
N3qsZ15zN2iZl5VlmDiMhSW6poFLY7SWuP4q53/2VVunYY2uFrkHAR8YyEXifF7p
xUoGBHSrXurDIMMeVbUrHDHbtA0GMdKoLvHNE08R+AlES8AWZLOHMXirGzoMG2K/
2BWRcdScqrNvSTI5qE9UnZ+3GSOaqEZdGE5fQARhhwsCNjtMnS9CBl0otOa4HzvI
Dm+yXFyKlNub2TF8KyUxh2JFwCMVGccrbIFpJK8r6ze41qLBynKmpL7wwr62ScFU
O1JRX/B7kdrcMXA1UL2y4M97PIa94tjez4wDvYy2giL5UVHTbiamy9OLOCHN+K4/
IPGhF3DCX066apBcoJj1YuuG7V4IaGHruI0/wUiW8yAfPJZ7tRx+MlglUATRRigi
MVrYs+jCd7VEA8lwR1p0q3356GlxQ77e0bEaLVc5REDiq+Tr4ywK9BNwFjhXy72l
uI2xgxooWpMZEFeXC/rmrYcH8DFf45mB0HHzwuki6TmmVm5PxoiCzAPvt1B79kgx
+pwhWQWNZuf3pkotVRvvMd2rzb2ngNx5h7xrecsSFZOZ5YLine5I2unvrqNzEm9F
fSE0m9Bu94AZhQxLiVXq0/qGRwoqdrzlvpmYBwuakn6HSbOOZsia4xNtC6jB7JsV
u8vawbm+7CJaMWHMEHDZwu4yleKbcjcCPh7skQ9RGfF7Z1uyAwgndkPCh5Kq9DcU
tX/sa41WY4iZlhH5YJnXQyUqdSq8YoAWf6eEuFlcZ60CEhuWFO0v7PYR6tg3i1ZT
LyeMZQQTfY6sux5FyNCEY92TI+O1HwWRYIIDLV23Tx+SWYAUDodgQQMZFg0Li4h8
woUuJFJkgHevAjpgCo1YZpD+DFFFW66Ae7tcPtdZJ5Z6C0DR/m4vPJUqV7FaLExc
iIGCWBydVA92P9bsXHKE/H11Vqf7xuQcs5zE5boi2frETmBWoW10wRO1ISJihslM
D8PcTeN6ym59gth7IgmMF0wHqnyOLOguHCac67C/AX1wC3zMSQ2w1cMY45kdyydH
nwk93R5BPOMdFECOnAviWewgKt0mhlUcX9GkerOO/3H0AUKl6Iw7QA45lz380yzX
wUPF385ZOvWcZfNaG0lACnT4mSjrjwgivE3KGfBhMvEmN3YUcKLi447JyTy+dIkU
L1c4xNuRVyeU/vmAEaEfXsoMmDPlMT9kmr/Az1wVcwWENZhrKH8x3SFRWkdmZrs/
Qrj2f+y5VBez9ntnXMXAumOTPoA+Y9aT0d9pp97CefuDw+DNPCMsPADohACyfzps
MQ0yS+37vZQ8QZukP7YSRbEqXpn+4GmPj769qhsJPBky5UUbMUZmDfy8QkX/n8hM
bN61yWaHpqZkV0ESiCe5qtgl5Tqv/5pHhox5GXeA50xtdwbw7PWzFCtHEk4QjY2O
jkoBK1CxVgOxnRWB19YzHGg/KzJWR+eGG9RMz/GiXIxV3cUOyKoJJD4hv67y4g7X
suklttb1/1P4CvCT7boeG7CXlDjqD8A8lRT1FIspOaavm64QFPYKVBQqcXnN0TUX
ffXl1PWe6DTR3siyN/N7hIrUi2FAj4Iv4oHDqIZcRcwp514U6VnXjrk57T6mNkgI
VUrEU4TonNoUfDdAhTOD5zvKuvHsm9aLBziyB8QhxCRgnbCdLwybbbYTMzSoiKtM
czRFJgP6JoSRjcnCZqRj5gJzN3kUF97+YIx47NpjTt/mykbOJ+6Pms9Z7d3SM5Q/
13xWjHVWf6E1BrcBWuctdXQgGiIRsHVwlZVpIZH7V2U4h99EJj+T/mVOf3wsRMhy
DKAW+uvnMsnJifrP9VOZDLGWVfpWV1jjRfW6eCdKkJg5rtdB9EuqNwZ59yK9oTYa
jxGlyGE0t2fDHirXVLpZIPdAoGlRe8ur9NdEFmxAmSH57L6GEQ2RCEVXUfNybvYl
VEqhYLOMvPAXjMfxH/BpL4wZdxCqx7Xu5UvGFqbc/9xStpiFGr8N598LI2arJksi
9qATGGJrLIJPLGAlcfeBVdQZgWS6JMIqWl9oCxtqy8M2LobjCJqF2r4hPIY2UHay
0SmkfkSvAH1U1nu4PO6LKhH8CIrcankxiYyXdvlE+GbuzZSnuqhvOmuC1o7ZisDc
H/vYw+h8hBOKe17JjOpG0KXGYwAf+tYQZm5DupvtPTFnkcreyS2AkkJaUgIZAnGO
naeTS+hoAPNkY9KPjYTCG9XpmPoFun4T+pvsL06NPo2bqMbgCzCNHYS5j0fYsCTe
ffkyUJ08tUrzhsoE0uM2ZU0txj2434HBvc7KZVljBXDNFyQVp86R1d4psiHs76h5
m/obbiG0Qn1EH7f5UFdK3sCQ4Av1ZMotD/w873kRJANjR06BcF58vhOIZtOCi/qK
H7gZ6UX2Bjciul10bayycDpXqGtCIz1M6waykhFQcbFeqdeN5UhP/ImOT213qAQw
HAXbpvQG80MZfg/0zzq8csyzxWr3OeXL0lgrE1YrQbigqbHt+/fJOF7J3KkBxl72
hM3RzBCnNmCYJGW0V0ChqwLyEnZZku+GlIErjKIWK62zbRJ0oN6SZOQA02IauROY
K6dnbV2EU/qcPeYjNbb41T4E8io5PzdRN0H9WuRAW+CJP3YIi1M7kYtZjj1lEvza
udiizGVOjQYN5lgejkHyHf6t5bHdGH+5m6qCYn327IwsoFq8YnstyF6ebu/c+kDy
jTAwq5yuC6hxdjDbhjNGIrWc14gD0YYWYGJfF3HFDrmlsp3lmTmeDZ2dSCqeb9Om
McRL5DHGxWPOOHDsZFVzxIGuM3M0gFw2OcLeWbzt+31CjYhhisl/tdASkZNwgsbM
DK/5ItCddUXjTtZUxSLM7dmzhrDkh7XDLcUzu0yWYv5erE3V5b1IZkQWw01Uflq3
PdDXhHfHQWuzqTzoubt5HPCvWMx228zVRk72f/RYnzHKf+kDs4bNPVOfZhSbpWIC
3wqNrE7yWU5E2RfwgyHHXfIOoxSJkv3TzmCbQDBuLv54xPuUVZX1bUJfeC3CfJjw
oEp1pOtvHPzylHbcidkjK+YfejlBTSbZkPOlRlLojxxNOTTuHWYYlM+bniM2c1rP
8+kmI9ZihMltQUcFzGBCw+6vLhXBjLQwUIK6nl8UO0APo6nYQKH+8Qpj2EctQRUf
g8RMxQNmJMrXKUtk4DgbCRPvc/Av5V7gLlm7WhkwmBkdpmr42pA8NH9cggrzC5qu
xGFnQuwrYBPXpyqWrwDzEJKDxLkMRBmgDxpuIbg7ugsNWrO1UFjhahi9CucoXlxq
wXybfeZwYYPHmaJGwF5jHPM8xHQC7g50JA6mv21WooosCKPV/b9YsyYnG+m1vCla
HntPfVkWXtjTe8wxJ4N3FknDxRQhyvgvsJlSUvxddTYqj38kXKdd4mwuPODhQJWT
8H8MLvBYeOduPT2YOcjHNz5WS76aeq3skKOkLRSdW07vF73r4d1tcBgICyVue8XY
SGWYdSgsiUlNaLUqLpnGeh7ULzSCGPXz06Bv6foLZ9vS41AINDpHV3qIZXWuYUjz
6yUla1eF5bj3I8kkkimp1ItFIaVy7yzd+MJZaYpmx+UxWMvjPRxm2zsWp9TQV8JY
GhPizt9NywC447m6gxYH+K17QaaIf5tZiMWiPen+hkRqmOP3mI92K68wQsZ6Wl+7
f6KktKrAu+LtsdoG/ReCbICiuZeqQGuU8HHQy/m806wfg+rJcjyuBaW0e/6s84ws
yDgRycFqMPIa1i7QDdhsqK10+eJjSezJBdbeyGrqLgY70Bc2/9Q+i+RZUWucNRkU
EJq7kUE0Qfp++dWhH2KTbDV8n+BSzl22MaYph5MV0Z5liRGwd4FIpEIgEXDhdrvi
ON2+VPjlzGvtedfpMLfoHuE0cir8h94/XAMvrv1aWShBLxH1ueS4afc45t69YL57
ntzN+oMu0LCU7HfbI7Cd8suHOFGdH09GRfzZw5nDJxQpoWWdB2vN0+6BiB+q6BKG
OXPFQreRvodA8P/kJACRGaFVjvH9BWjWcex6C9zCs/UWeXdpXtlzPdPnI/kMXJWk
9skxDeC0+4ried2uZfKGjdT+t9Dz4u61Ty6DXKZofh5SQyc2qywq3ijq6hmXd2KM
cvpzyf527LyebSgR4GY684TZrwmKaAkJxJK69L3SNCh0nECu7HBXDawN6r+A+BiS
4ZzM+ayhGeC4zmBriOkKDb4r39c0aPR4ynMqaHsHzK9RASlSDUSqtoi2i6bRvz3I
jhWWjzRkxJrJL4kevDAN6T0TYx/FpbMl9IRt+IG8A6BoHkOKHKy9Makg0Ohjc4qp
x0o6M1W01FewBkiir/7nbCWo4HrTDnya9ENgESwPgYuvRkutB0/7uU1NI1NKifTZ
Lfz0QatWKQ+3rIGbTqf72TpUdxSQmkPBsWPvhkWeBpVp4P4CqzMUMCnolUOb4Q83
aAYJwVjt7Az6G4qaMGE6j+uvEFbutVlBmu3M5OEWqAFLYUnw7zW6bXsHMYv3G4X7
DhwIBTfaIs75hfDYhR+r18EkwpqyrhZ6SFt2v1ZbLm29ADGYMbdZfv8qU8fCyNgu
As70M+V3Gn6Oqb9AI+SIbNT707d5WKKPG8oROGl9djZO5ifrBX1BOMSAGn2sqn7v
iV2aWY+UWyaSOpQZH5kEJyNyWFQ06j0y77sEibjvw3Dm/C/zfbOoK0uTGgzMkvQ1
4FkCRMRB0Y2pDBV7qKukOiFE5bYof7gh90c/0SPW0ATq0BjyOwluiAQiZG6lGGMl
EOsCc5LrDu91fGkJyTTymNv7R7Dx9zCv/ixkfaRjDz1EuwUFeFtXlVx4ZQOux3an
4d487HTLFeWEncNt/YVKvgW08sDv6ssztsNY2vCN3OfqxW6Wyy1oxWuGpwQ2m6WP
64PaChfknzA0Zy34A6+Gj/og5kluIWY+fKJE+07fRupOQZehJN/LAoDunaQ/tq3+
5yAnEcy9R8t5hU00K4RnDSbYvmxhnaSNW+Yoel31JEX3cvTQsnN1cdVXydS/2sAQ
oUxwIpiXBWID3njHeeRAnl18PbN/ujd+//Ti81EoLsV8Bfki/GIk6IMWKYNA1wWW
qkcPtPxkRo5PxSrFZ+q8gt8UjGoua8Xvh/ibYI+V9YQX3or/AI7SAsgEqsK0ewr7
O9NfOZcCxKQ85cHqTfKIlcfQpM4vmjUOCInurRAEt+TU9rnpvbH/CTJ6iRL0zs7I
141kvVxm/Yf1LSAQw4Izf3EO2lwBAP/WiDeMVfsFGmNm87VtVUegYeKIkyHgsXga
xpLb1gr8h7qOGsGiPL72Ai7rBNMjD/76GE/vlXto6cwqOwT6C0cS5RtcTAN5aQN/
aFHqfqtp8KWwJAcMV5jTILLzqtfYbW0SjRf8K989z0FY6dIumkrW+OjXqwWtqj9x
/tZn3nAFiwnAQmr8zxVhwxXyAnWnvCyh5kfOzVcIrP8ib/oVU4rMYq4+0yNc6Zks
fbekl26JQS/DW1yyKJamFQjerQq7QSk0SiY17AuKYGk1Qm3JY7pxL+TeflwZDr6R
joARX7SYsC8LyIG9C9iUX/euWz9zwc5Nqg61+J11zj9vVOJvHEp1hUpB1cHSSnb/
BIZm6GDOEKWKK1oQFKHiv6VtYQS8DiilfZuX0sQ/EkhcqEknIVfpiBCJTTlIZ1s/
lDH7nb7QsnJSLYRoRm/wzIKRU1aENGH1NBPOhkPOxg6fAsk/aj1WBdAT8MDhW8KZ
ROCge1ofT8ssTNDiLhXzJFKjBmpGDJteaVn8E8LpSdRXOf88/6yO2L3ZDmW6crjQ
WWHe54B/jFN86mtOpDoKiy4lShPmW2Zq0hSwDic9Nzi3D8oNt9sxiZ4ApWM9C0lz
W4tCbMp9K1+L/QqK6yhIpE7JISazbcUN9v89IN+ApMQBPJIRvh5VanhHmfqsLMxI
XAb5+8Cv0cj/8t/u+9CLSntaxY2ZB6GWb57KIq0SpD+TB3sMF+jKPLJgFUscNKTe
v9UDiBvl1H2pXoqTrI+IBL1KQiJBD4NNVN4cQifcYaoUiPP6vUIbWm1pYw4R6JSc
EYr7taIYscMJzyTocBfCueQizo/lGaH9w9KnmD1BZwqaQGfm2KHbTxxJGV+iPKrb
KYmqX2WcbsA+AeZLSRTbrjb1xyEB69POPbCBd9tmQMQzl8XBrq4ugYeqD/gbkawx
TevJAqiW6k7Kew6YzZu7z0LUEFiCk2sIoeZiRhyU4vnX9lb2u8SF7nOmIp4A/t0W
CjXvGSHeBSqm3CQgcmHy716awm5feSquIIlBCVGZM80ygIEbmBwGdsREQEWuGfLi
Ow1DqA+z5gynayHc17hOZlUH4s0BilljeFSlX7/0jnI2mtQLyiAp/ol9DORSVVrB
ob3m6GBTGeGW0CegdiSEvKndDrZPQ82vyNXPSBthMhaGFcoIfdzvmYvVJsj8ApcW
MLMizWeAc1Y92ZmY9IUd4BiB8+UawAxoa7tsB7XqFiMGHdefRIfRSy2vpYnFkTUk
A/dznjVZnyC3ILE7g7c9QHiyFdyiKDnZmThT/4lYEvi2n3LInkIiURMqiGR2tNQJ
arj9+oi0s2wC6S0Bl+ubqZUBCUxjkcMwSoYET0EOO72GsovveFXH2KZ09oitzMhC
Zo87yWJvI9HhvXWTtB/RCiNpkuTUTYsBTlSBGQN+N+PzivU4cs0Ggke9bdrbfmqV
4c51Lv458M6AcU7qhcIOZyDhoUXkzeILiS+CErGPMGoQ5oIi8W/iKY+FYAe9NDB3
NyLvZjCRAgyXxvVf1sH2JaHIvA5PGbV7DKwJm+nMYsWBx88AnKv9qc6LqcQJAHNe
gvGD6YHz1eByGcp5fHF+7K900nTsLPamuRgC94Lc5erOmr56p2MDtUU1xzsQUCD0
HGv3hhJFOp414z7+PToLW5FJWc6xUXZC0LKNZbTC21Iff3s8tdopE2FLdjxvIr3R
ZtUGgBVUz/ly5/ERxYXGwbSCaHJ0Z4QkZthUDXxCBHkGYWLrlnZ05k+5a9pqPDSV
NACaOfeLxo1y+JZ9Rtd4GaUp50n9IcRKVmp6UieogeaUyHfwHQrmc5bbfjI1iYzU
n7t5+lLQ31gaVWZ9gyOEqm90stycMsRsTX7rkIDzFJpmZAwx3ErFyCEoCD7l3GZ+
lyHCfsWNF2L9sSPttc2k9BNGHP1+9OWB+/bJCiefARM5wVso2qzPgAGxIFiIlDKK
rrZh/L4GFHqTB/gojZH12a/C7rFuMPYwKINPbNgiI879scsSA5bMQnf3k2/Rpgaa
ZZzqYr2z5iWKoFtQKS8jmnGZyY1t4CYVqwVlzHpL2ajSTDcihqfuVahjptONLpBV
99aIiOmYl8sFkRQExCr2L3a++GGFN3AR91K3VYIieenccw2b12eluZkyNvNnV5AT
bTbO38J1IsKXp/IJngWejf7J0aa9c5kExtuXC5jlF5/ZcpIKTtW8JVk+PIIqGEMN
zwWlaP27pBeOAB9MFT25sagVOiHLgsyufGsuuUNYr6n7funv6JemFQBuLGMmPNEj
E65FtCkaTlr5vVGiMR7or7uB8LiQcvgaBdvdOR99hJ/d9RIYF5YjnNveVWZ2IHSD
ocPRN9X1+leN0lPuVpfTapEZy3oYzU8DUvhztwCXMnX+Yy8p2QPUyQhKb4JBXa9+
GaW8Lb+b5opiM5DUWNkgUaFSNj3HI5Y0GoLKhc3110YikNoSd2DBNXa+bxa/e4//
AaEjh+94qCKa8b0cZ5mpweQhX1VYXQJpO44w/pD0EFqWpaYSFauOjcJZMk8dlo2q
LDML4QG6gw9jOZPYQzUsZ2SEyv1JxxZgY03NGFjd1IVxDg94n+zWTFFzrkuX1Vll
NtJmEKm5bQWtbm3OWvKIARlsTKuzQ8fir8GOwZcpY1YqGETshGiDy29PnPG5IGwN
/OefWXCkQH1zow/REF30Tq/AnSHBH3016Vhfe6DZuQxeyvxZUnvXVvA5o3uHwmzC
DtTWWjXhlQT49Pas1GfjzSDED6DmXKFRRKDrHUVP4GDt6O59YCHJwvE/YWox7PLc
vNI54wg/8TOZS9A3V1OPJav8q84wIzDba8/Dk67Qvfx7j3KZ9Lu4VoGE9N8yoeIz
YwtvJQxviyjzNwRSoYi/j87XnqyKNKOhsKHNNDXOlXaCCeyQM6y58TGLIntYUMQC
wxNVi9XcEygtQVhf/Hr0eBvKpzxrJk8rUbak/IkaybTQt2xAGyFouiNAHlW4mD6d
f1f9j5TPsan0zkTZsUFHK1U9xsN/CK2d3zAUvJx7RgSw/RvoS9y1CTcoWWrlGvZi
dZCMKlhkpgUcySXrcAccR6+QubdAi2Qnn3r+BD1V3YUfBViOajwOK/aPRK0rjRyH
+c7J7xsaIj5yh8+oZwzjjaki/TkXsajACoPMBdPI4N0EwMEgBQNexfCfIqi9LTrG
1yW2+q7ZyOQAUUEPAQwU+mwsIVl8YE09JAAkexNLnEToXft02qHqZkdMPoy/iUm6
i4lEMDbKqJxpIzw+x6B4/B+Dd/TgvIZss3F8qzXt711gGmryVA88pAkGQ3wOVQ1I
5SOiPzr2OA3jcicSqqfc+n6X/8PiLPrfys3e7ytopDD0y8tPS0Ko65H8vpwR+Aso
YSFANaHv4XA1e1UKyfhmfPTHSDv5rO2OcH7bhFAwTiimkgEC79raLCdJrle+8P/G
1wZ4nZl/kR2vzfPaDz6fjLEJBthfuhB3K/lym5z5pgr6fb7bfUJYoa4uA/TCW5Ot
LldCP8AsBWNq6oIk4nbgsPmVl1OpYP3bfLEMWswkgyuQXjasleJnrmb3RUIQIXhS
Lt6cikKMK8kvxZ5yRAM//xtb7SkV1X8wz3EmpSSuuqlkyoOZdCjA02jXiUrP96H2
AtMNBe8i9qWCWoUGw+IOahj3YTdKtKY5fzjkTEsA38Lcqup5pgj6hFvcFsPlj3jp
cthnN1Xm2slGU5XmVJIpD4RTAv7YzJFr04dQ750y6yXJSphpHrZZ01z76wd5C9TX
SDk0MeBg1DB293hf45741X/tIeCNSv8JLiYngcXhJjTzX7827uB8WHBC2oULoQu/
/2mKthWgfrVKP1jDKpI6Hnrq2ze55liJ1yqmmoOO2E0Lx9j92ZVjuiNgHyEHQyrj
YdGJVVn0GLEDVsFbFXxQ0qvKa6cy5RCOx6e119hkVe/cSVcBvHI3Idm+A9XNEIlB
/5bOW+9tamPgPbHkXBpaXTf3fHPwa/3Bf0ztJNq7cQBL7R0SNWzOiyNN70e27xYJ
78YM2D9a3GJ0QZsri9zOk+9BzfslXJf8zYebvpYN/8jhtTGqXgGayReyjJ/g2gFC
XEUG5IiHHbOE99Ib4yVlUg5Gsjz+nnMNtHN0Q8dtGyu4ZoXw4HJ0/EbOf2QO7IuZ
R4VteCOJ5N2ww4oHtJCY0qglk0ZNy0N4ipLNIBf0Q72Qn26wuRzYe5850BUyOiGE
qFACOwKlpFFDFo/cMj/nIxbheERjwLfcr4Iv/XYyrc2+UQ9wSKVjETpPob/vOz9h
JKwoHtaWVJahTZKNekeuITUYNY2UwYpcdCCqTBQzxXQOjpLZ98q4T65z3f70Nqra
PLsTPtBJohqYK1h5BSygndHhnWBaU/Ng5IlBLl28UbEdbNDmag9u/qHW/qcG3nGr
719NhZZFj336pa7CEqE/noSDby4bi5t/IoxLl6t5l/gN3zwDEDs99iJtYUFrvJxi
xMwDwo0YOvit3Fbtxcmb6s0r2SvGONBwxkZR4VddQqYV7iZ+TDtPC0+6Tleve7br
GnbssiGTSFCXg28pj2sxqZHJWufH60Gr5ysmuCiumVG7ul9QEwkPyhrrBITCFGf1
+aQ2BveIx0RGLE15HuRJFYPOnNcdT/QGIk6L4VnONIBO1ATZuvuYUjBPGElleHmM
ukSobZaQ3p451/ehYKargCCiNh4BOMHo/Mtx+6cjvPF0RShUzN5YPa8P79xDctwp
IZJG/XNtiDarVKVAp43Tupietc0DljYE96a0pIBaGT5nlhIJhlfG92lEn0kTGtQo
9YeIeaemLdc328DZMqYPPn36kRWGslgpfBpq+6uRhSMG2oIEEC0qF95KbHPK4d3k
AMQsqHAgArh5Jb8WEvM8ICKXlRbZJ6gicxvc9TP7VbuQcUo8gjKXulrTeMQ+bGYR
cgnpuANRzd/tkfID5a0bjoWwh9h/lCvXjdFu0nAahP+JCZeOEz1XzGwvqKfE0dva
ugI9jN8fiVTpa1MrIzkYQ2zC6QBoQWKlkqaIQc5zm5+7NAX42HOhaCGeSOu1xpcq
J4Rjlx6ahoDCWWlNqd05OPnOxGefPogM37vl51fp2RjJXLEEKBRChNUUWo7LCMgh
iBvfRvq8fp9ObxhfNbEGWwZH320k32bGlLaMu1ok5k3F479riaRLLQDeC6A5zKRp
JNyZfs6NxYPG36uZZAcxM+sRk4fymgNDj4+hIjdSmMBgAMMajDuo2USMasHOlZzC
zCt0wec3/fTYMSUTUbz3WX1Pmx8VSvmVpiB3SH8WUus+hQIV6HiViA56bVozNqmm
Pxf3PqgXcNeG7KWS1Qeq5zN5JdYRtaKl+iXmFMCcQ/pEWzVOiqbmsDs1sTPZ+Gd5
LhhsEqjpfeCoqSOtumpFhNzlfUXGRcn+ACH0KpLpRpBmkeMqm6/vfiKMBz5dbOnp
eDfFOi6kkFayuam7wMLg7qypdGNj62D85P4vLJ0TFwQvPflnckeVj93YHLLUo3ak
AvqdlKjpr4kjILL9zrJOC4ZKIgUF/92yBi0NJcmPP1CjbegHras8JLZJLzNQ/4Ew
78Pu1dabF07NfAp9wE5juZIuiyOBD3JcJ/z1YtacE0FQ1K4Zt/NTKKlCRDV8pqSM
FlmUD1PcEbFmlyGFa1GICJiQ3BdCB4XnAE219yvvzQfSU95F+wsIv9p2O166iFAh
MSkpBYQBzsK21sv0w76d87XVSIq+ughvcZUogmywDpZYl5yCOPVZfh9UQgj2Dz3I
71LaucE6+65UxjmdXzTu51mVuq6+R0mxnYbli2SWr4foE68d7iMGvZJvfaoB05Oy
MKvV+q6wKI+tUKrIy/SB6cN8q94ZdLhpq9Ihob5Vvmq4d42ADY2/9R7BQ6YAIDtt
28MOLQQBtOlC5UTCsLEjpynFjuhdAnoegnn5eyzmM4/fs/vIp2Gvrq2uoidShyDx
TDc6Yfk0mpVCzJw9SH9LxPPvruGqRHzkfM4kCfRnEVcSCXZlvKnSUN5QmjPULWq0
gADhdguutE3OXkPgviCNnWkovT+wGmyODuCYHdm6eSdoUPdmwY6j7d3wzkpqILY7
1tJRl5FEOhK2wUOzrJuXSPb43HoBYmOINtJAJgmE79OlXreyKrJ2TX6Hy5erx+Tn
QVpPrXhQUeMX4j2FZAMYW9CGpMJAwok24xOAXuhrsIFjo4VJmfKYmx83FIP+C+Hm
RjCKavorTOIXGOD3aLneQiOQsWEjLF7mypji8AWxvijfTF0v+5PX9xf9wn6EiBAg
WrgdsrJlZzvmaTjqQAMImtynpY45pGexOT3nApCKAsL8sNP0Ic34fEnQ3OdoDwpu
+/c9lv6WrhfcPQ9PPM3g5oDW+kQEley4zrQitqOJUMzYi5zxWCSpJSElGJv7brGo
8HiACivfnHCSvIx1NEmkNvxoTnQqGzuKnDsSNbzMb66fn9l/BDgHli0xbVOfuMOi
onmz3iPHBtTPsiTKF+XlgFro+hA/ZO8R7ArFUFCniR76G3neByr+Af7cxAom9opi
CBjbZAWpGoSEXb1SZ6AbDFLFh8OmaPoZM11pQjZhj8oB7F9eV51geSlA2IeZQqY+
/fTELLusoAFToP2MoKPmNWchHuwb+EmreNBWTwJKpeIae71/evS19dsAY2st2OrF
0Gviibu1VPZ5Ux6bodYO5c3/XDM2sYoCfYaFb9hp7xgphw243knWXF5l00h+/BKI
2kNlCEu4Twz/l9/iObk9X0RJ59BrMhaR6LbZwmMKJ5nilHz8SDRF0Bk//GaLvrKt
S62ilJT6+97JPEAkHWtiRE8pec7HIUOHjD9eQwumwu5Y+cbouuw0vNYVvTxluBZe
Rnni2qZkAnal/29lMWpCQKIDkeCp5tcHre4xrP7lpJMyHWSVPRQr3eeEfdeyfY9T
NwWlV6QLuCFoN88qIQ9zAuLdGfTlGsDjuto0yChyGtDMzAaSCG01Jx63AMDlIAYK
5M9YDFLDqgLlpIk44+8jTN2B0itJDI6nQC49QmWA/T9nUGOvNX8oTSYqA6VsWAnV
xFuwYAhlzk8bG8X0bOECpHoQ8kp58A3hS19B6NfIUQx4xg81aEpGmG1s+wXDFy4S
u4WaKf+yN6AtNpERhCbcpqKhWU3BwYMrRwGty3C7nHJeoPPr+EmpUvK3YwYZ4yXX
aDko+6TRQnEXxR+oT6ARxfAvuJSngVF3bgq3HYUWksswJ1f89rVMrS9du+yJ4U1q
R1dKA8MC8egMVbjBRCL0P6ygFA7SgNkY7Kpsisg3mthpZDBYW+rfGLjxxhq4dad/
379TAGvtixgTm3+TsO2vOKoGT9mw7q12ttruwUCptifvcm60rZjDjvgKcCFDAd0i
gTjVsGTC//N57o22/vK+BdW3++9Al34VC6PXqVV2BwyXbDsf3Y7iwpN3vfvpu6k4
iWyZ69ru2Iu2+nwvFAnuS5dyefSCeKNEFUiyg2g0Kx0kqFvCiWDtJFInEWb3jW8P
oYaEUTljYcXF3n2sbD4KkJHaPuIEqzqoDQjPbgzSINNRbcqCg29QdFHF5jn0qjVM
F3TgpvSDSdV3cecbyi4WwjrIklzt/M81I5N31nJBc1Wk4vjow189qZ/jjVA8/OrV
JMn5BKpfyzK//dOseQKhldkH4Twk8sO9ut8ORnCQCgiUQEmgLz90NiljQFHa8Scs
AG93bKQfiPg4z++/wEN4xRQOVu6vWtG9iqnPs8+HOm7wpnqs8z4gBSk73e4D1H/y
2ECYr3UPj+KbexeOMHDGyyzNFsAcMzU0FcygMJBgeKOCGBBDWEGKe8s7NYZQ5HWT
TEWM4EW+9BCroqEW958sgPgUoeyqg55gVsLrgIqS66GCvYfpixyuWvScZw49yhvD
rSvuQ0JC+10DxeVYm1xkqR3ygBeagLM6H3WAeJLkrUZMX+LCiktlIi7dNbL2csLa
ZEJEICASEyeahlCAkFytmfvZiiXp9VkhdoxzMOkK4p6NnJMlJvnZ/E3gfRrMe9Ql
wsJsgtH1Mfu1e+iwnKVUwoGifZywvAnXmECSnFHF/XFXqnVf5Lm+TGMIFRcK0KiL
Z+w7FU6fc9BfEHrlQvJc3Z0EXBfRiUNLdM0dhMdLzuuIIbE0f/r0Jbxhr+Jidi0Y
/H//zogXYD4HPEKCARrDM04rmu57VLAMkvB0Mg0fTC4ELgjXmeaKKsBp9uo5mPyy
hQZtYJQEtik8QT1ooZhvCd/OXbAAxcce4Cps7xHJfuoB4gb2o7vTPd3q54tRxw9b
fQRX3Rb4BnsphC+3K+QUTz/8EnZJg9n2IahIaoEnbcVKa3euFMFJUCbeFTwk0/i2
Wt3MS5Wi/jWt7pd5sUrHdQil3v7JIGxiziz9BetlFn/tSSlOF/GCpt3gobiv532/
kRazBtvsVau76pgMPz3tiIDZvvUaeefxEh4PeTekZBHr1kop6ao922erYLjcT79u
NFfViBthy54IqZWGScDb7ZQEVcwiXQL+ec6nWWaAOJfUqNKPOliIGP6c199R0CFh
fMSA3VUDez2aFwTOZmUe+U+fwylVa4RU9bvlAKLWCiomroHWqSiNX8LWt1z6tt6o
6ZdYqKAFD57ACDdoEuYRijDyjjaAh66eeO6ztkz4+xSq86NsnNOsW+8GAGs+5ou2
HtzRtyT1xwHpWVmAZXkT45yePrWCEn8BVl95UH9Hp8idXd+RvpE/4WVH7r1XPxrx
/64ZdGwVw86lyxj2H+I9LdX3/N5hFG84C83AItNI+1Gq5AAdS+yUInaawb2v5L2i
ZsMNB0BeMzkSHhi9IgVoqewvQOt+87dERvZv+5QZDAjtrTFLQ3GUshVRXQuSvubr
c93lq3rk0o+j+MJryzwSMYV2p66/ZrZHhWxnrEJgiSMzFbIEz77pgk0byaXqIDOo
0EZTE83BnnCMB17xi9sZbb+PrZiA1/lhiJWfPU2pZJa438O3kIgKs8YSISAAdIo9
ddKczxPbl+OYyBPYmKFnqFSWcXKxNe4OKaIKp0A9zKveQkq5665UeLiPOJokSUIg
lX/Tgp5PRVHuKQ8BD7UneDYXsM9e/K73GbwJeyGGhwQz3d+ODdpw+uY8dSuMoFNu
Vh1DRoR5oKenKStYd902mK5zaT1UkwhjpfGGrWC63d0A1UJD7fdEjQwT6KRXtGJS
8+uWaKMu8uQh1rEPbTUH7Ht5hOkVn4FMMpbzTziqnV7SSPCsjdaA65wH3Zscs6Gx
hFYbj0G7hq4QJidA+xGTxfHztN/o6mig4+f5gwjwUqI2g8EIp96C0sBdtJ2slT56
1FGt//X/J7PV2zMPzDD93RdWRB1+8f8Q7R/N5xtTw/sM0wmrgqOrwiApbT0VkPiT
OTMBpL0YFDTytntgDBKkNJmbwIROtrbjQQPBW5nl9mt2T8xwY+4/BJMIuFknyIUX
iZKnLWKFgFv+Q+VVT2csqeloKP2Btwhqs+d91kkLJhl12DLmCSU4+Ybti+kPat2K
8DZBJVVx1O0qgDnkXl7JHkuFw1LshDfgFI2xsI/VPhjSTHfQ+empNXAh3szx79Ov
gcjqyIzSos5LLVh8nYJBSzvEY3buEc18Cxpm7gpIv5PJbS1jV83s9rzg+a3uVz+p
zHskQFTs5/dsRmORERr941nP4q8VdeKtPD84qfb7KFq7eIqg0zl3ogYM/KKCoA8H
W6m9Dc1jykVoLr6Sj0ZlKIbEFV6V7c42Ri4yjKPuvimUT0TbyLeGfR8hl1MDC354
T97N5z4Z2lBnScUbVaKsjW/hBqFGfiVXHL3CDSgyPeWs7iVD9pS7YGrvDfLehJ44
bkWVbvN3kqtFf2bI/FOQfXdecMykKliuGVN7x/Mey+l/hr/1cxIhyAbFDPToIV3R
vwfVKmkO2D1mtTCDcimokeguudgZcuMkHKPGQB809EXBOrwwISRPRmbrh7oVSHxt
16v1rUcoSaEcwZIAxoGxNsn8PS0OwzoU4Db4eLZqx0PWyBP7JvYibRljyj5fxEiU
/kd0P7D6bGQaslR9X2RsurzUo6oRkrEVCUXgPUftiKtPrFt7XQU8YxPlclX5pou/
J8IH8q2k2f7Msgh75QXlj/RsF752NP1vKb+cgeAR/tUV8MA0hmOOhdspXBeFlktq
ivl/H4VYw5Am28cK09kIHNeIUhWXnQinUChqoY1/7Wc9fIo3u6UC/KaG8mzbBCn/
Vh76HdHZtU3gvSABH/FEVC9QRSV/IKVsCQXCDWcoVk9NsYIDV18LGqkVgd0ZZ1X8
UH6xnQsEW38BoUdXxJBbPEKGkMBQvzCNrvwP/TpxkuG1g7FWMW35xAB7fbIr8oJr
BMZR9YkBPGQL99YrlKtbKMOm0eSBhrV5rlIuZr/GWzZLIC8KrOyz2rwRts3CtKyL
Aw3gYK6YZCAHNTRl7xwpR31I2AEGIdho8HjaXA9O2HRxykAfD43ha5zeUi34UVAC
ml3RfDLZ7XreK9pS3BGgKuthvob0+M5+XuGgeDUBqoJzTt6CVgZXvv2IWM4DI4ju
vfhCKCc9QHmqS0151JdiBpJYWl0SrILsSD1sG2/U5OX+BPgVy3K3weDHwGM0IvnU
o6j1wuOfFpGtplMV7yq/O2RM+94Ip1stHM3+ryWAI8I/hEkXzMmfZLTHj2emTUSx
ttcM4mq/sAqyWHFaDggjRarTqytMlHuTV/0pA2hH+VKPk9+KkfBfSlmv8b8/ah75
PBKQAKS8Btb9t3+RQuCtJ+VURKzFgqZ5eWa+G3nNq+bHpxSdysNV9Cf1KhT4c+WU
VuxN7sFoYAseHBczDCkapx7PaEqmaOw27giG6MOph4hfSurgLhhNx9U7FuBshlPR
r/+0WW+EETrfF8cqp5T6bc1NZtWeAWD5xbc8RFPfmL5B9MiBSWN/dM5HB3AbobMK
6AHK61wMcOhFIsU0a3Gyzqni4+I0fYh9ghWy9vO2TgAHBFheB0GkvulNYMi9jZ0j
k3rQN/uPJptSEWPoocTwE79TIzR49/QF8A764JUpUwRlGbCOfsNeLSnnn31E9nWP
fHzPO2Xv9UlBf1rKiuFwvAPTaxgVfk3GDwBJ7Ko2zcvesRbpSy6ZZAMmjw8KwroN
xZSMpYNWe3NGPUmWdXxktCPpGEpHv4aKqD5mAsFz//J4BuuvOV9dmpPdVf+qRk+n
s3wnxPh3N82U75YLjyxm+kqoOF5LPTHBeVZow8ASO7HxPGPbkPf8AcLEbkSsD6gO
fZjsoTfteVREAnYtWiXf1EhMJVz/dPE8SakI+Mx9kEMmoFMzDFurRUhld5i6FZZs
sJezaZU1dvC/RH43CgR2tum42MlyKrYo+WVIwGqeDXupUD6tItIhL8BaUnS+yNVR
OobIjvqQNJ1OJl4kbBzN8XGjqA//U2gIBDz0kxH4sGE8VW9YQu+MxHHZva8r5hKB
fY40IpQ4dUhZo6emQfK5KUZt/gaBWDgh7Hwdmuk+Sntzr+LbUpUiYyEh5CFu8jrn
TQGtLEcXrhgzmiDbTbMbvAgbyVrUJKEdFkMp9eWfA914mCV+T3qul0bpV0MqPrvY
t+ah32iADUNAwSmV0qzX5nMfsUj5boFWL89Ez+mhCf4KewYTSXwkPGqtZakoqNi7
Sky9pHU8DITzr8WpkUijaDLOTid1OuNqETNwxgq6gWiQRxjJFgYDNEusjFJwLujF
cn/wLZqZSxGZzqqQIJzl52hp57cNYbNiychr0HUVSu9Cm0UAqYoiOzCjE4RTNWgG
83S0JQGm3W9QJ55UvLLMdE0zfMmLDmzuZmUkC0F++CvjVPL0878PTCliQ3rj+hso
P6S1yA6JTtITJnwnT+36pHLn0x7dExkj04T31nhMazNkUeoxQAqMxr0cVxr/0UEg
kDD5KJwrOxwtkPE90QC1d6EHU7b4OO28R/qmjlg+hVExxsisgdqm1IG1QqzNDrzj
c68I4vEV2baf0mXVrpwWkxrSTyvqlU9b1SP9TrZff/v7Ntf939UDu+/7C+N0rBlY
am2Vg5CHf+Iexx+fE0WAyOd7/Psq7iq5hmFndhLfTNbDoQTlvowLnDs4vuQ/x3VA
FoPZZ3Djh5f8pyxqF4ee3460m7/BRSjD9/0N/62nV9cs0+nHiNOcet0+oUE1gQId
dPcjr9+UrU3ibthaV7tEKe7vVLOoSqPI5COT6coITElA5C86fg7hWbvkrEDi4peG
LpK+K2Og9MjuwZUhi4waOATQoeSw1qmjd+iSUsGdJ3eDTfiV+NbD3xq7cdMl+Swk
DCHTbXUd5uz6h1bdcaqZ9fKNYnWIZwyfHOL/xPQK5bsoFaDYuLpCOVKvjHXj0WL+
AjmOKM2HxMvU5YQhs48W+ZfZzLrdwfHwadI7BWyuKlKMnAzGjVoDnBlcbL2keIoe
6O/pjyw12ZIisukQp04+YabuKuDNvwAZL85Q1my7pyC0/8OGAjN/Lnyyw08Jcb9W
Efi1dSN/kwMQ4FeG4a7KxOpAn4+EIDyGeP3udVFL4YLCNi8N4uEMiVuKuapU9CSK
6e2SHOGyJ5L9nZW+ajrEulFsFDgrOrJ5Uf/ZHrbnO1CX+RfXR3f6N7LICyUAfUvL
iBNdxPBIGhbNHcDii7IfPSe87Hb9E2Rgh+BpFTUSKhOwi9J67+r59bOBVQtUjrW+
YCduWvKVfrmsAk7CR2OIyuf0S8gJmjwC27bFqy5u6bLJe94LZ+uJgBFQH+jdalsy
pgdRkVf0wfB51ytZH3DePJZ27H2JCb1V+MkAIfrdVsyDcPBZ//mRbDgltVFhh9GP
Dz5cDIom4oIqA+WpZk7qoPOXkCOBmi27DcBAyFj7ijjzruZiii2SU5WejISEa9D6
UqGFkjnQx8gjo4OyJmJWv9T1c+xUAbxSBQhWkK8mKubgeET8bCvHVAM8pbOxNNFe
OLX2yoO7DvGoo/qRAlNINZS4mHbAJrVEl2FXjERXbl4l1XMNBhi1F+i4eqjytpyw
i33eFARIbsyyI674MYFFlUscyEid/h5qOU0GOVyXMaRIglzgoS7OapZJidZ8OMmQ
9J9vP2R1UWK12AYOZHJIwjltk2mP8zzLx9VvSItRMK7PKbmqqnoXv5og2Wb1wEzk
n0erXGnVuPXthH31dG1Q4JU5cB/bJXXCuA9BbMsYbVrTn62ie1dO/2xbUi5BTnJO
AtNE7zQLpy77dWX7fVyBJzpE4xFJ/TRFYKTzuAYuabz6/8vklsQy8SJGrtkA61uJ
f5nmQPVkQZivMYdur+BzICsaXat5QwdsZ4eJilY/d0bGCQxw+ueEFj9oSfZ6/HOE
wTaM0Wdwln0gAD1GfKr8ITbK1piakoFBpyPBknjyQoMHCMte1J/BN/tmMiHP//yu
osSFtZK3nTMs8yn7X/2q7/Xgjsrt4YMF7DdXArgYXG7dKiov7lbfseZB944Phs45
QNQRHlYs0URsqRrzyciZ3MuHdhIc9DhcKxzuRe6XDDmD/PhHKWuzQu7e5i6Cvqa1
pukGOUL/UT62R49oEB8/0QE8lhpDUQGxRIPxjGedO/2Unu9BDxOioOrlkGkm73ew
foDqKwsvZS9p5lTmkXnoYR68QDlvmZHK0dRgSUpH2N7Aoew18UScUb1oLsKuaaQK
pwv3/Aj4G0PthRu7mpsYAUodJ5vlHA4uobWsMcqrVKyQRv8pEg59nuMJEhHnBQr0
0Y2xMR3aRkRk2Bu/U3yrGC5ixmZ8EHHz1muw5es6GlvTqd9jtxE6rxN5ypo7ytt2
yIPGOCKrQZDGeqIi/PA1D9u79Rm4HE3QvS4AAYrBsAQHezIqbQYBWnUAPL/PIevR
QhYMFtHKx2o63L43QkePGnsNIlrBuDxo1FicM2xqVxDx33cp2G1D/J/Bj19DuNCU
wiS4To+co73kSSr/nl1hGdCx0Gc+MmIJ75NoHWgKP/hy4jv+MQfZLagvdphUsnN3
EbbWIIbyOAKhgR37eSltR2SvcaXw4yS6mKxpazAdVwGMBhSJKz4GCV9QRsvqY9Rl
zsVh8bwpSP+bg1k9u2Jhq6TFl2GgfVXTjN+ruf3Gl9lf9qVaxXP4xEd7rw1SqL3+
6RHU3hyHYj37qtI+1cEmmeN/33aC/+hpmveeQj3Z1x5f4CejOvLGyqK/hivAzyud
fJWkFEdw8dCXIGCRLy1g9YyqnfKbx7esHGKLBkmsRcxql6k6QOleadk/aBhDC7Ee
mjErMA4Gj9E/gSqiYS598Vy3pYiB2SOZxUGRUZbsJ3KWAGCvXNpHvamYbwiQIMP9
5YRziXpbVhVcSWHGN738ha7eiBMGO0jZOhgC8k8p4vJsqmNRGLiSpgyKLGM1hQDK
U3vre/CDBxwHOuVptVxRbsHP/qVSZPzjgXJaiUEcrXdDZ5s7iz9ejG7NJnRM9xbv
pB0cxd0EHifRBxq73d27tcZSS9e6e3OPWrioPEAr/LOrsEynT06DO2FVKJ1U/oUs
H+JGeK6k5WVeJcEbFEMoX9TsZurYbIn33HgxVjnt9NB8XPgAxyG/WeGUtZwvvpez
0wubUIAc/Bq2VUtQGxgxfssORGGzPxEfJZIq4Q/uCSEJvTGMUwQ4Bd95+6V7gBSO
gnIHaxI9hRfA2lIxxZOi+fNy7QwC8PW8cLGZV5NM1usvdlGsCdEHp+jK3/UndVDo
1s8bO/9Bl6BKJMo8Mr7F8N4/Hzxg46DpsaenW8Zm2qjkyPD5dA2w/SVpzldmzFQz
IAlREzdrWBbC0vxKLMI4XuPs/Rnhd9eMK5XXtdsaMYye6xNpjNPIpYLIKprsTqnD
6BGVsEQEc2PRnh+LU6XOb2VqcFd6NN0eU9q+SmRyKlN11ltmqS7xK4YXUkVi47ro
p+i2pKk+Atyb+nBLunrn/sJ7FMlJk6NRUKp7ag4mrocFwaJwaG+If8Umk9am+D7V
ovptzagcgmQ6rd+aCdL3Gu3JrMai+/HzCv7DUmkNNmhCLgBXjI3MvYUaiE2xZPSm
BE3yPDgmbMXpaFVjz+CU4ta/nZC+TFxsKj1AV3f38ltYOR4F/2UfupXytqYHSLDs
Zi9Vtb1DcyHI5Ou6q76mJcI3oq6skVAHYzTo1p58e2Z/y5ct2zxiRFB1EsYAvRgx
YTa65bz6qPUpubU/B7DCmOUJ9svxi0uCZlft8VsiiP2Pm9Z3mLC/4H8/1UqmJLQT
qHjvYMjmKJbqbDl/PjQhMcnqG8gPGLKZwaKTUjr33f/GFM8ZKyfEGHhaZky4j0On
tZlubnPbvKXiQ8u7yYG/ZYgCPLKB5eYpHxW2BHYmTOq6q9dsdp51iBQQo8uv7nuE
682mAwBA91why4+YNQO+Vc5SPuv0DkteFCok14sCFkHDBfxY2ahNZ2xnsRdo2eAd
UguCZx6qGSAt67Q23BvwEYkbA0Yvrftq78vv4JadzSin7mo2nipUp8H3dpFr5Ymd
wB/3XDEVEn/izegFbyl0PyImjI4PKFAEc571PbcBpHd/kzxwTG4jrNHE1obE/TDE
CJN7fEkgFY5/mLMO3BZL0jA7SLbo/+QUyOqr6E2dJdcbWqnbGkmD5A3RobYCImhd
BXIWbSjHhE6t9GY6oYeP0RVCvrJVrlc7SojsVFRUqOqYco9zyEMYdUAXagmc+icr
ne3wIW9/am1nN+tF58d7MOxaiAU1k/vgXoi6Qz7ou0Fi7I56f1fjXNnB/NxLys6b
ebisgluGD6yiQCUBfvncpmWGI/Nzah8D40164yXFxHKo4dL6SnKZBiJoexlL0rcU
jbo9ruTSSlg52rNAhUAWZ2GqGw085ZiNfQigNednCY8mG3RABOr8eFIEX19CLRqm
kSQmHEHOl15szTz70GcQF3JsHnnkgbFQRbACcBM3qlwR3STo/56Q4ynrziXBCmNf
jbN0bJ12+e2JdiKGnuBJQbltugsXsBrwOhyurTHz6RjQ01IS21kMOp0pQ/21/D4T
gb5dajvkxveMAVwvYhMR/632wvDWGsLasrKL/LbFsAYXB5GPjXlaqsBD5va19q+w
MlX0dKrsh6R/X4pI+QEuFHmiK3bRd1G8iuqickapoGtZCtJRXzjXupHNXBa/VLfP
SnNBFuj5p+ELEmNOnucVdAAktMAtsrPiOoCu1ozLgLYavn6jDw2gyuZMgHAjjRwp
n4iPj4urYtqOTlkgvTXiQUHS5oT7eFIF3GwXo04X/5aTVppRQvfh69O87yhE9hwD
MpNfx3jvUtTP2I8JOdffNhIcGGQb0C9D4HCTcUdi2fXO8CgdcjjMa+hJfL9PAiF9
WulaBfRsptdTlFzAZLsrna9HBa5KyJK+nbqqvj33pvr70Dh+dtvtHG95K1yFy7fo
Iscev8gLpknZcnIvOv3hNw7O69IibrhI0sxXeP2f5IiYfSDWnjLu9RWRk1UBcFq/
Nd1S59OezEGbJY71Hi29eSQLg6lcmyanczPLykl9185x7xaCLlMNY34MLbnxnler
wn+m6u7J/VwM5bsFnWMbyqjxC7TimHxGzFjNS85xxV4z+Gcu3SnXnzd77t6MDPZm
eVdB/qRBD7ntqA5rDWzYQI8gP7+PApa1CM326I/P0NlY5Qql5oekNftaOc1LFDZ1
Qm5dnfcbK6F0wP33jTsoVGaLkxV69BjngJvPpmfbZ0BtDD9qztoMvhKhtJKU/lFU
DY1/3s1Q1WOGEwS9HDdUZhTH2+dDdOeEM1Z32aJhyVRgm7cfNGFkzpW1EWImj59B
CPJR2WxddIIJEoNObIfshLFRDy8Fo1IOFC7re8qzED1v4M03+nmhUP5c6/jQOcYY
1CF9ECLwmF8SvAsk5hJ2TA5OODtq5iK8MsuDZ7zEiHE0+uUs4rgfJXo8msrjHrRo
t6QmQvCvbv+rtS1DalkDbmEP10l8t0g06vICD3Pcha/kuhLnQeXU8afhltGu3GZP
yk44I2FpgtaCHBHGSbVk8Nvamt7ScsTX9NNNT7VxKDL8cvRjyumfpht+Vx/eJ6Ci
hiruOYN8oF4us8hlrPkDlPmE9A0nsmk2dZkluqjv3AzMFl9FAh/0hrI2odbOIzkv
UkK+xxvx8+PWThGgc0kXle5mXb4GAKfGawVwuiH4TgI82lqmWf771ZZMBe00tAbA
rbyos7saG4VCFZArN+hMmqUs8A/5syFh5q7a0FXBwzVhCw5ICiq5a7z4fKKsMvMB
iaAfbhf4xcToohsGDTq3RxyoCtBqhSXn2YRlzY2Pr+HiJ52oS77anZFQoFtQQdjG
sCm1OXgHYrp/xBRgFJBvhE4NoRIJyAluHZsELtd6JLs/T4UVuXgGQj5Wc8CPWXhU
9miMRlcZLRDvZJUeSGONmoos2hjGi93WjMQW6PSjb71dytCf9bLJ22aFuQWYUADx
zXgHYlODsC8zxN5FEPmuQWOiqVN8ismC4NzeqP1I3A/JV86RM8hY/yFpOMeLeEdy
0hy1etWrF0VUxQT9JTFV3jycE2bqiPa+1nQM0VBi35JihkiEKtftiXG2A1nPA17T
ntawXXw/ZMQgyUB0j6++N3Pyc97wR2qZJY3H73hC5Wx2H95FVIDUkqi63t3ot10z
idEr9g9OjB7xozg8Rk3M7fS6nivdJC25vrrcMco7/C+HfuUjUh9SfU70pam4MNSQ
XtNnj69lYnDCWecvVCpYL5kH+3h71X2d0ZU/o/ygBKLoKY7vlNX8EsrgyOESnAWZ
tpW3HeUH9DuI1NfrWeQmYv5YQCetGYrfnbx7BBl0bHIuFtMIAruIuxhti6HYnxGg
2zRj7a4IlbwF7UCvBtNERB54h1ME6fTk7cfWR6HfWw3mhGLrI819fJ7x3trPJy+4
cp09ahcaqnkwYO1/47ZyFh6sBWqZyE1ejO7ZBLldx2arxVVTywIss947zcMSsmY8
21JC1FXW8QVnVPK4xMgclmh2MxC2K9scKra6DEi6nh13n+3GAri5vMuOJc6l+lAU
ulQoNmGJKABVhmURBhQE4QpwNz94CJ6oTEMx/tWPKhDUes2oe/xBT/DmJ0lOsjIX
NO6ACKTb+DP7f7rmLdAN76Jl5k7d72pOYjdyS9KCrzdfkIySOX3jcr75bADM5Kck
Qan0n7yzOdyGW4pz8LKs6vcrPlDbHkqOdglEQj4s3aSs6tge8ouHdSLt/K7qCTsB
sBdyqbSs3+8LKm4rc7liH8QoNXbvr8SpeQT/3DS+PWEyiX2xj5gs5JWHUwwJZaFA
2EmkVTyv7B65WtsVFTNeiUEXGZ/Gy8V37QR82S1VRosdUA5mLUcJNezCUizPruqB
78PWEx1GjUWlzPxpuR4ahGLTwPNvEfVD0aeKi/XgzIxJmjZFHyHL5K3wW22I++3b
X6772cdjE5MFotQK0xfcAvqR6fK41pB+6k/GJaPoKLecPi+V8+kME7Bj9AzyKUkG
zhFOc0Ny6lyaDEckgEzlzf0JJqoPmXJkSAy/LEcu6w/ANfr86k5BTXDV+aqfCYdA
NM5gDr5Ah8QM/PmQHAeIKwCPSdkCuu6x0YKcAAzVthPW9QAoY6CEJM8xfqMWkzOd
xWuZFxEk7FMrmEwYeGPms0dSNmPtqKordLViiIGemjaN2zlCJbsTSdrOFNOMJqOZ
ujMEQ9K53jLSpAlaLiS+3RIe2gw4BfO4idurhbnF7OGzmrpJh2hcKoHb6FK52LE0
d3G+bzThI7CxrlbiYwDJVWVlSFJFbV++gIwL36YY5LEsP0/i/n3+edxcUlfCTl1+
d5UkzWMKsga7dfPRSn+K1jHoCOeMH4vcIPRP7ZWrdLqoGrYkT3m4QjSS4Sgiijoc
rXFrvLNrQ/egui4EtYCY0zT90N6XPzQonICJbvTh66cj0u3emm3KJ8yXu7VBPKlx
XJsiR1ioGKcRet0TrFDajHs37DlwbtTSR2gNoV/QfrIJlyOfYPduParJPvVy/dcN
vajB8M57DQ2ol+QCeheTTu5IbZgPwA7C9u6IjqkX5hT+/4INQED3b7UJxEPXnJRP
rW2EBLJPRcf3gw/u+0zqw4EDeq3BVUbRnjfPIQiYSl6ZKEztPy605AlSz4y6yw1m
PdQYlOQRCVEolJ2Wg28Jk5kbGgORldkhpfdA/jBXzyVcLsnUJTdUlAhiPVpjOlJ7
PzD74W82Bb4REMIhYx8DmPYOZ4eca+b7ZYZ59Dw0d4EFCazUublWmdsD0pxar6LL
rQKlqH9IKb84iXk/lN7/hypDkny/UYhx08zBQ+KMMacLwpJ4PLi1U5jDpanUYAI2
yBMn4aQNxIG5V8OtV3JUhKmKYoX9wqZI6LCIGhDz/cEZ14aqtU3LLUtbnDroicn6
RBoXaoOAXTjoAgHLYwznPXxFdINH0rPtVQQWVqzCGgxRBV02l6x0kTermQJWZb1p
PvB+iqx6LHZOs8jbrlCD3VAL4MgS2w54q3gbM+GjfCw91Qrwr3rSKHBSbuoM5Urh
T23OFmq8LblUa08xLuQZBMKmsxvntnv0DAw5/qifL500tGmHCYq9HJT3VrQh4/nc
xFmIDROOPVnwRTrY3O5PliDC2B+qW3QsDh51+Cvfhhum2oVkMnqRasEoK0Y+bC41
+zOPguimc6uI1jX0FbkEU0uaKy9UNL8W9Hc0b3Jw4yeBfx24Xp46A+YErsr4IqXJ
RlfW/n0KLhdJ/VJy6+LwZss4lW//zT8SJxb1scsCDdUFE41l9r73n04OVBJ5uzeg
ZpJShy1c09R5KqfW5Lvct04OWS3dXU+i4GP75k+z5VnsKplQg6Nw3DRc3icSqjgi
Q6dOkCpH2x1aNnQowh0PzvLB/Wz/BbHfOSsz4lIldG2llFgEbqcCpEo6/4jhrNTH
cuaErAMEOAs4MBnr5+QW4NyLy6MjAdl+b6QM5NeUQNasolWcxtqjYv8BFROzDJrY
LMHLFJ19rxXGyFUHCnD2LeK5OzMpf1Zno/KV1DRKJtElaO7Rf1f1KSZAwkjL+jOY
2tIcbFZmlLbKHRf8csZdf96pfmhdqxrztSfK63ERKdhkZTcBqoL99dAZn9YPPbMp
2a4VlzioCvXaHc9RqSE78vli4GIS8VFDR8p/LUO/2iWB07jhSh363Q/4PUxIb5ll
m1WEaeDKb7i2oC7hjpFRvqoEGu1hsei7dqjH5xNXy3mIs86tqW8u1YgiFkj4VAaI
sOi1opRUzHwy1OJmhuLSse5h14thOHNhpPSbGrp3WWax27xzQHWgxeSPZkos8AsZ
nouxh6X4ApvyXmJtTlrjnM5fIIb/Q6EF4dfDcCQo4GBSTO2X0LH5iQmUzF/PKp9E
pThMQTJmQqnD/Ejbu6eDyZouV2jDStezE90UphHRTJWbGyGI2pN1PTbkxk3jAuJ/
1BOfGpiIazvnipnUPGi/Ldz2egAIqQ8PzZSgWyf1C0CIWSsuZ8RG49NEz2S0d3IK
5OHbJxOA2jCBCDXh9GrELLPy7/c7oosKgoAAgTMAxNh4VFR3ET9p35NwiAl5xIcN
J8WL1KriOkRagUhAOp7V/HLssJnwusdk9ky/3PJfLxl7sMGYZ6NNqeL0dYnItaAD
MggWNUMyHpAT2x2OgwND9y/hOhvFvuTW8/Fq3X2wbZcxBZHXfGd7VOu5nJE023SA
V+VUKB2vTa8Ao9pP8cTzk++K0W/jQzXVlh/Mehcx8V4khiK/4THk15+mRzSQnz7q
YQWcXuX9W5g0z5afzY8jExwbSEZFn9ePrzCRkcvekUtRXEWkDOOr0aWtnUZhpbp2
IZZRfR+WSiKD6lprdtnv4C38x/83ssqXp9rM+hSnTanBB33diQpuGOsAS5HrCEQ/
CueX7qJPmwVx06YRYpWuQ60NmTAS/pHr/DR+IHYN7a6+LN5ZNnIZ0pMWdOmJ2elS
+Lzo7lJdvlJLRMugA6q4WX8QdppZcYOgOZ1pDu2YfTTFaKtiVsKPdL0p+W+Rk7wD
UI2E6OIh8bbb9kfHrpJ34uwM0z+jTL5OV4yLvsWt7y6CEktqt6UNfGoTHLFaYbbI
zxLsOArFzad2F3IzkCfFSj+dFru226SPAWI5ZQKT1JrJ9Y6MD3sV7qJIjBZVmvf6
sR652XzUPEkLyv9eHoYLrGnh+ixsuMEcbkrgt1Epd48qVxuI7CF1oe6zQsyoFcwM
/VgCJGlKKLTyYZNjiI7Mi30C//JUHCFszBachcJvMkKCj7Uy4gvGZEiCfeI1c+2B
YKQdUqFixUPukNPbb0tEVK3y2QlVAYlgN6HTe8FE6n77GM7HEnS5g1MQh6zA6f+i
avBAv00I/yFR6m7mQGmDqjWe1YLYXsdc9aFX1hj2AMbUEIFRl3fIczJ42OH3n4wv
9xYValdNLwytAaOCi2MM5U1EHYyvDpf2kOjJWSEbneaEKPjKDqKQTc+o9yun+BrR
Fft6y2C/Igz4jRJcSMqk602Inx+9wn8dt02bZm6hge0NLOUxD9D1ZJZHZFlUq3od
vuEEs6hXA49lLtErVegECBdorEF9QRxetO8+f5upDYx5s22sVX6lfGp6X6Z12kMZ
0h6pDr86SrLcYwysfOHL84R6eVbztHhPJjhupkoq4LHNBqMXDiP4qFQ1euhzloR3
XPXlGLdR9GmxbeEhKEP6Xwwnf/7gsEH1n+UsIMfkbYaw0SntW7VIzuCkn1Vb3+iX
9jtQ6gAsLZgyv7uAF2oaC36r88UBEP/jLwAV5jox3k6aQLBNmeuau26hoCjUaXdE
YOkz89a+MSc+P9qCJuX1luuHR/AMo1RtAZuH9KoSQcVxvTced1yYomkpAI4yA7YR
4gMb/epbRu9Bmnx7pE97PWd58y1RQbyx2Ixv30RJrX4D912HWZ6hkhup0RgLTneb
7inNZhh5oe+03Jca+H8/8Ait/scGuzlMBfA8+NbQVfxn34eva/SoX/bLZLARns25
7ZKcC3+CmGNU+KQpSGZJybx+nAC2aoeWWE30regltrzUazXIrx7ymHjHvDb6SD44
NgS+kts941QmXdu8oDRPkRsqHU87dEEOTqP8ehFo/P7ZYhy0Nryg6/gvn/oGSs8l
xoxIocJiu5OannE6BGonJEMv71napjfty35Hm+vqIgcRNz18+5j40ouMvHNhG687
XeW2Q/eYiEiKyvfW/+4bjCGUtSSzB1Z55SDUtCMApHAswsBuBKPHnAUENXcoMjAC
RH+zet3a0u4ILPHlpCSCVnudM9TwwJ/AwbJ48Qboh7WIdJYpz3yCREfCAbgbHzFG
buO9Zgf2ZJF1wlnPpLFdROlw66yTjXOGqinNdHg5TgKxIlN4cqc8wh9wMWXbthOI
DOFTn+zpfEl6hweGn1rWMLxu9UzyidhCstbzmx6GpgvtuEfC23ZunT1hS6YVukFH
joKJKceboNy88FMDfCQO9AYd/Xbv/cP/+Kcjp6EpieEsNp+vhg5JU9nr/wO9gP+L
Tv51I26TTUhjbauwMO+Kn7CCb1VZWyltNTiOiigNNAzHBIV7Lk07o80cK313LNpT
Jnb+kMlisHKzE9TBv9sRT7UPTILEBnXfpIeiixHO7PWQ4oryk3bI8pcBLsoVQZ34
XawxGtIl4nkQq/gM/98D6fxmjUstnA7nNtbmunivBaFrj7hFh4QofjMjx9Bx/gp+
tqvfeGW3+hLvZekMoF+Pu1kn6sEWgNIIMgjKt7W+lSNXFC6gj9JlgPDMoA5R4dVa
JZBuxF2x6739vcHBIO8/d9Dhrhe84oMJIJPUtXC71NoBfkVnDo8eqdNbZfbTujX4
Bjally5e6yU4C8PZU5Q/6V6iNpaCOFKhPGag1LUVzcTY/2AzPAS2ELUZxPnoidST
CtGE5nMG4QH2y1mf/7/88S8AWAvSxagP7xlo0iV3PNP3Mp1SMUEBN1AbPDgV6/+F
KGTm4TitW9ppwG7afpfI7WcfgHhu2LdHSBWZri+3CvnYJDDmNcTONj607heC6xOy
qd311vSc6QAnx1+LMA1EJHqOtgQNGyXiwlA8pDv/C0U1otkxM7YIyn06FiA16byh
/i1GTGGHrG7rkkEirvM60q6ZTQA/9Vgp3ZSVqc8Kg6VmnuB7v5f5ppsMYMcrBWd7
zb5kUf4REZV1tiqPgG6BkXPrJJSx3s1Y8Cz49e00nOAqX467T0EyQLiWOG/NyQVk
5BaDiA3dHhNHllfgein8Rf4EkvLBdCTKJgZwI3B4L4LOd3jO2kP/NokGWqvpsGX3
KccVsPDGANQS6uYlEupALzSBtZ8Z1ToIeq6ZhJc23OG5eWSCJBcmW1viFPpEHsYK
avP/dEcpxwswyf1IyKEp92M01GbwZ1GQIsyhnGRvpkvCN7ZpCqfIsXjbLK8zm3XO
ZN8GhtN6+eH+cfL2kHCcAKiMrdxv3jZDrCvl104gH/wIG8MChZq6ZDhoZf0+7rQT
lOfbsK7K0Ts2hk6X/XwAklOUfz5HZp8OU+tyr3EjzMYiPTx7qA8LHgYrIwJzy7K5
5TBYbRQ23lIO9lS16l4HFaapiE8mcKL0CmAgPPStPcUaNKBYscsJyDVnMAhxuOUB
OiVrcpfI1sJZYzHkkum+oxwQcKgmGeQ6HexF9XIi+Wfh9GRstfA2Zuk+thG8z8kI
Rrvh40iQtZlcR8eiKBQkugrNemwa1hGKZeAtQIpBPBRBZklkLPAykwfnpWRUyltl
OcJzwHRmFBsZkAxD342+0a0JPVpig79nfT8jDAN0RfFNxqtjO9OYI2hIB+JfqDhl
Qf7b/+Hz3SkSGaQYI5yO0T5wNw1dPq1GenPrWmSyeJlDGrFT38wKa2tVB0Zninzy
Gy7dYz+suti4eQ401NQAp9KxemDx9a5HlWOdmiTuMeCrMVp5gTHbWFpAmVhp7/PZ
jOvSuJ2Swiv6/SPX2XzsRKVvXIThDvEdNnS3ICT+y2CMmZofJ8qouAsq577yFJRr
uRtyMofZ92Gsf7Cvjm9aquguJZG7bJksh9CurjUfdEbYRbK0A9vI6BY7EmV9Y9JT
O0E4eUKM0pI+8R2ZlCDmApq+nkfK7ipa7tOVLRHYBm2XNG3t4aIfSupMBY+jy4dY
exSp4ekHgAWPGV9H4/8l+PfEnQMU5I8qN2MIxnPLlcz+D8zp0rsK503EsoKGnaMb
5rrXKTbnsvk0VUKCboJj+s1u0NPzLIVHZ8GdH/r20oBqQMjrtg6AhujtnvxqL3hf
yteBC1e6tIJITUqffuT9Og1wlDT4EZWf+vyRiE/S4jW2M68AygsO0RO2GKAuILNd
Bduh5UTkU359DLvBNWpEQAkvglL0MemAX6I/xwOoUlutAc6p7S4PDxPV/oK2eR+x
ccPQhuTjDHqP2NCbYqjsQJyVtFrKQ73YiJp1HLHqpihRwT+2d7brQY4+PHW6kwsF
glmQyfE3p7CXmQRM+SshnrJZOFrxztA89jNMhOkEtiagRMRLX5LJxooI5ome/Pdu
gprzT7sntQJEe4MK71C+caoffadONv9wAKhuagsarIsSxGWgRIAzyeKmdtrstRbk
wkpezscfOb2X5giMEjZL54Cr6G2VO+YCZKW14BzvBS668RPasjSbGFGuYQWJ7r77
wHIz4xxc6nbU4+KGyEUHc1w+RKV/Z4pyfbg2WLCyw4dRz9HjWDhv194Pdwa1ZsaZ
zlknU5ocj7lthgEWSnzfwOY8u8KnMoQSD3ePD+bkv2Na4UkWIQXTX6f4FD0R2qRX
Lhfj4EIc3Ctp3qEie8HHkNjEYaneoO0uQjLQzQY+KDd6UfmCs+y6aXj5vQjkGZ1R
/O17PZMwlBCTBUxjnChUnyGY6fUBcS08DMka1Tn7ovdW4iiokwJzsZLmnCuBI4h2
Plb4oEzaTzArsGEGJi2ASvHC+YaxRbdPlIdk2Nhv9CtI/oSwTM86ITNn/QMbwhAs
JW4GLp5zam/4DiFWg1Gz4pvzcwqGAzBdEmVx9h6XaBSPVRf8/GoknIJbArMcPH0u
TQnOk0c4xnc4E6vmnSRvmvKTTsOIn6U1CHcSN9ksXGRj2exiDwp0cpZgJlEUE8Ec
4VgFkid0C9WUj3VPeLv3kdnKwYrhy+qhWDsQPhzr2u2y8dCE2sSfrMpGby+XpWgf
4kcA4SDjouWrBEYcQ/P81aaUhX+nlqhsL/NZHexxL4S3M4vmA0FgmhA3uekldMc/
4Xp8YzhoC08b6jtSPb97WwAuRPJFDMwpbm+1wkc4F4eOxXCC1V7SriYV53dyXqa2
dXIhjjtYgxZt+9O0HESfUYU5S4ubU9xKuoP8Uxa4yxKQnHVkYQFfM7vY1eZpyx02
uRJDDrpwoZlHYTjWLR7IWNf04ITYC8CD4BR+/zBMo/N2tmZLG/nIw6rws8MDQrnp
hgInsLUMan42cTxr3/aSZ1UrI3V8AVABn6VQHn24pbFIBC+VzEXgGb25Zy0MAb6c
T8X7+T2/9RJ7FvnGzmdBkqBTgu1RHQRgw7dDiwoOdRLCVfVyImFo9F/iHrhJorXo
t2pqO2lbOAzl9VkUl/BCd8+AJisOxEpTym/A3JFrxJ9HEsiWet6eXeemkZ0R0HmT
1KKBp3ZSEWT+M3rX8vwMIGyr7IAlva9iCJIX9CC1QCMvZNI9YVxQDe1wWig3zGzJ
bmDPNSmUILK1HyoEvUxWe303s9dEoe+p5m2XsGyM9m5rnfjkKF6mwgQOwLTPV6I7
eKkx1++CO4SyRWH0dpeb/D1nOiRXeYIXExZPRbMp64mHRGbL06ZtF5+Aj4VSqF6v
oynWgI4kab2VGxUTO55rYTX1bY9syZFHJDvpFsaEsRmjZ6AnPrnplefkTG+12C2L
cZ9T33OFSKOxTlmpqMcf7F3xyjlSJmeDE/KYSbM+6rPnIao3cmr1fkTH4+aZ3DlY
8uUPRcv5bBx6kzsCdUEyHdwVuEdw8B1qCJEWrb0/2MrXI18iZN7nfxy5ANumWaVo
s9Y1kaqMi/CB42p35zDgWUkAyIs0A7JmYF+EQMA4ZCS0DmmNdtk7bkWEM8ALkoX3
+dq2p7fwlBAVLeLsQMJ0sFR6xj2yveUb+vxO+NxBhv+BZhszFthIgIq9Us0rZLhk
DtKHRAqBQftOQuFDYQv2oDo9aW9+Nlcq7YX3N+ZSyK0a6EZqIQeftTTlkcuCARu1
aCHi9rP8od+Y0gqcthZ3IAqdV7YoHseO+tF4KYdauXrmMX1n8ocWSnUn5y/NIJRl
C5dVllRD7LkbgMtAVKmzPIPAMdXs4o8jPlCaF28nCn3nK2R9HNFxvJXnA61w+Hdi
U9dmCjysjFWrJO/qW2tAkObaotuAXGfBUbv4I4H3RBWbI3yH4eHASz3k0XaoUK9E
ifp6f3yz/IrIyzB8R4W3jPQ0utbSaCeCSDuQEJn8NqLnwyn9hjvMAI2K9d3bGmKI
/8SL+ZpO+woZAvxP1SEnqSItdzRbtUYXBw0KD81Pfutd+s77imx9qcDkCu4bfqkZ
Ts6B+r01CcUsZdRLewVrQScvS90JS89Hg6dEiJSvI4BGfmCNaHM3LQEGMImsZ3tc
kLbmCR2pKEjZbRPwK55XXjOkQdN30ZDQDvBTe7oY9h41x/KE24R9p2cfYBh/hRab
fEgfN8YI4pfu2whIGUQ05xN+pnXKkgkSaVw7Pc/1J3J2vHPTbnLp/kqMMXu8fexc
OBYSvHwKtuMPOdXn1FpOZdwUIYfZ1r6MYySDhVeHbJ9SqffhKqmHkgSQDwlEjv5+
AokoXEc9XDPVSyAj3WS0/AxqAVlkoZ1neyZC3ZIriMeZhvOGdt0p5P5EB1k9uAh5
AiZVffYpgJDF3LXTnEJcMLkDFvTkV4+NqTeH2XzbfdKsahPquYq6kZc5dA/ptbyp
MV5uQHiCcxaTTZqHcpvFI/2+Ne0/Xu0afZFwJL60ubU2sQSE7R04jkXMZQE98NQd
2rqqEAbMpX/xnXbqFsN6XmFZDuAEwV1m0FdDFBmU1DYb7rGa2xFA1ZspPNVbkp8s
B5LxJHKK/VNNukmuWSGshXfXVsmXEABoKknonNpuSPUPuXZrd6uQIcTscyj99aNF
THIQkqMh8M7Hl1zL5akXCirA16Olx+CdCpj9lpnGiTf6ANOETyYyr9GgPPi0p8sk
lAfZeOA9NJhSJiYra2YIV0WqQdk3phRGlZn8RbN+AJqiAXoIY1ve4ZqS+qDjtvX6
LMmZ3KROzQ2xvf6nOyYR1wvW7NtG/tjp+6grA3ZOdF+WuYgup1MkdNwunUj4XSem
fWR1NBfoS0RUM3y+p4kXZXagtNIgFPud+JuE1OV2HZslHEnF5GzBQhadFprNS+wa
8Q72jzcerBaMfBlpbI+Sya7Q9bV0dxwC0ndiMpzWTOZzh2F9fRK9fYj7qDA1n7k+
kRMY2GLs/k/3Y6u4pbX3/JyiERmKUyP1ZbWiA2/rW/IlyEnbO73Vg7u6Cp9QpwO3
OrRmB56K82szcSZtSLzYVl1cJklhfcA96MAelMGfvjpMftpbvZ55ivyh+TovcnSs
aT+3SLVu6MuJXaVRI4GysZxtoHTL88M0Nqo5Cg/WRdwjeW2ZCpX+3lEgsp4DPxCw
LelDArJaPf89ynHWcxwd3l6JF7wWZQkHwHKe2FXyUO1D3iAHDSKOFU1XyIu9RopO
d+AIYmq3WMOqv6E5AoTK92+eT5nZ16QHNLoCGPVF14QnJ0XXJFFmxsKYrLQRhWl7
PEfJEOLDH/2XkTQaPWzZzeYw8lTRwiJRG9+7kqsrnefPeKGA3VG7lBY1PQxMwkvr
UlmSislt3B9DIlt2LDkJCLaiyZPJGH681iQAv0DQJxig6VmDOD3nFJNCc0xfbT6Z
TEWLTlzUwP1Z6uUHyJ83agtaej2y4LGp+ilzdbpcKjyu9yzC3cYxfSvgVzr4oI8a
i70t2zrN1dVFsvVvZmOo1qLcz16mkRuE41Rjy3C+1OaRf6goWmnW74OSQr5Dlciw
39gQlpGxlKXO2EsSYc5IrOMGSBhtPAoK07UaUhFj3qRutm4yEKv3kdU6GsBA6Pf6
i3oXKgAuiFKE2ypofdm5bfzvusswQQVvtBH4rJlSPWgojgrtWYZwg8X4HOVfYc9s
spmJ4eKskse9s8nz9BpL4mJiwTFF7oR4lKoxjV9geD6OGlMgWKB28OuSRWAZSbbp
lgH4zC5wZPu4jujdSRdv/5yGA5Ew6T+weBPzJqLE3z+Hcksl/RiaByodYV9keqCG
gRsCu5QGdP8d5MOSV34gJRpEoo5HEblD/xbdVH/wL1sQ3skHu5s/KjnvAZQIevRU
gJs53BYOzRV4q/Ip7s2Qubbd/IiJjZ0HnJqVgDJKxfmBdIuM7i0qmOt1UwLtAww2
uS69UvnBF4hkJLMb3u2UJYN78RjGwDILsFhAddpc6090I2Yat6T0Yr2sM2ACmr8d
b70Vv+nhmx4Kr3G5nJ0VFClg3/lKLhNLo7l6ssE3NSB9WT6geTqmxjMWIOyMGeWw
PuUIehOlwekExFQidMyCq2tPEiRXi/UrXoKtXNLp7t6CiPFD1+ZU8cT+0IRYwmby
pfXzzI5tFea2tbsbjL14rBHpSh4vCzRCi2LUMg4byVxAsac4ElydXuThsw764vyR
bccyk8aKmodROe2pVTfVA3N4rqBeePd7YRYj4aoaUt4RVocgzw3FQHy+Tdd7Mo1H
Fss+0SIYbtD/lfKObet67SagjHBTgElisnvzIVH/rHHpCAl3H/0OEVeon9ejC/mc
QensrHxZOidrSox/fWzOVHC1/TjJZGb0k7eNq2am59k8lyf43pVXEaCOAx3nn589
Y101d2twiLXEJUetnZ58aa2cARsBCeTjCyHMCUIJAsC6yOQTx9qjJoU81TcwGfrb
/w7eZc25GaERQMGBIZze5pAPp3ZrloGxskP9URdaHxseVmktkSAjSZlVP8doTiNz
vUTv9FggULMuZRyWL6KEVzZrACK9Z4Gw6kPqDfdGoqJaWukyY19errGqR/3521J8
5NeEKn1Sh9mfzFswgSmUMKSnbSuSsPsynmE5dJvIfdozRqXjZ43CWomOt+daYvs3
zGLFZ/e0BpfBLAN/yWf/wVNXwk4P9r7w9QcD6rD+VzxGdKPAZ97gAcPbZq14R4h0
fCXYybymZoXuk4MBwYRlqdekDU3CnyxWBhMGTiOx37cKRE5wJO7tmzSKeu9PIfgO
hYW8X0sobJpzGZuBNCtJexUIgZW476UYp++JQ4DvuwngUVxlNfI+WhhfMjgS/PmJ
FB8Nnved/0DRFXMlYSk/XkG/FTxJTRpOddGR5oukS7W3DpPfJ38l9meOvBCs7tv9
2/kyArt8Gd0XugdQcMaJS/RjcILUKn6iI09qdDXbrIuOGcDRq+7GIy0CxVqqiWMY
H/ipgZcfAniwGSYPrZxAO8FYT+k2899FnfubMybit14xvxdLImCgY+mxLcWVB2aq
gilX++/J0LUB2P9cX1bi7PGrt1j5Fnzr/9gF9lId0xmNP5Beu1ZWfPxCtHgthfSy
Oak58GB6bFnTI6keBncqu0nwUVOPPnBrNxBoGSCAQ+dCNWC4yQljeDbx7rjyeANq
Csx/cm6pRQRGDnx0bsELB1zQp9Dms6d0HqUEGGM2sNnO4k9SF6CYZqqpfsZcm4TL
ReP1wUuUWUnqaqnbgrcWnEHvJDEVFvJiR9I1NhAkbMomp5eC0hfSeAZjWjaDRryG
Xl7xI94KkblpiEFLMpVFwnpPI2P4anFVz83UQFDtRSMQqOOboL+Jy8s3hTWV8MCg
1pWa9JoT4jbG4aHKpyJPTHeRwAx1eCDQDM+D4AwkvSugSAGmi9SFu37uJ5KY+mOE
khEtKbOgrSC2ScNi5dvOk+8ttRegINcDPpE2ZaCcy2lHVI0UbRishidzn+19tcfi
MLAJveFgyvXtLT5/zqU8QMlXBPOmacDw35DsUrpalJWk5FZ5AEZb2rFnUGH+CEO6
b8brYU7cVl90AKjTtkUsG1+W0ml0LTcx7UseTWsfL+vfWAKScpxAdDNE6bp+MP5W
BYokDnJR3UxFaDoeRbHGPWO/5udrigWtJnXKvPeBM6CDORxANUkMUXCGVZDZBmDB
o4kNG73QHv+tI5ReW8nzxYx0r4jdKlf/c9yzSNTDkMWnl6Z6rPkNAYkRzGgzB1yW
usUl9rVRquKSTFRjtILvwnzeO5uj6TD5XY6gH57xuJYSHE6ImKIl6sfqPBpHYx5S
9J9FiTMYQ35od85eRgKSGKmfwSd1I7NWtWwYBcaV/0Ky0NBx4ZTEoycW3qO679hG
khETmIVfBC9tRPHJ9r9skJm4jsAmzYIseaf4TZxhxPwUJk+UEhQ+PamAsVAMdise
KuuUBFBVAxuQ5fVxzcuMg9RRHfW6O6rqSiYARu4ro3OW7bOW1hMacuBLRZ0rxi7v
pfr9YtkiB2vhFkHUFBT9vf7bQ37g7eZG9PsrMx5QFkp6sDJSvKHqYu2/3ohFSdxq
YHBoC6mY7zCzhdhOElj9Att8bKCkkNHP7F6SZEgIfvQNa42FxZgkCcACb27Ariz6
auR3MfqD+QRKxgQRLRvcGNA2yCUeDFMfeQo9eVsDVm/mcO1Hp0fsTI6Ow1MuUuWN
4BSxErLq4h/b5DQk/geXjFZAXui6YFIzfxadaL7kzL5OdrU6C86idKXhQMJuth0Y
4qph23vSeQQ9+vmuogvhQCUt3t6ksh9YaYKzYP8nVEtMmdsBbyAZ9Z4z2eaj41g6
AAHy607GaRXFhCHImmCUzgRyt0TpyapaVLHbWtNOjO906gIOfAh9SS7TSdFys+Ai
LlB7r/huPsFyKNtRIsdhP3UYBYJvAHaevzU/H4jnf4Szpf89+6kI+6Y4gNbnk86c
tCXp3FYDEyls7VTDJkZunREto2mrHg7GbqsF+zCsWLg8kmwgzVe/7MkOgqK0dgcv
+qtik0GmKWe3G2KVgwIxhvV23yC2j260wfcPV6XpEWR4qZdlp3i7GOSlniZZB6W+
Sh1IRBC06VlQzb6UgjQsWZ87vweXl73ayovLCAlNR9IhVLR7Hh+xmusAHVK3sxE3
1l4Pzpqtj96YpMeSCuLJqV0eNQ0fBtHWGyqPkuv3uFmugtHi7t+UdO+djplx5LOI
kir3bu4eDp9sMtYZI5ET93HU357EdHRw77i4veHkyG+Ku3mradpLKDFTqPI6a7KE
JqIecPFq2kz9VqWbYxmaq7VsKLQB8nSfeXBZy8zTzUMBtalUGTIM1vchE26FqHC5
RbZrHheoWzQZVjkoC3N6GEH/XQMA4HYwymTD97PTAVQnYiW0bEZUcb2ii16dM+p6
rlcysR8p0wZ2HI6Z9OiaRK8fjzMtjqHVj9CqjiioKsrgyuAFlbsrc/AXZJVL+ila
BYOhABQlkckCyxS1RH5P+1mCla4JMADw7eHgr1x6rq/HZ6eg0gSL6TpJtnwZmhnX
N+fOBFI4UJgEm7PwhnXSmY4yLn53tdWsbHVy4FTDLDNvU7N0SGyOIEGODAUXzoi2
uiQyLf+idDHQkwSE7SFZJogkj0tbaFGpSKbPMn2ds3joqcq/DesOVTdMiJ1THvl0
UsGMTdis//G0ux1xupE8KbnqFqBddSdJuMp+hkvCKgXGrvwg3HFGErsV3jYBmP1S
fLpMC/64hr6X9ATU2vhiHmKRjNfgagmvs6IYtXVFT0ZZjwEwrH6x5rwTXlDBbE6V
OxtC1M5hDPdyoY8NRxxfHNroxaO6J6tc4W/qX9Pmut1F41lZMqshA+yPwEVyi1CG
F9SE8+lg++tL0hm2B2RVO7U5LAy9n7ECh03DPsGsPO19A81qTJRcqbKy4TMJmCAJ
64NinqDANmPwGXb/hbMOtklvu+yJhKrBxeAznt4ONck4bXqlrTon7blbUZbhp9wL
ZeT+s7WgMJWazLnYnL1JffQ+9lqOPRA0RrmeGkD2G9NOqtEwKKbGCWfYJpxHypG5
+2YmFmu8igiMNR8R6+r8H2ZUfvOc6eVixe7faPDWnguxEDbPFpxsBArkF0sHll1D
jRdAxTBKsMgaGGN1oahUNkZRQuyzRlHVG/K2QQI6UU4xB0vYABoOr3+DNOkPguJK
wD/aX7NqQ7rh1sScRjbvpQtZ3s7b1DcHLtr5OgKJjHkeTf4KjAzPDjv87G5TIemx
X4kbAg7CBGscqeUcrM2kzIEVW0DNxkMJILrm2i+gn0lWJNk6hz9P5WHdDr1wRF+t
W4p+Ub5yT+Jb5diDTbK1liOrtrZfcmGUx2nN2g0cAOpwHEjMNMygrvShivmZ2g/R
hAkSg5DQtwhxBmVpo8PU7PKgxKH3dBzKpnW2maHjCaq3EwbQFIip+7d20WxoAEmQ
2W0Vxqs4LBcrhnfmOWAfwjKhLlXcNrbtB20qDXVM8Ay3nHCR6w51TXmPcdk/prT8
PAUGPQqVhWzAr5cgXofzDn2zxgH2qa6rVsTMKN0LQeIamVGNgp2WyZYgLfz9JIcm
Ivvt6C+9BQnLV2YcrQF2bADQJ7HsZrKu20qcC2aY0pv+aCK2c2B6D4rLIxSf27oI
OuyL1FXPA6ogBnEjlUKtnkjUKvW9wGII6u9tXtg/pIOTrXFrO9itz2xlyQeRdiw6
Sid4LCxkgwRdj/Zu0nRcmFbuxnLkhxE6asBUhxo6Bj3jww3QTXDSmYKDlqnbi1xi
81xG2fwhyEA7bqjuqLww9rAkn/DsL7keGeJSad9ePMZ/dBCpcibf5nt4fgP0wUi/
ayHYL4qBNL/PIxcIDXC113wg5taspgtHDY9CEON6eHsa932gGFw9c1FAUuLPbgN2
uXJbVTg4/ZqsLHZ08VM7zDVMwj63EPh8TbYBGySEzxVjlbQj1sA6hrvU1ux3VRSA
IYopm7aqAb5NbbXGxpOa7irbcTQChcr9AucIzsZvG5HpNGfo31kAXjAxaSaKtuUW
mTlndDXI8Yjsw4ulOIW2/5RJrwbOqf1br7oQ/M+U0e8VvptULrBZJ9Weq1F4IWYU
vyf5CfcjJy/saQMJ1UNGdBWQfELXfwWSDtan19LjqjwufxX3zmYbPpD7wFXJTj6q
KF+WiGjBQEv6qEklEwF650zo5309SHrJh87nXiHe3Xu/z6NXvBSKvzusKjsR2M3r
goJze0EtbF40NJjJOaHQtKawbo1XRiQBxpgk0c+5+GG7nc4pkdeZvNV51UGicTwW
scApt8UpuUIEoMtfAkt0zqXHk5GmHNob3MJiMAtamICfkvZSWV8pACK+Dy1QmIdU
vlunoOZpT04QmK+t6IkLbjI8Eji66MMhO6cQcvj54Mw1f4mQOGwOtW5bZ5+SjKdb
UCm5/kQ6JXOYpQQ3uec6EAJJE8VcWD60jqsGS97pahLj7BhBn+As5eWTvSnxIB5N
/plDl5AswX9/nEwmKMhPvypNwON8i5Mi/JPIIfDrs0kjd/EFIUA9OyB97Xvmbrg2
RYcTPyxelvFEoE4MJHVV4rvYmC38+AL1vWRF16Vf3ewkVAaQu5v1h4nJByL1GtGt
LsfEGWPlm2gbAdmKDEnSfjJCQwDFYEPlUxzJ9PUg6ntgS1FHk7tZApnNSMqBTXR9
ogP33TqlTJOtEcaaBeLUeAwJ8TjPaNJcZbrsx8WAiIcMBxi7l2LA6ipMPqvqHiIn
5QKvYd6u27h8mnD4SllALj1bVlkUK6DktaCAk1T58e7rgjRvJEshkEbKjSEvIQFY
/qQeZrvj0kBmQmPv48TbOQo1ODc6fYzop/4aTdkHqpOXRjuGHuPhonw0P49LO1ZH
62VfwN3ymlxevigr5a+CGfBNpdEHAnkyYc8hzOxYs5SXbj/DQR+sWYy6wECTE6wJ
CPgCohHJUswi4dACuf42QBgf8FYiPBwUBQC81VO3gAwWfo0bHSTlG/1U4LLOkeCI
V2ko5WOihzyK5bAoTwHa4URwiek7h6hJicFB+upgxAc+GLpsUWciWr0bICc6WkIh
+9NNWxxCY/avoH32NdZhCcbhnX1g7qy79k60my/O0VttppePhZasG0vJawiE7xLe
a35mNoz8eNWpdVEWMagvhRYVrJhx9RaBzLvkpN5Z4ctV9iyrwO2CaqQWNm9DKid0
L9P9pCHoTTWd1huttPcnflSx1WXdckXg+jGemA9LG/BWjJwxemKbsDUMkpcS63c7
T7nHoLftS/aNn/uNdjUDvqjMRl6ve+N2ZOW7H/fEVEg46YwT/W1kAcB+Ve1IyIAX
BNEfwOU2L7DNZVuYr5pyWLR2mGjbW+VKbNhdwY3yVZWeW69VSuVy9m/hPXiKiJ1Y
6jxvmDVd+UMcP/rLhm+rW+2T1Xc95ljrnBfMS18cDpB3dAGrqc8g1fJGmu/aP19c
QdOren5AVk71gCd4v1R+PEmYMMEkdj70Df9U7/mHvbpcoAOPuAHICYcwJ2xqNaMw
xS7vnrRYLw6j+arjApLoqcYtWAj6WNiyIVmlbXYGdzk9he2qYrWlCP2gThAHHLTt
rjw+aWhK2scY+NmanjG7LQupYYuCH6JxjKxCT01l7DhVN8xJqygxHDXCFfnvdGmF
4veJhT0fMWk0/dZDwXsVatmGSxfdSEMleJ0U9rUnRd3Pq4ao42u1aoPHGcwnCASm
1VzG2IAdOZ0bFS3Z0pJEucPXwIBf3brk9C0l543wMu5TMnkdLGSnWWK6zvcuJ4+3
0ao4gctPgw6rz6Bim9zz0AzcSnSXvCP4Ex/cWoZY1UQKz2hhfAA3alUKAGeM9Dvh
ztYnNXCSchDVTeEHGVtGEGYQkHV+IWLdzqTN2HJV9R1wue5ab3+iP42t9G9Rm59z
qkzwhLYqbRh7pK0KFb1CCBsEJhM7HDVrtnJo8OC6yxUZa6xxicjMAS8Djd3Mj8h6
BOXQ9/NCdn8sOl5FSLNv5sVFHfElm9wDhTUMPphdo/4gh/Qmx/REiLrRA2fs/kYm
WXdnp996bh+WciUmF7Jylj3A6D5RRjNYIPfEHrVMEt62LT8l9g8R51GFYZTr5b4J
VfE+p/ol9C4E90k1x2L8Zmg2NeH/Zmoarpmg7Yd5T/ID6kqp4fGMw2oI8fdaEhln
F1kKysBulfeSvUTleDbRTIIe4PBDjpVClhiaxxEvo33SvOFHgUH+94ppU4xejb1g
MOXvh+bJm4caSqRu+T1iPlPn12a4oDOp+o9AUcKV6ZjuPJy1FcuABx+U3Siscahg
nO2hV7DaMMNRN8BtV/px5qiVx1E9OCLZ5T49JR8L2hqLZfsDSoXlnpmYVYB+aeKv
phnVMW6AjDX42NW+0QMA47vtEy9PL1JYOGiK6PwEoYFXAHp7MtxB2J3/fPGJpdOS
Jh6KA2bOmWPFeh+lMhXT8S+HIFL9hGpbRYssQBYjBHtgVIQ7sGI0csdNlPka8rS1
mwWaqxKVR+OblECFM/r8TY7SAmqSWh9zzNZvldct/MtH7nCpvV4rzEyHrTyAxzhe
fd/zR6g1Yhllyvdzdc6RXbnncXDbKkONzgNQ4r0vdIck/PseqMlr/f2o+t/jwJM8
9y/2RJK6uhz16QVPSsJqlC63VhsB3Tl0FKRQCCDgsHtxw6qfq+t40SH3YqAarqnn
ALnEX5x14oUhGB+1DtkqH3IbTs/Hd5dWoj0b1JkGJanY3F9l2mDhCKyMnrtkWPTA
VLLUhBAIqgznJ/tzKGvOdbrtgfG0AMzqqjhMbZklXSz4akqk4YXhTsSqr0nLPWsx
vz35lQDCXTecLYI9JvCuRunDa87FevBLDBMbjpkaCACyjcW7FwRvUEPJyvqu3Quv
+RGn52dsEfUTeBcpH+JrTzU/nOhPsmPCwL85diX4vreSaViK+tu5vxj/9j6thZyD
9gV6wF5ne4hMXfRqSDitaF/+4OFoDXBcJ/NdED1OiI3Bp4k7tqwzY0pDaSJEbFxF
EotZbCSIXV9DMH+UDh0rgePWB6GbfzouXj3pL7Tfp4tfqo69BchsNjYkHWhZQSqn
Kwb8pU6S5VPHxdwoU3TOljRN4WZG35ctsNLmYh6iOXoJw7it1KtklLxby1Kqk95f
4OQeVwpedhHH0tiPC0XzeLREmqFqTfYxcoXTlHsexMo5d8+VXnksVnpvrkleHnG1
/oBy4TF6G7RKZRwYzjIjLrK8q3BB97mpjgcL+lgAvmu+AKZzBeCBoprx2k/mGitK
sWk7R5foMHCLkxkAlJJSOjx4ItSktm2o05TQhA/JvT0nYNQYDRhLmALaDfTiPBJT
Phvj4V1gW5lgS5/xXmzPaYs3f8hSu8is+lInXLGATw8/uI/WEPw51xdK9BvH7gDr
6Hp463sNBU3qT2MDXwnFZaCnZN4fwDHIMIgn3HOi63Dd2CZzPpmk5I8bffqAfIfW
Bn9ugoJkGei5WjxJlK6ShW8xcYX+KWAoSJhj20TcJ7JYEF6SYev6ynh+fqKuXQgF
1365emXE4gGXKIrqzjM+Gs7tYG8MKNwQ8jilB1pVeHHN0Ia6JCUevV57akDwoexx
OK4WvBsf5vBN/h4Igam6ob27PygY9Ti7V2teEx6CD16NMT0z31jTbMdChFTptds4
9U307SQ3hH9Xd90yDIeCk/CEJ2vGQx9NT7hnOQ7gE77E0T6EQpCN0L/SI6UHHn6x
nnkCa2OgMIOaLecho72xihEHcijA/UfD3zRUnW9Oa9OQZFNAi+pKFC0TlHS4qy/d
XAG9KdZmhM4Wj+0UPibrcgl+/lhb5LDiEELxVfbYme/A4bNCod6nlNWdxNRPhIkT
AZ12ynpPl40fB7e2GkvR6BAGmYcS3p0rtHbJTAZEccmpM/CdSKT1eTehO4p0RCa0
Slaawax1073sfOCowOWavvUpoEpM7heXUPf7V8w652iQaxZpIBEo11IoHdDOo6Pn
SJg/5IfljAlXpsfm2WLpuufBzmLwQal6CanK3Fv59leODrn19nCTW59sC5wsBCbt
sEzkjmB560wPoHow9qmQkw3mqWOG5rNkzK4Fs3jVJqcs2QKlb4N3mUepN4VbUovm
cUfWjjrmVloYBGXEz73AyDEkbkVK/isczfuxW5MAoNqztjkYac+aHAEoZTzFvrQE
yYwTanoJlddh+ZNeG5eT1qkmxj0vFlwFCNhhZrnJEauVz/jj6lFRF8I+AROKsVWT
cBAoZfiEhl+1G9ZjWHZI+o3FMFUFCO6SpLzNOoRdcbp+/zaVK5MJXV7DeB4nQfmq
KLBvq0A6IiIx2fwtIjI3Yn2o4Rs82bAK1u7npDr/4NvYckN9zbcF8l3Xq5ovomC/
7XSnZnOMt/K/D7oREbFeNqDNLlnjXFSO1fTfpqCDcvHzcRvFSI+SMb8vbISbw3mZ
DfzJrqPYfITdOOr+eoJCZzyuHNOAjeR9qWzbhY8V5F6WMooK3OkmKvTYj+S/zYk3
PycYKCRr7Kevq3XrCVz6z1Dr2EeriU5ERU/T7yjuMr42VfS4GCZkRwXDxnma+g/f
WmHSYUNp6UzF8l3DoWqhC/dRzIAqHrGhbmaMd26Yv3hO5G3lHKNCMwseEuBjMfuw
xnpnF03rvQ2hctvMxRdQZqGxcEiWiowg4XO900dvw/TdLsh8k83zYAUZNxJfc+Mp
RSpysF0fzJpBZ21A0YDDymuuJfMP7vCIE3l3zlIhc2//Jpu7z/7oBRC8n/RsCFcl
E4ouHeuLfqclWeuWtNpN/IQqylP1msgBJ7MCQjZEHfavy8HovfBWG4tSzTIbVu7B
FaCvM/GwMgRZ7fnvI9zAWHE3HzkMLPmgU2VYXTbdUTHAE7liq8/4yK36gbKDY2O3
pgQpaOvjjbw61GQ+lDvfzaXuh67MxJNT4zwqPX727bszOa6pO+7XY929o24/qyTz
8CXEN4MODXIFGzWm6vrg9fcAZkS4YXgWDiDUNo/rleZL9ZkveOuMkfjJgwJ+cpA/
hzokjqU/I724tktynWZQqzSw444PsIqm5Q4zrfX3JeODPfCjelXxF/IsEo7BdxIH
MmdKPS/jqTPkbLuhjBePC6x/q0wSM9Da6X8PfS8tX+1a0LoYU3a1B0+j2brBulm0
cLMqoJBjc9Ogp9N7Xx1xG/AtIftgpdmgslLe+W1kXxdT1IPXkdCPbKnyzsYhKJCk
c6ekGFIG6K+ZWUMdktkmig3RAiymgsLKUMohXsy1nXfYV6psJacJpqbxdJiPjGy+
5fkxfsXUSrucUcL6rdWfrUeNlziiHycmgEq291wb25w66M+KCI3QjPj55q7UdGS4
cEthgSuEntPOT/dj/45N4EphD7Qh9eoOY3xmUrSq3qEGQpg45s4IOMAC2ebQqUmE
cEzRWKPEpRi7O+JeQSHYbSfd6bhF2CukwW/951zygRe6ucDLU9QO3tb3RVHCnaHP
pkJJGD8qbGeBMBgn8LSBfiPTI4ZrOfn4njxRxnPHchGki5EwNNZY/2rS6RgQJs3H
7oYXaoPsKEkyIQ2KgTbccLcx2Mxm0apBnPxGFM9LW9528VZnd2Bv6mIcydpXkxto
gSnR6oLfvG7H3Rd4eGfOcKjBLmQLJHagEIMR0J1H53A3OGz6gr+QOtKShf+tyQrE
HbbdgzCAG9LZsrmFqw3Wc/ByP2qmgCS5Qm+Mf37zkn9uKRmPJLAPGCSO3Xaw/1Pc
O/CEiEpTzwDiZzAft2tdnJGIkzZopy2rGRCZ7WCQ8vkawxiXWTqydFfko+Cgz0sD
ldQOSvfndYTRnY+XjM+xauarba42pk1TFVll0SJm0Q3gDuKq9jrVgqp8DT3izd21
Noi5fezTVbIHthd05BXQ8S630f/0peDFMbT7Zd+YyksLtxcxGoMsVCrns3JbRb22
LOknz5yk+NyNynF3qgPQoXFT3qwZi/gia9qUI0T+GXeThMIruZB7loj4x4HNdqJf
lh/LfY6hk6fYoag84/68dRrpHmP7uVqyWZGGyxDGGFs4UbEFZaY3gDVLC+xFjQpu
geFf7lD7QKAQp7vqVDjRdIHEfcLF+vUod2feQ8mn1BstluBA8f77nRp9qe+IfBYZ
QLYACUWBDNRmQhlMwsOVH8tgaiDLGKoGeI1iYh/4Kt/Mv/xjKIBG+jBTsmNChPPo
g4WG0pUOLPKAVYMc4/xfx228JeT3NWVtK4DSv7tGzVSy943qOFuxO9nZDcBDz+co
i8zv8whfMQbtIC5IBkOZ4Dkhs4ZSvQPG+9wYS1gxHopxYRlv6bkhAcs2GmeDlsCM
SN3N/62GwBX4dtxWzfW4uOzZqGu0k4DL2X2XrPag5PhsX/hMuZplobNIyrkHE+PS
UL9Csbs3jLmfiZ8N8Auiyg9S6Kd2L8pL1zAXvPSQU5pR2m6Vi2mP963i0mEQFP+a
GjQAlvarryIXP22z4aA97v550IKzO7tIsFBwApaXkl0+rfRif1Dw/gEPrxg5ftEH
UMTIqL9qHl1AqYVQuahC+85sO5KIIWb5sXoPOF43hPVR93WWG2ly/54p8Tdb5DsF
mDU0QrwOP2sODmUscqTG9L/2vA4b++YwwxpJd6dLWygntZLAzeiydsaqve70CUYL
Ve1E3K0S/Fm/hG+Bvn3GC3nyjATMeRG0UFVg0oxfxkyI4mlZp3lfpCYXB5brWsUa
hkRcquTrlKl23FIUwOALOc5+sPFbKzd7tXIfnLi3wzC3298Pdb7P5LSJDF3WF8Il
j3d2at+Sr1n4Y6Pinm23BhX+w6C0gYM8Jny9yfuWRzpGwrNctT7jIMs5CaxwLSPx
CSkIO+xSqL9LLylyfGNJxa0aCioxuv4mb96uvsB6r7LZBWcp4QL7BnBENA26B1sc
mZVDTCSceX3GkKoYP6sXGPtPgGQbghGBfK+MRdiUTixDlCOe96gbLVWhFmFZ3bwA
riEpsB1AverfZHOAnSlVWnKINL/fZzTkaSNfHLL73vEUyn1wREqvPl54n+xtyecf
UlY9B1NH7YVFkHCLOHhIZ+TH8Oc5+BZbyab30qFSvP5ZcdL+g5+PqNtOZAFixI+Z
BChr5OUI8Cu0dx1MDZicNdJEysGHGzqESl6iYgh2VnhJbeK+Yge+NrTglAsaoedt
C3iG27WuuJA40/tbal6xj2qS994t5TN/BDMrsaW9qR6kPlJYMRM9cYjpwtqz2yTr
Omq6tePhEmJ1g7GKsNNzo1jfPBEvgDTf0hOmScdsert+Gyx4Cree3RrUjrMYME36
pfcRPW4i+OmCtofXMnwTOgHhXvfll5L9pF7N0GK4OP4CUwj1GNRWV9NIjYQ11KU7
kVbJqCblBDpiJln2asJZCIyfPNIeKafH1QoKUGjQCSGFJhLds9yShq0u4RveKArt
TJqaJsDW/KD38hf1VcV+al09MZ9I48Eu3dozdRU63WuRwy4dCUFIXAKrx2kJyH/j
f5isZKxGLhJOZKDHx6Qta4CzP4KNLbv2BmCMIRHUi3495NxbSExGB3xyr8e4ZXhu
ohNPV9b1YTTaDGHpENz0V3f777GFVnA+q7QvdVFIKG0AYIfjoucuIlQrHjrmxWWQ
54tKkvRV/JpJR3S6tCvyEG3AT23i6XddeajsIcNUXBP4zcHJ6/MCWs7UVTsewdCI
xqyA0VvPBK2p5N4U3D/yNdX6g71hlPquNbba2/9wIrzT8HKmGYDOPMlNptyrWRXS
s8K3AhCCOLp9HyYQhPrP/Mj8MRd6Er7ZAfkgIHtyXYzPGQCeyy784WaYBe6VMgJZ
SkwCUCAml0F39UXAkwLtDJiPm1AU/yTABraIw6YKklEKYD6Sf6k2+ZXbngXc6KmJ
/PUtU5ZQEoYS4SLoZihRifqR/HM4NMInEzXAaUewZE5eSD+KTvUmmCjfOaaQaXVA
DO/XHt9TOhIknbeFbpiZNMfolE+DnktROmthTlJygHjuu/3z6rLhkJ/VEF5dWlAV
s9++3iR5Pn0yHxTaaMFRT8HaFLuP/0cQZD82NYOm02YGHgqqJRx2RA9yoDqbZ2+i
iVkDKXmVVrv7M/7rFXd9J8M8xEo7jo6fT0On6zcWcqjfqtI83GkBVQ5nCiWjBwB+
8odPC/06G5djX7Ikuf5xr1PZhUoytCYAZznZMSIrbVnFLavxjpAyRRnEJYzaFbWr
Kw5ZhvDX4dFi3/kHD8+VPb7fcS6ss6z2xq5ctZETbaKwkkytDsauS5o71Y89ieIp
DbKqxX7HY1DwOfM9IsiecTOxDR90PMIvZ4Sns6clwPb+howNy0dWYAQpXkWn1/LQ
rRxAdoG0Wv44fNRspmqM7OyDcSE7yuW5MO13R004t7Z1gpaai+kHf98rskdmJIfb
f4IYMBtTxwSxVzL5b4qxdykWods+QkGvr2PQKNEZRhags4gQtTs91MEvYxK/xyjI
u0dadcuAZ/HuneV5dRKMMDhkiL6fI1px46lljFuQTUWhUzk1p9VknGztgemP8bel
IgTSiRReyVQJfDPTsSgJP1NV4wY3R9ZPpNJJU6THJ9LUnVp2f2LVBvvhy7LxHkEZ
47+D06hLPrSaZ7fWw4pSakGqpMoCeV3uevUejBTT+OnpxvFdE2XI0EBcSW8U8lXZ
cyW6dLyNLx4icWkfzRgNPrNV2LW8Lsvyl32z6T+VB635yHlL8nOiI/BTaEDiyBx6
7r7Q47Q1gliaNnmR68PgXUspCEsNPKtB6KQHYJNGf2gsKzcUC7zIDpjaYE74M+kL
QgMfSGV5ZLRnuXkMAVeomolQDsx028Iz0qvOppMlREyTAnz+zmgYvft1flMPyoMZ
c5DAnm1MZs/VqCvlRG9gQA1kYPOwJgfPuh6iY3KkG1T/TrCMorAfuouCoMccLlPM
PiLJGLG1Pd3c7/V1vGuyoB3rKfGDyliFRrpQTV0hSWND9aJ8hf/9mIIeBQVFd36B
vmFc6WpgJDPGBftAlqKcTcXRXNo/HEyBXrdtDhDvoA/+Kv3hdX1gA4D332DMFq4+
Y71OceYQFAOv8xcFTTbVA/Awetp78CMjMrsX4R/ZiiioDxLKv5EQozhx4CdzeTEF
qun9rQvijt5+i8h7IEv4ijj1GOJxWIcovptGDOFjDsBxrJw8kr9er8rWw/GtFUuf
UXPYqSqldDH4rMxHE81SuRvCrz4FTIw47vdsLHyTqvAZ5mw48fvdKxLByWoCID6M
t+UU/nOiZM8L38Vja0gFvmWMO5CgIuvqWPcL23lCFmUzYZMl7VyomnGpLmmqlvfW
Tsj5z1duVY8XYYDSZnhzqml+jPh2n0aBmcf3j8Hw5q1UYGhMl6VUCcvs0m+8lJn9
0zqYYdIzvRr86Gs/Wd+L2qEAyWqXFglC/jziCsgE2+06yStZ+I67cgDqb/r12oxd
jQtWbOj0eZ7iF7W1B5fHu1Hvs+dCWmsKTQAW/HlBQIq6BYgHtHLfI8RiKGEbTS9u
TnvGdl52YOIOmxRAPClWQhWEmx+y3/WH/2gnYqbFNv6Y9H6KnS2LNx94hZbenHmA
7iA0DXugWAX6raZo4asHWC43UL2Eg7j+oRU5GN+JXS4eDem/iAB9/f6bgMXIQaY2
HwPKoDqoQ1P47y3/HQf7D1zmnGACeuFt6cIX7Ys9UMFI5Z5OIUxmPqNfa0hsX0dq
ZtM+8rNSugtKb+uFbxEPi7iqVcR8qYz0+BAp2p4VZs/XfjNLyAc0yWww1YdPeR6h
r4XN2pzQGJGYutBn+uDVNYrTWrWoBEGRtF7QmWEck/GgrGr8Yp2I3aEGuX8Zaxla
mp9IkzAV0chTKVVNiisOditHjMWWkeh/LrrfTz+uDAMuTe53Q0dMNgsQRxKQQESB
EZ5xJeEWOK85iKMUF4RCf1iR1pICH/hGU+eOKF7Aj1KiSKGgEDIGNdJhT165+3zH
+FmzoAf3DRmjESYUbTcTIMqQuEikHYVcXCFdyG3n1X2U9yhmQSMmC/QShKmyWBJY
QDh9V5dFLewfn4p8oP3kFgpYQjtug4apYtpAr26hiUsB2EvuLiq0ZQC8RDlIMfR/
QuQnbWc54v88OpgGxmc/isPe8hNpi8oGhWScS5nmaRu44BKY+lb0JXXustgbH2rj
18Yc0ys6twPQr7uUhYY1vjbeFJH5ZJr6yIuCIovau+pNpaD6e6He3Odt4wuw3fQa
mzIziRDFwe2ZFjOvsCTrsk5WYrKjds8xf3vQSJKnsPOdrZV8G3YACBZxvx01Xicz
DHl0tAI6+7fMiTq+OxGs0iFCgrd33B4U8nr7ihQGcnMbhfM2mR+M+H/YhLjedmYr
ZACMtCbucYTm1/snIzZUeCLCTrW356ibbm0n/NiyruAJkkAbnoBbooxHx9eqLni5
YzwSLpcqnbbihSVXLp/EfRUcR+Nz+bhSU2uI2DM2NLeJQRKLXWtCK8v1Zd2GrkvR
igfQA8byIfYG5/Z4J6O8HT8qnC8prQfLCaypa6X7wRRRCJA3Oo1f8hOu2Mm81CAs
y+orpIPh1gT9lhTDbkYULdHdVJpSBfxivDcHtje44y9vq1M036/18L2yDWxLCPMn
gijGofVessfO4wiW3jQ1UbNl+cyt63+svaFzmc1bWrs+ef+M58d1V/f7yKyzhkT5
RmLcj5ZefyyqTtdWD2Q7HaeW+NXop773E8CbQ3vXl8dK+KhHmX0gtdQ5ql5oACw8
CJdJ4llK3qrnLCop8RL2hB5yplxUMMcBmz+atfCeb1vEEN0i2sxGg4eJdpIlOQy6
2wLSrbyVpQJskp02fgdZraO8uoyceFLHOAHJZFOHlqsjLmfuJTLVG1uKcJzAQ4F5
Wueiih6LXQ7+mtQbYOgNTXrsfSx3IhgYM9sdhOy29RvvKa1JAayuQ7FIObdqEDPy
GNakzuXyO75qy6bfU5wA7ntf1ziXOWtEsg3tgNlZPrg3dR/66xuZYY6EsD/eN/vG
L53t4cu5xh9HdaroPlJU1fGvXMmvrahpcbDJ1Zu3C4nDtjLDblKAFZnRJAeFX/jK
9IgOIl3PpzPVjGcxdZsAN/gXN659o0JmtHpxhfdC/FQ/JReVZ5JeEOYpQ8YdwfM3
7xmFBocU18GwCF5E1X0a9YlY1U9pImZy1iaM3sk6YiiBCxeIJg4XCx1/9u1EegqX
LnBx5qlODaRqCM+z98x/KW5R0h4GFdDnUFiLSu2HLLhLOL179dadr33CmWCY6hl4
8g8FEV5YDoF2zIcPsbQe4CoJ+cEnevhd0/dEXo82U4ln6pRTbTIGD+AtnYEV6oNb
fQuh8nDqmCH5bmNbV4AxELUv598KwjYWEv9vDmwSHbuXIHRIMrT5VY3s0hRcQ8SN
KBXNjBcjndZRmI195RoL8Zis7kW/Ns4KF3k0qUL3SPQqfz9nCmcxv7t7dZUlQ+bp
V6cMPHN1kYEmTgQB5D9w8XaUUYUgkK2yBq6tH4Uh3mT0+IyMLJDet3oj9KWeJJrs
/BdNua1qPFYAo7PHbqZ9+ZD6A/Ha+Et2Hy85uivJ1uZ8A2on5yWnOH8/U1qdbx6k
QzB/sx93dJOu4+5dc2sKNy8IqN15jjkcRbsHhsfRfPvEgUi9zJJHvm1ORBo8icAz
LXDSgXIAmSXABzjA6soYUo1kyTJz3VB65j3PvIrrrimhJ/emS6SFMeyI+dHgrQ7w
MFRFCgVjU8zObZtyats3tb9gQVEeaWWVfcGWwS7cYjEvVbCVAlvictIMVokd31ut
YkVSXqwppiQUxIZpXuLv3lbSdKQ6HGjhYk2PfteLOx/iOQABJ4MJlnNklQ+IGogC
ExnKVCDIj0b535i1/z4KaeWndrPp0qVlgpclxhC48PDruACCLt3NLQw0+UDyN+1r
UPyu3ory465p5OnIF7VCY3r7bWiNygFmFmhEffOznVfcG/mCACkzGhfHC0xAuIeG
It+nMHaxl+id67rWsb84EFl/zPXrrlEq5TGcbm0jJzLsxw9myGwkB1KoTbr7WRwo
9yzVBQeDDL6Q/rBX5hWGOATw9MlchLeDbWHFDB1Ig0ofZW3F3CoWxz13DODgm+Jc
t7XJ5bXc8b2dFhIPoLoE4GT/yGCIDCbq8y1lfLOvC53VE5JzjL2IMgPMNDJJjOhL
oulRQU92Bt8VTGMrIqQrizKysIL9YuCpeC79bCi9uh2HPiLLN6VZrt+dgrd1sON9
iLahy/TXRVJkcZKnPpxbJDgiY7lbX0B0o5MuTyDOqSFSTZhofg8ms1Y5PReKTk+b
yh6go41mBHa2+L7888bYY0sGNDHXwC5nEJ/sou83tzp7nKb7Oe1ZH/GKVD1tQO1h
pd1SZXSO71OI0+BLbCWw17Ha5Sg6u61CxSs0zyHv3LyagxoupDG6mdH+PYg7rO0a
VBlm+kzAeZvTLQky0brcCg7IBsU36dgkwS86lAr1HJTAdxnciIjSCYn2bx0timQ7
BbMT4/0T4em0GB7/9wx/ll3jx9uH9oc+sIbB68jUo5NmGkYk3TRWmBrxsdzuh04k
RQ0cCeuOnVFYgDfhilM4i7kZUGvOY7RsdxclM4KlTOyjoZuUBa0RA4FSXyx11fRV
ZFPyfL34wIvV5e5t4PtC+gqVUVZGKImUsVDNAbZMc8WSjOtrHwoYGnyWBzMteKJ+
vb/ewQ6eHS7UiHyABKdTbPGoJSum0S+HHp/cCUPi3U2U+4rwDeH1hHfPC01CQ7PM
tLzAL2g4DgO4war/F89rmpFKilYf1Iwe3Oi4VO+d53Lt0FSvLN7Cg/JG3v0aRZFF
aupyAR4en62dzTNKxjByw+X5PODx8kht9XrPbtWxQbWT8pwghjkMNWKb3k0IAbup
YtJt9bBnVIa8h+ubFDGHpDaGB8xZFnvCj0bRDHUUewr5sRyw9gajlD1G6Juh4faJ
Q1cEXXh0xIeYjJGdkTjWL8YNlJMHxnueIgTNJiNn3DphPK17n+/9C2OzcGX9g04u
a+gJSTsikcTdiucpjjiNnS3w8T4GL3/Jk6aYAvF2gnA4IHJQSWxNu322A8/ou+Vz
nMXW/YlVw+JkinNocSC3WH5VRxD4cP0DcccROMxogZF6S5NR0kNz30tAF/al66QD
DaU5STlAkbEiho0obeoxaUxFRI9pWSaPiFl3/GGEToUhSJaF4b+kIew6jxyHPs6u
JkLALD6s4Q+pLzAve+ndTckopIfp4ZmAJcOHOmXUBMONLvVKaTWbdPf4tTy4Xrec
q6HDWbmeY1fB5HbO4KcqtV5MLqIRcpci95WHrP8pnpVzmUu4ggS4HcBKIiA1DAmy
szFI4WV0I1bBCUUgXsB1MIFAtOC1eFKzeChGhaOi0BoWuTJK8n2wmep68quN8f61
csOGJqnCM3iFF9fX0A8HC/nEZj3Am5fmLWp0HKnVeOrjIjUVIchwTQ90G7lL77bc
i37ZIICSHJ3Ly90Y+KqRnI0E9F2h5F1Sxhvh3margKzOojCnJJW+WLv+YLp2SLCe
5P+z7vNiaqXN5JCxl+FHirrhUc07girIpuOTBQRn0gAy876IO7+UOuV1kwsKFof0
QJJ+l+zEjUutqTZs30RDQB7O2TdgjHc+tV/wLzdjOklbpRaYyrbvjm6yYVyL4GBy
rJjEiAIvwMyuykTY6CkdvsUk8YC7hEbopqviRoNlptrKYDQp0i1XRWShS66/p31n
j0pL35lzDGJ0/WTzFedMUKpAXQizhsq6nYdxU5+G/5isBYD0dirfT5dcKTKhGaZz
yRNnEsQgbZYLwwvLxVDBxW6kG+lQy9yxy4RiHU7sjRvJmrryMBd6xB+FuVZOEyx3
PI+e+ZhiOf/sdOQopMz2hcK0VY1x6gIvmuYh5UWd9vlW+aQX085gHpnw9aI5w6K5
jsULWlk1bMVMKFhhlehmzbc0erkrrMBLBHHgY2hZa5fFOS91Fe/9Pqn4ySdiV/iE
Gwb2EZSWp+g03JMYtvD04nUJfP8PrfiVfyoW2owwLHxVeRZ2OfY06bmwz8DjANl+
GA5GZAiWggtT8rERyaU28gQUUQmaod3iX21uzUqt2/7GHQkKAg0ZxCutCwgFNmIQ
Y0a3b1byPycOBccml9otrV+43ndgGni//fWwjp2ulfhkLKNXvJsucEwM1xiam24I
XI5E9cKs/BXHuaKOo24goCkkkq+UOfG/5gWgGKeGq5JsPA4vGcTjrxrARwogDH0F
+tS7zjrsxu5yM+LeWva5AqfWtIRNOkSH+SOWdjUbAKaYcu68+xhqYLBVoPWPC0FR
O+BVA1yyVBXpSsRkf/rOrf69WvicYiwHsu4ywHP4DSAOvWbV0YtXgmG9kJvtyP0F
x/xX6LfF7VKO48USslioPXcIr3k9Z2qg8yBdOxIfMm6brMR/wGBeiBg02m0iNIo7
pYG2xu1A3tMVKBoKJB5jScnlIN2BWABdtQsDLq54UJOH3aDqPYqw+4zJnQBKKn+3
2f2VolX/x02CDfzc99LNyUtIPmyVUzPj0r6mVktgoaXXQMl3JxuXusd6DcgmCoet
1VA9C2FDOYlpFqcFFhhs6IChEV7TYx/Ky/wlOd3r6gtt5aAGbFb14soHutx2oFJ6
j/vB/ktYJ+bmA06V+8YHqtzc4ltAuxLegTlXStTHZkixXMs/57ijwZz9inuIVS9b
sD6oVPLwEM82E47dei62PdCErBxUvdS46MvpPTLf2WDyziIoD9ybnX9wfbmD8iQt
vhmOa0lgDFDKS4jzxi5v0hH01dhlFPvpVidzsV1f4onweHFFPdeomPbpQt22UJGh
CcdOPZ5IiuTq8eVjUaJXeAEOOHmV9BvtZ3SKwNaqweX/9X+ZTOoN0neEEXgiDvIF
MP/3WIi6mnlv06axRM8Z9h7x6yWymJC/Q/IAqGuaKNmsTYP4pduEw1OTGfhY2HoY
tr8kQIBA4HRV2ZlOVZ/KW/JhvfPx5ELCZxLzRYW6ZCLVyRv5UPZUk8VJs+VHbM5d
Vrwsc+XWS1LYAKFd9KsU+iY3/10Qne1+hOxVF6DNRht+1cO+xvQ71BDhRPl5Srs2
Uhg14VIhGl0G3VvgsPQWw9k3bjMDLRAXf3Zm5DcWnDmi++nmPLo8wWzei1cS8oBX
fjaksBuLNfKdbgaItxoBCJ9NnbOCYH3t84dQ/y8Wd+pGTC/YSTBHm/H/NwdPgAm1
1Fjajd5q3qf9UHIB5lAnqWmJ6+afrxAv660eEj7zP/f7wbL8HT4923/NuaI2Adz2
byVbo1hYKnf390KyWuzD4L7fjC+7yMgC+Z/qblsPQn7TjMZIHOgjNIKFE3KdgGoJ
e5Fw7Yyex47/L98q1QP4VLFT6uRMfT5dCWCVpQ2lbIrP4hgSHcoBF8nZmOQ2URdO
mneeBGxUqyIAtUeFH1wDacaCHLbQMPKMJUrAfCLg8K6XpibjQw55jyg1EWmB0xxo
WLjgZl9i7NMyAtytXM9WiujPqf6y9gfT/uLkwuq6HEAXXWB56oSXQjHQZYlv2y4d
lEpFn+GKSVzCpuFqOB/FbCc5GEFq+I12yWLaJmPifNfAQ4dHHjXH758z4myG1gDM
tNHwMtuzWgxV8PEtyqj1DbACDy2ZtFRTuAx1Qojv0lm0XQRY2E+BwO5uFf+2NRKl
LPuvxOsQnihBMhFJxtfBCdwxLjSKLsIB1bKdvyyqI5pQFCUhczq8hVpitEg70/dd
sCIy6hqB47BnGjjU4mW/bHvFPWnFczZjUC40esEqcNpQMW+bZd1dNCzxtVmlAObA
SBJL6PevBXFRfHcqRV92kmhLnR8neCJ9xdIBM4GlncVdJoC2+Ssh8StNGqQQeFoW
TNj1WXcf6VU6WeopEZ4zGrLi/HvDvt4yrLC7FCRtuVbOa2LDhRFrSnKCxP4jK88p
zIDbwMqkFfE+mcavDirBe1iH4eRaOachqSgYwbd2E4pHIi4xrvMAwefvLnwYMorS
psWXkcAIKBXji1razKPrLZ8G6Livitp9eopIvhaOuztpY6D075LUcMoY13KCygrI
vAi9kdQx8l/QjC577nech+jCeheDilh230YxhJzpCu8rocAntMzji8AqfOONuhOc
pQ9+fV5n2N3vcYEjLF6A2P2PJRfR6A2lszzWXZLI8D9K10bGBUjGJ0XADFEoX7q4
g4iX6vmlYeFHRKrEdJP6Bqc2KX4yv+GMbLN0C14Jk1vkZgpEGMFApkH4IddZC8rZ
Jk9K9waOyaenHWcnQALjISVeZtrdF50LCJHGs7TT+lvzTU/wz2A9gU9HEtMmIgXd
ZIEvhaiR3CWcH0Il+/56fjkFLZVjd0Sfw+CnDJsbWDC9lfDUP37HZA3D9uxX/em7
tAk2WvGE94weX34FhR/mUHvOvPDxIKowSuJdzT0sF+z9VcX3/N5L5Ca54XH3GM5K
X2Bw7GLlEO8WvJzV7rMGgfp4X6tEroWXW8nth81fSez2XLIc1jM/2IBukQO1Cme0
e0d1GyNjW328pYk3jP27sJA27yjJGAUFDaaNJ953okKMmbAaiWm5YlcySAxNzmCD
8S6liwdE3hGkiOIopwy36VFNqpR/vfBpu4cuA1Wzc0O6DUITaIx2UJ45W5S82XHm
iSa+pX5m8WfNQF1ikKA4VNHhT/6BT+x+iRmO+dZc0QJiivnpGtn2CwfPQTZ3amcf
W5YRJHq5fplmLeyDO9TnE3uugfQT06wkf6n/uIFhMapgj256/VGki3D45zvI3cZB
vn2swDTN+IGDqj4aHsdo0krLFZs27rZTIxlcZ7r7z7IcmTRCf7pwogSER48kJHye
RCTsTmvSkAaP1LEz6NFR0P2/95lm1af7UP2l7FcYJvgjrLt6PU66mSYpafugJcWc
BBJfYTCW3wlAbA8sSd+C/QJ6Ay1KPJaUcJRmYT57x4plgbFDnAIhVFUJPIvqTHNu
CqY31yhRCH54f1G6rnXLtI/VSttYnok+wJ86pNdQyvdHe4h29K/dvWz+VqWSSDxP
88BH1i7sVY5RFM+zhPCFZmPC2dE+THcoCtqMSXn2rVek50P/5zX3f5lHe1Kr8VHk
xFle2RFWI0y5ltsgVcADqHS8TlCXmNPb+s3DlZRCsZUjZWo61WPskPotGhuhirq8
e4Vvv9GL9UNQc2lfojPhxco1kPTj/njOynT6eGxH0H6zt1d7nWQnSznrvwih8MNQ
3wHP10dHogz7w/TYMmhXTq/0wVCosbQjKu6kfMusbCcc1hJdbVnbQVm0wBfHtbaA
UIOmeQ5BgaC6xkpAAWVsKsI9fei7VvKhdVR3IZA5ebmWyac8RGwjYgtu/rtSxmDw
Ie93SoEMVYZ4dj1rtQ0498ubfO7x4OuPNnDBcBsDJlrCXePKeRTOwSEwvKZF9f7e
rFtmEwY+M/xwWTeHaRKeRjQichrVkpQ3vXDDOy4qFFs5g32ssZq6Qjs0+GC0uzid
0YMEOvtMRsyWe/5c0BYnK0hOaidDI1zFxSyDRyfFg2gj1uhuF6lgrJda1+MIGhhf
gjSSvo9/zlOrvaS9o9UOpdRcSLYUbR9GazD5N4rUHC5fB0ehvVCddZiUh2M3agzq
dRENuJOINwor8HsRelRoWFAfLx5lwMbdzDZMzxCO/9qidBrDO4Y2E4Aj5uNpvCSk
1kY/fx032lAowdsCYeSbUeLd5Q0vnY2oBAWsxrVNkoeGB5rjXJMKTkZVgAlOsNEQ
M89THJtHV+jJEMhAeGzL9LrPv7pctDWSrq/QVKoejOj14zK94QrbXD1lijzjwYDG
4TrvU5URLmpoycO+JmysiyhIa26fKnYgwW5R6W55aktNR73BkG9VYZAtcd90yUlS
3bSHOldJanJKUkZ47GUDrdjzFfJi1VA+RwdvGCwYyW1vbLBdvI7WBhwvIwA9yF1v
D9cvqvbZ6pQ0YP+Kn+S0Fma302SggiXobcrfa/H7WbdnVb6ZOsh3RoAWYcMM4V5D
KGg3EgwmiS/0qIxL4EgNLW68xpB+s342juHIiBwnZJqqbtwODOslRafaRUuXCEcP
jiWF5YqxqI35BHqk6if3blz2j+CavTvloyLIhsI/vxTgkQdYQPTHhWEFUi6aNaFz
ywjGOLFB+55YUIHr3eFD6ycq9FK9Ie0HPNQrBg8NN7Efx5EfEOLlByXHsoYvjF38
WLBVPSb6pvemKfi1PyIE5MPF6v4uYI+9DSfO6PviYuElpuWO/uz17ZKlGoCow2TK
T1wzBY0M4BHpOUA4QamVDbYQO3nbICmvxv9acP+c+r15arNLJRK3zZbHn6bU+CMS
0v5w7SBxLwFXhwudYZvvVOUovL78/ev2t6++S5kbIMulNwor3GZ5vnxXAHRCAS1O
G201mTOnjYeFhOR4N1S7ypFcLdi5jE7ESOxrn1/9OPYWNdY5jf4tWk2egRtT3lvP
95CwsObaV7WD6kg9ub6T4fw4bDVjVMGfdUNCqfDwjy9ToKZlDi70J1GyW3T+3d5d
Rizr3zCeWuToQPFB9m7K5md+Vs5WclzMfKZ4AFHC0Op82Qg+vCnA7n8CuHpbJaYN
+nH3YHLifc8qmFRRDAPV064Z6mS7ywg+RBfUOJbvaWACd89aMJgvbt7FjWk/v4X5
NTbLvpHPRBU/6aQ9BWq329rRKRq3iyd21die71+WbTr5E/T1J0af1PP8qb4GCXmt
X5s4ou2QYQl4DflihZm4SdBZDsC2a5VNIKP9J3sGgDIgGaBUsNYMGnsZKxs4DiXR
K/0qNnMTtV3/Jjgc2/35wmfrF+VOi2Log/QNvFq2ks+PaefIKj/AAkZUf3/TuwxA
VNKWx7ltyq8+q25N/ik1ZN+eIulFNlkMudOt0KEU5DRlDXozzye7D0rfmlcTUvZ6
y97V6Mrn9QwH0mP8OrmdYNQBXUpSlIhvQnJoqR4f2qMFBd0EldEIrICgIldF+K/n
gaObGy8NG0NtnOz+31k0GOHbF9truLNRD//3DMtYaW1PKmlFwgTZ8Uv/sAoGmKeT
cZV4cv2FiHYPhw+WdOTIA8PvTsXE24s49GVOblxn2SDHisK/uH0tvXiBGWGN7tJx
E15fu6V7IL7z3T1Ecum9T69drXQ5wQijQqmGH1crJSgPZgK0p+MhlRcnVcftMCZn
8Lx4+Qg3P+dz1FXvyqi+4xyOgPo3TEcrO/BOACtmuLR2S0crDLgXwWwlRSjsjApd
DniqgGO63eAe4KwcE1hOkhS/lVamYthl/d/GdV2X0MU9M/3z9cXcb5VSb5JAC4M5
cmQgXz7vm11CZg7yU8olebmbZ9AC/wZ2X0+/fVeS1U2k+ygfLeOJ/rBsC2DREQWb
BUi+/uF5wUGwmQVUuyL4zH3VbY7yF1Fl+SLO899cuGoaukhheMGRwC+WxNJzUBnQ
n7DqAM6qTC6yEDBu6JfQbLxx6u8eMK8XuU35r6Gcr8qc+az7vjEtZEQhFjcHDRtj
V1xm6HOwjARzuk9OJ117QoxF+pwNGaHsztAqHYgc2kzS9TuvUXNw8uPbciq1+tBp
BsmVuVKamYP3JB2Xx8iA+RMyhvpX+ZqPIkokQVZWMmxIp2UwSwOu1TNLgtLzUa7a
a1a3+hRFC22A1aJ5fwD4/jGJbWo/bPBv63q8lNIlx0Ifl7GXr48ytLTlVeO/hw7T
8rUsLuEMEtTMJjaZQCYrplVN2fu8F1tIXtI2053bxwWLNSmqB7w8HQK8Fha048Rr
RB73eqprlR+Wl1sK+mrR1Ln6FLwdpUfCbUDvHDtHKW9eWaSryAQVOmDc8RKRVvks
H/p80hogjttMYzUW8gVQ65b0ahzZLHOzV4UeOAUoEDhNurDTLtubu8eK+MQZUzKF
/06Tdvqufo2QWnNiM5e3CGdW2Qdfwrwef9QaMC4YFOSXxz4OPKgYgu+M+uJ2M7+q
hk0zSF2msEZ2mNFNGoj8Hsyrndpt61L6Ub9uZQbJzqC+bmmPVGxVvfeewmpZ/Kop
uKJ3Y+Od5PWavRUvSTEK0xJ44GKJTrqbIuNTgVksz6znjXEJ5nj4duH5Y20qxZrO
8yaprbBsH5Y6+W+8YB9GPTUfJOgwHo54ohyE+FquLpH5M4y6hVCW9pFqg6oK5EJ4
rjT37lxS/B+USu1CUstvyIz6sexqEKpdZun+Hh0qppYPej6DcKaPcZVH9S8qqtac
qNziYRPqOoSDyRsqN4TmwXwh/aOmNXSL83PW3GReSat4bkbiceIlm5ftXC8fGwqQ
yWiT7zh7StlxPyVB98Yw38QOi19sbcvw4WhpsudHnQ2N/XW16glXy9vdQTH0AVDa
yClZ1FWEg9w/HxALPGjUs6wx/GAvIvqzzn6DdASIhWhPy8X6OjVHXpWCRMH4gDZl
Wc47lh0IJw9yMvAyNR49RhFO47ewSuAvKnVL5aVv2qkH17Igl88vwYLLM43IwC8m
2OMYHrjRdF1Mb2RD4fWi81WmVFCyK/ApTNCfHWKdZ0A8RfVUcxa7/ek+b0b0SqCm
L7CK34Qw1Wcdu3XHKlCNKbJwJepAWH//TpKsoseEH1f0MQBD3/mqwMeeSm+sEsWh
OFZLjSPaPCl5UpaGg2nV4VFVBAUbV8f9Gl7ot4rWa3zQlodNceCfrrYWJN0+HsV1
kF9g2/noEO3LtVl/SYkodEcuq5WtqJ/byvOogVcdzhGkXNG2QdhDuRiAqOtLlCI/
/sGpK3VU9/irMozTW90f213Ia78TJbnq8v/tmGDGF16Oq6lnXIsIkUmaAc4H8tI4
26pQCopQ6UbMSVP0cthew4y/dPwf1xu9NLw54RGR66sEOMQhYkfa2Hop4cs6u90U
ZwVcfXji3d0rOFUgfkj3o4CMMgd8+4BbGD6duvuD0YRSLbke1KmfGHjYGYcTnYRk
jHQ8C283DEnPn92H7BOsTrpLE+EblyYsoQ3MpPT9iBViVrB3j9Y5qlU3ngkzBWVv
PSiAEH7jEKnWZtFziwIXQ5i3Do/67LNutamyPe/OycNolrlXkLDAsrocPXuyf2GO
U7WGtQMrz0ILOvuIX5CLBOTpMGb6G02NCD+lCc98AIvB+upsFAxT2z+gAPR0u54d
FVPSFnWG+XGkHtHcdn2yro6nQzL1SXZOmI7EOW39J4amktjnZHk3SdBB5xPwwzJt
8C4s/GFWUKkr5Bbdt/9IDWql+867axGIqjTqtN8Nfe92nLTK/hVz7r8A3NO62DgI
3sDZj9Z1azLaUX1YPiQ1HoigWURTQp1BEQN7GKEyfWIenM1yYl5HGXCWNWKzc2Xs
IxcS4M2P3k3W8KEzsfODz/geftyyuSpaI1Ft6nulru2u3MtTWgE7RZQjmG3Wftap
BqPvb4ieWv315ukqN1MyRtOe6RgB0PfwNHRO9xrUIQ0pI8+1CLgbt9Bwa14i+wyr
0fkevnToFmhy48LT7/c7OL5sd08bvHUcGcJYPc6QBrUIvTsYdc7IumHZBV9+3Ql8
TV+qgxq8jd+7zPTyU59+Z/GHfdevGW6iE9QdhT8EtDzTpwRmNU1Ik51UwTw1tIIa
/6N+0MdjbX+tjIyDBnKm0Gf0/ncCR6IDw+AicjNMYw1V7p/xUmJB9E7E24E1THbF
tA/3wcrI9GOUfe+BlaSSK01FRf1ZOot5uIuQKqvW+J5n3zxpufGbn+TUWeSrIyhz
hEArlz1lDl6vsA9vw2LCJ7lFSHBO/Bqok4Pcbkbec5kHOCpaugbi40GMbGEYcKNv
UJfiPDVpBc5p43JbdC9207Pssydo0LBRH1akxmm6ilDgO2gUOZ66QYdqxcS70pnX
z0SwxdUNwoJyFIhl+UoXgDtpyKU1q22cltiBHJuowX9dfGfG46589e3i93heMdIK
iBa84rmbs8x+Aa62ZdLLc6fq4+Rf+PNPgg7uz1vS08m8IucH1CRMp0zKiq32uggR
TN23K0rvNhXdaudbKfgWiYeCk0rP7hABQLahFPEgEzVmUq985mMebxwqhr0HMSv6
KpmHoMWjprgR/YcXphQKJlqN4s8WuFsaeWfJyAGDcnWtQo5BCBvrI5LegkNb2uLc
9RCyIU9HyWszNO9bBfngN29Lg4Y4dRgAZ25QXAM3bimO18ovLVFwaLvuEZ3FjyAy
TcBpHIAjnlKRtAOh9+SQA6jEKrEWrZNPdq+YBgousLwRNtpHDiqUXkkiQmNAfNAB
OUTCm+f5xnLp6SogKvlJHnetomwJWj3FrNubyR6/4UXRYaZjP9gEKKEPMX2on8fv
IlyIpS6ZTXpBxq3c64olEGrBupJnE/oF1pIJdouCXjjCH90oMAhPPt31HAF6Zx4Q
3f5HzybR7vDIRsychLc++L5eHiBZDBXYSieXa0pmWCKyczUp13MUq7o/DXuPTkRl
KLIgIoBAAeN2zJjU/a+QeG6bxA/rBrFFzm5KZyRLMps4uauU8T+Ly7s2zLZZiHUB
4aflVI0vizg09rftR2ATNlURnKftRmM7jVa6aoek8+QFcm8naWdGIDF/tPhiNY9D
BRyC86JzqGBoOAnkJ5CTcniAqEy8URZ5M14rKDXNOybGG71NEpwdwZT13fBantEf
CBc+iXYb1TieNXQ3Mqh30DxQH33Xd7WQ3Wc1o7JWrIv8h1ALhns/SxhJgip3Of5I
DIxTnUx5uzXQpvtDrZKTSKpIWv+MyZp4JcB1l5TSxqdQyAMdj++E0tgYjelRULFI
leVKI/P4kiYnZm98jRxY88NkSvLSkKqnDKdR8Va+/CaprOUFm+JUkERquFMFEeHK
afniDkUh7YWzrs1IN/LZ6sr8xyoJrfOUQzSS193llb4cgqfcbM8wVPUZJ5JBqb/d
vLiSnCZQbGLSo7HhqKaVbRLnAKRQdYSHPktZ0nALUdNkGrVmjzG/xb2l0IMXxTGd
F6GmcMFIN3oQEryccn9RfSImF+R7JarVyDNJDn0W3aGwqa8nY+IyPt67jp9eaoVh
Qu2PXzvcbgdIGP7sKT5+WdGw8mmCwWBZGSI8nsjqPEBRPBGv3sa9bJOr9Yy4E49m
KRDki9vQ5EczwT+58dB7Dd5KRbQSA7EI2W8SWP1W3Tv88DQvuyQ6Uk4K8BxI8sB6
C00NuLoGC+gcha6xDKMKArC88mA90JnXCeSM/LIwmVTQgvf/HlfW85r5KnesX0Jx
7vUw3aB/3dVspncvXVVjSF4KfzgNDC4PKkd2NCqvvHXJLaeZzG/evy99zqYKGeiO
UJKVeSYc25PpGgOVrUSvSaz4tqLSCbjPtkPizNAkcVHzLdkbIQdx4Cw6Q3SRTYyl
8N6nK6f4C3PP8JUUC4BJXg86ASM+6ZuzfpxPBV+81G1BxvG2sUVtiuBrY/NfREkS
05OG+o4T+jDMs2zZ1gftkscnypsYUtWvKjWJInxzpp42avEpb1+RcHHktIPM1ACK
cmzZ+bdK/rpHOY5/oFJecMCU+YVX76HGvgEd1s7hMy8lfvRcC61imFJ49/3UzAWu
DfR/bC7asx6l5/Q1H6kXRJLV6aF341wOr/xa7NZNX0tUQAM/Cnytf+84uNSVsOxm
bUywKPtfyXFwOtXJJo81/qSypmWFN7ArSGVXvoHa8jprEFHPiV+wgz4Rd/lAc5E+
x2X8Gf+msuek+0f0tK5R1dWjTSTahqkvjcHMsOZwBWY0R1GoexlbW+kzSikU3V5g
hU2p62sIuaKo+IBnOOda7VpUZERUoVxzxI+KT/xisbdx086XY7nbd8LfGGC/1kCj
yoUFGlAifUDNI7vF8J9Tu90qNjFSFauIgWyLRnIAskXGLyHg1zuxPXtx53siv+T0
B23139xM7LPp8k+dgYdr7oXrVQXAyMOWtl9Ng528BOd6VTntT87D2YoutohFNrLs
ozfcZohevsl4uqGGy1C+bvwky+agmu8OY3WaSSEDR4rGTkEgFnvkZvl94Wat0tid
dltJOnt6+90VIplT+uOuINPMJJMb8JC+f3jdBY3a598Uhux3jNwsv55id0eY5/2M
XWovbxI/T4XXqcHLD9Uz9gMTCzLkqxBE1v35cvGK96KKgWbEpvsqcyNWHtJOItjV
7d/lYb2xSpMTjDxAHpvnbUD8oAzYTm+tg+6lsS0CzeNcbMCuGC8NGL/bEM8CixNB
la50/AVDeJYdr2w+qwVPYDixsf0OT1Kea+L1bd1GyftZUoBouY8IjMiGmRMDtOw7
DypP3pEw4Ii3nqywTVLpJspYybP+/nq5HzaMsMjqiLYo5NIxEHV5F3dqDSMY6p1/
LAJpeYv02jn5z7HOGTXoASzHsw0m/b86Iqj2Vg3rLK2kCHtgvXshN7fzvXbh9Mis
UTwTi5cCO1xPBJmsEHCPAUlqQ6TotHGplEYPIL9eLzZM94L4g58m8jRpltzOW3ND
g7Qu/3hXOuEPrZ58Rn6UyqhOCQwKtYKNxAHBw7JVva5GXZpBE89Ni40x1L3Ql4be
Ctpcx29h8DUdgEo+rZ2m7m2T+/HoYJBu7ve/oDRxIst/P6xsH+tXCQmRsUc29n7h
MMgO7ndYz27TIH0JolkcHBdii4MQjKmrgYfZ0zydD0WreHR2HvH4XKdLArEpcIUD
rOP2fFOoBKzw/XciZKkBPZKk4LfS/yQIcd5JfnjCaw8b9eWSMygM2WJHmtMxmt66
K6L7I4mAJWUCprwM+cVKfdJXfGb/61yP8DXZA84QuDy8SWVnquL62E5eAF83eqZh
q/q0g6HF+JaeXGBGPrjwKG2iQnnnTnYF5Zk1tWMDXoOLKCBGbv7RFaQP+7FqFRMY
dUFUTnQ6ORl8eexR7tgf4iDK1AItGgELMSRmrvYwjJ22Yunm5gY6wbGWIxVdgunC
m/L+LYcCr9agXEQeHFj2GE+1jfyEw1J1NjJClanoOhUThA/Qq9Yo+VOugzFUcDl/
0wyOFpkxKtQ9n56mfKxqoC+9IDuqvbmERlBnZ+6HQN1WHOEgFD58XrjASUV6rIcd
Vz0a4C9C3xvSEOWASL6Pc0N38KYvz4X91b3wPsHvEpuTIjERrxdRUxzHs/hqtazS
s6zDELd9nF2r/V4Y6WMOTlU+1G8pKTMwNzup1lwqQ6MdcPAZ00KdJ2vnVTDhGNuP
es0ZtnliE4Z52MbJo7Ox2hc6PMCNyXJKnrjq70rSA+ctA0YKLYPVo3O/BbqFld/+
2DKUUSOncuyQkKTVWFAYs5JjoLtTalIyK3SpP++YtnF9pGi+u5Q1aABKERate0KZ
vGy8UdCMMeFmUcY0RGGOC2pLsBWt7wjF2rdleApREBoxYXprFyFLMosqyVabckd/
s74zpRkDAMi4UrjTwUNe9FGPipgNYWvnO8qtetw9QUgUzfnU0GToVZ7JEMUiUboO
SyTbWkanmBEG6PIl+rumqXGS1pyWjO0jF+IptAD5uLQT5YmOWfdzxlwvzN64pxEd
NFYzjwRy5rIPhMeR0oTylviU8Rc2/FI+wZLFbubUlzL1g6pvcKffQmLVF/n7oitk
qbrTHamQ4ZhjiNRbDwAN2s/R2azq1BvTCZDLI7jeqfRhACnVyx7iFgpNViy7Io71
gkVOiOiKUNLhBfcCu+1aPovqmb63Xb/ojGCtdDKTEFFM7E2danCAQ2y7yqp9nlaj
AR44ZlzGf3hrWZxaYaDETQVxb8mnucN1RHq0UGAzKrb03/YzZkQI5kbYHMCh+dj5
b+6TR9IZ1TXkcEuKVNMMbNuNGmc0Kd2MSCr5rQ4JCjwgdPBAZddfeVUO3bqSniYu
BPQGT3Hs8ZfsBBMHqHGRCwa+bkpy7bwiMRh+Tix1OFQiaQ77eoGcNq8NnmcegPnw
cpT+YwigduAMc4o+v1LWQu5HnqBiPyEZ4RSxnB3GCtv8RKqMILgg6DqzYGs8mHv1
REIefja4esm7WFZOTV+GwqypvcWsFPqCb3ua87F4131sLzYGFswlIDIz+67cKoc1
wf1ttzu7RAjlipprjWh0GB/KgDyGkESKSIQfnnbRZa+N5Ub0sJLmZKFkPlSIMMFe
/qBaEqBi6uggKNbyQoSnZB4hTPcz+MMMbORf2nMlfH+m1Hy4Iu99lJ3xyFz1cVi0
uK2WekuVEcBnZyDCW7zLgApGp0V2IGiD/vr9GJ8MvWUsgDnr8hK7NW61snDW0KCn
YShbTen8cqxhkg5GVTHY5dHtyA2fxShHd8q+gk2d0e7sbDIz0LNVphIp1Q4xo+9v
szHKzKv99me8eWB5wrBlcX1r5hZ+RHw1ZBsPXiUJ8VIaReJu29EuaJqc4kDSal2D
eHP/u844YXDrG3Ph7Bnxl7QF7v0XVzcTVN/BZS2h2IFkN1XwL224So5F21vgWq25
HjNHXfaHC0HQIlgacGe2txxQQYWo5BlBkt1a2Rn1lwB1Yk3qQnhb6n03tGA83nCv
AGD26mia1kYwUKbZTWhvvyOp06VABILsanooONe3zDplpxOlCZJ+0KRbH3G8S7Eq
pDVFFmwwXgMn/oW6laYbvfUj3Q/rTRIJReiWvsYCy7S0QPUDCwYn/i4o1DlTfHnB
crdcL3/r1kCOTDoTLast8ccwZwfml0ASd2ExRyTGtjGfldGAQIfOyNHHklna3Ij5
SqpIJaLU/EhpN2aiMAjA1UJNOP11f+VtqP+32nAqifvUPSLfnGQqctZA7xyNeTyY
1Cv2tpPz3mvYRd/VjTVqJnVw1ob2XOVx9y1OpJ/ErDk+rhf03SYHB3Cph1kBw+cg
UC9ODueyTp1wfeV1zaHOxa2he+6zsFLp20OfYhodfeeE091MEOW4nZKLD6qA+FD5
exgFKy+PNt1IAeB9dJp/Ng4iITMMuTTj8fY+CcxBTum/UO9mauVinNECA5UjSZTm
eqD10mgiicBgvjmKcYjmkwQKexu2yekHxmQH4RMAX2bGIDhKzixE/liTSS0Irvur
yL/sa+Oj5a6fIqif3I7FvvnB//GXaKZ7Y9bUl5t+/FsQycDEvmhG+M2CbOXk+1LY
0tafpFichUw6eub+4MVk6dvnr9JiYQxFgfmaxpZcdedf3tqKchlDBoewJFBdD5Pq
DaG+XN4kuBatDaOxMc9Ts+mczsU+lDcJ75Cam2R9gkJmitWZgM1t9sf+v+UbBFq9
6UgG9EQpKZ7FK1yzwaC5Q3vC9DweSlLEqNlXiXEqUMT3manJT3hfSFNdhGZACgoF
YOF1DEq8hBLB9HL4x8EBSvVag+nZ/PNQKV3m7a77xYZFapNe1BfipjUqlChJJQ2E
pD4RrvHbzbDK2h5KZ8wZXpVrk4tRpzK7Gj8Y6CmtfTQ808+7Eoo+a/qcA8jVUIZt
yRIMMSUs7DDTgLhGQzx6SmLzbxA+9lfMIURE6SblPKMc+e/Ia+BOn7HSNbi5OsgV
eGliycIwHsDjppbn2RJe5GYOXKt9Qc2YaZzwKXNw7RFbxxgSstN6mC8tbm7Bwv1N
dEvwgGy+IGWwLxip970fxYNsx8m3uZ1HBKq5WzIX09ef8XD1lelbXO1uS2+hXDOd
alWbx+RewtNALoLOBsJ1fL1OoIavj4BdtLqdnasXok8ECUMQLVn1w2oq27RNsA4z
sa6kOcWEsWpeFc7YpmDGABUBiikdHF/vSPox94kjeyDrUo+5IVheq+khFsJqkGlo
5Jpg6amW9toT07+svK5VyjAKLagzSZNeL2O7YBdVop+M5pOAv9NzPAhPRM8kVQMF
fr6192pGw5PBdM7xqb7/+WBI+XycAoalEB5TbvWVY98ARqYIjqbn/iBBC4cTDR8D
VlVXs8vgZAGu1SrXJaRaT386vgZIw9JZhsS5vlPNbnS/DDmx6gf+EChr0VwAcQ7n
lGVbtii4slsCF8WlKp4NCMbxhV6ta3NEK7+L0JHeRY4i1/VuNUI2KSR8U4UcxBVS
aYhHvb2IMcu1fHo6GQ+XESDa/ZpghafV3Wv8AxyF9vceCiCVWLda9NKtB1RVtTJd
2H2j3UKeRHDASYKLlBpkU3X1zPcn+jMbXvEJZ0NizKDy9aeYRT94gxwAx/eAuqfV
iaxTTMowIEhduTFlNGTfjnHPAShzNJ4k0NaSWOGQgcMjoBOnOTdj4jpcV4jidLnb
xgBwUqntanp69b0MR2ftSxB78DeMyWlLJvpAJf+PpoSBRNpm40VY/4EbdA5/R0UR
ASkQW7pCKCKm7bH06Y7NJdtgB4gIjfHy4cMhZ++V5e3RSkBF0eft98EQqsb3N5l9
Xu9LCfTacrgxStVY34NuJT8O1+6ewQCunWJ1j3cGh4owMtoQ5hYWHseDgLRJppuh
OuKd7CjNGwOfCYjxQpYlxOprIY7mL+sWUHN5jo7kna/ywVwDaimq95lR5JamC15S
ekFOuKUbTZRl7DRw1rNMHZv35u7AJIfyooFjWLPTeX0defom2mHos5nP0n1dkieh
7uuRwovDp3TNNZE3GIjlwgHCSswhKr2LtloQnjJw7aT5y2d93IMoeaeymOC9J5sR
bQNRuyE25/Jcj5DlxjiXozxR0/J3hyn54hDRitpA8YnoBTSd3Jz4ggaDv2Q0blD2
CiXq9xHDIrtyoiMKaOLHQkwcuGxPIsq11W/scc6IrHVSLZocZ0guvpE4WX7ldiSH
g1RJnopuX3JtKj+2GstvmFywoj8IpgzReBCrlfyygL/4gf4abRmFXtsn1D3c9vVZ
4k6Vx1vcbARmIJcUvw5EzhBqc5Dd5jAHAGeH9l0ZUgZ2Lbs9EgMtceWXEZJtWR2O
/5CeNNI+FoQ5j5dB0YWz/l7cAfkRH/sFKE3iy+5nCzM3boAThwkg+O5RfBGj3C0b
eUrzYFU6vQFMP4GZgJqbWfRkGXH8i6cJrSkqzIH64AN+n5Cftb2VP6gMnlZu/OwM
oscW9+wtlTgAC9jyqIEPwjKxczBXbrXXkPq2Egw8Cd3AB87M5AlPatpnDsyYvsWP
iizGxInK6mMyOhevY2ShX7ZRAL710fLwUnbYjeMoGxjSmc20HD5MYHvjX0+2ffKL
02j0cAE98IXo2YgEsLD44yC+plXObXwYGgjW0iqpYWoBSm2IaOa4xVnB7QIxAOCd
VrenzRsQXspOBmzOROS34cu6m8tWBHtOsVGd7Nh2ix45xIL5KNTR3eKxqO6RJmWr
LBK7OyhUYz6vliXq7zIvkTCJsJhhauuhuAKupVVJ4rqjcPNxnmu5cggGQb9K11c4
I77PnLx8tkVyeYuz01Lx3Zt2wO7KTRN4o8k8xtsr8E3szAJCksyJ+PgV6EQ5GcUs
Oy8oC3p5M8iBej72HdhquDQa8KVzHvXICGYG4nCQwjobTCnYiEdV2budtPFP4M0y
w3syAMWFM7M9nu5/DxlzA+JKUorjK0vFBLs2TmzSJp6T11aIQv48hBYbXMKeovuB
xSMHvvj4G0nT+b0kgIZNLPb1TmKoVl3eOaXnGBkvqrTcAH41KJQWn58heBCFQ1OO
2jWjHqaUmLJTuZbrCAl5iVgohgwFHTgz2jcFKqscNGA5oMzK6PdnO3ZDaPaJM8Df
PcN0RGg5w4mkamcFxNY4EK249SvLj0I1iwrYXHqdyYt1Q7byZUXC+zOqo0rKgmKS
0K9DiIcLD5yFwDjHk0Iuw/mQd5yN929gVkwEeZTNinIup0Mbbml3FbNAJFFlVOlP
wjx8nS8f4WqI7TeYOGK8XfEKrAzT9kG+Z2ANzYe8utBcyDk6+mJ0EY0Cp0bDjsTq
4yLsa0vEva4TVsFS9byOjOrrjtizFJNd0GpSUp8ERIqpYHHndgN5paGltGQawbRv
2h26IWSACsmweSFc6qTZ4GQbw0NHM45MRv16g/C5vWB41UEEiEx7wy9OvFwfDen2
Z6G4stX1vf17dHx+Rs6BqTWbW5ntiPdjldGnna2Qdero1qPvekFZ1vwyOBDLNlNP
p3VjGNsszT0OPRkHjR1/g+iqNt3hgaF1aXIwRbnKi+DKZyDmzJo9DvreuhkWbOAn
myQ9bZqfFcMjlrYDedVO0Qek//JbQZvSfZ7uUVG5Q2d+RhjtAQZHySmQxUQoin5j
7jBdVrVoHbwZibGlUyIfrldv3/UOnujTN4svpiI6RBrxkhM8lMsOHy05F09NL7El
1CPRyuFviROAKC9/ehEJxoIDt5XJm3J/tms/qA+SLYZuVCYmW/ZwtK6utYJu/K3w
tW4bh8EN8+1Xl/A4iKF/th/Fbrf+ZmRVTJfbYYtJNUtyojUVZcdqOl2fSJd9rqau
tGxT5sS0ZH9U6U5NOXdMSU6o8PW93dks/Bvv8tmSdvoHyp1CrY/g/fzMlCYqvTjx
fLs/jMNSqWgNATPaDNyDU5jbT0/qk+Tvx0ZZuO0xRT002V8p3obrUztOX4zQgFYX
Ow4snofQuo8aFLbYJP1TrF7NsupaVuH0+IqIcyGqMEx6sh1uJfJNK/8IwIgAsw/x
xdhMUmZHyqxuY3+tT14eizzkcVXDJUEOg+mFkIJ1erYU7SeFxMhytSAAzI1dtK/W
ZFyDpAxpwH8KhYaPhBo1lEjKX0AYlxukDS5qanEOO7WkwaE4KSgfOqTIACUetCGB
P503VkZj80Jxz+gTz0Nw45ROt3nrNCAoE763tmKYDJeRYYPUrMKI4csNduA6dQ2X
4vPsmE5lfg4WOTbAUcQ2I2YOVwvX3UVOtWVPv27oOXtSrCb1L03CVXWmvK/nNa43
xXr5rr1mHdCXMzYNRqyzp5sWQjx5O0kH0K05IpbMBHruwejmit5/v+dscqW1yxgK
76Jj1mup+qxvRdoWPDCxgi4JgHW+E7rZEklaw5Oen+eHGXmXdKfS6Jc7CBb19qjD
8pP0UfIF5HgLH4BjCugfZvpbqyZFjK7Y+IPxh+KlIx4sYbgKn3fT81ssT9Bt7+JW
QAnd+RswvW0I3pR3oNv8RgmXPHEcyese6SDKF1n4KtJbJjmH6xL+Kz79a50Q3ISu
Dk/I2qQvSvd3mwmaXUC2KzTB2rq3A1SEgv2lfqItQPth36m945qzYsaWzr46otlX
+p6a3yIkVS06+DtPxBmPCH/Mc9C9/UtP/3hcvgUZwovAf3eeReneyTs87agsRg9Q
R5xtnmYXArZ4pg04/6yXs+Lju64vQmbL+aOHxNdKh2oMjmE/XHbms9iLYw7dcZ+F
9C+qe0dk9gs5kt9vGquI3Wj+jei7zp4X1oAaOJFI9Rl0w6YkJNhYhv7V9pDgpqbf
MNj9eDnDjNgrCZiPxm2DQFJALar6ytB+OSvBPfdjEvgR6YHGPxhn5izTR9mJI3Wd
bpOWq6lPjwEf45B2HNBdSDyfH35OuRUgDgxYn8FFelThtQhjU8gXnoTKoyK7xLSs
Q5qNxDRja80Rr/pINEolU6AQX7euSoj0UXyWuhoRwm/fC1i2N5maOLT9XEqWxrIk
7tI+OpuOaoxapIcSMFnpUxzoKKPBIMd5UJriQCE4ZBNCGPcZgpaTXWC4WfCXCqfC
ZFOQLf54df92MtsFTvJSQ710szDXmo6Z+63WS2HobLBLgOLMV7XlVM3T9kpINzZ2
u35wlV3L/RCzw6BYIyf1ZbotwF4r2nHmc80YHtbDswYjVLQx5W6XSc3sOuluxWNM
gQG7MVV/H9l4ouEOe34qdR4jXiV3cemxIPt/KSYeH1UThXpigrn2CqZGzXbo6D5u
xeVmB4dTjEdEkqnaRuk/HG1s505bBgjBZWSFbGaVw+oFwwLo8LKfLJSE4r9ezgib
UnG6T4qxPCp8QUXfNBW1uhIDwURHrEHJuR1zHxwaUtHdctmxJurpkVypxQAb/2zI
j1sMq6DcCEG5Fzpcs7us1dFK2PrDl04fAf6Kytew2YilejSKfP0FG2ZN6nKniho+
DPCWVnqkgbcoHnGHEN5ljDuf7UZHcgcI3A+LI4HJ5lC5ghbWXvnwSmyJZXFTsFZS
fvZaJI2Qgen0D2ka5WEBUegDzJ8DC4twNeGT/mRCrzgy0t+hBnS0aTqL4+iPTX/u
frgt//O6rjhqWG32Zgh3gZ2LlaX+/s2RgMI8LPNCbSj6gL+WoZdN5YdmSrtqaiT3
WD5BnbEYtWonfHtoBeCm17WJ8hdsJ8ZWZCCRfkbwOcWsgkqvgAMh1WjolOwN7Ppq
IDg52Q0jPVXrGqYJ2gegzVhCXBOTiXV3CisCRfMMwBYBlN0fVA+rxfrcBmgBAi/3
OnUJI+KbQJUw3WcYZbH9Nw+F0g+Tunk2t4EemYWEyYq9jMla29cDfMY08Ks3JRMh
Zv6o5LwqPR0tBGdro9mKIfxLQkIoTDwblvUJN6GDguHMFfYesGWdmgY7XNaDpiZZ
iCfO5R6GaoZcweC6uBFQh1h1UhlkjTNifdYZlv4rREBOGhij2id+hQw7d7tRDHun
UAakibDXpqPi0BFqIHOLiZBBea00fGaFdvLMH8vN7D9qfG56VDtqox25qX3IaO+h
y1FfkQ/t55k9mLo36oWKUnI8NCCD1dCw3XYLixCBploTWq2kVzpn7pmp2W6K8zJM
bqQZZsGfJy/jpGazMdB5Mbtv21FED7K90xr58z9hTBMAJ6iDmtrUA7ABqlcY4LPZ
GhcDh+yX8UcHocvD1MrQ86Rvu3J7weMuCU7Nl2FVlKUFGopiclWa3oucPzUQ+d5C
ZTWOi1VT38eOEvwWOmNczsT51fDPFYJyIDCa5n1VoMe1YngU5gxOvmgwxQXqPpuF
LCzAtn/ncfm2dqkOrSSjnASQK/KeIbkZjTfz8Q2wovXUSBBz5DupyfzV+0BEVY2k
ktD+DxnSxLbliAK+q/lJoXP5X64l3A8hCk0emSYgFTALQYQN3FxmXrVCIp/cF8gU
a9UM9AhAeM85smfSloEE1/ESqDOrpguBgTo8U0O8e5Cc9mmfr90bCh47LJJRV1ul
YvRlP30vQ3VmvKilHlDanu3jsIB7ql/ZlVmghbHzMDOmBRuCmS32VBntPypi9swb
uYQYfspJTylja6s2xqGvWF4gIsiH6bd6aF6qNDBeNl3s/TVO8bk6L2XEPgzGD0Bi
zdPZZJB9dhzOog64zKxutST73dZVWN7GSt5XDz75PxW7UJfH4+ShVQL7i6veSKK0
0uUZD5bZnQEcYNGKyTi8jG+jGON2Kv1RCT5ETD9ejvly9JSiAF1/6d3sYuNGs+UF
uidXfXx7/Ft25BwFHVzymix3F/blr1jcRwh7H0217KMdjrHz7yjHnBDTwTvnoCTK
RCNQIP+y9xpsD08GSskgBjUPY32MrzJFtvl54oa6B8gQeyqmmjdLOyZvLj1CeE+5
14bBOF1U/YZHKbAkLfDI5jtFmWDj3nwat/+C0D+yswOTSpXVFk3+39AHu0XN+cSO
HVAzL6xHlAKUzjZBoughhxARXoMffolGtEx0gys4xPqPq3nAflWWW1DSB87JZ5Vr
CrOBhmwOwMma92BD00Mf/FYEnQe14FvLi05kDXKHZMbywY07ooPNZSEge/lyy6I5
hQxbrooAVYjChdbxkTWoS875+fOTFVuPqy43WYtKFmcGCM1HQIfEpfIDwbPJPl01
t6ud+Zg8g6Xt410fMk5Ug5RHwxx3kUXU8K4/f7Abs758HlYIVw1R0/haoLTfM3r5
DPIrFlyf6gPT/9jFLTRtSHlCXA2PBGCI/pnTD4AZC3AQ+cwHXHaNvrZXQwE20zR5
+K+2NB20as5tONUlaVK67KShERRFGNK6avCfNukeegP+rkPrjnhl/8iNx7b3imyV
nww3LI6R5EsyHNnEC/WV2ydvbmW4vH+WsiGt+c3rHwjk+LZfGHhqw0+nR2W0VnoS
QhbKriJrQSJRdJplTwkY8VBSS42hC0KwBfLZPEOWTufGGDJ5yIEltf5RVVsmGS9Q
Mq1/f0sWYJVHxa0HR7FR4K3xDVKwLPS5i3gNLrpEdbCczNitvg1Rf0M5sCx2eLeW
CkTWOC0rgLQ7k68sH9i8Bw3O6OvEgzkSY8R20Ib/0VO6YIWJ7nFB0uyvuWL6vfsr
ol3k1lE/ef49qhOCGKow4vr2MKIV2tNglkF/PPSmTzG7NnOIMJqQrXH0BM7aOWPZ
gZhutJDTiZrTSCJBcEBjmlTIwbjMUNJU/w5nRK0Sbqp9DyQKgEsLsqdlf+qe5y16
m50bBmKrxy3JyAZdUu1eXnhCbq1mMLVMItoF404C7rX4Hm+EAqioC8Cz/bCbWE4c
tU9gZIRidUHnRFHny9bUJORIwMsr3UKVpzzjO6bx8kdsamuTJXb3LQVS4Y/YNN6D
gjc4PwZo8A0PnpgDBp5P1QaZm/CNdK1a1IF+yXN3cu2eC6vHs3mxCgIgs/M395gB
q7c8w5TEfsa9Rk9PXBNmDV71xH5jveLYMKMXgK5Rwo0tz+X30sDSyN4tLbSDnZU5
aqEtLTxXuXBo7Oi3yiYki0KUi5x9jvL0RY9emEt/3wMQbTBlY0Ex495iGbIiErbg
98pCxquWE/5Q7bC0CSFdCbix1DH0UrnPWUhgAVmdbvAGufGxsgiwsVa4/ozBTu+P
rlQo2upuxsct6gM5k7kglvQ8wKOXxpzblTgITVAvXjnoZdHKHrBMeIKVAqVEuUBc
Tl9xx/9kP0lIU/kWWom4lMJqwfTW7tCl93WW1hDsm3sdv7ZxI5g79bT7psPoInnz
L8ZNbBOzBrd8SxhY+47agtuUZOsu4tknAU8ECag5BRdL9UWSMv7KU7b6ADD3+lFC
wiZt5W6sGXlNOIwUM1wa2s9UsEsw1TQOp73hcwrBlOwY+EWXfFt3FqRibheVAH2i
WaRwGiQtsPW5qdwkIDS8XpBdfYOREoiBbtFaaV37xmctyx3kFZtG/tiKaejcZszK
oZ+fXRz3baeod0Vamm61abesWlVhvKjAJ1IKeddHJpX8rpa0IJOCYl7O+etsLJl+
dO7KHGmT4oGiH0HpnOTG59+1tSip/hK0M2f0h0fKvDGjP9ORRR7p+6Xf6yHjz+hT
k6Bf/U6s4AtzhQgtQaolfmL3dsuQbF0tEND5+YeuEf5vyWS6o7X+BQkuD1NSL0DU
B0PJT3UDjhNQXmcal6a5X35PavYuntfJQcT/dXtYYZsmzf0uuKZXqO+/b2SXQerx
imD2/MuKxY6hq3HXjwS9p/p1lsjhvZmUF6DxuNFKTk7obswjsyjpiXPVwMxabYlr
lFAhVWrZQcTZ//hFer/RUXkSsQ9KC430RUgICmaYuoSf8rxUF6clmCKdbXdqi7Ik
5SSE51hiAqVnMNck96T6rCLFoE/9rLoLioWXGmJuxydV8FoBdA4EJs04UfDXxDHh
yx54Hd/PDf4qj7XuTuq9Ma/rfZFP70w2wUSLJ2tU7h3v7a11fX4uBVd9n8choxXh
cf5MuT6fDuVl/lXwoCG6NTkpFtQ0tKSP4EWOaZZSCnSfWUi1SHhsqctdc66sKuIE
n0kGaXyPIo4zzBFOj0IyEMl0kr5f4ZgM0D2k5fwbO33fmUFt8ujsU+EiDrweBAXU
jdCBZ8K3jC0glwwLtT9Eg7JMeFcOXIHwXV81y4FBgNTGVzA4eKN5EkRe203HMb5H
+990W+BoTDJClMXuolYS0yF6PyLshaV/0wse/V1nKqM8vTKFgMxZMAWXBUm6fdB0
xtStV1cE26bduncpPVM6u0EKoJvVRGXpldAoLfaCVgK8XAgnS97cktAEpFg9mvKf
8fpu0qKV0F8C/h4HpGHXk7byp+4/xtAnCYBktEShJmTF84A6XOfDeopPp3pom2QZ
rp3kLD/2Mm7iTJihWH9DJ2wMPqdkQojVtx6hjNhq94RBrsYHV9H6efCfPDN/u/7n
ozuZc70gZyPee9WNfSe6sahfo+7xqhyro/ML5z/US5XybRO70kp0FxG8yBfiGdpz
UVdNDUWS5uDQy7NobnG49h/ucHRXO42+RkhUfYTtuxa6DzZxfy//qbg+HFWPxOon
2ykmNg+o7JbXeTgg0m8lys947/2+DH+0CB71Oga7Z6FMt2YFsJOGaGFur1971EoV
XHvRBeUj8TfAPIIdO/tCXA0WLZJd2GINJQtxh3TTICKLCXwGXK5i22EfusZOIces
+KBT6FRbg+8Z3xNGiHi8JvXafUqxd05Summ3O5eQaIahAVvUo25JJakXPqjx06Vy
DIS2hwg0VeDZd7SNSG+Otb1U3sAtHgNdDo4rd/twnkGEPgwwpqHlyLNbqOP8kIyw
kNTEIY+cilxBc0qYyq64/76D51KDZqQSOa/ZAzZrXmJ9HPVo3q+OCN0JQx/3rOmk
2PC0PCmR6uvNA0Thyx7+jU7V3LEfgE43nlMHCSeoAlLJpXiYRP/2gdh6vwj2T6Rf
0qIqgust6/9Sk3X0Hn6ICGneprd3hFMBVx5lCizgNzvPorf1Y5KrpFbkiEfVa0Dd
fnHx7dgzw/SBMC/X4vpahx1HUeBhgStTWKJHARMkDV8JJYDHMjirOD9bHS6VO573
KGMClI2praxQq2QWN+l0HgzGjCYtlABzjfrUw8krQasomD9xMUYvzLFwolSx2bt0
++plSr1FEnBZDwc3gYBzZchVRtxfuNFb/6vQO2WAdnOcJ4NGkL9Am8jpbuepc1qX
b4eKZDCt0JujhyVVvycutpjJkiyrn085SmL7CA4czv5UXuyVeZ1Mj/tauiSOSEPg
Sm7kUXnTAw3i1Kaj4BNEQAX1ic1Q/bgXPcHf5fhJ0xSVg6TQoaC/EsKE/6rMgIM9
OVaDwlMAVQ05jfOBNiWYPMelxfu/Tm4redVh4Uoh3fA4FJW+Vl+mV8klJ2++c1Te
aUmOVef35IMj5tsADbNOIkgj0pLxYD3PzaRKNBmqKVGLbM/PQMRcwOquZnRLW8K/
3/Qkh/fMQzwPrhSYZPVT5weZhcGTmIWV3h8UMpEOGWlBxD/U9jselIxX5ilBGJ0L
pyJuvj3tDunYWpOHbXjD0wu596COxBXqjxKfE6VVyaHXHpeMlIPEQVpvEBLpJITv
UWtFK6UfnQnuPxF+0tuzJ7V6EnWcaGy1CytJOtufYXYI9O0FV/2o0DlEbCEKA8Wp
+RLhWbiEP8ILnf9IOoshffvwxFb/XXsl8AVOKRJFRwy1YmVaSeYBfBvjJMcVgKKG
kU/AcaaqjUclYBebryqZz9LQLqb95j1hsHs/NaoiWzuJUg4dOO7Qgh8u1/8fz4rS
9amvmCoXRcaA6rK92uS2ZsbaYmLAChUin7TIYvsH2W0770bK+p5a4BY+PhV8n9R4
+Uv4jdxFhoCOy5TgrgF/nQbOy8DD892OjlgZMc+huEwAg6F0kYby78okm7K6ghZ+
T+C1EOM3IsXgEuFStCYCXTWXozWWN0fzT7vqyNluU+WEIIb8BApz3m+0vtKBSdYR
3YIi/EpvGrLPT14MM4iZ/VxrAAU85y0Eevbu1Z3I17qUg6QF7Wt8iC4Zf22iPr5F
TcYo/23brNjHoZSFLdynDHgHC9rFD+dGNwzoXurA/dsIFbYYKSQa9wFRIxlIwEJS
NeXTv+qWnLRHk8f+LdazFVmmjMiydBqgkXOMY5dNeg5gRK7AF8PqhFtgJ2LV3hEH
VaP0NgcSY9S1QS/tiEE71yiR89taTjKk20Exgp0TOctzH/dHeEvgxxIPD9bYEETH
2ivX+Cs892I2lYGQeP4l9SbRgmIi/c5gq7oR9PuA7rhK3pljsBcPSJpa//cLx3kA
FXu49LQfmabPKqdpaZTP0Lg7myInncTJyZnhgWlIhbi66AQ9xw/T3a9re8r08SGV
KIGHIFg4X49o3arsMItCzxCeFr0IqQfH1hKFvIeBSz/Z4ezWLk6A3MVRMkRNncxO
iOib8RQdJhWBP+TKl1sQpYSo8+eR9p4SmqVXn416G6PS2HJe/7N/WKxc8DJV1MqA
9SOMzsUuq3CSk9+M+Apq8CJ1hrd0juNubqxucu3drK3auYhfLwhNz6dCKVZQbS+G
T+wH+q7xTKxMFXwOa9pBxbo9X9S/sPRQI1AEmZwT6IzbTyDgcmeBS0EoUCdyJx9i
rcJQV/W6rQyQoBl0ufbG2S9IrMfIXO4AOvThRsQJ0M1Yn4MKAgjMU4N0l+2HL01J
ozQqh5FcB+xbW3i8nevV70u85fYyN8n+frUTC+PvAe4wcLwKgM8zU/67p2gj5dJ/
slQAi0SWAzW2yfvAZJwql2OLodr2+ee7++4Zb72t2Nb2N9x2EASroQiEHTmkNIx9
ks19ajcEP2/8sfHc+VG/PehfcxhRgc8NQFqMzuWUb86G7PPJF5d1RA4ASSteCY/f
7sGO3s9oNACMvHTQNKaCWLuOc71iLqnFMszmpzQSAfLLtbqtQ1Ph6CEjNuE5IF7p
4UrQFzQejBukJQRqZJqa1rFg0p9eR/3jnUW73vecw0vXj6+V6HLotzDIMTwLCuH7
BKJ3Gozmq/dNel9Hu2Sk/OdXNh/HmOVKpip5ck5J+yNen3Sa0GDs4bMYW10N9lce
9jqb/T0xcteSGV0Z3vU0QjVWB+GEaVFggYf+n7uxpZFABE9RD/G5W67q+Yoi8KHd
r4eWssA6doPJoLXcQqkhntzuE5FFcz3GuXgysKN7M3EpCBAHFpAheXiA2aUKrvvn
lDzWhY3CNDB4o7IuQARQpkFO7WmRLjaeziTq3AqUwh3Xzd16M2qEzmj08t9LrjzF
QWktIWxOj1L52Ult2A2zVcPorFMO85WlDYpF+B8xBW+U9o+d5gcf+DhkqOZFr5fb
HZ7qYNUx3S/75ZyKmYSBMwb3Z/YAZp41mqxiKJkvAbQNNfT281W0BiV78w5lAZ6B
a+xMQdW0FTYap/RWxxDnbMSoleIk+f1AVYcagLFmLEyeagkV4WNE1YG4oJTxqXvz
hKKwB3YGLPshB8WhQzJKyLezqRs1eQKtmLQVlrvqiincixR8ad7gJBzebJyupjNj
Ow2iaW8TkemI5fGihFFD0HpH86dGiSrZDNdbIq/z0TVB7sz2BQybWdGmnq1+tjjq
XgYs9m32WVE/IjpIlrSVm/s+3pb0rNKui03aCz9Gv5NMwSVuTNY4FPKzqAmiPUU6
LgHGiVJP+DaEcoDx4WtvH7p9qU+wEWo1pX0I+uzXs7i11lrphdRP47AtSj/Pxzg4
7XArcKKKsD0Z8D7RjEL4D0VAtgaO90vxccymoTLFuamM7GCvejDXJDX3PMk4MmH8
NGqIRy5JoTzy4ATMiCjIMZPBGHftHs5G+y+icFpN5AyE3+a35JV2nBc107zs9G8G
hZ1BXT2pPbQPXk5hAPmRMnsudPmvXOcEKGKIw2GKYdoLnfsEALWESEkPS4EEKcsU
InjpW95o8mdf8MEZlbkUmjXiGhi4/cI9iKcof8zcpUNdOyFzY5WDLjn2kDPspkR8
y6LpiogjPa589D+Ga9dLnpJdcCFE0inon3pmcuQtW84DtiVv8avhwX4L2zC+PAcJ
tKwKrxGZhuqLbUsWOod4F9wjl/9dK1D5jdYh5efCFK+u5hw6dT1r2q2Ro8KDOEFU
okh4O3qgGQ4odxwGhArwwuKOh5z9ZX2EwYhMDu1DSS7JZssw74z5PTKV0wu56JZW
QhnpyV6O6DrlVZLgAvdKQE6Of2L+RwMLaqmyj4q3X6e13/OCs/1hEIo1/HthMlRG
DqeONBRTLHKFYTRqEVGiiBXpBfZfamzk+CBx8LzssF1LNrWsxvL2av7gSMmfEuFT
hB8PEL3zkQMId6yLH3S/px0wWB+UOvr9VTQvusPAloCURzqL4U/WbLErmR24d07A
CfbuTfSvZRdL2bSJALViSwVSEMKad36N9Lzr95jbypKASeoTZf85T1BUNcOJW/Fi
SY70QDC7PcILpX/FoCKzsunTiiVVulWO/57oVytYifZY0gTShTILxPAbBE0UvZL2
2lOESbf9XdYuxDh7+GEgQ6AjxkGTQ0f48cUQkzZYue4NGEodiu0/AT/CxcZYDzjb
ZR6uga9nY91PlgssxzW2NzYXPz3VnKAsinbEr1wDAzPWadQzgH+nx0RWB6U6I8zb
S9HNvfN7HBp+onkWVqtyT4I5jw5zz7jFiSzgBmrALOv9v55o5RXvasrDQ476cZuO
2n8WiqOO2KgQKopUQ3pKfFys8LRXO8DNBq5xzlk4gwn+u1DAL6xjyq0OA8n7AfAI
ugPoNNbYdecwkEnR5cjZjEfqdK3pOxvTySppDJlUD+VeCaFoS6b7Sy6snqGwO5xj
fgBwxXWdno9FrfEaQfhBRvoYyXnuA/cuftMZZfEQkvhMgBGDlCm5gBkjZIAFD0u6
fQeRZyQRZZP/LXBiGyulHBpwukNBdk3CulCJdT4LqYcHU0jrBeziYdWWFPgmelNa
r2fAnam1zf2h90u/xX9QMgpJ0yfsG6CGuJGFAPsmcVUC202aa3H4gzGXH9udAN8b
CpP7W3hYf28zh7wLYhYg+swVCsEmfI3MJsSYqkQfcc+0sVyzVBcVzMN0ZewtKkmB
nBKS6U4yF03KYfk+PQp+r5xo59tAXFNOr529x/FtVteafiVFtf9nLuvegskq8Tut
cs7XpUyS0vADLH9c7zAhBZBJmkav/SVkYyd5SGCf53dsON1kjKydt0aZFD4a+gG6
19lg3cezJx4ZjPd8iP0l0R6NNDSoKEc/sYF8qZuLp2+uypxzu33pOCxec8dhtX2C
vRFuBoFmlTLtigQGLCKuyuHRgqJ0oztgTGBdZ2WoOnczWkUHtXiOTcJAVC8dcKIX
JyoModsC29wqXqQEeZBIN98NqV7/wvLjt2WF31Fq5BQ5xNjFwA8DuDUVScSY3E52
ZR4sO37uIAvGBld9wiXeWwfcMPJS7GtvbCbkDrtE38r0m3TbUwd3RLXoq8OO6sA1
B1pKzyuefVtc5Z78DPelhxUljyUWCogB2J+fXYMNBP3hAgVzRhaKmDZDuDNATmWG
XZsrwHf6ZttDoUyrI2rLk5HNBXaSUaBFRXpkx/bcLhkiJhHhswTSkj/5QkUbx9n7
ROv2Xm4HHoLNLwcPJ/7sW4NuBE/ak6n/nHO5hIcktX4Px6v5L5ImxU1McBsJ5N18
rCo6kH3XkCmAgwL3oSYmXC4fowrb9llYtYtnWbrH/WUx3FWc0fQVdbp2AjYubvmN
WvdUGI5AARj2GGHW/QDnjGIZooC3csF5FAAjgi7HUiBKA9pYucBdr6fEkcUbbh4d
iAFh7SnZ0Ek7GAX3rtIZWqe8im2vjntlFUVIT/hhAAIhcEzC4LtEp929mgfEBhEA
EZtyl12+yFwWXyMrT53IIuuHOm6sUswjitUZCTlK4frfhVAvvuvB8lGfWWnMGyOc
RTrjLP1I3kj6iMT5LQmhiXvetEDMbWe6dp1gaQ/pgRbrNjWX0uEThknfVohrNE4n
NA2/mTA/fHmw1zAzPL63UEI8NTHJ2RrD56k3FxeQNZTtQys42lyDnhxFp5/eq56X
NGvnNTRY/js2fTntFVWWQXZL29u4QO6CtrMKs2uO3hN0dupOifHg2wVDWAa0YYVU
i/DG/GMxFrj+PwFPIZJEo9pbGfxnUO572V4z5mUR5/wCny+ylGJmxW51QChc+hrB
j1p+9lwaGWGBf0zBN3rrP1DgN2P2wC8Cih7TQdUATrodX71GLCsE7DWWKbPuI2XB
aKIaVR2fb6B6FWiov/nD7lVTljzFMl/exNDFpa/7znCP5ZYmP3g0Vv71uFzW1iD9
1iKOchO85OzTZkdvt8+y4QBoZQNHqR1fjZu+QUCyogd9mf+RXVh3w3fc7cXWqJP7
EnV+nMLFvo0/SHaXvEWMunip6FLkGvv5mUix61j/FRsuBcro+KhGMnty0v2beolX
ae19IsH4k3plQUZEvr0/oKq3ru8CZhjcZ67mMVmSg2QcNudnzeQafZTBx4Jv1jgd
CvnEcuTfioxC1WC2Cs5ttV2flcRwplximQMC0R1FTBc6MWEfseIc+HplMNVYV5XB
a2DQvgCzaNVfqKRqPTMJbJVptMkCQ/gc4Ygo7OH2KILz3cnTcu4D5d8rBMQdeU/M
2tpMiqDuiE/CyPxEPkzTc1tw5frnofU4gEoNkcVE/WQ9K8OZJ61G64aH/5rm3sG6
XDPMOy9PQcHldRgvad7hHWodIXjqPlkTHQ1QVlwEqi3Tet4Kf4fVKZDjOXdlbARJ
eoSltkm5MpLRv9InBusux9QhQQ7LEKSyYkKuoYJAeEWJZZ3Fix5l1VdRnS5Wx0W9
z1MoKSt6mR+h+3sbLCocvriSWty4cRicWpiUn5yAVJt6o1tOfF6QFUzqlzfE8BXj
NvtMG5NzXMJVTt7TqjRrojioedZyd7n4oTY93AMAUyetTBL9lq4d/PhPmnNnHbRy
KI9I6cmQCRGiGA0NrCItE/KJimi7pyS8cSFbSMw6z2f6ruH6MIY7YH9SWdD5Legd
6ASG1cmUdQQs2jOcozwETfnWefcVnkXzC5Pd4NhzhdPAQFb8g0XtrP3O/9VrecRF
IwwP9aJD2+1cgjfXwnw5YujVBkbhz7i9Qa9LAFPty/Z17XH8oDqJyA6MV3k28xww
IN677Wg4lykXaRtb9fAxkJVwQj8eDzzmK9CZ09Vh9pwiQ8WEpz6LKGIuMCJjqQTj
qM79hgnbenPFB72eWgWS2GdqEZe3wLj1411fxKjkaxDg+igGvcCtLmUhvWNxyT3i
WK84GqbTq28yOQ4sn4apQ+3wls+8k+W68yMzsADfVhnJ9i5I9yC0RzsaH1gfdRLK
5sp46mpDzyhKTLIZVdXpRS1ekCRULZ6JSWnHt3D5C3tZhQKSrtYHv0KBdh31afVK
1oKoUR2A6qj7sbkonVJ/CBROYY9Oi85krKYYjbpB6PuNh7ZMqkJYBTiELqCRrkPs
HCCYNu0Bsp2b2ekk1dQzJovdTWo2Dkn51xMfexFLqUn6FwGe+3bTlFpgC/DCd3oQ
+N1Td+JC9tMQ+mqBLVLKFDmyukzY2kAdL+T3XoTH2PbZjBoDj66fcWR8V/2hflTO
D4J/zghcVDJZ+4Hk0PtlMyv7JoxNIs0TEyAaVujb/bRqlryFKpjrGD4lk76cxhBK
r8sXMniKlY6igHxeUCu9vwazetHjBcvM5VO/0YCsCUgqoqkQhq0A+hBfxpmg45cQ
7X1PndOgCmCVsrQS5RKX8V7EkGp8yFZ5PfjyfO11nz/FNQN8oZQugQ+gK2JH9JE3
TZgOEp9CDpZEpnpg8EMix0w1xx93+kRm9liGp+g16zPP7dRMuxW52ZKFabEG+BFP
iyrUSgRusGLE03EtGegL3BVswTRYUxYslhQoJTFOYhEJBZXLvOdcclRsbotGDc1D
6FnCFZS7ntbRs7KzPhu3aEIIO3MQMMYATnMc0qLrXa8UuZtr9cp2+QBtwbeH4Dcr
6OMRLGpn5juxti01EQDuqPzdCxiyk8LOm/QmSoSCHZP2FoHaMmnHgxfCDwg9K/YX
xDAx8pKaJDVMaYP8cCREZlfb/ZydyfnteQzppXyr+nl6jc1ptSzHr2OCgqzq3RLf
7+5ej5A2Dz5C8HSPf1vWAAYwZhLvYcu25uxO2zHUvT0E0P/i56p0dpxVBNL9pL9o
OQk9DaQq68obyP7GFXFuoE/QtyMG/cwVhUYn/cDKhpOyF0eoNfhxP6lwiDK6Td0s
S/qCGd5Q0jMEQPvN7x+YrONgeipuPRbLK6UdPM19Rfvk1dAU7lVJjyZrVfjTUgBX
/Hs2lGJeRTJA7r3dkM6z/rEmIP/8FfjLzZzWyTCRQSShd84M22e2IFdw/vVEcbMa
aOV7PNGZnz25V0LxdZvnd5iQJ9WIkm1P15HoM16FiEWEI8ftfN7CZ1IidkM6qoZX
hdFu+4AsRamgEO6GS61bNAsp1F0hCxcvQKBZLF1MbexFCuRzoEJnRTqxiuOwwxej
HjXLm7r4t4KG/UdDySZ40UxbWu80Hc5t/72DFPm3YWPQmY+zM/0+oNmsyfSM+Vo1
8PYREgEWVAMnz3pX3c0HvjTfISUSomZBbLgV2yqgvL+RYiI5uM8R+18Xl88gSl5p
qkyQ7lhzEeFaztpS6pA98vogJIxcj2cfwupx5LtL0PTYTEcXrDrZh7MusL9PR6RV
atkmdB7+ggTYON+VDgTmUR/ByCJWyigr3Zy4cIy68BAEICglXFTGA+o1veMvUXEp
JLBop0evc7NZCmKutM8EwYEWOPWqlMIt2pC/pOjHhngDY0Rn9SZEVOsC5WpfQJWd
CrXCpLmG8/cbATE+RgKGi1hGEh8TPzuvaYGE0nTy0dEGilUdE5gpqSWa/+/e1EuJ
wh3030ctICqoq92pLG3riu1NXcMamCLoUFXWrw5mL9PjV+e8BvkwDps8+uzewWAP
rY1wB2TrEnTKXBrGe7yixt22wyNXpyYnRhFg1+WrmukgpY+NqyzUG32htUd1b4Kg
NeQ1/S7n8FGxtcFCVBBba5Ta+PWwGK/0DRSoPFpZYVtgiAeDrpyvDNiA5ab3DgKZ
2OJ2Jo4h0K8UJ3z6lGyrFr9kdsjB7nqVQvxaNSebzgvh1fMypZ33J5xOsHmVCbCb
EI054h1FUql+SWZBZjPwpZTzDOAnyRasbPtr24626pbgICVsmZ9uuQPcSbmZu9yN
xoq7pWijRxIeKBr1PFsn8kitOfAvUELO3UwGHReu0fo6aOjU/V6EwYCkMefmqa0h
g6RuoMzSnRpFz+fsCN8mAW7Tp1gi55pYhdF53rAxUee7Yni/FDzT1N04UTzRx5+T
sH7LPRB9m7HUm5afm+4HT7aNNe/8Zjy0YrHeE1d90aLDmb/F84PWmbKomKQTBj+E
ORDufZ3xZ546u6PSuxKDYFgBkMHxRsRZxCO01BKKrbu5V3vDtup+lpILxporFAgP
3LydrHtgMy4lD9I70xmL+LwAs8mykUjSt8hVPNiE3NlKuKTB7fSo+tHfWLItqJEU
eblgZJmBI1jBfxtHvwTGgN8NvUcDVNECaWROLTamGU36S+tJ1qGj7jD5z1/iB8Mn
P12QFZLZBH/HbJiJEx601z1zknaU6QtxWpFnHDD8decXyHXyvns2OSu+aFlJVis/
MXTXH9ivPHdWAAElt2orRRBBchrTYYO2ymUTwL6FR6aPH9FPZ0cebNobuP0q5GCa
enmZfmfYbMN/IKKeeHlkS8KnwZysdl+Jymys7JZOFo7ReWR7l/6ddym/rbx+DLDr
2Aely42ZK5hKwmZHJbm8HY0xuQCroLNXHXJPgufQIAwNNUKQa8RPjiLujT2k+C8V
7N5Uu52nE0y94yxas/KqAj26n68aajzrLFHLkJGor++nR6gEkgMWlioQHzFbUrQU
Ab+x/gN8QOfnVwEe0yOslH7MUiYOsNOgs57su6TQSR067RtzRaf/Y9MClefEiuV5
TlQLlnRdd/Z2XNQ4U84IjhepIztlBoJvhvlAHOkR5u9PF3uGN3pTjTg6XhP0lNHA
PVJW/VJGkJ8+Hj3MQc0Nu9wo7dAsGd0K+YLPQVODUCut73xhBSZFZNde7G+D6Jzc
pOgwDhkheUwxhjaY+fnPN9V0/KDtxCtCVcQR4Rd5y2W2FtEAE1z5pcFsQuqXNs52
KGZmp/ZzI3EINfc0aLR3Ib4h4hbDFgzSpG5baj0hWcoQlbUM7Jy5LViVEng1gsQa
UY7ONz8vucs64IUQVer4vTDrT38+729c+AitiEmxLSQJE0RYeUESDTco096wzFCL
gHTwPuZtCdjpdkCvYPu1rCoOlIA7N+21XpXse/QA9Z8QW4bvbp4FVsTjbTXsx8jv
XUUOsBwo0AqTMD3MDCiQdD+lI6XFDpyB58xwFO3Yvg0bWDdsyyPidmhfd9QHGRBi
nebCvVuG04Ce524/OymgM5kSyxzOhm2ko4D/cBRyswQJBlrFjlBIdUhPKenvznDz
t0T4+PjxABQ6wHZtdlrgz6ygFMB0r6DJxXRN3cqgWFZIbvoHeipjEi8ZL3kREA0R
mQHoU/wKcEV6ohBK1od7B0RNCmwiTQqVUkxRCQRiJKMQ4XiGR2plPozhovfGz82m
6wcKrgitMItEX2zUp8mSe3c1OL29mLsfkAiqAOT8H/wjA/e+NmhEpe/IS+OKMQE8
NLEp6ILZOnVZm3uI8rX+zNBIzYFEnqSMQDkmi9D9CtCfLOFYkdMyzZknvDR+cPFL
QT0JKs7wYWoiuby5yl5+DiaOzTg0Nk8fmk91UGkqFMU9mUxZ8jArBMgS85t2dEhp
+91gltDFo80s9VkW+t+ldSwnRf+oJoKHYh7Jc2xLp7iYiaIrTRzWgzEbFg9i7Icw
idLkSOR99zAtkGWlyE9nLq2Ib2SwAJCaMxwzcztOef/YvviLif4/Kq0OEIk97QsT
+KSmForRKyqqJsJrPe2i/3j0fu+kzrlCyx/A+0SrHkWvAA/Yy77mjZk7gyRvZ8N+
7PH6uxkXwa7Ekyu6KQ7XMNTin6PowqOqMO/EJPorZ/fp9PfDKfOK8D4dE9kSksaR
KIaJWJOl/MS1Z3X01wkmkuecABU92ByY5krUDIi6MaeNvJ32hUafXx189vHtD2ff
BGnGGiQcUGoOezBJU+POYHD784EWKRYLNKk7tcg43op2RHZzJMMNjDt+WceVA9Km
bbdiDCIKSA/29hAqLhKSozhIbVKzzd/RHmM4m2ka3fA4jRQ86CubC9fgnS5C0aGP
psmh5gIusLPGhw9uCo/RRlQqpPuuq6i8hT9nOl+M36SYxeD9wdpO0Z1tJ/Eh4Hxm
Rf2y5+BWznHV7f8RZS4kpM9/5qj2DQeQhEa0akcYeWCCIvjf1fCoy7XYmmPNIc3c
WiGUlsaMgsB8zOjrxpPdt2VMnH7wMU1/BA0wgihyfILjuQISwn6zE52bp9JptrI7
VERyl3VardyDIUu4l5IMxNTXdFO6Gdxv8IGplgG4eWOHLKW3uJU4wgRU5Wh4xziM
lunIWztbJRjTgZI/YUXKCN/E3nGzfMhrp2AOg8bdZLlOqktXSjVRhhP0eV+R5Ez+
zTodFdhuQlf0/ReZQh4SM1DkWE1mW9dEsp4F4Q/0otIMjLij/2U0q3W8GsQnz5pp
noLflWQJCijl/r4Q8nPg4JgRVMwFLMVMhoe1XTa/mUP8n8mKiGGNXPmC47DDhjUn
cGWJjIddRDAqX5xupOIidunbVgqxB7JT+YKSLSS+bjfa/Hui5RNPTjGb8tLjXfWy
+8FatadoZOyfud3xvUXkNxp+XxvIANB9Aar1K1Ftu62zFN9Wh0tZKmaRHDd76s1W
YR0jFjeu3iNIcOWqR8y2F34i4cQXBbgoWkoBHvKmLLLTjrAuigDZjNm6OPHAq3ZV
rRWmkgLiKHmpDn5c9I46v/xlcWCecPUcbK74HsoY0+3zDsVNiUv7MJkOazmHH6gE
v/jfcj5/phpuPWEukPdF5lzeUjfLbTXts5ERFaKMBBDPvXGv0cldzQwNIPlw5WUq
TraQNc2lwJCBK4dCGC/946bKB6+prmUiBMo+izsFG6ZRpsJx/tnWtSyw92IMFOdQ
FPPDvz1Kv3Vwa7vD9ATIGuNqX8UAiB+PiJ6fLxm3h8FQGjTLuXu4GwLZ7sgk30Tr
oN0AlgZkcroBxaA5W5U7A21KbWMP+fLudGdOqOTJniXXRe+UIeSt6JASkPSqW1Yk
q4NVRl+4oH1hHpJmDMkje2zoskONw3/g8UTP6TUv+ANXhxJ2h5yXT6ToVJ1dyo0B
Su7q5OVT19pkqO0fbHV3UfPL6ILxXkQq4bc0iXuRosIPud/yO8qP+jlNeDjZQOW7
2NYM+B5LEnbtMVQzqwV+QekKQe+l90eZub9CnoGoTGfyqfoPpsbwFrLEGdzV3+b8
snYySgvoNy8wooY017+mGRfBDqn2dPB5mATORQ3lRGuB8Q6YrWTzYfBwXurZMYhn
fJl+tT6KEJloSzxVGEio13NpJkAJmN2rXydkuKpzMiwqwzZgQLT6ecReOEfWwokt
WLJuql/63lj9ByN5Gv77QTMfhFHCL6RNH7VpFyT4id3oPdXs97gqMI1yz3Z88Lek
lgDo4ls8TDP0ZVOgPo6/YmG4w+0UzIdHyLWYM2AbIBR5OpzrtXat08j8k9Lyp7ZQ
BTn+pvwKLqC5/8j8kFe5G5RznAXDwzxttQ1SO22gtGq63qdJIazt6v/MbQbOama3
MvgfqAkY3rkhGcqCx5YdDM6fvfEtLqbDu6FJxNx4tXsSrhB0ohBLDs0LZPzSa02j
oYGZnMgPpdNF9k9R21ZNP/C0v5dFuwFtiPi575gy7fbnSoNrWbPgdOjNOvmfZM45
kDEeZUX7j2bSQNaQirQjjBTpqKXw4YXq2e1jS4+bBRfkduaBCYCyFiBZrM+QZqxM
fMlMEEpCY78adPjLZGQJmWolYYHr8zGKHgeO0+LeGOneouV1ZSynYzqBkELXBsK9
e/R950D8O+WC6xjXPpILLdOCQsySjO9fRPFdN7fMBnNJrC6a28JNWRLmYI8lw6bT
ulBcvviN34aDX9EKaGkEInnvRXK56WZXAWDHdG9H5FroPoZMaz63Hsb8skTSVSVE
Pf3HjdGH2mSyuHVlOMnhsaiYTpq7HRpQ6WD6Xj4GL0LDtsgnSf5g5BDgFXs7Ox2b
6jIllkN2wl4cfeqtjEYRLkw/3VDyMAbXkC3Gb2kmaMvgaRiH3TyW2H8Me/3mQZg+
jCUeWrzQlv352iwDNAFYlNsy15l/waq0V7QkEFnmHEV/12ce1EKY7olXbVJGOea7
30uu3lN+2g9r2y78BgQY49CN7hKktcnstnWqoloxCje4dL5uqwU/HHGuPYmt2aC9
3hJCuI5YrkTVXT2dTQOsbpbQSXUA4SK3j550Q+lr497IcBpKMakYeXQZw0tXesFy
il7+8Ku5ZWin4x7t1jdLr0v9Q2R3/oUDqKODI/c9YmsHUu9+sgcqDMgDSFuZnnv6
9JNS139PbqGsERAdusJi2URVksBb60baGm/P9DcgSnWIRtJfxgzR1GDNULVWM6t1
WyxDnQxFroZ1wWYzbAAHu5pcs28wHgxO2OOIlfr/YhlzQR5QwNpuh6ZQHz2GjODP
8F2C/dU33VvEbH21E3OkIKVzWaOWAdaU2zdty/CI0YtpV322+AGG4VRbWVdf7BBv
ttFIdhvZ+wq4naqsFCYzeDo4fZ/nr3hXFifs3kAP98y8MJpwAO6ugFMjA/Z8yC4B
iN1j9UimIazG8cWKecZUrMFKu5pBZ+Sa+JVKqsGzSi08jSL8Inwcx6jVRtC86orZ
ABBSYgDD4r7E3KTzX/NbyGRXuMXWib/9IiP2lVpKKuqBr1x6UocLT+62PLQI8UeB
Mc6x5XJJTaeILw8W87s4vNM/tHQdG2v77nLPq+LrJ/ds1PKW6v/ShmdsglOclY3A
LC6P0M+Lgv7u2mD3SXKzTO0kFsEo2mWjBgz5PLdPlx/7xjMDSuQC2nwUQPyLUysw
21LAZKe8rGrSsRiuZzmNPgYVs0wkwzqBn4qZIjq0+TMATVaD0qG6vAIokeEm6QcD
mw8APIJ8tZNYEOrB3uerd+N3ktDaY1e0CBIywf6AT3K/0anoFkGf0J+0KVgg6Xsv
EV90sAfHFHuA9XstbNJhs3THZZM5B5OUv9HyTbbsBTkmirGIhB0klK281eJK9OYs
kuMzoECDGrdUSY31nigZO6CGifC6SJEW8akbhPU1IsQnfYTPaz7gh5Y1+yYKLkoY
26gNm0XriuFLgLhOYics3whaB4IvQBXerMMEoYtz69t0hXkWl38gqRnupRAgqOj2
o5uyDo7yj7SwM7lpSMHYyWqwpciKETCzOoIBONOk8c9+MyAr+poGeLAlUI16Dizj
bTavYqY7iRWYkihOLvgNPdZQSxax+SX/dQaI4Sn0gVUbdxfeW2phHrIuk4I7tVyt
YIsHko8APB4d71MYkGCWDi2Cp0qqR/ZwoPQqmuuKiVhe2A0D/m/7xBwU+/K4x0WC
djv7/sQDK/agRsiZ1IxhWb59L+evLzK8730cYN4cA1uWpO8WdLHPDW9j8jPDjChv
Ns5JHBm3C4LJHF8CB+BHrDWCFVbm5W8R3ENyHdAMV6i5sH0dvQvuWHv3/9me3y4/
Zst1YE10SOg9yLmRCpFxBCP1af5GWEK7ewiihnxpY+4arE50vRfLEQRoTAEHty3g
yEUWL7u3HUmhFzVzV0U6b7onLoD9Fjg7BSkNZduSuAyQgsCRZZhuuzmp3cnXWHV0
gGB5F2uzUA1EokwedRCjpXiF1IoNlVcnKi00fGqr1jd+8A+QjnJ9n78nZCPOfSOd
rLDru/DXn1gewvAP/PrhN07tJx9Gaikii0rbb464PNk7jk3wEhMzc/yAzqwC/CWi
EsR2xBNPbBK54CcV8ueaMEDnAyR86AfboXh5oziBxnjgF0XeLW07MMo7j+s7hZnC
GlZqJhtV7wIL9tkX2AjVsQ+DYL9HOOovs2i++t03kDld1H6Nr/rFKSVXjG9yyUP1
PyjU3S2nUongZCBarErq0YwF2AFsO8yBI1iMgxs3JXqaHA/zZ04f8RJKZOSr45Di
84LswzLkc6tRXbm8SUD6bUMgxC3mOd0fR8gM9o+63dWEi9GcQ3ZbUQp/V4XxC+jU
L0v/VteurAFSNSmFVuQXkbKBXCKz/6gd8kx5s9iVjLdeiT5btIOnNRi7XRbP7vy3
iXXzRdLfQbFzylYBdeX/OxCE5FtM4s5AK2mbbB7B1cg2gAUgYwRJRGqX8unRS8We
fmv9WkY0nI9tkQ8YcrxFcLBsN+GVxfQkI7lB0JwrrUHweBDMaMn8zrmE4lpwCC7m
2B+FAdSZ3rzvC9aaWnIUZlcscj0vWS7+8R1q5SAOYQfwswhbWGT+pXTNSvOdhbJg
8zDoHULNxk5R6XIw1Yen/JStcl9AmpN4GwzhJo4m+uKz+4+NxPYqK2rrymmTCapo
2ODUkbZngJkQrC+24VReFeoS1w2BIQQmAUKzZrXegX8ZAmDCpzNfAVrO/3EKj7ZF
fnN1CBGqWfGn4FLoqZSgG00B87u2JTJG9LFi0nLrPWA0KhDs4KB0l2DVj98le+v0
EPp73WAFOOLZmODwEk5+hwasHy4O7ldCT0cK7GY4dS2O5ytvQWVXbiFem6ZJvuw5
32KKh/2RktG2rezfRQj438kLKEcw1N6oTw0uMmt4hQVXhsWDbiyATQu+IXhKHsqj
8PENkIoXKtnG8zFQH+JsBwRpU6J9GNtAjlHhgBBumvKQqy4DazG7JM9hXKdu+XiX
/Fwk4FlGscMsWSPfh8ldfu51Pw1a8RHjFQS3SpgBWLojpcGV3Rqe6c2VM+H5Ql5x
Qtrw8n8fkKB7GMeG8MywUQM1ZWhvg+WPbD3owf1pBhgwPqsEmv13F7qJuy7bFpie
HnpwAfUVq2HGJNDlJGhkNCuA1NCNOjiZ2nOPpD0QoT7SMXnshPKmY1omkZLTputf
3YNyxEy0ax5fSXQyuGkbnQsfxSB/kNEBXSJjwNU7WX6XvBJVcOTIVwaRdKg2h9p8
O7TAxPp4gRtApza8MWsK2djdVmfGMIWdJxK5X2EYD9HlCN5Wa3jMBMOah8i0bOu0
Hzgc9CUC9m5sdWBWi3p1NKcEtNAfEuTXbgmppPdC04Hgc1o1hqlF5zFwAfWkC20Y
MMrAYupzkb5arSkaX0yo7DGNRjoZy3ibZoxu9bNZBmk7Z4cQhktsgYp0lZ+dpYRl
zx2Izr3vknt3/XVpxiigbYbTgb6dmBbrmX/H/gGuKsnuXUcmJcx8V9Wav58vZKdJ
g1yb+kXQiSA5rULKwgv6L6XmWe+BR4L4mOEcp420k9SXIw0YSDEWh7Fh86dNCOaZ
iruqk3h+jI/UsRvpVWB2HU9YyzVod+EBwSd0Ek84EMunTr5zCv158Co3ZWM4e8gn
SpJzFCs/dTRXpagA95V1ryAZ6lQfhIPBHmRLUhVLv0U3sXgzQi9ag8noMsf2eBu1
8uu7561hQE4LIBL7eX26J3KdX/LprZ7iFzt/Fiptk6aa4HDySS/mbLfskyQXwq68
ldKRdMOCzt/VIg6amuK+cnxqqvUoAUwzYQrZsOCKxlCMfbEs6vNPmi+nJg+7l4XJ
WMfPAdU8h5YBl+QQj7Oz9EYBXwmqHwWjGpwEeot2njrADvKOiVDfPX0y6CwsyfeF
ygr5r4xz/GSIxBsLkO2CRxevzIDlEmFM5ckV9jYsnoNpmsas67bz6g3CArfOQe8Y
XAenJ9t5QsBnJqTSCCamwqHbEoke92nr1h4Ej/WLM8biiLtA8e5EXumthQnLT5pH
sTQQNcICH1jBCfb8VFcadMhXabBEMKKrfuZMQMJ5VAw4WUDnfQXId40n3piVUewF
Z64qofAZSzlulXsI9mqvUWakgNAF/p6hVEbXzD6QPVs8zJ+Gd48RmLii3wZhHDbU
PxhWkO94nBIHFOcE6OYN9x1Yp49orjZMWcNN6/0d+nTw68MsJUsn1eSX4bgIV/Od
zz2ewNoD8yudjLBtCiAtxvefrOLlmxJksSGXJMUy0lZP64VmSV47OiZ0E3OlOz2f
CwRd8yFfngWxjV8HbSqLQzcfD/kvymcChrJ2uqgvHhPYVfQDraY0SNa657a7RVHx
VAbrQUL1oqmKXEpDKxKvKGYkmie3g4fyRBJ5coQhi/RZMhIOv61ygMgYuhcE81AP
uji3RYva76uM+TcBVckd54NvJGUfM2RICk9+y6xKtD2ETljvJaCqhVWyj9QNeFjj
r8bOf9BvOjR2iy+SrPGfsUuVSaeb+KhmtAcDTIU/+hc4XWBQHGRzC32bbCUgNWpL
oJiSM9sILf2oeOT5k+PD0qwQLFs0N4K2rydnwwXDXrJGPMvfhDQx6sDJ+VzDJ91X
SaLWXtd8iPR8VO0xpLD4iNeltvg2i0n8Ijq5ckiDO1zETw27o8/MJzxaIJkg1uRI
lpj4FDnXnIb5dIam0f0/rexZBOiWyFB92ThiYg7QTNOdri3V/9NUsLQuMv2tXMXW
C/e7FxYarkuipAlLEObC+cjWzOk5EKakna653NtULgfExgz89sHUYSsP6Y0WtDi/
+hYoYMymbFLKPsokB0s3UQ/vWp+laI4TQrqxpOdVS0nFMW2ESCsuXcGyKHci/RIu
p1nlx9hcaBA8blpfK1pgVsBfyf4OjWu6iPIuvH+L5PZBRJ02ClvIh833hSlHMR4v
8ozFB6qHq+7tXwwEX8lLRcVQZXitWGJ9s0Wo7e/nZsx3m8Ci0p7MKsA4blxrb/IK
uYJm1q6WioGPEnIl8G9DPxqWfLaC+uougRR7s94Xj9vfEoeYIRmOYupg2UV3a2xt
wtZP8xaNOz4fmqOh14oaMq7EzgI5uIgjQCW28IMRlS93/eTybUx0D8dxBp+mJN8i
B4oLPJQ0htSjAsnvm9Qofe0zjO7GgswOP5PhF3sQpr1L2+c93pbmB4lA1jCqeUxA
W7IHoUirYKk53t3DTXuWiWunYOKfgjSbK04hFSF5iiOz6vw/eBncmj79gGUgJpdN
p65Pka2fJYoXc3VfSX0bhGbIAHo06p2oU6MiffbYO/UAmtR+10rbFCiP5ym91I5e
UWlRc2neyKF89stUlHfOBqsPOd5oGrzUzQKYlYAE1yb+ODq3aoGOOhH4rBiwBeow
08lX0H+5xNxNG7GIKKpPDKRrc8rEpl6iD3qxmGpsRLD3fsZBvkjRecDaMeGzt4FN
DaK+RdqNcfRGKRDLqfvR7sOX1Q+5GsW2T2XTM7TGLrvR7ODoDpO46JNb/rxyUGYS
qHS6nZmn4bf+JxzAnUxpOwjQU3KoDkTw+4E2azf//goiXVMZmHcnJGbOEFQIFrW0
KsLpW4uc88h24kM3puZWTF5upCe2fpBHxn2YlXreqnFhdWE/d/cVmdE8RSy6RkqV
A3bOipcaeyWJezNPQS38xDcVkudlGIvcSgD/0snZLW1/afh1/FiroMb1UlFXTQmJ
5a1/4OrM0RF7S4e9TywfZf4vxGA/dY+4ohi2sxriuSK3IVJgKXlbgeG/1HHxjd90
DYT5ImSMlk9yuHn7+km4Xt0FS40dPaNiif5zvpLQjmGJpzBDy/UJs8kYbu6V8QjS
gjHQoye7BxkeNCGLM7FgOKMvYb0qlToqy9sKiRMIubRoMThkDYx2Lc/ZOR+Ka/LL
By0I4FyOO4/KY0iE2IOqYg9PQoRHsj1Ctl0yLmtlI8UG3NfsApOWQqP8N2H+r7b5
F+jrYXQOqg5XmbKwM5ZKcqwFFAMYsKZEAPFoxMWFlzurlLIno4AXsKy68ZLPycIT
q7r9QckyrwtTMyliPySfmBw94fy4cw50/mi3ZZ3rISKeEmSOyM+WWTGLqGvXI2uM
db0qGx+ZsNI6LHwvjOJYyTSnX5G8zUZxMEti11dvCA4u//GDFesMrqVhj+J+qsRh
XF3s1doGDHXuPxgWDlOotyoEJHgETM1+JTzvfiJ9zkVNA9BUksQbH/AE/iVCwZIT
s79249EmyP1hBLuPIm+hquW82xi4Mht1r+59lgs7l0DgFTazgpMwlyZxhSAd/OuK
s3d94s8Mow3Uq7AQ3GDaTgEdZFcPzluUng8jahrZDCRifYu+3sHir3d9KOtariOc
tSsqdH+WhJYC0NJMGtXhqMF9zGPV2iEmwK5TTrDo8lf5iElUULZ7njiGm6YA7/zx
fZR3HvHUioWMnv8uRWzuVXtcmiQfE0W4N5roFMpHuyqHfF8lEvVDGlUvtS0FrOOB
C7xYuGGpMDvBV/Fse1I4p1Dn2NBVohR3PdEybaWYJVaAMjD9Z9ICS198BpfLneT7
6HxUjsqKVWHGnvkMHJhGiICOVgsTTAE4776HLq6I2yY77y1xqdJh1mNicYhH0Mvo
2PFHusNmoy27BbZjJbVWRV5e+dppa/KVI8r6Kw1DqD+ve4ZT8Iv06n96yxYypFXL
4r69VAc9vkZPA5s/eQS0Xs8KbMQyc2rS6UJL+4rXNP9KggYyygOjzDulGX/u4KO6
Kvb6I0qeGBywBC/NOntQtECKKT/uAnaYTWwt72W3nRX3E6sMI6j103FVjGzcaOnf
mgXb+5L8KhzDUQaJVKf97C2yq+0N575kOJ7g9eTJGDy8JU49wgc/saz+lEO4Z5u6
CcVVd41P2X3C+RndNAHmcuJwwmedjXWDdOH4mg6kj5TUMq07azkhxMZewKlYGG3A
3Wkoq6PVliOOxypvg1viOX8bIKr+w7TrE3j266+TypWryIle9FGDrb8xdBy70SjE
24l5Aol5QQQzpkVCymHYyBA55syXkaw5C/zZ6a61w87xH7X/fg4Ilt2/KuEvDQpr
EqRlcS/fYEj5VmUEjru6svxzBM441cPtuP04lXWv3oTEXWMGlBKPG2bg0hyveNRH
CJhweI65cNV/SkhTaLbMSCy7En4TdpLa4G5w9WGkOOntktB+FfCuRs4omuwaSDGs
CaHdpD8AgdDJC/YmjpG9a9n/U4Ak4cu9kKIrWDQYvOHqh1a9IuUf3Re4NTWuApTb
p5oqLxwqgG7KwRRt+CQlktkSJRgeBjeAKQIPlNE7QpIU5OCOa7Tl25393tTidhEe
pYBasWfMskQvxLYcZlaihlbQmZH7j2kA/QrmONNJI9poyMaQvi7tk8i2EBWJoa4N
kUyrqYjRpzt/qqhM63fjBeZIB49EUAGzrjnhZrrCP7wDXSTqXbVWKGSXhebRahLU
IsIjympf7FW7GUFB/yvxk7zLqXY2IYQB5ZrDNba1ln1NvjR/izfS6gbXjIX4D4mG
Yn99XXr/1/qInoZDOTi76CqQgzYIWLkBSb05EUXcKLqdjux1qKrPommlavfppYxj
RHDUZ5R8iyJ+O0pCvxcffEJ/DKDdL8eMytZPInE0DkGkQgbPh6WtYCO6FqVBRiQH
Ry3y2UXmNqYMBgyTXC5lEzIa8lzqZa6hWFhbxwveOJAgPjRDrF0SSYLDqNeE6QnJ
Bzbb3KAPTRCbV+wuqqPun6eCITZ1otu5W1hpBTdmbSpjMG607cb3aj67DUr8tT33
w/m19SJ3CtEVKFOTNPqr1ItHLLtQUph4YAaqZhEnkdcxfbuTZhR2FEnx2p9XegOX
RvFZDvgS4BwRHxtQxfydBs+DIcK2X1FqSkdz9XNIdrmGbGXeucye70fVUoo6MwfW
/MeZ20w/xd1WCD/+v/YBDT/clg24Ob/dy9m4CSw+ObdT4LPUBYqSxVYQL+2k6RQt
TlxnHwf21r3JMsVTCQt3dfz2difqxvjLQdBrWHm9bYZ5z99FCXjh5mkBiyH9xfE4
7eyji/TXOUiab7nZ5+NFGNWsVdZSfz4UB/w5w7ZeuerL+wW9Yk2pLGz72EAjzwsH
LZ8oUNjlpej/vkMeTm5fATocgdn0QSr3IASjeWXQ1gS82p0QxjaE4xbwNu0QTAOP
uJalMqmkb6Ab35BPimh+xTJVMkyumE8Olxhi7xsMIOafH6pgVKuoAQXziAYoM5mr
jctFZuUtzXB+MCQwCksqp8ustMuFNpIttf5/+KZLbFpeARFEBapXxPFQxyEttoqJ
os6PGQPFKdJU48QeQ8ex/fjJnH/9pA6wR7FCszhdLA3BCJZzNdyxwxAcwxaCHNPq
VCg4BeBffcwBusAjaWveIejMCkH7OIS/6HOCtMii5UcDwVb02FXXgr5YRI9x1VkQ
zJq9j9NmVHBf0AP4A7hFE9UPZ5YLMb2n+lPQXDLree/WOJ5TRCGnLjbAjdwc/FVt
7R5KhPJZCl6vMQNo+fOPhE2ivE/JPp47yFIVU74N59BPqN/7n1onHXbmET+oIcAz
sUIo9YV3E9FKCS3StgSAyONR01V08wuAUakVQjUhBx1/uM3xjQ6nKOozjejk4ZH/
OfqfIaxK035S6o0jJbta+G41lywDJpJWVbPzL9RL2CgV5B9QJ3MXoG9Io4f3yYv5
+3n8UaOaHoyMdSDzACr529pKLsJSxY0QTqT+mvAlu5J0lLzQUcDa2xHDGZCsTL8F
IOZlxwkuSKCRH6cp9z/5yPYg2uBT6v8YhGCxjGhVBJ50dQlfu92PIpPBuxaJSWRf
RbyGRWi545U8mdFzPVnVZVWIpTVhwN2madpH0FJygvNQ6dvt1IfCZHUMwBmSqAzC
9Fsdi5k4YEWk7Qt7gH56EqS+kHZF1BK0y4pTDPe6yIUTF0eNvhnv/uuxZzoc0Llk
QB05qY1R3CL2qzUE07OdXfQrltdbCp3GO6R2CBTy1fyyniUGyqgTAnql0QK2Vwxw
fuaa5oRswfN8pjg4Cs9IAs7tJPC0FdtTEmZD+pud/nOkDiKgMYmUXbcNEt+lFC2V
V6aQIP8/laAOAXxDCFZBsK/dOKOjpXH0dd2rPY+Cl23rh2EKslxh8C4yqhmMYGbE
u8ZDBfOSoXm4/unswdZTnrzcSsguuv2TVmRKBFlxy9tkYiWQDzmjSfq7hbkeuVYd
NKd0/mtjFEkOQ/0/aI2njxEMXNC+PA4R98AWNtTCUYy0AQYf5dLRJ9IGkVUTTlE7
B5qqvZZ4FWG5wThkYB7HodAz4Qzn3Vw3dL2chKdAqFRe/40uBUH6VrBv89VOo6VE
GeRHPeR2+v4464kxnBKFgPTLpgyHdVkeXgPPWhW+11bFsGvkNV3Ca0NoSWXcprcG
m9LXA1aMQiTCqsddTOZ4FgFfsMrV8LP/dNIgzjAc/v5W+YQ4z147qdLE0NqGBk5r
A6VsE4oxfyyDSvAy5LdlHFfiKH7Sn4mejLpCNeGLqsuS2LBvy8vvyZU56Ik160EU
dVsZOmIT13aKjEg+gFXfXurk+hFtHlnlCy+h38/LWBk/d2qIB8Do01PAwPfmTa4l
u1W9SPEgecXATFQkRhqpRayR2WhhuQCd5rY7qqtsww9WoM796Elwqw0fQejWcI63
NmsW3fYzWcE0RgwMBbXa62SWNphiMt2SsSFsZdRmd7AH7mhicJzNRZy4rAbxSdPv
9lJxMvM29fsduVrXrcjC36DkEgCkUNbx3lL3K+kAkNwJe2YbUlNChDFn/n+GFWeW
v9YbV31JUqtD7j9IJjh8Z8UBGpA2jN9PEhIsgjV6adHSDqqMcpL3HKWh0v3P3gay
sYjAu4xj/cSPWYPb3y2+uI2GPCzfP3qvSZZ+47W5XrHHZaiYafX0EHlH4BC65YOE
0FJopBAfZSVFFBaLake0R1k/O5HTxNoC23F39aRSPbE4SG3azoKvN9Njy+qT/Gtv
QDOopjbm+Limm6fTnNmaTfwJBQF1WjimLOU9pJ9uvuYO0fGcC8faXrWId6uyszAz
+5cBd3hkh1rNWdfxC8JLhn73xcSn4GRTmKo6sDBQ/h0/Xtt/9aT3IslSjgwxayvO
s8pL+tgyEKip1pYmYhb7swzgKxzbSrQlP+RVbIOf2RNznT+xpMtgBFn7doUGHup7
5IkAiotKTwyhc9iA9ScqEBQXqWFniYNCKZq/5wX/7p0mP/wsxti4gL5HQEv1WRxc
CPbadYsTHAhqyZqDXDFaUoZArBUYzTWqJpytsEruphaSWktg/lYcIcJkybGoNsMq
OYb93Eg+Zs0md0UXUsGNrT12KCRhdLZqjA5NW8Aox4DN71TrgVizplt4rT3q+KeQ
6f3wHZw+JHjUtWAR27Id9/C+yGYEVY5hFw4eIN4NBGVwZxVxezhlHbjPYD8ZEFU8
JBX4yVXgMhJ/M5NPmhrhgwV4TLVYiEGXL9EqT/cwM3EF59o7WEJsBM8/pkMK+679
TLDAMzoCFDbOzxe5t+azqW7qprJBu4CF2Dk8i4ZZqsMfCewwHcEgqUMwdhYrpnyK
26WipuDvwz7A4Lvarx4RuotEKiTm+ZbJi4IwgMGEPDR86+MQuxFpHIf+F2+vkJb1
ZYrvWia6WiFN2EHtYPVXyvV6ZwbJXbisOkVGgtGYLbrnV7NejafuoagqMTrseTPh
F6YcnqcUtc9PmqlWyROF8pyy3p5pol11cm9SPKG6Glyn0GUeDKUHv5rV1nk227h4
d7u3nnpJdXy1SyHbui7O5tUxZmDIs56+vMPiONJHCs0UzpfuFjnJ10xLtrT3vn7t
RWh+Web0g7HBE7Q4K42xo860YsixiKHhAVFg5QfEn7+lK2cjSKQHJ+jT+XDSQ1Ez
oQEwv7x6N134v/kELDUwS2r4sLkyr7lGMa/Y1UtFRWZneEMSZCfe/SW5nVCAybkO
b5iVXBnR2ZsLhYtPtvhMXmoKjqBU8YeXIuwXsZRISbeUc3goMJy4IaH1Zbe4lyXc
ISXin1O8YZSs6s+EZOl1GzIlQUGaItsCetw6w4g2J7M5ESGwUqW/iBvZSuHdPQ2A
qVyUnfugGX9LBUA5gxxekh1J4VAckzFutJb/imS5gy4gqDif6ToL9pWNpNI/W/v6
NQsRih4lSZfZ7J9UZ6ZWBJxxr5/zZqVibceC5rVyVsTYg8rCGoaR+9gBfJUe2pQ+
7O/3ugTefV3SThjXNWlXZhh8+go1aUhCHiu5X34dv2aoskwPBZ15YbyQ/v3tHbvn
L4voP23TbvwQNvqZ8zhuxPht2F0U0ljMe0TOwdQ9A8/Jz/Jko9n8ZAKbqD7KBjj1
eks1wo7WYafFkeqKvOkALhNItS9TMz2VTdvqjGOBxlxgLzjaD3/J6WjRnAYEK0yd
3eF1mAJvDlU6PbHzkEwoS9IgiiVFK6RkFc/S/dKluTtukOpf2jSxCr+M/HGilY8p
+hnyNHqVfFozfUAgqzArPRXziabQjHtT6R7DC+7HndJBNEyGvXGCXeBh1zscWLxb
nxfo07Cx4rHWA/RGHs1/I9Pl8K/RoIIPi8KGNZgTaNy53hjaPMajunhFJS9QKIIf
YMa89m8B5eBEmOufOd65/ZOkGkuwSU3n5ynQM/J0Pi7+07E9t3fuzITj9E9I13X8
nopMmIesxBcwitKGFnOt2KV2gdyw/Yl6q6F4b+4evMAXIkuKISAEofAAGAktPe0X
uUbjKD06iG2NSuFQWFDx5Wc7TnS0YGTqXCoE+713m4sgiF+GzT21x0zsZWwJ1ZTg
LpW/XPkLVcgzr5H4JBP8IFkcmezB5BBS48MBiv6qKhXFo/awHzfykUUnIpO7AXmC
iQWbspN/zjfrenGSeFLS978b3ZG8ysgCUCMw103A/5s5mdYjO5CSLgKmLxzuTwxG
K3VXFYa+Rz9dAXxN1SWxs5MYl8nAhm331DNHJLikE6ewtSVuz+8y9beDgVFZjCnC
R2XI/56NZpyWIBI67fhtOs7EupAJIULxmEQi+RGsple6cP9nZvHrYJmsy97tOkyV
3RUnlYruv8kbwm9YPPQgXUazwc+29wF0qHy4j++dKILKo8RbOCDXJHhS9cY3PTMg
uNWgrNsjQXgzKOg6WMjFbAf5gYE+wccGXsF3FqqaY4CSK1oQMGhVIIpuDDiPReIV
Kr7zt9vBEOuufFw/CLfWI63HN3ezn7kS5Ya8lQJruBY6UL76LlpkhP7+WsJnVq+j
gdW3eO8h5F1LNKKdCxMiYcrPapWFHzjvb0tQ1PPDK3UE01NBqD40nADiTCf5O/s5
cceHqs8CmLWDejJb1XepATUMi6mQGytPbDSWv8q403lMprMfNrLuraiUaQgIrSMw
m6a9MkVjpQQWKqMS0KXV0k0ChWsLwMDynQXBk9dQ7zpi7eOAY272YcUNs8BFEI7k
FgExQ0Estv1r42nRrzx8V7nsGVsnrUWcMozAFjuiR9nUhkRfgd8fsj4ggvNSzOzf
BlBOtFBrrNYHZLMOW2XYzw70RJH2VWKvmf482L1gJmy1rCMuXus6K0ybdzPuupJ2
VXerTVSEYeeMz2D1EPtQozHoN/ase3CPlz1CMAoeSozoJbniAuiNyEGUmxXrgF7U
6+1noJd+GPU6QWmF8mOLH43mQR/YLN4nDwjwuHtnrYHLrYAb0l/ucLbxxQCJW06T
+C45qqXrr28MOe7R9AZJeZfT0Zi+HOsCgZzYl9JctcIK5hwpwxa0HhIq8FdG3KB9
1ATF308hETTvELv/3sDjiGwQ6K75JgWhW6Sw2CbqEgfzbAKmudxUnNKmuWTfG7si
JCPrx3VJJsJ8N+n8inG9VBnqqbkeL5SgcrrXvQAl8SIarV+RCBvzhGOzTm4DnXGe
NqBr4PA2VE0j0CD+fMgDyrl6b3r0GPA26YH1BRQl+XT6w8PXOUgEbtj1cLF+XG1Q
7XMbIDzyy+cSU2SJ5B7CYFVOZJwOMs+CNvhZGfGiN10Pt4+dtzaYNefSXomr4qPH
KOGVgPFaa3MVQhBNp9Pxj1xLhAFw6lCLeslmIMWO3ZGCj6V9X1u6xCYVhcw/YX4d
T2AcRPDyOlA0Xujs9a2XVHtbJeZ3C0vMXPlfqdYKZpHL5mzSdq5dbVXsxbcvV0IY
dq8n/af3681Lk6xF0XIsdPNi4FcBbnwiOvteSLCsfpXzslmjI5cgiYy6lOynRwVa
2wlKBZ2pXSHZxr2Hqse/suD2hFWRJXVEb/Ei6ACmXqpQGziegXh9oaI8Vioswpm6
as3X4q7gishm8jS8JaTIts/VRdlmzX0PKEo1pTJgnzjTxUxEGMpCa1q6cZxjCrnG
hOIfzOntZBQfzrh3e+4jxzhda8om/4IclVkkOMqo+fx581/XBelN0BFPTCodItN/
K1mjw8Dr95CmPxKkE6jVswQp+I61CRNs3XElGLtzEiGBdaNKYhv9n4pz+NRBVaF/
YoasmpEhlNSgq51wZ9wk8HufHJe0hihTqVnOyoSMbuAw1HFISPXYO3VE11VeGRuC
HXDlIVILYESOqHiI8nE/rtuDJtuVnygQvwtLajaNSSzoIdlDNctD9dVlsZkDC3rv
+rz/6dA+IflEJ5wfAUBZs0AkRs+ZyXpJKp6gGTGI9k/VfWxgWsJS1wmfJfp/+SRu
DBapH8DVcaZFKqSJBIp+KzHNhGAR2jEi0Zfd/xAfi7fNwqTupSVnGNGM1r4p4NpC
/SgzV9JQMj53ldpUNUdKn3PTHbwvxIJ+x22g8rkkm06XbrgEwb3sn80B8uDDm1mD
NRi2CWcqMFDuLRQxo5LJliyn6bVMGN90scJgmbG1xbF/wGA6V2mKhCanCp4fcxrU
ipZwbLsisl7Pf3ThZ2nfpQ0uwl8o3c4bgEQMozdORtFJsCXUrpJ8IYBYtaod1yXb
QNdqkoksStmwpHLFkSIh8Q7N07PznGl1qQclKU0cH4YyC3n1W4yY4QAUhWETcMA6
ByZQH5IKX//Xk4Xe2hzKpd1/Nj82pXV4+sNP7UQNP8Y7o73UnTwSaHVXy2miqZxZ
Nv166Mq6qau9nIQo/u0HTY6ppwQAgumjlngM0/5/odtN11wzUZiZPhlstrY1vbjH
cofvpINASWRqYNE2puoucGhyMTcGdZUR72wXm0EQGx+A+Uml4fC/+5nqRPjNNnMf
DUkFL+8+C7b82m3zsNTLUvHOc2kq9F81mZypv5s3FRlDxSNUMTZ3kSGa02hlptED
/pG/nCcMOkNmyqZqRl+myucom/qBtMESFX9D3xXfYaJY2mlRM6vIs1E4s3aRZLog
O6Y04PSUCPI+UTR0c6tCi8loZTSONQLVDy4dMeGLWnYuH8GXvHcw/MadmTiA22JN
U9H9LCodpRDiD4I9Kih/9DOYzwBg4NFWvMrmJG69cfMo7dfnCnbpH11ImlDktmyR
vxwqNVool5ApbYwqG26f3tkCUH4M/0Rk4xidTvof5Os+4c7ZcbQ/4PmvokE2rwg5
ZyiX5TDa7FhHnpsYwlz4JxH3pEOkxl8DeWcmThUUVLFaLHv0qeys8ANBXQrvK+Cw
Cjbh/xiiP288pMVSeV+fchTiPtgMmcoGB6IHVhDBKf0vhIZMyoj1tcZrrL+r5lS9
iOLppVlk8G0DIjeGETfKBoPdIwDsBWMO+6+EOBh1OUPgKKSoOUva65el1SytVGJX
jsRdL4gXSqFZQlu9IbhfXOev0GjDxETI4/XLENy6dII8oq6cctEYPCOOWUCU4/V/
0JL/A2xQ+4cD9ckedKHmQqM908Gkrq0fNceUqDy5uHVwFyZim36J6Zn/KonUx5Go
C7YrLe7gU6/H+TNMA2gl1fRkhK+Q90NOg8fkby/KoOilQ2sUeUp73p6ilkoCjuXT
CUggTBPNdUCmXE+lRUsGUUtMGkZgPRWwexU2w0iZChX0DWcn2g6k03yRiwJmSLvH
RuzeTArjB/eDv8JDPMy6Pt2LGS5RSMSj+5X/JkflxyM3xZ6UogEgvXl46gd6X1+q
Rflhh9VgiMjyIl8kPm8FFXo74BYbSvVHjcYmJlXBXk/W0WlnZB8nSxApsEoREjBE
kvPq7awyWWwl22dMWKf8AL0gltT/nBwYjBCYDr4jTiohWGwYlQ7trhBA3CI+2TZ+
MxGGi2kOmd74XWQO8NHxRLSMEPS0Z5LmxYEmjIs1T09+ax3S/ORDgVDQBTVJFJXH
EW7nSAMtI+y4uanuEif919fndZdBnXrgCqz6RYAQPieiTkroaSwEuhWQ2dHa9vxO
i9lwETKZsJSQ1T5iB/2+c2+hVvxLXec8fkDNqXrl+kcpKLZJ/TfRnvcZr16gJpcS
gxLZPOUZT9aNPSCBfQqtOPDwWiMojWBx8PxRsRGhG/UBNlSAtDhkeV5jj5aA3nk5
cR/A1Qh0N3bX3lTGzSpAPIeZdlx2Fr9/dmlvfwnjjgHmm363GB5kBwxQY6z7unUM
6+wqmJe2ge+E3VDukvVWPm/uWSTb+Rn8krJqeyRVETM6adytkG4iUK9IeppAmWV5
KHveVNycAyZX7nxZFn8dufsoRQI18TQjfYRMcAMFqj0fWbWsFLZqTTi8jR96jk+f
/xmhWuvvDTMvSlhZkMWOqUocoBNNHhba2meCBlMTNlyO8PQ9FSUzy+pO5/35h6u2
ftdDcq5/EYZfr3EcWFkJ3dQKCkXejaGklB0Wm7E5S3zizUvoSEV3nwNlU4EicmqV
ra410p4OqwTqLRZcPrly1gj/yy6RediPvErE4jUhpCPXeOLPBFvkHBtEWcpKhDSG
0gE2wQ9Hw/JEOOJh3vWk0CeHLv2s5gAEYefzfF9mNhfk+XYVcz8q6JJlbA1x+zD/
U3ajDHWf+nkwNzmGPOK1O/G3eTmXJH9BYbem5Eg1FDiWYvSUDu9nQDURROYAZ+eV
0llN0gBIVK9JJ/PpBZrvFXiUz0vZrQQJXhjEfR/MxGMIbxGeVpOxyGypxGvZ6+O6
qX3tmV4JUVpgvJRDkx93C8A9EGrjJ4K/h7zBf4sDIrhy4wSqqyz+lPyFG6fQMOji
veB/c3gBZkgOdQI4Jg0L8O/trTXpEIPEmbV8UchrQSPwxwCWKLxRHKq/iHFvo3dR
GGTTRxL7zKPH1CW63J4TnWDFJjtyIrnpJs3WR93HfeAIUJ/fs5s0vK6ok6Oka+eS
g34fnEgtIFyd2dMcMFSyaS7HRKUqiutTZT9Li2wxtFCHcnZ5qxStd2CeeGPYouQr
zRLD61evBm4ZJNvkVc/0vW9oBcmYpfguC5EtkhtwEZJv0jeV4/Wh6InWUtcfTZtC
82iiwB/KALiMM7DCdQ9VVLB6B11iqqvEnYmWxAWR67U8hxA2gJLa5Xz67hxTpuvm
mT7rTM0abMobqVxkL5PdHivOuGxZBsH8Yb+Ky0Hyldwrap/YBFtrR6IQLqNDDlp0
Xl/z6zr8mDUIr+6sVudkNmXm611jte2lmnKO8mUuWtFj+wQEmWnmXRiouHKLP2F2
Amv4S6TVcP6+y0v9flrIW4FU+uVIsg2kSLOE/mR+DYAtYpWInPgtklEE/buNtfSQ
s1t84Kq7ZSvRS9JRXWlobG73rl1Te/8C3M3CKitMO/CevC1WQBatD5cxJZo9KmyQ
sQlRX/b/7pDaieEgi/Gpm6A23QVz8EpzGcOlyiUxUzP4ivU8UtHz8ptGbH/cz+xn
CL7S+i7FvYytNI//+RkJiD/hpqAkeHaedx7K8Ag78CS/bpPlF5MAxjOZIQR0rQ9F
pgXFnV0hreHJCPjfG2F2FeTqagzMiOeAYzO9S3kkvWoPqzAtMRv9YdG/eEJsdXvX
1dWvfgOcf41Zv6HOkxCA5l2EX1gANLjWUmW0p5F1+UNX5k5TTUq3dqDsT51nnaXK
ISXrc5YpvSHbWsJi7qKV2PqFMY+aLggn0yR2znljb8EvYNnp1rgwyJ8ypwNKDPm/
LngQmEpQ8pjQv13Ha1zUBzp+UFrKEpF/rj/GUCqjrll6zq1UG/5JpCabHrQ6Ul7r
ASvSF7JB8CyBouh5EC0PEviqX4a7A6vbXEHHhKkZvXbiroL+ij8aPDaxO1BSNziH
y/6VMOOvIZ7j8/K6nvX6qj6bABfBFYn5fMJWvl4xr/YbhGLV/Ec5LOphETTlT4Ak
4RQTRccwzVBmU6BTmKNdPTtv5FfMzJNWQNET3Hnq3Ku0idx990C+2V+/tKwKfs8j
nkVAiJy+8RNswKb7Y3eXUPcyq8tEj4poPtVF3Xm/m8GzYyaKVjrkfQ1bP7TzF+TB
7TbG6z9wWiM6HMIcHLd2nBmofo4bRQiToBmCA8urFCrfppTqCFg2n1cmhRZKuxDm
c1VH4P1Y1G3wXpEDH81KOCvnwTsDQ3MShyA9EREG46mC9bh1B3ugBvTbgdqQshaJ
1MK/OOlQXMGGlHs1o1uQeV/DU4oleUOuWtB0qu2V6mWXvU3SuFxRcCX3+c9U8J7m
rYusoZkEuCT60U7A1t0LqUgj2P0x8bvl7owAaZw0MvwAlws61qbaKYd9uC0QHRsK
sHcy2i82SgYB4nquEa8/sREEJwI7qEIki6em/X9pQxhzekOUSC+2cNl1GOy7qx5H
u5CkyYkctuGO8FOYcRWQT1yqTtQSPi7MIX6n1ms0nlBw82y3lWINqdZqk2r73mCC
xRzIfTEFlwpXZbzwWam7lg8rz127/fl+ZJ1TkNTJhG+kfGiq1+DE16ErJY3I2c0v
8J9Q9tD+KHOw7+ngMlHzFJAskZzexiO9b1RVvZZcFQ3bdXUHsD4rw7JQDM1Mv27M
OtWl2ftH1NcdbJBjoCbzHzWPUycAZDx7qmBv7O/9vr0HZ5sIgaMv2xVgZE0f7euD
DNofDNUVbT7qdCrtQ3tO66rEppdmqp0gALeUtKslNAs188OBVovEsriVubiBe16r
gc4w60OCLBfnaHXx3gWAXPjtVbFQucbktguYwrRABLZXZiNq4l29cUOyE2idnn4H
sg3ALrvVG6jXCxd3n65k+gOzJCs152H2BGdTEuDHqBQTkR202lLu0zxGArLqZVUt
zmlZe1ZsS279BU4zjz4Nh+uXzFUzXQWrMJ0okPsQx4xSE2s5qOjy4MaFmiYZy+FT
GffeIj5rnicc4rCO4OABTBZzIrHR1qbglYwiFVAvE9OV5bS4r6s0sZcuGM2QGogL
uZuOGuHSa86zrFcK0Bqj909ru3pgHTtD3yO7P1w8i/OQUac1UVndgTrL1aQAtZMl
iItWATXZB9141Gwa2E+6aeU6P/AgNngXJCgpeaVCuudOrhC3htr56cxzI3d43iVc
pyDXQ+hmZ73iZ78kOFdT0QwYsRjY/FrRbMuC2sNDERklJCZTRQEBf2ddUPIOEFzW
DlH/W5h4CmYyX69DmdkDD4pJgTwJomhsSmH/eVUfkZLApvtZdiSk25Koko9Sqont
E8MZxP3T+1nx8s/7OmBYDzls1lNj1GiQYjpGx4dvmqA6NYQ70hFEtlFXOIpq0snK
UgBahRca5DRWFDiXLNxP+Xzs2mnSFtfhvXuNMmTVt7TdcUby/KY41DmCYRJgrj9N
1rBIKsNEVCnKSh65wijvVsv8Q6nOTjToOk+CA9eRu6TK5ISz5Tz2sQV1Drq1vrWf
XLtOnbmXWaqFPUCUSXW9KKm5+5VqUJ9q3nB534R4Uy/iXSlaJc5ACIuSvx/VxQsP
UyPkKlq8HLDpUUID/cyOpfn3Mg+AGAp6bXDf8OmOtDcCLXJsu+03ZG79pJnvTpNT
Uk0gFDuo+UjUkMLd99p0AYtJmP8gKV6DZxuHXQKqjEN/QZryL1BRqCCmIRBJEGtb
/POs0GxvqWBX4W50y1IWUBDjMZlU5ICmvtc5kBRZqT/K7CMdO9MDpAYrtbIFQh0D
a++6koYZPp7ulRALGdhuClKOrCgHfegoyJ6MuUmyW2rD5AJ40T41Ym+GR/mRzDRy
p19/XKy6oEeKLXzSmUb07hzIgVYDC/hCaDTgN8bdJK25PprwJskVS1NgxTTIeuU4
CrQBcMnz9jEaDVXRCpOhLFKXWAD5i6NmimrsuIeOBG5NnavQglPEbKyL5oUq+IJ8
EB4R/XDoFYPecpSpNDacViLzTe2uH30NodFHP6zqbSHZu0CV2gz2XRXPiIgoHr7S
z2AqTAIsm+5sg8WqmawEQfEyX39UR9ioKpynq+1yXpxZ9mnW/jbLc6wPZEPZfHf1
tMnW1jX8OqbuU5dQgYbk7k7vMV5oh4OoPLv1kB498//ZoeyU07lW1OxqsZSoAf7C
Qm5yi5y2ntYkOtJ9bnL8oASTJv8/ytFhCTG+NMpsSaxpaifFCDcOHM50bO1ROer7
byrl8HtvGG7LBWrOw7AgeBG8Mi4cGPO7PBkHr7OlvrBsNeajMD2+eAQ/730xaWV2
GRZqYFoDx65uFEy5E+4RrZaVKmC9G8Yxwm+x7SMmCVMjCUwEjwWGwfB/p3p1hrDn
kZ75wQJJXE5+gIFbLF05+8YEN/yS9wCvdQYpN9n+6LjSpNq3SywVhhGPb+h7PzV5
MtLYeqv4isS3o2MCVo5Rb4cWBSRkOxII39XK0a0OFv7lZsF8uOMJX0ColOtnZhS3
`protect end_protected
