-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
2n0ghNR3cK9Lb9C+G/m1AhnjRa0fhT/9dKh2eXTqO04+BOzUCosbGfQAAJSCt/AF
2jpZanbAdjVvprs8Bx1Zo73BJuY8dfTPTqCc2P9UzEniJMDL0s578Y1sjGsJBJDN
lYseUnYHXj4CoYdXj1J4TXoxuy+Y7NIBMRnn+Sh/J7dKrC3M9Vn9qQ==
--pragma protect end_key_block
--pragma protect digest_block
lY75ProVtPkdh3Sp9VVi2atJzqM=
--pragma protect end_digest_block
--pragma protect data_block
yOH9s3FDR957PycH2SJKS6jtjjDT7FtCTf/dNDx3HnJhK1oz0KMEsFkS1YuEtJ+U
a0H9ZCgtsIyW1GQ/FuZ+CCz2Lqi2K/InvRDq5Lj+iBBeR/+DHIZJ21OS11Ip3LFY
eVyvjmASGMhNrJc+0U2D2pIe03BWis93yBaFFBbYSZ0K+pBuJ7e1JJQYO8VF/aWb
s+9Ab4wRO2XUG8HnOcqwFItrQasADIaDGEgDOIZiRYhFm505lsr4qtAMoaP7Xy2o
JlPPB/x03IJhUeTPKF4vvwynQ6Sv8no9kuglu6I1S5nvP0IZm63dteB3kyWF+tL5
CdzEH+/udrEjtMjz+KinjhCUnF5vHPRd/dSUimEqClvCeETwCj8JBHtpRno3mCOM
/nLZnAzrgflrJL71xA56tEaRsY33laqviQFSzweM5Vunc5IasxYXyxpdxMFn4vJO
B/E3BP1SSxO1/BynoMcZBI8/Oo/B/1MLSzfxOAe2PdKGfN+4FaOJtfPMSXsKFWJ/
aV1Vrfz5E2gdC18My6I2Mo7Y0maZWYVuA+aiZOCauIJecwRXkgj6FJHI10Qa7IhN
h6zfrvjIKMZXAnJ+3LrOFtTbXrp+40Y0/zJd+HBFuBCtDQjcPh5AxoMmBgvyBXGL
4w2XBCnZt0Ss6hNuZZASUckIH7a9ZICX1Z5DhEsJsjM9Fb/WQpEj4qJfuSzEVpUg
6ShZ9qErfSO3ubAsKuOpe51QtMtExZb1kaTJOqGrB0P5IXsk7Els0iawt6/s+jRk
HvP4GzMtZHkOXG/En0jZRA3/4+DrJ9s+WmuJg5zWR18ioK8Q0ePFnLPGBiieqml0
UIpyLoB7AOLgs31gf6W2zXsDyqkXDim2QV1lgi3smSZqI4i2Ir/RXVdYJeDp7AZj
4hqDArjd6mgmx4x3dgxW/IM/hQLdAu0Wd84OipSLSr0S9v7iILDpPZKQd1FpC9Pm
rkkVIV3gUnI3scD9aZn33AOnt4E7Vcaxf9lI8LOIvZLPqxRunif53StJ0IUIZkSr
bEuIhpT6yBbIe/avhAUTJazmVsNosHEIyVWfHmq4hfn21MvogA2DJBqbvGXSwF6U
7g6+lsCSWDgHx5TpA8/M3vo5/OoQVK8L0OAkyns80bs6+SMKT72QXj2Z2Q3m3O5y
92ut1uIAONz6SNCXjLO0D5yhaPPkjYhOs4+9QLa9SgN/chvfgXGDoBQTJmuHtgeS
0RR6h9V0pUcC4iOf9eiH7pVZRxYgOJIWrAOUGLR823Y3JvtJpHa1MLVFFe7QR9O8
RNyciJ1NgRNVhKkom9AxWNzWZ8iMvnZVctLETGkLBFAxnbqnxb4ouNxpS0JfdH8X
jJqiiz2sAUdnwQ9XKNVf6DfL4bkZsjJR4JLb8bwq2EmXJOJz+4GpFq26lXpX+h4D
HhtRJ67okQCyhU/uvfVeYasUCdkhzA+h5RtYKW6E3NYoMUw/AoMaiGFJXyfmFc7A
yCchgD7+OB7vKeZkb7Ma15ZChQXUyBIGIw8TZhm/VCCR8V4VGr7nBMgWpy/0FiIy
8vZCfobaO9eCkZBK9Hks56mc7c0YKW6WdK9+vy2CRs9HKKfPnCIofaaOCFBV+0WQ
Mk1ok2OLlW2AqW091L0ppr/WbeQEIkoNVxeeWU98qO1I5BufIIe2LHv+T6LibqxY
ll6tITUshDJTgR+Lco4RG74HN0aySWW6wITOuGl0aFa/rn047THWmKTURTHEutcl
u6btYIK6Knbk8zFMQcqAyHL97uql2B9lwQmgUmMcyJOehlcR/MBpKMRc17zE77J5
myAnOWh4wvw3KUjx0FjDMERc+dBBc/4iqWTGV1vpvfA8Aglz7HLyBP7aofvkGG1X
rSynaKqV+QZg0jAkos4xv6UrKvFCZbON3MJHBASYC8AQaVhSXHKNqSrqvzV91VkB
org2e8v5Iyc+0ZKqAfCqYsUJqra6AS4qFCevLv2tUEbeikE4O7uqo/hZmnY7FB55
HSpVmuXRhOxVFMKN48OV/JoTGzfgXf0VN4o5jLsfCdbxHzSiWrNmTjxzIRmkyxr3
PooCnTyGzZutye85vI6TYTX/K3pk7jo5XoWOwxsEsnc2RCnM1N+lJ/yyQFeT0uVv
3Z7q4pFbocLxYOqs9zgQJ4yA/Po09Nl25OyyDkLp1SiQ7aJhpNMg7MohcxLXF49a
aH61xyodAR7krVFByAlkFZ8GyYsnOQ5Dn1NJejqtX34+6qpOtvOv/rYdmaK8Vy82
tHixn2I5QdwjectLCcg0odFQEiYgTmbls94y1OaWFcHPFHNFM8CC+qLskvHkFOy4
fxIp/0xHmfU6RhP2clyH9DwuDcQgxISUwdivYKKDFUrCxR7oLSPRjN5w2uZgngRT
3ijyJuHWsNoXYI0QpMdraa0GoXtFmj1DsLBrXBXtQshaFcr2RuKwD6+umk0XXROK
PNEBSjzj/froM6ht4VLaMCtPV09aoAOIa+9QLOXxCrqM8ETwYKJrjg+p/2XKVZpq
UoLgVgEZMYy4OOHNCzm/KM05fCwO2dz1FTwSYOjTVwlI2XY533x3SZjWEKxjxOzp
Tcxmmv2Gxi4j4/bJCfvDVRi9LgeDj5zMiZ9IFuXlr9AU6O+Ppl4W8psiWZtvakuf
57hozTTK5aSNqrBg8xeUMkOZ0x42X/73DioQwF/Ubf2PYTSuANPiQsG+Gf7ivTXZ
D2duzI3untB/IpQ8jdA0eDzk7HVBrkjgAoUPIm+xFmGacumLrB2ZN3CVpJGcChXU
Os5iSUgiATG/Dqye4CDP8Ke9uzc3LFGbcMfrloBzyqhOiu2RLVLkWwGpSjx/Hlrz
tM0kAjx2sWoSuZifVMXXncPVdEasMJCkGPeOQ8Q4AGHiTwAZtzSkXm7IVdy5rkXg
gZj517JdZdtjLTovwOO/Td7MpNsa4GOxG8Pl7iE9AJeeAbjY5ljBHWxxX+YSrhtM
2COV0rC7NP66ef7oqYVar0HH3KUECTdWpwCyotq9MQfQ1D1MJI7KLc6fBUbyuwVW
Y6kN3j3Cc1c7kFJ9/R/X1SHpF+chcvMchDhQSnWHVXSySIDkqbwc+xAL2URMIFfz
iP67JMMHRAWcXScCjQMXHgD+HlpN0hJcLw8sBY7Db2P5MKCjZjNh1nX/62BLnkIu
Fpu07HVUEnGSYpIFd/5rc9jb8/1wuh27rNJ2DX0TbLXs6KU0ug1af7PttO5AolHC
xUe4xk7ztvYTjs7fCLFgO1qJA13btdDIR+nL40KxagE3n8SPy4Fl/yspS0U4VI0o
lgZfHdPtO+vC89h+JW1dTD1yuLJQn2f2SruW6f4OO4jhTZqkjfwM7TNnCXILlbxX
VmLyT7dgHzwUaGONuSj+DMfxHWmepF3Bq0xbGu8kVh2xbfVEglb/x2qlRt7Mdr2U
v+Rpey3qwXcLPn42Az+0p920uborhes08NvBXmEwDB5CJIDB2ryMwS8JGZZfvija
BmWPMZ26u1OvrV7wZQPTpGA8m6xQntRfYohiPDYYk7Afmx+LXoSMU6I0Mga7KACz
+gkNV5vPnhJgep8uXeb4tz6QoJW0Y05G4TINm6HmC/OBCOzLaGGEHB1+T0Q1Sds4
9u+fXCqYq1qtgvqvH0HPXaR+LcRzh8W8pb1enqR4zOTvYx9KhiwU22nblZfCKp9w
5akcKMWIIncBP4lsVL6Wlip0cRmQ+T0OfUrq4udGH4vF8vEv9pIIoYyl2MZvAMyE
gL5g+oXiKTUT3aFmcRopU1ioga9ECV8dJ+E3fuPvPta/PV+j6QUuDDFGaMTYBL0U
j9QaQqhMvg6M6YEJFVeFsyrrf/meJQk2B76IWJdjLwWIRh++92CGh/AakcOxoGF2
Y3ty8KhQBb9to+jC6E8sKJ0atVlnxZJJsImPVB8h9TeYsS/YmRvUF8g9DGE8oXX+
IlytsVoVHsvPu8o0wJctN7e0r1wJBbOG4OmE5Hy0osmMJ6iDNIn6JEULW6bGdMYT
eqR8hOAxdfAax1bNVEfHUUNuCcE23XuCINw+SPH2ff2zCKC1awFATkewEu0rNdZt
gGgheC3VP9u3U+MOizuFhoG7krHvjVzaMsX/SUmOZ08uJUkzQLJD7g1N0zcCyMfo
iALKC8vvZrPVxraBjGT5GLTLnYe1n0woOe28ifrEl7M8QshIle6Bn9fAQ8h7xo5N
I/mP7ygQb5NH31Xwr0kJQWZ+Kwjsm8E5APc61zhqZYgF99PyiJXmFPznsU/6S0f8
Hu3d1voarPmtfp/BKy8pPxTxGOrJUbSr91c0ihqQMoStFKq3jmWEe6x34TMkFT6C
6NZPuS6Few0gNJpScFQxpy6NXKCjRSyQyR+r9KME8TfsycM5KfNYYzHf+eBrb1D8
TdTc9Rxv6vcRQdyUgXAG2NSOa2FuLwLMhepoye00rRTQ2K3f4HZIqd/AzAWn82Mw
J1qcV0NDe5mCm5mzA84U3DaBM0lKTIXgMRwuwwniJr0XFwPyX5PfFgLVB5/eKbBd
qBkY3QI6q5kDQhOHDh2J8DnjWbZJIyy4ANTAC5bP4AwYmTGNbZa9IgyZCYT/nsJf
EU47kaxrhW8DCaZASYKMfAC4vmif7nGJvNEXG78o8GXuV/ax2CbOPq4RX0cBELYs
fR7+BJyDdqkhg0etufpeLgqKBODVrC5Ye+QUWyyJAEomp4I0p5igR1Hmz0DXbClw
RJN9/YHeC97rYiMcvYLdPVXiaSsp8WUJVQkSDHcIoQQSkz1Zb2ufNQ8O3hY+si4v
iqXfokUak5yQ9AoJZrtaI0oaEQTW4VzV4Wm0430G3rpg+334jVfYXqKayqZDXDCm
b6HL9hk9GHz+envozxwCxxq/tF9tcWUcDgxbVbmqSmmpZmlzpZsiE4dHkq1cQEJw
v4fJ79xGqeTWyA3CCNG4He4V3+Kfuw9jrYNTu3YpTzkaNdPHz7Yrk8G4f8LD6oNm
P9M1uKlq5MzXq772LmNKqolenf3Izjt8YJAQ5qaYMiWtroIuF12pii20QmNySTdu
6a5lPpiOjpuNYwlKYkRQ03bUhYZUmtZnHbsTmBQ7cBxu2C/1a8QO8WJFIQ7J9kkx
B5bXcZDwceKG187pzwkHnLnQve3fi8PvEfqjXAYKwADDMd5LpbywXWpi/aNdHN04
YFsIfatdFF74nnjOkEN5yxp84JZwXsjYf0+3Iz77H9YkEQM3wh4UrKWj+Dk64ZiA
Y+C3NBX1wF+/AGwEoVkvI0XwD4feJ7iw83OS3mo9qMaVCBPdA4g4acNcA+jaK3zh
f3UACOKX6h5i4HbQ70O9vIEvTqEN2juxH7pmprpRxYXMai6JKXJMPDunAFIVW3i5
vHg1m555W72rq8i5LL9ehXMk4KH/r6P4g761OXcrN3obcDW92Ivr3Ft1hbFuXYUh
BO6cAcsGgACTq3N0s78wI36BsyIq25LyFvs5l3Siff19T+DCyBiNGESOufy81hNr
QJrbTgA+OPD7+xPx5wkkdQXK3ttmWUGgSW0Xlg36DI1teZ0wTFkClqvlJFQTzDSB
K3zY+cnpeIpBr9vQJ4YEWhonJIyyRrEHRnd+AtGpUHtF/27LNz3ty44cBadgSrE3
ziUMp6QwXrVMYQZF/YT0LHs8ulAuypeGRpmI4ufDrA5e13hTm0spZIUCyi/BoPNg
4U9dyZst3LVLl+PXi12TppvyJRWmnaOnlxTxyogXe+uv5u85rBXlxJns/CnrplWb
+HtEAyh4lykcR5IQNeezL0Td8xsUlmTvXBCS3mroWMV3qN4l7EkVqRfKOIUzt4fc
PkBqm+HhhqKkCutYqGMxYfBxVRqpXhGJfWZfnwxAb7783kqFiW9ZJbHuZyh2M2/f
MxewxkKdpq/52OSQ71PUQDAmdG/JGpD2GT4AZQah2CSJt0uGkdI2OUh98nJu/HDL
XSlo+kj09EpYnG/HC+h8Z/cOr+nH3SuSbQ7FtJJwF4zFTnvlFeOAiOwcVbUrNSvu
1ABdFHsx0M54mw7DvLLUNoAl9MrHgWpm64olSRvbhHB0RVl1xs6QPBg6LYRHWaah
a+db2aMBexoyryVnqzY2vrRP4tSi51RnJMdDI0WIQsZxhgPTXVeuMoxDeznJh/P/
vEqLVK8jvnQtdebDiZ9Pn+IwyKZIC4eUzIGtYY6vX+63IP7M0OZ1yDmIljfNbErM
GSvv4HVsfNTczOnN8B3+nU8p7jMix5C0mRgmtlyY/IKstnAlXjnDOCxH4RgffLEy
lsiECjwCNlQ8geh28uEKqmGOteoNf5/JpzGAFwqA+9sVkehd42ZQT17LV8/x+sOj
J7reYHJrROAwaO3/cPmou7bt9LSTygDg0ux9RmTKsa77zbrJdpVUNbj8fwOPugAM
uPy9LtfhCTrUKWrtYQUemUYYc9zKwGFZGWaRYxv+bSfdbG2kTZMV63FhvJLgK2Er
Lm/1jOHQvK9i7zPJbZYn9s0rjM7tHbmtx1pItkKu35Xd8Esy61cG3mXSF/a1onfl
XUH6CILIlYzJGUf60UzJPPz7aGI+9QA90j/mJZwzRCE/rK8U9BAB2j9pry0ED8Sl
S6KgwrFimIfvp7HZbqoVUCHWFuJchRnEZ3OhafQ7YHA4T4HOKd7PzPryDcixL9AS
NO1ilNgc2mxEc35LcsiQJZPZDg6kXZXpGVM/TDjmT00fEyD7v5slBMnSKjhebN/k
cWqZBsWhnE/m+GdUIlOt81oHptQmuVUD1OoGqaekwGpJnv9Czo6uizZGz2+Ca4wT
ICC8Qe3/zz/RG8fM5BtxMGFFCZJGTO1v5anR6NNSXd7ZyZgaaNW2odm2N1dQL4jB
DoXPxTBI898pwlRUBx0MvtkN2ampuCWfzeoO1uiqQsbXqtKlK5ADWNHkO5jB6LvW
F9ijiPnaS+G9mo09MTdYAG7EarVc0tzJjHGVMv/FaCpyWMi1nUv9crzbFqZEu5Jh
kZTN9bnS4jGANqWYPEWPMOAbDNrC1XjUhBHVhXqzNWhm/N+q1FRtSbZ2of5J3ldo
+4InzPf5DM6ISN/bYugPQvWbw9HX/CIuZdPNlVG0a5yJNAXxsHxvzKvOQPqWVc2h
kItSfZUVAMZzsyqB8dydd0pard4YJDqsK/DWrqfRxDDH1gxmxQyhatPktXFJ5P/Q
imWydo9Lhkl9C16EnvdKF304cYkpmSAl8ZExQcdUwyVJQrW5xKeyb5WOEquT+a3e
xtpOKVgTMP8aoymDK3NhcWaSoVoq+ih9CrjS09qvTxdYjt/S2PD97JWoy+ruqW5m
hXfsq3uO9z6XpriSNHKm7qJ401EIuRYBoFXmzmyf29YCvH+0E3NQ+vPUjfdKNqL3
wayYAARsS7PsU5SkO14QmnD17Haus7MoDnvHYr+2hjhTeSErTMh1cUdPfWaTWOtr
sibZ7ZhFeE1aBQCalxkb+4R9/166rFF0J+/Byd8w6chtoThZf9BL30+dcFZHaxyF
0vPBFnsNPIkuIN0kfVuKW8X0AlgjBPWDrZJ7JBOhR1w02/w4e9sQmPKDG59hv9Pt
MJD4Enm6oMkCpMDgs20dQzzGzhpEkr61VoLT5wcvF8wEFfLjRBu0jyt1ESmp6JrZ
2H4kzxQtDRoeQIEWiRen045F506mZasXv93ejBQlLoljcpaDbg+DB4CiUbf6aNDy
AGcRKze6AThqN77V4QN5sTZurcVwg5ptEdOfVN9DzyCd6NdI4uQgoDUEMp6cCRee
Q1kz9Mq0XzZFtsC2si+3D0np9FmVmxlA6f7nT6DFy8Fb9nJ3FnOSXDNNX8xAViH9
aqq3NHiQjXC/qU9jjBige0YLv4P8PYAjI2H808MYtkYj4w5ecrboPijwNvGYgQ3P
bJgEAYBi2mfc11Xlzn3/VEkwACtTLGhVMF0t1b8FlabyO942pAO9JktaE8IXuoyl
QV/zlCcSbRSPdYmnWawptT3fHtdlKA+t9vuSdovhGdqJxrjsfZWoemXukLmK1osl
kOBkARQmaCgnB949HIRVy0EIUwy6tq+dLOHzilbTBiSG4RQkEbztONzl1N4k7ZFq
YR4vbQOQCBZK4ghsdG7ydKo20va3V0OwlR2+wLjhhiQeh9Ha/2ry1hGR1zziMyGi
l+yH4+pNu+8UbwKuxc4NSRrG1gWTlkt+hvlaI489sDoz27jq0MnBKlO15z7HcLgh
zwYzoP6snNtE/rKVmz8PHjjAXB0HIVWZQ26L2P+rQbjC3c39uKdUmmzsqjZ4Iefh
fMlOKiPqpxU2338HrQwKDmIhjnEOaKyHraFhES0G7qWnBA+u0IXHpSPa2+M0+OSH
+2mlgl5cTvTJDu8+5nItsCRZbKRPQZNIYsUrvRSI7OF9hrQCI5l8wpUelBIMvFCW
6RkOlw8VXOPN8uNo94UCXZwFQOD45oe/9ScfiDTaQKEyDtbJrCo7pwnbohx7Uv7H
Ww+YYtuiAbNF4UPOGRPBwt3SmyX0AVDJULhAYpIz+J8TQNRBGLzck0+prcHTqX+P
pkfGxG9ITrAZMZ/xEBzknOmL27UKd//+fuhI9f2bQ431dH/fTu3hNCD3Kzbh3x75
OKfpG7Ta+Ja7R56nPWjhvVHYdR9IJ9W8SyOKPxqac42yDBsfspB4b9fVk+p9qjIo
KfHxG9VdQFPbrMqIHCsKAXSBlVGbtWHNyDF+tU8bD3mk1xwDvooPZzqVEn02hzGr
Ck7g6WgEVhUt3G4wxZTiBjiy9xkmDoT6z7jJAPyHD39YwD3l0FoZCal6/pKSHFAm
MjtPnhxjWDLNyQ73OEGEl5vPke2qxudS96c6Vo3xQKbk2x+nfovgUnPCZArtciVJ
V2IbXGz8F3XRwuhmDuaS7ngADaGM+R+X3EO8ZtTYnyThght/IjcJ7cbHXNPex/A/
r3VK+LpWCotYbQ3R8+T9N8RcB8jtD8Bh7wOpp2k/k+SG4iCVcNb0AcFmCqVaAJ42
SWpOPcn3IwU6YbkVYrA+ZfwrjuvTl5JrCTmRoJZMPvIjsBmRG+f3ExB9NLtqsBw2
E7clSTe7sAKUKoIeR3G8M1wNq8f0g+yleaGUVTssNFtB3YQ53q1Q1La0ich2yrX9
yniZQ/bNbFaBC+7ETB+GJL9b3YGSDwP5+JRuYrgiF/iHl1hZcG9Fzv4CkZsqgDcD
MrHj61TGk5BT+tFtVXKXPHOKEOCd9DB125shXvEfELM0mskp3hRc1dnbjBP3lKJQ
w/4G5RkasIg4NU3oPZ8an9QXyMa+Rmm7QKyQfzvLCpdR3T0b4hHqbQdP7t51zNTx
4kHkTGan08rTSgu62iTagT5jbxr17Wpf8MoV3hz9WwbVsF+LTy/OsvohtHyBea43
UnjKtU34pHqsoFLxsI9mhps8qhm5yPVmjRYnkDAAfyJoHNFx3DWzaLMf/tjC/o1O
OU4zeLX+cpqKnYFVf9La0t7EGCkfkhZ9cOhD+AmbK9rKOhEmVETpReJV6E9VO1G+
gFbCg/ZwNvDBPknSm4rdfOT6U9L2IgrYEXvD1m1FFlxmRu592kDW4g/dT4L8EHUw
xpuKOHpHiCafKAaip3Fs2FTGj1SLiJxdxtnpBrxiOFrMAw1goe34hQ+chSXWH5wU
LwMb1lPkw/RWFlLHtt3SoiOnvrKDOlAf8kkWUHzNVFhPY2d8ZjxiRBALBFD4phl/
ubccXOknSaOQ2m32FUtmOqVzVPG9EEOEIyfHsyXSjNCGI+YrwIAnPXKx8EiaejUV
U0ki0zUQLzo49ArDGc9kjmO9h4A7/0SpwGeZbKMR4SANohPbfh76L5/0V4T+zMSE
+wYoLpDuGJngCaJSo0uDXSlEb/TFfsWMHMb05NM91xmuCQJdRcdMEviQ20fcPaWw
pBjpqkNDrEsyao3seg1Jw1RWe2E+z4GoPwMMkroi2Zf0NeTtYNJzu1pvIkrSMozJ
EJm0fKp/XlMwSffWmrBz96liUnVTj5KSni6dvl0jcXGRUadTybWQumX4Uez3NH63
fz/ol5FeJEXrNbkMw+cAOtiakXjRKe9Z6deD5g+ftTCsLUhxA/1VtjnSvO7i8ctc
k4e6X2UbiwMTo3pd1p3zLZaPoHoHgq1J5xBtr09MbO3Abo4DxvpwLpxlkXGb/+OA
7D+oq9m1pSW6vA/HrKEVe/WEAKyn/R5tP/XXTdjBU5XixSIcDrzSevmMlAMDB6LB
ZievsknPSU+qWDos/r39XVDWB0S5vGU6HK/Z7gIVcFTwkL17E8W+nsPhq49ZFdLc
1wG7G7MGiEpQnTlYefLEHqFXkYV7zqb8I5qwGB3tmo3vQxJoCtstE4SFFALNOCWY
uZt1myw4Yig3BePi7bjYQx2UZNQPIELSOhSRXiVz3qMtc6qB5NskWE/yUR4kzLQO
tGLLWlQe6N7y9lH5g4zRRgDvPku/JnA6ThaQ1eOEb/LPoelCC/doDhtmLWLzFS0o
PDN7SZXjpXb7891z7ONfI3wvnix0QMxeOlCbetpT4fcyQ39sP3fKyVpXjtmNjiY6
V6aDThha+iEPxz6GVQt5XYgmRRV6qHB2i+yGKmKY/BOzdmha+axAlndxacubMG/p
eHurKmTdAb35CU59puvkqRwDeZUvVvZs1L/bAh9HxutOUxg3aNUvfhiUZxmfWvM0
tTrlwgmSrBzeC1OnmjmvR17rLF2ep4ZiqRP/J9bE7c4zCg6/dSiaQ7rYnd7xr2Xd
flor3XWcHJRbpwqXmtrlYfC2gMnJ+KYFb+kVIn8qn+XVqfaPql1qFJ+ikBBD5jy4
NCuIYdo/ifv3njJ67q+1Zt8PW/kYQV88V3lx9dSdEVeeIJPDCQVl1M0hPfLDymk6
G+cLx+17McXZpwHkpxmIQg9dhBH70ib89gRxp9d0AG72B/FLoDhN8bO7k1oF3Eh+
X7i0hrD7PA5LL0PX+aw36QW4TdOhUaNhb6xtxeNG3uX5CJc0Xc19EWLf0bV9+DSG
DzMXdOoArkOlPryo8pqQzX/MxSe2T7QO6LGpXhJpnWYxGs8SacgMbEhjKE9qOY1G
tQt2LXdyB8aI7RaAqx9EmltDbbz07w8Yp0Y7BMyM2ixzHLKSU3ZCUaHI3W24UH7J
RxYIm9KTrNb5zgOalvXUD1v+rQihHGzTUurnmjSK0W/bwVZKGjkBq51qyMX9oYjZ
n4h+XRSrwiCr/rrEQByhtlQALODEI9nOlQjTDv9r0F27vuUrTkCcHom3xM3IsMn+
BQVye06vAjlRmEGv5AyVGYd7kdUJKLESXs1nK9IR0pJXTf84uGxvK2hiyhzFDsOC
3qeJHk3kI2rc5qKfJdNQS6fLVjZN0DN6mYVO9GqGUi//1OBw+2ZrMqSZhRDYUmub
WTd4Fvq6hR8F+y0ITaI1XT32314NI3mspbW6VFKn4Fc/aYCAS4p6A9iHpZQnG2u/
Uh0WqpQ0Ub0QAUz7p3QtjZggShtpWdeq6lDM1It/wGWK6+oaWSvjlOhsnMffMOf9
a0r5FOUVSYQi9B3i09XiiNwA+ZkF+mW2q4tPIEYUl3Z5Fl5HFzilAiPot08m/H0T
hA0QYOe7ktPPYw0Y6cNAuKqxrX2CVTpUpa42iJa/c5SfLBU6tE7V87VRtXmAdlHU
5BVm4OLwBYh6F8vwCB8HYIGbwOV/pmuKhs9DTuRTCGANQKy8BOp149BPyUUzjkO0
Hj76B3ms2q6WRrwL9WKn0jHyPC3Ncol6z18rSU/7j9bw8Q0/hKZ2MHzVR/7ybe4A
hkMGNI2XzzfZZ/jDB5Lex0pvwRP0EwBrvcu+7K4ckpEdzKTazQYLcV4gyGA5/KYQ
6yJusUL/2tZlaxPf9cjj4pfoc0e5qYLbFLuOSNijGwywMjATwEW5N/9VsFsfF9iK
eC775yYBzb6Ik4vdNGUVJC/3BQ9jRCDhEmVKwgGQInHvTCcpHc2XyADh5nHVhfhm
z5f2D5vdNxl4sSGAHGMl4R7srHrRrR/FROJSJlRiNXck18NnoBA69r9k57ZiW+qn
uSTQxINnA6EYZcyv/ZCaL4j9myF5QdIvPHQwFdmuEb1WcUixCuzMiZKFWeXOo//T
yD97VBqFOc7DZc23kqQAzdbJ4ze5/okYbEwC/Yd/votI7oFXSl0VNllMM/wJM3MM
cLPc3pdBr9jPrKOnlWJMkAttcqvMopaiKpw4lCD9utkkf4Ne5HFGdnms62J/wp7R
rm51l/r2bMaET0TF3PNZqwy+zOb/AdXl7j4LtBJvik41Bdnw/uRvavvsUSQ7n0vS
g9lPvl6E92PnMrJmsfPuO99t5NrHUnIilSwISvaa7m8BnroIaHgkkjb8JfxJEQuJ
3268uoVflB3PhjBhndHR4d1GCeDF9BTFXCgDx0fhVs0L2WcD2a/GxDEXCejXizOt
gyvMC0zy5b/kZ1WfWPV2apfojSyokJOYAbVgVBxxVIC1gHgqR69rUXhvBE7NA/nK
JGq+lME7j7fBeajU1uQY8q4a1TQP+uookRd/efwumCf+QMOIrLbSSkOTl9/4D0xG
MTWOK0dNXR9Y90k4OS0trJfNUAoswRNrYYRNofrLW8kv78p8DNGiXOJspprv5YeZ
/FA714GdDm+JWZoS0Txc6UwmIYSwgrrOLikLjOYEEhgAnmhfUSxj3BoiZh+WXFLw
ivazTnDXC39ub/3qDzPaG9r6oASzyG3FL8w0C/coS75nQK/kcCGMy3OkHuzrxeFM
xd+F9VWtUlQdsTJuD8/i1chajScbuJadp+UM5ir0RCaDAuuanvxzqMqrB91Q9AhU
ZFUYjp8LX+vhAmlXYqf36PyGjWTrb92+vZLbVdPdOzW7yCQr7yS7A62R93vRnCxV
ftW4YJSnuu9/1G39ENXAECqyQcG5mrCJi7RDSSXcT0T58/UiE96QdDa2zmyC2SiX
qE39Gs8bsyp3G/3+YAvG6Z4lOKhUNahgnUC3otSkTVxxmHtU86qvPImfpDssp54w
eeHN/r/zlipcsDkaAUHvGhtgrtN0BR1pJyvpOgn9x+PKfZTipTGMIyXVG220f/E7
CIdrmTFAuRzkNcLw+TIC/PJNDmkDSW9tcS2Stm8w5ZKlFg8VQik/VldaDqQ7IgJV
n6cquyuP8TuN49SWCgl43hpnje4To+U2F47Hfkmqdktt4H0btVix/djyk2PNdql0
NBFfUi4RvZxWxkO5ROehqoGc55dKyFMNaX5A806zZcTtfPijtCZkwT+LlrdFu+7h
U7tOu26F41uHlEsxh+8ycCJJVKOOOKcYS3cgT+YdDSc8J2nBxANX7awfY8sISlWW
G5GK5+Qxj3u9mmKDZDLnXlH6ndoECPKHS90RZgMOodbGxKfOK40gXNSlDlO1DBKn
xYvhAIfethoN8DGKFzX6W4vw86pwLehgLIrTTW/BZn9+OYp2F8NzZOh6hkF/ly00
PMwkLvQ3VqkGofro+yZy1aCMFie669acvIT/635T1xX0NKh66pvGgYXARJ2JlBXW
HvTM3Umsti6OCPYwTE2Q+BCzJA8I7Hgj6XwPbjeuT0H9BfVTievpeVxSNu4qaqN5
qgXFkhlY/UQLyhVdImJXbxvuLy/ArRoXl+aReESJBHAogy2e7AKjfCZ0cjhC9/V6
lf4h1015AeuSFJEbGCPbTB/64batM+U938aZy6dtCfSUBqcPQn0o9wY9idqVwGrT
//zrmnLKAjrHaXwVWNCvXO8656LjvyTWG7FPnIKz2o6QabpMosuvyXkr5tlmUvB9
EhMLb1OmMLmcgPeHHjd+Ci3V2UzGkO0MzCJFyY7NDVEmKwMwcDPI4cFmDFg3oYW1
ok9MZfV7NQm+f+jUO9kh1w1xbejebWOXPsY92Xtw2ROfQZrAxFl6Kb/zYvf943mJ
Oi7WmGcm0GPOKM5pVvOzdFIHZY80NT9P5xMldlNhGvnKttpJvTk+ZMvF0oFfvcI+
Cxu46OPwfWgmIUa4JkNJ3jkqOZfE7vDE8fo1/Zl01sbbWAlNsMT3XzOj9rLZ8W0d
HIlIXjwHpfi7BQjnkgCAxkXp3iXCuGelNtUYFIvTqcNY7FFX7Lpp1K1BCYmAhNLp
8HktJaZPDa7Gaijph8datR98fqVr8A2E9BD4tMYMY0XtxRV2kKJ1ctXYk98d262a
7z9d5pELS3is0RyCxqWX4LA6Rrluca5cT0NsIGpWLQuHqsIORzOzszFgFCAk5APT
dWZ38ThcYTuY9J+7jzLdgVeXnC+lKYXBP2Jjc53WAaFl0CWcLkFTGetwO+xcLQ9z
ZU6eD7CHwlyZ/TmQJg1XljR3dfaVa7eJcCIxzisFLTNLemPmHJ/5IhGxrXAIccf4
sEYo1DLXHRaUWFZtWY7QryqkV84RIuQzRsk4c3p56xa7NOQPCVeLJvgVktaFb3Sg
HpXGjMXgwzTuz9HpRw+z5MckhO1FLAntXb+KHWj7W9hDyY8U7U6j0dAvoJP1aq/n
H2cHj/oqwZEyigNZDgxtN6EHztAKCGxxD+xZswxjQZQO3aOB8bkG7ubmZD2S6sip
lm2k+URR3j3NDdEKhDliyS3iT/2vT1BU4EVf/JUAQderd2DtDFCBlP1QVfA/6lam
l2uTkiFbHS0eYHZPOhgbaygO5C5nOV2uLapMSMTlh5dyutNxonDQ2cRynU+EmVaJ
dxjOFzZVy0Oi21U8M10CSD8waKhjlVHim4RlhQ+TPVBw8f1U0BBb2eM/IuPdjrs+
Nkspp2ERTkTjkslGVJC31Ul1KTHbYc05Ye4ovv2RIpRKX2/gqlx/Pp2dzd6bOfiA
CeiZI8946fZAHfckPEzruE6dDb4iEwlHwG6gUsKAnuNWUKPLkVzjFcghHsuF7A94
ghmRmyAmTSPH3RmNpMS+iFA9m5G16CEKCSmRKwRFFa+xHKHXXkdsoSbs33rwByXJ
v6ot+J57parTew97n1dOf4eQ8SXgN9tTwsW2FgR6qIrTKXoKe5B1k3pgz0U1Xovr
0UbzEoN49BThd7Gebeett6QNDItwT7L2sYXmS/TVcf2S3QslbbaMN9NKJgFZPt6i
Uud8hNxZQWCk5JshWBVDmeTM5VNhTOBfd9+rd1El/OUDcFNfmXr5EGqnbMtH1Dzj
Zdqi+YAt7oY+8npdiLnvCysIJCIwn62fS9UwHs6xBL/J2H51X9QwLsrXjvpogbe2
Q3axK/FjVJj39R9cPdLMFQq3NVgtN2xoBhtrkcCkdNCVboy4bt6nCSv29fS6yLj2
JAIL3jnzj3GPDVc+OvXVGthQbuL4NTI7IxfATSXoXw1Fnf1dkQixwYuraUqQOBcc
OH3DXBexZUYjv2olSsBcwUYFVgT0nwNXgseOzt2bTVPPVw9bV4SJTqHBHqH4gbgc
X7lLYSMUzrpPxOs5LYIBSsM0J1IOPn3UBQcrMP+tXnwuoqJtnXjv9OV91J/YvXYN
8taWBIK5j/hsEvf7DpC4047kNO2WsedOER0V0qj+bGzu0efUnIRCfqBoandD+wuo
ihIF9Wg83doYb/LvMKahjPQInPoeZNjULcvIRmJMfahe3xlGzeCgbCPcyDPUeGuG
ZoK2VBFdo9aScbVyu8jEThptpQvXJm3qxM2OCIgKG5WKvOcuvrtfaRrNuZcQjrMV
vZlC6O3bwJ5wF79KeLXv2oZT/mqn7DpxW3zvtvt5kjrelZ07Soac2rePb5PJo4wW
98fcbgndq6UxsRb2UvVIO5P75yr+jb+jjD7s12MVpukEIrpZjZLT+2gn/4LGODOe
HCLv8sYQMZpq8n668Ouhf5rjLx1gkOTayx2HtdHl500Nht9ryTL1D5sZ1ZibS+/K
LmkZbaKFwUz9VJzJesNT94hnKWzdwizgwy7FrEW1BhCah4or5Wjot2FnthLxDVrB
QEfBARiSQQSzQr3RNQ5dzPJBk04GyuNWWXVL+7VPoJoTryiZwojYvxnB8s0zv5Qc
NeVj42knJ0SrMao0maOJPBj8DcwdxJqG+ocrQIqX2g2dnWh8DDNvg7NAd2DCgRM2
oAi4O75cLk+16SiJZhRE1oyt1k35f4N7mBzB2NNwSXSrXoF9zIZTx5r8Wwc0REJc
PLyB/S5EBgGpahOkmyUFbEHqLEGbf08Vk7aIbGXTJYF7mO5dr0azqyUZQVRzEE7R
dj4W0mlbTvo8oRPqzQKh7EVny8ClpI/k/ySQcBk8lZebh3kbhcgVXFRuedLdoL4/
KjGUjKhvTPKtjbKzJoaXjcowrNWZ86/kA7YMF0wqUoB26K9sNegPkXxuPdUN/iBv
vtNFgcYp3RpTodBJ2ZD63kExeswCyAukpcotO6YeJJfY6OOk14KxuQ2/Qf2fU8Za
cNhvu/abdmcXIDClS0u82GFwqeIGU+vbjtv5Ov9mVqYyegXmfwsRscQ0beqxUlLg
zkV69oMdV+/o7HJVGWZ2G3q5A3goowpG4n+juV1gsvxeludXrSEAOn1NL2VqF//0
oN0vcnWr8DKIRARHfLBkFy/hCCcFR4fTwC6aStednP9ELY67dmMYmfi9QRZJGQs2
O1QPrHAGX+d/CTwmlQ3GfpBUDNsZJaSq91KtsmAPMrBQF+PXhC7hZzS/VnQeePp3
Q3TAuUkcSmSWwDL71lWScfBA4AH6yQvg6PijsZARzoKZMmuLOMhuKIhwiI2DovpP
teSypETYKXMWWmeA+YFxm7p474w/BpkGfQc3WhgLnS8JqjNw8HGORdWg2gw+e8sn
9LrMYzuf5hQWHbrgoFchjcIXeC0o3Hmk3ZWbKkMnCYpLlVUEiB3KjdaTdLTr/nD/
SnlUkKQ2YbCxiPs6JqpQfMIiwZPhZlZP8W5qsGqVE5Mwmx9UXQqMZ/pOEGw8Zznc
wkCjYtxRc7fFAnM+dmLuDTLHlzeoshqVMHJpJq0oR2zUjLjvihVfsRq+frOjXknS
b3QB4RJw4aBmwJm4kdmgaZ9M41O9XFw0pD9Bis0+nazlW764wOVUZ8dDO2ek+DUv
4E9JSfYOh8OUCXWxX992zSVX10+UqIBHl71vnMz45BfVwiVOJzOl12gUl3kqVj9q
kQGNYrLAeUicroU26CFM4NaoWSS4zdXg5ms9z/mypiA2RmAEWrAuDa2VKrSmrkpV
N+YZNWSJcl05SYY2007NfMOTooVWyAIhBRVdKQrzrMIbeQGsXCGfk3L3OSwGGV3C
PA0sjcG9XC/zVaawtcpM9DfpuGuVy+TxzNnT0kanCZ5WV1fb8lWwERXh70/iznY5
V564jo113TaA9Y8SpMLCE/ntjRJrM+onn8cn1cnJXQWlH2MhfFwGCx29iq0lzu11
NO8+nUEJCIOTYAwsMD84zUfcUA/yHhp3tbLoy1kwWA/9tv6v/S5nO6xyjcR7fcXH
Z1clco4vr0hZ+Cn2u2lFeciBBkegy1SMa1sIoe22ZEh5TWhLeMeIoDOQlJqc9bDb
0Q6VQjcHTNdmF1G19DqCYTO2RP7ziVzctl2qmyJGenL24bwnDmFWwwTTQPRrc6XZ
uAvluw+04yf/wckkVk01ryx8TKI/MFaDCz46h8fwYmLluq4Uda7Tp7n+5j3jndL6
22ql8Beh//BtRajI5Egtz/9Tgl/Vbu+DxE0E6fazxR8+XL02j5y8yVCf/KywhuxU
GwC5m3++oUv0hMiF4waxGJO6UhSZqHU8txWauXfo68FW0YodR1VmhysolKgekm+r
J2N/GSAWs5aDfiq/eEMhZHqiHQzZ6EuDjpJuP37TfSVC3R9WdFFtc2qB/zFZH/t8
k3YDOD8P5i0o1WHnamumjv3ppxNcf8E7F0UTcDPr+U9aNVtdec6vVQxAySoxGVo+
j1hfOUHEAk3a9WbxzZ0b6Q+2b+ioGF/ExvlBzTrOQrse/I4e64GcR1yFvSFtQ2WZ
mdZG/lS+OUrRB0q5M1pLfgfMSm/P2v8mrNzx3ZvKQb/m9NVZgqfpv06XErwDpi9b
BSAzLnl+HhQ12n7bFH8NeaGCqMGgAZmjmowd3CZTbO5jfvb//Da2EqrnSl8YiL/C
U3c4/XFl6r711SJ9LbtGCZD/tpdw/+nfQM7UxNeluL+wqBnD8q1ZYng2tvv/U+7T
a+vCImzdHLJhbVaEol0dDYOSwEcr3+fOP7mNMiHVd/07+jWAkxSCAXLSmvmb/MOQ
1cbZg7yex+XUDMNfufxocdB//t2SW6ZBAIFXpYLFgUYXd0XHHVJxlytq/t6R/ObH
P9yHBaz1/bnKJX7RUm4cJ+y57xrhatgdcERptohZZxRxyBukTEsoYzhKe+kPyFeI
3qkLscKqfM6HAVWIWxF79qZ4nTkwc6m2LNavGQZydPUNrbtROdoC6dyV0T5m4Vxg
4Pa80u0EbA9v2mXCGu4nEm28G4K64si0XWvQ/+4dd9I4dBOxFh1xd/06PkEbJiDE
JuiE6HYg/nBbHTpAs831GkvUZ10zwuryO7SsWsYi28tAWq23MYqhVgHxcZivwCjo
yD8dgjAiRRlDJUMKWYrFA2RORxMK3UoyPlxEXHHtbHrNuLNiL2PeRRSkQguAOJK7
+S/PajkvpkOd50faAW0QSBYn7TtYopreCX69RuolOiGwBCILmcux8SHBxkXMbOjP
GZCrFxpEBx68MJuUCUCpm02R4xgKeEBmgDE4FylXY7hpYCcoOCYRzIZwiy/gDbDR
3YfUhqmEnRMssFVcscBcD7YEngRhJ07YgUpeCq3JHRHWXKi0ckFhEP/bmiNv1rzk
eYZHD7g6G3GYBzcafWdY26mmweBYWqb533cWWdwpgQ3iAZ9guBNdUcqomkH16CGW
yF/wvAr4ZvlYhdsL9FxbuCpys1np4m6lk9UFRDG7iqiMWXc6gq80wymfzlgH6tJk
8peT+IH8RDpJqnuNR/3GTbmVIPHLPLL6bzhfp3aK4VCGtmqEVvz+Q1nEXjSc8HeD
c0fKeSzleNRVJSLXf3OOsk1NEZs8Lp78/uqBImwml5rY0VyuqbyjrrgK/KVrVAf7
6IOPD4K1tjaZ9cxPnEjcz4WqKyvJ1okwsL87AKHEIakBEh13cBNSGO8OsN1fd9ab
05ZZ51m+lPEz1jxwZArmcF2fhuAHTV3zyXU5IDOYXyy1HIo54Ru8YwCMc1fThMvG
xkz42ZZYSpccJtjdiMIZguntAAriHXAFCZvPXG2xu0CfPiSrP4t+ZZ89qmPtmOSr
KrpMRtqZFt3sG4LP1ZoWDuoWaYJwB3KyERUWC+FVdvPoegijyU2sJQB50KSanvHV
0E6KS24q8Vguha3IahJR1zk1OnZkrvscECHokUO1cTFEIgJ2WKvz2+P+jNE5tQxZ
451LT6rwd7lxucJV0nP7gNoITi7fr/T2opN3p/8qya6weXDM3a/eaZU1anXMr3Ve
b0kIyrQC9uVn3OFN7Nbw9x1TTfS61Db1tEX42VdGw2Dqn8MOrklaskdgPX6quDKc
+RrzpORsKDZYfjwQwahC99GF/bYY2rVIg4r8E6h/99NjpoBOrQHMXpbSl0p6kk8z
SivZrjy+Ue5wliVAgp/cdnjRu0uE77p+Qzmmf+d9JnmfiaUGT/lj7n+Ori9g3K1W
LgALCWe7gu05POP4xHLnc2VHFcKZgGCxo89tMWgso6FwfR92bkocA2unQ2KPxlXL
nDdVNxVE6p8zPzl9CYzchPxrftV5cPaAaiNBcGaLx6eFmSrWdJu3IzlKvgqQnW2p
ThzCmlNpCuWJCcvF4ePB0jd5n17Jn1ongo1mY0IbSgtGb9rVIbNihFateI7wwdhW
R8YJKkTKIwtNqTVbZwMSpDVHS96lDqRxTfsxoEIeuomJHb6vj5H61Nb1LrPKBPgk
AGER4L2l6U9rsIsyItS+uRJFzgVgRs0kXWBHIEVFUe0GsbD4Rsq/B92pcLGpcbO8
dBKwBnEEDVmSaUvdGpgBitoLFfNxtHwnYLERcMtpNOkSo/oZhEcUk12RjNy1xAfQ
k/vDBumBrYLCpMZURbCSkBfoqWMNe68mT+Te+ZtOZf6LaScmBtFrUOETNB9lmZ7K
LIFOgyr+qAYn5D0W3v0LPkZhGKBad/acVg7FzVf2SNYrx+7ZHzi+vxtx29807DRz
ged8rxeSOhwjcNhtbCmEF7EqrUbK7W0W40CldMv6opPkoXVuoPTKiLg1GM/k87XT
61XPrJIVbJs+A6VKS14yhnla5bjPiMZlEkKc8z0305jZDOmrx5n7nixid2p0xIUM
3baDsr56ScRDfWFWV8goip0VZABEdJ3AtVKDYv3/Sfgls6c8M8FwOLE/c7dwuB9m
JL6K3NER+tHiV396TxHC0l/ZN6EkG54IuFAU9UjMAjKAwSLdIoRxr5oNCYZTi3zZ
yRWXsgOwYPNSAqhS/sWa44TAqCJGxEf1Sutn1a0m5kYvbyCx4tcvmTp9ZZ7oT18W
iPW1i0w4pA0xRqAYJUD9lgMywEF3XR8pw8XvJUti4RbNl6GXbJYtdgptqTifb4se
EcM3VZv7qr7mvxLNN+YC3MPBZwrFHif14FVHa4ZDhdVeGWNghGF16mdHLRDq7tV4
rU427/VETYdKoWN4OkrnP2zHAFqaF4rAT9CHXeFAW36VZ7KMMV7fciwlyw0BkcH/
ZboPzivlWUBj9gNO5G87YpGVtEtnb+pwJ6sMU2tkCGXHvCoVOmINBIUDqier4Eh4
GqkYUFHGTcWblBocBwrXvnT2Uzj8xgZCKgAzLySvM2hUM7y4JpiZxOWRGk71revm
VLNwaVag9EwKfWHY+NJUPxvfC3UWQJvJs/vwOsxukJH/5O7U2IDXZO8uhmpQtsvn
lZVlDsCdL0UEPuIxiGoQZeOcCDmsfVK+AN7TJOZOFe13Pgooed219xDrGVdQQBBL
QD/EslofzL60pCgHN4Vqm+eZ6tDpIivHlyYk5ruU2/hRma9FpYd3vD6YNoCQARFG
0Z7qPpcLylcw0kjplmfCDuOIOn6sPhqQvBoWg0zsGKWUrUvwYD/hNycUaYKkSp1g
v0DBRxJbEELiot0tZAdvSsXu3vpeSHIsYKTYpI2Co42Z2I5jNsc74xLZo3q3/4cm
M675kaB0RSX2RPcdlOX6Clwyv2Jrjg1/jLJ+J+yl/RQeK21UE0ZBIhDmoaK+kQzD
L6O2xGjz1EoXsJOs9N23PRpzpmNMYnK6lo2eAC4IROkeGkbn0NiX7RihkqjHT5Z5
NdWOrjT9DkxPYJMMOEUO9mfAbbR+s8TqnsXAiBGkOZQxJAF27Ebaz+CRuOhsLnUa
QDfS6dkorqdeI6AeqvG+PeI14bnmqG7hziCNBJ7RIJYQs3GcU9Fhsz4puWSqyaMB
6xQ1pE9mL8YyIojpcU4Xy4C2yImpaUFsWqRSqaOt5F1eHhTJ+vdvitl8S03H7gwC
VAD/VoovVkrUAf9Eprtk8y/HUJQr31bzGk+0isWdGo69ZrvOyowwI8swXGWrBCl2
Mf+scwuVTW05wg+2Fymw6jAz6qTIRMHoqGxDlSvL6qJbfgwr2NIoaFjdiwj51jqw
5BTHYkJH5QPfh59urFUp95hXsPnMatyj+OwwaLfW53PusDf/6ZLi+i/F4s/9dv6s
7QFABbYtGRzqqej0r+dYpJkprxA+fIOHArrNINoRH+/FvZOfOB9OsBikGGOxSf6E
WZW5vHW0ycN79fezcZ8ehZp0JCLKaf/x/hl+KxDlZH5DzQGEa1BekI3aGj6e75sv
DPowJ5MSxhQRo0cc67oal+TjzGstW6Yz0eDmk3muhDTsKOrZw+Zzd5cWj8FfONoN
gWbSoal2ojZ9kfNKYMvqJ5XNquA5tag2T8oWIPZaorA1DG3TWcPhI80Ke8EfG7/E
+XC6Gf6IyHXPhIAuYZfeuaOwJM3B2VgWp+YnStagZNxl1nGsfsU6nYRegoxyurFT
hmhta1LRRtrzqyZlijkXY1zIzPol7DuQylFvdRUST8cea5CJ9ntyhNpgMflX/7Sj
/hXchu1QVMJ6YpKQgK6EoUXzx0sl3WE6WoCMqTLLt+ej5wTkySoibP6/eVMHGoH4
z3jFjNHvzKOvlbbEckvoEhBRxF9MZs49acA/7VkV/rsD/sNQjFnI+mEoInlAGC7c
NPBR7fmxLfUHh4KWDpp4hNnMMXN9v+daCOFrtipevW6dUP/r+ZYoD5/txuMWZTnC
8Cwiwf3L2EzqRxIMCSSAYghJEg/CDniSFqP2sT7+ng/GoQtWgsbNiRggfyT+8SK6
rltpYq/cNG+6jnc/7HYe+VE0MFweNjkSfDY98cNs+aBW4wAFuhfZ+3Rn4pLG3PZ0
y4taYeB6QQejavsImONM8lr+Syvj2eVA+9F+aBNw8wQmGW3GPYVJeBvHKiYL1VAV
RUn1qovbAWztlOe8X6vPImeekiMgYCmGVulLcS0VUyB5By+BS9acnme+vVRE1uG0
epxseVyw7/fRgEoaeghSimM+YBPbpIxwgAuB6fU52Dasq0/W8klpdH4N9K9XKNlT
Yk3YRMzXRuro45iO1rCmiyqmFXAtX0hGu8u8v7KOIpawZx6yxAAdUp548US1k6u8
vZIWZvYLqeBRwUS5Hu+4nu/Ev6CLJJb+6bDP8yPr+GDLthbAOjpR5WwZnDjWYjB8
agGszQ6osE979WZ31heX/QejW2Et0eZTA8DCzJyAhxbUZK449AzPELShGH8CXyBL
2016Jbaq5bKAQ5+xWe7uFcvk9XPVlSvbBIDjXfvJFFzcMorjeHbbUPZQwTcIgxuA
Jpf3DqkWiAlrFeAJ1r+ERb+jIgZfOpvAXM3bPEUu1YoyaVnpdO3nwr7hDrRvj/Nu
kUl5KkxCxm6/N3/Frwgk2frXsFVsM/VOp8tu9hhhXAv7eVLIoiKrAG8FOwLRHbfV
/cGQcBQTBMwsQ+yYxmTIBBf2eMLZpzh7gWnKIybXpzB6/SZRXIaa+H+ThhvNJ5RV
7LnxCXyg5TqrzauENhlr+aNShgV9yUBPMQhuI+7i/EpSz0PqWbYGfEYex/8sauLQ
H04nGNsXwUoobu6GzlfKoanEB7pcF+8YpKKTu60dIl7rZSyfvZEa87F6M/3HhAg0
a2VyimCLoSGvfMI2LbzM4sxuW0fQc7VNqal2pNO8Udd8ILtxYI0ab95htqEQmPFA
wPF6jBTyBmSx2+39zSdTd6i+IOoUPKYBJ5N3g+Jl6BzOOmG+u2PJ8YPxbeIXxMt8
mi/UYYTeaDFZjGT83ejpUNi4GQ2P/yTQFBvoy8PSIoChOMpb7pYMgxLK3cSws8vZ
oGCJH1SH50iakw4eeU0zSw2WRcD6ClWrv+FYw+AettIP1z41zOdRaYg0HJsMjvbd
aOohoXWXOQjwbBsV3qq8ajJ3upJNqo8G17VA1g9dHG+815LXupzdWGEIowuysgH7
H+9sNGWv983xp4QFWj4yFdZyUgDT292hWEJlt106LwanSlZCjvdlZhvk/J/vg4kT
xU6MMBIZRstfPsygXHp6CspIfuprWn7sZkoNy+hii5yNnHm2kuZ8WXk9b1MGVQQ/
8wib3jgwFlvxyfX0e1TpJlWINR5ZqCRZ5Qwc5qd4qsU+pml+f5VwxTBQyLLbO8Mz
sEixrjvbmhsLOTBXsG5D8h31BJ7/PcBcFJ290SZmhRxDY6S8exugoyx4w3q4LEFE
Qb67E1a2XTqLCwqs6enZAy88RxmJzxA6PJgFQm9JuPUhfRZqJ9K1WQEV6ZopVqaN
lAiwgyU3/CKxU4IoeCb8atTaHc3AUWntImhwZKju3AinUGibl1FepyBYk8SE6CnR
t/LKU/Uzwu0BDKStsx7vtEWbQU5BuRwHd1as+GIJ9xAjaA9G/5PhzGCJYtNFOdkA
nLG31vrgmHxksrYkrlCr1oAwSZ7ODSa8w16HMBlNsvbu5iMJ2mcJQlZPfGKSwTbX
oQJ+Xr2yd1FZIgYPQF5Thce/3X1uO5F13oknHbUJitIlBPGwvyGQlUeKHXB3VyNL
XN1O9jG7pHMPKAml0PuR+BXPoCUpjtYE973Ff9qAvjZ+icBKGEbqLtPZZzchnGWi
sbDPIYKHWsZRAlAEfI71MhQamy8VNAHN4UTvV1wy1aTDBSjAAL8oKSpU1NMe8/oi
JnIR6jhWraH0q60C+OUMjXv0EbVCX8HRMc9x6H+e7LDCGMVtN0l8eKa80Sf6YBGP
HZaK8wczh/mN/vDE2qVhGNylNzGZNlWzMmNSlUYnqmKyn5dZftexNIcjtp+smQyJ
ojaPMwFRwgp68ip36GGzg7cJ7Zp+J6OV9yX8BERmwLFA5Bf9Ulh20VRLDbCOcyjn
znkeyMzGV77hY1RjWp2UBmy7nnJCOr5B1ypSVKAcTy72XQqn+2n0xrZ0x9qHNG+E
8QQ6HhTD0zp85SIE+jnSfkw9VgIn5sicg7QAZJN5Nx6x6aU4f20/8fx2VUk6p0cu
blFO/mddkY3IjuLf9YifU3/DEfkYxXFEL9v5Wv5Cdva4Eg96bs3HXZxi+egY/l5+
oZJjZuf9x01a9sTB+9zeRsTF8QbN4Tck/KV5CXiErmevazYB4tK3ZFWl500NqVe8
H8w10A9BHvwdby2C2gqzx1I4XL2TYQ34PEzMMIr9MgpLDVfnhfHJ1qztXm6ddw5j
Ur0YFWA6STVB5GPq6W+pvBJZ13GsWuJQhbNBcE/9uDoKw9MAGX66UZ8BcqktKMjx
AlwTNjv1HUKiOfqUc0wcVujo+B6C5vC6X9k/5WA2KEIWrE7Jnm6RUZf0sGXY6/EK
8p3NiuV5C+K5oFbu3Y2MWmmTw6F2lHz3SbVAVvI2DbZbUOgZwTMINp78pN7apB02
1VVRspHKz2Z2o98KwVwC1erhFlaMykbi+oRmUy0v0zI0kr/x2zBKT/27Xqx9EVsP
fQTnaK48gxgBujFx0Lvb+V47JoOIeI3YvER8rTYUapSxg3CjB2nRhZv1VZtU/ghD
mqvNSIDjS+C7F8nxDirFvpIR2IhAQ0acN/DuDSgDUT4M6rwQFXKVrV5wrcP18rsu
GyUVXoPKfmpwTo8S9AnOm24UYxxGeD19XOgHSu46IlWz22gmGVYcceBr0T0plKe/
v6KE2mk9EkQeZnuXRjyHbZ5yTDYCChSQvXAvjIJoTpRQxjUv0NLACepNW/xrYiyI
ehdHnx2A9dydeWZ5vNNdD6f73WDbEtQf5UNXbnLb77xjUN+dyLbAapyBGkOKSDEt
G1nsLNO3L523l8LUaNi6i/CaNy0vbzfkLMcE61B1INDvNwOp81DCIOc4JiL3vTjg
Qvm5meami1VIWFogbEj+nKM8JEdG85cIcsvFO1f/w6GPkuZlwTE5Q3eFP9thLKQ2
cxDzGuGxi6SFCyPrStFOZsznzyKC+RA0F1UFeN0V5F5zmUqrvLgPAVNw9dX7QX6L
FF0vHk2VV/3KfHf7rwHxpKdJADF+XM61HUduF2hQJNfnEqtEzsFlfDL6Yh9fBHG8
50RgyhzbwZX4egzO51LVht3uTIuQ7vFBQw5DEKKtKRqhjLOZyk81WOvtLX6NnBs6
oDb49G+ewJQk9+ctJcmDobrMuT39zdsHz9FCUAoX004+u2sg+RlS7D6qto25wnga
7XRgud3N2mEY8sp/PNRpNxpUd8q8khkIz7jYpAIeWggcVn54jAYaBwiYKTKl+eF0
sA4af+tIHT/n8BWOEFQMjm7AR79569Iyd3cObkDm6erGBZ6wASoK8AC0aFp4LT5X
2aJ2aK83FK6ZN1Uwl6S1FpMCFLleL9Uj9zXKsMbQrdJK2jIG104hEvldWPx+fkLM
ndelqCkPVM39zR+R1wdBZqJdlvjxxFmQtYzogYUaPXk59dVpE5k6aH5HcwVhw4Sz
zvh7uq3W4wk5AOo20R0MnpZQGTQKtoZONnef6NkzcpzQHgXzdzuQVNZmN1bza0+R
GD+CB1Sl+Jro+gM8F9MNTvecy2a4dG1iHpT7dXz25WyVVAZLNKDask/qW8bP1HOO
R/ti2cFUiWPK+nvmU+OG6KKdItJmUzwHSYFTF7SBFoJKD5sH1Z2e5ThPTK+Ouy6g
Vf+wEQeucQnwENbor6pLhStLq33DR+V/1DJVbvZNsm4BqVAvdN/QkglSLuaS+hLj
75EbWtNvMyIB/Hf7387g1UPB6+dFrSE3CJvAzzC/2TZhv93C0hcpOQqlB7mbk8ZY
AYoOzgH7KCdUvSNeuKVLDHreaK1xySvAQiuoYos8gEz4Csnqjkrs0u+jNBmEkIEy
COe1JXvSrQUEmJDx/ZOo3+ZI5C96vL9arQiezVggbsI1hK2GzTNeGU8JBxq4HSJ1
oF23X9iHHy3UEEeiIupAgFTbIbWlfND5va/q835t4qBrhkz0Cd59iBNonF6U24BR
4yDInxjURsd3nUy1ssKku1MurMpZrx36GBv9Te++kVT+Y9b+/UK6+ESFFJI1LMMd
G8+KpSCatEEtqFZTdQCilVLUm5Ng8wBQyHMcwuyZNFMnY/UcrkXs8dOaBITISda9
pxPBari5pvhZtY8Tna+fz1TYidtTw2e6qKLYATJtvu4z+gSXUerrQtmUL+WASArC
xV64mKCdgyRrYrWUmMXpIDPus1EH5j4U8AkvSdbeI2yCqjMeY1HoUSdXyN68e+oj
xDccPvVYbf07VUuQGi8yPQz7zTr29ZThxilpeXNwhf85E0of8AT5dOsBP6PbNtM6
8H5+4LnwZPeHV+iRgdOc098p6Z/l00HgWiJ6T2JHNfp6wYlwZSycax4zMN+PF/DL
As9Sv30PtWGLP1nd/zANS4FZdtaVbeN3TFKpQyUAqCHA3tj0GY6AchqKp73yp4gC
9GOmisJj1ly8tdc+1LzcqqmmcIUeVXnb3oeU5FG3a+C8p7ZVXPkI9WSBzfVyydF4
66aD0htyXCsDNgNh1EqrRJOclCKdOq3HVtBJ9dvAMo6htFMjQPmrrFINsQyPix+G
4AYUf1ZhlN+tUf3ac9d8NTGzoPnEZo0LEGIVExXyf0Cqta7Uv4MkuRxuQDojx/Qn
p1rwnrNJTHlGktd9o4A1E78eoJ9aWLeT5apinGrVr5WPeCjixBARE16trK2JOIEf
Bqs5WIPrS9TDOJ8uOdsQSZ7FsDzfWH8KS0Qg7VXpaQNaOs1w5clpJvjcVCTZm9I4
lucKNEWahC2+uowzLYpBv31gBr+uwyp3aSAF7/O4N/KMPeDNqidNoVjgleVhOAio
/JXntwwt2J+aK5aLsEvgfa7hfr3gra24M8Fe9Pnq8AMSSGBPfc81wK/pekxFwceb
6srTNKhqkY2QSflxSy1IElN9M6iqgwS7FMwkeVnJZPUXn3PB15rMLdJDNKN226hZ
4pfdxC7VZn230ZPrlcjPtnNWhUWae8CfboyDhv6KsldR8rtN3eQJoV8o1cZfZpFh
bPo4vU9khAQ7Tt5in86GMsiece20qzdrTX96fa2oaldupxBmIDrTEInkpZnGwmra
oDsEgRE/Inv61JieLu0qntnMYHI+cG7r33r2VgbSpTdnGQOyy1sU+4s43MW+FAUM
4Yll6rT7Bjjfhcl3lRC625QjhhgKyylbmQSb4GsB2+9c0WeyaDj9/4j4837EOdpX
cMtXsBwjp17XxGdNYeYt2ZXvany+8UU9f+zCRLuLyy5OS698w4zI0LERZ67o+Jwy
yMBOlAO8PRTuakZrk4sy1MMIAOOnwaafiSnqimlmwJBgYhOwkBrgwQVdAZiThYSW
Zk9z01O712hiqkKvJcquJhkMTiyDTatuyiG0qzatn4mdAqG4zV2H7BBjShArfpf1
BohqRLUJtomCkDnXdd90ckv0Nheh6Tnxpy0Zb8pEPHfB8cVvXmTOjpdk/PTLUdVq
tw3IenUGDeZR6B2SPkAWHDJJeIc1nUlsDAMVg9YSIZnZzz3aA/PafMP2g9SaJ84s
NN+GxcHfQO1KZMKkw4oyBtDR2ubtWPZdL/INdXve1rxk082rsxtbIF+nbuy5Ccg+
I7yQ5dSJKH7Cx26QOjZqotD9WBSAtUWJUsBfrcJR1laHLzowSlj/Vo2XdcuAAmDP
rGcECoQkVqGwOqM3yoRVX6tb5x+oMgM6xxy6jzBCrMQ+c2jRuaEg/eF7YCUfcKKG
EVdH+oxXdi98OC9PjKdVvcK22UanSKBiIb0INhRrSiZrpnvGE+EwIAHosNsgliB0
gU1BBZk8vVEOIHQvFbwodbePS0Z5IoDQ5QQCoar35G1aXqk/PyFzviMqyp8Zdz/u
GC7LXTYWJlVBvLt+JTY4tEqxjdFTJDl/a2TRNWlGnSVDBEhSRscSDmCd5nXp3trg
ijVwXqpT0Bhb2+4r4NumwiGxatP4eeHoUot4O2+2MHAXqMNEGBqlAkY/jVA7x8QG
/P3hGiA3ZfPnl8Q5ActBcv5HjhNS3hgjOKkuhxshcYw1twFlzLbi96rR3Z7ip1m0
wSUHKDpneEM/IgZtmL4EEZCYaCSpSb42ZAnfaFgHMz8GE+KK66wo9LZThnZzXqWD
zG+ksdetYiEiVT2pNkDaGdZDziEobcUPeBU5YjnjFfBpgQUjPiXhSjZyIeg+KpY6
0Dh7ey7rbciiyvhanqmyr/5p8rERlbsLP2mID1SEB2cZag3qjMfkPFzY4JSaBg7z
sR0a+bposw3nI7GToeDcCs7iCqKJE6an3QDZl8YB5TloBk6RV1LrNmz2OLc5rK7c
rsYMKG3JhQKunZYFgpQlg0X8K6GtY6s1wFdxot2WkNg1yyzX9aHofOhcaBSCu3Rz
xTUYq0AnXWuSmxe1woM+JynBLD3535QZHfM5wZAwQQO7FZav34AE1eQVqlQle7vf
hTAGZrP/xZekBzUnd5ZBfgc99cHIP0FTZwj++11+DbddSpd+dgsRAapUH/oaMpoE
b/qi45u9xvXc/7mf9DV0cAm1NzLerNxkYNiTmy5ghgmoO0vIX/QR3NuRjGlFdNa7
L7Z372RktYpHEyq7jd2hNBsbKSSCB6tvwmGXnB9ymaxVpOOy7hxHClM21pSBLgtw
dXk6AXH4rOklM7KFgM1kCCUQarLo+Djm4TfwS9c2EO5Rw5JlPTB6V4thfqT+nEar
JgHptEIjeAMmAOGnIvSCy1wS6VeMktCH5xfFqxeOPObxjFNQ+Ss8MR4+eqgrVCmH
v4hfpQbfi5W1tmRYNtYRbCNW3aN0ZCEP225xmoxtsvkG/qt3AZ7q6JMjb6ourk+w
doKS3xw3HP2EnsnPDFvNjafVPolNr3swituoPkZ0C9FjCiXCLh23F3rWBJ3XImLQ
vw53DkoBWuSONoltYF2+TyrodEtARATfFGvX64ISIUfe2OsNzXV6Sk5whDi88Yif
7vb5T+65QZN5A6HjZekRMjZb6EnkqV0je3HsE9DeDU1Saj/JSSaGk5bqHPC107lE
K8Z9R/Dd7kXmw8WGXHR1xeJBtB3DQd97fAj79i2mk3e03d4wqZp7Ok1BfkOUrNXN
p8AqbGCoy3qdXmj+AkznValw58g7L5jypo2cDW//qUX9QBKkbry86uFY8nbnGhEK
CiRt2QoLT6rIazobgTECCEFVlPImPtW2zA8Z57jozIyH1xltyO3PIT1zVZUudkpr
vh+4xESzrMCWLLTBqZRxnJIrWtvqEPkreCd8j6d3HCoVDyeEvB+SlrePXlmdm5Aj
MX+5ZORNLD4po98rr3CHt8F8oOcMHVy5PdgbLvHNZzgV1C5FWrzuFhR/m1kw3NAV
Jwq4eZ/BKw+yP2CP+OlZiPvWxqP7MJ5UC8b0DERp0kubi+HpoC7xvr565HP/uMJ9
hTUksEGa3pZ+4lW6x9m1mj6rvH8NpcmMrlJUQjCRDgP/Pfs3CZOIQtX+JftTfq9K
hggYtn1R5aK4cOI98UPQNVmDZLKH4l4MqJrjwo0NO3MxoQoU4MfHypJvSauf0O4L
BGPAZNrhkVS/E/uTlUWuaqJjzEbAL8YCZFSkmow6OB2Yx9zg2B/A9ReGBGbCPVBe
68tOBecI6D6qqxa2AcxPb5on/7KIiIZ/ksCtqV6iMyicCwZpzL7MWhba5Bst4isB
IHuw8ABbyURNcBOHTEAdSoqqYaJFehtreoKtdwyUCFlDnH7yUd1ISeSCnjDDuxjy
hJWPu5Mx5taZDIyeJQiEn4wxKEhUSGOSceowLEkD5+trm6AU6Z0sMLVeut7XfLMJ
f5dmnG2pMOdYCzdNVcNxo9MXarFRRmGT6sX/OLgl8b2jYQR6Vv6JC5y6/VSiL84l
IKYdXA+xSlmEyY3QjWewvRomMBQ/nmSmFNqneU4M/UI7ubJkWiubHaoXb+PDK20x
byL/WCZ237MaEyi6mL2gfNh4V6GBz/h5Ni7oIYbomzvDXreNtl87YqaxwJA8R9bC
O7SSDQIudNbbHWAHPPFpErv97yMGiKCmO7Q3/Pl4SJ2L+Vpzg817XUNHWoM6nhy7
5S7e/QKLz4pIfNouwF+hlpazQyLZS/uUz9NerhxO+8QfT2GqayQ7INEYNc3ccTPE
QHvY6CSv48pSZYljt+FsJ+YG90uJMhnJWg5tk6TQwq/i8MVfbFQplhhpBwI6Dc19
XrtJlB0iQhikdTkA2GKCRRZmT8WExUcKc2ks1s1bnW+lyg96DoSeIV2L9IBx0y0k
U0YVuYX0QESNgf6En8LHffcz+GAcoRKjOYVJp43QsauOQZQy8CD7MobK3Mu4Baxg
XjlDYU0VW977NxwXoPtALmaVHVmaNUXcqNT92bKZ+b5ZhQceBkVRAAINMCm06n8Q
cuYtO7uJsjCku9jECrqysBZpQI+M9nVbNqfTNwrEW5/VeehOAloiiDKfVWKNWT3b
vPML96ZvSnVMq8KOFDAcfO36v1tOLfQw0rttFB1rVJqeZP5H9FZzMwKqNy4Olhe8
slV4+fLwYJgZNcnFPznMvB9pQfX6DOQI6Si1NIMkY09kU9nZRxtZYgqTzJz5vWvX
dGWqocE2Y4fouqcNP1RK9wj6bwbIbcy38gNwzvAacKvOtsqTR2vk5pIKJTHARrjN
qJLpFbOkplcZyovVDiomqv/Sk/osVc75iTAr4Y30bB9qLsb6aBT/LZswToIOSJZA
TIUFiohD8eYZQtGfmk9T8Kggc54qwAngPl+zOyAvcGYLUm5xo5AvDuy05BGVEGWr
u8e4NASBEjuMIn1RAF8/Hzq6jqY5VSEkmypwpHJavAouLRPAeBUlPTP7nmH5Ook8
Qhizi32jgHtwYbmruqrSkPbmiatAZlxUJl46TcYHDsvt9UebV90h1sd0myqmCtJ1
lTTbDFg1QjlTkcRkXO/QhLz0FvZA93RVSmftliwT+jA+rQTtR77z+nLxtvMqt25Y
WTZnc5bv2TjRSYMLtaogTE7b7mWQEWX9hwJSwRtlk5Nt458v3xQE8VzeddDYSLPU
jyzbPF8ZOJkINQ+Tp2U1yXzzcfVgMffpwMkFD1wYWrHNW79IQnFaOXyPW0WAXwOL
Mjuut2+2m7lZcBu2EWg8FQ89JtWblu/u7U+cxrn+qQeZHWexMZMu4P6QUmXpw127
LebMrhDR+oDlFBnEd0ezDGdabVm5ozzRDPK+4aRXJSNJmHaeOHiR4r3iQrDh8D2T
uq/ObN2244MyV2rzGx68z6b/YgWZ8sA1VAMGdNLZYJuaWKm6vZRtdRxT/iJVWZFh
bnQbXPlr4f9yRTcj0HqJkdKdZEqxp2N2xalKUTmLFtruPmQST4gHTuGPpevMV6v+
Wv1IF80Wm6vBA4KTwZPDAS0hVZfnuJqeqS0qwwq66A1htdm731Jo3yhiv1nCM/vm
PCSqajYUJiM0UTRzaQngxY7l3KDHk6pRmld/RLm5HN8s1JjNfL6D82Ts5KmZSDbl
bTbX4ItjXJXybWPfw/ILo172W0/GKfBLKwo3Lwrvc0zezsW+W/sMoQAqKj0NkMWe
I6vo2C+pmT40f7JPW9zKNf4ZX+OQsYXNlLuxTMdhBsVosUTQZy0vdwr5MZS7OTDX
/7Ywvz+rFl7YH9xryXKPhAZjZ0Um6ySAKLedbMpT6e3mRsbQQInLfBcv0UwZhA0/
iiT2xdUTL9z7ecUBpVMUryBJW4EDik4ILwZFBLjkIazWa/8r3yVXChn3pqRnq9fu
RGsMR4Ls21CSywymuynSxhBcq2AQxmgaroPKShZqa6NOHQbOMFM5azgLq7bHkt60
/BnyCR1ZDUK6/1+U/68jennwMR5Y09E3v9yEvbL/2WS9u/87SFlgb0J1ChWZSDCd
0/z6HgO2/r+CvGp+wpp9xd/C/7rcwvHQEk44cuzGcNOuxdp6FoLptUxaYE7JpwRZ
XLf0BwKgwKQe/DRHNSfozeaPmmaqbnWHI84kfqROZ3dyqg5zQh8uEAO08i/Ahql+
3zbtZvIY949M7PBMq7gOiYiswL+E3npvETOT+3XTxri11KYYRVi1l+IZ+IfNMeqi
IT0TMh7ueAtT8TW+w3emiG50eNodQ2cmbZk8iW04Ai0MtGew7UkRpQwBjYm8V6h+
XG4yr1e7DP/mQ7s1ZW5o2OUoNZL0EWLywt+SfCl7/cUbqVCZA6jyoq0/EMFPXbzs
E2DqmB3JFa1N2STHbXY4P4/AGaVJ5OC/02lHZzvpBEZ3BZ3WyBziIE5ITPRKn6P3
fEiimB/S4K3XEOLmeTrqSZk+QkhEazH40WcJnchwdD9MojcVW0gb1eB1cU8ZCNcz
4LNmaaCQr3jww2Ixji0FW7+q/xzVJEzCk9xI1oAJ/coUnLURtLlh/0HdDMqO+CaI
ma66ktQYvus7aq8BwsjMbLiGOnQD4Cgg4IX6T6KL373MzgXPd+MpR76tqw2CGrNT
oOU0+jesCfVLzPYoo+G801fN1Iwt2oyqS+bftkEtBxKl7b20xh0JjSDIB9oPRrwD
tfU8nu/aGHUPE/ResBRjc9JfFoMXzesNIMbvTdBYhR0ZXECW0f8QFaNNsFJsof2g
iS/0TGUYLqTNX+6i0hB7ZyxqYJi2TQrazR04vCjW1qLQnhURSKzaNosO1Lwks48t
QNlz66807ZGhJuMxjcthR/Gzt74QKgDY7Ho4KGpK9sOmr+MpsbSrtEIWhOQqzwXH
1P53dhOAUkEQuyBn4SyFDeL1fwCIevNjGqYYm5ckI6iYQxxgGpKok3cBrfOnbItw
Uak4q6RwcLcYdk65z8HrlPuidvjQcOGO85onpoEBeF4L7sDztnee64Eabn9WGJCw
7vuzvazrSz1Klgd8S7T9uRcrnH/6Ax4o/z1s7UUR1peE9JJDH03XTDNR2ErnMT7x
Oe739dhIuP/PNANcDTyqc3q2HKxkgHsEIIIbG4GZ8Xo4BbZ6BN0Nfa1aRi/YDXPL
t2CsXgUzr1Vs1KcuSYE+VoMKpFu9Ryg0Cc/POfNbendiy5Zmw1fzm1P86rOm9siE
o8o2IN92tRbKN34uYWPSYNEo0xr0ipqM/fmIx/DIot32g2hVc2mYFjJqQS1ytjQd
lSKBaxdNsvHR4E2LMspE+layVrJMvzDlb5HqK8Sm6lE8/vQQ6fLbATLQvZwvR9co
Z7XUA3DTCZKZ+WxRnPn3NR5uLLYDAZQK95PSrGTqcw8XgE8Jg1/WQXWvbyB1z+Jf
Vnb/Q+tpsN5HdI7WEAxU2QdvM0+Cvb4xMMR5wnyVQJpax6vd+/fNjxlvCmjJfrMp
13zWwFT7LODC+5AhR5foWPHY84dCe9MRqF7x/VgOiL4/tYiNmEuOB31BofZMsuYY
yE19qjRwroWSD9L7XlAQApL/cawbCtIsy2VuRm6rES29XxC5RQyo4mQofQuf8ULm
jKHAFlOWqm88Iingmy4TJNLpAZO4W23D2LcJK0HRVMb2i9x04Q18snjFiETRQVeH
e7n+sWQo8fi080JPN2Yji2BGmulXOg4pjw3VUqC1NWCONjphAm5JnVYPqOPp+yeN
wNvJwLBQhZ9ke8qnlFJ05mHTiYJCoqgCb2VA5jarAnAYWc/hUyONo/SiPK6VIKCw
GfMtWRJXvPOBUa40g+HlFBtD6Vut9vOBrISd7a/DYmh6Zc0WE6kkzPQzdhRz5JAT
fPSKQJVmsuHxdYOrieVyRHZCkHpoyVRyziHjITraBepDJTMmODy87CYiCFhcplUE
CvRrNYyg58W4zL43zsUISlxpXw7jgsmS2FvI4AFPA73f54XQ6sS5WUUnZX+scg2a
rStGwopkjNhkDeKVWZ6I2QjVNe71l5TOyjCHDkKinNWxq7S8mJ+MzBxJsFxsH03w
Wh8t1vidPn6C/z/7zxlZ8G8kuKdoi6QjViCB9/E2RFtnVPd7w5felghwcIar2Cx9
3QkhZBdm7Z/BKaRz0iHqizFmMhUi76mpGEnOSweKBYmfVX3k9Q/1t1BaiHWCifop
khW+G2DtISDg6CVNPqSyXUd7OVAc9mTAxuHdYVN6pS2Z6oFtC9nVuSxsJJRsK4ze
BK+jv1pahw7NbBM1Cv9cHqNtqwk3dHnceQGUK426X5dT/z5y5ek8P3oHkuiFEwLl
7c+p/P8n0FEKxcIcjjMeFClaaNe/z3Nn78+9kxtTCW3Dq2eHOnRGnqcdBP1qCuBz
g/FNYMoi6ZhH1J1r4EjQCkPFzpAeJMmX8blaRjIvXgH/lk56/BNqRpPlXzHLSsdt
uoqw9jggDKEfSnKcrroMESh0OtaC7aSCNxn/Eq7+M1eH/wAqvqLs8bJlD8/4lUyO
icIjQ1uPOkdKi5xIGDUIdUZxepVcfDbBiQFX/JxOIkDp07Jz1slQhdEHHvfeK7pB
xsEP598xAawnGzIuAQ8keBJRI45C5Ic5rNyE+qvlWGXhAxVxy77odyyzHa5ByIOp
R6fFwgwZJYZ9CwPbkz8lnv03S+4LOFqvoRDPFKbnC66OmkkzNWQL4Fc93dTlmoJz
rwHOuhEe5c4xg4/LqU1Dptfk2vAq+PNAJFawflDyiULQPSiN7F31TVdLEfpSBcfI
8B9JqUCsyJEyL7/tBLlEAl5slXfSbghgZYYNUXwPs+VwGqOHJZsgvzwSfmxONTc7
Ty+lcxKTnGI4iDGVFbJU9opD7hzDKfsc/HkSdIJ/bmX7eStIOUNiZR0GgbPbmwuv
65GM5dZnfZDafYHWQO3IlU8xI8OzPnEvPbLo18mMk4UUFyUata0si9GHDQWJ++Lh
DyX60wDT7xwibiMYWW9M6QktHwPu7OGCwYMcuzy1FhJoKD2MZal7gIZwtUB96sWh
QhSzSD5fS0GZ3RjOcyJ4b2NZv4B7LQ+AGnGSzaBP2egUNSQjQnHu5TNQgWKGoGBW
L6/gNzZEJLaIR0YLPhbQV3co2h54J932CCz1BkmFQuBMR6e2321J1hw/tl6TTO9x
ptqYJmNZjtDG+R+IvGfxfhwj3np8Qg+qmcifoJH1E0Jlh2SDdlI7N+2RRXSkoKw0
pjPIWlpb9wHXZFa40Qjs9uVtisXwF8MjtlQLE42eKqK02b7UxiQoNrdNhVLPkAdh
JCwUXWWUieXRBHYfK0G0sTvreH45S23rorw1wtfHFKz1+ka9yKlrD1l0X1cSuqad
rEwlvU5hlaA4S56k/Y33d83D2tIm4TvYp1efhvAQMhVj5QD4MHAwt6Co/jzlpb9v
YvA/QiIeVjphVSsQkK4tGMUvMI0qmSCGu4YNnWai8AfCQZ5maDN9lxQtMoRBCxbz
f7vNA9uvfPRY0LWc/bJLk2UnO2iLlrO1lvULjo1eJksXvwLTegC83k4wJKMqR1zm
5R32jJvzHbdGh8wmjRGbB+DF7jiBVhSqITLi9J2vqbU4pjjqFIm/nW/xpEDhNwah
ENRQnPviasWJTD9IPhVTPA5Cp+RpxgBoAFbyvTIuV223ON12khbJ/s4y4aqfAUVp
B0sIjthkrNzBQ6pvOOn5EBZXb34g0HRDMrnlOipen40YaivFw7RcnctjC05MlH4P
9LGkSNfwGxcmkfyEfQFRxbAPdNf5eirpy2RjGcrC7OUjFnSQZOdvqR0vH+zvOU0R
egzdmYi6iwgRKfSMVNENAQT1dKbDpNIA/XKHLfJ3Wy5XNIcG20SzD0ieqGCPQtkk
PvL5a9sH8fTtQ0mWJVV1bNqhTNdKRJevYJ8aWL3SIQC9V4XsMLN1C+MY1X6cZ/1g
n+Rs1MJhaDi33aH0OXltgKokztN0D2Ut+kvaZpH0cdlAvMaCe2INxIeTiAec9eFa
+NppJOJwusvK3nUViFKktClEMvHNeGPKCIepVxL0K4AuoUaqGKLNB1aS9Mu8xxEC
Dd2234uRtVvbmVxrEPphr8L8XRAmUgMmEe6U/l/RMXW35LT8s00SHUPS4D3tOYCz
keUJ3tNLC4q/Xkvigm2537yVTtfN3DT0XAtpDk8Y+oXsz7uLBM+zDvpAR9fyFzbr
5vzcFG5+ptrVnHbkVyd0/e4KRar9yZp9oocILwHWPxPKUIlcOFyt9gSf7azWDsNL
lC1aUzIboyZt/nrTb1Y6aCAiDEb3otMYoSLjRcOk355vBo/IfWxQIkFGhYMK1G7y
ApdMc8mi8DFHyMePo8OM3MoNTiSdFhdkj0V8ofTisRymPS/fycExsDwBoMxE8jy6
HD4+HJJbVPUtTPsGWj50SBAxQUr2+D0zWrs9K7OXym2BRHEV8Pqmj8dgILgmAc2p
CNHJsh1eKjrwQBn6NGpbBj9YUXb/lPZDWg7/Ep2X460acGUBAkpz8Rt28EOMiiDJ
hvkEQKX28RITExYRTCPSiAzltT6elf2xRfMU9wcUw3QJ3ZeYjBxjfX4xQ8ZweZcG
CK6081rRNaRLCTFUIWOnrSMAsNYa3bf7prU+YY5oFaN6W4k19vAfzdy452c+tvZO
n/UeFp2JGO1hDdpeJjGU/9rFQDQw/Waq4VQ2mctlCDlyASSnu9/4lcNJukwmjVn6
ktHNYyVJsAUCHejiQfazmcrVSXgBpINS04OszkEFh+VrjY2gjSuMppyocOaW//OX
mJ+z4+PUyI+HeotG+dQjoFPKllIY4okwQhCOrB+qODhDE/dQbzytWf8Zneiix01r
bDD34XgJj2hXCNPH+6eL+Ch73oYwWKDcz46MS0b7cUIHRiPLKdMcRADGOQH3AlKb
Mz42tgJRfCiDiUd85QJ7XOvFlbWRmII8ARMwIi0aLUQiTq5n9LbZemw8Okidp4y+
j1O/uUuO2Td98SVn13WH3S8lTBj8rv1bdhEowF9Pb0VzGXE378PvfzUSMuMdzSBe
UdOjzU66zcx6WWkGl7pNL163n/7jk5v7A06rZyXRswGxQQBSFeWrOlkwXbbGM1pm
fHTY3522pTCyoFUHytYhHI0eWCTpZtSFlMNJuXyxKMXQLLmHAUZISm9JMPUDZWkx
kEtRwznSAOs7XJ4pAdUIN/ow274or/d76D+Pcr/z7UwRqBSB0sPORiZjMZAsW+Ht
fuiq2umIuCPQCcbo1gWR4VlqbhLvhPfrq1YAzZwdabAy8BJ6FlF72xwpqen0Ur3y
4wyELNbowDNAply3GvSWs0FkXzlxpnv5+KeqqSRoIHNsEq0xUgC9XffqhchfLoGw
YRgajEOKQniw/yA+/Q33RUsSJYdms0KFcDstgE0ag5uOAdzp2dtVL0HyZntFm+Ia
arA8BJshCg3WY+f/K2yT4GUVAsy/1Fk409OtGeuNXJ9hhPewa1Cdr19rKyxLSkux
bIXyFoVXFKU6gzWerXblyiZOHH8Tqbq3oTlrexDk3vJKw2IyzfMqACpWwBC+AkOH
S/hnVicgsjPrHgdWLiDD6X022vr1ZyU9St54utMul0UVUPRdK85BEbqG6i5z8d2x
Yt0Yvs11cj2UK2aMqw7CDSQWzyHBCZPaNQ2ClaXRXUHz5aoCgIMN+nA6XrmoYdZU
RO0mczMKUbbYEWG6trLMGwDrv8ON7ENu9HaJliUCfR8N2uURAOzUdFLwterxCuNS
/ERVmVoOX+ANRoU1DmTkL3iJmpnnhe+S9lk6W7QhxNr7Xa04CHHsheC92CFU376x
vgq4nExt1ztAXWP5ecam95XXZ0BybSoVTEXGKDy3o0VBwz/w4YdO2/K4p/aI8feX
XwHZlosVOEvG7bWZB2bdKu1WQeQDjyuqWXoU+FH+lUdCqrv4wHLncVhXCNeQQijY
AodMQS9+RVjwIP1rhnZ90y83KArEHhihBYaRRVNEXfa9sUGyqnNdWmWGrXHdiXEc
nmG1aC7NKsJCAJQjwnPxj2rX3bnX0IsY/r/Xcg/XPY9ZpB0KZ3C2InHZD2IfTb7M
gkGq+IiOTd3CEmwuJC4G/w3NLapNepnydQXhbfrGJfTxwQinEju3cdynXtQUO9Ep
7Yz2W5c/SGfV7nrPuOPT8k5WbhOEKHHfd1js8fBgiObbZAHBU1w+p2Wcy8QxfPnN
F8OshjtmOsFSjUtJ3GFoj+kuQAubAS1+sxtG8Bu6nKnirsiqTDhQW98r8dCjuNWK
KjXwDmDFzhmbxj1RuMzxdN+WuQND2WV54On6CZ9jdXG0iOdUmcxxP1dO5YDaBTmg
te8UAPOTgmSybdpX0JueeKac8a6LDBMMBnWnguSDj3LP3VOcVKddgk++49BTFx3Q
J6faIyoxB2Cpf1iF7LHogGwso8fjqxhZ9LVEKP0SH/biPnygbpFEBbwVN8pbYCHF
iZzD9aO0bfNO4XEghrpO9aiSXpq/NvfTn44FcNLvoSHYah3v0QLpqmbvGohie76l
qyeFJkT+//D73GFt7hSOcMXqQeUylYRqER00qbNifXipLjAv+bB7D9ndpnzFnsgp
6PGLOmVKVtxQYnTjukd4xSK6eIgjDqGx1Ju2r1SbWh+7YWSvKyfdcdFAzlR5qSfl
AlFUGvxDs8i/sP0vfUml2ynPq3BZmG+PA+b3LNlLPX1c+cCkize4FzlnZEJhpeoC
UbeHDKWcEtKIR1uxbNBdYjjJZNu8Spb9sVNV4ZA+sFMrCuRTZWt8/H7FK06HygDf
TA6g6UCA+6Z5wqfr77u4AX4Lptvkub8B2tKUVHdR1jX5h/MSgoasBzsLGkUm1hrr
6wY7wiTGnaOs8mUvBPI0VjhHnHdmVwvs9UiEl5BlxLfzCxt/DzSv8GLnrdJ4B6H7
iUch624UxXp4kW87QcbYRy+oAO0bk3Fg2zzlEB/1sm5Hrldkek2Tcwiu2+wysFDO
z50XFQtS6ztkdzbJVHYqRUPZupuU0HzpBK2LaYCoErcreBlF7XG8IkehTe9ggPx/
9dDtfwbxYGAAPxISI+vOoPbUMkAH54t0QqupVSNmXVNyy0S+UYU97fU75BZP1Fcf
cKbFxFFfqFnIxZI+V75ls8tPcvhYXXIebVuxaKNqa2JmVjxixrnd/YPdtB69Kb22
lzEJDQ0ym0J5DE2BRmNc1rKZ6XkuERiHmXOQiZXcrBR5KRyplSDQHnu64T7VSjsG
pOUJgpwz1ZKexFyYhDJwcMH87uAUpT9UwgIWNF2GHYbwh43GG19+DYLc7yfMQgJ3
wbXL0l5YE5KZlC6FJ3B1FZ0X657AALONpYO7fpbUNtUay8aGSBr3gWieABsdc21c
7TI6PkCp/uAb6k5EtFNMGPZrUrbsdWt7f4g5owztDZEFgl51tYAR2V4AqMZ5tGJP
14u99MOT0PRqsPO6r1ffjjlQte74S3vfQrY1B2QE6TlLXzrMTk4nP0cC+lc/ONEp
W9ZRkt9eNOxHelXFFq03UO56bwEL6Gnh0VsS/DZJkgEhfxZmx4of2WCVZ9m+GMrI
GylMKPXOqcJrPK+l5bLroXQsdxPp7v/7eQzqQtjGyktY8VoriPbMRw6rF4wCEvwU
hnXddIHIM3NebTYlWQ1jdcyLWXkGx5BEDGl+Mj1PgUsJHNSUt9jNNWpBsGjbuund
p8k5xxpCvdxI5LwVndF0hey9jKQXH072dz3NwvztY27qkkveeCYGt8Un9rtl0fSy
UMWurr5rCiv4D0s2B0xE4nL0zJ5iDsxqeVlpSaLRbRCXFoUkZU4jdl6+gsrNlYeC
Z0f4z+VXMTt5iSxzh85MFyhDBwYEc+Mj/0CI9YZG2OHy4/tR+XoGCKOW7Aw4N7lO
UojJNBrt1U55C3bUGH2a/YbufM2nSOGWP8voM7wGC9mZm1Q/epUeH+XNwAeCWfwr
KcDctQ+WWd0nbb94NZFKHGB+Kl2PxYXMo2Hr+LLcM6iNmBTh48UdOHAQrW4+4UmP
anUccqke+nUX42qvfOjOnkQRK4qTMyrgO/IhLl0puIPbUFfSwjo+bHcO5qCOZPDn
dy2M7jOmEmwoxs/Fv5zk6OLRjfTQ5nfjzSf984yy0NWsaHpRhpoYtRxQ8f9+LVfV
j4k53+nkYr1qjBfKVltwMHxmGW3WlAetYped/kXTGtqYZuK8EisPbcfo09gh8rTJ
nLg7ygXJlk6YXQ+iGt6+ZkiWPjwM2Tb8XoZu5DSqS3SK2aHp4LuSJv88f0kNjpc9
s7P9pT6aO73mUGvDdD3i+rddtmEBUH8N/J/KXD4oi0CgP0d7UthMo4wQctJWBaiV
ad1xJ0HupJCuESgQEQ2DgoxcyZK3jGweKyIYrghy7c672G4MojM9ysEhijBJoLed
FVuPUFDDSDqsWyrvR7lZNUC5nr77jGQ7wFFOXqp4z/f/pr9RiPL2FSqI6vwQL+mQ
8fMzVM2w2RpODe5RxnhGehtdprXIkGLBK/FtuadwcvgmmfoJDy0RQr2eMMPxq8mR
+VFNbmHvipQnj+FrnI7WH5xyBh7ReKu6T4ZUxgRelUvXNpb7mYC/Wr/jx30YG+pu
/nCr/ol/wW2Xs+MJWJZ15czPpwWGAJTR2vRVHhDEMPtfc8P5A3MEKLjM+QyEOqM4
sA2EsQNLcUNpBki9Pap8uabPY6KQjwpAdNomq45CgiTr5h3mUhj3l4pxPTXwZIXa
CCFELrjofyaL0fx8a5pxq46SW6uT/KmrbDpn5zNMsNY1wAGJgp2g97NRLm6+Cw7m
hmrnS28NhS9/E4lNcyDfs0Gd4VxtbA1CFc5Ck5k9kEUA6GhyyAQC74RxnpzLLaeL
V9nb0qZRj0M2UJ5k8gKpjg+gX39kw5pml3K6S09Cgb9zO75H2fad/XIch2bLBzns
760vUw8v9Af4MUEp8YiEEIp1V5c65mvX1EbNqSgpw3XSok4XENlSaUnBtWnzZEjw
2j2BDMn3oXX4r+WS5cSek4eoy63G8MnyW60DJ8I+lchWutvS8ejnhdb8fWjmcANz
5DAkIOXsBIpo86DjcSzlKYKUwgyMQu8JAxVVzJGzx+7XM/jzuKxUBtPtzR160HeL
kiNrO+cFyTyMTFtZgDPQNP0DMgOgrZmFbQdsMT543h4LDvV55eLYgv80RnUxYq87
tcVMNwMfWMcqTDjuxanM7qqxYb9pNzhsjg9z/2pjiJ7Hg0w72NLh6aHCxRwMwOOO
TJRMY/catFoVa5xv+bIZc8SPCfxaEkUWomKVjQ7Ov81vZoutvs1RIZvSk+s33kte
396yylEZUiGmiGItILDPQN4G1P+S3F5TeoUxbttajCLsMiCGlrp0/XMVz9zJMNCR
/Kjz4a/LYaWKXAD0RlMbRLXY2fl7HMQIBEva6LcplvRDt6JVkVqh0Bes+i5SASVe
GbaprI+zY+rWr3wLr/sOMXcRrLuXiZLRx//5a6a9jgSAlqF9aB/VLcGRm/adIlJ+
ZKGRFZPNTcuxo+QFGynP0LbqKtZBpz3N7zH+72W7HltsagvcbeJlJcIRzVPUgCga
YrOPUZovagHIYGU7IZRVK1rpEQjRJrou+W5rMsquWfXEqXEg6OWXG5tM7iaXIMU/
Lqqt0Rtmnrxi6jscB4yy3qwtwwnnhhSfGlk4KVb8sN5DFl3TqGUcARkKF4NCf9qC
2/j7RI+flovFz47V/CUdYcFYEXe/3Z6XQvFHSeoaoRfqSYUUdd3HUl7eMnNUrjkO
iquEmAq8aweUVyoioI259bwzTU+76HUEi8Lvgusfn8uQoQ6x80gQEj23KU+ld6Kj
uDBD/rDWVNZLQqT3XhLEH9BRRU73410ic4PeFWtqk015riVXQ06R4SpMRRugkz0r
VB6PYnfpzaByrWTuenbU6PR3trGWY3yX5PWRPjTf915v3wrEXNOV3mo2H0hAxugO
VDKJgRIgbcI8GahIcHEXhF5zl2i1ywOyDuLIXwW9S/6M6Qx+XJRwg15AIEpFYh7B
B9r0CmJqrYAA+EBywhRGlrk3EeyxIY9bJ5DD2js1DETCzObvSqpc1wBr1/a6bobN
MDLx2xBZ2W3ChkAnB5PLg81KEnEBWBQKq4mAKCeB0HpWGNKuu4a3+Aap8RESr4qS
QVesIfbu8QAXYOx311waXlLhToREVKHjrbi9A0Q+KqURoSImmSjTnGeml7nF5vHA
rKFl65iTU91orUJVzumZsO6wqeHCfY4BYsWjJ8rx3OdDYJoD4O+pi7VFc4awX1eH
MgpQIqHMxLSYAIZo0CIQ4EnqGo/xkkusu6fXT9h2J6j70YW9qGDpOm3tbOuguVF3
wWrlRRVksD/7HmOamZ3VlrH5UhXO29e7jpUBdzNnLGbz4RtkeMxlTYnypCKbh17C
TBx10v7o88CrEMAlHShcq92GBTZZVS7iYOdjQWP5Wx6DYu0ITU9U24ECkvLBwOVJ
uM2hVBou3SXEij2T41XhGzfCwizRD2GN+gkuGBkdNDwwGjtqLjIslawLOVK1HgoZ
be9Xeg3mhgspK+B6wcYKBuad7Oq+02FQZXpOqPxcURyJRlqZ44GVBkJWe0saWJwI
b4CAVoGKZPb98JEph0SIdoJ93+nucQ5fCY1/3/XvM5lUNeCNNIiYAtpF95AWKFNT
pm5ATJEBaRZ5xzDq9Wf0mEvfvzWRH1wVXjsPfAoKSUbrxlzkA1xfzH+abv3iQnmo
ZqXDA12F8zTQBcFsFZX21M4UfOSIgyfbW2SUrbVsax8pxlcLBJ1YRAATfuQGMb1z
vsHbvGQ2eElmBco/RXbY74Hr2vccUxh029qqe/8RhEJgB+01rJZp6UC794fHiRQl
6dBR9UDkaqPWtPnoBRmLKt4w+BOVFunUXL/oC16/J5E1lu6s6UJuWdLXXZSTsUAs
fM295Fd5H9XQM/Ab0rvntocMD1iEH2yyZKbQ0SErnyeS4bQ8neLWyOo0+oeesQfp
mXRyzbvIavp/4uPGq9lEYNIq52irlpH783Bc2B0Ibef1wEFN7TdJha3FMSIH8GT3
5MNzu4E0Jx4acWNvj7RG6Vjs/AHyqZHiJhf7K6+RGNYTY/Xb0mNvHTzOu2mWFjuI
8uyZ58O9/coilfoZNBNUjOL4r+5SdIP67uXFcf7Z74BcMWmog7yzbm+qzlG/X/ZZ
MM0te8pvAUzH24D+A8+5RK1+UNS4MonURfCP9Xi5XcddxBri5eioI5P7xM07Vn/3
BHI4UQ2026oGMdTF8qiNuhfgccTY3nscjX4U7CGL6Q+KeI4IW3wo+L1HndTiuLYE
Hdm4Z2HEVNBSMxvc7tk3llS9ycX6kNM+YUHKhQ4W999lEDq7CYsb6Rv4uXp1a++/
qHvRYQ9hfoIEgOOehvlmhz9YTRlRGF1G0aVc19pW+9lKd3F5GLuBcHWxoJW2KGuo
wwLu7NBoFUEDcV162tQQrpAKLhL7firAhrwQQPdP2oAKE6rwS7uW7s4IhnEAqsS+
1PgOvzUYXo8ZVWjGMO+/MxUul0UUB6+M0L8M7K0dAbRxxYGVGrIYqAJctf06YvVn
XHs/gLYpWi1dWe7H82ef9zJJPiC9LTTf7APBJpd06rboF0AmwXUDrBoYM7u6owXp
KKCC4/sALjmzUO0M2+IJmeRc0xbsNxjjRV1lI0JE32/UUdzZ33S8pBqeKMdEQY2p
Eoug8t5fiaZFMqEtuGuOhO2/OY4zm08/Np5mdOBw3vuUBRHes9hOWZFQxD83TJjT
hkioYV3WwKfqtPydUnBOSa/YsDh2xDW8A5MO3Cw4BVPS92PhTqFB2E5LfXFHSDvD
dVtWva+Uu9B+w4wevmLeehzT5rkMzwcbC7Ewlu6eF0hMSkfDKq2jyNA6Mru7oHL/
AXrfS5bpc29F9Z/dKXaIyq5hkm0xFw9rvd81y07tpVvPaCa4VICSHPLrEI7VhNAu
/E6d50Tbzq+AVV/kW2XiYzCajVyIPv9qVQ5NEVBSsq7baTgGWWUV9sFPAJwItfkT
ghdkpYwVgBvucMCmVFZ3zqKwd0k5Y/rRHmETOq6+xRoMghdvwXc2pRRQN4CT9BLR
PJXuVIZYf/qI+PFpxFuyxvXgKx17tjFDyi6zMFnfA/1iBuMu4/jl3d1LexbAkYJ8
UFgr/bH7Qm4n8vvcCyUmBOIIgzCuxHi9jB9XzEpC5rxAmuX9IxaF/QYjQZdwqe8h
NZf3RSMX7/qRPtTFUMpj3ccXFw0Oo/ARbxtA919itJpUplMPG/0cFll/iLS8zaX8
zg7FJZlR8xKVyl3ny7FssXo19LYU35mug1aNjLSMPS/yboLv9zljNNah6f1qEzmL
TeKP8xfQJP+oSFLzE1xzRc4dIMR+WB9bHPLLKZuKPE72ffaoqtXw9DuE6FmEhiqY
cc6bruFY3W1MIGVjbvvYascg74mvaEfQdsmuV5MGi3D5hafggWw8+GvkVOzdlfFJ
N12BfUnR+X9bhUyJpmSriWmtkkPT7KnQVjGfBm+5EmDpvAzsJVK2jrKlJAhb87YQ
2EPrqhguHEul3SRszxTZcyss/hYDbXY3s7YUY4wHLTYDecHW+1s/DWj1w2g1kaai
f1/W7m5POLWvvcftolFLUHyqFPFkORa9byBps7HS1T7NGFLW20qOVhF+sPh5PGQs
qgTIiumq2ibFW3btA0/U0AOevWSR4lvJxFYGkH3WRtpqQvmSB/+d78EVX0uIVhRv
n9i9C/hbiX9zIQ3hjXTgE+TGCFXzB4GBn+lJnUVMeQXYNDvL/KoxEVAz5BehKSIc
F+XSi4rzLGAX12K5hSkDnYD1Hpp6ZMmS/SDwqU0pKtDI3lgJcPqIpO0yMC70AgVp
v29OKfgtbtoECJFFTA9DYj81nz0MnQIWVJp+sSFPjUww3B0U2D1atNz9Y5SvgQl9
D3WSvbm0lqEi1K+iafFFHYoEkqTH6FEBkrzzayz+576wHEinxkMclqck9ukqGY8M
kLlG+aMgN407DTDawrQLCRbyhFjq/SgXbsjjRoGot++uA7Z+wnryLr9cR/eg/nlu
8l/EwdYkdv736xR+NDfAcbmKnsLb0UdjivZ8rwMmGzUg6tLPSeQlNjGmmPmjQHJF
mS2A9FPeenvp6BYSt7p1OyRu5HAzrcaSIjG9rjjf0G4UZpsdjrYfZX4Ou68HjGqE
bKI2QAnup2VxO04BBQR8NtazH3vEjVN4QDDXWM01yyseOLPXjVdFOvvSYLO5Zi9E
krQV6ujWnarT/sBJd3Y/QHzIFxLcB+3zIbvXKDeCXdK0+UI7vNo6poyvRPHS0eIM
jtKECBoAoeG2TNdidRTD+f2H78qLvmrUlD+FFeQDrcDvyHuVCHB9ZedOGmDZt3L3
LMQnG+J8vNNOkK+iBNKiPPrlpWLB43ZJTHtawL5Az99clMKtRieEh7kn3sAhsddl
K1r1xVF476/TwwGFdH0qSlfIIrtCM1dvW00ql9LD0QiaidlUd+a50iXvdku/CRf5
+0Ub0r6XkLt6qfHxQQrjnUijTPo68YbDhzCHGO7BOXt5Pn7hX47t7sGxTNSrmNI8
16aLiKW3FJ3MPy4Xro4EtjRt7c2m5NJi7yq89Owuir05nyyu68A2w6P6W+ESnfuy
cKc2GcdswP2BwJ7CxDxQALg1nmzB/i+9BQJ1vLDqa2GS+M+/jZKMLnfkW3ikCg3r
LT9T+jvioijMfQOoMnt3L77h8X0G21I3PopcCziTan7ANV2w/YMfN2eJmmGqXPtO
0Eges17W+40ZZkIleC5ZLRwinQe/q+8c8gWpmesL3imdo4S8Y02i6Lc8VwQmbmEw
zXueSWaz470510aGA977sLa3Po0CDuJXMfxgULW5vSJPDSRO2KgQwOJRaRT9lfaj
jU1+YzjQhusU8wIY8rcK7S+0Ql6DBDEdN6TslFXbydFOMr8lDTBFF7yRRxwm5iLv
JN31ZGdDlwuL3o4eiZviRRn7OnVWz7KGr+5NDIe1PMQq8SOWMDuQQrwCasR4nVPp
7GXvj996fhD10F2TPbcD/ldvFofc/w4J6eWbfTtVrQ10eHhNf9j//q5tHbnh1BpY
81zolLzQyisX19Y42Qn2fIeOVpvsEzq/Cdxv5F/+Rdha/PI3AHMQ0KOthuEj7EJV
Tsw7GKovgDy1D4aZjhSOyMtQ4hESdDbmBL9MtYacI9aolVwskqnzGDLJxIfAbfIT
KW/fT8yPl2F+uHksVXa0ugF+GJBNIW3ykREra18wgzTqL28nRi28kCWnIF6IWhO6
yGUkOdrHt4/KO4PK/KNDz7E4fi6fTJMRtQvwn1Z98BenTNc+pLczeoorJ3j2+bj7
CeAayvGva43IdXIKaWBMfaoNWCQMn3mobWJWTWgkDO7heXEv9g/p1JZTGSMHwPc+
WfAvaZ6wGVEYtmJtLpakkO2APms9OjPyqLfj0UWCAgN/4oQaVAFL2n7PgwxMLZBC
VWoOyskz8WqSLuvIkdhAJqlKzwuo9LVPu5CNDdhG+S0mXhAw2HxZzMIH59hL1V5I
xUSsgeaYOLkv552pgDLqAjGm5ofavXoEt7S0soO8uw8TZRrwtz2dwuAGd0dpR4kw
cWbAYKn1CFegFFFsliJ6feojEjaUbi7lAF+8lFFhQe2qrpucpp9LbDzHKSCQoTeV
aBScc3XM2EVGaWibsJvDhXWWz+Tys+XjrG8I1wqkrJDSPyfGwUYnAPnrIJXyBJej
ZvWKyCNRmj6B6uzMKugXl5J2xp0YE3KFq8EsoXJEXeLez4fN2wutT+EdJ7f3tdQg
kBkKQJoUZgOr5r3uFs/cOug2Hyy6Hd/ezUWV9loAugfkNGVnq5an2OyLFM54pNZG
rfl90rMSBJ93CAcAkexwQxw263QVr9tWBc3JAi/XVDGP10eimADPxE4rhyHZda1G
7hzZwI0vOTWit6rrCSpABxlRQEc2sjzzislNzVlDPw2O//di6nm0nGSHGJf5XRHH
iweHfK21NWSv2Wx/pFirLx9ykG4G2+OGi8nh4xiItx9gjG5Fh4rGTS7f+Tccq0Kd
AYXp71hzucSujMFz/FFOi5GNjBDJ5yuXskFqKcUAePi7VUBJJRCOFWCshC2c0Bf6
+oNXnmYfNKr1QCmVmcXzFtalp3N2P34y8ByfcDTOx/WorOvOwxMDl/3mAyGVRWfm
KDXrysOvc27uymuDyq64OermN0PT736zL8r5eyiA/i1DM+pZL73jwf8h+7LyNYXW
AKQ23RABb4dthcZ2mjvoSBqgPLYzDYRIagZZs8E2J3sT/b1Sw+T3JfyUgsqx6p7H
9qviEsp/d+ntIEFyGi0rdr/4SKL7lByScWkgGo6jg76OPAhVrKi1UjVfeSpnq3Pn
8DyOdwRl2NshUWBgIEZegkUtug+LHwVdamqKJ6XWavaj1fR5D54JNWJwnjiyCu51
qp8sqAx25pCR0RC/K5R6eJVbl2b5odkyXBU3X5Fe2QN65AXrhbPMYMUqHDU8BAUS
dv8Fx9nZM3gP4XitA4mdWCHsnnpuqZ04lDWnNRO9g9P968dEhtMtfZRRLq8F4SCN
AgFGw4wAw4BQM2WFCaLaZQ91syDDxzRG3hbz5MaY4ooja6H/7xeuQq4RQ0RGJ4eE
8BYqDoKtWBxKE+rpc3/UbUo2f22DGlPbOnsUKs0mg4DA+cjTbxwwPoLcoFWVqAfS
pMofiWhX++7Zzwz+FuknBl6wNgP71hPs2whOcsG4LcB4A7/nbeekksl+DLPhl8r1
AIMpvlCmxoFdRFUuGw3Hw6H73NAHDkyS0oA9umlReXgPT/7572j2HKPWTmtTZsEP
rScwvbRzuHekFYbnfaQn5uEWlam1wk8jo12MHycL+SN6eoFnbGDlkgI7r1oxEIdE
3TdOnaozJR+K2Rn/TXodmVFvdylFj5FhbLupgZFnt61UJ8Sw0yiqb5E1FcDad6Zk
weKMjKU7Q/N8EqNbjqqHoM1DiZbXmlQ+ZUMWN3J1NxVOFuMkAb146Hfmafajq2LE
GlkpHId5t3rcTCkWXXn1xztW5vmmmkz7d3LkK+7XV35hvHhh6rpjp7Xr3vwHes3l
aOMEtQcrUvdmL78HwI9hnHzZSH6Z/+EioImQLkyrxqrlnd3Go7gphnojk3RT2WI+
V/8pTlOgPbsHIrfZ7v5FT+zKUeUqs6zSmrMBVfkFk9mZIVxhYvoEJlQALJ2ZGtk8
um0uOYmffFEf009hleiZV1a2FzEX78t28YM3bOCcgpO34wFt9S01FYT2Tu6RNqtP
rHwZbxHesux26vuHcY1gvcqhI4CFD7Lz5/wN9mwWF+XfzrT/rdzATyVjx7I883uf
M8izeXtBqbd0ettnML90ffUBzmf/UTi3fT5dR5v06N/tecZQeSa48cJPDR9rKr/g
jt2atxcNBdR/7UMkFloqxvW/XczxGiA5Z9CRrb1Pcx4/NMsxH5FYy0V2GrOHwtOj
IP7Hy+s090hsVqNDDn0xhA09RzDaucm322EBZKxIxgf811Y2nDOrCno9kdtuklDs
fpnay33+Ib8Jz5XmJdZlAcJNI9u6ymV+AxvUpoGDt98urAIspAadzKGwhlFCDisz
Q1q9hz/Iw96gbc1w8U3ezIuReERbWOEhbOeUQC5eusxGf0Fz8DeRrngz/S9XHMsu
8byOF4drHxXQZMpyAp3Aj2gTKfVop0WWf/EvXBcDXpYg8uWKzQOXl+LahtLekQnA
Zgu75e+ASrDRAHM5EwOyzb5XBDQvrcOOvkrpQBe0ggqL9lSp0QgKn1c9/5PQKVgf
csNLfI5L2M2wNgJhFKJT++I1F7UVvhHb58ZvxHSfraAnIpAS8Ur216zA3byXq3v+
UtJNDZ0ygttWl117g2CtqChmCL7fgmPIr0gN9ciiJj3L92vaUwcrdt1q9S8uAIEt
HZewUJFW3h+Dg+0VCyP4fM+DumuVcGrjzwCa6VQCz5QkcJoNvwCUPhXnVaToKJBT
07R/txDb5AL34+QdOIMKwk367IwwgUzJlza0ye05+JO5kxW5CYxe1Kfj9HcI4UrX
bD5CeKPTv5h6gyQutUElwfdSqnjfHUyESM12uTPVgf6a3HEaYB3O2vmRqh7sx2hH
mQsbQAZhWSdevl/N1/GiJ44KGothPknL5o3AJzgwdpjHmNehHRc5JjytKMP2ElZL
7iUDryo5szW69ketND6KxCNo4ETgyucZW49z/NZTF058ZgzgTo70IXq8Y08CqVbO
IRJvH8uueQiVNwAfYF+ZUCU4y5ydVdIwfAUPOaa7HO6sEUS3gcZ9k/8FI1pvUEHo
Zht/hDMT9SWmGLTYtEYx+3Kyt5i4V0BvDZTT2FsVmQrpvb5QCW95yceYlYPS7lwf
YMHMoupjflrmxHKcgBCFCtb0loQJz4b2w+pPHguHNkSP6lRWedvosJaYN+b0gbtJ
PlN1+UYscwncbq7Gpr6PFzYyBOiMMm/zNyrcL44FwAhg9WEgMjfiJ13sebPxdzpd
WMqYeyfd11azJl0AjngjaIP8wycWy9NQtAKM65EmbYZVjC9G2bvAzguF51SJmlvx
v8g5b2qRe9vIbdZMf87xubmaHG5PW/aGVGMvKYxxVlHR617Vj5BmBE0LGgg8hHqV
0OwGYdLZkGT/SXJOf6qL3VtGvcawzUwu4jAF3LTxXFqeAt8IxvSdoMtQEYtDwm3l
DnOwX7ae+IkZbnQSg2qELUFcPIELUVfirc3O2oLGRuspjb51QBHll3mIZzgr5OAw
C6h/cSf1r4l0tNCKHWc6ypdknMOERAluVszniRNugRbKrPjk1kmES/TssXGbQFvr
h9/5HTAUpCmYUSZ6K4ZhT83MaWcKAiGOYj2nwdZCUelqvv48BKCQlr5L148zyKCK
xdnbNzOyoAFVezshlVxN65VbuLnrYenXyZ4TnGywwg7btRQe5z2FxofAlz2yRq23
dzu5JM1ioETN8eZyO6+heJdfKoYTaDZhcJpi73FfpOX2E235dRPwAcP7PvT2ycBx
xXOf1Jyq7bABoQEe70TI5y4qCjn+X0q1GN/Sl7iDeDJTO876hEbeZzOplaH1Z9sN
XQj6l/qw9cD3j+fE6bFqDYt5yFGSM0hVUBXRkv7ntbGlxgHXceHa3s4E4I1W0R49
mnsebWTWAvunOCU4slhgy3tXNODhvp+gaH8573+7CesglH/JrCzBUZd+DxCoSe0z
yROnXjXmSdwl5/Fx8+QnSJOB2lKXE9QMlwFQqALAJCSz5SmZMaTp2Cl/aXXI3fjj
yXl/d6g3CEJdELsnDv8Q1iIyPFdMxrEy1MwEqiRNpPiZ9r2N/szTQJ5SM2++DBUK
T6jxRllYf029V2hdP5h7UaLUcs5vkf5F3E0EHN5AhHNZlgAw7xF7L8Gv6YQLPzMJ
Mw8mOJLxQxt7MXF7+iyaNkR/M1LxSu9UuM0IViODv1NjCVEiZMjFyU6hUo8eNwUo
cQieLilLpVwFgENyRzc8UVqm3ajQfTqziHcHKMdy98xgx2Ja4sfPV8k6s3ETtgMZ
usdEh31ZJ3aQhZcfA/hXPdCe00VLN4F7p3YIusDmcFsMLISiH6SC4QmDBmtRS1uA
x46mQ14H0DgLhrtYpsVv/9+RWQUQarMLJDR8DIAG/uXdEAKVjjV+L418BWOeHDUS
y2+7m3HF9PZNsovKctue9MZcOIsvNrLlbaGT33ykHXVJwzHpc7pxuiMEBHg1aSAP
PbrsSBuAtbkH9Rjw4xcnc3xH7hpLkwPAw+CEHNGNyDPajqhsAQ2yz5UJjsSagN+j
LUGlUmQZYoWoSzP+vnQMq+NDE5ZCEl6ve3iDo5/7PzuiYTiyqbEhJia6zwSpwhy2
uGHPUAM3WH7xNIFgzLgJG5y5YkK10WK34MPGG0hzxJxTYS2C3MiELsrhV2cRqRiZ
TXGyaDVE1u+RWoe2SDBA8vsOsfUEGT2+VVHeFLJ98bVdRS+EwTiW1eE6L+naPgIz
kRqy1ExjROdKyfZlQXqVaGn3ZLrieuRsvtPw91V3gGLcvUT/IHI7d8oFGkVZOFZ1
CwjqY8vnTgRNbqfxIw8pk4o7Xx3jNsRU45ke6MaXAXUfEl96irRgf77PsG3Qyxpk
Rz/43tx6F68IsVYdiA/fWR7YSABesgP2DoR4MqZTiMDAtYoP/PsrpA++s1DpqbT2
0oNA0yO200Ay5nzvORWaZDIWzyKilG72dP/e+ighpKats0iN//9kgWYLeYfMoYjC
eVvbPlNR6i1kZDxjUSKWPxQ+9VStA/hMfMvtKaemIZUYX74Cj5s917VNQkgMxcvL
/XxdFMPJRh3F5avf/8Cidm60X0zkLg8OJxghY3x4IIj3MU1bktWdOUDFa0lB3x1o
+fFG6eGmqNRA7Btb2BXwNTXuwX5Zvb1WhLQhCVmyuCW57Ui8xYuRxAoa0DZ3TffE
/VrCdG1DxZ/NMsRjboxSH0KpVne/qjlmy0bVYlQD7dMIfrTAP0ip53f6/DM51OkQ
wPfC3ERi5HYnT7xEBckLnp9e4t1ehb6BU39bRdLnSC4tRr881Pvhg+aY9M+pZ+V/
s7UshVP3wtA1+VLKTq52gcw675bFgy+GSis7or7aexHHwcPuBmLJ9J/Q911M9+kM
814oBfZ0xELZvN/HCR1sw+IXcdfauGCaolIwbLfsIJ2h4PSnd/eI4clZ+t3ta1oo
l2BwEse9flm3IPWD9Ys1hU1wkWzy87DozAbygN35IPfa8TwuxaY5U+x7LoNkmzbK
0IohCU5Pnx5IG6gjUXj5/s3wKfbS0A1x9ardQr6psHwqI3QmHoHLtptIFKaBWBnx
hDBtI81viWSvcPAu3cdflgu56v4zLfgsPlR4euvulF/5SnOlngc67ahpwA9pbP/P
CedU088TaXkxebPk4E7PD55q7hvjO6532INlzu2chM5S2Jvhm36k0s3fhvRgdjYh
zTHig/nzTJIwu1IygfEQ3HclckR6XyntKT1knW8SzME3cnE3s/hL1ThKZZNT3MTf
NY/6vj6pNcWwvBMM/79eXlrPpJSAtEplZEuM+pxJG4i+xtJ13MndKocb5yN11emL
tMiOc7WJY8MoJ+MVF7VkN2qIMysrXXRxyAzc8QwfSg8fqNfN+AtiBB0QHX0QQmDV
wlwfVTMIoSdWTu7yqqaboSjafRNL5FGRii7X/+k/Dcfehw8Chp9XcBP44UGb18Sp
Ycjw0B+35MeH7i5M8cZPnYbFqdHeecHGYIj1iTT1HtwMGx6wi8dO6hYoYIVRQpKM
cBaLprbgCLdnEg6OPXy8EuD8Y/Q6/DwCcnHQUrC/tnx9oP/dcjVUjGWTV1oJtuAK
iF4vEtsOxBUcExEaZguDQBVO2lhPn8JCmoHmQ6kXq4gAOIAFkM4ehoqaZ1xrjGgM
q6l+6qMoK7GruBdeHH8MLnf86I6Pmb3sLlX4gGl5zX1vS7u1nIaFotADEEvzzR56
z5IpPuhnbZojxUeJP3Es6Q101TMdDetiLOXee0l741V7UWbqPAKy7EsieZLeWhSZ
81ZiIA+iwH20Gclqw4cAoGelLGKywpXoF13JCgrPGFbOmgdAJwJrG4w+KOQ2Srm4
raAM8wSlF7Ge/8MHdhH2b3+4pj0kP8MS7nGC9xMxMqnvKxqy+0+DmpeNrMHcCOPj
QG26E5Iun5AhcD3JabNNxUJwKJEzyzxSQ9rN0YdPYwm4Zu86smrr4htlCnQWVNGX
FYVNXCrtHDc9LbBxYTpbCXMiAJecUVb84BZFdsTKckxVOfc1QgA4RWEOiUExF8X0
jLlEctP0K194xzOZlEFqb5FxHI8QqI6zxCi3L5m88bO1eFHgcsqtMVJ7VDYHX57P
juO4cJiKSYdvnRHholjw33MFYhBoeY8rfOiL0eK5YSQUDLY0quRroKSExaxicHdK
yo0U1nr58lK0hTy5P/U/EjVkuF/vvbpD76jG5G4bpwXxles/TlwmLLWVrlmEP5Da
Ze/fZi86ktv/QexLbOUs9BpZf3h4J4MBr4bTgN1ytNIpFwJYupTbLjHqvgTM65f5
cEqbIblr2cDZA9NtQraZRHP7g6NcjBfu5em4OZFXvGar73k29w8+/DSdhEN3NvDF
xvqtZCqsAZKo94kHKSCdr581kIfdkm9RwufzydOXp6L5yjTEaTC8WeStCjTnPo7m
c1/AwtEij5Ohgi+rEKmy7vUNlvxO2BzUp6ZbiNiTvvy3JuE7Ob7o3hUrL0ETfU4+
NcQ8hIk0kuPi95eRoOzZGfjHSSN3YR5Z0+TUzm7SoACQaZC9UQ6GeqD92UG/1pQq
dqs7zzstMjbWjAEYhprsErCT0/RCx+1sLIpoq+lcGAuIbNMRx9LHuQWlcvBL9ivU
JA05IWKFZN1ZGTUdhfQJTmYhw6v+u76xtdj7TkeidjMc/hANWdHAR9sosgIHN61R
jPva5dywMJ2QKVesl4dbBDJDZS7vmG+skTkMT+UYb5o6POW9SRROarKZpl9pGWvY
foVxw7bIh26Xm89tnyzEtLx/4lCuj7D3EhOrmwpGNZEUIUEaBRTC+gSecHdeT31w
/QeaNDItlwAAHseQiNxjxsJS6//VI5/uQSaKko/XsQRWTk5s3wEoVVgV5EWLZ1pW
kLMweFT3cg6heLsQvkM5i54gWdm1QUIbW/3hPaMCIfZdxnbXEr0z0lGp5aKLDBlF
hpSkx7GaVN1MRhsawJsuN3LM+lqxaZY7wRS5vDNw1l2Lgfc2Mb6lDlJpe9dOY8gt
HwLYUDUFA8ayA/4mMEXT1mKr8uwD2p7mwLaM44EIjRI40f41WjCdmePtsOZW+x/X
Kx2kGCJQlH50GVS1nxXwftZUPu12krRFdRuHkGfVENqyTPfinIbbN7r3FgKJwgI0
gCzqPipY53t8KL5gRjAv9C8fngk53QPnAq0ew0AKIsr1llFzLssdhxx5LskktXf1
xMumtZcPWNEusjiSFqpZMzIW+TQYV7W5Xc535l/bP/6aApMpB5lkOej88VywTnDU
S07nMoXJfAGdHTuG0HvdrdnjJ4IV9qC1MBcowfpAgV62KXSqKn8shjRpNRvXVrsC
Lp202heNVgyMR4iyt6B/zHYz1Axm464xStn9NPxI6ohqNQDr635x+4f3YIe4hmrs
SQw5ABgcHQb88mTF7mPM6pf+K0JEXfrLTZuQM/bsl1pPrx9zpeubUChc9IgqHCHb
CG20HdjIhiKSgqNwQKbBSPnPHrg+89zrmWPHwyvqGPhCfGVHdl8n80APDqnekqOU
ACiBi5OJbeUKpv3adifsZGhpMKpNFijZtwJDRPxAmnzGrHBK1BYhn7lJRU8lqDhg
wE46/rx6UL4dUSMZJVGsDJ+zSqcmbROf+XOHZWS9O3o5MphL9OgPYoEL8gZANGqC
EhDdQVyOF89I3EHeGBin6chJ8zxzId9PWeabkJVM+Cp2vAsxGp8Ln6CDSe0HOePz
+5MOWu0KfoP5rrXL/rVxWBU0O0iNXAf9zGPoHOyMFeYAeiwUN6S+66oOZAqfnZDz
62c+zypjDp3YRe8gQdSZ2zfQEiSY+rQeXWRZs9dfG8JNV8K/GN2jVIo/XEjFgGyB
MoywinMChg20Mp5HJ4shs0OKSG9SIUp89bCbN2/MxDnk3pBaPRKCGVpbdsw5O5GF
19KF+d/byEsI9yrQ7CTyRRUsA2963e9T+mBZUVp+lranp71YuaLqkRBOvz3C+aWi
l6EyvJv1kBBDLXwQVnyzFXiy91VCpu1pPn+sYgpbdoqd3nemAoLCrx0L6asK7mE0
uySwxJAeMsxeaEi2xn7JnNH5IK/4dqXp2PJcKkOaj/1Y+SDPX3I0OsWkTyjSEmW3
m5T0/ZCx1o1WRAJo7fyIDRdkvVdF5KiL6ucCOI7hNIzrTmlUE5D6WPMeX/YMDG+8
VtVuy9B5EMBew7GN2Z4x1eSZ7ZU4yMxY2z8j+AgBE8E5GZrxOwLDk9MsbI2aSeCm
5UVbqICW9mEC65rmUn/vFTEYwum26pIIM153uwG29VA4dI3+nt3ucvodSuT1Si3E
db/UQCGw5hLESS1/dxBkfVNOKs0HmRSRb7j7sC9bu+sO/V9kEKG24EACLZH9EDei
gBAilwXkklg2SaGsgr1sV5htAH2GDjag7aqUW3maTBPMyC+yfFWDmk6dCtMhl0Aj
5Dy8dh5AQ6C8G1eMhZQjRXMRibCO2z2YfqcHAI7lelLxumB8QzUrKEug0SsVnQMA
ATiNu2DQqQw1T4hB1blVJtvbXk3jfJCcnZCT2TtRfnJYWhCL2rQeZHA5gkfZJgy2
J+SPt72dxXiiG10Qy3siTS5viTVogNfmew/Pc9sTgWpB05tH6h146zMuSF2OW5bn
/GzeIXkxRFDiNFr8yEgz+OVHqzVHD7DQaaoDTjHitEs42nHemVsfRucyIQJRgDay
CVn/NvnpcjnAyLPb5304JDcD7rt/1rLoexpyf1dZ36TZSarbIRJ2x7w0SLFACXYl
O28B8h3lvZj4tpA3l2QQxalRMQQzTY7FUUcxoGMu3QTnYttvBTWShBh6gbiZzv6a
VBnJucgU5xomzF1YuBlfPbGznzuqACGDqVcA4p0bcG2L6QtfxaIscp25P52FxFkz
0AhNdurVDssuL5Vkl5HwRHrSVVmFYA+c08EkW98AohH9B+E4xDUDEhAh9vFdjOwS
Dd446pzOuIkgidk6HVNgmjyG0j74rQNnqyaXm+uY2j3+iKdmmn3K0din5uPirW+Z
g6rLcLx25jnbcaqYzPk1VCKl/6buQH2GzVSNJWViBuN44xABKlNnGH8DN6RIJEte
iQayNS7FwbcALuPibNGogKN3/2bCiVq/1yp0GSvDe6WM0vNPwQL/+sW6oxyDHcl/
QiXFc1WqKc4AqK97S55h+rAd1Zor5K2wvdod3G39sQkbxx0BKwfYzpJS+uPJb9gZ
he/nkfGdEQ/yG2vusB2kG9MGDaHmpf3/cledWVbl2PgJHJVSix9aIu0nPr93p9GX
8A2RMlL18s8QiXzgiezyxda9o9thKsmO1zo+TKBoQUwP2szTF6mVKXPPyAf2MnfL
N60Z4L7C/hZhQfPzTJDol7ksmEGkr3XGkNUtxBJ/xInZCpgP8fhu5cw9q789dByC
fnAAmph9hA6VzvoQANVcJV16mnOBdspp1LOrOMktI5ckkz5JsAw8iDaPINEhaSIJ
geOufPH8Ko3mi+DoocInZxhfHcDBDKOucKtVhnGje8Pjd8QvLE3staSYgfqpJI2O
U3zLD+6nr8icygPFHcWmuRLhhd+Vu16UWu3BlLYKywDCvRI1ZWB6+ShaBNXp3Bu8
KAfu7xKKnpxwxnvA1NvG8F27wy2vhtwH49INLn1+Sddy/nO3rtXdnWn63omrwkRR
nvJ1jgFnEBwr1DfQlw/HSXEszB0FIuu+z5Lo9y1+IBc1L8IcJ6vhg3nKwUmwD+eF
XTbfrX1DG4EeDUDcavDcZ1HS3yDDF6VZ2Go+59FATAM1eBGAyeHeeU4YfqqfLA02
LwcLzwQs+cgYrxtSwMZlD3bigXyqAJ4r3nPHyV1v0avENhLA1hsarbAk8oW/yg4d
3cmNPJdcnwS1SK/GvRZow1MeptMJXvIPAXPNAzkU7Sr/a6FyCnI3tYAesBmQgCbP
/LLQv9zX86+FLXiMIlrXHta6r9w4BwScVOepVDpUmSKG8QA0Eke2PbMX8hK7I7Gg
08UggvKwRw+61HEdEyJ8kZAgFVImRhjRyX3UvGlHu/FMbRgPOF0MbsPXvY92ETsV
cmug5HcrmeEenqs/W6b5ohQmOTFMQKOIm0oAPFxEHKpeYqiFPhQyO3du+tJO4m7r
WotO29tMZmIcixy2FYZfsCDL3K/Fb3K7EQ681fwnHYo8hf3L4p/uyL2VieS6FUM4
F9k58DUcaJUs0wJ4zVr7BEC8AukOoF4BN6ewHOsX+sgaoq8klfDZdq78aHrWhqu1
ZQJy6f783ldcVTGYoHb7ZukJlfMNjcScFIpOAcQ044rdhaHNHgoq6aHixySfBUZL
W3gRgelTT1ak80LyRuvxNdhLDBM7BIsuUH0nxfJLAJhjAuw5ZGt4wIuHpxUbnH8q
H2sD6QVYQUdXtWAHNhoZHUOo81AxFdBBzr6Ar58NAGFqhQiH862ga4kxiogsOS5o
8X4TRl5a+2ZxC8DKJUbRL2niJASQ0jtI7JiDUQSf2DYG+eIsiSavUJuMBV2NbBmS
z+2fk+lZtMwG4zkaEw14MOxvT2b619GQn90Zdft/Jv1fusUINTdZSMp/91ldR6aD
VwtWWqBzvWC8bPhq1s2hW+fRCjDvk6U++7RNWnATaQ2klcmN84i2jLeWKj9tYZ5k
xEZZXXYclMTZ3CVV2JCmbrG6WFmAxXG85DF2lnlqcDCDMcLorv5JNWBdcIDrwHP4
ncouS9lddMnXpDbR45ePstHSZammQh9E5pa8A2uIBIIquEsjFalJEESf1XQy5vsH
2itg+mKM362DSm/QRkDPaFqqSDLfCsH2YEvlVwhoNmylej/9UbxjTbhfMuvFO9Mq
YvODoNCAFwqdjZR1Xf/HzciE43sBjAOh1eDmlWSXzot4tHdh0XRhSfObznhjsmYo
xA2hn4Xcsa0/CEjBGyK1FSkbJVFXmvy3/HRb85hQJdZ/PgUntdEubH1IWtcW9bYi
TH7iMMZx0jhCx1pAAExC07D1BXTbub+1khTiTNQ9LhZWs/H4YC5jdDqpzMOJ5Yci
GQes8/curDEBn2PprdZln75BhCbvkxOf5uFFdnsTst3QUyjyzZqV9B50u8fgpTGX
J23Vf/SVYta0Ek2Dy33KF6iPw1F7vsKbmFRMansTcPemvu0VIA6UG3AlAXH9QRNc
2gzqx9scIgI81CtjnTflYKAopWkZCXQHlTVzC2eBNPspppvnLUAj1tl27/jmZ1an
YAm2ud/Ld4N5JX5kAS3v4Zwk+fkD1uFEMsK0aATFZw+JJgH+QaKr3Y8qM2j2qbsl
ocb+JU/9C/lHxLTB2svWUHClMc+gTxuBEHa/d34TtHE9+e7sEgrE/usnWJzUCUKL
QhFO+wTGfytxknXUNN6MxL9RRPkQ2ngNd1qNc/cj36KrNMWQ2nFrTjIAUfgc91GZ
hK/zQ5foYPy9sifW001zy3W9Ptf3vvtWzur9NnP/cGM1VjitcnFuMo20M9DLiC3O
62WmtR93rdxmY3JjmkpAsWT1mf+B2zjgReTLI96fxKWDKASWcDUhnl/842vnK/DD
MpSwcWosU2bO9HQsfRFniMDyb4O0Q/7jHD+M1NWDkQ8CIGRfALzgQmDny9jN6cXa
llIxkcVGNCDfreVFOIId8YfTfoeDu+UtB+Kt5EH2pu7j+qlQNU+6Sjx9QbB1JPsn
PAw2NHBgPntLqT3lHNRMHnFXSY5FPpjHKM5A9gTXRYw2dj8CbMbXADnapBAu4Uc4
10KQWGqk7o3KkYdSTM9VYUjb9kBTKG05FpFuExJJW+fYPIDD8osjxAD3teDcazsy
wDQR+skSofQJJKioLQXhgQ4MdMhQDCHL28ffAeOFwGYgP5N+rACnX7B0Pevd+nF2
TrMV1RlQGJmppM1eSL4mkJC3smV0tOrK2vwgWJjfLugEeA5yGMRFUOxZypRU+116
Mtyie7A/tUS29S3yp9fRDz6d08mnK8VTDtu8xncrpK4RiGusmw+T/J5/63DWgdtP
jR69+/894pqNew59EkpNIK3t96rqqOOUf19yAK1fHGpTkBZMOJI8CLxz4Lx5qmCt
MJL9AKiaa0QbmAbFzjg2f9xJNIEGmOrSRlZXXd/h9Cn72kjLAxrUAy+MMdCJpLUP
irjrrvMqRrYQzdOh8ZmwnLH6Xr0PGkTwRfMBwJkr2iXmGS4D1dWf9EF05UvhHBoR
9WHhJuzroDIsiKekgaaxVy5fP0tDTo+VgDvwaW0UJn8Nd2ZLp1x5UQ4COZ81Fmf3
SSoRxQOCxjeCmM4pm4ILyprSJ335kGO0fuzF6GCnI+3GcXonx4chhBx4diGtphl/
LAAV7jhmwAbWhWDWuPSkn806gHyQMGLKWrGsZbD/A9/veMhA0HoHUhhXMmu/Xz2y
4iuwTgpSJ75SfFM2Imfshh6fb91uxyYSJ2FeJbe6rBivTnvFb8biCHSgDteFPuyk
rJY80b/4FYv6csr6Jqwf3bMzMmPsDrN14aLQu9M2yYh/BqND4mq8crR3IigC5ovF
O6hfqbZxrqvM5hkUWEo/apX+IPMgR0WFrc6EZMIMDCNk2GZUm2rPl/tVQJZFNsOw
fViD+TBu4v8rmC+Sr2iA5srduIF4WGFivnss8OUisSpabBftFIsfBQ3I/y0L9aO3
N6V+r733bXqpzvTHfPgjDMWc0Bmi2gl8UsFPsqZp6LkIooxIGm4iTnqX2f+zLRZi
qawh3TAYDCHIatcNeie73d6fOs47GvSd46/4OZWoAaL1YB25yjuykmDUqjXHQ4pi
45pvW2v8/Ekp7Vy6KgDCQX6Q+anWS13u6EUnBQntWZwHv5DLnUVZ6IGFulhEpSsK
sUTauDFdmre3zXH5jWrNf3graIYMxzdNSCRJb1wkA4vP+j6NP9qQCxRP49Xq2Eb6
kSPW1JQJDkHtIQ2G3SHirulWvDZwRqc4zm8qIewlbZ2zQQ3YNnEvcckWJWh7YlOx
xMOnQeobex74m4PrOwUgQhE3ZC+bPInPC4dsB4DNkRbxOMI5gnfVefX2B9xykDom
TNmmKdYXeYRwpVDq2Ss5/24ABuDDC8JJS8g87KOjOQUxEKEJ/0WfKTJZng5L6o+L
kzz8SRLcVBflS4jwB4i9XaNui6bi5sVdQ2gnicdI1yEe/TnPx4maC823cW1W+Oss
ZsIGS/MksGIbxmIaNFCnK3cJsqus6QZRypROxGkPRonQ0IRKmBBCWTs8FJmhasbS
kNysYd7IIvyaSIqkZGIudIeNgM5O9juvgox+J46LoUER04A+/3DO2pUWyllWTQCQ
2Ui+hw1s0TCTKulicPtqRJeCiGcvGNpOSA5nUEhGfZnUF1TPaeVDuI0OMT3Vu8Ep
VVYP6Sjq1DVbR+TJi1CFGPwANtJOoPImDE2yDyk9F1niZ6RcFPdbMHMRcR0X8Kfp
QAMkdDsG+Xdlh6OOh7SWj0LLWLUBZNOjDgQgvogx94NOHB51SN16R/92MnL42zRH
uw/s/ohl0pNOIw/RNl2zi2fzR3VTBVD5sDVbGm3Snv/4bTkSAp4zeMsGI6xO3u2m
3k7J2hokE5iNpG+f/+fSaowxDlkEjDzy+Sux7Vu8emk0yDeyG6K2gKODAkLTaB96
bZmWDOaUc+HdBpcXSnVYPmDDysANDA6DvP6Rv+aRF5RmfjH8+uIG0z5sEqWyIMK5
fQEa1H9Ky26HHwseljkGZ4Y1pMLU5+CdiHokyQp7ms/mtFMjfR86MgWyDqmsa6pq
ocOwHIzN47nuTve0F/2ki7YrrPdx4RCPwZvpUX8QcKkoKwtfizj/Sohx8P8aHVlG
BeEbifpGespcYDIhtH5CmxEPMHL/fqXOYa6jsdMoAHLiZcWEvpMibBTL2BU314mP
6wUlYFwambUY29e0uPk5QaOr9W8aWLLZSvi1MCOZfekrTL6YsyYRes+U1RIE0ROH
g9ijqrRW0+nwvblUkQ7S1DImmrFHqwj4y+sDKWWyZOXu/dLWV0f4PYJrXkBPpT4p
Sh++iispi5lvF8MT77/oOXtLuN58ux4fD5jO0G+RNzkNpTlZd5TP9MWpkG0PKoNU
U95a3VyUghKBhwYOw/2OT1XlpP4LPButlVjOEBDrJ2ofAgssDfBklUn6PNrD7rqg
sCQ8kxl0WUzOfUujupwchlIIXnptBwm0BbhpsDvxFrQhXOoQDgzvha4SXng9qHKL
rsRwmieu1ekzHlOpaJRh6y9Y3hcvgecAYSsEimuHLE84U+ljGpHfuoD2gG6fJADt
1tTV4L5GsVolfMObDFkbnY/p0ofJiUTFTVsDay6G8XlW66eElSeCqlFit3DNW0Jw
4u5hQcWSoTYfS07WLTfmeSgglL8VfvcyFi5ddHjnSY4lJfrRYgde7WIhZmykXbsJ
/7MfG2Lah9Jyfvy7BXQIUu6qkKzIHmPyqystp9Rj9Zw2qVvtTYlJ8iyhlI5BTAec
Zm5eVRyjOCeE7tXnn+HdxXtMNfSWdNKiphZSsfvXwMp5Ov6lrAVITnhgHqv5M4la
yOGR4bNJs5wTFFJgRMAqQVQXo+pbhWRnWNZ7TvJE1F7KMYFS19JRnJV/m1qF+FgO
5PEAW0SLWYnYhV0+dEQTxJTyNpjVIg3y18v/CYTj+p5LkKj9sPG0lutYAaoGYnPM
jVk/SaSPd6Td5/+K60YR8FpyFC4t5ZWz8sDtDEGAPyUYv4tjj8E1T+JpUcwnJSaG
gL9rmkxxGfqWttgWx5iIudwEjvfLsCNDkxlZsYTqkptj1gRAg1LPqswNvkSYMZvM
qZsPitaq/PGWiW8Gid9XVhHqT7iCR7SGTDjKbVvIESr5ZMHRrFc/9a3sK3swzFeo
yPLMDNLpZzC7OMtPNtzgWxiRq3V/8y+OimFH++Wp8DH/ekMyg5z1lVmc1dK3QTMP
hopXjNll/CUOXcuKrsnq7HReRT1ZOR9lrSFdfvhIr0impFBM0sVETBHr4F0TM/OS
wmsx5JM1a8Kvd8fYc/sDsxPYr1A5CIubNG+mck4Fp8KyKTQYVN3Vnq2LYXzrwxML
BSouAtcrIeEEIo1jaf0JnlluKxBC57yZ1jwVNhqaqzQn7m21o2X7eEtMlV4FQdF9
SZ33ApvH3IJP4PcIXjUeVztqjN7bY1jC51KtNQhB9ZXiMI7XwHx44ujpKMOK7dw2
E7a2RedA+Mo5/TGw4wAqc2wu7AiFTeh3w+ZOaxeBnnHxYhhdUyN45KKtHtbEtT7K
js6l6pU8LCt6NsPhoGcA4dAV9QZkn56ctY5Ga5V3YOJy2CfuJk9mnlZwt3/Hl4an
gbwccU36NgkRLVQE0lY6pXJt2lcmKB9x5AeaCnCbVM9a+4F8NfNx8txSSWiWHydC
+ePZaHJf5u1j35mE+69keobU5YhUfQwdYkoicww2ghL31Nxed6RrbXZhrU6nc1OE
URIUlt6pNzd636MbpkVmpFznCFAYoGEwJdgRFaNJMWgJPnoCBos/KRMTDUPFrAbJ
WdKZphfGAmG4T/fgISvOD0tI/DnvoXXo6Coio3j3Rsi8iZhJOnZuvRI27TleJtv2
FDIRozYUlukVxJfQ1Flepv+xfvN0FdyhgR/+YLnRxW7C/FOSjkZLm069k9+2FQEr
ZDy8DVmMi3X6z3KzP+2tEv0YeWP6AxRZzk70d7Jt2hGcp4t9XmahVfkvVznmDy3+
TEYD7xaeWkzyS0P4CXLwqXQnE2JmV2AJsNxcFlM+vwY9rc6p83g7pG4KKMjHuK/2
xEfpAHIrgiwp94mKis2GMPeutWHRnzUKJGLmejnUZk6siJVlYGTw3PTB3grL7RE0
oHkoJktTyqmN4pOTDvxFtIZdEX9jlSucBs1J+3DA6SGLG1UDZu37O7zsWwQM079Z
tuIsj5kQMCA7NJ4mtxOePIRLtH2f8W6rOSE9mBDrbQorYa+qYYk+XwN+EfkLu9nl
saMItnu6bnjhSiAe5/OpauIlF55qF0Br2bK7AZf6sLjinWB1gn65jD8Pf++v9c+n
w1ajVpa9ND4qzB7+sbKexNHVZv+3fiERXdYsXkFGHU2tNg8MGuuKDHfFRdMolRzF
ZYUiZeHwTntrmz1+emQ4bp+gw/Td8SnnJAfSZYMrTICkRe3FpgiWwwQy13Fzrfh4
Z2Wq11MzHuyeponCt0rEtbAUOPh+3j92AwNhRwujGkWQeXvRfEn+b8mg84FKYbn5
obHRKNsRjInIUqc258lsPj7EcV7dz/mau1gX92yKVzjwGqIMInXkWGIhL6E93RMO
eipYpK9LvitqwUtjMH0OCHfERl47P7dxynIP5ULw3cI7S3SGY938yGbJPFE5W9+q
XwDgQhvry7bKpPT3M5CrOyDdiiEHyFHQy8BQGxWNTeNdSN4LfC9+D4KUq6H3GFz4
4w78rYIsZbnIj2rDaGcLQ5S/fPzE0UfI/vIwFk9LsI7q1sYZlLXgQ6i8v3fLtFC0
RLAJ4PsgF/WCFnbNQZg/A6/sgPfuXY/76VenIUtKHhgAiMVS29VvzrGfi8KJNaJI
0P15KSK0UKUvjZYa9ekjuNHIXSA7gvYQrM/Y2LWR4rVadNIOVUUkZT52S2YR5NQq
fc5AX6jfdkioLNDPtKluLXJQt6mwNqAfQo/fkjaEQbnc+uHFpr96TsV7LkdTBjJV
YUNenuAeReqYIycLbfTT6s0kARIQoe4CSW49dhP895W3aBSl0EBu563TQ5uD3GGO
4amPs4jidJGhDr5MhQfTmHD6rye02gorW+B06/0vqyDSGg3AnnX1nji1bh1L+1UC
df8gFOEw4mwSYQ2L0n/Eumb3AGWVDxvjOT8YVe/mUqkWxqixpObMcK1IjPvRfXNN
v2Zrel/7p/SevaOYGZtYJ+nznkSNc/Guj093FiFB6qj1/1WGox/0/NCCBvDhOOjE
47hPvJFK2s3SPx398OJDxAHE2bgxHbaWCSH9kxJOUY7o+n767WL0Wnn52ptM0oJc
x0V1IbfQDoBtqvyVwLohgmCJEx5BSYY1nT3arRK5rFWMdg1AKVzbWjW+RMJuESFQ
rU9VQC9ixbqgTcGnIBqiXNe7jlo7Oh8r687Vd2A5vk+sqY67SecY4yWAkpaSggr9
Z+4vHCj9Io/GY4VC0SeKX3cz3fhFX/sGJdurdWu4M1w0rR7NsGdSnIIC94upuqF0
qiI9JAd5BniDrfQzl/2IXl5n3MLuVxi080hoJ4aOOmmmyud3EBIQrdtvJbpFv5MW
L5KYbthfSZt8QTScCPtuydyaoeTB+KPTmyl/LfIf8jzM90A8p/6owak5GvBGLjg8
q7AHJeeRs6jQrcSMoQqATagpYT+MtW0jRLaDko/U8GLP1zzF4kVt4RnfJooBy06k
eflHPOhGPjlLI4vGurxN6BxrKxFYRCAg5FdrXwjC/8avsUFsT7IyBdS3Csc2WVLw
T2WDFrdJcv667dhfxOdw1Ojyk4MMKJ9bWMAS92PO0EacaoeoPi1maIkXRGOYfTGX
IwG6slBvd0BVmZC1NQyrmJgC9ANwMPDNBBLcV61acrxpK9k6vDRBbv2s6p5t/EoT
+JsLKzAsymCMTAwlzhBmnc1DTkmfckQeaDANbKxlxZYSW0E7t86AVwsVHwZDomJA
f94ptBb9oQdwI2MXoTBEceZkFLXfcYARREB+jxlweogw3zdtt6jD0MRWuiOFE6Vw
nQ9ra+9L7QdXH3KXSk5wwdaKoDL6D2cc93YovpkvRhTvCrua/YrYtYGo1X7/TLJ7
0u8LYig8rVoqlRIvrqbVd8+4ahv+PQT19F/e9DV61W0qxvUJjqLtmeiGMLa+YxM5
DIesaD+6O05hYPGAcSzt5YYFzm6KAoYJn1OXYC8A49MTpqxu2uUs/oEn/0gRcd/z
7AhF4fp10Cu10/nzlq5c6RPqlmo5Avd1bvhdD5jfGtXmWeHVR19UFpxEJnMbjR0x
Wusn557zL0XJCTHbkdLEB3KJIuXzwDfsg1KzQVhzkPeIjNdHiGdIgA2knWPzNvuu
sAah9Qu3DFwG5U+kFZuzr9jdNLtvbiM2xNPsnGNN8Wa7PPgqhfnM+z2wcN1uzoDV
Oy5Bs0ddkYXiPrcoGw7l9Eabv8iQys2eyAOfw6ONzeYHSzNe2m+NcqOX15cTj770
AznQ1tU2I3h+BpTa4OR8pnl1UoAeYF+f0r6MTdmx+W479O9uBbmTAQz78TkYuD/B
u5pupK8IpHVKsKF1zLzrhRhPH7LKdgSZ6ou1f6m9bce2x/t1VsvRtXcEUvR+NAPn
LGZ4o1nQO92ZhNDavkTDf8oAJOh9d4h7pg7b3ULImplzqdNNJDz0UDBzLB4hyFnn
4/zzhd5tRN9IXPmm12Qu5o+siJdRvhoBXVeH1q3tcOLCxD/Q5kMbgOWICwijXUKD
6mVTbtm0VFv259IUSAcIe/w9K2TxMFTRc2UavJkogHulJaHUri9G+ARnbM4lsPub
AGz95v8lvVFi247R12QKJkDUUMYDNXilY/k6Q6HO6EV21PpWuHyfKlRErQ5lPGjk
XpPt9HgTTDB8aGO36XXTcJmsAgYZvDMVHD5qOS+uGaA9YR+jV6x2zFFh2gCmJYvs
TsI/VB/ylh6vfkd6nsMa0CApcT1LuZfd4/UCr42tQv7eoum34H+iFCL/8Ka8Vz/K
Q5B6ZEgYH0nei5MkcCntXExFIU3UFH1JRcRxXFJxEVKZLqFZyMVzFlQCJ6yEit2/
KIYXKzAnZ8uVzEy7NWBTVBDUCTMngdzxF11RVwg6w3MT0L2pOn42qbBTNU/9Y90O
qP7TtDBI6qlZ/PnnGeGyp67jqgR11HpgZRjNGVG7+sN58ykDqr/uwqAueB0+8+Y5
YkEmxqldt6d2knyBwX3KtKO/XNSONlsBCq6QWfoHE8jKaCt1wn0tn/QEuFZ9Ivj9
E3pSXljDUDV9kdgV0k1SJsJQh7frVO0wRXODmSR9bV/zHFs/Y1BCIv59kcKJ1ClQ
NLhY346XGJZNLiV2YHfRQRLlVGX9ODBXRtbLGCKt25n63eAZk/roZZRZQ+wCYXQg
ea+3eOqWPONBGkUFwsxWpWYzH6kpb4s8WTKP1yhte3Iclijuy0LpR9F6RxkCaFLw
TcGIGzNx7Gz9w8DhXw4q2UfQwDdnZCk2tM8z2zx0KQApvZnluZq82q1knFrS69Xv
/qOzJ5rg1i1cWZqakdtgbFzOgjaDj0D6v98I1w/8irmUuPTUTFvCYmV04YYYCfwU
DkSD2YduAMZGLhLQQ5BwCOC2Zh23EVzIxknM0BSfKO7Wi/eiAWxoZnatxsvaIz/s
rsi6DdvbIqaJLztQ8RoYAXlCdSpSO1pQVQ9HQhY5xxp+p0dNQSpYVj0bI9zwhxCj
XuvXIisuRHT9hzYIzfC/wvAhHEbY9UC4lNwiJjjh7IZ6U0wvdYDUFEdR8jYvr0p+
7GfHy/yCMqpUQbeynwZLw82Ddn4ridi286SZE/kv+VjRj9DmP7uO7FvPCbWaPO8z
NyjYUVNGuiZhn5oHGZ0ZBklRpzPhTGNxEz0nlHLV4uXLcP310cZ6H9dgZwGnkOds
EjCSs2/FGT46MZ7mTws4m3XXBDrWsxVnzIO12h2+SxCTDErG8sNAO1DTq1LK7z8l
n1+BX/opCG6b7br1dtvkWYb7IbysFCOC5XWFDO3QPYtVCo3taj24vaEBEewCwPSA
+ysVtdXp8goqKmlv01ssuaTV9f7igp+FfVjMh+UmaQ0cu5gPe45rirPZ3EsStAi5
NJAW4GsBQF6STZO5Is/new8i5x3Q66QoJNxxFbohf3vLqRporNpnoD4HHcCywJCB
6RjsxcEUVF2Q/5Eeeo0IcaiaBc3SVh5zK528aQIw85nhUlZmfUhUYTbnojYUDer4
5te3QN6ArSeEl3MKO98wF8QhDFC7474MK/r7u4bBHejIUx6b1JiCIVTT+JiXjEf8
kl964ioGaI5ba8GM4UXyYTveKUitFuqpriUn0mtexUve8vigRZuOZtyJU6lMjn2v
xmXNDAlk4edprbjyAT4dMOlTLAdEAM8Vo0UGt0MSuwkg9sRsS/tnylHOjMMIAeBs
iE/DaWm8vbqHTjnmFpNRBBKfH8TMmyMyVL3kKvnSbBIaNnmDMXTDqjlLDLkUrhe+
nlV4meUkOHIUP3a0+zz91Tju3bK5hjEcl2hMGNBLvFzKLO4iafHWRMpGqjlyLCC3
WBuT7onVtajEBz7Go0gTxyFGqhnm7MZ542XeacD3ub4oz0o7HzEf1vvqVFNvvqcg
+ZInMs92H+QIRu0lbbtZglQER/zja/3HARs3OhEJCx8k60/AV0A9CGTqhU11Nqdq
/pCbVB1p3RnIpvP+8sIb9ilYrmxMLBqtDXM8Y+ePLTEobVRenCInJD0gRVvUoquW
cIIOmK6pr7DgsIlwSWX3fKORq3q4xjBF/vPzioXV9THNnWPXNqI4ujUR5mNdVAj2
MhalWeL6uuuSrnLIxPdLeu05ypEsDa3Eit6Z3ilfownYnULgzjKgm5NqsyozZhob
ddmVXXjzlbmI08t9Z9YdNLZ5MAD0gfbN1vF+N3ciRJ/HmfT2wMOp/PN1xG7U7Av3
mczvCLh7x75WViY2QXLfgyALIkyoMrLoB4kXk6T39roy0WI5Jb1W/3UH9ZbZJJxE
Axm5WmKNPc2oLevo4BKzhbJYDHJsGIby0rs2jpA2Dxpp92/mrimfqEVv/vVCfhoZ
3r5jG3F32kv6uWfXOkfdLxoPP4wJ2N19b7ZVX+szuKl5Ebl62sa5TGkziv3JTyUi
OlynzFA3Lw4O0iywSuShwUgjMvZDfPxFytFLx9L4rVmnhKLT5WIOiKCTLTslRpSK
gpj18KgDMz/ljOn4FzcBHwvg7Fx4TEsz9nEevAnuJjbK941ILD4J6pjXi8ZmvGQL
KPJ8yEhBMP8DAen/+QdPjKdU7wbjfqp4cis6ro58lTmnjvDwouZ8q/OTJ95JJ32K
3DSAwgdE7KN+U1vyGYkp3/34TLsBoxlnvK+ZPgcmXSmjTa//uKOg2G7zf28rx3vm
4Twv1f4Y+NrFSwCYORSM1MczepPfDRWviXStef3MrMM5VOhFL18I2tEVyb87ENAk
YQc7Es8Dm6IT+Fs/yaHaEb5WfmhTk4t7LawXIyhAatZ1iwB1t/apIItQRNFyDE41
qmlLQ5SFRZv27I8qqf6k8n/ZcYhyhoU+hbs+QXmA7eTVsWxRVC42w0jqMZAdGwZV
iDJE5AoPbadb2LvQAsNgYqI3juf/flPXNqjb+5+V+wxz994B1s+qlxls7QJf37/F
pS22Rgz7ioP/v3YYDssc4Gs+VHA0Xz/XloSRYC1bP8KINDd8cwFzZtFcS8K1A7GN
h0vFehQyn1syOy2uWxC24G5bTkKNld/QAUmqBC1l/uU/p9FePAwvpY5tzyGCnC9q
hW20cX9fSdntM6l1/dGILmfyDOHl0GCTmDSwtclQ5hBw6UeBWr96pSUvmLqc08aL
OrqDBOFHdII1nKV9EJYOjVgjDG5dXnIl/awD/Ao/uvZdQ9xTTaJvSbhi65jxu6Rh
jDeJWoYYACHXi2ir9ZZkSaAOQvfc76Uv0AirIq97GvhYjPkwfydNLQa15KPN4Spx
fz9Ctf711IJXAaKh9qp0sCLsSj1WtfvST4eveA6mu4hTaPy8lm+CX/rNaE/QUCg8
p8yhj8yOqxyVwkqpeDJZx34vv53vGCZkJXW/IXATMV1EcdZAJJk60gBjNhDgqK6O
s/7HmxN6NNttbG008zJvI1HfuJPfSo7HnnC2r6gRHUDf68MN/s9XgfbNL77F3BI0
2Cxw8xzqzjwesgznpakArP9Yd9nBTuFvufQD07XugzAOf64+eai0UWrpF4PC4FBX
TlhaycsPAsxaeU+o+1h2UMcxjBU0rLPDUPRqCVDL+WKu2poFL31LVTFqW4xw2+S/
1hBxr4RCsTFFe6+RHEHQgQFc80rg+1Eii/dJ+Sh/wLZbpRoKpb3wUD1BRZ+4JtUK
flRW7NEk4j2FV7+1TVPaQX6TF9ySQpWFPvviURQr2Wsepjm5oy88BGLpXje9GL2f
9aglPDXldtEQmMCasX9MHV0OU5HK0vMP5nsAZEa3jTSRMpnF1jQ/UIimhzvRYX3x
/OKZ8RRIu6UYZ5RmsHo9CQ7QLz1vZFv4t57KYCvY6gVeKDSOLyCxicnBmrUBvPmm
Y8AzM/1znb0wfBxD/7dMzlTX5kGdxpxgWI1Ax58CQ6fNy26a6C0kW+dpNMc2NsOR
Y63ofzxV/IMFBH6MDDeVXJI6Mtf+7ElbrzLvG4mXqDB4/MD85iAnNzv12NHQ8dLf
q1P+BxJz672nti8sQLyKIprdV5IYkGgOYujo28bVBYpJfy4LjYfIYm3NJ23bKJrl
7c2y/GHxJCjIbfF5gFpSJrLkh81mgU1dGGaSvjXSPq/8+9D8zqRXmyjf1NnHvBgM
IVz4cRaRKFSrIp67pWk+ovySsl2EB5jKRAuEOcIeejRthtbD3Ew6/g+AD36fl5no
lSmvolp80J0dJe8HeX6/4LF5Ij29QtAq0IOwsi0ntkszNgJVa07v2BoqMCNvCjFe
NENgr4NLoqFbQsMCiPcC5IZB2EBqZk08k4q7P6tE9hJ16Qvsy/sq2rjNn0zEX7d2
Xy8iTOteIoHEy1mSaJPD8yjqKfp4ErQ8jLrJ97d1/QGSJbGarhVceEGC2LztLzmn
ShFYCxyb1odvulVmiQ7o0PE17WqdeMp6X8OcKGlsFZHj96HOFwRXHurgkw/Oru+k
sC70E3rhg1j9cfWxdBRXmal55uZx6qvGEslbuQnnbGD8qrjqbOzUGb2rZzgSuD3j
1zwLAFocrT37eMkYVOByUIoWwgAcTHKLpfR7PA17zv6tiza++mUYEdpnlxJ5s+j+
JhE+RTYcu9x1HyRTBaZtM4bTenKeywCOtQe1QH1OV2f5hOC/XZgbHGvs+5OtqASA
wmOJss2zfOyJjvZwYU2dpv/F5eTqjV539wojTzuku2zU756kOLQ9+ADZ/mWtBEEV
kxxDkeJP8OPAbZVXc35+JbVQtwUhe9mcd9u9KlsAyvDJ4XjsBUSiufdl+dHYxSzO
5KTJ+v9BvnAJWokCRRj9y2QN8PqmWHS756E4ESPUfN4NyivyXMFUzCHsNuQuX/PE
h86c/GAkPZHx3qgep710yvS3G8O55/4Mram8dH4qKYcbJLuEUKDgdSeNnR71/XjM
hx6/n48tbcm1G+3nV8MlLkhXUHWTVkm4Bmph001ZbzBMR0Fx2fMmgUPzTDWLa/MT
bXZD9pcdUUZ6CfqJF9lttm4b6QYKxK4vKnmwCdUsy0VCXaHf2/0upVTyjfPx3so7
Y4jqUoL0gPwUhNtYqeWuXOqDkuUIAZvIrR3KDtM+RrDvYwIxflmeLhR7OVIaeVSn
XCsuIHQRg9ekQrzaEcD5Il4ij9SrG4p8eEjPeNzbN5PmqtZ/CRUe2ZArzGzJ40je
R8iV7ci2dzB7KE4rCKz7jEoLMa2kZ4iM6uxnJrJzlJi3kEXzk63hNKK6FgH0a5KL
SOcPd5uNuayvuPNoPhGDR/1oLFDLRHiTmbuPvg/5b34vQ0ofw3nLspBeNYEW8Iuy
ewqLMWhVxd/xhOCgIzrrdT8mdycgWxUw6PxycWW6LZyUeNNt50GbVFYfjKuTjeiz
cNNv6NzDndryBOUMhCWdBMpRR/m9P86qi7GtdHunwjM1fETGSzzlx6jT4JNGai7I
DbZytgDoOiX9yNfVk/ece/TvLmWqfem3+drFSNgkP7Tg2HkPQDIm2gIDeR7Gv6dL
o66FAzEvnMayl+GXLKKPbczfs4bNrQpc9G+Ft9cAnpepquiRb4popmVCDaPFKiAG
6eBCGVpq25X4Hiv8MoGyEisi+okPUg4Ovp/nZ4wdOlhZ2P2cZWIovjONdMDYZBeY
t+h8pYcBhHUZu+VmujGY477W4/n8OCYw0jN2D/acT23WaoyTHs0ROZIEn3qq9bwp
dfaP7VJkoRB91RUvXg5b+NM5J6PiCSepZE+BxkZkd2dwDZIsomV4IBt94MO7NnJG
wCqI8VghWgfw1cID9uyZQ+hjL92BdPfwBddgytt851bgraTEQ5aZalmKA88ZUXP0
Oadiw/NF0JbcAWpeHJJqSif9vYyqgUBvuxVH4HeZ8HiMJqBlfpl7xbTYzCtQ82bv
9Yw3sUrYDVbSTOc7zKNtDidPM+DeCL/qtu/tb2D/lLB8SsSY2DtV/xPGROH3SROw
Ck/e2VVlirlOm7qa5aop6LPJXwo++SJ7Yb/2SslSS0yNdwPoRUZM9VELhOmSw23n
HUPbf+9HOpIGKns/15MCbAvYqi47pqDvj+Kky/3BedQR7tBMr0c3esb6TFX0T1wh
E/z/1dtNzyeUUp868QtNtM7kkI7tOtm4NW3PkiNVqndgxZ3CgYcZ67Z+9/e+yHQE
dIo5kJxT4irgcaJhGmnWsL2GT4Wdi0+gdxz+WV4nC3WIBZ0F2+wiwGjwDymhYVRa
PjNKjUplj/oiKAw+ZGFHwjbTMLWbLPsP1tXmTg37R3SsqO9r2fxuOBqcTcF/2OVM
vRnSwedocVRHPfAr7/o4BstZeieAQI/9M1FnovclwIZjEuxuHGBlJ5FI4m5s0Tlo
g/kFmVEzBc6MWX3BDOJv0W5Kgb7dAObiM/MVUpGgXIP4FXD9+t3Npm/obEjzRUPU
cbXhQpjMfWno8/MFXAc93XWpLQn0vx+TYzKbUruH3W7cdT+xIpVyYP9zAfJqXYGW
k6jO1XlmayUa1naQ+11z7FIomGmUi4UneWVdqgFtGCymmHZxMzlOazp2QxOZk77U
5FLntAgq+FD1KhdZc6GlF68as25dkyw6xUU8u1t0/Evc4GBrEXpWq4+yN/zBa4MT
k+uiOXrpimqyJZIIQZYbmgwrrG6uRBUf4wIbSJpD9O9kJFt4VZtUvYweD7f00w+y
BsXIE5VXgKS7alyj4Nap9N5HVlxqofj8d8uXKNNyTeo8JMXQWZO2s3h/9lZllXP/
pvGW88imsqf+kLd0yBji0T/vugF9Iy6/hUT3joCIw76vNxNZNVhgDbdwmq74QYwN
Wt3F1JJeaxGKn95uoswevRu/LVy0WE7XnXJo2Mo31lJttIw5KpvZnepViC+6Qo7E
laDYF0/c1cAixj+m+nRSH0ur40+l4IcYxXy0BZb8TuqMxR0BO/2SoG6R0+VhM+GE
qvYc4IR8nf9tPnesNJv/opBOz2hIM0Pe3j+GLFRQnx14f9aRD7bNhcaKlxolVZFc
AlFuSdn++5fcaUkqP1jj4GB2mR/jh4MI1bHdY5iYidtmNFl1QR3ybrBRLetZh8sM
DReogiIYugFk7ITXnke4XMBSwj8aMhoLC6nUZTT1lr6r4DsyWNxWdv0xaEgOswmh
6vFviYtWEbf/xMqA/qqkKl/I1nbNWduLnoPD8SZraPjurQFZf2H8q7m61yaaaBvx
0sSZdfJTrKqA33kqj65uUkpVeN4wllflpc+FvU4YsirnfEl79zmQQMp9P0TzPhcq
mZChYOPeQViEF9l4+VyoI3MzmIYbT1IhWgpo2C1jIl9P2f4sHOmbrGg14mYqTTjj
vB15ZkpO9BFKAHHOHqa6VFt7bVq3TgW2Vj7miCSq6esnx8HuhlzSshOd/twWWkvc
RqIrN2NqrwhQeKQyIbAw7CKXt4km8MVklZu3Q5M2jhZOgz68O5vlNYlNefEd8sIP
tClJaYOe4SHXOwnkYZZn4NrinJ/8gzCYF4pyAlSNUnt4mMHFBVkh31XPOtH+NCzS
fSdMCg5uvjZ/oXFYlgYXAQq4wB77WB5CkejbpU+jONprBjDj3K+LomB188MB/Hik
ziCKTY/jMfvodJuxZlHcSnPDC/MgDyukCsqccjetwArlkFfMGGTT5Z0ZEG2lxef2
MCBb6dYJd6EHwc7JFrjZ0Tg5zH+RURBi/zduylwRnFG+W8IqgtLTELGklWI2QUY1
L/UtUH2qKFXmxyeovK3YGN4IARhNdFNWcmH9Z8sA/cHKBdtZGcjGEqAF9jFD3Oyy
KxVYeuj+7oeVVx4bhoUwugQFN2yH4F81gug+amC1AIlZ5c01y946LcsV+4h+Fh0B
Z0fw+sHcCU3N10OjBdOWuoDklU2SIK8AEnWK4YgJ1XWTNfQ2OHZBFgPTYZgdwm4L
AGkDE5dNSsyiNio4Q8l0RWS3PLRgNAfn0gj6EOJyjjUbEl8jREfhcJEL1AL5Qx/g
JPrt+q03N1dK92a1ZUY1bb8f0MJHavKWxTa6JhVAM6tHOywctj/lAZWlX5TXkwjW
+9YixMmX91ebFS/VTdI4dubPsNoVtJef+dnsF6KzepcpqxvQWgbdKvfip0WcrQAF
a5udHJTdDr2Cl2hJc1S0Gv8w1k1d22+wkufrDonDahaaNH/A9bIFQjgljXiQTdfI
alp2iuv6ZpSA2GYzE209YvqPSGNjMpzZYA386XNcmoBafYbE5rDOQD01D8Pqxidc
yETdD/VF2ZPqdXSAQDqlDpUsa83HtLvsEXfEEMH37DdMOLmmL3JzWiw/X0+go+A7
/h/m/yZZIukAGKuQkkWpXcqLDcXk3heA4CrkrTppPCPhgSHifOVZvEE5qOFOrSRu
Tnw6+oNJkU9Y3DChsW5iRy9a1QUEI0In9pi/8yvprgYe4SEJGvrIpX9Dh5MwLwe5
NddWvmnixYfT2iUgYUHGF+NV77a/sp8iL57ujbyfs+TLX+jNYSgZh97zmtlHAtuP
HQhE9/Lm/A2qIubnGBh5sIrmwy8wYbUK2tOcm3jsYW0/Rty5Ek02fwQEjQ/msjni
SoB7tUALXYWWGLDDNnMGlvHqAhzixX2QhHZDnF4GCBHpaZe9wu9HvUkGxiUOPJ4P
jph+jWVwqoKKspR7zXJU0SXJqScowCoRT9AWTTxqMl1dH4nzML1hul1dyjZMOS5Y
qF4bFBROEu8lxtsSJ0FdzWbI0DX3HpAWrZeCKoqHJYJ35+tDqMTXwEezxC76qqP9
gBw0g/y/5K0w6sA7/ZlyZO/LysSYMGyqefk8Owv7bndCnwJbeeGg/bz/xcpjjYuY
r1L3fB7qws5151uUkAgZTFgXqFLhdpby9xijR/Kzt+Cv9BqDnmJFKlL5cFtlHXix
2nQ35javFpFAdhuEhN1MDbP6huLrds5tpGpP5nJZ36Y5aGXhpC0HR5tEa/txLvbr
nhnHIg3I7pywePJZd1RYRFp9Ies0S+7H+sFN0zN/UA3U2Z2zlBehL3qMKA56DD49
55Oyt+qzEzgs6BDKkSH6cwYi4Loh1u+ta/Z51rdao8YqVbcPhhj9JMsVz8WXdK/D
YRu5c4cXy8KSRvT4MNOZRsDKaUCzopPzGL4WsHMcy3+1ljSuDDMWefnfMvfX+ePV
+KJcntKFwwe7wBlLHQutIFfTF1MQjCQ/m9cKafXgvpD/9uk0mobAcyqZhQF+xsPE
Jvmhu27jigzPerHMRTWTHQAy/nKl6u/AIHHW/haoxJYpNUaWV0I+jKPZHzYr30Mm
G51FYfa6O11r9+njY+wXMO+aBx91fc5aMo1wWuy+R+GaOazVHFMlFkeAUC2BBlRG
H0RDymbiHo0Wm/qlV4x2vDDj9DasPfoPQ8IB/z2mnH2DBLTmBE7mAQQOuGvJxEP5
jPimphAV4W5+aMP9mh75OCxQ3E3WJVdijVBIAffEDWlS0X0ZEafuoP5XfPjzFThD
W6alGb0m9wtUQHRSa6lla8pPds6hliIEM3kwyOsixRyasKz77Veip+TsYRKMofxA
pMA+Aq3caFgfF4jXlr9dE4w5FCx3pkwYzifGAppK8ZL91ZH4lfFCrSGFHkE5BhqU
P7LMsQOYfX3VhG1p4Sbx6YUFnrWyFs7MRl9qSWQvc10MZwpRl3j/f4rO7zornizB
I+59ArNIka92tzgNvihFEKz4AO79AXJSfn/N2/R2fIYnzDquQAS8CoQDm1SWN6nU
dC4tDCPIu85aeLsuH06QaQ7EKf4H8Sk2fW1xYtPfYmWdhyGs1xqr6UpjAYtnzO0O
FhRpgwfwUoVXO0y9TA4ZVX4C1VcjGk43wm5KIFZvss91WRX3PDYFOWCsPtjKCgcb
aqKPKpRsQRvyf+ftzQyraSXIJzypH50uJTOvEnCDlW2AKEPyy+gcBv/+PAtAd4oG
3RCYlWB5aPeyU99XhhTRonGB2fAqDj+TyX7/QNrXK8N5fffVVC/61LGNRObWJWe0
cQfiPANBzTF/+QnxDUzAR39HSCRJSW0hqRqn4d3dFoacxnl81k5wju+cZcrjUcdx
28wnh4rB3e/PAQ0ZRVC/Ff6NK5csOaeyVzInpnTyBWCTXy8iWHTMl5LlmTHGc37H
93B+hIdc/91K5WnD9WROiBYTzV8XEBPCa5rUzj1Vuc2DLXd49A2vEDvYhnhsM1xQ
2JqTCL1mUnno9xzftcUR6UmX9L7/q3jC1NKvdl81Y8fYF6kpG9t7mfxOqs6SNIB0
+4t2200i1zRHlZP/4nOUjK7b+1qfrzA9EP3pdYnVDAIaOy5GHJPg69S4nN9xgIzF
r6uK7xFdQxnhUwxvJw+jfL/A+oIeoHZ+5AqBCzOjX5ZBcrvuPyhUnPRQp4PQMgtk
6qAG3eoZHBhu5Mb0EUFb+SUMYrQH4ubfI1zbi5cb7vR7ZO6TIcRUE7aMjNdxA/A6
XwW1JtFHHtpwshbGwrhT7xqfuvNyU+OoSSivhePLE0T5ho5uoQWum9MdThKCTTU7
sry1XjMJupZlXQmtUQZYJEt4cULgt/LqxR/HHFjfa6rXH0FCdk5CXN5NudbWq8S/
7j/KvenRiOsiTc63VW5JXEU6Nyh7LrXHqIX1nac9SS6gUa+0O2EcUks3MipLriPB
nYDNHfxTirxJ2Mn4GLCGarySa7f2Q0lkQnyIt9aoY9cW7Ss2szBkWAxKfzNHjJDe
F/xrGoWCGmWlF865Egxeg/uWvQ3x1la/6BBF6NiNMVWmd+tK/1HZTwFcgaaH5mkv
udBV6QwwDA54R3WfWSRP1IyiGhNogs0snvJhb6sxcZWtVYZqN7MFmS/XbrxB0ArJ
Hl9vqf2cKu5fJEW6hXhKYa5K5EeCBf0PASFl6hQ7LHMuDpLSJLikhcLWvT+ouNia
9QYkVXscKvzSHwW8wT0JlzNOCN1l5lp7tvu6HPBjHEnYp4JMH8xTbsLKH4XLhZti
CGY3+8Pjx8sjRY2PZBw0g74BK9YH9TFwFnvxXtB2TZKBFpVxJ5E/e949Ai2ZwU1c
Tmo+O1ihwAELuzoIuF4H47Kni+AUzLxoBYI46d37UNec49wdyKPrVHucX1jhlog1
AMZGLNXKXP8x5QGmP11dsSrrFmGzGQrWprh4dnM/bmlmXr29CiuzRofNugf+JAyB
O0QAD2eOrWJod95TcwAxnALqgliuILgOvrHleEZ+OBd5PO+T6q4m+haxK8U44Hfc
fPVshC9DwNGT4JwYF2Zwf73yVhZVjqanEqDbU1zi/sfuP9YwebbUrigoeRRbXfel
RFSW1/NA3w5fMmHfVZBXaj8QMdEVnWBHxFP/QXwGb/q1gso7BbL/INdTfv7/Xl+S
8M/QoMb/hKTheT+moSheYykjlcPS8JZDtxe9VZuoxQQnNClLnW/C2fFWA989eGN1
2qX70U7uRJaFW+E5967cWC4gzzeED8Df8hjNwAuejpHgLl0eqFHyll8ClsiGueck
uAt5Myk2A4cHaFpLAJeZ7duRQGflLhLkExMLM1uy1cGPF0dinv8tgVewRPc+4KdI
RuTe+bCokVCrzsJ0vjG7YkO9XxQWuP078I0HLfULCRK2ARoo5WAH2JIane24KnfV
3iGCYsuOJv++7bLoNEIjfzjfzVwzX0yABg2onSz0plVTg5JkEMMr+rh3tBZXdcGZ
Cc9KcUNZNEGYw4kr28OZwzOZn72XCrHepL8R78xJhiqafQc+O5KSx1qpXV9VSZUu
0FW2CkiNZSHz8qkenIZO79U6Lg1PKMNCWCXeS1TGqgR4g+fXzH7ZpBpX7E6xdZsk
iwMvigTq3W9mq1VkGunbZoZIvnfJnB1pnkAWEw0Kf64oVlRu8WwROjg1Uzcf1KCQ
1ywWscv5G+PnYpS6stnD7+qA1cJgWtxVzMuxp002CPrUgL6IsK9SRKk0wItnYuA6
DWWlWulpJsTwq1a3wiLSTli2wfGqwnp6qEm5W9tG+LSzR/YDQz3VP1lN85YHkYse
M9NvlzN+NIQXs0ZBuu/cWxuf/IIITNbri1Cdc8AxmATRxRjneuEWem6mexOKzmLR
/dCpfhKiCfbhL9tcAImcmNhn7PNbKS5tYVVsivenKYJuGpDxFaPaVOW/96DdmulO
UzkjrzVAjN/QG0Y6blyf0VIBUqCV0f1WjhL1r0p7qYVGANLCdvfz2Z+VEaPQbk0h
MXtRWorcCLKI8hjmeCBSOEU7IRDyvreCCLOp0KStmsq5wnlepjSBikYuSZkXrvZx
yPtBXA/gyNEPXNiDzEI03jobrgvm8hFbiGlSMuWIvCa9k79s2VtfuCNrVbX8E3hc
7mo8J/4liCtsuVWkCI2fveufwfef1RFyZDH9TPE9dp3+2Gs8R/IgPDZzUOzrAmSd
AYBJpEjaLra0aXiXhcPMPFkgtTfJCCdGSIrz4sho00QqqsJJ0NdkfChTRSj18FsK
3+jqJgOFA9HLFY5+q5tH+/RYbQRxqob49bE5f3XC/VV971wxIYnYywKYJtXnoT/x
8wvTHeU+xzjRMicqhJQCzkk5tgVC1MpoNn1qvdXgCZGv1SPCn1gbIkcE4H+poP5s
rmqbc5d9Mfg5h612N8z7gYdGQYh50QQL8QTpqo5HlsFv9yNT3VrRRh2Zj3/x2NGC
39hbc+QGyEcLmET/zbKFvK2APNkrfOdRJGOAfRdg4yY59IGgR7LMKp+7V9SqOxDF
Zr3p8z/awzLPAnsUxuLtTvL8O6ZVKrboL6HH48GtKeEGkrsYMznuTYuuQlVpE/Ww
zgIALgjsYxXBJD1yPIKFM0Ux2CTT7JqmXz5lWg29qzZmwtKtLR8robxiN98dPDSQ
oX2+Vcx1DiL4fYFX+l4+YaU/weG3bU+zu+tpewAODVQ77QaCGtd2Pkb6wnhV2Wjy
18IndjNN9FJrsNdjcfOOpGOdQfHt2WFEdNrZxVBSfuE2fyn7QCXN2tbvcAkLHIYT
sx+74EvpjTyH5MQqhWGeJqjxF9NhQFyH3cR9epD87MX4BdqNUax2rm2muNpt2umO
+07voCFoiY8e3XW85jfTgSfX7wjsMkH4MlkUVq+iWWqeNb3gNcy1bvL9M4XLyhlM
kAHB5zkaHIQQijXvCGQxqvQ3dk7TQtjlkxoT+1/DsDYN4/l/vFi2NG5Bvygtgx9Y
ky91298jBrZ67vU8YUIHnvGAvzLH6rtfo6V/Y5+Gg8YCfy5YiJrdHGYSggnHEuWv
xUjtMPiJA5aDzSg/pfwrYxuU67YEeld2DZ9lj8CFYtj3u0ggHothPX+wFKd6PshE
LzHV90zpNEWHjCKuQjRb3l/7Fs4rB35mzoNnatKWHA4ak0mNKcsZ/HeLygkvYoAg
b6/gkEfra3ysPto+x7IjAXnsgGDmh29jiRIMe5zkqotnV2hui3SYlo8UyIUXA888
1LVXbZGpP/Wvoixon34p5u5rftGSRzHqWa8+ZV+0min4X2QuTTnQ0MYZkSMIoSsY
KFwTUCyPhJO5M85/j7+mjpAIRyitUTCsWo1c0wg3hLhzhq5wLQG2e6hcA2mCTXNe
Qhh2B5MN7jW0JE0EweaDN3HfPrU0bkMbZGCkmHpqGyqwVRoiEmNVrucWX11r1FpJ
GJRtnRZLBf+NAz7OmVaxUIs7RUqbt1+Z2EbSmDn2Zrua0zHmoP6ZhwFy1x4b13/g
nmcSGTwgti0eVsr7Fe6lVeOCK5cIJq7lH5x8nNslJckmOYFANMNFghtHhi0xT+g4
4YaPMDsa2D9VFwaLpziw5fiU5wPOqNc9as/c9ASBrsS1QISy9wEmXfUnxwGdImZg
FCIb1n67kNoHzCokDaDXzxvsDd+ncSE07ufal6uobX9FTDI0RI6KTE1eLlQKcW8L
WWa+DdbcLagTQbUCPiPQhrW3sOKLf17S4PHj+L/GKDntwmett0aTJl/6qDEfnIEX
UaJZLSY0euKq9UAzMCNiA1c0z3OLamchHKoHa5hA4P7PFfR6HrMA8OFV3oDPGpq5
le4IJOIRt0rHg5oTEv8h963vcslbHcd/14IFyr1BxijE688NgLuqpAl1UEURDX7h
hVZWl54dXl9U0HbG8koWiKYd3bNY8HdgpTNBkAVOvH4Uyi6Z9kqay4JZxJxOrlys
C9qixMjID7x/nG6ze8arIwQo0Yjrn8BXHkJyE8xvIKI4ijwierpd0D3B5a2+u4mU
BL4wiYSDAGjQCyOPo1s0eiZgVXZUsEAl7XVQBHTxHBYVjW5P2K7p1k95GuEfLj45
ObAXGHGXnY6oR/IfQe2QWlbOHgFEfIQrPgtKm7+m8sTLBv1YKFPbpxMX4t4ElpxK
OGbi+l09EUK+bTll7n6PMot0Y6nnpMZZo2F0qFeyDC8DCltuWJfJWmVET40k9f4e
hzWZU8U2gkAHntkkqmF9kAYjFRCZfN+sQmuZdWSlN941Cg1rILtqjAR2TNuNt18E
JWxmN/OeJ7s68BzPVfgws+ma/kjg3VHcykqE7URBAsICk4Q1DwmTvkx+N5AB2gIR
UsugC01QjcgrcUCRPodNkIrVoLlt6LxN+peWrA5k4+dLDcP9HeGFhAuo8/ayACX4
z67WMnWhV3qdy9IjAro5K8DDDF0L6ts4Z26nY4iVbOepudmzDrZsKasiM8rKM7jY
7XWdovq/I14y21RlBy3XuSJdDrFjX3weFzKE57suP1ReOMnE8Ubkx/f0geGVZWe1
SkZBjF7I0FykOUSGSuiOIUXek04u9cBs2Xqr9Dg/t5gtSt816k2aAWJM5h9L92So
BM2glVe7ec8wZ41x2+WmNPRw94DrLqQOggyCwX92CqGHAVuEUhsfcz0cok+eM2Gr
oH3xmEygqtwrrzWArydK1u6dnPgtslRIjYam4qyp58IkIR/JkzeKxK5xguc+WsTb
fGzLGKOvxJcd+0rexuMMKt4yDzUrGAe2yYbD9bCAD1jpITdFK1LX/3fausqYDFpo
cCKiLtDMOeVvbhiV2TQOTIAslTTGaeJA/kwdqy7+mBdNjJk3+2AX183xGlCdn5/A
01pktiQd4krzVOb5bO1X0SAxTrmzi2rAiZxMKe9Y4QxYNNK8AcLFts6qypd1sZZi
75TDyEaOvf3iFI7mRcjgR/ILBeQeF7zxIDNdqesDRDH5I71BPItKkQLkn96UN67Y
2N9Ayjy1D5OrNhzcvCmw0djVDesrUM/Oz1aOzx1PsSgp8Np+VIU631ibxasHJwsR
sI8vABe6/YTJZa9iNtMgcJF+8nbXLq+TQMNGae8xhoYAGquS2qV+BJ2SDgYlVanM
qauWlUxilcsdwYFH0VxNv3q2NYghKeErVVWJtkz0+H1+wqdo9FKmAGKPyR/tshEg
glGsjX3q2THQKS0hpt00XCeOb7+5TjUmTfRcrNPluPUNnkFd4oYyS9EpjzfA1+OU
An6WEQlNEoPgwhWoOspJlukmPyMcQQLFiNM+XxSfu5j8KZuVA5P+8E/cKtsgvsGQ
ezNdcdKd4qVygHY/EgZ+zCwQKUS56b79Q2wVbyg9xtOTne6iSW+6m1PQsqHHLL+s
ME9Lb6yhF20KN5+ViXTcBws2AkT2khkrIUMEhxUkf3/XZOZ8xtqpNJTHfzpFtVYr
dbpxBcvDAvz5DKpYwCWPUQKr6awm4N+OK9hq5JLkFyNQgk9GZhlcFVz/98nH8nUk
g0ADlo/0b49mb1Mb2hihPq+8pLxpucIETQOnNrMnT/j54rEHWC5h9D3M2FPW1+QJ
+UgSPiplBAypToueXP6WKZW5ZYRixIDHl/FtMj3oGcVnWBUqVJVA2aA8/qGjCpVz
VuFdeil5IeZDsuy+LtZCLfbLlN+xP4v8Tp0PP/wpliXwhamcS04k8Nr5LtDyltVv
Dm0MTKPiVTAfeUwHbMRzE63AZj+U/hGkuzS651fn8B81pAcxr1ndQX14Ld70G8wq
M9c9dPFT5DfVcHH+nFraZZycpgMj0yfiRJjecMAoqI4PdyHElg6fFuLjOVkzt/kL
nEy99GsawLPgiWAZYSEUr50ULlEExcb7Bc6RDpoLPra647C9f6Ei0sKCl/JWVQsW
w3CuDnSVzQeFT7T7YPPyLbTqUWcWqg97r3bCWmrLRG+hisD40FBaGRl69qvv0R/4
kyP2w1BDSbfiqAAS9GeEyRWM3XvH9e4AxCq0pxnEElt498p25vRkutI2hMBF5lQw
xtJ2Odt3ovs+4GrfvuvokqIHE9kf/d0dzDR7rSSmr5KIlEublAoqpaMIMDpo940F
wEee8rOZMeYxVCQUWKhCXXi/yIE9cuGmdSN6BMJwHU4uGqzeuVOwTAF4vPWjlKdy
WtDssa2LMPeTxEltiI6SCvgB3SdcyGyGD9BQJ+fVfyyhu0Zf6sriF3k8rGsfYX2M
zII6k1NPdef96aVPLMIbXi30Egd/GCaBbc3Gc81ZXI+Gj+x/7ZpZoCgrT0Mj90zx
k48vCmo2wQA8A6pymxIlzZiSQjQv32e4WuMcb5EJNK28V2AAhset2mG+4xFeyZFr
mb1Ua7N9BKZ489TcfF+sQsFgjTh3oEd+8x5SBvfRQVVF13sP7LwusZHsr+c+0I4J
aGzamV6P9A/QD8Kh+okMooeyD6VkpRNr3h+jxuZT6HUoRRgoRn4G3pg58hb44i8h
0BD0e5c9gFn5PZg6gVHz+Y+dPBHMDiaizwqgwuajtf1dE9W1Njg62iX9CHuKfQEI
uCOXamrsV7Hs6AovNzJzzHLVckZaBE9TIaO1FPIH5wIP8Lbmf2sTCsmV1gkjvjOS
6rLzZV/M5Vc2UY32ern/oav/op/7lFP3yTAv90NMmBuRK6EVu3OR+4LWU74if8hR
7Z26R+igiLMx5wAuvaVYZzMPTqInrZGQJz/UP5WvOuDvFq68oxgZw9WfltfYp+Dr
pSDKNjgjmUV4aZNfsUMnqBL62tmadC+DlXGG8DCLejFIXOMdivsGvLnfI49K63F5
wGhuWFwCAlf6LNjc4P7oWmslF/qzAPDAFuYMiEpMRk+4bZHO6U0I6QkUcLS0hBZZ
Jndrhku0ol1ojXE6LT/+wBqQnl4L3SMmWokFnbGYPTAU5d4yXiThDzslmOdwkbGm
yVmpNFpIHwSpZZVR6P2tRPQTTk+PP0RSIXdhN1AJ9A/OCk3Me8VDkn0KpQijbv/e
Yx196ysIxji+PkCnzGLK1IvW2JYcZDxxoxJrfnsqMTubHBPj4KC/cBHOGaOvTOYI
16anWpZhoiFAOGREyGuDA6KpLV54QJXxhvwh54g+kacGZMjAQnTVVKWGe9OqNDXV
jXgHUr8WC/PXWqPKQ0YQDXaNtJBY7+XtvQt2LsunT4M6A0cD5p4/q+/V2nnDnZ6Q
iIOXEHnxa7EU6n6Qy6xTMW58/7JsA8+Qt8TeDSuGogV+FsOO7Y7rdMbm2aCMJfbK
GBHeaoAIBXUpuWafbr84RtTb3bXrU9ks0tou7AdNpOuqHhtOvbmVm96QR3lmZRGA
vLvlmWK80C5dEl16v1vwZ87f7pH+sIc4cWqjyyfNkJnfivDUx6i6rfh/mNp4wcZD
90VWatM66gF4BJprASVu25/tcAKeKerOfVmJ3AfJ3Rj4KDTUveWvofDLVQGyPbta
BsSV0SSmRfghaXHMQryn7vjeF2AETjqncxEH71NGMQV/7O64ByLt7EWtMGWPMDDy
ZEgu8L6FvWg8JIGpNFZhfOQa+9SkPWJwA06oP/ocLjZ0nN7DMdfKX1Q2q/4cAe9C
Wl+Fcfx0pV6k70h+yvhkVsapRFWNe4EfhpLs1HCFKs/X0vxHKJ+GeA0LPKvywYSx
4+yebN7Hoh9OVKGqqAUoRQlJ1aRFXuqjeY8YTEYk3YRgkZBcecT4hW5rdq3BXi7D
Cm7P5wPWi3Wy6cJSDfAn/3vfF5VFdTh2WnskNWWpvIAmFOAHrbdbZZW4AQxKbb/R
mf6BtRRhJ5D0donrmTjRdPRqAwPvWCSRgJFp7i6VaVr3Z7jFl4JNOoXSJFFX4UXY
4wvQHK3q/7MS/D8xam3e7KaqdCEWmjk2srXa9EzNlotr6OZPD8XFQVl3ML+J696X
2DVTsM2o3Hk0DlVAD6u8FcFyH9VIlj7jypBW1kkiguvhecbY44wDq+hX9PRNBwxL
lNiJnasPcVN20cNoHp1/ipH/KT4zO9x2welWEbO8lgmpF4SxQzDDkUKbRarUJRtN
mVMuNg5LE58CttZLEJAj5WAskCLRHlG3n8ZHCLn3GF+Bubh2h47Q49dtRLyg0FRw
T7CcLbDLr33rRUFZ2Werj29IgXXP9F5zV0Wnc0/u+A9HjJuAb5sth4QXXEGXUr1N
DV7ggo08jY7XP2XaKN0JXpKFl+QDhQRlfIrQdISR7CnHUgGOnmcfP48kczc25L31
gkU4KV5l4k4eqdvtBSX7ZsQ96VTd+a+V+Pdxsw0FJPeEqMRzPmugJqUsxwdp/nO1
bj9Ip0xFLqS/ITLjx4U/WT5FQBwHdQdPwb0iAHY8IHLnFgMugxc9k+KI7ghwSvTl
O9wl0M3ULvqdsRflQFx40FFy9Aa7WH674UAl+qs97B8Z3u4J0Amyt2+9QrlGldNp
HNiNoC50bLwfaijK71P23N45hxshO3To4i3iSyEL1FQhmu4gc8HxoVdKzX1k2jKt
8vCm+D72s5PSOpt+nVr6Fi3L47zOMo1rSg7OBTKT7kF/QNz2JX/AUQZmCXjD68yy
TrGEvU/QYXdwSNN/6ucpLYDj/9RIvmRu0M0LsGrAFmn/tlcbGxBdyApwxMWq7PlE
7v14lir6Wzef2pV+3nZP9cw5TJJdgRY2Xrgl4VEVgymeye+ScY3WF3C4JSgAE0M2
F57az5QjHBHfpjoYiwJzi8x/QjHcSQgWSMOIBMwZWLygSrRCAlLfVqd2ireNHxd2
6zg6LAn2h/ukmNwIlSDgQGb36WP1QIHFvBT0bqinn5AFZ+YNrgzDE6AXF9x4efT0
tGZued2wRK/6e62BIA/SUQ5fQ2WJL/8gjxVSDSR2jKt+NZCI9YYw9QvyUxHRWH3x
qRRmVayJ58ZVLqfdLubg57QDJb4r6CrlJzJOC4BumzdNwY1bLMwMavTI4tCeybs+
ybR9f21/Qez1NjJ0MDrU0bFaU+dXfcJ1zD1u2zZaBpcXs+d6kzRPJsjUmuaZ6hkX
XSJ6XJY99i2DbmHLIwvM49K3B3cIARNmjGm/xrKTRlMl++mqhkW2jiaJK5PgxYHx
DNa7GS4zb2z7CFk5DzRIiOBd1JaxWkBz1HuKLJ2iegdJdtRljRGDW5i1VjwtW4Sr
txTraijjodjHUKTdM3D0cFMQLGmx57UrZrGnDOLNQ699qh5aAjv8o28ONZ2ZJVzG
GlTkQ6TFPNI/PsfTAIRk8hpdnEXJGnTAgo1GreK87DfyzehhMo09wd7FHiOJdsIj
rOSZt3cta9mIrNMQkVaVK+tK12w7Pc1AveESyn867G88MHeq0V+kt66x7IEULwPD
6MWAc2MYEEZDgbjVpb3sHqRXy14m+eysqJm7ATmff9g6yU2bEwDWICuXesYzM8pp
P/UPtcCaDzwLsOxSMSOV8kWDyUUFFL0asOPLls5HNqycdRK3i+JHvsFHYDWE5wOr
HEBWWquPp7CjvYno7l1vkM+B6m0h3S9p6i3/pI7a0MR545cJ7DqvT7q7XRhnqOFk
j8ctWt9MkEo1uimFp14/TeraMTnXQefRkiFez0phOzKzP2/SZc3KHnjvlplgr2pU
FnjvIYVFRQ9FIWG/hC7z5ZeEytWAbrqfaRsQS8IdyI4xiWkBxvYSFLfX9JgAygAk
wbVXSBlYjEVqH7/sHucZc9NdIKgmL+Z1sWy/g2gnEXy9vwhzWQt0gbOSRtyS+qaP
HQ0Ifyx9EIvgy3y6VLcLbjonViQhPc8+2iLiaaMIyiOoTv9rniUydadbkRan3MDm
3Y23Z/kDZ8eWukf2gZSIBb3iq7KuwtNjmdX3/JYL0Mlpmiy+qsTMFH/XzCMQJJ5g
GfYWT+O+yHfVoJSnTIYPppXd7LDWnvvL21KaId9oAIjk1Q5QyWbtgtXo0IT1NYRl
0BDQlyewi5NxjteEt8bffCtnB83mQ5eC5h5MdMbPgcz/jQB1tLRZwa7DHYXsJ8fB
Vv+F9L3p6qoh1aKh3Dgtr2A/hv4Ik3ms/eRhIoZ6zLS62/NSU3JjiwL+4OIZJmE5
PLzKDuXDKWqc2X2vkIx3Muq4z73BUsPhc0Z418QbmOFQFcXEqBZR8EIoFfQaWovs
Pi1lUcfvxQ/lc9d4VnqVDJ2vTYgiH8XDdpxYvwIME7HgiLXAIUz1ru3Pdga9+vau
ua+e5F945rIGD75ppeeaGVyBdO8bWMn4T70t9zGhdokgo+UJy/vFHxWPO5tAGPIP
5pcFSknLl3KmMNBcTiVx7HKGgv/aCsYhevWMfuQv2itwXMe+tSbG3fnRBaCDjdPS
XlHHr7WGRG/S+vJiABhE7etsdBoXgD4GsCqTNqGS03mptEP0t+FD+ipPB8LZpPUR
iRUypvkXtQ3x6E+o/+NEyvhlGEEYqhllNPR8UaQFjNqROu5LdAYrUOLywt6BZFMw
z3Z+BGTILAYvvI4sT1zL9vJjlGcAlcURkPvs3ruhW1gG9dV2NxBIY2L5k55pW0Vn
7YG3dbpqc/gsI56+wYSVDS7AqtPGEimN7vgi5MKEY8UhhBWr1hU4pDS0hRWMEgS8
Nt6vczE+717tjpeMnBsxrCLq51dDPWhg9ynzbk+2BQAF5tr+VhReJXBdGeMcS8JB
8x6DO0VdeEBZjild7Xog7bkcomLQ1ir7g3wjC2OPW7sy40kmmqUJrDMgGt6w4XEL
BWgUlA7CsYU7mqgLPrbr3xEas6Q1RO7ZVDAuN3WhZv2XgO7iVri8Q1qor46LwByk
rlN+SJA/e5VevVsUnMb7Mc0fEcui8I3zq/lgHvT97Y7+eaBs2UxmdLEKEFXdcAcP
JOw0J8YcR7GFdtJnYoAO3/gMgZq0asfYDQVGuCGMGyJX5H935Cc86VGMIUE3tXeK
gpPlg+BeBSefez5grRz+xGf1bRf5uLuL9kdxW3RivAAn+W3H6Ya47iMNX3IOG5kD
oubK4tFX7NZpdcmmG2WePcTUtZx7kZ0uTR6ReEu3d/bdZoaIenHc8aPtCl6NvYvB
x43NE9+T4yiVK/0ieqAhRJFoi3HLLeMqV1myZfMmp/6Q67oIZqq3tWk2QNfofst5
tHtF6We+lfWoOluNPI0yGtfMbcgdCIUvvpxZXJVu2zlr7ppJnZEzM+zRO3c2uDw0
mBNINcTMgQ5W5YBeDuEFOKcgIWoGcz/KE0w+nJRz4eQ3IRS4FH0yREnc3wlNLncU
GI0I4tqiFc1/HcTE6T3TP+oFHutJ6e59XgNLu85+nbEaXRNazAIQlteudZThJ58V
MJSG/9bIHjv2WKSF9M/8o7DpZBWcoYYt2bWFwff8eE+CaqiDhz9nOvpkiq5scxK2
lz8M0ZAlfyi0AdRVqQqb+pek3FwzwS3eXFABz05pAUB8AlozR1ZWyBmhHrOb62zM
QhPIvKAjrU7desgj3JJra8MOk0IjGvhaZFKsB6lcoiO/pKvLGhm5nhAoG18wXNP9
HlNEkI78vgT3UqN6v54YFdJpQZUYLaLLA5dkQ56FxUAcvaK8ttheNghjSKUQDEAF
PJAFgmgh4urN0KrDEqbBO1cRueXas9ArZvJd/qCL9204nbnhasX/uMR6Stfb2eB/
PibQttjQDrg5YbzZAEVIHFZmWSh1KJ1oXTvFQ25dsEloWNOH52fLHGCKAQyuT10p
KDzWO69GR+x7d94L4Lp8ViPRH11SL5QKZj4ABhQ+8iqZihpE+t8TQ6VZKqjsmAL4
ae/w4ktU8HXgcFoXbNUrodoBOaoFDuicwZvIXWdS5mLWivVDCOqxKWcezeN1nkIg
Rn5qwf7FaV8jX0aptKy2QNJMOO5lVPV5jik/hP8JSFNyGoXAV7biAET1IqLaeRrR
4y1YM9fI+qtnRm4B5jkuV8SWut4LMRVNNDtQhkIO7m2R1OYV7BQcmUnjyF4BZrYm
9f3ksFaCLZmfd7sJxCtXkt/7gAGNpHlYDv4E2/PUB9ZPEUhv7wZrCjWEl5OOpKYY
NGDWoFBYZDt9LJivN1I7/DUImRP+9nsAavGaGrvFvdxocZoEOZCmtzcHCk8lrrNr
WYoDa7e/8lYTItjTm9Xyy7iJ+ZkKeAB+puyBWoIniUoNIZhsNQg3UTQtwYNSmBnf
2Z8nANC0os99I5GG82lyDLgC4ibp+Ox6acyZQMDY4PuE+l+A1gLcI/8v5RvAn+A8
rQ5eIN3QwfYtHMgSEAnK7mme3ebpdIi6iVrOtH/sfnrA3ZtbGfsCTyeb+6YHUHzD
nFozPa4BPpaqMWj0QOpnXbGoZGL6NZuZWCfQomy0DLUbdUk4f2hWxYXBEiHLH/cA
a515Cbu0uqyvnnFAkJkIzPwx8vadO//jytdoeMsgZkOBoTjrmgayNtde7crjvd/J
pgs6/yYBCtxjwVQycTX4ft7I2ztZWObJa+dhvBySepi1IrGdLSyBYS+skzzVDDDk
h6lqOn0VJhTd/Mf9OQ6vKFKMLqYRuGiKnvpP5wGRmVNOrwWD3vrx/tb26/ZSU7/J
4DcKDJSxc8sQc/ONlW+onPBJjNmvQ6+mCV2/LK2216VJbagCHEzwJqVhh9E3//gp
5sgpnHQmSwlxxC+J4BrHg7ZdzT4EWSopgpR89K2IwYOhGJ9Twjt675XOoa+8HDzx
CFI+mJUx4bJeaqbFTJGicrAzIsvbKDpLIueysSl9Hg5dxQOqRvSNzm8UWwSZVAGy
vw/ohgUeYMUR/HAtwOcwgQiBpRbMb3jXt2ik6EQyfCVV/LZ5rkDJe+I/fPqgrnig
xGGGnkrOiQYQ0gCM9MCE58K+vKLoitpunvh/e5ohs24BKxMGlqMZtGhk/wxUAp7F
6KGZ7k1/0IAAfqEH55ueR5YD3l6DKUDiLxgQLHiH18NFI/SKiMEmbYkuYST8Pi5R
axuAzLKe8PbqwRi+0DJucrcFBUeKYxEtEAMrBtctSBDZAnn7dGvdNOjF29MySWhG
/YrjDaVu71dnn4FzrWrc8sTIUk5FJUOSIdio5/qwLACH1lh1joKQCjy51J6aC16j
qFC8UPSkk5BU3haNDz1j1L+GhlhjVjKvoB+GnksODIk5STUswb2PGP/n73BvTfvD
lI2dwvTJp3qHopRVDT8CQWxwFfiinbppoLpKzFYYaqb1ubMf8itpfWS7DIaqgqZc
Hts73xMw6YgqZr3vXH38mbhdQ4l9YLVJOIo24vE+jjdUJmil1WM20nZ91FyUVX3E
l75QXJ1ZjniKGcP9McTfGOfJfl5B89FHT6jgJAtwkIgX5sf9CvWat/ug+VpqHf5g
mjIQTazG60N7B4P97LXwKdcvl3ycQondMXMOqCJsGWgrUirD6b3VOTwqLnPeYmTh
efqp3zoB3MSp4LvFB2xchkdBMVl8QSJYnc/NCP2Q7xwLh9sLmJf8nTwpl1NK0eKf
c43OWhnvf2i8vC3wwO8jK3OqPWG9QaZ9c9jwBTCicERdTtcpqFvgm+stoQ9SjiFg
y6ScWEUCk857fuondBgt4Ply7tjKCZTZh8eEkfK2jzKEolhCuPvIlv3cPdl8gmoN
E/y/DQb8mnk02Nscr6AbEV+bzjqnFwROo49OrTi/+EpBiWm8R73wJpyXCDVBSbV4
u8qePh1PTC+PGQnexFx0sEddkRgPUPMbml0dcKOykCwa5xjqvFSygLRRa1vMysrK
5C2AFcXs8uQRH2owQrQWZea2UilomhyoKxWL8um2UIt6E3ySGgnQzu7pVWaaIYx5
yM3DanbpmSGgZGHTme1ljHjZe+jrO5cnwd5YIZ0yU87I5GdQVN4eZzYxL6A0lY0k
BuRX9EKZ81t7QoqmMImR0bGFhIirj76xu2eiK+XoGWLhuf9F0acpJFR6wPEQWmaZ
htYCUDjA3Rz0yFCRRRpJet72DRZTyO4fPewK75o19vf31eTT8gt6UR8JEfZgrWq6
H6KP/81TejNlpHepX3KTLzTnt6dkqBSHWTHzTOdR+fZ/EEXCBG4KO4k16eOg7C19
tCAIHhgxlEPPHtA/Us6d52zx6hiwrrByOI4mjx0uYQc4BiyN4z7U8weTP7fYFJaD
MHWLJ5qFSbXKuulQ/CINPwr7tsGTifBwXU85eAWJOV8XF/6CFQ60FxgErTneYhwg
kT7wVl2ldhz4DYS2lRo+yE1Jo7TuVc9oQH2lRIXkDZIG2I4NPPq4fqgy5bv10qup
aC8rjXJVKbAXfyEdz9IdI62zvrIInT4lDQ8kx4EhsO6TylnHn17lJPGDFbH9voO7
s05Ygt21yaPNYa4Ubn8+vhcJnCTk+8dwREDuWSoJCyEKDfGy5cEICNaoytW5p1za
wkuWqv07gz8ob2udx5CmPvF/O19mwX4pc/U0kyvh3CGFSWtXNoF8aQzEj7cNECpH
+EmOhEFLoAYmu/lFkn4BqznY3ez6p+yjhShUfaMnNuhu8WIPr2x8FlQKRf/jKi57
swVOqcPXQpuF0/RgZX/Mlz8SrasxjF1YLp5aHs7atQ4gj9rpAcBalBQVoZ9Tj3G8
JNHuKgEUEWmZqwVINtN2TpGuw3mtwxYPg1udbfXLL77VtQn7+nAIH3AQ6kXqSfP1
RSBT0r2MjIOhQWV4A9c4fSGVXsn/NgtmkJcoHf90rMUFrmmKwN6qKCUSkJUlnRsk
flAAvkrSr7yZfg1q9WjPnPbcwtfnSE6CZ9pvEwfOe6kyxlVSBmQ8Cgz0bY7feREi
HdTr5zxkYDkOUO1lMiEIxTreTVqmJsCTZr4QnXc4E6qjvFlgUoBcZbHyRdAXGUU+
cWFuCtlx0K/9Jf3HIZh2JqTxCROTJJQ63zjtkkSUKO/al/hp07mOVmvpY5zHqrpZ
X5MYw3U5WghHFxJ1XlTD+J5h+tO6rQOLOdEr/vmxEFdBvwU0Lev04cLHxVyZ/7nB
5qFyoZxIXCk73CEBT25267pUYqx7rrzaF1Bqs8lekxpgdXWzp++9i7xos+Ha9KoT
qAYWoPjAnxs0brRDv+p1pQ13agnMmZ2nN0ReHropIYNMfg5ZYEKChoftECAiqtvh
nJTuRyARGZp7Ss7/7yJ1R5tMsmIHAaX3TK9E9Q0YZWwkHzznQg24SDUT1TrYHYP8
6akiI8LY+zRP25v5r/+BOGXo2caAvL2PB/9THFXnRa3iQEJ67SFZlxigFvYli2Op
xiC63AtlmVB4SQCSkWeHLFgaaQeYCyedF6D6dRMrOKHM2XpQovqNTmr4Ee9GoLKJ
DWWSsLlvQm6VHbp3LMvq8e+IY1J8cmMfHwst91gJsKUBKK4hfGe7S8NAf6Y1Ne4h
B5GQuIbQYk46RlXK8LztbCi+ndiLG6Nani8E/TAAvd6uQD9/CxTVUZ23PM0cQtq2
UFpQWhix0EmJFqMc/jtoRTjqey5lv0TLsaxU0mStQ6cGOpIwQvGrQi2lhGBg+2ep
G0YnNxDIz/rHOBXlVAlHN2ADx3plt+r0oFhwghs0v1tts0j/xoTLVFINqzFDXSxs
onXqskw2ntCDMhJtzKB+VW7f7J54yBpruhz8p+zrKlwgw3vFZwmIMviz9OrR2Jnj
l5i2VLG8TYUY33uJrvDatrIgIi0MtfEkCN5MZQLf+BuC34Ld6sesYC4YorXag3iW
90FFNwO2mTNcmL1y+KaV4Z5jOSbnxw5vb/BsBnHjp+4naE91lT7IeS5CJg1iR6md
p0jjLuOYF0Jdja2W7NgTV3TceXOBYS0JBNHYx1ryWKSGXXRFaDV4R3grQDTVjMly
du/nQU95rrOnarRaHM/oixeCxQY/tWOalpoyNEP7hwUugMZjzc+AK7DkKCsLTls9
ZcAD1U2TV4RecxhlOvaCLDxmn2nLOV29BSuHSqvgf5C4KgX//2ppsZA52dH4MFXY
6L3r3UBWUSYlE1ZrKrYXb+8Fbc6YUXRoFNLms0YSW8aDAdEX9zzRS6uNH0c0LSqM
N/zxdIS0CCc9lVbGjZFPFFTTHKGqkwZde3li4QDgNjdxNEPeIbsk5xCtFgHNSiJt
t15vygBuxwZcWzJwDt7IPUOaqeZ6QBkmzJzGV6qsszGT4ZBfa+FWOp2JZTYvxeJ3
SJaQyVjuzQ3LcOumYpB8ag7GRsFGzKdeZCVW72d15sv1Qd18mHfycc18fxht+sEK
idqnOZm6Cy0IO3WkvgTJiKImRD45GHh436tS600MZxzd9f/BZByaH8wpSZAXgRzG
nuMZY92E3lhl86pJAn9qi5inK2u9Zn+vW1oooUifa3LXcqrqqIZnuxomqpv6hEd8
J6NKi0yzGW5DIYtdsFUg3bRWUQK/D2EuFGyiPVgiS85oJnRJbJ1eOXJABC8AaQIg
Rh917wZWDwupCTLk9PFSCdS1ozGitflrfpO9WBCkJt6dkvrXAocXS+hLOPHGV3os
HZpxeGDQMR8fXXTwu3YWbfwUE4GeFJ7Pw1grRGKsBX2qMCDRj4MPczH/X1CDwrgj
3kj22IimzzE3fzpJpA/sfOcIjw6DE58ppFzBgN5Hq7nxIWiMUdMvDiQ2qymQcbia
SSrq2xNVGIdfie8LeCeqt31mom5Omz1QozEA38KOKEyvkbyutEA5GZrrL4rs+4u0
Q9K9wsDumGdzL9LpD0lrAF7tONlqFLdccET+pk96ON8FpPn1/qyv5Xrn/7m7bN7C
FVQl2M0JZu5qZolHIEQ0E8NqZYWYJPePlNU4Jb1y7qqw7RqYoxdzitz0obZsPYCj
9mSA5xmPGbq85uoJDZt+DhBNm/hErNXTrJpCkArRAXivyaKu7NcFH9f3SGXa+zkg
K8imHCQy1ZdAmnpxm03yLunvgdawSlyPTu3Hag61BE9uVFKDYxyUmknI72earK4g
Ztka26e1iTkRJ4oSPMATTad2JSk6YCMSAMcscMOWYn7nBHKYbAh5K5km5oTvimhl
bOpEuDLG8WLODGN+fJg/EB/5WHWSB02nP4C73PozIpGFSJRu8y+tgfSYZ5wg5u0w
6lfbwB4EGtA+7EWaFJA6Qlj+jNxx6MqsC7ibZwqX5ibYEDuLlk0+cJaOBPozIQPK
gpq2cYQlVBRB3mKy+oaSX349aptX0J2SEN+TjFpPffYYYNLWb1M97AgB5Nnshkge
6HGVQMaVFoHyyF6nBTYhjTMPz7FkETQPdI8PFjZ6GH+/5cnWzRsNvmQl+KkLThcV
GJJbdj7aED+xsYjG4sG11mH9hz5jdRV84xJxb8zLssILzFXtjkyRjKYtWNg464F2
fmrRneK7r7b3yiUruKJlH/LRKfcPWbPIsXbh9Z3auf3p83KXzpUw63b4G23STQa4
E9rfR4T1LbXioX/6h6X8ynyju8oEyZE3WpYBE3K6yYS9LyCRZdq+vnOolfeXPlgk
T7h1hnTdrmgqvpAT7sskUkPfBiV21BMTTv/q8bWgwh3/fhW9qsPk7m38TcgWxdrT
IYKvnikQKrYUoZhLrsMK7nyboODx36MpwyfgUl+t3JU82B2H6JMRjp/dHNIO8pUP
h6L9nBiZt8fABCGbjdmquVHOfoTKrnBYkFkHJoT2vGX84cTncoEEgxibCUG3iuvf
Zh4vwCdDwOoCQCEhACiDCo74326LuNbMa91SxSgb2PrP+F/FeYgmWfSZrDolvrGj
7H1a+dZmcmurS5Ik1tvPjca28//y9htxH4cvD0RgesWFMt581ysJE3Y9nNk537MF
Hfk2nGLNINO8tCfgzRJbPN3Ny8EzXPe0iCKoJfsp0sptu84Dn/5s4XVLpZT9jBwk
lM6r6SnJ/TDeePT+REQPGEGL7GNI8r5D0gtwMSw68O2FnCW0aCo2J9QZqpg9gZls
6j51O4FRgYtOFhQTAmqkpVclhF932TAkyd9D903GbbFEaA1i6fqfSSbWx9vlUaSD
SwPxJKOR19LbjaXiu6JHTmat2YCUreOL3P/nh+qBL3mlMYf0NlOowgrQAXOG4Lnn
6LWFHaUsDWAQ2KxB3CgCtMppzkZcmSbkGf8iDCOUKd0N985NKPFWOHZtNaerAwH3
6MRac4ZVNvOTw+XXF+iA0ANy3w60I8EjHeX8bECWnb6rBN3BlKr5+9Aaw1mjtoSD
le9+WR8rENjzRQtA2l7ABFPsWkZR7J9Qy8RMKudo/e03AHYNvUKAfzhPqE/fklBa
P0uf0t9z7RUclOGIpZJs8HhyGcVWJgGBxr7MTzvpDXnaBaEx0Qi3M7alejtI3H4X
2g32D8pLdpbILzw9nbZb5pgEwAU6F1jrhHljbgizB888Pg3DJRU/B9JCi31k7wI3
hzpACDYfqJCEAD2sp/W69Y1dZgqrV+WIYM6QF780fsashYNNCFvzyupgxuhSBfzb
gwatIUc1tBOfehLz9rbITkfQ8cF8MUHtEkhEl//j2OOrIKNogFCfnRs1E4il1rAM
N7M8Iz8hsfqiYNR42UqpF/ufAvNjFFuXSdB9XDV+dDxZQjK5FaT2BVQeob9/vZOe
TZLrWsHAZVwjv6YAPUD+amnGNz6XcGVpixWtXOTWiejHCYrVXP1Avh0fxxSXaD1k
Qltw4mXWdZHYBhWwW2FYKIzzDcrlzUV7S9HhH3Drt+9m0XMeiVo15qGWoPIcbFk9
id7b72dPRb6//2h6hnTfHkKwd7nIindNr7N18tJqsNQ=
--pragma protect end_data_block
--pragma protect digest_block
zKbFXWosOR+IxyYPBGnhalvV+Zw=
--pragma protect end_digest_block
--pragma protect end_protected
