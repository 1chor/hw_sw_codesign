-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
A2xVM6lUbsRlKEX5iXO2d2+bCQVi5r/Be+yCbKKcp6HprMjOQmw+rkftCBlLtzoB
4Nuwr7ExBmd47VNQjrI8WM0yIsnq8urQRRRrRmLFQctseZ9O/LVPT6i1cS2QI5im
fw8gIS182lmCyWJUrZATxb20KgXiOgCvZuv/UgGuZgI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5600)

`protect DATA_BLOCK
yVPSvlYX2R391fkuAyfBAsGz/+DcPRCwRWAhTPss0o1Xb3gQtD6VcJ24Ihi86jW0
DtPGhOrT8MssbbeKid5jWMG0nqHWnaKNEC1YYfpaprECxtdSAZfXYkCVY0AQkf5/
/nAv3J4shI54urC+NuwMNiOUaOlADNEIYQ5QBHYkNDoI62EaXwFRovscnQYhFZU5
gyJSlr2DY3SeXj+C5+ALAlE8iHo+k5xYb/2EXxN7Xx8Eh7v2TRupr1hwgn9xH9u5
ZXN7v5ZcEmMGv3ibwfQP7BH24G+aY3I8LKZoeaOh8LaB5kPBIqp95uC/8YrTuj8m
mOW0lpeb/FWBf8DhA9FWvQtlAosBvFG/MVr8oJ9B6atVfsct94mkOtBLoPZyuCUM
iF5akHATVrR3bAaPNfROyXu6lcsHW14PNddgTuOvewinZOMxOa2BO/itDsMuxgbQ
DJSktlHKGVcC7TEfjF874sUrCKNUiFl5oeirPm7K9xhcQ0pjJEgy+W9+pVLRmrMx
gQMDWjdRbHKfoTXybIMGZYh16qOUuO5F/hisOP3hyZ5497Z4ac6T8MMrrkVD2mRm
EgOVfAXYdg6SXcz6kxjb958RIcR2qY3r9AANZcAh4lSZzhZXSiOg7mUvtScXdeQ0
i/ibtGpy4KxiZeRepBRBtu/qRdE9a6UCuUev2seDE0oe7Fy8+t7CtrW4N9xMK7fK
W+euLgesxGsAVjCTy5r1dAHEMhePYlqaS49REcNIigf/UMsMvn3eKjK/+aPb65Gd
effQePCBJGP0AZ74FV7xltXdFXANrHhRpifKORCes4fsz/aiMaYPg8Bt+GFXd3sp
M4nS/7xpz+MXeJ2Ad7fR+i9892KDMOddGDzi8y8zNqHdJhFg9MD2W6EKktDeexRS
OIF7wZDLJ+Nyhr+dFhhNRkAQb8rrU11TTo0gUp1IBngiKCub1CMRe3Lc/CVoTpiO
ci8ijj2SKYK0tmzhbzRMi1uHFKr5QYRFavwp+wE4tpApeKrMhdDVULw+BAYnu2fB
IYmgZV5kc6CzL+6XWCSCw4YyVmS1FVhbifKl7mhBk4+6leeuJ6jhLb5fcC6GHqg3
Sp8uvb4+hJwzKpWniom3T364jJiZt6Gri5XlSQtWSPVonW3z4vhVCPKgxYkG7GBR
y9R6u+vml6WwrPlPHz/07aTlvWlhHw1DiQ4P9aYCJfL/D6um/NaOSJnFhAh6NUS6
Vv5qUfIbfFgabUVXa8s5qknSq3EFsFU7SUpe5pzR2jQhIGFEw6kDjeltYfnKcJlH
4orSxwXrilvwJWuBoK6A1C/q7mM2cml+6jllbP1s9NDWyAeh6E85uPv2yf17y/Lj
RVNltJoQXnZ59RmyVD8mxpSjx92HmpSDI1CW2qU4KrtzDf+xR4fXoWh+CmTSQqpN
YAv2gnMP8ndXTl5CJJfBW/8nCzo0YqyvtAjPyE//jXMuPDL31gPKE85mQI4pvjbV
vuZYSpa/G5KdTfMs3VfYB06QdKENiHsU7B/zh7KJvlDb7fbQduRnHFM+B6Bo5sEX
AGOxqsma8eC1R5bRZBwhydpzrRIZGF/NE19AIfexBW9igqxEFYHgCKlbbIqQIBL7
f7hT7Jj8Hkvz7EJkKelOOYOB2KUbR684QNXhiEhZoe3ufXMSz7umVRStsxJQjC/s
a+YXlGXWtPRA9llnlFe/sDi9U/h5zpDommWrtMCCCnnFBdzHxy42hG4+P0RJ8zMI
NJZKLbiskKBYYMTPsKR7XKiWWsG1q+Ek0AgUpNTMKBUDnPBa/bpxD1yWaCvjf2jy
nNSxOqLmrFru0cVmrQO3DMsEejNsZnsRMxiA5sYbUMa5UUXpr4lDZgoB5/tmzVMo
1pi5f2XlSIc/EXnxKUHcebIh81smVmLYxBypQyC3AHu6nlKRQEEo9zS/tQin5MML
+t7PONTXSODQh6Ayok55U6sNMLdyyORJquf+UA4MtD84V6jW0UN+anpKtq1yX+fh
rFvckAK404+mT/a0N3cYMxsAqqy3uOXp7PjmYPqhoe11Ts7upm/xhK8JRpU09knl
l3F9rfItZvLGt43x5NOseg1/4nI3DUXUZqKKVL7g4fGL48ZfUlOcdkVUr095InXA
VYmXbQ9DYc39Y2+L1w5tyCBnRVLzTjEE1yhp15t5Fd3fF827bfcFk1Q/R1EZ7z4U
m6pEXxcIYXEoiM/qGdksjfey4jfSpyMGNufpnnlNsHptlI2HuYc3hDdJJQBHAt7i
2v75svK3VyhcjlK0q++ZAFnItuiAEEKCrpL+OBvE4zKt5h1Q7TehFryjV6nwVu3B
O+g+MdhBeaT98yGIqOg6MH5UWPrk/lwWdogSJQv25yRVpHv+oc6IfZj6RE4ib129
qQ6hQZm3EPIPeUdN0YFEZpqU3WZwPqls37FPvUO9PLT4O8z+a/jQwrTEo0fhtxO5
ZpIjatxN7EEOvf5iqwEPRhEBz1A8O+eqRCR1PdPAuywh26gIhmbTYa3F3nbxu5/J
4K5AToomjxlATxwyko+3a8uv9vQ0md7gSENSUhCKR11KsX8uSJ0iWQE0GtGc+Umc
ixpd5mkfmoPqBbkiEIVCIEs8owDkVOqyfe83vmij7lT+AXSYRSjXAW9LiI0bLRyH
Fsq7qf7uzWvfil15lL+6JdurKoQB7PCw+W04JXVNhxQfBHv6BAAFREKqg1xB5W4W
JXY66w6Bi0gxBCUtNNHArHGknXK44Y0tBtN/73PVdrxp4coWcTXPOQX4U5TcOOHM
HMfwi0Q3feb/9mmLYVWjnCo2S77bwfd5kYOcO4kldYelW3IzY3c1Q9AVJ1b+3BsC
YAxeVy+bXG7PpNU9YKRoaCiyzg+bzz0R8Yz9dml8KUNfLys8fwRjQgPwfHPWBD1C
uo9D9Hq765IcK+l0LrcVVCP3Jl+YOtWxC0a8NaYlGaPSYOzSEK1oiOfJhN+BquXG
z1mqhdWhM/gJHRiPLByEtTnw2FCjz7SXYr2GVDqVu38oMLrKZjxmIu91JGFkWBR3
ZIckI/4YGlINgk8My/44yAHW3PdDYpv7IxnrWQvzwoVDLOicQtxx/CTLBP5YZhdQ
a6Lj69xIeOX8H2dfXjXH5ipSyabtHziknCT34XIqbb4xSgUpf6naGuII3eV6NsoA
8ZjmyRMzsRvcTTrC9DzJ9GBH9f4Yn1sgx5cyNde0dy561csdMqT6Cd6kIajVrHRh
1oAGjDsv9AMoVBmh2nW52wCyP5mJIecZpGtracaJb8dasCmwax2tVN6xrXHd7ZII
BAThKzuBCb7fVXSJ76LSdtgdnTLUFIaEaOk5RVvDho9d64Keh6i7+StxRWA+bvce
YqU7QwyWVn7T627gZhgM3X2ECT3VEKxg5qXNw39YVh2yhCChkq5xiHe5oor+GGl5
QijLUXvpNAFAnGFn1yTw3DZl7FtMbgFbDnLlEEggYnogckm5nuW24/Cxgz5tOLgH
UpLDMqIZZK19MOV8vH20OW2m//r6SjsnaaZ418jIlGIMQNenErJxIK7YqwJL8VOH
/wld5HuqY3u05yYPeEluj1NyDCX0/G5ek5gEMecjIYIRJpIr2dow02o+8Uv3JC8L
RpBrkVbn42nrexx09OywSZqHO229P+rddx88+por24+kKxSXuMMIV4+g3lKiV7AT
xCdZOSwURcaigDp25nZjxBlP7yC/2GHMUG910lGioaNyWvWcuKReMOy60NQ56y7q
sXgMagoufT0MZ/VryZsMtBAB5jcTcpyVoygyu7+/i4ho62TwQSXCN5M0t1io1FxM
1aURzIyjjt2BbeLDo/d8WwbyaRHhMMk4u9Slj1Kgk8nAA90BkniLzANlbrXBJE/o
SaRSE5FsqkK3QSSk8LrJxOIg0mqc2hjdWBHetyU29u0NGcVrVpVG4T3ajRT8NhIp
ytyRPITfO8PPun+zw/qc2OWZyqM+/RME4UOgB2mNvOWbBsYedtp4s6JvyrMJbWPu
W8E6N1wQAb8DMPyUOZYPRS20jLWZ62c+EYmPx2kmniNg6SQV3QJiQTYBVpQUxUnE
BLTIkmEu7uqa+ihTnWp8aprA9E3+9FFJCnyAFnx4LY9FBixGIVRiDIhiYO4SYVBK
+EyAaDVe74WSSGDbYbilw/lNCMvtb4rnVuB6rx7WDaURIe4ljWaOtL+bbS/4CPBI
beVHt5JLV33ByiB6+rglfRW9cr3wsV+S/QMo2mE1/pqCMUTXD/F6IwHFzO4vhFGb
EC2cfRHzl0qqAmYqr0JQvitp62C0fcpgkMTRMlMltlqIYlJPWilgADf6QzhqtJ+/
pEl8eJtIMmwc/RNpbewwG79EcHlFTwhULxxtEkB0sUE+boYNAM9OWPsk1ox/hDVA
rXnKDt6XM58OdjHShd2bR1K08fnEdZxJagGrT8rZWm0q1e485WpRrb5e07NDXVzd
Py0ryhoXr4/7T2W/goII9vHnOyF7ooHF47FMEt0AzFOvE5nbk5iZtUgaKBTYPDln
mHVihNSW9Nhy3WCqJx72puWXt8Gzz0GMwJ/xBXnUeOx4wYSI6S/X7uASLwTWT/dx
nwxxs2wgekGp5Xmc4o4k3t6E8xysWwEv647ojyHiG9u+LF5eq8rBkYLUlx81J0vb
JgAhFp9ERv8gu6XmMoSdxaVAO7wJMfbjqdi2cvuSWsTo6VA65Bkwgt4KsvGeg7mW
XsbnxHmyfM782fbrc9O9BazYABMEUdZi1LzVenDr1bytH8CYwleB9ffb7lEKsAwM
pELwQHC8DKgUkeoTEid1iRP1+Uiyt5gBlWvxVZY786TLrYvRbPL/QExzx4n2w/II
c2pHMP3vlHQdb6L9xtaxpSvyj+2S+C7c0abkonhZA0Gop9TvSW7g2kJmjpDT2XfF
5tqLcoph4VH6L4G1voXNksdmf0t2B70UxAICpt+IjUDfm4TY/aVpbChmyrnjbDJK
mC7p8/OrP0pfnniFjgJiOts9WZrD7cDvQYf2gomKYb1SYDSO1RZIhnIXCm0AKckE
4ISBK0qhj1FRtDiH3aQcjoFIEah6WJ4G+JhL79Cet7RLWXmEWGAjxF5hZHh8ZbIQ
j1uDW4Ve0UeOZ1MWM9eJw/Hb18UXCuZWGPH8+n1E7bpCwgm9XwvHGZb0QrXkzRFM
8zToo3xGBzSqdL/r6Yyqs/LXiyDZMZPhiMp4wXXn8B0hWXrUyMj3O4695AjSIUgt
VkJ++NlLGi+t4ZPUvpe5ZIxlH54Jw61D/mZWj6zxGeujYCq+xX9fPOMWYWpmNhaG
LxMLrk//z/WQEVQ2bzswOiSwpWlZuBjXNFnSsdNvK7ds7f9oky/g0LNL/qPJtcLt
U51M9vVxw+5ynNxHxNBeD4zTUhvzs8kAOTmI+L6CW4iUOWElXx3tlj7abQvtCk9c
KPsKjyI2W5nx3PDEWRb8k6IxxwRr7AWO+xPEePEN6fdF8Q1o33DzvPajRjwlnf6o
2RCSCpkcgZ+KOiY/17SDPJmBoYSC9FhUbjg3fMSFezq2o7J+63IJ78gjUVfpfo2w
4Tt8dNYweZhSL4wcg3GKwJfAGws823luKpoK1RpLru5S7eSUra5oCBDZicucQiDc
9rNUE3/33wH/W9KC89I/7+rlFqbgjqjdHoPZPcY46p0CRipNc5+nHAnEJuoS1x86
INv7vZG9ABGZpptZoY5HSeYPG9Di0Panb++oshj5njY0U/06GPe45yqL6DApZcnl
oy5wFJj5hQ0j/6bqGkiggQZXggXaI3ch/SANMx/J9yOl1+FpzAq5prd9NpHG5IXu
72DEI/TAiFi2k3MEp7OWeZWTRNRh8qr6VMsnuPeBfyDGVCZhOUnaHfcKFXWItrGN
srHYfjFsnU+7eAwyX+kMoEsR7lj8GC+9m8mmLqe0BjUeHAmb2fAj0xRTYq+9ua9U
/6gHWiE40KYB1dUeDZFWwQ1Ekp8VhTax8NrXfF80dvATSPBzh83JXNSySiWtE5CV
1PRVEJeAL3mm/GY1a/OTqiFK0BbM2yeLy+MYpmy8okQXtf1AJ19egJP3HeSgbRye
X9cLva2pmaBlJMaDIdy//mBKuVSNFsDDOL/lcN7D0iJT8kwXleQg799i/AzZqrKR
GTuZjZtOUiK0AC/hVwlal1+vvwU3DRt7Vv661/ExjdoIDHso6h8x57eyamL7S/Bb
N0s0XGQUxeZN3EkI8BglE1tPYAfZnlg+kj/e6Y2BTHw7nNzeStRZtjGYptITUlRd
XjbhhuhBdRrbEGUqInv/eFwW9RANcNqxwjP6uSIVaZfN9Rh5CWKnLTV6eMVs7SBz
9VJDqdb+UIkEyk7flB4lr/sUvHWEaLyzLkC6RkyoCdMxL6BO5RsWfiwrp1IIQwUB
h8i3MUzGluOGje/GMEsfgHNW11QAOrem/yAXCKkAF1Fo+bWpYva8LJ/jL+0wCkAW
DNjxwc/dHSrg924xRJOKe5sObPenRvTqCzg+p7LgNNisSQw3/6rulk/1l5ShtRmI
R4NwDseSBULnDuYM0q77g5LGSmGQJ/etmIfZlg4+8gsYjtQ1yAgAYgyciArLHEyH
KJyHgNqj2XrcbWYpcD3YCI9IFNc9+LIRB5sjCrwFkt6LikbEbJZ6oLQatp7E9NT/
KuK/cJuBj4YPyVdLd25ZkLGG1VwWReQZ0oHOrcO19pCnWeocPFMQGJChVG13cHiJ
kfng7bZU+vaSaym4kxCpv4Mv447MTuUY1G3AyBOSzN39zdQJWsGISl+9ykQQhT+7
SMuhPgkNYcreG57Qjs/N+Ayji/2D9xsFdiqRc0huId/JtUJMbBSr0Llr3uMPiSSI
P3eO+9HTkd6oQfPv6uNdMZM6wtk8BNvn7U7GGHnWrrIxq9Lxu+r2NQ8G+sUsEW38
tkWqk8ANSOggAyJwKjuv11hRCFG7LMUuT5F6t711/0bLQJhTKekQ2N+ZY3gfHDIq
qt37vmYHABk/Pit6Guw+fHjAA31o64NcaZYa2kyVuPy0rE7UDrVY7SAF1c4IxmIN
SJ1K20Rlw1kkTN8BZwPUmTJ45E7sPE08coe1agWLvpG+w+He0N+eIcdW4mlN4Ia4
WiQXwR/MbAn5D0952wzjCI8D/c7lz1KJCTofUnSMD1tq/kpc+mw758/6RFjPqOST
sIFpz+uua2W0fYFj51xJBIhEDRh1qP9R2/3Z8umJE9g02Nb2ElYGcB/4w4NRFzre
yVT/csoI7Gm3FRKr1MkxbeEnKqap4T4xHWxJxIrubSGIdtR1RUoopA0bRP+u0RnQ
nT6aa9CoQz2v8XEgA1bXbhjbflUe9J0LFVqJHlDf68RAIG9Ckqy6b7NouSTc/nMx
kepUSPEN9TzuKjBQ6uyM6HEFPFo9jVkRDIY0aWxADWFVpQS6VtuQlbaimgjR2LY5
q3o4wrf6fEx1oD69wlz+a2oGH+P8j9D9Ywhy+tTYGKuIE+mroBv78x3O+AYOXNWm
3SuHLeCJ3tKjNtMCdNBnoqTH3kdrYEBbQAXmFkR3aqRp71tF5u51Hf0lAsKTMWej
wUAu0Bi2gbbkIH9MvXrFew==
`protect END_PROTECTED