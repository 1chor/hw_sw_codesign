-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
n5oiBxUKCT7ys7juDkz+46bEqFp3738l1maPbyO6bkHOXCno8/Yb5RFUucfJEqMKRC7O/fkLcAU2
u7Wy3z0RJEFpjukkBt69lzdtckdS05TodAYB0JmisbXB5Ug03nxTWNDE6aCQUMN8dxf9/r4EgE0T
nLfSoBP7f6/9PDRi2RVECnwdm61iqEIcYFvOhO/0mQS7+m98Lv3j//EGMDsn53t19ueyrg3TdyKL
B3hvD2VHLyzUdiKZRUmGoZq6ZDT1raJeweqvkSJpnLt5Bu9Nc3brG4ewHTGU2LZPSPDrWtn/lp8x
uOmQ/XOZ1/vWeRAMYFkDFFcgTD7D+YlwT9ErPQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20784)
`protect data_block
RHfMwwL0uj8vQIsIA30OPG4QcIYTkCF9nPw658oqh2BG23k9WvJ+LP7Y6N47Yf8nohPlpc77AjJI
iPOYzz5jZfcq501no0N+Pm+Vlki53i6SIrHoGRN6OuZMQRsoNq2l/VdbfHCl8IJqsAMFkk/Trfwm
HsMTEOqz+MSjpmfHzpvODz5VJ06LYvDno6ykczA+aIGCru81IjP5r3P9UY3p54UvZh8uHX/5vpbH
gB6P1VpzX6IgW19eLeVLNjVbqf2v85VVyf1tnWF2b1DfEReBp9+isaV8E+5aliN2UzGRVjLcUFo8
ulNW1GOHIu6IKUge4Ddgr99ARtZZN/MXB3J8wbalnz5qlYQbZjzJgMb9yx/v8RMQfLiJz2bOFdm8
P4lGRwAdMMDeZyvwAXdnmklirmZ4RoCJMALWm2gM5g+wa/vlYjIchXCySARa5GO4lG/n3RnfsPtR
XKlpXYWAPeRHWlVp6dUHzjNuH+bE2g7avpeNQAy0YPle4arjG6jv3BDEKfGmWR+fgSkHfPlkXVRw
8lJc1kgZxSyzWtEMonO7l/3/uUSioFEBQhJbaEjcyJ65QKEg2J7dzaycs0vLWSG3No3keOpxg7eo
mHqzWHT4cwQlEDg7cgDBeak4i5j6T8w1I7t7pK0Sg5YV2jNEkRkTjFZyHdSuOVsG6D3LDauiLMmM
IBEztXkJp8Lnkvgyz9963bVhA4Rv3wUR3EKqJZcz8xwPHWXW5WhsW/ir2cRWH2Na5mp0PHWKhqUz
cX2wctyI3UWvrSCm7p5mY2sJOCMwx/qFnDDcGzL2PrpwtlGa6S3cLtW0EtqaXErmeeWYT4rQdMB5
zrzUX33pc6jmpTvQYz1rJsd3PCfXQWOOf8scHmJAj8wtyN9x47UC3Nfhrgq21t1Kap7rX5iW3Qan
83dQwtWtn12kd5LztCbJpNYnMbuqiZnJL2lXeIDoptkpRx7QQvpzceLZJ6Tebo3wCxQyCzQq+HJj
I+9O+jcqwgyAQ52jPrf5SXv6EVvrskvs471YF5tapVXboZ9Kj8IvfqFNRmPbFFud/qLNzGijNnLA
q5XYpdXPEh2QZ9TR9jFej6mZedMiyI977oaT2zkiR99KtTtjMdTPhps3r8p9yi4F+af2r51aCk+i
CyW50It6dERt/OGY4qGudeP65AXhhmmwJrFQhSq4DYtHKFADj2nuV/86f60njTwUrFCrPY3W+H9W
WEpncEizbzm+C/VLGidripAvtfz3jQkEDoVyWY3hjD0mKpR35MzqmMQ2RDuUytiOsJH2Ag9BFQye
Oy44couVjslmwRrsMa1BSEKkuUk2nOMmK5B3PdXaTzcjm26yV6MpXwG9Pqr40reVyQP5NuXUJDwz
ZJsDwZLmEDePjAvPspm3hvx2GXy/8kY7e4UeLS4UxpI+GbWViVm0N68z1r3a++psR9kdNmXhkjwm
jqYqeb0Z+2ywKUi02fOM9+ocIoUTRkqie+hLsN3MrEtLEbPDGx0gkuazuUJeWJjthGt92R+unHHQ
ddOSJV5uaB3Nxdv72wavsCVVG9DHap9qYDzU8Q9YGyVqBMrME5bn0KUPMKpJXEez7QYEH+RORjh1
32wgAOOcIEf5tY1nXlfE4TLboKwWF47B223Uj5D2/9Bb+//NQmYooNTF3oyQ8RvNq+eZsT/yU1Kc
jlkANMinjD6mOr255Gn3/rpmvSUgy4MWtJxS4fHavftExztY8xTXYZgTFVXlZu2q8MNNvwBevEDB
CqfuLQfUYP/SmRXMKv+LyjTJwSBUOj91Lvfv7EtC4mVU/ocCgTg4WOWkv6VG5EF0NGYT7dUc5zNa
tWO4EEZyA6o08HKc0ji+qPJnK/tsx0tfY1HPz2NGZBPf0L6GnEKeLGYwsz7wZFOFcg7QqWh5ix3t
04KazY6JMswQUl6J0c6hlf3qqhNXMCB8bZj0/EMTefYS11GUt6DUQu4xOFjLBDDCwbKozqPoBx9r
IUAs/LInKVqh0zvSeWbNiCLC8CdrTm5IS1HkE9dVFabAby+2nqXacIW2JlWjF3XzipsifEawOBD5
3YZJ7I92Ww/EBKcepTJLVapsGUS/cDvONgEeuWEy5xaGt0oUTPuQaKeMH1CuxcswNZiLfc54TDM3
wE4yamxnpHmwIGVUc2aLOOPLoGQWnGF2N0KpGvAI1l2oLGickHc20T9bm2NAkTtQxHfKLtg+skZL
lbT8vb9fvQQBprqvwuuRrX7Pfu3XxfAdieUgi0s3FZXXdBdEtw4FI+zWg+FWGVWKP3RtcKrYi6Xu
N1ENcsgvGjjs1NIL/qpF3wa5UyMu0z5NpgbvAbE0b0W+Wb0KntdCDYmm4kZV3ZsLWxa5d0m3sYwF
sfChbGYD8IdRX+wOQDEM33DKebU1GSflJqOofDDsb9w0JICjTMeGZB6x+2oOJQTNXW6nzwd/nD/5
gN2QthY8R2Ak2cgKpiYbQa6vevoE2IAWKKGLJQJhdS/47Dl05LDU6OyUyQF/I2vKFAdf0ipDuea9
okGrcVaHtaps9Na6VIxb/EDLppYVmlOUAGu7pQy8UCftOKfwyH/kAm3BEXrZQzX2fyLnWdETFyUJ
4NjTLCqVqBpXk18/edowcEjL087C54/1mdnROasy3vqg2kwuhW1CWc7+36z5M1k/B6HnO89Pttwj
EWA8D2R+VenNW8QQW9FZ4FqcQzEasy4OAZlJ8WEk/hBqoq3gP4etNwDnTxGEQh6K2wnXHdJJcpzY
1EB+NLD9KV4s3+24DUd/6unDdUzSxL7crHnr/+PRfkTlsyRrwsZaNZii91xVeIVyKgJGZXWLpbQj
J7Cqh4N/Tsk0LZ9yTs1CjolmhXX6RliUzGZLvYuNGNQ/AJavZ6DnR6NM36fx/XrUlN9pX2y4rM3f
fTmbjiH8+ATZvaEX/t0DUkumsgVTYF8o5LRRtNJ63tu4l5sQU9euaT7bowFryGEAaKn2+AJGrvXZ
A+ap0KjQtb4TY1qe6etTTdCfSvSjM3MZsJryHkrg/Qv33Yt82lRcHta34brahtry6rKLijmKvAKh
jClrp/ypEYoE4j3kI8w51Oqf5PBqBVF4Q5KiRfANyoz2J5ccy7ikfZZerBkZR5OOfWumx/w6t61R
rWrWiD1MaZY1DNHd7dC6I1WPTHhNTh0A+HCsYaCYQXWWx/WCMoI+QamW7bD5CeY5sCAclLTuJ63o
DPLX4Iz3eM4ZEX1Mf+W02FJ8nT1P2dKg0M2agUVEoDs+vJnIbbXGIjJBjZtzFwVn3v8sfIX8OS7i
t3DggbBaJfb5cogi1KnC6R8QuQAq6uHJquOFaRMfb1Dk7BO5Xm71TfUAwJ9sT5Tm9Oy9f39Sp3Pk
WDOqNd9MVJWOuXdg+C7GEG4+N0ONvWMoF6SDAO7Rc0vbtfr4WEprcd5lT7k5/DvBCMAI0PKp7UpL
Iku1XPWg2/w4jRs3JQ0Yy0+WjWWRzRtD6b4SsOgb5qluSVpXa9z4eRu2e0jaId/3z8JK+y1pIh6R
1jutX+S2n08jumfWqaVZsBLT6eom6FIzzbcZEXnB2bpsJ0iA8RgIr8ax7oQ2MV4lY2726c9uUty6
p5YCgXhaSWrngtVhmAvbQeiIxiReha7liswqsVAXjiX/ySYYH4/ve+3BLjk3RWtt/W7I7QEV4QSm
J8x4ivq9I9rRC4OIGso99kGgD623LgTjyxRGC+ehE/RVI61/aBGdWLDI+2RXabOix5N67/oXkA8z
HGS+5We9kw9AHGYrRNb5e84U4v8gRy1T8iS6VqT2I/uNQKMdsuHehBM+D41+v0YeCuSZ3E0GrUGu
CskwVZ6zaqTnZOINZ1MgqymdGJ5tHEm+/Zw591KO4c4jB5gV6liPrvpQpwfWc9In6nrv3v93vFha
8kyoLSh33J6RAD7dEUHp492RZBBV2ZXr8GC1K5bo+z1oNpEbX5JRq4A8xRVwzN4KDG0vnOQehY+5
XZszWlRIyknvTOLyAmkTjs9CGLhhfBm2dCnYLxewLL9gcrWPbmMo70q0mezaIvvqi7JD8bhpnc5t
T6RgA0rH7aQd1srJTAYJdg/ZnruHkH7mi8pyM7JyoPaBCmaIynEmmlD9OWh5IQiWPLgx5rjbRDR/
mEuPPADk5S3EB/SQ0lQLvRloYgamSyjU6U86yiusymS8molprz/vfYG6Z9qn7AQVMGGCFOzZUlji
8RdUCemkGFakZtaUCNhXWLjinV4VmJrgHDfXBswLKE2QiKfnJ9H10n//WXSSG5em5srneo7/SsRB
v43y/sROxsUh7/MVr84XFTd6oPG1Bi4fNhp/qlrEUww4ZPC7f0DAAcogiK2LFhzDlnKUpFTQJFbh
qEcRMVf+zBLwbBqnLDCY+bD2vew0CYFCr207QuveThJnMCHyCSW4GDgmgGkMi/QAuU/XhOltgeqW
0kY02c+5wNawBDgO6BPmCL/Wqglg2aG+CbpKZI0z3yJMyS5HjFAQLdo/SNi2ZDdfQ9hABwYYIhqp
7EMbf+U4TtLWP9n33sFw/UmAsE6g0nLXKx1ajpc40T3B7dOUA4zVXkEITyl/pIRwFSZlUfwn3YnK
hRHC4yAVqCv3ZwaYdJLQvtKx6pp0AeZ1CJPnhcsXG3kKeD2M2AOn6oyQpo4nvjWU429ejhCy4O3E
LG1XlinT0ivfd7N2V/mO11fqy3Z13+pASau79oU8Y5MAvfZg3cV/K/NO9eUk1k48B2Jo0plbCrkX
IjT57mou2QDNeI8t0qhPHouzcVjbISTnfcgjbNCtzGEeIFKhKigFfqHvI7Jh5qNGrT9iabAFzCYB
DvPkBNfle29IxK1UhkJG/6teGuEghLXfIy/V+SgfwxKJq0Y7H+y9EwQvn0KL0DOgRoXylGyWIWd0
psDzilfsCAcg9H+wjWL5vENIUKOu++f0x0rmA65zAOsYd85MmQmZqBUdfCRhsneiJeF08sGrgObx
LjyUU2Pg6z8W0D6Kez+PWLa9bFtXSJiwX1DAEtSIZZ/aqJQF+zrFWjfA9ZzrJfGRuEUNVlbGKPEt
Ssgkm8OdTtftQVex8tynDEHwWaO2jM291N5zHSzcCNlvYBUJVByBq/wiDYcGNK4JU8/gu2yYMCAK
JLhXxbibzo6KExFPMwo6wUXl3gMWT9l1jQW/eLnvZbLCO8uXwuw3gsxznrJrPxNK3+RCFm4Tk24B
lPqAxmk2Wid00lxeYtqEeBuXuDhrHCUthtBspJqS/P2qJoJRdXXSxQ7sdMS736yHlMvisuhYzNtA
hCywtfdNedFymj9Pz84K1zIg+YqI+hUfG0VXmlG8Voj3wAnEqaNfTW/F0PMLUICek+m2jLYpepVE
yb0SkjfU2FAqw8iNxkfkE5GYsw7LrREF6NYIztoJXzst/5jklETqtlOlVKrpFCzTdpPkQ4FwCQuz
sNi4Ueaic6xF6DuA4+4VrqmvgbKeOnvr71fxEprVTP/HkXzAcAQsUpVQVuxfPrcy4588n+W16nKn
6Htdo2uMWF0s/AiwiGA2e4DTh8hxgfxsGUDz3B5l+irQ6H1uOHbfrCbmmZVoHhV5gxvlCl3sh74b
G7mcg6TFi0+0nRCLyxLQ5dlPCSm+Xc5x3EyNaHyUEAZ1+9gH8jPutXRakjfwvOScS9pB61Q74qCF
D/CV+ObkTm9oIBXrOjQMTSZ3UlB3+Bw3vW0CWJlQlDQ1FcXsN5r5ujWgl1vyaFQSceIg5w5ar5lP
eI58i8Csh9yJuO+UksHoyVCLdmrBetl/C3nGTd0Er23BfUzO0BxkHRTkK4ImJWYc+Nrbq/t1+UXj
q1Cvxx5sY8dAyC/M3AFIIb/A2gmFbImuZYJIqkzCW01jkfuN/g6p9hyB6xnhrNMZ0+CkHoeMV745
f7eutr2pkGlvsnKvX8giooShyPD9mI3NWPAQJVrANe2P7dQrnNFWSXSy0A91Tcsgtj6X5BZHSSEt
MPFVhdEOfCt3sVpKA8vP2IGqIXmSBocGAxwLDJi1zJikObM+MrMDUpC5SVtQ/a0o7/fPyzm9MSYo
9d1gYTCOxSKxV+ajcG1B6D+PXSe5t4MKdbilBvfyd/e8E+cIcujo9wZj6PlI2tU28YjsS/UfoFUK
iraxx8av1HYtsq6RVEpQcg8xGrHGkUKxwG3tWuX6pChsXgCWAIFxNN9ETJLAGA+VkTMkGZ8cCNac
GSMlUsfxtrbkeN2GkmnkMmGmJjbQulMcya3l1WbIlzX1MjGWZLqMNEeGiMSQZT9xplbI4hXsYOc+
syI+V70BcKbdi+u/IDRhqRZ5Xikan3tXHlrZm/k6TjxO03QUVHp7gGDEsZo6O8Vgt3dFr1UJz/n0
R50L0g/aPeo+I67AaSU38JnZnlbDPJ5NeMc9kSQeHNYoKsosXq7+43S0pEOE9mArfgq7bExwcRLg
1/rsTDDU4DaV460Mmo2+S1DuU+uo5EQbAvbAbHrKRZClJeLKRuQicjUlayQlC6LPD7lT3fuE+a6L
ZCJCWoyZ8Zbkgx69H6T21gldQYMvoXjsyxkY/8DF+ljQuUYVH4Y72a1KECJn4oAY1Vn55/M3S+jm
dYG9UHEZgBaIWnMIR3nxTecSJWDS3zk/rSfKmM528W/NsSBRGRO2fmczfr+BwYKLfskE39+rO9Us
hgHKi1y/SKvoQuqd7GT/OiFz1VHipLUVviWn09nQBtg+aJ0y2RRmatWI+yO8zL6WjPzP5wdinbXN
yfzC5oMyw0FqO+K5sFMBPur59gUqi/XrWTq9HU2/xuSXzOhP8UnOkYBBVURWe+pktv9iCkJD0ln2
poo8/xUngBJ4Ciduj4JIR3iCwMWK8ty7s0n6yXL6+a6qBK+EsAZQB7bkzlp2qAtfYg4lnf6/hbVM
m/4q3IlcH3707P4Cw5TayDSWiuad2Xn+mM1XVekgU5QfdxZBPbCLYbW2fd25/EKKNek9F+wZMdLn
Z546Slct44+CjZfssk4KyIeXQG2zuf06SGLxbv2HK8PQSH/4wZxxT25mrfYNRdks+Z0vCQgzqtFN
lqEe0o816gvYGoxB7/0W9QlEv09ZDsCCikVcGcuGCeIqvg+5mUg7IJOfZfPJr+Le1+B0wsvUW64P
b3kW3w0JGXULhLRdPX8A9t/iJ2uUVlKxnDeFdHyFZn1oxZXErQ0EEXMsWWtst1XNb/OkOruA9awr
gM2PuJWDDao07XEZztWk07dSdsGb8BrSwbg5CHsQaLikfWKmmXD2lvWlpXhzxXg0dfU9qi761yEb
VRbQQ1kysRMnsQR4gMSCg3gtJfR73mBByZ3C1URtlKTYlYI/YW8ExsA0qjLismXJMhomP3r9ntEy
GTbci1qL55uTisYoZ9gyrsUGCGorIYZ2vq8sqYQnWLzY4UfAxsxBQHGjqxLt9+eQYIiQkunWIqip
Ov1R9L2ihiq9WSVChfslo0hlxD8m3J2kfMgJroo4FCLNni0ipAkDWOcSpwiV5BLUPuqfqYS3d/wR
DfmikRD/+/IQGYRYa0+AM0zDMEDBqxQMoWYK/KorlIaZ5PsF+XRubEk06nSK/0DfOIq79NfGUaMe
TpEUMo/vLO3OsZfVqYbEmAta8D26zLdX0KlCaVRs6pMM2vqMp50Tv5oRkAQXnbYl6cgULvzVNOd2
qe7tPGKr8imGKkJ7s2uinBPmTHH2kSOz3pIoWxonG4RleTDyA0LlKn5O5UT+d71jGMUcs9neGlvf
55hSo/RMxIIq8doYD4+p8llq87wmXvdtx8cNCgYHFRfSm9ckH83NSDGO3jfTl2B3VhFa00UPQ+Kp
Ik5gskYpwGL3FnNBQqkbe6ReUkH/iSTvR2CMsCOjVOXXwGKAvRCeWHOdwgZ/ASq37vmSAi/z2TXy
QQI6LksbAGbjM7m3fzjgWHJWBZEM1YGCPKkbKaImTo5W14H6gjJN01Brc97b0aIRm4ozwm643L0I
d9EPQSb6+QvJ9S4GAb4PJ2NbUGoSlkeMBeztuNL06AfNvDxOTiDKaRej2Uf5KA4JRqDNOEfk0g8E
wdqzdDdOimKMrMffQAzUw/7/wlGmEQdLa+KlJap1L9QXrP1+vfnA0tZ0CHTakl4P//8d9bclj2hM
/gjnhdJvxwateMpXM+g5PVjzi5jSGzzZNg8zRDmJw2LhvB10pjHvLioFs93WxlxGThEgaRQ98iyT
ulskJ6zS/Ca0xSK++eOj5bVrFPQNQ4othxlfLpDE8R8depBdrV3G4cmTjkY8cvx1/8WEdKM6E/Vk
S5C3Wk00J/60X3NwyFLahOiIStxtmlAzHWNAcES11EzRsbZD17lz/pulAyogd5cKuDoQDpUMWHpL
Qr37wa9o+KAlKbiEDGsBMNWr8WFYy7kYJ9V6Lr+WH49PuPnhS2SuWzQTQxpMuhGuvkSu3pcMTOFz
M4Pc3Q0HPDx6nSOHG9OYFGrkmAjsFDxZjtvQDOlg+Okkz7Gqv+vEaKXsZcrnVZpKY1wWijtAC1J1
qQ4+yeaXCWmOj1Qe2M7DeAz5kv/pswXtMN6ys28kaTCjKvnyJbTFh/fou8WoNW24CXjaYu3luKXX
KJnwB68uYx0ZYOLMW4lZWy5i0IHgIyb+gtR4h5+PXdcS31m1InYzUYy8jYiYBQZB7SnBYpWqHLtq
IsF7M5sliM1BGCbWiGgJX+/NYU5/Te7b55GzxsK0nJKUjCxEUCyewpirglTUkOPsXgSPEWSwWiyi
HJi6ieiEBsJA/Px+AGfnyOmdGwMvSYOLEpYVZ3aNywGYUF9/f9K3fT2OsAp5bMzGtsMkp1TcR0DJ
SHYL1nt6DGEMrvsnDpCdXtmPHWFrbYp86umFlOrt+oePlmYRzvuV00+Jb7/fmBhNyqzVGHbx0p94
F9zL7dJCQ18kCJbkf8ZykxHHQecb/Qt8QZsFfdY7jvPAiMXyKOCBPOSuYRt9AHP1g1UIN8bYFxTZ
wAdC8z5AI/OxVRJOWs6wzuu2y1rwRirt9NKCrwhjLaIWIVHUMFZnOKrTNNnsslr6YpK1vVUza0x7
pSGq3Dm6q9yY+WUMqN2j073Qnd8R3SEIoVH+y5zFQWsrMl+NHu/b1jiIzcUVMOyNBY7Eiev6TpMp
GCLlqlNg+7DdnRB6LrR9HGM1HKC0lONOJbcenmABYiMgSlcilKkYJYABYmYGhIT8hxy3A4Sn+U4S
Ma1k7LkC/qolay1wlGDIcYjZ0FPNNeFedmdDSHtlRMQ0O+HkXvYjayXLrdp6Y6pzloqgaM/RDdbi
XO38oFus75JwMHj86lrQV5RITmfCcsPYYYJQc0bIfFDIuidBry/M7xzGUmoyKFdQuty97F9qiQeP
wTzr3iZBjRCv/dlaBHh9oj6sfTEodEe62MLQH4C4a+QfqcR5vIpz1RIf/aJ7HHPk+qNzZ06tO0uu
R5RdblBYmQ4ro4Sjv4xTM6kzfpK72fUICEtoStz441yilc0jzJmcQEFfB3KYvy8IUINoXe9TjIoa
SsPG8LVODOEtwNnE/gBE85WU4e6ZsDtzUHWsGjQZWmH6Ege/iksGFWrO9avkTPktf0VNFs7va1lj
Ez5kriUtyAIhFCDMq//PqVhL1hKRazQeSSMp/i+sTYNk1n0xr9xuwR7dWzsoCCiJYxGP65505hNY
xSy139k+i5j9eojSevcGGASSBi95qh7FBMvTheGw/KK6AS0xZ16tpOvaFCxKy26QQmVtsOkwYAoG
nxW+wRWymi/OEoaaaw3qM4DxVHGLWpC2QXX/t8tDY88le8bAyrFOXmuR2LzZ1QhjIXc8IxoRoi/q
Qfyz/wzMuIUyqcMthm9g2Co0ZP0YP/6N2mMGj3VfAg9xPI9Hm23pJP1E6ds1dCR17BQNxOef0YsH
GeZodBkf2Y3OXnYy4GnEQa5f+Wiz6LdHt+w27o21eGUvHHFuw9otj2A/yaBEy7xgASMOwzhfLzJN
EqdVN4meCcms77VNC6jqEu+Q2JT7CnM3AztmZBLAUmya5eK0Y52waITskNUgqDdz0h4xeoSBP3ai
DRN2C3mBABde4EWeScHN3K620+EabMFd9FlNhJS4opd2ht3T3MXTeqUlgRrer24lCLGMxdMon2Ka
QI+Dp6NpSEAj/heBFTzLbhcy3yMuzJXw1nxsMbiQ/Bb+YME6Cu/HX4XEMhZuheI3Bif6ZRTaaLcQ
fHhX75qTOyjyHuxvttcNB9Q+zJ5LNsOnqUQNLLDuI5oaAqAqt80Jo5OoP14LqyeaC/PsgFxQXhS0
5geIgOIL1RK0pnIaZyufLIqxSZCSCfPS8JJpVgvn/UzwNeQttuAwyMSadHEwvORikk/LDaEATgOV
7xKAOX1S+LAJmjcckMNKfSgLZhzk37Q39moTWBpHf1ty/b4wXYHDEcltyVwElDhLX0UFf3vEEtb4
Zp+1luEY/v1VUgo3yEkeq9cdMNC0beI4n/MbWBY+ak4uLUTrMQhS8sWYzbaRqpkwxXb4pArTNTQP
eKohIoevrTJve8NIma4xNoBgb27DiWo+ESJmkR24wSbb3xlCsRe+D4FzvXKgigc5ilXbczE939Zs
z0tsvatYZURRyORY4lpjI3YRbMYDSvb0y0RZXJGYVQL5WDnDMH97eOQHyvuL67uEXkCQrhXewS1A
/YOUbly3seRvo6BrGlkUERMDPJvlJu3/IZBKyaTWmzZ4EfFcB8D8jqE5UO2tQCVuqpLHUmhLgLfx
zCB8kpr65YzlejvT14GNFpJ1ezhEUna5pYW07O0Mjb8Y4I9I5vGCsfJTDC69lvuGZX4VKTddTC+k
S7aRcNF8S7wKn+UV3L8U9vZmeJFVQg83JApxqoEfNyzO3aDZCfWT7Qmc2pyLi7zfyijrM0gSey4b
5Tmx4Euz+MyY5ihnh0FvDKoh+wIfr+pFV6PRSNWN/gAY4k7ar/TNVr1RnyjwRcL/awJaskqEZFW2
vKeWIFrOzloADUS1kxV12RtubghqlG+9oW6UnlXC+zEMxNsURLCFipxAgQXabgnvxqyiufMu5ecI
/6OAlcTPnj2Df6kdZPcWE+o/PSJ8++ZEXchPKk8OzMSJlBSCysO9ewj2ic9DC2RFpDnPA96JzIfK
TA0eiholua3K9wggi7bX1FlpvqLGcLA2DY2gybDdgTetyl0SQImpJ3hByAOAfSxQ3qUX1vboyrza
cKtOkRNfbEDXYbz5heziRSfbn3u0pnp0luBcWbsI2kEgGRUJxcV90N/CMRB8jZ2vlG6hgXgOUSEs
wDDLOtv2X9GZk0Pg6FG0dEBwscQ/EYqU+zrBYIs6cQvdX3gzwu8XmLikinzAQunnGRhtN7t/naXq
deWdNzBqOZ+J6rR3tEuos2R6O0WdNCq+m9bpjUZW4zocwtwRh07OUYMoO7PAS+96/G+HUSTI1q+Z
Ka76FWtPF31GNXzjMLIx4LFSngvbEaLkdJK8b8T14fCAtvcaOmi63tzadxlr7lFpePOKjiNnTtjm
mkrRhXrdvmzUFGIcTfQhWguZkjQETjaVgBfY/riqezEwNWS6kCEJB7zaFn37qRJzZOQlUhtYMh5+
0NsstMClqos3p2SKK7nJxLO7jvt4ryxDtpjU+DjuY9yEPbaY4kBsyjLihKU4YI3mfYfBeLJv8SAT
2+6ScdqOykg/JhhSoYxlRRTZkzpg4Br5mxoWKpYqf6yNE0RseXp8HtpyvDCTz10hdKCQgULddUue
lYVHJxxY6oQSXgJN79VgT5wq+Wno7Q/3LR+pfMWy48aurzynsBGV0V9cq4Tul4z0f4B57LmXCWae
Q6H/9uwqy5rb1s3VGgz4D/4JMYoc58N87WILxYoyXJI6RTiHmuuNhUMu/9eP+zhYiGf68KM4rNsp
PU6tNSTDsv835Lb+0oOcj0wXXsaTHlUtIxBpIpZg8NdVoRQMoopg7d5M69Cxw4m+CuEliHst70uo
clbsDn4YZDB0u3+/EjE8DUZyJbe5hr980PE4fbqqIuAbnRKytU4Nf6xebfnahM9m76A1Eb0jzNh/
0drxTsyWu5YUMWtslgRn4TZyIxx8BREkDZMXY9x+SC0urWis7IjicYWoeMN1+kyF2f4WBw+9dq5x
QM8DbIkVQ8vC1wFmaIVUweFZQtj6nxEJTOXw+5x2I0pKmWhZrizsL8cfBkeca7M7r4PBy2b0jg44
OvUyoRW0EChAVigvjGNpBwN0he01ibIMfl8qQPxNmfhj1KFy6EflutJAyV3DJH4V2MdjVeJ0YJcq
4IVTaplCYh3c6QGhq+wLSU5beX5+87Ou/pmtjamPCH94j5QXU1EESTeyOC/Rqn0JPL/YSE74sDPB
+zZwmxRLmEDLtIB409tB3f2UywgR8TgQwgwzK4+PgB1Kv+BSJnqT7iI5UXLj/mPl6F4d/kg4LCdl
FX4VpI1oF7EuqXAvQg9JpFzMsmnr1Ud9eUctO38Wnp8XzxUK4h7pYWaMxoYb4jNrPdrg51LSeBE+
CUlbbAxUzFDPlBA4ZHY265BiXjm/OX9S974lNsmi6jVnfcxSxghykNapBtfpuqdxmqOe5WBexkvX
ty6PKwn7I5eXrkMwZc2tlGrne6+OwQTzjagih6ABbwdGYHRc+ezDM/V7OO6Mpfjil4i2BvZPnMcl
x+6sAFqHZDBmOKagUrLV0Hgt4A1zI6UvJagjd080cQIP45F/IXOJKhnqcxclvmlvxpSerXBjohSS
Qdhj8aBb5VcvWqpxVnEFO0NpJnnNIYNaTd6Z0KFgCtAKkLc+R0SUJG7GqEq0KdhRYW23WcIb6CVR
QYQAgScDQop6mrQ1NEwXCOEswzGDcOGa5VBVq11ggx0IKZqJHu835vt/lxfp/ZWAjM7WEUHLaRUF
nbsGS68SUqbPLcZjx6M66oPsv6xCEKIlS3W0BkJIn7qhXeztE+jHp8EMyA3St5dkyt+I1ZunEZjG
y3eQ0R5w8Msb2fcDwrU5pHhe/tkW0jc9944proeGFA0Fbxr9WTJpRIDuYlzFu/FUXF5T+5g6xq2r
4YfOE5yp4edDu6S1nsaPu7qO3A0UZwzsV6YWrPgIiSW1TffDQJSSXYtlkvuMzhy2OA8MhPbwm33g
eQmjTcs4WLF0RsLjnlrKQP2jDK+iQMJS8wbLCsP7BdM+CKoabMRMOGPPvg6hCD6ZcI23ovUzYfeM
1n5QMLiMlmRAmBTjztmd8rAP2lX646YwUmyjPwGL1yj6fjnUBre6IfnVM0mmgxUXZVwinUoE0UCi
oU9XVl3MqOtUzFcTOSJLfBqwOGQY8qValLkz9Q5/Y403vifrCbdTKXopNCnD8fgywBhSZ6qzsEfJ
zyCKuQUqIS0Uw/b+jwBi0sjvP0xWnnVG4buL12HHsIlavy3Rd4VT09PdUgy+i8cNfTytLoQ3gIL6
+CcRZGWO0LhRV7jJyuvT0d8cQU+nXAfJrozJOBixNAW02jFFpLAFWhkKV0ogIkyVAK4FxhdTj4EO
2BRT7udEz+GEIVz54SEEEfyO0B/319JDAEQvskmiac20xNeu32cvQW/fQ6GHPORUS4fesKkr9bAd
a3lqjII2KoIwtFHzg770V8RgdSmzKH2eruHc8Wi2eI/dKcQHIRLAuSiomIIYFMH50mfM7KVhp8Tm
8VakGXilHOtSlPixPqytdEOX/nr9hi9vo8ghwtz4LOzpODlDUBNu88jDxiRhesI6rvPB71ZlFtCC
/HqdEBkRGwHr507SKnEn63Tk1AEuW7K42wunU3RhEqS+ooqYoGXeZrxVkYFTVapwTxZiBhEUZAr5
iW9UqucFq1zpCMwE3odH0aVA6NNox51w3p1GmMF3JKyTwRkK3QPWMYX93hiwKyKevPZMJQp20P5r
U4xok5y5BxBPreSl2Te4AVtObPtafZi/FtaTowVszjrgpIE3GFSOYgNF3/zrPe/0+A/BSGPu7mU9
1+xoLTE7dB+eNJMX4jF+92O+SWfFuqZuqOx9FjDX9namajlcDeNCFoJQQtBCAi5TA5Gar8xPk37e
ZcEO8XfdBX//zf7Ye+vTMy8OGDW1FhcXqiP5h6LDhH7aUNMSIAmlfxRkFgVms+wJxorGtTJKOH0C
6RjiZwxOOSyF+HwEnbPPEAzTM9gaq6cs10w6EJnojnJIhw84WSk5BcAGhPsJixvQJW1k3Hpbx6IS
91tbBUK/kwXfU0J+2J7hZfRxSR+gXVf+S4qiQ++PuaQ/PeGHHcRiqTOkhsfWTZJR3V0LozyAy4yF
p1v4jZpkKvejvD+ggX0gHq4FMAv5aBXE8yVAcpOdOFUBDdGjKPdcLOzfGZIfTsVi0KEeGzxjxok+
xSN2xzA/2Afyol9Z5G0z/IoJYI6qohADyTpNTku8Ov8Ttvv1sn2NHQEh7uMsHJmAEreS2UA6DsMt
POUF15qCfo7z6bzilhlZhD/E5bbDGE0ETxdX6giUjW4/XGJyaFiI78DDn8GVKEoYw8FaP66Om8le
sLnbDY08TTS/3EDzegwRM5V0RKm4VfJYAVUxU0AmWp53tw4WViur2vkCduaZ75KOO4be9gfDfYTn
3LE3MRxWwqj9pHLVi71ikxNseNMdMUtBD2BooAFKmeqDJqLqWqklWMCgboeTm7T0U4XMhtg9p6qL
TWUATGQBktwozOswSiIAnx/ylcWaVSnX6yY/zYxOEwkaSXMZwqHcMpIzhc8241QgiB7e4enBHyUk
x6S27lwVYHy0iZX8qWzebjcbPFgKejAb0tTKSAq5Oh/jZAjcKK/2mGHgWjFTZb3wUOBcmM515ZiK
YLHn73m6q3eHXCpokbk3M61JjLaLOd0XShwwDlAMI0P7+e+QaLwuWskQx+dzj3oxtE36b43v7wcZ
EP8IEhGEMY291D6XclphSk1Ih87IQSy1rKDfgQXUpzbM8FY2QqXKyIRdLzCBnNV4Z21bxuqfE2aT
+kEXe1gKV37MPmE1gSPh8vazYYKgV8pyy7squloIXwoPKB4Kb3agxJQj69ykqV3WgMfTM9PasFmp
TzDiHG6U4tmErVFO/SyFvKoHacUShxzjAUXHDWOKVWNzxchfuwzhG6ajJl7cRhVI+PdBJF2rQi7x
Dons5PNejx0fmMvhErQKu4Yqe/INXp6ScP+IksFU15ko9wwzMbUSKfxaE9ZNaOYeIh4/c5kPRVqi
d7nUAmoa1PHt949sCsSkUwruGe7yzRq3hEU6tlrFe4S6rmfglKteHd9y6Ft+zCjwRJrHH/uXXG81
YSNnIEkHnOkhq9okMjh6muZTb8TeDVE3p93WnVYPopXWIbiuJM/Ckf6RGx309H4j5t/+JvJ4/jv9
xBlWd+D3cWn2QHzayqgf4ExN0AzClojxFCXA1s33uMUFIkts5cXeF+OObuhAMNJvS/gFvNal52hy
XKS9hI66JuV9BMZUiehUwy+CqeNHW14bokRaODP7wStTFi769uIcrOu4DxfYRTe3yqN/5ZorIqZp
GSMA9KsvGIpIFmPjzUh+0ikyvzJN/VERQp9CmWha630zDSQBmhvLN1TJ/QN6XG4FD+Va+j+YevnL
82oR2hlEi6myX4TbAUNov1y1B5mQR1xuwyWLcn6GkeCmFW0Ei0kieFViOcs3VENOqisvADrSiNHz
0CgLbKDt38U+EHhBvHn4ibc0LE0MZdK/Tl25RZeOG+s7uBcf705Uv8hpkKfrgJtwfugVTgLLJDld
elV6OkU5Y/nKgluCiWWx/oq7X2tI9at2FwaqlXTNB348GnT+c9bHkYWHS18l6YYWd1JLz0SmgsEv
b/vDfAnYvEwhud13ZQItUXIgE7V5kr20/9RdXiqCrNgWVR4Xh6H0NEKvnYM/dQ42AWjkEJMVmmqQ
/Pyxf71WLuSn6l3k8fmszTgatVhJBDB66ynvTH7nW5WdhC5KTOuwNzpOKwR427OldbyfMJE7IY98
NxJwVeaJEoTRRom/qTYua8rLfMaxfyrnAevEpgAO+IHEeRg/N33YvoHWWNF+oN86zscROvx4PHKl
U6SyKWnOnoEUk70scSwSC8pxAMhWbS9p43RUD5pCBTM2O4cP6HF/nxSEHSz3TzPrMGrKr0MAf0Zb
FaDbO+qYNFBB/I/PwhoucR9FSjwH152jh2vvuo+iquk+pvwBTapLlbbHf9QRWe+oIyxCduHv+nrA
qpNUCYAyU9CEK+drqYDDdXy3ecVily5BozRa7pJSIL0DfNnQc7kg7TJSWlstkwbi2Dl99kwByITK
co8KaVKw6krHimGb4F2rCshNiLCPFutAlvAKaZdG61eu79LQ3Qugf6g9n9bqZVdg+O+B4HEceioX
lhotcP0G1Ze+XjEIqwl/qX32YtcuMv/np8uMKTTRbATu+P8OSpnL4m+ipIcybYjufuJCiNyrgNgC
N2bu/PlxUa/oaS7Qj7PjlF3C8XrbtnvR3NQNMenVM0WWRbRuXkRh5XsSwpXMX8ohOsHnVnOqI4db
N8TBee4EC3WqqZ/JmIKg5wCHTaYWMRltVeilzV/X5SjZq6QJ9kSCTYnSnzG9wBBcVF7pE8j65uR/
xShT6ltj34qXqCrNrHyiTVQ8p2lYJddn33x/msgn/JMxcNGJKlFhqWPyj4O3mxkDKY3ZScTW0Jwh
LuZ2F7ROrdmui5od0rpI/MoII3pnCYI+eF2KhBBvBducnmqj5LMIDUDTUeNZ0DGuRLQywdr89r1u
pqcjQsXJbJ45LR+v5CG4lXAtrJlicDW1kvtCVKOSrNh8IHl3xHQ4j7Jij1CGmrZZNL4Bm98blnGR
p5BDaMGQmB6QxhnFYYHMWcE3PWhOj9Yt6NRCkTsKeSvWkN54IKU6WfY0Bw8c1D0ns+BaiMrNcAi8
ZcIMncc1KXQomReFFBid1CXkE0VzBxhI9KtB76EIpxHW9w03Z4xJyJHRv8oVVzEqVg46xf5q/Szt
bk5ROXRdOV84wtFpd+qXfK6WTIHd55ZxCKX8crAWXIfGBvjf77C7SM8pHGeoWSD0r1FzBoQs5uVT
XfwZrMafcqDuziOPOKNnwvT83+AMhEkSXCoeoSwwFX2KJt/4kqqhmZZOQJy/vQGF2bMr8WNT2ctj
pM3teNqnTnl6qUhEMt/GBApr0zAh01AClQ+/sblUUQOt7VNO3yjEAgbFVYuOLEjE0RVBypsYcdtE
BT6AzLDfx08zgHk/paTcWE7MXjr1H1EtdwjY9crT7y9nWEvN9s3Ls59/gtPcJcvtYLvIYzRsFBjO
/q8XmXAz1INqqjN69Clx7yQ4zTBsevPwbjvqu/zl5cSuOsdVyA5oI9auxaVwEZc9OVEV0/TufxNB
Je0u0q3XcDfo3c0YmNxoiWXwG7cigjzc4IXeDoxnaGKCezcrBBKWtsGknPFH+L5BNiNyR8qzGVsi
Jg6zVV81PpYahYvw50R5NFYEtBNG+N8CRMLsmLfX3gAOq+rwxUKQvJ1cEQMYpkZJO0RpIMwa7+rk
/0kRWoFm641c9boKqMCO0nIRI8EHTVT0yNK/NkJRDWVZ/L2wkI8wyo+C+Zdlhgi6RsMDqZ5Bb7hi
iwcyPG2yn6MFabc8FK9xUL+lJHisvnXZAFm4cCJi6kfBfI/MJdVfHwLBiznm7dzKjt7+n5JGzaLi
SWGwgADqWmFWLfrHaeFE871GX9R18xVFGpCCvDtf+IvPyTlDiknuQe2XT+yZow95WoQD3VHU7ox6
Xr3gNKHD9ZkuhDongkM3OWKZtywACHMNWwl8vis9fPBDWyxIdzIsZeUFe/SQCR79dCRNuC61fkVQ
tYBgV6VuD3Bts4qFChqsgL7nnJ6IPHiOWG4ph4KLJU583tCp2m4zCVqLPE5x0FpOXhf1DoIJ+At/
KMEwpZSXIoYivml2CwiYqQKyVKkpw3gsMTvsJPdJfXEr7GybYIpnUSKs02AVAenqV6m4/KWLkzbo
QW7gNFzAfvYH1AAqUmlpxbCW7/rxRoYkIFLnTCkkn6qhpHAjPKw57T1n5TrfROL5TnsWzR9By3wT
Li7odLcRQmJX3CreBSR4XGsz7iBpZStaYX9gctnuE54Dd1GAAu8piwTxq0b2BepdFXRo0fCSrW7L
CsfAd70PUqmFYifZvHuq445qcbOyugZEtg22oyf3dFYZ0CLlbX5PCkDSyuAyZSWG+4pUmvP8j+Cb
OH06ZPex0PD8wiUckesaifWLi0NUaZKSCVVK32dHVkr+74mmmBiJe90J2a0eDSVqSstStl65AElN
vQyxzjnLdNNsqpZuWON0DQ2E69bVBxTbX0eDnKozjk4jpnANNy28U64ILNOYnPuxLO7vK8yjBhIT
0NdHN61mxrpgtAC7nlNRoaLtccCjuBHMbLLezsuRYzTz6XAdQ2m94pY82Evuy4UOMO340lKxbes4
zCWq65cWj76qjHSv4f3BT/gbWRbnmliJGYBI4DI0Q9OZ+wdFXyCTN1sdM6MBbuyD68c8aif0uod1
ANN/ASXQ8/0xKDvKVWFxCZIyV1+6Ny7Ce1Kqve6IQw2h2o7Zxd5QOzPsb97kjI8SJit8LhqqFdAM
fysJ3NgH2drNb0mONSUotgPY7Wbwb30+vszuXQBjUBA8ZMrKz+KXQW+Du2hNShQ0tVMaZjDPcYhK
Y3ZheSQimyxNcauNXFI7elY9+KSK4h9BzXh2ae6xtNPrMgdsHAOlATTWcFLcoLisu55Iiu59xPhe
DKS/6ROrs8doMzJ4OYgh+pKG4ZuvVD1aKJtiNgZaKfkGeqfMyiuXW9d/Q9FMfZyGfXzg4AWLBdiO
ZI1iHWBAJTVqj1mD1TQXVitXT/lf2jXpYZNJUpe4qM1XqdnQwz3EPs8gaBGxsqqLIW2WtuwJBTbF
MyUssw3VONOjq+ojXV/olmnocLOPn8oMO8phVc/2eM4bCs18c9YbRC36G8MVDF08eOlKsafUj4cd
B8FM0EYkAhtpA8gRQTOYt7R2fTSn5MB3hl0NbshiiQOxjGiHmHhBmlr+vX8ykTLuWs4FnaZLuasx
QtE3VHYlbVYep1lICEoJhTTxOXthp+F5FNIbuOxpQPuSfvZah8+ph/D3Y1M1nWdDcJ94TLvArT1q
NDGuBPeVk2Lilrnc8H1KJ/ms7qZQ4bUpMV/Vf+6BbDtt1xP70jVMyGw4Tk78WEk+KqBeZHO8PymE
fbze7D0qHnSBWz1wB25IY6oUu3+0YrcTC593v1AMbJ+znLGekzljYyuBMKxdbImIyKj64sbHeLzg
giK1N621cXWpQ+uckVUXMqFHqC6e84ylgksgk3VbS2luqb8hYFcbUZuuiBfpw6wdLT6Fj5mA7Hbh
Q+fxZ+MOphEKtMp1gCzDEBk6nIta2lhEvxQa230gAYnakCuKdqRfN5kcl1P1ZdebeVwIvHQT3vjB
eAj9mEmaWujyFhNnTYgQtLKv5pzw5qWEszUAzV+UgWXvB8ymj22X3HT7vTHdsUTG8zDd3e5I1wM1
yZnKHYI1RZC6nfyqM+1SRycd3H8NijXP3PaXGhyZdl2snjIODsaLxDhpjoMxuQmQPRtdt6kdKEut
C947bWvwvrjUux9RAZkTS/Ios4NMq6wmMUvuL3n1zTdiNYX2/PVPnmHPwOeXIPD1zxCsXmjyRNnj
Y+htOaKnYl+P1BmVtveMym/Xe3XBkSliOvFXX+4gpmfBmL0lxYCzAWuAfW1W0FgCNtlTZq9dmtUu
CtGE+FqWHr7/GpQQlBNszCYDWo4pnD4bLGQbIbNxgXXOR+Iw/wgalvIg0USpS/L6FC8dyBlEsLyT
kcljL28CRQCkgv9xZ89x3QKzArTg2/PBHT0e3nDsXVMgkASYXHT4ZBS77qF4szrgE+XgMhAkVCQj
HH12lnT7UmSBZN2PSrChUDUcC4ZBlJZY8jwJOi9fvGskREejYcK3U7mLLxbGQkgyD1h+nT1RQKfS
XVHHZTTedAFM1OG14hwFN0Iu/eo4TThciyida12rk2Ffwq96Q3VPaRdbWW8NHc9DXOSwHvEqFU+k
InwUiUOI1NbOtAcJp2gNppXyD4HE8CUx4QCUvKIXf18Zjyovytfd0Lq8N8CPB+LWnqlNYZ68BbrK
89s0mqm3UTWk3sYhLMzNeYfsf+2uetJiYFQ104IE8MVmjLGQM3DQdg+tseYH6MVjm5+vZjkxUSAX
zUh9uPyH/gH82i3T1xJSCn5egOBWVbHdF7VUV1Ijb6YbLvVXDy6cVQORCa5Pe6OwltLyJ4mVa1GJ
JGNCXHMVQMxPNpRKEtiF1a/iFChFFDrf34GgkzpNbsDSG7xjUpGCxa13n5ru7/ZqlJdeCICZJwDM
724O5k0Zx7Vh3zCiMBiRh9E9/WlZTsBxMOJZse3NNrLjpEw4lFfxQeqiSCxlpqCMaCEgBZ303/D1
dT9jrVpYA9aFH+9Lt/ADvC+YXtWXThO3DcdXC91pfxxxr0tcZ3jxxuWOGNuLolDQJK8X4YwF38XJ
xM33P9Yddn5WSZbQPLA3FKMp35IYJvh65AECwBcHG6rfT6hUGP8dyCsvRXxJXsYr2lvoAAVO5TVl
fnPBQZGWVij7fqtTo0cgA9dOuhmDqpW3WvQTdE+XqV5xF8sLOGMY09l2/lij62gmOZVuqOET5mML
Ihttle5EBm6gTd2FU4h5Eg5mKa5+OCt/ye+r1XZ2LY77POdjb97fJnT10K+LW5+etwqmlcSVSOFz
pqEHPCdkfK4ZuXspA3TfWK/3seNbhrnP2RLGJhMBvJqZ+HJM2KrPqZs8IvTFbCUOvn7wWFkZGRVj
IjLdBrptdvyDvcZPczNBQGtZonRjDe8OOv4QocNNRqmeKdxuCrpA2aDS7Gg4XynNtBRbq4BHNk0s
87/qugmplECFm2slNNICDPc9L6owV09Y7mFNoK6z1IB4v0aWUtHSkiHTuoN+iql4WkHjtIpEbgx0
7y30WqS7o465oewl+RoBVHMeyujKZY5Swlwncuq0f7MbTbtk0vnniFMd6Xtp+Blgmwr02ib2TO4X
NymMVZ5oUWbpuLfcPdG8ZLRwo7uzHAkvjO4/xRJlTYsCPqDBfOWsu2J5vNpoHnD/0prSFkXx9hod
Tbr0mo/DdQPHDkS+mvUgHpAZ+kRyaw3aNfrsF6T+YU3INv+D4urPCAtQ+VAM4HDx0urIHEWvEPN0
U6dnHBVdHjQmZzwyfW12mQROc6/53QhZ4OhpkB8jOnzWDEQnHJ89g9BmayKMMIqzlztqyNsCmpc9
vNLMNsQBaOAvhCHQdp3+3KXuwU87HGt507lpnUGHKZeq9+C7GeuNWI7tUTuEbmeFG065USVvqG0M
rwY+Tm6IY12uLXrDXLAi+FxdqSUGIH0/5aj8NghY4eC1xH6iVZLjayGA8TcC6lkvyA6NGqITgnzJ
e1p5dEfOllVJ+s0JEcWiTc9CNlvDkfXGks04ZV8YSpMbpNlZVrGsAwumr42dO1ruVMDN6dXaqf1/
Hk0wlFN1bgs7mXpJCix7/c3VG6xZ6LgqZ6q4irYSm/TZ4TrVrf+kH3XWFlYrGzHfGtJapsJRWg3N
0oal4tsjLweVn8TvaxO05whualy2vZiYVqt65yaNFUIfq57QerI9TKVe5tJSeTILQ5CfiF7JSJrw
PD70xeamztaibV77SYkGzBAwbZrPAMXr38/b2Ozi/KGhA0eW2OTYGdK0LNgOXqO831VSh9PrFhHU
Dd292enJrF/I0wxZN/EMc6PHgI/YXNdpfASElUdlIb6b/bWgUep3W2k+R6aRecq7LjnPaID0bKXa
fOxx5NlekA+RfihN8M+Wnl3er6WxGSkH26sFUhQXntlL/Pm4kBqfWMSS5cEfnKp6G6mo9YUetrnm
up4MsrnGiiuQtW0wNonq5omPMsJykksBw2NqzvcfcPpqLF+Su+bTO13szbXyRHyV3E6Xst02sHHL
joNMhY1m1uS3KSYkPlZLa+jvAaiscMm4kVkcakAyFi1TVcNizyYT6mATKcbV25d3UMzjtfVg5NtC
1c7yLCsfm7MPIVRvLRPUGfk3LSJdc0P+rm3yhD8yUf887vrproou/i3pqzThsfHZ+X++Ur/uekgZ
8gaHC/xNxkG7znJEDtNeuK2ZOFoqT54cKSqgaklbnxRGwFDG9bAmCBUlFxqS5IKZXxGF4MrTjotK
USMBmD86pB8M+x5I+XUoxhIrJdTe/n6SQMWEAXZlQVhEEqMtebKrqQa5uDRNCcyPes3gBKh2vSkE
3a13D/SH1eHDIbLLOJWi0vc6s6fkxaMGjF2G/yfHPVkOs+1/YNIvpmS0E3RN2Uq1WoBNo58QFQll
+NayIiwx/klnFJEceueD7/84l7BjJl3zvwxiYfOe5va8vTgV1N66BaqSRjZ+wuGRINATJwFXAkCW
ltoH1rOiU7Geu8bG8LjufKEcgo4zCTSDILkWGf/pyfh25XBCmI6c98vJRm4uGfDHW5aSlERl9o7S
eHRiFGfsqNVQRo2Ojik1W7Ev+WDt1qPWSyKNY8r1lU13Ia/whOFtVCHfChmRC+JsOk4GGrGDo2Of
QRbwHPB32Ocqf+FhVaY2X9Uvw6MqzCcFNGupkTL4Bu5B2+0GoWhx74Els8ch+vYALtF7n7GgJt5K
szmJENRY1lvCWytd3CzbodZGwUuZh4q7vWh2IsUurNnycphg8CqvOV0NACxRsNRs+JMyKtojBCUN
rfARVb0cbtyEW1mab7J+le17Puc2PxiZYBFCd8IAJ4QvbkbqJ9CvIAfTsgGWLc8/vJbRg4jCQ627
+v9pIDJA2vyJHmiXradDv3yNhO0RkY8Ioy3da/sRHZAyh+Svub9nAmdBbTLG8zxvXz5Shupm2qol
hrbBErWul76hLahkzHV8xHcXEJYC/nVQiPbhTksahudgkDM1z7QaTx1uD3D/By+xaDgyGO78PTpi
crPybBO8zLIlrhTYqG1goflzlJqd5p1SJBYRAECzhM/nClqG+mt3KUq31DRbehZH19hH+wlsdSJs
8mZXWqfqlX5piBnGcp4h1fCgkWT9kDnmJut6k5Cb+RxrLn55QcOcuh4+cFFnkZeIQ2XYWfVwpJrg
pxunTU9+DmN9yBjbZDkPRBzTpoxZ5zjpxlNwSjmgLq9sursavz+PLRMtY3l490bX2U06FO2Db2a2
G8DGwsmDtWDmesO1yVy6H8tQX/g4fhM1idUpwtqC4On5svrscxGQyGS+GuMNmi6RAfRyEznH9w+9
H3CS1iOhE3/ANpvVUhotAnccGCJAOgDaGIGqbQ+ygTT5I4thSPJHfyrL+wly+ESuQKL+VL1UkGHA
OaQGNMONg3Ql37WIUEv4SmejPXtcCxAUant+9fYBcst+GXlvQZ8fdtLVvGFjOaGMZrJmTdz8GT+w
Wa1P3T+v/aI3I1/JkAEl1cqVZSkqlW5JIYuaKWEP8nUwOSyswrJNDjLYWAskn1zBaIFOCBY0Rrli
O2e2zmDmoaaAyU42v1GnMcWDOmM53x796JBw4eW27kdWRgMxXOftLbHFiQBaLt4bgJyakHeXOCPd
O64rHolnc+IKkb28ONOPSE+J+eqTTIdcEoKF4Y/FTsMOka5h5JxzOti2YrTUsZt6gbbt/YZM8+9X
MretMEvPeU/578kRqMAkO6etA7dAoh2sRM020o7GAoRQT1AAIF45oSXW/v9B82OK22FmC1dvzn3b
rFcnAYZCXIbcXW8TpONUKg1kj+szCg7DaYdb677qUq7JsTRbH4pgYz28BljEMnPGrix7NEPELMWb
GHDfJLYIS9pS5VJ64HOP79o12AzFoO0H8vZXewq9aSYssNCmSnSFKB27wv5z4Hmqcb9h93aH/0uG
07fALRpyFcphHm92cyWxl1ayDXOzzDB8k1jz01++/muq3rumWhTvlsvTnqLz8203GNZ7Z/pAI0oV
5847oetPy2ndEkpIWFfHax5WoQWfDBcuIReeqczmEMWEXg8I8Te+L5mv6GuTo2qJgNp6Z7/Tlnq+
+lR9zwfRAGir5DVqC/8LR5bz0q0AREKi3OLE9ruxa/OSAjtVMo2mPqguduwgXlswXq4v+JMZEV7+
bXPGI3/St+jE4t/MyYTouKpVsndmqYRsvgQ31zwNKb/QAhcjIgcUUIrxAab9rdHRAno5kvyfRGRv
16NghIymLhvCJEM/GaYH2ikG7hRyGVZYV699w8dqulRPXvnKsVNWDZye6nujDFHiBl4ByHR+ZcI2
KKB2papvXIkprVWtsXXizyJP7kM9zANuglxSiJdMfpnfmyKPoiL1sssajg6guWcvBMb2z/Vq+S+J
cieEs7v6hhi4yg3pjjo1h3INDXgSKXw3D8m5+xNOGKBqlWtB6F3Ob9f6ukqRGqKdkGZsste06yvg
7tfHSPDpU5gNbCT21n4Cmh1gIpJnX6sBOnWXyPPVtghHnlg7RaImShZ09eGyuUUAWGUUeEUEI/LJ
VDITN0SxsId62RrhiZT11m1LJAAtws5A6c/54qWZp4N/R1fI4Isg+UAcTx43ybqEWsgZ/Vogi/jy
zPvGK4oO9SIc9gtNFl8M3MYdCZr7KHZoZVtM9NOtUo2ytrUt+T1X8G+4RRIy9FpZr0Bz/77o6cjv
K+nJTxiktOrKNe493YDcYicAaju1XFOF0dIDW0J9Z6SB7GIrFZzVfQV1KzmkrHi01Pc/SrrOSrMI
5X9xVzPrbtbRNmsPYgLWZZEgVg/2Gd2KYzVulPdQ2y6wsavCs3f2l1jlbrG6g1Rv0LfG2DX1XtcV
mXGAZDKF+4TwDqbCnfASRuNg5+2eDbCnMGL4q23tZLr+2JHzshJcOS3JhuRV3yfF1yKdx2Bwn0OT
cjfK7eI4LVCJ0exPH7gNW0/4I8nH2YXLO+NAFg83OiRkUOTlVqVofxg2ZfWe2tDzhdfVTY+eKy+C
qMhDVxVWvx+ZzPx4QvESqbEQLlG0iveL9ZECtLEiOfAgj201g2Dfza/mNYmcI1edvntwsb964Gz3
BlwfpBvFYVhGMA0sxgq4F99rVQqRwyHPidk+RtlQklKP3T4SCoSSgX0wy5DhVfsWwDUoeyWc3tvP
6Qho99Xa0cJrLTARDR8focS4WGB/HwWzY2QkaMNKIUHAvP+6Uz/p/6LFaZOkwinkPCFe4L4yDQTm
GQsmtSUjdlwtKE3tZqM7Gb3pbNeDWVOmsdqCqH1oOk/rHf2oi9XQ1VGzfHZe7E32cGAr5Tqua9yw
dldyaT9vTuwcUzUx2hYBQLw8LOQUCApUZj0CrmQ3mBWFSUY3Ko0Tg9ABL0QsjZbuEWCRFLR/POyX
D5nN9tUBgcv76TcJjsiLlF0a6eA8/5NdGnvXt4s9Wy/vu+1ZRkUClNI+URWV+8EN86M3AUjGOmvK
dn3OzUInS1BVrEgK5QUJM9EuBfG0jZGh12JkAI6Mk/sURBqLBZ0zXXsyUR2M8kpaXoqSFPWxTKKt
LoElw5t/LFPT6k5bXewuVsDLtg31qD3hiIbM9Axgqs7g6OAYM6mp3eD1nY8ht5TBbYDbBIvPNlyN
JZUTdJpvmNBafusYb7TSyMVvHNqVkhIAyyTJaar6ZwEtYD+U/C69Vrnvi9qjlZ8voI8x5nUwEA0p
24aWWsrHS9JAIaOCdxXLjgL8KzS6dDw9lDTkUexiwCETVJa9CE5zOLC0kaBm2dEV1kuF0OMrUllx
Pbu3/+K+pcdHyhjTAFlJyP/ZlHaJLvpIFYHc0GRYXI0D8pgyzys29gY3J3IJBhIPJIJEbiFz/ubr
26Q/mopN28FxC513yIfDXsyxtqQ5xnf7/1KvZPRxaVCI+pDV/6msy55vVPlQ7svwCanjN4Gr4mJH
dqfpnMNgG2h4jzQl5NQrELTYvLf5McuMqCr5o8OBr8uDuTpFqVcLUQjvnRCBGlsq3mkkb4B5Sm5K
RpMccvhZFobma5g735FrwvE683Tb+bgRRkC0dksgKsp8ZLPVzV2opgRGiiEcBZLBRTN4EZ7Y0XDq
c4zsFcoC3ImUEhMN4ezBgNt8RbV9LKKOx5fn+qiK8nytYWA+9iMKhuml09qqFp2Pvp34X0kxBEbk
t3SYYtLm8MPIBbiCh0+HDxU5WlV3+e0Git+LkqqiAUmo9w/4YHr0ws48qvOZk0MsBf6R8Y/P7vb8
qRtjk82mcj4D4JX07Jth/Zu73mNIErF1xYttgSydBR8zY8ACYFkKAYV7sUCqFGxG/gKLFwo/lihP
GsZFMl3XTgLgUfKS/BC1VcY1bBziSJl4DlxXP4B9c/q3oM5r5h1vlCm0bFZbyiQA/qcDSOD0grKd
1UN1phyLYaaf6aegOI9A7M6LbYpMwC5uzKl0XaXlOuUCdVx1mWx/d6VZ65XgacvV0kTcyk3P1aZg
D9bpp2iteGWsPxiafaeVoLW/rTQOOwDjRYSnxaHI5yz3gQM5qOVI6ArZNMrMPBEE1WdCTWUvilEH
MfNyYqCLebSdcrpG8AgxRhP1jPfK6pAx/JeCY+4gb93Xw5KOxcLp2epuFdVuR+CxRlIWhtdJuqpv
i0nHq3geBPcaODsNd4wUMNAmZeFNAT0elf8iYZ1TILjK4t06F90Yqv63fF71i1moi+Fm0P0btw3j
sHdtOJzP/q55aKj7Hcso9l8lZhO/SJd2UC/04OMH/mBpuYmeijDCvjVebrPoUZh8rQibyc+fiSu4
h/ArYXgCxhSYbhLRW5Pkp3ye2EIKl0DqmPAOAEnyW2hzmvVrqEmKWY8QaBJL1YwREZ/b0LP4iUNT
/BlvyubPN+XnF6BnrphmotWC5mmEYk0AcWHRtNlbJboOqAkpanlz1DZynET/mj7sUD6tpmV3vHJ4
1A3Xy910N8oJ/lL1KFzBw01EpwxfTKCFAvpBl2UV4huEE8g29licXOzm9LqPabfm/UqfbpBWcZw0
hRJgcsEfl6su3sWm0xvXG6ItctQWGlgKEUgKzmn3E52ES1GsT/2Vdj24ykXQ6/uaJcw5O48vxpnb
k2+XQfgljq1X3Trb8uo42+QkMZ0f4Dzij5OA2MA5jI9RHxDjnb+t5ye+NOrmjv25jBS0Qws9ki2Y
suXmfKdicpjwdpGJ/zY5mZmSgCbroedWLpbL5/5EHlb7ALCIRL/Q2Y75bqP0sabLbzXZm1HC/Z9u
W2ueLQ6qlu6JhK01x38d7LGTlFKxqTa+pqs6czxOuWmL6r4iwVAaKiPRYT549kn1YP9078sWbHA/
Qy8SHvlBoqt6Tjxqq93Bq/vAwe8F65WqrPU+r7wKYZImbElhs3XUQThTYklClAZvRbLVY13bQjfU
w8Zvg8uuqZBd8P7PHeFPBgTxRDNALim2cVry7W3WpyxHkLA3pOe+F0YU31hkkljvQi5NMZPE8jZf
xMuv7yYouwQiAYs3VQxxu2AnsSaJvKYbn4LQUHAKW9S1Teieoeam4Lxwg/FqzR4ktZx1XoM7mf14
9DhDZKJPsSLHBGKhWcWnWQ82e6MkQzoHMnPY2OQnWq1tcc72MjAU0tYs2zKSkOoVsiYnih5pi3RS
POp/Y757pwFr5T9ismZY45edGzw8aoFXRG4zN5jFJMX9URrdVeqQUG6Q8+GwCvYlW5V2Ac5C1gAY
+FWD/L3EYWZ5mixYkaj2vzAUeV7mEQBzLKwbUJdc7l3qtfQ4IZOZEepT+qmfNVtwdn3osFFbNhk0
ZdGgt0DrCe/aVmIaVz6X+M73OziZvWgAW+BBIYbi3/YQz7tr5olMlUpQcAFTfFS6aokywvkhfoxk
x2g9hZhPEx/plB6tluJV/dHIoOxO0x4ZjqXmxaYxyJzM7NDRKEq1HvgAn4fwynVlCPJBQLCp09JK
8WVF8KcdE0vFBK8OFqC8q93PIni136wHmjRFN1Akc4vMIXOirPj8qi2f2I4xw5kRfrbXpRVm118U
QVwYmfmOq6q/lueSZS/JgyLIDMGRXrEBtKktZh3q8DNblaRj
`protect end_protected
