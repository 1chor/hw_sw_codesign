-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OGvF29BN0XjKt3FBotajsCKIVDdKnmcfAgK3NZ7H2zGehuWHVPUrzux0Rn/mlREjAzs2Xniy9AUR
5fUd9VBPyR1Z4IDVAow+RR6uL73ix7GRJfIB21tjeMIAArV/0Awaza0xYSFzZxhTDWE24rXkG0Xk
L7i+IRdt0s3GojrjKwub1wfuZbNlGS7zaPICK3tbcEuZ6b98iDa84ZKF+59leej7ecLauNuLkePA
shLZIcpYeYTBT+kH7lyarHURNB2eloJkd3nOmesa5Kj+XoXZ2OBsPAROnb7I0I+Bxq3ypcFFKupN
tNmwwflvAWXPbaTzX/m5BV2NOTAra+UlhO57CQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 29760)
`protect data_block
ZZr7855QtVoldId9WXsFk7riLmPrk4gJ3E+YcRHWAm/gT+3Ycw1kEL5VLST9MakTjcODPaWvCgzE
dzNJVnKkcNXySojulEvM57CyGE6uFoiqThQCB3xRa1vcyULeBuiz7w4yCbFDF8v2ly028Bn1838t
sNINng377IwCocrB41/hiOAbMLtHYKo9FQNn9NQmUerUUpG3DmD5agML9XRmJUALY1XqyENdeehX
ov0N07w8flcQWHqtbGn5vnlRegFpp67qx/XwnP4rdd7QGIMOceTpHmWZoMPvNeUIXLBBGBVqrJBe
gJERIwfcgfKJsTTEKscViVqMIh+xaHBFtxL95ef3Y8n5c6eAr38EBWUFdAif9pbS18gx9A2z3Ubl
m60+pKL7WW9tWV8HYLHYcrN8B0y8XbQvTQ8G/HE1hdHhPnArEyzbhcYjE8w19oCWS37akUnmBy0Q
2e74EhNlIJZjEdybsppqUcIFfEfH59JEkzHSEyLpKR0kDSqrrHtq66O0cYPUmy8T+iDsIvg+O04i
CEgAlI6YJX64f9ZVVNbLD4htm9miYF9LdI9+dHxh+JgnyuFvJPIezJuwEhttwD1lvI6QFZ+P2EMU
46/IwmPWFA5oubcY0vRbLnrbhQmDQpbaPergfZ1FYMnPjAbIOjpNCZdUh0iHjVZfubmj+z3XOlGT
0lnfn2N8E0Xvly7B2poVhM0vWQoBLhF+7wjlYKjXWfy2ezxUgp2Dlv6u3t9mS/mx5hxkg98cv1+Y
w8bGHJrjPzAl7Uvrdcuc8bNS/ycKKhB5DLs/zCqd080Z71lTzU1bCNjVoWE1A+BArIx44H/WcaBn
YyrE/UmMIjAWZHn1IHthQfEZyKlNED+uqmoRlTElEVVT4Mkj1yjJ6Wlec3jt4Y8Iyr+dILXHOEc0
4mk/nqKyor62zGvCOJwG72a3Tv2BtKuCjjcusgNvSi5oEMrbYCOSTt4I16mPU1jvxuEP0E3HYPw4
vep/TVhUkPK5QlOiLtUVwrGxL9S4eDJ4pBqVBoNb+R3HGYeyZRu9N09N/2Fgm10aHMOiWdOPSTeD
+3PGjZFG/ddZ0Ih+FGr7TmBvM82NAItXcXjTvjPMt1a5vNx9mll52lr6rdrcaTxvk8mHsjMBQV98
Zc5KfYl/RGbBwsvk30VL81dsyB8FSo+5UNi/mYF1BDiRqIjBTbyMI8rFhO91Ln4hgJkMIe/HDDEH
h4qU/ZOzK+I4HIxHO8ZDPb+oPcym4TYSsCXeadmsrobNCLLVWK5gsZaCdOOrTG+HqU6AHPaQV/cr
70KDJzJE4qDPxoln4LgPwW5U7kD1koQXoRmD/+xWEyeB/dNFqgBXvl5ZYlx6FiDzvbxKWuGHMZdZ
O6DmYB/PQexJO+V1Q5LcJBQmhctQcU84m96dXr6aVN9IsQ5C6F5kCeSpqvzAQfXZE6xOUfs77+Gk
Zzh6ZiXlvnUmqHxGxfXSktOw6CB14+28LeIeRMecoMpaIOy03Qt+HEq5ENCpLjtP7hH9Cj1Ethg6
NogxXw3uYUgSmOTG3T9RdrCENYtRADZosgxKSs9FpVsO4AyvSOHsQh/8GemI4HSU92QqA8utJ34b
WO59ECQqSJjlLhzoGncKE80OhYF+LPW0FVN1gUCNHzpmwyqxf4UbzVbRk5yyIY9kMTrmNwSZ3X0C
EYHMOJQlUEfGolR05cylRdUVxu8wrfgTgAiii7GZYUBUNS2O2G27LrWq26QgwUnofVyscizudryF
QCPvBXOLZLuukhUfMTDGgfsuXI2KKWoxKioED+6gNr24lOgttFs47MLlviljvgT7/OI7iqmlJPYt
QthVNM3696SJ45rMK+eWEgskM1BskQjlkkSRwQd7z8NKMbLYoZv3p9b4bNGwvVUUg7EkPOWNenMc
84Qtx+Axl3kgs5SwI0AIkJ0dPwjZSsVFTneXfzs0AxiysJ5IcXKs5qnNjL3JJULEYsHZtBquejL7
uE0dJFQzrz+quqHwVQyYPKQeBqRdH3x2mglTaglb3IhZTG62ZFTTdZ6L9kW1lgVwFK31lD+9oCJB
E4zH7fD54lKnOMTWf+T2cZqlvXoUXKNzBlKw9M+1YU7oaf6KQDh4B84BlJssef/P8OZvOrtoVzw1
eTtvMIKGTImQyu6vcXUVOuJcgptmoBzwS5n74sVXS9wZ2R/iHD4xJKwZqX6foFecL17gDOPCYIZB
tFpOHe+Mu3M/Sj9HiL+/f2t5GhzQzYKu7P4ktftQneNoDO3vmgrXTU+jkBDxzk25sGsqN7kHCOPN
H4rVAjdHIRJ8o16fKw3FSaTwRMBGpz0DoRWN6EMPMJPa05wvbvK1aYDHixy/eGDeRJ4SuBBBudLU
PrWeUpuakJJ/s2F2Y/J9O2Js7NKOMSbzJS2W5EYB7GXWgPbh7gK7VZCGIU5iOnsUU4vzK+D3WOQX
9RndO5hc0P8LAzB11sjHuuTh/kQbKV637DzBBU7xVXoyLb12y5t2yCKER74IxbygQ+6YGnwQGkbX
7lI1OqaUYbICt7TVpU1X+dDqzqmckpoeWQ2DPfp29Zwl6w6vml1iiYvCu1Gm/q/SgD8dLeA/Vb6Y
jJXQlw3SBngXxWh3Ksu0mNlt0AjSO8N4V4eSnKmlpYFDdccUACN3R5PkK+7Tht+5A1BC5Zdd3Xx+
/s/S8K9xj0cTuviLIBdigCPR+c5eOKM/1xYykaS5yqDFH0UFrs0ezOkrGgHO95VfO2ipo7KD1jFc
r+q2ygn4eicduOkDN5hp5SNMBN344qAG+p9qjmXb8GjXN5jG3LOQ1xZoHf/URfc2UeN0wPZ2lfTw
0n8j7tt1QJg2oUq2bm1O3maSdiFqX8sg8sFAhHNZ/GqwylnhJIlmMdxZB8bRpZ2YYwGebmcnUSOZ
RV9RLTyYVq0oeiEZG7SJIOiYqGahI5Ogz+d3Uckl8RyhUKlsjuJT1CdLjAXgr0A3HJZ5FZw5HBjZ
P9sTuBKsddNPiHbrQfhSlB09L9pdb6Dvg/w22+K2MXO1eXl6Bz4mAwEDXN7wMzR86Un9d8wnknud
fm3GVsLWnblRW41nxg7qkuY/p50jN1Z9XYWnSjo0UU8I5v+9C3idelca6qPk2Oz0elTr5payX5yR
Cs7q+sxIRNr6aUOH9oIxD7jgLL/0Nsqgqof48Qk/wi/kopz6A9IJWIC+g6h9N6AyjOip0PcNFqwv
n12DthtHicgq/FDz7Na0JKsjIDI335iXNig8++yN3uCb+KP62V2/I1moQ+v59xOhXGNPlpCFX31p
vP8kGR/bmyosXAZq8eh9HFE2QDMdpKi0HGO0fpeewUIhy/FCcKlNLqe08MvDmhiEN9DRZF/DfTBW
UlcmVd/joB2O+xb/Djv/iBaHQeJAN5Dp7k5XppG0BW5aq4jEfPaHKGV4RpkFiprNVsVsE5zOvvZ0
4mYheh/bwKbzGfpCIr0pWHqiKh7ukQvPebznBQGHVncJUR54X0egGf4sLKFO13v/BWmJV8W8sA90
uQSf84AxBB/4/1y4LK9pyImGjoc7/3HewbP+Qcj/K9pu04gi+4nZfnx8shkp/Ky7gwg14i+0JDee
gKRqw/sBucR0ASI7fEZN9HHsTbMUM95udSVkTvDdawC+P+BWZkAR6a9U6+HGtAfKP9uhgwH/trpJ
DczXqEtpGDZdUSrbM1lfALNX8CXjBom+0nXJnn/LMi3P4UBsiL3CXiIlGGzD9Gzivxty6AJe63Fd
lejIrk0pkb//SAj3xzx9Dy2XJSVvo72JDkTh2wFqhwtz05yKIR7mSVBG+TaKV+lpZ1B+w+//0gyx
tIDd1Ul7hTW04Q2Xo3jLggkY89GP74kEogfUTI+8Y/kdkbUVRjxO2VedPD27O4kZaVXtL7lci9aJ
q7n8JX+sz3YPhJRq6B3tVkpvCFtpGHzdsgMNfnXJlAJjWUgMgAHcviWBnxG5FBV+BGdKYiS1bLvb
26g5Gu765PxKHIze1C3HOgRQft1EmHCa37ZUMXLDVxfyuOSjwB8lcpaW688gtGJb4QhOTMJsZSN9
80mTGrni4WUyUYsbYcm+WXLUimhyzaG4VYzP0fEUawbpxBfTHgtvfdlt0Q5IRZOwRtnO1SGgzkXH
WR0xw+GYSaznEq+EwYQZWvdIJ54YUc3xQlhmEFrAgpl0xFlFnIlpBXdJNnFMKPnLDp1yBXoxC+JC
ck6aXvsBzgsw6VPsP2qZEoCGLy+XSBoriCONkYTkcoN7gy42GBtiPdtqGa5k+M5rPaKcPD2xnhwH
t0EyejJViamNacgewhDV2NlbwJrIsexHhxGtK5nArY7Xvd46yzq1aw+eZKV7NDImh7MIoT6MMe2+
CcA4qQHDK0SRGbrk4asOKFsjWp8b7WdWOYr8UlGvslLAFVJDhz9R/2nNfMzj4ppV3Ao3fqltvNPT
Dhcq0DA+bOw5L9SVXS/4OA8OqZ38NYtfkqtxX1CPoODK976Tk9AGPe8L2OkTZjZn4h/72OEz7zNq
4ite+xj//NLvSUJYVsPhYugyEN0NP0+cF6qfxi/b14MXrlJrRi72VSk2uNbX0I/fNd45m46xB8VX
EtOm9+rU4PzVQoiaHXeOXsdBZ7ph28uFA/tC+U80b8GC0NxTCmrZpMYQB7660GrYlTmD0AYZTEUN
GjwemB64PEFZAl71l+y59OAO1IlBhb2Zf5OVfNpDZlMup/H9GtQX73v7SUSk6uCWvMy5lQFvH2dO
G7zVkIdMU9yAGWqmI65wRTITgvgOfnGuIRebCh0k+ueELMPi1BMih3HSN1zA+8ulZixkuUDkw0Nf
oTHE2OEzE5N6+kAE6/uzrXiiNSdNzwhXq+RS4EOshwx1JfrT1kDl84NxWmvpDSaCO05ZLiBbXffr
sFmU9HZx4estjKg7PXyijHn743thYQa/EaoGbpjj81n+VLIaaYETvFToq00OQif2V1C5jv1lsBq4
LlgOcmYkgEfleNWWCb9psxMvAx5QzCrIuazpKvUSrPch1Qzz4MBoDSFH5t1lY2tIJcpZo4tpG5FB
blGqBZN/GOhDHsPhdwbGRrcpIDsswuUYeVhrCYqQHiXPDWkNvYFg0lbXSTW8SoPgLXF6GL340Wly
sCzg7SQ8TOUd+0pAhKUssZRRk3IkN1YmRVhHnH17qg1rtH6kaPXMp6GLZzOfYwqngi67pHPLNLXy
2e3jk4hBuEp7xd1hp9UdGWcj3MvxbrvxaXYIulv6lpGTURrxmeFzsa4zUU548pGXjule+7X5S8O1
GXnP5hRX/I3+09PzlFRgxsJPJjltuQ2Zgo346BccD+0mzAE872/KKyTck4eIKDekq7WTVotemSRg
V4c98DROWolyEodn0W1/O9CmUepPAOGp4gjOMtQPtQbaYaF9oDVqKdkRuKF3StaT46wRIX7ZeM7z
SekdId8LkDbrEBS0CbduVcsLW/RXujyCnoKgGiwkI5X7e1TSVbp2pxbiXXJeAFoprEQoJIOVWlB2
OUnNccgatHxOIoPRCcIdFoHMH/NIYamafAJsPkBhZat5E7Qh+07VzCjtl0tKL+YTU2iXVeeocFpr
byE5nzmnQSvb2F/oIifkixBUbC3QyxaI/zna6eJmPwKMjKccjCSnavgHH7EdwzhDISJp3ROhtxnq
hP8V3a86feuRKjz2AHHDYNzUgk56RktULG27xQAeR46cd+8uUaEcHtKeYFHcF5WhdmxNFDsKR37t
dLM9r/VEjAjHdmOpqugxMm447G7auAh5UPdxWZUQFnknloUzE2Ij7Qzl8aD4mUiIiKu6VDsEtTGT
wJAJ05O7RTg1o0tnMapNKOnriyNVGqjnIEeTxAKY6OYnT5mHLSMFYP92QiXNzDaStsUuPo42Ms6B
qXXkRkw5O/+f+ZBYvz4bCHLRyOmjE9ZgWh3myHwPk1T2BIxtPEGqn2RaH3wRD04OmISZ2PzfrcGu
LcaWK8AoNDqY6bxMUg+iOaYksEwWz2e4cnCKGrZg7Y9KtdMgHh6V4t74TjXweMnPqAHJ23mBNoJo
rkPSw8NcdlPYGf7YZ0TlqHZYDu2M8lWNVDJTiYIRNJyzcJLLXIyERhfnhzMNTE3I7iFTlRb49LDa
q2gZYlM1k35tmD7p/BMoB1g/JXuJSAoYlCzG6XaSqujNtIF+3U7NHo6gsWmQGvdDxjTAX/HXc+Vy
0DGoPrR+0Zl8oPT+u3nPnW6iZjzq76Cuu4pepY/cmF60oQW7nzddJM/H3nd0wzpYWyOhfUDe3vDP
0JQI1VJq8rctA7BU/Tc3E2s/tS7pOuXd7YpOt8JX+TgtxT/62J+vc41r2rfwXFpWoRpQFDgPi13w
tiHFqrdy8VTvVYZp9wzm4XxBg2I1iPp7rYkHeirfQqMFFajqWTFM8vY1AyC52tD8JzkUCi4NbmZg
ZHnl8mxcU/c3INum535d9t2NywMUxVv/WlcpE6dAi+kFcinoE43loA3JdfpbFLylkM0fi4lnVCCG
nAPiC3jfdVJJX/iEz3WXbO/4JoeB9/KSJJN151uq6RBVvnyCfXSLzDhwuTDPLJElWEde4AHz75HK
n9FHBz1FcL9oOGTBGoAEQvUtxqo0XE18Mkmpqm4BG+iJm7eVNGLIaLyhnBm/jnMAy6yJ/G4yew2F
76XNuMpluLc40hVXxwhm0XGOQ5cJQ+T3KRcweDKKb+4cEML/FdqGoWVprnATxNOaiOm7uMe/vhSJ
xH6RKpop+L93Ng9P9ER5QMSt64q3r8ZkwbBblGO03erE3vuY+nJa7ZXtQ71C7S5OSqV/nd1EKdIq
Lh3eFSAaVBHYkTR5KFzrAQHGPlag6miYmQFrV6N4bXZkvwJ1BmFMfqOSTD++L2qB6vBsURSVs28R
icekjYiuJGz9huTgFjsdAeKCBxpQ/QsjsEgWX6NzvrccN/SM2vOo2no9FzaiSNZOFNCqknsiGsGS
tT9fkdnOwxVt/CTPH6wrqYbID+nOMVhVFGsGxjzpAPZaUTHaNB/XHmFNnK9BP2MlK+z6MFYEVCSW
9BZhdk7uoaSe2soa51h6SdMbvdW+UiiP8kZmJcZR9IXpS21DA/8SZJfXXFAgWf3a/OP/uzpou/9r
+X5BZCHOgtyQAeN+GC5pu8qYbeb1rMMaZX2iJp+3Wcm/SOge80UxH4BJx1hj9EN8EBBOcnVTkgzJ
qTV+KHd0EVl/EKkEPMPICSuSO0kSBS/LY8hP99QcFrLDBQpiF1rb4+BLDchMOHL7jWe9hEDuuh7m
oclTfJaXiJpdqnluUFwDu8hyxlrsotDnKzsH7xAgWLUCRZTM32VByFGlLA+Ju3tIGydBcF2DhL0J
DA1EKDK76dHAmf4T80n5caLkSPxYPyGh3rDEIfZc7zcFeQvp3saeelW/oXHm+LZzHi6ACFkZ1dQ/
vyJzMd/AZ6gaaRIK8kwYU1ikc5brYgp5etRxWLDmsOBVTmS85oL1qEcpxhrYjRY44+LLhYzGdFWU
+D+XiGXuqyOniyHtqhBj3hyrxcPVJHCNbInCz29XjnGaNZbJtlmdvs3H8hysGTnlKkda4RKn1g/2
Ad9rk+Cf8s3ouaD89pbs6iNEhMCPU55XraMtRvyApfoX7ZR+UiMCmr5TRfDdvF23iLdM9avMUNPi
/8cAKmEaYPb/Dg0ZvmfHYJ1XbSk9/1mcJCCI+8Y4eD55X8CAL0VMGTk6cJjPHe7nNxm+1cGXw2To
l9J+0q+5Eg9n2GU6Xl0aeqNZMu2hEv5ZuhMpGKfd8qhLLbKzyezGHN+O7rrIdRywW7vOgXTgCL6F
kqp7Po9OepZseSXz9c7wui6HFS+NrY9LMcO8iLdF+LQz81QmFA7T5PnQTfQxzpbtdeMpLPllxSi/
vCMpADx4zq7v05vGLUumJnmz1GwT/ujEqBLmSWJqvtUGAJvtiTvj7Sy52meat39PKXlJLXTVsNn3
HXfF/cw3wWZfe8zQe/Oasi4JxMPXLLx6Z8mi22NlGGZTtW/MJ6j0HYQgp/HHugb3Y9uES+MAnMD4
Vpxy1CC6TErh+e3esEWpqN5GKlJwIiWqxgshlZrZOCNPww/0nUaLSufLOWdaVgZn4W2p8Mup+49U
Fb2G1B5RJ1H9omU51NDCRUBPsfArQapyBihFlo45D34/R0+XiWmJnY9hu4y6mTz91seZ3Gr1mxRl
zgJT5Vjc9k9VpXP7ngROr+F2xM7BrBhthrse26IUdLPQCkKp+NzHcbHxJUbQEJBgYs8g6/QE8gvf
nM/vn2cCte7L9KUdDXenKWS5ESINA+5xnkfQrBT79MK24+Kaj/KkiXSJdS7rfr3bWJXcX9l/XxwC
HoBJDtznVp6virKqjkFJN7vFX+P/C4rJe089YtG1gNP+ZhnZ/HAmURtLGRUryOPprfBp0nfEM95w
G4K3TFl1aamGkTb5bCb27lC6jwh+ciXylIR7giC/OfVSzU5DSt5djE/hW1xEI9nKozr4vrGRyny+
VmSFFlxTCs/Jq6tzDuXa2ST8wfYQGmDLIMx7Eupv3Mn0gPUdgK9ZlgzOTEUcQf8GmKcMchPBo9Rg
+plaFYR7ag2bPGc2B3k6z2ywYKsTzDotibK73SArALRhi32CLxEhsExfUvGWVMbchvU3Q2xOGZrj
0rmAd0ID2BavHwgtA7rrvjnkImk4Z2giF6tAZXmG2pfzx+Iow7h6ZinQJv0mbX8HoEjyGn3vjqIU
hl9TfLks4x8fK33Zdny34qcb2WoAq0UCc6vlzSA8q767H5rQ5dR5uKFuRi0WNTD+dweh80LjRJZh
8sfCFnGKi72XcOrM+w3uI4N1qrQGdqO/rziT/z+LZbg7Kjt+gqE+6x3UNAP6ic2FeTN3jPTO8Pkp
Qiw+Of0ma8ojQrGSA/PZ9dRnvIOK4oSRfllb/qTRaxtYWFm5F5v2dzIZcjbosbV6dG0PaiNZ66oi
RAQ87gEm8TnpSgHuC64R2W4QeZNg6RgS8B1fPodw9TIKQj0Hy2L6IFaVVN5ZvEuY4pzm/ChTrQLh
tsnC5sUUv7OO2QgA1vOjP8PR05FSVIk/O0HvlMz7RQjtUeB6NtMD7VNMYDDwnDKhXhWraWNm2CET
nuTmQvGtdOsCkJSHHRAth80H/UZYRGEmUNtlTbEtxM32MY0qOGwrmsOlaUN5Aw4gE3HgryijXzT1
HfGFoxWOsT5NqYWcW2DGqNjZnNPuhjhDYk/4EmXL/6SXUGn49k3mSNXoTVJq97MW+5o+B2x5u6kI
gyDvonZn+5gi2DV/9gYH+dkn4tleJIw16qW2nh7zlgb0zlCrEbaqUQR6Xn9D9DQs+/x93/9ei9fs
U0IHr2HNp1orp5ZoUYQaeXTid0XzXErq/6e7xE30PSb4i5e9dbmteUljPiK1Eg2uzJe892xDkqCm
Cwko/ScU1+169JYMkjG+voJAkRE/S7Huz3Ymji7kcZrLT5WoHRcDsf8mzusmpjInFNMy51bkAVtm
2DSji7kAONQYe+5/J02uPRPpWO1sktPzT/sTUAnhxCwmdpOv2JEIATwCrvucEWTmkln9pDGMt7bO
TFVdwZw4+aYemxXDl3gPMBS5+f4c3i4FGFP+GLJeRTmbaL0wfvtJVWGFggsNUUWAt9Igh4aXQ2sN
3I3lLyb9FXMsqda+5VS8vK5fgaNWX63DBGWPulraA0YzENkWztPNpT9BmaVOopPwYqUJUqBb9p3y
Qw+CsV6tBLDIBZ0UIub16GyI0zHBRCXVCCHEzIgDxLejIf5Xt6r1dEELllp3FbiVQd266uflruCD
N5XtMH3gvC4nCUpkDjBbh8JP90KvNNAlpdCsaB9KEfrU2eWRbh8pQUgivQQafYAyQ2pQeXmToMMs
2op3x5ZGxWy9kJT7Q4B/M3mo2mI3UF1ItgVxMc6KS++EYMn4lXOLa6wNTcYGtHhteKyo4W/5eSea
4Ys8G05Ts4eQh3jHXmvw728+QzzfiFjJriZUm8zKQxB3cFsD5F39nSId7FHiHjRCJwH/eLsqz2WC
/fF51LgfLXdeLBcSvX6ShIgM3qG8rWBpKT/mJPBdkGbfej4jR90nYz4dbcVurlcFwF2/i8ieOhfD
Jr0icLrlrp4p01H7sZ6Ex5FKWIqfAtKlkntpjjJH9GgmyvsRhryWJ8LbDeYUWR/dGUSqD80Ck58d
Z4IZkPMkxcKvDSCdi+sHtijrBFRW/ecy4RWoWHWo1TeJ6rf60DYyknf7BdjSwl3bN9z/HGMHc3LX
HmLMifdv8uGf+dBl3csr11j4fcqzmmkSjq++L2TKQoEJCUShJiV3oryic3wXvJJ9kJtYMsxSTfgM
B1FB8GtzAE2itt3gqVmjHsBiWOIKP6ZO/LffCXxc0Kah7SwbKrR7JZV1fwLC1G4y5GKSAVrlO0Be
DVlswX/jmdV+ACpglMwyZ/p2jBNblaa7LCTYPeR62h8dYJQ1tZ6FYvXRs68SwwjXsd2exyIrdGVV
2YhBep6mA51u+lVwV95K/lPZS4JmyURMu7WE8IJACxq1BG02rKfLV4UmtiUtsc8WoAaasELW1j32
ylBY8RoE+45/+KYn+YiOUSBfyh92Ujd2neqwhmOdDs6mb963nLoHolB5LJ+CJPbPYcRtNdbZ+Buw
VYYbF44W713Y/3nQ/58YoDRN5gSDrADdjHA55MBdaF6yaxOL6WhDpPytQjAQ9RRlz8h9qFi6GPSn
zlxqH5YvyL3pS2zf3QJx1ANL4NUiFSgB3a1mtVDUgjzKUzCpIAxpcZ62xHuQbFtPEo9VvPiiEj1v
KBwnlu05XCkur67IjdLmFG1pL85UnGIEbJrw0aQ/SqAN3LeFDeRSvmkOYJb7E8mqqK7J6KxkJZXQ
I3IDLCrTXm9fbP2x8Dc3P32mBYjWcCFMcCzdjPZeDhqP+CHpqs8uIShxgfr3rli1z0O42Zd0+M9B
uuCVMg1lSqV1hGZexOcF4o5j/g3aHNH5/I8nOOI/KPo8UOyoupgnrs0OPE3ujCiLLOxcjusasxQL
x7groNtbupt7W9wcupBdNwfGYqaY5V2WcX0itmeUa0OEgxH9DPLb0UtyBTd0KG3aqGUQCgeJfJol
nyTZtQG7KyanwBxUWjvTwf+2woIfC8w13ytntSAZJbSyqgBGqQUrSSGrwFRuFNNr4x5ICUo4Zgpm
xtiWptjlm6AesP0biRN74P8N3F4+KQ1ymyv/oVIDzG80UhSWAq/aA9q5qNosx6HTl/JnVePX91S8
cmV/gN3loc+m2Z5Ud4OleELtyat8gF/B75r4mytoK+D80c3Nj5hpnxoK1CWJ0ujIUCtb4qmB6GQa
tyiD7Z70pz7UU453ViG2cODq4NKiSxCO7+zR6YHkBxgKogyoBzNADs+QuOBKOsep8SeaKuNRD7Ei
24j4Yvbl+IZsRA/XDln0EWlMg/NcmhF6yWPlzQ594595Md3BahyAaKT3rDlk3Wq34t95+8HOUwo5
c+xZaxmJp2vvpoyWj6rde5av8vXSvMU6OmRRmnVJlof25GtIkiLbSqILgNDfSZwo5CetoK/o6Z+W
zqi0zQWrBNoK4M0TVEjZyyxsxZQchNQ6m4w9RxaFPjSAy4W4jAw8gXo4IL2+DXVLl0jKllLqVefm
KxLC14eUj/vJGlzcjX+ATKoRU0pdR8WdwurXzFd9lq8XQtISyyXZ55ZONaYEVXU29wBl7JAdn/Qy
ScnnD7AX00nxO+cZFiibwLGpT/pnLA2acxWL0uAJNkdamxu1HcKLm2+Y4jFal9oRQOD17XwNm7sD
enQ9ouufFEO0vBetObWLr+2o9U23O8CNHm3I62voVe+zxMKZeYPRShOV1gvh3bJvry26e4DvLkgh
1qFLEXImXHjuVxDk6OdL86tujlcPpJ5HOlIjmBJ3qH4bdAl6WDrg2tqAY90rxm5oU+onyw88xD7s
9Qf+P9HbQnCfEMbKWRxf6IMTUyO4229DVomQhGb58Hbiajnz94bqDDOfHwUnRKU1vqz4M9uQ0Ees
ZrnRR8jw7UDt61eEXtkI1ngGs3pUuU5prTVcA/h5sMlfSMckJxA6O1sNFZWHewSpBXfy+MVPSKrP
W//C0z61d4T8sTMnKXpbczxd++HpQ8T/IAO4I+IAMuqkixLwMVyNof6oEb3c+D9kERlzbYxba5+W
Teq9ub4dAa1qAAvmCIz2yyNZ85WMVa12KInfl8v1Txy6FjR8UnpK4/ryC2CLzlWokrTfgiPZb7BJ
2w9u17abhRM2F39S606idaE/40w6hxS0LJEz1oOth9yoEe5xM3tfvjBgS4TKHWwrvBWLwoc5Hc/r
iYxfOrocF1raBh8hwBS8konRGQGB0F7lLl2JsD8x9xu/8NV0ylMTCGi2PKu2N603hL2DGjcnezf8
zVvRRMB5VSkyOaRqH8sFgtvf7ZFMOBLGp7YQsgBctYmtoxccdirfP1uoCnwnJBKt83/7z9w9iLu6
gIEF2hJHD5wvJFSGpuF8R1aoUd3bWzd62jEzjWiOwu+O1d2qb/99VC1KwxG4uEbr8Bxnf2UQRnV7
vRE+Qn64fXklzBvV029j2ZRsVdatxXhM9+DwDVJ+y1xeo0De8C/4P7lYJUYLvUjbVvbBDI2Ioa7u
Jk68elJbTcJccnt7OQtDc5ey+2Grdua8MDjK0I65xWkWRs5cZHI95ZRsg9KybW5t2AYXB7i7FobP
/URpQZ2IPAQaRcI+gJEytF68d5LgoyQ0vAf0lPwZ1/HFt+TEHY3HB4mp0EIhLpLFUTUPFSgGuFZw
H0mIxamDjKdNdUuHJSANS7E+PzsnOHS4W3OcoPp788F5/p/nZ/SZgzzuZvtLrFufg0H4uxQDpUMi
1+WXwdA5c/feRx8GtPVD1g0MtFDefepu1QUpBHneB+EQC7/iOjWagUpI9GWDP+PxdH/fXLfN2/Yw
uGhoog/p+AR3QmINnTN3r3UxUSGx/MnlDMmaPiV1/uIHNYOd1XfDwj3ySa7bgb+aRFMs2zhx0N1J
7Ko9dqH5GdD28DXK4cbk8XwjSLjncM5oWAj3/LFxP57YlPyRvz5mwna0He/oFLLoAYS9cdxBhMKH
/UoMHTNypUU1qQdKetYVIk5Xlpr3MoqWoz44CG/TkNPYV4GclpWqoDS7u8SkSPfCMd2ECykNEiHG
MkkTAPhYd/xroaCfjU8aAPTDaWY6Ovf119Dm3ponDQ3pMlpP2iinV7kZpmY3AmwEmhEgi+nt8giL
e5Al+PqVUyf6l23V/7alsnepX/8fnLe4CqenwGYWp2Bgb+PKegwARc14yjBua37eDdHprP6diDOJ
tZYbGwoIdVn15XAZjVqVGb5QGm5UhkgM/CpafOXKeaxC9gGerJGFcvCFWWNKSl/JbauMPO9Pxczl
VYggEclJqRA8/N/g5mCjni54yeyKkfQ12srAwFLQu+2sJU3w05JjJ4GVGQFw8x/WE3Rn+Aouuc1H
y3ogZEy7cAgOby6bGrhpkfl0qDkQ/R81MwISbhlTynygRNxJg+sxM1FQcdvl0Qg1vDTm9D2MEYvn
T7GUIhqwtTx9boNapgrbzzSc+eMZSTiN+uZWbbNpCJtFy2KkZQvMdXi2ogIojj2m3IJ9tEE3v6vJ
cpTSYXAiG4Sq6UVO77jtTtKd6KQOsjkI5822lS1t7YUosNcnKEShID4K4geOMLZSkd7WwPWQLHU+
gtulUqB3fN1uVuO1DJ6tVrvh9Nrl4fqB1giaxTv8UkrlE2ii776oYbWK2ykbioKhJhFRapBtuF0m
X0jVUdKEkHvKjFEMpF64b3LBffcmosw2VrE8ycjAsbeLV3Ni8VF6zWTOnUFMjn3mBq37gRCq1fKG
dGhtAh+X0Q+Wa8JgonluZ1kjQjMlhotqAEIVOk3NJGjE0+O93vsG9jCPYXkZeInqUqwdDJWijG3S
piuN81mOWsuY7cNZl4SrnLXg/r3/O8YMWhE3h4biCxKx87DP2YL+QqHvUg0kZbm92wx7twhaY/Gu
0qnRadMvjXENY58Cc8DjxbW2w3PNF4sgBv5scdRSuJVBIcKMRgGueLnkZKufyCyHdtq0CRkW17cR
srO+ft8rLteAv5wiJFaTFD6FCvu2cjKbnpJ5b4Rq3PG31K+wY5U8FxRNKhZEw8WiwdrFK1C5Zcfw
WHa86Zbn0UL1diSWS8b43ok27F8XHN8vC4QoYtzuwPGi3mSzfyNuBFbryS1F2LWvD9xqthwOV7xy
sq1K1v6962VO12D5OtTRSRmrCVGJTXueSXI9lQoMgZOu6YHwctKdGgqkoxVPdUQyqJVj8KmJELMv
YhGuY/KlMzcsE3X6dQKNygaHw60MPOPcCilYkldyFRdfciawY+coxPCePBzhH6LI00lOkxImU2ch
lVPSLSg6foqy54HhAAk8YRmw6g09hK4LrgbveKXJIqSwMnEXhihJNp1IREwIPd2mk4lBekaX7e8Z
hqJNfm+dFh4WboFfGcwKCLTbg4yWN2sWUoZivKh7BbeURr9lGDqSXo27V33kcgzeTN3l7hr+NUhq
TV0o405t31J/VYFzza+R/1scHW8Rn1+pjqnSpzU8QoeSn/cZYDr+6IfcHWKasaL1eDs7dF4be51/
7KvWLtL8ekLmgUzkMfwoOG4JcYT/xQlOBpaU6/Qoi0b/+BFw8CqEZbF3R4rsjOt5NuAmp8lPotFV
/1AVwj6KOyOfPZ3VVZ+szkLWcXvguidJ4gOwGm++/vGQyeMnzKu1U3X++i4wlVY82vuXVJbMRbVE
ou++ke7u9bdIuXFPnsqmMlp9JXKsmLcSiY4ukyUj+bQqZDTM+neJMwLKEp7Md+sDi9Ta7bUW5IR2
qptolUQGonnmWXKf8VHu6TseBtYkGHRIq1z3nNO+NjY/RS4M65d3OwT1Quw0tkqT2WLOuk8zpR/Q
ReOy0VrtsiBhkrvUsw6JiGRMBq/EVwjnFQrTW3nw7KoRw5yLlR40Dd/KQjR57v8eSTaYn/TWvz2/
YDdDAEuqb3kqX/3xtZ1Q/87lJb2NH0z74KBaecJ2mY9676beZK2+WhA/WRVg2mMzBUcxD8cB3hRa
fbohTjUXzDXooU1xYskvbgz6Yu7XNQdjYS6v1fLmhz4jLzGd7soKOailopzD18B+Y/+3XnxluZTw
nICFwDw0Neo+ufMi0SJcfoi+kf9pdUS88s5ZN/rz6B1B8MVQyVG6SetbVbVqCUqQ2DlcYCjipaVz
ITGSma8NlcQS10EnRk/OW/qtGHIzHXyCEhy5uYwpSrURpI8HzXXn3RlGliQWhP3eaq0mj7jObzbY
qPCUx36bk7pg5FCHaiNtYfus0SMn51FoYlzxnb4X3LycGwtEvQ9hkEmL5HJk8cl+wInaUd1zdJmN
rJDakwvWa51tSeEJ7BR089ET/u5WTX7EZ554uoBDobfDQ2BC5zkGb+0qWaONHC60b/nep1qXKgC1
jK/COieHOyh+4q7psjd7FMlHmF1ROfPkjzcCxbOFXAS0cwLYqL7BJH2XhIWq/B9mrifT21VVEsq7
Zn9c1fHZXO4BzfXV5edtUAaI9MNV+AOWkYqvOd+THUyZC21CQgtMxhHir7TEsnTkz0zZRnvZK8Eu
fPSwDA24OrTR33nduAXIjU60kFBg4BO8IvLTlSrspPlhnl0myQTDz1Qtk3i/xh/amq9mt8bHeRR5
MuAdo8uaAU0q4dsWEiFc0cCypMObYhB5F69N2ANy7eM+ngflnrseLxi+8x+dX47vnE/FeLeGjnYJ
t3B7i/vtNa+hUK0SyzIwiTvuzd6LL5MvetI9LODA3lcQaFJbt5KVEe0AhyxEdqUJVt5WmRad/R89
ntf1mch5VEswr938jO0vaKFlMzvb1Eq9sRotSp4RTieduZuH9JbxM4Pjc3CRDPZEmnYjqi4S+4N4
jv39jgHTaMhBMKFUkcKleCM1+ajkV5A+xpx08TUHqqReS8/rvAQkUrWNL9vdyfYDPf+R2ja3y7KM
5gnhWL3K9OTHaHKhs2hNkVdJZ+DRywELNYyS42cK2F2NiW/Vt2rPzZYhlcgTeNl/Yygod6HfGLw7
6HWyFqI3AEJ55GH3iGb7BmNVal6YT0gZMYjIHuktpEbWzpNrnnMCJw7aGANNjmcRc7wJLgnvAVb9
UYydEIgX0eGwzc/BrQ1zKHrYt5CUWUDJ/3e25pVRwuVWO1xUipFn2k1ntxD7RfYvKhtpviRZbjtP
TUUpBsjG4vgOFba4f4a8WGg5PKcNrU0zawN+FmhdSOD8Im/IIhvzClN0LwFkBKJXPpBsjNAlbDaq
VxauBm1eyEBSKccDO4jfIilBnvXgOQlQUTXM/XSAJYBvR/JrW40GYSBCHgTtOTL/c2GpV2tUFdh4
kZhIP24kQw7xpCw95O8Omp7ppkq3oTjyHZ+GFCm8PphcsTCWDDNXIJ5k/kNBDynyYQocCof/UJqk
F2XxX4rGh006VR2Zw8nUTN6bHy/IkQNDcPh22zXUeXLyrCqu9Aza+9M1kYnxIRLkd5LjqNOL54Ct
ENS4Iqee1lb+5D5Q2YRfygOk1bYwAs2MxM63iZOiyYextKLM+nohKBk251kwTYn7akRrbCf76r3V
YgBDxQnqbhecv/nH5ueQ0ZF4aAN+rieNm0iFr90eHIeAJxwmxASttGqWQmzmyQg+iEqLSGOBwNt+
MQJ39KWPk98fjcyyDa0ekMmapU0bSIhoJazADDr+z+TmuVeKuwbEad6jjZPq2QjjilD7gHMBskik
sy5uFKvTMsJIeOT66gyJH1DStckxGtsR4ezwhfsgVNWp1d4+6lgWzaObdaFbfeuEmHzR/XtQHoys
IUcbXFLYygRRwYOBmJhZTrR/N1LkxWeHaVELplxWROn+kgp88yesXZ3q6rBOTz5YzMl00gx2nAxZ
3/cv6RxZgZ5X7kEjN2H1+At7BWPd8ucK/9XMGG7smf6mTGh+KEvS9e/O2aWPlygtjHxYHAMCM0YR
OlycFbxKwOnlCOlSd8/+eSXRjqe+5zJbLhtqoTuA7fkkyh9zw7Vx3uPB/+7zrsfFVbca+EdpKW9f
I0Fkzj57TuFGPHUN8p1rRTKctb4XweS47pGsv5I3SfJ6Y7AWkub/b+XcvoSxJtSfSgEvV3Y2/NlI
n7ZAyKWcEsTotCcKwUj/LVjL1WHyFqyujY/yVa/CRYkwjf0bL8sW40YYv8rplJ1Wfp/JUt6TOj5C
3JilGstd7AvaVa7z6GI99GwwPBlSt8bTARZ7w+Os3mVtzgUH/9v097r8YUl14vY6WK+txC9BjU3Y
VlqCkUz9V4lPMUH72yPwz1LwBrJJpFbnbT/C+8eWD5JRgPtlnaFT7xcOEpsoQoHLmkzzCC8qWHzl
iMMWMj7VQF8ugMSVIWJmBGr7Ncc7BQcCgd97ajf5erwhp3uU7toe9ZR4ryiGqXlhH6c+bul4cFyc
PXErDbjlm7M4NIcolcG7mSDa2LHuxk2zcL2sjVUGJewDYrplD2WD/Nfuh8TorU6XSd6ejjtB6VJn
2GEUSnLS7hBd7hO0b0QXuklNe98Aw7u93vWT3NkBXbBjS3Uqz9TB1vWH+7YRhAOXZDq0yPEb5K07
wik6KFyv4eNb9YvaOZ/qmVq3OhbzPbZOuPdcRynHWTFzGNOsgwF47RDyu4uldthfnD19n8XQa92W
vAZcIrbJlPqI/cZ3meGPynw0ioloYPZ+vr7O1+G5jcc7zqh8HB/PXO0PFXwvGxuNqzv+BmwhK9MM
eJsG3kBn8JpMobuoRBmKfI1irdomNmkoe+PvptJ/UxjSikZbUZmj/HJV+3/VLWGE+fSHtZn4O0Yc
2BGGXDiB/flWVyIt2GFI1IMuHqfoh6u8L4t1lPv3UUiZn/jHYOSk74VeqLZzustJT5uwPzixRyaB
bOOo7TLqDxy5ZDHOfOBraMSvt1RAjkReHvTEESFNAXIesBlerMJwQGBz98p/4hlRteA1YQ5KsmId
BKztdn7zq3BCgUGiqlxHbfDqfp3fT1A1AhR/KrvuRJCP4yvJBG9Q/Ojt8Eij3BXrjmUpesiCcVA5
tglGJjHNd5/rN6BSsdLhxEF0CobX69wFqWTR9ZmOGYzDMyRAqU3lcK/e2Tjt/Tzr3ZGyQ0FcM32F
w4pZdCDBw/u1/zmY8R+Qt1xtyya4c7kpu+YkLclezQOFq2xjYeCRDNC10z+03TIFDK6/ktQm6VX9
82BzxI600fSvREQudhghY1dW3jCNvU9TeLkO2+Wu4y2OXXRO48aJ19E6ovdmLJaHLOyrjMpCWHQ8
E611yS/sG5KdR7T18ZF5tF/rhJgErxWVVyDXr32GPLlqUp+mp62G3ioApsJv4eY1h55r7G6xZFNB
Ir9HYBvrmQICuBz6NBYoFTNBYkTsGZYYSMTdqoTnO6r9IinW5pJWpwuBq7E2SsO9SoHZaWasyZzu
CIeVZ4CEn5+0l2LKbvPC4Mb0UWmXSDHcJ6YJUtlBcrMj/QZW1cEiPczVpEEbmifTutMNNrmve9D9
PwYZQYDNyzHNPBC9Y5irbMavc6G0Oepm9BD74Qn7b6a7aS+TOamBnmpjUF2gOXS2MkU+noQRWrJH
U05fJ+c20/dt/CUFrxGZy8o0YJP/aYmQ9QoL2QnvnvPSmnQfTUE/jeCj0rWrRDFve0a52PKXEDb2
uXzwHyKBZjP8/7wa6eFLCcFQrif1kIKIzoGAydJPD7nP2I4aMUV8B/BLqcwRQIz28a6VqEDcQNps
/Lp/2dET5UWMfuhK2KfcrWwBQ0BkNKZlg5JVfKn59OvrJ6hJcY+ZUjEGPp5PqBf1dOafoAD09D9+
2CHUlzu/MHF5PJH/7hFqD3FOnkg8Cf1rHMCbbMwSCIpBpW1RmRDbQbM3N0uB5VpRTWEQQ/Gk79RC
xO1krCkUsAGzxQ6zTowXaR/dUmP99BmVn+RktfYDX2xg5saHOSuOrUU5avE/h3Vl80duxc80U9O1
DT+mnLKOKoZZX2QQGVKl0djsiQ6LWDoTXLOcaN4QmLaVVhAgX0vRdEppmTf90HYkJI/BZ0D8vTh3
Qq/4G7c7rZzWxhGHH6jLmLL9dCv73iusFi4VIXP5zUn5k/QY/IoSOPK6lDJM12NPr5rWE8hiw/fo
sMwMoT9Dm1rZSsuYfOGmiLeXU1RRZAOVhrBwNFc0lEQnWe9J/FPDbYfNjLBK6A70iU4QCRlqAJSq
+JAL0KTYDdgrRsmSnfFz0QUm5Z1PEE3Mjgra9EXGP7o0CBsqRtD9PAK/7YVMMWoe87BYOTtOdXyJ
Nf3q9Adj+ibz1Ujuv9C3VzKEjDuJjzHVJUwKN15i6LeU9YpHrXLHMwK55smWE304kM+2wl965seG
c/gXoOspkrofDm3vzzixzXREK2LE1hB23moJ+zTDCvLIgp6xx6VDqWV87LC+BjUaZwW5+iykc4EP
61P8ewdcwyOwWoQBkToNyNFZNfdDzXuaXcFtd+Wfcp4qV3oE/Zi0puv58/4UL+7eUmcThQK/BngX
7x6ihBkcSPkqM3GXw5vpAFmtbVEvYZ/LTccAwQ96qrZfeQmIkA0v64wWpohN5imk+as38ZPTNtw8
VaT+isVDBVwo1MbAoAUBccCFD4+4pXS53g66O8cFloKn2yD+cYaKSz27hPNRhqya3ldJJMkLxCZ3
P48fpzhGgldvj4BhKgeR2rPZla9UkDq5N/DRwN0y5RBxFleQ3B/yGzIzH4Pn3BUYTOOYml0/evSI
1OCPyHQGntyk4+rkubgy1Pv5qlp57iBFhHWxrX1oBv8+4hi5eqLBiVVAuzLu0xfsnsh9tEC6bvfJ
1S2TPIXeFiel670hEvNAR1g6OTH8xG1DfxrYCaOX0Ja91suKXNCc6NvGmVkyA9bFvEnpd364NdZm
8RX6AoPz3Njl9Hsdb850pt4nv5mwlzPD2GspBFkMsvzZbYELiDqmH422RBSB/zK+QTdeiD2tLuBK
kxgJwN93WmRKZrRLWfAUs0Su2jjGwSMMkUZZizXjcNhVRBVdKDjz5uh40C/0qFGyA7c4yZKzVAXe
fZR+hOFMnSNGOZOClV+jIJAFbEC7bwwg5tK65txw87qHXfOjkpA/nr6dAj4SUFk4jFpnZrVZr+MT
mcFLk6q2yl7u5fa4qlULmf+yTmSgNbmK2KFEPAe0eDsVxafWa+Hp1kA8PgzjRQ89RkqvZ6MGt1+Q
84gS1HchSZ6iLcLgQ/DzuY9aqo2JSLmyYcQV+Eb8pyQUsq9mU/0eAS+LIM3Dqjf+DY2TX88CbN3K
INm7hUVNpSiM2IBnCj0vmvajABqyNg+Jjm2OF2R+ty4wbtNePDenC6hELxdMr7C+toKfqwr9OidX
Ow4JFbLR2QRWy+ZHPYf17FtS1ktOoQwhG90TnFidBrOTRgdOSoGF7U+v2eKbp3ZRzuUL64RY1U93
RyO5t8wNtLu9z2D/IWudpBKIxQ6OUAfHS9bdU5EkxAyr8VLpFtbqbbrgycAmaHJVoKzpWeQnHFQT
Px8hhsqwrRDo1MSGUNyuIGtHYA1q2JKm0az/02E0QI1ugj7MZwvBV/TowjPzjdoLmj1rq2EJvXSx
glAiC8t4CTdIa9g/MI70tSGsDOOV/Bd79wzkEYFGIukwaGZ6wGfxSAVqdROdsAyooY26urBe8hwp
wKFSrDczgrsl5oGCZ99yiPF+I0OIwXfoe1+lwkTwuli7FW9eWocjO8Hgvb4PnaCMA3WSKedLdmm5
IOhs52wWXe3FeRkhsIikSWn/IdjhGlEYqIpuG832yJURtDuNi/n1hnFLcbgESDBfez26ARXhZJvM
+aOZolrK4BN7GE0nlBKJ06TvqB7SlwVKD00rspAEuw1tlD6C5aBoD/Aw9IKLbdLL9o412gDQyH9m
wju07UkcCYDWn0yqiISMh7BYiixtYsAefjCOU9Hm4KBudA6iCXlkItY80s+PkwU1xPLrNsZjrlLY
z7Q6FyF0kE35fUeg5+dwzWLVKpJUHQdAgW4iVr5k57kjQ9Qj6C0V8+ZmwfVhv948qX/ufTJxZqAG
P4EVaLcWovmDgiyJPe4MyOa43K3UHEiEt78tXCWnNZUnATniHraKtTPVqJ2hWniDaowp1NGPHnIY
BVAnuRLxgKNdUTRnOoeykSN1K9n4evtfi8TRxsE2DsOu0Ll5X7CRswfFJaf9Hs4ESxTyPThD5SxK
b3fHkRpv5pCgUZwFEMqeshltLg6HhO0BVBWt6Xi8Oc7rNKFICmFYtfMTEQD2N5KX1Gw9N8oz0BHa
KtUb8KAf6yuMCe2Tg7rZMs+eQddvMuZ9a0x7ayb42KOUj+tiBNfT2CwKyTt0QZxEmhgCeAFGmXh7
ikPbwJgpE4KsvPPHGhlY8TRgFCpkoLweb41B1E+L4dzRT/50gxYo/FxlRBB5/8tamGsRmHy35QL/
4o2k/eehxaPA0E5TLF9/a8r0Z7PjrRwghZ5vUMktTvekrMWv5OaqVthlGPZ9KulnhUT7ALR5mrt5
ugIA2vgYnV3TVGqbUhi3vbW4jJKCmQ9d+7m+8U7GHZTPrzBJf3/TdE6zYP+82mKADJIIYcQq/lJi
hDHA9uKPGQ/nehkyUcE9su4e4yc1eFoCcS6zbUqQVGZYNqGxrwbKaCDl8RWK/FEu0rlh+rXotc5m
Oetij/6JE5NUZ4Hx6FMD4g2Y5zMWYmcS0olsuennphEdSHFWLWbR60Of+kXSu1R8/onA1scWsjk1
bB7Nhr2nFqAxi06uXzONo3cIs2mTKgT6Mxrj7u0iiMsoc5BjcBdV2VTp/IAFz6de3HMlGpzGy61x
i8KSdCEui90ElyOB5DwsbmUpjYZyQRH0Lz1P+BA6WFrET6FFmY4lsAQCPV0q1fE7PTli4Uk+x5Sf
8i7CgTLRDJ2g5+qcTxB0L+BXJDhbrYMPDlNVq+aculBaOXDstA3SUvB169XWQXUrJ+Ro+lA8D23x
Ax8hFHT7yKg7lwk+qQvJq48UTIkCOIPoSqymrQHsle6jX7vyFqMCj1tLCy3AdJFhX41AX8gz7140
F9fP6RVX0c6wD7drzJ2LuQL6EPnfl9I3ExOZP7E0xKJxLJwXuOmKHF2yZD9IkcvYrWmEFaWuRBAw
3wtMi1AA7TKQQsC1Jd82fv21TdIS4fWLZZDc7eplM2FefZ286r+6CdaNMnyNV+16n/3ecvRfK5CF
1BQu/1HBggEAf2IQofwXBOTcQ3O31ZkMYymY+Nbw4layU9ixkrAulloawbt2oLc2z1vXM9K8gRbm
7w6fMhep1jrwWtPSpSatNJ5uTptm8pRE43u1YloT9L1NR/qXoXW1UrNWYS9gIFl6xGTAVurG1KcX
stPwzv4CIKRM161H4GhaQTsbMPM6Q63sD1kLrtgMZMZfbeEfcivFNQP3bTv/b1WiTahZF+r9oJCO
x3J5rBTWhn5n0pAz8QBPo7yNRJWlHedu/M9A5Cs/3Lcr+o3IpHHe9UeQxbSXtOmwG7JKGrfT7LAO
YijkuJ45ppCPoO6Y/hIASMmnp1+5rSYntN6hGi51QV8IjEA0kTuep/RwSie3Ggu+/Coqhx1jVstD
nPvpHM0JOIokhTW2VEOFqwrtvVROanGj81RabOjaRohK9vp7f8+X6Qwy/wc/afjchHTZdCVYmZHH
aETJYM+fs3NuQOaMS3LF0xAvcUjAA/QUgd2hrl133w+4LgPumia3qRld0zwmTDvkhIBVcESH3X1M
L/+vVrLf7CmOXgehOXSJwhc3Tgc/n/0ZnOlpnVJwLQGOgX6hzjnSE41Wyhwv0RrhZCsw16EfNW+y
OuI7sGTTXEygLHEYKy49rpp3SkOItbA5SZ1Bi+M3ADYbE/oyM4ye85HmX6ZdbUOK0AIHL/qzYjgs
suqotzTH8cnUGEcG3Yn8h9SntDGR6mzPTbRJAlNgYuZKjSb63Feefp0Gh1B4T2UoLjdY9gw2hinN
v10N1hKtKsqzqhBvI+caudzCL9QejTpc1B7ehSC11qiMuzhCIL+I8lDxO4HzK38IT+D3VU3KAz5I
odRGDfKRSoHqelsMBYrPcJjB4EYRM2T4wj20Y49nHYtsvyxZ+RGVSZk+jr/3ebjfEYyftD2JD/LH
zORje/cDG+l+/tJbCMa5CqbEEgwd55R4PxxvgnFY++8wjpLgKF5Ukp5cTj8yesAmGaioMLP8eOR6
jvj5oRLjQ7IRGPTbkvk18ifsaIJmA3k3glJJTFWh9C7lbwzp12qfMcMr2zHJzH67r51IehdQaLF7
+lua6aiJGBkgt30Mh7BKF77JhJxo10z9ZfN0yPF1dootiBYOUQ8f7VeAFSVKwmFI2yq7aTSsxSwS
govt2p+P7bjsC+4mCHaG7XNMAwNiJTbWQboSgGAGruDNLOcUNXxUbEUCEDcRCHa8O89e63lGGzkO
Q3n7Ug+eUR5uV5W5NRQ4itUvECvickzkAdU4cnftWk2P1zCOe298eDbk+BaM4K1oH6DVHSki8yyG
zfLWUPmxsAH0gnJQI1vxqJkQkEoNaF6nHxcyarDERGp7Evpuxf0blKJe9aeBGMTGP0sp4JWrgvp7
H8ia6NQTyjt20C4bAzl8xppGkyIr8G0Uk5BFB2DwwJklNU89+iAL46DoWMLZqHBrRmSBsxYF97eZ
6Q1qfhcgeuF6NzoP3noFp7Qu+VwuJe+CcLt3Ie0XkcIfjC7fYxO1KE2bWmNjWeO8mhSeUst7v3QZ
hXToYNHh7cCoiIA2YW3HdV9JY436hHr6qI77AgrFLicsXTrlzJL+gd1F4je1+LMgyUVQHJligiAS
A4ysZORxNz2qgNJOu20/4bcelJBuM3UCs9qT2Ar0yqQ+295hiTrig3Z02iEeodNrhb/JDvdWVcNe
k4Y/N+ZNPjeezPvomL2pHceC+uCvcpcZqv4cL2A8kqyZopVrTBf0bJ86Dse9fZHs5dlmwWhxB419
mEgqd+NwhD4mlzR3i/Hu88KiG+4uZjGhe2S6fsqWbEBme++oCfBAOGiPkGjaJrpUbugoMsQ4eE1W
qqsSnz4E/sFUsGVmr17DlI0rJFKA8cMgexETJMl+kGPz8oG8QQXuPU5lNo/ImcYZ3ilFsBEuewca
i/MZzBe+Z2Ze7jo1DH9jP4wxA5Ze2ST5tAxDSh7cUpjmIPHgNzbCRCZ6ct2NPMi36iwU48EoBxhx
bXXRkZWbvyb3h/qpJFzRyahkeyWgw1LI/hrakIdtloK1jtfgT7Y+ZKLwip3nGGNzQPD6Gb+MfNNn
vWij1YkK1yHsCDVXb0JnHAoYGqVsu2e0QlqegQ8d8jTH92QzFzqTefPw2YvsZ4u+iyjLAN6V98rD
nL7BuQawzbs9tCqIDGmbSiWftpGOKPoaxqhcefbLVNSFiAF86Mtv3d8LLTTp+r3mHjwFohmvgC1/
VsgyGCpIbZvI8Li3zc39BcHLk5Mzqs18PgagiLPF+qibPY4ofXp9UuncWp5XMmQXiAHT6xSRu2P+
lwlQebnHw2/q0uU5v38M+SYpgSTAZzK1eYGMcpJHcTH6u3LT9mqecxPaqDQOGzZj/f+IrLtRDkBy
fEO4wuZVXOOz2i1WnnTgJXUx22qSsneNSP+ZZcrctcFXNQZHutVEXdFNmF8PCJjXM7FKfX8OrOcX
xyUcJ9PNvaH0bZOM6JUOceXvjZw2q0UGGtaIvuyKJ6tUJt8RHWi4rhAaeIWhg95eu1PGzGY1X7jL
QG/hVkJHMJa/KA1fXN6ht13uCBS0BHXanE3/wt/Q01yCvBMvYwbNwUsUb3kVeaMF6nTcHkHmBWUI
Whfmxj2Th5sXWq2AG399UC21lPhEz4uDUNblmaYLQSnC00m7waxTIAiicJTWOjfox6ec7aV9cNxA
y2VDMPTb85DgoQ4vaExipF5uYHwUA/H+Iv0UQXpCAcN42Li6tmtKsc48O42oxx7oi+4NCahnZW5G
IGwnF+GbVjeOdkvzCuL+PPhPaazrmoMlreIQ/0PyiglIylD3TbQ0J1XFG/s/y9qsMouIXeXxQmYM
/zSvMz5sMBSymw63Nj9aL14QSYaIOq/RpedWkWmSX0a4WXMZDHIui239ofPPd3gpWCoYGCeGTPE8
qqATBAWbKzrcll9kF4EFZVbAouOYD82NhRccmy24IYxz1vSFUJWQnN/KGO9LkrX63sBRsH5yOWUA
YwufO5wz1bHQAzG7fgKZKAlll+vhmiWojMR/sFjcGzkH3tIxFULKQMNTxiVmJqBqW2Tz/KzCp4KP
FVqm8ZCmRwf7pH5mv5YK8U4nm2rLMMOIQUgg2+sKBd67/hKkr9KcFHClkujy7yGT+s8iY4ZnMunj
UOm0u38kszSl48ypMSExuTenxum5yKW5zXS0jvomHT7NqdE8oRun8jdGUz78yT/sZcIiiSYCHhir
pmHrGIIDKx+bbRfaP6gjn6RMxgvphLcUX8V3CxLweR/pgJMGmJLcGqv4eq+O8flKxg3VZmk3rzaF
UWfksS7sCsSuc2cmMRtmMXqmhpBsoUnBapOB7D3L5qNXllxkrzhH6AEAEZ3TBxw/nhOO/7E6AvCX
T4iE1pRS11BMZAiBzuNAsLymWksiyfzAG+WAPXp039WVjI9gCiwCu+wpTHQecS3BuJzbAXFWVoCY
kuO1ZFKZFCCkj/QpP7esoTgGJx2lFHqi8+E3BRhxL3QmrkU1lKwHoQbS+FSnxLCQ3a/NdfRe8dsW
S/iNrZ/a47cuUOmIi5WCw+2iSNrbnBFmx+Kn+SNy8O9X8K1wt6SK+3fHQTl/OyXKD1Uq7BGl+8+E
3Y4I5RtmF9DffY2Xnr3x5o2+AdUcGXSPtT6mhklgJus/pet/KCt3szxomTZUUWrMa/b/b+9d2QlZ
1726kxXOBesIaLfOrAYlIW8k3RQ/zhv7YEAry44cVzOxiSu2TjIv0Lt/IlFgIryXHyKMzI9BwXfQ
w+6jM8IEfebsoWtswQCgGtCSrq/9sdiTr1hk+UHHJzS0GMN7G9Za7WCPDLeBqe6zYP1eMkmfpebx
kDZxBU5l+YaU3HcsPoNNHYbKNFodb9jTynAJR+QisRo5tzp7UDmqED0utjtuSbbP0cA3aYW7bUcQ
xvL831C5lHfXnMqcflTndmZvPMwnX4pdYxVTxZR1bxQKtFfFMiwl5T0dgveatDD/vd9L9X9j9U0b
QnJryuPJODe1X1zNq1cHhTdgBqhZRnpEeatmwdoSbLF5Q2us2a6UfFJPWWFV0LMTNgmNH5o7C63X
EH/jWqdaukWJ8VTGk/xlfK2jhLZpUPTrwMJof0HzUnmcAuzVGXVcgVCxxqvMwX8RCSCOPklQJvEf
wqFQjKKgZB06L6jY8WvIxnb3Lvfym9FZerQdQfraYJU25reUyxeXbIzx7I9wB2uBUnHJamFDDIzs
4b3eQQWqrIG5T95/+X3KAfkQMcvwMhoPKcFiAqw7U29RgupHWn25cVW+Aqhb5k2zecaHU+0+8mj6
k8HBudfPZENBsy29qmpYwwKjian5YbATsmn7Cj1E2vEenvzwvNQ2GOw4YW2XtJ8BEy4Yq3lx1bSy
P6KSXGAYyn9YXwqDL/rpoXNYgI7ucqxPX+HKLF+uJ1H4YeKvr/4GgJXKWpusdkFTGcgNQgbXEiv3
kLk8rtINwKrzlRofHjzL86p/1qYzPPcJ9k7dqLQEUafHngAlOGUsqFQshsnXQ0I0W8f3dDLPHpHk
9aRTuMdnbs+LYZyXn5Zvdf34hg3UtnlFFKvU02t+dDBpjgROe+dqhLOaN926rrgPBkf5Q2dNXFJS
YvYMyHPr9yVDmDbq7Wa6bECE2JTGg7XG5vRmNZTU7gW4YEfADvZ5tBrVE6KOvMcWN/jBEvH2Y868
j0oBBc2HIOWcJpF/Up95hMCOFc6/pmnUyfCS28bzlGOtM4z8CtR8ZCkTsRTdtF/biJNNe2c5X1Ha
C0WJC3lW48HAlWtDksm04Vnl03ssvR50xsFUnAUkf6ou7cs9l4v5EOkRxg9bjCgFQ3J7GjHFZUBm
nh0scave01sOYb/Q5shwZpX4doqx4SLzBUqTpE/YFipaGIuU2FysdHqOLx7Fs8FdqB01F2wctJPd
bRDlYWZF94jTRVNWNAdDLTppiOf6lssPJaUwkaxVhnoSuM79BzjRbqAeIGfxfx0+LPyNLojFqKaf
D2yH9gkGQECYX/xkoHU82wtUdYsun+2GS+yZJTsM6OFfQH4GwYSg8QidxHWZ83q+SF+TFtZBJd1L
hXCYDTHs2osHgqyDq9QSB6iI+81/Me53hO2E8nghdY80ZItO95pjhZ1In2H0h/wteTMVMhXajE96
mjGPWqGOPz+/byt1F3sa8mAk9oj7A4yw3Mjc6XXro3ZAeNVibCWQMp4pe9XxbOncfCRtSFVWvwuz
FacIli4Whl1fc9ZIEIE4xqR2cTsiqMKGn8Ubm4hL8A+2ddLgflvUZ4nfdF6S5NN2O7WVgnHtSRFC
Br4Wa6IT7ZACtZtjOpXYRCRcoaGAe1Ed9Ta5E9kQbm6pPrwriMGi0E75g7+h1JGzrUs6F3DDhdI2
XMXVSYePI8ij3i8CprLgsX7P7a6scyb8Yx7x8G5wtTusIVa5AStzLu5eNv6hIYGv/e3lcqYTycDq
orKjJQkuFTd0wZOr/tQlP+6n2QfKjQ15AUp4S+Ml7XxNYhC4JeSv16ZP2Yt8RzeI8eIjmIhtd3Mb
KAn1OT3/Kpyoh8r4ZsRcQq1yOIvd7junqbheYaBSFgUya/49NyiTO1XIU3+oWU7BNxC6UJkQ+msh
86D7+u2SyN0n2RROhcV9uQwBO2dGJGZ65bOisNnoHKAyz1kZ9NgBpKvFANIaI2q19gfnGikMwMGZ
bv8fGCrgj9LFUUqKUW2xi5yxYsfsUsVzpYlV3vVkwxFy80aB5imTN0Gvg+88ZTFao+H/SFynwZ4f
oXIWiTKt03RUD4y4i4OCGSkUKo+8tn2NseKtTVuL2njZUm1PD1DLVW69/8i88N0sm7vhT3s9mhiP
J2yQN3WH0ykjnYdPkOSO+/U+kS3x1ZNweHAfsM7jRts22drHDg2Pvltgqpe+E8yC+G1Scul6x3a3
tCPc96hQ02G4je8TnAJ+peam76dtLsM7UcPsDTUgmRe9JAiUFMxhkoG8Mjn4Ge/Fgp0tYUZn6HP5
FXgZY0iLFIoFzGlHeLK8UE1PvSl8MJBK3NcxCkqIMxfYxnlI2hxEr/uTKpmIQg57fO3idCLcWOf4
Unn2x1jfUb0RoVYYWHLYrqmGqVi8hg2KYc9u3OeKfo5+8LMyeusTl0/Orzer0HqeFMBKtimaJ663
it/kbV6vl90/w9shrGHFoqn+H2aqTJhqxChvLQ/n6R+qXjCmYlI1EiNoeq5TK7DgbyNi5AtRpJZp
xmFWj72k9j6S2k1xKgYODydpWesvJukXtfTjUCvl9QuSKqtkxxyjtSmFGl+9ChbuRrx1cp/J11P0
cU/nzohy8JpamsD1c1ymRkpytkkuZKLSrAITHeY1wSg5kzU17zb/t5PTH/P+gACji4Nw9o1c5ivC
mAd/qOwaT6yYDHCctyOpxRLnuia9cUki2+tgr+8ec4YkUJenjVZA+DB9akBl4KxzsPrRr1YB+oEW
Y86y/BbhsYx3giVLTjgYu9TlUsmAKwSAilzyXXf6eS4qgavaFGOWHdUvuL76zg79KSZ1+FsjskIn
v9FddI62qM/xdxdyC4ygr47Ol/kmNW68JXpdpVZJnyFa+U5DjAiu9+GbBRdgVhmO9D+fMolS2ubv
NS14Fm4o7JwHMDbk9/M7WA+pv6sp2d9hivZ4ZR31nI/S2LYwgCXrgV+m2t/lfynHk9v3z4tfnyXN
ceZMzzMhsdG5Dm7c4yd3Ht/nnFPODFRiTbPE/HUw6RFhmmFHnvV5Mf17W47B8XGLd00eU5u+iqgh
UVJUrcRtn4oWX8mmWPrjIkRqOUVY6Hrp2f6vSNglKcOivyxylsQZ7qE/l66NuK4WSy3S0zQggUVm
NFbZyEy/fG70ArxBf49y0+4nvE5uVXQiUHnZ9d+/biECfq27vNbxkxn+HkxbDMCzy7H+XQBRAA9A
PEdfHGGIL9YYArNXPDS5juUT6205AuAk0+nqyD8DjlNtNIH5RddHJ2Ck7ly1EIwpjA/lH4CMyuWy
CTsdMAs89rBmjxk9aVC12KXIPntute6b+7NqZ8ISwej/6NpzhujfGb6Q4YSnVZBUYlPE15l0xqHq
YkJtfsPiquVjs+/Cr2YgoygPUrTf6+h+6WNSAyoQCwzRCts/2SCNSTMnS8gFaWys4tIky0xVPDZg
WFmLJPla5WArm6e3puaZ+cJktfFpo1DhGLJ5ROpfrH5AdUZhLiKlastKprFHrjd/CcIWMgBpklaZ
+vkHVgOXv4TWWaFrJQFORVMnNl7w6mOD7BlSxkuEX199ySaEgjZ9W8JeuUtfz+FfdotT+rwEmB/0
1SdrAcdmBK4dbdjvinfIYd1lLZf2AG0huyYDviIorgziGOnSJCZGJj2JI7WAgJtOl4rZp8D/Wbah
KSWozpRSMWP+mV4ZKdBzpuXB5vGLmXmG4rGWz3FcGfxzMpw/2WjjFPotb3csEFW/Fjnf6PGCQZ0A
JO+bC8GCwcHb/klhjBlePDL5SI6AGLAsZHWZxU2gw7d8Z7kmTrbi9CMN6QpMf5vaJUwjb7r4atri
kPPfRL9GnFtO+5DF6Bhw0zsV+iZTZOGxFMqWxG1NFbCrO9+pBN0EyK8FVcW/x90f6VcAK3XLafCU
J24ePVkSZCOsauG9d6fAO5X2fEA/5WFA1JMRfbVE3Q5JkpZx87BQ1B++f8nBDQSVjieQ9SeC1ToE
h7Ooe+N9yG2U7WH/PDw+1/hG+dTviLQb7yYvkQSfUG779QKfRgMogGF+6NXJgXEe5WPPyoL1s0zO
mgD+7ZQR6FbS7bQ3pTucOLz9wQgupK+m9+K7a2AGipcqeM6phHQXj7j7j4oTTLdovDCyoKjCBsoG
+lS6/rF5/B98pQ6tvuF5y3/NxfDSzCUV0SbmamiSeX49uVofsyU1w2YhNShcEDjeWKtUwupdPmDc
oS8PTQrf2P/JGmU1eq+dy5Fr8RgldGYZrWVk3y9unMFv/5o0ZatS+NkxfE4leNgmfS/0mlvJsgvH
xZE1tlCUILTRFzIFz88Ps5lKPV2CZnOK9kVQaM6sUMLpLaMm78+AebK1r4XG/YLBhOf4bSkW0t/M
SsWsPyW+qd2em1HsTHvGbU8PWIHO4AxcNYg4z1WXm5t1iRMwczjFpk2G+LGDM/kepQz9g/JcFNJO
jDd/2OYLaMihzqPRfUSwXWbDtlesgdGL/WSDs3bBHYzxLbBLXVhgUvkYOcs4JkUiBjXZj9sxh/va
XukrUfNPIa6hle0RuCfzfHOjxAmkWQAxJ7Cyu/8mS4Ix7CwVy8dJ/WXec/tIJ/2bO8i9TiL9m1tm
FAwhuL+d//sMUvzi0ICF/D8P3Hh9Ts/Rg8t9IoibrLYvmIBBFP9oWRYkBFvIKI/fhhHjLjTgWmcN
PcByvDqa9X6XXSMKiTwARCsjfbPMoAfhVhsiY0Zq/T/vB8NpduQC0h10J+rRtOmIcuxjqw2jR/R+
WdNrlWEHljdJFpIXQjVe2jRP8NYJ8/VmoOApgbiqP2b3g/t9ysZjSfi0KxFkHjG8uHu5mmg/ao3a
Oyquox797Ro5/9Oxh9x0VfAnb7NdTLG8vBVUQ7ncbJg472UNlGvNhxQnsZA7nFecXCiywozhC8xL
n6OPyssoSkqKzcr04TrKC9EQL4NgDWSCht9MYWTtHayEhzclE/4SYsfm8Mmbb6MJwdLzPn2VDR4f
X/vtourZ4SfPqDDCLeFaUjzXmS3+HRTGSIIRR7IgnSMVRVpB0v0vRJSdsnzaoOvyjYWRgldw+A/t
Krr6wmfki178bBb35o8eVC+sTDSnkozxvM9ulEoFU/PNUodnwCvrNQUqedbtI2KUh3VmnLS/5RdY
nJj4A1VXSqGV0ik2/lJmukBEiwJQ6ffV69ma/vh5q5JBsDabrP8I0kQO209ZvE8a8RSZQXBuZ2Dy
umndSRWm4InCM9bfeK2X4XGxR9nFS//MvWqRCJHHjkd5Lm7dKYUtTJyHzbzNbQzVPsI2oWMDOpyk
CIjKpX0N+/h7HIZGW9zxuAGRDxT2vC4RGr9pDsN6GSEfZLfrntIuSnVJ3UENoz43EoMnB45IplsW
tjhgGKxhvFWmkS43xaufjHCPSDlkZ5twaIXqerG5PJACcX2DKHSBdsGs7zESSuhfUoGBqJ9wWS+j
wlVt9PFrFnnPcH084tlMVqiXFPKteyw/I3wSdBhLr4a759v67mHviA4faJejOisC73BaHbQ+gYin
4UXj3wBjjkztYV2zj+NtM0trBKgJ+ALT1+FKhT4irAk9RjzRygO7NywaSvclGt0l+xGy0TaUFuj0
rWkQeOjVXoZAYCQj8WmXVYiAvOVEF8X3LqAzbVDReNG7gYhd+hjh8fOPtNXlc1TUZuW39vpBgJVr
41xbEEWY39FvpRpKbA6BF5hQL+quMuHi2elXI+dhfCO6U+Ex63HEAafzq4hChC7Bji4ZpvPlhZb0
WhMlOKshO+zF8iNgEHB46LA6DWDhjz4qes3PpfeSpoK9o/xsFNUJ+G3j1jQ91EP2605NRGNbMhWH
+yPghDZL81W0oPfoPqFL0dHBMM3KVntkp96+9XFQKecC94d9HuLYF0X2DcIflWrcges5aB9d4Lgs
leeUe2J2RWbYpKGjjQy9R6pfzYJ74FeDHYHAHBAmyBchgawOvTHxzl+Tus0yBBCPp08VnAB4c0gd
0Z5fFNte8MwEvoXSx12ELKWUeB81WN3NYUPSsptfEG4PdKDaC1GJRdjXc2RWrIZY1BMPkloggdgu
88h2q5rQPlin1GgTLk3b2gq0R1iVa0mhfzHNwb58cmCxvS1zjwwXojU/d/JoC28SaRfxjA/So0AE
+PM+nfaruvxQ4oCSsW+D7C+u+YvKqlaMfwwbE4MM7UCZn+JZwCkjC1IX8p+pfV5wAei26agrmLXr
kjBQ3EILA4dfArODSNUfi972yf9POE6ULxx9h3wv8kYnHhz/TXKNA4b65/ih9VSkGeqiBwbSCbGX
WLaYqFZTdzWRkr7EE9vakVUg2D5TwJQVnaeJeB9mMBD/g0OHjLPZdmpMFWTBMu3nAakZE5CQJ4Li
jVDRKLm8Xo2n6WKVSYqc0UXqVpVgxLAgyvoOVXTUb9+ErO4pxPR6RwXtIB/+0DxZKyzr97Cj2VeW
twFr2jK5ciCO8grnIdLx9GWQ9W9cqIlPRpzuGcpwyYCgD2OUjeFwnOsq5rsg8NaMqdT7c98mWIpB
TwECXSylseUlhryXWRtBSVS3fZIpH79mab+ZUwER+OOzGc0islVzw2f59AQZye6x580oH8dsuHdm
4kJnNqRiEXz43fN82u6gIVZt1cK7pkLKgl1ctfKfbo2Np8jA5Pns1qLLCUTZWxryzvL7W/aLZPns
900o1Sp80mjcJyFGbc/h//qpGewLnZCs7RBU4ucGCo7V4Qffb673oYIInW0kHnhHrWqEOeE6zIsP
ILghDifE9ezCXnu7zqN//I1p2hkfON+ImBfqwJiscpLni+S7p2rajkBgKaEBxvLDazJL5iz6ZtDx
Ldss2Pb4BMBnu8s5364bO8OinswCjAUJj9fkMSm3Ri3p7L0xsA6rP61H9s9UHi5/0ZIFFIxJxY8s
5wj4Ztrt5Le1TPSzWP5HLjBXiA8sxB6+tCNHrMwUaFHnPvp+Jl/Qt0i1PP84wJCiLZVH9+XaWqhj
zuisqR5ZHz/1XwVAbDdtKeL87GgTO7yjuHkTHeIzOeE4HCo+mzmSm22Y3a4/UxVZq0hbzoekFE95
Fp8JT0aRkevvZNjaIG/K+oYCNGEJ8pMVi9VGf/JBrlDz1ip/ma/TMHeMK8pveeRXtN+UNRo0WTNx
8iejEV8bHquDoO1ebDAGx2NYHaF9p5RAydGsp2HLasApiL9C7LGMWxo9Ca5zp2EBdIfRr7TeMko7
g6fVObEDPJ33bikFUj3hsL7s4n6BeHa4eZzkNBxLPMtEKdYunvL+WYLvC98WBlHX0G1iszUlQYY8
f0262PUhH13niYWh5QvwHoF8LJRldZEXugMpyraOYqvk1lacG21wGs7nifDnRKBx4OYAqgWkg/GW
fhnQil0QDFvg0cXpLZ8KACNIEXCBEAZcKRSg9MU4ANblYchDHyJfke+A5VfO66GXJcb/XW2avyUI
8IS+4XNu8OLUvwUWHIo9U51XVLORHRttD3jhvpmp9yHOTNobbxieCEJClm9eZdglu3cYum2jSN87
1jrlIgomzvKDIveTZ/Zvhzxeyx/iGTsCLjwVDX0JfkBSsgEW+U9ZxGiUOt7JD3XmCOZ/JV8YLCG3
6lRKrKzjmpdgcNeght0NBYsFSws4IfcXDmy8T+JLBwCnE0YH5Y7z8WRyCPV22hjKzsS5gZQywAN0
5c1AWMZSaJc5MhaDdigpA2aPbGv38AtZm+px+FCX/HRRPY8V/xx58Be7InzyEuFJnZR+Cc1+HpWP
gC7CSsPHfnG74nD2LJ9/d5rf9X4fQymkU+9/CbSGdjhcGX8z10qm/V9I+vzxz6/vg6T2zZedd0OF
dlm8VlwqLxElNi8gP4HSHq7MbVSko6DzHWwLY9bTfV8c+RHvtMXi/m4ILBK3o4rZRyOW7pG8qVQK
vpAgIcZdOici2xWz0n3cMexdq7chvrev76rACLzy0Fp65DGwMbjemsRmoddgoSxrW7Gup8LbufgU
KB9vnOa9OgceoCwIxxPlmwkZRF2uXxq32W1yCQVXiOj65t02SqURH+/iNJez+75EZAeg2yV3OkS9
wBJJDPGQ8z45pd+ZhlAShxh0xjTFK/iqXdZ1mpe1H691hQ9q5kES3jloJr8uGh/xryRNNRNntFKd
fRIGe2yV+luHq6ExHuamiaErkreJXddTZ9ywD6B8qRSHiF7f268rlYJARBvIXYqUMorDM5fHtEWM
ozGKGhyuvT7YgZcvhibRyk2T2UzIk+St5qkzldY+mjXsqlP1AglQZX2iDZcjYnwXX9NFu2lnIR6r
pS0qIyROurrJyv0OP2K9a5DxVZwTjfFpj4BMYtuoYd4aeBgZOCoVzCMw8DfncciIJAaS+++v7rmc
ifoBzIUtgg+TUH4WTfWH8QVVX/pQ3NnUzIZ0HtTXp1EqWEIc4SyRab4j2S3UeegoHRpFTgVxix8i
BnjJjwoQaoydq5wWAs00JuPLji9J7j7HEFnr4jKZJFooHMWwToQ8gjojgT18VhL1gN/jqNEDes48
/EGvtLzErPTzxtkH/xCo5UM+g9Z6PemqgfUVj625gFNsS4nHvuES8Pk8MyhPGnToTxdFVFkjTvhw
I7zHgPKLSvRWLrfNarQpUIbYxA3bxFutkhDOFZ36SfQcw4iMbz44zjFLTQ13OU+PyPyD/Jpaz1SV
Ss8bp2NDhcaPXQh0V+rx2w7Z6mm537xmmL+067bJu+hl5eQq8XZV5p1M969yiEgeUSf1iIfe6Bgh
/b/x52t6MzKSaqp5sb532URItrPwDuUBdhh1f2cBA3zeZGiDLKdmEC3lOyLIye31+rtjw57C6PpJ
MLEm6WjlLQsVhJtwtD+kChULTJCFIKUl06rBwv3nZlRgpz5n7BQwMokjvgjpnjenA7dMdltxi94Y
HEjUwOQIkEOL3tdy7hmEZf98M/0ow1FF84hzWQ2MfxMIPAUsuHHW8kb7ShyXtcQHw53e3XQjiXNr
++UaqxK+6OiOD/WItoJi2c6Ywe8A60zidHMkYhEbqdIrlbG3YjMBHVkevANiX2EhM0QV97LrsC8j
O1ryrw7Q1a0f/6sq/TzW03XQH4OVul+vKLlG3WwZ6wq8rHgvfDf0EbRw8koR1B2oXLaSGNJWni4j
aCoRr1O+Gqe1gE6i4CaShhnQfvfy9lGFnYJkv0G+9TjhzigZjDyxwHZDphDNEiznxiq1/xlQY7oj
om8+Vy49uZirpUezGNGetOOXLAgr+z6+CFwSNnkVnJ5jT5rE8CSxsqe6rBjGZnj36xE1ZCq6QKSp
nz6jSYyWWNqxeAz0/UjP69uxcEC0JzHC7nb7doM6LQzxKs5+8tyGY89azcNWmjbk+Rk5Z6elYZuN
cD1QD27mZrad1Bix6ozLhgzpH1iV3DULHtobKaz7bVX/jd2gaNUDq5bkY4xMO1EIVC8cF11eZ0Tj
o5vAxTzgmhsWjKB4NJxwIz0r9fcfno386s5H495zyjKWb9v+ulkscfR8SbsfO7hOVPMQE9TCL0JJ
t0o3wuKDTkGG+dXFlWEU27cPVIKBKVs/njzqikZN/rLS7dFCan/9LRwfV+BPjnRxtWCMeksrNT24
FkyAbeUOxh7/CZNhJWFwr9WE4FQtrW32thhtfdWSf0YLxLIH19QfhmaIUE3A9cRFQekSOV/CCHr8
v0sn1DFeO/cloKcu1cGsazHukjEMYJ0ET/2dEnjUdW4BEeAGNgy9ETCswe5BMwI7btRQagR43ZQ3
VM24/evHakUX2adGN23Fj/l+3KYWlxrvu4xUVbS+ylwGV3pcisxDBbxPrPQqiy85+LEBqRH8S8Rz
idpl/hLBDd8hfpfgr27qjIiTYFqBJI8YDtfvPdtNtMf05hzqzY3bk74fBTrrkpMS2e4BM5XeJM/E
akmicTSD6ICAVTuA11i8OHiqPPlZqd8chBSrQngCt5jEDvXWUfTDaAV82s8L0PsmW2w6tn1tcuVJ
RWNAw9gYhrxBr1Mqwb3wXgRahVVSMWLW7nj6vhZZol/54EJDheBkvOSzNhwr7GObSacX3AXtIVQq
vq4QVh5f/62M7nA/T85a4ku1oIobi6LQz7EEFmu9EW+uOH6RBcX1ew6WR+hXiYr2l4gWLA+mUqIF
rDXa/H9B+Q9NZ5De8lM/BqD45JAq6tiIjXWONgMjT8fuR5OWfSBGf6sk5loECGpgWGIx/YnsrZRz
P2n/DUlvWgFar7W02mspX+IyXdQjG0SLN4hqIdzFWq4hA64ysK4ocehFhrxInDrBJceFqvIjYjKH
mY4eklwK/GxFaHLyS2/1IxVifiHn6uItv9Wr/l8QQao5Ifq9+kA4GCAt3bJYQ+00H8sK2I5sHUJp
nM86pbG6pE/w80nufVZsF2hrqAQcbwoGtpqcgiwy+fjYZ/v89CXQyhhP0ieVZlY96vSn5YxIEmz8
nZLR4rHV6cN6BlOVLgYAduz4dNJMkApmbGPSv8PeHdNj8rnHKx12SFyHDJdXCZf18YktdR2OxjgA
77JvlkYjytMeXrogPamp/GPCr7ePHuSZ/OgnGbOMPioBLPsDV+CGf3Nvv9F5CcUEVpvYGG1SRUdp
O8SjBkatLN2RB/Iz9omtRsU5maGnKpOH6oUewmm4RHZLiHPnjhWJqRL9nctnCrteZvyN02Aglrls
zEcnOLqhEBji7QcFWDZ24vxPUMoGKRjSnTy2kAx64kDC9ystWhpizGkqFV/R4tBRW3QiuykgzzZo
QqWmbhzODqWSikERpCXharOvTyvpzSC736Zl4GW4TpG0yXfS03ybwDB7SjxyDyarSpXDeTePZGCS
zSYcDSHhHWs1Qeqhhs3RBBcSXfRsb2d630TgQ9zO32+QW3pxk6qsFjJqSUP/PL/V9KeF/eamETT9
l9HK4AbnychDsVyAh7MUTjW9j4AuHVPv6XTmGPy9d7f+YoFAhPuFEYb8kFgRMinznN7a1gijuiy3
y5iOjjCTS8aNIpqLuo3/JXO60vpwJKEn6uCMFymxQh1y6vi8ewTrBZkFlxfZfcyZw88ityrdXumg
6tzokJTN5MP/YsibnFdq73kcXKz9idpErup8rXEhwXYyLKxhXLWlLjOkt8Qbkrnv+qwDpBsBfhml
NjFfZY7teQg1CkDRB0NmAD0cNZgF+5J1bv2DgqTUproicSyzpAxO9oASaNpzSmldW526F+6GR2zC
wLr7Zw3UTl1RdMgQ0mARiuIfuKcyOhHifattriVt65SZuVEhUzyiziGbdgmwGtq92vZRfG49oUqn
0e9XQ5zbwcFUFpDWvBMk2vYK1tSpX0UusthGUj+NGAPtGGoVA485hvtEn6nX1J5vnFYCLzSZHhbK
WPx+QLpSeMMMYfnlDUnpqGi/Ntidao8YGYzmzxIasI6GoeaEzDaIPxehaAC5Sg5Ra5RnPWh3NAEK
WitTE1gzaRgbT+I6kLj5ODUu1iL/2edol0dljW+cBSBJ4k9R83qI8UXElogmZcInUfo2mP5nlPJO
igBGRnaCRIclnYMuwm462yUrZdRlrJbmmNrzH5H410unL5Fe8OSEkgShZHBu49eXtPoLck32Nfy4
O6ZgKyW8jWZ89B9aq6ezUAKwYrHl1Ucof/2zZtIrKAY6Po7ru0zDcQuyi2vuIkf/T2lhnTblmz6l
MH0VEGwwxNwfErHOk9ZcNq3gTr7W75oJCYzk+YBHS2+Qhx7hSY4ekqUiDeBJvz4FVSwNGBZxPAJ5
81u1tDw8jMzQ1m8uVQuiIaSscnoo2PKwYKybrLefWJ7Wqeyg89pl+wYvrlOEWS3D9MaBGsSU7lHW
KhrRdzhIFSSI+UekwFCgIQaPV6CFgZPUTAnxevqcJyoXN7yr4TbLYabKLAKC4EYNHofIfvFWWaN4
bi1/Y3a7DMrwRv5p9SgePet5QBrMxcu5jg1ozKi4Z2xJMa5tksW+4yenS9GipHes/2OlAjHYmjmF
sjVLeAhcx7MSWGJXOmzZo2vAYetPcMqc4/ibSAxr4T6k4TLR6wAqNwxugqJfyTlGFKoJM2+M0q4N
5A5Cd16jCmPT1BvJ5N6WOgu1G8QvBVx7G1c9CjAyyZ7N4wOnM6Dsx5TrrptS43LjlNqvEuwxDhyM
KtFcD0+MWjdhD/+SAB2DfLbVNQEatvgr8e9Bp7uJ8YNGb95PJVDrPPpnXG9qfKdktJCX4YrAdTpu
BboHc/8xW1B43KJZwxWBxVfxgdDfayfNWUAe9xu6p8dly/rctPS6oW1X46wMkip8vH30unJ+6EqP
+F2+BLVbEeO2cVJrVIU6AWs+7/nwQemOelIEWVhwI5OPVaGOsbEHw3f8Fk/CF9Vs3pAn2TaYPj+H
BSZG3lqA+JBLaPlVV8ww9D0bkw2D9OtoRkppPlHvg4BcYwWvZfW9q7heEGiJM1nEvxTIvMTTzjiV
+VVf6v1zJK4D5jK/TC2dWLfLntoyBJ6gp5PE+FPNqrBn9CqhvwtA0wKSIcHoMo9WJvziwxsAKTcQ
YzD/9pUdXDUd67QYizXhJrNFmUff1g0KTyN8U6tR3cclPzmJmveXgrEp+4a2qO2RGpH+0Iyax482
JUKBWaKE/ai9quQ9mqNH97BUeo900qvAn78Bki4LrkfATTe8erxyyQ9MRhut6elnJBBUzVGe27E0
u9oD7iDJnCKDgOtSkC0j04dWH67r5ggE4piLv083ermrfHvpYGeECM/gw6TBM/lpKGQ09O5GNYz+
g6A493jk7trQSNuudkzjV/HoOiolfDfYYowXx0txE1N415Cv18GMLCE/6T45qMhEigcUkfY/yAEM
QCwW/fwhWBmKyTP1V45tsLLxmXIk6rzXdaGs5JQOB1Sm6+YSp86sRPQzOdjnLwFu7YuX04W6AHir
CxNznb2sHeeNrIuQYcHFpjJ72zQUDgp7Z+xPdxvmTF6fG0fQQ8KZEguEnx3xms5+7bX4fEfN6zyu
SyfBWC0v0vm1OKoORBNX+jcNMzeGo6N3xaiSSBh8CrEQLu1glPx9pkphsxIjNuTpUD2KhPqLyTq9
B3GZl137P3hGEBUUBEPBJlFEfx21fGG/cdMtBoj6QUS0Ia0kAy1bHN4wNHt9s80Ooe6DyVT20whH
Wmv3OnS9kw/dl+wKo0Mb0aoD6C1yHeVP0BWfJtEUi98NqNNjP3d3sDGwgSANStas335dmb9fyoaF
KEuil/UEdKTdyqCGy3zyN42Jc8bsu9eVC5tv1ScgZspeURKfNn3zM47BlA5zuW6jkCjRQbdWoRKg
opLj6lIMcCudOk+5M3u/kY15RKf9uoj9wsiDdGfNfmuEKUhIy2Ra6IN+/VKBHziXt9pGfKcHAkb5
xGEEYdCiQ+LyaJxJH+UUBBL/vtI61fAzMcJu564b4eHNtNn1lgLQcYPmx8iKCxkSIKoHwU3NsrbX
4MMtt9MwyJWhxA4qQIbxJjsmjVmDOyPxeXxCoMEQRCyHVBtWt8Iy5UvI7DcGcB2bYJYB/kuqx1/V
4eB6ZkuOTJkcwaUpo9WSKBkZ4+CxJC2XQ6RJrjLzAooaDPROO8JbJZO1t7WfW01dpmCusPDW9tbe
3KKWqBOXrFmbcN1uM8TnM12ccyPXBoPMQutNvtEN+lQKIT4pWJVP5Xv9uPoDnOekx520KGlb466o
uTWkxn31u8qxMEn7ZQtsNPVCg1n3i/EQ5lvgcJc07ZART2kE5huPlEAbLHd5XBozkBAE6xn2Tlid
HniGRrqKHp48At61YRgv1Cx5dIUQJPrSApWdeRPhxwMqZyVc+jD50eHY0ajpSnm1nddJH65RJf9J
YvFXscBH66shy4FbOkttpywbl2EvaB87G9WV/Cnl37lRPwgjZkZ1PJB6LRKevKZGTCInd6gpJZAS
f7IV+gssKplQqjRqvrdXxJ2m7WktGjc81nx/r/NdJoLixmR+zfNTP9iu2enHAmioDJzV4DhG+DhT
BDpf5mvcm7jxR8hEqxaAT60X206SK2Lxib+Rtzw7jHYRYhEiCZAaXKe0bA67DfKqYado+oDWIRB3
tG95rsVcr4jVXQywJtprNMj+bSISp0+651hXO0th5lCLtri4aUrLebr70VAay7jk/UxcV1wzbWUj
jl16mXU4
`protect end_protected
