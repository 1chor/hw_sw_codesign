-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tMciMZ8IVuYzYJoNboPgXWIwSYVpXQrv3sOZO2eIVFzT0NDd9gC0bB6Hp5sdwRlBxgKvDKxw5RIi
mHYpiIG2ibbzM+ytuPyXwuUHdIkMtSHUEujWQa2Fmi/P6fPaz/B82wmj3u4uj/NV67yER58FoEFO
eqRqt8Gln1e5gapHTLcruD5wSrlW/4GveNSZKaClTwdtl5zTeGCEeVZBgM4OAEeFP/KTgaO8ojWe
YZo8lLM6RCIk/CinnQBfMU2YNg+LY4BQOOcAqEJ9Zdnh3h726Y/GLrAXzW54pr0Fvw2TEF1j7C3h
LJRq5OMKKiVI9Y90hET5Qkz6d9C6hKQgBrV8LQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11632)
`protect data_block
ZXIid5hdXa+o3CJE3rDMhMy5Iht0zEdPN11kMKr6TszpCBjU9v627xx0TdnMyIsZgVceA6v2JNoL
qtcEXUbqvswHM/5QJcOnn5WxsjF7a2ZlKkRMln0kuWGFHi3jlGGFuV1Ji++ZmILP/ucSnl6YaU9M
suDfueQPY9FcMMAWzZ2zbOFoB3AjyT3rqTEsxtJB/F5Ogmh17fweymwe1Cea5ko+wNLSSdDNyFAh
nkmCJ2+g/SYWg/TINXcASdhead/Cp8qjL5iGKBKufn6LEWskpxhYdwQ1ONiQIcf3C9l+EES9zsAs
Er97UeRqCOMyzopa03iy6zGCgElAnvhD19PdNFatDZulk2nZ71xaBskmw1tZpezw7qWvw3AKMkqQ
slJmn74bdlIt5RsyXYe1JEAkppZkT5ckFRBbAYvOBzAmQthojaPtAWbFAkCkxtFKdbQAvukt+x8B
Q/CUyJDddp6JM2qS6rHaGqt71cbmkg7B8WgQFPnPw5LwWFwn45uPwsx7DUl6hQmbYZ8jcgbq3rcA
l1dK+EQjk2hZItoXNlXy4U221Jpy6pT2Xavh3duZtsuXAXSh1q2T7ovTx2Cq51kOfA+l2njEUoJX
xcDag/Yl5Jn6cHfJCWLpAlJu6eFjQPoeDXzbUhT+fVHUg7cD4AU46dz7oZAB5dnxvWla+j24Z9xo
FcoX1amIifGXNraHft/EP5xGDmAJrDEVNZZIPFdKyquCpPvWKAv0vu/Y1e4FZacLg3y89ULHnB8+
Bi6OmCBOOi/4taRuKFWyfrOd8ie5N2ZRUXKSxvk/L8e1N+w4EuPnrrjOK8FjGYEqlCIQgSejOzNt
ber3+aOORvSePquBPKnElH7pumSy/a5uzqoFJt0zeJJ6Jo2zFjPK8S94F3x3qZ2cU3saf21CGhPY
ppo2CVdW5Aukwsy5k4CCulZbUpOn7yCzrjuNxSvWAnjoaq0lRAyVcsTQHDM/aL9ELIa+8Rfrv9l8
aBGnTgoFc+RB5Q4imC+Dk7W8GydLtp0H0eyZHXkhS+mXDgczH04paZ3Jbrfp3pZPPe1aUzKOqsvr
U3c+OvPIt4Sul7lQSZMpqvfTu+usYVY43IFFJHom9k7Vkg4lKPKFt9XhggiztNmNHhJM7m3LkvUy
38BQv239qzIftoqu7qg4UQz/HN4uxBbziFKdtcMAXdUkKJmwNssTrAHB9ZalHRLK4qs5G+2TYtLW
QwU2tnB1fmaFSHDjM8mCWTVlJhEY4F6Py/zktsE5Mlt66D+yX7uxwXUrFcHfM/pZlW8OuKLkAsVj
/GLZIuXXKEigSGIg76VkOuHtai3oDZItnfH8ABKqeHXO7wIfCJOhG4vm4UODJmzspvnzXpfbdrAm
9GCYUsI15KdwZt55QhE7xF3mtIab4RhtUj6BdaK7PL0qJ+oj38GM+JZVj2olGCTzoEqMl2zfcBbf
RGbSdXCo4MyM3EgfpS9CwwiA+3DXhKqmzc7jGXGqxBcKe++0fCFa1rP/Oy81Kd957fyIxxMGIfo8
8hSURWgMisd5GgyEttHIUOSnf3h2IwmphRLPUX1UeGF+254FsrJQEwWQw+3vheZ9TkSHaw/LCZCz
3GR8ewik9vd3uJNf0VnqvQ4AXG7sTYJlhD8/aIyxNCoz6g0o1TLxVzuOBO45kh3AYcr7WZIc3fB6
X6Fo8Rou6h45P4mTpL7dFwm/InJZ/cRJxFqmFOglYgBUXh4Rffqek8C1hyui9w/wHsXksgvKF/42
uOZs/HmOLnAtbrMq/NaCkY23y6LXivbze74kWg8JXClSex33CsVwTssm73eqMCd95XADV6ZaTjlh
Imgk7jNSGCP9Cmx22GS89ObVuShb11+asB+EXVOMaeqcexdIfwK0bJbBlWTWX4BPDSEiWoEtVQnB
ZXraDndujEleSnD5kq+3rkAhbFs7COpqWTJMrSeHSgL40eYjGYNIdJSgHVXcHAGzYlNxb+rW0ORK
Ek0i1DtF5vL1VZvcat+jfGxgKn26iMWurcI/zfUWtd/xyDKlPhJgU6jlLsmxcUF0x78frv6GRg0T
fIG9BtiYO4aSc0QZUqf9xOmHPnCz/iL1wxK4gI5BMW8WlnRQGUD+gzEUljjA4Xm9wwPbhIKN+rGQ
zlj0yzUFqS/CD93IziYZ8TqeUtD5ctRthEit+TetZQ3Dcea01CH0qpGw1RkM1OSxCCaE7HQTfsrd
gp7uavA/MGeTYetbttRSOHtUqtBQbwxu5e7yCLFse4dIcvhVdTjJ3TfFl2b2ZJVBKoLofbX2h83x
eeTXDAUI0XLdFo71Bagj3dsyKZN1o9R2meMf8IKK+ImimjobGK8Cb44uSGuRvF5nDxWDT6rtj0PS
1Zv6wzuLGVIOJ9BWGxHGmd7lDCwLdILBWcMlnxFcdSRSQKHxNOUnh5Udsg9PZ66rZn3t/2lpUfSH
JE+w1foKqF3xpV6TqnV1RtzsPP+nmoQVbrM+c4gLdwZqERrEN/PnOYT4Qo+OkHOaPqyztSjN6cAR
cHy/IeEW6oJz0+C58VOumrVRyrHzsA2F7Bmv35LEIF80Apy6wqeogISanLSiuEgDLRJa1ViNgE9q
fn1uXZC0OuneGIlw0sxH5Ske7zAb9vPNWH8ZSZPQcyPon2JD7VGElPFaGj9Oj1u3gCCtBGYGCLjx
dnFpmFAkkEh1TmBPHkepxSxjwZesZzgUOb/5iHaePy+5sR7taqZgFskZj0BYWCEvgZexGDDyfZuQ
sxmCnHl4jIOvp+Z+voN0657OgHV82aBslafkuWnwZa54p2ZWiAK9Te3wGJ9eoKdDFfCDZ8rkxp0t
b7IXG/1sNmL0qrqzAegGKIsgA3QdWonEhBcbYuwza5WXAhDWNthrdG98G7AIKhXg9aXNXOzt2el2
rJzCno2QWx6EHqu2HOS/9Hbz0egcJ/7vB50U4IOrPh9kOHSvzvRMSxLJwM6mExxaVUFh+Gnncwom
xXfpCiI1D6eBQEphQ8ouHwJFTIMVKIgZCvcYEdAD9b2hgbIC2jILiV/4aquBzeFvpONpPKMxk++L
J0ESLSKZBKbfAcwX/XN3mepvvv9fdMHVyMzCy8tD9QbntIX1ET+twR/bNdDkXRDC9mWle9sgslZa
IGL+GTVc8rmDJZ1cvi3tx55EC4JGNo7Nn2ZHfDRteXqoxb/9mCwWr4zJCM1YqBHNeiZ7mT/fXfD2
B7Md3GDxSANPhathP0D6oI0nWw3GOyLAxBoyRhEZb/hXPoRVHz36Dtgmx9dMWKM0PeqvnMEMfsOM
CjRmOiwxEnOulAqF0/5BMS2VwGzm3U2ZGbctBTqdCqMwFoWDCvB8I3VVmj/aSHYq6m/7nBiqg7d8
CNgpoxinSAhZYFI2cuuGmSIv3aRs9gssOGX1CgvzRz4WPqjhAr2+xVW1E9TUQHpmfgv+MrACDoAi
zjlkH8K3pAXZQapCln6I7NE8bU0hLsZQC5sE+qD/rOtGWzFhH1KV2UOP445aZ7qwu1gQos4pJTVq
jLq+vUiSoTKcMzmew60hT0lkNpVIw6v+935QKE5M5Dd64UoP0DAgb7ma6N3HB9f5DVy9az9NkDGb
Km2f5Z11yFt7O+3mabCeCc44OyflGnmaSqMmLntFGpfplfU6oboau33oT/QQjz/edpMPanhqr9J8
XVbLNq3SZxV8jqAI5xVZR0/912IwjAztLqlLJy5bSb1q1Ogv62twJgmAhifmvu64c/9g7jE15qNZ
iRPsvQOl5OsQ6P+HEzRiVgJSg94LByAI7b8aAUSS2pxZbgMapXvjMEa+5nSUma/PyhNgyrQg1qfM
YBbj5JiuNsepm5/EkUIjoh1fYO6N1fYOtaPJi0yMmsVBDqRni/QvGEH0XxqFqlx+82F2mE+cmmcw
zbJoqbu5Q1t+v3Mfe4EiS3QwxGCMVKYEKsfOc2OPKHQm39nLu0TVSMYebO+p9Bi8Vti+exaawO98
m0zGj5s4gEmDiaGlAxIysInlayCo+ipEmwOqQ/d0/ogxue9YGpau0cIiTsqLTzUBp09amlB+L8vK
LjEQWwtaaifNeGq8qCG4tI6B5/NX9toSg/I2V9r5CkJSPc5lVKQUAZJJ8+nd5HuDDODWTyvLhVak
aejkQjS6MxIriAi1mLlJ9kMdSuG3lXbjeX4ueEr4o30ctvhcq+PKNjNSrn1U80E56cHwCKQb9ne9
EqZVwWMxgCWVjLhMqCKVVOjlqT1IN6c1Wei32TUcLd3odVwgjD+vYrWy+5QkV/6bFkgq1G9VCWmX
6apD7v4N2b/OZDoiiCvfbArM5VSr1tYfHwrqN2zV+Tt+5uXLFq5WQB3VFc8YagKjDN8WCLhzzPn1
DUJs6e396E0VExESqhVU1/RpUYZ08ugjXHyT3VD8hEcXQyxo3Sd4Ay6DeAUI5hO3yY+j2cYmcHtQ
UGFkVeXzoRgzePi5otGjvao9z2wHhMhzcL7Wq0FYsi7z3yLph26PaIUItNxBJOSURLrnOsPDb5ju
lO1FIIWdOVfovt7ZF2tSXHdKWjv28vgMadXjc1fUM0paw5EqQN35+BZG/PIWH/vc9fLXgiMJrH2l
BsyvQN4Bg0+dXv6Wkj12IFZr2vUrZ79DFeOOsUSRxLs24zJ3g+jiotDoTh1HkPjkpWBySxAp3YGK
PVAz3DVcts4fqDqNgEaFFrbt040bNAJMKcOzvpWPPWJSU+jDMvBXzQ4/ffH4bKItY9LjZtmG5oJV
cm2/L/UbIJL0Q79r3Pfxz0R2DQJcg1XYbCODZDM7RXclNcv5ELlqnrfJNdMQqyvUqDsqy9hkFEj4
fx7SOwEvnO/qbqcjs5f8mFjGaOCTWnzoncOJg8Ch5TV8XkhMb0JHsEuVawfxjxqTk2ZkfVJH09EM
NbtXl/fk5sMfdcydKIUv1onnDwMdI9cmqXpPB5M7Up+zmS30j1W2zwSII9cgSLDWI6W3P5A5bGIi
92mncRJ+hMBLN09t+CgkqVb05ioEQPUyMpveCkw62N5X4cP2O35KX7q6iz5iVq9whS9w3e7SoNSS
ADe5V6Q9kV4JHbLFEkRXQw5njO/ERn2wGv2FYCRI8miyRdSVAMYN4hJ0Ahh5FycmMwnW6Xu/ipLY
ZwWMQl0I9B5CagzkJ4LZY4f85dH/pjRc5alEreZUqXX0+W0q51cm01Mk+o1ASkO8Qbi1rFkB6Jxj
aoUxe8qCqCpYLb5u4ixzdx0yzcR/YDULP687XUE0WGamr9RmY964Cm6wlT7f+lc3gRT2HDZIroa1
dmriEOVEvJNKS35QzUz0SHMxgf2ICXHEc5gKSUlRAQHvdgcXutYDO/Bu9VtutOI7Bb/FWBnjNpIJ
NBTWraBY/XpYQIT/OWwmy7Y7/UyMSZ8c+EDBeeb6YJ/hHnPdakzYllTISl9Mt4NALw98gVHXvJXF
r9mO9zVp/33PKJ9O72kTvcXlGVbrtmqOXnRrbkWTNp8bEc5xlNI3uWgTCVPoKC0kXflHelaz6cYI
ZcxvfY82yYyPY9xdUAvDnoOyfF7RjGUwOFT2dAydT51MhBopuIulu3jvucfwuoaNF6wC/zN5U1Rk
alVtMrXQ9qbZeGNtQlSsakA2WaDAE7nVngUdN4idwTOncKqhKqv5gHNg3lDh2xNEX4oxMt+654V5
Dy3Nu55V2IZgeWWMKzZ4rfZAuS3OW+wB3XElJeC3SCuUBHn3IAKZ1fcQuibDBGQvIfYfB65Zgo49
zY7ComyNUZezZsvVXlh4WDFwoHrhP7Qs0CGs7m9NI8uERiVwm/yYGj+5OMx851yUGs+eYzAtiEiP
hOnmBvb28RbazALfHejVjg04CJPVKP+HiP7qTj2E7C+qp1rllq+XbIN1yJpXRJDk9ECyMnTUUdKU
ksE7ASru9idE9obykahIfkS5saoywldp+wY8w4C7B7bvETm+Ar4Gajbk2+gdwxuDjaYX1ofmfoVp
FvaZM5foz3XKCWLQKUQtsjesbHncodz7yAX2HRbFBRzLd/ytrWRucCD6qrmCJDymPcIZalUTV1Zs
KKjOqRp0Hp7zonhECbU/QUnoJlLbnZ7LLmTy7Kp27dtM5nG9FpUyZhWGMjlgxl4AYhIUjBNhg2Iw
GYJDuwkjWqD+2sGeiV1isd8r6WeLDR8QANG4NHSCJZo97tyqM4OsJII+nl6ChUaW0urP4gs09hyQ
IgR+Och4s5G61ioZxqqRT86SmC6hRRP4nRIO6ez8X4WDOMaiUAjF7/CPjlhhRGRj5Ifml8/MiqEu
nModBs16Z6vfxtviUggk0pw8IBdl0FkDUMXsiAUEeJZ3Dq72URCbRezfYt3qu07VjofKllyNAC5s
gybd98oAUK79VotrNlZD4Wzv8PFj+lel1Tn7AEQKmIMA1dfmwreVQ/mQIQ7ObRfFiZcrFtmMbVI+
1ZFOHdgZ0SJnQwNTYoutZSkzn/qR6xQS9xsz91CGO2Q5aVKOvQ4TemhYH7uX0MJjwutbJ2TLYgOa
RJkNwl+TbCFLvEtZixIYk501I0lVxnlBoPiR/DsJ6AZljb74Xexf1Zfhj+z7e6jQvOVwRgTso7nx
OGHkW4ZfuYwpruSmYbtlz9NxUbrTzzrxiXCS+oLIeL+W/EkFEK+7bYU+EXasBf64XhtD1ed2KxSI
ohDmEI6e2qZ8fCvs4EeNK2a+v9kf+oMfi7tVjbxQxZ7dpZSXEBkHElgIEatVkUNtmkqRqiwTbXGu
78/Cl4+XiJ+B2+GzYHpYZ9lFi1DrnHoQBd4X7KgYUof3MKK7jjjOnZbsszAGI8/LPs1e5TkBzJn/
AZ1fJOi5JUuVN/G4a34jdLBChnPwdVflcofvqrS2aUuFN4v1GqfiCQl1cBKV/+A0QUZIPPtTV3uL
87YciF4huHKrX4LZGIVMbKZHoVHEFf+mmoSHh88rXgaZy5aK68rBAUtHKE29hNGOLYV7TUZ/DAdI
gmwqRaU/yPSXT15uS852kxzwuL01SKqanvqbrcgqaq5DDh5JqnZQ84hLfS/LgCySUsBRRRPo0ICp
OVi1uXnzlW+OVaB9C97zzKCTZXVcqRP2Mrfd/LQdFo6kPIJe0/iDn07YcHuGsNtyahFYHB4FFWKL
VnlsfA7kihCp/2oJNPdJkJ2le0Mt1o4iEDLIdQDVPzJC8Zl5A0dWMvjUH3Tky3x+yYfQOosP5Jfx
CkFkw/MWKXCEQdtVAa40aTz9hzu79+pnRgnaq0MJvplM4eRNmCEpjEfsIijYyg70oOQtpMdYIKek
60gPNTGBueQ1NGBR/g0EBWwi3j2QmSqgAr+a3+c9uXSP/q2IVLSRaWJdMo8Z93OCKSL7Q3erLadd
4TCvsTq9ERCDkvliW0nDLhzlj/cqqXhRCKHAeXVI0g61zv2vJv9kAGZ+PoSadO4OsWaoJ/R8SqT7
hf5TyRIpm8WE0G/IDaXTie7IdUhlrmjZgtEE/DB9jODRAdsBIU0cdzQinMmsWCUaNg+pewGgNhtP
kmOH1QOesPiEpeMOfxYPLFil5Dct+NWheyPq0h+MviTj7hNVJkllSkorQc0i/pA+94MKl5d48zi+
/Ag0YXed6dJ3F1oQLoqm+h3ujLGYVYpo/YySFb1/Je5kQeaktqt+U68fblEvezT9l/MSsvHoStut
Zt7zHPJbigN597W53poY7FmzQAEEnEMlhpgwk/8H/s0hdBtBEKxoytPHqhzKsJOtK0odwPwjXsvI
Asmc7x5aPwqwJe7wabpft2/mpUEDGmuzY2sifVCLbNmHpA3I9lVpZuypKfbr0rTiBN+jIhYXDDd5
hLCpt8wi9/2Kb9Hp98/TsudTJBTUkETdOiw/FcXpiu4t9fv4VR/loamArvX+ORUao5vx8M9LS5dU
2oTK4z+bz9rVlfjWV7+kg1lB9yO1A5DPW9p5eHXnWl6u68csEniqH/YMpLiBh4Ws3kdCexAzR5Ms
Nd+HeKVHy/Kdt+KI9TFZT3OwYlc4v4IjgKlM4NGZdiUSXJUGzWH5jXpUDEq3h+JUWnN/bREEyA8P
FLXIWh4TBWQfnLRcrwtAV0vKnDS3ot5PlfD9Yg5y/ptqLxgPp1q4rYx5H5r/ZQQDbjEyGu1q0zDe
AXZaOreLhAZQmkuwNEVFg8DJE2Lr93u8GRiV+SAzDTNX+kccTr8ZTzo6PMphWc1atPwhcTMQqr6z
7exkgCw+SDjRBEa8Y5oel/0yr/+j013zwNGYWhARZKgqlgtlFB6S9geKUl9T+IDl8ofBiofKLGFn
VswZAe/U+iu+0NyPN8MseXwB5CusZ3VVX8I8PPtT8qWT1B6h1KIY1a4y+hoV0Z5g3dbzu103i3W/
8ZrEiegCLtneltxWkgRZsW2XEiS0mK9zbHLqsmFSMwupvZktB402ozGIOymbyQdgk/8hFYRA3miG
W5FJQsPxS/Qx7+zLJl+kKpYdrlS/poSToiYlbODt3YTCGLP4buPKlN+gelaSLlOzyed6cREz8H0X
uywVD81Q+Wg1lpf0v98vCahvE7nqAyD486zFr4hmBEmrjDUgJBoYtLwDo7TuqA+vFsMToMbWIrX7
2T3/56aFiJvtU6EKtZ9DMxPY88fVMSAeNDldBYVvZ7uhDk9IoQE2wWjiCmaodK7piti9fWA5O+zG
ryJv3uf5sSXJZGrYvplML21A/rtHFOEphgKzPGa8mC2S1t+ud9lPxfAQQ+6mWrl71mQ8cmcfqwdQ
ZeUEnvlFVCSioY0RroAi61L/Ndc6ZIMVhr+uJHvHUC50ssNlySptx+/XEVDvL3DCC4P0Hksw0LJn
7QyMMvk+nRPKKqIr43CjnYf42FP7MQiNWplZt/++JD/2PcPJBb7ixleDBf1t73tm9ZL9ayFB7zZC
+yxmJ9p080fo/4CbRJw7dShG7ACphby8cOKhbHHN9mwRX3vhCDq28dSq4h8qV8PiYvKEbU+oUypb
o+bssc0p7lLERh/O2Y7njQ+R1c7Q3dCFDP9LZyFnosPKJSKTxLn3+qPtkB7gQf/bGCgfCUc7BuB9
7ucRd4x251wxZs7VwrCWRrWC8CeiQeXUYbnasTLsoEWBeRzI1UWnDDWQMzz/hZC2jsWBWfQjbSK5
xS3j02jufzdE3NA7YYUuuwFWyLIHV0QF1GC8HM/FkyuVn+y17m1FTxH4qbTQqmTIcG0D4noGJDg3
WEm++uB/PgQvYgjt5im3cmM5OOpcZX3tsZPFHdOf5VEg+ZLSKdBqcW39NA6D6mGdJS82UrU4lbi2
BB2ZdHw0CpedbkDj6l7ldXyMOcM7ShYotz+YVA5ZrQWMjhksa+Fcs9EutpZsBWHgn6ymLkhRmCeI
WsnxcryL0VfkQuxL322y0jcsQlei8w2BlscrZmOM/zYZ8J/C/j/WRoBL9GQcEnqjgVqLuohPUiy4
dgGe6OSDDNP3hgaNL/49HdE7+1LF6A3qldebQK1jj0CdYaj+TOOtQjo3PsMpQFX/7ef61ebPctFz
lmmy1hAqSxYYg0YFMgA8bBPyRu+EnVMH3ul8corNtz+Odz4+HDfTrE1U0m4o+x+22a0jvptsBrnJ
7LW11gkLJjdlEEyfFzHF+Chk53RGfdC7ycNBkYuh5Uq3OILhTH2i5v8p+wJi/3Oy55VHPsz4xG86
jbRe/QyMdMxxAHDRvC/yyna0aRpkwprb2y6VVKbz4n2xTFKZdHc9577NnMZfYc0qxyMf/o2+egpk
yVH1gwXymHEj2zQtE+x0mX/Lpro6aV/82QluTyQfMD7OGQF/Z9IqM0HvwROWDZochfBupe73wxY7
eJZ2G7A7SaPTqpdFB6d//iEFYZ8O1hUzChMwBAafqkenqLy/qxDRVl9FjCCu+6hSbUXCZbZ5uN0i
YKLJCKkGVHNYwrKVNd6PwWdgQ0b9lDx+Ppu9nKPSem7p8nobkUA0enjy/76jnpdu/XrCrcqM6RGi
0ybf5Hsx2eywH0stqDVXXGPmiXIOfEsI+1dCqgwt62L14fWUK96rXlg5+PFKyASm9gmGgX5iYuik
QLNgbDpk8ot4YcteEYDO7A38evpz1w4ovBhFAa1ZfFtYQtVU7VJNNq/HJHENmwTpnnXRQGexxait
rSTpXypw/3GuF0VK/h2sCAggvxuR8o2v3Hux3WQqq+VXS2Gh91ArjUao5urL0MXbY3gIo3RPQrTo
Ke9GT4v8rTAF2LqzgFTjjuwvrI7SnCs92OuZLXjdylN7vNd0GzOAQq/xhWGM6ACQkpYk7I3s6qlT
3NraFGAhkQnACelUbLHWSqUzzEqjXXBC7Wg/y2k7v9uzVo9MC/jSHuapi+9JCALU9Ed5RLsVQiYL
SgrdS+lQGaCaWYGYGuTGnoEsrXuwnX7nP5bsp8LlZP1dz2sy8Hlka3Bu6rjQBSZIGp5QVt8KeJVW
dKMmGJPtsNHJ9q80VYzLmBgtF71L6HQBXeQqPrQoqnskeG+fBUvAGFX+VjPqwgAjhE1LOAk7fR7N
OMCRdCfDAm/EYBYmEYtR3/sPHnag3iXSqCyVA9Nayqd/U2XcbBwA9u+nXejK0iYwGoqE9BeWf8gA
BNVs3ofHFk3XHbs5F22KWiDgYXuUaRF8iffZLP5o6eoSuoic4fPrCVaiMWOC0miF5/RUlvAH2CIK
5USeOx2fQDX+LgHgt7TeflBFDeOut93pM0VG8CTo0mEaG4oJRluOwxE9TYjfW45a0Smh7XMqcTpO
YatJqSblV1tpbNLYnEIGLT3nOfC5DEdoPE10FiVh+KHS6PWuN8lvebBQMKu+2FbIYlRYMTtZ4iWQ
tFPBg34vvjKnW84xY6d0/8c0k5h0BMw9PzE3E4KB507iwlbexbbBYIH0NfsbqJjFFfkjDS4sAdzu
T/XmH0x20u1n9CvGAHz49fndpvkdzZkkM5HVca3abuanNXiHQ8fTl9/lXgJi3AfxBfSpEsRzkmlJ
DW1VBM4Mx/RmCIoWTGP23R/Hz8OhRlAASsnoUP5dlPhCE1WaNfHBK6dOjFqDfkX3wkzG3d5uz71y
R90nsKoXOI8wZWdRBSG7Sx5ViXVkLwRGb0OhoSCwGnOZ9YT5KFwPkhjUS3gF3o0GDbfqhGAuMBHq
Bg2qE0FeAIkX8aVO45R7orOOVcX42EAAhd2whPrSAA2R24O/BWCEMFk6CEMT8aI1Z30Awkkg4hIZ
2kvAznmkaG+EAsvP7OKt9AzJK2PSn2XtMrGHwz9dQglw5H9hfJ10dBD2h6KwoRs4khf/UxDOVL5T
ErxJXyKr6OR4LYvLL6GdvLloFwAz1R9ERb8GVYbGPhtZqoEttfhJggYDv2SaNZW1em7g0/qHOCDw
MyjgXdmWf9bYXk1t5BcF3+DlS2vGD5P5mfBBABulSajMqy69mst0OalqnHOAKZsiNwWuLUWcniZ1
jrYS2SbtCizp4tNlV8xH2TZ/ii5WbmZwhFM2rpLG6HLBuojMNH+JP8HdJqgsC2XAxahTzN2l4Zpd
SflgUovvTJpQEvPlhVPZMocpwTY4CUxQw4rlwZ/5RDmuSfQNf9pMNVUxC6rWQ3Rp27by5i2G19yB
SKS49fOJI8v5Zvs69uEFdheOSeZ3K/zJqNxGNeP/v+4VR4GRGKeqOC/jD8L1xs18ECqFf7qinka3
S9KjEvPJq1szZeD0Y8o8Oj2LTVrjhfgdJCN56Qs3kqHLiuXqMGKH6zZGQPnfhsVvdnEqjdDPIJlY
fQ89pCSsHAES0aJqqsFcXu6zJwEwv53oZvqgaW7vBCB9RAqLcS+t5dM/9o1zI0Nn20Njt9loTLgM
hgyyZaNsFL7n1Og70Uj/9odmZzy0rGOqGMZvFbuPpwgTKE1G4VP1GWSZS/HBNenP0fN69/6d3uUO
TMQA1sjAQqTFOs/BXAm/bP3Az/W6YIkllBhpj/Z9pn5t/I0pMbvccI70Vok3A9+NgLCkirvqlKYC
0KREE0t3j03Gw80pDnUn7jfb2dbq3fnUWiWs4xeDdrYlDMN1tin5c3HJRnQkYF16Vregh/p9B2qX
9cYgW+p3736QIvVWx9jJiQICDoMu7J/Xt3X3a7JN3ASq5mFxSItyLN+vdiKRxgdGmID/bIoW84uQ
vFjVYWjLVchJZ6BvxskEDJTi1DeSN/4EtVSA6aqaTXnsPBfWkKlv0sDRZZaWGTObVyx0+3lkLcYg
R6Xv/sw6gdasmwRKh77ipJnbWszaVpi/G6wNTUMhHRUVisgOtR/AanDCgbABUDtzKHnj6cPa/vFe
h2lLQx5HIurTGQEh/nD0mDYgZH2xnOKeraG6bMEFXYbn/XSMBAXE58gv80d5vzrzmsCWMjRlSt/6
FlJ5gNjD9N5Co3dC//0vWrstQymnEDE5gg22W+iWUDuvJcplYbNEuaezSKjd11BHcKoC4O/z/iyo
RFYny3OTiUUqlMTMjhylTR7tgtmoPIyQy+VMot5m1mgzQhIz3bfCLdRgB72jyHVzdt9bPgZS9amV
TpHHD/Ut6/rN7p4HeNyURgKiydWmV/c8vtmwRiU9su7DUC5qc7gLS2dcmXszKnjytcRfom13r8g3
KdQOGiSwUGPOZjOAhFPDqDIs9egfL8lzQtSTp33WHhentxVeo12hX70oXG09G0rs8LzzfAKlIr32
kRAW72PMvgLhtmIGYB2ZQ8SkFfzqxWafBrxuphy+Y1GoeG5F/jWDF92N8sG3WxMubPt52J4wtDkn
nTHOZpGF+OKufHvLwSpyO0QCciwV+D+xBdCxZCsqoq7EEzVwRF1FWN3TO/SQvHQLzi0ApvsM595+
VJiWU1b6GwKpFZMzr49ejTZE/XlNu6laiGVKiyKXgaN4RZhBEUrezA/mlZBHIeTeGqhhAlPoDrUv
SxBKMfYsIPa+qQn2RBhGEDdGWoNxrzat61rj1I4kdnk89XkvfoffHNTGqul+0h/B5hVoLLERDDx+
lQJ59IViYxCSbDKypplHj4ChXBu/VHHVttDhRonaLsu5XejPtkJIPlnTQNZrm/GCHKQkLqtVCTza
Cdn/eaxZLAfFPV+McCEuG78DyibXIRxuNGqKv2boFnfSVpFfr6rLWZ99TmHs8kbl9O4utR5QtQpF
tCBkCopbVcMQx7S6Xj8besCw4bY2s36WRXeMLszFCkXbbqaoxe6wrWhVEjXqiO6NlPl2+TRr6SjM
DlHr5rKJDShWrvgJG+aPCureCGd8cWombsuedosP8RBcldLMypst6KcnEMZYuqSNMvwXydH3cq4B
uaNZvxnnqSVmjAxJzXjZ7sywwivORoCMHIeHsx9NG+C6NoE2f5RYH+E9ixmo4A92L717cPd8Cv32
NIWgiESshoxzFAdZJTphlp6p+OnV/b3EYhdYiuyWT9XrgxqQS2H/QXzywl1KRU4/0YEfFZ7udHcM
aQ6lVS523uEn5ljeqXlRAzh07zZ9RAsBHZk/AaYylj8U8LM1iyoNnnPQGlerzDRQAQFl6XV/50tQ
40YiV4mmX1VUH1XW6aUbKVtDh0gcAvrq1ahbDFYgIVDIVss+f1tWmQomQL6T7CxIhXHOR+isZF3J
VmYYK8ByGmN2Vq9Z2/ta8cCn/haZ+YyJjDvz1TzN9JqgGfLZA17PPl310QXmj7GzYgvUzzz4eBgZ
4ttI7vCgqXXF8ZsEiBKt7oSupLH6U/3yskPx7s/bWqyfIEKRhJK5tzlkbf3P7eCzRayR0cSu942x
IjRRn+khJtVPZIIrKKegF3+dyPxC7sLOJdtJgTnIPFhI7ddxpfn2f+oAVw+ETcn38oXVO6u4gFlN
q35H/H2dyURbZa1wUmVxkEiNr0j679jSR+mnl6w347L4t+a5HATPJf4RJQYciUpfwhP20h8AAJ+k
TWIvJnHzPy/NPlbXKE5Vv1qVV9xCW0YzBWt+ExnYWQMSPclyMI40ticSCXk6RngWWp5k9qQR1PVI
9F+d7JwFc5PN2L9gmaakbteHRETQ3oLo6k7CbfulrVXPBXxLupp3VkQ/y0KjE+C3foWQZLHGTAsM
7cW118uqdug9vZNQg7QYT3P2wvupUAlG3U7RQrFl3KtS0hJZ+bqHgsXddRJky+g8qz0eLlvtEdJC
8StogcyvSIVgKiJr+Ee7rKBIszTaM3SPWoh6xdbdCcKDDT3+Gs42muicJ40yxKfhQ8UacBLMIJB2
4MXRGQwuqmDMbpk7YhFS9hkiEzo6BR3KZmg7e5VE9UAfhRbii0S5yskoFnu2zZLhzNm5R/tTgcdI
zZv+mVxmDxgyOIvrDa1RiCe5uinAwkstV2evd15uh5mX0uuG5LxTousqcX3jAjlU5H3B6sctlgBv
7jPgWii9hcGHWiR3kVj6iJnSFoYFWRFxTM/akvdc4hidlBDVfBoVUuLcGiYFVXWvSjVipZ45orNa
x1fWKveRtFvA6FBu9B36MuTgoWUMDePz3inLljK+AqgJNp/VvBiSwXMN0/o9PJQ0UVGvqbo0lN9K
OjYhUb5X4jSV8XHhstuvN+OTq+FVXmSTpyoOga03JjrI8I00iNRKnKzhXHdwnXTdu3UEIdfy0VX6
CFw8Nmq7QzhKwl+8Bu/Z+4XfdAriSWQ0ZX0h4jj0hOWTmNJZv+eAqDUyWXho9+YUDcVnYQFpkZ0j
SZJZstWrkj8D9X5G5AkymUKEe7uHplkAEnauKWyHK7gAs+CDZVR3GmtY6mBrsuBeZtJ1kiy0oQat
/taHdl4L39IT6C5dkpRvVoPr8esXHNqTEOK4O4wWsfPpRBvCs6LmeayRtBDZZSfPgRtaNVCUa2Qy
/rgHFQuWqQpd6dpni2qXjnWBxlwT41HBwLpD4FwADKr5xEcogMRXh4BfmoCLmkC+vQGpUlPlBUoS
kqwijBEXZqqvLJc/QVrveQOfVHaGSRuyIJjTUOYBHM7VH/VD/bFd5vkWeBR+0ZGlzkMy79KAkajN
L1iVa9sCoHFqWuRHlozHgeW6wWHLJi2x7siG17SRGTvJ/xm+qSz7XnJHcSqimyOY4DZA3fZyHvSD
f+VufrM+JMu5LSjKlbucxfLMgwHp3cpQ8sdJ8PYZGTY0175W8EP9BPoI+VvPdVWhgaiyWNefBYPE
O94qWRWmb/qEyll+uHs19wMrrK3YUSwpxjz3tBAXvzdQp+Osq6aEGjHcn14gRNB+AfCidSLlc8Kq
JLzJ7gt5WAHqbnxaW0sZNHl/IyRSkVrtE7jkn+BsxLpdqV2fFSB+BHtfW/KadLnRDJsdlOfY0BJw
DEp1w75OHiWCsEb30mAgJVvQ8+3htEKIIIC4Gan+U/5YKlBnzUAL1/LqLJvYWxOQ+oi2tSkzmxfa
1U5XqYVlxkuUTMqaGitzKsIYG48cUTWVB9UZiumOA9EdMFFq64UXaVdSWhZDvy4lyQ/7uZ3nA34N
m7bMb75tVvD1kx2TSN6BNNrX2tm9sBWXS4mT7Fh1fegsyRYMczZ83NWJcv7PefjzKVHRaOZPg1FJ
YZ7Ge8wjYFNrfl+CYTDwtHjbo0BQ26RLVB6pj76JyV6cQwtUtwzM6iN22cPIJK1PUeshmaJf4ujr
vNWiqW7nvpEsof86gsGM6u3T0jmXFIySlXHNJX2F7D3ToFFwqaVsu7+QNBc2n6F2lTu4FyEfUUK6
hEz7nA==
`protect end_protected
