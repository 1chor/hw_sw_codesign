-- reverb_template.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity reverb_template is
	port (
		audio_ADCDAT                 : in    std_logic                     := '0';             --           audio.ADCDAT
		audio_ADCLRCK                : in    std_logic                     := '0';             --                .ADCLRCK
		audio_BCLK                   : in    std_logic                     := '0';             --                .BCLK
		audio_DACDAT                 : out   std_logic;                                        --                .DACDAT
		audio_DACLRCK                : in    std_logic                     := '0';             --                .DACLRCK
		audio_clk_clk                : out   std_logic;                                        --       audio_clk.clk
		audio_config_SDAT            : inout std_logic                     := '0';             --    audio_config.SDAT
		audio_config_SCLK            : out   std_logic;                                        --                .SCLK
		clk_clk                      : in    std_logic                     := '0';             --             clk.clk
		clk_125_clk                  : out   std_logic;                                        --         clk_125.clk
		clk_25_clk                   : out   std_logic;                                        --          clk_25.clk
		clk_2p5_clk                  : out   std_logic;                                        --         clk_2p5.clk
		reset_reset_n                : in    std_logic                     := '0';             --           reset.reset_n
		sdcard_b_SD_cmd              : inout std_logic                     := '0';             --          sdcard.b_SD_cmd
		sdcard_b_SD_dat              : inout std_logic                     := '0';             --                .b_SD_dat
		sdcard_b_SD_dat3             : inout std_logic                     := '0';             --                .b_SD_dat3
		sdcard_o_SD_clock            : out   std_logic;                                        --                .o_SD_clock
		sdram_addr                   : out   std_logic_vector(12 downto 0);                    --           sdram.addr
		sdram_ba                     : out   std_logic_vector(1 downto 0);                     --                .ba
		sdram_cas_n                  : out   std_logic;                                        --                .cas_n
		sdram_cke                    : out   std_logic;                                        --                .cke
		sdram_cs_n                   : out   std_logic;                                        --                .cs_n
		sdram_dq                     : inout std_logic_vector(31 downto 0) := (others => '0'); --                .dq
		sdram_dqm                    : out   std_logic_vector(3 downto 0);                     --                .dqm
		sdram_ras_n                  : out   std_logic;                                        --                .ras_n
		sdram_we_n                   : out   std_logic;                                        --                .we_n
		sdram_clk_clk                : out   std_logic;                                        --       sdram_clk.clk
		sram_DQ                      : inout std_logic_vector(15 downto 0) := (others => '0'); --            sram.DQ
		sram_ADDR                    : out   std_logic_vector(19 downto 0);                    --                .ADDR
		sram_LB_N                    : out   std_logic;                                        --                .LB_N
		sram_UB_N                    : out   std_logic;                                        --                .UB_N
		sram_CE_N                    : out   std_logic;                                        --                .CE_N
		sram_OE_N                    : out   std_logic;                                        --                .OE_N
		sram_WE_N                    : out   std_logic;                                        --                .WE_N
		textmode_b                   : out   std_logic_vector(7 downto 0);                     --        textmode.b
		textmode_den                 : out   std_logic;                                        --                .den
		textmode_g                   : out   std_logic_vector(7 downto 0);                     --                .g
		textmode_hd                  : out   std_logic;                                        --                .hd
		textmode_r                   : out   std_logic_vector(7 downto 0);                     --                .r
		textmode_vd                  : out   std_logic;                                        --                .vd
		textmode_grest               : out   std_logic;                                        --                .grest
		touch_cntrl_ext_adc_cs       : out   std_logic;                                        -- touch_cntrl_ext.adc_cs
		touch_cntrl_ext_adc_dclk     : out   std_logic;                                        --                .adc_dclk
		touch_cntrl_ext_adc_din      : out   std_logic;                                        --                .adc_din
		touch_cntrl_ext_adc_dout     : in    std_logic                     := '0';             --                .adc_dout
		touch_cntrl_ext_adc_penirq_n : in    std_logic                     := '0'              --                .adc_penirq_n
	);
end entity reverb_template;

architecture rtl of reverb_template is
	component reverb_template_altpll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X';             -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic                                         -- export
		);
	end component reverb_template_altpll;

	component reverb_template_altpll_sram is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component reverb_template_altpll_sram;

	component reverb_template_audio is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component reverb_template_audio;

	component reverb_template_audio_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component reverb_template_audio_pll;

	component reverb_template_av_config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component reverb_template_av_config;

	component fft_wrapper_header is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset_n     : in  std_logic                     := 'X';             -- reset_n
			stin_data   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			stin_valid  : in  std_logic                     := 'X';             -- valid
			stin_ready  : out std_logic;                                        -- ready
			stout_data  : out std_logic_vector(31 downto 0);                    -- data
			stout_ready : in  std_logic                     := 'X';             -- ready
			stout_valid : out std_logic;                                        -- valid
			inverse     : in  std_logic                     := 'X'              -- export
		);
	end component fft_wrapper_header;

	component fir is
		generic (
			NUM_COEFFICIENTS : positive := 512;
			DATA_WIDTH       : positive := 32;
			ADDR_WIDTH       : positive := 9
		);
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			stin_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			stin_valid   : in  std_logic                     := 'X';             -- valid
			stin_ready   : out std_logic;                                        -- ready
			res_n        : in  std_logic                     := 'X';             -- reset_n
			mm_address   : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			mm_write     : in  std_logic                     := 'X';             -- write
			mm_read      : in  std_logic                     := 'X';             -- read
			mm_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			stout_data   : out std_logic_vector(31 downto 0);                    -- data
			stout_ready  : in  std_logic                     := 'X';             -- ready
			stout_valid  : out std_logic                                         -- valid
		);
	end component fir;

	component mac_sram is
		port (
			clk             : in  std_logic                     := 'X';             -- clk
			res_n           : in  std_logic                     := 'X';             -- reset_n
			m_address       : out std_logic_vector(19 downto 0);                    -- address
			m_write         : out std_logic;                                        -- write
			m_read          : out std_logic;                                        -- read
			m_writedata     : out std_logic_vector(15 downto 0);                    -- writedata
			m_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			s_address       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			s_write         : in  std_logic                     := 'X';             -- write
			s_read          : in  std_logic                     := 'X';             -- read
			s_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			sel             : out std_logic                                         -- export
		);
	end component mac_sram;

	component reverb_template_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component reverb_template_jtag_uart;

	component reverb_template_m2s_fifo_ffth is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			reset_n                          : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonst_source_valid            : out std_logic;                                        -- valid
			avalonst_source_data             : out std_logic_vector(31 downto 0);                    -- data
			avalonst_source_ready            : in  std_logic                     := 'X'              -- ready
		);
	end component reverb_template_m2s_fifo_ffth;

	component reverb_template_m2s_fifo_fir_l is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			reset_n                          : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonst_source_valid            : out std_logic;                                        -- valid
			avalonst_source_data             : out std_logic_vector(31 downto 0);                    -- data
			avalonst_source_ready            : in  std_logic                     := 'X'              -- ready
		);
	end component reverb_template_m2s_fifo_fir_l;

	component multiplexer is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			s0_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s1_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			s1_write         : in  std_logic                     := 'X';             -- write
			s1_writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			s1_read          : in  std_logic                     := 'X';             -- read
			s1_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			s1_readdatavalid : out std_logic;                                        -- readdatavalid
			s1_byteanable    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			m_address        : out std_logic_vector(19 downto 0);                    -- address
			m_byteanable     : out std_logic_vector(1 downto 0);                     -- byteenable
			m_write          : out std_logic;                                        -- write
			m_writedata      : out std_logic_vector(15 downto 0);                    -- writedata
			m_read           : out std_logic;                                        -- read
			m_readdata       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m_readdatavalid  : in  std_logic                     := 'X';             -- readdatavalid
			res_n            : in  std_logic                     := 'X';             -- reset_n
			sel              : in  std_logic                     := 'X'              -- export
		);
	end component multiplexer;

	component reverb_template_nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component reverb_template_nios2;

	component reverb_template_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component reverb_template_pio_0;

	component reverb_template_s2m_fifo_ffth is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic                                         -- waitrequest
		);
	end component reverb_template_s2m_fifo_ffth;

	component reverb_template_s2m_fifo_fir_l is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic                                         -- waitrequest
		);
	end component reverb_template_s2m_fifo_fir_l;

	component Altera_UP_SD_Card_Avalon_Interface is
		port (
			i_avalon_chip_select : in    std_logic                     := 'X';             -- chipselect
			i_avalon_address     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			i_avalon_read        : in    std_logic                     := 'X';             -- read
			i_avalon_write       : in    std_logic                     := 'X';             -- write
			i_avalon_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest : out   std_logic;                                        -- waitrequest
			i_clock              : in    std_logic                     := 'X';             -- clk
			i_reset_n            : in    std_logic                     := 'X';             -- reset_n
			b_SD_cmd             : inout std_logic                     := 'X';             -- export
			b_SD_dat             : inout std_logic                     := 'X';             -- export
			b_SD_dat3            : inout std_logic                     := 'X';             -- export
			o_SD_clock           : out   std_logic                                         -- export
		);
	end component Altera_UP_SD_Card_Avalon_Interface;

	component reverb_template_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component reverb_template_sdram;

	component reverb_template_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component reverb_template_sram_0;

	component textmode_controller_avalon is
		generic (
			ROW_COUNT    : integer := 30;
			COLUMN_COUNT : integer := 100;
			CLK_FREQ     : integer := 25000000
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset_n   : in  std_logic                     := 'X';             -- reset_n
			address   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			write_n   : in  std_logic                     := 'X';             -- write_n
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			b         : out std_logic_vector(7 downto 0);                     -- b
			den       : out std_logic;                                        -- den
			g         : out std_logic_vector(7 downto 0);                     -- g
			hd        : out std_logic;                                        -- hd
			r         : out std_logic_vector(7 downto 0);                     -- r
			vd        : out std_logic;                                        -- vd
			grest     : out std_logic;                                        -- grest
			irq       : out std_logic                                         -- irq
		);
	end component textmode_controller_avalon;

	component avalon_touch_cntrl is
		generic (
			SYS_CLK : integer := 100000000
		);
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			adc_cs       : out std_logic;                                        -- adc_cs
			adc_dclk     : out std_logic;                                        -- adc_dclk
			adc_din      : out std_logic;                                        -- adc_din
			adc_dout     : in  std_logic                     := 'X';             -- adc_dout
			adc_penirq_n : in  std_logic                     := 'X';             -- adc_penirq_n
			irq          : out std_logic;                                        -- irq
			address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write        : in  std_logic                     := 'X';             -- write
			read         : in  std_logic                     := 'X';             -- read
			writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			res_n        : in  std_logic                     := 'X'              -- reset_n
		);
	end component avalon_touch_cntrl;

	component reverb_template_mm_interconnect_2 is
		port (
			altpll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			altpll_c2_clk                                            : in  std_logic                     := 'X';             -- clk
			altpll_sram_c0_clk                                       : in  std_logic                     := 'X';             -- clk
			sys_clk_clk_clk                                          : in  std_logic                     := 'X';             -- clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			audio_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			header_mac_0_reset_sink_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			nios2_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			sdcard_interface_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			textmode_controller_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			nios2_data_master_address                                : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest                            : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                                   : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_readdatavalid                          : out std_logic;                                        -- readdatavalid
			nios2_data_master_write                                  : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess                            : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address                         : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest                     : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read                            : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_instruction_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			altpll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			altpll_sram_pll_slave_address                            : out std_logic_vector(1 downto 0);                     -- address
			altpll_sram_pll_slave_write                              : out std_logic;                                        -- write
			altpll_sram_pll_slave_read                               : out std_logic;                                        -- read
			altpll_sram_pll_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_sram_pll_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			audio_avalon_audio_slave_address                         : out std_logic_vector(1 downto 0);                     -- address
			audio_avalon_audio_slave_write                           : out std_logic;                                        -- write
			audio_avalon_audio_slave_read                            : out std_logic;                                        -- read
			audio_avalon_audio_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_avalon_audio_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			audio_avalon_audio_slave_chipselect                      : out std_logic;                                        -- chipselect
			av_config_avalon_av_config_slave_address                 : out std_logic_vector(1 downto 0);                     -- address
			av_config_avalon_av_config_slave_write                   : out std_logic;                                        -- write
			av_config_avalon_av_config_slave_read                    : out std_logic;                                        -- read
			av_config_avalon_av_config_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_config_avalon_av_config_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			av_config_avalon_av_config_slave_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			av_config_avalon_av_config_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			fir_l_avalon_slave_0_address                             : out std_logic_vector(8 downto 0);                     -- address
			fir_l_avalon_slave_0_write                               : out std_logic;                                        -- write
			fir_l_avalon_slave_0_read                                : out std_logic;                                        -- read
			fir_l_avalon_slave_0_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fir_l_avalon_slave_0_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			fir_r_avalon_slave_0_address                             : out std_logic_vector(8 downto 0);                     -- address
			fir_r_avalon_slave_0_write                               : out std_logic;                                        -- write
			fir_r_avalon_slave_0_read                                : out std_logic;                                        -- read
			fir_r_avalon_slave_0_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fir_r_avalon_slave_0_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			header_mac_0_avalon_slave_address                        : out std_logic_vector(15 downto 0);                    -- address
			header_mac_0_avalon_slave_write                          : out std_logic;                                        -- write
			header_mac_0_avalon_slave_read                           : out std_logic;                                        -- read
			header_mac_0_avalon_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			header_mac_0_avalon_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			m2s_fifo_ffth_in_address                                 : out std_logic_vector(0 downto 0);                     -- address
			m2s_fifo_ffth_in_write                                   : out std_logic;                                        -- write
			m2s_fifo_ffth_in_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			m2s_fifo_ffth_in_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			m2s_fifo_fir_l_in_address                                : out std_logic_vector(0 downto 0);                     -- address
			m2s_fifo_fir_l_in_write                                  : out std_logic;                                        -- write
			m2s_fifo_fir_l_in_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			m2s_fifo_fir_l_in_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			m2s_fifo_fir_r_in_address                                : out std_logic_vector(0 downto 0);                     -- address
			m2s_fifo_fir_r_in_write                                  : out std_logic;                                        -- write
			m2s_fifo_fir_r_in_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			m2s_fifo_fir_r_in_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			multiplexer_sram_0_s1_address                            : out std_logic_vector(19 downto 0);                    -- address
			multiplexer_sram_0_s1_write                              : out std_logic;                                        -- write
			multiplexer_sram_0_s1_read                               : out std_logic;                                        -- read
			multiplexer_sram_0_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			multiplexer_sram_0_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			multiplexer_sram_0_s1_byteenable                         : out std_logic_vector(1 downto 0);                     -- byteenable
			multiplexer_sram_0_s1_readdatavalid                      : in  std_logic                     := 'X';             -- readdatavalid
			nios2_debug_mem_slave_address                            : out std_logic_vector(8 downto 0);                     -- address
			nios2_debug_mem_slave_write                              : out std_logic;                                        -- write
			nios2_debug_mem_slave_read                               : out std_logic;                                        -- read
			nios2_debug_mem_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_debug_mem_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_debug_mem_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_debug_mem_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			nios2_debug_mem_slave_debugaccess                        : out std_logic;                                        -- debugaccess
			pio_0_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			pio_0_s1_write                                           : out std_logic;                                        -- write
			pio_0_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                      : out std_logic;                                        -- chipselect
			s2m_fifo_ffth_out_address                                : out std_logic_vector(0 downto 0);                     -- address
			s2m_fifo_ffth_out_read                                   : out std_logic;                                        -- read
			s2m_fifo_ffth_out_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			s2m_fifo_ffth_out_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			s2m_fifo_fir_l_out_address                               : out std_logic_vector(0 downto 0);                     -- address
			s2m_fifo_fir_l_out_read                                  : out std_logic;                                        -- read
			s2m_fifo_fir_l_out_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			s2m_fifo_fir_l_out_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			s2m_fifo_fir_r_out_address                               : out std_logic_vector(0 downto 0);                     -- address
			s2m_fifo_fir_r_out_read                                  : out std_logic;                                        -- read
			s2m_fifo_fir_r_out_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			s2m_fifo_fir_r_out_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			sdcard_interface_avalon_sdcard_slave_address             : out std_logic_vector(7 downto 0);                     -- address
			sdcard_interface_avalon_sdcard_slave_write               : out std_logic;                                        -- write
			sdcard_interface_avalon_sdcard_slave_read                : out std_logic;                                        -- read
			sdcard_interface_avalon_sdcard_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdcard_interface_avalon_sdcard_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			sdcard_interface_avalon_sdcard_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			sdcard_interface_avalon_sdcard_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			sdcard_interface_avalon_sdcard_slave_chipselect          : out std_logic;                                        -- chipselect
			sdram_s1_address                                         : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                           : out std_logic;                                        -- write
			sdram_s1_read                                            : out std_logic;                                        -- read
			sdram_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_byteenable                                      : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                   : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                      : out std_logic;                                        -- chipselect
			textmode_controller_avalon_slave_address                 : out std_logic_vector(3 downto 0);                     -- address
			textmode_controller_avalon_slave_write                   : out std_logic;                                        -- write
			textmode_controller_avalon_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			textmode_controller_avalon_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			touch_cntrl_avalon_slave_address                         : out std_logic_vector(1 downto 0);                     -- address
			touch_cntrl_avalon_slave_write                           : out std_logic;                                        -- write
			touch_cntrl_avalon_slave_read                            : out std_logic;                                        -- read
			touch_cntrl_avalon_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			touch_cntrl_avalon_slave_writedata                       : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component reverb_template_mm_interconnect_2;

	component reverb_template_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component reverb_template_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component reverb_template_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component reverb_template_avalon_st_adapter;

	component reverb_template_avalon_st_adapter_003 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component reverb_template_avalon_st_adapter_003;

	component reverb_template_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component reverb_template_rst_controller;

	component reverb_template_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component reverb_template_rst_controller_001;

	signal multiplexer_sram_0_avalon_master_readdata                          : std_logic_vector(15 downto 0); -- sram_0:readdata -> multiplexer_sram_0:m_readdata
	signal multiplexer_sram_0_avalon_master_address                           : std_logic_vector(19 downto 0); -- multiplexer_sram_0:m_address -> sram_0:address
	signal multiplexer_sram_0_avalon_master_byteenable                        : std_logic_vector(1 downto 0);  -- multiplexer_sram_0:m_byteanable -> sram_0:byteenable
	signal multiplexer_sram_0_avalon_master_read                              : std_logic;                     -- multiplexer_sram_0:m_read -> sram_0:read
	signal multiplexer_sram_0_avalon_master_readdatavalid                     : std_logic;                     -- sram_0:readdatavalid -> multiplexer_sram_0:m_readdatavalid
	signal multiplexer_sram_0_avalon_master_write                             : std_logic;                     -- multiplexer_sram_0:m_write -> sram_0:write
	signal multiplexer_sram_0_avalon_master_writedata                         : std_logic_vector(15 downto 0); -- multiplexer_sram_0:m_writedata -> sram_0:writedata
	signal header_mac_0_avalon_master_readdata                                : std_logic_vector(15 downto 0); -- multiplexer_sram_0:s0_readdata -> header_mac_0:m_readdata
	signal header_mac_0_avalon_master_address                                 : std_logic_vector(19 downto 0); -- header_mac_0:m_address -> multiplexer_sram_0:s0_address
	signal header_mac_0_avalon_master_read                                    : std_logic;                     -- header_mac_0:m_read -> multiplexer_sram_0:s0_read
	signal header_mac_0_avalon_master_readdatavalid                           : std_logic;                     -- multiplexer_sram_0:s0_readdatavalid -> header_mac_0:m_readdatavalid
	signal header_mac_0_avalon_master_write                                   : std_logic;                     -- header_mac_0:m_write -> multiplexer_sram_0:s0_write
	signal header_mac_0_avalon_master_writedata                               : std_logic_vector(15 downto 0); -- header_mac_0:m_writedata -> multiplexer_sram_0:s0_writedata
	signal altpll_c0_clk                                                      : std_logic;                     -- altpll:c0 -> [sdram_clk_clk, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, avalon_st_adapter_002:in_clk_0_clk, avalon_st_adapter_003:in_clk_0_clk, avalon_st_adapter_004:in_clk_0_clk, avalon_st_adapter_005:in_clk_0_clk, fft_wrapper_header_0:clk, fir_l:clk, fir_r:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, m2s_fifo_ffth:wrclock, m2s_fifo_fir_l:wrclock, m2s_fifo_fir_r:wrclock, mm_interconnect_2:altpll_c0_clk, nios2:clk, pio_0:clk, rst_controller_002:clk, rst_controller_004:clk, s2m_fifo_ffth:wrclock, s2m_fifo_fir_l:wrclock, s2m_fifo_fir_r:wrclock, sdcard_interface:i_clock, sdram:clk, touch_cntrl:clk]
	signal altpll_sram_c0_clk                                                 : std_logic;                     -- altpll_sram:c0 -> [header_mac_0:clk, mm_interconnect_2:altpll_sram_c0_clk, multiplexer_sram_0:clk, rst_controller_003:clk, rst_controller_005:clk, sram_0:clk]
	signal altpll_c2_clk                                                      : std_logic;                     -- altpll:c2 -> [clk_25_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_2:altpll_c2_clk, rst_controller_006:clk, textmode_controller:clk]
	signal pio_0_external_connection_export                                   : std_logic;                     -- pio_0:out_port -> fft_wrapper_header_0:inverse
	signal header_mac_0_sel_export                                            : std_logic;                     -- header_mac_0:sel -> multiplexer_sram_0:sel
	signal nios2_data_master_readdata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                                      : std_logic;                     -- mm_interconnect_2:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                      : std_logic;                     -- nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_2:nios2_data_master_debugaccess
	signal nios2_data_master_address                                          : std_logic_vector(28 downto 0); -- nios2:d_address -> mm_interconnect_2:nios2_data_master_address
	signal nios2_data_master_byteenable                                       : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_2:nios2_data_master_byteenable
	signal nios2_data_master_read                                             : std_logic;                     -- nios2:d_read -> mm_interconnect_2:nios2_data_master_read
	signal nios2_data_master_readdatavalid                                    : std_logic;                     -- mm_interconnect_2:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	signal nios2_data_master_write                                            : std_logic;                     -- nios2:d_write -> mm_interconnect_2:nios2_data_master_write
	signal nios2_data_master_writedata                                        : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_2:nios2_data_master_writedata
	signal nios2_instruction_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                               : std_logic;                     -- mm_interconnect_2:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                                   : std_logic_vector(28 downto 0); -- nios2:i_address -> mm_interconnect_2:nios2_instruction_master_address
	signal nios2_instruction_master_read                                      : std_logic;                     -- nios2:i_read -> mm_interconnect_2:nios2_instruction_master_read
	signal nios2_instruction_master_readdatavalid                             : std_logic;                     -- mm_interconnect_2:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	signal mm_interconnect_2_audio_avalon_audio_slave_chipselect              : std_logic;                     -- mm_interconnect_2:audio_avalon_audio_slave_chipselect -> audio:chipselect
	signal mm_interconnect_2_audio_avalon_audio_slave_readdata                : std_logic_vector(31 downto 0); -- audio:readdata -> mm_interconnect_2:audio_avalon_audio_slave_readdata
	signal mm_interconnect_2_audio_avalon_audio_slave_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:audio_avalon_audio_slave_address -> audio:address
	signal mm_interconnect_2_audio_avalon_audio_slave_read                    : std_logic;                     -- mm_interconnect_2:audio_avalon_audio_slave_read -> audio:read
	signal mm_interconnect_2_audio_avalon_audio_slave_write                   : std_logic;                     -- mm_interconnect_2:audio_avalon_audio_slave_write -> audio:write
	signal mm_interconnect_2_audio_avalon_audio_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_2:audio_avalon_audio_slave_writedata -> audio:writedata
	signal mm_interconnect_2_av_config_avalon_av_config_slave_readdata        : std_logic_vector(31 downto 0); -- av_config:readdata -> mm_interconnect_2:av_config_avalon_av_config_slave_readdata
	signal mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest     : std_logic;                     -- av_config:waitrequest -> mm_interconnect_2:av_config_avalon_av_config_slave_waitrequest
	signal mm_interconnect_2_av_config_avalon_av_config_slave_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_2:av_config_avalon_av_config_slave_address -> av_config:address
	signal mm_interconnect_2_av_config_avalon_av_config_slave_read            : std_logic;                     -- mm_interconnect_2:av_config_avalon_av_config_slave_read -> av_config:read
	signal mm_interconnect_2_av_config_avalon_av_config_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_2:av_config_avalon_av_config_slave_byteenable -> av_config:byteenable
	signal mm_interconnect_2_av_config_avalon_av_config_slave_write           : std_logic;                     -- mm_interconnect_2:av_config_avalon_av_config_slave_write -> av_config:write
	signal mm_interconnect_2_av_config_avalon_av_config_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_2:av_config_avalon_av_config_slave_writedata -> av_config:writedata
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_2:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_2:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest          : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_2:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_2:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_2:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_2_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_2:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_2_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_2:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_chipselect  : std_logic;                     -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_chipselect -> sdcard_interface:i_avalon_chip_select
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_readdata    : std_logic_vector(31 downto 0); -- sdcard_interface:o_avalon_readdata -> mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_readdata
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_waitrequest : std_logic;                     -- sdcard_interface:o_avalon_waitrequest -> mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_waitrequest
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_address     : std_logic_vector(7 downto 0);  -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_address -> sdcard_interface:i_avalon_address
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_read        : std_logic;                     -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_read -> sdcard_interface:i_avalon_read
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_byteenable -> sdcard_interface:i_avalon_byteenable
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_write       : std_logic;                     -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_write -> sdcard_interface:i_avalon_write
	signal mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_2:sdcard_interface_avalon_sdcard_slave_writedata -> sdcard_interface:i_avalon_writedata
	signal mm_interconnect_2_textmode_controller_avalon_slave_readdata        : std_logic_vector(31 downto 0); -- textmode_controller:readdata -> mm_interconnect_2:textmode_controller_avalon_slave_readdata
	signal mm_interconnect_2_textmode_controller_avalon_slave_address         : std_logic_vector(3 downto 0);  -- mm_interconnect_2:textmode_controller_avalon_slave_address -> textmode_controller:address
	signal mm_interconnect_2_textmode_controller_avalon_slave_write           : std_logic;                     -- mm_interconnect_2:textmode_controller_avalon_slave_write -> mm_interconnect_2_textmode_controller_avalon_slave_write:in
	signal mm_interconnect_2_textmode_controller_avalon_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_2:textmode_controller_avalon_slave_writedata -> textmode_controller:writedata
	signal mm_interconnect_2_touch_cntrl_avalon_slave_readdata                : std_logic_vector(31 downto 0); -- touch_cntrl:readdata -> mm_interconnect_2:touch_cntrl_avalon_slave_readdata
	signal mm_interconnect_2_touch_cntrl_avalon_slave_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:touch_cntrl_avalon_slave_address -> touch_cntrl:address
	signal mm_interconnect_2_touch_cntrl_avalon_slave_read                    : std_logic;                     -- mm_interconnect_2:touch_cntrl_avalon_slave_read -> touch_cntrl:read
	signal mm_interconnect_2_touch_cntrl_avalon_slave_write                   : std_logic;                     -- mm_interconnect_2:touch_cntrl_avalon_slave_write -> touch_cntrl:write
	signal mm_interconnect_2_touch_cntrl_avalon_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_2:touch_cntrl_avalon_slave_writedata -> touch_cntrl:writedata
	signal mm_interconnect_2_header_mac_0_avalon_slave_readdata               : std_logic_vector(31 downto 0); -- header_mac_0:s_readdata -> mm_interconnect_2:header_mac_0_avalon_slave_readdata
	signal mm_interconnect_2_header_mac_0_avalon_slave_address                : std_logic_vector(15 downto 0); -- mm_interconnect_2:header_mac_0_avalon_slave_address -> header_mac_0:s_address
	signal mm_interconnect_2_header_mac_0_avalon_slave_read                   : std_logic;                     -- mm_interconnect_2:header_mac_0_avalon_slave_read -> header_mac_0:s_read
	signal mm_interconnect_2_header_mac_0_avalon_slave_write                  : std_logic;                     -- mm_interconnect_2:header_mac_0_avalon_slave_write -> header_mac_0:s_write
	signal mm_interconnect_2_header_mac_0_avalon_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_2:header_mac_0_avalon_slave_writedata -> header_mac_0:s_writedata
	signal mm_interconnect_2_fir_l_avalon_slave_0_readdata                    : std_logic_vector(31 downto 0); -- fir_l:mm_readdata -> mm_interconnect_2:fir_l_avalon_slave_0_readdata
	signal mm_interconnect_2_fir_l_avalon_slave_0_address                     : std_logic_vector(8 downto 0);  -- mm_interconnect_2:fir_l_avalon_slave_0_address -> fir_l:mm_address
	signal mm_interconnect_2_fir_l_avalon_slave_0_read                        : std_logic;                     -- mm_interconnect_2:fir_l_avalon_slave_0_read -> fir_l:mm_read
	signal mm_interconnect_2_fir_l_avalon_slave_0_write                       : std_logic;                     -- mm_interconnect_2:fir_l_avalon_slave_0_write -> fir_l:mm_write
	signal mm_interconnect_2_fir_l_avalon_slave_0_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_2:fir_l_avalon_slave_0_writedata -> fir_l:mm_writedata
	signal mm_interconnect_2_fir_r_avalon_slave_0_readdata                    : std_logic_vector(31 downto 0); -- fir_r:mm_readdata -> mm_interconnect_2:fir_r_avalon_slave_0_readdata
	signal mm_interconnect_2_fir_r_avalon_slave_0_address                     : std_logic_vector(8 downto 0);  -- mm_interconnect_2:fir_r_avalon_slave_0_address -> fir_r:mm_address
	signal mm_interconnect_2_fir_r_avalon_slave_0_read                        : std_logic;                     -- mm_interconnect_2:fir_r_avalon_slave_0_read -> fir_r:mm_read
	signal mm_interconnect_2_fir_r_avalon_slave_0_write                       : std_logic;                     -- mm_interconnect_2:fir_r_avalon_slave_0_write -> fir_r:mm_write
	signal mm_interconnect_2_fir_r_avalon_slave_0_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_2:fir_r_avalon_slave_0_writedata -> fir_r:mm_writedata
	signal mm_interconnect_2_nios2_debug_mem_slave_readdata                   : std_logic_vector(31 downto 0); -- nios2:debug_mem_slave_readdata -> mm_interconnect_2:nios2_debug_mem_slave_readdata
	signal mm_interconnect_2_nios2_debug_mem_slave_waitrequest                : std_logic;                     -- nios2:debug_mem_slave_waitrequest -> mm_interconnect_2:nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_2_nios2_debug_mem_slave_debugaccess                : std_logic;                     -- mm_interconnect_2:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_2_nios2_debug_mem_slave_address                    : std_logic_vector(8 downto 0);  -- mm_interconnect_2:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	signal mm_interconnect_2_nios2_debug_mem_slave_read                       : std_logic;                     -- mm_interconnect_2:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	signal mm_interconnect_2_nios2_debug_mem_slave_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_2:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	signal mm_interconnect_2_nios2_debug_mem_slave_write                      : std_logic;                     -- mm_interconnect_2:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	signal mm_interconnect_2_nios2_debug_mem_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	signal mm_interconnect_2_m2s_fifo_ffth_in_waitrequest                     : std_logic;                     -- m2s_fifo_ffth:avalonmm_write_slave_waitrequest -> mm_interconnect_2:m2s_fifo_ffth_in_waitrequest
	signal mm_interconnect_2_m2s_fifo_ffth_in_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_2:m2s_fifo_ffth_in_address -> m2s_fifo_ffth:avalonmm_write_slave_address
	signal mm_interconnect_2_m2s_fifo_ffth_in_write                           : std_logic;                     -- mm_interconnect_2:m2s_fifo_ffth_in_write -> m2s_fifo_ffth:avalonmm_write_slave_write
	signal mm_interconnect_2_m2s_fifo_ffth_in_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_2:m2s_fifo_ffth_in_writedata -> m2s_fifo_ffth:avalonmm_write_slave_writedata
	signal mm_interconnect_2_m2s_fifo_fir_l_in_waitrequest                    : std_logic;                     -- m2s_fifo_fir_l:avalonmm_write_slave_waitrequest -> mm_interconnect_2:m2s_fifo_fir_l_in_waitrequest
	signal mm_interconnect_2_m2s_fifo_fir_l_in_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_2:m2s_fifo_fir_l_in_address -> m2s_fifo_fir_l:avalonmm_write_slave_address
	signal mm_interconnect_2_m2s_fifo_fir_l_in_write                          : std_logic;                     -- mm_interconnect_2:m2s_fifo_fir_l_in_write -> m2s_fifo_fir_l:avalonmm_write_slave_write
	signal mm_interconnect_2_m2s_fifo_fir_l_in_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_2:m2s_fifo_fir_l_in_writedata -> m2s_fifo_fir_l:avalonmm_write_slave_writedata
	signal mm_interconnect_2_m2s_fifo_fir_r_in_waitrequest                    : std_logic;                     -- m2s_fifo_fir_r:avalonmm_write_slave_waitrequest -> mm_interconnect_2:m2s_fifo_fir_r_in_waitrequest
	signal mm_interconnect_2_m2s_fifo_fir_r_in_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_2:m2s_fifo_fir_r_in_address -> m2s_fifo_fir_r:avalonmm_write_slave_address
	signal mm_interconnect_2_m2s_fifo_fir_r_in_write                          : std_logic;                     -- mm_interconnect_2:m2s_fifo_fir_r_in_write -> m2s_fifo_fir_r:avalonmm_write_slave_write
	signal mm_interconnect_2_m2s_fifo_fir_r_in_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_2:m2s_fifo_fir_r_in_writedata -> m2s_fifo_fir_r:avalonmm_write_slave_writedata
	signal mm_interconnect_2_s2m_fifo_ffth_out_readdata                       : std_logic_vector(31 downto 0); -- s2m_fifo_ffth:avalonmm_read_slave_readdata -> mm_interconnect_2:s2m_fifo_ffth_out_readdata
	signal mm_interconnect_2_s2m_fifo_ffth_out_waitrequest                    : std_logic;                     -- s2m_fifo_ffth:avalonmm_read_slave_waitrequest -> mm_interconnect_2:s2m_fifo_ffth_out_waitrequest
	signal mm_interconnect_2_s2m_fifo_ffth_out_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_2:s2m_fifo_ffth_out_address -> s2m_fifo_ffth:avalonmm_read_slave_address
	signal mm_interconnect_2_s2m_fifo_ffth_out_read                           : std_logic;                     -- mm_interconnect_2:s2m_fifo_ffth_out_read -> s2m_fifo_ffth:avalonmm_read_slave_read
	signal mm_interconnect_2_s2m_fifo_fir_l_out_readdata                      : std_logic_vector(31 downto 0); -- s2m_fifo_fir_l:avalonmm_read_slave_readdata -> mm_interconnect_2:s2m_fifo_fir_l_out_readdata
	signal mm_interconnect_2_s2m_fifo_fir_l_out_waitrequest                   : std_logic;                     -- s2m_fifo_fir_l:avalonmm_read_slave_waitrequest -> mm_interconnect_2:s2m_fifo_fir_l_out_waitrequest
	signal mm_interconnect_2_s2m_fifo_fir_l_out_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_2:s2m_fifo_fir_l_out_address -> s2m_fifo_fir_l:avalonmm_read_slave_address
	signal mm_interconnect_2_s2m_fifo_fir_l_out_read                          : std_logic;                     -- mm_interconnect_2:s2m_fifo_fir_l_out_read -> s2m_fifo_fir_l:avalonmm_read_slave_read
	signal mm_interconnect_2_s2m_fifo_fir_r_out_readdata                      : std_logic_vector(31 downto 0); -- s2m_fifo_fir_r:avalonmm_read_slave_readdata -> mm_interconnect_2:s2m_fifo_fir_r_out_readdata
	signal mm_interconnect_2_s2m_fifo_fir_r_out_waitrequest                   : std_logic;                     -- s2m_fifo_fir_r:avalonmm_read_slave_waitrequest -> mm_interconnect_2:s2m_fifo_fir_r_out_waitrequest
	signal mm_interconnect_2_s2m_fifo_fir_r_out_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_2:s2m_fifo_fir_r_out_address -> s2m_fifo_fir_r:avalonmm_read_slave_address
	signal mm_interconnect_2_s2m_fifo_fir_r_out_read                          : std_logic;                     -- mm_interconnect_2:s2m_fifo_fir_r_out_read -> s2m_fifo_fir_r:avalonmm_read_slave_read
	signal mm_interconnect_2_altpll_sram_pll_slave_readdata                   : std_logic_vector(31 downto 0); -- altpll_sram:readdata -> mm_interconnect_2:altpll_sram_pll_slave_readdata
	signal mm_interconnect_2_altpll_sram_pll_slave_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_2:altpll_sram_pll_slave_address -> altpll_sram:address
	signal mm_interconnect_2_altpll_sram_pll_slave_read                       : std_logic;                     -- mm_interconnect_2:altpll_sram_pll_slave_read -> altpll_sram:read
	signal mm_interconnect_2_altpll_sram_pll_slave_write                      : std_logic;                     -- mm_interconnect_2:altpll_sram_pll_slave_write -> altpll_sram:write
	signal mm_interconnect_2_altpll_sram_pll_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_2:altpll_sram_pll_slave_writedata -> altpll_sram:writedata
	signal mm_interconnect_2_altpll_pll_slave_readdata                        : std_logic_vector(31 downto 0); -- altpll:readdata -> mm_interconnect_2:altpll_pll_slave_readdata
	signal mm_interconnect_2_altpll_pll_slave_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_2:altpll_pll_slave_address -> altpll:address
	signal mm_interconnect_2_altpll_pll_slave_read                            : std_logic;                     -- mm_interconnect_2:altpll_pll_slave_read -> altpll:read
	signal mm_interconnect_2_altpll_pll_slave_write                           : std_logic;                     -- mm_interconnect_2:altpll_pll_slave_write -> altpll:write
	signal mm_interconnect_2_altpll_pll_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_2:altpll_pll_slave_writedata -> altpll:writedata
	signal mm_interconnect_2_sdram_s1_chipselect                              : std_logic;                     -- mm_interconnect_2:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_2_sdram_s1_readdata                                : std_logic_vector(31 downto 0); -- sdram:za_data -> mm_interconnect_2:sdram_s1_readdata
	signal mm_interconnect_2_sdram_s1_waitrequest                             : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_2:sdram_s1_waitrequest
	signal mm_interconnect_2_sdram_s1_address                                 : std_logic_vector(24 downto 0); -- mm_interconnect_2:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_2_sdram_s1_read                                    : std_logic;                     -- mm_interconnect_2:sdram_s1_read -> mm_interconnect_2_sdram_s1_read:in
	signal mm_interconnect_2_sdram_s1_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_2:sdram_s1_byteenable -> mm_interconnect_2_sdram_s1_byteenable:in
	signal mm_interconnect_2_sdram_s1_readdatavalid                           : std_logic;                     -- sdram:za_valid -> mm_interconnect_2:sdram_s1_readdatavalid
	signal mm_interconnect_2_sdram_s1_write                                   : std_logic;                     -- mm_interconnect_2:sdram_s1_write -> mm_interconnect_2_sdram_s1_write:in
	signal mm_interconnect_2_sdram_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_2:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_2_pio_0_s1_chipselect                              : std_logic;                     -- mm_interconnect_2:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_2_pio_0_s1_readdata                                : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_2:pio_0_s1_readdata
	signal mm_interconnect_2_pio_0_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_2_pio_0_s1_write                                   : std_logic;                     -- mm_interconnect_2:pio_0_s1_write -> mm_interconnect_2_pio_0_s1_write:in
	signal mm_interconnect_2_pio_0_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_2:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_2_multiplexer_sram_0_s1_readdata                   : std_logic_vector(15 downto 0); -- multiplexer_sram_0:s1_readdata -> mm_interconnect_2:multiplexer_sram_0_s1_readdata
	signal mm_interconnect_2_multiplexer_sram_0_s1_address                    : std_logic_vector(19 downto 0); -- mm_interconnect_2:multiplexer_sram_0_s1_address -> multiplexer_sram_0:s1_address
	signal mm_interconnect_2_multiplexer_sram_0_s1_read                       : std_logic;                     -- mm_interconnect_2:multiplexer_sram_0_s1_read -> multiplexer_sram_0:s1_read
	signal mm_interconnect_2_multiplexer_sram_0_s1_byteenable                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:multiplexer_sram_0_s1_byteenable -> multiplexer_sram_0:s1_byteanable
	signal mm_interconnect_2_multiplexer_sram_0_s1_readdatavalid              : std_logic;                     -- multiplexer_sram_0:s1_readdatavalid -> mm_interconnect_2:multiplexer_sram_0_s1_readdatavalid
	signal mm_interconnect_2_multiplexer_sram_0_s1_write                      : std_logic;                     -- mm_interconnect_2:multiplexer_sram_0_s1_write -> multiplexer_sram_0:s1_write
	signal mm_interconnect_2_multiplexer_sram_0_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_2:multiplexer_sram_0_s1_writedata -> multiplexer_sram_0:s1_writedata
	signal irq_mapper_receiver2_irq                                           : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                           : std_logic;                     -- touch_cntrl:irq -> irq_mapper:receiver3_irq
	signal nios2_irq_irq                                                      : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:irq
	signal irq_mapper_receiver0_irq                                           : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                      : std_logic_vector(0 downto 0);  -- audio:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                           : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                                  : std_logic_vector(0 downto 0);  -- textmode_controller:irq -> irq_synchronizer_001:receiver_irq
	signal fft_wrapper_header_0_avalon_streaming_source_valid                 : std_logic;                     -- fft_wrapper_header_0:stout_valid -> avalon_st_adapter:in_0_valid
	signal fft_wrapper_header_0_avalon_streaming_source_data                  : std_logic_vector(31 downto 0); -- fft_wrapper_header_0:stout_data -> avalon_st_adapter:in_0_data
	signal fft_wrapper_header_0_avalon_streaming_source_ready                 : std_logic;                     -- avalon_st_adapter:in_0_ready -> fft_wrapper_header_0:stout_ready
	signal avalon_st_adapter_out_0_valid                                      : std_logic;                     -- avalon_st_adapter:out_0_valid -> s2m_fifo_ffth:avalonst_sink_valid
	signal avalon_st_adapter_out_0_data                                       : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> s2m_fifo_ffth:avalonst_sink_data
	signal avalon_st_adapter_out_0_ready                                      : std_logic;                     -- s2m_fifo_ffth:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	signal fir_l_avalon_streaming_source_valid                                : std_logic;                     -- fir_l:stout_valid -> avalon_st_adapter_001:in_0_valid
	signal fir_l_avalon_streaming_source_data                                 : std_logic_vector(31 downto 0); -- fir_l:stout_data -> avalon_st_adapter_001:in_0_data
	signal fir_l_avalon_streaming_source_ready                                : std_logic;                     -- avalon_st_adapter_001:in_0_ready -> fir_l:stout_ready
	signal avalon_st_adapter_001_out_0_valid                                  : std_logic;                     -- avalon_st_adapter_001:out_0_valid -> s2m_fifo_fir_l:avalonst_sink_valid
	signal avalon_st_adapter_001_out_0_data                                   : std_logic_vector(31 downto 0); -- avalon_st_adapter_001:out_0_data -> s2m_fifo_fir_l:avalonst_sink_data
	signal avalon_st_adapter_001_out_0_ready                                  : std_logic;                     -- s2m_fifo_fir_l:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	signal fir_r_avalon_streaming_source_valid                                : std_logic;                     -- fir_r:stout_valid -> avalon_st_adapter_002:in_0_valid
	signal fir_r_avalon_streaming_source_data                                 : std_logic_vector(31 downto 0); -- fir_r:stout_data -> avalon_st_adapter_002:in_0_data
	signal fir_r_avalon_streaming_source_ready                                : std_logic;                     -- avalon_st_adapter_002:in_0_ready -> fir_r:stout_ready
	signal avalon_st_adapter_002_out_0_valid                                  : std_logic;                     -- avalon_st_adapter_002:out_0_valid -> s2m_fifo_fir_r:avalonst_sink_valid
	signal avalon_st_adapter_002_out_0_data                                   : std_logic_vector(31 downto 0); -- avalon_st_adapter_002:out_0_data -> s2m_fifo_fir_r:avalonst_sink_data
	signal avalon_st_adapter_002_out_0_ready                                  : std_logic;                     -- s2m_fifo_fir_r:avalonst_sink_ready -> avalon_st_adapter_002:out_0_ready
	signal m2s_fifo_ffth_out_valid                                            : std_logic;                     -- m2s_fifo_ffth:avalonst_source_valid -> avalon_st_adapter_003:in_0_valid
	signal m2s_fifo_ffth_out_data                                             : std_logic_vector(31 downto 0); -- m2s_fifo_ffth:avalonst_source_data -> avalon_st_adapter_003:in_0_data
	signal m2s_fifo_ffth_out_ready                                            : std_logic;                     -- avalon_st_adapter_003:in_0_ready -> m2s_fifo_ffth:avalonst_source_ready
	signal avalon_st_adapter_003_out_0_valid                                  : std_logic;                     -- avalon_st_adapter_003:out_0_valid -> fft_wrapper_header_0:stin_valid
	signal avalon_st_adapter_003_out_0_data                                   : std_logic_vector(31 downto 0); -- avalon_st_adapter_003:out_0_data -> fft_wrapper_header_0:stin_data
	signal avalon_st_adapter_003_out_0_ready                                  : std_logic;                     -- fft_wrapper_header_0:stin_ready -> avalon_st_adapter_003:out_0_ready
	signal m2s_fifo_fir_l_out_valid                                           : std_logic;                     -- m2s_fifo_fir_l:avalonst_source_valid -> avalon_st_adapter_004:in_0_valid
	signal m2s_fifo_fir_l_out_data                                            : std_logic_vector(31 downto 0); -- m2s_fifo_fir_l:avalonst_source_data -> avalon_st_adapter_004:in_0_data
	signal m2s_fifo_fir_l_out_ready                                           : std_logic;                     -- avalon_st_adapter_004:in_0_ready -> m2s_fifo_fir_l:avalonst_source_ready
	signal avalon_st_adapter_004_out_0_valid                                  : std_logic;                     -- avalon_st_adapter_004:out_0_valid -> fir_l:stin_valid
	signal avalon_st_adapter_004_out_0_data                                   : std_logic_vector(31 downto 0); -- avalon_st_adapter_004:out_0_data -> fir_l:stin_data
	signal avalon_st_adapter_004_out_0_ready                                  : std_logic;                     -- fir_l:stin_ready -> avalon_st_adapter_004:out_0_ready
	signal m2s_fifo_fir_r_out_valid                                           : std_logic;                     -- m2s_fifo_fir_r:avalonst_source_valid -> avalon_st_adapter_005:in_0_valid
	signal m2s_fifo_fir_r_out_data                                            : std_logic_vector(31 downto 0); -- m2s_fifo_fir_r:avalonst_source_data -> avalon_st_adapter_005:in_0_data
	signal m2s_fifo_fir_r_out_ready                                           : std_logic;                     -- avalon_st_adapter_005:in_0_ready -> m2s_fifo_fir_r:avalonst_source_ready
	signal avalon_st_adapter_005_out_0_valid                                  : std_logic;                     -- avalon_st_adapter_005:out_0_valid -> fir_r:stin_valid
	signal avalon_st_adapter_005_out_0_data                                   : std_logic_vector(31 downto 0); -- avalon_st_adapter_005:out_0_data -> fir_r:stin_data
	signal avalon_st_adapter_005_out_0_ready                                  : std_logic;                     -- fir_r:stin_ready -> avalon_st_adapter_005:out_0_ready
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [altpll:reset, altpll_sram:reset, mm_interconnect_2:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal nios2_debug_reset_request_reset                                    : std_logic;                     -- nios2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1]
	signal rst_controller_001_reset_out_reset                                 : std_logic;                     -- rst_controller_001:reset_out -> [audio:reset, audio_pll:ref_reset_reset, av_config:reset, irq_synchronizer:receiver_reset, mm_interconnect_2:audio_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                                 : std_logic;                     -- rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, avalon_st_adapter_004:in_rst_0_reset, avalon_st_adapter_005:in_rst_0_reset, mm_interconnect_2:sdcard_interface_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                                 : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_2:header_mac_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal rst_controller_004_reset_out_reset                                 : std_logic;                     -- rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_2:nios2_reset_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in]
	signal rst_controller_005_reset_out_reset                                 : std_logic;                     -- rst_controller_005:reset_out -> sram_0:reset
	signal rst_controller_006_reset_out_reset                                 : std_logic;                     -- rst_controller_006:reset_out -> [irq_synchronizer_001:receiver_reset, mm_interconnect_2:textmode_controller_reset_reset_bridge_in_reset_reset, rst_controller_006_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0]
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_2_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_2_jtag_uart_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_2_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_2_textmode_controller_avalon_slave_write_ports_inv : std_logic;                     -- mm_interconnect_2_textmode_controller_avalon_slave_write:inv -> textmode_controller:write_n
	signal mm_interconnect_2_sdram_s1_read_ports_inv                          : std_logic;                     -- mm_interconnect_2_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_2_sdram_s1_byteenable_ports_inv                    : std_logic_vector(3 downto 0);  -- mm_interconnect_2_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_2_sdram_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_2_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_2_pio_0_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_2_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_002_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [fft_wrapper_header_0:reset_n, fir_l:res_n, fir_r:res_n, m2s_fifo_ffth:reset_n, m2s_fifo_fir_l:reset_n, m2s_fifo_fir_r:reset_n, pio_0:reset_n, s2m_fifo_ffth:reset_n, s2m_fifo_fir_l:reset_n, s2m_fifo_fir_r:reset_n, sdcard_interface:i_reset_n, sdram:reset_n, touch_cntrl:res_n]
	signal rst_controller_003_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> [header_mac_0:res_n, multiplexer_sram_0:res_n]
	signal rst_controller_004_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> [jtag_uart:rst_n, nios2:reset_n]
	signal rst_controller_006_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_006_reset_out_reset:inv -> textmode_controller:reset_n

begin

	altpll : component reverb_template_altpll
		port map (
			clk                => clk_clk,                                      --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,               -- inclk_interface_reset.reset
			read               => mm_interconnect_2_altpll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_2_altpll_pll_slave_write,     --                      .write
			address            => mm_interconnect_2_altpll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_2_altpll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_2_altpll_pll_slave_writedata, --                      .writedata
			c0                 => altpll_c0_clk,                                --                    c0.clk
			c1                 => clk_125_clk,                                  --                    c1.clk
			c2                 => altpll_c2_clk,                                --                    c2.clk
			c3                 => clk_2p5_clk,                                  --                    c3.clk
			scandone           => open,                                         --           (terminated)
			scandataout        => open,                                         --           (terminated)
			phasecounterselect => "0000",                                       --           (terminated)
			phaseupdown        => '0',                                          --           (terminated)
			phasestep          => '0',                                          --           (terminated)
			scanclk            => '0',                                          --           (terminated)
			scanclkena         => '0',                                          --           (terminated)
			scandata           => '0',                                          --           (terminated)
			configupdate       => '0',                                          --           (terminated)
			areset             => '0',                                          --           (terminated)
			locked             => open,                                         --           (terminated)
			phasedone          => open                                          --           (terminated)
		);

	altpll_sram : component reverb_template_altpll_sram
		port map (
			clk                => clk_clk,                                           --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                    -- inclk_interface_reset.reset
			read               => mm_interconnect_2_altpll_sram_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_2_altpll_sram_pll_slave_write,     --                      .write
			address            => mm_interconnect_2_altpll_sram_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_2_altpll_sram_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_2_altpll_sram_pll_slave_writedata, --                      .writedata
			c0                 => altpll_sram_c0_clk,                                --                    c0.clk
			scandone           => open,                                              --           (terminated)
			scandataout        => open,                                              --           (terminated)
			areset             => '0',                                               --           (terminated)
			locked             => open,                                              --           (terminated)
			phasedone          => open,                                              --           (terminated)
			phasecounterselect => "0000",                                            --           (terminated)
			phaseupdown        => '0',                                               --           (terminated)
			phasestep          => '0',                                               --           (terminated)
			scanclk            => '0',                                               --           (terminated)
			scanclkena         => '0',                                               --           (terminated)
			scandata           => '0',                                               --           (terminated)
			configupdate       => '0'                                                --           (terminated)
		);

	audio : component reverb_template_audio
		port map (
			clk         => clk_clk,                                               --                clk.clk
			reset       => rst_controller_001_reset_out_reset,                    --              reset.reset
			address     => mm_interconnect_2_audio_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_2_audio_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_2_audio_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_2_audio_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_2_audio_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_2_audio_avalon_audio_slave_readdata,   --                   .readdata
			irq         => irq_synchronizer_receiver_irq(0),                      --          interrupt.irq
			AUD_ADCDAT  => audio_ADCDAT,                                          -- external_interface.export
			AUD_ADCLRCK => audio_ADCLRCK,                                         --                   .export
			AUD_BCLK    => audio_BCLK,                                            --                   .export
			AUD_DACDAT  => audio_DACDAT,                                          --                   .export
			AUD_DACLRCK => audio_DACLRCK                                          --                   .export
		);

	audio_pll : component reverb_template_audio_pll
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			audio_clk_clk      => audio_clk_clk,                      --    audio_clk.clk
			reset_source_reset => open                                -- reset_source.reset
		);

	av_config : component reverb_template_av_config
		port map (
			clk         => clk_clk,                                                        --                    clk.clk
			reset       => rst_controller_001_reset_out_reset,                             --                  reset.reset
			address     => mm_interconnect_2_av_config_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_2_av_config_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_2_av_config_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_2_av_config_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_2_av_config_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_2_av_config_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_config_SDAT,                                              --     external_interface.export
			I2C_SCLK    => audio_config_SCLK                                               --                       .export
		);

	fft_wrapper_header_0 : component fft_wrapper_header
		port map (
			clk         => altpll_c0_clk,                                      --                   clock.clk
			reset_n     => rst_controller_002_reset_out_reset_ports_inv,       --                   reset.reset_n
			stin_data   => avalon_st_adapter_003_out_0_data,                   --   avalon_streaming_sink.data
			stin_valid  => avalon_st_adapter_003_out_0_valid,                  --                        .valid
			stin_ready  => avalon_st_adapter_003_out_0_ready,                  --                        .ready
			stout_data  => fft_wrapper_header_0_avalon_streaming_source_data,  -- avalon_streaming_source.data
			stout_ready => fft_wrapper_header_0_avalon_streaming_source_ready, --                        .ready
			stout_valid => fft_wrapper_header_0_avalon_streaming_source_valid, --                        .valid
			inverse     => pio_0_external_connection_export                    --                 inverse.export
		);

	fir_l : component fir
		generic map (
			NUM_COEFFICIENTS => 512,
			DATA_WIDTH       => 32,
			ADDR_WIDTH       => 9
		)
		port map (
			clk          => altpll_c0_clk,                                    --                   clock.clk
			stin_data    => avalon_st_adapter_004_out_0_data,                 --   avalon_streaming_sink.data
			stin_valid   => avalon_st_adapter_004_out_0_valid,                --                        .valid
			stin_ready   => avalon_st_adapter_004_out_0_ready,                --                        .ready
			res_n        => rst_controller_002_reset_out_reset_ports_inv,     --              reset_sink.reset_n
			mm_address   => mm_interconnect_2_fir_l_avalon_slave_0_address,   --          avalon_slave_0.address
			mm_write     => mm_interconnect_2_fir_l_avalon_slave_0_write,     --                        .write
			mm_read      => mm_interconnect_2_fir_l_avalon_slave_0_read,      --                        .read
			mm_writedata => mm_interconnect_2_fir_l_avalon_slave_0_writedata, --                        .writedata
			mm_readdata  => mm_interconnect_2_fir_l_avalon_slave_0_readdata,  --                        .readdata
			stout_data   => fir_l_avalon_streaming_source_data,               -- avalon_streaming_source.data
			stout_ready  => fir_l_avalon_streaming_source_ready,              --                        .ready
			stout_valid  => fir_l_avalon_streaming_source_valid               --                        .valid
		);

	fir_r : component fir
		generic map (
			NUM_COEFFICIENTS => 512,
			DATA_WIDTH       => 32,
			ADDR_WIDTH       => 9
		)
		port map (
			clk          => altpll_c0_clk,                                    --                   clock.clk
			stin_data    => avalon_st_adapter_005_out_0_data,                 --   avalon_streaming_sink.data
			stin_valid   => avalon_st_adapter_005_out_0_valid,                --                        .valid
			stin_ready   => avalon_st_adapter_005_out_0_ready,                --                        .ready
			res_n        => rst_controller_002_reset_out_reset_ports_inv,     --              reset_sink.reset_n
			mm_address   => mm_interconnect_2_fir_r_avalon_slave_0_address,   --          avalon_slave_0.address
			mm_write     => mm_interconnect_2_fir_r_avalon_slave_0_write,     --                        .write
			mm_read      => mm_interconnect_2_fir_r_avalon_slave_0_read,      --                        .read
			mm_writedata => mm_interconnect_2_fir_r_avalon_slave_0_writedata, --                        .writedata
			mm_readdata  => mm_interconnect_2_fir_r_avalon_slave_0_readdata,  --                        .readdata
			stout_data   => fir_r_avalon_streaming_source_data,               -- avalon_streaming_source.data
			stout_ready  => fir_r_avalon_streaming_source_ready,              --                        .ready
			stout_valid  => fir_r_avalon_streaming_source_valid               --                        .valid
		);

	header_mac_0 : component mac_sram
		port map (
			clk             => altpll_sram_c0_clk,                                    --         clock.clk
			res_n           => rst_controller_003_reset_out_reset_ports_inv,          --    reset_sink.reset_n
			m_address       => header_mac_0_avalon_master_address,                    -- avalon_master.address
			m_write         => header_mac_0_avalon_master_write,                      --              .write
			m_read          => header_mac_0_avalon_master_read,                       --              .read
			m_writedata     => header_mac_0_avalon_master_writedata,                  --              .writedata
			m_readdata      => header_mac_0_avalon_master_readdata,                   --              .readdata
			m_readdatavalid => header_mac_0_avalon_master_readdatavalid,              --              .readdatavalid
			s_address       => mm_interconnect_2_header_mac_0_avalon_slave_address,   --  avalon_slave.address
			s_write         => mm_interconnect_2_header_mac_0_avalon_slave_write,     --              .write
			s_read          => mm_interconnect_2_header_mac_0_avalon_slave_read,      --              .read
			s_writedata     => mm_interconnect_2_header_mac_0_avalon_slave_writedata, --              .writedata
			s_readdata      => mm_interconnect_2_header_mac_0_avalon_slave_readdata,  --              .readdata
			sel             => header_mac_0_sel_export                                --           sel.export
		);

	jtag_uart : component reverb_template_jtag_uart
		port map (
			clk            => altpll_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_004_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_2_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_2_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_2_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                       --               irq.irq
		);

	m2s_fifo_ffth : component reverb_template_m2s_fifo_ffth
		port map (
			wrclock                          => altpll_c0_clk,                                  --   clk_in.clk
			reset_n                          => rst_controller_002_reset_out_reset_ports_inv,   -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_2_m2s_fifo_ffth_in_writedata,   --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_2_m2s_fifo_ffth_in_write,       --         .write
			avalonmm_write_slave_address     => mm_interconnect_2_m2s_fifo_ffth_in_address(0),  --         .address
			avalonmm_write_slave_waitrequest => mm_interconnect_2_m2s_fifo_ffth_in_waitrequest, --         .waitrequest
			avalonst_source_valid            => m2s_fifo_ffth_out_valid,                        --      out.valid
			avalonst_source_data             => m2s_fifo_ffth_out_data,                         --         .data
			avalonst_source_ready            => m2s_fifo_ffth_out_ready                         --         .ready
		);

	m2s_fifo_fir_l : component reverb_template_m2s_fifo_fir_l
		port map (
			wrclock                          => altpll_c0_clk,                                   --   clk_in.clk
			reset_n                          => rst_controller_002_reset_out_reset_ports_inv,    -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_2_m2s_fifo_fir_l_in_writedata,   --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_2_m2s_fifo_fir_l_in_write,       --         .write
			avalonmm_write_slave_address     => mm_interconnect_2_m2s_fifo_fir_l_in_address(0),  --         .address
			avalonmm_write_slave_waitrequest => mm_interconnect_2_m2s_fifo_fir_l_in_waitrequest, --         .waitrequest
			avalonst_source_valid            => m2s_fifo_fir_l_out_valid,                        --      out.valid
			avalonst_source_data             => m2s_fifo_fir_l_out_data,                         --         .data
			avalonst_source_ready            => m2s_fifo_fir_l_out_ready                         --         .ready
		);

	m2s_fifo_fir_r : component reverb_template_m2s_fifo_fir_l
		port map (
			wrclock                          => altpll_c0_clk,                                   --   clk_in.clk
			reset_n                          => rst_controller_002_reset_out_reset_ports_inv,    -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_2_m2s_fifo_fir_r_in_writedata,   --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_2_m2s_fifo_fir_r_in_write,       --         .write
			avalonmm_write_slave_address     => mm_interconnect_2_m2s_fifo_fir_r_in_address(0),  --         .address
			avalonmm_write_slave_waitrequest => mm_interconnect_2_m2s_fifo_fir_r_in_waitrequest, --         .waitrequest
			avalonst_source_valid            => m2s_fifo_fir_r_out_valid,                        --      out.valid
			avalonst_source_data             => m2s_fifo_fir_r_out_data,                         --         .data
			avalonst_source_ready            => m2s_fifo_fir_r_out_ready                         --         .ready
		);

	multiplexer_sram_0 : component multiplexer
		port map (
			clk              => altpll_sram_c0_clk,                                    --         clock.clk
			s0_address       => header_mac_0_avalon_master_address,                    --            s0.address
			s0_write         => header_mac_0_avalon_master_write,                      --              .write
			s0_writedata     => header_mac_0_avalon_master_writedata,                  --              .writedata
			s0_read          => header_mac_0_avalon_master_read,                       --              .read
			s0_readdata      => header_mac_0_avalon_master_readdata,                   --              .readdata
			s0_readdatavalid => header_mac_0_avalon_master_readdatavalid,              --              .readdatavalid
			s1_address       => mm_interconnect_2_multiplexer_sram_0_s1_address,       --            s1.address
			s1_write         => mm_interconnect_2_multiplexer_sram_0_s1_write,         --              .write
			s1_writedata     => mm_interconnect_2_multiplexer_sram_0_s1_writedata,     --              .writedata
			s1_read          => mm_interconnect_2_multiplexer_sram_0_s1_read,          --              .read
			s1_readdata      => mm_interconnect_2_multiplexer_sram_0_s1_readdata,      --              .readdata
			s1_readdatavalid => mm_interconnect_2_multiplexer_sram_0_s1_readdatavalid, --              .readdatavalid
			s1_byteanable    => mm_interconnect_2_multiplexer_sram_0_s1_byteenable,    --              .byteenable
			m_address        => multiplexer_sram_0_avalon_master_address,              -- avalon_master.address
			m_byteanable     => multiplexer_sram_0_avalon_master_byteenable,           --              .byteenable
			m_write          => multiplexer_sram_0_avalon_master_write,                --              .write
			m_writedata      => multiplexer_sram_0_avalon_master_writedata,            --              .writedata
			m_read           => multiplexer_sram_0_avalon_master_read,                 --              .read
			m_readdata       => multiplexer_sram_0_avalon_master_readdata,             --              .readdata
			m_readdatavalid  => multiplexer_sram_0_avalon_master_readdatavalid,        --              .readdatavalid
			res_n            => rst_controller_003_reset_out_reset_ports_inv,          --    reset_sink.reset_n
			sel              => header_mac_0_sel_export                                --           sel.export
		);

	nios2 : component reverb_template_nios2
		port map (
			clk                                 => altpll_c0_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_004_reset_out_reset_ports_inv,        --                     reset.reset_n
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_2_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_2_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_2_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_2_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_2_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_2_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_2_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_2_nios2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	pio_0 : component reverb_template_pio_0
		port map (
			clk        => altpll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_0_s1_address,           --                  s1.address
			write_n    => mm_interconnect_2_pio_0_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_2_pio_0_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_2_pio_0_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_2_pio_0_s1_readdata,          --                    .readdata
			out_port   => pio_0_external_connection_export              -- external_connection.export
		);

	s2m_fifo_ffth : component reverb_template_s2m_fifo_ffth
		port map (
			wrclock                         => altpll_c0_clk,                                   --   clk_in.clk
			reset_n                         => rst_controller_002_reset_out_reset_ports_inv,    -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_out_0_valid,                   --       in.valid
			avalonst_sink_data              => avalon_st_adapter_out_0_data,                    --         .data
			avalonst_sink_ready             => avalon_st_adapter_out_0_ready,                   --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_2_s2m_fifo_ffth_out_readdata,    --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_2_s2m_fifo_ffth_out_read,        --         .read
			avalonmm_read_slave_address     => mm_interconnect_2_s2m_fifo_ffth_out_address(0),  --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_2_s2m_fifo_ffth_out_waitrequest  --         .waitrequest
		);

	s2m_fifo_fir_l : component reverb_template_s2m_fifo_fir_l
		port map (
			wrclock                         => altpll_c0_clk,                                    --   clk_in.clk
			reset_n                         => rst_controller_002_reset_out_reset_ports_inv,     -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_001_out_0_valid,                --       in.valid
			avalonst_sink_data              => avalon_st_adapter_001_out_0_data,                 --         .data
			avalonst_sink_ready             => avalon_st_adapter_001_out_0_ready,                --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_2_s2m_fifo_fir_l_out_readdata,    --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_2_s2m_fifo_fir_l_out_read,        --         .read
			avalonmm_read_slave_address     => mm_interconnect_2_s2m_fifo_fir_l_out_address(0),  --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_2_s2m_fifo_fir_l_out_waitrequest  --         .waitrequest
		);

	s2m_fifo_fir_r : component reverb_template_s2m_fifo_fir_l
		port map (
			wrclock                         => altpll_c0_clk,                                    --   clk_in.clk
			reset_n                         => rst_controller_002_reset_out_reset_ports_inv,     -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_002_out_0_valid,                --       in.valid
			avalonst_sink_data              => avalon_st_adapter_002_out_0_data,                 --         .data
			avalonst_sink_ready             => avalon_st_adapter_002_out_0_ready,                --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_2_s2m_fifo_fir_r_out_readdata,    --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_2_s2m_fifo_fir_r_out_read,        --         .read
			avalonmm_read_slave_address     => mm_interconnect_2_s2m_fifo_fir_r_out_address(0),  --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_2_s2m_fifo_fir_r_out_waitrequest  --         .waitrequest
		);

	sdcard_interface : component Altera_UP_SD_Card_Avalon_Interface
		port map (
			i_avalon_chip_select => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_chipselect,  -- avalon_sdcard_slave.chipselect
			i_avalon_address     => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_address,     --                    .address
			i_avalon_read        => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_read,        --                    .read
			i_avalon_write       => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_write,       --                    .write
			i_avalon_byteenable  => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_byteenable,  --                    .byteenable
			i_avalon_writedata   => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_writedata,   --                    .writedata
			o_avalon_readdata    => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_readdata,    --                    .readdata
			o_avalon_waitrequest => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_waitrequest, --                    .waitrequest
			i_clock              => altpll_c0_clk,                                                      --                 clk.clk
			i_reset_n            => rst_controller_002_reset_out_reset_ports_inv,                       --               reset.reset_n
			b_SD_cmd             => sdcard_b_SD_cmd,                                                    --         conduit_end.export
			b_SD_dat             => sdcard_b_SD_dat,                                                    --                    .export
			b_SD_dat3            => sdcard_b_SD_dat3,                                                   --                    .export
			o_SD_clock           => sdcard_o_SD_clock                                                   --                    .export
		);

	sdram : component reverb_template_sdram
		port map (
			clk            => altpll_c0_clk,                                   --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_2_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_2_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_2_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_2_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_2_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_2_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_2_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_2_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_2_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sram_0 : component reverb_template_sram_0
		port map (
			clk           => altpll_sram_c0_clk,                             --                clk.clk
			reset         => rst_controller_005_reset_out_reset,             --              reset.reset
			SRAM_DQ       => sram_DQ,                                        -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                      --                   .export
			SRAM_LB_N     => sram_LB_N,                                      --                   .export
			SRAM_UB_N     => sram_UB_N,                                      --                   .export
			SRAM_CE_N     => sram_CE_N,                                      --                   .export
			SRAM_OE_N     => sram_OE_N,                                      --                   .export
			SRAM_WE_N     => sram_WE_N,                                      --                   .export
			address       => multiplexer_sram_0_avalon_master_address,       --  avalon_sram_slave.address
			byteenable    => multiplexer_sram_0_avalon_master_byteenable,    --                   .byteenable
			read          => multiplexer_sram_0_avalon_master_read,          --                   .read
			write         => multiplexer_sram_0_avalon_master_write,         --                   .write
			writedata     => multiplexer_sram_0_avalon_master_writedata,     --                   .writedata
			readdata      => multiplexer_sram_0_avalon_master_readdata,      --                   .readdata
			readdatavalid => multiplexer_sram_0_avalon_master_readdatavalid  --                   .readdatavalid
		);

	textmode_controller : component textmode_controller_avalon
		generic map (
			ROW_COUNT    => 30,
			COLUMN_COUNT => 100,
			CLK_FREQ     => 25000000
		)
		port map (
			clk       => altpll_c2_clk,                                                      --        clock.clk
			reset_n   => rst_controller_006_reset_out_reset_ports_inv,                       --        reset.reset_n
			address   => mm_interconnect_2_textmode_controller_avalon_slave_address,         -- avalon_slave.address
			write_n   => mm_interconnect_2_textmode_controller_avalon_slave_write_ports_inv, --             .write_n
			writedata => mm_interconnect_2_textmode_controller_avalon_slave_writedata,       --             .writedata
			readdata  => mm_interconnect_2_textmode_controller_avalon_slave_readdata,        --             .readdata
			b         => textmode_b,                                                         --     conduits.b
			den       => textmode_den,                                                       --             .den
			g         => textmode_g,                                                         --             .g
			hd        => textmode_hd,                                                        --             .hd
			r         => textmode_r,                                                         --             .r
			vd        => textmode_vd,                                                        --             .vd
			grest     => textmode_grest,                                                     --             .grest
			irq       => irq_synchronizer_001_receiver_irq(0)                                --    interrupt.irq
		);

	touch_cntrl : component avalon_touch_cntrl
		generic map (
			SYS_CLK => 100000000
		)
		port map (
			clk          => altpll_c0_clk,                                        --        clock.clk
			adc_cs       => touch_cntrl_ext_adc_cs,                               --          ext.adc_cs
			adc_dclk     => touch_cntrl_ext_adc_dclk,                             --             .adc_dclk
			adc_din      => touch_cntrl_ext_adc_din,                              --             .adc_din
			adc_dout     => touch_cntrl_ext_adc_dout,                             --             .adc_dout
			adc_penirq_n => touch_cntrl_ext_adc_penirq_n,                         --             .adc_penirq_n
			irq          => irq_mapper_receiver3_irq,                             --          irq.irq
			address      => mm_interconnect_2_touch_cntrl_avalon_slave_address,   -- avalon_slave.address
			write        => mm_interconnect_2_touch_cntrl_avalon_slave_write,     --             .write
			read         => mm_interconnect_2_touch_cntrl_avalon_slave_read,      --             .read
			writedata    => mm_interconnect_2_touch_cntrl_avalon_slave_writedata, --             .writedata
			readdata     => mm_interconnect_2_touch_cntrl_avalon_slave_readdata,  --             .readdata
			res_n        => rst_controller_002_reset_out_reset_ports_inv          --        reset.reset_n
		);

	mm_interconnect_2 : component reverb_template_mm_interconnect_2
		port map (
			altpll_c0_clk                                            => altpll_c0_clk,                                                      --                                          altpll_c0.clk
			altpll_c2_clk                                            => altpll_c2_clk,                                                      --                                          altpll_c2.clk
			altpll_sram_c0_clk                                       => altpll_sram_c0_clk,                                                 --                                     altpll_sram_c0.clk
			sys_clk_clk_clk                                          => clk_clk,                                                            --                                        sys_clk_clk.clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                     -- altpll_inclk_interface_reset_reset_bridge_in_reset.reset
			audio_reset_reset_bridge_in_reset_reset                  => rst_controller_001_reset_out_reset,                                 --                  audio_reset_reset_bridge_in_reset.reset
			header_mac_0_reset_sink_reset_bridge_in_reset_reset      => rst_controller_003_reset_out_reset,                                 --      header_mac_0_reset_sink_reset_bridge_in_reset.reset
			nios2_reset_reset_bridge_in_reset_reset                  => rst_controller_004_reset_out_reset,                                 --                  nios2_reset_reset_bridge_in_reset.reset
			sdcard_interface_reset_reset_bridge_in_reset_reset       => rst_controller_002_reset_out_reset,                                 --       sdcard_interface_reset_reset_bridge_in_reset.reset
			textmode_controller_reset_reset_bridge_in_reset_reset    => rst_controller_006_reset_out_reset,                                 --    textmode_controller_reset_reset_bridge_in_reset.reset
			nios2_data_master_address                                => nios2_data_master_address,                                          --                                  nios2_data_master.address
			nios2_data_master_waitrequest                            => nios2_data_master_waitrequest,                                      --                                                   .waitrequest
			nios2_data_master_byteenable                             => nios2_data_master_byteenable,                                       --                                                   .byteenable
			nios2_data_master_read                                   => nios2_data_master_read,                                             --                                                   .read
			nios2_data_master_readdata                               => nios2_data_master_readdata,                                         --                                                   .readdata
			nios2_data_master_readdatavalid                          => nios2_data_master_readdatavalid,                                    --                                                   .readdatavalid
			nios2_data_master_write                                  => nios2_data_master_write,                                            --                                                   .write
			nios2_data_master_writedata                              => nios2_data_master_writedata,                                        --                                                   .writedata
			nios2_data_master_debugaccess                            => nios2_data_master_debugaccess,                                      --                                                   .debugaccess
			nios2_instruction_master_address                         => nios2_instruction_master_address,                                   --                           nios2_instruction_master.address
			nios2_instruction_master_waitrequest                     => nios2_instruction_master_waitrequest,                               --                                                   .waitrequest
			nios2_instruction_master_read                            => nios2_instruction_master_read,                                      --                                                   .read
			nios2_instruction_master_readdata                        => nios2_instruction_master_readdata,                                  --                                                   .readdata
			nios2_instruction_master_readdatavalid                   => nios2_instruction_master_readdatavalid,                             --                                                   .readdatavalid
			altpll_pll_slave_address                                 => mm_interconnect_2_altpll_pll_slave_address,                         --                                   altpll_pll_slave.address
			altpll_pll_slave_write                                   => mm_interconnect_2_altpll_pll_slave_write,                           --                                                   .write
			altpll_pll_slave_read                                    => mm_interconnect_2_altpll_pll_slave_read,                            --                                                   .read
			altpll_pll_slave_readdata                                => mm_interconnect_2_altpll_pll_slave_readdata,                        --                                                   .readdata
			altpll_pll_slave_writedata                               => mm_interconnect_2_altpll_pll_slave_writedata,                       --                                                   .writedata
			altpll_sram_pll_slave_address                            => mm_interconnect_2_altpll_sram_pll_slave_address,                    --                              altpll_sram_pll_slave.address
			altpll_sram_pll_slave_write                              => mm_interconnect_2_altpll_sram_pll_slave_write,                      --                                                   .write
			altpll_sram_pll_slave_read                               => mm_interconnect_2_altpll_sram_pll_slave_read,                       --                                                   .read
			altpll_sram_pll_slave_readdata                           => mm_interconnect_2_altpll_sram_pll_slave_readdata,                   --                                                   .readdata
			altpll_sram_pll_slave_writedata                          => mm_interconnect_2_altpll_sram_pll_slave_writedata,                  --                                                   .writedata
			audio_avalon_audio_slave_address                         => mm_interconnect_2_audio_avalon_audio_slave_address,                 --                           audio_avalon_audio_slave.address
			audio_avalon_audio_slave_write                           => mm_interconnect_2_audio_avalon_audio_slave_write,                   --                                                   .write
			audio_avalon_audio_slave_read                            => mm_interconnect_2_audio_avalon_audio_slave_read,                    --                                                   .read
			audio_avalon_audio_slave_readdata                        => mm_interconnect_2_audio_avalon_audio_slave_readdata,                --                                                   .readdata
			audio_avalon_audio_slave_writedata                       => mm_interconnect_2_audio_avalon_audio_slave_writedata,               --                                                   .writedata
			audio_avalon_audio_slave_chipselect                      => mm_interconnect_2_audio_avalon_audio_slave_chipselect,              --                                                   .chipselect
			av_config_avalon_av_config_slave_address                 => mm_interconnect_2_av_config_avalon_av_config_slave_address,         --                   av_config_avalon_av_config_slave.address
			av_config_avalon_av_config_slave_write                   => mm_interconnect_2_av_config_avalon_av_config_slave_write,           --                                                   .write
			av_config_avalon_av_config_slave_read                    => mm_interconnect_2_av_config_avalon_av_config_slave_read,            --                                                   .read
			av_config_avalon_av_config_slave_readdata                => mm_interconnect_2_av_config_avalon_av_config_slave_readdata,        --                                                   .readdata
			av_config_avalon_av_config_slave_writedata               => mm_interconnect_2_av_config_avalon_av_config_slave_writedata,       --                                                   .writedata
			av_config_avalon_av_config_slave_byteenable              => mm_interconnect_2_av_config_avalon_av_config_slave_byteenable,      --                                                   .byteenable
			av_config_avalon_av_config_slave_waitrequest             => mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest,     --                                                   .waitrequest
			fir_l_avalon_slave_0_address                             => mm_interconnect_2_fir_l_avalon_slave_0_address,                     --                               fir_l_avalon_slave_0.address
			fir_l_avalon_slave_0_write                               => mm_interconnect_2_fir_l_avalon_slave_0_write,                       --                                                   .write
			fir_l_avalon_slave_0_read                                => mm_interconnect_2_fir_l_avalon_slave_0_read,                        --                                                   .read
			fir_l_avalon_slave_0_readdata                            => mm_interconnect_2_fir_l_avalon_slave_0_readdata,                    --                                                   .readdata
			fir_l_avalon_slave_0_writedata                           => mm_interconnect_2_fir_l_avalon_slave_0_writedata,                   --                                                   .writedata
			fir_r_avalon_slave_0_address                             => mm_interconnect_2_fir_r_avalon_slave_0_address,                     --                               fir_r_avalon_slave_0.address
			fir_r_avalon_slave_0_write                               => mm_interconnect_2_fir_r_avalon_slave_0_write,                       --                                                   .write
			fir_r_avalon_slave_0_read                                => mm_interconnect_2_fir_r_avalon_slave_0_read,                        --                                                   .read
			fir_r_avalon_slave_0_readdata                            => mm_interconnect_2_fir_r_avalon_slave_0_readdata,                    --                                                   .readdata
			fir_r_avalon_slave_0_writedata                           => mm_interconnect_2_fir_r_avalon_slave_0_writedata,                   --                                                   .writedata
			header_mac_0_avalon_slave_address                        => mm_interconnect_2_header_mac_0_avalon_slave_address,                --                          header_mac_0_avalon_slave.address
			header_mac_0_avalon_slave_write                          => mm_interconnect_2_header_mac_0_avalon_slave_write,                  --                                                   .write
			header_mac_0_avalon_slave_read                           => mm_interconnect_2_header_mac_0_avalon_slave_read,                   --                                                   .read
			header_mac_0_avalon_slave_readdata                       => mm_interconnect_2_header_mac_0_avalon_slave_readdata,               --                                                   .readdata
			header_mac_0_avalon_slave_writedata                      => mm_interconnect_2_header_mac_0_avalon_slave_writedata,              --                                                   .writedata
			jtag_uart_avalon_jtag_slave_address                      => mm_interconnect_2_jtag_uart_avalon_jtag_slave_address,              --                        jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                        => mm_interconnect_2_jtag_uart_avalon_jtag_slave_write,                --                                                   .write
			jtag_uart_avalon_jtag_slave_read                         => mm_interconnect_2_jtag_uart_avalon_jtag_slave_read,                 --                                                   .read
			jtag_uart_avalon_jtag_slave_readdata                     => mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata,             --                                                   .readdata
			jtag_uart_avalon_jtag_slave_writedata                    => mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata,            --                                                   .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                  => mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest,          --                                                   .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                   => mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect,           --                                                   .chipselect
			m2s_fifo_ffth_in_address                                 => mm_interconnect_2_m2s_fifo_ffth_in_address,                         --                                   m2s_fifo_ffth_in.address
			m2s_fifo_ffth_in_write                                   => mm_interconnect_2_m2s_fifo_ffth_in_write,                           --                                                   .write
			m2s_fifo_ffth_in_writedata                               => mm_interconnect_2_m2s_fifo_ffth_in_writedata,                       --                                                   .writedata
			m2s_fifo_ffth_in_waitrequest                             => mm_interconnect_2_m2s_fifo_ffth_in_waitrequest,                     --                                                   .waitrequest
			m2s_fifo_fir_l_in_address                                => mm_interconnect_2_m2s_fifo_fir_l_in_address,                        --                                  m2s_fifo_fir_l_in.address
			m2s_fifo_fir_l_in_write                                  => mm_interconnect_2_m2s_fifo_fir_l_in_write,                          --                                                   .write
			m2s_fifo_fir_l_in_writedata                              => mm_interconnect_2_m2s_fifo_fir_l_in_writedata,                      --                                                   .writedata
			m2s_fifo_fir_l_in_waitrequest                            => mm_interconnect_2_m2s_fifo_fir_l_in_waitrequest,                    --                                                   .waitrequest
			m2s_fifo_fir_r_in_address                                => mm_interconnect_2_m2s_fifo_fir_r_in_address,                        --                                  m2s_fifo_fir_r_in.address
			m2s_fifo_fir_r_in_write                                  => mm_interconnect_2_m2s_fifo_fir_r_in_write,                          --                                                   .write
			m2s_fifo_fir_r_in_writedata                              => mm_interconnect_2_m2s_fifo_fir_r_in_writedata,                      --                                                   .writedata
			m2s_fifo_fir_r_in_waitrequest                            => mm_interconnect_2_m2s_fifo_fir_r_in_waitrequest,                    --                                                   .waitrequest
			multiplexer_sram_0_s1_address                            => mm_interconnect_2_multiplexer_sram_0_s1_address,                    --                              multiplexer_sram_0_s1.address
			multiplexer_sram_0_s1_write                              => mm_interconnect_2_multiplexer_sram_0_s1_write,                      --                                                   .write
			multiplexer_sram_0_s1_read                               => mm_interconnect_2_multiplexer_sram_0_s1_read,                       --                                                   .read
			multiplexer_sram_0_s1_readdata                           => mm_interconnect_2_multiplexer_sram_0_s1_readdata,                   --                                                   .readdata
			multiplexer_sram_0_s1_writedata                          => mm_interconnect_2_multiplexer_sram_0_s1_writedata,                  --                                                   .writedata
			multiplexer_sram_0_s1_byteenable                         => mm_interconnect_2_multiplexer_sram_0_s1_byteenable,                 --                                                   .byteenable
			multiplexer_sram_0_s1_readdatavalid                      => mm_interconnect_2_multiplexer_sram_0_s1_readdatavalid,              --                                                   .readdatavalid
			nios2_debug_mem_slave_address                            => mm_interconnect_2_nios2_debug_mem_slave_address,                    --                              nios2_debug_mem_slave.address
			nios2_debug_mem_slave_write                              => mm_interconnect_2_nios2_debug_mem_slave_write,                      --                                                   .write
			nios2_debug_mem_slave_read                               => mm_interconnect_2_nios2_debug_mem_slave_read,                       --                                                   .read
			nios2_debug_mem_slave_readdata                           => mm_interconnect_2_nios2_debug_mem_slave_readdata,                   --                                                   .readdata
			nios2_debug_mem_slave_writedata                          => mm_interconnect_2_nios2_debug_mem_slave_writedata,                  --                                                   .writedata
			nios2_debug_mem_slave_byteenable                         => mm_interconnect_2_nios2_debug_mem_slave_byteenable,                 --                                                   .byteenable
			nios2_debug_mem_slave_waitrequest                        => mm_interconnect_2_nios2_debug_mem_slave_waitrequest,                --                                                   .waitrequest
			nios2_debug_mem_slave_debugaccess                        => mm_interconnect_2_nios2_debug_mem_slave_debugaccess,                --                                                   .debugaccess
			pio_0_s1_address                                         => mm_interconnect_2_pio_0_s1_address,                                 --                                           pio_0_s1.address
			pio_0_s1_write                                           => mm_interconnect_2_pio_0_s1_write,                                   --                                                   .write
			pio_0_s1_readdata                                        => mm_interconnect_2_pio_0_s1_readdata,                                --                                                   .readdata
			pio_0_s1_writedata                                       => mm_interconnect_2_pio_0_s1_writedata,                               --                                                   .writedata
			pio_0_s1_chipselect                                      => mm_interconnect_2_pio_0_s1_chipselect,                              --                                                   .chipselect
			s2m_fifo_ffth_out_address                                => mm_interconnect_2_s2m_fifo_ffth_out_address,                        --                                  s2m_fifo_ffth_out.address
			s2m_fifo_ffth_out_read                                   => mm_interconnect_2_s2m_fifo_ffth_out_read,                           --                                                   .read
			s2m_fifo_ffth_out_readdata                               => mm_interconnect_2_s2m_fifo_ffth_out_readdata,                       --                                                   .readdata
			s2m_fifo_ffth_out_waitrequest                            => mm_interconnect_2_s2m_fifo_ffth_out_waitrequest,                    --                                                   .waitrequest
			s2m_fifo_fir_l_out_address                               => mm_interconnect_2_s2m_fifo_fir_l_out_address,                       --                                 s2m_fifo_fir_l_out.address
			s2m_fifo_fir_l_out_read                                  => mm_interconnect_2_s2m_fifo_fir_l_out_read,                          --                                                   .read
			s2m_fifo_fir_l_out_readdata                              => mm_interconnect_2_s2m_fifo_fir_l_out_readdata,                      --                                                   .readdata
			s2m_fifo_fir_l_out_waitrequest                           => mm_interconnect_2_s2m_fifo_fir_l_out_waitrequest,                   --                                                   .waitrequest
			s2m_fifo_fir_r_out_address                               => mm_interconnect_2_s2m_fifo_fir_r_out_address,                       --                                 s2m_fifo_fir_r_out.address
			s2m_fifo_fir_r_out_read                                  => mm_interconnect_2_s2m_fifo_fir_r_out_read,                          --                                                   .read
			s2m_fifo_fir_r_out_readdata                              => mm_interconnect_2_s2m_fifo_fir_r_out_readdata,                      --                                                   .readdata
			s2m_fifo_fir_r_out_waitrequest                           => mm_interconnect_2_s2m_fifo_fir_r_out_waitrequest,                   --                                                   .waitrequest
			sdcard_interface_avalon_sdcard_slave_address             => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_address,     --               sdcard_interface_avalon_sdcard_slave.address
			sdcard_interface_avalon_sdcard_slave_write               => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_write,       --                                                   .write
			sdcard_interface_avalon_sdcard_slave_read                => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_read,        --                                                   .read
			sdcard_interface_avalon_sdcard_slave_readdata            => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_readdata,    --                                                   .readdata
			sdcard_interface_avalon_sdcard_slave_writedata           => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_writedata,   --                                                   .writedata
			sdcard_interface_avalon_sdcard_slave_byteenable          => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_byteenable,  --                                                   .byteenable
			sdcard_interface_avalon_sdcard_slave_waitrequest         => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_waitrequest, --                                                   .waitrequest
			sdcard_interface_avalon_sdcard_slave_chipselect          => mm_interconnect_2_sdcard_interface_avalon_sdcard_slave_chipselect,  --                                                   .chipselect
			sdram_s1_address                                         => mm_interconnect_2_sdram_s1_address,                                 --                                           sdram_s1.address
			sdram_s1_write                                           => mm_interconnect_2_sdram_s1_write,                                   --                                                   .write
			sdram_s1_read                                            => mm_interconnect_2_sdram_s1_read,                                    --                                                   .read
			sdram_s1_readdata                                        => mm_interconnect_2_sdram_s1_readdata,                                --                                                   .readdata
			sdram_s1_writedata                                       => mm_interconnect_2_sdram_s1_writedata,                               --                                                   .writedata
			sdram_s1_byteenable                                      => mm_interconnect_2_sdram_s1_byteenable,                              --                                                   .byteenable
			sdram_s1_readdatavalid                                   => mm_interconnect_2_sdram_s1_readdatavalid,                           --                                                   .readdatavalid
			sdram_s1_waitrequest                                     => mm_interconnect_2_sdram_s1_waitrequest,                             --                                                   .waitrequest
			sdram_s1_chipselect                                      => mm_interconnect_2_sdram_s1_chipselect,                              --                                                   .chipselect
			textmode_controller_avalon_slave_address                 => mm_interconnect_2_textmode_controller_avalon_slave_address,         --                   textmode_controller_avalon_slave.address
			textmode_controller_avalon_slave_write                   => mm_interconnect_2_textmode_controller_avalon_slave_write,           --                                                   .write
			textmode_controller_avalon_slave_readdata                => mm_interconnect_2_textmode_controller_avalon_slave_readdata,        --                                                   .readdata
			textmode_controller_avalon_slave_writedata               => mm_interconnect_2_textmode_controller_avalon_slave_writedata,       --                                                   .writedata
			touch_cntrl_avalon_slave_address                         => mm_interconnect_2_touch_cntrl_avalon_slave_address,                 --                           touch_cntrl_avalon_slave.address
			touch_cntrl_avalon_slave_write                           => mm_interconnect_2_touch_cntrl_avalon_slave_write,                   --                                                   .write
			touch_cntrl_avalon_slave_read                            => mm_interconnect_2_touch_cntrl_avalon_slave_read,                    --                                                   .read
			touch_cntrl_avalon_slave_readdata                        => mm_interconnect_2_touch_cntrl_avalon_slave_readdata,                --                                                   .readdata
			touch_cntrl_avalon_slave_writedata                       => mm_interconnect_2_touch_cntrl_avalon_slave_writedata                --                                                   .writedata
		);

	irq_mapper : component reverb_template_irq_mapper
		port map (
			clk           => altpll_c0_clk,                      --       clk.clk
			reset         => rst_controller_004_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			sender_irq    => nios2_irq_irq                       --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => altpll_c0_clk,                      --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_004_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_c2_clk,                      --       receiver_clk.clk
			sender_clk     => altpll_c0_clk,                      --         sender_clk.clk
			receiver_reset => rst_controller_006_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_004_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	avalon_st_adapter : component reverb_template_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                                      -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset,                 -- in_rst_0.reset
			in_0_data      => fft_wrapper_header_0_avalon_streaming_source_data,  --     in_0.data
			in_0_valid     => fft_wrapper_header_0_avalon_streaming_source_valid, --         .valid
			in_0_ready     => fft_wrapper_header_0_avalon_streaming_source_ready, --         .ready
			out_0_data     => avalon_st_adapter_out_0_data,                       --    out_0.data
			out_0_valid    => avalon_st_adapter_out_0_valid,                      --         .valid
			out_0_ready    => avalon_st_adapter_out_0_ready                       --         .ready
		);

	avalon_st_adapter_001 : component reverb_template_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                       -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset,  -- in_rst_0.reset
			in_0_data      => fir_l_avalon_streaming_source_data,  --     in_0.data
			in_0_valid     => fir_l_avalon_streaming_source_valid, --         .valid
			in_0_ready     => fir_l_avalon_streaming_source_ready, --         .ready
			out_0_data     => avalon_st_adapter_001_out_0_data,    --    out_0.data
			out_0_valid    => avalon_st_adapter_001_out_0_valid,   --         .valid
			out_0_ready    => avalon_st_adapter_001_out_0_ready    --         .ready
		);

	avalon_st_adapter_002 : component reverb_template_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                       -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset,  -- in_rst_0.reset
			in_0_data      => fir_r_avalon_streaming_source_data,  --     in_0.data
			in_0_valid     => fir_r_avalon_streaming_source_valid, --         .valid
			in_0_ready     => fir_r_avalon_streaming_source_ready, --         .ready
			out_0_data     => avalon_st_adapter_002_out_0_data,    --    out_0.data
			out_0_valid    => avalon_st_adapter_002_out_0_valid,   --         .valid
			out_0_ready    => avalon_st_adapter_002_out_0_ready    --         .ready
		);

	avalon_st_adapter_003 : component reverb_template_avalon_st_adapter_003
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 1,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                      -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset, -- in_rst_0.reset
			in_0_data      => m2s_fifo_ffth_out_data,             --     in_0.data
			in_0_valid     => m2s_fifo_ffth_out_valid,            --         .valid
			in_0_ready     => m2s_fifo_ffth_out_ready,            --         .ready
			out_0_data     => avalon_st_adapter_003_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_003_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_003_out_0_ready   --         .ready
		);

	avalon_st_adapter_004 : component reverb_template_avalon_st_adapter_003
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 1,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                      -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset, -- in_rst_0.reset
			in_0_data      => m2s_fifo_fir_l_out_data,            --     in_0.data
			in_0_valid     => m2s_fifo_fir_l_out_valid,           --         .valid
			in_0_ready     => m2s_fifo_fir_l_out_ready,           --         .ready
			out_0_data     => avalon_st_adapter_004_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_004_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_004_out_0_ready   --         .ready
		);

	avalon_st_adapter_005 : component reverb_template_avalon_st_adapter_003
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 1,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => altpll_c0_clk,                      -- in_clk_0.clk
			in_rst_0_reset => rst_controller_002_reset_out_reset, -- in_rst_0.reset
			in_0_data      => m2s_fifo_fir_r_out_data,            --     in_0.data
			in_0_valid     => m2s_fifo_fir_r_out_valid,           --         .valid
			in_0_ready     => m2s_fifo_fir_r_out_ready,           --         .ready
			out_0_data     => avalon_st_adapter_005_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_005_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_005_out_0_ready   --         .ready
		);

	rst_controller : component reverb_template_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,         -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                            -- (terminated)
			reset_req_in0  => '0',                             -- (terminated)
			reset_req_in1  => '0',                             -- (terminated)
			reset_in2      => '0',                             -- (terminated)
			reset_req_in2  => '0',                             -- (terminated)
			reset_in3      => '0',                             -- (terminated)
			reset_req_in3  => '0',                             -- (terminated)
			reset_in4      => '0',                             -- (terminated)
			reset_req_in4  => '0',                             -- (terminated)
			reset_in5      => '0',                             -- (terminated)
			reset_req_in5  => '0',                             -- (terminated)
			reset_in6      => '0',                             -- (terminated)
			reset_req_in6  => '0',                             -- (terminated)
			reset_in7      => '0',                             -- (terminated)
			reset_req_in7  => '0',                             -- (terminated)
			reset_in8      => '0',                             -- (terminated)
			reset_req_in8  => '0',                             -- (terminated)
			reset_in9      => '0',                             -- (terminated)
			reset_req_in9  => '0',                             -- (terminated)
			reset_in10     => '0',                             -- (terminated)
			reset_req_in10 => '0',                             -- (terminated)
			reset_in11     => '0',                             -- (terminated)
			reset_req_in11 => '0',                             -- (terminated)
			reset_in12     => '0',                             -- (terminated)
			reset_req_in12 => '0',                             -- (terminated)
			reset_in13     => '0',                             -- (terminated)
			reset_req_in13 => '0',                             -- (terminated)
			reset_in14     => '0',                             -- (terminated)
			reset_req_in14 => '0',                             -- (terminated)
			reset_in15     => '0',                             -- (terminated)
			reset_req_in15 => '0'                              -- (terminated)
		);

	rst_controller_001 : component reverb_template_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component reverb_template_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_c0_clk,                      --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component reverb_template_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => altpll_sram_c0_clk,                 --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component reverb_template_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => altpll_c0_clk,                      --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_005 : component reverb_template_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_sram_c0_clk,                 --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_006 : component reverb_template_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_c2_clk,                      --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_2_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_2_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_2_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_2_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_2_textmode_controller_avalon_slave_write_ports_inv <= not mm_interconnect_2_textmode_controller_avalon_slave_write;

	mm_interconnect_2_sdram_s1_read_ports_inv <= not mm_interconnect_2_sdram_s1_read;

	mm_interconnect_2_sdram_s1_byteenable_ports_inv <= not mm_interconnect_2_sdram_s1_byteenable;

	mm_interconnect_2_sdram_s1_write_ports_inv <= not mm_interconnect_2_sdram_s1_write;

	mm_interconnect_2_pio_0_s1_write_ports_inv <= not mm_interconnect_2_pio_0_s1_write;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	rst_controller_006_reset_out_reset_ports_inv <= not rst_controller_006_reset_out_reset;

	sdram_clk_clk <= altpll_c0_clk;

	clk_25_clk <= altpll_c2_clk;

end architecture rtl; -- of reverb_template
