-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
C/Z2TeGf48OtnGsd5/8AXcZzQSg+Z6FO9SM1pyS0Mq63aAq4CRNQMlhpzc/exGTy
rPbN32pDW4APhMjemYNi/xzJkL0LGLpJctSMbujpwTLZ4cZV8odSBLQnu9VNcCqw
WpHpdpO55q96LOy7rqogJATTqG3etKlgRhaOw7GQ4X0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 34390)

`protect DATA_BLOCK
r3d448qR/3vGTy7gNeDuPvPMxIcOfiIbbJUAQAzsalcC0aZGs6INLBakpWRS3Rue
B5WdOD05GJZBOHYrKEhXloAxfgk3K6wWrSL8knP4dWGpl19VqfHmEsEyFICm6TWY
NL3OnbxeHS5ee7KRUm0NpO6toOLnMf3cz0xQU4Qy2a1QUTxVMX9FRHzqKqOZxZZ/
PIMQA5GVhZdXOqvPqbK6ER5PGZoRBM9kbxynTdXlKvfW0bBN8GJMIrVgn9dYQHS9
3T6y0P6MIcVSCEoSrziY7golvkhgtRDpcn/bOmBl8GGeAvoPyjrgAW4H8rY/TgwP
ZZX5BwPUWS0S7nLViDZxarLDuycktTyuGQfV9zOg1JLn1Hb564V3CfAgxrAMzF6m
Moup8i2QlQoUq4lWwVOQ+32bzLwHobh0XFt0g3qAgj++wguUngAn3WN3sAiKlpgh
oBkqWcKRkEOAQ2L7K9gVn7snxdOVyoS7PzSlWGRSz9m7Jpas3H9GSS+wga5FTa7S
sVZen8TQ2IE1dwTkRTHu516K6Z5SU335vf5hRfWN84GiJmFY0uBsiuTzJoDHLpu3
o5oQOdIyFqVXXM9MC5QeEGCU6xQSWQReN3Mc8St9tB74cfaDXxm8Z+9l/9lb3rI5
6kv+vk2OIPE+5IGaZpRWljrMzEtTPrMAVr8X/cyULNFYmFsNoZs0OxKhBP+buZaG
OqH+5wz9M5JeknS3iwIkOpaZ0Z2Y7dJ+8OBxtKG70vOI7vsG15Dyox+gD4NdHHCp
6HtMmYpsZAEC0r7zKMok9OOWhMthbllXyEbXrfjPUll0bjY6/76o3T5z+aE6pthw
rINlP/yNmrcCJ/bC8w6Govj/ni1xztHimZVDTV1OQ7BGaOSq7GAj6mrK/jjzVyaU
QfSH7yVlbeZ4LgoguRUzBbihI1nRtEuC2oJOX0gvMTAVIb2Bye4dJSULgCX0uIE0
ihYMqQteboD4lgqZGvfJTokm/+uVBX0w7rFXq3hWqRseA2sOLrIUXU/8Xc87GF7h
KrIElmptXi+IWbzT6Qe1XY06wc7Jl67kTNrj3RLss9Rmt7kMlUPh5OpTYtYWvmHE
2c3lv7u7YhI6jfClk4qLkBL1Xr4GdnOro3vRh/7oEAf3tU4pD90m18a4fl2DkQBW
V76a7cSqOYlCH4lgQG9gLQe81KgTrmcYR/4gIXerBXKOVu2K3srvEL83kFpDUxM+
I/6F60g6ILMFCz79GzAwGn4al9G8g5kJ+AomfRXP+kLPOelZrirFQmCv34ozfzGl
yHVLqu58lpw8ziGBfCGUXq0qyALY1huYmBR4uSwSlaY/EZPkaQgJZhfiqtK32xOA
vZMIbIIQTVoB5QkqNjXIcOEpYHGkEuh7ZLumMe/GSA+BbFUIhlzJv5DdMGOWQnzb
V+3m3XmYEiEwuWqhLIRRDz128+mMej8MEge7opY/MriOd9J0cbpCSeE6PtixBl+5
//4Sl8x2smcDiVxGs4lCMh/p2i0mnuPnpEc08+K+5QZCYX/FswZWN/Rpzg/2DiDl
tGyrEnYbWboDuV4TU74uQnlFBRhPf29molB5B7G44nJFjv0R2c96Gt0ucBKqXYlP
eXVOEsPaUEJnwSiH6iPdGXk6JHAqlm9qjLSQlRQNIX1N444r6YhZFgfjZffdnPSH
KQ5ifsBn01au7BiEy1F2aKy/JsqeDExLWoLRC4vL4SVOBNQLXfVq6Fe0jaEKD+WD
gyX6wnPOatMX2pYbQNtnrO9FEipKtD95J33O+BXX4RHPA35XFFNFNYIjqAzcZzjW
5munLT71MsliyDJiHArMMMfwcSae1h4cewIwH8P30qS/n3HDogZFuP2FgGcp6/Gz
sNflDrehN570kTYMy+NrkhQYs7rK8RrzIjLqeavnpOxKCjZaWIcH2OFLomENthRW
UxgNWIRIiexpPisL+p5pIQmxP8iccB9sDmJUathf0EynNTsWaZusSsPa3XnbGcCn
zFPXNoCa7gkVchuG49K3CzfI1dP1w/8a5VH9KoxcsNG8WOvYdY+SRi50Yx+rL2nI
qLcnhxMLZadIW0K/eDdkWnC5jVERSiFwPPCLYr0IimVL6nTVnOOnWGfA/wXt8jE+
uNYFj7aMPCAVFHJ7A7BEKvte3hnf4FuysmY/oPp8ZH3NtyRedCCHr47RkK6SDyAd
ZuRrjrBPECKgVXaP9NCKDcCSdz3W4SSKddJLP5NLwHzlzJEn8kVwBI+FgV3wvOAQ
HfIr5tsgWzMhhPjJJAlycuM9R4Esr40SyIFe01s2gqpuRgdrmfVfwskpANZDM5sq
W7BAu1/1EdciaH8Rh7++cNvIaHvlotBss4uOG1i2ibC1HQANn853MT4i9+yf3h/6
ZRcMcMZdjcdzIr1pWLLMepFiwUUpP1uK5wOe4BlXL6EtDe7g1xZfDi68IiGmwudv
oMdmPHE65rY9X3flgvJ+2UbN523wDce2QEl5l/WuWEvrfUcmNPZ9EqVWqQ+cnxZS
kFFQNaCAJxEVhT7Xr+y1IZ7XU+HdUh4TB2BJS8rLiWqimgFvqLnDEPDqO9uR7wBD
MRAZIsCKZaEqPCeOe8CgATAjoPiQhPeWUP+CHjwy0K3upGzYV8LtKflKoG0naC/W
LZCASE1J16PcZox6RnAEWXa37O4pclS+vbNmbiZOtvKxj3qyOyfkjj6YzTjqciqC
CZ/XdjBr8vluk1iCG7E9kF4/NZS+ZevFeMcsawtFT8WZU9jV9ZTM/6+LzArOGJ1i
e9qC2s+bjDLAce9GsZVpiFPrKoST9OehpZakMA0S/5wmScPosPcemwp/urmpzttN
TSa/dr54zCX4HZGKo+omCXKI1+IB/gKBhDJErF31AknJV3bK5NAmkiSp/iWNc1ZQ
dYyhzaKbnBD0uiLsORF0pGsIMRvgNS1LCINg1plnBHI1IeJavp1UX0+SWfcdpORE
tMayeM90BtkcJ5r4z/GFPLSePWwSTZXs1MjV9Vl+hL5Y7i89IMDWsPt2vb+uQedu
BmERaP3IGXeQmC8weEtwg2AbHtBPp3Sd2pcc0L7BSUCWYGCQqb9VHTy4rW5RuZLM
tK83PwVBugDFLWOjAEvvCl9kd/6kGNmDksvkGuHI96fjAWzI1a0ULbHFCbPAZHnx
OFxDqRHfJWjtX3LwOO2LqrtnFExysKFdGKdtm+wG/s4dSO5j7UjFpMCW9+o0RpRo
jfEMVKINsUyRJHyAVw5fYPINcHq0WAFB0jWdF5HKV1bLm1tJCAkjgLWvaw1ZeVFJ
O/3YYVrIJBj9BPsejcXWjM59oFNcL8w0oDX0Un06qUPpIqzwOgOPWm3JG00HOHCN
LwALf750lHTw4ygkbAVw4jLvccAHQsdeiGnphf+ZXqBQUtWBl8d9vDTDF9geYvqi
hRWc+rPDT771hG/a58oXA9qfgGgN1q+o+DkXFa+t0oGVcRIhlgoX9ZUK8Nji8Gke
00Ogd82wX/R0YnAXGt/2y8KuakjCUTgnzq+ALpzhLdV8EmP4isYU/ACctpAxPLyd
uCAQH9j2q8LFoyMqaDsaNyRIdE8U9CaSxoTdqIRUhm6/OqSKh1BsQVrtSJr+CAPG
8iVjS7MmSMp6DyfKLgypo/J8JoB8fp9NAL7jqlVakSTp76qgsSHtScQZitkMus3S
zT7eVi1O3KGVkHj4EXw7uAt7JRjXuHZjVPo6VXRDnJ8r00DurL4bM6dqcLWyNoXW
U2ATbpLGpNFIy5Wiy71cW3eZ4I8Zmnf8nEfYuywaJ7Ykqa50DmEvk9QDgKcjDMyt
UiXENnKCmsBc+V+iHDscpi3W6hnMh+v0wYLysLtVWNkgFiWUcfWahsUti6UiBZCh
m9eUJ25eoVOPFR6SzUKtrg8VAug6ElIwDwLy5n4rMk3OyOlZBWbw7CzGpx3sd05m
j7pu483YwnW9IunBlaO1pIAKiDFmKGsywrT+n4JgOUS7LE2hCV36NPxiaRF7SyUW
zUn2fyIlI6eUXwGSS0jvrnwnB35LHrpXYr/4IprdFjEvqDNB7bsHByCr9Ws0DP09
xTkKEkH05s5lF4lCJ/V6j1gFIU8fSZqnLVDyJI6C75ae0HV+v/VR20Ej8RChaiTX
N62vLyde/MA5bjHLGH18WTttjxDf6HjFCbnb3siDqmljmyyHpUDBjBN03kLCiC9O
14j1iRZQqKPIVubCHlf8sat73GstU6kcVFwyLpCwgNsptnqV0JNzomzO7PTvNRVq
IeZ3asqPVyNMglRyLyHWn8oKwwTbgw5F2ehaf5/2L5fmwA7jR6CtyJca5oi0dr3e
ll+ehJjkY1lVTeQwxoXafrWLdi//MVI4OWY57JCzy1GNcGf53djht2eTLf+02WH+
MVNSQtPwPEoex+Iif5b9IXIXlExzAIoCFP9H8a6hzWZDP8A1H4oOIjyM0R1Dwq+Q
+vaQL1EC+yqM2NGCBj1zaq5QuAYNclpXdZXwTksJO/cdh2d+W1AyXTlwFowYp4ih
LoGTmeukO0zCs90GbOoRMH4LVnUy8NKREBw2bIz9/hv6qWLw4B75wkx+rqpqzDpk
PJMiTs2MRvQdXQ7WjxXZawpihlHYeVY2Ut51IF848XJjUAv0vh8Y7m8ccPlDAiyC
Q0fj1cE8JBnoJrotou4XGTGF15EAnkdeCpJHUKbSnmQ7Lp7kbgi6wekjVgbzqiLY
mDPtFc65lAGQWERSm8T2TJduIX+RPsOfxK6JIwP+h+PRlgToeKEx0jyStGrUuLax
uctlghogQpdFhZ4bkIWIYb/CZiF5/ePDGCi1FqFEBMfxRwMq8lOrMcf0KFbdP9ca
CKMjVKvnWlRySif2WQamMqwAZqgP0GS0iUabVuDdniwwl0bMISyRa6Mn2EzmO6yi
AprJCci7C89W/J9mLeJHmqI4/I5Mc24V8G6yiKkLUbGFlN+3o57H9qsWw04f/v73
Fk33d5S2cepbDWv6MXvMPUjRekCy/9Qz2wUOlnDUn3dQoVgdquk5SzERUpZ+DlL0
GuSE6YuM9syMSVUBTyrJ0wZu8aJ2xz9Z4z7Kyn39ESyurkqnW4JtsvYr7CCbudHu
NXD3N02Fm1m4cUwj7bMeNuXJjCURkaP/fiMXgeP7nkoVDH3xQznmD0Mrtc7Plfqd
mhJAriFIOnUdPkl0G/4sc+fSdnhY/wvcGUq9YczI0sA7RG7d0Bt8VMR7QO5w+AFn
wzIRJxX0jHGYIxJuNhexY6xyEtxPNFzOPQl1WNMbLjIJzyfxoNq+BYhZvu47oOlv
oSQxk/f5fYiTeyAd8135kAjCPSxHZfBrlyqQF1iQsDAhWcPPwhU5N4iUsoK/RkO3
hBm4kN34vmERBbNIfh0eo9Ko/GDR2/C+PpP4+XF2THQwNaPLGe9vAVPutre26g48
6vZRYK9YGHHtQscs0xqL3o2QLtKo7USaZEWXHWo8kc/C5x0IAVaK+3NJat3Q/pZ+
tRsbJyyyS6wB8RhV3BDsLsUpy2AgafrhqTjZgcZ05+8vpctZKf1P7hmjCmVktDmt
trpEW+mdDssnjDCNOCcN9q1b8VVPT8Nxh04fV5PlF+NwI2fu6bjFg3J2rEfZQw0K
curax/frztVIlu5Z9kGo9l+oyCiIUShVRAvmfMcjY66zSt4LgLsZrztLXaFcB3rJ
IE76Xk9/KTyvGTysojDq8coZ529umwtQVM/gSBnRJo3V/ln0WoYRWtNfbcQbboU6
SdyHiNyxYPQf7g6jgK6DHG0sZmngIV3fi0KR969JbfSQUxB0x/LRRGE0/L8LQmpu
At6ff+BSZh05XxaeMTMF+6BjozVffeykTeNb4anQq0Kehl18AysYL8oRmr47Lksq
iyFmkYLFLyUO56c1emg6czNlpTWttOEyMLUNyemzscRYZgYl74AEudJ+Y17Niv3b
nlLDuf1R0nDUPztonxL0vLOXXFDhZDcHhA7SBfblCed1BfbDdHNR2hkdYxOFfSrd
LRjimyNfqOS9Cd+pin3UJR4ycLv1plCl+HefihZnagOBBnQzti8rveWeA7r3Fy4O
ZtGDGOgPO/BDXwjmTVBl3z/Blhd4rkIIq4INbcAT4jrDh/pT0TVP++KcX17qw7/E
GTffQRw4g54n7YHarHQgU/3skqBoR7BKyinWSV3xmjSLVwdj7R690x8eJzfYj84n
Ur5LbhWBnO7kVdiFlMcc2DG+E8OFX0x8gq6vSX7YaJXncV4D7gxnTGUVNolubCB9
xdDWZy70R6GIgSIGSBmButz4N+ynhpF0s/Ffy409OXR0UN7FCIZ64iHifyBfBX3A
P5i78zc6tewRKi6A1cxRnjSziesaDl4E17Up7KKocFuU2zqe8p1UCH/8v9pGQwpu
OIQeryvDU+unU5rlf8p5vF6wkyefAWbkN1sW65sVoObFZc6HHq8Y8NHFQYe513UT
MqKuvdj/BK0XhGfLZ5iWaBruuNVh5Cq0dtNjvEoEvG9aFqoH3o+lp0FlB0wVwCIl
5KjkQZhzJBk99AO/UyrRYZaAxtTaJrOxFowIEy3E2JFY+Xlg0zEo30aynoTgb46o
JA6Ktu6MI5Flg0P9YNKVuO3/eWnqor1c/GNXIV2hc7JhRH4f0kEnxNjlG0spcLit
ny9+k+arF0mk7vfeSiYpWo0T5JYeY0a+r6vfJ8Jzfedk92ZnDEUvK9tLs6XVD0Bh
7LuGkWRAeCXuXNMHqvuGcy7UcX7e1eNDHmn4JzYQRhvyYa2NeCUqUplTmUKl7jZ7
10d/aeW9GCwtWqnhQvF49JEQLcQUoPRFR8CC3WFM0RW1dNDY7QgrTrJ8nCrv2nVb
3wC1B0S1vjgsDeFuU5lz7jMKvbehQcdDwxa45nOyJjttC6cGPFTr64VNjZqCKYcN
/aOzo+DRUJVs6zE5osshJ7/U28yINkaGvh3ppgK72klSsaDgzHChvEadzD8vVRjX
OHrdPISxIkGXRLj5K+YZwau4s4Bjc4x9XP9flLk3OTR49kQbTvetJf0fdx+oIYTU
C05teaYanKpV4/BMkzayIvLqkyJ9NTcP5Q36tjMnU0rpNVLS3spAwEtiIdunE2gC
Pg0c+8C3eud5a1PORUkesQPjIAK5N2QzgCT8kK+IBVsGHv4dzxHlZaBFyIVRLIEy
/Rn0FkY+HrNjA+rEGzXr8M0wiXbHGnUNRMJXMSeice7CGwCtqkBYN9lC6piX2ZdB
dN6KIey155lazJ3cT5xzS8M16+FRKjxr1A7O/bthRgr9PaU5T6y+kEgKmxt6i93l
kqyamUqNikRNwlkBd9cFC7oM/U8Isv2bv47j6y8WBFB/JqhUcui9aqvmKoSRRn7K
gtyQmHr4gkNWicPKKElyINIOH/AA2EffVxP+Am1CunzjXbgERgt4H58bKh2VHFPd
fFXrZ21LRheS8ORQO3YszR69hRsWlYBEw3XD3oEgh6qiOwNuLa/Spwu2HJWAi1ht
f1rnwSToZVnKQ3A6n3A7+GrDo+sqndkcrXfnl+S/VQk+reKznp467zuQKCmi8fxC
7YoIcbsA8G8wUPXgtTstHUYLwTMx7T7fOjfzkqbb20vCPHLCIc3ft3+dcpwssSwP
hMUuHxa1S/bgSp/VsmkcDJy165Wy98DEXJObv6TrndCIWrh85LzCpBAROsvPQcn5
K4HYwOhNEumlEkQyCUrPVKWhoIk6i+p8PdPngrzAx7hnRlO/h+36miA89tjIPGzt
lK0hxUcvN6zWI8skNxUsfcIpwZq1tF214AS76CDBSi1QQmF0zC0Req3docDwy5Od
2L9Er8SdXU1LZVdNUsjTl7xKVz7v7musQQv2XRzQl9RQZyoqCfReMA41Nj3ARLyX
qqON9/fsN+Z27ftI0Gh0brH1OIXk4JnQEjoVcDgv9HCgQ2AQdzR3YUkMiZCtfR80
ZJOaaEKomrdxDmmgTc5eb9+DDjqcUZxcLN1kMBOOOxPwU4DSRpK9pf1i6YUvR8Ax
Nv0QhLEmElEuJnoHipl2d4kTnsrdaPBqnwDRkHsSy5C7oxOyNVAAKZ7wf7BWUbIi
a7R4R1GXH0zK4nvkOpXlxYdim3gX0Lb+kYyawntdHJBw9X2yFApnUq8mUL2CMfyn
fzbec4mFS8Jv7Uq5m1skFj28WnpjXZb//A7xopjdvAUysjfEfKSuFs7fx3hawmwK
4EvK2ywrt2kNEr2whMlEKrBD9RNLXbv0fI0j2TibHTvgVEvx+LUfZc1jImRpCfpH
L70PwLtKLqWTwjv1TUzpW+F6eTGAIBbGIz2kUXmI0rxVMTAz2+zYFwRtsDzpWmFI
zit9lDwXQb5u6BqoM90RHzR3WrRK9j3XyG+sypo/m+u8x92wds7w32rmgDybV/Qc
zENSCabW7IL/uQSXWEGdJo5RCcWMizy+HS7GLHXPwWmiunK3mVV2PUEtkaGqmROI
YZxsZ/zMae98uVx8kW9jPIMxF8CGwdqMm6KUReMJJ1JhnIX6/pdZE88cC6UTCi1s
usZPiLdjRZGT4cGgxlGxDkajJ3X2+/P0zEeGrUiHR36eTkxZ5o5Reny2kOvrK9yu
4gaIt9dGruYeOGnBdP0bhHMjiUx9IxC0KB8t0Og6wDd0vGyO1PW+fgluZL4M5cpl
1y2MUhvmeQ4JnU64d8esCnXj8wRfQvAWOn9z3DS+QjYN/1tgLAWsR0m98DCZrI+X
XsjA1g16ajDYspTCts4HfIE78hIqcIf5DoBZEA/bLDb7Xw4zHw/QKLkNl6o/3QBV
Emz6BHYqwpyrCzjxn/gPTfFWv4Ssr7zlOFh2sixLILSAV0H2+n2VQ36kaNEUO7tC
2EzryE1qCSWgp/HUg/v03CC0xb73J8kds0yHWwoGbpHEhrT72gVUObwrjOVmgRcC
BJ+3tD/rEWysla/WmF7F+5bJ0UNdXJ4+WOUtpV97QQxc0rno2fXqhqyHFWOpfu1X
LlZUhD2C2zYp6M2CEQI7barBIKN3ik/NQDsyh/AjpfPTjr3GJWgh7JOA0fcwLkiy
GOrdeq+7UWn3wBt5BZTkWy0YD0VVM6A2oT9y0COBrEzv/pNN2cABW3bAsXlnW4tP
IbwrRSInYWK+rkbKuiPKdjIro1uq9pzR1QMPpTNSEMpsBE2rSE5rOBaNdcotYDMj
22rBy8ci5db0cmNaHEJN3DCzthHGxzsW1lk4MFLGOfLNplEBdUrdPPYTdseO5Ljq
YpHqLuV7Pg6b92gRHeiGo8QQs6Whxw0QIEMHbBWHQqQlx53lb5IQ2c6VRiSSmyYl
kJr71ucMnftv47YWJ6abW+jiw2GYvUpRmn/uVmOZt6nSJmvuHo2wFfVfuxzQz2cc
GI6165XI04PNybzqBbwrIfWzH4gpsbtck/VdwN1BAIB8mBEPANqw8gINt8nBXa2e
e+S2U+wfI4rADXP/4a04WG9NpoK45f2ZgzHI6QWBox6zLFkFVV942H7qz0HnHE+U
Io3GeWAaohzL4tGmd4mQvPIQoI8WJw6vEAC7bNQmLTH3IHcUENKZQ3FYNWK14VYt
J1uwjnSsHzJfiYouQBKXaxC6osQScb/kUW20/hrQ+mYDeQIX7Hik4on+0RULf9+T
PHTVrosxghQLIE+NdlhpXS8Kn8AIJqi63u0PhMFcohcSROKQBdUtWzmCW+EcfXZs
YnzR6e8r+QrDMXLC9BYob1qdKlaWGB0p1YUMOU0axJKAEUDz/aTIXJSVQ7AONoHE
SG7Q4dBRv3KIihmoniNniXCbVG/D8vRoO/z5Eu6XQoTtiDbWEMxjGul5lNTtUk7S
ylauuP/XpQRG5RXFw0SNM5OOxxkKaO4YmqCtC5b2VnfS8jGiAPie8dIU7oxrhsKD
xDmBxg1ddi3eo4x1PrOqEu04JYw8xDJAkMT7qKWaxzWf0DSfXWdo5xbLskxwqXmG
1HfOxUpO6bi3NRzf9v1+6VqVu3Yz+6ujhVRaKaYBm8QZjUAfkBsLDM4/87+fX5Ub
nTiEtvWyNSxRwZg6QbbiyVCBuqsFC3Nmex6V3Yg8eEePlYNY2baoUexcqci66FJu
1lpuDsa/Jheq8Le6aMD2weonU0DtlUDY52kswWDqS1uBBlNRZEBPfbg4500Te6/s
ooVJKbSMggFGCirNSPXr5637rHm6rpaRYu2ZT9smjVO0onZ29vrbQq4rI5RAsSSL
eEIc1MkYkKpT88Uo/kMsj7EFYxfvnTh1d/mEzSFBMFmuF/NU4sbIx+YB5tsior3f
ioFGJaoX6th85LZAZq+Pp96KXcTmKQ0KUz4TykN1ITs1DpFUoukn+0muMnSwSbad
j3C4BrLoFNEE2DJdamDCWgSG0ha6usm98guYHpxt5quAMIS370482Xm0Wp99zQ+1
Wef1feVTJBW3PoXelUJSoqsUBLCMdWM7Lkkr03UuCGOXuNIUslwNXyBhLXjCc23P
OnQT4cPb21gvGYbbe2NNuVqhcLVh/jUHgmcAB7Dh0fLLIcC3MSKDmMS62uKfwgLb
Alhh7ioUEOusG8aANwLg+o51NWoI828h8DKHP2Sde7o47uf8HE4YseQg3p01KWXj
TGmZ2GxEj3xOVxP48Ljf8qF0TWsZDoTDz4eOTxGNi2qth+OyhbbEh78N0YY9JfOF
l2MukhJGckxpecsIYSljXA3FR1wqK0eW3QEk9c80ZvCaZtREefGxQ8DWD1GKChJh
/FYxzIshm4kTjMO+oGsIkl2H9CMRL+LBtHIqVkbKMtPq8Ldc9pJC6lIbkvkg3rUT
+QQ0T13bW51gMg0yEUD83NPXxSz0+jaXvpwRfJKdWDJpNFBWFKib628IZZpxZEbr
rSy5R1t6+uYlNtZxkJVun6y7Qm2whFVpwIA15kv1sj9gvwB8ok4I0yqplChXsBpl
5mU8oOr3Wtg6uZmA3b2u7SlfDPHi8S3Gox2Glcg1spVTf4FlZfEvRswTiyLyJREu
APXJjAEpA9Owjtvx88Nw3L9zofkquCeQdbjFZtnmwdWeC6yl92A35VelgemHi2UU
0Q0LJAGCLk1Nm1KHYPS08DuexKF+pyMtKf7XEUA4eMpu3x2riLHdDZ5pFT1rgv0B
pyRwDaZmTM84MGnMioLuPM924aD5vkNdgg+WQ5VjMo1/Jfwino8ZUC9gMErNpWl0
RHGRj1H2pXMiek8X+AirF0qWPVvnm8hQQQsNik/byyKZfrMHMucyqMRbj72G3Il/
DzGwi2ub0FApZAeCKHSh6cldDjxMefoja+4Ij3BbZDKPMXTfjT3Q+JDGGKcrAa/G
zKpkTnINy8K6lk/iZPnO0ByjYQ5d0l0irV/xMw4ojdvEfhrOK1jH/6GunJ3edOSe
YBUrYCvZzUFHeT0lOgZCuTmRWwIHmnP2s8XerwUOAJRXYMFpn1EBsCVQ0t54Kd3b
d/HuyhWQStO3sI9GBXdqu2hDvUZ5KFCWfOltHn+8Y7H/ZSmO2fqGkVgy8TtYE0RB
Wy6LEvViA7Ht3pJfRLXqFGEHQqvxW6WG0llu/dhUYonswQhVFEnlpG2AXhGpqMiC
jhRXdrlUOPdrG/2kvZpCxJgYLaxX4oEUkJQxaX7vrfuV9ipCVmw8hNivauE39ruC
QX/wLlZ+yt/AG5KVWLkJ/E54cuUTE8chDadDhlAE7lO9+GKPwX1U8jutKvhFxhN9
WuDCB2babxcZIZ1Z2A/Fb5T2eOzUFRFC9J8R79wqEr5UJNB4LvkZ2xjOYpQ5JHN/
F6py0M7AOTcNRS6GVr12uSqw929s5q4+0pKk4/KEhQy/85VWBCWxPyLYCIpzLP7K
+DK8eW+sUcSa3InEqyDATsNvsDpePh0BQdjkoEwCmYkpPzTUem620hV69/11S1sP
y1h/9U/kghWHFDD0GXuHsuGiOEXk9c1+Ay/t/r6JmB+LuEY/bd7WfS6SCvVBRuZS
0x7dI7e4GPiaeGHdj7AVV8YBovaV2OCNeS4PfHdUoXcz7L9W167KbIir3G8AAJRN
UC8mOWHaUl2jDpR/k8nXsFHT/uRNJamP2w6P8jBtEqKjAIIwmYu0TnJPvWbIPQRb
Yq2WmtrPagT12RAt983USHIJUptckBj0HYVnlwCgCVqYTUijWdRN5vWDCFDjdzbK
6y9AVrSpkO43rhUu7mlVXcdesPjphWsc/3BwNK6pm2/CopYxCc+vA69G+7ounmQA
Qbd5sVC4BuEDGqdnN6F8yuOqJ55SZu5HstWx3/B2XSQmEMQI0zWbfv69roYYlizw
lrrDH6sR6P+mNh3kgWhHL+FRVN5UYx/3rDzj87lxeMnwnAwTC/Rkyrn5WLtJzAcy
vkr8fBn9pKDFKJC0pkL7ffuGOe/6k1LDh8AB8NXoeGTKhGRKLpcuXjACk52jtkK7
/dGrpYgyFoFh61fHNlatW3rduSE4zujyHbkU8EqtRo/6YGGY8qKEOpha9llxbU6q
RqRHZ7/MdKQL2rv9cnh2SxFXzecNF4cSzWIvO02bDaaWi4jy/0Wzv0PXpW9ZUf0Y
Wlu8fDg9JdFzsDU3Ry7/5h77EyPf8zjScnA27MImHH4TaPZyJ3Fwp3un064zl0AX
MiypHW6ew6WEYoyR+0v4L2jC7yimCmgHw2rSCGtUrWCWS096MxFDMG7S/8J0rX5q
gq8GJaVuZBByUWoYNHASWC8CdX14aaXTsi3tx8JKw6oHzc2x2IKG+Hu/7Yh3Z27E
RobQj0icEL037pS4iJTC2MbWBFm7YgVcwgRoiXUqoE6SD9vr8yVJ44bJgiRYXWhi
HXI/QfrvitcXb9q5ae+ebMQKA2r9Vf7QvXfbKAOXryo+zSfS6t7VGlPoPEvIc1Kk
H0EhJ9h6Id9Wf8ry5/fPHQxo4GM6fyHc0Qd2vhtr/QyTMy2vBnsGL7nRucsF/qsu
moaZCCKCbaok1XL3kbm7ZcWJB241bU9eMDPHjnxmdeFR1dN8K2cA13DBuCpac5Z/
EFEMQ+WD2M3KlO7yczCSOTK2gAwNP8GXlIw8kogL/Uo6S6jvSn/K7BvJm3sNseO1
xveBu7s638VQCyBI6x/IbdFoU8UDylTyNQ2lC6+sNqVxaWHwhDnZHdDgbX5Qlr+s
VHkGOv5x7XK/V2mlmNnbBlMLnemjH4Xx5FiEWYYcn/RbFEWFnPHtPpQrVF2TLtFZ
M6IdfVE3xUu26yAoH5XAUWSV3GIJCgqta04sX/D3kZlBBuTvKgJ4YyHKOyrnbCnl
Rdg+1fQn2wxCJ2myj7z6qYIKCDCUE1vluSfqBor0zTL9NIY6wbbL5junQRd3lcZf
IpL1QI/Pd/lnriOCn94Y0gdk1dB8GzY+hp8pZ8fOPhqFDAabS/1ave+VaSW4GC3M
rVp6FhCJitE6Gsu1zS+i5y8aI83SMriW9qgnjEsuaYDCdVv8asvF8Yr08VllJHiM
EDF4qfQ4qjGosTN8Z3/W/or/ILI/5/Ms8WWKYhvJb88f1zss1XCUY8D5EKERiJMt
FY5KGA4tcbqrglgwQnZX4yky9FgHehWzeKITHein4WRelkZxPqlrWEo5UsZGZHzQ
Ic9xz5Uyi5ogB10PnwU5XKdH1F/odkx6kyOwUBMroTBPLCDHwdo1VnpZAN4L3rPB
e61d6TEQEilbgKOj2HVqWazCSppDUVP3IC+X+457DG+kQ+QYctjw2n9bGX9Xdcl4
1g3C5i3eATnD0UP5EJT5vYHsQ37N7G9o8D+mi7oxUUCt9zT83fpM3e3xjKjkZnyL
Np3iVOo72FH+DTNmRVqEV+SfKwkPS18mQuzFgkgZ8iWzgMA3MI/oeieTOrzmIk7w
iB+wJCrO6P8IeSqqq4qnbXJQwCvljgvPK+z+rZ8EdsNP5bPI7sxSC4nP2ww/CnOb
mM4a+Za4iB7ni8HXgF5Ik7hAoFl1j6puZwp/GEN1Cc4vL5yAVwyKvkY1Trh6rH54
/kQhGWkmnnnldnNqrPaQw7yOp1Za31egCU7pRJSAAlsxRABwgHWdpsrHlZ41lD/u
d2Qd+9pThvt3WGMYi8hthPzIUBqMrvRnSLmNaLz3T89ZwybSq735rJu9vcA+AlPm
8MDkUYvzw/VD+v5mTyUViBSgLw+8IuFGb8T4v8qxcnGkHC+OOkSeGfnqioCIpI9d
Jw4PNIOZqXxD/6dww01d73sqDNrwTLKgHGykQyLijZQXufqc+n/9pX9OrqYhkaPe
YTgdyVatccDhbFqUxVbYouUxDBc+1+R30Dn/qyK1ByU5dHUI3WqVbK7PYK0UQu+3
NuylThTQHrSK58tSRlE8w22vFckp1XEf7GalsxDkKTwZxZWfdipSxLIQnF0y+EmW
USXna7zMj/tF5KmYo4GFCkekqCo2ztbYHnGjdumYqA7xoUQhDkTzUuNP7mvlzgS0
OV/T/9mqd4r/57BEHVZwyubp4q4gUGBdY4MkNpfo86ztTyXTHFkOVzi5kB8Hxhrj
dydMhvJYSxjFHpvIthtzjM/YRYltfGsxEP2rNyosettNHmDbAr0FW792jYWM/dAa
BNSPt0ASIYxMqeyUmVgxyBqaqPyRivcJddhfpy9mZb4Zp2JNgMN1et3UXgha0WH9
9ZLK1ZAC4uToZ/lHFmIrLgKoLkhbTcT9uuLgLtEm+Fe4O/QUI8S8rzFLhTf/WGJC
uZ+7xb1rhlj9PoyPkDAH2TzZoJALe8rPOSSYsB4EbQ0CMwVfmCIr8OwzRL0PnA0F
uKC6duihltRwwoFXXnr1KZhGxN6b3yhTOqulOHpkhlk1T82XfWf1g1YurAgXeq4l
Eso9B+vjYDx3JRrrP4XERHWIMiI7d0DLpsVAhOod0dbp1ThCnjJzXrllVdrDhdXJ
9kOt0KJJbgwWFShJOZj/iUpYoaV5qvjbJAYNNo6YlQkEd7WSQzQTiYQ7sSlz6s6J
zCqToHZjifOzXVTVx7f7KXKBDoLdkMMPrx7EVqEDtMEScuHJ5j/icQArviDqiQjT
TTIqjZYpIyAsx4K4DYcXve0Z3UYMjlENB1ZYK1Bw6IMyxGrVP10ltuoQzsQTrnfv
daqwwVHQhrxQEGyUmLlFxmgkrMxObh1MyTy5bukUn2X9I+iMskugP5LJTM1fa8EK
GiVfPRLjA06QpEpCqbM91agDJcpzs8IUtTG/nuYOjLzPcddpZI/zpCU6LDDnX14O
Qq/1YNhfwyMUFODFIk0mjRiA84YS/pQGCHWTW/71Txp9LG342GS+JsCGg2jlSRTe
iWAIuCpcSasgpWlnUM570TKxHY+NKxOY7Yda+diDU741y+l8b6Cn1s/w9biHKBS3
ojDR+9JmqUTo5uFMMH/ltjD6fSWzu9Qm5XPznXR7JxJ6tDxaS9rP/I2o7qjFaf71
GKTROvH0pIbYGzAWFAAhhytPglPBRStXXbmJ+jmKnzZdJRbLtvndwiFPgG0q1y/l
zA7MrrvWrTC9n98Kh27Ey7TyJZlvqY16/jjUPMPhPdlhcIO+6CJNuNa1eqiSqhXh
Y1Y2tsu9eRygrUN4ada9kvdMglTPZKuvs//tFBMdXr2RL5Z51eCjucIQ8tL/F1FV
eKvszF0E/qHOKXzGa+7QMXOUJrSxkPGsExOV0MDzPESGnKyC6kBNJJLV6BQ/X5hI
hAxNt8UYbtEylYg0AWopB4gWRqwqWI1fauRuUk+mO2wfQbD/KeYah4IvGLok804H
18fkq1A6xB491ycyXqbxbL1uoxAeCxjlCUn4DeLaOEnimL9msDdQWQZWvYi+izpo
shg+N+LBwFCLyffd90i174UAtKHqDPY0cN/fXc+kFJe+gnljThMuNMgHpklLxMMT
1NkVO2puvXN8B05Gg4JIaZYAnWtbLTGpqpm3IJn/SNs3K40XekyNl6jzw3ZkrJ3l
Ge3GBqGLix9cm/Ux8MV3Tj2I/Xr9+bfN+8m/4tapNneoVAQWA5ifa3yuZ1zumlHv
ZHd/yWu22uw1Igfwm3j2KO9h1afRtqfPmWIRAxy5oDMJcbQ2MI4yBA5s0J0aK2H0
NBRFZ9WBxRuRM9T8egEVUwCaeuWTls/Na382tXOGcIG9QLj5ksr6Jtce1SZaLk0B
FC3QBN0AyoZPaClZW2LRsAm5JHhgWbsPtAMq9FBySZSC+/gIMcMeNK/8aJP7Domy
dIQbniKJLH1DLIOlflc8y2bZzgF3ev7fgLxjeN4Oq1kLiY31ZwQ1LzGML0tpxZym
fWV7iGGOf4IxLo+iwOqOnLun0SdSQBfWQa6MJCAgDLD5w3X8JJrIdjUWFQkkBFyS
1ZG9dM2op61biZAuDTPnuazjjdrK7Gu3Lp5nbmd+oOhIWEJ7SU4216Ux+kRKZJ8N
1wao2rTJavDocgz/2ZFqpr2ceCc/uJzJJaJAjZdD9+WcfmheBNFLJgjBZ4RWUtxW
1pT/ajAmNFGuq14vtGQ9W69Fn4Sp2VmQbt+Kv14fteQLPMh9k8OVCNHF9UFH0vJf
Ig1iEz2/EgsOgFFCHj5R9GNEZyNPhWxtSm2RinWcP/A4P3Gd7WUZJhPmhFsUhDu2
AL1VkVKI9880fgcBzG1TpreVdFJqoltcWA/mA6bebXaLySdn6tIsIoCCt/m00O8U
m0QJ9YdMNUKRlWGSBZI7R34apsyGBxfnR8It9r4vSY9q17L0+5deI9Kq8wxAH26V
UJ3/KOLiVcXX39rg/tctXax6Vj2h7X6UW+nKLDsoO452QU7iCFO8cbVX3ybDBG2A
ZKQ1hxNl2rBAeouch8y8gRxiVHMcmDtegjtzmf8Ceaq7o1Va9NVY5fvSvUe40SRa
Nvfq5pDg9O9337/Njv39kZnYrke0GSrRoNY6/XAPZ2y0LOWmvxpeRzI6peYmfR+f
XhvR3vGrQ5t1ilREV/GC7iRhejYUGTt01Hkyy96vJPIxujv9FLeInAgCJobaM+yy
c+y2FW3+iCG1fBKMDYHrV+2ornsxLuwKZRDmnV5Hh3rrpGoZJ8quBxIMNKauUqUC
lapc5v20+p+OEECp4qXmS1Boq/dBLhbnVnipYrfaW+2fA+Or73RPR6GooUxH7QFu
Z2HhmlvhrKHCqaGy6nV17tZtFDIXtu4QSAod6smPmdKxfDtNdXTi1nmPuUFrmMh9
iGllPr0YG4osxvpHr24cJH40B9hB5yPJpZHlwIKyw41bJGTeLIi2QxTYZRzwGNuO
GXDjrDNOGGUZpmApzUtHtDiYMpiAhykEnbD9tybxMvD3YtppcbsYpX8XVA01QmPR
CKv8wvksWXOcMQjasgGemyh1vy+RWQB3gN9vR9zj6Z65Q0Mymks3OSAutejus6tK
ti718omflQVETAyIRuMd1f/ajxuFKWobvVfkjTvFBUuZemV7ivSrzqJSnKgWOHSU
mMP4UXZ1TI4glHpijlVGvKVvWGIvYCndAZSqvRhRQs2i1BAYrG2le0SfbaPu8kZp
vrgw7QIQmtTRjXOYiEh2Te8OdvIntX4m5aVlDdX5SSccjz7XhwAD7Ip7yXJWFbbQ
oQwgzNuuoahd1v8HwM8Z1bhHPwqTMaidMEsdG7Csf5hQEBkuSgRaI0nBsSs9Gte6
95jr3PCxb25vMjxJNcXi2/Vjlkw8XuqrvcF2BhN8y4sW2w+APJ5HpXRfj9DXNcVi
pFfEqeC1U/rwpWlS7reaJB0KVIFtcBjWXg3lPTAczaBSdBuKDatLuBi9H0OwtYwk
2j0ukUyNR2nlOhtgZk3WFtAN6vcdyi1P62FtKIgxyIuhD4/6BSFionM80POWy6D4
LuQpJpgmZMKQe/JmwcxMdKym38m6qk/ZenhSP19/rQqVTO0TVFIk0F5Fgkd1HfBw
g5P6ZCg6sbg8a8aZyGwtW5MelTJL/tZTCFc42I4bJDr48cTrEKNMC5IfrttAnEh0
Yu/dSm1pA1zAZRZJCi2bd58t4HVbJB4wtK+0XbsvjdZGWM+vFp28WY9CtWhucma6
byEAhY2qlcbg0zKAGLuj0PoP2Vxb1CuIKjowEDB9g2OyGTJuYipAPmYqieTgsdQ0
jZZsWgtfa2gLSaWH8oVDiS69waQ4yUdum/6IEhOx4F8dl6pfm0VNcH+GGbITt1Q0
KDn2SKrSbk9U8Bu4u2fZnvs0ttiAEeQE8H7//7BZEH9uXEPNhmJLjdh+jcFX8zaN
cMOhlF8agUDP9zB5dLm/IaDvEwWyXdiAvIrDrNQQuUveWesQnTewGxyWOnpUJxro
qAiZd02qXkXvc8WgqnpK4MCsJ4yxNF4HkJeH4e3CSkHz7HHK3PCoTuQVSKbArlg6
3sSjFRB6tNIx/vTERc0ubzgQ5nQmvV8kVl3ND1YWtjtkipcxbM8V9AtnopPiGkoI
RSl0oqQ6Tdq0z2zO4w0bn5Qq6kFaSiUNIrskcCN6yDwvFeWTaI0AnnjZsHrqzSXg
sab3DfRRz8m9t6AvB5bnxOPQBILXOdaoVuQT63JGTvm+3HEfsKsHVY8CuWO1hGHL
LN4tYn+5x61m5zVgC3qM4AU+3h25UtVrMDWmwyAKC1DFGBderZdZ6DXW7X26gMzN
85LI658z2gW/VDg9Ovelk1WGDcJLofJ+7js5et5rQaEowZ7hCuk6HPekbH9gOatX
jOZ9B6/8ggDcJVIBDvMcLGps+aOjHGOhi2KmeDg+wYTT6v6hjyAIfx0iFR0Gl3vV
JzvhFOPIyfnEU9WQ8Xus6eeQTJ3lHONnJHhXlMINyRU3AW9+hx+zIxuRpQ5QD4qz
HDCJAJavGN8wlLBm8uh0J5JThsfMcCXLc7aW4hncS8s7f6G3odUqxxLNTRVt6NhT
QBaZh0n3N3QQuFpbRMbZaTwjqYOYlZ4o8FnE9VfiVejJfGPYsC/lzsg1gvWs5sRp
xQGqf354SELPp8py57HJXrolopFmgL2T4ueSg/k+GzLUwZqW7jybfmIXoFCtzn7J
O/y9PsCxVIWdnf1ksUEwhxJamk4s0cqmsLKBAvbGG+uubjy4eKRDg4jSHj09WWpu
FGxcRs/c87ALVwQMyOt7KJ6mfWW5vhqeeDouMN4y0PWbUgMk/dM/nUnDRCivi985
8/I/CjNS+xIukNEKbVdv3i/6gQbV7f2N6m51nJkXQAlQ2rJ86qiTa0ONliybhlMG
8hgeuOtM2e1LMkD0RLWKOm+LkSkySquKtg7Msz49bVn+dsUDry0EhSIn492BhzGx
TFpu/shT1M5lsdjKVRl3kl/e2sJvfYIjumoLBrjtmUwXLYx/vKe8zh5MoSoeeYSX
bEISxCQMx+LZvCdleiJlnyOdQkJdj6wbsT9Z/vf/QnYICDL0rbi/6aCeSL/tlJc8
NK5ycv3IF20nPcWQH580eZHAgYKKoGfDpBr3WXQy/dLRa/Rx+cF5lRnkCZgxC7EK
dOIAoAcKnVSHPXbHr9dhjsLsaU/Ca3dn+qSeFGns3a5Hgz9YF+rEXynvIowLez/3
nis8mTC7Us/nHIhMnRbUn9bxHlk5o4e1ZFqggebLclCLAHX/BECIP/86ryR2zHRD
b3Hpps437ZRdp4xBfMjpvMFa1+e6sELin8zm0xS21lLYR36fTYf/5IMyksJ0ZdFd
QvymIhT3HoizCvlYn9KhulIEKpXg9LPhzVyThyFtU+0x1QC18jXECi13LVwIvGen
AcX4UID22oM/HQMTARwPU4sOqNtekbv4N0yFu53V7VCGfaL6eFGhsXd6SHDUcxl5
a+ZvbkCsoKFM6DcNa4RlJfrMEwQBZzGUDthfsxan4V7Vsq+XkcNyjS8k7qP6HAEv
wxkjca1uWn/YaJsZOae/q7u132sMe+ESlL/OfktV+DKeUrWLLkPTDb5HQ8S/cVV9
mtL1QRao2gKXH+3r+ennpt8Y6ilfKFgamZ/aCeKlJtqOb6sjl+9N0S01Mi74mfjC
FYhRaDfR2X5r8+YYh+qZSoYnULSXFLsTlvgjnTyjk3c1nuyf4dFd8J5O9GpTsVAr
FiRbqZ5aFmyrGHuL2G33oyisoCc0lVSg8xTyyH4H/IfBVqIENUQt88jgktJdqt6/
/2j1F2NMKHOAMS+6+H2aaUOjB7pWJMBz7Eo7EB6XnTFhgrGWcNIbaV3FBN0Kq+C9
5r73iL0WS8MAwpOJrBsDfWZz9NMwIc7U6No8zIXVQDbvTJi4txgKfZiwJ/qAkuDy
4W6PyUbxfAaG4LmXgj7DJFfBDckgC88VZT9GIP454suDbRSki6KOO638WccUvOML
JzqELZPR5YW5i+SyvHhSPOKgg8HpRs8rkvsSoxSaFEHHX4IHF/eA5qEOKBBTBcgy
IR37P6eIOdK6/IDpUIo1R7rzDEFPZ7ia95TVDpe+n4e4lrYULpP+UiIgUn63Bj4Z
RbFuOPftmF5S3N7ZZC4zyrSOwi0LYCgQTg/brV8ZYw5OshRfTMVqBztoZ2b0jeZc
sYND59sxUBtcyq3dud78DUiIn3DU6IAHSE5FPXpLw9peQ0H1TjmbAPAxc8vUyDzJ
8NCGdEmWhTVJW3gVEOqptxVZGIPSyFe22EzwVGxAs9N36YNdAlsMdXigAOIHUhtQ
0LnLAXVrePsnt64blx4eSq3Z3sDH4dShy4umV73En5qdXlU4rWz6DcgxbuBW5lCw
gtPfNkpx7uvpkicNsmSY3YK66FTkfJ5VT6fH2PZJBUDDDc6J176lfcCxICTCGYlC
65u0DEfeQC088zJPtP2Z9BptjLvZdXAzaPgnj5Oxa4MIw7LmlHbItgmA6I00Iszc
zDZNjDeGvKD50Zmx2I38HVbegkrScQT3ruy8vUSgUEHqEvH25B8bCDCCC2+1Z+MM
G6ROv+7FGq3qtWhXqUsCAbdJcIdQgfijaKi1BuEeTnBVaazCL3CeT6s271cpJljE
eqfAOpozpWlWsQJWvlpEr9evUcBD4zz5hsnYDkcdQw04qPPlDffqQYvzqDAymaJg
sDWiZBaPmlF7hxigJpeitvC+IjrPnwTsC5t+i+jBVH5gLRs7eOHXABBagn2a8AZa
jIYE67wF9DlWI7IFxgg1y/UtzbARFGvsha30TeQDTi3S97lXTqjrQp6RgPTynSGV
odLY1TrX3b5TsUlokrmzLuBWxMHRgj+77NVIqCWEglHK0Z0HsBPUURWhh/hNEntE
5qQ9xkkAKhNuaMPYaqefD1c4O8y8fgpvmvArs91ySBpSwfdv87wqKbJuE/bRK7+D
11BFHtS5ZA4PkhdNTQvOpujvaVM6k7ac3JNG2wkBqibRVx3AD1VMTe6Fqf+mckNI
1ESrpBPku3emZjU/oK07mldER+mmCwGFGrttGqiFwoujMR0rGTkylTUbnUWt48uj
/lqBh0zZWmTEggVZBae1kVLVsXqZDx0G+2IHrsc4LD54U2uHeemcMmZEk8XaMFm0
jBmiOHUIhrkECxBxyMS0AI4ikL5Brz9gXLuTc8GB2pakvc06McC51rLuJaiNHqMo
c+BvxwvNxlBcH3kWXkfVACT8yuAeM1+mwcIqXyr1p4EbdkJTKbfhHSeHKb3zXXqo
NYG0UPFXTbT7doQ8/4TIRac0FGS+ivRXOtqMz5Jc0+LxLwn4gO/JEN5dQI2pB7KT
qeLvtxPsYLZdR+RdkmM9Q7/0/0LE0zD1MWeihT1wdBEDzRhVUic3C1TibAyWq8os
lmYbKDAu2qt02sB9tX4xf2wuQ/a9tjMJfvhFACvM2k+kl0sgqkLuslruUh9pSA3D
TExOPZoxyWqSd3Ex4qoronkNE5yWXCoXBXd/TVToRP9MXubOyzrDDFwvs5p8R1xl
tQULXcdYaT4FFgIBwvqProVdPxjhdrqDcirULgA9VCGg9xdQEkgaOqkRw4dioKht
n2OSl65egKQz5CGTskUzyJ9mRyjzhaCckPeBuvGlVt+jMf6LS44oyc4nJNzh/S45
SX4NQDLMJdc2/gnphxcQnixm/mUwVprsf0f6v0YBGjjPI7OP+jGOsWIN7KI+6pTA
OaQt9x0JfmAnu2AQz0pwGcOsujbwNlxLpaWXMZxtHKS2dNZNHlAPYb/RNNEzV7pk
Y6+pYr6pwS8XnNBTUNti7/oPGw17myQNNw7tDSZXFaQXr3ws8wULiePw8t5UMov6
aqpYtyu7Axu8rsz2tGfimL+u5pipW7msjQfJ5MJ0arKOMv4yS+tPskHsDCTxq1fC
L5fv8SRRK5YldcwjaE2NLMuMFshyesT5C7MfN1CY2fvDAJW+WueDb+zXYXl+sQ99
I+AwOE7z2/D5QvglYND8cfaRKe8odC3q0pXR9qHHVBB2mVdwvZSsMcihBlbudLFl
lCh+nGSKyS+xIM4RE2SvSHd3frqIzyq/lZcP+aB0ySCS25FKCXUrLcZzgueuC2On
vTAZFbmzP33kZvWmHvZ6SvQo4QvSErZc9siFtskGBsWNbQXIu4AgfPZtiykk6S7n
Rnp1ZXmFphh16ThdZnbf6isNcJgHYt3dTqycGwDBbiq0mlhtzIQVaXufISxZzWJx
AtdGTgIkNbISsZ49HYFdSKRuIN/yFIs2iNcxnR3y4ZVFAxtjwOhRpg+u/yOM5Pa3
WqUHYUlwB25SZ+veZd+UmuKN46am50IWbEukf25XdqkhjpZyhMjnx4C4E/E6cry8
/1UvRX7JxtO4FcMjnGDISaupeE2tIzfZcrntaP6B7n27sn/BxlRxDWntXVIpRZDX
a+rcGdqY3DImdSueCONKTXq10s6OmMfJZLxFj+mumhgzTwBLsd3Dw+Kf1KxTe5SZ
GtItmPhJl0wsXgZvrMXYPxx3H6hE+N/OUyY8LnKkPrhLo3znUKxjIQSquk/uGNcL
J6lQ4DP3mW9D6La/2CRVk0DHGK3H9HUVfVCFAr34W3ScfGwamH4d3wpknIg5toyT
9+1nns+oU7gsxQgN5ge5NoVsQjip1TGJIuab99k/0OeVcyF9+oRtAwwVZ2vYP5mH
VBWUMtJxtRQAZ9J7oajNU4zVcwVmLgE3tzHzxYOdlLfCqfokga2yOxICowB2b9Kn
K9Fru+u1w1iqgdjGd8oxqve1OgJbOhVaNmNrEzWhtWt2ekKxpeHmm2Cg1pnauSOE
j9wlviA6Ld3ZSNNYFgOO8Pv1cAKYhl2OPG5hWkV5EibrKmB16FYZiOioMB9lU1TF
y5tB+gYyLQ6W2U3ETcp/vRH97gMYpkdo21KUPumGFOzJyIiqSP7CYosUUZIEj8LR
rsEhxswCenT1EJlYfskE2qIYaEze+8Q/Bc2KvVdKtAPro13KpTJVuK/bvrIWgNzv
FHCZYXaF6GilvnExl8FN/ECwevGAX34b/mJa2B4fq6gw7xzz1XrEc/mQU/X26jnx
MEbvuMWWkwdjl+Qfnq4+ph91V5K0D43aTrhuQu9Z2BiSTvscPF7X9Ai6w2Y38eJt
eKx86ZxOngdF+gMxOFvpkjrdx8gm4OnekSJUbr4wr8GqZNEvqJ132xJ3qP4NoSZN
hphcoLb/pJFyFNf37aefuqvtmEDuh5LpHPUIT4SI60gR35qw7XEhlOuKrYYSgWhu
ISXi8/D2ALTI1vbpCCsz7cAj4DK1GqKUv9trKgoDrX3WyTuUCYNl7KT7+CRxjxyW
jzx9rJKqoIY+2QrgqvNRaLZFykkujpEY5Iai4kTjJR4F/+9A7QaaLbI3scYu80OB
PNx0s0yHFcUYnuIEXwXtcNQQKsoWM+3eL1YEa7pTpcbN0nRCxUYEJZKIgn4AOSWt
CJDnOSOxRVC/8W1aVzM+XhmnO5KNa0l2xnjT3QBKnsIXIWuzVnwX74j11weRBdZp
ESmqx9kpDAKOiMrG9XLgIEqVfypiNw3O2eSQnJTjX4Z7CwXjrqENtmtu1U8IvJmv
20r5YDc/AwxkfLtnpZeFmvQBGtXF84DR4VbPZZ319excmhjtcvPPDZ3eLTF/+nuJ
NB9mNfjOlK2ssBRYFZWOYhHT/uUYl5GDVwdC0ycgHz4rCcVKtVtN7UVjRQdknpVn
Ng/5UCRlN/ZUSRy7MP0ZpPiu1mRd91iiahhCH9JIWpPUep/EELsnMN6JNVHW3w+m
8ncvJX09dBX3JH2+7QDQ2mOg01KXHzLLVK0RXeL6d6PbABwiGrrLwqpVpCxKtNb/
ZDOTMa1zYUVMdWT0xRcJ9m/Upeb02luOBlhLkxB8l8Kse+TnglzM+hcMtwNJNGmu
EC+PGc8w+ongqEKCveNXc0Skov+reboU93vw8YLpy7rtOrcVebT/x7YdsnznNDDd
c6AkCngAaJj3Hm0LQmbKsPCoPtKc8edSy49zY3wGM1SkOIeZcR3UWpuoboc3RGxr
NqAGiy3kmjgBkIcX0dYeCu2sp9u99qiR1uHlXBEsS+HsaDB/w/PfgQuYyc00VdwW
xjG3xdaKuZlRfbx+ntGvhF53r9YuiBv17O3I0RK6WiXRg8PT+wmw5396RbayRSvS
YrkMTaa5hIg85g22rBPfQhEfJQ6fxSdV7x4jx8a1QlgFeDdVFQL96Y+faBa9XXXO
AYvEatQYTQSx8e+P2uG2jLy3I0cmITxaPnhZ8alWpqnaprKtZCG3503asun+2ttn
TN535G8xVLtzjo/ZOiT/qbM1aJEozchpVNjDUK1FABIuDgk4MwEGr2EYDjauZOnj
IA7py55QFrxyj55a3yqJPlGPyzA5Kn6vjkVr9v82eK5nZ7rtnWFKS3xsk2iHTTZV
AyVM9X1UTMRshKpvyMfJV+q9xDz03ZFEKRWeccJnGHQzpVvyxmRzbnnADmLtcD6K
9OEFtZA0AHoMZ7oASQQv/RGQnPHOOZE74tYdqjMp70+D807pSu2q+hKdymyNGrHO
IkizhL5CO/EfLeyDgr5CcXqpAZ8LKEHHDEFQsQM8YYdGn3wQPZqnwsrSh0Pswx3R
44ooljVmEQPLASipmWxXa4m74Jrc6ezCjuNXt/cdISRy9hwpwF68W18TXFGHXmuJ
XijaypOTW4aiPM4uZzLvp1oLMbT3u2a6wNuik0ZXZR6VU2ikShkdHONNDgTOIVQS
bPPzT9l6hjMh9fZmVBRCuYWg90kSk3Aary1jp0E//up7Iq4R+Uz5aKDWE3+Gd0Ln
n6NG8pRQjcYmIwmWwwyy6jP4rAnwWzk1H+/pgs1jPm/kBR4JUdfTSl3+Z0Ado43H
nLdwfl8NPt4UxWjeI2xqOoecuxscqfS1LNx6zElDD4SXnFXbHuk9Ff+2e6jCbVYc
MTCy90nqxy82wI1czd0yx3m765Q2W9VD3b67bNKN33EUkBsukFHCpt/siKow0LyD
n5c0OyJsUlEPjaGkJaLdoRFk5GVbkagsdKrlBaiOxDQd8e+aBAG9wczwou+EQLRb
R++LmCBocdpRXg2bZG0RaxGZ4u7XkoYLluPMOSXS3QvVfopdIoxuiDfvQwrgDccC
1kWPHc0vW6oCdpNqpwzXeFbbkpmXNF/h/xA22huNrkJKMM79QBvL5dLbX4NtSWc5
X6/GWvLRa5fybdUGqdQ5ZEcVi8rr/8ssovdP8a1P+Pkj+k4dy1rTYrZMmC9l3U7U
GCT3zM6OelkHSomywYyzCm0ZBLqrLeiKZk3VqxSY/BuWUX9PBAbWd3fNesWxgJws
hFLhH2A1Ox8tNYWH6S2WuS35yrfVHFRPYCo9EHfnxxKFYsRkYvt9BTCqVDCiegKw
7Sb+KrEu6xGTqaXQLsFV983XWUI4srQUGNQMNM51CjrA4OFRRR5Q4aGoWPtCP4B/
cfjW4M7LBa+qF6rnb4HPyffQaxxXRmpMGaCgyM6bOq68QVHgIWYpHqyVOiKxmxK4
8xeQKfI2ZYEM4W0QBiaBEquwtfu9LRYb0ebSVx/UY4TEKwSGgTHVoTOAxtMoH5Zx
9RD3xsyS1FsxqAo5CXe9tXhTqvgfvznfF+WbyvO8Hw9cIIfMidFXiWxbeuSOeHoq
/orP6DEK1qLE3wX85gGaPA0N5SmVAarb/oe9fOOsKcaxa1TW383/lIAcCTlPUgme
qwE7V7GJgySNwQu0fYxPX9cgM9TZYkCkcZE+rA5pV0aIFI8ShVWFHVzZtdkqDcXH
zf082J6HkhhiaksFu9yM0GO6QhAP5D09cxC2VwFTw/pASOG/uOUttKV8QZRzBh51
jW5xexUCy/Kl8p/8+Qk5Ie8VuGFd1XSQMkHHHpiBEjilj49/ZC0lRDyBvtxejXHP
tzJYE8ubqFxR5jhm27JFV77IVGne0lE87ebD6ER76bHZC4rqhlBvY5ZmbtpKpolb
TLXyut0lwAyBO2G61cQ5OAjl55q1+MOTwMvztvGc8mcRskAKylL1VTM+HwyW2HYH
AoPKGmXx6zbc095bc4UAu5Dez6ANbTDLejrPOgvHAM9Z1r/I9D8hQYrgjG5oIObF
6vwncpYqzG4WePO/6XiRZQNeWqbaZws1maRXuwqRT+ju+ksW/kKumFY2qFXnesSo
LZBW+fgEIjctPf7ehJqgn1S5Fdzl4sKWhOg12J72oBzWWZ/MFQgknNUyoIDGHooI
JPEf1Ons4ZUSqA+xAcrmbbznWDEkarnnLidg84H439wv/Ng3oncs05jdrnGnbjQT
MVHQSNzhadNdM4BeeYYsQ4YO2y8EGU3p1Ca8Ldl7bCDJ7W021jF3KVir2FMPcN5g
8q20gBQ7mGOtKqJKVQrFG/jDZWgSY9EIIVOismgS1LBlZKk3Ky6PmW2OkrKu9zeU
EQuP6RmXCyG4zTo83X/BTSgoFkPdpLMgUyjjhMbvACzNBxvjbl2BRSn9mXAsd3PI
nKx4ZTDwqtJs6TMtBUZRf7LCkpTchTmRelKQ/mzx3hgbxtb6Kdnd2jjD1fSmyqPA
X5Wooz31olawbJ0Ioz0dLSgHc25N2wI25qxdnsZyl6iN8EGJBb16C4pwSmBCivuf
ydSEjVmwJGRli80TmoUyZU2JqQgattDdFRMP6fN39579GtSo6lWjDnM1HY6KpiBo
hfalmahfT/jAhGCpdoOUnY/N3+1/5xcQ1IrZ7JdJEr7bC8sF3/QGvCwumgcCfIPi
BjRg0GZ+X3zJGZxYSqszI54ooS+vv1choViCI7srHzBS9KdZpuewinJ/zPBe9W9l
YlGfPiRQhljmvdmYaQXkVZKgCc7MuQab114NztAN7HAVkVx4aVyBhvZoL1RgRRmE
l+fIq89/eKMhB3ZrwoHcc+ghnmzA0OMDEUEc9oMoTP6J6Yf+4HgyjnomuBjWw0Kq
E8G3fKhOuzNWGYPk2FbpEntgOND3KVLyzp2d1pvc+rvJxMYemJpvMA275JIbgRSd
I7dv9L7pkfKTQzmPtNoNvsJuIVjzIqzO7SPYlBTVcFSfBgoNgwYelg+gtUjxNUPJ
WBhZKHRUsW7PCBjzV11G8BgvrM8Fte6tl5u3LqpSv2ueO21XuvJZNrejGIouP0fD
2USk0hm/LBPmtcBfTdOQ9mu4Y3Y9mqBL49KtkJ+1nz3/vPxSIkHtOt0cur52ne9X
QFx5u/IaEbolwsJ4Za8lOTQ/chtF0mDt7E8bxJycdOKWTuNS+2f/mJ002v+hySp4
1D2sTOFtkClh8TWTPJLHy/PxbYo0WA27FGS8YF2k8zPVxc8XdynCFKNZrw8U13Jn
1zcSDqVboL8Mmn9Kq7qHIIuElx3WI/ipWIbrSSNW+Yvle+HJBKslu+M1HESN7EFe
LKPVgyicPA187o/mi9u3+jLZomzXOg6IOI9OxYpRJY1Sud3AVTqsrZXEE9TDQ4VD
vr8IgUUwvkz/ibNxzidCD3vQZPjjvphfMI/CxyBUikjB3Ql9a2xUEVXpiR3OpPkt
z9Z3onLredFrZuifAlVB6NqUzeDoVVdPZDINcQAMjgnfrnEu8+t5u0pDYZVAW+8T
jGl8rdzQvm5+VLQsw7LyDvYFBAq1wqr8c4ZSWNye+LHNK6IH1TO3mWPhzP6tInlm
Jyp9VXyI0lAsoMkFWInM9raylgJ1m1MiveEFot9CKaTL4axmM3wcjMb4jbsSIPb1
BUm2/omxtB/TBj5L8lgEaZSVwyLU6ArBeMlGf7FQoDnEnKGBOGFR7QRnegWT4apC
NAmqOVEKiTkzDRnE4lHmcdB+MUjneCtInCwVTGSBFl+2acN8DG+WaDUDftH9Hfqs
BkxKHRwxXyoSOihyq8KA4LvZFYDIsI5QS7ssE4L6O0kdU/MXXCydag1qT1nwghof
FvyGoOmUzEmLVjBBDyUqIROgTMwJuYWqEO3+DmoxZjOVbL3u8FDT1oT79/R2Ei+P
+WUPhIm1AQsy4/g28kHJ4WpOEpinO/1miZ/R1XIrRR6UJBvtOh5OYsHMxwd8/VLH
UF+J4lPG7+34CcqI+IryniflPGJCAGS2FIPQVFDWtTgKNrhgTcG0QDdjIeVg1vqu
yMmnfL9xzY8UsJO//TFS102fHJ/5cgY5riDNESZv0xFg/usJ+R53X9uMuHHPXuFr
fPDoLLHwEqUagiykcxc95EcO/f28O9ppni8bnSV0+ngGriOAVoU/6jX+q4xpycOR
WtaxIVf+xzGdrYN9RVaN2Jnai5939KC2bMtGC/BmSb4CspBTq6iUN8vGHk78N1OD
aY/Fwkm2lPJeUUsPSRQ49D1A8enkmjQyFUUwYvLJiFnk1LM1Y9Prq5rL4J2ORVWf
g2N4cUL1Sg4gbb3kHAObibcG8L/tIflIbnzTeKPfInS3yi8Q0B6CJ0vDuzdMlWF4
s1IqSEHMhQfrBE5NOqfhNipxQzyMyMEqfu+y8Spo2vjcZZ7DRqjSPM4gKsf7L0qs
dxmx85TvtHYhDifsHP27DlwHPDarmSU13KBDH1vBee4hBt7z9x9xPRMGzjOPd9mS
FnhR7RBmGCK4Xa1tifXzSn4IdF3uDd/b5Iv23clfCP7vThdmodJa88TDQ+pDs0ld
x6erxojV+0oDwVExi/JrsTfxeYNKsroNq9xaPTYSCVu1VrIE6jzk4uxg8NxoreuW
xljZPMaXlTJspKGwBbuBcvj2TT4HGctKvjnNdTIx8srTIEq7BKwloN373hzOSyoH
dON9iHT+YGaj0y9Lv8Jsmr3hY5+k9FqE9BK4UA2/8k95A11X+I/n1KiLezCUJ/R7
v1qaaksd54vqs4lP/09u0p1UTGBddlHGNVgOiPZ8LUlGiq+fu4ec1Ftd9fc5JSSO
SATHVRewfN9pj2zanyyoCmfcF3LPQ10oURNAW04FPfiPW2ymmxDEPKtjAakR7EmZ
F/0yOYTKtf8qc6qBkV+oweIA0uQvO/gKWk4b1GqjKHuKTqFeKLpB4s8837yGYXjt
fTKAjYhaoLj8RPel306K845ZTPNhwpUIiAhW6HRALJVMDUHfYZSxAOiGk/bGJ/Vp
WMCLSXhVjmVnXReLtce7yclj/y45YcptmZQXfFVUoHUFACXGOmgoI2NqwX4BRFR3
SuXb1+/uxYkI9uAGz6FNeU9s8spvIwtKrLl4PXHffzSKbC6+iH4TnLNP/RVnBCTP
r3y6NU2QEwhonJlOgvoBDXBgICZlZhghUJKWBciR/68qjOFeT2Gkr8ERqHG5TODR
5Pg9GH8Cx3ysIxmpY8V/wbXuzqLh/tNWIzB85JwWVv3T72WKsB3HTCb3bzOEEzFF
J5dRPkexOCCa1naZ+e/hgdF48yy8FFXQPKNwjHDvNOy+D7HAIZO1rTULSHdEd0xv
7s0dyvl8oyNfR9T4OPlDGhout4Mn3H8KcxriseVll6sNrbr9K42RCIs0eH9hY1Kh
XE45YYQM4YpX/BYYP+vbKlZgrwmDaqqOTPx/Af8gwbqYXVTy/Wwo5xT3nDjAgy3X
qT/p5R6nl5r0T2XkD293cdRZiK19yGHc+7oqolFfElsCqjfrR4Lg+36jey2uOaeh
4GITUTdM0a6t8IMkziZc46TjeXLZ2UH1CacIVjMHHP2ABjT3rG4FqwshogUE/xIq
P5pp/5mQ3rVV0c7clDxobReJoDD9Sbei+hRJeeZmr7SgPrHbOVj8UbVIWedjGGw5
6rK3k6ToT1FNXFywTFIPRJcO7uqdZLyZuY3iCz4TDGbAPWI0GIFrDjiEzKKuiMYY
yoeJrYuIyvFgxaqst4FNAncTbtZucGV5b+Bk3w3aeUJarxlngi704vIJMCLxCqaz
oPeJDFL2QfuO91nd+IBlHgNJI17xaIAo9pfFCbhlA0u7ttgRPUpoH/mGWla3wPBd
ZhlSHAOOM2ZewX3/QZivBmfOcmV6H1TOZ4b7ukucLonkiw3kmwt0w7QlUqni3hxr
4qP9CcBuB1Tqpqmt15kyTfFK5ZbM+vChXnA1+4BYPJAq+D7tT0qQTEkJiA7UKqVZ
OSBiLCBnaMfGL7A+gfMIWVi3ub30pfea6juBkzTYAuvhXmrWNdgtXillwdAtAGjB
75LnHNj18gzszIZTa4jKqNrdsuVj/QTkW+qK936aITjaazGATiyz+YmneMSfGXyK
pHQLa1twT7IhbTgYdPz2KELHLNjdbh0uRngBoPukBZa+QHAiwVExXR0SUJZXJRkw
rSUTodkT5kfj0BRCsg0UIRDsB5HTdJ2zXSbmYnmh2M12BFMwslXMmhf/Ikbjh7kL
ZlvIL07kgRNq2Folt3q8vzA5ND1V5ju9XDaD6APez80qWeZkR8E4MaLz4e/Obw7T
Id4mq8IKDmgTxkuiDFOnkmf6BuQmcD9YPQ0whsW4KVesb0Aav4PLq2YcXMHOvXZE
MXP7xTMLvv8cXIg7VviIVikTN7BTC2sXEYbrNm06GxMSBC6C/r/y6kdAQS2LhGpu
h0mxghlXig905DdofSdvP58ABHT/Hudfb1qSwkhxpvRj1wpY5e8w3P2pmAoMrNlb
9Yp0siAJJ1tjHZBdpiolcx3RLt0In12F41sSvu/ohz/mQysYdieAc5lG5E2MPe9B
2ZXSM/pp9agO+6BuLbF57o2Lhy3cckBxUrvaUftUVYuedYWI9nExIemWHdzE6EM7
h+gXEnoY+sk6VtquwGjCOsBMA+0XESAj9EcdKjFGVw7xsX1N+DDHA2hmJjGOhezr
OcZoWtggPTObdHA91zbqJu8NLNEKocxjFaie4wG0rzYYI7m0k8QzKatdFC4K01RX
1zWnGBoaek8nGWIJ5GKpOLnafG/nVuui+RiUHq2d6AnEuaYBiDbkTzfQm3qEhsuT
GTcazstPQbL0gUn4MTnrMJ50bd7/EE8mYIjvGKP87eELlOHupe31/wvGQe4m+J61
wKA0l5fp+4m0RlhKDocGIDLxEpLg0fidfcxK1PvxfFHFsBKlKsd0Px4DZB0RQMrn
s81NKMTse74//GxU+GzXddKoEMWGMlXQfxB5qV9nsDeO9RumD/XI0hoHZzobHKiI
8XTZFKGxU6qfY42cwyeeWRp22T9lt0xJRAhViuKJjbD5AK6mCPpVwEaAAYMUCcWM
Nh9hemOsYOzd3yRMRwjMRTx3TE8WYrle9bOG89vMkeJa3aBU6orB9zxnPpfuUyBb
KeTQ1XMbnYNXpD7v3fWCPreCKHnckA/OFoqGGA0DZcA9Tn2WPYatwx8Sfw3gvME3
NhhVSusYNWjw3r/bmIrcu1peTTA/YsrDWEy/1lPq2ycf9bcgEbtIIJt+SFZBq0Te
wVNYwjZtrJnXb0yLG+jqb7VC4s+1HKYjeyoXzBZFMkgxrvNvngEjbe8SP/oqg1L9
bO7/I7culUGe6ichDHbq3ghtLymhf+CWU2LhVK4ANTuHowuLx5HSTOyXJYayjEA7
6bbw48HEZ1+Sk4k3dfPXAMq86Kr64KNyXck7VZNN0e1UJrF4ufy+BAE79r8wcY4y
l5ZllhItxauVxraWUNpXN86jyKt3uOIAUY+GzhOD+f2RLmDrcFoagSDsyx7kUBjK
mWqruaDcaq3qnykA6HzP/FA/HzXhqW45iXFNPABEnoTvNAgDe8EWh48m9oHJOp+L
GzJ9eQbH3gSe0+NmAPrJo6RL/aAvIWRGKa31bW9Oua5pyvphN0s9ZgkVISQlzsM7
b4iv/P1JFBu/3bRetr25fJrJye1xSmQH6qpUoel+TC8Fcr8u0WeRtzhk4J0wqGAZ
1Csot9PVmkXVV2KeMMBiWkE1MGo396sNDwbR8c8lbolNlbThMmepMhyxwktLJzXH
3LbOsW9vxETA2/35tg53B+G7Kt1iqr0KxTwihVUQTQC8ErydNU26C9JgodjnQ7bY
W7VdDBcaNmeaWhaYB8QGP1m6rCwVnG27jriu3CAhb17+fSwCu9OdtnvFnA4W/Wi7
vbQMdDl4w5IhfcQNZEwt4Vq1q3pOTvgHqDmNogKbUwG7KUZw6Ay9RaQoHQNsKWqH
EOjykC0djeRtFzuHTBiY8L1oFHnP78m/Jk8Ve3PE+oz8MCi0oDFwUjy9lhU1m0J5
ednad2tU4XXRfC3CpLFtkHRblpjYxO0sMoaia8BenxH0ybeTfCsZ/g9n9QZAkGxc
u87eslBL2gDYhfLaOuYfehW1GNQoJwsc7VNOxCEfMf4qiXtrvN9CZ4SNJgPaT4Q/
AGOrourVEmjRJNdvCM7rPM0lnlYhmSpyFYlb+tzGcwmL79LM3bhkn52IoWiPjjvJ
c6M8pmh6sQlXYwfuRE3jV7jwU6L4ZPzw15olFGGQoBLwRpyLkOLdYEfqtmGybRSF
LSCSpyNNS7fANibqBP2kw5Ebm6tnEpNhycXxtkjNkM3zL4QeOumEoseHRilVIWzE
yspuJqUD81IIcA8K3GWsj9OE8Fhq/62RApImuToi3FmdagmD4SXa+l5gCf147Mom
eWRbflb/f6NfbN6sAeJKnGfd69NvwQ7rOnymI4K0c6WEGhRXfdu86HDd2l8Nzq4Y
wNXwQI4B95mbMboSTnuYRCaj3Ki0AZZbazPygWgeI0M0ua+PUZh4rFbX4Lm4SGOz
GwKrF1CDE7TkRGvNfW/gIIqLSrSHZNEt3Dh5SuVBiNkpkDHX7o3cM2kO5QUrkoBM
F3WTCgwaYHtiF4HsFV+eFxIIu9KnI9Zk+sBQLSkQJDBwd94PcakpxasafJeUj4Ou
VEYEXoIZKkxBFWoF7bzz3tO1zx+lhrLGYglr5abZpURVOU81Qg8iids8/xilPB8B
38rHtmb5+EP7kjaJ8LoKXvlLymVyvlY3i1oHg+FTS0kzjq+izljPKOMIDo+rvwzf
wQhI3msi5pMWxibTqst8EfAY7tx0XUR3PuZNONxiLzHU7Mq6d0eTG/DmzaJdAO87
GDOVzu30aJX5y7VapS6q3FHNN9htX5PlJt+LY306mSX1TT0QVqIpVa1wtEnwkTIY
dGZMz86PpUWFUFSoXW3DgRGXqZOr+RZ1iYndN9bbTz2Wsmd2kEjgXogPI1ihBLqY
nxSqrsh/qKes3Qi4ZfodGEK6mI0sXAe49YAMhjdejTpU/iCzlTEM67x9130Wi7Tp
jYvxy12kPv1cdFdfdGQ/safTFtW+/se3A96omyXyGQqgwRo3m++d3d4wu4cbvvki
l6iNDCl7Ev+zp5Z9mfAjQQYWmu6w9JNneNmjAYQZhVbbAmLq6m446xZurWJRobMv
A0tL76Iudyr5zu/9Mm9ome0JA2jPygRJFjZrwF1pX1mWAyhmjeXDbSORtmV0G1Rn
mZWcSsegR7O9LnXVXN5hGp/uWIdEFbTOriPGta8Lwy5hF/lf9XyW7pd5i8U6JEVw
HK39ha0NMeqT9S2sonkZI+73SCWoGZKuci6KMl82eQL3OGtUFORoP1/YFrSCHZ2G
Hz9pVgyJkxtkIbOzb87TR8Kj52t6NdVQgsRH3Vxia7hdOk99TF3pkPmiUd5kbtnU
vtOWdUhz282vpmQb2LL1iEd3l2apeFeUVqzv0N+VP87XpUfdKUzP1lpbcbNDRPFe
KsQshG8GUiRxNYByxYtjK4lE8oS43sMq82+BlHnQkv7B5X3U396Morc4i77oBB66
sAJWSUf80hEFteHjWmWIooNvlCQ2hXVjZaF3oOJOv/TfGhtiIaU7frBcSHRBHUVP
8eIYJRzkOHJe4uLMef3FpG6sHtcH+0YAtGyK2XmsFJbUEq5evdVQbWFD3vE+6w0a
YpMa5G7GYSLrsMPQ7+DQ2XtYMlVoSneYY7oVP/JBnWxTUNBWPIeFg2uDZWuGtv3R
JX4ZaAfDpfxPO8d67iQP97f9e6mluWbkmVerH4ytRjFHAG3bIfDm/9iy7Vd30e/p
tkX/oOvD4j2lP6dLd/H+yvPHEQtSDYowfghUiV/fLYN40Slmg9pYHxeLP04I+cq7
Vv6eEfgL+u7PmbgVjs5g8Q17LQArp+bQlesVumedjG9w7TLjWCi4IOZtt7C/b+nh
a3YrEyg+1/aDgaG4IMWvIhME+NViCJuT5F2fRJZTivfbnA6Zh/ZDBC+xmeq6JzwU
6JBiVtf6SKUZ0Q+ARh9ZhtcEzzQXhuAtHsLUnX2E3NSjfTZUWteVbcKKqAq+NUCb
DMAkWkAlSKEQdiZybwsNtrlNlaC56ChBNHYGWuYXdMVpKcPRbdnlV5yxbwHKYMx4
5waah5nSerJv4KiFuNNrXWqJLSUZJoV2honzxdrLiSbykbXHpqql2SBbpgR0qpVr
KfKhHoksC3sRHbllhlTIX+hTGiIOK5tEKsKk4qAbkl3UEbFtH1eNM5CGPlm00vyo
rZJCntvpo8en0Ctu3CnB6r6kHdDlBmjqdhrTX4XfQV752qaxizEYOLYk7eKs2LIb
lXcJRHlYbaiv8S/SNM2kDhkfdpENaUSi9ulfoxq3y/EIRnZz3eK7aeOwb+/FPv51
RDXACFX5nAWDncupA8Rj6jjcnuR5oKbQp4QlSZQdA/x69jYrF/INnsAOQ+WVYSo0
W8TmeHtN8h9TbLoWeyFJjfuLKSWfn0vG0vXk1RcB1cD/Ak0jNfXi5JB9ofIDbi3i
L4X0bkc0XhjeVe4fH/Kp1ToYsT1uSaPv7h2jXBgevuFrd5JV0Dl/4NuyCTMtWIwJ
QVYgDUFpjiYhruPOaZfulnPvaQYulMqHbyTDTE+zv9QaWfCt07/lzUMej/x6Ez5t
uxQKxC/h6Qwx8AgPvYEKNikS/NwXMdNfpbujTLov5aiv1Oh4yXqXGAm+aHi9nUQ9
EP/nyT+wlsyYND8xSQ1aKASAvSCB1vuDUFO6fbH6h/r2vS8cneClhWlrEzxcm/KU
epHD/BybENWdGaWGNnLUZJR4fDd92k8GvTwpFVPEIG/EQTbfht2c7qnqdCn86OM6
ibL49P1wq+xagCyL6NJvD+y2GhSrixrIXDYRbYVw59chRVoajf9djsOnvxoOh5NC
JQBVPgjh3/L+py0EYUNqfTq7wYqdCRtRGrZipMQwGRlpKIgcHtzupaeN95WhoW/O
dtyfwtXLocJURyh1bWCYrgalYwgEISpjrbhNPA+UlChSSXfTP7IhXoydkN5xTOjo
rwip+5RzJPef8jXkvd5fN/oB01OK/HlOiFG/OXJdzIA54yu3KBFLYEiyRd6ZvYZt
WN9+90MQoqdZhoYHH+bf98mntPICaZbLVO/YzBp5Q8cqOpi8Rw4hbM0D0neTtknN
D7AFQtLIbZsi/fYT8tIHLzgAs1DYIIvZfaG1gbK6rVGyhwt9Z8+DPfTBXcna2X2M
BdDEnMKrk1MgSReXfR8KgYtBhh/9hznfDLv7gVOmJviTbQwiKTTjC2t6QdX0yFxv
/HWWV4pE90xok3nq8LzJioJIMelKBcBOTW6OUHFsQWRFvFECsvwb6nEOcSNJsXcM
Rm6LLcIT15e4DSKN3uDKKy0GHUQd1d4U89gOy5x8gLuVgm3Q2fT2cOrDFaRtQccs
sYmMWObSkqjcluSwi7vnjEOYuNOkODzg3SlxxRxlTeYgz6MK7e1iAAgoYUMEiisX
zsOA0dz8eNvk4d+3IxNrIcOmJAbbypSv3Xp38UTik3sDvxQP1grEL1hUBjdNQksF
AxMpM/rS9qs5HLaPcsvrFL/bl1lMxSUaibJYhW4FzXkF2EiVzd0K+JhgkopcA17S
LENZoJvY44JV/JgoYq6iZBG3sfP82H+sCq0bAyXGkBYpqY+LpV9gi2IVDuXAJliq
fYma+VqKdcUW5i/WLhSuPMIZaDAsN4LRhEbVytRlI+SjX5zW+LJ4HVB0QFfCjX1o
k39iRLuy1u+g8JdA0Jqedd2uQYdr0Av3tzyX571lhtokeMHK6WeTQeKHNjvWRCq5
QaoXE71/qeH/Nkl1mBpBMUl4EZjT1EP0/a6l0iDrGj7g2yT5I09d5y94v1Q6WOXk
SwBGdaMrXodH8w4CGyopYnn32qU1PjE9/CFYw7OsJBMm4jzefM5bp2+9OZWPZZ+t
fQQZNeKcSLiigFwHT/e5VSQwIcsDhvO8l4qw8qj+abzhYFd9QhF3HVYnS302M409
VBEymMB5VsB/wHdPJOk/y2OVgwCvvVxAbtudCvvAiooHWlVdR+kRWz9tKcwnFkn5
zcY001PQdagCus6thih6u+fcQV9OzLJeknqfAPGw6SFVEQv+iDiTqCHaPFaswBE5
AqnDUHv1WuECkNOrxEX7X3KlO7AuP1apEHbQkzfty7uGluJDlmFtFSz2vz++UTFi
dffEiS4xVj5CAZBsfEkxPpWzNKcRlwed8GyXKoWjyh7/ZOPMav9l5j4DMA4ZmoQA
ZRf4UTkz+JRslLEtgj3sO8l2VNFYc5yTVIbwvtdNNoeKmnIVbN2AjzozRmCBrAlv
2FVNGQ/M/tANJBRx+kYs/vrKDP+xNBsdx+m63h2z1cvnHHnvv4I1gFRAwE82j33q
UTqJyZG5RVlI6w53xQGeXliuqgZWmW7X0uqZdsO1j/J8vxYyB+lO0lFuhER4oA6x
9rsH+g96KDTw6QtApvbQ0rts8EjgFHznIRu1d0GSJn5HrGPC+c9DV2P/Pgwky9sC
X+pGUkP9URUpMnaVk/FNngsHZHQ1Z6OgDaaFgOlUu/vf/CQaS9kWAtGLOsu93oAU
sEW1gb/sx0FW+NiCc2mg/PFEOHlmMoJtKKI67psWbulv0y0KQkXTgK1AKALPHiWl
aez/4PsYaNCMvCwsaKgTZv4x0Y5FtCYFo5qS+ySDCDeVxok36i/FcjBbyovf53sG
5SqSHKHt6s9TtSD3Q0LzK8qsTz3pDWgtZhNbSolX5gclxCBNdnkdx87suqa9PnV7
3uYqg9JeCANzDDLzZGc2jp6dXeNP45n8yTW30elMEqJmYFFohgCpTEx8Iew5kF5b
gwEWo1FNaZJdOR484KihDZDjCHzHayme9q9rrtNlgo0wZgOq6yTHvSNK1b7P6G/x
LjIFOpPMe526itEUSYWnHzxMLbLXq9Z7AJWVUm+5Yh1QUoBeZ054v8+PKlJ0HPTF
2EqIWLn958CNjOiIo9J9C6Qx9+HMgSBd9JkESAKN0wnARPHUU6NlOSEXDq+LOE4S
7E0WSWms8yS0K1BI9Q65YCWz2NeJIm6CjCxodpAciPNwG7t04EuLBTvGJJfy5+ww
KP2Jz7qDYO2aTkCki7iOLqOk0bh3qKbxq0uHkl2ERJ/il1o0bShsNMSpfem2h+uO
46SPt/m9S5e2jktmlWlmrUJRfKn2YAEkJ7aqXSXdHMASxfyKqUj3IaDGi2DBqxiO
+44AsGZIFiuDqwHMnX+1lddTClLsaFGaxGC+M4A/bk05Dzxtz3SlG4vvF1k2zYQY
n0DZzgb+KHPiuRMfs9ipIRk09vjU+q2oEcwK1woqa+XBCVY3YCGDFMhHtn8oM4gI
kfyNabagE1L8qAtaKePysdhvOzy4o2Wu5zAsxZjv73qEv559oUGNcsORy12SsSNn
NMKfSyzdvQFhkBLVAeDthrbAgaE9rI4nCP4ORAR6YTQf/YHpW49eywsVFRfZSJ97
J+Q4Q6vx/cjdLBigstbloOW1fWd0HpDVaJsfGyWpLP0+4UVoNtSgz87MqJQRZI86
4aDrb7c/38M/WiDtJfy9F/1IVXvsQARIpN+2ZmuEf5V5ZJHYooKf1FR1yiXYVEen
fVyqDrqnwU96uZnITTyjXuFsQy66DC55il3M1RvxrLGe7QObuJwiuY7Y8dpBxrqh
UCedBx+N7pqNRNklnstpyu8LMQ6GdvtX2cn64DgmxvOk+0oSTOfOpModGIR4xlX7
9iiS5P3qQElAxP9Wja0Ktr42/28rLNuJuPHtKeWHvgXnYsI/Q/ZEiqRFbrZs4jI1
JLT+vJdgCxEAqcm+85fGvP9Lz6Mrv9zlf2Oa9jCJfIVN8RChKmD9dyCdzcrWazg6
YhH+eDcT3QD3Harx5gCzI/yoxOoIFHm1lKFpcjGF2k0KssLEW7OZzozxhWzQbAg3
cMfSRkWZPjSFdLAg8CgLUFdHLGD85U1Mows3TS6MJC+b1COPV4stQUd+xS8pY5vo
Pa5xJW0TXZQDDesZ6JE3VgMoT9XV+eAQN5zyjl0pQeNpiQRtvfcdmmr3E34D8CEn
WqN3AjHgYh0NLIEdn/fukzY9agjLd6COLaFLAlTACxSG5r7NXYLai0Xvj2g2VGuq
rpNPHj8rqPb8NJZaBAkcJGeW52Oa6EgaglMUugDrLZ+ODZcfI+XSFlHVoIQGTiPc
jvPGQXJmGFVpXj1pK+B2IzI+wLc6x3MxOBR/s/jIj4v2X1UzjScaJWyTW+3yH1mS
eZekgv4oOqHWIYLs8w6++f47KyqRFGYDXoy0oBswOXgMpyZS4IQmcepyJ7hKOlkZ
abiLX7nHq2PIBeqMgn12grzNLEbj9oDWx2W9xzDz/U46GicbL1lnfEgw4JGMYo5l
9PTh7QD4pRTw8/vE0XNvVoFiuoUDK6LOe8U4c61ZDAnGE8VT4woTB55y2znsXF5F
ZCYYaPwXXW+kNegij16FCsR5xQTBbaae6vFONubfIFDqf8Dy0cbAkPtmdA1XY0FX
Wga0Qu3OFZMSJz2G7MM1p9kC16eEa4OElIvckVvstzj2ctcKWx2JbfcRo6q2W6KD
mYP32Hsla93TvEXSbreegCvUWGtkJsitK35mF4NeZQY5QPHRFULY4LLolbhu1/Qj
TJarEUKqmgKcd9rvSQENb7FcxeQJlJJUFn2yvv2X/0mR7b1TaqbRp5XkSrLmgCOR
AlBCOesdo8ehfhUHe5jEWGmOyb9vY0tztA64qzSwucZf/bmlD9wR9RVLKf0BtItf
7C4ww/hurRu15C5etxuLZLz0zzNE0NfLrZ4rX8EBx8ySmd+OtJwvZ1hdwNA6pOa3
L3k3qEm1GISJiy6OFbg/WJZf5Mw92bgoa8b1L6WH8pr+G0qnVoQSb+amLB/a/wEf
Coe18fhq23i2/lraWc9Tjnjqh1XzToolDW5JxQYy5l3DcuWkIS95MbE1Y+7qIAf0
UF/rIT1ptQj23g3Dn5pJIs4wkrUbiHB7j6QUgXiBKjPEl65VcWr2AfgbK4tnsvSL
ey2NpYJZLduaxpWqotLPDiHqMuefSCIkxo1JNddRjVSN66OlL6NCtOANa0y2cXg2
QPSAuSCrv3Wv1x4QGrOw+6Z82K8PkCKkQMBvmO9gn5Ps19LwtjDNeCO8t/SQiaD1
OuOMt+DH/3YmBYmB2AgEu5Sgv9utR4wk4Ufv9vT7yZ28+bnRMl5RlIdUv+A9gRsm
YxxkOz8suf7kYI2G5vTDS9/WVN092fnPipxkw+udJb/0+saGMHdah9wXzQkXg1nQ
OanrIBW7RjtsLpdbqkit2kar0HheGYS7r3saw41ZfrcE2Zvedz6hEzKGbQm3v07X
O+dsCjo0KSRUx2oQbcYW/3K4Vfu9IBi8scAK69bTbBy9KXyWRfugQ5ejk4886pwr
rUw5x3GPuZ/o8iwCNFSUNJTy9ogMPKl1pJq71OWSRJJJBLg1M/D5/mOnQSeCHO5A
nuyld6z9KrTwM6QkzkrgXAk+j5dCFeiweKjlpaC9C94D3t2K3fEdKVqEGuz57K3s
YOFAu5ELPBgV9ZsUzNJn58ji7jCHxfJndOejR8pXkTIxJuKIWGDKi67MFWxtjMd0
YS7I5k780qSuTpc6POs2wSsYmmfdvv9PHXR76mVhVpNV0PlVHEpVv7ExEAUis+eU
aZvu0NqI/DKTM5gK9/4chPh+AZ5Lo2SZ7oriT6djoUqm2uir7UdZqQW2E4CklxXD
gxq0Vfm50Oycp0dlxbDleUUE09z7SY1Q8ENXHrdOWpuxjqX6Iv/1XUHX4ESdRlUH
+TMpxF3XTl0IylhHfF4ebZwW5GvM+oi3VDAEYTJc4Ek9td1oeFRHB3xZ8MugCRj2
a/dnWqdK5ywK53mQRRh1mUHtejyMj4LCeRYeP7q8Vhf/PSFVUNzIKCB4ky9nDqzP
mFUt8H/Xe6+ZsTHWBomkj9fZTVZWu1TYIMi5K0KkrfTB75ISazIx/8ywY9SvH6rz
euBlUjvp0S0zFLuwDdnudaAbsmVtL/aqem4O+kjOay9svedxNUvJ3xTUMEbeL0Sc
fvvIEV/+od4zxg55iBe5aL7w47D6nSFkVNmwGGwTYGEljbieBLXWzshXxoz19A+e
MyskhhSkCjHsK9TXNITFizu7GrNb10qDxzVxXK85cynp7wPPqcViCLpGvMMYdm7T
YXFxLe3AVoSE5YnT96c8pQaFSt1isz+dStCZPXoNEx0QAcJwN0GGYygXgh6puDgv
o+/VL25ck3XZkYWkPYh8g6N3CSohqsfS5cdp30Te5uGg0uYImf47cFOlC2Dkz79W
spYrHkCAvwRoYrBYaVAAU/gLaPwf0e6BOMB5coV0db6S1oTMnVZK/bvC2lQ5UYnt
MRJDpRDbw1bbBQQM0hYZv7W0SLyXSH+EdN5DZUQqt5NqU8vU1W4QJGa/MwoSwHEb
vKM4WaNCcVHxroxROLKOK6KyhEwMIdEMyk7e7M90h46Fx7fQMjnk9cIOg2qxeYQ3
pcunuPpAcLdtZ5XJxdV3ib41nMaC1pQOT9pGzhfsDAESpMec9v4DPkeQKnsSpidn
Q/XSQpMqPGaUqb6/eDBJmWNAf3QIN4BNhPxiKpAkoXGkXoEuXJzC3wB3GAWAZy1b
bojNI8b5BZTSNbyiDpQcSD0HVQaUm5dF+nsFx5yWsdvbybEApb6JbE8Lrd3mgaJP
pZrjYgOLu6H5v18vpLVbVk9g95ydW8H6B6CNR18z0jljPb7D5VGTbBHXOsaKToWM
Kq8lSta5JzcNQEIHnnpxG8a9gTDcCbj58MzVlRnnkRtfD7uvFCL6D3etWdvQScSG
hwPqr+QJ8AneEa8P2IHFuiAYHPcl7zJMTyUnGJiBxBGEjSCvcz46nYkxYCYMg5s1
bauDxv1j7hzBe4rNQmr4lx1gLjbGFu2/mEhTySBdM4WxcjHbL+pZLKV1EsikqPem
1GagrabZLdKD0AsugCkPn+5R4hGjLMfOkC4/OS5ItEuJpdus6Gmmil6rvVCeH4gE
0L8lra6638XqKPpUEB6DLLxwxtOQieQxlg01U7HgBVnLUMp0c8Z7QJbU0FQ6Hzpi
FDHgLIfcwF3ZztzbJOLtoSdAqZgUx+Quti8hYCY6P5nFHSNoN7fQx0LCcfYom0Om
qD692w6Gv0knQfCB+LkAwSTe+MWm0ExhCSinohXtpVOvgA1+1Fz7iCR4G8JdOwLO
g6QC/F8VNNke3HXfY/6wESmvi0hToqHtJiRf1c/N/WtVK1/FyEorcbEiJKxyLN0W
q/19ZfufeMI+SqJhw4ZQgiygg8lP1fL1ZqCNRS8mSofOwcvpKNEc+CXhQgoZW+U7
sBFjWBPg7ieHMM1IMG742dLHJxrhRxpa8Sq7UkSzmE/sd4l5tqatEMHdyXkbDCa3
oP3yT1ch4biF4XgQIq9N6WDrnjnlrDTXmKiDUeMI3mF2Vs1U6QTGoXA8OyBRNWI7
8SIU9hDR4snXx5YZV7NdJglaOEMJaKXFmsoDLuCHFq2y995VM8nRaKz3po4/HiD5
zxgQQWe8RVKdCzeg7kUUpb54u4UU5CHwgrafdvRdAwj3iQpBk5YI3mGrbwVyHs2M
C5p98mvQfRfRHEULaur+xwfK/roHFoAYCmleIMldFqxjzCEvpBr49mQTAGcs/qlG
FnSG4goHnCJgQBCI9BbtlwTZGk1zJVI53gD9apj4eb1v7kdEYbKkRQ/lRhCXemI/
OWXCkYI5ufqpZ2Za+wW55Hu+lYnXd7AY4yA0rLlfyNQ7jA+5iqgkv4H+yIeBLX2m
NwUx0lhcuzoYb3dWLMqjKnBYVkTjVCqRYFC5g4Z/1s9cBcIentLDDndSoUsDi5Jh
2sITyXPmfarAlqnIDPVfKkd+v9TPo3897aprDImzGsik4Hta1UzzeFH/qYCS9//b
z1iKXsbk3waKzIeEKFj5behQ+PHcO5nHUJ7dExh3bWSzXNKJQhwhGiWQ6V6/S+gK
sM/kGy+4Vee6QremnXazolgxvbHGcvVm0C8PjIfpvf942/7VGPNjw830VF0vECJZ
wGrkCgQeYVQFOOqSrYspGbZLuZuQVovWON7pHxKPrWvJchlDGSoYIewo6OAoe68u
8smUCy4K1J+YIxcWKFtJY1WV3/gveCf9yjsj0SNLHES8cfdycfAyTqY9E/1rGNbE
Oa2FYLzbo/TqYyOELKU1Xv6+J41Cb9ewOcb6yg5G0FdJU4zn7IDUItBMcNfViXcD
tE+KubOEg/0nioQjizUD2zlSpkg8033yWyQwAE0gzgH+laorkgKUXss1q5nxPfYp
dgosXdwm+9EvNLDX198pQX0LWwyp1ILtK63PTyKlLU9x5gRg2Rc/cauTRjRwYyCQ
UXi6kfT2iHWsFFlpJTmmwCTwJ8p9d7hvXh9MnvC+qyLsKFyaI0Oo+Glqfc8pBpXh
9RwaJqEwc7/rdPvH3CdiJm9EB3IYLpoO8Iue8uivN/SwftayjSVrquSBdy8J/BUo
UCINaTDsEaFz8UiAVK6GHUvaF65QxgigqmzTl1D2VDItglkP7+Im/f7RhKqH/HYY
XoUA1Y61ohAlCUdElcgBIvz5ZxzUr6jBq9Sc+XhY4Ex2MTahXWrdNDfHAxUbl86M
KsHNUwl8e2v1ZSxLTzNwZHbUTMTZqoX3udiU+DpI9HTDRcQFKfoVy/DWcxzFHiFc
qYi29BtGTN6IqXycpPJwid9gLJvmhn8TJsFapV8BnSHmTb0Mt77NsPxKK8xcxm+1
f30KhHfA0eyFi+gFcAxQATpdIOwEfLlxWYxauTLUPVOyskcQ2jpRsKlia4m7/kRJ
/DJld1arQrZmr6us5bO8JEwcWtWxVZgswkc5JwtleYFl36oqMSKMvoZbmgtgA17u
IJLE21+ukdxeAOP82b0fgTzNY8agV3D9FAzPQ+LHHQUAxqJ1KVn8UAc/dmTrvmYJ
SJ9az8C31nVnpsufuX6A3utbb5K8jHvbK2aN6c+ROfpIIn+PmtVhd1Q8nNxdfiyF
MowrVrCoRJrFovfMiiRpErLMq1iAwohPwrEy4e+5uEVoYWOytFNJrJ/IETGSacyd
HoBXqlPcR04rN3LbEnyCnMlatS0NkkcrS+gNtrhO4V/OEb9y46H3KJan2QxKDAFu
0qmq6WM1xhiLd5e+NsmaPg79QCEc5opt28CYOqY5U4u6ThK2cer84QXGk/BEV3A9
d9r48UIzb3KjRzu+iKgMnaZCams4c4hAdjunliAwcxoGFYWw2nQJoJ+wBQ8PPwtr
wTymNlTCTlc+WdmRRLmZBwI5NvesQdztNVr2QU7DqmEWShLRwnoV3hw4oEJUrG7u
ytRs0UCrAgrY0jgGvxAvfIpknBtgZH36lcUBQ1MRNTpOSSaDwZvWztQqvnqJAXNt
GnP7u7gwzCY5Ol5lQ/d+IyfMJZvVUuGRPObefe1mZmA9F/qDGVoPEQfJKIiBY3dU
xMywwZ1FQURm1mHJvocpA0oxasUE9jUAKfLfx9GCWqL/aXFOL/jZJ2N6dqFbVxSs
hbsXqXAYZs+IPAUXhYikbgowu0Qqe6gUEHGyTNUt8qHuZQRz2j2+lomGFdQU54Sk
1t04p8GUMCIyK+Wy69x1uX8wghzMLC1oYWiaLu7w9ak7SGOZDJBPAKy8DiZnZjMq
Xa6h7TyDpltk7FP1PJE+DRMb/t+Az/7Ez7w2JBQZUFDc6LEp8IFaqHQrjQ71Lp6Y
FjbNjN+7nOvODVY4gwhtf0hRHBPMrafXWwsXg4CLrcT8qe1YNM9zDal3CvY8baVc
Q60sa9Y9zjNvP8JafucWGN81Sfm9TGuPMuL6dZDXquE5bSqE+IRPE+JGmHn+XerV
ge5M6QoN+ZB9I2xMrcQm8qRe4Bt/Ft3SEoSCfGxs1uZAO5uc8I8w6J3B3mNj/AmB
I6JnOm+Wzc8p2kmmw/RX/sPNhug/QF38TXdRkdau6Ovj7/jkT7UNw9fEDL1K+PU2
VXh9BAMLq+mH/XLCLlS0zq1BCHysANxr15yxYojmBHd4rgNg4Ac0ncSHBfqK+ZYy
9dvYNOuQekkpAQMUxkM/qGMAzJqF5fgjO4+g/CFfPKxgKWh9jrjWsmgpMfd8p1H3
7GnWmNoUHWTRJVmYgy9kcg26Umpbl7BQiD+sg21lvn7sh4PwNPHSP5jGAwGmXi4X
I95up+FUmugKNaWXt4NRjyHxDdBuP3kjlt1P7caHmVK3jnI4BUotfr2/gZjMZ1zM
6+4kJR1uG4eA1DAac6yjZfrukW2bzcu9awp2Jr/yNN2jCCQIqp6stlG9Y8Ylbwpw
mileRO4A06dxP9Lv5lFNF0oEDBGtp6eNpJgd4+sitNeYuLKqeQsTnBfGpb/zQQNw
UUgBUgmlFebqKh7a6rV1a1o7DXgyT4V0HN1gsIlpbAvmwOb94QtNduJbaMN4aBMT
72wfn+OLrVidoESxUUIOXRdieNP7xYl7BmSw5kFgj0TibCrtIcMjCaChcfdJKBGP
RAH+Qys74uRMvAbVZII5M2ECtneIc718foVWodMHpI1d2SipVm3rPqM7OdTvvNDW
12OD8smlSffFuXuPzJ+fKltY9UD9/bz/vQ4heqCE2lwgYK6WU6iRfb1RNAHEbBsQ
8SGjRLNXbOHXEN3H9/KJ3Gu96L5DzIJ/h3P7dGugBuy3DI5v3wtlcD6mmPei8/ag
Qwa+9VNtegOoLzNHehIrG7K06zjUreUlKimEW5wzcm1JIiaAoj5288DSd80N0xXC
VfGYd14TMoVvcBsa/8nMYq3kJAr/tNxBRrlP22U9EezKOKl8cZSWHbdqbbWFOH5H
UQ3f9My1Nm1Eq1BqAAZmkC/wUEItcn7hsxhFKxrQnWfobWpdoZbEVEU/A2fv6ENu
eyWQcMaPF7eO6x13ydZH9YPizCROXeT6I3eombtoQC8qsVQ4198BTTawShBe3bMw
wtkX2j3zZx0YYmrO4nLOJZUAwLlN46qNe63BjmeGaf3HIB0gfo8B6fIuIYfnhftt
NQqe3kiHhvpUBsT/7IxmzSU7pzMwc/WSwAOTj6XdbrtbPMHpernI7zlag2JowuoM
dMpbrSr5PhWVVylG8/LqW4xSQcLuokpuU9DhH1ieOWEQ16OG50Y3gaAVCx5e259I
8/X+oXHfVDbFq9qinl8McZXi4NmIGgpLK9s4LcBOsOSW94mRPIs0TsbbOLs+zhvg
rGqHcOijifuioBIcv0ZDgq1luVt9FenqPpW6C2nElqo3LHb2CUT+OU5nMveQtLDv
fgNB8OKLPV8+OmqnOukut7QX//EfQO8qZNDN2/SVD8Yt1/IE5M+xQRiRkBxJF69C
w4Qxa0r5lkMODNwEbHwyohysoOLgGcEiI94xsb0FNIQPyV+I00K2fzpeC7+JzcOs
UNUCDgnZQOfUTk+50TrnBYTtvV8yBEDx1InVdabSwoZ8E4pszQo2jPr8CFaAnOwr
K6nnaFRdq7QAMF7/sqRB+9Q7FBOMUwZAyusjo+mh70bXMYSQyHf2wUgDu52zp6wA
Xc44mZNHMT4QSbTuegGrQwja9OuoJaukA+WQDv8ix1Zm48Y3yxoVhoDkYL2rgzuG
6EVLcEda3FWQdNWrVO1XO3XEr68WrnDN2eoO+7VUxEbPfKcD37gNUMuWhxoINjE/
GCznKPIn9XBM3AXOy1C0jSg2N6mZJAic4wtkrigCfMo5g7bqWJwZ5UuScVlK/4tT
x1g9/IGZ5uJsmWIKxr6RG6R+Tszvtd4T1CWkFXp2mG7LVsOamlf3fWQQGbwV/goS
c/O4qCRAM0D0Zr0wAIJh53pa8Ea+NWP0BUqBITbdhjkxxwEwSgNTnYZbjhnwfjTL
qaRW3fW5DLD7olFAzl8O1ZeowdF0p3KHB8ZFvUuja+jZMH0umgyaH0hTLR7eC210
`protect END_PROTECTED